`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fFqvKFp58Fh3Y178fi0vWZ6tepY/67QiS/LBcxeFE5qVhSzQqpFvg1gZJVCdiqlk
RR8UrZCYv5yO6KVkwulLmeoR9Eyy5LnSgHx1c91/ta2TnjIYHqjtm1T6KnV3PpD0
IeuznTZ3Zgxwz91vI8ekS6J3CkzPk17wA1XxUjJY+A7uqmclQAQj4jleav/MPIuc
6jeb3VQdYMXJcb9l3tBL295k4f5bfBWIzyqRZJEk8lJ2XpuTzT1ciXuUaQpO3wqG
Z02xzDzdEnQg7YAxJmhHCrDHqYq2lFc+eeYbA/EBvpa3fP/weby13tH8CEPLnjYr
/5ZzbkansAbSh3H+1oguksyzCI5/d70+f8f01ElAgjXoXCm8ao/hQUF0R9SM8849
LWRpka/tTCVtg6On7ions/6JuQ6WVVhsti1qC15foxWpr2VBAnOp50osqAOPyI8y
`protect END_PROTECTED
