`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTnkO2RpmJCMaHDDHB2mfVgpCuvOWkIjL7UUSnK2ivnjf1eQLDS7CNZTMKUijy/J
udLM7u1VYawRMzT2JVYxO7/vnJY9Ww3xZ+FegA6YMGygS6cHeWSO/Ou4BA098cDv
AS6agINhUDyMCm7Utdhyvo4GKG83ZgDYUDYji1zMXfieL5Bq37nXZAqmV23MPx1h
5pzlBAcME5LGY0Y0qa8gPVukkX5DuSnjfiEjarIDbBBK6dkkyIpXGcRGOiW/heIn
pDazCYEy0ZBM/m1xLMmws4sH58zLFyAXZsmKO/NefhXL95v0rJJIY7gG7mHXXDIg
Ixj15TaOcEfQWkeFhlw/x60LbXU6nVetqNITvcdtu0tENiPDC6IOZG/er7/OCcAc
ZZ+S2dPIb7kVDWv263qIUAmKgdD61si5M2uWXJ9QaPA=
`protect END_PROTECTED
