`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZPl+/zzrA2DETIEKjSdcH78SntJOrlRxa1FwzpbhzKC2kyuzu9xPdLAYjbxxse/5
Jf2KHuWcfn+6ae0C1oGCwrwZrSX0/Mg1FPCg85r2nFguNT6vKigPMowBl3kLV8hW
m/BREs1AhObc3BXA523Dp4KXNC4VMxFtaxYtOvk8CMQnrf2WF1nohQHTZi8Xvikd
nXPJIofQIfiJj+VaZBxu31NAtiC09FU9tiPdjC23vZQCZMv4IGaQ3s5wei03rvOu
sFlq7T1deMvpAs2DhkYXDlMUQkcw/9ahg3OLqKdLfJ8Qa4uqgKQXi6AZCBCKzABd
ym+pUNLF/xiJx49TDdAcky3+qg+BqVtvh+T+poeaaDcouj9a1zHttvWdkao/VXoX
uGTDo6sCi9OZi9WrbHc01OvTLAH6Yt3lPRtuq70N8k1gu6QtDsH1UBzOwD9M9nCH
FZSvx3teFRVHBUnhYEAL+vkNRSZ1qBHCMJOGb/9AJs8toO940SNRFkzq7f4oaZUa
7Z60jQuFTgrRPsoKKobfS2P0kvki99YcnyevNpCe00/N0jOMocf/xuhlsSEaykR0
W+T6YIoYeU6g0MGdO3VQ/g==
`protect END_PROTECTED
