`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWJGACRAoyaRpXwSw/CaVS9cxBB4uetuLGlWX7CimIkuzSMgYQwCDbDyL0VU3P47
w+AV7IOtRiYnqzRp4MO0E+yFRN8M0fI+R1+Bfxghb6gTf+YhQ2TQPmJ0i3V5dgDJ
/NXtHROTo9LHux0FPeweBJPTOZuGhY6rIvtwh04Rx7PlB1/Sx7gTBBXkIKuFdXuY
IZ8AMOm13pyBIWb70KOsApi1ojdl7ng6PsKrdvWqIfi1KS0X2zm6mqgaeAGUdgVE
`protect END_PROTECTED
