`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQ7urR18lLrixsN2pet18XD/gcdU6Myd98r93M/sniwqFPu3D8QMZoSVo8EcWaUI
Cbpgso3SawD7+ls2XSJhV14ZY5qaL3lp7pvKSXdCNc62Z4UeUOubYFwRQah/X5b2
HvYK3tSEh4wmBvTDcykGGTWe1nNlHXorpR08y0qTeBBA+ekqBiPzaNKsKte7T0QE
vIJ/76JZ614bwByfBXjlSRqvInwoNT6xMZ9niy82wwP1yiv6xB4balRWiiUVuvFc
tuPPzDoSq1OeQuk6q5EhHSS4HM1mB1xVXnLPusoy5lWlw4Ed6R/JA6Hz39lU3FcA
aOaPd9waHNPRADWy0pi91muYVhr7KEJj90klpYKDgL/yVHL4mMwgs2lN/5kINS1H
uaxOrg4mcIOLdhBUGSLIlFL4Bl8M54gcXAhGwAb7GMmBS1G9d8enLvdfmW2t79rp
feT9yK9bWY8t3944WFEtjA5zAvMEnSL7A31x0fTfegSMq1hfYJfvJ5Vph98asyAC
mtPUCZFMvFOzeuauFWjAA7FaX/HQyVBM/bE20M16+XxVIkjgwcW2bBGK0B2WmGj7
CvPzzjYCmCmaudw3zsP1UH23MeAugnZvlURKJSL8IKCX+zfCkjJDG4xsgjk2BoWF
7ypojvW7glUVjE3n+D0f3LOPmDaRJzCovXlU9k+hFhmyGpN2BbI/ZDl1jdAcYLuO
2kCVr7eVVsv1vSzjpC67W85YmePb0bf1UEUfIHLBN96T/DaMvyrPoWv3VXcGrKSj
rHrJZpF8yHG5HhcT9Eq6MPaTYLNByJ+eF7H84fHXfMeOX7ixVwwwhdwANGnVul3H
4xsOLTbxH7NDD34Wz2wm7mdqz6iSVWa09SFdu3rGv1w56WcPos0fydTAOeRQgAOG
8Gwa+CHYyNugUculB+igMzWu6segW5nzP3rjH0TzAML0xh+igKnYWfSKY9PJAdi/
SGG46WTVnfo+SOs8Yw3JO4DRGgf8yhzTof7muzvEB/hU2mye77ae0Vvmi/zPkVmX
YQImU0gDGqIJM6AuURiwrH+Db/aP/OjrzT+rTRSU2q4T2Sc3Qfb1iu3bl407fh+Z
NPGAykSMYQGfEJNI4Rg1sDuRxsEOe79MgHLbCvSAYzqScrOS2heI1A9gc8DXadSB
sLRrbUMrlD8ZfAyuuGetaY8nuEZnYtDGMCQKVdcfGAPkhqt7Lq0M8Id2lUSuQAeK
7pbuttuZZxpWWfxDUNmjKqWr9UXpLpq20bGov8FdKzmnV0d0USKD7APQUStfJtgC
HxrI+qtP9GGY1OiZHKW4eOtV+jHrmQ7UyJS/3zn/1tdkn4Mxx/TreZ5WtIB4HOVH
LbdXdpHyp++9aPkcy/5RhNYm8mI3GzpbJ7w3IhxXWWsJzVwFWcMCzGZSfDOqCPFB
5hnBYocxHmt4Kqrc3mLJodQxNyCuuIlle8OvXjbKti0zeLrBxjluUKLhWdh6S3E+
FXYmkUOKUn1EGz+ctfUtMqzK2kdtZmxFmFovyOsEAiehQkJxLeKVyQNRveuyxeUK
SfzeShwta3jophRJ3KmnShISfurFjxa3c9nSNX55QeFVY7EFG5VncTvIGIXXKQ6d
rl83TITReOjvCbetyqHYRyK+fhVZzDAQeT+lDFMmZBnLqM78vW67C4QlZ1byup68
UL0dldqvtNPrJntKopfCu69+5vuG6JiibzkAk+BL0mG+EJmSayqUMu9KwZEe8Pdt
2rqPOF5Xjd4T4dO6vI3iRxvSUU9RW3PstkuXUO/OVBvQZMIbsSwBbznazLwqibmS
26EnG0INXwsjbX9q/P4LUwdVBPB1KDO/x8o5hxR7K0nONHJF7yoFO1tvgsxwfRdv
wTfnAmM95EHuB/mno3JFNWwsZedNIv5rqjFAyjg60D2jfRadfanZJuwPT/2M5IRz
2VGQYcXxE8LoqOVNKpxWzTPuVzw9iSCQH49hDArxK7cX0uIx9yAveOT5S+k/xEyY
lr9TJzwWaeJptc6hSaZyrtCgzCalZUQjbmhMNsbi+mDyRyYlMOTIItq1diCfByPZ
R3AGzSgzX3o+gu4Y6jR3q/IkZY2Nvcpx8NVLdpYZGCPBp9x2q//0aFYJWpFb07bO
DATANd/hzDWuqqZyhywn9LLcBQpEpzQRE0afRIK02rx4W7NC5/saROfv8qDv3nMR
2OMEbU0Qd0Nhy3DKnvNEtJ2VpATYtw7wQPLWJdQ4FGxQF2B/x1tA6GVJ0aohllRU
q3g2ZvAefSroe6ydcIXoIbWY2CSw87kSc2b8bTt03Cf4Iti1mJq4Wy5o/cmtoqYk
wPRAHAPsyIn5RsAzNbR7uGYgD6PvzSfdFTm0SZlGh3JoA3gZdKytRGASlMSk4v/R
ZhTW8/mr0Kaqy84N2+8DadmVooBBVeP7rPfGLoEC6jKXZ8tLnVNuS9rptS0CAIXG
v3w5phFJAK0PF4q8x+f/3pxjF+fSWdP2/0cVVmu909eVwdP9Hj4a4AQR5hdFryxx
NLQEpj30UsJQ9vLUtVAE0ynT5bIjwPkTIkPR2VnQ61830yJxRUJQdND3CJirBavz
8vyvax6eDRI+28GpHor5h/u69RtmSLAsF+tBGIOfZ5E2tGJLELGJU7NAmvNyIstW
2GG/oSGOw5Jub6OlYktccF3KWaz+ROubN5k4ZGRcWaz6Wjk5MFa8G25teYUXkSh2
Dj9XH6FGYH6JpLNCrriF/XvzIV7R4Dnjz8u5zhsoK/0EeD7WSKW3Ukc6hqum5HZi
Bna3/hlvPvzsoHXxVSq1d27Ihfpd2RHqcxRn7tfsbgf9uAK+5jtnno3HoX7UkGMa
Ez1vuI3QoS/hd+Hte+I4DRUQyF1hChBH7z8LWd2VQD+Z6wWW20CK494m6mWDDoww
AOJw6cwvqakqhis8WZ1Gxis3Bv1JWvJNFixAB0mIAIBvVvtGPnBhGD/0aIHowtqy
tIi3EcUEtDuoYH4tQ8nCmRT9f2L5bkXH2W13udh4FqVjQv2rYqHClBkZ/WPLkEWm
FT5TltAZ29W2x3Mk3Br906d+voXDp/sRmP1wK/MbE4tqSCU1lamBWoDBHHeSbpUd
iyvi2dCEA+FWSMvWYeUWGIWAgtUb6R6+OUfs2RD/mo/Cs+f8nU5sgFiHUNuIozn6
rS882eOW+ugy+SAbmXwAzr+EZFT7mR6+pLYS9c1fvDxEqz9gnawKvWxpO8gZnnBy
hYbHwKw7Mi8wIvAo292noWaoQGFPilzZ3N4gvN37jyQ9RF3C4JIO7XE0wpXATTAz
iXQWNjJN2qRRboyfJcHwSCrak7KoBNzeBsX3AGMtWm4IIBRHSZY7dtVWMqbck1xL
OI2NcahpwEdDUyGy7WD6SXgLHE6j5GAFZO4eRwsE5K5PCBAeKjO7buTuNwqv4Xvw
E88ouF7JqLRqVkO6kswlj2Ap4fvJ+anGRIK/EF0SuXUsy0iSVH/ZQskueOckxfRP
Jpf10R6bNEdRZj0en0kB6p57801sMm1O78S9Gsp/MY2boh8rV8pI2LM4bDbiN5s8
mw8XbIwflmxa0GHzGqRuHfGmoZFwn4V3dSByW1g6RSwTDoU9oGwkhmQ56CFaDBZN
LEmayJdN0Cc9GkM29CLWXuQs/9Bw2n/nKz1x6qxcJpqaxXvZUFMNUAlueBhl3Lz0
2UIWMm9UvQDcD6V7GjTbliH8jwff+q18UZBJukOMJLfeqQPt/fcPp81izu+GXkV7
lytS5R8glLTXQowgdvxDp0j2WRNIa1B68f3KB27CR0rNyjFL962vyljqMnf2eXvd
+qkX03iyENAwtoiRszWN0mukzlGZdMfLNNdVcgQ1llQRQTCqlFlNLwbCuuLSE955
534Dni74AN/qmWeFdidZ2nufbuMD+gMNn5QTsbrx8jAZYVyLEj5IrTwaULGq7yyt
XQ/mLmnNW5teWLnLXW0V4FC1SB8X0Kf9Pw/XQTrrIiPO6e3K96noe07Of5vYBzJ+
T2zb9GoLtaiRFhk2e19lgt2/1AF2L8n3nbm4fOCwNtlzZEo3paneUlmhQD1XLq+8
j5bm3AdtOs3G2765Yp23jiRoUalLbKubmXq9mCYn0C0GZd6ywi1F9ARLzg9w/xXf
qlDAotfDJKjUNeENlRvwYCbU05ocxIILD9wq6lxopfOQi/5TJxGPNb7daYX9gIA6
NC/l6eNfUczTk7fms9dyNViLtN0rHkRTJb/KTtHJkHXvy9842mgN4FUcP3RzdEY3
y68xqWYfw1hvAH8e2/B5gYGJZK4SGk4GnGWVa1Jn7JFqKdD5fBtFxciTAfrWLjSr
w7abYpQBKx6kw62Ovm7jtHl5K0oJ7AfbCRITmoFemhrgbNJ6PUkda4IQ/oId4aYM
GRX7+7KXI1Y3hrIKh/W2LGubJQygnHdCjs0M5I87O+z7uR3gL8HIoGqEJPnKSSJD
wLJxqL4MOe4/pHwiw0B9hVKswm6Ph6/Qf8ZR/MKhrkvhncAY0wVNYapMnuD6HCiE
U6Jrhotf9RhVQSCg2VBy8MfiFQ8JrzmtPBywekCS62ojHCUZecN62ysXzZW2IvkK
lbus/WMLkkL1Ewvdz+fI8J40yvGr/M58UKw2s5uV8qp1fAH7MYqqEu0Rd9i+L/e2
ffesPLiO+Bo4iAfx/iRLPaUEkihRcjN1YFSbFXeDdQDrOKA6FHo9jUT7JtlVvo73
I/7KtbcyRhWNTe3rzV8hvC5qo1/BIruO7RZ+xTiUxObd3bAlaxQjlDFdW/VzbLfr
MyBbgnqNRKbfaZShhexkq6R6U21bhGeQEVwbr1oCzbBHaQgPonFjhnuyRTJICK//
mw9mVY+jwmOsDL7UDTsZ69EW9/EQMWqRTKJxkkvCf5+Ny2r5z1/NfuH8avlxYyOJ
kYTWVBcq/wqwmQ171hDUvrLbbZH3cCWpUJepwfjDE5A1Fa+OdcbJ2BpzWOnN+5CA
nLGzQFKQDlkBDeSi86ygls20pVsdnX4tQZjA1NdO2+8O1D7Woa5QEkMv51JZfmME
1Ye6/UVqH05f9HX6fM25J95xtTALzSVuZWIU3JgHSDNznsIwzkrTIzkv6ndePbdx
/KIQ/rKIoCsOqIwLf50ppzd8o9oclKJKR5vLlEdu83aD+RJPPZY5xOfirMBNJcjp
vliwqrup2Lzo3+HtJCLDPcX8Qt60moCYXbnJHFsmr7y8435IkalRSd3iPis8HgRm
vigukHX9vB0RFOYGohOVdIQ6nAYnf3EOWWoH8eALzGuTtvy3cgHQP7MNLVVFM8wi
x/J4sa6m1jnRoLByrIuUozKC2ZOztzLRL+k9wppYduibhGlhp/I9cpfjSq6G0Tln
JjwJNnV3XiKpfCjaiR4OR6mIBR8i1srmXDs3OMjfkJND749tBCFK0GcTGvF2Mtnl
YOzRVgbU/MPiAcMAJAucgzGLcqCfK1sGuYbVOqcwXjIhzb8l41zLH8xIfB/yt8/d
RBS/i1hbWIzJzw4FjcGPQEU1qfhww1WvIVYk1CX6RZQFTLTq2qeiE5i+7rb4r6k3
xEg3kb2BbuTvCDLmLmVz7KPuCf8BWZMk6lNueKmTX7L31ZrnY3KGjrBxLsuuGdbo
dtaZCfEIVJ4/gxYCumaRobQVYxDmn1TgxM15zvxPfs19H4poaYZ+H9drli3Rr0Zs
UP9iEWF50iWfikhYIrYIX3W9W/rG7zAF0z8pRVagjo7mfYSnLkDM+IswP4wtc+k/
FNtTubjSpZXbm7qhUnxRNUoTEqLe9WEapxnBgGSMwvWGuDLUWPFXedunNQf+J0G5
z1+wEz86uZ+sD6ja9wf9ow==
`protect END_PROTECTED
