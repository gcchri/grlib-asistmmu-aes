`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yA6/WwWYvon+ervDJXYfsIZ9nMCX7sSdqPVdCWaSFBXbTwfJVb7E8tgDe2iCqpIe
gDbgZPinPizHfwF5yqCkvylYLJBLHeqqJpRO1PFlKfDpnat5dRt4xl8dhd0OjfPz
PXpmNZ6krQd5hrQFaRn8hxCUi6NvNqX42GiYxYpH+fbnu2CIiCHYbwnnrpmX7W26
qfQIbSNiCFuKTm19FUFpL4IM9x+ABqH1lvkVhQddUACZ/S/LV6IXZURVj8S4RstU
r0NgmlZv1r9Hy8VHY/NvKCgIcgUJ/XWC7H1vaiiPlZ+07y+ed5DcepOt2aUbAUCI
FdYWTFuK8dNE9s5d41EKjA==
`protect END_PROTECTED
