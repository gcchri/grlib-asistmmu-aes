`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/nvZnVixU5dH+HJCzkzzjfqFqFu+TkhaeK4gap9nGKzNRHULW3epOU2TAl6igkRn
oyCkJuFuDPpqT/tjlmi3UxeEeTCDx433ZKQflg2rFfbl5lsm2PxzZyanG5zKioF4
tAdwQ1DOvPOkld7v97xz6sRrKKvWlmsHcBNNCzJHqCRD/8t5kApmUv6EfIoxLRKr
XVzpz156lWrk+jT7Ia66E3kFNtBhqEfpPqKq5fFo00gSbM/Y2VVQySXpt6ikHfPl
kDVtt2Dnnot6ZvIZ1yE6ekjnblw7crooSug0GJVpM7CrPfWZBfKufL+0aDzU5N4s
d0AuKx8+DHHWj89o+SzOttRBnLOTVyTU/upE+Ng046qBceyxEWO9PGMxM4YwovlC
`protect END_PROTECTED
