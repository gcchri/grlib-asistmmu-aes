`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rN2y0Ara1diWHxPyx+HcTsm9+lzyEOUlZ/YQamki/WzzAie8mVf/xRwI3EPC4bYc
GjtDJ+f/ddxxYG2xxZ5UVrHYocd63iZmtMGr/CYPQUN/tJA7X2AueHzXfAkgOVhg
jnaTROq/g1Vp2wVb+IjklY47800AHPF57LcIHUPvI5glhQfAGfSE4t6fwRkmNZ6r
FqHE4SCicndIPR3iRL5hnm9SysYr7YNgPndd9U5jLvK4jT9vZyxY68pi9+gaRXef
NYH8RNdS1rhVJio9AzD8BfF60A/vLlil5R4zkZa0zFL5YWdr/0AUrtpJVfmEVtVg
RO0FqLD9YaWPqlWhuYbLKkhKr6kM/RGHnaz+UWiOYSbU4+qKn7s+Ws+HYHzk6Bwf
AIA7SrvGXGkRd1UB32XBQanxmEURI0a+W1IKYyAFITf7rLeXmuAe/K5hYpK+vMLt
jTzhEFUWoAmEnhLjnJLkFGs7KVvRtehpEDRIouV1CwQZQdsthQz2gNWRDkPjRJbb
zHQJEsVp5Iv6JFQJN0ubSDBp8fWekSfIWttTW5b6bO+urWZu/TCyW1FEItgIp+Yo
RP+ZqYQbKDWYFVz9Z1RXN0KMRNLb3GpEBtMOrFVevAWW1StCW8TLUkTYS7eWqgnq
6JXYNI8EeuvVmcqD4OUWJMoIRj811lBSC3vCPqz1yl6LdYfbrSZc+lopV5OYmK3/
2zTQWA7zlRbWM0+YTsCvbqCKwoJD54zwdS1/BC3AcEQojzKpmYMgaMDBv89pNeTv
y1ARuJwWBP9X3/6TmW/uxFsZENg5QZs0tYJ/HpEQ32A=
`protect END_PROTECTED
