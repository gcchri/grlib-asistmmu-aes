`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Dr2CeLOZIbbgiM1QFSVnV2/RDc+teCrvcDDXpr7xj3twBUMVk5Xlhg6wnLlN8dM
2IJnGXO6MXerlYldEBYgEpe0j7hMebVvGAkb4C9Ks/psTNqF4zwIjxy/y+6iyhLV
KqhQfEut85/2ble3/XTjJLXFKzUwKLg/oyhqzi6ai2TfkxnDOhfzH4jpLLHu4PyX
QEIsZxP2HN2mRcXOqnhVXAoAlpDZrUsFQOpaRCRLIE0vNNJL+JCtiBfFCn0Kzngx
Z2UlrC/84+o9VvgpCaU0CICP5gmOXPgzoqCiX7wyuiqB0yzkc90vSX339eb2mXRw
/pqXnKRSnRNhELEH9TMWXnSyBI9fjC7dOD6Fu+xOWG9hTE+nW9DInIRjgQJ94xih
aB7JnN104NPYy0kAyaptarhuFtTrDSj5pVCah/0MQcnq48JAFFiwAg2yWpsdqCmi
9i0Gz9pbnlC9beQnc6oCBnhR3rpvKxG5yvJXEAyvHTCmg6P7y6Et8OmxuP18V6w6
ahvNThBpdhAbEa9Uu25vhXnpsQwy7riV7ObrkfapeQggS1OW+/0W5uDgPC5EF6oJ
WzHqvljA4CA1c7ijq95HULZyE25ZEqqh1enXFIv29oQ=
`protect END_PROTECTED
