`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/zK2F9M1ioKU8qXYeY0BrzTWoEOY3Pbvzoz3zIGACdeIq6stU3JObf42sd5Lwg3
bN7qPKUFW4wzm834NkNWaNjbrBdik2kw4/GBxTWSD2fC1o5rAQEMWkBT1k8g+crx
Uw6I3PyfHsuVgV2rvN/pENoMFgAss6Lj2+eoB+2HcSS/4cUwC8osGVmGA1cYg6Xy
tLEcr7ob/Y3TBtLql6Eij9mT7NdB7z7lkqNm37K0396utdCpFR6VafpcgR5cTDXn
rSuAFLnMYivbhLSDAMVQa5YuLWtufiWsXsKbQoksEY8wv9ZjygoCIkS+VIQYwLdi
wb7SAlO1IYiDqnrgYsDkl4t44T/UziXqglyWlOoJFzWpfqn+Hb0voUsFk3jsH7Sc
DZqIcgeWcvSzw2iijIwdpfujWDMWgi6sbwjk1hOfCR9MBZKHIVOSZ7Ej4oE2XcW/
J2LtKvyLfrdozgujSv2p6zkpCZUZT9Vo2I5+w7u9257PHAyBtoj9NrzCbisPj70P
+y9IGbhEEiO5YKzIn8xR/+M5wnKHjyNMl5kL9+Sp+EBnzL4YjL7A0TVerMhL7n3v
2DbOBxPYZDlrmf++7GtDs5mH3UTrK8QTSgVw30HQ0f4kAcdxiSmYEYPyQjtRO5Wn
U9mfcGm0crAu9sv3seG0tHKbqjRi9VArJ2s4mU4gYnmuUNqP5Gvd27kwHIU1wv4h
/W5UGrokcL4C6u+Uc9TcxgEc94llK3AWXB2twfghIYQWGKbBwg2f0yrexQeAFf4U
kUiDYBP5BU4HuzHk7/+bBA==
`protect END_PROTECTED
