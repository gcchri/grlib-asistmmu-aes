`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gkHz+ngpo3r9iZhldcJlTw9GFQDA/e8c9R4COUVJP6T1nQhRBP8zm7reJfujxZLw
ktC3qJ564I9rVGbk9InLzSR0fBByyL5Gnw7uEc5l+jwppJWHKmwk5VxaBSJdNpSx
zGFIaecytJPrLwbwMCaGLbD8pAA/so8XO+fnyC6AK+0hGOPfuVOVMxZO80UEptjO
BzeoGwx/k9BS5gzji8MP+a+KD5vPuF03tblNZ4SpV7JBFOc3+FPaRk8BT5op6FAC
2pmmzsrQRANso8tqmtn3Wj4AtkTMij6zWYk1wEvRXXEdBcfcXJz6urmjMQi1tKxQ
S0rnutKX+xmZcsLPotCZw3iFBveCeabNX9o9Y0GuvqoIumLvh7oqcjw8/J+9IWXn
5bhanxfSZVt2w2UHVcnnq7fQy+lpJNigeBUrn9/nXkaPpoL8AmS6E5omheKapJ6W
rOy1h1k768QpXCddRbzCJiEoVTFqbHjAXcZfjUUCqrw=
`protect END_PROTECTED
