`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlkmslcwuGT4djNtWMrYkZuH4aqBi63p7Jn4fwAdpn0gglA99I1koSER2pmo5piT
lIm0kp4a9uq+DKxH7TBPZL+7qdTdrvSPMP38gch9NgcCS3CbvC4/UAL+iKj+85h1
GQviM/fNJbKPmuhBkyyUeBNuwFxqcPculsisd0OBpBjqhjAa1qltywagCAnhQ1a/
mh0HpVQUKv/7LpQZV2c4isN1qSVI+0zjqUT+izKPzCsbMPaMHiqG0N23JSKqZ4oo
ocR12vjHpCk2D0Ia2Nt80891LFUzMf5zJL0+gbSKD6w=
`protect END_PROTECTED
