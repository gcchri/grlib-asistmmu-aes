`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Cq2Y6Cwa/v/zkIQFFYD614WXzbjCPQ9R9iKw/m2GwtjhoJ7/nqweNwDjIj9Z7gb
fcHUELxW7VtfU0AGGeVnKqRPYWy+F/NYIgCeaflZG4yERAemGOKLTyNYFuB6TkDc
OLzk3D0HY3FoEt67g4Mqk84k3G19bU+BG5cY0xy+bYdNTKHlMvUgvbc58oZPEbuA
+FpXoEt1dnk0lZGuriTSv08RiNJP3QikEsRlKQN62rE7zvZarofGhgVqbdmPjMIR
iQqXJPySBKyzUrFJtq7KeZL5vzGFwk6cOTg0PAM7b10TYI64QGUesKpq2WvMmPLn
Zk4o/Kef3qy2rEW7xQ0AS5P/GMbTgWprDq8AGTyjQOnZkQwlUfnkXuy9lyOK6Hyq
zw144W3TBHcK0D7xLlZEryQcHsyvMj0Jj75+kqIJ2WSpxkdNZxw2IfbhueHC4aJh
WtuGaJ3El/BryLeg0fiNSSFke1AvKFL8jcQqYT9jzYCrybpBE7TodQuoFbQDMDx6
45r7zdcEUIr/HbExbpaZn/2svGtXoqpEghRxJhcTJ3D7EjdsExJx6d/K7chq44vi
ZSUJvrJs5O5MdAKLZHrbLnwZzRKDjWP171GeDnvr0nQ=
`protect END_PROTECTED
