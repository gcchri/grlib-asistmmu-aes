`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gvnf9YmjCWCc5xW3sj9eibepsCakgWzBy2PsM5aHzHH7qmp3LsPjoLmIvO7PwDQg
WPQ9ZU9dC3J71CGrROSIgKD7+wh0biSacukG7ISITz2q8sqGU71g8fPdgbaucfWl
HzrjgtLMZkrMuFQocavW8oXXrK9BQauG2IyD72BOjFo0nY63Eq0bIKxu6cjTurjk
lUQsZV1LAU+bHpz4/StX0xGGjNcMgEtiSyJ5ehiMixFuHOXwptmPsNwnFuVeyd0L
tlyU9V6qzh2x2KLjVsn57Oa6uSDWOM4v3ldOIxz15PAmvrE5uWnONLx7iiOsH7N6
NB2MYOaN6lahreO3YMQnnq6tl8ud5WW2ndse7mrIeFWQQjNkNTZC2fC+/VCv/8wc
ntJh2ub2V6HhDnzmMQesWdvhIBxAvQetxbEbIdMtZ9hD2CXToeS3px7/3vRt98Qk
5LHQvDdU8y4t8c/bY1YPYlY+k0lFFrvprThc/GPjUOpoC5DFXJy22ueGV0u+3qEG
aLvAA04PpddYfTVAYVnPs9Oq10cFbzCu8QEC4gr1DXcuN2c4lonXtQM7wb3uaKOQ
`protect END_PROTECTED
