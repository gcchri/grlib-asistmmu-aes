`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kwwDPzIoeHRjewsOtyBb6aUjzZ1slux5GCXS5Si2Nlkt5O1YEJaT66292N1j9IOj
ts983t7cIEvTdQhHMVRAr2b6OVS5XZGVTWH5zz1LmQKW9lmi536JXWEj0EsyN8X+
UaM8LPFve70VrTaqtc9u3xnxOfcyyOo6Ki2pMc75/ikYotWWcyQ71WsYPtldDPN/
zkJ0oSNg33sEbus8l8btcdwuQZJng0YwXBd0mkFEPYz0mb6WyP8qfUepXnoQ57DY
1lU3KAPwvOI0vGmzNYgafhQBcUBog/CNULCrCEEt6IROwnZ9gqQzEI9UgAstZzoq
G/WRcUsxZmZKBZtJZZseLQhyWfnr6A33PhxzCmeAXRfTiU7H2MtoMf4q816SQT8d
daZp8l/eK+VylezTYD7pgvVa1y64nc51mCVvTOR9vThMotBEGchQblUph/msZNWf
M4JvmkUFpfz/8nRU5jWgdeXB/Zqa/5rMKZFLT3dAj2ADFKRN5filIhUQSNysXcmz
YY3yU+O9zKTPwRAPN6Z19wxuLXJinlNTxxodK0R7JWPEevt86445/M6tPBOz2gSn
sPRl0xBgdMQQ5oiPZb5/VvTfANhWhNOMJ0Wh7svdb71AXoUw1YgQVOL5Y+qCvAtL
LCFJaDLrlT6R5gpVGouMEQ==
`protect END_PROTECTED
