`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qY2MFtXvIERn4x4f0uJunNaQx6YMjrmAdEF2P/1JHWqgP1IaWEBWv1PhD5UKptHQ
6Ih/TAB+muV8EkRjI2OBp//4Ydz+rWFwu5tFZImH8GSh8ZHgCgoiuxlZHd8bZiGN
lwUIvD3IBa9gHkn7e7PxzCf4ct+Tbh5drZLrBDhIHwNS0oX/nQh6B5EW3HW3V7Ux
PxOy0uIwRPwIW+/n0edlX16t+8AbVMHFrxVFlHNEYifuSlgMhtX75OQQVQHiLFzV
lKPD3PGLCDtSpX3Sagci9OC0EQWq8RpZmVWkg2vuvptc65iRBv7J4geBmykEfG6d
Ip4FaWyEuknGGd91BcXCbsyV2W+ChfIyp8/YZcC1vHUgNXi4GINuSJWKM+8/Jkdk
Kdt63Mjs2ZJsfIEAq504hEL90PPkYsiN3ZC+6COnt+oH0h6LVQOefr54nbX26rTE
L6AbquRo3dgnbHdsgLOuw/uAzdFJ4FjmQ7IY/wLoA61rQu/JnED0H16CgqEbi8oy
rCcCWahtOpSE+usFtjpKAImj43Wmo8ZVcKRnlmnL//UUqXOfl4s5OktB4u5c25va
lOH6X97vt5jXvupthVF2dk4kDlaFGtxk0remAnpnokOxim99ZZCDXZj+vxKjU1UZ
BHADI3DREDKQSxmd45Hsb56W8r59NaRslmL43eox4UAqgA2kkR8JpoP3t1QF50vi
5mNJMnqbNqiXLLNgogQK7y3krzjlxgIg3c0yjKNk02vDD3Eo6r75j3sVr95MnS1o
PXEYjdJsCc8bpWyahuZLxL/rn6QXQXdzK1ZCpLtkAsCevF8d9M061EI+LiZnKwmy
UjpJx45W940OJ814Y8KHg/jyG4I4GUnOJsdOUhOOyhC0ktHqB4wjULuDbMvrPXxo
n1iZDQz08GAgJzz3868OLBPUDJxz8dxIW7GtTos2xumfJsrYzjsohYcPt2ueML6g
rUbWFmMYIWGp+II4RmzkTKc8J0gv5Od0PovuIWHLpBKUsX0GUk0ZZeQXYPZU9tRI
QR7FkoLAh298g9YlJYnOE7Hs+DbIYqISF2KDINqRd7s=
`protect END_PROTECTED
