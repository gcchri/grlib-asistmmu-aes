`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cPiBmPVqujP3h5gS6D561DLO5EJpwQjCablR5E3tLC4h//FN9NFc+vbEWfe2zC4f
+KslcYpFMuCI7dxli5lnXaL01PKYCRr+2cTYQuh0nxXr9WUbNNpdDJhbSmau24J8
MqxxU3t/4u4U4BEK7nHyC12aa7tBxecDmTPEK6IL2Y1QCnj1mT5+6jXT+PZM+RZQ
QtLIIt/7UtlQGIjC/R/R5eHjUpVbtlz4rLpN83dLrKMO/9ABUv70pUJLnYOQN27a
G4Zpn+1Xnebz3Jcjc0S6Wj0gBT0mYisKtbDXAenpnm6yE77+BrYQSFpMjj/SzkKv
fCSVLA437eyz7incsdUCewPblR5b1GvhpRedU2PBAcIqydEj2oECGgHtMrG+Csav
a91SDaeH06jI4Sui93Tn7hE9rlvMxSaRxyPosEO/VI797U5CU+w9ma8xT6dSLgUv
Xa9hp+sPSNlYu4akZ2TIOUAEuYfXYfscfP3ekbn4DYd0i6WFcxOAv5Esp9QyhgvR
`protect END_PROTECTED
