`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HqsSnoEyP/rMlHJSoyhRUfk/m0ITYaKIVCjZ2UUHOpo7sGEZOnM2rwnwfu3D7J5E
fXIld8TxNkD4q9Tjzi9ir7rSp/gfr30GHd/CU8VCaUUtP0V8peBZtbpJRvyQv58V
up0N7t3sZnYlrN3h0EQhaNgitOx/0zwbKu1/4cuP35r3qVmgl5AFrctzpHnMHtXl
c2fqFa5WnUHLXPKTm8jcWd6Avd3juxk++keXa1CkZ+yIyoW0oUaxv7y2eyTVZsY5
ecuk32y0bfKmQS1aZ7ilkoWmtb568GCym+YX9Pkr1lPMzMK9L+12wwOcqHdK+T0E
IKoQmE+0PqBmkKQmRKYs+SlVHVvEJ769zESjFp3da7W8ugERy5BPuQuXTwXEhBU2
3xgEnWbBIPvnz7f8wWdllFWMvjg7JkTNxLXjy/1nLBzLyFXKfI5YgWwvxyAlDeo5
F+qOLHKIw9bMUMrAxO8/+110FYfI35UJ3FdnvCCOTZ9viz8He8QW9y4RUHP5xvgd
MUWPegDJkAm16R1pC/rxtHclgPK9bnLI82oCRB4CuliLxoyC3xmyGqAdbz2c+Lu8
`protect END_PROTECTED
