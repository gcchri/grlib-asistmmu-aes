`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ex2dgBV9+a3RR1MQ4pK7iXw0Nw0G4V3ttAlJv4TydZvtUNBZf9p4lRL45d0RE60G
/1oRRd+dSONG/lgirg6ShF35+khY4wIpRkP9lvPKDWzsIVcLosTtpqVleGFQjQyW
RrnN7lTSp9DmFs41g8nDUvhime3nsL22eI/K09BOAHuGLaOPYZPM3jP3tIs9gpv+
yArbGDB0e9Jf9M0reUYcw9aIeiLw/LyC3OTi3p59Xzp5vNrFOLXIH5Hudn2egMnr
kiaG/pq6c0x8JjEWC1wC8L0KhbF0gUqM7TwqYrRjVVVri4a0wUil8q3mR91y3yDQ
6LionJoPbqUL1vx1FpvWQFkYI5SvXH4vD2W1y9PUslVUjpPCVVi28SmxLgRge+pl
LvHLdErbNisqKCDfoupSr2YVBjWHY0BB0El7ARPYpPD8SRkJbuwrO7BYCJm1JLiX
zEvUzw8NwxPvB6GbYUI91UtnkeG/fkuviXy8EWzbzRmVXstLDa/ktzcfzLbgabNK
xGukTw6QUGM1SxB5/AH1iWckSODV/hiVbqczJP7ETKgNQzGBAX8HFAUS8OVp+lcu
6wKQdcNeFaNxN2fsuDG5Y2PowinpJMDJ0x+DYYHFxrWx8nJO2wfSSGiYv+aMymEQ
F0Op6oDKxySB9E1H83CzP2Z5aC43/UeDoBCdoiMXVFZFR6FUZlP0+KqShyVGtFnX
qy7sp5UX3fWn4rH/AstUHw==
`protect END_PROTECTED
