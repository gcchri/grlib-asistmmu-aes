`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tyXDClaUijzQ6sE2PZNd0zQSgZ+RMgF5K5iACLxe/un+K/mGO5XozUz0vBW/f0/g
AF6ErDFDu0R7OrEzNfJccpSLVR6rgadvbP6F834pGJZtkLCBGRBvEoUs9sLvxqX1
p6M4gvfdEnmY6OeeTV9uhPj1OuMZgHtxLuqV9gIKQkJdIgo1NnYnpzsjCJjUo7Cn
MLB53/8AKStAFJT/nSXXJGSgD15JBXM/8PDgx82kxK6/yYRcX5uAWFJTERMytPQ5
8yqACDf/oNs//pj+ly1WqUm+FdXUOwzvyriszeaJ42BaneCqhxRk7+lC8EIlkEGD
VY0sUX9t6g4LT0L/etC0U2q0UWYUoi8mYpSeJj7tvLI5vvRNTr96h8H4aHdVJP//
N4BqCba9JLcm0MododL7BSARthjPqKX8BItSkQMqTV0fG6b1Co8HKnKwRDBJzYox
TOnL5xnBOHJiUpJlWzaanvdzplDLwE+IbyxxC2hAg22XqzlQInFicCRZp3yghagj
bloBRYM4QwQhWt9j5xXdClufHpzhl2I3SjumG/0pomUQdlihE+4mu0bYsg1bY8ou
2M4fYzktJebEN9T40YA91mkuXVMkRusdSD6VMEDh/EwtSH1B7rMfs2EBYhQKMLnl
NGFsBVtSncUjhKnArppQS2Bg5ZgG9FbI2dXHkU/oLAj1IWYAAjkz067kmAURr8h9
bwfyWUOoGJQb0FO5HFHCCFzi5OonkKHrcrSRdcEUpoDizzw+8c0P93sXmUzIqL7N
SBGOB6MEOTUtJ+Y9s5Z8ZiXkJAyYTvDBPMA+t9eoukRy+hxa2svIM2OhyUWMzfPy
HdGnY/DZVfjUD7Wwjx/oik49qKBXlxnP4LwH7ppqJ2kbdv2KtRuAUseJMs8W8Yx/
hWOrKUTqFrGDx0w3R04djA==
`protect END_PROTECTED
