`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1xQpsCjKQXDZ/zHLpNpZO5bCSqrZfC1auAX4LCokkL0k+5nNUdrqJQUUr7rkp7js
1K/quzwVyndn6rZfARXPbRA5jCOD7XIAqazWqkgfwe3tqVZ5oXACRldBwgqH4/aC
IFC9N1r9bcAyUXdzr42QIHrNIIp4UHcga+EYLocNS5HPYJSbL2kMZbAb9KUt8d8t
NBhb1vmAyfgez9mX28pU6Ev/fuKJaFW+q5drAYw/xkDosKn2oZm2o5DRWTAU8VON
MGDNmE7LxWOUS61x3k9c92/DYauN7v+5M2KtULKnQYgjr3NB/BB9zrmL0a3lmTXP
wpasqt4ZaVlhFWvRK1iTglbKZv4jkLXzaiwgojyJBUN2IViLdw2GBd5qCId9fhJn
r0RzPeG6OfzB9u083r8r546g8y81D7PA8QoYYTq8q8JX5iKFv1E15bFMqJ3ydBMM
jnl+FudZ9xrvhmHKwrnlU+3nfK8p0iXVUxjS8s9DvSuExwBbE5Iy1ycjcKfVrnpU
Hv6BAKzwOED4glkIuflfBne8zyWuQkdOHljvhhGwuWYHWgC80MCH1VB+Vo31DDl8
zt73ReWVfvGOtcZUiLPYftJV6Cz287zPlOjkCmmUcBPAEdHc3iSMvC9nVhBR5kzF
A5fnJTimBdPIXYsMFiBK5UHY1VmAEOGg+Sj+TPvkIK8=
`protect END_PROTECTED
