`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lICsICoWlCD/xMD9Aup1LSLHsJWlq4o2P+wQ4FI0yw619DOADp61EJeoLz9o9X0+
V6pMZy1Z5Vd1hdOKJVqI/l4JXET/W+5Qnz4txm+G+fve6BmM3V97j4ttm7ucyNnm
HApN/jaoI6ZnYe1SkElAg+TwCYOHVvkLWi0ozifH8N0ib5YFx9cUygxopd1jpF2X
gBRJ5NLgamjhcGAkRHwNoyj7FxscJnl7e+aeW9+gRWaL4h4GM0bmr8A9e6ToiMiR
+/AaDJoXSgPvuP9TIKo8NA==
`protect END_PROTECTED
