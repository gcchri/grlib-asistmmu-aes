`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U3mqx4uVbJP34NTm2fb5qQQD7eJEXhGTJY2Gblff5jWTl7JwBWIIFct4EQVcjwn5
nps64Czg8osN1OG7AvdYSx9R+eQJf2jimVR3AO6aRoSDHlvzGUotLok/7nJjPiLV
Y33DEzjxPNa7L9cJFj8BSWfuWPBBRu2LmF3YQrit+Ye9fJkDj8hFvdQK/RCA5Mu6
/nsyEu9Z1K0qRHxBYo94cbRgU7iOvNRHvPrLTf8GR6pZU6PiyqzC10uwxREMY3bV
gGTRq2F0hSJlLknYWEaL/Eevo6eIPlLNF5NgW6ORfAOgVNyx/xpSb1Q5mksWyFWC
gmCmytgRsVi0Shgm3XHo7bjhRZC/9SGE6o4w05MIVf5a46G5BIsYotT/xM2F1Ivl
ySlPV5H+PMeetWGCI0h0rnhkzichZVrp6a4XX0HbA5e8PWJyT/ML6VuhJGjJ36/e
fBeN8cqALqPwfPylXql0hJmq6jP7xW09P1ee8uj96ORLOV2aZO1DpOiW2H8Pa00S
`protect END_PROTECTED
