`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JM5rbxxwhWmFuaohQOBCM7oDSU90ahPZKRXwGVbT/Gk10uegamN1jcCB+pihQYuJ
/xcnE30F8I3Qdr6u0LIEWE/aEMJGrQNqQIZLxqUCvCzLkDsWgcO/NZQJJpea/G8h
I1x6KnybMVWvpmokuJq9nzV0vg4PKVDV0DKY/M0YN7RqzH05PUmThJK71lnuxfIH
2PwPi84kSyTETfgsfk2yCZLvxvYwtjNt0hSbSkv6uKcBruMuALOa11bnW4NtLT7W
1gERWdrfpxkOeNZ7IVfctZSOfHnZg7/ICIuHhS3nHbWi7kfYOAUXt/3DKC/lSMjx
MoCn518qQOlFX5FghcLPt14p+YUWF5jNHeWeMP0ij4Vr+7+MKf6idbUKuAAqCLCY
kLTfPiMwmxtGwolbokKafbVLnPxhC2cIEnZ+jzuezd+0rqo3rKfq1Cf+tc7kCsEn
DDYd1LUkQj1engLyGcW4Ooxzm4/RVILgRtzbtKlUqs/XZ9Kj4lVqlszX0TaxbNfr
9VQjZIbBkEoDyk6GCA8nStJbM/PGWjL+gxZmMQc8vdawK7qBe3KyGC8IlsRfeBFI
6G4OM/ZiLVE6zOuG3U7hA4zJOs5MrbTyXIltk0t7sL2+esoYwFM4h7onDcuPyPG7
NdsCmAeJJRzyhQiNyqtr1Le9WeNHqAcPaYDCIzJgkZ9j7D7qxN2Qke8Op9XbogJe
IDvV2Zjdd2qsiVNHDNZ+HYdy/MaOEdBIMgBYrsuMOucZc9fIFwYMH8F5Q3Q62xlO
tgG852rvxtuN0MNIeFVr2UMK+qXqKG2UE16yvNBxTld/s7IRpoiMQBU4ob9c+gYD
CLRJG0awFqaHV3MfKa3UxlYJaC1xXIWvwsn+SDo1v8lpbCP2voPF9EOrQeRo16Fn
JvBIJiKwtHh7oOspj7soLcXamdBN/GjTeOU7RGTXZK3OLOoaUwTpiynt9zdqWVT9
vwGkrxuCrBeBKOAa4P226G0b1/HXv98qjf0GQsdT9yl1ggv9+WtB1jGksf2kGSVj
lwB0b0bCY+HTYN/aCxKwAQ==
`protect END_PROTECTED
