`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
syXoK+87IG/v7MTTEXfCe32mj6yj2gBgM2/M8cn0mwbCN0q4aI+6kB1ptlwmgzgw
4g17V2m44q1k308/OIRwGteOBoUUgWP7g88yeCxtUxb5CU8vGjvb1U5ljzwpwhm6
PXmb66Sh/xXPwMQYlC/OBCx0qWIPkC3jQWJ2g+cYmM+GEtS9cIkq6bqHTdWf7RmD
i5De972lVeM3JXds18hvoZvl8LISu3scTg561Kst9BniiPocxeHae1Y5sJJgrsDy
`protect END_PROTECTED
