`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hqASFnaajOABId1AahIBxpvU+i/sFs586qYebeFmo+0zbZ0QnlkDZHq+2famLJTm
6WWkGqI69P7/3ugonkwUXebi51axnDMEGoGqMYSu6r2mAm3o60/CVMcDSsY2nlsN
PMP044wvcjbENR6rrlFlCNksvRCF9ZnbV1ceje3oJkOzxTPoaTAGEkExkpPG7O0r
AuttgZtLobOf/AeDfjQZlb+YGtqfsnm03Ajzmt1bQidgo6mgzwZG5VYgn+2mhG+M
bhJYrR3GDxpTJjfyYVVEPvp6kl6VG0YqtzTvmXJnTXKNgU1wTH0gbsQmtfInB0ni
C5jmWWETStKy1Bj4REe8gnSWw3+AEJrtYgjevFjg5EBYR3noC0WZNH1otm6cmAsH
hSUef4B6IngeZD0FQGfFNJWip9nwuaZ4nxSCDD5aIrrX+xBWkp0gPIkE9b0wERQf
DILyyaHaAf2YQGDn2lzJL8uQm8ORNLUUNpw8/s8W7+7b5ijSwlEwFryk6ItvmLiA
x1qP+0s3VsfkV4WTD3GTrCzkZXgGAuvjfJ7E7qPe1N8CPrfJLOTxOWUwldPHtLcq
mo8UaUlkUSTVjpStwbZzlLC6kMwG3NOZAg4tpX/FmN44rjFoj++QCuXfY4xGpL7c
scWGuGC/qgYSCgnuL7nU7NrtIFSg9mWrQk6xzn++A3VVYfgGrNn4+rihb9dq6G7P
tq5LUeDjfU1OnZiCBA0gik0IJKZsUw5lAPR+nzqZRgHTi+2EVn1qCLhol0H3uMPn
EquG6WB17A8nwQTuj9VFN4Q2/bUdmx3xfikShMzD3sn/+1sLri0uGDBgHe3D1mnI
dTz9sPJMC0E3rsAh+fXJoHVZ00NDeuWwo4M3nQ+64/9gGba6+5U00uJPi365j4XT
GTULogYp6lZJ1Bgq94yTUKvAYXn3sHCbZoG0D88EEXTBKjespku+5EOvP8GBHiwq
JUkap3xsvUDC7gW0xFPykkCIJnXsEHGg7sfwGcn+sBfXTHwl7h29w7wYC9eitwqp
ucNlUbZmTlDACCIhk2q0t/YI4KVxDnRRqQzbrG+5CyHRHCOTQNmMgSJOA27vMJpl
xth5WjnyP/+Lmz6md9cXroJpYucJE/h97PHTFk+7naPAqP37hc8ZHQdRg+YUaGVv
tgiW9puTdcF5f5uCirRaoox5WAwpXZOiFn1BYz2/3tx71hwvUYeD5Kjqw6hzGZvY
Ug572QzqNnD4HK96fPbid6j7ZYd/3XvTtKftIsyrwTiqQXFKKh12nm0CJl05znno
jkJhUSCGp9SDRBlwS6rsfCKOk4ykXwO8qRDffAxBhn+8/ZlydfMvOET/8z8Zq+65
MMPibqphrqhxG/Qm+Z0t4BaiUEDkvH52Vv6DjutbeDdl1EOehTOr0nRLkrM2MEt4
8VPogowckVWwekWMpiMSoMcSzddXJZwmK+97YJ7r4f5Wu7pJ+Hf9J5TapyzfYKxv
tu1lE6pRVj1DNrcy1M1N6qtf824qPOeyivOM03xYKSRwFhp930mQ46/9G/uJ0QqK
I7ca9T8TYh8+xHZfP+kwp53LQulgIniufW4twAYr4mRUI5TkVtzTJ5GR2i69G66y
MWzXcq0unZ33Kt3LKaRh93T1cyVUJentJ09Ldwj7OMilueYaIukcN51Wg/zA+glY
`protect END_PROTECTED
