`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMiLxMHxY1LKxHGB6779TweEn96ikX86EoHHOIhT9u8LjFjZq2thdIcDR6QfufdD
SislDC8s3Bp7PPxdHQrj+9pWg5IruEhxweKAuNuTeaq6PUpEyBYyUBg9mTBubvgN
wjWSjOB3bmLx1ZACBzTiB/y0PovOqz2L4igoh8Bd0rUBJfkdwoDmSl1d1e3ZEONS
nPiMX2SsKt4PqP2PRPECpKaB10/TewPU0OzpBuXyStbAmdtHt2pTkYQ0RIsu9qWm
zBcO+WTk2rclRT0TgcqhUyIw3aFPANrjjeLfl5y4r5rGRY/yPO/eOvp01BgPDzvI
AcxZ4p9AYSFiA6At3XYHcDB0eMvBUmeXfoKqcA7YPLvBMK3b8Df4h2B5JPk+BKmQ
A3hNY8RLYF0XGW9cCsC5IFG9CT7fijKa+Q/cLAcvoceA+P9UMQ0B9a6JryZdWqXg
ooWDNrMYBY0KXEEvdYFfTd8kKbFIuc2KHWMPMGpVWtqZTiirmhSt5LSoi9BRubVy
VcRlXtOmfi+w9iyOI/eirh8qIakXZSSFeTTwZypiumTrk4/D8QNdfZKDG5wkjjnO
U3JBIuTAznp7OFTRJRnpvVNffOKvrpZBPOfzi7rGiDSo7JnWVP4sfRFSKUJW8b8n
g0Q5w2Wk3W67XparJlObnDbENstfHmweWg52ml8iwTUyY3PHr9w/2MAkzTx52MpP
EAfAzTaylBxiibx797luOMvDQtCqp10LGTjS71bo0hScOcqPWyxZCm5KOAFAAf6f
vEMwvkPGUO6IY3ghaEY4KyWapU5n/wtAfDEUgpPsP/NCOc+buwf3W/4pkfLPKgOu
lYIWnZ2Mbk0i997rYdWgjYNfsXFunUjxb3ax1lixZWCILeAMf3gWE0KD4U2aSi6K
845uNxNXkre04aya0XfENNvlaOJmxA4YDYon6Gys+LXhw8RFI2AdhFFlE1+3FnMf
Sjc+dOjURKa27dbm5efPV3aNFbAyZnSQVB3IdIKgxM0TsoGQZU3fsATHkPQPL0xb
2KwRD3S62sO42ezil36W3NPrdL2ea431KYc7d2RzhKc=
`protect END_PROTECTED
