`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4ucZAi5zvT412vnmW1TnJ4v1zWaRatdmXpWSVCWU0hSA3khTCCOiQRCg6UdVcbj
xbAH5q5Bn0nskxQPlgBugayJcQz2ktqZp1lkNF39u7sSpcErjHBrUbeAPQs+mwju
YSecaYDy0fzx6rfucVZiGE15jsQpHR7oBvNFF8C3/YNnLCEiYRRhbqU86rSBVNNz
p6iZvw8Y83T7Jdf8g0etbZ6FL7KBFt7ZnSxPRiIyZcs+G6oQBOP+2tmEcfPgC6+f
ewsw/O2rfeReLwS+/4wzuFWt2OiTrlnMWmag0F2LOwagw70LRDTPCP4BxjWDHKJz
K7HRaexOMsR6j6eaVKSxQHndfPvs1UZcGRKi7BKu5+qdNXHLbulR6hmN5LrtBHGi
Sw9mPTO0KoKIpBASG+3C8jDVQNiYgQ9LUMvfMzceXmH3N83Oi/iHwhHYMpk7Dwk0
B8zw4xa0vfTFQy4cvWTPy/Hv9IWUx2+9wMsbFsddwP6JrEW/QnWUUW3CkFmf0jL8
1ACZK1YpzchCpHl8pzQx4tIsLVHmFPG8uat9nyP4uMliScylOprsfmop7Df7cDlZ
qn32/opDGfdeqhDnhFOUCnnvfKJWROHnMns+LMhOQe2+Vm0KWNkoRgcq7tjETiL0
2PbtkWgZyZDx4+d+ndSmEZufL5inqCemb5uJhS4M6IVSl9H0458RWHSb6oEbYUDv
YrPaZVAJGd0qL5aQ770M9sSs7poB80QzoYTDlkMKe7tvR6HgrNiotxMadI7b4VA6
4ZapZNSC1wZeHlBeP1N8X/csStDv+SuL9sP1D7Srej51/fFxKy7hLEhJPh4xtPl3
89QUmI9wUD8mLow0e2HfIWpbp7jVxH7ocHFpfMIFgDQOzH6MYiJXZuD2hmo4ZpVg
ILnNVSHtabYLLvnTS094MQnSK+x3/WKT80ULNOi/rt/77bkf1XHxQ1u2GQjNnS8x
OHAwChVtSpzHlySHS50F2aEV7GXAsecUWZ0LCMk6Fg0+Ehl9NPU612Flvp1zlcCV
K6RQyQjR3vVry+vYcz/hVAQVg2s9WXjMuKUuHmKXXisBe8VGDKEZIaeJpkGIcgB/
4b282X2ZnddP6cnEeECqlFM1Lk/eIYiim1qHS+buqpwfUbjYwALUufk2qJcvdTj/
PIiBbdDWzhME2JlQBRdcDX26IF2vFm5j7Nsn8D1CzPEb0QctCU+Fa5YOD90lwrgU
e84S9IfICM9bXpv/GqwCnMsoR4xFdO5a7B4l+uqwHpx3liBPCqtJ9hEzqCFadf2q
orjuArYvd1/cntIxQn5guAWkC3Tr8L9wcdWAFq3kAW7Ipe086DKq6AXKxJDSl3R+
VNRSgwPnqwDUqRvKJFQsKVhFvscZ7lquRETG3v8CG1ny/7ptliop2cQDwSUi6tnC
RY9VV1RJoJjKotqU5Su6LXF13DVQXY8YDekzI+vNpXiSou8Cmjh4LM8MaPaxGobN
v7e5jGrIGNTb637cMpFVIWNYUtVmkqEQpJiONpo3T3ZQ+yeApajxOpMQZR5KzK1t
8h3JWBUydi5ZncGJbyRlCRs+Ib9NL04yqzI1INO8jy4=
`protect END_PROTECTED
