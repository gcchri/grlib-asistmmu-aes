`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1McUzAO/lU5pH0i6YNAmp4aJEosesTB008+wTuFfA7ZeQV1PGXEBJ5Rq/0u+/yIh
oTtzW19kmtjKHCHue/BJG1tTOxyYq3CH2V+J5avBCXMPCnaL9TUh1d+qyEgZRrDk
gNz9tjhzGlVW0SM+X6nKUn39ueJuG71U7I2koTVFw2i65ibBTmnVNVuNjsxpz+0j
8fKWhY3sIbBBmNFFo85fruvILWiPL9Dq1dHGTNUySTfJzeI8mBVJZ4aGxLyfzn2e
CvToMwksaXntjBK3oiVIKaz9suNGSuuz+2MpbWzsdBg=
`protect END_PROTECTED
