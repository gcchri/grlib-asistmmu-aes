`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M2rM+B5tG++1nI0XnJyGO+H7J/CGbO+8V0bx6pGTDXTk+P04EHigsTLhgjWzz5pV
WMoAbrdq/9WmamCsLZ6dHYPXUBWJvQBf4WcB6TfWINNYswRLbmL4yF3PafUqW107
cwmioR0tUIqLBri7lXyriC6LrjWIr3MDPQpBXTCoAfke2M4Uj+a1kStn8nUoTdQw
zBe07kLnDzdcg185BHy6ovCB9Fj/hsSJ4XmQ0rZM/ndkjb+0teqtW/vcApgZwPYE
XLp+9+pAkAErbM8BLRTkrrgSx1bUGPGPbiQ0MsfEhpSsnYybDvmPTCili61dHEHQ
CGFj+CCHAdDGHVwFu1FNRERxhyGbRQpG2xOoIVxaShV3GiS5TfkMpUkCs6uRuhRL
IhWY98ANI8GL2VCcmStWusaxWYhqypM9HAfJUy4YTqgM8dIXPbzhuNj0Sk5FNuO+
EPCswfLWuRWxijHTh5tloMkOeqfIJLYlKSvvdJjIf/8SxvwWlIEERrsFMeIKP76a
eR4KsUd7RHYQv2dYkn457EvTXnXdbzepRfdg7v1wZjK4CfZ9S6U0K4kvt/mYUwQv
CLXThQR3gJyQkNp0Rf0GzrCA1XEv9DQjeFkaRAagvOPbeu3S3ZCgORTmHS6xpnXD
1ZmK/pmRCquiyHM3JnETuYtAAy5tOXvgD3U+s2swzWgypxX2MP4Mw8fwmVD/Y1PX
7eQ1p8M71n0XEXwkfvABta9Sff9YeXF2JbD4Y/CK7ZSTFBMb9uGBeU5V0CqLfUvO
`protect END_PROTECTED
