`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NdKn0N4vuIlj724O1zB6WS0u/ZNbsTGYDUkeOPc494b2rgHTejSfuhVU7jXaVDjs
r4d7Rsu+tJjlildrwyUK3TM37rQ1LChGtm4OAL8pgFn5xjHpkxS0iqLN460sxfvS
4RTU3oIoCXIKky94XeytOweGwW9F6hYUtYl+wqa05TzUcTzHD/2CA6hJde/A8uUY
LKX3ykuBZmxxVoDCN9Is5oqyM1ki7Ytqeg8LBVF3y9jNoh2oBnk19OYNMB+oimmL
91mWcZKXm1H75329oMobaeqOqYN99ulFxIzCzmZmVeg=
`protect END_PROTECTED
