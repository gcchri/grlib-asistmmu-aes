`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
riHnmYmW7VJd25SIBLzC8VsvsYJKMWjQq5oQnpOP4nGDLzzk6sGxAqfYY7XY5mGC
P6raMi5zsZ8n8WEsG3yB9uJBnkUiKKTbK5etgBL1AY2wU6KhqBh6+zsY+XEBkRMv
g82kZeta1k912velANrbmXaTADLTcJ9TeIAs5TPfgAjTPEajXLHtNt1OXEBEqJd1
bYSL/BuE9StwE+JrWS8ltzeErvzZ1uM3UlAOFnpjz8rBMEzbB4FuywiOKHZ9N/MN
qzKvZQCjocuv0t10heSuXEWbfoh6mShlRn7qlzV9XH1OxYiCMQZDJPiJ4QCgUNZo
KLClZRT8G1pPAQNEEKpQ5tFhvUwsY2flNoH4ZeDREDXUbWWzUtcp0j91RC4d4RlX
qeW+r/eAlS5pytjV6gYaHQYwGX5CkWJHRVH69eQeNDyj21FTwK6zpnGOGyBYKzwR
s5qaRQD/0o2u9qGttc5sIo375FLfsdV0NAQKK7xZgrE=
`protect END_PROTECTED
