`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsUaB+eWvENsSYnRDrucqjkrFx3szCNuw8bxrm6LF8SLGTmYSqhKbSx/mCOpaK8o
pxDqFExrSwzh+09CxM6BXi8FO8mSzT2xrULhoaR/A/kAA8YKHbWkTVd0ABTD8l1I
LOH2z55MXKje6WcsLqDIK7A6m/xpVEG1rjZgun5ZQ2W6zv5GzNfu7U1YjU23tkBJ
b+6a87s/hsKQ/uCfx2RrPIu3GmbYzghuWnfZY1tl4SiFRJj4qAmhL93mOC0zqlO8
1g8ap2TL+yL8IVCRCxK800Yn2BhzqpRlPmNJ2scraY/3b9wuo26cdJ9wP/S12tyb
KVZIBWID3ThTEKt5yzG0L4d9BwtCO2SLnFfkcytgPfuiYljNNPIwH1ybonqJfIoQ
C2eNXfmG5rV9DPatr2xQAgIRPtBd5NlC1Oz7N1Z4s+L3Kh6z73UaVT77ftWt1ABi
cTyOs3EBZiWWFIkVmdOPDX3yQhYy0TR6ZGF0OZowJcU8wFlvdXMCuzCk4vziWqM+
2oFjbBJMaSs7i83OG1qmMPssjjGit4XRBgBFAzjhazcWDQ2SRqCyj+5vmGrj2KoI
+WmKiqltiGwkCKOmBxmIcbBKMITFc3oS/6219fFTVSUCj2tSy3no9oTgeVIABuOK
p+hFnELaZ/rFeoz/hzKyJl7SJAz5NzIJHRNpJigvsmELE9L2ve59DPfc9trfjUOj
+5xOmajt3C/DHGRKt3VnsSACU6dwOvqHnX2SmEDJIKnMSTeibPLIQsy6+syaFR3D
n7rIGtIH74i/MHPtPOWaY+KCh3dIIH/7PCXWmYd6tDJmGRdO5yjUXakNkB2BguE/
vO6F6t24/RpWQaFoClFO4OMo8bnlH2BREs1fon3iMyW35CNooTgpAlgWE9ffatwn
4RMWRD2SwXUg/eBeVmTIrszlEabVsp7ZbQhCxzxtkxJk0oDtSUTzhkCoAqyRsgTr
UiKog8SBZqD1lQ+BxE/kOcbNC7n4xyGjTJggrs3ExFaDgYHElc4zfNzGUMeMKG0z
zxZFuSOyOO+vP28mnPp4ud7bprkOaLoahgXgLGBC3cKO1S+kKTTsRUUDuQE7Ewr1
fLqlXC99ipPJ3Q7Jsd8RZ21riprbI7O+XRY3Y//FH4Bp1ZNawCrs0vlVNmcXrwPw
++qjADIXezQ2uydicLjWkqMSWRMerCPvtgMHuFJUmQasRoa3/HH7vC0Gz+RQrH7u
ke3uHBqt7OAS3yalWj5fF04edXW6fC3mwVNo28u1E8FE33b65V4MgOyo8yI4y6OE
DlTdLokSwZV1c0eXG0J6RQyfkHNtAu8EAEAom1uWWmVDPShZ4kubGeik3zrAItSv
uzOxTIVsTofTOji/agdsrXYYd4DP40kblkNJUpAa7mRAgPaashiL4n3ximLNuKBf
oaQDbPuiVs+Yh8msX6BPA9BR8CKJ3KELBwV8vG6T9upp8RzuAuYZKfaFduXWhWh9
+/rG5hbjkQcXT8E2qFU1IWsInyZVHcr52aggLn1TT6Nv6aVAlv1JCUm9FegEFO4p
8CoSKMPu4Z8A0TkXOo1X6/9cpheTtc7f0FHvrigCmon2icUCxRjUwRRFO0cBhY+1
fitosaVsr7OZoSh+IvDOciD26R9OXS7o3NIYssdGTPp4HxWBn91YyBnn5MtbNjJ+
JSgAqi1p2vs6cRsTIjIZHrXU4p9B14M6uaYD/UxW/bL/nsW74nQ2M+5jbzrqfXFe
rFJ+Vsjd3jLR96SErW9ENd+v/pXBm0WwyIqtJsMxiz5h3qOpP2ZYIp4QIa7JLMWC
KyYJaNRYpEEL3yiRapeurCNPFuTrW7jAgjciJ7iqQBAO8zU5gLOptji/n3hlN9AK
4zbwT+RRGz7hVlXk+5qn52Tq+Lf82qiob8tokMMqdv5erYRewh0WvbBLSj8nfqiT
cvXYYBRKWhTMSzEn2eAI3/Gcm8oITV88Cgdn5acmVwmzkO006w6ULOYBkgd+cjjw
E5yLHT4VLasH5zldtsTp2VAmnk0PboN3WNDd2pKFo6i2AzuLP7IYYbLmKtPph4s5
c2nJmrHH3f5wV+zBk98AyC8BjWYrZyWr7+Ze67OAMeSzYV4OWi6fDTUGpOq6rNgL
s0xC5wM5dlqzEF6AjU9+CSFs6DosH6kxL9Z6g0BVN5Xf+uO2J0fZcZzSmDiGkSdS
12KgKGBB8AKcaOuQ0Jb64VCM/0mor3PJorH8wiFr6iOrqpwaulpdKPncVEI5c3x7
JI/ZWmJgHyqgc6YfCB/IV8Hh4Bs21xDAq0FwuLcLAdCJbKQ5hOgVa//t/2E0z++u
`protect END_PROTECTED
