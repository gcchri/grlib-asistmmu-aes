`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBzDvG+to5ZIrA97CPRhO18mNMdViG2I4qh8kKyts9MlDbTs9XcjeJ3DFImKzYh0
DaUc3GiLQEgczFGVWy6W6ITDQMzgWjHqLxAHOBIele0imVcZYIw1VfJrJyA+80Zj
2mrqOhPUa1QPyfVNc5MuxhS/fUFbShejSsuYtcubUVNZlr2kHzEp85FtojLyMi8H
WOEXRYyklOQUopDiL5XZDPqCr3PR918c8+3bGCBeHHbKAs5X7RaKFjMElnihMddb
fjgmBd/NMmb8VW+XY61F4fbn5gnGgRl1TmWLPZJIA1O3cvpMa9M2gj9MNsgnI+9V
JdqEZlLVJKbnFx7fpoXMXVnLNPT1XTd1hi9aNvBQf0BAUst4TpmMnyV3tQHFw00e
FRezbH9P0TYjX0T8XfU8Ra6LrdcvMyUShLEuSRn/MqEuV3uN+s5WRpXSbfG8/vhQ
WBJR2zgEzTW3naA4gc+qCvkChVnhp3H2HhlLHr1ArtiUvl6bv9G9ukd0qedAR5sR
6AYjtoiaAolJwYHVdiAsOC37xbouLx9M4Iifv5Cm7pHsBfwJAvW/OmCGkYyz/ejx
SgfyQTW72XGxiSXNln6loVi+0fy33YDWeHZ6htKxShWo6htgPXAGtdtMhyWjNSlS
sh366hhxa7c/97X3IIOuSpWhMZ4YoYGfjaQXlw6izLv2FOBQzOQPOodR3wsQGXRD
vc5o8MA46DyEzg/I2wvXzJo/7Bn0rrf3i1MDeYQL5xHx2eXL8c50AjidBWP5IMcp
fgRO6ILkvCf0x7wsTU2OuB3FMqOXzYntepmCaaoLvf01y6xUm6UiGzvHYcbITBnE
`protect END_PROTECTED
