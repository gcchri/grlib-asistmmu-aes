`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
47egHMTjlEwdm6/iEJc3PKrGyf3a+942kuMx+zQ7ktS6ak1HKS0O31A4YThGI0XS
EOWnkQ7jDmSCcUNsUDwtboCrLT7e3fVwOaPXYJtgNyCfLSgLi5OaOFn/onFDjq/u
5EOl5AqFvOF8pIib0JyGm4lnV9Xv0qmYMuELBptjvK5XmrSkjXU1u9RBainN6Hgu
8rCNdV+2X7cPmaDeFKUZ3oLr1l2lGNOtItzMwN9xEUVLZ9Y5jANqDJ0V9iHGzLeE
cInKnVJ4MeD3uMQIP157QELjPWTgRNMgT6pRQtCbYRWEUWJkeozE7fVNoNmZ27/f
jsTphxt8nJoP9Z+om/JIfGxTiJ0hsVmf5Ti9+dQqsrDJ9WulFzaYU4HebIuK50TD
1fh+9CKEir5scnvfiUGUCX0aEvRLCAn1SASpxqOb9nolD9Vc7q3wiinbi+8FJqFx
wq7sWZTjx7yc6OtH6Arx6eGW72Urc1IuMjSwCRbSQq89KuuP3MCEjzpOplLbfUr7
`protect END_PROTECTED
