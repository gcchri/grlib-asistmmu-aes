`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlLui1k+2YG2+KjY/+4QCmgWiSdfzhJKYN6I1HLqZU1BIyBE1qzRn15ISz5OJeng
yp6WXxukOeVzMYIn4VGoq8DrxDg0TP7q5gJsgbzm3YxnzND/X67t79h/dDLykutS
XuLpIIpvPz9fdU+ciB8NT9hWA1Q+vSQ2NXZyVUDrp9ZafzIdTncUhi2f7U6VgqxX
41iXIeE25Q7RnspdLfjsKPy6r6dBAsaAbFOkfq+RUkJp+wRa+/jigM6asqOaVoro
q2aG66TSZ4N5+/BQSRUixVtdIl5gAHUK70xBCQvh01hquY+Yxsu5x2kyRP47ErcE
i+B7qE8NyYN0fCHWsGRfw9EcrqdXcFX5BvpFSkBmoSYUjvHzxeYx1RaXWsZc5cNX
AGJPMourvG6P2L1C6hTVUQDG6YymEzT2WSWWwLZ51AhCpev2KpCRp8C92NkRzbA0
fX7RXLmVuA+KEgD4tiyqJGca+F4G/iDvVombQZl9B6V6SD59qWBVIla/BVc9vU4e
7/BhpkAPYa4t2nhwWDasOwyJU+BQiYBKhfeTA9dWthwgHpa/Dy+ZeO21MKWU93d/
VjBnmXeKx9CNkKaVEDp9uXG7kSd6MvdoK/VyNyCO+Jq7EoisgMEewkkyf4sfcw9N
JI8fNrQzEzxTeu+VOtUezwwj5mJRJIC0bVJj9NnEbBaqmL1I2uOTV+Y/I67xv1gw
hgra/tX7y2HgVPwdoL8MU7pD8yZmeG/IuiLgHA+xv+vPgt12PnkJ4VIui477IW8n
Qpkv/r3eZneOhksJLN9hvJRnAlKmVlttvTKH5qrn3qvBcbEUzaRP9Nsoh8H7a3Aa
VHor5tlBtvBeF1y3mzSFdZmXYFXdBaxcO1atyz/UQOOt7yBKqa4A8B5o3SyQZsx6
zoQ1iK4eHwz1KqHGvGD2Ldsk26x4+hmYAZyr/Z+0KvGOdbypXKajjVvwftoZ1Eny
Lpyg46wFSLZxOFH+EJi3OdDOxYXFeu5fJt5hIUzpzJCdHUumG7Ohl0fEqq2Eg06c
5gF7pffz/h+J//JfwDq1Gg0uURGvWhvUCIrBWpYy/jYMvga4ILwxPWT3Xa9h6Qkz
0VDOJ2a9MhXO9UC78nw/JbpaRpN4Ts8r9ZtDMyOWeoQmH2p/jMpPJaJHens1DjW0
/BX+R05cuqtsK4bNT5tALkjQd+MbQZAT2XxRhcWHHnO/zpcY2fhCDcwzYbBPU3NU
VPopk6IPbDcLTz42qZp7CiSkyg3VwVUTQBjVB8yL4OD3QU9+4yY3/NlFsgm89I7o
2VJDqfgb04d8vEfcR8E6hvHlvx4A7ZYX9KLxukU0bJBkpOzazUcZpxANTVlvfrVL
Fltb2KYnejQCBG3FezAXZGt0fk4rg6ZsoIWEoIiD64PgkeLgfaJbSMYL1pRDiu2P
69pyYbW3OuN45XPJO+SaSFBg0Au5qEPQEO4vh+NrFZK1nHC9w2y7DwqaL7WbYi3R
br6RQf/gxblw+pQHIAEh0yjB8H11T6Cnd+fsXhthAoFEsM/FKSo1YKw569UWIZ3n
+FBIJCl0xFz35D3Qt5wWvLnkHrvG2B2i+U9mc7aIhUXmhZarWvxjHLabRWTP3IES
HNf/hAeH1HNRGlc+4wItqQi3FEhLQDedHWJzKvSPY69EOe4cHa6mdKixU7racmaT
bTXhFwqSOcn2RsxuMbN/hxmaA8zTLbgDOc3u41UPhMcqLqT0v31OxZaV50mPcTTX
zGVRhHuayklIR9ICMt+/GYdIlUWErx7AdmFbGzpCzmNFuFWxvWqmGn8b6hmJE4IX
13oF9f/i0y8NT1SaDiDtm8aFtvcLobABOGfs5D1n35qLuZ6PuGeLDdg3EjqhDPXE
PW4SYlNzygFfrK259DRZp8A18HX9H2ZW7aWmeRcv+JJQANeQ3oPv7BYZBt2CH6qk
OaRAdPwelQl71xtxIHHLFTwQJynESPgTNntrssxiuoX22vdPGbUo5bpEa8Xzlfi8
U7PtThSz3LWgiGnh7xIGhrjJ6ConxrkU51DV9Pi3KW9FXtqfbhnd0LXhqj8CTn4l
rbmDXD0HnKMjdamgJxymsWdctINmaFnX1lU0Xz0VS21CdQ8Ou25mTpqJlGHCPZCm
DtmRmPtQ+PBPSUMHpxNLxEINgzyqoKXrfrucG0WAOYqOCNqAPGLcoFY66FE8+4bN
2zSiYcZDvAEHbFqhPrYDR1WwwUkeWeYoRrFU61Q2L9OGZQDOmcgA24DahPDBXaTF
rWgJB/lhr5i2xAUDS9WX7f4nMYtVFhQv03V+fYz7p99T3wTQD4V8fdbUbDxnzz9x
G1S51S2g/yj3CRflC1hupUvfZBlhQCEM7KP7HVXJ8ovhc7zecz0C1oTWyDYjx45I
`protect END_PROTECTED
