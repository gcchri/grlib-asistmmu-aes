`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgxNlG7NogHYlryYihQXpzvzZ2q/CvCQRec0t9vCZok2oRK33EDupxrakmstct80
UYRjnmvC1Hslh5Mo4s0o7jyTKvD45oVvcnSaXJDCkCxZRG0TS0cuwIn4X/Mh9ae8
TcG5SMgd6Eyp1Uermzo8XpJciLnugg/h5llqg/R6uJnktMCMY/4S//wSPyuTIo3A
Nq7HiTUZHbnkpjCnglNIutzgT0p9LKyTqp6orVaGJuWqNvugJ/dfCRxze2fLJHBz
y6tUIz9BPi07Du7maHZtanYwvUdCvZHA4kGqJRwjaxzJQAGccPosWqFkV8pUdYxn
PIsiIyG8kFyshNMGGLHkT23m7pI2Z/BAzaD4Vecx2eah/Tuh8Q7xmBnRAs4PFkcX
I1Ri0L6J8c5zFRx26PGApM16FCjSIqXpMXnyyK/iUic1tRxl48cinbbHMuHMGUXn
UaiiC7PbFLaR9Smzs1lFfCVW3naoTF0M7dFMSyvBx7NTXDAJ5+vny32weE1tlGd6
e3jMaIFRCSXEjIvytsETxC2kN283LWRmk3Q8VlceU0PDL5M9jh7Js8ebsfGOhTEQ
bHmUJQEa901vwhEofilF5Simu28kCAtpIEuRoNg2eczBOwMgVWmOjOqvfT728fag
NeUiPgImzX/IrAabpmH0/o055hfZrd8d4/+AQ2c4ppJV9RY5mpf/ZW+IT5prUHLa
`protect END_PROTECTED
