`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xGEN+bSt38J0stwK4h0j67pTka7YnQmPQwyeJ5ekSx1S51cKuVNIq/YYNxoZDj9D
ajstH+tVAeW9+Fgk88gxb+KUt84B4iR7MKZjKS12pIWYqI/UHlaejjk0HN5dgudj
OOA62B1qgsgmDxyC2RGFgITNmRGrl3vwBZaRldXRBmYVGYVrq2hO6wREu5lrmTu+
fmUXc0Siqtjg4AsE4t+XyxRFxTNVsiOcryBk3KE3IWcMDZbXuUCQEPVNkPFF7m3S
NYdusy6L6QE950xbY5nvZwawD1nG182VUbYcTmqYeTJKUioSeqHDSUpJvPzG79Gv
3FfZbJohDjCIyPPwru4NvpRLpXgrFYR5euBqalTZPzHNfxOc/HIw2M4fcqVjEcAx
FFEFX3zH1no83hmLHhSjcLtriGHR+B2m6t/IGEhpuJNKjANkRTV0CPKPfEYGIIAA
1a3z/axFmaBOJcDX1GakxduZeEba3sQP0tYPGS5WMs2gtAVMcpTsefUJhpbqqBjm
`protect END_PROTECTED
