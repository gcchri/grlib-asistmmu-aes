`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INhWsa1f5TvCYFJdt2EvsCj2U+P7xQ52QWaaJ5D8/D2jhVNHCwkFrusk5u3tmoaZ
Ebg/drZWosXTRpp7crnFYVAJdmQStXydOCdjaPJjs2oiV+24RTgG/R2qCWnacB4j
leyuwlM7xJZooG6BV0ZR0jmi44NUrl4wyTGm0Gw3uc+YQm4pXplSnjPN7WlcU8Ri
Jq/kw7DTKZIc5M8nKmEYwVuiGFilD1HkeWZa42MEJG91ik/xyxgn7BQy7LvHULI5
V8AlZD0C4GcsTUkyTVJwkEgM8vRvrn9NNxc9RcNL1Ybv/XKIGJxG2s51vVxaI65b
bv+lcx/OAYUnLDS0NrQ6ibx80LufEZulxEwBNs080kEOzNid/iB56gD2zY3hFCX2
2xxo/dMlXbEGV74k3j9vktPNuT/5bZqlyLy8we4YGBrF1LID/CSPZ3EEYS576AJg
CSv4uV39UK1S2QG4pKJjTdxClVXjDpieCWLgHZ/mFR7UB0ODEB7HGCYThqJr18qH
`protect END_PROTECTED
