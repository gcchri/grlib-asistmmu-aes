`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RTvlsFzKYUjTWjMXY97dP4Fl3isC/+SAaMoz75BI51Kd0yh8x6ayvOYgTHmKpaVc
jnJ7Nll5w0icQdQeyvpUDP5b0/ofSlQVqK7Zinjn9E1p2oGSMQ+F3xhwBHmwRwzW
LVTK/qxNehc4B4dVa1lkiiUDpZFm0EP/fpKPywz+hgR9N7w8GVlHBTUl92ToeEl1
OOAihq6H1X2G9LeFWuVceg+FadeS9oGAgdKSPrTIQYghohNevnF0skYAEX6LOuMY
mDaurz+LxVx9McdaF4E9+XFVY3hIk/rlNALtX5KYaS/rQepabIPYeaLRfgFlsO5b
3HFDvGE6P9NFSJimfVNJDw==
`protect END_PROTECTED
