`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzfgLYgOzRaPsjyVYavymVk+Y5yxU+JjdfeIDnCVwECHU1jjkCJDnNENiXZHbcJw
qsgWMvJAvMSrycZYxpLRx1tl6y+PiW6Ijh/6FdksJQxtWW9WLQUhnTcUFotisrpT
NJGkSnzuGTRk0T2+Zqm3cLEoaYQovNP2z/PmBjyxCxjCwip+GY68PsLOxluFxhcL
mepkfk0FKxSQT/QvisdQyt6/1RMZWEAoSjYyJ5u+m0xzyCYOGGwijQatGDJOp3rE
VuNpHhccvRSsc9poqltUBPJtYTh4G1Au/k7jrgVMkbTd38Lvl0vnJu8B9gkjo87U
hLjE/tA7kU8Q25wO4uDJ1KrCHqmFO79Y7MGMUDoBYrkEk3eJ2inEJek4hUDZxZgq
dxg83htnj4Y3dUTW2N2D8Yv1QwiuKAzPnUQOabUfy8H7muLAl8rNAzuoQnHb37FG
abcDpeCwF59TwQ1i32MW7Hn6jMuZiXdegpqJFpaaCRaghwixtuDNiWski5L3fRCb
ER0th2cjH8m1GhfYc+WPqKmfCLwhLhbUkI/365YfFdr2A7F2SpnIJhK7oWd2rheu
iBdawyz1QkxtxeSUGl+5/Z4yJdF/Jd+QC4nea/RmLCHny0g0O11WE3OGU2bhUw06
b73dHaKpJDR01UwV0TQfzKuXsw4I5SNwWG3M5xUEEZjUpjrG+jZo+A7isIHM/WUB
hL/ib8tF1dAtZrQ07YU4YR+MhYzhOz1rjmn4lKejwGTZ8HQUBrorDLlu/cVEQwZd
Jl6wlLI20uYPikqjpeJY8HLU06N+KgOGFYdoO3KhxWld7JwevXHucINQSeW+Q7uz
qUiOWo5QNA7pu2CZ3wVG3THWxLgOUWwKxqdJGVp0+x+NTUjgdsIUbKNZtSLO41/h
nkOdAxYqOGDUupmbOPPo/9InMl1cBTHf+eFhSv2IYm6NT87eQDya7vCSXfrZ5uF4
M/BLnikzhh9+b17OUQ0XbMglbksRAcNXoXYFsMD/rTxBFICoOi7mBU4fhTHXXvfY
/r3N/NLULkSIO8mkxHqCNCudhTqSVQRe+VwgBef3TCVX3n/B5mR69aUtaKAurrtD
t71V67ZByoslSgNa4gSg9fVeeS5oJNflnJldOF4Y2hOIHvd6k19HG7VmzHdk/mP7
c1iaHXvo1akA2rPR+M4YoT4iZAPpXW/yPACIJcT0R81zq9CwrCnrS35gDbmLPBC1
ZMGWojjkvtMyrrhYAVWYlmnCr2985maAVMFIDb9Lqkn7hrS6a4FWlH0Jr7fkUhrX
e53JkBXi+50Y+dZq0p5qUoKWFoSkEu/9uUJOys7bS54jAW4YBpmSbcEsDm0+jNL7
Gi2eB55LmQnGjNrHilmZKJgkIAE833vDpTAqKYT27dB1rXCpJdhEXeEvWJk3MgTE
oVeHKs6gubwk3Wjsc8G1YUHihvK4TcL2Wr2HDnRjB0JkncQuwg7TZmKpfpQVNL5P
lOt1HSsNOzsl9dq1i6MxgvVHgdbEDDZAdfYoHSEAt7SxO9Ion/TrpS0Yd4m0I4Hp
ld3J7rTMIZqZSscjF0c5Roswz5ZMiFpIQfcYOybAXa1Vp8kABQlIi5JLwnwQT4S3
ThVrrG5X3UuAqDfjc5bNU9zlOYL3WR9aifh7T48IMifiBAopftqvk036GRa7tZpZ
VMQcNV0fvdt15/lvvJX/BK/wDTTJwLKX/Bh17LRAohnTpjp6qAdeTiICZN+ycSAa
`protect END_PROTECTED
