`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r0KXwuoMY9ajJwbO0R+LU/ODOMIKa0EJYHHW+iCj7KeVGjJklQTKMlznU+Y7FsV2
t1J8MvmniocPcnuguwFUdQEych9YVSdYEAizL36JqS21pQA50IH1gQOT90eZd7kg
ST9EqDiw8hRNtzoeoKeyyAKmCVnUA9UEQFjjveEnczRt2wPFv36HZjJWRo/DH6VG
VkQELL0ETITM9S/cYvPin+qfdAYUCdYPMp7XiWSf1CKbINnyPaAU6+t3mExgzRCd
LWG6ECdYVOjUSp+ezx0LWEjkpsXQM86GhLw1lBuE8Tb2jMF+m1fQrwVnsvtLRUx5
zcUbzDpVRgdHRa/q4rL9zUzE6BoLxozFvsEfgck79JpmlMnqHSA7O5gpN3nRJMrG
7obHuJa6MP19471PW217qZe2aWBwOdY6HRPWdScHDEhAQ4KOyD4oV2iLfgDyc9QX
`protect END_PROTECTED
