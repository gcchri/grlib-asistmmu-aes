`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wWfXFJtNXLvclpOcdHIUu7BtS4JYGK9LPwLi5RpmQdrHT2xZH5CECyhamuCrInh
rgPd6uQBUD+9ckiU1bEhMCiqqstJ6v6TIPuNfH3OojjBsLwbDb2yh9rXgFbY06HC
t1+hPS3pwljR6/AklW7PVxRqE4Y3cnuvwpmJbQRZnk+nGXWswx/e9pn/d2030J/C
vrIn4rr2cHDdfAiBQlk0vSW/e8aIjs+KsydgrxQqDSFRG8oGC6W7kSYoQ+J4ESYo
FxR7+yYzwUlmqF0zEGa6/TK0eg9s5zgG8nRJNIwOqpKQ9mYzpv3QIO4vdtKlfJ5A
woP/HCUjGhM7+Hsrd0Va28dysgyinMfsAC+9Sb2n1dqE/68b5WJ8mNxUNedg80UM
FVSPro5h6CAYDrjM7z7GTq2vIw+JHog1ymE1wLG4WEnfLXHu/Mi8AQ3QPKJGX74v
+ngCgj3gSX38p19XQgAbDRU2Ke4a6bGVvftal4ZT8jKjXQND1b2nqVAUXiu0EEfy
3ybMi6jGPxCVRA7bP+SEoJMheEQO0B/JIVRRr/ATel3BzPRFqkU0jVly7lAxoD00
`protect END_PROTECTED
