`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gBvJ+8Tzwpfbdq03FPiRu3RFok8U7zAj/EkLy6FGQJwXOKaCzA5ltE9ONdaJr+Ay
lZ25uT1ofN0KECjNOJd6KHQvwh2npQFubh1V4dQJIvqbI1CMtc6AEYfybR8z6htB
xIeDsIylcM9vMEkYYXSSX6HclCHFE5OD9P8QXVt9MF5ztaLRzGStOEGarqSHksSz
X3GHnCPjjNCnE0GRVZ0BZlYnu6LZqsAj7W6i6yMYTHN9di+DppYQx3LGAVR9O20k
gCd5xsuuWy0JkwBZjm3v9ANqMxt4OVPquoqaGFpwNTslYuaES89jJuXC8BZFZokw
xQ211wB8ugvtW8xknkHM4/U7SocyD0iDIcBny5KtYXLoHSPB1Oa7aZl+9hJ+wXXx
lDuSAGBbrXkW112ex8AEaNA4l0j2Q7TDNYfNKvHI6SGqsd0gA3z0+qnlCvHYK36/
xNLPEhjInVPJVYPFEwAs6GMzbh3Ymhem1aS94r4b7Qh8y58uFbmkAm3lldLqVTK5
A5waimuH+ADfcp6P+Mlnk5Hiccayuxb3uNXDzXsvZ/K2ZUjyBMyhKNbKTV1w+a5R
v+URl6NHUSVDoIS9+xg84ZeDAm3XrJNeNLwAg0zbdUPkiRYXef676Cj4J4lwRrui
Bf9CA9NBFJJ1zY4vHWA4GoyvDlx/Hp3W8E/1ujHq/ReZZ119/aKz43gxMPYL5hC7
afSXGkfSoAN+4aDvLQfrDBEBS0+zPLJTPjEOw2tFRNv6yVac0z0FOYrqHq6gpc3s
+cWA6Hdp2gf/llX5FbJDxt8q0XQClzn0AFX7qA3LSdu92Ubfa+Ywc7EjuNQm0UUg
MEQDoQPe0/laguN+87OIByrs6MU09xu6+tltetdq86ZaiJQL6lOzYUJmFlcI4eEO
YWRQKakV7bxpUPBSEVqX2jpK/kjnvBQrLeBQN0pdyDOv6MnwrZBToQE+xakDyAzJ
jyd57CE4nIsverHSwRjwYuoGIDmWNlqdbggee3FBdVJ8VwpAi5GrpLiSLPHBTLTN
l9qhCee77TzfNrAJaxeO0IXJQKBB1Tww8uBcLmopXECOWqM4RzIbyHKubyDDMQbV
DvtbVUXsk2LRhsQB9OUffSsD3hsF40Sp1m5gPJf2/nmOSQYus/jxtQAWG7q0mfYA
w1qZbbLSqocMeo+iiGs8tLlKPyPZi/K7EMfarw9LNFnKY1AVvFbIY+T/9ZZHPJuz
kKBCDmdsrv25eEC4OEhzoxqktiVgFG3bS3aoUUrAuJWbBUig+VTNP+P3Df57YDEe
nXAl2H5c/t5KgMXkgvQNgesPOZ9NJKBLHLmzVEnlJ+7dYWiA8lR8VoyzPA7UJJ04
TfI2Rm+cFbCWeMOXwlUUmos8x3ioSRfIgWSweiaFCN10jGA1XmKaE1ZT3BJj/mnS
IcPeabYeWedxBaOI0Z5v+14A829bae3oAzD4ejbp2DWARGgd/JZWkbR4ri1EF/ni
kRv9Z8RiaEEWMKz8TJhrkbZZDPW4euywqVuQ8u4DgNsq6yZjhZQ4O4gtHBNvyaqO
47Vo3Dg3weK8vhU47qQu4Af2fcBTCf5YpTJcujOWUmDIxq1pne6CvXW9Or3jWfTc
jl3J8ZtZyc6PuAGE2MNJE6vqcs9QIcB1FnMdpS2Q11QpuERUItiXDwuRL79iURhh
ocMCmX/O11W7tuK36ogEd4zA4Jzww96t5Onx+fzHsaKHYCDV5KFhjlifB4sOK1Mb
Jm1txBfgCLBAMGa+WORr+QS8Buc1MJsKVWLOl5dVsrJfhCnzICYkM99Yw+cj3Fu9
LI0VsW1PR+ijyYpDf9VuEFqWA+4gR3nHrIGz+9sicbeVj9/n42BDbQcT6eV6yLCP
CyhzRzfzppeq0Mx6YYdfqDtlQ0jSJ/Lfvn6lawK5mLOmvoWRmeU7D31EeNZVDQWp
OXDp7drypHbDVaVSFUtxkvulmJCSxSGhyVpjIeaM57qJR9sVQ0IKxQVWIjvVwZZh
wOxWJgYCy0hFA7zy6QbxnAw48OKBdGcKLgBilTFzB4cy50NpUwQyp7ajcscCVqBe
0C29tGbHwD6ALNsQmF4lr1XoDgeD+wN+fbREP0jkuE0ktwCxXQYfknNPG1kDIUdR
cXZlL+Je4DnG013ezU5ZoU+jp1Ico7fsVm/2eiRja8Lgu9DjIzbtWmwqqm+jl2QX
1UFVrU8gRyg7QO7Aut7FnlnvWhNZpB7Jtn30GjzNYBQurEdxoPGDrqlsmijdXYiB
D6iqrfg2t9MTsrN1EMBtNGTbR5dVysef5ltARvMatQOLAGy8bmjH5uvEmFdOcpMr
VAWsd/KlAOcr/vmfOQnQTgDdKFIptfHIU2ptMyoFqRASSfF+GE9updGbNjnUphx+
fDRt/rdSyEJpl8d/yK5h2Y6uWbmopB84Pi/g7kyzHKdKGZhksgrqfu2o3+9nM7D3
megTqm4qXTyMYRIi9rCnuwjV8TL/b0ITFa75JDGyNQZA7ncnosGykX8LH19BYKtU
PWoDopaERdqNLMBKZMDf/LED6nqtq7sWUr9JZPi7EdrekS1CShANscVzKN8vH6Zp
IxB/umpimspS1z+FQ+JAMgXRQKAutTLKfNz8BBnlSqZXK2uDCFQF2GBntkk32ast
sT5eE0R1K4HqmbTMvd6V4/XEQXTxGMTs4hj4hb4xlJbZ4iJcJH8xuX4XvZ8sYebE
XN7oMDmy1SoTLqu8TOIKQxJWAfqjWHZhDvVWRE4b8ee123V5cMMM9zH/qnufT/b3
G0e2nvQTSHeCeTBbYyXkGkDpRy4WwqzqNkB6BrhzufEyaWI8pR4FWA0mofaQsFxU
iztL+Qjl3T1v8PqOkCO2F6Z/S0SUjITjg+NEKqTgG//aUNKxKtpJTdbQkeEZ9BtD
usnPP0jZ2cF8YBoA99u+Or0Yo5Jwh2kXkWk6qOk85hjm87yoOpW4JUWTd2FJnCZw
9ZgofodyfEoaXfpIsMXZG7/5/TAjhPVnB9PmdSRbGs23qewGQNXnjSECqDevRwea
jn/Sb6/mG55a3fy9EcZSSKKDCaVXq2KdHNwPzLetiAjxL8cUL6Izzz4uIZiR6gLg
IWJxvHSXnNVdoIc39Y9zjDJpTKwh0d4zFXrbdmsRIkj3G/YOaTJy8MFsxigwI+eV
V5HBRbzYdcs5nJTAQS75/RmF7rXt2nKHCBu/H4s8Y+ef3MQZXpzJ2JzxYkgcIwTq
GmV7A6qMiOfujz9Cy6rA1/vfjupWD1JrZPcVGXIGJHzZvpqdKw9nBRdaC3I2ThCn
7XqRcrHwqmQ9+ziu8ZEgSAlt4G+lZ0nepS/IZY1Txk80wqlBJRaL9uTkplmZExt/
nmaqxcWtKRJaQ13LyA7iTrS/uzNOLHjnquSI3OdoVLAN6HaldHHPClSNVrRN5XfO
5igGyFMjbZ1Ra4ExlLiCIdA0ikI/jdpfaA4/JmTY8x1HRe/H3/cZ6LLa05N9pzaS
KQ3CUsKSmlFFTtlGFSq+dJANr2vYJXGX7QZLBz1YtYMmRiHxr8MhHtYdOvifRZ9J
KZbZIqoLvg1+jIoBunoBm5ltYyKk9feT/OAwzrLuT0T4/RFF38e4UtAdDgk1sz/k
BZIg6dc0w/KNlKN1qvO+1bmHocZEShCPs3XZ0Gsp5noHkcMF3dtSlS1UH5s0mE8n
YgYhr25OGHHbRtUAGr6MfL2jIqMHkYjhm246AGqOEAJotbhrGK4n9hce2ZljSftU
IDjL+rAXVwuUwjfNm7hzOxFWbOrwMkmqGDK3DirnLHfzYPzq0oAz8V0mz//FGyUv
jUeeUNW8z010ptzg0wcpqXqSIxDiSlV770YPjnOL1Gbcr5yqNaoRXIGNCCh2lM0Z
gf/Nl860hDVW1UwrJX/89UpbFx5YTCLoUqfw1xJtIhwaqqOUl67pe8meK9P8AQFm
3q0fozb++vYvl1sBwC2TZyXIgxAVTyE+xKgXtYGlP9MM7u1r0A19tqtHRLZegwSQ
9NEYcje/z+syFNXFoR2B7+Bj70y6Xbq70zcPloOc8t+CDV2Ek1go0FZrEuxKl0YW
hp1jMX7DPp//giTV3pD0L+Yg82AyJbMpu+5EdTKKTYOm6OSaK3zrDNohObjOJzi8
wr6620Fj8tnTvAvUyI9h89SYcAuBgjIoECFVwRBCoFJG0zT6BfR9TDa/FHoZMknZ
MWmxdYE3gNFgRhXOGJBqyibSIbIpqSEZP9xdLqAfdgGzWOHB5Pk6dFTP3TIzAgPU
pnjLMUIZjyMugv2GuB/OSfwJCpNQEX0sAJ7sgu3hoVEagyXemI0q2+CqWkBtSD8R
eLAzu5vlxC5yc9qOntidQbuFk5r6mNlAKGwUOSG55fQ6lL/piMOFe1GN39Rcrv0h
fjQRpe+DiRMzeWrO+VOI3KKbx6PQevyXqyTOP8RL3HVdJC8wSkjzNylIsJOhMbvG
H9YCfQCObWDb6Psjztx49QSzJ9F0/6epesgp80xj8E6EGjn/USBFiO+snhz0pDL8
AYuWOJLATUis3L8dLN9M6TXgRtN/xEPQxEZ28h/eJPEk7ZcEW6un9/+MLBnVoSlJ
BrKs8bS2B/lxGzb4IQdbpQ==
`protect END_PROTECTED
