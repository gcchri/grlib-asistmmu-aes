`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UBm7kmuC1DiLX/49296AlErRco41SNOiL5xi2acsaUWWX1aSsCH2EInqjnaTWZL+
r49T+tvkOqFCao0UgnGgHpuVaWYOrdWE0DI1CaGplLK0JkIsVJ/vxJcshm/FD4FL
+KcBn76u4O2/4FfZkQFvC1JpxGHYUrHBXmUDZmLdQcAAs30I3uWEMY7a6XDFBECT
1kmx/bPbJyOo0DlEUDQhcdSF7k+W9xW2QHNo9gkJj2JCN8JlKJSXPaEcR6SU+BCO
q8wyo6DYYFzFzN8LVqdy4xUf74cHOZN+KAGi8euUHcg6heODiBIse1XnmouhQpsG
qLO7VFSCrk3K0txKoGtWF98LpFMNb4ygW4P1Ehd3C8pYGmTkJIebsZkvOVyu4moS
Bco5XaRw7930A0v8FJNAmgwKorF0Ut3J+Yi6H0tMa8okqBAdpXdQNlbfdomCZIZq
b0goJJ2yVo3LSBhYY98qWP4fZf3wbE5l1kdwQa68LxptXHo5SLVwa+biPnQWAcW9
QTHKt/9HaRQBagr3YpLNjBm8PirD9vKHEBdEN5eiJqIB4he3LeLVBGPcjQqeg2Rq
T7UQCCTQvnny4QoBENbbnaZHfNmKTX2VZvv5CuGdIgfmvwZ7sSsGhm/VQbZ/w8YI
/G2HBnaj1QV9dQnpPMccn/cTPK/LRJOn1QNDXztZPCYMttwNjY83uDsdZgDzQMpk
B1Qy9AgPyraTozZFvooN+8ZNzFXb4DEOMs0Oql79bghCDfNjziok2/zfWv0lJlXV
cjxdmlUbbdrq/OacHcGxbDxUDu6grplNfZroxvzgd3jv1GmLC5C+zqCEoPvRF+Kr
Yjah13pPdGK3UBS6QgRUrls0YGPvGkTMVpr64Nn709Ob3Uqfaenw80b43fofKMJG
K3es85Y6I5ltZyqBJlWndJnEIg8PPeNDrtMDnxI/o+vkO9oiNWLDo6gVcYQ/1iXr
Djh2ZcDD/B7UhzxVt2Mt+R+iYJ8H1+VhoVDTPbAY1s0T1b/GXCl3n/yk7xPHo8+Z
0eq1x1tR69iVHAAlbVbAFqpwwhVPenptVmH9EXnOxCV7wFoWUziXF3mdELx1hYYN
BH1/oqIZ5qaiREAeCkFXrEMZEzEMEOu2vHdfgn9vm4Fox5qZ3WXl9oLDtRS/3KGk
CsHLEfJKC4RJ1rirZeNOL4xynsDeRM/Zl8o1WCBHsNBAt00u3cIj/0Rk8v8iqw4F
DOD+nrI9ma/zMlGwcg6euM7U6ABsFopwOeDLCOKDHNHg2rHlQsALrP4IVVnN54CV
p5O1dsBsSoyrhSu2sB386uIUEdDwDhjUiXcJM9zQuErOBifvNbUfaR3jps3g88FR
ts907idi65UnmdpllCb1hybKYr7wQNtK0ubP/NJzev6aOHqdIXj+muKjcDwmEcmi
ebQTrpwdQoZISsa86LsRlTGzZxj2eaFWnhIYIabtIbDhaFs3yulVV+ME+fud1P1A
pwCr40NUoMFhukdtcX5dSwzjjLNZ7XCiWeTKYrkyrKoOHjWkO2Dme8DG4Q1PCVjq
P1nzIzn4+XBRtOrhASLPrI851/FYwC+qQeregGWmuBhbR7yvU62k+ydooo01zOvn
A3fgABoVUCHfkWqTp5Mi1jeRfndIxz7/LyGULCFR/9vkEPgiFp4mqRwSOsGTxqw+
f4qRW5g3JEQSyWlU3wc8aDTNXEdL78KCu00J9V06ZrHlR0XNssTlZsBAmwfG7Yy0
T5PAYioB3XJZQhWyQZ8ns/ebStKA+taj+9Py3UljyIBkPvhgerTupLq6On7dzC9u
YZsnwR3UMokTamPDWqVK7GJUwU/XBmNp9Xh1v+gdd3RjecRFuxYiszv6GGcFBmav
5AhXZxcA+tpyIvP+SSJNEnIvjCFeHofpYJHNBZ28VnETnemBQ75g+E4uWKtmlTYM
XBBAtbB+1Sy1m6IXdcFJdladLc5oh/xkF1QYkaB0J4wQPepO04/0fAgIBJxD9IRf
YSUSS5sWuYCNyQnWl+bONMDxTtFo9JqipGFb9nLcBNuWzXXdwPrjTjUvSCDUrNwW
idj/qFo6cnujpbE1MlYPOX8J7CnRKxvehZa4eujo/Pwq+byKS29UAOGtayxJ2/9w
YmfCfpreBrbnY0VwoAoOGo/wGrI06q+K0BjwvSf9PGzQd3bHjIC67qbp/+7E0DG6
0KZ6+iNLZjJcBYzrkUZAfT2kPIwQE+Qf9f3SIUTgL4rnx/7P1QS5GEhLhFQ2nrw1
i5h4tL24eQh0UUSmGqScmgXCdeHP80VLtLHii829QHMg4HyQmZybXTRBTOh6DBk6
zKUUUER5NDq+I1dIK6m/BZJ+3VGl9ZRXLoy6ahdpo/JKXQx9JCqKAVdxRKMsW1Ht
rfpPQKZ44acwGAVW/iszB8BVSdLz2piL1XDTc6S04IMB33OZYV8iCDAklDKzMuMR
H5BSCyECe5t+3hkbWL14LYc1TbpM9hZ7J8YdDuu2+Yh2Gd6UnbcAeLIkCwNOx3/G
IzkJp8mb42T0ZwcMKflkfj79fCIIbH1QsZhbdcA1YXNjqhhXquefR4QS3X/tcovd
Xg6wRYbPZva8iBWomZiQpvGcILebPM/Ffediv42D3iG4EnNdIFMl1ZiLtstCGQhw
P5euLiFkk5nfC9zvq/oStF+d1jNpEcCpOGDmdjI/+AFd4XdQjegStI4L2bFD1sfm
im4qu7Ec90Lj0nGAm455HLnrMeiEcYEP9skQ+GwzoS2NWmZ1A3GowJ23I+A12aA6
e8MdNqmwrCxwz9voAW8vkcjwufuip//l9na1vttYwCRt2wR+dUbgNqJYagpvoZ7q
XZZQxdcQCW876I2uCZGP5BIVIIapxiWbr0bYuE6sSVkU1rkGrMGHqIar7LgEF5Ct
9jPlFu3dFQ/Zn3bOrrtc4MxkSZsB+f19Wv1P4Bq3g+iPuDUHyhwzRdErSMMas3CE
mby2+tD7L/hb5JeAHsc/qEqsBQWyLf0NWvUjGYM6RuKzmmjGI9VVF/tTq9Ql3cP5
tKlQMZRrZHZ+Jq2yPQ1diVmDe7ItDx3j/R4dUoq8G2eyx3z58knhjQMOpRpXeB3r
ynoO5d2DwynW360DdsADcVPNdkslJpiwDpkwVJqK1n4KjuycXBuzvo2KnPy9mPut
fa6aTRiG/Pvl8lOWpclSU1wEZMEnMYCza6xbKgdMdr4bl1LtY9GuGJ9lntpdCwwn
PctUxIc/pE1qTUCMsu/Q7PD/pgUPnS6TkkB0ZDerLTWsaiJGPHot/RHWXas3rVau
Y8lQlkgd7nVPoQowamEasH6enmrFV9Cg7/JFfrsFO+LQRtC2F6g9MA+can5jQQ9F
EZKqeJCJs1QgWvHS7whdQjQa1FizWd9RCuMrbOEZkULfEkQsdNS/pW6MUySP6awh
JIkbv8RZ34t5eBiiyoMS9fBf+CLBlqMhF6JKdbcS6Y+x4UcTdTaE0SID6GLAMsRn
an4uxCTVzT7D68YY72WCYSJidUT0j92v6FzI3zye0UmA16R41KrlmfO0ASul+aYd
U0DNXjlrLTtKOeYJh34zG/6Nm9+A8QSm/LPnoG4nQ1k3Ha311dDS5it0fNQd2hBJ
Jk2jI8RNQOMCFtIZT7akCFg9y/96sLuqHPIHjzfi92WKvSTlFCiRlZCOTnA0TmdC
3W644GEaJFiePytRyr6ZNLVeu6hSjtByvAQ4jmz9G5pK1a9V5EOc2n/TLvKlAHff
VrXSglsL857e1GHE48CeV8Wtt0196/utVbHO7meCVIbgMIyoWAi2F4YDCHmAmIsS
hRuuv7+elQNMdOOyi4BpYK6ann1CrFu6mhTDwql8I2YK0+kbAhaDJd6x2eQ3tMw2
4t7ZuBD8vsYSHNk48U+/TPkmmUocILwrhPViqCsypmZoMiwLGqsgTK71LNr/WL5L
JvkOB7TUJ95vufSz0WQchAwvRWD3TmCfAevW/E3GXmKdjxit3ft5pMD/LRDAmQ5s
2RCclNCjiGqfe6Sa6fqL3BKxlskO21od6HCEgTptkklCgYXweBex1cV8zgC5DKcy
leRpOvvWBQz8ulVtHSsEPIX7YOR8zMXdwK+BJu3D/7KSN7ZyKlg+q5f3vSW7ULTY
7gwW2iMOsuah8edzvb7uSf82CYOOi73YLMdxXEaUdVYuNnJbLFa6/CNsrfhlpUJL
mcZPVpzH2c8NKOK9gg4ZHYCmVsRvyRohETvFqXeiGmOQY35o+sgS1Is8I4WvRMlr
IRAeNYhDm6q6hUoVmNJsJkMYK+H7WvQQldFoTthQ4pvC9wH2+AqeADpQ/pHiW2Ll
eRllbEmru4jdKDTuaPzV9S6cUq0ZaaAlrLxpsGMx2ISNUYsbXw5yvdtxw3aRq8C+
ZU/lwAD/jhU1y+SWw/cbjHaHtT6UhIuwS8MO+ZnTT6hb+XMLjYoU4rW8GnsgIS61
s4WPTsOipXbXfcSi/QTXvArFxSspoeXN5K7dc6rLkBPEKt4J3mKdCkgYHkuh/S2F
XeENt7mqkE8glSErEEWCkZkrDupGwU+mJ0FV3KpWdKTOQDNzZ3H9hGwFH6p79aSo
e+9FtH1P0iVZM+vo8I0+L6cbIbMXYMK3cKeNgBQEVYc7MAxOMBRRCsLOkownkD4o
N/JtGjfAwkEhYSmXo7whOyJvMqxOjnRs81tbSguOgJRUQv6zYawXYifZYI/aMoZX
1ChFggcxuWFLCOal5x5IJjsQZ1tVTT25Gwl86/X58gtGp8bvn22xJCnIX2C1cN32
1zORQ4OrmQGzScqkvIly1hbWNOnStPXah9lbDgH83OF2joon0MBSY/Y/aamfl64z
1GzoAUISge4W1B5vsDEPDj863FPhNjCM8kAPN23jtqT3kmQmnEylDwjjMSOxt43q
kvZ3hvaR35OGMKBkzF6EpZlyMDDnemh1q0fA+NeBWG+gZ+7EBfEGOxuDseWOhIjw
pUPI/QyDPcO3xuFzDezUL1/ypNwOTzNzdMwoK5xzTrJ0I9KAqvQMvzAp0HyNdfbd
A2n7SrmTeLClFh5d7D5HGgD1rYWf90GJO3tErnvrjCB8zA39haBdjYSHQofCPs9v
9RE/CZjMiQsj9Tx/klIfiM7abnFN3aWHeZbbXKxNOpN1C9AA3Sc0krXEOTVAP3ga
nM6SNlqPwVOzemL68kbV4o56g+ePQkoE05BYu6NKzmQEWMF5P46NH8sCINNYueI3
pBkVdua7VttxW9aeesW6jG2QkeoIPgk1l/1bt/Vp3DGhkeCpzph5PtQ6TS/tNZyK
WIRioWvo3vmBcC6SXs577/UYfaj+5NB1dT5xiXneQEvC0hOr4yNDzh4qw2XCsT2z
4xiP3XpgNeWwopI3h9BN6JMKN608uq0RGMAWt3C3EQ1n4p7iIpAEjEfNoCAMqWJ5
IeJQtyvhLZF2vA/ebK/FQ0XUHm5BLsHpoKUFW1isCGNOQdntX3Hkqyuc0Pi2aWn4
gOeldZg5KGXISvXfA2mmzQAbiYH0hG0y2K3KOGuh9hSzPGpWJTwJHBSvlIt4e+xG
xLC79YrHTufe9XhE7HCxl4bQA71E5MgJb26nWBoZTZsLE/GID2gJDgAlcOQgL/ue
VxHhBC4dvKHgOKvdcnedDhOI1MqdGpArkBasnMA0YeB0ZO0005AHlXG/uFfDBzWb
OJnFZcfvTOlRbuz9DebuSWyMZOAnxA2koh4x1p9O8Q9zy94deBUYQLqHXlAXrdGP
gsKP2iWJTF+T+Kl6Et17Q/M+e1pygUSMJ9udV4vZ5sTwWCeVazUEyiHjnrjTyorh
ZSd8D8AZsv1M/JDjpmsYgfPWt7es+Ny8XLH6uZON8rERg+xKTW3sAAfOhAKBjpD9
gpmCwCLsrBVn4Nf6k3xqjmOSsAN2kMhKtEMb+po3BioaM4EiyKdWTYgrqqJWRuvt
1kdZhQCV4ihjhnK9J9ZYzqHmrD3P6TMPoY2MAZVMBKm0sj4hO+DepFpufw7/XsIi
IkCocOpC49sW8nWhOpneV04HXnmIdxITjekXVyoDOho509noWBUtk/YEuBP4OTsx
Bve3Il7WZlljthl++tQ/k8i0OzZP/Y+g+TAvJ9uL4PF1V6gYfuCF+l8PwymbKUdK
ueMqqlpwtfgWHDUVtbOOXRLrGyWh0TI1UTJE9Aa8/d0QwDCaKCDrRX93isekrTgi
dwJwa9onMIb0CsUWh4HDAUhfOyZGc60lPC1Ujzk/LI9rfAtRM5wD9YPJkCDYMXrq
lFP4Fo3A1qLkzfCqyKqLNqSjgFrGYa8QjzehnfCErI9jTK/SiLW9hg1NOQCib7Iu
V4gAaQQ6DYGHNpH3Nj7ZC8lOKdfnapjKZm7Ctip9kLcsTTlnGnRQaGcmzWz6N5QV
cPhgxB0slXzWwu4QL1V+RJmXphERJQqXwj7CkB8X9FITsD7kChdKAXa2KSQA5Xmt
JLjNDWIHxwqG7C+OMBTgBCFNa4kVuW8joaTUWCt0qE3ogtD9PzJIEMDz/3sro12a
pztogGOu4Dscok4BU3JOB6yhRyogTSpYhHV2as5oIzPvDjHQcSmSDBRxOolOgZrH
oeU801svmWfZzPzlh2qQxZJpesudV3UtsBk3KErfjFN9JYm8iFryziRjQXU/rYGh
luLkRTwXCCY2IyZR4Lx0LH3iFCcKb7GhLvND1FkAtD1j25+L5x9orKcjDzn4SFoY
yOMfruTycjyitkC4rnGg/MANEYKMD/z5pWG/VxxQYUcuZL1B199b8gjj34WqqYl8
21Ds9vFosUlvcRhZersw3A2aDf3SPHiHjOI3WAzuoHljXtVY9nqER7BviRGBK7W4
WMc2zhGatdtZHRr+gMFgUO7/V52R83TDFTv50TqO7sVR83gb/LUGXp9wYZEBBhXo
U6r6PsKk/WlX4IzADmQrwe4iSX+t7bjy/MA7N8lXoH3FSMKRIhu4+SAJj3c5Vvh6
DG4JWaSLCPUEVuY33rUKVAkLveyF27t6WZdVPHceiNOPlwQVNRzmesgXhtTifnoN
nMvUFKbLvNLDb0gxMgY25G8nUWaIi3iwxFU1bxdbgJznFvsvK96CumeW7PADBFIs
ZQtjquWxtEI3MEZh/ZE8AQtiB1GfrOnzHrIF3jVKzt7DKXnRkNMsTJYDNg3jPlQ8
m2PnxrKRBtA8ODBPAe3cuPVcs/6GGhSPVHB9YgEF+PbqWhSEAevHPAgrgx/mRaqY
Q9r6G1JjILwpAS75fXr0x2NISERVKN5BOvpRNqzVQ2NN13Wn6ZsahakQtuZd8tUS
+/cu00YtYE9PBBQYTQNcvnFkkDkN6rjGJDkZAtA1fjbhUBozAxzAJT8H+q4tgsQN
c1MWa/PfcTC7OzhkVnhw0hhdGA5VdlID7jNVBfk8pLKOtWy3h3tCATcR08Y87GoO
2TkoqZjDWDtKGAgqXS7LRuY9r2esQ9PuRP14ewIpy7oBcuMEHglaJL7jb1Ixehd2
wVYZPoFy/WsFiJwJ+ltgoK5TEYu//CEnTviFVGHbU+8tgqKGqY/noJ6re+PGLVgl
R+UYtxoEliB8sR6B+PiBzCwxb1cd/Otu7uwjIljg/B51he2w2fXY+glkck1ISkhF
KP+5Ho8S6B792ExIOtQ6KGni8KO79PHL91o+aOKsKE+HBd4owNTIUcD6wUR42vUg
XtybG12q3PJlyiB+PUtfck51yxWqIH1srl2mgrzZHu4qxT6dwrTFuz3uRnPEzQ4l
VxODwd72DE7/cHD7okKI+J21/3vyyz66Wd2AIcFEMSeESNITZc95qJYm84nPMzU7
Mhg+xJYglA/GfkGg1/fOUtIHeff3O+4guXiD0oBeaAYarMGz7aUkcT2RghLbwu6G
2tkyxChGKxQ2dZ0wBfNA/FPUiPVdpWHiq/MoLjZXNmyj/lJQVoSz/DZhgHiL0kwe
oZBK0kY9CRXDQHs2vZzRSVT6wbcQ2oWBp0zCg6FXzZbSzxkychdUacV4bVwOpqPZ
giHCRiuWE0wWf3CrwiE9qUo8VjnbJ7mRHNXCRF/R7518bgk/fSGi7Hu2ScHH2R9q
Yu5gXPyEKCOXTglNSbCVeTimfxT15/IDDG4dcuq9UfGE3VZ5flAKhagahDAJbJch
n4Tem7uhWEedO+vNgZvG/s8gIdHdE6BnPvEz8wRNX7ISbAj/TPObFh4t/+yaYiY1
/Om6sffkezDr/LwbyxYpoB/l/HoE5iBkBJKGKvoOCIj+rj0/L8Z6sv/4dbYRLTAG
3UGhDB6a036P3zMRYrs1QMpbnlt8EiN1mPIzXc2QO0EXP2jpPg54qT/Wpse7o9nX
waO0i7kdovLbHiO+IYAsPSIUTd782NXyMyQqAitccefjOmtZxwSw5FzqjHAzJEf6
7zlXdUcBVDw24T+rU3L9B8HHHzmeWYyroURLZiI4TEsPZKBYK2X2ASXLbWTR2u+z
XUPZfU1hEeY1xs0gQSa9SxC35X4tliNFFdHqx9Mgj9O+Ag+FOkT86zEunfyVUG3V
b2P84T+9zywtqgdnk+/n3BxZtteVZmL7I5y//UYRN5Gk5dAA6Pya0d5UBtLIcswl
t9L7jJcU7LIv6uoqIzq+UdsJCoXgScFTmK+KdiuuZ/2JVjWtTMFEoBuFga4ICXDO
to9QuXeVcDLvEyxONsROVhrP/V4Drt/pxmilsyOj9NPFR+vDuItb50lgZSSm82nn
qmeSjIsJW0ftviWCslsRthKN5bmeXBq3DjClKoQDHH2LKnu/l6KBNnMBF8vwjNkL
b9So5+5FlidGemht7baS8H4YxvFBjId+bqqYXFKOzEXB1sxAalAQMy72JUgyyzsJ
dnVZqJYEXPsXBmDKruZUhL6k4ECZjt8eKMy6/3HnmWIAJvLIf7FfJPeVSTl0GJQq
vHpVQDXjfCwgoCwhJQUYEvpJRv01R2i4BXyNAGG0LX4R2kzEtZIxgpk2cZ4zICBp
wXfVNN2TPscniUx6DmqaWG7bC/29B3HX937VUMFVojkSyYhjcOoJTrMpb/X1C43S
vvW7ShDLTx20SGxKDwHuOhTJJo2ul9pwHVgXb8LOUsxPDJ7EQAJllNiXsKTMNCIc
teT9YQDgtWAAscM2YT5b7dvQLfvbJ2U8zRyEkJhe1tVLWGucf/W3hFRRkZsgdKAa
drdcs1gVCHPrzA2BYGnlm6GdQcnxq7jBioyfX1gc+x9TksIhTI9mfAFm5iinWw9e
ZcrGT+TQ/tx6aBJVqD0lyhMeNSzfbV7f6UGca1J1k3o1idvEKwCOS7ITs2tN7CnO
SCAyP74ykpFnqNkB414FTVyxXXnO0cKr29Rb3H3JknDG6/m0YahgHqK/Wm/xJxth
uedFpEFo9jqkiep8ijgbau5+uKAxnpoKRTHqk0hODVf+pXJkSv+QxfUQWVdHtS37
l9j8FtZckVRxp3xX6glDKYBvTsFPfsyQsHUW3AqHjDvs483J2XmSV1r3KGP5P6aS
5X8lLiKdBCzQD9CzjmnE1uKLlqMxt/VMggBiDTCZtpHDy7cqkoubZ+BYkB0EBdBp
CobyL6Q9cWClAd6gl5V040AkptES6DkIdLYVDrLdr9tqGfX5+rdWlHb4K5U6UoRM
ABjiwuHp5e+L4rdF1XALUpWRs0sKMa0+CeJL1qJnlF4Ym2i6XK4eJM1EYHKkp2Tj
UnMCgjJV2Sv8B6FLs46SDDn4ndM9RoiTS5zNuALVnOr2JruTP+y8TIQwGz0NxOZQ
9fDns1r4q+z4KdG5d7lds6LWsMqzZb2HZtYLurZP7h86s0Tkg7S1iNvbhGqqJ+Fg
68qzmPBAsE99T4P26T83xLuJr6idBEMCZk4AfXQ1uqO4RRa0FxG+hPn3U6leKeSB
SF7FNIhLXA9DrnLwPnd89JPq7gYHrOjO+TUywmLKJ5nDD5GCf2tcrj0DFng5xBtu
yEkKbp+/VevXZKJo1Xq3A+HWLvvR1scbXTeieFXcsMNbB4ytxoaYS/k5lSnRnql7
BVvMR/bNzzWxpEdDT4fbwTwRiN3PSEsSMKb1qsTG7sVFGBywXRHAwI8rXQDJTSYK
8SAiQYcoEK5iaScsYcI+PJS2LFIzDTchzhPnQ6YqwNXtGvJFP2+XbljnZ89QtEf2
G4bKsSQrQZAxYpacEOgu4AZmL2F8x2wEYHsENH/yn/zsp/d3k9xlv0cMffTKbaOu
FmH3hCdRXkTaX1V3fdfYqfP06f5czj/GNLp3kWRxjhETj3+DLQtAd9DW1TyiIo7n
sJnpzjkjbKxnWHpHvM4D8QpQZWwGLAdtHxSTQ66T63jx6o8CjDCjNHkZbEfN88SG
x1XOs9Biy2JhZcYZQb55ecKMwEVoVU/52eHz1w9XkAZztRX2Tse61RJRlgODdBZo
/Ohb2Ri7FHUqQjnY/ktL8hOX+GtxDZ6YjuD84ovLVW6C6pA1+h8K4uxDW0xViCYX
HWHvLBmOJNxCmESdTXFr3Q==
`protect END_PROTECTED
