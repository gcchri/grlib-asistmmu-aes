`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5q/ZyCChzaTaJme+WZTTPtLsoXCbn52e2J9cIKneqBWLp7iKbSdcQ9aesVzcKvTv
uX1J1mFg0LDB2BDUY9zlex0eODsJ5JLf+5PItsbrK8hbX7Y9UoX+PcedD1+xyTIA
/htGshpkxKycfxnTDblhX2v7Kh+fkCHIMHbXMH1r4W7Iuoe3dAmXGuAf1ecbz9D6
pDK+s+2hzcb+5H9L0bol/ZDTKhnt0TuSRi+cmL7ioqwi+VHeTtfGOI1uwwLxzUQ5
HwZeYhkYjYo/guz1pPeAtZORfvv6uYY08wpSW8kRkRBjThUCpkSjmWtn7mr1wJ9J
Itt38QC914Nk35pYjzGhRSECxAIAT6pHDJd6TakRZtitaBcJdYQE614eEVmnNpJC
pKS1TDk3GghthhGsIKc6gT5vxBgd8kwTewbvL7p0rGg=
`protect END_PROTECTED
