`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+jh3bK4RezNCNfc5Kn+S9N7W1wpwBFLnZ7hIF34Q2V+pmySlqhwJdKnAromuMAQs
DN6UwNkgh1mNhDdjMnjo3dtpGNrKU+UZ3WNo8G+OVHrNudiJ8brb9IVmIsKxDVyB
rcyGpFnRsed6Vp16SDq8jiLChCqf1v5D8ZLIFf4twPE3lTCSnIbeppyfZR7rjAcA
DOiHq2CRifMSUVFvxzRTiHcuC84dwYWYx4PLHtkzJiSGzzetuN0aOD6/9O9dXP1f
ys9k2Fz1q02bfR7kYTdrAFD7axuHZ23+vDaEy01s/7tzGii1qFT+eaO+34v1xsFt
BkJJUWCTOynd5oq/2vcLOmXNfXjYOmSmxdi7v6Aq8dpOGUHxC3Ab0EIsEJPW36FT
AO80BFpMa6gKjwvOGuofSDdSvoT8Roqov1I5CbX9DunyRjD2mVxMzEJqzLXueMWa
OLAW5qP6YjgtY8VsudiTrz7Cjr+bkTaNOcfMX0WEWReEvdNNnvdW8CV3GRdZmILH
a2Vv0O1s/Cp9X7vynS7vKjv48TiBZ7EAkXFfoF3utvyjE9VNnh/INg3Qs0jaX/hQ
sluHqNo9/99x6KMJ0SfZ9tpA7FY+Vyx75V44H6aLp24jffQsFKHf6/hn0Slw2Vbe
Wq9R6awwTxPi5h7B/+QEyag9pBztVpVZIcZ9KAIDg6F8aVPcKCf21Y4PL+w8XF/q
WA+Yz7XWfZ1aM9wAStOqR24FidYG3JVkoGOvYj0YM1THksWC/z8Zi6x15dOKohRr
DIaJqXClIPyxte75IVeKdg==
`protect END_PROTECTED
