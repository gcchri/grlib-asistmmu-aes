`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GhzAznT4Hq+oHzXoYzZo7INYZEs1bS3mO3vQussqF95ShVoDw7VMhShiO1o5wK3q
mu3kDejOwkWBUNxR/1IdUFvcNW3wl8b0dhCtH8yylP5tv49FYsyhVJH1t4nmrTen
XVgzamuTaqq7Ua8usuwHFusEQxJZwVfA4OIgx6FwKjT2JCjwlSgaAboip2Go8NU1
SLylvnXH9h4CmRszO22lZY46rOcyzHdUjg3QmYbQCWVMp3vrISO07FYuJgUgCMso
On0v9I5hQ7tTkfOV1ctAA5zqevTq2WTa8/e5RyLSmVkFRppiunBXySEaFqrUrDuA
tJiUfjlCwW4+qG4V6X5c0GT5zaByV4+9EwI0mZs5E3siR2pdqih1I2UYWWDH4Bmq
BK5bnqHj2tyfr2r8C52TFkqOHUIOCrdsQ5F9O3m5g9evc2Xcpt/06rocpMoLkMKu
FX9xNMZqDTHAOVWWDtl3VMma4SXYdZt+sSO/bMuoRVBf9f+oCS86SC2vgO44kb0t
bmCxpeG06hylaVVPcvAHp0Fgff/3lLvgWegPeDomKDLQU/bjpDpbU8fg7bw6fsez
fPFh05nwBIU8hGK3D3udv8Xkb42FJbqElbDlinEwgGo=
`protect END_PROTECTED
