`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9ylVxWhJkWs4ANwqzlliXQSZChVdUTVov4g0eweuyJ0VflSXqrP+gKsUjgm4Nvo
ChKVKZkQ/FBJ9VQ2kgkwpJeEdKsKLs78q43Xwke3VHSAEcS8q02p8uLAhtLoq3vW
hQtEKVzFBmgKvumZGhDZK3g+6NcE41pNx8H5e0qzU5OBGwjvH7yTpV9Eq1z5AZXG
X9dv0xYNOso6GhtOa0sErMuVUYWnj4t8OSVs64c4hPnCl+xJ3pYQ8nGe+NmFv0BV
Ol6g/9lPeT0EB7iuuLUvU25zfV+A54NBnZMeSRUhM9SohsoI4Nua8qqZyQEFgDOh
BKD2YQvQUtof2eyDohExzsNXHveC8a7RILY2C5EeHBSk2+z3rPJ0d1/44DlGafmy
u/qeWTSzH4pdqg5EkdU0M4wM92S//x4+80SzzfnVRrg=
`protect END_PROTECTED
