`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a5TY7/U0Soi5FV3E+NlS7lrkAnjFTBZe7qRmb4KOtfEs0OAv53vvtF+SYINVXH4y
AIcERG9gJDI7Nde+I/YxjZlEiDmoEip041wxTPe/zJe+k+DaajgCVzd5a+3VF9L3
BLjd97rQaxVXvbueMCcZW/l7PQn10CgMka/fYOj5WOfVFxqyu+xwS/abS34/J90V
xIvAgUqJM2jFiyat6S9H0X0ePoN+OuwP+xeWVwAKYGiM5bcRmXxxcuzsQH6Yt5EP
Vj9TkmYlzErCQ9XVFX95xg==
`protect END_PROTECTED
