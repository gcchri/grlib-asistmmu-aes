`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rpFVQIK36YLBSXxvCwZSYlvTLY2cVYjgxHxxCNW1NeVPyAT8APfJllV4YEfqVzgt
emcbTkX2qhWU8C6PmXEhWQ0jVrzJVGQqyVqEabCWx5opAezTEGdYecemTcHzB/tB
gWzB1DdPIBxxT6K45oDDQo4XIIFim4IKZk/yeT6ebb4N0yy5/zgwZdurazWKgTDL
8/SCaT4UDnKa1SQLyyz1XOF7xae4eCkR2vCnhVIfmbFf811qd0SYEPwyURgHRjXt
IY0LKWWokDFmskPnyZ1QX9vzhuRUgPUGU39i/L1g4zPblYx+WJcOPG5q8PFJYemJ
ZIqZI8tRpFA1IHyQORDST60v46jLLH3I47mW55KlTzQuvCFWMnIGIM0eHpXHkmAx
yigEIhh5qwZeARy81PYJlddCaXEu+W5iJSrLPOZNcgAnPUJyYpneHXWEUvCvtnfa
zs7owoZCyLdvkQO0n1NCCmfTT9HYMEOAxqEPqHAu/b9x44+ULK7QAy50CV0sjSNP
kATUETPWqfpw9jadjyNXHtlejMJPpQJTx+XMtBpRgnR0+izlhc34cNg5DxrNN4Oc
t6fsPbwIN1A7wpCCZLOE1N7Qw7zQ9T7ppnq0EQWpj1K04o/pnGpysLKqMDEbMmHA
KCaRhQqnfR6JV7L631NVyTwqQDPNENSv5sBUvXj1ThpmVYzzp/ucu6TFEGE04lnf
61pgnQM0WYTlB57auG2S0mMQ4y5pgGmr2dUPczhl78c=
`protect END_PROTECTED
