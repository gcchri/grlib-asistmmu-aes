`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4naX/5XcqGl82TkC5AliEAhyXkXUk9z4JcyTE8QvmB/S5mYIE7wabJMOrLu9TvQt
fw9T8PevQy58HrLHVHyQuLtyB8vyHV4I1REFM9eNqGkjJ3rwiD1dQFMl0oYU2Bdw
z3O1Pt6a6xvz6CH4QfzldNcHKmS97TQ714m4geGdc6tYMVHiPka8azlBmq9gAKPd
8UwS2AwS0/QxTKpCocUm89JV+7Y44/jGX0BubPEx7aGWjTDpDwVbdQyus6H/mogz
vL+uhwCjpb5oc1T/4n3LX+WHMafZshe7rqkd1Ye0kkG8wd7oVGkjH+07ZUByEUa+
MXLu3DSeeWvHAMvc5OG0z/ZHKJxlafMKUGx0WM1dTnKQADtwiSLs/l8cs0hk65O3
rdRITdkYsvWKAPzZsILuLEkyTozJll8QMO+a4Deh0E6Vt4myFj5E9oUOTG2mcmIp
89B6gX0acjUDLn2qF4H+DL4xjtZzPq/KMFKvsvt+KKq2/Iz1bbE7k7VBeQrXinPq
mLxGtggCBpRoZtaeHU/7adN2sBxIxtho+7dEdpSbvTYOxVAvyskHYAY4TTgFIdO+
MvHum/KdbCLSagTFdhNkwWaQmJZ05/ZaepErGoUR7we+GEuB0kxQeGuvDLch1SHB
eSO0AW8eQ6HlS5ahH/2OPcH+x0ggzlLfAx06eX3n0ywmWzIbErIM2xYmBaI6sQ7O
vGRgI3UwEZxxFZIaqz4udb+EF8WLTz9Fxz2IaGoqH7svxySg22M21Qx5tdFkVdIH
4zxJMnR/mf47C+RnTWZKhC4JCqO/18/k4KJ9VLU8Z9vyiv5J6HaDsKiE1lsw6HTR
IFGNzRAN0+OFMeSTl3J1whg6RGuniBHGYak5lC3Fgh/WOqGBDO/0VOLJeFFIvYmj
1LssPbkh3ggWpWx95W8dKKhZx+w88eIkIeaaBEYPUFYIrl2Opl0HbMD4LDK7zq4h
UNQvG9T7pGYM6CDg37MLfYyk3LNKq/Y2hmObANHVDA9/XyxPSihNsfvAGFSx5n7J
rmjahDwO9DZRpXhbduWWDl/4yjtQ2cx/JmUvxvhoToiejPcz806JIdZQAeIzPOSp
d3XuVNW4DHJmfERDN/JTZnHQiM/v/KIVVxU49aBKYrQ5s0E2fWBK6M8nMlLg6Op4
2WujTQhbS5isJgtw07Rqtahx18qYDBzuj9RGIZmOhALEB4gOOWcQ4CdGLqx95e3m
OiHH2ECDCFUcoJ9MSFfxU6/nuAIxSqG9hvH69qkVOp8cuaYp0vB1lIFM/yFv89Ni
kU5DNzhJCjZzIv8dXbBFSPS/A2OnWgd/+YqGM7gW+C8BoXZfw3LLwcaYx31aITkM
j0nelH01a5VW2JAFDkO00gEYL0i7+GKGWF9U6jezb8dWb1NpT99tq2HfKTbRZ7ju
2d63mnYQHItYpceubTMXaN6DUIaY7pUafWwx+usHTquV0GN6eLJqL1Ka5goq7YMi
Ng21APOn5I04CCQ1cgm+DyfpVi6wlDf8obwGB/jMNMttAXOVhgDfQJxTpKf52m1r
cf6r4iNEOmb0kiEKiUVRClK0tmhlVtri+EFKzJOUVf9SWU3Aygr3iBvi899plVIj
Mdqx+utcWtXYwuA5n+/II2BX4k6WgD73BvjEs9jfzYnG88w+yZ6/+av1FYfEjalz
XP8zUmvtAvWEQ2JUykKAmJRon3g/ZMQ+7eMVvuy2k03fP0pPsULp8jGbocT4ibuY
e9jfLkfcU5X5axxpmDNooDUTsRq0I9u+GqqFLLhU8+NiwH9euBWhPlC+KuXXtemV
EPTrEK6CxRrA0geIy1AHp3ybMo2enJDKvw/zgHblD6ad45ER+Gv1PxX+iAn8fkUm
5d5dOhgATKC/rGaVII3sQPuVGfnA+viWXAE4NXUYeho62BbzQeF/Dck4UUR4q3nW
wAYmjzaPOZpMZlc8IKg5w7Y0PWX8Jn3c8RvyijwB3Tc37TAesm05ephsKhRMAahY
NoSlAdRIgE1M74mAeX9cBKfpY60BKMcgu0SOnBkeT92PxGsKN/PxrFl2kb3+H7xs
i2vp7y+stI/wi/ZgmcMNpGwMUjkISuTmpzkThUW2aT6pE1KGEV8kPdcoITnbmsbN
+D7M+JP6G3ZNxHzNS0ivimeTQX9v6bkBMzE2MAY5+Xo3knTRiAz9/YEk1QutOl1T
cDcxrj6GQkSsIlFAAgF87qL2J1rpyrDkf8ZlTcPZIx7DEe4VdGkLUIYOXbaiGlh4
il8HgwVjKzO9PNZyHiGjiN8kTShmNYE0/mGvVRqcIVZYNXrlHBmkj7VU9HTTihEo
4Bnkpnprg8DlzNuvprBeTA4+BDV2OEMiE+YP1adpawLnphvylv3iKYbOdKMzS0mV
LzayWp11L0JKobNAEgKq3rKnW2iOutZVxp5nS3ZYGMbDKDF44kJHmWAdwlycAFUp
ECE4aYaR4A19qYSL9i7ewvOe3fVPFmkGOVR/sWiS6RgG24yoUy4+bf1iUUIPaYzv
mGPx2MzWXspQozvRXhHEMABGq5jm5hovoX3R6xMmK1hrPp9cLavL8MCLRRSuxnKy
DLD6V+7mhwMRX8mKQfSg5yZjbYBsSQTQSomiwrTmX4gqDcBNu6hq+5R1M3kLgeHm
ggzhpxKTTHYSwn7y1gs0xBKLd7DhFRKPHiJygpWC2AFOzJfNsQRGW9zRz+HQS+7D
/rTaViNvUYCa5/DQlNBoyQTm7ZUJwCLEZchypnQlw6i8+b8/xydprTAiqjA8lB3D
kbCsiu3cb2mld7f47bObVfmj4zsrvx6kdsG9yHg6ty+RjvnUDIclvR+GdxDxUVBh
1+YCymsKf4weiksK4nfcIOXBFjZ3EN8LPSoMZyo6fdMn/Zx4RDxpFyPtoGt3cmo3
JYa6V0LDGMFS8lO/4p8VUHTdpBurc/tUfnWxD03HXuc54ET2eL7mkvN2PiiieLVR
leo3WFpeI1+s8uygxRuf3eHwNVgLgIdZI1NYPNnF75nBVf2EKqLAtwS6NowJHcYB
1ydXbT2eooA4d7Xsot5RTEfga+DX/y2k0OgkjZwtZHoDEGNTJr+e6vNHSyzKxKvn
xCVFc+MlwbjvTc8GTk8G4CUxs1df0Punkp9y9PmxdkhEruIVJGMUkQ3aAMA4JIxd
P8CyWv+nAIMiIsUWZSWEuyXT/0Dsg1QiH/mCA4RUzCcMRKsQwE80EzhO5P/SVVeo
7+zMfr2N8fQoigpo98R4WFRniqnpu8k4ELAHCAW+K1J7YEXmdCBIuaTCE5FIqY5G
Amrr/duUfcZjFFvZ6mWVR0gqbNuE8PvGsoVBl2NPj6m4SZPbC5rBPYgc9AWRgBQB
SZkKF8fHLPkV6zo9f+7N8zNRjGBTPihamKKiQHItIjhG7CERmB/TqN6gWkONt9x0
y8yeCoH63HFl8QxHOypzq+ueucoaeh6xDVoRt7fpsV/iYtC3lDEEpi34PraNCelm
feefvWzAMKUVN/94Chx5WST15Ggrdy45EgqwnD6WflUlBmq+N3S2EN8PYqX0f29m
tQvL+/4QeX52GhNR5Vh92TUtXJ0V0SXwl8RHFfi/gBJ1rQvxDaK6CQyQjGtRVone
+ftGUcExswTpMyvdz8fZtePAs4o/bw42gFSs32K5Hh3NOt8kGlh00gU5pABlvMaH
VUuugc9oSHPLIOs2pX/ycROlzHVyOmclg2Ny4PsGsoHcilqSA2pz+uibGL3C281C
dhlA1ZrNdp6A0+cwTe9fCoN0YDNN8W5Lmw4nj2387Owaw5BU5GvBGP2C6hliS3X2
lf5zp1e3BTqhMEyzw6ulBEsF2H3q9JgkKxpKlN2kvubbZ6bA2BXnoSqtJrUILA4R
m/OPsCXdaKv6mmiVlL0x5dgGn/o1QqUy6mImpcqaM2KY7ETx/GLYtqlxqiQBWG4W
3QEJAUJHbT1kL2oFS5si1fnvaRli3ivhHN84RPXXl0O01mGSYOg9GUf83yYxJRcg
iE58q3lSFMuZIbI0E9Pc6aoT/eFrTw+LnzN3TOe81puMRz1jpSYtAONYirgeeyJY
q0WalZkcJoPWLwuReA1duSGk5WrnK6aKOfmKxSM502M8lzjueY1Bsw3V4R9Ex/gT
VrS/qkPhBTQe8fy7qcOYecDv+EnjC4TjfKnBv8e7ieKzBl4XmTon2pPHq8nh0lCE
7KRz4hb6nRvXafa+Vw3HxdCra3o88eKyF60vqx55LnmNrtcAiVrhz53NF81GwfTT
otBxqiFDu9ZIvFIFNtownD1zXQ55adSC6iZxKodMR5NM7q+N1XL0yWxLSwB99RgZ
2e2Db0RnWiI2eKNOIa+9vuYWNu4bu4S+I8Jod/bG244pge8WscBiE9lm1Qf0/rea
yX/hbX5ydjUCBew97TMxkS43+lSWMZm2QYCbqWlV9lE=
`protect END_PROTECTED
