`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
01UabDZtVNPjisyiMbvY0qitDjGvLmri4gP0W1n8920Okp982JM20yktScRGXQ2P
L50xQJBMU0ZAOYaf7m6/lDh0l6qfO6HOYNeZ43qWRSgxcNVAVrWxjFDmWdHPdiOp
+ipOfQAb/YU5445IOgQno9l1VFm8K9ZkeBkfteQtBn3loPa2TIFXsvO2Os9HYoge
WBRjyhz42XjyNsGS93qE4zdMsEwQsCQLHOl73LMN1uu+G5rJEtJ52eMziapzt9Hx
SBR9I/YJsfTO5BtlanURkvxwfTwmW2RDcr9fnEfFHyWZvylvy32JqI+xHBJ73gcS
k0xHoQQaIMZ1VAFoIWpfg4E4sUX6DV5Z1uFvQiV9Nt8oWt3GOJ+17LoyxYuECzB5
+WJHq4WM/b3SherTlc3CQ2VnZKA7yaPSLuR27nAFkjzxOC5EBJlh1d6A6mzgGHCH
Tb1xjV0+whmzozYQtZyUa/l7VuRhYCmJWFY4vpmbjbxLEiPKCWEbNtHM68P+ajNT
y7SH/YVzPQk1/jofL4eAiE0CvjOykg2zTMZAgHlJ1e850HUO0yNntOY0dPkREMkA
/Rkw7mbbAQrk/3GGN7PIt/vSYcoEt/AGKz5YY2myTKbGv+gUlTr/fKGz+G67yjBU
EMranD0or9s8m3utgK0B/i8Ef91RAaLIMHg049i0dAOafXAtc+U4uuBCyafMHm98
VfpY+voTEiMWIowaAMIgVjQLDzr2LfzvqEPsMAWwnFDPvEVF9SPCJxP3LEObC5rK
9ZFkhYZhBFrmqLCDXY17Kghbef/rpIUuESdg+XyOPjctRxL0dg2GLfRfHOHQf9VS
ei7bonGWOZQXBZFNh8uioDJxh/eqdRWeypnVdYY1Y5wZIIBcFzuO635lYt98U6wo
l2NKzVU/gLMIwxzOM+HewXJExAdQJZXQ+AHnBAXU5JcEjbEZR14zO0TgjQ5VvWHS
3kpgJ+hGFsl9RP+8+JgKOy918O9uUkvcwQS9ubSmDUTmbhQLpeb2PrRnz3r7vuGn
TqPt3AsOOC8RG4u9pUUIlSYiMEMSPRK4Svotn5f7wsIbcODjKKzbQlNpGW38z+bz
lTTSKuAMtEs16KWWiZnck7c7RqxZK7jfnNw01vXRGd7uECP0J/4Cl5C9Nu3JEOoF
NUY5q20vJHceHtbc+wMs7ODxZy1t7F368PYtkybFAhLwXiCKtGNzPvLTh8SQR04T
P6woX8Qlhg2M1Rp+9MIun9CwfqJTsBmqwAhcWw05HeqXD2qKgAQDelrWFNX5q4vW
wK+Tu2M/giINq9HOUTSJ4zc7OVXt+db8POggQrIWEZ8/OIZbVWg65SrzwJld8+/h
9wXA+3fGOB4rudjLAXEMGcYMB0lGxiBk44mKLrgWpZKvSQL3lJyNmm7nO8FLLBFT
jhjkXZbZIYwWzHKneQSVAN/Ny9pGQES0EORXi9uEn/wfruZReuNSLjyTzU8r7ySQ
NXtIs+WCSlO3et41SisRK45WjGuJt37vSE5mSnX8KQnHgDOqKRXgjnEbeixZ0aRJ
kClQEiSyWb9xhTe5adtz6vTvl/czCRJdcgbM3JlvvRjWmb4dEvJVtbdqAgYLYb/G
E0lh+IbWmB58xNCNBF6UZuvQ/tpynghhdo2LtsJsRh2rfRFfxxNCH0gzcNzZIgnj
xTq7yVsIytpc+dLyHsB8a5NFQHv9q/B3mQQXuvLXB1RW16qpR3zRFYl10hyr0LWx
k5WHyiyHB7uHh8Ed3dfhTiUGUjVTKdAOUe+tmVJPKyO7oEUm9S4C3rpXVrnp6tBZ
2o/6MD/SY2+Od6c6usFKPy0t0RMjYMP/wT2mEl9+d3qMc+VX1Vkdi/ApTfP4JJWd
xxIzfoaYY7q7TvP5n3Q2zYwSBS6bC/XZwqBAYNWnFXslfzl/sbJKBuADrGHawYgq
j2xaCd6baWTbCChJOsWHnalNjViHlaNPSOJj4uHUbiLcGWV5N35qZJ0B4fKSL/bw
NtLFX7x6u73WL56pcKRCwtojlqTviN75Dqe4QB22reUqecKgqhNsaYX8zOVZctTo
fTfC+k7rfaLt6GkXutgx4ArR43SZNdXs/vQJVpA5bbx3l5wCmjKZEmyUDuhT0leD
JRzmrvXDvH9ccmypeErauZeg3kv4NyHCgsezAHrn8vr05J+1M3GYqOKXCDB1i4kN
iwk3UFmmlKFI56rzKXey/voFWkXs1fx3E8d6RIXfpVxLxRWj/RPNc89zuieDCz7W
Xu+f4jI37egGmgRK/CsDYiKj12/YvERuloV2Jq0ZdcsxdDRjXyYDfWIyzQyo+TOH
Y6UmBPFMAZQZbS+/WW3qSp17+sBsjha73a3NV9Qs7CCvKxzSlNjrBBYApm5VSt6M
KVwOc353K2e+joUY7WJvCl0elwkYyZ9k/VL1yTXARw9fQqiKWVc12dLW+SfPbd/i
fFle/mr0zA7JMa053+nrHt5cNNqoBzCkYEH/LfhoLepiiy484uNxDg6i2M05ESp5
GyTOPmMHr8No6693Nx9dSVSkW3Jjh54P75Xxo/L41Ei8ajLEcWQBa2Twt0yS4tSv
FFEInq8wGS1ic8Yy9TYM2Em119UUY8WBLo/qT1WLLbxhUJD+4wN6LgeyTBK5WkRB
1ONqlYZXp4/6MruPQQMX0Z4YKBPt+Lr7+/i9yWY74Y932KF79/2re0AlRZ1/S/0M
x0DtBcA5YTfxaB4e/zPKi5268n5WUzV+smA2gATkjY87N1gn3p77sk5OKkk/utnM
c9CXjXsUJJAl6jNF8qoTI7B1Zskkn+j0JO7QBhN9mr8kFhzmsQjCj3/rdI2s83rI
4X00sbAcUuXnE1cEqx25TEg+rZmHzUY7a95FR5p7CENT57rF/lRAXvpf6VmZrP8A
eY9NdzR7HFfyLv4K4KtRDZuwgkAkoW2Uw2DGHhgxwyoVKNRwtnUjWjWkunsuoNkP
ICvvyqhKTpChG+N+00mJe0aPwXRTmxQwcrjMujcmaHIPVBMdTQgIOD3ePRQr2g3U
qmEQObN3TsTNugzRkiOM910IawEBpMF6og9L3vmR8mcN3ZFKfGtjWZjV7WsYfgO0
a7FF3DDr7INWiQmVvBh1gpyDoo6J60xTg0y6hTegnQ9LKaTg03VVZzzBnGoH2FbH
4iY3emM/ZzhmYZwa8e8vI7CB1Jeu5vUGkQkkFHfeGb4LHLwN15yVQJc937gTKIf4
kkod3jPeSqNWmgE4wWCBSsfISoLWAS/BSt20/LtYNebrWLMEdTXRSd//dHFa9J91
BDv4NGssUsO71s83QUIcK8Nd7yEuEu2NrKbWk+6MIYXjII4iVfjoT3Aw35ffzjMQ
QvmyUGO9hYvWIwQh1vrYppPbaMnoULAqG+qKUHT6C6c48/2jKoUGraXDvlWHX5+0
cDBxK7xVO6eqD5qxcMc2XLKe2xR1zKBm2i7bpowTVEWlt/SUxmqxIVv0frPSalia
A1SpLS2t/KTn/MPXaM+Gel7dU/Pl0HGIjoKnwhATeo92ck6BtN3w3VpR+swkyuuA
AIwMPRYweo+WRfPiM8e6kYsAzLC1emhkvrik+j/5dCnhUqs881up1aWPqGTTXpYD
ymEdhEfUePard4OLxgOcGWGcOXPyIYGXv8cJfDuP+lbSace6zrgVdgd0+DIG2iZX
ni/aTmD0VXYGx/NUzdERNliHa329vm+c3XYgZ97CdTNo/HMT+hUHwLb+KJj1ymT/
J3ACiG6GidNSFNzz7VdyXaY7ahgNL8JlW04b0PVOX8cOQKgzo1CrEzNyRpb0/DRg
BIEPAZB7ZID1uT7Fed+TwQRrHCFeuDbBzmjrVVcp45kcdKAzcsdvzA/pzjIZ0dgb
Az4tcViIcfQoruqI/WlX1IrgJkh4LXbixMYEvOhVakmY1LZucN6lRyWPep8yk7tH
pRnapUjCd39Kt05HPgCTs33qAYLVlydwYMt/cZzsTdcMbryAbEwq4Zd+Dz8KwEss
uXb0wYEW9/tYSJjZGtvM+3c9Ewoa7rEtIi3PGBHhQVPHMvwY0FjxyWBgLeCbxX1N
m1bQCrOnw78tADqgOaODuz2j/KD9Y8WcoZYz5F3c7jO+3fl2Mx5Kys3zrFIC+WIt
ixxErDv+LsmAwNDzu8Wddsj7XCI8pGOR6oE5n/3lGCr+WgmRSpbGLrs8l1GzfjVH
xZp4/8HLllqXn7Uo/sFR8aqtJxltdOrT9P1VcQ3p6HSQ/taycjqOMUP/il3jXcYg
pEeVpjQNqhD/cS9MWyispI6PIxG4c17rdGmhlzS7hSsHJDSSKY7sn2IP7TaSI6Ty
w12gJwMLvcPdSMJIcyej6LvocjFGYOb1wIJQT16JuR4POFDQkt4I5G/5PQxDpUz7
BPgrsuvyODnaDR5rECW+2po2nbVzgU35Yy4+966+rhEPnPdg1FhhcYOqlN+iy6Bj
bRl/AL/5ORWJCGQVC4PjUDgYJJkMnhKItPdlIMTZnUpboH1Z5byKpJ+qVgbwzk91
Ik3AaSLXxZNtucxHkDDMzxFRzJcRTuMw2/6y0P8SDwiiScHnOsMNrwo95W+5A0sN
/6ZbyUAZJ8dcNOOJltwq2aUVi3VH6gDXvCO//gjvsxzoNZjp7BwsXtlBz8lA6buT
ebiZRDQcP1Wn7DIeI5neSXotenUk//+31URyFuhVxiSptKoNOpwRApPb2hylhQB4
AiX43XUGDCLCsFRuw4LtLu9oGKHC0kqHen0WqL4OUKKMX7oIxhwx2iwF1SWwX3W6
UM8zosa8FXjqXoaC5tdRxF18u/MmZJewWBKPv4f9KSNpmg6V3QCMWnn/19Y7cD8e
vUXh6aHUsS+1J4urR57wyas+1qosiKm0BM9W7f1aQIO/vm06XRucvkshPRyKYs43
FHZaJ338Hg1MdvLJkiUWDuBwxkjoLGWx9ltM2YJokMJfrQzIiMQIa1SplAWc12WN
Xo9hVQ8KhVPenR275NnWsKs7ziM4MCh6d+jJ6Xha1+q+gBLfhiSiNGEVeevUyQj4
HsQ1AaEQ1IOlIP3Aq1kRcPGG/MsbmNByrtKODuyBvK0YH1skkMOGRz5njuH+0d3z
KpoXcEO1U2qA5ibssO3yytXXUiG/EGrLUjdTPueGWysNEQezgnoix6j8gWCQyuHh
feuQa42fjbkf0hGuW9roOd2yk5GbqjGBCiTns2qvI+HNpp0d8JV3SERhkaK3VHz5
de3/i4GJ9FnGh8khuZoxvztD6yv/BP3IJj2K503s8DwGnDkkuB/u4FoSHwyhQqH+
ZOkyiwT4/rLchasuECy5r1O/yizbzECjTc54xJjOv/R2zltGtxpeNe2aj+KrRND/
qAFELC/XYBiNYqcs6exFAJJTg8C2ghs9NJ0I6MfuxTRMqEO/uoI+M8p0tWcHeIYJ
qy5UiuR4tQcSsSL/LNUYNHTiJNR7E9iFLzTwxKcWbz3J6Yf9YnmeBZUW4Xoho9xU
dD6Co8HBDQrz+WB5puBJ+xsjDiNn1p2l8aXhYYMlCUFCy9X7yU5l1YVEedNSkCiW
x8/WDthMrg78X5YTb28SY3etto0ssoWoiIqd6pqVQeDGqxNXUirLnE7BvrIvlLhW
oxoHkMFiNFK0CQne0KIwIkVkBPAvpvpx2/vX3qhsxZkwMAPUPF7gvzepsDfLqktY
ucv0WDegRFKgi+jnaOypafFXIV6RbBeSfyAZeZPguXy5V+HwwdyW3jzwgm2ojc3B
vgWLIoVPcnLGs3VRC4yOAJHoOQa07Maq6KxAoKxpiZQm5RcGoc2GAHyFLMslf1IV
YbvY2DiN+sfsgdauzdBRkLLUh8qfgDULf8TvOoVR7X2ywgZorgTFcz6JrqdHrHqr
HZpTk76tLk8WpY1eMFTVNAK5OW3FY7fxP2Y+w9djBsY7SEOBfLx/DrAzG/R1G5+l
1OyX13iQYCnFxaehTqb9wdY8AKRsm78buIvplQNOnDVAfe700jOttkVe8J3vU2k4
Rml8RxbpnkqGVp/qYUpThjNg+JxnGPXE6cBa7yVl2eZpuvt/26Agx9Ka2sY6KDVO
rukXfhR2023+gb5BFX78Wf3nUQqTF/ECKYIgrcSfPOZhox864sbTcASvbw4KgLxv
0htTAbskPGVGnd2YxgmjjCntPxlemIOCYZEzDRjzKb4pcbYGQhyKHeR4qNsIP7nz
YNtN+mgaY5sXK5a2XSU9Ft06E0C8rnVohOSAQm+497ZRkLKKMpm7+45X5AyEx5hQ
Uq2Rt1k0ZtdRi0UUGFV5WgIPQLG+CrgAcCQNCvUJTvx0GATeDv/wwcsAu1z4MFcX
hUqfkLCIUd22l6awtCyVBat2Mfy+85P9HQkJADOpE7jqqxppQCL/YPvwOSxZHYoT
y5ubPuYW2NR4ZQLJYWgoSrlDkjgqrjxI4yvZYpJHXQgpIMSoCOfj7/CqJIBBLun3
BwDAEaxnsP0HxKLjHVRKtXAJIBse6fZsgs6RsK2rnfIS1QnSA6f5BydogoQYcoie
zQSGHgeCtMjyPWmigMuGQYpJ1WDCNQT8Mfc6peE7Rq/fc/VrDtXir9/kgva1stuv
1G99sVs+lfQMzOGuuMA50wCgPqO8yeUQVeQ6pKs1VkaiQNYtkEW3n7vyzHCeqJsw
SXgFWODaxZKpUOE0FVXofNeqGVwK2dQxhv7HHhsUUNF7y0qC+BrBBD9qnw0bgv9C
LtRL5B7GR3pkbKKGxEZx5QHQ53Z1kxZFdpVG3Sx7cvNIHwZIMPxfbiB1zEGWTV1U
NZF6YdzPTgRwnU/e0NOlKHIL25Zy4b9wXfB+AefVWi178E6OC0TZG525N5VPcnSG
u7oM6qdlSux9wSp9dvQvzjAW5EmgYhr1InD+tFL7d+ClxJa47ezClrLTZb8foQqz
iMe03LvmhXgQEOKi3DGazBla+/M37I4oPUQa5V6AvjkqhuSp6E1yiVdpNPU8gZzu
yFm/bZYJpnxuUMNMla8mHUNfGBV57qu9iru+Nb69s4zUbBQGOqgT5kQExvGck0gi
SxbkB2k5b82+n6WxPuU2cuB2f6EdknPl6lpyQ4GGh9BVqdZvfBJznSuVv38v8gDQ
G9/i1Z6eRqJ31eyxH9aZU02b8RJ3/usqdlHXKMewZpWycSkSSQebnjkHCyMBi1NU
QtxHHN2fFfOkhJf63NoVH0UkoSTHGbuYKK0l8vIMPXB6gpGu1upKRYxm9lbIGUk1
RaQQB/twRy+F785C3zRCMLt5YP6k5aRePwaotvyuMYM5BzCZyBi70qFc6pkamN4F
jvNqqWcpZ3XUkXU7bNk7l9KhUc1PVK6AjEAimIEqp1WWLpTYS55nJ4NWWteG3ZEf
ABP7nwriRdkGl3k3jnzV+vT/fCak9Z1cOShHcsdMfUYbdcXgoFeppwRV/SC3+Z0n
uXq3WANVQED6aFN/BBZ5lR/5C2qBVXLO8eU58BTyoOU0Q55OrVRx5v6u5H8c6bad
BZsDFKD8r9SjcYMGxsu9RgMcUS5nlxosG+Tc2LC+/tmKTdTwo9Zg+oavnpDaPkR8
ru5KRFuy1UlFlkmjudVGc/whunr3XhWq9dhd7xmeFKp1iGzj1p6x2NDEdmOvWpYd
AEjTRDMdznZo/Nw+wWsXdr+koC6gR4muEI2ZaGIv7Am6am0tyOjPAT7+j+j/gIbg
lV/aAmjrUkRYH9KoiuA/2ybXRC+b4Xef0zpj5sAI03pkA8bT6bBJspwTTvt9Estc
fdXB/1oV24qo4Jsr+TbKFJeAAYon51553NmI44HTXboo3bPZTrOFuJttylG9g+p0
vgQ1Wtaicxqmq2k3Z6zOPowWDGwYDa36E6OVDnV29+odPUvDyD6ZG/pi+Z3YO19e
KkSLggj6FXt6AR9TRhDgxVePVGl9unhP2lqDHLk62PXdmP1MXo6zM94xoSZT9rw2
q0yihAjtVXkfoUieh+9d1r08JNzJi/V2ILsyzU1/cnJQujycnrQeQoQYeq+s0CEI
2YcpeH8zYIqJ8p+3HxgnNEcK2FsF5Eq9A2Kdskb8gR6sB6ykYP6Dz688oOU+tA9g
LuO5EGJZ8YBloleRGKrMPx3D6s9L66vA6Z2rpVaLwd/7DtE+QA/zqRpft1Z3w8Rh
5AGtcbD7WCacDNc2wr9psVZv5VlpdJVVutXjCVxcPiAan/HgMQq0WOTJomT6IV4C
AN4pk0snvHPtiqSwBF4+wETaRDvvv4QA6KoN7l7kPayrt8dkHBd+wnvdu0OL79YT
rQGQEe7EC99TA1gc+RUEc+LxWpdBHV8qyfjbGrDVEIzDxIE28W2/W35DThL0Kqy/
6eZXrZiu4cLM3/0xDSR/oBMq3gh4weSacV9p2b7hpKWMZqefegtkUMQlVEUDb7/6
T44Lb+jVyL7U1hxe4CoxLsqIFKaXBbo/ZHF9a6f0ZmUNKN8BrtqqRHiNfgqWwlvi
vRhAlmJgEcqY5hd8VvVvS8LTSPxlyDS+r/ppljo2C/cTMSQ158Zg5uhpcFv7rk7W
n1SUrsNPQ7zGpLWURJnRIa2uIPyK5jXoqXQWxPRUhN/e6x7M3JGGzMgNCQHUNkG8
r8Hn/VEDj1KC43kHutdjgmv9hUgxXZ1EPaAC1cqTvboFIFuncABiSTWgk6ZYG3KL
m3GiCQccTSXvb2fJW6r9UmNrLm5NYpo/8FIU1kC+0X91orVbR6UnZaERIDCfySYC
zAJVk8ybP8R92gDRFv0jJivCkxrrV05WSsqFMxa8sCEXtv7/zhaPol1/AlzI8Uqu
XglrfzNJ4MR5ac2UOnZFmrCCZ648aTe50NY6HkVwjC+wh6JHzKHU81sxbZmW4/2s
rg7wwJ2S5jPQHkAYVQD6N5evzSxKJJGw+2aB2vHF0ze41koGgfVWycPMyGRH2+yO
VqHJmwnEVbgAajCA6LOH1Ifmw+uSOO8KLWH1YfzRekwTtmbB3WIdrmYVSQP6yuXS
JYuyJFlNZwjTNkWD6NkCsyD5X7DeBJ0GAhxJjdAuyl7pKvvua3sytAo4NLdtw7h8
Bot4gfSjXsY6e55Rc4jo2u/Rbolxa+bENbGFKrRsdQv2cAXH5mYO5gNYxMaHRlST
KmMVQaK+/6keVvXDBaCXFSK79ZQgYbb40fR2rt1GoR/wHJsCculpT/7OmMicXAN2
UTF/HO/RzNVkXGAkS5VnVVgR8DxF5VjQHEq/O2eZHS42m94sm0o2kl9XEqJCNdsV
4i3Uk9NUDcwsy/5VNu63N9ndW3kpGHbf6WXYK4KHUQHM7Gbqm652O/VQAZETgEv3
Wiq0+6W5YkzHf1d46RhAXsHn0aXDgRtEscd/797+EextW5RgjNNVFdlOF8fmXzLu
kdfPp3vAJFYENOLEJXyP86wm7VGeQM0vEq6s9+9VNQ4C9ls8Xv8dzA/9tvw/vjkX
kARGOay6Hzn5OYZklt6omlzl/HihVrBoIxWdscjgOMautucL/eVfnU+bmIBn5ByF
ITBhMGGIgKJRNgfdGp4n6h5V/1TJ0VdGUjhsIxGG8uxmcUcnsTMYugFq8diOv8u6
qegXVLz09N7CuSe0viIM3oo3epd2jcH0zY8xdxZEUcARW9JSx9pg/TB1pq9IMb8e
sCu6tQ0jtay0sXcA+rTf0YSsAS05O+IVDY3EQhEO7xUU5f6MEX6+U3vbmxK/Aej5
H19t46dmKdcLZTphRsvJvQk11O/30F0D18rPC7v/RsQRYAZZ5/9wYCKO8QhMv0Nt
IznNpH8CGsVZLk2SyXTkQ6yKSL42mYKR4RSOVbt12gwYVkXLs0fWlBamaa8p4I5b
6LO/GWGqUQ6DYag26YKLt52Uh+M4U45nT1PMRF+F6Uvukteis/pHZ9Yn2j1SiHvk
LqvwEAj6NuP0Kx4W4eKudO9aNsepmvAPlgwXxuPJWc4Y3+yhvtu5a+/Ljnx8fy6X
3VTkqSEc38vVzPSuop9wjz9q9xJ14yd4xUieuIPjRVjh7fb8Cc86ywdIPTwaNHmC
acN/PoIFFSeTipR7B8o+n9Fz+yv/hOvhIPIwtTdOIv6M+YE4d8VygaeJ47k71tDX
IgXvNxrwze+HZu0rOhzpewchoSLD7AIfbLEIY9l+jimkcmBj0Y6F/nK7yoGoE3H7
lhCVfTHs2ZjjKZ4zCM7fLAx4nmVlm8bgNCkwtnCmAOmQlxDEFykMxogxA4TFKtru
EviV1CXrH2rwN5Rb1kMtHqZyJhSDU2g/X8tBdPbHAPeJ2RIJoGxcBb3teb6uQJAC
+NaUfzUT8a+Cav91BOzVx25EFlPwgFYO6MEcLXmae5FmF7XSZZD4fIJR+ODq3sMa
sWmK6lcjrHj+74V+xpoqHPylfzw2X461r4FTDUE8xdqnpVpYqGzW5nnln2P0WU8Y
kYoyNFhG3ODxXjMDV7Yvj0oA5Veu2KgywWh3jsPjhuuTWepM8yvRq5CAvDNE5fZ5
bOrrpljMCeuqKQ9rsARBwpHbYFBnk0YT0dGHXlYoA+YpSh9pKK2ndYjTz1ggiqXg
C3PXLZj6FNovhKDLAMfwKFYtr8CzEuL775gs7TwQAj47y+bAAEJAlthRCqh4gwzZ
yUs7oMIDH+OUFZrOP3UKUOtkZt3oga+LZ6ocJl/l9MO8IEYrEwEAeqceOTw4b3bA
umCR23m9rqLCfxuhbr4nN3B75KVK9DvnOlMBQoDAcoeweK7v5eDnY6oYRfLR7gKi
XOCVVk8KFP245NaVuq2xpICZh40BwRlIspLKaR9SOIyYXuSpxKnU4ToxoC03IPdg
NBdZnc0qOmt2KsvtY0tt9ZeBa/4tK6vk/xVhh65ptiQIbBqgWe66XEXM1u8BQQM3
pa48bjwMEtF2f+gAIVGGt548ERDmIg70JnVKnL4dmZzRJ8Jq19k3QV+ozpeCO+3b
Vh/FsUtyzep1y45lWLy1bsVKtrYfnsM9qfb/nxAjxSutG5VzORbj1cCg11LH1l0S
CSGE5hQOyLCpuDspwwvJo08K8HVVf0g0imI6v4pUdOdA72rA7viHGiyyxJfApEj4
SY61MSL7BF9Rdn/ZHchoaI+/irdvGbgHHgficcKRDMwXR7BhsgUVhoBW+H1PcVxX
zUXCamTYie2MiuO8loInyKY2/rj+M3+oYsX8GI6C5HcfSVigWyIMZkbuViP6n1GL
ZEMtgzpm7lnGq/f1a/HJ4DUOnlIhJA7R+PfrdiurvWqN0V+RBVzsmNTuctzAVHoe
RTRXzwu0qiUb7R7HVesbq8SRj5p3UWL234LrVnBsY8fjFdBZj4CV0vN6dBQIZXsc
rNNbzOHzvD5JvQyTpwfs3ee0HZONw7EyL5WmUE4WPk5V9zE5bPA+v2SNNmhYcQVR
tN5zy6zAx6+1NCVN7lAYnejb+obraCdmpAFvtPwhzSebpqzP2jfXt9esL8HceVpu
ilu0jIixaaq3mk4C16jU+J63IQ1VbQLIATqLziFaPsVoA7T3v0/AxK93H47rOWm8
VCRRyEB1aZ1OygyqyJy90NaWkQ6oXyUUI6jrjeLQy9NVx7LlMGzaxTHOl+QP6IE/
Kw9T5AKBR4UE4iBxrQbCIPv1N6bSe1cs2TZaqIQ57nMGkpVy812nuzSFT+uqSN51
dWrmnfsIXF0whSLCCXFu6jzSo6T8VOYEztDyDoYZCHCb/gSBpCpbUi2Py19NGhJ5
aYqn8Teu7+UZojD/Ow3qpRf8QmppWNCaXhGsp+q1HgvyAL2B15oFsrU5QBIWzTmc
yZz0DVcjY0/pQg5xF8APbM26oFhBzH1DrSM1UOZ8ZWBAioBPX8cbMJdEve/1Wsqs
1f3tnKAhNAp26lOrChJp+liuLpW/itMa0GvaxOaCjhcT6uJAHyaFCkGAW7aq6GhM
x9uyuyk8bAowpBsqdCbEEpkEXqVhQ67ptTzUEXp0G6XWpYfQDFfmPMbx0KlvU839
qt1EAmTx/+295qcs8btkiard5jQLYJb8VdyycYAIxb7+7ERZCv1plZb9YKN0vF2B
wPuw7QpeMLI5mWmX816r/1cn0ncDDmBBvo46VBE/PTB0a3C1K00XPb48TPu1Cd77
FaIzqs03qhMwO4VprjqfzjXkh46Izu84HZHjcLFjDpk84/LC9yL0LXmfn4riaPvN
qLQWNqJZnLwG3oTgg+H6uq+nhdLt8hgemy2O/jne/Jq2FqUB88YFCiFIXHXZhvpB
irjms7seS1edYbMJDqW1AWG1ebSvDfdgdmXKgjdLe9tWTRVLXdZOlHhHfIrvjs1f
OiMkCWZyeaPBVLhYLTGznwKc4fxW+znoGjJB94Sbk7wloCzykyLcafZt42B898TG
5wpZ7ZfqaGN6sGe3pbHEEkQvfYHiWCW43DC3q7qkg5weE9M4klkTSXgBxJNI1jSr
7duOeC8bcfmt5Dt3bv+kOExrjnZwGkdEuLvm2MVVuXXSh2TRsNKtt8/dPuxIgGav
8UgL82FErwMZEMK98y6iOQxzUkRFQKL4CUs0inppJcvQT36Wxnk1M6mdc3tYHgaS
pL91FjoidyAB0/e6Stau+vhlQzP2Xiyb8phMLzORY4I+EAyZ51fDZPFf4tuIWk9E
4MiGSQQwx/OW6+OUQlwgIPglQO4Bj2Y3XXjjpStz5Xz0uakU/NjAs41Lt3H/xuLn
2vwDGpUtck+IljCTS5UgNOv9ZmcTp2FpcpgK8wtq2mBulL/Dg7/CLvcxucFu0h22
lgI5lzqAKZK1CRpRtZRb4aRsWmygkggRWsgQbUwtKEPzusELSLsGiEKOJZ+UKvOy
XW2Y1/klk+skzdqdZMGsWNqRHR+501vMUAkL+Ozs9OEUek2Rr6wp9JiX+F8MIqlB
lPWLl9h0FFcdagilaY0+HoiLjoSvcVHCMSTFpcgLV0l14MQkkXfyMFOgNjEzK97+
/aZgjC2C5n8L0tpLfJEGzJ0UDcoQwy4Hyi0+Vu/4fGPdkLkh2870bZIYrG16O8Gv
fvBqGwY1ou7TKmHSIHSN/fosKmO4nARvm9SFPifUJ7Ae4W3w3Cz9TaFrFL5JF9lK
Qj4W8UZkRmVu2m6WBg/dkY67ZCqNA4c7pQZlpXn1eQ/qRHwjG/WQDPboRCdvqb9n
iUQtWSNzLW0KBSwZKh2OrqXd9VudID26T7Iip2xf7RjxsprJiedkpzFXZ7Zav3UN
/xC7E/vSE/kpJLjH0NjXDZ9yqd50M8rp1YD1roTFE2HpgwGk3s8kcjv0aseq2P1y
sYesQ64SV9D12kwQsZgouAtgsvWGHBJMsIriZ/+qcLVVx6I9LqTJpmii+vqAjD7O
TcfpVu6JxJl3d1VQSy31ccIVaXkuZbyGxPf1JJO4WaJlz625NCjQAhhFS80eauqF
LDqQX+hH2zRyXgl+hbRvz1xNRCfUF8gvjeRbCQgoqe71R8APxAMBb0Ee1F6ws6EM
0aQfIT48td4xcLrQ++et8O5MWHe1uktuLQ5tG4OeMkdjyxIWITGZSfBJIpamTB5S
6m7a1l+mw2m1eCVAtSJXqCyQKFuD8jfAG6fS/hB98YJV+vc6JRV5jY/O6GPUH6H6
Ojj3Qb7reQW8iki/vTh27jahPRYj11WoDkD5N7aVYcErk9e/VW5qJfPvEHBaj6S3
75u5RVUnc7636blmOKiIVDtnmFx7zoRfekeWsJcCtq714zDOVBD9vLSFVrCfXodL
SKp36B2cUVxu3H2vg0MnIn5Yq0JKONoXsN48jZavOM8TePzr+jXM+GNR2pqHTWjj
4+9ULB/AgBrt79Z5p4LfgngkK8lBWTrMsEH13uHBFkYrpFnBuCONKa9eFmOYz7bn
uqpKuFP011JZ1tNaEiChTnhfQOU3n0I5+QHu4kAxzXG+V7nlMRCLko17ZRbTMBWb
/qkYAZjGIqTpnJ5M53yWQwf9CdODCVKMc38ZAbJHnydNLkhG/h+yAsTBFMzsoXXN
0678xRvUfI1pBW52qMnEm22kWJPtt68I5mpxfO5xO66+bZ+R4O/ivvGWZGzmWtDi
hjJUag39wtPExGGzCpfUX6oLBQ8b6iABjkUgyNgb9vNxqcvVVWc0EwfYflZlO6XS
ea5Ebe3mLGYZGpxvt2p6aN7JrHEdC59DZwljhp+EugQqVdY8Za5dNJkez9p5Q69i
/7hp25KHoe9Kvisp51/4utFMpll1e+t6ktXVBdzAwq8i7PjnSBDGxdNoRW6RSfXq
U9TOeSfSlC4CwIKIOKkWIdCDYhWIrhYS/EdLBOF+noDF5BEmDUKh9yzY6F2FNm/N
HMAzpuVrX+N5CWDCUbByvvdBwXqhwfcug+zzyMsrlngrQCvdKgylU/LuA8c4MmrB
LdWIoZY3+Sn1gzLWpr7fTU3AbrXG6tyI/yglHZLAQzsyyCqjrxA56eFxbkjUEos5
ul30tqKhX6jmstUsX+dBfr6etBKpQM5DYbTRMOzM0rTqufmhofVuO6oVe63g/4Po
+zsmxWAePzVKZmCLS73l43fkq9TCu+6KIv+B/DxlpzpmRu6C93BKnlJDUybIDAiq
NQ8Tja3zsdYBVAlXyAxzc3Al6rVLT1WZeJJrHC75MYMbDg1lL1Dv7GG+o+mXKRhE
4deA72YjsyAwjUAIDmOcVFXnoQ70DPt+TGJKqKpniIqKD2ziLWq+jUJn3G+YRU//
VNUISe+x5p2qrRrZdeVsDAY1wC4MAOIr3eq/sYdPQDJbIhm4NnUVIq+ed+0YTZ1/
XPpczkCkGMcxlrCJZIqLc+VVIV0n+2qasA4ugbvNYShoTai0MTkSnqxEDKcjSlz4
W5KGnb17x7m9gRvjPViq7fbSNsjnRKNTlBD9F7dYU0cTgdeRLrJTWyu16ZKrOfRL
14h1EeJnO3tzTLuihE26a/tt5iGI4aMkyaDobe5EME6tv/rA9F2+HanPdv7InsM9
Fa2zjRUR+fA7xBzssStqvzj+1vUVYL7lnEmlwp6m96Elrd6Cq85FGissvBTzuxK1
ZjQ+/ka7iMW7Fwxt8GnRsFnEpnQvpk3Qx19/Lw1HATYeMFJnL09AlZvOH3RX+lCK
1HWEwe5ZVRD6MubOtFmE3athFEgYh9t+2HoTPha6ssAITSW1cLaSq3kM52olUA5w
PtH9bqTt7IvSqBiD4SkPU/f6e+aT6nBDYHOvp1PUBw192vptOHcI59PGm777W4nr
bvDO6VnHWNtDuwydfQPZBeNUblos5t7mgRr67XtgQuUFBZzsWZ4PmRmCZMO2nZMe
vkBzQSof8Y5T4aMDu8tAhMYyhjb8JmEOJPvbEdMu77SYH2eiIMm/mal9cXm0l5Gv
hvS8vTQQo49M4e71LMaE4Z3JVJi1GuY7zE/dz95FXNFp/WunbR8wzsiveg+HD+V0
TrKByc36CkYYXN5Z2l8oYOXkyhmzmOoIKmzVZuacuivWiu8CSrkN1b/62NvVbXNJ
/YziRd4ft78z6k0Phe5D2s38rbYU5Zh/DRqOOVrhgMkbViOoO6Z8jRio5aNshx2U
r61vMjPb59dgdwWS+j/xkhmQW0ojkZfekJMhPanzjEbiNA01OxRCAtTw7KzpuQfD
+hvaMcTmdy+N+JZtiKP18ttBtTi0Ry/42Co246VtofDGuaKCDqP5u5wtDLzgTDSY
icm/nwjmWF1KJeaVHygVqufXTWa0aBLZRn+Ho1aKzFla5Tp6+NRJMdMbUHwuyAJ3
jgmuGuzE9toZJ4VcHucB6cfj3HkPttlZL+55bWGtkPJAEF7PHWHg8IQcXh2ziPG0
MdeDcEx7KXVeP+1VfNfAUSZrvDW6yV3US0KAGBAryj1vWFCLuMDL2i70Sl1Pn65P
7YJybxV3YsxuLGoLNoGoGTzt2ArHxK4uDDZ33BRKs62R5wDqqhEtSyGz1h906jfw
voYmCM+iuUFYLlgc4f1mHZ6oAuuBowS+eyLcHRLf3AymeUBEhZexoHpm73W1Ohw2
qJQYEm+RqZdTMNu+AuT4dRc+VU780b1gU9Npk3hdsvH4ORjS1F5jLn5xqMuY/G1V
Ei5f3M8owmHS6QdDN9wt9QdQ+noMx5iJ/uz8siMLsniLBr/Wes9Uh6OYFg/rh/4Q
+Mb9g+OuegteJdvYMFc3897JHCGmeLPWc0Wo/QiL13WwPhG8Vxt/h9WWojCWJG2+
L3eoARr51pWtfzDUki5JQZtGxQtFjM+uipTvlrx6yqmlRZUYoZfCGTUAsLEXKhfp
ZOZIqMuGnux5/N/d5EdI+wVk+ZJ1bSEH8BYIVe6jKa6UjAMEPfxmG+1tsVw4wTxv
/HCZGWXO48iPYvX3ZvBlcjwaZrz0gXQt9aGkmBh2X2+RuTwhIde08nAr1EAHRN0d
W7O4IUid++xYGtIOqcpEGsmxqJwCWSxfuFdAR3zaGBFy7dYmKc/NrQLYlQsGWYYG
H+2RXwUvhEL2aloawzh+by6ec/1FqLusRDCK2AM9jdLBY3NBXzzljGmPJcSMRcS2
qk1IZ8oq/WR1LgXulNS3Bld/B2A1LpduPgn7iGPSzHxWLposyCTwTkvfV8dqH+Zg
P8FBtnfzHkSeCN6TDVc0X9LA8sifjqBaEPrHxjS7aj9Q5I+RTtR+OCDsjvHaY9Ay
tIMu5c3Gjwpu8uSLHwLAWT+/tOzV3iZlD7fS4TURTrHSG09+SmaLnazFJ6XH+qD7
b2lfDrpeWQMXneX9ovLCOXhzjAybIl7sfnU/mEYWc/2Sk71kcCxUETmVO/AeFKO6
8t6Zd/UPSYzik+E7jygSsmzEZZtdBL4hQvSIXt5BYzCCSWZrACz0noAG9UZRy2wL
0a8LRgeMHbEQPOa1twfkqH+OMDO+/1gd34lR8dq7/AA3MGbnd2RGPMsRpNaC8r8l
N1lL+MuKtDYOvTZUjCg+3jXzg6aCnh/EFXUWwQ9c10Fl7meczS2385KhkhhVIx0y
Eq8UebV4Qf19kjBcu1palZNSaoFZs3FlHOYUK6Q/k/LY/DlJCJJYduGSltC7WzFt
Wlm+FCCuE/sH0pGscwquJrIIdetotgUkFOZXYrCJBJpa5BSBImuqIJ8R4oX1yo3C
QL4O4E2BxnjJPwJvapTB6HsG9yYRYUIqMDEaIROIIWMQefYfGxqTCz8sMEGohJF1
hNp5E5/CKu2OJaJMoho5gWHGqoyQ4HS4nUycqEX+TcfeooxfP6dgZ3miZWIPvY9S
eiFthGwwW3CLmgJpGEKIg9TatgVtUAzG3AOy/hxGJ19L6M/D+RWx14Vd6HZmnSJF
ty/XNJZ+aiGZ7U/T/0Tu4wXeEfrk7SWg4L5PEeVms93gwc/SDWtXKbZIr8houvyo
y1awUjwMFTif2oOJkL4ocwsKdcp1P0vTGb+fKZ81Sz+oqYyWx0ev/ka80zvonSyj
6duYQUm1pm9D0NCXTxKhLrl7FpOsdxcfb2xnvdHOHJmkJPOTj2EG9pC8zlTTLGt6
laABmPXYfzL7oOY+ibAKH94uOAFK6wiWYby6V7sp59BlVI/LaOcoO/h6z31edee8
kuEt89v5GseUGOjoLVAxKkmPz6n8w46HRx+janBljHFS9fWPxv8Vw9gmobaeyFjk
v6snztac6tae81R9EC1a6MlsfzFT53NwSZx9tTIWS7uQz7C9kze7YJlE3hVEE221
XvxaACrA0PpL083/hkaXYQphHjnn6VjJCQiMZ27AU4Vnj3z5bH5Ozf0aUO+u32qk
Fj7CFbMcPliDiA3iWTJfZLSinklLefZFmQVBszEOsalsG/o8/vX2i75uztMqIgdq
1rGkr8kyJBNvhMuQOJKQR9R0B9da/AlECSwYzYbOR5WyjJ73qkxZlu4ojdI2TvY6
HDtS7TIFkGNikRJsDwKTBo7BIqSunmGobuE8LW9+cwn5WYX8SC5xnhUZDYfmwcfA
vRJCmKW8AC+3RMWdH8TU/ti4nIIdztQzUTpYidPm5Qxkzd+oqW6i9MEgOgYcigk+
ZoTY9ZZ3nNS8MqQ/Qlt62bs7O6ViH3x7fxzrq+SiwV6z1e2DL0Dp9/rty7HNz870
QxrKIT3JUTikcQFjpN1Z9oRI3C1m6OPPra7wNBHUtPSuCj10NAP1qSqfoUl3rZM0
SpmyeBAzRnai/0b9I3MO6dPjRkjkWPq37xye02JfpMyrP1wRL14hXWFXRw2bfhrf
QYnYs9xoXeJuP+idyUr1nDZ6NNcPBxdWr7DNbCsxkTirDQpRKDEozseTCr7jrVIi
0iUv7tg/qZqxBEKP1iMR+BYwSBUJtwrxHsuzwIrteFA7xG7oU6DZFBMJ1lAOKHj7
hx4pn66F71LJoqFoR8tdi6ZW1yxyG/JBr1SCJh1WvvU9UV1SDzSQbR1VJQiypdo7
YrD8nBOta977+5VAMnSzqrYhscd6m5ze8l7HDpATfgTyZ8YzcaMSftADvb9Vmm2F
MfLlGk0T+UnvM66nwg+s5G8nPNmJGVzRwsPJj4bNsIQ=
`protect END_PROTECTED
