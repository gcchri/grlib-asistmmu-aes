`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8E4ypiOIgVaAsK/5+qy3F6DgF37JTtHmZN/nIDkQMQZ+kGxrip6O+o0rVaSJp3F
Ml0TQCccuPsg/1F/W58sf6kNrnsdqkIy9IU+5dkvJMU0otlevighlIvCPbU9IX4x
wFZ82XVF7dFjHNR4t8LINHPBtPXZPM9nVF+50C+yGYA=
`protect END_PROTECTED
