`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d+8g5NBgdw2Kg/pv2WoLfGkoMmSVLKrVTbiTLJFXDFY6LGvsBXjhWB8hWu+EhzPm
U2JaKXH9M7RFU+kad++UhCG2s2/eiwJaIz7t8TBv6drdk3FHD4/cGBKa99vm1LAm
EbzjgOGvOipLTxcBC3qSrjoN/zvKRIBqer3LkxMTTDdT8Mv5vYLONlPxp+KSDZWE
S9SMI3WsDROJhk4Fc/E9CALi/IlUvc24KFHtJeN4kMLx5VnGDKVkJkScJNa7I7/x
VkNhdo9uNGG/E41MQg3PDDaUMUc7q5bf8ghKpyZT4AsEaOJfL7+Sv4FGUW6tG4Ol
izTtHAgg2v0dmDWtBuWKYEqiRHPmzlluQKW71B7J6KTOFDxwO+Uk+Zo7BFO1z4aN
6cH1zwLHHRV6h9vYkQ9Nt4PXrkw30S2fhCMud7iGxcyxkt/zFZP+VdBqB19XHiPe
c/Pwzs/rAMNEBFINt7h1Aei23DJ3aZnJoVfugKlrZGavRCNprWg+r84HFQHngJnh
V4fP2K6iqdgEbtRDxrgKdRImLFaKGVwvjbaK4K2EwnGZRS81TkWi7Z/bWYVSmsud
p8u9rM7mzCIifGp0KQkiZ02b8A6xcBPcZCNsRgiWfxEcea32BB9ZiHjfN5APl8/5
9HNe40iPW3S9qCuN6+3ZBj1/F4u84piRelZpro7jrv9Jgyt9gVjz4A1g8iF48JWK
Q+glN4L8uZSTLsCioRDXGA==
`protect END_PROTECTED
