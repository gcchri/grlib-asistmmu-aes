`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n9QpytZywspshpDBTErpO9Cz9EZ0Sb5qzwpZv7i98zJW79gsysCt737JVZ1ia6zw
pg+rGPlVN9pb5ERkU8KptuiE0ff8yDBr5MbOCdFn/EkDl06a1A6PD6nYlbRY/yJK
ujKksTAyUauYM63NAlJc/UV82DITymbWGSkHjcPeB6W39BILGQQqMSPzJz9VXzH6
oGW4tTQz6KoxS9A0HakujdGXUI5nhC+TIlKq0uSyHsODs1dKkNEVRVu+SRG6OWec
O5C0ChA0jnrk+TNi0O+X1Fsa5GMlrby9xdVei7/1OukmhL92NZa0rppyE0RfgbKQ
OIn4yHEB3vRuP39N1P8ZFQB0Xj5DcsGbwfmhJl5Hpcb0U1zwYzzTmy6r0hre/MTo
4dwrdee5JPXSkiPELckdNGRmw46KFbbHhRhbcVydOHgD62HWoscVU5DzMGfRjHOU
KhPBlZs7t6uHw5J6/GgPlXiv1y+RslVESJ29A/t/R7XVfocRtyLrpUq2SycnOBuc
oa255NzFJMkjedKH+/2fxIn0zQHNG65qq00Wgu9iizPUusMxdShF64AHZ+IEUaBn
pnl5MkS9N9SUxJUGA0bC/2gMLhk0zi1HKwg5SnihrwfO+kXWciacg+zFq2oxmRwa
Cn3Xp9tLNY0iOtcQKJfGdfu1NJUNqjK87FP55VqFv7h9gbdmwIN7dKQGg9itbiEn
F2r6eg4Ztqn4xtj2ojAl0by5s6J9nhYRgPJon80yQrY=
`protect END_PROTECTED
