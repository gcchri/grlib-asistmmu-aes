`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/721qNdfxZOekETGAnnJ1Vd+imssaPU2Hwb86xemHeNY8b8A58/e2P2EYtxQ+UtX
SiKz6Uq0aUrbzgelM/pt+PXlYBmqdP+iMYXsMPuO3VXaFQy3Tjs9GqFgyvWqqUOc
h6PRjsDbmNSC8O1HpRuH3ElClGsP/kf1V0OqD+0VsK/LSgKbxfKxR60kNt4h7moc
5grfqFXguib7mw8crQgVLzpNdrLlQlRoKegLMZ3m3jOa7WRB0WEpzHUiFaTPFbd+
SWrG1UDqCvyShFhN3H55Uo9IvfU1aEvRgGTloCd8xSnMRj5PQNVmBKbaDhV14VOK
2k5LzDeM9kYlxLMonxffpfvwpLu9WnTVvJF3N4ZAHXYLmJY94aTTiyQi0OU/M0tY
g0aGxDeNe1+vBNdSd3mPqdHDL2nOyJ59Hzot/9enCo5RBji8pya7HwYSFtS8kFtW
GE6GtSWMx/1DBS7wzCYk0Q==
`protect END_PROTECTED
