`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OERZi0O1e0R2y2avWN/mNjdW9NtYlp8EpOXXjOH9tdS5Gcj2ClVY+QjfXtZ07qt1
xmMSoK38ScxjqXG3uVlAMKJW6mmz50kJSRdx8LxYHm9SNTD14hzmFPWpKuNF7I6L
yXA0nCLQcDMP60GsWP2g3P4s8/WlGZteSC/Blcc2xav06quGk3Kp6QlpdfE86hYE
sfSomDc4DEQdpprXXCbPIHyW9EIO7hLF+BN73WhO6x4qmZk5Fz5zZAwjCulSy6av
4GXxvkuJJEBbnco6KM6hJb4s+raO48btBUKUVPN5L8qAb5vxLJ4WdUpgsslWRqdH
rRRGp3iUZfuJwqQUoCeI0LFbMypGWf8ZCxbO+eS+ANsWKPLnYivoGzaJ505dPmHw
HjDegbiyH+SSSH5MpzKeqCHOecyqRp19IXnU5R4PPYSw+q/LttYLUrtt8+vdzDmC
/etq8kYlY04whF4zUXPqkEbWFL/zFMBej86/XgrfOlH+nDu/GJ/bKyqohJSormqc
IBXK8FkhlJ5uSe+hZWhYjoFNj+MoqLPLdZWd4Tz3rdP6hg14w27iFOEvzp1l7S/2
7ju2Z1fjFf/WLF+qPdFb7nOOnrleHzWyXMfEAgmVBC/yNBgg4pQDqMW/9pMJybg6
OGuQEHqootinlCuBmrF/TwKWPhp5gXp527K5RISHvQz6rlBLorEB5VoUKp8ssgQ0
h5Hf8wMSLal02bFP0ZOqK5eYOuM9O9jeaySJeZ4Z9/amEF6iUXTZiIA/aCTq6rxf
mnlrOBpdwcXecWQJgVGgZzg6xrjwsYy+Acp7cZSlSgK6VIa3I9yoYmpXmY9BTjSy
SQxWBy7WQhhwxXwCngTedZdwMQ6uduIYXjgboP0mGNNLkKtQdMo9nz4/bEX1Gg4a
FHt65hqHAx3wD6KMd8OlJRWu/HgD7EuUly2OY6GolVLnh4aCyXhsOPqdQq4J+IAT
vG4G4fLT6zfBMVYmtvYqst5xXr1pGjgbxKwDwqEGv1CKPZxg8NoGZPbLvbii7EvY
EOyp6EAm/lqBcgAkHDadMZ3nvDRPyWvedqYVvD/AASwPP00sgFUshJn5bpQdv/KD
YKDu8PMFtiPJFm1inxYMWFjM2yJnHsUG2p+Zjooe0XaH1YtalRFw5xPZ6aO2yUbO
VqxsmXTkIkiuGUVr7lH6Sg==
`protect END_PROTECTED
