`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGet8WAoox43dReL9T21207HDMcnw8u4h30RU0F3JYd/N7f6UgtLugr9f8qLJ9JN
u8LumdxwH+5WkB4vQySpwQ+DIIN0G8GjgrpWmHfT2fC/NOrbWPvs9Nx3E4EkoAdf
/h8YJK7DP5LNgmMTXdOvNAtj6RWz5vbD3M3arj8cPca1erNvhNrYKHKxI/txkqwN
bNmiuTHlUXx0BLxPBIzOZH93nPTyobyWOG8HyGkBSAEKieCf0ooc4LuSyb81EiJx
vSo8F8+5kojoFVLDS7fZljmAh8yyUoiVxlio2shA7T4r8ac3PGvnNrmW8Y+dx6Z1
B7Y1MYhnVSzdr5pGRVHvVCiZwaZX464fDHSbnFip8JWdQAal2aZ2xhB8ClIx/tR/
zFAnCjtArS1wlbhHyZ0J83ifO9Em4YJfDhYf9J4tX9UCZ+8PzrQNvfngtsmQjdqP
alGQRGpwS0q32xvKvRJHfoOiw2+b9RAdeiAYEzcmT51rfBSuuzcbyKvdhXGydngW
FBrVbLDA39qc/KdtvKCK3KcS2kOCtgC4TpsvjjiBzVTBhO1qrEX7Il27lSlpAQHE
IHZv+WuSU7280uvwgouYZHUHiMz6PMoCmyNbZHod9x0QxBMZwFHd5caTj9sf1qyW
ZSYcT70PEXuqBUD9te/EzaxvBl8k7TwpAc4nO7WXItn9CskRlRCSlDx7eiBWqtG2
UZ+NPkEnAcqDeKIeo65TcmyGhxo/67cNrntNQLgQU0zC85qvyZl3RQ8H6YR216az
g04vtCPUCZINdnRM1LY/Lyp/eTcnU5jjSP1B4sGupyd/H/zdpF4po5TJ5TSHgsgx
N4MzQBXoJih7sn2HGYYa+qZmZtWhLSaVQWvZmK8FvGlIJIaUmLTPHy4VTzH3MNdH
ix9sLBLH5Tp7v/NIZbZwYb68siqkAPfSOWDlvei+/jwkJ8gTTaBF1zrc19bDRypV
ufir8y9xZCB+7IArrAABGrRVT1eLOWTUtQF9f6fkqFebfrhn6KjGzxAH8RwD5QSm
HpYLLM8hV2AXMLyHpMDucNucWjqsx+omI5gEx3xIuAxPy5YRou7aVEqan3E7QB/Q
htMjbYvcDIhPbAQweZ8RJfu+DtAZgztN1wAEjpIl/anurFsQ0+YcUCY3MRRyT3og
IWMBTehhgprcsGItWpVq5xoMjXmA1G5pPXOhpfO/andxiyW0LqmLUAjM0wfVKjI2
/aXU2fHKjFfhJeaK1MEH+DRfhPj6/jVYhM5tp1x1F0fLxPU8HWyDP5MbE0jmjG9n
Sy/nWMLxuPXfYnhxRUpQamOojqFukwrnLOqyZtkcbdvJcl6qtO9ygWgAtQfaUxNa
g31qPOcroOvV4789jtPaSPqSImGmUrCyK0a4t/OUEAy2qJ3NCce4p7FBXI0x0mR2
gcZG4NmoVFoVCruUt0qpLrl45jMlMqIjNNFyQiiAWMk9/bZ7nO+Or730AVYjF2u/
0e9l5/TyvpcIlV4ObhNSO684OJJC7LqdqMwaj6New/ugfDCXfPGu5NXNfxdLOV+6
KckmViCEBqehmh91Sq5mOqlbxhDbmaeJmp5l9du6SzWYEcYKszTogBCC70miISmu
AUwCBkdn6zd6FCsXgokhSlNGiPwKfbTPMD+JRqohemKyvOJZH/MQWalXiY+/pg+M
gqwml7eeHrqhPnku6g/3ltIGrm5w6BQMDlMFNi3q0hBaax7ki7I3aJ4IizcjvqP8
oqA8vk/Fr3PED0Y5sj7Fttu+sW61azlY9/DmJbWxVJJ1W3u6TJ4WY5UVUY5ASri0
9vIqB0a51PxqCrLvpUKiU2uqIuzPCOKuz9yem8L45UtExVh0DxcWELBu3C224o0L
I3boTBGFH1hxoiqDtOC/jF5+lQOYak3oqCdjLoj0n8nhPdVARABFPOACbqshsdsx
jbr9JnBP+hA+gPa8WCCFcayuEa28y7yl0dBu9CdhcwTRLWSGhlHz1GrbZ9NkI//6
0C3501n+xhjEiSbE4t5WfL3+mn8oygmhwwUzIwYsFYISnEgOcChOl+UMMvzk5gwQ
SU2coBtDzB65pQ/ljtjrvh1jtlUG46RlQC8/q04dkNFkbl5VR6mag75FC/NBYCpl
LPNg1TJseooencsdBR8uRTrE9PZk2Gr5KZYA2wKWum1wyPeZmn4ykQOg/4GIz9BJ
D1GJd7JPMXQk9njO9IGRiW6nQ5hyoe9EZKM9axUobHDOd6Met+WTSjkdlSQmrFy4
44GatAWB5aQ1DbUM2wsja7D16QtR5W5K3PhvSeRVGLy5RTUlVw2ZdJoOpkXenMIP
Cu6Xiw1kICXM0+WI2mRhyDsYGXbmtlySuIOVpqKxu8RZAZ27063GuJtS/TFHPO9D
PU5336z+3K2qOs4/zqh06BIRlRNdnq6zDtDA7n1mWEHT9yosNnVaYTU3FtjdMJk2
Rww9qefnqHX4AL+enpVmTS4K4fvi+BxGKT2hY8D4XP2ghs8BbFeN04XgAY932ME0
q9Sv7T67L3I7eIW1944lMP2Rm8cGYhIn+z2tE4+rzmc=
`protect END_PROTECTED
