`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZSk8x6Uw838DeSBpzc/nMHdyQut2x/kF7bEJr1KRsXy9G/6z5TD+psnxvxLdBk3
VlipOzBYFdBZQDg4QU/5xVCGI6rdSCYT3Fpwk3P3Lf+GSFn3jy/ZRxV2iAK45XMZ
Fk/o0hOeBrZLGkSoQIiC0EOL69e5s348hiJkWeqrJuEMJn55prfHisXESMyUFPsT
BQpOaJRyA4qwz9vIYUlwvBJJSePXYOhVXkjCgGbLVGNGUWy1F9GNIuPBgVxj+FyQ
2s9ANOdIuEQEg8hoDUqtWg==
`protect END_PROTECTED
