`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
woMglsyZUEWw7yOQZrFMTu41MR8mJW6VLoiumR+e+GYJ+3tTjYs1KHpv1TycXSrD
SwWm+hzQ3ph36ZxTd01EWz0BMeD8jsm+0CRsoFQWP4KsS34uUi1uJdnbgdFeqbOg
uYdRKAp68ZE3ZEKMNU2vpYwjHyOpm9WMyL1xLe7sJtLLgSZBtGxS71b8xE9N95xM
BFbv5zgoG8cP9W4ZfQsx+vu2wWmUzl/CX9hdPKVhUV6InpAyJW3j3bsld71agvI/
A0hPcs2b42z/9/iB/qtGgPZ8NVExPfJnHy8lo0XelKmtCrdBXzMjZZb8nCY5Ojnk
aTm57nqDvTgkw5mYdetHrouopvtXNbZF7WCZNiGkxqpfE+hKoVgBlubrCFXu5SXO
r83OdeHSNL4PYaAN9fdkFZiFjed78nLmU7ZmMlV3pb9va+xt0hGo3mD9yKUiq7ly
kj5ZjPAS+ic0yxQSntNxawFC7hw5wlt9x3VlhqnSR5Ypt8MUZSI9na1b80fKinsa
ISVgUH5r4dmtdxzz8xSOBmFKV573SQdtxIJ30JsFFGu2Fqn+VdcprzktHhO0XcXJ
`protect END_PROTECTED
