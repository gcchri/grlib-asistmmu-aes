`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tklOcTMCQOIwyA5rljndaGNKiaWn86qBEbjKRo4FeLj/Y+UdeRCoumKpx2sNexNT
n5osa9bZTqlsvfqqNR8Z9hXm+5REj+cFehECHYbsC/HYVhMxQ0wx3NIwdhT6kgax
vHnnRNVLv25KSl+FPyxrVyJHE1YUwEHLvRA24V1uPheNSQPkqDbZ1Gci09gI3dUW
BdK5yN+Py/IuGtmkOeaA2kWOAqLZP+Cveg8abVPf5sri8w2q7KRdlmC+Y+Znd9N0
AkaUTZEAULVWLvxIjAuGjvdDRxw8fRJ8h868zHA+q2BdR/JFpYms1v2AOU4N0ZDv
VV2hfipW9ErQdRFJVcEo+os+y/wtYtRphTCB7V5oKFxFE9qDzBGXiJgCP22qvx+Z
HeSxyfTXNWAA/q2ekbEAFGeBPb9ABX6N7uAxr6r4/6g=
`protect END_PROTECTED
