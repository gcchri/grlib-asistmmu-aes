`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5Oi20djMyKaG2pbapXHir9gl7Zuq2M3O0VA7G8h207sxaGEx2mRmewLm9ZNy3z9
SWKQYG6senEnG747GbhTGyJGDx5pMmlFVmTYCDtGUgK20yxNtFW7ryZOkkPjc2jX
NYCEnvGbW2lrauR6+yIdCzjbyNSR5z8+35JCpqcCzR4S0G8Wnbv4ixOxIDAjhMPp
DvZ1+hGcH8b1l4JsxEvOrqSBh6NDyxgLSbGCaTojkCkftbpGCQyD2Cz5BIbs1es5
qrY5V7Y/+79tBIJ5MzmS4WIntrneKgWNC4BPD0hSqeeeLrUwjc74a9sUyqDPQd6x
AlsM90VHZMz9uoKjBvt22c61mvhfgJTo567RAhZ3YGs2dAmeXpl0CnNlXFyjEWa+
nQCjOx1bEtn3iUXm/u937aig6JJU53AiWZkZ5+JX+D2Uw37gnQj0hWUXNbhij7Wb
l6cbiZfLX4TsvA+J0ssfrDzx6Q6QYLjx19rQ2lesydeJOu5xLe76/eeuhQZbLwdJ
yoHTGDeuuk6ZE/OxCA37URSWCglMALrToXep0Lv6mNf/ZQ6PXXnXBbcas4k4jfx/
Y154R8l2rhr4BiOugvIZJ7AgApURpvs2SvW8Bo7JDzqWMsXz+fl5Y1SteC2SPVAY
u80oHOQ4V0WagHDJmAry8FuuYQ9z9kpoifr8e+FwG0gTxx2mvCfpYETqYqzgvvTI
fWxpJXYIxNM5iYU8bg/8BajfFUD8EBMmyuu4xF3H7jAqfTzjEjT6m6ixBHyCS3rh
8+QB4sGUY5w9sJ64iucCPA==
`protect END_PROTECTED
