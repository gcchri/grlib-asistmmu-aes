`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YreKea+rCIT2+WX3ZYvvUfoIldrM0kmFHccFPTL0WHYtZcE0/SK57saN01+fTBYv
Ur/svQ8QmR+w0CVmsSReH1KCAtovjjbEiyMS7aZh1Js4DLTz/mNzm35wB8dJ+k1m
dM2FgU7XRKRbG1kGAkasHHkeMuTyQogKA4QLyS4pDub7N+KBo+bUkzEKt2zGwP3Q
JoOynN13k72kz8tAWoskKzUTF0TV3Jw/FKPy4e1nuqUJCow1uC8E8ckO7zp4j6Mt
y+yo5NuIjpMIEEXdA0BaZf9PPbQJea4Sx5nCMTJMeZId79k9ZderdaBEwWC6RiZ4
mtq/Jmx4tIy3k9gx08MNT1dKq257+0Hndw3sz8ACtGmsHhvbnKC35fFI74vImhNb
MHe0rTxIR97Y1HT5uF0GpkOckpLA4y+DIx2lKB53EdiHFg/pO/ic+AgURPnebH/l
hrt37MIu/aQiSFS1YmphGL1JlEv7l8RWHQMhxpzcBJzCrB0kjuXnk6JgMJsisrOl
`protect END_PROTECTED
