`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BCBaccNvfnFOjbjFjjAwso8hc01eXwYleGfQNT5vjcBfxgxuUZGeTxVG3d9lKHZ9
diy/x+j6SgooHJwqMk0oFRScyVh8yV0HxLXL9+8ff7ss2uFPuO9VzAofI3WdB6vL
dhVLLLWfWGK9stwtK6THA8guEAuP8KpKRtAbHSv+zXf5IAv3dHZ6urM/c/1TEC8/
MWa/5ZE3Rg/oMGXfRezU22DSoZVNI/CaBc2PrVmCWHPDdZgv7j6L9OheiT6H+OCS
2dw8SVOwPHvSH7B6Ea3Mgg/25KhBnXxcnEjhsznqB05byCoNlfNOV0SvEvbryWbc
AKBk/Iu8ZxlwwetStUZkeg==
`protect END_PROTECTED
