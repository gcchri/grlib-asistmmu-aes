`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZqcBH7OHPs4itZ/vNAv/Jc4ZvVepOm7yww4P154nO80mE2JO20wuh5WM9hbTDLR
T0y4G3lkh6AcfreiH7rGjqI6bodIWXnwZMZ/aa+qEJsPFWzqucmJ0HFMbATSQNyk
vMSfMcy5jJEXvHs4Si3rXWemhxnC1gKuLVarO34UuS9Re7pTzHJUrDMY9SfRE3tC
vETXk69aWGFkOrgn2UMJDIi/aJgvM2ozYqD+ZhBusKyDBtz7QlRnEOGfiyV0PhbU
b8yd0CFU0p7WxzfH65af1LCo52r2TpLlZKlq1iodSMM+i5GiQiiS3ZwAb4AYvNLd
q42nhf1curneV+Si3UolBN74nOAFRS0H8N/S/ohWcNZJHgNlKNXXF3/7ZK6R5Wn3
GFS7NqUGp0JKjNpqXzkdz3RQ5Dvu1Ej/rDj5eOZ8ZyzMWTm6u7sHhQudrR/rAaya
ZcA3EvOfGP1uKAI3XZzMCYpHkilHMaE88U+D/wBg+cU=
`protect END_PROTECTED
