`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+r5YjblrjRLTnn7xdO/wxJNmQs9FiE5ELQF+Gr9xjrxLReBWdRtJuxucKt7cymV
vHAPDKMAUhdf9NjPe5jQ5NrIDNMHyJrIWtEnFM8T4bGbbtwCdMa35G3IBb2XTMQB
XJZZ2Q1LsYLpsN2pS86bbO01lNknAX0d98TpTtekx2k+QWZAGgrfk40PakQIXob2
oY7TA0GnuFCri7o+wWXXiGW0M9Hht6BojXvpyjEG92MSDKUOiVCKh1wss28QcGVr
L1kGpvtSIpWZPF8h9s1RDJp9tYpbW9zyOOL7wuIDCKIGj5xG5qzUWRxfiozvTIjE
D2DWhvaW3SlYfNTivaSDm3Y+m57HTKECeqWIqjuZBXzdXQ/5sXbAqAYZsVUz+T+8
0kxehNy7cq4U5f6nKaYmmdCrsnrspsx04yA3PVk+00vyMYThFkNTsVj2ZgfW0otO
FNPabXkpbEDffdKH1qLtMInT//nQeqahspvHrqAW4hpAOkMtpSRq4vR8m9HI56jM
HF138MguczSLjsLeuc+vO28qyI1cZVtP8nFGBLMHT1lPbwKFmzigsOyRJ3mS6toL
jofe/wUeT2UzAqCjURrklK5dh2Xf2kGOLJYdD5mEqjyyFUGUhgChAxGjmv0JRtWH
GeLmEMkR5XWqJYuD35NO2pv72HTebb3GG01Oqv8JDCCGmQAKS1NEzV2/5iFX/T6N
INX9S5nH6CSG3wffyZnB7yVBRSpx0hCxZNweTy0yjUsnM0tESv2y5izajj8837jf
`protect END_PROTECTED
