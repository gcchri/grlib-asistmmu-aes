`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KCxgXO3ADiJR5tt2Y7tTSqW21WTHE3K2MDXFdlRCiCUGYhvEnaLh8W9X84ejX04H
Arjh28RRtTgD8htApI8iLurixkfMvJvyt1CzzzA8ju8/fzBOhvQaLsiB0mgNyMpu
dPUshGuR7thr2apqS0KGZ6/jBR7lHbh0OKVR1XTepy7QFQE1CsO8Br2VSeLN63ie
xe+vufmyBrgD6Ngi7SEWVffUzAS5ztXM4axAHJYP5xtJSOY+roKWOc/EVjsyD6IS
2GjubJTCNMlhrcSuV2IaQ/6atmnyM8M+O4AXjn8tSV0YQNo9f6qWP8FphhO7Gzds
DYxA4KvwR1h64OeZAurhtMoMG4oTDjXUhi4wGRLwBUl7xL54qsHrw+VnexN51HJw
OK5sWS7otihZ/hdm22KeErWZrfU0ehLAT+qiFS8j8JBvrhHigt7iDF0PjzPsTrF8
`protect END_PROTECTED
