`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xGNjJ14X//TBocRV1BOLrrSGE27txFNpb2JAIJb/jXDpokr19IUB2pJS2VrC0dCD
xY9Y8mem90TsNz/eW7ng+tlN9kLB+G4ZjqKm+N8EJOB2b+1V6feHfTzLiWWn3NXv
Fi7asvPZahO2mYPB42OQG36Oz+XtaYr0PjH7iSUyqAkFMKWzxfnNx3IQyoAeHHbB
GI5es5nRIv1JWj9s0h0itSo2WgHWt8grIrUhQXRNxtWCyUlpuIuAiZJPAzAmXYv4
haAovDdurNSjvbMEuMZhwWUHMEE+yqXddhq5dgrLz2hbwkWNGq6ieCirFkWvjFNB
`protect END_PROTECTED
