`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LuSK0L2S9m0KIPFY7qWrW6ATkEuGHxk86fMPTfKtxLQ6aGOm26N/u7vOcW1vyfmK
5h4zms8nmFum2ON5ul5gKsKwRa1ZXnuowxpeYyPimH1f1pWA+FsYZYpMvB+GWlua
hc0otDeyTphCC3M4nPnSX6C3sb6ATy5Tz8XPyrPuE8UjdBZi74a1S06WDvF67RpI
pUrse2t8Wz67gzTOgJHAXA9fl1KelB6SBDShTdO3T/XtcfjiU/C1dsTR1uPe3oba
4cAbdz9uEdaklksorFr2//aCnpEawWHtLeWx+T2+y8VfwrK2Wk/9UCcxyI2LYLdP
s049QoNxWUe08LmuoZiEdA==
`protect END_PROTECTED
