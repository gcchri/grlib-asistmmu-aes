`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sciigKz9jQSjKaka7ZnEinkLU44iFMBGpAs42EJtoGE3v8vDnl8cP09uBhgssd6l
bkFvLgXhBtg9jWnMZS6f8Bbp9kgDrDd9ENy1tDia8DOhUOsEiecnyC8fg/Yi2tdr
KkgH0J6m4W5H1uIC21TOWtShA11f0iD/Q6H8e/ovby0tFk9rmgrUwmzyUqWadLSr
N+gOSYyiOxnsEbNTslK+KJ2H69PLmUAmuGcPu9GXv1rOK14cK2AF+hG5/phZQdgl
uAI/zcCcAHenL8/I3eJ8EikEnr/PqszTNffFAf7xzP+h2m2sNyuQ+kCDAwN5mdkd
cl6y4nboiokG4ZcqEdnu/bnUxG885X3YeXdZ6n79IrmrsIBaJEVuDc28H2Lw55Ai
EeJAg0+2mI4kGPfXBqZolx7fHQ5iOAU1GZTqv/TtRWYprpW+PsbuNWF/Mz7GjSGm
01F/mfyW6QbkEK3PbjhyPbpQx5BdGnwUFp2NthDNx/kSWcTc4Bk7+TfeounqMVdy
IV/shqVmybTW7ZopJQ+pkYWsEjLk+xdM/EjS6rF1MGKdWtG1v+ObGWtbTVRxSrz7
IvuJIRwOc17eSXmk3I24ndgf08wtTlPgcy+NzPmZBPC6UnTprg4AQB8u2i3YJ5kC
R5IQOd3oedQuMmaUAycdwA==
`protect END_PROTECTED
