`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iPeBBK99ZKdAfftAHLit2HY4YqzIYFjgyRe4Y2PAssYAerP3lqtSAXHKsNf3hpzX
woLh50s8y6cs4EKTBPBuTjYw+s1vCIYIuEOvP1HA27S6pcxUPDtzfCRqxAp6eAXG
NDh4UhUfEDNzeBJd9Bdfs6rQvKuG1I3Ff4TFTULJ4Ihupn2LOCEq46jcn0EX3ukT
/pFJ2k4meV48v5+glM2KNxzdCMMfRSHvkk3HX9KQFwzK/VRHiDy9/ACk2Q42AZD6
IlGwULv6gTg0DLAv+1VFx8l9LEsqYm4DJtqgf680chQNfo01rsHrw1MfbVnDXamc
IA+kG73svRHbmYYsNJQ1bQ==
`protect END_PROTECTED
