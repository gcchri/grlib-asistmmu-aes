`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BfSesJQrYbsTYRin/xser2zPUfJ/05QYnH2Zg9BbA8sL1xJ37JaE8lIDzglBnuCo
/eIvRIWq1CVRF13RrzYzz4O86tfJiuZNxPpNsNmau2ZBcQgHBwpWpisssSURIf+7
UU9jfLxnrIhbPam/GxYNcSK8t81E1iqcWYmDXiNX5nDj4t2CoS5AR8VB/twwuqsq
cprNMQ1+W0z5jd64wMsk/fQqJkClEw2LZyKOYTzJmW5L+wJFmil1AFwLHAssyyZJ
mGwGkjCBOvHd6BraJBBdWKNyd6geKcwrB1Cl+CCFHKh9p/cWj4+2CM1hAU7W1dyt
E1UgSRFjBRvS802Mh1TUiZIWQLlclyVqIwvvia7f93vrSlUVeZRD1X1aWMgvPrrE
kRUsc+dpSY2wkDJH/TXOwB5BWQ560FEKfRX1z1YBhSyE32z7C7rBgz0I+De9v4jY
ATf+N3OhKi0y8i5jmOwREryudGkcptsl2AxWA1SKSrt/YeynJPnEAfzcohir81Pt
foc95kK4zAGhZZU9i0uSbYei9+OotyCJGOiPVbeydIO9VQbpOiqhzTM/cM+Mfz9B
IsqQRbDmALRB/Gh3Usb+Cx74y71HyX8lXyaxHjcX6nuwQDU7EGEbeHdxvO/y1RlE
nZGbUtr7z/PRYZg6DOIH0/rVwdcaPWc7+znQf1La7AfTCp7dx8I/1cpUOgToscjS
VAnvys/fb5S4yToFVO8Sh7M+qNez36TVSoVLj1+ZKDSi0s9Y0mNj9csh9gHIb0Wy
PId7G176YuyPQvl9pi9WBQ==
`protect END_PROTECTED
