`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OzQHLIox+NoMOmB16yArcZ5ZPGdneUrR94VFbRoEWRVTPddk687xxP9FZri/oPwP
XUKDzmbXFHkEsS7FDDVjaURQPBnvW149p8gbQQvGesSaAXQL6fQpfVl2fObYGJzc
Iw0PyOr/cCmjOzjPFTS6ZM2W3hKLn5VpLMJ6ItbSJOcnjYbUqTlORaNQYja6KpOX
8cLf70aQFu8gXV/wl13BsOhk/AjJmFtusbnjtQghg0XOf9nuOWufnL1js5qjCosS
Nqhils48IhS7JUb7zdBi0QxMgS9JuAVpvfbpAAVwl8QsBd4EGq4O8sqbsStQqr4e
BabOfpRAZXgvwfHWEpjOOVBQfBTgII2pAFFuDM6kWYWeDaVkhcDnsazazHBszkk4
wZn6OpUfFNMKv+wUJ6aoUUCJmjLtSZYMmDjeChZysRxRJ1ndCwhb66yHxyqQpe6L
y7hODHu3UxbGmFkXwfCPvYXKkoTrOBw8j5meTXmASlDvjdBPWnZPRCgHYDDUFSFi
YaPrWv8WVRiB/9y8fP+Mcj1sxroe/H2lrbaec6+7mneBZHZRDQCW/camAnGek4ye
lsiqvFgi1lvpIyYCCJHr1JXTCWbEFDw9u7xL+8O0zEpr++dp9CD0RjnJ9Jkh7kvF
Wy5P1y2sb1tYJOY8aUJpeMc+LTmSukzN6CTntjHP7fyMPbgiu1zVh9LydABkN3/6
ki+gMRmuk3jUrtU31k70ubQO9gdGyiYFA8inAcUr0+B/yf+eEj8QXANxjsm4zn7Q
kds3y071BqyJtzJlgOG4mmbWYLps3myCXE7n7GRQjPKVw75PloC/4rC0I5Vyzyym
LXASVFTDcHebbiW6IcE2HMEY3DdxVAoSWIPzqg58qeec/MN2i0dbb9eKl7iug6TX
Nm4h0I1vUCkrnh4j4RZPAIYmpgCQMu2u/O7GHDnEfhKfQYZdMzTCKJaqbQtYsddQ
ty8CQHeN1lfkV53GigiOiWmyDh5bnxRYVHXx7o3HOCf2Zn+CAvZyoZeN7FMjbsUH
1omAIviyGxRX3A2jnlV1/eUQIvCoFI9oxVv+PCheNHpvi/4Kfo5Tdo5NjtoNXXmo
Qr/ViurB8cPq6rMnHVifIom65GPeeHrFkIQDihCJibfeIAqe9suxRBHIa0QjUQ/T
YR8uCVCTEfgoV2xtrE+8LdPo1PeauZiC3hJNPyFZ4/hQD/dnmHaszzDXK9Ba4Q9s
cshKN3zydFyNWWl1IuBkred0/T/buJ+9Kn7YobdVl8pCFCtZ8Xspgrqi4yqbL25l
mxGr9fFjAuAd90PnQTuW1rSaYwj5SiX26k0IGRIQhIgnLBTd9cIKrGARfBgvWHXf
lbDpxkyvH309NP2XxFVu8wKUSPBnS2YNhsujNrKPL8/IOQPQKIlI2ZxFHfkMc+AB
or//GDgGqC6VZcmXWjvOpvU+7SV3AW0Jdl/kfEM5BjA/AGt7RMNCfWKZcCeIrUC7
p5YdfU1vqqK0wXk7tLeGA2HrZpCrPUvKpRUR65RSvC0RpsxNebK3gpnMnrDWNH/C
pH9AOoH4qofTN4XaQRiIsYHj0rElQhLyBQdqbLfTir/4lMe9f3Pcg55zcz/Bfj2x
XqmwRvJL3XlzYiam6QfvG2EAXhlGSsVYa155UNt5BpEAU+Tmi+x94ym/bTJX5dPM
CehFwT7WIFM7BdI0+mmWZd+guvibShz8x6V4pmdC+sU5N9cAqmTWVApQ2tmvvpwm
15wIhFTzIvEl5R1sqvzD+0puoHBGb6Db6ZM6326pxCOziZplu8NjBUxvDILqhV/U
fuFBi9UrPhWxl3GHNCNJsEsGFCce7nFfySPTTlkEwea9sWpEKwbbkbXeNe0e00w1
TP7ZiL3/lhqV+K/ig2FJNOeKjUELxqkn1UU9+oPGpMOeI+8nRcLxA2hvazIRke5F
/IDgjYtkJ6UZPjTd1j9g1m2ODi5kFVvRSKEH5HK5AjW3qbMQgstH4Tr9vDzYpye0
wZfca7ptG1D0nRYbpKtkbRhVeX04yd2iYVWNR3+YYzzKinrURLFPWuS9WWRjF3Ze
r/9J/ru7HFSnx1RjOqN/5T20q9agC5HjP4/putM/sGOsG9QT0hcLlrErE7+dnpkP
wxZk58rCpyBGFhWWs8PEuUxV/gIfHVu3l9eseU+6xUd8RLXWz+uwjTTvRgxYDuB5
/BqfjCn8aEmasm6DMImb1HIQWAeSD9/3+ANTw9ZOy1ETeKWIDBvQ9e92Hnz2HQVK
wyTlBR/TKwg4hH1KhynZOOlRXtPS9FstGfmRsUsXtQoud+HAnwhniKlXdPluuGtf
I/hQz59gZ+O1dwnJM6p+h3UYhO1q8hDNKQLDAwaYWOIe+YUx9iFAnuW/KpcNvKnr
xbeZBhKd0Baj8+sQ5NcxVg/gY6u/BamE2S6hbsJ2I3nrObIh6i4QVvHTuSsTrSoI
bbowbdnZ8QJHvZu+aq6dXYVDxSGvsVrFiVRLjWiqGdypNRyAIKUf5AhBEFe/pYlT
8CkTZCTAS5cmy5Nanl0segwQxxTVwo4n+5+EEYtlRYX/nfmizwgZjyJT89T9qYk0
OibQE0vI139N2U5LsxhHaE9q+w4nNS/yHQN+ydl3XgP1Qxo0uRPfpLTOuh+w5YoU
aLiHgIQE9DLZtXFTy+B0MlSohDcFoF3ue1LDPmSuuiB1D4WnwXt/DYFLcAS603Sb
KLshJOaytPNnGXwjgbnKV/T7VwAODwcvH2I6ZTGPKpe9qkEI2vtQd9mB3GXKAFZ+
PO0MhW7JUSYEDa4lV6pcNW8txWjdrUNRUuxFkOGFaJ1TjM3uNZieTkzYVuLGyhNI
J41RLwkIR/Z4SGLhs0Y91LBb8GskMhxv2MAluKDGMW6FhmIxFCzYVxvjgOZZ1hW1
ndeC7DWYx7tknleEE7wL6yiYetU5d/9F3s0kqwGGNg7d04A6nXYKBQ24p6FSezUB
uhcZxQq7AAB0hPau4oK+GX7tZutgpikS2o/Y+ANs04TkcJ+ucggrTf78XvRWJXzd
d9PTNI/th/YXylpTkrbqUXDcFCHfvLNnzCIh1t85MFd51Aoo6Zwt5oTDmRkCVMbd
DIz9zpqSy4vzl/ycGUm0kKi00Q/DP+ouCsT66Q7nEjUAGr4nGlDicJV4/vRqR8Q5
F6mdjW2/bSqRL1fJZ6dUitSkGOa4Pa/ELS8hCmEzWl8yynZ2kYjT5hQ7GdHUZikV
66kdj5sAW8txcTSoeEWil/mKE3cKXrZ1PJNzUXWOExaoVq35YabQ6SVT6OxjND6u
`protect END_PROTECTED
