`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PbrFtrD6nZ76MF8IOB8uCjiN/lM9eKsAUtHxrWsY6+75rxJMPUA/VDlb7bUZN813
XskbFTKWW/OAwBqtHndU0JhlUfgETMCiTeoe3O+FpPfywjOVR87AbEz49sh1qZo4
fFAO4Kw5Uo+8CnysmMyrBb/1GlAvpFskYKLaBdaTsRrNwWd1Ex+K+Ev5e+XRUDpf
/RMBaB8S/1qotUFJy2ZO2OtIEUuHl8MOOyWCGXR+p2bCj8WUD5RuGUhw2FfwCVph
Jyf4TFVh61wXFawH0d82/F9e6VEoXQYVG0gg4DU80Sg848MK6mmbjCVUMDcQBQVQ
ETr2K0YcJEKM7zFla2QV9VQm2Eih6NAgin/TgkvIwUktXDEaMhPfzcYW+v3wpGA9
Rn/R2+oFbdxzFHNoUMQwppudltd+IB1768LIHOclk9KZGA8UgxNzgP5YaPfncZHN
oA/4soY5SGXhe+zmaSHTqdsf6pidT9//NC2aJZCQPmOogh8F3Oyu6ceuOcqf2QXe
mkmjbiNk6TcBcOdunG6TgbNubMkgcb54j66hGJA079mmhA0RngxnA1jIfXV/7koV
/yyLGrTI8zSL/HM0FUZUUQ42B+p41P7cYSMgtJNVx3e8mr8HPQaGGhULVEivqkDa
g5DAOL95BaUAO9mvGRZrEjErluyowtJ1mdJT5IjY4iLY0P5JL646VEzAMlwfvonB
JjF83xz7W1m4nLRKZEYXJeJa9+2HpqiDmyq2uL65HT0=
`protect END_PROTECTED
