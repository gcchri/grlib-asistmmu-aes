`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1deePJnQK7jXyHq2i3sFFp74n4zoHPIxCzBm9KU8qeggvMF+RcM9N95Nz0LW5r8
FS6zyHVbihpREGywHNd1aLjXHcy6a8cHIxJq0FzAGPmqNGFh9PEI89D86PQycpsZ
J/v292xtIvb1L+1EL1PrWJBin1Qp2t2zAb8X52dthRT6w9ZB3MD1t3r2ySl8kpOZ
GJvE3ovWv1jdc2ukXahXZHCzw5An+GfR46mDILV5sLBpox4OZHOtMkKa/tOtKhyn
kIjr0ezCs4VeoLFLrVVc7rX5thecoYSma8NJrLmYyS5xMnrFtyJOpzmPLJBPBKvd
O3t/6sbNSPN/mmVdpz4npL3IIS6FqWoxB9MQ1AIK/pd37jMZLBzFI4pcicGlhM1W
JY8T22QdH1kOviCVzdVjf9maIVq/6GzVxrE176/LLk62+kb85iEWzshqVO0NksS8
f4aKyg8qnXiPWEiNr2wBtmrYxrzCzL/69w4Ij5NDiU6iBL4NQJwOhKR4YuDZ4WEu
mBpSBqT6rVVbMvoyyMXxkP93m8i0hQllL5f+R2qnJ0EHkTTy2HXDc/gYwCJFyyoF
CqdaVTHxsr93IockfVc3WzT9cTFK8XLktEJ1zjDpTX4R/iYFewWafPy6937iDysU
tPvQgoH54UZRa7ecGhJ+NPCQlCBk9CJkp816jwmzr86cn04xx49jYGFfghzjtk4k
bmXZyqH8rkHj4FMrdIS9s3cWdmcK9G543XyaB5Jy7qvlLGQ5oWIn6Brflcypaptp
nLcQvZS+JUfZZKGpOXuvRgj7u0R6Sr3hDM1ZzdNVaV+/MAlOpIAlr4Xr6I3tKrvK
TUu8/iSC4E/F/4HAxeRWr9qEV+n6Tyaf40GheSluq3xAfCqXsfFEQTqfIWtoXukR
r9qFFUHJ5HcY59xiizy72QN+XzAuCnuFEMy5sc6mrVS9ef/IxL+1ELq5CE3U0hdm
feYgFPivub60CHY6kvzLwl9y1mtl5Zs0B4EwimGHTzycmBU3TiwjKPojgyk7lW5o
L63XAKOkfvMQG3AGpJKxdKf19cp/A9LhfYPkSbQC7doAtz3OmcZ/WbAXWWUGYsZW
PFmlCTwjYeNetYA3jOtckB70urYo2Mo9f4bWHAabOuu3F/yhQZiCrBC3XvkhQzIt
wXljjs0QiyJcRUtYONmBXoCNj5mVk0D3+5UCrvAqF9/A40562VoDdI76fhGDAGzl
zk4Sw2B3Z0o4gKS4y9xNYu8e5ZrtF4ecczuXoXs6P3q2TiLWnaXf4bucphMoG+iA
lq7HiGkZVpdgSxtiUf1DyoulCUvTiwavy9Ac61m9myJ22+baduyR3n2xIiE5h4W1
in/ffmAHdaQH1g+meP0RAX6mYCA+Mf3Itlr/NFkalGss2vhuwDrLS3F8wViUihiW
9Fb4rmRGNRMS4Ds0B0A9Ghp4hgRNh2i6yphxomk14ba73GG1S0jYd5B+fnj7EhML
RnpEzXf9Gtfei1kLN8NHfObnCdoiUUfBqGP6FLrCOwefMzLlit6vHa+7tphh2q1S
qLQapM69Sx60okFloVfvF6hhfzuN8GNUjQPvhIQwAZZZMoacubmtZBwjatgmcO7d
GXBZ1Bi0wDco3dfiTIetlOvzjyR9GPfsoPwMQxXEq1tE10ElkiSxVNbWnrQ0Q1FW
EmcOhAFXsno5UdL4cQtQ73k8MVWVJI9M+WHU2LsfIS0oAfTlR9QHVewyqF7w+ral
frAO37xUnUtr1oBVtmXNyvKwtv/IPtzG4louFdH7JExE73b3Yudub0eZ0eBDJuoq
gvoiJAvjXYxGQ3ua5+ypMhf74OxCM3oWehRvkXq6pG7f0xTSjwIvGbcH8UD6bVvc
T2Ns0t6F3+DJqk3fTqGgt4WjWZbHciRhDxbJYa6IEiJOw3tHBVe1F9eU+u1AvSUh
AKTttp6iwB5GjCUxLMPiLvDC9A+MX39AxtXidh59it99EGdVFYvSYBmfpEUEjGzY
+qrW4U+cK6IvQAVwBIHIJWjrVCs9q+gkLYY+U0W7E+ieo6s83SMq0Hrfxa+VV2Ac
X0B/jo4++NCNRMGaxeETMlYExEPBl7lrK0PY5wmf1OK/AQozZAcach13tAzIwZuh
jlyGQpOruFd7h25ZpeBnII0DIWRQUD2cb6lH5Ds6b0qtYCgEW2bRxC/3HQaaMSQe
mh4qZLh8HmWlcFHZEmEAt8X9ca9LIVCVU9i2ZQIYwgLI+e66l4vxC9RHKVzrlUkh
2rL7OKD3da9zFs/QO7WNiONgNM33194BuYuIcIWbx37tbXl9rTVISz1Iny/xrX1t
uT32mwVv+vz0PA7G3wAT1VbgDwoh/C+3yHYExbse5nqUFgTi1cUz6CuyqFzfK16G
lcbvl6NoE6rrvYgwpeNqmkLQ7g+DYj3d7olqPASjZ1/E86ODedGxGt5RICAYCWtJ
X6umdQXorADqkI7jybjRDB4WUYdtmqRu42Hnsh5NX4hsBJ0rld/lPiZE0JzFcK/d
j6wI7+Jaatdwm85wVizcesufSNbtHQfqg8S3WQB99j85qBHyLXkkKYo8xScACQa4
NRogPeJk9+tX+G4QxVEwbU0GFhobkhB25ObyyBkjWOxIi9FhOkSFGZYXDvNxo7+Q
q5X0P6RCBYHS7LJnl7XIRP8oECoC+0AxKN/MayEHirjyf+kriRjd+9oSzUJAiHlK
LDzCvaEjjLVnKu+n2nDdyRuFsdz7+1+DrWkbQoyW1KxbJkYUF9mG0JJ28WkWNwv9
Af5hk1f1k3oFdOzV04PVTfKs27bhciGb6pLOPAktOx+dmcob5ORYtartQ5pKKBPM
+0SmqbtoiinejxK9dNa0KHXZMHDp91IhT4buCQkXWqsVMM1wZ7ZksXJXOHNrLxyl
xtxk43RLk/DhT/vMV0jNbHNkCZZvoKCBRgzoMAU8/IIOC5k3BwjjCoINa4IbClJV
lb9Rqd1EE5BXC+F+EWSlvMYgCCz9eLyLHPvV7h1VCOUPxVrYTjtAhsbJ1Q9gw2vO
ZEhf3HsOPdq8e6wDpD/NeXhul78QufYHId4FMcJg3Z3hNtc3RCsN7BYyptouqDmR
T/Geoj/JEPN8CMTQ4nFF/8QhbwdKHU7eTNEUcxjY5TMrhRhiyYWkzKKDqU4xVJqC
giDNqt2STbFVKMAFgFSMaj1folFOzt5DkG4OTRxBogWwFkaDoa5iQQR6biVjLLi4
pwVrbv2D29gB+BP60vXfohWDQUaCh+p0g2HfoYvYSzV6jDLSS6yZQY6CwVJRczar
Y5zH8xXUTY8T+L/Ier0Aed7MQ4p2y+HT2WqMg7wAQXc/hjOAgKbOB9XXr99XrymC
xgDjB0D5wH5eaEcAuHHQw2kmYKdBWY5FSQCvTNWEYM73r8v1/yoH6WlHZaCGQGC9
Lm6UWsTg/DsP7s2co3m8Wgdlw+NTUUBrZI1WDsJgCq/u+gG14xLqC3v+GzYau2vB
c/QzVClg44QBbhcgTN5w6O2+s0bBzMzUFNYQbz5DXHpP9LwgdknUXh8zSjygnnas
osUxOfEN4rg9s+deic+4ijsVn6dcXvd8LzeM4rVnyrXQa4GmF4Ncp0bnOidZJTU5
as8vQlAztb/B7ugaRqMmIc1/b47Q1XR+JH6uhp0IPxfjQ8nTWqTftrL4I1XqB2m1
pOi/jUGCjxWt90fpfpaATpO/nNWfrOdo/DPpPSS/CBsWpxphKQSTKopvTQxoZMAl
nMC8cSQrz0H9NktBpitJk+6Wut+NEY/XI90U0DBgkLG8uLVeBePy5hgU6CoEv331
MBYnjAjrS9rr2rocBQZlaBit7Rxuoz1gvgsNf+VFvCJ+al00BO0dCjRwW47pmQR/
TK8QcYNFifHVIKzkKwWYDi8fHnjlxw1qSepV0PR+2I7DRb+vzxArXAxM2moiaLEW
eDUeZDqzc+zaxdM3GImo5HuDmOiRpUWyVS7gxw+FrZlrCcgPJ+vm6GB+rA3BY4RO
z5O4z4dYPAtpgVz+R0pVn7ku8qvtrUSXbPpzFszOVDox8vL2IRNTTRM6GoCAkrv6
asCxt4Q4r4+6LVBdkupP3rtDcXXfDez93SgHyaoCAO+hPJKNCUplX5I4A1eCQEKX
W6aLq9OlLuyH7HKknq3aqvwvLxkfsE+xN/0IwQxYhgIqgpncLDBRPDIkniF3Exgr
ITPpCLZIBy4gwsAj9CsipfRQYK8sq4qsHi/BnLhRDuasn9zCmtQPWzJnmmYCIFeO
QUO88mV3JHO36KaHlKjQN8kZZkAkgnfJUOyk9QN583FBfXPICtbXMeNXI0PKvVEx
nqRxolTkmdAhUWFGXWGZzu9G38xjAir48qRxFQ85FYdS0jb3ch7YzhbDijP/JYGE
PeSwh8aX7822M564LTzltDuhza0aQ5WYlaiFJTTv2TMngSkX8KppartYi0UDxDF1
o5fBSEMdDq3guLI6ADk2aS4KxqT6Daehu+SA3sAJONKHmtjGBNV3fD3uLdqj4nYV
PRwd1s9+r9/kQrCRPpTuf52QD4Xv01xaXOl4tcemwj6c2qZIEX0mXcvQWyU3Y3hq
sq9RPK9TEiytVnXS7UMLK65NgBGXQ1xIjqP17Hm+qy5ATJSf0BjsAq9HXNJv2nvI
Tt697vs8H4ULwmWzx6c1ZzlxZBOPU7PQFPbNMxMjdbiT+4C2Z+6YFHqls/HlLS32
aHQyjRY9bTpsYntohrLZN05CoH19zj607Z3HUxb7JaKoOJYkjOYttd1PuDnBU77R
QvkfYaqVXzYDVQcdfCAGGVpR8zRVCyAxB27Fw1uJy4STxx4zz7JbO1c64MpVbuGY
bptnh+yR7tIBKO9Eh9H/pp/CazAVs0wM2QSDx7r8RcAiLkmjnYwcf4Ch7iNKv1ZV
knLUQy09ye1O/p69vBzObNqoO6Xg1EY5InS+MFW0JRbUoXwK6eTmt7HBlc2CLS9O
KZGwyuvOqcF1r0wWoA7TTH+X6QrJq8KSKWjG+0ImML776e+ShxPjC6VlMFgU5JwP
2Z6iT7y1XXkDBV8qkv8pAJeLcuV16D0wM238OOpUMEjxqAct0KglQFJMCOY1j2+W
Bs5e7jnio3XpIgdUDgswrTBFWM4IUmvihRUnEvWRchKul2DDt4XRyUT0EUV2wVtF
o2WpDlCvoosTqP8vbBH6IF5lS1efzG6bqNOCNG4VbzzqMNad0KWqyRcv2MJYHkD0
HB93lPtOlZucRfJjlzYysdD+Cpe8aZFpZxpLz8x6KbqrZYHQjqLLJpwiFHmuLI95
fJlWlZbecJtwNKAxbSD9l5bvf/RXj5HWDDZY2keY6C0XmxQeFdMfv3lBovQzW+Fj
acrYt8YKTqcFW0aDIIHVilKcA9Kv2GuAUOjF/zVIcJtOR0ymtXku17j67u5tyLWj
SK1QshjSukeaTdRcA7NLWC7QqVJJRi2fSzuKErALQUjzshurDKW7+EwtRXH/yIWt
27kBloXXujG1DtllMVh0Rrh/fTNsPLDtzK1LO2oFui+UqzozTRT/g8mzdSeQilM6
qWeNqWktE6rsBWD0TwIy2y/vf+09zCRQ16LzGuz8WzpX+QxDiVPtMtQ6Skh6wV7R
y3XeyO/wq/iQx53bG119oQcxuUOh+jCQgEcCu1XCL/KwLK271WzWg9M/ECfLi9fK
BUNRJa7BrTqYSFxWwCqZjuSZxKWlqOcIewxJipahzGkwluVwHmkpzCZTvbzF4+dq
CF9YNPkGToFfrDZsOL7rq5jIvV50c+mCTb0HGTr600q7bfZIMVNkKa6xsuUTQsBU
ONyDtHzVCzBpniwgUWh2e+/epwuC2dOi88GRH+ShcNoECKAu8rKgkmiYcb2uHXmO
qhDjlSMoS25j0exN8F6gJGoqQExkOmyxpnPb4OvHo+qe+sLl1jfdXRFI7veUs9DL
dEEtIV3/e6LZogaa4cJfEVbDv3EIG9TxLqJhTbkLNJDxj7wvKBaAeYjzDy5lfOcI
01dBqkYF9KowXndHNtjOrrvxjP69G9SST5dCt7HeL418TWAkmzWfvB9cVD0HXPut
VOtzIyALINTgbxvDPdsBa4Wu/NjsnVR3yxp2PGvGGTU71pyweX2oX9ImJVMwix7r
C1evoYGfA0OI5CIn0TB+HH6S+HM5Tk6lJ+Dg+LjuMOoU0etkWPYnhm4pvfByqJ4B
s009bB0OlBs35+ucX6RPiWWnBFQjL+gweEHnLaIFi34VDaR0uv4MwKj8y4hgO6M8
4qxQ2B3R+SyFryvOIH/aLZ9H1uSnZO7auBSELX6Ekx3jOUI6tlqkWA+woPY9CtmK
ZZZzYj0NhMmw+//QCvMeYZ2CT7ShcW0iybL9quVFtHd6p7jMsLBvc6bIiZyMpW4Y
k7vZWJnB/6Ejc/IaHfSDobZjOshv/+niPE2dV3IvRE3G+p4aXEoYSzpleaF25RYn
Kc96ge0g8x6z4pRgG6KID7GSmav8GPuZdN2OD06E+r222PRVpM1m29SWCZXn9vlB
Vkq0rstyNAClgHjRfoajzSIrjn/sp9Yoo7JackX6Y/V8EKm6I8E/5L4N2MZ1mndt
9QS+vigPZf1fGmS0qOYByIwXqqOOGyQdsgR38xCuEX/BLB2/qgT4EO0ltoUc9jnx
Bcn1a13wWSwGals/CCnziNQRpOqkbMWG5dzxLohMILuolJvVCBP++V77ezwJd6es
JL0shPiuHka1ENvUuMsC8BUnNh0gPrXY1cMSbqCryQZiwh0TYq88D00F+HGnJ+86
b/ZPCkpo8QcUJfqsKp/HuNJlvX/XwLAh7rlAdv+TRZOan49KC9ADxId/oinQ2Cod
WZorBI7+yAHaJD4A9lMoOlJloOr7ghaNAx6KRRAMR4NP2lPTLTH1ao1q0AOguY7l
W9NsQ/BdtX7qFDOi9Wbe4zc7UhhlYNPh+/cqTZlurihW1QrKmg3z1PZtRa9+u/e2
xrrkUwiyQId4gNRGtDfAbGcm5eyZFas4Ed8WRdwtOYSV1EGI3Pg+vnONrPBhKvZW
KKiSTgTbaEsiY4aOX5oIDLrtEC34OSpdunJVysnmFywdU3pkNivaQiwXFTRy/HQF
cvnmmGU+gUoBaIbZQT3n8uXD/xcwLppH5BdVrwYuJWOHTAIV9lvt3WOEmcRyinLV
SZluZwR03iOI0AKq7M8DsjZwOki07whJ0WP13NrqKkj82vIdgBOF+NfK4HR3KGEY
isj2xX6XpLwzjlFXganad4Pj/vBGZCQwqH2ehKvheo91Wagr+c9vu8eoMuVYEr44
o18XCYx+K4qCsdRz4saRQV+tn0IGAAVD0q8C2rfJj8dRpa7x7cV9C5SimhTRtvOq
GQM4G9EMHsI/4bAUyckP2CZPeYg5bCJxZyAM4YEwYdT//hO+deinhUC1czLTKxed
reDGd2c4P18UTzAHNY8HV36LA+eyNvhMR7Bczy0yR6vmKcWpxUudtZAWPBZofC51
4pIg9OyTqD0JhnkgCVf2rXpThWjPDFi5+2iUQWwDTcMsNkObg+GANHg03R89Z++W
pidfa9L8EhmQlUtZLiXFo30p6xTNoADawPA65eJyfd4yjcJgs+5MA2wpKeP6yUJR
+0QQT24tFI3WTcsnenPY0C+MLUjoLdQmPe9Uti+LT/9xku4GZsShiohkeZpyWrsg
Rp6cT1uTHWgXHm+HKH78lb+7aOwR6ninvza3lYTF3+Vg8nWEVAg6nGGbP3IijXD/
IF6I/KyZuOBce2R/95sDxK75exSRZo/WDi1ad5EHuUVniSr/rg82Nm8w6aKXER4n
siJmSa7S+4QLYqy33GCYf3QRhduDNqGgPyYbNCE8V6OIoV4P6p8HwDkl34z4Zw34
MTpRx9fcn1aStcMw8Fy8XTaN2SLvZ1gcMdMMloqpkvaP2coKGujnGQT9/GDIVYoW
Mzwsfj83nnQfTzIKkBR8z17JOl/FtjvNU77/gV5o2MlstyX9WzNYjjbpQQ3VVkxF
mwYz5xuB55luxVGpZGPzEUrS6zRkCnwSiCBkEI/L6x5B070vBzz9McOTMTxiI/3X
1mmh9xJNRHonU3ZIXNqWo+UQG69aK9hU/Fczz9KyrKMBpaBFN7oED2jylw33/0lF
+S9Xg8kBn2s/BSomEF/RGr98X/vXj1FlDB9LoaTXA47x+/UtUJWXR6KUzkbHEAjB
eATSrTQC4itGCfjOJTHk70Nb+PTlhGSznca4OXiKUpKGNM9EBkEsQBy9FpETABKh
rVVZRx5DDhWBRXzVBSug+h232cAMzDsqviVK8aFzbKqIyZNsMKMMOX3IJojlxFro
BVsQxa1qj73jhvZ8I5+n2R9X2PKCZU0wxOKfjQXaS3yQ2doVXPUPVhQwjMtB7tQy
otryloriMRT46CvGbuIG1ZkP37VaKUdfuKkaDUCdccakoAm7xq1M4A4MQwW301Gf
S67gacDkBQrXaAPW9ptvRHVibbTjmOEV/sHFhEqYG6r1qOQEQ1Puj1jkNNWsNAlW
0qJL5YuvS2h8DBbMWp0QAhO2x4lV/aAMzdZLAp6xkk2+8i8tKsTKIpIuoLxDVbpN
Zh1ZpcWWK+JpRcuNxDwWY4RDrtqkpXaDRx+pPTaj4N2OL7OBBpwywJEuF045Dbn8
6UZ/DD97hojMg3nLT8+yQzWrfQqoxeUBi4U8kSGSOKHJaeR51rF+PVtFadhGsEA8
IigpiwJhRy3s9omNdlNUcdwukgT7rEbJtxRFZI7wcwhXGYfh809g1dsRKBWpUmY7
f8/IMLbW4ivyjGGKNDVjgXpXp9F+gZT1sIyPVrXhrP+H+SG9Z7qj0glDKndDNecR
ujoyHcWZr6aTuFCW1M9o5dLZxUGZZRL4it95cHmRwxoqKbhFeO0iKdL1ayFJvo5b
vxCJ8+GKBKCzsuT7zKccUQx2Nqxfoimh6sFhoGN4n94TWaN/hxnpj6EqcCzTpi5N
QBC3NG4RcpOxMdmGBdkP7Ko81mbZk44IW2jjE7hZxgyiz25JlPcsW21bLIEsLEH2
MViGWAPGfRnMMfon5QrJyRcpLGx0fewG+y901n76VW2NpLx7a+0RPciCDQNCYGlX
IVzSPWo/Fm+hGASkuo+sWjD5DdL0q8OzpC1Axk6gm3CEWdCB0IR2x7zMZlm5MfZ2
GJAqtq1y0n46AwSAb0TO5/BKx65dtZa6mXfNVEj7AGhsp5UQ3YTQTN2t/omQMra5
w7sBG0i9c1AhFjw53jDp9/5v3nT7zAEiufH+65I7DZL4vRF5BH05L8LMUXDW100f
LzS3Z0aZSFiHrf2TD1kz+pgDKTxIQNuVCATh0R+yZZitCOu9xV5a0M27QJ1fILUI
qLKsAnapfBBW7PXlxFYgpV4p/GzFTIWEji8wOi99KFhAjOqn/Np7O0aS/IRgPfJx
c4IRjJCMS7i1wp8W8Erh85RsyXP2uDJ1xVlB4CQAb3n8hR6DbVOiVH0H2LUfd7RD
M5pCpTqDfZgwyJAcq3p0GZYAmUodI3bBpmF0mkkZdSsfqyub+HGy5lo7EC1Qg90n
v6bZCBJ4DDlTm0MsD5nL7dd8imQIPTQIhSG7Ly0ucF23JJUBZgRo7Oi6hx2oQxxK
5sYZ5lK1MctdJHcxeBc3gDw0IF+QmgWzkmGhiwf/WTxi6pwrjneiegci+ghKPk5S
dzWXo4ydIQcex6B7Ve7Y3KSuvojvVMIR0b0scDwJVQqS42LB7Nx3F3EamyzqLYOE
QdPxHaFJLKj0OLaNmprNMYAcreJwsh3BBjQsbCgmiEAS2pKGtSO/VlgAMtEMw/fF
TYyXSFHkzo2LcCtRmfpDRDzSwAIekKV9hWgMqSSrwKbIe4M1tcfFmjPGvbNRJl5S
7z1lViGMS0ymL35K3uaJ8lTGQUuAIu6wNeZDditV9fo8bj9PIr/gvVRc/6JtwtC6
EhXvD4tRuoYVpCGi0DcNsW97CQxhUxTz1qNluW8c/kDutRRWXbnIAYfB1iK7pEtV
UGHo1nQ62PGD47NCLcaf42sE2SiX0gSSiS75ai6jePBmTfgGO5gr9QST4WYBihX6
Wy1mF7xFM4TP46a/qSej02g/WZ987qW2cX5712MobdEy7WoH9tLvR0eT86xeZOny
QzVTbRgFnZOlQ7hJVCIC25wytaN35wSOiLp4BpAtEy/fnBTjs3bX+1JkVj/VSryk
Q/oZZA7QSeloei2H6N3qxVYlEa3BvLbAL3xFGENncX3qUIjaCX11F8n8UF2Q+1Uu
d+FPZ3T14Nv6BOVqrA4IqFgTFquXvLJcIdLtS84uBGa+rdEmm1A9txPn6X2xmlN9
OFUNwoGa63Z6B/wq480KSUvhClcEaUEFdT72Ud8KaBgs6WQQKP/Agc1N0d06XDBK
ypI+pJLIRfJZaUTF/8OiCwtwL0BxZb11SlVUi5JXPff41AEP0P1lr/QBcgWzt/W6
7LpyUT06n7dPKrJ7h4C1ZoGoKjk52UKogDcMHd0+XxkD0FEcqLrzy88AM1HzxZiU
fXil4P6jE5If+CG3OHj8IXEKm5aFwhEXfxqfpLL2CU67nIMOd6mbgIi8C7odaz4B
Zs4kzwuSA/vS4J+CWuIIA4h63NCxANXtvrRQNh68LqmgYDQVjVrBrRb71pwW8h9M
P6WQmtAepRu1NGKrEmtTw4MBD9QMlYETUaTjkuUFJUxW3HOsLhYRsqzDQDCgzuTl
1fNaeSDIzepBHnth+3cKBDhbeRUKbnxbV6aDfCqgpz4+4MyXQ4zFJ9KncB0e5wPb
i6Yax+v0OP0IUx41zwXZ9oxVHC3ZuADAP4idzg3GlkeemEQC+QlLlFGF0PgKHBeq
5OEOL9MWn/zHJv0E/shS0sJSpWwJqkeLDjeAY05JjOiAO59opryu0ZpPpWnpo39N
B/u208dlMjHmB0HQlXSHuW1KITdTHqoQkvnrbfnhe/3pI/saNdob8873ASXD0+xA
MMSVDiQeEd/ol1QMJWhMPOdXyVJeW96OuUbG/CTkLD76GTZ/YtCi03aP0DFR5RUt
nXOzfV3WZNv22tVDipAtttYe0sCb4HzQn2hJaYa9Ckz4h3bjoEcDkfuy5shWxERw
YJxK1o3mQZkdD+wvJ3ROxFScq/x9pkvtk5AbQWHcxX0PZdwoWapFTYAnj1c6kClR
5unbRQbRfyAOUk6j4zPzzk62Prkpzs58o9Mpywqn8ftMOtvOgcNU2BUBrnffPoFs
NlO0IDAa75h7Hss7IOJB0tXX4ys61ZQHyanp9MHRvXIm8cm56ZnRzxUIQKc8SV+A
B2WL0Vx3MnC6kQ7xWwBj7girlbJWAredWLONc0h7a9Y1QR7Qko70zdMY/ijNFEAc
C2rX43vhTrbDZGFmGlGc1BtyZ4w9PA410z8kXP+TfAkqpQ0vL2omJx1WkRsdf/QV
DCkL7Rf+r18jOdANxYO4FsVhhzoEh4mjB3tlcwlD5XxOHicu5VxUw6zJCaRaRCgc
vG1YuMkTC4rVUnb7VmwOmtec0/VUCsJfmQ3OixwvnBLqy9JWVy+t5MdeIeXYAlC5
MxwCMzovoj6nuNvr4HYL5HwGO/htChf5h7q7k/knII8mnlZqmqnJKj7/PHeAtdi/
h3AchPrdJpkYI9zmfL4qsVbPX55iFWa4xaM34Ha7/4/80c6GugB8KRoOi626bQ3u
jw8MnmcnCWVGlR8Rbnx5WkagIlcp2xHA7rqJDTft1sn2UBUeapw05KNnkYTS5ACt
Vwx4hRDtn6ob/chAkw1l79ARdGCOst/68y/3+gn4poyTIfXYfUL4MZ6H6pzchb77
ki/956/bxTxmFAgaekck59Am3uNvtcKRl970RdbR1BXDWGt/ONG32mqP2vOD/a2x
S2UurONSzLZmC/CW+Kf5dq1NbucYcl85oKRUkS+YiMYxFRyDOS/qn+hylBSxtikb
dx4qLhluc3vjxyKY9bldgrvPsBBK6pFmGKDBd+p/4GDNSTBOu38vPV4lBPgQQmSF
JqUL45idV/GTxMV3X0YLdoxX6supGfSMO0up1NFO+/dWD5S43yaZayVJYettCmfu
FvVzGdHo9uS1GXisTY6yQteLocBrjIJZL+3enERQDlh+Jx3wuT8mV3SdK2Xk7O0x
w7oU6lvCEZN+ZI4dsNsXb/I6jtLoDsohN8tIROIrQ2CFyfV6KdNdd3FNO9sgOKP2
Q9rGkh2HchWNhvbEEVx+bWaQqDhaobeIuf3/WCYolY/0j9DVskiIJO8sCbTRA748
1mDzeYNZb+qjnk2l0pBjGsztN2c+Ht4k4dYX/NZXy9WdcOv2Z28qF6LYARVDagE1
yDH8WACeoNLWnOhfMEiZT+WZrWmmKWtcA75xv2cDbIdt3AxhhIEWkJS+876oSRLM
SRLmd/joOZlXnh2p9aOnKvAGpHI//dHH3iRoXp2GWtF5M1hbUo+jkQRd+xv5g+Tb
WdXzq2uuCiB3qiYeSxP0dWQMkHyl2BZgDGnMa2yGZFBE23zL/LHtX4xZFL2YaubA
grPf6OlT2Cg5VHxRxmhLTt/RdUipPhAGHCogFzkMOFNcM4UHZ0258hHUgd3S6DOk
+dNUZqamj9dUlnstb8cJAEw913bAnw2q7/4c7SDFAPXaDq4U+9IDUuM+hOVB2jE2
zmccnQUQtePPaFkHp57WWUpiGXl6uibPyYKmbfCQFI2CyRSpmM7HeaWEKoRaYXEE
7sh0mTILpE3fNxuCPiv7Y1J3VkiwCZ6pFZJcSRaEy58OfnQ2SXLffaenfwKKKF52
N0RWRxXL9drTjd8Ki5LeYxL5BBgv7+pAeFOy5R7VoXPpr0aA0CwXdCwUoGcuxo01
0Oai2XDGi0L5azQ/5cnGpTeXuWSKv/3bwaMxff1p/KZDOeMBG6yePxSu/XMW+3vZ
CFW0/Ul+or1qNFYvlcQd+9Q/jpsNQzMjO52XAOA/Q+QSGXw/RoSMovY1X/1eTsAe
7IjiYkJcyayDNOQYNsNJ/lqsn9MPPbvIjQY6gnwAmOalZWyIf2t9/A80p5LJ8gEH
lgD0ugu/znPO38iMGs/7r/57ldVgIg+FUN30orponOYUL/cr0hbwVhzzcFMxyNkM
4ZtoaG2xV+gP1JqWc+gmRGdVDS836yWyRF+el25ys3NBRkpokVEOveDdD+JncHd2
lVMU304E4UfLYF55xI5DmIHqD9HD4UldYAhf1rtgGC+p6Aj5J/Tvj+FQU2rDPUMs
URj+su9AkItUTeIIMeMzWA8xV9+ApOE4KFHRZd06kvwdKZM46Xf5IJ3ANhMAH/1P
WvStgvI+2NMy85bqYKxDqpRWEu6Cy0MAfHdUuKlF3fIFyfLLMyaGBTsH5ThtDAhM
NbP+pzM9krnCQB4umsA34icJp+N6G8dx9Xck8Do/dOOSQMX575AOXyMU9CtnCqOg
XAVFAyCIeZOyxjBHRNn6iZQU8mxMb6/PMYd7xuhu1EPes4/kPd5ErYzYQxpHY7re
jQGmvptkzMinndVF9oUdEQZamhnOIRPSQ/xabHKpZPvnROukjINkH9bQ9wtWhnTn
gBgzwQFy0USt33IgBBU38nteIv2gWwCB1XdHcCxrNzsrVVRebcPr44Q7Lons/MqQ
wr5x4cYZ++ulZ5zOebYA1AUD3DQqjwVQUjfK61VTSM5LM58wMmRm4pEkE6ZFFrxp
oMTg/tTmPs9wjYnW67pZ+Zk29U2kgsSj9lgg7BB7c13jD3vb1hipZsMCnXrFypVl
o4BFqlmz3DpInOOaG1xOiU1Ze/08O8tHgww9HiMdtORDlC0u2vOtUTW5+kq38o+r
zrPPR7d9a/K4k3DwU/Gtz3uE98s+kl3rQT//OHMmhzbcvNXs0kg5gsrEtgPewGxE
p1SYyMozDEc6VVxPblsGYplKq0051TDgvICsDlTpxaJqxP5pSZvngZ60Ipl8YV0n
UjTmDaLkaZ3ZdJx0skpEy1+/nAG/E++fdgnCW22y9ofmNxVt+KOEMpEfrJag0F/l
WkemWTQrBLamtcL4iPOHVcZsl9L+90Nm4lz5rBSiDRcY/H134rvYql00MccNNTl2
jc4KzgkmJ57Sg+g95iATHYGfMSA/EXusXpxJFOwTZEyAhB2e2XoZ1YMuKqQRLw5E
7mxzDm7K8zJHBBqLW6h56maBaYAOL/xgC9YNzgmhB7FHTIid9CvWd26LcTpSY/rt
GG9KnnAOrQLtlgy3Lfwe1fo+dwRxvI1Wllv6EHhKV+/C4rnD/VPDkW4r283xVQgk
jwBF99Z1CFmXTz8bOrqyIqqpsGkGsFnDgMUjo2XdAaO1LZ/fp3j5qqBQDDyuLExw
EDuBoN/NA1uEza+Vi5im8RIAMkeWBd4OhUY/3rVqKZRLZVS0KwPlPHWUj2TPVn/H
Ay4ccfLCNV3sGcTzVT67pq9s8sZA6+B5hJwYIpCYbPDO+iQ+yuAm4WlmE0p8mr/T
jBe6kCRLMp4WZ2ldOEQ37BVPZfmPgyZwA4V12+QAMfAoxIdM0+WruiX36z0hBpHa
xQEWtZUpuDk6NHC0qJmdYYWBmIRBTzdn0c8r7Y/GlGFRO+zrTzv1CQAbgQKpYxXQ
oTNpxot55jf7PREsH6H6Z+v0Nd+JER62PYvCK9jmFkY6gChHN3jcBaAoYxyzBJ7+
x1XIXR4wd+6QdYG3szhbS0HWGB2n9uR+UpH/zaqZOvbF7i5Aazi22kLpVH6/IJzf
s2dOrQoHcCrJ4q52kcLRTMqQZBH5BNsvQ+ZriRugS4p1JTx9P9IF9ra9Ly48uMfC
9GlN9lXxB6TX4K6ZYUubvfJyqZCz+kPVMApOkFA3A7s/Z+n+YDn6u/M9GaJLYvY0
VgBQfNa3XEB01q5TpFtaBgFQzyfKZkIH7bENTJw1aG+Y2m2K0aZy/nKavqe0FDDu
EKRo9uDDzDM2/5uAuVbRYHK49ONvmygRjD2V97Boai/2c/++wgNnfcynJx/fLHLy
nB3VvFHxn5PYDPxK6HssE0ei0ZcRHBerTnqqp+ucdOXIkkOxqa3olNUOlJwgIkxp
szn5mCIAMWXgHvaeqsQQjtM8Khs1DwTCWseqh7dwoC8+EInMtGg/f0WSXAcbeHFJ
Q+jLTyxoXqKcVGClRTNvKyB1nwDdThpPeNnCNVp4b5q7QYBPZHa0Wpom8PIoj2Gg
Tgq70NHKKZi9TDK19EqFG6qU/Fp+ugV/BCQW04LOo4ar38wCGlUvrm9Sw1XbXHIF
hszt6evHkLAlvZUcqf0FQALJEDaNKQexAZV2OU0O3mxUo8LU063bB1N8KqPReICX
r6fnaX2eZxY5R//TrOk4bUXsgTnRjRya4P0BSBPPYQnJ2sOMAaxmw6O9iw3bFB6C
M/KD6pyPoWs6lgK7vYbof2hW2vm+QO6umG4LWPCODpH/iGryWkpN81F4YjGq3FPM
+Cajh5hW4u30AUn92tm9tdrnV2lyq2SLY969livuc4TyR/lMTgxKrNVn37O+jM6B
6mkQWWFML66Cc5KoKbBDXiOAcGu+oGWdsyPGyFkd5aFSE57VjCGzZR28wVOLjLWf
NwGLvBGDOixdRaJphOe5kXAhF9FzoxSG275Zlx5D8zzJNwCXYqh/j21Pfrhpiyzm
1voaPzl2ZyK/Moo8tuXBVcr4lPJE86z5VBw0BYvGTLPe+cRWl73FkVTU9atQ89g5
HfrXLFwfL0M3em+KE+SrU6AaDucC3TWhn9ApfzX0vdN1kBiaUwi4J17jmrf45ztS
Pvorjg3Q5ETgr8326ReXBus6cTvpeIIooNoELue3rvg=
`protect END_PROTECTED
