`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkbNCNItTrIwcNTlMyoCtf9ZotMDjc87N3PS0oT98iX9shfW273jpcLCMez5gQgV
xQipzm46FKPBvdemjAV0gg9Y+j5V8FuS+pwIwjbo8EQH7TJrL0BvMeXJC5/8kFUr
qFi52e+87jHf/KmMDIMdWv3Dl+X3RyoTq58kbBbVrr6FHoqZcdsRYLBN3nwh2KLP
I4AGa0vDOb53+Nv0a0JjHiPCu0yxufMzBNhq8ziGjHVHwAn4/T2TymV2sNdt43Vr
QDoiSDs5W4Gh3cvw3TPa+ZaZPOh2WcvvHHuq9WEwOKbc7Xeep+xVDsizLdRNnKkF
gQfOCSoQR1slLwHiuzvXGVYvszyAnhCANM05jkIV1stqg0G6v+WuMolxUz6V00cK
T68Sp8OQ6Z5KbtBcfqxSgF0WLKYCb4oMQO+Wyx/9avd3oK48asR/fqh2W+CzL61X
/2ZFi/rMt86Xdb0C1PYXGxdsQz06hpZwfOSUOvEaN0hlF22F/SLtllT10UYdqMaS
Q196xPfwhftngd10tzU58vB8CCO+QF7WA9OFY3WZKYk=
`protect END_PROTECTED
