`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5LKvaO3f+pDVv23k4sb08jvjsJHjPMXxaa7FM6esGo9OTcEjP3pQID/kMpcvULRC
veo9C/3ZDR03VlF1H+Koq7yoVipNSDKQMudJfcnPOaaK9s9yzchovqxdXuLf5bv/
21AaVhgujKBVt6VHjSbATqqiSWaXa6woGDhvXr1jFQ/lATajTzRnOpVENTYSh7wU
dreAW9BtnZOtgzB1SXBvTr5QaxdUmIreobWHci3PG/t5heYqrRaDFIoKoaJOHpLv
jwZ+0MiHe6d7fQWYjQbsNo9Ahsaiz4YG88WZFu2Lo42J5id+s812fp+oU6DMmbxV
inw8PE6ks8WCua3XWIc7PmXKyvcZyAqa1fUb7sl7bEqwHOE0Hx6vEfEqpZw16+p8
TovhKtsqK/gh8pvjZ2nstiWQm8N/e7eMgODta1Zy3Ls=
`protect END_PROTECTED
