`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83Gm+tPkScah3rx3TNIJcY9OnuAhvPA5hnEEbbyCo8KzNIUE0GvxRMURuQGEWtDN
3j8cpj2b1rWk8mIzG4tgKQxC3Mw5D1fF/SP4EaRE4h/QFySuLdJYml93RXI9XXUW
yKN6KaZ/6mZnsI4KAuFvBV82TnOVLCGa59xWnUft/pHRkAMMah0xxEBdfT+FsZF0
gn4Ne7F4CrX/zOrPCXgikUmJ/VPXJY+wGpqlh8VJvaukf8JIMCggJlP3sXGCMra1
OO+XHdYJqOGJWyD4BIsDAMRMqT77rz+LJitnU3r2vsyfcnOR7/7TekU4HglVaxhX
juyiH4aWgesqEnOw0C1jt+ZJoQbVB7aM7k/UbK8LQcX7ctSkdE1BRtWDigIOFXdO
oovABezIU436AgMhH88LRlGCUK+a+m3AGR4p8zz2dsuipzYwuOEnnIEKLUtAgnL/
5H6FHfxJbEmjn2xo6URJblwUOEguPFjRutOoKNHUkZSi/auSzuZPjctI26O06fyi
sHMx8l3LncsGZIHYv2H3U0JPEp9JMbrg4zfEdj/V+61NiXB6WJBcD1NUfC7b8IEi
yN10V3h7dkEfw8YXjB8sjg==
`protect END_PROTECTED
