`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mH4OxLKmVI4fxVL44Lx+mEbKr5sd4uvBwntwZ/OHktsr6hnCCuKZKm67bkHDOBC4
VW6R68E9Jma/0IfMIwBM/JU/JfV+ziZpFUGULE7DGXY0j4hZ5i0ZvNvo6sPjPPjS
xNsOA4DFtomgFB2FwvIzFvR/wgH4s89vVHB998eBFkI3fMVg2ZpAec2gIAwGKWy4
mVocPyjgRfBGSdyW/Nvg4hT7CH0vxnWwrUQbg2WXf9QW7/tGbAFAJNjwHjdecyK8
IZsuzR0Ruw+X41WpIVbhcsih5qJYg5mpsF0Yd6PsEzs/3PWarQCqJPs3luweW+CZ
ApzE72eHqrlk5p83Dex0rCw0Q/ptLDXle0BF+XA0s49bLkTwUS/OVj5ZVjUQW186
`protect END_PROTECTED
