`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGvF4YGsgQ5tU/ofWcOd3gIvSgr0oEvVdzk25mT+CVH89Bo3L91tofPlgUxUylUF
YqFNJNorgsu8nyj28NTSWwMRrKpn+SvY3oFUeAXLZxnJCcq75xxXvxT9+g53EACM
lHmfIRJA6T0c3bkkVlH+TF6w3lukMW3/Fwf6weq4ndYb9zuhi7D9KnjGY4nhf7P0
ENgLa3zaILb4O/+dcw71JBbkngMOhg/evZJjZ9SXFPQTWuNDxhVqXEQ8lMYgFuPS
NhQNkgFbEUedaxv3VrQhhEFKw1x8m9TPqL6lWnyOlhH0/FpjuHmAVzLofBMsHU9E
iNdaS0/yXbTNvuBp0tJpBE6osMsAwCyAyaynySwaR3RRsWx6PtosttU62R4Yc45F
9E3M8y7wjDjuzPyMiM1EZ1hZZsNA2IMnkx1WXulbCcXS/QXmKsg+m1cV0Xif5c0I
DVUuzpWAqRiUf/FLKGJVG/iFjSpwffUgSuXGbO/QlqB3H2ZJ4jVotSkIy6GffJwG
DGDAJ3Rhd4whtRjoED56hhOYCKZC32ada3uFy81lXzZeDMS/asVmA9BE0MWdHfRR
6FJFFROPn67Fhiv3+LChbOpxZ/kK0hLXnBUfLSMVseCn0vB6qBJoRuwSoiEF93qc
bvX5ZXDo7XmvPgk9ZVScyaXiaEJVqcDL3g+G0uMXTtWlKO7GWtOQGrfyOF9IM5qe
2kU3F/dPUVx2quHj36y1WRacOJotj5QVXVPxhxyMG35Ly3ulrcyr1C2DEUWRBJ2p
jLeio0LXSPOVHMVgesK4PCfep333SVksIsq+S0H7Ar0melxvtao0G6DkVpVXXL9G
BVg91Ppwq/xT/1wyXaqLJ3OoGefrTPZaMUyxIlFZoMqqvuh6KsLOMdq5l89zCRf2
s1wBru53FUens933w1xCm/At4r0nbC9YXd+HCdBCPTUlRmQxzF7cHyYO3mxQ6Y3Q
`protect END_PROTECTED
