`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dtkF6gjSRBu1HUT3D9xS3V/YxbOaUnmUhPd5zQSGZmXKXAvxK5o0tQZEbqivRvEU
sdUqlThvWVy0aDqQSmuItBK0dbcfl7YUX6CZUJV6EMlB2xIgKfoRec3IOakkS58S
nQui7aNX4+6rwyYvLsZQxyKq4MlC2uiFrKVZF1avKUOYzQ0KC+WwkC1fIN1MG0bk
gvlRf2flgweqcrfWg8SMoVZ8aFuXCMx6I6Yqu03RD+fFu45T1OVwmE16YtxsGEe7
SV5i0GpIopbu667MWgjkDA==
`protect END_PROTECTED
