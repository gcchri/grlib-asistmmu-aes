`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
He+lklwuDZyCZ6pQkTFih7SdCFWqXwZbnHGvM603DVz4eK0nSdjk4URlsOFF+VNV
8gcxTCGzqRmpk24dQqLK8/FjPC/ThE7GbJLMSHTh83SM0sVC1KC9Y5vTkZYbq9Z2
eexrcNAb3g10XQGuUJOX7Cq56aN1fWl6ltTLcLVlmozGji+gAOSO72jb0A0sc8vF
XmRouw5wQ2g7y/9RkpX1wpYJWKsfe8GE2+i2VEpffm5Uo8prvYgX9LCQxARtC0t9
OU6vGeRD7QbPFpllyWOFtpL00cMTZsAgYDiq8sl0t0fs6H4r/7nfS8TmCf2zOWJH
R6qAAkLPSF74nC3BxY2LMF0y7hzXInEC9s8tU/HxgGBlPWxt45IxkEniJejGt/7n
ltMLTS1RxJMZBM3mOUBlUw7ml/3j9zTf9CbLMdTEWG8=
`protect END_PROTECTED
