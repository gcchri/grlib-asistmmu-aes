`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QZxEPXbpO199CNwS8XPhuOx1BpVu9ieFV4ES7N45fmlpQuGGETJusHtBD7w8XJJN
FEd2w2u2ceX5RTQto0sCrm9H50Yz4efcVKU9ctsCpyul7lcwv4E4iWve8Xj7gXti
ZfVbRCJX/Xohn+iSGvkqMB2eNB8TaqdyozuBXx2G5hJwgKZm9MnI/OjDN3nE0KRY
COiIfxBovMs7s9exDAD9XB9pM1HUq/UsYPOM5USJvLX6/vOADNh47aIvjUp/cGLZ
/KE0fXV3vM2iMoveai/11W35kV2/lvt6gRmegADCrCzd2cDSBbeb0c5EXnhO2ln9
YczJikrFwG+25QPQdNAbFyTNQTMl7iGV/Yf0i8M8nhOxfu4p6xbT8aikIlNtntYI
Ld66P3NzR5ro3wrkvBwRHSyC9pcLtUnVhcKLkl10YVhkDhOxlzo4A51pyKYn1cRc
K2qz9Ztf8ks2ClwUHWfWatIXVHhHXo50yUAuo+zxlAFTrnNbm0Clfr7c4Cjf+ckI
wILGYEuNH0hm57aKRD4PZTOyZ0Cv1PirL+dJbrTV7okI2k+UdlJW61J+6IJ+CZjM
uHqGwNN+AJorjzzkeNFcKJJL2cHuT7pIz/g2AG9148bpfDz0Di2D4TPrlycHP3wJ
E24n1dRL2lKauITbRBlkV7jKm1Axm0WXo4ohDjQAizqYmM02LOWF02HTKsqnB6T4
`protect END_PROTECTED
