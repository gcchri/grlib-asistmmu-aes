`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+nV+uoJjWZzQ88JQ6WLYOGPIn1Jm45RjHwYUiPS769siLutDWaVZ7JJuynV6F7U
D1Ug3o6o0zK/VjP6QOimFxcNBWuj5NpH7goJT963aUSywDAS8Qgu/QKjsVwh18oq
SV6jTESaeZYkl15x4vKkIosKeCXgShiKIBkvr8ZW0A2Ns3B9qOW0KzwdyoQsz+E2
qnT7LnoGbka4A2gx9zACXW2HPmhpBSsT9IDk0fX+vl2SFs/8kqY/e9XMKyO+6eBI
u2b7cK9dL8AsrWvtO7bOCIhRqAufa6N/wOw0Ni+zCPlravpo/gtf8RvXmLofiBBx
HQeYSuxNu6KyhblvXcI2rQ==
`protect END_PROTECTED
