`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aAPlfc5lN1vPXUUCEHyK2xucNt8OKqYEPsDDXzxdSBQyk7EmEwLvyNm0V4LI0bxV
AZ5DOiyux9PmY/C6FCERaACUldulSlZ+kn71oUDfTClzgwTa+lMg0OBb7zJBVppe
Tr+0y19IBkCEilWu2hU6af0wf0U4Cr4yQKljgyxIF8XBXcz1rxUpo2x/9kaZAg8B
UGgvKAErw9SrxfOZpF5SN3Hq76q94hA99/DyRQc/8CG/phMc01j/OTnLbdIc1cvr
ta39cJC+s/WpITovOzJB2GmMjYCby404gJa01fQ+snIbFhuTUdf7bLaNIUvVp3KB
7Vneqsvw0oYSlywEeN1XjR6P9G5/ZR+BgQvCwgduFSc=
`protect END_PROTECTED
