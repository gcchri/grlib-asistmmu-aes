`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DZyxtTsn6rxF6zOAlb7ZUwyVooUPQSuBl73o/imlQrmHX6D/zHmsoMQGLcR9vkCK
Jv9K5YmwmetiJK9pBtRswPMwJSCewrvRMcINaBkyB2CZJgVUqpd/fanf8cPHKk+P
dD54nSboF/xj9+C2ZmhZzpfLS6ufdTS2QjLtzSoJU/Ch9qY6xcXhKMJughSECfuS
qWup6Zv0bTjXuLZlr7Jy7DJ5fa7d7OmS1S668LiJZeVMp8DTKEOGtPEXceuqq9q6
9V7CqLMTpBvc1/Uvu+nekQ==
`protect END_PROTECTED
