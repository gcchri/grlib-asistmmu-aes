`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZeWi8zV2tb/f4FmqJ13pyRRm+nTPwpdUu/hDIxzjFneUVD+KTKBvOGZ0G01WFnPz
X6vxp6GOkWXc9vJ2GbOz1te7P1RDw5kidIKGa788DKrGHSXSfj6uAaXwjjrRvVpV
z/lOaqMAAm8ftdwGKXTtHDh7ocxj/tBWAoZOtEXAH4yFLFE72VrDzRqXftcoA1vz
h+wsE3IkHzRtdlakfV2gZN+vgE7LD9AtUIuchu6dO/gyFEZYPqXNTTOlO31G+Sss
j4c/5v83hkoVUuUlQwdPWR7YXxWAx7EoTs+ZBPJGsNg94twd7xZAGQCotQ9zcmz+
NEaeq+NyK21ZhI/kvnWnfT8cDBSACFHLQ6qZ1oEjYjdhFcJ6k+FbdFMwZhnT9Jwc
/hwlsnbgt2KSPgDifik/0kA7p3nMNB5fC+hVNZMrWHjoJlickbzO3+oHxaqv1E4L
BJyRUQmDz7Akes/mbQ/nb1s4IPVwo6KGFU86enUKBP+jAomar1EyR7QxQEcfASjr
ta6h1Tps2HYdp5Y/xMkxQ+3c1iB34xLf9OIFdvAFWfVpb2Zs9Vdev+P0RcRwN185
5xpZzPHyUG9fm+s0O6m3b+3hhRrf0HjulcaellChgTn1FCN9fMES8B6/lFWh2yye
GZ9As2MF4EF+oogU2Z1koGb0mp0ysfKXRFnl2RVTUrKAc81f72Mkgg84r2PFfoSL
hrwc5aM4lsGKoFxR2apkHiW5BdBSr4X/q+jpjY5B5FuO3VttPkER4hbBhy2Y5irF
KXIUAi4PGvftsHkfC3tBW5kEakU+NzDRwWILlPbD4d+rrR1/ewnZDPMAPHC3EDTX
a3GIEn3PqtvghjKn+m8RPx+f1I1Aqoj2jWiCgmvH7zA5RSj8vVIfWlgcYsSHS47N
VrEUMD9b1fIiu7/v08Mf8cXAYgMU0CyALrjSq7RPmprTuRPbw9G2qpv0532eMlF+
FdrDDOG5Oj91xPQ5yIWFKPtuzeA+hN6eqzUtuGhfnk94hposit8OftFjAXVxWeIz
Yd22UWV4evNggOH4L2FdOeVghme7tHJJF2N2agZjvJrVQZZmZfnN95V3LxRlfg3d
jtC3sB6aiczL8f8jWXmdeiAIi1FOwgVmdi8oGk1TElyqvzG0rPtSwH/I3agMC45b
k8rQCHm2uXxeqLzDT+wShVkoIovH/fHgV5iilswh1rUJUIICKZQbi9YdO4UdKWZZ
jKt8Y17yFwHyx7pYr241YpMsSw7nW+DoR023ml0BSTGbeo1k4yhVrK/P8krV9qPY
KclJCVHoq+z3T0qWeCKQx5vItQTIpI/lFwIKUdy1k3a5Jwv23e7+R7zqgBSlZZZs
Iw6qx89lP9PeNgdPyfRaoTK4mIUM7xNlSoup7KkMdGqY1Ak7z9i3SL9/XGJdoCW9
vs6RZ+ppWHgfD+GJgGANdJff/s8/jGG2ZC2n/Lz+zENN3vjq8LtBt+VRYR7z15IC
OiHzSqkcLjKTkWSUnuKWQAlaqEYCcnKes7V8zHf7AllNA6vjEvIJwoWelA9zXuMs
VhjLTUINqB7/PVrMnH6Iigegby/mfDQefkv77CsqcyjBtCa9DwU5IRr2f4SJC2Ng
1StYrtni7Fcrh8Ttuz9wa3jqKvAu1ak6Jm9KM38+BNxZY6goT7TCPAryRdTcSba3
qwV6rSyxT4dk2vSscFDNxltJxvfdsjZ3h5Pl/i99N2SxeHR9Yrt14+gD2302E3Xw
6W5Cf8dBnjKHZ2p1Ct1qkYFCOtF5Yd02FBbQZPWy/YiACUg8ed+YcfAlxmBkYdt0
vU8kTKOc3dYjrATBdgo+vfiSvsfojgo1JQy1REriyxSZTc65aN92KXMs2PaaDXIN
vX7K+V1piRUTbWnb/mycj+NWWPh2VIaEpWIygFwSw0mWXxC7hu1xgSLNhdUOa3Tn
WJLoXNWwOQnmzoePWyUaDR79i0EoBqsp9oMuZ4Lb3OikLN4htta65XfNYVdQhw7v
tNq1kct0zNHNpchpzzAdOGKTA3JRbwEKFgxWqk6xPkOcPcC7mZKl+l+NIOnuwnLd
cSKOj+armAqAqLupQJQqwJ2ILCu+wUjDIiSlu3d+htQrTHv+Md7RBZYDX31E4Bhs
1mLua7eMfIkgE1KgTNKF8wCkfyYfxKN9g7FI9aT8Dl2q0yfxF4xxNI6ineou5SHx
WWS2g56lYZnt3Jilo8rCMNabikxpmW+xInbT9D+A0IZePs/0/kTHYtEPJMFzox4T
70/6uaElzvaluGm67HzgDKhQ0vhEsq7MW7FB69wnRVElXeujgzDsD0qPw3o/Nl/I
z83FShBFfeoVHV+1AtQ0zo4UPDYu/stkiuDpaW+cbDlf/jK1H/8lWULXh7jL9xgw
H9qylA3qRLSVJi3EF2Hj2kE4feSnopFQH02YdiGqhQokl7sk1TwbzKf41EkvUzHW
z9gVB5C+R7uhnZia4mMefex9lP/DlNx4LdY3XyK3TAh+N5wISrmwZN9X1aHkrx6B
aCX/goNhXZMo+Ru88p30PpAmYOXGYaFtBDMDzB6FneeMVJWh3dbB5dATS+54TiSc
Em5rVcfSZjRNrno6SGsbtZ6EbuiCAoU+iF0jf+mW5oxwPPr3FzmikBGDjtPCM3vS
S/VFvn4/xvZsk39yXj0JJU7a0CVSLUmo3q3moUZj5zukDoFkhPqECDHdG4GtWh3S
ds480TVx1EdS85FqHl4z16XVxjCK4nEuXYUwEUNhhLQ59s25S5ToOm1jvsxnCuLB
KObACVZuEg8PJCr2YC/3Zsu1gR8nByLuYWvDaJKyIElNgV6hb1WT7Boeme8ztr7B
IJYQvMV72DqPElEEp9IGOnbibyziv9+9E+QC1XY4LiJ9ddVtMpjxpY69lFJULGYK
yv3URbks2qzF07B8gYsgesMUtMZBL/MBMDh/2RWElINcwfIa8f/YBohCjlhMZFT7
7Wj9W/zZPN1zbKndt0wmBsIolAYprS5/ZG5oiYUOXlgAKofdPNm8jD6IfFlMEtOk
Omq7bW8CLcpuXWNAnVmsMxlrRxFDRCxZyYAaOlOtrhZWJisKR/a/Gv38K/ivQ5w3
Z5D5BNEjkXrzlklIcHBHtyY90m9CpDCa70KjXEEe3bVegAmctmpI/IVeZNYAjOke
2ctp0kTaRatrKMj5A1mkr9ARzUpLk6/qNnB8El3ob9PN2yAfvMWYrmjyFc7KBGHh
sJXFo9Vk7jMyO4tiZRr1z7GU55lqlpYAQ4aNikw7Fg/kz3FnHOS1NkIo2CelFo6s
uSiwnbqlWP4tzN1gYSNtXAeQ4wLudWeaTNmkrsNxad9bpr9vPGpeRFLWLGX0A553
YQp1OgJTN6B/9XkWoUKTpilYPGKYJOUiJObB9qoyrZCP9apiIJ9ab8T07mVkVT8R
LBlfRVvQOUi3xmAf5EtjwzjSevyeIZbG6AZibOg5KvtyHNPU40RYB/CsFgnDU+f2
JgGCNUA0c8yTYoCQfIr3J6n86KWjmTfHEcHH/7kLjLgowGKPGoJNj6R2KHec0TRN
btHIrSUz5jcb+0Uvg3wYseYdPAnENpFrmpQsOxc24nsRUb3XO122Plsf/LEXaABG
jgbrAAWJW7kQyeFGpcZZt8e90O/F9LV5R5VZL7B/zrblfPxB9HcLt8zUB2XwyJ0G
3lJiZ7NN9uv9+u4ERqO8QcWXUrQlz5NKnZUnZaAd6V7k4DX89WZf9q38bvj5BGD6
8VLG+/o6kPUIRA8kX16jEfx8gIfP/qw19Lwvba2C5MC2KvplIXuMdOWkehpfuRg5
SmHphf6V0a+JcW49VIC4iPl1PeSVvNBziAAeuaVcd7tth0ZddSPPOQy+AJ1D7rag
PKQnphWje6cxygEQo97fLQnpbzdUuYudZUoiNbvpyfW24lkKjNOrFxwvDpnV0lLn
EhAQovXAHZ9FjLwwaNBRQkmbyv6+GZc4IpY2/ODRktl4midQoqkWDnKT12InqztN
IkVN20I4wXoR9RXhuuAkKqfo/mFNPua2dyZJtRoYGUTYDHaLX9duWhAoY/QyRzqf
91TamYe1qCY5QSz5tL1AoyBkaMIJgaHlxqIYPX69gxQr07zdLQNjnXnp+E5lEJm9
v/PP7xGUjvMqSMFxM/kwaNZnvTYGey5tpbGLrVjDy1d5BFU2+BwJW2W0bszHBY+6
kDMiIpqwf13Hl2wh47/NOm4tq0lyTuH7jPRovuQLRwb1pBIpxEx6TQQVO+q18c3p
UX5yS7Xx5vjZqfakK3qmPTqv8pcyNxKbV0cLjrysrKtd/jvKHr2iNDrO4vWruPGA
z9rKxhka7ZzR3pv52Vo73pSdDIJaQvbTlM2cVI67niez/GJ6oMFm66O/Eeo3JSiA
Gl06gmXCjXTYOVUZlWN6udCBEsNzsPSsf8tH/foME2tPb9gVF2c8Tfy5oWzMfJby
teKRL28GyprqQ4EnEU6WfIwceJSLgQJJ5rLQ9/jv7brCsl1kG82olaxg1uG1u9Ff
u0B2DXsKg3Pv5rrdgKBN9Fi22LM9Ge409RXNTHPaYrOeV9Oiv6ZngR77EoAyB6OE
/EK65/h+24J894q7KSL+iMxsMmk1YmlB7CxJUslkVb6k8QuHjSynFTr3foTfvikW
YU+I0xmCTSoFAqcq18+xWifAfzUeFngSPY8ofwkhj3w4v8+reRXHzDQVu0Nifejt
Ao1bShrRINvguxmS/eu3ElIPpwrXTKm37migggQHSXYp3Vs5+IWw68oYMaUzL62A
nu2L0a3YuSsW1HyXZ4wCQWeOIFCgPQxQJT93MlxDvA5KbJhnMoBZfxY1hKApj1Du
wMzGNrx5EC7SG5mpdIHbiYiJh2771/7ns1zvZNZrjzqdOjnJLendKpw2ZM8AR6MH
IBAon3yBLm0MPWNk5acUP+yqxtS8IdGYZDLKvn9IQZk9S/5mRigmDCdG/ftA0++Z
AtWiiPmjLbntGOwCsxjDG2Bxj5PtNjt/AeNKah0IKWEE7ht1cFsUhO0IsWhH89gI
ZtEw862Hw+byiLQst+Si17+dMG5akJ2O6YX2iMz7zIt6ZvzpEV9LgeRTb7txRcux
VNt/o//vu+AN0s1curloF+THlJdcErY/mDTnsAPislRWOkGpZlR+YC9gB2T7G/LB
IeI6lJYmt3FmWWtfDFvgyglXkwMjktLJ7osZwW+pEZstSeP+Nn3N8uTj1ANe4e7Z
9PbZSuhheqMXLuh/5LCoj0fMtbGueJ9ZflNXJY6+lDNtzS9tRqWgY7zOwoTEX5W3
kELe2TNnAKT8VohtkxcAGwcIneW5FCDfqm63rFcObUG5yJcmboicJxGanJTU9kU3
SB5PoCRd+D31nK9JUtsOJYvvDsMU4nmTC+LUhV37cFstZLrtmIxFToLRGzNlFsr1
JKEsbNF5cknyEZuqb0v1EvWC1UFEWZjf17pQeY5HGlFzXPzM3rShn8yezeAgyW8U
Mpi9qAqeC0RNjRqlkJSL/MIwhKeHuNhW5y7AEj7KTW+nd+tRGx1cuCCC0n8/pyhF
vey4mgry5Qdzwv/ZVnf4RTuRCzQtuhzeaLBX0W7+WfZ2HXlnHFgd65vdRKKkVClb
0cx6p8Gc1W6z5My7mS7J7gwaJg41pGVTabz7cwnyxYf9t8tiWH/7U089nCg6etWr
vtQ93Y+Qxu4HFviUVLn6PP82DuY+CRsrYqK3/wOBHn7f+HgKVQ+HyE835xUXtf4I
AY22a8TAK258gSBAbT/hJyimCiENZsg1nY4/roOfCsySLsGa9a3cNxSB5tY6CluH
lqLiMJEMU9VJTg4P6g5nqeYCk/y4tBLx24oVrXNwozCju5Qy+JxD5DLf2C4u0BMr
o52ihXe4T/4SWKvpxmY8SHKu28yFT8MJXDlKTIOA7Ifz9KtTxG10nt9Ft/MTyXJr
yxJcSeEqG0IsHhdt8ctaEQTsCQcdnMwy8sGjJ+ke1X3qDEZr3Lt/qVNDw7iH8Jao
8F3p/ZtxjtfK7NXlOgU4EOvKeYc/d9jDYgJUcECLs9gwr2Tc31ztXDAPjF67H6Qp
rFXzDlYHMBkUWONJAtbqc0wcKaBF/V86cN8JXSJnEVcr5LCQDs5y70dZRZm6AGFX
jkqJMGHVAKvL8/goJRUBQlqBKWzjv/1dld6rtl6ER6WnzquJWnd6vauu9Vm4Acqk
0TgzW0RWC+Kt987qi9FyfZgaesf/Dz4qFht1GdH2MjkIQ3fJsnn5w2FpwaDz+VMF
5MD56cw6P89v3OegCF+HqWC/0anvO/mcwL+lih3jZtklbScGC6qaKW2UoAbaCDeK
vsz2LzzmxIuBbNYWWEwIevFB7idBhCiaTPjPCDp8rCQKg6Amdk5VR9GsQc4ZLLFy
e8yJ2d+MzJMtxy+IAwEjNBy17Y18zPZxvsBfRBD0oqz9Z3e8RZX8Mj1DnJ9ay9AG
O12VZsIUFicMmVTNGKvYvi5GusohErPiMnNu0P04x05vNTVRJfIQNGF49Z+GC2iT
JMC59dU3O7xBgnfihWMkHiUh46CqIoYeK2+n1j99YouQzmj0HPivEHIzt5bzTNGQ
O02QBt5nYdiCew6/4FY96esCh/B1JFzGF56KZ/+AkXJNe4kVgh/YURdNkj5Xw4I+
11IflwccqX3Qs2m9xfY6X83amlNt8xIWMIC0pOObvoRIwcIkTGT/ZM7t14o0HHP2
TfuqunAmxhLsAmIdsnBLWOHXwV9Cyttp1e0PMax/jjqCa7hDpR3UfgAomOF1je71
GHrE2UEvIl/NHXuV0A1CEOqXnNC0CGZTtKIRlGc47zeiE9H2PPn9itwCefwncZQC
xvt0mARRGEZ3npGG6AVbeuY44BRSJtUrNxHMXvCpVGdWQWqGjRVRumbr5xkkq/eE
6yHgU6toJyL43x/vIoxaDCPjtiqyoJQMyk0tYMa2k6BWDwOvAcfECXkdr/AuDyL8
ZICXRnL1QU0iyuZCwsCk79+Lr8w3scyWEmMuPVYRstxeBdv2sKqC7OEDAn8tf1e7
ZLTmVWVddc1Hm+bKpT3eAplH8h92GQNoJtXtEjfYeHeplDfn4AIUI50g0JuNC2/3
gnmwkuEcdx9jh1ufmQ8UVBM18exdfPuNPm29rPOnEVeGBndymdPd5MhJpOenvH3l
5NY2qNXeLkUPPxD9Rhc7BsqTK7QWlm9NCLqCsBf/IgGwIdgjNUCMEADgg3IKO/a9
IcDZOyUyqV+pnRtraZGGXRzCMTvMmxoJNhzdtrW1mIKIRUBXKYNeQddLapkqIbPq
tfPd/GzlObQsqMS3gEOPxuIGZCjhfjHMjZ1CouW51ftGDW/PjZvWKnA8q6IFDBLq
GQ66VN2DivleFQuqY/6FSHddUYV0OsGkvmdIhCRWgUHfLqdcciODv/PoQmvLD9yH
Okwq0wF+BUY8j96MRN6ywI/Z21ljB+GFCuPbcGmOSIJw62DpJCzSaluV/tTfTFKM
vosHj3v9t9jztCT1T7r9N8RTI/dWA++m36XLonxVZsrCyIMsHMx60iiLa1sEoBOn
/qnZxH9rCCoRWbnNzyAGPg/bjqdBJdNIEg1I0vdtlM8LR5BLYvScbtSJrWueTTY9
1T2dhIrX6jhVyU9NTMShzZRfwH5wYOppiJ0dp8P+Zf6PWKDxZbXAtF0IP7G9bFnO
0ctfCn0uGsnSksoewBaEcoOyxJ7nypu0XlutLPfzs4Y2ybMq9xcZ+cFHJWT055Py
bPLq027F20YlpvvqsoylLDcUnm+hbPDkpEUAXlqb1caJbkVY8IOo5XspgaQbW6yS
Kd7+Tq+Rr9OmvY1D/yan+MNMwVeQBXCPxiibdRMwpVLTMDp8ZFOz++Gb8cIsKjtu
KfS1RFbgos0gDl6dJbkG5wU83wiC2GtVnJCvhAHzkMD7r+U/JUXvtkO78vYxALNT
a5TB53R55u3QnEndD1WHYA9DPZOngjV8Z7KvVxyrhwm6WckbcZGwnpritxXYcxTf
Mr13tFexe7C93bsdXngzUNtf2Kko4FMgSONWJdEtTGiWusKsP/gjkdc/ZfqTQr97
o1t6eFN11s99ELdlw2reG0FvXanfyQOEHyOYUqQbxX5sXRY8no6BqEOSg6LFT6cw
2Zsavu3ZKebV+0W5Bpu9iHSkbnyWRg1DL/KZM5m4iG9iVouNXzVSGnOKEdYyUywN
Hq47bGE1u6UQXCYd2WmkzfvycBZKxt6Mz49SZDX/vv8Q7v123SLJoLAa7VEQFYh4
UBBZZteG2xSwaUp4mR6De7LLxqfTQSs9FZqmoXYnVSM8pGR4hQZL1ZbIHcO38i3O
T3cL7eKZKV4gAVtAw++oL2F1h3YxGBcS2yIYnxpx2OM+wtw5DIVk37+hwrjnC6P3
fiPVzorPSVZAICwPiTMsBJPH1N6ONYd2H3uR2GavLuh/97YFG4lnpxsUT9AcxfHm
ySFVr4ytIWcCEa595qOZBDAYDlizQQan6lGvQLngCvWGzH9olMheFubOf5bDCrQX
5Ch7iow+WH61ebTIjcxCftYNIiJlBPhxNZOoqoD+YgMBnUXokfn4r28wkdftFzqA
kvbdMV6tBMrHGVZGppPbxByHjzdd4+eMaYn59FcgVSt/0O9DH1rD0a7twNElSowf
mZEecBowVV/VN4lN3DCUKPZey3NCibmZGEkGtAC6dx4qZ3pwPHDVG2QhQt4hALft
+sANayxYv/vmz3s/rUeE9pk8tLE7KtY8MWw3m3nOzEhk+6kg765E0ZbxYA7zJVT4
lWFcj33Mpm6hlb0D2U9i/aJhArVPZ2rn0t2P7GrfUeJrQ7Ce5eV0vFNrUaU6J5RQ
Tpj39XAuUuBMjo37ijSqMFobC5/KxD7t54+IUP3k/Xt/TWGzQ5By+PGpiGnrsy+/
QBx+TSpvKe5lI8SBB+NXo2592U7ZT6EoDrhFjvubej8YZdt/BsnSBW5+Tu4lbO+p
7eo2EghFLB8ZDSqYwcrJtEYTr+2EIwC/1p+Y1ETTm4L58vjVT/kv3XjG8Q9PUSro
Ew1HE8Ef8+VRocb+smdzsufptjO81Xmuk9TU+5t2EQ+GXfxILDlrYyub/w6WTeJT
Bzd/3vyPWaeFYHAV2od+KKLdgEZm9P5TOhyoYGtMjj/g+pK9GnH46L5hvISlYlQA
KOJojvF9m4gtDahG3tbZrLtaZHTkxsIhJNmZIsLvgg7n9R+1DE7lwwZ7rm1p5slA
T4lSZ6UNhVVrP5h2mukuzXVJ0SuRRJ2TTABTxWgjb8AMcBoyD87V+qe4LQOBeyor
WwfuSLBixISmgP7N/4HwunOkfAhpnxkZhTg+2wqb1xtylebWltZo5/TGYkZ2uNL9
RO0hsHR8j86BabdzW24IHryVTNgcrvW+M6ujS/J7L5LH0evI2rHsAqoRcYm7synu
TgqnzoDcdrwvW8mW1ntB+YzTdVIvLUJ4A+Zb2gbRUzTQMXNzajVla+9qg3a3jqMk
+9XfJPm0dH+fd0Sf0D7VmjKmuz2dMXlJ/nEI0iD8pSNB3pFzaUU29LPkCnc+B7u7
dy84IWDwbNOkdxEcSdM7O7Vxpwym9zZHo9iPGxnJFsgi5sjdQX09EzTki78r8HuU
Dl7Uu5XZvmbED0T55o93QXRi+Te2V3hQewHjI8pm4dMjJ0AeSqU2Ll2dfF/Yj/Lv
wz13lHMIyC53e1OqXL0CAa4/Rg8kFYfJz0difFT0wjrgwMF9TgnZlhKsMaUR54gB
/2RamOe0E7Nsya8yV6uuE0QIGzP0zgCPSLcBukP7O3cCBNCwYLfuUB4+RK//+10n
EQrF/0xbEw0RGtARhY301YxMSbEatvC0W19KUBFW4axGwxY89V2ykJX4CIAxs15K
zVDseNsEbPtvAWVQXCaskU9gAJ7MQswHTyMY1PVzix1tQy3+Bs5bHWD6jKr2f/Mc
i1L290w6/hHV4K6mSlRVtfPTnO8kr4pz4hgXwsy9kDTPZWgmzCICMrQCsTO9qyOf
JjDNf5ww0KsyiRGJCNZYbHPm0uSPgtEyBzEtyI1MQUlP6lRCscTWe8inUeGEY7wV
GkfDnaZWrgTKdWrnwkiS6UOqfDr/iwXlqA1iWBzVPvgBocDcIITEdo7MfOE11OtW
gwmKL77q23DP7P9uYiQrn5bz4UFrb1geYQEs7NlCz51nxqGKmjkkPptILOozESe1
EYGQtfe5QPkK0vYr2KAE7RqE68kN5OGYvztzQcDZD399hQ5Ftf3ce3eL9ExXQLut
1iANI1Rra/6OEBLD720sMTkHw7sCI9V0kcWVcw/D5vEGyPxwEgAR5KVoigKOlG2I
uTCLSYbyHstpuvhREPCZq+bGDU6g+PY0MgWCqXhb7Bb6T8MZcgGkYgdiTMrV+rgH
pjhkV9y7BmhOHk0XnuAMsR4Pz+KbBFKMuYk9EvmVHqTOxbycA8s/kNLAAulXRvP/
wid427qEo1fLiT8afNbrhADjNRrRWWFiGmqxHyyAe2z2dss5PdA6myYJsXAv2jc8
SLt86nStMoOYf9GFeewiPYu+r0pbaY9pKTF5pi+xSlM65lwQ7HwT7bqEBELNiug3
cOrumfV/J/N0OE/mEZ9n2/8wsY1ZxBdEjldpFpHYNJjiXNA7vjGyzhMqxiF+Z9eD
6mKTnH6qJ95rlIZhLA0Z/ahbD6KEzsD48NWBVzyNsZRLnWM7RDYijKqrH3L4I9Ri
Syb98S2Km8+LFUfeaZqLOS/BA2k1NnRCazYsn7wRhFTOfiQ6xnH02EOHY8Ijodyz
8WPM6ROyhzAO9QlKCITTDRznB+lLgO/vvSbPpmgcciHnA+Vx1Ly6sLvhke9bnp8P
GrWuQkAmjEY8uDDVjv+hc6XQ8wL3pVwgfheb+HweNkhMwOdspIyAfyQOCeiCGxpp
z42Qvn2KB9L0NbNCzT7bQt9mnKELqI1dteU2ui1O4DvzXPeoKxYnHlibTpH0Gy/X
64vbbk05W8nnxoRrLveoJdkSLQiU3PRsHcE5ykxcqJGqBuGf+imbugZJfRBq9qGl
7STdlhotaZGC06mw24zQ/oV1M6+EmrsV1l2pqIWmPJyoelVSBWX9WFgefgkVRN2g
JfU5BXJPVr0Pk92rcq/a/PkxLcqeT6QQyAzO+IZCFLGhhrCIvWzn18ArGnw4VbqT
LZHKLYdRbyFvp6oI3PxWKf2VVt5aeVy0Us+v+erM3Uodj3AiO2nm8yUP6Qj9aACh
fqG/C87g3z0tSvWpStByF/m6jPX7Bkez5X7o9B24VkyzO5RBnwiyalA98W0wsUNK
eSGtSRPPI8X+JcGVbs/XfTgdZvdweKCgoisdsDVSUAZVc1tq8m3TG36EGC8Q/hty
NpNApjvcCIUVHOWcZU1H+jqkgPuGN4lAGRiUv1DZi4o/4yppH2me909fhrRmrERV
ZGc1V1JYHkfImI+XFq3ZrPK4bPoTzPNBJrudQCQEc0Nopid+0EO/bZT4nrH5PahW
OFw5xU+iVJOStbCfPYHUL9dKryglUwgcW6N8VN0sJHZKhi7tuxbbhxSpsONJj11C
omsJrlaHYSL8NAlbdFfeSaZy6ngs8pzYFid6T+ULE+xZXlnZZCzvi5WJwCzlBmoH
5soVqOd/uef0o4f5qDhZBl5FKS+E+GtRrgqf8SAckBK3TV4Sgx79Uu6ZwdwJ7vDc
9D7LQstW3JoIKlPf/9d7W73kDzGllU+CkO34tKNrNwX6BQrEI/XH90rBRQbFIdd0
FUOajWX/FonM3XQBou9lt+ugiw/fitxmJQmt7nsqbJosWEDwq6iDUkcv9eUBNOxc
zsFg/ShcorEUaF/6gbDxPMNkwk4qaUb/qurVRTLVbnYU8ZZwOLlhmiXGmneBg0X1
cag7f8F+TjTTGLp70OquvPNCG6qSefFs4aDakt2/l/IF/HktxlJ5LzhtxQMDCuBM
TDovepHM87GlI5+PXAOala+C8kFj1x/s+HC2v2VTZ8vMiaj40cDbRJ7BqAwEm8mA
4JexJQZSZY7/9WkhhC2m5ojWTOKXt8icHuhhAEk0YVgPi2QRIaAzcTdM0gUKFUbj
yDi5Uh/n9WkPJYRvSJJRCccLMlM7t997lDE5MSiQZEVo3gL4bPUJqOby3nTSGVvi
RjiRv/TNRfnXtvJ+2wqGBYjyOTTa5DXVQfIIiP/1T3YVeU4sQ0/vSb4i/XIYZ3MI
lIqqD42kK3wLWC+OJbmQI97a2d9mqzQVm8pFYSJ53J6MudRK3RP5GUtGAQzs/+HC
1mb0UgNCyKxYm3bg3ll6pjQvVtZ6g10AGr4XlTpL9AdGlD9r29grpca5vCnJBJIg
CABCh/FeGR58CA/Rb+YWLewSZclUGNjeFlE5u91657O/obBWxl0jmVCMSSNOX1Mu
w/0jmsXd4BgRCwoqBH0rB9hmBdGMrPQSsx7JywwREDXfV2fn8lS+bYi3p3AcwGA3
jwbTvdb/l+GTL1g7WAinTL+XWB3Qn5TxAha4VfJBzVKHY67gwWIneuzl/49rzhAe
qyq85jLJfN9PF5U+bTCpAai/bLX+aiiz0EbtyNGQCS1dkJGB6lBsCE6pCro/MEie
zQlMUX305xDVAv36VsCTw6wEpwEhMlJ0FqAictqF6BEP1wPpqspI9VIZKkYzE4Uy
5NZ9dpDRR874W1PgPMdVVZ3kIEr9wABM3URNjpINLJv0un32CdUZ5OxMnqginRJ9
MgCnU7lC4612jIiPBaqSMrUstV+y33AD4AUrKX8hHZgyUDoQDIVH7MYlYbKwydNw
vusYMJLPVKZz7BlpFTRP7UyvIW8/TpHYe6UOEH0jdXDJXqfmv/Pb0q2j/L1/bBvl
VjkxkBUz4ATWn8VSAyTGU1HXZmTqTFJVxMJocwW0R8lEHqrJvd7FrjXqUoY/9BG0
pGFDVCJIE0tqR+SHmFu8k8X0GqEpN3Vn/VBU7rQZdDGfhMucuo8WubYxuF6iDwX7
e0/oMnv2yWIG+T/mp6pP9qJtYf6x6dyjWiVwDFjYpBStfUfQ9sCGBZQmE/IMSIwV
6DAe4Fp8Nb2c0yHCr9YUdTXXafl/U0S52Dgob6ko0zwK63zePOajhlrtxUwVyV8a
wcW+W4/hueQkO5pSDN7EoUSC+lvy7xLRH2n/cgSyQ9rip845av54PFOoZR4TMRAX
zXO/GiBsDy4r91So0twy8/AT7sDvcDK13jb0z/GODsetRCMXHMGgDcyD6oTU1xA6
IAPPbMCORyM2NomqQ0/BiR0zzmUqHFeC3h33lFrMlllS8RjhuIVjgHIWehLGcxPl
JyieHuJPAHQ9BEereQ/y3DXPiypYQCaGIIbYHrxgwgSErONZGCH+CnU9wV12Vl5S
1x1PUNEnQoikbektvqDB8q89vTeIWGsMyIV4E86upZN2v/tmxHRatUnzebH8qnzF
/7nCkvllZDBMjAFBhN5Kl0AAlek27tCnRwhCUmPWS7RaUlpTva32KSsmx0ucPz0g
zCrCt42CxM60o286C9DGaZ+a3fuvshRLPKQFoeY+St/qVfS+UFYyEPWDqVnKGxzp
PNK9kDZA7qo9101TewXtQc4A0H6TDyGxZDshh11/0LLyDz2XRvFe9eXmaQk626o4
RQ/kQ9Yh6a65YkjyUQlo3dl8nXkId5Oh4dHnZccWzvMzigUigzwZKxoYjnKixjXL
RjVoWfoIO9Dj6Nolp2ZMoL6MyMAcKKs6Yv64ybvhZEmnbdG2rAdjNyLoYj1cUEb4
S6J/MMyDSFUV2cmU8WSsQ9qwJnacTK/MyZW3gmaBsQMvae66UljaU28W/u7bA1jr
5wGGtK+BG1Y454L3ocrUzwm4WFRD2u8YdO+ovO/1Fb0OdmqFaHDBWy1dBzyQSZKy
YgaHod+Bk5HW3TqBhMYpTrIbmIdHvKmN3OqlqiDr1cBWOwqIJHopEYJXvJaOwpSd
9fR+OYMkndtIrqXPL7SGn/ZFpYn3ekw+xOpywjp02jpy0Vj4XwNQbsjGrMA7ugrf
ZeYq+rnudI0seA9Tniw3t98y4Bzjz8nl50NIlnRSvxnYn49ZJVTfxtKTMvyoPcWL
8i0UN8o8vluLrmlSpYxDx1lg3eDrk/EO8oJLiAroRKOEMzPKsT2unth1Yv5L9TUB
fogxs7rHnjNIhX8gHsUNIaFRdJB26hguY8ydkWy18zjHbQdqDZ9RonK0XNv3MfwO
esjhP90MKbj2nQRRzP9J8aCQ4Uo4KeQHvV3bIBVtkBgIsRY5r9mSWmdVTpNo8yCj
k3FceCuhjbDSam3Pv9kAEmt9+uxjA/FxX1ukAWIls+dJuqQ9dcKdau2l1XsrCF3L
DPPpz96zwzkOwMIqZLr4v7sK9/5t8YMkUNv0HCV03+W1p1KLCKpukkjq6lYfsKa0
k+P1y257tl8Y7qWa1t3wZi/hiyaDV3ff3tYhHIGeMOaWT9kDum+Ob8G2SI6NKC+E
KpannQ4qCg+sXyraMpuqzRwPfW7LA2NsuLYWFqBJORNHnukRF6gYheYNrgIEqkIe
K3k35ZzruQkvBTnCo0DG5ZnMLZTZjy4HLHEhKAEzFROfGIig+0Xlw7dU+N+h6giF
vjpOc/DCdxxND1kjWwB322Gp6CRR4GMHq7ZPnJeyJSaBkhubnUk4P1F1EB7D/2OY
6HAa/NI1EvZDl9pOVAO+EWdYSeHHoWSuRF/sRxss9VayCVNuqguny9uPOcvfOXIJ
nsyWw0JqOR8ytVAUoqqmK+L7+CyFkRPHvBRQpItcxt5QRLKdXwApA5EQluaReDxb
nDeLr+Bxn6ZiPCpymCJMWvAhekjh2H5SM3EvkCn/u+n1fvJL6QetJghRRH1yoi01
zsZUX2yleMHeCiD5gqIxsSdFkGUk8hpOec1nV+iFZcsqYaWWvmR/M9gssRmJk3Wf
zKbrM16JZ9HFQLBadfDMBcEE55+9VcEioKJZYif3lvcnjft/U01RCWLy4eXbxX2S
CBhYUKsLm2Qh1uth9LaoxsLlVwuKsDlWX/pQ+kkMOFgXe6qs07SCIzX+9flRJFUd
T0whjk/xxOf/9PwntNCb+KXwZIthS36wuSp/hF0wvxDCQxThR16CUgbIPFA9smO8
F+ZA5SpMt+YxfVevVKRMJUGl0SYMPSEq2FhvgBLwwv9t5y+mo1gdeltfpmP9fFIc
A/VDBiSffuUNTi+29J1k9KqTcMWIvbOwF1PYwklKwYSqCHTVjR8MQTQDGLv5iXIp
jMqdgenW+7Tkf06iUPsvz/r/Deuxc26XBYC5wj1mFvQvBSRA07SjofgQYeaOB1MX
rAAiSI8OBXIbrVDgJoG9pPfCLdjRYuJSfHUQFmSrOSra2c5FmKDsT0ZTafaSDpou
PRUvosFkWmoqg67160aG9VnFBcn6QchL8rrvRkdnQ/nl7PIkbTWFjsDkcmeJGA29
VNBWeNvTSq+BZ9aNObGKJYNiTRTHCdOhJKu1JLHWGLPPp7d0zWyNJfwzCST9iI7H
QFPPXOf64Dc08lCWC5PD6U7n2w2gqPQbV2K1gWaQp2AAmuMaraNfbvqfx1IN/lnH
RhVTIKu9wQMFEu6OEKIDMGZV/AZbFRYCMFo2Pzyi+smw2zqFHMSghAXbU3HOfN47
kzvaL5399t9bkDcx6+b5BR4JsLnvTYzdyVLS51Q/Yz6NrXUf2kE0JIqbCpINl4Zd
WwQ5tSeA9kQISZy4u/opV0aMKXB7pz0ac28a6RmI7VSFVv6Yixm7mgsUytLxZka4
bwEf8O2cmzPz+RcOO+NTJr7HEMM4W8z+kRRRyqYf/uY7VG62e+XKD9Keq8jH7LxI
RxRr17lxQ/qQmxVx1xjTKWXrHmWsmEKpwEfAAOUnEIbiDYmVf3/9UGVt8XhWuJ+X
+OwwAq0QyZy2Ey/B6Ce41b7+5f76ucZGRtFoXXNM6/WoLQZyCEwdRTXuDshX1QJD
cH9olGQNHxBBZP3osHZ37p/TuU9ThT7cRCadCs7E3n5hAZ1jNL5T09sDxTjUbuSO
kpmiKzUqs47vftDpgscfA8Q5uFkNihFCATIFJeHNv+QTXL9efxzwDDcbtYH5qkfN
sEY2LGbCIgwIIWKhSnfhLHl+9m8Qad+A4/7oj2DvLypah6HDXqcU5WDbTQQqsOez
Cp7X7D6KELTQ+T7cTvJQ3xMIyMTV2R5aYLaw85j8OucY7Hxc8wL3X9WNfp9QCIq/
PSAP2uzSY6u01HaiEMDO1M32+63GgYLBkXwUhlymy+HqJCY4CLzhsa3ijWTY94vI
uESiZLdY33TH1/dZVidf/sPcFYp5+K/YwuJnc5ol07oF0uFQFC8MmKH5wh1vfSbG
0gJISNbiVqrxCU0/wHgE50I9woRShGdc6SUcvFZPLt8O2rYhbFzd2k1o1bMD31sY
uGec6OkrjP1FgAppoBKKwg==
`protect END_PROTECTED
