`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+wZs5+365E4igECy1OUIEjKYrK5aS8BD51EljnolEBe5kdGS2V61lIsC5oUfWrQ
pGsGuBBrTjp7UtZRWipYaUMLwmXGz+S1ZJJvqVnjhwLdfT2TDvKu49ICsUzym/7d
xMBDGx7mWluS43xeyyv3H00FjTNHlwUPAYpzgiDpRzuBy773STS1iVpux1XoEAG+
/dV4HONxLeqyVexuUU75erP6O1DJUa7l6k17jFuyPaojbMW4nceHUfqcr9fNluZu
fQfDI37I20d66OZMZXAKA9xmHwq/6lZKN/FN+Cx1kg3M7c+wKg9tuTwwe7bwkzwQ
G+GklmzZK3u/IG3GVGtWaofpGez8hfnLkN2fPfs3BAzZqB9WXdrZttDgSat9xPRs
wYNSwnI3+HRxJSahoo1mOLv4yimLvrfWlYlJw7gZbjwX6GzvyHJnnBWuZ34PX/fF
w18AwApbynTkZJEoPy0lu+AhwPvUJG/tyiLxNzj3ZHhJseGqkHSRy+QSAL4ABYJ8
0caq79GMh8mHvgJYDiguym0OP8Dgg28xboa17DzUzC4yu55QPBsRaowWm/wZKPut
suBNZw6WfMyA8UAfJzIPEB/rrckZ7mvHbrUcSmZ4pfu53qKoGT5x9Q8jfog8rw7r
/yLu9F+jsA/TVCKpTp2M7NYZG0ezWWwLOPW6zcq0JdOaA0xqCAuLK1iV38bjGgmE
3Ke4AeeICQa2H2gOHK276tIqgI82czslAqw/Yyzu2FM+SCHFYkPwgrBHkG8QMGXp
`protect END_PROTECTED
