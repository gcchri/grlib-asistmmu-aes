`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
51xN7hFotkpHb7ksU5gOM/i2YpXJ9C7IXq+l8y7xGEgPQWYAtmKJsVFyyEX4GEvr
tMwYl3oa5vVYMCthlMpoKNQKkprgpheYKjl3EznoN1KJl5ROVrHWBItmGT2h1gH/
ogHIVt7OYRgRLn21Q55g79+/iyAeTCNKSbmajcSSGR0lCPNsFLU69g5jBrEBLoED
IfxCx+63gZsfyIRyFokjqk1oQABesfryAuEMBqqpZsbbBdOzoKRcmawga9vYmNaW
7REcGUrAbzK43kBhzGMNrkVXBMOcr/RgfE4MVIt7YHeVPx4ay1c2vD8Jrzz4ytLv
hh9QlQ+uxbVomBBqYzC41mxL27w0Z4YuhcpxvZBL1ZuF9yD7zcrlY7GRMY1RNf5v
QW1LQmle6lT+i7jpCr8QUy1iK3qH1HxnScorFDyZmx4WX0zmGR0D9H2cA9ntn+pf
5E3pRSxfMW8u5Yp+50NPAIMvsOfHor6gimhS4vUmi1A=
`protect END_PROTECTED
