`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/smfjoXzOr2taynKORX5mWPW9Fbdd/hcdqcS3QAyr5HB7FicxFG0fdS3t4YUPNz
7u9xyMEw9V2Gq47dkwa1P1xcmxfiliHYWOxFLO9rHG4bbGt4kyQ1cn54Aw+KWvuT
FPHTga+M0vmRk3mcxFNyh9qaG9or5QMwuV1hvhktPZCE45RYVnvUwhtqSEHVwl7s
MRYHnw2HIc85t6XFf/HqX2vDQ8/m2bWONZqNOOy3Kx8uhQZAv5o96Vuldumt0BLy
kKOLxzADsrNPGhZmiPqaHSa72Qu2N5C0pHTipCUZj78W1omLNypzLVxqoF5eZMny
95NcfhSDK69KUfYIdGPnpr/qeP7pS2MjL0PSA2rF11DzUEekbZXnaFPM4TnMcDQ6
THqMawD/cY3gLcVao4rmp88dNgo82g9XG6CerAoCwYwZOM1oro6rfykql0hNcL7p
KJtek1ipXwVjYSgZB4NW0eyevfPM/8+5Tw+g2pNG3c6+ttjre2fpGmRkWG5kaQ5h
zH8lwSTOnkrCLZWvd8vuMcuo7vhldXtfX5AiN3acDdg=
`protect END_PROTECTED
