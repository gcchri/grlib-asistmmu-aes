`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQCqMgVk1ReOVTjJTMPIKtNt0xh2LlQwlR/XaBijkINIs/ii7uTJJnnPcgxza0dY
AbxewiixbDjSnJqhMS/pDHgL3F5cfSHyKgBaKAhZCiIFlVm1fP5Xtv6Gp4WPNGjv
ttQ6Y15BVeB4KAAmom9wZtlG8WPqeLP/RanhyBBIbv/c/Wxah54o7WbC1kmXvGAB
TWn7MgGVTn5nyDl2CVXFBL9bqlCyAa+5I1w9rustekiuT6Co/3mB9GkNmS+cs7y2
ckxPC1JqsbrYbhjEEGLASt/SI3lTyS2BjcdBJaq25qa+N+eeZxTDJWoF0yzoexhE
j/Gz49bY/zyiVa8Ea8AP9gm/GshPJ8xTkliVGpcjLtSaMv50q1sqp9zPneKPNYyG
R7p8gTN4wuih9M0sno0UcNhFhjCsdiERDERBtXvJZqMhyiLozFjRb/+NqRtZS9yB
9pSQFHR14j5oELhhyq6CH3hinl6Uu0m0/gLS3llyAGOh1PcuvkBs9FZs04Xv2EBT
LZLOZbgtHzmfFnu4ZAB7Hfd/c9H5GaZdM8MGfAsxb+E3Tzy01Jen+oDhU/H3IaHR
`protect END_PROTECTED
