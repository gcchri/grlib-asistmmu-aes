`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/6pCY+0l9ijdrKdMWMw30SLo48Dk6iDry7luKO5srPzIerUUWp3FvhTx21DQ2VP
1jsrJO7GjpTSD9W9Fjsk+Q3sYd+vcWKqpeVtFfcoY8fyVIEhpZ18pWgms/EeItZc
1WqmXqhcvwA+dOjjDnRYyEVw1pXwjhmani6nhbWC5Ou+eWZEFMMOoQLhZBpeGwQY
B9fYlfTjTt9PmYQzAyK2man0yhG2kUd1YAcosdBnoy2u4N6ONfTwPlfppkLi4srF
6BWCO92N5pfsvT0026t/lx3joDY0hScPsAVIqkMYT9mWkzXkDV7CUvE1JWcRbzsT
ucGdZlWYoFT7c5h8IWdCx27KI4SVIb8h/1kdG8x0Mo2NZHLfkXq432StPT3DLBsB
SQw/+aQhtkp+xgfVKnPNjqK6E+kJXvuqd9jGP+gh8wpy3CzJhdxfzCiGzNpaojR6
BpkgHtzeGX7K9pQrZz6IoADlm/PZb8myAFr7a+MT2DIu5wy61oCnDUsVPxQH2jYB
jJ4XJMqk/uWkWmufM1T64wkyP++3qZ7NBvygGG+/GFazuSWIEBPfWLdEf4qruU8s
KCGMC1nwPjqPs1kpT0DBXmSCissWhXToTnm02x8YTeOpOruYATyf18myh3JjG9wk
REsLa9t3avDImzMx1Q1S4MlCfplyn0G7fOT6mLvXRlw6pZAB8nDLbdkNWCYA7PDr
jrbNJ1Ofb+uYjvplDk9NTF6c/pTF1pdDgywRwtw6l+iZSAnYaZCPyTI2YQKnyF5N
m3209/MHzLgcToLsv0iFc6s6rxUTWPNhKBM1Sw3JvkkOYvyR0VziE+Dam8vrZMIg
JXnQZ+rVca+jPoMPtIoCeJ3nIO6pDFem6BJBS7iyVXvaO7qxvUayL7uqhGCcSppF
3oSjskdN6khzcC4ttzjCt7kdFGSIEvVGKj6AcVgiRAmKySsvqo99jBXrDVDS2hQJ
fsCkM2G0/ehqNONT6RPGg0joBemYyZc6SCiRemMNLy1cskF8ewNVRMo/PjHAgWOJ
s+Mp4vynrOpr92wWU2SHEbvNMDytvZGnk+DjJwDJNlL2pB55d6/JApkCwxlWunq2
z/DapIQGPdIjIPJB3O7N6l4kDRS8k3zJ6+aVc/JwvMXbvzULlKyqoswfg/tSK93B
`protect END_PROTECTED
