`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZ2kjpLPL8IDPEvm4fZJLW1M0uk3qb9dDhTMsbNfeUyRMm1bBlEH55KfvnrW+dp0
0hY52fm3/7lp8IPhYi2fRH8qBur8VxP3GWVKtJTvq1uj/Rewak8uw0rCe0e4iiy0
wSVXQMQt4w1wX5+U6WO/ktpHljnazdv2T+ZccwoWlIcSR3NBCaKGptJD0ZsV/wiB
z59Amm9Ty5Ol1oq8AUyOWpm+aiDCg9ovh6OWgqQKt87YhbxEW4fO2W8ubsD7mcyZ
C/Bkl8/ZypC0euxwBPSJU8rj4lAetnJN7+abSa6jihyxBPzbyKuJBZKiqauaQ7oS
UdTma8l3VWCa05c+hejJwhwFvIcpCJyq0urhysZpu58adcDnWZl7PT9yjy7OyCJJ
Bc0hXyTj/UAl/s3NyA9sl+41ICBOT0pJd76wzQ2BSZ5Nxy1vs/fmV4Ei7urEz0oz
2l3OEyJROQv/wXEEYYf9GyMjaFGTUYxw7ZBuUI+gQOsZFiGQpHHqcqgcKyb+JZtz
mhBUrCq/27rE1wistUk/wWC0gPDRHwK2VJYPgju2oDScB7EFprta8TMQwDb8eNAO
Dl82cW5YEjo7FyaN/HDu8NRxm9vNKZXlOsQbQLVmJphL6PQLVqMAx08UxGU0cJjR
07GLqqWWhRO2HBpTmWnAsZYDOnsiEUs2P5mw5dEZl6mci++Bbagzidu1mY1x6JOq
2nGv6+gsrXTJOvTepjEGeHvjQBxEKQOeglUPHU8cEPeoNKf3UwZRSbHxVoDT4aS+
Mbkn2uF5/oh2IJOCaByOaZZLPHDXNbdO39zTgP/5n1NyHTgQsRj0pZ9M+rhKf6Od
GTz6VAw0r02b6PVrsRfv2EvIZHZgGsqHWVrGe15BvvRumBJGjFa79jg/PLSHDuMh
lQmOMKwHxWGO6B/Y/eixhbZ2TJFxRNjdL/o3KIx0GUO0vTfC4E2eRHSu1RYtlXC8
FS3nme+0aOWlXpHgLJjOJw==
`protect END_PROTECTED
