`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e/lMmsrlnTll5gYU2GsimKOiC/bQtjHgVtJdgtodcrDxpgriTV6OZG+Nl55Jjr8Y
sLSdAG7hHXkRnXzc1gomKMkc3BKDbjXTpLbwbavD0ZqfLcIGJcQWoA1V/pp+BQkK
6Zh5u3XU+4/3377FlGXA213WHpQy8DzeIbPzY8EWSS4ROMfHaovEwTIn+yuRtMLb
exMjMUrzXMJWfz487DQlwBhlJFTNkPeXRhpyZFKF8g/Z+ZlKrGieUmdd4WvqulFl
0ZKmuUu29U/+9+RJvwCodR3tZD3BDA7uDLVxsa8tpWDAEe5JACxJYpjdnpUBYVrN
0bIezyP2Ucs9NK+K97N2Ss1F6O3F4AxkCmEMwt+XKA0o3t83BgsLBlcb6ysm7yuq
MOzYtv9btnunWtly7WsQ60lCJHCn0NrlOhhaXnsDBDHtu0rE8AQu9/bR2y/F0vHF
NZrpsl2yenwz+avpory7jwA43bpIEmDMiTTkyE2IRI6p1BFahDbQxO7DMJHNu1ll
8/3di2HDyPj60TOyKmZnWL+fYxOvUfBWko7NM0lly5dZxrfdxYNWoPmcmE3pizn5
4BE0EeVoWmwvC/t1QntZYpthpzIKBjFAPiM/+G3SCdqI3DmsW1V94sennwBvk6em
Lg7dI1gX9oC+Nx4PAO8xA8lrl+ikL45eZHqdg6MYT4PaAaSr6gI4cmu0u0s2mgIn
CP/e8JpNLn1HfeRLa6XSf139Zpi8DobOQmNscBqgdLWBODpKqEtnG5zw8K6Tyq+o
OrbmDIg/qejirUPR8D1KQecEfxDPfS1jPXPUqKGnbKt54+Puy/ttS5WK7ZW7Qs81
tLyPIFihBES0O233ScC01DkRevBtjX95kRzvCl8GmWjmQKX9vPpUYCIpILion7+/
NlomjHoiOs9PZYeZkdfZLd7zHiixCk9Mb5HbAo7oi4A0xtuQhKkIoLXo+MRlw8ZM
Jedfy902ZWjfJbRQHrTjhHt7jUW99Dnuvcjn6NeKF5XlDlVFGu5tlMHIdbPlGEPL
RQOAqFn4DCwBZSlArc3CHa3rXfgBjrP0+HyPQtG55p8=
`protect END_PROTECTED
