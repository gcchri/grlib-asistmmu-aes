`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VE1mLvXfUQwE9dVkvtDco8dvKHsCbfnqMKbsv7ga54CsZjRMU2paCuCmZ7JSbaRX
nlVgqvG2gyZrwTzykieZbtA/QidCz0AzRxaSJV6SRnrE/Aj4P6bcLcSAaSBP+d3U
0SneghDsNIJ2K01uY9oHB4iEnzg8YQSq7kfdQMsPbRi4nL+/0b6i7GnKD7NV/f6k
NVRiwcdNPRj5X2AUN4RWYel4M/r24x+S1qc6uGeYgP837WbsQFAyhEzOMpu5VxYR
x+rLaoyVB7dfKDUg2HDCg5756PIeH3CgAwlPgSx7HhFHhKD0lgFHWZDJWBKeQc9i
zBeWlY/3830qMDSC4WRnJRy+z4cAzB0wI1/pHbFR8+BLv9A3NDv142/kswLRm3yT
EVjx4FEQJrgsfOzW2CNyrrD1F9HInvIhnb8mzMWJhYyZV4eGzJBPEu5fDD4E4aXK
Zmjw9BvpG6jtwQOr+MVLvktegLFoZ4pqjg8Ht4cD0wFbigir/jwUkl+YWLR/+i/A
kErHABssEi0X2V+SuDubuNhkg13gRcJRT/mxwN0KESB247W+YiEgYLOiQQaaEJnN
PzsQRMDXh8uoaX8/eEWtisQiYuTClAfvnIS9ymmUs1rNtyrDdFEFJT9uySTmH+4R
3E9z7yhcZW5JK3kEHvjlm1FWqN19pR0Mkn/jmcNLBVS36SGKA/yLDGfpoIT/PXUH
QcmrZ0Ls5VsUC0Knt0KA/MBcUQOhvPHVACULeaGLvPdb/qnimDDPXo6vOtj/+Wk5
5H9BTVYjjrxTPj+VT2UmmatJ/3nZm2DQzVE2O4ow7a5S1FwnoneHOMiMKV9iyb+a
95hW/cU/N8TVhC1U6x6SPwYWLpUaB/vQGls1jFWXuVymkUyO3xqpd55TVoPUFLZa
k8RO7TURiTnwehkLBX8XJZrK0xLZzEzPv2YI3xomlwCJvTdzd6GUYdYaMIvF8U1J
cBJTgeVAZVW8/y6SVGQa5w/1TgKQjx1B8FcVEmf12zYRaZzWSYrlhktSOk9759Tt
cifpska4e4q01A7GKaXknJl6c/dgo8YsOZfa8kpCBCAAGN3GMaXmGOAAU1TO8V3p
MnmSAv8ljd/qOjBa3nL1WqlG4J+gxaSwW1Hciir2e9ekF+0nv05CNQTAILoISOxw
66CZI5N33d7Dyziya2WdUtPIcPt1VOgKt4hjs3UmAACmNHYNoryBYczxedftMfj9
cdjh0KcHfPbqQx+YOo3LskRrBERFIXYFoeQ+yhay0CzBKs3Yg6x0TYpbUt6OHcXf
tsI+l2wEJKBhgKToRWWQd7MPKQSj0wvX26ukIJBTbrDL5SUACpF9oVnDSf7ub8Or
`protect END_PROTECTED
