`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ix1cNyg1IhN2f7lOi6w1VcicnenHvBFEOrduNAa0rsUrmWMdUPAd1rbYnTBXUG8/
Cl8AoSjFO2FOk8AD+m7qnPAE293/HcycwDDiQPRj+hXsUgUh1RZZk9XQ3DOCd1NO
etfBnut8LIRlizpRuE1OsjoWS2jn/18uUHp25rs3Fgb9Cg8kkSYNVpNsa7Zip91z
bhYeaxNNiohxumtRIV+HfSgdnv63TLt0UsFjd4Dp0FAkGWu9h7R4x94q1ncv6GD2
mNsiIzO25EGEjLm3h6j1qvzYnIfivrfC5zHq4MSSyWLV84mfxF+0pfU1aKNBwxdm
nemhUWzIGFTWsVE9UysTPqxZO/nPVIvwcAhgFJBeofTy0aJcS3z+1UZmMPN1SKtg
uB4uzU58H3LuVytTYMXvu8HLLedwXrqwEpjLoVwUcDk=
`protect END_PROTECTED
