`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wWIbba7hjXDGCTMhZoAmtZWxdeN4RSdSKPz3IJ+KSGvmV02+BNffnOoadSxwSof/
ORzWs7Nl7tjtUwUNOcWvctdSMIfYpvATLKyc6JxcnoWbOEzgMvCADHZG/5K0fd1W
WJuLS0bMjMW348DxKlepXwSi2mqWBsy9EaITYHzXQuLx5khixTgwQ1czkdWqk6TJ
AbIozjqtPP2j0PyBVJMgrSK67M49odyl9FEoRE3SVQCpo7n6KVGDceg8iZjf2gmc
nExEgvp4PwHxA9XSAmrclaofZrQb2ChWn6eRw7unBFcGEN27SOuDtXmqJhCT98JE
nRuLZRxF+fTiDT06HV3LLD78os4DOYTnxLHzR5osWscp4R/r9ByrkGLaCVGHwTGC
bWPp6oonxHEuuYCIrFeiPS8pQXRcaP2GUVtia1t0VU33F9488aVPrse8CRWP44a0
70EIn9wbk9L8XxNd1j1aZklsSGD1FuJVsFchzImJWhzyuH71diItEXWpBTJXqrXe
HncDHgH2FuxBVnUlfVXQGs8FVqs96PwQk6xYeDqwdjUqkV1pSX60iKvE49IUJ2nz
GBFBZKKK4+k7nXifBZOchYiP1zxY69Ujf3mIuhqfJACQ6hP475OV9ye68AJQZFFE
jxfJXZh/6hgQFLswy0lMgeDIpXHvmgWgqHlDxNO+0yW7eW+caFz830GMJkX1kr0X
fJ9Pv5CW6cFb4nLLIT7MpQFOJHUooNAgEItpZDetGWmtmhgnnVg8R4YZA8wOCT4+
jaWsPBGzCi3We5o6W17EfQs0/+01GufQkVAYusQgJkePqwnVHVa20BExJ3s6WMrB
wExrPJZtjSefNeGkXa5PWmbVRUXY7NIrKeAaHf+z2w9FYj+d2ELBiUCzi1kwt434
QjGoFq/y2m9/G7yCwIyYGBo0ZnN1cwb4o6vFr+1jq7IYwEQeODnLpoU9kMgMZlEb
RoXZ+SCqQVzc5ccPstITOd+tST3/cUItzRGDinIv/FpwxOgPwUAnJnBXghczN/kI
/JNxKq6AjPrVJWr7C5Ac7+CmAAjjJHJ5v/j/pRneENSkuwA9k/CjRA3nLcWvCit2
PQr2lI8IYWRs90NtRUPbmDsEqUFnf8sZpRYNbI4BobnAmOKnq3okroG5ZvC83K2e
y3uFAnvCFkR05FPUCF1jms0PP5yiR1V4VGtafR3abt2ODE7U+JJKd/YOqLCVdHdo
VXN+xOPQ3G7N2+hhJj9/3dfdQO9HvIXHkgYUvnllZKMTJHgod5tnO59GpoBtQz5e
6mv0WTPE2Yk5VC8krehcqHCC4cuGg03f0pIqx6es8QgG9H/TKBbTfc+jin+xhEE3
GJgPshR7E+nxaAlOm6N9uiDXYTOlGEHkKmqtkmI1CsI0O4pNuAXgu1Ov/N0uJSKu
L5z3WnLTIpOP9ews0QwNUD6QxSimkAd/UVpk3arz0YLQgDiLylECmAuapEUmzJgj
AkRXwP6GAZ8zKceLP0LpVSBYghtpzzD6sj62OgSdbJ+A9tSlpe3auzYZYsoIkdjX
JtykS9Edyy2UxxXrkf5JDAkbaR3YRKnRibpTu0gPWw+c01xK0majBIXqHOYoEG6P
xV7DE57GwnrBb+rnfuDPGr4dNnxoZBgJj9HlhFbg/QbMomaqmvJR6u2LDtUiI9Fx
WXFWrEWwBj1uSnqRi8665j1tFFtkfRT+2/wKXWyWVXy/FQ31tqEsCc4Ywuq9AecE
`protect END_PROTECTED
