`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/rfgmKEgp+bSuDRRWQjyGXMP4cqDLhaQF7CtuqvqsOb5UgIe9W/KJoNoQ5wTJKB6
zSjjAJg9aw/1gEDuvMCOBMCV8mtp34zZAlgXj1+vxqFpUy3xcJA2x+P/JHgNoHxu
sZscgR7WcQvZUecEKX9UlQVMwEztn5gXLC9x0ZnyVbmQR2t1E3kjA7M1tUpSAZkX
ifoUERSQ7hDf4vgLOd9t/C3rYhSbiWOXVqrF5HgGrDRP+xLqe1dRs9V+39UdSG93
Tj18RyFxLtRicwp7qxmNWZPXwxhHUI0rOGB2+ZFkQAu8zHjiS8qwx0wy2Wi7EGSQ
Hw6MaEZ+OTxWC36mNKVZqvePiCSdK3L9vvFd0azYBupMexrkdkEQ2jzdoY0FQZvf
sC+xfw5ProRXCI+tVhD3BTK3tuSh34RbyRb80abxrBvXDj1lYKb69sXxk0Iu5gKG
YmXhqw4JHlam3Q/rwnQ0VTjzqDMd0PWnkWbxkrH6+yTcPIshQMepYi39HHEKP1qv
200kDCBXWU/3Wo1au3MoeSLqzCAH+NLWKlFKLuVypZeg4W/nUQxsfVbW2d7vpCVp
eMNLq1DpEeDpe5NXAdigUpLwmQwxWs4RI/Kdom2oQYMr3bhqYVkgrOy8HYcQM/1t
8eXCNejPx3Ypeld69YA9r/V4rfyaNb5CyH+9jmhB5ohTTcIUDyGZGgTUmZeZc1mj
2oLDH9wV9Xu9bukE2+sKWeZvzF0oFFopBmNF44daIiKH39EHg8knFrKsfYdb+MvQ
YWAqUCelWxIvroaw0Uz3ILHmGS1ue4RHjaew9tio7zHMYK6rSWBrIltXmXLidhso
vc1n8uPwSYz0ROehg6wSM5VraAQFfayHm456SUomqm94STJFnyHa2dJUgaQhZSgH
N7cR8ns/oRNYn3nj82GcBupR0Q9ZqvfwE+UtqOeUYP9m+j2eUwZ15PNkh0bxneG8
mambY29txuh0elxXE40P3kcMsBWTNrk6NN8YqbToLW5S4jgUSghvYXqVHKzGeJQi
D19YH3Ddx8evieNy8cBAlt+s+6o9zjcgZYldEbJdUa1DxJaUr4WbT7X/j+EgvsFs
IUdncIolWvUPghw2ddvz8urya4nVJgmGoi6Rzsbqpe1vTj7t5YsoJtIp2l2DWo7F
9XTRueoNSyPJwPaIpGL6WtSjju+QoSUhIuQQ8v065HLWMHl4vJ2lipWEDzH2otjJ
6JzGfRrdWeHZVB/uFMY+hi01OWYL9HdOSDu6KqIaLwUgQFKi7Q62UiU9FDR6HY73
c/Qu1GH9G++K8b5cg2x4YPON0WjMTV1iECRnFHfaccr3I/ypjXOuJxvbnsqUhFKY
j9BQHMFL8b05AXbe1qKcXedFciCcL5uhA5RR9e8pnoreRMLDpfQfx7WGbo1pzxKP
XKFzA+5ANwl06EImmR6AAHgfmJdM6aoANpD/X4uznah/xAk+NKKrUV6cfR+K44SA
idigkekob0dZwg4Gm1LVRF5S1xQQqi2DFE/sPi4dBdxz/C5xE7UUat4dOxcGmRYF
LxgNOQVw9p3yv7WykOLlRiRRyFBOcLddtef+TTOkIF2T0MqJjb8D+4N00QYUBQIO
5k5TH3QdWk8Y4XpH90OOA+8Czy+Q54C7AyaFGHLzBzg0pgkJHlA3LaSWRIxKNHql
JLKlwwEZir+/GKp2OfUmIgJWMuPCHT9gvsk1bu8AjGjF4ZhHv0+cE2UMlXGFcPht
movaAheqR1SbAfVjNSpq7dBRev0bdG/E9jdKlYx6jLBP21bvlnVWzRSOdgcIOWXS
M3S3lu1Yha2tUSx43QJAePXabOVCTD8L87MEIlLM++pHgVsXv6p7719/8F8ogq7Y
dDvc46/3wnFhJ8Fb62QxKgpEFXkHUotoe2TKQNiRA3QavWJ9VIgkBdNFLKBnQbAJ
h2N81Wnn0k440LPaukL890tiqkQNAkaJZYsHszchVTIjKSBQeQ5IIC8JK2nhFfqB
xWmdIG/2AdJdO+oKnR4cV8WtlS5pc2H35FPZBD2NqvK0+zjDm3+ISpObTbEE2Mr8
L48UCeIMMzrhxPWdXjE5eufyn9+7pwTLHyY9NU1UstmhpZB1eSW9bjdH8+GsmAUb
EBax5J71DKmjZf+xFPEOZHfKUy9hsU4M5tPOFZIUG5kbGeLTApcxuX4IatEwTXEl
Lz75G50Cm8oIyNezov1ZiJL5RAFM19b/BVIT/zOAfvELrqAy9wmUVKcl5yOI0KpE
HU8AGGx2X09p1/Xi/uGc+JR8/W27rYeNMXbsEOPmxfmEZMhcTOjzlQR7wa4QuMzP
EcddTKUQTiYntzQlM/3R1/uanY1REfvXBPmDYTWty35esE2T/zm2yFvBuxI1H+lQ
rq1YXQzn1Ex1eg7ZYy7BqkNhAGSptYldHYuSidYdn/U2xdEQZhfadKSCMjWXg8xH
dFXD6q5l2djrX/0QPCmNV8wdzuBsqeTSDtoh2kPTVM386y1imLStxWSlX7HMGPz9
usXgXdSA5mIG9ktb7tu8wbo5vdrxNaeoyv2uC7qgD/FccOU3fUxEyhEjb+GIjNMZ
Eob9H5I810PL67u9UfQZ6vWeB+PJQJb8Rv+eDLFMBZiumPPIW1hIRAmc4isaxqLr
bBW3QTxQG68mcsvWTzFWco8kQftAx0roy/vdlbIfEMa3MzESMngeFkuCAKNe/H8S
LbN0/fp9svgdT18sAb4F2NUx39EAKHYR2B+9sHnPBdjTT9W4KBG9gBZZPCuXzjj3
51eH+qc4PGix/Oys8bsGbe4SX8z6oz48flwsM9QrPUaFKYFgI1pxfATol7PYawSC
7b8RY3fo2m+OhLrHtReQct1LtLFMFvAnW0sEJMLu/AyVjYeRje4JV2i1L5elRV9H
FyJ6WO1A+gxjnlpXZjKJKajYv+oOjKLjsWbiuwUI3UKmc2BZhsOQIHFDlSKC64/c
QiDFMCGPZvv3GkSS0/zbs7vePiCNfEAEZnYzvMEpvB7IEJZHeHIiA4M9qqTa1pSY
65yBkxcyV4YMe8vecQBoMNs65JbiHidfX7EFnD/qNgahMvWK7oDpIvsTis2SqhCI
UJ1QxkF2Vru3WVl3zk7YBjkRNkU8UxAQwGU+qCwlfonq1meVl1/JllZnDjRB7m1s
nbOHrs9cxmi1ajZIQotUEIZWWuLoHS8uZPdsIh48sdm/QWtAwl8kDSSsg75Hfwag
/2gwugx/Mdb4XZTaGZoD+szMYHbOYaMwKCM47tKiUGqDCmweY8CcAkVg4kf2Y+FF
YMhJawy6OY1wOLCjlOx+gh/Pwyt7xaHHKYul6wCLykc=
`protect END_PROTECTED
