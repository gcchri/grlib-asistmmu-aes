`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/gUYD5aLQQCkioAHO8JeFx3KMlnXmuDUl5RDqrF51IijCfUOCYfGuBn+ZDxq/Du5
YFVFlq6p2734IM7NRsT4TgEQ3v4gEmU1DjzbMb4VWm+iWc5VYd8o319zZqE3ihGN
asK+4FMHvTLgmu6a9If2HT2sJ8N1lpej9bCpc2lPuPLtybVbIAkJUVle9PFiSKPA
CS14hRCtJJyGSAGjrD9dVy2Iyr69gGOtDVJWkVzEhOcQ6Blb+s55kgd54r+qqk/x
/qqez/zlsjcOMsShphcSV33QjpWiPpGXh1MwyedgCt20nJG3sNJhdXy60FZHqARF
nYE6aQaOO+45dKHcWZ5+0W1bfMuVCcXXN0A4rr6W+C2vYwSuLTk0yM3h9Od+RShm
hcDYAQXgyf2yiBO6ixMsUjW0Z/77wHDugbHQgx5xpRsswhHOSyu8+Pitw+SdQGkZ
`protect END_PROTECTED
