`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KAsigZ9oeDLAgiIDdhEHljBxGH6VNwvzKlW5C2OcgwImaDZmN4Lp25Ga+w3/Gtqq
5NXP4CrrXE9vSNJ1OesQsZsj3jL74EsBag1qq9QUxQDDlBomy+ZY+I+uyh2K8T34
/chOmW8o5aPqdBOqjF5lNlcWYMBHW3tU3awZX9rykHYS8vb2jFtA2FcrJKa725DQ
fItwY3SxyD9p4joz3Tzzh/o8hpxotFgApK+BBImyYvZwVSBCbOuWTnqpM14oju2e
i/SFOW9MTzAM0Ds3kE8Wu17BO/2x5pgLZUmdlidmsJDfAtV7pAcDerojE/Y9GB5P
JghMrXekRmlFzTxROhra9A==
`protect END_PROTECTED
