`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Nq3PVowlxNH7yE1vc+Ickt8LlyZbOejpWM6WP8oLkN9HvlL6eRszG6crpxJbxdQ
tlQ9bYp94YJSAhIEP4nVk9tUrklizy1fhQhjGIHRJ94o1ZahnhRxvN/5Xz2bNSJf
qjt74DsBHMn42zaxEXCvN60Nji8j3hxk57abFKr7stkR+0ggY4vxKXysePl+EL0P
iGRaJ5MspmwCM/fSZkgxFaV942sg8y5I2aLb6XTC0g7nkFgCI1OUCxddw55/3oec
I6N362Kf4B//Fb1FAPizYu/pdzE7PF0+a7BHBuvwCLzg2dzfbQ6871iR5tmHNvLN
0NbqWyfL9gdHdybIbwUfrNFbfBPomyYhaIO9N1v4oytZ1xhPrkMIRCSOdUccZOdO
ItwZli/tIWKt8k+MG3f/K4NSmzbNMvA/Sf4JJzhlgMZy2MKMDRGSEe0tKbtkCW5C
HNeO44bwWBQRDy9JBuoMfPvcUA2Xh+wA6id6/dWk5cJEeveUk3vIEYHaqCsZB3I/
hRaqdqK23K64rm6tJKksacivnXyWEKdCA554C6g2eCnuDWZLVrmQlqSg6j7TntHy
8JjfyTGPPVojxC5wP4EU5Q9IPdqW4+2k4ec5CUHkXtKaxtR69ooxzTuIkHgsFDw9
awRinZsI2WOJsxGCCoXfYdB2n4TSMo4hcF4/mXgsgSMB00fCzpj9Aj0vM/heaZpk
QZHiPp2QAwiTHns+JDIwhMxLFy9vjAWO/5h4hgY7l0Hyjy32B7RcGUW3D8F0vtwO
TRp+nNkLhh5B7eG/gSsku7wArEYWMQMYsVNYQyANgZPlwRrpETtb9/8c7Ul2Olkh
yTdUpjL5nydzBFgAX93kzMI0Rs8tGsPgyoGpyZVk90ZcJ2RNJ1uEVFIj7KvF/6Ux
PhjFnYep1xcoE7U0vTePGp4B1GNjrp6ryvYfTDSdh38xCd5kvN0HeyfBPRTIgDJU
ZKfCxAu3NMdG126y6rOCo1AhQBaGWcsjcZHocunn873WdbV2O66bejsP3UtH2sYW
hyTPuZBOa+5zroRXhMmejueox0MWoofHp9EC74A+VSiaHmwiz2PkyGWhi0rsXFix
qfuTjMAgTeyfX4MzL9En3aRT97CDUmziau9rFJF2e3kjYuCaG/lvByxfmrAE2YEC
f5qRX7u+FOa8llo+UXxhCwInOtsDuf3c3ddVLiLK/Pt33HlhRp7MWrHnz9+FT+Mi
w4d7ESzBZY54SQXmDVGRTRfTXltB22V4TxE0D6L3pxUaqEToaQHqMDhxJzlqKtQR
B2tkkPX4loMM/y/RxahQutoZeYeEVxtrrqfQM2vvqED+7LfuOJAchvrnjRaP3EZE
SDecEaK1Q4mNEcML89l34D8uuKqkJMVGcf6e4lI+oLCThw+gj+e9OiP9HbT5b4gp
mT5efhRXogOEfADH8ougFpb4X8tQ8u4UT+7eE0pb7zSAjFPpoSxCaAbJq9aPMndY
Rv6Hmggm3WDgrtCoOai2BSQFZkcmuyoZr/y9pXtoneaCUpyfUH09IjZDa1rmYk+9
TCBgjZAH6wdBylfNKR23u4+iezgZ819ISjA9MlUvtMWXqOwRKnLA2mTaii5mcHf0
hDV3exU4YTzMhMw6QdfBcDW9zzGi9VppfVpiwcI0Jz9Nhyp3HaJhs0MPjvb2tWkW
WCcAACHqa36Vldh5qX7JOwM3G3FLx66uwjTviJ/XfRtXHsEZdfikgyxvXlKuDFe4
2+2VbX4Lc9+Z832maQMUiv+PWyZ6qPI8LUJjR7Mtzo148cU7vDY4wdfuFqukbri6
0IZv/8zK2iskmvROsJIm7QU5JjJB6hf+esD8K38+PpbWBBqjefta63XMMqLSsuGg
BG9WsZrByctVrGc9rj2UHC5LcrSvqNNcUUTP7Pb5FZY3SCZBrhEFMRPIxq7QPUfi
lGlhLvSJxq68cYpttMnuJh0DpXjHyr9cDCM43zXtWDTkDcVyP6RqkdXzio1RQvz0
Q3/whpQpAaz5E/v0huYsMxWp1SBdTVeVqMzZLnVUBaTNix6qy40soO1rh6mTDQIv
lt4SvMsphL957UH9JPDwU2ukJWt8eztr5D1UXby8zVrzjxs/71EiSwwyh+PPziOK
UTMdJOPTXI7nsz9hvZVOj3mdkp+7JrH0cy3JmyBL7v2vRAMpnokXyrlRMUCllHZl
PZKqGbY3ZY3uQUx5rG8XjZFupMfKh6vugi4C4vp0giVRuJNFJcen4Bgl3Xyr4WyR
B7MhXkUbKssWzdhg79T8DMCjECy0IilSvrFSerFwnkY7axQTzlVummXrTfQFZMIG
Erl5a23Xj31JvrvSPZvngIvXoiT/wI/3MphDYX9k8F9CO6BHtQbe5YA2QEyhxa/G
cidjVvwWUUFGm4fqzILX3+nsCIwVfEGz6djJ63PJx4UnS9hcWPooP6ACE1jYYpTu
ZXL8VuKoNDytyc2DRy5drEROAdpM3bXLvrE0uQzUOYs/iYknm8sI1tC02Igg8zRQ
UrsHkbhe6qN3TNkvqJ/fcAF9Nv9s69oAQwyqiugN++HXyGvPa7d64EFrANbTR3UK
P8DGPmQkz8CGD6rScRrx1xzr2CTQ8Diny42XWXEfOK0MUkY4mDedfalRZUzo0X9Y
M9c9VtFm/aGniY5hPmBY31uokEvUJoYX2rlIkqHHxVJ/Ru63uHl6PpvXO8eloZI3
wMQaNDL2bMtG8nh2dXC7aEPdoAlCTueDBER/yoakJAm4zf2CdKSWX2HyKpzJfdkl
X8GskCo5DP8NojWsEsuqMO5hKsSjn6NojZ/nljePpwa1ZgVqtpdYM5Rmra1m2Xlp
QRoNn9VW1R9WZI8K17kifgje8dVd3sdJfYyOy1U64x4hvtIRRO0XUA39oez6Khdd
Ipe9VhF0N34to2kUpX4A4iLm63QHXVo0KfqwNsgIAEGwyw4v8pc4/JMzreQGQ7bc
uT8euCdNXNjgPio/MlOviGgh43aEifcbnEUU34Hhtwwz5nqdErXoujxYdGS+af6m
vCecs+togDSZZVv3ahkVLQs5SGwNRLhLPf4OzVgspn5DN8kdDqaRWDUJ/P0fGkb2
2P9oplbFSVNmFgBt7cyNlZUrqi36j9veQ0yQi5GFnq0=
`protect END_PROTECTED
