`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0R1Rw6jQYc9XRdZ1FVB5ZXx32zR1F7sfKc5wKNXDBvbXw3bniDM8qkCKKYIPV3vp
+cCgVa2LDFLEyyfoDVSZucJO4CflcTtNgDynu27+Odf+WTam7m70Ppe0N4TlTTGW
cGK5VFnUOJZA6dnNC6z6RxGOqmBtv9fBksxdL/UhF1GFa/OLbRnziMAclJDBKXUo
aVWyBz+Ej47vU+X8dBkkh4oT1Y3v0cISYbZorXPZ6MmaJLtLMqEiYl4GgvkOU23p
suCpYGEULmv1pX1K3U206PjlcteyquWbb9U41YrPkRXZ/zVKyYP3OVk+7qGkYOIP
3qRqcf7cNH6CzB+/GGZlm/W9Wxl9wmMADYC+slgXKmaH57TYvnmwsbp1l7UQcKfU
zDGxnYa+0+Eda3z4X81ps8asmD6MeZDUkpJ61CuPtksNqXbnqCwJ3EcEZ9eOyzux
iq5cc+c1H134mucwuFlt8Cmix9Jg49+jF6kJH9mkOVc2tuFi4NL3k6XhnU9qP6qe
iS4T4Axou2jzYpuX8Zgf148YFycIK8MW0wYarRSAoKDjZWbznHjzDsEbOpboPzWN
d0a5aW7DVhkUIJ/YqQ3oIQ==
`protect END_PROTECTED
