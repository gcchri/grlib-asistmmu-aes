`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qkvFXf9GP3+9RsFOJJ0DqxP9v2MT+hSc5G4HdEbgxyooJ/FLQn9rAdyD0EIGbwHY
qDIEMLa2FrG0xodZaOvAcbeYRtrJSSHmxIiECG8ylP69AAe+nP2SaI2xUWzevXgE
UEbUPr5lpHZt8OLE4GS6TEuleSqMl9hWSTEczwhvLQts6fkOMWKeN7ZkD6IR58ST
iKJfvBJgM3qNvNU/HZIhKhOolpDoD/7WjtsJG4qSBectnnNAK0UG/RvWBKvGHtCB
oEncWh0yN47jsbIpfuu+8SovYP66jbDv/WcFutvxp0LneNT99bV27aJ9EuyWJtPA
ugfTU+i8Ssy2sl5zOntpNLWx1uZzQeDZY5LuOMvSTQMKhh8AC1TwZgsBgQJV2Sd4
zyNBx0s4AS06qnD2Ft9AS2dHAl2nL8k5NQo5JtAwJoRlbqYAgjg4M1HY7oiAjVSC
HGmmH9dDmcGv7B++95syhO2SayEfE0ocUR3I9X0Zfusg8wrDAzWa3PfL81DadTDS
IxeY2ETQVi+EFzIWqCtcgTnQJqxCOF+WKf/h08dVwLW06zNzKIVVENF3IqTa8AL4
i6XhvqqPMmJtnY3tBmpzAaFQU2ir8C+u1VB7Mz2ArIBZScEx7qC9K+yKBtCIR/Ck
xDT5IwAYthNF5dmFjqBE2UHj5k9eYqfRfSI8MiKlYaevRBVmucSrCMW65Qrspou/
E5F6TmfrdT844780d1/PBGxof5WG0MD+TARBFVjs+dD87eKASn5LNdKtzxv0of+4
`protect END_PROTECTED
