`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXoJ/D9ISPhNj6OV+J0TUuzYl/d8qy5kfDbbTEoToua3LAYNkfKFTqrOicVKka4F
XgIrP8t4CFmtkgfKrqafdCaJ/ccPLdErUR6DWMtQ9YAIZezK2u5tFe/nD0VnmqlK
cng2bM0TlJWP3i9OD/g7JR/6OdggK2g7RXompa5p/r3fF29pqVzJOzOKeZtJM6XR
CyK+4GXzkoQojwt168cvxYTHGED6Cd8oaGdrA/7unXK6Je/I5DOv9HzsjrxmRDRw
/px03LhUumgDqddOReHn5xIFuwC/8owPEbBcdazBvLUtlY6U9FS07M48Geabaptj
C5q1fYL1/ZXn8Q/qSuuesrvHf3rKdt5TZgOMUnwJNPnhj6N8LhdVQA4XhRHbqKpk
OupNfCIyLt0X0tpmBtLjG/ppvBggwKUZRLwF8JZo/oKolt8QLhaMZTwd0WElyxwy
NtFUBTf6GEbeGmwho35sfjOefsQkNAYINll3p28mjLER4DUQeR2RkeeMSEbm5xrt
4nCWw1g7hW/M05zgN7LmmU3ksUrGG4SUGQ43HKuefrldUdyKZuDbWE6GdAV1B/Hi
w3RlBGvRpg81cjg2FBzu26IOf/mpZEeFKEysvLs3eAsQdiK997Oct/PYxynLf74r
zF72H0tvAtuX20IEowrH9+rk7dwWPfztFSxfIPWXC3EF92b3O0pJ9Afiv+pUSfbZ
qipPYdpU4p2bYt4mPuv3VLIObfHEZk39xYVLn5+GWgybA04BzSiF3Mkad40LIDHr
EDF4Q7E7ZtCg+cBAmS8tYpjKHqqThtZZdkJeXzgbcTGMujd5RukCtfha3buddLRH
fXJv3Xnjddye0vAwxwZJFCq+hv7303knB9k2hxAw/yBjcPdeUFPrzFCgn70xlxBB
xDoxiA9XUhQFnIFpkU4XAWwKbJfQ4XJD9S6rY1OASQSRU5t1jDI8P5hzN4i0RpBu
uyi37HaKGtcFk0n88jTHelwAj80hVHfGDpCcvPbAyKoOBIAEz1L8eIGolBrKFW6S
vgNTvJkk3BkQoZJMyghJ9wfeZnJoAKvxvQZwv5ZQ5GcHOILSUHU8a7fTIZHZh7g6
0KrJTABSkPMiIJ6f/Wjoun1iZYSl+PKS4lqiUeRJbnaPKXQwSwboxkAG+PwWIx4E
WcOknM9pLAD2kG8MUgC/yky/wThF96fQTH94dkSjlroJ37NdVVx9ERZuIKogRXJZ
Ea3pz2J3O5krowdBv/c8RZyHNv1Fke3/qcZpXu/i5GMrrAOcFZr8b69E06iRsHYY
h7FnEgSZAseRXin923/tV3FqExq6EF7IcNPNnVvHLpWO2G+UjE7yYrpPISRDexLt
6tfHrydPT1u88uXUceevy8sIf6cEOBVtuhpLNo5BjoE1asvHv11dDWjREHrps4sB
gUiO0TS11/v5agvvIRrQAlzX3Rt8ukRd17YpYQYVlZoYGQ2S41evY7415ME8ih+m
AbCWZRoX2jvLgAc3OXkSQ+wPy+gxoWww63eVVEiUSk7gYiDVxxUJ4o69wwUT8W1u
8iN/8kLOVRnAnMPsZWBCYnwxi18sR4LowSKcW5Am5PsW04x1S7XktH0ssRK4ruVv
dO7OGrFyEYRzrp8sIlP7/gxwpUTMDhh4Iu05PUBAOEQRBGdQ2btEspDlwcXWsA4a
JYvnd3UqUMfDkQ6BmK7TqjotRpXjJ/vG2619gE1xueWxI0GZazEc+7onA87jsjow
FYTV+Qq/s83yuZ2N6qiJJvpIw4LgpCD18SdVFp9wONHEvxoLdKzYzlCc8/slver7
YtJJiuTJX0xkdCRSASz4o1FfvdjbzH1MXaUuWrjAj+0JBrRrzYNLOrSdtTGVYIyZ
gZ0wUQ/ewx6Scase8tji2pSdZyh5YqV1jsetW49vVPXCIxGRMuyGUZBkczhjn9Kx
VO7z/wzGSMPZzdklt8/fdoQ2YkQd25pa0kIs45joClHP8xzrH2u2iq/iVWKNDnFj
3ATAO9C0kZvAlfU1vJreEsJHlU+pKnMU+Qh5pAO1guT3D4t8GPjiLrULvq71kP/0
jQi00o1R0d3bfX1key/9B8dwoeyb6+MYgeq45wgV6ejZ7zVw4kz1uqsX1IRHOAVd
MekulpZNGj1UDDmVu5NGSYRfqR4yZqkEjrchAT+2/8Gy2dAiGTVdB3rliOUtMFhi
lvzHAZi3ITZqYN/ZG2F6dpESW2Xv1jcdA6npPQdd7iz3KBpNUeS4GzjaBlETrMNB
Z5QxeaKF72AwB6SwM9ay4w/TA8MDAZobDXApj3wOrWGLuzDttzm6BteGuJuO7euN
B5NtCwi7Wqg5AqgXp781PConlUgA201dqEfqGZsrV+HL3tXEvZ2aWuytTze481a6
fBVVeuVtmMGPwyW7bLykt3D9OV2K6FLSpO1FZRm7NIn5fS2CzHk4yf3wbEWDaA6c
Zq8iP5uT1fipRrRIST7+9rPxBmQoY9sUZ4pJMX7yGliGDU4SITOqFSD3vJWzgMUK
J4PxSoAHcCrx8h/3ZfxnyQF9UEN8fEGqwq3MR5LTT6ERTDn65pXt8JKn9RwWEpGM
Utu0K9F0pVbh8PADEtlQL0pOB20cDKvEeLNOiA+P7xx2ynve1+TV2r1qF8xbufCd
uiPtZtx2Wp6KcWRcDzxgrAU/vnBx1JAdT8eYAOmTV+XInOMtVNlJJdtnu3KwV262
e7dJclD3NXlsnZDoPHWRulxyoG+2/TChA0o/djM23K+1LT5CxD8IBYMoLuJS+gS8
/EkJ6SMzyW5t6+EjVp9X8gsD06W08rEOnfBuBjaEpotY7V/IqkL50gp1MTDH5nnc
UN52Tw30LB0qP7Nu93F6TieGPrHoK+PDvLVj5TYPud1P2B1EasQCbIngg+S50MYk
lgPWjzCx/AeQQp42ma9dhbPSXohXHcX2UCN6MSTQQAGrIitRPd5Xo/4yaH7KMARY
fEbmSvyBu/jXWarzr0RJ2qk1lhs0RA4YbfrZUD1dBW9YR/Dq/IhxnWbkaQfr1ENh
e7tvPQabrB8qoeUBKlRtp0TbPeGMNFizngKxc+K5YiDVu568w/uUM2G9mZSy4RAP
zqDxHhh9cWRVB3DsolEzUW3HGkRBJ+zfbq4SxNTrPBXFGK4c/6gZUKGdTZintPz0
Ujx9AEzS1dvwUTNj9lzYjPzEob4X56pOlkiwpP9WZx3MIpswf/vwN5z1pGnI6c8G
wgHenRCfvxS8ra4TlqE2ub03pRGCI8sVyYT5BXjEq44fLrkcTRDG4AA9Ds0BktCf
rRzpSDjwKGsotFLHLnRkc0g4sT8QK2R3JaSmDtPLDAWwl4cCmtcvw2t4jskb460f
OIgr46c7gZOIbC3s/1upQwBb1rMbNUoFFfsJ/1o447vSf1GrWMZNcatfwZMn0S1b
x+lIZPObTuOHGXhRWM5Xqf57Yq3bbdQPVVnjfXciHgJdATJZdHQDBOvcLxbqw7rP
XQRZZF3fnB915DrJBTWVJWA0uSegNCIlu9gPPQg2JfJH6aEaoaHBiDDmjlnltVGt
OvHSnw3XWx1TbA67aOdXqmXitI7DEHoCanETxrvxktDjyuJ9sl92x996EXOZZcRn
/AdNBwdq0oloImm9NUUWvix8JshrLT1HUj00aLhALzqh/Ex5pEMzDjPSNbaq0Joy
wzCtQuB11C7fmWU2pJzqALCMtnhLxvgl3Upv/JVmRlAKrQztntPFJ4JU4PZw7hI8
ihsvznSsSUP0sHX0m/QrSqO+QWU5HWEcvZM2kIErUA/qdww3fxJBzss1m0+0/ThI
gfqxcZ+cV+QwmEp1akjPgqftCAdcbFrBTK/DgyQm1LlUCE8W7Luu4pxc+ugpBN+v
G99/Ox7HK5iyx8UXkmAICtI7vjX02+Kv+bqI2Rp63hDCD0wXZCHGL/vEMDHjF/ZZ
oNwsobVmEEN1bb+PQuapMP0pTVZfGcwxmn42Np0MqJKdpI5mK97MY+L/+mOjWWWY
Uf/7i+98DMuRlkaPkFT0h3MGAx1bQY8r9HyuefbVMR+2RwW2weQ9WtvXXM4HvJ00
QCOvy+bQ8WCv82NzBC5ugPfo2nB7UeJW6CQV3lKwQPuamF1SIslXJ4BPk/LK9QP1
SsBUACIuoX/Psq82euWT7VQopVrv7F7Ztxoqv2VTINmHX60V5K4XlrsibpIswS4P
3Aa9PSy23P8zasQkv1vyyacS2EolYhuhLmmtcVVO3tbGLaMTTIi623rjaUjQNHqF
7lZNWBbeLEg+52BGPCgREgYn1g5oFPYoX5SYLFttHu9NLvDoljG3dSmgxfQdNcNH
q1f4z2eAfb3sOPHsSHslLwyXHYBeD/rmGxkOFaggPst5p3TcdO5Q93eC1GTcMP2s
GLUfPtScHM8GF1b9dfZmhIHNk615qgYLYIQ+iiFqujA4N1F9ypMgcdclKypOSNwG
In+lVudt1nmb1dOvKnNDYtexEO+3DyGMlpIRcaOR3r51ZcYSpYiIwSnhl453NXZP
rZHw93fep8aDog5sjlSYP4oMHyxrQXPV/m5bgzJpuus9XSWGDPga8swUlFN3m0Fi
gVA+1Tv+ivfDf7bLocirRo3PsYXsl5140nHQwtAe4DK60J4KKQCei97mF0H0NZFo
RdfGrr/lPl8RaYRZMStNIxqwt/QmjAbdlpRlDTCw7qz1rsqnDEyvfTTNRWA0FDfK
HmvcbiNEAl9Dj0nz/lcM0QC67J3o/yjDbu4Il6ya8meVC3toJa7pRkpbd3Hbf79E
ylxXjNyHdv3J07Pv1asEVh5xTGghSyEHXOM6gbdAAyNWcDADKfBrlpczw3NvY/1N
zjgYDyhQ2JBEB3ldeH1VIKGTxkACutcdzSGCbIDO7QLE9ZweWsu5S4xHQGQUqiOV
X35mxrrBj1GS2QwNiu49OGBGUPq0fOkzY+0DZ1gyVYQRZn5NPMMlcJOAerKL0/KV
VUOme44gZpUX8LJGYJQOXqlyQkIXqCaktUrDyaEym6+HRQw9+dQpkiUdcQtC6NAJ
+7kuQGuwUtCJkZo4P4y9BOYmzm+hPHO99J1oiOLFLDG+tsusMpzqfFO5nb9B87G7
MJzgix+A1UbtVXH4VvqnAY/wMrybihAPmn6UPjpyC3ZsmHWTIjBDSYYdkT0EVFXb
nahi6YGfZtCvphI+BXyUp5+yrWYKNQhFLodxN96VRe/ImHoFCWByGwUz+u+Tyj0C
1tn/rrz46XFibR58Npxoe1B77AHxomu2dTA5jZG56gbfrHY4xqjXLuDq5rThM5MB
6Ntz68sqj/Lh9rd9MWwao+a9poI612/1hsUshoot683YzjIcGnMoUOAyz7nyctWD
D1nZGUxxCSijhvY8N6Zsk9Z3RTwFI8lOq0qhzSpNs01hnp7x36y+JIFNpeRLk4F9
msHyo+CgYaB9CjZriOgk4mNyYSPWvDThm/cLMT0EGEjL2hZK4bnKyuGNAZe1SQhu
TnXvEYT2mnW9FW92mylfJV1Lv7MATwVd+hoAEl4VDwXQC6sDiUI/FsYVqX9QVq+V
iIvwnyDH7mU6ehyCIk+pdvibFzhWOpZb3JNz2isrzQVG1ccekfn8i22wld0mDttq
mBui6xB3J4LnFQElfWJyDONzPwBYdxZbgFidhaeRIaNLFpasEn8Rl19+8b9/DJ7p
WepmjKtw4cwueMIMVv2/p0lP9Y1LM8GrfwWCwnaL8G/c7K0CqSW3U5urpiXHb+aG
QaC6kk6hXGXAORUb5O7YYPIS261ywCa/Js/IjkaSL+g9h0LEm+yLt5vzTk+n6GzA
S8aAmXjpzoqQ1UfW68lHmgUl9D2CtSMpQjhoTFgdEUaf4IKcuzuPrRVYm3si/HCs
d04xTJeHvtdrNiSEex2vOqgaNbmDc6E/Y0iUn4yrz4gdxHx82qMfA3syf/jfsIwc
e7dO+JrJxCJGLidsehuG670hCpRCU1BZXmRQzIoZrK2jMHL845D5M45EMSyC71v/
89q0NxvYx6qfSwdHUs0ZPWuuQO2pf1vmpwqy8TFfuIkfDdvnARQKtWjyiD6b2Fam
USGunCZLUKtB7Ae/4uaHkiYSusBJ5BZKnu3Edj6DtyLmVlt9wd9RA8m8Z/bdordh
V6albhbpYAwnU+0dWaKtsphFGn1WGxAV/b8I+pCBbHSirCI2lRb8bhFjf5qfDtnJ
U/IGmCq4cSrFPhI+VTpejVijyLPYA2SJNb7axcHsKrpmw7MZdb1ShcwGRgNt0HQh
UJdWpiUX+e/Twi5mqQbYdjSCnosprTndSoHE0+Hbg+0VWJNx2LtECCQxi2Rd7VDZ
JHrWrIqp1b06cYiHWKUE4S/2U7dU9V8u1egdAbl6JShLWK7Yayf4QjmotpoS8bXo
CM43lufAyCzK2/ReytJmSt4RKulqiScQB2bWcGQH+yciljYb7f9Q0c6XLZnvZRGX
O20mav9oaYg4yohwSq+qJP2DOLwmA3xZmp7POiVX7oeJEC7/u0P63nXoZCRn6MTD
MsCU7AX0JTt/oteJZivWX+lEy2JlH+9jmMZSTiLnPpIdFB/gMf3AtF2DMWF+mCBf
T5ruWdb5i+u3aRg1Gq4IoNnAJo0EKn6WM8TuwiRl9UK7+osSpSjGxtzqZqmStYBw
pHnRQiHLMPzSSooI1xG9o41nNThQY8u32CaDmw5YUBvBGdgNp3zApuacQJkKSWfj
7WZIKNLhQPkWAbiAdOHqp/bmHkrC5iLMKzahZ0G73OqyGJVgXFhXI4iXkgoybHka
sawwjpmMbQREpY+i/KSc052q8BaWfp5ywY/4iD9eb1A1ug994TKH1kHvxoMv9Woz
SfkTQddTbfmWi61mVV/fcqHavmOBxqrkP5tIyGzAm3PmAJudLILoNRZb5jAOEZ0o
HUyFkSHt6NZWv9JNTDVr42mhmvr4HJEfvy+EvfHTPN1sXhoBOdIy5RymSgE8em0W
2CMnEjWWuZZdf3wXrP2CHyON91bQr1JX/dmtBCS2Oa+yuRx8MZHmLbntM8Az7OAj
ZqyltIvqqrSk8WDtHlsXAlKb34pADHwyF4k78svDZYoL9F7rQZFHT1H/OiduZdWg
D3SBsdrO1bHbOdMVp5X3+XXFvahpK6WnBDqc9XqJJvEPy5Ckg5E8hEk+aQjgYNZe
uWv6plwfKkGY9KLHUFNcsYDrlnymnIhlrZeQev2FyM6Gp0YPTEVINzjajbb17MC8
n4xYZJ15E6yVTEbmXRL8PPH+oOnToqRGvWGSgL6XFpsEr8Zm2jdr0LFV2QQsGLm7
+/NG1rMTdAwf7RcaSxpbz7itUA/5U8HW08N+pwtjyRRCfMWOrg7iEHbnnY8+ei7H
7FxSsM6YWeQoIJH7A3I7sP4WsNtFxNv6RABxokS0zAmYXmzYyhwn+FlhCXp7STUD
U9IJHAy8i+0Bv3CO8ssGxYwGxPWbn5uq1LVSkm0bpZQhOOs6u8kmg8ftkq+4G3T8
RzIPYgEUDcf0uovzIyXiOKtlE0QQLqhaYKJmJ5Wg2SOM/BZqB1FZvFiXO1zfHvSY
39iyaREOuuQCvqrkgvt18P6zw7a+RIlx9AvjHHiogz9ol+5BSPEDsaQWIeBPo2yv
4CDv29tDtKhGQKDwgYcpI36UuFUNMCWYL/wY6GlTMxCBAkkLpzTW6NBs3Dz8Vcl+
tXrTDlmCyaftflfXq4DwCrqFrLEM0xE50nLoYLJViIBG7szD8rmUGEA2iY0ontPg
OIi4/3hY85e8OCTzTG9CLaLOoKhnCSomw+Uh76Oe7rpCrB7i6QdX62iNakpzFOqS
ZUjdWVXVCbaJOE0iKKktqSBE87tjGTAjozUzMz81UlmHQ4qXIi1OL/kXJ0yLngEd
vzEuqOPbG4F31V3LgJqfRxyBuLH2Xl7bmsKGBAIhMkSk2PAjIHD+dZ6NW+cxKJCj
mD4REG6i/Brb7nN/z8MdjooRR//nKnzt3AUfqbEUOE/N8WxvVr6hKTs4MRhHWzFo
WO6j4a2EEFGfVQJbez5iY0T3JzK4weWPoLHTJnZCLDf7bWMjA2HqeA/nZmVZBoYI
655QB77gqFh4eCxhGuxArM/If1egjSSY+/4NT73hypRVAjLDYbmp/mX/gxjSux//
fPrN7KICJ8QaxfYgp9BcDCbSGdlOImj3Xw/itnPoLy4k0WYhHkoYVCdpnheIintE
Wl6P3S+gKEigvrn+V16mrXPbcrn3ARmNk+3vj9Te5CzFgPF1QwGwM55lO8RWaQ3i
CcXLgVU1b/Lhv/ZkmK9F4ObOj88XFE67humH/O4jcR3GlLdDld42XfHHF9BU8mzy
VwypgzdU+9e44kzrhTwj/8jzsOOQy71kzDNMkX20ekLS9V9yufb1qpE4v9zkD23P
vwlwRPX6Qn7Oy9NnU/hOzUFw2w0aDfvcFp7fncytg4noiBhBsLiVoiWzuciFbbTG
OP1q5LEMciqLRAOV1qihHnMLD7mAqgtyWX+ywLCN0kbKvv72piMaHLaPh/imp5h7
OHb4XeItadaIdpFUxVXb8mIdYkgZxPthUdML2pWaYv/of1Df0K0ifEZagDLQhQJb
COHy6Vq75cQlY5476Ympvhl2hgA2h51Zqt8E37IVjY6Rm3f606/4PN7AQZA5zSPk
3XEjbdbJMyIKj3VPyEdNSL4LvLQcF0C6zsiJkTRLSof1vnSmOVMIqGWXIitXh2e7
5PSNfuLPLfPDAeQYxieGAVzPDChKQGwXfnUYts+R7B5/WRgISyCs/TfIO823jscp
ACsP0/9oxAvXtuI/vMjxkasGsYXYzhHalEmJExmkArKGljwFScUNY+jWYKm0tw7I
DTYwPqV4e809CIcKSFwp/EL1gVTTUqCskcMVhEkgrUs28HQRVvNXS42nSkdo9rCA
e8ZuVfdCC7XMDCwoNIpH1FU8CmCQapcEGPJn8ftwJ7VMPrE6XxCrbaxU7MBa+cbi
KKMCUs70ADB9DsufO/SrrXf5MDV8Bi7rnx+br+ZFcmw3eWS6EP9rJNf0coZbLfby
acFzsnoodBOreXTUognQlKJuE1ttOgMTjX6gjZ/r01S5VgWkGn0yKHujuaKsu/wu
ZXQzSW/+w8+AvxikS27+wnJcoCPAPSe0PCJf3/LSKcmh6eMZ6D0+kG6EYxNfiQ9l
JXmyRtofWsvmLq5Xr6CF5cpHoDFJya/W2E5HMA2EejaoebdGJUqqWVLLGNtlzG8S
iHG3SoMB45J85DN/5zKWJMrNdn8XVYDcaJCJVoG/NrzoVdk9xlYvQGACWoUntDfk
185GP/2qts7tpBI2zIycEXiIqMQzpIambkXUydy+XAOo4U6n98UOXifY8kkEJHWb
v+EH1hc4T7thZQjXwazpt3ra2ButvkDhqKFgmTGjBHZKQwf50zATAsZrDbPKMMWw
F1EZ33auiQKgtire6hmKAXGy97nPazuAz//hifecUqJJVUuzkdYt41D02Y2zdmQr
92wGxYNFXTQB8+h+LAcsZZRDh3BrddK5PXZ1Wa2UqUOD74s5BrvtnkPRu9k2QTiT
HAPCnZ5KCGvLBGiw1LE8M681M2tN/5JK25wp0B/Bs/nKOg+23Ctl5oryrDjgKAuL
5+HE7eRG9JsvHFiDrqZTAjqUx3P2rLJb9qfmMtVrm9TyWdupBCmcPdNYIT+5X9gF
KaRmkqCn229j/sY0GLyk0cpZbKefdyuFE62n/rpqabNk4ce5VO9lOAX+lv9IxUYG
+qTE/8q8d5CVTkk4fx5bPSjKrYeJ8Yqkm5uffiasSgIKPlDWZwzndsHOB5G3uelK
Ym4fCPbN4seQjKkFt91Pq6s40q7oYR/uZZvoEQuqlDHyH67zdaDL9oCa/Rsewka9
8BbTZ7U5Qat9YT/nbmV00ytAAOJBlzHLZe+Vx2DtgV7dbxqOvay+M0A3RRchgMXP
GrtBztlOQ1vBUYvhY3PlvPAmz/X5qN4RldwRbzS1UP7T1V+mzKI41OODpgETz3q/
oHvaPECmuK+ija3yt8LYeH0amuKT3uDk9PmQuOmrqgfYHnakrZqRfj6gKksUOLCb
rFAfdMls+mB1whR5WcUx4r/3h4qYqVhjEegpfSlFBVUqQOBCMgatIx+uZn4tvHiq
J4o7e50FRbT+AYi/yTpogHDEefrdSkUsU+RkYwAidJ98N8aYGLSrS1pLBj+CuXws
kQuRRzNdhndlNY7s4tC/h5xiw2LSJSDDmM86PMmc+iwgnWJuFWgFJYObrY5szdYw
Q9OLJ8Poxj/+TstbIaHchq+/9JMcsAV5xcDC39Jnr+pxHhqMxAKBwvDGpXGmW8VH
+BfaFoBsjEsGATslYbQqV68iKbxvBktzk+vBU14iRJRdiNCqfhox7Fqjj9/H81Cy
NZnpEZNZ1gfksSA47cPRzFD/xVcEk59QFJ1KL9SR/eGcLTwweT2KzBXxGUBcNebl
T49DoKKRhhEMBvkOHv3Z+AZnewv/ZaDRH6dxGoLKqxtp5b+u32BUPU69I0FhOwnD
YmLvVH7Ukyyc1swUT9RkmlhVWW0FYHB53OG2hEsE5aQOedcTltB6/V8qZvU9ewYm
9EbC3Mfv8nufa4dD0Fir4TWK2Shr05duAN0VnLTXtZ5E3XmoFAlfODjL+asjnJfq
iGytr+/ByIfYwtRMEkWqhYte80xQ6HLHG0/FyTjcL5B8IGGMZXwim1vEhZeC2pEa
icBfY547W838a1b9f4UlYUA12uaMkOJxn6SjhtsKd0oU7DAq1FVR8GkOIPzhZpqs
+D0BIX9Xf6PY2WyqCTJZaMLWGADb4FEpNj7t2ZqqdJxINuEojaarC4cqKGV0yDqS
L4SFvJiGGS76kM0sTlZpfuiHIHbrvKX2fTN58LH2ZnKMMz5l+968lp0ZbGB+tNb6
FzZFN6+YgkBFZRjiLhh8/A6skeCwY8MEv8wkmXMGktmpc6Uc9ZgGAW53LWuorxBj
h0HijrOxJBTOOZ0IkMKXuYDbw3MSPwzq3+AqgX2v653pEzci406Wukab20FwB4uG
JqLJNXYF/NTfdt9+Ir1Zzuk+4pKGgEaV6ltlcoWR7v4Cyxov3Y1svLpOSa3SAwPh
GYLYEI9l2wbrzePpQTa1SfD14txSOzpJ0g1ajn2HEC6/lbH7sBJgwj7fzPmJTPOR
8WHTaroHFCTVBdDlZogwuRYyT16L6l6fBXCf8Md3KeTM2JBUa5qXw3b+E1ercb9y
A4vKZtsY9m6Hpz19loisDamQLIv6Td87vt+kLIi7kEi/l1qrjh2AQzFcclnm999q
+2CWRfUk6lttHzxT3TTaVfRJoVO909qBUDXnBsl8ROQ2Jykc7fyk2V4YPJqhvyCV
Ys1RJuHu0nf3SI+0cyIWrpamsGY/7AvmYVlCx5F+zJ39ROixilbIIDehvAr3a96v
vYlJGRXqjHhJu9q04SMM/8D6EhjeaPoEStfq+qCJ+jfe1MoOeoRYQvdgJpqGOkWE
6psQQy2KhOsVoKGRuPl+R01SQAmdAHlCvPARvIlFWWaPNixFmSbLHuLI2V17ZY8j
6ldw3PpX5Mm2zzXr1kUBn+nqbWfHejJFnNPGi8rN5gLy5DVkYcgGVM44yVooxTdL
S80otai0+lPtfPbqMj+wALOxnKwTI/g+iDWwmDjzsCLx3QpKbmD6+msNOSZgqJyo
fZwpA+zNqIUw9Ds9RyXP8Sn7a5IY0qb5KbjBWB5MaktPvUCT3ST5GWiav7fIPJVN
h5loSXbNySx+Z5DPwE1ej7QK4IhUXFea685huA907FSosyjPl4CAs9IjB3Mj5ecp
XLJsQmXMTbxktg55kax7Qk09dHfxQDZXzL8TH6zB7y4HGNb9DvDdCjuDeEzE4I3u
DW/FMa/QtYjfZS5kPwHOngg7A7nKYeZIIGjSwWhEStT/xVAOpN4Ng9u7Pl/S6tzE
tUdu2wmhEPmQYXL9Gn101FiHWngQ4HYgLvQntUQaGlRhxIuH9P7O4y4ijpODXJiR
zIR1HUaNCCWmbBq8HsM8MO8OFGK2GUUe07NRGGimWYPuB9kARthgcDnLeI7vwO7p
XiD24oRBesIcYdvRUT8lj5e9DGpPv3cioC5jE/zVwSBZDW8+FJ53hDC+EsLonpFd
UOpi64gi0IpyLkX4szqB2HGmsKDhacct5YZUbkviUF7T3PXGJV7349UppGQe1+tC
FSX0kTAVoOK6MR4iJXkjUKy3UctVBt8wCubAJl5JXUskzN6bnIGz+H/RfptxU5xL
lt/bmiD0NzYA9czHkX56eTJ0EU0Zt644gjmDk7HUMCoJDi6YssYX8O20ijRBibQa
l2pa9NabgHtzfFPuTyhoF7s5i/yh8KQoL2wwzXOZVtuSRDsMvaJOUPSRLpQNWH2P
+IfePdxEJpsjRRmqsOYv7LV/po9omau9zqjCy+QfRoc+udiKnWovnpMV0Nu3NPCY
t3GOhH+kslU8MOY/UcMBjaqZ9o6XfWTRIvZZA0HOyY9gXq/D331x9Kf/Jyr4Pw8W
ItLHFt30QFLxknUk6nmKbRF1ZsyFEWCuonPQvHP3I7lrKCmI6bQYHnQTcN9q0rfG
CZAhwCZQ0rV/uMqikeFrFiqHfX02KTOro7RPi5MBFuHRVqm/Q9TFu/1WErwchZUT
WuT3z82vY5c2lFaaXGZnWR4r9ttUebCOY2FfZYjQMh0jgyrpEl/EJKasjRs3A6Xx
9mH+Fyd0TF+i11Hkf1s3z//77QtMXhsq5wdCQIxQjgPFuBqSyyFZphZZQR2QwvNX
Xnq8d2RtFG3EGKBvCT15U+2K4I7LtP42bboy9J2C+3+0LMxbDlErcVVe7KV2k5mZ
DCNaG3GZFeBnCg9eoHEvBdeJ2Px972b5BPCql/YNm3PL2DEL6Ovir4tc/+GBrDVc
7wYjXF5iWakeUYCycNohvlJbmZ3veCHWiZk2IxFepfRTghqp153h5Q/KZqathz07
k5Oia24mg4/4QFcGuWdRgqW+6f3Z+iIh95JD8b61PvFuFwTfPianx98V4+XAemux
51fM/Y8w/PslXGjrXXskEpt568cLuTLe2ghYeblidLTdtVR/BDVoWq3cukUWcsoJ
nDkaBnDGeTFkxTF3sj8LUmKwramjCw+zT0hcQz/LurNiDas9Z1yu6+mWMRFyypJN
VtY2WyO8xbDXHS2pBhma02XcLQXJSqZxMOQJ3VrpUds0cigt1RsETGuE30DxrCze
2QTrjjFaY2qVxLF4aDGfglN6mbNEVpjN/QPxDDsmc8JIyTA8hzIpBp8MJwI9WLgy
s5Db+sPqhYsO1Zt0Tfim184zWKeg4weRoBoUpuRtDiV86QfiDZsDrjIdgeP+SzwW
Xx1Jtum4H+dBhMS8nw8k/1I4wTf3kph5nEELDcP1qMnXw2We8K5Zr2z8hC80CE3+
lpsx7y/jyfmS0vatZi+iVGAT71U7FDB5/wUOTYqELgpDK6xOF80Pnxy2UyFyLDAC
wmesvDW1AFyvHTgOJK1ZEnKjPYkOY5qTftUpdsiC8Z189FA//lVfoym2DJb3+0KE
yS5msGPIEEkKTSLTPBNUtVf74jA5i2ILhzizcPiDQHHRi6mPKDpNY1x9+CaKVCVj
dOeb1ahDJd18LzvGCk62wb9MzGjekX5hOSUl6eS8Q9hZsgozALrxl1dzDDmzCLm/
vVqnYwY+NXDHNFPBiiopfLz+ViFjJCwY0MU9I5v8eD7VvGNgp8MtldIM+LOFsQ77
864K9Am9P2e5eaVW1BP0qSA5IHXDbhKSy5zCtY6xtJff55sfB6MFbQFNvTmQKlmr
Js5gHmESRUOkWH5dkdhH3274WVlMYOhaX8aaP8WbrQ/+UMqWgfHYfZlewsHlUjx/
UyvYpwJ5F3jEBtm+b8QFeNtR1qr0IZcGzy+AMuaA/e7hnc1mHZp4hcLDn8FpKiID
m+PfKjjuDT1o0kyN4gbEZvTJ1BQDItW8kGtWSmrykV84BOPxAcjc7S5UImBxWCe0
iIQ/UEiqmFPu3e9iCRPul6DsOb2pEY7kUMIJI83aecukjx0yMCe+st4WqTgJiB5E
Crg4b/7Kj9GJE2eg2N7IlqtbWKbIX3DVTB5qqmLcvXVmPm85aR5CanHO2EESexfY
aYJTOiaeafDfOBW0F51Jf2ALV81d35GNnfPDpln4kcXMuR4bMoESd8SdoDbZNp5y
xy2G3YFIpDiWCD1QZJrH2Brk5YGnmBse6E5wNQfOksXB6gb8Da8NVDOXumCJ3ytc
Idv4alepkLm7Flo/Ge1JHABKRitvIpbJ+aetsHAs/fYE7l3Gv1TqO1nTWv5MjvVs
4Gfx/1hvRCtYCeqDHjislWTy40U6losTNOg577Mx+fHGG4AWZ3z8tm2EuJKdF5zh
sc/PDt6M8IHTaB0mwVJ9ens3rT87SnQooJ7iRI8te5jmUMf+/TfFogdP0y8QeMA0
77om9a5n4AGEcSmlzdBl3c9LAc1DekVbIXKLD91/yg5t4GtaD1QNJaKMTAxRjjBv
tjeF3jPp2feI1RzhY8P0J3qXJTnzpRPoTPIvwjbNQQI1FeL8teGBmm81PCc6Ja5Z
14EwGZh32QjR8/VO8SXQf1ycTI9ZwtSheHIkXMsyI4+MUB+IZX9GN7rTixC0dlX6
KaP7Hrdp3xuxpgkoFbmdguNtRcwomLL+Vkb36KYWcgOOcpqTu0WPXHOq+0ZTKh8J
l+060hRhkqyKfo3luE25oj/Lg/RT2vY5/deidVZobPicvkYpo9NgncMovxwTgFGN
llbSMzMUh5xzDUFhSQ1UrcOjoGk5YYpC9HS7cB/737kjorMAo6fmXUKSqx6pu27V
qPvdIHYwbt7+Y4FABiTKzr3RylaANziegtkehw+CJazzDBn1mucu+kmsKhCXN+sp
BDRtZQwox57jNUlhOXYU15/0i05CMYGZpIVYRBa+rrerRYkyl3fghf+6PcpE3viG
vpw50a/fQvC2Hew8AjUFGosSsnx9AnzK0+hIUiby/dTx/HjZBt3ShGx/3yNhL7Qp
CFGfcsQ5OHAS04r/Ss7ToW0HIRXZmIdg+xsWhZpW0xO4i9cgpbOZh8Guhj+POaVH
JHheK7kUCusRso+u+GHiAKpOZNrhp6Ea1CPG1iRAPLYYEP9qhwRnBrRzSgN2niQM
9rMpCgwlmeQb3XJNgtbHlOCOZykEV9qQpfQSy/Nt8IeVpX1Yb6qJ6GIidvAL3NgS
MvP/uQxBeP+alGyc8cHdn0ukSnCVpZqFl9ZpFUOmF/ylC0nIZaaeiDnWuoim4Pqb
hkVncfYWfSp2mQ8H8jOEmuOPYMKaBN4RaB9F2LvX+zMAALDlyqE4tFJX2LCIiH1R
Gx7dOiRxxDCo/XLrBnetUkHZTaFOk0QbYTCvQlCEmnyWhy70IccJLvzBMPErAJUX
v+PUqffkxvGsKgR2NoGUYfkzOygctQSf+LI0+72cotwwnqWoxH7YnbSkacieuuBH
JZZZtvdG0qS0jsSa8LojaVsk56UMMb26v3kxnTrXU97X8ulKVAe5EC05ak2Yf1iA
VqSBHW2wTx7f2hN+n4XfXrH2PvOIeIsBAo1LulDyx1xBcJ/ZgsR74VUSAHnLbyR5
Dtqy+F6aD/vglaJ0WF6fTGYMG4kkOHKn5PREAfDNWzioaSXLCnjMlEb46Is3H18e
JUytnEnzJ0DN0a5LRA8y+t691GCa/o7EKQTwuLubHQtmG+kiaTglf4DebRUbVKJy
msK7CwWo9V4UEY5BYYpqtVf2fzgK2U4u5jNf+k8idPlPFKCkb22uCUFXD4WG+mqm
+H681i94zGW3vNEPMl7DQ87dMQ5LlW5+p8XqZK4E/XafQKa+ZmrmtBxics8Xpjo5
y+73cYLBIz4GnYJpkp4fFgtOVTuK6OSnpiqD7e4xWDrPBIA/E6I9N/WZnuNWRmvX
cWW4BT7FTJS8PcT6U+RyIWqq5BDL0Aw+pwPYbjcs22e51J1Tlfs6IBYSy1ATosp2
DN1YEltKFtKi5hYr2x82RCKsHxz1/Gbnpsh7z7RcxwQG/AROdGJCpflfr6QLfbpl
gs4/TVUEGTUhfvJxIpwV1iog+d7BuEryrZNvLinHA/iyHqUhRlp8tAQxtEqBsQWo
MsfPnxQcrOz2Sz6MqoVqJyUuaTF1lxgnppyeaR6C3IrsOXjOQs/i3ob/qe8XXUaU
4RlVH8XQN/6ZSA6rS0RigAMHy6M1UssF7P029Ggq/LlEZYqRAT7TbYwTE7mmJlHR
IFrGeG/vG+aET0Fv7PBoJXTAnk03VIRRrK0Et518mhIFpoxDtGCTleogeob6DWYR
QvGJexTT+m6+l6NckJ06iC9uhpZEZmxJRLaC3MpJpAp0su+rsgU9XpKX9VTLvI73
r9HhbgF/ATGu/u4zqkfBblAu1moG2tkCxLuycbQzvIU/iDIJSBzDTWSMKN8f5PFm
2i6PQArKvN1cnIRNChPedNo4T9XNNmTnJFwVTFXLMHTLnfBSYMEnPrRTPFIvPmz8
rDvjBqWBD6HkKmygOXnPdJ/hxYme/dNlcuEtSKrScep/h9VRSVT6nnmT5LoWbK/L
x12fNnIZG6NNzgSZSKibCoYFUuPOzH4mUlLkp/GcWXJOQ1E/X/0xdXcRQEeMvg3M
Kl1RZNFWEA9aQ4bnfsSUuOabrL5LjvXJ6gfbrbXqOILVyeuCPZQJS3DnWotpKOL2
wFIEt1XKzL5d7N+qG4l/5khYpS/KqO3NN/IlJ+0qAuLNkvyzD2oy1o7rxqsLEvox
OW51KWAOEaZ/NeIWAZMas4fTrHV970H08K03uFU4QJBxF8XVhs0q2lliBsOd6rdc
51q89/H/3JY1BFCIOFEQ2ZMwdmXWE6ox9eedwxTx9XBfRMYVRR0htj3ZJ055j2LX
N6bv+5BrJVXA0CoqCIl1qCvij0mjOs5Q+Cikxt4XfNGuWH/tZsYwzZ1JGZ5aOfWe
zP6goJ8ntBOpy+CVxoNqzN/nNc2hn72mZ877hUCJ7vfeSlfP2wsE0tU+H7FCv2mX
IZREpaZZKs/DC9GpouYvpPpKtTIGtR4UTRfKWmePJxHThFbNDUUqP/qJpUQfeEEl
pAkMeNeM3R5zoeyP7uPe1hhfYB+GbHvpdxAcANGXomteYvx2ZpvhFBWutfRiqbIg
glMu4pm/9+xc0o1DD4bKuyTtkcrbeQ/9Yrcd3BraDBpnh28u6O46wIUT7Wzz0kyC
FqBkygT1kJ7sBJM6Qsnbxj+jT58m41skTUA17c13iYjl6vTZQJEkejtrqJJy0kau
+4OzJWI2vP1uux3l5x9M5dApGD4qDhFLT7hi4v35A6r68yRmjtwnSmlg99FZn81I
lrSE6aDLVvoOuDgUW89ncregKUSMfN50QMUbsSssQw/B/w+bPU2QpBH69HX7ola7
PTWMRhoJDaHOzNHMDy0HswujhFRTESjnjywUvuk0Ls56pzO+cSGAnVWcVGtqALf1
ouwYeYZ0uh6GMeZiauqBE8n5RESWTtspF27xtMilnDK9U1dhgqBbBQbXtCK2A7FZ
d2jfXNPxtbAZaxAX9xkFiVK8ERbBzc/+qnlRiJytTL3fuHv1VGjSvauQdF5kP3uM
Sq9jpxtxdw4BpeLQN9BHuoeOKvqGjUSxKb14jMy7BO72Bceh5XrJRTbwV9tQ3vFF
Q7nb3Ya/C+u31cDkIX9jw+RhIVNJMM315rLlgtPBLFtnbXmWx/vfUllwFbSk9ukk
dfyVQrDM87lf8eNLWD8nIHyoZX/AYWJo0BlgFP9es0jTRJBhxageKTht6tOaMVDi
fgh4Gc8nbaK6eE5AKVYG6G7e0uIoi1ktSIxH2amu/yK2DNV74itMPXnsYm+zQz0j
5l72wtlgghfbdPMbeAismOhFJ+qTuIYTJbABt6kj6RGSnoGBBwdogPaaXLv5YLxg
JycX+9uZnAfK1oMEgkHwmXIl/NKH8YmZAxq6CWAH0v9G6N7Z7KpHHRgCowz7bn5d
P1w4Sdkxfr5G1/ct5ceK0CJyFDamPr5EnrP67V96HhvNkRxPPEnNA0NS27vMEFB2
zg+q9Hdos4xD0u8Ft5Ts4RM/UKkR7snGXmaLdMxcpURxispvPz160rEpuPtJMKU7
MuiE4326JrdNkp31j4VqXdJggJQ85zT2yw+6Lcq++s6FUXqqFhdzl3XZBYLMgmiD
VU0/FFNU7lc0hmeUnAAlXg2nxwrYgQouXzMLWeL1I4lgQSpfsVgoLFaRW8yyXy6i
zJl++yG2bTdWZR/a57oJ7kg4l6rSR5ADPnvpGG9RM+ZP2qM+DVS7S1QYqn9Hw0s2
6mUzo6l5SCfkUwPw9QUGqwBMmifeRxtUOCJoNwiD1L8/bhC3UM68gYyZmT2306pB
6f++UhbpRfKl6UBpzbPUpLdSBmig763q/Xxvdl9ouu9MLN+p+mPz8rjKEVlRlGSQ
PzU7mmdY4P2fvHu3AzT/28sUJ+e+NmybY6B5JsVYXOqlm8GRZ2h6T32qrmgAXi15
gfgCPbmCPs0uUf2DXbZUtkaFNGaqsAWXM8fMdSKvm8t18n0bEmxyCx2BZ0fGKn9V
4TwdaNCFEebZqYPwZFFolsCNDQnDANNGKtse80MpPTtEcFzRsCuzjXw7VTYDcSid
f4dX/u02nDDWXNviaXCfveYLiMxubE6FO6h+f4ZQcx6puQHwxR6FPdmWB8qJLwjm
bBQm6yDQLetIlGCvSh1u3RPTPvbiDekZDED1XNeLqkfPG/7ju/gMEEESM6BJeTkM
QdlvwX5A7IR5omy528U0s092gkK4s/x7Euty+FH50W+pxTfHtuHhdw73qC+ICEyF
6RviuKvq8t7Lv2q+GHVR3tNn/YzUBLyAtR5tVt/b5EvQIyDDQQ99T9QP6MKeUFIJ
2kT1vWuVheofP62sL+hC/K0DENbGXxdAzwqGXVo6X4HVuMyASIBhaEG6+N6rq0Jb
BDYidlUNIl4qqUn7cgcIXfxdZyQRG5yLalQVHh6iGIF2yqn2PsmYjp5dyHwi87xr
bk+r6/9IWtnA0uJCdA1AuPzj1qMqSoCpnd1s9cBgNWfetF08i6ipzSAGVpulHBA5
E6hIYs4bRMqvnPfM24ZoOd9lCemYDZDA83b1AifKobASLFfqfd/mk5q6CGWO3zOI
J69VngzfV3zuLUzgy1pLUNXXkbpzN2LWznOP2DmhQG3DqpWmcSvQVMrP6W2k5CJD
FUFaqAuNYo7Q8DA1d5MAa766X05xHbIr03PMxVQDp8xWs9BE2wFcEEPcWEG+sGt9
G/2CjDwiKC1AUooeeEnazX48k9zDaK1HiSgW4VUEV93OiEHg4OvYRfSdaGAcIXdU
4354+MT3lYt1oLI1hWaRfLfqE02Qatvjza5AbeR+ofuGbZF/zNE2dLmD4zgG9JXL
x1cadFlFBPC5lSNJE+WLc8C48AHo3ONbY1D5qL3+MA9oLs6Q4UlK8Qd8Q5GQQwhj
lWK8/wma0mFw5niu7C44HwatvthatQ20A7lhBJaNsINborNJn+bTWIpWpzA3DZcu
JILQ2ZIUEu0m1z4grnt1VCajsd3FoSB988wv7UYPkNVwRTlaVjqjfQW3XBT9ey+N
lE51cAStSY7pAPN+3Ms9vfRFtmC6MamZoMR2my9ACVja7OPaLLPJEvFLa4PEKoTO
GgbtvhDKVm4i1MFA8Jf+xmPPICsvdEcpdnC1/X91OsphWmXjsIWLB4izPbixjo0g
R/161G8yTR4UA200H4qgKQICg9tgCf+zGraqgKeMQlE+ANoF8Cp8PRdFOEmFYDHn
O7LrBvV51BjeiCUxznsSwq1hQLfqnZBxdJFdCgAaSKB8u36E7kGHMSwccAEOwg6m
89+yitDwkx+BZrOnwI+HP777dTSh4Y4i5VDwDg6x21WWFt2It8MeF28qtq0pElM7
U+TtDXOyuRSXlA9ZDQ3o/3RdlJ3TbOB1mY9jWFqSxaM1eMEAeAM8uSx/RSkTc9g0
oil40zq2QZh04cq60kmov98oNc24ryqHrIkS1DOJuCsqufoJaS0YbWbS5NG5fK5b
oAQQLwf8Lu2MK4PQpBI7ruF24S0O97Ag0fzUlnxrnT7FskowuREYfGq2/VGv3c9F
FaaDvHcLJ24BAMhApzgckcamxg1uWMILl6iYvjbiNKsid2017yR++h9cjd1UShvO
EO5UdII1i953lo/ldY8krH6iny1JwhMvkd1to5jyOU2SWaULJ3SG+FyzEXmHXNyw
AwRRyf4vbm6jYoe0O2EMsJi+oxOwoIXiFOqaFVCoYiODnoHCrErV1C1EBN1gFCMp
iUmizLp7A3uLCAWy0xJNNQCoKl9qbG2G5f9jeRYdEZNtgReM3907dMcuhdYNIXml
hXVo7WHaic/8Nrabi6ocsDVz2y3qrwYkvUb9Qtk2nXKgCXNClmyl+k+slU7lSU75
6FxqW9RqkOIeZ7PywAi8ZEtL6RtHm+rB2pgHf1qeAynQGZSFNCDXM11llHkan+zo
V8adX+/shxvDT9k+f5Ypy9L1DdUwPii6HExxsdGd5e2N6XoileyuZWpbjwpoWamz
soVYhzvdk2SubpGz+dFwSGsvb9bt2OAPYpHcnh1Pb0n2ObpkpWpEz/6YgbQgB1Ki
dyIIRI2jATBC3YA/s1P43F64Tt7Mhzvz8UITHJwUTY+VAOsNLtqkjmxWydJlwXoo
huWWWQZhDvPmwwmfTTXCql6t1rBs0qqtx3FZ5BhsiHESaMTD/WeSteGvWjx2Xduj
qka6CNOapcNIm2X95LL5CD6StYRmoIgZ1wV9+RblquALSGWUZ8wVCcI00Vdd4jb8
8vLT6lWHKg05faUd6Fqelg2XDwr0uQLB3/2zym9ndy3wFWD/CjikNX1Vji6kCFzm
L1qhHkCm6kxTezd8HtPLPZYS0t6vzn7MWe0sBPTTRNzYx64VZSdT0aKblKEpuaj+
tmqRxoT0+lxMITJWwmV0/d75M7kaMubbQOu3q4FCFk/QTGTvjRzaV+MMeJysMzdZ
GT5gb2MlbwdcdFC5A5A8NgS8+jBiUUwgb31N537suV6rQrZ92kymekGb/oimBprA
/9FrCTAHukKALfqH/cS/dH+DkdZgJgii34HXvhBnpdeXm8LVp4OsGQ1LrezcICum
INQXbTwVCrNpFeD4ZJcEB89tPQA6z5uwnWshsLLKw465jr9ST+PBy0C1nimzILcA
By+YMcaY90pvyfHb6PTi7Fo25fv2In31sywucY4IB0ZVN6e+i2E+gbEZvX+Oeykf
d4b2oGcYzWHXuzKkS/By8tyUdwoZQsirfqLyz2ciykcHzQtu3L9sgOWZVDu6o51A
d8k4NPz7MqLIAfBlbCYQ3/JG5cnzMKR6vL2CZ+0Mt8lZaJVroN7iV5/xRnruyY97
0jdKEDcVeod6KS8mc7gUZyrDXXW7wD0QjFEGLX/38prmyGscCh07Ivz0Dz6Dqmd7
8v8Cwp6ChtEIHCYnAJ6B0qKxA4X7ruE1Cbw6CDvuXEGmNZpLnYdaEuwk3sxgJ781
j3Dcy4owkmBCWCjQHSUg9yKFKTEUtp0YpB/mD1TjkYgXOe44LirfjDn7z5DuW7oW
tNjM+deQ2uuGqfYZZR+mMl8NXDZFrW2afpSNzF9XVZ68qOhmUV6PedOcaYmn77j2
U6PNL2pakc+OkMFTcgeHGMSvLDPJuLgH1+vOKGvuTQ8xsDBaEQ7KYhiMd6QuZFMy
RgJBJPGwFwYiHcex2RnVZ8BW5kR+Ju7JjzCtg/IVG8HEa0CEksI9evSOE2FBsvak
DnFfBatN6sFPdPLoO0itC74j702mJnASWoYn2ydqWEE32z6SJIDOcACsqNx/0hcj
gbvxT0TcTX39JBiXYMG9RS7iYsjyQCiLmNV/f6kheiq26QoNC3p9UsJzrwJIJrz5
AfoEMbYF80XgWUFvCphir4s6JP0Nv5ksR3sa9cRl5z42BoBbDblVBB6MEJje+CcT
lyotORaKgRo+rInu5vx7HOP6ltfYjLip/UNDPZTLBeLMCAn6meWuXUlnU+nnvpYV
HdmYCpUtWAS6TA3ZZMinosXkuiUvCruVzbos5pAcYl1Gwcsa9Gjlp0ZxomcHBPcn
qMXgwgNA60J9rpC63g7jofOvnVYg5BO0ve0lGADBJ3/yJouXoW5HGoRZtWVzHrlQ
jNBb0XksO6LvS9juW4T7Ug0tkHpKpXGqj0ahIG4x91801E+28WGHwmw++eLCy7Ll
TfqDzwRKcgcux7W+aRXTEkI4Gd6rLmMuA+eSDXNskEMgZimOvdop/Ty+Flf4W/4Q
WGFmhVEE7SCPTs0l9toRsDEa8Wca5l/z9TDnm6m5R6lnWE2SyfZMKgoC44T2savU
8RvaFizivZuPcoQ20H3h6bzZlg5rZn/E6mPbh5IMUIfVacAgXWj+OZrq7Q2lgxDS
C/jPR9W8GO8APs0UymVTW7R3BH78RB7wA9XqxiFo82qEGefZMRuK3QPlO7eoMe1J
pa7iSjTp2m65oWgidf/Vns8tSqocINjlVGjOaNTtbPBvQ1fOC8yrZtMmAsFD86js
vYRPppdRPuf3JrZELZszN7w7HeKM3PtDkvLy7CjpID88emeuhOpea3vMy2vv3D1I
E2u2u7lb9xK+6LvvK6IjqfMWI0KlVqGRAsPcvam2j18X6cAlETAW3sCl+0TBgopL
/CTKyos5KUX/+KUE+w5FqkQoJrdRmBSA30yY9beXPP1GZC8iWqwlmkLBjBFrWfs5
ZRjAgfmF8DcMmWCoE6NtyG4Bxu+pxblz0jGhb9okm+IuaSVtjHbYXnaqAqHyotym
DaE+0W3iAGZr7FfAcILsTmBpZmBYi8w3dBTzMATA2fyezFO5lu3hmdArCuDjSws0
nLkNvC6VVRwrwN8ieZqIF04LQeVYNUOA6W7scNYYLCsgBS6kfv7SSK0FRa3w01q4
/Is00XZ3f0diCi/C6KhKurYfaQZUo5TMJ3JA+1KvzpythJVCWTa2Qn3+gd1VlgMI
97XXDkt5JPT1Uwtwvm0vjuOn5SSJO/atmxNxPHN/taznRzGA0LtD7YIDEldsLOKE
WaXVGoS6noP5Jou9GfY1dzGqXobeXKoYsUTgQcvPJJZ0/VXDSp7O0GWNOwGg56tE
hqmqTtVXBAfF9RjbwyV9HtKf5F2+UCaUXXmqur59YFxDdaBBd5n82RevgdH168Ho
AsERD6Ttb6GcguuohdISlILaI9urkJzzSJByIUFG/45DAgBmSQ3GmDWMjnsVis6o
ZNgbwQo/JuDopSuBqaa4P1jlEdrvEzTvPmwnWaUUg0VyMUJz01oQ/CcaPznyGrz7
yuDKGh9f7rWKR3uAlkGELm821iF2cL6RFg9RU1fWvPbkxL0toS9LalAaK4mdfwdV
MRZ3t5cu7B7zO5gnsx7u5pg4lK5d5uBTex0rThusqd7UPeWaQ4QuPsCECoGY9y/1
IRxRhm+cwdSDepkq6pHYCNZi/2nk6rlzU7/8x+R3/TTxWb2zBVWbZGpHlvtqIU+8
zVU9rtZq56zN0OG1lze5iUENvz3HPTWIXgvOeljlCEGf57Jy5+LHSn+xVGKK4J8l
tACXUhAtLyldZjlBL7p+W8WwJ6tcZq++uVLU7wnRXj1Q25rvl0pV5b0ryotO7Wrq
IwMomDE9X4Kaj6lElIEYLQDpg6ktYTSa0Asx3aB3N+yVncZKh+aSWBV2CuQL3QUU
pe4cjpX1Sl96cv0M46u3XBqOH7z/6ZxwHFHGghEiAQnrlT3uYLLMHpdMlaYvcf3T
PZ4Eq/1fGaBoA9bcxBfUarycdyG19Pvi9bYdH+Z+lNTtj38XkSg6KjX8ubrlSJ0V
h4eS6XDaQ1SJSjrJbiQ0WIPhGuriLWIypo7OMrVy4oN9hWLK73s1r56dOo4r1a9v
oNEQ4wXPJWus4zpa4vT10ua+q6qA9NnGImsCNjgNFXogTfYL6sLi6CiYV6J+lotL
LhDUfmhlrrx/kB3sWF0YIvfO42I1/ezuwgkc94jhbb26xi2vGNfHluStvF2JClF2
y25G9TeX+/4Ut0IX79K2nKdK413sGjlnldXVIfez7cadfvzHnrOiWbPGw02acZvI
bcRUvxjIwkICVTlu/ibv6J8Doni0FcRXRPI8xx37xHv/q5Q+y/aq46eq5/+1b/Xv
H6EJdeQ9F1sb2vw4E2Z7/HISHN6K7JDwtJXJJogIQtK6rIJgL/J1qcM/NkfuhkHm
8oKpPlmC3A891Lf17A0gzJbrxXrvgY7DxKSE+aL9EFdE+xGHJTyKp140bfyQILBf
RFBcQxg7tC0aeaL0AcV8JUhWvV6PbjKpPtaKbVrViCrmecOUrHnqn2HcVVgkpqsb
yLlqszw2tmkdEyYhIVqaq4BiQ91m+wEX45koELVdNfUecSisXyeWKvO68t+cJ9Uy
3JqjiYQvkYpUUKQQ4mbYkxBQFfmnHfd5ru1voe3juvfGkFdOcysipJP9dsNjgQV+
xNPWwBZqxOWnAuR7qzYHF3tY5EsGAuYA1fqJvdey3f3vjuEblzimlWyZKG0UiO2j
pboL3hIC6kpjpypD+P8irv/+5fwsEDoLLY8I5r12jtpC5wKZzp6LhDnNS4OP+zf7
vRCkyZB6XQHC6qjxHCRZsNuedodjILBefB6GV06SE0aMeuTQm4A0WX6YVT94SUBT
GYVRSw8DNeDjqdMwb01+iz8x6/poL/EQtGU5gfrr8buLpwdIUh2ybZEuel+MsDjn
UKmuMoo05q6uySQuqvcmTuuaQQA0UU+0oko+WY6mIOuff+sp2R5rPdY9Ek7aS7zJ
ZF0Hh9uWw6hswSYK5QaN0SX/hHeTPLWHgu+iKtgH1P9R4g75WqD10rHLkCgzFrsc
lwA0+DirZkPSv2kjw13GZw8zscsQrB6PiLcZv2ITA27L7Af8Jrj/bG+9afAgdB3l
lS/968Qp4wwWlytraRD0lSSMNRRWAUKMmzclFRhZcXVqvAnMT6XjarvkWFbJy2hl
X20WPrQ44wSts4N/YrOIQug1uyZ4d6Phu2IifusjM/R2zIbsYn+OM8F6K1edJQ+0
paqBTaaF7Bilq/BdEUEQRbH/zzNYmeh1/biVOR0RcxSldJq+p5uwsTVsZ1nsOq6Z
wiWeWq6H8J/5AWAY/ykUAPCDoodgCpKhkR7Sk79/D05MZtcqLDIGfU/98c/f5D6f
HXauxRGWBPYqPF7vEvqGwSkVe4rIpTySRPzsRUKN04l+ybGk/x5JFCwifm00q8ER
axOgNtKkVNDi0ZzKsXc+pqwb5bTNcGoJeXXjE+k58NLZYcieVoXQexImSnrOip0M
GrKLtC0ab519bg2IYX+YrN1Vcg+N5ZRWmJ2QnwKDivK9ESgj6c56sgum6C5/nAti
BacmPdG0dfTmdwhXNo2p+eSl2Aj5ZJnduB3kbPYMV0yL4G66hgmN9xxOMvcCTlZ1
FTVwTLPmHcQSU6wGwTKjIZ3tr7dFK1n+eHpEjJ1SCm0r4G50OAC7XqRjyoNtrP1w
/9fCG080OJ/FmGztGNy9UoXRS2N37S/9QPE+vkYiO3wvgzhGDG5761gN56JsgLQz
DdcjsTf3FyZhOvQ7ezFZ427PEMnQrLzjWAAPkz+/xeVYj0/ji/HaJlPmGendaFnn
QUa8TZyTsmGkoNvMj4OMYafybYZSjcU6xz9AknsS1Dm+GyAJReusvH2doA24I0tK
yXlWagxfGIiYV0RZYcHvJYuk+6juH+BaF8OmCkiHRgvX7Y7ujnLE1IxCZ8dnTRx2
bzZMQkBqPPbtjesIu5jlMuk9JTc0MMrKJbaXhHUa4pLK5sJsR/f07ac+FMs2gC1z
hh5OY84TTzgA1AT0KLzNmepj6Bo9U5JsxP1gzWJHrCoQbit6RSN2XUbMkOxCGcdQ
9KD2rWFWEM+y+/SpfBRKHHEcMwq/tzMGUZlqhxB1vhQXy56Tvj2gMHBZBWAqpk2n
UNISl5BHYbcNNOVVqUxXL/IdNQoGZ2BziV6rdkwB+TQXFEEzZbp5LaXVk6TlVdOn
VA1Cdb7+mWsR9PoIBIt77Is5iMupHlh4j9u5Z7rxqua+xZylfpveuH/auQN6TQUc
VaCs6uPXI08m+KIOjBWpPRvmCEQ47VMyvYFKpQZ00+xZYT65KMb/Qf2iiCS0QW+G
PuuiirNX4DzZSUtsAYbUAW0UTUbFGN3i637zwul/x/qjX09aFeKiEnBj3dbbN/C2
xCPnIutGQXlZTI7HuLnSwqFQQbYvERUbzv0OXJ3grQpeYY91Z/Rwz8S3i7flaCuE
QmMgW9aUlc+W0Scejcxw5jpnb3OScR8MKlHX+t3Oi4pWrp5a3emSEQPjT7P9xvk/
EXs+J3MEvsGmhIL/y9lGWuCcFoxflxVSDYxmh0Wg9lr4cBXPL+HDEKJLfdb5o7GX
2zPOTYhdrvqx0oDjKrUhSqr4albkxWrsORwf+U6RsBjlvLmEXQxbm89lu7UfpaTZ
fqTSQMGUk8OH19kAb4fySxCgCsoyeOmvDYMyAC7IdmLedcOA9c7jtU9SWBD6zxhB
xi6ruxbrQVb3nwDg5D+Hew3A85SjL9UmaMynLJFlDToa/6m1j5U8Z7Yhdosolvh/
uU+tQ7McOSgqlGa1Hyli0o1F9u5Ir86AeHY/GZd7NHMUYieeB9arAX0byMlGBf8X
cK/34FABt7ODBLr/weXM00dOfrzars0ML6L1PuWzFBPVHwkTyGEIFkYvEfnZFRtt
fUaDltkduBG+HO3FVFBGOed48FDVNpnXPCz6i2h41SV+2E1egR+oSpAmxbYWfdbB
Mv1+CecQEzyMS8esUzUHGfcxWberjs9NZWO5a6pjLSDM9u3IKkKe72GaTDeyNmUK
u4OEsfV2rUNpM81C9lmiOD1fYV70wyWym2k6AlnFQmwewDnaqzZ6V82UD8oITkuC
lqx6ifo0thApt7JFYjp8GV3+QbOLKxb41Xi7kXt+IKDffyrZTKoq8Ey3BWNkf6cj
/oiGTnMgv6yb5sA2GNQkjeKlsl/bk1h1WhTVmtCwAGYABmPkAfpXi2/28tUhPC9r
i/rPUUonY850vyacdUhi0RKRllRsGjrF9IhFBV7Q2E98YsMMneQIlaYFSZG840kr
Dtu6hl8oECNbT34uYF0xq1m/XJIimH/mqwx0CCYr2JSqLC/b4wj4YHEid49KbZtS
tP1ZqScFk6r66l98cBWmvNpwpE4w6lw+wOQWWesacuwpYWEopWc7J7zEf9qbVEeZ
/xi/PZL/P3ItiHDBlQvVkr1zv3Tg1f2fDxzYaqHROpQGpV8ojACqL1Gel1NcqXSc
g/CGmYgM+u9OnOPDHhPydwQWkpGZGNqs7Hy62WLXIDfJOXvU9sfZTvhDcwuiA3Ku
i3ZcYXuUzWneD5N849T37xzM7vnclnB3PNbZIVr8i1WQm4GjddibAr4hZHSF4l5A
/ebCmHB6WqyP2iK+yh5oGXehDyH9CoqFEglCt34il9TxCesD+2+UT6hO/YcmDnz5
nYffMJphcO30l/6ww1cpZPtdOPFQSmy57C1/qrvOslTYvFrzjA07zD6kPcTsUs5I
5YpQ5AZfBOswghbhaTt7TmdTNd6200uiI2V5HApOXyWGp5x0988FDIaiL/eCCX38
mM4CiXhbwyvgUtAyYHi688KzEX2hzoVdsD106A4UEiiKS1vGZgAwSG9OH3Bsnegj
AG5Ltf+ISNAtbB8ishzjIY6oTGHY7BFOzJ8IxfG/fdd7Bm+1jaljyxe7k/sYK3wL
Ih3Jr7pchKzwIw9zaZQBKdwJdFVu5As2Vl2koFUeYyEb/XLSDdvBvJGVDJDI3rDB
R9k1ePePN2R3riu+ZhOE681V5MS3x5uv57FSVyghb2k9saJkKDx//a/lxz/SXAts
bBQWy7CbDP79G3C9S4MEl7IDzowSVCTM212VS7acJAkQBaVr1gcCtg3ZWFq1BHaU
Jz+w549OCPj77bYUXFjjRVmlXIIfwTmuKOzBW5FQ97JnNaZ3WeYPZ/WY1sqV6XtX
t6NSC6EPynHM1S5M6dRdEdlfA+3CWcsSqw8T8LgVIrYAbT1/K6qmQ5MhkqPs6US2
LlOpwXJDPNdjkTOSLrB06LULbzdD2Md8JrQK69aJqgiAnGNY+ezaxjwbzNiH9ES/
pXbqQhvE4YZf2ixiIS/H9uaV17udZ9Cl7owAaaPJLXHSjY4fiS9CjSg09ePmlMYf
t7wa6XK8f6ZsC3023XVeQreKO/HE9rBTQqU75f0vygRYUI9lxU4XvxfLTLb+Jrn7
94OEb9jWaQvu1UvLoBGrttF47RpQKYWdcF71o5aW+t91rz9jj1Y3xXQ8s+cXje4q
k3WhNokPoI+s2wWXPUV0Vo/kn0gNL2DW89aEKBJcZlO2X6t3O0dTcTDSoQ5mplsq
P8ImHvqMXtJnaMVss5Y0FBslaeOsbPz9VPd6TXHCL9miknJ6D/NtyNF6+B0qaTmC
1VvFxchQWeALwtOoprbFkzbpVnW2LjJFsSgtkzRfm2mwb4oREpjBA+l3SnHKdB1v
C+wbXgLh5PEXFbUDWDe2VriY5/NpGAiHGvsHZ6hzgEJjdWVXk25v4RjGiNlAqHj1
iMXex5GmPJF4VFLe+dctmB7lI1+jnJ9o37Ztn69PO70X04zBJeT2cNsqacRSAkq1
cLO4WUtdTdEE9Kyl2N59UO9Pi1RtyGNIy8Ipw9BGU20Rw4NPL28kKOQnEDRHQY3o
LG6E0nNyYGt8lCIZebGfBZN6bGWsg4vVykaU4QSF3EH4mPxgZG78fMca3fIqddNb
DxN260BRE2TFWmU3fPIUXQ3JrxpfNXWGH9aHp2+s731pnX6zuh+nWnzWwm9GstqZ
Ds1P5fXQJWKymBjky5mCICByqBoZah87KOga1la9sbo0QHFcQHEBpFU27QurVksV
k60U3VcEv5NUMGp6NA9Ky0xu0JvxcAWlz5wqpMUkPESgQCCEJBF7SH0Uh8i9lUuj
ChKF9Na/EkHSNfdUK8MWSL0S3kqnU14RrvrXKZOtKl+0mWQt0l/mmxNEen0ts56C
s+VukCtZex5RooVggpIEvXJ0vg5pQFZum7i35ytrklbTUgECgOFMq5FpMS2DkVQK
Q8ZG2ByY+YeTc8npRwDib6xSjSS5WlPCL3/evPxf0xyE8FPcUgo6G4s8e5iQ5qo0
ESEBt8LLRqGWMcUmBIHA3rHkmEU/s/i9V37aG8zFbuXnoDEsvgKYQeEM4Qbztl2b
zabqE6XT+YH2VuWcGi0SRcAfnne57HLo7aMs1bycgHC5riRMkccgkmMk/qEfuJap
EqebtgJANAsbRuWJ57S16Tgage9qXv8DLqws3EcuLrsW2JsSmjKd/roOCUVem73a
nRvVEqD1o9R+Ej6NxuRrL4K7QAh/b9i05apoxuImXbP6nsYvGloCGB1ql4qaJH3u
oSuuwH1fGVljRZrqbipoCRayKiJAnKrD6rvU+ycUUt1fF88eyLqJ2bMCRZR9BQ4Q
qiS/j88s3Z9Vw+nEddkYKO8NMGomT5eajRuphhqCh7Idu4rj+ouYTwVyTtH4ElYe
/wcv57fc4K32xCcZwEDHC52SMJpasrMpAGD9qdQ2chC9+gktvVrAA/y2M4T9QAnB
Y80llBTL0Y03tIRdahZn3tgRxYpJx8EO759dS0MTBC9IBcztX5eJ3sgtS8Zu7Ijc
hcw6yj5aKvArE4kzA8cvK8+lTNkAU3UBusPAo/f9KGnQvFxJ7JsSSTCu7uNVl9Zk
dEXUUHA4JYHFsVSX9spOuE+e7U0s5cHR9kG1jsI9PahaHRsT4nAvS5IghrR6vH1s
aSoKcwkyu1+nucVZ6QHYO6gLL9628mgity5Mn1nyk3w1muH5x4X7g9wAaBkgzc0w
czCWRERDNW1hwJXJXU9NH6dqOJ3veT2dWHsCvcf83N7oX9qGj7+3OD01K1tEAhcV
uZvO1eDbo8+YYZKVnRgzTIE2bqAY/d0QYe8f49m25JcmNfAQIdDPMWYo+W54ndF/
AQqPxWBaixqSvuTSzLmfweqG+Tuv+sDKyqIjz4uPQQVq+evoKYXnEvKMmysg07rq
G1C5cAncJl+LXtQhRv6SJqWZPwu2N54L4mdTZ4IAk2xEQWBL8gFPwJLNOu4TUKA/
a62Yr0GHaZaFGSx02UbSEJg1JdlUYWqQlLdy+WEoYqiI/7hXdU9bOv3w61E4bV08
LsiHTzmIoBSNzTMv2yxJ3TeXZnPEkcIPSa3MbtvzUoW459lTQtpTg/QiwMl6SODj
iCFP0p7S9ZNSvoQSZONCXAqvJv3yVmHW01+VW1Kv9mLlVXSxKvKDjI40IWpwsQ37
FydPzN4Nn6rGX5PdY+rUXLQELocx3bNZJiQ6FaqZWWCt1aYLRyEUtSwpjLsoG1Mo
TYTiNyQNosF4DVlSX39kkPGv4ffW7Dwo3krKMJDS3SS/A0Mj1cJRAKE1qylDG5ye
e6I7iE8qlexyeiuY5zylxJahpgeI1s4bxaQaFasszNJ7Sz79sfJkK3daFJV4+CgO
nBFSziIOFNJj8/BdYBGT6IsywBVp0zXPzqVqMWzjuGR9qR9YH2ZiFAHOUczKvfGW
/JyHPcwYNnppadl3caqx4tm++7aOb5u8WEfNjXIz1L7TDxyDROtvsjb/h/TrDfoG
/+URfUcSTEDHq5j1e6hkg9vnc5sSwTLzR9/UQsWlXa2cchfuQQo7EArxT/fO/63/
c/KGis7iIMZqCSb9BktxvdIYjoX9sP649wkx/gvPY0glsZTDGqw1O7bN1g90aOJF
+6VgyFpgspe32dF3MhskydbnxLIDj7Nw0VgRcXFkn6rj/M94qBDxkV2WfDHHQ+zf
fAMaaxSPpuNh4kmsmGo+8euMaYLI9fgDiOJ2GB576GWN8Bu8i83wQUgLGmLtqyws
3+AoGehHMCUfpvpabjlayzTEeFte4zy7H65Tg1V7bGlE7UOLiBACSgRggRkOTmOo
tfbQSuGQyQC4TlMUQ2XPTeRrhR7kWgbFlPi4d2xIvW1weQM1Dj5CFfspyGapuG8L
`protect END_PROTECTED
