`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xMul0FHYaPtio8WtBZLmmGT2fAURyXUS2w7aF54x1kQ7sEr/k48O+GTEVVaTSVLz
/8aLflb5dX8KD4S4a7AMhAYdWN/2g/iFxgoTVXkDqWv8WPp1eSyGD1kejrAo6Mxw
2nT4dROpqK2AEnUAKpbRhgzlQiXaSyfR1q38Lmvfkc9ISWEdl88d5Lz7UYXnsipA
6MTcKTs7oV8IaumEHQ9TTu46zoI9HXN5ZVcLJt0k7+jkq3HsW876j1MYV7aQ8Cio
44sfYe2Z/5eWRhzaWtqwpvUR9EWDPEso2InHmOPP3AFS+c9jO376ijVCk7x6iFKA
/rgW9VpUhM0thtOa8J5eAA==
`protect END_PROTECTED
