`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ng7yqU4yEJIflcWzZKpyqEOvbzpFBrNf6tt5B5toD9SXabgqBL3BsECIBc0arSS6
FvJiwElxY68Tomf+ymPZKys/V97MqL9owOOebyzPYOKn/VcHiqBCuKAGPeX61bEN
gDx2xQqzjdBDJRErgZ1oZz/wdqkeYKxwX9Cjdvc1itpe75ZABUUfs3mnQg1D6k+0
YG19fYm5lSgUB5HtpWZxFPdVih2HUomBVncPiuJcYara9+VxnebmGt9mPFeChgHL
2nCO8ToFve4T52K9oneXjyLa0izjwnFz/h9FWR798tvbONGtT3GuR5FusHIg0UVx
EibLXC79fie2mUnNdpfyS3n0+gKY9+prX8ZRwkdZhwjQApCeMsfBIWfmX5qjUNvn
O0B6xr6E3k87o5CK5C4L01GasgwteMPTagVauGF1PKxg1mfhxXJTo+IlEpPMyXoO
G6+mxjKb8avlpDi2c4JDwEYkPZGFzJd/a6Jy7EF0kgbO1Ye9KPtocrDgtl/3IWnz
Ro8+G1/qFsZ+PFZozORjR9LEWoBKzk9zXOXxNa1cG82fKiQFxOKI5eTNo1dd9bCM
DuP3PkaewCP+JSIUiEl3JPdqRlbldnDEhdzrbws+oec=
`protect END_PROTECTED
