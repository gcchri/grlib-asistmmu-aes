`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8bTtJ9M0M4C578xmW+rfBv3dCNXKkTcw+p0n5+HDAYZGLGA0uUB0Ik34fyp2A6ZX
rHLOB/c3pdYatPpoQmmkYoQePce8tPvARaMA3skvPBXtE+GWTmWcriO3hQlSuT0X
UbEnXDP1SgtghYULy3Ij9pZkaDNjDNarNroz++yPshs9MfM863a3jkbCP8Xv7aS0
xCfNcNsyEeKa7eY5N5N7g3oG5EpsAkg2QB89m6FOUl2ASrzTeJ5wJYkCrBbifBoB
N5fagQdi9RCL8b00W2OeFqyFnuige3qukUqOkKb+APn5w817KA2tZo2/0H11K/ee
kcluDiEgD/l0Ui/qqO+SxaEsSq4aE6WYd668GeZVe4XtQiDo58VaYT5Qw+OOzlvQ
o3Q5VWnCM6jvlmZoSY+dyqcnXbDICNJ8dQF5Glbu7uDJlpI2/zg135egksusA/zv
bTQ5PvFdYOBPQhaOhcHIGM/xzImAVc9NqFY9dBWQ7YJlOftpawhhnd27ko/K9sez
OUn9SRrCO9VkKpWfJmc7hRSym/PPSiAtqxYs4qSTVf1I8x+OHNRBs/xrZtc+NHfh
gRUFtmudeaEQF9h3VMfvTrExOeL5AlikbaJZrgP2Uoq+ITBt3uw5hNNhnxO7Ucls
nd6umKsmpkqoPvkq/aRy3EGDPS85vp3UZICzH+wdEcOlEM5kCEv3K82doHfdWFqH
QGSjbGo/Ttyn95ramcjByMjsLY75KQWO+glSoy0yqQiscr3Ep8zIB0t1f/8TrdP6
xysWT07MyuAxn9i/rIbJQL+p91ij9fUHiWwQ40tYr2+FeOTgzkkegNpIvrcso+Zg
4B3GmE5uOvcSUZYPLIph4DOcyB+sou65UlB+o4/CdsTUHN1jKCTiaZOpf3Uy1HyT
Jdc1zZRQBrM2ougjMhnmk3aUQFwj8wug6UfcyMQUm+3aP5rk5CDT78U+Sokt0PEr
MYQeuA6RmvjjY4A49vGJYIVeTVL5n0uZHXSKA8jIP/cKKcvRfiO4Y59RE25buVf2
iHiO371oyVUFfbODVLhSon3aNEwl8faZQ8HLcNJ3VZRyZfRFP7XEDLRsE9l5YP5S
URUGQaaBnu08jzUAhrkAHwFtCmqdPfEop5TOXg1NlyS19N1DuWE0Xjz/TMWedpxt
`protect END_PROTECTED
