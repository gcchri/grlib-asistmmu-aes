`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQpYspGP+oI5EO9BPLHnlnuzmW5vb9PXyMVXlpQnNbqjY1AlW0eTdEFHX2V9Udmf
8X48cCK32TW9wVEus0VyqhTrkqLJe3/ad9n+wz82hLiliNpcMpXwq7qV6/LQ0yxx
gK2ERgo7A6f5MvZl6FaXMo+qfJtY6KmckLtB2HVPpuj1d6Oa4AiYCgUyhQ+mopPq
kNQzmCqaGTeGjYd1CzCbCflaqtyRkhsVaGF7aWquxnvYb6hHJSlEh2e0ULxGJC5S
JsEWRG1s3kwHOns/ZrkhnChF+OqA30Py4sWZqZkKtTX1e7YqCyBAXjajsgMVSVld
cuE6KFYv92J0Gvw107IRbUbY8tkBN6M3gcz3fl3GhJaS6z4bq6kB5mT21L8QvmTa
grThD2OItznUkGn41oEqe1MzUVa4TnLqrZzLdQsuvaGTOtGZeTJ/JWfc+sy2UUvB
`protect END_PROTECTED
