`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rfo4pKOBbLSBSa2FiCFVGNvzCZX3Zz0Pr2T/uKRaruxtdrgwaJizsFhYGyLIloAG
snGm+ubWYRb9IfeAla8ho5FdKD/o5zkUn8aSqvWza779dW0sbcpz8FQrAVmv2OrH
u7bSvmHhfN0TwZ/Lh692UghvmeW3Pce9QRgk79inHDmepTsJ6LHLWYcJzmqa6nGy
b45F0fOtdbnqIWqcLVSJjXm+8XMmaU1WKegF3Ptp6xTiQAW8QbCzmYguPJ0ju+Zi
TOqC2+1vqm4hSRmY78ZlElDg+lWofpVXwSTChGihNWCmR5Phgt95MNyVQvXq5tcF
Xwu+ZCbkLrp0L0ZgNQgVh9j+3oTFR6IVrUs7QTIcDTnnv2E9x2GWmzqr2QFncaDb
bH1QXv2jukIrhZ3Jgwf639XmxrSMoHotsUsxZeM4IN+67dAJhrHy44FDN/o6GjnC
YgiKNjlUapKUeWPpH4GwSEWwDfZgJNynwUc8W9pdTCrbIWUgCSiksERdlB+i09Ra
+t2w6h0pmTaEsK9XcHgW1HE1B33TAR8QM0etI0S8QV3L7MmXtIy9cyofFg9dKVCh
DrD4TO8L9JzjYWzuPbyNVne0WpWlRLqaE0VC2s8e89fWyi8Hpre2Q4AD6pYikiqV
dn97wHN1KH1eOs0yfCU1gix5Dvy/Gh1NLvAjY4HyyLF1QdSJQcvDAmfVhpulep5s
cERRtjy9esrZ/OFn0AxrTagAp05WRr5jY2wKoKeAI5h4uz9NmBB4l01GDuYFKnzh
ilmv5lKGztmBukuxhPzy3W5ZUpPUyYAgb0kHVxvTS334rPf79y0kfIJF7iO/j6PU
ABvR4j4PnhgGDXWiglLbLm8DWSAzKnuWoIls19N19Us=
`protect END_PROTECTED
