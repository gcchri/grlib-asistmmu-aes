`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wsgeF2iSAJzQDMeyYjf99hsAINVWJhSYKWnscEmqpMJZxV/ZBgxNGUmRTPTsCCx
neX+qsQe9/zD2AQLfvXFDHTlBrCegLO/NOT+WR3cwHcDw8m9QJ0PZTKyiPBx/8qu
U8kMEakiOzcUFJSFsI/mRDmmYGx72Ioz1ul/diBcsu7OpLn1KbNeY+VaCdgiVCgd
6qteVDPTuEugrrxW3PPNaZJf/2lPw7+utan/1AN5mUUa7K9A4AgF2ZqPXgbAsZ7l
xqJTIMp64GQNrO5yup/NZ+MN6L2Q0/neQzKk9eUKxyk5xSNfCvsmN+/iUkv2AQUN
QgcOcpqpJFhmJKEN6oxIAu/uDnXk/QAlsxBmRcYh+B0LH0JGY2mSbjI77H5ymnoK
D8H+UI8+ezH3KG99QHlF+bxT7pqQMPQ/a3dA4ZAvSIQ+K1uvFHYBmbhpMBOGeEd3
fcmM4lIbwYjTJZi1tWW90LTzoBpBTJcLp0gvfFpuU4Y9nAFRyc26MtQ6sdOzDfHX
3KMCJ3VjuA8iVzsIaF12yx4sjti6BWbzHSu4qpxrxlSceKQ2P9i8XiCwq+uwcTek
/U7t56P3wRngg8ym9ehMCDrXDa5o9wz6JbKnzodyk6EA3rZ0nlCV7fECGz53kfVW
SxTsRqiCq0tR0Ls/znqPc1VvfoKLy/fPW2bdF19Q1VtsEEr0QyO/4GtP3E9StNhX
XFpSsFAfw7u0n9wJfShVv3O8K65dtmjBe2tPFsXQBpmSc3w2rfNF2XRtdAjaAEqy
qGLvKRbZm5IRcOcL55F/Iytn3yTjSsEFlAROlgZ/wd4zhTHNkFq1mOF/2vcpIVd0
T0YKtebk/JGEbWcihJYMC+Gl9Kj7N3TrDhbIxIB1hNeIoow14XJXG2iqcUafv96S
6dDVccq06Qy+afKyniVjzE693VZEgUIsKjgU+MYoOiynpgSyttsSSTRWLvUcMloo
FlRsPFGXFvSaU+IbJOLzVNCqj25/DXeICye+1cUqw2rx9Q/S97udn1s31Js+XKRc
0zVuUHe21cuU8nEuS7uBZtfYV4YjM54ptIF5WAgyBb0OOs43D+bAv8U/3oGXN3lG
gjrVLGf0XaaJ9MC2OZECdQ==
`protect END_PROTECTED
