`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJ/Rn8u8sU08+yPFCLJ2fabn9APni2ZUQ2Wq1R5JDtWnA3Dcqj37ErHrem0QBMmB
nFCel/LeKzGZmol01Sk2V5z4upKW5CGWFyORhzpq0yMTXPiDEVeQd/cd4g4DxgsN
VBT2Zi4/EEZ5uZ0tWdEEdHieQSyebzqhYLGP4LOQZN343FHJh+JfBJgHpbGLedWE
/UDW9PIA9kYqhVvQDgcXAPmk3PtvSM62ll9jqY/byYzpNSMNonkF1BzFOZXpZ2rR
BQOCp4Dmxfkh9TFVW5TPXcBlzzTj2wIQQN736EowCzGnVyG4Xvknx8S7QDHe8jyP
WX5EbsSb1pmUoX5HkqxD3YQ2fMrM5PNucSsuA5kiMPENt6OOKgQxKjsQQZaKB5YL
An2OAwEnYsLsyjfpBPwTC/1+UKIBpEJYqoC7iRwCe+HWGVwPHxUOY9y/X5jTW9cE
iQ78g0JJT3LjzBc+32VEItuyo03G5DrSjzZdmuI8789zXqdfgoVCELJMf5jGfOEa
5vBz1vfJvru/xrlMpcNCDeujgjOHs3G1Oc1ShuGN3BsaDa4B2rJG4+AwyrvHOTM+
t7mu+wwKj5GVtMDiNklRO8KwiOKMjJIEgnSnm88qZVam2/f2CgO+ab3qdlVAOl0T
zCSzR1g7dhbLLoos6N+SDJosEUrIXjgD1WZWbia/A3dmpfk4TrBlE7o+zbfEpJSP
/gZ9bUibsiSPlWkwgHPzGiS1u2ciDWzPXm/Kv76cNrGbSlj6Of/R122pOnE6WvYk
lB6E3bz7Mlpuxmm6mpJx1Btpoi0B9ePJiI//IOK7++kdtCeyTTBB3rVCjrqLQk4q
vnXCyxQyMQ20BhRMSLuNoeIWEspY5B4CN5gnLCjNgsXCM6oqezlckI24iMoPRalG
VQgflf0KsuttJvl6sbRcYOXUgC5pCLo8jm1igaJh5c35KbpnFMleRVTre4q8tUw0
ffDSxgauRi54W+zJd6azackdUwuK26Pg59iNtV0G0kw3Bx5S9JIlVmAuYxk/+l/X
Yrgjf4/l9HXU1UDFwhvWIn8c3S/HbipMkBezR+NVtWNnxgrQsWR16DntBgktMASJ
O1vqTfZhU73pvk1v6r0c19xhfqt8qH4rusjddXN1yaXpwqND8TGGqKAdEQ9DkB3B
uQHjwJPJEdFNlfiuPpIUn81NHCdxXm+v6AGd/x075OLYzZp0+r+u3uE3vq2msI9d
5IgHi9PHt8IVLYu2ZUxb3hVjbQNognmkjEWuYhQqmBepp/WRFKpSm9OrIgrDhLk/
DI0yeMkjss7s6XI+7H6wNRTLmJLMW83CmGrrXiyFc2dSH8ZXuXOIbRb+iwvvvUHL
5/CTigd/qNAsK8QAOqi6kNjXXZE7E1SI3/6oy5bvMQEJmKMZMLYg9RyYD0JwfR8V
BFtf5aB3Upjw9RDLELkpKo9mYWCu1oByjOrBQAqrwTY7Cs3g/7E5uvMAHZL6vl1b
L/5MFuWb/o11JaTvAGPl7kykBhD7CkEr0PQh6+P25yTEgxGmFOSPBUVbHj0CpyAD
Ip8uRGq8I6HePda2iW33nFu53i4Ti68fw2TXqJQjYGI+YFyFBMmhjwB8KZWG5wjm
hISpxVhHe5sDZshqkSioHA+wppV+w2WjYoot6E4oDQ5IojNg4FzEWBbst93BrvW9
hsO6KQkE1HN9pusGC7j8o6VwPobSBNmDCv4jsNh2Ef3HusiJ7c9PBmpiXIXikBjp
mVxAcaQOEsj/gTO32Dgsygcoid/dQ7clZPO8wKn7NVQ1rT1l0w47ny6MS+mcrK7o
QmfojxTrAA2y31UUKMe+MiS7SY57TLsJsbffkHQPrTe1wsnZOkKNtkSGoj9qz4Pe
77aPmhPvwK4X2ohbMK/TQ9Ytxlf9KLUno9Go1XC+rU5HTbVDqNaJsxwOf+jooAVs
MweHSBDOIhcL6izlCthbdyTGMl8e3/BaUddcPymn5JDrlmrAySj0/ulBLG/tDxh4
oa7D1g476YdBgvIhLH4X+hfCvbADm1Ndaket0BJLkU35kTOV6G0/HPjB+Kv1k0k6
RZBjyxnxXtXGLptw3CHtSuid7T6Al8XiPF0q2IPj97sH/bweXhZ0VbTMQM6piBlj
/SKkdQqTEPym5n6KAlgY7bOj4kOAZ7R7sfw6wNfChpRdcTExBe3WALgUofcxOzdN
pMk2ezdJIC+ZPt8voLyE8mGYxnx5oztd/ZJTf8VNay1qjgqSmKZvNctwocLXU3Zl
YCuhpoZs1Zik/97KTvoYcV7E+oa0b3JL9dJN3PdaR7eI7VGCIMrpbJo+zxBHKSCq
nAvhWGwNhlcjX+0d1yKfKapJmJVoG1Z18a70Tg0ZLj15W1MORdRS85GUCYvbNprt
erpQAup4ODOlVuweid0qVwfAYW0Khfcj2p0W4l5kuF9ul9fwoM/g6cypCeCSQZaR
P2oG8IExtIEH0dsktaFQ8uRp1MUQxEmIOBgYIBSYKZ2cqpaMZ+xRrz4kvz20Wz6D
Kk7pTT+IHav3oe9K8sBR1OQVA797ohjbnQG0VGh+LyKV8Q19Y6zdEpOqxvb6M/ad
cAP1hJs/ccv7EnZwpRfciBiXiPrM4hoGVFJBHn8gV6u+L3JG6CakPW3gw/U7l7be
zzXsO52l7H6tmhVqdqitEUmgOJF9NVzRITIU5IGCc1qvqfvaBicgncFg4ho7FWUt
d3aZrxB2cAatDfAJGd9tx3jgLyuW7on2fIG8a0fOPtr5cITQ0vXGCkUbGKyGInm3
a19/kePBST0q7VMzYmixwTdMtRxstMJy+IyxnJzo9uT2/ZjcS4po5yB9w/E/tmkV
ZSQ02OU3BZ17zp+V2djh/GKC4516JgD/h861j1Xh2gc45YWb/921gtkEXFTdiJkF
oKPsMnV+ycmo8lqkZK7DXvYHtMlGsc4ZoNGTrj/vqyt0diNuxIWtMqpnemB452WX
finFwqYnL86fcl2bM5LYkXSr+9oN8JEC1Hk4+rfnTgvs4Rxzb0/KbKfbupalI6BQ
CYNpxn5lw3w5VuRXOIcxO9DBqhgXZ733gKY4I7YMjZUV9dqwg6NA+bA83gr21nxh
sbZ46lyJGISaNnBELyRP0+E+mtLvT169ToXcRI4bVl2YnDRJ6JdrCk2ng+4FQUcn
MGxKAkuDg8S1JpSYcegEdFqTQd8VGHQG+hZTROCFCkinG+32HZlw8AwnHqKtXlZS
Iyde38S/AU4Y7ViFy+0Ipdf2ZyZkpf3BGqYYobWNa6AvT3LQJRsY/mTj88Z0t4IM
dQi3iWzMlsdDpdD9iD7B4QYBpDkI724QvGkbyk3tnx/SnguaPjnZ6Uh3mh+bCW5z
L7u6/x0y1nvGArkCBxgEYiPyvOOB+AfCSFQ9ip3RWX1TX/4D6rNTNDCPqA9jlN4U
8WYikOoGirmJCn+p5eTaf0Am8h9mXeXLD48CiHX57AN8JzJaWxVX8CWWb1nVayAe
jUuBS1NP/97DwkRvITB3IP5da7dMcgrCGuzi4fmqp18+D/n6UunH3b7lyMSqPL99
4cPKr1P58FV5QgIMoXMbMMrSQazPCMMxWJYu8iOkj0hVauXAuMPW85IlGvOaTsuL
cAsU13JhJeBPm9E/hI0VsMyOfWjpSVDO2+CIK6e7Ka4xWo7hVuyHy26hIKO/cLmv
fbo45gfj5nBlFKdBlu/hqPFA4d/2iiM/ut1R5oMxsB6CjnHtnzgWGIhjDqAEmuOr
a9tQNGhmmQfkwvs+DI48vkl96mgPq9OFdoST85+s7x3Iwoo5LDp3m4rKvaJhxRrw
zRtnydDOAdrxLWid0nAeyGDDgIpE596eZftEqfaG1elUU1RPrrScYid5qi2e9fAh
I7Q5xWARxfWO4jVQ6PSQgKowHTLOYBx1USESTpyQfHGi8g2HVwnkJkclf6Io3ZvA
KwDeNPzsP38N9HqH8VpzBZ0mvn794lplgiTRXVtaUZq+oPTZna0TXRXtn2naZvLD
Z5nEMfg2pIIEdF9D/Z+XKoa19ZQf/g7sMWOhvTcMjeMtAwe/iKbR/o7PjiM/5ND2
XkNXkGNvYYSU9VZfDBWRTlILMyTrDnUb4b5iho33jmbiVWdciVX1eqOKQv8DD6N8
6Bs1MndF/kYigIRLD66PvQtBNT8nIkeiaLdaoARyNWIExULssLzvgJWcZt0wy4Iw
irDtcRp9KvO3DKZ4BuwY8WrPfEMtCTZMAMlRIhMhuwgsnqNO33zB7Imj0vNt5dQL
yJv5WjUfUl60Wip+4b7WeYo7BnIxtOIw+Nb8RTm2FJaheYvqFA93rau/IPcwqmg+
1Kkqk/3DdUF8xmCnesipa5juFakOz5RlLaaed0BduFSO7ydeGZodMzjqmRsyTvHg
msq8E10dpFQnhSeu8bOjv08CadvfX4fZ4McmYi9LrL+XvTQAx/JsCFhT1skTAflE
2z3KaDPmKEipmV4Tmtm+LiIJSOTa+cQN1wvg5Pt0FGqqj2yvYWBrcBLW38Vvr6JQ
TEkhuNWfpFXA+OYsdbx9yH+YUsdihNkeiMdNLUzNsESFaooTPV4sWQfmdr8l7Pn8
6vL5pPvKGQpCSJXGIlftOyNtsbgS65EaHeI3TKzjCmBH3P9m6rmaMB42dvxY4r6i
TJtg3OexodyUfRfNruXUq6a0mVyoW5N13eQuZpMQKxCvBk9EZYs8mo5P7IZtKNtI
VK2iUpOjSPaZd45Glm4dRr399Jk4YOS4rokXQCGgrabwKc/tYKG8g9+atOhNWvIs
ZFbgSDGQ+48e574vtV7Lfj9FG1pte5zu9qXyNF4wi5FGumpAsxBRIueesWRhtSBM
AvxwKRvqgIqAZQRHjt9XnzrTVErGh06RWKBO29fDqADYwMG6+MbTkx5kfrn5ZstG
yDdbVgiRXgCgzV6bqA72NcNHa8PyEM9645I1vtyzttdwS3KNI3Ss0aiVwTxCUMvv
MUFuVhl/vNLJSrUiRXJvQBJkzSJS9/ghXB7+Wo6XIVhZ4zAfcUdJ0MIQGp94d2dw
TYbiJglO20d404c0ewIjSFbnyTZbat4adRfmDvO8j9qrZoObCmGevXmXH9vAPEaz
0ZsNhFkTBj0FA7fZczTCEX+LY4sdaUDMIyghxDcoYOpQo78t7H3D8ia3uhqAxhHO
PNBgJjd5W2071Bk8S4DwvTyYHcIQGzuiv3Oyoq8BTXdBosbq2bW96/0tK97Zlgkl
UYLFRM1Lze9OeygmGL8OUwBlI5UPtl+2jnOCQ33KYobxFUnPmEetbyTnrvsET71e
Uz701V1+Q1V9odeTQrkmlMJf3BRyHuIVhp/PgCTkelfe83lGlfKp91UFJkedYiUf
flV8aVemxcaATTLdDExysnyqalOOCXhoUpqRCjBMUwmE1vy5xQviGClDryx44Yrd
5Y/VSZSDL4tyjVkdXHxy2czrOKxw2/2zbZ5B0vbMGPYwcaGjXC8w7Zrez4Y+37XK
yjZix1rhnKS0dVrSf0pKMdw6CrSvspOOXn2aFxjgiLK5l5X/fQzBNrPwu1KK7p2U
N4oOwjH1H06Zj5WRseTS5sH1XsZAyE6+z8zTqUMlcXdKklHmI8jmzsOQqHK4VAt+
ZNdI+O7rUcSaTBwHyTHze+xJSSsTP66ooNNe6Rn1Zv1mymIAZZdLeTzvUlgVbgU2
WDfB77FDbmTVgWCa9tuZLtlNAR+0oiIP3djR5HGfKKq8E1WoNT5DkgFqH9KF0R7C
GVBM4So3G+G90dDeN4T0Hy9tYivV1IAmZvP7+uhuwAx0ARKQfATZfv9g99kJCvPD
klR9YkFrd0gYZZuoC7WQvcMKv6A0vfRzE52E83UzFdhaI2iK5WttCOAUDkzE57TZ
Q+BTOlaQlc2Stn5zxq+YdceyFLu7hNFr8mudM8lCkQhigzyEOnmRMwVmznBKPE2l
v4IlvdH/UyUNjo7GljtGrfixmZilndIOTldTYbJ3r2vAl9d67iwWYhrh4mPYu4BF
yAEjhhOfq3/xruyHCfVBxN2alBht26lrmOnM2rAGwrw=
`protect END_PROTECTED
