`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXx4k2Dj9WQOcr/6NHnEVXMhnDo+A8ky3qCEvW96Sc9XA52kSu8/n5djiLjjyExD
bI6eyBGK1xK7j3lv18wLQsRu01GAGASasYn/r0Fz/xkOS9ShYlm4Ylc8Q4NUCAnm
cIvcx5TecmaLdP8AP/oRlWr3/prczpEkzni43L16Y6amDnpvEBhda/IrnouwTwWN
JFJmGUw+lpoLWgNro6fyZ+Frpa084ELOxgYuPPldNO7bp8oHNaSPB0edXHC06rib
+JfgZbk25n1qpeaOeHUSElEsr+iNtkj70RxKDt3GTbDuiFUkkDZdcnf+6CgA3Oey
M7CKHjEXG0vEaLIZytOffteM/nv/2PRmG/csyhXnOX6qz00nwo+wIAOU0FkyYDh4
`protect END_PROTECTED
