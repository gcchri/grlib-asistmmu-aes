`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlka5tRsy5BBuwdgaFuX3EcsFKfCMmlHnyuHPatvmNd1RsP5MAkTYiFF9Fju0wpM
QZ/LecQx233j/jjv/Jwi0xOQVxvUdEU43d5wUTDY4idoA/xJIUcIu808WVyOv0e2
dLp/5gT6tl+8VEccp8oj7ZqHDYPMPb7Bhfdj3UFbEs6Ea3HCfwSMnxu0B+tHuTZG
zu6iTDdJAiHOvsCpy0ZtgZ776vqnRkhS6T7hk3U//sXi91mpQ7iPimbgCHB6pbv7
khAJUe/VFN8sEvnT1G5SHsE4pNhccHRuYaQGNMdJ2XhlQ7y5l7Qu/JWSTwoD1O9V
ObExCPYd2HRs4LbUMXIHWo7vJtunIw7DNr3lHCyGMu3ztWV1cx/d/b/RHEwxi8Aj
/2ejlHts4dytMQM2CiLQxfZ72qLCFHdLkTvKXBWoluwRqc4wilIw5ExX8jayv7ES
9xpSJGLKeLnnIZL/ZuM+i1ilfE5+dJIib/mgnd3n4liUX2o1W4JedkSZwv5lfa1G
oundFuGYlqRI1g8btxzWRugFolvXT09qWl6RjPHvjSsNTS9LjxLzsmS6E6ExucdW
/HEM8r+FxpcRExC8owQlsSEbwbgri+2tAnfHCps7aum6vWC/ZVR6+lEBWFAovj97
5qFPR1Yqw3XaIn0ObCyUzC/7okE03IdfafxE9Pi/JXj4YR47d/kTuvts6jo9jFrJ
8FZ9Cc437eCUPYVsy37lGIe7PMauPN4khqgQPSgC7nHtuko0pUg8QNy5g3Eb1HGK
PNhJ0LdLG+ydMGgp8/vZa00ve6ULaKV+kOjPDHmoX3GhAeaoMcmjOg/K/+I66dac
jxEak/vsBcM9zcL/fW2gt/rBJwgFzPm3lc1tOLktY2heH9GMYhSSb1K4pP4WBoy3
Lowc0EE1NTLMe3+ucRTlM4HPAXTZeAP1p0MPlcNckQqIPFR7Sz5lWQT02cKaxp7z
`protect END_PROTECTED
