`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VuOsnSdiptACfx80aC3glFPZ0RTt9qsIVmmRt4JUNyMpc8ZaiSH0eLLT6+jpEAJM
wWo2crcaDjL4DKugMQ2nMonykgZh91uFsmCflWWXy4cn5OjRmIhtRhJbhTHxAtpl
lULLN3ZiV74AUm/srrKf1yI/g6rIAJIT+S7dyVUGJkbrmwEIxTdTioKSuyujW+8P
shpAM/6p+EZHzcUKjxwHZmK9I4JKFm8Hyvr6zGuAMOy77E1FHoq4DbdRcQwPXOoc
m6SVzq8mySxI00yGoTY3WAWRQYiWNCMkmj5BVSyVAulIKJ/nOCbttzlrBYuglVZ1
V71CeRpyjozzJH4hDKbHCu2k1X4HgAhLIM3Kbvo37dv4qX4DkbzFkPuLHS/UVH3f
jlAlNKNhp7plKlhYawxnd9LZsjyvb1bWIAkFC1bVMFTyppeIjl0rrFLF1lSCvgUe
zrf2UtvlS62Xrmm35XChYjSXvfCfOsoUP8iNgy4s46mfB7sQwd0tvhhYC1UFWe9K
EuE9n7QNIN2AbGe1c3tYqk2q8jltEwEbv8vThHE2ZbAS67hsRJOhsiXFNaFpxBYk
XsmTvOhxRdpysstu1GKwh7gbHioI1IhuZfjAkeEc1GGaLfyV3URyhdIboeTJL+t2
9fzTplmhSKf6ppcRI+KcuGnXSjIhdmxd+dszH2Q6a75kNW9p19AwDrzlnAZ0gEP/
hmKQQUpoEYyU8lwApglzvxnfg6uWo0rR+uz1nBxiODlPzoJoB7INwdr/+fbhjXlo
HBl/YzE4yua/Xv0RRfetjhfAa05Er0DqA9YFMwF7PgGinGHQUlxPhQVr0HIwhHXd
`protect END_PROTECTED
