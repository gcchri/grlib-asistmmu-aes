`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sLGBj0YIN/eVMAzrsSjdjt+RZkLSSMxwoUsDdV+nn8uwn6VLEKUVoG7DYyAAwdYE
vASfr5SGifBk8fe+k32d10/Sm5HVwv56bPD9x1OojzgCDFXeu26e4gfp7dPaK1rt
5JjhCLbL0J/fT8H3BItpuN7W6kLRk0FA9cyRC1prNc3rDeKAUP/dbdJ2HYFt34Sw
/bG25KmcXveZyvWTI5mulsQ+etNZrJK5RpwkVqAcN1c0LfZPAhMV+4mRCWhy3l6k
0hT20oo8W7T+p+W+MVv6S1id8q26PMQCuHfi5ffaKGj5i0coUXWgM8/YPwOUOU0s
tmpXLmijd+VO9A/KkdvZOKjYv0ni5Tvm+p4/Xhy6/yddB1ygHqCd0Ph9fdG5wjBW
O67R5/cG15RY3b+S0z39C12G6mZZLHrJfzTqvHvUwI4KL3qWzJ0xVA7SlZytQv0Q
4q+ba/MwGLt1GB+X1qkfGebwbVoQFeiZrRleL2lWeEV5vsIloDpZ7t2BEaVeBcDX
TIXXK7IGlorBJhXE6QcROGKCg1b1nmVthTks+qR3t0/yY/R6Fw/caiaGe1rvhsDq
sPf9TW2EI639QYiFYagjqcncjD6y95qnR23OlJaVXPX0c+qTrCmwmBf0djyt7dMR
aZPo1LkSjZ5C57RL+YYgWf+jiR4Crx2P4ojKBRJaVccMjFksocfbZZIrteErC1uM
ZhtCkiLpVTgKL5ElHA9QBrUDVT0zp4qNU4uIkzRjGVCTbgMxZN9Tb3hi/Ir1P8xE
2GcuLwZ6g32jqBLZ0yYe/9t5PvVa0lbnh8iXrWz7Yp2lrQu8Hohr5fI/PHw3Qi6X
iLpB5ApuLIJ49itvDVGriw/VpqCgTLkeuJa7RVMahg07NpaptuEwWvNm3lBpX31v
x217CGGzSUcnQMuGVxBKKr6a1DDCdBnX3tEshFuZrUnUZ91NaJG/DeOqspiU4dmz
V1vARUI/2vIIkEf/lUxX07V/fvdulId3SVbXnTSKahrDP0utneZRSLC6fvo2NZnn
eKPNHo/QYbVHQR4E/5QVDtYgEP9ahG41KuFZgiHza/b7FcqEAHOpy7PuEi5py0ie
x1MiEbOQzcLXMW2XsoYQwzWkJvzP+DI+VsCuxub4c5OvyByzkFdHB6Ckr9EFbIGi
6B6aHvxwT4TbH/i0DbgSdJLhBQULiXTZ0LVOYuDgxwiC8+DQYQO5ttGQFL5gx8g9
wYPzzt3Lrp1P4Vzo/RxaMPRynycVXQk0/oSLaIFrlNpckymr2f/b2SaIYKEc7SB7
gtQYkJcpOz4v/WplD/MadQuFeeDcZAXJEnhff4BuAMiSc9R6Bu51P5M4w0yrhGFJ
IdgbTSFodDWKRvxFVtwHalmu5iPpsTlvlOzVQVu43sPjnE7ng65i5N+20gPXPznO
pENvEXzzbePkNVNmUDShNhnplBqwhmsptKtI7T250eFyf9jjBy/jwW4yCsDQY0Uv
y+xaRMj0BzvpKg8lbLMwRDWYqZ4kdxeqCvfrOlegg9KHdvUYI3yLdX0bWLrQ1y8K
MXUIwR54JFabAM7MrM9hmXmnxqWeMuMVIbxZZ6lI8f8f+Bf7dRS/iCOxVIKorQXe
v9Esirq401goUzJpVaWk3s/CJ9DLlTa2i5mTbd5GkuVjFF0zEukfOJW5Hx1cGSyS
NZ/0jpJBaQbEq4Q+M+034TNi5smN73eVQVP8CtDN3rDeQuQYbvU8qUsVQlFhOf3O
TJqHA18zDyF18AOrkK8sc0TLN1ghMoKymrufUMBQNr7tFt+Ye6e8vkTW5AXxWEtP
G97mmxcBMKqQrpxAhfLFgnyZEcGaXFonkCJ8x8daZIwuyoglWq6yGhbGXrVfhYcr
JYcmHcsuK1Sd8EpAQtNnIFJ6uKrVJSCRtFJGz/rfhW4/CuqezHNYBG9gMJwd9bOW
i6QJjFQvl6BqywQYjRbJI+r4dT1nco26FAng8A9PCU8qpApWKMa8PCDe+RM8Bq6n
r1IkknzrdaM97NP2opaSv4ILKcFxG0Q3PIE+8isw/khL1SRJukf1OCTbCvsaHBWM
pB8dvMP1xi/cJ4rhnO2gFkF/soCF0Ac5zR1UQfWfPntstxRGJolhYwStjLZaIh8+
afkSL3YLwq+ARE/qUWEt6FOuOC5UV4pzJOz/j9gSX3p0CjPHDSuUAClLF79QwML9
BT3bvkFoSkc/ZFD0PxtEbJFQfQZLwUNCohTfbaMrG0nRwZtRd1xLUmr/9+tAfltk
CsSdFkJvsJY8kX8+cBiOS1PbpU8WE8ygoMaPue+fNl6fBN7bP3z4FyH7hBuehXt+
zINuBZJJrFHUhLhZ2XvP9szUDOAF9sHgJ+xi4Cn6mhcbN1GR++x/0W/SPjROXKg1
KURrNiquclrx3TWfxZiVrmrBCVGo5Rxb8YbfF1zCT6SKOPutd/qGzTfbk+8XSOha
sK0bjBPe/npPm0wuH8oBvnUvSouxGQWbLiSarHE8lPVVVMHSBYfz/mJetN/sZWDs
y0Uk9lk3YS5zXyNr+OSm3MqZwd/1E9hyKh9k83ytjeQY+4yLIGDnW5wJMJJKQkl6
Q8XlbtBsqkvVxpG8/BDKFwbdEV5wezkWfUVmop2e+nlKjp3rnknVByx2P+p5oRNr
0IIBPXaiKlRyQJde/FJOWb7yJ0EBWhrtGVFCvnWlSZY8c5glJqboc3NKFtTY7sjv
i5tFxT3LQySS66DH2kNfHM/FvgCeuksR9pgX/rydHgICpz7ofbFYQ20p20ej6Q0n
4PJX5OB/M02J42bAZqPmm4SFm3UDjpexotL1KdKlG9c=
`protect END_PROTECTED
