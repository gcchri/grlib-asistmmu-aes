`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3OilwxuUc4jHqn50WE+Z/kt1a3Q6n2eLVM6ChB9VsIWt8S0KjsBLSaR6RO9QOrC
z5UMtJCtBlcMVMuS7wVHcOt5oY8Ba9U9whmy4Ha1U18UAEvRi/lHAB1ZwNZwjmJc
/pubdUWBW08RUV11j/3k5hpjWLJfPWKgU6QldGNzaYqfrpxudFjLpPYEvtb3asow
Czu9oXcl5J4vxUarHW1OJO1Lk6eXyJnqRT6x/C4fgDrcE7JQaOcqY9VHUunn+hlw
chbK5KplKixf2/hIFCdHnF0dWW7Mcg58v7rCRlfYd0ciGXmYXwfa+EmkCV968GST
jLt4x8HvAu66rllp9ZdbsWavwMr0HzbviWFDTqujrCe+qUSNTCDrxsZNY1z6B4hm
fsdUer1ACOZflRYv//zI6uxRHZH4zo/DTwo4sAPKWwsWhOAYAEbDfNsd9YvY5ti5
2mYlhO7UlVcXPG0TX9kYE/QbTBQaRCOKFPc+ee5W9Hm2/BM+N6FXBSnpPMoyeYDY
692eSwuMNAnA+HSUQEnSKl9dPOcK1R9MyyaCSZLuZD2X/pXsquvoYpWCQpg5Hx0N
`protect END_PROTECTED
