`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7ijgozmGfizjxlXdLM6V4TRR4pLwZbuB1EHaD56/6rXeOenOTtDyWl7byVqJfW6
ZOLtFT9lKYuJrtK411B3yzdDAG2E+Y9Rdch1joMu91KmeVDXOwjKpnBKILn5BHSE
Q+yvx4givnCwI9rt+pLd2C3+yQgDCXK8AShysF5dtShtW31D5dXNLpJQ2nBVRvzK
2lkyaI2qQ2YOmNNNDQGlpol5OWDU+VcIzLuxJCIBvyMJryb32IBOj/wKz+EXkZTw
wDJ+afHQVOpebNaFttiXE4mClSVCDAAluq2o3dKnB1l0FH7tzt7MCnBek/KNKXrs
++xipp4j3S+2XGyOY8lPTxh4hk8hVhIUvZrVEQ3sWPUzSS03uGGfVA0UkjNECZLQ
zIkiS7kBx8P61Be3YvTPCSuc682lUtT1NcY2JxwVpq7ELzfWOaZvc4TtRMCVrpep
gJDIEMhBzWfsUwQV02isCk/8v9V7nt/70JBnX0/fKL+nqTHXngGBqHhAs8yrxG10
BLKNfxptYOh2xRrySTrTWTRFQpJGbDfPOQ7Llg588QikQI7cURnENwY0yOiujXW5
GPHeKvew9vqStEu0dzk47YQPGCcF94HQIJVDsh1s3MzovzdMFezDVR3EMfb+UUoD
wUfSalDT9qNbP+qBF/NLVdRSttP4z2ArHnO1AS1ml3k4C/aicC+eBuAzK3nsjvAM
/HHgDmZiXyQYJ/axJnPSRUkUjj95AZwTYI4xhHQkaX7wHCAv0VAv098kI/fLOeJp
3Hqn6WSE78z/FL1Q9OHQFB36DyzRAa3e7R6bngjDS8fQLiCUaVqZCE5z/5Ie/FDZ
BRYwlnJ9Ihe9PQf9zbF+OOwOYMonvIaTefmrEnDvTasspBibRLpogK2Lrh0qrpjL
n6jkiAsFgHR/sfN/y0u7lwT4fmrqR2eAKPZZyh8jFMwPbifUmCs1MpOGaoSw4oYk
l5p3ND4e71Mt/T6DmajZ2Q0W5t66n1Bcr+8o1pF0wm40O0b+oRnbyyLRBR2h7wil
+kaXrIzikht6B4w7ShNlHdLjGmWDWNJrVlWxVZ+rmf3Cnevy9yCQH4ZNeOcddcsN
ZrddYrtzDzdk0piIWWKM39mTy+uZB6A/Wc5Yde7jgC9+ehATc8rNWRZb531Oc3td
vOu+dSaUK0fubzOeazDmTGTc5Qbq8tlfUrDzzjPzCUCm03/gRVaWWkzXpPMjL2/4
8rKZXAn9HFpgrlVZQd7Hhosz+znmzDRtPwixVvPGz/kQPuH1/oQ7AZA2cN/HZiEa
nC+nzqtitiTJInHqGjc16lhqRHMIIWwPKqBuKEHLBGESrRvFv5A/xTjxmS7zs49e
UDFIOi5F9AxED7kGEHnIE1+Uc4/Ya+KwPOqepCHj0piMAlZqHbY1p9DT/1Qm7xQ+
/lvBl90y9kRHJJ04grhcmVrRYFgwnRCeuF2aHxmGie6B0osaKrVCcSiKPXxYUpkg
/JkB0wzywrM2bBO0AbdcYJyBuYFO8WRZlJkdH5YEZiNAP4hLVjDFq1Engj4blJUR
uA9G+XS2wu1s3qKa1fv3YvZ4/rPx3soL5qtULDQWWvD8rZP+OArAzDoX61BEw7Eq
tP08eV0xvWUVQfXuCXwXpemZitUCcSBaV8CdwCYf7OEwMNeTKqZslaQNXGWURtWp
9X13OHEVv3VXpTNz8WE3OYW2RrwsKTdgwYurwiYBeigCWcYAALVwS6V09s426cqB
KB24d3AFsw6jOZ9J20ur+buBCFDedMS52KEl8wY2YLo7ZcxeL5ZJdPKoPWw+9M16
xNQeCuib3ZTV65OjrQAr5sHZUKXO0ExbHES554IBZxppL+jJzsRLPGo1RnnwzSpg
F5pYpaJd15PBgjP607p4ga3y5bkAgdyrGaM9cG3g+eUQn+j18CP+V3PReyeFjoUX
dKmZkd9WARkpeiP2aAf0v6z6dsjitDQYsb8WYeG8Qm5iELjz9+qndGxqA2N3NhcK
Myw8WeH0R6EKoMbA4QCo5d25LOvqAKk0h/faiDMdzkZCxyaHmFeni6Ayw+BG6TMI
xCFMJJ8EWtZbYnpq/0t3F6tQHyZzK1SI453mxil2oJkB5/HLTNyM4Tp1m4zfEHF+
8Th/31WvT6ydMrfw150vWtPcZkXWclEBzTsqIOVVxAfKb+2y/eLLoPPoegyRCpcs
wt8gbH3jEFB2jBKe4GnPc+wyqB3njwuwzfU1jAixHr2hK6bAtZTz+JzpexvvAXyS
06AX3BY5FgZ7laa+MbiQeFViId6JbPLr5OLgJf7HYUQu5Fxm+SDuqkpqRcbZqhRa
pUVSh63EXDZIlqNulFCi8Vvvi/cMDi4k0QiDk1WXDqHnHDEJ5AgvBcOrlX0DRhvh
Mvjor4kKG4/4lsS+pgFUZ/+YiDPp881UECjHNgRqxDYjqA7gQlDT/QtCo1eYXANe
884SQyUoTeINeL77nHYgMUHJMYPjde9GFkZuXNHEL/GhIkQtcqC83oszKXEgGhsw
n03amwkvRy3lpPBcrSmMxbL2GMjfVJQkNgTRaL7bUP0mYIWw9yUYu198e+OwSbSj
xNX668fie8Wy0SQqp2jrgSHaxB6TuCkk7vIIIgwS3FDkBgwOKKoph3M9AY7xitU8
chdePh/S1fdOz0yV0IK7qfNKhz/tu7mQ8qk4oq+eixeTnzuxD/hObQ5A1QWYtlh8
y4QfOjQGbZHwijcxLtcTPpqqb9P5aNiYe+o89uHInm9e+GA9YIF6Mi8p4La8ARuX
Gek7nxTIZPeZMgkF35YlecVQ7s7kMYWB5hHzt9jBjdmb6UzeURIokp1jPyb0UB/m
32PU5dEiAc56D4x14gkjeYVSNI11IA0Caujjurl/s7yVsqD7cJ0/D+1Us+o6xbHe
6SiFommn4SOBKwc3kkcEwt0Cy1WtIm3vDudCDyTkRB9mDfwXljrRsLs9h8lcOPqF
d59iNVOJJMqvc/V4BotubbYHnkNCdazuKN/rOHVagbNRFhPc2l6CsqGudq5YMA9O
gQV9Os92WbbUcjLRbnRtjCz6g06dKbrXCi1buS20GB/86AlOrqY2onb3lMwIVjX2
GmzSpwqx2YSO88OSaTEbS2nNwAv6dmAYivSLaSJ5lZA3u3xwzB97dxHwn0JyRXak
huViFSMl7WtBkNCZZIc9uBfppM8g39+WAGoaFkk9PSAHat07cK2iS9/9HOivRmed
esi0qynuJTgKDhGu60MyUvgH5Z+Jj1S3iWevvJtT2tmI9UVmxl1DVs+ekzGdQw/f
1eF+S6U5lAu7fUTr18u4/5lWVrGF3icVXWRH0bfeiBALh/hav+NqzBBIpQwSwAiE
5aTB40lkCsxIzuwkUtH8lz+zzGNU6aOpysFnOuvg+aBEyWYhdK3RXHXdSetKlBpc
SgEGmNf7tI3H3BKVBoPGv7GynnUGSlE3RHaBGFOwjyDebltpfluGHLc7bkfGItHi
lXzERce8AgWwuZsz1aq5yUJczx34eWiUc47k7jPAUVt93RWMIIKGg421BdnVKXPM
DHUQGpjHRqopdYCqnYgSvtVkQlFgouiovx84Ez8Cqho6Gsdg14GBPYl1PVzRY0HW
97eeMUUHLeoz2IedqSXhQANJRmz4fMtq9lZ0oXb/cazRIUcg0A9MwNgO2Fnx4aor
jgrhayyajd1WWXSQfZpdOpHyzZRlSSKJJ+Qj40JzNSLn64v1bouCunddkI+UeeJB
xlWDfa4b1xUEZkCNcIQtDamBxZQq76nvb8QVs4KfO4NBfG0Aip5oPyQPSJN9A2ws
f+KqU0NY4WfT2s3SOSje1n8enQ+c3U7oWJPNywFAAbdlZmhxD5BKHqMKNyMXW2QF
ip0wL3oivtp2u35YvOsgeuVo8Uze6gFlhGya4kdydU6D2Ze1I2yFzGkaoRTrV/9W
Z+/gPYyZL6Ieybtb+0leeRDIZZIHBYnLJ5zbo8HAQzjmGyMkPaJw7erhYtFTSQxm
7pr1zPUCavmfwBn+D8RENYsG+8u1QjxljmbyL7eWg66j8plqYRD9LObnsgV90t8o
LMmjduNE1DsjbwJnmw2BFCRT4tqNsh69SjHrWfVr0lkzvDCdQGeNyMF4ZHx14KkW
uQSZDrYHwOoMhiyOvL8iWheMBQCt94q+Z91X6+/qzU8YxVZ8q2utRw+2gmftUfjr
3g35ozdkbDc4FK3CFS5Yb/YKz6pOa4k1TAvVZAvtAbRYHK9mKhGViEcOVCBDwrl0
gxvJ8LyBf9B3o5LRYLh1DfR6q5uHDR4gLns0Vtqfc5fq18Zo2bcJRKtip/FkzIuy
3YeF+aSDl4JC4poni9Ud/eAUpQR1HYnpNIaNH382yhrgMglY2ND3/Iws4Xnees6C
JHsbPHWqPN865Y4E4HZXIu3gQdMzCxrB+lXDgv5fDlkuSGl2oIvTg4NoEvCfSCct
mLk6Jkm3WI+1N/FlmFhgN3uV0pwgHGTtSbDPZrHJNBhGAKuPWH5rCgrOrn6TrtgO
GAMxwGZzlRJIDEnkHBi7WpsIqnwdoG6FpxcsfKjN5I9phjzSUOQzaab40hKlqtjx
tCMAg9QJ0nBQosVbHevV6ZwkRjTS/xH2f0srl56EQ3Wppm1HRDkS/2WmzKSTo1K4
x6LiqClBrtwNJu1UntERsMJQFA0m/zNWU9kjAWoXU9XcaHvpYJ+p2kMJk5MU+Kbe
lvfS9jbL2PzhG8zlxZ69iE8nD3y5CbKvuYeQACLWPS2WCPAisma5xL8snwDv8EY+
iVwFccb2GGE2XCq5lP/k0+BjOdDei/UqfnXSD/JKtZ1+ZPJA3g6qlKJn7WVveUwa
TZ098cVI3sMUWSNgqUxuJEzIUwV7ds64hUW1kTDeB76ZZBPULswI6t5XHJAECR4n
JgE8/H/43Jg7cRzNS7N0IkkXYa/5vezVffkjBnS1KVkQ5lAMJXpQTe7QWHQ2BrBo
8TjLmtA9gac8OLjyjZWTZJ7DOySwFY4FU2wsfD59RYyda5Czm0nliLluQCMlLPZM
LIRlPng0UrbpuIO/W7l0ueFbbtLrI877OX00NmYYrK6pFPmd5IW7mqv1i920rX4s
62ELQkmKNX4f33nrl7mpU6YckxO4UIjaXnSD0QauVCtCd/AQ3d4Q+1T6Edweuucn
LcH9WSCf43hOtli1CTVoDePaBKwI8ZmhN9VI8ooFICDL3i348nu6EbvmO9pwCjaz
350ADtfC3+9qdBRqE0rOPVBqym7t4wBuUso3sARX/Uyby2TpfdEi7ZLOZkowuYZr
ZYi7LbYf0AYjMtVkAlUviOXEIxjm/Avk8NDdJ49tFHl62r30TLZvMv8KI+TEmsYJ
AigUgt9fZACd+zZebw/7gK4hAEaOXNDZ/slbowVv7vIf8aqMdOBVRru2lZ6rScaa
DqGkWi2lEjnH5RORoQ7822MioWEiubzlS7YtmfU53RlMUL9E2BwPARtai0ZsX9kC
anXQPW+KDhHgmZnsvm0BThkCcQJBbpC1DzNdsPlra64c7NB3UEN6NCDYuGqYGKfU
uRSPfgUkdm5D04TQbv91ly2/ef+wrdxeFws9Vf0U3yDqxF4R7R+fxOHRQ1dZnhRk
i4sNzfw+UNc2kOGNBXDKjqRNwJTnwri95tvAXYEs3XaRAMuMNay1RuuTVJLMdeB4
2QvrjK0+/GTIGHF5ry6EDem1OMoD5zQ2j/kgeMc1eI/oYnbGrKQhEgJFDW0oxb8f
NzYli5dQ175bXr997iqRZE9TVWQpOHzjlD5Ysm1pmHMzjl6ffByERTK4rJimzM/Z
2PA/0hRTJ9+HQmXL9o4/OH9mbFolwE1olyNT5OrfKz8KDJgN5jOKmmM62qoJD5on
u/Xs0BAGxmqVfjSYAQhu7i2VtTe+h4qejg9yowxsmB53x7eAjDzaZO/VMLZVdcE5
NPd9N9CV1SgHt8O4Yv9lRx6HCH9SYnHyrascSYG+034KPl+NZWhWaasXSRm1TZZO
imLMdUgVWFWWFRkMY2w0z6Zikg/Xo9E6ACSY/Qlxj8o4noaT39VudmLiDIljlSyj
Grm7yvCfm5gsw4vnS2apmMCGTVtGOJmArckp96Yp0xXNdjPQWlYiBvg/8CBQgbaj
E1YudMUmDf7l8iIZpN635ksaa5yRPGnWEVDhZvEaSp6Pvrgf0bb1m3X9dzCIeB9c
9sTJzrbzzU2izM/22EAI0oBChojwOgEKeby8416OD1fNn2pskPUj0PBtV6tybWxb
Ogc9SY2S3GSgpSc8i1Yo7IY8mfTAozWRDf9Df/unUGXsN4oLldHNR/zFCvmi2RCx
GMFXw8PoHH+VJvXt9K0AqF99u54RyOr+NrGFKGPa5bpt4JHw42e3Zzf3zg+jREVI
XO5+mz1R2K0NdWimTk8hepB3TPxrJjEkympz2Bb3meuQCKgpwBwfG86S12ZCgVC3
3U1Cn+u90iCYQi7dfwnMfB4NArUO1EOXaqJjJxRF5rLP7BblvmfGvP4i3C5tUwmn
cJOYT1Hy5etuEfSmnc+LnrUpCjVrSpI0Zurslf4TSYFSHKLT7nGHQAOVIvEka2B9
D8Kyn4JDRMXQtuqKl4I4asZgByw/ZTvp/j3qgEQ9rAI=
`protect END_PROTECTED
