`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3S5dxPlYhCpTykwROBMoI8NLr3IjL+lMVOpIBWZb2dJC4zH/HEfPAk5zWw7aX5m+
ETGUpORCnbxjAEak3aOWErTRFgT5uLW3FaIJmF366Hhjs/k3HuvHygz9Vhvleyk5
UexfaX6hbAwLvL+gOFRz0z5R14Hjp9+SUzgdlHxHT9alX/yJW7okCXcKxgOUBg7+
UrQ9dOSEAqtwmKvrDfACm1KiS3O6PtPwr229FkXxZPVeZeLU/jFEFYyaUDX/jXyO
zFiWa1d5/hYCwOQ2a86aNEYH9G03zt/YxKgiWGeL57OPoRiD1w7Oi1+CuwlMuf52
fiTIY/MYFRM4TcBicuzMywVAliYUGZPuZTX406kaVrPbllpVbZJ2seo5qZtaCtnb
jClGiAi6MAHa8C7xMEl0ogrWGwsF0UOvDXLo9K4niMUArurtpQSZrZyk+HVnwxZ+
`protect END_PROTECTED
