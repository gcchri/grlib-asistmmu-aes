`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jb1nl2ZfBJXqdEz8oMD8Q0k80Fw5pDHwuoSPntHwVVMczZWke0j4EwEqoPcTNo4T
MMoFIWzAHCs0hPhYu2wVAD2IDjE3W1vJNo5H3nQRBbv06ldkjfSMKjPKjzWGaKJZ
GfB0jjfZUR+dUBCRNMZrpBnhLr+Gk9nCq2h1tKpJFZYPq9U3R35sketeifnvcOMx
Fi7MQiNFr9BAolSFvCA6UFzewKhHNZ2p3hLgOts73uolm1/mUpIxdQk6Lm7jdZtI
yliVgfeYV6ry66CUozRFh8ZC+bCo6e10tNpcoXH7W8q4ZkBa2+AAp9mEBtkax3Rb
Aq2gXu9Eiw/txXU9fhbypbnjki37UETncJSXcl/rjdmPL1Xdy2lVc39hsQz9zmQ6
XBPbJRere8qm8Au6LEruMIBe4k995Orbb3ki4jX0StvrdytVadsxRoChV0A3ASmR
Cf/zqkB+UVinAuKhhdfnRJxKMD6L/Lwe5ZabuSh2RSNyrgTBotLuvQNRjo/Pw5Nx
Z4jfbtLhg0gKOOMTqpW6QlmG66TLuxnqLBZdO6/+BJlBeE4ShcX4dPQc8mLBzbjh
Q5JHMi89lD6ViSd3EtqkkS/hl42q9rh+D2Yad3WDFX499ABTjszJ5FPrg25f+mTc
xtSBKoyfJpsGHQpL9B0iScxCXcyWa415VVJP2V1mk/l1rWSVyC5XjVseCoK6RrkF
`protect END_PROTECTED
