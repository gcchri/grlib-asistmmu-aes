`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+amHqTbWv+CUNhcdFRsxV7PxZ2KnlS2+tdag5eJp8YXlCctppl/OX88uSgLMkSM5
g6UVkbDO+vzGQIZ0a3ELmaxXvEhZN8HA/kaP1OsSILtj081EsHjMNI5wORMPUv0e
krvFCjyahs+2jMDvHdSaSZtxUICV5rfCGJWTcy75eQAvuyLMJZrbiaJe3jzFh9tW
Hv5DosDAqGl5FSG0SLbw+7z6eBPzrAepJX3y9KWZO/H7wQY5CsF/7CTgyLHwitqc
VIdDV/f9R7dcD+fAhX9HmCpzYBEWai9MoQ5VdyNktRAaaznj2eFOAnAeKWq0ZTNO
+pI/mw97X6xGP3tD0HZoDlw7O+y8y50K/xsI5hjOgLbF+0ST31vnXVvUB5MDGyzW
YIMWBOCuKdAou3H+85q/TvyPlYjF3QIc/2zUlPNDZypG3/p9wRVrhiuZynyoV8oN
HA3rDIxGwI38+bsob9YQ319eqjmoMxgaPM44uYHZ1NSnejaq72bCrtwEWEnABl7p
E6x4p8YYuX+OMvwex6hkPb/VxbXqrCKXfQzfa8V3z1RHThY6kvx2EI+x5DiwIasw
2DVrnzVstaPp80KcNmLRFODmadWTW/DkQIgp8xLByL9afJvGoa1EYW3psiOn7Mq0
k4cxSmyyxLZdXigziQrC11lQNzkb+efLsqJGDhE+WrKAdXMmqOlV0TH2fdSH0b33
HHsUjHjGe39ga0UehnDI9rvqGr8rM8+0dCbq40OxaazV1i4vZcPL8OzVCCImFw/D
hTdjVvT/ELMw8be7102wr/1THjkZX78NJMqiOBnE7MISxMjzCmmnasvuG6Aj+uMA
JCxsTDQVXhUvcXLxirjNcXc4rJBXAC3cvD0TYfTac/eNkEGFUeFyKz7oNskusTlp
9v1bRqfqfF80Cevkv9nuPw==
`protect END_PROTECTED
