`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bulhlL7hjq5zWB+6dCjRd3+dBfzT3IBWVeJbhagka5/p2WsfqBACw13YXj1qsXfv
+QLCBlyptGSIuPKHmnyoxrnvDdLKwX9hD1qh/90rnpNyFHggUmvuvxFooaJtaEfy
+0rYpqhDLF5YabQRYIJOK9wY1RCnuKjWqzxNGs0VARz26gwRKE2ITJhjxdp1n/1d
u0Bx2egb3vAtB4FI69s90wDLzFiCyk1vgOIyPs7bBzwxIUN9Mo5yZhY4OFWqO8cL
+s2uMsa4P2xETtwi98Ml1WQeD87swJwFO+WYxcLi7zotN39jfRmMA5GmMamfZl+x
wx9mJNbDE6bxSYLQiJE0honmcK8J0CFCeYzL0NxSjIutuuk9UYU/NWfsxQak0Jev
PFAdIEPy8sxwWjSNBJTU5lAfZazIWfbIEZE9BFekfhmNpbuHGc+YZGU4+jaMZBAn
2MNPU4IBDs+dWYlDIG9FcjHzmVQLoNWY5Mrz4ocF1/w4wF8ouOAIJ64Ro/MxcEQ+
U/TXXFroHxO/ZdR6Rk5XtJ1/iU7TJO8t3uDV3yd7kmSKyy+SsfUTm7x3XNVHG1pQ
cXdBC+hV3/ARdUA1xMTGDvK041B5KMNqM5EAcuCCBsFif6vsdeiLDjWFvW7zAE+a
/AXdqCe2Wj2R/f81GhWDJOkFdxXBPmXXmOdkcarq2C1DUnO+yqz9FxmOIRYjleun
V+kxo8xBCVQTyXpcRymcbSrCzy3O841+wb1ec/xicTxIwJWRgrvsXd8DpCteB2Mb
/5dWu/dFpbtNKG+NCqYuQA==
`protect END_PROTECTED
