`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1S4oxgnTcwzwnT7ykY9qt8Er00uDHeOq8GmQh7cmi2qjagNKSoKh4+t1mezaK27+
hmVZElLY7mLP9qmdfllIAdWIZW2BVlAB+/sLsin27u0JRhyhCGt2dmcfQTvbFtCA
ry2MmeYceQMobsgnfzBpQ4qER5TGdP+cbirjKVbn3x3L08VAlsnH+b0FnKfA8+bQ
WyYUhOv4Tu/sdT7apWjfwxM5gyVhD5FBL6TywM380Yt/Inaxfe4pXH08fVF+d+pt
CI+d2VqCqUmF0+76U96TO6pWBuSLxjQxRRfkUugTYfqy7+iTWLqxVDA4s9zvTi5g
jibFLi/5FfwyrPaGwVmpMLzx44zxVdlAiXqQ9ZUmYEBhn84ga5rXURN3EEnvNuyY
n0K0S9DOOnkFGEMua0wkzl9PLW3srqUxfAPZLUaPzvq3yLPUp7YdSiUHl4k15xNK
ZLwsbM7Ta2K4z2yyq6oQmT/Wj31lwXzBnY0/1enKFxZ+FoU+t8w7BlaTujx/I3/h
YvK76IceZH4pnSDVnS9XeS1oMM9vyruxIBypQHzATP8vSpEiATW88VEt4kMHR/Kp
t0VYR7Zlezbj85CaViV5HU31ClILj1U5o8vf+a2AShI=
`protect END_PROTECTED
