`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbLypFfUVMCG7HFh0xZ6mNJDsX616/9Q2hvUmwwSVEqdtvuGp6sL9WI/3rmWMsXe
UXkBwu3WstOKsPsg6K0gMJagDGu4pnwzHB2Mlvy4wFinA/WZnXk4NfEFxPjKWF3b
257uZWie0sXydas+HPFSoyS+NxCdXUuYfhJZibSPsOKZat5Vss/EL+mKdcpwRA8U
xPtCkygrJP2ydR+un5+p42MFb/y3a785at1FlsX5t7wAV9DiOZBYljfZR5iSDBQn
nfD4hNk2rRzzpPMjGltHlkasWJSz9v3iLsgmjSq1Qytq4siN9s1k9E1dyShyWRoC
3XyI3bGFjYcGCB8OMEfo9O8IF9YVbKSfDavupUG9AxzKc6s/8sFov0Owudwp616O
3S2W0ZQnFmHz6qDyjWuI6YsVUALb5YMr7/8oBMvApvlE6wpfyYjcAOoLosbc/7Jj
FmwZBTXvelsYYnfCCCAGeVIePJEApLNU2f+5OqylP7KCqbdG/0MkZlTA7UHgT/EZ
21EaICcrpzHzHYYBCtURMRlLdVvAOwi7FQnf3eK3xztdAcIq4fSIqcMlp3/j+LG8
xyOq+aYKx4up2K3/UnXakJEvZRNvF8L4tU0tD7E7Kp+xwA8yK/AePp7PYAGhsXCg
pCE7oWxDAHR13T1lhKeI3T2jNTvlE769pTVxUNUWnDkm5/erLtfOD/YxhA9vPr2P
TCPVGRvb4ZrZpRMUgr42m1LpqBYrbRUzKOEMXJtJnY1t4ap51N4bZZdl89DbDiRv
EEevfU/+Jbr17Ys2apNQvB9DlueZQblbFq0N7rWLsHxSqFurspa7GgajMMFHl9Tj
j85Xunbefa0mhT7HzrfI9hpWQJ2dkkFpELH9klkhLm4jHK17EwpAF/tiFPgiXZvA
ujPkMCvZkOa/4v1r5vuWUOoL1sBf/+L4PVZYui4APfo=
`protect END_PROTECTED
