`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gxJ/580HUoLcXNaVk258BcLgmhOQu20Y6mf4gnx88aEkln2GU+IGcfz89Vr9mxhq
iM98ZZSBJifdSasvJUuQLWjVAkt1VSloPjRGDGZ+unfR/TjRcVvxLMv2kEHhXaYA
YWpqqFXw9O5Z6SxLpNm2jaWXL09Rb21EhSWqSHRSQEVjb79+uLT/1m4HYOCv35/Q
6A8NK2j2r+r0bRqV/cPs1qICOsSWy+fUJ/glbVjZCjwgQG1Zl0gmjJEA6Jr2NKbX
kvrbz2LjQUqUTZhp9uFj+QQfJCYPCoGvYWf5cYw5j1gLHGt0icPf9uDYLgOhUJcH
pF6hWT8AxOtz/yZb+gWO7Mkbh5HJswflewe1u8IrNPCfSqS43IXQRfm/dYvRTzHz
UVoe8LbkDzgAlCFtUVjjpV4SmIDj3Zm1StnSFCLmPSj+kzVvYmBxhn05DDPu0eXe
jn17dJggjQ8QE/9hLTU7+ReqfPW52+1YxGD0sCh2RMFF4oamO8d0cEKJV34O7++A
qD11V0QNjmnnMUJ5JhBDkSaaIWAIyi3xkxesPw641M/GPq/LmSyxhnVIVCEJEFcY
/0BgjWj/MKfnhMaYlqbPY5ZCQVt+JWxUvSK+RHgZ167jfPF33ICEA2UOyIVwdh7v
YEen0o7UcVNL346l5tnTaNEU8TRRauwzgIeEHc8B4JziG1FNd9T/ei39/zWAMIbD
ZFb7m8RauPTLlgmcmOLnb5q5bnXO5QXbj08DL+IqFn/BbCyFQSQocTiq2B00r35d
y+3Yv9yudelciCX1raiTDhkieiJvgsWJ3HWmbhzdKZvIjTZXiuOYmxKWOx0yrZUY
vvTKZGmspRsmr6VgKLCx2mckLCE3FMrAJGqJxxnZXoa4kUjRa1/3BGH1efvxBqNj
e3v4fcFc7dlxB6QVxURZte/BAxl294/F9ZhJcISEK7D0oXOBp9C4iCusSejWTEDG
PO/PqEBtVM+ow2eABmtcimLkDt8arbota2/PVuM6R9YbpTRBLHNcv33bhnbPmXrw
JjErOJKfXCFVYRbP7IcWSEVGR1R+P4PUkZ9ntF8IroxdCIMuoJ2OD224xZkL+IlG
y3e8bre3InnWSSiHfjUwL19JR4QDatEgRrkq9QCzBn4J7sXxCcahUxFVQaVXxddo
ghfXw2nYSWO1pBjBQmADvzez4GIF3TY+mowfJT395HiNkgPOzApK/2be6NFCTC/w
tb/7JSTrdVicRvloPIILT5sg9kpwOKebYZUELqZ7jG9+3e3ZKHo8sgQouyBEUMTy
ZqKXUkzATn31FJvfX4MCB+PDUq3fYJ//cVeSWgZTj1SDhBN/A7Ytz6gXUzoHr9FV
APwu/2QP/pTWV9DEhDAf/m0F2RrSiysYRqZLI7J6f8gaZcxPnIHV8p7qI+jGdNjI
2JUhfWBlQ3t65PpJkgjJjtwC39ceTJXkNG5CRMtzsd5CUHnS3vNb+28kSjbbKQyG
wU2fU4+GPqsB/pBVdyhklQHtvHViXjLCIY398GniO45Jgo1/yyx9jPq6ya/iK9WR
7HcHZaMlOfb3sdnqOHddWM52lfD/ZQG6DxCkMa4/mNrUWPq1z/QVLj93CuJzxRtF
li75QpEb+8498r0OLxjFBwyMEKqC3hZ4Wt6qptZ2yGDDySUkPVakWnn7UmazSyjo
dloXCrUOo33X+CSojTTDwGB1qZYIxF9VLaKhrkNIiJv+D4SgbWuvMc+RKHe8Klh2
mheHlzCL0w7clsp9+wuKgf3MLHQyEYQJDtqupr60dhAE0fjyuxVFTi0wNyP5Y/HN
kEHauBFNg5xZst6cskjl4qAthBpd97Kk6d1aIo73WvK3qMwxNnBe9PmSrdUIsgYt
7GGya2v1ysqB68k4hrxL/D2QHALLBFYYzFakzfxNK6uy6tU0NVoViPxiK7tgqP0F
tmG91/wfOrV9+k78YbGU6TMo1SqGIRdLRJXfwftWr8nBGj/QGi+nUK3f5l8uPRL7
GxBY6/yx/7Ylis/aKJGN/K2lIQZLgTdQFsU/iVg2TcXI4ljfnOf5HT4j/yoLJw/m
WvsezRS8X8XlDR7/IvbDdmbtb6hb1JCCgiVry3PPlrKQnjaqQZ+toXvfvBc4PAzY
icmqCIjzFXtHaeC7pIUYm0Rbp38i4tJkw6PfQ0SZyMd8nZ1yCbsIpUyElWrDLK/g
79AIIEdEwIJqDs3svrciDAXrF/GaEticbDGn83xfIGldWAo0jXMTnxE66at6M3DL
joEf9vzGNh7dyAXhuQpifFwnCL9mF8SxfQLv+Zyg+wDvRSANBYQfaKNbr+DN7vjd
erONnBw0veN1Yj/XUa0neMOM9ynFCtqNwJjpr6KeBhbftn6LHK3YiYRRtqnugB49
BI7E9entu6mMAIb3dHjLpTKX68YpmwAldZvpy8drCluyl6BRAZ/81RpR1DXpbvbP
KQxY51SiMQlI7LYjC9EqzSFq1DYzYFFoUN/7O6VCoOmh1/vVm7V7SB305dzNaPO7
WAqGttcrukT4gIvufoPYpaKkGEcWweweW/EXxUpNtRdffiZVZsq7ojbWBYPDpEyf
oifcNPc1diqM+qfRrp2NVwa56p49mSIiJ8cElItwMYwNlYF7YwMdKoLSGnZvm8H9
8Gmv+Sp58qTvN5G5uk8x+eGNkpTOwJ02dGhKL5npJLzL4AMncFWURFM7Q49804BY
xtmeDZ+hhcnoZtFouTL1Gm/yzUk3VZUluP4kg8vwa3X+Zg86SfLzA1yfBZ6XHOVI
0u2jGMa/N38IL9j4MyiuahMZ2uKEduWWWr02/kvC8E+CviA6THimJzDELAaJjg5R
zQilzoPIYT1xV68NPClzKURz+uCwRPdMQjGxOSBAbDTQxqkFzfzYtTRWHDwzA3Gg
eOwH0Roc0rAz7paM1iqjUV+uxs4w4oeingPg6bI3I6ukCtGYVLEiu1n0Qnxx0o5L
/3rQ2+b1Bz6obl8HmN4EjUlzfuarzAE+fKPAY5rJh7kfQTsEw+tUQpn1TLrfUhtt
wPJk8s+pzDMWlgzHq+zo9a8KBk/0Zlf0XOaNBOFKKMzXsEvRI4+rZRMVDFWEirYP
DUoYJaWErLZuPhZtvDboR+oWdeUTq8CpGgFUYhznxmTXPeRHEtNqpGoe4IpSX2Ft
mpTAnFiPk5HiEcaoo5qeUw==
`protect END_PROTECTED
