`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3OXCZjSiaqWgIWuGRHnwngMh8nehpOWZrNwGTP9MBZDErYUSJqV6nqz4ZiuDfaqx
A398pZeQLAWEH+9Mne/rLE0AMjRSWIvHCLdT7kXOPKCAjD2uTwUbr1Jf1RlsEfCS
xSWcK3AZa25oYg11byuvhw4piLw3Np7Q5g5pII8rl76iwMIPusspOP0RbuOK92Ju
feldI96OTAANFMzpD3WFY8MEb2TWjoJoWIHsR35d940xFFizpjS+dicMTE8Juxqh
XDRwB98XDEIxHAoHOsWm4g==
`protect END_PROTECTED
