`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sLqnKH/ZgAc4QolmQimmO78hezoMG45MyA9pS3ywixbN512KMw1ttMZSiTZPRyUu
UvlhfsckS/7L2J3S4g0OOCSM9mI+LPkwHTLtUwr8wgPf6rx/oAwYsTR8wtt9nybe
8dJk5Xqkuff4rzwoGZIh/dV5Ym8lUTsY5EqY2ysl+fwMv2ZEiq8dndf4PQsM2nQR
t/9u+M5xsZbM1H6xbhWOogwmAjRR4xoJwTYD4w4sbW/Lu9Sbu04x+qpfPX6I+wRN
o3KwHf8Fmz2CThtx0uUtBdFa/Oec0cJrGVk4rsU7wG7m977P99q98kqcKG7RR7Gf
3meUHC9keQGkUEfrO2K5DhVmlnia6swZa0gZHxoB1ErGsclOLkxcEqzyeWlxm7mA
5IQcpLWAyjchE+OOYPrZ2TgXtrXWso3uUYHQ1CeTSqnMZfAfFaDFVlyDctwCjQ2i
`protect END_PROTECTED
