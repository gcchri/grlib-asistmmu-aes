`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EekjaWCjDf7fIlOz6js5z8hhllaQaTjKuhHZ/8LRrcHj6b8+7uNopfmTnFb7VjmU
9CVc2EXV/zS3cC46T6IKPLVbOtdohQxrekDPWY2ZBNzZhy25w80KCUYrf1bzKrTS
F/ez6DcNtfMyIIPGryuz7cdmR8WqeJKgslBsjLGOqAfWPizk1yFCrSenOH+l5Pp6
yy++DafPHqxDLvlGG+Fhy+3y2g7um5RvGuWMeaSWlQ11erqagVfcJ+dIn85K67P6
1RqOnkpqXVkZb58eoDUQ2gp1QVYbcjdE/du/Ci4xysCXJPG59323Fnvmjlt1DGG+
ak4FZenvHaz0dT+0fQNIoCTSQTQ1D4Mx04Wbz8tifFYyOm8BrTg5M5DNT2HxJake
q2YSQGIy4E4YSzGHujaFn9tbqGA+jjyOHx6bPI2Rj020HdKlMAMMPOleoQiDZk57
iV8APMTRz0zm+gUFmZWUPWWuttpgDF71xH1HBu8b5h2xmk0f6hFEuDfelCP91/Qh
z0KxVH4Wq5HDzDtLQ2KIN5Qc4SC+KofDsSa4VXWw16SdqoZnRpNoi7isrbA1QArE
ZXzpfQfKL6xEDlwJCc3iX9Ezy3NSp7wRw9BhPAMRYtYTia/C4YQDQKFiAnE8FP3x
qhlWwc7e1MvxoHLhlX+6xjhhDqNpa5z/5R4UpYRgXLuOB9mXbhsoxD8WlwJWNmGu
FT27Dl9l7hip0szvE8LjKASmIWNRm8rqxrFhuL8co26vW7FVU6RqvEVRafRXfYAu
qCnJ6sjxM+IGhfJFvCqq7vKUEF5/aE2etfKpKA2pLMkxLI4kQh6r5dRWoGxKl0+Y
YxkeZ3ytr9ntTML6P17COw==
`protect END_PROTECTED
