`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/vwcagHixpLOynoE31oCsMVQd+0SukTqXyX8nBWCBhpl/w/ELNbWfv2/ONgQkZH
VtOnxHrrYUz/2XHGu0uxh036vhsIf3N8YeuVZb2qa25BIaNSu9hLsTNZhWCXvB5i
Q2rOoTSej3ttebL25YRxHA5gFyxsnfnYVQIyBEtpuQOjom6Gt5Td7cp4UefpcN/i
AUBsr0ZrjeFBaaDLcbbYEEPnV6ntyK3lJccDgYAGGiGeSvf3+rlw6OZj2XT5fnoW
JFxUgN41bbAKX3bHua7ckEdI7si6MJhIyYfEske2hqnIos6FwwMpeheL/gpPGASH
kF4s6QXJuzSctrXDso+pBSG7w/+UlVz5JtEEtqnQ3lGTQJA4ryMnjgymKLeJWLWM
jGnNstkMpYwVnMwHVr9RAwQFTdAsnYvdT+vyhtLIO+zXy9x463qWAFBLIHdeUHkZ
gA+wPe8opzHgyePmBG8D3p0VYrR2EVAiEl/cJ/SUV2uLlkKlDqT5csRkQbjlgVbH
cc05kKfy9iZI4cmRfKrdhM7hWoyzUm5f9gVPJ16v2QtRJ3tQEbeF/dXxpsKyttfR
ZeD9qE3IKQUSlzCJzcDzr8Muk1j+CKihOiAOFmPO6CSzniYCb4tdS82E2wiTGU4a
no+QqbDEm3a0E1dIrnOjQyJ8qJTRefLCl7kfzFy8uUyU+46Y2SSxOfedetn08lpJ
hl17OR+znLMd2trweoJ/NJji5hM7v0Xci8lZItxLNbpjbAmwa95ylDzB57UAiDx7
Gr52mjMX4hY9XRRUpPwzLOlEUj1IGqwMp/UX7kw1cG0Tn0IKj7tPWOBdMJ9QYgFd
nIOTwUl/G+UDQzxezs8MdOu2bnXhSAnCkltDEzBsiFfYP8ilw7NJpbS2JAfigBq4
FQW/FNUzHpuVJxl1WyZpz2UuDRJQHxvn+O6yf5SR2zriW7LzmodA+H6ZCQ8dmONc
a3bzi3zsLPMn4Jdeoz1TyFsmLIKacVBpr2FNAPIZ1eArCu11hQrs72RIYEUA5bPy
k0aLfGfFBtjgH4ulHwG4DaAgMd9GsI/OO0NAYYpOxr6xSkpJhz1wLysF4BseUQLB
kZF0FbiH0TS8V7p7uxQPlQ9bibn6HQ3cnYvCSXxICcnqJowebV8drDZZbXZjzjoJ
6rd+Z+cQLweckTNPosvcIimix80reOx0RdotmXeWMgduH5ivgVXFDV7cz4Mn66Zu
jviRIpR5sPyAjZzq/pJXVKaEiTdRyrNPRl9CmYKnahv70zWJ0PMi6+8uckprNZ+z
8yWqpsPdIGpmIZIvhA9nJkl48x9M7/xtdtT9rfhVCmxW4lCEwspWp/I7P/L7yiOu
ISjhHerI/VpAKy1KG3D/nK2bwOB5L77gAJHBQYDhquKLtiC5HyZVLIArqVTwNaZM
CGKVYppC6mrWcBzoJN8jT+iFq1tDVHut79Mj7b5KUmlN3maTdWfQId9Gs9/+KIky
cbuczttVl07BHH2/Ek7FEazivrxWDYyzrnIALD5mxRP9JKjkISt7nqaO/DDbsDVp
4WmMynJcfbiuQRBZVDWZZlWPiyolg4ZwVSgvDcCeD8B06kAjPPZuvp3OAaq+vqE1
S6F3+iYoBtUSdXJIcDU1QKouRVtfBOV/jG9AGy5E4C18rOtAlN35Z7N7bZPyegjS
4ARPCEVmcKla9qvcnwOkrLgyLSim0R7lcaMIMYF/joQKdjKHF5tlsWQyYEmH0I90
i+NZHwHbq/Tylc2cr5jyGMUfl/f9xvmF2XcHe2DGZCRumRGBkSg3W49VFGtlPdaB
eHNdvEJkEzOmx2oL3eCwbG8Znw3kqxNnM84piCGU7h6QGB2ZSzHk0VoCjWcZ1lJh
DLzLnduRpcna9DLsGd06dyHyq/Rt1tXJ+4+5c9CAKJMxbUl4f2hlTIFynxIttG7H
20TvDvlHnnFDEIQkzB0xkyV6CB+cfAL71LQyPQh2u3aUv4jGLEX7d3lYTssc4KxL
V5mvKeW0sDar9e/wVafW10K17/7PkS5Ve+zUD9n/sTyJecwYidpK35qo82QdlQH/
zqh5HlraQVgA/wm7MWa4TLT5LF645PAAqT2TC98QHPHC/aiew2e6huIUfCr/ZkNn
bYeRsJ53HI5OxN+9paXFeqHD9eqi+o9PIylyMVJAXYY0Jy5ccPOqAGjy9A4bmDZq
bR9Bvzy/XHdaWg4kqxtofpyBPt3AbIr686fRuvVwzJ0+QcMitqvq4co77RKTZwZ+
I0yWwuaBeCdxdEJZEcLp41j66srVwO2beUwzS82bRL6sCrzTAjCtCOuEIGdPuep5
qRNzVC4cWqL+HQ9glWrgOPEC1wQhvvHkRVhSCsKcOVI/9tUsAQOKrcCYqq0YhfjJ
FVovfbNEzwQtOLtLlHNzevumDctprffeFL7FY2kwwx1QPpEOZMhz972p+EYFXcOM
g7hiya4RehAXGrIV5WPuuf2iXzmcqJtHVWoSkVziKXKZCrfzRkZVtFCDSvFrjw3Y
PsooCzIlTcqv15oN6nlQSGykPBNKT9x5+9zriCrO7rZJvBO86H3JHLRvliIP1Zg2
GyfUnk2X29eKHkAeE0WRDSkMiS94xW9mUcMwJyJxFLPVNIlQCGtfyMFKQoMHCPPF
PoSJENOLW+UT05fpCaiNQTYw39TZnVQHEZ+u58fay3oWYltWzwMzxUgVxQm+iaU1
Mu0RNqkG+TnN1mqcNLcQ6sxH4s83pisRiyHhknZrcLtJsJNA8yGkdVvy4frx52Gi
d0xl1oUrvQB/wC6cecqML9wFOKrb+UOiHFLqetKkDR4OqrtU+ezGgC4RQ2SecBQX
w39Eil35WNA5+H2gfjYsM2Nbory+157GHWL77/Noc0l2QQldQOjmfo99Lioz7cpN
5hrbPMpYYEcvSttNhm1L8qpllsMaeTx3u/FBLa8DNKGA4BTXNcbzsc7Rtn9vtIA3
h6N9teEr/ef1Vrwm4n6hiF/CGJBMqTM59DUZbmWFb+OvhE0iGAwh8yE+bsH47sge
pSa2yBphhy2iLQHsoDMrZvmOq1ZCn6HSDV4JzFtrJidf3rq5Jb+8+FKSf+XYUd9X
9J687pMV062rFxZuNm1kmWcWLFh/fnQn+c94MY6t3KyNHEG4UEnyMDbiqrWUZYES
A22dbb8vrEU/BXvAPvVFWuRJpgAVh8E73tmvxXM0Y7wf0lTpbEz+LSfiuGMeJyHv
AM4MgN9bj5QuPVqKYqifY/4lNHP+r/TFXroNrlmRMiocB4AGnOWXF+Bck+AlrCVp
R3EFJqc8AvOYHwPUo4tR0qL7/Cmg5itbH1Rkqb+EvGLqUQsDCM0368cvwR1NtZUD
A5qtOH6cTnGWalqMWHu6dVJD45E2b5O2IOCxgQ0jer670ljyF3jnD7EiqomniYwG
AiBQ6hDGQFoDHPmFZsr6y0CKpLF1q3MprbGKM/U9pCZ/wmD3JxyDpsbR5LIwtI1W
ZbRnQbNgvFynMa1eJVT+IyM/I69Row9POpQsNBBJU9FkwOR0GRA6akNAAf0M/ULC
WSPL8XM2XBucTCA24cgd3WXOyxtnUu7AEaWTVepK0tkFy0BJMtebGiFOSRp3bx4w
JWpCppixW+/frghlXZmOZ6MGLmJrIvSHR4pQ0xStaML1hGknsupwHjI0GSZsvOTJ
4jxV0exTfRHlcVPnaWkAz47iy+SnTBKixRbLjDQAY93XarH+booSwAXQQuUtHDhE
TsKJpLx1U5ZBaXuoAeOpENjqf1b95vja0uOg23L3trdclJ/ugmu9rN1ygnAZot0t
g/13yaeAzMOVUXmRUcrDYXql0LHLXMzfSTUKwBeexferlUx2P+ZLuH2rY3w5K+AN
XPgYG1/TEcdU+rMVjTpwjQ==
`protect END_PROTECTED
