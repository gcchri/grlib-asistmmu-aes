`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/aY9dZOvkF54YysqQ2Vj8YIhYhpaQ0Px5Qt2ECX9AJXPIraEq9ZJXF0hxlqXLA7
M3KeEtxiILN5BYIfAXKL4mMK7y7nxxws6yqoVnWjPumHDXWRp2jlagUtrGGrvy1s
es4VznU6JiuBUcAIU1SrEr2QCvgFkuXCnjYe8pY/PASVji9jY75vRIsa19XTYfZo
mDIosNKp5jVBSXxsbQEaygksAt+/P4FE+IzaFyooA/0AHG2nirHDfMBHtU2j0W6v
MTv1nX3OKnixvu3FomZxAbS3G5IgZmk32bSuO6xVc+9v+A3a4LdHZwh4AIILNGMO
oUZ8ZIOVRgtuSEFYgG2R9Rkl84Pt1ocwz2kjQZfpiWmeO7HLqWFKCbSbq75ts6IE
lk+E8W1E2YU/Ie5GIj/7kT1DJibZ23NZ/5GiWVZ6qFjkKcD/46J7BnqTGrtedZsm
UOxjNUY8Yag1fD6yRJflb9cuuMHkKVSlQKT5VWkPpANXpeIpX8/nx/Xf1Y4EcpkC
`protect END_PROTECTED
