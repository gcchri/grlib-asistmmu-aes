`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5iUbwIri+MEHP3dIcxSNYCANHFmwdb3HGs+s4Ni76sJ48+87vP8FUBC2tsSSzA9T
mx6bc42GOFD8Nx2iNnBerjv35kgO5Ww1+KY18efA+yzj6o8GpfDtXVq/8Ix2Py7Q
FxQF/ekMZV125XTW0dyvgohYYClm9TqN0mxKK6fADyXGvwa1S90corxLjuLiavpk
XchEiRlqnBzkJoOYoyxfX2H531Hu5h4PTI8WWHPQN26P4V4lCt4LS0RGzttHbx0o
OTktNG04inuEWedeL5vUYvcDEgg/z+2FeLy1CHKuTKQRNHDIl5Hp58/W9SAaUy/d
Ga/zKfDWvQhrJKO4uOpMqj5c/NZX4IdAg2eerSeA4qAYuR/Ze/nfzLxIgv82m0CP
tuZoRfNcGKu0MmGuufb8ig==
`protect END_PROTECTED
