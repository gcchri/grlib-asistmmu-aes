`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WxY9JseyorOgBZxv/coomaG0xB5LkrNJ3mDU2knz5qIbikZbdYc8eOu9uQdaExhW
9XCj5zQMzLfiom5g5NvNriKDVuu+sdhFEimuZVw5XFfDB7S9RQQ4gPDwM84Wtxza
O4DuBB/d8Ugmp4nnlQpbpSAVlB8vC9CzHj3mlenIwHxwfaDb+/ZGgoEcJSv/MTEM
KxhCexVS/VobZm65M8/gvZjrdnidLa66aHddPOX0pbrRUnJnVdN+tBkKvsw795pS
NoFdydfpcirJJpE80HBZsPGtEqXiM2y4isdjUib/NH8FVW0xqVO4EzoTfzgfYntW
8OhpbORzefQ989ftNlGiR40hJRydQZY9jq8UZKll7FZcutlCY4nl7OQ3BW2N8qrm
bvJ2zNQKiqUAxWLeBeH2I9+16etwBfs3iKcOB2k4u9CUWZm4GglV/hTbQXHywmY6
jr0yl/vkU9yB4yfXxVcZat7FBQoYKmCOEBf5yp219Igs2m1YTW3C/EuA2OjdWvNQ
62E3SMF/bokB/xnYzC6GV8kcS68ebpf2YazwsKZAAGJ4g9wzeKCDSwdj+Mq4Yqzl
O9O4yzlsIY/WMzqLWdUF6ymTly3fInczh9vJTe2FIxXE4Ek6kYDUDNPNZI0zAD+F
b0eyb+8kdcsQPLZBYAAIIO3JchuCNv9mhD7M2XxT0oOBsI1YMiywHqMT7x2ce4Zg
`protect END_PROTECTED
