`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Efu10oUa/pB0x0CGyFsRF7samP5ruzSi9Uqb6VQlrtKxwzeuIQzHXlQ1KcBJgDxY
2atDC0iTbGJFvFD3sNiDl0vPABrNThTQn+UzFNjG2qILdKVHluBT4lUv20EcyKFN
Z1d46dUnpd2Cr6tXIvcnxRrflMx6Fntmpb+E8dV9vRk5LOTwdThZhYzWKNIAjxmV
oOLgK37r1CAjZ98xdoQ5wB80Cs4Y/yYVZhIatqKBrUciL0mHpUvZ/4YReFJvH2n4
amucFWuJH1Ly74lKMF1kusZTzCEauSxrLjdex1HAb/Y9WVcqJqgdIl9OIxi253Ik
+LxEJasQL4IPeB9CXBx1jZFV4dAyVGcdWPAiOpSmMVZsHuplpj2E372Hb1suEdIJ
yHbu3nzmbV91ygdI6babA0yt5wHRaf1EA4fFi/R1iy62yJQn+t7yier2o9+qzAaF
Rt+/k7XvsRGyboGRu2Hs01x7j4Ar5rOHgJLLVt9bHDNTlv+x7inSDOzlSWaxsRnZ
TQX/4GOUXRIwiKWcxC33JLUI9GO7ooJlZ7Kqj84P1mZiUnn+8X61zwxfViBxCsFc
9ryiEzmXRZugs8VRYBcXmKvo7reg2ffGE0CI7D8LSVa4S38UpuQP0jXEswO2cW1V
of+v1hP2FcU6mXnH7kXmnrsmmn4FyEMJklHm6bhod/V1BoVafLwmJrTYn6/PBuke
6RSlbx/883kLErzidIVOS4hLvU0piITgoGidghWv0M+rPKtudQDVxoo9K2W6MZSS
JUA7oRCVOc3ay/KTdeNxUpfeLn549RPoXkijgDwJ84r/ojbD9DMmVKxqvqLZxiab
rIQEnqfim+QdsYg3R0+YNOk0I4fn7SXy1DCmA9rtouB5XlI7HHvWrcYq5MD9zho0
9Y/KUhv/oVRScHQl/5MFrZCNpmH5kTScVjbdpWrdLc4lJGgCK1sTHMKnRsVgWeUs
wD5pFIJwrSFqGcQjgOUVZQ6MWGkkgOmrv3zHZ9O2pEn679LSw+V2Owa6sWSONyfG
8BcVInNlgDHycLdhWsT+fQ==
`protect END_PROTECTED
