`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bW1vLLVsAIzwE2VSQujIGv3dC12sBro1jCJy4KRHZQzky3j0sfuj4oVWlzVhl4f9
uDJThXnco2Bg/S8uRsdX4UY7E/B/ZYSi1Gh/Uo71KNKTSo7zJ4mOatLgUJVwDl7U
jDgtzl1lye8Wj0V+QacMbWFrNcpARpqrL7/Gq1pYv2mCWT9eDx8EAE1yNjHCxB7D
URpxtflw4VKJOBrO9aZ60+hs/RI0dPRqIRfxeTegRGejX8tC2SYtcYD6AlJCh/mr
5/ZAGIZ37Hks2UyHArTIc9AdN/z0JVP+PxW2vKq7wO1sxJAvwu0roSgzW3uqeLYz
wvviItrPdabyZtSfsVJQ4EQaQTcklKW7Cmn9RmOAKBhKbt7ApDRstrnQmvMacRfz
J4gIgojs95oFjpTcr6w4vPR4ikCMJBR9sCTYdYuDXjPGnNDYilB0BO4HFuS6vWms
ErjCh5l1x/rLTpwnhHLPHmBMrcRhmAiF0km/+rh+x/0PRRKCj4X7Thfc3HhjS+a3
A8OCT/ChcjteD5vxTW1Bs260e8ndS/XQzUW2kvLr53TF1cdcJycfLv2lTZCkbe7N
Mn+J8haQq2Etb9ho1Y9q4uoHz+NrjGJiIBhmnn6Y2EZjzsfN2UM1L34pXpBQ8MUz
heaxKtkFS7XRrKe/kIznJYAwZBLhgK7Tf3/0Fdo5gwj0z8pUvTJg+FieuZQKiW9J
`protect END_PROTECTED
