`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrpP/0OM1+9EXw0uWS2fAz4tYqgaLQg5oy43iMm26VHdIwHX3xB8Ia0Ep6kFBObZ
crbFBP+m39gV9by+ZvRIRuwrZDARBnDYbDwHC3pGXW5TItCexcs8ws6z6Db8zuJt
lVFYjveQbCjf6EPYP6bvwTFa0Q3icebWH0cLUnwXrkD60j0HmjIhrN34S1uSLQzj
vNmS2SIjo6qfKibDBNy4kN6fn2bJqQ6ufQIXho/n2m1kxL4IV+pzdKE3uqYaWAFe
AUoZe5PZzdprVhi665PyjH/u8h14aQ+JRYErcsGnVYoMJMZXegYj5e+O699myT1s
90u+hyTPw9fbT/EnyzL8sJggUEpWX/v8d8PWXL1lKcPmJVrpxRhMzxMyaPY3r0BH
pGBt6Rjpe1+XqWGXltOpCYctcj8HVUZiOQNWGAevvf4o50CQ5QIkCbpy9DIhNeGM
uaTpApE6miCFhnu9DQAofGaDUuUOnWcQf8Y5fOyR5dm/PzWlcp/IW9CntkgpzNWc
3OWTX+CxFq3A6oNA8PTyNKm8ldOfe+Xa0f2/ULDSr+v4EsGxEEjg/4wcYlTKUwTj
yB9hQQDx0lGqqN9l02FxgAfcbEhFg6EVS9fl3Y38YbiPYV7K9GUXmt84R8j3iRz3
vZ54tEK407za4dALrK2E73XJ1SPVgixElUkOfYTEB9KR1UKIbJDY5YVk2NlORNvY
7pKAy32QceXHdz15WdlPfev/gnmsPRX857xND/5N30RROtgWOAiWoJBQvBLFOLgy
a8HCFhOFiaB6KQ0g4uke0w==
`protect END_PROTECTED
