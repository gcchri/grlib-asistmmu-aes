`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T19kTPdEuiuy5vdbJyvkroP21D99P06eKAmtTM+w/eTH54WOxeh3cMCEwr9T2c9b
IR47A2Zfy5YrnfNxlDlddom03uJnV5U4oF7X+RCUl7tJ1rILnGlIeLf1xVQvT9O1
hny2t1PTcRhuoauaU16sDZqX1ui6To9x5y2MH4XjszDy8dP+0ihYeroxvxf88E+3
lEq0aMtRc+uUTpnkiiPIi2yntu57xYROz4DKX67tiYXKXSsZ/dKvQ5DRrskN3CYR
Tg6gKPcovy25OziupO2IrXECRPVkPLJcoRVc0PDALOaPJmP4ASI7UEFqLClLJ9KS
Mlj2/PKW3yN/R8A9rQDoyOGsGGMU0gxDIDkKy6xpx9qtUonHJpz+xp5m0E2nC5+S
f43sotSMMQudsR2hhZgZdd5GH7jYQOF0sE0Pm7x2pU2AGTV33BqcrZ6+Sno7TV6M
eVf0gmo+Uvczn3Q/jS/+LIvR57epXET3dmJpolCpLuzExtyjmwIbxx32i5bHs/2n
AtuZUGKj2xbKTJXkq5Jaf0fT2P+kayicWb+JblmGGwry+bYkmgdAshCemEAovx+P
udpxND4lHwNXn8HG9dRrSyHBVozVRh1BMzUd4UfxLr8WK3mRCDONpyojAwg+Uxbx
M0RGuCoUt7PRvkMxC5+UTEBPgRttIfateWBMn3sYU6ZS/uJBy6d1BbS1VQzjtqsj
zGJR9CCvRi5cQJcvw0nZ5m1oyyZDpgZHAPMd49wU2uvgV9ISn0+K6QJz2F/CthgX
39r33jhAfjXFsKM5BskHNxIYJ1nn63E05xbLMld0bP3QI9M/exttFD671rL42Apx
vaMlrGAU88EUbG7PjeLMwcxtSPj6VSgqaK5p5z1zYfIVEsLfR7efoxoKRT7EOPk7
C94MVY84RP7mJexnW7RuJ+vIaoCjXvTdAPdjJlLyTXwreuWIY92YoPWjHhJikgO7
C2ORKdimt82DLCrMN+08He+N1tDptSODFaawrzExGKplhgADGpd8h4KErSUvNX/R
50j9agaR3HtMm1FrsjuaczQPYD8mf1NftYT9V2SXF64=
`protect END_PROTECTED
