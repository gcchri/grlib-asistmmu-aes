`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLwfCY3ekEKbUdhNktmPsaXWPJ633UcvEp4skh9cWV3Wmm13S+CcSY3R3p6pdHTl
h4XVXZdm2KzoY0gA4BVXaMQ7Dptna39cy/bidtY+e9uP5vvLE6DGoanWoNd6yib4
jMMY95fM7/z3VNQsM1jRJuBxQK32wJ0jEYKP7yUh+6LoEp7rAy2VIa91h4oG/dZJ
14inAVvlIBK2jxrVLbgH2Pt4PABXAn71E1GM/ulLwDH+rKGT4HlD+MxBVMExndfI
2QVE2mrFPdiam1FIMri4JyfaUVY+nCtnl1h8JQbvFtITK4UUy87tW4fEOUkLUlwM
E41M2W6RiPBrFZSLERmPv1CHkUKE3XK7PhTjS5I6UK/yW1Fyp1tz4uSZmFxjKgEd
e0oGAKFnH/XlxJ8Qy4LLcEEVs3srZbHioXhGWYNEP3accyNcjme9eHhhbdQt8WL5
omHN1701DYXlsGYuhpxjEqc2Eo+4RCgqXDamO/+uNhlModTXPoZh2eD5vxqQ8BZi
Yvjqawk3EWyUI969AwYsAnFMNiMZwRRuDnkTHOzbmHnnqeB2a5F/HMbXCo68fdrO
M1eS3OeSdc9Msfu1h6bfNn9o7Rffup23JhtaWUC/q67mfh7ISgDM4o3vTElqg6nU
1+DqkT2aBEUURjwdXmneynOw1/bM5W51v/oVEDC8fdQlceulVrEtQed22mQCiZtD
8zMIyuGbAnZ4pkdfKWWcoQ==
`protect END_PROTECTED
