`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKCso3+WjoTZwBRWIhqfRDcHwR9aO9D+h8WmDXdPDTZCXgMTvCuqEtKJlDald2EE
2kFtglUaiEF5lwaGP7x4sX0mmbgwTVk3etty437gxogeCb0t4dWi/XNG+t86+NPs
mYuWwSUcQceflHciRzeX/+TbPyqFuApVwWDATbnTNtMW+v45xqqqvc8PuDAxUB+i
Bn2n3my4RD3Vu8gXvngMrd+/f0f2LS9ScqrM6k0XktlXKSVV8tzgRvH96nY4hik8
OJe6a27ksaWPgOfmVrO7WftymvAysudZSbjg448puop8486Zr9wug31NEhg2+qHp
k++xaV9pR3pBbGZyq3Td8A4XjC3przphLVT//T+YAu5EG3s/9EPeNSQFvPyQb4Et
9IfL16zPH58UWwUULlHpqshMRpeu2NCzfGjy9i0G+Z7SXZ8NnhWh/jpkrSWpqi0h
u5eJXg1ztoPfYyKFEnImLHIKBmRL9XcV3L9PY+cvKukTzZRo37RBVet9QDTikkow
EBeDIGJ3yoX7UHJgA4+CXSm3pvDXlxtvDYBn3FB/jQfSI/1V+MBHxqINTopUyDnJ
VwsYqYjLeIjX8vc2ZJcSkCPMbDqg55sToXUyRbN/6xY=
`protect END_PROTECTED
