`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dkn4bp84TJ9ccUYsQEbmdE4E6yxonYXS8NHPhBFwougRsa2M+SDCsZGfWxH/3t31
9EEnBabEBDumWrb83A1Sm/NbO7SoyHWCsLpsjcfecQzLDEUFma/C+pL1huOw1Ynu
yaQbFDNtnXzghG20dnAXBW7OYrFDtZlxeQfvwxlzD3JqNKTZivhWpRd/S+hHASgS
vLvgqKJ139IlTM0icGeEud0h0hOoLqzzXcRUImUxf/0NTCJZAPRLmonT8aVTADY/
W7eAi9LUbKeSgt2nHeAjxhggQNTFzShu5Cs2vPU+2VSPufL4uCWaav+cDzzql4SL
F8DqyOeQjOPWQroTfVRibn0uPQGeIIsLoZ/HaKkpv3QTskK6wahynOETodoaYSDZ
TZfCAnsZvtVPTC91sMoUcJ/uTmdjGGdk5hpRO02M+NGBHmjs3/PJX/jRHdJ+2d8h
nGZQcRR5Lhd04l8+ZCMMpx/ksLYBDueVWvQrDcHnVss=
`protect END_PROTECTED
