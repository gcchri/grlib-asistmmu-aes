`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B7olFHfKzaw3QOL6ZA7rBVpNODDooLK0DAgIvAgAof7QjwnjoIiYRgpHebKX0vT9
D/wvBavTlP5CnPcSROQ94IcM3Lf1i31HUOgpJEBb2VSOfi0mjyZUiqIUjNUT/Bxq
wI/vtR270Ya1iYM8TZ5EHx9IahsavCchXdVIITz6pRGnhlrbdk4tzOlQo57OmCMf
GPTAfWiOSHNfFAzBccJhC75g5bn7tHD4zVAWzoSPYenJUiS1C2kSsx/4uJp9nOrl
5mCCNrpGWAltZ+W+lfYAsaTEiqnbJN4mhGm5075cWqMgH0UgspliOsMRUzxzA/Iy
g6g2aspH2tJyyRCWJkpSQF2/yHw3gplkU+yWE4jBdkjkWa1dWqqpACJNCNRGitJA
ybL51oZTAYvvzBKPA8bWs7JQ8heCRuoA7i+j7lKoyyl3HfF6u+7x0gFgc2ZaCZo/
5fUR9HLFsbH/7MuGPkds9ipgVP+kBA2AghK0btQ9ER87CinediTsArU6JIGtLcSS
zjc7kz0MLXxZCZjUw0D/m5BLuVfAWppnyZBae9Rf6xNkn07y9FM7dDIJ1BKcsKZI
4W0bErSW6tHEB6xwX5woMxelrwKsKerb7Xy6qlfU6vFDPSkrtmgh4h9COY68lxFH
+p6edbzZaswtyiOKVDS279ACpRN9CALjxIkqm9oiLExBDfhnAVUsVU9dZ547SFa4
JNSGDAY0vIcvA83ZVzsc7859KJmyNrnjGdAjWbo3ARAPCNmeCncCjpBFP0hKeWvJ
HEsCJUJ1PmJkhIThCSG+WQyueEMB7uHCJjAotYsRjp+jEKLr9H0pG0mqbFQkCdUc
MVNs9eAURNkKboO/VE4mBZg9ihAwI41V2yYH6qwjxPrP4A+JScG+pneyMxkzWExw
5FTgx4S/1T1eWbwQQhZB9VtOaY6Tzi8JfhjJoGk+9P6adEyyopOM8XGnkUGHtq3x
`protect END_PROTECTED
