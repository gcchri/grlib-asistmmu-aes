`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AtuetM53a/argyM3/11rvKW9MOgPd/HCHKNeh235CqkMvyg7doquHfcmlFtgSo0K
qQvB77b1LB7J08zmYgu7gqN5KtbuJkatOP4l9go8AxHA1Peolck/UxN8i0hm7mg0
xWJknGGgG9ZS7vWdus/0unbY6vufCmoXFJQQWzihm+af1S27O0sREbfdC9heW9tK
4KLqN0DTKMxiRe801pRAYD/2jPVKy7a7n6IfgTNovDsvT97VjuGqFul5qk8z3V6a
WNIIyiVC8ZMk6awv49Bw6kVzSldBwXz2i6hWv3n/MvuOpxk52m+yLlex0cnvmx55
sauLOlqECmpZKkzipCHFMHJKou4OY+/Dq4iEarN7bbrVvtrEpjLtR7Zk11O2Wbak
LJPRoOkxDlkCkzNudtLAGgf/PoWo5rheiwx8lLaaawHqAxJJaRUlDTLwjuNMuov/
k7U9QU9GVwRFsjMFYlYVTtjlxYiL8uqpP+qyEOQmxuI=
`protect END_PROTECTED
