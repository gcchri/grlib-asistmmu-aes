`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQY/ggcPV6jgLmz/tTN9gsyiNH9U0G1qZaTbAQhBabI6paPgApbnB+Xz2S7o74P0
4JLxY4PMcRQCwEB+igK6koHoIt7mfSxZZo2SJeh/unw9Vxo9PToTMxId8dZ8p9tE
nBimdzjOjqFN0cELCbj9R5dd+0JsZdpinFzWBQQjwm5ocVu/AZweHtQRcqTUA3Rv
yZOOC3W5FGYDKivB1g76WNKrNpkoXHIJUqef1YdzqRnfDWNrknXFjwmqTCxaDO38
y5Z15LlyW7p/dLsSckZvwimqhnoVRu6J1Hin7b3ES0zUE0rSURvBNKbuhQXbn+/Z
qhPwAvmPlsoWsJ8wZcNfaQOYOOfYKUZ6xdAt5/MYtnqYtk9W6fT3z2GBwettyFsD
+arCve8nSh++u4vUlad3mpwBtieUZbR4mbCnjXbPnyTU2VEDXx9R9aS8UIaA3+ng
NaJsTlxvuMEbT6MWT7QuluSZ+aKqm3Z3VnskLPgqDlhNrTLmPR0FX3MAuFsVjbZ7
OAWYRDgpVjCIBlJuKxF5YdPgussJ8MhAJ7UsApQWygHJ86Whg4WPNXuHvGj/p5Nn
glOnKunjgpYF3mJ2bLx2VXVkIlsaAvePoozarjkjKAP1PWIwbbi9+RTxJNEQEe8Q
Ehu0whM1i4uoCYPuJ/D3hkmJtHJH31xxe6VzxN4QKEBL2a8LX0gCITTkHFTda7us
4eFuK4QQyEV72Wbqjykyh4xv01gVEW04o7Ha+dp8eTazOuifgltiC7Jvb2OvJa5/
WGP5iIa1+hRAkytNeFCSwzLYBkBVdYQO5CKhi2vcqgSUYviIRAyTIr8p9sE3qgdl
96O0l1PV+14u+SPoyIBTU7/rz2ktCN2HKXVZ3wRZxOpfSDe3Vp9mniG0fcp/S6u0
Dd9W+zKI8pC4EBK6e5rbIoM1dauVJI1tEec6kc1KIjzjgk28Iq7wkulTj50A1PRx
7yrqTPzjPyh1Tm3h5TV5OMEluakwejVCUo6mZpBoQp2cc47UW5uwoTVimRT31YrI
vQXKhIdgYhL9MXwfL7AKl48pXb6vuF3Rdwj1Qu/Ca4HbmGAyPd1YovBd1mHqGHeo
7emaTrXjMwnPVg6Xq+jOd5qymojko2lJdiFHLM16ROZ9E559nqlKoDhDqewfCcXG
VLISUniPqNRdDrknwDEOZbG/hUBPQaPO4zHdRiNopmyywrK4zXCbQlw+II4NH89N
K6d6NVH71Czv1xAIwpgLZCh9+nQZpZGd/j7BLqHOO1YmwbFxnI+DjkBCGi8/WkTM
YdDrJFzjeAk1mXKfwQDLZjskOj71TOu67xXyrEXd7Y3jCxq0sAY2rpe3B7/rwJIN
x4EC7jTvdcKYIVZpJ1+TsSjtwD7ZCBJSZqMVaM4v+nC1v71oj4EMEtVB1GJQw9a3
HWZxwV+dgVSmNKWsUtSEBWKEoAD52m1jd1TqQZzp7x/ghojawy9NvnPzVfZ0x3VM
aV/ciuBkpvkXWsPKMh/rqAjZ82jbVVVCj+2usMqX1t5mB1E6pc1rS5pK/Nw3+09S
WeBRuDh4yK+jv9dsZqfJ0i8AjMC8H6YOACJEpKbVqPWZGoy5GiU0/EZwrxYFoCHZ
uU7fKLWbsBzOQZaZSd5ZdufcPTm2nO681WjkeCyn1P3ymvmNyaDmeYsB06W+Kc3G
vcK3aR14YOcR6o00jIepASUNeDCvdBSquiVkytLnw8OzAmwg8NWyCHERDuCCRiF/
EWYt/2mbwDrsknFlxpVZIiKivJrnTOzazmipThDCb2lGc7qJfBtzaw10NFWI3XEn
clQPkyQPiYmogEXfLhNhfKMuhXEhHV4LaDL8BidzMsLEQCAHE6arVsSFyvUj4mtl
sIFa9RKuqkH/Ol+Zu5foOWJysCRdhHr3r7aBQPdJvS42BQgYV6D2Fx6lPpx/OiTS
pM67WjleJeDib1xShmlF61uGFzY4KA+RrnJBTnJmfK50tItK/cc4AckERIMw4Ggi
7IV03gVFZLCZyIwpaKo7z+iQ/XjGb/XaB0IlNfI1QdS0yhTo+QXXWUJZ2a0ZrhuW
SvF1kMc83ABEpBBIVqfY6fcy8T2T7ph13rItNuKB8iFbRt3TbiuaTe/rL6mLMcWP
iTLXcadklnfKB3QC2U9+IBKQofJryTnzXHon8O8SkRoylCE5bEj52YxQy3u7SJhF
h+zt65chN5tdehNPvySYfR0Kvg/t8ws7/DceP5t5RlV+dmgJYI0G0NU4cKxwo86m
jRZo55lvmT02Yfckqe0NwC81XrBVXcd3OOJXxdcaFGT5JipH0y2vjD+2Fk3aAca2
4NHEJ3XUfb7+Q5fugpncNJf2vgu2lHoIDq3m10f9b6qXav032MKkoQPs8se4Hk/F
9ESdvG447CAjX/6wQZaSjgcR+2WMNwSP2GlBY1aFszwZUR7ajUHgmz1Hz/63zehB
C80vbmTk2LJb6ADEGsLqbHyUU5YWVbmxw0jbVElA73HRkzcbUfGp+4BlN2p3MBSd
a4QlUELgT3gnodRBJ/7QoE91W4Og83x0bnSGeTuR6L1qnwoQ93TvCn5fVHO0gshZ
5pHW+ElnpZi71AKwOC5q8FUJik5LGyEE8/EwTYUPMmMd1jOH5tQE9sfZ1oSlbVkL
xw2NbCBiNDVd7+JBE+ihlLYFoAKEiFGJ+CFlx/zEh7A3UewUMtSM1S9hggzQzWFq
qXeZS+9v4OcaV3hqgZchsfWpBu4YIMRfSb+BNE+lObgMiX/GMeBxSH7bRYf9hryD
38Hxcy7mHHLNbwrYIS/a175HHUbjv9pfoJ9K8bWgU+uu2q6hSM2Yv7f3XfGL7roA
r7bvKsE9DMoilEedJmSpqhzxVB9r1qmBSGhBvi0qIzfuV71LoCmgijVwKZ/zV1y3
HpWmuhgW2Ja3SbNVSHpg0U52tuFixQpzdDIo2kyXnGB8Qt4wiUBW/OtO/0XTx/Lb
Zp5R9pB1zybKOboQwkI9sXSgvx6rjYvfkLjtU5Z5YvqLZ0DtVDpy1reJgtBtf7Z+
RE6+b7DO8vDqLkhnd7l7ag8G2k5cpvnVYuJqgsCzZj58S+N3r0JtUm+WSOL/cfp5
wVfVAx9ffuWXQdHKaBPyyvn8ehKywAj+bJQdhzgGstJdEhM9X4uJBQOmz4j/2MQx
fD0aAb1aIlpcOywNt6lYQtP3naZDPPUatyRQzx4k2gOKeB9fvVKlydAh7AC7Rv4s
DGt8fDU3n9LqrvLHS6DrfUKahLzRySaLHI4P3xcvJm2Bu7jcQWDASocgH7J6iSBy
BBOxL9lEFFcGivi866GkBbLlxYxiVFcC3Il2HO9pfCCDc4mkMJgYuOmy84wqYF8t
33calvuMmjOuTH0vKSuHoqf2JWr8JjM/9ix0viQDeqzxGojOw6972uDYWfml8dBI
UukYDsiHjKk7oX7ska2Dm2Zpk8ANFzFOvkkm1mGg1ef91jFZkbUyxjtF1O8CkNGw
URs0+KGKHg1blqu0e/vNFvyYQMxDd14WwdeMYrDGuTc2TdwdYJ1f36MvJeRuP0i4
s08zcfIsP+WkNMWcCQUq3YTE74LnDmHlwKtexTWhl1XQsdoMu08r5OHBniDUTLr5
kjPOdvNxyslGFBlkohOJFfibl15G6y0oYqOo6lKy17R6B564YiiLmh5/bsy09Yo+
s+849GZueAR70EjZq8K8THZmIIOisY5bghr60kVjl1BxHUMn+bM1MDdDaSgCtfQE
cD7283cPoZ98svh5BcLoIHXdNI9FTIx+aIlSAQT3sJepSVzFtQncy/1cymTvFWKT
6XI/TGDblPwAMLBTH55zjFFJVwEjKo0GbLg3UOCXypmAvCEmz6aGIVv9rYDBYzWE
09uTyuCWWG8fNB2r+rW/P2rJQPzN3j/xDkdv8B/LhzsSiq2UYsoEdQ/eh3bjXze0
VrQtX3KtsyUSmFAHRENO+RttXkMOVepX+jWJZ2XsD16zyWqYmymT+Cros9Fue27z
vS7Izno6z8L0w93Jnc1U0cek+vinSZA5FQ2aSmKAcpq3fAV3rdPVa95NfX/YjzXs
y2lO32j3JefURL/tcCwzfTZYEYtGeViqQfrffDZpLuglT/p9E+mO1NbDFsX6aLVz
Jger+BS07RPQvXBZVGX6H1x35vtfgWlQ442IpyhKV4NCvF1XfvC0E9RlopW9avfv
BNi3gXzvsBGzf4ZynPWdlXm6VPCZqqE/YV1pLmusIHAqhYWLMpVVPi483MaqPyU4
nZbKyrVSMtCrXaNKlfHK87dy6OA7aLOYegNOinHQZX1ebbUNDQWbdM1S/7nFvXLF
S7PwyefQG0JsEOAyqlbpxG3B8UBTWfhkXAmrMJs697+OEBW2+crmui2hqkNdXv9C
ions+tGWUFfksPa6OuxDW2FYZbVJL40Ym+JqaS2fizBXui2RySOrcwxpe2PI+65/
1m4z4einuQZj/rxBen4psSznP1vqnKAtTv6BdCQRcRbO+sK1Qh+EHKz1+Da2e3Co
leCMbFA6HolgAK8RFnOoFszE1i6NyvAmvCUy7//V3IeIq0e1gc8rOuh9VaP5yr5k
PeIynIEgmegBvToaQpkTP0AobPpJZqIgyFop5JS+uDGL754aIzrAYN3ju3W8RQWo
D9mmw2hcWLup6hfMmWqk9RdBKu2Eot2aoYSuk8HRNFFImRJ3LmJAa+agzxYsd0tH
0f/7MU/gvr1ViYbqeOFi7l4krJtI3rjaQQIscSQjpmnuoof8UpdBSYW4LN0FsQvk
pq+kJVIoutOsrunCSqIq/GmePUfAOVa3+pQylIqiVnM3h1hA+GkQFJ2XW0QP5e1S
9fxkZe4vBigIdNIh3zextcn+htNEt8alaF7F3tRND5ktzd7BUU2lQBLs7YSlbV6t
H74jaK/9VNpDPGTE9gWFUULpGcbk00nAhitP72xC3/1B7D734ndAnPmpJEfxyOdL
z4Qcgink7JewlALAOjO6pp9vdeFQGykw+j8W9z7vQ0AsBP8zQKLdLCFmIpIfEQwC
o3BGlnkGDSY9XWWYRzNs7BTFbAG3fJT5sYZ+9SlnbLeVnhZO4YxCICOg9u3iaLoC
GHfwxw4URQ1H512eKy01bBYr/US9T8YjIPqHGCN4IFfx2VsAPLxNwYo5vimcsI/k
HatYM00af/MbkrK9vBEaUYPaU6nMzhEBdqoyonYDRx1zXf31OQEOa538KQgHHm/+
WIRcCBBugA+PhQluG1fbV0mdogybtZ3QwoRPAjIl3Wr3N4cPClHhpc+MppKF8f6C
xjvVEFDqR0w1dR1LniNrZp4msyVOtCXhhRX9aVZYRvaauREjl8BzGSkuH25mFkfV
KVk1/8zft3t60ZkV0wEMmap4zpovmecGhA0pHkOYIeTmuLwrHa1WG+bRaRdJivoG
+kX0m9PRmJJYoyJy6LtdqMvaDJ37VR0c5dF5Pjw9Fqe34fUtRh1hlf6hPRjk5w2f
/7MT5FFYhv8arLoplb1RJ8mYplZhotXWVp0CQsZYFMnO1BBihpxl8hVOjzQKsAA4
QS3ZtDwjJ/sdqZjPo0RA5qf7mtuSZ6OAiGxEflFuUSiZLqcwOOonnOSO6P8Otgsv
d0Pi9PNhJe78uxsWMFnR7Sz2UffNRvnOCK7dc/DzLQMuLDE5RQOArP2PycV3UhW4
RDhJjt6O2uzVWeu3q9ZL/4anrMxDdqcfEFDGhEtKfBt/303R22OUTJXbp8PDQZBn
BrpCeRRseU/91YNz/mOUqtelcx7fZ7FOHwIy37+NpKouMIyAUh+fhKioBgwMpxCG
Ot3HSdcRv+XNKBdPFgY3jmopZen0FaPSFKLHEwRO7N6XL/hu/9Az42KQxhwjq9Ey
g27He7lcHTt9IiTCLFIObjGsqEwrzLQL6nGhWG2grY/8iYhrqDuU2GtMtm4Wv5Qt
BZTalwtnoDAwz4pI+5soXbHGy/JznYzRzo6ma9Mxc6as0UI+BFozSFuOwlEJJVEL
rI5feKAhCIA50X/KdSV0RFiMMimc4cxZD46fZAZeFreuNcStMvKY35maelq2LNTa
cFPdYNkMumMEBU9Z2yaw4+5WLW/7M6F7gu17IfMMVsm2/wJl1YJ1g6G2lCdogQex
xL+peY0f1gUIf+AUV/ddiXUyE3UJ/MINJGEngyFVtOU8EUb3DYsLmdqR//Cbp7Se
NJEjyJjme0ki7pGjYDI84NgGWWgsFws9WerjiZBLrkCHcRl2NQQIGMMPns+L1HLV
fSoQXboI5k6kHSmqxNyCFtxUtnpGioirOddL8tZgQM+6IWSnOSyV6EqLixFgCSUR
Z0s+E1H3CaneCjw+lPrT8xpejO4qXFDbMk6jIWKcRh8RVjUhadBRxxW1OV/Zi0VS
atisSpYnZAHUE2Zzt1DARP/QDSkSDr+et6+aiWFHOzZY+mCEoWr4EzZTj2eQJ8J5
8isKkrzHwd6v+FAuuRf4bZr//MJgPHzlruQVbICgginJmJKFpmIORD2IB8Z17hJa
Y8rD3My97HPExkcKJAcsj5B2Zdft15J87tZe3SOrt3osfE4k6ugopPC7lwecgKr+
apw0pXfftgFP4g45t2ZG+p1RqOXDJafZpJOLd24CntSItQHEQVLMYfA6kShU7dXj
F7tbG5E8wRsPnYRRcadgXrsNUj81xmLQAgnWTms4iCV0awUXWlDfoz4Ob9gEQfBr
T52x2VnhcA2IO+S4+d1OmV0zH9h0siliY2K8l1IDVC0NJhQaGFwViGY5Z7XhvkDx
Gk9zTroYPNPiZXIZRO5A77P7qfgQCKDYaaYGjTdhpzAmL/0JuTPgFaMi+pjquqjD
U4c1YZwbjizHkwTIazHahY/IzgcylUh/ksOOvyIV0FO8jDOhXaQzQGkS9zpYAFoV
WoBCATQisIPFJD+6E9mFev1tCYL29gMu2noMyJ0mndEzuOhp6NlLKn1GCu245brx
a0u2L6PeWuixTd2gQlk8m+7fGEKo+v+clrWfHHoUuKGOOvS55F+qEWDLOnGOTy7j
Vc/AslbS3MROOvDmLiG40T4zxM8no6miezSs7ncikqWtRrOELyz787FR8YMg6jrc
RnompAtGQLT3Or1aRbwICtBgzk4/NgQ1ZOhnF5HtrN8VY5LBVQnWoA25FS5Qdbv0
LigeZ1B1yzC04AzE3xeJTKhrQeFklzmQ7r+5lA4E9z498VbgcdpUTw6Yp9k7Xt/T
NIEKHSPo8a/TcGt2AxC7C70+UL/s+g/EjOKAR2sniRvZQSJHQdVnY7kFRom7eLjk
WNQueMaOVIbwektmD/pwsHBAAbC8zV1kCsIrvbY6maN2GsgLhn9N+Hpvu+nQd8x7
/l4kHBCDS4j/xbYwvoK63w==
`protect END_PROTECTED
