`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rCrZKmQeKM6PZ8DNxz8QH7AIkP5ZrNg5fBa3yXLGqhpxS5zAdxZSOB9M15g5HRLN
gH0s4UZFzm6a2SeVEt0djHBmX+q02QoJd7ZRIKYHFSGlEmiJLOretakthkHW2YD2
QrsSrYZ/Uekkh2QAW9fq/hJE9N+YBweFMcAVxiePE0pJ2j+pRZVgj4kDYVQNPQ2q
QwIBe+06UlZYYHXo1xuiPlbT5SM3bJWiUId/TnGKuGqKhDi7YbYuQPIzWcthDPfl
SEmNnu2oxcuZiJTP6W4DoNl5/jj3TwP/jEgH5kMRHt3tUdXAhpyfX7k48ywDuvYF
lQcwUVJcbtr4x50j5ssPwhrQ9URw1tVujgsXKNK8xo6af9gnN+cIwHP0W1Z0lMkh
BN2k0O/ADHt8nLgdABEbSAH5WdFFwCBCMmKipaiiKYcSAK/tYRIGl+LJHKw6warD
mC15x+BmnEbVw0sYwfJNlZ2caNPHtJ0Nn+aHYFF8zd9TGje5r0IHSDQkKfOlg73k
77JDIuYP4GFQOABYW1SjPEJiiqWC5Upzd6EjWchCTRY=
`protect END_PROTECTED
