`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bXYdN9iKSXzSEGpvX9fpP0V+gASoX/1Fbc9KoKRMmpw3KOdpNuM5X/4r4M050yeS
0kE8sCShKvSGyTW6YfDcjJdKyQp6JIg73dZ2B9xaiNm3Y0v6KkH04YzOY2oHayMi
x99IU0Sq6Lay2OL1IJIdTEeZ5v07FfvmIKg5iULcRrOwr89hRsmUIYn7MsABPPWY
0/mcG09nMphf6DFaqVlZQcSmawr1dYinVyXzXrWLjnfCNqIo/hGbN2KVmr4Mil1n
1pTYo7QVclIwlr/5YeuGCU4C0Dfv3xmhiwBjk8o1OBfgb637H4pn6bZvlI/9aDwP
VYLPDlEFetEobCdVWRRbHHsTyI8+544aWJ7XB+4abYbfqSWFGcus/9PxiJjludLY
2gDgGNkEax8148DUh7TWoXdRrO28wmBYNU1NQ6GLSJwjbXgeypzk/mx/LPE1MA6/
a7n2zY6pKVdvmdfvA3Tu+/kDyTXpixn3hvr6kyUNJUvY5HMINJuU3Vo9hoEohALl
yOsYdPMY9lDmDdRqVfDz+MJpFNFNH+k9rqpBhccuLAH9bD4iUyiI8ZhCmBowyIJO
Sq5a0tMuEhVRjzFVZvy2kldEmmEl5sBwHMsyERajNC7bB0ELafIlCay6eeE7OT9O
NEx16nLjh5CWms3QB46+N31fPKZ4gAG0zTDAClGB+eofS0PV2RsltAUXuXcoSVke
f4bQcXfdTtaaKPWWj06ZDbHb+t/4qf8R8uXP6sY4nek4HAPvG3iabbbq63vFrTuM
FgWGv/02d7tz1eMw5MzqENxsRzCqPOrjOa0wDliZQw/tfemGffIVBGFglHDgBd9Q
oDJFm2/ofjNX5jS0DQM8JpzNcvbZHbkORaWC6iZz256oqJFawOWOLPMuXFyHY5i4
UFqBFewb0dfXTHJc8VMbNLAknVmc15Po6UvtbrsDh+vSYrqp7TJBT3ECoIgUHS4S
cJXwZALcBvqfgNI9AUsDyIuSxDEM0chk6NKjciZOH8h8C5JmezVyM/4tR7JF+In8
NcQloWm6nhcxBGqf6p4bKsgHjuU8c7D9pYxvrZBAmZdollf9Wuvnt+hxFoBZ9mJh
1eiy3o7QDzMxwa0va4lI9NklMYe0ig0uMtzIi8CYjz4gcmcPDu32fm/e6EmisBMG
jNRnRHpA4qqYBLYFH4nf8s76GznVMveNBIVT+uhJh1vJNpIq6v/atmTbPDFOJml8
HKSEua0zbJUR/CbeUl0GUO4OZDZpVVRtVDJdU5aU/UTS9YrjtXzM7tjR/SCO4BrN
J9RmLwTtsev6DL0P6P2vYZ9eOqevYgui6HMuttpEjfXdnyn6NHSgxBbIAPeSCRMS
ykTG1OKtbzXqUOscQruUeACT/jFgiwvujFWCnnzAyVGznKBzSJ3d6EH/XHq6OdGU
fd4ouFCZJPpEoi7lhHT/ljWi5vyVb3rbn4Jw41eE9DE9pTAuyY7XBHqqm8Ev9Qii
KkEaobeX8wUbHZQ0QEuJzk6n7CDgkeDCFWGizzixIUBdULZPGN7iUCdjcJ5tUWgI
6rJxOh+6B44xKPZJXs6hMOKb3/ADC1bTxtcHvVRD2Y47PvDzqppt8o1g3ve1UYy0
6ZhdNuJEpJqcN8Lsepi+JxHPraOMQMJR78cKlDWNDjGIuF8scRhlQpdPjNMDX4MK
1lUrjDDmAafaJWPbTmGuQqg6aRheSH0KJ65oAbC74nzA0pTT9bYPtnSIpsTGjgu3
o5XqmGd4jP87TAWEPafKYFAtigClJ52/jCz/ngy7aHfjuf3ZQ/hEeVQW4Ity+NT0
+h7dPriYqfHLjbP0hQvnW/BEvJTBbGMiaLrrAzVDNH0JNlFZqhIF/cFkgWyYniyJ
PuLDgmpi6TrQso95TUEXA0s1khHaiKvLUWpmHshw8y9p+DEkEl24fZIVwFWdZPmB
FoaHvITfr/lqGA6uk6t1KOX/GXJ8C9jaV6Pib7x0RQn7VpD1XRuouARF65umlmx/
oq62yaHUgyASvYZ5oyeNal83KVDQ2XfwPhTsDoI2AksjY/CxMkbgL5MJ5/X28N9B
RMJPpvGX7uZer3Kw38zNs1BKNRMWXajQZWauIwfHvX+CVb3VyEAWEgJBZYq+AHjI
KvHkO86tUi4Mgh59HA4FA5Aj3tlrJyhSqt2VqXi2T7Pj+Hq806rWcnzinLrgdUNZ
b5eRx4KYXCHuLhDJBxuiAEYgMyuUb86RM27Cwt1l/zZp4uYASSj5UvuBiDvJTTyG
laDUaDTrgpOjZ00VD996jzu2GBkBKyrkg+TrjOpj3/XkLRJYNMgUCRy8w+sD2M8e
S58J7+RRacYnKtfS0uJ9VMur2mqc1aBWQZ3+Ll7LDckDlm4D6KGoys0h6TM10oAX
B2vF0Qd11ci+F6pFkrZOelwwcuJRpASThlvygVFLRcw4Qtqdaoe6ZHbDj/kCCQEw
evsVXOmm4PCfv2CMtGNp8FHfL5vTT3DHq+xjg86Rpk1jvoTWi1KyFTwLidTaHKzu
6fsm/oo9Zgq5kMiO81BGA3KgEFlgR0kr27HAy/cgqaAy8ei20HTw8Ch3wFrZJyG8
pAsdZP8pLw8Zxx872zIEtO6CPc0WC7wWBZXbe7AmkfM3EQu0DqSe8gVWUaWM7udv
8ZnnTIPsggYLU080qPFV2HoqEKHHaz5G6vEF3WPpT51m/Bp8mTFTAsYZ+cF9WYTk
1zWL9sFj4AQnpSeyrTV2oQI/z6Dix4iQ0TB9IqbPvkpzDDE2BGbqitUgubj8Zokp
Bo7z5hEOSr43YRV9WuETsrtZn6KWC9MgadokCmRAKzCAYkjBIFZsCm3+ZToFGEpF
VGTK+KsXYvpoU2RZdqyN8N/7XeZK7/Xa7vA5kheez5lXMiaZu5Fra0btXTHOOTdX
UeB7vUW4RlaR0H/d88E7bh2H+LgqpTHZn7a5IQc4/5ol3zTcswsw+XLh5o+eqm2w
LFObRXao8CoE2BXOsSxAuZGEdE49PxsIz0lsADiklxc63Ck0J42M9uyiafOYH72f
Fuy8+VLX9CklYi5OWHz1STBKrc2A2AoK63jenZZznCq7mJOJfAr461bSHLr8ze9s
ywD6YXJZGUc01VeagYKTNWVfV3U1ts0qF7B7/EwB2kqzRElxA6nza2LH2QvreUad
j0U307Ol3i5vtSgnYbVWN3Rbi+tVC+LWyRiJWcdLUdArD8pEekSb36UvMll2TzU8
z7DvA92sxA5wTNZ6RFFezp712cHsdbdvacuZVPp180sjosvVrCyx83f8fuCH9Hpx
1Wzk/u7U9ySw4nKHLru77V7vEg2yUDiqCSEitxU0Yw39IrT9+bEiH4vu3mlwD878
j3P+BvlV9Ior/vV+4ma7dxIz/LWj0FpRgpV9ChCVcE2wj7z+0NkfLFp8iqJ6sO6u
2CHdhil53JnQEpAUn6kQUUjiby8IRJ6rpoV7K2RmIXVaMWOcCqYuwxGR5H29PEUf
5D8YpLv7ut7I6e4Ea3jBhqq/yeM9a2mihuyZjUXvMiCyP9LIjIB33kUaE4AfqLbY
qeu2ZlqmvTNfKa2vBGG+fqU2FDzwllQbY+ONXHQ/NbAeoXUb1zEC2H+oHVaKrHD2
UDgfrciIAv7noDuSUiG0IFrT+iQqtaPeKf6WgCMMxnSmwdWZPWLG3T7Y4vmyZgGe
zIYt+zPFvmtySXqlTE6J7cwBvjGcKF7aKp+3Rr0yPLwTkErdEETA2KEK2/UI/eVR
axWYNFCGkDNA18HteEXUFKhedaYZVU5oeOHss+oWhEGHfQmNrBOuvOKPHpkPZCh+
EY4pmSiq9QQvQM99fMOn5AcPii0msfKtOMOfQ6FAr3zSESJhN6B2c53sRTxYXJj9
ip+1j3IwSRZmL9ITEJZffMPQzAySbbBwh6KytNzviRy+NTviFnnbwGYnBXvJZqdJ
JjuNn6zLtgTHQJYz5nkskb9sUoNo20u06lssp7DnZrD+KC7e5tqw+wr10/QF0Koa
bHd6/gJmoPaIWu6FqB9ByN+yq7vwKHb5G5KIicgjFI54LKqcFSeJag3bfb4/whU1
u0etpbHjtY/yNrdSJyxIshomUqFG3Eb78W73u1DODB0Bw8GGLHWCc0CQRkFvgfYw
z1vFBLqnJGX0Ea1APqNRv8qAafIEgp0CwgLxVnjazhNo0ZYp8VvytRGFYZVh+m8M
1xOIbtkyq+SJdabQDykjSbQ5yCdLYoKUxgsF+TFzyW/n/oWWkwk5tOAJmmWcaQoC
hfphX1RbQcig5iErm+r3YkB+m59Ceg7zvMc4d0bXq00i5qyVHZ/aO7wUHvNvNYOh
iCoZrsDJ5iF0u85pazwHaZ6xaOLKLbIj6+Zy2Bq1ShsumbUmhQO4ZDGAqDRZFmJB
k/sakRCI4WhsHA9pdnqYRrLk1BbdH40uDsbNbv1tX2ftzSbv8QIFUSPS5l620vDL
monKj4kA29dn2RZaAyDQkoRoxaIUfqD9mXyqExe/5ABaanXOLyuJwNumzG2odYs6
7l+Jci5/BkBRYLmlvQ7OlscAnLQGOhpnvxVt2JLfP0PqN+tuXgZX3RkoRgO8B809
+msMlhEaZ6aAdkT368efFaWCJV38QIprNDqGb3cqLODGEdE6HBBx9RCPu5/tSqf1
mgGN+umk1vpCowiFIRZF49MfrK+S/G3R35ghQSn0NBqgU35AGqC07IBl73NVk6Va
VLOv64Bo/ryZIMMDUDtpz91hzKDLhzHUAqZYCWM6vNLApvQCCTJx/cY9OhWe9AKH
3MgGFHpFABdnl2xHA6Hd7QdFePODDTfsIHDUTB5tDIQBiNqVrkJz5ICEyNKvZ7V6
X9XcF+/ZX/eXq368o9xp5I6uUOrZrYFAJvC1+27CUtLO7mXnbRtss8kmRl2XRHgP
OwtaGyDDtZ+1olSHLBVmkmbEZ1J0rdVrKjk2tFCT1ZD0r0JSn6ZRpUvZohoQEFV/
a5vqMoMzEXrsbFJ2UmnDsVefR09cQruNRjl7sPixb//IEf4zpVkQ3zf1OjI5Yb5p
9/rUalslQlOLGxX5ZUOjoNSGJAJyZwm6UPrfTnHLcE81jB1n+y7jMDaDSpAo/Wie
Wdn6Yuj86UiOlWTJMm3uTpaY5d+NouATPIx27RrTteuwKpEx6LN2+Nveo5UPS4ws
CTxoVYLbJUmzb+gP844YmvE4IU9d9KahmkPx8ebl2v8Q/j1hzLyuY/PxA23sECdN
L+vwzD91F7GA8XrlY94O5VZFVVsQI8G2S7N3FJD1IUNp7mmfqL/1u4TzQKmS214t
i2LWm5iMxmEIgJhzpDHRZKNmtOsKQCQMdQ49LTlb7LWWGrwyJH/M3NRuR7++msnx
wx+X35OLwvwdqogSpVUP9DTodVZ+RGeG/ipg16LfemyC+bTdzD8Q4vYoX3STlOEA
oEksf7I5KtOYtrGEXNTZJ9+XiNmYfsRui/4qTyNk2nndESDkpN9VTbvsTQmiZa8f
D/bXR85m6hKzYAYMalKSoHxOUhnmLTvTSp4+K/BSJ+PmEYAI0T5vQWM4nxZs7W+c
XCw7PVT02V2fI/TvmnsGcYd9/DDFVuNjMlBE3x2dKyTupNevvoFYctawh+9ztLV6
PcufaB99fbHuATsTvGl8Lxw4bst/oj/1Hx6bLPAvysQRYCA0F3dwJOiGx1IEtrWd
sUzKrahQTtwxSZqiLkXFy0eDH+iHCBQD81hKYIzMuvxIaiXf3jWKSifu2qdopalX
UmIdOKP5AOARdguCfl/PX1lbytoOmT7Jo51yBjQixk41h8sm2KZZ3Z1ti28Qm9Xs
oNlfNX3wkq6JDWMF4YVHkIWfGmhrQZ0xyT99WgyEQtAXvX1Lv7BzKzUag/zKpasK
zF3/2KtGGxmPRESkN4nkNaB8BbaSFzWvIU5doKoVIllqD7+4u+lWZzvFWAaL2lWe
M+ZNw5NYeLW8yw4uUXAFsRvSRRIowDFkqeQ6MQHEQTMsbqeeA3wa1e5LFicXcv8V
tNan96w+uEPrj3o8fpSt2p/9n/E/cM66c8tx0iovBHtsEwTqfJ61zu5yhIrRkCBM
BgFz2scch+LmPxThoJFKyTD90SnKalBFaqOm4JI2KQgwjiu9/Anf93nGOS/Wk9b4
V+JCk1AIkgXpEmhAtfx+kZnJKkWSYou6EZBjnIKADHhMZKvZ8CbewxfOVIfIaP+c
cJcDFKraImsfWeX0EdVhuabqOtba53JN2t+EKeQJfwd+8RF4nmdm4h0h2+HiI0p2
wtDFcJmcPimd8RLegpjr6x3lm2ZEpn1lZu3eJQdXBWcBtG9PW7t7SPb4VXzBWogQ
z7a89s5fBrfiT1iR9OBJC1oixth/UHDAuQbv6AsiZhDj0POlZnwa3ObYESooj7Zf
v5LYXdEqyEuBs5hnrRXUQXW15VSoVz3nbuPd2c2Ajr2FE3pJaeTggIf/WFVV70f7
734qJ5y+kDNasTRLbhr3geeEaLwsnAh5tuhtfaNvocRRKh4vgbFE1PMQ+VMlVm9P
I7u8FZ0e1bpO5CB0LL5Ne9XGtbo15nA5OAUXTJzJ26JFWS7J37F8ksspwnOHHDVp
//SN/g4UkB8q01CWCMD4MPAbF9Et+vxlsDfA2p0qvsSnj6fMRw375NWX6VFNtagD
zYtBJcspP02jpkG/IhBK+TUGwsZnw/O+QovXwC5c67X1wSXvyKOTd5I+Hphsqw0g
9gcChjmsFScUsrS7vLwJw+W2guRGKHyye2SU7suodH8pFSgPrGNM4ubwVoFmPbEx
qFo/fiAWlvZUfnZekkH7n9dRTWMAMQdwUXud7Kqg2bfTLe3LP2lRpqdTreJ+uMwW
vfZf26pk472nFHZ36OrJC9Q5xnKlxSOnotm9Y/+ItYZGQD0iIConVP4/xrmW5bk3
M7xBOqc5t1IfRz+nvqoGpXMk8WZf/BAmngQHb27geLTdvaYkcz+50/jtfRlfx4kh
ipUnSOZzA/u7Rqe1eHYtuPdzZNRfO7XzPGkoPsk0b2OKhOKBPcnVAk0lDTRBNoa9
UeOqKPs/gTXJvNG+ObkFIw2KHSXt6ZMZuHWmvuLFyqxZJr8YJ3kpnD/aFbPyDCCn
IA15KvRtrDQuaRAogF2X40EoswCml9l2N7E/VySEfOJaz8qvbEer7gxfN9/uInvI
7GzGAMs2CjmngKGVitv2rwnp8/YGzfIbPrYlWrzMrdFkPqBtLGUn4jfHSM4ctjGM
3/hZlcUh3uSH4YMVKf+M6ppUPOfHHtmiEWw/1Zjf3V+luKelrwSEjjY5vOH5J2Fd
deEiHvFTNijF4QLM84DN31u1uAKgFkT0wBrBJzDJY6cNGRRk1oTiP46mA/gxBEKR
CY6k0MAuZrN+NgrenaYiboCg58718KaKwmIThmUrpS0hHyHAgo8YDunsbitBppOO
X4pVyrNpnHEUKFsLg+EUJH0dnvbksdX1nl/OlaWm7PcZrnFVmAkJFZ32ZXdufHpt
2YKfMTALRGim5+NmZXbvGqSPW3WaeFOuFEfJyilKI4qOoSi6gGOh+k7xRMIq4BTe
5jsKofujp42MHvGDd4wtuF0kT+2EK2XMVbJE34VhKTYyv+bA3vnh/m55jLZb20Yu
EOlUvI2dYKgSzBBlCf1GuCJLCt80sOY2+JeiqQVDlFDy74aVxLGfI4SXPUCo3+cV
631KyXGMtV18fvBEa8cL9z8Wrz9ZnQLUoRUxwRMDj5ZQRnRwxmn5SO9WXZPTjVw3
mocGU7+amQ34bNmNz/NbOHvEM3cRw1rzHvuGbehZvtvha5jCvk5LJT8p4EcDeliQ
VpKqsBVQ12tUvvjAEXDhexoo/avc6p8NJ81g61UQCU6h7KNYB+zpxwCx0ihrUFCr
lqvkzvv5Wt1hngg89P7mZhZSq2WLd33kRON+f9vHEKlMKbDSMY4ldlm8rqhQTjf5
bfoOD5nUGsEy0hy7tCsCcOmTLRqdpE+CsThBgKdoTnu8SSiEXOArtV7c1YkGRPa1
Ut1PVMO3zh58QIG0ajRmsFIlmZKCuW0aBXzvB4mVCgC/ZLeqILyNlHR7NfrUSQHK
cMoq4ZzMGi9sFI/jGDXd5lYJY2WItxXD2+j7pdZeT42eDspbb2FAuZWjdBHypIsT
4aYLujKEyiAhlKY0GnJu/s7loK68yFyZTuIqmnshTGd392X8K4KS1H0hke4jk800
V3tis9V5DLOpBrfEkQuztbx6AAprJXPClh8e7dD86YWPGFaGvsbvXN9X9xP6Keah
WxCoM7wGuUXJDiSjxB1DJR5jwYxbHMfcTNA0bERWU1jC+n//be2v5CBApa4O0VzM
PVGP5yxhrLXYuUcjr/BtdJd5bwh55Wf+R4wKRjxRUHEEDqr9JVs2w0tMzBlzsImZ
YAUdaKzQAjqnC9cf4ZUU4tFmTkjYiAw04QJRRSw+LbQY7ewYADHb2FwtcktWwbyj
EER/ZnWdo7NdfW5rvCde/fKCipHpftrBlrG3bpGU2z1HDQoYGwvYO/Jl9ukwfY38
nUFlylv/42HgKUY+msNkOpzaGZX/2JrIQoefHnyqWOryLKlB19azeXbZZs9v4Bac
icEDCCYwx5rBx28pwAhQHxrQgnxFWCl9dpxy/glIQzj++tvywkF8iQmmg1gHnBhD
sTmNu78qUrAp7KwvWfAo8xWFxmJxw2DYOHAUmZAgWKwWWxIiOgKE2XnN8sNiI7q5
0MGGC+35KY2xF7k0F2UlL2RPWlcCSFH/+Cl20h4Pq7+9mD3vdMLcJT4Q3kimpqtr
i0KLOHY8tJJZ1ga74bW6yygyKQ0BTLPpy9CrmjZtHdfZQrDEdvWGL+kKNzqLy4Th
PuNCvSkM5YhX5SvZQR83OEEFPtlV7PeU4RI/6KregyErXi30WEs4njY6PYiltB9Q
suMUIXUDgcDh9JF6iV9CyWxAe0QF7MnKEMP0ZSbXGim7BQWIKr4IMxb7qJvfre5e
T7z+KoorruFm43gG5JTuXzzYy8pMLsdGrUOHn+ozrtV77xKNLr8KzpT8DLfkdzbe
RsLLVatVNpr85HFxzAyREO71i1ppC9y9sonBRVxGn9UklODeP5PxPdrUx8QKOYJ3
za/4NFdiLXD59KSRZnYzPmdoxyUmerFTd9eQKCeRqs3PQTzToG5ix+IKPcIXERL+
CuETulfS4mmrZYzU/8XhMKqRlb4WqPrpx4l8SYf7UMP/18aFXi483HVsKzbCmagv
4nd/XuP8lHO04fkQ371IGne40x5X8sr/FWLsvjmdemHDLKk4dsK2hmbZTebMzB9E
YtCiu4eKEqzPTWDi8xhBAXmqGgDdLdbYqCld/UMJYptGNji/Fj3yd8rxaizmxKHN
7iiWn3bx4IFLL1oKyYzV0nZ/f/FTo6ncr3lRzdteOHWwdtBtdWdhuhXuAGK0GR7i
iKb3961ZZRRG5JhBXDM+Kbkbiv3oZpb7rjKmN7OCGd04QVui3bdYtSFFRyyge+FF
yatVk5amizO06Yk8i4gbrubMcaUYrvogqm5z/Qivtt/vlbx8NRwTEltUsjrkLZiS
s0JO04M89teuTz6L6aWmZNcUrD1aE6ruzqC49PIGarfVW8rquCLQD9rsMU3f3Y2+
zviEY4wv/PeWGyz/28y5EcumiVFAng7su8EhqFiODMtCVBMbocIcmuDjuaLqtr/0
wNAOUllTcyLo5wPhaqZzbxNR6El2CNmxyzCAr8TNY/JLRA7WSJ+QNhRW+I9ZWvPq
ElC/MsSkUQcIP2fcUA0dp/6zrt11OQwFT4WbAJGKvKTzTxmCQErzKfiUwi+Xao62
0yR0CHfb2l27mt+Ef+vnwju7D9wqDVJhR9iMb3QX86/Uot+o6dAEg9Iy+aA3desZ
KxV4bccAh1fFO3ka3IYkrOJNhDv8QoFjwyDGCNxFr834z2LK/PDAyL8bAskaqsSQ
4McRmAeUy5H4FhZeWUfiV6q+DVPAn/kWNCUv/uZuXAWL70OFQLNFkXV+qpcoRp/6
Q7fGxu1DkO3b9CYYiNwpxtgneQjPJk0Z/zaGORy/cLHgblIk2Z0AWUfBa78FLLBk
NkjWiYEd4mlJc3663If97BESibKR1ssErme1NziGBC26Cm9t9yAzo/wyi3KHnTSY
8aMk0RyGbcxVIw0mD4M6J6PaVt+7O4JnKjk0VhzMcBJmGSVnho8bzGZVH8TGTFz5
6cLHU8gdaXBiKgZAPO96g0EBI0dZG1p00c0jIElqtl+P+uvU5yX5skeJ8LJPprSY
EzXX8fd2djnWoDTSbRokgCQkj1D8cteOZWyk0LcY2AIwA8PDOX2Wi2ZNDU671w8B
GZrUcdbtHUYpZCvOhIErzDYCC49socUkl1dzLDpSleR4KgQ1EjwR6ibJZEEXZ+R6
9sPz1q3Hz7/VYmb1tw2twA4MjO8tJLL4Tc7fjox3PEBkLgeXoH2y6XjFL8iGs8Vg
LHFM6RqWosE0lYH+BoFc6hccVoQLthUjOfyWqRPqyvNDBrMMg8lIHzN+t1mWKCms
1Jr/1Ki9CmTeRQe8kPtMAWXBiP6doyBaXXhaqKmgMwl+xiKZC9uMGD402whRNkdz
4xmQ3iHx39nN1yJ6WfQtCK3ungISCYG6mIcpeU0Y9b8Sxy+uqc5TpHhi4MT1QzVM
z8kjfddQzYtr+gghuZs3X4S4cnujV/goRT81zw45fdFpHLu1Kfci0RGaVLi41jqn
O+J5FB/OyKd7wp6JHphqFF9RX6P8m7WHaOg6d3vi7jTTap8kHhoxUuqM2FFddnyH
+yEUO8+RtPiKhZaewZIR8blslHNtdEytKyzpQvQhlwQBS9erPMMmqJMof7XRUuK5
dRQLpnSahP5AM9iGDgHyqrIA+CWrKg82VxWtcF3RzUOUFtL/6r8Fiqd7yUkj+8qk
wfJDjnFHt4Gf4UQzGbSkvqwI0AkAKd7Gr6kvItNDlrj2lS33zDrRJ3cwvqhoWPgA
p9eDQiyZJEP2KqWIh1VATCUxp1DMBz9tM8AWOUQAA0CRqEbF9XXSGz/QUEgiTsrz
RYDjKgbGy3pV2uD8DLyuSTUMoOvTwwng7rLMigucmukA3A+7GHdfwL+Iuzw7Yfye
eCu9QjFZ50bWNDTfl9JC5IWzPv+zpnLhYpvkS8rKzLMZWWTLX4QUTA3jplDeWt+a
pxmXUzuKzO5tizeUS6DfuH3k+X43By2qp9Wed1tWXYOXZr2U1BT5QAiGTnFLv0qD
KbpERTRgLyNbNHBfrLSxdgHbaplmhMr+cnVVituVb6FjZObDFqECVRV0iQ7tdVGH
toG4By2+kiNq4R5KpVVgSDimCrRBrUWHk1F+fXSBRhT/ZVMOgSR8xGRbmkGWkz2m
kWKXKYHFanB60ZEY364qEXOmU7qU04Pa2QzCXN1KEFPiBua0Wic06YAeqHz84FO+
HVdVjONMffnB1Of5PeT+9PbnZoWs1SqNIP6pl+mjR8VVKftF3CuZaehXFyHYqdCM
aqqFUX/IyoM+DqROiskC/FpQ8yBN40H8JdiMEHwUNByyPneAXvyVBx5xlrLwDr+8
2rLDUPS9oFjLIABZTeVRAzaFIrMALpQivlITNgacPM0KNFMw4M0Nn/De3D+bdm/W
RDHR1YR8owKXrZzCVZw66Er3uCsOyjtBpyRBXEzoKFrJINPKljzzuTdIHf+BROwP
M39Pox3Z4gjpsdTcE1R9V4P21c+zo5bs6CR7sXS0SkHH9jKDaO7/0/NnoNLu0kuK
78NJN2k5cQBvxSWc6W/kmPKzh7rZP49nepJFSkh+QZFhX7y/k3koRUgWKX6TNWLx
XLiB9U2Z86FNi6HxTCvxdj1Nxwdx+Sf1wk0f8LwkvSfNFA4MQtIX3EZpDWTOIwbq
y10TrMmRzpazsM0EtKjplBGjHH1K2q2XKpFFdE+VcwuEKrXVrgMiW+YeNFHvGB8D
sW0b3AsBLPDgTqYAwvPkU7KEatyNq9JT8H/3i+JcZIH9RY9ax9OvlLQCZJ5mP6t/
z5M/8EFgc7W76q10WsRQwMWLNFeDZ50EeppH1pJiLOrIGobxgvTo2KZEoucPHY4D
btnm6U89YNta5jxqWXMYU6F+ZAo35aMEfh+p5v33wcyWWZij86C35ihdTcZ5e9Tn
MIg8QuWIl1FMlKsoX5Njz4r/D02PTxbhzIJSAV/gf91dY0PycVnbAmbEImp5aBdm
kVaFmcnNWa5tM2JD1wqvX9ZbUgNwN4SrxfvwuolIh7qFvhTY8s5Uk0JDcd1+5sy1
GtA+TdgcGH0fjJdiPJxJfy0Bhr3+OuH0cYQdAJGms+5vgsbRMGMv4bTQYW20YI44
d7+4vi0ZAf9xAieJm2BMfx1mzcAw/J6Z/xLIqaVNpVlGSleTwCtlAyMmEfM8T4on
/Kwuwhz1icgNoCSuh29M3l6EdzV4TVqJAGWYS8jdwIzLWHY+SkUA+/NiOcmAltZm
yLjo6+/XMdb41ZwhOsiNhBaNoE9GtkBtfzglTWepRpLasu+bMSQNn6E5XOJhFVGG
JQun3wvp1/bbQFe3JukQZGbUR9fxR5npuZLkbW/C6jFdgeefaV7DD9ZgTqGsBglG
VF9UtKQ3ztsIK/jvUkPxK7PgX5R/vV1FsH9K45uICvjgbfO2igkxVbviFFoB+Ybp
EVT6U2hbEA7EFmVssO6h5rgUqvD+gE7iwsHvs4OTwpfX7+jngHNAchP2kbTxIGOV
jNxQHJCGqmUIdcxpGnwJ0N2CcgGKwlBFP1B/YiOMinC3b9PZrAF4i3UUoDBXr1OX
jJx9nfJehkFZiYfzBI9dneflh+k24+ceKV5ZDKQuhOmOm3fBstqMBVNit34v28yf
cUljFCibaB9ngvwPQnvVRiwsoCYHkNYPXjcPalTzfteS7SXZcJySVoU17cZANG0q
3zz1zd7GbSjHSw/76dkb5zVBcmoohRFIElTCfQPL9TslIbMg7vmGhpjZ7RtYeOue
G31Q9SEtb0whAQWAAPm63SKKwt0D+h1hUZTMTyevEtu4HSIldnyoJV2lZRmb1eB+
K8gRPVo4IoiattBoRDvUsdto/h8aal0QjByToH8jChCHTVVbeaALrgDJSIr6NpUM
T5V2G4SEtO89kgb2g4wg4Y6djZIcn8CD/zqAn5iWylJSAM0xBJihbuDgvHqbPDL7
Ec4PfGaCsbEJ5cpSfhZGnGt0nX/1XbtMzfIifgywMHoT0yoa58PlM8aHywWuUFJS
noLgFXhk8kphEMSkWpwjspYGEP/UFdAbscUCaMWLOz0ur77DsTy6ucYf95ojqdyL
K0mv/KUoL6k65jq/dkiW6zh45bALl36HCra2SEvKl+/d4Rewz+Db1xRKvIn6Fml0
/7lsmTG8EZXTGduCyBE84spDyAYz4CZgIeXo2uhqyh95QTBAG+OzgULDyhluFQZ5
/uIPbl/XBdgri6eR7Dg3xGrme5Cz/EFFDrf0YCaV1xKtrZcnR74ce8JsnmjdDyou
kwYps54M5A1ui8lgBntPw606QUXeE2QXn7rb2JZXTsWUVBOqh8JUggRn8lxfZH5e
R+1B0mOpC8cJD9ZY5GQ3ef+35qhbsciqT2B+SJT3+xhuyIgArlV8Jje0397TTCMO
jMHMVBf4AHq16emv8tp4vNzOcdOhdUurAKcPeZK7S/Eh02ceYEzQu6zPocnvMAos
uia/Mfznc20JSFxeOepG3DKTOuZscB1NqmmxMvUTKKKrg4N83Ktopaz/NJamtt6J
9d7aGPDfZfIuONz06cJrJfm4R6j1a85lhMlKdtSDHhg7PSXRjb3jY5JyJxM8yBv+
eS2S2TqCti2euBnhM0lxdeZmbEuwnOyi3BdMC/tvKrXHAIEkMNSU8m+Z+SjqSoOh
KNSIlyjnKAaOCANRigg1rzZHaM+RRGvqLWmEHAYDbdnEjuXZz4LByzqsaeXfGtIw
V8cRi1RH+fvwjwBHuZB29/Hw8PpFqGmwA1Y3ulnhdQoaolrO22bqYhqmnqXrKD2P
ziMlb8CgFi6Sgl0ISuJVh5er8yWAkoRT8YulMcRbkDF81ir37Y7g5kCv3w4VW7ZP
XRXeNeC5tmxabjU69By+eBrzCXociqoJl+lgBtwsIqnhZBbd96l+PMj7ELrEA62o
nXu+MPXIKiqI55u+/L/bHovk4h+s4+Z0jHARrPw/+LDaVHuVj0+LJzLfhrQ6JEhz
iCXD/yPXyhXGXU1SoxR9HdMsEtrSQ5m8ubdIO6NpdhHYbJEFwZAwIEvTZiHrPvqn
SUTBYO3J0vTqaFQpOXO40K4WHJ66aseQn9qcIlO0MS1YnJwoVKfzLEEhQwTXXY3D
J4kJMFIaOdy1ymXcUtPkj382xc3L0A5gbYsdEWE9GX/9PZ9DbM10a+M3/KyJkmYb
wdm91ZKOASgOFPwcqzRhF9AgZJkVhq5GQudIRIMAzZZF8S2+3TYnHsEz5sudmgFH
v3KYEhZHdaGv0xMD/lrsohmt/HkKzRNActtKpiAxncmiUTXJdVDIk7JrHmVtO5vX
GTA+9nvmPumtarjz8jkbmQ02xJoz6VcK+z7oYfQQPrw38XVh+Sda6uQJsveOpGYg
KZ57sWABODwulxjJI+/BD/OF1+8fyegHlPUhnzeWIjEAyTa4QDF6fqDrYxWCjEJQ
nHv105aPDj+/PQXEoNebddnAXBklr0KgrV5YVnkJ58RWe1qkvKYU658039PDv1tO
NagzwoZf8R6NhxWePJPxhvGqMnUe4gk63iCS3qhKDSYz14k0UrEau1H4EZf0mX8u
gM3Nj2jo771eIYPdjsmCkeYtxG27aXIGYSy9EERyVhWyt6BT+/3ufFHU2sftxxMa
0BQjgodiyE+4oWZDEy3jZcMoP2qhObfOkfl2j7Wz0G4ECpixNO4biBDpzEW1My6V
TSs5vd5SBcEpF6ynUGmmu+HXOX2EiMmznTMj4z0+YrDYCiarp+AoUl69pnsayYuy
Mrqe9BV5Df9vyfxtO99Nezwfmd1V/mSgtnqht/7qc78VAODq2dUFK3kDUVIshARk
TljZQHYMOPrHXX0KYQ/OkDF+0+4fu44T/PNe3hiJprvd4mz7faqJV37zZZ82ieET
ex4IFnjkHEZZFS02gj9f5oFAKzIBvkubWyQa7hhxsaS24LReWdW/T9ZPImhSXP0o
9ETZbkRKChqI5SlLW8few3Or04je44z5VbggVdvov+DNcAsW1TOjU6k7VlWwJXKh
ofb2KYn2qHpaNkgIfw/viA/2AscclTqfx4zHrztyeCbqYbomjHYqmBS0EzBpgN65
hsV9mnY3stE8Au9omzBvGy9PJP9mVUYP/rmgLHSCnno5VgXhkLvht5uKp07Pz0f+
Qk+FKqMRrh8/TP1P0x5zTXkyxoUnM2q8P3W5lKY0T21GeN+nWB3rYjlHV04vIOFc
VuZZsHlZbL3iNMPOdRhKb9DgqP4I7rTO2/EeIqq3i7MEu6fHfWfzsQUiJVII1e6h
Jw8lAsWqyNohIYdCJOHddPGrjKOIWLDnlq5Tbw7Y+L4E7nDznhY/7yYmhTNGenAY
MFssUlkvu+xu9S6m56Ls9SfBmLq0aPQlxMVfIJqLP9eVZ9sriu0p/ZNHXvUiD/nS
/9RNipW9DPQtCh7OStYbk8iwALPZB9+teYQh1RkjE2jaPHGv5ewoA8mq0FqkowNA
78xkuVRpnBTh0Y0Hl7tBlekhElbRf5GHPGnGAo5fXpDxW67BF0GPvgbM2Aw1W5PJ
j9IAFMGAIpNiSbEfvP+u/aTl4m8MQZC6fHDkiRAmajr5f7wLtt9SXBeaGflA8CJc
j6Xrml0QR6EqxGnWBccsjTJ1Oo/ljU4ifXef5HFbzFbMSbutMYi3l4GX5s5FuwK3
fED5OaRRBUsEcD4yBHhvZGBu3zvPTYz/ImMxJrvc9heSzYXMC7sE+/DekmTzOM42
WE+kZqpMrcVNJsSKjxHPVg1kLQmRxdDXwTLvAocZ33Aedlej4hKHrdYkl4rbYHtT
R+yUqzDObM7V1IXtVzdQDxqlIuBsMJnNRtD8WsKnYjvlYBhekP0Oc/FdQEvEJtvd
rr78tXrQV6SjvUjQl1w9ZePmQiLgzpPuSflo6jswsA6zpBi9RI1cXQa2fNebwxhA
NhP2mQoCK3VC72MSVYf/2/sHh/XYB1fGRDwdtlFOgA3+unCoAODwRl3RorxZ56Yn
eC2Ludrp1qDv5+lK5okFtASVfJzcZNOD4chuer8VuMk2MJaoH8uNVPQsuEbVpXY8
Lk3ngLADllN77N3Zsl8pdR0zNzC0g1lFXY2Z1egfVCwaIoojTs79g2XTlhal4C1Q
TvC5FY3/6IJZxVjQF0x/UKoN/zW9qsvPggAjVBLPq/gtpT8ooHYt7MaHnPVJhhQX
v7k4P0qLamSq6oovtOrbJ+mFYg19/3VbsHYJVfb9lOa5H8EygUzNi8/RT511kBUs
6sYdqqw7CIZ75vlgCOWaT68sqxFQJMFlLKfe/4YwO4kZLiafPEV9VUjdeMQrbAVF
iF38jK+zhy2d+wkGztpuSfrmsUnLPCaScWa009mE1vakdHlCcWMgkGFBvSwvq/5F
Rk4FTrBAwoUbAW8oNSFSpxGyyTM2GUW+YLI3K0oTA8iIYva293GBTNYL/8G/NxXE
/JWeJwE7QLzaNvjOi1Gd9vdqfYyF8zrIU86hk+KR471MbDGyokfFP2EAb6HcyCTI
k+VAvF05I93iVMySogeslrUFlmK6a61fjLlcpqWnVHKNc/bnAviQRyvI8O/m8oA4
Oqf5kKSsYCRX3EusCbbEkmnlgv8PMZEy23/1X3+EaYpcOhQrUJ8Igz0unmlHmlw/
S0CqtQd41963bW683lnXMOvgjdeXA4/xn/4Z2WhrPuj5RWoGsFuqdynPMeXDsICW
DME8FpyCTbRxaDf5CWbBcH/pZggabhL5q6s6eLLVbN4v2hP9OZ2RO1HpxE1px3IY
8zg1bhtQqVTEHiZYQuL/iLdyeENtE0gG0Zfr11GvrUlsp8iqnwWenBe/5iR1xh8q
Hd1Y/0XfY1xIT3YAZ/ouhmpUCbbxw82IeD4CSTYwAgbks/t0wVlAHRjeZrkLdXjv
8CFQ+yTPBMZPdXoSRRr985KvS9w31hSpMZc5duvhK42XD9FELvaykbUmyr1Pg0AG
0NPnaudK5hy/wWh/6Jv7z30WGKbx9CmsQfVeWwjwChm+TaofWKFFdSPG9OFMRoc+
cCKxk2Zrd3wqWHCbJDH+lktjGQtcqJDF1CdEP9J5Flyjwbsp3rRqSgCvwmqqAq/g
Is5fsvw6xnc1GTcg0+O0GUaUy41fEQFo/UMcJuD3zw1zjUNnaxCXSAIv8pXqoM7O
z+MPybuIi6bVfL4Yp/IOujgqKGUho75ntGZVPbsekZtL1xk8D0yAz0KUU6rkPz4W
R9tG6pVh0VdtQMNxJCvx73NRI13fxSrbFU9pS959JKgXU5/zooqi27LXMy2DRCSb
0www+Aztp4Y+kHaQqm97+fgrlfLyGkwCEHAd69bvCpq/qiuCuCkS2JbV5fktCD6k
61s2lI8aEUDcSGoP8nfR15zLanyytF6SDAXsq656A8svebHKWDVXZd9TQ5H2nfxa
93DGIcGYCihG1BPWrB2K78+6QQHUUL7Zp7rVUz2vzBOq3yXCmXhFcqOLn6528Ibq
Gr0GgJb4w762xua7X98Zi80Qw06r/fRFAetmFAWBh9EBqXW+lvFfBTDLe5LkHvE3
bYMFCjwHm9P5iozKZ3yO7dTIi2kErIiocNHhYZ1a0yta505UemZcr/I6IP4Ik7BB
UPIG9cKtnfHo8zIktQe1JxUXD+0ThG6HctQDO57eqxu6+EJ0UMon5Krgtg1I0hhd
6eO3VkxLdPnbmsfOuSRituvRyl+UOnxIDEywYY0CN52c9K3ZT5Rm9f8LJ+TROTI/
VsPDthldnfLKhMfBPrZKV3HLFpBC4qMDfYQpeeWnkApuyIr17Or6aDUaVcut4Jl1
Pq5u7A3PMrzWWhCDTLVQP93ShR9N9HBeTcVN5lNkcEXpWL0mwaJODLcgZcZVq+Oa
RcXfZ7dlVujlH8+nj0xK9Em/dLHnwhxtrUR+LgD5wsCsU4effEL3tH44waVMzqpG
KcL+v2OwLU/bZlPVcTZ2U9NLmB6WuNoH7DL2EDH6WnqeeWHKY4W3f5ZPPDtGA0Uo
9SECJTSX+3xJq5enYgpdcREl9IHsuYop7j5yHcoHuBsTb9VSepfo3lajIj4qbZcJ
i9ZZ6lqTfTonlePMgPYEv9JQDDk3dJVmpmMqvw2B2fC2UdkcCIxeY7qcOXQ8lRRT
CZy6t8051y4nynVOYj+AEN9y6q+Dz/QcPynhWBfWX0MJgCuln7klTtBOpic7Cocz
fQBoPriq55PPXqLcb+l3L2ojlEh7C8Yzbxrv5v7YS7PUU9H2fbFLK2dadMXASgWx
SwTPctcQxepTVWuw5dgBBC9poSJQ05ayc3PV0DNrV4ZyXbZv4Y7k3WzQ1uSHtpin
nqMqluuycNMhPrPakLVoqDM2bkUv9zLDheT7ld/pdNuLzAlzT+yQD3U+M970FCDb
pb6DlLzLHfqTp+6IZCK3gW5tSekQxqv1aTOsDSv32T7HlWUghTEUE8c51RabxVOo
U4L9Z3VzoIEdCa4hhggGwsrxfCF+IJsC2I+2YKQvs5py+OH4KHy6PHSvUU9Gu4FD
8vOhxRDVnO4YnP4VVROn5lU3+EotNQNid1f6CVI+CrpIli/l5jZEZsoNkl7YvblV
Hhh70cdNpLASP513gaDtH3hB0Q9C9VY+jqlC7SBFCqCpXMD4NZAEUoQJ4oMZJTAS
5jiaQvNPu+ji+v0HjKzmEoEClzIHWXHR2VU772tNtLS3zYmc/SBqHx5snlfSfXD3
iGZ/mZ2EfRLovSVLUgARTvRCMrzrb3NDOkFnYztniMcO3ojwmFIOguMQaILgM8AY
ZMzKmKYbqoPIgoX0CZ93eJR/FM20v4fk/vo3nVb0fQmzGQ+IWMbfWN39Bi81+0bw
QspUh04cSTqDkXmtQ0Vduajbhphx31JEiJHnPkEPIJyBNarYtuxqwL5JaBpAO74k
tK3QpoYCWvFnK98rIN2rEDEG7LgA2oEgFmv6vFjeS7cNy6yKzvWJsrlQStTVwM7O
F6YuqV89AvV+HPWC9dn34kNE3bJVvx4HZBImvbkqVQXupglyzdvnpxuK9o7F8hdB
0hkJ8+CP1ynKbiPBtHmT9+PddnLetcirvWlkE6mqOd80RPIeqaRjtnjYaD5AGulV
sf1/x3A/r8cI+dheatycnAd/Lj6XueuI5zhrSiH4uPlMV3LI3aytUyRRKtAIUHyk
AhMzmF4eMQGIS8ZQyTIdD0i7jorzIXcKGx3coTzN71t1C0NNGz+BjVXkKPS2N2AA
Z5RyGi+MeoZx1dI4QE1221Cu8aaML7CTp6/cRRSq2KpjcNu8ZnK5BbLqCD96c4hp
RwmO880GG1O3+AqwaiykmhJzbIB6+nTxfeIFgAzBp9bjP8vCk/lB0OV7UlsZQ4xZ
yQnjkti2894Z5lHIPMYn69KDloRI38km9BsG8wPmPac/Q+9Q9/AwMJ82CVaBnOsO
ydfrLrgDrNCQ9pTdJ/Jb595Jk/drVJxaoI1gPWF5nkZlndPKJqtvYcMwwEUkjXC4
4rJ2yMnSUIBoUQYbvLTp0EJQCm+y8un5R5CEiZQuSIhclZFM7rJX7JRatrzeLrDp
c7+Afy0izwyq66sdtPUozZKZ0ngW5Th3lFw+NZmgUzyB/JF8rdAN/Z1PgzLGCani
Nu+DvL+YetgTZxVwU2t8RWqbHn2IPO17HjjxQr0Pgw34hVbX/yzt6JbkJU7/PMvC
zoZawQGTJaMDNQOu4slBMiknbx/enbF77UgExXMyJYt9eum5wBAiSh/gJzkrVJhc
VbRbaoCedJrsP7y5cpIJsTqV3QdAM4qXMxfW9r3znZt97xSm7Grul+ouBJWmgP5L
849Oe56E2XXmhQSUS/GiFqmSHgLhb/SQznZMQl9wrpdW6flOc48lw6sxw2blh+sb
zJiQtSGwbp+ybaojCiZ2fpgBWRJhm02PhVepWSMWSE9zPu/ygeVUJRiOfcP8Izar
IwDw6Ozq9iVQvZv6ggbS+DllGIRUl01wClQui8QQ4YoKQVPnufpvSoqjeTft+boG
zuXKS8hFdaH/wKT0y9il7YtD+loR2NvM6BFDvkpQbiZ1Ky54GKFFcMZr9TVcQDJQ
CtKfaivANiMi2ewOGe2rnHAsgeZeX0xfUgozYMQ4o3TnYFmC/tAgYoFhGrLMZM3x
Pcyb6pS4lmL4oEFQVOau0/TSxX1WUyRV6o//uS/KFYx9OHOGIGfYaKR7+64vzOI3
BCicUelUwr35JRoWdGgfyPSjHNu8CzQiYQWnNxPSg+TFCujXaa4l5VWojSkCREVG
D/kNmSJI0EHnSD0ZUloJaDdmmJLws2c4RC53eMNRDb1s+UgWZLaV0pLd640l/ayA
6LcsdYBm2Q3IGfvrC4JS7oF0GycLbSwXCLeXkKq6EPkOfxkuMc1VBLeY8lpUYNu+
N7qa9GHxoR70dq2/tX/r6jOZugX52u1Hipj7Z+IOH0DWYYRf4qASHWlKEuTCzlNN
IL2F7Cm7foJYt2Pv3YJ4pBWqGTJxdnkPXYPLGlinMYjkVHvTT5BEz3ADIobxUnqA
pcjfi4y3QbXmKi+UFd5cwR1RTSwmblccmDJ7+cY0bdfhe9o5K3vISVIHWzd+htGv
0doK+BhWCQmp7ZtdOaXDhjmUzFJm/ol6utalLvhdEwTIiC6FFjMeEyZdASxd9RzN
gB6UkIPyb5n+GgLUxjtGcfk6u/Mul5/gygMosxK6jzdEtgkpzhqVGi6DBGVjDRsl
hJENBNJbrS/cd2IVlHX7GnZAF3KUSkKD/JxGVJUA+BvybAfv7LjTecJgu34RieZh
km5w3oEnHkn2ofEhuh+ghz30kC5AcHg3wW5aL03tcc6kxCTzBEyt1iQBNsFmoMXk
Lk8f2wWr6YvouLwvy3PGZALz/NJqm4kf00BAJfEK3MKwYsBkQwNohJeOUo7q/Z9s
eDnyHz8LlRokk5aNngKI2FfwSNwrevMCIJEsAgW1NNC2WQHgSmFXZppCg29wlhwR
21hDmosvuZPAG9y7qCgkbqAQQxE7WU1UWBAM4PLK30axC/itJjDj3HKCKMRZUtL5
0IyyafewwiSqjMfLUfkOVRKOugzkvG/nbzaAOWAc/q6LE1EcDXz1/AkUK3RT+hw7
8hw4ubFi7DU/PfUlgw0/iGuUvNzYqlvz7s6k/XCht+fF+KT/K+h7MjnhfymCS4e3
0d8L4qMl7cvt3x2RsqBEOF7J87RyGMLSLxlkaNQzdKDeAdWZ+hoIa582eAD/rxzf
98/+hY3M5cAyVzSn/QQFHfkswB3xAEgJVuSCfYt62GOB5Iak8mArD2KsfcTXh3ie
8BNiPCRQ9W993EjgoX17Ci6lSNKhospooGG45/w0exHUbNRkdojkYW94MezEPSSe
6sPWWhQZrIPLJ3BsmzxNRi3MF2ICK7uZkW3FS5q6DA4xHapktXzebt7mgZonhTJo
jUmD0J47Y9ODvh9lHRhZEUOfExYD9zX59Z2rDrQ+zOW/rvW+LwEEMa0TkvM4xJT3
6OFeoacGJaP2VzgNWo7BmIZl/UFqyUVd03ITcD5zSLQ43KWPWRi1KRw61MxSFnsY
ow/xeqw+PjARloGJ5HrJ65GM/WbJ5/TcobO+zfpjvKNCRn4kmuL7S/YndLg++DRS
ziMlZo73s8CmZ5vQSynikCvINt/1vmoyq5g/p0tzo8xytKWTeQXV5uMb9QNGQJBX
MznZNbb5AnSV2/Qp5tYP3VSmHaF4pRpqUKHkO95ODiSNDzuFJJHyq3rVNuDqQ0G9
c96KvXsrqAT+zheyqXt8VbDdS7ndS3JsBde+jrCzAT+8gAU1HJEykXqUM7MhM0Ss
/LyUgq2JkJesopgNeVHKKGVtcTniuBl1eEjnBx0vy8HgNHBRPfRNOzjIxWRpdT0d
tF8xZW+zuyD2RmuptS3FCM/3n0sHjkBUcHJ0j8NvOmzrXs5DcitlRHX/jAq3CR6N
n5RNvBdnT5L5ng72bWFwhCbSNCPzVCQJslaBgQttcVINXR9yhJXHmZvuf7A04cm9
3pOGvfOZuSSMLij6mJ+1RMbpaIw6ZY0sEL6mTj60l3EZO5yi641D5IhHWs9WZgX/
q0Uf2pQuFI/LJ0TVxGTc6Py05ZV8jlt/oXu/C3wbnjTxbRHqYXBy64H9gb6u7vi7
CsQdJKm/8ofaNom7BAVpbTUw+TtVhSZJ5q1Ix1DkGydPafWXr9Ywkvasu4YlYh6H
tD0rnc9UGb17ct3Q7Qa8I1ez21HL4+Q8bnMDLB1abdyCbqg8pSXfev5VJby5/dGc
PVx9jLQMgnyT9Jf6XHuMZaFHQyCIrWHdwPwwawpNA73NNu4eQfgXvyC1ceFHmDQe
mVvDXLCVpHhiwKBq2DDrFOjLfNQDbL8BYN8ezczeABQXtVsPePoM4udVRGnow4SF
bym3AZi0r1bSRS71/Pkeoh7loWhyW9pAjNlDb/gZW+TfhR4gb/Zx36MafH9HOl8f
gMiTv4YtnQY+leFOLuSYz+5wgRcXzC8TrVPE0OaY6S2lsV4CxvaHePIkxatQtk/A
7lDDTzZgeHwpb49Rx2qMP3tB+DseSK2TvMfEM+XFTf+8E+QtL5uW6yTCmn3MbYej
bntTUTJ9BbnD83mMcg0JfoKpn9sERjMNKNndlXgDj5dDiONRX/pDtUVm6w2uVNCe
mcwmsxWwKIcuaLRIriRmqVkLMyFjDzzgdhUcUEWjM4zETb1olC0VnFLddUfLdTcR
+L2ic4xYCAE795SwKOIeqfpQkBaZHunbDFJbmxyPCj6w0yVeEO9n87mrheD2kGQQ
parWZhEGU7huVXqfRQAFDx2/VmL311Wq+eyhwGdR/pygpxamC3mzf4XT+L+QpodI
VFAVvPpiuvAyGHOtWJCBh4+SQSjNYeLac/HMnN8liMHapJB85UwuU2yJS9iWgiKF
tuZqbVvL3BuZjyIuEsqnYkDZue993WJtcjwoOUCC1YUsjlV8sdbMkpv3xQdSDuBB
RkVI0AnOtpzZoI1htMhlvreKXZ2qBJ9h/V/oivk4btGs0U+gfbVo1mIh0iNZ98H+
3o6vCS7nJeb+RXNREZhoxG4ncCR96cHAUT2xmPyBQ4bii/6AAI198HFaJ+F0HgEp
nrEf52pxXIfAYVfK+d318JEgId57lpGa4cNPv2JOT44gAn6jestZ4pzEY6KJl4Zc
/VO0tDChedrOqAJoJKo43a1Y1OUdF6xpH4+LeGO+IrNmCln55VKIKMnhzWlhqWRd
JvG99jVHLlm3Hr6QLbwRrml7aYdY0RIJttKJDCK5N9TzGmyYlg5PIw8CdWZqs/ir
xw5aRA29MPtBeIC0a8JPaPQsLGdHysieDke2GFKRAHIFsecuoNvCZ/mW8elbgWm8
XPTSxveNRIKZfOa1nzmhUYpCXp3v3NCz5oalQgVA6LF3brUD65tKMk6doGUy0WYM
9jRFSiefzG0tI6bxPiXnQpYGqyHih//4jbPhLutP+1Db/bLXiBZSKwsJOImkGhaw
E4egkB5REK4IhI2IeN9FfOKn945I9siTTWSNfyQMvVOlLXduqueV5ic+N2OSscE2
Le6Fx2/x6aWkoa4RA/9I8G3LEbeDPZhl0eeDXshQUc8ChkjYjcL2XyabTFg8kILB
WTWscfMeXvstwBI7rC71GKpeFz9NVj5YNdQHosxl+GALIEOMgKjiFnAuXT+vokq2
HIx8d1R379WmCBotaXMLfsDUHUNa84d+Zpc8eolYEQMaRU+FZ9E45qW9Za94uDgA
JUcyLf8tuTOf69H/+juA/1TCPtJVrRJnAi4yUqJviF1BrdYlBECbiA3Zu+g3XOJ6
jJQ5D1OECinJ+JsL1mMa5G09tSCvf8SEt+6gObCdru1bwbwS9W2CWBg00FciRCyR
Dw0IzQDWFSHKuk1iPcYDomEMfuecdxXlaEF5JLsjTt8F52sxU684GE/6slcfcQ50
JjzpyRjy4RE6QTXMG1M0wvDm19hLTJSdfF+wHm6DQbnWWdliMKDXkjN71MEGoz6C
5OD6rJfhkusbIgpJOfSpSqUSP5tMdLwiyfrNn1y6RMIa9gpn2ucJQHGA7bj3EpNS
pKX4Zc5USqx/ZzaVGzAp14n3P6PQ01GkkXyfFW8PeJlqdDkzbh1J3b+3wwnSr14P
5wBkA2jmyoCRNtj7jUk7MWaiMhEyyegB8ow/DsJxGFeujv65JDwYHW5RFI+Oh8r+
lxpsmB3hKw+JE9FOFnJJXpEcd/RsWrRdLvQcxvZYwoHICujDOA/aJA/wD30+onkJ
Pon3GsRqjnMvh1mpfgCCXpo/JcS/1vMxOg6LKJ5/qnZEVLIf/NKIQojuMxkth9qB
yFSXA2RiP+9rKNV33QP3WJQnD0/1dAF1gkDNOVOLBNZpA+7K74qexHZhJprKs73v
isPr9i38ePaeqR/G4gd2F2BJq2Xu+yDsbUgBWciWkw46Jv7p3NaNxFYi4y5iD2+e
Ahf7xOOG663JRhvOtgsSjYvxkOXL5bNU9TK49Y9c6CAoeBURDSc0hHD6/DIv1qad
icZeJfLSswJ8vGa/ypdIlxE90yA/ABpPpMDNcam4FDkGIHQMAg6KxpWjtaGrPwCy
oQIf9EK+7Jo+EjzCZlHT/OgYwkGqM+kI9fwJB/SRdhNAG0va8TG03flOwkstWntu
bWm9DnGBpR4MPdCa3GFQANWHKMSwGk+Sr/r8hJWH6NNK9PP6gFUgFaGOqaiH8w8w
sKJtYyeKvGfXNdGlYhD9CD9JdInvPhKuaJFc3SLL/fl2ALVtSYB8iir9vPfV7nSW
H20e2Ki7atYM6nVy/BAM90i040PJ+3G0n+MZIxmor2iJZcwMqnyj3FYRQkKW+lTj
PI0DbAGo4Hc1Z7SH1kk+6O1JNNWTD3bnEfEUepMkvIhKbprHhrJz3S+eZWeS9mSZ
gA0BQeWfU6AYVTjpNIxDGgrjkgV5MwjOXh7eHkvVDMxjQeQ5C5D65yozBh+ygCnc
snAACm6TkHx7lBxdF0wjXzc7bT8U1ufAGc2euOtwl2F/pPa2TOiuOE7LsFL+mpJZ
zLxK5ceKdJP/n84A0eLXXA88/DR9SIUPcJga320oWY+Wf0pEsbcim2S4n1QYoSxe
iLRhSdcBtXhklBBHD1UraJnyXZHCSOksljgTxyd33ynK98IHLrHUiZJkPiDgTn/x
dS1LkdoaCxjwFEPAHd1QEyeYFx/5aPW+t+ndgP7nELDgoa/2u2T/KkjZiT+NgxXY
8lm3HT8SvQ6iguXXpgA7dmGqAN2zMTx1qjwCEERucMI3WY+FBgYPFILwzCm+m+fG
L6gRhZwpJt4FCqbiaLXVy43Vz1sGJAPNxBHV6RTYxXAppA4ekDEElq6IZtANVvjk
Ve5JMsM62+eWmr5NAsAnbIZHUtTXxZi2jL4X6FC8sbpHlMduLqsml+SUqL5Vnp9U
Zrv8Lo/d2ii7vXS1PpooPkVI/94YwEj9cAJJu5lZEyoXW6zs057gRlluvhB/bWJf
uYqBU99Ti7gf/YJU/rRYDVpiWYGqIrSCBd/owQCZzfDqOhAFGuV/QuFlFV1yHJBp
n5iK1I4bvbxniIYJD2g4lzn0az0g72E/Ifgr8f1uMFrRXHNvr0uAVpdT/29cA3TC
fyb+X205F1sFOLxBE4Ii8T309eEddKuHPouDV9YCHl/DqFNX3SACvHr9b9cHjTlR
aHEiy8/g9/dMqaY4BpFBuQivbKxpjy0zIGflqfBy5DEmVrKDJTe0B302vnLNrtNt
8h9s58T3W1v4CUkvvJcYPtdGrkPUYcuLMOCmLAUtyVzOdwFgc1Fm1XOlOEJm37jz
QFsUZhR5oijRYgpIQ3bSrUZ5REa+XLNMrjyDKs7BO5tRXVG1c7ObC/P77AqZOcRL
opHMSv8EWbAzBuw+AUHxiGM74njUOjAtZzXVRFdPVeLw5ikYFftcOE1/PLvkAp9f
AjoyVzKo+r1kCMhiKvorR7HD55a01AGUNDVbCMwmA2tO2wDyNeADL3EaxX22ICsx
G1qiVpbvGsAJovZNSc+l6xoF2xOYbvAbiLiLDOVHMOI0+oq+2nCXm3dgKeon1r62
2h+iZ4W5GMfMHAQ+9Dd9MCEIOufB6n0c1ewe9U/nl6qp8xD3kN8LvBWNAKGUIZZq
iD9Nd15sorJZRNcU9fuZ4zEdK3Gr3H/hbKQNgyadl8fg7VvUugAC8Q2vnvE/e9aT
dBzbT/b1iCrKtGEyBmz2rYfB+geYx+gJnt3IClyDBKVUAz2MNdzyw8fJLS397LOb
6LthLZ1TGERA7iUwiM7JWqVTTUMQd6Tt1OaDG1i5r7UkxbPhjg6cbjo2OAEUnDJb
iyuxDdlhL0UtmDjqAcFnZtj4iYK5Com4Vx+1wjXS0JphIHNkaCvWnmMZnjYyklU6
6CKuv+iieCMzKiGf6HcVlZ11Z8mtesCYCavzzx4vVWA826j6mTIkt39gdUKXLNOk
Cmj8/XpJfrb25L3E+ATWBMVuf1wb2xc8Lx9DbLz++Ixeaf/YYOMYigfZST0W7Qdk
7xHHYZWa/CJDtF/fW34qfSB5dqdpRpHmfe7tXI2HpBHwitpfdbj/P0uJGumpHLNG
XIInjyJ+asVsiwlpNjKw8fs1pwqOkN7D5aVJLiALAlEjDBdsFGbUBI9d/nKNeNU9
u43es/FzXhNy5IOfVGt22lWSsiKKklBIoMhaDJ+haKBnv0/405CUJxqzHlQJdNXU
TlckpVdZXbtk15klqz22I65GRlMhZQIbrHigsWmfWaEwFyaoofIc9w0Ze/zcw1uF
k9q+KMFzzFgtKAgFM73oro0pUKpIxPeKxrdOyK2pt9DEl+9oYzQe5S+9Ylo6RqCA
44QvNlXTg4uTgv4Wvj+HVjDhVywHZ8BsIrOg5oGn179PXG2qd4NbaxB0eXBsJosN
Ch+v2c5Lxs3wmHYvAIN4Lmkj5E9ewrPNwb5O5XF7OFgkdce55d+XgYPdzVn9HWSf
VvB7IQ/6dBzDpRbooYfAsEWmIr0YPrVjGdDZfU/JB+RA+rODCQuL3asTAGQZVuNp
fCqWDAw7DCD78E4EwJHNs1AIpG/p8CDxLmgyzcKx4LuoTY5/yODoRkouO169vcfW
RpEsE+hKbmosYqy9sZSxM58eil/g0hBzonBW9rKYP0N1UDpQFM+xSBgDWeeR0PL5
vG11MfAme/SEss/QWZKSr1F6sdsHxLCwYSCE43tNkW6J3X69s+UD06wccfWlG9+y
KLmotbnJwU5mHVo6g6JGitTcg4kF3DywAQXJzRxFYZJ3/R6SGb+qCQ/XmRiH66+z
NuzhdsTNlqJY3CJ8kXhGQlmLQuTkUjKR+SUCMlGFcKwKjtMd64ZWMIFknCG5urjp
58G3rEJWiqz+LU2nByavThUduCF/rurxYaqbka6/YWuxwMWBCeDv0LZW3osq9hSZ
WLfSjqAUkXFw82wMvrqtaaiNeUtyB1wtNGrR+To/AtNOkUnf/e9KpJUJIYdTalq4
TUW9Evocr5RAUA/AAoMqCRUnYQFkGoSTdFPpMTw38wKF6yKpvTclPrXz12hc7lvo
mDqvWjkMErd0Mxli5+19M0KOoZsbTmbfOYOVQ2WPuOy5+0xStghSmaqxN5AGv+A9
PKCEC6B9VKoA8WoONjiUM5GTtx7YXHDWBwO8DoYYUCKPHUQQrwn2KZ+wkfhk/Ko2
IepW8B9OK9Sa9+726/GW8D1iUzogIaa8lgf1x2beIE43f4v3deijmF8vdXEbnHTC
984qfSjMsBDG2eFcxP+0pahqFIXUlohSpML7dMaj3Oay0lPYqp2+2eIAUkPEpXzY
xIdJGO2BjMzhTVQZU9MnuLxUdtMD2kW7bhIQjR+gZ/4iHhjJUgIvlDC5d40YrCOj
lnw3QnbAGOtJ88LJUoyHlXyosfxi2iqcJCBdI9idNVFeyQdjkv/FiJFeibGufRBN
qcxS1G+//xxrLWSTsjfzFTjFwlPQozv7nEwPyzYJyh715aUgFdfS+Zq2H782JLG1
FaretocBtH9LoD3/U5svKNCDRLDY6BoOBXi4LSQCB9wigh2sREfj1rz15SEPBO29
YD++XLAIR57j0fG6NsZEYJkGx+YHl6X7C+mvEmFp0I3UEVLHHNIHzzV96VZesqfG
Q3a4OkNJVyfO+rMUaS6ONbeRVtnOz9NJL/RLQSMsGKWa395pk9y4DoN18UmqfAix
CYywzh+Nn5tCtJMHKEptWW9PHaF+H5hZKhoiEU35amzBMBE2LBM3FwqPfGXpOQ9C
eI7Y0XAI0gLbjkzR3UKzmrnkFl5EXwgHLUcZi4lgr1w5k/2couVLNlIwgnCRZNWf
nsKbLIL1FEYxSvIM1n5S8qJQ8kTUTXO+TkVh99BGmuHLD1XxHMmXhxbgmKW9QsDM
nJr0AepNqxAnkrq37JIChkImEb7EfpRz2VkwYcYROdQLw4wqgWwTTI2fZGgeI/x2
N28abgvoKEW6R48Epqfdg5WnnLmf7B/npXB6K/e+ntYKoDLhrtIfGuVIrg1J8w2b
fb3oHN6rZtte55pcgBm/X12xnrEGPUHKqyIQHmPAE5OZSMR0bSdiPTDoQxXzloxs
Dz3rrM0rV6FZsp34ndIj5IMUf7t4Eu0Z/5Fy77mRgsZxTzZuVJSuu7mIS2ezcaMM
3pSYu8DhxOuID0lhULzD57m3Qm/UNUp9Bganh/JOj3ViDiv385VFm+fcLv04riRx
UwIowvUaWSLig825qz43LgYkOuA8XkkwJhL454xkyg7A+a9/syLPf/6LLRDk2NPv
LCszN39BBtpvJp7CMOQZXk09Z9MI8QL0x0mQMcDq/cPJQ32v3lPnylJMnEVOH3PS
oRRUpjEve2t8sK98jKFVUnHCY/CCSY/Own0lCyvyJgfBXunj0XOrgWRLoVTOgboD
hp3v2bP2vpu/ZMEWsPjveUL+C/KBEm1b+ixX6Ub4eMQwq9k/dhAoCeWZT3gs4Qvy
2ifVI8kV+D1H4QQtYUj9Ijy4CKQRZQgrHLGhzzLVxnGIMuMCm89WbS0kHUTGlj+f
trs4ms4ZRnEY6wnLLSNQylLxm9X00nLvdF7S7DqRSf7IRyodwKUWsJ6fQM/wMh0Q
/n9kaA6D7K5+iwC376BNlUIVseZlcwrZ2aqJGpt3RAPVswxaJgmfLUyZLncUolc/
qLjpuGa3cFinbhQJwznwqq+LjT5yP6XsYQe+odW0zOePraGNuGOVjCilFeKJ/NOz
gPd42yKs2/4BA28ak9NuX8LgqKMJi9e42ophggPqZ7TqzPt/uKAYE7+yB+yGWjoA
Ca5V0s/xE5U+FdJ7rZtX22If1ZpedJcjGxjjlTtSw5z2uAAZg1KKvkgU0EJm+tY6
Lq84Zr+HxybY9/8EfqRnOC8LxTKR9HgtxhdwVGPvqiskMvQ07Lo6dcfHCQw7tb+r
hAgTjStOCJ6EST5p8vf6BV2waWQ42OSfh7zG0zG77Mjaz3vAFmnA/19sZhINa+6z
f3RyOY/sXJygRP+pso2K91zwdlFTAr/3rHVond8qZi+bCy3KgdyW/ZYoSUkO92bp
nAxotWyD4ydYDUUd4uQZ49sJo+tOAKKJIcyX1C4Af9dJc7s6ip1pnysZsAzIrp0e
tAaLcdu/VALzzeUUYgT2jZ2xaws9aq19V1unlb1yoc3cPRlyQ53VMQu6My4gpweF
PWHZw+LMAYRq5desYsPdDj8wCRqnNtCSrk9FUquEhQp7nRpZKkesJ8trqYz/m45O
29xDUgqxDemrWHBpQu9iUA6JrzVHquArzPq/NO8zxJhmmLWLBXs8vxWqxh1DhqNX
qpNGMXBveoNEpzJ8GfTDS2IS8wrt/33drvHr8qQ6r2rHiXuDsYyvomMS914FDIM7
iamNv3MvjnHtbGVsBLxpS8J+m7+MtRml3JHNj5qSbFz0Yv5xDLSyAUwem3ftb4AL
c68Ji3mr63gX3b1nokXh02r1vAw70vMlt2NW0/ncLLQRd1FCNvZNlV8Ywry0HqwM
rA8VNwwmKh9UoBpvkQrvro5qbLlmBim9O2DS4xL0/+zl8jXz1ahX+mUL7/YBGIvi
tnC4VCnwFVCOZ3UlIBc/m+fVmn9gAYujBwrr+mbwZ3sccQucg2nLi6/4gj5VcFOn
6ufPbKi2MmcwT+HFGPPjyF3CqpZg1Ty3WNmEMT6eWTXPhghPmh7PCr4b6CcA/zcc
NDapQZZkKscstA4t2NwiB0FTdXefLp1zVhlWVoojDDpFQNVOOgbHnP5ETRMjSLO1
7J2XQwlFflezdzVyOW9jatqFEiLzoBFHVJYDXWCa79LBqhzLkDTIPUvNjw6Cqd1W
cc8MxicK6Ix8juFUbQLk1yzyt7HF1yM8J+ZyhpAwJK84/ajUqkXHa7Ax/w8ZXpcw
IyLE7uWU5vY7lMA/92Qex5JiTXHwG5+5kUwdkDuDLwJH4QBfvDGOijnB8n7xFAwF
TL3EhDTl1C3VDYkOWdvmvBBTlG+vk29a8RK3yWWQajM4gdsoUKYL+0UNG/mgTbjI
OztUejp25MUm2vJ/DS1peNePyJeD1YEi78pE/TsShLoMXKbJUBTBPfmSri4q/L3R
L2SU9bz/JDfitqQgq8+DmkEKPKzVvpE9fQZ3qw8l16gQxro5gcKS5/7DjToBfWtf
xJkcET5Q02SAcFMt39aoxUBXj4FwGyVNTTIpCjsly+OhwI9HzjzuGLKOFGQT/pOg
sJRojrR1kRbtDk1hP6vHnpNhEXVjJ4YMUW5Lx7otFJoURU4uEGzI0f7HGhYjLX1x
RCTm0g49YS+SI6DOK2aMZZIXC+hZ4DoYrla3iosvN4pQH/Iw2d1Z4x+ZBJ9d/uZU
g5cO0Fk+68c1XkP4OzPuiTO8eNBxp6tog4SCJbjQBbkUaCoLq6G8rSxKDUQGI1kb
+/da1lV7fOsCV8iBDV8ghuPMR/i16z85+9X6ylmwITditjooxQPd9Fr9FGqi0lXR
98JoETLLsFrhrM0xQe1JBXaAITWvzHe+PdYTZ+zfx6rDPU+EMrA+MO9y8xGLxnHA
QfqBabfigbpy/OUrhnOWPRYJISbL+Q5TDDcCxFR9wkfw1JSeaG2Z87lZveHNd97C
uhHMYxkylJcfYsPh8qeMBRbQwaGWt1Bq3Zfbz5Z9+cCNjajF+NINP8vP4/FfP/l4
sZTatwxCi0OMecr4lZjVkRqwEXT7pkwDosp3qKc540IUsSmfUFHylDe5VnZxHV4w
r/305VTqdZ8kXzY1SLLFu+v2ULO06prH9VRzv7qwZecpoHLo4jdyDWRLFGCyAGXo
WjVYHpCkSMHGyb/0C12ZLFqRcBTT/nuYLn9e6Yr5w1zJqXUN/Tfl8Y5KfpW1HjYN
IbtIw28cEIGwsyD/wzlwm088jdkzLjV4IX3rIGrFXmZAh96Tu5mcK4yRlnimX7vQ
uregOdbC6AK2NPGyDKGZ6S1JO6J/0dv6TGH1X18ZvlrjhYnEiue6OIVN7LRkKScg
pk+VwRhsbTy4OyMOKTD1HIc4hfq+TQECPMVLnaNeuy0KDRwKAka4xArq4YMKKa9K
taP1ZcicY2E0FSoxC4fuJ9xB7RhL39BcZERx/xAGqDphRB83l30Znsy4uWtAU2jA
TLtXgp4xz6r4dCxH1924NhhiHyx+TnY7uYKjuY3Zd+PEEtAMmVQrVlSff7o9MqY4
2opUOb6SQS/zsfKE7I22GJMDxnW14FdN1WwyiBWCJWjdpYA5lBRkFX2xeX3AdmMk
+rDuHf8a1WHQHOa+I1ZWWc0u6Ftdk6nGskzdaqs2ahSZiK5gq5paStO0I3pSXC+s
A+73C2I5TVTjSUSUwGUA29xceB1azz8eFBybf7lmj7qOhxcZMu0NPIwMqQFGpC9v
hoQe1mpLB+9HWrEZDoS1R8CQjhD0JiwL6NpWiNh3G7R+QoM0Mol6m32+DUIE1BFo
4AW4lkkyaNvKb9hILJAfrtBShqOOD/m8qwBvGROBa9zNOVYvpiRH+syDBLcBigap
iYPckLf+t/NQV4OF1JF/DlYczxJHklRWcJEcQwGD7st3MWHOaSfVY+X3A6Qz6HJX
HcaPOivNH1YV/wVjAIg3k2rBbUynP/S6SRZeaT6VkoYE7SJymKp23Ic1w9BOBCjS
kHlCwlBhePF01ZGIseRvoaIJh+ColxROmLTW+X1Z5XzZJhLtlM6OOsKbVy+9qJQi
69UuxTDRUyO/qoHsbWu+hrJFGINunPxCrKUsF2HIRKVu2Lm33rhmA+1qG0rT7iln
6WZ0/RFAkyyoKa+1NOFhBzPWqYZfIDSJi3vwubXJjZ3dhEXJZKqulKL7IxqhVc3l
1z8lMeyaXyQyyZSKqzKhiDDhi0p2O4+mgE0BUaa/S1pe3AxsC5G5l3xCDzxg2tim
ZgQ8jbTLaKMSD7XqRV0jy53dlrTE/mRmWxkReC83KTjfXgkG+pXoZhW60W5Z48NJ
XAf/qx9j3GKVfTwcelXQm+Kn2OiFPM38PKlr4Qy11GzApeAryK7f1SDDXBATTbHJ
PGBVwhn9iBWrFM35KyjkJL+Q1GPjvTtDqke66CwS8x/gDbHriBW4SxekXAyX3l0r
0cubUPe1/PVQRkOUs1Ij77huFGe56GyAkPa22xIjnHbCtqBVUlqNL/L7CaqVLJjZ
TEuiHYglwUw4D/eVp4MCKOEHb1v+KczJvd1M/jov1Dy90yHebg8Nwopvb4XXt+5u
1P1QDgj+/3qZE6yboXwzExySPIocVy508+0lnv3sqJbZDawpAd5lsY+nZjdzgn5a
W5MHerHXG9EYAizPJwk2HwRTj8B8/Q9EJSEmU/fPPVplid++xsQjoW0KaHHm2Slx
dTAeOFoBkMgSvAFH6iveRVRZp8sL9GUy6ZKHE4GfWQ6YL497breEeJ8Lp6dCxhvJ
YahBAhzSa/zW8AI31nPmtt2CR8xnfAoCnWsJwa30ltqCwJ/285NxuQvv1jSeFKA1
UNr59R5r1ycYvhl8egl+Oe1Q2z1ROgdQ1ZR6iHxMMRuGZBOgL0D6WR0vX+D2Zj4z
mOlGmzv8WUHGOoCAo2uLju7ROzKlo9FdG2RkCr4wkV84Sl+SC203zZJXGvsL99wX
mBUu36geOMYIX+JM3fifpEuVDYxCog4w68mE8OzAvAIgVK8tT1yVJ/VNTdQegV5E
460LHev+JNdtsjnW+TKQwjyjCduUO7nmnSDkHYfBPSXaQrLfJmxR+74Mpba71T69
lQrtduQ2usxc/KsHW7BoHuRlXBAmRYalqwWYuBpNGgALLKNXu83r+H2mP5lIfZSi
OYx/NfDWJ7ID7mOmRsESmy4TqQafMSlmsQOKHah/7PlVC+JZE3PexZ4HeOVeFKyq
dlZ1CXdBQ/z5Vbjs5j3Hjol1if0vfcYUx5khfqZcwmW/BdUsWX50g71dZCVpE6ja
5zEfEjjapJdMoWLfAMmUPh6O19IpSq1QTQPzG5aX3usBQzjbl4fV3351J0gk8ZLz
DIzLJuZzq2ynDzJVIWGM0HX6hNQtExPwl86fWm59zyzuhlGYugKkVdc7xkZnTxUt
TUg0KVSMuniuv9uc8dHiRSCg6Yj5PsmiRKz51WJb54lQ+OH0pWpK5zMlQmFMGILu
plIv3f4Qqq9sdZzquG5Q1BlY8IPt60BjCPXC658C9fooF0qorS/w6s4qrYFfABnh
J+XlidLAdxHl3IeVCeB6m/e1n2KHJfLVyLUFT86PTwLligEB5uBZYPzfP+cobVlI
TCadfVjEDuIGFX4Mq487tbFseUdcPY8/r2kExinoRWhFwgdFriojpOOReEbMU/Dx
Mwsm6HWx5ssFcvXXYXlJ/eNDHv9NMCm8QJppw+GSTCBf6dPLjmXfUznxAP4x0MB0
PKlTIjPcBA5s7XBkAPVhVzkaX5sXSHHairws4EahvZikwUQg1JN/tAsJU/ey/Tdj
c1MR/RBtVrZ7+lQjGdbwPGKfLKqe350EfvBdNyqPoZNRzGAy+Ke7ZJi+ebYEMk4l
0XyUavPhgQB00Xh8XBPxd9aeP2Kdts/4ZdeEPfjdjc7n9uffMY8FAalvnnW2yyEb
rV28XHWdmodeb/RptoLPW9l0HlpESJoIji7ZK8d6krdk5WwnUABgyPD2NhvuxR2u
Hx1uaM2HLtFW8H9z0LosWiiNUovcSrFgFX2h+OSNit8snXxZYIaUwo1hID8HCRZl
MtuBTBOwg25tg3D1Tvu4YE60PhGZam06HVPC81vPsbhoh8vlZecvLx6IhqgnMdIP
n8+KGxrSUKTZSg/ES4zvEMKNjQZURau4PjOUxxJnAKGad1ucI9GVUKAJiwexW2cr
ewgEQR1K0LsSW5XThv1opB4pkSCbH+K1Ul3OOfhMyRTFBiBvmge+bH/3svABvIvv
ya1nh8o97XGBPm0zVdggskyJTMHN+GM4B7IPjPcG76d5TJBDQnCPyAY2oRW6it5R
xmUAhEsRoJF8RM9K2Q69KkIneeFEw5kPKK0UnVfazp6fPPaphUmwbbyn2NYEmM7m
hkuLE1UQ8GQQ2ApVlmtIV7O9YcSvLSui9Qwzlz6Jwtb6KbFSYDC+w4RTyNr+vuVG
I08vNDzCh23nwLAQN2Hw40evHDvGvu1nytX+C2Cz1dcW0YZz5qBolZvl0OG8EMvA
VSuXIEMZYzHWvNBRmjdEdZbVmWMUhm86La8rDZdfIj2LekF6AA1ztzIZ3hAq+wGP
md2cyoztFgDXoV7qjz6reVJnFEiJe6+WU4xKMzSrVywiW2to1NbztqeVKvP3rW8D
0dMGZhs+xMiF46Gydtrur0ryFYclyn4cMlz2j3Vyw0H97Rxixv+MkMeEReZUB1Y1
IU8HzNt/y0nZVVJR09ruOmqXE7NkMhTmdxdWVReQ1eRKJaQrzzZHTxqFMlEnhZ6Y
QYBXj1CS8qqBoS9alEQOsHUEjn41m6EctiRWT+nULI0MdjtkkC3w8A9RMo9aTNPj
99+2cqAPh+1mvsXB21qQhesWcGJWvUhQDTjoFdmHcpJ779L3G5BMbDzZaVDRwEIT
G/p4/PeENffd1L+ILa8BVWkNRTtIBnVJqYlkHLbMYLC5hiyabqFVOgmyySBLpaJk
Pa44iJxmPMef6uOY7q5jYgtNxy65A2A/iqY6PAXSGR4fYguktyEQI3Yg/tsjS9PI
/7BD6R4kcA4D8ZRoKH5LDxSFN/xUSJCAOGUYc2YsCEahbwY6nUFwln+LRthSxKM/
Elscmp9t3jISjxs3HInffHj2djMJRMYxRPCBz7Wg4smumzr4Ly351FRxOp8t7woF
5E9WyX6fwTI+mNS7GH3qIf2anEdzpUs2Ct8ZuNXvxQuEyfHUaqC4urJSTHk9RZew
4GtrBgei1J1fqzH8FPtEof0jK5uUB8SZ/ZEsluNQh7BBmjpzrPeGHxO97jurHR7K
OfsggVQqfbMMFx8hZNbpFp1a6753fNcUtWnJX0iMkjwSOCObT6UAjlxr1kpNctHA
C2Xz2uXQ7YE1d5HmIf++MWBHVSazffboWp67AEvzqgaemo84e/ex5uHRz77Obfyr
k+ly/s0UaVTc/J7F1EUPjOWxnN66LbQySRpXXLkDvslCSmV3AO4+PeUdBavpwr38
/2kmYmRB9lAROXUcnA8dLbAACNp4RwF/w2rXOywwRz6kFZsEu5WU8uYF88JM/fNh
u5fS/PU926o+nln/Ut5fR7evxlTi4jSnSI8u/JZUsIwKTrEBHwU5ZAZ5nVmAEfJD
KTh2pyjKCh8U7SgA1GNNhGpRaEHhQy5jbdbP+gPVg1LWn2ACVMVbTHcQ2wSeHBfy
cWAsgAhQMhentdGZK7BCyUyB9pNtoT7wmymRzz65N7uR2TMaO87Qhu2zj9ciroxh
TshHB0hUIzQQGAC5rA3VsFegT11WEBPEZ27eu+1bxOKaz0OSSuZiKhhvYT+RbTM7
6Xci4FgKIDCtJdfA7cZieqm8wbyrMaMlhuT+c3oqh2o6kcllV8MyzQsCxY+qPLen
o8cqp6eihLxKfOk/u1xi1PmrEGmngfUjj2VkUO8e0CVWsZlSXUd3vMGykJSVLmqJ
6XKDJescA3lmpSHdaDdcy3rOvVpTf7GKyYi6XRzdXgGr/Y1uFAVly01S1fJrKTW9
0WAd8B7u332SP1Bka5JQHvqiE/H5Ycmflh3CBzTQMG1CNVfJdFkFLSqzoeyH3NvK
yX+lStB6wHskbAVM33Il071b8x0L/HMK2ioGpAaXqYDiLLNXoJe6rX9E/lcUhROe
dubQYjJFBu6U5lSt6iregWIDCY1JSgs2YbgGu39Ir9IsernSl23WXdAW2lekm9ty
OtIF4Y4XndNDpg+cYVkZPvcqg62r7uSBbB1JUAXtJwZEglvJJDvPyks27y4UNpbZ
kBPZIzX7DtoGxJ/S9bGiGZNg0YDnLSTBX7RugUq583pCCQtYAI+jcoqUedGqUJRI
5GwXdYR8kLaJbJbnHB4ZUaG3NmOdk4xALlyIJSjut/iMMKErrsgXGdp4D69GPEfT
O98qN+KyVJ/jdORxDG6p0AxOTzz21z4OTqKFLJgxNrfS6Ij4PIYgvAkMbYbd41LD
LIUEkG41T5Ei5OOFDuac77mX37Y/k2s/dNCf3HmQZksC17ghqtyK6Lto7503afy8
SYZrRttMdZSLdmyecJjh3ZH4LGkf1qm93/SDCjbaZ1uya1X3GNbHQXsTpsH/VTHM
jKN2Ym4PYJTmtW35UzuF25O+dMIKroKsjcClsdzJuljwHKGtdB7JbtIvZwMvDfFZ
4VyJCyB7sODTwcrFQDUtTrnJ47XGdBWxE2Mywva/JwPO8rYGeTEZbIIHMdy5I09P
hmRNOR3iBVv6DFnXyWGVHReffDmSxfjNsXyis19YHE3KV9DqbQL0yh+fs6FZBWiL
wSDZV40Y+w80vUxNHktwQwFpKK/p/fPqZ89R4pZEFCC5M969Q9vB3PwJ0q8EtIjH
K66iAhiF0n+EwGkcqGowKV+lLl2MO1MYuKvpAXlCNUQTKw2ILb69qSOZZ3nVxtiE
6V0q4Ug+s5/iAwSe/bCTXZkhEJv5YpQpB0vhM5OfttDvRsYOQT0Kpj2KMdu7BtTw
B4sR1jlQ8RQqBWC4qGAojhER0JB+A4CEeWDAr1CWqNi9VA7rb2vD//DTCbiqK3h8
/nWruUUpQxBy8oDmcR0FaaxbY+vxvqI6OT1xuc+6vxkrz3TlHdX58xaRAPoYkhHS
yT0kfMef8X39D/q32PrE1FaqpFSACRxefp6bRRlPWo5+0NjVqWM4dC+y1bwetw6n
Af+lLp3NqFco0k9hlIRHobCcInyV0W5wnsX046DNa3KuJAICfWWhPo1zPx3Esek6
J02NeqsiP3tTcP1DqoI+HlwhjdY62M8FckfYBD5WaqOvE2CfFLF4StS+LxYKangR
nggJ4njbax5WSISXuiJdqlAnyfBTzg/6Piwqccd2iCM6oB4/aak+F4WSmbDbk7OE
2h7FRIUxLiuKazQZHJMinSTkgGJrk74de71yyJdgrI51UaGk+hxmdNrEb+ouXEI8
6v85YksLSG64lpZrw3bhdUn/HYBKbFC1PvgNAvb5+UrqsaE+RZjxqI3jcykTyPt9
lDk0xqynBEjV0azDFfvcfMHUPyCzdSmWl5Nj+9IWvbBDo13zyyEG8VW/Mors+qmQ
/HYSIe09aVVTN3/3HJVoO+sH2vxa5RdSeGRcHHh+HqvXNOy2PlmO1E5sIQIKY3pj
I4QG7/XEPRnz4VvYQo9oqd32I79LpTDUqgItrWocf+eKgkXMsOd27mUaB/Q/o6w9
EToK+56pKOdC+tPYxFUIUG/CmMgbbdCfbs7pvoyOF3nu9u7rYawgu058IOQMCzaV
inFYRB6ofZNam82ZAcmFWBECyKkdUsybCSlFQdQCNKsId2tt4nbyHe12IFZS80MW
4aTJY4OoeukFr6GziNNkPbWNnZdQiqD5eK95wl8eKyQMvl4Y7CV/I/c8SjlmTAHI
1GXG9cWHjZBn2zTROzY6ul3Co4aes4ZWDAnvQkAEpHJGLrLubOvfoXZgQSuCZViY
5W91hF5Mf8lG67yj7J/o+K8DkYIQLQ0PHrWCqw+wFwxA1oDZDml83kmqWFu8iwfQ
Tbj9uX1S9OjQkcqmVkiH6ChWqFW+Pize6Ki1DN8MpYyn6RHrjbwjgvhsD990bLub
9hMDyJmM5PG5W/6b8tykUiKLxtx8adlkVZzhqmxP6P9iVt79bGTgOYIRkFw8jfZ/
PBS0cEZVo0cUrRjsvBFbfnAKpNRA29/2YboRcBZhydJ0KiE639Xq2BNzFBkVdGLF
hu+YbI/X6BgP6dAvaZ4Atcd0twT9cLtOoNScnlfLl3fQMQukqX/NDUaQsckZW+wl
B+5qRD8QuQMvW3rEVzOwBnzFr+CmQsJmJxc1DlcQ7OrS7rYzNyqrj8FzVfXtNzOA
Ie1IRio1whPF90C/uxq9usjfD8uYIbGq6I//+Zl53dGjIX1EgnSM2EyVI5by9YCj
dFFae1ZgJehSpP+FVtkC25z1FVmeosT44VU240BSQQidUdLvbqRZWBWoWZLDLyiE
89QoL8o7E17Rd2rlu//SM61szwf/WS82fb/ihKPvol/etNSKqL2SNiN1qYHpM/Cx
LmqFuBRyUwsnwOoNbbfXmCojtF1YJcpyZws0+qNwtoht8+wA6wg43mwupzAemG4d
NY9KmewKxMsFKg8vAky3651ph3UDgBw15qkDJXFt+XF7CiNk67uEIHaE9X8XxgBr
dO3BeRvYRQtYoBs24I6w7HTbr9HnXNooAfIP3nqKoWarFwf69RjabBn6TvHmZcFb
qzSgl5dQ7mJZCfRTOadl61Qax+X59e8JGB4siQeCxEehYRUXt5QSU7I2VyuxbLSL
HAXZeBIp3bjNIfWmtwMBW2z6g9u5ZHHLEI7hMw2sXuKDZC7c4sD0keRLj/a857dr
AxNvynVLY8osTgwsU8ZKia78nmVmbT+3Fonv1rv3ndvHuTnN89msU0HacqF+fPDT
xHnbV+YwL0u92dpLDRAZljxkFI/XRoBClEIJ+bO0M95NhXUsu2Vm6wLt+6q4iNHQ
w9z6RbIHvzFKEgBgQgEkf7ho6eLngy+P8DO2juC+RUqUPRb8GoxY+rnOys94B5Ag
c95BE0vGjqBuCuakuZX9KqepgAEX/r8k+Htuw4+zTBE3ZL0TF0hr9YMlc+Ej4QRf
fWBSSdKaJTeJUWvUXUvdQKwAaXY0a6tUPJZ9TQbnqW2b6fsxIryX/svEQBzOoPeJ
rCffu7hQBenqZgi3hIbcupyO4p4C/RDr5jpQuatdkXzll1J1Xg4Fg0GgWXEaWb5+
m/EfmCSVlRFhs5IBxCDgz5TBDX/anQhvMY1sA8Wrr4ru8MKs+ioLkUPWde6GpS6o
4K/741FJlg4wEP7FPgMooU52DgfgZVnfdSQzKhoNbYVEAarcjZkCcmLBp6JFKka2
JAbqq3w8qgPxF7qK719tPUeBpmeLLOZPTWE3Q1SZpqaGQ0BXyIXtTY8MeSEjqkZ3
pZ6ZvhgaXuZTmDN39f+8U7UDTQACMBGkxJaaVAVI6CUs5WP+gt3MyluVYfjw3JKc
pkoKQe4YQTMzz9cI6isGXmAR9BKkYCRjw+scXHpYkXhHlS++0VCtFMQHK++t4V+M
/ZihVApTei5x6tw1SFQONNL8x0m4OEPTeIQ80Iul4Q8TJUQ6jV5UsSLxAX0LakFO
znNvEj8jKQMN8z761PWZ+nYeoy31BhhwUu9KvnErST7yaOc9eCSLRjzepYEAQJ9R
6X5N/UvFS4q18vHBXyq29Hdl2/JCJneDLrfz3hXc14CigyoH9mBgyhokEtmsRjgJ
XwCW0zi87gPu0aCRrJA6XDRW6poKrQWSyj0BgRyX9ArOE02dD/7HkfrkvgQaRCFH
dP211bwz18F9DnScMf7GnjlQD83PfFcmhVdpKP4kbWnStlQ4LlcfsKN+05FOZCYD
agRaJ+Zmoq/HNIZ8QJhTOewlzNVThNxelUK2LhL4OF4xzUVL4BCrt43I/NzPYcL0
QWP0otc4hlSeDPbLuzofJRUtNGyYNrYIpzkw0dO/rzGzhOB+qc7sQiU2m/+kCuVu
ab/FebQSvKvC6kS6V0FxOjbBIuWR+o4R/jDaU//AMjHK/UdsXy9drHnPHt3yobXN
ULw0KOV0y5FrcLOqR3VFZRzLb74/xFPcsLCwFAPBLOp2wjQQJzlEFZSOR5XCbSA+
B4LcBe1lhV9TyfFht7ZI3HBDpWGFycxED2p/zjHuzBxmd2LW0aifFwh1O6DG+n7u
EmaPeVyRD6/gviX/wZS42M4XptyP/o+buikVekv6trAv54BfR181mCWjwMB05waC
/5rCuyKYjcPAhdEOW8DULZCNHYwb/JKul7ZGz6ObDGu578qTogsSdeyIroKZd/5+
udwqQrTjuwCzPF+jKBwEnsYkAgfsylMbKYnP7x+OHgpM62AbCw2mroIf47lHnJs5
KgPjcj3dFKBLicE/4SGvOis80w5Rxwv+A0w2PA82Gm72EhpvvW5qhFWVDLw2CrFn
OVdRunjtJUFDw2QNe97Il6B1cRn/BD6ldfiS+aqBK55S7wlx6GBmKZIqEsp8bCk9
Wv+jnPJxBEIhNEBjnTpIXL/N3jcpP/qvKyFPFasKiHmOlpPx/HI8OFQOhd145QND
c5UClPkvs26fF1ouR+B89q3UYhdm6vLia4FPjylfgwxE1cCBmxFb+Bz5uurywiEe
Ks9+/Puq8y0hnOgUNVwwrSL82R5jUT25i1xW9oZcS6RSbPBIV4MYG5fx8HWR1y7I
3UHHAZMhosyTKlwpI2Ua7mRH+g4vnYGlImnaotFenrtS3QBQ0seNHbGa96Qw4HUL
OVGU2Hnb3OaSZn9j+AtjEsx2SbWcqNgRQN5olrOvKPisHDyKzSEI9r2j6LJ01NhZ
4xT+Eoj2kk6pMQGXeXIoorotImg2BJ2hBOW+QSMp4cy9KlV816c6lt7fGYF0pD3G
C/73wKP+Jwv+j55OQGpO7zL9qrrGFv50i6Vi/VxSGI9oUAcUzvl5sAtj5x8E2z+Y
Jd3L5/k5c2Rv9GJSsVLY/RC+ZoLGsjrvuv3T8yHKDiWxMXu7wcS/+vRqbqnNfVqP
URMD6JifmZfPX1xHQ1km62otDTaYO39I7zkbNUh6GQR5YiQtvuCgsMqb7GWug2u8
FCRkicBRo7XDHf2VnFYaHv/HGjmWnc9OE0R0r85kWYp2cqHC4XiboGU+M84Q9s4v
tqqS9qFC0LQE2OzfLRMXv6q9CN/kz+O6YnSgpBijykHdxDJQSkLG2wa+/B4kN7+r
sVW7uUHxqILBDc/D3oF5GqNfKWj+Qk8QuChkIZFh2hZTP/8d+RAiwvj272HX0Hq7
u20Fb62NMYyszWvLkm4WW3qVftvyroyX0tjA0IyIF9XB0VMhLZY0RjubHuHHZIQj
Evm+CQSI70k6/5u4oc5xpWSmTr7Qfp13W6mDJXApnJc885rfZW2E6YoEtnHo4TWv
yVXzKXyJu1PcbIN+an1d6skLlNFkuj8F9Fb35Ul2BqGnK+9YfzVjK5T+fTe21hXO
cDsjui2sPkUjI80QJSZTqHInFKVgfTdL05DIUn7TDfowsyE0yy5bxhQ8rtuNtn8v
o6XwV373oDMyRjEOkBlyxjO9OCdcxeEIUe4viPiQw7crqwOuP+lkNwla75NPDnek
OOIwDJ4Yao5JrDKDTMDx84CZddN2AN58erELtGB8L2dRR7BGi+Tgebvuj17kx2HQ
ki4amPhnBk9doqm/hlgUwy8LV0dlH0aWlAj11c0aPVwV9cU8XQiJkLMpZVlh6/rX
PfVCjiHe1+S5IV50T6dN4U/KqwVAPebesqRcy0x6wZLJMbGe4cZuYQRdb26V22lJ
zAABjrVbOX33s+pqYMICuqPJ0OACE5VM5uLTUWAjTPeS8Tl3pto3bNIXuEXnV7d3
2qdnNdKktvCbKOMrhSJlKNa8VXb2aOjKt5GKd1tmtPkAscdeICb6VjQBPvSvdtH1
dXVsrYlNXQpJ7HKXkE0f3lzAjJ1YB68HN0OfvTbgRCJ8FM/LggWDdOLC++yEpS0h
uCXu9LZSIiJIbXNV2mr1VaIWB5plQW6z4he1j5Qsj1M8gyqy+K55lKesntYo1JIr
W2QwN0zyxaT//9tQsY2hXsZsxDsn9EkEj4NCJDkeQsAo96hhKVmo911B/SJ8SOQH
ci0D6p4XjPFzAq/IaaoQKFGdm2TCJd/vtIyaOH+nShu+ImyiqXZtxAExLZS15/Ps
Yz3GArOU9fv2j3Ojk4tUp+SOEcJXMxQgM2S+EnXxL4GG97kqxxb2wqqECvIUwH+K
y/DsKZq2jRgxNRXXFlz0zd9ZJ+N5yhY3T3uW0+f+UHm+rNCwDMkBceQQM7YYxUJX
suVKwLSRqqNp/obqTyWvPZL6ML9Gg/2JnQbRTTwNBce3IEgIDsBV8e8Dfoo6/QES
tkIB1j7bRAU/QpgPf9jxnVI+5qoTBJ7BBx5coGQ8N3hCJuAQsWQYYbP05fFbrP/c
xFKoSfef00HQTvqec6duQr0KRvawmZILH4Jer0gjv0c2PkNPKWwhH/xeT/mGAWOz
sestofF9yP1XallXfG4fQR+q9zva04ylp690dVUau1l4hqaCW/Lz1RMolgGJSqFa
jV1wL4CT/5O4SC3KB42VG5dr0kUyeg33nJUX1LD7KYWzoKF+QBH8XpvmL0NOCEBy
Eq/fui8cyb7vioAfV7whxoJlwxpAzexu9kIlvVJ31CTwGurz199MjDCKZS4B5ElW
3TBnp2s/tdBlopoVLDJALLswqaNjD3TfIdflbgfPCKnud3tfKT+FuR6xT1ZrkuMG
uxQSxudY7sdMWXIOorkZYTRKTkt68QQtv9JxYHATl4bzrNeqIOYAA2S5xPsTmwYs
o+EflIQeP071JD7VQABIVCSAiuVRg8LC7bBlUdsGD1YiIDmQ/k+IUII9aANn5Lv/
6H0/5buhHweucwP0WuwhaJTdt87p3MEc21wcjtdJO0w6qsgtoiKR7rnYEEnLU0Hr
LEhadJRIMfZLhImpC33un+GFDbrPoqfztuM0dlvYSJnD9nOHWdhM68rXxO+DZncU
mlj/WXUSq8jUOGx4opPy+h6adtiKYAYcuGCg36I9dozP9zgx0iP7HgmaH5HFH2lD
RNznbgcXkIZ6E4fhF+IRCWbTvMD46MqzgzFnpLyQ03y+aUlvFj0F5Sfqw07a+kN+
YIhrff+WtcSC8NtQ8RitTI1OL/pjGs3wwUoEqsn5UOFC2e39y2ubKXxg9zdJzsfY
2ctG21Jvs0U2F4dVOJcngB358iuVKbG9niQlWdCZU7gRtFEPtUQhvqLX94Wj2+/O
3b4oxmRM4mhT9CKXSzLcJ2l0kuJME7s3xePc2FcwDdCkvH9Hybc2ku7ObNb0nSh1
Z+wh/xNOwsm/cJHvJNUXnqZtIDOF0BqrpVbBrA9oDIKGbdUSD2kXhIEQGLWSok6O
i8l6pys4UCn6dqcwANSosKul48wz0NEjp9sFaWP//50Jy+zfRvYqEyojwIHO8xDa
5Xbv6Fr6z8hz+F54UPhIszGgpC3/L+R8ZIRL/A8mMH24TtcrsHbxuKWh+PYpqZHZ
+bijcbOL+vQ9Ruftk8fj7K3H5Y5JK8u0k8bVW2pGVSLhfGmQaTpNS0Krsg5e3OMZ
LBvBJPWQnaHZQJz5R1ULmXWBXf/wj0414wxFgrsGLsKSCmlgGXGNiSPD3d3BpUmw
OzBv5sBAYR5rdwhgF2tYfokkKkW8m9rlFY9nyDrsRrdBwHCvRE9hgmggcvzhl2tU
DHhPpZsc5569+3QauTQrSIT6/+T6grxYN9uFOOUgV+A8yqOWfwNEmRmq9zDuVMVR
O5RM1GETMXyPHwg1f6ORtV8yXEO1k60ZT8EAx1424CBtm2Mwo/F541wNjUqgP+NS
9zMcoPq8w1oVr7ZXqn223b4QK0H3xoqtf/ok353YVj7MDaFdKrWuo1sKPV8uGH7L
3Gty2+cyccKqB9f1yVReZxuKnoeBsKVXNopn2CaPmkh/ySKHewNREFyy4MXOinqb
FpKSsMLxMK19QssBYOiaVIAcTrJyouKJPIkkfId3ffLxKlfxJCINx1BHM80kv+OP
jBfzUbt7tK45Y/7t1HHU+XBhMydaRUV8ajBn/lVn8XLsFMVneVS0pT/9n2AZdLi9
Dq9R8GdONNjTSJpB9l/lv9uLHIfQ+kxuQms4mIMK/qy53DAqBgAkiCuJLJFMqplD
savneQnfDbEg5Dc/saJhOBiIIb2CcGG2dcVdZdXbjTzqp/R9LIz1VCxfsF6t9rya
AghXmTnOhO0k4NeS2biJuiqqbuLU2aTJpkqKD6AalVVioKWTAK76umT/3+Ly3AhK
SX6Oj8izUaWpEKuDpdtratS1KDLKPcNBQ39GyZJe2yKLx1gERzgdLfr2hvuepvnT
Zk5RCoW6CTlXkyZI9zQ601HpzD98T+yz5xhK4IiQHQUp3hMCUBrvqGFiuSAKwSP+
ZpUomhgn7TWlq/FwdqAc2rQ2DaxHjLu8kv9ecplpytD7rc26byym0y/jeddFgzke
x85hmn7gBg+guOxC3HcSqtu9i9LEgG56DYMCurHKrQizM9Y91NQ2NykcAYLLG8Y+
kD1B+Gc8YFPT5Ax6LA5hyFxHWuGrqeHq8xAg9un6//B5NOauZ3NLLYoyqKqUQ9xA
fiuucHEF7CZc/sWVkTXbUisV3VPvnzRdQOcKuSD7nfiwFUrCj789fAYKB637nRe3
cD+wQYIopGj6Jygf10Arte7fjVPkDE7KBkQ2s0gxsAwmox/knTr8+782ZfoYcXsG
74JN2v3dIIvkaPuTPEBSib/f1cJiUg/kjIS0cHyoRFdazTaIywk+40yjl+jSH9Gr
JyW5QMbwe3OzhcuLDQl6OHY7KTUl99Kr2xZPUrdzBDP+vUUltobK0DvEK5cnzvLH
P/L0Dk5sNB4ndLrmvnET3UFejih0hnKUcBxM844Zbo3m9tN/EiTZtNoNg+YzpV48
H1nv77i6nFxcE3nyS6tsiEiuUcHZzuGBS+UXB8bI3hlQYEHCo9A7ZRx3XEAW8F6o
F+glBbutC5N/VUhWjfMaYchlTHxI4hewET/rR4jWsYuLql1oDKvraGQP2RCS3ljd
FKfRzqoaP7nMvoWb2iT5+pyZvoYAk8J45fS19mTTCLTn14RDn9HUnzZ6pFKr1G/0
IpxaH0Z7K3xA1SvrTpICXScgCeQycOuZhkQS2m6F60TCD1xP5b8uV0cCRwXD8F3D
HPwRSX/jqjuGBoOgMW++8wMffpLCOZ/S07ejnWsigmc1kLt0qKqtRXBL2tbQ3s1Y
+uIZVt9G1tgfWqJ+i+PbpLcEKidMsIG6zixQ1pMlFkwvuIfPmMpxibcXMxC7eKrq
1arhANkEFXKUsgaba8iuIddgyIQIPne8lOxHCgLrQWDKXGJvq5n8zLgq66bj+tIf
DvhU9nFh4o1deVkPzjT5Y2NMMPVGGt/ysMXdlYQqFQIf+ktc00cb5tAN/zkidaL7
okqsmuEGpUujo4qe2oAQwqFcAWd/+G4Rg6LN0nvslN8/Nc/dajBE7r+frs1dQUmO
OWPzJNNwWGkQTRjWTAH4kuPE0n2R8lb6Tx6bL4iBkg3+xUtKtRVT0dx0dCSyxIG9
rARF1gNdgs7GpGY/L+D8iNB9w/uGVzfniv0lzt9YwTKExN3Hiajpj583/WN3dHMW
F0taINFCXZtOggLl2VuVZFSlflphwkpUE27wMXrM9IfxVxpGEg3c2cyW3etsk0dS
oQe0DLjfhHLXfYwRpmAobZn5p2kgXwx79TIAci8auwiWjWhNJz0M0nrbW4X8QOtm
zWGkjhdSNDHtg9vurSCV4LRMZjbpVlo3llHUMQVcPLTVKFeCk1yg70LbZsTihCvO
9m/ocs+gCM6TJV73JKHNwCCdKHXL/PXD/RZ0oGj4kwxNGMAcTDtq4+q6OhtBd31Z
qpagZ/uxQQcj/cnqyEjb3oh30CBRU17WYhiCBjY6cUCYhXNz/k4Z8jo2fdNY8KEv
rNfR82kmiCEl+5+Q27fM+FH0P+NdDrr0Zmu0tZzRlYYyaJ/V8wktd8wnMmVqSDoo
IPGkGr174B+jFz1H79Zb0OqyBqC3yuTUVG0jY1v5AKy+tVjyujbNEK9wDYZF3iwK
3v978wHwqcFBQEy/2bFuHRPDIIpc7W5dFJwIcts9ybrRZGtWahR2JPh6upocT6Lu
Q6jz6ajW74PDRlTO54wPnE7jbjTyl0sK7JwHMnKnYkj+uWDd0qcRxagLfQ2OF43d
C6LuCeFAVsr7FgxJkwSZsbzy+Q4Y4grqN7qXI7ecMY9Z8zgiJRAP6sECRpg5QnbQ
LFh5xBAYTRRao7RkdekniiS2jDMJd5Bi0ckpycB4NR8gEXH5ovTHKOp0rnXgKip3
NQgdXdQYa3ImA3wBrhO0jeqmD7fcdHqGXLryCuQhuJ5bWV/gxmQVkXkO2clQVmE1
ZqNCdHUFpfdBHCRxNoCuFpUj9D/VsCZc3IF4mpQZDULrt6pvYPyzi2W7V8zP+cJw
HBMGJiG3iNxYwQm+UrvhwRLluU/SAJjWC+iFOson035qmj/suZb16Yur/cHQhlBR
bSJcydS0CYWz33pbYHk+KKHMizBT27V6nX8aujroyDDGnpxBBuVQtDzY1xJ4eRTD
gl4uB8SZXKiJh0jmYinXsRThE0Nb36LroxVbSoId5EfIEeVlrsWjvSXSLKIRSFZA
lPZwzbosnAZUiq8pFgl8o3S9Wmq7RzyR00ANhACQFTayaSs5ELKqbB1DzPtnfFpZ
17pAVGBU7nbLDlbGiUA24K6DVI47F/grBsnyudCq7sIkgTxni/AcA1fY9T9v5mwT
VhwtVKtU914bMigvfyVAw4bNQT8OvqnX9SPFoe2JJutKavKXzwiw1URVEAZun26U
I8TUgPA5OMJmbFuh2QsYGRO2CS4dma2bCqSUHkHsiNPCFzCZg90pOUL6YE5nv2lc
R+JBuWWHpkcRoLcZwVbl6skGWiUGbZ1an2oFGtxFUu6Ha07g+57yf3eBxQ79Up4i
n9r/jkNmeRUD7J9R81jAvifxRb6xAawrgpX+xz//OXfH+hDl8/53o0/AyMbWv4HO
HZCrxNxELjm1fvPnaYCGCyTMYMszihi5kV/b1xyy2azELxhUFSF6uKGx5BFEnKT+
6PSQ9lA2Vk2HL2QZjDLd0gW4WKkPVYsj/JGPDQwSSrmrgg87j2p3MADbQ1Yv3Mej
Ruie+/oz6qGuDfbFuhhoZmm4ZZEyPdVXJMOMyNYDT2z1m9rwmQVgEzX60UfEwMoK
TfQiGXpwLhrEWzl9RZHt8nm2FDYX9luuvGdWdrp2enS7HEO68cqx0AldAXBxT+/B
lHx4TzcsqDexq4i7qR6POTv84N9oThZLrvdhZq42G8kGsB2xRLbbZIGkHQ1gK3SG
tmyyuBH46YZXAIJSrrBp8Tw16cC4TtqyrhCJRrOViZYFXPfwdAVRLNTBoNL2ssq8
YWqTkv5tMyi+ZBA/4pmDDqWLylPWmZGl7nHDfJFzx4Vc2cTrZdeZR0khK9vaK9yn
A3HSa2S2ZxNTYpwcLidU9vtqS+3nEwF5xpHdQ5wVsXWLGDehrGJJ7g3e+MQoJ/5o
XPCuQWcH03KXi64bX8HbtHiMb0ISJfORmJ20Ri67h1HtjbVRktJti0yLMaEewyGc
iRpsAtG3aUqm4seKWijNl+/Nr1FRkd4qGw4WfgWFQCjkjXw0StZCF8T5ka94+ZS0
oP15lchRU0aC6nbwse+XtEDEkh/Qh2j/cTN3GLWQ6zasKYk9XDagZnzgKXuXQoWN
CwonhqATtGc9XLDmqsu9/qr64FTUTk0WGsGyKggnxswrwviTOtLQbD62OP4RO9gx
WZdt2dbgdPGpfZWpMo2tOW0xskbhCYb8XGUvlYMWN6RJaUsKluonHACnIEQADagP
SyIIDqlCI0luTjv4L4wcQTE1/MtKEHcXGghuoWXlwA9PSwZBDeA1DsshlAW0xxMm
xEZ0v+2SPM1RECBbq1VBgRQDV7IUXxNyNWEbQQcDsGPhmRQ2bEnZ1OLFvdvNGDpJ
hSRsBkN4yl2LN9qPcZfJ4KbjLq40Hd4xjXXC1d1hGoe7fA3b8+8IolFDMXv/kehq
XHAYyu9EcAKZ9tJh9ESnW4i57IWKdAp4z6iBoZchSdKI4jGhB1S7cXYel0nWuuSi
f3svHeHNbpHDWyddFk+ygJ/pSNnWj+DsXN5HHeUgSCtmfUG3IbEs9Gn5Ikui3Mrx
ShbAijfpWKat90XTK+Ga559kxDfRTcU4ep/ttGwfKaJ9vaGPICnA61IXJiXRo3HF
gDVApWOiMt9kzoOgjFWozovGywRWjRtBY9YoiiGw6Ll3lieMLdyaof11gyWyxcGM
IpNSUTum36hGJiPIjxS/fjC2GzGDlXsqXJDcxiwa8q9Wn0oKRqI61f+JhlaxL+Mk
SWAh6p0V8p3pt8xXKbKC/bKz966la5UdUp8iHcBsE+iboPHotPjBoiutasa9/pnG
NTQSoam7AZZXAAYad+gdRnTthknaSjzids436y7pepzSpybCLtR20quIdpsYVJ79
XnGioZTxYj3kR2zbibdZ9abMHUMjPrR3Fy6QXm4gl3kcx0iL943f3gwbLHX9k1fT
YTDUR3od9eQAW0TcG6R5udmnsS3aB5vPA1jkTHkS7WaW7ycu75WqV46yUR7XyU6p
jXqe+/7y+ADoKMB6vxVA7IRWlb0TSlKiKj/NIKG04k1jvdCfPVxLdj+d1JVWvcsS
/8GpbXgOutmwj+KOGgMFeKfWeeW32tmbdNH+m17x1Tqf39Fkb+5jY1xjkb1tYJgR
4SXFpG1kiBMwd/Nam9IXq6O3sSiUPv+cNVBqdYFajm4N4dH8CZ36CjdEl583UCFb
4Yd36BnW8dNJWRjBjAhQE3h3W3yGnNtgk/zCg8KuDp5QpC5oVvExYUhW7eeob0Kj
5csay5R5uOcVXkUFGSGeK9VNzAjlFf/1jGHzxkYJiILqhFbGe6+UQUbRx8oaNUuK
kCN7pvAVCg74YEl87NQzVkdwUlEJaLLhqQsL6D7uDNUp9m+tRgl30uDxEQi7lu3e
qi9JiJuFBheKw4vOhbtAyTHmTTfD8l+ynv4Xpj2oK97IZkdAE4WCIOxBPIK++pbi
hjgQVZjqnLjgGU2H07T/9BHGZDVleFV8udZRwQOi+W38T774Xq7Y7d2BllySAVPp
BLK2soPIVl5C1f2l94q8wPDiGrAc2tYy8YoCL4AwTtlzhG1iI/xUKSkcMp0Dtf47
6WTw4nmkfCYf588Gp+2d7vWjFkBk+xxThc2vk9hjX7OUfmcUvFkxsuzIWiYDBvD6
uCEjAAoG0w+Ox35+Sjq13QuFIQ12S867mWAhNZiopumCe6W9e0sjPFFRbXU02GBv
BdSl/iUQlttTTQ7vaUSid05sUkhnKuQhTwF+5OanHK3DJJrbRWZFs/1mY2RZ5VsB
5z6KhJq4AtA/93phIB50+dNthkXmHIezo4fgoed8cs/KQUM29hXr77p1CuasMcxb
+9ZCd3EGiNojebTC/VcNpJ/CMi7lS3ciarsfYO+OZzZCGdRF8W7k4aTc2NRXbe4h
WB8esC9dJpiMZgtffwQrh4A96sNxZhx6Sgk1VixUamJsMP4BhtE99rewW+WuknL6
3rlxHlcbNKzAXdzpGD2s2ZFusl6VSvH5DnM35H7ZxX7yRVpiZaBoG9i7tSbWCHnw
794FIzOzLF7vBiuZkAxT3RP0DmZCyVDmHK9Iu8iX5DUixIXmpkmoBL1KjnmgVLK1
U3GTiYS0bqms7LWGMzlFT/pn335tYQqCgTCHWHVQ5q3HJEDtzuPNxjylmG2ZfKLR
kvVypoqWmHV8SDAYpapXtZrW5RAxMwrEtgj6MUYh9MPT3G+nqKsjpp3n9/Pfa3qT
V5FA5S0T93X2oDoj8bsZTMf7UJx1PmldHT2XwPRbRAVuT4Km8R8HXQXSOth5WJuA
P8XEyClikud9bSTSb5k9FSrvqqBvnrkVJI6w/kmtcIirVV3F5vumvq27SS2I/HpP
qAP1BajgfIKOGtrZ+c5wyaD+IIb/+dLBTTxsfQgTmonQlUzrr9yVnMDPRC1L1p4U
+FIu2c5mZE/OXCxVpGBFow7XN3BQ2ts3IoXIAU2t2rTKczOfNp53khLRRoCh7E/A
1/CMVLcYnSWYifdoMSZH1XwjzamWRLgnM5YFNwLqsTkqA0knnMt/K85KOYPu+RI1
BxPJoin18Yr0MaHGQWWVW/QThumqzB2v/B1JQ9RhCSbrscigjpfUmSsRe+Lwok4T
hN/dt0JHuRwzaiGrjKmzJJAzU+aFPygH7HkR6IV7pOtR8+4H0I7tmGcSk+v0KqN0
SCu/6kosy31RKhKmI5oTuAnzBIUZvGoFNxBGqKkUJkKFIabuOVXgWmBnhmFpfh02
5WZhzxVFpJZ+lNO3kSx/4fodLw0ckUEaJKxNX8gC6zEgPf6IE0forCskdWP9KL3X
+f/WXLTxJCKY5dfY5+HUZBPO3ajzNZj156t2VUayz4Mrnp57D4wYf7B4iga7sBM7
dWpgTAbkQKlYsKBLOixEBVCBW5mb0IG45yxPRgN2vG41luNwspUr6fLf8Dql/fdV
vklbY3yab0BpL2chBEhaNvXUZia6mbrjYglk4jpQWP15qI+WdUbA1vQeqv71iOKa
Bz2Fa8OrdmKUzc0ZVV0RhzBGdRaB3EGNas7UTHEdzG+Jvupm3lkAcCzUAD0/qpg4
ChcWt4pcDTSx8hMC34ZkU+ZU7P3HwMfXwpzFOUoj1A/kpcJRL9y3V9Nrm3rbiSjX
U3ow4kmQTCrVYAFPrHiojxoEf0uYf54+jtuw8155I+5qSi6E36Lv9K5i7xGiThmg
KYBBXFHqvemC+Jkp39jwVer1Ge3GQPgzgm5SaWV5ASV7eARWbHelvWSsN2ebV/fM
1NzWNvs2t24xfvuJ76gwP0lgxi2ASYITenFPdQ6IFA6+NmwIi2nlo84FeXAgbXM4
efCKqUcd1pNzCB9cNmQhnLNSb/MxSXLWmT9UkVxrdmvwbHy31LGnws4S8YBxFZtc
oAO5n/RQsYAYocaptKZOWjiDZBZoTkL5nzAeRZXgiDh7FfeKY99E6+Nz0T3yxaKZ
flgtjEh5wbHObLI739ymD2jtR/KvxnKHrodEiM4o30TfdQZTNWYOm0/8JWJuT/UE
lpRzMHhEvc0iqwlyxGDee2BegRt/FrVuPw7PEu4Hq0ty//TjlnBjCJSqAEA57PZH
KweqtTbWWb/fOCKhnLXNpUpqYdYiwvE5YU5bVTPntjrMi/faTc8UlJrnSt1WHQFF
JBoJWw+O0VOY7537XQf+STjJcSuDF+m80DHQD/ysRGDXAm22TCx7uIdJMO8riclp
80k4Njg6+fGPzKxM6Kep0jxBbOv/lJ2Rh3K3FSYQN4OIqyTE9m7wD+Z0HtkrvoFB
xhq3v3Azogo8T+pvTRzCzgYUyivNeyKdnI1OiMzThjibLaVZ8IVOfLsomm+zfmTm
W4D2knDQb9/5dfH7dUsmtbvPVg1U1CcTJxIw+LSw2AYXYy1xOfgwx7I932g345pR
67zvwm8Fi+07d4/NO8IcdTRaZvuK04t4bmNJ9E2guwTEQ+FcPdktDObKWRM+/HZS
pSWxoRhi0wj38L7ysgPOgsAKC+ZJ0od8kgo/u964Hky6lyRXpHfb5tRUO7OVq1cE
Be3gGOvjBghZOWoqcdRWXjR4dWFJwzaBY5EqET1gVbCRYn1l1MY/2umcHEzBwhyJ
CM7dPW5+IEnaA6m9t7xXRwOkScNp8D1kpnX8/0I64VjaeKo/Is3Oq7MFAMuibfgb
Rt9828kuDPl4I6C9kg5TDVT3AR3GSO9R8adC8rawk+AvsUi29yQoCZMMynaMQKzB
IbNlX4VNjhSlWPWcUu/gpTHPADdkeXMkQLXW6QCZPfXuNpJ5A8gpCVHeZRUKscp4
rbU+Und4cnDVizwuyDVPm4hrILfrHkDBC7MistInEjstUKSWfM2wxl45ZSaI7h+F
4dA/eVkRxYEq8ccLfEFXkKkh/WjxydnuhVjLBPUuSBO3mkIKFRc7m1lmJXIcGn+M
U1ajUVvDiB1PQdDhN6OEjQW1RtfCduAXAlOwCGdnbi6s9b5s+mCazdtCglaUHXob
0pI/oOkaWzSf2OeqFggYOQvQcczKkvAOoyfovhAGV4P6TbVYwoSoyTsG+4nViZfy
X7sRRytO6iiT+LyjeP/nbeT5LJ+qwDoleNTbkq7YhoQiZzRhqkgv2CvP53EJk74W
I1kh+TIdtjwg3yvjH8afqUsy0j4H2GjY2SWZFzfcduz1VIBtf5GTukOmewLnsqw3
2nBl76eYsJpqR7RserEWzb6/ZEz787Yweh7GHefW/q5lYIE6AVeOUxyqOs1YYKSM
uwPXkyqrtqS0Zzt8yFrUvuy8MDOejpVSS85fL+sM5MaW/ih7I9PjYqx2N4r7qgld
DSJVTGUnTbi5Bx4qiq3dd3RM7YHo6jDBPR8tJUHa1BehlUsBVF77O98mabl3qHTM
Erb6jI1Kgxlo4Z92nf8fWZyeVUHtcGrOuN9hc1Mt3CI9Kg4xVCbnqlLTk6lVlOuG
yb/Mmq1gmbz2GCAf3IDXSGOD5vFtK163C6N8CyLSzIRLS6TJYmlq+H5/L+QuQNEr
IV1ghPwyE7F6vykFmI02A6we0wGv0PDl8ltTy7N/bJxq5rY+yaVZzc8YbEchmv12
rZgZ+ldYt09aF+gcL/+5usXHCJVCmY+e6UalZTCTHRKsyRUfjQi2gdSta8/MNput
ZNsbvb0fCi1H668jGwgmOq3AuI8NdElBTyjTn39jz7TFUaRZp2dLZ/51unnWj/Te
F1aCMFBo8wcSWhgn73P/GHMiKrFcn37fZP/VtsdLRHver9sEdyjRgJetbLK+dgQw
LUds2PEgVIS3ZZlFscDBU9hklIonCKWnyeBBZh1Y8BVYJu0qt2jSknP+dIUOC2mJ
vl61LDre70aKQlNIarwIQNNZ1wk8m5BgOriQ6oxL9YmS0by1Zpt5ILsEuTcnfo5L
4T5C07oixML55rorOIZ1Gs71a+bnJaMfFFG4sd+R9e9D+yxNHgtX+bKvDix4wfGV
+ktQX3M8PV2ZL9zoN2D644eiAKd/bw97HooNApuZBoUN4uJcIpLyp8fgT9bKdbdT
3cxdRAer55685rH04WBe0Rany0n3+1bQUx880hTXweHKqBNORJgxTdxcFvKQPuoC
rlDSR6CAAk+XeHyx8tHxghJ4vtiDAKkGArIuUKEBol/xb6/q9yICFy7tN0RR7WnO
0+gOdCvKLbFqM78fkVjS+1OjRlP8SHvqGR9Q2FvuFiKz+Bujklo6CswTmJG4C3V4
SiQ0OQattiWSqcJs2LUEd7gHncQ8EoyB1v9NrtOaVBLnAJc0+sUM2MdO+dzt9Uys
nMxjpA6W7kFYqim2608fbNfoIY6a42oqAfDEwVH8WfRQNRRV7t3id/GyotmqZ/oF
/sdAodoTBkAIo0aF3CbDn/bwH+uwBQAnBu1RdhIAnuwgD1wwk9qYHkM8seaC+6hG
8JDEvJo5G28Xrq3fPi8skBWDQeoaCS+2i/vWfsUimQ1TY/nV+XNxbKAZFq72iDDM
6PDYx0ovA33Tjtl2NAlkyGIjp2EshC/2YEYhAllskMo4Dlg09U9Ns32ncDxDcJrh
ipWG6+SvAkCA7U2ZgR59L1/2fH9Q+qnDL6lj32/M2BchUkI1FakYijwbVc8JoA3G
9G331+PGl+dBNIYGZJLZH4f94t2t6HrwjJhNVsEEhH79JiFiGY8MkCbNhVfqHNE3
Tw1L3MnGuDE73jo3c1xaTh93ZHzKEOGvVC+1SaWKrNuwp1Uz+jDjRfV8Ga2fs1Ur
qq5iS8cvYUox4NX+Esz7/Zp8YusvRscewgiy64eTiwdTJEDZKsJ01jNpBiXCII/n
UYDd0VBbgK0VauPzLDxksGPpGFtMl/q2P/DoWd4NHueUb33ozi/P4vtWCWevROFj
9rxjPKdnTm4M7tJvhvbibi3ADlBjCoNDeJzmZPsYJg4ms4Dx6rN+4DXJQbEQ3W9Q
wwyChH3N2melbYsO27vJb5/lCDZtdtNbemeO9UvlXT2heQ4tAf0mLjo7xsPJ7i8L
wTh/CLbr4mTQEC8au7kugrxoohr4Apun01mFbPiwG8tfRzO3HnOrspaaVqzNn+x5
wOD9Lx+S6+BEHJ8wPrpHoKonLTdohQiYJZI+VJCNzRC96KIXe16iWXGhI6fI3Olp
c2Hquo9U/ooHse5+XbWsXcSuOJQBXPnnd/SJqtp5X93leXtJnsZSug9Vh5eDuTYN
Fd/SfHzz92fIAp06Ax+GPaH4pJ4EPA5j8fFY0NngIVWFQsThtxe+jgyVxCgJvnXA
27O1efAx3/eXmAjSVCFi8p26uXyeETMsE7yF7pBjrtS7px7wtYrBWuOJCj+VuS5A
Awgn4W9ApN5z86vlJmHMsn2Xp+m88h/d94IaN5X4zK12fmWo9Y/JsrTHQPLAnGms
Sn7OH42WZr4PiFOv498Febx44+isY8JmnNuoXpXsNHHowr0i+49LTrSi1ApkX5ra
BBQ/FtUluMbxhbiZhQm8FxJc4jrUiWVyXcVNyQc+x0DZNP/+1Zlb4GpgpQDMBhU7
lEjocRRTWvEopvkdVujSrXtjyH7FaiLnZFTx8uaAJYSkXKc001uau4UiudQ3cWgw
wkzseNKN6OH+3481xsSYSpAG8s4BMnEVRgXvH89rVl2qBtNgqipeCTJFdm6P8Plg
jO5btra8GdXhQj9/NE/2w04K3kEr/HPyFzzsRti+EmCRvqjIaZj2BXBb4F2LW9aN
E4Siu/4Sb9rBEgRf87DodkkS/7dtp1CLKVlPOuRxcRfJwM1T3y2NxBFcgDKDGZSY
oGZLu4lb5an9U1pOn5/E0T9+jrxblm2H6GORatO0PZKfrrNYPLZ5ceDmVBz6GOsF
N8frwpzgceLGYdanNx+8ine8SU92rcbm4QpmN3nUgkoQ5BOJLKUge1u2Nc6qi760
26nFouIMGCRhfF776+8ciu+Ux6vq+x8EVUWoEtKO+BphWuMqWc6FLRan1eoylV6O
O4SKda4KEbSdICGnZhLvtHOLx3tw3SSrE7KjsiRaFJXjtdQ/Lkxyv1z4RiDxH6Qt
EwdDMc8md3/wXNHPcYEbbk/fO8SiJAFUVpmuHfgYpfEnAJ7gthsgnv6dFYD/ovKW
2X44jO2kJiNQ8RgDogzXjoCw+rqYu/3Ms776DP9QKNEVpcObBneru2mHiDEs+LzI
JieIVG0neM9ALuh5EEPrpk+ypyWkfm7Q4pLGyGdL5OSpzEl6OozUsZsvO4FTdPvJ
ZPaEV9dXxC+y5qXgssKTTzTIYagORcbdDjJN8cedMwPMEmhs9IGqNpgSEGkhjsor
YPPbNZ6eLJhR9wJWeh1xfsv8t159UKwHg43jcpryspcjR/IMf6kFG5GZUxhUMUyF
KptQpMoXLjB5+naVzBcOjjXU3JtttE5zYkE0eUwSzIcY9iOyMl5PwFNWHanibrY1
o2jPwMdcfdCIn8PlyxdffgUGO3IAPREk98t9T26bJcu9m9GQlzroKocfx4tm2+9v
BnU5xw8vx56eGMF4+COra3TP6Ha6XR6QjYpWFInOGH/2L4OOiaYVhyqqrK0DC+QF
nURKgEK3xyFuB0oP2fu+ttJNJnvysCKQyPJfr4SqGPgCgehGDgMCi/Uh8dQG7sij
df1cSdM+VpzXAlkkvSOeJkVqFXjiLhG9qLSH0vEZuVEYVzvQTQYCqfdAwdNDUmF4
UbCpMbejLUcbvEgz9yQjtCiE9VspwxpkEdncTM/r7dkBVRnrMfzF4RlI59peJQrd
l0lZlmvjYcmjFl+nIgjlsU4ApTCF6xTSoRAbg58yU6J98Byc2NdK8C4QkXUfzPwu
MhDB2cCwOdTQVXHdHxxlGLdUSUjizyQ8FN5f3/SLHvQbtPNgOYbmBaCDP/C7Ax0D
N3Z7Od641dug36FL2n9t/6dFb4Nr7C1zvoqhLxRiIi/jMJFLzkCYPLjcm8Q7qE8V
GnegfK2HQjnlpKcGirSaLDy7EgpfA6cuGg5t5TaTf++uT0w7bKrDvPIiP/gWB/YH
5Xyam+ZZUA5+OYen9Na66VmDBJPpI1B0IG4H/1QaBFYTN+y+j2PAuQZjg4UnHp0R
UnHcVcLAyCTaTDchN1W54jwPQxbQy2JKQGprW7cIZUZews5HNaxMeCX5z/Z4e5cJ
7pr0xvfBnnSrRNVrnwKxOX5FfzJs2pB1J9UN5ijmdf8Unbjo2qNFHVVGpbGl5uj9
rUc40BNSjxZHp0YUrh6WApAXxeRzdmV2ZpjNhoqMliWDnXCnRyUBYH/F/N79HbFa
yx1l13nrqY1ha1Y4m9yZoqYksmiEZpwgXo/sKVtnchfHGWj9m5GMy6axHvvSnJHg
R1vbVlKv78gDy+H/4fdhrKrlZ4MwzoFoUg+liRuKJSpUIzGu35ro0shK9hKACkMs
+IshV9xyt9NsdN6DTeTmROSQ83mOmT65esa/hKzzz93xl0L0wzmX2mU4sHVKFlJC
1KbBZ3oSa7LSWjWHE7C5PFXudte5bIc+JyZ0OjeNEtF55E68hT/giGj1wXEqKYpG
jx4n6/v07r1d5AFhyIM1xCyk8jKXVto1G8qP25zWVQcJyHznflzU649qHdqYfK3i
ZqptCCpTxGKutEiC+Jlwg0LhJj494rSZdkSQuCKynuvKCmwB0v4JabmDlQhtjMQw
9StFUbi2XiidhVuTVowKkE6D2V/OKFP31RqVZlIc9pVWAr0vr6bV1oonRW2mJX8t
lgg90p/DboyzNRmyxvcFeUrf78RrwIv1p/2uefCwu4mY6uCnDfipr3NNlKHGy94V
neFOp2THff4TpjPf+fkgAp5Kg9UlcaKflxbiE32xxbXF9KVoErBPoDoQqyxRlpvS
s/YqUKZFB8/xcPdr81B52FqrM61hoRhDtasFJkRZwO7f3EtexRhild6en0cd1fPr
pQOsmJQVeGsIbb1lFELMF3nbIEVUvCfXr/5fJNcngFENCqCVAcvGlOcvHRpN/NMS
paIni8WRZoptwgjNUfq9FGDD33W8mQZq1jqxl+hTBjEZfrqjTWHeqOaSgGpEFmY1
8T8EMnj66hhRWPVJhiiNPCpt+/j/FBEqOgNn00eT538n/sDld1Jwwfac6hkCF8AN
yRTwK3FneNWu2m194kUJolDHBtxZCQXdeqKtqlwU/h121VnedFIo/TiBLA2rlkaa
q/9WBFMJvech1Zw499Ptwb3454Hvmvx0MNYlauNaotVFlhOZH9H+CSrsIuOFuM8Q
X/f54ITbQzxscWwukDfEuLIZ+j8gkiKIjvLK71oBK2rkAKu4/f+HcaD/dh0qU1eq
EHtnWDTWi7Uvbh2Nk4BcGkgsaGad0uJSlZKcmfLziZel44PI8yqspld2nImpS5gK
+0yvBBR4km6mkTLHsLI+S/49Ned0hDQQ9pz0+4HVB+NTgCEXGzaLlC3I/3n2RNY8
nyxawO3tcXhmNtME/82hlKePcp3LZP0ofqM3Pn0tD2bynH3/ow9X/pH+nEjhhoum
y2C/Qt6fDtS/IT9/8HpdVqyBTUhWKxM/Hth5iZLdlLtstw1QPz9F5+DdJOOtCF0H
T8b//37fBCCPuub0KkKW9M/zFQOf5mllIf8F39v8Tgm//zz/qapVbN1WdpQtc3d0
lcyQymiFzNUORSIex8hgkN4acpgyK90rpal3IfgRNQAS+P/sgftVyXHhsTvX0qPL
Jq4y7ZiLPwDH/dfteEJJkGPwsR58UYFbMbXaAIz0BqVC0yhbZR2SBSDhq0T/p2ap
t03TIxQKg/GUGuk/x/aQD90lLhe9bcAB6vAnZ18P4Ybfagwo/eywHKgeQM91s3Vu
3NZHrt8TlF4JRxGyJI882MRsekcnz2KkGcUVRzI4PKeeg65XSMXqXCce2LMQ5yy8
CRjsP8bJMCmLRH/NlyYa069T+gUdTIkYxBt8b8phyg1baLBA8eKMRr/NSnpz63Ta
VJ/Uhf1IjI9DZ9JRkiBxTRZ2XscWYKZEVjAQ4T7dZ8quo2YiUFHUc+0OiU39Mhpz
dMPZ8OrVwpjNoAzV+OX45+Qh6r0nucaYeQA9F4Jm8cRpE2rg8rPShOfA5UYokdkf
hZ8j6fmEspPlhI2d73EZVyQPWIfUqU8vsz59GWlYMZxNuR8t6b7wC1UGvdk5nULD
dj1atJCQzyuYICE4oeINkZGSwW8uRm8cC8JUSoaQnJaeAO76RDBFYYoB8/klngkt
2GCWcO6f/1DvgF7u5E+FPWsa078O+Ufi3QSsWrYj06GDN/3yHkEw+CDZwWDqDxTe
iLyZnav2R9J35SBWaMaYgDlTL6YxlwUtYD3Bbgv6/vEKmOlZMF1oPbHWAtVmFu1/
6hdVAzheZiJ82PoaGhrtVb0snaaXEKeXOphkiZvAtxxlzKd2ZRCA6Xkw7VxEIljI
o0UOcERhYI3RXCjCHyoEDgzDrSEMf49SuDd269c+19H7lmzNvZNYE0djIDfHhoPj
AsYZ4c1Fjbf/BFxtv3ChA5A1dABVtok3upGJEPSmp4DGjBx7RuezieFssDc1aF55
cMbF7hyiFhKvCPUu6EZRn8kcSFv6zXoCEOvzajV6JVrQohWJn6JxkCZbEIegPneb
r72BFRudXmS4Z7iJx6HmD3MzM1feXzXqjDxvzJqIKxaLtWdTEVHU+AsLLcC6bLJU
eVNcrb5/KM+liYYEIL1Z3XTqdSsipW/FtrxeQFIVrcBIQ4ng3a7PIwgPCkBEP2DI
0DFCI2OmP4lWviYK4z6bWe7HMBOBmuvSp6QX3u+cSKApCnNpU6VsWtWqZuRD+D92
Wa4ZPbIQRXJAa1eHn8LsJq6M/Q+UDqjHMNrz5SfMc9eyqnJ6PQcRtJ+MUcdozgeG
JwL7/ujUv/xTfnGVzhC2dmLlWOEOi6q5M/+4JFsPwn2NecPkoYSfSWkj9cHjDEoO
r1DHIsZ5Ul3t2FMIqBsJDVjEsnmGFxAq5PwFXBiscvCJYDiK/Oq6zp3W9jcUjF8J
exeDbYseDEWJT7KpuRA3O4mU2Th//RDHTLgi7hR7FDDxVJbQ5C146mvHza0mZZXB
36VKLvNxG1kli9M72bLn7yHrOokm93IxJhhuIXpFLEr9lGgu29JpjXf+XHajoGWd
S4a5dEzFgbeWBzlO588UK7R/E/jN6CnKDGQ901dBQzzqekDbtKRkdFTdsIolrtgQ
LY3zxsr5ozlYn4guTONOBQe8h4hA7TnGzCJp0L4heYyV8ZEHXfxq6RrbPYbmPMK9
DxbxaZ+uY6uBK6gcFFuy9e1hye4uiQkRH7gsZf5mOvxkdLSZHq+XFPEQdOQj69fJ
M19kNnrOZ9h6Au29zEaAO/pA/QUoPcuAUJOT4qBAkozWP8K6uzuGQazp3ROIvrf4
Zbp69FR++7Kze1h04QUYrFDEuQvG5EDLLb1OqI7MTpnWevIEvN+NAN9SUS6M6vU1
n1NTPJZc5Kp6JXOaj9uDPGAgcT81vxy1dvX6GsfY+RWThwLzM2wAlnNwWpI+g8tV
NrKpW80hBH2LFM5o2eccRM8PhbFD4X5zDy9a37KdpTgzUSOsCvDya7vNnHbOp4PK
rX2vGNNxsoclPBpTf5FiFKnCf70McI5N5Rvjx0TkLeUEfHNilT7M0Matfr4fs7fw
U12DB0d5p5nf+tS0zGMlDdanIbcb34hcGHQC7YteqdZAOOqjOUmx9hjx1+oFZRF6
fMADovYvwnck4uVAom3klTR94cWn2HVzBiRDhU2MYlxt/q+i789pkCDqwyWnw90W
092QaedcxG0r97nZ6Xjmq2polos3jr9arZGYiOJbxlHVTOLGWbygAl2sglOb7BwC
3TSsp46N0+xDjlI2KunJpLbTmXz4Rys8EHP7hVfvsVUk2KQKkpsv/TutjMimruo8
xniE0D9yNX7U/QNham3cNi3wlvHvi03xbj8HdBD9rKEqYGWJHEvewkgqh32UCwGn
W5CFrmptRWzR+IVfw5O0nHQmxcN0PZizE0J2TNbCSY5XIxeGeU7Rm5iHeLKZj/ry
o0oB0uDfuNnoiPQAMpu85iqjs29PbBUAsbmThdVU66CGUDEKGsgIUxJ4DTrkB9Bc
GDj5I/oZDTfMjnN49kn+wC6NMRRtmrnzDfkDVgIwO4EztLmFAT6xB31qMWdzSvCH
1LLEuy/g2btDjao1SR9yf/+ChBZaTnynMv9152NvVyZHkLYtqAK7HqSpK683aDUx
YQnJdgE2gKdN9k62ziInzu3V7N6i7AlsgF16wJEjV3J9hHrn4iQmMIZ7ksbmfNAa
q/7c3SpCHTfUkjeeCaW22bw8RjbQvbsbq9DFkER2Q9n4ozZFlqPCUfsDzrpJnAJF
m+5VEgx4KvpfY6anUqxTwR9Y+uSaspHgh7uOtffczDg5IsXP/8cQuZz4J73gJM/T
EgLI9B4ZPrdeqxCU3dx2DmKyHSHaqXsLt3dVG0TCsc1YSffTkR9+g/npz3JeiacK
+YqjKnb7d6iPZCK+ZkeZJqLDyM7QGk1k8yIirarHUATQ1V5yac1+1ox48QiC1tm0
251CdU4kXytHOSKARpISJGOHNdWVvpyN9tBPhEnywPHxFiwcbkmLjRz6pZpjGwJD
lOBdf06EYPzva2NvpTa+vNuK4e+/lMNlmCa1AkgS4WLwk4bbYNLpPNwfpLw8CGMB
i0J3eemaq+pGa/QutGFNI/sh4Z6SgKArVjKultI5UwI72L7yVfS7Ez2dzR7K68CU
VuobIRG21YFl5HVAM8enfnn32Clxaoo4FdFEaC8LDmNmLj1U/UEuLP7w2+bLyVSB
ykCz+EpAYoasuCXRmQuX9ysc9Xt7mwxBOxH7YRWi7oGWuYpGrm1TG3NAIS8Sru8q
A3o+giEpUQs+zYpoWheOBGxz/uedWv00Lsb0ByooqVXSJvuvan1EbBVWKsPf2zwK
TxDUj3IACyrSHl5dQtrMB15xxgTe6C23/5znM6p18AyNWYm8wnQSRTrH9EjbY6Ld
6Ei0p7Y3JRL/rZy+dCJkVDpeWgZBBFm9kzuUVYvqps4WBV09F4DCePzZgohP9iak
YAh1cnEjV75V3QkLsWDNZb/fvLb9JcCRFTDjS9x1y9OA5vUkIc6b85Nf4DYWGNlC
vWRMxasADuAv4MTDHEFDV0Wels8g+h1TT6a0tdNRQQZguVT1VHaw8ZMWhMHcfLLP
zO426zNZC/qIyJXu1Yl/6nUeNuUBzZB7gWaYayZldhluEoMg5EmXRE8R/2SKSCN5
LazT4Ybi+L4G1/l1gEpmJ0rqpfLJ2Ap0RsmGwzB/iwhW+a4s3s1M9m2b6a4K6rLr
Oz66fzSf9rzXGXTcbER9m3S1BgDgg2e7usejmzxA8GP0JXIVZ5YmvtfJUvei84mI
Y0pxyMGQn45XnQAMDMngI3E/6Dh0mnnMcpKT75uDINojJ6Xbl5nU5TAN1fOm0Fhw
Es1k/2ApKwrz7j/80JPb6zSARgB2bugc7Dedj2bZHg0Ia7Z0s+v6+RsWh5sy+kXl
ec1Nmex3RdGbPpP4wdfQ/N76LvT/QE35cULF4B+K9Ejn7aeC34Nl9wzifIhxgiNt
+mGOA623b2pyGSZQaSNnDwEY5459jGbjC3TZYed2X4RlEr7cae0CXu1UyMaEGwn5
iZLk9UG+7buglCE4itr+eT0UALU34KgmKn6CoaZRfpP/EDsMFww4g6T65dzybTGA
2jSbmmKSqPxusRRDCVJ+gOcRbzfTJnPIA3IlY9GakSstKiJiYQ8dmVdPiq50kYXI
H9tjp+ShvzwbwdLydJN52IOVKvQFEMZ0D8MrYAZ9GP+BxkyezfMX1TI5cqmGL3gE
cBu6XivPbOKLp8kHmolRswm5OgBtpfRMIoZvkS6CLGS498YLN6JNLbM3XhnPGN2p
SiDWeNv0Q95eT8QVtucjYeLU4/utSzXQwnhnjvM17FVbaZEPls6GLtsRy1Lkru3t
NtBlDu4jQuhAu5roJGcPqhnS2IDDr6V68RoAwHcVfNDbjqb1H+pPwPD1rwOYg50K
ciQn02QEpmfFLVNiSjkDetCIXfAbfQI1hRX+TICLL7D5nCaciIPfEgmpjTmEMR8A
S2zU+zdTn0TlrU2KdLs3ycGgxnZ7Y3PfKspODbGvzyjU03VUzLTdUE29P9SXwLlK
b26WTFbyPk2diDx1DfGgOUaU2uvSbzx3ZPY1pyu0Ii0mckRogMUIXaPmRqmkQ+ZA
yjDxAPRlo57igB/bR9o64oCgpdX5WGpBQDDpf9vzjhzZl3k7Yyt//CKi/AGFn+kV
sHjgfmZ006Wk9Hp1AIZucW4Xtd61JNChL8woU3zHV5vlTzfECoP/MSmJLYT3PlEf
NQKZknWBkB/hrsQBE57vyXWp/RaqytM2wm/FFSy2DdJdNeifF24dxLM7YylFdBrm
H2p67FUVn3+d+n0HsWFB6g+7NxT59PCIxomycSe8Rat4ahatJTzO1YEhTC43SY4q
HVzVTGtirU3HEM8fn2Tj8MKhWHXxYEc45CzVx5SC07iguqQ7qPhJBnkggMgPFoj1
uhxdxcuGw96jSvTDAs9w1u0zAo8LwTMH/l6AhbMNpHmJcuxJXInmzK/bnR2nq+kz
tHl5iAIiHQiD3q0H/7Hpi/vdJaD3a9D62rGcvZw7Ht30MPlJVj04AzIxaSXOQaey
OVizqGX4IeL0UVbwRrdAm9veOFi3uqjTBZzJwxu69AX8FLU8TFmSWV4G91x0aJt2
KG1nY9R8u6YNxCFxtDb+wAvn8o710gi1uFXA/n00OiCP/GfKUGH7ybsm7lej2nNU
IT29yNXEJwyld/5El/BAC3HSbs53fIboFeT0O/SZz3Srfa8Fpa8q/AnGNFTdky49
og3n/9bijqrRA78rDyYUUVXARnMfzufqJwAo6veKVNkif1IxhfXaQQWeDn6Z6U8E
L1Ztmc/Xvq+VytEqbW0nPdKLsKR2+7wZLVkIGy+Df6ml1NVSJOJ3Dq8kiJP9NvL1
9HMhPSmIJuc1A7hBg1BzqiyGNJtkTekUDnTHngckBSPcueVu/rsXEfV3U4rbzJ4Z
GbB6UYIbNYU9uYH4ZvyRbH5h2q9UEve6Alng4fzqAIU9iLtnBuQfybGkk4IA7eiD
zHH5G+TfURaF4c2Fy8Mz8E0NVrBpZuF4sjAqbo5lc27vizgRhLDFCI/m9oyNltwl
JmtwvtmfPeXbTZSL55XK1MxmMLABM1sb3443njP7xpXLRgFJljpOVg3eV2l7+D2d
lUG10YhS2nUP3Sdz1lzZ0o095yaUb421P0JlUdKU6MLqfln1FL0nqsoCNE1nQoyc
kemUf8qnR0rb5J1gBdOUgNbQky6kTKpW7LweB3hzeECt8mJnGReEEtl/bq/xQLvi
NJ7bYxCGK14CLhb6a+cf0fjeZkTIPoJyBoC9zL7zXie0iQA5bOFErtAZFgSqR4F2
2rRg1/0fhzQbLIWI2MSfEClBNNEvWUMSuTq+JZzaljr+MryioXnawcoDvD4pdrZL
ZUyZ0Rxt6e7mqJy/BOvZwYkFxp9lJUIAcL4UL3dwzDNR9i+VUNHbordb3qInJfCx
3ie3+fHzBEFIdLDQG1FOPUJc0IVy/FjhZaQAyEHpAmVJWf/YGN7FxTwkCbBjDUs6
lrPleGo6ONkl/CbeWbcLD4v9gM4Rqys5WnIE6zhe6SFR5ybEg7dZw6VRl8HIvIqm
ksXxHboC5nF4/VpSgHRkWDhO2UcElgjJPL4MplJOdCvZv+tn6zL+GDmELSfiO+K7
mRDmfKLM+UBNwp0eSHgYne5V+LajS8Rx/kB84C3j8JeLhM/aAYi3KRtB6PHB0yk8
l60+gwgveVKCt9DIa+Hf+VDbGtge8j86rN4bokeAWpXaUgpzLK1cZvQEVdP6MVyx
/wzQmrqUQNSqTtD32Woyz1PRBRa/pxPy2eWG3FRLAdWufXQRwv8POLV7yI7vq5yz
Snb16LVrG3kkPgAyHygU+gBsWg29QcuOM3tCX7/H5fjlbMijuv9i25bEveZxHfY2
rV2EdeMf4m+RYcojlqigbmFHldrU1wg+9/MxVl/WZTSC0IHqOWyRHrKWKXyqqAU0
cVy7Zk7xcBZZIEMLX/H/rz/bbQhY0pJ2yvHjxojFW3bzb4MNold8dSiXbDG5qteV
RxRqjY62fxQWhwIiv7CGfaqWegc0n6JzVkVo5i9Pm+vXol0UtZ9WF3v5ipFaiy0r
nSjXvnzf7NeOb7b+knHKb75rj8XpRXHzrZ5N1GwwYmppthPifnn1QTlBBrIeC4T0
kJNK1QRRNslXz3Kn9COlvrHykbI71p80Us6BVrBiiUnlLHm3Mmg4uk6HJO9Qqfjc
UqyODWrzd4HjZK/cUDIjvv6GVJFU9818/et4VZf/k7xhxh7L1RIQVEhNG4K2kFcw
BLlMlHkOviTX3ZRdYkXC5mMOm1DwkFNch1oGXhKeXK6JO4yfOcGjxCt7UeRR1Ir/
Sy7ghktmKUqZTv1PCrztpLEZzOrr/jRqniutsmuXyrJPJ3YiPYRvgfXVXa+cGf4N
AKtLj2Q7RdAzYQb414B6uxkg3o1QMmFakqunMaI7UYlYy0gMTeLv9xR79wVZT6H+
BelM/QxpaiFeDYq8QHvlMIgDErzIMyuVzFjeTVZGoXCVjZR0bMbve9y/0lXnBpR3
CO3nlCmo6HF6RUVdCTw0MaeKGu3NjEUF+EOM9MmOf8aLm+21+vniR326AoiNHqMl
s6NgLbu/XUwjHqVl40HlqXU85ERD/u7yIyno40X9cScFigXzjwxeCIoInZX28AWA
auouxx+b5JkpZiNaPFc/QXlBimrSag3CBAm7lbuEOv3wH2jcIPjBi993rv7Rx7Vc
qCBqzuIEKouUspuF6xNbgQFWBTu2VX0sizDq63T8SYRKWW89xgxjZMnRUujQVygf
1/KrokoH72fA/BNbNgGJQAft37dNjHiV4959K3vt3UCBCPtyR290I5TI/ZMm8krI
teEKrBoDeQjTnLVePgmrZEq4Gx6Ai82wsOtNhJ2mydhsSXxvVfrvfZLNhRt7Opju
XzwQX0az8cKGu/ub4NAGkQvlsEhNFJG0ls3ha6DpAYMerS9qOXwGxWct4dwlt1VX
G6dRNq/S5OuLSNCD+IK9MM+YvsiTkWpMoQqBuJ2v5uNNDWdpZ4QsgXGwKSgdXAxl
MZ/RKZF3nBgGyZMUMn/F+5f61NfmojrcYrzn8EcKo8zSeNi04/uLiz8r7wn0WhAM
1AaYBoRlX04Em91oQRb3zikYL2NQtfLYLhXoq6t1/GhaaPlhRV5x/M+1X6j6NGOt
5Vtvz443qGGxJby7F3J4Sz2Garnups8ziHJRsP2jszoTg41GiyN95pwK0Td/84qE
Cil+CvYN12yw5a5tS4+ivxs8q0iR8WT98doQnqms24oOLJ+1VPhrSwRkOUYo3qnC
PoHz5ZtBIquB74sFYLAF/vs3VluZGMWoUTlKFrEwTV88Dn72+PjgjhhYQBzk3E8p
bZrWCrqLsD8vqyCrdEcXfquD/0gLgUYqmUkVylQ7GNLT6NvFuubdsJfzn0ussQq7
qXXOBzGi5nvvVoAjGkLDLE0pjW+oICQpt74S/BA8uG4yFT5Ty3brd/pCxyQ7ErDK
gQKdmcEfbFcIUBC0Zvl1M7oZZdV0t3kzaKK1J6SawmpteFWwzqLMmGFSBl0Ov9lb
cSMHeLP5rtwRqjOk8AIVEaaP5tfxC9KxSGk5CG6tsDmb3F8+ZCDHKkIS9BdgNbwJ
5rU4HpuFkjgb+aAl2xhmVh0QjGdLWcqGCnTKaGzDdKfZVnWDzqpGjyNYX5I4B1qP
hhhN35Ezz2aGitNTfeiT4XD2hMvPCUQ0mKTqMOKWnmz3eTHTfF31yvwBQmv2eK3b
QPXXgA48vpdahjNnIDHpKLZRBPUBwPyvNIIgwvhNPtXapEkocyoZgv9jFK+iRXIH
kHuQ3wY2/MfN3AtlM+3vB0PhsvrjTt52v4XGx05JYOTo7y2wywVBeLcgdydiXhTP
ao4Fa1IIEiIZ/gfDGPXyrR3RlHNtwoPfavv6UB99Flt6mrB8YUCi9PWXjSufKcXO
Gg/vWeF6V6VuKAMwg09VYSpGknsXuEk2RbIrjhQFfTj3/urzBgN85ZE7txv+IUME
IhqdlvQXBkD6ZRFkALIRH5/YrFyPulwK0D0eQ70g6yXaAaJ3E363s2UIUTXpwLby
I0Re3zNarBkoqkHyKxyR7P0ssDrSljJrH3Pu6E4trf6VT0VCuygYlq9NYvrAGfTb
rEWKZBNY7OHeAQm5iHfoE0rVp46NJyk5kQo5XJwzosyt5RnEj7PA777B8g90ZvUF
mDnyhOv87S+lsZJYj9U2abiMrizxj1j3OR03bpeuA3o5szUKg5Bbp0HR94vvmzRh
1Th/x+w/CvVLSG1pld7fIGMLaap87xibqbuvZbECI5tcy2c+WVM2a/F1AAJ8fGPr
0ZUXHmThVfG2DUfXan8xRD1SqB+zb66x377t8HodlG2KbN5a6puwuEbD36gXGU1o
Z/urGNEaWooV+932NfvKoiEbflG/jy2pAbOPo2o6y7CYRLxJ6EzRreUSALT1fTAS
rDWvZAO2f8zn7Jti7LdMp2NBZTQCJniSsdIY0D3KjFJGjftj6dsEzOlMF56wVLRc
in9fuKCtXsnJuYb0P0zjqVU5zE0P5wbhWr3S0swCpbUaALs3mCyZRNuB73QhW/gH
pV4y6sHjYj2Oy602oY1AUom5xM/TkgV+HNLlQimvWOiq/JtumAr6DV7N/gv3O6kW
N17TQehmp6Xxy0QoKvYW7S578oBn2f3g+kyruMxlX+h7hKQEg9liU33OvCVt2lSP
aQ/mMUTZK5wC/G/aKM7WMq0iR33SiSfVQ7dQj8Hn7/BV1rYul0gpafhvLl62MO/w
w5te7vN8cf2X3YsIvrqIBlOw3fPZvknNnY9W4gYzQ0QmVTEBFd/G56YZqm7twWP3
jA+u5yew4Hp1teW6no324tOqAJ5MrZ1/frGEKf/T3JBjAdBMfHyl91pCLbT7eB7O
qiYFBPvk774NO9YRLPexOMj5YgV4Q9ateq7s4ika8Ol3GzlsUlgI3l0LhuxJ2UGl
bjz2j0/+7YUfAzDg1pbWLZ32PkNJBi1efsmEdoop6H5dQNNz99GVXCbjW1QyKpS8
a08uZFJkKx6SfAa7A2ktq0tSSBuMGQ5XGxJ1Yiv4FOttqGHPrJjOFIk1zIWGcIJ5
aLr9x7uRNLTQxHqWzZgfo4MZnbQ05NpPrHBTu+4lF6zP6e4tnYSUChKQLnrjV7ue
n5Zgx//5oXF9ujdHY8bP7Fvf59MOvI1BrMaQKDqPBheFGH8RKvZWbJQ/H1ExFpax
s0udXoM6ibs9duHlxO/U4qFRIhK+7JaltSSTyDgAMBvDdtDA9EA7VNwS+TXbGMSZ
he4BBSxe5szblHJ/A7vUqKUJ1hpYHzThO7UCQYRLtkZKDI0oO0IjCa1+lQOhxd2G
cb96KXVMocLWmQqPBM8Wermg9FxP5CbbtCD18nCIjuuaOADlysTVtpvNAxUMnFPj
BPKasImsWmlfcHrd17s5S4DmSKeH991408WbP5fFcE4/hv5x3oEWl83X/VAHZw/w
LDzWoXZl1jVUsqfhgE+Pb+7zkzBrFVE028+IbI8RV6YnYB8Q4d86DA2Yf6YliegD
nqr001/rL+G4zaf+eNnZsCDRxr/zFjB8rzCQiR1FZKs56FDDVDHTEMP2IWsNm2zI
3idpyxQ4Fwvjq1WHMONlXjLk6eJ6N5uAh+Ct/QTMB+ylYe1u2F1mVIBo1yizMqQ3
qlI48ptqs2DW+fCuTsUno8VufzP1GVCWDJcfPxlZbjhW/obpbyccGxTRcgPjmvcC
pmlXBYidbHSVmp1kFu10kwJoSrPEudJaD7PTZ6g+h0AERrITvtnwPOMZ7cKnKYVy
G1fxzl80d0bvPIq9jyWHGLG+HpiW4GKccS8J8Ffkqo/EBHJORiPKzs/IFD8oLdg1
zBqnoWqR5eK4zBjXieY3SgDqHLhyBB9ZcPiOTops8NSMrLVhi5UnpQDqcgDgD6Wt
iIfF7h3w/Jhe+lHE/6+IHIqMU9eLw0+PXFd8GsBFWL0f/7RMRqG816iLno5Ph1Dn
PfogF5uzjECT/cEpvVo6hxzorg1MoTxbToYH7zEZ2aw45MPFOKozrtuniUCZWZbO
DVtWMzYNoMtzsV6gDsQL2PyT4shNF0M7lALo8CDpuvf7Os5UtxBExYFhMACik1Iu
kcRhx07n9Eie2PvQ9VszK1liHKKTnga1GdB8drSnvvDVL+JwdtwO9Ch7KY5D2XEO
pDpkEzUBlf0aCRa2FiGpZ+R9kma8IclY9BPttGzx+aUrScyRX0pU/meBTdLtwyD6
Y2N7mDmMI/tKqFbfDvtBxrAkSJoghXatEHcoWVJhKe6KyU3yix4tcqTB1Y25kzai
msZkhUhHHmXc6gD0Hm5B7U5VC9lFBzq0czTvAyKIdw02aMXo5IIy96d90gwztVAD
tAw959gbv4t5LZmDNIdnz+1+CFoOiuQBHSTzRjYnrxuYyq0UtYIeDgf0vHabuWwi
a3HqBgATETrfPYXZpaXhNc94ACMqD2wIgf4c+XyNFFR6pitCXu7oZtpYTpE8AImC
e+T9WaUufHO0s1XHilnRTiiVnm/Nk2BcILUJq4wyjC/31gN4huxxdjig9PcIxk/P
i/tS+ViM6wqnw9PjAHELOrIW5vxrR9ZTo6R1HJlaT0IKRvVmKzERUHBwlelq76oG
5317W13MXjpDoCI6Vduqsvjmto3+FE2qFH1a0loOQG77RGejAOLWoRxtJ6nETR6P
A06HucnxvjA/SLwMWnLazrDjbvQGqyKD08a7j2zh6ZbDBLDQjdl/Bc9o6Mj4Ta+U
89fkwi/MRPsthi7g9t0E74kuXFLe5jDJWYg65XiyITYxd78MSqMfkohacfi4gpl2
ZuembEThbokq2Ywx+3PfgGI4zJLoOG8qRLm+shjOBWT1CDBu8i4Ag8pKMgc41mF8
OdMgDdTm/JBfuDlfmJAb2vVBHeZjmyW3vJefPkj47xXqDjNX2CV2bjYALHJUXDwE
N7gK+btIXiodZ6/5t5I3x26Cc4c33hPai+tkDF2vA7dekITPlbAI5k+GdXfiDix3
eLuzMpIA3zsXJrS/YMMIft3kSUcQtYb3kkvtlka1binwveAUB2fpuOQ63yIAW0U2
tZpnbYUVNJozQAyuCwVyuPHr8fw3lcrsFLiHNR+0hhB6yIu1Njtspd0vtWjBXkY3
aX8ccBRWS5N44YywKIp3QO5kgvJB0kp2qkkxqnN2/WdAynLEo443uydW/3iTzdbZ
80PZKiMQfKnqOCZD4zl5fmhT/DEAwIPk91kaO7yvyDnvj3dTK27bv0dkp04m7q0l
gi91MK/wKjJJ1pwUzyuWdDA316oGcVvRm+N7qgX8NPxZES/bf5AK3YWrJ5FuoFxT
l1pcwAU8y3Y0t9Jp6ILYQg79752YHNbU6Szk7/thXaSMm7uHBywAkZonMRtzdr8X
ruBIa9ELjrrmajCB65EKIA9ljhCscoLDgJgUD96C2HFf6GY0c+qZuW35XoujzroD
bvb5jCX41yg8keaMb1rSpQMbO0EP82DpYrifMJvaEIXL2QCnTdBsfy0JEH34p7R4
ypTkhrCDSCogwiso/SbGcx4Uyr/bDtMv3odwKBerTQcALsJbEDPUhE/IIQAtWjaV
OB4CL082bOwIivCRvJg9JBOk34jNc8a/pY8+1hxpCbGlFkEZTu+C12m0TniauYLN
+nup8IhpHClbKnqT61Gpflz5Gp1Vm0u7kl0sbHGd28OIxWPYlZZ30S+KRAj48Mgs
m4Gdnn29Sk/HkCUi1aLLvamy+f9DhN/e+xtE3nrsflY4QzAGJ4TCmKQ5bIssiIt4
bOmPOITFCFNyROowBEHmT6UUsfVvqjYvmeqZuXgNCRZ3esKNcwej6B4DvBgMeBYH
NWLlfPuQi9/MBw/WmtQ0h9ImthHsvhtmsQTUOoxWcZytNK8baI99sXAEZ6nTypZO
mI6Bhal9ivOyaUQwJyOuhapJc1N110aPG4vMKw6QQoLdH+fCIuBBd+FEt3Eb8PtI
l7AB4PMxO/cXH6WlQ59AoUMUai9pxszZSci23vmcp0/vfuVx0hdVYNO2i6G7QNk5
5PKIiXlP0h7KeuOLZq9gj7R5faT8wLBudjHR7lgA4kno75ESFw3bd/jLFQYcv9BD
03MRliqLpQbkgFfMOkMh190+WfQvN+j1hMbJfnESIjhjGkCyHSB/xQ1tNuNluqKv
Mhj5VgiWEG9/l+xweVh6PiirscPVKAWV2TOz0s0zKxONydhkrwlwq1ddNrAJb+Yw
rhVuRtFoku7Lg0PbASvWY8HJnzVT0UMowFS8bAtQ9MIvyyQXJtLCvg4qOUzpv7Kr
apyY4gb10Mk79nAlMUMuFguPhh0kvaJhqL1lHIKeb6X/0xrQkhB5imjDQJ5+CwoW
ztcAlCp2BicFAg08I52sxsYHmGco+jS6STTaRpG8JJRMbhf0JUN7jL2beCBBp0/O
skiLvV+snaOYq6vQkK24xAMaTjFr/sxxopBahwGCEvPHKuG7wgAXD7uYwA+UynYy
E7P/JcD18MWgq4l/wjMrNIiTkkX1l1EYJv2b0FlqCoGUNxtqmNHMZ5SrF98UAl7c
AuOnY6gbmkqwZiR9xuIYV9G0Lp6NjvLbDNIc9pZTr15RMcjLHtb05dSr+gY4Mrmk
c2o/OHoG9caU+/DOkxxmPZ446vLsZry4tSi3DIwK5HztCHqrXqGzhg0kC1odo98z
N9bCg4Owu3YXOPwZwBA6NWv+XqIoDcvLhqeFN5Ebdm+/qoko7NEd6HF4x7x0kXmN
6PQWVvNxi16iT+4ww0VJV9QwxxJws8SvYTbiViqosNgtmKPtJo0/8dI4/4JWwAnX
MIi1oDZAEh+9NdP/eMX1GjAyyGQsBnepX41qoq2LpOc/3zHOpK8u9ZMr0j8A9e3K
AdHQHj6HBdHq9wVAJ2jERz8bRyfuZBY0bos2tyIBop/RHIqjrK8ZPBBtj64xeu31
mTFegcnD6gYTRb41BxgdlmavwM3ehPrjiEQsG76AascYvM4T3x87wqWwrZRKCr+S
irHu7V7T6dTpVH2bMLF5w6Bl43wBzrtMHq/f8RGithBI7tTgAK1gk8zJeusG/LOe
ck57GJ99uqUeuGpi5F9WUl8QCdrMx/eXvvKkfvE5oXps/tSXRp4OQPg/d9Eq/lbO
HjZwG2ZnGjldh/XcebVf5vx063A/D6krkWrjF9VXxXFnK7MiMe8hZXbfgSzH77oZ
pIoEtYADG4KUjKhkKlRqfrFA+gGrw1hYE69rnCPWOxVqD8jkcUYSOtRIS6SCPyng
nvS/3hdZ072KapzJpjChUAYPluA7pPgmG/ZHaJMPm0/M78JkByrkBaL8nMUrj2xN
hU0VkZ3jR+amK/RCVAkDEiJaLdwqcx+rX6ALhVw54DgTEZ7HoEMehgJEqn983CuX
e8zfe/E6yQZtulZLz+bAcIX332Puk21Jj8GFF6hHdfqN3bhTyC+zML4zk7Z3W4IK
pTW4ROGUdIK9yMIZOCObZrCUQyWOc3eWkdbXMb8WSVolHgXWfDuEZjCEZJ8vZSM2
pvFVKwo6nI96tGNZxaAp30HBXuD4PHdRIuI8obIOP3if8HsO2E1XC/7VS7La3jUj
aIAu8cU1qfjHtvP3py00QFCHjtF8fzcj/1Xg/cB7fFehS4EJcrfwHJy/IfkoUcWx
NRjDogd+FIIjk1oa451rvZ7Z7zOigFWg4hpwxQI98pnml/LD3Xmy2scuQchSXEZ3
Jq7zG1szN5v2tkeZ/BU5NJb8ZAhHAkXwnbO8M8iw4cvS3IwCtNiVwtP4aNp58I3u
mzQHFNqWd67/imPSDH4PCj0snFuNObCbL+dpDIk/8+Enq4hxpmZZDBfxeLLTKfHR
63zCFSRSYRs/vQjSPvdbozAeAeGyYqX4Ss3BjQmbRaXYIRvCnMo5vwrkwet8RIJB
QGdzYbnZ1HCKrJXh6IILM9ODwZYt8x4rK6fgGD8t7fY9OAm8kYhSayFQy3y5VXEJ
JoMkhlikd1ChIaEG6prutx52wS9sbNDBhsq+TsAZtTAH8sKeY8sLTo47qnptlXF/
R5A+8KpFw9Hn44cSB2RcBRhI4RnGCo4teqQkp0m7E25n/3FZ3D5Tb+2ZNacnc5v8
n3CKqDforY32i4gGCh7MOAiYsbBUia+I8kYpfTOrCpPEA7wFqiw/G/BJ092otxz0
LcCnPrwxLvgXbZJnVhuKUKNIUmGJ27ZBpT6ehoq8Fw68gil6aaT8RTOSwqL5k54C
KhMPAQFqyKuNnZiHCxw2hFshNgH83OUYdSL9kesa5bQZhimlpFU1liMyWddnGpFD
hYa+4m+x7uLxDXQT3Mx/0fUID9ij5mYHqw5lpW2MoPK0NzOO8P2PRjBHBnEorJLa
5W8h4MeQfeaVggkpAioTP2Mu4JxhwIvzf4qT9og2IoUk0XODQ9AHfyZZ6ZUgly/D
XoLFtV6+2QL43dHkH4LGy7M77bb5swD9ENpJVqtiV+9Q+1REHyGm/bEyONZUlErX
4Twsbo6vwe1IG8aWoDUFndfJenLatSKFd+I5n5IHI3OTIEBsjluwAUseC6ajDa9h
eoqagVWo0kYmqoW5zxeh7y5LD9KadXA7w+T8QQ7sBhVgwWF5J5zxo/8GlXEQM85s
bwzGAVrypALyvmhmveOp62DEk51uy+JPlwQnI3KFAO+cLroYJ9WMz6L4gTwMETTf
WYK3L0Bx+or9IKjpnGKU/lvURuhIeeHLvUrPaCw8MeN8PwEM55+af0BxOqRTJi0h
Pt86MFTbD3JvWF1pXe8MFg+axBrNypniEU8CloZYt+lOdKJFrfBBuM4Ses7+pzcO
2TD4VN8NtFFxkYDfzMeSM15n9xrDeo8VdLiiZgaeWUV2wMvL0h+J3qqWheNf2fh+
eKnGD4lNA5/gYIeUVF9QR3oKa+dIYbjpfpKNdN9I1gij7BxKVOHtwkW7HkNd4P91
Tm93EJyLv32LIhE7t17UETZLzf4vmIYcDNrXH/1rIsruUl31E9a1Nn3PcojbaAuk
KUbd273Aa59BgC62vEmCZgMl7B5fdPFfRs+nrA4KlyisbdR+EbhpbxjIV9XD8Nwc
YaZjseytanrnSCYWJZ9l0dZmr4sgYd+Eolnk66jmozPaogrqwxch9CPl5Vz9iCKM
hmuUCp87FxN3IUyvV3HB+aI9iRWQtqbFZFP3RrPRkLtrvmq9gI3udqXW3N8mewdH
3zSis5HVMsKOZs138ClIX+dprKx0I4RCixf4JAFEL2kdfNPVAgls/XipZ+mnebNX
5quPFBczuZfrM0enxhGpi9D4ig2zHYs643oh3khS4dJbrFd2PtgQnDB6mn5so8jw
5Occ3lAiF8FvzZwETbRSUV6YtOUoGnqYKcttnajeJz/JOg2OHK5bqfG9nq+RytHb
7ftaDn+0t/m17Bfin3LhjxO6itG3xBocIHiBkD9z0CGP1eb0d3AhYSIi0PA1HulR
IrroJtPx5iuvOiIwSMOS6VkmQqjk54mTPBpIsoe5HVKrzcMDPahuDef+HvY28bs+
8tu1A8CHOr7Tl1HV/BcX5HQCFxyvHS4UXukN4xedq5Bwk3KIqnJghAA/IVXj13ek
2D6hbGR1+wy3sz68ynzqr53h3ab7S1CsqSAJErvggNPsnWyUM4C2PNqK9POY62Pe
jPa2xD44NYyppR/ka46Mig7mHDE2VjN75GO6j674hGFJd+SUAjM/zfIezAESp6gY
WODPamqj79NC33UFO1uEfEzeKdOYVtADAOllYqXz0eaPtmSBPj8HDwGutmHheUpS
MiwT4ckqMlD1oaiwDWNNahy+nr2NG2LqdWCdRiXWZlxDp3MTMTpHi+mDWE5Q6LtA
LG84Ljsgu8XcPgO+hqXmcwGfJKimbKtoZwm+WfbBKeYDcCMKIJU/C8htjl8ihnyW
00cPCtBmUmD6rN7aEqHgUqxZ2H20GYQFQeKR/YMCdyKph5sbN9NQf5t/2CzSNAnW
1EXrRkhzKlzuD41FMrK4CgTLtZJwl0Mq31tJVryGlzUiL7T9iTCuc5u3MDGtGIo9
/dJuqPvjhoxVxB87ncXQHsVh6HX81goqR5GX6g4H/tLePVE9AYnxS27Lya7vmdrZ
jIXv2gGK6ALojla3YhTGRfm/yhKBbfKHFn+zvVmqRUUnrV+T/pyDFq/luRyRugXf
OWOeIG0iK3zNHystQ9fg1d2T3OMdSwuH/TqQ0sjJRoWxWbpspTY9VMONWSxl9VqD
RkoSn1K7M/kWtbkiaPLmTjlvpOYz+TCCp+qO6RgJNzHJ+MKiY+xmV3QnBbmG8eSs
rXaU8dJ643/aXa3peIgMIULwbYv2mUJ7UB4SNnLeqdhTNBGzmcfCTSiJr6l3LKSG
zhAvwQ8DmgK3L85PvwPMsvgt66Zil7huklDcJEatf+CEk8+BpmnfEXhMPDgpyr2G
rZM3QuIWQ+v65mS3wFq4NLhVt84+IcGAk2Vsi5nMj7jW4EFy9qLFSz3+RM9Mt3nJ
pEdVaOrW9SKcGUIgHxHF9G8VFQdJ1y179nyR8Orpk7ZFae6TU3wgyYhXoFRyNuwo
wvCFLKvQuCTRWvJQOgwHoGlfvmiy67a8HWMbN2XrjaToRlSzUGcQ/Tm0n9yOZRMI
vZvCrQOVcLFu+qeOIRACGZQ4yfuZEqWr3KMjl2pNNdhshraALF+dOOgR96EDKvxF
GAB74N+w3dNPAYPhMquv+yQOKL6WagPWIGMk1mLaxw2cRxOCqnbCdjXWZis80TZ8
RjWqVaZzATKYQ5fiOfQrx7AJbtWigQTa9xOOIevd0xM7BncTzsjhjFX2C0pPAkEk
dSmhUFMDInCG7fG/n4FOz0wxJsISfadzlee+XlX8gwgnaGj1HMAU88FGZtiCD48Q
1hZLOQgKMsDP47ezTR1JfYRfXnjTslrpO77EtcIQBbILi+GkIkjvIpbbysaXlzrx
pPsNOxUVeeJ1TrovxX/4OGER03c0FxJMfanOSwGjw4l6uDHRH6d1UAt7b67cv5XY
RqSwjoziSqquSCzjlfaDbKagrrit0dS5f7CchNplmPbmnr+ntr69dloSCuL5VWEW
yA0AfnkTPb3bmeFB0a1ULcilZwN8s2AIQMPLCPuq2TvakTaxIDeJOiY+FMBdazVP
zAHsN7MRBLIlHcTm8vH6sJvq/utxDFKKR7lzjUFwZmQxobvFRbCpAzeiyhlxojCh
g125b1v4+ojw4Y28qjcp0yDBB167WuKEN0WGnxzn32zuNcHdW3wgqHzdFIeQxam9
fUBFNKnCtdsr9fjBl1epJgoJBacsA/wmJkODq5eCv084lMFBtmRwGs1wdoUcWLAq
UFZO0Hl6qSbl1ouHvDgXh+KiqcNi5n9GSFC4VZbiUKDLms0dWtV2RONaY5b1VxNY
GFWAtfgDrTpKfzWVdlfIxcB40jqmP06vbzZqnP13JFUeuUDySqMMcy+M6jMYrj2/
6j4OB1pSwBYItPzT3SvA34qhsaK6am6gurt2+un8m05BGFErL2IsVqmh3iKEwwl2
ur8IcdYFLYzFLwxAlc3Fuo3MrLUOptriCxQz0VR5wwRrCMixLY9n8VRk/S+/Z2b7
VL3VNP1lbzomy1qq2wj7h1yhyjeJL9jgoMUFgArTLA2h+/GQoiSIZqXxR0AS50x2
MsnmOuJPJ0B67dVBWzLfueyZarPO2LXmX9XQk+JBLZtpRyaE6rIpvRWRY+vwkOpy
6+1BDGRFKHxsny70s8SWArHH0lC7lk6dxkPvKYLwTdqsEIGWIP+2tQZxGUhWZaF4
5vKROsUfodj46MugEGL0MgaDkWjS5uzcEeWQlwV2soIw0VOCcEO7XR7+j0LCKgGU
KLTjqefF5xie0TBL5inUAj6mDm1NqHYzbW7bKMrWI9vYsQcmEvbFBx1+X1dgnO7f
enusDiCZXy4mQ5TQU+S2ccQAdUvwKSzw0xPBblMSpSkWRf79NXd9sj0h2B7SyiZ5
oPm5gMHmEf2OP0zKV8Yzi8CYqAFF3Rij0K8slX71bv2ewrp45TMmA+KxpJVa521W
no2lnjV4uu9Befs+LTkb5BRK2rf1NkXXD9ezeldbmFwFUItHAcibPjPhCVdK1rSL
PwrKVywQrV6zf4xReo6u6uFC2Cqe/OpplFGiV2l/OEloZi1w356/DFSEtmh7Ay6J
1Z//rAi4di4CuQBMlXmX/6vxJn4dEgy9OV1/GYXKqYp2rp/RFApsvXOZZxXPyzrN
XryVPsmO/6/QGoq4eSzbJ4to79f+rj+55c5T8CKzNTpqdf8MsH1tlvdzyF/mLbpX
V8FrpWEf+ZT2pnJCixSXrvQU/EDAepTOuD7bmJvnei8Jl/5gEzBmvyHvJBTKyOBg
CEf2gbj74cEGXkHG30bzhLg7d5qOpOpbHJSTFCRI9RKqVx5LkA68RtGwH2L4Z1XE
fQeURMQNr/lEO/Ho39Udgf1vqkURzchvpAgvAKWv+GJmpnUiYfApduopU/dQlXUy
oUjh3uKOsAf/ImrjGF5RIBiSzA/rsoaQsPuHbA8UIADIYzelRc3/vzhfZI4FO2pM
uDOX/UbPxPtQ+U2G1BYdZcAft4AwE8NIaXxlnCT3aq5DLcusyarnxJQmJ83J/NlX
p5e5UrEJLadxfXHXLq6FExPgOSO0RGBiRpYTkNmSU+ZDak4A9DSLq43k/eSBxkMQ
pSympHGVqX/BzHkXPkctBNGR8hjOmDXzJNR2r6Wwr9sYX5zmnW21cPYn9sLjZRif
3cb56QB2HspUzZ9u3Rx21E4L4Oy5eX8H4hhmY2lDoKgqcSI+XmzO9BgoD0QdRBOx
0VvoO6f1KGGmEtRA6NX7vQJJAbkZc13T17fR66hknsKSUhPGn5FEWJwi79JjFa49
MnYl7k7KJmK9kYFkcCaj08eYk+/QMaeZUpETIVIk5lMB/azbfS5hzafFpkrUnu0T
Uw/e5D7zgXetmKbk2xI3fpTPiIKTSPDWKMAXiOHsWPcO6OxzjlJ3XoQbPTPVDN1j
esdVnIBdGFuUDCsyqh1gP6/NsCTRVfNgcdUrQ4lQhZsWYVc0nWk4oiS1OlG2i48k
K4wer9Ql6oKY9y1mXWBQ2nfUk/k8rSJe5AJrq6lR2wIrkdmudofdGfPg/tyf/T+r
tGh8ZrPejDWBuTDHQUJWnL1Z7AIMO3p4ifDUNw8ejXG+BLaVd8CGgmXEJerxYrH7
7n5HAjcmpitCCg0Z7HTCXUITbK7JLx7SSR1tSetWfVUrVQokq/m06Kue+eocrM48
zJjuI7aVElr23470v4jhNfitm54ObW6f3J+5iC36fw8KH7xD7SgVxB0PxEjK6OSJ
Foe0HWj8s4I7vBRcWEdna/ua2IHt0utuxCQmk5IuoSg9fBzVITzJwFhlOMsHY6Se
xG9d2fQtYRWTDDdKJCsecMYBTc3KtqAvrNn4DGdKwuc5l0eiKayQghZ85JPVgrK4
VjyZOdYIgGyhWpaG1mJhRBQfpEE2tr7QKDgFjwnqg6i16yhR+IymigCkSZ5v7KES
e3ESkdeJ33gk4JCjB7xx8EOOfK9Vlff+p9S0gMWIX68yDoTmOFSJr+UG8M7Z3nwk
xaK3VS0jg7ss3fFIhGoHJrwqGGFSFFVmZ2tn1neRLvURbI1ttP92Et7VbXQfYr7i
Y5xYb0cC6oE0z5R0IBJiSrdG4CI9tTRRnCkFUDfzJ0uu+ymUx/l1EwnIWeDIyXLN
YTVXVnuDpgV5xbb4AFyvOERnOD74tyWD/G3Hm46tpG53FC5Qnu6gtYFF0YKFkG3y
LDS+FZVc+LveSS30weFDYew5thtRfTcJTtVwSBoHxYUZF2D+GStL4Vf1d/K41acF
ad9E22eFiwojNyMOSoBjcHaYV91yIywPPyhu84m90yTeLUl/Jj0qywmQk9JnQ9Zq
Cjbzing9JpMj3ZaKH0U62SgJ7w2Cpk1cz2zXyzkOS5NPg13PVQ0vKzmQ+vi2eoUg
4Dka4iD/ptMBMa3//pk13a87U5AWaXJZEdZaToQoUhzP5H6QaL1w7B9UPoYAl4cX
PEs3/1x8IC+QwV8w7x6vhgLRRH4k5BaCG0w4pJFUEWsToo4ius0o6f16gYmeUEUf
81qx57ncObogQeVSlAl7hkORM30HGddC/WznH0hJhL9nIiGacBFrawAnLkP/kLF5
RGT3QhJGS1tqoFNP9joqNhgCFG6Kuc0lvSRiDKHA0f3tIYmSWmasesXkCUmT2ptJ
0wXNFNkUBe97PnHr5EqgcTy3gs3k/1J9/F+lSR7H458tGm5QuOUs5bllMTFZSTbC
f4X4frI0MndYAj/1RXk6wWdCUjgx3pSjWJ7YggDJjwl9nffgI78Bj/XZxUJfV824
3RAILEhIkdDqwjQmAQfJThGG/GC7eYbAsiG4JvIJHzqbxk9ZpOQvrrZvcSx1c2PM
QH3Dq/YQVC03fhM9OY/JnykGVeWLTOIYN4wn3dJGYV6mbmQ30mH8l/aNy5eZ1Wvc
MbV2UHFtZ/zIuSJXbnx7Hdab+3GzMOmkxnzDrOXf42EBydhAlocqFxrc6QUn82qv
h4GtK7tE2d9RWbUvCgxB4OADXSE8Y5TNECoiHFhkD6HrgxFJzJd3Qik8lIt2Q0iV
VslHRqbsOZ0/aNmwpm3xq5iO0b2z9QM8VgGFE1GJh1ZxZeLgj7h/RqYW30lprY9E
xIf5hFWqrFn1DAY8JzTV0baBszfRplqZZByev8gTuaRo9afeeGDkNTCDuFWorHB5
ZA3tG3hON1zl0Oz0JiovoNoznw0RZyNYgz6Oh+n07lRGYyOSCUy8lcHW7dpvY+iW
z+o3HS+agovMMCSePv2px4dMiuULwk0BGGkihd2NRwMde9e8BEOoQsWOWWrrYoTp
4q9qRHJ1nSVIMrzI3u/QZ4pl0VCO0z5HWGCw7E1YUYtpuwE9cMFa+xmMy6h2TNOb
4KLcEx4cqOY1yhqKwuTTeNSSHA2M4sE5JX2/BRp+bkmDH5gQ++VZo0FI/++XyP9g
Fad6EpPatp9/erXl2uD8P/RcOiRkyz6VHhJe1wtP0XUodXgH7HmEJe3HeGslo6TN
13zjg9rbuQVbHjtFRHCIoNAECkDSMCoeTrvVAx15cy0bmzShAlBR1nT2UpD0ReAb
VsNb4+SCObkFtri3yPgDcwkfGxYaOQLkUMvLE5yEvhYev8w7F3lzeW+RSGtyTCiD
GZ5buVXfmxqrOxPR4UT0EummUUhKVdFnmLRUrM+7vb3jXGDI5NiIoyRuvEQXFzWs
zNczJ/Tzkou9Zj8o5X4ttwC5qKoUNTdFL5TDeY89qp8tnOpLKzuXLaqIo20zTKIF
41XB9omYUxKTv7MKbV0bGs9scNFE7HI44GzQRH0BwIuIKppzs5WisjGYXoYLd8i0
H5kikrdsnvbdmDAYhoBfwTQuR6j6AzPStCwxkpMwxlkIrqNQ+srAvqqJr+LKHnuO
kEpfOyVcx+mqALb3CF2gGnBuayOIUGlMJmc6gBB4t14cWhLp/kf/c7N04nIQ1Ftl
cvH+xgpq4Jvbsk9NAnXrMZPPkPJDSVUsL1AVIax+0bu2bue4KmTvrGxVhnCimCLK
9/hufNeQ55Hhhciuo7U3/JCzcdct7xA01tU9PaVANYewWTIBFrUziAxt12fzVdDy
oeexOPK2rQ0gKRTr3hSuRtnpCWDedUhW2LPKf1OQ00LdMXituZuSdH2YLRzGC869
sf86n14sLUBeTl0nfC0WSJp4+7OAK3ajxEzIe0UtDF0D1GMPBPfBTZJpcbdDRMgH
ZSCeCQA9xUIWYCQAGqYD1mikDhbg3T63IPaQgmKcNOZOZMmbrQF9tFTqAFgyQdZQ
0bsW/LDRVd74NrcxfcYO1niPb1vvrWFMfyC5m6fh/C3VR2ULfdzAfKqhhtHhJI0G
DgY1t/YN8IFnJum03/n8Gzlajy87V6ISyg6XLdXBldoWg3+OkN9azgWvF9YE9zb8
EKT+ayBx8L0Jb691DDQofH9h+5zbq1GzHdup4xEkjxdk/tXEOvrm1kfXkFWzVp15
iMoRdg7ci1iwpd+Y7ptzKaZP6JW3+skuOyOBvqO+2ke5aQxrXq4L2SA3y1LfcGWh
2PElv2SFwIQbJr/ucKM6i730LpD3A8DcdsMzMWd2FXdSrEHbhYCgv9ZWXOu7FtkG
9rVTOy3t5JL8hIcFfZslZ65CGpyB0DRY52OvzaBXJNt3+mVelULnP1/rHlOHnruO
eO5npqFb+Jma3XiL91hx2WKBdPdF+iVrK7s7pYfCt33X1Nb5p10STqffl7mQJjCm
k5jeS4q3UjNkT9yopjlrGXEZzsOr4rN5O2TyQ1pjxGKM2LipCZX2GPtFb66Jf5z/
WyDiKam5qS3cizlimhuUistPLV3ftBSAW3+FQSIugLn2N1/b13cXkOstRVAZ8mOv
3GfeWULZ30zz1NbfnJtQwomE+9jRqCwpxgJu1Ccepq6G9LELT35fdi1yS/XpFTmQ
4MQdZ81ILNMq5Nng6n2ziu1VM9Zv9/nyXCYTMxuYSg4zV/AAoZ6qkVy7C6dd7wHl
MSZvDmKPa+nUrM/VeRF6w36Mfp9ObnrbqRbhpwwSTAwBYh0XrqcpWcuGOtwibzNO
N+Xym9yTUaJi6o9MYpiR3rJInrPMWH34+zCU+jm7BdFsKQZY4ak6zhDd8J17vggV
4J7uDJ+6MS6ZHbgkf27sbatbw3xm9WqBBkDWioxyPvcmC4VYplBA97MwO9h+bJbj
gXDNZwzZj7DhaJ5e8DAEc5yUQzeK/3YoHGOGpr/KqOpSEIDclcTVV25QSCFuUuMJ
Vv00rnUKLum3C1b8pKyo7hi3U//UxdWSTB7VKLnAcSsm+vGsIyRqBGZ2nUJmTXw0
UYR9gcK0OqhFn6JvRQcvpFpKHbTM2HCMlGtAMqL4nJzBG21b9H2kNYI/CaxnWR26
IS8lM/RK2hfnJbbdmtI+DJZkGPDq/AuM49b2n6uVlV8VuHHlJo0j03SgK4ntXsoy
G9nKqZ7DenbQF4MKdHoPOvsU4KOekI9OikQ4vvwb9HsgUgqFxf9G2INKoUh4IBqG
F9REtUqXDNIldcttcjuWeKEYqTCcmFnRvyoqIbVTibR3Mr4UzDkdIBlKNQYfviDF
btSauNDPlrXEGm3et7P46V39AM+g1VjEfSr1Vpuj7YrgYvb8nuNA+yDd5g67ahqY
L2PnBVu3CQJnBK5Nwzs0bSB5Vh1F3FkTWbs8HKxVgI71ubo1hFm6xtOGPPxQoS8/
cI7XefNkEW+dB3qS+tZ33xnr7C0iv6qQ1ituFxS37B2E8g+dJPBIOrWhMNZAhJRQ
h14WFRAsgot+G+shUlmOAdx1tHsV5AcXFxtrhfapfnth76ce+d53NpXCBLHzZa65
Yoml3WunnFNw5aoztN5ZJbdyhxvs5BXUVY4skSoABHYz4QF/+rsvGg2/FPj8SEB3
nKJNYgT6CVbsqTSV/Bzf26nILQjePNEzU3MmryoKIbonDRup44EcasjzDQlxQ5tc
M92o6GXA23G+h4TljZu/LFBW0kwh8wPYSWLQ+fJgFl+iH48vX6Td4iaELYgyg+Mu
Td/nH+UXMe62BHI5ONqr6xLvf+vf2CCq7gGWlFI2zYuiJnNFHfsYCPHas/Ry+E4p
mp2K9zt6hYUJE8oCNntrUpVjU/jJXEcbJXAxW/5/jyKXAFEPYY1gKRdcJGYrTHIy
77vQKIg9ZUsmFMvWHc62jPyinBOwbG5SdDAYqsu34cXSoT97ttUc30qEupSrFJnF
xNk8A8ILcldF/nmznRJ5bP02CGsy+eF5bVW82AFrIGJfDOfQXkccEZo0rxCim1la
AVD2cofcoBgvi/qLMdgc22psRKmO40jB1XWm6kkDUwoLsiozYMsD9RqqD3z/S8My
NtcgzEm9Hp52Xp3zkj1WoqvCd361U1aXuAGQbq1xCJIATOOD/7kkOhbv65iYuF+z
0yPXc0u0Uan5GLitZbbiGyHkRDMPiLmkYZFlZhWlphtDqznjvaUTanob7wsko0aK
NUpykArqz00Igj3HLMQAjF6nyjv2/7ATW/MW0jzV8COpIisyei01FP6xGr0s62ac
+bMoIiZjDlnzag1Khlyp5GsGF5r8/jL/J4uAD6Y1Jyls3C4CitcYYGyeBs4TXn0V
mAOahSYmLI5upRLhZO85K26QWVxwrloWUuXWT42NJaRJqMySjTh6xCnkFNeOn9Te
c2maIcrzaPBcy8HFh0+Ohx17B+580zd84DhAETcFBHqA7aurgRMO8ERXxjNXPjg7
L/WytT1t5D7bVPfx3LTlPJrcZg3seAU7UJP1bQ02YkWQFRzPyM4MZTdDdhA5I56L
EQrp8nekOUY+4tnvIg09NZFmbklV1VA6B0C9allWLFhhYhRAWLdM4gd1MKWw8p/J
nIbaEt6XgF78EevqD4BjL+KqB9Qrme96GjnPmvKV/Qka8BGbFP9SYCiUkULzKdZQ
r/QHJQdMdVm28oC/93XzKxkFBwbqJW6RDrliFyTNltegpu41+pGjqX7zgB3dC60g
GAy2O8/ivfvAzyczA20NzYeGZn6Bx7892Wsk6tmJURHszRlbzfk7Hr7d9xxXMXW9
FOmLW2hFQE6TsXLzeVOi8BpJajRLDMJvloqzVbOGNp+JV5HYFoq8k94iEv9mCQSI
fyX87ep3Kj7Chk6LsrNyIZCnWkJtPIlysWLEF1/gir0lzXmDLk1eRhDfBkxiFyb1
ugJ0UrUwBVlPmDLntibmfkJU3PEzlYXENfZgTDc7RRPWH6Myj8cdMYmA0e1w2dNF
ye7iCStr4oVvYILa6OU+au7pRdnqFhwhrKcXMnXEnXFNtfKC/zcIUWuzz+nAhMj8
LYvAnBROqhHnO99+Coo+7xR+xd3jyw0rKtPNSWpLjdY4m6D6bEqIpvO2O1lg/BkX
OAD/WW1xyEQN63D0gSXpdgDxUJKmMrcCoX534T17mFDk4GuyCKMdFICKYdtxWQ5o
mHTZNPvcg4hj43rWWUa+MOabVeJLVH4qhWdye61rg+2G3MWzM/JfsxicZpQVov/e
teFfcNyrexOaJgJs3xnRlM3YBkO+dg3f23DU4W0JwebqFO17B6neOCJ3KnkpkD6P
qxcsONx+Numha36INwhgSmq+ait3+/XxeDzJJlGNrbsn0sEGcbhj5TRwwB0yNjYu
gsx9vNl02GffXEYbgHsoXdfXiVlWsot3Ii8LnrbGQg4cs5IKcbYyubBSiSpsBW/8
wDu9KLcW1vEL5oysBRnByk/YzeYXDPDi+hgA3G8lLpCkgIAXzO6pog0BNY+SVaWC
bfXXJmfw9dli/GL3xqXyegfs41VP2crXJ8deFQWRfSfa+y6h/llsKzly2RSLgtSn
j2rxOlm4Gefe8CRe0Fpp8zkoZU4oegD92xmaIJU+2aOJEs33ZGSKfYLTNPHU6OgT
oExjSqSXCmPK5x8h+X3xIBX55XOMz3D3Nhv7xtyqUuyylddYUQLAjCVBxaFGEb6D
kxUJxUSn2q6FHuA4kdEvVLjA+KNORnHVD6YvDFvICKTo6oZif5uNqODSTt2qxUc4
VhuKkBSJV1btpWkBFXLu/zh8T0UmV8LLE0MjRrXel5XN9p/9PQD7eEB6ehtKFEiT
QoviXGx8Ug92bNP2U5M0sqQpwe8WYMFOaS7ReytWnMEtOON4QeoC6i/X+Vzal5C8
xrjME/u2JqyKsH+KxobTrQc8p18vvCjcULRUDNc6uYb29hGsXjVX75NdOlvTXZLX
iFLyAyqf22GNwmLghzG+s26pMlGtxcvMMhaY4RZjLJVN8BarVbJbGrfVPCekj3yN
Ji7mNfAAXNxEL6p/Q/f9hchxPInecN7IQ6Ly5+k34X9Mgh5xvPRwMaUO/yWDISj6
5sj0Jlzhj4xsiJl/zhnNG8RVCyneJPHzHGA6Gt3i5gpiK3fN60R3fdju4Puoo3/E
TLvLZWh8NNEhXf4ctAndK+I22uBcwdUxFJ8SwjylFLwd3mV8VyeMOWQN5JKm2yNY
RJeVaUPD2sTNNvIBhiWPVpjep/RkXUriPvEji2CIyB1TYEQWZL9607dBU+WX5jtd
RTuRM5A974K4YnxCKvHHjJERyIKkZTvj3jx7pBvdbzqY+gsjr/EfZ8HJg7tL2p95
PFj98lM180tdXo8kJfR8dhADgxNNZrKuJyiPxWQIPEGuG/sOap1qcO/eiefuZYPs
YPUftgWpecqka+JsmmeA0lQZbpmKv+re9fo+6AdKf1h2a0k9WH02Hivmq976i/31
FF6R+GDwLRe52miMgm+oYgkPlMCTNMZtktSDuw0q9+uYp5LSaVJcuyCknyMCBaoL
AxPdpcKhJkdH/1xbSvjoBdiF2okTLzKFNCYzaCGomsLq8Iy7/1N6lmpbopfvKtgn
/rLKJJ1X60lkfD3AI5uEDFhWDBOqqGJv00cMoool5oU480DmG18bT2VkHD+QX1lC
GIIu8XaxeLrgYYyetod+MMMwIBvh/NCctAVrWkgqyjVRZLy5DliTjcx/ukjQMWQF
3ekTFWR/dH8cz0u/KBOI4nz+HJi+uwvWPhI8+t8R3gZjoBFutTphRwJUtnIWpz9Y
TVd+ET2Tu0YobFj5F2rKyeEYgdnMSkZwHXus2e1EMmrBdvPcteoHarzmes7A+Pcn
Y3hHrc5Hv2qJbTR8Exg/8PLQ3HxZvGuFA3sJVjru4SVJqasnjXZJfar+QQI924ve
OI4cJ8ZtQ8WwGaSGqAEvAKES/msxrrr83tXeAmMhAh/NZgyuJsEW0Gcf5pHbwSUt
W7RuJkTDfO3cexihLSpx9SoLL/oXudXvMS8ynq9XWRY1/oteqXIiPoS3Br//DXvN
eFW6tvFfLOQSQMolCXZLJbAikfVlslotcN9hmOAGk3BbhdhdYlEPesqLcYO8f78W
NQmUa0AEAe254poXxlRWRzIrDk3CR60ToTt3qr6Vj+LajMwpAefc9iJuM+WQHrIx
nCeWg36JLGudZgQyLqrw9a0SM/u1hvBoKVrApp8JUpJRyprmMlkXjQvtlFZhknRl
V8mKwIFy6c2HyKEFqInG24EOc2I5WNq2uh3x4jFEztCDAQBHPPri1S20rj4pDi68
3Hn7KYioorzEawWjlVRRbPOrGO5U7/hAe/h14nialOuF/6u7vkxdmDlzjPI+Vyui
NUI8bVLPUAAjWIv9znlWVasZo93uORfcD3o54bHKGK2bfiphtNfccK/IgaJsxrlo
Y/OwGITCftIKi5k/nUMiN7Mb7QDZfaG7JGQRXGNhsnNgXWYMGQrCtZxYW8ITT8wk
J3tct35WY16fzMF7EyM1Vj/r12sN4i9gFd9yEfyKH14vcougHx7SMKnIDV8w05ep
o3y4bChbLNqyo/XldMT0JazWoVp81fhSOGkC2JS6UGPdTuRn7GcJz/AASiBFa+0L
qJ6GZ+qpwkihO/J0n0LoW5Cv1Veyb+y+n5Qvh/k2KkJUAtzgyB+XKAnDl8pQlAlJ
3NrGBoq0AiPSdWU2yjDdS+HEFst38Y7YQGO92QuUct3cP/GRIUc8Aj3kAScfH8e2
E4ay+2pKGxDK1+g4ZkuiUSC5Reayv/E7TFqNz2xzdA9Tkd0xxHvJO+zui9QgCjYq
J2w2JL5e0jHC38g0glGD2f1Y2+vuSS+hzWgOi7KUfQy41ibDpdz5AEN50UsamgcE
Wau/z2NXWkdYnnSwHnivczDxuk6wvvzWiU5ZF4mhYB53qrZ82j9/TfwGMcqQRJUM
b6oDvJWAElL5a9HpVmbLoXOayKj5wno7k2KNQDg3psLnJ2w/0uX8K4GWeoaQN/yZ
tWxSQO9b7VlGrpzBMPcdCQi+kdIBZ0DpAuTK0iZJ/vCwb2AGBtF1TcPC28xi1DgK
joR7oUZrkyHyjGU9h3vfcWM8sr4EVyDN4QvwtOzn9kJV2UU67uhn8eZ9amPIz8HT
ipy/jlN9Qyb5Fa1ajy9FVrh2LTeVlRK+WKhrO8x0AoV//UG5KYAXZ/rYykZCTYgV
XOwX6tRERAxB4vGA/ExS+QjO3MgjDKVEwWPM+ksUx+v6vz7vb/j7Bze3QlKcoFv4
rj8Uv3IhdhraOcAxj3+oJsfqyKSliNQgTv70qXaBv+EURvc4KcfdZ7xeBaC+Yavv
cAK2VF+/IjKEPxuFJeJ+jkfd5JDHm9njoqIz9KKTIF9DR86Jc6foegGVSTyvvmO8
da2a5tyklsF62RCyD6RkBx1jIAexiSpzoDZf9W5OPfS+9Hx7wouk7GEnjb1xiguf
MNDXXWjSUhSqfDah+lsEcEgL3nnwyWKkZH19nRoJdtDlZrZqYXjfFaFq0aXVgj8L
RwW1lUGYua30YbbucdjL4yz85xVm+EuxpofTDWjFq7xkBh1nUGxzd4+Fcq2UZNkp
C+wHa/5AfYVkV+GCJQGXP5q7sjTMVafaoLRUGbRK/MKdS8sMcq2WmdkW+Kfyor1D
jL0xOTRy7r3YruHJIceBEZ/xDWXbUvIz17jmjtHCvsC5FHCi3bAOPsPfGWHs9miq
qFyXyTHFq3gSGcmWNlgjqzC25N+VRZzU5Uc7gQS9iLDmRXeuNt+QgmLu1+44BJb2
ePtzQOAFO2OY3qV4Al3nAzZ3W6cRbMSi4xNldPs4YiEGmhRhSZRmy9FjvjMqH6yo
IqP1/WZ4g0vAdD3i2ra6jx1B+SRFcZrig7PD3koAqNZZkNEIJdVNTrIdhGwRl8ip
Dwq/moOr/+Lsijto1FeG4mhwOVpELi4uN9ScJg0B0SZLFhZUw9Q5bP2O0uciQlC6
FIq71pb1WcbGRF8aANF5P1cC1BKuSRCxqO14N2eLlobOZMlwGFv8OO0N7sI6hWQZ
sTeya9S6n88G8NZT9OeamKEkf64dGpN3D6LMop8kc+rsgip0XFf8xeLXDgPcf/V6
J5ooWEAQDfSWp13t/lwyoRkQox4bue59RcjALJWys2BsvbxjAG2E5HMAStuQ3C/E
iDOBmlfQSH6jYtNpnr54ZU9cg+2RLhK2UHrK6C59LwPWAmx4QWXudklh2DlZl0nG
37AHNzPvKr+s4/E5/lLu7evNMWghTXDN/bZ2d/c3QOtoWZ7ObTkzdgJc3vBJDkSR
hF13B4+gABcV/cyaPqC+Jm5Rk5icY1AC792V3z9H5q2JQ+LBohhz+UsxlZZedZLA
8hnUIzxDpBAr7KRFF7Gj7yh2TlA41CbiaQkQcHNVe1R8TrA+Yhx73+AxnQtIKAX/
Zf7A0vYoqsuTs9FPdq8iJLNTzfSvFl/UH1HDsO78ZskMU149VJAnoXCl4CUPuKa7
TxqlQe3KadR+aZNsR4aZZmQ4vm9/1Ts5DvJ1tmKV1wc9hezYN457JvV0/k07t9gG
Q9329nG/VnZ6BD6lDEmsyeWurg9nyW8X3abFwaxKCLsQStnsClW2vgtIqyyY+nv3
F9pLbLIJ18YGQZxjHDaRjw3WNkJV+y8oJo448UIXayAY9nLCSw/dCyAMNlRIXjos
aB72TmD5ujzQcyljrtyiwbppAcxchtxI7F2wN6OOzvI4NfDE5PfE1Yc1BN6hM7ku
/RMd3O0iNhYmOy8mKOh6NKroRwhxxOPN+fzmxLtymWCaF1uV2HBmWNDL2HaUh0B8
s5AyBnXhEZWp66pWDhd3/05pfoS+n0LubR0tJsgwp3jggEQyL4TrxEeJbVyNKQoc
KAaS4fXCn7mO+U+Qi64t0KVycAXxRHYUbRqINHg/674h7crtq91ZKbQKJBK7NIJ/
n1lVR/uss6soqT4u+V4fV6yIBTc+6zaYRBJOE7vVk8gG2YErQ/0mnZcHeyPLYAi0
oq4BC15Sq5bGcbirvmoJS+dGFF+PdM4y/RBPDgsjKPrbcKKGsIJxMepl4yxHQ9Uu
BAWCdAGJutFQ0ydR048/DKIKJBX8U48Ao6hwhPK/yW6OQaaip0K0+2AWHRYTJ6Qh
XXPeGMLKxfXu8VBblk6WVY3uT9rl/6KOxPIe/fmD0L8NZozms5C7/61yWkCZMvnv
r0yKY7Epo7RLVQ08zU6so+awpSptCt4l7OKz4N/giUtRn8r8UqbyXVcMMOepzmMF
aWUa+Oza74SX2sAw8jFqlMUZ4MglVhV4ut+7dyjjC9XNiNyIdb8jnzJfouWR7Luz
xkJyEDIv8SVNj/iY3Exl+Trq/dl2k43GEh7BUNJyPccvflvaL6suXtAOM4Z5kcK/
Ztir9xZS6p5OWfYc1mDLgSicp8TRDqTJFHfwiO1KqHW31n/7AAua3IhLj6/2N+m3
RPXDWZgg2MG6/JbnRWAxLUM6WlD+h/aWvZxm+46xD0fqgnCwhq0+etDWPtRIcCf0
CDqDc3jwwzFOMIuuyxCvy0l4kIeSkuo9EMgUnsXv+BYLnwvGBlE67hZuDH/T0bNC
5aLo5WxGTFJJynA3lR08Zlc7/Rws3LP3zvh4HA/U3QSfljaZq7VHQQtapzk8Q1y3
MWcT+CGpv/KtAIeS/L0YBidAuBwcyrtXU4Mzj3UmqgtqXh08VzWUSZivq5tl9AcF
cjWJyQE4mW+QRBIwYeHPo/E+zEhTCqwW5z6vnZWtxRtx99SOuPMotN6N/1bwWNdj
4oYRc0G4ZWOGQSvucl/2lp7VlbqC7BH4wD0OVSZu+CEzPEaL3qNOam4jhw2GhzNz
/ZsEeMeV29CJEXuOL5rEK3D4eIg/utgWKqJFYXfmpRSc+Zc5cZt+1bTyRQg38Ml3
DENrmGIwRDQN2mbnBVaqjpbHn/ekxkgPp7xWzGuLUHcs/J7TcEbDrsTxmC3A2EaD
GJi4mCt/W0a6NkaXr9siOAs3/M31EFt9vQeDij4V711h0F9fV5Y4ZNb37BS8K/s2
SVpfx3xc4uzlkc+L/dIyEvARFG4zzd7N0eC53mXGyKBu8CBSDzg4YgyJi2e6mFUU
tcs8Z/Ezp/9FxIkGvGcaAHq8ru1CvR4zQwQNYmyL4X+YHFjMWsvQscQOOdAZGt0K
m/q9JGgiKldfc/16Q6GTcB+pZmYO8kvMXF0hE8S80x2DT5l+X/l3I1cCsA4GTqwS
uwJA/XvqurXcQotAz35tOxIqsBsZWFSWwGCmstOEpGOJLuxmkG04mlDgDeA6a0Zs
TM23xPBbRx55W3EU3ECa4WaOvTHMGQN+KwzTtd/5R0DmRD3z81SxxtyGhH+3W7qD
nKswixlIHL8Qtll7E5MQdQHsfOldJ+nUpWZLgJlzYg9Ij4KlLyVeXarBp5xVqKiJ
kDS37Ai5uXkSbV8wZjLbYgWPr47btFDSk9VAnBE0sXx/00v/VVl0x/6SKxRl2qCA
Ujz64keyonPvwuAUW+HHT1vkLdTO3CTFgo9DLWGQPJ10RK1cHzBTp7iGlxLWpAvf
Q/oagRnSHwWIgkznyhRHtJul0UrnlAaSOSv9wFFYDc1H4YjFTOlywJvh4h1QE01W
OYAwBX7CY2mRXDVPH+cMRG2aZvpy4U5fzgq938WYqc9D9fd3qcYlEchTGjSCjCM5
rMVT5URVrHw6GEBoK27mT6VYVG/bhBRXTrpC0NyqRlHHjwW5WauH8Qw78By7hyoX
C/slbmrrKP4UY0PgEOqVDIRL59YAgerDmN3b5uh+bp57oMZprCwW7wGTnX9wiBmM
ZlI6gF4U3xsdDcPWV9VUhQ1xpxF50QSb6O0wRaNy4Ymknzz760k2bJqLQCVWnWGk
OFHW4MHzhq4yt4cBl5/jLqC2jxBZH01TSRRKrkINBnUs8BxkPFOVw6nvZ5P3drEi
ACodUae+Nxoqjju2cyEzrW9pwjbPdzZSekHJaqHJ2cC80zl9w9vbAw7JKBpAMx2D
xC90HxQ9O0s5yWgyXdRGRPobov2b8Pi0th5ide5gMf0IWZ8gD9zPzuc4E2r6x/9Y
DwzT0nkDeHboiHLGumv39w5TTSW2qryLjcB3bJxmaavFtzsCH85A+jfE3vuaRVtF
lSdFytrASjyLilEAgaVOcqbK3fR/tlm3Q6FeTdbIKAZjKCK6yBulGWbJoel/e5vr
u9kWc1qLJE3l65XzIjlr9YrJW4yLPtPA7FuC6Yi3hHMpKwaMgR84k5yKJiiINvlW
OtNwSeXM3wOQTL7ZaTjHVRYJnA57TH7Eqg//Y4U6eI+w5Vo8Yrt+/aDeZF0fuXrT
rAXlM++vgN36XljiAHjCvv8Gw1655I38kZ8FnYemTvqDNWjDXQnkzqXUdsnbMuka
XDVJJ6LuOmVeYxFiTuE/yIBxFHzSR9PzWOBg4wITGSNVJJToj34GM+vrTPazmvTl
x/Emcx+JntIV25l/25UZqk58IgdWefuJJrNhvH3OLA2yJ9WGeF+rFuDXkS2vij3J
hsBcA6M7ufggdmRKk4JTidIggVsbLcr7aT3bZqi6IH0nQtL8ICVNuqDKASzgHTSc
IB1+VXyyPr7O6nW/uLDP24PTKWhrvJV2NE8OhhoRwiTrTRMCuEN4rv/ftcMR+cLn
hkEhpe40+e9CYeZUnP5Uk4/0Bs/krBOKv8oujK5nKl/TywoSMllOpOxmWy/m+ckB
Lhl4gJ3leWiuNyTfQejYSKujVL/a1+eErICbywRcej78V7kUvxuCsiqGITdoYpZw
9gpGR9YdLyBQ/oVqmG/IN2853tLLKZOSmL2bkfTfhq3bhonqo+v9wfHBhZwft9J+
QEySm3yzkab4nox2gLmVQwyVuyk66vveVVwo8MZadrLySn/SIdrjbafDo+tJsQF0
atQiZe0oLVXUbD3LtoBDpO/FNfB5falAgaXhEnyABC2nrhn13pc+xhLIn5ppfSyW
JsyDa1IqqiA/Tphhind70JKWSrAGRu1PQ3l4wIJ/uG03tMYNsDpyuNQ861uGm5Kg
Cb6CiX/wdqslqDbQGVqu3BUd0hPs/7wyDBmlrtA0rGj4y8R//+FK5fbokPPz2jC3
IuUNQst9TR1eal6KDa/CaVH33i7qhhawzI9PR3pbab3QtWMh6heFOpgy6RtAhMMv
GkRVqvPZRyonsy17lawkm5bTRIYLmn52BeVP5X+frZNiVtpKeGen8agf9NHlWQhn
cMMwFWm+2Bv8Woc/NDykU10VeUBg8vwSW5bJBpp4/Bh6JMTTUMiLDFMsqAMwDA6T
rKlw5z7fojlVvQeH8boPcG6lOPpeoQJxsP5BkMsvEzlhDCqrE2tlzudDUClN59I/
vpoLuCItUpCrOM8eMFmpp5ZjyedSCdeKXhohCK6b0uIX+NjVgn6cPKe3NBSzHu3c
718MTVJAzlObsVTGzlYUqSpn7JZ+qHGldE0LesoceeMjLfuawnAqJg0uz7M94zCY
QNKn6tVLcpqU89gc0Aeso6CRRVb2j/x1WugQbsBmNaMWFrbPbQwgcS9+67/9oU5L
MoCmlo3DXtR+03fzHbTnVC4CWyyN0UTrr3Lzr6YsfRE3CiIcht1jWLtVIPzFJmP5
RKoWsJQ63Reef2pHlpZ5Lf4C+hLKwwGrlacayV6tBMh8JuRR0W7e1P23QIQzN3ae
DlmJmKzvY5awIfnh7OAaJvujxccLVqIRZHivJ4cGKjicgGuvp5c+IHnLJlqPOLFA
KlyJs7fLgVHoIWoOhBKJd5P3UaPooiLSLqAdWY7fBHsF11v0sHsBQpr9Of1HfjYi
BBao8+yUMoidlVVfy0cWeG7tspkB17NX3lXJlxtEfQbzmcAxA2HzIdRQkNPBBkXZ
6FhWuCHFKAjzHeeEQO/5oqnB82iVlciLoIAGgOjKc3W+at2IoRQJWKGcup9XU7cJ
IGJU1BrZ1hCHkpdhGX5ANz5BIfqUCkVjrzYe63yGe1j5KnqU6ub9DUfpp+OISAqA
pv0HGZB4SUkD9WIaAFCfsCmGrxvnn5h+5p7wyVacsjuo1equOFoFAaDcGEaJEkyy
C4VUwl7XqE82qu3ZIjqiEXbfHOialvhXuWNXThI4jlGwY3tz0FrQHRvvUB06vjdS
z5uNtONO+16HPZ6PrMAFUqF7czlsU/QcKn+4NRZvI/0xQR699gaDknaNAYyPfJaB
JPlrspz6p89/GH4nI00ocxiXqD0Mw8pCEqofHtiBgIo1qGrCxsSykRZFjw3y7ubx
xsKMNF2C72tr5wLO4bn5Py/Hjl7VwnBGjxuBgfQmbsmcpXO9ycKLfV8MjGhjBFYq
kkBdt7Wc0+YscvllIHHdAWAd7zEeuVtz3P9CXrLUZwhah4lXBFr+X5/ESYp0GLN8
M2cJ2CgOSmMmaWgK6rj3KtIsMrZG4t4NlZDvJhR6f6wrVol22eX6yc0onYRdgs+i
64efeQwOx9lqmsjCPuL9Di9i11oFr7LJ4t5EnmWKklxRmjVlkci8lHaUhbD1xJjf
lrJKr+gPmnKmmggS5nxRZFxKqhJl2jMRILinuEa3IOc0PoRhyArhglKC0utUFRLC
ZO63CbAHWy+gbG+BfwTrGWuHqBVl6F+7X3mSBrkt+M5AbvbQ01+g++mq4hjA/tqm
unLY9Va2PoaxwiF3+m6IGJ0h4hFZqKlVvGbNMEERtaW/a4IuINuKIOOVjKLgZ7jM
byj5I1kc3hclzb5EXNwlZrH4e2U657aERMkiXMsWkotwxLIAs5BCFD0nH00Bpyg7
A8obxp2fssBRJZWxkvxsTcXleDqF/2fXpwV3ETkfSBgEFAtXZ86C3oX/9qpvRTOx
JwLwqp3gPoqeaS9/nMpEB9lH3SJBDq4vl+BudeOkjqRpPlFfRaVSfOLe76OdE2ix
0HfVcgEAWxC4Tea9y99fJWw3NbLI7KLqSi4Z6meMDF10OoPtg5067W685nPrnFC+
DA9HWH/uY+wL+zTuJ2hcioz9SAmnL7mcbyn6/EfZpoMeX9crUWOV674Ed3dxI1VJ
D55UvPmRMf3AhempLOsB+kwem0De25CRksgc8YaTfa4toou4OYptOpJ1ua96pGEb
fzCIaeNpbVolu1c307e4LXpkzInydY9/JX6d5rwStnRrytyQdV7uav+bI/KGppdd
iN1fM4tYkH87O0V6iDXlCCgphEhPsoDaO+AIJtMhrPT1OdhDGwaD1L6KQUfXf6iD
rNt4fyEl9jZqQMu3KR/n588+jm1byWh/2WLuDySLoxJE5NdkdVVyqR+zrcaqt87o
E16XVPyWKWqwpNdlcA3GfgLhhe3XuYIQ11Idl68BCVTTXoO4elSqdEBjKDqLENvF
TqJJ0/r+TvtSek9nkaUkxdtKUcsyyOIHJrl4vDLwmz3Xd+iEl69zdmdwW1DTJcig
2IBOVHmsY03N/kopDU+WELEDtJr6RvMuZlH4l8nXF2WvdHAHXwfimpgworAvBUPa
bVKvHmQtX5PMROdN88fjtStAgoVNRE87JVIyGCnt16WI2YQ1J3pzNOE/p5WsoRkJ
eO59kUKfRC9tgwM05NPXB0HbPvfrxT4HJyd3+nRopfTYi48hRmWAkVVuTHuPB/FV
ZIkfOk3G1Fxt1P0bzGrSYv+RQw2iN+P6Pcf/Cjzjymh1+YohMy6qyGoQtdQW4L1E
SAD7qQJaEath5GnWIeRMtz0WUKk+Qvg3Lm99U79f7ShfkYhHY8gEccA82TfPyirx
gkbqbAKLwkCwztk/V7oflWpbxvWUPRJ0bagCkS1QjF/im8ukeR1TucqHNqYaGqak
iLZqKIdJUNzGSdwxCQ6ljeOS5BlpXv+vARDBQwPBBernnrolk7itZ7ATygVfHRUg
YcA7PDc78AhoUZ69PAguM5AitnJ22Wt0aeBKv5WhR8TQ7ia4Wpnn5Dm3MsVHZ9ni
vLNI/CdVLuu2t0pQDfHI7q3487yrF03EAA++HLF61zN/f7KGSlN0L/sSVJhHs8aC
E8vvqOfJ66BaJjOCiQhSAZB9l4LgHH/anOKprHFEiVZ2dgY13LgJxpfiDrMKUjoh
fWJXkK+f4eEOkcshWRz+eY9Sj7moEyytVDtEvqBxgHNvgkhwDR5j0TaEJ+POwSyt
P/Gs0ALmABVvtCjliAHVjJ79vvbDdCVfp6VG2PxtQGYCrUQBC9vjJ42Yck0f9iQ8
BQZA+Y2VAE2KoYlXZqSvKH2GFZUPFEr16Kf/WMDnY5xnuT9mgPAwa6YJQ6AuULt4
SX9et7iuxN669ssgYz80/LKH7wC4SBC2MyeVZ9den/SV9632qqMAws7M0FCKCIlJ
GjNd8Ob6J/dnPb4rcG/PLE80aMrozBO3pE9quhcUleGpm3ZSB4OTWJmhDJG1LEsg
JQtizKges85SN0MnV678MDa+UaSZ9BdZDaFzNmlMwmLhIYxFjf9zPMn4tSjcPZ+q
ilZn35u1F7K30/deIiu19/HazQz+aIue+pXRqDXDHK0XQVlv09xm/ZQoTb3By5TL
2spC6BLJt5LFw0eyxILi+dT1/ttUiDC1n98pGX5X92nbQXMT7QCBigiobWaI/GTG
H7Em3g8nR7Lfa0qy+4zuEecNIBhI2ysLKas5Iq7NpSdgN6agNlYsv4/PyorzZ+U7
i3fDN1BmSK0hzQKddHUs6G5WrYYrWzab9jtMlTsnouaRY95qSFtGWS9yJA3HzTJw
xpPFp2kysgDxE9yX2m8Re0Ezm3mntJzfKXL1B5mpJIGyo6SkbRqj/ZRmhOq67QbI
oOvbCB/UmhScYEpIyTvEoDdxoBVrNJJyfmNpWdehylAyKUw9frQ6mR0upHlaLTDh
Kw/FyikUHcDk4z2DW9ztqlb4rWBFm05SEF3JJnRfUgjga8BZqeof2eMxbrfVTUl7
OvjsQnFo5MlyeyXMoHmuYbNyLZz3Zlum8o28mZZPYxZvZrmxACofbfo8OwA3jJV4
aACxuvMNctom2Yh64KxqJq1idiCn8ajenS1f+TvqhdrekilO24tlEsQt8tNV133A
sroqacbmB5yGWI4vn8+qKXbyWl3L3qqQOQXgfQ913Tbm2rLsqLZYUXhWkhorqnbB
HFVV79BeGO0PWcsPU9C/5pNVfW7n6yuZEbPTFm8uZV/Wd20TODgw58bqUUC4fRqy
UfwX2hulrfMKQRpGCneFwmpeSfnF/k+w+ldyn9kZUYRGvbje8M3u2ciNjwv1tOei
CSidUEs8SPogXcX3js1OGztj7QbSt7g5t2oSiLY4kq0OCFZsRWSgMXQob4B7Mc6P
ga1a51yTnna5TnZBM3Ga/cLifW2kg8tpZOctrNCeNTNLLYpfb02V8Zyvb1JlaZy2
AQcC68eVw4bz75UEkHI6dEy5DRNJLvhPrufHv6DV5xY1/yqOxJaTVn+cb+2Eulnv
JxKIbggBkQI/JW7pkCXeSM3PvETannZcnJ+tVHbyo3ymnA/ROG6PzlyjVaCOSckT
EbvY++3AAI7KA1b5VMYda7EaSky570HBXsLHgurD2WkTNMMep2r6e+3ekP7wnA05
ez8NN8nVs/75765FXRy7bXtip4MxfhnW7UuuxfNqoRZpgGlSS/mrIXstkT8uAjKF
6lhsOo/0chLzvLo1LS/YxMIjYgEY90iJfVEjdvthRkVMXzvcgRJjV5bulONCMeNU
4vJ79VgiYxedwq3E3rUQr27HNKpji4QcP/tjPyMja2c8YxOnipnOgr43yyUX1Uhl
rtlBVLR2rapVXRiWl8ecXVNnC7im6aO71fKNpJE1h4XoyyW4J1JHal0tEP5BHUov
g2aynp83+UySlhPXXYYIPU/2TYnTnCrtFJ/ZXhwOxLMHcjaFyxe5lcwzG+F/2fqS
Cd4kDZil4VQYzYXJQfyZdGhrqSBEKv0S0aLL3wUJ430yRzYttWL32hghmvadB2+i
tDGBhiAipDnk67Q9pfr2pQIYQuPhJ7d+P11XplJfTEFvAgkdVsQJuFQy5XZoGaXZ
BG/2BZeQ371hN6pXf1szEZldJZRhQU1tzNlEZS+sIcZUPezf+oBliMgUy+H+nouN
b2lnt+eQ0toIq/CuZ5tNREucC3ETFTmnquKKneXHsxODbg0yILbd3NXUOzESUWlG
evNRdU34oqlzAdWAJr3UyxRQY6fVadHMwtsI2PkNKGiyP7pWUxWkl1ZFXAzOElQm
APCahpO5HzgougNOr5FsHTkbyzvPwkYIQ9Ree9NyvecveQCKuNDuEv1CES2TU5I1
YfRj6/vFxGzI3a/PRzvItqPUrhaBKp6YUgSVh5acYQMSd7WSz67zjwVMUUkrlhVq
AX+1j2TT8D6XwaQYmiYZ2yRgItdAMOqX8tNLk29dhH/wneFPSnF9eo7mv63P0v44
IBdy7/5iW3zLATxitSbQmVSYfxUj2AEaxQer911Jn0oqag4NMZ5mNF9apdBKLBJD
LrDSjIZpTRCMjV4NqNMsKHXPX2X6NtDk9ig2le/fyKGOyF6/TuMBAhaREynjETj5
SdkK05i1BIGyHEJbFMWylv7M7MA7IsBky3rmeV97BAH0MHW3tBQ3t+B3w6UOYfyo
ALKkEJPWC6UTvvX4cXBcAAaNDr6/dWtOWtBtB09rhqds3EJ6o3d3HM0vUUSzA+Tw
4jpHqoXBHKXIi6E3ertdsNIg74T2HCUi8t37MqiorBxP12A6vT2bhkuu1Xlj8btN
5Y4gR/EcMrpa9Gkn+uEdZrDUjhn4jGimk7tO3n7Ra7uDYwWLkHj0Og27wKGI+EZ+
v7NGyzYyADtY1/bOivOyfOis0OSMVF9rDzrZHGdDaxIcrxq27gQhs8qQM3K5EIbn
EN8VN8ee0qgTUsbpU6YXwlgQKQb9iUlxyAy06ykFMtIUcW5/bpn+RBrMwODzXtHF
j2z45cGNimolMDB7Xk02W56MoQ+MvPavwvti1NPUAPnwZXJ1TxYBFMAKLFGBxLHw
62ka6Rd1teeXPE/QSOtd/0DJWEqtEiFP91ZR6ljrpEHCT9lUykZ+SGr2Mi0tDmS1
xFu3ZjdQkEgrknZvm4BL70GjcEdrZ1zbCnTwKYq7R1XE1WAepT+EsC1bR2e7aFVe
/6cwWYQ260oaMSLv4KdG1BCK7lYxJVOKEO/b1Lu/H80AKtStEJCTH4wncmugZPbg
7b0ctE4T+sSc7VAjQ+C+9l57PtUYL5R6Ho5Vv+3u0zzoWPsOyjyyhGcyH82io/Jn
u8tz0ON9n2j1X5FG5UOVu6KZGuwKbfWc62cjttTIQ9MWKH9i1BhSB0PrK89AK6Gx
JgOkUYXsa0xnHigVQfHeL/riWzW9L7NdyqV5AEa1QwDiyZObaIncI+/aWLybcxA1
YKm2rpvhGVzuq0f+OnxOfAp7pji48bhWhjCQfnNfo3Ty6u8YB5qxCGaPCg4gUkJr
TSBONjkT+U0fDtsbs8uBjIg3nUaO78pjme8Fjj+NICHVeutL//RbrwVEzY0bs3t2
e+rQiSso2E+g5CfHZQpP2GhI6O3GjYFFQdKoHcWsOt7msfwQdkcRzj82n6zNhUen
peEjz2cySfj2mvY482+FZipmH9lGtWG9b7yqBGJPq07yBVZbREAdtANTWFo0LF0W
XK/P30dMz09X/Zaa2t9wQxikuWWXkVyndSoDs2n39wTajVibGNEeo9pYOeQGzJfM
iFxBVdwMWm/6stjd+n7hMxJZkiRd29gFWlJDRBv3cQwdRSG42EV0spHjy/thCpdx
CzpBJHwE51S4cmWjNCCdXjC2WAZzJOEoVIIFtkMPj4NUdD1XAD52hndAjgAgUoN7
OazwCRNu0kwQ+hkO9wZYqtMPzBB5dHUAVKPSn97J8pR2VESw7rvGryAp9BrXsmUq
NaiGJSJNcu8RqFyqgk7tZAkDiALzDPrmBV1egzMpM6gKbgIA0HLAQNG2XKwexR+h
KQKZYYM/owCcMv7c66lPzOmkEe3weuAwsyheokMIEmt6dPmx0tTjVuFPvTWTBBVO
LUJvPpSHF8lpz1d0xK1ddvNAF1T062sqgXGkAQmOw9XHa2XQ3nQoZEpO7qPlDJMC
OgKEWutncvRGrZsBya1aKx6vWxkpyCmdTX+BSU5N6SpttBDZdXO1hZ5nknM0Na3O
cuPLVQnAgqhS/YKiWaXGe9TMTGKuqlKbcGZjeevGcWIvfMrgJcGa3V8AokigrHRc
yz32OEU9zN8KyjCpBxI6vAxwszClIihbEBVewEEfDSpANGzKj+XGyU5wIUso7wGY
KYFVmytqYsFozTF2zlRTfffu6WYn31Ab//05aef7GyvizAATxES7G3P+r6dsIMM4
m3XMTXqMnv7xsBXAorHlQ8BZ5xs3XmdhC9wPbUS2BugKgCdsIx2qnm1JDmOwr1t7
8ZuHLTDHM8fM1ydhw8BKtGAmaiTkS3v8IcQGDUjf97iVZqLKVq4r5GmOFZ/89MwY
CNVf1bjC3yiJz0Gy7VBKZXLGLJsUiAcGK3ifnKrqkmg+YFo2UOdvU43xLrJzVlEX
JD0ZBdTlKnr50oC2DAN5ObeAyerKSPBvwPgCAmX4BGKScepOlz6fBjhOAC1BeF6v
6+z6Mq9q4sEbQKEERHr5Dols0tG56Zj1jAikKpAX6N3Z1oyr6keiVGB4x3I2TT3k
WS2Y0nj/NRjfpmyWa5wCKkmhRyP93tL97MQ2crpuj4lmLgu9n6jrVUmEiwK6zBgn
++7s2zkzDmXNXsJjgC7FWx8mSosjUg407KY7urvGslqZlOQNa8Deix5c5AfZ43cV
X2FtvU+2ayb8JKusuPLwETZ7MH+YgrbeoLv5f1cIALs6W3j/isVcIY0rmlJ2g+kt
8xVv/qekrOy5VMDwaFU+WN2SmWYyoyDiNBso9N9DahFTN3erCfZoohGF5UoqFf6N
2z/CCbvf8YhigPZBBaAt8HUvXQNlMxiz5fJc5Im6EwqoYecdnUY+iUXuEu2GNI39
dEUvjJUKbrHuXxOWAo04KsMiKb1Ll9i5YMq6QqPYjipl6zgX0pAsbyZTKvjp3jum
yjuvm7rWZVR6U3rlPpf1c+FpSgs4sPVjmBmvWiVKPaW55mqdzw5gDinhXMUmomC5
c6sBLBa2uqp/BNuRyxMlPUnKNAcVLTlpBdxzc84bPPVAd1vm7eCiiNhIO7fx6uZN
vYIvqXP7j12qtAhZ8ct/M87NPdzGLJebAbFSDOIhP6eiY+o97li/fVvv7JDMvdQC
4KVYTtZwwtRdi7Cqy/Qnjk6OB1v0FkgTmCxDbpW2dbU4IMP3502WpdKvxSGvEaLo
oJKW6QUATtYPMQ4/d4revTEsm+KQ0Fr4Qq5z6HiDxTo0QFt45XW8Ht3RgMpl33vk
a7HuoSDyA8/QAOwOjL5k/rsp9bqC5Knn7iBxEkQCiEFisB2gylNkz44TEfB8M0q+
j0kVTsvrZy2Q3NQx+wEXydlMQYB0qloOtpzCG0yKNEbvASkki3cYinoJbJ5yzzvR
SHF632vsQjLMOtIdfVdkFijHZoDXE3aKrfY4iFeGiokjsdU4OyQs7KyO3aZa08tO
1lcZVMO0ZDg6GwHBa2Pf5EHUTz0aYlkuvbibFRkHmLJTCCZWtlQ8+IDc1AQMyVNZ
AgqS9UeevYRkA5hKTpL5EaAeouwr7XsX46lXmjTYhAoU14u88Gpla9geXtEHwAH7
EJK9MVOC/wrC1LlmDpLda0K7s4OQS8cBzsLbAMo0e3lIH/zZIibxEvEG7BfK3rkf
EIkuBgyY9eZkUQbR/SRpzPUr9y+itHXQfykiaqyIpJJngsGGHSfP4OO6MHTkowYO
yrV29jRH9mq3wlkNfbTbzaPQScDN1WP0wxCW5+pjuWCIZnYlE+XzRhor71DdqkNL
8t2+bHUBFoY1RNIB4ix+/yXuBHCwmqk+OlHuGnKG9w6do0QqzDKl7kKdJQbSGpCa
VHDR6YpqMa5nIdqw9YwZHYBz9GlEzIjWe3Nb6l8YMnI8VBIUC4hNK4wVuCxARB/2
Oqv/1sc4r2DFrcrON2pLfjQ9FiXOVFCcWSWwe8rqacqRCnZwrlhZTqGGETlDOw0L
zXTJJQDWs1lMhqd6KO1or7wJY7alfsSXMcrTK2HCPb2ObrW9LabDqjWLbQ1/D+f6
1m6NypImGdNbZGHsxQV3oX3NLn85fhlofzCzlKS978CCvq6pDAXNq2MwEJT06jQY
gppFrrUyGWkZpcYiuBNuPtT5JeGltTd3C+Gn2X6O5Vgc1v5HeKzlclvUsvy/75Ff
IeveOgA5kefe90lo/TY5mZZUvhNDyiHBuzfoyOZ3t7fFC4AUbgRw38ytyCgySR62
2TyNyM+wS8fH0LLv7P7N7F4CwMUK+2KXtrsccR2tfsuGgt+ZQfpArh80yl16QV4i
pc7sJQ5tL7hIoppts0RxvyRYfwRUYAnN3MbdvHkjAVHPFVDDAaN6qUVmnx9l7wHC
PR09fY8cxox9yNHJC7GjEPJ9A4Vyb01uzN8e6Mstmsuxzi06OVaFCF9Bue5CGCb6
L7rtBbDwWT05uRT+LIDFWSTtep0Ddh0++jk0NRSkbdKG7UFsHzQpffyOA7QifbFh
OFSid6Mw5CEhDzhOd0Ri7GwvMDsBn9iiCRpKAVPDAEJTjPbWwX36sXZXcak3Dgo+
OqjWaf8cCQJLMQb+JfLzXU4dR6+sFiRNfjFOD1OuHWP/W9yOxl4XtXI4LDIuUky8
Swku7cUDylcSb+EQCiVkUaVJdmElX1N9/bjaGt4RUsKVzwzQchV88CG6jSuS9ZDi
MreKFk/JHqo9+YrtVQ9P9rVShdQ1kR5jmz3HlUKZiBnlLLDx5vXmIgq4G1hO4b2n
fQ/YGt7TCInbNEAvOqQEsG7R4vNgAhl0syr5GBu13rcekYhCorri7wQyLrG0oRpz
wqso1i9cvON4JjpKWU9PDBfKsdnNn8nueu9jbn2TwmHyM7rq3lw0V+7FvydI3ur3
G2Kfr+RYrWpgO13+1TfcrK0KvbsgDRx1lujSmxzPq+OrbLPVFhzFSKfZo4hvgudI
qDGqPINUWYarov2LofG3B3whSIrzMrVjgGhYuYD2zV4Hb5t0EbzkwohciGfhDWhi
2/NxXxtpAj+OS4OuuqqBeHXvsDzU9PR2SkWk82o6NMC74qbzvWUDcNCiNiL9xq8p
STztzx2BCcYSaMno4CiycaKgycGW/EtdEoL9Y/4r5xuoqm7L70g7KQDWUDfZjLDY
pPdznNMxewPQuZ6hn9DugU11H6HQbR7jZwbai8PFrFs4Y8WoWiqIxPYg4S5AjfbV
ilReU8683ar4YnREUty1egPl3B8wYkLV74yShX3MfzZP1fydFhbfaaIuuIl9T/eV
qxToygiYn+gdFAdIcWGKMDV6Iz1dRvdtFnvbQTkt7YGQl5oFd5bacxSsfB7p9cTW
a8Z3s7yT8mfYxN1t1RK4e6kXa+dK7vs7S791XabUXD84+iHHwBmbveZwJ3yLz7yP
p2q8S9V8EFKwshKRvDmYeL5hyB34BaTB5xqyoUmIxSp6MLffge3zRLo+uJyWUqy4
RvFWljPryAkgUUyP6cUHuIYkOmKyRKnNAWVFqETKjJFatllgOnGXla7JZKkF43/E
xCim13fkKuIW9ycH98TMlsXpImHOmWn8SpAA+myfMCobcZ/xIXKuc02lVBITCGwP
hu6xWZvtVTuToxTVTdk5OUwWXIwXr2wUAyDzK6rIe34qAWIJa0QLwaa58E+H+Ykc
eR1KpiCmcYngj/mK/nPU5WfEIGydEiY3SDMsFShrgiI0drdvjdfWHU10gLHmNrNF
kOdPaDpIXE6/2PdVXO9RmkXHyJAOgkm23jPAQiYnluuqbYxIioaWMlIWvMeGZLrw
qHBUqT8b5ePIzuT2J3TP+n0A9CaSn2mhABsSKCV4iQoh7f4a+JZ2hMoKYa8/JDSl
zw80AcaULsJKcmY0bzjtk0bHIyWULbgH5xYwFzlvRZuuWZ1gnqVihcNujEhZH+5N
e45+iPKD6sMcraae0R2HklxZm6e06TE4tlrHbMIFa6yLbLOuEwIR1WGnFRkOkOEe
GiZMgJFUEc1bXX7tJSv1WMDC5e/UNOfrL0Lq9I7ytbg/huX0tzZw3+MktziDWyw3
6V3jiwn3TIEUoiU6z2h9NvtgOOGs2jT+a59crY7+8XPW6RneySAt2U8D4eN6saeh
8sohziTJljdNVEmxUXOG2pW5oIUmOewaeZg3eHKz2rXnoSCOyzI8qoQzWcudVcmC
lsAAty3LOWklXN4aTp3ad7wZFWAMSQh9shAa5AK+xZZicom6JF1Kw9oYUSlJ+781
4HKXzi6WPwh2OJIBW9Fgkf3CBKa0RTgo7dplTyazE1A5WBVlIFG07jXrxI92z3va
DLtakkedas1O5jhxX8BRxJHa/7oQfApOQTlOmSMVKsvHpCZ8mPVB00EeNCsxuNbZ
TtjJeI+cLhe3YlaTHNWr+DsqJfdrCKWj+wCGnBjsPqHatdq5pOyRHU6QktUz1+Gq
LfEJPB6eiujvJKDaBI/+/7h4q2szFO5AeoeZVywW06WDSppqY+rIuRheDO9VwcfV
ucDZIw58d4ljYEED3B/emCy6oKuNCD5kV/5qrMngFjdrZOBBdTB+9+HXFdaZiebS
DNZCrBXi6LdNJlwkJm5IaOMDs+Cf2YOAaHNYH4p4mo8jmC7Nyo1i7aMFUzlCLQ8T
MOY3T0Ze9S4z7bl5xjHlcc1ZW9QbWdyvf2QXfSxswA7q5BbEZtIfnDMhawKhaW79
lUW6YX7lQnK/Wthpzqbde9akD0s6/mGyU6WghCfxGs9LODIDRm0BqkTxjSf3H3ek
S2VZ9KN3FEW2F5dgwRKuc5LBdTo4IyMPbRvmmX8rZJray9RARhrhqiO2ECnbBd19
TzYF/uL2fLewGroZsrcWxUnEXqYKIH76jHzKhICgIShvCrKWQeAFHe5IMQo5krbd
82jK51zO0+cug8Ql80CTMeb7hbTMpEI8cPyTESk1FElniQ6vZ2gSMNT16hR1jVuW
Jjb1e9jP3HBSWBNiqnTgz3Gxs364q8Jg3sB5ZnG3OGopS/bQqlYN0DRoH5pVQBWA
tqUf/35IacjApOYlDMnQ8nE4H24bt9JT9Tc9kZXPnzJGMgQC2Vo6Ma5WVQ9sEK+j
qUU38UPOOuffQIYDL7cP9SEPBHPGFdldlCsoxKMVxMmB8QOqrc4Bp3WRlUxA2PlZ
OwukVdmBT2OROJmCrbOZ8V+p7JXEcD4+48zv3hmYvWcPGozt4BZHxaA3qh2Ju+eu
a8SJr+LwFTysIuyWuWsk9UMe2cD00d8mVE1G2EzzkbeTPc4l1KQz/ePMr575zGLN
mbXNW9UNoIK3LbUS8l2EuwQaCkPIEHc1Zn2pdJAJhWHC12It85hkRvZdmEme/DNq
p9In3xd5kfaGlLu+TjTjTWCCuq2d+NII9U9TgpJMWx3JITmwrBoCjZZ1s+AskRpH
S/rIcmhnh/PvxOQl7nxVA1BAqEJGllIxJfyC5QmYedzkBalHqoTkzYSCp8ztgyQt
qtm0e51+Zag14plWAFuf5gJhkmMrDDmXPhiOzt68Srlxn9JmprfRDJi+Jg+8jI6K
wqmIN3kAVxB4TdqPI1P3J6NZVmt5XrAg8547qj2QWtFVM+fOGeJ0hyoQfJ4rL9+0
Z13LKEgA7H41W09+U8TuHnPtNzoroffgOcusqIkTiVLAeU77PVRybhojyRcVBLMw
MjIqszrd2eF4ARF1ZAGvdnfOlK6j0uNtcbBHHJTQE3x5Jds5++TOcrST6B49cZ9J
FbYRc1/V0jgf8lrWHvQ34hKBtyaSTfdnogYe47KC8jjlSsrm8faG6iZoGogWZzv0
/Q1jbpt6d2YXoTDhnNtigpBS9c2vGaIZcpgBfyEt3rsgtNQG3WfTURWaLm4GN4oa
BPlqnzqdTlfvJOht3ekzVI6FBFN7yyz156WxJv/78cFYcjeR9pUiNrne7E76kYCs
9JCjfXnBzJHN76Z1GZa+FKRKmb6qMg0koBSADqwNPadytoOVMhXIc+xecbmANV2g
vPXvZUlw+7aIWd19KAYub4+VYBnnvC3hJAmKl2Py1WrKCngiemJF63Py4UnZ+7Pw
r9GUfq+/W50ZKji+nZvcr9+PVbJALjIV8x0yhBdG2TZkvFnitfe52pyTWB/Yj6cP
qVpGGd0ERpgNqbZlbTy3h9s3x+V1tdwC12MVH2m0Ndhqfs0RGuWsjTvGrzR1Zrvx
AZI83jIPRga20jqmoao30OMxMSQs9O/aDCw1JfR1jBvLSVycinn/bX1Az0HSKn/H
G5gAxcb8GzeqXYra63zpTZnL3s1XOLwN6Qhy7ng37O8+ZBzCMHpK0RtG9qWHwEix
bGlVxog/7K9XneztaV+HMdoRL8+kOaFX3bHudpXJ6fpGuAeswqXO4S+iDhed4tnQ
zFT/hZXrcuTGOeQNa8FZ8QlSVST0m+3PNmeEeZPFIl6ZikGdUEwmNdJKQX4/xLff
2p09HOR4tIXkw0hN7YUQqy/vBIsAKbuyvSnzJ3E0rn3DojbNp8YWr7bb3lb3kJ0+
DpDoYMgf0Dcs+PI4HJnb1WovnNhlGrKSzCdqL+7XCffcZBuVu/1I0p+kjg0T/B68
hR1LKOe+L9I4cTXMUxV9MGodNNInPNxCELHr0I6nHv2vswLrIy2gAdGCxCGXiJS8
/UMCSS5eqPhok8LlJu4ZcUoPdiNwm8WKPMJ+ZyuTPN3tGQEkKVaw+UslPQUm7dhj
B7Nj4Gf0VJ1VhLhl5m5kDJjIIb70FmP9pF900Vpngg0KKkW5HsttS1/gg4iTjQQT
2QsKMIA382RDrkiZVnsUOrLN1NI98IlrM27KO/lIJQ8/nwhnIhRmCnaExl1G2P8P
BsoarDkO9SPitWY2f9N/8VTT2Rg59opZBdXH6ymxHLw8JZhtdvaRbsNUs/WTKGXj
TUXnmzs5Fz+O4fe9QBNWZYabCMTVI2gE2UQmthlvPQtWubyKKadPidVQj3/e+Mo7
PX3cLOFc7e2FAbbTVBUItEcQ76d5/Op8eg8iDpPi+YwKLoFogH/gkLDMk85tecEp
jLuJvU2d+xSJZGfks653vIeTV+AYiGGPAwvqSuXBz2kcvBQOTs5cAJ4ZIhgpWMO8
3oH3RgegPRhINKA7SSie2iVKEWrzBVzizcrD+8xjf4ME2d/q7dCR6xSJKa4q3OKU
haga6uGuGa/gZ/+AGppyTb/6Uwgl4afHodemCP+BuJ8YOe3ga560P5LD83Xfp9H1
sEvGr8EMOxIW4yOdpfPEDnyTllAWoBLsv2Ht9QDxNVxUyxS1fOW0D2KJmvrbQR6g
cZC5Na2pitfnVWVZgKpVmuvYrPWZg5S7V9JV5pzyxRlPY7JdQ9AXxKOmz2qZgRxn
2kNGpe8fdbFk16pQIutV1YLeUAe+6bJ7RKMzew1M6GEdf3qyqXxvx/8qMZsQydEK
pw3rK+SsMaxVGc2SNcXsZ9pk6qddu9Z+bet8q5vS5CBAnVryN2Rzysabi7nnUXGe
i2+r5XOQVZmMHzStY9EiqmIkXxrt8EkttFZ54bUopRvTGzBZ22tFL7trxRnAloYB
zrgzn56JMfMRSIUa1Wi8wK5m0taW3Zwhb8IGHu2usn75uSxnZjrKe5x+H1zp7B/E
AKRDbOPCbHyPA8ICJn7qILP34gZLKLsU60rGLnw1KuhZRlG4DL4CSD2nOhfpgAgH
MclhSQggoUPExpf/Hm5EOKh9gTgUG8y+7ufiR9s5FUwgN2ZPYk73QYKAdCnMfQao
KTC1m86lpPXU81Ntp4teILEewn1Jyd5tglEegDF5exgSRIo4IAP/B+vFB5mIsOZj
OtsFRfo6b4mrlp2Ce2wocoqvAxlEtGCeEirjjt6e/XCwSWAXQAQrfyUUlQWcyf45
7r4MZ7rByl8Veo2vg5KMCi5kUGxpzPH/xKKzS+ygsk3uvW3Izx1kYVDFJsGqEL1u
HgXd+0lJ0nCD+nQ409Xm6zBUKtYOHWT1QDZ8kRQKT3DUQarKOoKw2uU8eRPu8hGk
GBjEQ+7nmWMfOzD1/9o0AYdrfAO92boSVdx4VpoW7vFbrdCUtZOiQQVMm7dgKIxo
jmStd+NJt+YUy8jrc1Tny3f4ZZwlkAKlNdOLjHGaGKSNdEKMgY1BK92RS3+jRBOR
bEB5quRD7CrUdiPhIwnPn9+fYDVaAr7pk7QHlINre3GrGGLalaoOPBqgGHnhH9xL
O+1zmuZa3F+C78d0QHhSIsTcEMGMbvPD+4mTh7fC+wOUinGg4aag0/Kr6axqnRyk
iNXvODUOPNBQDW56ElVq+NrD9NU4m7Fe+t1BuXVLh0oVzaJPwdGauSNBVmuFkYbM
NejSnh70hoj7cV4w6IQlgPs+CLQUsvRnR1HBOrfJ5T5971MKNzPPTLvIHJcGpzuq
hQRBRXrDEUpw0LvGntAz46hj/UtpJOGxnqGXcwMnKIECHivhaVnkcDyU0UUCNHsb
NIYovqndv2KdVasLpnfKLbsvB0lk00sTiQPJdjqiNJ6POFMWTl/bWtCT5lQCMnYQ
14vQCwQKIa+D17DCylbSk4ZozoFMch4Mv12TRB1PwM5+xvMsGNAfdNJ36amtc31Y
oSi3/pbEa9n7Qkqt6McckxqAOPXx1cRl4w8hdmqF6hK28ofJgqEsVQ6Lg58R8u4i
rztUQtn+yH8Lb8LOFfbFxjVgVlhOr19CDL5bov2qHR0fVs9rLENuqYqMAOcMPxdS
bMsYvUdZUlZMDm94uDcG3tjat66jlqVi4VtaJdW4TCnLrZoKrB1xBXSA7bLM/3Lt
B9INNxlA++y/KnKTExpELV8wnVlyp8WLVm6+XCG4U0/igVcnP9plnKuB+NuB3JvW
DxF76VDAtalaqVBXTSAR0/aYXNJsFV3zBbaPJGoEAOTHftpq7ghibWUIBGZ90k/y
kMAQQh7W2XRh+L87Z0+AyCb76csdMexceTsqHqh9vP3ohOVHwup/7g4W/uTu2+9V
TFD7EgE9+j2WcMkG8ROjd8ZDDKxHOc+KZbP1NsmoABUB39OPs5Q87f86uM4bEvd0
CgaLG9e0YYUQKkGJ9+8nlD6WQ6aBFHG/QeyvpJS99TQnh9DiJwXsqz9mcG3Ywvav
qN3yd6NRAj597WOKkfforQ4WkFLVCOhP2Or6WskH7sXentFH8pBbAY8O0XGpqjmm
6kqt1cncMrlxcA6dTSXC+AbzcGvtx31ZiqhxIgPxNW83kCVFa1LZtv9ldVd1ZGfx
O1CMXDc8Cat5JXWbijsYBIlH+oo37rhDMCBShqxtxe0FI1n/QJcLL578iCnsukXp
awM0J3Dr4YkfonDTHGUD7uUy593w9cR9YoM9aVdUPjxmdxVD4m3wTml2n9bYnL1x
P/M6xYcH5HHXWbO65qI+7XzcZ1w/t51AU2ttb2LWcTFkbro0g+MSPVNNNmCCmPo6
RkNAvZUuO+5pWvZqoJ2IzulBQUiVnKTAF3osPU7cNdlKnkZ/aV4u47+/yxnJdXKv
TYHAVFlOR4CJR8JaCu0HRFL1X20pfwk4TsaKo1wQmJ/a9WeKyW6BMd1TP+H7i6DW
BFkSOgVET94hlDYnil+qxzeEM44VY8oZINuKTDEooV7x90HKV5tPAP02PGe9ywD9
7hH14VU/OR2MWa64/arEZDrIv6kf8HELz5B9XgaYJPdLb1YXvG65J1yTuwPTGqtc
UKixziT3kOmHsYvgVvmxmOl7fzH6AER2OJHSDZHzr/r3fW84PWvyAyF3Fg8dZ84X
hxFI95ItUM/mhdxPnOLty3FSz3WwNrEt/+5QMDqn/hF6vyWFju7AGsfVgkMEG9VQ
IYVTfGMUCWTCTUmUdPRGEiYz4466IXAKmvW/8lDldQq6tqmfyuXHWkWYTUUQWCEt
APc61odi3lJ9yoht251tNtcexnBE+jefwtudGtOEDjqxtLix6YmEGQzGWFsj7NwJ
UlPbBD0/Djlh+tBnQB3k4eEPlXl95CPIHAdfEW6lwgA2hQOU3BQwjQvtiLD8XRUJ
r+sKfHbjxR7WsQYsTc1UAdkPvK/KUug1P1jSVvEFK5I3AYfrSrX1t0VKbNBRXCfH
hPRt2Smn3IjCigQZzXayHTBg/J9Zgs8hQe5NI/EYe5GUD/uKV5JG0LQTK58EUuMp
SQbBQazz5/XfMwLtI+32jAaGcYF5q5A+pNeeynDinrX9AVP3XwI9OO18A6Lu7NhU
725eWuvWV4DBkshWJKRCdVK3KxU1qYNhh8faKk5K7d5cGaVFIfFDkHfvBIg8a+dy
GjPpX1I96Nc3rvxmvFfGCs01ZYGWU/733pcLQtPIT+P1oUHo++gIegpMIPHd/yqM
mCSpVURxRC1WHEHYS6NyrzaSSYKpbIpf4EPPZi5fNPhoOkMOndcdz1tfge3XPGyl
zUbzaugi+/i+Rhy/woBq0rN0fFn42w4QpAgTUF4sbSGGqX6kNRZr0xfhl2X5ZQJ+
EgtkpI0vDpY5Kv/hWk58us+2vH52Ft7Tu1BNPdGnw1Qe90JPymCNgCwQ474p/80g
XPMS7xm+0GPf7zFzOqCxSKwkYyH1oUEB/8/x5rFc7JfDo2K5nEGPABc6abuI7WTz
saTAz1YD1Db36u157QvU1A0MK8mfC5GXf5aHnPWMwpVSVforsDoUO0vEIWzY6+Xd
WBBML3iOMGXOlmqtT6b8Q/yY4NiFyOFFNP5SszWHP4lsCBxrpCVzlZ2EOIJLRqYf
5/49i/shOg8eySUjXXr2p/X1L4jFt3Mg7qRLMRc4nMX+fxj1EhSkt+hs3EwOOdAm
fV7vEAI35/yZieCjJfs/jI2Tk8P+jde3/FAONLNw+VledYpuczuArFs2NkIsJQ/k
UO9VisjTZkYuPJG6qlAbrVq2RgtKmieonnqGnZARvgLvEYh0Z+nGFu+Muaz9pmaB
CMHxDLNUHbjJigAFz3vDSw65u8NHMkoVK6rrLHhYJzMpeUTHDld0AdD4UzBk5fw3
OfbXw8FrTPXRBE//w8B/fa02+B13u7YtcTy4hcvgoxCm7Pn5F6Kyyl75yIZuhtzY
3R8e68oBZcYGRL3SJh/tHBedn0QH+QlV00+3juDGOrcasSVwNlVkYxhCKjeequ0/
QwqU2xqGSOrh+DkWNERGqf7UvrACShU9H8/wLiXF6bpDtoGiVyi4Ype9ZlbrI8n8
6i0NNSHp9b4krYX1MzIQF1EjQVEIH+UmxqPhetwUI23JNe21tzXWnkNHaLRK4iru
EFAsKxECvL5xJzqaHtuyigFWp18jptt4E6lt5lpfsOti7HmnobKddyhaypn9hds0
JwjEMrjgT4JXO5Ky+3j5uX6JTl41T+5yuvxv0L9rwNdOglaEV6OoAQJAEKelfYOC
qu7SHIvrqCzXB62u+rHRX2wjkeiYOpBQ3PAJNfwYa/fS+PaLsdkXot9wSm2SmQfg
vi6+p01xAKbpKJp000krrhaOObrPLVDfsowV2g7NJnI5YSqXeRYIbRdggOyQtp/v
npAstzl8XmnmEp7SPGq6pz1PIvQaIRduPxwENx9rVzcoG7MJerAyWpWMFO4Ow0H5
0aj8AhVdprPdwzxC+6uRk38hGeHNW5aLNYYZaI0Y+W9AdDWQcGBpTwNvJ3hYqHby
39cFjARzTLfT29lKGiaVwUL8hvdaOQW9WSwCHbHjk1/ns//2ILGIENE16liTEOO7
qFT/e9XWO9CAcIALVKLAhK3Ee7sEYNY7ga/cDwDmeugOFno98ArvlZUr7gyE7+bj
dZOCk6VKo3pYvcCppPfTRv9rBtT7Lhy9tbfd1T0NHhi6yHEnkIBkOg4lAQH+afay
HguWmTPm9WpOK70A5MET5w619RxRFWYAABDa4JEG1i4XZ708NZkCz1apRpkEYfjU
qX2cvtoaPksadjZhseV2a1JRvg+ywiPn2hpTqqJk/QlwTaHG0w5/bTTkDuQNgIEJ
6qhfs0fetTbVFk2SvdtL3iXS67umBaW/zpmxG6AJ2Bu9xdADMHkm0YcrhIfAXwHI
+EYGaXmp3hgImDGuTaNr/Nrjcg3v13AcISFmUAeQYHSjmKEZKzk2SMmnSc32zHy6
vF4ClZceoSYqcluCuXaIeFhwoe3RMTN1VG59AZ2dD/rQ1E3jO6TBY7K5G6ttFTRO
Hh2kGVpPDOltTH6MPqMYxb1+SZmupn+yVn4nGaCketZQKGKvZfMr6RoilWtytrgd
CzxHqe0KmyyakE1sMbwBp6u+dceP23GqMYasj3/Pem1UeweO3wh9d29caK/rHLWO
DoNUPSjPV+nViEtSjWIhQgr2gBlSdHr+MHV40HWbXgj2v0PT8Fkxi7dbhqKplzeV
LCkUOSYLKHfmQTT1vu4HJSdpYOCIUgdBWrfeFyY9sHsnTEd8D8nwQwnOI961I+2h
7aE2QB+MwBl7NiehTkoNm4uLq5wD9YIR35PKMVoRz4uG3Hfcu3wBJrvHvPvvAAJk
ik93JV9+EE6jbnhv9seYrDE8AKzj9K+EO2otqUhrRum0BoQe6wUZdfXNRxK6046i
J+X/Yz0+ybpkym08QkKRp86vuNNcQmw5Wdf1chnOBzzicwiQ00tGi70z8PWz3Dv+
P49PTHcj6RJe2az2l7HUy/3O6FwBOhjuO9I+J4KKod/4EM8RmwqjPRoz1aphVIrq
wNGHwuenpnqdtB4bfVftxO4Kyvt651DfKPntuxqmydFCLYfIGgPvhPtSj87zUB0Y
FA7OkRJCiMgav7yDajgjmpgfcksZn6GbYKad9xNyCMbHeU5lH1tQcm+x5r1Xo07F
M9h1F6V0WVQBxw9LIz1NcqrWyn8KQZD/jIeqVbp05kjbyNrQM99ZeolsMUEDHdnW
0KsxMogsG5Ce1dxPYsGfvnQ9oUQ0jNp5qzTcFziOCLP74MZNyxHaPYCMGboeqYBV
QO9PiRhyJlTDPLWyxQYmtsrbzhIdBhEgBHwn2EZqGxY/xMFucw3NYIrlQyFzHA0o
vPK7r2Uocn1LVu/wP16Qw6rDDamkhrnJRBuxGo8Jxczuhj9+Db6Da1WEXYARPksP
F7wZVRGdluVbztam1jvvy/pbSPYcd/NfVLevfYkQxfLdBx9WdMbDPPvFTShPiaAG
7bp5NZuoSEordzJCkchpPnLosGRDca9rI928wLzjwTA+gw2L+hLx0wvGZM6FbLMW
2Y0uwiAc1Ht1cuxxtK/YmPqfi6F2PHC+kOY+zv3tD3T9KrypARPvK9jyxYYQZoF3
42RdxmFnDMCgvifirE1/ScCK71SAQ5r1USW+XcylmIMeDA35+LifYIWuucCZ8WP7
uiLUy7c1TC2XSuRi5jGO/5H8FomalfTmhQKHULa9ltvXo/QTqPcreR3sap3Mh4dt
ara6iA8eQPcBOS0OK7ajocgzXHF7wyOH47kDrZUiildgTVGdkbhngQU12+i7/if/
VX3yO4wRFkDTlPvUS2SDAwcE7jtsXy0bvdi45WxBZ+oz8s0p2ljKNQic7TUAEtwm
JS8wo/ZvKosazej7FpWevdg6w/xdya3h4Od6C8hhz+dHQGeHY9jzupN1IhIlvXW7
dX4EKOm5HGu61X31SiUetDbG0xOJIGmDjodoYpDrpWj0TO2vbjYhLIOblBF+ZlD+
hhj6fCp4KG3NJURDt1W1/NENW3DzIMsGeTNra/XJabShXHkEhP9lsB9rqAHQgruz
PRMQrecHpDIDGxVli2YA6D+E9ftC3HfHRlYIG2DaLm3eiPin05v3HYbV9qDZUCSj
9i2TX1wWDkjwsWHoT5WT5B2Hs3u+Uo7RdGZDrnLGTU1HCZId/YTkbgt1pwofx6J5
Izd2dpKrjCXrB2tYA4WR9TuVlffJ50sZVJPwyyMV6mPMr8Vqdm+8v0MA37KmVb6R
W6kQCGhL8xIEsZePmN8VLEuoHRK7q6yDQSfDlu3ZiKh0TdAES6hxPNavC1ZyvPA3
lcJ+nJIS8pzQV+qqF0pQbaEqhD1OXvaE7U8FxyHXa6p1lx5SlrzFFVI/u1SM6ACW
cZEYcMl+skRWaWueoGWORg3HoL78q6+2OkDeeIEBRawdA0WsUKjmbzpCPMDOBHhI
DaI9C/uM7x5qOWHlzMaEnlKr3jWJl2YWTMZgzfjvycl+sfps8dRn+qgnmEcTUxfM
xwRLPFSFfc6cqBxok7tElMYOdQPDRCl1j5cthoQ737Q9i2cFGZ7Bl7y29/dRIPeo
vu6SVZNYxLSmxAuvaEehU4ptS5jWVliOhzpXT4lIBeVhv1E5cbwOZt/a16cUXman
0WmmMeHNg1qawzrgtZs7DIQ8xYH7XTBlDPlVKdEvJHOuU7cgqx328h4xKckBetyp
tbQtjCbcQHh+0tD4jS8R8leVwEuKs9+Y7YR9a3sM5MVFL0+Ifg4g/XUYzSJvUQEp
sIeV2bQVNFdQ7SafZ7cIakaZFzlHQS8dPrYG5Bb5+6E5NvF21PTimDPnRBsrPpoM
s/WJtty3ALJ0qm61OrmdoN3Ty0QDBTwTELUf0ACTWCwx65NkWFFcbfGrVCmw7FzY
vnrJId9reStAVHIuy7IAH4Hp5dcxzNvSuvqUrbmHXVkWytSmRX8VNhrjmMVjCf37
oRzZFOrDAm8/1zAc6K3G/4C9wpoYMzmrG8bcnTW7MVtaYPoEVH/+NkeQSsgPl/7f
x/5bC6QfLHe/QNwNbtPkCBItUnzyouAJiCS42Z7r4l1IWjLoET35bf1ARTxKciQU
lKFF0ZeBgN0E4PiDqlPMI//x9wFv/4tlKkdybXxeyW3K9GUXLN5SrUmNQnfIQnqM
ZQ65ae9fKu9aQEyQe4k75dN/sheptsTafzhcxmaXE4DHXLPV97UoONDF36ejkQRJ
owugQbWq7Kpo3d4oQDJQpi9WyGVo77IVidft05dKtqmIPHL6GrZtOuppKvEDsypL
rmB3Y/JxvxGYJRyMbop5emjMA9VVL2nYxb4bB4RdIqNFlyZkv2uZKXS9vGhT58el
ThbPoDYQbGoKJy2I2p1qVby05v/b1eht5SaHBAKDoA6M4j/RyqxsNfY3VTTH0zO0
bjo5CmxIQYxO1DqKyOFllxz4nNLDxE070WrVKZEEtPESWBikfC3U4ry8h1fIkSD0
O6JjcyzC0DT5YTwQCHWtQ3K/QhzMSgK4KkMhmxLtC7ZdbJnLMtnd5KfnSRcMQVcI
bwt873wE2AU3/MRnVSy1JBCWgiPD24moU4fSJpwwJX+CENsSsibkKATfmVeZnJ/R
1NpGAZQS1OCQoK82AtHEDM+WAlC4IT1sJMddD1INW5Rvml/r6hJdxzelSLkP+HNX
T1LGdXeCAhJSIlGJsS0DI9WAXrnPKKIvBSWzod6SaBTK+Bjqo95k+eqYaqdE1xuL
BLabE/+/qx9cVdOpyz0oMXtokDqORlUrX0W3Luk4wKbIDOBr39qruPTYDFeIk4YM
imSMvYJDgaIGFHw1GuwDnI+pvXm8Wks6RzS1JF8mOE0MA1zWZkRnpBXALhYK6Ax6
1NPy8TK6crRe6sEM8yl59lyS/YhxdiVWiL3w8oEKz006xR4deMixy8I8QVX22ChL
Dv2LJhjIaMwmRj0lY4mzfg8aNLWwqAOgy1ULsyP+wFZCD9y0iJjVILvhOGJvEEMm
KDeH2ZPaotrQ+yXl2oD7Td8OrizIIw9ahXiu+q0/DzZ3NAwawIuu8eqA0Y4UL+Oe
Z3FJnt2jCfIICiHiCXTNlA7bFsMMQfLAoWV8mLbbUqR9v4Ts6XIwh/7NhiyyFE2q
nwwQyz+eRi5K5tgEN5afZS16N/L2II4bnyCYfATF7bZgSaDlwuisM7RTHASIrsNq
BWf0SLCfrdodjxzUzTAQpXDKBRovRrgYve708XS6uTda/YomvXRX0xuooJWvKlUD
1U1PpS1EVdSHA5EGBZzuo9iFvO7H0nQROJ8nTcwUOk3rJWzhQXXxxFWkoRSQ7+cT
2GaJ0Y0aRB43OHgbpa8TIqwfr+DAQ90nK15VUQ7y+5ZiOcSzpLMMmd8F+J03rHZ2
JtgSWI1SNWHe3L5KQDtYzzRqwWsKIc00HIt/lcf4h1Qer4hWmcdpI+o25+yYFtmH
oZZTHSE5zKqQfF0lIWJ0bBDb37UYZ1GiCiCfE0ZXIZ6G7wVl6oWgqwDGqZfcSR94
CQupv4MWXX/8eKS7+CXDdJ3MLnqhiSsmNjsghITPXnCGRg2kYnet6aZJT2p7j0WI
AiPRiUJUh0/0fnTVKVflTRVI2N/GEbnFdd/Ds2BzMdw79U/5jmp+QTK6ihKiuP+E
61Av2l7VKAngeRwrjCfgkNpX68+i1dAuJ178Nt5HYMGmbFs/AIpwcIDKSYpUBlfS
gwqgjnuQDOdZD20pxMEPMi6XNga1fRLgxMJ8QbMtlcCtLTsR9114uR8qKeJ/TN5v
5EVXjdqqgibb9SI2llVz0PHzW7zfThfh4616KXBIyvmTx5xJy8KYca+ZdFok1NMe
18TkECVpXkMD9yBGLYoz0OrhTT1PJSsmnyWiq2EY/MDteA5Y8W62VWSCjNTjI6LA
4pm7uGXM+2Xc3s5W95s2o91vqopwuD64rhywaHUqaB9vo1RwVH4pCU13kSnYg1jK
lqjw4B5cJYGFjZOPHz6XQ8Ux54SGHfxYI4R9YlVABQqy+TWbSrDTnZmfHuIbqek4
YNLnQOlZdWSxUyJ98TTKztRxqd9UsifN7r6ZzaKxqKidg1F4WZc4z+zbM8CTC28Y
UldscgpClutm0HKxmRVFb8vjIuvjeRr4Rh/+PorD9YWbbMwsqDjbPUIgnoqVT6xA
XASuBBvTDGa5Y+axaxfEQH7+MvCp23W6y0/WX+O8yxz84OWBjyXBv8QYv5RKISkp
1EjWBMt7zD4yVqY8WUnT2LtYxW1Bh9bVOxNj717gtlGvv+nQuVPHS9ZNBs/ViySS
5dco7fDm44BF6bvtDrpNIJIWHCScluVkfXcneq2KlcQyzNMxnfDQcFd+2x5a0uye
nLD5KyB1fsa3LitG805C/R7L+vr7nVXRCCBfpsG4SB7yl4aG7cZhCK04dDcuXAnC
/Eo+6glTmgFkXHfECXa95ijEsOtQX4mP74CoHzVOS9VvcqT9kt+4bTiAPRYgkNhC
NsyHzj80Xys19gqQMj5qBwiFNNDGiuO3Xyno2xLxiWgpmHu0FixToih/A8J0VfJI
k/mENTPemmj9Ii2Sbwjd9H9JrqZyZidgqkQ/cmdQ9d9oyPdQ6MfJ2nwlsthisKyT
VJf7fDnbiuJhcc/+l3vUIOwpZtl7N0KocPVDlthQcOxF4su8CGyzYHA4dr9Lv9QH
3udB7glu1Wdt4NhWSEStLfpyCtHrefIPtCmRZQAd3eIPYw//17A/wk2PU69rcAD2
KOliUV2GPzlE7aDrObcabjGvBhNkUPESxnrNTMfREygWi/5TC9sjTGJNEBwsfRjd
vdSEbfI3zwjanlWoZOIV7FyY2MKxaAM+clzOoM40ilZKWw4h5R+b1ZYuZnVOg18s
pc2FWHiou/5tAsACOKE4HWQ1h0+t/IRUHDJq28s/HNbnqVgPEfUFzv/Ji1tQTvae
osmj3pJFzWJIFu9/9RcZ5eGuwhBI/TK7dFk6hWSGoXKQTSaJ2/pQENS48qPihE1l
SuXDU8+PZnhFUL95cmN3w/xc9NNUDEl1FUO53KNEjvCpEe5n6T10IJ6I+lYwasGP
4TvtX+ruNlmY2Tqft3MgOUiyzqB5yeEZ1BX+eKGuCVewU0bC1G/LlyeJD/hiaVaX
f0UOgn+jJF+ojB+37p8asfSMrrj8ldoqgUcPiW4A4nU8pfGTDAkVPdtqEIJoBiC5
SV+9BM4X4NYnqEA2/juhB83YmYxQbvx4acioWoPSx0UKHLZtdoBRX3JY1s89Cmhw
HqYXo109glzH6nlsRGfH0rE68qA2NFMH12/8/PZz38n8fKXebpudrzDLjlMp56+V
ptg11f45I1pmz0x3RPooRUKN8wLtvSpah1OofXWSFTWJgVC/PoojOhj68MAyNyYg
RM5b1daizx7OgxVpre9YfrRHonocCHGv7iIb3E5Nnbv1P8Iq9XA0N8SQPBTilt2o
+0yD4ELvoFlJ1022TDPvNX0aGgUgmlBtf4D1hO/zA3uyBOSU06LA1EIoCfeawLGp
dOaTov4fBrG24w/eB3vIkKYp/TS25obT8WyEaArDkiEiDlPKNuB6lL2FjLS2I2ni
HJaouAiWNmMoPNQQPzRHIL2RgFmvpH7UOwvur0d7nHI7tTlGHNpV+4yp1rz4qz7B
IDtKOiJWzyiFluzLb2d+U82Cj/VBOPiVQ9EQvsSJHzOkqcTXc4uEPMGGGiYD91iT
T5L1dpWiDIS34M0dTQAqQDWPnT+QIrlGcNrDyFODFsxf6SOY64EhFA8X//cAOEKw
tWdqvnn0rZpt9c6vYKDr7zXMQsRRWAfmAub/1sQeFejrY1uoUMz9QonBQ80gvdVR
FbzrfP5qH/oY6BtxOo2cvgbuWyAq90sZGK5+gbmBpEutMoGAnmNeK8vifueVprVO
PWz6t6G0+0qoWiwlijmENo8z4IP54ZaGcB3P3xdykOTSnId8liq25J088OVkSLPr
lLQ83k4wgVf2SYkGzhWvvBhOXSHhZqnw/d9CAsgU5yKC/UPl0Sh9m4p/7b0JMzyG
rkjQnF3LPY/uL72UzJ09xjv2tg5xlJC2i0LmdNoMY5TgIP3Px/szpKt/Y+HhFbDd
b7EkWXcfq964doTo+eTQCmQAT/U/olsQ9KOggf1xfecU0XDH+JqTdE7v4nzxhA+t
vAnXxN3cGKS5aUPlJJElhv3PUl3hB14yMIOBTnwemQGrPt4drPla7C7jLdBBgPkI
xoJ10Eikc5dlkMdkDD1omlYJG4R2SO7T8CZ2m15pIUw9DmMWC65Um7eefmeyiy+Y
ADh/jFOgk0vZWL6PKqvQff6D/q+8RUTsE+Y44PDx34nvqC+wj5YS/ScqBdFUX8rI
2OEAZrlTVcz3qVB7uYWYpzGsTK/qmRsVGnzV7HzFLK19psqBC/IIQljLgtMrF4fL
5b4YKiCIrC3ZoEIdjOdy2bk9wjup0e61B+ixcCRf8kJKIZc+OEOWNN0PMzXLAO/y
D5ecH1YXwyETf79WWFnZhiQP/DLc++ffZUjnhEc+sQADnKPgOY4FLekYZh97KHk8
KkzLBLIxoIgQXB4Ro2vp24uw5sy7SzWT/9UwtJ1olaY2AlA3zKet28yc7TyRrFjq
Exw5a+0m3xvc8Kab0mXlH9dd8WJUc/RiOZTdoXoUrJaStGYczw1z+OHBBlImgcfn
70v3tMU+ClSjgrSS7MitBvyN/usXiBn25HS6PHJcyCk1xchM0fq4o70+6YcKPlZO
fcrZLVEDnd8sySXsR6fO/75G3wTKL5tsprnpZUlh+KWQ+177j4xuXYEMn1V3fiQ8
CNeeAop2gCwFFpW8uH3E2AUbJCBKv6ELGJ28fxTinTMwo84NIQhEGlVPesk951bz
bEaU//QrCUTWkfoQaLuESeT5XzJAtjUriBQUIEhsH6tcgdNyndTPc4D4UzFlmBeQ
rQvnZJuHqoa8hBZtnTrgOk7jI5oLXKy7sd/qByJ1RO+0elckbC3FrRecvGs6qjzL
DEP38ZREVW54xbAXkI32kHgLRGgs+gzG7WEaON1r2xiOm+/2PyAzLCoE4N0PDgPT
ZD9CzcU9iMamLWLi1D5FyLMn9a6dnxvycII+bWnj5R6ELDOo3y1FYriYQ8fSf+e6
WV005UKyyYuZHqKkZ6niqnOnbzRql2q+aTGM9fJgl1fM09298IrFLw1h47u8xnzj
u7JpFps8sXDR60QCyadvC/WEAuBN6GuoioZpt3wt7oajKePIRf/NCF0D5bB5Ctna
wWfnK9rMYCypFeGAqMh4nL6UtyaWURj6vQ+H8ZTb4QMAZ2FhGWE+HwgYSJM1jihP
4aNrMDiz1MpbAzZChivz2ipyye8asakbV5z329fIGALacwQu96ZLmiZiVXul31+I
5K6ko5I4vTzMiyADsm7PNxqRt5Jl1tCICsek8q4L80W5MomCRpjfVYSmUw7Xy6cx
5LDhZYZn+ETm8WJw5xW3lB7iH0RY5XPdXOCC31nqTDC7khzJswV1kyhCNgFJMWTs
EYWgAJ553eKIGr1t+2ELLlSzNLFgNhd2ObiyRVq8DawORROx0/QEA+Betjkc4vto
2J7Y3JzpPsCx0+pJ+7+glfnoJ6qzHT0Cl57M3caxlm7LNuZdGDO4nz5kJJayw/BY
Oyr2J3ZYypcCJbg0+yBrAMClsSeGzrzXJSC3rYHolcRkUpJFCc4aOFPCQWDFj1ay
J8e3jrsYzjEdrCnxExPKPhfKJBT2bfliah+BqoLDbp5y3CUiAILo2zcjsNFkbYAg
2KiYui/EpFDn2skr/Hj7yuGyvzAFcJ5kCqqSVj2rf4UlSDQhvAaSrc91vn4YcJxD
7fv7m4/T84y18FBbqYlLKvTzijy4b7CwdzKuI8tVPztD33WKJ/+ULC2kBLY6n4Gc
tGrkYr3POj8RW68AtixygwHiU5fl0GHbBM1qDdpR5OQaWszcfVGrPtnOGD9988H3
85xXrmnpMpoyjKCS6K2JQ6WGNtS6Y9BjKIHqUo8zbqZYSP9AU3jZPoHXCRIIEMK1
Q6IXtTX495NBavr5FLvTVXCChpOFjhCQafRwtLE6Bn/Bc0h+owuLMw3/PtlM+hGb
Wvp9ep38IKfuSWJbiDwowQF3cUScdOlP9rBKARiL2+AlgsNJuswK3puEM497+6DA
SlArMH7qc7lUgqk0/7w4RPDzfTuDFs6dvZxk2pTnyZY4pax2+aAte63ipF0ENw6+
70EzBxMsjIrzYSXUZt4+P9zHcSERZxWZMdIdGG51hJ9nocccFpAjiGlGJ0O9+hlk
pOYg73tc15kHqR7sEMVzsHnlnalwVDFW/6QD+IoB2VRGCKdmvL+Y/jM5l+CFzkAs
TPEH0N//SEmEpFXfpLa3kY7YotX8KTHw1pRFku1ANZZm3SfTskcGe+hh1DiNeKlY
iBoZ+S/2KF8NGuOxb+8f4Fz94b/jWrgrB0YiFYHzHhMARz/g2IRnu4RsNhCel38g
U1tpQiqIcxNOEgDjlC3tAfAW8XABfozPbr1s8zMjuzNsNSfn/g2HtQ03RqASZ+a0
AGFxjOUc0z3BNis8n8dwWxaNZbD3ZhFC8KvB8MacfY6CEE//vtMhH6kjtbCdDrt5
zQRY/SzAFg9tsX6Od0XAA03Nt8q+8UbQ3o5gr9KfYjdy2xvq3THsKHIZXx0svoPu
zY89bXCyb0taU+pTd4D7qZdqswohkVAd0UkEZpFGGaCMqwDMnDAGAzWlgQ97mHb0
W4M1hd2zeipnrgmeaVsMSrxyBYdusei28B1nCxVKJDZgFQFggB066Urf9699jPwF
ec9O7CoRyLOvSnQtzxMTpE6PsvhP8pmSZhZ82tabg1Yl1hPBzo1mdlIeGw3Db/du
kZLrGwgf4vJx6lrlDEZr1Ykm57UQpkEBLGiaXMItiPOI+MBuuILV3wvUveFncVV/
CFVktaWdhDs8GIABhOLTov+wBsYY6ndbTn3Agq+eV+S5aoDZJl/eW2Q7gUzZbf1U
x54qmkei0Rlomm0+S8/4QaCdwtLQBCMJbI6i7mVNIhREjAsE7+D1w2J+QObDTws9
VmOVBuGYNProoaf1z5G/JqZN2HorrhTRWn7Hfvka9XJU/tXZGFBETrCskitrAxDJ
9kgEeXbiPZY+vqEt+Yx73Ir8CmX3xYQ1Sce5OCKC1u+xY07Xg56EPqUeTHXh9RLz
tsDlFNZXo0/OkxF1FE/JWVO8BO8ZaQOuqacKGAOgRe4iok1ujVzj2iLvS4AWm4ea
GEE1CMZLhBOjjprY0MZ3Hi+fyHS5dEuL3PVfhoRmSPqO/V26Et2Kt5+Fnf3PE96m
SdnLG65JoLLtPMnyTJBRDGbqC09TskEde6jjvsS3DKKx6jFH2YftnbMVee9lVrVB
mgSsL4nS69QcbIrpENYB3iI4/plc4E75qM3E9Z7zJ4zmxAAapBezg9EjfDyz7QVk
5d80CHFetP+RW/4+PG2ho071SEnPGuDWszTz1Sg9BVeLtgmKThKzfWu2kl3lMmPK
6L6PIzcIvoTeqheEgMXN2CAKO0G2Gat0DwZA9q18Y/A7Jb1u5iUku8TZ9tBuB63Y
MM0fldmQ/rHVAVyDj78SQHycpkLXAp8E1yfZqHWWtB6gqGutga50S9CmhGhdv3kN
152u8H08B8TPSGj1Ik1g8hK+PSEIf+0ymH92KSx4k1iPVwlxVXIxoYl2ceFdsgFs
G14k00swevuh3ZaIJiHm9nbvUJqWDUxudEnIdAuustNN7KQGnVBCPc7WyOEcr2X9
gFrf9Mv5RkLuTxH0sOUh9+Vm9iIGJS5ezB72eX+h+8IPTaeAqkwMtgjplG6HlTny
T4ZLN7EYgi8G3TJYJ0HsC9DokvHk9xjNOHhE1CDjliTbGgTyAVXMzQCU0mc+bVg8
sChYPhDTL1ovBuwvdGK7iCMFsN4FPI2xWceCUO7h4B2GUg7HkJUbdLs3wt1ouBru
/Fmo8Ua63owYx+RmfgujQ+rDfS1aloifLrzWIBHaNw+jM6faHDXGmjP7JqrdpULD
mSmrpVj/znPAakrhDNLzUAIvk20zMLS45kn4j7UE3FoQOLFldMdb+qrlTEhhACHu
UxhYurSRz23vaqgRGQRrHDk9Ixk/MNbIhQYLzV5hgZHQMpn0jDdf5mWPybYGucN/
Ug/G8GGlmJ2zQCaNnXR9xmBjrgiemTfbNmVdSlecDTrtIX//T6uM4fRiCRzzEBXx
m2o7TUHweZuVzPyf13Ih/zfmP3ZlP/PCJbcv6kj3bCKXmeUxc6iO6fJ2AkcU8le0
LqwqtAFstaASOTGF6PIULcCrE7JUHL+6KyokA3gVcDZW6DNkxA17PLO//rVydvar
p8LevK0UViBXYWF5i5sHlu12dEQ0YmThsLtPAwri14iEygzCAYpubDdBTRGqUmTe
UGIOepPk0H33FK9bYANANESnl7LCpkKDDF4180YVZ8yFrxtRMlQn19W9xTtU77Bx
7akcIaNFrb+2SHcinp5lOAP6WZB3msPcKSy1vCX0k6b+g42z9wjmi8/SoTn/cwO0
vKwQ6GXuBMdQrGmhSGSqIzMhmwnpzYP4CdYt0u0fSzuLuD1/hpqUNdgkaUlox4uI
noJ/AJowz/ks4wS1jjp0zEqlDIWme5CdUuDFjYEBLIVKEE1Np1bewFGT/dUNKfCP
1k0z///TIASoQ541G5MxwlN80WEkCz9WvdlrenresxtsGG+c9N6tcGoYkCKgkIXe
8Hxj7QH2LtjJneii6KEpJHUReT/7xURna/MTGdK0xIzQ3xrlBFPPjDm38u49VhgN
btwavVSPSfC/kwRpDKvBpZUpypHI4bQr94DHMpmQ3lFfE8sS4/23hZ3hYygX0e1P
mBXjJymPlKRUltYHA1X2HftUsH4JD1a/eiI270nWSD/QJJKHK3IEsf76of8vSsWR
boUInHmQJhtaparp27yibHPV0gHX5etgItH8zasWJ+hnr96C4oR9TVxTh72A+/27
HaiLQmiEG5JSgTIBAf2Vn7smKcC3BMGH1A24LusbA8BevvKqnv+x5xhh/HdorAK9
cVFbQj0HcMCIx9NrUAO3r7aKFM42qB4c51Dd02PCOIKBb/DdF7JbAzAdfeuns71m
vcDKo5olqjGCdr8SNaLluqvUMV+1IRIogjsCax8DjYjjHa88QC3cEZHbaq1KocTc
6SS1wSG6Kcb1Vk30vlT/cIxtMA/lM8cCqiOV1amnVrD0UBrkHeIahRSdAllEn1i7
MfA477Rukg3KSs9k+2OIwhnlx/yZM2MCer92ZgoKKqCSEArcIT9gR/x6M9LWn7X0
BMbY+9HvmkWe/Key8HWNTrKkT27IEnH4iLjLguzROldTT/Ztcg4fyA+t+mi+CEwc
qKAwijLyn/Gha3g7vSz/6NqB7/R33v3QXA4Qvu3XhH45ZwvM6aAeUnNGZyx0NfMw
HsFQebpFOcly5/2HjY32kwpTZ6/BsMTwRQ+p4HlJA0X4wXBvcqY1Tduvh0/mS7tS
WsNgE54BbukiJYhQJjFLsM2HSDQk+n3ss8OIRsAhrfaGd/NC61+bFnS/QCZehhwO
Hy4rCkJZ7WAB/DD1kaishCb9Det3ippvR80NIdRSBoVpGHSo246IZc935Ya0L1OR
ke5cdein9kgACboZH5Y2Ct/nmVkGKS6shYHjIHnnXJIzOerpvPJLYqlpi01aGyIe
p4pmZ54bd8nIrkuCC3gLTE2/P2I3H1O6DWGZkMulHGY34BvOcnVcfNm5U7McAqBX
eFnVVrjBlj5QwIWADMNk0sfy5o5tviWfHxaHZWVrnIyxhEJoK6j9Lnukd4Gtb6en
sp+Du94rUc9i9+8AGapxlR3SXPbhe7oKSkN6/XUQSKoxwGvxde35LBkulK+7Pm21
oyIiNcm4DoJMc0NaeTxln+3VLu9FfSDfUO54leloEH7C3h4iOAP2hIPkkda9dicG
8vY7Tv4xj63VSyarMWrjpwLSjsVEt7pBbrc9dHAjef8I+JDWB7fLX6vPzae+9m+T
8FeecSgsrxv7C+ffvOI+GOZzhnmYVYFuUjrdgsiqoQvw002Wtc4mBiE9Q3bJhhD3
T9E/5YwrF821FWLhPlSCpYh5Obplbt/75ubHNsz+L5DXfZ0I8ru3i0ceLjo1+tG8
mu3kj4RJO5eG1ihaX/UW4xIeKXmM0Rp1wxi7lRP1A/I0Pay26KaBzIojrUeHP9OQ
7YgHTCReZGtCO0RPjeOR1R1woGVtVu/QsRt/i3aYTkLDiVBe0pA+28u1Ex6zwPYf
NmTf0AWutIOD/k/geMSM949l+VGzvc+k4zWz8m3A6M1Lk7IAB+PfZbQJ+OhXA74w
Do/dTuAC/3WlqXU2AVY5VhH6U6LeGy+SDtnTWRMn/DX6R2QPgeBk140BEa6rZ/Aj
rWMLKO7tZT1/9yKFZ898O4IvSxlTOsDWtpt9MefGBD1id+mlMUb9DlaGCLmbTM/A
oDaZf80IlH7ZRNOKXILS/iskni7yI4QIOVkdDOvbICKm4mwj+4CLXB6sDh0a6Jeq
6tLpoMtohI4jH6LdZGUrtLQZrom8NJE2C52Fq93i5NcpQr4vT9owImkn/Te4oNKM
0ov8plxhXO6LRR016lnKir2Y7BQ5AvuIZlZDKeLpYpYesU/BPklsUYWmXu4YTyXr
bO5gV+X3L/RcMayhGUum55yc+AhkpPc0/M5FoRpZrehVnpw4FHeQjddlw4/wjsnp
cUiJNM4RK67ctdT3AK0AykrX3cbOSxEHfEP6lJikC6OmgJLcZddrDjVs/9ji8hSi
kH0Or+9CGGsJkxWByiakvI4yVKGcUB10802mOdfaLkgSQKBxP2OYTFUG5PRm/ExA
JcGLZdKpYxira5Vh/v1DTDGIxRmUCgF8be1nIpVPfX0bKyQAzz6h6MXNYCO1VGg6
ODWbGc9JAg++XM1fKrJhuhlHvDaixqe6MRnwR0Ttk2TJeN/FR/5K/EhQvVVIFL9J
DMBjO1wOdyHgVRMN7xTLTVPaLLsvDIqUI3mkjpjsY/0Ri09dMCl21cZrSw9Fkwee
D8P300ZD3Pt8cyVTOrmB6+2Z6amX4clYLMQYta+V5YDvWkKBpry+HPft5VFHm/sC
PJege7OQ4DQZtbppo9Ddptfhkd38Z+KQBpMfY8g1A2SdA+LnPF9aDfZCGqugRRhE
E1hWvCWTD0LX2dYW5QDgTeO/jIVwAvVOL5JVVyV7W4eZbaUz5+VZfI8O9gHY1e2X
CZaySdBhK/wogyNhENNCt8cH1HpBZ2xiBdqv0qxkCcENfXvsBStS0HSLh6YdNDoY
GF8NwtGUieKXu2fxlTxGDu7v8N96ToVomOWnhpJpdFP2e3NkaTCuB9AHzi5K1Adq
vFe4EGOhfVbPbBk0GQbzFEV0u7sSoA6ol2Umw6QVtdPRd2xlhycqs5L/zQGQjQC0
f2Sd+zKculeU+y7PPWBlisvCFVr9h0XszWiRrZMYnEhDChmcP9PvxnVsalKTO2AW
TkogrMZDFZlHZBRq6A7Dt96aStc/MN8jSwBeb7yRYZGa8UIiM7czGoQC6i1a3GI+
x+DJmQwHZxiIgx1Q1ONbkDzS6Y5A1oS0hEdkwa2VgBzEizWCeeP0lqdVmxLU0VvV
+Q6JfqXKqdu6tUA5l2SWYKKB553ZtxLvbq++lqpokS4D8FYlBVssDYh8sPXdgge0
sPwaXC91LagC5Bn4vOPqPGBAWWI/bO2pDwRceoXRX4sbVp6qiw6AxeBveIX42C+Y
ezIwEuhATcpZnRLDKADxhInaGRJYCISED2HfrB7OCfuBRAisWjLWGZsATBQROuTz
OjiiRmNdPmtHvepBE3Bod+rMYjBgGxRwgYxy0TDCv59SmHRleMiMesCjNSZ0Zh0G
9IQT/z5hGBbSIkzSTq9Kg9nQ2a6KjLj38DqSXmRotwUJEeFWNrFieLTDMGtYJk0S
Tog8nvM0JL8gHrZ0dfBhVTXhNS5B0FMuYEqDGiBzbv+4x06PSLL/kGqXwoGwlbp3
k6+3LNzF0iNezWSDqLtnftLkrBAV2qK4oSk+51IX0+cbwpT/KYpoUnbCmrftbEbE
P/Tw9i0Z+TM/zwLNr00UajxK0a0I12WVijNKXsD+Gdh8ELp3KDNbmkRnUyt4YvO8
lTo0efOcCER/MaTUeaYxVOesmdaOlC+1TlgQwJ23RtLP2fjd/Cfv0WaalsBJmuE4
D6W/d4btqwyH38fP85NWkks19g8hsXx+/qI7XpITG2IAtHUgEPcQH1JZfFhwxaOw
PZ4CqFBs8IYdP64hZvRMOb1uCa8DUEDBH10bTPQYOC84VdeMZBB61ixjgeTL4Ah7
QxQ0KrGEa+2st4IDPUs6uidlCmdG1hCihYW1LDgQsqbesdFJF2VqvDV2g6pTuQaD
ZPUDaH8HU/s39X2GRRDTmrIi4/1gBaIlfQgJmOMS9i99hQUOwwzlSzhIB8QythD5
TGaHcGKrbuuerx95FGGik1ufgCzWH6QPO3uj5Tna25kQXPFSmDUrJ4613h+g9DHu
72mBP7knejwXdaKUuXpcFp1NRgNVhGGbCmbMIaW0deyI1R7Sb6Cq/PSKTg61EYSY
k2FGWSUqQwiWsROoMa29ts3Df2vu862K8lYpZEWcEsRlMu6ubH4ib9x5YvERTq61
tFaV0OxzmIjYFSNkpU74ryAXsTkJb6rXyrZkqtm8BDnsuq2sH/HRk9gLFmkjZ2a1
Q2h6iG3ZmP7SS0Xfl0fNCaaQ1+CnjLByaWDcrWbJYvcnM8qzc5K62KqFYADf4/X9
upogfbFg1KBTDWHD5FUZcwAeRXrpdO5nKIeTh7dcEQPLTXPqgEk/pAz5wqTozakV
T02aXshe90oH54I5zuB68JDyeoqBBvYMDfQePzL6WjKxSL6Zjf1OchAsiv4+0sF3
0bWb7NAKW+kIiF69yvlfPPJRFD1r1EUdA2T2BaMbHLX6sWJt8NzmP/GGlqd0it2V
9tRzfnPP4E7bPtRnOSVkUumOWHtB2C0JOphBjWosMUwRDycOUjrKmuVXj77tL0+1
SCDSSoCxDoUEO5yL4Qie7q5KmWCRSkyWRq8ey1RfHIrltMf+qM+k5Kb5iGnoQ7zJ
HTvPNZoVyaj/b9QgnShk2zMvLRPtv2m5MqTY5jvMHEf1luxZPyhPkIra79mLDkgJ
SG3XdYmivzYeRKXHRnOXYarJLR6Xkm6X2Ndi9RVjWLUS1A0jYFdDvYKIZ988VxUl
d6wif0GeQkK/5/hhAA66+jy5w/159YCHvTNQQ0Hugwd6qammNN/amtQOgwYsvrb2
jwXLnQH7jw9c3TEDZtwTS8ML9QDypEVE7gNEg0x7p7SLJgVKr5BoRPfYOzqb1XiW
clso8YX/sbyLe+dtSX2+MwP+SDY5TIDU0Lu/L3Is3JaFM8VO9r4QBZZg2IQEAskO
TC/eJpuQ+aBWzCFoGyZWjr1hWiLc//bYVK8yR5uhpwP8T59iTrFF/H2l959xC6DX
iM6NmyeNKMAqi3qyx09lVyjoumGRSBkFoRfT5L54ptBjLSPF9ZtZATfZJ/CfI+aU
B4PBrlRhDz+TPrKDF13SZfnaT4iUELRxS3K7ry9k0PKDMIXDK2COYe7LDYehnOkg
3xKo6mlWH3qqp6UWysxPv404qfh1G1H9MobB6sc2SY7OcxRoufnrZn6CT6pJiR//
s2w698jI0wu0IGi7RwvxcnzGS0UcYl4aS9YXDHfsiAnyuLrR6CyMnX7mfXVQ/IN+
Qjm35YgWkCecR9JdEtfvx+x/dMNY10E+LWFruuo6RdALPoijW58cmgO/mzajATGb
boqljTqD/PXnlw/hz6wLTnvFLXTWehtpOTuVo+BY3YwqVu3d7E4jLX3rqUnDjL3I
sCNU5SQFWS4vbenUaeCC4dir3mWRa0CbSWXw6+1RlKhGjH9QI6t5fHR7h5zbw/UC
k6mDP1qZd1PTgIjiJQykAXA9qDFUluo2gny6fBVKHdXgctt2cE1uwbKAAoMOGxpI
zP7ZnWWlfWJzuB2IlDI2H2NDmXPJfHayvTDcURC7lwBVmh7GVaJTW5V2xvjJzph5
9jTJSJbSwgdeQEHIqD8gUA/QgihAKeKpsxjHREggbUTG3IkpmISOw2p6Fg0F1L7R
EMP+ymYFfUUVv3sCdZHwnNut8Xre21nlYD+Oh9+fg+7RuCyqmKFYqfuj9Ht8L022
nOSttU4OPR1Q4OZokn3BGcIEgCFJBaO7d9yaReTc2NlvGt6fJLaSr2tvCWb8ruHy
+nYyg4+1EPB5Kqn7gbnYz5yGPEHFfufLNUM0ui02lCj/+fm3y+fq8Xm9dAOuhdrF
1Lw3OlloFLu0DgB7t2ERX9X807ss3Q4DTV6C9SeZ/UMptx+LBXTVtsx5+V4LW9hf
9B8i2G/JbjG6IT7G1AzXuz87qAux342x3qM7WcnVnovVCM9E7Qr4JOgBxMqJl0yz
rXKuuZWPCFooh0ngeHSsAIwKra/WmK9kyWosx7ypi7J/71eKKidh/Wxglhj0vmI2
cHZtGRyDtaJFQQvUVFansIqJmk/TvD88MCWNrnV37+wTx1RdnkNwoiwMu8jQ484C
sNUiq4XcktygWfvgGmnEkhYHuUni03Fo3fs68o0o4xbsG30CafQ8M6s7Hlzhyia2
BSBk0HL2aB1MUAwaM6RSZFsy8Cf+MF9Vd8Th/uZ2MRcVIwwXXCpcgCnVoOUxTRE3
z1Us4bQkdubqZW8+EAIEO5Ql5Vlre289DDkxK6+p8Kw6tLhefWwlNIPNGz9PpesZ
fHO2BZDt9ks5eJVzbtSUq823GG8hfkwEMP969mHn168eFMo55e6parlmdQw6Gzus
9Y8iTTeks6x1SSv9FCF1s/bTNevPS5mBDRsi/iMdNHuJgHtCDLqTi5ruE5DN/Y11
BmSVzfEMll4Fs248B2cCg++hKrWdZZKcIewm6LcYpsmK+3f/lbqQMm6rwJpvoa74
LNWl1BaqyWzLcmf5FTKYnondLvpfWvb/CUvBz1qM2ozD1PI4VFgPqvmIl8ou2Ncq
qOoLI2IdWhs2xlOQLanf5BZtz3Bor8AWLqVN7u0vEhlZsuSQ2AF3w+aWLmglgY+F
QDQeZTHxWYHd3orbSJQYKhyDtX24dDbnk5walkgBRPNNDYrCXtJ9WlA2n7ynrVaV
jYMopnoUmHKiW4eN8nNKzMTfr+Qz5uJS7NsH5YR1GYgZebEhEeI2PYHHNb+RU2jT
HBOli59ohsVnuLY9FIVMUHat1RqdmLZnvixFBh22jzNbxVKrC5j2bE7qUlTACD8Q
k0vWPlQYFDGjIugjSTZ1F99Tf91pxSLEx2KoBQjDGxmGoI+MOG1YjqfihSOvXfBP
AVpRgrgy8OQe3ETkw0SlOcNz6nujAESCjdRi/hMdzFLafo35ZuhHas7s1iQY2cFt
RxfDB2VGEbuKjRBEFAnl4Laair1DPL8dj0gSAOcWcx8bd1jkUpxDDiK/dmTHEJix
xBDDo3+GEFYkKyQnN7yZ4XiF8D7v2yYIl+XY0+nqQPiIvufWdAxdIfrKJqICBORr
wM9Gexwi6KdIr7KllkOeg/LC5T03epullS9MItDzV72FMQOpyQBdpKqgcVuywwOd
qbv43ui6V7TcSB7bIbYKj6sZL3leDWzO+OJwiU6SpEFkOERIQGmCoDFvSDy2sehp
CyeokG8Fe6GICJeszuLSPeQYRa361f+Kd7ji2RqauO3OnfVAAdDfIxnROqCyZs+s
jYVJV1V2EILvtthF8bVoHIdrc0kU3zarUY50jfb1cdv57fYofSs2ObtVv8Q6zOvS
4VsMci0s5xiPbT0gRpphczS53q5QJJ08qoMlgtKsWGxC7zqGH6b8bdsT/5PpdYtd
h6+ZTCR3Kz7C+5hAdKks0jr/731DGr1k78fp92/+jSZYNzVOb9v6ebqFZgSkKWXC
kuoHALdiNdGolf/A/RN0TID4DYP4CVmg4vM29lrcqJBmhlRy4K7BS1Vn5VB1wM2G
b19Y4vvpi1hrUUeqNfSbCsrlXyXTaNBq52tPgA2CP/2zjdaHkzemXgNsj6y2wQpd
H5RncPBHYExL8gB77EbI36a88O/h1+5saAyOjYs8ZdIdZFywMp5IgK65/zgMf/M1
X5MXCcsCxYbEwvITBNQHn8yo8tqKJcuDEIFKs4ZfyTuVbxtjDzH/UwgOxOi6tN5P
wNIfVwPNnrGmB1/r8vktNjvAsxel0X9xyQQ/1kE9JBsKyWKz7p7ba651rGeV84d9
wpLrnfGYN2lTJli4enGjgEg4yDUTUzZ84i32ZCGwqykIo//LtcwwzhNTAm7eup4+
5X3i2Eq6gZKJuxs6RWZh5v2A8/PMVBzj6H/Mexov6HSsGJx5eO6fvKvWV+qN61hi
Ok4boGHZSBj3cG/uk0Qq8Haew5A4zXvEq83Q3/SBW32l6WL2kQQyGFoUzPO7+c78
2YwPVjDe6XzqTP1ZzUfSYeaNjXHyX4oeSDPw7nwAahrgYdi/SzZduRLx70I3RjK8
cHGh+EEzSM6wI8LKFeaM/KP8DG8yDX2bzx+ZDSKEM6YILGjn9DrCXIuOn01OG4mi
AQ9pRE0znVYf0rts8XGMdeWV+XHXPzfjm0ZcwVJA7Hp8rUFPPjhe+N7DXzabaYv3
Gxy93BFinwZV50BUSMdklhSx+W9XBQIJ1p6V9+22ZMj/hdBYyudnilYLUqNumCOl
3NhnyFurLHwCoYQ2mrw+izRVLJVsHSeOK1+s3kOBoxWQrecMkVCbGZd7RoOollgj
TBc2mKWFQX+hXeNyzBel1gKJS0g+2QzpjSuk+AIBVUfbWYcNX8x0l/bQck7d+LCn
GuQCG29Ch+UrNDMC44Ul6VHPVORLWO6qnb74Vmr76TLu/aGB6IgqQQF3XGtJQatY
9h3fLKYIVJcJ2BC6WzGh/RhTtp4POAtBstWi6P6vS5/FytT69NFDFC/R3lYQUmN4
/2rlb40fgo3RIcfLt4DElzPhQ+9zjoKM1H7V9Vr8bPFUDVAVxgUiivw8WgovtzEB
apNknIVt0SgE20njDxwdlfHlIg+/cFPfhIVKXfaCYvPFNebj66e8pBfhGwCRdn9F
b2hlxQKQS5go050E7KlJuhnDYMJAYsC5S5HxFUI8blJP+i0tXUtQULFa6qNgdCTf
dMC8daRrNcW4deAvXZOCtKpyyOW2Xl1nAooyq/PS/yhuVDKih50UoUJpAUA0o51D
1JpX/B4uBMgF3B7KbYGLXM0t9ulaedDNwojKLcQP6A/3tqbEiAAs5/b9O7BZhkrv
yEhxuGdXCiWci8fzi5PPiZz3eb+95+cQqZq35mL80WMcEYx8uWkGP7HTfMiK85mp
Jz0GPhMXbCaWXkdyIYvt7wax0seiefpNyTkniNg3elPOcs4goYqXUs0v7mkC63IN
wIIYsSgL4yveZZXKytT9yZ+/wWJ8LW+9FabDZh4Eky1clEoOFSh1HdzYMf80IQ3x
nqrY8EleiAKZtVivQocdiEOwIx/vMTkFopGa7CeTbJFrgXQ6aJD1EegYNnYRaHaN
a5YMWj022ItGiMx29erVWTAwh1GdjQryr2UgBy2SzLnCFqq8WH6GqM9CLD2CynNp
V9D1L8Jk0nHNTKCUQV+LNZ/h11QsF7YrCtInGlg7VTFR21yHKZMmpIygaFx209QW
74YEuLjO48fL4/NzTSiaFH75aCZo6FFZvZoIHyA5t42Ak+ftd51aRQ0hc+gVsmqT
/yOFoRC7gMPeSHWrie4HERPgslHbQeUUG6lqAWpLZ1BHfHVT1Sa+cFMB9wCAyQhk
5PtL3Lu8aXSMFUHtM7pLmn+xd32RjlfDuAzwzZcm2VJuQ6dl93zrrn+NIWj7AzMV
sHizjzg83PHWuScPWk2+2vAUivEo1gSibaesnN4JYCP8b2zW0DR7Y9IwX9fU5Cv6
WamezKcYrBgSoqjZ+Y3o983sedjfu09oTLTvQUZl5tnvbKFiSGSnss+OPuDKLcmU
vtbl4p1S0JQ4T6jzQ/B0Cwm77T17urb+Hlm4F6TbLVsLRwxx+bIdK8ifnnWYyHmr
dPSyQ0JsJPmnOSEVR6IhLjUdbnYTfGtjA/ypHQ7yxmRsrd1z0zjlJd6RHunOsUi3
IxOcx6bT1aNsieI3vAFDZTWAKP5I32wVAJXFZHvt1c6OKrXL+1JeG47KGvx/7ce1
FiS9GviSU4zdKdKvpaYe6hmMInJciQWAMypQQGKyg350/PXcX2GrNOKUmiN+IU/i
5rdsqi3PYezovzqfxnv6eVNV+7SZTkXUw4ugkLoqFLgXqAZeWOmQeHgFW1Zrqkkq
QB2oHK+acCYBeh49/L/OS/aIKXygmoI3Vg7suGjcXynJdFj/C6VfQuFnXxNd43wQ
GRnnOB+p/Ct1IuM5vsvCR8nXJl/Rss7J7YveSg++tNnuYVbScirJYieQc6+KGRmX
LMqDtrrGu5cUYJyRHwJVbFB1iMOlbIzFoIL1yfWSqluG2YiPWRk+JjWSMgIqLhWo
nTb1aeQEmWJjebKpHB72o/FAZqEZZ27ak5wymAZQiuVhwfz6QGlhMbOXpE/FOkjn
aukYJUSfXNE0yqH4tIhBVgX3B7n35vTmAuymBsqTxOjCnlgIWd0r9I/HrHO3LNOY
uAby6FvMDjSh+j/LnrnANeH0TwOeVQk/+wC76yEKD4BVJI17QFRcUqeWC2gY5r0p
szOjzi4V4RowtKUkv8EDIUYbK9ZT/0y2ot3t5fqU1wbQHeOf7W1SN/TH11UKuH6C
0O/Imhl2XffkCLsPKY2xd0nU3QWwzAFRlEIdBwx1fGTlax8YIyuCrVYpOIw5uLK4
0ymvnnD2Jl04fKdRb5wANc2nCpOV50NFqRovI7J7yA4Cc3JTNJCoI10RylvJMGDj
gqqwPsoAnKj5SusDXYd/Hae+8s6o+k7ZMhpY6VZ71FMYgGo1MLRQBXO7MXKRc+KD
GLRmaFVf3coAjjO3rdAAqqpi+8WMGT3zKtYogY51SX44PlB+3jm3gh2ir0CXGniU
eIuya5xdAfygEKEgCDOrGlGwN2uBDcexT6Tsq6hQlkScWc16UQ244q1FMmfMNmuI
qNbIswXIxvjcHR12+DCrp6274rhdphel7qDzVMWjd5nbcM97h/A1d2xEv65hpP+3
eSRHrux+ddeXccjdtJ/hez/xaCo4y1/s8ZU5LhPtBk03VtVVTnkSjYwCTQ7F6paT
2QNqkjfFntkz0jdwFIkI8uWuHUJZ94veHKWI7cq+rEy1PHXeTvql0sLz3nNXh92U
JMwnIEOBoRkfbbwBEHTvKveci4bkJ3JXorlEhdmM+O2nSYEGHIdfC7IiiP9tjpU4
uY6/HnS6AuD/sY6/BKVHO8xjNMVr899fekc3cRC2CFQc9H6bSTNmi/0Z2ffu8l1T
jdoZcYBvBBNLyjT7hSJ9PV469HVIp28noB7TLlJ2CsjWLPxWxgOwDaywlUYyAQTi
FLtKkqOvxfli7at2DtiMYJsqyoO5mEbC24eoV0LJ/5arDRsMWH8eU64wkqJwh1JF
Qao751XS3b66cac8dhp9PXE5s3+PFi5pOV2cSZOmHu1plh1rdZeKmQwv3wlIQavY
xvYdZl4i/7RP5X89Ae8ZhEazCe1jTF73QLQZX3HN0/tH+Fr6vDW455T4W/yre+qx
8ySa+e754itKQ87rQ3afWWziA0QMHUml8F9RXtCNy5Cpn4z5GA4Cxdn+PkM1RYOg
7kESSlKdxej2HGIw72+Oyb+EFj6oDzRTCtw0QN6GpSFbbD/+of1JPMO/gSL8tkWX
Bctjh7WB/JjiodUGVibfvzwBjv0veogOIEON3FgKDYVKiKqy/OAMbNlUlcFyWbWe
EBFr4A2aYOQJ4FJ2MtMF9EKD74ABV/HN33A9yVVdgnU94h4ffj+UxWcqUsq2VMMG
4zR1F+/xx2MZmdjNOOIOg0q6PRtCY5pZHpI+3zTkvj+STC2qF6XbMfwMjNAprfMh
VaiTqseYnzRZXg49bmCukfJJIXBcVmMwppj87CCxZKKM9s/2bzoDQYnII9YPRrDb
C9PSJcbZqk34Mf2YOWqXelKmY9sqCygcRbUvyuzNdBr9/TY1kfIoQMLR5bTWhdTP
H4zmJBQSR1OfzAaf9UwEBDH6HVWCneoqgV7/D/p+YcPmkIKizMjekwjC2k0Z9+IV
GdT66E6jkrIt3KclUQLUJNosJfquVn7w7qEvX6Sw/CficnjEMJjjWkOz32yqPxnE
gaxw3TbdwMprPBbnWxrrULDbWtd0/V7htK/r0cpCGD0FVogVnXHReD64PsTmlUmA
EnCfFsZJUtD6WvwJ0h9SgzjiX6QknlU7pxxPKrxMS6eEP28H/df4jf3EBrN7ggbA
DnpAn+Efx/+cfgnV+rH9kluJ3WB8th7JMHsaiXyP1LGhbwru3OXZx1XMJ/hUZJjl
ruSoEBUdxJVEZZpmstCZixC/7wEa3o/tE65iIfP+/8LOGzm8Z5JR7WmdxU0OV0Xt
2S4hQUhMjQOXLK2Z80NhlW6QxAKQuD3dNVkThWZtQklWqbrAeTH4UmdJpqeT++hE
49c57z+vfb7b6sbv8wZXSOuiZPiFaV9x982L5FxCDiBivT7VPnjR7z5cmTf+Hl9I
YHARCGJcLvOyYkn89PRBHMuMmU0dUFthJLWOwijsAHDZFU8XBlGRNtmqLBDx50VE
8QRCfn+AkaKh2pkGPycBelfYB702f4extZGoRhmnjNyoVzeFb7DpIgH1h5T9cau2
B7/mLmgCwlrTaMY+TnULpM1DJpyJq1J+sn9gI+O9PBvyGXMswvPi6IZyOHW5xWcA
MtEM5VlLgnX6+K+ZVyeIQX9NRS2UBHD2/yD1Hj0IXRjcnG+GZGojwZ7vb/hNquzb
DVJ5HkCdiYtWk81b4dxsMwx5i6HNhP9GAmQxmaqDPujYzX3Qqu4/+HlXZ6CuIIEI
ZXoa2jrDRJecRk/LRvU/hngd/nTjUeICSbduLptUvvunWTcZ+T0uufIm6b+5iLAO
/SrhqrfadLgIfqUmbaQ1oVhQu0K/bUiyZ9X5VJLAPWJwFyEFNNJEYv5gt04JQYfY
Ib316YkiO7hoI1TQAnafszxo1/WpcYnBWtNIA4hh8p8GnKAKP876UO02ucHvIu9y
ZIqCLZfHvGY+/YtBvieekC4awlPeP2c2sCFIKg7HgYjRztQ2Gbp1Lzdv5E8ejkZv
Lh1fodZOjJP8vCcgTeMefMecRxKMnvdADTwiV/w+n335/pXJxkdf0AwWHvbjlke5
DkxDMcvHzLptT9A4w96U+BGPNKOgweNUQVVPzWcAU6gALPXMwNLC3yNB7atgaUhh
bdoklpbXsu9fxRtfRBhBGQKuvPxSk+t/qxQYSJ01d1/3iJjTad4yEPcUnhRBsQOf
cfSDMZjFg7BnIywu+7+On2DYj9aKHpxUNCh6NJ7onz2zvE/EeRcOugEe/MjMS/G+
76oSpK2wRjC7ieJbTNDwXGGFp4RcDEVa5+dvTwMBCC9g3nQEho7ABx9wzlaRcthI
kfKIOPcyF/xVCJGtYd3AQuTyZm8BeX3R4easmWocR75tW6x90eyARdVygdF0DJD+
n8aYZwe3xE0eYf+Z2Y1T72okmrxugUA0pltZrUVZg5qPtLC026ldAwEIhqawvnQj
XGjkKR2YmfAzOzgblTOSFLNneOKzfSXvbBrq9LsO9uMKwkBq1fZbNXBgK70NDXww
dP/ii5yfLHOkb3YUDB/wdCGkSztU6WMd6H2oXBWcHE0YusiLZZ1B/yOxiPoW1/Cb
jDEOR3QlsDA3xrGWAIKDbrUsi3EKUSQ0lCzlEMv2tAWvwzAZHp0DoPZvsLy1ssig
0VTekDNgx5dtUE0CgyRVPj3zaJcdX3TNbcxIEHiebZYvqjVzfykrhHaNr/M2zzsb
qiJbUPeLnZ+IbR+mAN7+DjZ8NQxJ/mdlo7fKXsm824w+faLNYmLKPOXway+LpHPt
GfTTYeHeT+NybYmNgMHP55Ozturmb0HSwNMbAjlSVN5DAfc3NISgcuYEPqmXNMuC
bbe6tHZBwGNyYd779ZsLbjvAW4KIg342MQpSL9EfjG0AA9gBECqDe/2s6m3khk2k
t1jqCWCu9H+pkNhBIRU5Lp/5gu/ENx8yvfHxR36C+zFdvzjxTKzGvvVADLpUJpAi
G/IAbL2gyLO+9W44dz1M+NZ4+WbklWaFEysL0/w9NHvenBFkkgfIvxjq1CgSUAb1
PKcLXyn9Fr4gxbTOWXxBqdsy2+A+qbQvdiElox/tdY82MNoORxNqkG+N0WSzuTkh
DynTIgTkLRNKzua2jgWBIKcApfA302nYpymim/cs4eVBFFGnbDgEIc938g/KIjxQ
6kHJRNfQuAEe450iIr2XWTwN+DVoD2+ShTyVAHWYrmJbA/m75J5VZOVKCzxzN+Oo
Owe3nwBfiHVCfX1QNjlDy8rB8jXkIyW0MEUjD5YniHSxuBd9Rx/3+4tjIGOYzKJp
yJgi1X5+rkBgigmT3Br8p67bfpvvaXF9WBj/1Be97BtnKF7qvIlG2tS/RV79PTT0
vWMYdzNP/DsBLiM965JEhQp7RWXyJwfQ6Xpzi3pQ6umgUacSg1CsS1wBHnJ026AK
Nq4TXFyMB7uCIIMX/CVTP6pcm2rQjtohXkltGtz8tmYL+/IxD3qcgr7Tw9fy8yqs
XfXj5waprk9QH4KSLG6yBYpHLvr9YK/ZMbKJVJbll68GZA0beeeOst/KlwLPlT+y
+Sba7xnQUkH1l9rqdyhNRm7Gj9aPcNkdlnR5Hqx8eOouLMiyzerVCc/uh88vNZK0
Zi0WpnMszVFu47b6v6fmQvoyarE6i+Ir7XAQoqQm4CUwRrqKRccac5yrwfegdBEA
PZWJqWgFqTvc8w1ftov/dOfqPE8Z5Q2zmELt3sIm0X/BkpthRXLb5e1k+gFLQFA/
vl5FSb95CF3HTxRj2r7EGT74WaOAYEd03pqHoHDzzcWjA6VpUVOMdisfxZOEfMOZ
iwr3MKS6KZ+8A31sRBsvnMOWXtLt8oAsz+VBILvrP5RXd/OfFejNqsFhDqbk92l2
RHite5uwD5IgYz4mPYzGkoAfJ3/zFoK8JOyOzKb12Dncs23iTlkQA5dfvBtCQmXK
AfeZGC9X//0+bYmGMiOuSZYSDJilFS87YMiyAPrwELWh/TQXNjT/hLSOQBjSzDl4
iHQ8k6j3P1/kisrBn1picWt6LY52jhEj56BzQHBYTU+8hLB0vtt1xsy+r1fboD8y
Y4LoHMqCPZXkVFHfyqnxkQyYybM2Z26rMeVeORjhSoXIjB5l/oF62yrTH9Sg1/Ye
qsCWRFgIBZhiERfaEnAFkHgxTQjn0pv1y1caTZU/J/d+LFyzBwC0gSdfFC1h/syp
ZD04ZuUD8s81x58ioFa00laiFd2esB6LGLIN1QeK3Q7nxUhtaaraKB0ChjxjJaiC
SzaC7+5NK20bcr7dx+mza7b4g8JnsRVueACz/dpqTPXGwRhBdFUNNa+PA7d82F6k
q4th/jboOtQsZnEogg2Fh0s6wvnjKyebfBN08chpSYEul4xEQcRZEfpidmH5DhYB
F1AmSvzXWgRSmHe0hM0vXXMHcIDIkXW/ew0ptHWt3SRLFuTSTUZJmLBTJEzNkn5v
pSIhgfVjuST7GOPlNsWSEfd64cxEF2yaOj5yX9B/MqGmsbzdTqY9xwc55smHhoxu
75lXDdUp5azfRDLJ8jvrKBx7HQOG3ZXqUamWi4HinFvfRAfjFpMCbOYtQZ9u6meK
aefFGAA68+NDgtTOCeFH3wYP2XsPoIpmQioyWwlCNWG8dvZAmNAvAmrMgnfHIGPq
USRhWED/Da4IefHUAeMsA9ZQ4mTkOjiwjwd38EV1bfubZTpNnjP+1aQoAVWmqG8x
YtJzou8HQPmp6+Xv7jZ+Bz0abK4CkzfAmdrYa2aYvF1bq9vcI8Tt/y0bCREAgsRU
lLHud34pYzUvdage46o7BKCHBtmZ4PqmTY01b2P2fkqUExOBe87nFbwNh+IDlKCB
CYGEvaD3ZRXyESGaORvxBfSTgBip9yMOsw5OtOQxl3nmRalxKNWrQArDUd1Ujdoa
onW9PUh/ssl8pnuf55ljRECulPH0mdabBScg0MZVLlc/y408/YxWJVSfJacy3QZL
YAV67MZqE9vsQfrtpT7dtKygmkVO6eWGSykSyEtjfPJu8r+TRDApBhHG/EwXhjd/
M7YZFJIUKK+edrRq4G2MHVDVyuZW1ESRAPHYJvvcTU4QGYjEc9Jh5UFBg1CxdZUu
xC8ktMrHkpi3zNDHWGcaEnEDjLB6bpqSpK3QWqcfmJZ4VEFh9C+2MNGxY+HwCUZV
m8oJ+PyaA/tb2MA4GdwcJIjZMq4iPWgQFxa8DK3//vTCs+KyfjC4PxGAXfJKp7+x
yoaJz9OTA+o/Lw6DaPC+4DCsLRlwtZGzSfhQJ97eROf5HrOSBjThen1/TotIMMHW
sDHXe4Sr7QBMlfHcyhL3e17K4NWtLMKxrNI53CphIphNPEmpi+iv8rPbHwxJnDZw
ZAsrVX25zIVdqqHJYwkQEYm4zusGk7JIfDXIGa0FHye0OiIH5Y7SJrz1WgDn7Ugc
lMF/3YU+G9daCQoexi4DF8dMjsq6lgPVDLBCIXLWrCegqYE7vvPhSIAhwqzo3Gs4
oLOrvb1utP6ChypDkgqJRIPOvK9uKi4NfxBzVo6HDyMeJr6AndQ5aw4y7N85WXK+
Tg1aSXLrSosz5f+5wGY5A00u0T3aaRVn45vru5ec2gijK2bgeW9Iks+AwcXRLjlg
JcWXoXtvsLdsSNuF4jn1uFyi/TiN8RK7hWcc+O3OgDvTJF3mVsAMAbmpPO44Zj0N
JnfNvknWBT7nF8r7QXmAOUGBkdCVZB4mX+tRPVDsb0QmsnQwcFtoGjs0liP+qtM5
fpV5sCU5/lWFtjetJmg7vC1W/6MqL/yMzt3BhH31yWSSk7sA11/RE37YImm0TApY
0PVJgkb7ab0v9orQCKxy6CU+f2KMbC7fL3Gdxu+tbPYTHPo5FlsxrucHzvUDRVPv
tltxQuDju5129+OscqE1mb93SUgOhw22rXwPeb/PuDQOg9w+wfQtxvXcxi0pmOJG
Hz1AukYPT1YTEfuWqtv3lVWnnL4ogukUw8kb74kZ/y0LMgFiMlpXAeDes7mlDYlN
am/YLTnI/NZEHZ3aPhzCwVS+s2wRRPCc7VW4DRh4Q5E+K2J/j1fq+zMWKXLjAqTi
apXd63EIHASLdyM8/gcoc6UtbQ5SKqzGmmMyLUSXvR0x9WATYt5gqV2HHq6/imD4
cqgkfbc84QZ1xWMuTtM4VIbaP2NbuHEwq5JAmpikuYSgmb7DdjaflxhwYjLfHoDh
esrmphWSb7AaKawLHAkIF08xYLWr2QBUuKjWD4jqi7qlKX5wIDIajaa31Onm+Cjq
/gLmUHcV8Cv+jqsBvScRUrFUTrIuKv3wRIn5lxCzf7GTy/HxfQXWqOiGiz93mrCJ
5yTzM1NkR9eaLbNmJJQzVCUMe9yt7bRxL1reUN046YwFvFZu9+i6eOqQ2eCwlfPo
79MK3gNolU4eLlSK732G3Ys2qDHpAVrZf1u215bTpx5AWFvLrc4ZoibpYrMbDl6D
6DIAy89WPQdvzMbKml1hnqxPINPG2G8ztgdXT2qZjLd4rGVK+LKsCmeb485QUC1/
bFGFW5AfeBnwncEzkJDC0VQYoFuWuXT/r0Mx8BPVZt+H9znllYKZtd1rfgcrdwa+
+p+QD8vW7fJtBCC9ufrG26VjfNoUwgatpZuJYm0CQ1DK3sGXX0rydH0mov2ZWagd
HoD5BY0g9sjoQbEOCfDEeuzZQX54ixy9F28NTC9OZ3kppOTf2hAUmk4+GIq5niqx
VZ0i0Ivi2x06W2Fz0Jwl2I7GRD9YDg4eOy65OyJT3HWRqxeXnRLfm1O3Smyh/0wp
PidcqgRw5CiG5e4VXKUJUu3jYGcAGL6pCdOYe1aFEte62Yj2jgJF9mRzQD5xaVuy
twAvGSk7azvYwyfzehlpDJdHRTQlwVTIUwFwD1tUSCCc4nGBHx5HYT87LymDXEB5
L9bQmGfnhgfnWH0/G/nDb0VK+aYO6OkKG/k9B08e+r3zAntg2fi1ONG58DFbSuA5
M67TsMVnxFJ7UFw3ywWII5nTbn567dr09+a96fMl/Mt+riU2DXXE0q6OiUhSj+1c
FW8Wn6zTdGiOm7Ofj6VXMbyoy7MEvVbtIJKoVq5yDwBYJ5OI2S4N+8k6XXMlCKbd
5qcyMEqhkWGT9wON/cLOt7CHwMcuUb2n/qjsi6jNwFZXO6x8BxFK7j38h/c2nctW
7tggyPXZz6mEw7LU7I7nEvFjZA8afrVSQZH2Nypms6YQHrnk4YnDb9mE3WnNelIB
kk6nJX+kPDkU9qDz8F6VooykDKdG5zCpJNDdPIyMZHKDWM9F1KthHPgKoq/VVkgk
0kaKhHdKk2stnF3+RH+5T0DLj50kkN/xSnIwfisOYLqi8L4l/wBQp1NX8nb6huBP
5YMEzkM1ohYXyH09w0g2d8f+Kaebuh3asoVDMuwdHnl8qxzearg4hyzqhbdIzgbT
xr4OjEMR5ERLXykUBjBB7xumORluQPij9kd4t8sVuPEQhPG/bzukAxpiEyXCAYQ3
46jxD5OFOpl9Qh6EyIvtauriZo2kr4bMq5JUr8Z3NU3LXaaKOfh86/a2oTiULVFt
fqCE04h4hOEYt/PBkCqhutqN+86bXdQ75o44XvitmvP1BHifTGRspxTaKNRwWc4N
Lw9VsJ/LTlyO02F+m4PpfKINR2cG+bkzNPQ9hAWYeqnHNC2a+cLkZ3XiCLIfcsNi
6zgWJ4GLeC5WaRDBw3u4XjlachkSi+UsGS+JYW1UZcnmANYvTc5mUIrdgnupRf5L
Kw6UoUTFv3bsH8jjfQfoPxf8Dq96BhUrZapTuojLHT4S6I2k4yPnhoxnqlmmcDFp
SBABUtkPk3DyyHxzyTwE43Alp3wCB8Axh7+CIqWwDsUgfA5ufFV4Iuo4Y3wTr/9b
H/g7DeOOYiZcZ47VFhlg+szcj6VrD8Mnnr7hfktOwIqJyLXmFKEEa+Nbtiyb+zB8
tT3O3sU7+/eX0tebFCpGB94ctKqnCQaxZaUEbl/XxA9NksXsnxZO6sYLnafXXg8w
K/qnnUqLVyRsA9pGos7JWqf5ik57UF2cvnfMrGezyAWGTv1pio1zEUitajCBGleS
XFSVJ6hNDohkfON2P2zQ/3hwXsVMjO3mvco/CH8ls3YKcAAB/mzEsd5sFTJW5ukx
btkBXn7tUSQxbJhZBtEof0l5V/J+PHnl0MKVSDE6wED1H/sALFDgfEIBIIXUw8Rn
nAPzl0Zqtf70tkQeeSooCFtIyq9Pk4C1FvZrKUCR8RAZqtFLBuIhpKpBtO3sriQv
0bpncoSzhHcd6rZ/5FUYZEu98AJwAH6I+CXxYkeTiL6bDTTJl7cm4Q1+TutC+Vz3
vCsf0N16LrIKbfL7WPqa2v0ntsAHL48VqnFGQvNf8V6nqUUBUHRS9KSf8cpr6d2A
roOQiZHlBYHtqCvSnWK7RhqQZ4lu9qycW/qiQFqjxbx/+HQKFCew4Ffxl5rvycLG
SQf4ni4d1zxyD8C9DNIU8CAow1eyARMgdvROSYKn7G0nxVTI6U0FULpKlMd9K/wq
ULEdLoNAnXSLb15Ri1garhifm4BvdbyXd4P5yQnvjyneRrg/XSbuwk6QHovgh5Pk
aJ2oTaKlXlCwh091hCJgepB6ez9GpRaEmOyqmNSwQ7HXY/NnbhWAUuSnp92lz9g2
o4vaUwR8Zyj4xDfleTJP1zNO94nsFZ9GiyxQoLpCa7EJMG2lj9TKjsqnIMs9wy+s
tvc2JzlSdQQOydPd6IWocSnp2hYOdvdGK70CF3JxmZz7CHSftsG3oL/SYYAdmazI
mJeIDdtXEQjeGS+qhfaUCXP8msVbmHwpOeK044H2fOiwpPCLd7F7FqenLWjmNqyV
l9ey+NwQOR7Zg2Pp+9xygt/92MucfkTzsPjrezEBiAOdtnOCMffe5qDoERH2NQEM
Ay6VKuDM42VZmgjTfa582uy0uWBimvykeN1ccA3WXnf99wva45+do6v6fFwfCVdr
jeL5oPMWhwp/Mna/fETOyqnzqRxvUR/AeijpFDM+Gnh8/NciEGofQmVhkhjClcNp
Hh6ZKy6VTgVnvO4hTFyIerY2ChdeI/9L9GlrQyG5jNCPDrX+yKbNBGQxBvapB/vT
mDisH6aD2I4w1yPvlOEp42FMN/q6vDWvUbKxSlk1VkYWi6PE1dHzIQpYVE6HuDYA
XNuDLuKQgi9JOcD9hcn8n1QiLm41z+b5X4T4WUL8ROHOVXPc4legSN2D+w/tMYGU
ZOosX9nHXfoIIuOIioTow8oVpEtw0cp0EjsnmebrmtJYC2c/I7v/O23CpLU+sv8C
JC1LolVnTHRWkA9thBUszMxkegfpjIDv7diEaf+XkRwJhVk7YKBGjY5J187cW8KB
wq3XCVjrCP9+j5W+tjV9rdZGjlzFMMLysG4PzLAMyMKqTfAVIXnJglQ0FuSMLEt2
l2GGnmkXiZFk07dQH5CEiCU7GBTCiqchm9r7vfcDGVXCfaeI4fGXfdyHpH5sT7Gp
2YQk+rciM9KQLhGYzlbcYWiB5oy1AuGiKS4D1SWlYgSIRKpqg6SDKzTEj35pM9wM
zTZznzfalB/e3A7mIUqOCYxrdUscxCQV/njhiN+IdnppjezGRyg4y76K2HyTXYNy
qpxb0oLNEtairMRgL9Xvr4sBVgzSAubz5lTm3t79EC3JE2Nf87ZG1NZB4LGbmDPf
TPfGZ9qJHvhR6gDBHEd1c4RKiItwu7frCv0U+eQyiE99SRb87orSWLfXiCebj4zX
yDCORJnbRtiEkpNvPFw7PpDgjjAIX8UVkcmoLMq9T+WaRm/P9Y6FJ7lowZ3xvgDY
nfArEOM+74fqQof92eD+5cxpG1oRq3XFMiL9Q4SmAPMDD9L/SK2wTi4UUaPVovcH
/PRMoBFlj2stnqHaWoaxEjnXvL/CPk36kQ8Go6c/MzYfkWkrIdo1ujrCB+fWtEqN
cFhHwoVUxZZfJ+YT7mBvOhDRqS4SeHVX4erZ5CoZducFg0E+Ye1IMmsauuy0ORSd
nkMMygSy0a1Iigwd5pTqRFe2xoqq0ffjyJlYYt0JXqKfVe6GV3N6Bfg8NST++gOX
nryJ53c2iiovONVag9fnicAE7HAny34nN74ceUx/BfmofxJS+6atI8wof0HBV4bq
prT0tN6+rg57zNglDqXoNA1Xqf9HIe81Q1bTv4UeYBhka4pCA00sbBSnQcKM3M1g
psRNfE9NGrudCWeNWUd/Gc2ANmwJosnn7m/YcCf/HTQg6Wb9Yll9OxFVzZSMC6cW
juwAuqZNmc9d1MLFpKwsy1xyH8yhEwPsS8dAgRwv6x/Re4Ytp4YkI9KY14JbUrWK
eF3d0/561iQ/Gq3SXZylHm423U2Pv21XdGsm1ehcoadm7pftdaOsDyVGyiV+xGZ1
CmV1cBSZieUIfhwBv6+i7gvUDLhEEGK9M+AO1C8nkqrJQwAEZm9q7mFO5zsGchKb
ipiE67wdG337REmmtcUAY1UCzBlp1P3lUGhwLKShoDdLz9AaGRxSj7XgGJL8w/tz
Vg94LHHPbC+cu0KInjDi7nvqRL85ZXKz4sbQGyBF9DxwyAdjGOHs+ySGJRe8Uaqw
jSKyQXh7jS3aAa4PyQ3hTJVug5Sdc5kjkhGbAWuCJO9zLkFx9ymr6mFMB2EgUHH5
1A7SMbWzVOhBXj70rV3pNSLd0EuwEOmmoQAOU/6P7asHOlFXbslgAQ2oZtgvdFhA
+eRm+xfcrDUtAie1+/ws29qaeDeyRy7/eESoiAD01GDpjc7lnPKdEVw9WbhJ45Cj
sgiVZReSbja35XP5E+qWpVo3pUUiX3lstZ4i0EhYimN/x2myOJ9/XpnGmyowNBWN
WiMGEkj6Muc1ILISA/bsKmRRFIcvUKiuHlBMh/okT1y3rZUKXzwuEKQFkopNxOsa
v0G02/N2K+GyNHGVYMryUlWgcfYVnqlzdtvNibP4dY89CBzElhwXK7oeBwaLH02N
I0Py9MpA1tBZYzsr5lKWu8DTCSBTa74+DRiuyRSYeawhSyAPHMGNcGjTrGGQjVUh
Qx/vq/D39nFY37mPi8xba/TVUgsW78MHWXtcAJF5KzXiBhFlplBnD2jfQh6BTvW5
P53bNGhuTkpYTPwm+xv6Q+l92RwAdYADH13ijCDyi1C/FClmmoVQguInzPF6JCX2
bLMRH4Pecx4EzWqGPTwmVhpwFYZ9mkeLWCKfB8lzUAYNnaVQdLa9UtcX7hrQnCSp
4AF/tGy2fODG9b7CpuxEyJV+hQP1ru6dIRIpgc6LRobDw9uYeBZlL6qujdz5mNH6
CjiBjvpOwz60oMAdqqy/V2GKTy5foBYrEa7jUI3LIcELM+4nOMynETxOZaWoIwIT
Xx8UkU54TJpGWKWmEZrVZONQyLRm3p8AF5WwBGox/hThJUXlOuPb99EVFmsvHssW
rUftJpvVYRngeV1bSpYAnnU9WL2SAcg6uHhtqHnD/o2oXm8Z7HifLwgqEHRLKQdb
twjDCkcLPyGpIEQn7DA70YgxxTmFoAeo5nTPgyEHwKi2gXxG4EPO5i68qPN23dBH
fbGOf/h0vasI+B9CNQ61TX4e56scy2U/o5BQ/k6HHHS/4VNyOio4h6Z2s0oQYo/O
rTYB/Ax7TyjD9kFEfmmw3ijTY+JPNEO0ZSUEPHML9PFyu8scRrRdkEikR+ahjE13
OgPXRfsix0dMgsJ39NKvYddpQpjcpGm/Xsbbamsra2i19otBZ8J1Sq2ZfB9X4dTi
hIGzmtux5A4lT7elDFM418VYD3h7S5vF15xtKPRmOOxmSOU994kg2F2t29AC3Gye
OJShDkckbWP3Wzwz4D4qQRtJAA0swW276Ku5DZTh99B9arAFCJ9AGHMdjyy0gyQm
hGRf2he+ZDe+gq5LQAKpbReca/J3le32s9eQljmac3orQvX6c1O/eUataucllKam
k6Y5goQ4ilfeOQrG91kkCmumDJSHy2MKHGDESAmUfrFqEqxtB03GIRzzTiYiRRy4
Ws/56DFF3cYQLEnQ2UiyQf0eo5D+H03N6SRTczl3WztkG7n/E3vhl+9F8z8c2HHT
fklWMQg5f4RtU9qVekOwXhq83o6ls6M9lp5/0erFJA24EzcASrzlbInHZnPrvpO2
IXbavAxtyComZM9NMQLkjJdp2zFUY3mreG41v/1FFG5zUpmug2yqKaAixKnLSLLS
oE2CcPRm6/Et1VuCtbWx2hdK3lBVSfUx+1bcTqyBux/m1giH6vkkWqWzY4/G7uSw
XRvuCWraZz9wnmhri2fx1rvfveZIqN6FjJiZFFXWXfTNxS0847oiv/VhM+O8hG9r
g6dR4wOkTBkOhlxOcaBCsgf/rZXC7wLQOEl5VXhJzCL+xxz2M7ShzKVuYh/NukKz
VJbUtCbcXhPmRV0RBtiPeGmDR0iFcw8nmODqVmO9owFJClucrhkuDux5dwmXd14c
Z50bCy/NUODWxe+UUh2ckfyZzrzJGGoNnCAD6hNnIEfl6NYUKoZ0tCSXTrE2ayOr
83+7t10vg3yXn1ZG+z+038flh2pOJeywuEQmGDJYcu52DIBvv+lE1mKW215Geq3d
Wao0pucv1xk53ZIVAeltX78lBjOdcFnzVzb7RoEQi+2jEZWgfsNmDzLRxW+H+q92
AkAA3onzMUheMLD20Us4MgWKbmzkKK8x5y/WvI8eSWsJvamaVHUa8dPaF5qIfbWN
ZJH9v3TEGQfZOpef4v/DhMPUc77nfXNgEc2T8drftSt6hJtzERUdmwv8i+V1NNOk
axiK/yps9Gqj5s+xAJOEIj0vx+aPRhJKmOf8thsXwyf8qXkSwM9j/3NCDTMLaYmL
tkRUmyobszRqLdTTEuFllbZHk1kTgg0AcoCyZHBepmUa38RmCB+zVzPFH0t0czod
4A43nv1pe8PrVuMK4v68czEDgi/v9N06bOxsjUSiXfP/7bZ3o4dxHyDk2gnUOPL8
Z5x8SIP6A8PSqgwn3OwTdyrkHJjtU+dSP9Gh4NYFBCQ6ELq2MHH3bc17bRLkysGz
30vT8QaQUdYGFBj/3UXJR2n5p/HHFvdOSDQSPVRU6aI5dYoc7pWCIms/uQtAcMex
mFCbECLzo10HM0I/JNGdp6AuvV3hj/e+Xe6LImr+Abb1IGYlIBO+zKp/dSTdPMH4
Rra4RWvgePnN5eI+2jA/kANnOZN4PPkY1pbTz0CQgDiX4IRmR0+t39wChKv+JjXL
7ZfJlaKHeMVUQ7m+FZ7AM3wWiCrAXHmcoy2OD3tASgJ0ftnszwZfePXgtp+O5Ygb
fSLUfgXiA+Ssk5KS3255lizQ4LMaG2LgU7QwPF/PRC5v+pxLNCgEwdMUrNEACbmw
nj9YReXRS8TAlvXDTj0htN6+mMBFEmyJrPh97Vb3RqozdkQeAqfwXb0+s9Y49Pre
A7PRGsvBH/hIcccWJHgCCyF2TS3AAivLJL5YydW22k5RX8Nu9cxUbx5C8GV2JyXG
XyfvrwWymvukUdnqqal4MwJKVjWX416dL2jTD9jEPZGZ6maCz3CFUSepZ5Is7PAQ
/XV7qsbMBCXVfrqGM4pkXf8Kn7fuQelFFKvWoYd8IovmNzVbkZ/C0k5hdv8+Pe71
Nh0OUKzAyHltmyE+RAtb9hxpd/6Fr0eZzd7I/jR9b/n+AHTSOnSa8ehXZKjxNovR
AQ1gVh1vUyb/W5gOcsZSiv8bpPhpo6xhNBy9vgTp7uqXufUL/60lBoNXMdcnTi5f
9mIKkjshaIH29SI8MWUbuloyeNbz4j+2F+iH3Pc7NOavCqId/L8qqat3XQMBFp0h
QmYcaiZBXmvMWjrxFVyDfjBgt7LRvStd8YCRMcuzlfGkfxrjA+aTM/hiW4Mpz7JQ
gn0B269OdQDzms40j/VsP5yV4b1XbK2DlTsiMlilnbb4wBijcI66Di1+rxT2/zfG
Nwm/29Pc3BS2FUEmwmk060FLxT6luNH+/lRf4ItnwDV4g7UwNGJzF4/xTV3l7hXm
pJv4Xu6MrLDDUtHXjW+sxTJ/ZRI4RZQSrxh4qg6cMmozhfJYbTluVzgyeDiioOJ8
BZH7AQJfEq49Y3pYYCVIR1fJ/lsioJ/7R/HuGeepYClrFbsiRhktJzn7TMBFU1MA
McMyiOJrwYtELnoczKwo586f5bOzeA2dkvsCKvsxB/3dCN4jqV4clOOKS1Zaevze
cIWrjhfyvqngD950mMUJRUcZXBhBKaEI+6+xQlxodeGvycWHX8NfnT7V+cMHJvqB
RlSgXfKUjygCdZfxTQlyg8yeQZriMqymmy41bF83bnqcW6T0PByrmqrC9+vbTFx3
CzkG4WNm4vYK0BDD2mQLeGKCIPJ6uS1NXRw9EjcorZb7F1LzbrYBitcVDpJBrbq/
W2I5hYICt5YPCRF9/XYQTSnNUzfbJegNcI50VtWr4fdKqVGZwkgcKz2tO7ymZaqa
vdkdDxAFCyJr6ogii5aGkcSkm3tFbFQ4BNsZATr2IZmrz9dGHYQFHYIT5Uhq75pw
jydkqaNKCG8rCFnbw8Q+KXHz5OnX0lkIPhNJW9sqx00iTZ8wFrqrVItF2/Y6iCzy
5St0En9SoGQSg1ol256LXlbkjTtzpcTSbtJzEJVGvzh4jLF7uxyjHPqwO6xa5c8K
37vZ5VR51ez1zbdM1pEVO0dM0TlY4A4W98tReq7gBgmTqsv3sTEp3AWchTjSACPe
GCNIUu9sKy23gnNDawrTn75s1uPOoJ5+ijj39nL/37tmRbQaaCr7fbhNT73rLA7E
R1JJVcjj9ss7Fk2KjjKq5d0djBZYt9yXReC4YtsX1VTRQY7fvzUZwbZPoN8EV392
6CgyCArmNTRjHk7cxFQGHmAWV06kCVKLWDJfNH+HpqdXyb2TumCU6wzwFW/E2R51
xYLajy6xx8DaeCwLp2ObVD3IaF+kO5ZN4W9Pfew2ZnQ+f3ZLvLefNNKvGjnNyM76
iE/YDpp066qEckFM3hOhlX/bAFCH57Dcng5Ib+TgMQCatjAG6IVGvJGVkYF4N39P
aSvgQa7DDMSK1pvDNvoZz549nNrjDIs6Anpgy48/i+kO+wdcnNWK5Q0POxlV0i5s
dEmNvbozQ7cgMMgK14A+Ob34brseDr1rAwo59L9dRbcClRC/UOtfV3KfB0D8L+Ow
OM4odj4T4Wk2As08EoM2jErah5ZJxagBddSggZ2AVNHULGyK4HyScWmrNxXG6PE2
fu93DE9W+ctUJHJMcEOQSnHNbsjsQppcL9TElmJh4QoK2SN0ux7rFwufgMy02c4o
Kzolk/bcYC/ZqzYENm7AsWfHvesqVS+tShhm4qiFrxc9vO022B6tKkXNkFsTJEu+
xKGBW/8CjoJ6w86oudrOTzUw+nRNX8UXAXF/66bueuUz5ipcYJIASPXjqPqR7uiy
vesOaxoc/f8lMFPbG1TYxDMI9fGzj8CCEy/sFpE1vjixB5vJjhERFTSv+tsO8Ukl
4FXgm656lMp5lSMvIA7pqGHQ+IjozFh52EPwGnGRskjNGJNOYjgMES6YN+0Aw668
hauajUVHSA7cdZce72txYDNf1nnOeuDd/l6T2cZd6UyVN27tc8jE4RHxqIL3aD8s
uIi6oAxhFyJwoo2gaw/EcOJkFWcqfRnUmHHjxVMg/Gl9+8tctSGMEJTdk4Y9brYR
QlE/427nrquQKH6JIrrhHGp5st38HVyI8QFGYvuMDR6pF1Qs3LSxJn+KhqT5ZLqM
UTP6D2OdBkXanXnZW9ibgjgx3AumbQkr6KKw6XKoXFSGlGQvWRuysstwt8+ad09c
+DPGmjbK6+tnCobe6vVTNAHvjTJJHzZw4zEIigyjd7BdGroz5lMcbvCYOD+8cfa7
0PdsI1tLU0A9xkB+gNsS0N1PQCmgM8kufy3CrUL81ovudiS486LvXGkOqxzZRfrZ
Q6UIqqqqWw3Skc6cCdHH6glzgZF7BGKWc9o9C3ffy6HC07lTOxoIia214PVsx56/
3lAlYpp+2uWJhkp6/vvKrw7ggP3XRzGzs5IgPuHYTMhSE6EjR6OqwzDA74x5TbSl
PjZl1eVH/nv+CnhF6mWqBqCzdUoyVPEAPTRpTOLjZPnVNOPErf0kQmMKhTlyoBxx
4l9kZlK9VhloB7bBO3PNi2hCyEfEydQ+F5MMOwm35jbpv7hdpbhKjkHQVvO4jkHi
TZ5HLFDl3RUsiGX/rWoq+OH9cIShGarR4IvyDblVk5E84KU+lksbDeVcG1KIMYU1
ekKn0IVVPHdbXKLFBS4uVXlTLdd2K+A3H2oNWcqEj56gEaF4jN9MnMMR05ZXFhx3
ZM8cUZQdqcl5b8iu920dvhGCMLUTJozgL8x/ltAvM4LQUsizaO9fZFbeeYyHxsUv
YcEbYyaD2h/D9FBbb377OgDuoO9IZarHVtDdn25CBFMZYJgCDE5RpJXatfLlrd57
S6vTkEB/vcfxEWwfwJC6ynuUfCkOaizohsTNirHPZ98ldA83eeqeCVss+nCIeQG7
JcZwG6/BNqCv1hdrYkGiVpA1s5fcz0mRsbPabQ9BvLUpQN+Jgc1uf0aNiVdaIlhy
eLp2CFPXVz6WVEkahMbYK6rR1X5An1kQxoBeNhzURhk03uuzEc+HMH1GMc1s8Hr+
OaaGCUy0OCxRypVOeujENVQVuDon3vwJi/X/i29dY2qhSQc/QX2b1StSQ7zaoHf8
sVvrXz2pvwSJk+9FDM0FGUGKDfXylqPoxkbRjAQzoa5KYoXPb6qWNGAY0kt8IWSA
Y/geAy1KDTZNDsvyctfnSOISSG3xWhNol0ECw6S2cV7v9qtKej3uNCtDvPUrtSk/
s/zIi8JlDZtGkpwHJusIYgkUXvo3vK3On3M31c398XHgJKFxrriKYoEm/QW7LMff
iDYeSVXdEBltZa4zR5Rurn7g2nDKqONA0QTdDi9/pqHxBAgx61051DCTQLFDOEF0
YDcBxmicPz36GrgViFk+do3V076/QNuU8Sjd0p/K1/36F8DJECUWvrlZY7PjPlFS
laCY5SZJWva3tapMJO0oEHMqDs3RaCSUhe1VTapsCESaKuVIqGyv1KajCS5tQagq
Xr8dGKJWGIQvKEcZr2dYcP44T8qdPezvu5BMo8QQrkFYGg1/AJ0M1kqakZW/G/2J
lJI2iry3kJmsRfzLHzMe6fp5RayGF4bLzfG5TFeAnRNsEZZu+zjQqHK7vjd1pc62
aRzxGDxoXPVj0PwH3y4Wi8Bd7ybSynJphpSsgZa3U1h+3AuDHXcRZ6EZhAY8a+pc
cyJ3pU+gqTUuLS1g9QPSjbLL5kn4oWi9YYqOVxt09epTG+cyRJNzAp4ZZhMG+43S
T8kyb4SA4LhWI3NOTYMnk5tuk31rMoF2P3VFdL01oXnTHVF5N5OAfhp6OsAlm8sq
matxVQMJbmdPuOxLBMeKM0yM7tPuNUgH2xbyvhqmXagCHX96Be7de1Sb5pFmPGqj
0+FeV456tA2eT9xO3ws0xdq6tCMJ9at9/rkIlW+KLHLnK2jZvgRdSBosX1sdQA5i
Lh4IwruvLxdMv6xUMgSdoZJqHQS5nBODKHLnjHAqcHGA7lZFaV8SgJ9i7c5LU2vE
sOaviueSWb0H+YqTj38S3CnunuCtDOCjmMYMENkFEUPCSS9Pllti3eCOjj3uLbu4
v0KJ/R2IHwX8KUddllvkHNCD03Og+B74X8EoGHgOk1RhjNsjXgX0UF1laOVl6dUZ
OgZDR7EBQVyNdR5bW04/A5OwYxY6ejaae9e2rmZkZr9BP+2u/RwfxtZH2poQPHi+
SjcxvlXKsQ6Ap5NKvDlYnAG2pcXbdUSdv1romKJHqVeuFVyhJZLD0MVqVCUsb1QB
XynF7DKonDaAy4IG7nadcAyjDBK/8SqvTWrqrfmCFrYccH1q72cnaMvbA66PkZNa
XamqmPT9TBHrDPJo5viBruC5ulFXzrBEh4IVYhFTeKa78d2VDJSRshw1rVX1Ypzw
ipvmKHdMdzyUhZaYB337Vl4Va9zG+4jG+UeWzQJhjSrFwE30PStLz06yzeweuu0M
0oSa4lbjaGDMYojx5IlK17K+LaIhiVJFwvBAcYt1+FmgcbOwYjP+qhUFan+ECqjq
VMhJpJ9v9S4FUlymsWHAmILK60C2INJOLQ4a5MWZqjXFkbcCzgkkqSe2NempYh1+
mbTuqafgZKlqUadmJn2rlViY7CWHTsouuNNjxGfRZMpJSoOhhnImhs5uDydZZO+1
t5nqwX+Ih7Rbp9KVdGAa/e97RD0b1OJgHp67OSan7ynBi4um2naiP4drrvsXRECY
VgJ2IK+D0laZpFjmpcJEMfVTYQ435vyAMk/N0d790+Mya64Zj7L2gfxTKG0vBHOt
NfkjrjKdUuEs700zTtpre/+pP3ad453R3U8xkv+tyiU7NHDANtRF2M/4EgvnMThX
1bNc+KS8ASG+gSRlJ35X0UGPpiyDVPX6nONJ+fzfnlfqh6HfA3PNiHWvXBdpbcff
ksosGHzbbrQ/2sSoR4TFPE/2yCiz/0ineSMppZNq5etEvkFPT6paZpwzDrQDsyKP
WnGK8lQz5w6zca2nIqbrtikVC8YKUO+a5U11/bSXnrJCmsUENDVMpwJiXqF+8vx6
EDMYrUHaolxJi7xCEOozhuO42EqWfWsnLAQQHFhZfz3azRuRSWV8BIKmVctjAq7F
HrIypZ5r3B8RK79ofDMl5ECICkP2RN0/6WUzHYddskSrTS8/kVeDy9B/0eH8FNui
rYx3eJi8FclzCd2GoyW10Vk0D0TmEyzvAfeOz0yIpiRpMSnXIyRjMkAix0s756Ty
28qnYQ6O67FfEpBk3GnhRrU5HZJHYynhbF7WRDKfSNb+IHfrzSNZ0nR6QMU2St71
JmADu85qWdvoAaP0vx//McUgQv2wjl8aWXoZaoJQuh5jydk9q+IzWey6ID8mu8ER
ACh+7VppKy/1gZ4TCP3xI47mGqWn581SBB5/xKbjJrS3kJUJDlcSPYXJ3XuQeFa1
aWUC+I9Mq/hx7+u2Lx9fh/RfohCZvveltMgKj0lcWArCM8Ymj+VPLTLdAIxBAUFO
bDQnzP2s5ObPggF1hF+l01bD9dA7fv1l1jSCP3VMg6ZyZuccrFlQpqMHxPpYd3+Y
iIzoGNIITU/SjvolrflSIJXUjeCeY4jt1xwfzMASYNjThX65bCLXF9Ijmq7X9UWp
9ugf+uoqPUtIypdXMnHLOcrBwKx3Hlhd//b7drfHtA6wyO/8h7+ltBYix969ecwI
YgtbH7eeCLv3v7U/23QG3gJUecVrVosJaVSj+dCRKER/esvvshCisQ+3LfWjM0v5
mqJrIk1TbPsG99f2lZNfFm3J3i8yanuE9LEP1sDQpLpaZIAcZlVIAHYGTfjY9d/v
H/6ulXr3IlNAX3aXoKyd2jKENxNCI9f+cVU5RfhRNDVKstEj+8k7uPEw15vb0TeU
sqBuqzEjYz4yN2LXQO0U3YYeAPpPxf1HnW+exLF1999gjW9cfWs0scNSXBGenGV9
BpX4Sn9WFcJPL2s0b6CuZitsqKPjWbjXA1t+qZpih20zZuPNG/rKxIUhVZP2rzgr
1KRZHToSr1x+wzbyqONfkSDmTG9wZqcJ9fnNurzL6K+Q6qd+fILLQJT1b3rJ8X1A
aDbfCs7ZynFX65V7/IrieZu2qkivrr6FgsXvjewD1lMWTUQOcZNlgjzkdjGCSG1u
m2oEMQhDwCbCtFwFaT5Y0n5bFvcIfwgdZAaXmvk3R9eFbyd1/vKj2T1fgzGEfpMq
hRf4MCudaqEDRqMPFYW+pZPzvMf36yRxloB1rOLNYdMeCyug2/6dJYhk1SGXd61b
5LuVfk1vUw/FGiMANGyb0PVLaKbEhNDwUKGbijlUHknQVpZIzmWIH0MfNo1fyqlq
6Y+B7x6vs2p7p1E56sOlFCu3wBBlZzeDSFfHCjD/kTb2qFUl11zDB4tMSZOZU7/X
xAvdCCkxNBWtXAgRKglt3bwyqDJKlnrOYUvmAnfKIcSm/3VOuwXdX0ffEigD8DLo
iP/LT4zLUX1Q+ilQZSfug6FvDTclpGtAvOVtGU3BaEOVvJuR+PqNU0K/MIr3QYzm
DsbgMbpl+JZ/0d+iesYDQdRmZLHXM/SsDdM14y1z9AX5nw38L0OcjSw4U22bKDv2
NUZh5SmJYUky/20mB/BJ9mU7VAaOsO/h68uJuWYPIIXrRYSHkK7oOxecbZmm6wBc
eJHUf1FJ5fxYjJcz+ustO8/IIJoHtlmK2A2shgDNVyPdFyLgo8J8kOxAAGAfNWfI
ggtZt2BQDFtaMYsV2a+6JrnyvBfUoKglkyE/vMxWvx3mPinf+zX0gvQDLwtIqjRj
HWoBva3HtpzqXSyuql+Y8TD2WuCG4jHyxDeDhvmKDHQkVYUbY3TVcNI0UE0E4bLb
F3xpquKvsyQ1mjYWVMv4qoudaswNkb7wVBS2TdYWzhDF41JWEirzO2DujqHT8AVW
z6HDCc42Q3BiQYpnSdb6ddKIJwEZkAaZ7gMPKiJB3568lYFgUs5gpNKy0phMLc8J
xw1MGuTV964TZJ/SNvAbsp10XVGINuB+6bOcAMO51TMedrvxWXmjBhyCPCY6ku2y
tetL9SpKLqLzj2FQ+LCdOni3Jb04DxtK68QjcSLQHTYo94ls6Q3qkfOeJ3kFsCMX
yZ31sN0ros287Tqp5Gpk9XFvRQVmVvoYOgqcKbZXFGlcKpsg32bwEaLGTtCoYY5S
+S6nTWCgZUhjFSjC0NsF7TwYVZLrsgOJ3mLfGqCX0dWgPwRTtjSlbVcz1MufVxSv
xAbpTDQuUyLV9OGoSqjWKTNs/p15avyIIL2xNALQehthta40YiwopnZs2CqXLG6f
aU4M8D+antCJu8q2dLWgRxQwjAEPfS3gmJ7Ke+Cy+SX/7ZV8yZhfzBNwo1fWCW/V
ZmUJQBremSNucJl1FNT8jh2v2DBTO6affMpOnc+cUQN/vV1xQTjZsM0dZKAby2k0
ywfQfn3cVoCwB7daTENXa7VAysI7lofdtZJuwVw6Qoq4x9Dz0yeV3LQ5yyoG9uCE
s/rcns7GRcnx7jENBcONKf5dp2uQzxMaDu0sDR0fpwnARBakRg4nu245xvxTpgaJ
8K4i3afWQ99MZDntxOscgXdgRAvHtbtVnjtxSqL8JWek4czvFlcmNKLe31h5oKXD
yeRSXWI5D0d9q446h7Fc8d2p/l1FPGHU0GGuXhAe/Tv1YIs8gTqTs4kO1bawk3eB
CrwIGU+M5SziKv1vzqeK3dKH8OViKzKkyFXWiJlX4JJRritcMIBCNRt6r1pi0+nU
imHj+95BOVKmeuVXMeWY0Gc/Gpl8ce03D6YsgZFQuE/RdRUaxi9h1exNuSS31kxj
0LcWeY5bO+wj4mAtX1Qowt5jI+PjaJIrCG6suRUwh/PLI708GUWKc76o7lo0EYWq
uhqEehLkzadrRVja3C4tsHq60xzQeaepRnLJLQkobMEE/NHjnOqoAJZ5eQ9fCKRW
9X23DSroCT1RnisrSXlqsR1zvx2o7lzW4USnk+gQV6mTFSJde54ivtx12QtdgdX/
kUUiGur6zYVDnFPgVYhFI/etuSrcxfOWg5TPeBKoA3BSFFtPijv0N9pas/ez/wef
UE5+LRdqM4B4aJeGt0HhAZid1XnTVQBQd+3B3bEiDi+hY0Z4lUptJav6ju64H9M8
jlY44mU64ZX5jIOR1d6kaV3pAdoQ3uSfP61J+k02T7b5fg7IoT/Ncky8dWPOyeHz
3ivzAOhJpM+7S+xZL5Qf1t++IGsHgM/CB6kmGe2gHQ0aawPMmuzGT1J+RZQU01ar
L+7nhUBe6kh03B13DgRnnI9axm8lMjZX8mqbVN7jMKHnEGKPwNkLUy8lWwcASzbX
UlzRURRgmaZZeoJGY3mDQS0fZnQXwXbpOnMyAnEiFb9/+52Lb6nZLglwhutqj4+j
Wcpu57/AdMtoGMpl3RdDhIMovVn1tJYC0gy2gDgoz0yhafsCh2AGo9y388T62oAc
/XuaLq8OYZKt73Kav77uRSQ1UA6XhHapVglOXE0t60lZu2urWS1OknIy4fbRlNgV
5K9k33Fp0YstsbWuKAp6jtsyW8pvq4ZGp5C4FvCyTYG1I6ubeRCabNMHIkyQCzgQ
922dtBzQuvYxMiJiAvzXyLc8YqSfphOU64P0lNA5+yBo93UHXo+DWQ+Ocmxt2A2h
COVzG1vBFs7A2gdYgp2Bu7C4WVouN33I0wY0CxU8MDEiKyPdLh3YqJ49tTPDc+y2
w5WEhZlTvmK9ZU4U5YYMQRFaPXIrUnTnl/xMq8mpEYAsQGZ5K9Q5V33EL2zoThC/
b+NYWOYjjVDKFl4HLuVDlHsw+EAOximF3ylTaw3cDzd33haimIyQDsVJce9XpEwn
2ie97KXZCLPBjpum/R46h3Q/7ANCNz+z12Sbr7QqUrHswHX3LdQdqJxIecg4Tepq
3Y9DikgwSEMIwKInvu/wppb4BwbUqCDi+IhLDiYFzWrKvTuUgCNIZ869z+SSfg1C
+EFjxydRCTBtQhiCjHNLCvfd408KcXFH9q2F5XzeXE5QvxiAEZVS2O2FENThuI+c
VR6sox2qBVKf/fuU9kg129/hRAK/lwrrd/rjj+fpt4sRlB0AprS+VJIMRIAPXPfx
EY5ygQejOZXMFK9V4MeGN7j76T0t1os/mO6hfFAvuASQDungxDH1rYOldgL4eSt0
bPv1cYbq0MkCvTTvKI1DuORqcli9ekqFThf+5N0uSumLg9DJkgchEa/VCGaShKIV
dPZKmURMoUI/bPhoCz3XO0NslzwaMMErWJOxRuFdH7+w0018rSBOjoNHeg40HQE8
0XuXMOAejuOwINkbKHcLpUL5m3ELvrT7dF3JsxncQJo5B1p8bRZui+AB5lMos3Q9
x9YPmEN4/AaTbZTnBtaWOo4L9jfvzbigAXm9tClcGnX7q004enMBWMei7mueJEL5
OYujC93Q0Zd8p4CRpICBkO1jLNkLN9azWUCeIObcbICZlJjtxlK8zn6y1N0akBCo
fcsSY3Hmuj4VcW7A+yZ0PDpc+dVv92bl/QgxS0C7WhoI5Mu2BZk+9mbggm39Iohb
IrI3up1nNYh9aDb7+LbUZogzey+a/bU4KyEomLgSshuJtOUCcrBtfbgjdIG2QPRO
KItFDmwwyHPVICDKqTMrfvLTV8JDPnxzrkiu9B19+BVKDNcKYjETlCE8IPO3tBX2
TBFInW4qOZ5piRZALmg2t/uW0ltsFnkg1sXrtougvSmhjbp1s9Q8dayfApSzUEbs
GJLIJOC4GQ1UveX0WSIUzCYWroDE4NfbbWcIjNAcDICeeWQ3XPHyRELshAaaKUYG
IQBw4NL7N9ResCD9el//SxPNMDtx0LXOy1LChAnb4Vl8swQzdA2AkTUsHsgURObl
YcsDaaDCUvzfKMb06we8KkGcaVD5oDoAWBNbPhLWgZ1vsTffgTu2lhatR5rYkNpe
T3nlo+TdQgrKqUxfMwD0UPb5GbgSSRD8Z3mF4jGAqg/gPgtE0ne4Ob6LDH9P+Cly
nwykHdLi6ncSFqGx2P3Nkgnw5+J7EG2gRZ3mrdOvWDoCTbRnOL5Yn1ObsP3LXZbd
1Kx0ZPtuCgHH2t3OASccT5RTSNnp+4E2FgnYrD2VP5LB3++rpD9H4tjT0ts6BQk9
LFmbWi/yKPCHfXs/UwnsW/W9JADjFyulwUUZAwr7UFToIjdLd7+zFB8hEfamYb3T
ocr+zM5ZvngMOPweIO8DdrbHK0KQbZedGy7mgo9pHK+PJ8V1rR/W++acoa0WdDUI
jlpe54jvcYJS7ZUWYiBDqCPXW1DaZRLF0SHDio2HDvYvbImJlettw8adKpgDqjpD
GI3+Qjl7dJdp2u4IbKjUGQYji27Bc1gU1gexUu9dfQWFc56K+oP7x4QK25kTQHDE
os8UO2mXetBzwKUHMfsLmxyEcWpkqXM9muQZeJOJ6CVKWne9UwVOOX2A9vtATF5h
Bg1uftUo1EIOeHA1ChL2Dn1fuzYQ8QN+jQc9/B8KGoGAbVNoAkj8J+ZVYjnSAOtm
3DxOoskbj/rUG3FYaHYgLJGzBgP28s+7f86iStm1d3J0LydPVtvpeGcSx2wlLlkp
87MBFOOQ8gpwCWWvkcTGzEQ150Lrm7otVfrdAvOVFDnpc3B62Dyk42lQRhBl02B5
zn7wX3HyHu8Uk0L8uQlVvqWr4cJXkYkH9YB5fCFl3W1zGfEXEl+6/lG9whqKCakL
za9fzZN+LO3JdW1C88kiQaT6yqR6+fCVqFkk44xGDMzcfWQiNMs6cBPyvbdTD8DH
hjCIkUoA0M9PhQ+5o0rK/XQ+wDirC+81hHfDCXtvhq9tPgIvttz+pMJiPDIn8sv9
d7hen3Lux5xXP78rEO7sfLGEaNNhHRJ7zENHvChZAnQPQmj/KEchx6ctns9R9JUC
zPi1ufkQwNehnwd9LRDrdYWYJ6HMgE6ug5YvknEBHzuIX0MLbANKeG59VPJ3xywg
oPS3VpkA/46VTlZ7cLrA3y8PN1DYEMYb0rBjSXqFjCWU+b5ntVKsQIoaCq6y4YW6
eI37HmSyy22NN8sSOVkoeTnnBsKHt6D2qbb8gYScP/YBaiABrjfJWlQ1ACUvQcEh
42PhUEmKCb9tQViACAoN+86CAEPuO4vnDmZsYAlK63UCBd3s+a8ByUNxpvASos5q
OsznSbMZvcFaWLpekL+bel1K6oNHN6pS1D76AQPzo8koqQGwU2XfQx52xT/NBtkD
ix2mrn2phHnwQwkyRT8wVkJVf730hDymQxUK8vCfkp0zunYy3e8UDLekA0VrRR0J
CtyAyRkTEC/tvkIBbDXCKbsVgaqNM/ahbZO4cF56RNl7VThXj2B0msfYmdosAh6S
Mm6Oki7MgppqGUc1tDa7PFYDMiCzB7F11EtVTfikj5bhaVsu3ogBTvLnYZ7oCDU7
BBJpqoE0IzTt73hElAUgUVC+61DT7Ue6UfVmXCeq7/QeGnKUf/sBUoHpcD0T3ceC
zdRwZd/OpsbojHWJ7mH14eh/tdCbRLXf1T/Wlw283+yJRJ5t2FzEICIcMsE9SuFV
DXsumdhm34N2FMJ7FpCU8kom5hm3WMUAlqHlOcSwI6IUQ0UcfP4dDGJdto+0ARNH
c26j4xFutvz/HkxqdrlPaLI6+nXFYyRVKYMWcp0F5CVD8ScSFmIHPn8OlF517lww
aSw5xGMRX5688c5r962EwxT8uLW8B5nl88IIwnHB+33NwhlSQVh33oDAhb62R/t9
3f2E4MFr9+U4BlU+HLPSqqtWNKpj6SLJk5q/qjgqflI4wkpAczrwzG+JCWXgK9t8
vZT20WrkkFoSSKNRmB7m3CPl/6hY75pE83hkRaSljATREMv5z/fDdHnCggO1XWcn
PGni8yq+aIy+5Ly0KnvcH545Soe6VHqAiqKc9eDFOKBy1yLqfoonv/syokzeR5Wf
SG2/tLbGjYAPxnc7AmM76ZNDfoMLdtSO7Oqj+D1MpQJdz0NdBcEA6PA8RuQZbUWk
EMRCJaMshQAAtxklR+0kDc41VzhCm3+bAi3sWq7M68cg5TtRLhCbfAL9/iEVXITt
vut6SCkOpynnbmRD+YQIZH3mHXKp3u2WT6AY5CKF5/R6oPbwr7HC/RaKcoAGG/Is
uqiY/fv2x4BRv+QJBO7xDjE6SsnujM18h8rkkc182vCiK0lQP/0RAlliRTKdajpD
+Etssk0n6AD6v5FStemo6nMwv2L6c/n/+2g73lvoOIRMlUIjPirs2jVlI97t+vBB
ev2QEH1eQ4lgzX+kBipiKiYAujAcfjZnQkpkH6+P+6Xeqa062z4nRvevkymXAEvf
ZzM9sj6sBWkmp5KlqyU88hU+m5/3SWYUoZWI95xAnKnBKTTpbBIiEqCfUdqPjesN
iNgzjnUJ5vUC4yA1rv0SgNjwEoJF59sqONvvSyGxfmv5tquJHVjurg8Zrad8kvab
uGke8cGxslh57AabO3NC+2TEkzxW2JKE6LsfDuE2YC2O9/e8opxknCJq2V82XmEP
l8fSgohnXFAuhc5pnoUNF9JIevrc5CTWYEQDWPT4ucSNrIqF4SWOvvO3j8GSKqb7
stoMlThwkp7ZPEW8oVT7Z5Dqn30+jrW0ZEoDdA+K8bSHwf5KXeY5hOE5FfuU8pSK
3NjicMXrF4ipdMPcIaQbzXhuVH5n5HZNCuMvqvgZRTC3gLQKtc3idLyMUJnuZvzE
XiDdcdqy6Yu9rC1cuCmDyvN1emYohjO4SETocMlv0WyoiimTxk7AyRmflKS5MpwZ
91RSK3UCx47yhKlZ1n5cogw5OCm8c7C4c6M8UW8hkT1Insdg7Tor1vl5YxfhwE6Q
Lbm+F53Ub1eAqDfOVtvxg9P/w7/hfS3SpuBx9ID82XpKHCywJlU1ANZn1R93lYnO
84x1TwPB4RlWXUDkRmT4nz2mD6YA3mGyNRloUIhzAKYsty/lSHiAaO0Z+0WXSHuK
vZUVxyLfYKPcKyalRgv5Hth7d7mXYZGe6v+fxuZ9dLuGHfM/m3mFMwnbRps/UfaW
KoUPq7zlgUwVbanHqdPw0rVozzXCOrmVoVEu84Vne2ksLB1Lbzq4oOcfixJoRl/W
fSPPrbUT5F9yec5gSXqx0CTsL32f7BDP1rTEUGdIOxP8apTP06V52xdHepKtIXjE
T9Yi6S3bj0OpHMuZQfPma+JLBNTqrr8/ARVOlaixGwoEJ0xxqVzf1Uvf4UQDGWAC
BDK6unnO5csWQkWCsQczSSik4Fi4QTAb7llAHFJxmHhGsb8PEbPNh5yIWrVH+SnF
aOn36AsXvEEu4QGECCzjsoglfu9vXqf+Bfk8BlY/n+AehVb4GtsLoYgHh+MZYaZA
qBQkiXXzvcAdrFp7SdBZ2i9iBajfxiCKEJRY3QlP/+GOFHUgCEXf5/HF5c8cwdIN
TOov0M0hZX/qF0Upi5GEkSfEKb38Y5C1gt0PoRCIld7mcPnQQDJ306d7LK7mGnJP
TYBMKWFhSepe0JIaukg8KVdH070GhUM3aFx1ZrQJ/2oLTQpuy1oZflGC1JDSUnBr
57BIK2BYtCX4W6wkz5syZHUtK1YCQmPReMI+7AvlQqPzQEICgPC5sOkWetxo+V0j
pqjKdPVw/u5Kcxy9CzpneIV9wAZpP2Sk2gqPk+7iHqwuFVztzORmjiDDlox7MZVK
eO+VUs2idtYxZJEyVGOhCLDJYm+PesRz8AI+Ly10Boh0ZMns2FEzNh/WfgkCXTVe
eCZYxyeVb8W8MQboAJgkKKeobEXVy3Mw9qxDOnWH+U9mX2hgD3RD2t4siaOtm+vi
Oes+ecWztQpfqtiyxIJlbZsDYY84XJAZVJfGU8q7i7NGJXS+F6kVhDtzt92Hma9/
Qrtvhrn8BUOjy8mR67zXpgdQjhiMwntATbN/wL6/Z1ZxLzVl03A0hUPbD0mqsM3B
bVW5eZc10DRolzT4y7Ei8PXWCB94YgAqi47i6LDG/uJi1+w5Ia4zo+wkilUh/pzy
1tzxJBgFiuGEaQo9KdccKWb8NPsSSpQ7BprVnuhTHzPfJPnEt7nQ8lAvjyZ9d6sA
boq3mwk2zJnLsJCNIhY6yJpdlehj2ri4qvOlxhx6NdLRl8eOknapTTbGYvGIY4ur
qpSqdIys1AoHX4pKqiLJqj6FSMa3wQDCpLI3f0030AVBRaorL79lsi6haN8GN0D5
rLP7WhBIAh0gB5KgB7qPY4gulI8QWt8vQdcW8YIvl3oI3dEgrVBMeBoZz6UBf0dW
9RjlEUerwmgMioqcthWRkDBswCkfTCcpy1GB4gmRQRoOMDvBER5BG+lVk39RJ+qe
4+WSnvUYdY+JHTV6i8HIf4dOngRuygGCfjeW8Eu9OugBM+8K+IDrFoVg5ZU5GFUf
R4pyXHj42Po1+fIPjOOBEQLR6/Hd53/3ja4SyEdeHl+6W5T5JfNIXghGOvMbSVDc
JqoW3aH9sl6ntwPFyiUM6z+lYUubb/OJx9iZsLR/1duFemd4lwF9DI68Atej4Tzm
3dyv1M1doXuwjK7GtZylaeeCkmp/HNIEyX6igwrj9seGC5pf7HiXfm7BGmvXHxiL
0oKxa4nAfbQ8HaNf251ZNLVTONkftylmdteG4ZEggetdpaGFxFyOIDPl01Ia9XAC
H3XsoETPAQqAL754Pe7qhJD822lLPxj2MVXz7TNha4BXAL9xXQ6VFzi89UfhNgyg
fzrHBk/QIr7M1y3friz3QpSqv5f+DHeGZmXewhGPlslRxhohpeXFcTcs8doGhXkO
3GY86Rl7T2QuT9oPUfxOFO1KoucO0zSPnqS204G4aJVK8aO34A2Y0jiKMgXEnEUO
wio3bijuYQq78EpLab+7bxAqpTXyPyYYHxLh6rXRXvEXokJW4Fo+tR5Az3vbX2Wd
INduH+9+pQgGV1KI4NPNIpvGypsmwJZbTO/BERMW5rYkW1lLfrufDIYgOC3B3oWX
zjEyy4Bq/94NUIMFvYC2SrslvR8b3JA/T1lmryUzEwNR10c/va0XxtEjXJKh4pAa
Zh7EpjaOvpoO7xDcj161FYZc4XEHZlRNGLTrGJ6USqPpOtH3rPYl2NE4Gk2uYSXM
aTpYg659RgiSOEnCPpW335N1fyscAwgKetBVETp8fE8qaakf5Ol2VeZe6SWlPxk0
i5ded4EPpasrW7IDGOQuSnkVx0VHVQKW+hfIH4qIEoCDfx+U3kvBBCZappKx9kSh
HWwFtPJNBMhP4cnqTCdFjo+QWCMjYkKrf2AxA16N0ee4K3Do47krOVXxBAyfocYU
dhorX3S9nrw/Fq8FyL19NRkvM155SUdMXxfa/SPuduSr741ffBiQW7yAWxN3Ni98
OuVn7EDBiSg/6Sf59IVgj46p439Mn8Z9HGnfV/OXJQ/XWeCobASGLbcGLfM7n5s0
aYlb/uZjX2+ktA5ybGqLzttySBwUTGqzn5m4Cg9PD2ccX2nN2v+lIFT/iOnVrisF
ABqBd6RRNDf+Y+eTL9X55suomFhiP/852tZLTQJTzMDl0/yCAxekiRJqTkKIqa+J
elL9G1r0IM2/zfT6rNCrYS6hHF7y49G9gdUK/oAkl1htpmigl5D5iTU757MK9ixm
r5n6a3uCvXhzWXI+RQecOCMLIWzDMyodvfu1oUA7ynshJoZS+76OTXSSMk0XmNAS
+1Y59FwSV/Mzwj2X/RiqQaV2cwi8omFcVXUyRvSEhpJZGQCGlhoZq6MMJmBQA9hc
CgCgVW7xd1Skz3eyKfH4FWNx8Zxm55sHEvX6hza9n87RqHAJd+pekr3rsSE388BY
5ggzoaoPsVrNTiRFrAOAGwKKfWKxkghJqygho+T3RcaIzDvB8hifAu7ZnoYK+K5b
i5jsVmy5sG2lvBC/jL7cIsUDMJ3MRTEvTOXwtM9/nU2ZdAjt6lEMtOcYRgGL3uxk
agh/EEqSEOZhU+RCuAE/1XYFD3eM8e7CPA2R9v1s20B611qrT8U7fbWLmH0vfvsc
UR4S/i+3UbJ+3qEWoyupsAT3uTYmNr/4tnX/a4WO6OGvGfNXfGxDOdOMV7pOiGs8
kNJANNr/5ifAMcW6zPuxg0lXZpcLmLdPgmO5fzdZfCHv4v6vFBev6lWpKRQxfphd
IREjQ7DNN7V1V3+3gAGApXR04mVBjvgc8C4nv7P6IHRpLv1U8400V5H/a3D2tdJJ
oypP0/XKT+y3kS3LRnQX1MOxije0T7cRhaRgzgNS3iYBBDihYyWFzpTe3vu2YrAe
inMVLj4/fdLSu4SPd/b0JJnwZkXJ01vgDpLGC7uCCoc5vYCD9KsYdM6aAUAvvLHv
Sv59vr4Sd753lglZ6ApBbJbO4CMextbhIvBEZ+vEmKlEunyHQ8vj5OzERHGDB4u4
Zq1omr1Nt/QTT1yiSyQkrnwzsETVSanLXVr2c3L4o3MtYzGt5YHOeN2jZuirCXcf
5zMed3MC4/67mTGQ+OpQjTw3+TLAVLfschUOCUr/yxtYMa3VvpgjkS3cDv7FVbzN
jC+aTptG5i4HAKZcQJkg/w8r/TusPBK402oX2GztqLtOdfL2adrNpUtTwbsLnFpg
g2X2yO43lQJ3g9cs9e9w4YOx6/p4jtfiSCVQbQrc94Qjd3et+PHB53ltE3MfhtEy
9i8jqsKBGKqkOEBcG/aEN+em1yfYVNqC2kZ5Yl8opDIfM5xqLWwUeNZNM6FxzoC8
GddYxQ7JK8JeVJVjYK+Xj8X99IEzIR2b9seV+1vDYu6sX7jO8egz6VIvA6wi0ER+
ARBN6GYat1Dnan1z+OzXhkTt4WMf02W+lbeFrI9BDZvoJ8Iqb/+HdnZ+P1kR7mMQ
OR7k+3wml01eRHgYUV51581+YAzEhaTV+pkh+xsQbmzL3TECp+CBR9EL0HnBDvY4
GjNl50BxJJiFBQnqnfXbsKIolnOibeI1dtRPcLCMPNtCO3OC0B6jgt8KKPs2Vwpc
3oI2UqCMiWDJQZnm02OoX6iWKSEh+6ReV6Elic4aowc0eedcBRK56qivKeOdM4pM
AotUH4PiX7TRlRw97+JKifGtyb/My052FwQIQGhB2aPkzkKo9VXUJTpeuaW2fmVy
Zl1x5SA0IW85IU1vcA0sHJBLA7M7XAEIbDm1JA8ikkZ2HqaMqYeeOK+1HTmoc7Br
XDTjm3eGoWw/u5ZwzOcA+h/Zm29bsHmE5v/CQQNksY+zT5TAn4zCvkOaEFZWSgZ1
a9FJ15+qZ8U5Pq0iZaJDJ3n+zYa3tkTXcrF3iRmeX9Ng4bO5Y67wLk8xV2x1cZ+g
LsTYrLY/fGR3DvmxuuJDV42tHSGMS0jqPBaHM3D78m3Pu+z6/GXq3J9PAEnpbGVS
3qC0bwrO0+ljL+1pTyRP11RQFD0Uoby46FnA+AflCADSin4/ABD4oR86ln4O434U
8NUIfM9+sULejiBrdW55h32VjXvxhor1yvf8s+z23r6KYPTxF0b2qTCGRv3x7A7u
qidwiy88T1OlWNDFuR5yQvJZ9n+gHMAAFgiGY/4wFSso0uTNHarMQgIfufVoqWK4
4GMX2CIogFeBLU5Y1fGHIDkqBrp4vj3ihVWMsr/oOJ9P+fyRpEBO8c7xDJhhIw4K
ljLIyZQZ5KTjpx9Qxt5k5Y6FQYeZhuU1HXpAVJX2t6AqIoGEydGDh8n+7F89jMaZ
WlW5fSvwTOi5i5MJFH0pcMceFctCc+Z5zm2DELfiPUmv87bCyjXMn4Qo2e67jUMN
5RS4Bu0mjh0+U1UyoHyg8uGM62cjWTUBJV3pxTIvni1YSYrMjfzF0hJiw0UbDZEk
B1znngXtZ+0kdeNaJqMMq+E4dYd4MicLGfbV02O1FbZXbCNNF+3HJg+qJziTD3An
dvfQwM2xFB1LgMeH5SE8IM7xMtM1+vcwqwp1aAf7frmOZPQSjayMhhBWKqiavy0t
ooDesi6y+FEOp61sKLyonG+rLPN5mEA2RlM0nS0tizi4LBg38Vyxqn9U3kiNKHcP
a/J4CyEK0F82vCULeu0QrTr+DM5ZAB1vArqPAHddN2c8xjVu6+f+Rk+39WGmaVbo
1mpTV91/MR57b1CsiER/+7patnuOK5j6pJl7ytZeh9MumX6+9Ua2ovvopNMQbTOo
fEMun/04jbcgCY9i3oigZ5gzhqn+5a/ihamCNS0IZ101S0PhPXbdESUYEaXo/FiJ
upbj18Vhj+pk9vcjaYv+CVIJlJ/MEQM6wObl6fGp86n8NIxY70Rzvk3a0BaPK6RA
yIcLtJchfTdhXI/ELick8zchUDHl73cT5j4yDssckRd+AIoyLPIa0CTQMTCSg+j4
3hcjK+9PKSOsPn+hNsQ8xMMHWb97zxFCh0QC824TAsLTmUfd8sfKGQMYalNl2z0h
5ukAXjPf0f7J9zBL4gsIUOh68/59ON0BuShvnhiSiB6cyziv41WBFW3Eyh8wlt12
09oWGUJpPaMDxEtv1pJ1AXjnPnMINq04pJfAqA7zzOc436VxYg0Lv1RjfyMsGk61
uRs0OR/CRootJariP+lv5lyh+EBo9NhEhUnOh/cM6lAtBRQFP3Wf5eUSwRZ3bj3y
seozfnO6tQPk4s8K640RcpJ2+V5vOx78uvQ2gow31ppDfwwLBW58yk85Nkir0Rtm
46MYvIH3lHA/aIdFMbg+ZxEMiXo1l4KoGUMgwlIOLx/jyfHmKnLctoATRjfGD+Zk
XrrWDErmuQsjmHVwd+Wn0H/oJA66iiqLWtrBNonSle8Sl5UUjiiOoQYIU6WZ1Ryk
7q7EgYP2yyV0aKEZGFDU19Db/JACobqjWz4Mj5pQMJDrrJrTEXn43SqTn/GSxf37
Ka9zWMZWwFzuDMi3YmLgrB3N7VjyZ9F3MaaP9XGG3iInELy2hhlR39CZbfsBoae8
NUSgCQ5nFQOkuAYhZr7iU5RXa8rGeNS/M6DBMakfsHM5Qqkl8BZXRQLL40L4bss/
O5oJUQNX+cU+xbnc1y9oljOn0iFwRa+cViJeaWOdiozAdqp7ElybVJHjgK+mWe0v
3GE1KPPYQ88yTPzrt66H0e6ekhOvcn0ZK6syldNdhK8S+JuV6Ap+wzurEwrbJsZY
fuTUaKDCK1VTK8esBDHWMR2H8xpkc5Wsys04kRCbjGT4OJAF2kGQXyHuYgNP2pzK
nx73uUbxo956oAoMrBi+xIHuKX6XdrromMapiw7A1Ps+F2zHij8gj9Vy4SUngQ9u
pOfNYV3lpEbwfw98zjc+CMhlV3hOibCTjtctMt319p6bGVY7+DVscIk2X9OA80oy
BHM89BdDW9n/DB57oQMsPbyJ0EYhVYvqTevt2W1559p8u5QDySCZsnGuX3wTMgK3
r07zZmS8EJrRv1kph1ck9nE/qyIdQLnkGHWeJccB4oJexWeRiY/DK4nsHL7V2GBP
jQHPUiBjNCeLaOCJ8roow8LigYzdOBOQbxjyjrI3TG2fEp1o/KjCltVj3/BuEdTo
AadRQwrjaejonrOag91/G7lsYdpdbJboR5MmU3u/QgY4sZf/646T+Q29JX8+HHul
5YS8hU9j8BsRzp4NhZ2B2bkSKc5wsr6214VReNpOVFlkOjSKaEDgcGNu2Oi6h7aa
iekbVb4eWs1WvFgNLAO0vAsndVmeVlchVBl5/dN62n4Lx4aD/411rl6A7Lhog6IW
QHOlG7NpPU0gZwMRuAPPn4BtpYZIQjPpLXZlt7eHjGYJ0WB1piWKguEVkkq4kgfe
y9HpHQG1/Rt7lLDdy7kk46/ovnEBFK2kcGhbou24xXKPTSsUVaNsyFqm5QO2QpzF
7bHDoPcWTum2aV0axyQqYFhQXMCaxcGqq42t1DkysIBEIXrXkQLTrhmm1HIJHJBV
BB4Fyzoj0xWByx3LkhwzlsmkNDmGAZF8BFy57rIbKjHk7+3T5WAIogjzep3bB6iZ
2b7DZlZJY5J32ZN7Ad33IUZYPk3afxwFXU1YokN+B4PXJnodoKrUPSo98gmKPwbl
y75OP5K5HaM/Z4Uzm7+QgGeJOUHxfyeTBwnrXw8F/YeFyy9ilzAkl6huZriiC8y8
nePOyvtC3CApECiq7Yh+Q2QnHTxbA08kOSnD+Q8NPgLhKcKtyh99a1A0Zbddycjd
lXYvaoGTaylrqtHN/ODY/F6OmwfNB/brfIM+5mi5l7H1n3rQgTH7RldICzubllMr
6u6w/edcs0fTmBnTdr7vONeKkHZN/DcGuLoaoDzSwDzE+Ll/nYXgrEA+bYYnXJxV
7dCEVjtKcJ388c0xiLMl+LnobPk/zCUkdwH/nsyol7Q8mAQgnwCTlUvCux+mGmso
JohbSRT0c8DjCM9QbFvC8kAJjc00NeIH3g9lyKLZ7Pux8631iBxm7QeoXJUdfHMh
fJcNaS/VfLWp9pIzhnWNvRUWJklNCZEADAX1X5gwYouTaGbdtlZZYdqVBqnrdbiL
Zyq2z4SbCWZ4nbohBansupwPqeiQeWWgjChDXDOh1CKsDtpSbx1bcfas646tNBcP
gVlKgp/2YDUYsW4etIBXpv8U54AMKI1TSlGn+ey0ZaV4DwTwWKAyCuMImrjk/iJa
9GoCO9lDD6tnejchSqbkWwOnDVFWBdsQcgXOTBGThWt6qdqNRosTkVYE8DSiFKVx
bDv32m+fJJbOQENsettgb+XuNNk8iIFfn2K9e0eHDwC+d1hG5ZgvG7ngRlmW3wuz
sWo/QBerlVHJZsX4vCq5Eu44VCsffGGaUVmelV6MiXzN7OXRrmHnJg3V+g8+n0P1
KoTJrke8dgfj6PM3a+wwQxM0u7VEHazhr1yowQ5Y9G96ZZvaELE+ZnT0W2SxZ7ks
7Ox+/yGT3htHAGe22NZIkZu0UFGeGVJlY7OEwIvR1St9YRXyQHa/P7GEWJFaCRXt
E3yCTtRPrDJjkCiOn60Q2ogIhnLxLkcw7HpHaQfxzQdlt9xsJBzGfchhhMG+c9aA
Q1puLXU2g8n++l8z5xLQMtmazqsS/+UVsF/avgnYgzb2d8BSUgxgE3gGrEQFi2/K
DcvCL1cObH4ngn22V8ynNT8V2K0rod3xMnSAjKXV+wnMlfWtWKX4Y3KMQRWwx8RD
r0GFecmRbqCP2LaA3Wgbuwd8KHqv3ps/G0TLDWMpisi2wMt9pZHdfu434s8BIkDh
4Hrb2SdHfnA+ADd4iJsMZiIJgVfO5B+EU/3Nzso0C1KKvyIoel4dsIWFWH+RGhU4
RL1gNcuo3ah4jk5Vgzv1J61v1nIv+xYrDvDrcUOIXUkJHe1GcmIpZAsPYFUvVfvX
SbDAo3sRpgdOKyetLJnejyWJAXtfr51xc94iKwQKIfDvR2Zw3ebwHAb9H3SPvetc
uYFZZagqaXBOkxSQnSWS5sjX205BLYpBfCUH87aO9f2tzc9QEQPTXWbibCrAZ+a4
/mUsRA3mhT63uJbkrUMWhwflM1IZCNqe0x9lEyaefw6VQfvSR+RchDsIaScIFiNV
8pOk7D0Im5+iWNdVDoQZBIJq67csy76vLAU2w5gcEuKAGkqKPsxTSPvD69IFkGwA
CJ4AqmfTmKmPc5KWF5AjE9toA33wmwyPdcimMT/7XWIEaJoa5hqruxIWiKv+UHil
3UldJrIRLRbdW7O7zGDI42BqEHZf0cxFK+wTWosnnOk+ayr/ixhcP/jCDaoN9bGZ
oKj0ExsTE8sV0p/Eot61CjTqyP65VLcE63S+E4LziWnbOrecARL1RemkB+yay2Cx
5p/bvbSxapAmDqCkackPjfbpUX426Rh+LL8ETIRKNfbRtIdXiV8fvCS6aFGCW3B2
WDegIJMqluEiaT9fK6owfE9rux1sAxayXuMRI092kU/tlxGtLjohKcZYbSMLYyvj
actm/EYc3WKG8tkP7P1xVzdrEM55hLKeKaxhS7ExVBR4f+T1gEmSxNTKHjYSyzao
IWepNSNbbjvtwhS+fTynGE4N4vqpIWfALIPWtszG3GzwC1qQPa/6KrDs9r9ha1cT
iCXF756Hhjl8FeqzWPAZnbuEV6Is1QxiPqheElTstSDJTJ8Cuh8FMT13OsmJbKZ8
SInuT94kuXpTbw/UN1/qzzmef8ky2TU/fHRapJ5KV+zXwJmhe5rPUHtF1L5bt9lZ
vvD74c2VRXm1H74KRaxskoDoV7L9aJYgmLfL87Ab3V+rQ0/LnCl385kOj5d4JVOc
nl+/s6S9U9j62YVPCtQnk9UcytIp3E6wJuFL2amkhxCPqjdkVGoj71ukLZh24S8f
xTLu/oMmk3RQ9F0m+IcTWnfuHTjV2tDCOpcXGbr9Ge667MvDEy8J0n33WccYUK8a
0NXNj5mQuHmNkEXZ9n3j3CdDViJnUmp0O3622lBNnh50NX/BZpglo1FY4ogDfywH
9oCgYOl5BQwjSc1E2Qee6J0Yxhfi+pD5qa+vrCv9olC4u1KjnTJTAn5kGs7OlJTK
wAEQXE0cwqWqo6vUlAeUYYenEnDUzJ0PA1SgKtLplTUrKCgbPOt0vjNNsxNL/Wgr
t9KGUjY3H13TZGhuRZ210HEGmAs02qfzav1DQ/5KH3cBkQD9a7tx+HpazP8bxtLO
KxqB3JLuF87bkm97fgYTdqyg22qqHOc1Pk+WL/bKy1hg1eKSPec8WUM7y66EtTms
CAwWK4HQS3mCzgjv7veFAj1Eq7txRAE/DeNFDMcDQy99+zJ/dwVkqB997+r8vWRQ
+KpTn7jqpK+TOLj9PHiups+sDah73V8x3075bhCdAYLTzd9pMZifEcP9GaE6ldWj
QcVNj6ql30iHPoBFIc+G1grc88URqiVfZJy9F9kC/GcPpVm7KJX4CZWzCKmGzxnP
JhbRaCD5j5eKcW3bsBm0M6OxZNkreGFBD/aOpoInzkmPOt8LuJjf6WnpMjXLE8LZ
s5MbB9+bHuMjud0I1N0uI+O0r28V4/svzNyQVJ9zFUki8jYyH7xzCv3K6/ihKIua
7dQ51yknm5kLkayat9rujMi1gd56qMAMhp1VljoiE0YuH6DK9+xIkW5lTdWKnEDk
UBGizj2EBjPlt3aBxd1Y2XT4mhJfd/ZQp7h+WkrZkJu5RgctehBGPj89KD0dmN1n
n6fKF2g87uD8XE80g+qyXSezBj8/DxCHhN/uKxioJm9ANuk/+hXi+bpMuguubTAJ
Ghul6Pbl54E5+EMmwiXPd6ZUnby4sF4ls47NFn/y4FBYA2XgTIJEV7pSLiBUVHHw
hXflazb+7GWi8/r6rKzaunK9p0qo0P2VxllyxlNwEYUC9DhwKa1fHDWEYg15Dlg9
dc0vjmbUVcmuZCC3noFZI4yIi+AiNcl2Yh7BhzEz2sf5F86Pvg589akKAH8x9z8t
B7Q8hoEx6Uizcb24HDtytu5ARiAOlECVdwpEHUL7Y0ZvI46MwO2xxbwI3IQVKQra
P8uC0A5ZW864cETFRLyFtpWgbENxWWgLne+DgFlEEEt5nvNDO4nGWPtv73pW7E2Z
/YLpOfZfX3qK179isz+9a7Ljw3200NGeVjrvwMdVwl/6hI6PIr4xXOgeKp/gXjBj
EN/t1NqQH2LYHrHCnzUlEkoYlf2F8o/4orB8hyZ4b9TV/LT/8gJX896vqYgShE8W
/m7jVZRFyxyyfwCGdZUHs0Jw5B+eev/GDca3eVeR1gMWJqTqM9liNLvIz0d9VGZ/
Xuhm2tmC17Ztv/8PPBTrOdqCpsWV/BzBoskjdjUeMk9j/sRingYT5Ow+JTipdfGU
jw+mkc6gPyE/I+OQeEdC9nPBlA7D8wpELPgCS4Az3LImWQS5ep/uOmrpkUoYXAPA
RSWgIINgp8wL/8B3fEYTEtekcXUa1Rg6sFsyYTRfC6uOq7Qaz4k6rNn/1YpwmqDL
FN+jRXpFz5CVrp+8p1bPBHjRAQXVTNuiMAnjD4yJqqQyiwYpaohoP58WYgrwjnT/
hltpKFKtkA/bEWcpaypNwNgtthMZ9CM9LtKRC3CVPFJHmaXwCipgkaBVQ0R+7K0v
RMrvjvIEAUl8ljM+5wI5cJHdmRW0hH/IjFF/gsbrYfFob2Zr76PZ7AXK0zCrzk8w
JdsFNUapgRC1invNBrZZIX0pCAhvNukdWLGrE6FB7kL56mMcHhtEH/JKKAQSszLE
N0NjxXCa6uZNHNLtsqrvk4laNjep2CdEjaRTDZIqWOzHM5+ykzH4eWJ9DXXAhVLP
Tv0PATwFyv59tk1Eqvweq2k3frDKM0PKK8jyYfHbTLIAVhkHf9g+Kvfi3j1JgY7E
5TqikA3L7+V5W3y9TYeU+xlVnJwV0/lK752OxXmYsURk0gkNnwGHeYA5mWNbFxbB
jMv5by2Z3hbLv6Jro8pqWHyqKdsDV6e3AaAa058Trky5zF6SLUvqnE6G52NOMooh
FNPB6YUToxHPcWz0R74IKuUTbqtv7whzi6muiHQtYQ0fFGQb/ypbNhG0goW70ubl
6Lyj9om+ovbmdn500zBp4AxPRWyUPO8Bb+IdV9jDeHzMWscDVRglSbibMbZpR0aZ
SAqLCYQ2C5rJS1o4Eyo1VWU/QYnRpdKP5oJFLA3StWhDS3zskDIuyQrsLG/o2iny
X6THxfwCDkyaP9rCg2SN87ag6WdG8szYihelFgZZThY4/OIbRKCMP87Jfto4xzRJ
0Cd4zuSHCfKohw53Xi56shyZ0zwDM0876USnPSL9zcG337pPsMFSg/3stCIUl1wj
ZXud0LKqvgV/KYx/UZd18/bSOYR7lfk/H4ZpiqJjP5s2/KBeqp8gt11lGjqtzBe2
C5hKawcInyJnrm64mP+f83jD7ZebvjV6hDgFNHNfd1v36EfnZQikrVQqEFVEH3a7
ObIoFK6tPvFiSPIsS86zFmTwPJaOk4WIgwNvkIrAf4luSf8rUhAt4Jj42198uOsR
pZi9/mZyerilPR1P8InDbKVHH1GBaHqx6UPUK1BvtHQO7rSWslGmJ78Klz1Y3JTH
nB6MVdXGnsNlCNxBIlGpf7gbDavsuumMJ+XJp5yH6xHC63z+SymrDPp7JtKNyXwN
Vsnz2tlQVzMpub8GicZlkode05xci4ekxGhBiRlldBt9e52JTm0ggUyIXfd2uYwd
49iNJmM4vhECKZ72qMYBfYemgSHZJZ80NMAmTU/2FrHzfKTNqJ1CGrEgsqAlcc3C
XAUEnseO9a6KKPjEAvGNXrACBNPs9rKrZnjOskMpg7nli2p8NsouHa+5xFe9cLLd
/hchYD2qERUpERes/jSFV8mxhJwahNt95ud9epPLp1IKxXqplPcR/GCUbz6r17Gg
zRWGeI61Ejdhukgfx49oVZpxaEc9DeBod+/RnCeDOv+8cZbDzN1N+3IEJPU/vAYE
F4bvw+5MULlp9htnBdjapdWkr3oUHXmpkb2O8eMcGiancjwFkSz9KwQzqe01+908
e2GYhB9OMKJZADihGXlDa/lRvdsSBme2Mlp0eA+459ZBGmh+7MrNQ7hHm8kzPqsx
8ooL+d5iNLHOfLeZUjAntg90XL88j2M++iUjXDdc2Qidvy/UpUCs1E8MYeIOqjWJ
FOiX3wlFN1zaiAPCkd2OBfsDvEIW2gORQVLyS+iy/kznI+3j090Omay0grPj1gW/
D8SGsUwv2otaXU7jQf+GKKi+nshlj1c2cSbH+06WmJBKrNc8yDVTSBhrWOSFqSpX
0Xzu0u54E67HrV1sEx8eZBQ2XShyCvyN1xIxPJjQ62xLQEJrwBsUnlUZ7yU8zvp8
nZDhvyRPhxIjwFJM0wizwLOOlc06wHiTEwl4xx+bRZIVb61x/sOexsRZywuPgsV2
p2iOjW7A1z4vauLmTAimzbCf7nytiNG5oyCWYvB0WNM7Db7xWSZm5kQZ5CEa6B3k
Hm+s1fKL+WQb/OnjO29B0NwFOpRtvRk3Sb28pePrLntQF/xTi6Rgu5FRXJBjRGZ7
tJ2mW1emcOFQwk7sXU9lNJmwtMjZ01UvX+fjiJBfLkx0DUshJJWSrwhLFr9pwNfe
N9cQINKKlNphs054KGIJY/Vl1E6VBahev9SQ47zZvaHi/VmDa7SwqD9rt2lrec8H
hdLN0dSS8Q5g+79gY/y+LC3e9E0o9rzWRQjr0Rt3Mvj8aGNxGuEO/EQXVc7+Yvt7
Ge92oYXCN++COCzRjQr1bp2Ebcqn/yyR3OliWI+BJeAKNzSYEj+dJMQjSdtlpbgg
xooofNNV1VCP+NSvDRqSsge7H7NrOZfjNfBUzJOwfYrJWZgodwFcmpn8P5Qyz1MR
iVZTxgzdoFuUnIG3Iv/u5hJRgXxW433Jyx+F4UgPmKAVex+TYsmH+/wUjKfon2xG
WxlZ4cUZe1IhGWMQDPdHNmka4e2pUCX0+lmzvan9UnoQMvcqgRz+bL5LGMUSbzio
YSBAAnbF0y4I5sXBoSOqnMIOa8BySE5mlOjhe7cn7uu4F298brp144T8MwwIBQlW
Mz0Ijqe2pYe4hE+EAW0LKWllCjqck9DL5g5pYKSVNnntSDYx4CrBZVC63cymdB64
yjWbUB+eWvjjoLk2iabIjRVNXEkEg35ubjwzDkuC9AgaBBcQRi+4qqNpz7tsVMTl
7GusbD4isV061YezkpQgF0Oenj76UUYn23GrO0QiWvcRWxaVuE7bjJxe6JE5Iy7i
W6woVrwAb8hpId1sIFUMgWb2tAJvN1F/aA+xvNRk7FqiDC5Nwcwzf6FgYvEtas6/
3UiOQTnFEOTQ8b3mcr2VpoDZlMbu5yykL0OzXYDEEqGdlhix7UoTM81p652xWvMm
OsiNTBEXA+ZcS8/9gkFrTDXSGTLwtRL7b4uLqIJw3tRmHIG8oNCrkEHrN9rfDQGJ
I38I0M4Odf6INMILuMe/AgXxzCtKDGsbhaCj1v5idAm0FUKrUFgx0GK4vxnZATBX
pmkme4qWA9tR5TjHH4PXln9cFV1Tld93sjdSOJghbtaFvhbR11wHRntSoyYMtsFE
cE0DHP2mwJViBznHuLgNtgJj76CYp61NWfvQieYoAiABMXKJP2waWDTqKc2K3jI/
i1v4XYXw82wuTCskpYEgRhfNGN6IMP7nKgaSjYqhs6Jo7IY6Rs0gjzuUFJ04Wyqy
lu4OR7li6XNtIp7ot7vz28NyWQkJHYE8N99+CJImwX08jtXEVYQqbN0C+vVyK4Pn
zqQi7ON4kvjvwQSV45HcXR0qVMHMD9gzECxUJTrc4obDL2DZz+/Yz6UJkJN8gpm2
e4Pn5sTbrqwFapfUS553t23f19JqMZuVp17uEnlvwmxY4eFLr2FeNWtpLB+sV89c
yIhTTt7DIzYPvrlaaoxTxmNpM9kyr63UPNWJP/xArF1KdJkYGbYQHkCIVGTY0ESP
PdmY+6i+PpMpXMkxZXSp7Yh2R8a+U8HDkG7DEdEHkh/BmgCXYMaITdf2nli3grvN
mxhMieYELTemdgoIo4+I97Zojsbon80JcmcS51i8s43df/mXrTmtAvuX1BZa83Ge
tThEd5ogwOuQyiwmPN6pjmDz0VCpi3uhovZK8Rn5p7kI5+ktyOSfqeYge87erawV
Q4ZRq8m/wm1YwewWVQPiaMTu2BmPZglg/Dpfy0RRRCPlytkcAsjJwnq4qr3uMCeY
ZC0EuDuKBpmlilMQa86OE9cTYS9tWhdz82SVHm0HPLIKnC1QY1guuZVx2JXl9If0
3D6eUgm9ExuVqK4tdwRra8aXRkoFzWx6/FV9oSpKtdkimRiE1hREhbip8fxU1tke
R3n/gijuFfwKp1E1QaPGS3uPAzPIlRWpKfYqkZE9aYCrLzJbRiRwdHJer/7miujD
WOzq0WqyhRGY/Bis7iVnd5fZIS6uEl+xHa8UKiA2CRG4zgjOKLoE74MeWCyknIdr
Hm/ZFrJQHbZOERNG3R6JqG7FDI7+YYiOZwOwdnQT7umXiHx3TBMMs78PzwaYE0xg
2riK4newTCqIRMo29OR2AkamLP+zvIUpV3EH1njnuKQ/+YNKjsxfnPfJ/cZm7DUW
8099sxdlMl4U6Efx2JLQmlN1jTSwGw4QFJPFhTHL6DPy5W5x9z3Gtfq35o/l0WLR
z7r3SSiNZ5zAUjOHQmQ0zqyES4nTwUl7Ibmru7T3TSTUhhBU7q0uzeYGiDq1FaGg
/4ORPr55kT06v5HzlYrKzdZT46LloGS+s4pjmng+MIz/ZUnAMQiqzAQNkOjRPXiy
K7r5KIMrMxr7+nJ61LRfbwWvvgHkAMzebYkvupQWqa0aj14BHKHm0pvrCQf4W6Iv
hK1EhpdD0pVgvPKXQ7mvJ4KkyzmRYiyZ6cHhhfpnBRWiWyC4oxOlvgpCKRYVoudb
kcqtkWs9hF4erIuNWcpgxkwIAp3L5trs9BWSFoji1+exRBL8p1Pew1qW5f0TsNRb
zkYk0mDDZ0mjJjLdxYX8UF3uFOG6jr3v9b0OM6gqC+Y5A8HMy/kGPeTioSktNXtr
1v1oyZ2XoHUlez5eMvsD1y6RCBm+j+6CezAATHz5OqnmJ5ZSTzGsnUJaEdvZQU6f
G00dVk3XDQlCwjF+3cdFXVYC0XEJgxZOyKXdKXUu0xp3FL3bKMUy7QT1eHts+Kgt
WtMfPx7c5I41+/Z/lNypPuNa+A/n7Y5tQr+/NZGkD6bK3iuXzabMOjn8MFg1TcnM
65qgE/Aw4efKVvX6LLfdpNmkOja4i97ObG5W3FzDgTUlY44LCB4k7q7bFIaCMrF6
RhISPRj9CpxO0+QSCsNCHmwunUryNyD0lxYnq8BdyGoq5HWleDxozRw92Z/kqqKA
hf9edX9/gcsmGgZhy+KI/LtfLqmEhWCqgO5PuZ0LI2oPMSkAY8Iq6xaHJr5Q+Agz
0DhpkGn02FwC20RN9uoeVar+6XwBngjBhfVVM1DDYB1ykoA1diuG5D0zJObnRFeD
o3GmH/mmqv5TRCl1vlLS/yjx0URy8tXi5Zg5GXDsSMXXPLOXwqh3TG0eV+NWw/c7
AW+91Cdr1stKSo8gdPocyO23BPpcyfiexyBwJ/LWvZmLlqYdOMt1dwuhk1RucWCa
lgEFIfbZ5KMmiOxz4p4IWbue9SV869pnuDxPneuIDSQogZVvGCcePAMAJxKZAxN+
TF7Pl+9b+SrU0q+ZDUrpqfiRfzknYjVh/DPEFz4/rVHHmz3lrIc/0eZRJlMNNEfB
g5FFB8UAqVU0f7eLwfU9A38ol7bkauF7vUkdZ4w0xgjyPzUc//OYKZ1rUHMAnKBJ
A8FduB/1/tCBxcvBav7AxRg3DwN4P/gSGfZM2CFGvMwxZdtzWyuX/WeYlaAGs63o
bP4GlzlEEY5noLdY3+UuLj4E0JWPmFzfaR38VUWdU5m2toDIko7H3Dze07YGIfJ5
jHtlWJ2gbhH3Ty3wKzx9X0hTOaom0YKJyZv2m4f5NrisjxkWzhcG1zxrWkoYobfz
Th/BcUIhBVoN3vSs/oA0FQRC+D9a27y88vs5rNUTHVtXUl6Ii3KmTNabTt6T+Hod
OmKwwMOGwVVg8FOR623OpD+Ezt2wf7TTnlndFgInNmd9Ew6EU9AOpTQq2jHVfrgV
YW9zp3L8oXcFLUqopydF4g/lOOaCCHGv2RE8O5TIqAhtytoHV3wepP9ct0FFgqsU
iW+I6PkvlcjyZmn2A9pwS4+NsBo5SVVfBnzL14jieNfY8wrrQ+Axhu5vV8DWCEYC
MR5BZEMcWcW4idgMpi1LW6kxhfFMqogfKFv188oZQk05bfIsx9rbHrIIBMrorfYS
n8n4VAGfImV3JV8fKX0aXu+sADGGt4txiRKkULBwBj9e7ENJjjwnXePiD6w/SHy4
o24adSByUCmT5TOCZA+vnQy7AhOqAzk3rPqpActMdZCA4G4eI9jF6zn6ECnYXb/j
SEta21c4Ez+cC0GRQ81NrII+KGJs2WKXTi81mC5wAubdPq6axZj3JxszWTJRuEa1
g8IBv0eM9xhuJNZMa2smIYmQBvDzzKqhGUjFa6NFETa2l7htAPh6LvScDj66qOlY
Z+oMZA8j/oHCu40yRAvjUg4wC2+PkYX5me2cLSK6uub8I9JWXbSWXxVMC6frAjCF
fO/JcMU5/gbN4vEqXjYZ7fmDxHds+TZKNJoayU/NLpmxrgxkwWIalaaSJ2mXnf//
ugwVX03Y3chdran+LjMBOHyIgnEfL1pmeeyGlfTrBW/FyqoWpRNqC1b7BGywEnfG
A3571VKpUQ5tpDoi+Kq97rFSCGqwA/Gc6x37VJMsy54wFQ2fPBs7GPg+wZTvpkrA
BJAWJZl1XTRKGjjflTO82FQMHFpM79OnYre0QdjRf7+I4S1LnW4WqBPMAw1Vubpr
KYqp58nQRvplZ+DUgslMbWGo7i9HP0da/H1l453OJdZDOJlJcyUT8+DJR1A6yN0f
ku2TFJPGnBNyuxGpzbITVYFkeZS4CX0CU1DQ14NvHPBItfCfodlEewlH9aiu9DqY
vPVKrvPryUQwRa63P1oTWTbA/GPN9mcRnL1fXv7/CISMDzIoIALbHqUzt6ws2V4W
RFVxDBD3UezS9jJIdqQom78JaLrxe2xoOdSRFLJJFbmEdSWaN35IVMt59M03JXHb
1rq2nAwBXE55y1CyhxPnp5sQ7W1FeIqOJlbZ8ty3cfxgciorSpRr7SJo1BNYbJaC
kdjtngzPeWUntv7wZph8xXwHcmLcApU/p9HGzkqU1abaDuVbdTbGo6W5Bs+vZDox
GcgrfZa7I0LitNg1Qljc1uVON7cvU4esK+whIAsG4SZE08uKtet8W1vPj6u2LHMM
BTWDxpi6uF/iAgCWtvFuKEgDBn3MbEkMDwzYgexCmhMdsV/eBrHxkM8UETyu0e/M
qHE+iYrebQ0VSOO+b4mfipq6v2XneKPoLE6hyfArLDtIVcHuLm47XcgGywTf8Wrq
5ucu14sYx3Dq46/rqYQ3K/69Iu42KwSvwBGuoUyE6xGDuPzKTV5guhP3I8GVEl++
kH1rWhh55VPYYaqoW9nfi8YzSpGBfdXgUl2DucpYb/xYjtIKrMSDHFhkdXjR0QE6
gASmKj7baNtoIkQBmsPoBxqG32mTyLVfguWzBEO9/yBvAW4F+CXWjxoW0s8SLTic
dxcRQi+uQEUGgPW1k3mYQ03Q+5bxcsomaS6mpBGPKDYsK6MAbLDnj/XcgPOn8lLD
OjCxhB/XajQ4LqUg4awFAFMAPu41Wrcl06rCnQ++j2FXVoiSlO9OuqGOfNbCmK9J
r5eQP0wUQxkHQdOMHZp84J41TQzRHtzPnVe5+fS03ASakNvvL67o23JPDent0Dha
dxAyvqRY9YU36ID5T2/eobXHv1YbJkmDOX78p4MGYpqIwgVAO0CYdZkFEch1TjOO
hc/36yVhQN9IMexdmRFpAjZDrlIFnGe+xoHzh2PurN/j/9fiZZmyFHIqtPEyaKCD
zId3TUe8qleAkggw4tg2I1kANSjMNCW5esWgkrOUz4Z/KxaZmZDuD5lX2iwRcceV
Axspo8Yuc4c5WAU1HDXSJ8qDqSUfgcihp2D2uUKf8Vyh3Icth9OfSnMbrCjZUCVv
D9ki9E1IUbaYQRomDXDlBmGGcgA9dXvtU4L5h1eMU0PxtAywsjl+FtYJMWDxA+vL
1lLX7zKOMEYCdssN2xztaJIDJhWW08ZOddp+xMcohSkoWwhV91m8o3j7kct0zklM
aO5CI9gAhWmuCXm4V5CNQvZ9vq7nRnhS7/u2XMYZAuEJfx8saaCdwOKzGd1ACUxG
vIqixyTRhYjf/OmgNTqdNGKVhJVl+iYNgvxWUntmOflxKQi0PsaoznneKP8KDqHc
vzjWhmHI1wLO0Y5OfLrAY9kF2regISJT2UuXmrewsjIVsSTVlgqHAz3oeVbrbutQ
pZg7BlMaIVnAomCbnv0TuvB0LwLEYEuzktEljnruB4ACvpCbpRnBAtbeLxatZtfH
puIQs8VVATtxMzEfmHbgvZLy+p0YGHXNri6mF6xHB7gZGBoJK4ioSd6hD8GPLt9r
a9ZEXZ73j95SpqqzqEAm0hJjX3QjIxbuZiAOZB0krCkv375ClGcPjtqrI19Cctgl
1IcwLfMngyu33gJTIX2pW3JwiiN0SAzh50AlLQa1ISOkyH7KGMe7rmxutUxH3Kr/
DFkZj9s6KqN0FGQKBbTgux+AVvAXZNsbhZX8j9aORYLzNORRVNQTkROxRS4zABzm
ioFSM2yPReDRA91GDStYIyIE7Y5OIVxsoE6eM9iyGJXkslG2o79XjYFDUpgNma2k
rFqI0B7Xv+F1udiYf2U7Ya1egGpxza25+B3A7Z9aXvU5iG6UGIQn1YxdHnrUy15M
oSik367qlaTBo3LxOhBbjk20U79dyZ3yQSfzqBjEkR/DP7jaB17HsA7BKK/wJFg9
hJvBNvAONROdkev3HcV7av2RmTIH2NDXumCqmMKQ5idSfuQgLamEgmzugoZyszeA
q+EIFU2wuJe5dx/HpvC1DzAuZ3oFSoYKWALL6lET1MlafDMv8RpW3by/iN2TP0JM
i0PBh3gSWxoJ4MRLZ/fdZTU8JDBc51zsnpB43df2OOF4znW6pHukXDniO9RPnN0Q
DKW3W56DIu0C8U43RQXCCSDwz5AvLqrFaRi+bZnGnz0wTvF1RD41clitLuAGPUSh
zOBcUccuxqz+UrJjU7vPYGiwLnm2A1eumb/2DXY12cRBPvsSNFpRqGvLm1Bielxb
8WfcixQy1f6VLjK5CtQHYI4l6XdsOauA/cNtIknZrwxi+GIwM2+FEMBW6MaCvo8h
hmmfXkrTQfpPqLTZJmC16WAmEH+QdPH1Wel/8JltaNEyN5y4ufGLAWGLaNbqqHyg
kh0x9iDofsgJi39MEGSb+e69lKFwwMmmzhstZiRN4279bQBK6hsKZjws1Jep55L7
oyZrpe2aWumXy9km2tgkBpz2KqgVymZ0nfEBCMFUr7ftVnhlm302+AEiF6Fqc7vh
w99+dy7kNWKNnPiCqn1sYt0DGDA+m8tEEeyw1ITKBgEe4+Xbor+E8UG2pI9SkKr6
BwGV0bBViEhHIMvjmpwz0J+t6epKnPJkjBWBjM4EbRDS7OObEGhGmD9loc9oUHiW
pWd0EvdEAXbEclWlJS5qLXMbQZVgMiCQE0UPBFU4fOG2ZkGRUQjlNIHiFy92keuw
FYPUTSnL2sY1y8R6PbwhBIxMW/6h7vxoIfb9KLzUK6hObaCQCD1lCzAvWiJnEA0I
D0HrmC1KlgQD1uiO9a6GHXeATqTNd2oLu/bK5oowxLNrOrJMqtsirafM3ZE9IuTZ
TIqOd/sJUe+HPF60uCfk7o1/Woci/h2hwcrB3bNtmuU4QwIeN1dZ65caYUFhBBjd
3dgW0SnePnBAxmi/bnW4yXwLr+h8692vZIcAUCOEjDeFyciBqmfPOF/yVY8iZfxW
BDKX3Iw+a01RINU5vilSJGkF8aDZ/67zV9NnQ1zOwLfaUw7HhNlCMG89UxRXOBBt
r2WyyPZPRBQRZmqvDtdegnzmaZK0WgSkDt/bkgx3nO8qKaQq2xWX5KpsuS3IVD4u
XT4eWr+mdpDtHymTC5bggG4Qh4x9bEllT53EY0xVNYsXI0TbNPVSz8wQx5KqQp2t
1Ifc7qhMwL5PC/4E3AlgKs8aTQBpu18p51+0k49wNaDLOKmfboWJ+pril44YNXa6
56zzhZmcHO4DR4M2dtSG0gOtsGBsycRZCKGwdMYXtKZ8IO2rvhenZPWCgEuLpo3V
YnrRTvzUwz+XNq/bh8x4FfuYscj4fLwlQ0V2QixX3rPqkeh+xuVjS41GdxQHiVbS
0b00mce1LPjBOdHGHrCZPuXM92JRqz/QjUPLmGC74WnTdzOOuHYmzNxD+r27MSSq
DVzsPdO8PBXUmgpodvHCDIuSyV5MVGSr2cb/MNl4kf4fJk/qTEkM8iTXcj5kUlle
hQNM0jtslaVrvIhk4rQaW2xsgg3zOqqZK1qmiFS5DPADUsTrn40GzMTdrX3GTvp8
DjG5oqLuLZM4sjvnvhfZFe4pLq2zz4cYQVpOPNp+NC9OAhWLf71tU5gYH1x8tjZj
rwxERl0XuwD7PZrYJgMdZbSsSBpGK5/XxwwARUAsa9he7XSlsxtJZps2wEHupMvv
3Nqyaera+wT2yF9Z19mMz94P0oIbyccAHGsHKBhyIo2TJO14HhFZ1EcU//46p/X8
RNdCJ0cFNvu6Xzsm/xeba/2LScDhU3ybtBJAaFW66IfmIhonSofJr6IcLlFoAgHm
1HIpOeJ8dqgWPwefpS24LjbmL49uq5N2xfO6B6tm91MNktIUzzNewGly7PC+7onH
dNM7kjWYd+5Zm01HBpvQGtA+y5XqD/EvwdlG0hZquGiLv3QzrsaxTtcGEut6h0MP
soFuQwueQJrFGMkNPmD9o8P/r+EZfO84EHQdCtdni3n+g3we9rA1J7Ol1oPfTqDg
iPUSzq+BSPh0eai+K6XsZi7kABx+02xdO//GyfxkB8WIAitUkUcWV8odWyQhn69N
79o3q6t+XB7a2Nj8PRDwbS8kJylt2u2WjAvSC8dcCSMIazV0c2Vrb8wJeIyAaxxb
IR+ZiVAZo7ISAEa9D3jH9EBcRCe8UHrFcfAN4zXUsK0zYox7AYVuiHo3RppYS1Mn
cQVDSMbXneyrMv9+1DetQUd6v/RQ2ZOg+OK+8ReeR3VY40dwInbzmHIFRiLCDZip
7X1PN8nViTng9yizR/ZowlacZHn42LWb3HDNeBzhv5CpS8mAff4+lOdVtEMu3Fl1
45rInzCHSIOkZR1qo77S6eMDW3eJXJW1gO/VA6XYa/f7NgPGO7oKyDbjOs93sOXE
X57ILgFOP7iwTOyqs6Upm596i/Ohy8wNbydPHMo5uY1zzpNLs4CMI7m8mmrFiSWM
yQ+EzhuLDpPlJb9F4oeIh+mybR6M9JjvoRgoR8J0fowjGnOX6h5/Gwi4mGNKwIQB
RjwN6b10RSIVbe/AgFKrTU885pLIempr/oMz7xr+hmW7RmQPOMjyNRzORoJP9d7D
fVv1njT8YpPtGNLBkdbjuNxGzB/vF2V7dAqQJAEauZxN43klVDUnpEAM7qwj1QkI
2vlTswpyRXPPxAcQ+rE5X6iAoyDzGduzGrC8+B237Rce9HO3nnivfNeqTgfopl2j
C2G4vS6SP/DQJrkT7AXk755+hzvHM8BlqRS6SynLvtmjdcqqmSRdFuR+W0t/JtV7
vTERiA/JtB1lXlMNQ30Y4MCnR1gUi1UHLKjmsNFWc9CIBtoFkcK7TQVsfGuPD0sr
rdHLir3ir45irAWO7Ciylm077WnhZ5enghA+5/RZVcdVY1DqONrdcJwPiBsrWQ7Z
kfvjzUbpe0iFVJov6meII4IYo6kVMWtnccjfSszd+H4gHpSKAGWlAI/N3z8S8sIU
MVB6OKwqUTyxHAdiI5GJpI5TLQlixtUS+Zdoalk610oMh2w/dsqT1OsXpV5XPo31
Q90oYBaJhSbbOwVNXqvm2fr+gqTs+Kdi7ffwMh7gnLAwQXmDTrizlqJspQbQxOSW
X1P6LoRxyM5j1BueEHH+rn7ibN3XV04un2kao9lCHDYnXzpbbDmRfxF3IXhF+7FG
OC4kujS/jwl7sihKfTYhCi39RwQOU61lNFf0naLx/YhtjijJJOg7ig/WRGg5f6Wk
MmlI9uix0WNV711aandfWmJ3YCwrONr6bay0GAeDM/W2PdPVnjUF2q3mW9XrPWpL
SxrsdFiHqCq+LqB1PCC3aywW5sszs3kN3UOd7lXp5dKQldbKS+lpuQYuPiTyc8bW
jE/eiQEEHy0Osp7BrvExHg6kML6CbnYjLkRxGgf1NFpJCOeATk89J0yrKVT9WSlv
wIDFv60n5aE/6xrVMzAcF05iZUdp9lVvFE453QX/pyZODotWTtXJdC/rzlZbCt5F
5Ha/KoW7A+oO2gtf4nAVJlXY7owupTulrnLXEujuPxvG/gMj/tRfKd+QWnYLeU7R
xCVNnQII300rsV1IwrK7nSnoSUwZ3/2WgCBeVtNvhpJ8UNVMo3pG0qluDcv91bGI
3MBuAxvSWMTWekwxBlI8+tanSM3ZtMfe6KUPfpbv39OPGRVI7y+q7FoYgvTd//H/
6eemSRZqBJHKQ9UoPnT3ed1odBFTG9qiJ8di9TLQq9IjGzSV16+4a3JnhGdvx8ZG
Y2R+XqKbTzXSW/4RrmWZhlZ0w/NvvcsGzqZ1E2RhriDD2ZwRmpwaPisfkQrMWMEy
85y2QqLpqKVl8rFBq6cH2EpMLMI6STWIfXmuJBnCnbJPXxtjan8GQHCnhTRBMaPK
AR0lLvlgnffsL7yoc4wNX75SYXz4BG/DgpjQ5lgPsgtbQNVwQMVKOGG0MRjA2m9y
Wf0fFysmHBNOJ4b86SP5m7R8WQKY2fVDO0vFdvkK1Vxc0zxlfZ8RjPBPkOtV+V2Y
a5pO7TdxGI1b+cY1mMidz5iFt5bu8F/sfhDWyc3xacM8KLQZQ/ZfXTkjXj4uokhw
eCOFqnFrAvTauVx7XIxQYC/C51DUScZEdsJDCiayOMC5uPahBvzyLLALi4Htd1hI
KSNIKe0/OG1LNynQp+krv+azSaBXWxq2PR1ayxIBr7aoRer8UfkRHlUofluKwcmR
7fyCITEUzNoh47JUFCYNTmhIKPQdf0bfLKqmDBdhwFLrMYWzxYgCv92PMl4ttJK9
UBmf4SaV7OGN06dLFIfzHjQBCnXhAU7eifAhVCtSjXT9NdVHaMicckz7pz0rW5V/
f/IosNMpmJWADnWWIPbZ+b5LFwSBnMkb6ZfYPInVxLOW2NbCAJyA+NLIGpLgMSqU
03S/9fUl911fopRz9U+XeMmAegufiCJNWjK9rYN7c1Unnecgv9Fp/WgON7i4wTPl
4bM728/SyO90PZZAirQeJ37cfB09dtpvBYipHTopSQV7SQH0BpZooawejuiLrcY5
g6CVp1IUcpeGPS7vaYnxrozc4bTcDUu5Tl5a/YYOzYsioDdWo8odC34jsSw8ULxr
AJFsbg2jXbndKCQFu4J3cYWtAt+USSVtBrjJtbVmvvPU1MALsu+NmgYFHMtXnL4F
Q0bSBTvHwEF17kb0hMHoJ4X0BBLeAQD02nj/1nwmo4wjo6JzquLDON42/fY8pwuF
cFxkX09b7LVdOcc00OcWzLcIQ1e1p3dfvPEe/MQL3d/LAfd1oSBjv9AVN7BB8D7O
ozKRfiQ/XCBe/nIZRRDB8o/zGBp4NS4pNe21iJBX8JdugRYT7Nl+V4L27KGKHnw0
nSpy81NHYuSXwjwlc5ZFjWZNi/2aT+8vryU0/+tLfjhnn5Z2kFL77B3ORQwci69X
h+Phu9lFtPxpG/498XKPPj+IL/+aJOxgCb+YgNiNjngW4MccVottcorPcB1x9meE
LTwA/ms1PN+0kpVmf2BMD5yKkY7wMD/COzj0fzpFKg2iCmhQLffGY6O8IBobj4mI
IXbZIh9UZ74p/UPsRo1EsECJ7WT9LYZOZTBWPjMHOsSQPGydjwYMeQx6A8jBBUGh
fijF7AzyquFVPNmvJfU9Z77aZT3mDOuPokFkLjJlv8lWAygm4pk6YofYDkCXqXZV
x9Uo3GmMFlriKiPd+H/gfIDW83ic+YyKD+oa+QQe1wkrSqgkf0idZ3wQ4vZA3KOL
b2Kfl6O3WkToeULzGghOQecE+qzW4unV0l2SN7amlTJRCYNshLV5lckxXOYT1ARH
2WyKuM4jHmq9S3QeVLGx4+SnZGfC91N7V4ubOyXHmaAXhn0gihhUiZ1LNhJVemCT
rmK4q/LdSShA6MWvJnzATthCk9bjoo7mUF12YGYs2T39BhHZHA+WwWTkUfNZtb0V
jfgvb9D5Ig1x9+nYgveKJtTEwz3WaBLAOSF4nIh/3o24pCHZ1nNPEbWBDLPBmjkm
KwuwTUyDK28vk6iSeF3p5rsf6Q/J9NWV4yg2p8cDCbVqZRlXK91zU5T+/AgIupdr
ZesUEEfJYPscH37Zqw6Y9uJl5lrsozD7Naj6Z3xFYwsnSBmlL80Q4n29yOCE7jCX
2r6uRh4R59ZT6bwIk94OArCZ7mXLmHnq/MQIi1d2VKUYYeMaQ7//memiTMeDEc7S
ha614KHjG7B3ySeeuHUXNm+Rl0+kd3brAAQCBT7OrkgorFgb95ytLIpGG0u7sKng
zG4xge68gP+ubE3ZuFiEqqxnAz/sP1mFxDrfhmLWKMLjpvDRDc6M4KxjOlEZFFZ/
MhQDzsPWOFz6bAbCXhZSHmc2hS5d+Ey48TL27enkTXVXYPozGIWQivXOIEIxQwAx
7eDUw3SJhEmjyPoNHrP9OIuQatGrnpNSlEO99XOgv0dZA47yJL6W7T+3bm2hzWRM
x7gEzQ8gkRxQk+kuviyfrK6qyUK1nT3EYGHBe9KGQccIvuaNnmO+4YCXiJ72aaeR
40Ap3mKzT7A9rK6Rm5HjucBw3O3xXtiBEDpfcTPERjIaZMtz91krubLDlMPrWnEh
FvpUfHao45tYtKmJF7DQGCKBpyRm3MRutPwETVkhX+pu7QwBFNOjXAvmHrnh76IU
gg5bMeROqiToPKuwx6s9Fq9L9cVOaaiz/8T81tz8rOZKMZ2jN36tBh5K17jH9NhG
NtJaTfks8RDz3xNzYGjOe3MXgRdCwRfUazMjwJyF3mwOhtUUT/gE+OXqW7DU/Fqu
v0ntnpg0t7CRmrPKF2P1bO41ePkwy+PTi6NiJ0IwM44F6W5bzgLsg42S1+pXncui
yNlbHjHe8QFnbcEm+iMmvB8/DX+KS+GRXuRptZmAgUpgmFMB/koK8iLBcOHki8is
mic82fKPd7qAud3C5cEPhA/zG83mC0SOiE2LfGE15eMDeo1OauN5+z9gUQ37Ct5d
7uZLByHTiOvDANZYDGvRGNrwTQGJizkv9dE5VxNpD1i+tSy1+oY/77BwfI/HguXt
AV9+FHgnsE/QwmLwgfCPO1CQI3S7xrdSfSPYBgwrC/I+m7M5sFsVMo/zR6UHPe5U
QfdYnGQbXJdcwKk04rqU+2YsyLPofSt5WU/mt3Ftn9U7dqlvESFXK73RucAt1sjH
tc2VzAhxfvqmBQufCDA5yYgOYEipV9DtOWKl9g+8Hx57Uecs8Lhkz3z6QYasEyf8
StfawE53XPXShHL2OZG+7W9hGibjONMAYEzIwYwoC8OLXPe2NNRIXZssVQlUFEaM
Kxv0aB16ALXiKmNfTvn0bAV81+u6rXd4QKK02bsoiTTdgW6MTsDI2ErVMGCjhK6y
lNw8vrFXN6aOV5zDH4gwOMguQdm+rmUGc9cEnDIbhCL2fiKYCfQS7fM7B2IZU9yh
aQBoj1SYuLIvo19Tt7OCMZDhBEL2R0hAwCFhtHXmV7dlsALoi1/lHqyoS//DwYEM
RhT3PfNlVk/tiUJvVVFn9EQ09+3qeAdC+Nh9hs4NlMEfu+fo0X9NMtx1tSHP44eM
nX9iV3YwXPYoy9BBKRVQ0RCtUpuS6ewIFm8+2gfFaUCqsb8zfxQdLhtsFprpKBP6
ro4kWH4ABTm1oatXMzg/kRMWd+UZlFCbhn4tU2C20E6+4WdG7bm8a/vBCRVYrXMw
lHwRyUY0KYSjbJ6KJ2GkKuwYz3Oe5uzOmoLqy7u9hImAGwXkE+i3UISj8Z395XvV
9321wJoPk3hC3gy3fGTGmepthphuXD6iXk9BFI0UNjd5FrRhyb08CDOamMkiDNhz
ZB3jwoEL3tSLu9N+9noai5kpIQmbKhwKVMJkp80RlgSXQ1Gj4y8Vkq3vn4XY73Ay
GjQ/iLDMFs8GzMabSRz6vk6B69wvUFxCpq2p0EnUERhuOBP1SyXxdhhdSkL8/nT3
Jsbd/55IU1N0aWVEGjmkqqK02+xYkR/iEGUCtAPHGvHhU/TnKfgPa8VF0T6+BuRX
iRo2NBu4U3Ys0ishGSExdkIWMnUla7crza6TstY1ZrlyZVb58C2+DOCz3zhmW+TH
iyh8+jnT+eCQq2jk+COdsGSW/0aO1IzIIpQh/GYUurozgWXREiGOUaR2Y4cD1GXJ
YooWrikalMdY+gpKKtRrtHK2TJhZaZEetzqdJHk8UhnLfVegVmWKeCSlrbc7DxiK
TDY76KUp4+4T/c+Gopek+cNxsV6wywF08BNbUEwtvTggMAvd6oyHyCYVxqwpQ+bP
S556wCQgZhAeTDkNq4IBGY9bGgqlFIE3/7viGJmnFX+etw+eOIMKxVhGrfyOEv1g
5bbjoh4g3Yc1mUADmLoK1QqNn5UBFtt1xfesTW/iOlDFN+UK9SvllWA0nCn15Z/x
6HE5RTtuaiOtc2M8M9elAauPxsL4RjLTqbJqlCLJtHCAlow20yRitIYY3AAreHnh
f/jYsmmlEBDAXFt70zgNP4MBip3eR68aS0NFrqmGJQ+7tFLmQ5AycK5nOxVCGfmY
Hhw6AQaQoSP7SrVqG5ugYSWBjVfg8khTd/Hjfi845Q/4QKokWBkI8yKRMZ4LHboS
x4g/gZUUivZJOlRYbpyvx+sUDn1xOUOZn5Ik+PUnMZ6K49D9h5Su4Zk24/VHx9Rd
rjhQN2WWSOG7oJOrL2FnUpU6abcAluRtaRoEKCMSYKSa58WdifhmhcjIoX8ZEugE
6odqd0VvLWTAxj6/Bb676a4/1+nVqutpdRlM+nld0Eab6ppKneuwhF++d5FigFXJ
qTd6cxiM278+vh/7jPZ0fG57GbJMlP4V2kgu0V+vvMpIlDIN4xzDynES4Bdbr6bj
v+GsODlh82Nah5UAtZ33eDzKUv5eel8IA0el0lXKPZ/yb1o2aIso0bgleYhA9rcT
pXHIRBYSTqIhYJumzZgim2Z1O14RqITPMzmm3GhqEXwlNyLpecX9vbQPr7Gfvr7I
TYUhx0km8UtTlnc1D0uVUXqzXsE465PnYB+aK5RiXxmSePEjm5nP1m91QA/atuyt
mllFpbS2SB7sQl2OnkEO6LukiPKEJdpPITwnOYaYBwpMycoF3sJ8IrX2Bix/IfoN
5tFj7QfhfIu5Yo1S7j5y5PI3oFnikY0lW1JvqWFYDpqSDZ/4bQ3dJULqDys06uH2
SbhJhHz0ZtcP26BEXIDwXkJYzMvCW70xbTuAk6myOxU+9w0AO7TaQdW/p21XE7fL
YsypDtZhZg+oixycJn3H7DaIDaNCP98E4O3VIxHFEC97W07cGnuD2lJ7aLD6pZPC
zh3bNOhHXjBbBE9jQcANWgr+RcgCErLpwoYZKrcosgkjbooHvFK75fifaVj/AqeI
eCDcmxHSHOcOOM7BBBfwuaewBBsPRqmK+wLAz6cHct1yqGMotkHFRg3wPcKQaNuP
5wk98/FH5X76Q/kxpzTr62Bnlj0KhPFC1OXDAof+rUW7hBrJPa4wdZz5l1vfyVin
8kwmURTRR3tQVQlX2wqIoPL9iOgP5UseMZbrxOfC5guAfRaGdxex2e+ywveJFbFl
HDwyezwwfNz2iu8mhj0XRgHIyDvgToDYnwhiwCc3neiyR2p8KlWaI/L/LOzBfpC5
iiFAssNniwXBiXtgO2lqjsibb5hVQHol4lEd5F31d7DiyYp7krDPy+DOyNeIC807
ut9FaNYedrdcedU1aiYX4It6wayylSl3B9j/Y5nBVCnbe8WgrIHI9uCAHWZ4Ykmt
Yo/EOvj8GvtSRU95o41IQJ8y+ve0sc+kKL50V2mANHeJ7SdI+BdCSV0llZ/eLtTh
8WGwsIOoGLj5n3aDrCsiDNd/hIw901gMDlnao0TipxjeGADidwYVuG3q6ql/D6CQ
n2okimxQTvQFReyG5U2JqFhp8Lh+xBR5uZBlQLzBkSdFnFn048Yg5/fvAjOPfMa9
YY0JLCZq5lWAEMiOZBezfox83baiKHZF+FRmxysD+sdh449NdXxEq91R5R4VBfTT
CX70STZF+6f3o+WNaZxI31NgA0Z0Z3WR6G88m06UZ4aqnu6qc0+xNOOpRtc3DC8Z
37fkIpKLm0vozj1cjF6SCQCwaxpRM5GD7LRuu9bV9hLeH1qg8odFCpf+5g1lEz4D
aNngcg+RKW+5xtsMlhgP4ZxtP3DKknHB41LvrzBdRbL0L1GyxZFp+IvJHXf5Xao5
L3bzpps2aOgHWTZrcRPc9nWlqns59UDG/vlfRRLpV1NQ3MDcHPrA1YL2EgQbguKK
lD4WW0k98GY/SLH9lCsUXuORYJqLgRfTZcbHZVi1vdws5oGJCt4X+rmIqzdjQRpr
RrnqZjMiyTXK99XB9pyKa+K6nyH4HBFgkEUfnpHedver1LX4rLNAqO6r4UDvPmPI
80fp3vV9v6Tq3jK58ivMtxwpNu3qB+MhW/w5IUZsw2d1P1aXpPPrM2ITVxMqe9Ts
DIqDnoLFKcnWvhRYjVCTFdvTdzk2p8HeMQSicoLVfcObyDRV0yPPd+8hQ3G7WFMl
OdO2MB7/H07S3BsslGdIduCPQoEWKmKEwAtbLJtuFKza67w9Exe/F5ouGMu5gb+c
hu5AXmCAQc0VFTUo1S5wPGkR6AUt3l/rppvyzMocN2RrLCCjP59DGJaEYMh8QaC3
W0yLi/F0UD6qiY8eYJefZdj2fJQfuG/gJtYHUIqD5kdTt2ei7o3/yoCnnC+XqFh1
Wzk3jwJqARWHj/UYitzjlLzUrDu0MjrZWz58bsrO/YSQugAu2R4blNDWZczhkW81
IpL+8tgEGar9Pv9EDyYXdzCXs5QuJBTVStAGY54IYsxbhFlbOxNN8Bom2ygUGSHj
vZEV9BAmnzfjRyA0ox7EyVo9Ho0rLmKzT0bgi3fq5YHAdgDA6qC/AymYDrnblIle
f8QhfyoI3a6v9xOH80ZAIrMOIOvDrmKF1CSmAzcuuV+7rSm6i+Z0LDT9yzm76h93
nE4ET8i9cSRRMMKwIzPdmxlayKtpRaQDZy6ZBcWifx/Htieg4LTtXv/ScW6zxnci
LyjRmV+Fmk9HTnZYr8LGcqsJFGpGs2M9pWEImkPnNR7uBO3f9GNf+UxD14TCB8vb
mmIyQeF8ZTgGzbeoiRPmPlQ4KtIu9KIklXbdiH+71lSpgoLyOYze+W4OIUaFKPkD
NEXwWhU2Z78CdZqJyQpsFPSvh/jXzN4xzO6eJYiQurJnUUmIDM9OTq8+1BO1Tf2M
DzNf85g5hwy2t7ia9F7U8ANjNRROjYR/LkXXHFjJHCeCo62MCApljZVZLL2YnGE/
4m1h7el3fPUMtKdTRCRm6KVs0NOS2uCtj8dDjjT8D+/qq5ufX9UFrwT5i+bV5etw
9SLOguL3b9xJM+0yotk81s3Pp7FGdA+Diuo9Svd4DtRPIAvWOo+LzH6Un5qiokdt
U0Y5zHKlcZN6XNk/016lKJUbjQ8NqjVUFLZOtxNFeE0CHB7bSDGWQLhqiUD/AHzR
U2Y8oetR1slOnCfNW9T0gO6gGJ1o9heZbf9lCcYz0OxlvsuBJEZu5LWwo8LeCSVE
W1hpb7Yw3rPSgEyTR+2PathCpLqTN5dyfpbFbsDJE0lheKFF9z93RejUZVqDZBrO
0XMoIBAVPUXkwRyBsMV0FbSRO8MmzdU6wk9aDKY0IxPUJ561oQXDVLSgOtB7SIET
7Gy6ptKcd5Hq9qagNkY+eTrGEct8J4Wt/m6dQK4HIlIBg3N6ktd7fCwK12cG7qzo
7e3Jiz7Fe/MAQB3kH4n8aGDvmFcorpg8yhOQSqQp/0wPFAKtb2xPGx1STCCtVOYo
K4NoCKF37zhUfSftGG8hxLsqfZgtiG3JyyW90hUpEm0KAnwcVNTjK2uymuCrUtDv
FllmuOI+tVLtYn4wdo+GJCZ4RLqspqY2BVSG4MMQBmPlU7OiQsTTLjfNfHQQi/0f
V6kO3m51j4RtCCzwr+9UkarRyuQ2GIKYMbnZ9Ap5pe6m9YblDN+bnl3J6RT3//l+
VfXcLiex6lVBmsWt3VzTTwGS1wGm8GxYqJo6G88tG8+3h+EmZ52TvKvX0CQPWWdD
MHzYnSn/WnxGKEW16R/TmEG7FgYXW0oP6U1f1+yx0rlbgtdgQJC7Anxt5nYP/fes
cv2i8fOI2RyAX55ig5tYLamiqQ3sp5fj8gH5qihEapccpVxLgKPVdu3kwsuSjOPV
fFZHyRC7OffdcvGAf2DJ6bKnxJ2Qy+xsn0q5Dw0Br4ChZzM+b3ebklfEenXhra/b
mGzq4f4r06vPyIuxioA7zRyBqrNCjfKUlaLxG6c/B2MLThOh3IwM8XQsVP7rN1ja
EHROIW2aiVjbvy4qsa18WqIBpBydvF62dN6VUiyqBLZMHLfA7+BL3TZUOAed/dxh
fSuGsT1yYtN6UiyjnDoqdJ7QhR67xC8KnRWM4K/G6Qm8uWLT9US4vqTIcN86bTy4
n2Au2OCurtFmdRGlGQH6MGohLaRMeRlOOnegd5GaIWEqkcUAhesFhRieUMPCWixB
yLZrb2Ds3/N7gDfIynypnIyzkE65nYaE0Ax+SVJn1FJZ3I3gkNOzM47v/QX6x3bd
TnGmmCtQOZ9uwXR8fTdW7ZbE0aifzAmXr8x7RWPJCZ9lQxZPojjJLoK3xyAHqz8F
KIRNXz03Bi+PtBTQ53J3dfdJYNKr8o8eJEA8UPjmWcP5rXQXnucYeRriCRwNu/J+
nQ155kkytX9m9+ECLBPh8ndYz2lbjQMoxXIw5oRk/A6HH958QFbELsrTYucEoxMj
dM1K5zzogGHJMexkPTX9xViSQPAPjRDDXpYmGTtzjv+r34ftJ0MFuf4ypY00gU7Q
xIuWe8UWc4TS+uYQ5SBffA0TP2c0Sf5xL12fxrS6WbD8mt2RFvmap7/BhCzIVBur
tT4zqbeXnH0lEgMmztuqHXHcYGpHJjf1lCbYzYCgj9mlLs2Fi+5mkyWPgR/KwJLw
fi+P3Snm2OlG3VO67e6lmF1a/avbqy8zi7R5XtY+dHxxuITozoQ8HkQCkWZU3eB0
zhSbVo+k0iOUKeW5grQuWlcLQ2HnP5mm0O/IKZfgFyguBAgXHtAyQpRodu+RLvRQ
f/CsQifbRC3DpbbrPHEsfH1qxX3psSc1xc1hIPiBOLLd9Zfpg7sdSbQF6UG5rXyf
7mU9OcQlM3c8hO0IFcXYO63u3SsFEJfjSVpHk9gG0u0YNQAucpmal6DE0mNaYc+x
4rE55u8eV6nN/acLZ1xiX9+PgSWySWnb53e/LARL8llPMVnRDl3UNegGSKEE2f93
Qrjnl0LL4wXMZx9d8KZOBkMvzo9rYgFQdxtDARxDnHtbkY/bwK2PG6aeMQ6XMr/q
L2+l8cmNpH/rh6I2JXRi34qOxVmwEZ7jJdUXWIFzGkvq4ll5jVE0JAwaiwkbXbBL
lagQJCAj/QFC/ECMdUf+/Sszc2TG2MXSw5gPk+7+HYxMtW97MRiPV6UQ8xXqd9vv
oma2BWjm7MeXVmG+3bT//giyiI4STWCGxlGIY+N7lUEjLqxym9rIFCvM8s12ha1A
58x1eg5uFa2xsgAkGuXoyU5NlG07HLMlDNr1QpYxA5AAMxoH/vz0HFago4zef+PJ
9yzjHEomhPj6cYoijnjKi/7h5Iq3Sl1PQwmnnWbW/Qik1FGQW7m5B4DoCXZAYpC7
aANRNxCsHoKPdGgx/Lwo8ANT+PdIVmH/TcDXgnmRZi6QJc3edjSeGlHeCtkpBj7w
IgGpoGrrUUbXXL9wr88rJ2YaOYLepY7kM2/mFK0CJZano6as4jABUJaML66V5x/9
8HIpao3y8aUxyQrOKjomySapVDrNhLs7PrYwrcYRUn/NPIJVBaw+eoE9Bgr6D2g2
0v9c0ANgwyP+6XL/7oDyyrTm2kOkeLYEzdyC8teBh0lSBrEYNwSgro2u3OMWqAkz
dJYx+miUGSG1xC0dJf8uub2ndd4DJj6rBRqeN9VwH3ZHc0+YhPc9AbFd40TcvcDc
8WINr7sO7Yn1xQgDVNZan0oE3y9vB/7oRmJ7EMrqq/LAU0aIu1s7y+OBh122Ud5y
Gw3wg/YnJq5rS9paT/toR3BIxmOb7uacmVAQdjkg2UDYEiA2PTpUkhh/HawZvyq9
OuA0QRNcCfy+jJlGN3zIMBJahaCwJ3bqy7lY0SSVIMfIBzf7hmrc4g1KHCDroM5R
uNiMcqBWDO7mEUgBMK2FgJqQrthbAVLmMvV/zT69EFiXwALo+gGcWZLd/SMMXtSv
IzrivkwIbe4xxsDityuJjaZRY4u5ez+4anl4E0xvChMNQIArgkm1k6R+5yJ+6hD5
+rOfek4ke7zlnR/CqiHJOVIYN9k92G9xe+7YOwMGppvuKlYVCdOKzBZDwHsK0GfV
ENZ0DvP224nXu3ZomnEwU0mE3NsKZGp9lDJtGq702RDPXFje/oIs+9KwaBW0VC0P
WOuxiGrZiuRPamvZ40EjpLJJpc9S3YocXno8v0WqkUDjPRy7qNJcYKjFDDiDY3mM
lCH/qzNfi1p3br2lJIgiHb5C8sXuHinSztjzkUYnm3m00OwRo+l9px8g2QyRtBQ0
WlIS+q7vmmhG8yh2i7bnbYM9Oq36o0ZpSmt7iSepAHW9yWnFMhy0kdDxK5ifl5G/
VaKWSQhRmCtrVowB2OmiAC+PU6hOMslmyBS4VP4wTG4H6+1RX2JulATWbdn2ZdzE
X3533hjVr/61o5CReJM4tKfiQvBdMgNk2X8nPkmh06XkHq7qiqRVbQ9gvDwMtGDb
TS+iQv8fXyN+A6Gpxww3+pRSgSwnmqyagsw33TDokJXEdwlM3CPf5o6w5CH1RNWX
WmOcfY2hnHLSEL9QM51cClYZY5a2CJqWHsBpzbJxzcX7LWEd3vn+ICd1s2X7kq6g
i33sme9v0+mEFlsSJXcwh+DRlIAtRulr9m2OjrNUXNl6BA1TZ0ZSm7d6BgoeFWTw
Y1avwGYeRuJWv69HfReSzPW+XvCnOsxFsiL/rV1t7W7SbXKIUBklBZIxneNRFzo8
VVNCZW4K0PmX9h2WG9pHfsrFJhV6P6b+N5q0gS4EEkSQk82UTX8P+ZyiIY6eiLAU
kxs/Yt3dajt3PNT4kkvuakpSYf2RaftF35+VWhG2cBCoQ5DLOrSPouatf+YU4cBw
2JP5Vr4o4aYLMb3txxxfK87W7t+BoLv0dKvg4cwpc/1IFHq2plLSGstbf10jmlpO
sht7KQmhE/go5ef++MS9uQYhxew4TaGCEPuSTSZPLREwRcsUi5PEsAzqt3vyc6df
p4oSa20KNIpI5WTHm0B07kWyXxMUacgSfFYFjoTlPUSuPlQJm6+NeLvUp/Llbxf1
ToE/q39maijEk59IgvDQLg7KVjkLcQsSUeaT7IaeynM7qrsYIRRmY9lvZpB2bsaJ
X/hgSv6M+uL10uGvE7E9Txxe05+4ouReTsF+JW5lmOkea+pCBavj330mxfBe7AP3
/D1TKELf0y6qU4qyYLZ/Pswgbda3qLLoJA3sztIB212Cyd5gCsPxQ9k/15UsBZCl
xEroWvTxIFd46axyC7clpFjtDI8y/QO9bfFGQZHIsSEAZIpBqFDc9jaW/YwH16CY
rwT1nqOkN1F9aWF6cRY98pKt9SbV/yIP7wxLASUJVkM0YsfX0zHCRDi56FcHJ8F7
6c2BFcdBtyg89dmC6LBeHkbcNBTkk3zvvyQzpSrJxYBZ+BHjPc4NMGcHT2hLCtuB
qtcIOFYCo0vUbCccyrG5AEcTWMKKQaPkq/6KOZFIs5PuXHgUYXHKCl51L+PJZzW4
XUTV0TihGAZ/ajUXxKI6D+EEAqks+rXcXDBLd1b5LrHdVEPV0e23wkyetplMmFBV
hayeY+uMgxr81Tc2Obzsh6LkOrH8jTyJsDP8i/HXTRnyEs2609MTQ122A6i4ZLr8
R0LAKYxmluwvfkZ1WieeXGqO83NrBaeEYBSSmA8JEdNHWzjKSQ1Mjp+Y8DwkGiSX
QlIiq4s1V3v3BYyHls6J7RaDigWar4W6h7jcpDOJOYhYgm1fPbH+ig3uCe7QN7GW
2FkfLeCBjAPO2SEd3R7cDOiqBNTmmEDFE13P4DeWFSRmywwb6gOrQsCE/cilyDQy
8ZOzMp/USjGidZvUl/eDw6IjVM1V+DStL6Itv+dxAaev4tf/rc0A864EcHXCiKSH
T2KPT2I7JLihAcfY2kjmhkgWKLwFL77OhyGLhlg53Zq2Pta1Z64TIoEWhpLu56yw
OMZICRgc5vCgUWA4snMgf1blaC28lcaNoVmhs+xlcpKoOyuitNqzV08g4lXdejVd
RJDGEzpT2RhMdTpn9AAyR4Z1Bnac3LAI5yFc0g5OD9dfdmg8RNMU/+nkaRC5l7Pb
muHm2BxTrWTcywP20tefXysBM3o5rENsztIYAmLEjKJXfF2FfusBUloXnTExOY12
zb/bVXvJYo0YBtn70qr7AnY21RCk4yUFtcsWqpq+6SthJtM5oiqlIcaLy5Qb3uBa
DEww9CwKZ/1zbyXWBaQfOT4RebCe97NN9qH+TMFm2p04cBTfsuHOG6nm71s9413Q
2Pj5sIEQdXJkJCS0GJZHxnfDz/TXvCdK9ux26EGmiZrQDwkKTkBxFV9zmcY91n1W
UM+srj46N1xkaW5phW6cqso2aXf1a+bx1IyLuyk7W+G+G80HODl9L5eF92MqEPMH
pxTx/QIVup0H51i+2lA4NdRNfyr6Vrt0TUILosqqABm/91BKdZso0EJno0ZYtN4X
ZTcf+QyHVnTxN94gb/2bzRmsJd8WeJDALRGyGz7rPp2RlYXkrmuyLvrjrIj3jbs4
7saJPm2e/FwzFb8xRTIhGt85n2NhE+3dtLLtARntlRtKVBRX2vcW6OyKwhZYlgKg
JEPdg/fjGFRHCGB5MH83R+ixFe2mwZlSGofncWLOBWqoQCrVO2wabRyRwZOiSWfM
wnnaxnawsh01xMSUn66HnM7VtMX660UJhxdtihPLHfXZTuNw1C01oQOULOz/f8Xq
uoi1bYHbjuhAqgFFsWjmv20/YF+inlA+si1NZKqkEDsj+JwCP0c0WH4yiKV8g+YO
OZeh+He6n9RACswoPkyOcdf/gYL5YPI2Nc6KvmBoVlKtIa9kCS8XtNhvtC31QaA6
bjy1woQygbJN9MknPkFQHcheChizQCshwEhkd9EqMyugDYk1Dlfl3fLBGF2SITQk
gO4KsB7eYU33oDnHNnouvQ/eHHIduyzdg3aszjm9VKND3DC3F2qfZ2aO5D3P3wt8
iiALpwOYtje9kJNv4z/Nesmq7I3EUsLheh/dZ/HH4i+t2AYc52NyUkUMXvpfchMO
xljQZYuBZVL0L7HPUcmZUwwrEHyhSAnBssJPcRdp3Q8Wirb0b9aEekTCRBuzr7b0
E6+3A/4DrI/CW4mgP7jWVvwX5Gtf67VBsArgXEBOJN+zFmRCTQqb6X3Z4MyLUamK
pJMpfJNSx43JM6pJfeiP2XQwCI5XHz2JQozKbzlOqRZdFx8YIeR/cOHNgJaX9DD8
+EsGSsL5GwQj+TKitAttJVmUCVTSz3WZsKBOIirK2DsBTzaiSDpOCIIOkYJuqtaz
Plzky6sD2yAXCqvn7fIoEzayBEaxPnynGSWyGSypT8ajdenh6W6VUpboURiRDJBY
Wo/zPSO63BAEonv/maRcTwdFotNnUihesvcpZWepDbXYEvpiNxhopudtrNUuzwWN
gB/WpvgEH6LYbXcii4yaXzaCYLo8xHeM6oYuMqViWQi7tMYlSdsEAv1rzVdOkr8d
e6wirTqtU8DBOuZZ9Ha6fmw4PWroVrx65Y+YkcGKl+vfv7eWyHReC2qxePC2y+3u
kl3+RMXrE6731uppcIkylLiWzCuKVnUwOu5twgDmPT8Ig6gK08gvrmlj57jMSLpP
iWTUZi2iARIp0Fp7qb/TqPBM5ZLHu2GQ4vKBn6HQdZ4ui51I5MydYemNnAEzSD2e
Xb7te3G518+Spt10sxlYBTMyxGZ63m9MULLz5wOCgcDeFVJxFO4LFZTtTBsqSZHi
jWs7bqhuKJ83XjUYIiltk5UDJhlKFGuyEMXGwcq3GLbGD7IZIjBrnVwa/AGIblka
Gn37WIZow5dg3ah23Lw3QhDajgAmFLEfN5CgjIquc+fI1uxm7Lvp5gdGhGy0ETie
HSsLP4TjARyYBoEKap3c7vLi31i7RcbItr6kZ0jLjoXWezldxDX5IxjGhFoiOA95
BrRPd9CYCakgWhT0a/e3s0/R5i/QJ1Dspq55g90GkuBuwziOzwxfTT0AAvH1ReAy
JhY7IfaMIVCkjzkjIXqjpXpuUn6csimMYIZllliCb2jsv5oF76Awsze7/s/ab08z
XzWetGbDqV/E6avcouhsIN2uE7h0jT3rfM+btwuWm2IQyiHdvRYCThjX38oANKvY
a+pdx/fmeSG+4kCOs7ztfk0dtgxTuv2O6+3U1OwBaejc5T9BrZy6/vVmig7kHtGQ
Od3cghnLbrW4T5Q5MmsumDeD+/IS9F9h6Mu7HtAioKm+62G+NAHDSV7FSXeW0/o4
B9x/Vokzszza+uB7kSwUj3mLK4hafHIwmknU3rfqWhJGDPrT+3p/f+ADp5iGlVgu
d+csJrAkCC84RiVjFrGcXka3zxQ9VZBwC1RsnWwHZPKtSl1g2tSOxGSBV+2jJKZ8
1+b4JJsypKFIAGHF72kNyALVlM0uWUtrtCZNq5Mnhzc3v4Rv/MnnHn4iRAz59lgh
UuOKdeeSEuqmKe6TEpBfBCyO2TYdPoN2FbKuH7O1uKW4YF+3kRAytzkLVGzP0pcT
4vnWhyGjTSiHnC5n/13tJgvefWJ9SyQJSMuhHQRqbPz6R8mgonmOkZ/XcOZiUiYF
AUF0xmK+eSBESB6wB9JOKlUPcwscdvcD3aqJvKG1YWLhkSwhceEsSf+UsWU46T10
E484uewdHbt3oHaoLIXM+nz97hhzOPRDapINf1up71CuXKBKcbEmq1BWeTaZNaYx
XQdBeRJk7fnVoSa7i8ZVZNTLdWn3ZpCYbL4U7tWeIQXgfA4szYuU76Xx08ZAXlfm
Y3+pmXVnrcvDA1LA8/u0c5dNb4nXP+ZSH3i6OfZK3SDEYvdaYE/cz+Dw7/7LJmGF
gTfkcTI8DysCkHGDK1g+5shCDsYAGahTfYjYxTvd2rUdel7w5Pp1pLmljUND+/xR
x6SDhVaJU0esEobfqFjVq2uQeGBE5Wfv3/7phlfdhTYnCuNx9gK4LH+5GWx/JKrP
KAk4mkXbRT5YGbL3B44GTlTd3qLlrCvbSDhjNfM4cpQ7KzNjll7kPmXNSYd71iUA
K3ny6yUQtkJ5//F+KQkYWIb/yzeL5enLs9h15nbWnTbD06sPpuRC11p3xq4vKEyc
hqWsZk7yx5bDzZ5JPlb8r0qF5iUr4NT+P2WAOvawGFjy1JbsgsMQo2n+Vqmhbbad
yyL0cZNg2jIoN7Ku7VkFpWI9+T0EkTfCDK5r13v4prlcE/zIvc5Ba1dlkQKSpbff
y3T27uMY+o3siksRhz6xscZXNQOG5xd0MSsq+GSeoTOd1K+ew7XftIwjBKsPpD3S
LbcaDwTm75pdO32v9lXIuve7zY+iZkeA7yO3LQrDImmxmH/yD+MJJYhcvMrddMp0
ZQFtj+e1msT27GekbLK/jJiUoyN1Y7OqXFXr1cPx52MkslfT3nYAbqEynmWp5cGI
FIENl8d1kRLqQfqHXzBaCxnRUokxL3WxsaaVMNQoHvs49o1JiDLu5/Ef4UTax+f8
q8LtWR8Mpf/ATsIgL+QshtUxgH8NIRcBD4GuPO6TPTOAgvN4E+/Lrm6I3GqcK8cV
d4CGBoNkklUPUjKnyg/tWC9mkgCTdDxTbjvE66jltGUNXK1EzAyrXxKlOmASwquJ
TYi8sN78N6BKqFAvYQ+B9l3OKUpXTHWrcrFONM3iN0HbLjn1sqZoDBeCMoz3q9cU
FAyh5j8d0uOsvssQ7MuQCuxkR1w34+cxdO/3Q+uLCl+erHJCnen+XKSLKAYzJl2c
Pl5zveDcryHRDsFa63lJ1hAxKgar9o/1OTY2y4em5XUT83zaG2PZWdloRJYKi2Ak
1fadLYg8QQMA4eD2BBjf84xwzZGqR7BcMS4VeNuQ4G6NPCYCqs10uYoD3/CR/EXP
DuNQvHC3CwhR35ztho7/bU3dj08oCzL2+dbf5mqjqR+PEHDRLd7AjdF+SFsttnrh
Qp9eegMVUrTo6ed/Xd6veJSBPjU+/5JlvmMsVAIVPtd2xfgMv5iF9+cJpyG2i3ml
72+HNX4rqP+XlF0EoyNmZPi3R9z772xLK+wx3FaoJGnqaUDcsTrI9s3OBs5tQiE0
6gUpvshIVbCtICfgNru70OH2NaIHFcz1KgOmTu8oa+CKAdzy/j/a7GSLJIQcgjLI
GsbQJYFoNJ3sLjCLUzEfPwIB/mJiINxX3eciNU4yiiju1XTHP0qEqBjWYBNUd2/9
uktnfEVOFByxtDEFM1+2eqdcP7Kmk8GObVCS6VpEbPZwKHQ5UGq2m5H/I5UyvgqK
NjmIJjsmlp4N6Ukn4h2f4+/DvD2K80c3o1qMG8g+HSh9EnvJar0cMxy0fJ5uzQsI
DnJopE0mNd55geKKlTmRRpXwpC7srB+QXSmR06aahe1PEKCDgCoqz8gI+9duu7H3
cRn4i6ClwwfE9JyYqPeUL+PD8XSsgCZyjZLwtEcVBwz+OXXEei3zuQNqzz4Fq6EX
uUqaVV0b26kAM2Vzi8i9PQAMhD/6fXyoVCDmvu5BhBGyk6BPOI0oEhK1omlpuU98
QDwBUVKC5uwd8+/1Z5Foc1229zP+NZX6NbLWLXWKgARl5OdD9ZwuQRe0ZOfK5Iid
mJZXxAhzCNlJmOK2q9ZC5+kL4+DEhSRtCyhM+bu9Oqw=
`protect END_PROTECTED
