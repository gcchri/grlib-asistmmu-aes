`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17XyZuUeldiBC1la9wGF7aIo7R20YeJAFJbTi6bva1IzKXZVqbOzHmqyFrzTZYlJ
UYszU6IQ5F89vaN+FjtdS+sjf241UR+60QhKiMfnfFe8VUaNGNLp4Ztl7aJQ26q3
aP0FJ2am7mh9wA7ZvQc0YexTaZsOxp8A3QK/xZslVNry7ipxMtZWrCmfRtPYS+z+
9StPtxNn0i5YGZSf4IGsSyah6uR4CeZKtbDRVeSIO3WDqDgOJYzgTC1eBLRCE+az
LoRWK4whgCRSR3BdkjoZJb+t8wgv1pH2J/tdQnUG+o/0YtcU0i+a/0TqAwcWEa5E
zZxPFnxfhpwDE52TyxU/GuLsThnkXpAmWdFi9RQNxfY2GXP4llNa4GI1s7HBli6U
sSj9+evJ17H2y2E0UeHQvXXMPQ4es5JJjwYJL8YYyFraFe7QaXB5ah0xSsD76X8Z
FlghkVCbpblvYKfiUWdpZixUQVY4drIP9Y4AyN5a4qFXwd9g5ScZ1wtpmKeywBvy
03tUDuiupzebBEJlDdZd1EtW61EAFlvQ8+WCmRZUBdYjAH0Eku2zdUkkw9S9Oc78
DazaLnUj26ZbPED6COM4MQrJWFeYTkLIfgxer4JRCnY0kNr6Fp2+MkQTtL9QaXs6
tnld2a6+2nbK8iECuWgZ01J5Vs5/O5HENzUC6SZaYluEhJXgnZCDkh3PU7dT5s+n
i+fIIlzED6tlCOV++O8mYkVeJkRdTkHeQL9ksvC10RDIO9PvP38XvRTXWy5R02i7
b6k2sAcBVkBIzT1QGOsf32Njj4C3agH9rcW0Z9X9kacbqqlROsWsP1DZ4alUuQvj
hOfsmxpmkJB9ysri3K6DlREvEZJKFTbLFDRrdeN3/iD+pjxZVj2HQjn51wz8or0N
nxN2k7qSWVH4jGOg43+64jS/m3JI79XAlMRbF07MDHeDUi1XNJZj3t5WfHW96VmS
6MyrGKwdsxfHrYn6dzJ8ICMGnCcGtKVOTZsbabYF9RU8TysLyphNu4Wy4Gt+yOaG
tMSMM2ZZu1xkznIO04M3TkXkv1COz8GOqSVEW5UQPumL/RGB7GsoEeQk+a9wAg8K
MIYbLzc7Oi4HThzjRJRrqYgVDs45dVmS2LMMeEh8GxxuKaYt0Qg6T/qIIELFEC86
p6WAD4QRTpUT1JjWm0mvv5hdIlVrcBt6Yc3VbfRisKimOWkTuD0z6+aYwRLsJqt2
G8c/Z3AN+cDwRpPROFpsn4BzgbkQWK4E+5kqFuWKIf+3nGvNtxKlHzkD2HjKC7zc
J1NQeit9bLlV0hMrbNAsgV0p8QZ2QB2ZhnLjDWkrDsigyIy2wWXneaA+IMOeASJE
Sfdj16kJNCtjACFmSTYq/Ebi3U7WVJBcuWRGz5TpvGMSZL97p6u4FSqXtrwTL2Op
aFZ5zPqT/PaNfP27IzcsNAXAZ0ilKOjzD6ogO8q2RH75lh5CBKwmhpHyAT+QBlbk
NSsPCPSNNKkZ8/tGtnPBFg6iUeRT9dSXN/NqYoOrE4woht4a0osGwEmOy81trrc+
cG6QfPkMSSy8efObY8vk3NF++3eOX0QRMriLyinGiMuNcE7FyfOQkG9GT+y2K1dI
/zwgEfz0nl531SqC0Tg2Afz3KFAQdscaWbi5f5j9fuiP392W+YAG3pmXwmiv/a2D
KQ3v80z8KDlC35IEIF+Qk2axsp/72y9qu/7c/8EW86UVr79ZPwcPlDDi5exj899G
57gO5RDDl4W9EEUubAKn0gWNzEHj2G5uhtRIsNgmFCOlrvja4yzjR9Paxyy2Jln5
jd+V7+xeFjVBwOTOPEtey8AdxufFk8BwNK790zmLlwCp098Rs+nd7VQA2yhOhXlu
Ik1lN8Xi6J3r0y74uLKIDHOM3lMxbOKPqdKwlRYochMen07YZXPyLs8kC271Dg8B
`protect END_PROTECTED
