`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBqeQNNcX1l19WoYoI3FEKP90tOy4pf4hfygYto3KhyEvsBH15HHwGuNPEzW5XYP
8osWIZMACJgP0djAkIkGmemtsdXOHtQRkhMtUVTlLkh/a/2ccY9FN/EuO+WYQI8/
ewv3zLsrh4Z2debrD3QomnsB65SN5jmVtPT2LGTZn4bvyGcSX5b4PRCSWLrOoLto
0aUcmzA2YyY5OfpU9tEkhwzjKBzlsHMnhXieoNJpAwW5voJN5Z8RJpNNpKOfbu0H
/ptmmEhM6l1GKYr53l5++M3cJinrXGewvDYmBDSqOcotccf+3ZGcspN85bxjKnsE
cf2eGeHAo6tqAcV5oqyF+nmIYPuzQMuvtQ/EgqHt0dqdJdE/8GhQgKLejM0f9cMR
aE63xIeh8iCYSVKQq24OOsT6oXggF0NOCnZ38lSOMTcKaPwhHcjnG9H+xrPRzJj+
`protect END_PROTECTED
