`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3F5TmjYp/2RuU23e+BbVyT53teKuQgtMmKAVbq0hoptvRap1T1KqDyvrnM+AbZ2j
DV1FknIHkmFw+eZwwEA6PtwaJjpIO61NiwtBWFmWcC8N679yVvnPNnDUXwCtXcic
eDAaH9KlBQ++T2VcEt5w4UFQywzIqaSas+lcOedfvgf0NTO4Q9RHjTFq8sVzDS7j
MMZdDTQO31mUQlBCItgZTSs6kI1hGSI5ehOj1NAJcUoTqIaGPtdbTRNATrwzwJYE
SuzEDzVtBO5myUa7kM404YHFF7tzYxU9/zbvCPWYwzavZxvwql+RJhSgEmLbq7Vp
oG3BUW1bJHWiXtxRyHQau/10Zp6hQe6LcM8ASJY0FR+u7da6svxxkHXApwbcDdFR
URzFx5ZF2hOpLqEMj3E4mTCvxe0FXb86wjoeQmxzSXPO0HF6cUmzbecCdQ6LH+dt
HQmjMJugkz+xQE52GCO0bhxow2sYxwZ/gStbON8keSQiPGql/sMmtR7COV+mJ0Ma
6NRQnipLHxC4zMyAMEC6l5ESsWEGE6lvCRXstiGMn4V8E3PZpCqfCKat1xCZifp9
Iyd8DRbvTWyNMxZlbRNdPAaoYMci33uiGQxDi28kFqZVNJ7r8CbEgZto2ZXNph99
YaaRovwrJbx10Y/cfPVwAw==
`protect END_PROTECTED
