`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gt2oxwqNoWRTzDUe/Q9mqZVB1/37DmgCeiVL/WAdH+7a6hLBnYQrvt1lO+llO1eI
oOyqUurmQO+44GiWNSmvF3FAWa6LRpVMF1rVkAjMd5XR3LXWdfZ1dycEWufhnkku
ybwHmvYHfNWbBqIYBWw8uZ5lvChCmCVotzOdO4GLohmJN7WTUvaI02cpR6C99qxn
ZA7NGswpjU0FMNTJpkp+V2mGHh78M9kFwhJVfgDrB3SOH1xEt5Ytq8iExguu5VH0
PE4ZC3l+kKnMA/luxsZddA==
`protect END_PROTECTED
