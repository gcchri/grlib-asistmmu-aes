`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1q+aqilcACJBrCSuszgwHMJVKgjQCGJTxW1C94W9JRKnZV7AqTuI98JLcmdH71p
WvbyxxCumwqBUdTwBFHXcC3sfFPmplu09UpgaITSNCxHFPVBZP+/moUUn6m8/jh2
dnxN/LrRk7txAZJ7/LSNYmVlIhGN/bkismd9Ror5oFwRnaItE/A9v+C0uqPU/Gii
30AjHNBykQZQo5yQoVsOAvbq/AwTbDARPEvibLnAF67tiiMevohK5XpNYkYym5ob
4m0JHO/O6wT0CoC5whXNIu5/sGGZi8sm1SoEuV+0Vn3JQirsGoZhEHyziMCDiY2F
BYjsmNhPG9a9Hy4auCzx5DbvrMUP3ZU2BBppnqNpfPgwdI2X4h0lu6A8qCFgqjZj
quHlhfblcdZ6f3w+w6tOpK8rkPXd2M/qzy7x7ABJAC2tzcxtbaSKz6s8nRvCaKDp
DSsiBeto49sFUrILaBcGj2Ee5w/oHS6uaeuGmVaPr+H5eiTldXgtFUrt/Z/VdFI/
7P8W1HCR8xbu4FTHmd0OnQ==
`protect END_PROTECTED
