`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cLuQtjKDoQLS4Qr71y+xdNWSsg6zsm56ebs3holhoiQp1tMOrMKKxlfyto8v7FY
rl9smErlF4zS2+TRV92G1IGIaiUSOHbh86N9Z0PRfTI6PxfMbizCns3zyJR9HyOC
vAb4R7jMI0wrkNxMn+tynZ2xnlIKeqdlnghT0f58qrVWZRscw8tsTJSW8w/J2Uu0
OYLdVJ1xV2zdwfzkx8gaUyKCf9ltOdhEi7nrD8iqyWD79V5ukvBxqOBnTP0cITtJ
FY6c8o4xT+LirXdhCrSHgNAhJ/qe2cfMA71zcO+CyL9Dj1P3LvCSfuPvNgnMe6t0
WLIvw1Wee8HMK1sghCQkHEXKhYhLAG2HkXX5NrsSBdquOszfdxBxz58VD0j0kp0z
wuRjvG9pmv4e/MvmzDGz25lAFRhhOGfM2Ut3pPjMuRLITGRhcyD/FoVj4Rn1AgPS
6Ox620klmzpwsv4Fv4IGAKPCU6oIYES7Y75f3TYbLOV+Hrx+OBSD/bhfd9UOFqk5
TpERvQpWBpFoCEGWpEpaoxHbvxlQCNV9NuXW5ExvY1wD89BNfsCLp5YEPVRdtTKf
oNs2SC31vuocRolVqx1efoepHjZur9trrQeyg6XYttihG+CclLDmthLmUxA1X+4X
8V5QhIVvXngD1g0BP/oYJc4HZiE8XASQkeQPwnkM2OEBNnziSxycq/t8O7LaWr41
VKgnMbC49Up2au/R/J9u2wf/5ppY2Lefzc5K5mFFmNo0SPZhRynfCIajmLiJ1DtN
A613D+XH2lfr/5gSVEGMx7xzbCho4WpYtoQoK4ibzl01oM1UaUBzMYTvieZjSahK
nAm40kEaMEvieg+Rp9F94d+uuLeAS6TDi3Yea4J0BusM+cowBAxS0J//PiK2qqFV
z+MlLy4iwj6CuU8GR/1SIWgRtkdw4rj1oh5cT2yX90zoG5Ea2eeSY3Ke40HCS9gX
Zo+F6OrBnVAPTamt8bvXKg9ueJbMCe1BCol6OGQ3aaIiiZeJXil4H1VJSNco5ZHu
m7NqxdM/BISVYGSXkkPl0TleVZFwicUQrUgY51XYs+c4j18K5NM19Cy0jRkckEm9
+8oYjOz+zlO3bIhoPzOYR4n5wqvJ1r5aXY9o7izKU4jWXBKjBADFVqsJvUmWZUr2
Rp49yEo5MRRRmOu4QlsJXY5IrUkKbqeS6iy8kTVQ5U9si5mA9+Jwll/yXbsbNjUr
fQ0fevn9JVcu03+oyslgSKwvp6rP28pDPITXPf4s5hU=
`protect END_PROTECTED
