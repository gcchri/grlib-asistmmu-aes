`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
elHUZxtocvpKWDbpOY7D4bpJmqElVMqhIvnKY432LN+JB3vv/fGnyXSVxvFJ/T88
NRzn7Z4s1K83YNz22EhgehjUpRF6CcRMfDUXe23EPoOIU0D09Bq8a2U3qIFt3/gv
9cuLMt6G0X9GfBpcrbx23Uc8x99ZPTGoXOw3h0ZLTjZXrRcTGp2zGdW0ayMmJDyD
GvIVHcinYHWNkzEZz9s9kvGW88lbqqswhmZrutLaqw4ehHaRhv90bt6K6LfMJNCH
lYiW/pytfFCILCZNDDIzdEpUYWWVqSPc/AtrKTeL2p3G/uFkWWHhtZiX2fRcSy/P
zzfMieHktTWBiTQGX2NhRMyTKLBdNM3liULEG9QOVhI=
`protect END_PROTECTED
