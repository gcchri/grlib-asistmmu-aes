`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1q0KfM/wotRwsEfDTuaVfpu4VzFj5bZLf0fGep/COD5d5OboTuxy6g3bB6Uz5tzd
TWD12uh1hB28I+X0e96Nea5FZOOC9bTkEYBITK/im2W0mr52gXNIYHY5KqA+tqSD
bPwUBRj3VJSHufqDD4Hpucga1uBh6I8Za9pygpRFw6UF4pxW9yZM+sugo0SzgXKe
FI5NaTG0EpsZSY49Hb4KszZJnJEmFGhMbrV5fiV0PLPs/qYamUYwLsYZSuqHlZRr
Mpg7P1fqVBZBY9EvFokbZdia5GM4pVMWtAle+RGv/Nqr/HXIZlyv7RXK28KJhxDK
6ALDBp96Lc8+WwsT740F4dXa+JE+lOLlKzyOy8xLjaWHbwxrN9xWSZNC328YTbdt
uxZEZCnMddp1DaI04z1fSxdlm3nBbNbvMcDGCaFV3sLV7P1ngGyZHfmvX3dztKrm
DNkjOxWcL4Nlu2uOXwbIH40xGjT0S9Rd8xiPiuiwTAAxP/xzl5R1v6sVD/SXUaMN
MulOph3Fr5RpCiiGMZoD7C42Jj2ziffajCo1jukUAOn1A3PtaRjGhYT8Jzjya2xx
`protect END_PROTECTED
