`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2L44x6EjhgJEtQHE/rBwN5um4du244XoT8h9Ho1zsMSH2OBN7E1u+mNkGCVD5xv
yQWjw9yX0yEE2klY0jpjO7iKP4yM9+mkxJwVd0sLqjVKFSrsG9bpSU8rzPL1sg8y
TzPg96pXZvSW3HAZqUA91ME2Bbsc2ZkorJOa96umYA7LbbS1Iit0r7DAtnfbUDIU
VCylvKgxfDQ3Up4rsyT4UrXJ6cIHhuLXMUGn8Z7x8AH5f+g+L5k9xqgjOGzJkleO
JjVJXWl71MvBq50j9S+N1EhEEmWZUukH7XqVRWGEP0SZl6/H64gHhS7KnlivFPWG
HOk7LCgmgiwFjeDltsm7nJe9gGC4qt5AVG8sC0sKGvuorpPrZWEGkDFwA6kT/2C2
GF+jMQHiS2FuZZ662R7LrPg1GJQHHiETcqoSlwOwO08ZthwPIISGr0dDk42EfJk3
/Su3KvienvWnTOe0MS4FUbTDmCnmVvZcApo7cq4toqkNIyeivPTIxGgpiGmDyCgj
PNnqSFI36n0svCrMfcjBL5dQLtzEgn2MObROIZlMvfssX8tF4j0IK0cEBi2CVdzs
eyCICS08t8XsYqYpSWyQr91mk1Wfy0xjlbfHye67KeFcKpvyPE9DspLkuKXkKsxg
0IhiJS4Q3FpXscQmr1BP8O/ezxnopAECzdNDsF+TAulplaV2FqapQsM6JVufXkjx
niUMDX5xwj2Hqxp7S6vYYXQylPO/LFBx2ADUZQweV435Vdt4SOstmPGMca6Sjkzc
URCZMkqA6E9E9vtJh6rJk2VVStTPqhX76iQyliTvmgjWf/tY849ltMMvaQH4Jrsd
saf/5tjqNwMEGq8CqiPXe0VE1rMowBeUkm3DLWvvasyTCrp2B2yRzqA6jfWT0AkS
7TyKwjPTHwPat5vQmBNsvKzb2gcraofdxQilFujbvhWIxBV0c8/gnYX1/BwXms8y
NmhyWlBa6MAwt+PBFtcyd9vRZHBY2icvmzL/JG4JigLX35bGo4bYX5wRbSEwFGMu
NV3G6J5oiXx2j/OXswmQRtzETKD1M2J1Ki0qLR0yAFbUB5oN9uVloJhWAzn9wsu6
4+LsABJLEZKYIpDfQ001kMb+63/7LRiUstoOpHtCG0vsYo2J0QdKB1d78heGOJY4
xsIWmNwvTpAvYM2lNKZhA2QFH/tW1nEzfiUqCgalgBjbNbMgr5omVHaDlxzlr0BG
c6lUH2PW2ibCb8i0iX175g097Bg3+Qv3BHmAZZlxlwx7DUbo4vKawfcx/dbsKJBk
Lb2QoiQ2X0pNHkmTN4X7OA==
`protect END_PROTECTED
