library verilog;
use verilog.vl_types.all;
entity SIP_IN_FIFO is
    port(
        ALMOST_EMPTY_VALUE: in     vl_logic_vector(7 downto 0);
        ALMOST_FULL_VALUE: in     vl_logic_vector(7 downto 0);
        ARRAY_MODE      : in     vl_logic;
        SLOW_RD_CLK     : in     vl_logic;
        SLOW_WR_CLK     : in     vl_logic;
        SPARE           : in     vl_logic_vector(3 downto 0);
        SYNCHRONOUS_MODE: in     vl_logic;
        ALMOSTEMPTY     : out    vl_logic;
        ALMOSTFULL      : out    vl_logic;
        EMPTY           : out    vl_logic;
        FULL            : out    vl_logic;
        Q0              : out    vl_logic_vector(7 downto 0);
        Q1              : out    vl_logic_vector(7 downto 0);
        Q2              : out    vl_logic_vector(7 downto 0);
        Q3              : out    vl_logic_vector(7 downto 0);
        Q4              : out    vl_logic_vector(7 downto 0);
        Q5              : out    vl_logic_vector(7 downto 0);
        Q6              : out    vl_logic_vector(7 downto 0);
        Q7              : out    vl_logic_vector(7 downto 0);
        Q8              : out    vl_logic_vector(7 downto 0);
        Q9              : out    vl_logic_vector(7 downto 0);
        SCANOUT         : out    vl_logic_vector(3 downto 0);
        D0              : in     vl_logic_vector(3 downto 0);
        D1              : in     vl_logic_vector(3 downto 0);
        D2              : in     vl_logic_vector(3 downto 0);
        D3              : in     vl_logic_vector(3 downto 0);
        D4              : in     vl_logic_vector(3 downto 0);
        D5              : in     vl_logic_vector(7 downto 0);
        D6              : in     vl_logic_vector(7 downto 0);
        D7              : in     vl_logic_vector(3 downto 0);
        D8              : in     vl_logic_vector(3 downto 0);
        D9              : in     vl_logic_vector(3 downto 0);
        RDCLK           : in     vl_logic;
        RDEN            : in     vl_logic;
        RESET           : in     vl_logic;
        SCANENB         : in     vl_logic;
        SCANIN          : in     vl_logic_vector(3 downto 0);
        TESTMODEB       : in     vl_logic;
        TESTREADDISB    : in     vl_logic;
        TESTWRITEDISB   : in     vl_logic;
        WRCLK           : in     vl_logic;
        WREN            : in     vl_logic;
        GSR             : in     vl_logic
    );
end SIP_IN_FIFO;
