`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVb24A8cpqxU81X44YhJ9WUf2epWvSNRqFAz9iFqlEH9A8OQo9I0u7U2RiaTxA/r
YrZdyK63nx+dFkcauskijmqOnKZKiqOf5eIGCxaD3dkxNJTkeYNCXrqvHA27zf/G
5XyUGRcxYhWwmwAR+y/kDJmFnoDQ4vGjCRf/EBNupMvW8EEjoBTou0Mh1gJyRpy1
34J3DbbvtU39MgwUWPXskixMbNzK1lf48tVAY6yuzYqQ5qLnWCLseAF583zi+4BC
WPf7jDY4888Qn0fUdq/kxtCf1KKLDn/02R51SH1f3eMuM4T6IqzBBTEGpLzVmyoJ
/h7Kd3FASGlQCKqxn8X+wo21yH+zAZE0MOka0pEvgaYZhkL1VXU/j3LWlzo5zydS
qZjIpyp4N8mU6ZZ+F1NRMAuy7jO7SOqdZF6bEc94pi3ds6zfVFPecSNG4izHehnK
xzBd6conIbWHSYM96gUqUvFnRWKTJ8RFQg8xFBjZb0oHb/7tp6OW5EQczjhTPNdw
qCwmieLzilfS/FAlV8wKjEK3J62gnuGw1IXEpJmx5553gdBU+Iu2ha/SrQZXlB3Z
nxVq30hY8Q7J+wQgf9GIZqulfD0l+RnTNpCRHoobBENh4z3N2NvIGKCzOSfbD4mf
1Xu/UnCAaC1WGnrmIQMjUZH7ycqssdIbVOIybMkiPxGBLPWgFK/lX9frTfUa01eh
jQgZke9DBjKeggZNor1WAXjKNx92sgTB5xGHzJw48DiU0FS+5YBLoLh9tDnhJk3t
dvoOieM5jTJk3Svu+pjrplnLKwnDifMnHZdNSAIdq+PPa2xijakug81SQivOQp3H
925bWhM90cBdrsDuUIDaytj/FW2k4RP4au2VwmFHh1/yM+UM/uxeF4VWnukQokUR
Fw17RhbXiwa/rdC7tPsFMnq0CIDND2kdjJ76c6P+WJ2ShT0Z2gIu4UXOuDD8NWqa
Owjr+naYZiHdAdK+ItS1DdQJ/95+BUfWFSoR5UxOC/bNf5mB/sWcXj3y2Pv1gPXb
c8Th5ZfpmChG7OPBZ4kArIPrl7Gol3Qsqlb6UNsDm7HEjH5aI4FL1eEzvE/09Q7J
aoOOZnbQJyWN3tPkJnUtVv7usVHImsvd9/zqdZyG8VCAlzJ89nQj+fKQ15/y5v2b
v0yajoUeeTs7AfGJ2+/b2XcsugSlK7sF3feoMmeu8Ew=
`protect END_PROTECTED
