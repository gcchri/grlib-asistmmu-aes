`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jrRESEgB8Kgd5RVS3s8kA2rW9ymN4sugSGnu/CWr699YeHqLYa5mND5s6I5JvqV1
RoGxFq55nkStRP8PE06dTATsE8xa2JI9Pg9Ncwpp2uHWSj1ayPXbG+IJ2GKInFS+
cS0+FKzSc9QTl9ihY8lNBOgSZyqvoCT3eum4VjeLLGLEx5YIQm/wL//NnYh9Troo
IEqlxzfYgHuLzHJ++kI04yn1nXtBEusoQMLYLERxpT+d7YRtKVkExr0h6bKj6fMu
uw+wGCZ1ebYdq/uT0IUe+C9zNDgk0chQua9PC4HKzTt3tQiucyG2sWrXcFkJ2QHP
6YTUZ5aTqYn1/dpMdmv423Rc8H8PdDaEdF0jaSaYWZPkjWj3pmgtIAS04f5nLCVv
qJ555gh3nGECqsgYNC/mMjzU3YYGV5/LK1J7IQwseYhlAh/t0Qn37CKY3aiqkGKH
Dkhkgfbnkn9tPEE+hdy75nSPU6W9B7cMWdwdrUDdOb7Ztqhzhw4zhHYrvDeArL0F
sGWPcWwkfnuazuAW4e9+rw5YCMecyx35EQ04FPLxU+KW+nnQaPeRzS1aJ1rrYH0P
3dPlh+U40tc2cnc8OQT3U703hOtD4hYndyp0CSSaJ0wiChYDeAAuj3obUEVy4Cvo
FA5LyXn23VNo+122k5/Ndg==
`protect END_PROTECTED
