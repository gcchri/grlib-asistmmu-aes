`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LcXzmEVbGuqS6Fo1j00ivISDUO49exmWwAO31fof2IWWv/p00gzImCzape5q1+kH
tWfyiZeM/UcbwO/mFze3Wbe/HDIxxEzP6o0Y64OWni/eX54rp5EvdikrKXMCPjO5
UUYfxFpTMhJvb63sHF6eFKsvGf7S5PIu5F2Bv9zS+YuXgaaCjg5kxN6DNAHs6EUP
nUlZGWZ1/Yf1cv/GZoq7xzom+t2KVrC0XW8pFrNHaIRsUazds9BwP1k72Sk4QMYO
57bLA/rY/POPrMBtCPLk8acwK5r3US6Dk2JojDkYchumD7cWBSCmH4LGRO/yfFFl
l1v6O5NeAlJBH1HTHp1bGeujv61rrt+oh7/9+k9yj4WmqBkpJg7n8SrWtVcL5JEi
zNBXlShSIxZdhDvor4TGPVgCzskI6MfW9QAdFcdVXCxsLXZnukN4fbiLybKH7ZoF
H3ltmZ4R2B6M1xG/Qr2bPKNyYv77znumEY7OjxBjdCGW8go/zR9n+aNcSyWR/QDC
HNhFGN6iz1cx57/NMKwMssaIrHqDHg0yShD5jSqWKG7bRlKShxTDoAL1H0RKStNx
AvQYxj1jwVNqHGYnWK/X2vrImEfwuGOBKiERiQUbMws06Yh4ec0q+l1tBiINRS9W
werSUGqcET26BQZUWhHWeTU+AUX8Y7OQV4kExYMn3IxW8r1Gz1ISNFYed+yHiJ15
4cpdFgtUK2mIYva8bmd9aTgRhNjXD8tv7s7F2FQTkEdj48E6AfcAdxj4GYJTdaVr
q5tlydFW2LhmsC98HP1jkDwxBuSFaM20uxsmo/t3hiYp/wE7sCGG7fQmOLKC6XbS
9Hwbi2o80Lh1G5+VoonA124P8MWHQxgGfSY5raI8kDlLdMb1woKaDszAh375pfEs
6fHgVYd5oB5n+Rmn2Ayt5E2R9L55fxUzgY3Vk4Ib91CzYgAsiEN0cA9Sur/JC7uE
NvRksX7Zh1bGHY4xDhZbbnYdXjim7vOk1aAAwHdNpAKFRCG27LMP1ElRFA3zHpdz
E2+J0wOP2em/rDsYPPwvDa8pYWkCTC/Ql7E9luTFF5uvaf3BYBCkvAJh8MW95qr7
6ASSaxK6BybaBYY0eTD8Stlp+KPW5/7zgquVAfmOwJvK34cjexvDaNsMa22OPWSa
opDJAgGWiQxP7KbVZVJkB7WCGEFz8fU0Ree0PtyeQGueyzBkiz2Lq0c4AEkpc42s
eDkQ3TXvDpeq7UBj8+diu1+xEU9vk8BS0DUgiw9U3DcT7QB9X/8UlR20muf7sgiS
pqpOdO+tg6uWHDSbfor8uWVQXAconNwyiRCTllENzTKMMdhYovWgw8yme3v8yVN6
fOoMe62b4Rjn4i2sfWpkDTMfLC2FLNmoLvDRUXTSYR6E1y2rB8sFcKBkDlhCOtgy
PPlJ22mibtGSGuTpX79uUQeUsc/FQ+CNvnyEONq27AkdxGQrLgrx5pDl2Ajiv2dS
QlJE0OeqQy+IJ/INHpjK4f1S74GmB3vtEXeTLTumsR9TK+ONGJPsbDRtVwc3czcx
MyIT8dIhDLkbtf0nfIo3X5YL2gSaRKaRhIIQQ/jIdpiSETSxeUcA/ayePFwYh7Wf
bP+SY3soy/qDp5XlYkNKjzEMCajjRPokvuAfe55Ww1dICEDt7tb6rhixD4J2u7qM
m37NcDq7OSaaV3BjAyNVectFBHeJwss0riTG233aFB8aE0r636Unaz9mKXzC46xi
YT8pWTCLtLqD8TanEBicAviVu1234rQ217+liLZszdEKmtErIQOyc78gcoFo1ZUf
1XIwoF+gbXr7UTIa5UBz/5N+ccLzBVMoiOFoPeq/zclzXcqtpIQ2uPsZxCVN1qk9
KIxLItCqlvTha/nOo6SgiK8HnDdpcUX/FhrK1E0sPYipzsYXVqCCyq3GihzHYXaq
WRNexuuj6k0Kmxbk3LBn2egUf202NdzFZiPVhncjlB6rhnq5DVd0x+KZnEonQ6hO
dKY1+3C2NUUN8UIx++i7EIUlBxt4mpdu6qVnUcUizla7Qh5DS/MzyOruAg1R92oM
Oi6C0CTj5D0ea+rVO+F/7Z9H59Wa8345wv+gnCrSjfWAJ5K7Ir3NCuPudo2FbhNq
4oFJguuHB7o0JXgUUVDVj9YCgIw1e4R3qHtg0WZvk0DFTXLUlntIQfUud44m0xrF
eoRrV9MQmbN3AP/28R4GChAAO8ExwQNJre18hh+7+7vwhyEhrWhd5mbrKNmpRRhl
7TU+z6YPpwOPDui/9rYLM3x+pOX1zFLhlGi1E065vvRHwSWbeEpd1E+jBYpJGPcc
cJCQUhWb5jtnsAtwBhMNSBeUkFtnmzZCfyQa6urokhN/u19VRj1K6enpC6Qj1HPd
RqzbnRWBE2MkCgjYiXrzM3q3c6OAO4BKOjBBL8+i4LypZGXOdWo8VquucXakOLBJ
xtF/EIt7r6LqmAXFzoQn6xpHd5lEvY2jL9cb4zkq625c+GDbzyFTie82Gq8DdH6u
r3LAsM4+VPO5jQ7gfeLJOYMNFdTOMe6z6S+qVjrysdDt5u3S471CffBQCzX3WLLx
dyuHQ9AZvGxOnLCdv6EDjPAXv7uIJXdiUBTl4JCpWQSpYB+pA4GWQzw3ImDn/A2A
jKN+o5gLpLSlanxBBWBBgNvm+Vi3v9Fja39d74COF3LP0/4vjO0HhfYbIMFTy+71
FaPI861K/1eVl0cJbIySD8FqoX6172Kc9/unzafvjDvZISZBgaMgECadsyJ8nAXF
QB5eJWss6jva+5xa6CiG94jjBL1i65/rIa3TWOibxE5M6jyj4Q+H2ZZqLatirqiU
Sp+5nwDOMfAKx2uweaAL1jsDTXH8sPB7nCQ4tHWe1XiZnxy9PxJcGCJQwxLm7J5s
IjvCQWISFDp6l5UTOBG9ZyO1ulG037QH6WcWKNr8pqEgPJOvr764aPCFg6eTddQk
Fh9f9W3+nSRSknIAf+4KOZIWLI6wQyFq/d1jZhKZ6P+7ehYW/JwRuhfQHaOZpSzC
heI/c8RNWfh+rO8H4j25xs/QRuw/ituLwBWAzz5fkRT3Mm/F9RQkSdvoEz4IdvaY
WP418bH3gJvG5eEpOoNe0XpdxbnImHBAS6q4hFcQrw/uHBYYpiGVE2c7V+pQovkb
ETn1jny9ZKE5M863iXmKTjYjjHqRF4E/Y/vNYEtokbY/MwxaLC5FgTo3ev/Bkxfj
bA68spJTulyxFvV/k6Ev6iltHTRRQGhAoI8CrM2emC4MVXKuHKgdF3GfEf146+bZ
uP+BDXWan5y5fbZdpD5awWMIqkeW+274xbDFmkHdHHeCFSh5Kn++PZvk8iqbCIQL
x0lrr9JM5ztWFd/bB4pUhviLmFbon5FhYzThcvIRkhsalmC218zxvHBpjgl7owqf
KJMsESKOn9TEzk91GgILEzs19+DE+rJTK6AA27WYZ5Ct3BHSgkUUoJPKqEkIRDtv
+9vl+jmdsIW6D1/P3Vjp52IwBX6YG2mCLfnn+qZwEjtdokuYRhE16gACnUg9KsU0
/MOoSsVHaiIARkvNoB4GJPF9wexy+Q2NlCAO+3jMDpaNXNtPm8L2sl306JbeHSZL
9tJASjujJ07DVqOXG/bT1IBaEW8uhQ62YGVsDK9RCeJH1rYQyA3HleJ8gZqGIEgE
Wj9KqKMSUzyMeoVHTiKvZCZrvVO89N+FsXy83RG5nJly3PSo4Y9iVITLfm2Ig6y+
6U6RYvueqXo65ZIwN8XY+xs2d7HvPT9ynGsFZW7rz2QVIRHNQe2QnAaB5CSXSg3b
9fO+GQBTGmfnrrxdtzxkxL5AcRcE9jUNIusFi7onRvZ+NF9VelzYGCX/nm6aBVPo
eqsHOIe3vmtunDdY8qZwiChGp7muHx2Chc2oPzFj+hIl8nxN9ip0bcAelbgzzAAn
0RC2Q75l9yBU2+/C0RwZC+XZCskKbmJAQKTyPBFZAyGGIL5KyqP3LxPAmneVIcdU
MFU/GA8JrQcbezjEA7SpN4FzjwD7sJUV01LRuUrRMPS26JJt75+jQ+QnLdW6WXX8
8GdPjVQMKbH/AEHkXmTN86/IW92yASot+XzMPeHpaVjjvHKOC/bfcSXO01I28b10
TuYELeLMFknhrRuvUVfHcR7AnNaDPQ9AwYHzbzh04R8+PXWZlRzTHRWaPRBUf8SJ
003rjoHwOL6KmMO32qKMcAOFgM21bK2jwSkq85FtSt+y+ek6HXY3+rIIl9yROvBQ
+RFaPNXVIMbx4IEdP55Q/gWhYoBhXPVxs/7G8w29246vdJvqEEKDl7iU1K4Njzb9
x1ArVn90RAnUoi5oPALvtOyAF44e1Y4uY8dFeq1yReKO/i5CpmQfJu+mKzli+qMt
eFEGZxIhJTt7TvpNG7ovNhErHp/Ii+QYgrq+XmQcbR+I2/x7B1Cy5RkSlNRhamxl
UW8d3nm/S5t3AvOb9FykePnpJgg6qUqoJ6Yi/GFRDQiYVmdzfYz32uJ39PS2lLDe
wxDVBkahWSsQvB1/Ex2o6DZPHMjeawbuZB5Mcf2lqcliU696J2LcV6mKd7lnxXSY
OvA+kFnSXZhJAquWd7F2Xc09VoSsKM7inUE4iV3Q+mfAyZKBni5MRrEJ/Gd2hxhD
WbS92/jj3c9KKthahSqKQSk4pYhj4LJKSv0GL2UBGsTOtXI5WtdX9nD5kuo3UvWb
zyPdGu464aPjI4Qxbfaogay5f5IJ88SxrDmkfJr+TX87u/Xekd8fYn1YIWeYXPkh
et2+NT9c++xbQgcXXJgmcalcs9VktJfDnUVQngywhJFvvWnQNs2KsisAXuSMbW3P
MnrRmjZxvrYtlIda1HqD1NhSsqs77nKBDxqww9cjmVjhwACFGQKLGKxv8fkZPCQt
Bo6xEWtppCKs3DOvaMt2QUGskb0V0bDBt7+8aXtdgWoG+XWXhLo03EJQdttOLVB1
JRlBGQz5Mm7EkiKOYaI/s3h0I4FMY4CvEro1QdXUmQJJSQuknmemymaRIEpk5T1o
vqCAokrg9IHkegGGAxGdhmIB2YrBLf+b14ZToszK9nVr+/L4qmt4xZQ7zctVdl59
gNxzxQsBS1+Yp0fXUhG99GooDfox70GoKy0vRgg2Vwwujlx/j12kW4FWltfO9sXb
UtTHt1dKOXsvZ2KK+Ib+CTCHd7pOYxau0DK1mLZXox2C5e2Aj9rz5m92cC1SLKwC
hjij3v/qY+rxyHtbBW05tWSxsvWAhJ6/NxZghhP15oayclwElfx+hyIuP3GtjniE
z/MLAjaAG1AfOFA+WEcmd5M2I016QH4Wjf8Fot/LTfMHcm/P5wQUw8SOQrhWnjrf
bp9BVga2ESnAXXjtACnQHSTb7Ntlei9nLLBhaMtCoHT6lXttz7OxUP263iTzQ6N7
4MORDO0hpifX51CiOLsxV0J8NAn3mqLRQMNmY7k0PQW9I0JP85lA287cwwreIjx3
Nqj278AcduV0rxBBNLINfkz3f9xevAW+pW2V5d3+AcMhWvL2IuZjvvElSTMBomBr
7rOzmkvMbxPGNUI6m4aZbyEZbPLswvDLfaMRkxshwkGXIsEwz9PbF/MNYKlfOZQB
O2fha5IsJQ2HiUZVHpd6X1J+ud4JBj2NOlKD0dl+3JX8hyiRlmut9i1zlkUHsQFH
KN7ar1CqtT+61sD1HuQWufvv6VcgApdB5RbAYrm47aIGCvTDqG1gn/Wti/XCnRlT
tSu/nyZTqegrnt9C4f/5l9k3Sac2nokyXqxPxJ6EM9Zch4jkKn/JJScxD0y2WueO
qXYtNpAJclPe2Fn33FBX8wfll9bUmZBFjDEWTJMWX29/WP8Enu4KAfx38s43/Ndq
z7C4F4GSzGEAmacs4LkLi61jzs9ICfdnTXapTZV6w+ia8z1hLLV2pFnWiISewRVx
c7hQfg7kwRGJtUIGcRf07O7NxN3gewhYmVoU+JdGmRQWLswxrDDvAwGFJvvzpY4E
cT04Fz39e/wAq6dOwP29NvRO7oO6b9wBsfQ5jmpnvdGiK1ziMUKDM6hCljnYzlsG
Y1Exr/OnfFCyKzT2QYnUva+/jz7P08iXyIq4p0hnqSA7FMm4n0Ek1R9kc5cFnEsu
38Zd96Z3dxev+oRmKv3XQehz9YVaYmUp6/JdI/q3e7w7xni/89Pm237aXSBc5jwG
I8LLLepXFkEFu0FnC8ufTU80cW9kOmIQfYhYs/CIPadpgbaF+Tcf4Sh4FhqPdiCl
rv6baPvYvzoA7KOEMiKCOA+eAG0nhEyDyUODGIH1rYZRNyBgKeX3Yn3+ExkkuhJB
MNOHl2A1ZJvvqJU0KLaq7SCrQ7K2ywNY/G7c8t3MBzu4CzjLm8l84QocLJ/FCZOy
0nzaJLMlXY7iDD2W0RuPyIcOdSft9reXriOYw7F2fLe1CZVF3OYIyIS1Ll9UELDM
0Qnq0ge/QHRFRXZJyipygkbSgjzfUwrrsz9q9FsGZBdlcqKa9AIX8GcoCEit6VRz
PEKdZBkWkrH5adv0Xp1O0Gj3u8tGwrIVbipKns91Ba7Jp2zc12j50eQPjvBkoT3b
rE206jEL8vCcTDuz1SaZhHlNxwY5wqiuDCsUBFg8YyK7+okBHWEW6FMz89owJfuH
SbRhCBqJuelTBHsV9ghE/vWnI8RqkkqLEvDrdOX9QwfnXkQfXSpf8JscDDQpzFC9
IDrpzF4IB0rquXgEPk7MjdA9COLQzWPagcGYjEei0UicLLgx9y9YHnasIBT9K6Mb
z6JOn/A2aFCJAy3XYhAuKJlQz4+82Wa73a0FDyKMo4Z70vdO5Xm69VD0zBnJDjAq
tFUlveGdxrgUSG1ErRH7I1s2BxHONAhCAve7bpylia/Ymlt4dQ54u65247z/QReE
uRxT9i0dtBcV40xrgA6aUtWDAl9BtQSvfvavpXuJ7TyG5cg6n9W6qjX949sCd6Qm
grUFDu1efyeBMK8MjIr8TA+cgIIBO3mawjTNY9wWkK6Knr6kODsRz1FmbklEvrTf
iq9K0xB3jRYVtjW2/mR1hXBU6GTfgPvwv1OgAlpTPKfxunpYLPAQL1yVlgCMxSjD
8hwkPlv5M2pMldOASt5jLmO+2LaHCur0BaiCCg7Ng0az9+4JHv9r6k63GcXjQyyp
gvpKKVpPoh1gFMW9jh6fHZyZApgzXX2UiWJ3XhJba1yPPFasvGTjQSpSGP9FrjqS
v5/O54q4DFQNFFJMMPQ2rRwPG2I/yW3VokgRrgFgNeBWCeHgY6OIqTZLLXR8HD4f
FGG7KQ7Bqz/2ZtvfmfzfPKZ0QODQK/ef+tyQq9fbT6jDEqYDLZ5lNQ+OXmrxiV12
KnwSYjUrax6T7JKElu6kBheVJq+as0E5yG8wbrzXuXRKZgpiS6ZbUtdmK6yiZexh
7bi2aOuXO1hc/UN5yd8RR5lRlhL9RWuo+fLi9GSZyw/XgHpt6iqF14Qm43O5bXbR
Tdt1WR5+7K9YhIYQHcaHghc0Cv2b0up8IEkme76MWwKY9dDso4rmIq+wkKsuO8z0
LckIn5QCDRlyowloew7pj+cpbAYNyI7aSarUVp/h7I964Tueg7wxR6woZYoroy41
6zQmcZN/wiI99BSLw0k5X0HBNI7ZhaDuGyqTpdAwCguhmk7aA3R4xW6mV4k1mX/v
E+xrA/MFmvJpZWUXt7m/S6MDKN2W9VgvhZp935AQbvScOWLyWpfq+VxRC6aAxyQm
QA8Z/ydLVMRSqlTp42y+Cc5o15PtKjwbFj2HYHqI904KhVP4digPDE//h4FEU30s
XqlNHvjLwhhdICxBqtOKhhpyH5cEKdhT1Da8bo9qV2eJZL5ok4XJTRMSXdIp8uem
uAa2UyEo8MAAu89Hgw2FgrkELSCYFAjfE7UT8sDUHIcudMz3RtrQbDt5MUT2xn3F
qQKN6Fo8UTSL6954JGPSwCAR3RbfjB7BJgSluvFis1nqNaNjiUcGzlUs3afth4AG
n9EAvytncZFGk+fe05edXqjT2r7OVPTxagrDSXS4zHnnuMk0UqGX4XLXzP71+bOV
CaY8QNRJbe68uJ5+IulZEaR+8w6CR05I/N8B4FGy2Es9ZQ7kGWGN7cCH1TAQnPgL
pn5TYgXdiLCogi0Bj+bLdB1nV0ZD/7d2vtcSFddNH6LdApt4d7WV3z1fMOXrIIcX
grbEusWRlyaRoNnjgg7e6DMdqdI1lQu8G8JmfjsS50RIWBHmVZ/vnpCfUS7soHYZ
O2Wul6BZOgqva4FUObmYwFrNCKs4/FjycybfFT21iIvNiTfjumtP65TO1c14M58h
vHzsj9acJ1buCw6NMxvu9z5+vbM040SAvKYf8f6t0lZ8I+5fBqSzApKEVSSwQ/gz
8hOqwmJB8mPMDVmDQbRM/zVXXyZV/mNfcj1jcXm2EmOQkJ2GDmg+j76jY5rAmZ4P
Pck2WKZhm737C//M48sb33JjjkcqiSb6Cht14H6ZGkVoEuSgJMPSjzn9J2ZfJTf0
0HxxX286GFRNHM70KdV4x6UqL7z3DzC1ffhZ+7diqoVVxGzZVpyeI8TTsIyPv2Nn
jeRkpQ6dmwiQQHy4SOZQmQNc1n0powu+L+jDhXPazsOdzNyxBVQ/yPcC8K0YdE+Q
BJHfLmgHVsdfo1HLylDbmCmhRkpIHfAjG97nXh8regFdpj1ydj0SnvJXk4F0QjkU
Ve49ke+sl+5wABWipZwjlqNyrMy6HSpJ5WBLjmGz9hLdWBoj6Ps/SLKrltI5L81r
wxdcKM999tDhMa6y6X5UAvpeHzxrCv6lHu8tlFsenunJgFkfArRNvQHhiDFftM1u
rJeoZsAoKvsnm85fwtK6g/J/lJ0BXBbxmdyDH/tmhfkx3qtY6zH2AIWMMzebnw1e
8wNEE1160s/4s7zNa2b6lOXsQnXKgRUxThlWsyY2YzpflRPz89lhdZeQKSVE3W+O
CVJKzCgsHu5ti1ZGrTD0+kk0Zc6jHVPGTK+GtIxuYsZh9Uv246WiL1Q4yUjH/VSn
xNAe5ip3CeyWUbfxkWnWxrJFw3OHms4RWA8iNjq876Fw7ghkzHdcPe5RXoxJG55p
s1HcUZmozc7Po+5ahBvB2y5dygjuOyjyb3232N4stVOmqLMmlyIQTndn9PmBJLwC
IvMggBYHRKGquVLQBcRNyVAqoyEkYPQjjr1JlDUkBZLBY6lt7vzWjMxqkaPEL8bi
MIhY82q+NzamXYI7Oze+Yo/XTkAMhVyJrCUoC/DKVea6TDyVRjbc4Irl/fdg+eik
gFTouDzJjEJCNo5KqGMftJKKi3/L8sT0+9nBR4tzO/KHPTZI5p+8ep5ikC4/EFZZ
Qpk4FCJ0lap8QnJxF/dV2xhyP0UTPYKX2DJd+ARGeMEIAdFjl9mCnPTH1501mqLu
PeaRdvgXsyuHykR5BHISleqhxRuCIqWQMJWMBKPgfrLcSUcyLV6KIt2DzjXPr5Z6
oUsfGLf7VmsFqdHLOITLLdjRbDIkT5CKdRSKw6OcG61qytklh2RsGmhxRZWpIWBZ
/JWzBz/9b0Qs8KdJNKYch0Z7YT/R2JUgW9gfONufwtdaNJNjrF7tczrjIviY1m+2
TDptKPJ5Uf5WIWK0hIarla07BlHVgCScdpvoiDL/nhlGZtXop6dZj2HRpv3uw3Z2
3NosBCfioDw9j2pVa2fXK4Vc+ZH4BvJxBg9BpzydCkhFJLe+AEWQSAN9fk4IDGKP
6CBfbIB5gY3EQuFDv+qEe++cYTJDH0nlcAdJTOekchjJVejTVE5yuKtqJXpC/Yv+
CFcXUted4HPqZxgBRkquG38LB1ug3JxwlX++Cf5Vy/CKYuberuXt2Q1vbsjYBzNc
3jd0GSgfVXtpS2esSLKMb/4KQoW904N9T0kgIGfU+YjHRVjBl15dB84xJ0qZpUdn
pCp9vjbba+EGQH5Ka/89k3j7iIrHoLuNn04qEpbzrjovacVCE6Uy1UEKxwnE8o4a
20xuaiosYTTS+9pYARlmwxSxh1nfnzW2MOiwwvdC8GE5zfphxI2yaw9x2bDprIDT
kxbOhuEXLckPHUv53806rW8XxgUjAavDif/CevRdc/kpzpR1imtLoH3+/T6ax1Wt
xL7qP+HTb3TX3WTl9oTri87swBqT+WTL7RpY4kGY6FFcjtFB7idliffD1XxiGCqI
hAyCin8GMd3Rcx7JfDfDWNoO9wLUwxjxLm79v6jCStnnMwrFmGtZ98xtUS4Pq4xP
KmwPfJG1EhKWpTHY9ZrSs1wNN0k8OBFc1UnKyv+S7klZQi7frfnBfLPUa7Lfsmc4
oCAMBtSfT8onQLQ9y4hbrORIHUlPqSUOtIWO7Ww6hFoHwsgznSalmeJPSRD5eozS
Mg53BG3Z4NpiUTmQxEk9kyABoILSZEvQohzTcKFEZLqk5WTjh0S+bDHI49+ELEOh
43tIQS5cOlMo5nWmykX+hupZReSFXPLGvPMY2yFWmqL4nrGvEa21FKydiUDYCGeo
Jw15te8mInQeSXHkP/B3DIzgEWFu6b6WeeAqygaejSjKfRgYwf5FN0GEDnf/zAEf
n+Zs7Mj6LPBc2BubGOfJ5XPZbLFb2bZtpmImfMlw5/wN47aMpzgyjag6BL/ejaHk
d/6dF8wiIuGMie5notJ8cHZgJ7S+mjGCRfaCTMTQsy4v2QbWAq3UouAdBdjUwKLK
/lUdVGpG6ngsp79po/d9RlQzFM+83UVW6NGQCLY/RRCOaqn9B2cwXzs7r7YTGlNu
ESVP7KsVxlZomFhETD+wmxQmCzp1y0+0OKilNNeA1tkAk5PN0vBS/N3R8iAbRDrl
UCrFr4/Y6nIJHo3JZEvjc+zeN4uj0dMIoGlddWAWlbKRJR714e9FsgGbwR8Lb3ON
1jEYFQuVBgS1Fw7VDT7mwQUhKwMtAW8iuqd06zfd0X7j2H+JFaIFd8k1slryymYb
5WSfKR/qbMF8IaHPA8tfj8xuWI+Brk4v6x88vgRgMdY0noCeQHttLx5KKMi0A9So
6FDIEexd+5czS6rM0i3sJmnqfpjLKSkFRALUls8SDHYY/XPufBZgT4Rt7iVI4kLS
FLjMaTVj9J9HykwWDG1acnKOZuXMo4XeJeidF8mseTimu6a32VBWbgatPotOUE8d
VbbkbSq6SkBrh/aGBeE4xrofy6yeTEVGXlSnHecs5Gx5ywus+rWSLCZ7un9odNKe
A5wqu0obsUOKmCyRlsCAKmGpCnG5noVbgxOdvkcpRAXM9mZosZN1tUNdTxcLHXFl
8fSl1KixTwJw+GjWXj3PBZGd9j3oUo3m9cdA+wbLikb/VvL4zbyzOMxVmRNOxTHE
hHZTTGZ9HM8c9FzrZdkyZM7v6IFT379YEKlSAtPA241L8J857MuFD18LFSFBhWUM
A90F4IlAoS159Hq2do3UDqmOb2HEBNOB+RKvSMqCP79H/D2ebpjLgT8dlpvTK9Be
AdBDl1HSOSXNKsWnPUhrOob8ncaKDG5e34QDjsmx4kLv9MXzGTzi0OgvFRDMKhwY
ObkfxcYRIANkS6OXJHLxs3GZSZOk+HU7fFgz6PLUjMcRzM6D0P0Sfw4mjbNGaVMM
E8mdmzIKXd+srFo67t8cpND2zAO8mNqUGPFSDnWx4BBClFn+djX3Xi1rCJgTFl+G
TpxcVzz014W6I5FuFPKlioI9O1Y02qBAkePXGDxqxUrQ62RmAEUlVlw6b/Oj5Zlz
eCR43UHdITQHVJeF0om/hxeg15eCwscDXhE272mtTLgnPJkO8u74NveD+fNxu3PF
+8I/9wW1pdv+Dv0FX+cclw7NLiaw1MzVepQdeI9o8ojB3WIORN6qi8ZF+haEF4wC
B68+ydgZIFm+4ZsEhxk2xBjSM9sZpNFjW88g3KtfFGe5SuvdmwYj2yZS3uXRFn6U
aSnFBOuIO/h6YVpnJtFbOxl6nvdt15BnkXHYJMn374F/LfYlajhlwReYFmCNJe/C
TMcw5oKh2l7lhrwMWf/TNmRUsG2Vxqoj1jDFXZd9vIQJjxLvMyqp1KlDewt6btOy
igG14dsS3RlpXH28AFO8pW90nt0WsNwKVvYxXOpEblPYG0MkdGCFcG9hZdXg19ab
R8eDS+4g54m0Wm72YHndyPCVr6RsoeTioFaehOdD/pt4vpw3++FLhmOlyBDG6dJx
pwLO6Z0edgiZNAOqCilMTJFr4L8PXLEBRdDe37xQsDO7Zq0K6x0Da69S6+virbyU
3710hl3Ept8uC/wwz5uKVNthjqpc1otQSJyPaymkZBtKHEl1NHH5aqN8bo4Pq2r+
2yObk/I629fZX1DLzogZDilanPBCutoC0IiEhois2RBX88wULU5PoNLm/YMZZIZW
q7kla+ygbAG9794P79NNHQQI0uy7/vsrCEgv42EF+Wxoel0gV3P2f/xdi/CPIdJt
gIX+C17VIo4NCqXdXVAWoSAG0e61T3G3HJDszJiz2zei9fTbYxFPzQwmtirfAz2B
7ksFKBfJUsLHkEOgfFggUMB0OIHPua2Rz3C3wPrNlo4SEVYXJTN980/ukw6HM38k
BHhgmnh6k0xPD/urCyhaeaMv8Ki1Nd79e5Fwf4rhFynkm4zwAooRya9LKIFqdfco
d4Sp19vbLKrHVV/2xrTlCXG0PLibKbDknT/hRGqRHJM4bTSEZF1xbW5hMilioTRj
t+Po8YTEPuPcuXUDK9iC9KZ35p/5RHJ1Sp4j2lOKwcY=
`protect END_PROTECTED
