`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5IIiQVpbznhz25wRMcOBMhLtjEwHAWgzpa0mxQBYzNR9z3RFkawXtwZMK0VHFBZ
oMmKUqJxoyJqjNAYRrCyrl2xdxXH4TRL2W/yNKAHrDalhk08gQ2UQNBN5mKhRfNg
FjYaGH76w06aefqVFmA3e5OcqyaGZlnQZRXacF4FMYosA8/J9b7UfSFbqvch33x8
7BMezxLVEAycajt0uz+6wG4iJ//lSL1AGR3beX16tJMjwJhfFmh9702+8MCbSrWT
zh3H9hbtCSUuFUF+1Tt1yfnLzBtUM1SFA+Iecri5Tg4BG6FxjqM6OSkFalJrV4XI
C+N5J+4N5LzcsyospYObyOlOM9CK4Uj4b74D+bAR/a7DkiM7isQUEvVIwTFsin9+
D/z+K+uNvHc3eOo8eXpcLfGyBIKCdaKftKgkWTP60sLoowGGFxSd2aJ/AkN9TRFk
k/Ay+tap/KBW2X9w4/1PToiRUHDPEf6yrfvKUiqNkxZCbP/0j4PNMLn9EslOSN/N
g38/U+kTJePxJjIHqNC0m/Xr727HB2t/RLn8k1Pul+GiQs0j6Y4riA6SSZ7emkSu
+vsCBR31CvBt0iQog4o+njJbV+mcdKVS916c1XjSDVSsMqS4ML7qVQRkKuePi3zo
9yRPEiaVKNac/kEZM5geHc6vfa4V4X+2YAKSUlnznwe/2ioW4hlYgOCb3FHic1kM
BNfvmVwW5cbc2jeTHBaIIQ==
`protect END_PROTECTED
