`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A7xDdByUo2qzUcZ3j5J+UD8mqboPkmny524xpfrnr1zJ/TybBt5WZSrZrU9GqKmH
6ZrAqNCwzzvcsHkNGIxH1JBUslI1t/tJQWGwr2U7t6/sH6u/cczZCbDNN66Apatu
hrouT4c8+DwOzZTC69GtWkJD1mNKOY9nTlEHRXVEBIFl7hPJH8079gJHjfYhA5re
FKoAUEAtqxtiaQ2l9y2arxsqUD4zO09cDxHpGZYxGfUmkfTnr9SGClC8Xgb5axNa
AExSiQrGlSUabu9UHXC61GAB/Cdj0qfXJkwHsF/qEIsFW7Aj4H9+/oKJviDlZgyA
QUg1stZwZ5jTLeUWztWtARhvoG0irQS/iDOUoiRTyrok7vUfCyEOikOEzxEDsT56
cAMpiM/1Akfs571AZlxaqrd+W64cc+LOKDJDnapX7TO0dNX+3RzoXu/KZ0ni3WTV
`protect END_PROTECTED
