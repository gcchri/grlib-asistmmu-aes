`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrLumzHY3jGs8s4bqL3HLoUnFU2HfquDVnQSn6iBakOkhZa0O/yW+5iC6EIf4Uyx
V5qS2rgOwFpXt9OMBWkFqHAkcOM1c8GWWu0P/rIxb9bbL1i9yjMZt29zBtG4jjIO
SUp5Gyc93GwcsGXvBE4D8aNwPfO8NLirQkDbDybkF/L3Zc81g+kb8hV61kO7vG0W
KQBXepzkhVM4pTP97/GbdGPVDxbkQvHgGgHJFTmL6te78Kzu1UFk0JDWmoGK9/W/
ZKpaCoBjfbeznzf7XSfeL5MAOVvLuC4OKIRD8/c70CmABiTwCV2Xx5/LCx+UJNoJ
BRYWNJepe+W60UV500wIwZ8yuKpEbIbsDqgrM5Ec5gnPEgOfvJdfSx9YnVQ2jwhy
u5SBHhAsTa4p6SPKDQ7KCgFupJBhmgBCvaoEycnP0oRsd3RedPo1LGAR5Y+1kBGe
sDiGSg+QGvYwL+6/w5oXpNXM5WFY21Fb6VAa/axutoIgdDQ8GH8TGQiAnRgWt3Io
V9AjhZbEGyiyZXIofRSDtv8J7gxFB6Z+1gGOx6FYnawzzfv6x8wzO5npHwIfnRJS
+Gr6EfFM/ufqa/nPUVxG4H31YOTr0DiPlt8IJuYYs9uLUmziQb9bjWXbEyEm5iP3
eg/1zg64ND0K9P/Oy00MsQ==
`protect END_PROTECTED
