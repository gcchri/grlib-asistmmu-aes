`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vaZXVUGcBEcaXxpAy2URYybLBAbrHrPC5436FqahieL0Als+cnNaUdONoLyUedMQ
aAQCZeipB/QmKI0jDcX6mgn9VGOgHOX1N3c2nHseR2uqtkXaA7CXkrh8gRRHTOMa
bVUtIMAvbKVlGcr7UHwawRWz4uZlqluf+M4CigKeFuV0K4Z7xjb++48UFHxxi4eP
0G3mlk1IJNkT7dHrB1ODfKmx3ZbabuIiggf4CGJE7WJ+ejmdHW4vYXzDZivZmntk
iaWrxf0+JbNovkbZoQGDVDJqpW/7wNz4RoYW+vSc4Is9ZvvYjoIOvmfTAkk4zh4g
qSRwolL2KfDfpJMdvFZ0Cg==
`protect END_PROTECTED
