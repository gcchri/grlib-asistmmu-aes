`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TG2wEXNaJ2vT6cwIXTrpZCsHtIEypCJ9nPvVkaOmqIFBV364AVaDVRPPeqkhgjSC
cWupvA/rePi4ncake3otKHbstDsY5G2ML3CGczPoriHW8EZCyxpGG2cER7rJaQUX
UdgtrdIGIp4imvqmyxmv4sdqmcFg7IDCuIEE/4EaCaQHAOQ4GYSkrfgsQE+P+iR9
LNugGzmccfBSoufl4JxOmm8qYiDvYfmOzx9AJabUhif4ZPF8IF40SGfw7q0fcDO9
pNCmw6b4BfRYvmJE1g3g6Hmt586drwJtd3fSSv5bzdNoXtCyg9Il4dJdZCijzJNe
m7bYqk1fmXSgAcF4nVg+8E5Lz76CCuki4/8ptF3NPS+6dVkEnmuYSShc5JC8IIAJ
`protect END_PROTECTED
