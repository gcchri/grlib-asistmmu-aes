`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zC8YG65s40jfcW9Oih2n5gbF83DGO/u1VwTIskeZ9sOleqcQSCv01JQzSmvsfAD7
dtQqiQpbWpjJ4lWnbH/MvGhoAf8dsXzGwmPQ2v6z/6TCVuWyqB+jE2jzAd67lrzj
tyZDt9gGFimNUUCWVDAF7xE2BR5KNpJXIrF+vO3QnsrIB9S7Lm1HeuwxuHKUK++f
lCcN7ur/4H3o5VpB+2GO7L3+8ayS/93oMXkwU3ptaSpmmM7LboABwbRqqLTQMEjO
o9ytyB94cDSwQbtO+Qn2R6EeYAciD5Bd3a6re4In3UAqSZQXAzJ11zgY8mu/y9Mm
T4slR8RVCLchPpOeJa/Gzt3g2qIA+41dy9/Bw2QqmVycJHHKmin3BThFyAcU3y8h
goFW6mMwIfRLOipbl6wQDfCvw5u+CjkL13ZiAcOvpmMtiuC85EPsZpk3YRpbTz/I
phiW6PqY6k+AHsGNj5NXS1JWZtDGFXVehg8fk9gKbUsL+yz74wNYMocfDOZCUBGH
DDnZxEce5MAn4WFA9d90S5IfTU/YN6BPCDA9YDO4AkHj9ZTliKvD6EUmv5w+6Mg5
wiaQEwm6XFTun9hi4cHyRkGCtfSJGlLFcFmsIc0D0b6rdUR7IKmh31ZsZaftMlP5
fZcGEQLfAOkbKQhvOCX16ZlEkeQ+JxEcDdIfEGnuUF9K3m+YRZeZn/vGRCuxcpa2
vMZpb+TyCrIARwJlDfYKCzanIkRU7S1Rh4k2e+28S3QFL0OfznY5CzroNXzrbhqn
LfGT4GY/Qs2hrCXrvXYZZA==
`protect END_PROTECTED
