`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYMC/Ae79vL8dJJ3CLzJW2BMUNbZePhRQ4NY9SG8ZtQxA65hcuWkxqu5GM+4oCUs
snB67+jQTnSGTv4zPjvspZiSAsIGP2hJG4JBjan//DTX/C/R+b7/lBDGlWiv+SX0
fqGHdrv8vUzmVII2oCHjzBCUckNVSnB3xLhxG+lJ3tJhu77QK9krkNWG+7bOUnTy
CrMOxmJ+mvmnTDkoz4bFDwf2s8GlrWDibh0Nu6y8lR1vo8VdUz39lVKjNiKDyGcI
Z6AIYxTtsxRdbR5pfi6f+oiCJGhgtH3oI08RPmmsUshjhOZOSwbiWuq0G0Ls6WHd
JyP0oHigQin/NmRWELOLKiWNOwzphc/zxAksA5p4y7cYxCbBs8CDL+7a3xuVcdxa
JaVYIMwI2CxoB1XlmpXje+tSG6xgx6lsxj7zuWpO9T+Sx6QN6bHmTFCGFl90AhyE
EFRsiU0MtQXJMGEB7EuAMSj7YBX+0d1rcQxbIkWGOpumWuvyk0lmMbKawGCTKXzb
DuUJb+Ij7BdoZJOY+Y9XMVKMDRq4si77MgjxM8xM87mOk0zluUVuZpuR0DfPWpZo
b3TVYnSd4MYMwASdCO/0KJWkcH6+5hBpQ4MAkgFZ60unLzAGdtINOYr/Qayya0NW
h2V5HebLeQzgU8YJw6Ldz13Hh3U/LK1qOGCNNsiM5drJfN1o/+Ga8ye2jLTQCj2X
K7MdFtOVuOkovBaHfavoLOFwvBC2pBmsLtHeXuMqoVbdz4LTVSqvcs6QPvENeSdU
5AHsXLdbNpq2tjUamQQkgtpMZCZ+BuU9UwS339eap9Jd6Tvtt7qE8zPQuZD58bOa
dBdT62aUbarfjb529OPWO2Rw7s1axkNCEu28JKZmDzIAUmCV0NRku7VqV0QGNx9D
ONEg3h+sDniTjfDqT7pdfIJDo4lHuRsqjLcXnbKoykl0YiPf5UlXshhySQKIYGzF
CCY2SuJkgjLKo/oMy0NGQA==
`protect END_PROTECTED
