`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ay+YCj71KX5r0w8T7gpmBZMmPZ5AvyDI75KhTUbAJUcoVqqpypT678YrhMiFEkRf
XxHUxq9kKY80VJ6jAxt2akt061nPUvTA7gVYAj7vwmGwaZrOIa/MknqeeE96l67S
apWOLP7uXA5n/sgu4hKvBQxY51DDbxMRs2f8RnnTXPluHTduHPz7dQcB/Cji9XCj
BZn/TTnY4qIy6nQHP0kew9GmXGc7y1PYMyLbUPsl+x1MQbfrRaTAmSZsr58OMgyu
ddcW+Pvrso8of2x1DBcLjsHzHu6TrbFDRN4qL6aOE3uuoK0Naf/MPnpttuBhB9Wz
`protect END_PROTECTED
