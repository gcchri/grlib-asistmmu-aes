`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEsTqb3KudX+fIuAjEuKX96Zsn1yS2DAyBFdGg7oOA41tXsp79fFbkegVw57CsZK
ez4P0hbilsNX5MBASSnlLlCJPWL0n/PqdJHLJam6qCatM/sUhq0/wOukmhsOpoJR
yVVZbA+5ru7lJsAUK4imkZTEJM75AdMlnmGKo6JtsCzniwaYTEcVv8zZWJVgF+1l
FU1FUlc6DPvP0qpfn2CRpZLCjAmCpO2sQ9EvvHwb6D0Uszx2HIezX7u9xETmsagO
oeJvkxkrGnf5CU80oAJVEReiy9rIz1mdECvU6pEg2/emKXfc6SKbLQy3Krjl2Olp
y989o0FueDJ1QhwhYu2UN/LlQbxQIrs44rzWenHKQIZACLd2hvNWx+CnuKKHH65l
PDZvRSLVxgDlXS7ZT6KS561xTFUqfSqlSBeqVrZL7IUDryB8RncYZHLSPq7BYXuP
l9xZWn86Wel+gJIrO9b9BB3ximRq24VZ9hryXTIBBBUd8ZY/tN8hilbGC9n5AmZS
WfsZQoGa3U9pw99YrKZ9VUB2yvMzhLJ0jKb94ksdxCmwdnJLA+qt1gr+KC/+xU+5
C8/aA8dIDJt0zhPGlMcA2nIel9DJAh6jzZvGaWoWopT7vWLdoC1PWwGHXCldbTY5
gMEsMlSh6nMEHUeouKIqX7doseXMKXBRCmkEuT0QsdYj2WNqrCAOw5efeJym/X4/
2jp2WTcgvRraDNz/kIG3YfJv9tD9ec6cdys/hIHuG5kAqbUIqywdMe7aTGZJ541y
nvgzwBM76gFUMbcpOkSIz5esrcSu7m8gob1l4EtgRTozY+9M9rWZaXUreBfv99L2
EZvp6GB0kCjcthbEQh4dGM+stccIJqda6infBwfy4kHQTvGVZt2Eo5vLNtYb1c5/
nq+OYooroS7/IQuJaPr4LcCqSBP0nNAsFbVOQbPmhXKWI3jXFFDX8Toeqg5PZYdy
zKYQHoBAQIYBsFSD6puLJWWERfYKg9mSuJptreubnCkwWA5BR2AhOWdlNyRFw+Mp
0uToSNTiMV5S+mWD9UH84OhUQ+wVgE0P2I3k/msRXWio8m6ixj1RSvbveHUKEkq2
uutcdXsP1Z+SeM3x+I7t/5fbPSnAUIG/7UWecxGiyAiRpNf2UqgzqvCNU6QD2lF1
kCjzF8acfKDWJzdN9pBu9o/s8ZCVXSSZoZEIUbdc3MfPllzOSOzZS4F5ZYMJrR0l
vqy6PV0a2QdU2iEOTLwSuN1/1c46+vHEnkEMzc+FA4qsXeAELhNKvzqsGFolNi96
rI2mz8bmuMgJoeCitQNiZaWcLK/apojQuOgYep0S1+yBLoGZWLqS0fN2h9FU/4Jo
t8zdMnCOVTPXW6pLq2h5BL8CriLnsygcaUSynY1uao9ssi7+gbvJ+J6YmF0iNHhx
ammTNRZoa6GEVAgOBow3qVrnCRQiRzeo9gdmUl03j8ZpeHuB2O9b+IupC6VyEAIp
i8IX4aZWeLFjd9Xzsm8DVOfKw7W9G6GpqZLbWn6PaC5g4xd2ipcwZUQXokBLR/iy
U5VUcltUZxLhkehbCSOXnZHn+JwzPwxAFrIymEOhJOnu5mUnI6SWNT8hAjnmMGbM
eb2TigJ7EzwJW2nH1DvC3icCXnnH1OWdidSuFuxxWNLR1urInYfQeflwsOFSk2g3
Gxv6x9VId4U/a9uAVeX1zcPzoXief94IwuhgT2jMUxnW3BT5tZOypcJxj/Q/5m7r
exTvPbXzuA5efR6Yc09HeCBu/AoRgxc2lUBB0k0sW6xq/Xv8POey/sYT3gnwcwzP
xRTSvf8Qg47C2RedYb+q/SA0xzQo5v7k6IIuzuGDnPQU9VUAdKeCFyqXY2R2nRt8
cjwBACwl7A6q/oiITRzavwY31ynSz33kkV8q2kZhVmRqaA3f4i9SgY5kOzJwI2d1
ccoFXhEFY7/TSkBDyECLKiNhCC5ODyDwDlKcwlj9ql/F8cTfAFHGPLy0QraZUsNr
yN0vqfAOJWcVP9sJ7nVdU/Uv80IUN05ahZ1YDXsf82Ch8V81OPxGwq+66rq4CSdl
MXUbRWrH7unFr3hReNY/bVpwZn5DPlgV5dBy/dlwG2Cma5jyJR6c4xucmM5AfxgW
VuMCUQBUY/sxzwAvP+LGzf+k07+MsIrOCPihgNFd/mSWiY2LE7FNkZ7O+zutRGqy
p2M3yVC6I2TIDWYAsi9M9tdEgU7E+LpWpg0yCBToXqVhTsj955k47GhA9P/XsFOp
Iv7kADMwra1HZOfASYrryVkfHDL5SCSpPF3v+pa8rnlpM4RselO+nJrXzUzQjZG/
fS7fAMo3iVnkqY0w3/md6WVwDomtWozHZaVOKP3RKU+/k98iyA54SfnoC2RByOrc
xahUHlzrCs8ntooJ7WDAySYSc3tfbnIsib5ZomBs1IOMJXqAzXCHrBck8QPrY2ZF
BJfXIJyUQH/6MCbl93g1EZKs0XUcI+C3PzEL2rZzsm06PZj+7+LBQ8tl7fHj6syJ
Ezn6aHDCgMY/7DmesahvZQukEKStcyFldvM6nN16TeV211bR2uRYuQKURaOKv++R
Pk41PrVOMDCy1yUN6uBxN6ZJP/llyhtpJvv4ZDCth1O2z7ReTCArmHN0Hj2sT340
HDf02nAV7eev/NlyL8yEdwfv0+l5inB6xwIz57yeocFrPAbVdIC5EpJGQyBCS0CP
68z1mYtugBy/k20UPJ5vM8PGfkLrJGPdJuXWtgRVdhWA24DEAyePZoF7kiS+mXTh
eEyYheC4RSBPv0PIUoL5cCRmspzAt3Q3gUXLopx1IoNp4eG3ZMiSzd/jVlyvc5+2
7qqznYe6C+hQAYDpIRjxlVh/hMI0Tj+IpHT/4MYLgxJuwPjl/LAqiR72lMT2mjAB
6ATmve4WO+b5mvYmZfmuEErb4rBQ+YJqn4IyhrZWgxozd+SPZ28j53GQpyzU4l2W
+tSNfC0oIBmeDbeuJ7VTGuT2t4HfKSzPr+uk3xPJ8F+BiJCutyut56cj0V+AEorA
mumEeknrO7eSVMeLUby2VDxCQDspz4xbPeNFqwlCpc2tNECYOxGa/+/5stmeHHZM
+eta5aLbNdBebm02Fc0VmM1wF8X2ZcL9/Dcs4LhvmRUtxVzqI9zzdhadSsFfGksG
nVTI5VUWvwreTXkNKJe3SY4gVor/7uiTy5WvD4sHkvN/dUf7gWKpnUZ21Y02zWZK
owxeZMb+SIhJJoDlcbQqeFJk8aZHxgUNd7YRU0H2LMax3qm2qPlrimc0p73SG+u3
4my7nRvkUWUtX64vpM1OP5wXFrXFSNWFzEtfvI6BREyVWFFG3cun7Skqrbu/v8of
S0SxonUtzCRJvusHpK1yawbj7Or0wNrIexQdAhF3KCZKdrl9USuBbjU/twpJxfrK
j3nzPVa8STXo+5O2uoS+ScWMujcu1mrpJCzT+zVaUBGoHGkAcmGJSJsrla5E4a3q
XgdgjNY+7/T1O5QR7iI+NpIOYuDi1KQSTL1/qS6hRNDf9v/uiUuPp65GNQgbg2kQ
g6Y02G2D2COK8P5Omu8zG2qi2v7k03hzEeJTzNDO6qfU2CChRNYE/r2yRv1hLKEw
HjgEIbOpdWUvcTSp4Jzl3Q+DMaqO/diKTI05zi7tGqFsPsww3o6RU2SxAgoILFV3
hg+7sTnm/SWeym5rHeOxnU2XcrplVnMp8Lt/m9BM+r4TkEwl2U/laHJDFRS2NXEk
YKCSPAGivtYKUqdf1VsUXCTTuPTVgkvS35LTUq90v9+qJyocJAtyHwE9ZAzSGx4j
UxkCpjbdkTmjL31buABJQybe/mOJ/FKIWdLm0zpkGI2BC1iq+euRXGlHmTyksY97
5Dg9xi9cikV8nNs0Amm3C7MoYdRQf+WSwF12eTGVHjkgPlOfKZLbTxny9SKBQHab
l55NNN0f9evA7UM1xDCR6Hgz8/zvVLzT03LClHDnvCBOlEQo3dAE9KouFT0xZLyA
hBTOGg0inSAJgFUxO/CsyfLV6kxCyKVIzVF967/v3X/yB6bPMnV7Xat6rvpvGe5m
`protect END_PROTECTED
