`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TS2Z+wc5YaUXdrFuPKGskMhWRhkygfnlntcv8yEmJ2xvM+TAIMCX2PvHyYD1oG5x
LfLiEIqvuGmVfiwmEPm0YuYgvX6oOu1r5ps9lK5maKjuSHP29AFJXiE/rP9df6AL
4Av5dTio3Yfe9BmxLbqRtb2iU23S1rPL3/BK6uzy5jYbxA8+fsm/JhcHQ5kjxvYA
1Ujz/HpmGSA2qxOrzbPNWr6OKZK0stPUFX3IlhQpktoAzScYPNPrkwE+DgTrRMyh
nrP7sS+49bbu66f8UCHJutHVWZDbgRtmCkLE0I49LhBqZbN5PwrWko+TZsvVowF5
GjGb7d1CVDsA0nV1OQR9eR74D6u7rF9ojYLPh5CErZv1nHcgZz838yXSPtgr6SFQ
`protect END_PROTECTED
