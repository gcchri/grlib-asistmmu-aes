`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZPlVQgMoD6DEVJ0e6KQXEeA3xm1guxNkccku45HRXeWTPHR76fW4fuP6tsc24l2
+vReszPSfBl0fURcIUmikz525rOipKjXGLMuMihDAc/Y9CJREaSE5Q9ElJC/t/rw
gNPSSGKKYpTKjsP2cGv+agofHt4LzMfVGG6sNg9KJI77RWr3nc0T2COQUWSRzHAV
oxVZqT9Jpm4o0BsPS3+TdcT+kzpQMWJlwW4HpARsnC4XL1UhwDfdVLUw8eNgbrIw
M598OCWaSOiTiHSc0BmRAcFM47yPnmURkRQieS9OwI2G+zWS+22gbPbzG1Z1SELQ
xYMJV0XOzwak1YqaakNAaBYSD03JnMvVo7bFExin4wjv59fJRM2B5exqdX4HfUS9
6oxL4Exkc31ITzuwVlUfG1eYl2nnpIRZrZgHqC3AQOqDP/0W2sOSXNm8AoHkb8x2
iOcUa3dhzZ9vqlU8/eDGj1Us05FDbk4lms+19NSBfPN+96DPOdEgw+344tLJb+4V
A3H1le0oM8MnmoZ5aM5HTQYu4aUy0KSrn/dl+I2yLoUGE9MJMC5Hfo6KrK9sKcBS
+dLrykm2OH0UNuKy1Ja53uvTdDmnjM/Gn/EZ+Zitv+f6mYnpWjNztEdUCC2/gR7W
ex43NEiY0Cp1r4UPauuPdA==
`protect END_PROTECTED
