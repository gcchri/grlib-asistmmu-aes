`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B726QUJRZreRlLkz9DIQnLjKsfLJyTuKtt4cxutdNKaQnZtJLxWT3L+KuGSPyyin
6yW/anqRPpFOH2ml//rjRwdUFC38ERmMpA2h/CQByS6uqCtL+RygQi3peGjDcmdN
QvMNh+SxY42BOs/mhSJYMMn7MYOJZnL3JEonNIODNV8Tjl2bC1A2X8kOo8Y7RjVb
FI1wO+jDjoAZ+1+PfwBgQt+JPGqidxPBWJzKxr6qAPiSEtXrg4DawQqdJg1UGvR3
5ChB3RvzixQCB/X0Ch9KEaAD8AEoZeCiTGWUsLT6A0fc/VEkGHA5kDohP67H5HaS
HYygmD+EBnBJVqboVwYv8L0l6v1ayEi59HMk7NryiUeykEVDIX/C526v2NL2w3vb
+rvVENIBVuUovs6O3OijsIWfbMhUfsq6FrzxFm9/W/+gf4NWIownCS1ehl3e92oM
G1H3OvRd9jsKSl4udwBMvOdn5yDYv7X/rO3RWL1bbqAgJpdL3lklFXbd7TiEo9KS
7PUJ9LNUfRWYykkud+r26isCwAVoXTK3bbQINU6PP2pJtt8iXlSVrzzjnNCysg6G
`protect END_PROTECTED
