`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rIiVxAK7iM+NsPETfz/ix3DhsJOIUNwABlTJyQzl/KFsTA6HEGLVoNSs0Zg8eDWn
BKrZ7xdegfOqr3FUG2ekSOdz2juQsAjwRW55OfL5oTZIaRlDlM2V7VYwIw0uYQwU
ZRyMICiSpJbc9CyPv/aj2g2doC0Y65u1qTnjIomI0GF7giZku4bA4igr210LKb4N
jLwmv4SGCaMM048NQw0agIvl+nQF6dL7W6bJRwqeVDnBPAYDKs9kUTh6JqwQJeuk
8exaoSzmlPvJwuAoZLD0LGJQIzTBHMWIHHs5HbJOWo/ZzxZcgthdMI0+rpEhP4Ua
BAYmAqvFrUd7B1v8go01DqY9KaLG4uhTsZRngZ8EazsYUw0nfCmPG1TlChx119LR
RLtXmR25KL8OJc+YQBhnPUjQ6R8ZrMAKLLUIBMI6/XLrqSqEfGV0Thl1+W6+CDfK
sBy71tri/B/8c7gIaSL3PlS6qOrJYVZHd6iqPodeKaSEz8E5M5m+8CCGQQxVeHSS
nWyMZiK/ecug5VJqWHAvpN/khWWQww9fmN0YBvx3Q9WqWJjIxQoka+77x0gyO4Z7
cQqBBVeLnKJ7Vm1SodRgO1+Y8Rknv3nIiLlC8jl769JVh1gQ+BPCHlj5lmnj2OD9
sONnEi32SaRMdwOSEIyyaqUf49+JZBgYopEQ6awR+yGUinzINQUnRvW+nU2IkBO7
crV5jNpNWnrlA3GuobhEvmnzlhp2M0ncedHn99p5qD0kvtiZBbcs5sO+x+vlLRfG
l2Et7cJFtbCU7AOkU/y2W55kM56EmBVCJIFtIVolskCdKQz/6gcqCinLvJbvWiVV
lFx3/GsUqrwYGpz38Tw0E+FWcNgnqwByxZsCxGAJ+baB8C2e22yIIB0ZsKmFfsBQ
2LrpAxk2zcasxk4LmyOXfKMvUJVKnvemL0q3AGTjYpUV1rdnrJFPHxyB/kd5bII0
YRTV1rcY4/RIu4cNzLw3ke0/C6sJiyrpnmR72KunbiKPybi/aGLgPDmex33kg9X3
73g/c2KHPLT1VM4bGP6LT3kEGil3uP7rHG0Td8corq4J7+b5hQ1OZ+6FY76Yvql7
ipHKVRc4+oF42CNwrmLfYqL0SDs7FuXjfMp68kUsvavFGxyQXsuxBS76rNXykfD3
viKNutrTrLzZsNBzWkpYrkIKlxxY45Fs5xsAuKullVo0is+vO8iloHtyHsxrr9x+
1GCjex064yGDHJPtTWO3+70S8ZUMtLNhgx9seE1+6MnHeqO0g9Y/Mdu4HN8pJYHC
Fe73UfDCrPp7QWdoSqgo8BtMHxmryDtOCgQdVPRAin/Annrx81YF+BE8to5IlwzM
VtY0bJQvtccLrBxrr7oImGc77qXsNahtFrUoF6LSAjzalTabC+2MbvL15+VgCMXd
NrHu0XogXGAwbaUej3K2Y2V5gDwcpAZQO1J9V3l7WFz4rc/SJBEVT1YMRxtoQQHY
nb9rOYaxySNQCHgZ1ndGw2KshtTTlywEjfm0NdK6xMEUBe4ep3tZHHmt7HTgjD+U
5o5qATaDJee3wJKo5hLPlexqOBckjDzDrxyNt5k+4EgyZCrhkyQLLxG4nmiEieR4
cqORh8qrl5l4WSjimN/k1t6sEgf66WaL0CwsmqttFe9YKWYqHXjgouVpKoTv0BFs
m0DPhcZUq5Iy/2oe7Pd1hLK98FKe1PuyYaOe5qEAVncrrTugcQbAC0PjdZOR2owV
f3GFjSxt/6K56ZH84rBUwKqI3qv7IXWmE3rDotBbztc85EhOxpAy8v5oRyCSlGZD
2UojDURAyD4ZvjFCr+JQmIYiqauvb+lEHF4HmrO8HNKyUd08FG2/Q52BXT5Hb71/
Pjhbb/HXf4Y/uKnJVMfr6K3cX+Ys1ByAaUsqdTKV7RvwjG/d6mY+YA13wvPs30tI
4mcGJyyTRtL3lUZXyL+CBu/YMzlzjpbLRPIO3cSfT+PV/SqDw5r1/spQ867goNc0
3Q2XnVFl2BFjYyWiAvpHxBVDpx6hfeEIDpH874aJIkeiP2UiQeJNrrWmcx/X+jwu
2JC62tuEnhhdKi35FiVCMNR/Mi7qGmWMPuWV7OXIoVj3J4Fqw2OSiw9vP598RaQi
UcpzleJu1AqoB3dkaG+9ip9ZX+zuYRsy/Yp8o+txmY9BcVkjshZ0ybqKI2T5hBSB
DkL+9pkphTP0JpwDcgfBhhKT3LLWKVG0gSr+KGbymGdprJQhRcKyvONRtEwiVK02
P6VaHxmoRGQeRAcOakI5pbHV0a0J2URs8oj/oUQQUA3vT8Jasz8iSSNLPzEdM10O
0NlPmUVC9q6zOQm/2AI4iUcNovw9+uIYzgWxArq5JIutOTgPQrAe0uCLE+JT0UM4
lupQXPNSpnuP6WPLpP1KcPl+misuLPQ9Y96dxbk/Ik5KFmtYHK+pwkUdCp1b83K/
Y7skTSDY8yzeQSwJwtd4mNqqKV4B65QRPQ4LI/mKNsMy48tCMvy5SDau4NUgNLT1
8kC5+INS/ppq4kbGMVVtXmx1Jouh6PaGNNGNran3a/AeRkmjz5nTKnpEhsEjL+wM
taeuQZ2gcdF2QGJI3bcUqwEJVrWQ8enlOoEWTaoUr/qHG9Yk/x3irx1au7oVeAkO
tFHlzmxweyVedUsI/59pPRj24RB870wv834dbuWodMLe0uRHdYp3uxSM2xKYYfJ4
ogJLBjlnroZIY2vpbz3uOVO+wCAb0OXHBtHJQs+SzjiNMaW0Lbri8IfXsbXMPrH1
JwSUbR2hxbvJxrh1OtaEJlFWoxJw58VM3b8xkIJIfqhy7F3m6ZDHbyzICTvXOmMC
RIjNYAClGr3RozEI3GF11vcroqPmQ+p8H7ijLRCZcVA2pBKnvALqUlQvACAhA/NQ
v6A4swgemcEY0XYZJjZk/wvHMwDpKGLKquLID3AjY44NQ7MOlIFC3W2TDDur8VU5
HIN1MXvUOqcCUW/C181evwUFXBdgOyG5bX0UlAze+6zsGG58oaHfbrop+Be5lYZm
htZ6urdch0QRoF2vbBqXOhnggFW+hla9rZrV3yFw9akCrhsVy3jdu6v1M5fd6Cnn
n+gzmB0evl07bZW5oReb9r/VazJeUM6j3+FtgKupfPvHkiKtHWkiNm4TiZkLYY6C
87hnOej76vyuSNtbR+OENY9Cy97MslZ4VVmO39xolzAD8B72fcV4cbU4F2AtXZVI
aRbh6E1acSVCO/CHKwFz/sjRoMsAtJhQ3oyJOEEmO+Vh/Z8egETidKj+Qic1iTHm
ixl8QNrmNQK2ZjItMyclEw+UKfF/Lxe9fyae1psp9RnerMbUYF9nw92C07wWG6UC
sdSP0BVeSRXPOSJwty+nPKgqIu/lC4TO+QJ5V//FbLD6E2DxZJ0j33TtFbFNgpCe
pnTaSEvGAbBu1ITyzQGdOX38kYtnDmRQuP99Gmp2CJQwQYw09FkWJPx/MBMZ7Fdm
Ouw9nia2AaVm3RyJPWVcXEwsSjcOcQ5A3rDxR3C/reZGS9P1JLty1MVx4pIt2M4v
FFwD9LxT2tP7sf8OO1w4Xmyqit+Ov8H0pp0o0C3Ar7kFf1npADWJrGVikZ1F1rLF
zHdizWXVxtk8J0M0XfPkWLQd87S+8cbwjmQAPIIkXUR15F4t+xS16q80Lwizuy5W
xHVkG+raZ6HrcIuX8yxeklNR7ikOLENYc0mZgjBZJu4lNHYQFkTYuP2y0ztyVOHh
QaVnDq1FZwU5HW57k0osYhuijqajAWIn/KLCsxGA1MjHqONal7LVU1ckr/TuijRc
nweu03OB2EYBufNmwpyDrzFAM0KbVAT7BOKCzwy1UW3BjprP3iJaOZQ8vBeqb+Gq
vmSdpINjAamLQVVYOFcTJS6LvyM7ere+QigjQ7aIz9HedzOhAnvqX556afg7ltNr
ZpxGf6yYkUFtvxZ7kd4xtKNOphimgcqL/Uop02qOXibA7w8Zcls49ry7zcIPiF/O
aF2uIf/TED2Bhzs0WPFc1H+M/BB9PsLJnzD4+MQpasInUWb6hcAukqGZPq3yo3sr
HPFCdMQ2zUq29K6UOgsS00FSSseMw4a8rPWCWl6gVP5pc1YrTzg55a8Vm39EBndX
zErxqOLH1lyX5uibo3rOTJscD9AygHpSEwWQOZbGmSbQcPp3ZawpEhkJicOBYBfC
qO2Ccux7sv8SqP7xdufBVvYmXwTBS0YHhhNjPo9Vg+O97n6UqzbZhCX0B+M/G3VS
uPInNk+/V11FUwNMIs7tYrddiz3nAziIYmp7QoDksfGaNrwPueK8r1Nl8xu4BOWj
iGXeiE22N8p83E+advtSVE2VB2rkHj+uVCbV7Xu+xerOd3Q4kQ82NMgvXRI/8Z0N
xf4KsWMwX/vKQEznqXVOY95hTaZ/F49JMLlN8J80ddNoGkXcOW8MpLS/d7/P9pCG
v1IeAmg2Rv5a/eL14zw2NicEISmIqgiigOI/qLZa/KBU7yk9aY3yoJdedJAqLsFg
sd+/MJArGMtC+uHB78YGOd4iVW9UcE0iMgS1kAirGVlkBWnhbjJI5troxk7nmIrL
MeRUuaaaCMFTmnLQ6vFtr2bEfQj52fe6SoLCn7TYPuEZpmTcXFyHtI1fqFGfVIUH
fr02CcYhw0cpIIKVqtgaPNwfkw9casuAE13/Hk0v4o9u6m5ZCpnAFcrB/Cv+AU1C
xRdDdFva/P0lLqH+N0ya14Y3OqSfBKHab6A6yUCKAQz4DvDIWqKUfg82RUM8dydZ
ydTkmpR99tYUxViRFB1Gu95lEtPSY0cR796pDJ+WOXVhA/m+tfmLBW0Xq/JQU82T
vlkV9K2cVGZgN8et35j10UlJswDJ0B/q/GJgohPMmEfqS8lOwdxuHOO97XMcNJ74
5qa3neoVkWSJqc6QnbzOfcaGW8IP1ZVK3ejrJHqYa2LNHB13NxtdWUsCh93W9Ghx
1LKvQ4awg9Rbnp6V5apGMWLN/MvuPml2NxfHHFynrdoxnanBe9E5aJfYGhKlTN8m
0v4kEzB/+7tkKJKudKk7r5QFzlnEGidN+WDCPpo6rgEpRSKIYZQsTVDCy3oyrjE7
wRHH1CGSsC3uYLwV9MhYZ2T5M0nHttfgoQGp785p7LJ7wFqGzI88DtVVVE94ybWG
kPTLnIvTxQnbK6TDjUHJ7fYMObXk8VeUe2rYs/ZYwQOuZpsFI+44qkuBbX6cNIHd
0p8/qfiC2Szuw16Jt1K51TLCsrd5xJaFiiG6O/V2+tvYwhdSV8DVD+D1kMiAM27P
AeJ2sF1KSGnlrxZktu4gVFq8RxUZPdh89qMsubiN/1pja9ww/n7iRslpOG68vXDO
t+BRDiUyvH3GfCj1CC1Pvyd7fnLf63drP3pSntSacIgxDtvoXDKfVEaBxiGOhUzg
ZsRnOm8dZLIT5wrEme8EoyzjdXYuUlW8n2OPHDSQEBHqwLAfAZ9APf34rb6hhV3Z
071Ws9luppJpLHLcux3azOC7+1OPf/AltdBlNaRoJ1/Dksk8p+iHmCokgtnS1zgu
vMbhD+NS8oIRA7CJxIeE4PFci5U2dJTlhTeKSLKt60yTrbmKnWoVlp8epXkZH0fo
dL9NPssrITkdct3ZicCHSXaClLCnpTMbrhEqKR0H/m9sz/LqLO8R/CebeUiCD50B
PS2ZFIshSTE4igm0fyGqa2i5SCLnQNXJAG8gNJzG8uO60zaecViwj/xWNqmu2kpC
VD14xBduS6asd83h7Hs8NSCJAmLRPqUyeoLANB3gUGONfeBTQsNMTWUOlC54mqj7
5+OPLXBK3CT5vNR3rJlUxnN8GSNJaQuuy48DAHlb19e1Kqkjk1Qj4ytApauhmIpo
3M2CKm1yrmN/ucLHzBdJ75iN7Zzeu2JhSEAW2VaBFhayIXkiND3q3FfGBJHbVnDn
BwSBE10AfHTFQKjo9VlQSgazWDvCkO1h4azJL4GAYhblguJm4x14Brt/Ci70G+qn
6P/S4Cc3PvExpXvwZjuugewyGm5HLOCPz8aWnBFLijHLPxR5GOfpcHKas9lukJF1
FMMr+Uf8kbQ64fG5kwg4HHGKkSX+nWh2fvMm5Z/Ey0sOx9/Dkwf/h/5q1G3jz9RB
Nh++cvB5a1inPTj0+jSTImBRTPfuIxnnA9VmdcfAZvFrCEELftqakZjQl4AMYruj
OXMWyjQpXdicj7K8HJ5l+VLZPE0KHk2l/aTv9qEn5PPeB42yS7GXNt+LQ7A1Cu5s
jYCf698VebKiM77MqgVsTDPMFhoMoHkue04oFdnD0dVOy/KiEAzTBizrO7sLObld
2Hn92lpSeVuaTanDQblf+4nLiOGPNdu7pl8rM1QHDyiOP2K/zvSW+GDgZ8ebbx+g
Z8o+ukXw+BbZ8mIfFdWAihPVAMl3gA79Fj8TJ3Jpa5DrAbZLT97ZdwX7dGNqcEO3
4uOunUUn718W8ecA4TVlMlcg1382wiou2bGvGZy8vTXsauS+wR81RNAUx5KrgidQ
S/LVY70Wgd8P6vADQ/qT72ROBNdJCDt6zbxRHE3xhrdwF0Xb+kDDUcvY9AgvAOMe
FTtrYowRbjefb4QGlicQ9f8JWTf/frwfjCwNsg2WoAP9lgD3ElSx0V+hFaRfSnKK
LuqQ/fqeT8JcRoLR6xJuCiEO3enGCrSZmv87aaVpZdDjIvCYYGs7emWgrScxi+ve
+CntSq5boT7oNGqo4s3lZz6AY/aI0by7XVdEu01N2n1uibq4UexutykFp+O4MBU7
fdrE6K6exM2iNPnOiFPy9P/ZIsxOzH1592KB/CwxDoTl2fZjLAdEK1ozVeTTIdN4
Mk2mLYzMLEXAwBDInWT0+9Sqi/XleOivukvCR7Lo2TvJdke24NbAE6+pOzQvIXBr
bXslXq3vWbvMt8Livdj/lDHyAXMBxdklosSvNyipK1qbq2tJw8h+hZ0XFaP9NOYY
p00ghSiD188JhMg+8KKx84iZp6J3xn/7csym2teqQeGLWI0yYzQ/a8PBwuIvF1vC
hE+T2U1VYFy89OXu7sTbl7W8c5Yoo/q4L/LCDv3wu2HeCXp4gyaC5T6jD+nXnlCM
rjKcD6A3VdCns0myYuEfl8YhEj3vc3yi3HqvM3Kvld4+yKDNmK2zSuUtc8jf6VdX
Hx08CW5YXC3WchJhQlLEfUihQRUAUC/A6bCpqGfbEmIwFBsUetCl/wcXdQvXoIB5
HUl9OiajACmvSzlkpYD3qHvV44a1AtCOjYhmN+J9nd4xWSNQRXxPZWRloCMoUqg2
nm6kKcT+QPPuwEMt5f3+Obss9B2UM+36p8C4pmMPIRAg8dE2cCaFZFkvw75KyAHR
awEBxno3OvubGTif3MLjFez6+fJDVBgtD67wsRy0m8XqmR2SK/384707z4dhreah
BHzg4KnC0Mh9AOpNZcAWzq3BOWJJdu+SHVTNBnWPf42kbcgL/eO/wWknpn0yjNp4
MayKNZQxoXTrJsgefIbLgW9IB+e0YQVjcXXbWWi9WdZiAi1/LwdWbqp5FfLd6S4B
9uVqjSvaKR0Zrqx5ZXKYzMaD0lm7QSh80LxZCJTInHsRVkX+sUriN/iB70vjlRAL
LI/kbzQrDn0bx19Eb/USVEVrd5sWNQq2GaJvVuzszynWjoRVB3+BEgjCOnJZc8A8
cx7XLBFg2elJV0b9bZDarvZwX8SOCNCmFSmwKdQ6HcsZk1RKRJbsxMZXbIgLY4FE
6iQ5lDj6HndHSJ2jUnoX6zaQpcD542QGOPScW7BVxJCFFBQrtur05gSJjmsWjlQl
9u07MnRQINiRx11hDT4Bv9DpUDPG28PFjxbwKLNy4CdrnRiNuE2b4713Lhyx0mYF
+oGplg4Jc20EmOxLRgt+5xr/R/zgxJUvZxE8WF+mPO7G85Z7Bh3a/K/98DAdbQBb
J81uYVxVl1BHVpw8fUcfZA1p9Z+G8dajR59LNUolCaZ9Q69TGnoHhyQzuDHoiSdt
aJTz7rmIjh3VzUzFFhL6sivNBL8HVezLgX86Oy+rtvZ/z3VO4ICxaj0ZyVuRSJZM
611jd53cYjRkfE6BAgOQbANRp8IgIq1bTSWcxYq/ZNhWqvdG5V/qEAVLWi8neRae
ScDjP15c/ABTlY78rDMYqfsY3WZ1kcJh1w9/bLiJtcx26btO7IDKHpGv/CWfvDdU
FbJ8ZVRsh5sxkblrtx0UNgNylh/h7E2qb+4hEPv2i3zSHTxnGgZyztvKddeZRjNQ
t9zSnFA1HnMFDJU+jA0OArjfgKwlVT2+iNq86Ep25342LpjDVjw4Wfaqx5RKPmAX
h+a/X8qeQ8wp0runy71/eQW5o3TEBFzbJWmDJZxLjcK2qgZIh0qLkn3hbIFA1Q/u
PRgI0qSG0V+KR2yzpna4ZJw5IJNBFbcTmqc9BM2kd00G67V2WYWLqcYJt0q6gCoT
iKOhnM2sG5xMnARHeAOPZbx0xL/KlaXWhqv/dINoqus6Z9JpmkUmqKnYs6L358T8
JV0pULuuCDkF/ak5+YKuMAoIvkPmmx1L6LbtOzkY1n78ZX0ZaUha2nqgs+I8Py3S
LR8gRSbr0tze2UbKjl0Qn6zhkjkty0+hridUBtvMmsHSTO9oRRiJHiRDAi4LV5CS
LVJTcPnUBK1l7Liwwh5YLi2ltRQAPQwBdILCEUyC5mNwwnfJmeKbAEW0GYlApD6p
lkMc/KSZAmrxqFwmQUWN1V1iCet0wuirLxTKugKsjqI/QgK36yOLdihMZyLsoj9N
NSCM7Kqeq1kMciVA7e3NCFCfGQDNve24tnnwpwAnpoJg5gzgYPZ+PHAP7OJsfV1r
m7iTQnQXCteHFjSVij7jtnVdw1BeUg4fFMWWCF5MEDiNlaq2oBjBj9tn1UP+XzH7
hWBtOok0zQKi++AQUWb6ePqJrjSNj5KR3IOBkJswdetkZUG3K9RRcKEHg8pWfQq6
QumC0a5n9yGCB+DqU0XS0WUKPL/rTaPFeQzkmT0asOTPzbcmomMudgjFL+DFNqAK
D2t2nUXAbL4O6wP3Aw+O/uJKg/daWaKra+MvIiI8BwUy+skAx8CE5DUVaW/dEemC
DfXYTZFVzfCSnnMWIHec+YzeyUs7t9mKkA0pykS3Ezele47M9bz28dyNeCwksbNP
TWIVLLwHAVgHegBTNXted8acyOd5K7J3qHemuhPiNBj7w0ZeevQF92V24Fb1cWaG
VUp1NNgEu7up8kPQCofIZzrs8gtS1zGJq4/tYOu5HO6q0VL/FxLvDpzARlk6QkLH
O4i7nN35sFmQVY5ghcZ/byblnEV07mTIZNefdCBLGYkSnRvTBbM1YOfdxz3NoM/U
crSQHtPrWelziGvA1tb9mxLe049EgYST4PQuXfvXXt8K7VBnN+3Tgf8NTWr6vkxb
Qd41IQjW6eCKfmz9oZ2XmlQFmvKS2TIcyyWzFBfnWtBWej/8Kz6CIoPl0fSmwC7F
0x1t+CWgU46m4XwNpQQgoDmxOjXpbRJp5IOdhqqEB7mlpMzehZ2+fZBGoDzpsDY3
eDpS6ielriDomBHcCDoCjqdQR1aJHn5rtsda9kf6n3F0TXE2uT71L2wWrrpsbG0F
Ts8i9AC8KbZdxsgBFToeX45h4Snw8GfqdzeVqaw5lfAjWl6oCid9wnc4tdQRzwA1
jrWEz1sKRXAaHETGay34hQDjAko6iOJzC8VPFAHCWUle/4dm2g6bq4/GNB8rutFI
xrLP2FOPN9BdQhRXsfgPxnZvUajl2RrP4ThSUBYPhNQ86ud7i7+Ticlu34hevTf0
X/A9C8v7otiCazApdp4xTJJwymtURI4yBrItpm139guSyDU5PPOpFoKv1JU6zZIK
KSaARHSnVn6axowyE2rrxyb+bJBtgqmETU3gFwr6Eh4mGeqEv9zdreo0nMCpbSbw
JF6OkW1BUbXDt1Av+snUAYj2M72+zEPWDDbi7YuY4+LCb5/DGzNaHi2YPhRKT2YR
D5xE6fNjTgFp2aVR2AsGRhkUmzcKYJA5XoJ0i1mlGj4ThXUJSo6R2hC0Z8Hm+ZSY
IgRETd/wlKldT5Nz/EoWp2WVcKOiZxLLzLELlAW7k/EW9Vk5dr2xcjhgZDJUZTCy
IaXIBdWqQpWx5sEp4l5MyKaqsWMJTsRfEUwPKJRwH0Z0u6FyHcitL1WM0FvldWHS
nb6H87JAT5bqxN0w5ZdN+VJm9rTHIijP90WzlN5v/RleY7AB9NISCL3+kZugaxZK
bvy7jUPkKoEqPfXIaUEGYHwyarh+rMsSpani18gQHdo1Fqnl5Zjhw3NnjCxa3g5s
5lC9yJrriqIzTjXbcXZA8mivOD96On/BnqYpZNgovDtgr5ohIesgMM2MhQAa7JZS
KA1PZddXmfOKHEBWz6SL4WlorDO4vqw33moVhgWp56RrAaYUR57i1x3GeubZqoDT
rXyZ5DjGfyHx9rZp/TEN1Jcz5eqbsq4R7Dh6+X85dzEKT0VMNxBdljcNooTZg1Ij
J01kfw+q+w5hghxWQxGA/lBRsmfUIYEm5x+Rasu7kptMbQRV2WclA6rsSXpATLdm
FXrZ3iM8ugkqr94IijeNNnXhZeNyR93iX8LtKfE5iIumdTVWmO3Zac/VlWzpuM5/
ky1RGVM6l+mrjkzI8QYd+9lsIJv1+7dUPMZJmGuep9UBWlGZZH6BbaEIcCJ9u205
5n1r6aR/ltDls6+GrhwKSkEpc9nvaYBp6zKz8/DcV19F+x5jTld1Llgo+Xlr+JH7
+19ELETSjQfIgCbvbujS9V/LRrfBJqtyrjor+FxuSe58hi+3fOZAi3hihKeh/0y0
Znv/oduRa7QPI5KoTQy3OVI4g3jhBK3eN0o66Oj/xwadVYO9ZmqaFOmfrcdWwiiV
1Kg4RwGZSXwrsU/QO9HqRuKv5/NVw8GicDBL/FhgYJ5bnUZ+ojQKFyzm/doWgJQn
Mkn0uc0AqUZD6RmxpGl9kIDaLQV6o3CttoIbcAj2IwlRNT8H+ON3okiVF1ffeMUN
ZPV9u/o7sUM8GoJSN9jBgtPQlbbWla3FJVlG5s2byKxwl0Ds6Y2O2GtL6smPBMzl
cjru1+f2SSUHhcGcqSYhGLk+ybOqChW3MF9qtIK8JCruk49SGMksnxJPgkKyIOT2
YWVThehIXSVK2w7B84oAyAZwGC+6fkTLoVOEpCCqRgEh3zQ4xUvYr+sKbj+5s80k
5n8Olv4oilt7bssXV53WLiz7oLN38EQVVzDy4D2ZkZuDmILVFcLbqHEwR1UpVqlV
iobjUdPOAUeH4YW7X/ST5c/x5RkMhZ/xzESQor74t4LQ3mxKhPz4v3QFrAjQJT3h
+oZNWTaagtj9t4votK9kcRv+xS0UIvhOEdc7En+QRrSjHdzHd7eK6C0X00AiixQg
WXMKhZHLhdMgu8hKvrAqQnYsQn12It9S285qyN/S7fVuNkx0ua09rFA8NKI/I/7Z
AjBeL0FpvQ3i98UYYb4JVG8/Hqtp+aBpDLmRI/tO19Pf4lapB9T1H7emCH2FN2x2
TJhagBm0kxbdYEH/8HpoQ2TCO7PPRBXsLMu6YKjCZfTVKlvimxbRmUoNhnhb88p0
1tOnZLlKXvSHIdIKiqh7JvwwW8DgCTV8yf2oORUdZWuywAHTyiTgFNtQFNTKPc9i
JojB6zcVP12vgm5dlS7DMAhhcS946LwtXUz4NqHRT9+BOaJ5z4i9s5e0os+yrjBs
oQyyAQX0PigY3zGmE6aaFvtgFSydKs2OIDkBzhsg66pg+K5Bvi4Y+3Y6Zvx0q0I0
lZeVnXiDI+I+Xn5Ed9j1Bh14s2msMlOUxn0IXouP2QOsSpd/Z8H7+HXREGJgttlp
JRVgIx146onOXGUUsDmWwkQYAoDDmrTVXQDFQ1OV2KAX16uNjK5ZUpzUnAqlj07m
bTuoj6rvu19CFk3+TVz3P063UXsAitIsUyQiAuZDYZQmPvOoewOrqc3f8AfjOVe+
fuQDBmkgBp3WtqFlKantePZNmT/z0S1sjfdqv7qcvGaCSqVZT5i86WiDzlxjm+as
cRbmtH5lQIklw4i5D++DT5bzRQ0dqyJhACqtt35bhPQf8cll0aVRTcyLpoXtncvE
aPboT63ASbF6QuoB+WBgz737LTwlQk2RYX0NiHyXwNN3R6zBikY82x9aeQT18YL8
M69x1OSYDuzl8QUr8v1TOTVRINCFqJSFnHCiLawo2D4Ncb4mfs49UR1G/PTckHL6
HTL81Lw/KW64RcmVwVJOOlSOH4eWV5Db8CgMMVp359H8MtMoTjrMYKmhhMhAecpO
Y61qsp0qevmz5rBlPVgD8eT8JCfkFnvB2w2AOUUV3BoVO7/KAdeM/c7PJ8sUP/Lf
K7OgCQv9m1EhKLKGepRFvgGFdItK6rSJvzG7k9cCUodbDWDIgi8UnD1cvxEzIhQA
BKzVYpJ34TV/PnxijNBfv0+13ODyIBhfKkGtPQ5DdOFpuL8k5IOG/d+JHexhH0Pu
eeTB4l9gMm6Hh5kxy+6tFp9gvRRes20b0I218QjAgnXSOpnGk+FrE1ed1siD/fvt
kW8hv3n8cQLBrMeYB16XuJTxvse1re9LZ6zlIqmzygCEIQfHXzT6eJ70aRMk1V8r
B4S1tEcvxb1BWZ6j80kfg0R7wsePLIfhAcc4IlOPctrEAEILj68TH7neGjZsa7/Q
aT9P+s2oozLC4AbJEEC4Wkkbb/iJBlD6LI+TFHs2HcoJvJYvKi2l+f2Wih4XeoM6
QiNDs7hh5EU2K/mYzboFjgTe87nUxKu7SKojoTaMlORbNIkjAnt9RwPERCOzfYos
7gqGY0nyzT/pIt/Qy3jJPidKHVnWlK34phLSSejQYFEpkOhXGb03MuBf4HQ6b++X
xMupIufSKwcOywOg0U0sKOeBAtGLuQnl3JkwRoJ/cwi8YhHwFqk7/HOohqdK94zx
dwiZfPnXtCDo8eHP+fBAy7wVjN21U13MMytX2FHk9Op/d42h9SUzsE8ZlSkk5QmS
sc30kIUjIZwAbOLWAUKBbYe6/cfrL1QC96aqO/t51pGlkRnU+7fBrRzD+/OdeNoy
KRwPvsxnlej2pZBw0CZ54miGqnTCgQ8Aw6+HE3Iq8bo6gNbWo4uNefnDYbuikVig
j35b/GLHTjVQc85P03ZI/WYhuFq9ELrP7GTn82ndXO1jz3ZUaVWoAkyWpnsDR94n
ZLKd8zesGiMWIOMm+0cFAR3KjuuHmkzvszerRc7bfgpwInZAtkt1cHB04FFIqrri
gt55mtdU5RL3wSCyMGEhMyafUAtKFvBRkdLM6Hs2cTq4vjc67i5Nf2jqQSdPDZTH
TwDT6oHhaB+xln0lkO2dOBkpfTMuXJC6dm+cf4Xzf51yg9UrAoRRCAd42tfcD4lB
nUrtZamGpX4WOFAT5WycQb7xAB0EmFy+Ix9ckuhuETsWfiJnRmnERBov2tOaD2as
S4eD+EPQl8kgwzwQqryVkAQYdlicSqc0VtUUxP0NbRLX/iJaZCWRb5gaJZYPB9Cr
uXGM6EHp/zSBY1yTvCD3TPY8A3swUYddRwIrehzCOUiDimXSVXBa6MvrqEPGn2bQ
Y8PU0G2+l4lHxGzzDoMFrGfe2D34Kr8CE/E4kX8QMBhH1che++tGANgwoYKeI+zh
1si8WTH9Flf3+VnqJOgmtwkqa5B5Y+4n10tNymngsYeFTNSfGBdKfNOIbJ2wkaZn
fqFmJdGa33nTEvO1ZzC15fBy1ujOnXdbwMV9C7vO96/81eNVbHy5j0j+0Cdwz9Tk
/Z1OVuWz2KAXT2G6Nxyk2kYCSyq6BQVu6we87sHGYe7CoH9gUlFDwugksz1EW9Ha
vW52P/6Po3iaqchK3RVjxkxXqCS7L9QWzkSlzOGe3+r65AA4n58IlSuK3omtK3oH
1a2LGmqO9W5806khLwl67rDqDktlqrcdz2ZDAqF0NQWfCdkZwsO+ya99ql+ON3IJ
pTU3SbD1ACS0+l898pD0fXfX0YpFrDjgKbfFJE/bnfCC7VL5lu5YcBbshQI9JPJB
eaxTGuYmuPdxGt2/LgXwWi8ilbiPKLyP5mGWgg7e3u6hTrE0gLpIw0RYpiFnl4Ik
K3NMCEfX3oEH0+5GNWTL15sZsM/ba5EmTT6LVLlDapHuTgwsAjc4/Uv0fzlVIqdc
LBhsJ14l95IHzg7CQzwpvqLZ53u1splKtnDeJJtkwJy2/K8kcjOdoo5xQRotr8k4
P3DgV75CT+lzquoRuWwKxo3Kf+YtE4fuNFy38xZXim/Z3Tppz/kDA+8spWe50pkR
fJoXWSf7SaoIHmQ6LgOQtBF06dWyyI+egskoUPH7gN9Y1oqQNz30jI9ScunJLhKH
R+0EdzqUVZrLhsMyHSFW/PEb3yx21qfohfyoU7Gi87sL3+CjGDWP2o5aN7KHdXzc
ldhR4gX3Zc+sJ4YmHin+fuHigpYLKwvQf+B0B2dro/zIniU+YFjRrPexO9PsAKQV
oOzAy+/VOh3/It1NkmlPm6/nDdmExPsQAW0eueYwajMh3FMN/kRiI9dsH/J5I3Nd
ddg782j0+XtwhE2Tc4ancsbeHdT6CVBMP6p58mbWEqKBGep7yJvSgCn8mh8jBB2J
ORuQPLXFt/EV8pl7u5rRhB8+AM51VDsUViXmaOpRwPBWgl/QOW+Om0wVjGxPd9GB
NgjXKSA04W8BT/pbPlD/Fga80V1T7R4klhxQGZ+yxoARKW2MPpU32ybgEnc9/Dc/
5Ijk/GyPZrAgb2O30Bk9GsOBvVxwMCYS2pkqfU1Xu6ChEVz+Ox7+SLPsrp8b/ln8
ja36MmQqb5ParlBwgrP/F+RAkGNv1JSrK2Pj6CTl26AyyHSbc+CS420Fjs6xFqPi
gl3acEqfyzUYFwiNVcXQ/fL8Mh0raHrghZ/a7RWomyW9WI0WKU83kjFKeMUfT3Ov
KcycrwkFlBiZ9eOf9B0sxbqu74PupSC1HXgkL6jSUT1hqnwockHZWsgx2g06v0ij
dNttEUxcxiqfZAxmhco7FoFH3aVtQwF4iX5G52BX5dQmBDsWGCdGrDpeGhDWUhyf
6qPVp4ZT3MdOKRSL3MEPZZhknM/yb4RBrBugi0s5S9ruk8ArFu6oXO+Y/mePi6rG
uvi+uhRZwVHo/HQw+OkvUb8WO2vRR1yiNnVNooeVqNmVTIdcIf+LvpbLFaG4+rCj
bW8FHXkFrnAAW6qPOM3UruyDvZni2L7Mt6zZtr4AKMG3Wpc5hxENlgEZ1mEybWSd
n+I0rattRF43GXt9u7rYsPVD3OMw4znmvEHkTFndGtAhqLMx6TII7oi9+6vY1J4R
h2+3iKYRWzEcgdv+Uoyluf4oB7F9leHm8wF/EI6RPQ6iHFQqVF2iSia+WrUGT0kz
fSAS0sUKnD++8hLx1OMLa2WY4s1n41GYb2H4kA8IaAT0l8Z6KhoKQN1ccczSS3PU
7TTnfHKpHGqLfVJJ2XboVbUUxpw3aKKh8+Q2G+CHcpcdmndyv4hA4ttJgXz51MHk
iPGflPdqLl5RFl7jS2jVs9LENMohyDgsgMwki5opIdvLbaK1xNPRxtWJX8rs2TgV
GjD1PiAhr1YUbD0cEWBuRBHNoRaSVpKOtj/SYXg2QJc3xi39TNPEFtAmdbqy7SZZ
GP4B9hqzz4uIB38gkSaQgf7Udk5n/1piw0kgOmgKHFW9sItyxFbs6f2QX9su4sWG
O/35el1tvVvl0stDxskHiw6ntJ0FB1KgOfH4Gd+quIkMz0BLyI8cbNEsCnhrdFb5
A49iObApc9+oFhqG336iPmp3hpkwLo7+i0o/sR9pQdM4dRR+Lk0WtTVd5vXIJOWt
Y0E94qeK3ipYb1/bR3zKoP6r/36uqB4i8d8BEKzotfItn3w8jE+Dg2PZ2S8GIsO8
G+TY6FhfmqQorLSqSRTZvDXFOPEEzHTxcSB2VaS96BQyDVWpgc9YCNT9C/czE8Mo
SL4UdJkKGZEuy96TsNquVF/KW0/Kw2G1e4VjULvoZtmWUElBI49LR9h9S9EXre0/
GH6QtwWFWk7K0Wlrzq9JMqruMXrgmIQ/R0Iw9zqL3n9oTBlSjSphGmVt1eGk4QoN
gRO5b5ETrwfUqnJmdtoS1H6QPLGmsCS/aOnbFfDyUfDkypL3CiQcETgHKu6Loxoc
jXHYzpOP7LoBuzG6ZpfXff/FzOwb7IjtMSSpyUxHrtINWerYATNciMHoeFnt+ad5
Jb09avdN9nj7wealJMFZRiQAC5fxrKm1Sd91LPwsHH4hh33WZxDD/1xJvpbzGKFo
88PG85fw5g/aSdfMMjbZr9liNFO+w9jQKzCnDn/+kaP/jsEFTQt7IgXas8g5HNYi
GXYeQ7kuN5AarzRv89G/5DBmc6MVMMAtq9dOim0tQtFN17Sk5ptVH8GGyi5dk94B
xThVGaJ5G0jXAYXQvYXGqtifsCOeAZ/V2I2+0pUW1KhEeAcFdGz0tfET9K5s3SAe
m8Nuzwh9hezgcefAF3SsGK53D24KEE8eLd0gGWsPvjOP9wPQB7sJRSiQfPW2Uemp
50WSxIJEbFwAxwBQm+NQPkvik52az5/nMRRlq9I0VoDwUF7klcaxLAK4ZqvgRVvB
4XrBP0BPkFS/8rJyFrdr4n29SLSgJQvH/NnPoVl+Pp/v6Wb/SeU4+sW3Sm3bLcXF
YKaNUiGO+tcSbTtazU+BOu9Ro6aaNpFSkoyOFknCj5wr3J3JEIoueFivdJWgUmYd
2Ln+3r5bWHh7vcVxKTLzp00TfcdU+FKY1hsBREynNMJIniNZNrNuPY8omDJLuvvn
NI3m6gd3onhBpT2e7k08CNtebC1+oPcAp+ixCJZT/S+167TY3oBBdDeC5yCHYTJd
D1yPTS5vs6H6Ly+s+XWoiElO2f/pi6OfLLaoMEFMONJNa7DpZ7zZLK20CmNTj8sV
o/pP2BDkT2nxJoHkIcrBZz2ltxXaU31gq8cBZnUO0eOhOHb1UBRiL6ywofaVF2X8
OmtMb4xg0Keh+utyvwLVvywbEcHpTj/EkJ1j5PpyxnSSmR3bTHLX7lld1FQajM51
pjke61UxjzhqWaifracCeFC/rk6GNuJhazbigV6F9eMQL6ISUlp0ms29xMlfE/Zj
/CNqMAfSZMipOMxbc7KK0yLE+y7QFbt+mfc9iie5CRl5I6genzdC0cufc8n2vBA/
G9RgXP2Vdexi5OUSD26OwtQB0fYdWyfbbnR0viE5s5tEyJfRQxWMXVzS0jSCW2EV
rtST4XwrR9azUwMaG1FwQXp/BrmncSgT3dN8QawMLygZVr7QpREs2ygaH8KaaBAV
ZW4H31lN07KUisBNPL7WJpcgrVMaKlM1HhWec+gUb6V4C3nm//YPwTPLSskVjW20
gPPI2ymk2YPC4E3O1gCA8gylU7DdpRUnG0vdNSDoKz2hfjc/GIH/UdGUV6ZWcItQ
3/OhVI6wKcCYJHaXuFHool0LwXRuuES3nEJJkrZienGhtq8/44m5NxPCyTreMiA3
tezVCSGms54yYJ/KTbJm67uAcCewy2mxxiCKMH7QQlDoLOAW6MNF3tlYKjl3kZ6G
Da/TS5vRjbiQFn2q2MhKHkfiUujv0NmoZYwUsoacLXWMDogyNobAuRsuA+A0U5CX
GOByzlOkWxDn9Nw9GuYdYGF7DC5O9RckYFz2B0WeDZn4lwBAPVLzPdw5mh/F1fEH
5HTbgZsqvNL98AHAZ3t7vRxNKJs3358/gN8Xy1W/EaNeIKkQ8z61rP9ARXzWfGta
FCpJj+oH1W1wUAuXZB1bXjk1v5TDpLYxP6DWF1u/usA3T2TuXGeR2GXrLZv6vuh2
cU2uQaeD//LTp+OXrY4dV1+Tq5KJYiBTPYzMHgQ48PiMFLwntbm/biKpft4koTqX
pTXKhFiG48BFx+7+rw3HI1qkU87dMfpgS4txpjd91H3+DF1kkAl/2EI3oEtNK9Lg
TmxeljLNU/c99V5Z6thQIKhLRIiC3Cn7sJ1WUmZwQdBkFgo6jlBmOqHi3hkC1kg/
OUFFFzRmXYIdh3J+JRJd3fOR3wt7brVbwTYG9SLifk159K77/4jEXTmiOdx6vSpM
BFvr/IZzRtmtdx5+xi2CNxoT6cMg8LZIATHwGd4gFTVyWHlpVi8HHehiLmrKcQmC
VPEQh7MPJBxKJUQLyouAcazKBLuIYn592HEl1rwWvFjx5NxT/g4yyvblwVEhKXtR
r1wB0xol1iC92Py9rd23BP/AifTON7gHFEEc9+Ffaeaz4QQaK8lPP7yVPa60ECij
RppiPP49d/9QlhnDRlWcrM98ozZcSYBcUKII4hPino9J0BGM61ilq6jDfnnn8Jx+
ZHDs9WMNRMii5LFYEBsUvlTNDwiWbzw2MuH/9kkXRPFdiJxz7Yxuh95Cyqj8Mw/I
adPvrde/gJ3M+MyEHReL0eiRnCJ/biuZlMtvd+NqlSSbgTcFlR26wetJVl2a1YmW
9S2HYHmQlTlk53Ik1Q3H293RDp1mrsJN4eN2FgP39ZG+i0OsdSgAwmjyiIxqhya2
G3h2OOUl2unpyUmO7aB2tEeE+am4CTc8xGqU9W+psTGZAfnQ3wR1geZWfewSkn/c
qYsMbfETRAZ5zSy7x7uHgl/iCGByZ1v6yD4EZH9VUGzEjllTNDQZkhoukCPhRVr0
/RiMJCPbePOWYU/A1ut8YOZiOmagA0vVvQAhLZ2qwvbYorpcb5RneW4X8M6TEojm
sOmCdj/naEwIeKmTtJH30rvhaubRo+GBXoyHgQQ0orgJWUgYMeU9ukq0dMXlWMvT
j98FEItVGP4yjesSPPRKq3pyRv11cAXzgqoOZ3R+75bAlRE2Bos4XCXyKz8ppmsE
vi6Oe6oOzUgZhR/dRYueD7rVHsuTZzSSU1SsC9OZLiDr+eTyiq+U6hWQdsF44K4S
cGQoSVasoCs+Q3OeG+Hx8hDdRpV08DLX3Cln7IDAYtisHougmwlFBtNkILLxWmPA
M9FX1U7gG9jCusMyxd+R2pM7rCHYb86sc0jd2oPzJ62VclpcSRQO+m43sy7UIbhK
FcU6si/EarqCphEB0R3E21pHi7zlcdqiWWtSt8VxoPflQjBiRRZp9K0Jh5JAL+Je
1HTF3Da6aPTwD7siD/d0XGuXgrK4T10s0y6wxzXWGT56qlczkbjx/pN0hy9MW05y
9o+5/2dcmP+JAxTV4LgqIQ743ye2PYUZ7mS4rVrbjJhwBpDsuV+cxj76It7sKnLl
xVwUEQNKa92IAaPVmbxxJgv29Ps8YFJaPQdFroMeLrlknj3NzAyX1XkwRX/fzM8w
PvnWjqtc3oIvOEDN/qgFFW7yTlJ0gQpdJYiGSvNoQJD5Zeg7K0lSpiZeUy2MQcsO
U3YQyRtgUrDK6ZdlGYxDZ5r6M/h4WSK/iu2iBdzLab4DrTBs4JcHoLLvgu6l6CNj
/h8sE3A1Lg6wDGMAFROvkED0cVc6VIO1mdQOfXHSR3EbtG1rxYj8Ztf49UKKOE0I
5htRWbiHEJeURMh8KE0SO88vwaaDYHSjSMfIpIJtcSVutpMwiALwoWzGvznFoM+/
xaVRogLWbQq540Ih8QBZa95I1tALgHT/tq+uyRBqFWm9V0PS9tnhXj/yi5X9r4Ge
xwjzMpSbCuL2+uwthHKN9WEwi8GY4uQOD8EHLlcaJx43vQzTRs2OjiIYan2Cl+02
3uaAZdrxqPcZNwUZedvaewasBNSPW9R1YE1Ze5nur6/q8+f3StzPg6FZZE03IW/Q
luCD7BOYiCDwnaeGAC2FkLqsgIwezodcQBsgRVRcgmPsHc7C1NJoNwwXM7E0ehXL
cJDkmvmNFTDhT+RXuMYd9Yyza7ipot9+4KmS4EFg8e3lFJl8WnurHGYKdD7mEkXt
zo4dY4JkmIs11DLyMltWqYbISdvT2ODOFWNlrvFsgwXdlsw0ccbRNt3XCplDDful
VTcaGA/I8kPx5kfGXEJyhJsaeztXkYL6J11eXpaITMOxFePQTRwLzSmUNpvbcyaM
jz24UWv5JhMtXaJ2ZHQ818OOKNxIxedh1tSilbZTy9rLize0DSkOH79gkdEP74Gc
c0vrJwsYCclaRbFyqo1Mty9jE5MuXj4GalPRU5BXl+CaPpM+rh3bdR0uxEcJ4xBA
oWJw1TnhLdy7ejDT2YDSk/C+ykhccMX3gp3PqAmAAvSmSCqJGJBl5+YrL3U0gwGo
gP+2BKNYlaVMQecKAuZZtY9BlYgJ5YdsfWnv13MeL/Ap0OugEL310AfHyYD0DwVJ
SBVCQ0SkegJfp/2ckSvkWfSQvdnY+t8kLoEnUvY/+e9qZNWQ5uiyWZjbHxuRHKht
VSknxvjK/KdD5IrKuNcxbBHLto2ofqQLHUr1TKNQGjKXHDpdVUTmVoSny8tXUSU/
wmcSOae7wycuo6vDwFnJB0sZEsEB0WdhaxNC1JeVTXgGDRWWZd7NHUGwawNEnn8Q
VnhhzwfzdvjjRzP1kihvd/EHcJQdCMAxn/7wBwBEPEvHE8w/tKjptWgBFzxul39K
4IX7d+niHdNk4TEyI39e0jDSaEsSq0MMi33hlTW3ylOkaPD0nvkUH2YL4UBsfU6/
R8cY7XkW7Oq9z5QWktHenIT+pBHWwLkAB15nKfWTc5MUk0TU/+dUEJ04KU4YjdNt
4kl+AzUeX2ihKZAR4xfJfk+HtPKltplIM8lRvucIDbaQfe7iuuheCprg1cJYJBIN
vWPDSJ9nQNRdlW0Iahc5EY0Btm2WjioO/aR5zIDd8zSNQ+iRVyDaNvLp+tPxIRpN
ozl1mHGrA05iD7PQfV/z0IREEnTQI0QK8/ze5xIvCYQh/CmYZPIxojj7tJkvctTV
3zVkNI7TDNEmcy6688jm3dzTtNGhHM5XefMJ992+a4IXmJaKw344pHt0SHpkYGM3
LXWZJud6C9qixNC/+M2B+nFJiOC35UMOZU5RWecMuslyT7svMpgt7NKmgCIL3g2h
68MyrevNgTfl1sKsdlvjvFRUxNEs6lrk7Ig3p4bKhJx1s4RWz6wyoGL2pSWSq4W1
uwShjPXBx6BNO6yuRzw/pVpexfGwEyvN4QROYmmSJ+M4xpRB2jn5F0vdu/fQiiZ+
TCHwMeJA5Y4QS0KUkJnTPWQ1fuBxcT+n5KGBXZqbCbLPYpLsJvKDPxFwpo3wziDy
5R2zge/LmQQ6ARMOjwyYOyq/PR1w/9HVzhbPZzpxfHqPGm8dPrEviNRWm6UOink9
VyTvvJQWyYHYCOg4MzE4UJ07geIWAAJ6xltPgSS7U+aVvmkrTj5GUfooQyjMj1xX
rOtM6DD1vtOX2XuJIzi7fvq38ASSvtVGuzx+FkUPw+hGd7As8ZQgcmR30rAOAJja
wtv8KxdBXzL0vrqZp/m51UE9SZgNSK/5vfYvC5YhnDoCn6nYrdgOniaq8ew/NT1M
UsdLBETFHb/WRkDQtXSXv93tYIk1JDrihB317Z6xK2wgSaMqbVdVsU51Xme27VDz
N7dm+Yzr6lgTSYU1Ik72i/y+r9GnivAYFrZTfx98gaNUiInOoPSsFeAWOTGX6Iyt
AoWAgGwIs6u8Uci3/fFDSzVUxVE0KdUJnMSkogYppaRXmVKyz/4DsWK8Kqo6CVMl
EuXb+N8/r3VEYscPNlIZD7erTzlkAxIbU4K0x3oCYuUzarTD8tiy1pIuYp1ZLv2E
pNGCR0gksIxqpJg33UH0WADnPLiVekp2i8NXXAs9+W9SAG/3ulnglIJjp6W9pd/j
fTtCGy/2+QZIVRWxr+R/Tsk7nMMbAW0OzjF5f1clFllvXp7VIhHfsHOwZjQ97A+4
lcI3UyQuobsROJbWunFuzRba9nWj+FoVtRLhjncqAOKJbMYxz2SSYHVTBp7U4DAO
eD7w56RWvptRmPNpbZH9AlWjy3Un4RH2FIFZqrsIDNGBVpY2BhWvCWs4/RHGcRzp
PMeRgqjiuWtzixifaJ3wxfp4RTcdZNrvB74QAwaH73m+tOvcFvFboem0fXfx0Ta5
gNh9Sb1/PmrfWHc9DDyVLUEMHQ0Kny8VY6TtDmwGn4MZQUiF9uFC73Bpy/L0ZNGi
HhiuLNFZvAfOc6URGYtnNRuei8FC2CpA3BAbdg+NPWZu6ddJqZk4Es+Lj7e24QLm
BiXntdTcZK0UyXO6G3l/VDdd/fVsDUifgSXYCC9qdJqqyoPROG1glzBR3pm3hkL1
7lMJq6llLaDqyoK3/KbUM0v7Sa6GLoWcbTihREc89U/2MiAVqJM+pfU5ktiUdSsM
RJ4cSc9uSMtdMM0jsGZXSFdX+YrIJ4k9hq8mOzZKyVsJbXQBnLqVvkD3du1NqBnm
tZHibcUroxAxeasv21JW8eJPrFu64mosyu0EbXeLLV6uJoTqsxMNmpJ5LZJ2yEaL
GjaFqLTA10GZAyOml79ESodjT37ogPCOiw/ei5m5ZiGjZI79/3u1xceuHCuNM41o
x5X5FyS+WYIED+9J4CmaOvnOX5brjbd2+I6L5gdaVjUA7XOACnlZ8OvqM2wy/AuJ
VV9jk3fekeYFQacLtf04WvmPYSfjt3+0Vih4HFXuBiqDkqJ8Q06zAJ4kSlgrnIwg
yM9UKYWmzlabmstxWk8KjTjWyxQdXh2Ula46W/GAOUiANn3fvacfNX05yYHCSlsQ
6CEGP+Zw3lHK9N+/2XTBAtjk3yIxXJyQ/g2JFr6A8QE6/z2Hv9tlL7+41NTBeEO1
lgVE/c1su84FuYxwdJblpcD0TLMc7PsmmSfd8kwC3Svy92DqrYguHbgwLg0ijSWM
zGgGfPex1Z8Z9M21d8qYwPh7/4Hl9LqRrD+ZMgshtkzJEvw6HiSvxpTbiKlACeGD
yeA+oIMaXLp6Wuh3g2OZWsa/JRTzjhAwUMJLyqSQyjeZialNXEKyqw8hZ3TKhgco
hJiITjwr2sD9d7I+30ES8tDnjj9g9Epe4I5/QprQVwb3Py4InTsd/yroQmxRU6Zv
LmtRWdcHDyk8oCOebB3RhQ79/sgrdStJqXJVubWvAy4vyAFxxrEyXteUNSMgolI5
fNGqJ2v2LLmriDavt4E4cFO59Z/xWAFbomqnZZahnHhUf9/KX7eFuCAljGDD5HX6
TFE3ZAvOzzJ1EO9rG4ALf6hk/psLixvm5P5iSCREGA+QjAhjW433OmoVSoKRtf15
xE9qvsBJ0xqFbm+/QFXZlELs5w2F7m/QB+r/sisfbpVZ0aCujuUmkE8/OqV/wCIT
PdeSV46ZGv3PYfWipvp/LPgJcbLsa0m2/8vOFbdIHrD94nJnVAcInIIDRXN3JL2s
rG4NvgEuYWoTSG4T0xNGA40D7DKONyGnUSk3N/945NWepQkaI0+d0SwAjslFWZRc
gJBu76yMpTBMnrhMXqK7Ej+UGiUq08i08/0MLY4VZdW0Gyd5G4bj0nXM2JusuhGK
bIEQ4g9WHzdZLx4KY1FQeo5PnE5VSDmLqZnJoofmKiTuqgt/IDZVTNh/6WF1Pbq8
o8Fx2W/hpX6rLwNL4zqWVASdxKijziwt10/Ymgkk+qWBbasEzZof+hWn35EJyu97
o3qPBB5FH+Z2ej7T48Zealp12cbEtVqvVkakO+5k8ntuQ2rulrXBdBmpBSm4i1f3
ZwcGtpgVul9R7zcSbzgpH3kpDSjxxyJvXO29CXBYprpoDCb4MNqXHXTvbSurYHOL
IEgAVDKzgo4fusckR0Lns39QfrvO0xk2hrrlNTNUqCS8TnMkLsu9s63BEs9lnIS0
j6U1aONGirpiga72E3nI8BXu2YN/m8kDwfuKNlmHsTkIbc6ni0EEaPXylAj5jL10
uvzeE/75G2MjPDpY7Nv8xjuuNwWWhwshYrmyZvdkf+p85ZNsFy+s7CXjZZS/LmKB
YjeXrnjaifJ0BWOyCIpQB3z2hM/v1VO8+A4i+IZdqKT9JvrDqkXh3lfXKfwtUBTv
4j47pRSg805tnsmguvX8DRSuCEmO+BvSFSyI4rEv6iu+rHJgOuFCUk2a+3dSEf6P
oAQa5JektBGimcPwqt9g7YtCXAd95NtGXpXL7mhNCSnT0Rbxg6V642vbPDuqbwLQ
W8j4Tvaalb1nA32nSa5PZclZ1/pfD+vDMNzKDSK53V+0q1wn9Pj2k7lqFXEbuuDC
fD6gb5/tn8Cx8A58nvV3Qux7XW3Qyy7UgLQ7D4VaeO0POjWvO9BawQgAJ1IyFGrY
IL8QMbJChLwV32OEIFGZbDUHDZ39RA+H+zMGKz28bQqv0K2I/PvauhrF1GaIJFur
wcMrRwaUO9HcE+iUeg4Jr8BAyi+OD+J9xWkbABzXVkrFyhhh9fAvJfnA2tJyK4db
BknjgecY8KWvjO+rpF7HCBLA1/vBXYUkJgWlbvbVSvPikYJGl4Hht9Q82vNLGubF
QJHhm9lnLfAsnoL6du11JsDxhBeDuGrv+Y7mqIEVy+1X8yuxhgAODgiuqTvn5xov
6nOmGtCGyVy+UtZFuRTqN4u9i4e36WgbceexXJLZ5HIIWWprXN1jvQsQ9T6eF7fD
lC+64uyD0MBt79zAa1bIyajLNzWo6Mi04uw+fkdacqDxRJ8niSufmQiceF6yq5wP
TrEqzBBELt7/4O8WZe9kGByWarOOchtJ/rWYtRUmog7FYGzcfd4JRuHZQzoMiPv2
983cg/x+J/vUbgSHlmsdXTWmxYmQ09RAZn4YP9Xxfy1vXXX7V6flkFm0STnmtQx9
VVOlru5qMr+iluMxVABbiZ/ssw4hvlLFIi63dIU0XLldOdBLPyENyeAYaxZ5Nbxc
S/ZQOkvaOcHQgdWaXRgOl/njx/Pwp+mXYNkVW2eABTay/99SKTLf/7/1+qkr5TfK
iwjFYx+Wt/JGHwTcmd0gI/3Po0L/SS78wmTQKtbLb4YZcBCRsB6ol3Mjqixt7tFp
j83roq9iFLkKJvqaKuI9D3syZhVhgUpCLzdRDa8hD/zCdrOMJrwknXjNAZFKo+3z
HOCOMsA+IyqZyboGZppR0F3fZss6YPbaKCz6E8bcEIRY2jEIOoIEK1Q4bodozSKM
eH2of5v3cb51x2ogtLFd8Y53nHIk/5jW9Xss1dU0K6vIbekoKmfB8PMN8v2wGE8I
sBKI0vV6C3kI1tUAn+k1IU/lyjUW1JSrXd7JGTUcmnHQT0sGBG0AiLlJqMLFDM86
bNgoRgOUQPNjchzBEE4VAdylt587BMJDh40Z9ozl8CfdPhdhY+xK8xG3DX2UOZ1R
bbVZlGHJJXMZ2MRB6vVJFUoZkqBYkgLcga8YonsGm3eO0rRV7nBs9/4JTLlIMmNK
/8973O/wOR4w+q07p5M90jpRXPxFX60x4GclquoCnaXwdz0CGyT9VlINKaDS7yUM
xHQtvcIWWcNTWFBTAgDKHdiRs8cL7UuZ7cLVfX3Kz3rx7H6hcAAbdNro8NCWKlem
G45U29Q281QhIDg5Cux9rHge+/ua2/Nkn+iwhpNuIJYVQR7thLbAcqEHVsNw5CIt
U4Zqf3UMwgbXCuvQ3k4/zJBgpfDH4FHCinyQBXHFgHbmtE51ZhYxb3VqoCOztLOe
cS/+Z5bpbWavXuliY4DQ2DSv6hR4ovQdYk7/34N/+u5B6GVeU63xAuNsRnRkMvB9
D39IyrT3i/BqB9XzHN+DN3PmDHGRbEkEea6xD1nh6rMxz9kxfve2IbtRDcqyuALr
jBAZiIPFc9CyP4mMh/RDDbkmJdsvrQmmymfHO29WwaX2im4yR5u1UcJXNGzLE4Em
PEmazBg37LfouEZ7P9lK5r9/dddY/cJM6+ORAYDwJV4oJOtAH1xEXThM5MX2fMvR
+qbyslhy5QVgJITVN/CZKQVM4u7jAuj5JM/J1s8AGQO4MwOWy84RDe7n+S/jg5MZ
58HdvPJUCSk3qKQH5q8GhukFbFgxfjogNCiB+KSQS1I0Gaz1vgmHqfxIaMGa6lbJ
v6MtV/bmB3ZkkmEUXmX40fuZOmBbAhDrBC8Z4ntl6VUyxLAolnRkmTMNO0WagcR9
PlzvRU4pTigNME0D13k3SK1TvHO8LDYTvbFfIam3YzXL3qoCtUG4bTEIA1K3iyaL
437EHNyPDOyb/IL+D9TIpxBiSPK9q6c0BvB4U7bFK4Ap9NqomNPd59wwcPOwZevb
OErbCKGPnrXZRUBK7g8USUmmzazKv5fS3IfbcCXi/Ml6Pmj34/QpEDHajt4ddKGB
/LcRu0wCnSuVwLwBJrHmobnu1DsGpMaF5MRaNYVjGmhVZz3VLLG3jyub/R/ifUXW
LWmYEqRwj78it7egd6CXKa2BTLFQOXfbBoliP7sRn2CcJz2B+xvcr66XjzthNDah
7QBm6/WFCbVBZipavIaIL10VHet8bCr3kXZH2F1xzhfGZw0jTA+mX/1BKS0Enk8Z
Nc92jTmyfLFkGotSQLlew4x5loKNHvy/W6/WX1UWtrdtF2PKDSI9aoeO7ngNmRXf
EAYcy2n0jlqjUx7ML10TSPNMe8UYJ5HQ9i2MiE9l5tlLVxs17U432t+0HZoS++FT
RtF3HH2Tm9d2V7p+aeC4aP+A5Qyp5Wkp6VjmaLGD+SsN05m04BJDKiQwuh6BA8J/
AdePq3i5OFyEfg5sr8tCi5SViSgZNPcMy/IP1dTlwkAVouEay7nJ0gRpjVlRWRvU
Mfr6jGyn/0V6BifwuR3oDCl0uqAuQhuZKw/1E6ss0QswoOMNHrf85SKbGHIj7Co7
rwEsV53lGdaaeQgaKg8KccwKDR+d/crhhAAHnTehBCf02MIyRRQ/sxqJXVQv/uXT
HjTPATl9xP6FFTflj2aRx4juITK63h6bKmaG7n5byT/XeCJnbca3nAufTJavBnBb
B3sT1wHGOToXBrw3IQWdiT7+SVvvpD42lJzeB2dbBEX7wv6huH+/qlaeJekckak/
dTRSOr40dOSvDvi+CaQV0Ig/We+O4h2kpkEyuZfhwHCzn9DAm4abmpD9Hbz7qBxf
WPsHKdqwRDTXVPDD8TJ2htzj6Qnxm+IV2hNglYlFNByWHxz9Ofkps9aWUVee7t9M
Us2Z3Nyvl/Lnm2UBuFAP7jWWMD5PeAdCSzaIqumvi/uaBMQi9Jro2rrn72nrhwxi
A9JV/6XBoXpcCV++zFRNXlWM4GVs5lpJgt04fZJ7QDLvAX5hAQOsun6zOchn/1G3
FqdNDKBEZIC2XPy0t6pkgijTAthV28igJCNywlqIEz48TCAef0teEbiuwqP3R8u4
oVEbT+RlaloSM1xqSZENI4cb8EHUIK2piVEvuGVWSrwltM6WKtAnIeS48rxbuZzH
dDbmSERZ71cmluPhpMlTX8DGYNXVhvyt/XyUrwm8fEJc14kJ+yC+kTitdCdZZkKQ
A80ZIdH5iK0olDlcvuujQ+bPNEm6Ub3obqmrNUDEwo4r9b1rXAubC9poNfyTxDpl
vZgSO+wTEltjgIas+sJkV3SmDmxs3Ta5KTymgXJYfZyC+nkUL9wYctlVEzQRtkam
YfhFEOCQCDR3aQZp80YESASFEb+tr1eJFc2jbXy74OLDZflg6C/qsaSJ1xbCw9ck
Dng+SDG1LqCsg8So1wdoAKcvyh2pXi2w5CmzdFU4rj17I7ChcSfNyV2zOLUHorxz
XsaueECYmZDoCZKzx6nNP4kivj1DwiuZAZAv9GhPWKob4hoO9m88pJQkCWzzkB9T
v+LopGNIh86YMdTHTLxUq7ZN6a+yM4dkLx0JO+2c5r1aYKgVrwHx4p7xM8HECLOk
FZTa0nIBam/TVUPMylqfhoe+/E56cGBhh7ruvaMYSkGSEAOqLh5mmOuxXWGV6bVW
mQw86TwA+NUOnzj8wsHL7Cf5evENQPZsqocoJSev2EAMsALLzMs4xZMLkdlF0Zhj
P3/BFyPg0vCUTRdYjtz5GYsuYvJM+gZIMVxXum3tBvenuWjhxfWfT59IIrnOAOdn
hG6XKsE0ywWs442z2xofpdHs2bD5pMJMtUm5AQrG+gYHy6H7+kapVWTxGFtK2AeM
1/pLPGoVFchYzEbwHXdw/RRc9L5YdtnSfXTzmBXkfdmONQubGpoou/N/RWBAxlg9
gajhQTRQIX5JPSVu15glBEpSSecv5ZWDPS6osbJKbfZaQLs3IUyqiXhMsjp3Nzca
yZ9uj/Um0LJUmihwD3BG60Ueb3bMf5MRIPvvfqiGPb4U4OaevzMJoWXmsDi9GyAe
n3Z/92N4lVMr9xzHrAOyzN97rYfgRhXLXtEONDCkzvCefpMVnujftiu+L8yEf55v
0y+QNWvYZT7d4UKuWGalJbCBdpefCstUFYYy1SRfl3pb/XjF0IueXNEoZJmPCPgC
1GZDcJfv2LPs8/opZTY9pB0ru8sMOf3yFYiMKRbo1ZrfPlro1sDCsiD3IKMfs4mf
bgop3MqxeF+EsXoi1qpZtUyEFhcs1zJWIveco4rQF1VwD8whjDVDICNc5bvVoIt/
MDHzometFdj5sX3l1PbysLD64WYgUkvivYQxTL6PUfcKf/GmNnPx38QdlfV+HbMR
g89Mqxn/B551nTRP3QIcVIfRwKf9C4GI4Hvaysdv0q6y8BD3U7R0sWlmpcpZ2+7Q
HvK7d+FvekmMx+ROil0ERhLVSouf5kOy8vc3/d8v0PP4TPVzYovpFn/Sv9IFuc37
/tIK+MeVzkSWQzTyx0mfqRo9/m/3T8ihq2kyXNbP3nYfAIJ+2iBUGB5iHjpq/ypR
ToXjhtipjXCm1cyn88Eb0dNba6yoFkCTJLXQCymmdUKljQG0uC58To836ztX/yWq
cL1TUvZn62h32Mjorv0MefX0ug773wPfBkRTKh3uxhUzid9thnIu9FkE/aCOfVuc
H5V3OiciJJgGNbvjt4iCkVHHDC0QA8//fxMF6NFn9NhnAEktvGDtgiOMBl+cG4DX
Pp3uGrNfcC584+RO9VoHxuB5kG8bPAXC6nlMXx6npItyfSK8xYVlSioC1vsc5sNV
iaFq3Z3/lRe9x/0L7e4dga3/Pf3XEKAzHvxqiR+TrUOWTENzRocU/7afDw/2lx/7
p7MQMF+XV/h79iD4dxWNLtkdTsmXnE4KZxp/J5xrggn90k5hq0gjbqs02djavZLD
48Rso9Q071HIuguAaAQk5Wm+CQwRsb89i2A1dlZgzBLunH9IB6L8GAGsMxCC4wps
CeWIzFkxLorN10KyUIQKpfn/ZgzdmUk5tLF9IZdr3eddFLgc6J+DrywkZTBQowWB
19QMmyt+H83h2R+JDBv8wyB90Rr+gEOpVVmPYNdCryKSSGpV7LpmbeXrIU7WPZOU
lBl3IBFSFcQjrNC3GVpHFStsW4jliioecSaK0tzfHB4EQjJjn3GyGRnzE2YDM9f9
XChaZ3RGhaXtTxKV+XnkpHkpBViGmsn6m3xN2NBTX8hKQLXiHCaAM+xMKw/47uNi
hY2fuXKDQyOhZHuiEuI4xVNyoKyn0Fs5QHxUReJBLu95aAFYe8Q2vihgQsRxmf7o
cz1t974pew5wngw4qFXpa3Fbax6kmUKV7NZOAA73CtgSMYk6P4Y4ekbAkjc+WmGe
N+77lEHKR4vKQdwxffR+IcbagTUi0/kuYkBW8VfyIALYComwgBv2RdRPHnPsC48e
NCiggqVnMrF56hJrgzIDdiADX7c9yr5MmP4P9U6BohP/mOquvm4TuLqav6q9TJ7c
720O7dvgM1Dpql87/GoGquAAt20gxsP8apxBQJ/jORJETSIAxteKShVLWh+G41zP
oCaYxD5f9v92WAwpBciPj3zqyfe8RWu76wxxYCWd0M07b1032uF932nPW5E0ZAxy
VrdrBT28XiX8hxiGn+6eLSq9MtonDG6f6oQLPRKmhuMYc26QA4KjYGFWvsDf/B5X
bSyV0xjpzk7ut6jChgi+fybMmEMDdqpyZBx21YKI3QZ/kn7sXaJjuBUUzgldWiOt
T1mtWmCPClK+A1NS46dhKIhqRo0cizQ5dkjuhgPfvHqiX6DEcUHVpHVClOzqWerf
uchb2W8V+2YO6PVS8ABUGgHM00Af5p/fK/VCBTU8x2ulBW7U46ncYaPb1n7Q15Su
iO+3d9vU4VotH6J/3qrvjPXD70lCQcvDohNdGtvN9lPaAVnCzKxSfwfdAxeYS7ys
mbOLkmxOKiH+rJgMEHmUrqsZDW9E/LLo1/puDYtETgzEG9/hM+pIuBDkqJe/iZma
/rwQWf39UZuBovR1cEydMQ1jYV0kEKbdtL56l+eyKdpwI/A/CRZW+DbpbPeCwGKZ
b4u6ZOlBAT1bbIHcsozfVz3PF4z8DkbQL0U9Wp5v1Ao5j0lIKSsLi2ZFp7c1tY+m
z2rs1JKRD4KG7Eble3oMzrX75zFvpAqtqIdpAkvegUvGiGqS+UOYl52w4XqRZPEA
c4+x62L4OmViGVSu/O5lj9wp9kuTPXUChniZWwg2FAmXUcS6yfHoEEU46OUqE7jv
BKx13gxyRZ7RUqgJoB8vUsCVrtsJ1UZq7k8TgPCNBYdiffhTJ33q97K0C7Eo2lyA
xzkuXjvSAlZNxvbWcWTy9C+yD3JVEreavblpLZ8L05tKk32xLKGD/0AS5LA32C4o
wDzRWWMs/CIIpdEpOGzCkGVSIoP29hRjkHvUA9izMHjVLTgiLAgwh+mQ1jLFU0hS
xJphvjNa/PEdD428Bp9XI+BVlfuEDozSWlI6c0OrKFZpOiQMsd9QU1Pln1C4hVWD
46RqcBIGvY79ERL68BSFNDgVYtn81zNWXxqRgCNSf3rs8kSqTDsN+gkJ1H/qf8q1
sfJmJzjZOLULFqVLAy+kqVQ1v+ufzH5pzcGJOVU2Vh5AJVIdRnMfmFD0reHM+eq2
8VvVzt4NDwNiuC3UtWP+2q/kPdd1Vh6OddALmPRxBeE8qvQ/+zScEorCCZsd/M9e
Wxv40ZMIUXTgW7D5ldky5qQ8KB2GhZiWnmupBj2S3aPA8Tjm3C350VtEToiOtMEk
OEM7SfeOC5fXz+jvEyfa/BvGqIMddRSZwpbK2smhPohTXU4vVKfosjWjjiSHsgUh
tZF6zB3YBhUzw/M/T6wkzQ26YaUmd1DJmLewCxuhcnp/Or4vIAl0um2ffOFZeeFj
8b+0WVJsqBXhUBscVdusnY6YFmk7GwWeHv72JZEPR94CtHYF+pjPkLU593C+YDQ3
BNMo9lxsEido71qbk+XH7oomJp2kHr3GC1GxWp4EAzMfgKlce1P5cIjFKN5SnesF
DECjgu9vKX2v4IvOfH4UX9BupdnclDs2ERqorhO0iUfr6qpW8oroEZQtmQUYI8K5
/FQPmDKqn/OiMVJibn4p+WXfRbTBtujSKCP7FtdnJwpv/dda8eZy0tC2jgA/AnHx
Cvd7tUq16rxjeonzSy7xn9MYM/ZnmkJopG5NLR3jkjdmzXvTduNfaJlNTTIHlY1G
BBjiCOF8iOaA77Es7k+04FKvO/ZLUtvhtWG6l4K1assL7MqMx7RU1xae5FIKNKuF
L2UIrOsASMVxkTyZzY74Xz5MbdC/BHXmVj235UXJiynRhjSr7Yh3XaLSQy8kZ4z8
L2YdCmdGX8G1hvauuRG5Feomzf+857E3NOiYz/ANYLv07QVJGaHxRZmmSNveJyO2
X/cDH7DOb5Rv5+iGThdxxA5MJ9kDhG0SZbt5IJX7e1XiCabQUAR18a9zrQMGFQdt
0MHMmVrx4j5mCrI7b4FSaizqq3+HW/HHdevF0mmDwi4N/jvxhGeHp77aGzzqsYcJ
22Pr/KCgBjlpmcdg6PhGIwn+Xk5+rxT4kcLaAkJnsismxcZ643Br/yOR7g6I504d
+i5/Cs+ldpcslCf7MMraVdbw2ZWTlZ+fT35LwgY3CiH3eCJX8O3VLQZiAn7pF1ff
7xlFo0/KsFJEH+SfhegfwWdMdRoMQPkUGZ5XXq8m2yc8fNWR9WEDtUOZAjWG/StP
tjr/mcLG//UzkdFtX7OOxQXaMeNaS0LVXSxqWl044EEBxiTZkOFOQXEGACQIvbzJ
2jWeWPO2W3jbbEVSd3e59rEkMgoxQlKFR4ve9RuDimM87sryJX/VCJ2t6YluWObi
CztlDg2Qsf1CySFQQOxv+cPeVul5MxoFEgcRlJNAYeCyzfQFNDdyi36Q8Z0CRjA9
wJ8pWb55dsuYipRM3+5nWIjFZtyyB+3EVvIntRyeCZnmTBCxaZ0gAhsDkp7NIVCV
kaWzH05RLUc7/VA2zQMBl5MaXG2d4ZJ07yFXrn1sJq9FFVNysXmreDQKOhXea/UM
aYbPMl3Rhl42DJGncX6lKqxeRkMSYpcVggvGGuICKwyNJagskqaQnyhJwzZ7TQHg
BFENUH6+QL6Eo8HpraHvGsbxsr6GRNt9aPqnkzYLK+6F1GGun2bDQ4I1V7uzQLTk
IUE5cMAb5xzFuFnZq4MBTxr1rb44bPqLoMIjItILXBM3b67PztEwGEP7Toi+N7CS
paRGQ8v2UdJU8jVyU8+Ea3RvScmMnV0lMlzGg1bgVofHXKBHv684NQgmG3ClWdWs
vt10bkea6jnoXvsHwWVubUj0MV9+OmSALde0uMgCbSDfpfSPP2DrBF61N58QIao3
xOGCcUBt6kUD4ASg7uGRGCoKmMAdLJgE9AdOTS34aDAN3rX6zq/pmiDppCxk/421
3nE89k1Ii4O1bahazNqzsJi5WLD8iOA+BvoiGA90w/K3OLi42pvGchGQBNTkD4Fg
rVqdplw3nT2P8fgZWhTdpiAms/+U01U7J46RtyCueq1cp54PwZUMx0yEvEF5eFRA
u5k3jtDr4PlJswffoPKU4xizcLJInnaZLc7kQsq9EGyYn+xWyR8imIwsHfobcwzK
fa7rx8h8GElOWNGRgWptSqpuN8a7db+nKzYjRXhneVOiOAi6cSQdTrPqsjI2Sszq
9pO8E2jtV7HdSZzk4z/qBncGDDaN+iKLOks/wbh70/yz3Y5lha4SGQEmi2crgxVR
8l99QYNBAqz8kj2yfYx4N9tTwaEhSzpSGR8PD/85NWV3IFNGzVI49dE8CijGNsWJ
OP8k1kgP4Pru6PIx4XkFnhjVq/LP5KYZgyBLKzuf3CXZ0j6JmmU5NJlMMbR9fS4x
3Y3y4gxzTNLn15ebDazFkysq6NnJSyY5YrI16TpZ/ke5pUq23cnoqZIt5Vnwp9xG
0eEPWuHyz/WGtYwkv8jtx4LEccEPPIAkmF5MzqA5BundsP6RR1JEeVTdUlc4wpmY
ull3xuGbp11LU0beyrZ8ByZCuBXWY5Gmmye9157lV5CuJaW6Mp7z3DqGvVK25FFE
VD1exRs2eJVLOijEwnKSH0YZC1Ea2pYBtA6vaPhicgQCezVNjOsd1dhU2q3hukFa
vhEuBWmOFeRuVLkZL8fRV1k4soZHc8iQJAkooFMDQ1jPaY8Aw/9+2Q2b9WUlv6Ej
sPs6AI/IBxhzSwsU6OMz6WTUYk4ppOEL8f2HjerTcpdV9y7iy3TUKRKlaQqj8Ko2
7BVolR+4/50g8qsYZJvCr/iD6ojCiSuhItt2Yf3TGQq0GFTbXtByewDs0JX5CCz0
vJOxuZQMMP7sziln9XNyBOkUA2kmg9T8u3NjLtq1JfbpxJ1w3TtKKtox/Sl0e8dC
c/S3VkJsj9pT89gqzXwngDNaC1zhwg7tDfx4zXIulFiuOgiFHyz/miQNEGGWPDV1
QjTOOGiw4Bxp3Q3zHFiEe1wROR9asHPNSMqIoV4ddpOL+Gba14HNKVXm3IY+3UC7
b5OOsc4DyeQhYcDbdST8R1Qmoo0zyH5GC9rwnh48k7UrHv7YoXsCPBZYTYZdterE
ecZEtYtBXne8C7/e6P63aBPQ0weMhTyO/Vba9cvnl5eZhNUVW6T3DijUAQXoSpYs
KQUT8zEQpRLRTu3ZiMlaKMyvwe2Fh6g4Zf3lNrANLKxjRuwb/89RfqbXwNY3Nqkg
0FHI0aYowc351lEqaJ2PMFgFNiG/3Gq8ylrlrNdJ6QaAiZ1G0Xie+6VHFqYU/u++
OF46FOQc9kc2/FEYa75GCtY0+IzvIvQXgAkiIGT5mn6d0U+Z90Cl/XmcvVFDy6jp
CKCncdYUrP0N7osA7fmhNlYE+CQd5og2hCwCpOAjFawkf3ng+N8EizgnBPaK+SyE
ze4g5CWlMqvkgJUcWyM14JXh19ORPcwrSUV8fOuF0X7wpfa2U031e9HjAosOxuty
WgEUujAJ6CzCAHO2gF2jcI/MK3wCCnzcFv0mcfpNW/G7Hex/hZ3jNQ2x5wqifImb
5rsrpU8rEkh8xonBZGdGXxOeeJqsQwPF32VEOIsRFhfg9kcQJgv6x+3O8+bmb2mh
Mcr4gU8ir2oNkb5SMtgp6MiaNd0+NkdCRFZRQ1Q+WwBJfuUJ2iv9Bk4P6XL7M5Vh
J3ye1gDLUTbP4BxOJLdYTI16wH2AIns4X1JeYCF2F0SdVqEK12AcJ/Irycw0KwJs
7Ul5J3/IzSxxkHKDoaqEE0Xk4UBdHyiGb4PuzbZujMdxpI+o8bZ+XXX+TeDns3mh
nMX+ydHjYhdPziJc/S5giGR5peM6IdOB6Cl1c6ZXV9HLfVuqaWNoSMpGy0B7hhNQ
1uRmqSeV6kAtCK3Misrd55ne9tE0D/X8J0c9ItWloNQi1+qV5LDImTglAueHKoHD
cbr6HDqwRcxhDBWOs0rjpillYpzjZ5vBPRqACR7ZzlnBpanudgXc719SokLsNA4R
2vKid1ys93eu0XhNOGSJ7fSHCT043iJhoAOxe8hA7c9CUXQD8SnUVtC+y2TdzhLg
cuCUbhR7Pkn/ghvSiRay7Qzz9s6Y08xE9g7gF73wF+/paD9oVhT6exXfoxlSlkNW
U2ziIgu8vVHpaH3BqHL+dhI3tSG8aA30dhMeLCosokQBQArP55PxkPU6Qu53cBwU
yHb8i4+GzsSLW5pEOvrXAdjR8j2mBMPEiO2za4zMa1RIIhQYj/XrMsS70GOZ8AXn
ViPFOsid4yEbLZ2zfXxeqArxJQ6/HCXzS+ccImMkSAVtK1idwAYB1uUVtOt0z8UB
FClvzN8AjM8OUwtqtvTn4Y5eCVKziRywjNGV2NDWZrmS9SLyKz9rBo/EtGwSvZxr
PuNovfSDGgS220z9EiZP0dIVW4wN7GJXkQB5GAS7BrRjU7RhUu8/rOBDlgX9BFGH
Sa1VUEg/e1YFlx1t+Jvxu2L5jww1xTyQ7Be7GuFegjMQp57Lw7zA2o5q+l03JtjC
/ZQTIB87hlrOXKCk0CNzgMEEG2zWYHGSC5ujubEBw+tkmpC2ZkfkuaBzY75d4NQJ
VZu+xv1mTuRY/2mBbzHaVWx4nJo1vIUbiPS14UwNVqVQy3DOLdUU3cCNvbCMbjeF
fAbYagxf9eLI6Dzqbkh+MRA6ZV6vUllc3rH87nTdLHb+1XBufZL6MLGqTvrcEI8g
s1GyJmTnLPINkq9FqiHKP9X5M8/JaOIWDS+e7A/vgecXd6zBZ3aeId64/DEa5dkt
Chcw8Pq29ANdyvsFby9nzOJqFqgeo7vL2piGt9Uh8tSrrTtrEOthaVwfvWnmV6tT
juPK8mqv16scKSpHkFbaCo31V5K7qDAhnFDD7pmaJKCfc+U5tX7ju83IZlvkuAuh
RdPQxAwumzUoBdHKKWNPsmYy/1SfSkfJcT0mDwSHMBen/4ia0y1xkE8foabxt+hB
m9NIHSK1mWiSK13T8nBpm/lSv6zHhgZDREn0gdIY61WqVpqEPU/nwEyr+nBZ+v4F
rssoYXIHIT0jOui/tLLnxkb84rRSkyPovG4aja6Ulqcx3rl7TXWH9iIY2cuCxItS
OkRjAtlq6gGFa5ENWjgC3XIdshkW/LQ6JAQshbEY3XGQE9gJqErD66Tfy/H3KEDv
FK0asPVq+XpJ5WeECsMqWTSWy9gdzGTV9GF7THbVyzVNTV3LX3qScSsVIr+Y8bxG
t+9SYPuaPOqJHzwr3Qv6Hs6FlT8YrQrEe5mq2O3bo9R5BQNCjlDF0ct6JvAffeXi
QAQCdE6DuLSj6NjFVC1MSYoLBZfuoQgdOZJgRzjiYl2txIhrYYBAJXffaY/lTJ7O
YPWE3Rr5f9alLSTvLgQ2Lvx3qElnWGq6vXhNYJqqL13R8AH9d3RWqij5C8uOgcQX
zSuPemiuhUAuvIBDEgl3uCnWWArM81UNj0k9Mdi34bXYzW3pnpTbj/UPAg0donqK
JF+/9RuJfinvXjD2jryZBQuU3+Yr78GGN2u6qtykfTVjY3/x1opKlo1NqHi0k9gr
2MyGXUZ2RWYdp1NBdvcM+ZwpHIYujWMJLCW44p4AnUJjKT6VEJxg14329+9ZfFcK
7gaKGo4l6g23uX4Gj5ecqDYcVlR+v9K7Tr7HYOTAzp7YVJbHWOilDDUFB5wigK3s
sPgrtsFHhvUzI4UhmKsjq8FmQ4PxoDN/o02VFTFTfbEQfClHY/Zu4oDpuBAFfnf6
nrm1OtjA6OWPsUV5uXRxjIoeheDIMJLbVMO5fDUOf8JoVbHYkeF4+uXryKrStNAK
EmRzRDZa0DTGJoggyIt0uo/9wtvYF9Q1GPp1bCMaXnGa8cVb40sTZhnpJ/nbwrJS
0F0PFiWYZKixs8PL2C19BdSGJ1pBnznkg+50nQPMN3zz2Ha+z5Jk1x07gCF0yiih
zipY7H51bB4W75HIxeg9gBHB8KL8XXLvQSXVP4Uuz9NDQAXDWh4Z559ps0kT/eW7
TrNPYbRBbkTeDilIWo1hh23e4myn3omvEnhKBgDHnbe2ydmxZf2b1f7r1axTp/fh
oeGJeWNxCTadekBK0RkJgqLbENUgUPJpJ9iq9656ngaK2P+GmhiJrjqjT29jZQNc
+iMDlPvvHQu3vXNyTEsa1/4g6SNzAiLd/hRzY3xyLdC9suy3EQnwI/aLZnMGUAru
q2LbwnAEgweBH85f3YwO8NhG5ylK4lccFB6ruDiQULF8md62HE3T033Y/3nXWM39
oIm+Z3TBJYPsJH03HhXd2bXN+5g1OHI/Dz/NEluOWfYSeYxaQ0g9jQq5RC07RORI
YJReQ2dpNhUp38Fm9uJLSMHXbcoFN89QpIrvkXxfYTyvVvj0x/0JN3rmScn+qswW
bNvkaWXS43vsMAM6OGkIzVoToVqzA6iHaq/23DRdkiK1Cd1e7a0qc1Yv3/a7eLHb
SF5u+IetNWFeJ13zHoVr3UEFFyBU9WPNxx4D85Cb8AOxKi6tFpUdYVueDy2w6ypD
GhDQxeFO/rzlFE+QoFm1L9ZmFv3bTJfbeEwJDsiadXhCQeHcyuo4W1ocH7Mq9OuC
/TMkq8zZlf27XjNMsKjDOlULFQnut327jWXy8Ao6acOBwH5vt+Mr41eZ+SNVzXWD
8Tsv1LnygbkF6Zjm2w7Ckdhn8jrwAedfg/vgNGcoJufBB7VHWERvVfoqTeFwoeUf
v+3gDqyZpkVfjlqCt0qnsxFnDp4cDNOKoX6rw2nhkpBsXha8lixF3Ajo/AVw3jYI
mBUBAF+U/sdnxAijAeLlfKMG+xfWugZk9uLvP+M1G5hDfFiHfVtl9mXUpxObgjUT
YvbhV5XekI8eFm84OeK4khdVSpj7+wqzwmiAJNNiQFGuyNrBUSsmmMAbo4KtOA0N
BIeTMHOLa8jcSPSxaHIzSkVB7lugyPJo/QexVTmJPi3l5FH4Kx5x+FYl2P9tm/wM
nbN+bn2wkU3I4J6tCeZ9mPeUl9zI2q2jV3mhRUpiuaL8C2W/UCaWE2Z7zmIepSsO
8z4oqClHHCCGAK7arg8anc+Mvs4/hGNV2UHx0QhT3v4ycq7rLJDafRoMQ7+nQ8tT
63qAb7aABz6ii8pQ429oMsKJKA9gl0kbm6cA2tVom3mko3vS5rOZcfaC+Sr9eEVE
BpB3eDIKjdrWZRs/H6AOrnqSVf4jJyRg/L0C9hZfQ/fyITT2UA3+r68L4F34pEcH
KgCfz5FJXwHhDDWlLBzlhePfPZIA4ClTwrLdHPCmxKqhnGLhoDOtHtNzdLjGmBoO
LBwJkS+G+bi3dzk1oOk/REM0f6U28LsDzMbHykj3aaq3MTXEWNG0tSiZha2kd3WG
XZPHl8328Ko/idYIX0D6Bz4wZuNBwMHGf0bEr9OTPlqdbHQL3TZ0cCu4UT8qgTjL
/sO5Q9Z5NLn+LVL2RkEl0grb1T+NMwjxELSvKwAwCmOR4sJjUwxMJxqwR12dRC0b
kwt9nPp2HdXHiK14Wi+/btRR6VMPl5NqFk96p7LgftplzABRaSjCEGjawqf0YBwZ
2BfyJ5PpaROybdidAk39E3lL2Yd0VzIOK1L4/aFqXStDFqw44M5tAqxTI3GPlulw
XmqhLTt4snN5GglLaxPIQdCwGd7X3gsYKu6xu3T61U7MCQfLs3n3pCNhScGDehaQ
628N8S59xoCu5mnkrVDoXFddS/ZAtVt47zwQJx5jdZ2GdAFzUs6kyxIXIylCRles
rKBG8xiyPY++nnWquNvD4t1R3BOhkebFujfCWhO/nI68Pdn3mVoigjyiyVydpKqT
I1x4uo+iSispdO56tGHnCSYct3UdJsurfVKg9bM8K8iMhQXbhPOPagu6+1aH0BNa
rtnnaILlkQDrAQgzDevLi3rUyDjFisJOTJFGCeYMo2ry72zPNOBK+becZFq3BViZ
2afgtGFsW3lys1T/CRyG7lfg7FzntWS8y7n+1dBko4W3M+JBG5zR2IfALjbkb7xZ
fqus0G1n1iunJ6RI30WyIEc6Er+Z3XoaH3WxN7IIAbou4LhiBQ0cINtvlcVQZT1f
2VN/xAK8VYsuUPw26C81uJw76blQG0ZS8il6v2HHqIGBqlfypZw0j+FxRiYNL9jf
gqEjMiAccoR2hrhKIs78+Swvg85OIEttifsirFl7zwu/JBCUw5gABiwMbhjycxSz
VoQFMbaaChh22NM+afsm8eWBI/cGJCHbjk+7a16ibJETjNqVD5xfnzqRhaKWEXq/
dL6z1bRRy8hYj8pnWZDTd5h62g58lw0oj4ToPOYfgo1b3vt+Y2eyxxdbAEcudaS8
xD8RTYy8Y3CTJXcxP71Y07c4GzcHpma7h9MjwkUCB4xLF1vX7pgFBlO8J8/0cbNs
ZnPSjrv5DtRHbjOqe1QnfA5t+S+oVIxsHFbqB3iC2KUm0nnINiZRU3nHpXt0o+FU
vaeRCol7WtoghBFurzGCzpbzET91QbYgKBTCC2LZXK3T2NliTWRvNpHrBw0A24H6
lMQQ8VlIL9kgi35a7LsihMUtE+JJyeDHaRR+jvCzvgc33Q/OC91C4rCkPllpO2DU
1Nh7OPU9ukiPOKCLU2u97y/7OoLhesLcYRJ9mvPYCoDTT2SF3y6GadgEEwptTI2u
9NPyGluj0pmtDw5MVKU41/PDyTOaKJFCadehT84DrZRyC1QqD0iv8VpMjldkrnYv
njxOp7iDero0DlBruh2pzBImUlWP9dOvURVvD+bzCkl3HG9TN9/+iRTHjojCe20l
I5WMmr10I7gTVqi+llRThY4tGuvSbNAP0wXl9So78TVyNrvlvvNwOFuqrJ3cVBaZ
bBpkGRkUY9zRhWFlXWnaLMoZwJPSKpHJyj1DUw2yAMXdm3xuPcXfrjkdL4CY22JP
wj53ejYMghbslAnuPfEhu7Wh9AsQjGKiad/Qy8vV+Csgw6RsjOqZwjgHGqqSZP5p
tXqOXePPxROZ3PkqfuV9mHsK7pI5TN+nNUSRq2vFBp6ywIeCSi5Y/cWVNCV00kdi
eOl02VTlWsUOp91UTNTMo7+uNDZJqAL8YgZRxt9gk6s61dvR9ZtA2PJqYRyUcD1w
pp47ymN4cB/Jss/3kQuq4vW5cL2Oo3mw3mTr8yyKtTueZkZZ3LNvL3R88rEYjrMk
Hgz4rX8zN69eqaFPZBt7TyH5qIzA2xO9QweYTrLwnriBG2ufI0zKXNM1ieI2+bkr
i7dtneVSIxMCL4CmKxQFCYzP4RGhgR8MJFllveNHC57DyyAba7bGHhF/K+rIs3Gn
Km9AJxMBPWeKWKyyuPEOQrv8OyWCDEo37LpWu2yfp2ZHjE+YaV2asTXoXwu3Yy78
xpAFOyCLn6saKlVTjQu4HAQ6lwPNSZNZ9zh4co/80HB1kAZcluy/PlqiwDP2oO9S
uCGYj+96moVwcyUEnUk/HCaTq1ePVUl2svuwBjl541NYFhWvCiwIBY2xUsKdTJQ7
4lXRmP3MfJlIjkqJzBUZdvBtwtxb7Zxy+Qo6jVZg+TMcs9OjCQywnpT80gp7LsAb
a5KuGgJupr45OGQTNvwECgjcO1vCxXg8AMlIgmE6XZLo1WI58rOHjMuILH4dEiIP
JLJy3vi8qA6Jvy1cFwrvcOUb8kybDOPYjD1QmsEXujx60/yjCZxy9G/dwckxNKx/
VeHIYGixjnwWIzqB+cLMEXhMU0HQu3nKG2a0W5Z+TrNMdy5Gg3yDvUkLmFPFZn35
Mds6Gby/AtxbBW51Q8aen2xpqM9KX6n8aeGjupcpiOAKgepfKyMgM3Djw38WJIP1
wGljkjNMWPRtyS1m+bkCiHQP/ShAxdKRFhCkl2qD9yeTCyEE4hoeccE90E/FLtal
HiUzBJ/8KHddbTZIKpZQVjMYRSFWocNHa8i2opWSHIDrwnGT9Nj4XHwj8T2YLaNJ
Uo07H0hR+9/AOd1cA9i6kFOn8x9S/fWRX4tBkvA0op7qM4Uw5Cx/7t7GLp6cd4T+
WS1VopFnfH06tS0qRHXm2//KOHnagPuUGWaoeLqgN7ZZLXP8tHgELAnIawWU0A/f
VdKOtmVh1vRU9jtjxodKsjM/Xy0UgUNDz93e9BrKcO5zaBsFDRu40eWn+v/5/xlp
u9BCqlH9jRk8ww8/6HYnW/s9Zprw47uJMx3uRSxKakMMrQDS8+KHYgNQzQaHdjTx
xrXd93pW54Ogz5UWas0PJp3/oSnBj+7pd9PemRw1OL9YEHQUjTjdNP3Txy7QJi2M
pniw0QwRiZoyAJAJEE6STPgsBuf3RRJykk+pY5n3uduoLArRnzv/2hH8DfO4gTsq
65JZ+FMZBdXCE4VNzKl2yKo6es1yqejRRdRTrGkFZJs6jzHhdfL5J3sqAioYGhBW
0kxUAsIU+rXIQgstk21j+NbY6UXGkfvRY0BDagXDiB+zZNgEyi030NfblePmwPyl
xgnvJ8grpJFhXx+lhIfprekJodh92PMHichZ6DaHWd0Q5x5Eve5M9l0wbySYSL00
MEb8XXd35cbwciBxD4IltK5bwrTe91L8W0qKmZ/SAcnVxUuqLElOcQwpgrmcMqeG
nOMemOuzrNtrqbN2HnrJ7MHKGplDWbMY0w+gQmDqQ5IfPs77L9aCJukTm/ieq0zm
85GvtRXgVB6ZHcLa9eYYI7XVTpkjQLP++WluQEkKkegIa5gNDZQ04mKFwk6YjAT7
CAzoHC5G6wM15uD9nnCoLo0CuqoTVbj+DAUCcGlsIzMdnfnvPKjAWqa+Q66rmgp5
wS1aNNqAhCk8L9XTjaIa4f0qzEs6dLZo83Qvx7TzxeWj9OD+ghvERJbhxKveR/QY
XEqGuWg6F/Nv+4g0GYRBItnmYJoHNYD2yDBb5M8v1bzVnky8EZ8ZSnR73HT8qSL0
Pe3rwA6k/GA4FxvkLubxkBrPjD9MwYoGuZUuE8aCfDo6zSzZC+CJSpFzolywoQP0
W7cpICaz+SqdmXzH2ocNYnTgfTU8/CMNJj0WGPFXOjvQU9UaG7/xees+5YG1JjKz
lG8drYyqAgyjMJfpQyo5AoyM+rBGIe5ieYJUK45g3FMGTykoEk8KiaxePtcP+kOF
hLZseX0AdjRzKKHTrMPK/D1wamIzq6+fwZvv1S0okVRXtaGI8aMM6lVaQOLKuekN
jRsf+2fVLyRWXvGj/6E3eAwhj/h+/KDQ6iozrETgBbEyBpAAUNBYXqD5+lpve/dO
6FoahFlTijS2U3IhJa239en97hQnlxRaJLfPKlC5MMkIbZWwcAUoSIGHbmYk+ryn
8UwQqbwdoqCV76Gc6vM05B6KuYS/9mcVBGkv2TLsDo/dsQ4FQFAahk7Dh72GyXiu
QZT6eEW8qYL9Ob5eEFnnfm1j8YDjXH0xfHxigXHCI3NeGlpVGdA6naOgurVdYOUL
NyqNceQF6nIOTCgC13Y1B0uMnBxy2enhBYzWWrePTZYokJrwZoxVVSJ5f6aivFOo
3YBUD9f+6NphXisQW9RgA5+dfy54o45ixeYvym5QcUAAlw2oACjw62B/pMWyj1kp
yWV+UgLv6UwVKbGxT8hJHOHDd6+A6BJpMMC6doyx/r5rSlFzf5KZR3HAFIJCbom3
S0h08gjFbHd++EI35JeZL1PapAnWc/eo7AYWiQ9nugng20Z2FaC6o2EN7YXOzE8d
zR1jRSUCMeUn4VtkhrvttUAaTLuFWwg+ARUGBpHCphIksLGJRsEsLrWAhkWRsLcf
72P25I+U1uet3L+LbEuwsRx2YESrRBG8jlZSa8wK1gumC3nalYjhlqdL14lIU2sh
mwSRo4sCCDuaB2I5rIpIwVFNIcLWuKNZ9dgiYqAuF+PYJjOUCZkg2seN/3e0jbBn
hlFYyrASh3totvNPLRXHxVlk/1uo8rVuCsK6wBP8qhlvNaCvwE/LmvcXG+TC4j1n
lfRnoYs0/Y1ZP8Gmo3sSYeKRpFfp+ubqQZTg5VEsIP3tzyNe1aHFF3wmVMuPC0rs
VLNXdKsVW3Wzo+mJ+Tanc+4IrP6uqYAAWZDciuJxGEKjuaJlTIQD6qBs5zAmBuhZ
WYN+tfRc544S9xTHmAAkfePA4h3PQ+utmwGQqw7retd8l+nUGAwWN5QoqNlfchNW
QV8e/Z4fpgKqjUUVyW7bJBze8Z7x8VBcVgTcp20KuywKshpRFzrtklJ2TOCfATf+
040ID2abWnFvJZFlcJHZlfeejOMs3GvTMwY5ZOf05mvw1kO5nkzO6adR0EmxHYGB
En/YzmozpdMJDLPHKmO4qv2L9iVKhfkToBo+Y7N7mHgFCx61FJHmdL4IvTckzi2b
J3F+npwPI82RhfTsiZ6R0TaXZBlvAThoN7XEMupwWVt+tL+jz2UK+t7LngLPVt0/
PS74H1ON8aflKDdY9wjkpiz+mRCi4E+pWa6HrVEksKbMHJS8soMPGk8v/MO8WIPH
wpBt1GkOxxuSLuTiLTuj/uagtS+mpWIyIJ5u1wxurNaQ8LlpmtIu0IEVZ/93j3gi
4mS0WvUJC0Crl2BEM7tDE/dwTWdCewGi0K27nRH1yrglh014A//DbxU2jcGk6siQ
Em7PPn3Fo6qgSKjbGMRXTDXsSSRQwq9HEzSJ+TcBMKnFE14Sug2PG3vv9BCUjXug
Tx50mixeBG/UUw3yGtLa42hQ16X+810QFbJcAmfxa3LPWUvwLoxUx2Ce8oYkhhBM
CzrSv2oD8783yhO30lxTa+9umGaGVKKAQk8bRSXKqex3RX8uVDhHB9zsarzZVsc0
je6A5ADajWgmX1U6mX9MZ95nBsRFJP39Pc72khDZ6ewwvylSka3jcgwLozEdJ+6z
kp09zpC46oNOKtxepfDda1RmN9vBulEUrUEkrj33bOINvZRi6MH1vjIWDWnV+Hbg
NRCtoIlWQO0PHp1Y4YZSZkCN+rHWLpYs/OuINzmD0s0X9nunB1UDYs5Tf+nciowo
eqk9R+iPIAolNqWhN5T1//9+X+UPkfpgyhR4zHHzWQvSx8tZC4M153WONGozPQUz
cTVZeuXjkMRfTkSL9eBmyqlopA7Y1bvcBJqYcl3H/72ZlTTIu3BQm6MLIT58GD99
8xvvlokv+bQssqjTSRDA37NJ6ZXoqXgaDgv7QudPsBcYIg+ou1bSVZdWn9I/qYn8
6GsUUTJpG5CmMIqdcKW7Nt46U6LSKRsd6y27y64qN11EVaf+RMVZtaZAFfYJpQK6
CoEWzVqBNX5SKndy4PdmqcgqzkI54g9sNxTP7ZG02u3JyqiQ5mv/hYcHdXDiqejy
FGGdMNUf5TaAwSdK8tU9xxilPXTbKHiurkQRwlrHgKDvs2HroftKhuiT7Az8loBA
SY5HJDzbZE6iFAgnWZ/arj8Ht32qq1lBwIhjuLyzyKGssfqdihDHN4KhhfLDU4zp
+lIxwIxe0TsKUOvApA9E022Jhw9R4Sv1c7Y9e6zxMB2PzCRzAF//lCjHHn9h0T+p
IdhDL3rqmTJ4j7oix3Nlcwnb7MyLR9rzQo+VMyQPCcEYiIhHvrne8M/RQW/zVpFV
xZpFJviBf44OzL/MIY8c1C92uA+ACsqy2BdCqWDXWYVZNEemXnbUJE8gywXpOAT5
hm0FJIifo3GrKqpoKPzL79aKU2BZQc3+kUC2I2ohQ041mWBkj/ACvTxheHkPHS2w
9DgX46oCkBU9W7NP7CXdFFPlUVpWvl3xFkOsKQh+PsHsDvf8i2jxpcWp51oJ4I8l
BAwMdk+VaV9xgOuWnUoy2Oz4Zthz0BI3+fprzufQo1mfOzy4EDZTEZs8vvIZb9Ig
a1TIoCa7lz1rmXi+IBkvMxeZbjOk4T9fVK9xo9527ZqtIMgN8baahQfHWBU2AqSE
QVkdDQjcmlbr4pQ7sTA02O8Dnsj7pIJb4ectk696MC/Xsr7d8KFHMKpRj9NzPzsD
QQmkhjqVhb4lZDimiZHMon8gkHOMu6iSSesNk6tnxHSsSVjZxmm2TRxO3XqsV+CR
PzRy6mNIq9zHlsFfxfkga1FcNOXo/bRTaK8gcFanAMaZUrIqMvtHjbkkM+pziMpH
AKM4kfYMqR//Z5KW1BSPtnJSbHidGFJNX918uCTjFY5I1rrTwh3GWiibpsXw/VNl
Caqa0rUN7t7TnUFbiqUkR2q47F3cGHjvLqIsovG8gNAq2Gke1KhEf+2Gg2lNCa4l
sA0WHQ/8b7JXgsL8XqQtPOxLbSPSnwxdcyGFwxphrCUtf6wHpHzrWJW9Mjg2e0Wd
JicYjAQerT0AkJNbYnBunwd5zxxKwbgH3cuNJbZz0ZscgDFN5IAuJFuISZLEshkF
L7qK5ct8T7hrhc/oSw+SWqoxMtpO10ZjPJPRwkZV0wmQ/tKzUmO8lr+lwveSdOTd
id3GVrthmR7iApAjkbGC6iXV+Nt5Bfc5CgmGDx01HkpGYY90FCdSx4Me2MlhYBap
u0V+U2p+MR0tC/LtCjas4t/IOtoGlHixCbbW3TWCL9XtS/y7ByibVnQ73PWh48eE
ejhikCcUvZ239U+K0qrFxdRTwuiH+O/pt8A4T8WUUlsbB8+SeiLwQXocqgW8TFxt
lZuT2YXKaXozTL8Tkxm6Bb7pbNGoyqvJqHD5AqyDXA4QjKQjEsDWjwZ0giuD//zR
pbp4ewRW/aiL3+cW0VcBulMp674CpFeOlGbmNa9VQMrtHAmMtgorql3Xay9SjYH9
eteYkWhKWM4eTv2O2VmZmLZQNBGTIz2R9AfhuKxvJ1UVhbZenyRbQyfxOroNSiDu
IKk91Bh46+MYtmi/Rsn79oECpOQ3L5esZvwVKq9WdMvlBSpPb5gqyN+2ikS3vhH+
XT7P7rIBXgb07WlntEDpCVkBIrhtKZ73rsHTgEfL+u9B1F2ZWq63/iQ0RFpvYVP2
f9IuAaDoVxSjKMzGQWxnxvhhcNWeZfk4E4Ap3Ls3MfcgNJ0NqbdyzYlOgfGWyYKU
vMzmP2sYym1iYjCig5d7pNOXOaqU1Z45h2NH4oI9yZvyPpr/CLYJlMNf9J9Mpwk1
B5/k5/0sACzPHym4V2Ir+U9aK9olfYJlZhr52v9ZNc+wvNioPWmrNxfoD7wFF8sn
mB2jYZU63/FAplf8neln4lz6ini/XxjaFzbByZvym9IOCLC+kzKOU9kRSvYWp1vS
embGEiXoK3vQ/RNx6CcKawlwLc2+7TYDhFj0u+ruFayyrYMlrBISg4yxqvQuTaD7
zvBh45HULNuyWunqscVRvvk6CpZQr8hyKIDe9JzC1q4vqDvDGwx7pXXI2Sj4+5rP
gk+WQQv9FJi4uC44SWdbN394KOX6zAZP3KmoSk6wOgqRAToaK7OH2Pzpvb0H7i4k
6EiAzmUWdlbQtnj948tpqiYhQHfsANkSsnE3wXnj4/48X2McPZAcTU++h1Klny6x
ekaRpK1L26avK+/vSTuhR00WSWnPKzHpxPAdbl5agl0w+6+XhWXsJZHxbELNUozo
TMudTzrgk0ZRI1mZNtukWGEww/65QmLZY4LmoSAL1hv4U7YEn5B8PIrc8qwXFwDT
vRDsu144Vp0MBXddOxeBb2LHmp3DTgcwZHgjzdIjnWYcpVrYeGit2mIkc2dxLvGT
Lud7cM8M+KP2jTiw3ypagtlUPyBx/NtImEZqoTPWGz4c9YK/8G3veX/ChE8hOht3
qkVg6+2zEkZjAbXOcHhjerg2GNOtjOILTMnoGuhi8IRTUGBDRK6xwYV+0fEyOJDq
hMtpRwuxtlKu7Fhh8xS3e3X9tADv4viQwQlCILoWsJEsknmPPNUx/p5yy6M4jHWR
P34EJ352uKgfeC2fH5TQuR8uBe6xPJH0thVawdvT1Ph52UCtYo5TDlkSL8uPEgPz
Fg9FmHezmtKu3FQSesImcA2To+3qL+tIYNPG600YTwricz+2ezMr1coILfOm79tX
q5vriqK1YMozZf7UmjpO9J1QwPUm9IawCw/0MtsTMad5BemYCCYWbZKTNIwAgPFE
R0YexPJE2ooZAb3/j74/8qmfFpfysd4uOkSSGACWi7uLjOOyy6tuXfLFdDI5M1DG
5xYfYxjf/QtKaV0JfA1xSINoAFzH3rp6InTqdKTimsoXzTIZOIf9A2N+dx1QvS9Z
Y8d+srUWnkFkdveAgWITVhyhHj1WYQ/ILRv03aYBwkmAo7pNVO/glQrOXZxnq0Na
wDTbgx2E3nUGwML703Urg3fF418IFAxLPNz5gOtg6iJ6Yun1zwMdVkBWFBWl6T1U
wSnDCK8pcHtrpd0kfb6IcAPUFq6Ms6a9YUZ8fbO2Qxl2SZxN2ABj+gJjZGS8Kg/C
UtydV1cxXHLdFUtQyW+Wt8I7UbsvFpvUJW98ucaxZ+EQ6n5ZfWoRwvkyYyw8zy10
UQ8tPPe+nlU9DMVSz2o173K9fWkigH4HUG58Dw1Ej5vvEJpaFfNHatmgJbsCDXfA
uaG1Q6V7TNNCyzDQRp6Twktv6QOSk0CZ6woQFLKbBDG5T2s1rxpZmOQHa8YjE/W7
pOLNwu0mJioxDrEglUKpYbiNn4uiXqEHrh/vYntj+WPgkXBqqrtzQLYG/yHD0RYk
Qy/nNCk81FdqTBIDi8hDiIulumOTQetRKmCtME+nVFuyTSm0GgpcpFLRL0Q4sRjb
z+jBj4qMaZsw89g5ewF3YYcII+jCkL2UqpNinURVA3v+SGvu+4PElkVYT7pK46ws
arMAQ+Eg5DgXKvnOmV/TpS/Rz4RLQDY7bTQ75Wv/Z7oQs7qwzMQ/MgzXcaEpiIjn
1S8QJIS8wW2YM+OQ3u5UnF8ForshQbLloJHU0ObcitfzCUy+nKYeRskNbRPJOLED
lFDeBQhwLyUIeUS+JdGjcWtkHWeqfsrBVL+woG81cwhV67euOqW8fZC3CSRzN+1H
2HA0BsvtvbyzycJtMj2Yl1BHEPjulkLY+Z+qP0hsTOgzhyQXkKnvitZECryc+Ek4
h59BnBG5L2J2sjxcFNtLyd17cBDu/EP1N3DjTC2xa//SbtGa4neATDcVGVFbtZUJ
lhW0LhV3jyMxqc2fjo9KTKW8NEaNU9kCpTX5nGWWilbXq1gRVRtU8+bAwVAT7nv3
gLTIf2W4HXtQ8u7qPZTedstCGojwAToHtDPSch6zCiS14w5RQa3VwbthmjgR4J6O
LB2VIsqtXL/b6sx/IGSgLI2PTSUY33i/uelkKcMGniV8UHRMw+FCSn3E2YCjRuat
d0+Z6xvOBylTxdu80onG+isQboiuPcoLT4ytD2qraMuRozfhJYepYWPwIqEAkbeF
qmFNz0IVN/rdawQUG/WBdaR5lkEYV8HJGt4kPNaNkdo/BHtdTVTrpd6wXzylTMY6
K24GSr7xN763vMN0OAltECDF7SuAwPER+XGu0p7SCwDAI1/ZBiByKAAKupB/0mfX
iOM7514sn/dYB8Qj6oepTyBv5ddwMzyiMi8Q5+JTWE5leHKIUIf/YQfZbq9qwhki
eUvqqyD+gGkRxzxCCqZiTmk/Oe9UkYjpNRs9Hr8tVygsxS02g2cPu0wrME1fY/cP
Ee7J+ReoFsbW5onY0AOBoC+WCnXlxQeODlhDeFuR9fMtbZ1ANPAe5CZ+xDuW63di
Pb4f1I67ElijdguhaNJdhAb2LynsPHQ/J4A3u8ZBN2nwSmhRMe1/qVdT5dgDwWvL
GSr6w8YfZBBQGBsBaqIzK1sxgr9t1r/CtNlj3ZdBo+mqPg85pb410PfTgkUHTIwY
SouEfNFh7irXSEYZZU/3ZaYs0lXJGWLB11EvLEyq9Ifafv4UQm92Grbsj15PXxzU
RuVrEXTbAotvMBHj6ewqK/2MMzAt2ohbJQwU0q7ANOHJ3YwJZGobs71N+2xmW2pg
wyzcWGPvnmXZ6tPBNnh0sbNl/7MhzznIszh6xeeIKhPWEm1Dg84qvjfuz1lHVuSn
0+FB1xtLzuECWtf6XyFP9g==
`protect END_PROTECTED
