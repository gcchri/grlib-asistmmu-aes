`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0d/x1BtqHpqY/JURcrKgmgOJzqverHnABMOLtlPUbE7sBYkyrDWDiyLBPQ32qZYq
MZxBAOBMAzVMWUEYVEIPvh9uMim9xay9fj+S7Xybk5OLuBOQmwy6C+dCO0nCaLfy
Rx4HRu3r+wSaVLI2ngYFqsvN07vxT9oUZFStW875WfO0cAlDMwpXNlWCJTjlwUBa
x4kDrmdYE2vYvyjD7lH13d45HN7orh/7V4h1CkKFqUDykIoMyz40djmexCxCqh41
4rK5j9flVT8VWSdssKrsKL37XOXUCX/1ADqtvcoynrmuo35LagJe8HLffKKSwVfs
`protect END_PROTECTED
