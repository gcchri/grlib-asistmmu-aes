`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RQeUhFK8L+CN7wIRfEG85NksVhrI5YDN9bJFQU6T+T+Kkci0Tq3dm4j96wMIybtR
MJx8pDkdCNIrmNBxSOxliphgXGjHblWGZAOcFNEyUVbIEVrvn8L1fTCPwdVzOFSk
h5yun7Y30158DtHY2vPEf/xTTcypA8/6VBeJKJQyCyDOM3/Rt9Z7UdG4bOl23E3U
2Ijrpg9cMe1RZZ60gIMPtgRu2kKbJePHKUIgl7d/hoTI7PdyGKQ3Nl0Y711u3D+Z
+ZFxD0LlSvYh9MoQSw46Y8oHikDpGNIciIGGpSheQiAmXkOb3zmm1r19W1BXgnUY
elPb/dPdUkEoLqhzUjJ+WimavSsZsAv9iyRB187ijIn8CA+IWgDeo6svJqfYzvBR
QO54vt4hlSTWv2B7Ezati5fj5kAk31Ny1RU3/4C9Tsmk/vRBomMUUeGxsRJt3+O8
JamT6nroi602KYIxcUL/dsuquXm3R/GFRkA+muDjsMXENy36qRDXx65vvdsVkooZ
ROFgB82O4V1Wd42+WbEStiEePpmuhCegWLMDLpwOWCfiNMT9f3ukXZ1u0weWsnMJ
v212evQ71TOve13kKkpYhSWcQvzY2hhAu+uA04t1eVNgtcZgPAfxSRVbFBTMc580
t1mTfA/lBTR4fZHkTdfkmEY7JUC8Z+Pj/raqw2vyh5AZWRJRcqpcRDYDM/7ZmpFP
esp7rMbWk132CzplaHDSc4B2pEK2vJxKaPxWt0uodAHBjx9jNa1ByR7tJptZJmHb
KMaHOe+9Mt7T1pBKSP8apthCTY72/KPcQBEUAtUt3+ebyndJG3HgO/8f41YFsCGx
kkNaISUufDA95TQHIvPfXRC8HUZgovW32pwZ+zGC8XsVJEj5HgS2w/UgsirKhYkc
RZphouTOyAFg+7IuFW8UcanJHt5NOzFwpbFLZeVs1cQ7DeoLyEh5XPh6PNmdZd48
hrlAitlqUI9/9mBGD/KlrrGQFUIURBmGMoUN0netuYmQmNLLgNpnWJMPcJor1Bt4
MkxTSeX4t9eMTQa8kJagPawl1Im5g+3xshBBdcXFb/ZvAx5dEFoZNVBNZ17BNhf0
V4Cp782JAUggjiPCjQy1kxPRuAwbRYKCTbjzPBtwj1s3M0kuFke76P/SkiYOKC3C
GSwNG3BAsQG699C3vUSK0Q==
`protect END_PROTECTED
