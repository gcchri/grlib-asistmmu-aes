`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dBKF3vhQcKBdWdbxubAHS7eDaV2SI2DAp1fXqj8gGjthfPHz4g8k1WOOh1gP/FT0
zcBd2RVOIvtD7l1PUVQe6y4wJKDgkx7Udb0FzJLuAUUso7UtsuOaVBXiTOQMiAl0
AVBho9F0SON8VEHg1oua0v6onezKA4qWM/w69ZZODA4AnTf1bp4W9UpFIikT/ec3
QFHf3YdJa7p2rEWUdDQhq8ltsYxAw3vXAxlpmQ5lX56gkLIOnPG1aUEsAvyCk7RT
CndzqEClaPv5OSfGd5cmTx+BD37MwDxj5SZoyZZlUgRHoRL40WKclza8fJ7g8Q7c
fgvb4vzmngVtdc9BzN7v24HioklEmYT6VW/hd5GVutj8pxiI8ctFglllN7nNS1Nt
GH2Iqs3T+HvWfc7KTFqWl5wWpUIOeKiDEI44BMBFHKndNNWQvYvXQCEk4QjajrBJ
Vy8nJhMBusoeyseamt2iCjq8Ote6YRR1hHsp2O6B5tVFg/IBlu8Uge3IqZxp6Ww6
5eNwqDUvbxxZVE8y4frjslLzkEr+gAU4sMc/ZzWmEvg4xmGnMx1+WoTnMKuAZ84p
`protect END_PROTECTED
