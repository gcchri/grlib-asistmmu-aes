`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
quftGPV40DaXxWsYsis60o9L4G2vvT0aRNNScd48Fayx8uef9NRYS14Z/TezWYtv
iHsBrir01E8twf3aL/kMdG0TUt5Bv1qbTbgs/rCwJ0z+atklB+PRt35X7BBMSLfH
FH+AX26iuEXbt4bxZYmo9c1HhJDV2GZxo0cPl4hgeblCE914wuVpVcoq2F3WKqsz
b0wKjLRO5aZTF8TH7MA1Xww+R5TaEk0NEOGYS/S0j60MKMJrAI/FKLJqTo0zo3MP
3oCFIYwkxj5/KgJhitey+BPyGnYwJKgEyBw6ZABgv85UBx/b1CM8dSibz7VXXYlx
pd02/Zvr/BSp4Z3o7HEPTIhBwDRFqHknASHo9WPCbdYDjupSYNpPndTk2fWlTvFh
bXu0Ia4qhfaR+Gsoo3jktuK4bQc9ou3dsHM1F+RHxzk=
`protect END_PROTECTED
