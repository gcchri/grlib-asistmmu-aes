`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B6apDyOynV3NdS1KZCf7i9m8D0Dnlg2aTLYgv2pzrPoqlNYK7UjjGrr9qGueLUIp
2glSM24Oizza5PxUmk1Q/k2dGQq/6E3lu0p8Q/wGY8wGSqvc3qy/8CAG3lpNSHbL
5m13n8SqghzVXhBjPyKkM3Qc+zY7mVwDhxlStntvqlsCSDv7LtRvhdJqkASQdChk
bVGfb+5P8Ft+vTbVTIe8ePmNEtXd2UMr49fa/5+QnQNOgtIguxYiQomj143SnGQi
Qb5d53l+cNhnFc4c6Zlt/FN2zONIEuI2Oylm9+v9jZw=
`protect END_PROTECTED
