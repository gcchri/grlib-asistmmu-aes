`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G7HmhPPcyO6srmH/ZSNJoEJLNzKi7wDw1BA6KfqFakWOm48gBPuz9IYsw3jnGv8V
uS1/QBevrIWiYmrV+GL8HLKIIzXVcYQ66ZaJ82FT6f7AWnYFMRI/OcYIa2G5gUtH
PLzlN2pyobRUndaneukPvZaNEML8r0GUvcX3efn+5MhZomKTo9b30LaEGG97wxxB
+FTrj69Eun1cEMR5d6CpaBLl5etWZ9+mTcGklOpDAvdm9JXT3tp96IM2wAuPqtxF
4LfsxgxCEaMmaoj5BfF0I/aAC3HWZ/HWoH2pyBYEPXh7SyJkjP+Tl16G+ZOG95Ue
YcXopMG9n8x6N+LmSoZE8EpV6h3Y7YV2C9IDXIQyhwPWdviEXCyLCseM0JV+gs7+
oxFq0wyiolwIM+DpPsq2U5P725Du2qiKPZG5BG9ZgnJdzLe5RBbJhjI9x/2Kn+QU
pYxz90t5+MgSVMKyFWOHKSo4bbpoERt6/z+EmzJziimCidShu6hN1GxnvIljRDzO
rY7e1jivh2Pbm1Pv52lwAhu+mTzBIxRjTSqWXLMERdFTAbMpHrA8OKYqTxBQJuNB
7w0s3AmF03qEC8CE98CL0g==
`protect END_PROTECTED
