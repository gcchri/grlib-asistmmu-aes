`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uexupefzNqz7ASAEh98QPGMeFjN+mcsY1k3PIuL3J4q4ZxrHjTZzbNLvNIki2A8m
l9HFZ6oANttrpLvpKTHP6xQE7R0oruZBUudAkYHUuSiDloJhuR1Xtz1d3vL2xHul
c9bPnLPiAEriCtUwmRNfLNAhoWPNZcZBmXVhNHrutnPXyvkkwPTG3/xglzkLX3sg
MNrl2oEnVmmRLeqa0dVAB8axLXxWpNV9tEVyPeDmUVuW7sACYWD5OoCyWxAjhfxU
qgRuE0BrjL/U/dPKYBc1G+JpdW1cCZ6EMWZTP+22cKmz3PxfBZ63u/kpFnkkP3fm
UKQI4ro9b2hKHBXljcTMIe5edDaE1aXg6nHzyWUvITtyIj9Jpe4PuzYg+WYByn67
0j0nwOaCCz4KZ71gVtQHbjecdvjxfnjWHbmQ/ZgzsLgXoxba5RXez+XFRbn9q0+R
1BX1TmM4H8wou7TZR4qpCM+yhtFCMRVqAdychgR9vpRzC1ksAbN6SzcsoQte3nIz
kIAcU9I+5VTd7OVl0nZfZoyNrT86C9u3+ikzf71xQE9VltmGLq5rJG9sYIAo91fZ
p7A9P70kbTT463OiK5cz49q+WMGdDUJHZR/PtLAJ7fHC0/9BowJsRg6AfrOotw+h
dcrWWQpxjGig7FwVChVAD0iY6F9J7oV4FSsPmRYR2gHR9ZzHZzVrzypIvlsboewe
TF9Qn38I9GYW0SolKn47BxpU4PwIqhXCFy8slmn614UT3oo+y9dI87w/dX0G5L0a
24IfkYI0IQVc/2bvjWgTLsZbDonJ7bd+UpdhRKfxFJRWXftD2muVCYJRV1igt8Rt
wzU4N06dLNgOEMPZ2+ZOxBr3dFS7LofyIOVZ8bmnY07hd7yBKrHv1jXKhsE8K/pd
k6c4ZKs7L7YHk/SKGl316zda3tWBy+Gf9y+Jd6gpoefnhRHhG8CsdZFud3s5UxAd
UwIOGweHxXl1F1w093ZL7sYsVM3m8dupyLDNJfD7A4PJjUCuIujUca0TJeURNHog
YnXu91elHL3X+e2/Zv8uIQs3mzi20YsC8qsUHvnDBJIUCVsImCEvCcnNz9gMkGyQ
rwPusDdTD4arE9R2a+3Jcdnnc1q7uchuZVxzlVM6vqhdhuOWXAMbnHZpbN3P4JAS
MhZkb8SE6uBfpitIzCzjyJ4yNQ0J16X5uW8ejLOMSqYq6QuVlgg5cxFhQfmfA3cw
xrExvrBeZ0KDywDg2H00HTVCq/yCy3E+o8W7beVxsRBvW0r4xCnUfbDVpY2Insjb
`protect END_PROTECTED
