`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yvaOwM+5RgykALep2ekgW7k/A9P3hdt3DUs+ihe00FZH25BdQVfXLAw6478tfRcI
8F49gxjhSWwN73xygp9klCnN4+lrGUdf6ZGwlj7cBnejEiIbtCZSCWcimUtRtksQ
nTjTWap8wl+9HiGudAw3Mn07jXN6NReQna+jgPxCBvVs0/hlBM2/g3WqqRALQ+Qn
0IDEML2eOy8WRhEol2rZj7eZFIUl7aaGBzba3QGfkm8euuGlwWLw3UCowqRRxFkf
HeqGERR9OasHppKixUa18g5SG91mfwxhF20XR6bjAqFMyDzYbhWBvh+PrcoQlz/t
ILSp9ktSAtTdXoFu+FSoAeCn/euGEDdBACCDBYFTWSEfXUTTAWwS1RNqe9DNoNDB
f8ywOUV2mnT0PqCLd30VXmSNJbXZU3//bZ8OfLyLjevUrHwVaxXPaHidtMZp+r7x
NEghu345zIHYZ5CJodQp31hTbFYXAKo3FasRcpetfNh79hCsJ+CLe5AfSHfG+6AB
4YrDyBYMSOFtu+SJ3P7EKDQUOz7csHVBIcx/aYbwuAXXoBXrF5hmQ1DveqIqBKka
HpscAGivhoFmNIGOIA2BYWj3ayd0oU8YIgSX9DIYJ843YkLpOsSSKWCW7NpC+cfz
HAI7KKt8vlgcPuJthObpuHTVs5dDMc2Xs6S0nuG4CzIkMIZvs++yp8lK0+uTs+hJ
KbOWH+NQwoyojI6mboNBpdVPNXQewLnFnazHV5dTSV2osNm0aQj6xgqX9jp1c9Sl
DExaKv838MBo9tDITra81P06KX+XPM3OcWgpDEbRRSv3+zxkZdnx+uQS2vXpzozY
n2M+XxO5danEQHvho53Q3TFkThMsWYo6WcS6GxySANYN5CmBCFniMRLpY/48ZQcm
hGN/lPmK1zHKfRnp+IEMWZJMzAEHDTRoiiw87TNRYtBvpq5gDnAYYV6vteP3/fdT
63ZdPZo571H3dROJ78MFheGbY4tYx5IaCPbcFoMpQYCMNrLFKAjNXQ7A2UK2A1hd
Dqs/Fhu73E1RmENr4wqkAvtYTY1PrvfiLRUkGGdEzHoJAxqVn1HLq6mxr6G0rG6K
SQzyJ3uqKxSHljMedkaPJp/towNmdEgNXktMzFKUoW2Be1JFSv0+8wsg1tZzQmPF
2ZjPgT34YUfd92l/TRyrNfCgb7U5PaeOJRpr5cl0dcphXX55B8rpWEU+S4ofpO0E
dqv517gHHaPoPoS9r62GJR4n7EFbvM9v0ax1bH4Gkxv5GuK0xI+bWkHjboFcDc4c
AwWV6FcPL69gPmnbnIJvy5LN0fPduIUnd2w/w3GXri7w7Tf07xhHfBGEDx6oQeN1
pUSFh1fazvHdH8sdxlpIIf15HR/CfNQfOACCeYIK/+83W1fsYUwX+dhZxTKSUAyT
ALw+tf+eWFyLVdu+VMGXvelf3F0pc3lxV727CEIWcHnSUHfQElM52QEVmDJUqGMr
bMGxRibxuxFdboEMwelpNpGHJrWGXhF/CBKhu6J/BuktdD0SNltVRWZJUZZoxGdO
VZGDwNTkv7l8GykmvrpGWLHjmw0uJJGlrRJ1539E0TL9wLEUt42++igTrCywlIR/
HMMDomoXOgB7lTGqaN75Rq8T/Lqlw0tsdCa75Wln1WaqGhILQaB1AY5Jliy5oOtn
nzp/rVWhTC8StAyaXvcoa7EylGTlTt3p+2SfEFkYTpNhkeI+zvg2VEn+0GNK+Hnf
VrO7D89ph1iBrgw8TFpPwyaXMIp76RBfz5JjNbr/Fh0FrMaFGruWjB8LXQNYskfL
7jlbYXNnX3mryVNfjpg1ZunZuM3oLnt/04puHixs6QTHjcTdVniVblmhUdLnwexu
XpbmAyYdKGxoT5+uS5Rk8uHuDdJkubsIb889S7CAckEjPzwMjxQSEZvmjj0eZP2R
RW/9dNa05MpBEqsKC7vhPsUeHgZAdiNR2ywc9nP2hLsJgq2aGJ9XY64XgeElRV7o
rvaEYyoFsUfqMlvT1FMT9rPphzGs25uObL9khVhsrjTWlLgBnxIe9vnK4cF4wpIc
8fpTylQAd7TFei/KX1iylZuR+nj3CnKP9H+5c0Nia4tQ7QhTqQ1CwHvX+ugFTbfM
LBxBJsG46qaeA4X/aqEw6RDHBhtz0sE6xu9OCak0gMpdzV759qGQtbJDPVXaQs6q
pS5XTSZcMH2hI3uyZWH8WH36G7/8pWuGpWwhAbCQ47RClyRM4Jh5+GuyhTxsu2lt
rth/EA2DRECZKb/GbhCESn09WCbchvWC7vqISpf069ROXpPM2ywQBIzs+OFy3gsp
UTkdgxoWxJMZtnfToWSLwbvOCkt0DsdXZpdzwPG8EqlqU5jz5rYLhW43drTPmHBN
WaMvtnBVlmEzvVnOR7vwFM68BjkOc5CrGMO5WgguWaLDAraDnsyC/mZJN/0li89L
a1KjfhoEdNrTWq7wn16hWkNgtR+AnSAa4F3WVEvnnOaspdOZ9fLGhbe7MtG9NT2o
n00W4cIB+Na97wExQhvpQjb3wH4L8BVM2iFIqSLSMI35ZsayAam5g/memLHYfpFa
Y4YOzpZqNoLsCkpJ1/AmBLSm5qabE8/AFYNHcEEhwN/d5NnAO1Hy4QlBp+CLfHA7
gMJOxWQCj0E4x5CX9x8pZKtwOgcUZ9x+rRLNLIyq6sbqqM+6onBramO1Tvm8lOXk
eK87IqVN8wP2oOdrpP2LfgEPNcH9wnNA0iM5IGBkwO3Pq1GWsSFruGxEG5hNW3Gm
YrfYJlZzN6/x95gX7MR/SP18c1blxi6851K4qW4B041gGP1PIIPDkDT6TiqdHTKM
61MPFQFJJKZ6XNkweYyW1SLX6V/GBkzh/X/ZjBM8jLdCrVxkBVI7F3of7FsJYNhD
qVDGZK+YmZf4rerd9IZgXy77lTn/6VcwcIWDrJGGmkHF0mDLnWg20zi/1s/IcS3h
M5ihevQKstK6Av9rN8qEeRLWm01g42p2oDswh67ui41HtV18LzSuboW1GgFNo0On
jwiJgiSOFHQ0tB7b6Ial8oISm9MUWwAB4419N0cqExAkCcnxVSSFEVXCUvrTqY+/
RPtE6emqbOZmYb1xCQxFff1/fgWC0ahwihl7Z2ay2tA1hil38VpQ16BO3hafmoNO
3uFXWqWMp7T6hKH/c7rY/PkGW8fh6tQ/Ufz1NCOLKcMEdtg7/ukHP32HgTU7zkdv
VPteilY+adx2CeLamzTCbtT/wI3sTFQJ15pyllzHw49JY18LNfIFHRCgN5ASI9CZ
14RpxLJlhNo+5nC/sDeKyweT/KL2tTZQ+AFhyu4kXgvNm5LQMTJbqTkspp5C6vVi
X7artaIAUDPv33izwK5Fr0eToJ6mb4M+yg2Ebw+eyy9WYFBHuJA05ADWGeiyDR/r
L67gcXBS3K9dhnHQZ/LRpA7sl35LrHvra2dIaS9/w4FOnBsgHURASZBwjatwjzRk
gjmLpJjUmHbw8uFDo41HxlMcpI3L2vcNEdeK6bvQ78IAji240NoE4ZWR2+8zT5RM
CLwESnZRyivpz9nORSL/xYOCvX9POI5wAf5ccea8ZLvuOo30dsTZ6fOyIMh69iPa
k8Lz7f9UwBWERvMhO+8UVQxqQlqQDxCIYebMua8ZwQ9dJlGEGoOTBJAj0GWPHNJ1
bB3p4FRuCTEZX3y25PpPhKm+eKkA377aVQO8peWlmycufzPxjUocKXeD8yXKTLz1
ejk9IHpkBNh1mT6xGHF5M0S/M5V20HlfrNa6ukYJt72IemF6dHAVhf3OoOA4i/e/
jcFveZaWdUzwB9iS9ESwadeT0T8FFe36Jasx+zidTRrWGdrA2g5XZTaHudmIxPTQ
XUcmk55oKePbIZq9hTukf/O/kRikna1g4+9Gz7uoBEa5risKPUZaC13PcdZd4e/i
y3fuwuCNDWJYo2Wwqi9rzWW0AGIg5y7Fbp5yKAGMX3S3DHGFuOhhg/KU56TqUD3D
rV+HqW1YTQPcw/x9l6SywwrGi0MlMYdbT80vtGEJJir6RKfC+CwaBor3wkBj0Rsz
gnufatXJgI7fH2KK+wapRXpweM2VOo4yFms+VmLilDGewJwaUB+gnzJ0RcJK/UI5
dMooU/U4VnPllo6WYrwUGTfyufgA0YCPMvD09G4JHXDcA0xF7ZF3QCUwyDVfk3zY
R75QZzMKC5CX60+eVOJn1zzen1bWM/7Bz6+e5CgqAZ/tYlHXgdvs7NI7fl/z58D5
zAk5QY13wXU6IG2/Pu82gPV6Pu5wVErCXSSwQjxCATjQJtloP5tF6w5l1pNoVDRa
hpXO9MHg8bNrS0qfHcRZCKUwyWAFRFig6BjZLfRYH8qsGgZzSdW3h32b7BdC2l95
AsxETglGJ5SVcbTi9FhR/vl4b5t56K7W2hZrx8Tqj0Hhh2coRMk28zX3BBGepGTX
E1vysKiCbUETUj3wR1LK23N3syenxJFbMSWfM2d+2qMb8s5By2j1GNLzcC7wuGyz
I3l6zgyPlJoA0vt7sYtZRzWsy/Pq0lViNFsn4GsUz+SFyk71bstqsObRvXIcfzUA
W0Yd8hRwGdiffhDU9gZ0Z6T851wkVMf94zOVNY6+NCYaTZMDci3PkAHrUjcva6ix
22NtPPXb2ZiYm6ieaaJItb/QAzYDw4C2fpIgZsldrTX5c7HhclciubzcyHM72jsD
LoCxGjf9/tn02ze7EiP2e3ToGl4TjSzQS3CGZ0sysw2TMdIk0Q16zT5auE6DErrW
W2q+cHcxzk/m3Afd/lkDuwe489rY5W0GdQm3KnM1yq6z9h9XB1advaET4Xoadlsq
Q87+49o7nQNoLBlt1JdvuQrDS/pxt7KjcF0d+M/cHc3H7e62GsATox9DF9EHSqPS
NNsf8otrZbkGnTwT0oMS1TERnSdPUmQgb+v1K0WztSKEYQah5FBXtc1XXRoRg+t8
W4BJqDJVi8zO4JURPBW0Ht1rSPP4VNWug5Yt+uRexjEB2ItFBF6WCoDrBu7huACz
CrdSIToxdg871Bb23y2K9UKlFUY5RRRY9VgdwpwN7P73ac8H24kctliM9hSwSC0I
tO2cBG7v/KAlKyAnIyars13rPqV3qBHXO2NTXttvIfxhof30xmnPMujv1N+CDPv8
Vor+5TQeZD+UZMlxUbxhs5xT4DZ5mahug0ooRpmC/CatmkXK0CUNTvy0BhRBOFXR
SP6gmqRnUh3SZyfNTFnXNuegvjg6nIowMYxwTT/iFdwnlba3DzgbDus6xt1KJxq5
LkAVevrD3uH8EQsIxeNwCSj76etWGLl8kcSQEvY6n2xxisLq8cswaLwX0PYUKt2Q
OY+ossQp7GzsMdE6+rmLAHoEZX1Xkdc4zzHcU02jslHZ1eaEbPN9gp1U1q3b4nYL
wI83ZtvyTDaL1M+rVgxvli94GTqxxPVGp314E6+9h08g0q8dS0flGYR6mUPInyik
/Nl49FSRE3ezqH0ydZo+viJUmLFBvBj+BGxt/1uSDZbQdNVOC+pVBhulkVTrDn4N
PrOjwGl7h7jnRpT2klagX09WtX4n4hX1+lS6mdRy0rxwaXoDKsULUMTWT6MGFduJ
FeSKPUocIj3xGmLLKeElmh3+89pi6Mv+EJlJ+ykq47rVaONTRYRyu0gYE3G/1VHs
kZf3tv49etpcPKtTkrlPEdCifqYtg5Ribw6bbyAXR8NDGmqcj2rSCLs9JS5yd3po
9HQ+Rs+CrxlWFAEqhk1+CTgbj13eeIQoZJZyKevaVLis7/IPchlE2+5AMdB0mVOF
DGxmTlHqf0FaNTkMH6seuElFlLUFbqsFrvtKGwayGlP5x9sKRKsyYcifNGQZ1caE
zoPTHcX09mNjeilLH2A3VuNP+3tTKAbmpiUpsqcqhHfu0x88VTMmzytMxqhjFC15
dH7jEeGBKhzb42nuSUN1k4EB+0CJgGFkVkM95aB7z+TYX7NC4HNBtIzMyetyaKah
xIxkSFkdwNlSmw5FrGY1bUBybyzCycPe9bFjgUuNla22I4FkIl8aGNQHzeiCxxNf
llPsd4BoNPhLvxJ2WmJGms27WlMTPD+p/Noa0Q+QLL2K6M3MxxkiOmiBqUPSw1eg
2KjiWnei0FQwsRCidflD69VpQzJio+835GRZwrf2fREzBS8gRB9UFimGJOxIEv4P
VUj4ALprI/1N5poUh8wnoMZ7X0CF7V983KnSRYgL4cJiTcLodyknpldffhDjP3vI
3tSn7H1iSsq3KllEEMDudEvtMlIs5zhR0h6V9WKPm+h33CQY4Wpq+QN6mHluSdCt
5CMuGHQBayYq23rDvJUgq+C2r+2Fwp+NXwaurZ9SZzknwNBYZb2Abu0TVgSyoIoD
b2exAVTxTS0AcdV4WrNh7HcVL8E+xLsduzJiE3Sns9QHWOE75r5fSY7YDWmLo0lb
KbeJ2RotwOOms4mKoaUCC2oQJ0pEJb/SXWLD7KQ5T5LxiH8itZKLJyjbB//PlI/O
Pxgyyd5YGicZxWZb9snRzgDTwLWDyiw6rA3KnlA57ZYi9Tyzse6Ol5n1BUS6q0+0
IxyMLRuXK5KTiGWdfzTXd5GXpUo82RL9sYSJ/XIlsbBUuvcgo+Q/WMNVca7dWNMV
3JgwUupGqaxkXMSnR7gZOk0ELKovkPrDgQOJS02eTa+XbyEbjygGMz4MsRtm0taP
YPRYYDKKBLev3LrmhTZda7C7xfp3UfoIrVGID+gDr/jTFjT4toBQBWnTZL3sEY9v
Om6ccjFVVcsTKm36/9exd55Zvzn2qowhMs1MYh9R/FlTZO/WjC6tmbOb7XAYOGPe
dNV1YVt42eHPMrJzAGb72rlLRkloxGGC1C5JJ2sUXJqdiwO+T6fCBOEktxtXNDfB
9VFNJI3RxZt70N8cBmdVuG0DPFrEUJhK9d9wbqnVJzolhc1zTXIYyxWTbtSRWHya
pS9Hv1M4pP+aH97JLhjknx9PO3DreXRxFTVqPu5XKld2fXYc5Ky/oGRyJyRuMD4/
iit41Ie/VA2Nu9uYx5+zUIHpr+pr4VHp9zknwi+ySXsrTIJpHpfNpAFBtzYwo5A0
hu9xaDedT5QRzBCkCCkhn1+lnz+gGAk3I+xyiJv2UnN7EU9qy/K0G/HbgCTX5188
WJtAx8V2tPk+yD6cP3e5V7LJCV+xVowFF6pw98TwrPXMUlH4PurZSvZ5aZzIw3OF
Rpp9XLwdKJSksiZouR8Ropau9msOuXMr5rLxVs4viASJ/NBHpxbB3N6bDn+BCUFv
KaO40jI4QVBDtv5ojPBIbEaodtlmBvln497eIi5TwRbYq+VpJwSpegZotXBIoJkS
ZVYDtdYrx/F/btZHPKG5++gwfD2yt9tqV9vw5TtgjXCxAnj4hj/UoIfXUhTnROv2
83M4h123peetZD8VCMwSGDjs+uQi0JZWimHQEvUlFI5ZixE2L5nToFo4B4sNa3M0
0gMvxTNXw7k4/bbqc7Qgp+yptrJsKj9G3yR5cppHDr2NdHUzUXFlOdgcrCc/1q+o
+G3FE1IaTGI0uWFOmMslc2/SWedO+uqJzEMh2lr3ttjHbdvz5QFEvJt8qvIEswXn
hQ7KMChZrJZ8Oj7UepjfOOzB1nq6cE8nOzSec8Jvl24oYeH65bciSsugYYzWOHiF
g1+kdz7N8YiTbbxqurikwCEjejk32e0Z+MFZyOpYYTa/DEYIG7fmdl0U1pVMIWMt
q1izcRb0n0bpTHE1nO7PnZIGUoEMWzRSCEyBQ0X62wM=
`protect END_PROTECTED
