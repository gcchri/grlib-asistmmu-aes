`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eb0J0zhNIiRICs+1MAN4iD0Kx+1rsggSefPut+syjhdI23uTJYNT5qysVGSL+yhv
YxLtFh/H1GgzKSvovvcg+Veh9VN7svj+DlOZSu/3Sg0iMUZQ4OQxaV+87lB3VpJg
T/Kc+dlp6YZnqNpCgm6rFUFUVnveFIq4WbJB2QdILrLd9DYmorDFcEM0ZLhOHddT
BIps4Y6KjO2j1cZ5Rd4zj6e+49T+Vzq/2mJGrLIOdHUxYeOhpYiOHPvxoTiw2mHs
JhWY2rE3LvRHYzy/9srW+XUoeAUX3qTbTghe9hz9JuM0ObeL2RZmWCSd/I5XpXmd
`protect END_PROTECTED
