`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MPuLzh/Cs/ukaJsx7fTb4ruBW3OPSp0E8QF1/CV2FV7DqlzHSUf1+y75dv7y8+dD
Nxq9XAOpX7IMvp7cJFWMMT92lWwOaDD9I2gnVH4RZAloO3bJLDCOc5r3L5NpXh23
8YN2RVM7FmQWjEsr8OJ1fZO/Tx1ElVrHI8z2nE19ZnnzsUmq67H6VjqXyLFV+ZdU
mdCaDRt3Q4Q6RGUJMsVbdl8s5uaIYmxzT1GmBc1Q5UHQEcOzpsfVozS6UzHlbUxC
DJvMJE7Z4rk6jNglFnsCsTBpS1uY5XmOHvgisGwQFTi+PbALkiTb0kjQ1c/exTop
3z+lb3QnK23CjJTEHi/mOwHXmmkYO+OdONhJzhkg1D7UdO+MLD+hqtE2FRChQuRZ
QLTfflRW6QM62ve4aTax8YJMPpMLBmFhMgBm7NbxSK4=
`protect END_PROTECTED
