`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7UC6sOdv1/tpDIZSOmy4AnhSJlExsaFoSESkRsmY5wC0ot1k3Q9YpvqVNAxX3rq
cxMQtZ4HmAHV9li+rBXF9NSyPDgVaaMkZVOYz5f7nMQRGCkpOdLLfwU4AJ5ku3t4
9puXtLRMmBj4FE/K2HSGF4QM4VfwBN/0g+6aZ+rHN881Yt8LYWFmK8YtJIucQtdG
vR4y/8kbMqU95P4DZinoj9XycnMohamNqwgNX49YzjibVFp2e8Y+0bRk+JiH3oqD
6R/UXmQBIjuX99IhAgwqKsA+11b2dGWjDLrXzHQBXFJ9mbPTf8I5kJG1UyuUeX7B
uHqRpnzGU1fcKQcggJP0Jetvi7NvbedElXuAFPfaNNke/2Ol0KyrEgbkpHomxWq9
BmDxfGmugULilJb/8YFqwRcbu3BYukZ95yOAjBQzNWY6kFj6S7I8uqwFqfD40hMB
Jbwq8KXm2sXXlfELDjhLvCveWtPp000PuG065sfNx0mbzzXEmQ79C3AdaxCj92Mi
e4m+GkoM9qZkN1bHCPuIqTZ6Jcos/+tGiE1tNxIaFbhtquIkNeKHAUnCAvb1DOwp
nFJbzcFIk/mRWWhTK5B9BQFR+qH1BAbOogXXrv+77KVl7Cqfzcto83E4JZyLreDX
+40ZTg/OZB+i8OYWl6ulIMs4hkhcOePoLJX/m6SYrNvezzbw7FdMXU05o0fdaz5p
8D+Q9BBgf+a7kmYfQRg77GPeLBUgrSejd2rv1Ud0u5Hwqmg7X/LIREAO4dJcAhV7
3Xa7ZlmNj7051HYJxOS+l/Of1cuppI5UnTDREXB2wK5U0XQeGsgugMvH9Dn/xaoJ
zi0szAepAPSAGz2jROGiHpbc4+xZpS1SzTrY0mBoetxFfobDyTtfxZuMz5WsNi/S
vLrA7edOkainzLOqzc8rxRAHeiz3CMeR/l8AK6IgwSNsMUmd0F5EECyjVLdwi33C
RbGTRURjlnp8o0YJbPqbY6Db042DUwlx1DJGuoUhjPmX8Q+Y6sAH2tpy4omaLWZH
1AciXPpC02lNSHMGpUETcCmgYYfcbro2f8msNTsb08eHLiX10URWLkfIVJWI4AvZ
p4Yx7AVJjsuajvJfP344el1iQhP3tlN/yrwPUmUrIPDNzJMiSiZiIIHo4ZeB6i4d
x9G4Ynf2pNV6FxNusEBAYGjk3KhWS7pqfN5dT1Gwc3SEnKwuL1fHoJCn0kZhgXrZ
jzbr1rjUp2F9qWJ0mjEV/ay5DlUDokdmvb8sTN07T+QlOcbf2qhJ5ook7Nu2px2N
c2CbVY7pi6sGoBE8KN/MZIuoZFWEoLDLzZ6vvga85UG4gZDqKzNFXatxWsXp5z4y
G6EdLr6hWrOjn0Yxi2IDM6ySF54yHfjypzAFAASYS9g=
`protect END_PROTECTED
