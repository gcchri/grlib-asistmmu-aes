`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BKjGBEde7du+rdGQw6GhKePCgNYa2U3tKFUpKIP5fP8ClaoHq5wwt2IrvuvVh8Fo
F8tPp3I1GlqajE5f4bBj7mlCDLsanDCiFPCTVGtBEp3jHEHbO7mq8bqiIjL8ReMp
Whi7Y4K/Q1XPiknaU+FICc4Ji6YkGrRrcrLWWZ5wO/x2LTBJMWvgi7Gqm7YeKPZm
/W3iCQrE7bbpt8m+GnOEl2Z7BcsgI10mvyC3yr8ZM3F8TshMWSWNx6xBZKn9VLtn
22OsIi8p2hqcXkOVANF7RrZXQyh7NYm6kvykVCjKq0B01oQhxIPje8czDKQ3Imle
u/io7/66z2Gt4fp24HoolqBTRepO1mXc7dJ5Oiste/Pdg17fnHpRPEbRBZanmOEe
xg9EhbJGSL+KAwYazsmMaQ==
`protect END_PROTECTED
