`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJQqygT4iP0+VLojqS0s3bG5wXN6a1IHcSQsP82Z36XJMJvvxckiKgl4j7aKIX6i
16GsiWxDvI7myg7ox+UQ7uxpGwZZJPtpBeCJBGUUzdCdGKYrK1E0ZKxynnEuTZVy
2M5iPlmipZE7D+JW1gulqppWiUlmiMr6XRG+0Lm+rFfwNIWL2KEMQ4TDZaYEVCz1
FXd68LkEChE6ked7wXe0TMzviQXrcrHmhmXRIyAr6fggmP1dNZmjNPiA7E1RKZzR
K/ixjUzeNkpJo2ftC2lfVxUAHnlxMzRvyKfcSDi03fkTROtAou16QAvkXhcFDU8i
YH4k+CrPSPU1mdKYy1WbuCcPkKozL+9VvN0VaWYWaGeMbPpuZVWRyuK5TSRjB0wm
qz+9CLudS8EuLNB980uahtZz8KMNu+Alz2XZCnS8GPHj6Vfgt9DglPppXyqYdb1l
3fwvVt+bwF+Kg+pg0h1KQAvtqsA2FFDr1+GtAmFN78qFqAx/E2Lnrt8dhyzG6sZY
hiK7DGL1k2wkmYV450osFfqKLMhtX6+g/Rf9v3tSMM/kqNS1mP5Jq631WDBxvJra
iAaN1F2OferuTcch1yvXYU34nofP898JSipfwBrR1QFZ0KBhYde7U0EM4M0MhSon
E/57ojGGn8urT84CprNLLlNHkX77dth67B1dPuJ0fbA4Ng1bTrJ+IMUsFTtIuoWK
nPtCKGilAs95sM/lQKZiiO50Q7io7XeKSHXvHs2z3dIdQdLAHdVoWowWw/yJFEMg
FAq6BRcoaaG+74CQRkpw8/kh6A1hLTIpRQqiHFBRFaFVkeFAWfqrt7gznBPfzldQ
+SuIbsdtOEWQj+IopvhKcRjxHYVX2X5LRe3qDebulPdIvuAEcxTa2qDNQBrybFlV
MPHiDQ/hL9SEkvAInCgFqybHj7bgLzF4vZMBO8L/9fVz3Zmp6upPxHUj5w0JIQ92
tza7anDq+NZes6JFZPaS6TAAEg8xxbTUXtgiushxsNI/zgJSI8mjOuyxMv9g01X1
`protect END_PROTECTED
