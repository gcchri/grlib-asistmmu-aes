`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9F2REcGgZ3d+58D6VZUrR5E9krHKPtihg+ByhF6w5IGg6afMgYeSWr6J21iwCwRz
CAqNEvfj52HyiMTvpC/HzP02Pjs7uSv/jN4O9hWodhzgwIZwJ2tHhRFWwe4nW+kY
Q22Hr7KlRnME5ynunBZPasJwNCWvW+Ep3W7FOvglotJZDk9XnIvzZnQuEQgz8TUf
CmezFh0hVkicLUKcnecPjRafTuWJT/mNW+N2p6/tNIfOo+dRvvNJlIHWsc7kHE3v
UsZZZrn+zeCSGlwTtkZKPw5uRpbuLbdXM8pEqktljmmVrMgN8VnEh66Iwhey3kN5
crfiU6J/VnYA3CmqvJNovICBiQ+6HZ6HohaRwjjCWZ6Pt1rYd3or5LKDKxZKAx2x
FDQoB7HCVgN9p1CWUZw23DXRlcNpBJWf+iDKw00uI3EdRQm/9j1cuGxkBg4rqagY
mv5xlHNtzGA/Ua0j4Meta637GYZsHOBOhhTJZPQyeZPdiTk7iQk37VLlmXBlQDR2
Z4qPL5QLtmWe0OYttXzkkpN1YyeC7GrtgfemjdZPDgBTjUV8MnvZSaSx18QcVZdc
nz9r7bxpXyLH3gCyyEkH2jIfTv+xF5FQgGJTpTGq0Xs=
`protect END_PROTECTED
