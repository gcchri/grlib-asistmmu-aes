`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J1ek2scDdn3RE9bRHD1kRGzSyTujVoAbiEREc05YkiWA9Ehlu4bn9GfzDcz98GAG
ITXYXa2gtl3tsVPf6vFfKBYVme4aUI0wekd9fVY3UfSVvcGdm4y3PCocOqL1Yw0c
VUC29qmtiz0CfYA3VW6f369HSqcnMVZq0+5FEIW+NXsukYrmdN3J6le5Hj2vKGgn
h9yyITfj/I7nEXVL3I5yAhiRs1QyQ/gMXuO5dG8I2TCs1p4lUt2C9btLMg3fYoez
DryJH9OeuPju9BnpEETbQHHeUtUX8MIBpZIwTHPxneKGRoGl65yehSAqYAEm3pvj
zqOH5u7Fsl+1mELPJflaFGZ/r0lGBQ8u87jlBzXX84z/q1JxXbUZpt25gLkkcGlP
ve+B8Wc1ouLxzTjscrar1UxFGYooX6Ne47CFSUmwIF3QZR9i2qMrgdlgNiGNS7NA
a9+KAdZCVphkVNttdQl2kRAnGdilBD0p7e3YIO0KewHo9HIFujyfpMd3MPJ96pB1
ZShvw8/qVBYEC1Dd6YmD0t4YlDiDU6jT2iR1yYqz01QuJow8IAScEr7qycLTJO3A
MbAFhoS3Nc5UrMw+vb6GSPSfyl+M8dJ7f/vEcex7WBBRPLartQAVaSG3n2NfZC74
kSnkkEjSqq0s/SQoiq/8a81vpMXpN9h9HLqLZbZfPhk=
`protect END_PROTECTED
