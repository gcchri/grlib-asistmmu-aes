`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bTT71/TdEn/wVdvjT4MbFPwebP9tWXVkFazVleMOkTFg9xRBZJCukrlV2047wr9y
qGRHxqRbO5go2GbA99u8Icm3o9wA/gN5KQlVU0oPlbnfBD+q3r3o7ROI11KmlWSf
eiEUP0oj1d52OGz87Ox0eMVAyDqhNf1QmzSOtRCZi0VwdvONQvGpee9VoXRVSsYY
uX4AMu0Wz0zHbBCUxsFjtDVlIr6sTviXHCWbPiujq8KeJwkmOF2GCIWkrdSz0plj
TwAWN39M2IMqxC5KPvJTbeIJYwHmuh3tlP8GM6CmRm5+nJ303efREt9eAtCW0Zfc
CJL4xtM4zhctxFVFGPstm6R1hy9cVH7rFy0sz6woL0B+fiMgQ1QrPu64bBn0+iSB
mMX4HuySe/daC4DIxjhESytIiIaNVoxQ5yMxbJOcqdKt8hS31MjVnl6m+oeK9rk3
nsdCyKg6+kxd1W7NdyzLLM6NuaFMRE/Nka0RfeQhNGWBhkrw5scvr0gX1cxpjaPF
9RwkqUdUhlW1tNJGdiPvp8MdWE0wWereAVWec9cBlT27jjiRnArLBTvAD4wIdZJP
vzN61cjkMyS4DqlMXyn9BqViOb94H8GfjcmpqCmQpVQcwFmj89dW9pAi+p4hbbKK
zvdQ058djl9FRc0L9Py2Zw==
`protect END_PROTECTED
