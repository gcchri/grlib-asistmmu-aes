`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
noi9AcfWnF9MS5s0tx4FtSxPfgg9g9uiayUZ4hfRxO7grMAdUFF2MqnZEbh2+iTJ
t/DTcSEfRYf5fCjVY6CKBajFLzTHPPesV4E3GeuhDvHlcA/Gj0dHN0dUpIKP6Zxb
16L6/sFoBx5BWYBZ2TXdaBmwU37l+evV7ANYCPKUgScevHKBwKpkQawJD7lVI5uC
kjcoY3qyBIal67NvawhLOdkFQywWWCZGEgX6Act13PUCZ9TKK9UgqizEHw23MJ/t
KsZUhBHCMBXrvLbr6Tz6L01hbXyq3oUHal18RnsoObQXiBZM0jKCrhFc0IZRD9/r
6VCMC8+XxhYy4F+HdvvZEKPPgbHjori6S91h+e/B0WPJdZFF5ZFQxF+W11Iu+jLc
G788BXQt0N/pfHBl4baFLbvr9Dq+NYnCWNj41F1HO24kzr3QnlqBqUW+XVQNb/6G
uT9+KJtsTgktmLDEUAaK4bxgUrX28NOUF/Jg4vy5LF6DPwCebcfCbjkMs7Vq+24U
`protect END_PROTECTED
