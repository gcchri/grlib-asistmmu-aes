`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IPuvCPdLE7ra33ubQC12MZCjjHh553qnOzx2+eh9UH7Zz8mm0maeMQ68NTCa/61+
IgjvQoud0uTFzDBqtBeitVVAUl8XmW/F3lUs8utZwbXef4eDTPFmYFVAU+XOcVuk
T7LjVyrSM53ZtY+1u6wVJFrWtyspe1Cme7JTHezl1lgu5usplcak9cM34bWNhLp3
rZfdEt194C8AqI3I+aPWpfB0CigoTykDyQXrUYkKbsxb5016WGoglJlF4QwL07lN
Hs/USQF6Lo5Qy2vNy8aTwwkmj4epbgbePj4gSf0ASm4LhqmsRdfyNDhmz6jdzaTr
B32sth/N1gk70JVR4B841rmMp+oAIIKBJ8raKraxsQxnhq9HvvA12OWpQNbqOP4c
0uN6Er/ElvyNdQGwxL92A44cSBI/F1HJi1R3mO5CUFtKxZNWkDtAGHo9evbipGrZ
tMb6pPX/Cf2PC9Ppkx881XyojiVQvbxATYmF8X2qagttXadKYf0biuKIYhe/DNTo
`protect END_PROTECTED
