`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
revUFmQj73KhEfe43GYTF8PkAnUggIrwkDNPWl8CAZ684b7egawJStyNUl/ZUw7v
ej+bDwcS7SSrRnfYH2vMZmVznGrfaddb5DjqF/QjWlAeu6dT2nc+S33MvBxdzGTE
doM0UHAZBUzjhiEC+lSwhObamWIqQCu/wOp9KkcVGTC1Yv+oq4TYsJhClGjCPfWj
4qeJE61zSP3dYaeIA/TTAJRUVh0nGkCwcyZOJLeb8JkEMeRuxTqHx0NSqDtJfB0L
JTtUfuKHJ5DAggQ8xVjMhcIoQq8DXO1zk7k9XUiXcck+xnbb1C180A/6kRJNlNSE
7UL1RdQyrEMyycgYgsA7Z4BIXkCZ4aGlqCQeCfWgx/woqVWt8Y8NBI/9lG+rRbDN
oX4IO84th0rspI/PeWnTSwfJcu9mDAXREPktqGIqDA8UO1YDPPWYp7uEObRzGYSV
jerx5M9B2k3ESsjCDfHr2JtbFqcOtnS5vl5khnNHzUNq1uHs/b3vq7hLW51bnp1S
NiqyKoZlcD1BboiUnQ2eJdrSUCfcOLiaJo677yXYj00uT+Fckj7ynXECzAoMiUog
9QfBZKjOTfCX1OPuiFPyIg==
`protect END_PROTECTED
