`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/pi53Iisr8/y2X8aMoS7FOnbgtVMj23ebBa8LxQz6YVXm+wP/EqxgvBkOQnqquNK
1g0ijfzGmt/ftOYZApOP75t5rr3beJY8A8Q+V+B9LJIb15x6KuBkeXZZF+wuF6yS
CQtFqfix86+Csve+m6PT32uclPXAumzcTwCFgOggx818lahZwm6wjJZgjOw8/7Gf
sY1uvZcEC7R1Xqi/yUVezy1J5SuOjOn632LL4ykpXdDQcuqf+LfPofMVq1Bi3Mg+
hlaFAaICi0qOrneGO9JrRzIH0MfXVWRF9dOaPRvkS6rVnIRezu+PHImxv8Jpy3rk
pukRvG35I87o9uowIH+ASwoVoa5sf5YZ3BKxpZErPNymp7zo1Xtp1rEpFxjjh/bv
RxbtSo3UQCCbmnXO8URG32ETVKE1wOyoPpSVt5HJyVkNSdFtly3QiCTbkUUNnpLV
jUOGYZJewQGCevjAptNstmQCqyA1Qs3DpbxQFQHa9mXgENCKb9Jn6IdaoOEWnSty
8wP1BNomjCRuxEutzIudCs4W1om/cAQv2MZ9vXJRJcML4UIpq8459YPXJ9N8vSCO
qwirIngLw4qH9IT9TWIZmfiiks803e8QhHa9t8NZGGqtSWtCNmdQlT5rgSI+BMI5
7Wuy2KRueGbhQiYkWYfy++4N5KIWV/vJSYNT0Td6rj8cuZjvFTFg7/dVoPfjsHS7
7XQNiNVR/0RoQG3klOWxF9ZKc5AeDtCMk7bkb3F9ygJg9stSyGN8Z2QJfMcD+AA3
kVQhz5cxq4eay8S7O0RB3Ji+YwlmOUpeYJMsZwJE7P9LalbU7T74jM/YgnYouK/z
IysSyQwfPGysTL8ND9Pfu9mx6gY1BwqQnn4QTJVJzBMJPorRNFAiLtKrsO0/3d5K
q8gLLrRkWuonibZcIqwbnAxlkDYiC/0/nGcvnldSUNBoqbcYtqOxxnv1GR4kHoeA
d/gVzj261ZehBNBW76hbQzRKkbbEjRleUYaKwy72xyh+hBFBTMBgShz08K6ethQJ
xoftT8awFJW9NIMEf87wKLNq1dl3rRcwdU1nVFEQCrofNLVzLXzVwU9XY5fXZlk9
BvTuzg8sA4YqrXIm5gam5CKwQARK89DO8Jy5XxuuAPyajWy06dMlmziS8gEcKoqz
YWWC4UMS9MdKmSh062TuU74qFc1bbWUxl5fF5FZmrl0tteJRiC7I1sCHSgjTqeJe
CBftALyRlDXIPwho80mp288hvrjHZdRTe9Wjuc1/fk79SjOXmTtsWTRr+1T5j6Ij
xtmYAs//8II6K5TYPWTqjWaHMgmtGe1Qehv5Hv++/GkgJycHnFpUfwsPuY+lSKYP
uLhCNBLcfWzhvXoDt2wt0YU6JiW4AnrAvBgi898y6/6LSUTN0JmTTYhkjUz8aKMz
TB4ByPg/BbplIbByKskmt+dvu2HaZobpdlszBK8DRsW6IgHHITgbmC0gfBxcVKzl
KES4Pxo6+Boq9+ahveRmTwIf7Z+JztP9xqAbS+V5Ck+v6a4t4HzuGjAb6Ef1xfUz
GsVoKxtK3OyNgxLJP6tMRV+a3NV6NJenI7aUtcR7WrGqrB+F+pfSswvXWzxM0QnR
AqOo+S+vWwdo46NhoUJEIiRJxj7CtJoN1x/+4WzzaO5ykVHFN8pE2dPq2UdEi2JJ
4MzOXnAbkEs3mEMGMDjWiOKhyNacxkSkPdoK2TGAIZzgM3DOHe9+OvLvD98AetvR
RhcQuPaRu6/lDqeC9kWXv7qbdo2ZgAwnsrYe5WUriqqYGNhfBGrG//43HHEyycxt
YRy7gWJP8KtzEWbKgx24mR2L/+uvQdA0zxIAIqp1KF8AdUHFRP/Pa6BxIXgzp+U3
Z0k7J04hBHxtdosm53P8FC+EXwcfK9u3kkaoii3cK1lhUXmvmUwkQ/TRLSg0XPpI
qE8U5qGxnt1UOMXZ26k9nDvbxPvkiqTgK2wnT+8ZJvBqnUZDJniblMlXSaLEDvz4
`protect END_PROTECTED
