`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jw/pQ+iRDcGEJPVyRbMn9yNjmRatX5t8VYY46c/yB3Nh8VBZf8CutsedeZstEI9D
2EuCiEJRwrqhJhMzXp4M7ElcB3VhSoLIS/V2c4GJx66ecnkopS8cmktxlNazi9hd
WIeAf7F87KPRW+NyLz8R3XP0u7KT4m5uzga70gQaKITy6YgOtY4zmbG63DMvNke5
SH3ebAnteory9KVVVwHhqzP0JU5Caqt/Cax8Wbi3iY6aV0do3PjmrKfTxWcgauDG
yFJfRzpLJbMmB0UZ7zlJJGCtOeT/VN9DVPJeezMkk2s=
`protect END_PROTECTED
