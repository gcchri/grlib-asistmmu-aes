`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DBy9wPfGGnelDvXgucDlOgm0GGC+JSTQHjEeSdZvc0S4o1Z3XdGgaD/dnTTfovdj
lSsI/5qtLhyMur6bgOVvvmw2UOTjIUK7xQ/P4XPwrCAFSzL6NlI0FLabPbhVq5aj
q03/DRvaTBSj+TO/XbCGoj6W8Ix6zbCFvWwVP/qYeOSzAC1B1oPjguCjBOdLLMd/
L7cm4qObNt++urADH2GjRv8O/1OiD6tGx7JccskjeI7SWXLgQVF7SOtJDGwco4Cw
W5rMuuUnikMsdZp0XyhxTm79aVwWQAhG5mm8XOVW7q7OmwctqdBEo8bSyiWWd1WW
IEfMHwSlJ0bJXWKs0o/NW0Qyz5TD8BuJ0YGXnTm9fJy6epF+e/hMCypHGpt5xfeF
cfTuWyfe4lqXVxOgr0hH2p9yJVVEerQulYE8Xr2WJMWLhUYsIL11Nk5HphU8sgmd
r+UfiTFdK8WNO6+cezLzBnPGv0KT6VL/vvIsQmuTEqHJ3cON1DNLJJjbTSS1m4Hj
jqnbXX8tsFCljzzn5QQfjOLDGcLIy3GoPlVsyHxiR33wZgDXaV3hqbJLT3JC9YPK
7GJTOFt7MLPt18IjJNf7vhsYBgnPtFSFZq6YHEwdNMJaUdtYP8Rv1KQOK7iPtiYW
`protect END_PROTECTED
