`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GwkX2gMwa2ZmzgvlJSxlEBFqgUhUSFv3GgdG6iWb4rL0dpumBVKkgHErgJ24GHYN
Jufo4rD6KidOTR1s6tRDdE7ANtzAKNXyGh6h4kjA7s6Q9pl6icuKCxTxngDeMpvS
V5ZlfwgRjUtAWdFNzyycai2nWtaRijkvHyFOukAX5l9sLniLCjkhrK7Wq4MGVYzO
Tzdt1TAsTmBFW80Is406U6fDjxbMd945cWBwyuIIrpJzLL0SoVU4OaLQxjMgs8uS
xfE4nM9VMuip10v6h/Fr41nJwlrsPOzxhRrL3bz8AYhKGmLqqtEOnQ0eI7tJoyxb
D9icJFpT3rVvAnHtmVH7okVKW63hrH28kA0IDSj9eIwP2qdXF8mVT/27gtWtnyop
6eBBt69nTn8YYPX8DYMEyYcVAD/V3fikZB2EHqcDC5ur2Cwd1X+Lc2X8trokUXfn
IlIfsB9zvtijNUel0ZAqvUaZcDvXIRuxlcW1bgDeNQVcGRHl9359URocdorbOXJ9
QjIrr1oHPqu5MaXcphHLEeZU1dHIteAJJCgdRgiDzkoAJCtrs8sZ3kAAwbXt9p81
WJZFAPhCTn1rG6K5V1UAeJ3t26IHOc3ioXoNmLJ6euVz/lJ70XVE+flt1q3GIR2o
5/TEgPjQKm+0JQCot/M3xBus+e3FBHsp7IB5rz7prWJD9TzpTaqPqSaMv4omuxIX
RaxyUd1JZJvNhONm45YAwJkQZ/ZFVvq0i3pkunoG4V9v8x/SZUAIOPeKwcp5vQ6b
C4BqHUwUIESR1SzQgvS2aEPxsrgA2+G2xfYVKwEKBKNLE7i8qPMWPPvUCwbtbtyQ
`protect END_PROTECTED
