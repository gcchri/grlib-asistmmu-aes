`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/u5UzFM65rNR2fKUxNL6M/otQ3uHL4AcLPlLsrb0vhz2q1LcDpP+hOxpCmjjwi9A
9OszZY5HwZAPc47QK7q3BxZJJgptBi6lE0qkbCtRHjvdxjARyJooEUsbpXqrOONw
4ZfkKq1dzzX2pHVopWcmZp1xhFCghmFvviWqWoHm13Hp9CSJ+zVd3GwLeMK2PZS3
YJ6Rt6b7VsHevsmMk/z070bbBrdCiOyPupym1Fz+f79ubg57e5sISqyaA/q2wj1z
YiXL09F+kU1PnhYaQ8WVjIsjf3uF9aiVzwlvijPdH6PgMd7qGu/UMwzStTP2K4i5
C1Do0tTiKUXBm8JiEj7rNCvvVcn01zpCH1c9vustYviY9xEdVc7fR3ZNeCcsGnXm
dNaUTSg9dqNUFlDiiKfGyGE5H6Zm/lsI6Y/WUeyuYelFMlLoO4jj39Apu4IHV8U1
5AIC94wuo7iOLuP8KxHlGoxAVjW8N5ZDThvG7alKPxdWdPxCZW3N/MsymkBA0a5G
qDz6iuSA9+Mdo4dkOighQRVTjBmZezCMjnlP9pcMn3m7VgN2rnGiXJ0fn64VVHFl
DexsN/rTI5DxE95Z8hHnHMSjhr3Of44WCelwmHY1LHI=
`protect END_PROTECTED
