`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tZAfwDp4NhocOpZ60zSyOTcfe6sR+9+ZzqbjRK2y45HQpxT3k4FrgvyYDqYkhj1K
2pWNvsQHOTAR3jUMHcqWuezfheYhkdgTf1EzR6uIoCZu3EGFyM/iUej/V4e1xbkZ
jYWISGGRxD0L0T4sAv8b5JCp+v+Lo+L/mWXkXGNEkZfu2YMMyWOxOz819rVVSl6K
cQF5leNG+cDis7PK0OmApA/TUm+ZxnJ5qNOMD9tCbERCy8q7cPnC9k+kUiDuPRUY
od1w786Nav19n6pbk2pQ3bXh+Yt2HxSkZZZZKd7iby2v7eYrerUFOrwHY3U7nNeU
Y3kezw+EXpaZlsjZMJqWAVLFbbiuv48s9wDGVC1PTH+QOHnq0hErNoTyTcpxPr/N
mT2RZDkOj3Uiv9uZTBJOPbaJBGY1qlYsUr5KFs99j6CC9UTTDiPtRpkgUy/ucl+n
JlPpxahnZabJJ2jsWPFfFz5BqO++d2O5k0zJKWOG2gPoabvolFy9HBccubBis0AH
/J3trcu+vxncPL6qTTCJEK53GOVn7kQiffJvsPoDPsw=
`protect END_PROTECTED
