`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ily1OyPVQpqbfaZZJsfFt7gX4vx1at58M2XtXr1D/8C1eMAAWZGIDP5uksPRlIit
F2CyQNGaEbVU90lSNTXyI2OjReGaah4AuNAR3aCLdRoNZgaOcs+mtLRLAVdyLpVD
7TvNYvd3Fe5FYY6aHjbueX2Y+6zjCmj1fFTUQ6hOlQB9/XHXIOz0d9x5JWqIOx1a
NSf8xDJpYLHWrlk88DHTqWMa16dL7Mp5U1jsYnNx5jaC1C0jvvhok/8Wfb3X5MYS
wFCCpWxdg0HqKsVDFic5pScbvEBhvTqo2akNYwE28ffq2R+VL92m8TDgT+yptKKG
wdviIrjJObqffHgVrCONF6IPyRqwhF3RtAIuFBiDSDTO16XInU7nqKNsLWNEmimQ
Nq9vU8bwJB9HogPj+zgnKRaklBdVZ6LLfSvSS89wSfQACVcoGNDkVYD/f8Zb+mvL
a9qRK/XQuJY4FQbEK1gjDQ==
`protect END_PROTECTED
