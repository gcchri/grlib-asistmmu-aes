`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+bMAP0aokv0uG/yXAj0GE0jYHpdFqy114QHbHEjMkVGl9/p4cg1pKrg12kDbfHx
zdc8PJFObBLWYhd2OiWU5NE0dmb8UbaGCy5BpNH/+WsDHzmn3pusRrrBFzXjdg8S
K+LT1HsedS/jnH30XGqwkEC9UJ5hbZbk0k1gzYessYk2i5Z8qKoPpW1LJE+uUSUA
1Yvdll5hFS/3gkyyTflAHW+VWrZvE1aNSkNXVERKkAtfuAj5tzbrUwsNHKM1rs4U
EeGPSrcnHzky1CzRhcruxvcmFs6oJnfwh6C4s/aea2KsRwa1ahZl7O/pb3awWs98
Lq2JfCei0ORicF0XW64MswTQCtehmWgQSE9CvVulIhjBX8FAU67nLO2bxFE1Jl+P
4jyP27L64f82+Xx/NjT7WS1yjA9Y0e3VdJrZL7HAAJr6/aBD+Ic8AzdmJ0zGZohR
A31MfHrtaPOGJC+x59uGpcWtHVwoFahOmC/tGWp4VPxu/2q1BCUWGgeoGOekiKfl
r6VR2Hx0Bkl+VEXXTWJhpCZgKtWObqv3ZlvckhIiEc3MERzn+JlEIoLEUOieWdkN
vqX32L8qu+HlOti+X6lhoNFkpIJb3jRoLOY0q+8GVcCgQppu77KhNLaCXDGBfBAo
FWbXHMGGVvoqIUs8E0Ux/Bu14HepV+bx+2GxWfjBeNip4AgIWjVzoZpBdrm03xmR
T2oIqF6ZOmZ45/LbX/EZv9AFpBYC9XFKGqCPVTEzDBE3sVDhK6DVOXcmhD2so/0x
iJjCpH6oh3yyNV4SJTz64nTbAXgmEoS5anYDCH1zBQG8sb+nBK0t61qJLWElLbgy
XZBtPe2ni4OIbCjTUQIsVPcTT7ZDR92EH8ETc5X4U9G+TCY+xx4fw4mdRuJQwY4U
8wfAZ5a4yW8iUe1MRiIfC06A86PF7LKwhbNbg7w6SIqzYEfnJC/yjO+K3Vguzlpe
b/UhOZ+1d3ygncGZmuxGvj/57y12sCivVBTOWGExtOrnt3cSh5yTsLDDWGPI7gz9
ocj6NQLbR6PPuKzTnVN9p1gZ03SR0C6IDi2OAvz83702FITiDo+m+/WRE43GxMp8
+ULH7Dz6R9DUmwcdDGtyGA9QLD3F8VWdyrrCpTF4ViFkFXEgxrUUpPxJ/lgXeU8T
7eu9yVarpz8UJnsywbRR4N+AbAntn1sSUzNngrxh+sCqNcx2eVlFNa3EHtQMgluN
qpAIzKbfpHDC8fCJls7S/9p83J2h4XUJpkIjWu6lLXKxTpDn6aqdJcl7mEJlOX6e
1GEFTgyIPJE8vbuwMVZkWks80sxU0nnxrXMm9xH5M6JHH3eBjnrVMMNX5weChyM4
3BU3H84AnyWPlVXg9AN5hyR70ClWqfWmD2fxN8nPhUsPpCbfjgor10TNiLZYlbOM
yym4+UW+zn+RdiU52QpSraflYBkYK3SHB+FHFK1VKz0katVxlw9QigC/VwMMqOCL
kkgZy76CmtT3iMAiN9dwf9xM+3scJoz9aG3xTTj8hno8SnSj7IqETEcJTIqPynt+
nr/KsjVyOpienkOoqtf5CPlmtwkmEfOdq9D02QQt7o5nTzCyH3vb79Xx0Eav2Y7o
UzmYWamGw/ndwP3Hs0TgmmESNJYsnwVUubf5nJ/t8pkkuGD4uc7M0wx2Z1fTUrZQ
Y2ej6GXkKJyQTRtBmdNDAjxsfygt+lQ8lXdg91lWEZo2vf3Syyipv2wGovXzxKX9
WkOPO7XoI0QslVF3Eu2p8mDfeCCO9l0YBDR/pGLlHcxRUi9RCg2fV+yDB6X6p6r4
X7QwFY4NazXalT9cocShM9J4cz/n7a07s/lSQDtl9oqQFGKW5aISSXMQOguoJc6S
TIp2G59ANBXo8Wg1W/ISmJtZdjVOojLA4NSU6+WuUGK1Hy8AGaPieVINCVDHUh0g
dmww/weZE2rzItugQMaQqGHk2MCFVGIEozwOzi/7jpn1F4SmHovYK0vaQzT3BQQA
ryWMBOYHVrsbWAtLUZBuvfMjj+RwS7/qYZQLSB7IaynTMtXSWbj4s/3JZtoUlWUg
BkLFeE4gHjcvHOxWn5FsQqQtL7/yiCn5ltkRmmqAg4hXJ60ZjjDFh10XnYqBUYMB
sks7SnmRbR51yhs7NFBvElnqC3xZCgpSQh2B0gwU9FDxNITC3EsTiq4HbLsrnq68
SAKgKIv9VUldOoRTt8MR6I5D197aZbUXF0aQ3Rc/iOaWWa/BJplzPAlk8h4ZGC7C
gJjPYHwSfVYCf4PT2G42uMhMJKmxvTcGyr91U3AE/5/X10LvG/qgMHFGY3vAHjLJ
blP0NqbrhtXl6re9GF7Lszzok3JcTH9lbEPQo+VEUgj1O0qcFB5gozqUAb+haJGK
FEa+E0zMYXTuXH1LxmIQABnyfs6+lHgg0onGsYBfGiKmFGFr+pOUOC7e1HsLNjuB
wt68vIh++bc34ZP/yjSFINcUfKOyGB7VVzIDf8A3kw12vtgkHvRRwHbjwoRexMTU
6bXJwXlze3waL9g2VJZeEJ2k+zDFxWRGu26mQ5yrc/cbbT+IDNpXLS+eKMtQwjVD
fil4WvBNbXG3v/xTqoCdite9aCRwRIST4Agvh2KYLrxwdGenkD+t1egIsXW/NKmc
3P2NZR+tgO5Wetlm7QLTTXNNDILkAf42wanUGQrQ18bkH8zdkSxCc8y5Y6S9t565
Tm0LqHYWeuNjnrYSTc0ObHkUNs7mZY/ybGURmdbg0FQV2XzZKZmlY3vbIfbOAy95
bskXk1xQBlP3QqS9U680ESyhUNuMIzik8hfO0CC0pvnMJ9OPKewGMnjbiQycvDwO
QbmBSolJcNmWJN86g//nrVf6kU4ANfMzWLRz6s6uKLePEepFMygIKJP84aj+fi1K
MAWzA75Pq2AiNzcucopul62Ogce1RY0HIR5GJjGj+MvJFsf/DGG3B8ic4EvHPnbB
s22LbOMupIjz53lmrA3XOP8eQ0Il9ds9TjyBhcffrA5+Rw/MyerANei6klSto0qb
xe5NXwFf78wCQ+8wmwDDhPOGTnIyNeBep/R2NmymxjDsJxQ7TE/C70KBmUvuoP5/
Y78zZc1VlhQF4rf3AzDCQMMEMmtqEYhWt6r/1SuO6DYR7y/gf063++k3/C+rNfWx
pNTTc0qQbCBpwRjtINibTF2eJlfOcXryhO4qFkpIMbCef1RRMbRbE8fUHlOt8yn0
Pnp1IjoPBfbcMnd90QmYAHyiP2nYDXSvdVGRoYH6Mey0OX5tncHuC5Znddl/f+d1
n8zGPIkvO//rmL1dmRzs8CmpPeD3yPi6loVa+vEgeR7MmO+jNPh3VeAuXQe6Bqna
X3KkbjwMh9+n2TTtyP+dTm9642+uuzPCuiFY3kToKzdV5oZL5pGHmnDMDGj4J1ur
dEgTQQsxSj880kiF/GPKfsEhfnT/Wohn+IEO9P16fDz57ubndAZwQRzzP/A/OhbE
b8w//FOGLGgMePycJ0BPEdmANgSKp5Y2UpYLDxatxPlcUYA4dAxZrv2pAiI7PLg9
jLcHoh/N5pfELu96b+eIzizqaU9UyiP9cnv89efsC9iFqS+HK4M1g6y+hZ73ql3E
qAOGVLSmVJWHS5Lf68Q21R8aXNDy8MSzoBUohMLZ/l56OmUPQpHsJtjDc4Ex9ie8
dRiFD8eoL8krd+ZtcPg6UeoQAb1KXQ6VPsZ2U6BY54nTEDW1F7ylBLKTy5z7vNB8
QVXyKD0L8UisVs9O4EYexxaNN/cA0E7tLeMvWtHzgxusxV34Xsy7fSdJRq7wGyq5
daudfmynA1BadX27T1h1sXGjcBNwUczRJ3pLnVMpFiMpvkyWqB4AIfQtDe69NzKt
gbnZ9Mv+KrKitV6XToVduNZ4b9Qu8dfuAyuazD0Nqbg6WcJjbOfscOEory1bIhg8
eEME2uINXmfAqzFNHgK8pKRZf46TsPmC3qABIljbJoYAKy0KAsqh8r2o4gY/OpS9
pRYrrJo/JsV92QCVXT9vp1QajBLTcDO0jlNNh8Hdw+UWSBo+LecKf7l+QIsUtyav
6/0TVzgI1oTbHzJCBeqU74jjLS83rBkwYX1WuXC+COardMq8/pLUIPu7zJ8tclPO
fm39/tuKEb9MtOOC6HZ7XzGPPJJc2dvQjFLYIp2G5QVDm4AygHLLWwxKui9T7dme
LtEyUo8sCWTJYstgREsny7ZbWSu/FdI/Msi1+EAyCcGLurVeD27jHQhlHD7RagM5
IlIJMrdlQvosXEH5D/rotaFuRL1uOnXcgOpK10lrKiizSSiTGIokKLKbzVdX9A//
D0+QK5ecTmLIhp5jMD4H71rBvUZRBpCRFe8nSrYWLqsflRdZ//EFPOXq4KJ0WsPs
4lfQoid4kK3gN3ptUcsgl2yj5+yRhe9ebxTtwAxUxajnegYUH56L/dVteaPbcD+u
lGp0SdqgItUT0qUz3bQyufyBchrNRxfgOMegvc/8h5KqTXjsGVgS4yvC73rCfLDs
bXHQJ6zPt/mZcO89aflNCFz1YUowkzOw5cvlrTBv5/QV/G3QNle7o9xfbm87U0Yx
JP6h1eEBwnLFRHYTB25mHnNZJ2ZQqixbKvER82nvXjFnLuxak7OEWl9tM8IAMmps
aC/epDjaWMJgnG5g6seUZU7Lyy+kvMx0mJacDGmx8jaNRwydwN/rt6DiPXWqdpRB
kEltfnfFeNMR42gXocHVrbw6nVYdHdwx50mBoADyHllhOHZJzK9Z6GuFKyZLtsrl
GMsZ3hplquhvM0Jyq5MH5ikt203rqS7x9dzTsv5QLRyHRXCZNTBJd8TNhDoYcPrb
l3XQHO73vAKNonLu+5g4Mi+OxlmYYzdvlokysBmvuKXaAsNvV8OLOXQ2DebNyKQI
lrLvFxBigWGVynSixazUHXFXVaMnF5cZFMMY+UgVjlkWVSwDPMFQRZBBrIgVYA8J
LFkhz0skS/MZXkpoyUFXdKFL1aiuLuHKhnf3f0uTH1Q3uf4idS+sOEUsNrOVciXh
6qxH78cKgvxYJmonI7QtLGw4PvA6RMaB4icwkxGKtYMtBMWJC3XcDtoutR2LCCcL
6NftPmncMXh6AYj372oVnJiVSl+1h5FFXSuHDto9Rf6M1xm0xHh200XzPYjXiQ0P
gNMjjLXFubClh/KZqY3Iq8iHJqqCwalY68daYwvVqkQRfZntlvjCPD97WWDlNfqa
EqBxOnvoivTHgrOelmbRYvnFr3Eejq2xmwKFNp+b94k4USJqm83z0SPg5LYP7cdV
BBbbCYrdkF26KeFYP5pQrvojEGcoBzDGpVA3VBtGhcImychbKhZerC9vd/XoChxF
mfXdlEgFrkuuLxThMotp737/rHB11e97iKIz5LKbuV9WsaBDtBz+hfVWICOVtnzz
fp3To6iU2XBJXNPlYKSh6kNCXCbVBhCywkwuRI50BaxZpexd3d0/AA4TRSQDtOE/
SRpfbcd0hTjS62u7202pgG80jNEpc7GbmcLDqAYb9kSHcQ0yyGPaLGRsssXbNsXy
814Er2TrgUbQicXDgSVO1BfrT+VcYn021/SwUu73BCxcj3dPAVdfvwVMCGbTWaLQ
T9UN5kHspjRArOzEn6bUtR6U8MkTVhKeD2YONcZPZ2fFKFhfEaJjo43fGgMDY9O/
2WpVU13pzRVGfwWM8NpNZ/NPiVBtCwVuHYoOD45qTppp8J8ZeWM3UucoR2M49EnO
8OFTXm1oho0oURKPmPMZS4loPPDJO+E8IZE3o+nf9HAy6+kh90SfUY+zgsESfwaP
NNajuqdrr7Cvw21yDqWCtqLPaWjBotXhbhjnGV9AZBQQK9NwEHijr+Xx/YuGCM++
PDGfshjKQEWlCXs9VZIEYRUlVDMvlA/p4yPR/CSzNCtcQMuMxRQFOqhmr8iS4MmS
LI1UQfJz1LmNOxOlM9UZTjuTqY46A+pcqPQ+GovwA2YpfY86bLWIMPq3cH6PNEDz
IePENOqMoUuQtb+JIa7ey+cGgV1/FH7rJZpYEBrUj0lptMKMNKbybL7Wf/ojA4VS
tnWttZhssPzWW3RlvF6mqVEu9Wjb7gmH7xIQKwpoGLt09EkUr721xSOcoZHIVEAr
e5FfEBobMNoU5wAQqZBcgGUqrraYWC+ue2QE9/36BhNd5h2eQZbD2s/0VqqbGKRJ
XM+9dg3pl1yR92aXD6Odm3yK/9awI/SIGEfWwxOBVFFRFWFQNwhtmSPdG17byJ9w
OhCHsXJwuy7WFOILpGsiSIgAS+fVBHaG/ffFNHO9/2J5Ypc1ZYLl3E1daBLpRhjF
Aotz2ceHnBi90VtDqhQ/CELTw1dg7KICN0fmu4Kh8TC9XTT+9cgjEg6xTw/GvPAl
3Qh4FlbuoZdIemIJVd4OKmgsa5R3SupPCmLqtBAWTOTyhsV4CVYQvGTVxJZ2XbnH
3TZC5DAwbNy8B4HqEoIE0NiCQXo+AZM7+GgE/G8nGADkC4px5qyWJ3FNXikNeYPn
mclYglvw8x+nafducAHyn9UPZI2/G2gmkYu+NYkvOf3tESikwSNEepqRAKuT8hkH
bhCfkVa3R17aiEim8sPeUjZp+QCEiyGSLnaRPcXEBgN1I8kzHFbc3/1GTKSDkP9w
ZOcFPuJXVLHz6zub5oI2efKt99QZR9a3HX56AVHxyIWUlt9zoOra450JPUvNYWl6
6wHNKczDL3bNDZJEbPRMUSgwNWLW6lZ18e8mxnxBzQANai4STJB2Ux+JWmonX20p
2qK7PIMegYeD1SEafSr1W4o9uq2jBxnco3f6CvCZwAxjRglxCYmJhhQLtUCvwy2Y
r4nJLnH5NVWvqbqtINjXvg7av5JBZ3VY2CiJY9MykHl0oL5DrCF9Fu2ULbgLNuPj
Zw0PrugBvEigOYeRkpZvO+nJiO1MPFbNbp0HgvxudWdzJnR2SJ0Un5uFmx6wbn0l
NIi4XtFcKd7nXTXqhwQkXB6aBB+Ik6/556axipZcKDz1zE7GNnrdNPWoSs169aJC
V62zJy/hUyoP0jMkeCUnNi+/JbXmyIZtPthtid5La23U/cF0LyZNdPOneiPI3PTR
S+comh7qJD4s7pdhFaC4Q1+A1kvtrqcmVMxnfvDwLwTGL7uFttypUTFdjSq7R57F
fjf3NE4QWxahZjHgjmM/SSwMESCxtadbhRaHLxUzTFIJ20UOuV1/lFb26Hb+53c6
zJRd39wZF0Uk0ZkpZdJKHVj8DgUyM9xjBghNaSip78MKy5C2/u7D+Bxs8M6Iv/mT
aIvm8dW7tRWI1SrMfKcyBwZv7+kpmNcQSIf7aRG/mUJNBV9coellTwNr+P6Ww4+G
K6dtRDv+T0jfCkilm49Esp1pGQmhhlU23LaIXDjjbITl7oB+lSLP2tFcrAaKQWBJ
vYju04wXd3B5yLl97G0SZyLFxWuHzIRwaFM4K5w2fRoMiZ5TgDvt9G7Wj0xwCy8I
K1F9RBY696Y9J09rnYAT/DajPc6SbRFt06vb9ln2o0sb64t2qiUwSE3b77yV8/Bp
jIjG8d5ujcZ2bvj4OKGKLCF797faB16qOVHamkg8MJmap1uS1jGSpLMpjk7SwMZU
DocO7dVVMDYhHLI/TJADcuYbyD1bJCBmL0q8Lp/mfsvlZDmJsV4N/Ie9cwJH2zz5
6P6eVzKvyCzRNb404XqzEFJBtatGRrCpC2wA6mW4X9kodiwiJFlDObzBQSgrsr+D
Y0r8AxYNSd1VpNC/mrnwLQxynp/1b3rKa7PjHImHQl84Xg7tUgNx5TgkyIEQP2pp
aBTfpLBr3mK7odDf6L3YThcQcGeauLsCUiMspyYxBMraR3zCYHbx3s+tmaV6lMVU
cgDSmPJo7Dkst6dSFPWG+uDaNRpIFFvj8ZCT9titwzyfmLr55t7fPYfdI0sInnhI
gHJ4RlxLK2Tw4++CD1YeeZ1stIWVBuf9tXz2mtqYGSN+E+jgEJa1s3WD/8+lj0R5
qwLVGaDKMh/FPlQdpg5gdjxNxsg7cxDUsqN4khcAXv3V+BsZh8Y7ZWE88BIQRlii
pnRBHmKNQg+k9tFcvuLKeruN9MCBBUe7ZyATJ6aTlv4MLa7wZxrX+2l6Bw0xyPIl
TIWJR7jG/F8QyLYo7PLSCeROv35lJSfc0Z7Fec24DmdVaojDvN8lNhUSToWFRjST
NvCgNK6jyxvN4Sv8ltxrQ43UFcSkgukuWrYt1oSR/pSvtSX070ST38f45fvYZNBq
32UuX6frSLOHONngZ/qgvf/S45CFDIrEjrn6bb9yrtuERljVwywNsi4TknqciQvI
ido//KRcl4O6n7fV62zc5lVFthIi/BF30Ci+i3hR+rX5ph1jwMJ6dkMVgK+yQQv4
xBdMu0NJrgnMifUhcV15kQRSoUbUwYCpjCEFiPCYgJLWaASHh7O7y+6jx3ULAR+D
jYEOFL5o3FhKW/uEmRg7h6bNGRiHDjmr5Ny0lvtXYlit0WhzLw5dmyyWvVyru5Ft
uSlKpe8r0frUsQwD3qX6ME7gZpt+5Kmyio1kZkkQ9eg4st8k5VonatrjWeN25RmH
3tmY58ZqDU+LA4Nq+h72DpRx392Gv1IWOdGOuEpsN0ej4+XX9fKKCpOTanD6lRG2
2R7kSPVmQU14Yqfk7zPRSDW6ERPJyeh7Sjy5dgmcqObXHOebz/aSua5MKR3MiZK8
xhGjbXBDJXYGHTwZow4+nGXbT5+MdIeCnNfMlqowOlM4F0vsscQ+valyvZc209T/
nDZ+5t3KR75gEOcjjoJSTF3FdJ+My71crm02rjnzR5NzTdNGxfgd2GpNaZBTVzCk
MwJTM+RKXoyAOra1hFUK/10Y7h0xbEc8qgYUq3Leo3v1RDwW8itAD0UvTSJJWZnV
X1MQL1EHWB3lmWYPFCOZ5ykeGHbpHJFVq55h6wE0DMA3tHN2LnzXb+KRZTO56rdo
MkWhl8lqvVFSKNmseRuI+EV29F725LILTJPTDC+zYtsfesFKlntnMW7X/B3YRKip
iVgTSTCbpvXjyf5qmKSj+K7X0o1mwdgjSWt6OKb9uzikAr46rKAoVNZ4ZHzUoMzP
dSBLZgqnLBnlLUEAC9KHd0nL0MKGJ7UpM0ye5AkQjKXgGhz54o+FMP5BtzaZe0TA
97yj1hlQn8NzFziozWwmojOZluE0Yo0ZBH+70kRuTqGg5N1PTxFWSKPyr+PLemXB
MFpEVGob/wHJZSxgc7jDC42Ino7nKCdYqZJluo4pJv1Dl+ElYgvmu4d3AyY/ykQJ
QmXiiuhioOwBJT9ngo68RqIWV1VsgAc2YhFo2fXmCJf4K+WKwEnkgt45vS+r62X3
IG34jH/8vqcIVAaj20HOhvofcZGv2s+cFKPqNV2a4eJFb96YrQe0kZS5emhWURmI
akFm1IO9QZV0wIl0YIv8ZDEmsm/u9ymHMLV70gocfSXs3iRLYW1cw02/yXUo4n2j
CGsnevFRNzaQIYtspAMP2VVpXEv2TC8oqSZJJgl5j1/LzMqvk+bX+CTDtqtT3WBV
BjUf2c0Qp+Fs3SwKNcGdBBvnB2Z636zLEnRaY4OkfZFbcRDznABSQ4SvakFzlC/7
Eis4Hu61ME1UMECA3+dw56cJ01Im0dAMYi9cRI/0AhOGKavU4p2Dm/vrCxrnzC2v
A+zAjLOT54USala7m+5aqxn2WbWKDo8eDckmhHh7XLctrGGEKqPKrgMDS14Io/BF
ibPiEAXgi6Z7iBZf6mxLXahHgZTQNxHXNIykj6pL/D+HDTCOR6xiUtiMqrmoT4Ym
OnpD6Gnj5cC11972Ezsq75Rym/4jmY236sYFSR/rM6kHi0HVi0kMGO3sxXUMrvSN
QzabrDnijNdlXojT68fSUg2vxYAkcqYjvp62aqzVXVUjGviRZuVns/gIrmVEt7PD
4kwyyLqT4Kjzq7M+49sG+oQ3TanpPmq1hoMU944Mv/3GYmzq8+M7UmFjqlb03N/K
pX4cDi1QdTBjmmPjYVJ1yi414zr9BvsbtyZ1J9W6uraqzGZw83uNFPunwie72Mxw
eUJioypNQxlXhIx/z9XG3Z61e+kH63MAqeBQtTjxx7ilDRM5RyV4TLlJzyfoaqIt
JKceXLJMqViKWkPe3ThttnsKI7c4BUOwLYa5SupwVJzZppztg3VE/T+jZ9b/j2Rn
/oUhGgY2776NPk2lK0UPDEdaoVqSxUwxLab85/SYx+C11E8HS7ZAL1zQ01QlL3Fu
LQ9A1NjzggAw4uF7dZPKlmsXAtNW5zdIKMtRUQCVulLMudZvNmtolDaSY23RWepA
VEeDUOuejcQM002NAllMI8H0pseIKLRd579Z4X6XuV8vqstcPe7NWDIhVWhoHgw0
4s0gWoMonv5vl7haWimZl3aoyRCSYRkTBRs7OvoAxSkr6orf9Ai5TunvD4pKKAGh
rxkPXE8yehm1Arcch2FsNil/o+yPL9pWPLXWOZvG3lQaL4sQ4bjkdIIhKVnZq4nP
Bg8RLX0eVpK1bo+voKkGAGNRkvFMsjDSK+IMatRQJ62579/YN44idNVUjg7zMpIU
SDmlSooDHQ9iP08/xLnRIGRd1uWH9HYFtjBW+uAJClV4vgjGDaMZ1xWhNVNSYCyh
ILFL40TWez7y/R49j/Zd/7rp9n1y4MhsAXAXKXHwj8QEg1cd2zMxrqT5b/OHLCza
u/0QVxOd+R0nNHIbkPpsIN64F8clnAID0OtGkCK5jawhEh/lgJN49Kq9MMAFLT2H
6hunCphQaJNiOhZr+ablJa/vzBw15J7sVzc7KxHVJjCjiNXo/BEE1QhDyoXwI0Y3
7cSe8/L9yBijPLBc5LZB4OKpqFADB1Wm9grwKZ3DonV5+OXb5tar79tJyg3X3gL/
qSFXFt9lAKXBJhgRO3LbBrOy+n40d+SIyiTJCdDUyufQVRaA3hT3xmGxoBEUmoLL
8CXMe8rqpfhtqPFVwPhngNEDpT7LL1yP9Uqts4o1IYqlOOmxSbEGwky914Cwlz4h
oTtYP4VjEJpLg4VXodnC9nFDkS5Z+S5VCkOJLZpDOvxRVnAGITlGHjZdJ5I4OUq+
Fd3Wd1rQHzbe0lyET2Vy8qHSTHaj/iNzIGIA//hV5/X5B1Yp88BTzlQVlwzYn4Eh
VvTcaEbvLdqCLf/kdj6UDYu3SdL3NZv0BKyITcNjHcF37EZpEbtO32PN/RJeVk+R
olMG3m7xQzdWt9fftqmbTSX4TzWaTp1tlyMhLnphUVyptghpzBGAAKQBHJNfTkC8
74jCGYJHPduXkDW+hPcE/JOxhOUJuS/jf6WW2D1ztfJkzAZVFdmJNNH0nBhsHa3Z
sfc97ZWjC3YlvJnnYqTY92ob4REstFCkyyJXiO5sZrDGw3zsd3t1ESi2Cug0f0hP
lkl0IhIThU6Nl9ZIdSkOFdRf7sPDF3wV3cVjDFnG5wBcXo9TOjs9NR/MttZcbEyy
MvHyitIMlSapgusMxh+/raNeQlOZmDHEYvGdq1LUBHAS59wRYAnupw7IHRFFS03S
Dt39Tmt99co5O6dOke89ES2qL/P2Rt4Ku2sD5XLjWPPQQQaGdM4cP0HotLvvADYm
kTXEijTpAsSPaEN4YP/Fiqa4i5hTBkYr4cnMrF4xN0vUxi/YUunqlz3tPJcnDOv9
oIa5pp7uv1t0qMlk0auxIe5+ww4vRXWGrWfwMxTmCMJ80Dv5lcvjH1iykTjcSP4i
uR4dv7WycA7VpXOLd8DgqYw4mBKUcFn4JYrc9BJXyQNzQbx8jWHfDs00cP5JzbmH
Fl1T+8yupNJhDrPQwLENi04xOHDkZzxa025fBNgkNE4HmiG66na8w1fg4w05BkxR
BDTf5zZGdVZkMLZjFX8PWMu2yg/b6hjzTe0SE3CXPCUe2p8yAeXBw6Y2BE6xDegs
J+7fujPtwg1gAZh4q5u6CXkA9AMQh957E6tc2yuuwqYpcPj8zpLBRIdmP752CcSx
+DYeDKsMlBmeLQBcNbIyUSf7U51k3ck8HOP+q4gUQDuxeT+6p8jJ+K/PS/suK2lk
hH4yvjhfZBrUjwht0Nko/oLcMISFLWfYUuHJhDjF1qzCuNh8ga7ilvFtVDHm5tkx
JrIViav6OlBCRvQh7rDqMLxmhGkkvUIzf3SzxC88bDhR6yaGuZ0mLDTNT6VraYLT
qompUx10VkAiuZAKE3pa7z6HP6wnkKkAmQzmSQhxLoEBpTOXLBMGIzs9gUpsFyjP
4UyoKrz55+ucC0k5Wa6ca3FbKL3J7GHNJ4UjDBxOJXQHVgiOTwKlNkbZPP055UMv
MAEJ6Zeb8SHcM/uwABVESxtx2OFrpTDyoFDQDZ+meJPh+IBvSAZVUfgW+J0gHbHg
UmUFnLoDcpx1l1TPC0O3TlY/idWP+696fPg917XcCdRqGVroYTd2kc9rogtTnN7M
PFniM86gO+M5/sbV39n9jXEpIr2Amu+y9BAC0OlFVXaH4kNawbH2FjnP+egHz9Sx
Ho+Y7PmeSX9/wfWa/u3UHrvwDZ6dcTcpz95ZAN3TEQAZHauEtCuNSW7nMjTPvtja
k/tCZguFzv050O89vtvIkBO6ByFjOpVHg5NpKWUe31nocoGcniLphzH9CtewTb42
3sqQX1ryCZ7BtSao0vdJyTKRm0jdzpTbRJXx5OSAaAJelvhdZCxRiItETU9ijn5N
i9zTBJcP8OHm+PWlTsJkBVlCxLf/Xg9rLNcReTFGxEk0/i2wxJhOM2Y+UcgnSbr0
EDeUaep65vd7GxWbT/sNN1SqFUulY7gKZaQUdl3PgD0WyTxT64jW5wZR91ZWtKK6
55pIVx78fPjVc0mtrzjCVFjvmAtrolCis4UV3UOMf3I5COUlAh+YyjcJpU3G+E8K
sfh2iMP/lJnUlW26Bg/GIYP7VFsPYL/q03EMJyqO//rubw23vryWw4I1h9723CN+
xx/OuUA9VDXWLFGn1G+1ijw1Udp/NVFCfEJ9gtBVfOtwqeXLByjsbADJDJa/Lqqa
ckGqzus0QfitAn/MXd/VRGpOzBEn9w9qMr32etoLKxj0V+i9Jye3j15AjKQfb4QS
42nJf7WSMdS/B/5hurhOnbYh3kgxVELOjgHDfZCfbMXchMOL1zGgdiNTB9zzm8Ed
0/m+OT+GD7bhrGlYJqbApr+kKBA93tlQ3KC2eE+/ezWN+eRV05HhDGwdiqbcS1Q9
6ZdzNl2RKPFbVAMLtV1jhaSJY8JltF9t8uA1Vxk/rx3Jx+G9mqjuLRNpJW2OgGV4
DYZzKNwJeM/TbAcrkTLf5AZNrIduWWPe7mGB2c0RtPGoDKCaLt38rHVNtXOkeeSl
H8zhvZTY1lOX/iVF/+0nVg9nAliCrJqy1dIZiWh9QB02ETnuou9+dzGJpNvl8VLE
ActT5ilGBRWqbFtuwo5BLsr9nt3wlXgvS0VY6EE5tIP1zecZhjWvaGE/kodqLfEk
V4xj/jBnYDgITfFKyS+BFQUUc6Gg8yY41CEGo8mx0tcrlo2xo/OSnul1xZpjyOqb
P4x1TXQ+APj8ZEjhUWvZLned9sU4K6Rgtvm/TcDc4HjU0Oj1Uy9YbCaIBMHedfgG
HqEKD4gza2BAH75j1EFMNZorNipFCb1spHLm2w0vvm5qVQh45if5ifmrgJE27IZt
vdVF2j+zZEcAOHZLwMnKoFNxBn7EbrN8pxbaYwXgKzVsLvaAiLIoTfy8WTRy8t3N
Hy2WwOxqag1Em0RTotOrwq7b7u3CCKd0oRHkMibpewAIgxV5ptPyPMS87sa9mEX6
HJ6WfRCQIJibeJQbrqykFXPPjBXpGA0DBJ/aMxUITt2Rvy11dxvEAkWUHpgQMUNP
Ba4ebfPzlFsH0SFgHi3IY/Q0qV2GLAp/VEn/+oSssDOWTLwpB5Klhrahc7VEarK4
T8gEGj9YS9+Fqh8BX3dosnk/XQMWxwu6I+DUBw+jJ06qU2yE8MwMudXEEsmQUqvp
QFWPrxTLmOqEanGzEWxTd9MozgHjagTznc6rSNglqoOKErHB9yaL7X+394Z/Of+R
kpJt5ZNwT3/U4TONsXK4vVA34gGCPlKepaEBKiURM4SYP/c/FOR0KQ38Brka3QaN
97ZYHR2RW0u8XFgvvQde66rrWdm7Ej5gG/VsWZUuiypcZPHunR8YeROOpZK1x2o4
tvKqGrQ/ecT/TEjrhnNWTLKs3XNSG/0i52wg/bxJOarOI/ya3770nTXzwmMEIOKa
5nWkiTVHr9anOH+pAeqLCU7mYDG404f2yg9VP1/ukkXpE6hdQYYwoeS2AM3ePSej
2VEAcrJ2OJkVP62Avo33+DXplrgeTJp2FtqNmJSVwDiv4KnHTa6D2lB5PnTI1WJS
1UXgRZhWw0QXYlzmpkP7F+AHwZOQVPUXpgme/q+Wenuh2erVgY5MV0ujJG9FvG3G
e+MN7TG27QqKtQh/wFuFDCQmLZIj0xplxzF6S4Y8GzYLwzre13m8HIgcPeH/d+vc
CYM/5zi5mFWvykZwZbdTCgZm+o1NoMeBu3Pstp5TkKleB/LnBewrcbF4qpbHWwDa
CwrpsTCEh/E1ieFCMC4bKej7BTMTwNTpOSfzR1tEq+SjeODNtczGCjlcPR22BLTW
7fIMgK/7FGV22VWIdfxUvc5C5S4ok4aTV1+kAKSjSrmZSHYZHcryz9uSzwobD5Os
9RoP9bLUXFBxWIIxDvzqjK2sxhnwP7p7MyxX4zgm20oQiEzGr+gBpt9zldMGVh+r
D9+LT/xIprOwFyS+jCEn48TnT/x98GNlrBw+CgQKnF72V7vTQo8UE5nRIM0QYlKX
agp3u5SqjXYqp5/bVr73ILNW35v+MdrjhYZ90dj6XMSaV2IyZeAmRa76jVxd67l6
KEmagRY/SZrp0pLOTl28wbCK/ar1Qpa8NryZw7SagLWhybNO+8vq7uG0oXofbaHy
AGt1Aa3fcOdm6X9nfWMLPje0nNe6la9U6MAOv6hQYNh316sr2VW9eIiM9OnzhI9o
TR05sNpXNDyqNJpXMrAdDsaxPv9Y5hwEGeAoSox2rN6zeozwjeqr/YT5uLlQCiCd
icI7370SL1YC914/lgQKjtLTo//FNUeymZfcO7zVfsdFJlYzXb2dmtNt+W3PPgeS
5OSWB9b6HNzJs5RAzPf3miF8XszD0OC1TyE0zVkTXt4bbDJ0aThQ57bj/xOhMAVC
v5S7wxCWy0z4T7cRYaMEf2L5Iptc3Gk0vqAQe6InOZbzexjKCiUnFGBoI+TIN4Xf
+KZM1yzAJ9P0LG9LicNVMOUJLYrQonil7gTxuYCV8p6Nwb2Jnv3FseQxRLR+Cl5I
eWhnI+6VpakkCsVTFzBf5KZPLmPkE18ZF0tmbJ8NayfJdn/nd+68i7VWw5ykdwXh
NpeUapu300g5MzvgqymtIfJofia6hvVOB+kKMBAgWoR3rS0e+X/pMHo8CYRUsh4q
DA9yAV5ROw2mSNzsmNP2ht82RC9c/a2UB8o30ilNok4EghgurKDwMnk7vOjt1vMv
tTUqdw3T/zr/YgIPW1wkJyowd5bT5pytIjNUGz0g3j3eG91KnQ48QIHwg6zwMLj5
cnJeIrCW1YCvC+TdNaE7ZqXDGhiZi3fRTj0lZOlMcEDI8gtcpQiYDkOS+DFNUDq6
49qIgEmxQnyBsSSqyRWL0NsGShvzT881fB/0QfDRPpD+iWNZMxI7U7xPwv+enRvj
99p3LtEsAY/jhfTKe9uzYf72WHXwfHsbj1HeGbTGpARyaeWARqh/7ZoJEO7YY9hH
gbaviWwRb7fYihzzpawepuO5xbFkYGbepCTBGJhUOahwLGPOFwd+PeuLWzPKjSyG
x2/EI7xgDR/SQ4zZrW9AmdGgXOr7WRhnPJ/SolGw8nsbTI7YZCfATBoxpt8qEH9X
ph+6/BmXmPKz5WwNPvnUfnZZDzD1GZ0MZq9mQfz0TDD1yAp4a7jcVbkWoOhv+Qt1
kd8LRf47EAl7zm4av+64sofNxPU4JGM8WNUya7i/YC4mOszlAEo//h+RDLdQ+ZCR
eYvgkH9UZsfi5eVGvwdog9cduo6B4on6/DJxpiMareqVQOjOkCi9jQHjwXVub6O0
Lg7NTv+WqNEj3PADq6f+oFOLV8WHR/buIp1beYnDmiCb8BH/bCEtfyazLpQ9tpzX
P/DgFYSc0h8ZmDm+G10PNrRKCz/URqycyJ+5IACamNkTup8s9PqqH6sWt+kgnInf
t/ro7emq20hkfg/jS7LwaM+DiVET/KgeVZklQkEXhVE0sUN/RhlRNGnJEBtnPTyP
QlBKiJai9iFBpn3TwMZDDduurYenExZs7CQEJOdn9sUraZsoowm51yeHVgqlRyot
xXq0T0w6kqXZy9hl8NVX7r8Cs/CvFdZqunHOyX5s1Jfvx4R6aR36MTq88Yf63cDE
V9IX1835XsAICgrl73X4vFpnUZrPJ094TtP+LkJi/z+y2N5w8R6ZXwCWXVCldbTW
IJemLI63wncvcIevLIcf00O9ncrGkXuVD7cKWaRJPhlPzqO/yxi/SDNWsHyd6sZS
00JRXWDvOnaCBTXe1cdXZ7UYu9ESeSN8z9iG83V2/aiMTFdR9PjR4PFqrFGFPLXF
YlvuaBbByGjkWfT0etfFxRRHFjxrvn4gOSltRJwp1C98ff84lr5k+wFsUGrB7Jl8
mSyBldfNWJ7C4Jv3udYN7K+v4kfH0FrdE01JVvdOXk4bcxSYdxFPJ2auQl8uZt6h
b7b5wPAEHnHQPt80dtRqiMl0eqEJV7RclCuRV8A306Qmdi+oh+/ze8ucXbrmAXIk
`protect END_PROTECTED
