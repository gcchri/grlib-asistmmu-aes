`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5rCg7gLSkUqWdgH+Tw5CsJXDmJ2y/7VLLAi8kkZjjWKlvwmhZaNLkhDTwSG6PSo
xMfA+QUTTSwaUuxUop6mC1tjAnpBL7TCSoKhn5G06LngS+DMctpL5LFhvPWcEAcT
VbHBwk+Kuxm411TFtRs/BqHsjSrKqycqGcF7O0QZHQeetqMygdCkpV5+58Q6X0Em
H4oQmbaDC9OkTAaMcz5B24d7DySEf6m99G8MQwWgVGqFwm3tc1+clv5NYm5ZbwgJ
r7ibvxbu+hwtnTTNMbN3TJStpLhCqmJOepeieahctL4Pe7+50hVvQ0/EMhIfchCS
G5WSFR/JqgSdHCNoMOaZRzoh2kixMuhE6OsB+rzB8AF/1xC0PqrU6s7kQ29byFOD
avV1B2FCfrVUZttZ8byeETG3I13hq4YIXtjPhwhXsgB+4473baVWs01ltOUuuPpM
CpQw1d52MJInxCAl9zuDo+cDkCba75+qTzVnpA7BTwaPMxkEjBI5s8fbeLKubuJJ
eyEmYYreTRMxJf406JidS6+e+3GjhrF4Xfb0/+gY7FWuAGRX0nR1iDGxrwB23OBY
N4c7henrC/xwh0Auk0m4KbX8untN5EtkUZqsvcnqnnsyGcixNnrZaeV5+4upvozc
9pLeRbJAQg5uvbcdu5NWushoDAT9iv6FesZVmyWbwpISKn5gODZpVEzSlNqofAt7
XLbXl3Yyif3VWl12KziFLJw9E1UdlFmvl/jbuSXpfJOsPnomow5enbXT8K2F9a97
w4Tm6ORirsR6UErcB/HeR4g50YrOqIX+m0yGkUtTFGve3gn83IFrr2q2D1mN24ju
xXeKQ8IjLZfLAM+virWJuO66G2bV+Js0G7IorAZJh8RqCiEJsgtXlKKxYLx71314
Cq+StYjSfkAdTHVs+2SXI9+dve9ORTnA82ic1bImOFscs/FXu7htCnWS0jrXO+vG
GH6mSbMT3drLwdaIRf4WMW6d3Gpl+eN2Kq7bIhzbQFjtvBgGt/rswcLLo7wbG9VS
RfeRk9+n5RHelu7t2qHvwvcoyvXJ0zC1pP4UmYaEf3qMqDQQAVxhTQBjdaMsSGjn
KMYRHC0rYXws8ZY8+0NTJaIXE9XjyurRRJt2mhnFrCtqVUlN5L46l8RPTBbEJOl5
TuIlgbgfl7BrhDorigfWwiMZhL4o+erPgrYpkzZbFeyoroI+Zyj/CHIKPROcjiTG
YhkZ+0qIMkPvd/pmX21WlevxFZm5CYAMWmfUraz9HrXxrKS1uOs/cX1aR0jH0KyX
ofmMN22H1jH0cR6He/oYF8n2impS1zmsyl40RE6I2iTPAsPW8npyCd4IHArcrhjc
iVFPq5tPLVI2GLg60xJ/PEqBgTiD57xeNav0nPpxASHdZEiT/wWDnjCmTRz5YK2+
+PNKvel0BWax4xYisDNCbAdv7kKWcg/6LfbL2fUthmbErv8MDP7AXfGzmUvM2O9n
LpJfe9x45lSpTupvzABsaAcehX50BP/sP5d6moUTaLl063bUMBjFcaqoMsVs9Wls
iP7Ja4CkHC7aI0SOz63ZmG38o3bqB8dzywEfemzOnJPcKxHQ7VCUEeOL2S+Q22aa
8t6wQ6CvG2OVGU/XsWgFJI1Xt6bOn3s23J+lYF5I4Ulw/u6wPkEiyPQMyOXp2Obd
rvp4Tj0I8Ktqf98dqvcH35sm8F/dRUk1Euy3DCV19numPV9jbZg64ALZXCrsDFLm
kfMjJ6hjyN8S25lNPE7YxRiIab6vphbr4QLD1bRsTfRSvHd8UW/SGhML8rIA25qe
263N+8eAKZzIa/zySMR+rldL7xJ0smU/oLdiA7Jxp335tgW8TKY0e42S+tlNn1d3
wJn7aXmkLwNGvZ6S2ec+nH0FmP779gY6D2jm7PtVPnPm3U0SP176YfdBdLG5hT8T
t2FG5/NzuN8jjCRbNeJudjmBE3ynBGw5lL53ng9/EcwmACxYas9I96JZMJTlXfh2
waPQzeLij2dS009xCl6Eglru0s+XGmq7Geu84bYNzwjuB3+/N/y+0a7dUsR7a1ao
UeFc31wFPPp7sVo9m8zLb6U2Q1Mmd1r4yJ7ZOIWXoccNLFwGglRHbu1Pc1guiJ5M
PtW9Tz7wYe6DsMbwK0XSNH+GeW106bKhuOXgS9VffzcMDe1aHzORgO/+eytkrI4V
+c5UyY5dZJh3xcwm7AGDknC6ptLCfSnRC2dH3UZFEqYiUIo7DpIqDiwDQ4k+9jdG
aupO7d20O6zWniiSBfTCxB8XZhTA3fc26CpjrrPsmwGSyEE0Cug7Ckh3TQBYNMqh
Me9UVL7DvhRBruh/tN9uKMQqnmZcFUYmcYky1zv25VyuwzLBngdkqoh7dcqyI0yx
W3y16497pI6ETC65BDjc6RVHtb7j4g/uDQua2lDvRw2DGC9P4YT37S83qKa1RU1D
KtA1zoU/ZPQyn/5/Bu3oJoejL5SJo24xMzZJC/QzQ7JAmZDqwHvbaPaRHq1nUIuF
rsfwhD67tMrvrx3n91zFm6Z/cosmmW5iCZLMTnbCr+w/A+S0GcLFMWBdZiN5s9iO
7S/e+cMv7i0/0MEmwtS4lZvq9M+uaPZcWGHjIYJR3McvfCU+cNpaPMZCwH5yzFfJ
Z/9RuTaoyoJI6+SnLoB/b1I4JRmhBWGX/bzWylGzBz1WZGTOUgCivZjpzcc2st9Z
NGhj9nRSM5Qk8bNZEh7VG0bMzINnR6z0e3ODBmNHSRq85t+8HxZr6AAJQGBQJZ4F
h9NXG4Ds1A4xLNLquopLjb0MRsOP/agI5J9tu9NUXRGWnB1F8okzpElk+Mdqpgro
SJFp187oYy0TRL0yW4yLg7vt4PbHe3OCFAw3vtB0O8PmMRv4C4rj25HMzux5fxM2
XuOY/EUTJxHRqtLj83n8GDdxf9sF+060F5qLJ8ZG5Bb+A2BKusHP6+RDZXuIWE/f
E/5zIvcL46uoT6zh2+2dZSb9Ug/ip35P4IVUz/FRGZKxupl6sCsAfEv0oEJsDY1B
DGGbQc1mPY+Frl+hYxJSSE+pTT+Aw3pkdXiubmFSXPKEIx+BxPkkNw0b4bZFWIxd
pZ/wcJlQy6CG23gCSWc9jVvx3gOj1iIpHIhDlWEvPuIxCA5fOIwTh8+4/PKue98g
/A6uyTEtqhXdFBc6dJrhp/IILwC60NZIinPRW0d7zBDF/xJwrnlOHYRTSHjdnVjR
Bve577e/beUmwg63chKQzoNDoyw4Er49515VEOZwb+wC6lCgTQnsA2YENO81AVLw
DikKRpHqGOHPiCabKi4aH8uJ1lSPgGDd1AjPUDBYIPzrqfdNxCLpKTDNCrQ6dcfu
bKipnVBDRktO/iw8pJSeEqaIhukXvT6SKp36mk2HouGNma2mArHAAVBVAhodMyJd
VNNijiRybdwa+87LSrEiCdk3DNBIcVFnX7yOhXGQhwvvDpGDy/5bgRmo/mMDhDgo
0g3LfKzmOz8HbESONtJtj3N825c8Zb+ulm+bNgLBLXsGODU3yjP+I+b+zN4pXhg9
ROsoPj24olHlTlOK2ARSsaf2F1ETPiXBPD41wZUmlVBpxA0t+iLbe85BBPZTZtTe
CEjxcZVgKLDVryNA4AACZC36JnUjxoZFv39YNPXZNID/6+XeEpA6kfyu1MeDcNNV
mD4lqPYqlKaR8OtuDbw+kL/l6FbXyTWOI5MZ1UYr9vRu7cgJaH/aFpbRSosizEIP
+EUtOnV9RJPb4RLfadRkcNL8jAZg2mzWFRy3Gn11WxPr0gUQlYp1BIjHRZKDSrHc
b2rra2KEt4JpI2XAlgPqgglPSp8LjDI1pr72XUt0NYWfYK/iE5iqPU5xmvpnX1s2
1QGh0fNfFOWjPBrvKv7CXK2c16+6IQEIk9uRpkj27zU2OqqUzfubhk/wt+7cbD4a
WWlliHJ0p4gtRj1/z/VuedS40C59hCDr1BXBKONEreWHsllLUFa+cF7DKqAWyR9I
9ol3COEe3pq9AHusVn9qC4IHL5bxHwmKG8zFdfzXbxEJGmm94BSUPvrP0yisVqrf
iogKTLJ9zX2oU00LZyEE2lRc9TSGghcKX0KAHEgcsU+UjZD64zR9G/S8Vy68RJfL
eKedXyk7fJ+ppdaJ1A3OXRkFrwarP2yOSwcFpQ9WdSqu123ZIZj9FZGmzcTEZ9l1
b0vrMHE4J7npU+Rnq5fmW1ugtVLCVRyohpziEoyFCosfn7lrNXB+0ZhnHfIANWAT
QztQ+LEplpg9B6Snn0IQmCOxHwaAwNe6tGqCiGrqqq5DhtUlKFbtKoseoD+0kG1y
HX2u0to5LB+uX+SfpFXFqLK7Sjueht/RT3dTczaCupveCDFLaONFk4vceTKNsG0d
9XKyV0OOXvKQH5UhtDME1FtkDIEVVtoJ4OIysbRU54YCzwk244IGQf7vzQxISRYL
xeCmC9nx4PvW7/TN0TY7gfsm36HDmDXgtvBn3X4/HEdK2JDkx7WQW0EMMkmTZjfG
us42tAfhvpwCkGfGOpW6vA66KFeR6uBy88ZjnLZpUejh8czy3r8n3kTPz1rLkidS
Z5X6AVkRet1ORX+FZNgy7QVS9uQXth9BXGUhJ7YWQaCdDmqvrMwEl9XohNUz3cjo
9pdhhEh/ivfRn8wIQ9UMd1Ix0excPd8OfGWLMuiVN50a4yXX7UKcyFpJuts1rU6L
sltmloU1x7JNOvL5kw2mpZ+vt16fzsCvfBEMdqnI5z7hK33O9cErg0R9JfEN/b0I
Q+WLJLWdwc5VBjneSDmyYkqNMkCbiBdkU/PW8HsACsfrWkeJgpUzVICXGhZYB/Sr
jo4sTvGZGvi2aM6IO1FUfTCgMSebPyzDbs3JhzJ0IiNRiImS2kq9ASfxFymrr3d7
S6jrDB1vuQ41KvdpYhKz/fnaRPRNTksSF1e8+nTz96TazrcczhEosWdjp8b/n6k3
4gX8miZqyqaJOMbPVj1uWdDFKdjkR+DqsqIzCL+TQmTmv1Xn3OrL+P/lMtqj9ZGU
qJFYR7lUm8INvv9K3yCXGiTk1jjduwhf6iZFzZ6wHziZVLjY3EwlQf8Xd+ZqdQIt
2aiiq28m3fes3O79THqGAt3MkE5qLq+beZutpISwp6fKpETl1SPU6CC7raK+9nGj
XA4ZdWPl/hDc+TBiK9JN6p3xQvfG7C5bKIqFvowK8ougLSvWmACQRVhYkfWYXMdF
iYPPZKHR+OJy1u6Gz29UoSkTKWWeVJbxuLy1EBjARX7Ym/szCfTYU8RDiV7fzmry
a4+QcwmL6vTr+FGZ5i+XYo3R0tFMAzNPt7w4RfhruLaSk+FqXHZg9ZyfJJPvBcEI
fE8lZt79yYv3jc96x/6453m975PhMRYGXwGgFNYaE9w4s+bFGgXI9fJIGsNECoG+
YYSAQeQWyRWVpT8gpB795cniGImLClWuNGGk6cjshQRtwCpdvAQnS3ihFl7pBbxq
ZyveDa0wgI1Kir5IYH/TZCbxmfcO1a6x0ea7C/exDMzDkRVrwd7DDABH2VvRI3fO
8WjFDjFMjB4N+pcRVww8jTj6nEy0g2+VeDqjH5vR5RfXqyIPZqc0T2h4VsH/h1Ie
uj3hSE/A1XtIK9MaRIqHr4A937PsG2WNXJ20wlcqw05N9ILTOOmx7B1F/gG53KpN
gsWib8k+cNRjiu+dWzCqOEU71GJUzkVw6ow118Y7Z5pF2mcR/OcVoNzSBhjxaBqB
Co6lEh/abWS6KwebHWZaJEKqeYecrcvp8lV7Mc4bhxXvGEf4361tI67l00iI9+Lo
ikyNPW7YttR2/n2YPmJcIp6DLkwsFazQi4AUSm8lH9f/3h/tqZoduCQbnBNTfKjG
zMoLKER3iKK3BY06NgqLyMpASYqWi3h+uedRAmispadWbuxnc89MoqvDb5L8G9yP
m2R2LfVA5KvSnM9eyale0tAi0JtR7HrOwx1QcDJ9isl1we4dB2IKqI7fqTKURPaG
PNgunoZ2IGtSUeMZaz91io/iFmmWfTLEsux8cks/fj4fg0FzHQFPItZ/POJTh6FP
uQJBaHZ2MtP6rIGG5A3exB12jbDN2T1jOkArC7oggQcGu8KK/dO6w9bULrsFEgmm
`protect END_PROTECTED
