`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpDiClFItjQTKNx2af+7q9LfERQ8/1yhysnRtQdj1CqrK4Dop8Vga8BeD2jC9LFo
qOez47kxde+oYvKYH7nmFo2lYtpgyKb4akhpWJ9vvEZFQdelkBXzcBZ2njC5BQJF
I5PC2ZW5OxlJYGV3ZHdYAS8NXhVB3PdU5kbma4QyP3VeCAiyDF0wZucMEv1UspYX
uxqvdQx4CFXxt4RIFpDOLyLJQoGnkAb+a6CPo8w842WMGeSjIduyU3lh8Cp1gkVa
5ctt0FdVAdNn8l369AKzrSTQlXhAswTwOMCjMZuPjFXCl/SqzfUkN8kWXMb4cGwG
a/ZKqsW5cLKXyVzBKtTt4hcL5Wl23lAHWwv34Q9jh4dlt0yS2LO42+nvnHYOvNl2
NkN4ySU1F6K6GsVJgYtbw2w2U8felIHhrcZK+PhPkjFUbwfT/pWwOfcTzXYoNE4m
0cLggfS1VDq4x64JOSEu+J0Tup5U1RA/7U7Xupw1/Xl7hxg9zFswvN4Ruqbxi7G4
YzKvOqUSd1QroxAD1TY2jkHqA+moEZY3KCUe/jJfhnNnM0TFYl+ZbihyPiiuybXt
sSOlf2zmVoprmjS1/D4g2bOlchWvZ7pV6NHJQP+Czy412WBypCcfP7cXsC2shIj9
1Ta+ST22I8lQk15AQ2o3BjfYaAKKN9MnEOkkEX9cXxz73+8i+AWgwkycVxwOenW2
yEpdWDE24GNTycogBd03En+pOWPvovWdA/ewrTqOyDMEn4j/VcWKufc1NVY2xcEw
gzukgk2xIGwVSWTTZD6alLY46Rvtie6vdeX4H3B86Wu0vinfozT18PvgTcnpUw2V
JiougMN6MUAylyV5hXlyBc+Ee7Qt8YZiEOA5Rsv/bJM33Cy5YCgX6sLsF6vm9lvu
C/IFLqVAefyMfpXq3v+MC6Ynk8qz/PJoZY4QO1xQWpvZ/Hvf74ZEDLYp6ySw16JF
fGt4OIOvh0RQuLD71EGUittiu9w/xuBztKljGGdbxm26gFQVjCxDYLFwf7843q8h
dNb+9pVnJ2cg/RbxyQ8H/MtwVlejuw1F/dY3Iy2C65vM7uigzk6C+uWTXFtFWOg6
DL2nvKZBzQyCqaXztrY1XdNwr5aw2jdYTwSVdH0aMclFcBmgqYTnU8UZfuwYpDEw
bXsZr/8Ye5T1YFPtGBvHQ6kP5K7/5bdv+h21O6P14XyzjOpWlSYQtb2tgSBwEq+/
cgMc2uzJv8DMQz7pvqm3hXvIlD13DG+e8KgDcmh5mtilWyGvQN84P0s+Oq/P0IhY
NOw+u1NvmXeYj84g+XPKUWIAj0+R6z3gz0wknSYGdaIFxz6Go7Akj7TF7mSaJJay
XYRS6bZrz5jGilnX3dPbTGcHNziTjmXdiAHLLSjPC6U=
`protect END_PROTECTED
