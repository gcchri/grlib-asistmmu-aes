`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4MoWNDBZcHD1QGsQsQ/rdPIsYO59KSUo4c8sznDg/xodkNm7LeH+gJZ98qLWmpjU
49y6wthJtI1v6IeV+++A98BTGjKdzPvsG5drh3NF4UdPRg9kn5ou+YH8MgMYH6Jj
jLoXkCxdGB/brFwfU2e4x4dCAdZhTgFULDIUIFSy+7eQYK/6zoBrLsD9SyjVy/7W
xW67UcnSWNuiiJ5IVm8sUyLJvwXgUk5csUrs/+imZyJkRIgpmxsYIwh7t7BqNVFq
p9nuLpyGmJRUuVTmkWgKE8HMO+vtVMAjWObN6chCbNpZyCmOdvhKDhhIQND26PyD
RolXdyX2TMdaq0i1ymfq7LgQT9PztCBAZEl2SMFRl0fTN0zA8nFJJoM6bZyoe4cr
KXMQLeZg4jUC4BZfEA8rug==
`protect END_PROTECTED
