`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T883hIFd9Qr/UHFAAZ4QxD8RnSZHsr7iDFy7Yxd+LlL2D3ASelmWpnkKmveMrj4c
xcXUpMmuRGq6jaBS5fcXqxOy+HG6POe2awQ6RkxPsH2qCi316ExKPQhgotgr1ul2
adr3GAdK8y3pbbVUaZs7BhwcG4TQBbpxZyERsMZY/pJiR0dO3jhMKD+4Eokf6NAf
SZwXJfuKk78KX3MUWkbMlhu1S8rEiZWhzOXeb0yTrpIgmE4NsvNlOSsorHHkQowP
dEBZA7zpu/X888zmEzJhrR+zWhpvNANGSFkPWN28RQDigVHHArXMhmmmnScEUKwi
zBB0MXVGiuKEMKEGGo+QNB2l+9xw4iAHXYcEzqn4ikwCGcOxYS6sUYOu8/TZFI9b
lfNL3QN8pD04uekN8scO0WeJXPhT1AfWdTzfXjOOduVGN+Q6dYXkmwZsRttpM+ZK
3Lx5L31h5FEZD5Vz4xHON2kSrWO5hQ7rkkGgxXwEpq+iTKI3O0OdD0sDsq0ZnyV3
RddPI4RYPuAFr+EsgvjTuzxDOrgN8Ltf7EFwleGS1G8=
`protect END_PROTECTED
