`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y5zGxm9CoCgzmyuKc0+Ls2/PRRx+i3aXyrail7s2O+ZmsmJLbgRnjQBHbkYrQ6SI
3bbTR+rZ7gyacKweXJmZHr1N7jo65DRVwOwhONw2Kl4kJ9IQ9Radeu3YsneoA7V9
cRcDvLE86pPfXEGkdNow9qSvme24QcInf/0SlSJCiH0DMPygauKi/hNZsL9mtJmi
HYWtoDfrfXmC9ICA1HptQPi6CJ7uJt/2VAbbAy2XjUuvWrP1UlwOP1mcWW2jcOf3
KVTCZrUvuWAzyZWmZs2Kvf1RbZkTppHqRox+C37/Kz+tJedPEtEl5DYUbn6ggkfr
QkkWdEMDC7QsfiUc1LWTK2Y90mrYxbCQV8ZWYExwtyty8c3F2SYeT7woq066TUna
aBJaiSmKCU5pbWVUIasV6+y8qYJI/WBPuEQmiORywawtsRpZnvoygs1/JwQKqaAW
mN0k0ffBtb/3TUAC2QXabLdH3GlcuIiLKvUChKgO5YQvtTOsmb7zymgUFA34Cz3N
FRokqCDcombnBbR1O2D9aUmQm7h5QI6eUwLBb6HSmJk5ZjCIchq4Z/g/SDEyrbE1
4UAuqgPEYFjoSkj3isEU5ojjx8qC1Tv2wXKH3hEG/giiWxn4Can2RmDARERAGD6u
wi6N7d4Ukmi8rtIKUUwYdbkuYPxtYkKNFFr5NYxl7WTWfmm/C4Fz5uWTdAVCenvn
p3PkCp72ZqQem15vtu9pQD0L2Gk1yOMQuJZknpBnMoV9lJhIMtEDnc9HFM/JXa6e
Tn0WHjbswxgORGNfcCdUGNblVdMqrLpd1m3teKKOnAF6uJSmU1adCnYrPJ3k3E7m
y4ch77SzMSATI77Xu1oDfeabrStS3eZD3k+1Ba6Brhkk5b8A/aSBReQprxJPkmTH
xqTMstJ01RCzbuYiyUqUSoQNlcVrqc4VKT8G86y2/qtrSFGEWAMniduNq4kwXUlW
WwHIJxT2IErxC9l3+GCuFBy3JDntY0qdLO7oBmmXpOHFIJqMooBdweMJqZZlL0Si
cmslH1vUHbeHUIYk7W8Xgl05y545YKWYcLDQkRly68PFMHa/y01y/Ad7gWLa/RBa
TM3Hz6CRXH6x89GQdUz1l5Bo85F9i7AKV3AIzGkoieqDeEeQnuBiukP2Uz4aLOlG
fce9dGkApxicN2HHSQ2YXmH+uHt0WmtpLd/a3/fmMsTT0hMLtqQSuKQbZWtyOL+g
EI8i5cCBUrR2hAl1OZHukHRCNvTJBl5CqSfuyGtph+JcxXeLa1STNcaic/XL5Jl7
V5SSN2MnSa+WZpQ07inDh+CuOp1LOgDswHdjmKo5gUKvJsHaCss32AIEeaq/xyGt
PrJfdqnuv27HN6ZANp1jLg/OmTgZzKAeL4Yu7sP/8aPkvcEppLSIK2U3KKnNxuP8
Btnp6x7FITMV+ThhejbvOhT5Wb5UJi9UIk3EKNC/4WTAAxH8I6hqTLSH9Q/IbQqW
DmjgkVJfRTwLr9AjmYxM04WwfQV8s23g5lnrAzz6YqbGfFF+n1W+X8VWaEQpP9bP
xfT0FzAPZFYRY6JzBeWoNIBZV9VcsXX5tY+a8+G1WgOsJuT5spwnwVHNtkbeuG9v
3X2et21jgbK70M5eSs0nEr3oFNE8Ecq8kepwr/myZkkngera35Qsct9IpdAztvqq
sP3CydADHKYgLZ9WwSzVgKngj/S8ZvQM9T/1OMib+RF3y8k1JZRk5f6PNyC9evvu
Yz7cc/VFKDwvbscb3s9C99nBCOYcF2uhaWApo5XHxo8OAr1Ypg2IWNj51aND9XD2
DTWTmKqqUbXbqfJTFQiVT5yevQOt7DkzumN81rJr5YQuSrxN69/CTkU3TThme05E
DQtrjPvAK9zjgG5+gFPod3Ndl3mIusgrIqw4nq+0516VkoOro4KY2rTQTfWiZ+C0
vXG2ejpEVC5g2rFOeBMe/+LaYluftF00HRMKPyvx5CB60gbkd8UKuLxPT4OppI6x
HuLkR//8mWO8UjsfOb9mlezIHSPhudKprpBPW4IMPveVyZZ/hh0yD9qsnZxtsEUc
+JjgpgR+G13MdI7lB2HjHnmNH0pB4n9hlnR0k6ZtQUAYecbE/3/c0683nru4k2L9
oXEg+ZIZgCXhbYlL83ARygrsFHM6sBshDeDliEYYyZOg0QUDTWFqKei1jzohRom9
sD39Mmt4WN6fSZbtd/oi1ifXj7V4jzeX/mmr7Usx07gAYLYs80OEaPWBhzMRuxZJ
F/3h96AfoRQXwSrnqbH9sRdzeGLSJ+QAOuS331Fsm4cGBPY67AbxsHeLXNFwY8pw
VrH0KL+Cmq6MXq5/Sy7m+DTyyAey6Q8pbN9uSArJ+pOv4YSct0B31N14ECAWgRZi
M6qBlhGQL3Bu610w/NqaO3gSw3lolYc+oFdvIAMNBn9LJqIexVgvokwlaVp+8aTh
AzO/lemg8CHekQrdfTmGu3Dm99XQKuklNk45SMuH58xAfLmDLSXOQB8vr4gFekAy
se6tqNkocVwg/UP+nWAcfyW1LX6zV1dRHZ9eo5Wnxi2mHjTM3JrddNZImXgXiOdC
Q8sbyDxRqfrWLWmHsnp0MV0p4npGNIjDiT/QlF9Z9dFXVqvm8sNQMAEhYA1zOmQJ
eA76m61VvybSJu/4SzIcnQ==
`protect END_PROTECTED
