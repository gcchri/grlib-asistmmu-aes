`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iM8f3yguLxe7t3fmNy1Nvxvw6SyiqOYIPRrlNO7pZEgqV17JvupN80gLmHgwDf60
TW2BDQJzZDLYRM82dMP0uk2/ULIEXqR/ppMXtBf5yl4QS+cIdG9++H0rsfX8RsN9
0qv4Yu0IMZ3tuAF+3gLPls63nUvYqd6ka8XFEbp0Y3gEHC1rTpu6212WkHebpidN
H4HYAqooysAJLZQxk5BxEi+0jANEjf5eoDk4ZWeZEyRo5Oe2xMxYycBNb63rCBjK
nScpm0wbG19ZaQ917vID4Yf0eGDVGKfVbAs17SFLwnNIGSE+AivIQEgLCQ6QfOwn
K0SoI2FF3kqSeav4mBXUUMoD4lFl7jBpsU+KwSUGNqLdyjU6V9ltLSF7is4pAoQ1
gBj1plrZW9VSwCI3LZUWWrnL3YBAy2y1drZohRXpQSQ=
`protect END_PROTECTED
