`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
azugFOmsfKbs8hzzMs4ARt4jouJFprdv50YTH/HHDF4uj7nOTnFs/JSKn5fM3qY6
WB09qA/N0FsuHHCRsfprU26i4KlO/HjMPFsb5reBGwGIyE3MtGol1aJMeP2F8I0w
cpx2khUM48ZcpdP/x7w+jQgcae/ggSwqnSVKK0kNOTZwo9lBxMVG8SXVejaSKKF1
KckZ0dKOO6kdFgtL8m5gooktCqwUDMfkecJlsuhx8PIvwcaeDxClOYKjAxBvBjFC
SzxHaT57Ye01GFCAmTiCpyA5RvwVNQ0/iSH+v0bmGtc=
`protect END_PROTECTED
