`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SDdrokWZD8q54d6D9oBWeYUUTVIC7W2ARMTWKWgi/k7nHnY4ePdSMRGiLdIINXzc
H/meob7yn22TYDC58Max4KX37ENeRkXwLeSQI0otEhVASBoCx8ntPRasC20DG9Nq
xBlTFKvZkl50Xvq+4v2tJ2Xhj+GiWhwNNWWA86/0AidO5m5F6dWbMR+So2vmusR3
FTdcTV+quchX9fuDw8OZDfRQ0HoZN+p7QLpyS0yupy3O9RXSUx0rTNk1eJfeGAeR
JyoKfzdoG+Pv8Rlz9Nv2VY32de7GnsnGIzQLjb34mXZ4LIPFaq+osfqZ7lXo/txV
ICiIeXQyflm6ytoqCyyCP0CwFrn/1BOso4u5LmPW+xJL490ZLNd+U3FkUoumJzHX
T0Rtkc8Zw9aKgVProbIU3g5VscN97ct+GEKBFbz6ShFmFm4VRT/iSM9H4e1BGCpH
`protect END_PROTECTED
