`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sTavMy0TgX6hdvvA/uN0ZHyZMcQ2C7+6Ak0IGQpFFiejeqKmOFx1K7SSpRD1VJ0
OK3xRLJux818k9mcvnyX5WAKOw+wTKSS452KwNc1E/Dl7rI77+sVcc+abYTTlqI1
Qr7SkvtgU2XO+sumo6pYvf+U0+esdZutKslwjWooPac+pvayJU7Z9huHvlgIPvCh
0MaYVZsL3c2x5BirlS585TQ9lvEJ9Ocskgq4+gq03bSRJZdLfW/4VKEVt7quIsA7
4ehhcw7Wtltdm2vrSRdKE4tce476enB7bj3YDDyXTkS2/3ZYJmj9rTcSlG4/uYSZ
ovMbV6J1sWeDUsf3AtzZ9z4ZX1j0E7PKAHhGxSjX0Yauu9Jf/kb+PJciLv6yDR8z
CEC0vVfVOkmlxZqQd2dN7C73TQ1GE8jRBtKNdWZsqOlMEvTfBkriGFDtqVaCtg/C
E9KXP38XCc4Ne2ibBQ+296tl7nzxsOfWp/2WFqCwfOWpi4dp32OxT6FmmZdfrugv
`protect END_PROTECTED
