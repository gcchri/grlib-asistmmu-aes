`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LYcYgRk0WlNyIM3SK3TX/Pa4tJRch95uLoKJj19mHK68gBMOqCw6u3IMWkYzQZVi
LCXpJyuljm9r4n4eHSBALcshJf9VfyljUY4H7ltvY0gdq+trcqGoGwD/ikWMBO5W
uk5NRTFKyShHOq8EbW2adlccCqW8ihs0bBrOWN6iLbgd1Ubm6uAmctMyRru7e1ci
q/LM19Zu9dDeDCaqL2U1v82adEkjkke1+2b6DfXJDdLtzYXrQ7/OMxMDWRiOdG7O
`protect END_PROTECTED
