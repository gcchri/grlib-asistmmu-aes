`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ukr7sim6jpA0g2U/SLV3eSD15JbuXPn+vcXQWmK+BB5/p53VQ/Dic5IpIikZmLxf
jLXRfh4MrVV6YKyYtehqTHLKpykVZbop7YQe0qnJMzCQB1itojp0GwI/YL5uiNW0
HpvMMd+yQuiOKM8px4YENE4XGyJVVCE/xn2ffa1dvLvYrmAm/lWRM0IQbsJnhKk5
UVJpeq4B2Y1AdtTWQvfGk/QPYYpeKGdmgXw+Eo8mw+xz5Td8UVX4mkhwbT36VJ9S
31vvHOZoePufnMCzAz5e+eQRsjC5Cc/fjArLxFikiv2XeDjQPP3JME/h7CUB65w0
bHxKgyHQL+A8vrfTubAo6hOKv1iyPoFaKZcAn1VFE3H6CtJySHbJ7irZnNVyTEQx
`protect END_PROTECTED
