`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zK26+oYxuiDkpEgD9xCFFTjkMjEOiKQemdsRYoQroBNdbmRZTlyhHIRglIXL4aOb
ke6WPzrwWiKikMh7vcsiH4jwh/Z7dO8sAPAvUxKVHp7fJ+5umQbWXtZ0ZIP7yAJM
0PwcmZtKk2092JgzLw9RhCMJAdMNrULEHi3GXoj6Jf+rJgAsKHlrBettHDN8tmiw
DwPqU6f1CER+zjWcKeOnSpfNZpp8kuUd3NDb7OGByQCaNQ6NnlDNyZxp2XViLD4l
VMUzOaghVLGVfJ1akZZQGRvCUXInJCirPFh3XccI/rd/+6DtvssqqmTfTT/MEzNP
cUu3wIuQ19sDmeC8N+hXQNmVRoYAZkFkNgZvG0ujN6FPLQKaAWYaGal8cHq/uqL8
Y+MyK58rceLr2q2Sj+UohsdrauNXTNzsR+/WegeWagBHz7lAnSz7sUjiehav6qbK
KjsBfIGZb1p5Y2Ow8Ofg58DJTsc5ghjotfbzSOo0Pjg=
`protect END_PROTECTED
