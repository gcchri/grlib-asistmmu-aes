`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j5nj3lnlhRb6LShbv4Mzf6OeXqEDCbeKwmbIT61lCrstln2eD63l9gFHr8bSSetA
L8JWT/4P+19QVQFhcpe9U4+5l7gaWCk3S0+zz4QUG2kdNuoF2W2DI7qjtR3mC0VS
pT4GG5yTKvou50/c7VHWhqdEyIzK2D7IGwNreIG2GhNN8y/GIOvdxDVYc6OZdMmL
Gty58SkWnaAc1lPlj4zqCKVy24JNs6OuGoJkMYI9aZsS1t5Cgu+MOvs5xn5SFd4L
qz9Z3+M7FJLz6kNgKaZ72zLxOGArfN2UNr2qYivmNTFNkJIOGqij8AlWq0evi5op
6jQVKE/dIzVSAfwZZ/0K7aXmAnhlnvcCFle3kDEcX7Ci5SnnC7TcSdtOiGnQ5vkr
78QABvPi6bOHovReW75B13ZU/2yqO6sKlLPXr4+iqy0mELuBoR52mT+2IIfr7/ye
k7kUmtyIWTDEXRlY5mckRiN25jXo0S/IqqS6BXTrpeingGnL9qjmvSFPG/DfWwAP
+M5QPJ5vo5eqbpl/r/+oPl/pyhvJVFi0RLm5e1Yq0A9oOMnq4a2fZ3ZJS6l7xZkA
dK3643OCb/0NY8MyBdDH931Gq8q52PFxpZ+hYAIDIKkzs3ObWMQGK5WH2ONjc/e8
OyBDVfrbd+S8534Ie6jrgwM9ZyqomqWAePzRROzsk3hKAb3yyVBoJ6ztqWKW8k/S
YaFw6H/B+qVAa/g/UV+2+8Xde7zvduKnx8r+AhqsjUDV14+h7ykGLScCBLY9JR4w
1+kvybC3xJvZzhX9EF0Y3NvVA/6+sIX+qXr3WlOPikH4XnsYXQ8Fx+nb8+4R6WM5
hDoixCGiQ6NJJSF9/uQJnYYPJc4id5yXFd+ffr+rqgCPTmbeTXOBGE/IgkYIq8NK
KqJSCYPhLVmPpU4Ghm3nkR8ur4vAFC7ZKv3lXdJNL09CrlwWZS3EiMUyldJbWR5y
pQnMCl5g+I1BhvIPv6n98cSSGBKLWBI/XFWO8NG76zrkzN3sR6Dw60FwkPcnSEzX
TqwW57vs6dpv0a3BsnCybKvpRICqFsXpHgaI4lTgiDdvgLDjQbyUzZ8L80oYYlJM
xBsnSO3yQG0NeVSpU9ZoK47y/sAsoYbLN7hy//Mq4QrZzU+8c9Tc+AZyxztPPezH
NJKo5I5YF/OqbBZ/3AlPKA==
`protect END_PROTECTED
