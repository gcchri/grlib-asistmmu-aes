`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z28STo+1y9Y5nudDLKZYE2iwCSFI1kd7fohP2GtHhT3eYokRLbLivPQ7hy1A5Y1L
s9y5rMBkRGVdLzp6zPfFi1lKaVQrsdDfEnDDg2Rsn/m4hEPKFW5R9I41Vn6gP5Wm
tpwnqZ+OxwdNHzfPm7vFTy6xXirhCUnDT/8NPeTzplTi03xk/DlIKfxVeAaDZSUS
1KS2loDZl/837WL2wn8Mm7aikqNaEpXfKUXrrDycC4sU98tiT4Svox36akMAffXo
WPkoVpNpCD57OKtwy4Sj1HVn5A6l3ZCFCCHyJhJjIMl/mbDiSKL03KzUFO96pHGi
cbqREWHzdth/1APNN7u1O3EXaTd783dCsiN+vLp6iANiu0iaer51KNteoYI6c0Qv
UXUscpzm69O2ZOu7xYKP7dgyz5AAqirLnuJ9bdhQNvhvXeDHCrNtGOfeEMrNx0Ug
R3QsH1cthFXVM82NZ4QvNYDKgyvmljP86exccaQK5RBQLj8RNDrSLJ5Bsr/gMNr4
AUsy2cvz10G9r2ZoSD/p2N0+B05TD8aklFFDfbx2eoz/VW41YSMBLjdYcfEw6Bfp
EPvrvecNKqnhg32OaVRZRAGXpd3aHmdH/VZKqvcvY/EsxiTvnSZ6CGNHnVRlRrGW
St0o0Pp2NwA8w19zV9pxVzVTedgcS6GjHrkvQLQLXjHHQ4cPEEIKkbfGkhWSBkmI
`protect END_PROTECTED
