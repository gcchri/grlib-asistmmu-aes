`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/8dptVq/8a8bXDwL46qGpq415bfR3Nu7WeRYZl7c6jY6jksNMkvfP1WGJQkoib0
ynLhSKcgSniEFDK2BhjbV0wWg1WOW+92z6Vs90gnWOA5BjC90yvwOKsdgdxtAcF6
WHyZigvpzXk39cN0mqcUPdFvotsF3vPKrnWG1+rdbBAAuSwSmB5zdLbRZFuAz2Am
YPzFQt1xr0GdkADcJALUOSAWHHC0k5l7g57go3KaGcyiUAPWTA4P2W8yZpTSNVml
v5J6eJnsfkIdKQc9c1Xa1SG1yKyZhu1aPh/dcJe+5dud7swt/fM1g1BisAnBStlo
w2LgZE/jm8eitsrGimFeqOAJLr2EsDFQk7oZUC1owuUoHTTK4L0aDCIM4xZQDvn7
1GHJx43eJczgES2p7KYpD/SDr/yeFndkNtTioe99scAJY5gn6yxTCzLYbNFokLLy
CLs9Z8Bs1qL+1yqARpnmoBeXwVUkQzeK+9Ys8PYyKHQkCHxmjrNSF3xMBaYGVfU4
l+gRr0vr/TrYcyOcXZ4Up8aV6myldZoS/4hRBO+x3VdUfU9xDo/xEiFIHmdVl243
AbkibLc3riHa8SF5TZcS1h75H6z5no+/1wCbmt8dvbx+PVU5K1o8jJSUYJ0Sz06c
UDqHlrGpt5Jvjkdi75WF4M8bf8OklvO8VZ56BApGNuk=
`protect END_PROTECTED
