`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EiakeZw5swnz8kf1iDHLHZjsxSK/F3une3Cj2zZ4vSne0Ov+iLsnMVctHnSdFmWc
25ARqn08BlsRG1LKidyzJDYH/R0o91+lsTK+4hqc7f3AbI2eoJdyAsIrkQU4rGnq
ZVt0Y3dJUXmVhCUIJ6nlR6lGpZVotJLXBqbwk3ebEOLNJqfhtNfEsiGTOyZs25Es
gm8ekfWvJ+bQJwcZt/bgTDt/ujCN2v3nruxgQpMsBnbs49sHEmy45Wa4SjdU2D8o
ELSjfwtcAkE6b8ndMBCrgA8/R8bwCWJZqqhyJj0Fm2ErYkbZHHJ2eGb4lZBm9jev
3/ymBVLpQ3qEW1k88imGBGNJhGHIu8/Q0CCigdzpV4qlbENrbCwUnRzY3DXlzaO6
0xlNJBc/E/DFvKVs+iX/X1YsqQObZ33yPqPh5f/s3FbqAW9xdA9/Jtbtq7Q9dxic
RUbM1+H/SFTsHZfdU53VqlJ24NI5oqPah4BWPeuyT9ShiuQuYEuoAhbBbIqQI4DQ
ktRk/SZnexmtBha2vGHxhukssEMUb7F6IuZ7F9aTpWEwZvwOcDxNa3cIxkimCWg1
9PLgDqITBjq1XmIq/yb3rnBN0aolftH0LtzzEkOCayK3EQnFhkIjEE1EtL22SwZt
EtTXMgrpqOMEWbnLreb0Tnrgs3klG0/H9nz8+S0ZAwm8EwSLv3zVgWQP2aJHc8RJ
De7ADFtBlD0BZmkKbTOT8FNul0kvDOZzDNJOTkKEWHxBkfCgR8NjNQkohNmwZi9p
tKsVT6LXpkyqzFLenQBqHYwwP6UNHHTEXBI5DUHW4mBfLoOXPEQMzkziLzuqx+r5
z099fOZX/1nmVBPEYXc7j/eeGuyenfbgV228ZgFDWiafwa2DinP1Kz1BwmmtBLnx
M0jaPsCIccpnljKnEK17dw==
`protect END_PROTECTED
