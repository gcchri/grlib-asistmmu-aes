`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hzugOU/C+vlhKjozJd/ll9ZA5qpt3vIcMXcKwctgwGPP3y06to7fScwBoxm9woUF
n5ydBFowjfJmeMr1DTyoPRNobxexhIH6H4zvRJ7Kv2GP5He0hZEsIri+jff8+zCQ
1pnGCWsTpl4rfvK6WGzjo+kOfmXyHLDVBx1dFl8TV2PZ3hh0RkFR92bnUG8d/osl
eMx4X2thz25/t7wfU5NxH5qnAeD7pxwAjLnqSb/l5JyVlAbm+/AfCgLlaKUwswFI
kO9BOWzdBnaoP1xZ3x66/GU2M9pwrOofe1DvgDYAzsUfMdWsrBFAFaxhqtrIClN/
w4Lhx85XcPBwCMcwjC16RE7FerHaWkb6GZsx6vIptDtcxpOJo61sJM7mJoKRcInh
aOQ/PtPXAzFsG8u4ijKWpIVLi70IVRTCUMhmKql4JZN6AnFU20cnco6h9Noa1Nvg
XJBn2we3muKAewlCd0SVI7tlTfZBl9DmvKb2Ge8WHvI=
`protect END_PROTECTED
