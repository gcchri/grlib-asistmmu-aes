`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/x0rKfhauzHblYkGd/p1KLwvrW1CkJje0iBrVshOTV0Zj9uNAgy1apbgOEoEus5
h3cvSvkC3mksTrM6lNHP/pjVjv9UzYBWh8c6POe8UTHmyhLk2sVgEa1G19ZkHFrJ
vwylijF7YYLDRyUUCylYW7LULTnIPUadoRiaIaXBAEIcjeNLEbVx0NUnX5uqRMF9
ehBfdYAjI1QjOFv8ICMIhdJgD6f6p1pgHYcPWT9sAirV7bUTPpMI9dQBcXM7yVei
LOZpV3hzR342BWWay/Hp83QLPDRbF60s8KG53llHVKioUcmcpK/a7Th5JBjrXt7h
BV6ercZ9GwG8qKIrttplCyAK1+ZYUAefplLTZh9Uy1A=
`protect END_PROTECTED
