`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWPFHLcxOQaW88HKDWucaTOkRMWK+/APIO3xkKz4pSq4jCcy30wAlKZMCvUcyV06
TF1QkNxAisrargAkE1XFzz6MLaWVTLGJceoPXGDwKkOaySxgoMRkrw5YUsj/ueSZ
a5cbO3X6ZAbllozXRExG3X1PchN50NDkikeYQtZQpwV+hGDS3Da7qEBr0B0kE6uE
2Pg7KNZI6AkCCxe5Rqa6QTdl1Za7qmdzpFVWa51YmyWA8EqyGFOxPnQbKXNjTCti
e48kC9kcqX2Gw8CjePr9qTxq0IRrUSS2xSy8PaIq/+8sL+VzVodUtt4RLb9qBUBC
`protect END_PROTECTED
