`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jTIZb7+ln4oWzeDBH5+esu93qmenPueS1K1ptatOCsMBSpvZYWACKV3dSf+0V9K5
zJB11UuRPdKRyQHLgVsO9eOmS6r1L67X88lcshXRpc+uKeBjNGlGCJ6V8HrtMFEX
EbMBg8T1X+s1MseMnvHm0yRfvVeEOtYN6npO4P6v/UKbw+i5mzhmSCZT9MD0gu7C
Sq+zi2EV8Ghq9q/ljBI2PARzdrDtCRwruUheKMMDzYtaOSplWgUQW8x2HAyy6sY7
5lE8i289Vf5lqxCSo8f1KOlKjc+LTQmmp1C8VccIlzDfHq9HZJQPkYjBUYEf0p9D
mZWMthOWVkmH5S07RvCp4KdXeSGI4Gin7N4JjhMgLwWETIRtPo9YFPdK24h+DaBa
n4HxOtooJYut785sQlMZR8NdUKbMGOVB3wuPlxYQV9gr6Q8Qng1e5Xy1t1RlPLo8
5gRg/bZVG3vKoGqJNCK0hMMvdVqgDGKp0Wof377Oxg52XEclPW0xUniFSftbOPl8
D9K6BAXfZ5CrtyFYaVLEFw==
`protect END_PROTECTED
