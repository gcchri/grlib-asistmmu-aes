`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b24/IogNK4bk2V25Oiz+8cYpq/+TOwn1yVvLcU7dW8bqT1CA0JeHLAqvWPVrJMPm
khyVGcXNClv3d4XAgu2Dqf9VXnABVrTZ6ZzFYbWQwyrdZXRepIq0CyAa7XyQ2qhB
PpcPgRXV8SXNl2zOA7ipIJKrp8hZs7sqoUAlwCnXaCXagNKwR1pY979iGGd+CzF9
oLituyUZbVp6Uvg2t5vxUUKktun1mm4RgiFOCwhcH11lB5YnxYAku2dfFHkmKvvs
/2TGi2Y1vN4fD2Gysjve+bjL4YihPaFLfoDzqusgnFgkHtvTnsT1cRkKHnvgLiSd
cQarvYgEM4VF5H78boE78g==
`protect END_PROTECTED
