`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5lTpFqcHuzMGDau/T+daKqhcT3xgfqKDxgYo5vMAhA62Mz25xcHuHwZsJ7c9UfDN
Uam+OO7jguRLjmIqjBtiflgoNlpDEgaMAHhc4ZSu2cHRfQl7rWd3BcmjiyW8khgB
3s19+IRXeIWhxIZCQ49894AXSUe5dm9dAoczA3zRQ27px7jq3Eh11RESUVQGF1Sl
jmrumHSutnOCZYKMzQeFddKJ57CjBNwENgcxnrhTiOmWWjzbfADgXCR/9MGYfeqz
LFizmBR9Tfmj+o1M1315kruqVLP4mu0dWCR8qqvdKfHM5khi7JsHezTBUx6+DbJf
kZ5KYKMSvN+AdGdNoRymLPBwJCx+uLTwDe1R7u4osu8cLitQNZT8Zpg3eq8HI0ON
P4xXM6aEO3k+QD1DKr0pJ7r7fCxDi4PCxvqKT6TTQeioOxxnjzHO+OpOKKyeavtT
DoMhhyrFclQo8F7YGkgMlUX2VscE7ntoBsKDhuO8fUJn7URhxJYJIqo2BDGeoCSe
4LWL+zTNVO0CYU0D11BSud1SrWZRcKuwaUKoIjOS/W6G7+R0ZE/QEnPlp68dfCgR
mmy+d5GkMQ/8xAYT0VVLvMyh/QuYiOtKuDb1tBxV+ZUo7r+pHVAhrwQhITj7yH7z
I3F40EKqjOLkXUvdzZEzww+NSOanUFHt4OCBzLF/Ti+Y42QoWHmNs2ihF2KhJ5/a
WEZL+RvNx8aQ0P2QgrNOCas/nZ2RC5uEfx34fk6/RYyt9L6dlXALXZVDmaFt+fTf
jpEfj91dFAfVKMLGx6iqJIHmitawwQUloMn1B8IyKWlN7TapY/eqZrzaOTEV7bcM
INDw54tBUfB+zCv89jfFjR3l2+0XuxaRbCtCLldK3V2xrrCrygTG/w1XC6ztxHyM
BeIchx3uJiC9/xWtswkSdqm+b4XU7RQO6g41Slvfmvfg8PRGNZKeoGTjXWjiUyGM
NlBTPmgnZzjhlvfKfPGvglfZfdSILmU6R7cy+fEPXHkqe70rzZQdN4PNljckYuyL
60xAWjySISvhoK+WxTuIyKQOiJw4TEMbMiATI/yv1EzKd2N6L4gZuCuLmvOEHNhT
YhxBzPQvj8RCtiFCid88WV0ZW5VS5n0+F7k64eWN5xqQob3uueViwZiKpjehzsnL
I4TsDXmOZPJOKVq1EaTNjnjr7ij03mV92m5k2oYOPwh9cs2i6D0aX1PNerEKjCGO
pOGHyW3yEXYfLSj6C5FC3y4f9SCWrTyCei+SNBEaHTQ=
`protect END_PROTECTED
