`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMQiXyAQyCW2l/kS/sj0LrYjmf1Rw2zNznGjzoRffqf/C8GllnR2weKZS8GBGIz0
vQe5C2h5xjbBPIYzoecQyhICvn6q8NRedsWu9X/QQWWDi53/FrMTgsV9worp/nXX
2w7fGMNAUVPt7EDPglW5IlpO7B+hZWNnMdQMNJCdx8myJJ7nciCme3HV2nH4RUqO
xn2oLyXW0/fHuYheagJ0vVic8wvhljbhyn3CjfesDXj0OsQ1sNPRpSL2X1iVbkeL
xdOZP2G0lzQaox1lxAGRe3e+HATwFcYmlq+dbLVNfF8wwLkrmZkpJ6CUUxIRkhLo
DZQGD8yo4fqwCPAM5+HfKBDipNiL8Lfg6MI6E8e0dgxOXyXi+ag49YDwg4MS7S4C
`protect END_PROTECTED
