`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9SE4ARCVkPZj0z2teNQ2TEMneTh9xHMFRlVIqReV0s4py9w3LKfsNHIFyQZyaNV
IhBkJbG2vZJCTNWXFUloktA1xzShIwQahHsNpw1Xv6u+6H6WQzIrsFx7WLps6qrK
gTjaV9RdOeHh1KFA8b3Gh6jKXX1lvMov9N059dqz0MTcEwA/0jEMlEiQzrj4js+/
ucq5JEFIv9jcnmbqRpI7VQhI9wFCLv2k4Ki5be9vr0jjndfDfOuBQZFPUJVNK6tm
whyo6DtIcIvsHXJUIy0GnRIbO9J0OsdOx9UZwcxXUhcQIe69MDmpGEn1YfTym9Ha
tlMIwuYMroUSnVbQbwZXoVzsHFquaU9jM+mAiiIo9TYvihVAUlB9MavzQBHihBQl
pPu3tp9t26meNjc8SbwI6hozpC4QnKZJupOI4E/tI4eL2queB88jnjVM7hCnBXE2
`protect END_PROTECTED
