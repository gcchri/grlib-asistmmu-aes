`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WcsIkWFZMWE9lQuZAjws2IhTuz/5sKXpgXp0g3j95pKF7atWtejNvZHyNyUDxKue
gZmLqsiErs0Dkw0ispPymzI8K4Gs/gEjEUqyk4P8eHDUBqkTqQT/f2nE9KE3HF/B
0lSHuc72IpRuP/bHW3TpB6zuT/jHsgzp9rXtcTgNv3LdqOmZ+3ATYCCZkenULydO
Om/jU8uN05yHF7yQC8aMxaloiBN/mAS07XRpUKe+BAc0Ky0sHdOvpxDGZROno3CA
D0coaoEt/lmRX8HyV61fVhNPUcl/m6JRTRntbZ+h2d84kiK4CWyDhJQF48JcwwzM
hNCY67Ucqo1Y16xiCzN/SjLqh6Qnva1DkZMvqDsYIBh3EQL/hOXPISOr1wS1zYCl
6LfPRf2IS8e5rxa92BA126JIPdMz+eN7+CWt6cTU9oqZLKc55SNU9aq4F6omYOJt
YPqTqGhcfBUaaqgyLREEeekcIoRxX41sMCyUtHYpBa7scO5XveHLPH532kVGxLu3
iWsRUT+wIcACOyas0yUAj5b2UmCXGqwpAqZHqvX1RSx/oKmMPsZ3gfulSureIgxg
cWoy+UOcazAu3iN4F1C9ug==
`protect END_PROTECTED
