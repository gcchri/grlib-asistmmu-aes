`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z0GFHtbVB+gVOT2utgc8bNRZGu1B32jK78emAvXCxgWTqTFr1P77QkbWSGLjJLq4
vTGkb2BF0vFfn5DL8wZUEJ8MjcxsJEqCGiZ1ApgIs0K4+FUoAWY8OFjEcc+A2VtH
q1wzQwMcXp1kDQLcaYjSdpHFWoEB4c8nbs5RMBlI7JMSQ6tuTwMnRRrbf9bjom1N
VC9GV9FNxKw/3koVxrB+NSk4hfPTUQCQNjYjU5OCB1/QzxxxXszIEsEWyq+bGI14
ybn0LxRqf2TAb/R9BZoDxbiQ0m3iGVNvn/JRBb+8s1N777QbXVq7yoFQx8ZbR/JC
iR6d6KHjT8BPt7wNBBquUJYydJ7uhd9u9eHS4NVmbk4RDIAp/OMf2B7Jz3o/q+3q
4mNm5RUol9ZVwwiltbgIo0JdffLK0JA/9c1acDt5O+6WPI2q6xEK7e+1/snoYXXP
gCeerck6ORhD/bfUZ3mwiGUExUGZTw+9MQyThhyvhmrCVhgdXhYXmPqgJvtQlU7p
FzVhwqR7uN5K2/QLvzo5cMNbHqYbVSUbEiZ7RuoYm3MquGf35cXk0A9ILlvMMbcq
tip0VDJwT+IKcHc1XAMVwg==
`protect END_PROTECTED
