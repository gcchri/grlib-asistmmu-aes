`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rp71/jsN58wOtjMZCuP+lCfIGMp2nzfjCKULn7eiac3tRG/CGsn4uQQYgAUBRamX
cI2RZczk6EMNXYsKePrU//q7VlKJEj/tjE0OCnAlPDFgQBrvoOUU+Gct5mPW7Q3i
/XWJP2t7kBs7iy8m7ia3A9xXZOaiBzmRyACcHUbnL7dPGaFalVeoVyWN8hoX7FVy
oUphlxULH/1wGf51K6CCgqruzkCoGhobguwr8Srs207HSjB3ChefHilwLrCEFIQW
nCXPp1ho3jFQukpx/Z8ElJ8tgp5INo/Htv8loWdBc68lUhubnZPsFzPdLWu4A4q5
zQM1ykuQweFC/umfz4z8/fp4Gb1uQc9X03a6hnjKzvBMFZ7BKbRTy0+SZjaZQMZU
P2aw1pm1sg4/YvxC0V/xfHdclz4WKwRhLwDBi1m+/4/nM1cHdorG80p2Oj77+hfb
s+1gPe/ztFGZGff0QqydeJeV17MBipq3WdhrGAeyzuhMWt9S6fEZ6kXGpmB4tBEt
1JIuDuG5yWm/IlECs2Jj0TUoavhaVvk5iQs1VWSYZKralOkpE19l8f5FFG5r4G7s
Hp7nLA7iiY0xc9StBfUZu5rR9JnFmXADMc+oOMG80b0bPpb5gNTKn5WxyRavVi7t
AQmB2lExVKWm2//zzbY1Yg==
`protect END_PROTECTED
