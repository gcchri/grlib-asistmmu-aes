`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ys+gmdWHd1nYUb4+lcaFLjTRz3tVTD+Lms0SRFGtBd1JTnK104HByidlytlLLdb5
AN3W5LaBg2RCX1z9dpz/u+h74oarn38UgW3aKQFSIQmp1d7z25RWEtWXN49WPqpA
nrLyTGQIrbLauv5ZNF8DZHf5a0UuW9sQO343Ss9Dyl8QzWnISAwb1RiRP9ssxuk+
8wpYUxV17eVf3IJ4W7IM8OFkrriGaMj697WuJNHIH348XeH3/2h8uJ9TTSRRGWR7
Syyu51kGmbOJqNSYJ7N6mhHwLqjXFPjibRRW5JLJcjQ0QZMgjuYnSCrpYF7jFzWB
Sodd3PVyufDJ1+M4DKg96Vv6wxwXY36wt3acYHoKgjSONrXva4dohwwqlr1piFxM
Mz9ku6sCjW8GsjMJYzA7q3p2+muTipK2PST78A+8zWtY8GRr5gpiLlOfJdmsh4C2
E6/MlmHNH/6Sa+ekwTqJky2FXRTJBe4g7N79PZeZ+wLBPB/KFbDjWzuUKFMIAVEq
u9NP57VOrgXp341AqJbwF9VPT0XHTJyw/PL02eWzD+Mghrmul2bEvVuATETzZoGi
Qke0dOHJXADpWiUmiv/m2LhMmjwH468eWiAJVm7wkA6Cg15P8poq7fX8ADZY6Bec
2FLBcYTs6AZG4fjn9KYdDw==
`protect END_PROTECTED
