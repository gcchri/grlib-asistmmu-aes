`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kBgUpyxnXdRYFjl1qRjeHLh2YSnLQNRxSGohUTGfHuDfixtt5rlLuJDtrniv7S9W
SOeqnAp9rYjw5uwxThEjQuMGDmgr9MIsEY3Jhr0jcZVKrolz/yMyeqsSyanV1wEb
8QEHjsS6dzdzDmPyzBs9pMN6B9zFElgqUWUi7AHqgKuwibdjeYR5Mf603eI1JEv7
u/QL7LX/XiHACHovBoHz7XR16HZQs0mr0frnMyYjtkid03G/aZ9eHyprxmprd0o2
dY8IMduE3a3CydCNBmwW1Pv5otEkERHRzMLMw5u+jxa0qprjt8N3u8+I25AAi7Bo
HiEQdmETDXLTdpdXX16ATl1SEDM6BDhjyhXf5suet4gMlvkXbO0Z3ra1vDVEVytR
LzOa+Utfs28AOUNuK0XzCaMW/p7nlMlRx+XZKKHgGnAjgTlt1JkLSIIBX2wPuIZ8
UP4FAp0pZe1zp7+/B0VSh/okD0eb+jbzPXGhhDIAFL12HuQzzyfjM8CxeyVDBZYL
`protect END_PROTECTED
