`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/Za4P/2zOVo/fzxIZckUe2UezvWHEwXTroLGnnNUD9ggcuHH46c0YWBpxgpaMGn
SHqJCNf/Bzlj+kt6Ss5UNDH5i2WRNEgRR/HhT6/jg15W1S4L5v4XFaV0uArCydLM
3dFoCUtmrDLVbv0EtN3fFnReSYUKT30Yyrf0C7neoquRitI31p765UIWjk0byqU9
LhFTThmFOSwGgvM2OPVlZ0CeoumayxZgxM8/KLwyqV1lyAojPmvcP+bBMk93xlPd
S51aAmn6Pu+hudq7S47hKZIjW6mEH41TNz6O33f+lTFwLlGgKVWgnvanglCAK0G5
ARBEpvtczHp/fUH87jgt3mH/jSa488vjzawuS1duNF85xZgdzDVoIHvMwgSyOEDx
F2AWxVojZOQhGQ8RYC4+fztLV1Er15J8h1BdrWvcH4FnyNYbgtCuc1i0YGjmCR1u
FhCwI2+HF1xRBp7Ve25TtqvxpagxqRjB7YxgR3Cz3BQOXjsi7a95Gc0adesQCFog
BZJ3ze9rZIB9SrxxtMBmHiinKLM7zhK21Ob+5apm+9gDm5uSABP4aMZAealceQq2
buS+NSZJaKisiPqx8z4phLD+kjVGap/uE0FosiJ0rVM=
`protect END_PROTECTED
