`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
STAdqD0lNN4dwioblyl4H2ML1c2Pno+90aPROGcflUDFUXVDKB7jrfKVL8w3q25c
dTAGOPWgf4Dxn8PD7LmPllGTw9p30Zfzwu0/sM6o+cSqGgnDgy4VvwDYl9Ps6nky
K6v9aKFi97vCYqlKuR9B6uI6fgrk1yN24sd4s9jvvO5+uSqk+c1dr6ve0jH+OHVo
ADTNQnqSKsR+rWUIVHyqkZ1stZ9chND764ZOi782n0iIiyxCJKdPAKZK7G7fJ7sV
v9O0AJ5vq75k4uOQN1Y4smLda9PBApOv/ILB0/mFKEM3lfJbzhGPyFsAgE997IZQ
/iVZ6qYIL6nEweZgMRDbEgB8ZIrOycVvDUtqGJ1Hu8DRezhaV+/wR3jAvxrEB5gX
1GVowlr80QDdiz8wt62/E+CFNmYg0yIPkpzF1+NV2qvOOh+N3UkB7qx3mbqXSlze
mt1Zm9dCaWA53bkNZyFSxKxDxPyEVA60bpWIFixvwiVP2IRbI905nBku3pqq4uOB
FsUYfzrYJXKp348lGc9YGsEbRr2tVyyasnq9uHBKOg+GH0MvwWOKtdNAnvGvPPPs
k0rfatNR/O9aY1iVZl73dcbLZxTmKxrovtYPIujW81F/1/TEc9YgLAoG4la0gmkX
QN/EyrvIwEaAYmWu+RrFmwXBIOEJ4hpjUi7MhwupsO68zsR8EsESrIr1tup8wYyo
VIUEBijUGFWsyUod19Ua7yy+QEG+yxKmmAZAOxgw0HzaENyLX7LB/HTSLyyzdQV3
QFJjudkb+XhGt8fqLwazI5zL/keHFAbvnehhz64c9R2HnO2VE6osUp1fOJcVwoTd
mj12YVEfKKxaDcu41bsiuEUksl3b9sNVf/1Mj8fl6UmGRVesetGl1uYEomYEChmI
J/dRv9YDrSPBcNBYTxkKN6735A0aE4W5UWb6QqXmffpSTCLEhEsZtywh17j293s8
TyzQGe/TuCE53jj5BTwZhd5I7YILe8I2RK4X3KW0oADFFYKJ3RiPUrnc6OjQIYQm
466wl1glJnVA97NXneTmjh/Vd6IaTCL0qgTmVFxZdmcFXEdnrmp3x3nAFWg65l3E
xDAhrgw2o4szm9HECkRUtBWVhBKZattdt2iZNPr2buvuxzNFV/4ftz3GoSJJFEMC
+Jd/jfzb5VGbbVSFHD/lwHzLrW5mzdcp2m1Ro1ixk0qH+QgbkR3IDWQ2HBr5E1m6
`protect END_PROTECTED
