`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZGD+h2PPF5n3SjfzV7ZJrCiqkX/x5gLv0Jc4GMwoYfokKL46eDxwn0FgqOgiotF
0Bo4cv3xA1A9wITAvjMOy74QhvL17Vju9JZ/0reS48OrwWDjDsKkEKXXAny5hRsg
rRvVmVtbExgAsnuZoHP9dO/r+miLvlkSI8ApNCiCZnvOZ+9NI0xz/oleXIU5KwUx
ZhH2NVXFNt1KrICsyNcqgZrI97h3T6PP2UmlDCPvUOkK/pdV69xy3TvBFvgzJFx7
xWhb7K4ChGq8Mmfi3Hv021iQ0SbklEMGAdwkRDPts3As5f6EnGFzIAQJ1hTkjGgN
kFrBU9/H5nV8E0n8EG6rn0lZtLNI8Vv8pX0STUwwdDo6ZisbH1+delME3xTefth8
`protect END_PROTECTED
