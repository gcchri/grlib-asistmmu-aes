`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHImwKU21RHn2/AGbBqhmCd8hoIn6kYpESniIO6Lx9Qup9R53mqZAeKNXlu5uMGw
+M9azmqEK+GDIrEW8J24Jbyuex58VofiSorVU+NktC5lNed9kjVijdDkM2voOp9K
NfhraCODJEJb75tRX1ZamElNzQgPkBwRGORYcTCROuJ1jCDPLZNTtVD9IZzm8LeH
JrFOutAS+wp0nywrpYyWk305Y8C88IxfyI67lBfWST3zUp8M0vleHePKpC3roYVY
cWsR2by5XisH+nIkGPLv1jrJIj9aYMpguSY1wm7HPOabPSKRPEDLb7vz4cnkywDB
1vLiLymh3qhJ6fakcYYj5qofL9ZFBUy2ap3EIujKxrIhmrC6NKeJADuDf0oP65Xv
MJ7vrklJy4ylkOSRWcKpDSusRAZTL/Lsf3ug2/oAtO6/rWVw3q3zMyMx+I1pzXN8
K/Slp95eqgCxydekLMuh7dWzyEX74fP85LanksS7Q+NsSkYNOE7AA9q0ewVNQ3zh
uwX0Qtl6uOJAoylCGwkIYNVsvLWAfql70IK4sHwUjQUTrRXgGPW5iADOiGZZlMBL
aAvCUGBIlL9Hq+6OQIkj9S5T1wk2lne7+hNhGkKG/Ds3uH2fVMg+pbZSCnc44e/u
ZaXQ7y+Ej7+2CgYr7QwsUq6SFAmaJheG7bABQBXPcP3kVoAh/M4cDB4JtthwGgz1
hJZuOb4hUkSPZ1ygyM3exjUDz+IEFSASO5wXB+w7AtR5TbAlNQExbmslEi2j6S2k
jQD9i28ZhukSwVqiPKvt0l8IHnUTG7aOFRd8wf+TAWmALnJPShYV7kqVn31eU4hV
tIVwESof3vuBXJ49L9XVNddZPf28NK7g736/9FFLCv8SrO/zsaXLbSMHcnZ9QXHB
xJrV+JHEOFIxyIJxXunJoQ==
`protect END_PROTECTED
