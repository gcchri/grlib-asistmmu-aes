`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
myJ+MSZlvrD/JCpMLxJ/QC+rQyAMXPYrfU3gVMCSTzRiYJ1e30xFA9Z359q93LHs
onstH2GvFVO+4J1X14ZuV2mzkknzX04ot0vcvf9ArRTiAQrfXANJbQXb56YJ1T+p
jtxcFZV26ylvisMW/i9n+Poxd7FHTq1MCEW8XuRbL6dL4QdzdGw95kFEATnWCGc3
i6HuHaJvm3WBgl3TonPpcYTJZLbJiNNvJp5ERAJwG5AWI9k9KjP57HQ3s+QCLWyz
DYONyx3P+TcIe9j6SCuD5ow4cdyewg+x9zqF5GuUWMh2KIiO1cZK4U+UX8Nj7nz8
n30OTR+NfVwRtSuEcNd/cgboxD2n+lcXOYPCyHb5zGGZMbPVE5s8SzO2LSXqbszj
bhv+rCIGtCYOHZYLLGljKyzJ8JX25zOorGOMxCFt/iIBCKmOZmTYX7+sZBzSlQfS
BBBnBcXN4qvf5zRDXAsWKLGPTfxhuEWcbC4CfcbG2RFK+Rhfop2N010cKfvpTvi0
`protect END_PROTECTED
