`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MblcXxkbp1S7QwPdyHYq1EUcGq10pvuVaWfyPFdA+oZOAxGz6oZ8HBvftHJstlOx
pF4AzLs9hS+FLLYGfYWXj4khl2d7GiDk+7TXYrhPMyVQZ8bddZXRf4BdVXxLj0DE
xFR5oHbJTn3XXTFxPdJj+v32Pu4goBTobMQdfqcZ5QR+4tTa8P6Xzvfj/5lF1BYo
g197mCmFTSur81HSBueDBFsIxfJaPdTnv91nygwpeFdrftpXZDnT3BvP+iq/FeiJ
uome2WyglkSaNAdV9XWtWVoQpU71EzFuDCNSA5w89bimvd2rdO9rMgImSpRjRvFt
gAIzLpZIq4QdB2u/il8xzXy0mYiSBnsLN5uUZyiV4nYcrtc+tMyqcJt86lj6CDiy
ecLeLyj5CUJ25Rdhfs/g4RStdLCYdupdaxE/kcFHyzfVTIjg5meItMhkpjtf3Szc
`protect END_PROTECTED
