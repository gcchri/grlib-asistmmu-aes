`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bf2vzMdJ19cPjhzMyioijijNfO1z3zx41CvrC/WJeYy3qtRWhWAkCvunq53hYFr+
UBRdsZmGRWmj5GV9Bmuh2L38dSnS1/4PlfBTCeIbC967FlEv3Eju+Xw6KNKp+YG/
cM66hfVatn5HVn4YEVIGe42VCjsKa/CVxpti/EyWnx3oz90yG1RDBHwWN+D49BOw
5xa2LBsfB8dtRel1bttSmcEpGqaDUDvBPPXj4+iUYtxGayPW6SsGNm7ynTmRpGph
dTo7TiTYcPh3yvaCKaN9HcrU8vREdCXJVXy0ulBhRDL6M3Of7xi2gRrYtLowlGq4
60ue1Vd27X5KmWwP4U1GkiDbLPaZ/o4CMo57T5Vy7C8Ll9V4QJr18GzgGrcv0J3a
XQW9Vfog2pourBxYIiNSnKtQ3BargPI617xg9mn3dFc/9mELg19EFgjOBD1sQeEs
UOrw6wpI8UktC6HyfN/nIAFymN7BUf5efBRcpgbKbVUxbfKm4yvahcMCUqiPEmPJ
iyIEaKF/G+kbF8ZI59cfxyExVmmZxfKmOEq96hNYnoDRNkIFVdsSnWAN7I/ciFuF
jJxoEQNyZG7/220qCbyiXfdrpJYHK+bHxnLWj1wOtxK6IRVRScw9Kln9CCAoo95p
4rHsKmZJOz4iWqcEGBhVitBZA2wub8p9y31HWLqEvjDqgEZvjrAaf1QOnEkmKrNg
tsybaBaIGwOVBTdQ+LQoTtocHHaEbYSWW5EKQ8DoYqKPU5GJWRFpqSetmOOxS5zc
ZRtkHeTdSl27Z9IYcYDKHGpAIWZpISz8mUsQdxZojEVtNZ/DJdl06NCVNNb9cKNW
ggck5jAXgmr64R7uOfdklo27pvdU2OYb7ORwbafKBVaQgB777VJ6RrQIsNVrhV3+
UmE9MWxf+p6N5qtu3ifUBw==
`protect END_PROTECTED
