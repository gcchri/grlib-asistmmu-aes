`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jabqOKJcEWLeWUanUlQn27TCYhGsTCVtaFESrWDvJpfy8KULLbDB2TfCofIUwyit
aOBPeu5jeoDr7bSCcXMR0H8bMOA3x9YlLWo9/vZ1jnkclRlscPIYeh4ojeFZ/p4l
+WCn66NmIdxgHHnuAYP4w+oiuJBScfvexRjgVqPbUhMkz43BySGhNSYVIaoT0qHZ
6gG4I5csuGE+bXfsSth6wX8I9iGAC1OQC/EQbsvJp6oa3CkUQXwXX6sJGtPaBiBc
1S0N88G3WLK+kXxKRLqpwUTWJG80T0sOZdIwYvax2p7KhXSOYECPF6hMDRKocC8G
`protect END_PROTECTED
