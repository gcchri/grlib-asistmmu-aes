`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
esTwPYxqMIcdQHYU1euq827Olj/7OXrECiB5nTUAMokx0uV95wPoU3iIHhl3ms6S
amUMxCYkytDZQLOSBUd/6y0CXplsvrxnD40Ps0OS3y1CV/Ud7TL3FpiLlq1d/Tie
s2n8CbjduxJl7d5xlr9VPnUp06+IVcvvitnxL/EdKblUit6PUycT73NnCs3Rw+KZ
CfvrclBTeLzjJnjzQzzk9qsEuDRvKVLBeJehTv8lMtDF2saj8F+YvSvYBOYyhei4
LW+psp1DqXIN+ueig3r/fqrL6DDmQd74FSSVTiO1kZhjYpvZi4h9PDd47GmJNKWZ
UkrcU3YEcL5bEA4IqiFOPC9CCO7xxpBO0Ze3OvNhULKco4xAlcWOpmuAUnku8PZ1
WY/aklupJiPvf8azNpqtzfPWPaIypisZSr+OoXrLl4SLE7uWztwrb5fsvqD/rca/
`protect END_PROTECTED
