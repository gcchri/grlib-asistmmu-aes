`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2Rw7M3pVVO4b4+Aml/ie+4+NeWByFpv0Wp8AIN37DJZinp+y2pbiMXI9ZN1jYcK
BeGwq5QspseqdhEms3mpaW3Uf8Y2um71m+/2vNXRoEV8NXOScFv9fSvYMO7DMYym
gFXDl5xE6P7iNn7PlfgukfWzx28IfHtAaPmMmqeWV3RP/epxNP+azcYQHfr2qvQ0
zifLRQ6WOp98Tfo9YeSphXGkUrKxiLQ8kiG1UoCbs+0qH5YP6V6mj1cTsp7WAI+Y
IcTyyPXKDIUSWMfJ4yZ070n4x0YEYnzJVqyPmQb3J2WZ3KEzMSeFf3mfZkl7lnoF
S6xLC+M0E87J0WauDJhJA8rU7e1/Avy4pcjp22t3oxRHY1h1euBrJ+sxixCtIkfn
0x4uiQRQKt405acGBfnbfALAAozMpNxVIosyOual4G2NOHKLPFMpVL0QtkXaYxJZ
1LU+/Nl/9Jg1nAZFlsgkwkAEtRWC56gPpp3p/YlLTrn+0znipLaKavh/1oPL14cE
`protect END_PROTECTED
