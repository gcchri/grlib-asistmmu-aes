`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j8IGClLv6XFEBuSz8XxDFplFfIDn3ToZMttOpcNRhCvjUrBz+Jn0R5QubBvLz6w7
LJKyFymRZ2RubQmOYb0yf500aiiUdBFtUVLFYRlblc5Ma40yHyLzx2J7vWWSbXjz
julB3Z2OK/HelKxaeW7gyZc/uX2BJ8sT+zrzWODhWjOM0VF12vRkfAH3JbPVQKYt
ewC5y7/Qe0+CO7e3JSl0DflLxDqHVXx2v1h2X4j9DOvOqopvL9JZGSCCysSjnEyf
I+nITp8xRd5eY0fKg6d0fYFU5/rARMserCy0rH18tIhFPyeqAhBSqYz6odUMJrkz
BYid9f7RCG/RozJHFQV9jVtO0tqHES+y8tDrJ53l415oSo6CCdI3WJc8e9ArMBzr
mf6p5q+2fH/J/47AHenVb2HX+NIniLucpVeLY8oc+LtR7CU9fJ+BQfbCpuBj986A
ziIc7qZkZ6iwZ6mBGbjvRu0mQS051O8JtWR7icN/Zcw9YMas5stMwOZOER70u815
si951hBlwa1z9hIDPfM0mwtZMWew0Ltrz02OsJPcJbNjezc15j7UolXr02F802Rw
ka0+aJVI4emAMBNru/PQecyvejymIrUKv7FUr5aWnIMoOInJiT3kR5xOb6whyXBc
hdB6s/ItjwCA1CR0HANeKh4A6xjCERMoRLzdTXdcUt2YWSpFgo5X5m0Evu6rEllD
K2jEDYxQE8eh/Y+WThuTur5psWoeIQES509197JDGPXfwsDwbSrAkcvHWJvgv9MO
b78ZBWjnasK+BlbJdBPMAqtyktSmcUKoEEdFaww1yrOrUM0yUqWIbaadaIsXmT/V
Bh5KDSuxiIcedLcJrvg9BgEuSc6ROT3s/3wAr5VjQg2M4k4C5V1oZVLUC+/NpbQw
MgZeaQb3M9vgF1I5ofuOImI3wf5fLnCxYpaPOMm4Y1FoNXpkRLbhlPGMI0lX//En
c5MrJeOpvKevpPNe4qiDB203GSYvvNKfzfDNsh/Tt1AzW+0sFzSH4Qy7qBaQZiGP
iQxzmkduZiVyfxrD3PSAE9KChdidLRxHP0B0hA7y2wgclzZ9qaNRHOD+Tnr5YcOX
bc/kes3qgROzyG/OXc/N0hhDBafc2YcKOrUeQn57/3q7JAJtDS5eFKoHHhooK8Wv
MsnclZOuCibDpz0ypoQK9uUnD6YKoneK2T/rRZAfgFtqxeh3poAkTZT29rkKr0rt
uC5uBqx7iDyt1Twx7TIKKxIQgJO8f/byPwQaF8x43SgIjaZ6VWFD9TDqzarn1b9e
PGKG97TxNcAdG0sVEPZKup5fS1flSQ8T2nnYnu5g/o8EPvqKCQyn3o8BhAC2X73c
GJUmGhCJLAQgbUJJJmI07nEOkfNgUyotuj0fvMhLQPPF7gkQpK/7yzDFumXw1mOk
/AWEdrp6pLcja3DPVVaUXVt4XUhsV9kP3iw6fO/a7GFBaGzk1reNt1AAm+Z8HFwv
KZ9JDmAJuEA/EkPsqjQ4lh8JT9YRjD3pEaiStx5fdVXX5QOeYWKNaKG5fK+5Fs2T
Hg5RfF47IDNromkP/aWlV2pkq5swF0dAPdowaCzjs8UtLgum49lK9XUs5chasbu2
CmHhnpPdaLiRvBxdLYweH8+031BsAN+GJ74clQSylXmv/rQGDiUlraqubNuLafxj
SzeYCC2NbGltPHhTgrTGYVkUmREnhCACI8+7wVTTeZSZXl8m2IRmNXzq7WQUob/J
Hdl/KSvYwdioAkbt8/MT2MQqshlRtA1YDDrA8TLF6H7ZSTHwXd3SKN61M1HUKyrp
VArbZTfI0OECfKHh9hqULLfhmiHkpOPphwwUhdqVuDU1lryCiCWkxO82V18ydXGp
Okjf6LlfY87i4zX+wqOS2s6pRSOQ+iDN4qx4jsWrAoXz4FwHdaW9Cev10TG5v8nT
iRuJC/qc17UrGVM9YJFY5Ogec24ioprx5AavyDFYK0Mx7+JQ4zufKAR0IddjllD6
JDQUcbOSi5CrJEr2GrDm4Io5Co9E0JcIQtHNuYK5fjGfGJuqjzNHF4vPppkRfSlM
vRQLw3tFfHH+57ASdThs1QhzVLLdD7jML+U+/FD/Vdr7kuJ8Olvv+LVLMDRraVoY
SlaNFMVOeOW81z6u7AVdE46YA8gJyqrMdLCdqAJ0IB1nEXK96XiV5HMZrAAZD+3y
+kJN4De5xQYr7DKIgUADVK3QiOPGaCjJf5CGy8qRfhyuGal6Shjf5Rb8ZKAPIrSR
vy/AaspfO6dypC9xsQ5JbwKZ20PiYNsnrbCbIUGdgt6jAtNxo5QPYGd35IlyMGwA
IfJy4WX3JwwNgQ/81hbqSjW9oGk+/9dfr4k56cpPABOlDDd+uGvslLSwGuGJqH71
FpNcQ5Lgr3nRB7Omz6bUROIgAHyibOZwfDKwC6MhCm4w6ex6nl0Df3zPAsk7ux7R
a3HUcXyv5D+pPmw0XIcU+0/5y+UbF7uTak9zskYDMPcRQlIBmG2+gBqMI4F3J2bL
AskfxnYWm3biuPT4ionkrcYNT7mhNLtHvdldFLQ8jxnsNJX1ks+efaqVcJE8esfr
wHdgmiRF0R9/whl1/N6Jk5R/ZKKY8bRUQX0qH3Tc2yEvMHmxraxmy/Vhqu2wt3Ue
GH2qyfb32rWuLuSmR0WcRGlP3+VKsezsZ1gULaqX5qeFJXzoGdpKJ5MNAx9vfthz
IKMTPQ8Lxjbjw7tsE4zT10ErHYd6xqJiDS9xUIcX5r1BujIoYcw58FWqlPDFoPZX
IsGDp3ZOxxLYVUzjwLs4ko1aS8k23HxS5Q563IdHMN9rblIFZEKfmMSvLzLiceuU
RNqvz+qFsNLplDut8Lf+lQmJa7QVzkDEaHbFF8H9Zo2jMDDpBexYzEleS/kgQh90
hlsit1vLKjxRc7jJrbVWMzciZheN/xY3Aof+ocLWaKWA2Vec7pehOEkU6dDLB6H6
9hynMYFpYwVG6N3ZbBTPs3NhpJyZyNJ+VjdPr3JgMgMpoyYapGLECRW11izYnw4+
UrYjAfLUCRY0ifM/CSVXkfLXItah4g95i7tpaozc9X8MCYdL8rxNVGNRxwQtqDtp
8a/EnOoZp6we4QCfQhOFytzHduTsnQRfA6T3wKSplIwXdmnG1JW6Fbes09Z650wI
wgsmmgNsNfGXljuGL/Sx/vObhb6hzH1h/NriZ7B6Qis9M0fniLLbj5vbM2eagrT1
gYvsdWbTomBn4xME5KqYlC/pjM+QRoMgM+zQ1ZRVY5bMNb/aMTnNuNf65XDuFGKK
RnsFbEh+SPDuxghUCwGPKZTNM7Jdmj6Wggux1Fu9Rj35GnshwjGvd8zCgJr6E0JX
lA7f3tNuRD9tC70y1g17lV28mOyaTrf+lOwisMpY66pUNsGMe6/iBUiE3JdVuX7T
Q5cX1a2dSSIbsEJnUaArsFWpjzuVQudfhdRT06Wq+ahfP/sdqInsB0vAHX01gDP+
iBE0Xc1ZyRwS9IKStFuvCtJVEdJO0kG+dza7CHn+tL12MymOJG+ENO0Q/0mWesAf
ESI94bslK3HErSANye9/k8STUn4Pniecb0KbRNf/aD+0LpcdHYEjgg2vNwi08bQX
EZ77bTfuoG7I6gpwfOqhG4x7Ahc4m0xkUkIwnkPFQP3Q8J4rXSyEH0iJ3dVZYcT3
giNB5hol6NMIkBr3B4QxoNEprvJsGeg/izuWBj4biOwNJ+oeoqt8Adw5OzFAdw3/
ZGlE+OEg5Hz82rXE1t0G9MgXnrrC/v1PWNI62cscnabtOTJSbP91DSIg7TXbvmTC
Mm/Q+AUSiWZC0OMd7DAARmeiDTNTOWho7PrBUnhqkZPnpAPNzRHVUdIDY+5vnCRo
CQmVKKH5viYvl+5yoXro8eUy+L4K9r0MyE8uSE3XnSX2sFeU3Yl2sRJVF1SVqm9F
2w9GTsdNNs3kyJ6GjjlJro8jzVCL1YcycN3CrvUlJQ/A5KO/5bLugA+hi/2zZobp
imlXafPzwLqjMNcN5b6kLKts6Nc2uDFo1pG3K+JDy4Il83B5lLK+SyoXWOtvlH2R
P6i7JazMl4+1oi3SZJfxXXMNDP6vummyEFpQTLg23vaIb/KX9pdcd6v1UOwTNsfe
S8iafqLsARRKPBC8icyj10wgJil3FdEIJYlk2B40v/KnU22rdVXqZyGw85ugD0PA
LcV49hA5o2Sx2npVkd8g1PT7JTEOg1jINTbTHuiHvjLzRDWY2hub3RJ7M9MNvwSA
xIbE9JIIbeEy34jJZVRYKb82EEJVHq1fK8uC4qCQEIzEsh3wAhIXgOwT9TrEfq8x
4jmYKQWg24C7Y6YK1Qs/Zzmwhe54H3DJ18qbz1Zv5QBHA0gW7axsFEo0i8uGBPvC
35Xc6nrxD0+0Cek1+bg6MB+bDwygBolhJo3HS6q+6E7oghMqhIY3P8WPbKckEyFi
+bvsRR0vKI1icOJxGSm5DRAJ9GkFXole4KVWjtgoWfDW4l+Af68NkgRALzH493XP
7Ksc3crV8zsWf3CmCjoLC95epuKc3G4xAKRAygUaF3OkwvkvI+9TInwGr4iiJQY2
0p8gFkdtWsOPqQJuLWol1GnAgtCVtRLzUuj3DQBqQYJ2hwWmIqJZ6zmGqvhNvgPR
ta3HEJsSxQuHubHtipDiYQA5K6xkq5XBxAVEqZlUKXOXWKyTT4DM6kdUwyZDRz63
d7TRxZvIhYGSBT30+Ud7+dr61E4cjbe0iqxnTuZ4pvi7bhB4JGxBvnVq22QUNuku
Ts25M4jJ4xSlGkOUQGQKhl58K9myHqwmdAKu/oEfHFoV6uX8eifKEmOK95e0oydh
xJrOy+WuZjomsd9pWTYpJFjIHWntETO6zCSj1uC4gQTvnNplRBnwQQ7Y1nKKGEa0
ARfEKqprI5zj8dKFfkUp7cgAaNt02CyYz1X5pxSMpDIdnjqLgkE6gdia7f/UeEug
vmCqOEWr8t99ppiwpjaYoB9+q2FQWrTW1+M6qKyFvGZ71JwyWFHeyqjeEXDz5C90
QhJVXBUKSvWCTlMLjm+9bXG/OtYTIW01TvfjayEMqGJS/kKCmQ47yHlLNtF1S5yx
/75L+YNHK/Yh+mRhu+LxDB7OoOx0Ue2cY3BObXsyIlK2WMJSXFrXNR9d1lokSc5W
JPmrwQ8+Hjks/oXCpt1yBz0G4pntfTuW9/2nuVJeBdA+JLrKMCQKXjp+luEjJIZU
SwmqI99RiMytXEbsJ9XqmzhddaOeJgM8aYHyZ4r2Z+H8zgIHSn1+cV1jggRaTaag
qa1t7BOEAggeZqK6ON1evj33oj/97K5uBsjX7NSGW5nBnpsPbFicYjth4NyWzhSh
mpT0XLPmLgnab0e5wVz7az7klFWZsVdvG4bGyZDa4WLMIEjNSGOAwraL7jMtmPmM
kca7lA4rW78rXO/C312CjdbdUSeVuwnyVGYDS7rCFzIebe8jg8FcSEY+dpcMsX5E
6MniKgGJP5HBelFhr1FrHXWm9So4+zRKM/LG5q/acyjrxveyTFs8mIivvuIs/b4t
V64oPbsB3Ig3mIlVyyjWmptNCwjRIePfiQJX+kl+kNeSTHoRuJVRvL+0i26XL7+9
1aQv5o/pqPbRykIhfzQPME2mzMdmlcUKvkbCSF0+fTwuE6DcYVzIQJTqQbpbZpM+
ijMJxMEAnoy6RKBQU4ZWkoiaX8mBylBbRg6nq03tNTivSXIR/6Kuj+QIvaTo+ZmB
ouSdLVd+yWbSwMYwnEqkj/BKAhWB574eWaHSx2PHRfXNks7EJthlGNrNOBy8eHyi
hhV4YMFag0sq61yXr7ce7T2+Rw0pi8C3E9qm7tNtSqhn7sbNxSRbKgxyJk3yeb/Y
CoHnKHet2S51dJo9kVai+W7nY4Gkt1Bb5a/StPjRhe0W7EOm/J9BRorjSuycPzG9
kNXa/0+iE+1aIjGIWvbE5P/uAwIUsX63cifHC60f4Tc7WjZ/Fif2pKW+SuAyHLoJ
d97TiLgFO7gT4pFp40l6no4TNICID1z6nIGEsY0NwpgedSiDQHWWKPfUGFts47wJ
eYvZlJ7FfXQxPn5oqDTw3B6qBz0sSqKUaMbu1dDmLZIl5du5FreMDKJQdp196jRG
aOV/aLR3qvILK6tOqeF4Qj6uILNkOV3Jo3tmjCP2BlE82LTux03iyldaWxSr6ezp
8tTk7XLEl/oP8PKKJqXiV7SBEAHBnXcCzxobaJTb1ciWuJgAqOqH9O0abeO9ub3t
a3SyqoO6jlNUli/drXwptscAoATCEOFNYJnMlURZ8CnIPlYIGyzh23wq/6lftm+P
EVWdQpzTM+qbZN6Tmu/Z0E7DQsf6ne9X4hJA3EfjuCJgtOlcZCsHfK26m1pMS0oX
W4EI4QieAybhonV3GKuck/ceqf7JOAeaxx2ULsMgqx0I/WCW/pcRlDpP5BFlT+g9
P1RLjAUAXQbotFsJ4YZh0qAQIPQOoWbGhGpc6GRC7GO2td4Gh/OR9HRsh2WIlx0e
56hQuk/u9YYlx1BQde808TCT86WD/kMF/gvZX0KFCH8dqcRPVOzj50CT1PLniRQx
tF5Uu70iyhD4itzdALl77J743W2IKEWC00F9SqLzlkCcAQbZdctvmkjTJw/EcJ2G
y7p/+oRJDQY99jL2JD0VnGDpWPUoII5r/JtAu4Xel0h2KxQ+WK5pL/7wZ5XVo19l
rQ/o1EAuaReHQHGTlUVPh0wcNA8Nc4FW/l0T/YBSPdr7vltb0nQUK5ikwTpmiFoZ
wT/jlv2KoFGbGmuxLrKeOBlHPumXdOBlPctpDoIPaa/ulqsT3FYH8Bs6BnUSh4CK
S5b4qHlXfyQt7d1pn+sy4V7Gi9adWT7kcJQr+6i8GQCoKaVOrW+64L9x8tSM4avG
mSJK2rbsvsVVMvYIHL3N4Ldg4FSrT1XCgMjyo+ttUZPpEYmdBPgeVCdhi68dXQ9s
dU7wbBd3iB2dQJfWrrjXLvslXp56dWqlOSM3KKXZy2hLAdL6IcoOZrZsUqxqxTQp
yDy6Dz2HOVhQKm3ZRQUB1+ntuvB2Z7GANUonV3wvWrWx6TN23QQSbWJWnOKbtIne
W0p0N08EzkZ1JRueo2HI64/xJk0OC8sQOXDjIldr8a2+HjpAgwm+LMtx4yOK5a6R
7QGIHWAANsOntTXAo0uA4WqWYjDBkjfe7w6W0owTWfhk7Noa5G3oUqAY4NDKUFWh
NGP5vIv9LTq1poNOu602OACY1Kope64hkCJ11DkdhcecYA8mJ9NttC499/yuYwtW
5eusvT3Mfx07W+sgQP0+g3DQ043dQ9ktbODtICgRgwakWBXPHtNixonzbDcVieZB
QwMUB//+LaVSqbQ/pw9pacvtJt8049CWkdeJ/HHqwQbsQCVSLsJD1BGdBhnB+5Uj
WQox60U58ckQKltOPkuA3kkgx1Dq/LsuL9FKnSoTtXj7uu/z4iqKIuN7p6A5cSKW
rOfukQ0ckD2MYj9QZrxFmI09MeBghHRYZLxDJvzPg0z3a/Ks0En8SOU5ABX+AueZ
SQIHgOWr1a2WJySnv4xQeBU3P9NoqPNCfWd3tp/vCtOEEIbTfNQpwEXQ/1WJunZU
euLtm+QeaGUPuTue/CPa7Jnn6iyRQEj9SU+euksUq8HLkJ9UlghXbcunucq4Q4ma
RiOsCLsHH3VN3UeBI2rnn+B+Q51NW+9OCS7osuSzhzGyx3H2TQUl90HDLx3fVOge
6HTbMrxoDMdbyXnHiM6T+ZQ6Z8wYNtqQR5NY1OrX0TOO2EVcFdv3JrkYZWHmJCW1
0rk7Ur2458uQopYNavocmrZ67Lilv+TrdTnJhxtg4eGwPbeuU/PQ1m5EuN6xdwzH
4Bz3sEZdnIutvAWi4XpvG37dqKg4Z/QJARygwJuBKAUIX41dtO3RP8ieobL78jlh
K4SN8DEeRVlUt/T/5UpsKpGoR8fFdW7zFaNhYPfKMFE9FL8beBRZi4e0s68ZUEcX
KH4DYr7e3A1W/sUe3mwDenLZVNPA0ayTvydI3tVWbdzRmqgzMk7gtVGs9JUMu0ap
BSJNOpMxRMi4dKTer3meGS23a/hJQ6nyva9B1sqD//kZIdQtAz5iIqmSnA55yI8h
zOXTpd9KOjRUHWQ9ANbi2UEiJ5wcZjyDnIUd4wFiK5c7WfFbpk1zVhS9/T3wKPot
kAzPUKzkKOcQENCsCnFEgiriPC7+k3aA7MjLeApnb8faUXWghW8T5ACW7JsFKANU
RL2bs9E1A7TsBcy8teE8L2r7i5fYiCnlVMNj/+xeA3dtarXs38esCF9GCDihJtlr
pvdy+qsgA5FY787eUsO9lWK8foQeI0U6tA5Rrl26BYcCZU37xmzgOSYOjEs9/QIF
4Ts6wgsejNESydwyWUNqcR/kdwf//wzCeiGUY35E+3iskDD1hUU61bAib84jgFBU
J58nWzH0BHRdA7lodljxEkNSN5LUAs1tYPsmWHfMGtX67G55qpQdSr7em3VPhPdA
XNnmsbLacNZDh8av7Ix9IrNLmbh9kYg3VLCCDDCD8Jvotzevafh9SWC98U6yYs8e
siI2k+RW6yv0+eW4OYSGWCoSTgk1kluTaz6HMWfsYGjJdALZSS3BCqQBqnHdW7uP
N68eVb1FHlc5A4kBV4vY8aJvJ2N2Y2Oe940hlL3m6BhhQMu8rTjYy92f3p3KeFYL
EHjg0pJE+NmF6L+6fGA7+nUSF8V3XtQBX5/75tBpXZ1iLY+kBDudZnVRRkc/y2t+
CI2pKorjoOSaMiok/OZdOoDR6yRBJVm+55G9KD1N5ezY3visIIYrd2Bd4bRr4rpy
zreZK+yImJ/LCEte3KISCZV/p8HSPMo+8xPEWUwIZ9mF8SUC3ps7mEkCDQMZXllX
LkGIfvVndvEFkyF6Bblp2nyIMgg2s1rJBLtsbh8ogr9kYO3jk7mipuwQhEFi4zJ5
28Ey6zG/RI3DTs6loV02TvSPJEjRQ7kw0m0Dg1buowODwYS1fG9PmZu5XCEfZYlD
5/a7k5b90mUlI0KmJsr1uU33P/jjHA53mDo5FnNBhcPDXsy8n2JlM1P2DEqg0lWL
IBXxOCNckyNd8WsCIkzKHSGv9MVZPBze7NICqFUT8917FqnEWUH8qIP06vT5ref9
LwLZitCWFWRUpY0cL9ls0r1GTL5f4bBpzXMdf7/qiC9+xjoOXtmtHW1FaZZxozAM
YaRYbUtRrvYlAvtq8I0nqAKDsuFQXw2MzBlVVTzWB562oKtZMzP59Cxz6zPWlygb
qxGkJUK9kkOXIgH0vPxUFIoBxwuMcU8mmY0XhK6N4WQ5vjv8c9/h3XJBSHIoMOyR
fZAqWXsLWjYLnU2+XazALp45tC7KJR+Rro7QQxp79P5AAO/SAozn3kISYgNW5E+c
ntsaSovBB3JlxBQsBhhdf3A42Fi78t6+iQ7fnXyWp715H9V43OKTUZx3TvNCZsB8
rhP83FZr70gZ7wivr0UhDahk0NSbhHlSKWQeqok3INBSmMYL5KbxceW1CLefWXVe
s8FjJ3F8W5TODUdwhPtyHPKI93jq1M4zR1RjgSB0t+rN/Dh1ptvEw+Ql3EzQZRBp
D42Nkn8dFgWzHtooKl/ZPUxia/qz2GcHb/jcmXN1Idpa3udboLwTh+1wVR0GGPAi
iiRN532Xger5znGATYiKNueVSvq0j8snXiGAJ2LVpp7f/DmewCFYG7tLbCVRHT0o
8vyazwWqRVoQe7pTh7QKSfNcB9/BwykgPNZ95EQFM6hk34tvjpIGkOCbl8fEzmST
ByXZjG3h+KC5J+fCn4XjzzXLGI6fJnyquFM8Gj5MHGYaS9vZxgwWIo7EPQ3XD7NO
CSshxiPEeNqFvmKbAcnhVicroRdSHb2i6SvNPQiRRSXhgQX/lM8UaOTSUwnmhcjl
78Cd81ESlp4ZDp7GOXygQV27/loK2AO2av/slH9EkEQZ9rpG7ln4a0K6N4VQE8SG
3OgbFphN0DQwxfetdGKroOR58+5uQA4UY2aaBOLsw1j2nVlDjdjatZ73xgf6561q
V0k2u++W7tG1G1R8rdR5bbHClvCi0RoY9zo8WTLWTGRwUvrTWZevdvaEOsa2nRXQ
zb8ZoWMd7o//biPAXligJ58cSof+QXD/n4wXQRxeD+DaC4UMcfUK1WIxmfNPKMgS
HBu/EGH876JiHN/Z/rdHfiVr3qEF2YNk8fctYMIFgKTElF8yaP7WFzRFmNmNXu/f
GMFO1CMRbJngeDHppksOxCrxDUe/oRs/EcT3au01OK7MBgQGUommw1Yq2C1iIZSE
PjjiL0J0HkunjEZk8CZOwABP1EfKyL3x4r7S5chyeao8uLJB/ZC+osma+/OGzV67
cQlVmR7dEKjopBb9M9IIQ1B09qUpE0Ho3ttTMUYDNCB1C4BlVUnBlYsxJNBkfhLz
lkjvDRNyjnGUvBSgC6C5Ogpg0JGCFk3YcMNEMvtR8Ve5bNgfw6LwVLsgxF5r4+qb
Aoc7tlKMCsG2bk0gD5+5/QuHLUmwAqJzWf7wXxS/Us9DVSNomSLaFosnRZMheoS9
YsRW/IoXu4ltiZr03ENfvcJG+6eL0njGAds3lWsif8u4bCfQkFF/SI1nLoXG/MSW
Hgv/E/glBXMpmrh7qMzm3TDo5cHn5hIysFRR8flTso/9ayj/MpYiMw56997mDLcR
td6xEbx0dldsYEVMWgoKc2PjG1jTpXZeNwuNgd/dUzk6kA0d1lsZuB/+7zfL0JuO
f/3beKUQitx3ckTK0mb00Xrdpxdq2Slbyq4YXgdSHjeWYNm5OayKC03LZryoDpYc
5A5kkga/dXkkS2qnutzJX9pC2zosCHrphtO13GErigo8lx4njRhO5z+fdketU44h
vWbUrptC4nURYgrXsMB6J2FPSFALqRCKvVHGouX8tg6r3cdw7RuR22/J/2l8GQf4
HsAo56EwyX+mC1e+TXqDnka6jOLiN1XQGUvfS6l1GNUCVr/oUCKYcPWzL7pvk2KC
eHlGzSUumGLN8+yL5Ws5/xsuy5Fs701NLdltHDFhxXMpHBktjd6sOOTUsNO/rEnz
dDq0F2zaIsfWdRudxmwZWVhgnnE4qNkUn89BAlbkiYrabq1842KCtLyO39UBCkZK
AJvFeiqxTjzphGiPMIKvQQ0i0o8aDQUPD5RZuEiz4hb4LM1qAdAr/57m2imPb9bb
FVT21D1HofKutTPBDzl9F9TiMVMuwU3/MaXVgn92uu5BMDeYGu5FnIChjD6ZL6T0
dftJckox9c0imn6xTgtyCGYGaiwerEP4EbVPW4cUB9ziiamiiFTjAGJjlgalvy++
uj7b1d1KPSJpVpvgwk5ZI5fv3J/0Mc7rywH5j5UUu+0JjfpmgRjPEawnbiLWswki
Q+IgCmW407+GNQhcVQFoH6r9FlCWxe6+VML0rfS5L0SngX26oXHBvejA237n2VNS
o8RtJrjMFehddC+fMdYnr+SrAdEcIo2+3MTO9Z7lngQ6Caap86TkyShhERPNE2yl
Y0fKNA+sCakI0U1/sSHoOMxdU1JOoe5Pwdjf8iRxcUMfQ0gD87Balegv7wD4r8x3
qsWqwXr7/bA8NLQ0C4gnK9soDDLLQDTcjGv7Yv8vMd9NRnrQ8Psst1xnvu4X1GNW
sLzldCv7KXEsGJDI6a1bomIQpp+qMszH0rYU0QEre3N8kPFDNiz93yaUn+mfTDsh
SOceA4QQ3GzVoTZJebuysNZ8BW+HlyJ9D0265euO+ogBF/h1XMrLPPTnqRPXH4C3
LYUfONwdoREAIf3YEAGO6qK5KV5JGDBM73wyTSL0K370pbc9Wbg7PM77DdRLQVG6
6D/HS+ewnEJbiNcg0DxFEubbQuBrD4J657VT8eunLxChDoDmY1PfHION2vfXhFR2
1AH6yQaIx4Ue9nHY7SmLphr5OMATviv/H2BLCKbViUUl/5GIcc2glKDM3KOIMUjZ
ZUG5pthJKsXRHnmf/aJWiMwnmKPxcXPh2FMg6LHqht4R0qWz2O//OYrmC3ghks6S
LX8VCp3BC5g2s9eN+zDl31V3n6ZEl1yMMGLeSfAmM+pDvFmcgpG6gypa0FmeY8dL
p1219ikJnrD8A/iEOsi5xCxDed8MPIh0IWIK40DGSntANL5DoCdapEZiF937zJT3
0Ss1UMN0r3TEkV38a4/qvQhBug3ma/gXTBhhDFzDa2CZfnF6FTaxA96goi8BLT0f
QS9eJyuBltO2DZZymyqVLRbPFLA/OonxKXaJ8iKnE2e1BU78MNEs+K4z7z2wGi9c
j2kb4Cq8vDSicSphL/7QYdV0UYc8e75K7+/7v+1bKUBDwNpz3LFziK4zeeyR6zH/
J1QkoEuNnZOmuEfjkZyhDAf8Biw6fP5K1kjyNB49wELOnd4wJce3ryWdrSJ9xtRE
TtD+9JiPT/oulgJFk1dRC2DSnsVcFD0uudZjuO27ucc=
`protect END_PROTECTED
