`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tq9x0ebzrN/2RLtK0Wpzckrk2CacAwCU/ogE1kmxhbuefCYaYTakSAqvslwkH27w
T/ahsc/H8jrfeb/OkBJg4UGO2LmTwQ0bEgXLTQqODFCaINQk1sqwbD8km22bNdlX
BARufWajDvktCCgsakanpR/g+r38Srs955jpvxe+lCOH/eYCG6KQTX72VxuGGzI1
OqNO7PhdywNnCTyZuv088kPWL4kNn8VbjBRInUrsmDiq58ZU94xE81eaGPlUOYJE
O2JS6kB4NSFVbTthDs8A7lyBLkCJGEGrVdRtGhPEceYW+MbWTSCVznMJwczp1EOT
L2ag2uQO8uI95jmy3OqvE0c/FELcvSSvPCDq92C+KDYzKRLOQGd88fB5Xx4xkXRc
JY3VGXgUOtog2z8SzbkQtug5mLbPhNY7JtO1fJKLIdU=
`protect END_PROTECTED
