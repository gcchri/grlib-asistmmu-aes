`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjwnQt7GqofB9ITlyPIqEoUGibC2LrXs5nuozoGqYqE7u1zOJ7uvzqiIWhQV3BcK
ifDAsizaTpLcwK3AJQKkq64PShwW3z2KSb1VLiXcvVJyxZc6ONqXr6g91TVAPszL
+1HsUpZ/GZ8baV2dUEl44CnVf9k70eU5t0vMAJtXJXIUyJ+FkfeRgs/V+/D1cumm
XQDXiigHa7Pm8qou6jmTXsLbeVRZdNYe+eizsv9zAgmYbeggkwrkzSKS2G4p8egX
ZnB0abaQHZRrv9QySJeFzIOjPMpsvjxH2Dxz4Z6GXoueaGj7FrVwIVcf5IhMgT0w
gJ4HnS5ADeFQ666xY+WhY27QO1zjxg5hFn5Wdy/Ewqn7lyAfF7GB5FZzgHYQHoM9
cUSUh3ly5TPUfRThsYWJUNU8nMQSDlKARsAXrK3vR1Uy94nVPwS11ppFdvj6ymqt
JbUE7RYC34D7HqiTZyiXbX4IvhnVSUd9TT5VxbQong7w7hIv38xVOLwSsvLZB6Ap
`protect END_PROTECTED
