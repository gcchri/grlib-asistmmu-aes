`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JeuvfBQBISvlIKDLUS85/HA1OKr/tDIErovrputmBRvXEb3VxpsEJCdOVdrJOI4p
6BOsl33Yiql65MqGZe71Wyqkp0y8MzxkKM+GvK6qMRzvBW19CbaerSK0oTrt66c0
8LJ2NfLet2msBfPniFdgsPOeUiKfyKy/QzaQqEdDGQy2phE6vTlv4B6t9NuDFKx4
fYDvnWmmhXzB8P08LWGY4HL9E24rV1S9jqNzBCraHcbsMiSwM11C8Ug7ZdsVfUpR
1lgm6Snz4w+dtE68+z0ZyA==
`protect END_PROTECTED
