`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PhPVZU8zqoBHREz3DQXFLnGghV+GWS3oYZcmkLNbKPG1SEhUmHKNpmXQAHfjpXQV
caCriTrwjIikkGiCEHzXB/3jsYeu/7YJdam3btmYn7ePnaHflUcHzcxJJpe3FFSV
YGms4WzI9nBrQoUtvFuD2dms2FbXfMHEQWk6j68j7NSLnKkHI5kT2iO7jf4chtRv
tDm+1V7oB/n3p5OrR/lSPxH8cT1b8B9j2xnll8LXCbQ27a1KCHurhsnE7jLuE4Wm
HySCSUtAnsV1ejUBVtJvzx3/deVslQgLJh4I5b3U21pwqdcDe1l5lFjfriZ3hB7x
VVfQ84MuhmtFJ9+Y1sKhVsUrSvpaUqC2nZ9PmPoKHaVCeHUpBlCPJ77rSqWIki6P
COwdE+xCk+OWSybJFyGd1qlTggPNkeEuVc75V684u/pC9gtmxWqzU1hTw0uRNcwZ
OUR2jk8wgakw+94ltCjdXRKsMmVfOViWVYhuFeAhujtaBWi16aCFh7Z+NcB+4FBt
ed3Hj/R8oOQmaOB4ExtuKAGyXBuW+piSAas/u9ntuQlVy0FfBlZZ0d0aHY/mXNcw
eq4ByFIZ8CZTHxAkBZ0eehprTOwXRGfeenlGPxmZ+xho4ATJGkJye7UVfP7SQKGp
7/nFQqkm7sDci5fWUk/Qo7E8n4LQGxBZVS9tPEf0Wgcw41PAax5iO85vD9oHpclf
gJo7rHyVVUJQ50Sft9O8M8RE0HJ11o6nbBad3le+qyILWjpN3sLEds/Co2KTOv/w
mCqMqXuWnfDvFi21l3W4gA8StN7jS+h0Qbi5cPpmRRspjfhokceiNqcR6CM8q3IJ
Vy8aYGmIJOqH+4m0ijMnNPPvdW5ChHBEWtQ9eUUJFvtcKmo8CckXcO0XLSQkL7p0
lCt4tqqOx3ObtTA9j+ja8+pecQtsqRNhdgMFJdatXjUYyvpl4yzV1Qvfydwrwtu1
`protect END_PROTECTED
