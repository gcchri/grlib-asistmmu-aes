`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgYrknRYFRreJWPanJnNo+gqnl8HJ34fK3/a8+YUXSKohOTBe9W5tKHpTVKKI0Sx
EvFH6hLuvJnn7DOlp84qSlcTdH6o8wp7IdrXIDFp+JBC+FlAxZz74y3gwQxrlsB/
lV7wQJyyNzFKy6E7Fv9CDyaptqCShfmMtOYfMErrQeAPe/e/1LoNdFwzvFCylAqt
htJa9tbQOd/mI0/icf+s3MmpjrzjfsXnQrlGIlKeTkwXXCkoeDD5/EA8xBwjcxXS
uweZnN/lai9BhAeYD1xScu+Dkt9O2Gre+PJ7J97cIBut8XYoJdAKPes7KNrDrCMX
99BF68TKPOxLe8aTeFRcJw==
`protect END_PROTECTED
