`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tB6TlLhZ0u0xb4Pcejm6taYrnIl16HCZLIFhP9YV4SzO7XPe+yMeGNmiZfV3AM9+
fLvRCYvYmY3lIxxIw1UstZYY821SJtBPH7zJibfSEpe91IfSm8MkJHAx+H0G7Jq+
AjgepBopaINonQGi6VncHm4KJ2ULInQUTvzrVRDMweRxyyrbq02q8hBf39cqcjMi
MN4zaFHvKXT5fMxKyuGqIo/s1HccdxGR+WefNqcHyqtwYzUeFwFAnTI8yokJsDER
CL9qV9ayZgxoC3hOL3nrKQwRDlH7F06hDNF8Y3kWsObW6QEPjVFlVtyPy3rWews8
Lr8NUa+Nybi9LkarQCu9JEiegfWY2AdJsmtTBI4AMyxljiHrmuGLHz05Vm1axfkA
Gddd/wX+uIMZ08qh+9Zf6erYSJid0/xQSxXMTdEPWjmQL0nyREhYHmWOIe9A3k4h
eDCAPeV4CTsMo+yxkr4mrikIMPlXMQ9gXbbRWb3PWeS3afRZjwtJRo0WFppTHqnp
lpyfSZ42NKxju95t55TRjpxvHKhGWOQcJ69TOAYtWMWcdY7nXbs/TZJB8Qiijo48
sVoYzPrfdR3GbtTga/uLFQ==
`protect END_PROTECTED
