`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IgPBAMrv0CfLsPloFxy5JF4PRPjU2LRvXyrdvF1Z3XtNdse8x2cpp3Pjc2pic+l2
WXmNe4PK42FU7eDjPNv5gGchjl8ywCKsqH11rK+uua8/XAOC44Av2XCjmX5HaG6x
ywb/QGRTzv+dGVM81P7ytJbwjJLDzhg9sv1xaQ+z15xfuAsR7I4m51tf+uiPUi1D
Duh0J+w0WVMGo0YhFhRBISWijnknuiL/u3TItHedjic2s00sTX9J2Fhn7aH40HIA
lVfUDQ6CrNSe8zjefuo2JWMjrlXXZZ9l22RHbCIj6w3zLsxmOxtw+Ymp2lQoUFtS
udGe2RMyZDd9HktP6rpS4nhM0eznhBkiYKCoB4oG41aPGfgK8Y7mvehIDJEPAWVG
0WQeP54HjnrClmuS7REd4tWUTElhnJ5NtmzFxy0xSrvYs5GycfjvxtS2yG2q8TNW
ZlODlewkZc9fnWhRZfc0Pd3+Xatq5dx51qGg3G8t3HaMhDX94PkoIGGlf4TGjRTI
76lrpcHixPsuH7tnKOPtI+LovChZ6bSTeIaRj7eQHum3us7j1EaQcOIz5AfdBPv6
7+i4CCRUmPwjQUiawuHu1wsOclU5YEuCrQ7uP3kdN3o0C6/7akyfnpzptZkuyQUe
6BJ9RQ2GU3sCkI56vIcqVgjyW0E0HF399jUtNYiI6775wfkE3jr2gRZa4omQIJZw
i5SoNqXR8voA6PwvckEfYqLugXCDoGUlACyjU98VTV7LcNnkgrvkIdcOc1JXeSkY
TO+PR12u+n8IdLaMUsYXdfMDjTNrjCpV/Udhedk5XRdZlBCwO93FKR+3X+Sssqd8
4J1WpwGjv3bXoV1IdtgRpkM2Nqcxq5noux8L7qHys6GBE6aPWDs9hOwnsvOsz28v
DQFCve5vKzuGuoRGWjP4DFzWxpOfHy3wutBKsiXbtMg5ZCl8KFvbm3/XJIehULIl
J741wPC07wyESRu2/l7rtqyDjpEKNqWx15yCFsXXaF/WXDRJqfMZQvWIskRz6/0T
UiR+yJ9zJbw5amJ4kg7O7g9t3B0O3yPVYky0iLvD32E=
`protect END_PROTECTED
