`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ZfXnDRFXRr4EAhKFCnZddz4tI970qCM13NOWQBJpHzEkHFa32zPVnH/Nt1kuAzI
k9LoPKx/fK+DEBrj9OnYlOicQLVx2+xtkqlq8ueZ1qye0DkjPDQE+37nKJNbkxdg
4zXSViJMEExEL+wf5ZCw4FNRa2VTp3bfDBLrvyC3kxV3iIPoJec+7FNTdXXBMcH4
awXib+H3O+sqYW1/Es0mRjVQ9v868md1Ac2z1q1GXIsXxj4hLtGfsBKklcWrwX33
hbjErAyYi3K+u7yOFghugoRUZrVq4YOLqc8NaoV2M9EZDL/GLZqA73DilWfeCOGG
C50wE5E63KQdrDcIoR7LEj7yJy/CTlg8mekR0JaHPqf9DIOLQCYa3MjO+0uF/TXv
KbGDcom+jvK7wQJU4tItPYgs7GCrLKXALvwTWyQXxDTq0Qu9/ro+JoO4+bTGkCG2
g4BgUTB0ScpPUA6xfeSMtw/xBg+HuTCRhvfMN+90SRxp1k2l1el6FZgxzMhRw3Aw
vG4ClJxSLkbqwx8X9vzxUU3Dln7TC3GSCrm9dquxw4bIeM9afAJofcx2W1KsBclm
XzUrKx9kSaxZyBJf9wn0VAOh3CBZdUgweK+1NQ5TsbO6a0nV3mdRhe0w97xHSWPl
V+Tvt5U70bZ20wX0RdjEb2pIailijLUlHvy8CVA1L0LyEgVXTaefOlkDwKtX4PRL
vGmx24Q4hZOtpJRb1AEsqKq8T9gX2zQL6ZKBMNyGJZC7VNS3qVqoCuvE7DcJWK8/
37c08mEYVBp7yIubEG6HIPbzDXszPEO7TqJJ0+8PHi9bjdDUkgPdGAKUYgUyv78X
RdbluY+d6slC5/nR9fbzMusc73XT90inLAamYsA9Sg5RDsfhP+l08laKlUEwOz7n
KK7B2zOIeT8/gObrl2kbDsi2/ZyxVKJ0f8IgrtzlTOphAbaF6ayu0N8bY0jDej7n
MY2YwCK41t5Po+2yY0oeYRVXm0uMC7eRDl00PgLikXLEXr9mBtPoxH/bsq0MtHJp
COkf1BRkbudOdA2siQZrePUZiFB8eJ+pPv+HCRmoBaWtN/zfefk0luBCDW1lp1O/
o7T26oaIR2fnJRXGWucHODNLWy3DyEcSBEzUdvEJGMdgNb/jZnnhLzQAos73jHCT
bzEQU7HXwt5XoJMRiOHSmBgEb+qzb4U6snVU3G8f354=
`protect END_PROTECTED
