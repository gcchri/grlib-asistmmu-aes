`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ADS9IBLFYxoOL6fuO+H+a2SoCUEcLwpNmJZOUDH4rv2SWny9i0M+FuwOaqCuzzjW
OMtBbO0WwhFZIC5BU5zQXfgOreTHVIaC6MdsxK2S11qtkxj/gHIoTgxnCg7dic69
0Haqim4oKJQFEPDMr3bgWWKwZ5Gr82qEVB/L51pHLuKVbQ6KUBZ0Sg43UcOEYpLc
VppPJexvkp34KpRa5jPRGutl9ZhDyc4b+u5SHDeRIkRPH+Y0uQv0OTGux+DLjGbU
IJMR4unI/jWNduusjadJxbUZIlS1DAiT6B4go9TEAzqP68GbAYuZ2/I3BIkZSsRE
gsDlzcvV+jALo5JnhSfwOYL4JMtxKIZh+k25i4bA4LSE/C8xssJazL/CC3VTT7Qn
PsKTw89CAiKDuf8LgF1a9kYhzPRWxXC9tL5hldUV86nnxEsiAUrA1HuVQcYRsPGQ
4F+yJEtsyrrkhCmY1hm2lID98l/CleFPHkxXsAD9/ze70vRvHwdxfShJAOt8dU70
16z4XUOyyUG+tCmG/FS890hDD8YyCHrTDLSfrXLbFmRpLbzX4CV8YDz5uZaXUKLH
B/+qKle0b1o/41kSTEWeda3zwc1Wbby8A5OOSZuL10tcZIUNfYKrftL7IjYWEMtI
wcqEOZFCV+0aAg7ymp1J5d3ffP0PqCs61i37A6pJnYY7K2Sxl4miWaNObiIPC5XH
bOBOi5WOJwQqNZTyq1uRrhDbjGNCxo30r/LB3IV78SsEEDo5/1k5PPZYMF9FcVL4
4KLYnE5+peBCulgqxnc9mBweGcGr8nN62Yz2C/W9eRVqrQSERNmh4GYEZke9ehN1
Oj40he8qh/OAGGryJ0+rQ5yfK9belGdxpCckNPS0Jui9a6qBfw3zbb91SeMS3Vhf
fUxrcIyIr7hnOvdu/jXGeUJp5/VrkM8ztJrCduo8oaTCHeCXsE9yRg2q83P57x3s
vcDDg79wSTiTtqdbCG0A93c9pFFCLarcD3nqZ3PEyDmxVxx9HDmsL2lOAtceSmGl
8JAHFL0GyU04nVEJB5K+9l9N3hNhSFYH0hIC2w2blnwuSRL3hD9PVHHbVCJ6ovDL
5qN/KyHDRKcxWghA7Eyg06Hqguek636Y/NGX3S3OYoAz9r5bDGuOYHKF85s+vqce
oRTvkkmg3+VmZn1459jfGjNqQ602esTs/P0U4c/q6i4=
`protect END_PROTECTED
