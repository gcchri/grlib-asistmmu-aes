`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/z8p+/rZvQopgrK6rkrbIzRTSrrlZnOlZQDtFUFAnDd7F8dC4F+Wt2uwCLKWksrz
mIkegSrLug9/ix5VI5NdrXCw3UKXwwto1GQ/BwNqZsf2kw3TFVZHs3PRKB660W9X
+K0Rr4jkhiU0Vs4B2ckX//yVtRW5zBr44jmFJvyKmVZ79pCig27mq/MORykbVLG+
/hoEUeZlY5Vu9JbSqwjoQoEQJ9Lxxga05FiLcEvfx+Jm5z1zSn997l18z3T2CSgx
K2ckjV1EmyvkhOaxCeVeJakdq32znbNVIaHC73YR4wyCUW4khFuFPdJU3XiMlBoJ
nfFEHnZgsTNkatavOrir4XL9tUShazoL4mVERU3eFLHZtNExIEZUgpZTPq7lgzTP
VrNb6uauRGUFxZaG+PCO7DOpctA8a3K+Vgh4SIITT0Fwnlkd4p5/RPPFvas9cRMK
cN5uIlFSCCKfhRzmPiJaQeiaT/u/X0AinaL9HJ6whAxWtodk4jHuBPBRpAF/dxsf
0CkhEvS6Df5Wpau564QeR2VWLRst51+yFUR3rQBY8Lc0q50YOcEiqh78BUhQiloj
bnn7PjRRA197fR/JSAl8HiA1uPoJ3/B0yNMc8C4cPI9KziTgzUmPgCwaKXBgeURj
1M67HhYoypJKl3PoayXtK6e/T9XqQc2ZYJYArCJOI10=
`protect END_PROTECTED
