`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5iVAHgejeAH9H+Nnd+gALgBxx+oojM8UB5e0lh7EDdYqqW/kREf+QEkvVhqi3Axy
q3s4Fw5DI73d2SOkS6v4IIgozjFprzNqTEUd6E6D/hWzc+fGTLqXgfLFFdiXM6Ay
rWhnQH0+LK9Dwk4aVjxKK5fZm6jTbsqVYbr1PSvZUA8Yj6ymY6Y6Vgkd2KsYV9o0
go5QSSE9eM8NugmYnIUOgk9gny+WuD9kGDOLEwV22l/m0BPrgc4PefkxvWW3GwTM
R6KQ6xJhT1YqK+vlmoHKeQInDhTCoI62uSdEdazdhlCfrVGWtXVlDc47YylxDAfB
m3abPM/lhU2IoDyGD/fqKYtOZKU9CUyqI1xyAn7I2g5bV/XLIDBZ0/kwS18e77Qf
4ur6v2ZAIr9caxL2/ygOCx7Jn+9HvetPX9tnDmaN9kr25/vGfAnfs33bHMTJbeGx
m6GJJIrPOhskX6+746eLDbWUrJniGaq18YcU5IdJFylTjwMO+dGgKE51PsTkDOlE
0Qe5issK/T29KoZxJ9yAMVleshEioPy1o9AYB5kD9RY=
`protect END_PROTECTED
