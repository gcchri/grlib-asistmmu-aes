`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/imJDb9d3QMeQxF44d9r1J4GSyZG6iHmw/NIqC8tQhYiXtaaBCh8Atm1jJ70pioS
K8eKiBodARkPC9mo4/xJ4dqgszANaQISqnahrTfccGw++wQO3kat3u+janc3dwzA
PI86aMDU1MaaZBHHYLL8QwGP1rpN48/KQ/LF6R4cAlLgucT3JJ6rXk1py3CV70FE
DTajBNrV1c2FyG4Hm1BK/yFA2gqIEBwY3ZUP/cDZqATbptKj1PGeiU7o0sE97V9F
TtpNR7l4wLANQ/a0f5p4Ig7VH0CT9e65rUrD8sk5I9rv2PXs/K7gn1M5MfUYGLOS
WsSPJPXUFayMI1mcRPMKiVP/+WJHFRomGOqQiXwI1NGnWlkjqsxhFFYy7BEBWcGF
FMUyizTzmdpNZ1vfaXXHTWCY06QnzmfjcHxBoW+31KW4CfZuwvNNRA+ACxo63HdY
`protect END_PROTECTED
