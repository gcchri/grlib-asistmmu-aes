`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lBbl+PhNGLJFbTef5pjXT7CrUwpufCa9sZect8G4CThNW5BcHT9fEUug6vLh/1+e
nsxnA77BsMI4Bj3hR6NvxhuqhhJtgreTVC5s3NY7HhjEbHQOb2MnHAFkVl/Gd2mY
jRQ2l7lxW4x0BH9mZ2wa5ce/U4KYOpwxs98ReATmYenQkSDnXCulTTDtaYfYc3ey
USpfPpmaHxCgrDF6LcastJa5KHHMdRNpG4GuI4TCBwi4hmrf9u8cEHc2cPH7nuEF
YanPeqt1h++LDingbq6RkOeIvvhPqQsXKY5H5n68Hq15R1eC89hBKuyt9joqLkFf
S08KZOSjVEIxmMsFYFPywbW/4NSRwMzlPi6N40fo/uB5nh6DSpcQqLoJLC3bKHxs
7BGC6O8YwC9i73oKhizd+e/yYCmcuOttUZ+XiwEn8CBaBkRjWnPoxR7yU9dD4Bpj
FlrBcfnNkjshDdYVhT9i3jRUu+2cV1zXqeZZBED8oeM1lskwzUP+WIrtulaGx3HD
FTjpOYkyrTBfkC5JPBWJK9oH1a2mlKmmub/gEdNK1DcpOIMfNqBll0kh85wnZUzb
jelHRqFQO24d/QUTObPr4uoJbhXzmNrEB06jZz6n8D1r+WQgHH7VoWonSGgmDSUj
yZhzoHKIExYEpy9sGUyCDcpPB+poYoF455919SmjZmRQBKt4bkq+Cguuo8jZhur4
gP3SMJ1T/97a2hT8FThWXdQJrlwu/QyADq6CMYuztUI4/QjWQQysZzJfs9SC3LQJ
n2UyM6PWSVqpP6oVFnVrhZ3KZISPjglMPTAaBUm4YBb9K5Pi+rzm7JUqjs6O7AAK
y02fOu+ZwPoidg/dLKLIsbsnJ9lV95Pemv69wif9zIO787sTi6QKQaKXChxvZ1nW
VOUf68WmJQjH15bD4pteBKanZO5AcZckALGYFP+VGBsQBLno5+F1Mjf26O3Idj/8
yReJGQW8Bz85UvV3EHPyYLMDnaNroLeDPe8NkriOwn6/1NLAJJE1qD1bO5/O4ECr
v5L2beuo/EMRBsPOXtylP7VTY7YjU6IUAUmoAoSBZz6leAlInnwW29GbKrtAs19A
OJYeXb6SroHxHfE6/D+z3u4KJtPPSX8pskuLxYp0blPGWTDY1XnT2oWlL1Bm8595
/M+qQGo43tYiiAnQDUnmpuV8115O1CPBjGaIFwIGGvahtdO6A9zkqqBjBI+FFRYK
ArHoIAwv6ss5sX6S79kswK8TS6apWhYcxS3ZqApzToHpq4TZu40QfzueDKNXw/KY
CcSN/WqoaFhJQHYSjg3hGLq7xgLmVgRa6aCk9v9z1GqbRXjXVaziO4xayBjkmGDZ
Q220FKpkO0jyEyye4WqLzFlGPSu2POHekRf0R2luZbS6xY3cfMIAiKRyOEHQXcCm
O89I3RAdi+FYRsvy8wE6WAT4jWNwxLMfN3gqgkPO36rmPVkGo32Si8sLnPIe1G0n
oXEbEp1wMQqM047QZscA5sNZsVXwykn2ayVBpBmVIzBexbbu3fLPPb9IEOojkbUM
f8d30eRObGZWXUWyqPuGL1LiEM7ZMCusAFdMKOQlW5Um4cr5GAjLaBtXYmhPKAhj
dm8tRJI8RfXn5YK/Fn9aof+PGsS5Tbn4ljfgSaNE6CojGFj1vYNLQdkjfG7Qv8Va
Zf33QisB46RsUx9vWhJ+tA==
`protect END_PROTECTED
