`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMKyRPskQHH0+Ho/w1WG4XQAM+6aCirLK550dTIMcvVm6/uzYdzAoHAmwRBpqsHB
D7fYEAPv2jV1/LUjxkb0uUrZtcAkME2XWknQh/DiwDs9S/k03dyjdnFURkcAaInn
qISQdfsoAs49B4o30kzAzskCsyw99Sd5GCh89r35B8MQwC9CMAS2ZzFvOzcoOAR8
l9ZOloQ573ps/J0cYUEcs8gRp4MyygtuCSK2x6LpaOggHmskRYPhhc4FGEUHZOXb
HAWg/ydTzT1E4IlAJbKuwPKkZQvfJZCWj2ycOFR86I+eIg5CT6J/RRYyDEtm846f
egoQeQq/plzqlkQUVqtAwQJNluz1sZkPsk4QqxgHwE2v7bO9xxj25IG0w5g6tg5R
qd1CsD6T4zOVB6UKQQpSFC1z4O9woZ3ct4vezs9PZHqyOpv8B556NTUDW4o6dIfm
H0fAzYQWba69CO8hBjiHzxpPBFrPLU+qZFA2FnFcYkBl7h6BdKSC2eSVRxpJztun
fv4WbYTSJMeHWOnP9QBkQXBcywTQwnL8sa5JJURiO0sYgmwCJe6u0P+jldidmg5j
72OZj2BCOb0O+wKrWwQKDrC/PvXTTVHVImRN01O+cvyYBGX6GoqgXotCXhZeVQVA
cb52DByb/JpBrbXLR1PlCIRF1C26Z6FqZfAu6o0+9BhXPQITxFOgE7VScIBslMxP
fmyCXbYcijgRzcAIFlHacg==
`protect END_PROTECTED
