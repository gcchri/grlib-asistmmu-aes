`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSd/uVswMArmfNBhTIW7J5TCiAuzeBeGVCyLDxxEmDYK81q3Rh9P/6l/ofpO5OrZ
83BeyivmJDmSeZWBXZ1Lce2jMywaE2X/phbfulWgkpxci054Y88Iz1w+EamfWwGv
ynFtReySfQfQy47yJi1GjEihsPb+GiBePdy1yeDs56+JIk42v5lS71t+CwDr3lwh
x7Qeptu0XkYqMgTsQQqROUpQW4hWuni+fbahiyseb8lqmOGixlmJ2tTI/z2dlTxa
5Oos/s43oSqjE/7TwjYB9rJ1Fd6W9ItF8fScCuh8L6GhnkkIujjnMIJYTUL9dhrO
p3AvaN7WR9sSp40zfdG82xfptsXq7Tn/KNvH9pHVZT181PMTAP7tjCTEIPpJuG7P
tNtoi1zlk6jevE41c3jUawM9zLvPEzlnIcMq1Z9LfO9zm5DQW1iGDXZEWa3bdR9N
VktleXp70FzCbKs7jwnZqv4613T7ebiR9wmb0CIZ3YLS7BcV0S+g7VsnmRAo3Xpe
IaGXWZqqTNAhUOzipXJC/ypfw44Mm8Q4+mswaIKlDnmWI3CkneGwTZNZzU6qcS7J
9vE972/qLoH8xf2+d23wmUU+YUq/dL97IbmHUX3WPAT1UUCxJrbTq+FjiP94R6N2
wqo/RO8mTh9/ZRqPPq3z67BgI7+O+L+nNXOP4fOxlRYMrDEWwC1kIcEj/xi789/C
W4lUuIuu+VwPRX9D1Du9tblsWyXnpEvqiXsPPCvM5zMgQaU5vqlPqxt4ypB17HVq
UAqLQ7iUuTshFUv+Txp3F845CQRpYiR489svPHiG7xK9xBmPC3iS8loF/0NV3GMQ
vyfSzXej9XLi2Ldv4fK9Hr8J0Thv0/yOuk3e96z9mS+cfXTkauJaDcnfJ5WCnMXr
m+LgWdpwWWWkZ4wZpwaBTH4NS2QkaHFhp3TNsH7U21M+YrgKDD/tWKhevKCO8Lws
/dbd3DIW4S49yXZjYw1Tqx/ZC7rr1fs+FiQ054sQZchmDQXB5e3tCGcloo/1R7ZH
R6dhcGcQiW5QvYJK2MecK6cBG2aOHZ5gsIpFGIfooV83ou9M7POZDYn1NLGDa4NW
g6NDPh+wBu5nHz2F3XzFuhYi2uP3oqCPcSt6UU+IgbOIf6OPLDAxIlyG73idFefz
UV2iGJsBNwz3Nu8Abc0OwuAlWS0QLa4ERhZvMrG6Qfi9zmiHlUZ5bp2durdvDPU4
mwG5jEGC3XlattWqbpUCw9tSpBreMamVMTiOXCMHbx2ZGVKBr/+2grxRk6gKXpmt
wmq9u6FnBJVP0vErYEm5Bxk9ZUM/YYHY9v81xViTrohoUGwMoEEvwQhXumSTuW5G
7SCyJlDi0JLsbhtSJSROTIQRPUjyWjgzpZwu4FGmu2t0uxGmYNt0nn3GdekdQvvM
TmXh0JQ4Nj2r8zjozyoWi2Fttf61Or6JBEHmnT5hSOl3ctYOIRzMGCGSP1T79+fs
ztcgh5eqCC+bH3QMwq1Ci/osrtW9bbFwjBX/C0Oy/0u7ieoNKB/36LGoOFKPo1x8
RqssVpR1/8D1ODYonhTlBj0mIAQIopTANHa/RiCEWAi6L0BJwvcIq3L7DEZw2DSs
6a3Tc880RDq2BJ+YxmKnhqJbZB/ldRETXwyzXuSOZ9zonCVgaM/duMgPPb6tlGmR
MuhszR+1TovvQtDWs2piOays3MFa/J6BqWgRLL7lXiGsUlK9k2WU++NUJpQC3H8J
5CrvbRJyZHflJe2tVzznlrDwXm7BZQoVz/keviRp0EhqbavJRFf1jdMo695O1NRg
f3qoe+X6f0lYINX2VHZgti71Qnl3try96i6pg+cgLgwB0sgwXV48YEjZ+q4b/L+B
SNhbaDWJP7Lmmwc/Omfn1hsH8jZy5rSshkQHq8c/xfrxrLY9H6TeWuO8T8tl3zkk
mj10SsU6fpsSOZeBgsbHSeXFyQlU/UboO36HnuEBYLKyZRBn5PdQw/sboVZH/e7x
b0XKyzf0iFYuuH9AJObX6L7jJbvd0oal2Lg50yuDGLV6Xqo5dGA142GGLtcFkKQB
aRiDRxi9iSDjOrAo9+aX4Z5WusKBYLxw1Z+ECHI2Wy2FlIBy/eyUxXOvalUxfXCz
mhxffIxWAPMccOJW2giNISPX4hxjPsBtRnrd4VBFspdnMMf+AbW9TQcu3lciGUI2
`protect END_PROTECTED
