`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rpvYPcX6+kspBWIGXLuZ7PJ/gPQkRcw550y79+BB2eWQxbcbhF2OZRn9+LziS8BT
bqvX7sn77pwUyJfkaAdPRDFdMK0AtEz51njPXENxDaUzFID7iGhVWmgLVYOZwdhr
Z9arwfEZZAgTqOzWV5WiyzyoXUulKacRoebyx8KVZL9zo1p2g2Ecuoz5WmiD5ACl
EAAAIB/Gwu6eQTNTDBqg/JZPJJli1DZSbYUTAmk8YJDbRhyuxusIkqlUFgmVtyhT
uhpEXDADz2Qc2Jojb1RSo0yiNIlexqmZ5zsvAiL4YdgQyu2BQL4kz1vzckpzB377
DPgDKUzWsPdS2LLe4/Ztn/QrCJOz1a7JiYXq026kupvQx3B1L0j4ovJ8S99pyrRC
`protect END_PROTECTED
