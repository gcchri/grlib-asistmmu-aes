`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCdkK0G74Hyq/4EkPpH0zOtn/s+vF3rfshAHs36HGNS7o4N+aP2diM6NZbJJ9kQY
HKZKCVQqJS+IfpnvxmK+KWPIGlHT2WYXbNSedCJQmyl+KIyxvo3mABwgfszLTXf1
pxmWa14Jr/tvLDCKHGfKWKzlQDbUu5sNZx3QffLF7juGKEzAnLU2Xjg8jhLhSVdJ
a/m2rj5GN9ma/WOvQPTDXAec/urm7WwGz5B6fX6KHsreWqX2kEaBTXU2LuqvWnb0
v0avo8Fij8yV+4oEC1IOWCISHWcynpt3z4w2T1J06WFdRQjnN4s4MRSaZ+ZcaEOQ
v0GBIC5hIhr1/I5RBDGKkU1vJm2a+vse0a/ix89iv9ReA6KihMRUiauA+20PYhx+
U/6R3Sjju+8jyKqHPDT2DwnRbANUYV1CcK7C//UKfq8=
`protect END_PROTECTED
