`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7OrzSjb3IqkDkjtjqqgqMpQgIdDlQahvqCp6ibIATdUw+dmKOtL7MIMdveotvwV
TtjUp4L83LrhN0sZxQSp/7F20cp9/3frqGu0D4kYQSHilE5yJvzosscZaChjqV7r
G11Vs6IOQZ8qtI3mSXUsIqQ9NisEtq8KQ4hFBWgMHQlWuPm645X0xcBtmzPfQ0jW
YFvYNi9fFSm/S/Snr64A+fGgFsPuwtvzmS9GW3OfEmugUqesGcW/NtIrHXOyM94k
U7jkmmeQaEjUhnE3oP8adzhMroz6Xo/CyddWQ+VbP9i3xKexam3mOPVRizmI9GhV
hO0tU3p0DLVVeZPuHAvY/g==
`protect END_PROTECTED
