`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETuC+mBSQUFACgKhvcSu8PwrzJOC7db5oVPF+vQ/RkScRMfPm9tbNNUoaWqOZ+rD
/w21ZkHryr25k+dzpndP8YOl9wub0RTeORHWLwKcQa83RYMnTev3bjbULY4ATd04
4dsFLDwFu8r+e1eXd3QAdaYqkyttWpWmCUmisA4hba/5XTMZ05CYibAXWUEZR5lS
LpD2Xp56VpfmwWDqpKNZSU9v2nx+U0o1zVH9ZIpg31fD60476RSgfoyJ8Dxyx+hA
LuL4sxL7PNjOpI/nXaQ9tjK7QOFx0o7rYBACMSGcpPtyxo/UKIKLPlTUH6jsFZmj
ChxU1ROpzD3kyQjNKYmgAcax3/iXkMbOYo2UJ7bLldOU3VWcL72dfuOGlFWbNWOm
zyDausDlA878Fga/TNt+O43LLJte8h4g85nCCjlK6oDFiupeCxagei2ZH6litzLi
`protect END_PROTECTED
