`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8qoPbnR6qFk1R+G+o/e0CVnjmPrPkvpljuSyxrkXk7mX8ts/azK1aC4R7ZIjM2H
qIQICgiOofxwoMp6M28SAs4/a8XDQ/wOTw22dUL7zjXVZ+S28C68mgkld5tGobDw
8SkgKPZSvsu+7yEfSNpUCMpliNUj5UrhWIaDu/JGyexEm25JOfIFEgzfkhspRGkR
B/Y3rj1zXrxIBgJSvQusVMsAIz32RP2pNsO7XJ9OAMTuKfMww3+y42dLOahk+Uik
0pH4fyc+3aUFDcrgqL6ODvwaR0GmjD6ewaWtxYB4JE6HYsnh3wnA6h/Wh/fcsQ6/
u/10HldKaHcgwt8r6LJJlMJfSJEeNkT8suvcOIS92EWkUvr04TeiyvkEGJpeKTDg
3i0TUCSZP7BcWzBm/7wBA4fBpeRbECl3DuTQW3KBd5/pSYXS7LC/ffG3J/MoR0qp
Sy8cniO5ogJEfYpvvm0knKT0SL5Ry/fp4EFP0L6r11ManZzSs+kiAgm4OD8webfo
rbM3ZL1amT7pUglG+QPg+H8LtDCqtB6tFQKeuZSBQRNXgdHCY926blLA/P2vszFe
T25tZk9t8sY319gdpLdQktDr6t5se3IDKFujsv12TiEH98vcVhOl9CrOc1chO4X1
MRqyzm9XxZwAChTMCCHkX6jo3HPkDTKbtrCZkZnrF3qz5bLLSBKd8xwmOq++y0TX
5+I3WnnThL//Ddd0Sb+LVFdKETUbeSMZw9q/z/65ddBvXE1qFjSqcsK+dSLnGr4x
7psGqPhy8xc3UjKp+ab4mm6oe0t/gf18F701WHlAP+z+DUKtuKuyqE9LQ64V4ieG
rKImdbtwjepvolcxq9FPEp3hR+Q1tj25oXJVF7vq5q0uJBEqMQ5Ab1SOGF7J5OIi
h8o4Vssw3eG5YAZxa7sQngd6CA/v1kIeH/2feqPEJsKMM1zrPxZdMTRAv5RWS9Y7
`protect END_PROTECTED
