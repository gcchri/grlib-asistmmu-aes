`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ouG9vOtMlZIxQekpq0m9UahnLj5+LjZsrxLWmyqq0WBF5gLhajMzVmVwldXvIzTy
lYLkx3ywEaTYHfIOPHAxGuc0OZLmMdtOk5fNnwnKZMaVreYAQGiWOFCMFyGjqHPr
/gMKKpFSYI7uWxmkQhqJLsXP9xrB6B1GJoNz6jXs8IXONOu5gwVq1vkKD7yMjJur
zTCt6zGPBqSihCz3hdgC3dIf0Eta6r9RVqcXnrC9nWcf8X/ejnt11lwOjoaNJOyd
FxdLCJh2UKW/R0xFgCEcKAI7oH08eWWOu01V20/txhLGYUWt6xJ/z6YaBRjtoB+R
RLgZuIS/HmRyWhRbm4v8iw==
`protect END_PROTECTED
