`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvYLt0lou/6sIGcth0TyUw9NzCo9fcliGFYavmHntxkWB92IZuN4i00u3sCUn9Xb
jJgq4LUP7gkMWowagphFBCwUdIKuuWKyBBEpjOZ7ukA0GduVPzZNKXX8Mxsp3kJI
YXHSpf317dxUlFg2mLQy2QSEGtqMIHemUiHlyVsnN+EVAKbzFL6XuwVrRKfTQARK
OzD+1vOFrAgUAiKDE1Qp5S41tNX4HzQhp+UdumacA0nh0oz7IEliBQBwAK0uXcIP
hn7+clIsntmeHL9IEl50vN2BlI8iDCr+/bBbiIEnlJcsptLxqzp8yVND0dFlmDDW
vdsU8jHSeUZiKcstFwhAXlRa8uNWlKDNiMdUv1wp5vnVJo+F05A54ld8HWT485Si
wyhVgckaI8ka719znygSvkUHDK5ppiNbw3iD0NkHR5k34T0ZOhjfbPVH5emZE5J0
N3hr7yHulFi6Y1buwhdPlDTC4Jyj33dtajUFQBWFwNg=
`protect END_PROTECTED
