`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sAPe1Q3kbevEb82Na/4HBpbUkaR5A0k2y1W+7BYKo7YsJcx9vOSdS6wq3hC9ksIZ
QI0qI3zVS8oxQurCfSDOPRJIzSghwaD2s3TQ+n0Lv4NBUTusOfRD8ovY6Nfc51XU
7wRuqnlhHov3WuTamis4qAWP3D84UoygnFF78lOEwVywKIonKnG1WnbpX4TvzfFN
CRzxxnRupCMq0NEIWhc1BpBGNdtaTCfst96QCreEHkwjLZoIoffyJlbm66NUsX+k
Nqjr2MlyOduaysM4JLTip/UA6dGL84XlCuaCaFqZnpCNOt1nNusOu2QzBDNkD3JA
3UjuZLxey4ERb+TNTjRnjOsoWW5rcV6A3cCgiuOSq4aHhdeuu6sNYJgWpun1qFMe
F9Y9Ppouq7Qd4aVH5jzgQt3LYGLAT4zpckoXTG7pNg+88dborODbGoJwZfc4MWfS
+iZ3sz+1ZNgd+PUAWUuuvDpRIJdQOucCyO2St5Pw+30vrVx2ERfD/rgcJnbvQDPT
`protect END_PROTECTED
