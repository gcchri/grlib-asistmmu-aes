`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mi5OcT1bg7fWagoaoMWR+/XHHn+HMDzlMbl/90Rgsz8NhAHkA3/cnzBf+k/j4V8Y
ieWP3+cQev5MGROoyAAN/zYHkWe/Ry2f6l34XNhKq5TsywR9hNRhgN1kKm3rWzfR
PjSJ9vJfqJH/PiLX6744oZvg//qkToP3Mr3KIzKqANLGLXgq+OH/dukqZW07yVPp
/9vaa3X2c1J12+dGQJzIlZrhqSIRmCW4T00XgRkRVj9UaTyM1KcjTIAKR1gqLmer
YguBkcT70zwFH1ZUucG4bXhKw8fPonMclLaNqHxPdWQgHhmVxEbG/dWW0Yq6abOI
cCQagnTwByFHyCGrjunWAjRrLCuqvgNQObGvK4r7pelz27SPiZb3MMbT5saF5ktD
V84loskaiNILgxgzMNRco+jee8TAcjrVUhSqxBq6Y4tyF+IUaDV7coIiF9FtpECu
dfaDyiepglyyQaYrEwqd0Dkv0S3B2NG3zGbVZ8hnhW/56dIA3NQQlbeHg21T3jr2
sIXjKl8GHC0miW1Tj8icOdONBoe1QzdERVhVG229sN0FoMX+SarHupKn5S8c52ET
Ps5zzJUQnlbSNwFR4T2bi7oE3I+v2pi9APLOUpvXNjBKKJvqWWIN4gXEBOqKur8Z
mWv2pYlK7S3dyEwYcj++kg==
`protect END_PROTECTED
