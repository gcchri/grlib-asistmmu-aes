`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXCD7mMwEI1L/l0o5kNIKZQBJr/5gUSVqH08yv6OHKrZTMVaFqQoxrgcVW+J7K7/
yg1WLM+msmZ7IjdFlSVbwWM9khLM1S4wK97HBSVYVtu2csMJUoJ6/qNIuroR5NQU
7hYeCFN/5bQYGsEkWFfuVmAv8eKEEP8Y1u+pIKVgzeWcTGka0QTofYxPipkniBFY
JjV09BVktr3CRSra2AVNddz6rxOuZwY3paRJb29uL6v7q8RHNCAA0pqpifvpiJIE
2O9EPlBszU0LQSxKMfS9wrEpeAph44Dvjh1NF9mRipcWbggNdFN2+OlTBu5QFagB
O0pSBcavyxkjgIBbhuvMJuYps6w9UozNq11T0/vuhL23xfrsk9yuEk7jY5HSk6Uc
zib6WH5hshJqvYx4Zn/X4KOMeeAJ08xZm8ownEatnzljEEotTtvFeBOoNrL4e3TO
kLYOt2/I7YD5BhQ1+pZ7jkaLs5/krlAjWru41s9Kjz+iI8XYFAHJJVTfx753i/M5
Q7Bi02e8xaBPW0n7/JJbHm5GxMRjah6NcgtzkZ0VFjCCvr2MGXD8umbIOlZPfIjP
H28745RZn8T/YVrNlsjShQV0V4K11nBNfMmfW7jfibyASXZmCCSJhIOcHPQ1Mr3r
0r4ax3TKF7SUSitGnsH6BkswTVGKGwZmdOSSpZ78QxIyB7jitfi86mkWUwdnUPi8
4sALyYKJGgOD1Ao9TkRVkf4mLK6N4ygYO4WakzaNVNo4aRN1I/XJgNedkCsC7cIa
e1gb3yi8PsLywyJ6OkBBe9it77M76xtCvH4rup92Gv1zm/Lh8quuKwaue+7rBGBq
QJDmVPdVI1cyhr2wWIrHWRcdKNCaQF8hoUtPrDfDKm1queJFQDdyAO+YUry4tSlb
NuliQxwGbe7tUL25FVVzYLyy8wnyfNON3NC9ij+lxDleAi2Ph8PJ1/3CBkUS9Vo0
6Wjwk8lEpOg2qw1cv8NY27yWLJ5xv9Nm9EbpI3kEW/PhevPlPZQmrMjfl2pW8tZP
6EwezHRke2o4xTU9Qf5F7WxBm1JKX7+WavCnn2oj+jYBUqOJPbj2MMpS41UbXx32
258dkhqC7SEFi/vmUTL2GgXPgSegeFX6ppAgMQJ/QI9ljzL2taFuYepxdp4poRIz
9GC7oDpQbfNoi1+ipRieOFg/83doo5hZSaBcFxV9GYtsbaVvPW65nzWRnc6G7bSk
ZPDmi6/1FfZHVaERlah0FqFbapVky5iWYDxRYE51mNv9NCNoWm1L1ewl1tP2Q0qJ
7y7+gAGgoKrdItQvCDIXAxEyuWFQtw0up0anznJAqY19H2pwYRmdyMQUXUBFvnpe
0gDcQ29IFl5jvAmvESsEZdLjQIxKmqIUoJJaIi+7/vSYHLkJP+U0Qj5pYXvYmvJu
r+9og98FPMIhGUr+lcNElP5SNsnBA8bfwy+gqc1cNIiLTOleGd7XCGlMftYQ5Yjh
nC807vAQuVqgC5ejYHUrEBdqg0QB/8mRhh0WtO/kGZjYl5+ImSgDnbsV9dDW7e7I
vUiE+jZ6Jha34LYYQVx1PLdeawbrNWoc3I1+Rl0Cb2w2V9wgf0DTPcf7K+/N7KQu
CqzemoDq6X7HCNrkELDlFNTWVDL1kq/BOzqhWESY9nDYFP6U8Qc4VaGz0K4OFxgn
KVDafXsGhtcYLrcPRhIKUKtixzbabT/fKPx8GdC6U9w=
`protect END_PROTECTED
