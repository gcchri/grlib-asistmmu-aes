`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHp9PM5kbgCv/wWgnfrRkHiUjkt3hvQv8WIEtxK4ZS9OPRvlDf6+dYnm3JjNzGx7
HmzXjXD8D4nJYEnJSjVlZc8PV33KonGqiVK3Np2VRxWYzSjFLWjQrYR455MoFIrT
Sk9Os6WA0h1ZUsSangmHagBpM7YVmXQwof2kn6La5yzoVfDCWuPP/MFRlOi9E2Ig
q2zeKL6lLY9Va7Bt8kYH4tmGievIzty4ZzJOXT/8DFplNDDuBspjTVfeKqeMnE+B
TzT5StYFEFCjA5y7SDmugNkb29zyFPJgnTxppmVoRs2eC8/EmVa29eavDPxn+Tr4
rjuctndIGVjA0BpNXFgfOcJlL+PeEXshLYUn7BlFifKCE8nUWUGD7X+KyYnsO7+y
iS/BE3ELTNNLwfhILXNW2UOdvCYuzidTDpxEdYn0H3jr5fpxdqiFW5XEHnDatAUB
AimAIoLiyFY6uupXqL5T5Rhgas7TbsUqqWHl/vyMU70uZnCJl31sirElSvA+Avv1
`protect END_PROTECTED
