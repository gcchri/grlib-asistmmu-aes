`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txQfeSipjnpIXmUJ9MV0phVQDcmaTJmrRoYHAzs4NGGiZk1N8p2YPBC+nKqgT1Uq
WBaFzR8QPK7a3JPY+Hhgof4nO43UQGc92EN+nWxFnD//usqmdHBMDdP1c3ZKnavV
gKo6eIDfHDpOToGNgvCiTNClZ06hXa9+T7OJmh8QP9oSFb5OaGdsAb1cP+hvYNIJ
sq9O7zvvQnpzyEA+DNQgQRnsQlbtE2nfv5JGV+E1YfIx8v/vBXYiL7B9LrC19/Fo
KUbqi1TqPJNV8FbeXZuNRozAXDdDP7aNVxmpkrNpICoAPSf+YtonwwQT4OnN2Fnd
TT/dVdUCiVXKBaBjhdE7ImXGVc2lzRqS5RlRLntjywDJconUh5ckmkNt7hG9ZV5B
`protect END_PROTECTED
