`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RadepYbYFA12ELci6eM5L/y59qXL7tGoUHNbQHqqo36ejhUeGyVHbcdsX8vHBdS5
VmUC65qtFjFxD2SBMQG/sE6ezMNzIE45I/98RyfMm64nPAGtpVmefmUVagcFsoHN
0hXSBgt10KTVVhb0kI0God2HIZ3ekPtAXO+xEbVwn8nsFpybtPzo0k53PCy4TToS
ZlFKxNfbKZZilhE/mOwMTTR4U6kBp44kG3iLArEpCuSibcy1bMVMnC7QrgeeAdgV
HjfAosV9zfWwHv+QFSSk5LixBg60sip9lf1j0ujQ8YfB582BD8dIbR/S2FcnoTrD
IezzKtJ8pYQsAMsZ/7R+jmFui5eMLvxs3qR0aE0jCA7lD7A5jm1yahl1sURB7kPU
Hp9Qll+wGEHVhek2FKIrGY3NKd2qBH0e1sfmjg55Ny0mdmN0uU4WmWSN7W3GWd3q
by2VJoIqPobvcD5JDMLxLeWNyz81XvSsmN4ynN2ruvY=
`protect END_PROTECTED
