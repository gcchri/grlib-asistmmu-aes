`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnnvbHp73qGJgXmVUkZqNppKSspIREq7sGFPO9b1nOgfZGt1VgkAsZ3ngSEK0vHK
zuukcnWTOhruCEOwiTPBqiaMTtN39yOL7BnAts39awy7k2ShrrSxH7XK7Tk0Qj1V
1w+mLOEINcXmohO3bIAD62YFaC4rk/GUa43mRyavoyReAkS5+/12V4f6s7qGc/3w
OMo6Jj16q7fO10w9SRJKlF+EPTfcT9QDPVFhmdWjDHx5CEwnbNKX3BKEK9FyuIxy
XO4+VEM3FKeKshR9EreG5hw+xV/wcx+CIFzfBobAZLF85uT0kEWE8PMR4PZYe9h/
cDP3q7tJslvbb+uzWvIdwpEToIrJRlnDYip5jP2V2H6l3xD2Utk+D8vzyqC53qH4
egPYDQDGCJUyg8quq4EPAV+rGhFNPgvNL3lk4vMNoi5JOELWhMQ5dK2CCQsAqpvR
`protect END_PROTECTED
