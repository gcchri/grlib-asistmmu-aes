`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpNgvWzw+OU/S/sxwXjq417X/1nfp+z8UZREuYtX+Q1OkznPsdH8MLbcjXy+FIsK
7IMebxyYsp4j9dbNvaJBIthUaxP52G7vlKYA6pjee5ytYpjbZQfhAzMsXMKWAMao
358fo0wRzuw6S6xA4SU8xAosrpbZQQD3sxI/6JZF7Wfa2dWfyix6B3599VYxv9kx
37RIvnjwJB9t7VV2uMlbE/YnCLZ9gzDu5iLCnsi8XVltgpl8ByX5pS0s0gvbr56r
i85vyFSmWtuYDzxWqYLusA==
`protect END_PROTECTED
