`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCQdU0nn61BI+geT4PogTbXFZXN96+B8kNebXxZxLRYD0qioHOB+kgBYWkB4fUGF
iOiUcPQRp4MTjCvcO0Y4UkcS8ujHh7u3t6OZQx5qKcvJxcpOp0zvBtW7ENgjtAqG
lSXgVhWimuLBSguiBkSdOTq2PIM3bhjSprqm5sJsMGxUJRnR2VvPlNBNb7bxSQ9v
WlJfpjBKJVPNzBnOy6sJugwvGOolxX9YQv+pZSjIGjVYTk9Rg/h8dVSEPopSOomh
YXXEirX6daaP2t13VAB2AZzmywNc5B4b9n1cGa6+vuX9LEN+gZYIdqlec8CL3F4F
Kst2tK8JspEcYlNhanhE5Qn78nshAlVrUpQnfzcfCVpyxR3k19iDAAJLpOh6VNf2
rQwyIVfI+IEuxwYWlUXjEM928vHCIyDUzvXG0LD0ZPM=
`protect END_PROTECTED
