`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N2KCqebIJSBGIjXhp8gUrNY9XsPsx2E0OMvhPZVBCRnIsDRpiVZeq6t8t2RfrZao
d91pTRzbrYRNVPLFHFcymKu87DskzCYc5MziVWQIAMcCKkvELZwuEBwRHMop7H8Y
HRZCMN7AQk4czPZXFbvkhRdZmJ+MrILhz74C+teUF83QgGGjAD4K4xz6tnp4TeJf
/V9R3wKt4CZnosbxdPUBoYBCsilX6Y+wDRIzpCfi33GeLVwC1nKaHke91BJA0XtH
LncW5cd2fJ90bXE8AucwwAmJYWw6sr1GzRiD/GKhMI5sGEofvtkOBs0z3Q3YRbd7
xhW1pTOJjXF4O1pAXucnMJ6qYJWAfa/ia58azZsaHg7/bs6GGV26EMiXhtIBGXL+
SP8ddHM5ep9OMeKi0qJx26KA3FVlyzCwC28UQiq2DezQbwDD8RDodSozsPJxkVnP
KB6pfaO0OA6ywoqcssUvNiNSF5NWWC45Ywdinh5/bvT+wpzFnGUicNfP9hcPEVQq
T7TNsYuRbOtClosoe4iwrUfs1tMrk1i7fiB1rK7tP9FZXQ8/Wks15yIr70itU6y9
GykBk0J91GvcDQxgRaip1sWgtXyekgY94uzL8hq9g+o=
`protect END_PROTECTED
