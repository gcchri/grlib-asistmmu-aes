`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EjIoO5pPLMMLT/PbR+bhee6cCISHeEr81OPqycCCENYtCdRGGje+1IpxAs/p2T/7
Bl0Y22S5Ey0gjJnv6irYAOfkKLY7oLL4sXji+iDumzADURsdMnr5phCn/igvS29i
U7RStoOJQv2wGIOX3lwx3CrICt+ninmRTPWt/4LNlJBZPXEyRoFtcI9SZPdRHGAb
+N1v1o/qKO7kIrnjA2gp3C91Z36VZsXJAgvOUU2TnrdJWQ8e+B2vv0lI08n1J6st
oIfcDtHRKxlB6w5XUjGjm8aTR+EOqkvU1vGmpmt8b/78L2RHdHryy4eP323nWqGg
wfWhGABEQ/JY93yK1N81V0GyoUgAIQ5g3XBL1fnwc7vj5MdiOIbRqXrEM9j2KEKi
VnuNBt6FRV1imlQYd9UlZHhQwcWwL8/svirOXnFlW2KPGv7lMbAR+lIgGSBjZrvk
eT7BBkcoDJWqY8Qqs9I3px9wYPnkmVGrsjPaozeFL5rCtxvESHMSlNiaxgdL2ElU
izHVHI55qRRnJ17hWshqTmpDUOpArW3Mclxsn2xqwzX4tI2bWOmtPw7tVOlrHaos
Mv+dz8Q2R7ZtAqNk3AI9VMO+NehZ5RAsmraT4peGgER8ucfhXiLcR8FXdyiiXWJ0
x+xRrVVoQcXeUZwYtJdKKEqLQNZUatG4yi/hFh5hZj4ZtlmhsiUKD0NuMqCvZvfQ
vIp1M3rNmypQVqrI1rzd8u/PYQYk2+eUKFDTPkIPBI8=
`protect END_PROTECTED
