`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0H+A+L4n4adAw6ymdhhyqUydPlkPQKjBcFJYPapZWxz3nn4jSgPnGYuzZWrr2ayY
Rh46hq3LodelJpUnvNohEh2lXQs4n5S7OeZUUJA5B6ykUQC3qCizBQ9+bQRZf/Wh
aLqwDFoklgRv07OFVO9bgj1K3pONp8hKlSuTU1KtI3f4Hb770fkM4wCJWQgGl97e
QaldyASqtaGg9wWGLHX3gLyjdUhClKN35E1EPSTeWQaW96cdrStzWXYQmETM8gKB
1y61sLqzyVNvV8Bq9Fk/ZNQ0HGZx1mc+NVfxuQdEHMANPUL9GftYdNxKcQkma6Mm
vatwB+Tikews91ThGHPEqLz/Re78W0Jxb4RC0mlVH7I812ch4nSW+njg3cB23aoK
Oct1HQ0uI7IJ3KPDFVO8Xg==
`protect END_PROTECTED
