`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NVe0/GrnFph2tRKX8pTfzn4IGNaqGO6xiEaA559RegmYzBYKjPQvehziMbDp+NXB
kTcC501qLfAOUwyPkV5mb2QW3d+avfdVfFbYy+QpeVGRySev00vmOcXgslAYtiSW
lqqUdIps2IFulZadXXfPQM3uTjrtmjeJMq9as526kl6C/n2EQlrzOhz1DbpI/799
YPlJ0MEkgGO5QrMPGsC8SC1AeMXI9jEceNfqrKtBtISBBi4dGxeOYSRV0qjSeguq
RIzgRiarGF31/J5WRR34Lv0oXpUaFq4Uc6N812qI1PZen+UVeY2L4BJS2rlBKLEG
ZDhV7PjydQ44SixrC0hiOnaxIUKUQgu1bOZ1hsdYb2Pgc0JTzgS1mazd16VW4rCg
MdpN2XnmdmgpID7D2cUpW7USPJwyOeGSEuWwQl4CaCE=
`protect END_PROTECTED
