`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tRpfKZ+M25XymxWQSxfXZUYzToarsFkienvcNMQTl92ib/lJvQP8vQdxlEFAJDZe
KKxygNdsrlpE7tadqbwqCoTRVovatJzpYQXZxYbPrwOvVgX0o0aBH/Bfg4KFAkc7
VaneMLjjE9r7WyDuKbkQ23tpUehE0nL4mIjqmSXboP/Vw0XiWQK08DR7v3V5sXqe
woaeFT8hyZ2NH2VyJpzlaaW4eURpRI+6tYmq0UyNzbzWCNRCZrRzmfo3QA7/nooQ
3moCTN/Nlyhktxzs985CSly+xpIik7Knts/csPUMufsTdSHSwCuewlCfAGlyBwBX
5jF/HJiWv5Y50rk9Lds4MQ==
`protect END_PROTECTED
