`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ma5JmMvipMQTaFU396PaA+eBmXo9uvlFMBa2uU0DAB3hXw0qJlLB1QMlELJMkTSE
CWG05FLRI+LAViwoCu9v08xq/wel1bTrvvEJ2t2aSpZG/9DPe3mKVPBBBZyff0k0
CmQJFly06qDd0ePRb6xhSbfwfc11trhO50x4s8W5Hs3JI9zNg9dsrERqabpKucJ8
ZIKMFukN0YWP5QNF1n52mIu1bg4WlJ3nd4TAfRm6fBfW5CfT+b5IaXgO8+IpQcVw
NgkWVkceM/hzmB2zWFF7/jhyv21POckDISS4BQ+yldmhPlYOQ55NAOdOY5JDcW1x
yNJ/E6P0IukA6wMi09qW/B9KM/ZiiZ1R/lsTrnzVT1ifztpLzg8G9TMorihmMMvp
qGOfMfcxCkRE0j4xlfXnfRwZosLvV7T91Y/jqKtMLaa41MllIbkmKioMDSuE+NAR
ffwPJ9n01g4ExF7R+47cB5pz/+wc9XxXjlyysZxBSbjN3Wua1alEzG+CEYsHDdoy
wUcTqnI/Ft9GBX86TvTRVrbgc9OE2w48zFTH1vMX37smNptnU06jFvzgO4bqJuyZ
p19OGQPSS+266Fi0YcOo/lz/i4HRTEtU1PGWRwBOhEZUVw+kShgLW8Feq8LgJZBK
OcICQ1omHngxRiydpM1kVlTGM5Vge3i8M4ekw27MWmk0TCP4NoU9En0MmgsFJzaq
SfHosuobrJSLoS5iJxhqJe5cr0FxXUFTWlKt4RQZU8ubTLe2TBixjaex2KVQB73H
tyOY7sQQfdJHgoDTa6wei5H4pwEjlt/4uInxAFgX5fA/xFuk5G1k75Arz6eunTeK
FtFEubylHmI8nupmG6g/x1eN0cOhTrbXX9SArbrPNLVzCpCIfXfgrOqzV8HE21gu
GtPu1QZ6Dxd3cmotJN9Kdg2LX5ZpNdfNMTqopJjXfEz0wOYW+cR8hv4MgowhnTrn
+0pfAXYF544/Es6+k3rw/V8iSTLSm7lZpTbSkUamDkRk4JdptpiApz1Urr6FYEFq
BNBrffLVkW3gwlOZszvCZ18zwPWC6B39Ft+XRkzgiZGtZrJ9tRNLY1ExKOHMKCr4
iJzIQpWVYgOk9XQxfRinrrb868WiN6PZPlfE1gSydnuZD3CyS8eTCTzb+938tsDz
ijgG5B2HlRelm72OHA72lXVup3pfPpjCMwy0a5A1FhKXBfC8eaakokppdXFK81ff
oS6lChxeapvcRcQH5/5pyFh2co1T7eF/l++K4B2Kj0Nsx81q4OUYyK6S/Wbn0HZ7
+2g3CQKc3A57CyzyTr2LwEmFp5m2VJkRrtcuMgGYaX1n254MOqiNvMBroHd6vuIQ
8km9OTFc5Sh1ZgeOvfXijfyOEHdBfWH0xZeyO1Fo1uTKLuLd6eDdHH5QgMb/nV07
FEsTJhK8X+w1Q4qRMgUlAcgkZ0gD5oF6sCBRFsA2aVZd5USLT7g61nB8Ez0tzxTU
P6oRU4IViS5XkGNRaiAbkOSod+03qDZDyNBG1KrHsJsoPGAfjVTdDzg2Zb3+jhNQ
u7vjwerCdepz/NNpzfmOGpFxSWwz4wJ7dFu8HWlbgknqGfxiW1Rd7HKlM0awTzVU
wLl1EXHbPicnJbbqgWX9SLkjzHebSuspsSVspRhirJ75LHg/0XXIseC/MLmQDuYo
QqP6zPP9m1V4PdPx65HWioDj2N9RvnAa1ANKv29Z4cvykyjEgtIIvw5ccQx1lQxJ
ZzB/lyRqb6sGIug5W0YlsFy9cAVju/E0O0Q50irqrE2ZGU0GM+xdIfJaq6wMYmzf
u8pFeqfy2rl+9pE5aI2ecIjUoWn1xkRkhnT6NfMjj2pFo0wZSVTDreFZQKqd8vcF
a2MZ52JDHuOgpAqHKS5koyuHQwFgBe13mx95r0RPar89RRKAa/N0o5nNQuW+3jJj
5KBgw7Wz6l6JSjEmSio4n0YUXdWSce7o+UWEIuGTDeDxdWHmf7WRtRuQ+CD8mpSn
AxtDAfshGfryHGcEM30QmzmDzonlhus/5EshuERAjtarPtwpmI5+HBwj67k6P6n8
Rn4Q/4EPviGy2BYtJiMM3kigPKdB2xjn9fa5zOZfDtjf/AuS6tZJTdZap835hLFH
rLy55751e8hMsnFhuGEfDg90EUWJzxQft6GlhqAAn4Pkl8lvqKJlXmfQPekzWdkD
Nn8+7JOpe1mSlfgFWjIj6bikGshGQuGdmLklyrVxORcYhC5liJEuOCzn9PetbhjG
ce4ZY9O+AqU6L6IuMimNl1zelBKtH7pgs2ks8bJtHZpGgCa90TOlIMPqSyrvQKnY
B+5fszLWnNwsxACFtymOPYhmYBVugB7gZ0NvJlPFMEjX5sfEIFuPd/JaKhPob5Oc
3wI+CGxVwu+pqegjlIAhSXxHiip1WqjktkcA9wYpGIS1L6zyvYLYXYIwEymHePMi
gCGHEfYnmXX1yW1TgrFjMs7Nb5hMcjmZPCHpRIuK+73kDu443+dUAAqdSkDEUOCh
mvREbbs1cMnNV5nRdMkXjWVPNhbc1Z3pujdGGf90lGbZaIufBkw75uJEj+Rjq368
3+0FNRLaVaZntgndQp/h6yqoHlt4m4PQCC7cfC9xQz5BbxQ3IAFBYXIn19J7hslk
/KN8CgBDf4FdnuKKvJYYKD0bclRYrGSVS/NME+VsGmu9boSvsUfpVmX0Z2uarx8+
SizRF0RKr//qKUoMFk9qgw==
`protect END_PROTECTED
