`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jk2kTMeVBN5lvxe+Y5p5a3VnZIfv3z7q/24f5Zjhrqhv3/ylk2haIfXmzLT5FV2r
aLBvsn9Mayatx8Yt9u3rdnhNuDycIXxBno8caqSCslSUooY83pfG8dgWzNw+PUem
bLS680ESxUukVI1O2H5SrXP6SgN+qZBXMArYsw6d1Qj3DKjoaRTgR/LfMliYIX4x
GTXDiWh9cmE6h+jMlWHWkqLnVJk7FGHJiIO+mBppROhxnTmDVULHtaJfyeTvfXd4
VzsW3aM2EAYrl/5F+ltir1cYy3LuwVg7rBCBhRO6Rp/vIVfmzGGnMn2nt2vIsPHL
aVrd/taObVl3zd6nlEHn23ZKarDR+PKIJ1AMFMyF/5UTQkew6Y44wqa7kAYV6ri6
iMzFRKtK1uZFZk3B8TzRNDflvPIB71J0ng5ttbbWOUpB0klLNEjZixC3XCZAXin5
`protect END_PROTECTED
