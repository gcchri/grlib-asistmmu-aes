`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZKk45zFaT6oXaoyEqcvuMVRo2pzAco64HnojCjp7fa4GSPnXoc+wcb7QlrBcbfJu
MeHJ47ppmP0T9YR8k++zLAEu66FTfYpQJngWNPhEvI3lWLQZhzAfdMUEE4utYaBS
vVM+ORkyr4jG5/ZBWiZTRA7k8d9SO95vJpBeSz1Icgh9PDtHQjKeTf1JTTF2bjGa
AOZjJbNqZBiwBXaAFrj8h+KMzHcpJwZcb9AZY+Rpg7Kr95Q0v6Lzb0TVqm0Doe4k
tOYXH/J+5G8A4us+3S12hRTFTJF9kT32vz5ySj4O3unCKhHgZsBGFJ0sGjXpyD6V
k9Lmiv2GiUgBhHcFBXRW6LxC5BPG/5F/orbMv1gGrSz145UYaG2drnC3rmpFRq69
6QsdR5V1pvT4YEMk0tfssCQyVSEPGzlLPzw3NYMphOum4oYY8HffBRoE39/+HIqe
G53sy7TR5Bh34+34TBdwSUok5ha0UQa4bnZsaV82hq7Eg/buoatvNCM3jZlv274D
rgxU38kxkzgKyfrEae/5YkrsW3rLxuYwb8YpBPF1yRApECY7lU2NincxDCpOZWb4
`protect END_PROTECTED
