`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C8foVVTz7o/2314rCnSnnHuhBl9eJCyzb93vXAAxDsKWFXbLJ8w7a4aUCWz12WNP
ftSOfGoGNB0p+t/NHfZ4/vqSUTIDddUaDH1tbSfnWz6y0jGpMdTI7B61WzULXek7
xSllOzlzEdIhpl5kKF55cIvcIL86vdBSNBDcMxuCJus7vu+bP4MObvjug+V/yj5b
HQfWkNlRVSK64iL3bvOhDjQLLhPIaCFJEEPqmPRednyKFLUwttmqM7asdWvkHKTl
5x6r85lEHnmLqc6QncBcxQiA4tKhGNSazhNFBwyTwpO2QUqBWkkQpnFius3C+2Hj
m0O/mQZS5bm0Mnaly36uO3sh+M/rS1RgGN4d+/H402+sCkc6Qj5Bo7L3e/lSvbVP
lBFbcPAB6Z+hZ3RQwbVgGsN6M77VTL912eAhXstUFcUtA6E26x2Do4HaThEzIIoM
cvhKbqKuKRGlUPHLuJGez/biAun1uyEwUNv3XLMtzzQ6cEQ4FHiac0ysXtq2sKQX
3oKY+zVX7Bc6wraXd52rHGToOPsJIGl8Lday0rGK7/08PJFyMg/cveXcvELzv8tf
8xxHieZCPmUOo+0uY0BBf+AMmjIqfFNqQCXbhRCYLpGZ7a9ptLPs5OyYTJJW5Bhe
pbrNmqwrszVSIQ6PqzlvGpAFm7lxaBXVxhE7S/4q/wFHF+Gf2kjcQaAOdm7xDWrT
qeCgGoE07MQuwpMETspKiTJIs9elyvfBlLIA5C/2B/JseKYlmKedsmb1UwmK+HA+
D3lRovfUk6yLsmKq+LxMvOn1tv9w34Peoe6ywuHiNxayUDqmL0CTizK41LGPPBh6
EKuUdyk4iTsVC7TtrAz/28wjig+W3aAdsjJXnM0AkH8EIW4WuUuW2Q/AYXrIgAKT
24tnXAToAW2tV6naCz8UmA==
`protect END_PROTECTED
