`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q04B5BwCx3q6OvWtoJnkj6foH01ohNWcLLvrbyjPCnQGZKgHCxEXz/DbwhWSRgtV
rBhthNM8pmWVFsciIUYyd02K/flm2b7AdKCkh16KJZMXXpUQYKVYYBDpRuHUrtAP
O5OpE9q46gnozZXnXP0CKlSdIteijYa52FdwsM2q8EUCcutFVm2cDOkdEH/AyxDe
pWP9YYZjfUnMjTpM9ClTAWve9vdamWOnt3Xg1vn8Qyp5P42ObIELPtj+qpFcPU3g
1bEMvAVNbsSQh2dryF/yNgIkjwDvNor96PAjlh/0oWdScbydsowsBvYJvSwIyKa6
bCBs9n5PpQFr4Q0WIQFWlR9V5MlOPmSfViZmdy2yQVHt92OTsekjWHjv/cfqhIvZ
KDsb48WyFEgzS71JVi2KT0qtKLhIulb0VhMQLZjOecxLUL+HEOg57efR9KLWBpBL
2dGqvPCM61UwF9XN/q2DJ/MzPzEBopQiCkjyFUzbSH4dEXK8Wjj+7r3iYN7WeoRS
I+VqT61FWzsq/Zy7XmNJa+u93N1aJFxCaj0tv80YDuJbt8uT2jSBlwi32xF5VDVZ
HEpQMDNj12/nddzsan7HJIdpaOne+4nmLNPxiMRN/ppqmFXyC+Ol0Qy7Z0bjAw8e
eRVYVW5b4WzM0Opx+/6O31+w86oOq5ZGh1fK2zqxBfdD4qFoKNtgs2NUT5ko3TPR
Ec/g9j08s+nVLdqmVVs7kdPamnR6e3vKc4sGh1Xnq6fxDlrZSG29a9UfW0d2LCXs
LZnvZUbOkVW8DrDmQt6Zj9y6jiC6Ghj/TQk/sOC7719f20jhEwRw9DAqQuy675Rh
Lb0ST7ho4wWCaF63jLeRiyFine10YA2KokK58kYRmUpV37DoMnxOq3lMsDOdCliz
KpndkHbjYX/LMf+oVALzW+d2U7QHpE8DfpfBBniNd3Ocr32zzCxg0Dv5IXCSpAY1
wEfEF3wh6wOBj7dmqp0aixnuOfXqs+kk8fe6Sk8l9bqESLk1Ja/9sU7FI1kZtjqW
xkl8BYxsVRUn9TiEnFIJjo5ciMaXeYtQM9KBKuWBOnUoZpf3YYREMy2eDH1vzMKy
UoQ6WOdRXRuUwAD7Hk85e38ovmv4XQi+CsyET87FtJN/JPuJwdPPyi65Bz/IXw24
pa3uFbQDdMtFX0LSQmTpRwUNIYJdJanVEEYKjxNiwcftbKli/p20ePh50H/qJTD6
87UbsN2Axb5wk9V+key5CA4bmNkWwMRGlf4BCUQJ5v0VWJV693QE+pt5kUAzhiI9
eUTJ34S98biw/12f5MlF+xbjFCO8sDA7F45kSzZ/IkmmlOUOXouDavrZcIqwWJQc
P/zX6XKOXJG11VFSxpLeFrONlhCY4RuqAThXqv67FTLj3C7Fm+C6f/96kkUMH0lh
O/RyGY+3IeU19hm9sVbpgI27nM2bR8qxfca/9whzE96u2V+Fzz8TXPvVvNWM9XS1
0PZkl6xKLfq8+v8ZrzE24itvgdA7M5sVmLGBHj7jcHSWQxreib5JI6wkrwOFqTs6
+VKHxep8ivnD+JvaAQwR2GkFw5hfLwWeVjPYq5/Zdrk887HW/TaSkK7ZeJSLMUYf
8sgd9xAcnggWyoz+ROHKEEFX/Ehy0xomiISnDnosnJDDKmo0nhYs9kuDMft4fbGY
acMywjRQmqFTSuQgMYka6CG51RKwt7XAXirwl0fMPkU20Qg6ytaTKElWw+Yp5iku
ZBclYY1QOjfiqWeUDhFUufhXMPvxEXhwRDC7O+HDjO5CGYpdPzCZUUTzuRjuXC/7
bx5SPUNJUsDpKAEvro/A57FpXkVYODg6uFjiqf5Lhs2tNSFA0kh26doVb4EtlFGd
DYaKbpM5zWz1BJsMyQcEM/12ZLHVlbrY4iGGHFAPPwTdggFdknIqV5EuPjWJB5Sl
N9vNfmS3sHwcSJ/zs4eGY32vH6oHlkuhtdd+nwzJ2VvJ/soxVJJzVxI7ALGDr93d
6tbmksDWfvUZj+YGvFWyzhrOWmJBqdyCRlp87N0Qwld0n3YFcCGbIhWaeGhXI40B
D2J6YKgm+fiVIWh4IYiwVxJHOclOiNx5vf6CUH2/XSnkW/wx9TVDYluBHKWw9dEJ
dFiq1XnZGwPNyxoqxc4BplmPkJasBUAV8ovw2g92PAO8n4m7Edoir1hpUNZq5LCW
/WFeRI2XnSJHz/WlPg8Ly9PjZcxYC7Eaf77LOwQewmFhlIYPGWdKeEnzdy6Aj9Kn
jQwVf5IWf1TEoyC7KoMqCGnmLaAxpma42xESE5dOP76RvFXjCmsBe8Fj0QKIcnXC
1R84o5GNTLdVOuZnYCc9M6BrQbpcfWXN/qsgiHdE5rM1AQN+KxQD+HeDe8ui4fNF
mJbGAJvdkyO9xQ2fDmXQ3/C3aCxleN0YOftOVrzasxDYTOaIl/brr1mbCuppiUlI
oZglAShzu5MVxukos0Y7LN1bUHi/TwfCEhwo25QtVjVjmrcqodCPYw9nR24yxwPU
`protect END_PROTECTED
