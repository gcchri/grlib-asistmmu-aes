`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VIf3rRmSRVX1q0dT+FkvAhdAt1cTfHtACHSerViNMyXJG0XEanP3PWYXv3n7sgVI
YidV1f7VAfsuR3Lv4t2Lsjq4uySYTJD2MfAf2kTpXpVj7AdF3l2ywNTAwJLQW/9O
0SG8itJZn+EBi1Iyrj3v1qVUXI2PA1dHsthsRweWadXNKKnH7YycUwxn2QUHYg70
3SANLdxeAWWXTdSendIxd0Ug6xTownElyVqSAv7O8QCAjcxAcyYu1ygZ0G8LOY09
t8CY+xjxNQgG7Ed0ti8r2SAiCkMAXq7UmClWIBfEQvMtYtMy9Q/MEI7XLXSNFfZO
o2wgrHimhar+BfZpQnQV8ODKNSGoUaeYFC5thYxtwNVNAxD/ulpWN5UqALVZ1l4l
9T+yQ3p6JBmxkwEC+7i0/xFHlYEBJU4ZiH1AiClPPfMkHD9K6y77rWYTriXyLXTP
`protect END_PROTECTED
