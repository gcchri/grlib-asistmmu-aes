`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wj0Anfef/gSoumOn/+3Qaj4njHPHWkUvwM7erv+wdFKDxGSUxzBraG3lSI2QWinq
mQ62eZpwUNX5G7PoSItVCAznHWwZS+3dCpWRflSihdMddpfO9QJtHVIlQoruvBrT
M3aB18rtYKkgUajPafmdPlqdshDdFdXnQO2Qn0dEeXnqLjgnDa3q9SCJPWPosCB5
HLzo8w5UlqreC35efZ0uZGM9lfTxqgB3NipBhf/cq0JTZRtO6HImlS7VQKO3Xv05
th51rKoaKe4v4ccSw27mrI4gtZDZn+Hn+voSa40eUubW331OvY+28VP0BpDu2str
BAxfXruBMHG3i4z1VvnomTBvdynHHBhyrZ+f3O6RWvVNFZZ1AoDbkrtj7M4b4+Om
GW0jm+g2HHE/ncFEPEQBd0LliuaL6/JBxtK39k/vHI8yiG+XMBshfeHZKX4MVIlH
QRZlTiaSsBvFac1r5MdU/UmoZlS+TFj/NIKXdMx3weAMmFKyxfCLsdebhUgmjzd3
ATXsdkeW4agYRqwqkk2RJbo4mnUigHTYdTRsDROopdBAQN/b9Lkrzfz0dimSBBW2
T03dEk8vkfPwegzfNKZzWPCHNEdq27+vbn1jvmEZwtKMxyJ76U1q2JMjijq7/gk3
60F1mD9RkGUWWeiyoMfHFC39+1/d03VcVYVMs8/IRrOh2WUUvqPBT5hItlUtt2im
kV3vDg9J56JNpjOXJx2sTfT8uLXMtX1CX8hH3y+wdssK1X7ykub5zNQ5Ig4BSgJV
N+pOXw5tp+EUg8BQIEUpVR8yuKR0tV8ZaZBFr+mxz0JMLvqrplAhNwy4KEUjOnhk
BwL7ekcnLGNVXxHPawX4nYeunHg1hIzZjm0uhZMMe7bxFeC9ThdLTt3YdB5A/Bih
1DMBfjh+M8IKHCFTtF7U5R0bSFNWtEQzdKPyVKfxfs96Z9hZvizFZNsqr605KJT6
IX5NVxcoFcdlk5J8D29J5xOyfiawvNILzmpK9OYF1aB1PqvUdEp9NkpIM09kGu+V
VZs+Ok3gjiFlhJZSTLlgNSBcHjEX9UZpwqh+XMyTBpTFcHnqqBFsvUR2757lRGcq
7/Zkaoni0s89r65U3wcaklPeVAkoUt5CFK4O8kcXgaCsp8bUzC3GxwFpLX48LW3x
7xOBi3fyxVIn1RI/PcZb1e1uBzVtmj1e8aYlgffQ3vXOKT53bok6PrGo74kNuoaf
4q0gMTf0gsXUbdvBpp9E/9GGff9HGhprFAn2+Jt8oU0VJNCkXgGQXU107Gek1cAi
VapST/kyllXh/18KouetWeELXNat2redbsdONwvxADRAZ6ab2kTERkd6f9ZaRxHD
rMxuzJxhmhqN/zu5vKeFsLgX2On17+P13Gjt1Cl2xaU=
`protect END_PROTECTED
