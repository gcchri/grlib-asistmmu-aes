`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mfa8JjIu1oJ+1tcj+QqrMJqaQCcu7yFOSPE6z36w13on63Lj17kvbJIThKT2N/pI
7TQU547OfDfgb9cc8Xkgmij/mFjzwfR70QLk9Z+mFCuEm75vezYzulsLim/Pt4+O
DSi+mm2yJ1mCibUGpmjHZJ83U0GE2V5O6cM50DmSJGA0PDyZVspbPLej/ti9eM/2
KLwdiGmFPxIfkKjf+LidAQDlyoJ8Gb17JzzoIRiX/Gy3gduzxqovKNREquhg4kZ7
prDeXf3Q5OC95PKgrRVvGhplnZ/GEe0B/Ale/1/l4j6du4osGzcETl1tIYZEomP1
5foBD+js+HssThliSWSrpx/C7zzQfSUjBaSpAoWi+zSi5f8W5jU1dLvDxg6+yABs
m+Wy+thuDlflC/s5ng0pHxMAZ7Jt/eTaT073J8Z/2MVTY3kmllfDQ9vfd2CL5xZ3
XVd8P4lxEVcPpZgm7AulWIs0DCRXuMDNJVX/phS/5XnGvlt+AeYWQA/eY08uLhty
bukvbO1oK13vFU9Wa47qITPgVb36kEDrDy9gabRUdDeE0uBun+TR9ouk8djrR4Nu
iQzYLCTgdHnOEzA++CJQCvWfe8QWsS/kZle8cDcbhbvHTUhUL0dby0QoFjSQ/Un0
whBLVQeWTIuKneRy+L2yfRtLlKuM8D1CGr9b+csweKeAgbd5qw5Wb56+ivAS87Ts
Gc2XRn2JRSS/ycFGmWQPmmLw+/c5yngR4qCp8o8tJmlSSlkxWJlL6O1JoNlziQZ+
lCXpkRwfrWOak5CXgL2ngtUY3m+uoMQy4+fvV/IxxSuo9PYgaPGEkQfj7evYNHEa
RpRbM3TP9Gacw+P+YwVTk+Up4UTRjOA/SRzTL24IvDzhusWMosEK+fZsj5r0WFgj
GLPAQXBEfHJggV/ainPg5HOQmsLIELa4yF80DQVk0vTvNgumUETuzmqk9dMjMuPM
5/InI/vYqxXRICPGfV5yR9fk2StXDORrFHEspTPIVyyx+yDkh6+RRVPDfCcFx747
ylM0RdUF6v2LuyLKLS49zJqzk5zOHCjrYxeufXK6Qd+BO1dGF3tBQ0mHRIbT1E+o
krQVNHDjRGr4ivbFSc6fEwe802vQpVqywsh0A7f6igLaVqUX6OrEBdDYy8MQvE72
L9zwv7oNVfI69hK/6eQFyJxdbE753jNukc/4hZ08wggIZdkvq9VwphR1bE7N8Ap+
c3rtPQsk2uhAxxMnAhvb1g2bfm7G/DgzoBntvbaTbpCz4HKl6eWeFC6b8B9haRkl
CUOXDIrQQTxLbs9eeTJzeHwqJ8yKHzv6V/7PKCOjoU5BXnqWHPTRAKi5S9Vqm5ku
jYsuBILzLCXMyzkgIWOI3E0tTclN64suVyqRUfUepv2DmQyFhyJ9qjxM3ILPBFej
lRfvq7tez9KmPORAXLYv97r98wAeBRPUHIgch8kkovc7p5ElTioY1I/WeH5t0dG9
hi/NdSwsrkS/DoPxPnMrCrdQ3aWCDYN97Nv2pbq75qarwdhIlT4HFVjEY3PIvJTc
Bvj045KrvgrBv/V3ucnYzUbhxw85S3kYIHZcjhtfIeN9Gp395uQg+Rxjv/x6RGcW
gPLokUyAeM6zup3kVb0SQSBMolPEQfGkWfsTfeJUO0EGaGpkt2NqYB4/YkEm3Uzs
evzcIpOdXY+qOQg3EVEcIQIRmzC0WztLRLAZiMorS1T7HP3iCZ9OnTyNp0L2p1IG
KUqO5P0sv+fD06UZyMidPgmAsMMlPHsodtRjNKuJm/j8PWBayk9xDZgBRz3QNVyt
4wni0H6H1lqldfnK9Gwb+uMVysbn2AC7vE1BVx2HRv5QF37lZAQzRX/3oWIj9t6/
5PRz3xinJWcgXDVsg21hDtGxreDvf7FwzA0QilHGkp+3YQTFQGZjN3NUBKTtnQsn
MkBdHK5VE8HlANaBNJHNioH70tGF0wHlNN8EssHWyJBXlMU0Nu8gh5lsGqx1VKuE
wvU5Q57ZSDtsRnHassTFJ0wXVfdr9YeVw5nZm0T57mEQRZnii25r6qN2lKKRZb1A
POyAs2GiFOQv1kk8EdkYWHR5KtMb8s9pPOpZXbQ7ZvAqQ8G40tbEiV/tE04l5cYr
L2v6iEvP9L1RHv1VSeoK8jC4pKqNTMsadg78khCMFqj9IYubZGg/UYGqpx+209j+
Q7s1/EqPrGV7hO51lX3ifg==
`protect END_PROTECTED
