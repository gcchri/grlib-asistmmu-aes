`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwWECeBSX4j08nA5SrQz80vBlTxBkx+7E69SSSu68io0XUbofJBNlM9p2/GcdODO
VvjduTBFtDskkurX4hrV26yhLXAUNPfdvvPNBGNKEjb8cTNJ5hPaslxUrPe+5lTn
fqr1RE+mdd1MHA2vMqgS7eiWa/FAAclu77E53wgRMD/z/Zn3jBC0hA/TztWwSZRV
DKckMPBAcQ9QjeAfhrFrQYFpioexb44yYJYiJVNgkSmhUa2vFQ0X9URTN8Y8DZFT
0BslFgbLbT1nuUvfYj3HGdpTT7QnADhy9OirTO3hYt3fYHfjUxNRZIP+dSsdkgBc
Bo+JLm11WrMhq4D++jQeDcQ4e+W9/Sbbe/U5nFN8CZ4wT4aLDlzSVSJiLZ7IZGK8
9sZhnEQXRQ9hvXG8ICV9PazCqb+0UFYrCCtEKNni9UfPuFTj3V7js0nmBVPepWng
hQJYqdaih99+zM1268NFCli2ays5/V8p4gw7HtGm7zOQ+M+56lzSVjAiUTlcoQXq
MrX7Ug02LoGroGFC0ckNCnYAc4ugY+bGOOVi68FXMFv/nSOsnBY4xL8sZ3rUGu2H
j/eutrR9cPiNjWKeyZojkJzdlHtztw/4kprmHr9wLlEdWSb97TkyBkTT8x6V0C/1
cH2b29I7l1wh3UOz2jouMK5/ijbDb5z88jwCWEbo1sOeadasGpTjC7zf6igXF9v7
V9cPF8qvW1FpToXWnzIqHM92hVS67RN660RYQ5O0mwKyZB4VfsA9ZNZv/73hXbwn
ZGTXJhujJPKQYr05S5rTRHlkodgjhsmfh658U0IcYhnJf7FlO/pIDd8Cu/F32NkE
f9YG/5qL/7miafQ69x0olzBAaQeuMLVJahdj9GoVaDY+/DWkpvDgG+Zc8RNuwm+n
L4nKhSHYXSaFBCaeLyu95ZexSo8H7Kw7jpSu6xp/3O89+hOYtC0Dq2yrk1LZye8d
0e7IsT9qtQ4lM1TYcuamxKpCppL8s4F4WgLJ843SLo3Uwt/uiieYoQk299M5YQUN
NwV7Tu5l2yY9+RZwEPCsO1vYBBg4YmAW+WB7mccTBpM46DjAHdb7TtMdbgBVhSVH
ORTgjglspfsdG3VzPL9ZJxz9d/srqdeTJY9AkOGt3n5NH5Jnr4JpvykZWtxc0oiz
2g9pQVtkVzR00AnC2dbwWaNAYZknZfOnpvSJGEUgDI3WLx49uW2Bi9HXDnOR4/6p
z58FLU21ykRVHzMOWnBjwH963waD72/JfkTJ+CRMBQyOoFCTrZP6h22mQwEVyEV9
VDas9zD0/dcYd8q2phf/yoSmhcALJrkoNzC2jIZLNVXVJrc9uI2HHUlKzksldROs
GhuHuWcW0X/RhkDH4zTrzGVmKu3QaxGQp3/w1SrSREuD+ngNhizR948c4d0DOnFU
tt6xSCelnj9UbvqF5Ol9aXct5aJZK8RT2Ndw+2T+3qRxc+FUzedj1AeaCpvwoyBw
eGSxprmojFD8BfiEckUOg/wAxNqprkGHkMnarkRL/5H9QcbObxxnVEvqwB0nqttU
MUK3MnuDvlYobZdYVDcTJHdLcNSBYETwGnd4zc7KK9P4ZgANN2Qdv7PXdmp6RBG7
BRS3Yf/mreaVB8SV1DmEjToh+s2NSWbELmI6kWbwVRtAtXK0syNioSP5KJuovYMV
XqCCYthe7CbrvwtbQ32dtnArtDE4gVZjn6Hck0ZyrDh36W4TdxuF0uv2m05TubP8
2K66E42lvOoNqEfUyZSuD5/6FtkTQkKPCZILlxkYfYOF00jFfAMOM+t7uRecDL2u
ublYCkpOHdZcWKYDAZl5NXf3hRwywYv6D7Ouu9LvNqhYO+PnT60kU0SR2TbhM8Si
mFQ3g5FBZsSxhu7tYhQnMsNbI9dHgs8SAkwh0ekL4izrOZGc78rM9Ti9e26lP4/D
k4Ttf4N/ZRcILzcI7RcNiAke9gXcu2BwLnXzPohOitLrJhS6srnxICG/nsG43Gae
wmQoaUHAD4RyDDScY6EifQYAeCfNsKJqJ7JvRxX74vrVBmJjpyBbbMw6Oe4cMsn2
ZJNuzWb3ajRSD7Bx8uhTXoIiuhfyWwkQU1BJtre/Mrk=
`protect END_PROTECTED
