`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Ck45AWY3BZDo7voY5CxUS0CmrGcf1fxefKuRi2mSsGHG2y6cGRAfUTS4Un9Mnpz
XEbnSD6S0/Wbm7lqQH/HJTwdVs4QiuLkvVrmjZabyCsPUCSKPqfU/HCDWh10Mmm1
T22ykQqlGdcxzFxXm5E2InMNjO46X1OSKxkqMi4pOghAdQypc8gzhubxI0wQDKJu
OzSCNMqWVyt/tGmrVsljXnmETc1rJv0yOOEn599YtNRuUcZnRyShT8AQKnYmG9dQ
FFwvXfhvHKCHDCKpMzw+GLEtsCGGvARlzjxsc/khl2pxXYIj2Dv8TxoRj/EeNmI4
oPkIcuUE/HYuNXB9Wet1JVF383VGuO+TlkUbRuFhJVI2ZtMXyuyS3wKaW+ISZq2+
BA3ZB7tgAvFjsOKzxPr89c6LloNuX8iWCs6q2+UFLUC3WbLw3lUN4etoNnz2HlKf
RwfbnSsf11PDgFrX5LjrVbU+M9YMkcBpSz/CVGeDHJMFQEPu9D0/5ZevbJdSIUbY
JqaDuZYyIHpRM3NMd6rmiXQhFrjkG3qZoRTrfR5XTaQHvlNifFBcvVe49ipsY0DS
yI+X9DAatgQFmljnzC3v7SaqJQtvGyvYte4NQzHnuBOOz5jnezElDhhfn1h8nfL3
dm3PeeikQayFCjqyUjmdL7e3yN9pwDX/jnE9gMAyYTJE9sCp3Yqo2095B1vVDtqJ
SGavWtn6l+3Ah8NG68/0z+KtrnWArHYfgKO4FuKfkMg=
`protect END_PROTECTED
