`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLsxRNMJkylTpJxQIQhQPdqlhrv91bfKIeq6hFouXwfFLVKGFcDjy9DOAj1AsUWf
MYOk6IKzAi7XGbZYqP4FFmaOUHU+G1oYiHMsuOmnFT/unzu4WvdZAZ6bZxiwf4Vp
eDeSChbgZH6ZKhsoz4QcphZ2OFuaAuWng7N/n5tRP/z9wl6uzBuIzsl6mTp8QAN3
LxPk9gV6yPjaHCewZoI8/nTc7ZcjFql75Cs1IaKqfybeVHsQc8a5D18k46VjQB33
lbaxPzVMzcX1rU88A5DK6IcYpOfzoY5BMixwmnmfhl2iATliC2f9ZE3/VM0yj8aY
bBN8hctD2T7THf3tcyakIwO+3cyVXsSwIS7AHMjY1vC0mp5e/1RNanl8gXYOKxUc
zCwG6xPvTDZhKh5LSJDOQuVTmhXfLflB1qtWPiK3u4R05e+ZjTz5L/dVAoL7Ynv7
H6D/WegWxUY/JDaCq+A+tzB9xiTKRB67m4sESmv+eg2WKCTIwH58UDr9UaOlubXQ
yLxuZPqFahDUyqE4qIRDAjrcjB5Ebv3F3wzL9feDqErUHasURwyyMuIzFyCirjMf
PPBeZ9XBnf4VJ0n1redMdlYiNFBJjiUPE/M88Ml2//LY11SBXjdiyGhfJM2XESno
VMi4KElS2mlbnX9hT0JwEcsu9r82hxQO9JslWp3LoQJ5B/OQcdk0PWaSpD7G5E0t
gGL8/Ln+CSBWXd8F/UI2ZhozwUvz6nD2Yk+B+TEAeRPXT4EaKuBHV2Ij8eTg+9Sr
Klw+C7iOjgT44LEtmp8Aa1TD1enF63/U1beRJ5iYRC5fZt77Zzcbb0+ZV4KhV6zz
uJo8mWtyB+2VxiijBYUJccRm0LC+aPRYbAgpvHP4ogE=
`protect END_PROTECTED
