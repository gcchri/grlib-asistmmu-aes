`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bl/365YqpcRB/eGd35iLrt3Ox41wnPHumSJc0K+siSjuojchuU+vNpGhu6YwoXhW
fmWtaHUoKtRm/mP36q0FUOHHXLM6sUV8DxltBZ4MC3BMtxlTRMWb4TBr7a5FpdnP
0PnCIyHQTH9kDfHAuu7FhfQzG8iz8JLyPAX87keoS+cdMFMjLM9SdM9/PnKooG8m
5YD7yTOU+RR54S2yj/KENFCaAzBQzSCxhlvkPFzlq6Lx7NEcehStTh1JRISCmIM1
3O9QS7b4MAx5DvaYQGXkYcQ4StLjv3CRHwnQ00kbyrdQPidBTie4/nYT/7hEv8w4
kPBalQPQDTSUBRkcZ+YfJhnQtmAwqCU1PLferXqdqyii4X3qQj/lzCRDSbnPh3Zf
SBiPtxE1p4pMeGxyMTZ4uw==
`protect END_PROTECTED
