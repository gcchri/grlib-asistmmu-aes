`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qm8AVCdaUUPuxR0rMICQI4sNZJNTwVY3CSUHMuGx56CrVUuvKdoyWaIcxmX2GJNL
U1kbc53899Cx8kpIKmtWPtsLwpNe+tG4iT78TNxpOpeesG0wlsQewrFRBZU/V4IZ
/R89jtdgy/Nq+D37+Xjshkg8jA8j+caBocM6R7jDX4jW+GEx9E7VtNydCdLllm3a
x7y6S8T0S0YTdYJmHhmQH3QsQi3F3phUQPe0uDdPwMfLKaEPuj7tWltGH92to4NW
01qA8iuW+LYx070qvenIzHHJ5lmc5N9cWYSukYMpOerBXtfO88cSXTJFKP9Twc2T
crd7QItgRBnpd8I2RcjHi2y2CRm2/ZTVKTLG9bJ6FYR6CNHn37aEWVRNL6K1C8Ne
X71bQbn3ZIId5cNK3QhwRt7rfSO29PzItNmLszW8PTfav0p76yc7LN9SVx0e3GwZ
itY+sP0KSnqtX3qNMBkBaAUOIy9M7ARLcpEnhtiKKTBlAZOeL4yupcP+U5zbmHwF
Oxs2fYhmtYdH7bHvZfdh17HPFzK3H4MMuJGBqBXNSgG2F2F6JaMwhCZXfiFDypZE
oLm9n7Wp3Se0pHgoy+YMBKkATu+CygVS8AZGeliHvQXfKRhkNRR6O/PaQvvn1vaO
faWQz5x1zbSQHtXOf+9mnRZUYcEOb6WCc8mP6lxZ4gfXDRUa+qdjrZ4dGeUuOhVH
vyiNr6p0+8KSlHKmaXB/Dez4wVtQPAs38gs7Z0agT3G0j8YOTQCpQmN+6VHDbCT8
`protect END_PROTECTED
