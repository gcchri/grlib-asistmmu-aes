`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xdLpyxjBtFwkoCDBuC1vPTUAFMviKMLdlO7k7ztnZXEGwoLlFVSg6yuFU148YLK
jVozvSwqvMjVbs2B6brU9eipt3TcecU7u7OV7a0seU8pBKlNcEmUgKF671ajbTmn
ST7eBqIC3RdwepyoA3+l6vdAVL3zJ9iqsRetwCuC/qu0PLbdK7n9nCasCcLX+WtB
Jo5ZE9ORj2RKhxcIx9vX4Rh9M5CyJCgCkcYw2QTvPTv1VRuy5fwxVkZqamQxO1Gl
mt4Q9R6d0b88P6vW7aDShcFTQACDq8H7ySD6hhCBcwa5hW3iLq+IJJ4b9NE14XcB
kzLUR9ljduyglJSUqMG4lEcphpILgw2zTEPVV8Mcyz5bHIGGoTcmo/NGJGBLSURW
QJ/uvWz4LFwzRUfQDn7JmTj5Dr44IAmodQnqA9p87/NoJEPqRIFF4gi0lLLSfCi3
dnrctbSFuXqYA2el0iDzJZCFdODkuNU//mwuLBb0zNime/FAat5LZuXnnGjvI8yo
2B7v6nU7n2rrYtAKgBPueUcN7ljXrp5ySoZn/ycNyQ0oxCFA+As+HW8K0RwjTL96
kaHgPwLh+GNlJx1MPRSmt+bt0zk0A2JWVt1S1TaXsq+1MdAjzICew+mYG6alovpg
+pjkLCk3frqjXUEO3aFlnBnGHHCyhiAB9TKa1VLy/K8QmojBqMTGakanmEsyAQOv
ucBoOpcN0cI/xCfwl9TFYgw19e2I0Pk9nTUDT20IHB3AyeQjND0w8HymxHYkStwx
o+lHEKMi58BfR5939JoYSp2SSTDXvZGuD0Lmjb/j+/dbheWaK8NseS1/jWD8CRFB
CbRUMFaBLKQIk+YwKUYdqxS7Pi1Wc0Hd4NwZYLYcAYbiemvG4TkgOf4APm5GbB19
GHe4tf26ZCozQqQza7+XJC+NptSz6G21v6cNeFhthSGEm9ATzeiOjX0dPqEYoWCF
2RGD3xOWx3sySgrpnLuN88DzNqmwhAm+XnmXFu/++GRNckUyke8Br48/NzlNifIQ
BWZkGbNkC3c7GBypXCHiBSwVnEkeqjlUS7c4QQNANPicA9ACF3JZ7puvbzF0ewgs
3bhhv6rrpdI4Acb9LUe3qr1+LlWa3XlIojUYzSh7KIf3k+sOtKfsS0i+Ye4yPzEz
D/BUYSb/F5sPq1TOYeqJqTHsw7Z8wVPXeh9DYAG8wLf/kVBOBIS+8qQox0CnbFAR
R1T5O08ez2dxQUZss5EItIpUuI7lNIFHWUrMneRzPsckOyuPIUKtLJ4cLJKwmWNW
76gvQKJ98DPzcu5XeBJkrcAZINE4elhvKKQyCFAhwnk6uSCQtFC0HXEUm02FUNx2
JEUn+1t0xB5yBL35/lnyRMaIkobm2ek02EHyo2mvD2gZeaMtJIxbEwp2PFscpxKS
NzBsAM5aBcZdS9Gxm2/8o2tc7CS9F224HY/KePA11KqFiAa1zz583b3w7hivagqi
ndfr4hqPB1Uty5fdDhXE3ovA4BQfVjykxtTHMLFavz/EHco/Z/46xKmtLTPPP/4O
4r7DBgH4sddCq+3ynGf6VANP7bYTb1h0KmZMzSG+eWv692W/TGsb1l5gGjHg86xc
pAO4Ivj76yZd4pofKK9+H/rEGLE8TqG7CFPRun+2ZAU4vrfe+M34b3ByiLI1wvey
5QXzHKBFxPIiMP3iNxGb9PL5SY4EwICo+j/6ZZ+ogCIMYejUeIOc5XvP8mjfgDpt
KjJXuSydYeEbR/bdJ4bmdwsXx/r1lvFM3Zyi2ib9CPTBWooPO1AQ7/gbggv5cJiq
fXq04aCsmtQBwnWUYNqtHFP+1LBuBvhLOJdv37/4mHxzRGtO4q9BcsFevHyM1WaT
XA0TSB1WnEuZoxsGQMhwr4c1aCctRhEo5SpmUSp5uJC3RQ/KdMT8n/Grf143PbpS
Z+2IIuS4lkTJs3ohluzJrApYmutbYZpxpYVvkJjnQVT+y9rAQUUdBhHBwuG3jBEK
DjsD0YkgJykD1HkZaqOPUPv0kvWjinOrzCcjDeA0ySmDXnehepwIVpKuNLAQv0ZO
HaCQGNE+K+/02pE8L4LF8kqG6ba6+01ZvflfIEDXcVysPCWfmpg8NQ0lyrWDYpW6
egCROKJhvUn+DoHrctzQyHfsrTchNxcOnVxO9AskykNwRNMfH0r2DH8rGRD2BhlX
zO3qQI+nmBUqWlJCogB7S9vasqUgEJt145eodKdJ+LasOITBIXq9vl1u6/RwySyp
hVwHb+pc61JfQ3iEN/2t8PC5MjXOlJ8kXKHRW0DaDeeyES528Bk1wKoyV5imLqXL
1Trl8RXsbOvLxqkjTS8CmwcqpwXr7Q8DJYVyqAGS8vH1wn0lWZJnrHkAnMiQMUrR
ATxI6mFvsdVgHVX8m0idEUjkTNryixVQ2zcHdN12XRarh9nku8t6ehu2kdKXdTrr
gJGNmzR8UokfdoMf1lojoTl/XPv8pHxy3xmC3AjsPZT2LKZk4ZicvOwDzaXHLk4q
bm1Ij1ABt2cWedNC4CRmuU05x+59yXXgtum+VEp7oaVpUN5Usoydn3JdQdMfJO3Q
Jm3xbisx/1k5K3hIzdEZ0MVSZn96kFz1RUcWEsNhBwCzUqRZ3fuZci6s3LPcVGYH
0uT8St6NtRm2jTf1NatSqIMeNVcRFcmc/jO9/Ky4JOv9TUImvLdt+InqozvXr4J+
RiCUNcwzbKudmLx6XZOoW2T7LZj79zFrDAhbkXoPQ4LQLk4rdasA/bD7WAtriB/6
gno1xdhJsMcoNs+wbg/ldwaPHy+TJAl+Rb8VlK/msG6jiohGL8WzNK2w+V8RCvLt
hWV0hSWBg7udQXAOosUmToLbFERGXAgyT3hZXDtsa2CjBGA2ZDGF6zK8sbMhhb+m
1UFndUPd4PQrU0jhy/aMP8tKq1ul7wRVnB8FukbGhWD+IKoRsY+lND4YTp7EZqTK
JdoMNqjkQzYqgEOQIOGfGKCdlu1/jXiEy2Ooa/3M3zAhS3WAPdMDCE811kPvBqgT
SOGbosBs7m/a4OU4lzIxgrntymxfZ36ClU5HzTnfJnS+9pSQjzs7Fvub3/alcQRW
jNKGgtakzwlbEJ6VRv++OBDiXAcqeS39pVd78+Hn0AVEadrUR3gyWZp62+zhg8T7
GT7RDKb360K/SLAQPc/g4RzltlwC/gZOYnrb+QdzP9o=
`protect END_PROTECTED
