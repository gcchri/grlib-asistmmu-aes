`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qpVb0FN470KPhEgsgoHZ3LjMmu94b+xRPxs0N58DuAWQHv+PFGjMeP7wV/lhwjn
J3DJWbSWssqM+ax4hBHMXfD8lBt1rpbmLIQAgA5OeUYjESw5pfzkYKAlnzd7daGN
mRNuyzpbPkCU/7jVp4m0g52XqA+wNZ4HkhPcfaJI99jrILFELyrA/8a2bUvMx/7i
MPhQxvaJ78wzbP04liGT5lG0d/GmUfglE9gqJuhcNFrRu1uHlvPAk/nWWaONxFxr
z7/Q4AoDbpmOJbqxmo2quW+0oaqbeRcfBZEfxXFRTke/CpIbTcdCcPNLVXADAkgv
36icgN8AtX9F5OzJAWd8y2LHb/vnyU1sYkNf1M6GGcUBr1LC68HJ63U2NEvv3xy1
9RHt6m4Y6wYviUzTpeSZntJqYI+Oy13ox/ADT40BSIqKrsUi7/QrfP0YeEfScOoH
0FKJhrMyld7MYp+H3fLqvA9VkSd1EqVNVIhcu20sovsOfQ10Xr5EsV3veblLG14p
/RAPU4oCklfkxyM1OlfTPEyV1U+F0fC1zM24IJT2G3shJL/YteqY3CQwlI/b0mj9
T0QV+1XJ+B47jKM6txlzBxYNrpdJ6VsFhnLfIJjRReiP7CcFa1t2Wbdo4OBa+8Lj
YcIiboii6uRKVPdKuB0uCWqX8FPP+4ML5TbOqnZ/D3xpjl9Jp4vZPOA/KQQ9sWUt
QPPZZ63o/2b1JdS3FtAfZtOvVI61FF79E5WCySQDpNwGH4dXnFSm4dNgv4CxidFe
n/+XmmTJbGXcBgBYynGkswUj7K3K0fU4dY5Np/7gQe0aLxdovEOdLjtEerQJ7FT0
qccyVPIYSVWlMR7ae68A9iN56/x+rw+KlbROLl8dDF7RPzXOhfsyKUZi+tGObnx1
vTdXwxhQCwYWZGekr7jY1Qu43KfqQE4gRkmIR8SlsBTlbN8cA/igfPm740LcOFQY
QkLoRPZLTiQUI3MfhVwR6EnXjfrTuP9PcMx7B4uuovU1zuhBv40bIjW1wrJ5jrMA
/vR4YEG8YCh61HOLDLbKytgnhZqdsl5xy0VR+rKliK1k1A+88MqEfPz0L2e4U2el
aErJUdrrW8UUDrCY0ujq37kR2aWiqwhrqSYILaG+z0Cd6mboF4IZhutWqdn8XfiI
nMzQJefz2UkaDJ3ugTpxBD6BkNytg2+jK45ZAblbLekc9A9GUpmVrHoKdke6yJyU
7Qss/++fsA054prbXgBNiNFLAcgBzSLgElQNwR9mJVmGMneh8Ub2zIEuoAWlv++9
9H9R8Etosu1Uu3Z4QKuUj48DahYv8voDIJWfxptKVsFfe8W4XBysGsplwNpWniK/
zosxXLzoAWJBP+3wHqos4haxXMJ6/dvPm7DZSPvtFXdC4PeRi3KQXOvlm3cIvpkJ
k3bbh4gJs9xVkYPJgmfV/TRFc92hPZBlAxsKwSdsBW1MClhzoUaxBxNIdaXyCFSw
MTe875BbSY31Pa6yuaYx2QUGMrQIiYMvQB0cylmh+qrWIldjHNG1lEqMbmvV9aLp
wEaRKKcYgh9sbkgJj+u0qt6tnwKQTwe7F1fP+Kyf3qRVyvLRXRG0VOb6amAV/bJh
VNlvTvFIXxmQkMieYpJGWNJVseLlssv8pwJoGu/IgY7u+pqu6iytPPkRlpDM9sCJ
wyfADcSXKO6O4XllKqOl88z+XBw43oU41Gbgf0JIgCbjBb2GCaza8aNugjI+9liR
rKVx3b1rFenompmHgRGLf9zMEyt+XMIWfhns61j8AvtcwY/xL1LZdJ/1rYn7TUni
iad+EBGzAXoZWHEfpIwstG/NUePbc9uBGgLqWlgKroAF5dSUq8FFlIBylRfJXJSG
LkDe/V+W8bZlJh9vw4VZMCAFFqFwokIDvu2SE/md2a1zr9dd8VB5j8DuFTjlvyQF
VYl3iTDHsnP1fQM3+rjyr/Xiv8ISohe/2InPmPittYTeT4fi1NnTpdElivUx+xxq
uD70uRjqM0TSADACQ3LJcQSUNoKV9q7Fes3rT1rl5TDeY1PrzvijQI3R+Swpcpg5
fedtOwCX90to2Vq3C+MbUdZDgh447CBwI3VR7g71f+UMRRM3NJGU0oePSTT6oOiF
Z6IPgKnVwuaVRctZRsOXY7NUD6Zk9uuQ3H8xPUa011VW4F/QNNzaDQyQlHgEcD6a
V0WU2X8KIBZMyuqPwo7tYyBnmA0wcRmzdWLm5nypBhzGW7OMqosDNsq71aGRQQjM
Fq27vnYi6vUbhYcAz5Xw0YKeqUBwUfjVaLhzhZGj2XPztDN06f+fkQ9mKBFTX0f7
MGbgwaiKrGC9uFG/b+joSEs2EkmQzBM5zN++56lb89W+Yjpmmern1nEzgK8GYDcN
9WugDIRtbL6XuDvqqUvEpzc/oB91cVoOaIxkN7FPbh/slUDA40uyrsBcTVTNIwic
K+mLl4IM+tcG7JurTqiZrVIbcKzpMqQgcs5q6zVopM6YzJ0jmApBFCRAqHT+5eEw
lnhC6CbEbj/7xfhn/qOH7tB3boZ29tXEkZPAO4I1gzMSxyejMycWkBpMlTE/uM7N
3VBayDK/aKr0LVL/9yL3M46769RkxIEmusOdhEQjAnNuqaXzB+bxw5A7B2pVzWzu
uwD9jfXGDwHG3ya7khalrn+RtDFTrc02+G+hNVWurInj3uht+1gBHaG7JyiZ9hGm
M+cfYMasEX+kQUkHhH5SAfiLBQ3dzDMS8GRJEOfxOVqzHfEPAtQRT9d0i2HxSGYz
t/j0Mbl2Es22+SUOLxu9CiSHB0ooISPxNwceht/uenhy8fItoo5UiPOVno7rgltC
9B9Qn9rahacGbGicuJiYuQoZwyVyBSzeInfPMD7Is/E3FrQo9s1Dnaxr5L0C0EJn
+zCIK0EfYNb3xKxLOSPQgyGysD2QWPzMsF7Po2FN2ATmvMZFPTr61e5i38E2l7XL
ZXGawTIo+v5WAjL7cUBp9RU9UpZhuuAwU3QdLiYrRUSMx3fhAIKSFQF/IIc4liHM
v2O0ISFa9JL+RV12DNjVWdKPNGO3p7/RkNk+D2ei8Xrau21yDKPEPNgzTG6h+ioV
x2gSNp9L3iqPMgUDBT6CQQ6Y/gaoBl/rYN1/OF/gyuq3GhumTl30LxIPivhU4WYT
zqcOieRoPTEKvH/N0+r/XcOdmvCvF98cdJLt/PpoPKI27pcA1MIGL2jUcf08mHsI
/3dDeCuQaOAtBm/B7APs9Fpa0Y7HIOPpPNBvcualQwyR3q/Yv5t2mfF2dqE3r4gu
AjDCwvRB5CZ7whoy9+rl/QO2uHm8nV9BDPSTmGxbKOZFKUQmJWqWPu60UiuaTzlD
AioYeO7RVsJQ4qQ9WJEIRs7idak88T0quYGvPtZWxtJm4+mqLLK4nRL0qUPb39pK
AqbIS1rpizWPVytRiWGi2Xq0cVQQwe8e9uSY82MZZyFT4BNXjJGQS7luDPl+4LtB
RvGmPYBXX3ya9V0bD6twJOW2Et4GBm69qaJLuH6UNjQLN7N6r+m+d8q03pUH8Dsr
mEUmmuG5CLE92g+7H9RaXoxKo1P0tT4L79OQ8IIGGnNrT9okZ8mSrXwcpw3Z/80k
OJACz+f81RqMBkOmThImzkk5GMMvpebrjdJ8gbVZ4X+4ShEqoTFvFhHqnPg8+kc3
NRT9I7inxvdZw5IfY3U7FN8PJZOCEDQsRP7rD/OJo/+nZvKhIIB0WIN9BXtZVyAf
w8Q8e4PPAUINZnnjjfIi4QpfQxL8kyCx2peejCLcd8Pm2nqlleIla9E0fxhRTcHI
FkcaYB4x7uySUSoSQ53KRijgpHNyzosT33ks+1YDdRYRDmkSOTr2Y+2sw7Nz4UMT
Nes2IO8auZfyQt8WwagCYDmYfZnGLUAaUqTLvjvGmucmAq/iFnofHQTCsxi115a5
naquctLtdRHYIH8yDgMcB0Nh04fLVAgQcIF6r0A/wsfGVBYrkdOqULkXhGXDlaPJ
G5+CsICXXpWEFvfQmkk/9jKIXLljPoNsWLmtGryEoUveAmy1idTXw38yWGcEQity
bp14ECPJF341mnp5HQQ10n3Q/AtLt7TmUKbvz3umFq4V/YSjj7TytQxPJd/i+ylv
GZzP1e9xXaXi+65zh5XoFQss6ohs1WSWE0uO9een+WaJzkkC/1a87ALURzUtlU8q
bR3goVZpjZW9LJVRzueM4GUjZq83hyt6hwhdfjy1eVkzcLHZSLHfqjwC+7LMmRzE
AtuN/JS2p60EUke2pexd7mGJO4OfkV6vxWuVOkVkuIdaGMNqlb8fSSUbpxT4+I0g
TFk6urZ1JBpGdYIEWERkJcV0vZ9RH0Ms4AyL6Ftf1FuqcV7X+NodfeHfdD3fe1bt
Bq5ZtganLceV4USQJtb185v0BSk5lYGfUscGvH/dU7WdvIDxQs2oxeGvkrvdo20Y
ZtETKee7uv11CDjCVWXWNi4saReznH5RvhyVuasRGWr3PDDitP5CUwnVsasvX6GQ
FP6x3eYb/1/dAop2Q8PgJFP58Pk8WKy3ThHDC2TO3WIbKBWsFwOmngUcbOFkBYKr
CGw+s6lmOeEGA2ppZD+cT7gIg/ZbLL5quDTsfZWFEUEUo52dvzQzG8TcH8rWbD4F
9Ad4lKbOXZAmzxqyhUN9FIO8EtINRXY5khSjGp/5d0qyvrvcmhyKCwnQI8gmqjvm
ICdFuJCvQtyIJMqGX8kgPyJFalnh3hEYFXCOkdw5rjri0arKwTh9uMqZEFmUuF0H
OfN5vsq/pz5b+lhQZSAKkOCqXXCMC9EbB4CIt0d7U7ol91Xg7mhdXPEIJhfXYYbC
2Uh9jnKB9RWu3R64QQun9KxkyNp4aJ0GoeuWy//PRc5E+6Dmz1cw0N3nPz7l4w6H
VQX3j6d6uSpMX3GcoAnqUk0hKlBnu5ho24c1kW5hDmLl8uaAFgFJQ52oN0Vt7m8s
CRIjoV40ZI9+1YUrPIr88LhMm5DUo3Y1vNRuaAqCKIwN1jGh49c3mpG1QT3x8/h4
vTliFnyqRG5SHliuOKDNUg==
`protect END_PROTECTED
