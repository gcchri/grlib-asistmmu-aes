`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gW7aWXkXHqZWE1G5RtJWB4h0tsVjfUPfgaNW/h/GrFSUI54JvpcZPzVs1QZxFvJd
rsj46sfWQdvmQr3klujImdoTLPAJ1VUWF/J7ekzKkHkU1VW08K2EMJtW/DLc4G1a
5RxU/+enNKR+7U8+haWBF1IlHTxkkKXbwyeLDi62beD8f/AR1C9qOCiiUF38Z3g2
nt3tUyOdEeVpyFioRqIo9xPFeSAeM7TGzoGITWM7p9in5v4sCd83w49KQXLoWlbk
yJ0WnWWa4uq4x0O3cZuIuv7QogdNKxx6kMmrLceF4HgvVbPBe6oHoUvsv0ER9I+n
Ki+mbXLAClVg+iXK3KmZm0rPR5lS3rF0BhVu2CmTRhm5hJPIwaCAc6PiT7nxyFFi
sECE/zL8OAPvO8YKf+rEq9Q1oU2wMFubvsWnfexRWuMlbN+khcZTXX+irVMdAGaq
YrHgcR4lVYz0OtWx47tiiNJAK5C5lh79D8RwaUYq5bGM1BajY5lY/ZguPL8zelhB
HlFQUB9x4plI/PkAJNhVSq8ivZ2KUKn7s4Syq5X9eY6WtFHkjB5besBd9hxU3JnB
Ju+1v7qeg/YEUYg2hcpvJ3G+VJmUIXP08Ir6JDiDZVxgzssSHFjS8UQX4r92UgX0
Ur5Cxdx/8aRj3YExknyLFLp732y4bX8/eo2tNVVLNzpa4z4C6sLmP3l3pdDuVZ3Z
B06OeFXisG2TmjRM8Q3kDkijvURUrIy67zFSbFIiQyOvuKGw6Fm/C/pupktLvG3/
8KXdJR9vLerIFSgANPkibL+D3r3lENb6XDA6YHremJaWAhKuXZlElIlDCxcW7YyQ
QZ3b4//BwBL5GsQ9SyrJ/KjnQ2ktaOiGFdN7+SEizGJFlXMCbMOJfMSV9WwbsAxU
WWgjy8GspCkCKOKT6Hmqrsj7iDP3rtMgTUMWHf8aNGXQx8ijfK8oLy8wndX4nKKG
`protect END_PROTECTED
