`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j/jLBFkwGeIzLnir35mtlsa6Vv6piaO9c07ArenMW3ka0C57dtXpAKCPGlAiytEW
W/QPlZuj/bK41T40ba43Z5F/HA6CNTKVxGBeRfxl8VTUlTrfRnD3rX/YU/JeuVEJ
myyt/UVtyQROEICT/UhJHFmW3uxzSrzfmLWu0eTO1SH6tzhGHO2ccAGa0Ae8VXr1
ZEZq02Doje5swCucUcIAs3qIJFcZy0aNWE7UJg/NwWUSzvhCPlR9e9hvCjtN/Shs
9aaoTkhZddPXr3V5ccOmJ+YHUAIZUnnLAsyjgcbdQKz5+X6FwQzlxfyAQUR9hvNB
0IEirL/uFg5zhYYNUhD3Ar2bDO2gzBBa0LWImgnVdJ7o+sfwskMVRof8W1oApuwr
UoUw+jeWj2dij8xuGuByRA==
`protect END_PROTECTED
