`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5RQwD0RaxYc/Nh8I4dQyhH/hv6p0Sk9zVWiqI1Y1fE2siIH+zdGkY9iN0kvx/vx
ZcaRP2BYcHSzi+ZbJk2SO741ftLs4MqFmo6v6jpC+N3O5krRsW9EmL5m/02AsleQ
9tzSBdX8nyyQjAybQWzYNk/TYzoUc/1BaBJL4iD8J1XyYq2T79qpO3/ZiLM7PjsO
EA4kxm2u2M3rm/VpptChRl3ks0MULw6K7lKhf3dBbyZB5YJf6ic+vzGgD3VySVJO
45BQ9nqeNebnJO4xUJVISkydCFGHS8KCXPEL6alZ1vZPwImVxAxMGwGDH5c/g5vu
+57YRTds4IU92omZ6qfcOvTyG2Vsoo8L6+MQaWPKau4PeUcuJ9j4/oa7RbBhJVoc
EgZJjovgjpfsDrYa6R1hPB66YGW4FI1MovTy+qjAi2cBpoOCWO1kMlQ2AXjmalDs
+CzjlsVg7gWT3rpfuiYWMHnqVoeLO2ENhzk2GYdL8iHgBJRo35I8OqC1utEyTdtM
AUrNZV73hqAM9wS8s8e9kajRecpmJXrUflmoICJVKy38vSoyCNwYDXlxVIG5n041
bgM6GePX9ihYSduuJ4m4HS333P1s4i5RYbsRoze/JF1RVMJ+m3VfVtPKNQPZF/NR
hb9CVVxWT5m+t9ezqBUPe4NqSa3frZ1V69T9tdoXSvxo6pA9+8sXSs6GHmqtctsD
JkZMLuoJ8K5vpnTgaZ7d0+15cedHIqnr1HR2JKZ/nAF6idLqhbaoClV5CGiS565V
SjjNF7x71cgWORmSSCci8LWpvOjnsmU2zMet93DBbWvW6LNy6nrgpwYCBVBNUloh
ONYb2J2laWNhCYpSWOXZaEEKz+bDGng07jrPw8L20BfnHM5KadOE7TJgFwXWFJ0L
NPW6SCp23fjFNVGIemT6AJyUySRE7stU28v1crJvaxTXd/LIMbQYdHARrjRnCCoA
ejOc8lnr87bT11MnTudIK3guuO8bLosXSjIFjtGQqoAFlZnKiRtR7/aA3BvWYYpS
ZdebBndI/F6xkLFanWjITWLcE6VcxJHjUja/mMwB4u2nITlEP6V5ITI43KkBy9Ex
klFKVsnp/DQqrLl6l0RwNRPOBJb6KTW1mi6gro1jY5A=
`protect END_PROTECTED
