`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AgjqW1c0FCNTKpL2PA0SSxfuHBQuh/+7g3PvmtcF8vPpWf73tkIZGTvdOHHtjW12
egHshsnJSylBecyZ55BRuH0JqqZF9/WLASGMkSK4K5nWuHsQp1NImAfqNujfDe3s
Rvs8Y08q20iGteBs3zUQ3so/Bzi3AczbOoF6zEDMx0/hQIwaWaz3DDgIzSfVGbUM
At6l5X4Ng4OTy2PnbpJoeBr/fOdbxVNvr9boDeAN0oEziBVOSfVcFf/G+vhH+3Sg
wHYpX20++mPmG2DlzN2NdfepPxnN0ofZH4NtNrcBjgv1Hzqdk6NkcM0nEZD/YeqI
+AUEfbsHNXEJwP7FG/mSAhxryET4EF2bS4XmO2jmWVHCkokhQkpOXjuo4XhHTLmI
P8aJwmJC4p3Q+rcqYv93nAWEA4xNMg8S3iNOUM48+MK5GZkh0NJA0PQLg28yplVu
QD5S6k8hJ9MvCnmxIN8eC0GO3Ofy4fHw8CXACHgCRNynGPRfxIJOA8UYVZzif/XE
oFqn43E2VbVB3I4Rk/Y6iLKCc0niFTw8D9P5bS44CvzMiDzchVEiCspypkTEG8v0
OL4QMdZTnigeuMrEnZz4AS3wGEPpq2R34neSSFOobcWcbKS/hc9LBJoZaG0UAL7X
8UtGc77s0M7D7jKOFRY4Srwxw53lm+DBGu7IvKYxh8MmpxlV75z7P4KRAUKYC9y8
PjEW14s1nTALwpcgHCSQZ/A5sGC8Tf9Z5USguzGcfhgSddHkBbtSDvW7XW6ubxH8
`protect END_PROTECTED
