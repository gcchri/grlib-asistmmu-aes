`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+3/Ik/yLmZyMmaiB1CB5aN6pZ2WJtv0XinfDNkYevfQkAcKtYTMxnCjFITI76he
W6lJoN6spkvUYe8L2r/6NGSZ3t665FR4XMvtg+Ult3Xf2dc6nyBu+lk9uT1msUqe
M1pxPRMQOYXqr23tqQ+AvG9yG9bqi6khrtvROhKVYJ20MBnHiV/60YM7IdxYGeQv
RTFL9szjoDptnl5/AyRGYtyYzy49aKnAP5drYI9Y091aTWuD9MEaCLnBjU3j+1fk
WklOQCljYTvJDYjjfOQHfQ==
`protect END_PROTECTED
