`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2N51Fic3fgq1J6TYQ7gr6qdxeQOVv4JlPfMPzjZ+Hc8wPew5ootEs4VE4HrFS17
jX+FiitN1llf+BqVPyL6p0+gHvrKvUOTyg714X9opPwrHZMidfMDm32EUxDD/PMY
cyM0NsoNUtvFCZa7STJ3+1PS23Y1Tm9Hf4lHZF1bxKGpEhbDrhnIV1Gaf61ZVCDu
+S7hvEhzNF2d8lHPYcFhyhJT1qMZhorlP2wtyjXfDCWQV05j9vmSkS/EOwbFDo6/
DNJY5A7HQymGufmHXpfS3zF44vzKJMDoYHbfv3+tVzKtTlGPzE9bVen9NSu4W7WN
48nqDrHILnuxqviABP0xonBi2e0Bs2pbmy/EeuUgsJzeBVGMYBmX5XdssJtKpRpW
fn3DtJ9C7JBxe7DiadysDwtBBhmlrElmCjn3h6wgQDK7xaJlYym6D+c6A02uxhMe
KWzYeYxDA3+cHUDJ6lKXImsgbHmJFtHngfD8bFGV+feIHx8Eu0UJdMwGEyBC+twe
43WjN11Join1LPVIwcmTP4AzRYSuk8zNbn+If4ORGQjawbMitbWXTPMS7cfHO7HH
iDpfDxV1PgahBu1oViezPYtZAUOqIV3pLdEKIwa4UGH/4Hlv/sZCGW23tVknL0JX
Upoq7Lt89OAyqPkOGMNJCDfKGea0S81F1LkkLP+7/Z1k6lKGKkR/COjnOti79Xui
HBuEW3AcOZ9Ni85W8GLlJfiCbfvfDA88Ei9MLVXm4GFi4Z7MfgUEdg0F1EjMUxnD
V16KF0Ol6CbbRWva9361ccprvgywxAw0W3WtNvIJb+HGofiyAlwaMDHRRVwbpOvc
bqehJTELvLS3ZSRjabMl0E1wD8tKvGYZQ/ec5UhfvOeNzJT7XW3M2qNCPJlS0SbM
3Uw2PIGmZw6h+Sub30B5dEJwMzR1CKQrNFtEcF/njB6xhY3b4NmM/5HvN4OtH8lX
A6E3gGE3w9SZ2T+oJHlbWkh3aqRhudzSCLvroiELg1wWEKXjfvgJW9ZEfqP5tPD1
96+43nzlBLHmTWx2rBDagcZLOPr8RpKJkbz8+fFAHvH+NBXa/p/Z2p/zV71mF/JY
O28E0+lqjguSB3ckWnZYMIP0N0VUrLKi7ah6SyERtfFMkZz7QF3/F+oGPvJ02dH0
0IzG7+Ecmam8gPi8M4fg3A==
`protect END_PROTECTED
