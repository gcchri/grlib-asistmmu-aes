`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mMxfi2I8UAv1CEMzK19AcwuqntdS436LOzh19rqMNWXyYzSxMQoKUrxM9gUAaW70
XAJA5+PkLYDfIoLRhOGxMFTw3hPuOnJVMDjRyvzTnlw8dB7P89dlLFBsQgtAteBv
Eowh4mbUqNCL9nc7anEsecYxDNTsO39mi8zwypLRbAAdJQ5kUsvDIjbhmOUi4N09
/gdQiqnqztdeanSQA8M8Ryj6QqtmgOIHg2VE/2X+KyLU8PKfDV5CkiHLZwE4Yb7v
fQR475Vh72vqvO2AapdnS1QALCfKnre+wyu7islrmS63joHPlaaaWaj28LdrmaJL
zo5W2W/EWzAAyuk3LEpdD0odbzsIGAPmGtLX9uuiHbu9DzktDhPywSwQnTLE2Otr
CLrxaq6Lr8q7WPioE0+1+w==
`protect END_PROTECTED
