`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/m0yIc3IBwsA8cvHOK3ykOBUBaj3Z+UHJd688abnFppNTZwzlRXVVZYOlylMLf5
yeMpVQd6itdFQ0/tYkXTQJM8q9gy2p7qIeFJbYa+gopVdBQr5UNu/vkFEnBnRqLS
BpKHTOvnQ/c96w6MgV77P/TbIP3zhZ8pLaw1BPkbqR5jFSJA6L/eLl+gblYuGMai
CN7YX8Ea0RaYvtVczYLBFQtMavmRhGx4M5rKGLZZBlLkbVb0R2lfPW+J/IE3rrkI
WPAUijDhuPqaQmLq5JepSJ0eIHD2Wk7n1g8DGi1hNL0xFVvfi1LJlafCp7Bv3AHK
+JEEmlzq88BldH1dlL/AgCNidS6aP0XVLG4ymlJV0sc8Y4+HuH5vc2htzIOVdxmC
jQFPvdoF53+4OPWGIUWma+sQJaEVT4r74eRAupGYXqNDENhN3C1246suE/vyrMKo
YBktmEyVWKf5cDrrVsZlBvtrSM/RXndAUbAUmg1gCrpSHo6aI9y9V96hP7Klvas0
G13dimFZL4vB97KF+MZRNDTE3Cc7yr7WoVCLN/MX6RW9M0EKCtogVzlojLvTPaWD
mJLIP50G2/aAvNHjva7BZIALpLP5Us3/8hCBuwETZGRbxdUjoDrlolpJ+IosQZlL
3GJbnJViKGriI0yFF2YCIRsxmWJNAN3KtGJKk2KgtnxD7Q3ueVnrjKlriWzLN8aY
jFqUfM5eyRSKbkmXg/TRRmndVbex6BFaq0AiExmC6js=
`protect END_PROTECTED
