`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
23Z4L6dJeU4aGMIbpFfHaKTfikbYHJUP5KJOHBC+R0HRU2JsHdjDRi0voekIrpIS
46M5feJ6QHD8gOwDM0KOFrSG3juQP0lU/lKkZ4kK/6zzAAgZInL+Yj/EpJcGf3gN
J2mfeAIOFl0cuvmP/KRgQcw4/dCXndwlgw+jw1ql0685y122eTFJQXR6cwmKh08U
rxZaOSmVbAkgfSWHgOOXBy3OZ+juxZcx951KXNXen6xGi7raBj1uQe/Ksw3Z8Svb
0SH/S1ZTm5ewvmMyZvsNTq1WQZRpz0MbkFX2m+1NCqUTNzwSECQrXP+vnzJdanP3
a4KSdow7JWTU+5nUvp7MpLVxI+2dkvRwNac7mM29yT0KmsEL/K7VcRRI4eCQLCix
Q1Ywz9ua57uUSc4YGSBfa13B2ybbbyDOPey7X3gS5nKAYPp6Fx8mjZq4OuiWTP2L
mYg/mJZLKwmL2DUvGf5x3crfA4kjA2DBUlT3DtMOhJL7aG8PiU698VR+EFNQx/HL
zT0eeHj8moLXIbKuwWv9UeBzVKQv/f078Nh79XvyvGg=
`protect END_PROTECTED
