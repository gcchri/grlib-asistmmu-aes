`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BnNOXkanBo9RmIhnBGqjHFMZ66GvecJVZq4DnuWG9RvI1mJX08FOjOW7biJx9tlW
ROoUYG9fvtEwRBPO48z+iYMFqBoMpl7sqJDi3x23MmMqG5iuVodBS7kl7o52KvYx
x3TbvLMUBwFn8LMHPXphHsOtiFZ931n/Rxfagy5OLbtybCpARoXtpd6d0u9a2yGu
4iEHi0/CVVeo5Ot4q0ugk1jUGzJmec+fVKvN+f4eMIfQW6H/ZLf7IN1dj02CDu4/
Ubnx95Pch4cqGneDs2ZZJ3CLBs4BN6gypyhwluKiT309mNgP29cJtrcbEhcYM88T
WHFs5Oqa9awAdUpVP9dTkYbacAdWB+2Z3fwKzz7p2bFLWYkwR80Nl6K2c7oZMkZW
1rWzifGIFHPdqFYYopj3CZLvegGTthvDjc2+1k4UDko=
`protect END_PROTECTED
