`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bj/oQkyIjmrbr6x2rUhKOAE4WYMLs0Cx1hzp0OZtnVBq8TyuLmlywrsSPz161ggt
iK2GNTGAfq7h9pdRppvwe7fQRC3Vzn9FOp8xCe9LklgsUr8SPWbUtv7y7nTreZa+
URpd1Ro2fO8rwCgOWyvEhVN0O3RoQZMpVTxXISVNKrsokc2auH7sP4hjahp0x5S6
EGv773sJP/4VwQr9Pnu988o2gn3FRfOG2l1dELw2m/Niu/pj2GqqNK6fmqdRzBgC
/9zV86oZQR2Firz1EQJTzSEpsTTvXkvvARcv0srA8nKGbuFtKJTu+aGTeVs8szH5
tUMXEsLcANplUO4+cqqJtgM5cdI3+aK5ZhNFNEAb0pwFGTGsEpW/8VhkpV3slKIy
CdWEFfY0W8KKkkoFzFEzRMRpQR1yQjFAlrx8or5nj1G1aRqTXhoyg9f/6Ewqj/so
Plmb7M/QuOHsA5uvpBc9RTdDgdkZE2t50fhSZlDsxXP+6zfX3E3TIPKP3reTYEJF
x//yHawKQjfwq4it6xj6CC8INPIfudExFKJbQilp0g1iW61eLwR7RvsKcTjMLoeJ
iodPzNq0SdQpFlLQQFnXDpA+5ob8bPp48WbBEgTYOm6uiKQ9VJHRlR/AIJgtbyLf
njKWL9MqHwWVNrgnXfgRIIxV09GIba7zxlo6PtfHlI1MZU5Fcpy+sRHo6wmHJaJl
WfVA+gSga5v7Y8ZTq8aZFxrjIO8101QrNhIU2Hg6kIEVNqHs/Srg60jNb7JiS+w1
6w1GlbJANzaFMS3VlWDBWzTdh87scfv8b/f5f5YLZ92fTGGFhES0RUEK2ZHynyGx
QsuGE6nqTHTxz83+flS7V0pRfEmHgAftEHvIvnWg2ips12/KiSABtxLILpPo4hML
gKOFdizVls9+bRcrspdXz1o0MWVcz/vaabTlMvDjyYeQhcqJCkfSmPvyMGuiy6v2
DU6xS/aSYoGd/XIChtMB/zns7cbtnkO20QBROeZN5s2D9+Vt++8YEuwyoSQBiyi3
QRRlkWVo9nll59tmIwsM6lLhvvxf938q1Ft5+AL7AT65X4obQqJYm88DZiG6FeZL
Avtblm1SEr9aQFBZ+r3tnh0ZlUVkRXjWEvkayEQLwCs=
`protect END_PROTECTED
