`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1t+ru87D7TvCM7UraaUSehE9I9NbKyCQm8v3MuaafwVLVok3ELJ0tVKpNAig1zQb
Rjzb4Cd4L2q7rKViABKpdGXxt8BAmd7JqsETi4fZ9xi0yvgcccWzzeIdx7735Vhj
Pwi8LRSQVuwWR6xsDZRVzpvu0i7exwX5N7cjKLmA2QXKBecU2WxwRvBZ2hNIA2YT
bj51jX9JbEDsMVQjSeUYTZJS3xo4PdA44cmDhCmDHF5kk78QtAVZN2rhL8moo+/Q
yBqQkOJVo8BYuZf2uq0/OLJ6b/y656GdG6MfVkcOVXmWVXN8ZU6IE9R4cuG4c25v
4r8p6xp4rr12k1Q2pznKZGRnuh1da3MD0EywbPDSm/EgbdeL2FidEW5JvgitWhf6
AKtX3c3ffD8lJKFo11KtHZmiAvXdj8XyC2r7Ps9E5SxYU+DiwYF4LWbdeyc7s/My
uQ4ZSzLZzxPmm5qGY9WQOw==
`protect END_PROTECTED
