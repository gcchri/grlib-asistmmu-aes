`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
57Lw4JvNiKa1HXrK5P/eXzpWhVTVvIUlcwdPxFHHgWQJlZb2GQXd6Zg3o8ZXSTt+
+qmqi9vRh2nHl/Ic5fGJC+AKB5C208gRDKfd559VBdX8V4fkggGX0themorK80xz
xXulMcWYf1cz9rTi07BMz6Pk0oiIndKiMo2AQv5zI/zcoTh/Xb5nk4P/q/l+A+3y
CkL/0cfgfGWIn/W0uNJ7wOBEDE/he98Xd9h96OW7rihO82FKxh8OfMKwSp1HV338
9QFAJVVEgH0fCuq0nWNHOpxMfF9e/Ym3lxcytXpCgh0XYoQlgcLob2m3VGO2U8Zu
nOOIN/3JMvpLw2XMiSzR20B89SHCGbakHf1O/S2hFvWiXfXeCBja11t3gCX+O1js
ohDyqhS9xl07u54COo5J0B2CBCo6ZYTm2RB10c65jkY=
`protect END_PROTECTED
