`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T2Fm/wTrtVfMARg1wvPOcUf2RhnrVCU9K935n7xhSJ3AarLLx5Zr4qqDwHkKCcH0
EEALa0R9Jw8JF2crpYjI6+cQriIcJ5uO8SayBMbRnYv0dz8grHZqsjpb43ZR9PGY
IxdGuLPT5frZd6mNzyQW+2JGVPo3RgtYaxhhsGNac1B5GaYx/7gyl3KgelPc/e7v
7zhINgRcnVykEIrrn4a/B9HoQmyk3wMn0TxNux/QX5OSXDPe7QHDu7G4eX4M8rmJ
G4ZYuubF7K/IVp7uqieBEla83jEoDIxS6s1Va2iHeeDuRZXRc8lHpR7vnpQ9lpym
JSlHfeMWhJsi9sNFyvUtdA==
`protect END_PROTECTED
