`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZW87IAIfurffug4hcjsLBxXKicRQ5ayyazw2nRzJXWN/SnSf8WtrV7x+bU9gYJq
mOGI2RTyIDNaPIKG3sfHZRE23fSYAgKzBBPbg1iG4tPLb5kIhQ/drwOwt6EYQwqI
xFRLkbBlZctylw1YWW34kqorw5W5ZHMJdnjg/J2fy/YxikbAq6VCgJOTLZh9Q0uF
F13XW0B4y+zh2uer5Zk96gjvWuLoadSOL6qZ5vklMlr7pwYJDxvE7RwhtFkd3tv/
dmH80vU9HcHB8Tdil+mGeGRNXzlFnLjb1zcHu3dFVd3b/4H27u9z92JTa8Nwvr43
eMdp+0ul8MZjdsSDsO2efrABcBuXZirLKE89xUO42rSXKarRv2rLJEqHsTR5RGmT
ph1X/F69OmeIjgxLKvzD/H0XF25sDVJBefz23sqh3VYtX8MFBhF4qD9epqG/o4ze
C2jCDpiqzjHpsD/9cnCuA/Dk6LV3PXPO41meELBxLmHszZ6kTYS96mA9lrBiyoTi
KhhJkaxd79ktlj78luMONSBtSTL8G6nbKjkq3S+RjwktZkQowAy/ejoxno0lVVxt
xPk3xb7mTTC3jjHklPm7sCppFBPhCPmlyV4aW+8378w8SoVDs0IpU7SWQH+HmFpk
Fcm0E4StoYavg0p/Y5HihfKXa+p3L5bpHvISOwW371vR2diZXrhn0mvlYovSzEcm
spopP1gNNwhscc+mXo5bWJKPZWuM7XQ7RL+SHWIZf6THKmWpjxze7OMupaFr4zqp
8sHAs8WGDXWUn1skEU/shRMcjeeYLga3yl0VROVCwHpm3H9LRUDnvw+isYi64zZ5
RbtwhkrW+2p3A1sY9j1aci8tyHs/9MTjHo9Q+f45ngnV7/0vfR9CP/0b9H9yZskA
oz4brlGznz354IsQPi+HWBJ6SryuO6pjMtlgZ/pZ6Jtk8QDuTvcSjtPxpoW1WgQo
2tfcZXB2G9NNyIZrhGI3RB/hRa6kEC/fHY1sBWrNmK4zRVUZBB7oh/HvfXsOWmgw
jYnFxhHHYT88HsEBbWVWDs5fwnOzcTdpcznhpdxd3m3aB8Dw8nzSnnaV0Tc5Ywm1
zYGdjme9bWsvkVHCNbO+sob3e31vy1ghaL3A7yO8wJFaFtXXM7Yd3CYEfxJKyAF5
dVJiCKDQMyFNVxkVItpFbgW46mHapd5FcfSSM7Mc1v1aR/elXj0eOpCee2RTR+cr
vGFsnp9PAkY2ybGEDwcmvzsC1mOTG4i+peQqXzEER8weGw6ZDp1zv/yq0spkU26L
zjmkKlU+YV4zsgAF9vZ5Ajumi2QUkW6zkW5ntIm4PVMKE9ZW9UrU7O/pvC36eqdC
s//D/zukDVhe6BC3PPDAG80xiEKwaPa+i2jm/tPEvaQ9KAgjnxmxfcxmD3aer2hw
je00pBH6+JYEYGVfirgeh6ZK10/dEmWBidaIY44sXI51XsBWvLEweivCuXCmHNL9
imE/xAJ1rwvRsGDMMLHuYHlPv9AqmimRMryBV+N5n/V1Dg+MPDPbg6kHfYwsKifO
MUBWm+4oZenYDt0UHeBL5cMnU8j5fE9PWiPIHQjO8YNzsitC7f5+IJtItGYdAsAG
6pR2YeIet0q7JDU9BnhBn2emMEXV8IA+P2Mx6c8LaLY8lAEYwIjBNowDwELm1VDW
FieSN2vcJ/Rtw6sR5caEUznku2CBEcvWIlcm3GFULeXMQhrOBgBKHAfVSmyq/6b6
o4H/PhVHrl9TVeT1/R8T8DnEwBCtMqSkGEjz/89/alC0K1b4Muw+3ItrQOvtpQSG
jiJmTtrNbdGbio1qUqEqMPEVv7h7s6wAVTJyOxrvn+eXGe7p0RT5bxq0LJ2AY/Wi
ybgIXFon3POB0wc/r5J/PVybsPBXrmyL+IIKX20X9OwoFvEgD6DJvwu6MouzAsyX
gjjgsXMoryXNBMGMDYfextnfZTVq6qsVE2o+BNKhMTyER02nQX6QULixSvDzwAZO
pIRvIVfdSqCg7vQPMwsHQFLthRGdkhtmzAGM7OchjRu/aQWWoamShOOv+kARJm89
JimlWAp7pPreYo27nmQqd+1aiBYxhXjskY2pNukPDwvYFHjhLM4l/lwWjBChsdqL
RLeWJ2YhaMmiYRz+/xy950njY1PCETC20hsPgykECIPsURPU4hwczBuVGAFCo+IJ
5SnA5YDB3Yx/+foI1nzr32rTs02hEa/TNoC8Al5+XWKSjQ0SpLgoDQf2R76wGva+
EGIpd2ilzKtByfRol+z0A1l4GTvrMTACYUC+b6vE+LSe5lO2I7uHjzWPXmR1l5gu
Z+p6z5lipHXe5tX/bg3AaKSaVAJeS5Uqf8bvAHdHzQYLdp9swC2t9xWof5pz/Ws4
DenJJ/eAdtVNVutp8yLQXxJdmTpbE+VnLcOwQhWCCGIpDBXprXncDYJUfCypxlsG
+0NtOJ9qyrGz/ZXv41THaXia11GRsaazp5lXK2QTvE1niUPFj8TR8pH10o/RpTfY
euGo3LObNfcBkFFbZ7E8BID8qhSnk1AOIYiXzhd9SNGyljglGkWgutK0PF0manbV
uvAAvy5/DoKbf/TxjfThhynM8vJ5smXbbFD7TVx8wirsQ0NNaEeZ6l57wfOoEMrr
cuWsngasJXZ/HGx2TfTN6Ri7xLSnIN9yvIeTkV12r39Dts86Ij6LBBnk0XEERD3r
ehDBAZPngEVJ1aFMNeybrL6eBgd59xjCNt30ONMPhAGDrPENwknFnBGOkwQ3TQK6
xzcsVWR/DCdhxX9GLJQjAsJP7/zVk1jfCYPC5WzyqCUoRKWeH+FDTDyioRQnOSNq
eBKBNgX8zInRl1X3lbJrxWCZEch5Q7MhpSfSSSuIaRDwN44F1S9i8OTd2Ll+QdDf
MhBwO6rLqXK6JD1Wtacl5a84EVE5mqf+4wj0I0+Dq05XC/nkFaOHlMLaUEOWelAm
rcP6aKx5e008OXgCVe8eCgro+YYGlUBaQfY5kF6M/PYjZVIeHDKShK3wC6JrPpFa
0TJNPfBWbq+cuQpHMjzgRlemEYScOp/TVmAbqQtCKPPFYaCMkMP2buYMol/fAPaD
dLBUUTOxfOVhReIqi0GE+bLTPV6zms2zditTGl0IEQS559LBVV8lBrCdOQKmtoes
Pb+2M6SuH07mJFi/WCQKxRYNnphJoa7Ij9NKRPgq2Civ+Chd+omSVC6YGAf2rSA7
gRZ6MWOAVEiCtiRs9D4RPE9+qLz5ALLOZQnnFA1Lzgh30yLZc40Ujgj4RAMde7oE
S5F6q7HKyKjB55EjCzSwIeOfup9x3D+e8SWRNp9pnxMTglgLpkgcpEggHiGhQX1J
u2QJrIPu1TJQyX9pqptiyaPYFq3u998hIkp/GicAbhJyniOQBJMeFxj/vLAm/7aD
hhxwDB1uDGXeFZbQgXJuXViNm6lCyMDPuPThq0MxGfBCWNIlKEmkvehmhw0ZSJTl
nKJBTRpqCDeGe6oWRe8Mm8PLWQE//+kceD6VdTX7fYuKlMMKRsEE/mrZa55u62oX
+st6iSAv1F8JaFl2ZO01Uww7zID7DqO4raVoKE9UXvyfKk/ApEkNOe/dekQel5GL
jjK4pt6EHcelhPFg4S+jhStJGrJXGWagw9DPOSZWuk1s3QSTqXI+6o6UvsUZN/9P
T1wIcT7+Ticy69dNImqJk2ML98JBuGkeziYTITwRgnfZdSOsQbt+ejV9lOq18gPU
KjtyWYDI7fFAAUgwdk2gm8sGzrVhKxpTUrfNYYxTyorNkn4+t4bOZzAshSY24LH2
k6GHUQm92SsVN8WoLYwjLw6TPy5yFaBwM7u3U+gPZpkUMDQA/jl3iYp0NOLUfwO7
Bt61UTuBeSGnoNPtyJ4eanBe6GBEKaXDNHzvSKx2ZNawssWzY8LOq7fQddB/ZAxH
jsC7kypslVta7ZZtygzmnnoCQ3b8S4BJDrhWAAoLXZMlwckIf/2zpNyIYS/QGoFj
+vwuOUAD28UEn6DIkX+GYWz0ElFAYpLj3h78y1tuRy2zY6LX7zJ5s+03GvzxqQpH
unl1rxoFhfRAK8CVbhSvSA31YHk5tJKR6cG+cFUYDHI9SzFAulfbZOlKQZ30pZ5n
W7IXp/mvHsmd+/A7Dy3UgYcPHPOO/mZCWoh/iExuOHovVUlyvlSrRqmvbgiAsKWJ
iwnzlbIxZVH84ht5zmj8f8n77gh/vNmTiPCiyxZs9zu32BOEOaztNS/MU5vtD9Fl
3vMK3Wj1y3mpwzvZblVMbBmagsZpIz8LnmmqVcP2LvejJxYgJ4890mUHChbnAfAS
3yD3D0FK71vjgSndHMRannuGrAVTsR/gCc9W1NWw0zvhnlODhi1zzW6ki9OEmt0Z
nWNUrgWrhH/XEjI22YyYVLB8s3qsJzDv7qxdn012x46vNHdzyAikhOGHLo5mQaKr
WrlS3rjTvD0ZQjoC+FTkhh0tVC/Igo94uRfBhDj/EF5r8gkS4xRtNqQCBGQP+6CV
TwlsSz/VoStoABewic9JorM+FWysLAsV/+GpWRh9XRklkvPEn65S2ClZurl0vX3y
Kg495pS0Ad9hqLyN7yCM/pRWrJVcqbiejaCk0tnMkIDU+FUhKYlQGhjiXrgGCUi+
izJYRenDvbJ+Hcg/ei+4Xj7FctUqCSvoEQ9spmuIRGoSlJWXsqQ35BKabzi6kKW8
dd8Gdk84v8/zLPqf1Ry3N4gC2je7x63oVXqo9uV4oL+mKG2xG1wSOK9Q3mJbThbb
ZzYkZor6ZStW51ZRq9bxLe06OLeP4cFB8bumJQ9dQg1CnSksL8C8lwV78owLnAh/
sbheUmrTtpVahRege5lroaIfaM7rzdtrivXJVzBXllQCEtJ2guJ2w9aQkM0TMIcY
QsZVvo6Td1Qlg4+T545oRbYPEqH0SGqmke6l39bTiuhDX8uqEAiKwz6STWAHpANt
TMvE3NetLUQXYbq1U3JwWtsHZP/11TnEGkjKCiZ1ByJTmumaGRnI6hso9nUOgR2Q
cRb3Sdf8VNGX5kbk5DpucplLohs1ei5xPVrDboH0jtqIsNIVwSKmPTujV84t2Vju
dySFtEGpCXAfyXT/wrKN/7AstUB1lnG1ThKyLsaKOEd1DIMgay2yDBAtlLdVhs7W
Uet3ePS90NeIP+No1ZYQokb/qiSTut72I+mGprEa7iOCFQlnf1bdmehpcsX/gnep
DFxkoUXVqiExCArRFQA7lLfb5BOJfaFSmmwzwTH/Y08SEFTw0tE3MOT/cLKTWouw
A11BoVjurjavVWcwzd8DGCxRxlZBwMLBqe0CFOtKUtRXaKVdxCSq2dVT1Ruzm4tB
BRBoqDmwQI9ibf3ZpotzPbhNxwOnIUwclcVXOKGrmoG6yah69Xte9p1p9EYJaT6f
BluUYKDi0OIlkG49DqPiHwb26KB5WYZ/CelfCrstDjYQmeRsouqICDkjd2DePuy5
7vxqpgjeGWofIFy/5ch1RJd/wsXTjuxdI37zKO2w3nmsnK4TfoqdjrvK11X6v3Sv
68VYHNni8i9TCHcl1J5xggJ+Xrkv3eLuSftY+pCv9Ot6kWfGpSJBIuFMHmefOcOZ
dPk7WEAHtP1ba74A88poZg8PBovOwm9vec1v7RjOcEDbOzEuzJhUNa8J0ijMKqpG
ZyIbvn85jR5BcP2VWY3swpM2JpxqUdqqwL5wxomAba4RJ09bUPAE4H9CuRKmRvgJ
mdEqKGj0SoP2ve+TdDr9TdeZZYM2KwNH93ECAeYYVkIztdAA0Z3vqLazeCsWeQSV
NgLcaX1tuR/TTu4mwSTCUO5123yRmxPUapoBIMAZR1HDK/GJiAAWOfotEvM0grEg
wkcTZ5gmwqGRNtMJiswIA3UZX095KnaHzH9YXuvi+9fC6b9F8FR5CaOpKO5GeIuN
Zr22+4oYW+XJtswwI2nJeuNgbraMlnaYTp0xmckUTjz13hJ30fNANajuiSA+EXKf
UvD5XXfKnWlIez6d0JSyzpBVYJT6ya/eVYt3YqibwFDMCjVaYtWIn1FW15mxOvtm
w4MPpbbfaCKg8exj0GDhkVkeWpzQ7rcjsbL6+unye5q70rtGG0wvBVgRtPSHuuLv
wyKYE1HhU2s82PNfJ164mWpKLzAkfQZMxoB4TSBMkS4mrG9nz8nuyEL92oWHNVqt
3bhMe8m6nkJdCGrPx5EmW08leNqzjIRrlVZE5dCu10RNXpBzVFALcKWbsrbx730f
tHlxewpWmUdC+hwVMHn5o4ZtD+dN1gXj120MOlBb2DH0J/Wr9fR7kNmOyLG5CJF2
z5f6Gvo3MJZ96Rb76HdAKKgKOAUuiHg8Lx+DaF525D+ibDI9+yO4Mqc4p3RhITO3
RToBk5mJ4j0edQwOpdnmX5nIdLGNZMVCJFXKIb76ZFRoTW4R5gq0gNsMq98DD40q
uk+uC59wv4V4aoB3V1fJIoZVNmRDk5YR3b+Ldt5491kf6Hpk4iZF2iuODDP3dIpn
WJCPZq6/guTfFRjijt3HZbI4KWvHpqEO6twyxb94XKIEwR/o2fqrAuckzdIwqjlN
cbolt4SXiDcyuz5oP6Xa8qPzYRicmrK0smhBDd1yN0uj0FGioY7MeV/lhphmAZhS
XyfDfag5c04OZsvYRSsuLLrRG19uRPIFFRtxKHxrn5nI5PIrBfhaLMXMclYWWtzZ
61G9ECjY/4Z9MnJAkoKdYpxd/80U/Casgy8UAVJ4RvDWZP14zVLDf+NWAvgenP6e
VrPL+RFX8jMg/A+0Qd4JbGLgcQwRbH0ieXl2BGVz1HdMnTCQODyiyItwegkMnM7T
LmTQQrV0O8G+UJzDWV06+IjkLDrWYZvw/RYYHUyGk+5ahFu7GdOWXpILpo1jnMpJ
TtPog1S+FGxLfUj0S07mwxyuqpiyb3B2UI80FPB/jpvRhCWMS3uHJEYUlU9MPIgo
/9p+cTdQ+WU/Anr7It9P2xWc76nKUObDNql/m6jHsHQEd6bf1kWJ7plMl0Y2H2Q9
livLPvCQYaHNQ7KDoLnCAZEDvR+1rsxS+X7lchfTJnCKbd9X7my2TZSPaORhYQNV
H9+aV49hrdEP12KxB5476OcVzexD3nvTnwgQMzwkXEPFiNEhOgXXlWNWULRQYon7
JFCjdPpmtEBnikxYe2Z5rTyO5hTNuzUWnw8tScbKN81m2GnjUK+DeOkAZofX5aBH
0YAFHSM7uht36MH/h8onLh2ACOmYf3FTD/4cFOEKYZ+/Y0lVp0Ch8Bj2/sZdHdXO
71Km0fdnwq6kZ/Fw14PIbtK11d1U4JAmnR/nvh30P7MIa9uobIJsYMUNg2GSd2lK
ZGiP7Cgm8eCR8fX+CKfP+2H//pZdPXZIhzUnS1vGzsQG+bnMB49VD/8UtGVcoPU3
H2iPTX216UepZXP5Sh77a2zNtvUZW60uh/66Wb/QLGq0YHo5euhBBxn1PxJ5gyzo
1D/VEzpEVgECbkPZLRGhkD1INeDqjcrfVnvlyo0Tb0FG/EhnJgDAzf3X3j5WmTU/
d158MRrD9SLqoocj3xuVy8GwHSfbceB9654TYe+VZSKMQ9BNH5xhfQL0EdKQU5C7
p0ONyk265Nt8hBLY5ceWyr1an3y6EGmFL5dId7QH/5hmObfcWvDs/8dvWuNNjrwv
faeynJRurDtEd3EryIh/LvxJt5U1ifilHc4RpUYGRWUHz83dKhmflgEXbKrfwVCD
nb42NjfQ3Oe/UhZQ502PSrAh7aEkMPldBMBNoFrSD4sCx4RCxEKX8PuVBSaLw8bo
Vm7RWUutH4hFtkI9H/rouVScvZoncq6ObyymjS+tR61rPNjwGw10mZDlIOKQGITy
pQAPon2P4/Bii0Pq5ZSZ1lgYdfvumbR7lp9rIYU9Diq5uSYE/P/NASDscKgmD0ie
2Vc/TuHGm9GdmONP7MKmEmZJmuqDMr2tIXfPW8tFD8mU/tg9KrdLh1GuwITtGrf7
yCkuk+tvB4AsJCk0CaJj/F7TRquphCYNYnv/WMNoB+yJlRL3gSqApVWa6a7p4svG
uJQBjLIwE/xTeGOSWMcLen7uOgAJ6xmH993RGHUNv5m3oZGN40e1FNuHT5wR36sy
9Elo1l0KVYKbl/bG53TuIWVhvRX1/Ma014BuOATSBxqvG7ub+kM0zsLvPiL8sSy4
eUqUoOlLmWJveBD7YoVo/8wWuwtY9ZKn7hKmvQWRk8CRnfSFPQntbshIf2uWJBPe
GZc+SLTtyVGKqs0qtVtv0aR65WclLa8hQLFJHwkL7yyhIHw3yGyaTd1aCHW+052w
VsCkVAS5QTwp9fujmPtBDm/vEn+6CRNs+UYzMkKX3pbkOpGW9dUCbzUayf/5lApH
njBV8UX6SwXW7M20t10kimCKG/x8LJc91F8ZGyqpIGGfO+4tXVOyLYsn5KK0NPbD
XU3Z9IdTnxbFCqlhR7xGfjWBDMXcNXtnAgV++wEzNpF4QY25P5GbHnl8UAo9Ptqd
YxsxR/L7cCs/MdNSbqbq0Gnuoph18dr4Zih5C4503K6pAM1acQt+ZTH4MM81uXuV
Vqi1zzIwDaziXdJI6kp3qHYlMzGquw4B5yuZ9hX1QMQBMZi4gsroe9gWa/RmnO5C
6MH71eZCkbMb8dpdGtnm5Yr8dwGClaoq1OcJrC3j9O+a44H1zmzhLz0vtnxZkjE4
HXTofHWygJKx0NH1bI+tbcp2LM36ZJLIsvKGWfLdFh8aZ882bYmVKH2SmfuuuNfG
Wf9rTuVKkr/8gfocvsyCuTFzTDSkEvunXgtb83EruAd+2ZaDQH1fFFV3PcCavVz9
NtFAgwGANjCz3nX+ibQaW5kqGkCIlgRtm6Cz5ds+1v6jMT3o7ISfz1G8mwXWHlzF
/nyzb6rWXuCvSMh/TyCw7iufZQ3dbRZcNtd67ck2WxmKz1TiYkZzC0Se/ZtShUiC
L/kKCmmyxmzZ26/8NBXuCqiTEMpZ6o9wMi7TogZYx3JMHeNWRfukPIb3VR8FACwl
XXr632CVrs6rVzVxRjYf0CRqJuaFVuYXQQ4iPqKUDIhRvVFKfTR09ovgFiNZtlpO
Pn6DZhYQf3t+5gAkI5jFbXtMUJLhpoj57yZIyC9ascu+bkkhpVHv7L60Gh3rtnjk
W7iXtSfq2GsU/ADatiLA9fEFjZiJ/U2HduFAf+MIWnfUYtfe902vF5Eyh4RKt8rL
RsM/IJ9msrdwhpNo40DwCdLuWwWeM5WGedkjd/Dis1Ysq9BcS1J+D5uiK8aIw12C
Tpc3VpvCXSbzBwnl9QLR4sUks74M2tPa5AxNDzeIxpq0VzGX3GD6y2xwUtCqYMmE
Pd5p8qiNNcUstD9nqMoTAscVK4hEYUd3xPTHcZrbs+NTA8U9q/gMfLFEiNhsfSkb
xIecovuAoEliLDz827BZzp/yka0rGu/3vEOVaGvdDbgWF9UgKSX8xQTcW8oRaf1g
GXCKgn5m2FU6KxM93B1i3EciCnruPF1QWNWTS2K844WPA8PWWByd5ip7lbsB2vF+
Q+v5eWt8+ksj0D5a72TKrT8RzteLpxPTyUUeS39yFCahQaqbPihcFkz9u0W5D5zv
tYq5yxG3pEVGVB4ziwR4liwuduf2FpwFbDMiMQmZ9hx3b9E//TZ/BpzAw3NEM76g
DR/BUoDL8xnLWV4bRRg4L790LQHzIRprbXPrMFeWLcBBgd2RxzHpu4nw16+xOBw6
9TCpCIp7nHu8mLOWFCKU0u6TtnpEsrzfP/HeaAQT4IBt9a58Zzcshmn+YvZ6rlT8
8OuSe5nsMh1sfP3Sch8tKt+XQMM9W0DpAoXui8J8gzX5Zl1s1j3YhJ+eztF8TYWe
5O2BxrA2dYNj5FIfbpUVc4kguC6S2xPfWdb3FteYdtgnBnT0Wxlarrht3pHNKcBh
U/xYgEuNNLQcxuek48Lmif4YYSDVFO2ZytXrAkGndEuyDmgGn17A4TQHANjIM6ZC
AhSUgmxLicnDi/OmrPqNaJzC1S5HqjPSBQNxGc5OOPh3Ik251xRctOOvqkhuiIyv
9PIig8jP0Lrmsg65Qc9bUdCJBiJbrcGyF0WuK+SizGO4f+VPvRMUQRUeMCc63BBE
5cMD7S3bghtcXNVugeiVtK7ibxg/Jy/wfXgbrHTowhddLx3FHad7oL7Hj6Nvwbak
5iKj86F1X+I3Z2sCB2VuIM5kwenJXJaJ28zOD1WgeiEXgRnVBoih+NtBYmaP5Ywi
YWI0dSzu+1hgq4+mw06Dt9pQZ3grzrSU67vmhgLFdkQZQalTMXwKESz6YGjP45xu
tSLKIxmQimXQGe02qh19JWGI086rGBTVsM9y1BqaW+xWeKvjhj3qLBDuoQlhzPet
QlmomzwoKVX/uBrDvlkHiRnlRmCh29qUkB1v33JF1ZfokPsHRjYx3Ddy3rLtJX4Y
jGR2/oIrLI5/NpMA4mGUlSbH2uP4hKiSJjvPyCtxNgKVnuaPqM16Cy7gi1EM/M8/
Z6LDEk53e5Mu0ksH04jkG6CiPRkslcR6Us5NW/II9Y+NQcmwCAfo/pMQx/rh6Gag
OwFn2uXONeX7uRubCLCTOvoGWiwFAd/uizTS85yAgSvOk1cL/wNDfaRPHcaf78du
olzCkiSNLnR+oJUqd7M2/PuYFudTq3k16nJcjVxB5jKzoFBiRUdQ1DukPwIx2zFI
V/TmMgoXpQlsd2LuTb47CGKvSht+pI7T/38BClsWQOWNKJqpRnbtu2ITcKMnwRo7
0x1+2iB7Yfn/vuYflMDt9yyRpDicoQow1RRzccA37G8OJenAH00gkbaUlCexmooD
u6VkrhX53tE33U8lUYOrrPC8Q/BGCWHaPr48x/BLUwt8M+sMo0mTY6v9Rz3ZBXkG
XkX5l6WTojvJx8p4kKyrCSngFPMfmPXI20y6W5/kDYJE0HyDdr5yTim6R7ftQ2Tn
QpIYdYOf+QFAexRcRDyaApvmcqLs1IMgRgGVhyng1muVz2ER4g0UIMlC0cFdTtra
Fddg12goP/4Xl4ENOtZlOqaPGDN3KphsBZ88a69pUuRRMatCwVQPQR4jE+iaq5/A
KxLZTF6sR83Wt7WX1EuvG69thaygPGeciM8fuf70NDtktfNNa1NhynbVOIpfcTOj
9A+9R5bnvU2/q2khURuGLCMIx80HpQhAEBMLbxIbvIClSLXKQs/nZ5Ylt7SjCeuq
IqeAkZuXxdpswD0mWwXYj+XziNqwpo5eWZlYltT6YMmkheyVoOXYyvQaxKsk79GJ
d3EXbnEytYhdXpw0nUmiF48v28guJOrsLoetpCX6c5kLl/TQ/unQnklbrTh1utYG
pRrrB+/uDGeHTzoRwBjZZPfZzHcXPdEqfAb22LmV/tKwaYRNDVXOMKA2BuNbt9Q1
M9Rp0fz+M0JLiAD5WGypAiG6kbNny0u51BP4NfEH6aXly+eaaWCSR6z1/MNKivnx
5g+/6UpY+vvBX4bZVBD0sKtIuQ3oSnaicNedg620qvJHyBKY0l57WLWJQul+jXJf
WWdkbssy8Tg8Ernb973LBq2hKmBkCHNpUkgqWiGdjwLBCbFf+gubZLYcx5cbM7tL
rzmZGmyjhlE1J/8O2i6IhlJ4SE6QwViMfTki95o4p9Km4xi875lrftPJjMGBgJpL
7YwhyaklA6XMKsPLLSP8AClPAg4bsQH7nBmMOBSi9vpz6hDzwku+ubmxHCHF+lVp
2UCdHeNDElOTpXnob8JnaBnSwnGMRoJqff22BGmv9tmn5Mvvh9W/Myi2VJyUEEkk
1lNHY14tUv5UIgZsK7SEdgkjMlSynxZ5Mq0kB1dAKs0FISxfc422ZLj8ZBjzRrm/
+lXb+JKStCAIeHmBWZxD8cA0zBR+JhXzYeUA81ENKrBMNRVoAYpWv72Gj0SigCjc
m6LZKsYkS1ygn+h4I9JhI+3pihT+b7NCpWqjICT5mWbK7HWNt/6T6G3TWWTXlyIP
eqYGYecQijg3xyJfcuH/jKif21YFCIYFayzlv+Y9TUR1/tz47igLUIHpGL09YO40
Gxd+/lz4G1TSR7mEchNnnf0fr8dVfrVyEFGUtIa/HNm+ssRNKdAwsD/pYSttmsLD
Ee00vUX5RgnKd/V5IuHr/7Aj4Szuub81RGLwi2YmWOibX/VJA6gMKKU8YdlvkJjP
Elrwsx0QKprmaR8fJRYJpzEJVBvpOtzf0FTqPdjZxYITK8xBJ96nInVRdXmIyg6p
2VV1POLGvcEgAmZBgtvVznYe75rCFqwKDBK2sk5uqxYJm08PRQkQRh+6kerdStqZ
AHce+9B5NYPwNm/MDcOTqPN59Eiykc8i68jp7EejNEbqY7C8dJyKIHDKASPHnGL8
oKvcGNFjU0Owc7iKTGb0NomUoCq/2XbRd4Wuvj16POpfkt5qk0Ql2SdU/LywjM8q
g3sTkjnvbVeZ2xe7mYrKquuR/WuDMbTiU9e+KUkqElHXAEJrw6F2KVlbYs3WxlIp
Tq7pBPcXNzAe4vH4YGLCXdCJdGnp0cnK1J6gJ7LVUm5f9157QeVRm7uTM2+34c9l
P/P8MAl3FGiKg1wnIBnst9Kl/x1n8NFvhnBzgxUmUh58SrJiEBIrtKFWeIxU4V8O
feRuqugItNnmmrBwxoFun0UI0ns/A51GIbXzHC2B74SefPkb40sg/HtNyijuuIHN
z0Vpaj6f75n6A4xsoFFmtfNOk28suQM64Pr3An+q4skgQBMLGIBpzbrWVpBBu/un
y1osWa/O1QQNID6UnhnqnQqBxBnyIwVuy3O1dxLwtRcoU8JU85shvgSIiCkOSK0w
`protect END_PROTECTED
