`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/cJVsI8qUSmAQmYz/JsdDGzae5YhFTS/HgI87KB5LzpO2dM/22bvNjvOeRA4gLm
gKVq2EBmg293wnsJ1SWMFziYz4nugL0lDBUMBURvxa3na1Mqw2viyEmHRkmK2xO4
Dve+g2+dEH0521EmjpRUT0yLTgytfsjeU0wQkGC3l1HXDi1k6UX8SUg67TFzwp2j
svP8VFAvF5Qp0+OGHU6qyVnvnNVftbtCm0MV6UYkNf4wW2cilsBFba80HshPlNlw
qemO7uLbbTqWfiNDlvJWS+s1d8lHT4fEsP9Kt8VFlFj58FNaPhUsVQ1nXduJniqH
4dLt1O/eqD4L83mHg4iA0UPE2EHDQKRa1Uk1ObEJRL+cX6xyPdCGzfjd2BGaVmVP
SF6SrdWDxO5YPMyCdnWC3bo9xi9v18XONahtw6ey3jPYCM/3OJfe9LasMGDhnP6a
ZxNi6EP99EtJUnRhEDTCvhcozUFeeQplwcMheq8ITdHKe5N41e30PpSNaYXxk7G5
jQajZkuF00oMcSg9c++mJY6IGpIcGdEdxNuSrHXMwKbmooqCapTmyl4OsaHYQ8oF
W2pwXtPRtc6fE1U7xAhwMBZt++yvE+but4PEQ0m9ZqMtecmn/nG7GtBjOOh09gm3
FvpVwGpuxDezO1widkidd3ZRAD1/qKMXZ8YciZdonEiikEfeUq9yaQt/TEorF+h+
Nh3TwZ87OlLDZUynUmDYyxNfebuY5mC2Ar28MwKHppfqZrJkd8x6IBOE7+t2miLf
HV9RwqEy0JqxaxHsOSAU76wulhPFHFJ+4Rrdx79Wz5kFM+rLHklFRGi6ubYV/MMu
KxYZFcOJUFu2Kr4HohMnUF3Ov6RsbRJGWF/n08cpkSM=
`protect END_PROTECTED
