`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+D3b6fdvx0j94YPDrUcNp2VV7jTTk41k6zAn1OY0TGf7I1O4+EP68SAnqOODZ+hV
uJgIepR2LiCs8t0opZ25int+s75MFrqTP0DA/h+zdlawQIqWm6Ll8xkIzil0UPGu
keF4slnbJ3yKoQy46jIyD4ZtJSjdkGSu7ndvVtyYfZqyrkvl0v+NYfNKzbc1FqCL
VvLqHQ/sWiuSq43GauU6GFzgEyvmDVJIZ+Tyl9U55AylF6wR7YsqG+2548Voc9yr
InKcnoHPbwz2YrH28i16kB8jEOVcPZJ98zLwfGlKPf+6Tf0QSpfg/pnJcHTxky4p
qS6U1NSAx2SXPXBhZEAe6CMBNZOp5iYjCPpvOWjQ4DzTxjsOpXFqfivlWHxP15gP
rTyVfYCPPzh15SGM6VDp/O7KQ/QFEsxdFk5Jy5Fu7uy9d3po/4Vm48Z9NO5nkGzG
QuUKt5JU91RqpAAlJSzxMxnlW2Qk3oPZjkRhp4mUqsHve+ikkSnX4kkQ27a8sbgY
TzEhQPFZt2o1GRxlfDC5KOctlWWVcErG7kC3M/nYSsa1/HWWbWp/CQfDJrXKwT44
9M2PTwJI2twPfrcgBD08rXreFp3+BZCthcIF+saXcgO0CmPlvAuY4v9nKdtiTDzA
JCEzu0NtMM0jmcKdQvRehoEh/Mr1c2icxhGWAlojdy48+R5+elSbtbC/fZjIQ05N
3TmCiPHuCab0EbLsgiA+BjDCKEtVxEUeOWSd/TsKdX1fLP5gyP6twLaBNAk6Y8yx
8WTfeaSJBaNYHawp33Pca2u9S7eO3i2CK+aK4EVkvaDL2nl3/XOl2wU5nbhlqllk
PwsLuJnkFZic5M/uaSZEiuVWnWlqoFmJWBfN57UbUlSOG7vyydgHXNaLuLoZ0JZr
nu3G1KuMKBGIG6Ucy2onaqAOVFhC5NCUAhguNZ/IeAOBF75Xy4VECbXOGwIm0LQd
e70wsGYmNy+iAW0dtGYqEE9nluXA3rbqCwwakMVyjhxUU1jfU9KCJfzCfi0Gb0os
dbJq4G6lPL5dxAIfpLoUqHfm3sFL20NW9uby8cOHY0XysXiwWCYkEgDju/7vZnFX
6cha7kU8NlRvymVqgrM37UWG1Nq0kPws6MoBl9JgWjcUNRV/B/9Wxr3iovgooduh
I5ir40h73EV4HDaolKuYn5pqF2IJv0l9y235b6dKirvXL1Jnb/M7S9vXYLjKL4LZ
TfZgn7OxoHMGxH/k0e+i/iFWIsLDoSrxBJu1QnRFu/q5z5Mw9Ali/mRVfp/lSO7x
EnO+cgTWwPeulgw5LI+dXttDQMyHTRDfPIqc08js0Htw0KSBppUWlwq4PQURPHVI
zODDpQ4VlpE0A2k957nW/r0Vd8xrLTtMUSfXmzERn3/HugROcTF/3NZZblHRRDA9
BXl0qvw26CHbLxI/NX9Z5h65N9gAJ5w1Y48BjZCGBOSshCP2E0NCsjHJOzJ8WH3h
zHosyW9deoZt5VzJy5lfS/3fFvMZ3j4k421mrIvJDoUCifAQay0qKp0x8WmkDNBc
lPVAUbGb3cjYcZGqAFnrLPHTiquyUqecp+noqeH6zQlQuBsNn6ToSWvb1HQpfdoL
aIcO05hc+sWiMMYVkC/Wf9WddGmQ0HFkCBwXpxIt3SLl6rq62+VZYgtJZu4Habw2
CmXcCElIF0OstzvDkQxKqOLaX4uPK93HVOb4AsIh3JtiX939hJoFPhcyyH8BMSnF
N1z1G6gjWUtznp46ZUpGkL4bhW5Yj4ZhHOvWjH0mj3o=
`protect END_PROTECTED
