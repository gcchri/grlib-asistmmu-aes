`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kD4nNIJcoF30UVteHHRGWiMArprw0VM5GE6IedTaUht3SESvhSPMawd40aRL37ZL
/EepYKjcx5fHb+RVnjrXnjl+POxrKcc08Am9cR4LrtIbKkfyZLH46gOcINd8MaC8
+9LdNo51IDJbxcovWLZZLMwYILZOfIAh6FAJ1lHk5gTrFjcujpfpA2EHRt/1kwek
b4uXLU+tCTmXYtDa486Egr/+sTgoo5j4nOD6WwUtmeaxF2RsGl+lqM1RvSuJJbBt
IztnkRslfLH0vO/xD5diuT8AhSpm1/0QsO/WsCxqwwqV31YAkDdANafUHtrI0QTA
iY/pnnjs8XQuKtUZzJr63SQhENypeKZ6p8T4q8wicupa1k8mc4p2rqAuYVFsSsEh
5ftMcYGocluiYD2ZiSneGLtGTit0+xEQTjk0MBKrDzbFssrhjxiYAXBC1SfQZi0A
WL3rOBHeQbVmx5ISrCOYjVsGEXWJSDvAXEcE2aB7RP8twNXzXqnv8TMGm5ljLZjp
PaFHftSx9mlS+b0LTPC7o7cHJDZxfU+ohp3AFiT+g2bX0cNaXHKRm5UNDH7N6cn1
MR/sahSojT02vXdZNEsNkx5wVWzqD3x2/oT+/0n4XRNp0aiOMsmiNV6RSSqD9lS9
LrZxBJizCaf1N7pB8uoKCs60NfCWSEXAw1GESNNRbcwKSryaWuqLkOyqowgWO1e3
qg0iW2AUBHHVkueuQG78rUApMiY1SgGSwPymOBkOxsF/lovlElTB3N/5oo00hJ3L
D2QQrQ62W38y4IWkQcMwu/JKAB7SQReZZIj6qahRgj2tfHx1KT9KcJ/VHqSxtfcv
orAMNVYQteRhIo3aRUQSCn0P/XuVMpRSrFYDaMcSRUSoVwb/C6vxzX343o69bjPq
A7jpOoEnt4e6C37OdRAQwHybrUaevxmNIE34pQQJU2sjuuXDF/QMZw8PIkaaJi2b
BccjRaQ1D8WeCcIdcjbeCBzjlkWI969ENgs+IsLQTpkWulVLZrshr8KUG1JqY//x
uoU+3Zd4ZivGsLPoDWzG00ExIQdYs0e7PIPTmvXnRNv+1nMnjXg07Zc47e9n2hYv
7wjAxu5fTsWi2H+PU0fffl1e0WsdAswXBEtIh9BUyLYiozLM9QrE2zDHboa6/Gxd
UyDGpD4QvpMz0aQnHea8oMR1BCgjbzLs+7NTDFn9WbSQWd2Rj5zSj7+66aacvSs/
v3DymIg36R4/kBF7n80U9kEYN5kOsbfaZHH8XIaiEz/ozWQppTatFanhvUmVqrlA
A+uBKyAVnp6CYamzjDKJNm0q+/fkb4ONoZ/2cVRvuwDrz0ZH6no/CNmkzFh/XxnH
WB5qbhwd2Uryj4VgphJXAeV/QdWhsqZ2zEhLUCwXoQ3sL1gcNXZAAh4sBMCZOuF8
o1BuEUrOpFQRmBEpQEHXGV5maiaAWR5/55GY/jLWK1O6Y13Q77IiA6LoOipHYvjM
joSeSdnpLr62lDAeV5+ItdtC9UAYV92YA6K9FpJ3EvAgAC+7qs4Z5BbGus0mKiSn
/33/PUdMu8QcFO7rYqL1HB1UZkqA7VOcw67uJ1MzY92nhg9QhBYgotI/3CpK6gDE
n+FbDHoWVnL93feQgDQ1jp5robUI6x5VM0HLsIQREUGrJLllqFhJiTk+tjSd2Nik
DLAtCK+3ncZ+VEtrcIjSdIwh+D1Qv35UKNSS+Fo4vCg4lfg1F7Bi2eVhEKMC0cKe
Aqk51/VGXbWfSZEhZ3iyx5VHyPHBK4MQpMcpm8JGhC5NK6QZLJPpw04dAh3lBtkq
4eGI32Cvr2eKG/BgEwSKcpR1ODOWeT3olLTZC6QwVcMjmAtsmS6ZyTC2Fu4Gr3qs
vtuiVzeJ0NDQTyNU7yUSIU/K6j9V3Z0VgsEiSwzg8FtwHEW0T58LIwxXIeqBTF1K
F1sIPwwWd5CxhDo0WTRf8qJkPqaq2elIOU3eNNHT8ovfKJVaP+A+Sn0akSWJN6B3
KEyxIR/sHgvJn0zSlboP0QNyopR84fv5GGz5VR4pGlOolaubcQSrTrGa8BWtcE6G
i4bVvyWIVMlcAyYkUUtFakZVSApCoAbEQad11NmCLedlMj7YLg9ENIUFcWYzemki
BhA6cEnxW+PllI85yrAMPbX5C3XcfsEqYLMfnIvfg1+RLb0pzOxZpxDU18atSCS3
O/wJ8Cesj5a4oi7fVw5FoXml/mnJPXM+idxsMjaMeyvyhHlRzTEDIIcWh0YQ2ws8
bCXj/wux5FOtbd42RxLD5f6kbLn8UbzU38ZRzAU8fv+LdyDfWcltmyAtsJufdh8H
1qMdUw770VB7Tat3+Dags20Xim4g6NuETo96+Qd18ZkcGlwZwUNGljptwmsCzP9t
/pwvRxsH3TbPV6ZnWxrLZTSfpjDRUrSbcc9eIPW3cdEOunjHqKthA7zym5JGlZX9
hsmpBH17HeUUEKja6k9U8q6Sx2CRHMVI2aXkQ/gjnJuBNZGvop51b4r+/qzDcybJ
uLB297vU3jFn7B5sciDLwhZLQK2Xt+NhjZ9Q07Qh7ISKx1HlA8V15ZezJq0GDGD8
t0iw5RSmG08KyYAk7yJQlBLYEhrK4z8NLh62YhhNUcsME1QSJe4Vg5XIY2xWKzMK
dPqdoL+6JjSgrFHtDRlCVDTs03wvYFYQLLydPg3EQPJaFf6sV8GtWyu9Z4q315xc
dZAwkoYiTkbIDnnhbqtMqq+lO0jnLWOxN2lH/TDQy24CxWxT0DcAsURDxo+l6Ih2
ZrWs/7c2MEi0VAEcbPFXjg==
`protect END_PROTECTED
