`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUNwke8YsQEpVhp6k3NhxM3Y6ov+lvK4kc4z6/N7DWJzWL0WvdmbemiFcZY81FzG
tB38W50hUTD9UJowQfujEFwheNBCWKNVZW9n8NCh9T0IBjJEhU36Bjbqe5d5NQIE
/89JvbHvg3t41LikgKgpgGv6QLeGIU3P/Fl4RI5ZE6KW8Nr5ljxK7EXq1T6uwdvo
xgbx4up7pusVAxO1sZ2SUIgIw5AcqWcklM23VOQom/pPYeKBaUztF6jKGcC45MO6
lb6nRuqvcMYOoOc1eFxbsy3lweLswRRHBrpI8FGvtYkKaCD3qc+HYTOrW0rhkqpL
IKqLlpDcntvGQEykv0yyfYfV+q7DBNv770LzHEi6OBz2JcUiRItlEe118Cx4p9Wz
CFdHgE2Gp72inDJvePcqOvbEPmDdlkXCCWKMD1eCqPekvJRyPUip9H2v2qWhXhtp
kFACfXveVeKS+IJuvCenJUtZCnxAz2wQF7UOe3HzeFrLxnwiEsUYSDK+6xakEKBv
6tQrRcHkLH1dxJYInNj60TaEslvAnj0nizq0ONcmz2e/KBPG1aYrFSC9tlUHj+yb
ytocuOvVzrif08oVL3N2Q2Sbmt4Y1CA6wBVy/cy8iNt8j0LyXQK3fxOATtDt96fr
ViEPHkX4QXdYpdoA+XdqJqEZlLBPZMN2/7XhUZIzRqBu1KJq1bhHf++YWtwm36ei
krJATW2ngu39HsXwKz6xVqoB/r2IJUTIqegMLizGT/VKTklI6GDBPhLGhilrRFu5
FcEU5nWDuWK/d79Ts+XadCeEdLQqIU9sDec1cbeEOKRZMKnZKHfaM0cCyvnlNQ6x
T48O2cj71ORUUpB+IqVRU4vVUEkDARZH1Bum99fBk/uLj8gT83x6/EXHQZ6iZGyK
S0npkHX13hTyrR+tlaG2CHhu12cPE9SyrCU/y/+/dmGPg+4MF/osyNbWC7pY3QZU
gJDk82ivQRFU4J0mPqPz8hPWMVSoA3QIERICkibB2E1z9svnm+sTrpsGC6T6eeQU
j4+Z5/ptySeJQx6v73lt0A==
`protect END_PROTECTED
