`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UHYK49kAywW5VyW0xXibjxlTptj3LDDXNV5bxFsIREeVSR/1r2eE3sVceuu4QwPN
m3l2N66DLzh3MNGHUBl/b87ORB3f6u2mWD1jbfEQ6szEX0ONZfgIWSzt4GJ/g5Ny
Gtk0h99v91MaxeJipdB4Iy5TKP3rqAZGMEkaq3SZn2snSKnhnkHT6M5EJsSo4a1V
0GsvMfK4/oqU+RUJlEGglkr4sOqeZAy7azH5ucX4bJfE0yT+QURPYlaCg3cUw6yM
7B1jF2F1ECR7DJ/S6VvkRNtj75+WL44AZ82P53dyFlTZ9/1LDXapxrb5ESP59gGl
d3YpQv+Z/vLkEv/fZPKhxVn4hJoq86D7swGnVW3Ul2MYSWfVmccRovZ5w+wvlUK3
SYLUkzmti8uL1yOUTu7BAtjg0CHPgCAYGqfR0xP/ZPjPk2TZU/f6qr9zNl47PmKb
x41VxDkyfCAp4viukUA6NA==
`protect END_PROTECTED
