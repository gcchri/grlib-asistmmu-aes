`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbkWxRa1z0u15TxgMi/LDAtUykvj1/N/RlHZyr3YBP6WSD3KZWzBf6NOnkPLvLDr
vugoUj7KW9nXmGFfcQJ9progwDD5S4Bj7VW4b5MbTXFIrsnOIzx+qjI1t4PUK2O2
qefieCSwhU3o0z0Tig97TjzDL5OTPtrYU3DvWOo5zvMw+Jh4M2ITvxVcTnDjNGka
xvB5YpzqXP0mZn2GyDBm5aeXeoaK5+Ifg++E8OvzHz1Q77bwza/AUzI1LqKC9Qqc
i4QUuMlJFpryw2GE1uO7k3ieN9dR0YNYHPLdRmlogrYoPmt+X1UWRnkGVRW8pic0
emCNsh5LyDzjGC3JFWCxgNmryyjGKXoto67657GJyYiniOK7p1OBidg0DUk/VUct
GC9AtoB/UmPVQ6vCsQFzzgt0YAemhSSykVzBIhM+gecClDj27KXTNUjXp/yA1NvX
Q0bWGoW4t/YmCtFmLv18BtC3Xadm/wiOP50D/E6cY7YgNWqcVe9E1cD/dVg+L3/F
x3/KBL/wu8NsaKRwbJmWs46iubNB2oUPT2O1rU/k34NM4eXrakANn9PEA6609jez
j++RtP7ADq2Ht8on+kpmvC5+39mbumDoGIvNkjkHP/cMqjMtDsNoN9DjultiCJw1
4nZh09GmbqK8kC0JHGrgPX8KVE5cACJLZuPBE7jEynI=
`protect END_PROTECTED
