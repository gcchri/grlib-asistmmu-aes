`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJsSkG0smYQkdzrlb/5EYtKSw3UkYQ09yLtD15lY6C6nzId1s6kqbpL6C6pCss4E
mt3xSuBGHPYC1nJoYrCiDk8Nq/J3+e3OiDhSeIzxKsffSKMIENdMik/h2N26Edbp
u76iPJcktscYC5dCGFUdtBiMRrtqNJYKEGi4mTKTJgF0KiXP2bfey1GqmGOsP3ao
5fyWJwL6/HJIWInMBauN4hoIr5KF6D1RMgg/byuGVzWjGihKIXdjD7aKrBl126zt
MVl5UdFKLg4skJP8LogM1A==
`protect END_PROTECTED
