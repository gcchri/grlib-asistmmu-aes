`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8TVyZzbd5yg8yGD/JyrdlvdCw50XnwpWcsfz9C5MPs24L5Cg3Hp9/5MLwe0CR9G5
g09I1Ms+8YQ4oD5JxJLBFB/qDSC/KCekzd3l3cuQAKHQFw7+QbHhxuLcCQYdqj+g
6APKFLo/OGse3nxoIHY5Hx/gS4GHB3xQbKwpNQ7KjYL7z/nR3jM+U1DdXs3rFrMJ
DKjIzz/MWkc3XGoswu11uozh5Yn+JLigMHmG2pW3cQsLpA1q36eeriFEk2v8OJ14
vMaK1Fi3Hz8Naj1EPVffCWBrGxzSFmCdPasglR76k95ocj9ObMbwQYL2FaKltIaN
kZKg0YzkcpHSn/qZg2B3L6bmMpiENRlv3xZJ/Rb9YyjeDKn9c43/NMs6rJlr/70g
CCkgadbLaLMtwMlg6wp3AOwM4/0lj5gG63sElZVLRgKRBMHaMiSP0F6OrKVx6Xxz
XqMminbCBR0E0c2TvnDeupgpKxMjGZIsNLNT5ETtJuXaUTi63SzfNLO938VA3UP9
i+Iwl/cDgXojK/9AHoPqL8d5E4fpFrtQoKqwjwaZdIAld/+nDj/A8D1lqoQI7bU2
eNKncyZJTvQTTnHD7Xmay1TnYLk//S/pc8NJXdqRzLMZBhmF4DLs65tbggkslr4N
44H/Q8lRmMKLucgv0qrgmTTETy6VUHi7C/ewjlxG+YXIcqC98+/7mMIU1mRqhn3X
`protect END_PROTECTED
