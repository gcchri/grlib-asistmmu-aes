`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7M9KNGfLhWq/dqFB4mEfBiKdHUJFV1BrvwYDgaORjoWdo7LNx2srfB25B8YuDhGC
jRI2nMx856cR7QdcSa/kpSRszJnD5kKKfjWJHUaY8mMjKqvFWvib7C2OfNFXZpAs
GTLvPz7qiFrQF2jjhc/xUbbvHgi27i+9rfeh9IZBmJH39T0Yj1F8WQnorpTNQhiu
zx9K7Ms8Ww406BPuubao4k4pEnOdLhodZKipx6FruQCPauSAlKqNpvABk19tZVoR
cwlZPDReDtqzT7c6DPCWTyEj3umJfHJ9EK1Ismw1tqZcQawWHVmH0pOd1qebZidL
RiWkv5QjjPm7n5jZ0WcWDgFkba8jiSqBHcGPCwhUkDkVxzxptzIiUOS7r1sI5/Zt
lHoOk8av16buUPY4eRNC5bx4GCKdLfQgwbGhdHz/FH6bPwpeoXDDA2KYPWNGg4mk
hGH859jmfMTzHB3j1Z+lCmTuj8t3PSMJk6t95tSdPbx+rL+fIkZN4lKfP217Zycl
sgi0SGySY9S6E/08V/DLm5bqhJyfccniGqouI7/NcZ9xJBTGZXg+yJlwU0VqKzcb
JG26efhC6BEv9W/EGWa2SNP7viRK2osyxkrEzuYiRRvwBD51j4APR6wDBG3jhVal
ZHVOU/mamxI/+0R5vsoJmD2fDL2GGiRT5x1dNSa4wl1zCVb6AiX+5+c4Ocx3+DhK
wxNLDHAVHa7tmT5k8XLkkqpsKwkf8NepESr7zbv7WGUXOn5OFfmfQ7jcbizT/lEZ
ieqSQYdUnpjgYqYbtnAYlL1bh03rvJjLCDR42wv7hd8CyqwcNkWAlsESASiw0H7F
/RAzxPPN/9GJ8y6YorxGfWMreSkaUHOSbWggLV4T30DnOG7+JR6eTnmYIpyR0aab
Wzk21Q02QMm1niXz5mOsMpRwOmyrT2K8281+k+hnu4PJBmvDsdeMcT0trHBVCQV3
U0rcmMI5hJIt0Hix5KrBNjyGwvSexGXsAwlBvR2ZFxaIaSbw7YP1CYBE+zUVMpwF
13vmFkOqKcBvVeGdoz4g7WO1DbtpP58wdsM1Ho0tj1zSwL+tqcdFaOAqxZ8+an9d
0laEAO8SFZgt/1C/dv4wW1r0ZPQwUewWuV1l0xAjmkIo2D6+dA+9fudFvjbD9Pxj
F90r9+9qyICw2Tli8E/4M1f08nNME39deXtUlsmTQyKaILV2VKZOQm3RK0FFClWR
zpmTHmwgiNmr5BPy3f3Jsh7sLFC0uvXF89O0Zg3iiUfU6kNEAPIYTpxEpiHnlU6J
ndYnxYCOhfmw67/AU2H5C8P1d51aukDlEklzpoXe2onGIcwudfCu+YdIni7PsqQC
xkeX6ZJMT8dlplAy0VcgdUa8y82hz3Xen20qlZDMwisHTz7PL0NGkg1/YGGX4hBZ
XtyEsM1sQ3D7vvgNNVb7IUJXA1x1r+STTu0Uzc1wWYzKg2BL68bTTHj/RSvQR9sn
9J64thA+/+WmTaOodfjyfr2oAuvORN+MeWe68/LfqKSBLw26MoMOdKEApZeUK/S7
iRmYawPe6wl8bvO/G1BXLVLBzkPvr8rbsgZqQ+S/UH54gm1grCxDY7OeciF3uYdX
v2R+VBAkL4SYJhIdoNHSe4gz6tcIfe9Eo8D9LDMNa8YDeqMQP9PwSX0k3/VlS+49
jOzeMxLkuoPIn7DlFETYfVDB18SgpocMV8wdMUfzhGdNPvpZ46zcTrRz+sIw3zXa
XVpshi0/sROqd4WGvnTtc78xr02l7Q6KKapl5nPcvBh6QFX6poRHo9TQ0MTR1g1o
zkJdeaOjEPZAs4eGNLG3y5IC0sVn0o+WzOSubvywlRtVRzZoxrVEvPisNNZVVXLy
5lZKeV+rAQpAenHR+1GB98+0aBPmcBubMpKffUQUP68Bgv9VGvmBGWUNQDm4mCDr
Q8UKIb9/a8g2rsLYBrDy7bSt7oZeqAa0vEoOmebfE2JEAVEqTmDxrJ6706wPGpNP
Z64VBLMgLEkhBqfp6ipeTsNiOWuUTWYstylZGsyt9Z26nJ0f23khYv+bl8FkKMPv
5iuIu2O/dB/1E27jrvKkZxYdxQ5fhtBadkxym2Fvc9KRxQOuHabvyFkJoZn/U3Hy
3DE7cVO4RZb2g2YYZYdVBzaeBLXWwkiF+qNHKJo4mJOkbi7CWkgUcE7JUe+Rp9mt
fRNfb3vqND8cNTkerq8EQ/wqfX/Ylwu45Ouo8sl+JbELcUReIvdPQtmxR+BQmFt7
cgyUEk+uxZP95L+mp9GUO6KUSQmka/mAayjfpV0k/o6ws8/i+4pJvkWEk8R5snjC
hBCgd+D5J3FMMHTkBPrFDvP+zKHYNa/kqDwyQlTEIa0KiTrrBKIYM0zr/Z1wg/86
`protect END_PROTECTED
