`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Ila2Bpgu5Jpqejnt3rHxqxvo6xPqZeQ3d+0Kl617zdcwcgYv/np8KAIOzGpsCgM
QxIhc/FlHy7n5rIRHgmY3WJUAu6/rhVBbCODLdxyQGlrM35uFEOuUC+v+Ve0XiIK
8hUIsUubXvvTP9/MfADHMDdy1NerhxYuON9JgjAopdTNAmeMPMOH7T42Y9c6Pvex
CsiLtUFrVws0AM+pLqMWg1zgnbXLpQz8VbMYyBkvt3AzwCRjd/qGIEhkQmi6XeOA
ig8sN8uJrvZ/VKr+ZNiVye4IvifJM4Ep85imi8yUHobKLIE0KClXw88OL34IiVHr
`protect END_PROTECTED
