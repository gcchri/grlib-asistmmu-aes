`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ka6lfxrx/H6yJydbSKSPMyELsse2unQoNVHDts2d7N8WzKqkQMJlsqmX5ngWCeAl
qjIyheM6lFCt36KyAr84HQH7PgSNkfHhhLZdIlzEuyEemJsrvqVl9xyU5E6o1Frx
GmhOtjaE5w5t20nl1384zY8aWgu1LsGHYif+uCoPcTvtMth+Wzl/y1CwZwlWPLkC
3sc2FB8Hrz6u+HstBAL1EEHt/GHThWe/W1lH/ALUpTwZaVF+HLrY9lfeczscpMp9
5eOTg0skoBE42M63YyOMpWjDLC3cP6zLQwCxx5iY25TeKDvTBkrGJ5Fg09V/iCAf
Q/woDe0kReoxuMdtTvq4a40e5VGQsSpXSGYJa1Gkowxb5DBVNEonY+z2Acx4Ygk8
riclP9PsKF9ZMdFnRRqDJX3MN8R+VRf3X6bo3PS2e95wAkBjxoekuFDQJ5XqlsvM
ekGGwgbnoAnsKjIKUmHuQg8IjpeD1U2pOBQpr381tGA=
`protect END_PROTECTED
