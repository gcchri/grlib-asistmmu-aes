`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIVGGhNIN9BjJWn7rFncaYAs24cye+a0X7bkQeC9JSbNrSojajVzOYrG69VT+O/K
Z3+brwBPc5OvO1hEY+Lt+yiygJDLgfMHIdbkjniCT2KcCWxzErXk/++oN/HAwjhM
AJWnpVLPN8KTnu2iZmsnUyv0fPgISbtiJT/7KN9SQPR6h7E6PFaYuKT9C4A4kdpW
bZceirgUabwILCz8Jkq7lD0RKBTw3H772OOYEdvlIiLgHEZ1cvu+QE+YTGHlRmoD
2P2tS1kfU60SN4QnLt8fuA==
`protect END_PROTECTED
