`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXsIoD4kK1YV513CA++6hRmnplRIrjQiDuHz4yYVP5yB8HMJT8yvW0Sn03hBsH0J
TRC3JgUMwJkrKg/piibSAiDn9I+ezs0ZFORFuNS7siWfg1osCFZSt+eOJNK4I9y/
1Djc2gKtZMStVwCac3Z7jKmSOgU07o7YZD2A6O/LXyIojDtwolRbG3MO6rhQxCUV
2bjbF+cz375z6dhoYcEvHTwoLtyTWId1XK4tGpWclShiROxBBz/E8Nwj7hCrfekh
AD+V+pYPtjlCy59Cn10oUDQesXZ82g5+zdxAvRfWaw5lC76BWGKHCxl3oToV4bWH
MabmJil9Kkx7KMeRvyP6GP/+E6GKHQZz7JNgQHZmCdE+q6DiwO1RWBgxM3gnnpG0
qtngZofrJI2zTnEcIYpmiGhAEtCb/L7IOdNFZYKHREeBjI7UkF9/40OF05ZGyCvY
LVB77RkLcPFbSlcOhadnClsgAxzqp6KPJYnZMUmxrD7CHKgrrFYfZElBPjUtMfAI
ZFTWBvN2WrOr4GN1vNi1msJtpmzN52k5wxDsecMwP8B/2pfjKPIkSXEEJLe3AH2Q
6HaYf9S3w3vHc1Ue+/V60Vj09gFQZcjaLZXpZ9R+oxkHdJJ3iuZ6z4BCtWIgPlkh
z7T9oFpq72OSwiJpQBfijlnkHM/3C0959LVoJ4Cgk0ALa1Zl99kaXD/pzwVn3dVx
hHbw/1COzWTPORzggRgYP6ei+SP0EqpQPWX+JXmaRmRsvaIMi/r/WpAmqXpGx/if
9t+Lw91+EZXBDT2oFYbgGCNGgsLZy6l3RcGKL9GVd539OSUKJ697D1jiwPKLa09W
FhDSWyuPiOv5Qb4RwrWSlCxRaubBRmLRMBYUyrKxaCcXYfxUxcjIQLayLhkKlinW
5Al79x4ackRSitxh2XZiokNM0Qg3PqZ3GyQIiS+WKGdvqskHIvv6BkIa/7ntVifT
j7Y62fAYAe90mYiqm2Yqg+PfT8evpR1nApYFDwzEdIA=
`protect END_PROTECTED
