`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lWUOdUuwVyZYrm5pZrCQE2priuFhZqkYfkw9HcaF+Xg0D8+GmZipc1l3EuQ+/6b8
8PuPdmdqxzsmlVZb3v7Fn1jSGsbOl5AwKJFq3IW/Ya+XxZOEjEWSRx7UZOXIzJfK
bxUn53sw95IMoaoGFo1D6WqcjvMarH5T956HGtVIfNHhKPXxzcHSuk8d+npLDl5Z
IwYU/Z85HsQbz/WxqVzuk7xTyYCHG8hYyJoKqQA3zjcgNvnhwyRSq4noJbszL5p9
NdAvbfC8u9fa1YsP23FAkv5CwHguYY3JSM5GnvllH/4hid+HjktMFxd2yIimyb1u
IM19Ij87pHZ6ODxNya91aR40Vd59TqsuDVLGjJlf6iNSNsJUqvA6pNuaiH+VeeqO
x/r2zDbRTt5Wxvggdmpmlg==
`protect END_PROTECTED
