`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NE3raNNBEIHclCeLzGy9v8WDUUNnCcwuYW3RThCeEQka1Z4Gox/tRUuGXAvUVP3O
q8KPJbiJNtnlHix5t6YFaWwYtrw7dUarllq6hvpKdgVouwSbLpigtpRATof7FNp8
UgkK41F1TZwJwFUefuWSxkyUsgfgeBK/ZdCKhxzOGoei7nK1UnxUMX4Mkev5Ov5S
3POYJaW05KkUj8ec6cDjO22rLHhYqimyl85y/MJA15c1DwPQy8KL/xYZO88sORjC
Y0+ter0bwlHo6FHV9lKiHWojYvq46KEsOAa8dz2Ykit589kz3Sxv8PuYEkFUmPbW
CTFx7+SLwrqaxGJKXhb9lBN2aSx8CNTgn7gymayTXA3eYBkg4I6S/2STbQqqcw/E
8PG0ZO43xxlhUOUNfDON0pHW8f4pU3MnVRTI2btxqkOTlq73QlOkmn53ABcsxStX
sTtTUcUuwJyK33GEnzhMUmfWuDlMY3HwZjM4BMr+beRHKvAf/WJUzqhIjbVwbDPh
K8h2Ti3GOrC1Y1k67Dkj5+CNGlhAXLRovA8WG3sDqRCkQJ1BO6fhVTeNviGd9Kem
+/+Cq6U6zuvm1D/zsh4wnZKG1CxQZzXxnbYMgrL3g4rD9EmX5285L45RCPmFX9JL
3LSFzrnEU/1hInF5MLn5XlVe62OInKlgiAj9NPKvl4bQ7GOLheSx1v5WQhSUOFDw
OOtNnDAriQtEQVhOmhpCET/dpRNzIzcS3DZfXdKrUQP5k0+WnogG9SgzxZ383T/o
vtuaRuY6OZYAWinlbAnjW7H1zQsdq1WkXLNCBM7d01Ov/cKpLUN17n9LGBGeXWM/
K8hlCDUF7SzmHdUuqSJ5yJj71dkunNmD1VUFvGk3MkanIELi0IjWOLy72jrLBenV
S3Fbc1aksNWlKh/Y45ZAcoDm8POOn2pc8MXdM3rIXKDMXgjssvVgeE5jTHee9Xmu
OSWGvs+65vT4qoqaE4OlDXwq4M5ZUKhWU8OCSDcbITpNIDFENGEkMBdlUuc57TuU
QEHIxukzPguZeai/DSeMaeijN5VxZobdOLV28GK8p+x6IqSdJParFfbLJKyvqYmO
xxB3j8s58Ksjw7HLcHrVIfykNSp/HHcMCm60wAD4rF3KNzOoYiKtXrrEBOPi0hCo
URHZna1jlW79Qlvxw0z8LtW/tnEnBKQA/DoNWmvXoakhZ/RNxFYiFL0GDW6jQRme
HfWr2K+k4IY3OSukDTPSl/7pKysdj7WAVfiQiG5DrjklsiSg9YYcYTs0hDrQWKVf
r4GVUcCY1QWUsq3nk14tyyCJo+yXIE9kQBTLaQopJ+XT27Lac3tahj/ZuECG1jJc
A4nwRjxM04MUpYf+C00FxMUaRXVlvkqETRO0C2OY1CQ=
`protect END_PROTECTED
