`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/krjRN7fxWEGyErCDXsud/Pl0vW+TAIJM1LAqPIw9oUMTAkddcyHA+6IQALXAmpt
VF1SYHCD4opxWsejxiQ7oAambF1gplC86TDNru6sJnhiQ4h8ZuPIXuF4vL4pE+jy
uKw3+/FUvsHwjy9fKmfyPhGcfetDRwrU02Sfz8MeA64yoGSSgJ41t0ern3tHDMpy
abRXC0vQMldnr5Ns781Uw0zHtgmdqdGg5mDWFDmTHQhVMTcmVcc5zLA5e/XHIDD4
qx1sRTVNSmjr5Faqa2KjBQhhRfWcYUSS0h1DGu47Lq8=
`protect END_PROTECTED
