`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RawMmwZssSmgIlcbZVkchTbCxW5iq3swSEuGahqbx1wtelbbL3enK90Y1nnjtwnB
1JmRxVJweBbz01kIrjaz59IB9BL08CA9AJjEomb3d9r/rdtwgBIPIFj4hCTQs4mR
pd/p/IWHH8YAZGq+ybUDDQZi77olRwIU0MDcnzw23cdx6XJixlLM93rzgLcyBTdF
Z0nkiS7X9N6gf4EZqj4ukVVyKV8TsgjeAoaTvcw8DWwtpUuj6gqpUol2dt/JkEmP
hbj078Oi2Uif1AF40De2OcDg+H+ZuH7B9KmzVFNEz/6XYlEdQYj8ygI+t+ub0zWD
7yJWWcQ19sgMKMr8Y1s17vjAIZ1Ci6n8Psg31Jfj4rKUp957m5lN7NyI2DOwR3pu
cXr7elkQvcLe8Fdn88j9hllWfmj29o2KsAi4UFrbWdVuu+CG/ttaADThLh+6qMEM
7qvhCy4ThGleYXwagznEywoH2wv/8QcV1XstddzLk1zWwkAiXBot6YViEWmVLIDd
xTisy/8iEiSAUhivjicyQppBq0Uu8l8MphiTLFM0HHY=
`protect END_PROTECTED
