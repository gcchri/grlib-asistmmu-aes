`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g3LAsqtO1162bEhw8Gd2UN7B3Fev/UhVcK7JJNJM4uCJFpybm8nMxSGptHlsHdyE
dPCvZO8xn1MfTTISylrvgutP8Zru1OE5uGRH9e00+EanN4xrLt7ekx30JQIi1/8h
xK0tMwKuClQOccsO6B3QA5VhbopG2MF8cZvtxufZ50WPci5EOmhx/GJvpcMxY57X
fJVv7G7apOwfEUvQFHB2gsCa67Me6abaAtgRZzfAneA9OQgf1P8ovoJz5iFAgqQQ
WCRAiIzGF6MBAbBCIMnnI0rA/fza+6hhn7Dt0moqwqUnxGkeRDzycW8blJJTqs0C
kPOsoodcIOdzztOVYQknDUJFwSutvvRjLSvzlRGCDxKUzXMmaUk2/BGtqm7eGNme
srWXzg4erF6QweU04ZoEbeKqqM/RdHoZOjHFyrrDYAjeSq/CvPmN4ylaOrqiBHUN
sbLY3EaEAh24V+xqXU5+OnoS8kwjHYLDYnDzSlXFQwUOjojTOe+RZIQkw8nVYdXY
ePHBaBMjOwTZbKvHlXf8xJT6oWuNRNMbGTp+ECm9BcRaaFILLXnJEBmXI1rlArVi
xRy9v+VmVWCbHnBx0c5zZatOdynusw4fQZNKVR93AKyy9MuT0IPpiUqTpr7HQWZW
h2F301wCiCBxFEdhVXnHQuMA45vA6BQFY94p11GCAGmXJof1s8duUWbB9jvwp5zn
UcHzCN9FF5KZmiYpRDOr3dkZC8jekKDJqa4fMKjfmKdIQ1UjpqAoKTkJI/jm/iXh
R2O02gLQn7ssekQXfqCyudXmPgDjjVgt6//+AMbwxW4=
`protect END_PROTECTED
