`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLt1gXvnvl4LlDXMNxovb49mNOXiKGMt6FpuoP41nNcJb4Kh+stJZJ0LrRH8o6d3
qObz7IHvO8DNd8v4WL9HYlx2PxHGTcdpz84NZNtxjK5v/elTS4X6Qqas8WRwlGyL
WPKsamk6p1AHrqvpCptFPYM+BOwVeyIzphFVU0vxZwajuXD2i+hhv4vyt0BZLFP2
lKQw5MhN9gF03Ew9aKknz867/oN33nAIFc67j4IX/C1SeiteIlEkXCFFP3s5eNcI
byavJxZ3Ddo+/P/++PLF9QyFOWzprt4hY7Qm8PQWm1iz6S2lNzFRxW2SrClv+I3a
NeBqFbeKyn7vyqlfSaNVBVQcPrMpFOpjjeDfixZUM01PC8dYk31ILyta82eVC9j9
Afhkpz1BTO3z5pqvOtJMivjxdvMy1iuk4JrXmJJfjLZtw9pj2TFLmAr/XfC25XIw
YlKhcjsiIuALtJdvnTU75mA2XQdaczvhpsdAUMD8pHxdnxMErU2WWIwUL532n+S5
vr8iIFfGy2Awppcj+DOUg5e9m1jDLPAlh2LRoPIFba2K7fiZr/OvhNOsYLmXr/rA
`protect END_PROTECTED
