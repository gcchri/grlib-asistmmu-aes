`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INmEBF96SEwfjvbfdHgIYhx9GuBxF/vJAdU8Eo37sioRj9KdGglbsVYs0mYMd3XT
Zp3veAfhtDBFsgR85jJJMrrA++ym0hU+F/TFNYbUpnvQFcKUqut9HsaCupYrlf1b
P8rEAPF0zpK7anL/pzCKIP4anj7fpQKc0/SG8E19F1FcDyYfUkHKd35iETa1N1wG
WwgYAh/zny2m4vaVmxrVtm7jJGwzj7TurC3WUDYxak74vcw5kPb+scTiDu/nrQfH
Y/XQl8psAbriSz/E2UPW0YuU3+nPKssAKx4II7OXCsOdyqqhZGi4TRRBgZNRamEi
DqNMUX+SWBvIfJu6/WvDCzgvGnUlX0/KYa+1stpiVHcftFw7wdhPI0BtECD3EjCP
sQw05eXni4Nac2vY12mDH0MNBVrQ1Yp0R7AllcX7C6qKsUyAidAeIa4tSSVq4jOt
1AImQc1eMw0D//naHO+m0ZGElJHWX7PwFvkvMqcvw4oT/A9beJRsueO9v4GdDqj1
WTbkiqBzU7OdlEtWujzBLn09rVLzSPSrRXINrtenKMJT80cYiHx1APBE2xQOxk6f
5sW02Qqj5qTyE0p2nrrhzKQHBeuj+m67FjBkybPNqjL78wG+WM3AgLN9iogvGDYH
5lULBj3SCIzWPi1kDwh7M2It8R/6u2Bk3MwvCy+QplqmDF6TTkKvRKzBff1V8uhh
biRxQYXqyAwXOY/LRZM1h0mi5tbMsINDOjulA8MVXLz+gpt5GWV5Pgrk/xBopZw2
bnT53YikHVQFsYVmHLYGzdcxOysELLZKs9ri6/O3Z8fvDNuxyhdDXesOJG5p3ebl
wrEcXiijOWEbQ6a81NuqoQ==
`protect END_PROTECTED
