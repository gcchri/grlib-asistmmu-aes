`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4edduL1AtTonhIbFvvmxnjXjzzRxCUJ+KiZSEgimfrmJtnVJalTK5/LgirbYWQSn
yaV4LS4Tur21Zr9ew3kX4iXluW3DGrgbqFKg4qfKWyZNPWjmyHNjBKgYbT+EXjaL
WpZVkRCuNjl7VfUJ3faxUNidlPRvsczIZAs+N5e0fQinFhnK7/BREbukaPlreySx
VXxxNqFZNnALuyaNapmNVOn6DjcQSFhaCrqB/Zqmps/9AAUsvmSL9mDhmA0hd5gg
gT7nQISh5TbrSVestoTrCMYYxUsZY3JCDDRe91Pnc3+OB/3h7am/cvYK6ki1kZqs
e6EfEOFPmj2JoeA3EZybsZtYA4qFl8KcPeuW9U6ToPWaBQNshxMMOR+/sYd4mbEr
dduYfPSYjgySN3ubW4PTLCTJmT0ATHYMg0tQJQ/36kM9JcUiXDL1VdLooREmm2/w
G1Z/8OV7siWQZrStE2rfajull6+yYVh2waQx18PGAXFaKkEJ2qPCcrbZA/ryfwAN
lUrXEAoNA67UNltalN64ywBZGy+eZKteBbblAPjZXtYap2qPRnKKjbAsRtvuWC9J
7kM80GdyuZ/o5gTu0WyS/5th7J3/kPCgD0U7jaaMZwV27QqyEaBEmfICMa1WSydI
3z0BRiPoBiaecwOTdFrSZKDe+vY1rxResn0zAr1hf1XsABzRSrniAMrTLSKloV/6
FXV3sz85AMw8hjh9RO8IpH6jNkLYoU+0nmhk70sBzetLta6UtGmHyoyFMvTiQl+u
xTBAvTuPve/VvLOpFRmN8o2J4SPtTnHgqxC2PIM8S/6CsDuMOxp6cS7HDTEnOiKV
fz1mAiifFYgJpX+uzLmpsTmiTEumhvJHt9W259OBK4DBbLlXhWc57XxZz5ACGrna
P1nvvO1jLyylk9WTwC+lOJoAMvjlYegNcW6+f9fHZfqR/OF8jI9gnUyR+7y8t+rs
JKIAa2oHbHbOjzed8XQ9tdcg7/k1vYc3dCYuSiGkkRO8IKQs3HDiLOMe1hQETjzj
Lk+57bQIchapsNNH67eS6tTZgdQgJYOt9fDJfxtlm+cK2MqdqiPOGWrvKFbHVgas
LVxv5d5ke1X48BShCseUAJ07NmlGAuox1EBJ6SeXLP1rzr3vNzWAfQXlPpVgGykU
Uq7eDSm8UwYh7D5FyuR7MTVFQJ/WmnDasWdk2Rb2Rzlvrav7vKF4KnJH/slUvRJZ
gILk9bvsabbsU1SF8H9Zva5HSV8jxjfXcLEjWEvjEc8DgK+djeY/AuWNNt4rK86I
tn2exXOKLqK3kXcC/TAwFq5Tx/IS2GmNxU5mJyfhmMZlZm9r1M58m+hBWFPHWofe
4cnUtGeHEAxKairYxH7G13n7lccJ6DCq4/zHKDddanpWdmJV8rJ3NnST63K7ph8V
XbhODXr9H4qhxVCpKzjx+9hVl44BdO+gduadhjAIG7oO5++8/s/CPLrWzWPMD3i6
xaREqArRxVWUmxhprAXT+seTiN6tP9n8MY7RNBVwb3XxuaUJ5IO/ALCGC41mAvNJ
bbByPAK6ZVbDpd+xu+u0adTgafEtY1aLU7ZAMSaw9XptaXoAruiD4yrmZj9K3uD6
4Nsku+Cg5dTOK8I8aabclZCE8ff9Z9pFZFPb92icRh/3qZTAqEvzerWbVgarFTks
HH2yvEkxQPY+DC3/f4itg1Doy4jo3on5iZKVIZRbANKpa002cuIeMBTxrPQO70DZ
BtEBpDUhHNmNpP4mS8clWVtGGma5yRIJA8LXKCy6w9m+BDM8Ya7ECNjLmxOYosOH
r7u4BV1KP2gabrQ3AoLPYvRu0qF/B8EFtWNUeBaplop1MKa4tttVgsJmMWMKjuuX
ibGFidfudXzVh5PyzhAXVFRXYggcUj8htRU8OdOssQuthotQrJXkftCz55e7U7qP
4KVaFNp9MniPVbwU+K+rfHTMFGTAOX9/gL+n7s0F/+VwkrIVuliZ3qVcQTpeAkhh
06tMXWwmtySdBIKdqWClsmoCeuNyz+3xm+ZE+Qy8LYeVEP4q1eSM5siTj8A4bnyC
4fnWkQEEex4eoReP3ftTc4H9anayY9kb5i4HSlOLb1F2HlHAx8cvYr5k4ElZp1Va
Xrw/KtUXX02fX6J/x9DEnLqna/ZG2rsh1hvbcfMT5rRBQaBnHLUn0yvbIS+8sHAB
pZbHIJJTY30u/fsNffR0EVljFdrIeWu2lUjSRTxh2fCmANR8Yfm6flJAPTZIwqi3
5eY3IJNTwZ6mWDiF0VwwK/RD3eTW5fPVxwJEh3TQOTE364PMWCLJXCE4+Pv1iXCf
reiz56KWHVz8LgQIifuuQ25sEupBRHKFD3EHlBloyUzEsixXFiOOS6+Tb+KNWMds
YpLS+sMIcBH9pmN5aUDDSaSyrOUN/VCZJCoT15NtlNupxdl2z3vUPrWi8plaw03x
r3agpSSlgKNUBoQMCxb42Klvh8neQAU+ZtBJwT0kkBP6ovqCQ0wgXGqOB+piEA2X
p2781I/7JE7ewODNHm3BQxbbTU8AeDLvDjRRRPfInqk0tIIYq8Q9yu4ww8U9RQdk
1jK9QuM0o17gwIlo18aoP7LiXSf4HGUbjwQdW8wIA5y60a7VipI92uoUPphO2onC
a5rwukpKVhq3scMbvkrspF2MoOoYOSTRcRpR1FscIagme0chV5LlrDBImc7R30kM
HtWQ1VfUsRXCCJDOKgGXNRSNiLlQpyKtecdhEbK9Zek4dBcUnlUHJ766jvMW8IsX
FOKFgLSoz3gR/PqAd0FSYL+XNVtaXI1RkQTdkAakDDtw7kpoqug3ibXiPvYj+La0
jhlLhrxBi8gs9+WXva01ESEIAccZqJPJkcAzGQmLLW6WOylP6JGS6n+EuQBffJKu
eI+oEQmv357zOn5u+2GvAYBF/VMNxzVl4gZAbceIPBl2kEzAYDtImHAC9FCpk2VV
enK32JT7Tdqfs8ktFKluVZM5ZTnQiBo4UMHitNMQuYdoiIWw0cxuBCZzEQsnR66D
dh/mjm8ksVl/hN+q8L56SqPzomZilbTl7eifSbvkvmjZ8sax0w5Onkvcxh8D0KsI
ojxmYwNXAuNGsTbMm7xqlm9HbdK+zS/kse3ZccVy6jaXOEu3YF1p83XQSLfineSE
4SGknENz0QblGA3bEfX+OnyYXiVPAysXrmyQ7WXrbjG0M8rm1yjmTmsYrS1RC8L2
Cw01QkkKtex6um1Ht2+C6L1jmKobVZIg044ozbIb8iQHlKWTVvZ+R4WfMjTDVJjp
bq7hIxGA25rhbQZbhGK3ahlu1fgNgAzcH5o89mkKQsQ7w0beLKv4Jl+pH3Umnm8z
wbSviUBMEl+lYFUVnf+OKRjQqDW8rlHqCJaskZ5XVNBCVbcoPbloKQ2+h8MNZcPm
vtBeesduZyUzeU7RIefiT/CsKykURRhceFe+a4/x2yCci8MmebA6wfwntD0z7GXt
RjMcfWqiMRIWlBZIktVZbFqoR416mnEr3YqmbfgE+7AG5ANPUTetKjDIizrw4oDn
eeZbpK8DpTJ3wrvwl/jTE3+f1kC9wyUY1iWlnBIxOysy4zMmwCvCabXnGBRrVRW8
yEJZ2tmS0gJBiVqTDOgdNwzNl8nVm5lv8QnrBk+yvclXM5fU50KgU9U1npdvPOmK
tolas905LLyUc+pGXm8JcGjN/GOsS4MlLc51OgiZgrDr2bT2ZCUFeRLmuMBV4Q3s
/jIyGhQRs2lyVL/PTazwMzwPa+0ap+e7bajxhyHQo6vDW08cQ3IeNdArA86H0+5I
q5+M6gNAuLMOFelNvsvRbpjTzwQDg1Lv/eFAwqkJn61etw2oP2/ohpZ+idPJTIGB
J3WzWkAYXOzmVkJOtD/CzDOXvD3wZpCqUXCRsbyCI5WbzshvMuGsat8CV4pbEv82
eicqZj0OMRpBvSHyZ/ZsgB2H/NH+YRuVOB+zBhyYIe2m+AnIzRLJ9QI/VHNiuShn
fVoFoPgcXLp6gl9OVnMyyOFoSyNnu8j7PT4Y1xdh9ayrBSHBoM3aAex0OQPMPpYt
NQF5lRzH/R8+DlEK6/46QJhNR+knpTLgMr3UVDO8EhB+oslwx0LaH3qD1xR0rZFY
EqmSRDbHyENQz3nyDBF1ZyY2HJb+CoNwt1IG41mU2U6mYG0MkNhzXzG9uIoLqIXb
`protect END_PROTECTED
