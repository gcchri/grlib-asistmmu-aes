`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbrHI0w6nClXDkcaSUqGAxTfLZHiBN+AUHJX6Ti4rr164b/MVYq7ZvMuGo3r866Q
AjrnDWk2JFRVrl3G9IYJoU5SXqu3F/NpsokuWt5t6y8TPnrPrjS0AkD6Gt9jPPHo
Nyur8HaJCNVQXJCkyoZd4LVQUYsHo1x2T49mhH396Bx+sYM012lehEq6he30KTCb
gQJjUJjQwKLl/V2XxAd1FJvIIuE9rXE3b8QX7Ek6gOmK+PY6xo+VfPidtSC0PvZ9
0d81fcfyig3iibvLVfsmWA==
`protect END_PROTECTED
