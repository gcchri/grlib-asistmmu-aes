`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UenY3xS4jdEi/an3MyoTFN3oaZmdEB7HadtoEXA8I9u94Ra8sw7emb7uTvyWhXje
zqaOm/IldiPDnPPz1pz6l2nTMKQftUsHNVYHPi7tcOp6XTgo2p9yY8EAWevKOKOj
pO0ewNaSpk7TP1X3VUtvys3B+WyQDBJBwQTJ+IKmTi5J+IEqYOF3tShYgBI8Im5g
+poh1V5jLPv5tV5N9/GxaG2qpE/QnMu5RsjIbIZMfNtqJ0WFSEq/xmWfpOVX7KFi
hW4OkiBSeNk1JZptFFByX24N0SMIjEyR9rCVu9C31aRhemTs9hVq97eaKNzzhrXU
84lgsATObgY1boVpFfj4o809W0h1gy5pftmOgWJTTZfXU4jLWlOAWc2BFvcmsGLB
UBKFfu2JpWE0TvKwG/dRN5Ojs+8o1hL7b8e/c5Q/pzraCHibuOvpGvuY7Yx2aJy1
V7IhUP/Vmla8JFrb3u+kvaDtRa377YCzAn1Vg+ig9mivzdY9A5ytNG/jy5ulX4HL
SNBIvz4+V7+6NcNpDJniNt/MeUQqIp/cgS6iv+9u0mX/uDMt00obD5KtOxvg01DW
fnXlnnJz2FcXaD+HX7+53DNpc13zs6l5PdkZbGRSvTt3jd7kLVMVLqGLleHQ2p7c
/rIdLZMdoE0L8yWhV2qZfX+S1BJoMs4rE7zbeJF/etI=
`protect END_PROTECTED
