`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2oaXAvAH0L1xK5Ehe99APHzoexnIBjnyl9C+jCWAy+smDdw+oliTnFCNuDJhNTx
jof7s7aqZSCG/5jUJYXJlstdDx6pE6zcTqoFubul1L+1RiiYH29G70jClW8BcKcQ
DQMBDx49/p3QzEgFnNOCF6yI5jso1lYqryjXXsNGB1v7xFk2zC/gin+Y+hP+Vlvn
gbIycnZfzyeoPQbN4rUIktRbYgpO8aSv9HqjXlO6IytSQrYdC1+RBQPtnhTK5tVJ
T//VZFAn+i4wPA/m1FLSjSCrHq61tRojHODsOrk5fbGtFralvSshQ+a8K8JVrUM+
B6UbmQTg+6famAx78QzvNtjxpAq3MlsyvEp81s6FTrJPi3L/o/N7FTP4P1Tql8j+
CVfQTb7LuBgfGaOE0AmBd6qQ+tFzpkc3ACwNGXGurp4ODHouvnH28r2iPdJRfjlp
/azpkr1zzUHF019XSzfUk57jZISLqPkMQ9h4dOOdRY3TpYlDXD/iv98DggHtCvjr
wiLR3dxtyN+YmvHQvK9IDhxbvJ+kEY0rfA+FMekfavzGSUf08F/Oa+wn6AAhkY4L
3yyEALPCstypAVaz+awBgw==
`protect END_PROTECTED
