`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dY5O/Dw/4qcXsagRaiWGvzUTD2MqYCpzuPD5hj81kAHThOxgHpR8jFIEsGjhBaiI
/MX7eeuJb65D7Ddv6vAmkwiSI4p5p1k+nEZMQf9l4VZ/l/8KdnbcpGoglFvqUFPz
mSSR7+G1SKUuSB8Mkn2L92Jfjr0hcrhLAGZomS55VrB8YChFe9uTUuWyFCk5xxYS
eh6pT+Y5Ef+fkxGxlF5boHVtHz6Vzkfky6ocUB4HkGteVSLXS92y5p2IomFi0Kzv
xCDXrm8xg24mCDB3DlJXvkQhjDQWj39VWA2hYEV164dl56WEzIh7sjVJzXkcH7nS
9mINLjmRnThbRaHCL549mw==
`protect END_PROTECTED
