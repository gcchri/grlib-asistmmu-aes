`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0YxgE0ABbjARPFdKzflKsWGwD0EeV54J11D3vjiUcgVV6j6rAWflZoLT0nm1ZVkX
/Q9UPngeGDoq2VX5XAxvc63LBoY3E4+NnK5uyxtErNa8n9ZsT1lFHOsepGLhxUvC
T6RWqrE4A6W4KIZUmdTQ1Xx+HL3JsbJgBljWlWyiS1WSoZuu7hTFDZYPo1znYWEZ
jSPFrwdYcyWRpZEILlH6KgwcqUL4gWGgvH9fufcDM7w8duwLxx32kZwsmg+LO7ph
sODCbUPRk8BlPSn5/Q2Hwg==
`protect END_PROTECTED
