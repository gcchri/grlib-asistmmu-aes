`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tqPs7T3TXEii1sR1Hr6/r/HjelTJt3JJUbpceTU+7QiKVC1f8aW4Di4sof3zq0wI
CD+c3RKNszBjruB2hQXzMFLHu6mvy718DIQjbe82Xy2TnT+3L1LV/QBR7dY5FxhV
/4Buli7iRCpjsOg4a2Cgv+QMaKuhhfz3OflNz2HdDpprrUd+zHFP+PDHRqJDA+9l
zx1bQhRQxraSdciIT+vTuEIsWC9IpKWpKIQhIdBeXHkvx3nwLkAHwBJQA+TDjhhC
tsHVLm6rBBImBoQU1kj4sAfpC2X+dT4eN0du/tzdxG0++qS1dBynud38Agrb7TrO
jhNSHbMtr6SIakBvpSsh1w==
`protect END_PROTECTED
