`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3H9STuN8xij9ah4DHl86fJItkfqNOuutqTO5NUWtgWd9/KDycyHpz9V6NfZ6aOfT
aWwH7/NOAxv+GiQJs1qcdTaEEKqRfHg9XD6XDkFYrnDPLNZ2USAqgqQ5jPo0yuGg
hV39HzKz3zx6WqgdQBIHLlGvh++KsS/oHvSgjcowbo61xcsYCcYPi68/hCZYIfch
rpN06hrbaX7YYXnH5klwHGsjymVdysavH53Fr+6CMJC/VrevR192ecUHdy081vvs
hkVy7VsGFX5dEsRF0qnQ5zsDfa0Ro6ppEjd0Yf06wQ5PGTOg59aUJYnUTKimMaT1
vudLjwPomvsw1c2BfOVBJ2/6ggwlQfRJrLkb3N6hoCkjRTP9IY0Tby/t62CafI8T
pCpm7A50PHnFz0m4ZaLL7zeT3zrOCceeFlFS/8TlkcjlbfSBTu6fbsLbplTE3MzD
8MxQqX3cuWRyRKdcVTKqJwIE/jsDAXAqCyNpPS1FPXe0scNorsi7GrT6MNVVqdhQ
72FDKFalC5bGWx1+NkRCPQiLs4q8tUp4QkjSeIifrOKuenAu+/HiZX+1fIRGUMhC
DX1+brJpf958QgmEP3V+lhpIvi8nH0uEsku1rH3iPIPcbnd4JXUFVn/SmbAfwMKU
tNHb0AStsyl3ffxwxlT0jPCOXLQS+594kgLQ4pCqLVWp+8RW4LA2acSI3xj2cAj8
fk3+my0Lmhxp9WRRbpf/NPOoiZ53TAl3g1caY0vIGIi10QtzXsbtaSaJgEJjmamI
zpM0bo3k9nqlbnmFuVZRYwHsQma6vlgJuBoN90A+qaYwaGgNzCV6DNCCf7CqX0cz
Zl1fYeqrgJ9nG/AyLLAJinY6u4blNgDsA/y5ChWaC8hvfn7VyRcb4YZXIMqMoY6m
+djapdsYolwKRLi7TlgLDwPWHMYCZV3jv/Rmc91R93k5u3SrAAswg09B0tpNkvke
rr/drspNkkZQv7gS98xN+eEo0w36KbRj1aJRaOyyenlAX/7Yzc0rkK62641YBA1F
qyYEYI95UTaBvq7bmQ9Zg34ZgJxZlfTk/JWerB9GT9PIAnsJidBweDtoapOkZB2p
vIBQ9+ID3q5VqWueFFZR9PoITyw0JNkkY6UYS+KCij5H1Ej2X5QyyCvF09CaNK08
VlXb19uNlq0bfeN0xikWATA5fUg+wNbVuIJCM6jQC0+GXtFSGzilPwPxcEsovxj/
rvq231458voLJgt2U8pAZhbdaSy5x04mOAtL/urXfBp0c4BRL0H6KUzTDT9nQbZc
I3jhrI0bWYWwjRuVyiMULY6R1MgQVFY0BEu8QDW4q/O7LU8l+CXDLCAfYLxir7ph
mkzrBfnC+si1XoaZPTCn6BmQJ4p3OtWn+88SF1iAyJwQRFTuWVXwnHldOXyA2Vv7
9V1r2eJ9ru3u0UPUtCM8Z3DvCFvbqflGJMf01dp4IWD2NqsMeaDIzTxOexA1C55v
pbLlyL35zx1dJUSMdI5PiPtwbWg9C6YMkVx9rwguMQwCxsq07n9riaRGU+LXz+SC
/rhoq6EluEqf0ssV9R27OhHA5YrZEVtrG+nXVHZDlbXBQ48yM3wW5QxJWm77ZWLi
o/ZvmCL2hwjLpdoTasELqCypS7FN7SRb84Pa5PWMoe/4MB0AKEgb6g+SBXhwFZYR
iFW4/n/5UyU2nGIJRF0LarQmyjFWizu5zlUdqJhjgunVfbdNIq7MoMQWK3zfmK7q
5Ti7+Xb7B+I4duflcY/OejY7enu7c/Vwj48dJjqGQLJNCZiDtECAC4fJS7LNAOOV
0okippzU5zYIot9VCIn/2ryvnKHevOf3SnDinM78idUej8zq2kTfMAXTZ71xZLD6
/orKKcdZfi6whtaXssgr/bTl9O72OA0ygngGQNOt1mWfr2K7N0D2n7I8oVgK22Qf
iS4lP8eWjZOZ+ZN9Z2vtqL0VOEXjjSkhwUMzkEYtX+Q2EnOYbkhd4UfaABElLh8c
HApHJwrPLew8sUhgWSaTEcrlDF2eV9Fxyzv6jfiZtOmWRVAEx52RMSniPHZQ0yw8
2R/b0og2m3UTNIlfOuYpYSBUjl3nabx4xzs3MZwEHOdzkqnpmSed/onS+n5ZV0t+
SBGrl7k0aYFrl7/vrwoxKZf8JiU6huO6naG9AJVANC8VLZJ7JDIQU7yfnEw2RBW6
NHAsTxKakPh7udN9P/B75mxckmnZkXtU3fWjKOS5Ky3h2QcA0yk/JKmwsIA4jPYG
igYtcvKxqiVRa2CQhK7XGAtnUi2rYAaLsu0mznBArM5dc9fE8P03vxJkR13jXwB9
q8YE0FoE4pmbvEM3SH2lb2vHidirZ8rZolIjDu2Dtjh4464TSOBY3uMBdufaK6xP
/Owpzb7kqY1mDN/NhswAnXeAwfJ7DhWGNOq1A5RkAgyy6VEaTCzbck0QQW4QVEYO
TbaDMENNVzvXoj/ANH14JjAvC8QewJIr9hFKACwLJE5ndgWbQ8+tuNNlTLUuCczA
yTEntG7c+vUs+47aeTVRuRySIFXYCq6F5wloXhnJa9FaDNsDC+wzMmCYmkjEuTdF
o3W1ksfd3gmP4mH2/mA4+A0LuL1ujWvQWgFy0ZaI1yg90uz6oPtc70fTeI9qDU+S
OA7YKDSZz702dxzm/MSDPEziWgT21XM2C9iDEu+xM8ePM672Z2K4gbFaxEU5LR8M
qSKlgn3dEu7c4ZbadF7dEdH872IC7/uek4VRGx6MGyJNUA1ncKHDG7AClSDk8u47
RGE75FN2FrZCIDpVDNOJfctal9zzK27RXpZBrvSq/0M5V+DEWHi1HH+xk8+Etk7K
rIfibYFaARKCqljYSkPfE1vr3iYgM4vP1ZXLCgj5Tpp+7uaQ19aJCnrPxhpeuMN/
98uM2E9ZIDW/UjuBMB0B81r99BGfnldGrmxVqzquOt3NKpEcVhmQ2A8aex/5NRhA
JbK/gpCe+3nJ4WE/WkNumMwxxjTo6Uei57IcJ4LUxTimX26WAnUPa+kJYvcRByfN
MtkaAvwnLLd0ovCCCStUW9F+kCrcvQKjK6k6AvjDUH8moUP6Wq6jW95UOSsLS7rz
B2e7w0GrMx/W1VGWhWVg/mafnmTFOdl09U9zQuDwTokCSNz7478wgjaOqpup9BAA
kviLNgqhBnxbcLLRAFAerSBJzhET5wOVwbQ2IH7vKYRLsn0OWdzeZRtqX0uiLOZd
qTSnA+Q3A+mzWWnBdGvmqskwF04RXSqs3mEPOzjOAcrdbjQEiRLKpPFQxYifnWYp
D9Svld6ukTUaGeK+dUGcmj41XBmQRVNP/H9tb268P567hMgxyheFryAhHt5JI0Dr
wUSWBHlAA456MaZV0pGBbUSrV0tG+S6q6wUdjP3WkLqWkM4fbZMBtXXQ1VoDb6lw
nRSXiMBIxRqxTk4QGiLD4KgMaAu+HibgseMjPfN8HY7C5YEtvDD5UvpRsC2ohdlu
vm11N5ZJo5WyW78Re6yrdpSuFy00zN+QGN4Wes+yocugyp9htSsgdIVRCmuCrHgu
UNBjzQtccvPuD78oySnEVMcF+V5QtPAJ3rhn/CwZH32D8Oj+qQd81vqlqt30vQpu
fZAm1zYAAqWryMGB9+Mao6cXGtcJXaQl9zMx/OOizK454ijgH6KVVTd92NkL4Lbr
2aB8gcmrtXOWIEsGFV1ZCHEdEHJiSISALn0sNBxMa7GDxIJ4JX/1Md+agjd9+rQc
J3LLrwyAAupTL7BOdUKkLUn6bBjxE6pZH7XkNKRO+6hEg7JTZH9xzgPp3fFeoP/4
qy2pep/Jp+asiHMEG+CkGEEINN6k2PlDpKJnmBaMn7jWG+BxWhBIG+LyCwJc0kye
c08Nvt4n5droeuOnzCizo8Pm7fCraGVFAMNCacHSlvuZYqfIFLIQHbHi4fp8Hss8
JCIUgtZ2t0ybtfgw9AAdy1c9c8o60iYW71r6Th45BrVeXYjnymQqRv+VQcCaejAS
b6YU7vJ5YatR9jOL+N5km5uQRwppJDgxWUjXdl/iQwAdaiIJ5j7WpUQhcMlIc/Xr
moXLPe5eAoh4NfqfIvFtSzNDBlcWW7IfW3eMe8XmoBvNDdXtT3BLZvSRchYYZFIk
fBm1sotqvvbm/LR5xdAOrg1I7K5C3PwMSpTmH1WUx3nIbRuvuKYbFyBABoXsm0ti
rlzAsY3efLcqOvHWlO+EDIR5QYZzXahE9oUygLdIIbLTwsSu0dIHqCSQHolQfvcv
2c8V9qomWEmnvBfrSldnVRW/fk8rcMj3DoiQ9M2hTPecurxV1Ycex57c3j0tpLfa
Dk/k8VNe3M5KHXbBd1s74BREJhQuIcqY8/fDSiXum0SyyynqjZQOV/DWaS2Mis2/
aZ8Q50Yo1JJZwJWXGgaWjwl19dCwKQ/9m7E83pEHIPPZbo2xtQnVgpja8jciZsFT
hIbxsYMtE9qSuR/8vx/5SCawndjQcEtWIBLFTzdTgCRlv8I1DhFcZDrrvSTtZAZT
U9Wxpzd8olIey1PDSqrj+LrYJ3pVMw0jOtQK8V0R8pYTeBxayj+sRN2A6uFQ1KY9
k6ZCvBsWIS4PCQmzYs6GmnoBd/fqo6VaKNtLNq7JjbHgwdbtuCtyfjvWfBQDsH6Q
hr30ry0e81lBm8klkC2PdWgXGaMjZupPVkfHyZ4KbhozvX9Lu3bDsq2csr2dLYf6
FsGeYoqUWCxzRbSiiX+OhgK6S3xmbFfK5MmtDbq2IjwNcG+OQ7XvUlLlFHGDEvEa
RP8PKwpECE3Le3/oZgVF/o0D1OJoI0QXqdwI2wTtgrVetaPuSp+ahYQkygdsCZ31
ZYXq7XGuAWmgPk3EGA/Lw+quaYitnhEQeN1waYdR4Ja5s2OaWJsZ9WkEjxDgnCTB
XIioAcl58SDd+7SHUCXQM4bJ9sEdVsUfPo3PkKkbVvXBr4h8WEhhTCwYjEqvpK8f
U7oN/+aDhzn9jwmzz3QNnIcSMdokLtPAecV7OkE5TFiJ+EhRYNGzkf/qS3E2y/q6
ohxpxPN/YukxgXISubT7Q0P5ftPRf4H+4Jip6hpkMzaqg/o86H9knz4fOLiG+ESE
QdIZ84jn1NMTob77NKwQyorh/PzlXw6xCeUZVz7o0+TeA+/L0B5nq7ZVDLdvlKQQ
DhJ4YfbjLp+Ro1XFS3WzU2JCe6yvtMaH4Pd59eU/9NWrPDaCGP05Tam9nx7h2U+o
Q6c5fO5yBXy3hrTf9qLYVCztp7MZhRDAj+E/GlJbDIoupPOjIP/InSYInpKjgfpA
t7lIBiZRISOSzeb3RKWSLqqOXgMJ3qrjEasMONxin4GxDkUt+1sOuR/xEqq/mUn/
Dcp+zx0PVYpKHjd8EqE7/Vq2RPIc+XWPz8WLZFoAVvI7zNAC1TEdd3gByh93hRVf
B0F538wZGE6WdihAvwkkGxooI9biTJX6txa+XYJ5R3RfkQDyUr9fCGvZvFVXE1Re
`protect END_PROTECTED
