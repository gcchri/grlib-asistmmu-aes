`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fm6MhwSVBN/EdPWJ4xn28ZjJrQbWMGcQw9w51GjxQfxAkJcR3MnmfaYKRU2YkIWZ
DclA4e2rX8WePp/pFLUdptBGuZg+Omi3RCd3S5MffSrjKQ14alU8UBeUv4Gdxtj9
MaimC8QRJgK6B4BtqcEhOYMwKWxvGIBBdl+fExIgs395NDbALgeILQ9yXnsGjC4C
n07aCYpiRlrAGjJMGSoltwHLsWWRQtkM5A7rAsZmCuFwC1g9YCzqADGb//NzkiYa
A3qxsZn43mtm+K3ib2y7qoKlnxHC52q4WzTKF3XM8Bp1dk6MSL6QUT2r+ntw/tBt
pwy0ymc5dg7UDc1SlbLliwgfSZhsF3CHhHYeWN9Qw9TUDKRFGq8My49xBkWzdgZZ
Q3kfDrIg6bxGxFk1ejQhvA==
`protect END_PROTECTED
