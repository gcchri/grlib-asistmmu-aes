`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sF9LBoiMRTdPxUhC3M9IY38poifBGoNNOASLlvOfcoNtyTkcfsvpy9vXHlNMPTZK
UpJfH0WorWmhnFLVcd9K8lBKjeqV4CRBTryqbg5I9DZBxNfovT3y+MuPYapnYXod
AgjGPr11O/4hPtE/Pp+iIrF2JPbswUslnTl0uysdViM2dQ3Q8HDtcAjK4AIue2I1
Bd+1mnz3NjFNbbKFUjGGHoK47xNLfPVu8K8VdoswnQknHAx1TmYSmhUbrxWI26Uf
00JrfEwy5cpmPSRPxDTvp9xGXmrzEG3Z916imgpZj98o8UDE73qyBSj2JEIf61Yi
9c4ZrQcCjEIBtlNUklgbRcHkvy+vCQWEw7jzgGwVHNflo+hNhpb+Th/5BJFSHqCa
k9S2HDxaKtI92NeBwr3/2y8xI1RqyRhCsdiFs2gBgdrDhO+UZ+ezPtpFZM3ehZZ/
5uad5QjByG1XUnKA9SJpBV19y+VmSQ0xtPcGtXWO+BEA8MGJS3dqhErlhuiJ5n+l
1A17IROeSHT+ON6X4nBhboG4Avl6Nc1zauOCwOiA5sw=
`protect END_PROTECTED
