`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/dPDJufKNnx5JIgJifbZud3+5QXzuTA3PYVJ1+3tYNA4nSFdzyt7HKxUfD7rRiE3
tqwD7DnyCjWodsEb+5BaLlPx2mhvm9pG5ReZO8uVlijuu4sp30Kovqqz6vzYKFnv
1rjl5FHZor1EzDN3OkaLGY91qqIJ68kHbJm3RiVDV/xYFz2ptPUz74646ZNznm3u
UX+6ZX08lCRJHT3k7vtU24vC+gumnyiaRJ5iBQ/6OzA/YMvIgaBOpRnxpLOB8FhX
e0BIA5u5nbiXxrv4gSeajNnauQDFTz7qqIQf29wKSizv3HYth+dQYSxPW8AJhiBi
bnYXGP7szPY0K+AiuibFhAiyYLVZLL3Y+AWBNMwHBq96vs0FyWi2aOgc2IeDbQn/
9fL3mRgVHWnt237So+g+7pxhRyLMR4YsJnEL8X6hkTeGSQFL6lNTUQnXcVSv7Lqd
vRYodH9caYS5luNjmcuau61Shd8i8CHnjUDYXz9mpzWQdWn4VBKEmqnErc3WFOoq
ZJeWvEe4WFf6OD33T71L5pCq8BoUDvhOXluOGXaamT6Wf3vP4zJJHdELhuof0JzR
snh6ITRbMsZOnJ+mMnNKX+iGTMxxOlML6RFKwWflOWVfL1u2D8CEcnqb8LsE3u6D
4WmrC5HIrb0FWxHaT7pI0cLBo58ki901JmdiwiOv85nERmiosUQbiZC0OSS6HpPT
M5Qn8UCMfwGTYJdvROIRZ0jIh1dWyBke4/NWDItXm4ILb7obLZ+F7575SdOahWAk
iRhCkEy1lE4LuAqUNCRJK1TmTkCUN0dZe9dIvaaOrpVAflEFWp8IcuHK43Fhu42O
uzdJp1SrAmzuKoCZXCzf/8XdA3lF3wVkt5eTa4gk2gzEX530CGa4rQzz+S89douK
kOcpEUqHeXWWsZ2pzPT1RBOBHcumzCFQO+5VMOxMe62wjCZk00bRoRduWuwKINSX
HYPnOvfPZAEVeJ/f0ERnfA==
`protect END_PROTECTED
