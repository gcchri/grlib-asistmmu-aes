`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FtYQDKeV1Xd3/7ZvhOUZ9R/l6kotcDGFRlkNpx0fKPu/wbe6/XY0LKo3U3bQmAm
KdNhP1WvT62/xgGCoAIT/1IWtZYMt6FprwueWu+fU5r4lAql1Z89gIDisS6cLmEI
akT/+gW70KMRf9frq4xXFzJYQJovH1sYyd81g/ChTCAyDhnBU3RCEEjam77UrXr7
+XBMH3sq1Pg9aMrxGMzyzPuJwXv3QZTudaM76podrsQ5WU8IbhIscDUSxYnUeTOl
J3ELiB4MCh4ki39VYkRyX3WzBWjkq8fi6CZPa751ARe+W/Y18NUj+lOFHXtFqrFv
zWS8i45Lugrk7rn/qdK2x+28CIh7G34LICNXfEBBzNVTwohMJt8TrlrRdxAFOT9G
8dP3UzZlHQxjM/viOtVgCVfax8xS9rrQ7vdsd6hkKr75mYKIMK5TqKnTLQSEr3Jx
YZU8KYnrs+Cc+hwIJJr1VCY+OFngaEtLSxPdMmv8wRZSeZpuohFmvLnFOAN0FK42
95nEbtfyL4dIYeihxtPyJM6zLE1XH7wlC/CP/h3/W7MpuhpFKoLs5gxO+BeMYGR2
UpneqvBvjUAv16ubXPYm1jlRoOBN22NubkkMZIQg1JBubMJwlyKH3INSPFOJUAHJ
u2PfRvwF8osS0oh/tTtOPEonqdXN/EcR4/+X/54OLilX7h3JzTqqFDgaNW55mUg9
mjrBRi4xAdr4kwUHg99n/ZQyAvyhDv631sxtL3+qFOVnuRJnkW4Tx8pPxktAI4ZX
ymOmsxNghLPUnMIw0o/828PAno/7bM7hc8d/wxhJ2fuCokQX0js+B5PB3bx+mKeP
8WTXSCLc6//u9R6tKuXx+d3OEe2h97FqIcBmkX2IUVBykrveg7Ixf2zVlm0tNaNb
Tc1Y8bNTJTFRwzVHRHWSmUxQwclu54p3++NzbJ5Nc66scwX1cJs8pNenBghdvlHe
rfe2FQYR75aG4QOuGgpQks5+MlISOo3jmMo2xPZvKZEYG+iH5rDPBkDq/e6w2ilq
NopGPzZRzSKVS4mYuF+6sFrkljSzr7pSgI6WR04FVuHZq3ds5J8bBT93VYX1XJ7C
xyajNCzNdrRNt2q7L7aZKKIYIf6Q21B5/GXt4ULUYniIBOWRUXOTDJ6L42Cf8/rr
GNtlAYuPxIa7iHHfv5GOmjuXKRSoTsM5GfAE8tn5i14NPwMdpyzJapJRB9+WO4XI
6CrBdkXGGlU4z1O812gRzZKZKtbeh33DKr3YW1w17+WA8CSAmJ26aaq3NzG96Noq
whWC5lACtYkR/mTk6QHAImCTgc05s6kZt4y558+yWgwaerDKUFax73Ad12uDhPnq
`protect END_PROTECTED
