`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fy+do/fnOQuU5WoiqKPrT7Y2oUoHSMHYDyciUUqhj5mj5gVwreVceTwSopaMO7D3
UyPbPUuppkG3LjpCH2f9+EGTF4X5r03sCEzcgXTiTZgJXIaBz59CYyVGUC1G6him
k6hXUmZkYjnBeKGdOWXc0yBLxpKnEf/S0gCDRyktMy1Os3M8Y2fFN0mkwmjZ8XPp
8BNIPfDzJp/qdqDvZ04zapndBaDcc5aoyBCfI7KHxKr1jO3D8nj9C/k/UjYF1sgp
mf7GlhZpEtM8eHYW26jOiaAmFem4dImRzzrWxC0LirwmvKtVb+bvtbOwOuEOkA1a
AFN7fW2VuWOJB4Z8RNQ2KYCHQaJf0EdwU6OxuoEz6OCYAJDLT6N/nRMuvH5GcGi/
u5dtJpyTSaI4nUNuwmsWlbAT5bIzwTxNcX2aff+O6bYcMzFYJF/nfEX3xgfsAq8N
RvqB9HxTrjwDqy3LVepEJ8X8yKrqGpl+tn6s9lFw0fXdczGZ+KI+IWL/56MyQUAj
YxttG0ThndxSfheh42skNIC9eplZVSPUvoPf2VKomQsblniByVMaDsbHpfvwzhXL
d35q7Kr7JaQRpzt7e7jf5Q==
`protect END_PROTECTED
