`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PumgZIZNzDT1tszBSvD1n363l/5X5re1NwuNXgROIHWn9KQ4AvB+87Gxg4SMZvcL
w/bzD7uA1Pitc0mqKvHtWvb5uV5VwsChnOiq4tJwE1uYXYJK6enJYKzR6Oxv+ssA
kngieuTPO31tjvIO4rVv3iZSK9sRAoS1TBy9WVUntTGA9YxG8/APhzkmhJbBA/tF
4n00ooYrlAwmShPRgrPJUuZ5AWG7Qx3Il8laMCprUzj3ZUbgAGl/ALBq6roWlTBg
dVx46BDjewsSDbQwQYhPvCiCHQexs5pUZOA8Hpm75kfPThuAeupBDKKc9XAGdhub
Vdbqz5VZuiPTXgFoi0TNu4+yTgcsPilAsspO05oimt3ZB6KV7xBMyPRLboDaLzBr
Oz2RxQackAuoLyN2cMe+dYbXczsUePh7UqCn7tP1oCpM8bDRlYbCvhp6884BX9SG
Z9QxKqVTd96D2qJMSX4gjCTM8YY6yAv7Em3qb65Iegz1MXzeW4hPtfOdKZwC32YW
95nesitIRFSGnPJ2phaThBTx8ygZ0SbbMudFaBCP8qzMk6EWx3D7X84IFOyTojuc
qQFRB78AyACso006ZPk/8VysdRCs5QD52eCTitswbLvPkqt4j1fDxyys+rsTF90R
IZQ3co/E+9+TZczCY8++LXUJsCfaOar+nFvv/QdHCBgs4GOrtSqmjfKQPqhVZlH4
Ff+ESNyfRnXsHE7RIJZfQ8rsFyMkD1OUbSYZSzvJ5bgSieX+dwQheerPCemeiexW
kVMpSFo/9UuKY+dJXkIOjoey95k77uijcLMJiVVbWG3mtyXhIszqJ/NEnnpqxTXr
uBnKSSibVyrj2x5UeFr9OOSew1hBBqJnZGDfmYmsfFsCQO2q3f+3HWRPXJqgGMqN
ocGQDh6Ef2ZBCFT0CVQrOm+6iFB0Omr6hm+eaiie6iou3/+9uOtlgnDhvRdIVBng
GVmwYYhUKQNhH62S3MwwAc0ImGtw6eCfUNq2ZlmAyO7/laIK5IGjfm2+ffv7+Y0e
FpZnigEI71rzimfOzqhvIofO81kpl65J114ZgQSoDd4m3v2C0f6n3j2Nd/msbWpx
gu3Zed0zy+zgmiaYfCThYJjxfWCEaDx1mVSKTgXYE9kMjHtq3g3LWTduHkTaHaT6
2i3Th4vf+FSL8aAcwKu76ceCtBZWTLbkMoZSA5j02GATN7d72OlSWt2ddDbJqMex
/G3ggFrOdyNI5bQdAbtmXFm9azIdS1UCgUxb4rR/UL9wJ850Z8/kGb5r7WsGVMdz
ZCZtevcAQppLqEyIfleed0iT7LqqRHlNGrfYBcMhHL/4tchJSpu2cWvg7MIjcG+K
N2aGLO4jLRheUgIneVYjtFGTxl0ZD41gMF1UHakQZDKRjIuk+E8pUMW9ayyrmbEx
tgq4JaJ+6Tls7+SVMEhUfXYrUdV93Kv4RGZFBOUklJdKfJXemZgFGAyuQqL/VZ1E
MHSdF6YfiXDDM7H5I9y1FKMFU9u3LEGpsZi2iqTk+dSTDOFsDFJobmXjpVtJaad2
KaZgugJpFo6B66SXcfA1ZXlXxiI6YvtBZV0tuoRBFJMu7pjKqaH2+i03r1miBF2l
WEmT6b2ubf/0EoJUg0/TkL1vFvvHwxduqOHc8bTWkr+qJytTe3dseQycwt7ODSMB
x7KPxNo+jEoD9SY0CFJGZDznxlSURCZ74fBzaG29KUpb3uOmbMcU+NoUsGycXvol
PWCx2fK56JoT8YTNM3mmrzoUrPNR7TWOKOxk3y9AyAWowJ8ioIfyaDsx7B39ktNT
EiJi8B9YyiYwAtzSbYBd1zfP5kZwga673K4PUjog+XJ2ne2Nn/pchpvtuKwpl5Qi
5pUtINNjiEZuL/Xkc+2tij5uY2IG2GOWJN0605DGkPC7UQkMz0hlywgQbE+ikxnZ
3eGRDeAy1mDQYbV35dyqOG6ubGsZYxs5ULszX/2neTajXnLG1b3WoAb3c+LSO3i8
0VjgsEQBp1Eg/WRTLeuE5sepWTMDT323urgHjkL9MuHlZLncJJMuS2aUyLdeg//A
MA5Ht6F8gF9GOmyQZw7RzOGbUeG7Z6OuZX/T2Ii7Do6nZ52xI7fbdAWARWs7Rtt4
pg14AYxczIvxrQyrf/2h9lj17p15JXmfKVtLN6oqKFLK6gsZVVEpup1zxMd0uKoQ
5EnlB3OWM/IT5awYnP8RAtvS7lT70p02R0Ia7GdApIfLfylrXpd3PauuDa/cuL3g
dD/q6qU4+8226ZJMR8A3aMRX5oxOtWgUSWMn6RMAd2+CKqdHjuJGQbvx9wjgtvEv
SqWELf4sPPp/JYqsldYeUdmHVLxNvN2ldF8J9PaLCrswRUoZpr8h+Ou6v3gjb5PA
21SrGWxq8rdSfZlRotrQhK0GA38LO/un3wPezEVMdQ4b0rYlmxrau4O3aQDm28aL
4XAYHhEtR4BkYkZvT4Yr+0ESUf6V58q6jU1rFleuJ+iK6rB/TUu30W5U59yk96zP
yb+pG3FsO0PYXHEKc2hMQpAJiGTIpbzPO9zyql8DVomjULbTGUJJvJvmQF8fvo2/
MjFIMUihtL+jv8t+L4phktVX2OLnyAyQcgi5zxVJKNz44P1IlODvLi9GhL00R1bc
lx1lkJAxeEFWLsgNGdnyxH9cFJPNauFhMqFlFh3xyNuT0Cj55g22QiSBEbHrSCWV
2bOMnkRMqCH+uqRhiHU+JlmyEqtvmDo807/h0diWlFu5ibp91PLyU0NGD50QtC0z
eeLkG+nWKXcnoxBlUCmFZ8hH7qN6b8jYk7iMgPPu9kw5FOCKRUtMde/NB0JAAU4V
F4n+yhbbeJqSovMo1hzqzK5Wjjd3qBG/Dip8WY+fg0R6Nasc7dAHi4PUUnI40D4+
XXnkqj6TYlrx5XtTGM00nfFY07cZirDO5uiRnP03Q9it3XHPXrOZRBS6nihhV2ra
f8JTcbMNmuBXg6tE1npltvFu2Qt0oxwxIrawsPTqgXh7QJGMKL39NUKI6Qpc982a
3zm59DSRqZQVEsWc8umQMgHh5CvfQr9TNQQT9hF5m7aZ/KWns/ET2X/GdXX+UVU+
vALDI6c60mG1j+EwxsMrnvbZzYqpZhlTf+DvIC/pJ0nt5UlR3rGt+OnlKP/H+pcd
DrOSR845GVpOJdYUolD4UoUae5O8HCVmCltFFvdc9S/iYOo2RfVo+CMoXrljZ+Ad
GBFzb39+C78TstBh9XZFq7xF1J310Cu3iDP+OIVobBbX9ARImLvBqJH3fJmpDj6K
mwl5LnFZ6V1dlpxc0qUVgiRnhXab0kdcuA0x+akhsv50V9ZOlUg9rxoMtKJSNByM
zcP+q8fFajREq2M9ESih6IpMXdEnTzM7BvZ9XPAuhXlR4TCJsYwzjkebrSlnNFd8
C8ONQkbPXFHWKK/tYYYenWvUSMYjN510sdlTMtWNx56WCOQuy4RfxboDS6BQCrZ6
tZ9CXLCVKaXpO841safM2R+dcS75QTUNLvCp6sIkYeMrsswDp65IhvwRR1WMu/Yj
JD2NWojlF6WioFGPsUH6LHilSUSnA4BrpDJVjc6QcUk4M5AmPgfrm1+8vkkF4o3E
dHjfeDQrJg903ryFSG/2Fq9/lJMgx9h6aSUHAiC+Q5a0nD0+QcSD9x44jT+q6VWM
RJq2gVXF4u2ZKucZ7nXk7egtktnP7Dw3gCcQMMepLxVVCWLo2UEDm5hYNLq6wkZu
CLegPQQa1L6zKpGZtTgO1nq+32hjW5OMlJ8tNsdtMYG34VCKSse+rNF0ZLi/5QMC
PcxsWqAzdJfYp3aLmW7fwfoldPrvLNEwRA3DEejMhhZ0peTjF10g5ack1FzTS7v/
RPG4EuiVr3cBsHDYBiaEg+Q3neZH5G61VZV+plSI8OLCOkrARRtrWJ2ldGb9skzU
pp0jufwapZzIy6i1IDEgu7iQfnQbXAw+nubQnd8bhlhpt8GE8WTXCZsjBlD7Dm4b
N5ylbrxH99yWt+QpDcgQkP2jHumipEAQEViH/b/sWfXSamNcM40J9pu+OwN/tRjX
ugB1IzMxRxp6LE7XI/jPn8IHYOZ3Mfd1n+w0byZtpbg6J5o3M0RCB5TFrMt3PT/L
sXALvpOebM7eocu2tBpI7oeS8C5DUWJCunC5c2493uMfza/jRH8S63rB8kKzrmSN
6yA96CvR8zjghlbb/RJp6g2pIqeuj3NwXAhFVFpbXayf6WStwWDdm1kmCdH9Phs6
wCYgrwpo9yRiBPTEPYT7Bno0wHnu580WRhJQ0eNy+cgF750Dj9I+bTpvKb3m0mqf
/fW0XJ3G5GiR12KfGlNzZu5IjzDAS+aaq7EP9jts1FtV3DFpCsy6yS6Uen9s9D7T
Pw5uxmOQOH9EFq4mKIsheGkFoBsa7l+ibRqBiPuyYeK5cboT+dZa606OhXq0TC1+
mLcwvWa67KkVoGHlK2VXF4n+A1fdk2gULwaAkwHVmH0Err6kvNSlyikEPaIdjLnv
uVSTgOPCkm5S30WXWJtccpRRc8iILLW6zJx0d3ruyJV3srPgLvqaL7fprIM/S53i
1E//VX4g4izT+6jhRDWMeC+I/tcRZ9XZhbY7fclFLreV3RKdvj7pQV8JtjjyVYN6
5fI0ihZCj3ZLoHtmSc1TE2tbdGbAxRKktY/qiCuxTLsGX1LsWQD8ahdLfM3lrg3Q
+0J22WGFBBmxtvfk+Xd62fGP/sCSDdhuy7lzDX/hLTTyjTUN8D5Bs3i6eOOXCN/Z
a4WiAyWRHHdsaPp3JWy4Qbg7ReUxD6p+qGTnxT/uJSPA2vDg68qYTzKfLe23lxy1
8XfB41zMlB5xYA5midETg6porsCe0CBb4itsojflCSod5oDMsDsLtyMs8rydrNSK
/XS7lMgow8Y8TxRultYVczWLEEliVK3Gk9pPTclzYUbNsxb6Mv3nLRmUqXSGWxCn
zfgBw7oqflhRXdBoPz4JTABcrCoT26tpIKHEMhdzRJA65TOYLrr+UO3ra7beaJGd
JpM3AaTCtQOgbpic9S3VncJ0dm5T9sCWSfvTZ1Zi1yUz1BlqYOmqpYMnka9sDzOM
E9jX1ry6q+9iT+1aWjzgfiViXAzZoxXnTBTAYBgv09g2c+Z9F3dFGcOC9wEFLvXK
9h2H3+bJHRPfgmsoL0+sp/v5Ftvp42gPIi/edkYAzEJh9DiE/fRN97rAzrhZgc41
ZkAuB69mYnqjqWIFdo/VtqUlikwjaLQk77MmbwG2SgqrpnNFVFE4CImxFz3nyTRs
S4osiN2Ob4cwKSjRWE1SU0V8F7mX9W2DrBX6024bIHbzYhPXJuoCUUCPuSHN507q
Em/dg0tK9J/P6UcBfkSezuzUejEvAjAqoN4PjGTg00Au9J5hV5OBjsH7JMNlbA9N
OxAAiHBzefyIHAfjRYpzMvoDn8l6fW8G5qqjpe5bIWx7cFj8t6TqJXFuLgcYsmh4
x8QYHDeEL2iXTW1Tl1Cn2My2QsRaI0pkobwIG6vLtltetajmUN6RE2QoVSQpSvhI
CrnVzJ/YBaxlXEBChhGGAplD2I4LRXIfmhM+1A9lpO0skBmZ1qMeJH32uGLD6Eyr
PkWQ7XT4vBYEJ14LIS4IIxl8tewTpWbqxDAFY/uz/h6I/LlHPONa7UAfrTmt5t4W
WsKNbX046785hYKBWKm3IsmdPtSXji6xnJOc6P/O7UuBkhOmkrmuVDGN2XLSSHpW
P0w8ce8AmSHEy/W+cApSCr1caAY3XMSsr0JUvBJevLhmRdLSiW29MP6T7Og6ub4c
kr0rPrm/aGYYMZOEhPaatPINDwmjxYFITnETQrTYioyJrqtFbBBgMLyuj62Vz24+
EA9DZy+UPUmQMxN4WL7w8BXkNtKgq7S0Ah6FqeywyAMEC41Qck5GeD4vb5tD5YwF
Jo2RwG+7ugsKe2x9pdexZX/GKRvvBW46FlSpxd5bjDSPVU8PJzomJ345bVnVKT1h
/xW21j34A26TmZm2jdxTINp/y7Yw18yGljse/La+8CImyncCVRMPiz/HhJE3MAzk
CD4QTkCwHeMargYkcWpYyMhvAt1xa2RAzsz7OkLMwB5alO2xpf6cO/uI8fCyh1rk
oAJRXuYUbxQJu3coDRn8ACWvBJ3rBlT9AzQGUuxcNmXpAhKOmQ4XwMkih/Zc//x6
xOl5bPp/0E3wiCMGfQyqoK6CFfoEe7+AQzfYHfk41yRI5odJjSQ290Rdesf8IIsk
Hy7a9igu4xvgRXMjud2Ji2MlK0zku50qR9kIG4wW8UhgY/juOp4LlEWr2ADvbf6F
vQP5gf2JSNpHdS6eSQgZMSUujFD4irf3pVW6E81OD2hKdBXFY556Cd8SFJn3J6nm
yvEIsMiZRTvUx2v9Be/FWiKOU2acvdofrdlm8Fhx4WtJrEuhH7Ym/q3P/rMbwELF
LmmxsJ6lclvH+ti7hLcM/X+F6ali37oAY7BCi6hAONnucSMrInYthVrnWaBFOmDm
CWNs953UFMTYbZFSOyJ332aUqlTwR3NQOhBYfRLD3qio8CLHlA4nPKbJh7X0+l8j
q6YAFKc73UA8vdPUX5MV/kQSJw6pBhbaB5JyKAXU1lFTiNl35HivIcd082D1c4qZ
5OQBQ1daSGt6RTcRvTdSYoW0K3X9TD4sjkIgglQw0/bkMNMbH9hrL+G4AivlMpOn
vfft35NCkifwHBPS6+KBdteFavQEoBz1n6dy2u9IolQhgXqP1QeNKuBHWdnr6aGw
9z/ovrbkGF5A9udrPSYm9zjpnWali1Q5F/OU9SY9akKmcXgHfqAzqci4Wqb4JG5g
iNvmAQG0qqkPlnhpOCnlniTSpFvdtkEAaJi119FZzO67b3PGN6yJpirVUT69eSQT
TeF5ASury9DVurfCP8pRwL/A2cYiEUXW4emkcw9rg8QMK45XndTL2xenmP/3Ub7E
q23sageh8hdXoZqzdI3mgQlmFRpZEv2955u+cbLBcUbtX98l8le5O22AcfuHfBJC
MRYGvmIa7M/g+QYZI6OKrwoce2ROFY1t69e1+UZ05CkIkNFBvX4YV39MfgFzDOsh
iJrn/fsgE/uH4rZZjSx5VOc1jICURlqE0QFoklNGb7E7ts3BkExP1dErbGocB9Qr
LoETVklghUESkhEtBF+fFTMArar3nm4lKuam9a008IuNPLl+OFIkSMOwCiQZmwsI
Hr4C6MUINELtfMqM7bP1zRwFMlQ/FBJypps1oUWg1NzOvJw1W5gOk5jFVnN/fsbp
WgB/DOCFT5tUWIOkRPBXQx0Uh2udhHikETehvDR4lTySACz5NcbATvlql33sMOQs
CJP++C28vPM6Kf2Jk3YfDmTSof6N8wEWbXmCJk8hfBUSprHgyV88PsCaxluXVGMB
oVBRRwlJMOuSbQoDVp2dJXZEOSQPIwT64GnH+hiaYyR2j9yp0pWGE/PNN9p2z66u
5kudHL35VNTcT2V/YINfCtJIn4j3KuCBgN4GvFXoZcRThzvMaF+OXG6PsOh3vt+A
gpcqQS33PVpj4B5nUxGHPWIvIA80DH3bP/IM1aDKA5A+QbMylFzIWsUFqoDmzpqY
3Ngn7oviSs9sUVvdO4+kHcyJhIbuQ4Fu1BgKkb5Hu4OQ+jYcRyfqK8y37FEpYoqd
J0aM6MEzIJ9Voqm4oAZDpew1gRDMxRWGMI5gI4NZnltUhX+I2OFiH/JV7rV7xORQ
wTiSUw+Lo9vcRblWKkya6hOye8wwrOi7H2sEzCmIW81rHWPn/PEcqC+pyOPoLsZQ
ViS8WX0IHOY/vwVQJmgGbUUkBFvHyTThlpflJ7amNOyttV/cDaI0kfmuEkyC/PpN
Jtv6jrHRFKLWWpscAJP+7oKlrblktR1kAimuA1TqhaHdzP9xhS3r3mSVYKQMMX+k
RTeyTsuE1kSR/CkCfEjh/DbFFR/EgHfjT/2eWq9taNGZsCWCtpWFIGIKW3RvNWTe
sCaUEehSlpI6TWP8DYWqDoXHpJQMfxKaTxmNdvQM9GUiDY8UfBcije5+J2I6nqpx
5mzRxj+cPeB935KwxPp2yYOFusRCI85qd++mpL8ytornGtkevtJJ1hVimFJihiYd
HrbrqicVGCLtwD0BPo7xV3yeqUlYMtzCLGJS5nLblc+16LoJpD7KpL0DeYOzKOtT
KSPxWH0xUkabcZcANZiZAIQqqwCr9LIlZdGQuGSThqZ7FtwDpB7bAIGsP6jL8fAp
UHLOLVS2GBMy1icJolONLROY22/olKDFT64as3WqhduHF5mnQzeqmZ+AfjgNTSVC
OmXCNVKWztKOG9mrXSZfXdTaadEexf36BnwJxfZYBmpLfD9cIuanReAupl8TTghq
MnhjqGisdIpgtirEiekWDCUaTGrprz7kGC5W/Go6lsG/sOxzLeF3b3QtxSQ4ZdS4
2R60n1Rh44prMuDv4aQhfqgdO0vbyaoSx7zSQ0wUMDB8IEhmEDk/gPL9JvPNSpaY
0bLX2ACkWX5mcFR2bLzV+SUB/CjK5KMU2niSRM9DpoGiQEB/quC0ibNRy5cCWMZu
BJKei4iTaXrwXFsco7RIzBqAx0IzrM56A4Xrk6HWZMPbVW3j78vK+VmvTYTaS5SJ
fc9QlpZS4+wRm7H+jEXCfWSIfb2IEmImCakMOPWUCzBAUWaPYK6cs/TlsaPCOWFH
6vhMAPMO388DLAxV8zitGOnrScQfFfBzC9vAFHxJFwNJLowp7J5t974hHMUNRjtC
gqNXFanGYQj3h0S/v+PBfWmQRuAP5XU50ykDR+z0H0wgRarK8ywU1V/1fAcEG9h0
lL6RWmymQE0KNPi2zF1ZwByoc8VIBniVsCZwBA5k+Mdr0v6SBcHZaUsXBOCkdEIA
g2+/1pWuERU9iC7PZ2N3V3Bq7sqUEOnmBlnShYCZqCQ75djcXYuo1jBZfol5L8a7
QvA/3F1FPs8sYc16tJ6JYOknqXnjsU3CBuE13WGEwpGYYuT8C6J5+Ysb7N+cetYV
0jMI1zsWRssLUIgOqRhAcjNkXYVy4WDwpE4m+AC2+33SlYOVDBdMB3TOFgO4eCtL
8Hp4E+ga/yQ0f2mb8+NiLF32lOvHty+e7Z300sPfhpl4vqYlBs4Ii/36tuyvCFOM
zReDF5eKMw6OlKX02XrD235nRt4u0gp9xblHIPDiUEz7Jd3dOzU1WSSsGGMF5DGb
Lhq+YGN8Vm7wjZm7T/VeAg97sZxdRU1kiOPGISNq28OhZtpGGRo2/KtJXZdghEgU
4xkbP+DlI6oo2wNZz2K5ja3DUCYX+LF3hDGonrErF364f7PG3UkEuyOyXDvhgtPJ
VkyXMFx5LdUnHztEroT8yg/G9IuyRNVZwBWGcORUiZfigkb0dAAkqBvBB1c1HImX
aCCvWKQgKKodfxDHDjb12PrwEz74OcX2ekSXX2q9fEr0A89nF0a6wqP+33wlPHRI
OJZivd0OAusGAmh1j4qihyQrIzcTbudXMUJevSCBKEvZnHdOR2tURZ/L6TzDWcXf
HMxdZK15vbXyX0LoLR1H5frp+n68tPKtOjoNNeIyxBFg5LJBswre2xMKT6oJcSrq
BjOPrp/e2RngcjUrfN1HML0kNKskqIdYHN2tJvDDn4YWi5hTYe4kE9b+snuNpJMz
3ftZMc4Yh/TrA/hA1ogaZV9LHrx2o7ho0I/QA3ToL8kdz4lbHKd8EUGeVAA7KFiF
yYAegCmjRFPS97zzckDiQRIJVYWvLAI9VKH2pxhOfbIW53Q9Q+NyZhgfFQUOSoV3
XpvK8FFSVZRV+9GLNO4l+ZbYpJfrUu8nlgYM05ce34zmNENbV6NsYxbn0pFGCBHG
qRz2W3ag0tXLa+ZfhfvSTFXYX71QgvsvERgdZYOuE3L1DQaslKP/0JIiJtX82xBY
rteZHfdPGbAZhRKbHXSb1vv3LED/CBAFVokeBZb/sDTbPLw4qOWEr9nDQe0VflbM
mtoHnEXO7j7uaVOUIUxgS/yWqogNL0bheNovlcxsuLAsfPFOx2L/W1GdVEv8kmNQ
uzEFlSdiM0rWUOZscEOmjq7VydK8fi16sCz4R+VIci58t2z1bXxkPjE+TiL0n+ES
eGTJVjpXx1PC4/czzE/vAfQDnKZuObzfyc1veLBp10tggy35UgwRPw4boPMNj6kX
tW9kzWW7T2MMfrAFUzbedRkRHxgHojYrgpXVVM5g0q2IcClJKcZ3Aq448684QjmI
vgXp1F/UVhrt7hbyzGdhJIjYlbFueFoEhWwBpyvr/ZILuHg8P++9HOg4GndDffoD
n9+z35ESOmvGmd4dpkcocoMlok6gOywh8frbWtQ1T0eM7bxIOqrUb8+ubTDuiNNO
vF+OzLLNyahJGaJ8MGcGpxwNpN2FH51zgW340a5bd0c07WDeQusQ0Y/+zyedCia/
ucqN7hsVqMzDT5YF+BuchNwE9yVns5F0yMTex1C7ORtk3EAWWYNEYv4foqcC/tQi
Stjh56D7o7RkI53NUVX/jiqjnMG1OkeVHp4eGbJLyURBYxjkP979IRPVUvroBdBV
jm4Rv7Toi9MLsTK5Xxfn+1d/SFMWbxlVQlF6ABYLJhwbzyLhhaCaoJVHz/hY64nc
31P73a4lm7kCKHaEr9Lokc7pOa+lWaDNLgiNxjtfobGB573t/AJLYRitNF6FPpk9
ZY1tpWPp2LXMOJh2vWfO0qkL9hKlurNAGk7PIpDlGcVydw+VgAksJT2YtTd4+AEK
+BzUDeww5EQkm/Zn/t0XadzaeoJ8t1wV8BfYDX4H+/Ll7vCZXuzxMvirtKv3lsVB
pPifDd7q3AfNcPfHgZIpTQTx7LVkHLjeqMEd9I6SdcFo66S/AtsJc5z4prdzA17d
+9NmMaJ0tg2XFtnZSqKmrlwYIXqWLNFWx1GFuOVZGhbJo/SFlZOYAxBNzjHTyKlB
BZsV+PWl4D0yoeUExviNnw==
`protect END_PROTECTED
