`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JeM0fXYj7QwtiGQLEC0G0EwDhbIsx5XzapkR1sL+4KL2XIB3/YTd1BF7P/sB16dC
Nigm/DqDjiG+eLhLVzYWjpQZVxkmOpvlLVveeFi9JR9rnYV2G/1hZoLdHHg3Ez7N
NOGqUEC0OdCsmno/h8se7FR0WB2hc4T4mduyOP2fIu/r31nTUubnAco+HJFgiPng
mIfITNs83t6hDfOFPbp/SG+u1Tp01t+ohnvZPLQ+pRwuE3syJCFePduu+SEX7WDA
mZauz1jcg/fnrdvPCv0UXbdbJpMBDf97lt4XPB1D59zB654Dt0G4CsakmTQzBujJ
xbMbWwpSMzTFdsUFnu8BJ+LXfAh1BNHV0nSOZ4QqVl92lBR2kaoxJ8tOLOgBfSVj
hV8L+b5dJrzQ7ELGi2QhXyvG7zHBm+qGtIaSCQmL0A0B+VCklqHnfkVdbR+th9jr
e28UxPnuHias3yKJVkKUTg2I5+WleZcQGY1drDoDvLHmNaExMAoqfyhh6YnMy/rV
`protect END_PROTECTED
