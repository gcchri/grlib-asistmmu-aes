`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Ou/vtEREsCKttGou6EA3VbjCytDEwBJDMo6njEyegE3QEHX0p8TY8WWT1J2MoVi
3yyDZ5Ekye6WxTidCMGdQw3/5THc5wyaD4stHawgxrKPajgnM0lHSgD+rG6huN/A
vW9ORXW8YKW6X2EYRj82sNaN2fBuPjyiTtMNAzFVpcODnw/SsPdSLmulRnrc38aq
CB1vFrX/RcLlE8k3SiLb5s8Pf/ONVauN5quQwTUorLId4yICBPqo4NXsgD/CjjBX
tHYRn6LNBm7tOOS5JX5jXPPORmYVheQwLeMFmhBN/Ejm72hFMx28fdI5ed8bE8Bx
5b0TaUG/sDhpU5YWwCBIiuLUOln2EFIt0Y5p4mm3W7M+FEElxVSreSR4pFGgJX5O
h9MxJHOh1AS1ieto2w0TvM+W0Sn44UNP48gefKEnt0eNCSn/LnVfo4Ks+OzyjMp8
0p0pG3H9H8jFUQ4eoVjRHcMy0V/Wb+LmCR01Hrc7e4YPSue9nvCv04GmYBwECjOh
6kzL/wc8qCQG2Nu2e1R8d/p59ufBOekXkqzzRG1rRQMqw/z+mmq/fJx8Q+NMaBbJ
GxYr9cKmHq/aLcv6f5KIxMPwbzRbkfcECcyONl928cX3vf/+xVSjE06CBWCgSy7o
z+m/MXVNYYWQOkgVk1ZHWxLBi9Ebn+fc7h+KxJPneZ3XrM98AWyUDiDcxLnnJiv/
uCFAMiSmryuHfUugg28TMgX6bGATEziFw2FOoxOoKQ1gMrBEwQewNr8/K8de38sL
1bUGL6Z/HsLpRpliEz1SvAv81PF0cNljKiNc/y0GMo6hFq0PeVOs2tTSzKEofr5g
NZnxXcb/MmhJ/i14COyo0RziSEivHQiD8OB6OBzsLB9tKCYWjHmkoCgwP6pIeYkE
xex9khf6jugZ6NEBC7ktFxGiviiirvYdEa+Eh+Lu4A9qo4pfgZlFYMmrQf5fZ7QR
H9tpE9khQg1e39EwbXOFWV2o2F7VriHrEOT/s5mpEjMI5RnLk+aF/Rnj278TYtiH
tKLKM0KmPmMxO8shD+G9mU0J6RWlwweh7+ThwpZBzjPTCKgGDaMrQjp7QC9w81iP
2lnEq68oKn8bx6PP08AwI7E9x2PPK8HjT4o4TB1W4hcpgc01lC861NDEvYnWL1L6
7r0Q9MMimKb0Rr7yNSXXD2C2xhkh62Nw+XwkCav+xBvJy1iAqfrJ8N1xsPR4ULzq
3mvqmYQdhrCsyePa01azJVLTm4hgtrebuEFHsFbrPD+mOc9YzkXDXeNFn9GrT+eX
YPlrxkCRaz+pDk6C5KwnyGL8ko9PcU9KWaAznQq7AYzEN5YJeqljh1ESlqOTzG3g
Qg5oevLFy9C11npzQbo/IeYWYt3ptx2v2bW81MVqg51OSN5BXNikAgKe6KChPsIe
K7rjc1OEonZ2InvokQBQ/4m7+sBNdTP36Lc+SF8ue3sMPoMabl49MxS+3Xbj4MyU
DJRRBR41R7BkquLH9nQyI4TGYVoqN2fOEWZfHTMcezxauLKAonHJotq1cVN8J3YS
Am3uDIXGRDiMVzmSVB9oNlMbaCahbsM4u/ofzT6oZspU8qic4R4gZODNX8sM/9YE
SnV02EZjFI5iT49/AHfuTXSujt6aJnxvy00F98b4b0afT/buEW+4Iw5YgeIdCQdz
BOOCb9PtDfcLv822avt0DX6RdawraLnenq1FNz6HgJ0rNVP/u7vl4IBlOMgpo9tM
oWdRE7UkOevZLpZXaT3b+oR2y2JS57lVDifo5dzFL0yTUwmAPRTULJpDof9hTwqA
5Rs8+l0DNiMKji/gVdMUxfa/lvb2o6cheCbG+56EJgwrqqQQ21VixB3VZQbb5WMq
p9lM2Jp9bXnC/kZU2JRZ8d3o5Frs6XjLrTpjgmitU30Wy2/J+Y8FInGehAXtq843
pscI/Z+WbkqaSYcxHrPeSrPsAOoPIMSsw6sC1nIwmCGVhhFnZVT/fYmlbbNAtVqR
a8pwWURFQl4G05zfzaNijc+ACTE19eeUZj5AmnNuwhwN7aco632Ogxp7qoXrC4P3
5z2DAwb1b0wxjCdIjLS+Q9OXj5+TY8J03c9OqA6q67610mr2+PJtkk6COiykQ7ap
5OrfNsubdEg246dEVqJe5hEkdKpzjVoRoNMSGSf6+aobTuSDoj1OiB53VfGvgrLQ
D/TKe0tdtMFoXRSB7wS/ZqftdAywE0qTIFH48tIXbITV/BQd5v8SmZbssWqBavL6
Jy6BBs+gdUp7AvxxGz68xiy9ciFomHVrf6sqGbTaE/+w9D6IIvZ6nVA6Ry33Pod4
WJLNLYo6DOJ9LjqkjQBgozUZOinywWEJ1NLwu9n/xnnNbEnSGlWTZTc7PvRMJPOl
b6/yQWsqaZMA74NuXVZA344igWn3DDTP00TCsKaHvFMed1G1S1FD+jr0skTo63Ra
KPshw3JtKQgcepCyvxvRm+QUQbVUatfB5nQ74aiQJ7LneonxVaTChbPc8xvc6WVa
wqujkc5v+nCzn3kJzbDEmW6JXIm5yGNbxdksZxuQqF41zEaZYgBmeV8uVo3mGEKc
eNBRGxbZkBzokQWd5v6RyCiAUnpU3mXiRBqr7kTEvYzTLyq5DtwbO1PRFeb/u0fk
eSa5hB/+IKaPPrHRdJPOFxSQyN6dsb4uWLCxva/85pZ/zEXm1la0dPjgY8ZlJp6Y
X8akVOI2irnnXYAcjHhjM9RRze81LEWfpxUb9Fuz8zXZlxT25XOcm3LjIwVxfsxy
5BDZOYTfiC3Pff15DtJ6uoRIKmx9Cw+Muh6ZIuABqvKlrOjkUf/zuHihG3QO2KWB
KNjQeoSR/jvSonGxqerWD1yKm09B7bsnlblwoBAaSTH3nRNk20sUdbeAIAlD7mZ1
NsRzHrqdyrJt09flygpj6kDyLZ1csNZyBV7CJTrrhYAaZNQueM+km9qSwxH5qy3S
l8B+5+CVFL9HIJLMPOhYbt5N6TkMUowlnmGefrNdNFE/dKyQfFZif0IJnd3aAVnz
tbufSCuCV41l1CQZlwbolPRH/F49KjhQpRsMXeWL0Ev4ds8xGbvJnpsZeIOWXC+j
V8cHXvz/vUBlLiANyYOklMcljEVH4SGSH+7FptSpkzL8Ih9+PMoZtnZYhfIaZJGO
Gc+bovU5t/2Y5eApmm7z+00RzTv1IlpRdZGQfvw34ltbUWl3C/SPEerUoAtT8FsG
cIkf3+2pikVVA9t7FO+X9F9X0El6XnB96ETo7CU9iDcStlF014t3WBqoxN/voxoL
/Htis1O7HOiooEk+l0acEfa2/eQbuyEYjRxxgidMXGE67T+bijESe51chVY628iK
XGUCgRDmfCHWqh9aVgBBcX3w5pkepyttDwzi/rL06+wDFfTPVq7t2jDHYCHBHJvq
E8EnliwJcRwbjSkoS5JsiXrrpl179ZzHvfzInX1pKExaAYTkO4ZVvkF2+voQM7xK
yJFt4gsPMGh2yWlZfPk1gcK/TXvSvOqkSGRDv/+sAVrB/ho0c8OwgmyVmNO6etkX
HjrvWlehyKXWVBJAjyYEK+xcH4Kiud5tw2SmFH3UTd0SlHT3G1DYdgTZ+DvzLHsy
oFd/PJ/j+4BmuYxnJdLziLLTdFl9RkUPUQ4dTrNBwH1KL/rZAQD0wnrVBzILtee0
35tHR0TyQ+nWcyp5x3uVo7SV4+DdRGO9rUxtWE0tHiLZ+9g9mYIPkKRMjNJZsSQa
npCl+p0dEnNCM26pWAXuuGbwqJN7aKst9ARJ86iFcbsWWmTLuiz69L7Yt3OY1Wy9
hj+0lfBEop4F8Z/bfHB3SQ==
`protect END_PROTECTED
