`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xwgVvbHlDSP2ErCqzKNHXcgkxX3Xu5ePTBYMOqnp23b27gNm89qmD6fcpvltTgRy
nUAzzgIT5u/Y8KWuyVPph34NAao/QNayFNEyKYSpYUSeavxbDwVfojhCDb03ixFk
XVUMDKOx8VIoU50pHwu01V4x1QBP53FlGOmEt3zRINkMrFlEjwa7cSAYbU844+P4
3wJGxxGg9tRQZjcT7eqSTlyN6GhXbK7eimT1kPllcaTOcOM4lQBab9nqW0ZvgV4Z
Xg4k9qTnor3d7jG6fB0yVhPrfhQdHX3jLJxOkB/yRJQiftNK4uz3jF5Zt4rlje/W
5nAbppSeUdpbvemZb/OGqM4JVobm1wYktlHPd8smwuhy5cKj6kADOQhpkjKSX+vd
N8D4yLmcrUOEca8rsfZN5PgUAY24vLzbLYHaFv9CBFFn0WMBsGokwOP2Fd3rZcJD
0V/C2XMZfvKS37A+hS8kmHJaHxyn2qKeXl9spSuDRuqk6altA0G6o3qUgLQvuj0F
8YtnsJmCLpIj8ZTBqavLESTRJ9ZeybjO58o6gbqP4EQDGjoGFAb1POnHFLd3/hM6
`protect END_PROTECTED
