`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
066fkmGopsKqwfs+k7q5KVvufrVyu9660KLH8IiWvxUsBcXtcfL3Tkcz4pKMonHW
detXUPsyfpkv+mfeeDLw+1BTCnExA43WaZJaiRe8tKLezsDlXBeNVORJAokz/8S2
oVPGv7gcCqz7vt1wkUUvjByTNEZpfbfRV2c1uF8x7VhgY2XpT2gcCQIYZ1vRphI9
2xswbcHUXti0peSdWtlReFgqm9aadieKqDSzXfxghmvOTXMAib+Ws2HlpbuUdGUA
9BppQg1HKG10pxpIsxaquTSuQqBwNxIZNv7zzygnCmXVGo5qSUzfbUqJ10/TB77+
yJ6sHmOb9IMuS9+ocktGsqm+MbFUAVH36XgqixGsb95cDFEpafC86duKvSfyF9hy
EkSUn4kD1ij1FR4EnWl0gpZqJvS7YWnXxWvqKCeDXL7Nq+GI3XSSe0Qfa9ct7OCb
5VJFvJfICEXrf7U8Jy8yXhzbb7JVVM8zJ++VCFS1l8EESSzE2kXoJXq90RqAe6Bx
S4XhiZEVpK4UzbYhDbBq3Pg5gnFiCHqgItnaKaZ5Fx3OTNDLMFaw+dobkNaQ7x3E
eDNbKt3nYwxXroTG1o1oq9yFNLWBs/R0WJcwZ2q0Dm0PHVQeFkRZRwq1rR3YRU+v
o4kQ7xiztlEPgzHu0p9hhZV9AVfzLIaM8wLjpWhAhnDmOMYNOW+hcnY43vDnvwep
A3kJqc2DZi+TI7A5XtJPZrkWziSsri2fCGkChhFiI9k=
`protect END_PROTECTED
