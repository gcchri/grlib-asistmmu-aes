`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXQxFLtZJGnDR2Jn3tMsYM3lnqPJ6+/cjCs7x39YQkF9txSt0wuPYFkM5U8BfAEa
dDbrO5yhb2dpSuhSu+KhjZ2e5VDirthGFC/SGi9bL9X52cqgfUdVCPmcoY1CtOKN
dfV/diJw84pu9PNI7HbcmgfNZa7J3mDEBlD9zJlWXUFqrvPVXgDiq1sLlu0P3Uqt
bG28mFyaJsAx0yXJw4lmmqH/1huaSDqT9LlVI7wgirDAK66UOGxPTkwqeu2AK7rb
O0VqZc75FTjVC7z3af69aE6Kkp2FfE0gL7IguENqHA68YkbLbdgOEFB3sMliCwhL
8LJ3bSymyePVmY2iy+hDBU9TPN/OYbXSvoGbd4aAWh8=
`protect END_PROTECTED
