`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mVIwmYrkHt+nsA2hiBTlDe28nPE2xMiXtw3cYgtUpnknqetlYSPpANvGUJqFrnlx
uCp5X1xcvhTaV+lDB10yh8rhZdENFjkqqRDomKCIGToDqK1Tm9GOXzYhRDLF4PUI
tT6yGRUYUZ6vcvmY1DtKflGFPyPNmT4TpWDysoT5PbHRhv7SiJXjTxvo0QvMjz0A
CXilD+irhST3hKgtzU2hOYXoR90U8LNu+QxM4kpJDF5FuhvlvKdmlMq/+3qzfNlZ
Bfdi+llUKwsQHG2T2haJvoz22romgUIjxfm5si2JD5CrrdH9uQhR4nVu9ZthY4C/
csO9WjeKyyOlVPlfTQWWv3kftLdjsaLPuWsFxb8vImAJLnWAwaq33xj1Dc7API6I
qe/H/tl+1fG+VWLMHcLrti2NNx5R5y0M/XeJwhqNhHI=
`protect END_PROTECTED
