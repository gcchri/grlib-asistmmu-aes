`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOYzodkFdUTDPDSaQitFZIp9rBvUyL2qhjKUVmROtT88gaVrGlt7FRlJ3/iiN+7S
UPCOqy1De9duLcAxUHE2MAx8dq0k4SlSFTBLTCjptfu7Zga3FyAkuGajRirT4pEJ
fmRneLlJIUpg3b5a/wBVwHqqfGncDbKMwoLzP8cKD8P3QLWmSgR+13a6fAqy/COC
0vZawsy+QxEbwt0NTDV2Jm5fxXnYEIZgVYDjA9QzZbTWguRyuePyuTrU+vK+vgyi
tqcFQXYxtacD8EkQTcfmwiMXp8IXYb43Up2EZKtJeMAIDtvS6FCxwmkFj121wclv
yBF+DuoEvu7N/CUNnHxHTigTGIBDZ97LRDJnIHc+rlo=
`protect END_PROTECTED
