`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vYmWcI4vwmWnwYQdyR8gHLsanPQl4PG5/jdFZqF1EiNcKAqP1HgHIQ3X7nutVhPr
brz5b5UuD6SwIGjzpoiKVs+kDtfgDkYr7XUA+NFJLV0wTfHrpdwptULNHYXTah6U
XZTJY9PhOdd7hpeD5YXyvorC/oJVxdl+w34GoaGkhLV914k/lMTGaNfmfSPo1jPh
C7OdjGmoqFtP0Sd9Fho+nvATxDQHuRjuCUUCzdHh+sD5arrAdE6avAhx4yq6dkSF
HxVQ2PxMwLkzjiTwPz/YVA3WteDaDO7vxmQd12/x9MxlQ7yCnMDfvHG/wSABjN2f
UaPY+SfYWRC6Hu/oyUrOD+7ZEhjlh4xs9qiKifQDj27L5FdJPNopINihnMmlvzlY
cPzrg28MAsby/pyT7Tetz8x6tJK1/c+MBXYK+MUuUgw58u8dBaKYPSrthuVav6Mj
pb9udPYzD41/K9KuOR8HWNyFjCL7qOUGKQEOqLomAot2McUtA5vw63xjYmyLU6oA
NvNFUorYVwYl6X47KxMt0GUQmc/KDvZRJJSJxSA31c/k2bUy3403tXXuytjsbEyo
mWWzx5BXBtivHJhlPvRxnPeFkiYqjhBYe4uW+IrFpXSwP1e4nzhpMqjUifFze0Dm
0ByKjxpRU4801Ly3Z6mxqw==
`protect END_PROTECTED
