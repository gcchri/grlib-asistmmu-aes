`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/k3vkSggFhKrXZ8XX+Abpz7oTzFtESPR/yssTvxOFNWx7xPfS/6AMd273+rrn+b6
DwF4oY3u9/JAOqg1LqDCKG4fiYsObxCpEJzACw1gWI3YUvYf20UPj+S9rJ8/GxHn
ewLEl4SR93wuKWNoGPaSosvbMGRZd5hzPffl/9c5P7O54AUdpW9DOH4yJqS2u2N1
Y6xlsHZg9vPuOZQeqq/PlW2+p+OJmKArTw7ZzIQtDqU+Xdxm1JXfF1elFPVQ+N0P
CiRAyhGwPxaweWeE3ZiNszQUEg23aenA7LQpnIBUPePSUTDzHKFanQrDfmSoFspH
B9FPRK8ebowVQB6KqK0liNKKmM1s1sHQCfna2xZQ+1XxI8i7zr5DJyU9O5xZTJ+H
Su1jgaCdFdQnNgXwICTrCROfZUg8p+BWUuzlRGxd7seaxNRdk7C1My4hjZjrnXLe
w1NAz+z+5ccX+nd7sSG37E3KwngFDB7rXldmRb3OrVl0j6akdKM3EDf8x4SJt6aN
S0OIrq1nVwUxuIAb+nJDlfQvcYosAW1LJsl0q7UwDpFsaIO0PJbhVsdOBTtpy/N/
QHd1qsgTAiri3U/v/NcPeKsL88/kcwwPKWo1YmLHgaD5UPETscqMtqtSYVq1NqnV
txK9qKA85gAE4lsyrT7QigphT3IWrqSdV7GKvEhc8nHt3y01bqQHocM+yr6v+Rm6
n/bcjDuWGei1zrhpEOrcz8E+kqPtt78GnFqbPjd3/zSh2hbyR+5LmGmw5gUBS5Dy
YgiqSMn9B4ydV7bPyN5H4YrTR+h3Z3kuZf7w2FjhIezk1RHwL2A26btwyaAOWFge
uJfo2Rm36gCj1oAbMhPUNicqjAfwZ320HUeb7weckKJdHH4hTqNu1ErGjOuAiBgJ
GjS9L++wgPtue3bKcsfa1JuIAQlPs+paw1reG+wh0Nv9HROWlUUEzIvYIKPRHPyH
jTqpDOB5QkmH0A+neH8pgXls7gXTj8dH9nh6j/6wVd2X5qXzLP8JomUre9SOtD0Q
QH6pIAnaLH93XZBzciMZQ9QbEEx06HEWv1hzyNjdxTwNQm6kBf4yzcxK5TTAk2bJ
EvgHa5jutQdn+ECA+PdjkoMbw5xQODi7P/eKxCYnp/JzjuOwKccAPHlhzlhIEmx5
PR3p1jmOmIuFq/88DMWTguKxFfh8H2i+kHUUNGf7Mpi+GdoypqGQsbVYFaA87FdE
xuweEyKJC2JqDvvnf/lKA43P3rWI9J77wd5TEXJF35jBnWFfdzqwVRT9lU7WbZ34
0Flw9ttw+YuRg5pkEEJ/jUXUZ9JwJ7Wi9EtY7MWlcj5LUKYF+6cIqEFGzSS9rFiE
MOO0NtexrDHQ5yZp974HQBuq7Ly5kvvEFVoJB3waLLhL83tF6cjGm5SCTtZ/WKJY
RHmTIlo6Kk89uGEmCPZVVYptBmII4sC9FyJOr3l37ZeGe120pkhar1oD4J5qYrmJ
xL74HP6aQ5tUYrHcj+IwyjLXZCFdpbhq/ng/CiudilTha6S+pmkQf81ThatVgTWI
cE6hO0sGzogQJA2yGpm3yGupuxx5GIn4Nnccfukae3fHCjLd/SZ1FhKFFplXwiWP
6Giw3hxH/qTVA7MduSqAxPItgOOW87WKAqUpwt20sUI1ZuntZse338OWmtExvGd5
CURH/a7x+DIdMnaezVemsnlmhgZlGw6o0WIGp4mA/mEuuintCD091ZrSe58pyx+x
0xcwdhhWfEMzVmVcRmpFk5rJJzPV++CPSLlgXOURQwB57emzj2N5YyGIlqBigm7+
EAzaFIoZMramGx1ATbAug0WtE0mL7cArR2Wi8D7NFcSY+7x/k23yQvnYM8i3qv0i
Taq3vIp+6XQJejGooxR6YGGFkpWYrXTBLnoaNsqYxtYZKAun+4djt2UmaQpHYtGh
Lm8yIcG19I2/6shuRGjWy1Z4hUfXGUnSoFKhHXoSfaRGgkwbzhEJnY5S6i1gD0qv
fdznOem9GWJDhpMXUO3lR6A0nEgMbZ95zw9Ai2WB9tTZ31iTSsdeNhCpqfgYLn2R
m/frl4avk81rtKRemPlEy/Wa9atHodOK55N6kWjvd5JSKFc+5eZNFdaonmkb+I01
WvDRFxnshhPWmcVc1+gSO097lMpZshqXhHI8l8HPMzRQcSvfmlb2sfZ6X069IfOv
DTIXXiZ+290wg6+jdXQw4yHe8FR/CxO3H+1yXbui8DHcZUN311zcmsKxxtphrG2Q
+6cV4H6g3ZM/ey4LgGPs2O/kBmftOBfL/QUZ7ZfpG+Bx/67Uap3Zj+HTCX2Ie3Re
OrdGxXvjiHFDHg4I+hW8FUgXrY1X1VhskzgQj7FP6k9OZFK6XIvQ0rr4oHObYuOE
P2+zNehWMx9iW1P8ReZbZqIjK2PxTABhUl0NBKdR8RPjc1O9oONWBvG0fG+K+3oW
jZKH8Ld4x9QAWLY1/HQBPeyO+x+MIXLNl46KqkgdXzlpJK6zlSiDHDislIxP/erM
pip5QwG2mIP/YwkGKpcBoBjWU3gFT0Uvn3ZS4YPOlpu9icaXqguNGMbEkFG2BBaE
GASPCfo1uM2NsUOl6ZuDwAu40n8Eb8fg0v/aECGu6Pgj64HWBeqNUYA97ee9r2FQ
uFg31zvkYpm7U/dfqgqU/aO4zvBzCuZwDOm/7U3FLGRKfw+dGurwUbh251Fg24Fv
5+Tddttuq8yhDaKFSgos3bylQb1Hu5CEymn+2ef7jmCdGCcVV0+TsYfYk5Jl/BvK
kwJnxjK09wYf1SsJ0nCqx6SwCbfuijp1mZWoNXISxArl7CFZ77MnEuVfE3YuihCM
7S01fhYzh0DAmdsQwNzj37raBMyukPX/aecCrA6EZRTBtWzwjDJnjmQP9izrJm3q
Ry6safAiJfrhsuJ2AhtJzOjYbDV2lDrGpmHLra5qEHeAUFFfg35SmjpqKIJz8fMk
kz62QYQ/M+TP6t2fL7zUg5O9X3IFLCjrWeghDp6JxgeHJUvoNJL40Tu5gZsaeMI8
zJoCULlwsJkSRgN2Zw/8Ee5p13cjFL9k5XS1FPK1ksuw6vgOCD6DSyIffOoPCU/T
Xjt5Dqd0sOTD2V706WkUxT30OOs2gvjSkAbQ3S4/Rr4IGRrvqB6Kr9Iebm6EJe0o
9nDKazslP3wvTSgh/t/H4LUeDMSHpVDU5rqyQ5YsQiAlt7+hgEPoQP6RHZsjelQm
5Jz2paesVLZDA44DWtyJOoan2lX7eIZEQm+ZMKjIU+plbpe7MoDJXLRlcZsMBdtt
U2VtQEUjPTruAxJ8WbQhAUVVr60AbJtMs/c8sk4K3EPbG8MUss24EcHXKLyvPk6S
p6foRZ3+TIuD5PUPn4VMxi0oeQrESu+Ki/c2Bw/QahWkL/Lbg4IlnmDZLPggLvOP
AJtFIlIzdH3Tm3ZHxEBlKYmA8BXJgb9Sg0WbAKZTQXUkqThyDWd93SP/PJHYWshQ
c9tWsq76Q3U2bCRyWVdRgTqUFsn6UBE/UvoejfZUQ5fRFEIFPcBntxNfKdq/6O+f
5fIZzzdNWm/A3TiDCxpJ073jysFK9eNZ+IBZAjAzSF6oUKrf22cIKHlndyQMMOgt
tNZUVwwXuYl5//Tv/XqVPLcUKQztY5wDt0I5g8rykO3KXdDPPmNrVwYOuZDFTEcA
9WUvfDKSFiWFOuhabPAdpzt/F3We5V6LulbgGj5RNGy7JAimw6pEXm4DJt5aasSM
kIevd/8HNeLM/QZbg8ZehWK4CtlyOgZH3mYNL7DcPWPa19m9b+1Mz0ngO/GnNT1m
iDMsqO9piVcWdVvePd9VUWK+uhRwVg+kzYnY8JUIQZmqreyYlAtu/aIdta/3bZ7q
MdSs96Kan3ltI8A1fpf+CffmDUo5fI+FVdGR3orznd9NB0rBs/TpxwSBwakIKWbK
cFPni9VmAN9sivauCcPnDnaxJRSNy2bjXFnHJtLTgGX6tECNbvcxMIj/N3HjOpw7
6DlZEtqMuL2v83yKZist7RslyM+8lsRS+oS/VykZw4b9dJPG1wwSoxCUi/M9oRLC
Hi7eXjx6cGWrU94XhQCuDv+XUHHeUQcNBTytEMiMcCaZ7yvlZu0U+u4VAAk6xEyA
HG+AIRpd5tcGibivbeSIB8Xs97ekUx6XWHO46aq97jQEikf1vOS5tGSpVP8O783y
2kSFMAO4/7k1mqplmf5Y7gkTMrRIHvU51t1EIXODrmpfiwVMs4LzgvPx6LaOrsQZ
lcEE4mxdH47t6z8S9Rd5QGyb24jpV6j1NdJ9nnL91WJcTVWkYdxraZMmuweSzuHy
NbU0moB5YC1togDuTCHQCDmxauPY1X+PZEq+TcPnz+UpR73zSGzNdOzGxtNk8hDB
ypG87lv7bMqpTpEuqAqKKakDcNDnvAOeDms3y5C5AR5E70DpjEAdWt+jiFdh5Xu7
dwy+qHfv/tskvZ6XSsocIbGIrgeUx7T9yTBf1zt1BANLlJCyCd49ql546n/uVw1S
B95XBT93tXg8dLKJaNZ83/9gGbHryCQv1FMwTCtqendanGQ9YzgN1nDIhIszgYec
vlqqe59TBOUigF14upNx1ygvWUul+C8xnsLQb8cKqk4Rsvm+x56CRTveJKsjURYg
ZDJPTBMxQW1alH3glo1M3iOAQJUavLHMHZvLMKzrIHk+h/t47M45CcarsiXkPvSn
JzmcxdIo5Hue8GFF181/t0pyieIAa2ft45NawxmvXBY/t7zLZkMsuluWVfrCuv3x
M013mNgIUk2jKIQGrmZ8aDzaTUIyP5ExVqmER87JorN+C7zbGoMRiZEUrO2Hu59O
ROFltDqXbkVpsLJEUMgOCZjQ4YoaZjHqi7nZak1LRajkiTQDhFXK2SL4xKzVglCz
ZkIydM3JCJeeAuoTdfbgEoXOOvvpSDO+LlOxWqmPZy2sKk/6xYd+m1uCR7WS1eN3
SXJ/Q2Sl/3u8B7kn+q5kQglblMJb76iY14gUxi0T2tflfGvNbomfsyfXQ/0LbNst
2Y7uAa62NDK9PDkfADTLmuXlTBMim99q5H4r4z0CY5VXShq6GWhMGBaPvrXSvTI8
RVYroO3UtBiA1lg8UW4xla/TDJAZUU6Daowx9BDEzfiNOT0GTU2e9NiOY7KwA9YW
8MLVbn2F46JIOBBmaFTikNUwnWgTINhAETnLYCe1flPiSi8EEAN4A7o4VcsUDWlm
JAPi8N4DkLRUw/4YtuquplvsIq20V2dTPihny4UxQRmFGjZIl3IxFybYFl3Gshj+
SH7OeGRs+Q3hWtx6duT2P2Qlrk4+4GFc4IujmZMOfvCy1n8y9lodHg6h8I/jrA3m
+0SqsUG4+wPFnLggj97U3dsWu8nGPGt06WU6BRFaW0ueiLlDvzhzfladMTiM51ak
iQAcxptGEGPCUDdL6Bx6/d4WtlqOMBGGx7MYeSrMhGW+S61lQuv4e8ZfPicqL9L1
o5YG2ntWUXA+te67MnhFTou9yoV/wtGKWIKBx2B1/SO54u6AMN7n1nDI2bMJZsZL
PhHrxBw3foCl5aF6/FJYqIg0qVGMeFvWbWgjJvw22lhQcvbvl8JCWaKHLtRTzude
nLPxLfDccEuH8qAwodEq3I9AGsnIopCpeEcro5YEOBWr4qGBv7uf6QQuqFH0tvgV
Ct258JzgBK3aTv7ErpkOHoWvZCQufRoxIXId7D7uG463l9h0xtaFrPghz9g216/I
oq29lpCPGE/Ewq5PZURhlKJTxPG/f5VKU83o3/VxLXS+6BniBKu5c9mm738UL9SM
2f3219jHRkG7I4hv28JVCq24qShytA2fRINMxi0VugmzZ13Y04PMJod5cDJdeD7i
SL+F3wVl3hTXbReFEobvYkAAO+8Wy1zPNEufh1npJXIXUT2uDgKR/19Alb/hCax8
2GHhctwI4cV4vf5pOBF5/S+VYG94Nurmmaq0LUodhMu29iniGigdBebde7Ljsrmb
1iCVrwg+Z5LUVmtPUtNqsmh8xWz6Yuq4Pqq3PU6nY1zt5UXbev2VtSo6ImkclDMS
WfaU7QoKsEZdge1kSvxmi7ACsOZhoxfp3u09OmGhUUeklSEhoVkqU47yIxUA5rBk
z2i+04sWZOAw+E7FWHMqgQMpAmNVAKOcV5xQ1M67XlSKlYxv7wVwdsJisftF8Jxr
nF1vhoo+ByC1vu9wAt3r6BzvwSiPXFnvUD5dmxcPpR7JYkY2EwePuLk8e4YOMFdz
NRjdLryDbZhrpcS8nw3ZSjyDV/ToEmUpzav6FWHzQ34/PgfAozuy5XK/0HRRZi76
6/Q03inAunj/M2+Lc0ScWlc1szKP8w/E67ca8dwNKRxfjx6BlW0hLcj9f2SbWi/9
xg8jzrruVV1uS02fa44FkhT0ngOyw5jx2lRJbcO3VjKv/qxvMwJx3+QLoaHZhimG
K3J3doMq4qCt1coluq+lqkRmAlZdezycKZyuJCCt9OZThYYC2MlQ6FgjxEG/Lh+5
vcbcB/ub8gqf+RsrxtLOFf4q2bhKPOfJmJqtvDMKn8/hGfjRhnK4sojstVjHOzZh
1qVeFXrT8QKbnfLy4xVPEDpNZBop63Q4qHoC79RlTU8op/A5Eg1IkS8G7BEnyj/x
d+mzDaaPZcxB9xNUCHxsyr9Fl1DbK8utJJASosScLqMOKYV+nAgk+3JW3PjREgrl
wbfk9wl+Q2g5k1b2hM7fooyukPADSyCRLDvPamQA8GSbYNSqyN+v6mOuMzwIYrrj
jlb4z9wM9XJqyk6Nbj5iavxaqtBGXDMOkJLr6kpcpThSSEm16dwbNUbeWbJ1EY2A
zW89hNGr0Oh86sucFYx6vbBrXVIxs20Ql5DHEsxxOEy2aTNuoyN+GSdeJocmSX54
fMRHdbb0JY934+YDmLUjE27zixgMaM/DCklO/5Wd+RlXKCySFhwT6kSXY0TuVX0w
Y7NFqpQItYMK0QxfwZwTySOGd26hLdMq2h7HDbRkosa6mLUZ7JdiPhWDlJg+QTpB
3/W5J9CpPPvZSEwky7WPGrpHZHLpzs+zvqxlIqw6of9vXOQyXsAkk1dr2st1fl7h
8zA/anuiXMwwU7kWvw0MY1C1hG5llE338Qjd9pL/lS7+gJBfvUel4mW27eCcdNvb
gO6nlUttMXYc3+FZMSMe6xtH6SfTminTu25ianWdAQQS4iun005NK+IhO2Sm6i4j
V1N0Zoai/QFP8ChPF6o8xQ==
`protect END_PROTECTED
