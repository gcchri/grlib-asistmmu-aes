`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TiiCCcKaAS+TarCgI1Mcs4NJSTPLNw09aYUXHu7kcHb8yMtsr7O0WoKmzlgFEvd9
K7tZO2E+jr9CbPLTk4/ONbYgrB2W4zQZfF4Q0K0A5PtBTvYD5lkq+WX4z4A6O0Et
/ccJ5S+R94Q4cIDzJhYA9uC+umcyFCuogTNVxL9X5dQRHNLCCgX2mCZQSPJo94Xg
XOfdeb1TeqdCP+fjAuhuBYpc+qTylayZH6082BFafR/Y6yI99NyswVgg3nHqSjgD
NA4jm7V5Cld0AnLD15XS7wnLyBLp57kq/rHD0oIW9Vx250soYgNQ2CAX458w3qbJ
Y31ddNuVHFAGsUU0zeVNpBZWR2izOKT4vZWaRWihg+g=
`protect END_PROTECTED
