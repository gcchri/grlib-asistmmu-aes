`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pr/1QJAEg/Z2l7JYWg6BEwHMoROFxYuAhgTQHCflaMyuIRUPpW4YZet+pp0weggi
imqwL6648Lf5tQEbJqWZtH5f5e4h9fbr+VK0++YSCqrZuGehUY/jr0iJSIhZxX6F
/w4ZaH3+OslGPTdaCxp8s2dA6KnwEwasRbMt0TQCqg3jtTxEvbXCcIcDHZPSL0/U
bYxofxmBOVyXe1OldzVjnq5392kILYSU/VLTN8l7DyEq6wv1mMRRrljcql6Idr3G
EsUZYKiZgZhOHVJrNZCvFix7bLSrmI3eihlr9baqJQlCeAGtIP0qk6ti82LIIY6/
3ZMXQ1Ws4r/rycEo2UQHFrXQ5GUBPFW45BA/bK50fIXwKOr46y4P+vaeKx2Ldigl
ay+C7xdVhlaHygcHmKNhZK0MZKulHfX7rN/O7j5csyoGBFDSuhj9XmPyY8Fk5vKc
wRtzFnAfSonyLLjFabfw1EZS/MMb8bYj6pDC5ZyK23I0YlM+TZAZ9F1Jz3uduvuT
uPZGqu4UvzbCLI03PASDHlgW256+YYzz6rk4Yon2YTDuVCd/DFLuYVMD1cfM/MWE
B8V8XTM948Er1USwrwu34L304TfkOVN1T5dt66hAl+3wYo+KmJ2j3fUcby+ge93l
dEP83WqDdHI4yfpR9BTSlLaqb7Exh0ElZJpNmYRFTmwulODp9UquV4fKZaPlF5+n
AyooN5ABReYkIcJDC8Athm89yXXYIe5Qn6GSDKHsImMmVGz3JK3DlKxEX8KcJQ8/
9zqF0eYOwdnTQP6k+gwPknV47GPVy6fLihceKn6gGVEofe5+1Peya+B8ykgNww0w
pn5g7m4t3U7m2n3XarmZZYu/Dah0PODxjMwI1Q2vxpoLBZ3D6ZWrE4U/4itl3KkG
wfRPBGMuztD4vv+Tvg+UEm2JFM7OLGwGjHYSDTvx74ovlthnrJKY/NgM0E9hoah0
qakPKToy4pz2wehG97vf8g==
`protect END_PROTECTED
