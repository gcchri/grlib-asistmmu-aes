`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNRW7q0SF9JwfBxD0518us9WsMcqJgx3tnyqJ90to4/1CfJmUzz7YA7NtONGkCcu
dCq1StNClhFS0dwd088NA8twFYyDMyurHDLTooiGqHvqCMwuqm/JXOsxTK/TleGX
WgZiqiO46HyUN6bTCdLddm4dtaMsEN3kffxyv2WXm/gpxP5aMpWLOTN76LTywUmk
B9glhbh/wE/uOEj02vWHegRQobuSsZuVTZTFM6UDX65tIR3yqTQChm0aPuNTPmKV
rBH04NeBM3LBASQxRTkjUkfzVUOOL+uF/90dP8U+5eZELnunzE0tH5f/h97f6v1Z
xap03/4M1qsmd2gcEErSr9kAOfojwldcDQDY2ZFwutg+pZmS5LDLfN8uAvRgQwiy
dZf0EqOFQ8/9Vusj6R3LztNXl7/YWZ76XT9JGHhwnmM=
`protect END_PROTECTED
