`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HodmaXgAJbbQLu28y6LkTUIc5te9xNnBerGk4HhqO9u3e6GfNnhgi+wXovykPh0q
/NAy1lVdg4LG5XoLE3eVmK6Lhicy1tus6CPsZ/oYBujnBzRUF83OnkjrSvX63Lfj
hEqsh0tmXU8rCKrqQaWEzBf0ccfnBJ9QIxgKvJKsyZElArkzWHfRDF8jHYq++d+t
N78eFLS0EROW0x9rLXiBImDevtofsXl6FcwGjuC9hEcg5bUd4WLhxjqxJ+6jtbaG
hh1r97qFhLj0qKUIgsig0G6IMI+v4egUFKEYiYxYVA6JoW6AjN7g4y6raqI5mBdF
oXw/FUMIVA/Pjb8j0G3Uo9yBA8OaZUFCiaylSVDgzMQM6dRo1+KLt5PFpgqqNCbi
ADl9ujWO3LN9kipRn85rjBUMhCDNGYtv1ExKI1E+/RYwUTzhYrG/rGPmnX0EP192
9BVd8V3Gvws97HmaAcxXjPlul8cMTPz/MgaxBlWFdE8nQLkBocsSkclwOvedSXIk
HjBmZQO5B4Yz/p1ajaybh0m+w5Fi6AuQsIiMbY8/cEw+ZdBYmE35TTTxd9hOB+2b
P43ekQl/WyMFD3x7Ua1T7x5z5pG2z2jEhyMW7YwIX9oUJWNZFpEB7hRSrLArrQLn
a5GF1jK13akoz/XHlVdNpaLtyL/51lqr1ylD+m80y2W/xCqfv61kuI8DmN1nSIdP
t6+qUC644lZ7feFbsHOAlt+yiU6SWgPiSDtXSjEq4Wkdvub6Yg7drhgkhOVEFGyw
BfR7yxFTuaO+twUvDUQ/yWPMYuphqteYNo9XxEzAlG77sCmeZIAtbH8ULFcc57XT
HFxvWpP0a4nA7b412iX98ox+M1vGqqgrgDwv58WM0lHyJd/HgwHUdXKigxMjmmCE
1ucD1CEDgSRryCAS+0PNfvIhSGykefl72boWXc3oRYVjEde11d1gArwivc2YKjJi
OUYOEM+Qu32VDKLEyL83HO7KkgwuvaVZak53knGVAtsi+Iajt7sWfXVi7+DZ0mBp
d8Mu4Z1yyrZf3akJshrnh6KgJPsNqTLIMjA1Ae0c9xQ16Xq1fxvmBjNicvR40Clf
rDWWGhZcHpqiPGC2+yvQDsepaIGW9jgm73az6RjGTNvcP6UrXmhnM0EOh5IEuUua
2GdcQqvg8IlrJPTqSI4gD377NsIaH4cbMpTtTeDg68anJwOxPvxfpflRpp20H72j
RlaUUNMXod90hZf6LXa2E4gXxRaSWqoMrzy4cmcWZUitERXnRF6taM3kqHkmfJCn
ZOfkxn+q98vvpxqn2L/6gafCt8a6o91swv7yAbF+b+8L/auaN/LKHPvX+IeF4yWR
JMEswO4ibtMKzNcQCPVvAvt5UGfZpB9fVXcfcVIZX3+HRcZkcdhPhXj/zf7E1wT7
/509qiLMq7TcWrpl1LIR1feZ+T9c6vChPztCsuGDliZNr8HEehu9gHnI7WIKS0gZ
3Xy4I0OwYCgyMtc9nVUkldumaxYC+aZ0cElIWD/ZXUAT4Ur6mrsb9U11BHhv2RWA
RqYKuKazRn1z8x+TnR7oBaEc4W9/oNfFWq6ihu6aM6U+CTpboWqBt1I7Bd0C+hYt
xWcFZlgygSGvjfZduh19HZfVyLoo6EDc6DHLn2Y2RmUtBKALu6sb209m5U39tw5j
fRwbAH4EhZYpYyvkuTaDmUx5PrwxpdzQz1I7UyBEC8zS4Hu+VAl8pnv+av43O9Qz
6h7hGUUqNq7lp4dm4p803E7Omh84t4yvuhaBxz1gK23WU2YePUiZ9BR1uoKnsmO3
lCWw9FX1M2xSWOsZgHhBAp7hWpThxRLPXKMtOrSXPMeeoqc4w1GAoZVMm/pUfrjH
SrfPRoodzlpfYRnGGD4PNN5LNn/ilwkWgkle8vnV301j0f9s8tmeivD9OUwdhO/H
JrzqOHyrtgCx0ca/uhhKaaNs3sZbanX4MUfOtBac1Hplk77nl5DcG8f/4y1XRavr
EjGvZgA9qhcgFD/vUy7pCLVv4zFUFP6e2FsUYo/iZEuouIDBmF5YwGblGJE1GOI/
IpaglqKEvP/9btTXYsigX3X51RaNiqwKEIr9ueNQXrexp+V4CQqmky+seB/aPTYx
h4J63DVj7OWzaI84YLCUZyF/3YrQy9BcZPU3R23M5X8+o3oc4mhHCj5kPaW7nL0f
9cxtKpoxCX2QzYe7/Sa0e7i/yhGs5YHfjHtdXUSllYH2mKYU2q4emJ2rSq0JXNMR
7CPN4e9LqdIYH9/n3ZPYVg4m91XOwiq7bQWqBOyt8MlAk4/RGBphy7vquTr+9T6U
yKhhlJAmgoIj9cIJlCoNzYxmZ3CkgsIGdp0mRR8Sc9DN+y4sMArx9HIZ0KdsdEXu
9/ZgHpCIk7xLVGA9+U7CDSM6haJuc4qa9tBZkoud6UiL9qLWrMBWwSicBhdS92kW
zXANkT8+xgwMzCNq6JkiZtWUyzHQ6Jlx4nKY9fv/cZ+JoaTWwi74GQZ7e16VLACq
RwjGwEfrawtDKOFPHS3O+fcGiG7LwtJ0rlsASbFO3KYRT8/JUt/uhAQCTfW1kabu
LnztjOngTQFyXjYtvoBS9uVJtXi6j/ZaoEifyavM4Rl/erImXd+sgC1sGlNdxncW
eDnagbYNFdbqSQ4dX2pHCAzKRjpYWvZpf72PiaoZ+I7cIMugiv0PSDx4fFzJAEsg
TG5UDxjQ6Df+V1e2oF765IR9xn3iDy62iaIW01ad1fTMyCzTXtsqDKE3X80sqsaH
dGwbV0msj+ect5PgR40Hv6qvHLmO8FGj8e48n2WgZUJcQF+vdWSp6A9XlFmzE9kb
rXV75MLBlXvM6pb9+PiXe6kttj9o6ASaXJGQYcL1G0c+g7hJQeHq4Y34N/o/ADfm
ALvz77ZwvKlikRz/93rL3F4P3xWNaYH1gimWUB1eAxOK1EZtImRg0od6hwZF5KP+
1GU7d14bFdBiMjX2O88RzJDi6BFB5JP64Ck8BP674FITf66U27I3IE6t5YwRvjt9
j+DeB/cKlgCPL1Ez1aU90KrzW3vIiHyfRgZoujvFAUxir0bRyaao2nLFF2CZu7U2
J++6Al7j5O69VBczGMIizlHsBWIUtvT70y538lG7n2GS9kP7e8FOahH6AMDEZNUe
pVc4EN9rm+J/vp/QShuS255ZKZpwoTdEZ+BH6UXuy8WiR27xweF69q0ZRnURc+ys
0Rnix9usSqnHOPkGjkK36FN5TG9Nq0bZ/XmzJj9bWLxkSj6io4rV4JUsfe7C+f7p
NCITLLd4UQQYHV2Rb3vyH5ErVmgTvZjDDErk7mDDTRS7fhKE3NF7PUjoXfnHz8KX
SF7WLDOCL2VH6lRhIolnPLSOyoV+/LCU2amH6sWbA5u9+0fBG5Wv8XZW93kOLnhM
YjyMSaAzMBROh/GO7syQo1un4bogSbCv0+tqC1vtg6gKJmD0nyMWuXyhvpytp2B1
TTcngnZu47nHz4jhb/KsZXh9ES46D76t6fUYeMXNnxOgjBietZzbErzww2voy88h
dBW5ZeKbwUa71a6/068wo1GiYbfudHYQJwF/I0vozdcHqv9A2sOo5HjuLcTZzsA+
QaOv3x4lubgnXgJfM01SRiz7CtHWboUOCB2C3Mm+mmduZDh+loOqIQsA8ZlhYHSj
kpJ3WoGYk/VU+vM0c4ZdN2nnSEGSc6WkqczFHnyMBw8XylEsHKMuH+t7ddCkl1FP
dcibR8pVPVzrEzyQVzr32x9S+/a/AbZCggK0K8HKcbw8IYDTBuZJt+kaakPPDHIN
0ObI2PVnNArdymPiyu/eKhSARDtrnxLU2YiVAYBLBnlne3dJEOyHhhljEPCIn6Lg
LWpXHn6gwpLDG+YwTD57oILJX7s9fXjeJwnaoHNlc2MiiK/Rbu5px+ORd6ttgTi0
Hj58EogCiHbqt9u37d4jZXocvXf8FLUo44ATEOv8bmxNhJzYOUYh9gafaX4KPO+C
icwRaQrGXlCKqvnagU9+vd1e4j4g8VPyHPZlEUByO4aZ1lb0baagQJ+3y8oFGvxX
65rLHA+i43IKLPrXh+6PnrznNR/eHbtzV3cPhIzsF7J2T69m0kdKnuvZOND8oXhI
2LV4Rmej2YEK5F74Sqe/gE2BdRmUdVDLjuUwDvE+78/MpT75AAAdAf4VEvxmmOCu
ILHQ5QjILpkMj6firDnI+B3PYDCpgOJ4KT+PquLuX7198uzwTxb36zOSjg0tViE+
NTBspO1hiRa6Uu1pwRXtA87OCOiQKCCcy6GOowXUbc+8bqA073CXHfW7sffmkQ83
Tfam1/5PWLMB5RVS6zx3vNqU+UXnzhf1LttMFSkceRRFGV9KQTQFoZPiXRAY5UGu
D3A4CEz1LaSNa22MGxaBwRcs/sM7GivlygZIB7TWeDJKlzw4ZGBcNatdLS6oeAJz
nl/kKKAyOKXH9GRbMnNgDi4umvJ7w94oARMqhhp7Fu8RNOAMjuXnEFVlX4q+OEbY
rK0xxqwGkL6B1ALeSPfYYuI87CN8h3mMiYecyloCVUxCBBi7qSjdNc7toO8Fim7s
sU/NCcRJvAoI9udEJHBxWrhew6bCprT/XG1UxHIrTC7lmoDgcMqpBf6P8N27+Vrh
5/kEB4Mp56ZPQTmVS73CR5FZz+sVxNnZ96MRA9qeXXctEEVd/D7n0WEg4pKnkDeu
rYbZXIFf97tUDAHWtnbcCgpyd9+9svX5E3lHx724svO5Z8SM33AzcJku10dM/sSs
NSLgFw+UXXg6CFsb1/dBnh9YcsDD9gAzMRBCPA3PpxnrpLJiNLyIb3ZYn0cKBBzz
3qjRacdjGOqiiNc3bVrvFa5ravZO5q/9HlNQ8SzKqgLZar4gFAOrkplpAgOBTSh9
rs4s5enmEnzul8ZkVxHZoYsueZERoK12U4U01/PRmxcBbW96XaZhTLccNjcQb1GI
5Fsok1J0ZEc6ahoNtkeoniID3mP5u2JHlpA1rXuG69J8PQoxWI+e+bvcCzUucGv2
7PX4TJgV/C2srJM924psLoLFg0CArSadhnguQ1onUZmTQ/GyShiNnVsMkUtj8wHI
Jc7ikvh2huHXyOE2Xr+LgeTGOjubiESYg746dsf79rwFdBe0vubgkAukhGFZkl2U
/TApEwLWXwYOJY6QPIxLrlxCoj0P/r5pBXUwtdvsbd1lzYrkSFyy9QHcBPvXtEO4
EyC9w6S8RlSAgXBn6uRsr+LSuBdH8zeH6whxUC5QsM9BrO0XzfD2Fc9UDTL5XM5I
VNP94RUScfDe2cZ4bNlumaEqIaEY7ZOI58K8QrDOHIsI6USmA2k7fQ/D6mTvt/kg
qmjBXSF8JgA2vJ/iCklOO2RgpbQ7wzyUlLGYPgO5ouHhpScOojavdt24hq1PxyDE
eECD2I5gnewfMN9AF2K5pFZvxDgjusYgQu0Qrm7n1e6fG+bKT7nAkYKsJ78h3P7b
eOqDW7okESYPFlRwAA4+8MLvCIDMRYLMJZYmlEb/+PGCxgRsRp5wCwaU4AGQ4Q0h
gafOjHovgc8fQmyAnQojH2KW/QGywV2f6LY74kPcrob4BaR/ML5LmopQAcEXkuzB
VdsrrB/42V+6EvKJ8z2c5miO9rL+aaW0X9O6Sx2lUFLGVVe1IFSgC/xTA8Ybq3oN
S/qB3EMWW7OCza7NVCMTagr6rK1dpW8pygXGq04frojWV4qWeOdsDeeH2yVPgmSp
+9WKhnOsf/rP8FNcP4FybebTcv7yM4yACdSzhU8CmoEYhGI7RLgVtxHEgzFzCbEL
mnEvnlqSdkA+jABocExWIbslW0Y5fxzL7KIeetwAlLvB5+q298FxeYBrIzaXONf8
mLMWi1hmKq05YUhk8AD4wVFx3Kecuhm6DZW7nqX1ejaI2OQkxlcN0UMzjSQZOvSN
F3DbdYAljcnA8sFFnqVSG5OcG/hIx+yZ4TlYzp+XJyVRqQ+UjeyjWwTiqFJ8Rqsc
fWcKLoIkXC4utRxDJGwcY0u7QIlNocA119PPlv9VYWDJs4e/nzR6uzS5FRWe6cby
W4gKz5KGWZgKsK44yat3BVIjkH70Bg1xlK89P+XV/NdaCkVrScRhHtfRtq+k65tf
3VGdGWqar3wKOaTEmDvVRiwK0fm0TEdgv4NbcDDB2Zbx/YqFgT3XUuRgrb9EhqVJ
zCm7GSUP/Vn9EdPg+eo0RucfcPzYhAEthZ1oTxaTNvNqBoO4xIjFJts6/zb48Cfk
gShqGXOJ26ybXokmzKpFipZ726seK9QkpQYJ9E6C/IssMAjT7Lay78RSHN/cfpHk
Jl+JqdosZMpKToV6SfxaSMPsv3pR07kBlhKa9Fx6yuPaVRu2xqO6V+bg+D7SDbS5
poeF1xDI7vNfqu3+keujIorm7vFw/FuWTY2IxcRILQAV4YoJ92RoEv/9RZ8rTF33
RRrLxY+W8oaG02/x/Z0K9kOSDi2cx3j8LmK35DQLXtHzqN5hxA+yetsJhNO866iN
2PcZT7trxfkoCWQtlo5d96W6JIbHWiofoM03juIH7ou5+08auBV/Ib6fBRiacN1R
OhAdXkZczpS9qfDlMTGiTrKyXwm1ViZk9IZVF4HofoBaqewHfJO+aK18nQ83sk86
EEKp0705t6qnldIMlExBpmhB3LuQ+RFMmhhlLOvHdCNKCJPKG+MNRdssLih7kmSF
eQdB3kZPKYahopnBbwaeJksxYA1pMPeSUn6B+2d/svEjo3Lz+ikvLq1LTYcrI5Rm
E5fBIBl9oJmqlwsJ/pGT1dSHujzewXQrxlcRgag3O74NstirWWfmc4dJUEtbPDY5
XnIwYChdtlebRkDmxNiA4oCxDicznxwiMPacUs0Rkk+SitfE2+hMUbO29w9LvizL
Ik6jU4nVlAImoxkVNSNSU8txOCcJUMXekSizy0CwW4ab+KgyY2UM10VXW5zyeNuw
FjJBGzXkAI+CZaIyx7dUp8CEgdbeGupZOuvQJgGQy7k/5XzB61ynTM9LewwT/XL+
VXYRKwxDQkzFjbdmzFLHJxex/2znDQhu45paVfasO+IkbkaNFabecQmICDWfd/UH
ymzXJiZhmLofHHNZj08OlAK+biX7RfMm7L4ZKD8T1uvQ8Ig+AJZIcgFjFfl0iM2w
9LRrVMTAVjLgOwKG9Sk+6Pf8BUOSh2uvufiLOtdCM7baPCUB3gJQjrOci+MnfJKE
UDAMsWhpUUlGSfs8s/1Ai9Es/BOCUya1eRrgiGVrQufzGBjfmLyx9wvL0VSLkXnX
99OWh0ujYn/X8yXBH12KqHTBfan53MfIV3AtxC5zXTYAv22+tFxQs/oPAcmwJR4k
OWj1iY0ggChimYc860Fg/LrQj54HmD2rgOUgFCHMUkHDkR0HeYXQRQ3kTjChj1Cj
JXdtYkMiaXt24NBwUDLnUc4I2Rzm69B+azLcBGUNawjBsxrhrvgkqNE9b07mC/V1
jHbC7EgppVBXwPSGOsu99Ve8Bclau1CBRqeeWBGEh8cZ2SaOXIvIO0dkfOvHQQmp
mha/XHvxGXpCbjAWB9H++sfI2aVnJ5PF46U4PaR0RKGzVdHE5qEff8/geYN3DL1Z
3P058NERHgEpcSKnf5jU9ilE1in43TUNg6iLs5MRS8rabw17gZwE3nlGXc1d6ovd
GIBKA9wEmgwJ7EKocQbbHm0UgNscmUyNToqxYuQXIWHhAaptp1+YM0AVNNPRDn4H
klaoitilaSGx3lJf00W/p7JBvM+vzfMoR/myjljARkhFQ1nrm/I6n0ysm3vlS1GW
ww+lJVJ9zXrBmwk/VAmCWzLVS3JOISrPF3UDrwJmew9+tJRFmL8LwKlF8RZlAVYN
PEu/OOsF2VRyIIDbEyKUSMXB8c/ttCTapJ756LgQivuJ0oMBp9RgvsDZ+RS4W21m
HevKCMNzrqwY8QQSHTZA3MFExGTMXQ1PapWy/Qw1ZPnCUPj5rP2sfB98JWM/Fxjx
g0iE/0SFr7RHM6tcnzjhW6ssjPoTi8DaHSMpk71MqbOQPr8WIcp6zO1bATXyB+kc
wAw5uUhmrs7UkGLYvoSRs90UWxd7HtrpXIDDcPXs5KH7hJ+wE2K3XHKMjjsSc7oh
fDPr5QgZvl85xBVJlPAZYB4e+gJpEy+RpQtjyBGgdzGVay5HS5hqdjUuz/zmbJlF
53FPgiojF1TenKXKPqrfsGrWCf0r7Qgr/Oj41vy4+Y04CJpNdm6yhTQ3kW4lu+gN
o2hTYSATN7DHu4R+8fcYrpBnSwgebDvwFUliARLG6lruSS6ScpAHhx3qeDku0EfL
ayp0RFrXI5K/NLdFmkMfv9XD014LcZtL2b+eqQ4b1WMyTuQI+TCOITz+W7W7d9Ty
SQlXsiL9UsEeJut0ph3MzVvSUGAMKLL1F0xCVcokuhvYeVF+8U97hwumVKKflHBQ
gDI9gA9RQcpdahgjC7rl/4Egxv5qEWShbj2CYGl1SdP8VHlh64mUO3gQqiX3oa0n
OIVd/YFMVSxG1Yoxt0rlR5WdIGkC9I8qqithNHWcgkBCCOSg/9IjFEv4VWxFnA5C
K/x68tJTVSK9m4Z87UoVWMjXfQbASnKEWYtrdrwnLgK7HSpQO2eO8EbnrHGwJ5+n
m0zDjAZkAc1kYzLOsrlaRqjV2FkU7u5yxDnGfODyc83m6vozH2SrcldYkTROT+YS
o833vngq3cQDXuWWRFFg8OaUFjkMlOa+EtYxypI+BrGJkcrrp6Sel2iJGcP4tUU9
8ynDMIsqUWAsvBC4n6SGBFycjADigtyclbCeWy+xB+9glL0SFl6MoDa88CqGdozU
6qpUf/SvpJEDJ9R6I32DMLpawXgAza0CCZsRLVemgrUP4/qEaWeiKLli2ykHfSzk
icBrH3CsIin3Etu61uP+ilPTx+LH+TLJ0mCEbUZhK8Tpnai82MMMaiPXwedc+XyI
DMieglIfvJcBxeUQ4WyEogA38PPifWY+0tqOstm5rwxi77eUo8jNbjkgXxGhTxF0
xw4DNaTA0r12OwlvQE4aoUh2gd/4+/rPGbe/C1J+uttYH4x4JnORdI1gWB4hpkiB
UqHkgmqL2YiK9OHVPsnAgI/NSIiE4YLPJEqPUqUxsWOO/8Z7GAYAUpqzt//m01ml
2+Ix6/OniyRaFH3rbF3ON8u9ljCh2P777zD6/xGv8ofeUoh7cRB1d3RzIOS61PRO
A/7hzEaQzT0Oh4IUNxJcH3bReIdezZYqnv2QvjIujqymOX6Ez7a3IGlOSgUSD6T3
OkgR3e+g4b+UB405GyLlAlpKMnyeFmbdCwYvBVzNq36zpfqEd2/a+tRFwa53iTdH
Kb/KBIhkFyL/wki37g6IecDNKjqmdV2/lmnN/dG61ARwRgT3bDhL7ji4NMx+1NLh
8j0aNC3kXltqWwnGjeWlD4BHkR9ETtzk3zf+BmrI3q8+afeQb1bnbsfMoaD+9wyz
VyLdpX3q+MIPomFiI5Rxi7ucZ0O8CPsK6jcriSlP+9BGzWHNbhW234B1WAVI9Ggq
v0XXeX+KMIvNW05oZ7sau6J5tyixoaNPW3foH8Bpb2WhxKjH6bAQ2NGf3F8qfGgw
9mhk06pnNVMOhUKwTnW7Z0JeoWOweGrOnkxhZ91WLaknT445Kdkp6OxDKr1aOAEz
ZptHoebozCK85rNZqjusNN5Rdq4KA+HmqkwEDIiXtHDUSuJrtVCkeOqEJuadliDA
3GLKIo13/0/DaTifU8/4GLhpkdaprUBkW1+FwIybTYEZOfQc4yuMRz0zV9Abjy9f
DxXRMhKTy6V8m4wY59eUTX850bM5oVCkzFsWYtxQZe0LJrBnpse4n9vu8XR6HACR
XlTlGf/RBaqJvxeYSnuqll9/0F/mogJh+/w2NlAmq6qZuCcMLfJ3vJkg8R7jTE9C
/m8o9Jc4BtBRaMa9h/AmsWbLNJkPmQiSe5kPAFa3HwpX9wiNDzxk87vMbKM+nDMq
cVgb6n34THVgK0RBEHC2Rz6jtFE/EN7nly2FghwGb4xx+PUsrkZRIMBIPzkiN/72
4Iz12nRHbzZECDfl46fAxEJtuhehdsqBVT9nD2fMql4d+aClO1WC+SkyHPuD8p6M
ez7Vdq150XPxlxDBh2Q7Qmg6Cebkep4U6kBEXL4RjMAdEz7vDRae5vkLP4KVPjRU
c7u3N0zCE31PUQzTvVSNaCrNPhhOARwlZ675nAYZXQZciZJ+mvEohhdMX/Gw+f/h
9CgH4h6GTWfsfRbS6aVBRW6KD6SI/IqPpgn2CTLtDhy0JYm2NHyRCodFzK4S1neu
skmtD9aMJFjA5mEEEHuNGCKwgs2Lb2SjQFjuTz0MLPiYEf4WgI/mL5p63mdRLeol
RcJCr1DaHwUmiVV2ctgDeuHSNa0lAAis0hobrwDB1Hun/9h3uTvW4fMRsGl9Plzb
LdgYMfa7MKhZAcLQvXhi8Db1IFZ3vOm77qxSV+S3EPYfgvjlriOuq553CSK/fVep
GP6EgHju5ORRpUFBo3AC6qvyNF4x9SJxOoh4PgnUSSJNu3gJ/V7/8WrInSBQlyLn
POyzSHOjGiumbb6mBuLDqjEDttpM3kMpSM3m3HgemwmiCxMbTj9XtNWKT5uXaHp5
ZyqDaKioYTOPU+mpj6YnH7igEYnLfYfCKFb5n5kIbqo6NSKQnjXxqNqsN0e//W1A
RyHieWAI1EJ9o41ObQJbg8k3b7WXRtRN8GtpSpBM2m6F7YGrohgJwCk667TgProb
q7kLM8OZ9EKzLxWugCuxbtlV740hPZ6eCBdj1LsZpO8CGzNuIPLMtdmdZmTrbflv
QLrUP54vOSQbxSGOD/TTJ0djwueqxYSaczhQ20r21jFOYHOgqiCKJkcTo9PO3obk
3KPGa5u7d+/h7x/d2ZZp3gDKJjfrHry1r3KKvc8cJ4vK34qx+js7Wp6Bm3plW3us
SQcmNO3MSHeJkRlHuMl0TMoKZyZh0TW9jRaoms0gIuCvo9yKRWLHABP3osWWIB5s
JrNS897ZTXY5a+l6U3W6JX1QU7HSnhi+WkrNYZXSwLpZUqYDrr5pAvyjBk6d77tU
LzVOV9i1YVsPyOEO8bOXueXd9hm5R4qfzgcEKYTNxCpPk4KaJRHhAbZX4bkxrgx/
YkjM2+8mTmEOdI+e6+XiiO/hXfWoWlRWL6CVnrCzfSRnOxAYopXcluuc5wMbd8qv
mltb4zxdepV/F7HNRrfsuOib9T70flCyBD7swkiN1M6Xuas4Stbke9wH6rcK2ov4
VOC6qmay2r84MobMCNTtZgqW2qdt33gSTljZF04/YIkVPYiF3nJv0TwWXAcGSyYJ
vPuSlGJrMFJMTNzQ0la45mUNulaogfMY1R4jvcrEhpgrSskK4pml2K+JQu6ZX+/4
haU0UkIh6Jlk/RkY9uk3ng0ZO7FC35WWUvywrZsgoOxcXJ33L4ueNKx/2QDPHPH+
+gidlrIo10f05F/FCsEIKzr4hFifJtBsl0mvM2pwLx2XiOp5uSf607recm/dORJ7
8poEwqMyF/seizfG+n5qAEtpQLaYIeGO/wbLy54W1AL4aVr0vzPzJD0dpDDl4Ge5
IUwYrOEXCckfr/A6D0QgRypYOX8C/fj64iF0esLxiM8wt2ltpNnVTlxePtsdYPD+
uLiN9zqFwnLCmRaraSYokgj3pCEemxH3mUSB4TBsj46Xrz0VB6WbhAATpwxXm74N
gz5T7UdwMoJG+TctudOZMOQYCWi3Bd9DRSaAya+CIYPH9mLWByFj/qEHW3RSJP+v
F73vevCEbthqndy6MmbcaZLoMFFQrTU8D6PgpWq4QGVp/LNKuIy+oTiwg8MVPBiD
wa13cBfaFw3uTlesDtpN8aaDug5lya6oXLRsxDAY+anjG40raPaM1OoXdluT80as
H44+Po2AFnQu8O5TY8qcd1wDWOJP1cAwyotJCIpDj8Zb0RTFj39y5eiYM68q5cw5
ycTHqePS81YbxVZhIqF3qfZPTs/biOlKStiG6js6SvkEyRXy839MQOxHSRZLx9Tb
0y5cecg7O6BiVcZQqC3ywGFmoNHNxA6usrFH2OyB2nhkCPgUZwVmllME9cDMCZ/B
sTmeTi+1/dD3nsUAe93TP6SXI4m5Iv3bqqYOeX0Bl0bCJgtmdXelyVa4CDGZgqH2
oE7JeCaR3WJmuO3AORo1ppraSgoa6zBe4z4wJji9YOiNt5/g1D5/3kqbJ+cXrY6h
1LcszPmKcvE74wQZWo1i4ZD+ujbTd6fZgQUmFT4Ob3t4hAu8jsHVX0C69iilNwGa
EtuF3pszh6sCm62qiK51nZ9MUOhongt+DsiQvaq85893VOwrvz5pBnWkH6NGFiGj
N1MINVP/0FSAlZldOLQQa03c1WeNodYsv1UnljXMqCsE6H0cKduB0zcst8OSCSYP
22tarFJaCDOPed/rWBKbqKImOZOvnhGMZrUyl3iBVatQwkqCRdOtwcZA1CPMdA/V
m1g+HE7ejP36TC2YRltatiKt2kp4sKGn1nQMKgMysn7fHZ+zf0YcrRziLR6OKs0z
tL1OmIzTtsitskx6z2UiXaJp0eshhNpTXekKe5D9bOminnWH3FuxQ3MEAfNKf1R3
i/rk6CfXQ6Y70/eoRqpxiBxPx3Q+Xu7pvWIkRhMHmpUaLkOTfiPTV8C5og1N7HWF
n3SpguhzEK6TlinOyvdLBPO8n7t3eTF3rPCV1uCwgo6bAV9E/b/Tg8oajWwEjuay
MV9HtDBl51rJLcDJNOYyfnOIDe2EOCtZ58OynW4Ny+riDPzOmEreAY/R0Fb/450m
9ze5Y5f6q3/FMHYTps9SGpd4ucnVo/eXKsVebslM8GzXr/fjsJnB5+gzPxwci03t
iUaFG/hLiM2RT/rFtafDklxIi+5L+HmknCXg2aLX5IKGhEOaT2/P+mTLb68jVtxm
haasSbv9iTjm3eqdpf4UcgghyFc/Tp1cLFFarPdnU0QV4nbtqSchrZbUBR+IfnVX
sRKbMd7vUK6S1wg6u7TxGReiIW8ICjafXwAZTraYJ34i6xHPPzc26/Mf0XBOLuvS
FlELSyBXD03Q0i6cMtiRdkdiBlUOcJsQqV/fqX1QP3MawYOlXivR9pKJfmiktp+l
5PhDtfaDYsXHBMpv+eTPhrLi8l8OXwaJIltFR9cnmfGB+YSjFFnZEyCYZub4HfPo
5j0ncN5bwxpBRJdX5SDfO97eAhKRgAn8xStRDd3/31Or41BygcqUHeeNxoYQZVIU
TZ+HCUrZnJ/uHooOrFTwAxruPnDv2Wh9uFL263ocgRoW5aryREDGE0prqDHa+GYT
J8RcZZhYqu74hmASGZsBMyiXWTlC5p5rElEqrxzOC7j/9N+9oJhoXwjr5TI7QANl
EgYw+wxgUCzJg+H8AZLOPPSKlZp/oiHLi0nROGtjC5wolF3nlNO+1rrb1ZaUEBN/
ERDBfcwpqU6PdbDq0hP5MXDYMGk1CWK5h0GY01q4D9ja1TjdWcUOXuJkJD2kGoKa
tylgKtQTqY49b+R0Hr+IbFY34u+cxlqJvH6Knro1yECrROVxFYwtQrhH8y+kz2BJ
Z2xpOC4EQvWk3Rza+cPUYSXGVH3EW3d9zqqcJEiPsWkpRuqN2Mb9y5uRDRaxXC3B
3LIIS2ZtuWFVQVNAEkZBfTdtMEq+FOpjHwhxF/d1fqGpJqasrGX+WT/inKMUDUwz
l4f2B+aU6NdrJ9UjOK3kHxVOjM3hNjeRKFs7aMenu0X6BRHOdyRdWzWRPA2NcRcX
no/invv7g6h7/BFSP/RZjfRFjOkldEOEr17j0Fyff/r3iEBWUnUA6uSD2Bwd9azy
jzGBbB+Guuf5ywBhBKofb1m3+lNIooq93sreT/92x7gX16Mz+V/Fptj7NBqcpN1W
UniifPfvausYJRYQ2oG5Uwt8rnBkD+JCZ6lNEOykmUAC84bHmGfz8nsDmhtHnGbD
e4GhDPIjZrOSgo7HFCMMkaRUVZB87JcE7CdPTzSBrZw8X9S5tetBJu8K7SWzJNm/
Zu7gjCkL4Ka2dWEdNZHQrYdMQU3oneK5YdZLsPUyEl3qccRgXPIDnDNVxYFtqHW+
qEGBC/5Qo1BhpzqwhJkrlSeWfjxkJbBaMdAL1RrXPltDqrD9CgEAlvo/GXkYwFjv
hPW74/q1IF2Pqi1z3thJxANtA3e2HDtvfNDfjXfHyuiA+3lECMNcDumflG+OWdpH
7a+zVmogUhQWgd8uLvNlrxppzEMO4VtjKrMVTDX829/I8PK3Z3OM4Ksi6c+/aC3x
54rtcpBywqfIxkr7/nTbOCNtZfC802NYjoFRmnK6DmC+tWG427KWpA9vSf2gglvb
roxVKFcfLFkJH0PLxlU8fzhEhP3XZB2SlbUFmS34cUkWCMTLDOuq/JRtmfVIo/1Y
t16Zlq9MuR+R73LaluspUNfXLsB+aW1Em5Fjf6xAaCU1o4zjVzKqy/AREZIs5m9M
r3cha26+VtfjJZ9ZjcPaZkdTG0rQvg2iGSl55eAwQXeNakf5Q2sLW4z26sC8umW+
n093JUv6kLme8ntJ1DbLhqJULhZZDfBYsxPdxOL85X7DQ0NRo6ZAZVB4dPk42FxD
LVuAgTWR/6OyyQa1w81kobcKL+kNpbUYvLwVdoNABN807OamM5vVX+QML0dKpf2Y
PYTmup9wlcTJEyZ7fSVB30SvQvCYFZ+jVneBrokRxHuptFEPrWs5QAQ7JnyDZkr/
uylXJ9/h1ZSfuX7WJiJWglVM+MZ4Wk48Lhrn+BRNgN6f/bcEqy0ZyP9/vhBVVoUs
Lgo4YJ75QOjfpMTelD3BQ2hZOUUgOv/ZldLBXumlm/yy0Ig5aJTx2Xv4UDV3Lwg1
g20ACpmuiX5ALAVh5a1TtUjNbeVAyd7QUKTBGuYGEIPsk8aoQd+hi2GZJ3lrlY4p
P/pFj5YMyA4/L4mlXOmsxzsTtE1vFi/7pzIdFJmPFc2Vi8xCLaDj0f51YhomacKh
MdI53M6rQ3kZbzEzah0XtA4B0iKHMroyWQ3Vb5KCdHTsBalE6DPZXXegBVtkNR6W
jfpXOz4GXGzwGEIYqRwlGZKtZ2IWPLppY//8zNKOGud4vWb3e2jkjVb1TAf+rOW6
p78dWiyMsUVnAw/Q46ilXbpBuI/AWl93PE7r2KLxqblsBR2UvzcDisvx4875ABlI
X7xXa/Z1XAqb/Waxrcu2drMHfXN5Zuu5Q5eOkejK3DFdKsOEfaFUrw0VPixPqKW4
OxBvZLEM5GZ6VYI8zSSpZfjKeQ/iTe7TJfQku6dutrmsN+ejHbqZOV7qODnqYGKn
UqRJX4/J9QyJGs6KW9uMLgwDCKMpb6ebC0oyamzzptNmz1vB0w3iqSaUcJMe9qlg
dWzavwzpQVJlZXPos7nwuDPlMmgsmkwgAJRkJut1HNc14CdKGMOGbzMuRftVFjNH
25zmOMyT0Q6hPH4q2+AeOg9+uMkNXhTphzsqKrRelT1gCFq4xC8HwwhiMbMbhCfn
EHTzxGW6pGh82bSQ9vDerDaJ/MSvjLQnxa1l8jX9PcvIljs9SbGyqAxGT34AZe0M
MwpaMmxtYVizg1TSd8ynA+J3GU8621Ne6j0A6goBwK0NV7dX2Hv2o0THbaVOnuHP
CWyF50YJmMywpMDJIxxl9rQTkoNQOChWd4nX/TaeL6RiW8J8uPZlKf7Puzn0IWXk
b2OJTkjAlfSFz3gCTYRgKMWT/A3qZTOZdbbbApr7axl5GQbY7O7X/KCZ9ahjrooj
ucTW3K9RJlCRd65R1sabQrktQZbEmCHt6Fh1hz3Q/05+MMISdrtemivyB664oCg+
zzvNaEyHo7feLRdnn2lbuT20sn7o9uKeEdxHV6edMyENIkgcaJhdeJaUZDty6iJc
/iThzUPVWIV0HRpny1YpKy1UI6MVD6TmYwGLoBNAV93kXb+FJkoECLPIXjt6K14Y
k2QbvMiLSZxGHyu5uCEzxsyOONmIBVDoaxreGUW1lyE3ifjZt64kjt5k6XOJpovh
yU+Lfc85r0mAMuUU5UA54/xIw9/wCcKE+9wLi0auIXbTq8yNWs6j72Z0WmlFxaUh
AihltcpNW6TrLm8zY4CGKgpHUXRxoMuYcf2om0UUV3a4oVlxhIKimF+6ytW1Uhtk
4JNrvQ6Srv67zE8a2VkH4FEnRB1GUz2nEANrmT6u96i1jNp6pUjBB3kFFGkPA74E
n2WmJUvZYQhV9unU5tZWmDy8hRzQp2OggRC5/LYkxEZbBUYyJmSXJJbZ6ZG6r2h1
CssjyFIsuwUG+yAhJ6alXI2fZY3EgnvAWdg+PgwhwzvjDHO74A4Jl/xCye0D11rZ
psP/hIhppJqpHIlafsF8jomEpKa+Gu3elg0O2CGj6oPxEB3qJxGh4hf6rNOuquKM
aVQoKW5+sciTcIhDHiB1n8Tj5rfEf7qYvL6+1NIijC84bhfp9tBGa9fT443h4flx
DQre10qtDPv0mVL8byGU6h4IdemDvEVyW2HKRKGF9bJ4jMP+BJ/EJyJBiY3jkz1e
jpZeVxHwgTwrFspV/ehqZhdIhexV7i0RA8+02lRQVaxA3f7yMyzs7zAAC8cAxiuz
FT43BGS3sFcSWU7dw8CjY1yXidmBKtHYZbSi5xRydhyLgdPYwBhaPfnnfBkv+cb5
hJpn1eCMtQpeyYTAXRYRR6imu5ilbux5rs8gmLugLdQl43WkXr0aOkp8otJR5ZGA
G9bup1j/QwVtelDOxsuGXWH4T54VDkU/A3LPnQUCukGxfsTctO5ahBNbFfZHAPog
bDU0u1q2MuDa8awHLLZF6XfKaJHHYWdqeMw0uc8PspERaOIr4bnY1xA0oIp6MjnS
nWorRUWi4biI1xGvzIw4+IvdIK1/yHvLuONXZaMa19YOURqY4TlbyR89bcWtkT9b
8q4/O0eV81GLyjM/1/QCrEAWTC7kAch+P/L2lokgV05dbV9VBUQe/ONnZgdrSl5p
xOwPw2gGwSkbU6K8DEVjaYNv7n8TN4V8yGjeX+Q13Tn0MlCdvU4wQQuzBWzmj9/H
YjIkvO7VbWdnIO127qKSYovi2j+2e41tpDhBITMzbWY62LTwRncJrdod6gklDrpS
CGJQn3IMkGktuiPBvi7DUMDa9DWhkuKGs2pnbCIZ11dPX7+aE1xlfuFEqaFCaaKB
v5P3iT5cIkdsjxsWmvrLBRbFt7nvlnRo+xgyzSXa1/9PvWI13i3n2735yc8sF2Pi
iQjURRuUrAjrmUL07qqLLiMx4ssIX/EbQlXIuQjK7YjDKq68Y/0aIj3EraX/HymN
K/KyRVG4Q67PxLM7EvQY6XLuwSWpFyHwygcFIGGNuZkhSIKmR8/1Xc98bzfeX+D8
lJwXrxYgsBChgj3SAPxllR2sn1mnSCz7HG+x80pTM2o6W2tDVlzAwY3vAPUtaLRB
eDUx32gRdkU/kZ+rPKq/sUTxfeUG3Pj7OHppxTykxEddfQFb30vIT2lXrlJ/vy2Z
+1pJWaShMwV9r5TvkD+Bjh6VmBnncmRmm+i1vFoJTaZYkQWWUqGNByQvfUBhQC7/
pZaDrA2NaAnWbpxiaxo1Szp2NEPGGnPNB0lsd2VWIO0yyN7fqeELc3zFaXbDAwU5
rX1+8OPv0Ix0xT5tLSdt3edLfSqHctoDStXKXxJZ8nQe7ML/l22iejV5RDYl2Bn7
usLKR3OdFbDFmo3y1vydDusmPbeTs7n85pz6ZcgM4un3eg73MpkiI8WLOSZ/ty0w
3SK4fasj2wffTqheOSgQK6MkCeykaEhMrcWCGT84xSkfvVL2HTs5weZ1Z0ZQF1cD
9tLdes676WJMx/X0D4NoorCdwFuOGef02UP5j/aX7iTHmZVnyiAJfoyPE37ePAhS
pRQ/rH45IQc54E0iRclBhGQAI0yiYU7yP53wdxbDv3D/EHt8pXxQCzM3BKnPIe/k
k/2TjWj8daiSzI0ZAVrEP8ZRQUfyfShCYzDzaOrWdXGVaGZBGo7SF4LkSQ9qck33
Q1Vkz36nuFuXbHNvd2iPZYqaekwIJ0KOrU0g4anc7mM=
`protect END_PROTECTED
