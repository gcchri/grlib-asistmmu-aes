`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/VuxAgjuyrRXigYcvtV1hgY6+W3WnHB1Jn5R1wlpu0OGA0fzei0ZGDewWi0ZpOG
L7AuYup+xe1OJIs5/Ppk7vuA3FPk9KhoAzOuHpR+HtYCwDMjcdOZf2aLo00WPdfp
hX3p+mxsYbYYFfu72B+7s9QYlT9gfxoClPSyLmNgJzVnhuzLmxWdtITDtMhsgnvm
S/tsbcIqgoR4ftiTlLSfeLNVoHP92kEcqClhqNOF24piaOvejzrsiuYvCEscqikd
s2ndvZZl/5GLea7GrEicQCyhtN5ElayYBiQcR+uudJWm0HXX1FEv4RGo4UudlwsM
cTR1yI3TfDiki5ZV31WbEYrUc2ap6MYcBL4JKclSAS1d6zYuRWMQ9Px+jJtPuS2b
meB4AM6a2QOXyl0VSEY6MmaH/EVs3LmKsYglZWH82qXw3UdddnxRRKwJ33A47xL9
AFx951cNTOVfbVp5MN0Jy7oayzvmp7Zy9pnk3F36PgK2aR+8r/Et9ggeLBD7aNQ9
rPPEEhFn7zUECeoOxMNISg==
`protect END_PROTECTED
