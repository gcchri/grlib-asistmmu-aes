`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQBUB3kEFG9yPHz1yKORGZ8QoTXPdXUQ53LyXEfF5rcXDKWWaRQFsVsEseUxLLsC
95mhlmxCwpSxCSGk5v0Jq3FHY59r4RFuO0PMBRxEyPDeLGaQ54DPin+g6Ptdi76d
oRBCxalD04BzOECSRjp121DXodwU6bA/1HGwF4B9nLyKB5A2gJbOAS62bwk8+oVN
oJNUBZ9I/4lJA6RSZV8t6EhPXZu561kxFpN605fKXbzXaPj8UDpDHbP2tDvYcF8g
iH3c2FcrpzgwtmOjH0Xe0h/+DY/JVOLOjfF9sN0g4xJ2zb2tlePjolbi/wQxKKAc
a1mwczI8PsFYJlmQ8+D0LUBH9D/k5uwle1bvJN7QVngaC6tZ8Nhv5TmBZ3ZbLVeL
Rv5ca87Aaw1j3hWofkri2mnCW4BJ5sVt+w7GgH4A9hZcfJDsYWF32TNoEoSSkkGg
MhUVF7GoIZnarZyY59OHVoLjiC/Vlwcd/4tZyPpvo19qxjLyGQXiaMkWJGd/jXt8
vh2eibP5Y1WeIWQeZG/dRnu1nmGXrzqKcd0KymkCHJkiJYIU6gwEdZCiAfhesOB9
2FwyhCN1Vpms/PTOfGe+exjf7g9VjVKB5uW76OA3jtpHGrvFt8nLwINuNClcSJry
yV8YeC3+wWWqgSIMJvBTbrA/KlNFHJrGZpB/MTvmOIUoqiE5YT8yWVT8XsFRLZgj
69ifpOPjg8s4/E4l0synCePYZn+3ew6UxZTfJXXtAft1Q85dMdjbVqj7AcmulCR2
zyRgErGWNQWJgg/5+EL7ESadDarhkogPJBvRiHscbsjYRHT/DY+SleN43QK2cd1e
+yrdYkKiJWEFwtQeGl5IQvZJ9qE1gEPbcXWGUm0CpI+4EF+xgloIXhjIN/gFlc/G
mdwRTnmJ0qOku0JOE4NdMTvZYAiHMsQEu88gwPpjF/qQYxxL+9OqMrljyGVoqFsg
TFJDP2Dwz74dkXcEelSluLvbuuM25BDTFUcVrOhTkGOW7b27T5HrknxrN6N6OjaX
`protect END_PROTECTED
