`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xiwUShED0fu3exhRuPVv676jBpo/MAzLxFblSowxvDC0Gukq1x2H9e29rpigHP9Z
V/q87bmthJs5Q+o5xyW14bOBNp2ftBDFo/ioQEFvQBzWFurwE+wOWrvyjVb1sL0z
ZHs0Gt5TAlzzm/QNMCYnQXK2oKzFYADO4G8QgKprOq+NtHIMSighjcM41PtcCbmS
6QTxHmWrM0LppOva4b//2J2CgsSedRlUwMZpx541xRc3OY5M2/Ir4gUBPY+Kzn++
ASPv1w7LmtFKya6wGVlhTUxfeub6kOOnfKxgpjSGbFoL7X3ELJqYktnKS7QtuudI
K/w0obtHdIlpqlfVRt/PANCDnsqi9oFnUt0UMrYoFavEOkuJ/nLdLUq4hrkpdDRf
Y22+kUykfXBu1KX24Kr9T9MkYJlXE2bkN8KcIVPTCq64lIy+zu5zvCt2sfmLUIy0
JK7Q6vEhevr92gjFyejgZuy5tK7rSeL0BwNPIT7QIH1DnzHTpzJaUbITyIQ/xrTW
Itsf/8j19H1y+xXVhOmVHMaxMOQXuFHx15SDTrLWWsbJsU7+nJ76tjAWRTeBj5aG
94L5+C0oE9UkMij4clCWB8f3Y86F9rlIIm5t1n8Yo6UirAlV8oAs/JoWbjK02CC2
/F+WahT+M2u4ImKYHAWtX4XSonHXrB9Knt56v6omYCPWZ6MVpCwmkPKAVnY9z3Og
Nb5A7nRxebS43U9Fent8n1X+pK5ULI+c5LahHMoNm40SH5VrfBe859gxrU1q+iBK
sYRbClVdHiWG8UwWIlPWTxuy5TmHRdNTUXKrjoHwRhIy9CqiGkuZFiuhOEDvinKI
VNIpYfMBl8HEEEHqmOkC6n8X/z5sl2eCTxn/yUV6GyivFQWepq8nkyqFGbhJ4eZB
w77CYleAhMuS2GlI9+GPbguG/NRkU+j9WhrPMD67pMqJ/cJxCJP/fR6xFns7z1Fh
`protect END_PROTECTED
