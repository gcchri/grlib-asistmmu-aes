`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWLwFCkCJhDfKOoTub5y6IopMorKgs4LP6uerRtb3HXqqFsM2CKH2gulI1vb3342
UhIk0KltufRLieVgg7zBKFpnyGUmeIpBR1Pi+ZR66Wa8ZNc8Cpp6s116ZFTMvXh0
9a3kEolAyo6Fc/7oyEjik+6a6rpA998P6mMG8HAfqywGNd0pyZaE1OPSylsvAuNR
8Plw/upL7eBZMS5Yq/oeVXS6ONL0VD4Z2fmh/WN4sqlUSM4rAEjGpXHKAd9ZoXtr
VCQOaEeNN0oJUtPtgEKSfg==
`protect END_PROTECTED
