`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8NmwJsLhTi4dtEI1NCs2y9N8ZrivyWoK9sGF49f/+250LWHuCKNNbZnP9aQN/0c
QMW67e20129bpq2zqwyIxK3dvmJThqoB2PK49zonmR13wBfakqOFgow676V8YmLi
TyMDMqiA0/OYuClDLa86jt80vz7VihxMByuzGG/51E3h62a8m5MbzTKwuKc62c6m
GbD2ZHJPXgP+5XPv/bLGwPriMNiToTPSBjczmkvRQrd1AP5+cqaT8lZDpFe2TWmW
+UoBENwRxqksnhnGsibUGaj3M64Jg5NgXbSHnrygqwqyRUjCGWu4N/oxk84xCYFk
VcA9lxfoXecBv8aY6r5e6g==
`protect END_PROTECTED
