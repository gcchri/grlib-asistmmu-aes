`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ST/R8xr7rQgqxMrefpkvJaU2zfFlC1bDWTS5GPiNG/zeAV+H65Kbukf8dSmwA3a
013k8GzcoghdQGHpkTSt29FO0eEwrTp+nX4Su6A7SyrXknAnXNsz0OMnJnmCefIe
yKnqE3onHvrGrGOhpq3XhHzA3AuBuNrQDYtSaxSVyKGE9Ju+YSIa75hZT5qf4Opw
oeIquiS+uGmz1mIO/jK7ZvRWjC4MMVochVd6dt5OxFnSVllCUXrimOzBCva9THHH
oXIa5BF7EYslkiYxv8lRyXBm7Ztdmh4dlOwNxMi3HfqsRgUVW0KnxtnFuCy/m8Ox
pn7l8sgzopi0f6KJFF8lGoAPoENvS5XnTI3E7H2O53/5NY/KrXbmKnFlp7vYBhys
CH+3FxWnOTv7HEvv49Jaboxm6EoPXDRdCIEBd/NUZaSTzrZz/wnGbuUXzlDGLT+r
+C89ApMMdyJg6wvWzVurbnVjx7pn+hrmvij3qW+7+ehWGKw/aWnKQqNfXREI1yta
pdnKrwK61ov14C9t0TVvk5ig701xhfU0F0Ggu+6dm5ttQeafhOVhKb/hxyrQOAYh
5ru5OmcP18cvzaCG3VKUzk3C8ym8bIJgHXz7Ce32oVb+FDZycs0c9adEl6zhPIsV
r6aUsAi1ySQiqEMDb5SsS7UbxpfhPeAw0dxTEOZVf9xyCsnmGx5UXBYR/5oTyEQi
2I9MC7HSLlrn3FW0sC5vmT/ipT4fZxcjfsXFGc8yM6yI/t+7/MpEVs8IN/naBm7j
iYUlzN2KJPsp6CJc3e2sI8yeb9ww3R2/I+SgzYVfGN/feyu8+d1Bs8FHDaOv2oko
d01ickwvulH2IfXjhzBdVSNkswCDh21sxzYGgSytsJGOrqs59oSGFB6DlDvc1Xej
x7F++gTk81gCfpuUT/YKQZ9axmp4fC5sg/73v4mz+c4gtZkjswrWERzJ/rpgOaix
X7CNdwed7R0zbG8yy0ZjCv1yzVF2s5r8inNd5a9qgkL3xiEv0YhKqqWhE8ed6Z8O
Kk6ZAZu+SnwA+Ywe+zOIipS8okTIgNR8aWRdjNEreG+XGyjanKOleZ7khKsQlMVS
0O9uE6IqOrZrIe/r1oGD5OmEPBwEzc+3G8VYYcIQtmXyJ9Anixv8+vA2YLVHegFY
5Zu2Mrz1mSiMSi3Yj1LN36EGJY+6s1KuOE+ANSo/P6rIlixn/NuBKEFtziuXhlmN
gN4xsLgic01+5t9h/As7yaJUO/Q6jQbfeNbgt8JsRx1fClVUIHtmbcCG8wcFG1uO
MZg/bSHAcEUcKVeLVvvUN2U/BOdbDz4dh/IscJL22z7EOpLcnyyheXrvL3Dfz3/6
tB7jjkSgx+w5R6VogmVOPg==
`protect END_PROTECTED
