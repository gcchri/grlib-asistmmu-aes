`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vMSvfbfFXsUvVuWoCl/K4rFvpP1pOzbtST2Fphay5F7tXZ8K3s+kR7z3cEKWEKI2
F1RoZlExaxf6LTenZa7ndN+2YeezK4lscu0/t/6YZi3QBt1LnAN3U4kP82toGlYg
emskKdVWVf52UIBumUIUAo/Nx0RCa0n60+/JTyn1Kp6iHbYZ/rzyDsR0a/d20cEm
WuagHyGVyIjw7tFAgiYoWh6wZJRF0s1/MtaIFQcjK8FAjR/LB1CwTMwnGXSJveQT
wA9vTC20sIYiedLjYRycztOrGYdE+2tYXJYqjCnWVsTMaBAkk6MKoxV9BLgbnrxm
8Hs6EAvE3aYMxN5Stj4tb+QoF46Ywm07Ss0LfJgy4Er1O3bWrHMhV9AMJnmPzJ2J
Xx6rucOnGl+FS9XmzwuY2FtoWKlYArVx4Cfl0P6kpqHuAu6THJ4QXj3HQXhO4QRI
grch8vlovya31y2o9PkhC1Huy0MQoWuJFq0rOWRTrv28N/qTV8gcOTpY2EU+Gmw7
CQrvjJIn2ORWwdgJoePjdj4sYy/WdyiWsCmIhgDg+Hw=
`protect END_PROTECTED
