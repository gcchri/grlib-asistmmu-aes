`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5TthtB3hUeLGaZzFXtxqptmCH4SEfC/xro8OX1MW1dVAL3DWYvDzofvSEIMayk5
RhtpT9P9a1TqZKpJcYs7Rq/Odbc7YmkXgTWMBgQfrcEKjCU14AZfEYt2FTxGZuth
J6Obr+eBuovoyvgtxG0l0qHnFN3vcUwK7OYODkKM++Ki0AM7T3m+q5X5JouokLbT
2c32Bs6v9JCRhucPtpdJqzpl7vsEoZjkif203i3SdwDTAlzW1WXfgBTy/tBc8rjv
`protect END_PROTECTED
