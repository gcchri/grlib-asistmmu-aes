`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vl3YmsjJPq8i9/WpVlyA2C1q5AQweBfTrBC9BJLXEsPBoU1mlnfNb4z9egbc7DaC
T2z+pa/5Fy9WwdP19DgKIb9t7jLU7jdLwjR/DDUzZFGlG+dhd0WRMbsAFDXILAI0
UssMgErc89GYnFiE9APhky82DPAj/kgShKLpx6/89p7koAO0uYZtLVnymsr+t93a
G3B/Dczw+PK5CB9GBQ4GN3/VLNXhOuH+9wGyzccPQMoppIZ7X5XgeQ5wv4Dw3R9y
V0J35hu/hYNlP9bxguRjbk2zOC1KGUfMMvdBXSU6wWi+j+AzCGWav25oAnoYaHfh
wZe74fNhkjCElTXlfH2n9cHI1Rq6bpFjAMff6QC/BIhlU5vbq3fRZjXLC23XhYit
nXcckBUrcoxySFo3Iug8rtfjmpAQMZy7n1IJrSk1+6iZPa0iU4t/n9sp8342C/CI
C3/vE1Dc8tkPHPHF3MSumD/RU1zQ6WDDtm3wu/FwDJ0lW82kahglAmLYj5i2de5x
4CER3slzeWm107WBSr49/328P7mpZBGHRCxFMHwKxLU=
`protect END_PROTECTED
