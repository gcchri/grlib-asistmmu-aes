`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4uEyaPT1k7neJO7HgAZ7RpIr5dIGVd/1LLlt2fsooXg8Y/IAJHz7PAz95uZJX3K
gf0X3L6SObmzv78tBsR5emxh3hC34+qfrOz8yibIN51/0eYM+JsimwW4vMkWfa7f
Vp21feBdlUaQU07xUqC2Oi7jtkwT8IsZs+S1NryQNnsAztbIXHqvNX0ljgSuFe7E
8UzRMIB8qISeou4wjXuYRVMy4CFhaQpDgAsG0MAxjoG6aw/XNzwrzEuwJCkh9Kvw
iEHUwrkfLtIjY8DvkOiu5q91gQWw7E6xBCTgvLX52nc=
`protect END_PROTECTED
