`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gxa6Dc8NNJ2YoCVGtVPRneBuwY+pM0ScgCtzhptXPoxMs65zl5H2Ui3RUVEJ6fdt
7LxaM94c31AQ+WYcwaohdkHJIJT2AqqWwWn40Kjc6KSj2mc1Nl5hHE5IS/HPxkfR
VtE2lwe9nNAWNbRseeDCBOAkzyEOEdXEDO25tbLA6UPG0fYVovVc2dUOfLbPQeED
KTpEl7gnlwGbcN9crdRO08HZHmKIYRpgmShpVaKTHcRR817sSKhNS/ryW8lrar39
iN7l3yWfwZ4yFn9ijBvoyvjtGsLUbP7HiVV2HdARdBgACe+79r9Uv2o6MIxzVKyO
C5xfJTOVOjHRfDFNyKdS/fDKdyksJLaAiJoUp3we+QFZhrLRXjpT66rcNggjvKnb
KgpT8lV6KM75a0+oFKLLOkAltwmf9hFQr8wrBsB8E/qGR38DNdXFwTvb8+pyoo0g
BjExngK43n1z6OmH8OJL3OX0mladgSRJ4h9o6njPVhw=
`protect END_PROTECTED
