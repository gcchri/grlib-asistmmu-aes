`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSIjJ0/Nwsqng27to5JPRCM6Oy2cj7yWvDNxbkM86J+q0Mam9ax/Hl1r2oJeo/de
l/GHawIuER1B1VQ0425Fi28TctCkwG0XHoyqULAUS6hsEhTrpJoWd/lqIUo1fVHp
uhKkKxeMpoFfPBxQCmp14ji5O+FQmW8XqoxQLSHfjL9/DY2CZXaZkBvJxHtNZXvI
fo1rmvLz42OW3oqCIwNn/YqRscpNOQ5gQChnwC63CQn4pd1NAeGPrrrwbxTRE9LV
/OubmpupV7GIJTzz9z2u8Q5zXtOWkS/WWoquq+QhQS8=
`protect END_PROTECTED
