`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+nV2JZdc89L73JRU4JJNuzzFVpC6WiLJq6t8glLwaO/bc64JD0HZ3Oy945z6Ew7
H3zjPD0lUIQ1QIc5owirAA0BqPNu5Lf1iOwfJyFX0AxZTQwjuGoyo/RpEOksQjg3
RopuXTUWiLDmzmD51sIa/ywGRv7x34XoH2XlKUaFbRrv5gS/+DBfr4h/0ScZpndn
xS9X7hox5i/RfebX/H92/InMEKy9VJz9tpieZrSLJ16GKgqujAod6aL+PmX/ppYz
IwghZK0fcCBfH2Ov5e+IQ6NZtnBbzWhcOhe2LOe9wrhLaeUyAmdiTjm+DcKOnjNa
7bAhATgNh0c+pb7406xonOQ0FDh0EhVLAOzc1VyREfrEMgEF8wme3X+HvTzVjZmR
SF9inTgKt74lnYNRG7eHKte5sHbSawASDwxblLkCEZmDf7jIvDQCDgn0Emr1WQP+
yCkinMZ9IhADJdDfjXGQPYjPBZU+soFVBsyc4cnG7e30r0NB2CvR4cok6e+qLWqy
03CwX2QjCiKco2nqrat8fa4hggJSi+aEa5jEbRD1Cf5j2Nz6CI+tGdf/qsWgItyz
RdvQmyM2KkoUZsK3lVDOirZfj2Glw+VgLIq9aEeroC6TSQUHvvvD76hJ9TI4qP5I
ZLE2wcMP8Wqt64u1+PgCX/mtPE5u3RH0NwnW4guaIYeoe0DSdHewyCNz0R2V/uBk
IWQGfOKGrvm/eqY/evfcnjdcaIvmg/ZHyW07L2Ltt/GTvKIJZRZAaQR/nXg9Nrlj
4tDbD8w/By8uSvSElTfc9dFMKdE/UJLETtVQAflyuA4QXPd/RIbBPk3b2iwevMk9
L3WbtjArryzTs8lfoLI60JmSOCAubUnQG+JxBh/r3psKHNZruHpZDgSQXvlhH/w/
YyA2WXXH6mE7u07e4ZLie3d69setZCImcWAnzhPnjUABLrSqLm90uAb0iUJ+gA8z
FoPlh0h1duj9looyVEDSmKbYBTXr6AgJ8ydgHpoO8KbmHd3SHgnTYBLSGd+HiXjj
GEDU3+VHiPQKQbmRuY0P8mPqRfgnLkXKj54zyLa2EPRqgSY9ISxcdmPSzcLbc3t0
c9KJ+J2QxraG8YHYsMSugajqB3f6ydeF0yddNZFJ6LCEOexKXT0QGYb2QGkD/RHo
0dEzbdVj2NHWjT50zJYGmId4cksSthGIMh0j27o6jYQDHpuAXhDmGj5gWwiAZoN6
ojCxd0gEf49OjUZhfJpBbgFY9mjwcKJqEiG+d0EYydGP4UU+pF4qGRi3hrMFcaG7
+HyqYgSPrxDwfmBBYBAg14agYFvqRf/6Oa7E/NNDeWEi3QNIAlmOiIM+wkslDwrr
Tv5CidvDCYzGlfbT4HFsLfz5R13Hot11VKJ2FP6FedsU0jLO2x+tGNRZSGASfRhw
dx6t6kEZhii/p5P8WiWwqkNxQWnZpXDZSe3fJW47O5KqSgTuhcY/UFocATt8kVur
qCA7P3jy3DB6/VQBO6ms3LQqdX3bGoo7fcIQ7vjoCqGhDedpxgJ7xDCe88bwTQpY
7LYyMqL3IJGSODB1ZjszNEsjvB9BTDwaJx+M+co0KJoEiAB4nAny8RLYSn4YsYdW
`protect END_PROTECTED
