`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B38Tw3BHMYyxkeZC8zgNHz1jdoy0DTRDbuTMmtlRdeWSLcS9nClNZUXJOOKTZo0q
biShiPusuEax0GlfjFyoQzL6MQaGCW21dkp7cBK+6dVi4e9fxnuPdEMi6LvLnJYN
p/zccbjdk9uJ9DtD+HWdhSj/LHEHnmnTlK88TBS+GXGiegPjCnHuwMOEAauXOVxc
lYPK7vc9yAb+ic76lWPYsurG4IZ8FK/f1KElaoO6YscL6EVsowWM3Kic2MOvc5eU
OEUmHTzJWNaclJkHdyS6/g==
`protect END_PROTECTED
