`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwKNFm5TOiou0Llrzcj4Bk249xybmRcpEq95PrSZAzyRK9J5NX2PnMzYu+136VNn
fk+X5hJyQgIvb50ApPMCvsOgPsEbS5Rule5LhGBl84Hb1qB+/iv0wI6qon6J5hhu
FyqUTvAYiDoqViy+YN4d5BMpd98h+39orZvsk/Pdrafpm2PJtM3uYelO7AwPcpig
+NjaAAXXHpSk0fGchjWDqEj+zARkEGiKptTU9rtJIl1sCs2uHTPn4sSPQ+EVmown
FCmz9qzCs6HLBX2boldeUrmjnLU8v15KYBfBvZO93EtlWeTo81rDBlivvI8rwZQw
oTslGkzWwJZpGu3jmFQyZORJib7ZxC84S3GIaQCcyizD64B0ZMNOKAqW55A+ozyA
tJNy+VusIMsu1JTIOhg7WicGEpbL0ONQAEj1tpg1zA+JWNSQVq8kI13xNa1LmL90
VkH3MJIc41yqss8pjzQRJW5sNeRIglzP9IloSrEIP6aL+gfWxtbuAmJ/HjrIemIp
IGDQ8vXQIgg/OconOGHYpQlIrdcXdLGu1z0ScDaU3Ix4Qn0pW3ttaUAEzHMbwKcg
WNJFUH32ulEHIikivLAqNZ21+iQE/y7q+WYKme5QBCVJyBkHilGR31AVGLegJCqg
gbrTkZOqdiSZTi5vvJCaSZI2H9taAJeMLBpgemhp/hOOJSw/0PEc7E9lC/e3Z6V/
nWoJBZHdhtV5GsTraOYGhUdy9DNvOvhGxfG7GIMiGA8LJ42CDswu36vhXV6rTfoo
wNrmh5icWj6ML8O/rwvClgtUKgxv7rTKHLIGLBNpAq+Am9iXTYNScC4c+yFWiq+B
oScEoGCZgtXC2+1e2tnhh+PsVF6suOMHOzggmQQI+aCfQCvhu+1DOuLKzKWWCJni
0U2JiTxM/UKueStnK/yTJNMCrWhgkr719Lbp/oBx4aHdKIQUrHMgwIIml4x+DC1i
zQev3K+rQT4bGcl1S9pMdapekAOq8EtGtwlnOCNZs7cuKkfC0Spr7x7n44FmO3Hd
qJrA8FrvH7mo+Lal0cZXgMSK3i0Rfn8FosrYbQKvfzL/rymF1Qlaui2wMxRCswMU
o7YUDDwtzakCL9z8Ht81u/6i8n/5x/XPLq2OUw5SBRpJqHuToH+oAGw50xGy1jfm
03urLNb4KjSjJkzyzm/8oas63+/Q+pZTxWu/Dre5zoIBoRYtlW9JxBrjF11UCfq/
/Mm8HlPN29MczCM1ENbJx1stlLv7ycDWNEPTN8wzbM4=
`protect END_PROTECTED
