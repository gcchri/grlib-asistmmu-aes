`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WIpgUByRJTArm9HHgAzweeDlz49K+ChZWCA6AC99RQJdxuz6vj8ZmWYAeJ82zzwM
e703/CvBl5ZEmRBYxwNBg85sNtB2oqv95Owkp8IRahCUSbo79teAa7450idJFJFi
KQzXO4TQVsDjQIdNTXTFbfPUs6P4KSF1qRroXbWx7WQFWfO8x0jCId2tg8dutB9r
I/DIonm1sFMnZEaQ2OHus6uDAoFNSM5C02c02V/nIB2enp2dRRJDJtsyQoof2qLd
Hqb6KOhLa9/7d7y/78BWvXjxEbzCD5kEwlYn3djBJZq3eZKrQz2gHAxqyCeBcCCT
QeL/G/IYW8itdLtb/2Si1RBOPjURJGnoruCnQSUuFfiuZxgEoPAZlWQBhcMDixV4
dIqYpjQJIuhJKG+PbUU5+gh9P/1Ks+j160nmgPJzywWBBOzH8+26LO7kPkX6f52Q
6D8gBKJHaGuj3Maoz2jvUifWcAmZyPW7P30519gWwmHSFp+8AO7CBG/WY2czAWue
PiTFnPiEGwDOJlHw5fiPbdvqlrcDiRw/y5htzc/5t5rVwO1LtNSuYplWPknbfpgQ
czR3ZyTMOp2dWs6Ox5sVYw==
`protect END_PROTECTED
