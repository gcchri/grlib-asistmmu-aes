`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GToh3wfp9R437tXNaG79ooA3wu2LSSfTxmMyfEidCwz08M751vkbXpHTINpg5/bu
KyBxYL0Ny0Q+AgXyqWT/galpC1lBlEyQe44F1A4s9bsu+21ll/Tpw5IddEQBJiHl
7CrvjM+Qw7BuFpG1qL+RvMT6InyjCOHPyGEnhtF4vZb788dvNKSdeLBAzxr4Cw2O
lqb00Q4J9QdKvF998S43hrF2ZNHgMFFBbX74+nKNHC1SbgQQwwIyqJar2qAzTt/u
XWbB6RoERENq0nqXxuPo55WOH3qq4mjD3ooif+dWE3iHh2Lj1AjUBWaWoy4SFNWJ
nfVsamKpjqP+NMLMpxWdfM6JAjGumTFFObEShxalOeP1H/ls30Mx84Cnh90xF5am
3+7YOWqQFw2cB3TIVfPd8cZ+WDBr1DfYpv+yPzsQH9Y6l4JA4OX454J+2geiR5cU
AzboaHsqcpFqdP+ozDJU9+PbSH8Cir0X9qOT8tQ9/4L/ZVJAd0PKIAjMn2nBgIfh
Mgft/RWgrlyVR/rAMTgJGGFv7UxQ2rMpNXIM8CoJQko3gbS4jd0jegtinwsYLqF0
/B2dkafCkQBejvJzaeezR/3IpZAzATORDKGs0/eK7SLGnJEumKeDTZI7xhkmsrgy
nnWPo65k7vZwI7sKtJrO6hFQ6sg5Y+koy18ejSw4icEXltpUFkkPy17Ikpqjej4m
RbZu/H94QdjjABGarAj2kaH+7cJMRHfFtbDY2owdpUTxFbCa4DSwEkZZHozZ0EgW
69+8hDlzktc6Td1vrpMp2XLUQVwOrWnLcB30HisdzHIrCQdQ8tzIvBY0QxysEA/c
1euGofcFZPTDQ0wadiJRiJbFhjJAi66jql2oFFauysILGCba7mn8nR4efv5hPgB4
MPaE8RXhc1yZRyMEFz0ITvzDo1RwwB8Lz2yODWL6CR9BZBA2s6srppDO2FG/CjXd
OR58DBEpVDVXGwCkQtcWEuXH+Ye2hDuYewAZ/RosQFKguzBKoyRqm1liBjFsF4bO
tgDA3xq6yUpmhklApO4g2dOMw0PQeo5cE7FqCQpnq5XBvSNe5o4kSSZOGVUbp0vo
pSB1AvpaGDxNAY5FbH0afoTvfViEAKDg/G1EwQNVCInx367i+aoA4GCa0ZFfmhgB
Etn2k9upWrTFAdZX3SbMmxx+JJbk/RyPIGHrnyJTX5D9EwC1pifo6+jcZ4uTnSzI
bedR9dL8dkHqw2P+VYusy2jtTxjXtPbOKfahDeD8sQiy2PN+FS3accXS7/PEh//J
HV6fd+CPLEQm0OgyXYTF+/WuHJA8ukJLrOVcHmgVr0doaOlAvH/YoLtq0AIjTMMG
qNIwCH6sI7qfmeQF3fkdbWJlJYtWgHnChGUtdJ7FN7fMK77xqQcwIwIlzhjQGbjt
OshzhTZDZ59jyqBxpgJTddffH99lMZwvZ5vB31w7j71HPHOSBce1Ma/f0JeDBPUd
X5PfxpEq2cmrNfVHetidlx3Re+a/CZWihXLszSYA1kgQpripRBj8mmNynLAVIIm+
9jU6PPvUy6qzJSnIRdWwIIHhMrt/HvPWs7YiXnH7XewAOZ8Lhn0KZWU5QnusJJ99
oVs1+DN8wifLUNI58zyWc3nNj8DnPTTOPT2K7EqkQAyTe+dP9iyQIwRSgYek5bg1
x1KH9RK9cqh0yK1D4XF6w4wNBx1/bhHWJ27+msgNo/rgygxGHE0RMjLRNqYKmeCM
OvVmvyqyX3IO4kpHJ5VXyB7FENJFfkCHYM+0gDl+eP5EqNfGSPYpA1I5o+UWafom
gqELDSV2L1RrTPENRDlhr280HY2LYZjei25F8KozpNrv+dfHVKElAumAzToViGDz
S4vkcf/3zkU8umk6NIzv6Mos8scYFHo5Nb/mEmWH2ClwekY+bihpb/YQTdv6d9zj
es/YyuxHMZlJpkOoJq6gjO8LuBUvCsEl1ZGWFDjU4k68xfNJb8mXumHu6ksYZ5Fl
DbFVLG9lXaz7opUcMmZHNfpkxQh9gChshov6cnZSVJw2lw8A06FZOoOFB5VAptnP
XOsmTegbR4YHTFdZAInxL5dlHEpXRnIa7zrdamqqyHeQFAiT1YEd696vSKiXCQpr
6i9Muwj7WJn2x7iSXJCvfNA4b/gh1K192YkFQDCJH/cvTnGTRTULn1zk7mK+9rx2
XQDs69KPS6RueADjcvMeTLYM4c0XBlzpWT5bey5bmdmTiHhckFgS3kyMY+8/w0sE
9nTbFxsHHvteBR7CR2nnhE6UddZGcq1IWzPE90uvyGWhiVi96xZFpGbdTUA8u6hd
gagRWcL7LAAZRwRc4vS7Y81lm+qB6a76pDmBYvYOPeau6gu2194mL5FJBHJUUAzU
r307nf1r91mLs15Z88nAWYQYbUFh0fdoxgGsM96sGWO3xXHoHjLjggX5aU/9HGZH
HXe1Uolmyy3KtauzDlIE4MjWZIVXMswRSYaNQD8fNHu6kpGtBTfAppuPRMS075q5
kYJAu6gVpu5pmsLfnOQfKFSXBrclv4E2w2UmAfxameaBy0NGzqsmtiawt0TuuyGA
IbCFBxRFc1sKf3ZP40WEMQd/M/74W3xbMHrVniBVZKdDCKm4oiOiD9x0lT9otnaZ
EjdII3JstxubtGx9lzzS6hJD2dBg/8VrLiBc6lbGUzdjicvGPXMm0IRzIdPhy4LB
5ZzE4VGkzUAs4413lh7li2Xu7PI+jcT1kGFVlOD5gJ/WogtYFadoYQVHk+OOYNJZ
UXyLl0kel+VYb0oB4k2NlpfWMo1eN5FFYaI+gJTD0yE8XtZWNt21yKvNlU8o0W2J
fAN30TbXsuYc/1hycEieLx29BUk5oLL5lUaJeqTssRw=
`protect END_PROTECTED
