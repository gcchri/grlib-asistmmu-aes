`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QrXMNCU5hn4aj+KqzA3M4iRhKKqraq1V/b4htIXbHKr/fkLh02V0Y0dxayEEgrTF
GD8ZHEpUuEYgzxbdIZu9eCG5Tf3De3K/MpapNfxuxFe6TTBHhGKKwN41sXKNDrja
R2DGqaEGcZr8qFw282/IR6hySG3V9dR6GCyGTnWlnHCjYbuZ3kppN63rXjK1AOe3
X9GZdGY4YwMLXRxawHHGJhjVSa3Msqv4uBnbj2ZzYMtPOOJ9KpJQJNyMAfCh2ojT
UpyISs3L2+JXJSxpbJri51Ks0jrmzG9IA0a/05osWH0ig8QujYxClCiUsQszTv1+
qMuQjj2wVnrOErZQrEkNsIzkRWfALqvvKZ71Rsj49dk356PfV0MoJVgjKC60o3ac
AtuOX4Xt1GvmQGmanDIb4PJcVLqHYylFGp9An6/NYEt908+0WS4cqckNisFNrxMl
Ks67wqKigg6hgLXm1I2a1TAf0uUh2NIFcGhvkk9d/EOTKUR4L6YyRDRh70oGCUH9
Gg6NP+TqTBmZPYztmneGJoVZMVqanZt/YzrhJ2vccfV8TgkjE1OIfDzMcE1NNxOY
xQfY2xkKMcHN3qFYIIbzTGYtBcfRCibbHWMRpobT6rM3Wr8wuI+1SB2r3aiMObeZ
jvFK08qL3vqmWTmwiUNaN7x6JcPayPHVDD4LoT/IkbYzAo1DKGVeHlbPnO+AaxVQ
kUL6tj4k1+zPe/hDLzB6Q7CXU1qnO79S4djVOEY8BFfuCi6w2RsbqLn0udKFrKrB
rTrslhvLDEBfNuVNI+DmlN5bsVlFHUcKr9Muiz10OvRHQZ5eXPgrN6mYDpSAznET
Xz3qD1D/rmb9emE+0pkIXmvGiPwkXONNV3VsokQ7AKq9gzCJcpSBJcHgHd+1kvbS
CxG8Gx15smgfy4RXQk0bi4lr6fLtpqkso3u9X6gC/ELfFloiXnBCPvFpw7OXl4RQ
fOuYqu97aIfMlfRBk2kSeqSK/+qLg9875jVFZL+cLR0sulo+q0aBmSLnfYZ/Su3V
ftetP11DGNci5S7bh5OlEhgJsop3SZ4zqfDRX73TNcNOTYdvD4JQJ2wMTR9UidW1
9ntO9MS4u8vJ+ABxJEYAtrhwjrBDSDvsjTWFFVrl8Pw3OpSLzXgA7LaoT6Swte7o
b+1tDkCKz5Y2UsFdYZucKBAgtFqv1IWN++iaaaiQ0X74oEoHGxzCZt/3i9MUINR7
L+2RM0FTIQylkiDkVuVoE8foAdhZIUPbm34ii8KfGmgmeaIhaoZFyZzKe9i8Q+67
413N2ag3wNxufFGqA4+5nCLuGt08XaJ0ZR0hBRJHfx2A4af0IHqz2YDjkltOqplK
KUgEkN58MsWjIEy07ILZuW+DjyPqKs4QNQWrU+55a867MJTZqrf6xBvWgrF96I+c
pYMQ1N8Dybw//1EJQ0wJTlIHu2hqzDBz3wVUijA7CiiuVnh+0z9DlkHt7QOn9XaK
2GDLJPwB6cBlKgkSo2HFDYIfBaUoDE97RTWqCKu3+Q2cXrnZLZsLacYdeyI31wVD
9NGwLmOwn0FlhUUBBLWNdWaLfWxrGldmnY4ensqnmObBeqHDRNKlSBbhqrnaGoLZ
qRAYZVVeGQhTXqC3Ml+Xcr+IdqbTHoytZnU0V/qhWt5npjFqd7KQ2TrBTp6nxCfe
RqyW4log19WO9uJkURKvOa0Smp/1kb88bjZ8MnJhpOm6Qpwm10AwJ89IkhIr6SJl
I+mCV8X1Lo7YWx696Hu6u7es4GzUPnkGsErkDIxZGNRf63BH8NNno21CIypyX4Tw
1foOqualizbHU+HcGqUH6Jg9SlL2cyT1pS7M9Hsjik/4po0oo2t2UixLk9V2NLcL
vV2+tYoqJDq2+Q5RRrfQ+Cgerk3ToFBEu8LBe1oTEeU=
`protect END_PROTECTED
