`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lc+g9pPPCUc9zpyvRvw2SXKBpOto9sAjw1o9RpVvFEWWiInbD7ygz7uAU608xMEJ
07Sw+nSYBR1brKhcG7qZwf3Gzs65Zvzw+Rv0H7UEL9dEMkZnTwUg3JoIkvwf/P9i
oXWl9Umq7mb3SPQfJEj6/jxFwxkgtYtSqy+Ebgg6nMJ5WNXgAegsWoGbt1Vv9laj
UDolvKyf4bOKTRrdgN3KQ+ON6aodsbQMmDRRdtx7F9N20GXF2/MYwDRH08N+/Nk2
1dTl5Exe3Oyz3VzYKUSflp7FzNsVgG23juuvDWcgPxKDP3T97zO7uj6Syvz2SFtA
aFbLKsxhnCv7r7AmmuAiy0qVUupbvx6Grt8aoXROCLoQOpU9VLHIXA/knwFpf/Ge
TrxRGahfpT5nuoEPqD4GneRO4IGgqTT6qSHBTIeih2yDf+aFXhKl10oZuPk5lakB
TWevoHjdxFJ9iO3a7fEgWjds+AaPMF8xISAF3FQP+6gaOi7vGDu3MGwottZYlq/P
lOVv21xpRLVWMNpyzfNSxa+52nTKi8lC6nxkaW0Y0PgFpZkkjawUjBzRuq5hm4EM
cuJENQsGYbDY4UV9iRwMq3wGO3ZdJUWFzeyzQd5FRC/HeEeTO7BwBxU5jv3Qwl2S
Pj0QgmEPQqHCjf7hqNuDDXnLk6hqojqFKNmNgeshyoxzXIyz1shUw/y7zct3yHJg
DyrnqLmFOKRa6Werf9gCd86Ikui8IryNsujFXi5Nnp+CbxPoN8qxn4xbN44E3txO
jtWcp15Ncn/kYON0ALCz45Foms0IkTp05GcW5sw9R0/YCJ5zYpWJOfl5PQMlf43e
xGmpU32533KweO/DLQd7okGnfeLo1XeYlbSMIQ0dkjgwWImXVVxvIsshB16jWC5j
/PVHONxEWcQ8MAisUa6QDbY7IdXG6OrbV7imqSs091npCeVJnpIlSY1nC/OMy0RY
OKXxYXjqd6TmoKQTG1QA7WJtO9MmoBNL8L2fmlhwKoJ/Eyp1ZK1PeFDSLdPg2Hu+
aDQv8mXyRwx9MGgoO1pDnZ2rLZt11JO+VRDBWbt+UjbZa/j8nTxRsJT4F9BgkkZ8
EOy6qp8NpuS+3BM1FTF9R1KnQ2SccOV33eoyxrThSRMr04gLH91ezETX5PEL9aTw
gwm+yEy0Lt50BOZ8UMTYH4CONWZmuqy521Ag9sXin9Csw17BzbZTgC4TkFHkMUHf
/+0Zx26TfNYJ+JDBWgPXfwzfGKtUcWpZMh7VQDMkO7JLe96Q6Xitv2M8erRGZ13g
N1MaZInbg/q5H+LFCjaDNkqapBRv5B+y819lvhHtpuVppgPWYMyb+f9eEYmQBEvZ
2+KBtSwoiBKLjZXO2DGz5xlPJz1iHc0QcY/SE3pWgRuN9vQJRvH/c89tcN8xB7PG
+02ulCPkRjfihN1vOfnksqRdJ6hUK4eJ4FQ5NgHMgN9Euahovi4HXO+nNDzEHOlV
BKxEUrOesHpAWBgDAdQXkMQJ1jyAmyr7e09KztemjgH48K2gKY5WD/G0I6kjflou
`protect END_PROTECTED
