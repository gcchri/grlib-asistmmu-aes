`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OfuMdivNnOb0P7LyBx8nhMOct37nihJJwkd19RdlRbljHiTSJZh3TxZE/kfuzhM7
CCDDKDns0ZlvGZSFZ/0bPtpRLMWBJlWDau/lp9jEisGdNUm53KHjjki1bmKzNUPl
MxbzYmz6/Nsj+ibcTrXjs0cl1YWy2y6A2rI9BoI6+JEtmiXUArjmOdNq8HQLGgtg
52laBjf0iJlZq0/DcfogHk/i0igMxXcUlE3cb3eV8wpnL3nzrvFOucyHrWjqZd4/
XEdmLQzqNwf1zEvgbPYWohPAy4irYouzPndYB31zZW+Mdk33WCKHXcafkjrzrgs5
DF9vOACOLR53bKdP3UqHCp5XRvuC9h4fkyaS21AR/Gai1Oq4eEHXEW5uJsPIXN4S
7SqGEhbFeX0FBfbywln4Tg6taPBOqkPCDY2anDiGsa0fRaMr8R5bY1WsZ0icq3A+
`protect END_PROTECTED
