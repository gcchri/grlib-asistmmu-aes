`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZkNRimU83ThrY/bTWBijGoKH2Etp9/v0kA1BHuXxgo7X+AF5P1iIhlRCteiZThBZ
NsosToVLvO+qQ9g9XA2HxRQNEA58ptYKySN4YQQov6NGTsJ1hH3kMjfsSBHM36h0
YazKRzn0b59CmOuM0k82PL7QO4r6GGeYqUGXjgCq3j4RmVH0njAVW1f3aJJEkEVC
CzKEqPAneuia5/6CSSOdaGKqkPpDojELyeMjoXcYEd55iJLdV8zgHyB6PycKZEnM
EPYE482tYxKnRAfeLYPIi2CBo7zhycxgrYsFr688BkzaeSLLrGfLkfXQcd7OybDn
Bf1nlHtKRTyGYtsjgG1cv4z8WZm0bhNqGlRHLclLUOoYLm+Bro7TVFrnjAOaTzPk
L9KiACTe2y7GW1TBYpnxpU0NySUj0agRRj1PdZ3EoNDf8qruADJhRbVYaK3STen7
sucUCTg0EqcSrVMZEf2YsIXzlf5qZ83+uQCVEFVzFPkh/VBzLyRtfOZSmT3G3dE6
Q5jxpQny0i5SjoDLtlOdq9WG3qdPZQVgShXU6mXM4WjrL9mDJJIPD04CmVYkab32
BeXMyDS4DybbyQWnHy28c83E5Ii4+9Ytkn0rJVGATkaZeFBNQdn2BdPOmivmq30V
u4vFZAS+fPDmYpnUELd8UBTTyr/M7zD0L/CCxHvr51ZYT73bvdzg0umOozLG/MfH
DiNGOyZ0RduFLqBh4p9m2j4ZsrbEehhGJGs/BQ45nuNt7P1xqg8tVPN85+GVKgwH
bU8hONtlGfjjgoM3V5gIz2NIYHkghZlQOo2nCvJwIUFh9ymrTUaq0s3EAekos76p
kmH76iTDvuQo520QXG/lAln0+fWbjSt1Mgfj6VYdX9OTqdSYehGR2DxIm588FtCQ
+CFfy9T6jnVfJA15je3AUT5/R0rUPIOE/adv8a7OE/J/qCJL6jubIttkcL0UZM3J
zp4fJnleuNWZVwEKA/9TTXxPTNCtSAy9WlpdwCxHBffhjmIcf1lukkrflwoDs5pX
sOxjb1motjS3u5hwgD1IbyGZqBieDu8I6XzfahsrCZdzVIuRAgUE0/oUYnq/XTye
urt0bcA8BDLpb1usznbxdm3O/Jy0uJ4TRrmr5vMpwzL9P+FnOjTWAafRjm7hp1iV
ukLjibIPo9ydBQA+6iJmcflrWrHKpSP8n8vXs3PsjdaVXoXt/hg54Wo4f/1iRpOo
okD+Tw9sOoBoDP1Ivt2gxLd7jJlsLfBlMQkGhlWVEZnPy9N+bu+4jyA26VJW8L5W
QCjmsqJXx27qP44h65faieMPixWTiTypTjJlsFqK8TEwAKt79gk45mpGrPeBUXwz
fKjMfHy8yYRJN3QiRn/sRwNefA9w8xWGslpAlukCm6UlLdGbAKaZmSU+uyUSXnYN
qH8WtCxZGMiBWd9Stp034ZVWLUgNh6178xn20Dg+jxbv4HG1XzardLwR3EKek0Gs
fi7B0BZkK8bF4EMRGeAOg8sMuxTcyc7CaSIi8MwD5ovCreYyS9Faz4bcx1tcbNt2
2eze9vrgIMydGg+AGGqRIFOgnBn9hfmbmGlvNaV3xkCV+DGksUp9rcbJong3aD1q
ohEP8IzDb4pSbAti5Q8LzA8IRo47U6WbYaXy4DyWUMYUKHQmsd93Qwy4gpXgCVeT
Zs6LMWWZH0BIvVuIDVdYGORVPVkTL5bzacLiiCOJmkgTuQOqkSRs0+WmseghX+nY
9z+MRPE2uWEVWYiWxlNHFkafbbcq0J/k0uK0dwVxDde3zvd23uWKs7YZXzKT1hRx
ktwrAd0OuPfyaH1wEuokJ783ezZRX3eYfgXNLGpEfPGHXp6zagNFpyGKlrn7M0D7
dnzvAg0eAH1M9qLH8GdNazcvtdpl3O2NAqgwTr/krtxc7khI/coZ7t1YmCql3h4i
P8uTpH/IpQ00Y1VLXtKqCRpzRiqNHd1PjUEsuVjGiz7etmPFPFvdwSc0DP0Zp0po
3zcjWKpSyeYUw0ubo3gCwt0OGEva1tIT/2G9Kc5/kSfZy7zBVDfp91xGGsylj3x1
uBhCF7Z+fiRPvzFUu1//90anQ5Os42WuaA4ECUSVUD7uTgahKFMRfzof2FTwvR2E
WGua38zqATNmtSzHlqJbfSMOZBzBFi852bOa+1lXg4MKHModSwnswzDb8lR4Jb/O
7XfsvuBWkfa1SD/4C1dMadjQwevSLIIBy3LBnd1gAS+EK06NxrhiAdnVusQDnL+i
4bskjd97DfpNIYuNxtZsZ+0RWn1BNshJk3fMdps0LbI0lw7LvclIweTJzK2Hc3h0
dzxkr+xSRK8cOAWFEWOJ27M9D2zRwGq8ufApu5M+LdRP1IZDLDk20FNxtl3g5p2Q
TWlKDDkiEq3pSetht5L4UXE6ddfQpi/ckXmIARv+2ISXcUcTPJVtgGKxhsYOxgb2
gPxokZ2x5ZGsUHbxxpQPUKqel73CLHHpjiBP0xUEIUhPvoDM7nOi//tVIHiPGVjm
KQoc16b8eCqN5Js+/BuK6AqWqm9GbYyaZ3oknvOrk/7wDD1TKs8jXAw+TOPoY9sP
y7lEH5xbBKuxKP1yM3CrftOWRUcAVkgP+19G7bgmYFPnTMIrarM8hWvCyfi2+QA3
FVCzUZTc6RMXfhLqnoeJCjQbdpaBY5l39EAEPxnwu7XFZSxVOF8ob8Nwt4hQ5l7Y
ajiZnfirr/IlAR2GKeRYT5++eueew6GgNBn5cjzK0t9ulm3zFWW+tqNepVhHqesf
2m7OeHe+9AHgXex9+ndhn3NYglFSqXBy6uj3WMKMnpdijA+JaqCfIIphyQEQ4tPs
nuAFRcngR/iqC9vIqv18jbMDahjNMjVSj+SmzEG7QKodHun51GKxc1YULOHULE++
Pi1nPiqqCFZr0Am356ZdgyiLZFhT3tcSWNaBjw+t0mhRzNZyAOfJQR8IlotIzas0
ZFyJbgZ3hlFEhtHXGzdXepMZmAS99woQmC1dUqpGg26qqPt4Qd5zGkXL8f7aV0eb
`protect END_PROTECTED
