`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gZlUgaRBFJVusmyHTvbfO5EecmFp7eDdkHwxDncbxaSy8dRnYU6RoUaCnR9Mv9a8
DqpzlXfdLq3zRqT+t8jh/X5FwYdHJ5DKTQFkpsB+vCQkl5/aTzZQekZScDBqT2Wg
FpY3Ci9W1CsZ88lRmZC9tD+sNe59F3Y1SStbKRmGyv+iGrB4Kkq6G99k2iaTihPA
3gs88gWfS8kQOgx0+hn4Pymc4I8GYXVdsGr5qSg5OTIkIUK0r9kpJcTXulunYVyS
DEO+g0QHUGi/RIReQvzCJS9GD5oyjrVhj1JFP7WlOCYGFLrS/BP9nNbNfJnf4oDx
yXw5ou7YH153NkuJgIgZy4LKTD2mBD/CN57TznQp4h5ENy5kxIASAS/tGhDoj+vF
VlRS7TFHz6/APwKjlikCsO3G5vLFi+4n0kfr5/jWc6f56YLRxMJk2CjtIjH41h7d
2sCUDmIXTdUqCU9xAgARS5X58xNEJwl9IqZtkWWexGZJFz5Xc1UrzXzBcmb2gTw2
BpW44ajegDxIfm7hN4OZ+/EEV0zer6C5dyH8n+3Euopf8ELh4hDPfOx/wcHb57t/
`protect END_PROTECTED
