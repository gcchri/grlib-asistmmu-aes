`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7f+YkKT4xFmbAsRvvFzjPzaa6bSxJI05Uofa2DfflsKsoFe2ee05QqUoVsXH49wb
6XyRXh7679quH2na41VaUJugpVqo8tBOWL6uNIiLryQZ8pm8tWw+0zsWTtMFydfn
3zsXRjCPXzAOTmCPrDK5yez0A2jvRl8uE/qqvYhJ8ZUDkVb3t+5+l812BSgqfBQ3
964LmvdD6on+FO9+4T5v2azPU4ox3ZrVq0W4Nh67hoqniIlFtnXnASTMuCkW641b
s9C6gwiRR0qdzxdFb7Zp/IOGHKbz44Hz8rbjyC4qf59YYH8rc6pxd1H5S3n+H3EZ
I7S9AbMhls6lOJPfB13Wa9LZIox1E/r8j22Dk1pRFR97H8ioiXxw1cGMaDk/Yu4C
cDrpIA0B7AUA9WEyZvea1AjW7J93ZovlIC7VCiV/FxIGu1cupi0+dJ/wRndCRg2a
3Nh9hNtqYiFdnxp5iGEx/gmQedgkmAVKXYZWs14TGlnJz36IfCrqWzpjRVCHkIeC
uuMcJk55UPYmT1wcEDrk7mU+yXThsbbCyh+FuK+mA3ukMgrTrNk8fkDzfbIuhLrX
8KTCwpKzu/7FK9KWV/j7PAyNPbORDxZeHT7cA5FHOskt3b2sna7CmHTHpP4QjYKp
I0n5L+CKDo4B9bSfKcoT4u87cyOp+hK0kKzFmFTygyIKb+kjlIa60ksYgvACKkl8
zN/cXhpTtjXDmx3ty88j5PyoqVTTzM1E4qhXS5/eCTCkVm/MQDub6fFm8oEXnzGe
iSYsV+uVNlDiaF1EqRr9rtFAvnaiiZa8FyMh3nviwvhVwdft7UM1vn7TrmRV75Q9
HIWuSvTkVyrGNREcP9gfZ35GKlF5QsMb5SeGJgppaCVlhI86KttMOIQdEYD8FFbe
Msq4+ycyX1dv/l+plTyn56+ptRSrvZe9YGixPr8xGPRrkZuVZUQ8uKvvFlS0b9je
e9J9cfS3tVf1AWDoXNHJtylJu9Y/P1tVtn7spPBP1bkXGOb2UDcFvFe6qrBYvmr/
3W3Lf5prW7N4m52M2WvpRIdd3gSWuBRVxLm69RNO0XijQ/6VPZdK2tuCBKrXW0YM
NMeSTZWvN8Y+JvStVYiyumz0/4mtzFvHd3C3otyTcthx+wo1Xvdq6XnnlkMmj4FT
cuI+MvGFmU+QNACimReaAf5GvsnFyYa/4InFUkdugF27AylE39/bUukXCqqniMwm
XZX20HJTH6/wVB/JflSeS2Do7pRcDLi1iBNHb1CN91ylIejkAstTgCRh4f0QLyhd
gEqebGQM8ZdI1XSvwoxbkxWJW4kUthLKXlMvj6Y8izSUvIp8pdkcCwQNSHLeO2ES
k0rjWv/GymqrrmD4pzKEr0k9KsK4DCuyYDrUkZJk6lgSiUycc0qomnWckvedFAAW
51wEsda4wK3yUvAzMgKPDr6Q4Yp+1CuDsX55vhNRv+7sB0n6JgxOv56zBoeXjUw5
CmStXmx12/uzi+YRImryYCQNJtElFX2tWQzUBLBJ63S2ybOtxFsSDbE3T31Y61yD
snlgiAOyDA4dxhv4FC1JNGX1g4rV9NItTtn0T/zhOQKLX9ovMs5xoveEhuvbuF5q
D3emcG8sLSYxq7TFvfxbK69GSW6n/DGbZUyV87ajnthnR9jiLdhl/UdUy4AjZXnp
ieNh2hpuuG5nTLOJ+VpxW2oXN70o3NYBqXqMke93SZCPSjHXVO6Xu4ER2ziLlk3W
oK5C2bKWS7EeaNNOu4tzMN+l8d4ngh2/No47a9MXZIj5J5NirhqUFpEly6ZCeMDL
r44BY0huR/HjlmYRXnexkgYsaeTI4Zh4Ht3LE3l49OGA9gpyNHml+ZrNdras7Aq/
vxkXWf/mp+DOLEQW8HqHnEN84z1ygWa2ZwYsc3Yi1En1vQJ4rbe46gKxGq1e4ITW
6SJa4EflcNHBdfs3jc4nz/Khe66TfGbIXj9Jo8Yb127bkQxpBuQUbKYeSsCOBVsX
lqE8TwDMH3ApVifLfleyG7829qkZrkGuGwNrqmd2RgFccDrfe56eFk6ooRc8Hjoi
Q6aeBss32tiGVpuIHjE2pQpCIfJGlGR0F99ShGUEaDK+nFABYjs3XKXh6I82GHiw
vhKjPoOeX32wnqD3wL3Hc4zG+mBTrEjU8+gqGvDEzbEOQHjSLh+MmTfyzMXXTYmz
engJwyl26i9mBSMVD1wwRXUSNiw95vqrlrlacl6nN2AxTkr0qR/8D3GJVteJTOic
ujygAVNV3w2vGZy3ZrIwkExG6RR6hxp39DRSMglHqZtiFcWNRShAg/B6LvoKjmQj
qhDmqBDAx2FyOD3U/NG3pB1Aw00tdUfpc1mUNfAnjAA81OkWIUlH1FROvdUwJyhR
tJnqExYYRRWoh+VVQ+w2DKXscFQQctlRpPfYBLjII7kdFhXybsMFhqdr0rOeBbqf
7Y4pIYcPOQmHNtsbAl7iACRaYwybb9lChtlP8YbCzdG0kF35zrE6Ny1FPH+gjm1V
rcNIbiNgu6Y4eBgAHcbD6tW3x+NuYM76tWoxSbuOmVEf44EvBGTp17DikDZhiv1e
XnqI0Uj7VjtQupyhV7yVZveH0Tc1PfkX3KgnjFDOulxrQupn5jcrMD6a06xgPMDf
vMefKsqByPxQQiBnbZjPofFd3ahvVvWlpFHblQB1CTyCWBsK/sGwTHbj+sqc4rGf
zN8Jn3+iNzv1Lq2iv5uWet6Vo0cPoGi88BFbSXfjfAE0j11tHg3oFFF9vsAm+s2A
CbwzuUZ9Mvef/CtqyMo3V2axv9gwds9vHxpvSHCMF3jXW0w3QRusdgq5FH9ioAg9
V+RldoTmrDPnJ0n5ZUI9wg/e/24Ie31GjqfDzc5Fc1k=
`protect END_PROTECTED
