`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zavl7/JCpaJhXyA7N1QSxuUF2jnlEPrmkFA2datCinl+/rUrtDiHd5uChlmvknAW
I+hXvtDl9s9IErY9A8VaX81MJh9+f+sI6NzJlI4YMbw+QtFdxnGPN1TksrlHoEH+
e6lm/ajA4vwhDKdYhQ++k0JVjQ+GKQC5rrVyeMLxXOdKK4ZLq4eQvbzwFyqjzfRs
ntTweFBgZk9/2I1m9eSksBwyujPUOKkNv7MrVju3UQiH8hZEW4B1CmMycyDwEqol
asZQpmsDFC744wbbgjcWtsVIm8cJAK+QvFtYbcih8kPFrWEoIGfPrgSa5EgCjEq7
StxfaOOFI4fnpy3cMlXKff/p8+L9ETJgIDhjL9DergAFJUbCku3TlpicQQ1a2ZDi
tETEnVnn6Wq/ibFb6AIm3wWDJetWvqv66IoYyq37KmuSWtkPzDKWrNGjkOZhIVo9
o0RrVCpImj1SWuTX29uqwcgJb5WlA0s9Re173J5zjvoZjaetYGwhzWS5kufZ127I
YZeApxvBJvrWHlwhQi8VT4vky03/S0xI3cH39oe5nhWVnxr365E1obzxWDTd0oXM
NnijHfAyJY17h4Xf6oZMzlGVe/64/v3gUefgyMh9oDp7kQ4w64ODteH2anSwRzNm
HJOcZKSYJ2xMrgjmzz/wpWE1cLlqNyJtxqDBdmsOLCxWsukZp2N/qL93021e0QEw
PKuUxNxKBsKzKDBKSBMaPvMr8uj/OxuaHqIppMuZKj1b3G7f8XqoUFrOu2QQoITO
JI7jrF4uf0IWa/ug+DFNpu00kTk6xge5vN287PEEzfkXZoyYnMzUW+Aeyp9ofCQR
fMyAmsbpg5mxc7+3CuRRVUUyEAfpMnRjabpQAHNAhtADJF1qoSiWkwjmo++ShiSg
hwvHoEtxXcBSa0a2bOYs5f1O6svBanVBP3kzG2wo2MOuMX5IGkFetZi2YIbyfzRQ
FfxTLi5a4m1Ch+eB5vX2AHSKgVkI0T6Drd9kJQ5n7/RnD2/Z8J2T7Vo0a1n6WAX1
oNLcbDGNEfVS1osXW9wtwvYIOOBv96RkXTOi0/KWf+3TTVkoATxoIieYTRYUKxUL
T7fNbNhBo3+tZAgY1SfMD8Tk4YfqC6sqdDcUBdBf422veDnP0on4MtaUp8bEGBCT
bjQhogiqaF1W5E8f+gZblRm2uf1Gkm9nodqqm2ALnvkdN2RaUbZV19y3m556pGZ/
ElKFxrze+kxEAiuYiAM21fiUGqmMJvSU97G3M/J5D9jBgtMk9/CCYDmDbXjbRTeR
cHtj0C8xkKlNfaDh0zgFddhaABHruKmnUrvyI2tOHI8Zaqmbd4P9qp0/ArFs92F6
GzDAYAfk3dd+CXMmy2hI271kNlvg2vKMSWGkS5EdLwustWnlb6RFzr2SiVJCSRpC
3FtaWjBr1q7rin45m9xRhTKkCyt6VYaRw6kuV8OJL0jhV+16qwk/jEdPg+/vpWJ5
w8CgmcudM02U3/OX1kYKJ8XfgYo+hbG2cxk9AbBEE5A88wu+OkMHCxXY7TkzA8h/
anKra3jvs/pQfBqy7BqpNOnUFnvRz3QHrwM3q/64F3v5Nm5b8RmHy/SjdNOiv5Jm
3uzzSYZeVZFCwpnYgoCfK1dFOGFQWu++e2kWLvieokZP/wElpJzONpysIqY7DR5s
3SKDOdbDaIpfezsRWSRK+DrqgZpHSvITML3rf7FI1v0NxNpuy3G7mceh27JjfurI
bJ0EYf75Vk9htjLVwinUumuxJuQbQKjDlT4VNT7UcQC0xnIQdF+gi5xmlQfunCu2
2kzlGkoRTFGmQ4JOe3FUJUxJzg0S/VMa9ZCUalovan3O7Oi1YlwvmCkbuU3PZV9J
e2lDn1XLWYu/pT8Il4AdzO/0n0OXxbxQobO3KRxY4uesSO8Bn6K0GRGfKQWOPuB+
dBVlufW0TAT7+YWfsJ2fGDlOq3LX7G4Q2BWXTPl1MiRzp8yPWF+S6AFoAzY4QI/k
kgXzvJgXGt2UP5Y5/C59D5Nws93UZvU0d7b23pVuXPV6W8vxgANmVWknHKdKeGAI
7iI9NqftpZpL5yscrjY/H8bM0UKaBUgKEcNrT00I3xLiXRhl4Ll9UjoL9MS8l4M3
zYn8UYtD9AGks3OAI++eNdZVZHW+PDcysTHsftzmqoraRVQoLLWPkjUDOdOQq/E0
t2tdrFWG47nTUXel4Q+mymTH/xG1Wa18QsPcJ/ylKq2C58bJqFvJ0iEeqdjZlMPP
j8lREuJkU9cZPInmO6BcWc3CvYLu8oQ7lknd2LA/YPkP7OrPZO+jjYxysbdShjBz
53utT7FM/81YBUq0RZ8azxO4SRssyecDSzeKbiQ4oyYBsaa9mz040tIr4WCQCeEu
0Qr8mM2XjPXPEYVRMstt/zYq5BmSF7t93PO0NzLSwX2Vrl1/t3f3BJYkjfKB83K6
dyVTShXLOo/6t6rfE+3yjgKzP9NU1dr2iP78aRBgoL/POMq+DNB4XmKcDYwt26nJ
bInPqMn2v6Xwmos0bhH158R0LcR91BBZqqJKEgGtVIBO2qoPvPsiyxVAFrG3/diT
VUTePSPee+HR+3LNEPQTkRH7BMSEgcy+vwyGeAiXTAhku9NnW49ZGqVOcLdcZCtI
QBq/POMU4Sjyrq5EVcCHFUewYSYe02IX62TKC8PzhD12XXQsuK2fz0sB/fblkNdJ
/prdEBzaKtiX6GgmznX/c+V5xnFhgbx1HzAmdermeULRZsju2FKoSI2G469Gd2Ar
WH4s1Ko6jn1uvmoc0nGGHs/sGaEkpVtNLeRTJI3n/VdIasz86o2xDVM6ega/2R7w
jVPQw3gfkPwr9N2NWPXa9wH67umjzlGxKOoADuSUlyPHS39KxaKtUDiBsOBHHwty
Us4avG2jiY9+rqcSTyy+aIfIvysHYkmqvt8ovGJ7ZuoSccazpc6m42ANPm3vca4N
o2J+iwc46BXjp619W6lpaWD9lGvCy3bkXR79yeMNqwbQBFnmTvHul6W/QOsBsiEd
bQipFaItZe+RYzh4Ump5zjvqwLpoRHbiOU5XjcVQPg53kV0zDYO8Yc17vsaoNjxG
NFNvvOLjWK58v667NxhKUzOnC2XAYEeoawEZ1Zd3oy2TNkN9LAEnI51hjOw8k/JW
cv1tG/0+EgtHnh+JJ3buoA/ScVEsZ8xAfbkzK74Nf9kI8MfKXDLlKd+kDCMzQ9Qq
KtcMrxfLoTeHEKXrvQRo/afd/iMk0m6uoz2Ra6FEyIA5gLW1zASNKapbBS2rchM9
1sGYApZn2vNLvI1+ecL0oaaFwBsaRKuOv8AukTH67A9UXf9jG4hha8Fk3HnrDX2h
iq4l8BHRJEgmkDpZjIBdvjOF63fJJv6hqLMVLMXI1hFLZ2LrM6B3kMF36t3ZcYJ0
KBW7+OBxp0XlHw4GIV2uXcOcSv6fdUzxonWRl4GjJoV+Vq5bzoWjJcG/9lgiBlGc
MAG8UGkr4Lq9CrVGkmIJFAV/nLhjgRvqmGcjVxfV1KpvuQ+MfafjOGISqdTtRiRo
3NTzbDaIng/pyOTiZ0MuXE2G5EU73OOCA3bxElJPT9IpnZ4UWxiGowpubNcPiraa
0S+Xxk0ICDxug2AHKPtMNPKiyls0OZX98wTO3rfD1pILqpIufvcrBeYZg/g8FP3z
Oz058/LJlP3bO8rfNct7X6RZqEetpBQeHCAmmFcht2BuQdzioRYtjtvVUGxIOoUH
YXycE1o/M6xsEqsVQPBXEtTtHG3v/HxhzemubTtdQPCBuTZpwVBCaQzDSv9IWOdV
NV15deHyF62J+MZ7TAARqj6RAB1mbEg8IDNFVWMmE0b1v7SWr63VShYXmyn8U6y2
LiV+AVp1YllcSEu3Z8wh4OJxuB5vsohl9F6kko12Lm0KDZVjSRyu/3MLAD7V8/7W
IohriNq3LbxEozgfifs57rfa6wNfmdtjHGb5w+NEdYlNOpsO+2lYmpANbtHpd2c1
opi8YYuhamSUA19FdXGFybKIRm1bOFWexp2qQeJNkqxPPxKZNIYJV+Mtzj0MUi6T
VDGe0vVT+aW/3WVkRCz8Rbc65V1shIwXDnrpzsimyB/CvvXrZSd+PEmRPi4NIp81
dGMQRJLYFPS5hlgYgrh7YxxeCsdsIt2jj4KYLmI/nUuBdJaDRVx3HTfVk+GNkbAQ
H8h97JuVm/u2Fe7YxSy0CvM5il5QtoXMBwbTM6q/LpZTEFljjiKt2j8mp9hDYs9K
p8NjKFeIow7E9WA0uWcJdtAZiRCmqlrXINRM9/6QUyz8dTkzv0kSbdJztY5dxjrF
dkau7599obEz7t+cmwyTnGPGiMu5/PamBJdM/yUS94nuBmyzRGqZgGFWaNYEJA4o
pLnVk6GstwqRHSrxnAk3iLFq22UwY2yD9J1zV+w+PnT6ArzNGNEIrAYJr4WSUaOH
8rfAHWBjE4IsuhYljPrM5V/bKJsTt6wsTOx7qF5Gy7DK867fFtgcHXZ/qHJ/noUw
CVd3coxnaRZOIG5TeeqJVMD8LMqZRYgCW6hy53+dEhnavOH7yuJ4OmuWR4ug4GU+
GqcsPsMZjiIiX2440ChqkZTBMnXG/jqwJo23HdTccoxz0z8wMbJkYz+BzVHf+lzO
fWOG2bQGexvZtDtlCxW8BmR5aG7/E2naPTnB0qUyTpoKSIDGFNRzJRT1ChBfo00R
3Jx0lg2vCfg9eVU0BvsnfUSKu5N3Bl5OUbsu6psrTG7fNiZIGcssE8ZecQOohgNF
9io1U/S5UAFZOrOjrPzhYyD8+pY9TrVTcy5ztZsR9eh+0flc05zDT28Ak01WOyE6
TMWq1C/zIjyv/Xl7R2P4ZCHw59opOPI6ZIGwzqtBs2mSHtq323R1x8Yji7SxWARE
0kU0Gqcqy4bxwzHv96KcRr9KTA9GB2fWR/rbPUG3XMcO4fsVbiPkin0wnRNiWDAh
b4+fKMOn4YT8D5RXWcsQwtwE4UFEDma9TIguWmV9+rFpS6k7A8kyURAajh9W+Zb5
+5XPJGlxyy7NTPOrtXZM8DT2cRTNfdeYNFOmQJ6ww6y1vCTlEyIcwwFB/2t/0+Gb
sjJfXIEWt8rl4kZaX7VhUDvo0P0DA5MHVIJUB61cGsV0eQ8fTSGBVafrrzXINxI4
Bw1bdYcdJYB/HemkdytEHoQ2GNPE2/FMWMts/sz9Jxpf2fuGKcQPHaOYuxY+bZ2H
wZEDs+l7F9mNH6qmaZ0H9YDwd4+/v5NNUx0x7jek5+J6hHqb+krNK7/l11iZs6mH
PIvv0Qj6d8J38W0DWdJG2ypdThZEKj8IqGAuyPnU0WjdLdSq0TB7CPLV8Meg3Oph
9mh7OFTVwNx9OUYo9JPe7g1w+ADaj6eRGPz03o9wrVFI02bMOJ5VcjLLE7nqKOw2
HlfguIT5VqkICdE+currGtaqjZJd//vh6zR4ZiovwgC8VcvOY2iM/RVMJRLuFVG2
rjOF3xphubBWTL6hPWdngPKp5D8ZVPhZFqdDwXBSBT4HCsic/leRpHpOtLTvQLxQ
F1WECYLmtd5YXudLqmtxU/9hq5HEs7tnDu5DusJctFPbZR0GiIcJlrbsuuH/M401
56dVGikaj3duZ1nSLv8XrwsADk3O9TFQte16BbtZuuoSZd/weSnmtklOxqBdhUc2
ljwzURk3A+2d0S1QpeYeZg==
`protect END_PROTECTED
