`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7lYRRYxE8l294w/vTs+425TCwkmfdqDYtyKTYs28BaFbNIwh/QnpmpnSJRa9JNVX
n1xiejZcA3IpwV8wspkqTZ8LMNVPxIEFI4atmQgwfw8icwk3nKl084b0CJ0C5XEI
CBZtJ1pwyH7FcEgjsugWHdVKBWoNjjFt+R9IfPfC+zIR1sODZRUrjmLiI/BIR72Y
5FxI5mG/l0gTLlyiSLKDcRBct49F5ovFfNl2t2w6EOXqvXgWpu7hF/d8v6un7oWH
YxAF/cFE1PwbqyN0tduFvgss8ThbatmR7PJCR1ZqMuVEM3uX22JG3BE7JUjinaY7
ZwFEaVmPbti9t7iGkCLI/dj06CYn5ViKHlC/nb9Keq1Zj5byNwMEXn/dUfYCLsQL
ZPo4XVFBsqmcaW1r0vehknKgtUAuVXOdPrkCi6k4jvNCLB011+YV7NsCfJufwnxS
7FBJnLklC76MpBFhooHioup3s+dpLYXzLaS1rkVABIl56ygftZuP+3kjEaJ7fkRP
iOA1pqPG4rsdJMt6149K4dWw0ev6jYfnUVJoya7/VdwI2JL+WL/bG3ggSgJetULl
TvAOnXP6yzHEmGCJDHMqE9FZ6gxa+GT+glHMCcY8sOKuIbaBeRrfVL3I/UFqe/Vn
EF0+pCXQk6p/itMpC72GZtqnW+ipo8sJKJu7HsLcso9kiMjggIX7hTWV/f4tT2W6
6VfnRIwiUcExn1FpIAOwcKN3DKi6dYPwueb9ET7AXofVF/aqyVfwzazq4a1ZwH8J
lL3Oakl0knzc1WM0KV53Gv0lv2s9zmVnME/Da2WbZ/6UQTISxMPQBGYqIhU9GGjn
izc0m3MYwkfX247LTC+kZSxErF6pNPWLg2XBH2LkRHAtXQ3Bxa1CxXC8sjwadXUR
qqQUSuAmTRIUAmgFETxlKF5X3CW0AFGoSKG6lC6BhBi4tK17N31A8pUyQJbu+0CK
rjrAMT5pBxrVTFDvgqtXEd5mWImceeLoA4tYG5/wWn7vLwNunRCFlgdpCY31MYLZ
9gdW0C5Y5S6vAsZIGW//7XiHpqznGibBN5a7GOyx15r/Sp1fWDroLOqU+p8EuCXU
FKzSb3bdaf74RQ8FYwgpjQ/bWTQUdsF6hNnyrdxaIG93dkVVi8BQXrxeS67iHgIu
uDZzydSH3yJcfiv9qenT5ucY5uDSrXbrYEklQcG9dTSSjDMz81QYjuAnHEBha5GA
4En3Dj3An/x4us6L6wY4Ty2vDekV0lVCsNjCOlroUkp+6qjru/Iyti3l8ueNAbnp
LHGlIBZJAspGydR44l2el184Ds39gttibOG/KqtvEBGDyrqAG38qRQX0M0VAYhzb
w9QBBGoOIt4RJuAkb1iXAqB1s7Y+xHRjS7B/pf4UY7GuuejomDyo0C1lBzCITbuq
+gZZhYEwxdjneZdcrSijWGr3rGvNQlSSp0P3h1KwMMkpctJcISHwHr/Rny4gEhQr
LO/tWuHlHAIzvqn7qH/QzKEsrqLlj1NZN3cjG+7hCkA=
`protect END_PROTECTED
