`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0B1U/RreqPJk8fShGhxcPFRpqVeNth3xT5HvWjZTecrFL7WHjrSH4Lwr1f5Zr0BE
DatyUzGfHjGX29W8YbmfZf7unGm79Qz6VaDiGin02H5QiAb+UULCeOZTRk35v8tm
gQAxrwsLbWkvR46zaJ0UVgxFF9bSZi3hVHVuLoxu/ejtL1aD9YuvLSf/iCUSGXI1
+ijt6Y6V7FvNVfpEgGYhycUlGw8ct8tzb4e665H3eSEpDeuzvi6D85mivObAhssv
92wzZQuChHr6MLr9GM1ElWmhnFwFMUWeTUkvh6lFNRSOsjfZMgd0JLhBACzL8Hiw
grjoyQsxlOqt9w2DXXSxR190p4f9RxDrjCzbn/+KNiSinuGE4oLbQ6RKToYmHh1W
2IfOhw2GEJnI+tf6wti1pMkoV+JIfjZzSBdq6/9N9hwwwmhO8mra96ZbgCsy4ihj
`protect END_PROTECTED
