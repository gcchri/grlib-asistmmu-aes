`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wsJKEe9yWS2wqG7mbriZgtGIrCHE6w6tsWzvUSxEvE27KLk1349WU/Ezmxp6fAw9
eLSXxi75731K5Q+6p/SRcDgATVCacwSnVLrmyRb069elJawX2eAz964zZ3pNj8H3
ZbxRwcy8abdoIDQLLG24C3kPTdoOclHEontkvrCL/H1GNuLm4IBNIJiF+Lizo9jn
z829dGnSLL9EnUgenaM9UnJqmZRd3TDc6dfz2GXoI1+08g8863JQn/cFBQsVO4MN
OMp8HqMo/W3k6j3MAlSo0ki39+yhckhIMX6xsrYfJwNgvBZ9e4kpiB1L51k28/qY
IL5pAysdSR91e3CLp8GQTtjpVybJqfvHXfsAXADmW1eXyQkUB+aAfjt14USZoKAz
bo+ou1VrvR56P8AK2U5TgjNEfbjymTCKOhuIgHREnrglf8B4O/F65895TzF7WhIQ
XOvQAEU/J4ZQtfwfSGnCUDgu3A0gvQ6HrpRYDDBR4qM5lV6MDDdHI6VAcWJqnfXJ
hX9XNPfmrA3wuaR3Ou59juoGtD4IwdUFmIjAXTj6izAl2fhfOi0X9hqMOHMcF6gl
vdl/qhUR1UhDkrRVzh9hDENot8BbzLYeQSBfeanrVtnG8tl1vKZKY69RtPp54nxF
HsamTJd0Bx5kdr9al8FKDXTx3YXI3Lku1sm13ly2dfpRtqnhVzZ6+zO1JUgMAU23
FMC6Qk7VNA4jsD1Zx4jFai4SuHvFzKTqGxq9Y3SVvMpEzNop4dzx/xQfy7pC1rBY
lrHR5qm59u8n9c+X2aoiHYhaXEc3qzsySr24Us2TwE+rgi8XF29hj7GbY5+dRfik
NLmNeXU0XDIK9f85xUYugmR87v/csBdaRn+8z+H3AD8DwUWxpAQVVMckDVIIUlvr
0t2J/nC2D+fdZ4ZQXtOSQEAKL36aw/zAh+JDFx7IdMBHIJ1BgK2t77oGn9H/aP+Q
6RsQ4tkrovGl/Z8kOKMAQMq8OOJtJZJ5zp0eTOoZkzItWjeePTneQ52F3kWNmBM5
4l1nLp9Sa2NOr2pLrBJjhw==
`protect END_PROTECTED
