`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I43pv0zLBuhpvHWvnv1Kb85d2hrd/a/ZcYEVxeeLFd3EBHUvV9GppmDp6r1VEiwg
+ync5bX8wXaXr56mvHDLhHIj5PTSI3gfjhIMQ9ky4XaQ5VnlqGj8nYAhC/UR6ovL
w6fP1oxs846iXduFUTCKIToAgaqCzb02rCBXkeIuPzC+K46JkSNFah/wr7MEXwl7
oBc5yVQXDHiDG8DusdzE8ZCpfCmCQP6THVysIJY9fyzGOAxyvSAD2CT/zHPy/z9A
puPHzo7EGjoPKiBNw2YASP2xF+o2o1MU1OLLriEZBo6lrCS8q1OfytgOKYubyZVO
9vD/RToL+vH+xUaGsfuXQjycbLFkNQUKaZ+kfsrxuAF4i/jox0oEDC4Mh1cVxxOk
oZles7zp0k3LLPxT3X9wBjYtrEq3rMgy5mt7Q+sURCT5XZg61UbLn3O7PTdfrqOp
UCbcdcjQmxfUPHfqL9HBnmoDH05F1dzHQRI1hKsG2QwIOLYqBaFWEEOEzB8cyiE0
vNddokxrDDnLx+H4Zm2jS3gHXA7ZdyxEiPBqoocZpheoe9XoXT8VkAdmreAABR1A
+U/Dsyw68Xn8AStphP5Vjs/oB4ofGvisAEihCOGd/IdulNmtcE9i+qOxziDuhgl7
`protect END_PROTECTED
