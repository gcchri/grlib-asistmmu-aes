`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7RkTQnkfCLbkmJ03BWldCz4UCBJeuuRr5mEcrx+CZ+2vAh9MjrQEBS89Bi+T+1X
hbuaamsZJNmK0U08IW1muiQ3yB5ub46vI2KSMmP26rSfoaemqU+OKu/ZkZszmtoN
FQY2gLmp3DLwRSU1urZvpkFbOlvpGJr4kz/0iE4DEMfoyiO3P2x++OtU+8JOivwq
7zstssCF9YIgumG5HLhNbM/beP7Rj9HX5t834dLOvXjiBkrYBO3nxqG6RK9yF8FV
46rRmC8hJFqGTTrty1pXr5NgTNcnJqJiQO8UTPMuekgk4HayTRy5MbjWO/49pGKE
U6Yq7UNr3znDJ+i/qXzzYvTYXfviA3/yLB3A9BMfId0B0AvjsItWBAj1QVUiUMlD
GEBErxjkIZWw6KQ/hmvkZ2vS259GZ0IJr5hr71DjYw4=
`protect END_PROTECTED
