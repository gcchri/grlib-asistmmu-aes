`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c67TxFsUzf2wHYP8DTK01Imx6W3UvGFtogn5nzd4jtO3/1P1pmjjT2O7OO8WV8bi
oRtH2YNCdIIvdG0sVYkMMJS/DhbCkj39wcjLZHtCQ6GR5C3JOFI2vUCLzBw8XEq8
03XQ9qCQ4WNAtWfPTzVaaViMaJ7jjCLLoa3MIZPtn02px3moCAwcGq8840J2Ak+j
qYoa/VHaxADHbFcEAwQKIdZ/KhX9mIkcbT/K5GGxjMHQYQwmwI8einhn3iM7ISaT
g4445+ResubMJscx6VJGKJFFISCnu/BQptbHImIBl2T6dCenMheerhuBdfXzfhxJ
7kZIBdpRpLmfEVQblqNrb4/HuZqMk2p43eUICyLzniAIDNSJR7m2Za+3NcOPhhyC
g1CZNKO3k/dgC6kd/k9Luaz8admYOypR1ogLXewIgLvVJq2mpnI2KO/2LAy0NCD3
C6YoiOZvXkJcRXCdnksa1BaUQFHh7VlJJDCqgP1lvL8ctNfnd4o5csFAv06JZrfY
`protect END_PROTECTED
