`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5q1v0kQjJGQW2AHVfxFv5awA9rS6UJonBHO2AQRb6nkOlfCDtH9l1ootlVp5UA5I
cC4WS2uRrc6ogicI80NUg6CrdU4Ay65iZQ4M2R3xOuX3eF7fzOyCIaxl/XJePI4v
1rYashdpHwUNDvRaYTiGLeCuzSg7ZV3rF58cf/MbI5iVJ/QWfDtb8R7+ubjFOm2H
bT7AGz2DyYxOvTb2aWvvrcUliU/GiJX9q9juW5N2UuX/iGchgl8p4UlSiXy16YVp
nKQBfVSxxox1XmC38nXtemRcZj2hpswV3plGRI8Wd97VHKB9HliULUdYYxIVLUea
vCPZwYOqEXctyP6ASLa3EuNsKKDGdOKWBeetv1avXSCRrE6dvOCx9kebreQTDhPj
92RgF3zDSQGz/HQbH4mOOi+vAqoG1oL66w2ObCO0koK9MbOIklbuVgVG39QyL0Cy
qCAXMhZXAxtZlAeyw/POeC3ivTZBAG3H3fs5tM+f4NeiDSONY+7sjDwMOW7gTvs+
ZPh0yZtb5IDjzmAnXObiLETNCDOoI8uJ7M2sLLjkQONRQPz7/a6m5EfVhp/7+VgJ
fC50zAFswsYyPY46UWrkTNTSqZ2OwE3utZQEWC5gaIBHgPgDn+SYXBzfRha0Wpwi
ao0ieNz4yM6ktwiafjpI/3eWcwo0iEHWRDrECQFM0mg=
`protect END_PROTECTED
