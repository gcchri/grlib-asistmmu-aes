`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qxc71dtb7SO1XanYDZgFTIcKhwOK54GELLesnnOS9kzlj0cw9cg5hNCK6go1rKaX
Z3EubLdnXlc9VqF+n+xcQY87NRU7SJdh5IaldunoFjL+QEx3tENUYLbppt7DpMKT
1J38U0Ci8jDdpuP1n/eG9ZTqWnf1eYteonwvXbyVuy4XRNc2y+CSWhvf38vwADg+
9AomyNfa9uNZ8T+Ytb2GKVlF7jtOLTI7K6mE04dVOSd40OXorDmS0BCznUSZJo9l
OSIs/n8yGh0R5Q7avnoasPGgk5w1ZpZtZBpsK0+lfjabZEVjo+e2JwD1NbPlvCpI
g2I8M5E801UGnqydwEN8fw==
`protect END_PROTECTED
