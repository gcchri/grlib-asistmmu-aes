`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3WzJes0evn3j1Q67RUc4mkgr58MnOUPTJxJKafWyXUUMtqsTTrfb08ONvqquJwa2
8eKnz6fPh2wItdtHT3riC+8dvD+C5Sk1rMxK4GsJA7yIh1igQfDxGTpKN6WQDLiR
papR3BKU1D37MpU/tULGvnZp07YAXaQBiM7Xx0Z3bf2CedQV+WB86T1pVBd9jmv4
yWogsPLbGmrjVe58zXeioNRJO0vLnbm4Dv9bR6NlQv+5QRx5sAG0wq6RFCm44XpO
Y6ILIfrAqWTmmhZh3Q6nA55VsbetNtvzAUmb737GGfBWzhkxyC9y+qkBaBg6vGOZ
HkQg1B9rKC8JSA995lFimskJDIOBuurP9QUYpDYv7fjSTyV2qDUp/NFFbq5Bd2hT
FaoGarqTtf4Kyk9h+EDQiM20JvuTWQwQY0yBP864xf0z+cvGxJJPq2OwmzRBr9H0
dKyKxXyI07rWDcxcVGASGxtiwyeQqbndrNtB6NlbXaCHQQIC7rfhL+jSpkPBkARg
PKL1I7ieTLIvqHGLGj4DWVP7OZBNx6/WpdmPuNM3uWMBykKich9eAMIO1yX3zbhO
dVaYqEpNLqT4Wo+iHaV+2Dmbutxfholpgk6Lu2iqTAPJ68hY7ZHZ0WMV7hunSk1C
d8WqyWzvAOzT2FdcGd162P2rf1Yh78bOMCuseeczxEtclPmkCbeTOFgm/MczSIKM
JPvquxF2LqqvwKIO2LPPJ0zEMZ33NMNVMCeoQHee+2TrmGk0n8T/rkHAmryWP3Sc
HSKNCvV3KUpO+tsibj0SfaDXJ9jyCa0MVxwjsOb39sM4C55z/w+Pzw0u5K31kkZV
/ooRdDIhWH2ZvLpqjajp0HGhWRRzkvmyG2rxOn8K9+SrBXdv8iWHBFyius0Y9Hiz
fMJ3LEc/IeE3l2ueL70ZKQD9k/P/cPXEb19ToaWWVq3dk4AJ1uh9vuT9Dr6vVXCL
71KTG9p6xzNfiB73tCF2r7c2ZDVcXGIuXZ2H4GqaLci+hvg/qAPWy6QY5RidS6K9
sthAQechHyBBJBFPVd+lJ7STOxbqxebrcSCMpBBPLsuL508h4YdQQxMMVwLqfHTf
BtVPrztIDomHaxab/eD2a2Z5pR/LwMj2fuvbwbbWv+EJl0FyJKJeu6BUdujWWwEe
72lkADfrJZrW5PbhtJuk9zQB3Rm0kQHvHZ5rpKJffpuzdoCRCqwesI+fv1FEMUe1
Mz2mhNYj8jbVV1zS+x4LOaKnMP6Ny76EggYZGN21N2OjBjHc0CaprSAvEkU9H0J2
jKa/sfoaIvGZHO6PugYjYIkUThbiyi5Rw/P1f5Mw7+0TB/ejxjwgXppEh17/4i/O
nrqSuYmrZWdMF2YAXFkiGzwaQYQSIzbUlcXClPUDix6Tql39AvPuonIUkVTST013
N5z4AMdtO3Ry/yWQweQ8wgUz59fDqDi4m/8RP2Jeg3uvEW8lazwVF4U2woINKciX
ux5ylgux1qWwDaokJxa3t4gaJqZiaZE7EW62YxUENVDLhWfl+V3loRZuZz+1sr8p
h5iuhklphQg/IqnTYmBeZFu0fD5ds+z8ssxZ4iuvB8JJ1SnZVmwpVOv+xK6sHmIP
FLinwVfmFyOf6cVCZN2HuKKETXQJMlmdnW/CQVFJKiVTOQbjzte1dQTqodAA5yFH
Hm0h35m4IaJXYZrbNsaMEGzMtSUWKLiXUdfxaiDfyRlrHJFKlvbMGG5w+PRktThM
9+So5p3KuC5BEkkOuwSCVT0I08MYDJrrkdZnJy8Nf3tbkUoFxvcltBuj+QxBC3kD
DelDrITD81YcbSh2mvy6cXbuhXjQMp5pzvnodbbDpX7jUkouGw6qOHVOyOfjE3oU
8Ce0nArQMpJ0fm4JIT6dWeYMi+ZVMtZnaYBoin8gpXxxmYY85pbmbvjsBS4xPflt
UsVsz8saEDCwcU6oqIjZml55tHUr31QY/rRUg/Cx3B0wEd1BeoOXGwjQaG6t/ZJV
jDVliQXVPI6Eu9yEvUdBhySUldcohd5xR8gjm2LZyVE09ptdILgMfiNVHzN9dvUZ
sjLZKoa/dkx9HtqwVXts2W67CjRvUuLrMFOEgINlUioViwfhrUmt06R+JWDYoUhw
RSRRfLDlgo+1f9+Z6Z8sRlJH9KIPzX5lSWOtwrv7dd6z/sprxYJ83X5vhenBxJvK
Ur1a2Qu3N99f5sG6ve2xXQcItu5buaoxY+J8CVLc0JJ9bL0uBF9qQ3ZyIAw7QOoq
ytdqJc0uqMFzGTd5Sp4zJi6yvKwEbaxEl58DeZlsU+blSc0NIKLGQKMusJ10KZQy
tREIlwuafLXODK3MwZyN2b/dXJYdSVLDuqx9lql6WUevLlwiaSMXM76gHr/X9e1e
+T0C50VISlyWKIyY+xxqyhRDAmaS5IYS/f6kYSzlNMmV3MA6JGb9UWqMXZKvAxtk
NjGTthjWXxejl+trQLPpOTTcVrohF3gKorcLyQt+z9sK8bruDxhkbr4Fp65+SpEu
PRiHodPO3xT3ZQmYmuN5uHbeac1CJ1PgkpGQ+X0dWtUQCEIRQvjpETUQWOU/2lRD
io9/iIgvsMGDsjF/PvsixtXxdcn0SO85htMU4SkkcMt+mRAIdv1rf/vonLJTg7HB
27S2VnSP/egwBuPltEf74XoFtQ/LGtTnBan6vGz8fWJV/Q+jhdVz0AKXmYYEZfuv
CvR4IB+p6h754QPFmZe7wJ5gPlFN9EQYfIC8D0aX2VFUu+pKf6k5JJEqTdrD2wM6
6g+GJv9G8bY+/3saooUFunmchY0KVtzuE76N8j76bTHFdU9MeqFlnBvqafo/MgQL
5oTeCO7iOr72B/iod4mb3DrUn5cqovQw7gz2pBVnjHeNhuhBijhwInagfbixHq03
mPA46El+6166lJQptYt+bxQ5V9TEfN7EGC8DpNJv6fxrCTvT9vC91/hX5poWugZG
gqzTPWh4ZPZyThhztI0MAsUc4Bb3xkuFLLuWTQSr7LetAkCbpa496W1YU1F9M2Q2
Hx5PFkRy4wkSTmNRp9L6ox0GGtB0IFJ8XZKcunBGcPgYmo8kcET82dIoJLtioTlC
O9ai7GvfGSTxSWq/Hx1a1GrlU6y0xuvCjT/oXbkUMeZQCLr1KxY4nNtvj3/bYeh2
JEsuLr7LnIRe2iU2zDja1JvCiEWsakDG83D+AQfmgCuDjmxvdBsQAhOXf8/tmpCp
6sOu4sikFj39eh5vETM7u5Poe1QcrnliUp8k69UuA67RpnhB+sXGZAb7XN6A0Pw5
Vw2x+I3U1fV3Wm2+LNfDjNdXkC5Oj/lYhJi7ayeZ3Ysl1HQmNCs1MIWOIPiB7OtV
Ew/icMMaVEieevVklGbmLnbnEaPndmxYfx90YhV1XoG/+wYTua9icy/hU1o1a/vX
CoaIM7MqtytzohLllnR2zJIIeQOIHYLq7bq6MXYslAZnJOJxHBwVjuvcCS09B1Ox
Bb18ISyYgLx3cxfnsWPdWTOoUPuP7ltv3REO6c2+qbxRgTMaY6K/xU42Anhrw2UW
hWI9GxXa2kGEJCGZqMyjcG20UpaBfSnOY9APzfp/O29Vs5spR/AqmOKTypjL9xVv
Qx9aUgAL5glFjsTgIrs/BUgzmX99UuucnnOC+HYL/lXk5md21sv0SYuSBz73quLf
DlZwbp5SnDTyMWVW1zvzMDjpdQ1jQO8eZMNxflB4qwg/Z09lCmgUL7QffMPoreLS
yvp/hT3pJPfXMKkLB2FZo4VYvX9hKGI6ZcBjjYmW7uOrVPiBaWA6HhYzjSZIP+fg
TlwC/r8BWGz3/wDTdDXi7OYuT/sSKfFG4tUH5MTjdfuakuj/wFoBxutgQTfc1Z2h
qW1/WPVcBwSqhGTHgkKzIqEgqWZ4yVWdclhiwF3K4ZixrFy9eLGUilBeCrNK7lAY
VUkEvTANIKWPUeUYYX2aYqpgeqwgHJX/1rNWwNE7eJEWIh+yi3PGSweIbReOCdku
nDjb4AHOGY08onLN9EU5BFJrnbZ+BnOj4VKTnE2tpOunpR51G3HDVRizha3e2Yxz
3Z+h/xctXrW6gMNTpP6qO0afii5nj2IR+zreeMN9iwl8UCzndiPA7tT16JvXlo8M
wLBNiYHoAlLsEvY3QjE6Fko8cw/wiDreVl1dTgZpFYRLvkl2hoZD7bwWyotgkLS1
5X+spXEx0wR0y2PE9KLMdAf9W26GjUUdsamXv8fL3HMVXMgCrxU8P2gzU4fChUpK
ZjkKT49F/t5HP0d1KJTvA004hqbdJXBrewz2Au47bLz36f/x/4U1cBwpRUn1vMsV
UjSYByynP5vhMpn08S2VLludBTTurT5DtxiCOvuKnL6HiuyU+RAnmi5qzvSjX9mu
dPFvVkRp+M2dOnlg9aCFgsANm2CqEI7aSA4jFJcUibntfFeFznmzrGeaEleYL63V
w8QDm2jtJlaeOFL9gleV6DXt3N1kiYt7B/S8JcSbvTK1Eb9/S3JEOo4U+IYhQ1cP
ew+0+qOEGkeKwbZO0lkhikdrZw3QAHq3lgGtchG6ulnjWn2OuXX+tzW2bvDahDYV
2Ku2108lQ1yfcSxuCouoc4s3dfTV8cMmSLLiOyCQj4Nrr95E4nOjgzpxvKYVO5TO
vC7LjwyWhupsv01pvGssHcCWb9hm+C7c8/ORBLAHM5bC67cEiJc3SBUzGrXW/kJL
nwExm4j0JYe/W+HGrxmFBth95pbGWZLzSBrvLa4LsiogiJrQnjkkUiEV5Y9ge7sp
fMQY8OuE/b/0tpQAbqKyh3ArCCNxN4jZQkoWbAnQZ+ed45MbGwCGAgLxdyiRjvY6
kn2LUartorwAKZanSHBnUJnl7qhz7tXpjkISFETZKnMRM8IsNeprusboBObkNfg9
smavoeqyzERLTq0JuvfYjL11DKukGVB+zGu/UbFZnKMh7yITQSHo/tvrl32uiuIB
Gq3MOlIrW/RGVhJjMxs9Il57+VueJtwfZHocY1/AZrfVOm8LhA9XD1ExlGeNzvlQ
tRV0S95iwXRAG4a5SLx31OJvVX2jFgoN9fT3MLTYrPQ=
`protect END_PROTECTED
