`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nm/FPxd+r/EHr0ZqSHXB1jdOva32tgX/iPfU7sWHV1NLs3JSvQbi238gWVUYyR36
7ijyQWiC0VOGljSDnGGimMHajVU1ECXcT2ZFWpbCKCQNEn6ov8116NA9xO8+vTHQ
COinYNImWSPw+bZDsx897dvSQXHxg7cRMur5BncUzHL1NZBLNqzzsGJS3lHf+MrU
tMVEkqT99FwaBATPaRTZoY+Wj4pY6bJttlODPJOS2+9f5whc4WBF0Uja1yAEFHu4
YTyTG13Xt2QsxDK0PuOvPg==
`protect END_PROTECTED
