`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LJ/mwMFzUP1UdwJNpotWhHZ92bztH5YE8QZq4gxcg3VTOavmvGon9QyyFb03L4rm
m3WeExKfdj/Vhxmnng9VcLgfWaujNOx2DbUM+OxQrgQ8JZYNskKkUrWOKHLF/m+z
TopiBic1A/JmNoFUPLVpg15imlLxqyk6Tpsh7xfPJBn4JCtSj/XV2wuXZFKXIila
s4he+hhH7xqjMy8k5/HPe4Bi5iu6hjaFOBU48YsSLAvsUfJFwAZ0aM7pxYQKI/T9
ny1XwvSN02EX4zq3LRUw/8m7kW//K0obJ4BYcNT4z8YVtVp/TUqqiD/P9htBK6ym
OQFpySlpYchXE/18QyyXamrOtWnrNwreMv/kMuxKWtUSZe/286M6KhoPKs72cHjo
`protect END_PROTECTED
