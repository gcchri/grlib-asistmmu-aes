`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yPOXfj0qVp+mFytC6ku8z2VUmD1ONreBN1MdvHQVDskKyTHMRjQLU+Kzgt83TLX3
CWM0GY9/a4f6EvSQQ4QpK7K7FSyVPJQeVxTDdVdVe7VTpQ3lS00rGMvnBS6nKrhC
aNPCsvnPgCoVyV7Q8Cmzxlu0X1ypPmz0wKs/PvRoStN0YCgoKlb0BhZd6INfq7VL
w4DxL3aUlTSXFjIuHtcfBZ2sG/ErgpziZW+C6tjlvkwBnLVvR6ZMJ7lXUMtBvCC9
UD4VWXsHPCfrC8QqTJSOdr51RuVqCzVIZyyFmbrY1QolHbiurm3xM5qd0ycZdat9
07njy9LbAlyyUsReHACKugIOlUe9c54QpurkBh5eZb+O57TlnkYjU43EEt9oANqO
2KtWD9bitAXT7ktopwNCk25Vy7mNoeaFLeOMHlMPMukvnA4CqdJQ02zncCkieU4f
j6rlUXqBu22R6MLv+5keD6fngC94Zz4SjdKM+Xfo30jMKneRV9vCpc8sErEBRE0s
eCPtxC2S558rVIKG9YS4tCKuAVbT2xww+vTDQHC9WWCcFeuu0p0iR8v7RprfNsOd
SFPBRcXw3Ou0JGNgCg46WWolHVgOP1MCX4f+fyoy5uVeqJ+Kranh/Oha/dxr8Bmh
I5nwvTxFqGZ2QcdBH1kV4j5VL/ElkE6y9dUjR0y5xLfiyuUVlvZPD3cQMdyUbQI9
0SzVemsr581J+FSmevti/yUhRnTkiUIghZiAHUPAY845Cc4JXoby5kLu9EVE0s5s
GRGZ9cv0Gcp+TnSQ3Kf0redkVVq4EX7UJqf3dW2tQh6DTHpc8WtnrVO4IMeEO7BL
dF39iG8DzuXM5Yl2qPLvlwCOPmnZKKiuGBGepKTqcsH28d2NIkZTxULCmmE6eW3P
Y8XDPH0AaJJyk+MX8QZ25YYaIMn8lX+WbeZYOEZlYlc=
`protect END_PROTECTED
