`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PQbnSW9zzsOwZxisjpn5l78bxz1di68GeJbBOSNzy+8rg3s3acAIn+ynVOky4RV8
exbUDTO9jhdv8nUAspAYPzOltjdRppUhPh5jBXOA5zjOOKqdyRzXQVKkKzPN7edS
fSZfzJbVi3OhiaLVeghtxqz+nYRoo5c1/Yadr1yZbvK2iO43AP+9w9XFtd5ZJPBP
vfotlyjRd4LRxkuy5eRdD60++StApEIWTdRAztiPtRAKDhyUaGbIDSETCX1KJYTL
Tt2yuIfVVlxyHo+jgkzMTGUuW9CXcW2hlxvp7bOQ2Y5UncogY0IrENwbfyJNMw6J
E9bJhKU49BqEWvD9ifl5Xw==
`protect END_PROTECTED
