`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AL4BRhJaC2Er+T3JI3l9nAl6Pq5HsfGaqRhe2fbC5NNQUTQDx0Rzc7vy5oMKGnXA
AMOpP8O1S1hv5avXZe0j2K0Vs9z5I5y3m2kUz5XlHqiWO18t+IVFk8UUt4SMLE1e
zvsF8tenKlTqW3FKIcWlUYDNXxtN/nafLdG5YsyswYlowH1gRzUl2pI+laV9VfAl
NuDdTctxeQnFbIKl/3Matq+83lv4Ohg0f6lqvRYLoIpV93L8a+8WsfJFlmtQ32r7
N2uOfsT9ROzPEyDQVarmBTHAt8sMzVrfC+DlPqmq8UtudK9o5uHm0MfQJUwSpLnw
`protect END_PROTECTED
