`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eSabUEHCAIvJW37F4Ojvh1SFj7ACD3A7Y7M7ujBdk1WAoo9HAJs4L7lFI2reT3IH
qcmw8iGGcEupsXYcs8U/vf3/IGx2+wBanDXisgj2TSflkxF89qD9SCiVvdBccnha
nNFoEYfYMjvSiSuxqMtQU0uKsuNwSqZJJy/d8qTukLzUJ/fMhDZaLyEQFfTsWIsW
UnIDS+JiokJB9xsJc7H1Fb8rhYcXSkpPhTD+p6jqnbZKWvlHrb2o+HPnalbbrp6R
8brbWbrvFUTH+iD1/wrws6sVkWVROJNswNE+fuTP6dpjM6JBRv67zrTpfWzbX7W+
ctkBpRD26zRfk+JoglPTNnNXRC3PE0NxJoW4f7Ozw8JgmGmxM36Hg7wuzHSQlLbN
cqZua8S6oRGMD167a5uR4g==
`protect END_PROTECTED
