`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYyzIf+zmv5fbcmLcTs2Xv+Y92RaEJMDguI83jemeQ8Yl0Seu5OKNk0XG3AdVmZg
NG9+vYz6tdtITuBzxxt2b45SohZlYmwNfYuIjBymNEUklqjxF0Qq5EB0gHJ1WEeB
/ReEVa2tt7sn4ExGVPJR0/eo8CMNTooUzLh2r0X9zSm0xV/8HA8S641Zmf0wU+Ik
UGQCKDQdb1bL9y0MCuUyPdIctBILQ/I0hY7kaTt5hcYTZvuEKQn5tUe+Wbl3+sxb
AecyVt60E9yWJZuvetfJzcH1E2dNC2eobzPIGBRxyK1AQXk62z3kPdWAPlYryg/d
ypTAvk+HD7HWhs2j9qeacOQEg9F2ADcugGRUKUkrt04nikdnveT/yBLF75Sahhw1
exQf93nu6xSq0KLQzA1BcksmNX3//OMcm6aMrB7/nYG4uwOjn54Jjqmw2U8wJPuP
dpOjF+wNPcoawJlNmR1gf1QI6kLGqaAhPPMsY5SqlKdhSd0wJwngyG+m96kLZNWg
XZnfpMX2dwEfuWZbd8ueOQ1PVDR2bDMRIFiv9/O7KXhRCjjfoHKYRxdLWcw7SWjX
AW99Hk7AB2Nsz2fB1+6BBzqkKOUHV7QFujSf2pk+F8JPMZmM8vx7EF7gw4T/kwus
/F0hgu9E6/Xujk6L+dMnYc/jgaRbhRdC8Fxvl5pwkZyons6qHX/IbhurEfk8m287
13u4iUW5T62fA3WJalPvihdR5DydDmaXbProvilIeFLEIBazBedoiNSFznPXcHVX
ACdapinTfyi785Oo1au5CBrU9yZbGLRVmGLBkc1HagoS5Yt0uFCPsHvLZEP0yqwg
yTQAKNgxPmf597hy4Vpwmsu7bAOFh+SJX2PHp+w1kb2yHCCPQA88OJ7x1xgVM1Xt
Acqra8ah1h+71zEUj1wsHz1wukPHefS/0M3wkWINBvLaymFyqnkRc7F1MxU87pRx
qQlZmc8NET8mEQ6RhOHLNPN6Xfd7tOz2W00nkkpcGLuiFIINumQpsjTrXFbjpb+W
EU723hIE7YQmHWs2id0nkHQ3RDxGUwxcmzCAOQ4SQAt38iji7IDNLGql3CMNmhWN
3Eg3g8WL6ExdFRvld/i8RpMwDi7na7Cks6pru1q5m0pp6Os2wQvOy6QG4+t5xTzo
xdNMTQmgFYLIpnJIwHQF9WlsuOx3VxqxDxSDmvSbLa5hhvOZgG5K1Iw81BKHtJei
wo+c+62AgkaBKrXAa8qTsJtIkz2uzbyv5KQBdI1yo7E51pSfi1qVYAxiEM0ymooe
/Z8mH987AeqIHkDV8InBdg==
`protect END_PROTECTED
