`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n0n9ENOjsO6qrI3DH8emQLZtg1YWj3HibRmlIDUXrVDL/Y0o2Dzz1xw9zVvCUHst
zQdxXcimhUv2MySjUlTY/pVxTbA2YaLz/UhAzVwVmMcO6fHC3b7qZm69hKhkqJW1
O+1TwuWGMtcHlp0j2nb4BKbVxgQuaApmZtTO8Pvz8aU7rHHn4xzZcp+eVhYlF9th
nz617TP042IWKSDycvEsi//m3Gmnlcer86frftlAc+TLy2pQ7QqwW5vbiZ/ilU23
AuC6b6oT6VCxhFDrvv97yUszLx+Wnb5OjBLugKQxSPvDy0XYeI7UiHIgpxx6xFjC
14ICKOcaeubUVXG/TWe9BYjZ0flpj+hpCGCHpeKIsk8WTJ9vy4dRGmMaSdqR1ese
oMPu60ITql2cR7yV+YVw36IW2YYWqr0Pfg3KbfRi/q3eMeK7L2ctPvdC1i40h3fp
cuhvd10F/UYe54ApIMQJznR9/xmY97UMOxonQgYPAw4Mwt0aEBHg5Fyg6yih+Q/5
t0GEwPqIDoJAoF7Z+d2XxOU8edmtPvpSeyHeKzvvAK5YF40Y/QUssp2NktQQXcKq
YfcqB7sPlrQhXrKRlkZCt9GmsMBfVF9h+MlmuzDTYBnubEV/wVUImRzjEnH+q7Nv
BkZRB98GqukiKxC7vj3HZvtLwBio9ZmVA3Yogte2joGg4PYSou3v4Opz5plN5qej
w9KGck/3wYNlR6NM+YHKginRKk6sXDoE6+TG3EhSRuGNLzekuFwVlPX9p+0jdaWe
xgZnFUSQdkMxYpJLgUxkMxQY4iXueW//cAf1A9cQb5vSEkh+zh0RaYH08+vq9ak/
MMBEpENTWVi+qCS0f9LUAMBCqtqaBwdyfdlGi+XmNbzJmQ7nchwCtBQYdC5NxPnB
tMfBxYcYWy0hJNMl/TKu9fghI+/zAbiR55shoFEYZ7oTZH5Adg5aLHE6luPl4jaN
JoXdi1WnQyzvgCCyYZvRqIg2ciyzHiSqSVy/Ha7xcIN00gh70X79T+Gxme0ORUTe
65jOtNQt/Ax17j0ixU6TdW7RGn3V5qcO96YlGCcSc/BksEZ2lT8Kt4sqHCeQsUjP
QPYRt4sxpXhn1L/ozc2Xmm+oWI0XwLU9G8gq7qnszNpZCaq19oseeqYVXU5X80Vb
joISMJKi+0w5seX19L51kXPlsfVBcZT2GJv9BIfXqj0/xwLHjOQTKc82tBjLLkCl
/YQJjzOV+/FsrKdnXNwD6LZMYUJuENRTrCymH2LtsWR0JVMRjfQzJcOGnFTHMb6c
Ug8NCurscpfsTFn7G92yxr7hRX9Acvq/SUGd+JZmcfHFMm0fZqIrJcuHNkJ/ugwI
naNyCBX0bGeuh+0Jvrpp+UlKHyg9o1C4V24f/LB9XgfrXKQobqdUmeuspC32S9Bn
hwBqbf13Xds/AC/6Lg/YtFG7aRJ9c0nW8Ukf73BDOZBDfhZGHUItBx4OqSlVWi3v
IkQ84BET7yy/Lbukezd2JaLQDYOGG92N2fWkGtdt9XlGqHytc46e3jeTX3Vxb6eg
nA1KCbq7itvNZBhuGU0fKL7qPQ5iHqivs3OJhRgF94cqcKSd8PR8hV5LtpzsZKeN
dcEuaKp7msaLLzgzzg8ffMcy3Ljv9PbAMvV4/C94x0GWD2l22MR5XlmK6T2x0vYm
qgAOh5nDYN5R9JRqBF7diL2KpDN+6y0L2VPXpfXi5YDJg6dJ047fwj3/mKOyqAUn
BBu/XwbHYE0MNtlG2uwk9Bc+FbCheV2FsVNEAQbSuEvq3cG1+adH/CZ6RJgt48N+
1OHLUF2+qFPCFRi1odHOkTDj9uZHZuvRaZDSFHeb/om2vvXcKKacVQhAjWwNcoUZ
BPoTf8c1Kdiov4Nm7GaypnbT5OkIOf+Pc4U36p3QFeOR1bb4KNT6acWH7rIj8mRV
ICnhVwK3DRsJsK8fYQE8hwXED3j0jhtiXgH4DerFHKkfebJT7QdLbyVo6x0WdICZ
Z0idxKoOw04zYgaXeFz+vg==
`protect END_PROTECTED
