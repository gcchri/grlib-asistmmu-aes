`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HQvTONTaGvfk+fQBNQnqr2zbnUUmKJ8vRgyoydBJN/mACrZbEyeShJJUwoYLnvCL
GF33Y+5w7A3wAowGLNXaj5r0htFDkJEVbHmSH0bMJzdbGzHT4+/a6w/1g7Q9U4sw
R0r392ekctrC228Czt3h6tzAH6ZUyRSiGYtzXIrHDbgAAIOdUWP9hN0j5eWV4tlU
ctZpFRX+jdrmLB2gz3FboFOh8alIJOVL0epxDZ174Kg1wDyBOQxofJ8COQXgW5h+
VrlhQYj3xOne70SlSNFQ7MBKXIeyjIM4xS4FVD6ZfP5XN6v0DpFYh0MwJVdG9RX5
VAuHkPC8crUNEU6hgkJEUUEq6zav9Dy880EiLWUmNyHBF3t7BI6Q9PK83XsRJLaG
GbCEQSB0nVDM7zYyvcxWPUn2dInzNotLbbbaH275eBI0fgwjh2pmkze46dK5RHO8
62uNKKXhKP6P/H7eH696KcnUmNQTitmWvix1Q+1swilPnquOYEo17VwHHXvjL1aW
CIzqpbpeUHoYOW/IuUWOaBVfbM+CjwJFc+b/0E+B7hJb4P7YhIUobTAaNaOplr2t
`protect END_PROTECTED
