`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J5Y0gEPlTmFmQ7lZYBQRhMtUrXDZ+oK5CLLsiAWWnvdrN+H39SgEoWQBj3X7GGcg
274uWl74IaCMVNbkCZNZXoDkowAN6FI08qmOJmajwyC/x0SU4FF6DjYBuIELTYsu
Zl0qm6s4NrBzXe/uJtpF6iGY1mnqV2yTRwiw8JX3EebDXGrCzAq+8jOgdk+AH3wB
22PvU9ywTuWJJ3vp2JwiP7r/+oRIb7syXTsxPPt7UqiXIhE+dhKFDk9Qc8RhccUU
x5fsH/NE3542MXmFCAB87TkOU3dg0yKtvZHfLd0bj88A6t4tDe88k6LXphHXD7mp
YdHwUMUO9yx/dQ4N+b4CBGXhfQZVUp6rhs4PkOHYvbGwFp6N6SxwAqAB1OoDD5UY
D+l132FJJtCa6/vNnLmVD3Syg4o8Q72F1oXrC1t7AHw=
`protect END_PROTECTED
