`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z3SptlfXAkAy4wbIf/ZwvlaCjn8Abe1veqYpnlaeOw8zNZhI0cYJLiFetQx5GsAI
7U7OUmg4XiZTlGpGuKU5dNGrQ80E7K0l/wJfA3KprZLEbzN6lj5wDgOMXouipRCe
37fQscFoyJf5vj0UIlKFE2plK6vuA6Vi50vvC1BOZh1DvPtjxJL6qRYEd3sJRP0V
mqpUrjyGoGIQUq0dRlhEeSdUDy/6h+c0SPTbTN7Mt+TZ1ZIYhuIKYqZkesw0fO6N
8dVuIt1TL7J0r0PyvZtVqQg0R88c7uuVUNFVTGV9L6csw4NRtTsMJrLimP4lin2/
Jp1K4uAKD0vom7u4J+yBm1UFOvOL1pkWvK1Y4Zpf5Z0=
`protect END_PROTECTED
