`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cpn/qpQvMOYZwP+mbpJDbfybquaDrUvV6kOE0TpWfW/qIaaqOoPUk77xdUZaUWcM
fvp+HXglWNRwa1kgE3WB2yqvxKgTT2IvlrnYmpmKA7g6aUvUk4nYphCLAsu0ADqm
MVdlJvu6GLpo7Djx1l6NwCETvPePVtrtTAOWsQjlmL2R6tgrjP9To1NM3wNuU2wj
fMcVPFLYNkiUpuayhuODAzNoheLGCU0K/5fTE6rabn2NkS2RXVY1zmxb/ps4xBGN
8iZJlqEMQ7KMPXtbX2TSK9gAnizWO6YfVxvqVk8fKxPm3h0Bso/zUnYZiS5DkDGV
O2CgNlyNPD2TSku6cnU9pyy/mH0AFoROXG/0DJnbIPOI16QvRTvHBergfZ8qDlZ+
vXOFfmGnXsrzx5yjoxg4Sxlnir9p2Gnc0/hEDOVuQiQ5bAwLa620ty9mO0LRnj4z
fmcexkU4IddQ+J5ysE3tixsfCmCYlSqez46N2usXbub1n+x5nNdHsLqxrOhbsfl4
iqU8TGrD14JvrSjO0GzjILp1rSS60IW86k1cNBNbJN+f/KbFliX0YYDva8CJZ+Zm
zm7gwKE4TTgODl5yf1nYjRIxVQcAqwqGoG657dlwDJdQB6zP7bSJf0pH3z4rf3rh
Fp/E91BnbSM0rM6CfiDp7Q==
`protect END_PROTECTED
