`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1dmDoKvY2zx8PR8w6WOXAEsrqNDlmF4wpvxIsMEZMWAvUQclKq13GQ0z3ui1KRO
D66CJ/D9CnkKEtagn9l3kd/kMgunIbA1579wfa8QjIuABfaKLllNhlExGNA6SfO9
DY8RQjmHn7mRgeYFCMfcPSp7YUI593KN4UQNfZ0zgg8xMgbEKrJ9Wc5Fqp4LuHz3
HuJaycTeRKAfjlj1U6b6hhp0jVHzSleMT7DobT3lQOK8aCEVdYAFl6oFKyP4NZgM
aKBiidvFuaxa386PdIf2lFrdNVDVaezW3BXbK4+BfDyaNOhN/BpX2Ne3idEl+Pxb
AezdCGVvspQ4CaH4O7xNlsvgDmKHuE8fEUexPxD88yC3vAySCbE1Z1VHcYVZc91g
rhZgi/EkNQmN5sPyV2UONw==
`protect END_PROTECTED
