`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Btil9fXxl/7VQNXf2wBf70OCS+gq7XqsZpVzuLPNmaHAGzK9F3nXyvl+JQl+8vBn
j/whWaB2pN9/qQyQyEy3VgQnaQLYuKuu0ZXjl+xacYwP+8raJIgzaY/VGcKPyrFK
rxJRPx6zmgfayXa/FZ1i43vSrNsoTtK4RxtHQ41VAtPN8Zzgsgep3P8rMfWV2KK5
44hmd5G1J5Lmdv/mSCrkVyLgeBIp28Fy/C0PO2xW/4Q+8knvl4j2/YpCclOMIMtQ
CURY0r44jNvl48U/dlbUvLpFnZZw9FpZHzuYPgFAg7JUWGyV1gLOr43d7kQiahHq
0pHnbNyOUa+P0T+wkg0p6qmNwkdYVnogi40waPJ2JmR8ta5Tu7jrJCSPtyt/qpep
Ui7yLWAr0qwNHNrQGAq7MPpOqluacca+kr1yKzq5Z3KiXd7H2BeuupjAhbpZcHT0
AAI8YJLVHKeEJYErt9Wluk7oL7Uq4xefserAyW/QrkILHZbtThQBsByciegp9q+k
HzU0t7xIJyus8qqyq/+8djpsnEm86KMd2BjkUtB4zPnvWQr+i/FPdVg32lNEjsrl
UP7wuS6vsYEuv/wC9eRKTkaTGM9rEeDIH94mSD0bNJs0IAqZl5/pOEDF8tOKgksC
27R1OyhfHKDJCU+/shLW0PJuxTKscRpF+/Gl7ZXwCd1omC+mv1PTi97hUJHh9sjF
PR4ubjHgO6uDZ+2CUUTlgNKULa0m4bZmSUrQR8OtmwyKdI9Yagn9nyC5PuduiNQ6
rcH6pI7e2P+D0vC+WOHPvpLicoL1kyuCY2j1WCJDyqMeJs7IAXO8zyEfvUlpj+lu
mIPouJ0Kp7NhyAhLJuBkKlfNUSw6dj5mzTdrYDwiQGE=
`protect END_PROTECTED
