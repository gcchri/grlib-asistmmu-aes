`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XnPlo0F9KPblUhVGbksUeRExn6UjKkwx3jKMqXyOVZd1NyEmPRoFLRhPDgm8v+bH
mo8QMfHSiEECOb7nnWqB9dsyeimyocxuAig+LJELEfvRVcBvijuUfIJ+Dw59LVpy
dTT4Bit/EsJMnN1lCyRDhR53L3X/JfX2EegxenGb4WSaUymqBapxJG8JaYk/vyWb
NC8WO414wHwvRMjnAf7i+mmPu9BV2GoQ2d9ytKokHbTM4r3XNUrJrS53u9xv7xfZ
zDC2jqmn6khZJl5W7/26wvAfFL8kFhBMjz8hW+m+H7k4oC3ug9lBfmmQ3+9aehrM
VPu4+uxcRehyahJpLG+buRarp0GQYZEREDzANcoY5f1ytpbXLS7Gn7JQC5Onm/gb
MDOhRDczjfm7b9gCj4PNpfh7jl4IZnZMMKZS86supmClrAhFG0QLLZ6UX5xrOAnb
K6Ypuz0pmDSlqpxI3LgsdQToZBhJV7bRlz1gAOwXzyoXILapr64XU7xaIPZ+6DJ1
hZL2ZmAHf/ozTnzBD6aAA5F+WJcbqAKXlJMtHvKRM4QGWuaidcI5Hh9xVXV1vQh2
x7ZgSpiG5JSJNck/ulr+gEi8iN3FJcpVmupWjBVeWjeYuqkGmyW4O3OpFrQNQoGn
xvJFGWH7OjHc53UGWuoNaXNA6gqwd6QRmXiWXpA7FRvoiwjzYC36hdEnrZpgZ4aR
E/YdnJdhgInr8pFY2PIAe7ef9UBzv9sNaAyscZZZF6WsLoAKz1hFqObwyoQ8GCv1
dA1gcDKO8nUWn4QuROo1sGB2l4S92vx18XW8js+Gdo7xhKywBwqwPKoLzlxAkyFJ
CtyMJ+bjw4O6UF9XbwJfoKOjfr/D70aLKLtv2/2Is/CgijElIdWyF2ksCPtZYS5M
1GAbgFnALhGHdzgy/STJuTnV2IW8N4z1GCbRfLM8787rfo+DtyQtvqiGT2hQnPZ3
g+B9cKi0ZNvovY0ptBi9RYv7DApiUWKgJEVrC7cSn4vfB5bORvkZyTNQtrrZkhqQ
PeV09LZUyWg5qYTGtydTeA5eyi5t37zjSF5rc8stKxGJMm0sZOEVBjbPpTYjVO1T
/DqbN/EcWAGSeAfFEMdtI4UxhNWf7kC+sgAoy3nheor/+m81h3QrLY33K0Q633tJ
VMUMWHrpIIGFRnSnr4gv32HR9l851on1sKxTz+M53cME5prOvbZ8q3XBQwpguxX7
igX058qRg8eA3D49wLLLWyZx13yvZ88irnpibb9Ae4kfrUJ50W0YISw8BmUTeane
v7g8y7F4tLUwtfKpiKO1PB1wahJXH3vq5+7agSKMyhYtBXdOLlJwZucFv6ajnSJp
ol6nkupLztTmrTOJbJi5pe39ezMNuahAyMEbnsLCNkZ8DAg1GzfOnAJRdR0YXgPs
l7YdLqoPs3Rfeb61strk1PTF+W92WMrnCHg9XXa3j4Vf0+3nr3Nu7SA5NXqneTWf
HdDPWBGqafwXc938I2tVFEEjKg25wSTpEqGRK27o7/Ts/03P1U21l6T36BwtE8UK
dalJ5vEer/kMu3StPhly7tDzwxtmpYynmI2KRMA3NlCEUy0+RGpDxhA4CswanTjL
fHPpGPy1vzS9jhWThNZfIAh4YTsvNCxuOvsdMIK1VXNSnKaHi2DYdMBVTL8IR1qm
w/h5dBsmmUfkeNsu7pRopZg9/7nM3ohA5zL8fPNbE7ux37j3oZzuvDNnQCNVMjHF
huXrzADGpEe114thqU4cuTrZUyKYfrXvPuDHwTcVREpWym5IHM2ww42KJ9o4T0Cd
pG/elJTTSxVFRgdt7gy/iRrkjyA+aRhe3rWk567PohlHK4p9sA1m18jTYR98/22y
hcsIF3iYQieNfLH0IZdtIFw14zPkrPVfNdHhFe9VecRP3EyhwAupN5/tqAaBQ7yH
MmTQ0PZql4iWNOLDTLJWBg2XGM54SaPGqsMYwZs8LBxOJ17lGlUQqFsUSd56u+s4
k7/zgxCVV6GXC5T4frbXNLSS3KhmeYGAv2yL7IVZpSCCbzp3SdI3LfuRwkW5S4mS
zAoevO1yIMCDXztKU2MgX3c/NdGQQzYrIiaGSotBu7WIzAmdTGKHj+zLXUetLtmh
/IfUrh4heYXhFEnIBMk9WIEaN/iy2PixKxIHyv7YA9q2ipDy95zRHz/QSAtddND5
+cieb1l+zvyVqoCVWZdzOwgQaJKvUXJAu2n0CpIXZmnx/pIxvOt5tVT/kFCzpUcb
9C6/NYCdiBvEcD54SWbNPovMnV8HXZxxak7Uncm0hvwLx5Hn7z+B+fbh6lXtF00v
dn37zbmQERTh/7OQYUxi3P6HI1Ahlso/3s3ZrzPqpC8n6wpcREtssHWDudG8VmLH
HJB2HdWL/F5xm5ULLZU5IJISEFPusctIyCS3UEHRroj6YlPDbQGx4LWikhiRJ+Z6
K79sS6HpufR0wHU0mqADUpjpG9f5vNcmwYNGwGvtF6wmLSUoPviYYWD8umMj4riE
PRrZcB8TjBR5U8GyHOlqBCRyPJATEUacemVR2O1ChLT8vfhHiIYoiCIaUonMGHa1
cNCpWjDNgOeS4OMVJKJnKvTKDMozIJZ3M0Iqcw+AenwOsleO7bIllaXZCL6KqHvx
UNxUPhETPHq4ZbDfAtVytl92lvgZvZVfSVRw+44W7KteaKYb+iEsxAxjD459g2Km
nWHbNlmJO4iVDB5gPQ2vsK1wIgirz94xzl6TqS+5FAaxIcRKXCQIVqc2h44TTvbX
d0et264iU4FMVpglXyR2MGobJ5euqLhPgsj9Wav1Us+oudIN3cJseFg7H9ZWiNsR
wvoirRwFsj6Xogfo32v87skW+gw19t/p5feFYiS4GQZlCB+RQPTrOwls4mlQOjl9
wSCbuJQI0Ul7nLMQi/lmmT5oYSpcxF/QrjlkxjzxT10LTcxf2moGLLaUGE//im/G
LP84f5pxbDp/GDQEraP8j2HK2xbnpV1rUUnneFnTlfGg3e4TTvHoz5BPop1R3pC5
Zd/htgnnGTxGnnO9g4T3b2X4OcBlmJevIWUmg2/jLUr9WIYBm14hS+3gwl2SREcJ
8+pcJJYTlN5f3recNUiVY/+0yszvKKYZZXur4hTrdHmS6UjB0p9BFqfd4hdBf+Du
0HYhle07io74b1q8kuaVthYyWOpf3Mm7Hs7tBSxq3OENOlB9CKlul+WedBqvpy4q
13idhqLnPAo7048Q6Tw4P9vkXFO5ptEyM6hMOtExDHx7Smj16zSS4a1OvLe/92vf
stQtVpOCqf2I/1DwykZPhhRFqi38d6qz3wbmr62thMQtquXOgs0tgb5JJUIMIjuK
yibOonAwDc/oJbKeYfPR+jZAT5yKeOSkR4rX1nqy0/Aor2sa+MX2LnYHQUQXYqbt
MhCdUUeFcMgMM00XW7ZkyE0hlLWQJBDBbpTNi0nwQPHq2hesOJzHNr+qNV45fhx0
JOjdZwnoUBdEEjXO8t3F2JMWBvetVRVlV4KEggKxsT1Heccft2sw7dk6/A0/+Afr
sBYIMlvdxgL7syDfus2OBohoPAh2vxfHllZEegXeQ/W1pXVLXtFN/+kv2KiYiH0/
0y8ABq10JrigseITDjcK1JWkbIFWBg8N5GnINnTLAzqsT4FkoOVhvHAdHeNcjMXk
PwWqmThDHcBoI1FeVtQKZu5QOjxSQfcaUSrIv5W1DOxf4jIIH3YZB7iNHcUAWlVd
4+qf78ZASwVYNdNInXsZx8AaGn8c5UMZN6OBw7g7rT5wEvgaP3RblG3of4RauqpY
yIY2OuDGqsELTtn0gcOy22W/gF2KITHqxVSEGFxxEBHm4CE5ULSVBLFEFetysIG8
IhFIXv/DCiwK93LbVDcaFa6NJ8tXRDfz/ejOGMhUWACakev98H+++Tw0GuJHPEnw
ESw1bEuADku6bFfvNXZLFoaRQ9gK443OXDC0+2XAhfUxeMyujDfoE8XbBBauXTJp
XN4APggc0tBJIKdf8PuzzVrIBkT++P44mfjYEGckrNFi0cDVGH2wdxmakeatk9im
orYHEAXItbm/2cTxYwY1X56W0MJGfj4A29n/JwwbfJSZIWxxzhE25mKRs6p5m7vB
otzCIkjHMV2T+ueWax4XZTMUSg5OC8TeVHyMNfdGUX6FJC474LfgoRetIfWyYg9L
O7MFg8oTJ/XJyu2kUryUFaEoPep8Q1cQt/2iaodKKDii8QDCUCalal1VznydbJBU
2tom9JFnVz4I9lv+IUofB23/r245YSvktMbFSLiVrQIRxMfesPQICNB4ni3aoqPN
f3gLsFUT7438PFikTZoRH9ydlWaLQu2sAGyqU7ng8mQNHdwZbNCiBb7o06tXFr5S
QKS74Akca257Wjv4CbWgS3Lv/4Fkul4mHNjGu8+Q6OSDRXGcd07KECu6g2gfl7wa
3Rskd8PDdhg/SO6w/B73dGiALEBnQbJHpVZAv9Bw5Moe2QZCDZKnFAFS4KfGwauj
hdD0DiCQHfN3GLx0j6aC9HEObWESgdMOKJRL0pUeRY/wmQPSebtzAy4bvRY38GPr
VI2sJw9UHKLCsHL28bAr63ZDGasW6b+YIK43zcSM9eVOBevBxEIbCuRlcApfG+CF
ckGpYHdVdFMIy2w0L9VjfyvPPcpeupHJ0MK1MY7bHH1ZmWLXUcQ28wWxPL4svuLt
HGci3W6AS4EiT9rjXJAuo3bgM5gPQUD+7xJUjR9YNeTVlKbpjpUbAEwzX6EZxho6
HCo5o8p1Q3WyQijl6ywyNiM44J+CnXsU4HjiS2S97oJG3ZCCVwhrPJbaF92KO3Fy
XrVCsfbspyNWC3OcMrc20iTLMiPQLQqN7LskFd4bDJSRojJ5l7oQ+ARq7/TrsIa/
n7rYp7FVGaQK7DvfR6kDJiIw93jT6wJ8xhtseDMcTchHaZhj1OmWYphQODlPwRti
y5GqCBASmBdy2VsZ/z9FAUnNGt8ArZM66dbf+1zJ1F8fTE1VqkRVm9k23zG54eDP
4n9zljNAqXoDUyECg4xwZEHiWHPNke+0AEeHR9wBb7NmvvkuWMfyjy2h5FMGG/ZZ
YCQxFb6xa0VqsWVzBfMafriH7uo6aww2jd+3hZCe/vD5LmIkiK3bkUZCcJMQvhqr
pDsq6abf43uJRGBO9qH5XBXhBKk0jlESnhN/bPftMy26donuOZJqb8i/Xla6UpOz
8l65nXzGP62wrX4huBJz98zS60uG2NChsxZhHPtrVeVZebezoeZSiqY2x5ud7oPw
F/gLNltFdTPeM7dOYQy+kjGMRIK3y2q0Vs/NAT8A2lS0oOSc4uxRInEpO1WBtCBN
x5OAY/dHZVYYPYR5VNdaU59xZ6AJ+UQC1JMZzpSX/4Uk9ByK71x6v8hZkUX/njAV
4KbdBnKpeh3yS6l2H+ZJbOJzEI5CnTbMUIP+OUjnO5dHXfPjNGurEYTMbeiHf64A
s/7E6KHdY5KKETasttLnEYB9+lHLqn1ABIWWdskWFQ+bkaVJsRWLInOJ6WJxAqz3
XEBKvl8J8eQL7H5AQQ47EP4RDhGbeBw1/2K6wZhHBbY=
`protect END_PROTECTED
