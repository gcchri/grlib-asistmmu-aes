`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaGKBWEBHHRUEv+pL9O6zL1i9aw3t9P66I5NTAEsdC/pRSfWTG3wZ9S6hR0WJ3KN
UOAn/Xo++b06QDKwDZ16Gx1drMUebHy0d4ZSG0w+9CElBVAa4D+AfLwaYHMlm2Zb
p/h9+PI3sbt8QJcvUURmh0T2ledg3TKO2HdJcAQqmMKk3wHNJOe6+l/gAqurjcri
dgQG3gs6+1ceafbus3zPg7AlYZcPiYULDddYCmxBmBdHTOJLSjLOE+RBLIDUWRhV
ki5LunTJsn/Jafjqnb/I+Z6kBfdhE60QwNWpHg5BFTJkoqacZ5iu/oOijLlWZBPQ
iYxAo4DsUs7xAEo/tKMiFg==
`protect END_PROTECTED
