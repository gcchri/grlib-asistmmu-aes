`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9uB6lKDFJG4FGi6v40NpThGYAlWzl/6KILpT2ql5rfzDuqhhnsy9mtpqNbNZBGqP
aArz1WmK606cPrmTsNPp2NizX9J+AuNJ8zfcStGXtDSljmoC3bQJv9tse1gaWBHX
pNzPqcfHJqZu9vC8nif+CweO83UiMNl6lEOsJFO/mvFlt8cABwYx8mMRUFiBaKWY
o95uCla9suF0lRDqwDP6T5Onicl5EOZ5uOEebXOqajQIqwoQvtDaje4rxPpDmuIJ
XlsnuM31xbnzCbzkC/AJj2nJMkywadDJ+oX++V81RSiSPKdnHkeO7LUsHQR9Mt9a
aps0bOE/4o073Zu3U+bG0yhVsjTlNE/pWfjHcFwp54SHOpl9GydqPc/65J5lITkl
cnYZD02bUGrU5b/hLauPHL2BUEOQ4ASoUvm8SL7GJ0LpvMcAPUr5RQhw0AdaNcT0
WxQaHAcP1PGiawHpD26PHGpUvSe9pB49y1297WAJg9YdpDXHI+eb2XlmaOlZb/Fc
fUZ1/IAcnjPxRhpG2sFtM6eG7FPyAvuSWSAIzhH167s=
`protect END_PROTECTED
