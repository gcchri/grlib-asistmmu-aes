`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHzxBtFO0HnLgmrTqVXhTy4oiS/QYiQFu3thMOli/RSwqYOCbkuSofNF1DmNolwz
YMDdM9GCXmNuZja/4WfOu8oWutQny006Nf/wQrL0wT5KAmgwQAdwN4b209bwkeC7
cCe9YhxAB8p5l7cgSg7TRzuRQnLKQh/MlbUmeA/Zo6XU4329zq3nRtN2hkkkZYX7
1tm0hSG6WASjKtOKW0zqYrJxX4E4xUUu/JqMfkon8RVHvxAdAsmMyX4NVNt7850K
KSRS60nCansj0yg2Zb9f6+7uxdWo7JN/o/434HmMRyfKAjwJAivh38jbNZc4AeId
gl24ggn0AIi51mf/4WSvaHlmWlgx4Ddxka3QXdon1chTBgO9X+m0Ntj7//no+9JZ
+yI9ZOMWAN5rtmOyIdVBVwwFQ6yn4A7M+zVQcAPzc1z0DXYOfwqJPpPnb7oN6dG3
8mnHw01bQWBnIouGLIr3UyDHlcE2k1GbRHQkYpIYAqojt4pFDGAxqSGkooPdG3/T
zFZIDhuxvrbsugfa1rSk0mDbAQnRuvwq0+DZmlZ00we15B5PfBDUawmWKjbmpVa4
`protect END_PROTECTED
