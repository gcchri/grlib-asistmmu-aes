`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAj4jMIaY7DuGtGphQrlq1IolJVUUgeqjlpKY2pI3m30Dtkr97PGJU3iLtG1FFN5
FAzB4qaQilJBCx3V4dS03NNpVN/WXUTrBxtDwd5o3KH2Hvf1TIsHpyvk7/Y5O/p1
wExQ0LKwlQABFBplGT/OSxe01p3ffAzcMG1zJ80D05Y1Fe0QL/1hMPL+ClfMIxUW
Psj7i3AZGUnzMLOT4j3+H5iPT1lVBUv2epUADaVQWcs22vlZHjzSCgzxytOS1+Bn
g5Sy35LWoYBbS3AHPzG/DYtSW3kGF8V74Eu26sKbqGjPgkrI25zg0eCfWOkRTxiG
`protect END_PROTECTED
