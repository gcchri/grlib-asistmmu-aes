`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wsS61hTSa4mzpmorV+lq7GpAKpHtZLRP61qY5HgaTSY8HTlLa6+elco7Qkc7sHR3
kqvc1/MLbhxyMhoLVV6fMjsx+mHA6JkLVIAzhPt94tA7wAHlHZh558Rt0EUhTH3g
u5xQXrTWQo4RqEQBUWvx0qvCo7AUDY4l/Dp/gVSIgz3ke1Zbd9fSSn1abEZblL7Z
oUfnH7HaeHOvPJv4WqpwAZrSZkjbXCA0AES1mySDdU1aI9XgcKRlXm85YmH4r6EC
HDGQRlbFc2IQyHxpnK+OPBnsdk9TrJw0Fn6MmaTA5+ufRV6SgZ5/MvzK5UcA9UNW
zlOYc7eO3HZpejoDBot7vcp/5L8co3kxUIAV0LjoWUtK7wbP9x+wBOCPOgOKm1aG
y3c01OmPREtdxXGX3bLlyCrhCYluKTCGKDWjOq1pEsC+ExAgComdndVfAolmTSeB
UEgMXYqjMnValTvT8Jd985kWXL0bZVCcNOveHaW5XDcLS6TutDIOAlGeAEsbtmzm
vNRc4YBoVl5XPl+LYDmfyf7s3TEGo1W3V6WRmnvDSVYp323fekoV+6iO3m73xPzb
2oNGpQJaAw1BhShDjdg/lRgTXntJF6LGI3HTL7JVfHcPMhSuE6B1OiU/7E03439/
9HbcoZsPscTpoTCdydcHIxRxlFJ4c88MheC9WJ5nAvs=
`protect END_PROTECTED
