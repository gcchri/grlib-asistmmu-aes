`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zz9yI8shg8GM2hRNrMMDt0AxfaJwtDqTLCIoA8srIKBaP6AOBnwx28srxnBaJAEO
QV2ZS7+ajnBKYdfLMWZklgAvWZbZ4m5iCQ0wI7IyXHfxOcpI1T7W5YiYrjmWTLJd
MrYYobptfrvsyEFRGVZARwMYZn0knYbMx2fMmZ3TsKJyBC08P9RxHtoiZEFOVybl
d6ooXH9Fslc2k6q2d6s2Nzn9f14dTqnRdJWmRsmxU2h0rbkYIaS2oLEqHhqmy6ga
RlmUTB5/70ppLHfkkn6JadDS81u8sSHcURMF2rqe+c+D6Kae7XTx1ZDaoXAyD+1Y
T1Niv5Ln+EqtLLslOiwjO2hzY86n8SIHZ/i0Os4yq1gYFYTZSKa1Na06C5s4sQ0n
2k5FSHVBGP64itS4zqQeKYrfjxIl/hIdhOFnKXhGv7aRNV5OLNmDBiNLExwtDq+V
cHQ8m+SsDthYQWWWEQrQv0b7JWg/kzHAaVQIRHyfchusoBz3/jcS54PPCiAnMIQ1
dLtX/ziP0G4VO7lF1Gz2S8dAC6DR47STPzLpQPC1vznHYZkvdrVRlfBzvIBeliq6
ZMvrOp7uCaOnIrAp7LCy/XfZRbhErXGNHEByUphD/cxXhpS17kWdEjXh9av6l+xi
YiDDFyHEZqEQzWjLUQjYyXgwnNjDS+Yla6D4R88Eye4FqIP7ewoa4VjKfApoarUR
+r8qjkRP3xYP8FJNmWhym6aagx44Z7W0p7rvZY6hsoiydzrQrBKrf0TJGoHSqWHI
bki/r3u4yDj/TEwlaCV2cQTJ+RWLzK92Xi5adrl3RWYSNTX0z6BF+7KPGpUNIzeQ
GOXweWKLRLhcQ/5r8MtWtULawVq+jlKMqzVeKGOfrJFFMgnFdNnfuvIBj6ZHWmzB
j6F49fsHpXTGzIAcaGDSPbyNGOjwoVReqK9ocUlcV8dAj2yIfoVyrRBWMngTQZe4
2yLWTsupF8cS42E4hU5eT2mSTRzsAl9JAEr7B7ildwB9UHdsx7QLCTF3QagWFZiZ
7Uq0wCv3Cnf80aLKKHC7hJDDh46plMskXLZZvkdmUwMt4ROksx1HK/b3YIont7r1
l9f7JpHRtPdsjJAJNgrVDEW5PwRfr6TwlSoxoVrU2wZ4e7tKIZTEpVFDwXlzeKzY
GSeGahxDly11BBt8oCjGcl+7mb2XdlrmNjG3M6WOirYZV0BC4lrLCWpI2tuN/4H1
9dwPkBvFTl6cxDBkV1//oWBE9FBwnCNO6glyywlpd/mM4KhpvBWV0fYLW4EO4WQ+
6d22nHIzzKTIxHqjHLxYKhq7bThOcHyl4i1PhMfJc0BPd4eROoIWM4oifAIeQryi
uVIFKm4i5KM6mwKzLJmYA4QXVFgrW3IH6JtBjHYTCD40ZRzx6WC08ODa3QvhOXov
mI/NsHR1lNKrqwDkSU3SgFUMdQSQKO/2dfGkMc+OE9ddC76hr+ufbqb+uWpfLnAV
dPxSukBO114u2wCIpb1xAhAw5hT+svQ4P7ORhVtPgXH0FIu++6UatCEgVfUsZXhP
2tfepR1H3ksV4bpcqPOOnCsTbyyaD051Q1fzsUHOfs2GjIIqnM76bEu5sIf/zBBG
vDeVbCHtWCGozVqRpTwZQBkUn8MJNteIcXViPnZ5GF+C+QiB7h2HjTwMDcj39/Hd
MJr67vmvXZaSExnnkD2+xpiUyG0oKsPeTfwWmAYnJmWECI1XZfQ0ZHckhgyErA3S
4qwL5F8waTM0D2qqxrfbWSttNBleDerebHFaRYMn94q/euifAy2JQS5XIPETQdgQ
mYuFGaxaDG2q1CqwjQ9zR5t+s64jainRJAwDrfzq3UqkWhBf/8juYi0azGi8aKx2
rVI4Vc7CxLjdAiEsL5LYjRclOmu4Oa9elcrcUVItOncEyDZUTtNhb9UKJuO/1K4i
zqPsxi82jG4AoUdIHIRraob2hNl0ViUwa0hNq0gWBpHwXIpjbY9H/Fcu2VuQKmI1
IkpHYRdXkt+ePWLzZ8QVb7Ra09gApM6ChGJ/jrxvICynBs9Ko8/Ni1aBVc++iZEM
wWLGRZkEfmcCPTYpQWGdVke69F0ut/Oe4epvAaOo04EJSf4bxqq3IBgzh17S5MVz
6l2LnIO86yBNi6JYz4EAWEv+uoB2A1hdH+29MNJtaZJF5N0LP2pc3rhnglJWD17T
/RPpCFLUzTDK1S96IMfGqZJEOyFIXrqsU+ChWnzKCIagaKJ50p2fpLI5Bxel1kir
QD7Ka1cl1oUUIOscpfu93WwEpo3W+BTzNHIWbm49wthfRyOExODVwwuxeNzL/fuQ
N05UcT0Y6ZWfGpqk4eSUN9LDjpBUfexig2ebNlZ9sfax/oZfQxeNzz8D5yoTcb0s
IbIP+CO84biIwmIHrhEoRk9K+NB9CWP3d+qTr+XBFRPt6vgy05YHoR850/64eMBR
oiqRF+s38/s8+g5T+bO2IdqgC7U3lc/6AiHtKWhZxwlAMeFgDgWfmumatGlJqFNx
pLndCcwJZRPXiA3pdxjYXUMSMAUNngE5tGd8FFSMIdrB26W+Neuwr2F+kdUkk908
w4ktMppgfrMNR/cqLLZDpt7TUkVyHDoMPqhA1D/OmC9dqHWXKGQ48EksjVSORRZr
94kHdSpgygabKiqaw27iC52j0cCcwW3hX+9lhRYY8iqVRgHf/rqZtLORD6YMl7Pk
bzGKPdptRdOGxNB+RriYgwqWLuAk3N2S41MZHkNFXIYKgJElk8TU3ty6hLEPcn2d
SPREAfy87rpPZAdP5T+95WsMXeW9sUaX/XbNXftRBkebDSnX7Xo8ECmoY61inXsX
AuETuTZ8fXUccKlTpNcQxa6OhqhxbK8RVE1+woJEtzTaCkV/Sl/kPv9S2ZxHByqV
hF2dtAogUxfsvy2f5fONwusZrdNPZhhksAoxnmqL8+aX9JcRyaU8BO9FGjmJAZKU
8RvmQMnRwpO8widMv37Xiey1SCLO+6CTUB8wLp7+Pc/XsTwR/aX84+JDZUC8hw5F
U+goGENJgZo5NTdqekDh7cepMHceSWzhBuCoIRPt7s5k5BqXGBytfBxAbwZLCsGc
WgQek3dm0o/adq0b3L329dFIxYGoHi63CJQWez4HRg4Eb0lsQTbQdodGk5Sge2VS
0QaP2CidiL34BIt6SLO319+VuzpiY+FM47EEelLZi4qJknhnjG57ybWbogITOGqg
64TNyZvR1XU3Ll91t6NRJQbIXPTI33DbJId3TtPakxRNbhJTzWyv6ZKm3F3R54C7
ICy8xNTGOD54uwtcXXwEP2tbvhE+wm+fqVS8SfcnyM3+hX2CDX9VZskN2R/CSOMr
1HrjuzpnhBDrCGwWDA6GP/MKgbkVklSuVzCmFSvOtiegr8HlqKmoMebehFxDaHGX
XRaxWQ5rTSZpVGuOoPYIWyC1ZR/OUywvgvbI3I/S1VgPPdNVclcRsGgGKlPYjVEq
szg392ZBjczgUkMzhdA+PGQBOWch/6NpMi822pBBi1vu58E7ISBj5L3nRZtjd5mF
48PtypUuQCDQCsL7jAlzZT0tfqCexJuqzph2OtN9+Uvf9OSur/qrn+JbA6UVx2su
TKq/UfJey6EgEaG7SSK7S7UM5RXrz60AslsZ441xeJG13fcQx1DGR5tnHP+/IAJo
xF+mzbAOQhygDSPDd/fwSkNtrpE48uyKA4rSurQx6paKyYopyi1wYzMrQK3MO8fQ
N2m/9kxsnwtXh+paB5K5uzfqo+BHX87+Gh3K3BRaFpNJbZV2gk7LGoK7AGC0wokh
ycTqXsjyW6v9RAvFBLQz2QsnZuFV8vEhrtlcazxaaJzzJDs+2IMMqFWGTNoC4r4Z
k07Tv3eX9HTtKm6zlqY6bW13Z8VKuVMMZhIKUg8DHHivxHKeE/9A1g6pm60lKClK
bVfZ7OSsmN1d59Qxp2/MUqUTHSnqb5jI8yqH0ccNLyl92RvC+Onfoy2mgZ2dYbUs
R0Dj/avsVJw6e1gZp9zNPH0Rkk29kn8kbBFg+5jry8ivaKZ53TDlAIdtZMA6vjSJ
f/KyncsiLmP+U66Qzk1VLL29+qPuNb/sJZqpRpSgDytHaR6rVDn/G0ePVqQWmGsU
wtmyGZ0SwO3vWsUKPUu9PhbKZm9ojzJZp3Jaz9uAJE2UECifNE816SmgQArdSPOk
C6s8KUxCxTGxaNnFC5ApwJV9RsH6ccbwEpv57nbbWAARp6vJ7m7P03FM6DUERBf3
69eLO6vlafsrmSwu+KGDHvSbAPTL57sRZHlvSSGQ2zGglmBytsG9EThXPbDvewug
nWXg56GvV9SBENMdByatT8vBryYtun7Re+Z82BcGBxGO406hf1R/xwPgaW5PMEFj
yzTgsWLfNXqnYvHf3SOgUT6bG6qy3BeRbEHfiO0ksUBEsp7ebZ0903HpMtaHZpM/
0pfo+PPVF8IOJ3knHQoulBD7WahJwjdWtqrFfZN7gXRt4mJNj6CreccaMa0mJuzb
niZXwYpOFq+y3dGlNApfqaA9BNDwrkyIPv/drtCgDiNOA99gnRETTPhVyf1oopac
MOWsZm58wMwCa7TAiYxwe6rI0bOJj+ol7jHyydJuhdAAQ90VUacITk+/MD9fxXy8
0T/VSkfZcwl4zzKD3GhbhIizUSFpG7MSrRkZnmVcqYy92rjHeUq6DJfaub8Vn1pN
+5dl7QDOrWb7FtZ2+T+ftTIpW/9SOG1KUlnqjFM55WskFMlLz7Wcvk4wENLkMUbg
ahmqFNzzsS8ihfov3arN5dtDxJLc9571NozhyqYddt6yIKRcIIUJtTl0oToHDrjX
utUVPVfnsoujl4RUfBPpxdHFjXWqdanhaU9+s15V02wc7Z6h3OaNP7Y43iVkjTFn
i1xaCudQvupSpx3jiFNE46CUS4Arn+8dfZhPv5z+QSqYYRum1D2ixZ7gtkdMlFhE
yl8yvniHgELjkwqW8e4jqclTKa5FiGVmTT14WK6foXb6MHmR9b/0BHo6KZDtHrEo
rO5GZxdLYDQJIh766AE5eFpuWf8ssR0REkcEHOKa9JLd+Eg0uy0QorAkLTxp2Oah
3ya9tJj68CTjVOr6Ws6Y4PI1k8+jb6ZkQk+CEpRk5lSiIKd2LJ04gl9yvxwgnrmm
5uLFnJQmwJwWhdcAWkwwhXPX+f5mCIvoRLdsnqKUCkQ4vyFijiRZMssnl8A9ZtJO
4MXx5rRs93NvzihKGGVQ1O2XstMz9GUdOvXA0HX3iUNxEdEQnKltqdCJCjANdY3G
0xRisZcv1sx/6wn4X/uNqEWsY7qG0brubxnNa1ndusWnT+6D0cEFoKaU9/NJcX4o
m9F/jaSiaic4r1zjXLV/nn3mbER8d/3jjMnkRPxH5fkBRxwwJ02lYpXkHA5n+VHg
gakniT/oxKzMLOC5ef2zUi/Yu9N+qM3nGpkDevhcmPFuL8x58bR4NAcXmZXJxaI6
A6IJf+2B4K8bHTt+/cNRrQrabQEVb1n9JSOOAzb5FyvpBu4TuSuorMIQz//YwNpC
1hKGl5r5uBEYz1bUd6IYCOL/Uu5FaYkK9CLfDuFBhJKxAkoGpnndLRmeJAxsntT6
xzXpNoOr8+I/7H8Hu5vGI7oS55alX+oeut/LSzDNGtHl4uNvpdFxsYGZKXOJQP7p
ClhR9FUQdx05zFMIpp2v/bLDzlj66/+7iMfCeXCQtvlRVUtm9fsNymKtf+zfrTeY
A5p1j2RBny3ajnLnqfid5/hndvnHqkKRWYm2FcbRV6q7qf9HSVAcEXZx4dY4S73u
FAhOC8meh7CjzfKOWo/FNbJqZy1Zg6+lTk2PhCRFGov+p6A2A6rdZCApZxKa3h/b
J5g1Qlw5dYUxeb6/Ac/ddn/n0GTn67plAHH5aYtRJg6VybyxIZVOjcEelfjF/038
CBqZ63IKbOhjjhN2VS2i3Kk8dAP4QMXMSZkiOEKw+RduD7i+/kf0LQYxDD9Y8iS4
0jdKKaRP7+4ER4ZJEPqPtgWJwlsaiG7jebpadpQYCRm8wQcL9Fm8MtFUZ9ElnH1r
pQLlvEDjGGzAn+dMr/S6qYX/dWKS5BUG+gi10BAXCQYg5G/Dh/+mq5Mg9M9q355h
n/Sj3KtsPV1l2PiH5FNCs2nO1xT0Rdo4X6sW1EJNaBmxblG5ywz7xLTCwuXcODSl
Gcf3QpS48C8k5BFmJwTHNKlidtjY5+froBp3lh3g5wQ0UAkEplCRsv/oedrE4K8W
6S7Act2/pIOryVKLUKQJaCOd931R67Df5vPG4xoD25BZjgRiMVU97y6W+yEg1twu
6br202OEmzo8HaU2lU59bTTijjOGEF4ou5aOOmibtPIq3nDeLkHkq9Br+wYR4ZWF
AAKL11viorztu6mXBfnzGtpryvW20qIXa83OmRIvKAJ0TpPD9N3AkGphawko9p33
2siEQbkvR4rSWXAj4Kp15x26ugcSWzg/qcRA1m3Mstiubpsy1tRYqZXBHSzA63nT
8PMIzDS01v7U5Ef2oBawiUyJKYXh9UIhGXkdfX1SFLM2alvDNh4gPhq5ZMOY40ug
fds9CfXXuSJAi40360JfrHo7sUU3YHu5idjpg/UjfhTFbjK1Fj3Cuydwc5vKcVZS
am4N3oLyq+RC8F3/bT+KrsvrQefchZ3ePNDODxSk7joNIpiG8JF3/3gP7bDYNLQH
r7izZT+u103XeeLqwE7N0oN351PLQ6PFxt2owOi7ZCgrtaZt7kZo2uEkQppzdzkI
10yg5bjOr6X+bJ0riZMqw7XBEucK/JYuH3SxmW2Tl4j7KdNcUG3cIM/DH9IIctKQ
0Jsa2jGHTPsfTkVAXxfI7K0Kb3y3rTPrNzQVCWvhUSrXIUBuN3jdjCFm4ClMc1Ts
RFAW8NbaKMdQoUa/WWkjntu1sWPBPWk3xGGnYs+mlJgVXtz5eJlku0jgEHmKD52f
vCM2mII2PJHabFUcxrcXF4lNG2gdVNvktiYR4j8TRsKpiJsr1Nh2XYIPw+tGdt+V
qn4Myu9xOBbq1o6tDwDQWAgHYip1GSZIlvhhpIPIJId6+auyhajhtvFrtQGccnHP
tq8ZNrkuAl4BYUMl0tJsre2s147usNC8SDQgP0KCnHvCzTnhFvu1KPM3b+SCIBmV
v4Ekm1R9Rtj7DLrpoP7mu9Oi4k8jeuiZaZeMgbuxNxVoRCJvPTptJi4H8RM8MmBN
BvbpbWrVGPr+8fusJIWfjEX4Aw6jS+qPJInJPHPONu1grasmoUVJooY3WiCa4O3k
DuVIo0VNbi1xeB3SH5mPG/CThH5ZmmSEcDnnvuiPJZUpQNdqEIlrGAbezKSM0wt9
payuAilMXbhW+b0sE2qup3s43BvAq4FvvWB0vEG/teOqDmxXY6w2GRMapQyHatlq
ewGXK7oANNUsHf77+m5TwZWC/TM29AP9xfMWX7nHZ+0+ADA26Eld2HIVI2aOp8SJ
oavh8KE3hY/1opY3+LN9ZhOXATLEY878rF3HegbKm/TpWlYUu8/MdaOCHEW480Af
ppNTjASeWcKQtiHQIOThVT3E46qQNgaGTuyMwZ7OAK2aHJCS1KzNInBlBjnnrg0v
8E2gvluNizf5KehXQ90xFJQh9tO1jzThQnjvXoPENQyMcHBJCE1qbW45I/+sPAZt
UmyeqYA0Y3ufIPlPM7E0XJiPxH1G7QRhzBxeKOBh24OPavFi3CwyLR0ArwBxC/t4
zVnaXy90OSPeslFp38XK9CzFVHgdOyFsIBQLbqxLG/NAGpnfOESQR2urRJf7JODt
QHULp1FDyy+j/DUGNZjvZi3BitQ+VrHupMSO5zXdvMYEfWoZnrw9iVHexjcuZVLN
j9YZCCyjUBFs1Q2s1SD/kRKTYMq5Zu8H+bMck6m47xryNSNUXuKS/8Nq9qvbPrhO
exFizB4mRI3aRZ/+lLTv11mcYDmeBxrR1OtjMeWFYQ0iMnfqtZuR0lLbk2oXEcEJ
Fq35qWJI5mWcCjThygra6z6iWR/LHoNdUf0ce8UpfWWzS/pVnymkX/CEaX+Nf9Hj
JEs1a3AvZWCcCd8ibaqvSWX4GShuIaI+LsIni2c3kKVSL/B99gBW+LkoOZ2SEIN/
cDVOJocvOn4hH6jzCcxThmcJCq1fLOmDCs36FWB9qtktp6U3aM/GeV5G540E6By4
O0+UfCjwOe1wNF6DJtaMEs2Vh0wR+A8YF4ZY8Iczt5tiXzlP/LbBG50IDiL5hNnh
XwEZ2DRuzJq6O2YyfgYfYIsO6Q2cBPCPHlEVeVi+UQmwOHfeXUM2t236xu5Fut68
UGbtyoatLCvtdBenXLn85x+UrDy1M2DhMJZZKsGmNLMxEUU3mEUXCdaVYOEzyhGS
Le4LBKmVW4rYYGySHut0rnCxK35S7cxnXl50+JKqamgYmxEhPU4dlGSiKvv72XjZ
7ymSSobUBKvgbYcMx7MedBms4MuNnbZsqdmVF/iUaIgTLyO0lX0bvJGYSBiWPTxo
ObfSGmJXsIsapzZzzxJfwKuvaalXRE3AlRkGqjD9+fPoquzbceUlzAb3MBRl7wQX
HDKzH/fOej6kHgZAGQK6ykeZQKQNsevXHHR6+Ju0Zg9XwS+sbilXB/o5WbtWj8E1
NqWfMeaMg54tMfJpdZFeMg6IAtzd6Pc8rjgrJiaLJWw15IaV0IkiJyDKfuqO6gyd
jo31vw77BmvbPyW3V61Ptq/mKBo7h9YD0U0XBqxlxkZ/wljO9ptgGW4zWN9q3hZu
DuQJDZGwoWn1/SsGfTdyerc07OB3n+FoRaNtb2X9au/OMuIIoNnQclm9aFBsjnBz
JHfc4odZJ+CygNPbKetoRk3PJIylCBnpEv9pcRVX/oWkBLto8qcJk7o5I1WG8krK
TKN96w5hD/fYghLQ6+p7x28ErEUMJ1ZE28+IwiAWJMrbMA8X5AZ1CrJvTijrSVbg
RP8LsxEANHiQR0HaN3iXEW03OUUFeggtL5oYy1bh5nP5GJo5DVy7/0SrEw3FeCc+
hHOE7BRk2X3iZfWR+cY6amySaiwdUQlTGqZ9dVPUBa6pnWPnFXzp2UUlsvrcU2Kt
dsFL3aP4VjVewIMZZ2u7evlt4CR5LE9WVqajsdQc9N9Bcal3Ido2eWTGF6MIUds0
vRBHY8C7xDGo1Ebc34O1uQOi5ImjXTKN6OYfYPxbGMTi6FSzuDQf5w2xD1B36RbI
XDfUcUdkC8iulkiI+miD7cj/w8y+qalgWlBXcb0rfxYv5Gwzut12Z2cgx7vV/gy4
w53BPnJrH0XfhX5ydCH8+IFMmMnqiv+X+XWR1fpy2cwbE47or+a2JxxtEz3nwNXU
bFkxSV4xfXAOVeybbCmu+CRLKL05jVceis5LhqAZaB/iU0xzXe069+QNkcJew6gv
DUOFAmBN9Bs86F6hjMiSd7EHeWTmJ+xjWdCk7A3xsg0ZLtBEIkjkA6amzVlCKIA0
erWBMyqmYz1h2WOkY7wV5pWT/N1ikoGzOG/vXQ0ihQDv7sgIZC84Y/HeGwb+9m4E
/6XEprT5m/jSEDZh7vRTRHDnoSIOHd9PGWMQ5tkyggtX1U8VaAUGSfzDEoCdPSPZ
qCYGlIDRito3UY+MKSclbbJFLU4+cyVLe7bYFI/OWzU2aZ+BxVPvCdBKDvU9NKWA
pCm/+i6D2CnsiwxHy+82UToRg05HzNxUjT8183SbQOqGn2Rx3AUCwnd7NBriOQyE
PVvOjL8DdNnR1UUrwmlFh4bzPZolwkQc+7zwdY+paGruxuSvCmPdMzw9tr5Dj6cv
x/oEShJORTiEqzKurTGE1l5t2Sh5fnNKvftfkQhg3jsTSo588nvSZoLW7z1ZKTM0
tdAxuz8Zna0TY3wwFJylZtKZ2qorPCRGU80oBG8HKcz/9iwc2fxqpDtpIEj/JNSK
evc4R8WrOPfi7NpQchDEz5se1CfjsPW8wzBdIaEyb871WkGLmnlRKxOx2ZguOSZb
gu5jnZciLVsbtTn+PQFPT6lmWRWV5EyQohMjgWuGv2w4Fy8fBbnfzFC0XhCuuxnM
07IK7t1gjQlFlhcKq0ouPQ==
`protect END_PROTECTED
