`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f0O3KXj4OYL681rozv1szP5VQmQp/naAodG3Pqn5fbGoqHeCUmB2gE8lu8+LjH9M
sf9IxXEtwU1bpxBBxa0X9x7EDiC+gQfTr5fcH6UroMM7zQCIpfCt38VoENXIBoY0
L54p3M8SCWQgoAoTNBlLO1W1+kajpGdSBsBMhTPsibzin9vI4kNE78Q+doe7PG3y
Bwt+VFnhURiP1Hbu2/rXhKd+ANTdTn7yTIosIhZ/ieTvFvKLMU/7qqizN8V2K1z6
GEe6aT+oF8kktNKE4ylF8/uC/coG9PVuGlNR2hSkKb6xIgV2TK8RiLrzdP2nI0Vg
nVVF4c+Kl5L6a75Us8nZZm37TwY5Aa58i9TCH6qRDj2M0ie2QS6bTTGCBY0sJPL4
Zai1TvrZmGC6H34T98nE2kkso3Cr0egei8uXQHtN2hyKJsP4g9y/0zs789nHg9qJ
sAt2+4zkwbU8MMN1WMamgPiqLqb7YgGSYwH2okPqL5PBJlt+bAw8crBdQyGZZraK
AKg2ArBjRZmK8vCWHZBNEJ+Q1k4FQfT4ZUd4z+TsvLHWqXB/7FvB29Ek0X8NWEef
YadwYoPa5kpYwql0+h/HShBe5UYrnZKNV594GYCBaj8ePMfofSYeGTujja3ZnzeY
k9FZ4h5Hu6gAzLkUx+v7e/gwdLo5QfkeRlyWCeYd+w+ja311PHH6CLL0xVs+sey3
wuda2/27KhA/sYzIicLM5tj7hhbTJPKApfCPu7DCFqJnGq56DFbNqHCbe55vjIqT
Y+WjyYVN5/4ZvY5kqIwN5KziE+8Q3y4OsDKo8yQdTvPB2Uh2mnbh5f7KwKsBNh24
Hbw4dgMeVh+rBhC53amsFfwF396H80bRG9tbwpJ00xup9XNE6VVpA/Z2tWQOssf0
SoWoFX3r7R5/v7zbvIY7L3/+G8MlljKdXqt4IBsfksaBzbNeEgEbjBAscUVv/8aX
kNeY/7YBpagV0APlT8SiFf8SumfWubApiP8rIMY8A3MJ9fyBo/CA4eCMxYSAm1dk
QhcdFXiNs7HjhQaMHWv5J6CiUVxUr3GWsQoFhUj4cry7hELdyxg10Tg71533fw+4
x7JDbnH/DuvFgndXhjoUgetJEZZS3xNXOnjTf3lhIefIgHNLC9v8p9Z14o8QV4KB
jU8t4iPg/GDubHw/VH3QasWBlDV0JnNbioPHdD14mqRZ3O+aG8IZjCisZJsPJVxL
CVXR+LCAkgkRWvvjprCUmwJLXBcI+8kiEnDbpcDGTASGb7eSwH8mAmtzi81WTrpc
OPCmhH/pR7ol+Smg364n2kS/FaFRlRPHYD1F6gzZKjrE500BN/kxh+vcB6WehdjU
8pwiYIsb2J/qCy/p/WKY2DwYto23NpPEg7UUQlfCToq1yVm1V1RwzJfJp5UP5aam
Bw1jb2VdDC9aOsughqgXaxb2ptibk1Qh846HcDXNq40jC8LOIaVcHHwh9WirEBUo
5+714SYX6AwDXZ73aqwqckC8WmDD8pLzcImbMz2+5vujoSFmiipabAlP/pf/4xyO
Rt8KoU/T5T33dzLf1/p2sQ3cEEtpSIvioWosojLR9m41TS8I92O14poKxymEzkhO
D9ET+vo+XqKbDTVss+oIBbDYZ7hjb06NqBpE70Fiu5NMQcyejNwveny+Y6AO4ETw
vcMbafnnoT2tBQcsqjBzgFgezUcy+6fCHYjcd3Itkw6708OxxmOQUiqoY2dMkoQR
WWg3osadbo9SMqEX2Xk0IW/Mn489KxTLXryh8NIA61xgA02bku8Hg8z43MYJWslQ
Orv9mo3LY1+fyr1cBYrTBx+6SFIdDusIccY0kiBw7m7NdswiNjmNU76kaWCnog5W
QQIfPpda6wdfVWZajYCvCA+IRug9A43d6efMGPrTCYhF0aCAo35q6Zq+gX8pcfjH
P3obXZZkiJFgr9kGtvjjoODswtiK4GvyxOcZmux21n3HzhZx4YOAJbYRSAnVG2p9
lYLfN+EY+YyK4D5zD1FYKHmXOo9gzHuCeIR0PNWW7KJXQlO3rU7saVWxHIVvjN56
brg4puKTYMbXbqGG2m7gnZabJ46A9qSeu1bL8X2a6/PbVbInWFucU8jUwAJqbsgU
X1qt8b2yQSaiARYSoa8x56g952vv7ifVJzbU8vYaeXNVA4Op2PSEEeV8uLnUSUNe
oOQ9C//dBUuu14vfjA9ioWlZ5Fk2Qr3q8EeCQkTOFnTqsPflRepx0y+W1fS9jgeE
`protect END_PROTECTED
