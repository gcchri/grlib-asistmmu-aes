`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lNLZfEtpmMU2CuWrTWGgwqjbx0Dh73xcAzWIAHF9skYmkbeadYYaA+OpoidW1mLr
FEjxgvlh6+/plsGlSJv3u3Bu0xb6oxUMsLai1RMlY7Za1FxxyQsITvLTi86RV09i
1/gDDy3H3Tcy6/B2pZFcFS/cRN6En6B4eKPpobGucezJJTr1lfo5F0zY2Sr28GrK
Ob65M11jWmonBaaphyn3Rl767yb75Jgu/ojPdCM/eZvHbXyecuP5Nej7lxEEQ/Zv
K3lYbk1fky4fOhYGV6D+B6AwYb9u68Ok/rYEcXa2sWDzJNH/Fwk2Kp8UWo1pyCF2
`protect END_PROTECTED
