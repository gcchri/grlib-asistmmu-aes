`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K7iy0nXKQJOXI6qh7Kw90zKepwijfGVBxK0dIvvOka2tLybI1rUJ8BogKAzj0LaG
c28hmIY3QwhrgLgE1LJTtHjkm9nk/eGTiCZxcbrTa5Y+IXq4ussCa32nBu+NgNKj
e+TUT4Le3bO7euXzNJJEmJeSs2aGxoeywTMMw+0t8SLJWfHHW1T6V1byNlZ6PIv0
gtz5PXeTIpR9Fl78Ocs37uGk6K1vBmxNkaoaOvrsSrZHkEyenGHeXC+3VsdkaQIi
oiFT5Xu90bveCoAEy6sHXkeB5fDejlUFGUbsUH7UpXYYPa/61xWf35dvN5vSVlUY
hfPwT9hZPxL5IqNoBFvVZjUmrU+4KgiTtqx2ipco6q0lvUn2NS2CLdzm4luMZDEG
+nZWB+8K7bfnkssNNbD62hNvS2KIjteEdVO7iirxbudsgSoYOqpigqxWiUDeMWrE
`protect END_PROTECTED
