`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NLI4hh3v/qgKM56DFx4KYEhdROaO9f7lGT+tkDwI8hQj2VSV5tQnUea8Wi95WJxp
jKSmXUfKHvv10T/YmcOh8Ngne97vnVW1XgIz2cnHLbOOs7FJl+pHuYsadi6Rd37z
fiFKaE/MHatT1H2EPHJ5ge/DVSdLz1V1kfIXfbMOfASoLhe188/RneJpzyxizB1W
6fm6FxLyEhheddYl3Ux2qP9lSaTcSqrUlbFSge2vdwGctUx3TuYyJtPd7nBRA1xo
qv6OndMoK3URJnrmVQOJmtb9Qi0qAs0A9y43qGRrMF9HzJtF3xTbW2p9mhnhMgmc
HCx/iKhYmaSEKvAjlViGCm4SrK5uho4bDnoc114mVxFSBAVDLSbEEE33s/nnbGFO
Ug1JNTDjvRs3BxGHNsNrjuvq1wJ7vnTN33bXJzWIpN8C0MNKAoAJVtdutvqTIPYo
2RdEvfZIXS1wpHbpvuQJ6x74+GqFAeuYwz7v9uuH4SfE+2SFXfYZ5CpGNyv6U/H7
TNKRV1cyomD4zm8oZ2PB7rrZzTbhW0YTN1cL6VvBihhOKHhjnqoqJ3MXKE9mIy7a
OnKv19Wa4Pu8eJ8MjjnmbBbomUeiycGXWhLfy3tb8BiAxIChgGKw9bl/ygRv885r
SfiQNXzW87vHK0GTDLnNvNdMgiD0nURYV0iqJAfgQJ4cfKb7xP8tMy3yYWU2k8YG
7rvmc8pFCztpIlrB5It5Jcqr3LNKEbhjnRcIHwmNvkK6FhJ2B2CJdtgNZ7rVmRAV
cUDJD3pVO8zYiIaTJvwHunhJMk3km8DDcl9AMQWP6FN/J0KxWGOcZ6lWPqhXFQ46
JBIf6j4uRiG2tYSbhOuIBuEbXkAM904LbhC03/Mf5pPwf0kpJJoMW+NzypS8qfxE
XXl0Ouqx5ntGfvxZ0ocBSZEUlhsP7OQLUHjO0rzVmBGQ9lWX3n1czEByXbrb0xpR
4jJxPHJAJCN6XTxfIeftbaFO2wEVVPDNLvpbi+jUDQrmMihBsgEBOlqMogNu2PNA
QYT99heD9ElDQXG1STPpJwrYN3mTRfh9CzsnILQhOzbq9DHJTauXhR/MyssAbMHJ
mc/00cu6mrMILtYoJ2CS3HRlNLkd9rv7xWUBmz0kTrlJ36Tl2Tjvwb5Eo/Fyayr3
Pmcvr8NtVjvy/Kpe2RSiCTqlGrQis0UB5G0KQYATwGSScSDPmqAYfwpLRKWLMPjv
iLlWQvHOURHXBAlsYCOW0qzxOOr0LYcGg+pSmNRSYMT/JGUkBhjlFewXDcCfcSMW
zTPJ3tHs0dTJcKQUErfiwNIrvfAclGo6YCVPUjwVnOErDsYzUoKLDTqLsrb9cpyV
ZA8FuVnJZ98/k2BgdmF5otAljTFnNZIau/eEiW1C2T7EzFNihpZtwTKPQgg4kOuc
laDQVrHII3BoQkyqnsFkAJDRzgxGAzE66s/P/hE0KTbhhi4aSOWaSmYPxuzJ3MoQ
bE+3GcFUU5UYYmk5Br6kPS0+h+CG4MvWuNLVdni6LMifzEgq8AAjlw1DyQI/JMrs
p0g1fly5yD2wUfp9GmY6tbNRrqjTPpsUkQOjD7mnJGcH2VPg+a9Nh9VcaNx3dprA
Letn3QgFrWglWY7oRLX2bXXPv460mkPQgE2jH0LD+d+hdDHtpFaY1zXb2Vi7ORiW
vLiFqttRrn4JG+AiHOtir5VkRn0jzNK01H8AjM5IPqp4mo5aN1H4Qk6QSi6YKNDu
B/QI49Mw5bnl+NybeDz2HogxHR2lbzM94y/a/FbCFKeMB3VCzVlXZ6kBdeD5rb8I
gmEOzfyQaE7g1WUHivxjD3ELlut2Bq0lt1RP64oKYVP7/XFWV/QheMJNFyJMi1qy
3iDou1w0MavssdL7640k7aUesfcGpiclfXjBpd7QsV8D2A1yuQLSYtgGCg2DAE44
GQGp2e3SSFy57cL4t+7yDv+gk996DfmQQez4Ca5ARyNh5fPvaw6aLjsdv7vW+Jrz
HuU1M9PUBwGpo//yKAcqhnrtoKqHcli7DzMgw8cepTpvpmR9GxeaeM56tvT4oktZ
j+6hw6SefOrGLdeo/oRT36bN9vOwiHzahZd3czUPsyczgFrbjD3YTkttjq0KdjeX
sYuY+DkKU6uiN6Dt/AyicdMhuyIbG1CKsFztoTldzjioXue8CDR9WrlLVjDSSSAT
ScA50uw3vDJinUk3ZF8Ip7+deGb2cyOdrwa5RVb8E8wgvpUFxdOpUrHeq4FhU+6s
3JPz2FxAQzrl3NENIiUuq3jCJC2++Xcr7LusbYmKWYRxgRmOEK46ohN8jPb3+KzB
16IhbjT5Q0+dBwjlwlJOII3K1W4j3ozgK6qPMeW+G+TBpExew6fjTyJVtxm+8cNT
+r5sgh2cEnqaLFbFGMD0HVX77Lg1MNR54l0pQ3kj0XoWv+gcBCq10tm7FzeK4r5b
x964Ij+ZaqXQmdU2o1O6QbGUhSnhQZXga4HjgYEwEvCIDXA9TCEvk1f5bCc2IiNI
ns13qXvBYv9o7EDhfI24uWtJFDKXoNfVKWk/YXQ11r4NJ83Bt9SvJPmT1gbYtzPZ
7N1JwgKsBORVIJzqRzNH2y5MKXROWj1+UZ6X5XWaBcNuJqoKfLNMwORqQrRWHKk+
vKfrSaudQWuNTA7fRZHFcq4tJuuIUjEykem4Cs8/mDqqyFXvnEKPqbkiRWQ7MPqG
m5FDhHk7rk+VjVRoB553R6xG+WDk/3Ww78UcjoJq6mlzKvAJDrSFycgzRKp2Neft
MnKU2Rkv8p1IR9TcA/x352/EIWv7zYu0bzHIzbJl+y8ZwvpWEVk9aQB0oKkhF+mT
28Sw5SmmyVvl8Bv8mf4FfeFJ/H8hHWqemPnmh4yXnt0W3QeO+d6B6caXhiPQaA8l
qq5+QqTNVReCwtiud0AtpIV1dDLQinN60yfM60SRpZUoUY+BftmtpnKLEEDTJSqc
7F3H4qBLFbc3ALX4R2euwS1DSekQ1qhg+CiIfMtGeZB0j6p+mgUumKL5FCU2PEwm
VSN8DTMTuQ2xg5ZsfGCodvITsKIbMWIwN1uEglO5yhludXfj3cd321/TvcYJnOFK
`protect END_PROTECTED
