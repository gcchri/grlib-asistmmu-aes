`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
og2T4luBfXpKsx74cKlyZy9JV9Dhs9M6cASsYhdWmqZBIMf5Z09kOw/YWRkf2bOZ
TCyXwd3ZM5nJRY3SLuBttPbMBQv/wxVWjoTA28qEnzXGRrGCggF/8qt+p4aIzrUU
i9KcxCx1eMx/J92X4cd3O0RI9/kmvUijJfT28mpjzMazVJHaC7eexVqCkBSNZq+P
djGROSUYXW/oct+JjJKw+U1NtQcSYCnnkHA/v0UV6TgVsgBIotZ4XoMWx/1ru8bU
4c2fJqVrLTuSpwhSwiKuMKtyLucDXqtTpbHQgQ1LMEqXaBuNYPpfprP09IIegyZs
J2fvOeUfl0/QXBxefviJ/nuJEdpOrT8L/+p2UwbKdD6u+Gd5SgL2JZqPLxcWMl33
WQJ3mK6oZgHGF50ZDbMe5yl0yZRbuDqB37jG+hawNj9RKTOjWPuHBD3DN5hf1nen
Bi9g+a0dZ8BocgS+Abfc9h6pFPmIEUd/jb9QHj2fdUInU57sv/G6LT2D5phB5Ckt
`protect END_PROTECTED
