`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJy+ThLwWZR+7HDPEiEu4wYLTC7bEPGogDs9PKrqGKPJzWcSjmxMbJq3QQhClCA2
2NzXyhhZWO6TWSRglZeQ01SNf/Zq0Kvi8BotB+9mtqmrEv2KMnKS6gGRGH99SznE
mpE63EB/1PAHDDAa5FB4sHdqW1diKsWY6rLfB3AEJQBY6+Np9YTDR2Iiog5M7lM/
U/y713TFDbBXT7zcLzp7aWT4JkaqsIx7rsSCE9D/ChM1xv/CBpY2qUH0qYVROp5l
kQzXx0bAoj6iQ0j4aRobvw9P0pUg+f8t2AIGCBrwqkPz/5YJkefyvDj95DhNUhtb
D6lDuXjuJj5K2TLyyfuz3VSCEeYY81hRpWnVfc2TqzfoHgBxmVkqfOTfViz+O4GR
98xeJdQTTvFfG1Ex0BAIrswxJ5N7rgK62guusps2w1o=
`protect END_PROTECTED
