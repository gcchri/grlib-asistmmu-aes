`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wsp/9KT7/XkcvEGJJOrYXJ1CvW7TFgRIqQKXqxOhNnRom5xWkZrFCfZnFvW7A71w
qiPJ/CkjDEXBQc56AlrQdG+iJh8LSZOglLalRbc7hIKXRnyenAsVkxEQnx+of3su
TzPzRtfOSchT0bhPayYhQBHDod9qWgsSQJFbWR0L/hpWVGCJu+0OifrpXwcUPlcU
TcekERKgaIVPQpEqQ4BZ5g==
`protect END_PROTECTED
