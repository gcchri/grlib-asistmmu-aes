`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vv3lEs2gFNqJ1x8aAO3S/xXIeNvjy5g0oHaKNhj0zXFsxyo6bswoVhKwU9OffziF
t0jnrqp8UgkgffPQGWO4WT1B8I0bBKSndq394zuA+OcUuXXh4SHb6aVuol2DQc1R
5Vz54Pe7HCSTXw0fEgW5oJtGjcfHp4AOpKA+iibtzycoWWIv0brNfcV8hKn0xiz1
XVglP2CQaawB/8ZdwAQwETHOPjTjdIsdyCMY/hACwdOCIOBoSn1EhA3fq1MSjSeW
NQORBB3PQ1Xd20/uzwqV+8dPkWST0EIo8DexVAVDRE55omOKlloMfcyZRvQmCfQt
n4HtcAuLq0jAbphZtYT11epPoBMwdr2PfdrtisiE+0ajCgxtyeFJBmDhVhSwNaXV
IlZrQf+oytQWS62ZtWZKr9+PgedA2tWlWFwThBw03SZpF3BWu1q57ngqEfoyjUHN
MIHQjOscx6ajXVsftaS9tBSn5j/64EJc7QFG/SxVJxNg6Hk+G1oIKhEEt3E5g4sG
MRsA3FPLeZxjOG3T9xuF/+ouTZrwE1GThXN2NmEBChYgLKJvS7hE6RXolDMvDBQe
TGETiELH5lAVuKF7Y43OYJu2hdwen0nMypA7zroqD0WqL3nN89uMkHB92iSiS5QP
I6FmkoAAd0MJ9jpxWOnLKWjFaN6Mjx6KRXJQ53df2cYCntc/iCS25In3slLLzs48
AH+E91Wkk+iDlneUJbFUznzFDvTolsqJyGpGF50M6opJzUhYlnyBt0dhu4ASYHh7
fPe1AFQo5nbgzd1WV3yaZZJxMCDZAu/lsWcHWEcgbeyH/bTq/XGoVd9mMVykv85w
ArjBWjSjace25e7cqpeYuZyz0eeFqo3GpQcc+qKSZFa6o/0wy2JeGEUzPu4Sw1ob
k54UMH6Jatfv2XOgrCN6d3WcGn2UgHFOfuGT2HnmPuj8QIe5lIUY8roR+9JtHBCm
xR+4xzz294r3m9pE3HqkyXJ4IYnANufbv2Niq5DV7BWEQgz1ZNZ0USx9zsQx2QvK
YaWnvtYDB6xlcqnJ2pDc9jXo7nkvSG+SD6UOliWjU0QxAWGwUaNXIj3sdBh0uJIE
rWldIkWHLhu5S+Riq17Fh2ZJY5xGGlk41djlYO4tjt+xzSCGGnYbfu+5eTIhZjct
NeMWHkGpTFqj+dmcssC7baKvl5ox2BYkpMpToc588mB09NT0cRtkoCZJHovOlXEi
bCkKyLXaHsQOCpRuM1Ig44WinclnWqs0vXlPTBAQt1rbh/rtu+VCEavYFa0I6Xg1
6F2bVhNdsETyrKxqQztphGs5+J/4CZgC/0ct9DZjEtCpfxxcrceFRosZ0lRDW1BJ
P7g+3xRolKM6zSBRL3AP8J5xH3ly+pJP916Fh1n5X3IToGqwPuYIazNl84ijpX6c
T0FHpuyKcI9Kedc0hZ/CUX7xea7NLeZITKWgBqFNku3Uq7wqC3PsGMBfucsMQa8G
+WYWACF9+RSG+eU7LedCDYH0W6rSF5gpGy2xEu1lpyNkwXnMEJDiAIy3h0PoUgec
Rwcx2YPH3sLN5iCeqq4n0F5UnUIFes6SNiuaZKMmIQB7ZLq3/0cobSWMaWlaWiNW
dxYwWvOGNBvhWA2WfPkIPOg3rMiPc4PS2zYWdoCWehQqbuISehsRB7mWLkOeXCzC
/C2EJVhSqb/qt06XVdn/c9GP6zFOplVfNTVjiWFTr8wLCVOUyrXVIEebpy+hC5XF
d5xRMKuqafJdhu2g6anLcg1EJsqALrBM1ivdT+nBWBnpVW3ky1dCA1Spy/yh1PV3
lQoNP81iL+rakWieQQiW7iQAXe5WEgtEeBTXrHMvSMsU8dDjxvdQ8B8+JIRb5d2O
G/Vl/vDGzLLpNK3MPakxY/txbNNfWm0vWPoxuSFjjdb37HcBr68uo3yK2+lPmgkR
sNXsMJnD9FS6ahYEI3cAh6u5rFzcK3ASQC3S3BrQxKRnwqFa/gq0uvZqaAXM88tt
r+TfFupefVifoOc0hifBXgs513eMc+f0l759lB7c0oIosQi3cepbNOXZFbacSqGi
fmJ88Rs0N9B+og+FFAVxFslP2iZtTTafzNdwkwGUXSuBHYhKbBKLxFb5S6WaUAah
CxrKXcTcoivgaN8+A6EbA83x10IuBMzZSw0G738vgEuhNN2ZaYk7E46wkqtPUxrH
t+Rw9TxtGfycz7zBf4cUBJTa/Yqkuesq6ZTNA8Z02WTWzIlsz1zfJcRtQx/pkWJm
9DZEtdCHpO0CK4D5qWtarHNWLZae9eBZdclKycjigtMz+qAHM3TfBe/00kw6ukge
cBW8tjE6baSYpofMozdZfRWTCP7apRcPTQQXBTwOSnKzamRvGLRuG2gzxuwUMnB5
0W4dx6by/zWg6H+QDYnc2KRJG3XfsqYxKDveHrthaIMRjbdi4BQuzC0NpJvvZD7z
9x5pEYv5BpVk4ZmTmxsHGnR8TiVzt3ttG9gqxSfNd2NLNpYQU6x0EO9Aime7ot5v
8VCfC1K+dOGGuL98f13WOMCVzKkvwa5CdFt9U/g0PgxPYV2ksYYnq7HfLB4/Gc2n
Gj/DPmBWiA8phrZe+2jNZBd0OGczdLlgJ/KOb3TTyF1kgkEzDOcvDW/MwXxK/taF
lD/mPdcr7TOL6n62sky2a+Egel7NISH4XxJVz6/IgT3MioXTn/5TKhDUOhILCKhQ
iwNJERrvvXMi287gS6rq/EZc8+uQ3ISUhUUCcQAYmpEFyUDAJtbOopw+FrtvP4Qx
vhJn/U1Z0myDIUJh7zp4b8ldYP0q+7zMgd9rdkEy/dXiOpcLMqK2OdvHwl6ApePD
qvpn4/pPY9z65Qbipi8W58JO9JTYQawN5mPHX4Qx5jI=
`protect END_PROTECTED
