`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgh8pxlcCh1h2AuKAzfzUokIKs5sPQiMOGYX6itjKnnShzLrscGf4Jh4nshzrDhG
z659sptQNdnzM2WcRbxVUlVTmjulGrD5RAc7LD9qedh0kFXnYzwNAiyf9qm8kZn7
phT4SnHIfRpoISxoPfi8zdTNq4sl8JWUBqKqRvu/mQ9yD9LwCW6pKs6q74iHeSmQ
OHj3q6Aq/4jE+oJ5ayjy9Fbjcbx04ZhRKGIZ5/5Gdpf7A66LQ8XwHMCVQkcdHPiP
VEJrbeLkGMc4HVk+ZVJnfgOx/mx8aObJvufoy16UEnQmvlPqgkxBboNlsJs5swHM
bOfoHyECEPowE9I2dXW0kT/Cman3erofI7DW2L1ao5OSMRNUkV8quF3fDsTfZm+3
D2jAKkvXMTaKhzyGhX+aXg==
`protect END_PROTECTED
