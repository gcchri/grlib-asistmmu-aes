`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
22ceoIu1lHrr0zlAkNbH30wFDRVYSf6KUJigtVjriaWoiiZLjOQm6sgH8Bt7xhzV
CUDreuLytE0QOdJcnsrLLXh1JJH4BLq8RqNVSNgok0DaeVdmCpPr6f1Jwkuh7b3w
wcSqtJCArvI1V4jY17H94Py21qChDc5YqmjXDEomJdhKgflIWSyxB4wCiB6NxNct
SA+EeVePJg7xaarIo0B5pVw42Z/bmuxSCo3KOG8GDBrN8hiDhE7JbM20Z0SrU2jn
+vuI7gIZBbIiN5lLQuou7Mof9WrNZ3Tm2Ed1WpYxEnkQ4X/WPKn/EmGy6YqagFce
`protect END_PROTECTED
