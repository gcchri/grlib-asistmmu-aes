`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BsQgTAcUxfyC7VeNu4hCSE5xnGRv3XquqR04SEA4ejHHARLuQ8Zmj1RTlADnBk4x
yJn7RSRUSk5DhYUjsN2KZ5dSgy+Vf6yVc8ZvVOeHKHz1HHBAfsKPtKy7GcWbWWxB
2YfoRqIt26DZCSieYQmvi/KNiV+8nSHBmYVbozxxgv2+4AIZbuPooVoTpBMMmS98
BdUpxVmKpYyXi3BkzW3l2DzONNUAd57Y9QNIvhEjct/iFleoipl6TY27WDQPkIPx
Q0viL5jJiogDwS87u3qYuQ==
`protect END_PROTECTED
