`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MNJh/Gae9sGqEHAe2g9SOHmW1EDxJWkAKQj88p/+QG+XYYnOSnSeJ6iEticdtXUv
h5uSedrBYWhDm2DciZtHIOTUczX5Jc+GYs7qAipB3d3pDFr9et9B1fr69NpJeXk8
7Vzwv6kMKmUqiDBV2eHUAisHbPv+B0hqicdYGNECZ/nxU5vdxiXzLqX0/NzAU9iY
8lNl4Uff8KJwW1IsKDQCkwLrm9kLtmo/mKou+QJPqLYvG7pgfvmNoKdJzbB8fxSs
YbFE43qIuKsm5Q8CD6XbWNomC5VoXNRTV6BXD0a5WgLO3d4KytUSnmfrOXY2DDDw
IcGwsWb3xIqK0BntBF10Jib+/eBJYG3+uMDhDNJ5EugFdrlXENAzbOXtvxqkmRnZ
E/GloXXPZogNMHeYzJpYv/4Y3Kz+oIGbA0L/lurh1LZmFgsHwmiEJZX2DNe7c4CL
xKYfCGFKIrnjbdGp+bIFAVan7cxRBbGrP7KPoYUvhneQVz01JVtG7Mrr4DBDLRRP
`protect END_PROTECTED
