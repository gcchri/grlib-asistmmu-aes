`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VTeX1rSTsqcmnmXsynQMN43AA/EZ7DJvpOvdux/rMbeR+KN5Z3fFG4Qt0dzftpfZ
TE7vQgbs11wCVWZC7rEI4SB6ZdhpMrVGCur+ejqBHLSdW4s+3Ai2l/m31btb+wsf
0TBgCMAknIP+33ui8jaMDZrDcLxbs5+3uTitmoighLPjgIaTAtZVYPJq975LEGjU
zwEqETs9gA7S+Sdh9tdbSsSa3+ORrCG0pofbphmRSDQiFSr59rNlU3MO5xO9PDM9
Xi0I0rI9H6XYNK/HuV1Dg1uSePztKwVOe+K4Q4soQGn1UFzXRaQO20cOhDqy7Z1T
PEUPq5qX21+9RBtIFtrRhxgW8HhU6SakPxGXqAOy5ONYjepiuqbZeAQtRT2enXm1
+nSKbBIUnXgVp0d6fVMYhw0TcbydVoZBhmf7htgnQk56op2RKyOeRwRQ02Vwe6VG
LGrVAdh6tnl9ZlS4bW7DNpcd82XPGnXp8QwwO/o45N62T3DN56rppgP5U+zcIZcD
0jD/epoQ8PgBMLUIbO8XDw==
`protect END_PROTECTED
