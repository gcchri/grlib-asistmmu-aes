`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zxXsxT1XXCwAuuz6VFbWYutWlx7VuylvRXX9xDVEsMzXoApKjCG6NtP3fSV0NBmx
f3ReQywOCBBStME9llkQS+KfQ1RTsqkUyOFpAW82PPqWzp+di4PKrAQ3HiZrirGK
e1CXXiM3HZ//7LNcF7JibsZ6eYDvbzg9HzFyv0Iu8DlYSguLOWNhXlBWO5/clGKs
dK5jtv4nbeFkozoxgiKsBOh8ARab493RMhAIFsdF0T4BrdEf3RHR0Zxt0ynsvqDV
7Hc2q3HvSkiR1pg6ra+dDWsS/y7rBGRdq5NE8e/LtPGV8Gk+O9mbbqJGgvsfnTor
W3k8ssZvRoIqQc3dx8vQkRueJHIG1x+COJQX9mvw21Wn/WwAUZVGSyVbVYsYp9UO
4tUI7HY0IfT+FAyc34erqoB1iJ6kvv6q8ixcU9uVZPxJSy8LvHhY51b6f8RsZli4
YI7A32iEJxP6kdmC61eTCNe1+fuzPlJb27lMXf9TULORsovXUNczxUftSm3VsddM
1hZtaenNvd3KI0khu5NC+DcDMZ/oXtBuwk9CXhlfv2LOyfsx/VSnLZ4apVaVIrtC
c99DKlLXwqIBFeL9DXtna5oSUIeW+ZIwrb/0BolLgnAmGO4jN6HcUtRLeSInT8d3
/kcUETjcxo1gC8B7cUvhNzvcqHlBLmeF9ZIuF9SSFAYRTc0vn/o4EbF8GiGBvqPf
ujiWVQG/Q3Cwgsl/3MDGsL6gFXWMzsVzaJSy8blger1uY5+Da+T4EOXnw54vVt43
eSQLAaerlYeaxxUxgD3Sgif+9WaJyTRMSAH9Q4OmRP0G5cJXMPdt5OnmDUjW+1oC
SEp3sEfOrmhGQP1WORb48sP8lo+iKa6aqzXxSy+okB0qdOKUTjeAJ3UNN57i+hyw
urjoCEZPaCR3vFoTP1aUKodM1Ajs0Dg5mQmniT6RqpiS9/JoJ65QozLS2zb/32fP
IXqQ+qWItk0DbkYZ5qnKXf4jskF3J77DL1uGCTllUqHW72SudSn1b8zvF3NnvPEY
WHP2vIEuO56pdxMxcjUd8s7V1tEpfTokkChl9n97+b64InTtc7z0tXwNw0yaqHYK
BCsixO3J6GL9I9fF58KmiVqsPonYwAO/jh3/1bjwxT4YTWC7RjjD1Yi+kUfIs6bW
6kIwuFI/9nwMgkw7loeTeF0WUwdqibefCP8Ucz1OIE/yQ5mExYMPdb37g3C8ygWL
V0V8TYUl5omgteWX87D7E8k1b5V4GEha/5RG56tZMdrFORRMOK+2E7zo7X4UaA5S
ajXsBTkm+DRqnSD6QKwd8iqTthuUxUtgjBMoVbD9CiyvCzGVmTLNpPt4rTNrIK5n
HwNW7nX8F5PMCiZNdg/t56j3EfZSEIpJjNaJTySlYITb9gmAiP0t3EWTGl7zIzEG
ACqAHfQ4mznr3QrklPYlTNaTnPMRyZUrLFvG+og5BPunSkdbk8pjBpuc5b/o16K+
73jSltzfbw+vn0HobrccoaSEC6xeAdn0QW+H07RNa+G64u0glqyna0xKkQfRnZFY
NLnQIq9bKl/8mGdo7957oskcFLsE/0wEPrNpglCTImESkvKPlD6ocfByCqAKw85p
PzuWceFY0mhqKZCbB0hxIppMbCT/H8bgnN4EA8vksGFLzlVyG6gDSNBTALH7AJnl
XbOikmL9iutymoRlGzmILImQ+z5toY9TI4DCq+FGU8tIfLXRA3+VfIay4lv/FxON
GaiYCeBWSzY5dQRsB02UTwpMgJYsRhkPWDn3Ta3IPJ7a4SLjgZZxRb12UIAiImJO
rduepGg2NZBjdcteYpZJJLD94BSCR5MR1sSjzd59ZXjfVhktLq0z7RhnoopruuV4
juZ2GmNt5VFAof62lUycafkhfIFcgSnm10q5aeso7M39F7KULA2O2PIin+66x9aV
z9iVb6hWoBHIf5/rYUL77dfYGkULX9gulXi806Zk+HLaW+DgvmgOlpGkC3FGp9zz
cHwK9DRL198XPqRb+HT7WFQzlYLrdBWqae+BSAgYa9IMYzBiRpkEu0ZYP1n0NMBP
KsvdKuE6m6yuY0UBfhM2YeCSv9a0ubfhEJeURyKRP0K48OfTaTIfqJWQke4mROk3
CobEANaX4ptsXh8+0msG+2aASOFpN8uzBuSTn6UJSbRqB/yRkcvFbkGErlWU7M+C
Z7+Cbctvo4I5awbwiyL6SnW7/JpKZaUxCIDRWcEfRdIYofmPV4kESjBG4BX9UF5+
6pwCJ+R0rl5Bq7vlnTLwIPtBarRqnHgdeDxDdNodXi/b3fRZe7sAEr0wcfAL0eyn
hUNs5gvC8xzycNjuqK/kzBh0+u0ZXb0sKKYMbfHLAunxQipOUi+5s4ZDHL8m32/q
uV1gflWx9a3mnRi3oZsGATisDfTbdVHZzQW1Dtj8GjalY/TFE+/tAll87Q7QbD0C
HfrL5rGelRnT0xqfY0VC2zHQyVNOTTYQkOq1/Wv5FbzmhB59Ovot4xEFXz8LwWiJ
f3qBNcp8aERCna4j9rHleYpd0Oy+j3Z5q7ScdvjvfTbttYNFlnuqtimHqAkUug97
FW788XwaGaliEpFQUy5HTAPTRs72rdzLYVkbGWtNUF49ciVn8MlEqilqqcTDQ6aP
1+J0tiPFlBM2U4w8n7lNq48/5/Hhyuvj0zxxmV5BkLAVHjzJwMuHDHMT7IgU3Xg/
jsr81TjtpoMD/N0mfEOnoJnC8BO6o7cUenXvKInpd7V0l2FegsJxpQaCT7G8rZ8H
aYQeahGSm/fA9l48z9aqBr0AeHZWNSe8gOGlwE5DXEF4Iv8kqGP5n64afUmOqbqm
d3FB0Rr4g92olmKYqonSQ+z+iHbmK5JIyL/zVEFH9WALcTYDIurvw+LlxLMGa3NO
BT29igiCWJAlmylAC52SMUeXEXgLMXLBK75rG7xM5HYAYpwd7mxY1JSnrG2NUQ2j
AzSL81OnF+K8nBPS1EXnaFexYulu9LV5AqhSm7JFKZZMDx3YoxMnnoGTHQmIevKR
vsV2Ky3u0EM9fxEtKgUtLBa1VDJuogFgxU3wbDbPk69eFWtWYaaWsOSLFnQYb/Mt
ifgLX3e0oS1ibzO9ibi+HiaP7D83oXxobfaW/zZXsjTstZJ54ItrO5HxlAojNeFK
3OkOnPZ1BR2UuUqhqMLIYvOxbw4Muu6/B+OPMNwTZ7FAjNGkWEfq/Mob+yUHp7gj
r+/ibkkUoCPRmBb5+1/lSHB5qbN96f58APGMDXulnyhT/6uOPNAcXITdmPSCHIyE
0sxyj23tBeH4sWXalpJgt8uYOkU8kpdsQn+SEL2qWgb+E6jh73AG7kpQEsFcaVBl
J2fo1J8k2JUYecKInIcFGybXGfE0VcZIA4K3vQT96forV6DuI4oNtBIe6cXKLiF8
bwYw7CPojHiH1Vq8BW2o0TCK/GoXDTQJXgu/mLMc3JH5b3S/rWn5UlmbKy4tjzGr
DNo6lIk0IV9/GncEAy4wDdG54ce1Wae9XNYEEOFDbObJLvkzAmfhgapbuMw8Voca
XmyR87/zrcVbmj596OyLHUbrkljl/Uh5d8uEld79H7PAhjLqc+TgRXhayI1Ucui3
+zUz4mZgg8PvXUZ2jCPG8LIIU1vxKqHe1i2P19A0VjbJDEqLyrOuEbArbOeiToGn
PjMaYdDHzzbC0PX/FN64aXBV+AJ8Ccq1C2iKJ9Cdx52D2V7d757njx3Iz1WGEJkj
uNIfChAKZqjgHyvMtOg7Kyi3w+m2vQ1bNCJeZ9cC5WLVlTrmHvUpFSSQg1dlYAg1
msBbF0BtaAP0Aw+v7UgQxjledkkKqK3OG5rgtm+8L8uSAcqMe77IBARGpBbjWIb+
g5jOVA6hhcQ5vDlUFK/pG0OisGIiSWMCOVbP2heKPyGraUaiNcL+vPWM6nczqwSS
9ACMXS7X1kdoVmzF9deuiIx0wlSbZorvY1wPJAghe7hB0N4/eF4mhAtKSLTaajR5
AZ7VuyKakecDWw18QeAvUoOD7yg0mkhXMLabN1IQjXKTrf2Y0V7/9iOjVpgJthaG
Wj0pMultMXrUTf9XPslwJ8UDLCx6AKqInDbec+FbLaIWIJi0e5U1Fsv7x3IU/+nZ
wXPbzXgQzWMaSFItI9bIwaFL6eGU/xLsVmRCYq6lIdmcYpM3UTrumQ4w9DpBOJZD
JUxO1XxNbkGOO34NK96ZDzK7Hh0crlM8d0LoE4hH6f+ebxcO4F+10UUx04vUtDSv
ZQwdAVhRfH4zUwxFrvLrlMop1dlikE8D54D8pOIOOFSPQpiXuCbPXL4YbFEMmScJ
brpCwtlnJCz4Ymd2f+b1knyNdilCVnLOK5zitlIXKyywH1RKw4JV1DQEP+E4gmnf
XC+CkPrJSE2ZBWe+snBmAUCc/yOZQDg2TWG+05nz64wM7Sm1V31sLr+nOatu8aBQ
eFN4neLpV6womLNHZyxrWpkv4xSr9ccjORdVjhJmgUA+eBCFEx1AFKa/RShkEeoE
FfM57pCqI9ar1ZkMcaFHZRaYh8TJwRHPRCmNvIcaIUeWmJnWNtufs/cHeYacMPPI
UgNQgdyX7HMWMQ21J0agWj+/Zod//ICPCwmt0Oa9fADicUcADBiqC49gh57533yP
33HCV6ZHF/Z/1USmx6BnX7pwnPhoUgplouDe7z5umRKrBmjLH0uGquMsCqAA7ik7
pVB6+x51H6eUef/9S3i6ei9HQ7DX/HT49hBHmR9JNATPq1y6KobGMLfuXubVQwlE
qoX4AvsPG/tdsZ8f1R8J8UjlWhTPE7lEG3iy1f01YNpWxgRnlHcWT1fLt6JAn8Nt
AA/kRq8vQgNam1AQGq4NI/mILwmD6dTDj2mKLZivb1DYVTZsda8+ZQviqhNv42zs
Qfi9DBZo4dysl4Gs/nHSOEePbdMNsBZhRYQUAlXLh8gj75ssz9HL/QMnQ3TRnVVp
iK7DAhLHXOyoK/NEtrs0rkpooesVjrPU2pztTpl6sc1/+c6glwBLCimPiXt8tACD
pckIG9/EvjB0Y3d3SBMVGne6Yn9Ni2D2uHOFswGbNK6QjlljlwwsdWlKjJkmOSJ3
yaSJMU/i+JziVg3S8vDBOPU4NYsKBGt5tUwYJRcxr3U6y/4eFB8PkCPtURzwEjk+
jOYk1WgUypfCOcB4dicJ56ZcbFpdyoW21gDwP0GIoNkPtUw4XCRLO1YCo0JtmMNO
OjBOYQfeCOLcvmDImZ1KJP9KBjY8pBmxsWqVakeOHIaTJd8PSOZzcuQlAnH7Y8N6
HsW0lQE/9bn/zJpEBInvMu09o42pVGM61uPILQ91nwpWj8gAA4rcasFD0leZWR+c
xp7qVLBEVi7Uc1Ry2+rVae76hPWaVrEoDhEwRydxxr63TNaWBtQemCvbRA5Q9L1+
xKpQnlH+vYZRdfGaFOrEUerF6JZK1NEVtGP9q7/gu0GIJ5VAhHaiVWJznRzlZzd6
kkXdQ1ApOIIDytdWo2iNVX+O1O/cXpI2nutPqZyLcWM5Yly1+sSUjzAEvGO9rdAD
PSnFzlyLr9vcmB8vMAnT3C2rbanjkVs2kv7wZ5qVTVGdMZAgfRFwYCbYH8+gdyfn
eRU8ANW2IYoYLEhRRUaAwSN7o9E88fUhRy1qSAbGolQKOgxNiNAyWvO1kijQDRct
SaYa2Zm34CohAHf2cOEnJr6shyZ57q89xu6MXMX9z41d4ac2RS2JehX6OEFKmKiJ
pvqFmkPrrRCC4cwqo3A3vRFVqDveoWLY5VW8A+84NbijLQ81v220pwapZIVho4Aa
hdvEirw5atb/i6fyHDaFN3mJibxPkYJuCu1okU3z1gLQXhelPjfTWxgHWG8HaChD
Z103UdQsHhz1fFh5cYTP/n5W52/IJpM9Vlxe98s0C4vahqLwGbBcbSLolrJoMV9P
i2R+BnauibfW/iMm33iu9romvunnyiNHRg6eKqeqT3BrUXxZfxuEk1ogZX5nFLlT
9nxYfApBRcuSRZwCgUCbxrakOOysqKgsvOC41+dYvejyPrZ9hv0E93PQWujt79qH
JxAr0nlMthXfmjTN//K8TlWQ6FBedMvvVvkC6BmR4oV+sJjCFXT4gHmtCfW+ohdM
aPuVnDGy0qjA+i2Oaxd1PaNc21uJ76ss7Bb5MIYR3EE+mncFmUwNU4PySCE9Pb98
CLTH9QSrbRifktSUwSxA1EQBc/ihVjiMnzcbYDO/04ky4uXEjTw3kL3hT3N7IMuf
81tTqLBxfUyeIB+d5H709bI6EmmBEjV1wAY9LL3u2Lq8v+xomp60y4h3av/o7ruJ
5KJE7mILCgOcFZ4TUBTDDZWOzRjwKCsWLkmkOxAZfQMt82+Y2q1u7u9Jlnmhq30x
gTQthr5cl4WdBHHQUN1gzIBbhTzxDy83AN22QOu0fN04hSHniAcEjD0UQxMvyD+X
KnX/WYv49PFthZCjgzJOmf2G1N9wtKKPSP+jDdvpPGHnmTNUIpzgkYbIEAP2VNEt
CUaMl5yZB2QMez1J7QvcSDZO0H5xctRVrrTKoHswF1UAhM9cwTR/G30iZOo9UabC
ijOTeT9jkGU3F1q1Dmu+fAF+DCcgQ/0bVLOPp9+2Bc6JcczMiHTsALYkPDqxy+WD
O0yZByhAgCjexxoO7hFJWSAiosMeqFJa4W/tyXbu5dLFHglftJ5idTP7Db9IJt5q
1i054dJo43Nr4H3fPaPyr5NiUOz5dnQihujpErcxskKkAij/AQxAxCJA7W7FOmW0
ZypMIqM0v1Us+gBtsodWJqqJ+MV4aCKJijMDj1xe59C1MOfKZy+dTVeQj6LQJZYw
Eg5SAf5hSmKZ0fo7nnkn7lNc93jKjr7PLEMWV0dR8BiYGTEgzIK1eULTLUaLFhV3
Jh3zDyJdwNdECOtFim9k17+pcqeVUlSRFyQ8/KxyH0AUuL+Tjfn2lLfDTftzR2Yg
FB9XaZy/o+6nNo+CKrYE054AjHC9wAxxWbsPscUQQ8oSv8o/5Q/FXos6Ct99g3uG
Nibu1OUiz2mnfMnH9Ra+bpgNzgsGjOEm0jL9LTQQX40HBcjWgHEVS9HzOFZPipDi
Iiux4yzWQRLw6NL+BivB1pu4nzRKaZ7enYc3kCxFuNfIo/McmqHkoCaO1kYxkRuR
JjN5AxJWKztT5VKdrHSHmdLE9LFQqNjxTG4D/GJruDt0FipIl21tQzferFQ+/lw/
75UBtGlz/bqYbNuiLq+q0+f0crYC5zhMEbqVRRfSN+MMef05IQp+lP57CtWepKCG
9PtpP6LnpYSlrIAnR0nez/f8xBJBgCz1viXUg+pVXlnrzykSGde4A0axZl1R3ebC
Eym/nWX6OTsmZxyJ5E2YMqH2dYPj+mluyPzY0bN3tiUGmpgMvhg/f+hobi7iMN+z
QWZkEgMqlujyJTLQlZUgkAlMopXMviuMpyEA8yk/q2lZEg/lVDLh8/11Eu/Rzcci
eOgyfcRaZ0kUJAIy6PDUNEFh43rg+2WDwPFgLus0Ve8GLDTueLDwmeG3NxdvEno2
RpnAisyfsfIxOpt1Mr6SuefN2EnURFjfrkLoJqTtJ3Uqt78m6YgRWBxz+qmei9EC
rM+yrC3t/yEjZloGZU5CH3lW42llrPTW7lQ/CYPcJkmaAr+0KHhFZtUMvQGxfvBs
7LDLeYKnVpbN5IANK4uytoaozXCymx6PVemj832bhvWgc/R43LkraQQHOObAkorW
lWX1CnOkzH/mRC2O6Rzf5EzkQL3TishWDHENlGNBXM/EmXQoN/ZuUlRZ0UAZiRnW
6uhoAuNh6b40S2P1pBX2+Eg28htpL3YSJMixH0pi90N6E97Ypm1WMshXBBE6X2y5
TKJaIeUCvVN5ThuCv71H+A==
`protect END_PROTECTED
