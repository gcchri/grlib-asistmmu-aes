`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9daWqJPZ9PzFxz9NeEfayDp1yJKzkgoaJUR7Byc9R8e+Bes2paEzXCeeyptjaK9I
VAxApnJq4CU/YSGvBWffpQbekmajQBZWPV3c+TEWgmGqKlLiJ++grhRkkQDOEDf3
dAiSDqK8seukecnM7YNExmhn9hsV1lL546CZpaG0t5woTM2mXsYgt5lnh9LfK6O6
jU1DadgTruhAuRzBJ6f0Tq1VQ7mPbeiVUchduFQtOzOmdzoqL1rb39E9EQO8PDuC
YbK74ikL+K59A5DuQ+3uYm05v7sJb6G2yUVH5BiGhnZ2uRSjt1Riu0AX+TQVm+zl
nKnobthgIHxQQZC1HAs9Uz2M77B+DXNfd7RI5XgG1L2rTYjl8BvR5HEtM/zFGDxa
+daBpprWwmE5vEJorpeAAA==
`protect END_PROTECTED
