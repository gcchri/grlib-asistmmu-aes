`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9jRJkUtU0bczWWNq6WlGx5JJkVGI0AWN3K7GB3BiO5iNj1LrFYPwcj58zST15S5d
ATpbKyl+wsh2hb70yNgOBprIIMsqlRZgHvpRF7t1oqbUAbttzKVkIZfIcQg6DWy3
kEFM4EFQuf0eE3mqFKdeynj0Xm94/pYM0tofOah9lqV4F+5YLAaBMMlPHqwFqirm
I2XwyYo49hSFER82rupn9/qYqc3VKLe0iYeXWeWKuKO8Ngi5Cn8eMjFSF4S/XfyV
XbRjE9xjZQr3OTlUFYHAYJSLHj/YOFsUk0mhLI5637+ckP12l56T4T4/LJlWmwzv
uyH2FMfWlEKHlS8/lUAJxXi2jzcjbVBNrt4KpuFPB5Gi2oGcY2JZzgtapEfj4NIo
RCPP9feylcMsfdJZ89t2gcACMg2OZeyYQRRbyG09zunqbWvpjhPKL5chyFdgwrdZ
ImRSdrQQtcfCQKz00XWcEU9fanWyYz+0Fh1sWYHBNEWfxQt6oDhxq/GjlW/4y5US
VXDxi8pc6ion+qW9srIQOs88lDPPfFAZsX06MSLIFg0n5Tt/TmifBh5GuRm+2ouh
75t8BotiGPetFS8ZpJQ4tKL2GsIuP96Q2K1Qwo7drt+vp2yy61MM2UZ+H3eFQDWX
JtBPvUbuTBigFOrmv6Iw109nvqYsMB+gLveyloKNtL2zeMLvs5kPOeWNZ7fzX34+
AXuRqnXOQN1kidVoA62eEIWa247KnKnkKR0EJCJj5cg0OKsdzwFz7InybB05cmon
OXg0SXjq/X8E+ViDo4MnYm590DbGBXPI+wZ9n7kXttsRl9TJyUqOZ5NYdUnb9DvC
/DccJQb/bN9QoK5+mf1csII3mxIt8bDz+Ye8x0LMdL1RIhhyCFM5rLiloi624Rmw
RwEuGDV7KxNKDUNR2a877sI1tvjSC4/tXdBntm8CtIoTbIxksMeqNcdplIBdgIL+
M3hb/fX3d9h3PpgJWf+4Tu61jVrWFl72uWe237ekqmpU2ZMB93kvs3SoArFw2ezc
If/kLNTF171xQpxJ7E3LzIYzDapX5Gt+Twfx393zyloqt2AQg1wO20nQzkdsarTc
efMNg6uMRoSJ2bFdYHoPJmFuK5OStAXU1aCPtq9IUP0=
`protect END_PROTECTED
