`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
srtf8Ynt1tuI6bNnoVYSg0WPBWXlqBiGWH4pn7lp1csIMqPAfCtGFP4DMDAQT0l0
TXjcPZXxCUDi9zsx9dveUGyiQUyUk3R7alGnyXyJO4LzpPAst98Rvtvi/vBxVsFt
33SfoI0JoaqeKIonpVh+Jzkc7BjHp81yEdVfLcPLAH25BnLoiwnE0yCVyC/D6v9v
1vKu3EhNPhJrYZML6EdbIL2CpvdRX8ionCPwPN0WLbMgtqy3M+1BSZx2zzgYWrrl
`protect END_PROTECTED
