`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3z8zVYVRjd/AjmI/x9uDf6mF+k+yS2xVG7TIIQ0KDd9Ub8G2sSKzrxqqxLVMpmjJ
/hyJ7rGq1h00vFzAsc/lq40IEue79wb8mvkyy8qpQhATSPMEDajLWIxWg7IlOTVJ
Ar1M8VhtMyDX7JDLvnmWQbNfpDC82EZtgXm/NGdUT30mUayJs70kJGFrRlPPKR23
m5Dd0RPrENqDgcDiLhCN69ToUCMF/TVS0IR3KtlA9Los47j95xJcT9oO9ZGBRO4d
sT/FCEsaHo+PhIUvz5gJW2RKrMUU9KTD6UaOzEVKxDjEdKoJ8A4h7xsN07PQytm6
`protect END_PROTECTED
