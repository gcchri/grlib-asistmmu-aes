`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tn81GZKsro+W0SSkOs2FgXSpXwT0fyjWsbEUTTcWXD7TBjE7hVUwMOptqt2Uz2SP
Zxo1ygDwJhbaq5xwdD5DF30u3atlwgtb8mMEZKnw/ubMNkhOav/bkQKrJYxeLGtK
CAheioZtvQZCk82hATjVdx5kB5C+r4ghyCMZVUhFdLVqge7ANrD/JVMdG27LHyHG
8L4pReGkNtBTjxoNhaIkU2VD5cG2pKIgWXVqvBocNbbzRkqqJZpAJBRiwGgrr3uW
T8JvgAnDhAZ187OYbMPNPQY6DzhRoVRUK7c4OylKyJfMlXb1JvvA0SLAwd0MIRKV
XHeto4SZq6yyXFUbSoILqHkh1oIJ0VXqpyzzhCnvLj2sjWESmWsMHQw21REYrFTw
VCqhyldT8KzZaYqDPUh23MAuG1ZUrvE172e4f1iIQoI=
`protect END_PROTECTED
