`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sPKKGXKVBcxAhmGVg39Ygw6jiOh7LptY8Dl5jhVzv/piqdvnBAn84aJLpCxL57ec
ZbRh5708bj08YbY4kD3XEvYTtwJqlThchPrDj39cobw6PpJ9K9nw2/lXtYSUmvlS
VtX2vmuUu8F353XENmMZUt1+jvwvoCxG1jNS6ps6tjfzyYSUnzXVwiRrevwFHOF4
VTxQjBwuepMydo7RIosZsTx1IFD5B5BRSMhTYJXNTCBWZHDwkE0rNVbBdpW6Nhkn
3ArqpuxY94vcQef9pJKYNQ==
`protect END_PROTECTED
