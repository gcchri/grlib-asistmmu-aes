`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Fy1UnkcD5wqZl9b2AkWeIuBuPfoCTCyWKFzmbIVozlV7c/EyYcD7uM3qSMFoiEt
4TOrs9ztYWdIv050ULHBKPVO/8mzz8CU9bswAz607Ciz9KZpS3i8rmdh7+V08i4K
ohnUJfomP6+VNMo6sCRh7plU0oBFPcPh6Esatr88BgpFm5Ne4vIzMHMfjAef4crn
0+EnGeB08K3+9Lg1AOZdHi0e8fsaWvDABTzfgw4dZ9Y0IkEHJjh76wt+CYZIxKOg
mpHa4Dw3dE3HxeUWBy+07btlkrYSROOwvHWdA1Tu/cLG0R9UnbgiDqYDITZsixlK
OemuM4hS+j0kzMJ2kiVmcrB4+703HNm4aOcJutthB3Ivm2no63PWaP9nJBbhPIr3
1XiXfVOiN/ALUuYFAwQfRd3zMVGPA/VUX/18GMEKC41bR7F0gPbVRpmUmo95hSUY
Kcrc8Pi9LZ2sT3OXBD0mPECWrGH9vK+RCOfAXg4OToIwUSQL7eBTJN1KHGquU09e
K3zxBDaGez/gBpuXRZBkVl7+nJ0yp9t40XFF2LMQ/O6QbM9jge3P9j015t83NwXJ
g8Qzc3ZyaaK3HCCvj8zUN5apReJjmDGLT5B/rTbcRTZiOHGRVkzmU4iGPM/YgMmN
xcUms/pOwKgKaN4YJq97zDQepzcr0YD5NDlsXgjcUFZL4lb/k7NUxuuVYnax2rYq
sRDdSv8EGOAlx/20F/dpPt9Z2Qi/vnAnefnZ6RdH3tQKXfEU1ODHy3hWqrqMUZqG
og3NXk7qMnbvUvqWGYrTb44AF6bMZVflPcVnF18IxF/9UseIS7mV8J1dYHVbxZJe
ejkUQ/vRFFU7jKV9Rf49RbynusF+sRadccADyFRPOay9VlcFhpqOQVKAcLXm023a
eG4AHeQW+N/NRpq+zi/h3Y/tNlD86c0I+ipbta9Qsxd+8SivrQaFR8no58yBeVs+
vvi/0Nqm8K7LgfwayJzkyQUaJBlLONGVU5X9CKEOI3sXgHgum+xKCKXQBzUlMxpk
0IBPE7q7mOyeVQHAd2gULY9vxQchKA0FeRW5zs5LjClXIPVsCiTcKO7LjnLegN7y
QyUWvW2jn7JqDckmxaU1njPFW9mu/+XleWNM2XPytt/SchCumPh5WoigjSfC+9Us
`protect END_PROTECTED
