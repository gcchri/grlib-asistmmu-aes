`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cWFAJiN9JDDytt835uMJoc2PHF8skrKBKw9e6PbY3ytr2VfZdtxcEi1cWSX1seTn
Pg2Se3+p8Yh+fERnyQSY6abtHbmaQxjuqUKnPNKNrb4eszeWd0Psb3Q28JEa4nT+
LSpJ3KrTR9AjiguGma299QBRY7kNHzH6FBJDFZj/y+JQp6i4mXPj5arDpY3847jV
NxYF3B4MMgM0wx2wNs06eZjJwJbzFpiV9CNekApr6JxU6i1Y5xKwzN/xrpKBu6Me
SHhcXFB2/K5Q1fj+3vSMGQuTRbdcGkgD1BVHiWDtNmU1JTFmfe2amh/4clpsMB68
ExP6cUri0zhRYTOYoPML6LWMynS32rWFIYISzypqTSWzceoyQ7MSHIOZuuEtx1If
0PAfNUkexzFg4XI6c6lCm+SStx40fxve7K47g0EW7sIQF+KiagNEvRmcwRu55cyJ
vbvL0ozA7gBppr6veVI69a4XuO8wuCeFpOSYZsuArg2Zvwc8RahdQ8Kw2harEhRQ
ZxmWq4BxkPebjb6sUo58MVKGElmW41XU2R06/HwlDfjNzUyeLpHY4yEp2b7dgV9T
wrEIwDag9ClWNBCVX8/eUG0Ogqx+7aKmhATZ4nm9kxlwIsrBfBLTHXzGvoOeRymi
F6hH4ksqlVwFPttLDt6VzI38rz+OFlLVU6p06M+JVko=
`protect END_PROTECTED
