`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
12f+Vv6QHT4Lxc/ijrUoC6WrR4zKtRm7rHbo7K32UgNIAp68VIgmlgJGO+KHU03Y
bWeKni8JHxLH0HAFOYgIzZ9RqXygGyPfn5TYm7YBq2tR9TlxX6GlqfJe0+oDi+dT
bAQ62uSBEU5thjD1mx/4Dtjxtx7EKT3ChWCbcpZonJgj3h3nUHAlf5KWDITvFZ56
aW29d3d4ZJIA+GMRJRcF1xzxbfHWMaIVtHGla27ffJG8ij9Gb9Ow5CrILLJjjrNI
EJMItHSJyA+ap4iRilrjPFp6F9yuHd1fg0voKDIm3fDYqln/4fqAh1KZDxiPkeDe
GDg4O5/TNCph42BSlzmLEGVFTp3j+y3qw6X3XvW8bAEroCV1CSfFUcOsirZz4kro
7b5ZLDCCdMBu1A/OXmRcn1J6a8h9rDRYAicoXxzho6+WxFaxdbMiPlbLoOq3CkQW
TfuFxILV/P3Hb/YXqMVpr/gljtM+CaU4rFmriIXQJ8ousqxugCYfYA7eTH4gSs1A
Na8hwte9BEwVtdggY/zPbYCOT3dKJDSmv7NkHSs6Ip/5k0fVaKZjPEK/NKAlCyyT
owZR8yC+CNkPcJpHUBfFNGEvwsCjaGPP6psyBc+O+brJ+QmRuYfz9pMLAR/E7aGh
oFfVzDcVqNfu7BAf/cOebtFwgCDPRR8St/jUP7l0QjRo9qTZOKdEfN9EsbD+LCQ7
ZI2LG7uuSsmcbd23naTlmUJasQI4pdwn55mVs8mNHQ++rIbmLEZ0+Objvhbdyqlf
dYJ8dsqH/wjVUYwRtYIQ1tasN2KQThD3+HMYk1KkbcBWVOz0xgfGrISO188f/yBT
VG6c8KZi8eqtuwil5INRKvJNX4RKaej9ZsUx++Qct5XAR/0NISuMKtdmzaIFVEU5
Uc6mPpyBXdAq5S+d8+RU6MRopI2pD5VhC8TNTgNPZ2KAJXpIzAvcENq7G7Wi+QKm
BG9ycM/NUl5CIiMEgReAn0OKfXP22DI/txHzWb76/VmFzMFkvYLFFxM2Qrl00hFg
UAYLEeqO2GSVBWpe6hrCAqV1qrFJq6u3Sp9zgMfqH7s5z1OZlOrKdB8+OPUj1SeC
CqnZ+LbD1bMavvAaxhR+o3mVrk1q6x8iIRmH9/yxiP3WfPhHfYCBbTda0EU0JF8h
RlEoqxmtIci/IPSm9X2gwpGUsqLr+E8ntpSkxT8pVkzJyd0wzbu6FJ/+2jIZqD3M
8deRf+Jb6yKAuB9z4i+7GgxPzHgkxHlqWP9HB6V5GYGQRvUuptukUwytn1kIQYuc
jwNuxis+x89Uh5X4q3Hz9oyvudsEBB3jwISwP1AFewc4c2VEQSxX903avi0V6jg9
vPEFgb/ue2GHR5Jsdjklr4Of7wUzXRXtRPBatLz4C0hhneWNDNjnZNt3fnn4vePs
iPJD8xXXzMomu1C8Yd68G6KU6tE6BGWUOjkN7fr873jgSZ+KDlqrLVvXg7zX64CO
Xic+n6FkXNjhsyD55Va9P2ys/r62dEFePfOk1nI4w4GwFlMtTxrzOS3k4SB4XpeJ
8HvsBR2wAETfphpwMNzovgbr9ZCq0UREbUaFcT7LuLYKofEI8PhQGvt1FzvZxoR3
BUEbOhw738IFddor5QP5RPTM03XuRfm/BBnWlW/DWYDN9hmHJrPH+HA5W+cro5Wn
twaEycKbj8+H2UQ83DC6BIoTbl4/r4soeWWVYTjuR/MCPtxNm56r0blWGWCqpIug
BsMKNYQJkwNmRY25svBIfUQos1eH2iwPl1MhVSUQMsflLHV2hzGvxZpSb05ny+CT
oCgzmZi8WefoRt1bzHnbEZGjULryBx3V0+FST/IZKmlXe1U/IvsuPdFGo2ajX3t3
N3NaeFCw2dRIuzUorUAjNWAt+XkoCrIG7JOlPypGTgl94uPoprnMGdKp3VeBb1jQ
NXt3M0iPxjAby5BxEc8aGR9aIRr9RMQwcKZfmEzsW9efSAosvmbvB+pSDQIBaj7J
OLJvafBDbL8twT56COpBJTdxME4LHrk34s2/H3Gs74Ax7tDVMjq+37cbmVDhCYaH
nGSYHRAQnswiovLHwl2KdUfyia9I6nO1wEaiFFGO8lPfWw7Inmj9QYFd83dkt18r
bnmzLzszMUJxytcM0WZH0p/soSNkGxDcHPmOr3RPZXBK52TIoX6gjyo66IO/rHOB
FMDLTE6oi8sZnr+HSM1YRy3b+c6nL74ZO6HhgFG4B3Zkmye0XRbbA18eKMN7ESQT
w+WriwCMem7jZPxCyY44EHWzhisGui1ZmLTHfWaX0ACFgselNtZIOH4q9iPMnfw9
fRIB99o2/cd2nI2+2hpUzSjLMCc/hk+HX9gu3ihbEA3jjZvsAl1ZT+ML3e/ymU37
vDOLJtkHtURVZQwuj1oWGoDZm5WVCFhITmHmAVdLz6O7nXYU2qJB9VsDBKkGZ+N1
eq2zGOghKXXkDrQDynNKF/ycKy7Gi6xYDw7Svhrt4LO7SJ1i9V9Iiu97A7BR80Pa
6i3y7wQ/qOz8kDdlosNUjfEryNK9E28K+UrS9gojP7g9+Alwqv9sjTVJRDOjXcZH
tlDrIU+pNKQxBdjxWO3RuigvxltdtIYOcxKcE1XpT9jR/NKN4R4Yn0bqGR/SGyqK
ysLY+hD7bDsQzJUqGXVKoitlom0WQ6jlLJHaO9lki4NV7Y+DsLdkQ2nbvI0Q7pQR
c7CP+j8z2hi787yddpZw67m9rXpSi2KCeXcmR/9bNNBab94YJX61EvXUv4vnZHk4
uNoQphynEGuEsRP7q3XcpARhPg20hY/9W67YCYftdsArZZmub3RccoQ9KqKeyWjc
rlV6RAtJChfh9p30nAjZP5849gNjlOUJ4c9vH1EcigNpHT1pNHPjXgXsvDrXqibG
VwfV/gw5XNhz9uDvoZsHIU9+4B9AhHcqzyog6LZf/LJIgV+HDZ9OPKWH+DIfX9Ps
/F8lIz9DqG35C2m14yPm4nvriI0sFMsFGEayltkKWnUz8ARwgqo0uXY0c9IrvtBX
mgpwoFB9qNciAk9WzMXRVlTMfZVAFzO1f7c6VR62Ie2NYFIDVpLxdkhESxQExYVT
zoqupKwvC9Eb18U8P8FHgg==
`protect END_PROTECTED
