`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BcC7AOdLS5Ho6G4dHLfrajn4iOg7yIAz6tpDaUXN2SDHlBWoxr2wm+MOm/tEY6XG
Gkc7xoeiMrYyIMQb6G4HqC9QudTpb18vwe1M+n3Ql9ClDZ3nFWP1NG2VBn++Z7F/
PFstG7MPt+lL7qTSekmaPBUL9LvB3bNu9QPCyvnG2uDt2wyDvnnxgnMybyjuUo/o
kE2Tc6BW6nLCmeJ/KsQuOPyZ91vXc2Jc5ADD5vT+76t8lWnhaujdQVSkRj6PVf0u
WL5xqdLQ21zASPjPRtv3RYfk/uKsK8oTxw5fa/EQpebbpOOCqzyshKdqcDyQ2Zac
5pP9/NzSIRdGVd+rsK4ha9Dy9amB7YJiGijZ1e+jZLp5hdm7sC2/njENJpfdx+Bb
6948S2cu1rpG1TN9ryIpNDYQeehwV4eORltuQkKKYoOPqUfe5MtusrRTaA7Xf6d9
QmillAfzZ6JqBBlXDJP4ei8CRdTAw1wGnYR5e28Yroo5IOvg7oFB8s5Srgs9C3oa
n2GJqF3ZutLBDF3L4ty6QV5uqZEo+Sd75/C028PfxuPb+zn3MWJrz8N0oyQOiuou
28UG/7OmOqhCvcA4k1NcRDtQS8pHcEj5BqYMsLmx/6c=
`protect END_PROTECTED
