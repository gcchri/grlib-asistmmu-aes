`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdsHOQfdQjUJVu9Uit/+e7JiTrvwQCeZXE7R/tjCDcuYgDSRfmci5h5sH2F+dgkW
3nm+I+0EdxHFXiEqmtPwrNOwL7/HLg+sK57OIDzXy32dWBEye3fk2qWn+m5KYbLQ
DyswUn/xDgu23RYaN5u2TyY5JpoNXU4SWfyuCFVC17rc0rJQlZYYR5cx4qeybVL0
IPaBg5/Vg5X+eSfGyuIW93an+5mdp701KIEF5WLHz4jUYMjWriVXL4vV/oJvCTUT
0LphdyJrCj6eUUEyNq6mtruGj/Qda2cR+1qiq50nzCXMhd0gJ5rccjpGs9TqK8f9
`protect END_PROTECTED
