`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bshjguWBkR9NxFrG1PpAjAvxglnvtw/Fu99VgWOvISo8SgcCcwQY3MBa8n5C0xSp
6g6ZNouMdYC1yJFDi15fA57VLmkDBTxWAx133EprVx0Hm7MIJmZ/1c0q1rTX6OdC
sRXxOh8Zwij7Mf5ahS9PQgOg2RFTJdIshp4AWwVvD3kKE6POg1e66cMqzJmfBUPh
z59RhxI2vS6jnNZYTQyEaTUqD7CcF1kb9KRtWqjrQzHMU0+8TlfFfL6pYKZJarLM
fsN8z0g6k7ZIso0eQz/+3zjOLrCbN2vIGYn1p+6UBII3MnTtT5KiBHJyIoGYefxz
7XFs+x45PAytyuX97Nu5hCf/ZabAzegkJ1OC+/F82dcgSg01fXJN/TtE5JKa1hjx
qplBffCtsuZIGXlnbLYa+R0+RtxxdrjSuDLT+xB32gPU6H9f2OpuJJYxrdOOaNWU
/PN5+ge1D1fZ6qMg/NF/NkZS1i5e3uZ6YdphePTilPIHjCwTk+kbvb40lg+/HeAl
R7GNhHurlYdensUDRYFilMjPJfU/y+t2ZVZtqtBWRPVJNIMWn+C9KHzarikzX082
2LCCAXbZwWJFRIKLJ4nmwwXVuZjtcVdq0twIE0xaB+xJF30C/i+MINSw6X1sjv4N
PTSKo3KMx7NWBnKAI+utNh4wdvq1Lz7ChhmEp9NtRQUU0EFRh+E6uGZUuciRF3NE
taKh9BhTPD5rpfkf66yr+mADWORvg9RnfpzPsTWuRh4zZW6yIVObP26G9mtTaS8q
yllLKF9c3w0bef+HPOKnfKpgaIC8t9J4cA03f1w17f0tFUTOkMlW1KrUwtjpMnIC
94cMucBkhihjJmFkmVhE0o5nTJilCc6PSEHQtuDD8OStRwIF/CdDJoSUPBdJxhzG
BM2Wn2CL51pMLtMVSnQ7TZOAFx/4VznpROGVy8ZQbaoYoxZ+qIy/Yi3Kl5vFL6JX
k7NYUIQYV65hnf1rNQTAMpLM+eM7SZFhtsihDLLQYYx6ACgEZhQJDKTeGFmmYnkL
3DfGgo/Q0ACkYBVXoQXfjNOjwgjRhineVZT76R5AToOL74cX+mIN0OYkvggNG+bU
SWUiECfFeXJbxPajhJJLyAIdur7B/wQikGU9+ICO0qxGZaQllVKbrP6RWeD4Vppk
wpIz2hZizuFaeD9UHNh4MrEql5+wjRqft8Ok8h3T697MzQsKFVHkUZUHdl9ZTvSf
6H/J0PfSaKnPEGw1N4pnQp/8kIBr5NPGZyThqtLCU28D0dBRFiSY6+rvu7AdehYD
PZEBtazclaP1fdMfyC/sDXpXLAEMcUch9yG5uEPpiMq7Ylc9KVYR/hkwM4v8lH1T
vWoHWbemBbFgyKEkOdiRrGue5RRhEgTtvXcbhJ+7/RL3qRc0DOatdd0reaq1Mzox
suufrw9rfPk6uacIE/Bgw6F59BbTDW2GYKmDq/LLn66PGcnro4w2b7fCvAYRot5g
0dR1VaHlyHPfZ+rY+jVYlKWl9scijbzhyg8ilM7tQDEimKl6bR4e7oXtXk3OWl4X
/WOo95iGNo/vhBNboFJUVQDiaM/zx15fRZXsdF/ofRAeAh9R9li32dI4ht4AEmGP
6CeAH0/1ASf1hOhQBEYtHNG7H2kEnIALDN/+OnaGLnwGXavhrVhk3VMKPWA20a0M
HqcWDU7fYPj58TIObwOgjzpFt6j9bpG45hK8Xc7HzGzfTYP6XoP4yMrMXj8BEiBZ
/A8/B+jzbMgjpH2bonBVJ69cx8RE4wIYBl2yFkCcYrFSdDzdjXo7AbuvvkzFUlCu
x7fa79QpoexNANs3FDBkrgYiYad76dr/HpvVnix/CMRul6a9a9yAn94obdB8j/6Q
9agjTi2bHnFLwpBkl8guLOA6dtSLJdXI/E+xLhzpDqocf0gJQvCviltjk7o9E8BV
P1bM/24gdORVlYE0Is+nbjF0ZWRpvN99BvIi8qyep0A3fjQC78yOaVXEvVZ5IyAr
SzcACDkrQhloDjnFPlt+JG7/ABDd2qWphzMB4gJZlQqvBkrDXjwspM+cEBpVXfrp
o6WnJzQcobQ005PRdN5fbUfEcHgiHXvBrepaaVr8JQfKj6zrZ3sKbCI3dN96od39
zy8uq+FYWXpzqWUIsY/Y0irQWBuOSChDClYVrwOSmA/wJ2+uJZ0TNLm3vi6ckBHK
lu/ec9ghTgzP71KKiiqcKsZy5oo3brZuCz3DTCNTqzzBs0BT+Y+0MYakidV2vQOd
HZ/xFmkwkq4C1Xm/hWG5jyrQ8LT9V//tSrXe2frXQdjsLTp9pH9TMQ9i2sxbKuog
TViekMdVJM7R/Ym1vjLCCU//lwDkiMc4gM8o05OH49jonqPL5ZMHy+O7WfI/WlUs
eG7hCVWAh2LpbnWStRsHG6Zz8ByNl1CVGlhivPqaRHTp5yLsjqCjB+wuFcNgMov1
5P6Io9QiXScOnqZCyam4/UsVJWM6deAxEeT4YRg2VHSKjKCoRfyF1XYUp3Dg5EZQ
Y6HRaACuI4DJCJ+Zuy1H+nBqQdgdg1t4ZFMH2UZjvW3xcQTnccS9htsx1HNU84Vu
80Mkb43iOgD5zQubb38ycVMM0sWfrMv/TIhwcsUby5MyVjybwgOslcvUgWiBEeHt
nQ3JrfKEYMFfEIxRxTlgbX9W9zpnnLlSnu1sB03h0Atqs8o0HbeLRdjkFTQCuTZ2
IN/BbWzLqMcHgPAOl2Cmr8L3miiPSMtNoLAWd/Jxh3a8FyTvvCUkeAx2D7/KOz/1
W7R3RGW7DoV9+1bvy8woxhSGkwCGEPcL8x3GsX4Eo/TxiS7knw+Iu1LPKzOnTO3I
Z5JTX7ipMmMhUm4qT6sTEkGYasSOThkVTTTw6mftJxjvRFymXBnIddsl0tFs3Bdl
MmAu1L2/39cIOsbBEsrgyBHgIISjkFdvTsKj5Vtb+p7ZjW3fngJHFWnuma7nHusA
2ePt+WAwGVQaC4ogGonQETVGnrGlE7NZBzwFl7tzzYvEa0BpeQNwuFainESPYgKF
w3THPkvg1xx2v5qIHTZmfov62rFpzMQcstJHICFFBIw5HAWEg5K78V4KpXku+XXC
ZHcD46eusM6hpJeYPqvYnPxLKOx4Rqanoo+HDmX64q9KtGHsPA9O74qXLyaNJx6i
pmWFnA3DZyCq6KG3TKhLzTL2cY2ILfR36fHdTAvVXOwEXFHot6V2EcABDQlmxdky
3AzDLYp6z+uF8NxYooD6YUO69+lMwmcVNdc+nw1B/+Q9N0QhwNOQOSAHOSpkLoxa
iaAs43F0/NrHgDrRN92pNYB2oJrIWSv7RLu+WZRCKnsd5SFOYosjo28HnzGv9lwO
m3PVnSPpdkavTdIj1shpnzSmCi40I8LByFO9GczVozq1o+01Qh+L3U5NS+OinipN
JWZ+wgsfDIsNoB0X9dt/oc07ihulER8psUZh5ynwwb70C1eFhBiGW0RqE9jR4LV6
eveOMNMs/WCPDDmGXRnMIbcSBJgfM7fhGN+tQikwyZA4KdG/GdI0S4izigK1i3Jk
t51ocSZhP+EiM23wpcwjt32sqCRk6VkSDgNG4OoRQg4hF53wH/TfwTSIDBYs89jX
wms7R87w8xj5RaIIT1zOPe90POKsXcHZIwRu5+3qOFcrnDvqEkb5Pvqc8yrEiZ8v
Noz1Ru8B92bf910aoHusFVwDWl4JvIgsPP4PSpvn4uup70kyxYiOJkdLpYAfN6V0
eliMThk1QANUl3y2fYvd//egRwGpIrP9EccHObpXG0ZzHcJZKA03vqcWtZjLmmsq
JJccETr/aGbgWbaiajPa2PINndflX2iL+IdjVVkGRqKvfQC7IUO90Uy3rsL7hCLc
+/+Mn3iNVainzHi1wPq956Wuy+7vVQrJuwD3a3xnMJGua1huHJHdodakFeIAZhVj
RtJOI/Dd/gEAQh9xChQqgulfV5EITyPbRemShl6bsR5y5/BbqomhTZELo2NJRBiv
jYSC3ttJsYPWoYyLPN9UZaEVZgQY5jBG4YGyZ1ZrKyDBiaSQ6yeuCe5WfN8lvzuG
OHPMDV3pk25vfJjOAovXEnGnaq4+7HHlY5zW4KErtLsHWJYz6Le16T74eM14uuow
8Vf37GT9fVl4UwBkO3bck4SWVvtkN8zHmiI0wNp8QiERbvjJkmQUpgpa0I7Tr1FY
Dxhdels4oSkOZu6PAhYWpuvtzngoInEEGQiT+0nCUgxAjkmW6ksuySnidUnO1LYy
cpTP5acoZP1zszPcHxcYq7fUgsQ7MBXnDdLt1TYh3XS+PRqxKIbuQiSDRMRFOu7P
DWyhMtnb/Ka3z63sT7H5FTAf5aF5UM9nqZYMZEIwVZOBD1AoDWflPZIx+h2weuQC
EPoYny0tWhHvDQc/Y1G4pCYuGIzV7sPNyHnKqIymRGsTSX+xCd3BcvG3WiS52JMP
X4lnHEBwsUvudHRBTZmOlWH56mVCaxBNKl7LpBMdJzA2TFAFWCtWHFv+GkgiGsZY
a950uKAXfj5p2Y9Ih/9f00OV4ffDhk0Y6/lVidqXb9eN6xz9yHeAbitaZllmWdJa
eLF1GgGOOJ2mTP7+1VZpQox4Ns79wBVnVkVnuksGUXsjXTAVg9EsW2lpzTuQbLIm
8s6eiHA5wW9CvqlFgnnRq1WeixDKBrkf2jAEzdYKxSnVgTAaSbsPcU15gEAlzFMG
0bgwXBZxkGzu49gPCG/q1rf+TO+mZ7n9PUU+0EIvIMWFWuJBYD9QB5mI/zhdPRSc
3fPDt1pBmhxY8jkQKN4BFhIGO5EuG0C6L7uSRf7ra7ImybobE0Pks1fSXqc3XVZz
KT8pg9F/q3E80w5iDWYN/LTGtBhDENdmrpZpqri6vwnFIKHfpGQdN3eWxbFGdJbG
fBRkaXvsHBP7YdYfGr96x2mPgSQh1L+EGnn6co55+WimSlysIQiOtZRRYoj6qKdh
FigGXdwQYWOhr7konTRwOW+1uai5AlFAFHPG69TrXyDV9GV5/eEUlNQf/UGC5eFx
1qX/l9ZqxITEhII3oEft3oeYSIAK3pgdnG81wAr/8s4poR90Zw5P9Rbndq0wZSKU
82nolcphcK6Es3PXDACJXtzARboSYqb9ovVvi3kiZ2drRkp5Z1Ruq4rvM8hFBr5z
Mh8OeKLk/vcaoYZFyJzQSgDCmmy2IbS1snzrI/zeLFYuHMdUtTPuyOrXJNak7Djp
248mS5Gv3MuF2Z0J6g4e4h9rEl4coyhGmtk2XeUukB6phMqoQM9BwBqkobyQjMzi
ZT8Yxb4nQ/kLqlgbVSASNqeU70KK5YKyizQKwPYs/2ydVexrYvDSnIQPLX2jHnFF
Ls33WZQYCwvR0WPYarcV+pAAdesTL2KT9vQRjKyx2gAMN5VVPsR7tdHyro4/8+6Q
PiTy/8G1WdGjnlZ8ClVI+NiHKqDee61BEReyjdkAV+YPWNY5HvL9iG38meJ8JcKJ
JrdoAC27/KXKdBRCpZYuOlMh8fL6wzpix+a5dFSzRtiBtrdSJ59Lp1/APRyx11Vc
ZENkkl95izvbGkiZnJ39UAPqYIqzZ2Djfrw9n/VKXKC9mQsyRoh2kWmM3p8IJnUO
HlkddcnEpnikP6nHVHrgqQ2AY9/BiaxoxagAlDyxwfqsLnhkyYmwZNHYZQgubAdY
pGRe+Nz5cgzSMo4WDJokbBEDq+q9velEfdaHLUCeaOAOoP8Im2bl3jXJYEMp0Ss+
wl1QE5mkXT1ekgML9g/vmeUH/hJpTVWTyrPBzxj+epoJghvF2JD4hKW1JBUpcFOe
6SkZ/r/ajhGujvadhtnthoxiwjBGo3ukmUF2QZwv3lWNSj+SJ6KTNZGvAjJL0kck
P9GCihUBpnXqj4WVEFVUrtkxIwKtRF4UMxnAUyqlwpe0bkrFQkziwpKNnVxdvc2J
Mc2VhzECZlfucPVUp4MSCe4l79FTc4r/CTx632gFtSpVmNnz1UyKnD2J6eJH2VRW
5VOujWFVPSZ0V/siAaP9znX0NK9K9RdaNbuDpTpVoieiEuknwHNb7tNma0B1jXLm
/oN8lic+VX0Lg0qrwck1yIRnn1JKj9RsBMJ0EQVpx8Fu6piPQABXITFKizbxf/yX
R4ROMlQzSEEUt4CEs4bviv9z7Jnz1frBbHKtWWQmymMgLBkM/Pcuo2vZ4uhl+tSb
/8U+P6KG/mAigeneY+FG2aB7Ks5X0S+83caw+ja/oZBWnzLH+JrWWptUjOaV3WAI
P2AzWgilxC2OXJFvJxK+2V/o6CF0DqqkLV5XkRPSsWWOqLV9ncmSdx1I+bX0TeWU
/7njFwbXc64ouaaEY0kH+dJ3ugTWbwdcySLDEQ/mzs3cBcY7NQFBvOPgtb+O9F6/
SJOWVSoW6ZZ3vsus/F6KLyOQiuE4lTWLcKiuhDsJPjyA3KYirc8PGllcQWAN712z
Jl7+wNgeiCxAOGZaLMyiw8Xa2CHdEaxawOwEb5I4/SgF2CkRsrwmjIbv9nDjLlka
SJSRWO2I0YBl3K8hN1FjbvmfCc+41zvngNB9Ekyd7+koDLcxMYc6tile29KZ4V68
mYl9uP706UdwLUrrDjA6GRd6VfqRJuxvHWtaXorFnYhfajT1a8CJYTv0GVSVIj6I
XstCiQkZM3q4Ecb3Q63V7xJTsohI/lSqwGSRG4l4wVVvMkyxzolAT/JnBBSLQvdJ
f1GMRDEn2eBMtx6GGXcAeeMJw53Zi94VrxeUSxxnNGLx/pDhHfn/abZomK2oZKDs
WVrRRXCjioGIuQRf9IcYDfxjv1aj8HFWHrEI1be3vROiEYTA8Jso+2oFlHtfNGA0
4ZX/0apjgrh8C7rAEoTOHATG8Rc3Xuqr/ideSHllWBVbIBXDga0rSlZwsUPMoJNx
jab4d4nwBNp/cUFtWu8wX8tFlCIvGK1oi0Zeut/RUjjYBtSNy6Q0X7C2KGCYIpSW
rfbbj3zhZkL3gmAqJHJ7kFFOPQlkRxIm2MJzkH9PADrygppmKL/m2wF9UQlWOPEp
XmogNWI41U+Fa8E6MPKPeNCbK6Rs31VKdFLF7Fv0MRK+JmDU8GGfKcLpcYUNv7uH
GuZkDxVydVu+188sfFT7XcyuBSmu3Lhp+qeZfmh/tA9SJ7JVRQrZRZZWATZztVZ7
BP8pcME1CiROZ5SvyFIgsc+YZbjFAXAdABOqg+SF/s40UY2FudtLdHuyxrmKX8Oo
tLrLw25rLbpwx9/GaEQXC+1mRKn2F4j0OPKn8YN/xDRlpP9xkQ7LB/WLdD+HpFy9
XEjhZ8Z/olkNNoJRASFjO9XrkdHG6oMD1DHVmX6wLojDjVix6EucqS5icIwgmoQm
h4fXadTcR9TCg3s5c5dxZLrgxbCsh//2Vdy869hP1iDpIchaqvySAVYrMwV5+ZPc
lYCiDK4StdfGv24S92LVaJgWObnqXQmY9wRM4oeOfNAura3CZdeEqNDJ8XRB8C/Z
0weg8K8wKZcxJEY9lzubE8AoZm5XfhNo3RFvSvUlWaxDtDiwcFk55VX+BD2xswbC
15+fnbSGw2/AAibaJP08jzX2XRU5K5NAmWiD6bElh42oLzdJK2B4aYabE28oudTN
t8fVhXR51en4UXvcfzrM9d0ixIdhEnmFOybWvyyQul8KSjj9IYGuY7sxro3FkNXn
je8zst5dG9V5El+jEb9Qb46QYCNfFxmOZUdtQfvYvnXzIBU4qJVjcziFMCKmduqd
y8uDQRp98i/9PZwgh866eOPAQmbGK9J+6U9nmBqwmQSfH8DveNrMLVEG9bcObFaE
XkVJ4nS1UBFosN+SHfswNk/LCvq18/OvBw0yBeJs2sYzRO+bfWIMqQdUAtNLiM4S
uFAIzL619xVKSV0zTwuoYIAFIAaPrRIoHIjj4Zjkw873WVVJMMBzJtiyYY+VN4CY
Cw9S9HcM8ITpwkLL3SIjy9K3udox5JbgLF0KbRzmLNxTRg27Y+auDan0ZiazuO4U
ObvcMp4k+fw+2ICIuoGTeOuU/4BD0kCppx98EM5av8of2SkoSUIs9nM0WnjQq3X/
v3CF+cWPMfmY9HaobH/opFd+FoW3MQnwUkZqSOJENFYjhOS+z2JNaBNqp9fRC1Hj
+lyzRRtTjpJnwGJ29Ts76GywhkiFiyxXV+y20fv5dJ4hJAHOhMqhkBJbFvDuGWYv
TH3yMYQdxxTeFxXz3Ci4nNmTGEKJlQiIZDe0esPvAeLSoiwFqfkcWgFoUhDyslbn
zi1YrXXitJii6jCB5cydMddIRd4028NRaGN5ASBimEa3fa8d0mXASuN6z5HkP/F1
W7JAXZqr2Nc7ZqO9Nk9RpbkqB1qREusCH6c9rxgKNJT2Aw7u1FB5WD0ciM3oMJza
XWWFL/zQQA4MNeabcajjor1Via2VVb/RgMiE7ACj7mL5BMU4O6jD7LCTF/+fyZ3s
++MosQfFSy0SjwUKA3EBwf1gaMegAQzejCXSn/g0rV+pcSFMfwPBoELTStPok2Fc
mKBITtkWmHqQs0H/DPSyYJiiZt6qL8FaijBAtrd1ViCs6X4DDO5ckScrZWO1GXn+
aNdbALzUribhPMlQoTv/GofW8QdK7ki3a8RyL3nB7oGoh8paYo5rnjcHrVgeGGau
IWQcL6oe8CW0bVzRLWvKZADrRTMi/wu45D1KOjlYGE3KdVPMD1DLGRxaQnpG1A4S
ecSZrjhzH6IhBX6lB6YbvKndAnDgs0egP05FxJEhBwlxetkaNk7cP0BwWqiQaGqb
ZvRwqKtl48hWDkWlDd7QDTm3lVDs5rSe4EJi7dmZlObPO+w5Tdc/UUVPifSSBEdg
prowmDIn7rHViXPd9Y9CABH+fXZdN56ZSKSjutqpMLEDZAtegj90ArL4KU1GgluS
9zUMt7pml65Sx4ZWRr1My9JX4DiVHyO05W2b0sR4S32txrBeZD0gH2aRmBJwQYCZ
FL5lYiujHsIDFp6ZBCI8Pwj3WYIWAzgOH2QJa3F7Eq6/xWBgyw10d8WmO4j9iDwV
AF2c9VGZESVXUJ1d5Pf9TX7olDO3Yk1zmM5kQyDq34/iPzXnTY/NwWRp2t8Yg4aJ
f3LlKqG2rWg0G+ZL1jC5A4BQ0SIUFX+CabIgiVZWzaaYEOF4hBe/YsVpGXM6QJjB
uNb6hG//DMaBc5a7x4mzGCcBhJ94gyHNtgdkvhelTZNRfLic+pR0p52iS+agGqon
d+All5jXX4DSPmm6QiIq0DVnOwW93dJ/P143IenQbdAo7vqIRfzPtuRebL6TClVe
YaYvSEh3e8GglakZqoFqkDZS5n9VxZLcSfmVC0cq9NGG4KhGgQ5nWDZMjTdyq/3w
TTlq9qXP2jL1LdRUuXFRtqxY6ZWXOewCawAsZSdc4i3CVgdVn4ZrOUvAh+dCwbp+
LxTeEF1r8UCgjBf+7mft16bz6/Qg+p72JmYD5ymnutMLfWe/P8Fmd8qxC1EK5xN4
vTu5vuzURXzVO7q5kCXj2LmOccya4CFo/OfUqORyzxONWeozoo7XEA1lQnecZRdW
ekrRsYEIKbAB67HCHy2k94HYLhRjUufLKmXvYWN/BRkvjsH8rrWPmD0BzfCs0oGs
TPSFV+PxP0GoFzLNLoFzy52go+Wh9ZP1s7qui6hldmxyUgX4sTQviJKtXUN7a7c1
EaMHtu6L/M55LfEwM0wawwnRjltcsVGTmoRePvAVnkgW38CvhG+fS1AiPjkuOBm9
O5zSZhiPoyJSZua8CJPuD0Ssqo5afj8L9+hkKVQ+cFTWbowVXxiZimEgWSUrH3Dh
NPIQo95Mu7YkdEIuvHas/AUki8pgwq3j6zTzGIJmwrqk6Qa6ZyuLuBwR2BO+466n
x10eNvOr61eo91D2RZdwXpkoYZs3IajBS+dKXXuMaKOocVg9+QEWxZefkZXw6gbG
sqBQ8WbnEpk6vxfb/BX8KvS0uLVEaCWwiMCyhkWN9bFDFHXxzMAueaiCCUG1/FL+
8lEQwW2gNVH7Z7lmKVEKwO+Te1bmH0kKdOZXHC02/avvDXSJ2HVWcvarBbH4DQ7Q
OlQzBH15iqn/AhRVi9aRbI4uxbT/SmaxxJVAcjQYx5j+uZAfgbcGJDtkqBr5i/Ww
XbtoIM8td1blPznNRw9FgyOVFARD49r79US+m3s0z7rAUKcp1G3S+tBqfAexTA2b
N3iMyZVPDKRQygJCuD/bDh883SDZwqUzGdG1zzsemlcAUy00MPAPMj4VwP3vC/ZB
DsOIULofHx2p3wy4iWwFmbw7QnsKz48KqxcV+HXPQn3oik5J4hH4jTJnTQn7YYAQ
MC2l29TCBqKPEhKolOWd+zu2xu+gtLqTmusHyDFuWc13EHkDk8ipXrDZEYPWaiMU
Q0ntsj+DUjZo21Wtmcguw5bKvjAtHElpFfJmO5KjmDw9OXsVFgP3oT0PZrZwxLvv
lzIn8JN9CUPAkh0UF7iYXiszG8WAkgQOnOlIRG9GM3Awea8NQeppkroCgxWF/rrp
TTlnv2vCd8m4YXH2Emv8LHtKGL/TZu77xLgJKfHIxY61vfTMvgbUkbuxUHEaH+Da
PittgRvLsWZ1esHKJOzcO3NaLl+uxQEtXjc9lE4LKryLaRr9BwXczQuCF5hFz6tT
4zzQrAStsDqj9ehe8AMQ0BADJSt8EyXThwtJi+SwMN2YK64zYTEJ85CLak5w6cNm
ZWwa4o0c+PRRKML/WGQyuTEEyw1D7sgiIvR1z1cl/i8cBwyNYk4gTmkuRlXqNX0y
uzal5veC8IRZU/9USCdP16rGFBfirpR+/nEJJm+4IIvcRamNEy2+qE3FBK8gmn1o
WIuXMpb0Dobtu+nFiEOlYHQExHxksLfC28fEKH7YkZD1XYB9Fc94GU9sGIKQrK4y
jbBy4LsDAWS7bLXUeDpUg5lzYNhDwY08sb8wqUkWQ3Hnwx/xIyjPoN73X6kT3T21
Ao+rc1XTfyHQd6ZYn3AhNFqIgJ7qzPE8F5D/hRVcNQRsEbBmcFghlUfRfNIYpWsE
B4rreWeIHTbyWkO2N+I4YtSeeR0psnfPAFb7vY1L3O5DqIEtILZ+kIT5QVYJJiD+
iVJfuZgZ1Mlyt8JPCCeNjOGgfqrxOyTa9yOPSTC3mvR0nGLTEZ2txysx2SCpVsob
b4Xo8EZsiG7XIaikPDB9nbxfmTtCDPA+VafvCZhbOhhj8WLEb1LU+5VVrZVlpZJK
4YitF43LEr/BMjBV3kMak0SmgaNEEB3ElrlldA/XUErXPC0tV8mAdahapOzbwPs1
ujuynmj3HwZE9VA6KTNM8a1PRJTEYE2KrnCAvZPQ4XKUDFsu6hsCzkRXuXnFwQBC
YwXU3Pn1+m4URp0H/6L28Uq0unfEdFFaItQTggAwoRUbnlOPhp1IxXqY2KCunLAr
C9PEU2RTBp4o0ElgKAxSuKga6ANXtzJxh3Y+QINpC5e/jf8LVI2ziVxH4nvPZzYM
575IKHe9lEiju5wTrYyUddAmMee0xzqU+Jyasor+jjw4h0rw1X7hMCXP9gXoK7Gd
oPkgrLHlR/IhsUT4w4NSDoGyEl6wkawKKyDh++ZEFN4/akKhgXfrmEdYgFb8p70d
YdX1Whz5thzMeS9ulmAr+og+a3TB02brtsBG6+GEDXbxX5wnwCAp7lnEMKWaHb/M
L9suqymnyiH0M4IiK3zFHDlVXsTYerldCptIEx1XT3gRB2KYx5SKw4O+3xQuFBb0
HUZYI9L6vnzNtoPl+vCgTtuefZz3yzorCP8y3y9hOSzkqalusj4aGnwiDcgfE7bw
ZB/54YIgAJ9ACgZ/9+L7eXDBdAsmkU4DQ4AHTlqcjNHxtFc8Z18/nek/qhVgAMbB
0Zqmuvi8Aw4a495LT2kyH2lLgMJTOI313hDpBBvHfRAxgakwMpK1GUJ6dOXjvdEb
u2IaJxFv0Iu2gLY4hYYJEA7Vb7Cl4CO5yQKnVArJ+bj4POVa7ZkO3GhH7K35tYWO
w8Z17PWiNe1jgc1pT7XbT9piqbOgxZuWZBoc6q4a16jUhyDFTKBdc+SNkYIShGM2
+6fvKJGhOdrZYos6oEVhMVZ4O8w7hkwEJnLvP1NXXEhjCzZQojcUYTrqIaMXzV2h
EdczI3pS5p6R0wxPJun1NfBneuA8BZMw9Vteef3uNROLfyomUr2D/fF7m3wSw2gt
H1oDSwb6nY49ewHEEnJpe+HvbY5GkYe+Ea8iqhC9llP9JEJePi/424OBp/30zNoS
rAaxIQAYWso2beyYHJdmRcU8sMaj4SY4a9heHJhyvMuJM1yXVEoX6JQT5228xrR8
iSE/cirPNI/ZTSv3ZAwikcQ+yfJ9orM2d4QIivQFaEUfWMB44j5aGEvYFctUbdM0
J2bOWHT5q6G53IdPYit6slwGcjPqHTe/+pDkSR8rqHc13DX7LZqTa8YEQ9Txng4v
08ALxM6MwbJ/j+lMvRxhStYHl+WQUndQua043S54eq+pqtpxxPqxjjVNtTeWCtlg
vpiTeZCLjz2/iyOnPMhpDrS00YXX2AFfMK6hZ1/KvNftmm9XzOIMh5wXRfhp0hoU
2u5CtA4OIK3ZY1RULSdAEjz1yYrpyEPCjLT88Ml+bdV0Ya3Bs3hUZKe9qWkZ4jDF
HplhrtfbmZ6zTeEC2PoUBOs1J6K4e4O/MTrQMl6vbqoRE63CtIHOx+F7D7jljorl
hOI9891ChLYbbAYbzk/GbvHO4jr8bSnUlTMQ934D09ZyuZyPp24XRorybVCP820B
+Rml+opHSoLK53JneafMKdHk9KKu/2gQXRMYz1cucYSMCLwwcF8Tf9OYv/6dE7jl
Djx1VXqFw4YpFiCGF4JEhETilVvmbMFgsK3Z6ZrZfY05xCvooZWurqqU6Qk0mA7/
3raYV8YB+dnxtq5sl6lmGXjabfk/trvIJvMcTKw6afIe9CsCuujABYwiHZoYAgTM
YrdT99taonDFfjjR6lOHcSbC3UFL51RcSPE1U+z8QNoOrd/ixox28sPZecRobR5v
SUJ+od2hHHeQI9gqedGK4LN/OhLh7ZYM8iyOwPNdsKlsLX8jOzfBlYdojDEHiJN+
JArIMECIAw/GWcDVEBygqdqpLxI646dJjmU5AYCcUGvnRL3PoNA4c0B16rz6LMsq
Wa9SwUzDDY0HozRxTbNKKSdj8EhYd9CwPlcwryGqtVwJ5pZ27I7R0NeaCHC59eTA
R8hWZ/NjHsZ5N9Juu6UVWDQio+LK8g3tKYn7fJ0zxwhJJGSEc0STE2FbKd5HwLLx
RFK/tWOHDcHHTXd1fTU2jtIsGddWHzP5xCbTfD/T8RVxlZNUYWCnni7bI0+JX85d
R7svwKhqe9S40NNQUbzkqHu5SdrSM34zz4je4XLzMoS46f1iHaFzX4V8897km3rX
dFAzMhP9vuQu1CkPl9TUJRR95N9A9J++q6ObZl+Or4DJWCtRSP0dHvEDuCEYBxvl
7CsNzj9PLTA7SSyyqixpcbZt+GqZBTXJzYPEUdOQi38znxga9CU7hZPBaNPUgRou
V2+FOzVZRMjnhqa1yiPkjX7d/hlwGmtcUHScQJif+Uz446qwric/e6/bSbpR873U
gYMsObUL3OjjMs/hAOQGq0CZdxozy+v97/5HG4nwYnu9n9ZioVlku6dLJi9XFrVy
LT/XWW9bGPdL+dzFDyBSsILkEAyNAyNxdYRf1/sYw2gZ/roomfqIxnYtU7Ohmr6m
hT+xSIjEunIQaW1gOBpyDtJ94mwiFfG2sG7oGBs3RBuWnuJs5XZ1kNJA66evAryR
Sx0uX65Tnk0RyXMvAbFk8KCozIrCKl9GgkXumf92gXrYbLX1a+LaLHrhfMRECxhW
bJ3N+xHYBwFXhxuViTlSrpkA6sWlUlXHJ/dexCJPr4ImQ94vb2fWIXz4faWCFE70
XhtMbvtSDgE/JSYK0yk9uXpw7RIYLY25XviIFIgl6a3GGKtlDVj760r5h41NUuQW
fJReRkeo8Ja0j46sWPvyCwbjITSnu5XWtAfID/l8XGsjT9qWJIu3rookvfJ3BSJd
BzLEMyGwTOrbEvrUei4ekVz1qDCFHBmnfVecTJBblfPK2wv0iVzjckvIo7wbYSI/
g0KXcbEaubHIyVAIA0DuVqXIj+KkrhAY/Kk3xQOloGqi5T9a2raDHYy5TPFa6OIq
MC1UykmtvI/k9FvogWNlxIfGyiC8S9UOq+WTpXkDiVCdyJr9WKk209XPvIt+MlPl
wBTtuD1aLDaEGwKtaQBehKEq3BBEvtUzO73yiZ3cbCOMX4m5hAcmHdedUuWmgbnl
Dku3Lu3LeBMYUj6mrhgfDHiMXEPtdF3BuJj7bgxaMtvjGRqYkPF1vyvBcSYj5+Uq
aYyMPg1wjaEcSinSNksTwBlkCGeNg4Icufqoi/nyUTIruzgXBgYWOe54cJa79hx6
+M4hyMcIa6ofSsnPxLp3ffeR9BRwypwTrJbnnZJTdZwHI9vQhVEXihslA3zF6Amt
DfoPA0HIESZrEjpN0EJAgCtbxBK+7/hKp8dklpabSRDP98aY5Ie6bUUCdzS/3ir5
d4bs4yv8FP6FnV9Z3uzMey0MUZ6zfXT8Ic9mykemidbPTD/+mgqCGjmV0sbj7mfM
Zhw7Qb+ySat9iaa74tjCq7qJJnE6FyABwuIL1br9xWyUOpeNnvq+7PjCblMQmCOC
mtgc2S1t5IOHAHp3L6AkGkKXUbgQPWeml2xY37T7ayHwI/mQ7jeYd9wP6jw1hOqN
wU9EmAJVAmOgw9/srQtCDN0EDuxvv1zE5JkoA/92PoTNRhX6P+6o/B/j8LrJIGBa
GALGWVtxtUvAEhzuo0XD2Qgr2DW7zNHpfaau6tYao8GQQDIFynQ44fNq1jG25MQz
jrttAuXYEQ1LOAh5Ldm/sL1EiRSLBHT9GrtME5g2RMh6YDKjvMeo9qQaujNtfq/z
dUwpTWVUKtXmPnSvWoRchP7Zi1B77VPMvEpLxIRnknSoigKslTM6ngbjyyp4wSMD
kUMnQuLHU9k7nxtPgLFPDRd+aVolwUtCCTEfe/vOMBYyeD4xxA2U+kLtbkNMj0Si
xq7eK0kx00Kh5gwYrzH3QwHfu4kGYfCSIPy/F2ocW5XCkpCW3yQfG4Bku5JvL5gV
xUNsHFfeGd1opl+erbZICvTmt2EAuP1b9TBaHe4V3R6bjSzyxCOAuIVHElSULwiO
bf6AsG42H9sg6zwmLdEiPuYqoG5M735RqbVhbqKaOoIQhcrCX3iLEFJaizOP5yJu
FgxzFpj9Y6dkCQrxcsruV7MNztY/gg0Ib37q+/ZZdRx2RrOBbnWFn/b7hM5FNSaX
c9a7LfcER6MK5fNEJWgq8LMQZp0I4PddaJR+r1wwBsom+hPtuKa8v9x6JSP8vlt9
nTimlRMgLI/JLDeY40jHblkTNqRQgeGDFsKeYOFZLykI0dZoDzK/0xD0MbD/nl0H
YRY3fILPM9+7+AO5yvk0MOd+CamjeubUmspKCs9Mrc1CIKapO5tIng6H864AGO5+
BbP2BCddSAPWLmjuELJR4neItqGQ2Eo1/aX+7JZGbXNvPjL0vjxtH1usWINH4G2a
OSTeI1QGUaE6Dm3erlI1tPbsTtDnwcoz2VF6eS86tjudqGrghWh/ApkFsa9k51eS
6Wj0H8YhwmlF/ML1HE9cooe4PpV1E1zaauOsEr0+z+7BwdsvDe8JHfo2zDDQabAQ
NlUREDwYJdKXDzwUt/MsIPJNm3n8LRJI20/fsBcgFBGzuwep4XWTeKWL+9y1gx16
6ZBnZSh2+kW2z+naakocd9MG9wV3JKwhf9vJGcmzID0zJ1EwJLjSzpFw//EPsTX6
JZrK3IwiCj99ekJ2V3Vs3qEMtyHAmgyuHsQAoUA+K7+GSBUh8EKRErIlNRxRmL0z
GJ0RRZtF2S15Ow8M69vF716h+u2hCZN8HwOsnJP57Op4nwwfAofrFBRyRNVr4hIS
PCNToRgqH/S0rrvNIdlyGVq1rneV9851+dw/iNiidW5dShG+0YEQhz/7udNpjFhU
JdxFljXWQoRPYDm1OhNcrVYADvrphC40REQjOlK5SntLs3vXeA545kA4M5oicwDg
5P95Ac435qH4dvx+ZwmaJPkyEMpBaNx0QpwlGmXcqMgpQKfS7iltwByElh5nx1M2
Y0uo839JwTH+FQWbCwuPHYO94HOKuxVOyusA2Ndd89GcqUSlMYiLuAP7FecxEMpb
CUYHQxUp+P4R1KkMgNNe2qRb1MYuZxeqBtrUTcRb+lLjAMD3zlN5hF1wEazB94IO
5JryL+4uAbT+w4bTcXtjL0xtZNZgZ8CA2RH2cR+rcJGx3hdxZUu7irhFglyHwjPR
1hHuGh8O7LsI1LaYT/nT4Q8T8VVYT+Tx39FzPYLKXSNhXnFLCNO61udISmddcK+7
tUYuDXU4/OSZWt4UH54Ylw4FcD9VKwtQrzmtqeWZ85MYJYxUqVCLKVtGBV4AxFN4
wd29Vui2GWFjHtJ/gQzssXErhQvieNx8ZZ3VyJyHtfq9f/RciR2vB8iMHdJ7EfrU
/mNW/g9BIjyERvmHW7k57c+X4enagPqkcHQ4GNLfGwTWLvtMJ4M6DMFJ8x0BAkT/
FEeMMuOkC2Bltlaob73UblyGX6krqepacgHobUNXqeqvsXEPPjHuugOmi1UcVvVn
UUGn8nxo/dJLojGDJBPTOc5GwKDGYdISn2E49VgmPZ093xCCWBiaSDPlhhGTUdPn
D4qdLVP0qafQ/L93uLIDsIfThprGfs4CQwQ3yQ4P2w3Ny7dFgsebQbWHlub4KJSs
E77QuxxJq3EjTwnri03vQS5DTdNCvgykooLmSbqT66607C9oSGb2rxga/NaxOVwQ
rZLTUU3gVZV8KhRMFymrvbOjC6UjwN8FPyQmVtaq/M/y1zI3O3IKk6XA17r0Y1zE
Y86pKFX0UCljl9ijfQ1DXWwA8Kqu8iHdoHlefvHknnFm7vPu7iUmaHTNcHlHSlcF
qdntIqXPWXDnnXsKn0Js6ZR/EBnf2VkmwZqQz0RLxIV1g1DalxUIpmmgOBJCc4Qx
kTsTOF3/iJTgXMzPbs/Canvxk+FZ76FMk1+78n8iuJGbgvLs/1ccWPQbpHIDn2wd
NYkljEbgW1/HfTF7fCYKFR4Vk53vgg3Xzw63ots/wfEuMLzf/XzoeCLpUDNL78k1
LRkflc4eUg1n8JuzUiEkJBZZkk3k0FI7ys1QpamO3yS2lNeS2ewAjMVoovSYlCTF
nUNbTVJl1WMpxvXufSlsepeEuyJie9LAa9ug6pxi7HBgN0rygZhsRqpehgo8oRB4
O0YE9sjpXtBNuMIZCCbgkw5C1xbBagHe8A/gb6/G0bxVgZ8S96dmJ08/5K1VnXXW
eDdZ2yuXl468bnWNgp9ihV4ve0zHRbhHhn77czS5v1pS8nXMzggTWuG4iWwl8s/P
SEeLqexf3btn8aswBmBzLV4t6Y3SxQtK8ofDQTPz7dSy9zaDxqG7h/2LcNcDEb/V
UFzkIOYqZx/1AF4Wwpniru3Y5K5ll+aHC+Akn0c4oi0SNbJay2BdRjLdgSY5ysl4
WVQRNpcx/g6/cRjfYTGJ5n5PWTXKSrBNv3j1OjMlFp7hKwdAmpVljp1YNp9bv6WK
HoGtEJsqC13W2N+Tb+iLDfXPVS1FIhFodC3arHkmyU1ZS1zkzzucBuQ08zl2uPK6
QXo38JG18Uj5vUnZZBRpWsARo43/y1B+fXBjgptM3v+TNIGcSgW4sPDFAuF5r8q+
CNB0KKCJCubMQjEB6AibJpa3U9wA31zrWAU878rP3bkR0LOpt1dOofjFF0z3CgJo
cIUKkMB92G5q2VNxjSVtCZJ5zzx9qGsGUUET0wX8YTSyJ/C4uXFjwaxKgu9FYsYu
/He4gTjHaqFFA/PTHeWLavb/qs5yuKVpwMraDeilEwGLP/viQR+F2ETAQ/Rk0Znh
cTI/YYw3QCD4UiRzT3WyYY3ndbgFbQ6zJ27Z4dlg51zkncz0a8j+Cr8yAtoak3py
TkprzNr3Vu/v4qBJjB3WeFbQPjBDUKKkO6oAR/cW9yiuDzyId8wBgdMAa6yLyQkl
4sruob8tVf/bErujPbMl/xNoROpkHO9uAY1HF3HHmDPkUtPFuyAU/zf8vxtk/Hpl
9E6t2JtiwrQyjpslSk0MbfC6f3UPKXv9ZsXhSXFwtbMiCraHBMMSF5hI3qB5Orc4
zXV2GUmRudQrf4ls+An5AddbDhGu3EE2l4Ci4MX5QOiiVTTj8L6puoa7x+bldpWq
qyfFZpsn8KBeXxX7kZx/vMIsHoLv1JS2m/L1LpMD19ppt1q2Jl8UVWCfqTdmCuRq
VD+LH7r26ZmeymRhWtSUf64t2Nvi5dfFJ/RUT6I5DFhiok68Rx61QLxDqPc/x6n5
zvXP4WW15rOpDvqKLj4JeDGCWjPpoCY0xqxabrmj+e41+jV72BdnF4ttGpuP5iZ9
kCBscieEFEj4VArZ/MGhUh4I2a/5eISs+GpVNyr8jplMGsYtpAwMBjygDhWxROoi
nGjFNQLMQrrEw+kppUOD7RUf4jIP8BsxZoGTwg4OHUT+xw4i/MdZJbO+qDmoUxTV
oso/iVrGcRtMR/uFlS8U69nMlAHlPqjteo48OOl6DQHz0AnbUy5OxAsSXX9NaaUv
Pox3GpGYifDdbEV4umycKNX6Yfo/Ol0pqwIbQ1GhNDCy0OIMwxO2koghQy8Mu5OD
pZBzD0aJP/2MvWgV/SZLD5NepoHe2n2v5AUkVXTMq2I8hzEhCqL3kNrw3A4v6RuG
KCq9o/ud6m2CQZr6p+BxmS+tImSguzDDZ/eQLnxsbolyKxllucD4QoQ67tvnsUFE
cSUwzSlO0c53EsNT4YqiNtpIVUzeMJj7rwW33rORmU9Kp3wyBV5UTGqFZ7bSdGlB
zEvQqj+IwB8NwmsHyJpUH770d8+cRl0WCSDsAhekiDvB+65FwbZk9/XbduMQslXo
HaduHGtJqyvP0JpJBVGncU6kmkrrOOCF0CgGPnHUUEHMTrRIZnt4YUQ3w4U5KawJ
5crsJBHjrWsHx9RtG4Wh4RTfo/sB+LP3j/8iILWKmPCZPSEQldGAWSCW4Vd8F4/b
A3yM9HPjFb2Pg+MZ7nzHbcjtyXS8vAEtnP4grdv6sUEKu4P+ZdhZS4ojwiotR+Iq
5w2NFajTXoOLBDl/AHzlKjqn1C+kndnrVrpTUeqC0f0laGhG5p7ZZ8vxHTLOUD6w
/h+9DDoqhPMNsDx4t7VRqSQpywZjVQXmJq60ME0yinekNO8vhLmadjYyC81g6t3+
XvwZoEL4Mn406KfEX6Cd+bJDNtDHFfnhbxb4nhVbH8/1awlcOQgnv4Qg5kS8W8Uh
/FkLIRv29NEEURqeN2o/e+d4ILEO4Xsn5i6+uB9MBtYO7hBxgb6jDA8eHV2rYqhg
vG2mdCIaIj7ezDGQHMvXZ4H9a9Nsf2oyJ9IjeuTtBHqDc0RQyrAODG5lDj1Q0rOT
tF8M1krZL19PJ2YleVSE+3FLxGjWZRoFxqwSjRUrj1l9df+rxEt72TY4np8wOcjb
bge+ZYpIlb1dM/08/SzcstmCATVjq4mmRgSN98vPY9wiO6vwdC2Dy+03uQKJdUIT
/007bDj9blzOif3GBJM++r3ZsKPg6V1q3qlDs9+QNZJebKrKDjQN6orG+27REOV+
qcRi4GI4WU0o+T4ftz+SZbMTQNzqy2LGJFAsLQvQyMNGaYeifft8zZ7tBM6TRZlh
0aaW2GQCMj0+jzKEDJO+hJaehB+plWxf4NiwLLQimbLk9IlcrzHpmnuRXyFeOGRv
JteSD+x1okyCX2+gN5Wqkg0jShTyh9BfrO4yaf94ULFLdPj8i79hiKi9FMOwqPGh
babLT5bOtVqP+F5qxZh+C32fOCHTyimNb3Sli17MWmIy6c/GN0cm2wawyXZ+95yx
eFb/pPEY8C1VncA+g1h86Z0pGoTLOdAt3YjgQU1I9ZxMh3b4t5P0AS6Cv9xVRQ4i
sziYBAV/NdqAkROGg5NhCZaqroREiF6e3EK/3xiBEpzNmEqsN7lPBLRVYQ/ptKLM
AfGGveOzaBzC/fJUqBoEsqLXJtrsPdJlEFXKs4ysT250KBut8aXDS08FiXZO6FVt
cfgj/UaKB+miq88xGHHzr0nBJBrNxW75sY/yYUAWzggwvjAEUVLCP4uXLVWVwisM
1vDpSqyZVbr/z6jrpk6UqhHnb0M+/8A6vZAT+PFpLxC5p73OAmXeFjOE0IbQcopt
psd12bcrcD/ewFrA1URrSIppLie4f9cs5nHaoMGcJZIhvEknr+/fp/mM5FQ4TMg2
1QFhisvvjhAQ6wPtxKY13JeEAjSsZhJVn1aXZicbaPYpQNzobKI5M9ooKDMK5nvP
Ai7wjGx0E6SZ8XcjuvauHfjBpVk6l1xWztWjW/XC1WriNWqeiQAkyzQ3DDbd3D3Q
R7sPSqkl75fubJBSjmBtHOopvsWo/ykClKxThnBD3H82Z+o+YHdGNTvVWtsNQDNU
d2KzMDB3YGl6IY5QGbgoo3PqedQ9NMkOx4Q7fDrvWAsXjFi5UDkIdd7KsaObUvJh
2q9gnMYKIwqLwKmqQdOl9fOWR8asMqzSX6G0ya9p14faNK1sobMf2XFQHCpzG3/m
sZ+ZApsc7Z49/jLnviyBSHbUiKVg11fcxjGT6SU6XlwLqH3e6B0+FpHIJvOX9xN4
iF8AG6ZXPexJIDAzewWSi4dI9/yRNDBQn6XKdWQdxJs0NGXu3V926dHZkmdXFxzq
kfUYTHIE/pmT2t+8ogQsynmDO6Nk8gkAT2uerYLv9rFj34ttoGOd9zr/esBxT/7R
kA0xeLUw/tBXR9e1DpJnIGiQwsF5oeV4QOZiK4ZOEYi07qeYHmcW4GjeJz6qW0ai
9ee0oYKg1fphsRPdUgZ7shwd7H7tTRsTH2KrBPtlatBtgXhl9k7R6gR9mhuk8AmR
vM8243EOtMPjnZmB2ckY6Zf+jcekioRZKZtfN9WFD9s8hJuGXG5GPVdEHoLmcsJp
1XyIo6+6mOpmZd7+0iEsaqHAQPYaObt6fbyTXuTDtuaYmimUjj8wGrzU7o9HgHTL
mTSVR7AQMLiAkLZF8fGlsv6FV5Pkp9iDDonDr3bAgWaqU3DoPm/kv+903wdK1/ui
4paRUQeaHnAoh9SN2wkZ0SW9xjQYg0lrwLTX6Umc+1g1D+wzzND4qQ5IzJ0iwrhk
aFwIIp3EV65e1YvlmZH9oA9GvjY67oUdEaenx/csl+PLKA8VreTpdq9ArrMsI/k3
d/q6G0cb8x3j7fhg3UCszP5pyBobn0sQKKZBXFu1+dFgzVnwPkSz+P43n7JPaOET
eL5uEOsilq+m65jLAhEUDSIJe41ouEe354amsTttDzxPVTIJcxzUZHcEjXnPgPrU
cbRVwxAcrLQt1Ruz7+vG3voVsX+HoR2pnHVYOHvRRLG4OqLikmTZRuaPUxXvjLSD
WTU3M9cWJ8DG/mGxbeqS+6Odacuwhcgy2BNT/WSukMzd20RtXh2XHvTA1wEMi6B4
druOcOOhOoIkNhMLWazR6cq1SZJpkbqeXgqbeoem8v3JWKkZzYWXV/SmqzRxASLj
HQT+lZ1GlIMn/gEshoesTBnTWNKx4cjqGBfUcyoSHYs0FooT5PRCBnJ2QYiU3GRW
7OpwYUyzoXUvuw682lxJemrJZBEhu/pCamGFM0sPvZHiaJF0AIg6WQsUeKsVkCXy
3zvifZSg/sBn/BKEERqw0ZRIWI6rTxQRUhLyob0qbR+nM3dRvPOuTycQW8fCbLAN
1bysZFIzFa5sEFkh1Boc86xDaf9QhrjMuKZsoIyEFr7MvVy8B93tCBmzClG5qW8J
QHjHxIX7eEJ1T8h/ia3BfiYxTYhho2NnzuaoTgTBeKnq8sLzg8lo6Rs4UIKUY/dr
e5u8g1xZV1xQGKzd9OkWFMuo0zZXphapdWiF5YobjtiubnzIt6/lxlZs0KxcTo37
pBrJrMgj4arQmxIYpuArf/ASYQWxGtLISOjUAUyxrys0TKd/of/zIBnoK89ZPZK/
t3qyR30GiXHtwKJLu431NK+B2GWLag5xbkGAXFjRU3OJfzMvHbC7gYL4z80g01C5
KFI+rNFLOdqxYnx5qCenhIOm+QdLUcD6YCRkpg+wFjeh71Rnb9wMFhAEywRdm9eY
/cinp3Vuw0uYnsQxcMMOheU3a0OsW52SXquxAYucBlwMY/+RjOr1ScJv+cbSzWak
nLRDrlukbJGm6MQexSeNyf4oSiql0WXXAe8xVhaMLN6LXEBzwNw23sidcjpEcOQJ
xKgzzadionEqNEtNTIsm4kAYChlU2F4cOWbI1Voo1j7MLC9JWWvibFixdAPL3ZIl
SSnZIgmgnQkMD9RALZ+FUhxgnr7nMHd7jNv0mqRHL0vvaAoXwmOUCrL4//64cJZL
OyRcFdl2SwYdtu/O9kj/9XFKzvBr9fHN3dXGqf8xhi3HUG7Gkk5+jW/5wMMTzSHu
twCJxzsYJ2xu9zGfPCDIwoNopVcD1mEKj5ZYlnwaH8Ah0cMvqsTbrTWItf4jiA74
3Q2wWhi8s9jXkQZw1srMGyhb8vPA3Xv57gA1wPZGeqqIQ7/YAjSYS4CMMT0FdvCr
B74mqrRSPP9BxMAqTkgfKduWiWsS0w4vZKzpqO24CUoP5Axg2EGUtKcU27YUFCZI
Fr3mGqEm82HrtlY79ef3OyXZkEJ8qn5CCXCjKQUp1ELUnyDXJjF1mj9JSTf8ZS33
ePiATXtWD6sEUXZCcntRItf1o3X4PeySU8Qrg3+BtcoFyhXcQc38BclSrBDdtP/m
mUj5TMCDcMTamqq/xQhDJByYwUYU2oNPPY3o3+zFVkrAJkyTQP9S2ioGmcAXfaSS
tKyCb4SeCTntjs9dOLaS1iB+0cy0L+RqLwk9sgxXr51m3iDcssMEGbcDA3/4mxT6
XI0yBSFipT/0EOVZp4aXEWOs1aOtScf/sYK8DZLHDHJ8EQF8PoSj8BUvil6ofu9I
Bjv29OTKLgypsBFseqdVMDO/Hxbv1bSADm3JcHbirvKko8Vev5ClLfGK27McvKzK
+uFH88Y8PoD5x0pPXAaE/xpF7+TQ/MB1CLGA+OmheNs0SZHOUINZqVGYuldUCPmQ
C6GT22B6uiaVCT/SQ1V7/jZ7yJe24hVsIV2Gsj/cqBCjqI9mwSK4JzSIwIwuejmD
eI05Jy1iaF0LbqPVG+FSotTjXyEL1LY6nx5LEJbqc0c0v9CIXjk0N/kghqGQ65tq
gekH+qnY002iItwlvzrPJTJvxxsBTnuZe44AU1UhGwP+gC3FTzbQ/IcZezUQa9P9
ZxiJPaK1JjswL3E+I1WbJe7f/kL6c95BpnUFaB4H8UT5oz/34PJ4OpmeEmhLITrz
1o1f/YPRvXwxM4vGGad0nevy6A4tY+YH8U3nG8HHMQENEVo09YrpMctsd6V1oMiJ
9Ml0E4N71HJOA13MBZ4ArGIyT46nvd9/b8h9aqvd5StBeTuS1Ui42X8b8wrT6e64
/4/uxBWxNgU6omEUr+XMsS571XeNINtJdzJPxJQqOAK5LL3KZjTQGJeGIVJlIrrq
QSTBKitg0JEcPJHZBvD3p3F2StJryLOPaHYhzWJ/yNXnDnvkDun6MifmhPNwywGh
LyH0BNe8R5mQeuYVJU63dPML+uyK6NpkN9p5ylQoHJ8ai+Qc927GNdqaWwWR6aCr
GiMwSfaNfL3DBSDTxu+AfvakhpF0yPI5EwUdm7PEa89yItzyjpcgi6jwmDwgUDXA
oI3abm5l0aghh+ADIb9vrXFRxDH9q1ehaKodMl9Hhp4/q9+mjN0oav2e1svndf5a
YfK2PNuSnBKB5dIa1RbMS+KHvHVRBE60KlRuaVUHQJfzO1XVWFskiyidLJWYD1Mp
UzYP42xD0vi45JNBD4/JkGqbxQ1/scpTTMQ9smtqzc2F8w8AYKX6RwqwnZW8ucNA
aq7B5IxI0xow4pR93T02DzXco1FZP2CKHmxPLIM0BZzklALewFnYC3NmdacoD9a+
fITQkq9FC7RMpy6JzDLbFiqHX2D/xaqLpyQL41ztr5urMzPrcw3gdfYO9U95tuKV
yx4V+rpNK44gXvXREwJzGPKSL8Rlt9G+q3H/Xs2aIM1hqpgQgzM1VmbwXbKsy134
G3jNZaXq8FrpOMWCwfYwLIETKfNsTaPnUo6L6upf6sfbyyp4jA0Li30hT0EHybMG
HIuDrtwkCjQ2VNZxS5BWpR7jiXplzxR6hfe0l6keNL+qExxwOMnp35Pb6l/2HmJn
1jbeA5FfcbaJQsDxToos4eQQ4A+PyHVUYYMZNcjLve37wjBt2sceGMqeigYT8epL
fagGTvDEQaQeUCX323uCyApGF1WfTdu3KEtCmU7CwFVxjmfwV20d9utHZimq0qiA
VdASItx5peISJuWTS5zqxneC6/M6ew07ODfWiMsv34GgcSjZUKuAN95BUtbQsEAZ
VInZUaY2RvdLBHKqBGP5BmC0gaQmrXhjr1Zq24tP+swHDYmmw3g1W9u2yCpZMBC6
sRgRqbzdvG4A99Rxi6QFZ9lAeNMZ896y71J0kfHMnjpt0muoLOJrYAMrqN5tcSAA
S0qb66OEKIfztsbMd/UhkMJsmik8idJT7jK2ZPY9eHUVvBgOgbDVH2aj3XiqMlQe
e75RnHhqi5OI1ekvRmZ6GacDqstWuUp3U4BM1o2VS308Opmn95XQmys7xcQEYosG
GEr6MQkTnon/dPYhI4CwSmnDBSnT1kiGqS4oBIPrsY5bZRztUxdljj5wqfVabuzl
4vTVz2rDWjb/5A9QHgcnZvP8H5fACWG7S/TRZvnHABoDRMXwGENCLT4RF+xqiMII
fIN9SKsuLHaPkClA+aqUYhhnRYAgIpzJH8gth9EOCR30H8WoQ0/xnHNx8OM3rOyv
ZOMNsrJbI+nronymcNle5vo10u24MPbF5xP6R60beCi/sGI0+oGRERcERt/gA4SU
oOJYC/ML7Ck7GPkg/wxGWGhQB6sCNRqoFBR+iKNLq8g57iIuQCY8IjkqFZiwCu5G
EEWLB1/hC+2ZBnVJt7WvkqU1c57sQ3Rp60uHhryRnceP/iX/JWELwTL129eMXdc5
apns8Ef0toVyeSFhlfexq2LeDhTPiKOjJ4aKpYprNqN/gvTQRPbdKcYv9DTTOP/9
dwXhq0v9UK3A3HindMu1hkKYkOrbhFmuBUOqmRZy13lBjJ+RSiVg7Nq8zBJqmmtX
f/KKRBJ+jhVzAn6fmVFhjoloEDLPEqQUo3/kwaB43HdmSpdvG84Z8Ea3ETzDonvW
py/2iXg4HoKvYs2CAalJqq1lE38s0z5Lzy2Y2M6xCkqpT6wbId+7+E2JwODsng5f
4W0xTZdls11539v9y2lEwaqCNchgrDjJsdq7jEc5yLChx/3N3izNuwVknQoO+3wK
da4K+muAD5jvNo4gnoqmw2mZaBzR0of6IzElSCWJNWBVZa5neyiQwBJdAD4FN0Ju
Ethz47HYLABjn0T3SzmfnLMeixdi6cZOhgLSmIE4blTcml1+0wXDFTgX3EQNszKI
gq53QhMWJsOsmAJeV207c0q9Jjm7C4ud2iCLRpaK6uKQdxlTdO9TZ2nuBluNMsnc
pGHHxMqIF/pgeZvcXE5xGQYPjeUpqrbOT8qFDVIas852hW0UyVgCHLLY+mDb/vAT
eXzq4yeQpTsZZ2BTSn0XD1q8R6Ld95YeDlygc5wCwMoEAfKZ5u5jlzCn435rdnnT
lQbv3RqbdB48+9jii0c72tN5WbpO0st3iQhs1bNr8tV92twyjQ6uZF+0bAK/FMDt
DlhoN//6bVcDyLVRxAnM7nqoB5lF4S1ky1MX3x7ZynJXkdiM+lz7kxqhsx5lcgJG
39qnRA8CgdjLsbtBo7pw2z0v/gqn/FY5RMGqkKPEHtU/UNdWWjuJ7NGf9kHRx9We
kgSXnqxpuVhmqZo/W/IT6oPa/KkUi24t7G79GJcurvjcRGEHG3DJFPVZ/K/BQQc/
NT2WqaA2/hasRqAS8uMZ5Dp8gtLGguIf72y/3M1rFzGnmuXSNtdOe7GpvzRlTHf8
ua9S7Dghl8/FYugGsq25ot4qMRXjBURxIu+6JoeFJQlvdLx02GhboqQiXAZk0IfY
TOAC3/4NEpO7tEc9POAjexb3+fxd0YZ0UhF1i5dNLSvBFeJJRWMJKZQjU+zOoFmm
/xu9Ie0hPLWFqvLqsvSQr/8JfArgWXDVfD1yB7PL2VHyQQHvJQyMeFjIsL9lDk1Q
t1JE4KBFkZPHO5lXx0BcewSob9waO8tmYvIjwIs2jl39gFve6QwjK5F1Wj2ufO8u
/L/udKPJL/u45rQKJ41VmAZKhH65OXeB2koTiEmAsLW6PbOBtsyOplAGTwSQRnZ0
Qg1QFBCCk9Pl45z5SXgZbN9aDdjsW5CC0szvxo3j7TQIZSZHyXS08b+C0KA1lwpE
/UXzElvHwpJ9tsaG+OLrLu596JDpe5F4UKtAvQ0YuPQXY6A0E6i68dT9C7SErAGe
2KJzOhiAstDNBFkpjBgdSQuCRD5YwdE9ip1MbW/IEHLy2UQ6mQE4hcr3utClGMSU
jiDujiUZwFclQpajguYQilK4zZ2QS4+PY43MivV9SHsF33+XH3YCL49YWRFtkQh6
h2Q4G2dKbhv+MdN3DLVZuqC6/CsFvfFTns1wTXle8I6m80bs1v0IrHmPrfKYju2t
MZUO/mYyyEQ7KN3eS79NcMFwYyFHD/6Z9jk0lSBCP3ZpjjiTF5WewM17fzrO/qx+
S25gOiP2wXAVG90PH9rLKYnWtLiKlhxZ5DJFtMRYW6M5OlES2qF6fcpCKsE9lUOg
OB4DGiSslqyx4y1eW40++yPnWvpAjQWP4wFRk75r9kZu6TJKrAnzzoZPOTwgm43S
cSMD9QTDZ2nWsmPYoY/edmadMfoXB+17uxhl8qNMeIXkNxG9X5KkBhhWgK23CQIA
z68wplxudhRVPtEoKm8xij314HVp6JuEslAP2uwXs90Halcds47MOZQlJPut2vce
RnjfDYLBygrbcYaCqFvp+BYwiwvjNelPnLsc7WUm2Kob32URl1PO4mEJwQvmyvm/
bX9cU34FS5YJq4ihhGBH5qXGdhUa7OmtrAhbVnupwWe1KZK15pP17UCGbYlumygb
rVo6aoV7hq9AKd9E6o4UyIgCi/U1/uKteQrJ6eFOlJzsbvIzXYUxD+cXk53zGKxs
HlGUlR6Hs/EGJvlOyiewE2mGSD9OLjK0Q3TWTpxDW1MIONexvheRyaTVe0shvabo
ww8ihN2iWlm8g/R6XAZ3NcNvIIyGJhxbdaKS+7gRHXTeQxH5lIGfpyzqaAickflu
vbdRTE+7UNKYtwSqOg95G7YC+CVe2CLE9TVutqn6O6cd6LPerLm24VnUwZp4WW4k
nU3lJAbnBS3jCzcmJPJKfCawRJiYd5wJDaPWtS/CTwDZ+cOv2tJAkaZzHOz2it4E
z/EfRActYCgsGfJxEhV8I+TsXSX8pEmqgE5fic3OkXWbQUCyT9Al6JMQeySZVs50
p8J0X7zcFeYp/zKVlLNiu+azI/CAL5kiA5mkN7jyhKTR0W7LCvuskJCI33SZZgZK
emyDFHaL/0kNyhzDePCdGOtyj0tM2sMqsGaqBq6XCEKEk+CSjmVUwJsDdBNsayGd
iKV9xcG+yogTABdbdNiS1Bd3iSzAhNderqvsEpq8DMBuub1KMjLFOaKuYqHRA9aI
FhlIdkeJSQQhpM31wz9YInRVQ+gDuD9kul8SfdtICu+DxZnaPjnqEuLSZfVEjY8B
0I3OUE1Mrvvll34v+vPkAm0Uu3rXpylCsLuW18eEpE4lN17g3ce7WQGqVTj1hDZN
+mbpM4h4B1Kq7Xfqe+x6zc0Z3xR7WPHYRgGZT/K9My90l+I/U5ZYzvA+iMbWNl8t
vQMF6b8UCKXrPcTicoUNADBgsMkwZ9+oYy/J4Jate1iFAJA4vjPX2alF8GlRjjvc
+hoqCIYmcbeB7nM/IshJ57R4uLCBYO24v04ldTlpf4lwQ6olGZ/UILBTk4OL3yxw
2PdkTBrbVU+/nZ+Zzi4RELeIm/BixIXRmtIsUQGjycc5dy6D4Vz/Iom4166ZPqKd
Bx0MkX6KMxrpV/Tznal/JeCikYEhyctrgLh4wDg/+l80nzLqJ5NVCtmUDVL+I6RM
V+dUhZMF0gzAGNEY1xCUoXgKpSDc0/r2cWIytpJKZxKtcHe6tNp+8VwPEOO+wHjM
gevVuRewoGG5xCj7tbL3hoIe+qGxlSbDem9Fux3/2AhvwsWOziH7QU9p/oz3zEuS
MuNRVQdAm2BWx7nYP6JgnTNp86NoANkaNJ2cN/y8tppn1NutvG3Sb0Atf/DOso0T
8Hoo7qDOl7dkfYajr2ryfhVrvNQ5LwlRn0150AkJUesJTx3MMdxuERJZrOUtYScC
g9qtGBjZ4IUx/tnzh04SL+CaZW809NBAWoFYHXoGnFq5qbl12QUYGccYwMSCkjye
WhUTyTraiWPhRwM8neJxeXp5F84dgXqT7pLbzJXtMxZ50DwA1xr64qFX9GkA9aw5
Iw/QweCAIiKG59Y6JEqnTFqKDpclQybinqKAsVPIm4I6gpSeFKLWJDy7AantpOfs
tRWXg6IMD8OJ22bMYPz1DCjiD59VbfhjSpmlX56SZ1+vjVNH7O+mQnz7aseprET1
SzkPNyyDtKc5FrXaHzNx17ylr7H8P//KUnzbpe50RazhUgY6BwESSW0T5FkY+7xl
ZoXRP9deVYKJWITJBwfzndTEEYZPkETbS1GlsEFWnNJAn7AnABXDHkqajvDNLk/D
1cM3LPMLsFZvU5tB7F4KXL6ATw+v47jU9u+fS0wFZELuvxtfkwGibLJfnnEN64AT
O8lVvlN+gl4X91rMWLTKKa3ib3Fl59/ipL2IwgwdZfV12velqJb1uTE4yV6hSWgk
sUDVvHTTsGpprrSvT/9xCPZQXJTPx0lawXN68Km9xqyaiQCZu8+l2QaPqbF1nQok
JYJAKMsd7kk2YJVRH4HbZ0SWTK0oRlQv3tRREoZZFbUmWFb74SbHq2dLSPXgxEYr
GDFSQofRdcRbmXLmrPHSZSS1COBi0mm+K5MXxvv4HMkOo3HUNYHQWoyOM7tDGTHF
vj1L/TdZnAq/SJWxI1igKk38oCPNCbpFtH14TBVWPrhzCP401Lr16n/CIJwXn9Rt
IVIj7CxjFKkFX1akRsWBBvaPMXxhjrAw+7zRgtORv64IF0jGOvTzmCgLfwsVE+r5
BgQSskTP1lP/wvo8Sy9hxchlwFt8Z8u0a+GgbW9g+T2k1JmEHFAU+o4/zOgnB7vh
glSlfatsOhk9/kwcdxb0F7/xo4jkPv0PtcTud4it4TDbXzwPHDwtlHwszyWK887W
KZMC+dwUOPK+aAqN/sINRo9eAt20Yy7nOsi8pO5FBOOsc2lP+3WRKVwJYTG++JFN
EgNVxTDNgUeeOIvTwEXO/qgcNtDVTYjHrMVfIWqayXOf/YkJN9P7krnwVPKmzKAL
ZlmXTH3g9W6r2FryHQQ7dAuE+V4o7hNpf09eo4YTOEicJ+fdiEqt4piABxOMO5Sb
xJxrg01Jw3m3PTxnHpMGIcq3gNvMKqhKvP35JjvbIG44brxiQbIJfaob8MQJuhqz
jNlLJRg6ELVOWwPN2k6rJWsxgVGUQlGvAenVZeNH5F+rfaIQtlgAi+0CB8g+G6e3
A4Ffp6DOo2SY67a0nm8fNDqMlUyYiA0U1G1T3lf7YTFafH3vit+f3//mNHuOul7u
Dwr9Od8gel5tjeDhU632Y9u2YveAUzgBNB75AOfC+eVa82CNxTTg3UW4uwo3pUN/
qBJl09Mu1XavvRbgExcv4CWjvSQV2RbfZeyJlAwjBB+Anre1x+2yGJ8i5m4byLTZ
S1r1+LkfFWMsbg52lvlo5FFtEwLhRprmdsvZDYPBJSpFfhfxxxgZVA+jDHKbqgV4
ro5xZFSHdA/quATFaiLdTLI/VOH9WcDK9ylvfuXTzl8YzNXKQfuxxu1R3moddIWq
WuiCfmHN3kMRmC64qsV2eC+qqTw9KpmF0axHdI88uY4dJUxJ14Lm9nFEclg7+/Vb
ulpHigBc+VDF5ouYeuNXNvkQDk/djc+mygq/FC0VK4Q/yHGNj6N/r9vOmEbTO2jw
pVpo/gunqU6Lj5YJgTOmzUR+iiwNyREnYwjDJ5LOPDb8YJGHGbAMLvMef6lA1v3y
DZX+DGcB7UCR5qMMyCpcGFhnIRiGOVJP5iOkHF7ZoreKlrU7+F+oEDv7IaL5UN3j
h8iDXGOgyaP8u0hr3FTpZe9xmFgNUTb3wI7HBPpom4JHAp5pJYT+OECwLneTDlCQ
aieXmKuf6EbjNCLYScxrYiNRdy1dgkNJvGg86FiKIFZq3eSChQB45HNWZ+cuurOI
rM+RGsJj9rKKmE3l6VfQjTcGx75trUb/I0xGDOlkUlrrWKk19/sNYEmLNRvjnk4t
udsBlc+vnRY3uTNMWRPEMySOE9woC1Q1EhxfxOpqDvIcoEBII9K1a77H0NMeEWbO
TTUhojXVyBpNiI4bGr0aq3ZDV1IfON/FgNEp89Eo17nAl7gkoI+vgs983gJJNcHy
d0ODfxQmVz+d3U+cvagxiCZCn2iX3XeTnrzZm39tCS5Lm9i4YnqfDuBGllIL3TgK
h4c1BRsA9QVz7SU7CLYMuLIqVPFq65OUPW58mqixSGRVJ6J1i1taV8B1sCAZQ+5m
+PT84+da7hvz+7rPrPZQSdU/o8rmWnM88p32XJmtrK2DQq3xg2FIdQxRFYDmYOc3
S2FcHMb+q2C5gu58eGY3bEnFEVZ2vpjzMmtJshmiYYNBl2FqVO2p313X8UBWGRqi
GCdHrHflV/0w0VC+JDUQ4fRMSEbsGNQr4ECgSMwED/OxDVLJwxVBi9pgnxLrwkYA
fMVxWYXpr2DHh9lJyl9+Rm2Ibf1jXIBKKC0zaMvDPyig6qoKDu1Dykw9Rv1usqpS
/35i/sS0zr6QmhrRKuxBcEy98MEg0pYEngkB4VVQiGSYNbrV0QYexfrb8CgBKeOO
uxu8iFL01v7FlR+s48NCrKFYwfY+MnL/GXMMrUTFqrsp/+r/yoBxitTZfpFuorFV
vISnmQJazGGXLpI85s2/3CacVGrYEIF1qfZIw4Nd7TzxEtikKQ3nBBpfLeujRXdo
iRulbU46o6v9b1So+Fvp25ilDqiXQBexPAY6nsS96RjMeF90K+iIu7K61oRLBoFA
4VzyqecB61NFcqpQfx5VA33mCe5ZpbgLKT35oxL8sqG/pD0Ig7e3vLCocLLPsE1i
rAeN7h3lexiuCbsT+1+kkwj0F1I8qPPlohPQHcaYMK1TAXguI3gP3jiepSHp9klr
jrM7aKl+s9zJOAIBI0e5fA9JAuWsrMp69usBCBzXpv/pCbUh6nIgvJY2GTuAzeJd
ULQ1PV7R5afe1s/xGWiS3OjyupAZvfMj18EyqIIdHNOQB6/MpFGEdjSHv8brr1tE
9MxGGNHDfAZces44V/DCA4vz4cGyuvyDgcZRtZdTNVQ46Y/W/3rR4j0DLQlEk+uK
k2cCyxz+ACqAKeqQfF173+W+G+4YnF3bSW2eNpUhz3+p0f8EC6ES5FAPDwpNvYos
0DJylgQB8KN0b/fRW4HiVFhA9UHY3tGi0jZ1udqlOQttmuroDO1e9CsPior/P38s
H4j3oK60rfTsq4f3YigirE2LdsQruG5IlqsgyCw4i46myq01Hmi/DPAm+LcJxlJT
BgwDv/jtg/RDKi5Koy2uxXVL+UXhR44x68duVHsHTdcgm5jHawU4sHUKn94c5rB3
+Ej00HNiF6m7KPht8rhNJNKRqsYgqJABvuioo000pu8OwMk2NLZpojzByKXcV14P
Z5mlIxgYy0w3mI7WVlg6StV/55Fr8VbGlP6jvMbpYkAAo9oj01J1fuevYym+k9u2
Wb083o8A9veOEUUv/3dcc1oZ3CCpY1nXNYbopFU9vjFG6yd7/lmJ0dGATB+85TG4
QehYKXyzVaAF500Jo3EmRNR4QbQ8XxI6GYPyPCvB92B0KQFq2HSEx/ue46uR7Csc
7xfSSWb5MnxLDdFa189DTMFxzbAlyNtvvaeSuVnG+pZTI38UZwskS7spfX46D2my
RVsw10t4JVA5P6KgkhrlJARZX6r49zPj77FY/Fi4Avd36dakFLl1IYWiNI4bNoWv
9Ek//k3JLb+fiKoz32PJdMh9XGbNskXAAVu3+CNHzfmcggO1FZoIzmQ6VkdOKOVm
aOxSCtAqknmMZPZhMmYqjoHk2XBeqIJgxvOhm78UR9o9WcgPCvG1Um3b1HqSkIHI
ovxxEsap2E+QWd8+LEmNwL34JYE26mQV1PdQGAaHJ/GbjyulkfkdTiAGYvGm4ATw
d5t+/I7zxIua0ThcVWwyZNoja8vw1UjOyQ2ZEtucCmkjfc5LlMSKMBbN42VbkRwm
KaDmWaJLim4PEpt9AR2qze/ihn2GshZpEASyck/uIiLQetgqdH43js3DWem4sJwc
U3WmPB46BOhBkumRSXltrJN1Tlcn1s3SXo5s2wbY8tSUkIXaFnocRYYBXF1xw4i8
t2Oz3SwPYofZPTtcR4198QhYSEpzlnfOyem77JowU+tqbgyeJZzqkBCXwq0IQg8Z
Fm6ccHtL3sq6ha8KQ7kW67OIDpJtkYNJ8FdawI+P2IXo5+PDQPZFh//qs+gwPAGk
KdwSluvkYN7uKqDlcwNAKQYFzW7KMLT4pX39I0GAH7RJDfqsZYTSLckss6oYTcXJ
y7FXlQFWecl3lBrXW5m33SD9/VLQd8gGEGsbKQftzMFkqAeblDoblccY7NQMRcTa
2Lk/AGSBvkDOsCJKhPhXWQnCt9VR/APjzD660LJdRLqQlCdUejXIcxK8wmfhJUHP
JuO+5PoLrxCe+J79942tdaRH5wkEK+k/c8ZWqDuTY5PbT23Sf+nEOwclNeC5W31y
OsnLvZ9lYTKo7mIckzJiLs3cQqrplj1avIlp+pKy86TjI4qbYFu5Pd4CaGuA5XU+
UPneVf0uFyz64xl1SzfS8Oro44MvmhmOos98Inf9cz0mxneD9IWRcW02eFyGt343
Iqyo7mapLQlTRhO9F+nv/adrYgclApwzxF60ieZFt4B8OmJ1usGUBL5wk33xi4YB
/75NNXmGQHmKoeqt5OwJqkIHFtBBtA4AM8PReMOq66wk7dghcHCSLDHvGHgQ6LOO
CF7o2xvKc8a/LSoZ4dnEl8rstTqSiAVtyt4GFSQ5OZn2KOSYAUbOvybp0dN5loBO
zu/gHse+DMFiTkyIp3b7+bncYsCK+rsRHWftiXmzEgdMLAnKzukt3Qf5ZWfCsvQS
neOF/t5Fv/NmknUB0Fmb3b3d7lYHw+S+IT6ktwHCQvUoDtsRChYs+86qGA/Cb5RY
Qp5RM4UZ188gi9N6KKXh7ClqOPs/5rM8239j3TvXGCPFPMhbw3a3zZy4hcXnV7bd
vaYcVoLxuTRyyroYms244vCaD202zy/8Xfv1/fP/Y1khxltlH0lV1x5c/DML3XYJ
PrpRurzn0nfQ6ZGtFbVi1dpOirJ9RNIDqAH90c3f2LDPCOSsXt8Ore7oKcnBP+/u
rjePk2koBStE35baHWFhtIqsoG2pxWUMaUn1Yr4xKLlzhL/8KEhjLio/zJO7sGBI
D3VEj85KVJGSeLjLZS2oI4v7XVKWS9LaG6TI1gUet6K4ufRChMBe2SJvXeTzgqj+
hqbkK1q2hH2lZ48YnHqxSavlJamYb1yuaYiXmML58vWw5eTyaVTwQKZTvC6BnoJC
jKidzHwryCdoN+kxNckZ6KmVlw/yOAOHu4DljweMGN3cbELPbWVKU1gtpcjTrg+O
Ko2+0CHGFZ5M58L5jEvF40Dis1HuKJIb615G/ACQb4GYOATU/Et8BS7+I0Bsr/7t
eXd17Vltb9nz84QbVEYHZKcLwTj2m3y1jh5lVFZlQZSb+9cEW8wArDc6eORvlWil
24edNSBD7vdSeqko14dnMYWFI+4l42crS9nyavxz1nqHAw4ki3Pfl1m1vnPru1l0
MvU8QEzWS8EVsiGp7skbftJ7UIF9GhhNmNRNei0W6xrLuP+qbfq/6TCuc0lOwIKS
wgXi2aDu4JLW8WxuWrkJ7DMu3X+7CMs+TNwvwNsHp7VH7B43zRnlhLcqIfqrKidG
D4cSajt2EFRrxqbWjQkabmGFYe4I2HXaug0P1ZrXjGp7Nvkl2vmP00nevGnBSE/O
ij/yBGxYXCOu4cODWZS126bNAal/Io6QN7p9fPHbi82xniHDz5utEAquRyk1gywo
PQSAdJ9JioRL4g3gRwDg5Z2yFGHdY9VVt3Xyt6dGwBvtIDVAXoC8gnKUaHK8gw5k
EmA6RL7ZM4jP+WmZquTUueJ3wC17Ve6PkF3JtGRRt0/qh+wfOAh7P2GhD5U4eFUH
jsYNyFTT3Ym72OldhvA2ZhuA6brxLTPXScUkpjvRi4+BZrEMUH/WBM+VTtzp9Y6L
DbkayRuv8lHi/JGfrOUKeAeGL+VU72yZwzhjo2W1OIb5ljJqA607T6DIIvdvyLZd
i0QFcXkNyso93+t921nnPnsFh8+d1llPDy6Piu67HwbIisxWe1W61edYZ5YtLjIH
wSWKY/DuVslw1aGDRSXT7DXDWCy9h7w6q7916wVtK+e9rYpPFFdyPHUSGqSQjgTZ
xT9ccJKcOjQc+r5j6lJVjx9x8zGQ/Jrpx9+iGir0rZ9SycWkGX6iHd62bhT6hO+q
cqYI19GlIi5dY2j1Wgr+z1KJf8Nlu9vkbA0aNzfcmGWhB6byJD4UaqbhWbPknDAw
GwCVcyzDCX1OnmBPURaUfpNKnLZH9K/TMYRrVYnPSWY1zdUtpeUHCPWQQNIxlKFi
w6/afW5HupMyA0akx51hIU1Ut5Rpy7DB8gP+hhbawHdnn2gSrO+TF7xos4VZjzql
x0f898Lvq6xJey0HEq8QfaLxhbyUsKlJduOoAVzke4chS8aP9Z1nHa/hXw1SmFLI
lhIEZmudNieUgMrINb/D2gdGPYigQdxoagEYcg4yIRufHOYjBhDGa1WcCaPYQr4P
61VjckV/rzxcxCy11eWHAFc/DjA488c750t0vuxZLIkTHiLkJypChJUS4NyaOOPV
LTX7yhJVJlTXZAmNXo6hSCYSTFyOecDzU4731MJCxqgGk3OPURo+DM1N7v4pKfZ/
Qzt6WaCZpcyxzh4e3u8JthRdB1UpR5PMp7XtDQ3ipnqq/XyMsvH3Wjy9hZP7Wy3I
9apJ4q+v2cTKMFViiDMbhH6k4oZLybcOKVY2EJj+D4S+uDXutG3dPn1X6ijlCfAW
oqHHr+IImAYQ6li1XJTEykwjPIn34F6wN1zngoQC44ss7YlYNnys8XlUD10cGKl/
Yni875n/QJa8tzhT6cAeyhdWfhccdGePuRhiyWlsQSmq/+S83MUffCwFfJidcNTg
bPrZ2BntijUVnzY5r6yadwcY70teoxjfKXTNDVPLgQhm/ByEDWQYuV2P+LI1iJns
Ss1pzTVGxaJtkts0u1YN3oO9t8p0DeTNSqMNo0/4RtZA78XxMRBoDK5epcuNAUAv
jPkSOTyKfbO/Hmm7/LhiDWOErOoulveRarTLtMFM5rezOp4VC/W3s0EY0PENuDCc
NYpwHzMKKv9NYS0IuP28ooGTk6VNd5W4rJPmgiF0AgzM31T7Azr9iiYZUBgdLD5n
IFCjyv2NxAEFRuDf08Vst4vOuOEI6QlRDpua6//51rzJG4iRpBIyApx9vCc8CCuA
MRb6EKbK569dD6s9YGuzTbYFDAEy1sjqO6Bx5FbbtoFefoDc5SgupLTu3gRVz/om
ckdRieS4dNx0qHDfFSFNt7DcUQt4K7QsIyAoIQjNx6SWWuKSqQkBriT2K29YKRni
/DDpM0t7IAr7ScUquoX5ZmgQ9o0odDBv8PLHkZRWmrkM3wGQ/FlurO5Da525EsCp
tpoxIE7DefgYXSeh0s2VVhkZtr3o9TnmXrJst/FY7ejYb7Mqo94+LGtrcuznbh0z
UwG158p7qgPD6S7pKI2XVkfDRNhmRTdB799wHqewV8nXSGXO/lXaB123VEs2lGM5
dFjihuvWl4nR2ke8y9YdO4bSGltydl6+DETSaCcFgbXSAY/lWebkTqLlVcwo6pLI
4s9exYp/yGYfQ9xKuQ+esDM/XQfXRZdHhyDMT5nBGIBp3zRM1KSfz9HBSG7/598x
G68YAn7APCWYHNYeM1F/ill8udTULcRyINegxR5qvvcjpZjJ6tzSzihbHtsOAFEb
HUmk6kxr7iPyq8AdMbP6HmlwoatihfpT13lnJefOjbLD7Xc9uVe8uVQS/MlwH9A3
DH4s8BZ/bw7mCkFErcEDsqheXhR/JFHm1q73d+hu63wo5zKom6yuRJ2tvkamK1bc
KKLpithurgtYuzLAWtvuWo8g2tEPQqSFmYp7doXRcUXF4mjPpES/6/fGWIqhzLKT
orpNKrgGizlN0ozA0vxfQRi+wz/O7DCqBx1wHkNbdpuav2Gz3LQnK3JvTcVBqbAD
srTT349TBqWkwVmbm19ShrNw99lZDtbz+ipg48yPyxa5QNIx6zEVecyvVxd/EsFP
OmAzUaN1Xo0IyVTVex0UnRnBqLbQTBQ41+uhy82HaSEcTTAUQ7nLG+2Oi0iWSpCf
Q5BthL+i2jUYiiRLVrXGAuhWlt5yNldT/j9wskgRxH11kkxweB7E+wk5UNZWGBND
nF6DDbHV7m48hDR77t8Hc89uN+86/jnqMJw6x/UqNyJqVRaI1NcXgN/4UWLRQtlj
d8acvPpR7B5xRSwNf2qzSbKWbMzOHqnr96/BgyF7WenY4TNY2OJhSiHrwuIWL5Qb
35kMVUFbIWQkXGAGS18aa557rNqnrKJz0bFafw5/4wP0SPTjI3UYWr2ezjFQNb4c
gm0XVsSR7XkfgXZicZcozzKjqLcPeVV1YHZwtAKfMWUuuDWbKhz8w6E0+CY+VjJj
o5ogj5n1igb0lZCpJybPjKNzRfUwd/PnZN0Nal1GvqnP5vdQ9KYxNA/OOeLdPgml
ZGeSpMPRVq4iu2D+8SYVKSzhTWLEow6lsHFLppx/t9OVKAvV/Y1x7sy117rwEI5U
OMIbEb1jXkk5TIHzBfXgCQemKGLAS04PdfDoJBDVbuRWBeyDuaoxBGCBjmpFVFBY
IzSTnlZGwzp4m010oqdyL4NV9qXpqUUkiHhIrnUHp7PjgnQWtPxrYMmtxrhudYuE
I3klPyfhfh9HHSl8qrspDlwx3oAE6OtxnAysjhODkorzH0NvBwl3XG7HhaIjiWcN
V+mUdyzaA3sfB7RAkOnh58Wb4XN+i5O6F74TGCoo/2l022go6C7U6jUtgFGV7ty/
bXocsrUK2brPG+e6hd5qmuz2DOxc2DQYfhJ8dgGxKlVI2iGfWrA9K9pRblRx+i10
VDtxVeGZJVk1nN7DzUjRbukOcjvuJL7mGf8EP5RNB6hEOSwPewCvIOf3IVLRJuug
KGGaPeEKV7e3V0llE+iuZt+y3VEY0HUEdPCn2Pj7/+fQeQnbQPvyqlv2wmQLATUK
4wvfAOO24fIJayE+crBwXAA4JyhViMr9ypXhUVIdtYNZL/+bBZaii9hkOzt+vDOA
nKbkMfcUWKIKNh9qhFHlK1kmxFzbP7T5PlHz7H49+3RKwuy0vGM5En49bPengsUa
xW6xjFmz8F80SKQBOpuJIBK55Z2TbK8H8ZMo2Zo7z+Cy2CYehm/9JAcHLh9Rc91V
Iqlwuiq7Stnjy4l2j5m10QYFNs9G0mSqrOti2DKDlwE9F4KDVI0qzuoKsmKfYhJM
cGUqMheNchxMDQi5s0XULGt14PIYeBPB/l6NyDWpZG/ovkJB+mjVerzxOmNv+NAu
atxcHcKRjU6q9T8slbO1ZeUCYSxE6RayOi6lJtXRdgjeh4qX1z46gzDOQ3KkGgbm
QyW44rEGDSbMt3tJEqddSXK9xfjDAMNCkAW4uaF3CM7x9I2fayt9RENHfiaeO3ny
ts61Vkcj1NImriFGf1IctTrNqKYOFsQKHgbtmf4X66Q9Z4THaiKz4xuFDqi1AzkW
LjmG7NSbXHcGp4dehiO6w1/GcSVMUGuNqj7w67t692A2QI0OOi7m8vxOZwZXVs/2
5HW528VAGaRaO0Lf8e37SBgCHfDvIfk+in32CKU9zqb0MiX02iHGVqdTPq8Y5ISC
prtwDyWY3yzBpsjN1r2yLUChOnoYD4J8+zj9GCzuCI9CvKFkPr7lZ1AfeVTIudip
PQNnYkdi8hipvrgFcnu6kG/CIVbD2AeVc7fiWxMWQCeL2JaGVQvLLMPZvLxvcY3T
qzqy/yqO0gQj/qrql0R3sXm5A3l18F7hofDzu7IBIOCva2+rDHo2zIXGP/UsqqtK
95x7iW2XXNkQx3ZlTOK7Qz17zW7RGNTJ2n3CSp1Lu5X2M7U/urRVwfAiOt+BWY6P
IcN7ztiiC/6btaBvWJOTRTsKg5OIFakr/evI/uC4nbB3KuGv4ZogRhp7XTfS6hIl
3a9YSGvo2g3xQxJSbOEEjyK+1Dp+RFn3GWJSQpTNCY0vQziQai4uu3984JKTLCkh
y2FDtRfmRMV8fUlaeCkEelTChdOEgZ1LA4c5FQdNWBARG6SgVDLudbMYuTuayidr
Sl+NCq6K+NR70+mwRyq+vyAmXwUQArEEQCCIxKcQY2Au3NbadbSZhgoERqQtfedg
iarNYwo3CJBc/kv7AWk3RoPsKTdpTMNwmfowOCZmDerd6LJzlq6vKHKtwt2WTTP8
mzK5/Vz3efA533J/eC7ixebLYasj3rahInh4IrcwRDE36R6dPpgMk6+ovs7kXC5z
C9nxVr5BMD39oXrxF3517GYOVqb8jphE/FjbikJXNFZyHunkwY/q7FA2VXyyFNFE
roma815zrmVUpWyv1SjnO55coUomNcrP++Hr0azozNT6ceq8Qxr1BioRYS2t91JX
PC13KK79O76qXzk7xgunfqi++fmwZPVKjPZqBXvQlB6wx1WTAggfzSueWBHZPHQT
wMTDA1xgvYB3bfoEwB2+o+BcN+alO0RHsmRI4GSY3dCHMz/l36J4qigLkXU5xxte
zhVUw004uyBr+7YNxu3KsH2WjCthvwBfoAsH7VMccLdwzJfev53jNHCKCJH1OT8R
5YR3KTj62+5re5kxdSaiUPDAHxDxm9LTFjFJWbOnr15z1djXInm6uJBc5dCbLFgZ
tT2Skg/fPlJTyu2vJM1xlpktUwJ2ZNApEIvtmOXwZFVw5a7SSh75mxG17iH0RwAh
fcw0ag8dtHOp4m6fApcWGxpG1go8qJ67WJIhfPXDkGeO5oiSxIBXhFhFeFQLCDM1
p0ZQhsNN3snVtdYk7LJLWpIoAXTxaudo3l88X/HGXt9ehQvefQONnn1O7X3WvNhL
YH9Q3/6NX8MxcqKBFxSMm+018R7OGn94Wy8kFy3H1lZKtrSRJmWO+3lsQzTqIKGZ
HkE01ylHVJkp4Sbi1QTE0njmY2/NDYXx5Cw+XyGmtvEzLylxgVlRaqXvUYPR4uqP
8bEh+XC5Dc2THTrH3d2K3dVYOLYs14GpKjKoVBSy0I9n2IqnOqqzXUQ+wUwP3Fce
wVHP0mEQ405fUq3T4yxbY8/9WAl1YuXMrm501ITAO9/Bon2S6P5zsPdwS4zwtO18
Wry4Oyy2XVddPl73pKZZ32OA4ePAVXf2rd2YIz9NkQYxPKUSESJF/oQp53epx+OT
xo69U+FxBsujE+nqZ+kNdMM5Zy7UWG+//rL4bUvw7mPgXmN+7yF2dWu8Mce1GPa4
DF0jDP2keTD9o1f198exrpwnufqDZFgNMe5inc1K2oFGos9Tu5dszVgZPbWfEo99
RxITBZuP5/15z4c+ovZpqjsE4rAVZFR/9jjeP4kLgyX/XSebwvoWogxiLWoElAQ5
RF2lxu0ukUDPKS37PqO5y0b3/sVhSJWknCT7pS0Jx6IFkGtQm3trlhYRtEQcdDUN
iPnjPtXwHmCnIMmWGKB6NCtrG5bncqLblGG/k9qjKd2NtQ9kGw0SKtU/WlY0zLaF
La8WMNHAzUG9lWPFqLimzonL0MmQEdaLUqZTYMQPi96+6GVfbLgQOlQRDNoOksrg
DTTah0MRM+DN1UnSilpEaLndNI+Cn6QplnQ5es73PcNt6vRfhKVZb7B+YjIBxls5
KVetK7HROo2LBNxlAafZ+10z7yAOkTGGuRPsr2cXfhcXgUJLaOtouKiR/znQcWE0
3buYtkTf/Xjp371lT9H65AxXuDaqY+wcMzLzyoaScY4bmmWu8i/bRfrmXttP8C8A
ObHyG16ve4xX7/KrPfWN9fpZs+i/bcDEZyUd5o0PBImJufvWjVjJIWlWoLTYx8yu
Zde1Q+BCUfsPEzgakVJTjg0HqoGGgpEpDrtcScE4QkuseVEoTf1aEMK4yH7k++5O
qPZ5FjLienUlAMVxOV8pEUHFHDCWikzA9pC+WSyg7DtWNF0kzypOz4zA9aBtSo4s
b93x87z6hXVqr1lf/rtbnkqbWfXCtU9VgSJsAIwiBKUE+zmHGZV1pmXy1OdjUBnO
8SotgabKy5w/sK/68zcGDYGmVDnupqWT4bk9E8mPctns1JNB8i3BrdZY4e6eetoU
iWxsUKzWRDEH+W+84YzicbmDQztDjVnb6l+OTXPEV021bSw8ZtXub2DqW9xicIrp
tUJqjm+eYLeC1HT2VoazcIAOVdaY8JtSoIH+qZDl1DkrpdOSEreUlQlJfASqHBCy
K/IVhewQ0zLEMZxBYK8IF+QqqBzbqFAZAEN+UkBbNvbRFatQGszwsBlURur/ine7
K+ef2eBeUdiqt4wVfDushaoIz5qZHkyShce8uMKbKPDOvVwasJutVR3muWv3eQY/
rmVmUMUxrOwZaLoMirp/6VU7rwaKUUvqC/UEoLYAceQfPKntMQHshRtvHcSij2d1
pzQYnqE7qs5Y4HXmIBdSQeC0yls13L1/BhvaQk3MThMcvzRezA6/z/qV+FuwhmEf
6zmu0GmX01udhxcoF7H1TAWQHDrsuxfqlITSTg6xVUlyDjnlvyqxOJ8h7q1kcVZz
/rwDsUjre9jhJSYAStt9qH9VsDcVpUnDFd8xiK42yUr4F+B4d/gU9EkZNJQyFmta
fpanIhJ8vKSahu4RH6KhXuu55IXPbLhTkrmW2yXTz8jbcALNz0cnggkUV5ZQD3nm
knO9r7ikbakQartrAw4J/VtpKBnBOypFa9tigWAGeIGiIFcG39WI480y/hLJ9Qcp
QUlFnsQ+kf2MGwgZutEAbMsDqCem3RJZ5amsFNCZsVv8D+M/xlAQj3Nsj5X6JYqY
YBfFhqX7rCRkB+CidowZCuT9LVJWn8aXPzrlYX9FWWzPwGaDYZaiTEsTJgx8VG6x
Ax3fiof4kLAitEi/zPS5prqRNxsiTfBkouXEs55SjZB7NllGgFJ9MyPz9ZqenQEt
pOr/0Z9niZtAFqwgQARKCwDxL83otMEY7aJTySPviAa/0X6rkIJFttyw/GsL1gH7
odoOhE2MEW9M65ALbZeXIRPnaM2pT4y2fnn/JCYG0obGKvVY4wHDKNySsCq2s8ld
d4ZwPVsmkaPYzikvckij96NLfERYfTPpn8ry6raITks63H9U7cjvF19nV+6lNEei
Myo5GFXKuAR3+f//FCnIadMCeoyuHmhSxguxZrvuTp+wB0VG5Vj3U2cVmIKroOST
dtrLY7OC/6HpKhuRUTe2448yjPtlRssZKMedBuBSSjdMzsegyk01jtZx1pFA+5Dy
w6VncvIOxW+w6pq5B11rqF/ikd+wpDdiNKXyX7SixWGYD71kamLAbiYNAiRSiZ3r
GB154vuH5loOIw1Osy5Vyk/o/LMpDAx0sX0qpWvbm+d+eJ7HevIDi82BbX2jCjeP
ZHo/xRYuAmfI1EfBZL6vddRCTilxd8j8tqoqHqZK7BxWxEgln7RfpaG/A/SV5lcJ
VWI4rmDk7E4naOCIrdCvSM/azcPQ8+tnPsqU9xeP5cPIQOWMFnShYX4glgW1v0pr
zX0CtKlzai5EXmh9lp70dY0yaTie9Tx+kmAz9dKfQsiSbZLy5TZHQyT6z6aDDPmQ
FO2Fvl/t9v30zsKj5qkLOzis2MN+/1vrbeJylJpkv2wwoNXAvNK58kpQ7hiaZq8J
k4gTSN2mCZIz7xDVyd7QJ6pFKJZU29j4HUmLkU0PY64pP3NcTOaT/CbNIjs6R2AG
pq85qNZPPhRZEaH8fcLHmkPv4gdjYmYrx3v1I8gBkKi9CYh91CKDAsDLlL0JFjc7
KmcpNK4k0qKnuHvCkfKHUeLsDOmZwJ7f0F3BERq0MOLRfQ64BnW0NvwrI+ngVPkX
Oq3S4ICl79X56IFe97b8bo9MXnmI3o9/YgCpahoG/X+e6Wb3z3zxUtsYrP2HYx3a
2WF4sfco6sqWt3Zds3CzXltek6UGOU106lBTNoq731R08soPh8ia/ArJAgU9THjp
eNZMacO0Zw64Nf+AwVS95VIsmMG8JME1wlRxSarJi4/iTalNaImjORDJ5dU74Oxv
7INO364LxSc4m/2MO/5/CATyR0sQQMabYR8DC9Ue6wZvT5w5EEW9Qch+oHUzMl4Q
r/dxIbJnIFzsGGRcIZfbOvWrAEzAsDDiAB8VhF3kj5pbhp8KIx2IGJmthuIjhBXs
GD4v0hBJY/MakbeozDqZqD+S8VmmttCXDEHrbyWPGb27Az/g/PPM5AG34uHKn/+O
ZnRy3tq8tN03ccfkZDUpev1crtZVbFVju72u0/kQZ6g+QHFHySSWqlLLnjTkgBHk
UfET2IkKfiYUy/e2+pKPy2HFFg+F60Slp2D5C43jNZKkYXbrqluNRxaM63t2skOs
5gEIJbgXVUmr3v6NzpXvDkIarkohVedLVmc2fP3Ef0ZKmkDWTTUxAI34Uk847YCh
CaSOA95kGDtmKN80uhyhiU2sABA32Lzq6qKkxYnZz0zDui94edy9pXiO2RZwIO/3
MUuaz8jCl17LQ2BSbE5Y3i/a2omjN+VmvgGghiKlnkPyqztDnRPNI7icvT8zofHC
ZahjtDzkhu907MluUvU9vbdcDZyqSWeJa4WUOJ6eguJf00uNbW1LX+wrvJJQ1JOL
QxtzhI19bn3SUaTDjo2X05aA2Q9Cajh/D9xKr+itj0ZXQx77ruUjlljmwU+Pm0gs
fhO4wyM0AiVkPT3zlrtZJ/kogA8ST6xg2gKGzrtbaRUZDzAd/LsRYSgQJ6mzdsN/
ByUlOiuHlRkYqkIdNtkTlPTq++VlJEUv1sS+kPzMEPQwFWZkfKYO3FhQBzj9RDK7
S/72lfZ2pMMvam/ypjS5mqIB0g47tOah7TEvO46qeQWSTALQ+8TxGGt49fHX6Ife
FoHazpsUD0YZdPBK472LY7Ve2sNKB7VparGlTzth0QY2VmcIyIJLk7SymIVQHysV
027oP8qDMMyMfEoYxZzKE0vaXlZzhxt7MUQ4ruGBIVb6mFa1aZBTN7zIKfED+gXQ
f4q1zrzB607Sv8Aslc9Lqo5atpZ5MDBYz89GlMuveH9akvRpqTQaj3g1q5o5BenE
x+/7J+sxQaP+/MNChO9BE6AYaRyIbkiF8cGH2Wgm3uH3Q+iV96sj6Jf2TkD02xUR
K3meXvR0xC3motlwelSSMxUNVXx1OtogrKTzSgnW/Angx7w4HUNoknFXSsMcdLXU
6r3oA6hlGE2LTD2hUydDt1dG+TAXm3wyyK7wnnlN5TBTPbXWZ8PTkTBOZWlJIMcO
DV0w67DahownyLDzSercJxMLs9s1PoFLSODJFZg7LSt8zEOLpjTOX7mMZfZ469tC
5meVpxfHCOxJcASbuIn3pCk6K8WBO08MFmB0yUTFvFZsQ/YI2OzC7uff2saClCGz
mFEarOm5jXXENBYwT7B0WFAFksVppiu5udt9M9BATJ9QgiZkeiQR8ZhaiPDIdkgP
jxv8XmYPY+dZsoj3AGjeTERfido4IvavV4IeIbOoML10/LI9pU6x4HPPZZjIfG79
NpPVecP5dIy5xh6f4u5MFu13fdv4kq0E+sLYUUnD2mBtIv6UU3fe+cYoyPH1lDgF
Y1XM+2wne7v0yNH4ABbN7SzEoACo7TfeP3lzpKaDO+sLjUMRqvFPH2q85g0m4KyM
m4i8Hll4Rb1n7ITEnMQKUEI+nrAtY3S429SQSPBoLZsvXZr59m6UPelpn7pEiMhb
d6Tr5Y9+B+6uHjJkpTAndnbyqbJ5599M0IevB+mdwv0Qmc7pJH7bnr7P4NhpkwiH
peiPUPnn8yLnfgnclRYaLfXGdFpoqhf2VWFiPlw+LXk8kc1T9MvRJlrwQwAZodJW
QillPPocNUAdZQgVzYbTjPqsnGf1Q0y+22eBMPecaf/e35tvKD/SfEq2iCHuaRs7
HfrJ6tg2z6iLMtJj9dUS7YycPp04qed/Id36SAib5XTqCVOD3KMmDKZ8Ryo8v1FV
q6gcbJLeQy4Vs0/ZBKLxcP5YKeu2rKBOCXqxhkeSERTmml2HKBC9NZQ1clM2k75R
JzAEiPbPjnaXR+/UKcgomR7VbY/gp72FH8hzsDTsNAJTUjQ9kZMSwIsIh2CGCmsB
6RXiBHr428nb8RW17G5NU2immVhVq64b1ZfEPu2W1kmlOJPAQxWEkLMqnrX1freB
7AljnfMQsEVznE/rBiamC4hsCWGFSlN49Hcl5oh6dFWLXpocXsE/oiuwJakjN6Mf
pRkMDY6ioVFajyJgRpWtDXhNAKuIhvBCjgtpBBeWmk6JVsyY40mkX2e2Olq4254r
+sr0g64Ouq8VJk6R8ufFuJAiBv03BNfqs+hEE7+x6utbSUujmGu7MgPB0Qr97TTS
Stj76j3+In9sejXMzKl0qNP8pttqv6PLHoUdvnlZfEfJMB7hxbMjFM/mJS2b5jet
g/i+olDkcAcLNybxeWIAcHBRTakYVQfsKDhpFl8tGw8vfo14+gHsBIdF/uxRrTX5
dbT9G3NIj8BNt6zkM0NTQMDGw1Z8KZljvlPLw7mikqWwI5aeBz/eWsljG1Hdxg5w
mIXEFlrdHZlqPO4t+ohv0d5HFVDSbSR9fcD3mHp0dohcB3UT5a6ywAj3WoiOtsZG
Q+o49FfKneGCZlx7LYpNXlKZdvUT1lhDHg2F27vQvVN38sY9zPvl1dAD0JukBIWZ
7RTeWQrWrnX7PUSZJIY2HSM3PNS0AjSuid6KuhO70YAVYaT+w+eYAQ9UmWsUfT+P
XD0LYn1AL+gZtRXoADL2hQhMQkLsoULZac0e5GM5lwo8+F39h8BihwGVcPKmjkcU
aqH7coy3SAL1q8GsIRjd+4VAOEZIh7EgnPr19NegwRhsfKyn7p8K92gchsktG1dm
OTsUnN2CR7ZYM+VNIbRogFSHpPYf1jZVZvJ5Ka8NLHT0MHfN1H1Ay/o2XaK2EuNu
DcMHLvAqogeTAFZQXrfsRXNe/CKR8bUKWoNI5df364lOaefdPOPpyzuKj6E1GA+q
vqFbiXvrHEmFlzVDmoAip0Id85BE0qG76pTmIHHFwjcB5HMtDRsBDTK4LUBgPIly
N1o4S2G45ibl2Qu5eO0h2dSAX5fapUTJ0PQ6BvXcLadG16nKXgNxasfIhGkjWI8/
/rRbdbxZNUy9w3XJ1QMzUMc3CFfeACN6IhcIIvr90nX6aC0nVpxiaFB5B93qdA+M
lJDeP0nqWPVJwIfhBedZwIM/oyv3mRWGkFxbbQQpLZ5QvD1rl6TMSjkPKJH2A+k9
To9P81OFqrX2eX14JUGiC+fp9R6pMrEuUrsFStJzeD5B6ucf73RFhy32jxz6AgC8
rfWNlYkd3D3gvac3JclxQNy5+afbKfZqcrGfLlAmo+dYcjBNmIuNw2TBTKAge8tu
FTlI0UC0ij20mYJesHEwVMS3PcA/nwl1nz8l6K8syudOE8kVs+XSmoZ1r0hWbn/a
xEn9an4vrgDWO73676SXbnu+3oNyCCT0i0TppxOSHkKuK9uRl9noMtWqsCI0kiZl
mmyB5gNlg8VJogcBxqANVoOJxMEvOUfuSHPNXsSORDWHk3zG8xbCOBIfXmNk1gxb
+c4Rx35LR3gajLk0jkYBNTxTwudfqrWrXAqvbjybrzGAqk59QRGgCZLac5bT2yJV
ICQAJPwd/IAhargsHSM0y2wCRBJIH9ZkYlA9ZP9vr9Z7+s3FS1kYGhR/SenslG0p
+0W7Wb6EnL7yyCsMFaAxQLU5s2UgzyTGPvRf4PWTAdwxkKqHPNgJrZ2bfJx6pZMT
fy8H8PeAfDQe30TE86+7JlCcoUybpoKeBzphxxn8lymaOEtF+iWfD5Z8Moc4VwAK
x3Ek6fEEeG5H1mB/C9hahcchFwOqbFrmjN68nrO535aagcAkBfb0KyfSi1DZ4DuC
bCaSsEPHx0qUSMIVxEqPXqaYYL2Fxdj0hevgfPrtKu9erReULHh2+ZKHJ4zGEhVM
VU9sHbksfbWzwnMjtJKu2KTsBU/sfP2TfZXXpbzXlv+p3jvCy3Kfj6oX5C/rdqed
uLaCdjnFNxbHbUSS1cDpypNKhdS+C9WVaOE8Lcc4amN3uIZ1c6HY4mpSmh0BPmZe
HoXW1ieMSd/5oj9rmeF47ntPR/WWC/RGoFl4BUct90IqE2qgfPyxPE+QPqwyJmVj
hV4+kacwX7PRw0FFEz6DGU1qrjihYWMyKdSZyLb9r2wB6YlB+kMSOKsUe63nOmZT
bfu8lMZiwgH2sjedTtKF+Mt+7AvEKcoxJ66Ri4d9zs78CkIGoe5h6gjhvCJZ8cR1
IaoqCrSEgpHdmV9P6o+Vg3OXllKioXnZAqfiJMVEsALfFvrQuRAyexhm2R4QY/It
zH32td6kB94/SJQ8ENGYbZ592G5d5U0SWG0xA0A4xzRk4cXaA0bG5tQK1Jz+0FLb
hDLdY5/ljduhdNCDCOfjT0udCXVRCSvc3n51vbFWGD4MGh+LQOnLrdOFX1Cokt2m
/6Lok7l1jMpMrN44fJqfcrC9iAT3oON4ZQQMzo0FDDfX2and0z3/KCTIh6CsVg4z
DCG+KPM2Uly+CUMMWz6ZuZY+wGJr/3EqgTQkhGWfv91UYvj9aifJ72q+WDBITqBw
5lwkgrOlGIK9P3EceGKrovoYdgNuPtyVp+5SIw4RoZWeDPZd4aFQtCZTrN2Y3/Hl
BEpb9ZJ7UH2wiRswl25YZ6Fg1YEvke8ZEimlqDAN6895OuZOKOG1tC9FOVoQVlnk
JAKcv6BmDxmEyyNNraMzXL5WgWzfpfQud/ik7Tt/HlXA+rL99Vm8LCZ0iynEDqry
vAdSC3zGm/4znY7NlxDUiEcPzs4qKiVuxHKzb4qfi6HdPx+rtGRTn+jHICzylMHw
25W5mLEDD7yvq1Uhczw9Nek5Lm7YJn08OyuOkUrE56I8M3GOpIeXJTPxAcsZVO9P
PgajdFJ/yUE+FoG+63KhIJdCKyoSRoHSYRG5YbKAdOW8+gXwsIN1wnkyZwydBWB1
ubczcrnBao8FY+IyPA1PI37QCLAKYIFDVEfX/5yEgyWwE+LoviWawJ7Jz2ZhtM39
C/vDWSQXyZzxEAX8KhxT9oor+iOpePib9HS4enY+zFev1FgbuE13TAdWS6n+zrXN
VTu27aHoZ/u4n+AC67m2U833kgrMMiHGCACzeMgengibT8oZchQVI8h8Ptu3IwTb
eGOYIgeH2b5RJi7Ccm9YFkks0gkXwS++FGnYnUVmQvzHPM6Rth178z823/7IUSUF
eqyPwU7Ald96ckGsW4tm4E4H4eE/xpARO/3y1bjb3QpNevCh/hzstRT7hGtFulVl
XuAuHCc81Bcjv443TTzfcyW8XFX+1fB4oKa8coQXkdnmDFIaDATXZpmhlXhz338C
gEGRArTtUQgn8tZaR/7oDdebkS23WZCsGxI+JQOAGHPn6ZgfyxvxPwBjU64y61fD
zgbSPusVWVwBG6TOeUsqQs24cBYz/Iutj7vcVRYSSW8CPyapZSouWpikngcy6O14
9evPg6ToPii8uaYHUskKEGbBRlYkVCBMVCEdW2oGaV1yUrNGgngSbtgHgI0BqYaB
8M65AseQHQWnsOyfTyocRJ3aeGIEjFzLyBL6TrPhSJW8JRxWddzqaFOLBWKonBMl
noOXtNCFSBQPXJA4NUjWzFSmCWpYPCUSagSjglTzNq4/zhnW9nV3FD9FWmqUOMnD
d0BnjPuQ1vvUPhe8bzC92m3hjwl37T0/z63mPOzRR3T7ogj+UhVcv+Cghg2K/JgA
KAaoM0RoY8q5xK75CtYyMiJDQST8I8+RfNliqcUq01e+CjtU4XlmWVL/yPEdJVg0
pjpPP51MFhioYELmF2fc+IzNuEsigccKDQOJSEPc6HG//51K/qbOIamwWYrWBms+
XiEMkkxRZ9MltXJupWDdQvBgqbBLCpH1wvayJQNUfUqQnaNu75d4Yq5OSvPPUMfR
`protect END_PROTECTED
