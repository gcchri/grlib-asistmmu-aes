`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EKfg0QM8mzL5eR0fPO0GNzdzOEZOPJ5IQBO73x79gT8ElLH4n6HDMCy5n11oo1L8
OOPh0bEgAJSpJ5pkIQdz7e77a7xivjeCCitVSZ+AkWItEUdAs4Xa9KKEuZEfP8Gz
JvDjy3u44i/J8ko9ATfHVebw6C1idOv/s86Wg8VDYB3cVkf9afxW6NXD1r6HNqn+
jqOOZEty4kzpAK7b7s30dHH1D0Ylwq//jzmzb6owOaxSu558dpKg+9S9/26Jz7wi
1maP3essOem/+wM9/kjrw7jugons7gFZKwAU/E69yB7+Wi6Xrtxml+PF7AIEcqGC
eS9N+tF5NyNMo4R1J8zZk57z80Y8sDPtCZ+AkZ26e/WRRWhsuO9yzvLnx0+5ZGLg
B19Sdo3n9Q+DkYIFk2e3ugCYzmYVDAHSAFRvmyfazLqG8lxQ/c1Ng/lmQg+/g/Se
g7QT5O475YVEziCRpsQU3YPk6hc5hD9j3wX74RIdHR/IXoEB6YbI0g+fb1SvA/i5
3CI+HgExsOl5CUSg+dGDcv5KDpipA696dg+/qZqgYxy1m2vxrPv2sA8PKPFfzxqg
ccFphhrwnQ+PQvCz52KVh3VlZXlc4KgmaImLJjd5sFSxvpOx2jTa4MOj5dawkSab
uGqyBIjSqaVZf1y5iNTkvp+UxMVcDewM2an9PblvI8oKXf2MhFDwkBSVR/8sEQRp
k5/jt7svZwvw1EaNF5WqWVeNto9faTaPGGPNep4QR2L78KPg4FOef1/GCRr+Z/kz
LuTO2IlU+pS8DWdj8PNeBVXBxzZOg1BArJcAanLOmmckSAtoXs4aq8BlG2tchzal
/AJWkZCGKQeaskDa0HqeMz9uBqg5fRL+WKSUa1t7ywzOMS7m+4yVgiLL0Bxle1/a
AwwftVHnpwjLFXtChlUJvVofTzkaImP9Uwl/0JezRfwkJXwrP6fLIIQd5y6wr6I6
7RR/9/k9yn60aR35nR0EAnOUVUNj052X7RCd/R3pCnZYvGjb5yfeq/xHvQ0tFOi1
CVcs8+hSd6Gvi7Q0sUqz4dZWFbD41ynbCSmTbJu5J49irVQ6sLIi5AaU54k458J2
7YMzDHIRzBIdTWI9EaGufGXbCc+7os/P5EsZKWCJpSuiXT0jw9zPCctbBnTt730W
HlQLlqBIVURTNTUMWiPv6P/98KGvv+MCDY37y1liJ9CJY4fwTj6Q+AM5NBJCA65q
tWGcZNDiRBugipOsXknnyGej5V4ZHH48tGTXTYAlkBRrpVxoYKDIFGXDPBK8659M
gftmrH4Um/UjPeggoXENaV3TMdTLIS+s0XmkR0swUtDBFxWDZIc6YCotgx/NoOof
j8Szdbf2YNy4oFaZ21VYE/002j1a6wliIP++uPgFySAn2W+KXUxK1lxRpbZvlmmJ
/syXunrCZjaZVAfoW3uetaT9HP3rZsEQQtjdpO1BypOnkvGNT0Mg6TLoGjGoezwS
LM/xUe6G3CbUeKq3DgOwkZBS6Hw87JdfFOGozOPs72l2rQCEdL9S2uAVeP7PxGmQ
wu1PblP1aCqk4dIOy37s1KTJYWPgjOUl3J7Y50ccngXml2RFAPAITWd8fqrEToOg
+W85bIH80wOA+b3hrOAfeV6CfjVlHPRQIgDPezAz9W+ewX6d9bG2C7iL2wbAhcpa
o1El/hisuuXEvhF6rC55ArDkvDZSBLQADd0MOgGwWvgmCzWn15GZKTVG9c1wsLy/
fbTqH+Z5gTai8Exu1GOJaKk0z+mZShikShIoFh9Fa46VkOXV12b9DsBhOT/VpyD/
EClAdI3wHaeISETpeSuUs9YOP8KjCPomoHam+Ig2qJyVV64zNKVAdJINtB9Iyqyk
ATxYZ2OR89VkwBkG//3E/mWsC72TfeyWrK3FgdRO4F2K5tmD2KUJJzOIpBADf8Nv
O5laK2c1+Ayz8gpk0KXpyzrJqYY/XjqpVYi3/zPzE7Nf5f3sq3znLBHpom+ickmh
AntaF9LS8T1XOshsdWTmutfzMqTJ/xYUOhSWqGmbLtjUUEgk5jdrOGWhY+V5cMbR
bHApihvPFk+/vHtCIIbhpyn9QuuTweVJe61ye9+L5on7Gf7OUz0UrKi9EMpvMVCh
I5OOLW2u+DthBt6bGhDaB68cAXNhtEjQvZk+QOpdTH+nZWPHO7fpuNZKPJhZLXt1
OQbVuYIm9k2TGurVQfmbFC15qhV4mK0ScuJEtm+FbOCkAvZg1Sr3T9H+McC22lqY
Smw3rC/zWAH2NMX/ECxQGRKV2O8TjR2/fMlsvmoUNsoN/4JL0IQPpQK2my0+v5hV
Sk9W+eFhP6PSmnwMm5AIncA6QiQ6UDcC9d+fEkwRRF8auGnq5t8x4ib4cpZpLqrr
iZdmSjryei/RQRkezarEBsolm/KDiRC96APEewO1ZghIShtGKyjOgHJgVXGGAPcg
B2Shpj9pg+X99QewdJ39x1xxgOX7vYh0TckFCIqc7HVTXXOFStTRJ/cdxTX91ztb
D4DLNyxR1vzhvaaJXwwz2J1NOs/SPpeefSrHAfFJIugwbPvnKSFYd5J0cW0BN2jY
I643pk+q7qCg3ofnCjOSm/YsP2qHc5E0GtRN3EJ+Y0PfJXEwCVORIXBMVaI/fUek
DSJH5PNn+VPcYSea/3RjajtfIU98jgXMyW2Ogeti6FzNNVSgwmIUuux/yiGj4NVR
Bv3PjvUYBv6+raIpHIOfxTmQIsfbSepiIXkT4yHJKU3y07LYHHFpns1TlXm+TJwZ
DU4/MOClNlUOEJLE6udMHADzoY1BZiZrsVN+1LeBzg3prQKApcU5GHkDlVwQe2i1
rPjea6crnZUkXdZ+fImk9n2flHoa3xHEj24tpjx9xptpNbJHP1VyRZyM7Z2C7DJO
uJ/7DGDvBANhiGjiUIMCLWq1fhSpjQLdegzt1V9XqnCKQ2qvUBfectVBChRrobOf
0d35z8WqEMYV8k1qe06WFDQ7waKTiW2ZTs9f1B4QuCw2X84mFZL8a+M5imNez8Da
coKbRhCjrkwkAd7DEQjtAspsbuC3yEaQcYiT99zaaXwBuYRclEhaNcDtJIwjKEI5
6aX8vLNhR+dtQ2KdF/exyAtIr58EWnW5NXeyfowFRwmXXf16nf0KFFXetGhbm0Bz
C4avkJknf9m7+POu+MLaTz1XYtJglAp+i0v5IiIDg972l+7nJrhVla+Mhbu9HCxr
BhhtrymeTdHM4PtzDvU/389l4tokK0tUoeYUCfTGLg//Qqpa1y3yf0fB8D7uekCE
Mbta1kX68zziPKckStOt25FsiplE5nOpIpaKP0JTGsmDjUFZAQnPm5yy1KwZHU6/
CXZoe2aOvueb1AkYMfuMp4NO/f01YK2uU0yENwK+yZOx6CL5qPYGXyIhPMVSBFIN
ugA+wshjhLjRK5cNDfVP7h5Ql/uvieHN8zmkANh3LUdJZLCboMRw4yUWRTAnb907
AegEu+5NcYb8V1Lu7hHlhqWLPZwi8IGXtj0ZTF3K3oduEkW8KgYTHCEl3amwOH39
WkNmcVIU9321lADgXdoPUwvKpDhG3cP3C40MpKJeih7iOg6Ka57AdLQXzzGN5swW
xXjcykROEyI5/OtpNOgwkrdMtk7+8v2srlaDvJwE4XUuRPs6tGgZGjd8i4dD/RhO
86Lf3/J/p361+bL3dplH8rn0yyBfNbkjQmCIXnBVCtkfFNgUFX1OrByN2qsZxJ9z
EE9msSOzvgKEN/gsscgG3MODEzL1KCDptHNn83SRjyQHk23tLs/De0w2DCAppCGG
0B/M9YYKBTrFTmmjkRPJ0TS1DdKmrQdPPRkHsJ5psB3DNMqfa9Y0JzQREnUsrFTu
MLFOe54Q2uF9CqXAqsaTmuOAgbHufg1GB9Xc+YqSLyO+IetyAiUx0B/KcaZGnCmf
IfKPkRRLmdjBCFFS5xlj4EzPRh4E4AKCZr/UYfOp5praF/iPD6Jka4kCFaiUw3ug
8dL9TCAxVfWmI6L1CfRnWjc0aknWX+Ak5pfqshouZUDPaaOMUAOyb1KuQwaQiEUT
2gCmXfprHdVcmIRKzs8oteieWLVZaRky1IRSS65NqTjMgsv9oYuhxKMSA5JJiU5U
UYU/AJ98Fi5urtqbz2JQ7g2wAJe41MNV8rqmjYCXEq6MS8vyLYCAlyYwg9/sd8Mz
aOKXZFUrvasOe3lMlUgMFKaMpOpfSxMcr5VME+e3sXLRwUYNW4+j8aQ8G4DVhERy
KXlfybBEsBvLDL68nvalSYN72oqgd4hpJBNBvF6y0sZfdbzKYjWeTTOEFdgj2f8h
CvzSt7rc0gvM/8bRCU2lvCpisDDsel8H5sz7zB9J8dk8k7qyA3D9tH96MqyoewFL
gQ1E4aNstsh0lAUXwc5kfBXDbZguq2NlVIWLLNlu2NwiAAC5vA7qmnHoEBIChmWG
u2YpWwFoYbW5IaiSO9HeQ3uGP7LSdyLzxvPMvBH405CktDAmtvD7KSaY+KpOwqiF
cfHSMLViyUdUOeyfUp5ZSNDbeUdPV3muJx3esBH5Mu+UKCs6HsysPlRJ/7OxV6fO
3mfIUDdOFA6vR2/0NyKI6LfBQ8bclPaXVzFVVgPT3U6/DjYTHzZuArLFItqps593
2og+5lfoVOoKhDXguMI56e+lI4ZQ0HPb4RppZ4UCGlAWMRsmoaGi20T1ykeOaTvx
gQHciROSmV59ZDXI8aVDvYFRyazKp/KCFuqb5G53DfhH3LVXyPzoUaK5e8ZLYgO1
5mWa2uWCteB4wxTOd0MndWW6aVaiQioweiAAi+DtCymA6fgP2tAl0eO3sc8CLDrm
QVeOg/3eg+g6JVTW0S5FK0d66TatHpJpIz+NOuL0gtigXKxFeW3P2VOPOP52PUI5
fShjbEx7Z3DIYvUcX4VxIWmuy5ZfyD3MROVPtc/6Ogz+yXrrWwmCTIciSKG8rLad
EVSMOGlFYNyABTurNiKjjSgie6tDSd6DtfgVhnwy4cBh1wjS+K/Fn5zz9sTmMCRc
GwPPSLXmDlyur5hHP1CriG1K2Bs4JsZqeIUb6WgSh4mbRxcJmhtI/DgZd+clg1II
z0yIkQZ3RcMFEPjGSNUnm2K1FYPAqXlaPsl5z3KMt+YW325gL/jJ/+jJk4PbpGF1
FBWq3LP94PdiXMhg1x2o45szfvIWOPLQecOtS06LzLXdrp16iEpChY1LxHVPuCLe
LQQon13pD9Vs0JV7GmKBIG6rjYuWevi/nO2zuudKA065UpAXPnvMzA//GZTBr5qi
MDoVArFhYXEQzAhxMdFSmRAazsSu4rtpKVWvMSuGdhbmJlMN4KEYI9zpOQD4BXi5
QfQuPYWLCn7OXovDN6mj6+zTMv+Mqa7eKrPM7FEQCcoJbk4pyAkiHbG6x1GiIJuS
Ww50djFfSKIEmMgOMWnGmVUxUo3eC2mnA0KeXO9X+nnPy0q2nzQIafEstoixjNBm
Jldzb01MhwdqoHTnCPQZiIE6ePS/GQGnsW4W5RutyTbB81yZIe5U/UBSwLfUVItb
rBfqZ9fHaCpsVIv3yMSz1NvUJm9C6xVM/RID3GpubDTvlhirayHWDQ3YK9z0+/uz
EzyouPk5znOCH0BZbeLTyl7ufclXcnMW+1O0f8c6dID9vIGPyT65KpG2k64jBvb5
kwZfoC0Y5SFvjaLFLuXrJll0LqB8QYpHtjHsWDOJ/N/dfpWqtqgkZuCZWQ7i5M8X
bWfn8k1oaR35D4Rnhq3o/HvXCWRzjvH7iv7/LX/hQ/TXPEnoNsi+q9f92t8O+5yE
KVLaSh+PuRY5oAZWh5ZKAXcxsr/Qgp7XZrT2yeuXCz63+g0a06JFjdv5WE+uPK3R
vo+FyIlxUwKI6jTlgu3SILEvnVVTm19u8rxMxeEFdeFyichPKqfC67az6OFjUTHL
dVEa1zqJCy+LcZhSf98TpiFIEYKRjt2WsRfjUHCZgKlU9ggSxCEcptCINBGo8S6o
9KzonTg80QTKIVSRHRUt4KTuEqS4cDLv/qfOb7LN8r0snSwDNXcy8IvaIx/kUDFZ
Lob8sdViVq913vYK5oozRe6NG/+WQP3V+PCDdsC15K+3Q7N/wWepaOJvlkwB0p/2
x2+iwca62Eq1g0Vjeuy54M0LBjR1SWTjmZQCKf3qf65448Q7q3vF4NjAz+TOYzjd
OSPHTfSHioJnSMiiTceSk7m0jY5s8nTTsPWOfcMhVJNopf6W83FFovRovPIMKdUt
Ro0UhVzUEJDVhv9LwnfRenvkMTb53D0nL7ZI4SaMZUTMwFYzYIdvOmAz6Kp4YoVh
i94o63YTA9J3Za7Z4SsyCFYhqcZrI7x94Y2on1XSujLqmdJpUUxO4t4KSxjbHUB0
/iWQaii6z2Tk/gqOsfPVc6444J+9VkecoArcr1hC93QUAUmJ5Ei9uxNWEDPsG/xu
YZ7h8lfvJKjRkVXvfRRe/QjlRsqHTb/xfTtLFF0sHNWq7TtuS58dq1/4pKkS3oGK
YrRuJrVpRrE3AeFK5K5RvMYdOd0qY8tfDh9Lt8E2TpVEYjFi+HCY3O2NQjO+Ught
BePtJMoYXRU21B+EP4stDi6RL3ezDC0kytbHfetE8Qhijbi6QrXPzaWEwgWCOkcg
Nx+oWXxkto8CplIM4gF3ud9r8T3So3SbqOGzptlLwgUGTLEjfLNiOSMtvnlluomS
QfbSwQdSY1huzwy+rbXQ9uKgw6yc99dELf64KnQBf+ZmRJRexP7qF3tiO0IkAlFw
m+z9/xIczOmreLEEP7pMUe4gkpreE9aqgjNB2RRPoF7wAdipFBKaaa6Rnip7vPVX
7bAL87CuZ7zRQ5imyMNmgDv9RZhtktTHcdqEWbXa/uF5m0i93fId1dN2vGho2DSo
ycOs8guxNQMJt4ee17Sw/+NLnIhNlG1lALA4he8NLoIvLKJb0Uba/pIOERp4krEf
8UipVnbX2akEdd7xEcuv+iw+nQmSa5jHqRj/WmOg/R6yw0Nzozxeg0GXpMivnbdT
DS4ydNleMCHxYHXUYeXJH0bq4gdhFmrpg2uHJD1BB0FRzSb7sEggM1olpIww3Ee8
Wiw8PLUdnyyQ+pLOILQnrc/3KF38RQxIVY0ccXenDqfRm0msPoVCGF2K0auKWiO+
xdiwjLZhLnvyd+dYJ2Rk1Q5VmCEZR6xkyF+1zclVsOKEb46Cke/RuEKl/ttpynK6
xIDROxUEXP6lt56ouAXc4ic47BbapjbL12JwrDmB4qZHf/w44R5P7zGX0S/Z+n4f
VzogC4GkZu4SJPGFzvpi/BFA3ONa92AXIu8zEMlAQ1ixnJ/SKCu3kp3RL8hW+Kyk
2LeAwqgw4M4eWJpqX6nIq8MEOZG0nQngpdoNw5uVxYYW3xy6lDr2yIAu9cH6zMx7
9X17Fg9L2dvR3EvHxUofjptx/gob2GTdASJTj1jtuJ4=
`protect END_PROTECTED
