`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ybhFFseYgxEgyKy6V0j8YvMFkx0EiJ9aQeLXNJejKzOH9wXvl/xWpRoIbtyBjLo
XF6Lcdr5RHYBhx5bP+SSjY57TqIBSldb1/srQvySG6uHlrgsl4bHUcU/iouaiO7l
BVyL+uUR5tP202TT7/Dn9nH7dzzSAP0C4X3aGE+8vrdekeBZT7k9EkWbmHbO38Wu
SyLnvD6+PZ4t61a61FA+JCbU2xtjtxoHLFlt237mlZa/w2TGgqhKfZcAZ27v2M6/
WpDgxQ/Z1+6NBzI9XhMumidwFiCg0x9mYrmXWmhGyysvbtSuKQc0wWlChP8EjgoO
TCeNJepIE7UIpEwjMebriqk8WsKDk1ovkfam4t2DYKfsIGdZlaOtbJkr4yAS3xiS
k+MCHQzhk4bsejbttkIwuvQW5WHQGimu5biQdys0ALIo6IFQcpvWvqq7q/4/Xb//
CEtZuTkhE+0GQVV2F3ypmgO0v+QtjYczIPgl7tz6jJVlG+6nd61hf/R+oOewv6Jm
LejKWe3dQnsuTXXD952mTVTC9oW+f3E2gZdZMVazv9NSTnfu4b61kyS2VbEj8oSO
PUJGNfjtFDjLiDE+tnZXRtd4m0FyCAgW7PE3507yAmrYlxqY6b+XSocWsK+5+c1K
YGwXq2diCrgFvSGKYC5fRBedkAmbkcO9UkQgFiT4t0T4eS5dYxJ5Q8AFvFJt0phi
zvu8e9pPttV5fdd2njHAtg==
`protect END_PROTECTED
