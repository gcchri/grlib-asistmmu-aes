`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lNH22yFrCbstyOoJIV5JVk8tYHWyp2HLRxWdk1B7DRMw7jXdqP49qDlEgChJp70b
eFmBc+pVfAOC7JCYam24/wvidN3PmAEMzD2yO+49bYZKSNpxtkWWhy16tZwuKosV
rAu39BRb3bbLOMAM1bOItaf9FuxvvCYYijCMeTg1uywEE7WeEzDdsoZu0dYD7x7A
XLCoiJF+oRLpXlKktnZHcn+wSqb6AsRyFfFpYKz3BbdBHt/e+r4btc2oFPq3wfIN
VdcaE1S8SFQ1JEqar67nYGNyWJhThePHzqE/PLdjV4OPfU1NJtzg/5hGgoFCgp3Y
ucGMGSFSd0ak5aePkM9tSg==
`protect END_PROTECTED
