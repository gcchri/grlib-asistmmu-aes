`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F5UOhD6Lr4qSDI6lFTHhSqyeOplmoSRXVMGmKSddRc1mML4HdlUi8GPq0c6hRNfc
80ZZB7aTDMN9ZBntx8R12DdE74ykyqwbGTnIM9ikgOlmGUost1yCZemkLdGxfjsb
tcerWdIPZoEV4hEmaIWrLlkfMqzS51biZUUgCSR5X0ErLuenvVJu8RblZrfRuyxL
8rMFsW8//RLcBMqy/yJLZdQHLHmMxCVliPn3C+8dNaOt5maSInvZmswnmHH9i26I
vk/HIdRgNuZDCzMsI01PsZRShdOzYHH/z4jF5t1GMvA9C65Ho7Tm7FqFcZ7JInh0
lLm7MoKRVXQ7DKgFByol8sGjNzmmoFWUigv0bm6SRQTA4J1d/rcHv/PNpfs6X9Bh
`protect END_PROTECTED
