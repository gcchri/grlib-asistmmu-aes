`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5eyx+dGKOyvS3Wtn+ULGbonchyDoWWa/WPu8+RSTcRyZ4Zq72ZL23DRXkeFC/9TY
gRb6r8H3ELCJR+OoPyIN9Nm8zLvqO/OqiaNjpCjpO86gcuP6M8uqtbMpP7a8Ou3l
mL7UNrMo0Fmlm3eUF9kJIZ0W/SCWhIZOQcsafLW82wsmHfZEU19N54j6VMSuRlPO
vp7yTpJhKrX85KuURKEDVWTh6mlL1OzpQk41K+UpDQaVOJpI/828sBNoLrjIrXYF
OX9zQABUVM7ad2f4/oSamwDIvDACTfHCBpGpicwPRbcTGm1uDvz8XduIQB2ax/Fb
1W6AlH07OFXJjQ6NOkpQuQ==
`protect END_PROTECTED
