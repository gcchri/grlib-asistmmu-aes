`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J1EQCsIRkd3/aYWzsz9xmtDbbOlARXlXhNNwn0tIKUJ0poGaA2bfZfoDtrzKDNK6
GqSGa6mG0FTpw6qqhCN2v42el510qAboV1lwlA203SV2KyZTguCPNXhhSzaYaNNg
74Cyo4tknM6TqFiQchU+p0qBsQuFcxNPuLOkNLJ2ridkpOFCTdPpl1S/SgCPyroi
c/rj1WF6Uhj7tbS3kym/NfdJl7PGoxjYNNPhNoiD6ROl51c0+2udZqxDEN9vdyAE
ThIgHCImg8LAljviDGi2jFJNsfRcDC72AtQs5f+CKJtVrRRYaSoSF5MzptLSLFXh
OaJthn/Ha0VDuXaNGbU3vWh5uKtZPhmd14yzExc239dkkPtHwid2LQ30JhUD75Eo
CAMvG42pWCxiL2B8GMKZgt1qcX3EE2eAHMhi/DlTcYPfkKKkz+xbxm8iNRc+A7+s
uCmYmTgZIj68Hl37sT+cdAs44wfbyouL9giNU/CeT6H3fvBzYyVMli1IQ7ckAA6j
HWQRcSR0/JDC4H80SaP+CINyjIKT1oCZxQdcEM+H2FeQnSPu78zCQhFFb9FSQbmt
F4+7ICYCmwzoQ+r5rw17ZKvlp4zChL6CzIdPTkpETX2cKifIRZhZuJVZvmdoEPcg
lgTUAS1lHyXwnkgRXYgmn6301w8OCbm0zS85J1M1vbIa7e1rEhC5xUtXvZzz1RSq
0snzxc1WqnLFTa1liUILXg1aV4T5GJFwAQyYTIEtRw0oycMAyBVW4wq+nN7yB1i9
sBSzqcdtqcqr5pRt8WoUZQ==
`protect END_PROTECTED
