`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HP4QxaKGog/cvDsJT9I3N2ugMCjg5nnEJxpgT6hc5gn2cRp+A6HHaQ0Q/jX+fYS7
TDc481unqfru/JUtkY286GzyDb94ERvQDtJtn+TXTJRAfh7x5KFh/oJoz/w9iThT
Nqg0jz2bxjY+2urM2NIM3fezWup+MDw1Z11333Cwp3zlPhzTEEfpCPVw8GbZ9Oey
1jk4VVO1Nb1Os2qFXTMWubeFQJih3YPwprt5+/B/EYPM0LQxrg4+1zBjE7nHCncf
pmqiEhSh64zNDBZxKQNbfCbeGyUdPujFXUuPqiBSQbIgzyvNCLZCzgNCqqt4ikLY
Q/a+TlxBDxXfp9ciYiXcykQ3iyYtbfcfoDMBqtcHlsnWTq9o9D6sK0YNJ7m5WosD
oWUjKtQJS2Ndntzy14nwe2VIFCnAerNoKe0lK0Hioim0UCeCUfVZ/vLe8f2XWQqh
mKdV57uPKVFXT6XS5u9pbAKz074Kk+eoiscg1FPp6vySqw1MEPTSNur+ZnMD5N1M
`protect END_PROTECTED
