`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BkJP+R7sdOagxLqWQiPcJajoCAVCAGaRsYFPGXJepQdCydVAa6BqJ/fqdRPIIBh5
D1mvmWeK2qzS+CSxfzWk32C1QzV9ZjI4oANfCHc1u/rowo3NMal+BLfFUfrgHCoZ
t9Vz3SIptOCOTQ/y+6tyxzltK72YVCo/VxMFUR7s/7Ol4lG6v0225fZ/fBVMfWv5
3hUgekhwaCRRIAxdo6C6HhRri/LLNdfZ6ojyYNO/gvkMytIE4JUPMoL47w/FWzdx
2o2iBYKv2f6p5r3HVxY1mXI43kVvbw63A9fEvXgtvi4PAcb5Nh/lTAGQZnDH7lqL
F8XEHvDGm8WEDOWFh/ATyjznjqXTjT1qVaKhsiA3IEz0VfuiLjMeJXbCwlHog5nF
3ZerFZ1lJMnBD5uU1iyCnADSxks4zAQ6YvrhZZr8sfW4ynzKotJ8xGJgM5qy473i
`protect END_PROTECTED
