`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0LimcRjHoQUtMxWkTwxuVzpjhXnsEawrcQ5XRJMYR3qpszqC0xXcVg17wMoe+eDX
rvqRS0ZJC+VcqWD9G3YDNsyu6esSQ1Sz+j1tXhPUlORzTMOYMtagkanfDkV2kCGW
VGV4yq2k67i/e1VH0yTMO/T3S4NTCVqM5UJSvWNh9g6pOLXQw/52VhtA5atm258x
jnf5y1eN0b5y6ZKLatJd8ViFqDq63Z+aQx3K/VLSWzHPxf/tkZdRtdFktzpQf+wq
NGycP+zydtQodoMMkYJV6svfaDGA0ETrhx91FxoChx2elHvxjOGpi0dLRS9Qc56C
WU8FFg/aAJW1W3N9YsmXZ12ZKLPGI1uq7bwQZEwHva6Gfq8QWkDmdDEdFQHgsVlL
2H6DTVOAdDBX8Mmd9QP48olY3fwQnvLNVInvJ3PBJSQWCh2k5ozUb9wb/q0hZNZf
fyMrFoBCPlfq77mpwlKjqzdCUcPZ8P8kHswPG9AV1jiErDCIhIDjGjLkzwCJ2xqy
KYNVAIu83cIJvZieah0o8ujLrZS7KlCnq4DCQXemZZdCXoYOwd9m+W/rj0AZtdIX
5dDgJH6Z3cVYf/ageMH1cLb6NEyOA5sUnsHroUjDPbYkT6icIfJO+as9dce3DomO
vqAEktxu0LssPGWwl/VFPm+7Rdt/Xtxi7FBls6dL5gi0qhNGE5iXQjMxjkhBlPyQ
sojvkgaKoIoBcn1AvP6id7W+uoFh65mZ1DHlgoZD7zHQh5QT6OuoQ0/W6QPpYiwI
R5oIMDbey6vES79QweEWUA==
`protect END_PROTECTED
