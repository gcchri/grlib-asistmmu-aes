`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P13oVwOOU1WQPN5HGtJMVwst/a61EenvjeORZMXL1Cu9JV0Py2m3P8PuQ9F3yHAk
AbmdLjidCI6hvmwP4JUj24/9od9gIhg7ijLW2ZjfpkzV5ZhSDeqbKc1ujfy5gjOk
axs1x7ay+5Tqra7+OhIBgqCwOQiKh8Sz+D42D2ok6JT6X7l/jDdppY5wBJHDhFmp
pSZQzInDrpNpXRXrorKFTtpN4VQVoNqe4WN9FJnBnRpbc7QdWFhEDTo+q43Ku9wY
ieEEhPGub/mWu3Ps0/1/fpm0K+30OWTzOSQ4w5UVgUj+bpj0eUPhlmdBfdO8vVmj
jtFuic9uFI2VFqCfYyG9Wj9pwz7+coCYxexQGBmWGE+sdo0C4n92XIzT6RWuFJT6
CYS1LUcZnoAyVkvCfzvHPRNYJ7E6vV3vHXCrL+Pg5KLa3nVC0ilKGrlsuW2OvOj3
rTDUD5za1WtRtXFk6msvy+9AeSXzZGqRf5fh1Lpb8E1FsFMwV73XQjxmunSrFf+A
XYy1Qq1agp3lE6EPYVYELnPSCTc5nHpnod5Ye9w6O07BXMewveq/lbTwQp8+PMkU
J9gbj5N6rgxCLjLY1gkq/wXf3V378cFcr+YuKBXcVx/eaNwk6YF71FODt1Dx8zmi
R4uMYdFcRHLcxcJi+oQbAdIehL/1ebzBqp0FzmIaTZwqwdntMGBNcpmnph0AKikc
85itkJ3D9pCTCRY/vL1K6z1lAJFbLZy1QiJGpNkm9HF+QmxfF+iZ+ZCLbpgDFLj5
XU7nxqVuknqwVihoKLTrMBX5+cD1Pyl2+7S43gmHHZy8JngpyGVXM530dDoIOgXd
XQEAbnbLwHOeBza8RYWsnhbbPocYLn43BuPT8n/Bi5ewOhIJ75Z4eN1b7IvcIYeV
ijWodYaWsymMnr6QmKt9s5lTzpDqkPk1LUf05X067Z9s+iytwfqZZD8DMH8teHCa
m32OC4nhLJT2brktFAARJpfCAWpMLwwKmSC1fKvDvN9gNX8zV9tCnk63aNolYDl7
JB7ClzP81W9n7YTvyz+JtBnqFWA8HM2yIQV/+h5vV9E9JKYUasGQ9qGTGDcvgH5r
XPOv3YDQQ7Nn1lOsccjDjpajzJBM0/dp2aVp8IqRsnS6OFIsIgpAZ4E/NGH2e4UY
/y1dwfC5vspjEixeD05Q0GB5h0lbvtYyg08gJARtHmCrcYl0pdkBD9yc9vVboTja
YTVFuansafQ8RMAukzhA3UTQxt7SjuT8ckiakg/boqmFrGvxdlPgTHynL7tqB1ap
y9IG9cdM6rptxfP5W28O7r0CDNDaFMVfOL0DZhxqp09mRPGGxiZZZUZb094YRNuK
NJTfAbUG8OSNo6Ayzx3lyGcQ0AYISIkXNF+N+c9vlsiP475gu3gKUF745Q2CUrOq
eggbkHx7PHZnqGXMyWum1TqqRX+0ZXJmmSb47E3jOwbwh3gVI8MRVjxjFLG7a+UR
1FFSamhCTtf1q+sBPCioIjy6h2Lw5Lgvtl5BbJxvsJT9lQGJgkbIXMjQpaSM4ong
kDx42CPcYwL/zMndRV2zFstoodlKWWzTCMlBGWBM999bJBk7tIG/riIy701jYFTG
TCapGKOZ6EcpPVsDTGn/romkaMHPgJ0TdtgIVotNojosXUe4w5O1LpYl41M1wCSq
rXn5uvTFc/3JgYbzgew9GTRxCFzeP3emTL3pf6YVEEWkwdIX0yYxSn+g4ZeudpoV
aIebfrHQnIMdGmKKum3+HF2BLIWTBECqvvA+KMWHo7iKmGT7SftO+tNrUVcKomxv
UkNuKPw8r+hKuzfsHbGT/JRfblMWnux7uYOyJUc3msBKZxGri77AbNjrgQ2ekS+Q
ANKYCyUl0jU8u10Crhns39S//X9GjDJxVKte5G+VVTWFkgedE/lVII/d7KeQnj1B
CR6ESJ9x4Xp1WfY30H8wgykLNitoHKdTdbQZTFnf59EDXB8g6EfVSV7OX4HHCm30
ALJwPQ9xYMSOuh5uR1ylkIK0yMvIHYLwBnczii0KWH8WQ/gYnPl88OsRelJVdYTU
ACo9/e8jgm4B7uCZ/RoizvQGreTJuy8I+WyZ/GShuZ5/CNxKi4tSVfW3ajPn5cas
wCDQEQ5NFFLLJWWf+yxq19gpW45LVtGAuXnxX0Sm2Ty8ZgTqoMkZTlDWNTwUr5s8
bdvhtFnrGvvzfe3iBi5iVsHxJ9SUxiBgj97x4pKDrFNP8s3SNKmAJtKr3Pl7UC/B
e6b7dUp1u2gc9q1Xmfbt9QEEoYvi573uzpTBhg/jcbDDvx6RzzDdR1x/6LP3VG2M
MTXVH36Plhe/l190T9KHHASLZHjED0bFhleoYMaaMwO1UjnwovzsBTS7cmgh6h5J
R6NPUOII+iwMs7KXU/BeAdIs/gn9DZsNqGK+KOeMJj1LLFd3iWuZUE9/ISeZyi78
9NwHTxMQuk8+B+422VFvROYGM//ZAR7yq3UTkW0BnVhNmlNo1LYrJwhj97o1C0Ve
Rf1DiwYgJpo469vUWYrI5GdqenjIaBUkZuURekYrWvTW1pmMmeJ3jTUNR/x7GOnJ
PVczqSP929Tq0Mymxha5kGvI1wZNwX834uW4f+k4ySYsb9BuGfm2MWk7K7aYWQqD
aCq/P0H8j+RQgh8ZYpuC+1qmh4zBkQnzHG+IFIKq8tSj/Vd4WyvIZXIoMe8yXfhX
+XpCS5LB1N6GXu/Bsw5usCeE/QoUPgp5vPFTz3pO4iXYazBwz8CaCTxLSrtk+7xj
7OJXZ1pQwoloUJRZ6a0z9p2K0InRQpFk6bydMmhU3iXLFdPzZFeMWEsSQCxfWK9w
K3RukgTKjSFD4/BmkcYulL2RfBf8cKrQLkDP9eGZpEHYl+8RSjjrXqRYaCv/kP8e
NzjteYPljrIsuBITxyKTPRQcKyvs45brNBdpWr6wOgMTxQzP9wOAjmy7l/hk+Ttk
zcOGt5INGHqjovaairQyPGxXvnQkGyMwdEgR54LTQFGfL5eVAdAOonh381EnR6wx
zb6NVB2JL1txmEHjuVge6FqV9YTtyFGX8O8IAMaEv2ZPE6ZebaeraD+4M6xrR2kq
q8ZW0FXaCHAQf8adoMP63kPHqiGqMhGEZn+rVgS8iWIjVBadh7vLdvMkQK1kBYnu
ardh2ihNbdVKk6PKhAVQfOxsfoFD3t57RaDc46KFcof/mgLaDbfHyLEXTHnX8dNV
unytvyxW4An9cdTN22yAfQ==
`protect END_PROTECTED
