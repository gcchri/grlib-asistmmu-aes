`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BA1gZRnCQv6IPPKOG1PXmirdncEzDgeyylKUm8kx2aH2C7QLJfBGXFJm8pJjkX5A
oESxjoKcsQbRS3j2MLy5O5n+eyTfioK6QBS0BHNo6Yee/RPdc4weEMYgpI4zzvkz
cK/RbuHQ0ebi6AvNuoVjDM6wMr75yGuqHH3wiEJw+s93mSXCKBMNT/E8ncaowrFJ
7231FO8alchjtKmJbaungUpgmiGHhuXq8mOY0wgYPOkrxT4r+ibvjD02K66tmzpq
E7PJcc8AzdD2dCfK4PG+OLiuO03CgYjKjIiU07Hhnh0UV5S/y872rbHIXNYajGGG
h/E/LMpcrQbirJ9xm2JddJe5XgMI5BRoLIjBNivwtxxfDRWHENX8PJhMqztY60id
lRsmdEjft999EODg6c29C5IpnNlE+s79Mt3D5uv1BTv/Lpnb4Zd/GQk7+aN9zgAu
aukU9SCpyKVQ8/2D+NxK6XFVsSG+gBMegKxPtwejLraFxo2Wzk7a+GI/jfExsgwp
0CgXbajFBVj48m/wmeBqCBfbJMLoG9NgUkzFya0jSxl3wwDA1KJ3OMLWOiAd7fCQ
lEYfUkDdiAWpatFbPRLDzSRjKhytgycFj2pDgtXlijRHdd5Abmg/7ppdZ9GcFHAy
kfTPUQdKcljcYsD4Sf8o/qjtlw906XzaYfhXYx5siTWnDjIMlXDD33DtclJM73Y7
Sp0zoTURkjGxeK9G2alJweXm4VkCrjH3CMAK5caArpo5jwDCnXZHs5QAIHctKRrX
0cnbLzpeEvUEz49Vyx02UV73CcD9rZOsbbIn6Sgcja4tFrUgqspXxa0jhNPR1CPe
vQyCBmhTRYc/K1lyzsA7loQeXhqyg3TNEAZOXBoy5qByYPkvR47boS5I6ge2hFV2
yypfEq5ZKyc/WviA6EvFnq4D4XE1w9LJ4dod2mTYqIqtN0oQUgl1uNBuCAdzTlV+
Fvtzyz6ZhZYVqttuCG5YFRUEL6uQWr+MGuletVncnuhB0FbwEwx8MJq3KvOBqz22
gmZamNwuA2QwLnbbIi2ZHU6cSrMEJx3cPtpmkGUWrJMae9jypP09SLwambrqISfX
G+UPXu8S2lSXlkehtI4bMzHoaA7Kpfk5pjHt7d9IwMCglUPVEkg44KpuYzQKlTHC
9omjl/JfY+6YQyTqCRhmVN+Y9XzSYqf6cJHU4MsZeCOeInpzJ5jla3+WMpA91Sq7
cYwvUvMDU2ntN3pNM5o1eVmhuF6GZdDi3bZNZDX1cXXqI8IWL1nRjsYV+YlbAU+E
0mjwK9jKjjVBs8cQqTINmOFWtnDQbuw21rnjBi7Kz9/BpS1TakGx7LnoM3+VNxQL
WmknqXxzAK2sf4TMggp7nQpaDqmZ8Oqerq7Mb4rmp11gFYzm6HejktcS3ah2Q/2B
SCsqoegyInBtIxeoDadzOu7J6M7/Q5h88cMTxe2zNTQ97n2s911Iu592ypGRj6yd
3lyYYpVjGHJkBkLH7Dg7pDum2oG0apYGfiRS9SpRGzRSOe53DOLhDDH1HTcPkX3g
V3dh837PNCkYMQSRzcvfhYe9pyXjP3ZElfmbvtAt/WxzimjIJfwg7jur9QqIcYXO
G97TKnR8nv6JwiFXeY0cIObP/TwXkA6sAEFUWMTNqtWRjgFKzjLaDi50o2rxaV4F
kelzWpXecVzb5XrNk1IdXvpghphq6qd+Eu06nUU72DjCce+Uxzf0um6bH8mpW/kX
WSKc4CeVJts+mNDOVw4//q3aTKv59ngo7CUIfGJGPZ0X9syzy+E+qNoHPDjJFG8G
FyBUeY6duf6AhPHpU8vnMgrSRTys1J5Tx7tk0ZIU984vrCaI4bFtbNxgzDVKUuEu
qUGiDybYxhQfJANlug8gv7Gd+gjtNURNlvCF1DftZj4sCP//m6ilSNXTmJEYZemj
PDa1P67GRJRzHD83aN65B/R3T49qzroHm3JD0IDvQAWTWNtpkVuK57SL0Ea4jxmt
T3bbfOIUKgrXL6b0x0T118RJHPelB++Lr4aEldOQsetNWSAzYRkfRIHwTZ0aE8mr
GJg0IPmMywMF8WZniLm4hhVUqF5QKxVJZrqhbSrr9+vDNjHimpD16fenz34lyAi1
nQbFpbX0QS2haRdf+6udWMELIGbJNuyXvbq4Evsx2/lkoyIm/ncoI+qpc5im0V+V
7zqCqsS4rrt7NCuZLvdKd/D29JLBSR6bfsQ0O+B+p1TmMlUqCoZSU69SfoWbWs2m
VUFVRaxltPeJ141yZE4bGi3I/I8CbKqLRvxAvOg4g2ZXdsKUej89BQ3Lz/EXRF//
RiM+2MJq2G//vwuEhui/z1nM3xtp20V9lsCOsGR/HaWMPK0/E/LQGdkZOx9RBTKj
jQMQRRFIGfrtQrZ4l4GZPVziuB/TaDNDi0g4S5zLhvu9Oz+VLcs6vN2FB6PqoApF
nHHVofEyrR0tHZzBRqsgSqhmqw5ejwC50iPlzIu9+mHuPPL63F1ipQMqIhDhZy52
ncBBS8c3nG6HnvaXUdIM3w==
`protect END_PROTECTED
