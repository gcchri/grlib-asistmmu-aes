`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yeb8uG+JaT74QjGFb40ACyDXx8WgYmXekuUP60YcoDEtEtEEN9NlB3sLKGbkfa+L
PGNspYE3zN2TEgVAxwxLKlLmnsGAL2dH7wJb27o/IAG7r6WjgH4PdBtCcdjyAjrc
gxHW4SHlPi6ah58vHGkcyiPRYvnY6dpasLUJrUQ8XTR/wgKn8cWjebGVDIjlITOL
L5rrTo/PwOLdn1ifJCiXQhZrCRmV0dlShvqHkVbgfy5EnwP+Zd4olzIhwwAvgTNe
VTRwZIV+b2VJafijuC0DVWFfNd4qxDbqFlqDUs78UE/iOewArZZAXKloGladqA8k
ckwQ9VTsN88mBf8vNZvUhKD272KyLH2N69mGHoMyxmidhuxO3e34AUUdWAdZZVE3
LV+M1NesObG6OzqtW5/ppBa5uV+SJTFFrTNo/+IUiV9CM3q9N1nLJHjYH5f0mqA1
L6A3rYoI33P5s6t//MqnFl7dQtcEN9PmFupxJJdHBTtwILUbR8uOA0q+jXzXAI8O
Hsof9MtPKVeKLLoDaiNGonQ8mA0oAowOCPVI+iil4No4N4ERqm38POtsrWME6Gk8
vXABcA/MsH3oE9MaoL5V/k7xzzbb47biOfWMJiUQBpSrHC7ZiNChb+1ArcTpRanK
PVIeLLWNUcZT1MakA2J0LQ==
`protect END_PROTECTED
