`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tL90rXCg5+2eXRlJ+h4ozcO0bxlii5HMIMWcVldCG1i50AUk95VfwnO2GxdmUi3
ZWSop1XEQYkUaZzo6yPu6AbUGgyCEpvuR7eDjTfM1UA+lf1nenpnP71JduXF95jn
xIh9SoVtpiprN4MjnbMbLXBaR/A9wJ8pYyz23lBx8Hfk92CErpuxuB5gc/VJTey5
hQ0PXWpUpoibX3D40uvDQMTL3fNz0rxRs8E5Pj71Ky7cSrOz67d6tHVZIXtXSorU
MBoBxoWdbkramM68fKICnw69Ip2svJXY1QG/rcTWTdeERvF6T9j0F+ZyjjGG4PTw
pka8gKYyT9G2mUyjX7dfQdn+B2+mpyBg18Fx5XbhyolarTJ9IMAs+CXstY3PK72y
3S6obeUf2PicwurPJjBWOaYMC06EoIyXHkazkq0ke9ce9Zl5EH9B3WxuQA3KcH+x
/P2z0uyHHawTBxKFYWQTQQ==
`protect END_PROTECTED
