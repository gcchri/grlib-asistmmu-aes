`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSTZIdNK2MkhWRgFKuSGths7EX7e+qlky9SLe4Ghxgid24s9qg9GUB5hdNtaIT8h
6Jn6R1MZoxtaQ8Aabk6zLgraTm+8L1UYZFsXV1boe9eEZYO/n5gjZtziM7sUBfD9
emhGgCsb5GTYf90NDpjs7cPbOS1Vul/uJoVPh6Jn3FaG5+wx5YeiMC5mcpMYlkRA
InsPrPtseBRjU8vPmP3T5IcUIbJ2wB/74BCYHgHXMCj0gJmhSpGxSzfYfRaBdJTY
KphUSXKKsbZg8NZpOG1lt2P/dHD9krjGYVQhCKGfOzoEdx2WgKftoBZjzOS6T9Ez
ftErDvW+10jTLZ7QZHnRmQoSF1bbuB0vFIP4owBXGJKrzki/azwicL+w0fXsazPx
`protect END_PROTECTED
