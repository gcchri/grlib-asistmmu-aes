`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AY7b4RuwXSrCIFcx2gKb6LfcZi3xQ7XcJnqlp6gP8vEgwiSFIjJgRwAbbepPDjYH
t5OtrzQ+LNM4NwEY0PgzWJ/Hcji2pONfVFPOgbI88wrtDawDugGpCJmkdA5SfXN8
vc6n78sLZNM1B2b93L08tlWMhh7lPpggmp5+ypWCnGyvN7lsTBEPUWGyqJ3wRdyq
Jz92LAyBjpAmemefkS9PEyRVZWhaG/qCUZnKjG/xRldxQUAr90Bc0FnusqdL/p1f
kf016nK6SsMl5Srx89pBtsSMFTlNdopdRtncjtYX5+YHdO89wxxle+nL93t9WDht
D8gTkE2n4VpY3UQ08yyiWCwP+62p97cYW3T/1KqNaLbM2/bzTU1MX6rl1eDDcMsg
Y2wW3WaAohCUPaKHWO6EW9Zf+uzHXE4gFcL6kfp6DJFOVxwCvbs5PBqo0bh8oAr8
PFR7GJJ8cA0V0it0oooTSmqk4ZEdjeSs0tzgZmyG3o+eBDwVyR/aCWAyzOvkMjKp
QSkVyxGOLuhgtmLilqQF79vcuHWScwdvemLcTqztICpeu8U8OFmnteeC61B1p5bV
bVUWIkRDnecXIPx3P+YupX24vMF+vtc96G/B852vc0zsmFllshH3Mie46e+bJnL9
X411eYSHj9zryzcQHxPA2mEznlAyGkRCOlurpGnWm1hBgBpN1A71Qx1GAH2KKNBU
L+DWu8geDM+K2wulKGYdloE/5e5nX1vzdcKNvE/7/LvZD2uTMhrbW/7YYOd9HQRf
YaeqzYjm9q/u+gr68Ay/8aezffGS/pNUjBTXdtZlm4iq3AVCjsIYNUM327gCvIfC
p0Aml4wZJsTD4ZYH8pwjSU33sbfx+9Sbhi89qgtQxLJOT98rrhYZiWjgNOZIHLAw
l+b+KKkzjFdTHAOVJ7BChn7Hirkxh/GIxgWZCa+Q5nSH2UO6GK/nZwjpRVEYcKGg
RXpqyVbqEYdj0tBDv2H8YL+HDvmTHOJrSJpHimb+XlUpkMAxK9n2suUehnMOqThl
Azhk+aVQBN12DKFu3JTkc8FWjFsHrkAxs1UXOQtTyx8wvWyCE0uLppFDwbrdPfD8
8CT/o8LmmzoBrX1f4uwekcmElpDMB5X/fWkIFYGTiUSjk501ufjBtqQbrI1G8mr8
I6nabStIomhe2jWzHtuEtXTcn0IH6FjrfKH76/wopDf4o9vxFYAjdQ6pR3wd1Kwg
TLI3DQ6D6++saShXPA17/0E8kG1/+TERQxKcbouPx78ipQBAa1LZ8I+0goJXvWg5
MVrr7b5tM74P00bJOm2vjJvGQp9mJ3uae1EBuRWwfB+auxGkg4+F3U6rJoGW60JN
76cY3aSyp4900RQcf00g0M5WPKqNZO2ziohQgvMK31wB5BWoMl/VfnZHbHyDIsdt
v71rW+sYylVcm8k+MwATliITDUGjwaEGoW1ANXWQCJeY0M3LlRNQtRRsc2PMgR4w
QIK+e0I7jDuNyfqGTe68ag==
`protect END_PROTECTED
