`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmAXiCMTSB/4RQHjpND4BJEJkyazOIaOjf7hejXtxkpS19MWTmKQmQSN9/49aRny
5kWtXwFJVYCtaf+jWjuwKlnc8o1W5lx4toaZqnURfIIB7F9HLvJTcuKOXm3Es9RH
O80MT7Ayno42Fx8+9aKd196p8mvSpyGn0jf1imKVvpTHqPd6Cf0rt65QYhgWNoW2
137ULbioaJTZATIEW6cwfP8eqmFsMN+6j7ZWba772Khk2RUcWFlz01qDXMWxifRe
HISA+H1Iq3hYjTmzmQlwymjHD6xWbOd58kYn/XE6c8ZIxKQ450nQyRfGeZIYrGfQ
bd0CBPG5QpgkXX61b0b5175tnezzwM2UDle9A0ddobEJc9isl7AF4H++rwO0eEy/
p0//QAelm27hOf1clbTh77WXxaVAIcqEvuXGoSYarn26nKN7XVCmdncf/aHPJ/5x
PEmnedfj954K/xExdy6RzkUP2urE+43AHnZwUZpWt9lz0fV2JNPN3Tk7btUW0GIF
+Kr7gY+it53IxXrXz+fmfbwXsaeVt7d5ecsaB7k/YDdgJlGgOq+NJwcqYSVTNPrW
t4Xnty0C6F+0p34hql4+gGcpi1+qHNfAzN2OeaOpA/602Bp4Yhgy2I2UZMfa95AV
yIdolKhWHOsi+LX9XLumvziOTgHcLRrqNrNvcuzuPlFmekVxYF+2V4DXlxw0covI
vcOcM/2HIv91p6bgAhTvl2UdC2fibPemZM4qyh/TAzp+FUFFYRjXbSNip7wTOhzM
uMuy+gOGfS9fQBb642VjKe5qV8tSZ7SuBHe1Kt8DE6pW7uXWTst+gsNWAcRPhYxo
n0jORstXQ51NHFBx8CIqOoSTNlErEApY9mC7v1ejrcEtWf0OAHocwbAp0Tx+R7ou
zMG4iEtfbkvoEVWkA6mjgg562HRSQ7AG9rmp5hteF2GRM19X9Ju9msXTYjYIG/OD
+NlZzafGCipRi7aqoU9PL9k68XH4+T1Iw/OyQteXX1iepOmHq+1BIo8WlD5SKy8W
UFFHMBpabDAklJ8Ag7agorPk0IiW4Sbf+DPrcRTRupv7G+J603uy34KeuQjdtcsv
xQDzdFkTrSr3QAvkHCcFAd5AwB04pQZy3P/6ohejWA/OJa5XSX+CgPH4RGcyhwM/
GQfPKLlIKCUQ/sgN+ZjpEKnmDYIgjjoPIG4O+zQv5EpLn01+moaN2+MFklAdXzfl
4FcGNDFzF4rVHuRPwwZOz/koTmtFlJ8k7WjC3aTK9AstXZE0mR2SsZyXVzZb4aue
DBswlc6NDLCxzJq5LJyF0JTvlUn8tx95VDjHxiD1bnWi9F7FwWiT/AmsVeS05kSA
pdcDksZogudfUyzbWgIuC8618vtq91bSEsDGxi0RX3QgLhHhJDf+vj+3q6il0UQH
qJZzmTcVZFrsRt2nDa922i9VPuqeCngAkV/14Jedgz29TsA6hm2NuNbycNITyOlL
jV4i4XIqEquPo90Ub2L8yPx80vnIRugQukcI8T/QlmqLZLPSYVpfiozRVRNmFN16
Xkb3/JGqJUpfmfl68mIOfu9VimHbfbdBpIlxKM3C56pf4XMZQyks9ngFocMGqebN
cdXSvg9axIKuA2UQ6V4vmJIfQ/OUpuLSl5FhsqBxOm/+gy+TsJhsyFHkni9MlfNq
KYZ7JnW6TVqPJT+8eHDR2Yo1Yn1ILaMjhomVgGQ0w/1lNZcQJq3nzzNWmZxcN9ec
D1wvAt1hrHVEmoxmVPW1354DQXhp2EVz7FY/Je9WhAPHl8NPIs5IwgNgMkdWrmFV
APlW9dayCLcBTCn1BaUcBQOykuZ6fD7DY3lufE57SCd1J8ByxMVSkq+SjNpywdAu
/jz9sLl+m3ZI4ZE89HnqHGkU/G8w6uVnvIM2TF/6/lQnp9TtOxSSUxYle/t5kwrO
7Dnpc9/yqPXdgrwTUgP64isyIzQFO4VrWA9gLGtFi+ZI1pjeEBS62eADqja5N0XZ
j0WRw/0TrpCLvlME3Tk1vqI/Y7tUWr5O7kZ+Nv/GO5R8qdIhYqZeLnxoF2VJ8Y2H
xU1cdkOU5owLd2+7fUGPqb4Tz+6612bUl5bxYteKl/UPY64BRWteCSZLiz9fASTC
U19z5ZqIftbm8nzypByDd3EdxwL2TwEZ0SXJEabUTfzzGgberFD0vU+XJlhQKmFY
OKqbSJhg5YorENQXD1TWJoENyfOAtARIKMVVMAVkhvKrTd0LAQitGvrntdbMzIWX
CwG4rghUu4GZliqU3dL/3u56zYYZjB3X5RVjxv9hq76BB/DGVUSZEVxu89wyNwDS
8ulsOWN4sP80XyWsm8msVaKFzBuImii/w9HNg6wnNwxDAUyv3ZUowP7eGOUdZvxn
MP/cOz0Fp8WegeH3WxsGISJ5DnakIQTECT4GO3giNX8/E42uISMiRBvCPrOTo5O4
z9P+6kXl6+9zoyoq0N/jUc56ns70h1Zes/8mkv2ZwPMl2jiJSdTavZOyPQdM/0d6
3r8LkuncgCYJsMqYQ0ktls8xKZ4LQH9NflJA4INqmjllDgCU46/QayxyAtg3r3+z
AIj5RyjNN0mWBcVpuPdwlM2HCYamG2I9A/a6B+70q8axZA69zzcC8g+bfDPVu2Hg
/k6Pu0c9b4W07XOqlMUPh46480CGheCx9VINRRJhpPaEsGp7p/Nih5laGakM9fbJ
bEIDiYUnM5CooKqFvJmIvCqQvLO7equW8q43LMr47kxw5ZfqvqGq9Scgn3AQUzZ1
VW9hqhECwQcH/soLQwodUb6JjUgeIyMD58QVC9JlYZ8oruiSRwikJl47fS+2EUzY
KWgMupaNKmwxwfM3lAKbE74WFOA128rmYzezrX4N+ll47v7W4jHefj8HQKBxCUoa
k4CM07KBYgjcNxn/im/pCo5qa42sMHDTyYEaRaTu0fZvhO4cOcvMcISJjDAQUbGI
DwrQSWJ5nNKjn43YEWIvKTnR2LERWmS/D5Na5yAnblPsVjLudalynyLt/GfrBuxN
wqbjEg/YiI9VYtrHeyDaeOja56MVvzBCUZSNRr9MIxHaenH4aHs7005ZgfvmiRc5
yojcXgz9S/tFUjimzAe/WQjLUC5EEa3k4Wq6qcw4lKCLzwmJAInnd4bKEWnDygfa
VB+N6IEC3wirJdzP9S104bmYCmHUUL7CWw27pI6i2kyyMAD1G5iMgJSi0lAJuvpK
8+Bynfcss15UOA+IGWIBfLoAZJGDWnsa6NbFle+iIrCWDqmc3dy0PN7RZzqYGnWO
0BppDkkePn9b8TL6Ke3iHm6Y59uRU/jzfyj89eBLDua0JcblvGF0njtiq9hflqCq
kq4KGy2HcFxb4/mR9J0y3jqQ+coL7kP5PVXgIk6mUTPIN2vbcNGPRPwCDO89aAz/
MNvimjciPYMT+sXa+/Xfd2dTOg3lCz0FmlqwHsyfZrbImTqyQKfabxjgaRjma4gR
1v4m0SELyifQjrbMLyeXmzdY8YbGvKqQszTd4ZJl7BiOT55t5CYFqxAerF1ZqnWs
hiN+8ag+iwW79VSqkYgImEAjx6p5fFkgeMzgjah+HCATNzjTVl85pEZ1XNQ+vLu7
H9bycBm+AJnFp+wS/yaGso9KQaDZmEC3qQg50OTPYh1I91rGvEcwlLqgu1lRQmBA
l0PAQTmt60C0LpGr57xAjNslUjfLWVQRIpwYYd7ZD2Wec1cUSi3BtmUybNHoo2Us
wE/mTrk+0/gWZTMtFK79W40+MD9OlK2hxPL5yl449pdFB0Wg8bxBxULU+jDkaO2W
RhGYxXXKExfJZq/ooYIgZoOattyRnl4Cv1OJycAn8OdeYjIl3NCDeqTafLVTYwtB
WguXAkBDECFFau/JV8rGzsQDtEXn2f1DrxRSdOd1iqB4XOPCHONp80nlONOp82EY
jnqJUObd3qubQxHqSRSz1mN2y+ngoUsHbkeKM9jO7lubMU7/YkYPJ0e/aGBHA7Ai
KiYRoZVm3I8Y0SaXImRRDAf2PZSgPvmliyLw0oRQqoNWjfduhNmyk4nlJconfKb7
TE48JP2fSySjuZs7iNGU9Kb/8BDEv+BUjP9UGZmsp7unhZumlL+AzwjtV6OxwvnW
E4ga5e7gjDHmBLZ/b2FSvE37fm9L+Se2tIpU2QlXPGoCRwsK3MDpoxXezKbeuAq1
+LHmGhebJOJsEljDO7fFl1Cy3JV6D1uxyRcZHCITpDl58o7i2KH5/DJCl1n/AdC/
cx20bDiPgGjBWvN/w8Vvbn7yWDGSLFMYoeM/mfWccws1iBBAciFh5kOijDVx+ozo
RgS9wl9oxfSvuAO8tX4rIuoakI+44jSN7H531qy9gPjqP25MLan4nGDOSA5qn6kc
gL2n1jFxELbRGdFUcxke6OHlsZH6n4hi1mEArB1aGLv5MVs8fGW03jddkxeeQkD5
uMT1ehc/egWmnwF4agcF3kWm2Yfx3gGF++agVMuDF82Uj5mL727lYmsmeOrTtiJV
yVJ7rlB+vxS082ZOwydZCoYZ3JRcGzRqAEfgH98JYupNcxNKOgRtSTwivrbjkrVt
OVRZQcTi7Ub5e4KkF7q6bXDjOoOQVaeGkoLhEYKc2yodBTaw2w2oVr20zMd5+j2X
j81sTYlBqtR5yTRLH2BBNzjUqyRvn2W/CoxsCpPfBZflodl0RUUokm8RiVKyADqA
e1tAVAoN6ks7vKfsTZyRL5VYGQBqopVk1GKZE2Y09iVtaHXPCHggp6DqsfZDg298
GCO0I4ckbYoNZYsfvhML2hQ9qP9dwvxBroWzE2nWfDo0Xe8yP3DR87c/SiXpC+Dj
epXv7xfBaw5M0aLO93xDlJX8MvMHskdOTFsMjtYjBljNjYNg7PgQsXTIvn5PYWtF
8c+4K5H9DwGb71g0Axn9ybVVZr/SlLagg11eLyA0Tz1fv/VCHvFHBJ8buCPcUopw
EPfFJO1h6v3GJwy3D9tVyFCpd8A0cbFKmy9rLiAWXi4pxADy8RhxDD3uUBjD9gHI
FjHjv5dn4qRj9//M3hV+SR2zFvB4kdM18dMNn7MkrIiKlSAxIt7bblnZczV7ZXLn
lULEX8YhvaZUkycNMyCTMr/pzFWkcGW0Q5AKW3n82x6tp7sZdmw2KAyW9wrMpuMw
SzoTZO3Xhi2eJV9RfiCzVJwM9d7F+C2G3Tx1ptYlt4ttvAtA/32sOOgxkmZ+aVmd
DKYToqwhMqMdfaYDVfvSV7Jh5zib8u9+7leyMVTI5MHujEYLn5SeueBQPQPxjbOC
zRiRbVGZ5u60tOIrQECyn3081qHZb3MO5qXfi18d4QpBmEfY09lXGGHORfVdjoQ7
Hc9x2uDHdzdE6/m225Ye5rV8WOfeA1p7G/cZ1lzq0Ykbs28WLREdcvSz+6Fl5mmT
pG7jctK7NUE1032hDnB5sGKtzzi8EohaoIUtxnIc2TZt+pxg8VWd5fi81NCSt86j
BQCMvgjBU3aiix1C0yjBpYakpqgOiovoBT2P0TSd12xdE0fGgVFX5dQRb+LSZcEI
P2WXFDcf+PXjhIYKPadruCMMAEmI0GLAzgN02He4IIo55ZXWEx7rTaOc2OPnNGCH
++BuRHLT22M5+VrWULiY2caMO9L21wCjVS7kUNU0j4BhaFFAmKXkUQradeWTHqet
XQ3YvpZHA/PgW5UVtQBq/JRXU64wHHFtDrKxPDKquF61OtsHle4DllU8jTibue+k
ka6IsWthdMGM4QP8zF1CPXAhSJVN5ouVtWhiOrUnX8kUN/5O64oV5wy/r+ZRz/MV
hL7WMUSXc3iG6YN2fcZ2dhvvqPkiAJVTFokVZ/GYtsKUSky3ypQWBVMdyQmZEY7g
crSbvm4A2KqzcguSVB6Dfujl+fMoRtGEAG2PCbt6LqLTBCPfCtL5GgPQu3we7V1I
FP0hh3d5JRTmCs9YfePssXsi80rxsr6XHPaZz0zeuUddQC420cyX5Wa7g3ziNOkS
00+Oxo73BGhWyUsxf1NSXYqu7o9K15zG2g782L/gW2DdXCIiKr/jZqiKkyKIUdlq
RYya0yQbDLM+BLEZN6EdRAZFUF29ZGUYeWjqodYcp5ZOINhTpARGwYx2KNtSXrtD
bKsvM6XwhfFILfU+NOsIlSNJcpLtjEPUXLydyDyuP6tjvb3giNEXTPWvgjdN+Kxn
MwSqCM4pg3Pz/y7cK3XLqc6hgRHle/raurwLr8S08+mZfcs66TiM4YGB7Hqno2ug
dCsdC3t1goVu7mXTPnV2qvLxyrAIYEYB8gsfxS2F22UnJkbqMzx8P0QvHajUWoKF
7AHPpR/SX2Rf4EaQ4f+XXhxhzQ+rFxzGl8hqWYNcnrps8WloHBnNM2tHSDenxTbM
ZLvvEZ//kF4imGGS2u7Qsp/ZEGyNax+uwZa30Is4GCGhONLJ3gID6zFM64EN+E8C
bFgP7aoJu1j3IPzxUyF1Sl8ytNWp+YfJBxKQyL10bT/cmXbW1/PWLDWSKwFAi8oh
oowubwwGAAqYUULsodsrvrva1Be+fHP98MNaCfcvYPL1k2bYDkunZTDdEFYEZ8ND
oVMxgLFMKL9ThK2U/TJmg087wrjxLNOx3HvGxQVgwj9x8eCTOBkeYY06LpuBH/6n
ugRyxdTjl+EBX/yfkicD8BohqcLIemMwmER0UuTYwX7GGoY0b3oJB8dletmzjuoX
ABS7HjFzoF6QTow1hOSUfP6NEjENx+CiaCiPZdxBj2qNSx72OhRshwOgrpXRNAjd
PjfSeidrYS2lLo1xt/tZeRrs8Ai+4omf6kMFohusxb1/VfFjaU45dYyCwKodH298
A1429otcXPYJuiCil+BpQoVx95+tY/LyuyQgmEWXrNGF8nK254oy8iiW6nuW+5Bw
x54336pvKAe/cK6oKPn+uqsIHBOfLIhio7NDyomNZ9jjybN45VunvSi8XlDkxWqO
skLFTW9WfqUWF5Exz6I4XY0/wZM+USfj9OO3PGdlXeYZ6pgNpYNMWyAHYyqdh2SB
p3keXFLyswTA5FEZktT3Rjkb/RhNzbKQfQ2pyz20H+nCE3MAniFxsu6CS9mI1Z1e
GAplai7kZRpbRrOT8sSLbz6/Ze4kgG6WXcbiE5TClvgMypeDVnfLEbAG9I7rkUbk
jjyBnp87UgsprOG1gBTgZOZZxQnaMvVpkkGKTqe5QjTkiDznf+co+1MYFs2i++Zc
A79LevDoFvc5nDE+Ew4roPN7z5HtWrqW3YLHYUrAryqbph5uBgoOWzll0fyDFe5j
vQmKZiQvkvwFIX9KTa/C0eNPTBuhH/wBiCuJJsQAHdtI3xFF279enszsKWkc0Ru4
oPyu39AaL+aaxtDdut92+hzQ3XBqc0p7DojTbc4GVfLUB35OJY0Rk7zkcEXgh6Sg
Yj5XktXfyfiFtWaCUN1K+KRwWAhieDrH2HGvBPqjTKI3nOvlaO5vTaMqHkQbBhPd
RZzi3dLSaewZzGupzbtkX1UICPQYLrrKOHxTZfuM0AjV3cxlr3BcFF1Vj205J+TQ
1dLu2FlH5p6AxcEzDNg5LxVJ9FxDAmRzT87nrq8NgKRP8HPmiLpC0ESOQWTF2mZp
1VNLyUERMAVU2Dbw5TChz37RNEN/0tKxrKvPy/dxyUwOcS+KgymyWN1vwk1Z6mNQ
ggzxNfAKx2rA3omynniwZPjp0DmfOo+xttxJQzEhHhe/IcNV6rQQCI6r+H47ioyV
P+mmXveRaAQtT1/dj4C0OJNETj4ZimkbgY8cmqjgLXbt35YgJ8Uo4VvKdwB/Yymx
tUWPK9zrzwxHcOwG7pjJhITys0rRBgk94ma50pRXd6J6nJDwQS4dOTXMobAYyMVC
ol84m5Z+5m2IglbOa4HXQPmAlI51158Xlhyjy8HNyckjjcu59DtosxEtooy8EV0X
FNuNb0ptxrv4o369vWtoEwRawWreJ0rTBjXnLIpcMHPMjiaQLCY/8VsK4F9H0QT/
toZ1J9qjvLo0xAMdtoFzayKEWgkxhQg9aAFs5/6BArpWj8tbdS0zAU+YwewI8XY2
mQAdFsLabFwqMFIkSUfmhedf93ZjXPiP1XQmXY4csDvX2abVrVOEdG3w74t4/aGB
ZI1qE3kuxNxI2nUvXvtutoTGsVEhUMsHtJnFjo/3fikBu9YCf8Kg46C+grLMCTdi
Lr33Ogt9MIenaNfk/XgOtILa8wWltO0vZIlxjjFB8E4eKEcSn0F2Bit2RUMsgK/2
ekMgD2DNlg5TUbBGTQwRZt0HcYAUXIynP/A4GHeO5G4Oau4tIIlOmSba8P+qp9t5
MmmQozaE5KdBcatrzjRINQdas05IWTLbgE0/v9l8czanUFRqDqBHV8TrgrkL4aYp
fqQ17UHXslUO+90hXw8R3+VyGbsvSvUkzLGYQ4Oac+7TtF2T91byRfVCcx8wRuL6
V8VecjlbZNNDv9hbdX8Jtb/qOhEKHO+CdKyY8aqU5GfTkdCgZnxn/u9DaLY/3z9Y
fhxVNux5vM37kod6TxkPRN5M/N+7sKbEZTZb+fLurs5cIU+UdQEv6wWqqH2C7Svq
tVS3I/91GcwLVPnpuptTTuwMTEgSh7TY4jKCDYiC+8qEo9i7o3dxSzt7vO6zuspI
36bsXzcVO+2feLRNKKS/5DT+n8C9dCY5LaEmLYudoziA6XCGHYMZMI3dlMHtLEMM
5NPlO9LfQLT5+qpqKklU9XxwT0XbkSPguDmzxJMAV6RBITeRYIg/SYiO8+8OOI9R
uSKmzruMlFjywEvcLPfHasTzshRgvyOXcz8j6gEiHi6a4PKIjEllxSidahQvNTob
obZhRgRXUrsc9RhYqpBU3SLbZHZ6G1nf0KnEMEFrQIBa3ZDS8mCSIEwidD9FEmAO
kxG/8Qzo8SAp8cSFnJIlcdbDh518oS25iNbhKTVPuNUdEAUSU5qr5c+ioLZ9FEy/
e9dZpnfFslA5eCjvqvgpY0o1PC2P0c6EB30NzlkXF9pMv9QWJFbkqQXyJ7rrARwT
3hRAZCpLy+P/R9etkQqe0ZB0npDECi2U2FFL24PKZMgEcpYCUtgVTHkjLELy3rx4
EhjF/EWPllad/JM/fUEVIk4Ixpi5RO8XH0BEgmBy2ySYtAbtlERlIInSh4ou5Str
NO0dowsCyiQYz0FxdApxThLxB0E3+mLeLkTU6+xf+dzkPBpE07JJu2EyPj7vcKYy
UxrsC9U0UdBQr9DYA35gc0rP8Km9jf56X5SSprkFyAOEd01uR+Ez56FN/RrLpkYH
C4W05HjMix5g0kh35qk119d0ysFCX4eI6v5LrlWC8hxOkNmK4QhI0R3gREyxrrV7
yUQ5F8HnFqvpocHU0kYt5daz+NHWh/TTZ1Xnb8vRnVvy2T8JovlmlUzSVKYQnWw4
YqXmn3lvD68mHS9Bs2mvswzBSB5tCfG35/5lEr+jXIrgDF6pLD2tMMRXTXrIxFtF
yiTaMPthy5dqkqWvDsxOAnGwQdpl0C+3z1zXiANIfeOIF6HA/8qcG06CneQMyAGV
r8Qmj0mFyIaAC0Z5zDevT70w1POi5Pt5En9wSf9pzXL2rjhN2ZRuXoX5H2XNSxen
o2fp2kLWNbOgoX6+mpo7HCY78J1HW5qwM6PFrUwc/XGwJEwEydod4EqxUimxNsdc
Jx2W4GeUYDIxJThCKR5aGC6OcNA2CHjAiAD6ucZKMBTrSbYm10yZW8whIlcCS+3O
oqodp+R3FcZaKk6nuWnJhcpQeVk4ahzPbYgBh1TZ2S4K1U9ZqBRPo15seFkylMnN
JCjS6LRt7OKpFshHpv/GDgqcO7HURc3O9Shv3pJMRrxIxBwtixoanpfaoe0kWpNw
D0QvUumzvDC6PMlYbOJEro4WXgH9SOXhi71vrc+9+OCmichgafpXtTxQ/rh30Ps+
BQPi+ZVSaA5IOu74bCo8IWYrjz2kqcywR9pLI6IwyPltm+MhbwqOSm3wfK6xSrz/
sIwiqqwDOtGrS/HDZNi4iQx28cCb7wteu8y9LNOuogHQrDAUTZxCJd0VMLv6Wo+j
Mm67ahq/bY6gq1cTFbdiDp5T0SP3j5GVQ7CQq7jUY+1Vnq1AyyJ88z88mAOoJt06
LFQQlei3Dy3pTmBDs+KdZP36KjN/OHH6v2zdeTe1RmHsXdD5mr/lzT5n+T5bijJo
8zdTl5SHDsj4EfKVLKOD6cDiZE2X/qIFQK2F3Nw9VKUGfSa8tUs7ZRTo90CK/AoE
yNdCeaT+TzMLDtIdf/6fCHJPkWhZqzo6wej8r6wQTtp2xPuqirl25oQyJb64rkQD
/mHX7ICVEvFh0Ho5pJG4i2PSiQ6uey+hbGTcyfQ64abJoEEwSUFTk+5dkqf6qeZu
yq0ip8NfdYm6AblFdzyiB91/UXCxSg52nD1OyxR2k+Tp0MTXYGOl4KB29VyyFpB0
mJ2lUDRxPLmSFHxHpBB/GxKDPD5lHVs7lQ4E5Qffo+Y0SE+y3IbENrYx7w//Krff
mLqRXi59Jg9YwqXwTpKG/59cMrmPdYPrS7iQH/ospPxnjgNx9xiqpMyXliH+YKtc
fNPRA819AHM0l+QkgMKyezMgm2xZ0AT2eFqyxnwetoVMQfG6v6Je77hV2csLcw/s
FIQNX7In5JLQahcDiJoQO0j0bFVaPE62NWlXhYrTwcEl7z7DNCEissHRc9i5/wbN
Ph7Qjk1s/LAmuJt+Koe3dkIrgj6gpaFmvupQFldvd36FdZKB+St+gSRBq3R3+qMY
H0rFo7wqUN1oDLzyKnp2yu08cmCXn5/8goWGMGZp4piW1t/P/gG7MqJxGkECjAcC
e8lIQjDFTFmz6cTyaYeiZI/wlNNivM7fRFlYPVKXIRHHn5XHaGugT8lZOezYOSra
P2Oklk6rlPqIzR85fCdrFidd6Wh19I8AfHkOB2pri6n1t/70bfJoC20bXl4ty748
7D0WhFbXj5rQJNwKZrJrI3AWeFTFCXgAwBUK2P8cElPGQRPEsKRW1lv3JzV5mrL9
augPbwQjXvphyLJ71gCcW9Zo+6OzcKxtTJQNypZ3dP4o5UkP4cyMLTKEEEy0FUZG
zB989a6Gj3P2nUoLt0lttR9SSMHBwLpDFL8KuKqsSC6PuUljiqOALlHInwxRk1RF
gWR1Y82/okCerzBKzo/VxGBlHaVgsmzX8oh6m4JdkgydbkkxOs/3ZfGoK/Pg5aC2
LE/OhEM9Z0IUeNmg2AB9wkglBpTt1fcr/7NPf2A/5ACUEiWO7RdeBHJhZnSGCqed
nZ+fgAKb/zOlgxG6v6h5P74rUjSPmk2kVDpvQ765HBH16WrZKvtSV8KW0JHY4uMS
/jSpeaMuyhdei6cUKOFf+qgM7e0EqQ75qiymw1m7uwYMK1szWxxyB/pIXvi1pDcc
yLRdF741tqn/28x1q17wuYfVP3bpZI28avA9tqXwCL1pJc7QuMtMoflb84IQ8v4R
ji77nSXGBTUVAmPLptvzP7jnsiqPMaKRXNTFGDUsEiAJQjy4+TQOXHQwaSXCD3Vg
5pexiaXZNKRJXtbNCgnhdzGFg2rnqoRFzWnY2Ep3oyLlSUGpMMw/yhAdaSyQZJi4
EWGDTWPND0p78VJHzqHRZLn6RHGO+72oyfSGrFcxUDwWPry9nPy6O2UbROBlOGmp
Ax0tUeD8Zeyc0jhWrNC/HXiqj4SORuBoY4Ygs1MlrYczugkysnQGPYuOkcOyE1bQ
BTmDTqzHW7FNy29bGaFhrOylq76H7JA/Zi1rbnTYSAK14nkpCxBiSiLh0QYQs4hB
I6tX9LOrsOwbFO3y0qeNgm0NukjznhKdqM7JSpKKqiOnce7I1xijQVOel6JfcFcO
5qwxraib092Eo3A/SDybYvcfHMGbBHqB93E9znDOA0iSE/NX0TM4B4FXxJb+h6yj
WrbFrAii8GIBqb9lN3gkJ1KE8yDcMZTHCzSJYdsSN6l6OhqKNmv1oCKgg6u54CD+
z8m4GcHHJ2RRa+8ADqZYnHaq8++vLgPbM+Xm/9tiW12J12l+q9AE4PrUFGpzJ0lX
/muFvXXKBYI1mR24CQ3D2Ct/EEoftM0CzoZtEVtU0vBFycrgZIBmWrY2sR1OVnFD
ilk/+vWw3ZkCn1eQ8iUXGyz1C3UwuQy1XobzfkB1qbti78FX63kpmIk0E79V6a98
6EhWw52GAtaNsf8DEkuQt16f1jjp487X0WJW1RWXn5hvhZRoCf7KQULJ2G+nB7IW
VdQsZngiArUTL+YNNi93shvmjT+xFBwdj3oSgrcF1dbpYrZJ6DUFv5MrsuqrOJqi
yYsi09VkReVhP5875TQmqTor7LAq6XkYy4n3HgPR2YGMYxCP0XanFAE6Sp+vP65j
ki709VT2OKeBMohPTo9gcnqjcpKjd186w0sqiWV1/lvTNZ6Vm2eeNMQq03zOfiGO
POE/KEl79sXPHAWVq0XmlWBk06s5DEe4vsbBYNpeBo/S0FMuicWKzzk50VvE4rWG
8JCeoBTCmGWTy+WdeZeKvWJrVhlhMQW9lWl6DmxRqYObWIYMLS0vBZa5SqnXDloW
l/2WQWgvTKoKtBzm3VwAA3+sgNZTqJxL0xzi4HP1EaAdjSBCXZQ+LpeRzYSwCijP
v+MySUyjES4CLDEK8K+fvX8UezBM0OU7KeDUjwqx+5n135xxkes6QEhKHUcESPd2
IYP8io1iFMCLNFaI8LlMIcQV37cZhsctJoWGeqGm2ma7MkD6ZOi7ddu6nc+S+gCZ
KVXXk4Ab0ZcvZSZohIbl7Ils3rK4C2+7j+BZVMN2Tj8ZGfHOuUmAlPpbgV9wEFCM
JMDCAUnmgHQum5UOntyoDVxazXUedh/VwLv25n/0yqwxgwJomz/uK7NESdRX/854
Y0F4cA+AE3Dk1ydAcxbKLFzT08ctd5adP2QrrKXhST+xCHS1BeQCrTVIyI6QaeJp
i8uLzb/OX2w+nGaEPhKPxHc37mwYk/JzYLWF58QjjmbfJccXwjPtrAZAkaKKwt4T
UGUx7msxN8mqNNPKMCtt7Sag+r0fWsgCHzdssgImPr4GdHwASawcfH4PirGJiGRP
BOERbkw+nLbcJy9tfrmhzqss2eK3SDFyfDuKWQ7+PamQblrUD7UxOsvE/5YF2E7d
WtTr3Qk368PmdKMuU5QiBzl/3qkiMcMqSE4bkl2TUn6tWMLF01yHXZPhTS/Rn95k
9Iz9i0jwlfHLIps3RqUFWGULfe2D4HVdApvKCr1kxS3Jhss81fXhkTPGGmB8rajQ
nXbsRpVK8DL6zaLex41axKw2hjUJFI06JSH0SL7qeHl3t0fzBajs31AqlWUb5GxJ
cbd/Osuwvahy25B3ikMyn1Om17lE7gmHgmxTG9Bj1/q13aqUhVtHkePl+Ki/d2gv
cA0/3DLGSaDJDdhlm/MwEtKJdPiKZh2dMuw2lJVFbpAhgL1Yh5Od9znLhHF0tion
VmwShnwRa6FBjBX1jpudNELlphbaSXdlVcdlIA8rBxaufrgECBv8xm/dm4I0W7wb
3GN3JrwFOEQeWnd551x8Y43CQqsrMASYFL0rVt0nniJtyWZ26hAI1Wpy7U6HkJpw
iGol+OytxaZQACNpSQnNQZ0zzzO/ER1NfPkAXEuIEUOJLy8dzgemwZVzN3YeikdM
tCGTO2xOoAreecI5V3Oerqk4u0YLE9gM3Jj6GW3sxgj7Rg5knQMklBCB7bFe/ApP
kpnXvochQiaifXK7LTi8vH0Sz5FtI7tTwwOAsRk+zknAmEJlPF743Po/Hz40VlUN
Vol2C+CFhQFg8Gf+7ArtmaS5FY7bFu5cHi2RnYj4ed3+N58EIcQwqlbye/A9LbBM
RsXW3oF1MZc/rk8AHTh2Z9RwPs15E5WHRW+Q8oNMDDkvb6RW2G+vtM3IytfXZp+S
QB5GmPkww88qi2bj5luMSrGN9vA/fqzAbv/+x6wIM3LQ9F51jQpXcRpYKZH79ogX
S+ywUyJJxDqhdo2hcj1aKCG5LY+iYEIeRqXSpus6WrWKSzyDYsQOcnsXNJBIfH+t
oREmrrYSfTjjOo724ofeIzdoQKqSHC92NIxmm/p713wOY1EOvRdBNtTte2KtkLFl
G/LPQaB+JwZrOD2/aOU1rWrVMH3+GTyaS2f9h5xFg14tet3bmW9QvQebdkOE0sKH
cC2rFdo8tbYbwXkx6uorY4DJD3Igars3rSKTA8gE/8GBYSgZGoCJDF+glPF6HsG2
y48eRTNEVe/f+gMRY8N2mSFXdNbt2uyLQAkAZcaLiThJD9A7l/8j8KO0qu36FPTZ
TRnhUkOadm/Wm29YAfjmDbhZzY6s4SF4ZCZ9JpdkKLZbkKalK4Po7Ayd02FjrRE2
ZLahi072dG+o6LS9VvgLXkwfLEWnbQ0gTbZES0Wuz3WUENxCQcZyNEuyz8p7TxLG
RM+xWapqdnY1M07hWfbIEBHhmNmsqjOrehy4HYIY7vFoGPTQVv66NTi1gIiDktl/
7ueE4UM6lVjXax7GGtbdRJxeGuwGRRgeTLuSjCrBf+HtDlYWWUWEJRnpA4TQZkze
gshWdTOhsdotefFN7/UaGAziPOm5sMqZ7iLtWHs+uvJR3U1EtvjBOua9Mx/LcGjc
qp90ckSybZNOb2xDY11dVpvRtBnD2771h3to6SC+B3hOsUXG0Hu/75P2RlpXlFuX
qyzX8poH1SM+m5sYI7cFEGzY4ISWdFBW0DGHvupm8qnL9zlKkYewFnwz0SkePtLQ
j7Fc8wPuvwUf9oUzCPK4HYfNhOITzzjyf9yZqkMriAwWXubu3Yj1gkiQ+tmd3arr
Psi9WZpDy4yKBsrL9RcltjU8SXqoeqxmgrouu75E9C+26tY//WHRzYANgdloGmf4
DvAPHfP4ZIxqCNzjLnnrREotZ+fYQcwwy7jGFEWcD/TyVYHL0jKWFVYzWJSMdj5G
hDkZNNycPldiDFDjNC54AW74B2Wps3OmwBl3Jmio38hlRwnMKsX5iWtLBSCp/mFW
q2kNaJa9osRGTq0YxE3d/W0dOVTsw3F+QkZtqgngo//jJc2QO13hwofFG6FOcD2N
ji5NXiUAtTGLQ6aMipllwMbh+RIJ+ShAl9JzGerxSS7NuVn49Plq76uvTH7M/hkC
PUNRApy38tx9uPAhmrlrYLrD65Z36usPrnfVPwKXcmo0Yk4Z8KVTjzPNilT9Vgcu
ZfBC3WF9b70eUq1JCDXnJFZ3+FKyOmzPtCrhSqeL1mapwE8p3DQSaQ5SIGhR4mZl
JpgWaWQieeo5off1Bc/hIZe/+67wfXf9NGXJUKwiMoQ5+EdNC4FTJ7N/khObDrn2
3cPm5HndCQEAomrN1P3IQjyw4r/RC/USVYg+hF2EfMTLFRvcrX/Hh3bf4lZfDA+K
i2z7FSL+8lM7EbF46zSmWb4Ur0eiAtbKKPGkwJ+1sM8511HrmVbim4XICHMpGzx3
AgBlaDwEEpO1SESp33rR+GjUiAqMlTbrOsBDOrPurxirayJkMtqtiH0jNJ4GPGJ2
mkzg2uvpPT5o06oug5OqBc5F2YUglzl7bty8c5veyCbBWWgEMuP4Qq98hj9hhea5
v4bpbBVJEE+Rqbnr9LRak6R4H0NKBLcwU9RShaZFF1jBoJE2CZoG9dU9xychM2DG
kjxlhT+ZxCSO1MSc/FlG/Y8CVGzYROaIF8oIlXjm7SfdQtsEYzIDzvh8DjQHm3/a
NP3CVXuQ2melBjFtO8JxIsfC3Gg+nxoVl/Siiw265qPRrE+1vCjAcdv0DBNBOMvQ
ZRfN1CYgF+b7v4pIKlgjAhIREXGLvBiQnIs1mYelpnODfj4YPlJ7VDmB5C8bHek0
nh0JFthSeJQNDhqNwakuoUWx9E9apr2G4SnDTHKJB3mNMg50ZRBEfFOprjT1XWin
dOGvB5dE6fFz1E/AsS0QUErGZbg4zYn3R70h870ig0OuqLA9/zbQ/jnOqZC0J8Yr
sWxObP3XHjgMgiG/mnSlyeDl8cORNh+zEC7LRluQYjNnKDOCrM9JBNm5gPQB4e2B
FQbD5SMSrYmvLZCj8aIkVyXZSQohzlpoAnT/wPwVQUBMSV6lOPbQCPK8uvKytflG
vSgJM+0h4yBYw8xvVN0ClOdhUIJhy6dyuAOpouzcWaCF+kytmRMSuQiSXvER+vFO
9v1ByMKh+X7SkZDzYXljOWkP5zwY06QZ0/hNzlXAHeEzdyF/xuxWXZpIQ11HQ6Ee
BXgwtLHHjgtUWwEmLlFbQcN8TxsEm6VZQPkv30GyCb4hL0gyN1JVGo7UNMyaEDX5
VE7L+CJAs/GfJt300YyJyDpt570A3mUnGSIp/j37hQztcDlwAo9aodoKqtmsmOcN
GW/6MD9BOlRdh4n431Tr5J2ZkupLeBpI1BKaiaXJxUPooF8yLdp9wOVyeK88/jGg
uAvoU3vnFtzv+Qd7PyW+zvom8wKWvAsaosPs59zYzSD6sZ+cirUMG7rVsy6xK0Es
hFxs0zuOJlcEVzm/rd+nhALvaSgozmyba9fhYDdK0nJsGqp1o/sz/LYBCsTlSjsR
GPRCP/4kbuabMH3Jysjva5UoW87xCLJAlcCwhyo8bos44vSjMHIBe9hV4kK04bad
+M8OcYWiK1RpQAjZIEC4/3AKKBDQhNrgJxQnVy8guYpMQOthU2jPXXyji1XZVgJu
oN99cO68w5Yv8bfIjfPF4qR1Q7LaSgQHu+G2fBbBu6SRFeFN7/coqrg4nsiooq14
+1XG0PNsqdcSgtqHlQHalz15asmnXOnaE9SRuBJWJ4rR6ng4U0XiRCuBWdYIvQ0a
XcF+6o/mGJFqRf7Z/ZWlcck6I2/507UPpUdcQ7HHijtD6+s1WCDAWj+7Dcd6YlS8
tl/gai5Mpp96yqPJN6hvCcx7A+1Gtgt5yKLYcq9FbdsDUYxjV3DJ8k+slrvgiwNJ
yELChqnxvklAEewIUthgGzLhdoyLTHRoe5UZysYKmGotFytPqNtOJ8oshXgDb0e6
++ensRJhWu8tcw/XmaaTxTfpwwadR5vk293OZhMRsgv+BHcM5/JAWHNMm7wtK4ik
Ia2lmtAe25ynDQPRjYVJ5GTzCqSAow3ymGgTsC8Hm5H0XmWHxlKqUO3nEW8X6H0B
k9aD/jE4rCVJSH+9ppDqawevtdEvk4qyKJlMEPTXqlQcTuV9D23ZqZx+egKD6Nwx
3NOeszcyHMCzHyqoW99KsVYji6SRqr9e5BqSK5jDW6LY+gDPVkKb0l/4PEYeYdET
3DEB7CcEL2e0QxFlJXF2KX9Dou55dSzNCg+GKL3h7gaWpQ73H/lv8U3z1LpI+wpu
Mxc2JTn3M2UkK0j5Cs/vMARBXGgOkd6n9ZsoF/H1HcRK+6bn8rcnhDNoHdLT0Lm+
QFSu4hgnqEJ1xW7JqQwH3ZH384SISLW90b4+gF2TqvdpR/AjzWBYa0RW5Z6MK856
lLFdDZ3WXqMOjoDOQTlszR7CkNzZRxFCN5hM2wueFic/6oGjSq29O7bV9JhplEeG
woWQSKEub/T35aCDrOxB0XkGsw1XkQiBQHEHUU5+cf8wXPc+P77DfwSwZhRVOsfy
ftrV2su0L7mEu+Q3Zm0DQdj3ghrITVg+CMm3nSYvkLL9Cl+OLOg5FT6qTveO1sx8
yyyvoODAvMS9/+Afupk7a5fl9OPIi2T9Fwx1o6gIGXXw0D2Zv2APFedirdYmOYOA
j7bpFOtLXM/Av/1lDTXnpz2uc3bBNv40y5stAuDVggk8c6QlHbBSF3B0DXNmUTsN
qlyzjxfOc8SJ0G7/yn4HFdPAXIWCGEXHQlMvmIuut60Udz0GX3e39cbE/CxkZKeI
kx6Xuq63y4zZ5aeOjH4hh2yTYriiZu4W7ika0mvEnvJq6nUBNVc8BKnOQdMfXadq
UhERoh1vPk9TkCH5sIudGd9ESx63C65HnA1doUls9+psnP8hhWtOLW4HIMPgSuTV
ipClikv86FziZ78vnh5ij5oYvg3Ju/BCwy7s9J+VqIE4QIIukpjgg67IpCBDscCB
bxaCiF9bqw0OWmPZMcFuDVHNFQZGDDjsyAKsPSm8qMfKXk2OGHlToxTfeq3a1dpx
mgSdu4cpZ8RadTZowQRgZoqJjZ7Lf4rzkIfn8R7o0t6cC+vGu2GYi8uY2CWFR1xM
gPS70PNGTVzQBwW3Jf4WbrXnHLM26pcdtpGSVF41i+j3zARCZGoZcUOcWqg79h0m
h+pMtM3lmdLP+WcrB7cTtsvdTyJ6s9YmFpa5rnfVeZGfCjcIGjPDChllqlciZ+dr
5jURryUcAJkbPZ5lP1Dh+8nsA18fqsSznR2ycIir/SQw+M5bGxHMF22pzPgYyEc9
i0fgJzUJC1fwjbRSMRqVUCH1trjK+W/2Y+LM1X/fnwVlgSKNKspp2PjEt4fKRNvh
u+E/rnkhuFuNNxlMrSmhRfBeP0e6U7VR9C7hIMFb+NroWhkpIX0rv3Icsn3aR1GN
fmc7KPx1jJvqDyg2TGa/vKpa5jD+l8k1CLjhatMpTvZ4HA0gSrBltIMV+uQdgIRw
RVxz0ngHqfSFeQwymA+sH8sk0FkZn5X10njcEn/FiJ44on2YUIFOtTn4BqPjd5V9
+JbL2mW1LDzAtZzUTcFD38gkDN3l8eQJeiL8lHe1fnVzSh36SwP9b61l0sACF4x8
0an7Lk9TxRbB9lcvhWXaoEsaJeslc763A959w7E3YrK+tttcYTNFl0bvD26ZXM3u
DDvOMYgG3CDsyrYJ2WTvAfgwWLpXqPHsxs1d7WY5rzsGK7G9WcKmnZCWS+PLf91T
XMWB6Un8LAQbge34mnhNmVIAOzbVAkx/6b6p3Z6+b4+ZViBrWQLvlVnU5Ai/isZH
L9diVuDfy+4my10qFopZVBbybUkqpysTOhlrABiKPZNKGpkjaEW1iL7xLhsakORj
r1fc9hysIoqivnr1yo8xUDOLiX5WR/4ImEx53NgFSmMjGmPDWK7IoBftIdFp9g/Y
YBDwFLeo6/gTll1/NXDCQ/E1yUrqRVURx6unU3Aedw/zNMV3HEDbGj8ilNlMGyaR
LbZ+sqT+NUospEP8Gt4lHOQaFZ9bMHh9AfDhYTnKWHXmxvvRdvLyc00HTTEGAQxA
omkY1nwBOsnAMpCZzHYRGvJzoFHeAANB43J4W+rdiKNhLXQl6/wbUBEWmNztPmfb
Lr6a2LrDHlNNYFeORiMR4JRm8S2a3aK9SNxG2hofGrF/vX2dmnLYyGJx0NX+uwIU
NPeBAB8rlSkHQWi+Ti0j6fYKnus+z496nKQgMMTUuCcDpPUG0DWNnhP8nTM6wSSf
Yu9379QoMmeqCtqxphk+7+xruluPMQ8AKeX27bzpu97EYhz3fMjgrYG23LvLbHHv
IXQVgC73pkjJhnQQr+yEfjCzE9sxgVTtKDg7BDclq3LitvqsY4Owf4Fq6b9p2wY3
sw1MflXlz2CBfyPHDZnJ1F5TBNKJi0B8ztXzre+lXGK7+Td9aNrviSDzNy5JOGfo
G/7pv7hV1qJXGqQMHXRcA/ANQUOauS7wmE0qDhcD52EDsNhjkeqFZeSfwNQt71G+
wxcHHi1gvA3CWSv67fSWpLp3qKweUQICUm3O+Okl1O3gsCMsW4C+YQrjePJpCR9a
K5ISu+OQKmotgexVJlL1wK0g+kt/gq8Fdeot07SfHAmRFY16ShcMw6c2aEttJ20I
lwrEfX5ALAlGu1b8vPoXjGu+H2UbbeYuwG60mUCcXH/Xh2grJWCKxqAm4FfxwQrG
bqzThVn7bqbN6P1IWF5+s72z1eCeusguujZOW201fHp+IGOTrqUAihuf68nOWe2t
5Sn8taus+eF5L3VTj2nI8FHrVlCn7U3CV9PVMuB/do15mYx+dhzTjP7nPlHH9/Xa
4GFFENM24jMg+KoSqVORWVGl0JTqWNqZjuOHpGOQ4k1eP6ayaJCCFa7HqS53/st3
pa1WDVNz+LG8x49x9NMIx+KxuutqDueF117ywNbqjCptkgh6OQb/QXk9U33q5KY2
OCAnfk/HsIjIG6sE9xN6Rhwgmq/9iMHXoGO0PbjOVUua6j3o5g0ceHtf8hgVL0az
AcrdrnKANiCXAEKjSo502wTqRTpwwAwj++9HHYGNgoiDhWpBaefT43XWn9ZoA3i+
rhvqqOVhLDTRAOE068QzL6pPLUpfyQ9TbYwrn0omg+wMeDzx3Ni2QSy4IWhKU6Ka
9f5yIr36/882jzsAAfQQos/euvvRgN0sEdMilGFBcJvtvU/ttF3mH1rHSPFul/3r
q7OTm0DMcVCjNedt/6nafPcABcOV4PcHwij/FExAV1Ft1jvs1LTMI+UPm6D+RceC
rysp0D3QIjDCBU2v/PSUeA+SA3ZuQi7IV1ms7hH/E5hMCDaCx2TgAJOKaHT0vcta
jZCj0GokKX6887XLKHCTnRmpKERRXshQnO7VtqYSQLDHsKeu+jXGiIRjSP4AEF6y
SC1pZmPSyIEnSzLqCYTsVBXKNu2U+u85Nagt+I+DX/sJ7A+f2UhZYcDVqydG7u7j
9ewQbifmRqI/AZcWUHBqrNPWAPD1XyIeQMQFhlWHecG73dNGH6CmtZMFU396dKco
xjJ22r72tOa0TuINDK+I0pBTRHmYCJSGY1JK4R1QFrkrnmaltJp9fQ3FAuQOAwQC
RwOhfZlDaMlkHiyddJjzYs8lcKHGLd/zAHb5QhxxCxJzl8boCyvrJ108GG0DU7+B
wohSjb32WR5dE3AaOLuMnowZBgb9TygIDwoqwwEhbgaeJud2cx7Rg9fUBD7TOzOf
OlztiaFeefCZOKzdL6s0eIMTT/NFIpJhbGqfR7oKW/7J1rzkUCPdW2aaf45M2QYC
yCbbRTMtWGqRG8k0WcW1MeW9/DLH5p8sEamTv0wLSPX36acvTy98TqCeYvieiMpQ
SNKHGm4Nm1vrb5R/i2Nt/HEMOcF86tPc5wxn4hpnMIxI3+Pi0v8GJ7wdS3Zy0XAN
c6rNab1cnT52SUijgFYhBPCFHs7xWUX8ivwFXIz1GU8iW1oB0PPVtYacrzmXYvYw
kcjWuutvltKFbWpSo5I3K/Amuubm8X12uxxnjYRbDpAxtlnOLEWERmpxzw4HRXnY
BWiMKUPHZ19lMiFOX+t/JZLXdxduGaOIIYUjaoL3c+UHg7LaFe7VUmwCqNmONXqA
igH5jl3ScVNA92R6HZta8jWzlKtY2vm9SaycWkXTdFQVG+aribo2MfUjwdHTg1hx
f3iKMR7Q8Bnl8MIpxP/W96bgPPFtQyTC2fjRHmCVfZoeTvwcBk9j08GDKsrcS3ck
RjiTcNujogLohXtLiyPAoOhALHfhEJ8Jop1yXkLjQZZd4JzGJaccAWoyjIZKQ90Y
Wbe8eVoL7lOFqtKO80xTCUQ2E48IDaPGC9loi24ngQN8yEwi0cuKBsWLXbyDGIsf
ytTZi1cX4tjZ+IvtrTvRiUNZjD7ruL9UzFqOSssiiIkzgWJzuKOPQQrB/ALzQrBi
yzehiQ7pVQiKPLvny1X3Ufm3cmPqj1yzonQ9c4KdlL3PVfgUihoQx0KGNfQHtDJy
DBzXAuBymcvTcgZgRJ0nkwIWsXUNblllMDeHU/h6ekOkehCV7Cz+YKsJSvcn2BIr
suN/AjDs67m0uxVD9lGb38AwA8bwQrQvkhDX1mIKWfWXQqKSNikbm/nV+9x4XZg1
KBa0SD7ds4xFZ2AV69lXyaxABYyaWjHqJZQfSvGczaW/Q273tpOzwZHbf4On7LJb
ABgGBqiKodXdNvFxzsG11fe3+zsvMgYq01fWcZ9TBBogl3T8kAKHkABrFVc/q/bv
/pQ0tIkM9ufdOIjd7Lh5xCcwMGqeMHLsVVdlsKJhG6M6rs13wcyTF25bmjah9HpO
Uibz5aPda+qk1dt+BzLJI7oSCdWZboAWVnyCig2i0bVKJP+poXPMzxzFttNLIDYs
4DO3dEu4pBBpRGqoM4suY5lSxcj3O1rquwPkizDspu8p6JH1mVjd+TeMg05/kAqg
teAs3Uy081q0ACOrgbuGI+66xJDVzC2SfbgGEf9JFjSbE83tJwHTEUFr+99YhYj7
/3oEFMazzutBzq0TVluYlDA71iljczd5mlNiSYjrLqjP5DQAW+NZYVD9p8NNgfYn
S/nep5qa5/dVTSGQ4KCSRiRwT9KAPMcdKZwf32EEJ7YFecaTcU9WV46KmOBdRmn3
4D0GtLIj1Qb2ecloreW81SoZLKTLJdui/6p0Ma0ShtOgfh8uhwyFSmraEu5ou3kJ
Z36OgrFJ/iRTof18dor6gPbnEn5L1BqLGLMECZlBEOmpDYOAA26tOb2wJFj6641E
XRIYQBsY+QvDWJqP5UIp+LjGkTQwRECjKMpuYyw2roApXIUD3RNpLXjx3aLH97w1
d+q1otFRzsmdvu79Z+TFpDZb5mKfBqY+frWCE0fnWjZ6YPXPUhBVTxiHwqru1Can
ONkSCHtTGgHw5P1uAEwZYppb2e3elbGHJZVyTzjWtfcECEZeOtXqBIDGk4Vxhayg
tXQlyakWSEmyaTf9uGTgTxdTbmGbxbJ69eW1vfnj7GwS25c1Q2MRbIMz1EPmBQOc
GZ/sCONmb91yrYoQxgn2KD/oRL/KnPZR1AEBmICajV1QfIu1I8nZJvTa10odkxpg
DZK2lLsVbsq1YG0KOg+7Bwm6Y/zrNt0rnR166IVMpeAJxuhsBFkqe29Y6SrSNVW1
B+UYuLPmpf56q8fUGsVy9q2vi0Z+Z6eSh4iIyQTBGh7u2fMWLlXhnzLZ+gEwtZI4
vggwK5c3Av+pKbGotAKtDd8RycVRYHL4a61FzvVcBMKL4PpHC4dlLpEL6xvy31aw
Khsuki5UHLO7e1QxKJ3Bgz7s+q1krgnLvhzayUbjCnDEEZ0qivZjU69vy8xvA5lN
fqq3NpfNw6Tdlb5Angdk1PTwev6ys91oXKH/O64t51b9bju1WfavAkXz49/udSeU
6UxjwFCuNqrxTv2UUjGF33iA3qbg+/LkmZIs4lEyFruE/TNmgFhu6f1LKyxQijRo
Swjy/ibZX7S35LdjXJAiUhL8XNSCZdv2IsddgT1l11KrCYJuPlddmRPEcen/WauA
jRs/wv7sNa3RP6PwOfc+lJeeaR1e8qTkm+HUt9iXc1+Tphc0DgpZtYKH4NoksNKm
Dmz6icHT20WOQbvnNKrv7IYb/PLwGv0mmjpeHa74My+0lSj4BQLpN3fjdeHjMfg2
bze/dJvqETWKqKTMubgmHawYlRggnFzaKpHPwbjcvQMFM6gMs2Ie03fdx+B3Anlf
cRdTyc/38khV+4SMgGjnMJjHFTSkKdfnLAnhwy2SV6vSyy1Me3zW0++QmHPI0tKn
ow4R2n1yqpd5BSuuEvshFCvkPhum74yLnYYorLnu/8/xSkB2tic1xyPboItikjcR
QVP2sbw8zmhoh1wwOB5E/7wCeptuHlyspSTERicvz4mEl0WkuO3WXqDCpqiPt3Y+
as/cgnouXHtUDdWyz2oCfHA41Y4AZCpH6VrwDV9Ff4AlmTtiro8ysZX5EPyLXqp0
/6ljeiO5GYOi7fwl++J1dLv3lLrJ9YYC/QoLD/1UvPmi1cwUoOKW7G12GTotUcQc
wtewe096Gz/kq2uCYVXUotmCth5WeG8+mX3iCbonlbD7Osl8jLSfA/eKklw9sEtB
g3yyyr6imx7MPcwl56lofExpgu4CXnUKSrvc9UUIGcy7bR3PCzLBP+lJAn6c4nuu
Q4yQri4WRNtf1zHOMovrpIBT7ro8psp6ufxpn5S8cfKco6bUkC5FeREp+5+I3HOw
1R8AE8Y7jtUo+d7KR4asPa+46jK4DHmKvD/c816UiJUeby3Uv9y8QSosx9zzo4hJ
HsDoxjcpMN1tK8xQP4Hx+/z0HzjTwM5lr1PgWLL2IRTO3r+yYK/tytq8L3zdIpuR
6okHiiqIxywp8Vhq/3l7GMW0reeJkPnRJFmek+VaK2MeCCZMsvtJBurPf+QkAq7b
prifbLETtcUrFnCoP2EKe0CXUkTMqmF+IgOSbxeAenXL/NldnO20yZitjPcr1SZX
T+SubXV9wI64SrFQPSLPedJFVtwdNnX9IQPVq61m+P6J+NQvg6DOon7ziGUvKVnH
G2dG3/qFOCS8jb4F6n6HpVuhwyEVKMnL5oKInCjGb9qxuFR+OQOwVLPHwQyl1y4d
MaG8miVmJ73Rj+8hezqiHaDA3PPdQQsfTkEkpuWDC62N+cV5t4OvyfhzzfcV5u2x
RAbuq/r+RBQELZdqD6mR5rFWDZIiSu+lw+rKodUV/EwlEcTrQ7cayUsscTpFMFBf
pWPl3hrPmg22jKrI9mbejGRkQ6pnv1X5qiESWBMx9kwLORODpiMg5sFflpTkMZl2
bw8/THSCcoFJvh7Y2YtvJVA0IGeT0ERoh992yl3Qk5cHeEA2qm1UVOa/FQt/34mC
w7X599OiJ3euzhXvBJo0/rhZPL3bYvIODs0QfJh8IPYCa2YqJJ08CCKjmPQOJmNA
bE2Kbr+svFASEqloY4GRa0q4j0QEqf9bnbssX6j0ZRLO2o25SNgRb1NZ1MlNOpvc
j1f8njdObFT5KEz8JZ8G8LJNOoMdr1cW2DJUfv5g0/o9WxXnI8PTB6ZIhjRFPf4L
VRbTecu4vCSqzo/r/V2NgYPZ9E/318/Q8QtwhLn3xKRUVJ/h1ijN4jlBBSqyqeK4
oRXwTBC1fRPJDLYsikc4dPYK6B2VvShiWYOADBWlV5dwtzDSfXGeJqc/FgQVEn2s
tk+je2yoNtNolEprpi4s8wxcAXzHtNn2Ek5cgvlWukURhEWagoJOdpkZ5zV4GnvP
/D1PsrK9tcBiwFiBMvaT/kO6w+GaGvuUeWR2VXQYTD3qT894tHnC4xBY4l50CP1s
Ik+rDQvY9wrSpf2L1QTBtc1MWsz2K/1UaRKTFUXWUP5JXhcvzbGiynRJl7nLRdnH
zFYj66D12c7c3n1jewYfqLS11d7K8GPAoE++FAaiB0LDuIW7MfYTkq77tVHzldFR
JAwBC12nX9SXnLVXzE9SqggFvasm3ZixoGLcIwMRELekqwRoTbX5pgg8bz3siM7O
ca6vhyG0y391n3XTJbOyVPghED5ZZy+0LZCOqKxqE/83Mq9+1FPvkRv+0rL4MHA2
VwEGDceR0ZxQQbd3boLraFj4ZkOYHfg2YcniWb1VC5U5C2+LjsmzNdrYoVUfYsPe
p+383s2TzzWTeORx4Bmbr8JuDsAg7BLypi3ZwWb0VoBhPTfs3CiLJjvstHJHdE84
6DL8PapD+XmHApRhRkeOThVbs31XFfITT5Q9q1aKHjb06TCbrxE9o/b+KjdZ+cfL
3U9KUTI7PMWqeUvYdAxkzPQNv2bdRT4BqJU5hSP59R2W2OiuLIAOP6kPq7g2XvNY
z8vgUbnakiHpsH8RavZnp6nPAWdijAWsYZkjnAHZB6O2ZJFTjxdWpxh1DujVRLup
4MP8diHDRkdGBriUimAteojuKiVJ0mo4dufoHIue2W7EQ0HpfPJ2OBdptinRr8m+
23LqkuZKBzA5J4sS9sfBMNW8pfrFLXC3QUzT2BZivOTQ9qkeOO9/ihYII4HT5bKF
kgCtpzSFp4WCHdSdRu/y1c7bXtI9avkQdd+84CnByiDlGAJIKMwZujXNd+FlIucE
HqQQtaFmzp8rc19Lb4Dzcx3SlFk6aCmO9L5VufEIbkNaamHd8xQc+6a0XTEoquqq
z4OVmT8UBpuuVzKyAHbuP+8MH6v3A+PFk3gAGUM306rXcbggGXumx/uMgt6YWNCJ
iPCr7YJEiFDf+UUXdpOU5jYdMhlt0uFuyzmIzX7vFW2573am3tFmLsEkutn2luVT
qdd8fsDZsoGEPtLIzXDxqPMqNTw28y3ifg4KXGwhILjcmX6w6yq9i6pSAgp45i8/
mr6nMY/+Y1tleSwRaJS0ibCvrn7NgIq3EeznwWhQHstmE/4KE1cYf2oEBHLoICZn
zpe4e9UIq5BErS6pCXPf8XAEzaZ4rPvpUaAqH3BTV5Sio+fjbjVN+VVpZGlnzk4q
hw5EQkJPQdVJ9Kwd1t8F1QtPC1u0SXyX+jdhxTnSjZEQqyHmsrgzs6jb8ME+sQu7
BbJtoYc7e7y2tkBzno5Sr0huR7M6vap/1dwbBkbMjEdjGmtUecmMSvzvd2XSatFj
Ky3tZteXzMXmq+fdu89Gy4AjE2esa+R0OreUrFjKpFOo1huG92a1FMcwh5IZRiR8
qRkWRTLXJao1M+Cu8RCjQg/Juw4Un+blc9vDN1If+J1GFbK1qNOXNp20LyzQSitJ
LNpLCrqRFEjv16tKMR42selD+7Cf/ZRdlRRTYcvvID2MLxZ/ff942bhYfOE35AHN
0xzypiY6Iqxklc7RHVpk+uZoeajrpDoRdk+0aV26tNh9Gg2nAKkJBk6MBI1brKEH
A7cPyUhFyNOeAZMbSp9Yj36oXQbTelMokyN3IbunzKoM5TvHh3jN4aZUKHM+HwJe
WmE+v2VYAQ/8JH0gtjBdWmacdqIZxxp+14Tq0bziFWNDUe11Zp2/oEDaD+beFiC1
niGpt5gjrfJOGhf25eHoDXnLeNZYllClEpPlhXky17VKyGFYMJ4wd0134wXGQPDr
Eto92UOeHx0B1lATKNw+RWmxpDcUutRxn7CFHqtUfAHSQt958NWbTE8leFRqE+du
uVViVkUu5svrLuFOx99MK5FqSkH48TJXVSK7NVYzfaZA631rXdgVk3COeLlrj3vT
RJ0jmEYSUEWecLAY1Oeec6aWEBuMmO012uie1H9uLTMuV6DNCspyNparx6SaYQRi
OpxfAhVM0uVUp2NiLfdDk6mwM9Rn9LHrXFRQl+7h8VM4xORchHWD/xi2DahIVjeM
MrPbhz4EG2M3jPOg3cygkmWxDZIonwtKYa16w1KW4iHjHNnp9MVYDzOsJSHH7V1w
vq2GTJNp1fuA97N8iSZEPIp53O4X0nYMT5eyw5Ghq8ogxb7GGYb9UQZ4+qJyoeAk
knj6G1+Y6RyiTM+nMBaAY66JvxZfFqRm09qxJP23rSFyW0qd6ht+oT4UYc+baeqa
8bn+snKEkP3g1fpLXVuKlU1D4ruftIxigPqLclxeZnhQAlUTwg/2VqlOoVfQH0PT
NAExC5ffuvVIXCNTF54ccNchPVa5ueFLi2GNq39XPouA1yNwE3j2POAoz14LoQsY
faF+LyhUq6xGl00sWtv42H7DNYjkvZoTCuclTuIeKWXqm0meSZCiQGhCLYf8nvMO
g0k/6w8xo7o6BtJxPJmeOLcAoQhUUtxlVAYy1nMG7P1yvg08+dbKQCLgqaGoapqN
V3ggw/qLvVcnEEjbYfYwcE863btAP+8jvaNkjvVkIiyuXtRkLtlzGAYr/g87UO1g
jxqtcFUSKEO+Mj9bA3MyLwROE+BK/pM7ic8JBw/9zYK+S7o93cikClX56RlqPcp8
sweHqDXW99El0yk4LDF5CcJjyiu8joRyIcBa/RQIfLSBZvrM3gB3T7/XTIu310SB
MhPeSHq8ghLLfl4SYTn1m+C+wc/xG4wUqSj3P/KFXF7adF7EH+7mO5fYRnnTJNhR
sQRIoGy5PLBIqkcQ8QfEMdcXhyyeUp7/th7MO7thOIGQTirjSwYaQzMUayq4CltP
/Eg64TTprxJyCf44KI0ZIigCW9VEoiwkmu7PTjTDhWLsWMI5y0jGFLQUYh/5dug3
DtEAdEs0QugkBqMP4J7o2bHev0RnTPw21c++mZD1uIWvp/5TqDVnqntdvjh37puA
e8Vzov5YSKcEcaBB3m7tSMtERfKInHZlK0f6F9Siy77TcD2o/kD5L1aLMWmFs9Eo
JU3uD1Q5x34N/dZ7vUXNoXgScGQxBxicCnXePfEeiEch1xZnOLFcuNLWoJmH0I9a
Yhc6+rFV/F6FTE1vnTDIbejgxRx8Ns5+6dhicqb4QiWYY80bPfRHt+FFd1JupMQ/
cDOljJi5t56YHxWxYrSpImLBagvvDczZv18rPpwaX6+q0bg9mMFHpIn7uB9BMq3j
2/+uHH2MbR68PtgKmu5gQKUuVjI81rHIoDUOOFe6zHmXqOLAu7Awx25jA6SVIEnH
7AXGzjHwCIB83L+qezoHIvKJGubHinoFfbL8jB84LEFpbdi67oRIdJ2TooUmhYsV
hbtyGn3jBHWWCcqONlvXmer2/621fvdPO5MyuwM7kh6bO20T9crid3QLlG7mMlly
AtgOAFthI+hjOwkRjiD1eT7sdc9uiY6fjk+XOqjfcM28ULzzthuIaQKZ4EbyTq8M
POrNzgybtbYvRhtwur7yszqTItVHC6YmoWlar7pzonVI7tC3jCLP2NvutJIVCyuo
UOF8qhnVg5fh9NrBgNOWuyBafyMU5bAHFcaCKtVwHNiXtU0eXBoTMvwMP4ZJ+uxd
/XvGxTscTu/jAAE4yduu8+WBMeAZK4V7Ce2VITLkKBfkBhG+ypgOYXmMTYd1LTn8
mwAGPZWYQ6YdX3qRNEyYlLgISfMSSXpH0rRd/duZcJiDMB3tQNSFuP5KieuRfm5P
CiOhBERxYLmYAcD8aD8yL4DgLj3mu9bQyvwCduawq8hfQMZgmS/LEKMBsj2HFdNQ
z2z49cghy4COEH69yn9+Db9H4+u1IDNJpUtBQmDp3bpSP52Euv6TL9eyjzUM51gJ
rL3/5B5jiQJNtER8kgw9h+pg2NFU5E06D4zxUhvipru3hXKZJYSyPl6cZjgi8MhZ
NT8xg2QceMOVzqVYMowECRKHcfYVmLTMRtusof5+0qkiBlRWm9/k2WMVnIK751Ov
Qqo+ud+M7WpOQHFO/sl8Fo22lw0lKKW9AXJehVv2//AhelPAeqUShB3CrkxdGrHj
B+B0RBa9XpuA8MrkPwQdg8lGD+0CeXbM6KvDcBi1gEfZRCjc74kif9kEhOpX2FV5
dZxeLvxWbnmWpKZcff/2/WYUJ4AYnjKbUyfqoug/e2ah3fU98F/WMwTVY1eWBQ8G
KKFiWxvMGP86YWcfP1++Vp1lDJhlKAenaPRxDwr6bKnLb/yfT01hxSij+tVq7my2
9JvaVf8unyfUEZShWqhdFTCNwOFxJCCytNpJDM+BbblWSrxCBRSc9ZbVaTa/HOaX
A4DjfNirsnnevmhT+6z0LTsCmgwyOAnfQaU0aLFDyOkLzKWMGziuUAIH3dIfZe3A
dwlLNMSm5PJ5M59qi0/mk/HgliyNni2miNs4w4Ce3v6CH1eLQPZSCJXSrcwoA7SV
RJtvQ9UWJ+apRwiV/mfwemRYwDszLDCCYVjsxcmFNUblVzlPIq4RYsw+ljFmZevr
gbY9zw+4/PEgiWoUOxnbWqy1iFPuZA9ytiq+tdOw/2zKSGYz0iGZdDbhfX0OjbFA
UmpkkrY68oy4uArQzONlucZ5/DJpn7Ej2peepgZbSg7xj6GBtuyB3pG+daLu1gSn
PjCLg2oUpEQylovC8jCFY5+H6+7tVZentK/cr7I6bto9FOvX93/Xu+VAFYxyCjgg
SBvl3BFIRYpzzyNLnMuxh96URaCy8pW4ARGbm/z0EtuvQ2B85jasfy23SUofImuo
EKdkUfpc3y9pmlc1lpW3w4V76NIXXUMpwT02pum1RNll4V6gPVulThvB7uRsXRn6
q9+YpDYRFocTl5ajJVagIuoDyMgsgoL09n6gphZhENZ0Yyqp5GgbeLIjly+zHNab
obQGZlzCVZamnie/Z7GRK38O8M77scOuk/Pyi1E8UGp66a+e0pRaXBzmkPwxriCJ
Lu8zCCXzyoxObOctN8mud4YOcpGvPKl8teK8ImQ3hBKDEg2/g2TB9/Mp1WQlNmqt
hifVWInqJBhU+k12Z5tXA8n0LQoSgclAGOiKng8KyOYw6Oiv/aGqHn3SG1uDqgVn
7OAnP1g8/Z249ycriBT49XnBLlUvrSwYqqjvTSDkd4pO2sSHtZDM5Taa8nyi4WE3
tHF3iYkduzUzdGga0nF9gn4kIaPPwuJql45zvKNaRC5Ej4KEYqve2GLCijqMuz6E
i6SR38MCHodrR8cs51wInV1VSmD04lfkauu3Ozc4dvHseQJijAAUQKecISgNPDvu
7kmZmzlwO8gXNA/VQtR/fso+jcI28VnR5xPg5LAYAI2Q8cBihsiyeblWGfyDuDTa
UtwpMvGWOh73CsQ1i5o0tci+i4us2Hr7z8jyXGJ2FqTnNUKryw0NakSW4wPUXWw1
5PwYX5iBDgzTIMjzyN7OW+9MQ2rdP2dQlTh5b2pAMU8yfru+lSIHuqFsV98o22Q3
AkyliP4L6NjbNKzLh/w8q3FsJO1mcSake1c86CVWTgO/gCXqb3yH5z9p8518kvjv
5IZv3+u2VGnsoKaNubIp5fRYLf8CwGHhUxQuqEyw9Wc4bla3kpsTVlG/ZyOUpCpV
froOW3XGvV/KGNbDq+lRZrRDNzesypwHqmyqAA2A5pXh+W356ZOJ0J+qgXdJ1u+o
Aefu7JEDp1GgjQfeuD91HhNRqMfDlHnJObD2iIT1jlfoHJgrO3xKmhelmEJIh4kz
rbkGXwZAPfECYeaDA4AeWz2bLOZQoiNRLn5TwLNH07KfhjBFDzVoJsgms/jRCTsi
5nNDYODRTgvxP0MFNkQuldj2ObjGTW9uYIwOxJkatKa8UZtxiwS22n8eqLxYSZYc
X5ygqbjQu+op9U+9Yy6SF6d2wIR06CK2wPjsbIfjNpWDbjDz9aMyoDUAtYjFYIXM
mV/zdFJ783hZrx+45eUvXAaoiZrpevvDhglH5usHufoGvfsFedX+PCPiYeICFBlb
j0STOl1cN/ISstILotXZd6dpAzC+7/6R8kQgc06RK81tXj6WFhKDOCEcG6Gaepjs
vbsK/3OYg3GPyj5J81cD6C4aK0wNXrQ4hokc/SvO7DTrO4dUh1NplLmf61owF6ec
D7ur/SMBASwGD1v3sUbcN398dvhRMGQJupMStoPY+M6FPGjpX8uMntbPJZ1VhKsd
tDR3yJrIJ1EGVwsEy9NFAz/wW3ai8bLP7DAyhs1i8tzIxtkpN+aHX7OkQEFdX9uW
ZGeeAfqxkNFeMOU7/BpISaBFURZmSF7n4gs2k07exqNJHIyyulg6vNOqUzHyM8sW
WOTTjvoWinwp+ybXafGme44mlFR6sj674RnMBqM9Q0tu+Hhb984G+TT9LNkWKwi2
QANHoB8DIVx882ULSP9fuvkkqF/wRFZnHyDzjwoJeXnG5SPBpky5yBJD3DJzBa/Z
LUrz1kLhg/9aJ2V82rsIacrrzJ61CO5RN+eai0Hp36FqOz8d7+Zz++0sSPHP1cVw
Ct2qGRo9jTw0v051Oa7x7Gsn74DSElhgburjgjXYyF9ROQ+V4PcJeDDQWYAKYDob
H24uTj3TjNiJV+c0faH1poJgkZ8c+7zY0y8Xjn8edKAATbzsJIcSNEiqvflQ+PSA
xy0cotWxdiRT0wi2PaHucb21qE9ctuxOd5DvLUTedlOO1wGzzkbiTDwJFGOKJd8D
mvtDSZRCWph3ApsiIkrKLleD5ysBcEbkEImbJYf0K0EVR2Jkwd7yW8z/WHpFpc8m
YzhqBX6qp4b8ESVU/F4eQ8wrWYzNiLJ7SoUFSnyZg+0aalIkZUd2EpZ9SSGbmXOT
7uCCYvZYXrJq2dt79a7s7x/PmAPRCExNyJHlgQsAndx4HTr+S8Dlkf3PR9KND9Jn
pz8l6gJgNm7pnDGN7UNjXEu61Wn4ApLJWhe6j88+GziLTSKuGRG0bGDqIkJj5g5W
MZDk2byVp4v0g1SqVknREXrdUvTxdC5GRLwjZOGjQhFKd5TpfTxeYcXg3aOVsCZS
FSDAZhSTBCTGaw6qOm0kvE0oZ0kiV+wDzgBbNapXwS+e/pRe39oe5rcdFTeFgGa+
jDAW6z14XGpzwqeBytQWWRk34p1rAc2crOxhgVnOzg8RgAJHsfqHwgnhT4DfwrUV
NYq2DARpWccFsFaGswckESJNfv0X9A49/kCEdUKeV+hBHiLd4+l41PdW+IB4pwMz
US5VV700qSTVBiXVY5bbQW/NV7JywcnjRfSSAaSPRwDzxRFS9y+Axc0OgwkMzIj6
3CUL2Zv9eA6JryjzomO9kY6m4DroirNHYwlzwhLnZTp7QTF7EgVHvICdNunsWUoJ
kkXK+KJakEJyWbLacJrlXAsjJsil4jhQy7sL4zzXUNTILUY820C2rlJcawusmLRR
elk4zwlDjESxgMISN8bD0jBbVbeqeiIkaNzdt1cctz5P90KbJZUPREAsvKT9Q3Zz
AVUtvjqXkyYKxozTDyvTUqEkoVUwgePxnFmXrOjGH8pP3r4Hms5PymsZrB+vMjm0
ExnvVn+gUsWSKSHc18nqe1M4YlPtC2OyjbT6qp5cxUBtXBODvY6OfLoW/eqGJOzm
WuMoDQA6xBwA04Ur3UBw+yanu9ttMve8ELbsJROdRGcOpoVE7Qu0imjifq3rjA9/
TAXzuk/mUYMgeRyGA8aa1cacfC7iJ+l2wjO6RNLYJJE1ZuUM8+yzYUIP+w5Wruv+
sOizX8sgBURsE0PlqdFprCJWmqWVaSdr/xZ7uVgYeP72cth5b7SgBLl3O4EVsK4h
vELDafAdDDx7oO34C3MX19NLRzrrNDMLvCDfEQr4tYXKAZ9bAVCGI2k+Om66FgZT
aNpZjfomcsDVsEpoLdGmk9OQXZ2MxjyhL214qrnpTqczylWw2LXksEhgOSxCaNqV
4gVQJ12/ItV70+5FIjWa1DtjfwFqwwSpz2ljH+4DpbvV+sCd+qi1VADbm4f0vEsa
132pC+tYZ6lHjeINeJ29+yHu5ngUSx7XAWCiFq14WUr4VRnhDaJ/Xnr8lHJze+i3
jF69Zb4mzaFODhs3D10iscZgVXa9kfgN0xW6KyGjQiUFs6ODOnNsE+XEC71NKi6I
wkINgRJlOevS3xsoO0Kpx3CZbf+89MvNS+R6nX5jmg4oi/ihNJl1zQc2eezyZILL
/FaQBD7H0ziKYsspBv8TEzpZ4yzxM/yv+gxcXjHmnO2+uL/VfTBozaw3jCF6OqaR
WaqJeKmtAeulvlumXiHXtbAHE/qecLBw3bNib26ypUbmc3UhemZ3gzgfdb8/BMME
B85TDZdF3IofKmhidHCpM1M2ZJegmr/Ay3ZSfUtfuoOBw8lPTUvxRMD8STRtPvKa
vsvcYJQK6PRKpGjfv798RC0pITi2Tdl3xI9YQ+n9j1XBzTkChFvH5FlDc/BWt90g
2ogjIlnS+thC56eSQ9m7vFJXZWW7ySoBfnF1s14p6l3LFs+9CQDikUivgUmaj88F
YCcvTburb+w99Hk1ijTSVibOj6HE35cjpk0ZU86jd8WX/TuI9kGeZrkwdYgU+cb8
kJ5zg/T15zrQLPFyZyqaW5TPvI9cVRtOAVUr5UJre4i9VwRK+8yAplsVhtQC/VZ5
CaAEW7weMQw5+tKqfxtTbXcZeRUYgQQe4/kFMQ6lY4WBA/AJB4RoMZ8oDl9BSezR
BFv55LSJESkAYo5XMR1A7BuwMOPWFCCIaeIueD5qrwTnzqXxakj1NydLvFWlawhx
ZRTKWjHFK/4ssvg1FtnJ2ggrVVwDDnKXhhIeK1EOtCrc21YHoLuFG+YvrH2l/ClP
A7QVlJ8NCX3o/7HNQVT4pwpBDf0QvqoDpyeXEXbea4/XZI4qGy+rXJfQRCElePb4
0ON3TF2wxx+MeXlNbqgQcU85Mt00HPNWJxb8N89EAlT32yngmDOFibX/B1fv2dae
cAOK99qdtDSb2ePdXjyZm5D7YIC7Nw+VBRW8/C5mXMLb9MXWrQLbK6yb85H5FQIx
IPZ1FiiS3a7X7qdRoU6FhjK0aXehkyMBHbqdKX++coTEguyRMX2QjTAOlV92AGIz
qwBslzgit6AFkgax6yHxNO0OLibMS0st4Ckk2VFUGIcF6+/OfOMYSCf4z2GElj/6
aNIy6/MSzSAF0EoIDIhYpwzV+vtq5AWIeuZ4Bs3c1+NiW0DZKBG3CTzMhvu6d8k3
Lbx93lvtAaXnHnTanDACx6OWOxdi9H0CVNihN7ocJo07InuoTBs/VtIaQigujVCh
U37cvcdOmPPR8VRhq1AnQ3AIhvDRbt08RWbaib9H/HWOfKrL9tpNd8uxkbBMWhRx
OHqxZdYKClIaIZ/0hF4qpYy7t1vRas1XBqXYBvV8DqiWUAXb50D5GnGa+HVKdV2Z
Tfyz+rRj2NlXMInBgMMN/AglRYPXkarrneigFwwaotfCkuQ8m66ff7jBi7dueWad
m8yP0h/tq3RjHNeYhEGqjPgoSe62NqPfGJfyfQS1kRE6Kv2Em90WwzJm9kCOKYdH
FCpljTHJa7LL9B6kVp8p5ufgDx2GlTmuS6jQsiXNG2yAHTRSH207dI4Iuv0W71w0
pp4YhWn5S0XIr7u7raz8Yy5wK48FEr4GRD6Zjug8tFw48afEqu1wI+12hbS9E+pY
wBdx/TCXBlfOcXWdBxbSR+GOZBgIwExzl4lvSa5siQE/qLF4ggHlTAoqDhLx+F7w
KC+7HvPSjLsSZQO0XZXNDuPGGXX43AKzHmF2TS8i9AFU1j3WRxtnkpvbqwo05eat
ZKXlOjKuH7dXZQjV46LminEt41l/UybIGNtC9eBilgDgx2krePwThPIpx4uaoPt5
qOs3xjIoqia74dG50tASfESVPV2dN/M/LBETcCERlKFm3YqbQM3rGjcApnD1LUWL
J8TrFWeus+rUpf3zeoSF2uTfQe+dfyCxGzF8b1UKLXFIui06jdy350lyi4BiBTC7
MzeAEyoGXejgAp+Yxq4Iqja3uSUsqBfZJrUEL6USwL6nKk5gJMUkT7bw3yxNRsIl
n5mQdXdEwSddUyQDtddInUVl6LTzjdBKcAA/J92OExGnnj5QF9ECCuiIHgGGEMlb
xEvKKEZNfII8EXOuoZhWg+E9fICXvGCLmR8PACmcl825ep43+0bcxwze1dpbPbAp
kvpe95NosqWGFeEkiI4ZSbsUgFiKOcg5+loqPq7xndG4cKDDh86Poi+UurbJYD8z
MfSQzNB0UKHreQo8+ggrrZ3Yv0FUx+mWk2qe85cImqgJiETtMq3ZWiE66eNJ1P/0
+g3XfHzjTKMwWZfs5KuHFpu+umUg06U7hwPh9i0xyrP+g8vYZy+bx3mXM7YaGbah
K741Q1IbIZ99h2kpfJQDKydbCDb7n0ThwaWh85HgqCARyUiOoTh2qgQTCFNuPhaL
erDjzmctuuWMWlEYO22ks0NS5teiY1/Kg9vYbm6v1O9cz+AAAK0O9wo+UjLIxRvM
1/EJinohog4PJNbkSVH6NI7X/K3YO1lo/aiFdRc4ZVZdUvugRcOmMqIAHnSv9wKZ
mU1DyD/tQyp+ZqZFo9QPh8Lwq3p65rQxQG8dD+uf41snHjpFcA5G7AxzaOh851ng
fOIwTLqVfNggHkBESJt/eJBx4AhJFKFQJ1QX2hPtK2QDd9q5nrov//AR/aeLe+oX
5DrovacDyU8a8k7jWoUc5tOceki6p+2CT43lcjfrDD5bVOZTJcIXGOYreWBkw/HG
1Ww9kE2g+9vRXUsfnLjujj5CUo2FFKIgmQ9ZRyISoBrbOZeIRz/RBNimwIbI5Q73
lXRQUM2iydki5Ou6zEbLeSRBgw3qDJKODp+BRrzzKbgRJXuxP4GTcjj9HBFz8+xB
cQAvR2WJgkQFtjd8eBwDTJ/fMTcl+8VSguE/n7IjR7jXQ6SraS+oFkCLm9EYthde
kxj451H1DHnT36lj7MxLrjWhOC08a2ImbDCLem9w2hVFXtsXzfiRRjPohAgdHzm2
PZGHBcQmjKGsp/VhQHfSkyKWQSSZNvB+1nI92ziZquLpZ2NPZ3CiLZJyeKGSEGIw
evEfKJ2+cKgQ3MVZ4B82REG17gMXJfcnYmAmaIk0LZBXtRHzY0WYVPtF1QZAyrbz
s5/90gYfib/XxnBSNRNznwFsrZM3tEM3ZZqqWtmMHoYjloamijGyY3GG05zsSnVP
Ljy3kMgIoqQsdk6dAkmBzPXTRUw8b5iY6SEqp+sT1O0aY1f+xcf8rVaVjjjgNELn
6IVWh/OFfAQ4v+AwhXhp+jHF+DJ80i2ZlJ3Qt6dvd2sKoPydyZctp7r4Ne3gl7vl
rZhosi5OZKkovGVDrYpWD6ViVGg3NEzLaIah1l9fzIG6c6tMacj45xYURfPWihsA
1dXzFHlxT/lwilOmfWG28O1WEzehNExiGhgjmshjt/NHDyRGYA9EUdRRTfpcSO5b
rrVwpwsGCVEJAFAgIRd3NGsqtoqR+YvGS/3hpgX3S2B4gVOMrx+2aCkQ3KGHuhr4
CdKM7mN48hHrbrAjO7TMfGdryaomjwfLn5YQqPupqwE3MVD2equO1386sngZjNT9
uh5g91S7mBG3jp8T7YPFQUSZGs9hpTquWNKqYvPuTMv4/crgi1k5UrmUtDlxIcon
xblSi0zsbGCMyQ4ci00XtZwgI0Oz4Q5w8rRU2Q1G0oGfMH7F4yrk0lwRwJ1f2VR+
i7YhDPGO5mEQGni7DceDXjd+PC0ozRLoLCzBxrAVrXLQ8WyOzfkxyoX8HVl5uB+Z
8kQ5PQZPH867eLclNQyK4Wlp8R3dbFtXG6j355OYTtXTA3vQBiW5Vclkoddxl5gz
w3CGzVKRglrUKmuN9zv+dhvwdH98K/4+vuMeDvdbItPZfiVs+n976aQbRulxgRKr
/LTPJAxNVRwcHwpyEx/38OxDx4jrrJSyslUTQT72BnKr0K3kGLk92pKFQXfoN+QX
r5SaeilVXzPcQ7z/Pdb7sb/oGRR+e3wmKy2Ap2gLPnqPUKoOA6xbfpnSPlHl/7y0
MqX/H+vJxJzCRpj5URrf/WSU5NOu9JXgEqgXMj79u7BZQ//nVCgrsRcbVFfdi7Px
ymfJ++KCAbdRcxdXgeuIAezQZ+RJTPub1LcRAjLJXp6tkjlIIBaO8yAr1v5t8YwV
eKeORS/fZRDn2Mz4DgfVfvgiUdFqhTSKz+e5NwmMJmCnNqFzzobOOnZkXcTHukQW
798srAej0E2dOegDAr7c+H3sidzC90GSBGZqi+HNvwaJQntXpmRXpOxsmY3b7ECG
BagTN3Un3Rcs8rSLDZGy1Hj7aEdCnbNda0xOvy/LRNXEt08zsglEgskAqdOnHgBY
sjKUOfzU3AeXdTkh4lNd4qA7ltyfEK797Pj2EloNNtJYa2rDD5Kvr/bXi1FHWJMI
k67CJ7mxNLoGBrn/N2LQcNgQv2U5Mnk9WupC7bPVIhITPoYrxqMlUOURv9thN9N5
qf6R4jhqkqsGN4c2UgKfS1vZm0jRQlk1S9hGe8YdzXctEdf4PVCb+Fc+ar70lXdx
XZRbeZRK8N4/UemwThyqhdN2WWZfMutcF7k9aT2vUnnimbTMa8vJ9sCnwjM9WXlh
Doh4iaIT2eA1fg5zmO7BpyxrioYaruNPMKD198YeTbuwAks8K74z+JTj2wWm6IfH
FIKTvIjrHRHyXu2yw3WY1yOM/Jpyre8XERF84DZ5bDDKUumjck21uJjw0EiUKdqy
MbxPqm6KQvih+ChcXxi/V0bm47gteSAH5pgNwW49VPd4BFtpk8GXSeQJoZl93Jfk
j07E+C3TzHH9qEkvQcsL92GdMt9QnSJ81SA96l6SyDy5s2+c+ZiTRfPzQJTryQ8I
/UyoNGQ6MGipi/7Hn0EoZTTWULmBH942QIXms+SXGlbRqbDzWqCwI9dMkkU439nP
bByf7ipt5DlSvq/B55HxyofnGeXzqYmwnJ6nu6S8XJaHR6QDYzMEtoaCblm9nk2x
AcQmVVNBOjEQzP/YmGcu/kw5vrNWPLUcxYLJL0oSgnGk2HHcc+CMPR7sZ3oSIox3
9Gla9lo9eWJ2vgYRZvsI20Nz+STwsVDbJrbZLYP360mS//LXvTxW7FR6rr6MdT3l
IBSnSAtsqM00GghXbTD3GgzO7fkv2sF+floBtkePnJWh3WlWFh005FAstXFrFZi5
i2bB/d2uqzkp6aYbyBZWmVxAUX17lq9budssrb/Pwg1eC+0jxmduJ/obiCdq4AEg
TM4AXQhe5e6n2E+tI1ciFCXFWN5iB8xVN3w4tcmp4f3zY0/3s0K43az2MghtxgzP
quVKZy5yDtZ+XEUAUSNUvnSgvPEMhaug7BGbeIzFOPxRReM9Hq5mOq6eq+e5TbwE
GRIbXkxHGhJ1u2gBIwL1DlvKOSagaFiTJJHhqpRELR9syoPI5m6zmyVmRRNTLpHJ
c51foU6DR1hNXN8Axbw7idOO9QMMgvGe4y/VDh19m1ISsipgkxKUxvcWa0C3krSi
uLP3BgG80cnmNc6N/vZGK85LFxohFFXY13zPcwAxr2chk1l6LpXZqY37zrf3jjOD
CzQ10EYaNV9iMWIYFoLukTJHzRA1Lb6KbURkMLmfyHT7CZhUUJaGPSeaMOoZ+r6B
EQRNsA0I55mlykPnzCg4faW+JyhJDXOfUa/p8zo79rEGVjO+SkJ6+VO37QuBPvuH
/7KYlCEPYbr+hDYyhLbMs3FD2QGH8hqgcR/P09I6sqgYfQ+hFbVbb2/OahgB8GSG
Es96UBXzjVqbb0n4t1CRVSRfNB7jIx46nZr5FFlkf8yzwRV3WyriDWlpk7Gy5KkS
ddlc7ez8RclvTChJNAFG4Wm9sy06w7JoH4MFQCMwgy4SEfv0UboGoG6gpIOtCjxW
oRUgAkaJ0pTeYuWelH9OE9MHjdJHh0lAb4iH9wLprtvNA0gxuJTctEAYgLPn+7Ka
ingNBjP5/SjoYhqnl2B7xokHLTsFktzHnfIgzcQg5XgraWCqHN6sGNg00dBhGRby
GPKyIJ18wBPZIe6bDxR5fdJQBgtq3btwv12M9ITJ+c2wYVpbXiv6HUKwuHFLzDW8
ZNytd4sWzjFn74I/WmYUNLnr9UFMxDMVJR9zxNFBnMGv55UOoBaGL6LPvsAxOj8c
rbhXE4rQ6vZQMR4ltICKsEWZxf6BOq+wqZlMo5NhGxLgP9La7vQKkNseoOV+v24E
+YHGHAdfSpAUSFZQdL933JvAuZCDEknQIzwW849NM0BdKhCM/qFNb1eJxmWpjjGf
mfyhzb5iDLLGK+wAq+Upu/dTt8SsnuoW3CVYv7sF6NyvRzmufdJyoLAe3pdZSW6A
Uu15Hk/PwM1vTLJSgV4aoV4YzStrz2YA+/NklsR2VGuUx3VreAdw4nn/83TOov0O
BjLDk03k9Um+M8JYEwFbgU8Rnf+YtPYNezCrXXkl8oQQAzxXCaXF1UgPXlrpLqay
a6TDZHOHeXy0TDVD4LVW/+czwYYfFk20SNoZtB+Aq0s81TSIOnC4f0nF0AZUaZZc
NOuXoCjZT68aWJlJw1I4Z5Dkun9yu7CxrCcChzvn+Ohh41sUXXQz3HwMswq8UMMV
JwCFUCBuxAv3ywfx5OQDTFNzpVScVM7lC7Cxwkxu/r9JOTf1f7LcA+vwEyRBsGao
K+cqy3NkI4Xin8HJG0H1zOI9Q2EAO1ANpfHDDr1fEzdcXQ+pf0hXab6W7+lzUrYj
4fYvQBBF2DDPeXJcbqR7R5M0TCEhNfOkHbQ4ysjMjNgDqhZek/ZlkIJDXY+7qM2m
Vr6L6q0WoktVOWwconcnB888sgBy2YLQKE3YmvRaKUh1Ilwbkb23GpE3t2ejDpNO
aKTOZmyZzNZCzNjcWtMzw+aDYcfeIoLgLZVgh4nOWbejKpm7RDbElhTXTPh1Mj/i
5ag2OvrEigi4eTRIWl0Eyh1pP1xAmeV+pV0YJRCgYmL2Q2xsfwrRymM6SIKxTu1Y
IfxbIqnHoWfDP5B/R9tk9cXU6gHkf9BMYoY4pjJC5kSb1QS/vMuCTrvDuqtGEBf4
fP9TaMYXiSoOUsKzgGlDmnd4cnhLJgXskHC6KKsFInCCFvEyiFXODw2G7HUYmFXy
GfbTCA/fsRCVJndMquhytlJXx2rYB3W/uvz2OdMAnZ7m88/L3E0akWbHD0Hqe8S2
Tv8zXLrnmrzdOA7uroSN1XGLjf+lCG0EDVBVioBUD0MG2FpeK/R3vt40Mi5RjF3p
+w8kWyrisHDPaAtx+YcSJ0h1bBxuCdRsCKARzQJUCU8qdTItMOnhHsbTI1oyo36O
7NFo/hfU/SBG2nBjUZnKM7EA2WP/t+6+HUY7RAqwi+GocL7szZxMigQFZj7CZRDx
U1vKlil1YKaAyGf2dHHyyT/KocGRPgDnlj237TCyil3H9ydQaYRR88oWD9j/JLoL
43H9xjqB24qIpxeQ9FcVO+wfdXRf+BywQp9UVH96a7qvJgyTz3EByeVF3LwmjNY1
bSdQqBRwM2mvKMsIMlxt22aBFP5L/WZAAyhIO8nWp5ZDsCYSLIWANtEa1b2rc5S8
TZFHfl5XK4RpoD1AyVZjLn2XqfgJ3UNVH1Qy9KrZM5cWau4ttaeNv5SNlYYdTbNk
CPi/8704JY4Ikr14bP+F4KRSZV7xuxu9eY1LaLwybH6kPyknFI3+vwJT4gk6oO3w
qrZzfyD7mdC571/yO6nC4YzFhbYvW4lhxWhPI55GDjk8tPyeyH21iZsnIPZYUqRC
cGPLDBL6ZfV1CPRTJMl1W45irrssxAi5kczl+lyd1qKD6BT/TFgQOuGnfJ5J0noo
Tx7m5QEy26Anlr6NbQq3THSh/H7VQYFQcgoLNnrYckNbo2gPFXdwL3etmW9cZmnX
4L0DDdFnsCI8cSty4PT23tH9KpiEfgQKFPcoe5s2I4Iq624IJ2BQsHMTEB/h202k
dcKOlTrtjer6l5XrEq+C++HcO+nyhSbZPoYzGuoRdnMA0066mPL0G/ZiW5TyxVgJ
qOOVWhcwZqYDbSPY58b1VejO2qmF31yXQr2pPvo/dsfzpmOIpuq05+tL8vVxFwUZ
X9CrAzYUheN4rSSTfSEALjV7RPYqowm/d9FycJY45aSyJ01AAvhemQKDSltMN1ZA
DRX0/kZK1lHhkK41iKJbcWPfpBV1GP5gKv1t4nxCKiSlTEDRNqA2wTybsIP9pOIH
bJZ2Du136l2pP+9B1lT6QdERb0P07MrMlBcAohuKeOw/PeisC7m4WpPikD6+RYCh
gyEyCOKd6GKJFmRXoyABn+0bskACdm5TYqh5V3ItFAmnsr7Emee72tg22XZsfCKd
sPv6x1clz/CS7/+NgyJMWSttzqQfjQWPn37KivIbwO7UjHarUHmPeR2ecgbu6OzJ
BfIUtzCk6p/eLFFjtZvd0B/t9M99+8wVH6A5cavY5QLnWhLhf53g3+qO0IlnY5Po
H+NmC4L9jaQC4tXk9IGigdlWfPcJHFD7Ai94ytidYzIRl3MJJ08wZybmV2/YRCOj
uM7p7FU9vZj+jo4gj0ZrKyLT1YM2qeb2KCQV5Dus8NJ4nLJ+z4vUJoUgt1adPkM1
YnXAWzVkGozVHAbly3xPkplzYeXMOiDfQP390+W2f97PfGfdTm6LDpaViTHroqRN
1Dzs3wyM8OnCtPgQ4Qb5d6fdCm/HYZrDezjGhhiNetiS3o5oABNgfCOW1ooNoLKC
AIkMnoaiM2eOvJOt+Bpmj/NfHrJ/FT1QTe11RwExd+HkuaOBCQq4b81UVql0jWvC
+FCUphqyoYpulK2CrCZOhOX/8NXFOYxagySego631omTbCaAfq53fOHpRT8hza/m
usy8s1p/JFqK90dyaPlPwAjexTBY97kv5TkAonNr2KoLds3GrnfgCvn4weJGXJYS
hbdqDGq8Q9FDg5akwg2rlueNf5YA4xaiZVnAzby8mBhiinLr5m8Os6ZUaez1pd5S
KvcyHS3zoncxG02oDXzINtpJYRzIKuo/HRgg46MPctFuid/BSjbbG3hzhEEobfC3
yUhCsXNnTiyrrJCBfUdNZkkd0YxqujKmfXPSd7U9dOwgpDNcHtOVX7Fo7JXEHE2e
ZVxApqYoF0Fl2uEayboDXqbKnNpfIjq60937QxnMKTFvZT5Ip4a6THn5dwXXk37Q
M4JblROjfnCpDAvT33NOE1gsvqQ+hGVKr/xqr9CNzhj1IPcuILnlJeVVfp+Sltn7
aaZjo0u1fpOly+0aovbsXNM1pJi4m8H6gwJ0DlqaVcWTmV8bnHjOkZrzPqw56zvs
YPU3B6/+1yHHWCirHoF41wIdbzCRKFdm2s71e/pnv3pRcK0hsOuxWjtYX/PqButo
fQW4NYVOZHZGqtcAx74TWifst98tsPvHbhzoqAQkdrvFBTF1XFdjPIM4jx30AUaH
25WOh+A81vLQy74M4gf+mwgCV2YQhfkGmK78+CXNBNVNaCT0mIAZKbchQ7q2i1Ku
AnveDP/f93x2MIFhQpuRmERaMjyo1prp+QBuBe7n4e9YpNq2zZLlWbc4Q867NWm0
Uc0QUulFCGfaiMdS+eLfRWMgCACzcKLlBxBykcByZdY4pQjsUgENUlJJAIuk94mc
zcWACPJ/Wm2/w+8giw7diyXQXClT+Bz2afF74onWgn7VbiiQi2dYWe+W5uxkG/LN
0DoXur695At88r+RqEkTnb6P34Vebaqt+jL/EVMvh5PmMgAqb2/TNk3xKkDenGIM
9E7d+ueJwKVl9s8kqb8A/Ts2X/LGfZ/0jI1OBIlEnPK0T/BVDDqlMj3u/DZYW3Ou
9eGeNEBPIvI0WU101ltPBEqMPy9DXHqoktu8TDuQR5b3z7hoCk6RbiSyTOhtdMNB
calpSV63kr3IZ4fEb2kCNx0bacAWySBgYrrgMVf7H0LPk2Iw4V7YyipbFxVAhm0I
ERguw+5mG+50/VaL1/idVorC0q5ohKgd4MWlLiIu4ot5j+jNFDfOIZ7iVO6gNxIR
CEuoMP7su2qfotvN/dYvIPSLzCW8Ey4PNYUOt+zoZNV2mQncUNosPsrlMjxqpMsv
qmu7qhSzfN/7L47BSBmFUVGCBwxhmUhaIjwhQ6AeeAMiN1gmoChjANVNKpSnR71b
ovh3xFoP20wLudM6pJY6Mc1YG8CdD2bTAuBOjObqqpsJK21EH7WLDmet2eGYm/R7
1Q+n2lv8MSIfTYtdriDJ/70cnJML6GLggzz4KBLcMQ16aRATOiN5TuBITJKAkUiX
s52ptacyrT5swfFnB8Sb5oqNeZysyF30nuQfiu3OgBePsFvplXPXLcvOb90QCiRV
kLKWt7wxthiJWUm4qTZ9EEa4UJ4jqXKxHiTVNAvF1IVPPZ9mdFUT+Y8ftXDRPwmC
SgSw2vHKcKbUIG3472pKIyXor5A938+Yl3Uy9cG8JwhSePom9tBrdoT+uMwBNJfo
r2WODoylVN63kk/mFqEWNI0ZXwA+Ox2IJ+vMxrji7r20l6RDzyclv/mVcCYzuvDd
nIHVQ6kziak4KiBWkPVcQeOVSxwqkG7COGzpov6MPPwGr9mzIoQgR0nSMzFj010s
EpXsoVJbEVv4mUPWnzJWrHDaKRSWh4cKfax+Cvz1hx01BSkjIDr4F896uZSzWBy0
bHXtxD9YTGml3Um8RCzdcHbaYV7EUlIYaoUwCY8oGh/ajuivbR842AxZUv4XeXGQ
hP2E/7GTsRJolblyLnweOdW4Sr+4Zt4IWneAoOW7V0YVh8W1WbfNWiRzmg2nm1Xe
pollbdzFqH7BxnEh5pUUD0ORpkGGAJyAk4cCRhIw96eu2ve5NcpQOiRpiSwDzqhp
HmQznN7Fong/DtX3gwey4fJahsao7sEdj35L02vu04sDpjQfN/OXu9RowMATuT4r
xgMKInzucM+AD2RYoUUJ1YoxknywOudCtNujWl8F50wdCiYhCKYosEG1CDD5/M32
X2XXdQyxHO0Les1mMF4kWABSAwU7WOcz+D3PhFSi1Q+hnc6w5boG8jFDGBe9gSpa
JW8pYVdBCRpKSEbe8fe2M5kIqK6snZql8P2J/nCVqUisKkLVISXhKvFdsfL8QpsD
Qn8gq3mqmrAZK9Vf+1WuRjdFO0HbAucsqsup8eoaBuob6kAHcFJlQYZnPQ83PF3w
8HRymuTjGzhEu/xMwUL2PgdNKhIHlZBCHy/xAlxIxpX9Axi4xGvm+7+g7xb5oABc
bieV9GsR/hMxzUhmTl5ZI4Y2shZz2ZIA8BsK536b0IDF5jQ7PBBDimq2uTL7vS3B
4dH+5WvNe3s5z+qtP2UtAKG6TKMBm871bVzeLfj/A+tg15m2BK0R5cYEZFbH4R4P
Zl2VBq0YdGU7V5iGCjbKLi/bBiq1pT9EyetC9lMxnch17C7V6QH5w9gT42XmElo3
R11VP3bNZW45zv2bIVP8vGE5yQXgAqqFqIgAiFS4kxwaRX4fjDUaNA4TxcNnjwzi
QUUMHAnqLxlRr1b83nlzCyMlSwt0WnzbqKwz4WHK7ZihIIatnZKCyl/wzYhM7xsW
74dqvnMbPgn77oFm+VhOlfglCADhW1Zym2feGBpWPooksY02LcvuenFhKl6aTzqP
D8zyEYSVtZGfV3YEo5w7Jl85xPHiC7QRNRWLCOzIaQ02PdOeOpi5Zfd4ce0LKK2T
oMb/ij9WbSyb8e9GnRoj6hskwBLP/8lQZ7kxq/dMfg/1+cVfhl87y2zmAKCZfhWp
7nm355fLhQpnkHsYV0pI6dAniKMRJmT8ImC7Ea5PbwXrUWmw1DwifbpVV0b4ZHeY
k3Et3Ol2njSdS7f1+gRmAK9zXxGWKy/NE23E9qISdRzQQgv1ZPmYn0Ga1AYttGBV
SJXSVrCySjxf8+WB37uy82lrvUs4IvXiW1V8Rq3pgdvVSadSqBAn1yArKnlvpvDW
UukkM9WftZFlEPnX+0RVsngPso2stF5AWAJMVdAj3Irk8oTDNrscaOtvPt9hbwMz
KjKEqZJqe78ivs0BpbAJJtypbYr5HXbeJdCHjuWBwP6vPfqVqY/twlC1f354D7uE
c3Kv2j4RUrV+COjxZcDVopvRhzTDIgM09Y6YmEZCHHtVYEtz5x4o6CX6xa02Brbd
a4ALQK/3AgOTNOv3WJctoprGuS1UzwonYMLdZuv9j3sM3VoOVYkmJtRsyOusRZYO
diw9QWNISSnmHktee1I8GtqfI/22qJ3tixJC2OJJ55QZCPgp0iPNCvbswKHUy/VG
a7JayrEC2cL526HAKDYJwgSofLwuXPkPegtqNYplcYER9q6XL8pMjXiwa+jzM8yo
xpGKwIHuJoXe60WnaOVsxAfb8pswBCaOnRybRKlSPm/61lHU0OTOUSHJ2LfPh6CN
y16BoJgQ/nb+YBPZApfOaJFLqvrTnHBha+F4Lm7UaatupZ/hrtmR8WunD4pQcRsI
jWTXuLwLnEjByBoCOI+pYihMG9WzNAhjKWP+l+abLKGzhnL9bFiGfaB/wt/7NtZH
qEEMiCp+Kai9qEm+JL871FMu0ck2+x+XvF1boYwttJBCYa/RgeEm8niUodof/5Vl
Ko5diJXWWac3HbJNzOBKNSO/Sez1fY9TKvN1nzB5aLnc2j1x2VbxqF/F63/fbp8c
nFesSX50FXK+eEPjYjiOi2hHXWiUAnCwZUc0rjDkvmYgjuvg9UA1TyFUXNpiEoar
Yu/E62aP522lRFcPLhV3JYvt423WJvmnvlhZQ9o+GybTDLhnFvU9A7ob9nh+0+eW
SHzR++YbZ1rvIqXpqYQbKQ/IUfHwKWWfXsf6iMHdLJZ+SpetcxgXJ64Ktz8I4YKu
TNVhLFvqrXcIGdBAnD2vVmLpr7N/SAflV+Y5RZ8jYa4JkDLFBGnbWOpZ4ynQs5qR
QnBXMD5QTcfliya4AT0lk77m1sO8UqXw7R79kEqD5plYqJ3XLJ+1Z9jCXK1MdQ1D
oG6A3mG3Ar7H3q3bu4UU3r6zeLVy0D5BLjb3kkYwHasPGIOACkRH+wbNXn2kXRQJ
0Tv13f/BkYNJ83pwT47zegBuIA4sbuA1QQzOXPPGfKNv8sJevlOgOvPaIacGBfas
p4MgYKQqGOC8pQEn5gjCHBEua6KMI9nkJefSHRQ4QUly9mSUOp/u49zediqRm45K
RKP7xwS1cXapJlXB19ucHC0Fcorb9PBBHjSWTUM65tNrb8P6BlJlJ8Ae/WJsejum
Uoa3+CM4iPrvcaQbXfCphkqj3atNuWVAbb/SPtXLLlVpEljhQBgVWTvHoBYB5zES
FkhicL9BNIWC+Y/66WEzKnHjzsrDJKtRgpMizzxmX9znsiGD+4ijsQrD623W6h7h
1zFCpxQxle77Ic1JfM6fAJw1vFFlNjcvTCH4JNJt8XRUqw2vYx6rdUag0+Ht8qc4
ZvyAce7y4cav9HRnLPF7HRqeDh9dZ9M15HBn9TDKy2CI65gv5GGjRfYvbT2L64nY
/ZVr9HoHbiJLtzIdrVbPG50YF1DyhI22y5Rm2zaROvarzCV05WHbfC//9JrFiuti
Jo0cY7CO3MS2Vwqk4+Qzwtcrx7i3x78H04qiPvZZocnEdj6PFn400QtYXgKhGE81
PEK66+DcWMWeK1ApmoCmTIdSFFINrw41Lykj4FoxXR7lKEFNnf8FspiDLN3VkA2O
IZJMD+pCj0Gw47TU5fEqxIiWJ5xwG5yMAhJP+clWbX6DLCnz23nL0dm/te7l3PYF
YMTFiNjLDeoclJic3JkxR625bmKePikwPpRH7gPcUUTVjk3kc2FyYSheZRPdK7uy
n+IVWS1aGLlyWtmyjQSHu5FMQ5Uk1duSO04uYEJkT6GS7ywGwGuCQpHr7nUNc2bP
vXwXGwkvKsz686eBPIEKYULa7YmYlUGBuLLUhs1J3rDXMOer+Vf40YhuvSGtmeVi
1aicNtQJDF/4t64NZ0UKVwl/UT64zu3fO9+IKva1rhjZfGsqzZGh+FI9/EVG1qTX
D7eHHCZWC0Prxqbe4OKIzy3MvREP0vaQgdwkI7Oh6cbaphk2gHC5GR2boXol77ui
qRtc/CK1shY/0gMU1AYwY4ajKNgueC0+Bk59vNdJA1u4IaBnNlOCN42Sjib8Y5A0
QX4AXfo7HgLOqJ/nKOlydSBtML0OOPkxIECAk+du9wlT3BwBMTS5QQHm5B3vGaVK
8LO9ydoININlkd2MA1FVesCtxM0KQtc0Qvejt3kCU374w+75axvfoX8eMrv9MBWq
FCnl9JqFiJl/p9TfqE5uwvs6Hk8z3jS3sz+xnpueBngO2XO2HaxzWSgY01fi1ADj
i3Jk81uSLVeUOklbrQEW4ABDPJhGi1A+q8G0Kv2tEXMS10M3j/lbeqxiJDmlV0lY
OZ0fco2S/t1hC3YMO7Z7qqb79Nnx07HKiQ5kvCBmurv5efaxKcNi2TfDde+bI5af
yvPEIE6Qp76DhuYzW1n3gGCL+LdBVK0UeaVD0xKJPRTRheZj4sLFAZh7L0j0AM6+
3YpYDTkaUPbnasMTwMpxzXGgclN+Gh0QM4CQ7N4sFbf1EDAYTcKsQUqs2MIpekiu
HSsAbLLcpgfoCdwlEQRzrOH7BCGQcB+/N+i9n9rGhV9OtUwoYKW/OfFbXOwq+m5m
UQ09WbzzFJLhNkqmmmuJv0Fa1RczYaZr50dNoCZybot7sT2YP+mNCaQA+Nr1dGsv
5zAjQYE8AqBt/NheV9+Xx79htNIAR/BmzXFRXSjlGIncNlJ2rGDYNbjETKr+dcSQ
OY8BBdhOqL+DdHJ7417TgYmojw/DVts0OM1hW4PSJdmrGSErVvQsAd3T0H1IooIY
vaP7jPxZnB0+0MHkKQrklvJJ9EmFoe2hRr3rrIuu5MmWlmJBwRNmYhpOywd/oj8l
mbVVyuDiVjDlDvpSRlDqU7NjUqPhE8ZM3jvWrFhTUoaS051xNIyGTcAeBdIpyYG9
ss7HrqUwIyQt5hCqhASN2wsfy/ZfVvNbLaoTIO4SVge+UGkTkeKrxdYyBof0SEtZ
pV+mBk/np9dYjii9yp2zSy6irJuI9jqCrkvH9Q8JLI+BYvw0S7MEXc/LfzTOamTt
x0ufOUEbdNLivFn+T5FIVuzp3vBZjS78ShZxM6uKUfzFLy/3akVa8VJPh0e7bwfj
kYlpxmAzRrmR6d0o97oLO3EDw9mNhY0kyNN3+P5QgDgZs09TQ0FdG2Imw8m/LM/T
GzyVBOhpenGghKl4yGmlAtD5CCk0NEi0m3mz6qAL7HGS8KDVSiiaMrx1KHYDmwVg
/V+ynclaPK1k3dApt/Hisz084AU+0D1umrBuaiX0apj9SBMUL0AYnqDS4Nf1yQWX
bsAV3auBDmsRs5gQ3fhRSnYCdw2OKWXTjHvWZILY+hcMQowd6YV49BViBYXAvrWh
/T/U3XpLvAI9HfZ2P4a5AqPSm0+OubyqlS2RB3C9+XgvhqOjwMxeUUNcP4AZLEt0
NZ2KjYYem7OcgG+KRZVgaoJn7HT87tS2ei0HmcQZixnKx7fysMi8ZddH/nKxM/Db
cntrMx3rX9D34HnhuuMvSRXXWoRuH0t8qn0n1ez9SQT0iDCXeblPvXlRDius1IyG
tMUl04c3ipmkaMRjHeljjLXFjjrZI2wo3UJR601d05554HwQR2P8cbZZxIOThQvJ
PIqi3ZItMx68RyVN8hJpaLS3M1aRWZRYwJ9/ktD8E1HTEdo8zSjQUduu3RSQUIC2
EdI6sHJyljFh08nfRZL+OgZP0U/PpdVsMQwPLhtuor4YzNfsE3sDs7wUtBcgzpnu
AH+o16ICQHO71PJ0kTk7NRDZSU6ts4gKCIznITCPV81Ki/Rb8bn2D1pQgqvVc3Nv
+F9WAt+ykcvo7hklX5iAuQ2VADZrM1fdDeAt6Q+P2BqDthfwH+oK5Wz/+9u6PWhX
3G8Q2Ws6p1//m2ExOYeo82HciG+PCHkhYzYsdavx1G0st6DWY/r+WhS10/2GLiiR
NgnlIXfyW3BXTSSGmVyo3vCuPIaJEUmcbC+TrLeKaR1DLK0ATJOJWtw/bf9EiFnR
5ZkhXma5UAMIY+CPFs+GE92a1k/eVQIOAChdluhvoxZQIpV8S9mQIZajF7MOW9Vj
ebIo6lB8ZPCMujT+BUB3qXeizh3Bcvn5kXs4FcPE8Nz7PinCk/mtLQURpgXNvZSp
8586QJqVKa/4Wvu6u+6bRYVRqGZp9pkz2CMZn93iIhHx0cOUuPtpPes/ZdUVDd9r
h/+Hb8Y40i43atouLDnGyTe5krhRxsa3jugDTkunTOADOAeXmFEOGZ81CWK5q6qy
NBO/CzYJvqIm/n4M2+66v/QR1r6Z8BF73/tKL2810hcLgPgsfebZgU+8AMjXb5wP
m0EMOEZJOe6HWJeqnVRzlxiSf4Zc1xeOxRe0SwBZnRAMoLCt2Uq+shRfuZIRkBt0
cr84v18EkAgFZ9xGCeOOCrZGmv1yiHH2yT+4MgqrE+jsWxvDcg8m22t1PgSuducZ
eOy6WmhjenWWf80FK8QHwfOZ5D594QmJKQgI1d4QsW+XZaOKD0BkdJp9Y+l+wKCb
L35twrC/b2C54/OrIVJWnGxEI5qH5hGt6eFzub80Cp6zQm3B51yvmcbowrAee58X
0eIXp/Ny3jFXR/92JM/Gy1lZxTOmRx9ynW0+OzFrGOgHxlnXjXXp8tnFQJzZFjbe
1blTyJjv8C01XoiEvNOAjDH4ORKdvrtD0bqRvt8B3uCBOwosNAaNv5Gxbr4wZurI
02TK7Jp9FxgkqpaE/9T2Ku66hecN5v3oBJSqdrJuh50n4b6Si9Flb4KJTNt3jcec
45u0Olntz/bvTkcisdpxzcNqllHD5HfDWZICQbqsi6pny+QNZ87u5eihafsQj/+a
tUZx5bXBU1k+QSsq1e7CbL5UgF6wI/+OolsvKSCyCB6op8jD5cmrUD0/cfYK5Ui9
SDw7UVH99irPwfMJaqLV7H5FltEEWNNHqQN9LwbIRoDhwrjlFiUuqHhzhqr75SZi
WyrqVcuE0FgzjBIeTY+4AQoiC+rTM+lYa0/2mSW8pv9eQtTGuz+qA1GQ0F4hPjNa
Irw2c9+YybUKqiHj258cbSzIkSquZq6LGaEE/Df5nlegOdADUXSRqmvICtGxgf4f
MA4sJGkglMF+LTUHztp10x+aqz8y7q5EukBtkJgR5k8yCVS+Uen4pPAe4V8F4jsm
r7oegVOg/ody8sc0+bv0wKFDCqWP3yO2S6UMLjGlOQUk+ShKaEAdF5rA8I0N/MU8
CYnCAcHHrsbSKTRmipx51GLBHpIG8MAuo7ig3hts80OU5M5npfB2L2fEASAhMw/S
QLibtFw9ZjaLymfwtIcvQ5q7SRTlJrNpMgj4avXUIEa4foBdye9lhhnAAHd1iwpz
BSe9/4BmNQWew0Zu8ecloinGj0LwmSEJsXxL5oWREiwoQEH+H15JAYyyRDEheiVm
u2FyzsZFY0p8c1Xnvk+Sty0iqPMHAIh2tQHonin7uP4Gf4ndwoH/iCjHqLtSuepE
lYzKnXRJTv2coM5XHJju7SzKUGuh4GkQjv6xjNEIwcsxYD3RXZWi9t/+GPV1gFzn
+0Pt3nzvyVsFQ/ga5dTkJ3zXDwptQW6oaNzfSuHsJzpaGD3u9imj7lfhlRzuDAoM
GcAjJS53hHLsvk100d1DwVLEyF6VoFTVGKOsf2DfU8UopP8suPSqR7wcIVGgA9MA
QTFcYZj67aJRdbElHThnGIKG+7SMUEPK+Kuc9v4Wnnop14BU1doB1PBj02NtwJEM
9HKmiPDx2E/oslZkdt3/qMm4nnPDgV0hFPphG5/aFqHMOXeMypw2es3FqybZd5sU
V1Qsd7r9kOGlUpMiHDZ3AlyCy1svmk5kfhV0Iar86KcqbYlalUFA1OPONu9SqiVM
x0bkCjal5/a7xTVuQh+JNEUmT/gBTKPFRFuGuVEjwArN4lsxS81Of/XVCEIWHM7M
/vjW/q3heJq6+l76njYx8niJu7DuUlWK7a2m9s8IBhhcNEVR5P6y7LCYASo0TVCE
9Ucy8FJJtjc/uS/vfsZFgXRYQcPIbgXrn2T7b96nmW9AblctZ18C93ZmuMLHkY2T
DaQTFALHtz5D3oaI64ho2ThCglWzSkcN3VSEKF9hXeCAg7tlF+1JGrUL/mGDX8xg
RyW/8YR1eJHUsA041R+uag5YvHHyfpAmT7xAv1yWJIUZZNUskkV9runCHHhbe07R
oyPmQ0G/gord23601c2SXVpmsO63mUULHd3y35cDEz+aA1TobWCkj/4BTfDKfMEy
RZ34MyxC3cRlWX8vsx0Tt0WwiTK8uqRj1N1ddiAw6a1s5q6CHrDZpRBEEI02IqwZ
jfjseG4wO9z6r+xaonZPRdaThmsI7ApQrY7wlEuAkVjMZTuyQ0UdaEO5rcusZXDX
s6YJcyUsmnQPCcVozw4Ytb9k9hOb2UR9TwSG7FC633tk66bxK5VLnrau5YhUbAC7
Q3nJMMfSRgCsvDX6YwpMJ94FNWDHacrImCT7+Zmm2bDjm0VD2t7JgT27g0ovdNze
Z5/2EM+WhL30J8dBELCb9woTv3P+rbkb0Arkz8Jw41cIFdixLdsqY+r0sihfRQT8
IxG51sDLLFsIIi7srhnuy/OvDgJ/bal9X0jNTQWGXa5qAtciziQ4f99Y2nb2Zmxy
dI0Xok8zEGqxJlzXbDXEvroo4D1K9TONqjbwFB1tFIKGzlmvQjTYUy4eakq7ixUG
8ZIZyiESOfiUcWU/I9PuTvjlFNEdhgTsMIwsnVeduWGtveICdWG2DFQIsF5LAFIB
D0iBIzYA3lw5SadFQwayT5IcCoui/cRhFo0p7BQx+V537nHCrmB4WyYev2oCul/S
Q8QvpCaH/xqViSxc3jRcFf0MHi8FvyE/aUZf9zww0PvUQyS8L8CbGDF6tjugnXtD
8Law8LT57GJV+tBp299yRlWx3LDi8FRppoxWNkcvYfHH0dNI2TOk2UkMk6BqQnRB
w4d0onvTxI7pkPAZBX6eMZVHBjKF6ttWGPKFqj0a+Hpygn2H8wOG1qI0PiwAokGI
koGiXqYm+8nMQGZNJOZhqdBCHFTzLOc07/fnFvWPVErmrYStmGvUbopWFcOOTxuC
tPOM71lNGkCQ7YD2sP+9Pl0xQy5ovk93z92TKzpM9lE8DcdYXd9hiAzQXkOsyvca
A+oLionbDPGIPzH3/FH8Xy77ulKvgrD+cHp4rZzqEMJm6VskFepF/5SsoCpiSufU
BPaUzsUSRmyU6MnJ7Mx73RbGQiM6k6mKaEiE3cuXXM31yfJ911+s8VhbjuW4I3rJ
afB2TF4Z5IpwQGsGtYOTjO29pd2U5xxSoqzsUTny2DiOL38oDz5ShUwJek+4ITLI
ihA9mMaMc0vIsAoQ6pvtBJ/EAw4rGlM5mi711mKHS/gzlnRtvSP/33USg+lnA7al
tiLJ4Ba1K8Il3hvdLlek1S7dEhhmDqT4fLKBypfun1HGxptLr8d8C1+2GeUuUxPn
kcBI6cAjHdqov+3M3It9ByX5R3d/MRFePHhx7e02o6T1kwqDaU9FAlMI8pGvumE1
T35MwHOzhwfjq7nQGGFrr0qWOLSarZAymMGMPiVKZPZI+VZ0mXbWIvpYEoVAuAWj
f0st3HzTtLFfR2VqqIlnrDUoKwez8mFakCH5iGR6isi1MG/O2yMjpMv0k4yHlii6
NpgPoH5aE0KiMRXu9EbogO7u52TImVZtnU7+bEvQxF6NJWKS1RqeCuOE5LgBT3Jy
SX+stO5POojpHe3Akq5e5gv1B6Cu3xnvmapAqKsj2O0MbWLihcv1fSAlvAapQei5
MU4i7/CPQ8d3D5DNRXJP0AhXCWKkQpzBYbYzRppKGfpLzQwJWAKfGF81Im4KFJY9
pVhrxJdhOo4Q6ptzEUcVJYU5Xa60X+VRqsJ0cW3F/HAk5YB/3ifioRvvrlXZc8+f
7WgIF6Lc0dh2O/NBzn3Avli23MLOKV6XVe8jAei4zziFHd4UhXa2ENw1/yORTMfx
e/ikoiUJHAvWsxLRlG8akHqMQ3+eYQ2GRRmU5xG98qfjAyL+nJlnd8JBSlup09sA
0I1IntHoi/JIQXHJHEAEVhyDh4+i3InasD6vt/BCa9UqFmkvB6q+g1H2Y7n+ywxr
Q5+8W4wGoVkd/E3fapXYuSlm7O9P8X8CfT+Uxf87ZgkJECFzFbuvbg2UyAiKFfNJ
Dn4gxkgqwoTg47RWE6XIQw//WU7bsOLq9DHKG938amKO1vml8Vjum6VLAGu+O+GA
SMHn9vLBDUhh1Blpy/vpK+T9VLolDDJ8G+/quctJnXPqdXlmiSwYBs5xnBteaEDi
UIu2xYFbO+v+3WvI+k4hJ6Traw7U7dFACOgaR8ph2Yi2J7xEiceji2LaP0OaeUEi
bncGj2XKnSTvZO7e1pHmiM4ul6XRVDcHOFL65eyYsmZUXT43lZYO9PVtuINuJN02
10IVRKB1d4bhlZQxUm2NanlOBA57qslW6OujMP6WAveYEJbB5lHD2vQ6rLyuMcU6
hCjB46ISaJo0l8LxRPmghOIlXXMsaJ9DH/hawjJhqBDLbXkxt/kYhtTFXdTCtkQ1
Yl2jqilsLNwTZ4igTeU6o6fxbPM8uzgn42tTahO7ZtoBNJJWA3Y2YVTEPowu1CAH
/mlUg70KZxppleF9gTD1+RB2/Uq3Nw6PqkNL567iLVgs+bqa8ugqSkjwWAlsARwl
In4tcIhy/5j2SbALGNKT2ZKKnudm/ccs240FZPsupU1knpVvYOw6ieZI8K68z8BI
/dfxr1RJdVF9CW1j2gxCsJOPbKkPTiJXCq8Sde9eiwNrvFDhiaWZ2hqjX8OJ5evv
wdwDKIYyQQOQIWxXuy5A0HF3vi8B/nUIggRjgv8c77p3go7ORQrrnPjhSsX9yQWU
ycJOAjJxi5nOfOtC5w7V/O3iiVVmkFXyQeBmUl6rIkI3YXHMujoADS+R4PT1VlGj
TtmYRIDNqm7UBjLTYoJOMwna8pF/CJadz6Fx6vJFDAi302aXP901Swx9P7uLaV/C
kYRt4oZ/qw+CPH7eNVUpJY/07x0ykR1qvGIJIrohr5ZEW+tZzkKYcL4REr6ZMTCd
qKZSXHpN7/wce2wJqSiy1gHGRlX7/msR0twDk52BycsbUOxWSOue3kTbT/KdbAdG
ZAV1z0nrurCbK093Zo8obllEqVaF5PoRHS16lqMiGB0VZO9gT7YkdDIZx2LdsVo+
gqb7+uYzJrGaK+TT4Ld2nlOdIUp/8hBu2+Tp2yZZkTLm0NHtTrOklDeg3y/rGjMO
nFgwz1iKmh3KwdCAswrn3LHJ4B6xsLVq5oyrlGFifAGHDfiK1cvE/BBx3h6uPiNk
1otlmlB3o99NnDluRxaE6mlCAS/gT6PByGFlbaKGgnEJ/y9O5c8+AQ1HTNEcZvIy
QnLSy9CMq8i0Kxv+cbgk2Xmg4+PiX7tEDn/IbCtmQYIrD1hZuMKIp7xtbBVpS+/k
c2xTvX2LBrozX4Tt5Wpnjmw1aHCgkHVvimpoUxkC2Y36NO7LTxqIW6aq4EjydaMd
O1nMDDnH8RtkWCy3SSMli3nOUMUNrirU95AyZnYXfakXvvqYhJysYNjZNFnP9A34
m/RcYTnwxePp8+2Mjta/PGNETXG0W5x8UatuURXyd2BQ+IUIZoMA1lNA4HwPQbZY
5HNhLGYOh+VOQO76FtI93tDZgAZBpPPuvPN8zWKOD38C7jJ8Ap7pZ5a6jKokyKS8
NTOpUiCp0uTD1KSstPv1b1K89acE0uBIFBcm6yhg0+3bP6foe+pi9EmMhuumR/2X
Q1ADuKvM7mOjDkvPRIWgJs3tlM4wx9efyYhOJ7o1iElwTZ75QExRwWMxDSz5F5H5
vKCt10wcbZ1MhLaHmmhSdacTs3OEhBXmYw3QUeAoua1eYEUmvtBVBsiLpeQieQt3
7nlWz6fdFVGynmhIOUMOdNHwxr8B1z1DZHuUEEDlY9VDgHhYoJVjaGl9h7o5AIfj
mCxRlHAu/bNpm1FMMv5NwxzHhPwQ1iCK5JTrGjQj4YqekVVPzZNLEH8SZ8sJaa4H
I6/uTiCluAcg88QW5iMvdXCKM8DhIIxPwwC5QPkKoAzf6BvW2ICkwhWdwrVocJNW
dPgqb6dS/jr9zNjYHR6nGAdx/8Znqc/NQeOxgznyzsL1IBsDgnT49JPlr/WYNOuL
2NYQhN6ppukogAPVfqHS6YTZ5Gz+lyFUwqmH0OnW+NW+jJlq1+WmVCXbQ63HbJem
jWLim64zW2QC/uF3p5vxfPi8IOC2quvuunl25Hf00VRbX6WwCgnxM3WCjdGaKYEf
XWEt8WXIAGrL1iEDu3mxn9v0QeAJdZj1r9eI1LWX95I+X2NftLHv2aaRN0H1G5wj
UIJ23oilFzeDaR8zVGiH1T28W3FCyoifHKlF2RdACSsSGO4/TtS1YE7dtdk0w8Xm
6fL6sr0VzqPKq/bUhNb2NdsmXWj3exJwxYtQ+gmM+0i/krKV8DUtPumFjm4bw/G5
w74BMwhzK3Rbcri/KvqcLTjvGKjkdWlBdqIaCCtRkJ1WY+iB6YTG/HzblKndaq1C
YX34rfKr81ls7aI7jeqKESgLJPrNDOv8vf3j7o00zX4cBBJoteDEqDYwpPgcJ/gD
EHWaKXeD7McWRqEACwmu88lKT0A9wfMBX9EJO/zOgWh3/NEXdYyyVInILJ1p8kB7
Eq89tjFBMr+Emrmx5AN4j2jAYUWJexnSvGVJq2M1mkmTKd3/6wH4UgiDoIu6B/py
jWJAQooEBuC4R3+vVEBORGnVTBsaNLwhfPCUXbWDOJgy05uCA0mAHJ2E8oiIBEE5
VYXnFUEtKKWmsZ3kT5XIW+fJ4fQZZ1LDtG8fBeeq29GhoSvkJabGdV2qGpBLSrwx
d2h37q7fOaWet8wKL1mJjp13vRM2ucv8OuAKyKEcNcOKQondnYdVQTqnHB/Dryen
w0qyEg1OiBSyb3YAeYa4rVYbEefnBPaj17RUdFmWdvKsSRhQGxJPFILBGjwOn97M
JIBW13NL3j0MNdDhqDk8Jf0QqGSwxKXSZjXc9hVh9klhM/hGvrt0eblEKO5EVFgl
Jo2Tu0e8Pt4S0eGVcBgIJ3eXpJS/hTtDuKH2hvGybvbfN7yG8b0YrHmgX93Q4t6t
TuaWEV8C+IhoUaZIp5fTqPyrzNtFi99pXVZXFgro43uEF2ulyY08ow/gspYTRCBd
6mdWlzVa0MB12+fIKSSlhXmbRk0Ov/Pg/tINglOAWDqs9a6D0luVP/Nxy9EOAABW
y4KAyeBZBZmVtm808GIarFg7WF5V8yJvMKVKGNLG3A6zV+udAgIg0tswIQPyd5pz
vI7qxecT9shvmGHpMgc3Sb5NR6P10Yn2IRuCxgdqQGYBVqBPx61/flc6BFNbXqT5
06bV8hbt+VCDXzGTOU2Gb3kn/IH/Esb6AO7wHgUkBPFydvBTRHlHFWRtVB/Np4Sr
CE0VGTKLysfvcYhCdmZSAy6v6unj+dn6sYVWmZneAocbM3qA3Z2IAUmy+Qc7HmNk
E4Ja90JVRImLCGbtu0sFju0KLqvdFTjBeWCVB5372OOXw31zw5HHucVF4LI6Eyqv
jzF+zKHhYADea5M7XzHtVKY42YJZHJqIyA3EQa6avDjnoYQKkbxkOsokuuXsLWR4
z/sZrcuFZ7bDPlsetDJrIgDIJVCkBVpz+LlpeqI/7xoRNd9fofNDRsPH2UvGU7De
suV3nqXGoahVmH9f4dJeD2/3tg4qpQzUcOhHnsGbjxFYxcKIg5XRKKjVsYGfmKj+
9Gmdo0goXuI5IgPzP1Uo7dCobHCtx8jbNNczktBcEkf7prl4xlT01jEOgbIEaIB4
XIJVnJ1psjVH1CxVAjx+LVCUIE8O5R6X3NWaT5vbagNAwJOVMRzC+UL63nIIE/Br
ST0xdnnSSXXFQVY9z+LuoKsX+8t9YXJiWj6JSpo/EwJb6jIeM4b0wKV7OQqLNTmh
ZUgESxJue83jef+nPjA311eJkBHREgWjl89BFm6wta2ra2mJVaTTC8UGZscyttI2
Y/8HwSxqwU9CXbMqrFtyOe8UqGHtUHONGPR4oN1QXs6TuoAjHDZei3NthGkLuJ5w
r4kJa0PKaw2uyUhpZcrywwj6pVceVnak17M1q9d9Fs0K9pRBCK3xtHoGSCh41jCU
IHTF0ttYrEnlV9XjYZD95Q+3VMD86Vvfh+2QH/Uks3LxBzeWQxUmwv/wcxHEaw8/
b594x8kZQLkIjP22e13JDe4U2AqqsdXkET7LAE/lce99EI3iB3ACMnleUIHK2XS8
41Lf0VTaise63BhOFjEB8i007dVGyllNIz/j3T1G/uMHiz1ytUGpiHyC0o+xqW3M
bX+GcxjXvwaSvJhWJopZE5l6AxEfV9w2m3K5NAXg297VyfctaxX5X07Ik8ahTTjo
TovVPoPqAViRWerLDgvHYWptkffjV1+cEZO5Q0JFnxTuRLXyo4ACMNunrw7EOrnj
PUfVXi++EXTP6lsgVIuRux4kFVKhSV0r+4eGq94WALtNQel7W5/UbnREx7ENYEva
RiuEiRY6u9hIZ8UGg8Uv7XxStyy6y8O4dw6ai8XcZDfHDZwltqwtSKjN5YYDqYkk
s0vfCSSIaZauwQYNMZEZ9e1B2xGlvlw0aPbIRKkjczn2ronKv49aLINQDHQxuT3H
2cSvaS/IbDiayh48a9+8aKPhkeD2UJfc6Uu+EzmT77Aw8wT6IHI6XFkLRPD7mIVu
wOO2kn6mzOxhWxPrKwrk3n3ysB+iH1wMe3aQsH+dDHSuFT0/Ck0l51Sq2xaQI6qs
LhHjcc4GgSFK8W+6J6BY4K/NKr6vLOh+8r56ELDvkrmQ/ZuKUB1XEq7YZqawsv+e
TzfAfpXewRBs0aMqq0koKriO4Fw7/T72Up1lDK/ZKkP8VqJbf70OVnln/jQ9V/SL
F+3psZU3yhRdDUvEQvhc97f3r83FYv9/UH9ghs8mKBwUbSLIoZRbEKiLOlr470nv
XOq7f2MXJJ2DnQX6qiM9HcdVJjKO753rZZM2zdBNki5BDBoQQoDwjw7BCDNXaqan
jsY2EYCB5HiOZoxnwD2pmnb+d/e+Eje0bl7EvMNdcCBaWTd/DBHhnHZRSB05y39P
DuaA/sLGQuDrcZ2ceYHn9x8jkzYjGzRB7BbI+A0szJKSy1XafkvLM/DG8qnhSqXO
xlUpNtcJnm3Io+J/HTURCVkI/KbvLOKeYlPdNKT1jqYsRFsufY5lXegDkMp8f2rX
ie6klib10TnK9s+N+T3wmA+rzAEQDW+GZ3+qpRzBNQ+QHFxAKgoJPWDh/l8lUNVR
H6JZqzdo7GrPLXaRb0cGzc6bRsT/VMO2t0/4JZA7YHPvN7jc1Mt6WS3iRO8AhG1q
0w2Gk/nYZEdxiRFELDcHsgRQuoKFQrHcGq7EaGCOrrUD2XQkW1/1zI9S3Bpj+h1+
FQGMoficqJlf5nTdeMHdxmxkYOCVjEJNDHNk1HuTah824iCQ1hMsMjIORILeNy/c
L4JfmDM3iSkxSKjmbbxptGyrYQwsdJbSaYXTzThU4FftUTQdoMlqxm0Xs98L3bbj
8nrpbaZeFR9cNre0mw3vD6DHxAIxg8DK9MnbxSbNt+qWOaQd7xZuX+mm1sK7UOCf
ZcqWfkqJfPLDO3E58ZzY/4Rph0hWtx6tTDlNGqHkLtzlctjGI+JEjXk1WwfzC37a
L0ulCex/yr8Ty8+kxMI7TNSolRuADB410rfXqwQHpIzyUpLPvraqZsZvU3wFYUNa
cONMcD5tJU/JK21SMZ534ZJHtcV5UvdjKaFu1AdLhzYfAAXBTSgQFi3ucndD944H
BZmZgu4mWggdojmZgGvGuFtdPPhSllGkW/JX1iL76d9/8PmVx8PwPu25ljSjA5nT
FZinyFSVr03OmVeJ20zShYUeKap8zDiHGCc2P76ljViGh/zDEFKXCUpgNXz+Mjhu
8XXDdH4mlWQGt++MJduNwah1icR2mKY7RUuH+xp73Nk5ktLdWuO8w7lmx78SxNPN
9VtCZgyQDT0rG1Yq9zieGq0vFDh50Jf3LJbp0j62rVeXkxs/FJvob7WGJQB6Swke
ugnHaLnjlR6ujZP4uHtFyARc11pLGkxFikFvThQcW59PfwKzmCxvGN5oPRme3sEW
7ViOfINQq0y8hthfxSAfG6T9aWFI2moes0jPuZIbfmc4n88Qn+XABGBaVN9spRt1
atN3NEpskXFsQOhj4LgGMvjnvVTvZdyYWiCrqn1Dwb7OnFAkOsnA+tRzHQXS23TY
a7eIBtW5Cme14nChrrPmDu93XSP3r+ohrvpJXpR+vSRZihQLFRZphkX8NSJXAwda
vNrinchvCPqlHH2r8M8yg4YgJW018CzzYz4MPGwSVeGOdOP0TkiZS6625zDrZrga
wErNGVyxA8ymDBUaS6PdQBHq5Er603K4e2pMPVHXOJpV+BufLgLiMh+jCPg0uV1c
LSASBo8x8P1kFWZRzUQv1rUCL+OVqvly2Or8jqdkPrRproZ5q7CNyZ24OIj4rNmJ
IFFEmj1p+KGT3EkunsSMIe387DlCmo6xnt6Jt/XtRLywUiDqtwbzxckGmwz544Iz
ap9l0fGJW78b9hO37CiiYTqAYBEAbXcbHjQrZhuarQozIL6zYqszVyHf7cuBWizB
fk2sy5Ff+Iqzs11jYAaZpZttaC3BVyl9bqzMpEL4V5utk/D6PdIoqUKhaDPsWlsg
UYFIHUXdg2s20gZ10yU+v8Lk9Z3p9D5q+Hou0MYsMUwrvcGeY6VuWqBbAFeem4S2
EwoSSJ7Xl164KAyaeGlri9ZmjGaE9eqm1S/Ut6+ERSnrrrbX30Uitt9cC9uoiYwv
run+0MK6PapjJTIfwmQuWZKiplCtyH0tVYxsB7b11pKuRdeGgqyqyaut549gtjBK
fH51wC4Lw10SZzODun+CquFRcCOwi9lJRRdqSbM4TJ42dOQtKLRuZz/1g5nnf1YD
qDVuHnxc977XBT5TZhHiH1N9jIhHkaxuukzh/0UQNUwqmIXbtHIJ9hUAlUs1rGW0
UyUAwbplK+0rb7l5ZOj+fclL0f5dFXNne4P0O5Pb0lfZrOsmi8FkE+wwESPmME2l
UByh39/Awbs3nqhZjac/kUenrJA0BZCLXY/Prti2b9RqnX24f3/GWA/bYc2lalt8
aP5uw9tvTv2ATMDnvLX4TP3a909n+vJo/U2QSVGmSKZM5YMJ7N4IlYzqNPEhkq6a
KrucoRRqQIeHqo7CCgkz8vPugfdD2AzOPSm7Oi3lplCGLQNHrANVSroBQEby2Jib
+5aj5yQo3i61Cm2m+bBNv33b0/RBPXXwDcLcBv09uHkcvToTT8CrCLPHA68jFPCq
PqEpjcXbWeysO1Pd0pVhlrj+znWe9xKb4mh20cWKr9XVmVqCRa3CUMqK6kBE3ZDj
9ILHTRlp3xpH8CLQ+AB/k2CnTAufgESdISzsEAKU7/24gaFrSaBRFZxX5UQYAD6B
jdqHg8CCoEX64Z9M8eVgIHBwPyJbQN6HwNd5O2FaZ/VCcTca1tk4TYTLmCNTvgII
tjZ0AkaDlHcx4ML1XAPtaGwJkvrNyEDaCcjv0WAggC5e3hmwIb5FwZ+C5/topcME
AUSHW34ehcPUxwb9925CmdHYH+iXlwn3yYIKvBT2uCBddNm7PP5gj89nd9zAQMVk
Z9WrRkYW3FezZFQw5X0/Rqg/IAsbBmVT2tiD6dh2h0ZQn1r7M0cG2uo2wVR4wOBS
qgqs3zQhoeBHN39TcXeLU301FN0wSFFmKzlrGsVgW13lfOHGueB5HbocCMc4w32I
UFil3hwuMo3PMt9C4fbKAEkrOilIYjLtN9eK+F/O4XmBXqsu0gc0UijoDYPdF2fJ
RuoN2HAxf3EhUSWd5O50pdUnZp5SjlQZQLBHEePBr42pIRnbJRqnc8xKUpz0bKNJ
uSRa46E6JKOcT5Eitj8K6mSjk2FYqAtPx/TlaBEAHHPwRbCmpTAcIktkuJukoN5t
diGsgSKUucBNDMlY8KYNgXkqOWvZV3D5txqvu5s20QxOKaka9x8O/qeyTgkqMuLM
tv2iY3JLaSEEulRwbw2UBatQckcIB6GAy6ixl/vKJKDU8eR8poP1Hvsfnz6urL+3
dI1CmjF4Hla89E94tKsrGUwQnVGj11KbtHWOxuCM+pHPXQz8K72gplOe5X00l8Q9
3QJrpM5FPeTrkAT9tMyAtaCZHV0Tq58OzdfVigl0SusP7Jy1e6zrqinxqWNQIfYf
0vU4xoY0syJJIO0xhVi50dnI6uHxbfG4beKwFpwANdVDgvu6gXaWtK45zqdjiMpQ
VjHUust1LOGkMN/A62hDjAlxpB8TCT/KRyb05FuOC9BoLDNpkoB45IvE8Xi3uPtY
N62d1YpZ89UsJk/Z7U+DqTHMUVFXAqp2DRilqnh7awzIOFKQh0xYpuIvRFu0dALY
xMO3I7X5vTJypHkalK2LI/RBhTnK9huBDTwk7wrNboir40A4MywtB9Ljpl7jE2ao
eeaelYVvm1cECxwiRA47qfING+bNsgpVXAFtf4qGWEFx6F4HxFjZ2Q11BQyhbopP
MLC5oP4E6q49vT0Ni0Oe4S4byKt0MEUe4qAxaBxb6eMtUqhZR/Jm7JKvm+Uf8I7W
Pix661WdMQM3lIBuJp7yQn0BCtFrif6DpiLyNpRqUEwfORZ4qQzS88Vsg0n1ZjLA
9EIj7zayuqrPZUXtP08HhBqAVS/EabnirojtSYsjqnB7Jkd50jTx0pG4GhJgDy6d
UvVs0576FvJ522Vn9uUBgqyBR9qFnGX5OwVL+mnk3y0t2PrRVPgtCRhYvlXPQsqI
EYAOxaQJ3bQ7+RMvdY9iP/gt1ZQ2YzoTpc0O/36sXqVR0ZXfEwvnWB1ihkJGjY8T
Y2h9Dm4dRl7J9ussxFrVgwGYQRJ1xVS6Tv7ovH2mZ9BCD7FgTJR0djiYajoLM7/I
elIuySqaQZhtwJf56CMBTHAYT++M3rzMML9o/qBG4jTKQ1R3nldOhs1SPkdmZXoS
Gj1gItQNuDxbFa4Mnvo+sUVdPkTy+OcVaKWGRWOMPnxD8LaIVYEaoLMr6xHo1/83
tbPTH/SxNaPTtvOZoit7by0AHcteW2B9Y/ves1zKjTX/FQLaABembaJNgnRLIrjT
HU8RQTXUHJURBSTg4jzzbDKFGZmia47DyLB6YqIBa4v3JhishBedMCWvd+Om6jed
lFnJplHu4AYj1+bvXGrbfdsW31JtO0IhIuCGsMJsC0ZDGKZR5fUi5AlmoVm8ixFA
tt0ROEel6xqeIvNf6wzKpxuJ4QL2dcT3eZYu36nIz2Uh5u44tZUrGcLqT+UoeU7l
SO2TtBqlP4xjbivPyI8/fzSquz9F5IzdiOpmfhYRY6Flgf+/Q6wPSWEisFLDSWya
J4reNkB2xRcVhwTt1Nu+qp0pDbO8zVDc28GLRwdlWNsQl6JAZ0rfImsPuq5YIMUi
HJdXz3MVwGlth34du3OYMz7j/kLIIed/N9ksOxeYg3mQg992A3718fO7jlmL9Z/S
ws9QBXCqAXYQvh0SD3JCgpt5wM6SEJnXD551FfX0bhyQDhPKt0eoY1WDCuLRLs4L
bExqID5goyr0u4B4ZAZ0+n01f/73gnHb9mHRy77lznAhbGmgg68+0WoUhyyiXo8G
YItayLYrJYkZQzLO5fHOezpMcqp6ufXpVhxV7wyOYPH8+Ol5QzewzLbnyo5BTP0g
eh994YwcR4OYPO3e5HwodQEb0JEk136h9oRGqF4bH+LlOHpxr8IkQOxu1QVOUQl8
HQwBBPdp5FZsxXB1ZcrCo0GG5wPXgyxntgtsy4t+DeXPKhUNORjFBVBU0MBWhMHq
C+IL/YViR9zYONhX9+0XG35oRRAce061aPWikcKkZ37CmufKM0s4fZDpLTeHnhDu
Rsk6DsqbNpRzKTrwUnTeyKdRZjVt4z+0VgnosMQhXXrbMrXOCx7NvcKHgooVhlQx
5UTvC3JKaVO6FklMxy/O/RBKg4DaWztMUOVG1VsoBZyGByFz2/qSnntvit9cXEeb
YBEnozwuxGK+d1aQtUafiRuff6dPpATDtFcH541DfxXWK+C8pAeWD6ytxhKeJaZE
5RGTMUa5rUdgt6cl5vpI9tjuga1am8CpAjNbL46dNkHqJNv6afG4ZjXYRZqtIORn
uFAnrUn5jUWJt/X2AbMM0CYauPG3bbL7lCEwUnbdWacYWoshPAbRal8VQ+TmjnLF
Gl5KAiC+ujuZ9ZpfwcmHy1u2G+4NJ94P0NbCj2OmMREkm5uUQjUiln9jF/8Woh9T
u4pIJmebvq7Wuu1l5tyxEYCLqt3nNlDkl7c7aYCvbL45i1vPKV3GWm6ORa+4nzu1
MQZyU+CxKgfVuviwUMEogac9YZzPutKLOE2Wfvp3tc/H6R7W/xPXADPbwmJzFyip
Unpmxt3qbayYATUyaqzherhc7qNW+4Wg9SgvXDEmN/6VMygdBI/TRivsxNAlNZ9d
TsWtRar2qpDNmFFHAaaHEVu/vvXcA91wpUp5OyU8v9aU3j6KLNRgCbEEyU5GXYk/
6Bw5I1xSMNSITLyFAmtfxUAcDB9uKqLpYYj5poDK+Tj9pV0N1Or1OAmefbX1kl7T
d+EEsbG5QS4fNmhXpIjqz5i9a1RalerUzI3LRwzMz49hssPL6G4GSjAJxTt6PRHP
gVe5lPoYUoLPMzV4v0i043X9aIoDMY35OPFOLYH6Ib2mrdbAWsa9k2IeEGa8jyp6
gPIoO9v8t362SUI2OFRECCoZUExGHBnYi0ZW1zak8qYea33tXzPhKwGLLczS7+ux
OJzIIJIYOLojqqUMV0ITaqwJcBpsWivEmhEzty55bhT7fo1buwTjTJce5Sz1cTgZ
/BWWtUNemuiLWoEDEM5YBzk82JXLO/WREl/p2LDEce/XzNrGAgEA6W2FZJL+5Z7g
9D5Oc2Bcb/+qCf/OmK1x80aEJWdtj+wxdoWIpe1zem/3yuS5Qqbj/Jltruw/F1HH
AQ5Aoj56fOhIi9HJnU0n4m7VXEjLyxKxFNMwLe3IX67njCXJ62EwlzpDpyFe8MRp
vaosQRfb5bk8uK/H/f2UWgZQizjWQYmwBbGrebCobxajYgbLB4S+okB4eR82wFtT
OmxPUH04rnaa7YmWLJv6utDBIiXLy8BCEXLcveblj3PLJkd3xJsK3PfIhdcoG4UC
k3POEHMzvStYR08Bh/6RAQJYVFeT88D89rle2DxcCAGY3XECYXj4moy/xJwLyFsw
p9ioh0JBiFd/4N768L6llDm23rCXgFxdOx2ia3QS9AmQmkx/BXCpu0TAWBZbaR0J
UlX/ry9HZDThzQKlm7G6faHYsVBjvoHRuDQ4Fq279Jri9IxQ7WjKkGN1vGFq6E0T
PEkzoGu9N86Vi5BkN5u1j5rXfXXHlHH6R6o+O289X48HQbTNKFW/TyC/L5UxT/bT
LS4R9OicTttCGH5Qf/Rhpksayba7VMI3nFuoJRKnEZYQy5EpNAtvHfNHIonZIeQZ
k21P8b1eN/+E0tHEGz4WTdGKd+mK71Yypy4Amgth3kGQDRTZoRp8lmI3ytKA51Qo
ceZ9RYcjcQOk36lFIlEq752qF/TTMJzxvR9QGb9GaWVKBaWIPHKJx5X/NvxmB6o9
KcDVtvoRBt8OwJbKmd4o+xtIFF+K+lAOAm4jd6KsET+J8/SrAGBErOJcMQQqVLaU
0rQxPOVs1FS7n9S3CScqr+gL66E4VwIg2DNKQQ5bMT9Hujt3AozhGyXiDToOfaew
Niw1sLHDydgb7jl66W/xRjUVwZ6AO6jU7PJt4uSUzVJDCp40miVqZZRBj6k21vMN
TPW11f0/N6bw241ds+il2bbB/HPY05JmOa6Q6G+ce9AHIzTAg4DHfj2ZEjuqRu2W
HmIcf5Gdkm/YV3oBlkqaQSfmGGDD5fYWJG3g4zddQxUXK7Z7n26PlaPEy4aDJfGh
8DDCFMvRUU/0KTW12J4gx+z/BiqPHDCiLIJPn3fV+Hlctl5tFA/nJtFpQMrlRXJU
fQtzzugZxB/s/xV3h4oUGrWD7ob49hSjF4CWW0/fXZAIpuMK0iFa3L8xJ1hKcmUI
NQY+mdysozrxC7LwZN0xsx+O9P9ldIVJzoNMWvWOcMPVElcgjPBH4lIR1/IRh8B3
Nhl6jVsE+XdtexSozqpvr1LfK49Bs+nkxrhaKnQ441TxZ0217je5Ot0hBSSB/y+A
IF2rS2luBnShw18SwXyq3iTnPCYXXaYxnZHHeD+Yqsmtgu6BjpEXkmzEB7qA+xmt
Odt4aTVACC7TxtByjw8pdPxqHzYMrfnMWSohOps1bctN+4bJivcjr35EgZ5V0kWl
8OK/vTfB3k5Sc8fpzEZCnW4Rj7R6+zMh2hN3+yW66WY4KYEy0n7wIz6IX8/Wxma3
Pl+xWnNGTm2W9E+OUN3Y4YKok/fanO+a7bFYZ3ET1wbVfKsg4dNJ74iGP9TwPsfT
SZWYWZQdINkzDIqvdunPvjqsSIwwvdBtozT9Rpb20NpPfctjyx1vFGIVbz1YBmDd
xMsaBU3wcaCQ5QSQm0Bz4Rlwtvc64Ru+Ow0KV+qgGWY97xVepsv7zpJqiL1g3tSp
OAGY1cbXSvRrvBhugpvjiaexKcuh9aIB4afqj0OOnPT9JEoMMWdWydzzEIr0KmoB
wvOT7mXLmxuTYqjnBSwgwn4ufEPUyGT+DCrQoLQd5zQrVYiYczXh+sVYM39r9d4D
lD/AjuZIJAQgcIhyHZhLqDN2CmbnUsNMn1gwSmsxh1/rqdzHkiXg1ODoDkIFFEaK
a3ha4KUkdJhs2UOuDXvhww74AXnAz3QmkWi2k4ftMsjmwCWBrx7VcN008MIZY+0h
tiajYmyDFdw+y6HqKiX09n84Zex8o9iyA8RhJmB+aKaXdeYZWRaApRzGmcfgnahz
rsXgGbjDpd6zOui5YUwTtiuwvQnQlDiWCK+hH0cyllK3XJIMTg4lIpMTur3kw1JW
N44nfwxLYhH6QovKXkXFGU9iJbVSZ78Y1mvl7NlwCX9Jrmw8iF1ENbs4rBtoaqWS
nh0z6tdOUt7G7YgpglefLIoPNpN6cP5v7mCodLiNK615J4diJTslSpxn1QDgrzvA
ddo7++GJpd3+60iOAX8O2ipwHLKmRwtFdqki1pas8XDt/fB3vsiSrw8yYn4qNzlE
VklZZZTB3wykCQYvfB88ftSxpTXDQCrcNIqyDZinPX4yEC8s/pIwQXrJ89TSTcmw
MB9fuXHGyom9HQpt/o056r8bF1CUm80/Qy3QdDwLs4Ls9bgLsh/AUIaGjMUZqjAI
jn5fYMFADcgg5eGBHOaXkhU6DP+tBUYIs548WVVK94Zc8NTkTs4V/5MmpDMiK9Nr
s/OV6/l0tM2c2S/Vlkxd86GnZ1VdHNJA4E56b73S81Xhi3b7hh+jIcGLonLom+Eu
B4cFjsnuN2bMflTN7IjJeqliuxVoVwjulTbMerl6KIBXG02UnlcRgg7/gkNRFbbV
BDLQG6gZhI5v07NDdSqjsK1jeVvCTUdpnZhAxp3u/xvnjEXw7+PMXwmd1ParAW0W
wt52AFd8XgLOumjBS9ZZ6Tn2GaHHsVa6LDK0nrXudMPTu3hLzC8DdmvZ88R0yUEo
LOSr/dujJ6jmBkadlmBQVv6Lgg0c6561OcQ792UPNrhFXSEn5U4PLa+PntGXM7Oc
JNhwEPZ1Q/YQLdN+h9lb86/ZYyHXEeDKJlWyrirFADbvJfGklC41LudnBBzGLX7K
CR9F1445uhRYvOX5e9+ETHN7X7r/pyv6NayBS1Vs5wWGgyPPDE8c0BhNUtm8Wzq3
zcVDnWp8zd3qA1onsbCS4csDZPGi5RNToYHlbDqhMH2ab2pzDnxkF8AwQW0xW6/h
r9mzGrWRoytK9/u5I1SX0e3oOOdlRdnz7h4wneUjFIOrNEAeUpRDgfS/vNXOiEhK
Qm/bmMhCz1Y8ZnULLq/9Ln2IbSVKQdXYpk9jJbPaybFXO3dS+66OACzkKs7vwOZt
tYRVEOOLcS++Tlo6uoa/sEuE+E0W3kabUqsSCGSNoS25mNoCUlfyPYJ7Mi20zhxX
1NfYOdntgFZob697OhXN9k7vuTFX3e8rF3qhUihxeEryVbQzZu5Tb+anZkt2Kdw1
g27RiUc823wDmmATqRRdBqCj0U0FAzqHEFpBIeag/UJmBegyYBHT/QCGG2SiFR+D
x6yal97FPENptecvCif/w8u0s5BAjo/6CtAdbWiWEBZQMGRFF483CTuF3CeDrZm2
RAXTho6Ow+lHmCdve0yqvhlXVuSg0Mm75dWeBHfissS0j7o0oxsQ5uecDGCuR1Rh
M22THXpD6NZ3On5dOwm3RGXzKIeMEzW7GBb2eqtHTuPciESSpmDWVn8M2i+I/w2+
TXbqZhqnb21NUHl8dHY0Q2uPne3vAHaJQV+I7qpDe3QUhBpHqCrSgdqsKUVaR9aU
Xmjp6IrlmqqzXzggRODqRs1lAD58Tb86wZqKf4gBfIycT8tBf107lV1cMFE2VJ66
88MoMRmG6sNYR8ZnUueZxFsVI+D2GxwmS6cwOUAopAYLutNBUX89SeTIct1bc5vm
sqOTiAcVkOdpjINK0n8Tg1CMhmyPEclA1xtrpylwuyhvAi7SoZvHJQJONRhda/5g
QYqXU/gD7cPo+C5/O+tZ5zt0NT84LkTXh440z3xOmkQQS4VXH/7jzL6lSP8//dLf
LqjrQSSlWKZEIkdvj019YlboD0tb+mgnLxzhFuCm3rmTa7N0pq8A8UypZ4B+/Yiu
gS9PslMVmAs1XUo1N72re4ka2SmIvQKGdVV/Dlho8iAfNHe2Yt5PC3Xiy2f7cuJv
bGj+0rQu7AjsDylxJzrQa4MGHgiQIugvOT7giIQKLbIlkYQAOQeaYRWHFuONUn1w
Y+GvdvRp8ghtu+zGRTl8au10Rly2Um/R87mZnHmOLSr7HN3bWo9E4Y/JuoWKSvgf
Oai8cwV6ZYOtenm3mmCQXq1V3BmWKsOxCSVJq9P4/0eLR2C7E6wPrlDfOXAeunXx
EwSwEvc5WTyJ+IM2Z24Wmyri7q6rBj8NTYGD5KsFDkQ0EP75SV17znSRnsQ6yJJL
WM5gdC4XhQcdJYebFg3S/ueMgNEHcVn0MfGEimDUkK5chi9Bn2Z/xeqr60w2tN91
lNKo6rwPO/yf8wy0kPdk20r5C3EEGC+UrokdcINCy1M55D/yCm85kQE61ODOeGl8
/vsbbqicXEx2SqWxLuDNo9ArMHsVrriSfwf+2R18o5T5iA/w5KydMYoC2j2pjtXu
HQPerJC85KWPEikSlUc9YRnwEJndWR2zwZwzOkTYSFUvEFGT7xhI+U3pr42N7jpa
GuZGLfY/4ji6J8PWBGFl0H/n4fvS13uXz5ssoHZep20eUeqxNvsdDSV6m7ajfXWc
OUmmc3CYa9p0Jun0uiFXKFKrgNmT+5ZAOSugMZUaAlfKGk9A9/xRogIrIPC7HHMB
PnjejLkvK4KaMEjdIGjiHHv0jWAp0ga4AiaIwbafVnPvIR367ZqQZrXoJIHEWcvt
g0JoVcWLdfLaFmK9m/IKu9xHI7pj53K2lY0NxGhjwv8c/M6phTe0q/ETssu0MPUv
Y4yjBmSfuoVnUegQlENn4Fgqyoe+RzHnxDg4hTvH4Z6/UkvqSx7/mFobx0Rd9kaE
qN/ORz0YMhm+afpioNdQxq7LVreRCRtlPgyNTM7Wg9YHENfLMvGb7PHzhQpK+7AW
ijDaXm0QIEGorVROkhPakwl7MPdRXhKRYjrcAwthpOfMmu3vIcfFSpdss57LHdvW
ziIrkDdoI0ye5+VtzxksR0GRT81MFKN/krkNAwX0SUClKsAgWxgVjQSWM64qXTpv
fH+nSTszFRRPTjiqarSf2hEWdw9Q5DHWQphDPaljciC3kJJpLMOPOuWPyk7kXXDn
plt2WtJismnzmjKE/gy6PaaDCGtCDIAVcoQK2zfHJWcahelXKbzG1DmNC+KS9fK1
aqaFSjVCLXGF/cEndZJ0vWJ6BKo8Afjb42L+VL9fUHgm5HkdVJNaHMgKM/REaPx8
SpzZahQXywA/8rN4z+n6GhTMJSEEbnSUGhzc5epSu4ulbtR1ZeNJR0RZJaBor1Ta
hTAfJGs8sZ8tGo/IBeEuhFBcsKz+YsW+EbsFAFRXAJfT0qrDrVO87nf0NzhPSUA3
Kl0zGjkkph5XpGaLno/51f7LEDTxzv+B8gsTCgzJ4VFths0bROae5dkwooXZai9u
NWwM0JAZBwdchHvAZA3LtybeF+ei2pW4KcVzvAamaXyg4Vc3efMiVo/678tMqfEi
hiYghTMLeKUuAoBpgqS/HlrqaGw4Ec5ckEI8bBXmbzlmjfy68KTPOK6vMXVhyY2X
jQPDy3PVUPpOEOspwxL86PE03QfksMfUaIolUwxGDi4dEKQPGvuhVAP6YDeMlGFP
YKFszQqnMrBypteEBmpxEAik7oBjOeNbmF4gZGa1vC7x5Qqo21O4yZAtG8crPiDA
4tD9vUjRosNSVCMA3cXfBPVBsDGHpEdSXAdJ3UyMNR0lNq3FNpwbl9LXjqIYIwpP
32D/7EYSPpjeIharJLgncKhBfIXE7v8neHLAV2Lr64Ch1fgUGIzAii6ZFJdJzQU9
aL5HYJuCHt2LHFrUmgF4jAwQTuNY17JKf6lrdfg/mZ51Vb017IA6IyoR03bYsRhB
lqPy0opaThKA1Pea47ByV9wVmF4UsjOre/TbHAlW6gs0+1k9kn38lJWfB00GRsEp
voQ0+BGUbyhHGFHx6spA3RzIrmvWIxO8BMm1+7Zhgl8NI5ookTP498yKS/6qtbl5
qWg0LFh7VjuhJjBTibOvFnEkNuvsu0YwtxywpcyJrfI91YMrM0k/H6BahjnbVaVL
QI1b4Vnut7C4LnBj4yZ9yonu7gO6r6lad97TBOk6k9krYQStHhI+9DNHv9MAaZl6
sqKthvBUJZf5m5pmRL+wR21zic4318yVP9LCTliht87tbyEPWvJpUq1XxP8IoB6u
1kSD1VO8XhDhnRrIyOacIlCcEJeahaQFVpGH/nlHXdlm4kh3O8k4DqvLqLmuI/4h
V3x5OxwmPODusf5LLiYKvKTqi5eQ9QQjGJDGJwVuJ+Bf6IzLEpNlCqeDlPwuEbkM
pGtL9GaxnjdzrfVNPQU4TJwW+NDe2Bw9i8fhXoGuSnMJKiAV0plZ8pbbgd0zGPFv
ewYk637Y9padFdUc3EHU72FPIi0iBH29y1jyCt7JIyVT/jb1T3lC2XLDZTSmJqkX
/AUDPzTYQQF55bjbUuDbBgITHtNpFZejG87zcOzBGxZn9Uq9QD7lvEO8DJVG7bqA
vdjMiujMX54olrkcE4KwkDM6XeVrfO4ZmfwkZ3dBEeYGGIvdd9SWf8HsFztNd/xB
lRkCXoeH+4wqCOFJHajeCA8u3G9K1OZxH6CvhU3madp8BLEiuYJss9H1/ubMnd5y
f3QAz8WpydeA3qDadaeEDCaPZEk/og2j3W5EzBwh7apoyNo6624ZqFLYdgJz9UWE
n3LzFZSqceVW88YhV221PgfuSOzJXo6hw8tC4gcAQBTszSAyYAX/OJAJTm0ay3Ww
psKGCEyvpUYj/twJ0B1JemP2poecJzdLN9pAQ15oUV94HaQlKdK9m/BrRUDhNQP6
tWbc0LlxoQSJweuiryvdSYdghZKaxr9Uxnf9npNBfEG1eMC4XKs0y/Xqiw5SGZty
KFyRO3AcCibQCIc47kbRBxtSb03u1YKlYmAKfk1qjaww65neI1FaxpQMDKlFJZZJ
j4cxD9OWL/3eqVAMTItdsatalM1swVrMyXtlF5yJo+hGqZAyfcRQpz9iZKTK3vqn
GpONxqK4BCKx4G9yilYue9R6/QO0i7gs/xAfue4KtLJQSra07x4y2ISOuSUoJJcI
m+gO+TFcZDGZmBE8arm9sitUGu1QWJkLpRsvZFGWNuQZQj+bHhVGyD2d/i1zsSBf
mfhnge/I6hqsIa8Wz/eqxcWAqm9hudKeZOl6TVB/Os06OEWRqwlIdinIapfOWHYK
XBGFObBAF1tjgw9EoL4dJ2eU1BpCJz7A157gKeu+TM8TlBUUMsqcnRz8i+v8ExqD
A6cLR+kVMYZLYJnVzvLFgUfrT39CuYAcgR2hz4n+yuOacodACc/XtOc1nn8aQfoG
b7eDChKLi/FJ3gFI3Z/KufSE8OaQUyWqBQGOs6r1aeOiQB/T4Pd9eEchJbrEyzAe
XPVMhHYOKALbwhfwui77MY2KEvX5KEI0Ic2new1/s5m2hstD9NTzlX8w/I/XYiHM
Ld7IOxR0IFF9u7nPqax566QueDEYjgvpncJ2iULFmw6YdmQyqs3B2MmYD7DO07F9
kEuHM3HD83TuSJt/+wvqFHFGNyb0FEmRBZYVa0yQE3PfY4QX+UES6ZpkImngL8GM
q83VWogKNUWmxOECwoVSTwyrxEp+RLDhgf7EzpQW/2G8ACATh2Xpi2vz0rFI08On
JsDw03QotbrVB05C7XOdzJnhxtC7/2ffqFygMBg6lzGNZBmuuEHCyYvUqyaRZMsU
OM5p0jRhgiLIvYfiqasX61OSyz7Rm8Ra4LtqWzX2k0WTlbOUASZjxyvcnrhMXTmk
L/HKyfB90IHjsNur9bN45mTDHBpk1pbNzmuNhomXk3YDO010qiLphCFvU6c8MV40
VgVUY0E8ETFHxbsBUU5257KVZudzoEMuRgySUgRTkdqybtpyefMKrD0vBli8+Pci
J6gIthXni2hq3FX1fTqGyVvsIiq3Gzml7GVhoNULBeHsR14NZidX1min5uirN0Fr
9GXuz1mIaJzVGFsSXRmhm4Dz7kxWB2RRD9NZhKFByLakxffPRMCjmHS2Uh9YOoS9
bOOlbQnjLSxUigSwF4etTeQ9EykFyp2OMaCt7lKEMhHSiDVMFMV6pqHt3CbGPGK3
8xcD0Dwq6Y9G8xlGuWRQQcQoskk1jKmDCasm/Yb9Tj9IKaflyllAZE3QkenijwSi
IxgWfY3GYUjkF2YoPdywXBG3Q3r+PZYCMvgmEPUR0wTh6/vBwPdQcULKSuuT6PhE
Up/8nat2hU2gK4UQdxwr46zhfLESuHcPaCt1cORO7BQYfPBN1r5FeQdxHW11dM7O
mkJsPmygq3fO2BFXdQWdcpgWj404pfbfAwTOGlo+jjRZ3R869nZ2D7QTFLzrfXm1
+Il6+2RgFGFnr/kzl2JYVU0oQnK4fn/16luDEZLPjyPrI7EmxWQeNawOLPZbQND4
T8x8DaQchYszU2g4KujjUfNX9JYXp/t0UuNGAkTZrtb7vOyZ06qv6eLhxbVWc+On
E6dt/0mzSIKJlWTwQJ8uhcCFZgzsQoO9k+CIV2y6V3VmH0k/8GtyfnO11VU+mi0P
JOBdrE5RiJ0Gj1BAk3VQSH+lql2krtk3YnJO7Huhhk+KGp7ROq9Jd0viQwEc2aU+
eWx0D5fyDtm/5uprl8aAgovnse9SYia4lg6ESLH+6hjRYWqkChpPHsOVwIAj1o2r
iestVjgvGcp+3UbkfXrsKppadvm2SRRtoGeL9RvULx9eUStwSZ7W2jd2tV3rURDa
VCIl8CTVDa2d4wqUcHCADfYtxrHNqT7/v3Dut4aivmYK+bcxogJJTYxM5n6kNDbL
EnzCzY2wTy+vfEWkQ+NtalbRBZdhM9/LN6qFsjhxysuaJxGtkcc8B8Mq0S1eCFg/
lwlASu2WUBuAj5X1HU3VkI0IP3ZH1QGxSJR50PZ31wwA7oDG6QIgbwZh7ojVDXUC
jpRg+V56i3lXZ3+Ia5AClgQgqVSG72qgAfp+umdPFBbx1LMNhLVJzXAY3h6S3gyW
WIU40XoJb0NvUXFW9Up5sSeueh3oGqvY95egdZA+zIit9zBSHlWhJ3tcSZa79ogX
vKSHxgkrkbPTl7qSR1c0pQ97Xw3lWJVo4IGtuOzjSf5H80pYOoDhJhuaDXAkBJHk
382IKS+muhdqO9S8SoiP/8QCIg5nzH0wdgf9ZNw90XGZ6R7LJHC/CU6zbW0+GNj3
do6W396O+FRYcJiiYYBeyz+ZvQlx8bmOm2ii/GIJZosb5DcYOByQ52CAVtroBPS6
2DoQFz1zHTJQ4Jy+a2YERwhQ43Z79wc1O7sfj5ZVq5wMg1e1UczWPqPnbFr6jj0P
4tar1tZmFrt+fp7/GAE05bCkbI6qN0wUhQtI3e+V1FDxxpGdpfir1kBhWo25dnuM
wF74seIiMSTUkZvkZRtEBA1H7XQoNnrYN+G6gRsImZawj4qra5xVcqQtXnQ+IpRi
a2M36M3q2/ZjcDMvODB+abTYZ8qkvE6W+yZFqrnGV+oXBG1pfCYKOGOI7AM2ABCl
1nEWV+0Cqrk2Tz33tuI/0UBy23cSyFzxCbmOQKeCwBnvtyk4KF97QEmBajO6VNrR
9159IqpkuSvwwtpCSl1aPTkif89LdfnJ5Y+ViiTsY54FHohRX1edCiASuA0CGSMj
7y26k0UC5tXmT/EScpXwpXra0EhBu54XX6tdIL5JeS5mB3jGwYtmfH3yXpqhdpw7
TJrdg15WX0W7l1uU6Pv1heFNzvdjhknWFT0YS41O6S5u8c04RSu4YBl5bc4iP/Tc
FXtG09+f8ECy4qxmtsmq3IjnmHefHtVopHkdLL3UOvncSpcStX6tEaElUyeyoJgw
hafsO0f8lOddHkOptiSAO8Ocpx/ya/MEv6+JI9aG0V4+RjcBlyctIF2mP+DGGqyU
Mx/oBcG/9kurWyXiKhsTjZ80yUt35dYrG5m6+7fqyjY9NmqWERITKk9RlN2uYmgq
+1IiuaddD1XYoG9/Vm7gYdTebi/wwFvbNPqcjDriNzTepZjTI9bYtqjgoeCUqN/u
RXvBCF+gqSulootIDST/fFtJwJJ67R2JnxrMjC2/q/mzTvPxIj1KtmxrLzvO2bZI
50WLDX8Lo34bo964TkiLvwifGj2fLCXPuymjEBIETKrgsYm1uwunW9dySg2bl1vQ
CdvM+x4U+dgG9FML9w5nAblNQFFr4RYAIckgnf9us/IWjYj0ErlqLcWftFGHJ64T
p/sIvSizAtH7lDAe+xCYxo4v4r3S/C9CE+gN7V/tW3r3wqV+68CyB3RAqbuAzL07
wnKdD+WZ06EFFJWKBfzJSMXkme782JAPD7NCZJNl+Xoue0s4qmMRnf6qQimu4sM9
PVQ5ycJnJKVh1hZGWyT2nQiR3WxAu+DSNhGbaQ6H5TZFGcyGftnKCHRMkyKKFhEN
jyPRAKRVD9WtxeiOGnaJUbUcOp0+qs5glgyNwfzplskrfwt+rc8sD/fW0tafITay
YHbjvoxC+lf3mVrvB0eSHlH7NcgbSJV5aOrPmLIuT2zyIlGM000HyHlnsGTCzfLN
28MmEhzGdfD/kXeUINvGiGASmA4dn3C5tS0ELbwmCnSwdCSTs8qSBb393eGTd+pR
i2s8AbVSydV9DzrAjcuUt/HaduBu+H7kG8xIHexe8QLegXXZhB4xCdlvtplAwMes
yPFN8SLORBZpk3wPhdieayluPchZEBnutbnmvYoICpaS153xdZmpKshsIxfbyBel
e/eLG2va2V7JLGzon5K8jgfrrHneOnYc9HiIlxOVVG6vs8Zy/GrwW2a3QS+5IbPs
dTZ3u8mGJiuUpyI3T9Hx37M3ERHGSN/kwfJQ5qkTDD3tgb+/ZlNdyLObvXJ2Jpyb
hcdNo/1TpE+2KL8M35CqV1DZF3QjOh6EGSNetXulT7Pi1aDdeNZtI3iP84F3ySrB
Je0YfNv8k+8XrhcWGvkdDTUkfzKtXW0tJAj/DwTTrzWz9ofIJpxvVqaj38dtpLex
4GjlPJiu8ns658O2lU2f39CDZNRQmlJ2gqDiYzmC+z4outDOjWevP7OYM/arhxzv
V9C0elcTF0h/9N4ONYvvk5VlYdQN3Y9YDZX8hl4RK3tiYIErexQ4qeXFZXo7hlHd
uadLBBVc7cszu0UwP8gf+I70/ClyTpj9aRuv09b7WCH/tFfRoMWzwL8sU/4XW7KH
PR04JDj+zRRG0GhXyh1SS7k/P8DStKUQ3IPEoMJiwl7js/PM8mrfY8QCql5WrWRA
xn7OV0TaSgggOLuMAVMB5qB2BO79xBigXXmdY6no4RZQ6RrC376v1lZqkLZCXO3h
ciLuYppf84ci6UpNxsBUqUMJWiBbl0l18rj77hHeaqplyxQtTQwDEtkK8H/EiLR/
3ipCTi/P2xJz5uRhRFW/SrN/zqRQEGOgcEEJZKrRaiNct/k8+bh9laoOJqZiwbON
hrUzfSp+qAeVVitUr3zZ7IjV/TKqXBL8g1hAP+UYA6xJVA6GmlPa4ar+nW8XOcO7
0is9BBMWM8ZLSC+m+Fgbxjs0kv/OPWQeJrdApcVXX5XqXz4TXVirklo/rL+e+Kfl
MRjXmodhSIdg+vX5h3S/uVSYV23aES73dM3cXai8p6O9p0iJTBb63H+9XPwd/tPF
GbsrR9TW9W0TpOK3OMjVZdrhx9ITmFLd+jJi3PF9I5X477/ClI9LRlkftA2ppNqf
eQMCv0QOSiPee1i0aw6nUASsplTVaUwl5sKiScP02u+C/04IWswrQbgb2EYueWsT
KPb30ECaQgl4+yxxw/ewiiiDvyZCE5gPLMI70bPguUzVh8uDbYUuXi5AVvedJVAC
SxIpy0o/ZKWFcbHQWxmk42C5O6SOyiYaoHgYzOxIlkaYkGRwRBqPaCSZQcRsYFAz
1lj2is03pzQFcZYp/+PpBrBgoegGvHSkPUREVGTn+srvFOd6sLuCEnkcUZ9+XNWJ
CbWw9J+X1uleTgnaDZszs+QD8EIHT20eLH2hfDMn8lFhrPrHPDef0QJ8csFXLIui
xitqSdUW5BhH0eJCFX1g6cYwcJf3DFsG4GdI3A1sa1AknWuQSdMYCAyBa2qc6+mX
4j2u8R1pJboFKGULK7qgMCoHTyhe9ixEw+IJ9RjMhqYI4VDnR33bQ+FKqvBAc6y7
rAtDHip8YmWUCliGwQau0EJ/rCy3GlVrn+hy96lwWPp2KcTZDT/5shc8auxaG2V6
YOlECmoWLZOjduTUOwuZ8JNXCiMEpEAOr3O/LnPNC/LWdazjlsZo/G/4PxDuhAbX
oxvMv2yVInCBpv234wcPUxNEBmGzGtjuaVUsoCQRHooGJEUxnebybkeyNOu+MMt3
ExjCf09GeA0ANOyE72qP5Cs3o6LkLNwqSuC2N3+3n/jyo3Yfl7KCmSvFZfp5feAY
fJUep6TudH8Bl1o4DgO43Hpa1RRAQcxjvp8/GSeVucYpAeYsLXF3ruRtV7hwXXJ5
cMXRiAWpiiuI0vtb4PYXoT8FQjWfdeS/D7lFmaqjeIyQRzmvb0q6Ie1Cak5xSW/v
bb785OLHt/n42d7H+QXSUuYpD38t9ATaX5nWi8cUq66AE2Gcuk2NcvOcA4Uer9OE
sqrEA5tLGTC+nUtb/btQOvHNELbVno7p+6BoYffHSUs1NwsmvqfqiVtSNp+drF2r
ouC2w5yBVG9bkNTGujE46i6dwatkGfFgE+53P1doaEQyZjS4jRH9l0skVoFKMUoE
r0J98hsU3BYOX28jiKL0NhD/tFkRZ32LDAKBYiefY20CXX1KgZ/9X2b6YvIKm7wt
YKpIXnNKJuZu0fZsVTc4iKcBuK44wmBcamuRyUide66ug2Vk5vLmF68dDJvIMwxS
L+2LmUQjF9kDJc3gFrogPYQat3emtomdm6b+KWZzi6xyQpPtBWpRhUZuCVDY5Oki
sooXusnmKVUFrDogmz7bJbgPdpEgXSewGE3EvPlug6ldKfe7l+LaVRvlfHN1wGiT
Ucm+nHMjCCuBRBHEDEYaeo9g2XPKy+VPg+wI/GZ56XSm3kYPK4dTxg69NLM1u/18
j2COC4JwM13PovP9KguiOOmiqVCKEBTrQk6eqIT4QT/yTK+Mi8Hl8vqJ47vy0Zf1
RZN5DgRbsKqpNazoYxgiwnbrj8dnvMxdHmUd2iTtqIu4Y+TzPltmC/2IRLHGAEkT
ZTh08rjFbvMIBoWoYFToFPk45kvIXp2//qTTp0kvfhqTGJCzRuvPlJBelZgAHobH
3M7wmC9at6uJbtAZP7SabRqMlDYW5tr/3eiDJ0gou64qherORMzyRo9nxCwt4RwS
6kxiD+LmI9nOoa08By1jmhilxy0arZ0vFsGYipjhfbtWC40WCGYlm0BmtXTYE98J
9PGcX5P8+5KfNwyRG4p8aiRxjLfOnRNF0mw/zjmmCjRh8HZVpr9Tg8n6lTxndGVR
nQnLmoHUaVsDHzY9PLRk1j+P1vwsyNNTprGq1fZm5lzS80Kczxgm+9hRBavt3DGY
wULNWuCjILxGW+69eJTB2uhvRQDgtiVKUJeE8EwQpktCCdcwWtpsfjsmzpJuIiqY
AfcEsjj2t1zx7Run5/7tZjzvaAyB/BQzQQ55elNEcGIECwtcE540MFgPvfJP4dAx
jY2dVH8R98rzPOyW3pjqaTmO8PjDxHVCi7m3oh5vRdHbpuprTf60weanNklHqxzZ
eKAQVHqE4qzqRnIGZGWC1ai3JwfD/I+XRgjRdM9OgGgS61OOP/Nwjtm2v3IavK5q
Ft8jFp6PoRm/aQtwP+V39XoNxLR3FGaY/Mh9kHLBO3rWv6JrJScnDTxgPcwKNVjc
HHjv77q4+nywmnxYnvxVPtDwVEzws+joqfPwwTTB7XIjRkiESRJePdwmD8o8Hg9F
P62nVXkDItbiOSkUaM46v+zNkNzyslsNzCrlHL0rL3xoGNQRrcksAc6+I2T19/h1
IzIYcfSULt2Ik91zjZNvBef1teZCBkv66TXtjBFuw348bBiQsMtSjkJN5e3e7JIf
iKwFe2KcijkBWfahcOB9JQVfCoaquJxjlxSasscODYBTGS+lFIP4sdeVXNukoO21
yB8qqh9K5EUDePuLPCxa+BPNfqzHoDq2THOBlIa68ZWt4r30slKm1vViY99S85Iq
RYlM3/542edkZAK8PYhhdIOMPc0vQ04BBCC5cf6yhD8ZpRAZWO36ylFrYGfJnx+j
JjtWCjUL7NXxJKedh2QAck4k+88Q2bbb/ecQr+BVx3Get4SrGArUVlwubLGphgDF
ICuXSASIsZFsHVX8waTQN3z4WhhuuLb/kEDNjpnrJf3SaKJah2D9l6dXXk4mvpRu
sGAPfaBQJLLGaSvKQSLJZwjD5FTSI/EoV6tPOKwqqf0Ll3+QXh5A8kpgPxBrcMx9
wihlpGkgjmSuIXet9Evq2NgeuSbNGTMpWd9nHTvaIDBLaixZt8EUZIUEoTdEarzA
WzaLZhRJWk/h4gQLdYQERKE4LrfViXGTQPVAELBJ5PyF0uQum+l87Onhk6kAwIfk
QOfLWnRzNfEojHzarYVmvctcFqu0cvVp+Znu9a30GUZ5PDhBYydfGsnP0v/4FNvi
8xHcAM8um2coyIyuwz1Mr4sHVn+eVXfye3HnGsMVxaZJ8VC4MXyMQIVFEjI4QtRI
cOljtGkZfpEOT6ztD6fkZgqq5EmmaNInOPCOEn7THvm+OgN1Svf1yMMA+uKbt5DK
6ebfXXHNgqCAUpI4IValSqe5mOB1MhPeKVD1jJNzz63+omMm5XhOLALCW/OIlqFc
ZlySjd4owdwiajC8auNdDFN9C3siD89mFxaWo8g752N4/owCuZQC75/6EGYRAoES
/6W840Wvhtrk7DAa2qXlIgzjY2O4NdM3TBdmugVTfzkP4XwiBuEt61cHt+xA/Q84
SkDajZdigKoQ4sH2pdZi3YbPxyWrMyToHfVBvfve3jV7uXl1PTZx+DzzQ2iGUMgY
roLQB66eLgwsUYo4mv7gctGqSgp0H3vVDU5NtC75fdZSV/8AA3kgILtcr4F+gGUV
trmzQoO2RN4cRPTe5D1KZMmQvpS13utXJpAp8N06CfhddGn6uKBw+3ck91OR1kE4
shTIVIL7gl08+aAp6CROV1VPWRRHdxDZiT3ZKQ+nx4pf418BWdIiq2FGoKdvj8vx
MKJ2so0tjqXyBcyTYKS/aWTdoPH4YxL195Dd/bkJn5VUQdMLwTuGQcDjwiKxNmb4
BdwJTGSf2TvEes2ynoOikRMlsbFx9jR2qRMt+iry98dj1Jzc7WXDqfiZN3sb67lX
jXlnWVB9uhTTkTip0b+SKpUnKwBSfg/oh5MUJlMow3wEEkRCPmN8YEoErLLnqaBo
Nv+VdL1LC/YblluLlfmpF+ASxEmddcnnhEpFezdRhUT60Aq07SOzNlrc5YjKU9nH
eVGD+1bb/0hydpHAYGPKbSTcWdxFnBPVodbJR2Smah1wrakwM5DMusYh8+BYL2r3
if9bpeMQTKPor6mV5DnQs3uEOXdRlRLAvk/aW0+kVL6KDziYpHWk3egTeFCvTpy2
IqIZBbgQ0t1yL8YLra7+nUIena7KQn26PG9h8VLyemaJM1O5Ll7EaKXdyDoPvqS4
31S+vUoIK7xLhXoiAoPx3HA8JcaKsTwyuodHFr4/x+5/yYEzO7tPgRuIV5g8bFos
WX36+jAGdpj6A0WauXu526ehK+LZ8WgkbacZPtal0XfYgXz98IwKneSMxYAZPwPB
7cVygS1ROm3U6rmYe1hQ4Oz5JYL6J9w5D/QES7TcuGf6dxWZZLsGpLxLTieJbe0/
+5QtjUCKm5LJpmjwU043/orUJl1FK7RBOR9/fKneLaIa1E0GpoMALAKX43BEfOg8
PUudiiEztWOVXG0GdbSdsNO5F/2K7i5wJxihW+8GotQwpuV71VQoXZXpBnsaR1qa
c7jDUEBTttqIiQPLIb5zBH4ulcnRXg4qoTgfGt462POXaSXvoTH6DfWRLMFyAW2f
r91p7gkTjDSN1L9F+4QXGcSUSmEdfWVElQhJtgsTpEqIy/0yPtfEGbV6p2SUk8Y0
fQt4+S8PfmcDQRvNcfSXt8ozxNX7pF0VXOQNkzRt9ctI6WB47zsFAKCw9VI+hoTb
MND4xC3osHc8DuZOhlUpEZvfDj0E3R1tznUCR4G5LzBlvwdT3uuRdTndDWYZGlum
I2vmQsaipWAW6j5qXKGKsN8+snv98BTc2uWGe2bENSASfGTBGvVBQhfa8tn0qQ5I
zDF9EFKxhe20s3X9dxuyrEvUdRokA1vNut7f83A7PIk6TMZSQufRDmfL83NsTsAf
+owsGROWig21YpmHIks84HGb9WiS5nJ7e/AHgWzElnUAINXQkf/GaUssrnEfQsNG
zyc7+QqCdx9XddrxaBQoOKec9yAUumlOb2KA2vuUB7P96OQt7+5yWmjGfZBkv/hu
xsLjagB/8OX0IswAoUk0qiztdQAJsXhxstSp7HQ5GXUDzJw2dh8dakMJBfnr2VDW
WC5lKKbU5DUaoDAH9/H1TQ2w+3dWJqX6crFMa4ebj6J9ySohypKEuemXwq+ZkTvL
ufCSOevC8pI4/qNhZlP1QvubR1umkA8TmElpeTTMaSH25yqJIm39uXzO9KilaDeP
4qLrg6WRi/B9mOXw2r34/lGe2lhcgqs96MBFuWSeojzmXjkFZFCEjR/DYEZ+ybXL
TpznpA7jx5yty6Z6bqbJGoISgU0bJ/9v6oeSFhSkcj4U19fZUVgkr2/Xk2I73jRK
uP2fHMOSghcP/ph1FfHvquFd01kY2JzJO6cbVP3AeIm+GeWaqBbCj13a0DfyfXkL
DeAMTrLL9wjxTDqB8q8srRPriZA/hYhJsrPl5LUYMhr9wn15ww+l52WhILnDzREx
JY9sJvr+ItcXffh9gKSgm8+IvovCD0xGlns6kUr5uVZ2B5KUh4HOLh5DnGWNsunz
vQJ3zBaWdtTzAHEw6MgA5g7ZoaKFWTpaYgExBZy2H9RlinZtq9o+67nd6ORrdhwA
PftViY1vPKdurZc7XKHTzezcBG8m1py5qePZn8CfumV4480q6RbQYuHDJTq0eizj
aVzDv3PCp2gKCyI243uTk3+nCMaxU0AXQV8YwzayK78eQtoQLz7AslEjbIxy7m/1
e76qR1V1MclJnod08h6Q+7xHuUpH/gfmBvIDgvk25/06Lbx1jxlvFTe5FZaowoZj
P3np4VyOMJziIdQeCkgIOt4+7Jqb8xRGKS5tLN/DZ1ynYh4qohaShNIClA5DyhUQ
BxasdekXTz8F+Tgdx1exZW58O9UTDzWdH8B7K4WJsDPnCtsLiXk7T+KAs6cetc7p
OKpueX8/sB9/ghKY7vtSu6qkGjtXH8DHdH+mUSwZYtU70zdtd6WtTiDJmZjuBNRl
PgWkGm/My61w8Q5GFh+uemxAWz6cJ9mAD2IE+lLhzxd4Cfr5du3DQ1725hdTEVXS
lffLb3tCOBtEUnCgDwmIvoatQqN8gkdvYlJwPvonMGNozXdJj/YoxN5FVJLCd2AF
AkjQcssc56PLkxEJCoKQWtYLqSw/IceJ0mfi3U+N94dUNu8j2blzvw89cderbtaR
VBi5EXtjZDVMt24i9MaODFEOdrHtDoKF2N1t5cMsmhsfTjlrKE7osXrt+mMjYpzc
PVzU0Vz1UF8gqrVkAuSLEd5nePa6NP4iwHzNT8DVN1FWPL8pVwuVAd6vZggYXECA
5s5gplz3PQi6I5QbsejqUeO/q8wnBq/W35JwPRhwC7Ce9G3l5OiQ4WCqoUPY8L0/
djppJ65S2Z/0bxc7MX65rVYyIy3nVSDq5KUZkrjn5jnG25TMNKBqP45zvqcY3DfR
L2nxtqKDx1UxuMwTZjEtnqgSeMQDnPwkzVMprf/3GXamGW7sPf923WjJse1asZZW
Ay+8ZBsyRFTBkn97kq1i8ppO+3emPSy2kJ/o101y5B/boR4GXAoum/1dOgf8ss70
vH6jMQKZLNpTjIe2EE/bhQ9SYO/NeubDATzXFpCW/31DJt+IjsLD6fkvdWklpg1m
CvrGoRerYYo7uVB270+ChnCzNzXBEZp3SSvpq78zVFFUPg7QrzF/mBn22k0sdcSS
AKacY0mJMLMA17XIdc62EZo8TQWxR7FCmkc6UQUIxX/6JtWKJyDUgNA+pymZzGT1
wDqafbcyCi9yitt2EgXbIPIeCREKedcIvY7XTaXdDg/rhq8dJVay1bH8eFGhJLPJ
1PKhWymlcQ48+NlkydtUoFWBLsHPu1TffFhh1zD10UkEXpOHNh1D7jfx9fj0XJp4
0qeIZblPAjEwPaPZNLYTo/AYSCG2dsE2gng7krpCv/jDZHD0/c0+uZimsXFzra16
RQcCSB1qWz/Truwpse2ALEFU6XXDmzlMsBBFwQguVluvZG+wKlLshRwIF5P0YOHm
KwSl/KHGNN7bd7UDX1xxriwq4CVjQUE34hYGiYzdrdahWQIGuVpUvDQ97ooOL1d9
m+sNt5QAF5r0XhTJ0hc8BR9T9Qw7eWsxXFuXxgYfdsatXzyyk//otDcjvuzHonpi
5FJa/Bkhx8jF6clq9ytIk6ZP13O9YIweR7OhvDyDsZjnYLJ+woPN3tXC6FDJBhEN
FuleI1ILDqIziz5z8SvhPT+1DwoN85tQNqaQre8O9U4NB0t83/ZZjIMEhCt1ATmT
aukw9+8UmsvP9PY0H+TdFprr7UNysMYUA08kuoZ1AKGXO+QgigHLoYmnuOxRBY18
0liQX2Azk/COcRaiaI7ukUDmOTJY7PTdC9LIFv4y3kiBt1B1IvzC88hI8/qygf6w
jjTodoLnU4FK3loPlHH18bDGW1M2VryMwkopeaz/c9qoC4dxWnai177/lF9nDZTu
X7fW3w0bBzia2PRYSE7SO9gPOAnAA/zERoK3dGEtetIc99nvFebf7zrez3Md28PP
B3x81kpFRsTXZ1Algu/zdmpIWVaTnbNYZVlXZ0aC+CFrPhXWSN2Ulyi18dhxwf6H
cqL2jL5GvLH/h03YsmSE3iy0KwI438FLUBDHaA2KbN9U96YBf4fjqsgbJn7h3PDN
oafqGyzl5m/OT44EVGfPcNP/MQuxbw0D4Q/4VBFCXuK/oqykk5jlrGCwlSFBxafN
nbFKzizgfQZBfYhhdIcs4/dpytMolJE26jmNzmtzb3t150a4jiEPuVBgiJL5UDuX
l+MeN5WAAADY4Qd4uPVY6FMf2bsVVGVh8Ly3k7F0Wzg5XPu97jtuziECbhQc65I0
Rs3c17tNq3zDFcJSC4J2klIoLb35qqG6f1El71xPEvinQqXPTOjT4RJJts2L+49n
cByrGOpuX9cHGsKgaB235RBv+5uvDgQdZvXEce3zofwuN1+H6bUXORZ11fqjbmyE
Us1tNeETTDvVZ87wKoCP1ET2HYCbouUSfkHVCQ3paVc/FJcDnKi8yyrm5Jj4pOR0
zMDu9wJftDqvhtiQPuZG5afMO87lNWLv4SY+96Kfy/RUAnKIreYrLGgiSfd1vEZR
perbbt/sbaS4RRNwBhqREEh9INmd9h8V5IWi1xLBmhkeCO9yuyEr28NdCWxPoy7n
vIiuafbl7DkL13t+vZI+/jIH4mXMx4G10awh48cZZwRbSYsPnPejls8nNOe+8u1W
DucUusJaPzL2ffqwPD9yITWMtEcgrnQLNJDFxwG/1Fr4Ai6XAR+02qij475w/phx
GoSRJUSNBQTsFwiBIoYhdmp8+FQysM2jh4bt5qwJaCC8Je+8W3m1N7I660foOLsk
cA3EBs4jg/mweO5aSIIulDs6cYNDBXGe98WfnCZK7hNZG3AkdrqfI+nlgWpa+lKq
dVIEwU2Vi/q+/u42IlDOJmw03qLl5ZjjXLkfaE5PKdf5Jo6na6xXa7s3eYjWphBs
iPwOi4GlX4Rv0p1zKySGpnK51xqc7jqoIg3RyftfwMEfa2m8o0UmoyXKNhXAgBrO
pY4lKiyG5yLKRT0dzubTqwutU1ONAaN3goiQ9ssZioNYpsPBKZIpU6ADFrb/iFaz
W5Tre8ZLzd0Rf90MJEfOKVKD3lXJdMDLqHZMjNJ416amY1SKBGdNsPFjx3TwwBlO
BkBQaAR14afEiC1qKa2QvUQ7MkmsZx0M3tY1pllBItxdnGWNnnPjIVxhRnaPy7In
tn0z+UkBkZjfzqVlLchHuRyu/brxzCzICIqUwxiCehcALLCM6B7RnF41FKEPtlPj
xx9pSFYylh9cGGH0m7bblmoHILAJX51CH7yH4E2+STHqpp5v2RmWa++hDYOKR1V7
zFUvKY3/jrKaZraniIjhsGhEw9ijwASfjQ7M8FhUE1/u/2fGfuzlKXqjU1y+ek2p
PvrvCpBluFTH617fNbS6XYY+/3gVFhr2uVm8lFWWKKafRBrA8Ry5js9HfVop623U
RSTBzFoNbdFzo3VcT0DRVFzB0ss4DKRnQJP2dkzGk2DvxSa46vikYXWmyxeTnM4l
hIGsTeLE/SbqljoLKvg8y3rLkM9p343w2XMeDe8H2dTFoUysqE0PklQWrprivmqj
t0T/d4CBYX30NNjOuXGGPJCy7nk8xOq2oe8TNfOu6OWgrNLGYvwvtHq+klKEcsUz
ZHMC9m7Bo6Vh4WeS782HxPqlRbdto/XcnobQ85RtRbZ+VnY2hyzNHg/BEtLILC0P
BMFsXfZ792B4vpQkUm+nVXz4etJuFKfqEuN/lkPnRBzNhBC5qTogV1LSY4pvaHGr
fE4ZfBPhyuasIPsz4HsvoPvnHPTI/INxhAfrFp92qh8gwxEpO1EiWnuNPtgZ3DXj
Eia4Oi4ss/jo3txyuGmIbK4uO7jxCMbxevDH4DQ0x2XFrdu+Zrz5OnOJVNPsxOS3
R5s28qd33BDy9nxdEbaZbCS3YaPBSuGE4kvLZjGI9EJrnL4WmJkLKYga4eQm4qLE
Wh1aMYSQ3tnfsm0DKYVRYnkE3xQ602teLl6NeMdKJ5PiVcoWLZwcHmtVZqVqZJ15
UjPFtCQ/p86cPZ+owqP81JACqeXYZyPqdGP12UZwe004E02hy6J2iJcwD8x35wbY
l4NAHY6AFyHHSCiFZp0DnPJSzMB/YThGwmYQb3tMQfNgm9Q846CB7eFz+DRSKE+Z
bMS5PbwEB2IiI8wC4H69AM2r4Gluawblqve1OwWr/668A+5e5HdrJwC2WdDCAjLJ
WFEMkvlLlo7yglKED7CXwqnwuWKPb3TI21NOODkhAlsUmtf2xXw6a0/wKIBw2sTU
RmdR+lL8uNX3g/gI4K+JOr0xpifx9Oor0KIoHw7qMF5hMNUu2mX6yQ0SRvMyjhyy
u6QgJucwpq+Ut48atsV5xQxL/qDmoHLLmPMgxfyxuQJCvyxtC3wjCrMhaNYGDXqz
aY3ExnOFH1mqEvmJHSP6AEqTXI1B+oCkmZJ1IShIDspcKnDCrVZMNTT5a5euErA9
dMyN3GWHH6RUrHsvPvHh648tyMT7ZzMO1nxT4bl8WmWKehDaSdT+PPPRrAzBJB9H
XZ83Jofd8enP36c4TEOe9GP/cXeS4XGiDwVFF7qdz6o2QC7FFwj9HQ3yd8hhbkw5
ACM9sKXR3tt2Fv9iI102vqJSDy84TyOL4akTqanbG+sD0KRZdP+yrvqbMPLBaoIm
D/BL+3nE25yxqX8nI7IRU+IOlOEZ1+9Iv/mFcepf4BAbGnjdpu7ApyGt1nTdAB7o
Ro8oNO6lnQwtOrxleWT0LWD3ExnYrANPBi6AJgZ4IScF1qZ66EEapFqjyc6jUqi8
/JP0we0Sm++Wuu4idATeY9zQJokI0JuLpNe3Png3Q4XvlbGdyE/Gr8o0H16fCNSJ
PP5r5ddFInnZ1sFYE4afmXFzWAC1znEo9yN2rvjY9e/9ULps8HG6vYhODk7EBogQ
zKfMTjT3UYoFo3g4W5bZAzuhpGY2I+7pDkTQf1M4geV86j4xFs7soQCFCNLdca0A
P8IlNz3DLfMSZs32AjdQaa/CQPV49E2/y9PDg5dddxX0LbDwCoc2+ZCqkGtk53HK
4bda5RjQAzY8CG4Y/CWWQwE9mhpqrdP2JxgJu+HHYbruLMi+ldQ1G7zu6RVb+KE2
3pzTgOXQQK6XZScpmOGwPPtBUT++9IyhsP3NVdwDPyMdWP7kN9/LEuCLMOrGICOI
RZM0/iW2IEabcTXRqYUsnB7y9RHoP8MEFXBb6dmThAXX2kqa5Mao6A2i0VHeZVov
/ak+dJEMkCCn3iBP+OtW2ZT2mosyY16G57hpeJsofFaIBPYspn+Q7mox3+q2A0Ls
TwQC6juOpdYEC3wTPwDnMfrX1TuajpjC9zTaPM5vj1yW305TQvUfOr2yigUnPoNG
ctRVx1QNhI0MqEQft5jZKlsZtPfVRZroHaEY5Cg62w5MJpYqesXgribXzYYRQDlw
Itz+7V4uSfGcit/NufYpGYspXK0He0s+TVasv8kO5EE9RgVtVNuFmBmKOk+JXO36
CeQviWcDAZN3z1ScwxFk5R0L8tvW2DC1cBaQmCE6n0bFjR60xByW6/DSD36Gmegg
AzLL3S1cxtCX7A1LeuyLJeiHbC0s8DoBZ3gQ980X0qVASWX3fzYirh+fVrmAwaC1
V57WDQ6vrLS59d+pG98sn+n43F5stKXX2C1h23HK5PnEqT0X5iXqNcokyKp9OBT0
CS0cGajRFfy6QGgb2MLhpfeP/PHUOVKe0O7Fylt6OZojqMRi5LoO5ruppHjl4PU8
Pdhb8cAYUky+0C+r/GXon5GZz68PqV5GqBwfEHb9jgGGl1A1Vom3DjAXlzxJM/G3
4F6ir2SG3ZdTvbOfz6vlCfEG8YR4c9K+CMo/fCumQKX+CfvCjgB1IM07bZ1q94SC
eU1ezhlUqO83d0Sgo2dg2GmnaPoZ6XPhXsdj4koQRELXH/iQ/HkIo3x34kPvXC+r
+8IgvJlvqkm09JdQGXh/G4AL+zw4sVrk8yIOjTAezIbFeGm5yiyVN8R96qwSmyXO
Bl4tOykT/FHzYXtdt4IqXZzbuxuqgaCuA7xp1nkQHD/euikmZsFRdNOA0tGDp8Ng
MvJk7HvthFwI0qZ96tRJy61zoFv1sJaJbR95UpYr1p+HQ3kD6buXBrLYq5+tCqdF
17+tAJ1FD1uco/F1AX9AJmDvufjT+Iz/4zWBi75DSvIUotzrH6bKpX1whU+G4+lO
4eOD9AAIuwSMIgZSs01GuOKmFu0jEqga1lex51WnYeFoslMsQsg74lap+D5weYCX
GsE0QMUlSTT4FfKFL3NNNh8mzTbAdr6QSxyKK0SU+sHG+4RTEwY4LfBWXTCnJQrY
zDkW6eC//Qx2kd4U00aw22wwMZkTIECwDbMky9KE5itZQ+CDTPl8CwX6wDpw0Fik
cutU0O8gqevL7VHxP+8OEeTHSSLbU6jsSL5AgSXukxBYL8IPqEDlQLwplYIW3d/3
98DitIw+sqlk39mPKOI8zNLBCSttOIuid+LIyeW9cffCgS9+mL5/iuAbdxowT00F
VeTevQmpCXdIz5Omaco7iiBsW3dAUKHM36aXXu1Xq0cb5BtQ1kgl8R1Jwtl7kma7
Gq5BxnWWKGJ3qxHA+N1VozlSv5NzgSlrpNpddasbvbh7SVeJbX4OCRryXZ63y3WW
DFcuWByhhbImPH7WJblKFDikcQmYWHus9xiLSgPGtcSbnDXUh63y8WOA7W8x1EzD
+x5FAPKqyYi/ogC29z4KL+mGJqNf+k9f6K7J/uzSSuV1tLkZw5pKBCjpIYh3beUC
wyPYLMwUwbAzSG1J4dOMjMosR/DwM1JUmD+O3H9ZGidKhiPh1zQ3/4WucYhTL+sq
VGZXJwZotO9/l9kf1/32czIGgJdXHe+/AtUGzEYzthMxSsavWEFMg6W4DkoTGzET
JS6c3NUbC8LKdtIwH2jOT8amFWF+A5Hv0P+tzcXKR5ZwqeaQnXwoowphHYxl60H6
ZM5ObQbV94l5SC3RLihxDCIhVNBPwHqaXPC8DzOQftO/qx6VMGXFJlAWV6cogoXZ
WaJmzWM0coUYQ0gKlezNTfLPbPaLLO+SSV3CSm4FWGJQUBg5JME0bVeQQVKJeGnX
NI9GHbnzUTGrvZN5jxVtQ5+3yPhf77bCMpSCfiGVTCNdMslANWNMZFeTQmLiYrY7
S/TLav4RXHWxxXwzHb5efg6SeZnC3o8P1T3W7v8oQtNBTkyG/D3eNIWF8Uv0cJ6y
B7inyL/nEnAGxFop2NAQn8p2iA3ZViV3mVHlpVwu3DsUe61btVSR1H9qVL4l5mnh
qMF/8hmGUtXXskBBZ0L2rDnKpYlPOouqvEb6xf0fWTy7NKqi3QxLa2sRS9YneDCV
lY/rFaTEhasMLX/6+p99NNKtQiBulFUU6nHlkUwV8HZsBkc3Kihz4TOK7Tf2HeYX
F5lWMaHBP3glp1egJ3406DhGsG3Gi6pH19WrSlN1pgFTdlejTwlzxsmZQk8qz5xm
LC56HaJ/wImh9+Ub6DIS5BukM7afkuXn4F1O61/BUXRM4GhX0QsWMoPfd45PCJxV
nHkZ2UnJec3+a3G8N3i3SRU30e05EhzehIde/fbWUmXrSOZzHC73S1sdLK6TIG4q
BLhrjqmaYYEywjgHyc2pYVEnS/kA5Uo1w0x/TfWGycXPK06+On6KiGxsYIshVnD1
FdjvNJI12bLu8xbNuMHZHaSGGXuGS2nd8A5Us+gTK3cLjIS8VwjvhPru59vC+u3O
C4twYlp0xzUaDNTdRSN3U9AqB50CGuy5lberUw6op1ysboQ5IDsaU5AGuyGJa7uU
2wMXYssaBchwWgS55OXxys9PvjSGBbK3TTujFYp37JUok537A6tW1mAcIzCM2G8u
t3P5aDvJssKvFpAEwgE8QGl9lKShAvN43j7gtdra9R2omIJ6dL4RxsEty9T8kUXN
ucCsIL0lOh/vApdjnJNL6X1nvHVKURybAOngQBTKVqC7VKJyW+fQcznFqmY0+9XO
gnnWE/DHxEEgfjn66jk6MxUw1KoFHfHYx99y8b7SngvuSgrQsYaLTLQZflnbpol4
ZtaW+pfgtFiTjXWQSnhffnvPrJ8zkINmCDEOeBFnoiWtIXgjEKXmmLliT2WjuchL
k+OHVL0Em3Yu/BVy+BrkAoa7RqV/o0jwmhtIBfqQcOrniOmv16eyGPUYfHysUEvk
u7Pkw/NVjNumJ1ZOyyeZhxceWNHqpT6fL8quKoFOn5Nw9PuxP76p6q8IOb1Um9Tb
lf14YxKZZTEh9ulJ1I2Hz3XtKNkmKHXX96LeX5BScb4xRGUrb4tFRzDzsqDHJhU6
/WCHV8uJ87+Byf/DgV5dUb57SoJSQKMQLaYzmI6kcZaZlf+NuD6NKE8cPYundYnK
UAUL7jG8yYg40i9kvmLapCob7DNuj0LoQeILSsd4EO3E45/HQ/29sI1tPkCT4PN2
Y5Le3zlqSWSX6nwWcLDSWBfs+gz+d8VDajXcSDcbIeMSX7sq45j2rRiZb5z/YhF7
C0RuJ33Yk2RawieB43JvU6f37L3zI3eROlIGoFqevWSLOw7bUEDuecBnzf6KDC6U
V+BFblRrcpM0YaBJpzbMrubjdD/Mh+S9zwAIKt9LFnvkFR/yQT/3tsUtUGi2tmak
/fYU6i9ZXyJorM/xYj23GthDcV3Bmr2GCOjXZuqK5IJwKnLH7o0miH6t8BaN1B3X
GZLEO0jNCdAlLa8okuogY8e3QvbKt/Q1y+zVXdlEAWtf8REsAJTcM1VBxxhJYKi5
6uN3Ol8CuVOo9LbPY//YAC643zjyWmtnNxiZfivGDA6cDraA0uPzM9dJBw1IWJbH
zxqoyKgsgqlsJtC2zfsHjeDr5bVoh9zINlWlRtJRTFx+PAWxRpyv9tLC3ozBMReo
GTpRjR/6H78+hEkKZU2f24IbiaLU/ITOZYmC1nhKmh/+iwKdbPIiYy5X52U+Mz5R
JRl/MvonwfH3hxz1eSv3FZ2GNm4R1fRNDfkvQoWch0K2Ig6LIzi4yiZKZp2bIbg6
Cx2A3BdkI85jAhnWFxovBTKjTPaOy2fh12elBzua0EK0G/gmX2Io2IJb9mxaPshC
41aW1SoOnKkBEohleB/C2LsN9ljM8Pygr3ZcL7xKqNqV4e89gpmOj9MauvLQls8z
J6NS9MmSpdLIEeSUmxknFtw3LmNhvjKnA/GtLdSgLATxhb3C1BWXUewYSd8e8HDp
9JJ31fZYAVHvsDOCPOFsNKd6dXtII4pL3BOsMCHCUGhulc+hnpwcqfMk11v0scn3
vSA/Yso/O8ufv7XghabTw2nBT25CzNWyW7xNagAcv/7wA21RdbCfxwBuMT802FCR
OWbqk3Y1iPzwNayJyxnMOxz/2VK3edjS/vsSYp0oSpAqRXBbbEGdCPa5tJnYViSP
KMIYHD/MCYD+P2tiyz5ZX4Tb58PaJsNC1yTlhkeVal1OieaxxFo9UuQGudJJqczs
1hQM3uZMRpm6QhaFr93tB40wLppmlm8YKqGtUjodtJU3E+nZ2DK8lvHsK+6CmeZK
AFx7Th6xiRCm/BBEgFMHH0BMxkA2Yk6CEqfnwhn/YwhX6FOtvMHLSZ04nZvRmQGp
ORsAbJyeWgw5goJHaLh72Z6ifz9iKyURcNVpnr5gKdfubk9drydsO3RWwm4WWcWf
Sm7lakXGtB846p1b11ax80E8rWVQR0a0u2Fgk2PVTu79YTa+nGyf7pAmtzM46W+x
nK+j83Wps7ypMKx4j2QmmaqBLgQqHMqKVBLLy+qw4lbuhfLyitIOnP3HbNljyr42
CjhSzXTRZTooCuPKFmDzsMTbxJoMkxt4qewvPkegcBXAlkF/7G2+rOdZq0QC/fih
D5fzGci5v3Gi8OcA8QK1uQvJkLEqfu7Q7Rwy9YSPO4FVhWhWHwMOc8K2DfjCmpMU
fdUTdXUyMn73wlEwXNF+iWt+zWYgDOid7Rnh2oNphdcZLo1ehQeMtRFBjJ+vZliS
uL8nOIRo4LU+4eLR5g5AgTIr4NsHng+kDOvj44cFoFiGuFy1xpA0XHuSeyFuYBoF
3wfsO/bCrus5TXZr6Q1LFbOBxcFAxmzQwILIwvFQPDQyuek+sKGrgTLPrLngIL8o
1B3C4GYpzw652zGR88QS/4/qPuq7avO6L2W7iTrQ0SfZTkZ6qwqn2gJoZoTQsCnQ
z9DWGh0jtfCvZIJhLDKhqxh8Q1dJ/dycbMgJQBpZgaT6VABiblRQQM5QiLvj+NJi
JYr1+xu5BoQ3ux1WJ9mQAkLvfa+/Vuy0xmntpd5B3M4mUddFh5YExEm/wVLgF4lI
R8+wsXi8UcexQEg2qSNBBogRbZJ7wzlfF6g1jF+0+40cLH68x1Rx9A9UqccATCj5
df8NIBE5sJkhgd/15B1VH/H0oD1bH0qDMgEpqNm60Gz+mFpyDl5U2CosPzhsPoNz
FHc4frgoNvVqGAVo36w4Fe2H/JFv/VPWy5jNrA6zBJ1tZsfCN/bAmi+0B2S5NlmP
lsz3m2ZOjqkqfoA7YP8nVswhvpQoUQ+32qIqgu7shVWJuim4txDJ45ITD08RueSw
43Vqm0s1kqgJRKz0qyL4p5iFgy7phAS25RhSIERq7ripiNUx7yTBcGD8WT6Mw3gE
CyvruHUU4RYtH6lmraHaC4LdOO2B2sMVXwo5CZcJIBfzHPbWfpQRQnN5XhB3GZMA
fnqU1+iQSjZsrdO8SxO+pwpa5gqwmsrXuEWd0PjxutQda1AvxOhj4k6QTZFNoCwq
yz89F2lh+SzNwvT9NYYj0C/wcL3EAeOuupPnJqatlKJhllW6GjIGN0+hVTDsDyYR
ENXBd5FNqSy8msxI/HFIn4DucEkypSYtInpvAawLhno1tFrM2452fRxDfa1ChH4Z
1rEZlnPkvj/s0iM8BQTMAF5HqcEDiSq2Dq2Ykkm6zEMRS6XTYnIYN9pYHAwJ6/UY
9TbY21YCHurOsOMII8gvidNEGFok5aqJ2aq0lyF1scVQBDfJfbhAens0qL5juqwV
Wb58MT4aRKb+ugswmunrheIAGtU31trFeze5WhgYGFF6tWPyrDvXxDmnpoZ9/q2I
TVc4YBBougUUuFMW7JUGisKqlTSLrgSDnBtJpPFKuCz0AzTtJAoTPprdmwXMbS+U
A+8yj+CjDq17lPXaML1Kx7zlwIWm3i48i7t+P0OV3hCWPOmd1EXgaqTdjDd9O5r1
vLll2EslJs17MsXNt9UJHPRSB0jwFQ/u/6F5UxJ1P9j+/jaASM4OnQ5dZ4xcEnfB
7wp0doyVKPTDBxXTe2URlBr8Hsn+I/gmGCDgJ/S07EHzPgaU8y4EqZugB8sCabI8
oPM3mpmoQxUthAMeZN7Si6cHit31taz+MuvKhhMBskwFWr6D/hjNZcvZjsll/4Od
4cXLszpnAyZOD3+J6I/y+kubxV/H0JY22eIITFE+ITrWGS3/4NUs9DPagEgt0DOl
VB6NyGAG1V/qisHmTfl/uF3LB9vOHrQdF96lH863HIQ3UmqZ+PM8b5H6khtXGciT
iQIGbN6R3aG06X2YCkNZFJl9cTC4qWlT2hx4aWpWDMgUtHqLUr21b1pbzmtEZH+D
dyhMXb+Isvl6pWSotNdCnJ4RcZbuPNVeLl5GgKQk5wkjW3W/yRccEytl0yyoK41H
hPCmrWAS5tsLm8+ghAgansesew3qSGco2HSDCYUbGsA3gMJ4hX1TlwScJW5SeVic
EwsEq9/5cegU3p6JahaEFGmfuEl9lhgUgz88yHuQHjwksXwSaVul0Zj8H/+6kbwY
r8gPv//5VqYOt8YYIOlZvMaa3GxCfe0oFtGMObtpzgjdXTRIxFX8frAWk3oIMLS2
E/ObQebVUKIUdBYY1tn3zYbcu+XlwamhAHRCo8D88AQkFHCwLozHOMdEl+521RKY
KWg+jidpc5c/GLXzzh+pc6GqC9by4ADSR7TlQYVh0BitGWVy8hmaPYpMMxjmPtyi
B1wUz82TMHJvFnxNxAkV6EUo+Bu2wfoV+u7uWrmKKj5gC94D/YDiNwzUqrpLexxw
HYkieKcTFwPxEbGQ+8SfGATw4ZtuuZIqW//ZnsqNnY2ZuVye60w/9ELW6NfD3Y/8
8DUsHK3rMr2eq0yxSyPd8rseeFk9cp9335U+bH96FRHp1mb3BowMew+PdNi2cwld
j8H0jTKAanzMtgCuYPoERkl06obD5QuxfL7r/glTVMUNUCRsAA4BhDpojetl9zz5
ksTidJgFISFY0zPPQGjFKYq6FpePm/wrmKKYNYvdns8BENGJdAJ21VV0GZHl9fqy
yA/DyUWvMehpegiUeVP8WAxlk14MownwKx4jeK+MJM6BPaHXm6Uq2GtTMnki/74x
ni4NKrn2Dmcjxglp1ehzhAFbRxUwUIOseejmceFVm8bFHjuwjPdeVIqFam8kICTU
NixV/9Yb9Rp51TArkLlaKzsOORZ1Rd+st5QgZ9kc89fIsFwo2FGCQMpfZepbk5YX
X+jfsfDgT70Of3E3baM+otrwKLGChIujDMvqObyg6wnNqaOUZjxHwAX5sGxz2jK0
je4Bs5RA1IH/iN0e0K+V/ByfR0CNKYxqmX0+vB2LPyRf2hpXmqdNRZOy1xUj7eor
8GnWJtSUTW00nvW70lTt+t7hSGYC4uehtzmHBc0OTxgpIM4xybmFA/g+lYowzpIy
jWcvw/03qMciN6HmKacCtCciSdWnipoGEwIh8OFsqeBtLnlICTeZjGigFFP3TxE/
EdWTElYhj3zrJ0zexGSm34nYoj+fpsjYhOHWdh0utxgYIgyn8H1YROuPLenB8gzt
O0y4GgpEADQVn+kHtnic2TlIr6OPX7b0KT3+YVIfJh+MP+HAzej4b8blCziA6CtI
3z0fFv6zA3jcV8bNMOx8YmGdnBHycd3yB5MM/SJ8a7mWqTJ0VH1KhNEyqWXYt9Pn
e95Bjm+3cBX/qdPeV0l4ayIBRihY0WwGOrY0wfIBAz4YDkwTs1r+XDqv1kVkMQut
xrBqwe5YL8neun73VgHGgZrD9aCjUFqdbC4onTtMIzTlaE/KRz5FEf7tODsQKVbS
dGRHQw6WFAUQwf+yjhRavt4RY969LhmeTX2Me5gVkhqkClvRXqKDRRIGy2ThJUfi
O1enL4Q1iYr5nl8B01+75sW11QX2z079/ZljRZTze9vBV9ct/uIGwMELWx1nePpY
vrPZJxFv+Y01uIef5bopEamJ1uy/x7scsk/ZcJI5Jg7nyHOObXW2xibreB5Djkty
Ugw6GKtmLRfC8HU2DmmZbZf/ViA5s+NTu0Pv6dVXaNMOhkcxiiKbEJDgHAbZMAzs
3enAwzjvSufXZoH3gQE+XNI5KwhynDZlF7TnTYFridu69oSqc4+l0cWn7BlBX9/1
JiZrgebwoMJBLIUhc+y8z3NcsrCw3cPnKnbmcPPVN+Ib7YF7M1r7jkw7knvVNTo8
54ymQ3fFsBus3C0Y6rwirn1yrp00PqivhQ5WLd+IzwDuJqwWVbbOq76BPuhbw2Hi
cfCXttN8wCPDrelpJKjrdOZ1Xi+3KG4sJdx+I8kTsiOOyYtizbm3rIJlCxuEj34U
p4+7EM/LBkrOjhaI4pDpBfPZDH34hpim82E66lpUmOaawQn2kvlYdNiTMObprpIb
Bw+pt4ImQ70pEK/EX0Njc0/2OU3ZlI1aYJY198y+yS2x1SvQfYjORW7blrHP7vac
P5Dz3Qb4q8V3Aln5y8Ualk9cecxKI6xf/NQbADM7lDegr3s9LbZazd9qjw2f0ajK
l3obZ7GmK47xpHla/iqEG5wfcxifDq92XC4Dc33XzCqiPBuCUMFfI4QbWNSx9dAi
i4uHEeWXwsaL6rDBnYcj57nIX085+Tl1VqTT6YNN7tG50rDzV1CswZzNMMXjXwI1
0kyPwiLvTUHaFGRcvsoj4i8RBP9zbaYLX1emhJWzxaBdj7awTckJULXXPX0qzNvL
wkPPwwGpgWx1OtXWBassdQtoOLUNEE9wtlUhcWHX/BeeuWLOg6UnlRb6Q7dTyeU1
H4QUhmCRTYOkmtIiiZ9WsURnve25Rim4lE1iAaEpPx3lCOecmpOBWf+Z81zUZ8P+
ajYaDTuAaGJGCLd5Q8+C0xiyJPMX12P5nzEdWPggFDB/Mbz4fmIhXv7BPmVW+Xy2
H+L0ihJHKgJR4nrIfa7nkQLQmkypSGlRrtH+kIzRW2BghwbGo6gWhbvMzq7Rrv8E
BaIkqet2tiU2G2J8vX83LcvoOJzhp+0/TKCptNAYtbXSiTul2fv7onJknXA52h6a
ySbhhsREFjMJmdXeBs/e8B9sKJsDOmckVXKha+A7VH5FFnlHHruQPlaZUeWUi/AW
qHOtaoc5M+aGcz1bh2IaIn7U4wotqkmBqJfZUlTFYns1zVVMXw9ToHWBedYsAd3z
zdZExycf1vqu7peTbPcdnL2DUH4oV+h/gc5u/q8QUb+InQNAZdabZ05ySbPSqIeR
Xhr0QzjO8VUIm5CvRkbcyBmyvzgyp9iOdAtJsGMMDXscB1PkhPxBnTKPRcejQvwk
bArklP771RDVPJJvWzXNRwPIouMaLjbxlV7VIwNuv/dyJdXBedaHcqAd0yH8MtSU
mnfqmcj6sbUvVigVZZ7oc6OGYWmGwYF+y4/biRSuYqUex35AVkW0Wem1CkcgB0NA
bdqSkSoabFONhnQTE7GoPmQ+GkCk7KpCmxDyqLadgj55DidUTpC/Hr33kHf4D969
6BChKmrYrEytHGYInYNlRUG1uCAA7rM+Byxaw+ZikAphGAuwUHglf8wcXSKzpIXO
AlhMiHzVOjy2pcHBLP+6rFvOJfXAQWvRzQjkw6ae+Wc47wzAuIRMxxUU5fnnaJ37
2Ia8stgWv4YXP6vTsXNQQzpHAENVtM281x8M7bUl1pSzm7vqpLXdgJjSJ+RZIYS5
eujwU0HLn/FJFoFT3ziDxSr/XzYFz+ixW7kZDqi4HSbKNwWRbb4+cNcUUUCnrwaF
Lc5N35ZiGNxDFbYUlnoJavRip1+UKUEAdMizrB4rq0ZsOqlxaVGM3ZrUpDbf0bcp
BEpkB/+O1jOQRj6wRQKc1+VVqpX6RU/T9mQCjopAsy4sdo1IABbvzq+vnLwfJHsV
GCMGdCBx88tULmFs8miPzg7RsnMm89qg6iRQ5XiknBYIT3S7hxa59LKMIiaKv+Ip
e+pv/u9K3MZrck3Jc5Px4nvrhEq+dpq4cV7BGhVEDETN/c/de3Gm8KMPbOLOm+s7
pUtdCpskDBlhf9ukRSjaZyPgErMA1Z5+0ZlNB+jlxAFDZf3y+47oVrR7WrmuV7Ok
BlowWWpdhyzy5h7XaHvgeemyoDJi95G/ToJz9GaejgP0Hz1wdEWc5SaoqD5M5fmt
lSKGzn1fanYSqj6dggS78Bk2SIyRUKsZ3wKRxncdtuFHAIYoljLnnazOBpTGzGku
lIwr7mwfzJQzv9j8ZxqAvDQgTCa0Mwbojw/ZuWhis3wtX1l41jre8Sa48c/PFrM9
DIjvqIYo9Pudp+AJChvaCDrOpHWYcuXdQqKi0rDTsNOBCVq+jWGnRr3uz1vad9ik
cVqSR1bQeKeD0EUlQ3KyrPur6b0PHp3kS0cgQaSwkUJo/k2y39yT4VdYn2uRwpQO
tIQZAp/OhgTKYE/vTSN1+uUTy6A8JgPs5Sou/siKSbtPXVsyryCAI3RZt7UC/tqk
l++LSQuuWnTd89RaZyPMCTR3EDFBUu2GdNgCJHx2mVzvNjxBBOriokfuu5wcdlfP
nduZ7KyGpeukqWvc4n8XjKujEmCwde3/hQbudXlPO+1R1Jf1mnt1Vbx9J2VDbwQk
nWZTbeFDatzCCXcF48ns596jm645AqPY3LfR8S8iscAdiLLHKUhGsvSlYH+pYEqK
TfLAXgE8O9871PwHyqlCNW1v8eO+IOW5yyy+pW2W2mVcNol/vqIu1uc3W/LabQVr
hAsssFrfj89jxsz8OhpSjSWg+YFMYGMDWM8cHGaC3c4KQUbL9GEPGyKs0U5Y9ybW
1npWZ1sGRXhN5O/Psn3nbAKuUxlrMiLEQX79CtqPT0YHplY1bZPcz99LGT3ldali
CW2tToxArCLSD5gUa8suHAkSy5TXxuUeiYz3kkbSCOssNH3qtXXwlftH+eUKOeR8
dUUVRzKccx067Tk3+67UxlPa5B6Bbpzi3jSYkAFtG15SuyktuuG6Yfv1MCVup6//
jp7DCa1TqW2tt2QaygGPxpT4W5xaAGIHG7riGYhXpLLtWLIw+//y80sBuoRdEs30
TLD3MiJxljM73A/UV0qwusyDpfp94otnCv8cjSdn/lfdevpXZ60dKayCl7gQnzL8
nGOSmN1SI+6SHbaGO3v2S5Aera8VwGLCw9nNxKCvEt2QzGtP5H34ui7X+AK69iH0
7kbejvx3q3JDIM7G+RlISx6224dUchH1e02DhR+O7LtmZSMXUgMbkNqmncUESv/r
PkW9/9GCJQCeLlOoc8IkuUmnEVm9Haz98QyC0acxn2O2Tu41pDT/bhorM1W20gvL
6cbV0Go/0APXIfwMGRDg/x0cpaUaP4bRG5zVnydlCLm7uIfAQ3sRW9d67gOPNWLa
C44lZf+wvQFcaDfAAVZBD7GCAlXaHJRvM9CxgbKhTflHkuKMSAVSD/SMQrqdp5QP
0HKVF4oq7AYLS0DQcpNn+EwFJi/k7tMnd/eUuxGUyhF1ZstztEB555qaA8Dtld0R
UcEQIXYg0T7OQDjF1vzL7f9rpqHE91HN+ftiSsTX+SECdYLo+SVv9u3BiD9/xm7D
Hckur6pfja6GKPZVLujElKuR2ParrTYUP2tg1zjp/EZ+8f3DiMimLXpRLsFaWeNq
NF1SYcUsnReBjHfvqEPl8w+pAjhqBZud+VaBwXHSbGwrI0TqpcBLSSqavQx2ACeu
iB9esh3eez2WPHXGqWVscxebDb5j478R01g8F4szTgl2j93YvHylzikGtgumeVXY
bq8gdgAPSq4isqje2ybxQATtLhkLnGfl+y2T0NQRUlPiiMxnbgmSssh33q9yd9lE
522066a2zO7OS2ETyrfUVWLg+Y8aZHpYJBRtGXGL0LAMoxiydxab80hg+rFv+/t9
qEKtxdzE9gvR/qQ/AEGDOIUVDnlmgtkG+5g6T5MyIU1gP4Mi6utNivShjcfeE3fx
ChNOnT4fEDYqKiRZfVL3OLHR4hlPg+gPC5MbyaXNXu8AcKxgOcbvh+KnQGA3x8+0
4rHL8CcxXSuJkSR4pE/ZvqNr5Ur2SAgJYh3/LYFM8wCCmxg+AZyAnjfpJdryZSUw
zvw0dsPZfbsrshTpuaZSUwwp0VHug9GbDWXlrCTT6T/ABPolj2gJUc7feDOxlCa8
hg1qto8mytE4UlcQ3tl5yQrpPVZVI+z+M9QPNcGPYzMtKUPMq2Oq06YnkS/JqNQx
5QNlm6Glj+F0QWcuhOYi9uHNcNXa8fJ5JrQYLqfw8uvY9tViJoloVv65wOOoR/Ze
uLIaA3gWGkK9wiNK6obVVh2JcaEIwH+kgxk1q/2wjwe2p/oPz6cpvvxxD52BGqVu
sr9hk9zMZbLI30BT2ze4hYNG4MeHfnRh+OaIVLX7MEqS615L0TQe0ktc+wT85oHa
x0JCj3Vt3u3y6W0DTnQzODmjqHYD91FZWdXFbhUK0nHQ2AU+XQXiOoMdPBzZO92l
6qYewDD9+re9UM0mrMvb2ek9OAHoUTUa4V/mZRT4hJYvWq2jaTnSfOmAkt7QXMof
QngPpAfIYHnXqiy1W2wvWWGm6ca2vm+5VIDGQKfoqJ29DFlNh4TtNpUUHIGcadS4
Lbgsvj1z+hSDfss40LwHLmYdh6NqfXins+PP+AnJUot6P7CvRRvBjIr3xxDTXpRj
MI6kAZqbkya5pdGrT8FFceWFrZZ7u5BDa2WAyf5oidNrtXmWFUxJj35ZnGur9IDU
lobmqHblbzf0hJ4OobbkMvdwlnBXA9mQ5ydN02KHoZmY86XBcnSl4wi5Qdc3kRLi
Gr+coKPuxW4xhkmq4fLbUlV9JF2FsRW9p0tWMxDzLNEdlOZpro7mm0xEKTO3Sp81
pFk8idFQ2bYPPFwfY0j5LTf2KWwicAhrOKe2EV/d5ii3bD2H+nXwnq8JXoikInaB
2w6bkMVUBKo5hDwfqGOmVJzucIAtFyiKU4bDZxDt09MKNqLPKiB4B0NvzdfomizP
a/2lKhM8nw4tBGtKgkFTVMK2YhKd3++1yfLMBXLsXVKtK4wlar+PyP5x9e/Mi0sB
reFNfhDAZ4D7I1e7xfpqEP6Tn2Q2GsH84i0u2NhnKEwZ8xyumOI2t176PymCODmX
Sd7+Rx9HxiViHURIZW4ToVi+vfYHyzRaoVMm8jpxPtQSS6eUnQ9VT/WfCzRJj1t0
zKm9isX3YJLoJduz2wAYyXkb008SZ0Zz6pfhrZnQq4nZDHwbtKgoA0NCXlPv6p8e
dSwP0E51f0Xlz9ZY6dMq413qelc5qwOwmk81wK8WE4XXNt8IV7ov9zugMVqdg5zv
Eva6No/2ym2PEDAa3X1nih6xK9/zwlq7CfsiPcreSZAz3CznFH22yU8aVDf3svDA
6JJVxJMC5BFFCM7POjXCLgfSz4JI4UPb1tmkFHeOb//3Gtfg1pziKOfQFc2aGp97
AUDJcggnOA56vIeNXKtumPHrc2WxtWUygDaIikd5knaRBqk1buzal5DYT1fjEdix
oCfkVkqzpi6yFynqaGEWlARvECZDTc+TD5stUDrbgWdTmmg7C7ZUo6b265kfBrop
LzrL5fYGbnrUtXlOAVDRYpHiER8xTYq6sHFwBrm55qHW7KZjkcpoowu2pNjGToR+
WyQCMQBJVw6xOWpSz6f7TnseOaYclHPHbJ0FseOOG+xkVbQcxTT4qrteqMOkBJfi
UPmliv9RcuXR1Fpa4q6jPTjfGWQX9tuKQjnXRv8G7b6SrbcCN9MJJJbWntFmh/g4
lSCQB4iYV2hUqdFukvd8a/2pKVu+EtEXWVA5q12XJbEPVopaSbIuJMPLHCAC0dBX
geu3wi2fqrKbuFFXmISYduK1R6yWWmNAv//AFIgRixmCwxTVkwPEBbbLLOAVtQyu
JcrZnG/iR83csG4qaTZS2pl/jRgicJCM/XavGx99ktW7XDA6t0waFWFrJL7Pfnup
GAaO1R7QvCXYxG6B1Cqu8l4TAKnb9qsYrta62jaYPCAD+6cg8GZ/w75EKbcHaFui
BggdEuLOcT0YQ6b1QUE+yklCcZ5wbFYpkIzjFxmjJnvSkmJB86fqsnWzX9FhYWDf
PJ1zxTqMKXmg8UMHdcioLRs4FHN6HnZvNmLbiB4vt4TjZAB4Ca/tfrNHoOMidmxd
cS2UD2pJxnPRESrJ3Adied82b2u/0nskNnsCOFG6/MWh8y01XMvuupodRmgra6tK
KzZyApvW8/xepq6wXBi+qp8G1j/TFW810btpEByC/2v2diTc9CeAHnsImSjPZdp0
w9wWYS0wTIzNqwUhxnYvFinyThBwXBEc2J3JAr7GKe7l0I8FsrGguP6EEVC9TsHc
pfN5xkLJ8CUmFBWWQz3jyDx6kUAolgCwsr4kmpsAc917O6wVeqD2QwL6I9I+r0IF
01gcyGS6upfBb8uKCRlDrMz3FeD3nctAUU9wP6zrcHHWiAa0//tNStoI8wNl6E5D
d6+O6u9zLfpF5QSSVv3NVfyE37WnSE2/tpXyr8VWIskmyDo2PBzlKudqeG2BpypM
3jU5/kbIJ0crhnvKPI7oxyXsI7iccSslCH9YayNldMANYdevdTQjfuwXnNRAmoJa
+74TTNGk9XdZF+NL8FStLAmE76P+3cNiGaciaH+DXYE5vbjZwPcA9bj1DuyCYz8r
mZbZCRHD4Zi1QF8RqSsv9uRtJdt5lQNuZGRj4PqoO8+kIRD3cRof/NO0zr3RAGa8
Dn7h+6xmWuAtxocLNb/atvQb/S/aaJdWU9ZK00KJFfsCN5fxwVFaVsmeCPokbl0C
0EWkYUhEbdRSPHcYvJQr9ZOZNrtcDpz+CR/vkWWe1JPnwSg1j6tJ3xgnfpjk+3qf
cx5y8MllmmLDDDRBOu/xYsl0kIm/GtjUJ9Bjs6w3MHi1lzOhgZqh5oHH08qHRq8h
dX1RQgg1zcLs46+iozzklQLK+B+EHwU+kin2Em9OcP7EtEhKo4Zz7uXuyIJYWbU7
+ahrD+iH+s91Nyj00ln4Lp/+JuaRJzzDHhCPcVnMSs8XqpNaT23J5cLSxu5s2Cmo
5rwz0jfsfGHwJ48sVuRnFnGnn4DUIemROjrEvQkHwGaa3onfwgTPsgfsJkVXqSXA
OFpH3VM0efVafq4PfP5QuW8exw4EJCn1aVgCmrgFQEzN6/hGa6Y59ckF9OVJEPdm
KhXZnLi/udgD3h0mvvaM+g==
`protect END_PROTECTED
