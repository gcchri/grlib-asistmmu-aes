`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEToL1QcLuwk6IM5pCFd0mLkIc9GZvmQjIGGU9KDgprnFe4YEKBTYFHYlirnJbO6
7jQIhV3X9XiKcSmDPbCgL5oyuOuMqoINM1mKackuvVRS1TIvfDo/8eaDkTB98CxG
PgKSm10U0hd9qx1vNUOPY+Jh1uINeXyW0KeJYO7khVb+ukGlFeghilC/REozNEMg
QCfwasJgb3dvKCMGDZWeOzZd59U9E6imrulFoZOL1tSoiDMvYHQEbfzpnCmaZN9q
unc5WW+1n5IjsS41owliML96nEpLMdJPz+Jt709VwoQwphqTSqJowuxJslem/6NK
+S/DcU9Fw3W6CercPyVB3kr8+svgiNn/2hiW/qGvIkrSyAvZmMizs5NIPJ7vnzDr
/LzaRCqvWgUgRh1G7ZKnn2M+cLopyuv840Bm8qesNnqTeNiulaVvHGY6bOROJKGF
6DT/csB86Ker07fSPBHxj9WzmmAbfvW0mC6wvdVNkDuJiSo7MT8gsfFDJnVbFyaN
Vs5I0/nKzDi67Fi77IQMmHmzUXDbncMJXFP9DlY+Ah+sg33f533WLg9pZxbyDu5P
7pYQSUkmbzfEg0cjBmYRk17wJ5TXHmEuptFBSJ6IXbfSphZdjqDc/JmML9xh5dgL
6klMxAj4gCwu5bGCD1NWxEm70Uapbt9ndpSyKRP7ZrnMqr4tsMXM9cY+1tw6a5WK
Ju0Fbt/mhIie6JSjjoJ5SIVUuK9l/Ekz6Zmf6J6s+IvmGl4IKzzh08VDsYrBtT3s
OsW07Oz+b3hPmbGagUcXm/MJrG4CBfubxona7QxHfajdhxKe7bR6pGe8KD0rUexj
xalJZBbFzOyoBlDAQwet705qNrRZz4MRW1ovKcUwGF7WPh2Thyy2eRIXwSVbyODm
M/1jPolM5GzaDCiPA7/1lqoWcRJnfbzE5eMLvPnlECw=
`protect END_PROTECTED
