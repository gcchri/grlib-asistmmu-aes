`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2F8tri0JDJu4tRBu5BEItPsQJRa+2otjbThBNQavrJhUwikwWmb/pv95goSTyHV
IdbE0w+8ee3NWSMw3f7yzedj4jU2mU/cmB7yKYdUr6HzamPJhGF9G3ZYHdYGE2KI
jQ/xPkgC3U871D2q3Q6nKaETjLF0dVzel7dU/ggoIzSotDC6djReiOWIrKTlsKfp
bXBorlG4rKG0c2giO1jCPSBELycyppr415pqwta8oEOQ6XGhNANZvznMCQWBhBDW
oV/+oCn99lFhxnqcYfDzdsL2Rjwcr/+zfWTul8wwoeYcxSodmg9ljS+Hb9x7XozT
nTmMw9JQ3T3LP8dO8ICPtfGddKo02PaBFNE187NYAh7Udut0prh5VBHF6I1ryFLw
nnzIMMVvkx9kVigolxHDbuVWdd9XiAr7VAXAySYVylj2+kiwqkOCiotBLEagV12i
XthKhR3qa3Mm1G716MO2OtF+D8NKYBqUgqVi1ds1PRE2OayIs9HLl2d/oNcuEv3f
DBBpurtiI0Eby8IaGO64JIZFJIm9fsGLvYhoYyfrB5bB9JxZNm761A5DVme9zr8Q
wLChLQsaNXPGICdaFYGGLaU6Lu7DCDHAcp8AeXqKAQYvD3T3dDmlJX/O8m89G8jC
nxDaSFIaoWqdQoVnPuDzXUYy8m4CSJYJT7eXu5T5rcj5BEjPBk7A1uYtdRMGj12a
iJX7i/libbAsLi1jbqB3cGfZ6PNIl3O74g+tZlpznzMHtRsM6svXt5a5IwfnKyzP
hWc+AunD+gMrb/tDfdiVaeoR6bqlxxfuALEwS9roMktUPnhR7vW7OISjuC+wp2L/
37VAsztfaRI/JVGJtNPET6QsWDuwgwAp6QYdwo6R3sE8i0khYUbahQn9OcDXwkXU
cdZBUrjYHVEzZRdWqzuY+hcPvRia8E9HKozOt1YpZ3Q9CMMpUXyR8YomHSN8kuLR
/ENiM7wWyFY8r1quwgs1VKcjQBnomht1+rhCmTSiiCow+NunH9qv6BZxSfZIyYO3
iIGkeMyhA4czXb6FrL/7R3qmuOjOQfs6IzkD0Dq3mvqxlL1zPEgUrb4SJr+tBh1h
`protect END_PROTECTED
