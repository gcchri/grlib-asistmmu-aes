`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFF06QmvOPjRY8r8zIkfhK/paCxJoE7RDK3qjEVQLF0fEiVM6F3jqF+UgUjuUzqK
24vuFyE4ZS15vqbTNYrF9dlNRfCluhFQm0nwL+ALC6oubuV4ueqic7Rgg+8VrD6o
mhif4k6c517hBma1mJPNGDGvzuZfzCo2a3TH9eFioyBSn/uzfFxU113cJZjkeI1h
ptGHEFr/wysSMF3EjcxU0HYx3k17HN37j89Ua160v7/+ggQU4+BKdEo/2QekiAzg
CKE1ibjjtGEY2d9j2JVE0GtXWnkyx8sccXVrVNERcyqZ+e34crxR03+qaXC/tewt
QJ3POKJadOoK7T7GeADZHPbOJTmtU6ON6+ON1OnoHsHteq3EYOr9fdkJRRwQkLWI
6M4bZnOuFho8gpCKh6PJnag0pYf9bG1CKv3oYwhvrHWpY+rLRnVcUMGl+OIt8Xcs
NGnpmkib51vpwePob/rPGSHQSsmZpHxiEJNesZI8iqV4nzczNE1SCKbNGwRy9Zoo
GmNd3SP8NByQrt9bSOGoMP2j9snbJBqXDlmlvizyIaWOpyzJh1GslZ1wd7AIc73V
6RWd97TcZuigq6C4/385GwMbA1Hn1rmZQMFWSPRDzGmpRbacsgGz18Xp9T1kFglw
LZdW4Cz/4U+3Ao7FS/PthwvVX3TvAzl88PWpws607cg=
`protect END_PROTECTED
