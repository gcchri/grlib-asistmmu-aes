`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D28JoUMQVFetelVmUuZBNc79Z2RgFfToSayOPjv6l0pGP6ns2kMjjp1UY1+ESakc
e55M7id294Pi3KCI0KlQp8EcjbhlTneXPU/LASi7v7V6dKzKG7FsDG5E3tXq3Jle
T7PBfhROgb4NEz60vXqQW5BlED06MQNPpuZ63RiqJBD/BS40jsPq4kYdIEk9q9Al
ga73LiOobjhe8jljaalXnLNjokpR3X5/sKT3U9JnCxO4b/PQEUTPYxqc6O97rcvT
YWYtnEukqWooXuo8ehgGFJtu5wFqXPbioZzaj0CpN7As8NsbxgkyXgI76yFT2l4d
DXVBqFxUqJgUGfNbPc2UVF2IwZE6JCm+gGTgMdCe0IY4yAq4PL3Jj/5GGdDTHIi4
DgCh2FFxisOwYhCMQSSUTL2MophyEvqRn7A7bDOEs2HjpG7xrxFb5TeNMkEoxz1o
Rwxq5EsMUz8R2uCTl7kBTPS9QO+tOS7di4fCfVXFloZPwmqeK7m9qUMhDsap9gDX
LYGClA8CeTGzzE/OZS84hljjGSsNGSLlCgLD7LpicetM1jJUFSLuhEybAayZAPjD
XIaJuvAGQNnTnN26CWabWY8p9vFgQenHAptXvDyn+6mltKTNb/bgHLsPwT54INju
S2iidxNqwJhiXsXyu3VkyJZeQJzkQHm8CwkZxMvv7LPju2rNRNU9nILvEq23FQdN
`protect END_PROTECTED
