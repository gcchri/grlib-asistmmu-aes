`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rOQhRZnW0GsJacO8vA3T8CapsUIFo8oclqrOlHuKtF9vCIiw9r/yl9yc4c7/II1c
69wrJQrUdyBJswoJDjZDD9pZXxVgdEdfHo1QmUyySIhnBfhtAlW9QZ9GlOPxIq/r
dSe7k52plDI/n2vS6O/ylpZM50NFmb2KqPsfKKUjG20Y7vN6ZU/G6Xhs763N8H5Q
xkT2o0EaWzFvY8glkv5xDAxvHHxhuKQFhtbeh4Hjtc33FY4KnPRNFRyVVciOHhVG
6Ivl1nRu8ZlWO1BYlUZFvnh6s7pGWSFZMdhmQWoES3Kv9rNWFwHKDUzpcAj9ClMa
1gtcVJqaB+/vfJn1fkdjCHfQ2SB3h7HJ8ILqymL5cSCyJlEfpgl5TB2LyXSogq5F
5ptJrUC2i3ijPRLir8UBGXi9jynYjDwAMzzSmLyz/yxPyJLkOqFwBysrwqqxEfCg
p1F8XztpKYeWfhD9LoT0jOY9bHsZbLAV2CEtcgh/aWrt5gwpLG1JzAzg44ZDhpMc
qyF89cRYcXijnUyvKcK8EezD1Tyk5M5w/HYIKWZSyYoLBGyelvaNYd+eAp02Mb2f
`protect END_PROTECTED
