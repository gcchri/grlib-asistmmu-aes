`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6VVbDDVhvVuaK5A3KEzuTPHbNgiH91UweJKZEVnLNhLaiuZOGSiYINkvCRPTfSX
bfHeKv8opnlkFGubKa0glwEX+ebiqXdEU8HzZKMXo59QpaFWCeLf7t58lS4ovBaK
0xFe0xJTWwQeB1/z99y/IbWu5kQExZZ96cAlYMGCc05grcMsMUuWBm9h3aKhpikR
qes3avTt3ss+maduOUX/BcJRw+0BoNTR6gmlN9loX+CqYpZwlqLP1AKYHw8uOb0T
aR7uHxHeYgq8LzsFVlwgHe4kGNc7diAo6mmXOBa94GBlmoqarFGB7bRZSxBkAScr
Ou7f3h3K1q8+lNoZf7SJEiccowNL5NwaUbnuhsf83SjwyME7jOAJHEEZCyRCV7Yh
eDdrGL5v1I8pvr+Sh+uLgmF/AMlAFB408IpZ2Wh2JaKVEjnxq0PIltQYF9cbwiIU
4FlW12DJMfMI8mkEEUkZa8k7GLgoLo/9A4HM9wf8tKChjhl53OECokXOEvsrn+ov
fcXz+LynBjzmITGBqgHQAMXeHKifXDEpEp8jWM6WvOsikdeUenwI1/Aeb9T8xqOW
ZMbF4fVUHIIaLXtKXiPBt8C773A01lVSJCzaXwkf57uZHKMY8fQdv0ewoyzI7JcY
5opwFWJBFBb/ts2S2OF2JZG9foR9RsuDNFOwsDQryguoMLIM7vRY3gL4Ndd4cnS+
QJ25ROntp9DpyPRa14lSw8kCrVfbTWSpzQa0i7W0kkL2ijz7WohuXzCmfVKQz0Fb
GU+CWOqgAb+ZQxAj1fGgnTCclEt6UhNeddqonJnaWqjzlP6iT3Y7Dd/HlugIYe4U
jWvQLimJOI09YXn5MdLl7Vq4sF6YmxVnIlOOUakBEuact7F2KNn18kEDlXyKNDMh
7Iw5q1z12n+p1kn1BWqDoSCE88AGWnQNQT0+8G+n9/ikT2/pdWVMvCz9+rP+d7Sx
bJa9HbVOkwhNsZhd46kGj9gfVOoWFg/0yfYXzLzNFS2dD5HGNYQBum+gLl4K/idh
gq61OsQ/Cqt/aCumzi9lhH3jMQ72wTaeSVG0GdeLL/tyDTaNpWcxZ4TnDhoajGPE
0d1/W6RJp26fgsvh8KgSl96QEbpcpsaTnLWYNSZniTVFF1uAkdurliUOFMg6zHnb
5JxPxF1o8M+rrxBAs722t1sJua7dtXhyb1WefMunOJID/FBD8z1DPBYO7mYPe9IZ
DM7pbSBBqMW61CprfedrSz3KFLm4raXK8O4XswoIGxdqkBibY14p8Fqjm1KpCylu
8zBXTjmqrPrjc0KxRfyDm1rqxEOGRhLEym3OpgAZopUBqDpSH7Twq7pP/5T/xQsc
EmMzyEC/UnMpL72tSg3uVcuR9Fs3h1L9Yq/ddtL8xqcwrBjKQgOeE+4tt7+vpDAu
HPKDIPoduA/mct2r5hi7P2zqXK9WSWw9rnrn5ybSmp8t38GLzuxQcC8kqs2vnQwY
1AdwjxcOZK3ErsxlQOyhvQtBXESjBUKXrSc3MQVblSPvXQRTqOIhE7WHHLb6vkA4
D+duFYFRi3o9mHyCru8YYbxpYnRSpI4xkms4HVZ4xawsRrA+2gkFjbJmgi4QNRS2
R9mfyPIAA3JsrGFZHfPnXHEtmzQQ25dlMyUQiof4dagkg1by+5u3J961T5dj9jGG
K3mBW4/VhHzZee6yaylZVfr0mxiTVVUkGhiiQ4rZ2SggTZUNYFZgJ2smlau7neCj
VkkOodnU/VVFQr01E9+5t9fGXHQQckzBaW6rGgQMMi+iuwAnKVqatYRwi7GgOJ82
stBjtRXY8JdP1VFVwtf0l0I0s1CYHxA6MRzOTH+hHGWERmp1AiVB6fd5LYYSomE/
PtQelZ9tu/BRM6JqbEjviXiXVHTzPoUvAMweVmrr31uPbo77e7Sw4JAieJPjj8kC
FSY6eoujs2QuIXc/NnSykAIABjCC6T4s17oOccHvJVBGf/WYa3BPcjtIpkvikDt5
doAsfSSaq8dJx3X4yx7K3mACi16wH56HblnTMxCQXDHYwupvyXhTsZhZD4sa7KiO
ecOVyHUrdHZJKE6XfYrNpexVRmjoQxEXZuCW6Mf9QdyvHJyzrCL494FQHRSn27jM
IOo4uKPiMoS7Q9DeosrYsbz/GYzkKsRvYFAc73uDGWw/lbO8NqkkD5DvKUncyfUQ
zyEcCblO7Tymzpo5VcIjhxGNfEgnCnEVqjU8sLszj+O/LPXhuvVI9PpuPPCRn6X/
JBxg94v3K70sXKsztujN6O2UCDagmgeAAhM4n3Mlseu5skkyIRDMFgJOdASAxpvV
yiOk05FPpSpuhbvzIA15fQ==
`protect END_PROTECTED
