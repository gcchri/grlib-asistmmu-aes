`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OfQ1x4XJS3B2XUxDBwKV77RLV4VZgzGj/Idb9ibdXbciqnHbqjz22k56eMc/1kXo
lOrHJQVj6jPA6/Pw5+JS4yjglmtEIMgv0191+IWdTKo9S2V5GfB1Te+ZnRalFnJI
ZarTHgPKbOv5Np6CjVgwO/nXUqaITpnH0FG/QhXHgZOt7fMz/KPEWwhvsq4jOAVI
AM7zJgPnHTLF21oaDG7h/BHKxuEkBaVKIH283ea2fnJYNQq3HqXXkjv6lIeMCc8+
O7bnSxRGJz2xnI2aEnMjD3d3yzhQbiUaJVW8f0OknEAxKsd8wHGziOjP2bV4bN6t
y7b5KAaYU0Z7XsICrPO6CLVug+q+TgVabXV6o0FFA6F5ogC81SlV7J0t0FyTITYy
c+JU/l8U8ZSsyAcgkBptZavQvP/VK7Fzij+pLaz7lKMz0RuxTDZf/cXG4O06FWh8
G5HA2mR/ruqzNGQRS8Ppe86A1kC8rMIFKj4yZx1FxKfYVN0mEbFzeBcpOraiM/fh
FFEV+xt8zo7ZKeb/EDtf5C47ubyWrurTeJil7m+8Y3cSFfvynFKse44zUgdER0Yh
OSQ7jQ5JIgKp2y/wpDgXeya5mlh4/2xxs2dHcinM3WW3wdD764obb5oMjhYEkoG9
+jfClHplBUzED5mkVlCvLGte980Z+1mveFZ+o5AWOkJvMrrP9QkVAIaLMRnV+5PO
MSkojwQEWeTZ4fIJoVVociHIZTiqKUDZttAdqzVx11PuSKL/U+fCa5Tyb1p+KriV
KQOYPs2wQVWUdfmr7BiYvjd5osZ1Qy2cPOL8iOzEGWLip/OBe2k5JECP1nJ+IxFS
i9tT5g1vF6508uIOldKHDN6SOPWcKwXkI/+5++5oVfCLT+LR091BPNs0j1bn/1MW
t5qmDGzFrp32Q4pnnqcNNbDQJ2SP0yBjVZTECcnxFVX/VKrdDI3es/o9EBTJlckG
`protect END_PROTECTED
