`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NOb6D/W3dqqaYRC5j6dJo7bhFrignaj9dBiMDbrKcIX0694AxWHo3JwQ8wsLMaaZ
bbeu9H/Qm72ZBF1QHzhfxvM0hY3k+46WGULkjpFMCy+3LwsNKffbJ3k8BJvcQD1M
YblQul7j26qfLE+2pvFHe8QIjpn1sB0zeaPPxGU7xyHS+OjqqzFkuiNphJEojVeg
jrcU+05xvRE3UUEY5tPondBp26L4r6l2FXC0ivKxku1Vl/BiLU3E90GVgFx23wFc
17NYhDsONn6NeaBRkqmQEeINTBYNJ1sR62HyvNVpm/E0AutBkpMD6lVpkZywTsMO
LqYH7K8a24q9ut/07FCQQnBZodILohsW7H+Qi7KtjKf0p1tdvXr+k4y0iz5DIR1V
JymZESkwTd4gJA8P4pTTm8OKQ5NVih+ojAFzWZ8S+2NW7jHtIc2WWmFd8ZnOPPYH
AjjCRdxWM1LWfhZdFaAllpsTylMAunON86ePBcAD0xN/dqFgYwBu2C7m5V9EGIRY
NlBz2CQllQQoZZiy5ptQKKP28ZPT/pBRI8qGFO5pKE7C+cjTYuBIR4dW2iNGpA61
kyYOSjJdnU40w/JpAXr8trPbKDOxNtvCsHn1MSLXnwOx6jVWaVAeWbdiG3OLIeov
c8Xs3GQZkf7S1mHNYPNJ6w==
`protect END_PROTECTED
