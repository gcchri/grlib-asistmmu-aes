`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7q6oKAjLCUvgO39W3w0B/qi1KdoAQO6BRnIXrBAApAfKN3GOsJfOnKg8SpnH+1LF
D/xDbESq53V6ED/xjb9hgr/cyRRILV8V0mSt4qmrrJNCJeWQXiGLSYdvNfUwMKV9
0yeGGZgxk2kawcFWycKLoI9AL/CpF06Fe2bICMtVLKVjNtyn0vCznz+NGNxCg6UB
tID1dMJ9MoQape4AjxYIcnivpXDyDK+G7PipgZeBeH8O3eVV8ghAnDQcmS27/Q7R
zjqEfTitUFdVJfjE3asN4oyOyqYX+gEnIINknP+DJidEiwqb9ed3TsVYmMqUFCCr
oejLeGmNaV7+o86HBpkUcA==
`protect END_PROTECTED
