`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZJ/L6H5bsIQlB2AtK+AiwEO2Jk4OxEj5aHw3ZgSCpKdAq4Tx6QMbWHjNDkp4/WC
z1ttON3SwjRD9Qmi64h8PJ+A1I/dtpGxPWIgTnIzZhx1TqVujS9chSFsBjnfvUVY
R+muG7B7L/sg7SWZP6ozu1nG7R4Nbfiht5d/5ON6+hksem9QpTGP/WFB/C6KCxyR
b2Ttw2MEgksYMJZoeX0K+2TmRbifYNBgJrvw4sVmLsCBlhPjAWra8Ui9MaRHXRwS
EFJ6olGdLVUHcl6Vgl/As21D/U8O64P08TBuigMs2v0r0Aud9QbytYBnQq6N7MvH
K2v+rSvvQNoJw5c7n01sPTD74vfXqWe+YOWyheNi4LntVIlZt3dtJcTmpXPitNzz
v+ypIXzNJ0P51CVEe4Fn7K24S7S6pn8htcly++snC8mUMPZd1fUD/hAmNLjT7zS1
tgPlx6yOmxkUXxOQlGdu6e+dTqnq4ik2hg5SSQWEmtP+RW+StIPKkU3PcGmX+3CB
Z6e7WK7r4Q3jiOi041K6FyqaYcu4pxSOoxaNcdqRrXS4xxEAxatEkJzcgokx8g1b
kykiqZmGKO4wvUavYC/21ILmcla6vubeQJXr8Fy7oqWEdl1kqnGZYLLeL9ZRC9+S
Y9JYlsLhlnlCs9evLR5s0k7e4fqAunzJMWpJX/RXOiBgVeV0wwCmqycxjw+xtvEr
3z8CH39MnOsx9pKfNcsltwt5ZSu2QnP9XlyirpbMDT7TZNFMF6F4YY23ybW7MOJu
Sws4RVKOef66JIieofOj6Stp3RJRez1XrbXKyq1e9gYZbcev2gBB5fX3dHi/sk0x
rSR7K2Ffmi6QRibkW2HW/johmDx1NooA5qKeE123akgXwKQbAagV3ZtTkc/mVVFu
N/0PtDm8DvFuyxuLlZ3g5Q==
`protect END_PROTECTED
