`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eF7sweHEWfbTTOcLm+b7w+EqPevFaRLNgJQ7XcfSL5W5DzAgnfYcRiwxXcnu4K9o
WnAy1o8hRQcp7vvqxkK7c5X5gsGPKETQYHaYQOVr5kVcqKWzOBjDspZev0R1CDPX
irqrwYwlDgbL+B1mvCBQqlTev/wOZyZuJd4Qg2/mIcyLp5CeeybgV59J8JRWVlHi
NkOlibFu3U8KTAwMqwTcnK/AjDusszt0AzF6J7KMkzJipjL4shqwTYiisD9BFPz+
NGkod9Dhc8NAA3SzyXS+MAxtc+iHDK9aeMgMgI3EMAMD22BFd4YB+FL3neKbyXuH
Ihc/BZyKk+ZSXpi44T08qApGv+djoYDLQDRH0JhBSeD4zaWTXEr4FENLIaZID1sZ
MjNMj0HmCUfIfdgsA5Jjg12vBFDCFcrUIPinomQ0W5b1ax7aSr5DZbdmoxtfq9ha
28ipbRv29mohxQhbeUKMYRTnNU7FwvaGEB6q4Ign5/vR9iwF/R1+cSxagxUPU+GD
JQfpzuWS5J/kXreUYgi5yjZ/AwwclBR00uYma4bBq2R0PCUiXGVGEewli5BxTaBV
wTOy/NCL4JdlDY1tbDEGQUmYdyY4zD3PvrbAQtV2ttTTsfoFOEYu47K0T+sxc44c
SGImNFYogWW5ioojfM4h74kuyVhR2tx68DgPYAPKegWC/zACYUzS/1VMzY4yYsyS
8ji4oZLyf+Llx8J51AZ92kR9VTpaiGtcZaPiP0woZIE=
`protect END_PROTECTED
