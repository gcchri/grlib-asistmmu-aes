`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3bSIP/0NYURqxFUrwA3V4tD5AdCoMaS4j+tdzTUk5gHgxZ9ne4wtrsxwYwhvz4l
uFHYTcR0B0l5rHpX96zp9hY281ASytJ9cofT9Lcj6ozL8zIjwkgmOtdqmX3Aopei
9nvFdzE6mogTwnxgCiwT97M/2kW1hY5gqBEauvlRZZ+vVb4+mjRbgZmqSrQimrT9
IKdFdseRXmY3DuSbmk07CpEc4Kk1r6gcwwN28OBblr10MMPgGSgR2iNcTlTipZss
0yV1pxyNWQJ8wGBYIPRKDltZzY0wQiI/5vpDh/wYPlbW8fLlOYpVFawGl8vNjKci
K70wDxpZKHTkFJVfP91sYhgWETVjIH0Lier+GjTDPuO5PMWbpuy3d/DkvgfEG1eA
tbnCK7m/bmKkACya+WSeU6esSnIMNNDiSQjE+CIA9l9nirOcyr/zFJdGSUwOywcS
U5osWvpVFJqH3e6aNniQK2aS+FkkviAVNQana71wzR/wExNPeo4rJ2Bxsb1ZRCiF
Je1yYC/KUWc4paPDNECfYLMJ7SR2ZQFxLj7wO4POV5wVl9QOHDmyEewj5S4YeKus
UHITjsnA1E5aIYFzHYMW7YhINsDFVzLvKRh6LHLt9RDJonqnjnctX7rlwl4PHxqk
lgoMd7K97feIITWylnMg/WMlV+XK3CaYL+P32GH9bI0=
`protect END_PROTECTED
