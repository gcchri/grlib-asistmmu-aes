`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYccaN6gx2J7QckO7YCbXwjYA3EB7QcNTUuZ+uJueHZOMsjP+OVUch8NE1EvPQ1+
rmuCVWroscUXZTcFbu6grivgwL/s+yfn48bFg2jMfbTsz31QZuZIY+5o8226CId6
s5r5j21YUb+zEqqpW/xefUs9i/H/opmlPWAR49BEi3mavU8KnyZkN1A7OHzZ4vKf
gvZpyT9M92viUJDPusgQktomA2LcO7KzY2NbdJlExKluJUgFXTn5O0PlvjnZnCC3
7I7C5RnX+N+u3kjMmlS8WQCZii18YaFX4OD9MXtepittP8SnmDB8EAAiQZQNlhbV
9TczGhinVp0NYeY7QF8ZWalj+3AQkuNnrreDlmBFiq+FS/BFwv//zVv1kGNSGwwh
mWsTRHROW9zJgyFpgYtTPcuwQoKuse/kXXp5wNNtON4EBXjqGkbDI3lD+vIhVpTg
DWA/e0TeC314K6HZxL3aWg==
`protect END_PROTECTED
