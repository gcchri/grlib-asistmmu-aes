`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqOg5y7F1kCOhY2iPD/8fZeJ+fEjGKBZglm+Kftv5nceM/7zvlHEDaUrqQulCT5s
azVhCnfxRNOl/7+zaeT/wbA4k4aeqrFVq1/3aihkOKkTVfdodM1shyPNJmbamhkE
yIVddpXEFCH0I9xdsDEjFnzMlPP7jFbAa1jpzi+sEuNYq+8rc4/JiBEXuu4XfHCJ
ZmqxeoaQNK9jWE4irTDb88s+WY6lqpE+56ejEsCNkQKbQ2oIG2jqsncFJk7BnFhM
OcPYLjHw4LZkKVhsiAUpbbMS5PxoxKgyBYvFO7bUxzYNrll/q5e87IRxhJ0RrWQF
IWe0/C1KqN7DpKR3zHRkYA2O+Gi67hWl2NNp0IszV1lC0yQ8s0z0te8l9S4/I3kT
FKEi8AoYpUhC3u5nXkoP1yBG0DaklwcE6QRSsLGu41PHITaY9PGEMocsnfqb1UIn
5KUe4jKxiiIh6O1r+4m2agUrCf26DVRET3bewRNJ+CzvdjyK4PeH879w02GhI2Zf
`protect END_PROTECTED
