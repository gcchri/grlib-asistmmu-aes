`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yoIeteIMIPj+Xf8QlZNpUwHB8XPn8aqmwyXbhEinjHnca6eGlkvrf+P4Ke50T4W8
PQvLNGdDxWHPJ5pTmOyBOPrbEkqXh1UAgJZX6Wnd9UFdTzqKMiLyr+4CpVim1uZl
zAT/+LPZyEv38zfVaNseEQckL/Rwqh4suYa6NHcJg8xbolGHQSF/0RHcMopFUIuh
wFu0hDtsXZ8ocu9FHFZfk4hGV7iPlKgRwgq4YtGYhbDxMxm3HFsK6apvZGjva6Qn
U3MY3l3vh8UZYgQb7EwIoylsLGGPRHQwlfwmMRwsE+ZcIWHRM2obIKNlW/n6ZZFO
yTz6z79fdSlsxRJwyEp3iM/l9vF/PEzqDP5VQfs1d1/+8XpJgRf68bJ+7dvcU6An
/+gN+geXMAJiTwzovXmNYpXpwgLCS4KeiOIQckpdtm/8jxpdoU3gJvmr0s3g1KJZ
svO6PJp4JK20bkP+P6BnVUuBEm4FEb7F1Sx2xyORIS2mwyCFif82whvK3U3k9FrT
i8sMXLcdd02YazhDSTxCj+oet/RZdJmv+kh4rEg+fwIHuLIMmo1ZFM4b/E6bmyih
UgwZvji+MJSUs3rtyWCHAPIOKMBfHWne5g73ytkALZsFD1Zd2t9EcjTkfj1odTav
jq6hPv5P+yVDa3Etc1+H1GLgZDOVwspS5/00lAh/Ih7YHjgDvpXzQVtVdT0SoDEt
fYOvxoY0JGLyKBwElzMDVjFaqOaX/bmjPWZaw4BupnUj6Y//troh3m+8QAEv15mS
OD5nLQ9fFdnCVfMphNljTyNGUPWEE1Y0uzsG+emg5OH+rbpE4mXU3cgjaHO4PBig
QgYZ0VpY6aSzM20NnFTryfLR8etf8gZHZkBFSxZr8Kzj2FPsGIOmR84oHQY3c/Ev
gi4n2txFb1AQZ7ZEx4JPKVpBa9uk0i4EcXhewELNqAnLL4Ikx6TY5zzHYvXLryTv
4M3+JYSXeDdrVvvH0JkuhgSG9niHHFA2l2f9YGmMG6waDVIL/ehqQro9LMIorJi9
qP/fydHZpngv02IwzvrLHYPiDCHW/udXVMORTrX+VakiJ4kUYG9KhGaf1E8q8N4t
tWGfxc5hCpVT+nvvS7i+7O31rHWeS7LemRRsO/VhGE87cN2d6qB9/eYWT6d52Rqc
4T9nkUSKLC8QH66u9Dy/JnnRoFLoHzGxYF+y9h85OKE89mCQaqJqUpCSsTeG/cV1
1Y6/s5JvN9JPJ6SGnJG36wo8ZiJZLUFqKPqyFzT3rH/3BCjzbZxHux6H5QyZfTD4
86XouU5LHZRkn+vw778cuMhn0xDn8+YmKPQvw7w6Ya4=
`protect END_PROTECTED
