`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qAprRx42t20KBzCw2nfsoL7X/WbUf8oI+TBP6ybZ5SPpZNntvrbjRBG4W9i6MEk+
RAS5aMuX4gRtvsx58/jP6guWlecQtK8/pBhG9u95ndJaMYN4am8Ks5MIIRb9/xvk
/285+w1h04sebRdX0q1g24l00pThfl4GI/9SdySVKQDOX3k8oVlAPBc6oPxC7OH2
Zi5JB45sgysE1s47+koZET32Lwk9yS1Pj+HegMFU6YEh/q1KQIqUxPAurnA7U7+x
7x7J1KIPqzbtrzpZpMwpsU4HSsfZa9qDakmMQ/pH+imFnT3IWQKsiQRWb4h8shal
4q8OG4wIKtbKYRa5tSFPLaZNVs5fzbJ9h5OBWLhzK7LdHaePXnEhtJS27mjgLIFP
WN+0VuSYpaDPVGi5m0KA+linbm2oldWNERHrht63yDPliI2mY3E7ak1OYxexQqXg
hIPDU5BLb1i8WorgxnZyJp0c8s35gK2vv0oH1pdhm3eQeQs3T+gCUzrLMlHR8I1V
RA4m0TnlURQreDmCLF0A9Ha17VMUxXZh5onTXQ8FAy+v0qIRfvOLgfaHXh22wq/a
kjrcxeTYbWuphSXpIHiVvZ2qAdZazgUOOGuQNISSK7az0HVCf+1sE4M4MB0FI8AN
f/dMvXV7g6P8zLCMBN2PAyRzlDkR52AF1B8i0ZNEOxbt2MVGIG66/MEtAihjEmU0
OgRsEUaxSlBY4pqCYlj4L/CUA3uiLmla3bikgHiXyD7GfQHoTX9aeD0ziju8nyx9
fr17RZVJ2P378sY0jFlehSMnLf9GUXEl0RGKU8N7IEKVtND7iPagLMfcyj59X+o7
bNYDVkpuzndGWKr1FoIa29dd84f2YzjOcnlN8zrbc1UrPK/wiZEOQv8FyA2YOOFu
yj9Q64ERCkvpx155M0XAVAeNEdR17xBVFf3JZAHsM6U+50nuUMiylnEPw3FoyXY9
NpOzh9WfNoWxZWFYGLRZAvXV0wfYNi9yiPgcM0W2RbWeBSdsyNr5T3eLHtp03tlx
KWt6tZ5azI1c9V9xXmFXLnvVYL6Jrgst+lDE33DRxGwwm9wTDU7iNdR1HTR7KBuA
iv3jac7JDYnj4Qkp39eAwA==
`protect END_PROTECTED
