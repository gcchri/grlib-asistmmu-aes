`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UIy9pHJba6GdvO7xBet3yCUnAxmXTFoqN6lNzzc6VhSlm8207ErTVWA/FlkNcakn
A0XnIMVDniTzkCQXbapIzlZEvoMrcC8fiMNzd2ZZiBZjLxQ5axcgdTxdmFmdMCnf
DIYFuJMUxg61ebawY9SGoWow7403BncS0wMnokQwGp6VjI2yMLKzX/lMD5jLb1eV
mRBEhy9z/51KWz0WYnoj1a6qjqn2vnfoXjIN8rlGD5M3F9DWY7KEZrelM4qPaYTX
eNoXfmPyQiLZGtHIC0WKh37x1e+SGUlCZBB1KdDi6Q+4kx2lnB0TYAKX711Lj789
3WAm6gaHMj6I5OAxnqs+qetcZsxKqFlzN/OAlhNglKhJdht37wwMg3AYDW5YO9dS
hFzhEFJE8eChk+1vMBAvfRvEOvUOBCnqb9zqplNui6cZY8qlV6LUSDJ4ymNCAWcX
cljIDbk5HlhbLPWb8rMqPf1yjmgxw9M0/wETRUGVO5jlu3zUzCptxR4ZUOQd8pUM
Z2m2YFfDDpyXaFW+xMUKn/+KcMCTY1NxWZf6c4yCBxrm5fcJM4HX1+2EDhEn9AYc
8qVAU+8zxKx4w7OgT3Vlt0Euj6XxmVMrrh4MGdUE3wPmkGfd8WX66GjAi/UUegqd
XF2SSzPoyWEIeGXQ/uACxg==
`protect END_PROTECTED
