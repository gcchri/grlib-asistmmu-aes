`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2FIsi410PuBxc1J1cr9RmNhzI6tDzY8DTn0AXfSQ8KAj0vuZIlaLeFgByubR5tpc
Y8xr7wkhVz2eixd02lwZ278Zc/eCfVMYlQlt3CNkaC4s/9mguUmbT6aM6/eHdYIb
L3hQw04aXKLUCedMk05SyoQk/J7ihET9qaQoIiTaH1Vv5h9ydJV+CBq5jpk7Bl7i
Qr9GoVGuPg+8657UqVGrYlyy0CKXz3a1gV60mTuu6/ZCktePhlBM4Rmu2zi7vn6e
xp6U5Yi7xLCeHHn3p+wdbXZCbsogda/q5RgAcarAgeYSN0SEveT/R8V1zC1I0OSN
qe2bz2fX73iDkq+TQtPr/JnCGoW6ibU8LLwroFT5DXs7AXn+mq1BK0RnTaNqiwXx
r0iTqiKFQ07Zlg8I+O7ne98XTB85SHx++VfFSnUZotsohdVx3y6jWDgETjJ0Te4d
gD66waowfVSQ8bzn4UWKPwnL1EeDS84ZiH4bvK2EPRMtiYxe7CVjrl6YSVIXjzbs
mCQyad7albt7KjGrxWFTt8Jb8JfDWRvdg0aAGpYZ4jENeLkryKe0OYUoxWhqW+Dy
lCikUGcADID9jBkhRmeOCQ==
`protect END_PROTECTED
