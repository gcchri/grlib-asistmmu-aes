`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Qugkq5NezbMil0/6vnaPicvJZdh3GSUMcdJ6dBVm2cC9dc8APRclSogZi+z+xOD
vwO/5zvGyxtNx/KpxTyUTcA/ZKrEJ2xL9w8xvBago+rnzZ8U0MNSxeVYgnVeJ+CJ
0AvzyCe4LkSuYbKqBjFIJ5jLIgXQVD5w+M7UYyuRTClP7NlzPK/hWA8/6PHWtyHP
vwonVMG6jzrBQmq5LxwYf3ufy7IwxM6G9BfxQzF4Q5PBfDgleUiE1wZGzjmHsKYd
5xlMn7cc39LTBTbYweAoe33pLm6Wt2kbYKLziAWUtzwBj8MoKjR4UqTksU9IdSb0
o9miij0cCJ4ORmVd/R11+X8BPrD8M1lJg+zEpbFJuzrETXz37RwMq87344UMXEjF
zhcznQ6fAfYB2ZEQYRfm0w==
`protect END_PROTECTED
