`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vmuy6qyNRaTipZmVZrG4uhLO635eIb9uBaC/+rUzRfQkGWL31iHNRZcCepPKXkEt
f5BMBmpgFmZdGd1EbCDT+rLyQNYRSTEnK8m9Lno8plcpzfRmhMdBeRg1v+zmVFPL
exBEEk0rV1pMfSvdC8igCrGJ9goN9T+fwrIQuEkpj1PrB3QRzgC4mMLI2SyH+ZyP
CzN2XMvcyzlw2RldtSCX7Ojkk1EiCjVSpttUe3pwDcs+xHugDbdn4wFSe9nEXVjo
V2buz5ULTP98QvL8OB15bJ+mHkvSviZo0EmLVG/LthIvcJXrpaHYF+XmwT3zSF3p
c5BIBhMhbJhBuqs5Ytr6UkMPiIlnDz7t8XgA6n6AS8QyAqMD8Ndok/V0CLbr+zhd
P/fKw0SrK7UJQsVcp3HSX4FCCu4E61ht68qWvi8bvWX92kzlTqP218War4FI9Ak6
P3PTzb3yZIOTSZr5Na6s14TneqWIcWCjFdK5MVVOV4z+JKIen8BRlGzjgmrArVLT
CkHD3KJHnUVVCuVQ/t0+aRA2b25CRlG1d7tNMHHFlG8KPJHcJb/Ikwxwb6R6zm//
DSRemYskMhIS0FWQhx43VvbLgi+qwoSv8UoypbjrDYKNxMTBbnGWpETD6fuLys3i
4Mjwol+/2qeqR9zEVNLu3ppk9FRHJ1NV3DHZui5jUn5ZwRfRfQtPBkBHuiUEPIJm
9dE47VHKK7JiKqwbd41i1dKlMvUWpDe8DNsYw2JtilqmKFSSLNSVh4IjNkyBxtlA
mSmYDuaUTc8CJNCAxBiefDRSOHnenbF/6uQfhtGG/uyNfaowdENywFuqaaUDKfrv
OkFcovX1Obfa6Eo20WKbycV/pzfpsyw9nWz74CDsO6kCJMsgqBY0tk3Lw6srCRF1
ei5ZUzd6FD6REMFkgTyXToVCEbHHbPL2RDGP+2Hn16qxSflXpkqkjq5Aj+FW3Ikx
91ZvWpsXAEcekMVl/ITBuRu8z7gOQj0WRCj3K8kUOpRuXbtBiIzmIHEmu+xydWgZ
OxFrE3m0ZWrWINb7NhjQ3SSrfeqld6mH5imwZaH93+YGoaVNtslTYgG/R0VfxMBr
2jLj4yAfdBT2s3FowEaIbbW+6x2/L82fwNDHS/0OwDa5y3w7Vjji9egMn4aQmpy/
1/7TwKopb4gvZav8ysWu6lx6oZVNTJzGPTK6yLlrcAdKWCBvgosmbaaLKcuQBjl0
qdz+rH2qPGDruGL8kp+uLdDZv5PuA4uS+vE7amAcBGd5+5O8GDL21WVMROqr8Lzl
FtUdsqOWrvU1n2nGb0IV2mh5ggthrOFZEtKIxb+lAx6aJfAT66pT6C88gKM70wIl
dUB8A8OHYnNAaY09hjvGk9ZVxjardmLv7X4zCIJmGWLNzrB/m4IggRFhfp/zkK+S
1rBF9nHL6xILJrokOW/0ZGP4Lb9Td5qNzB2ZTkrW6iEu/e1zf5WyzwrZVO2mRxTC
1uOsVv6mDqNcgw82PQwaXeHCuoC0WVf5cYn5d5rzFt6RsuIy4UKs1XTTfTbZPNJT
CFgKJx256VkrwxmBY8yCFzFy9hWNnt+4Y8jf2GMy5XYniPrxCxcfwZHSleMvm4jy
6hV5Oj5s7KOlPiiAZI7j1v0Xoc04D2g9+MLzJqd1Rd19qu9NdKycG0yMGBP4d3ZS
S1v5BprhjDqXBPkIdHxI7EgZ1p1dSEnUGk3lRvSZN//Luu2+S/2dPUPdc8wRh1Oj
tSul4PCRT28vF3JGpDvEtwCKrHO9Kbq760nak3sYVz4GPI/fQf6rumEfV0Gobc9M
5TUexnjzHIjGGJIFgMr0Anl3dQnfdXkrzy7U2W90R0DY40IqSvihOY0hE0YI/rK9
k+NVv4G+Bf8/3ZH/7Zjm1RcbBZvJgADgXteMw4Ofx4ps11wtSbHilS/zTYcQtqRL
OObAXhxB67F+NRkkXAE34Op1JM18CgXnTv8j6Uyl+LNj1YdVx0I4dUD+d8pMasHd
3oBBjevLQ5oICCyVifWLyzRNwrl1uAArxP9mLLWrq64uhjt5S3KcsRjrGEDRV0I4
9hfrYGufKodqv3fievtYRRSlZDakrqtcD5cJHZtlP9Gg4VvNEdYtvcBDCNrGBSaz
c4LeExvIqNRHSitja8Fh8wS3kzbQTbzs29mjnLGzTtDCWlYQWFyLJtXaZE0K0D3Z
/NGI3ZQpLrAk0vwm42A6KSq5lVf0McSGTqbhuIJhnQRwRaMdbwEPWhiOL5jK3jvb
F8wazUkXWf/uTUJbzcpPwqlnmU0QcNQEzVh8jlXLKcJVBlvzW1ljrL/AHO1F+aLz
tGHguxuvc3gy5uMtUKqIfSrBMkK+Vu1kVPluR/gPPITumy5XyXuK5Rx5KE0ondiN
jw1dhC20jzshbw1qz1DY+NNwHLClQrAD5cjIJ+IE02H/MXFBlhpcjdez7c4DkjNs
TSD8r+fTKpIm/9Fup2/god/0w7SvyV5ovOARbYhlnX4eqwdWgGCxumXP0pKWZ13J
IkJZA3zQc7hEOY+Kb2loe9SBl3jTHNPHJY/UcKBGDVIu0qsZjosORKUQg9PF2V+t
ESsqOWER62uptJ3cVTo2vJpwDQxbgjYZXF8tvViBXF8Eg+UGLd/8xcZGdJUJdG2e
VYVLEmp2h6cqEz+mKsHi3enyVEn/2lv+O8b//vZD4r1Xu8IDNAlWBrciEkPrPGNB
RD7SC5V1DF7u7PCdp4Js081S2LhfK5FJdoYgie1c/7hjzFL98N3kC0J+E1AtR4dE
NHi4bZpIRkVDcRu2lWliUEznCS5ZFfv4X67uNiUcaDHFz50TGM7nHTQS+jnly7mc
sWYvOV8UUJ/06GQFjvu9ag23xYZZFEVK1qKmpRUHfYPO3+/gs+U2GEfwCLww5gf1
NtjRrB9JTqYqDFCP6w9mzxVd1v0kI6qxqbi2R/npwQ4FbC3DfYr2IWCxf0G74mkh
Rs+fmyYcKNY4ncOjfobCcMx3SipXrc00GtMwIltZoX6k2NQpb7BhLLRA4fOzJttY
yiRNiISYfVb5A2MD/uUWi84flHt9NgFxlroZnJc+8Jj6LKoKJw9jjOhZKRGkNyaC
/5r3606nKAoO8Pu9Yw16n52fN2pp/frlytpcbBWyS9JajUlS+fIfr/zhfwWxgiAt
9PlHByk9p74lNGZ6Rko4trpOp+gPBrUJZqSAPd3cWqCFjpjU0mIBDlw3mX8hTmn0
STntDHJAttELuNYpB0T0aIEs8LH5ldHJPR60D5d7xDEf73V9SZniWjDUwBRE2KtE
uRcpfakKOPA7i/6iKGHRgqMT0RU8feeE7QfiDsoandhsIuSs6eDQzlnEBIQmJxt/
9ygwE8ujiYTwV7BhVDeGnPwGuQWg1iUuyskvGgmfi4TjUiCfeo5rzkFmVym1FbHI
SW6lxCIabYWamBWMEYWNMl1uwpfb2Cf4lp3cCQ7CtYrJoZ0IGf1JSmE1jUcafzIq
WSlCYwquyzPKZjyBSXsrnPagr7L51QhS+iFJwKiq+uE6aa7+ZqeuVDaJZbtxhbBU
T6KpO1rz4nkfoaHA8XzDjfEGtj5WDbJ79uhDdGkkPfSbi3S1PJ+KGdxivq0QrVYw
QoAd/APveWUHb4UptKWeC8pPqNUI2wxvPsBjEd0KN8YkLDzeDKGUVrijDuNRu5l7
mk1mQFxC10HE/WbEP3MS8xFLUOTlhTilbU41itqZjW93bSc1qf+SOo/F7cipgRrx
O/zjPbH5ytPlhEP9K7t3/WrWCy2S5IrIv/+aM8g8kzSPTpPFTdhE39xUp8mXFcTN
7Y7wUqnBtGyUGaW95KdPkZs8rWy21G6SzKKblvWPBwzlZHbnxbHMECxrt5ljHDLG
vUp5dnEJAXv2Hs0V2+lhwZHWhOFS7ga4Kr4Eiiiptuwh9Rjw/gHHKE8eC6yz/p7c
AVO2a6f8cW/zdA1eBV1FPlvzEwX1b3ewgRWOj6kyMIETlluyKOrMrVT4410zANCA
9PqHmsxbY132sECoXv9W+kYwcWX9kdWEC3pyxDoxCG0LntiAFDArF2x97Ue1++PH
16owZGoBwlkBBEY1kCwYSN82thv2lYxZvCWC/6KLOpq/1GdaJ3rlfBpLL1gCrjbW
LE7LXHpv7CMS1F6Le72BUHYH2K3q39Tsii1nSsrs1SgM7cyVfZKv5EoUC60r63Jy
3cZYH7+mIHdvI6bt71WKltzOHKyPt6cl2hfWKQug/Oifk8VUQwtEEw4DQEmNyud0
lcYjuaa/5hAIglSFiGxkPGcVuMekE/iz5zclk6uw+/o56aAWooyTVaJz8VrnzY+v
69OHX0k9ROhQFku+SumfE1vRtb4dSwv8vRn3gGB8ZdtBXNvjuwvDSdxehjSSM7KQ
+B28HQ7CaQAZuz2K/O/UuRMhuxbi+YKQAabGUOHGOVG4EE/NyRff+OBnLtq2Mw3Q
m6XtEl2j/a9vNmFNHZ6QvubuxVCWtdOfyYsYJDrUTVoDVZaRF4N9MEQlN6l+/ZRm
mfJC9vI9aRuaP0pqz25DPZi7i6wZdA/UOiMiv0cGFtEwZPy+tPGjxyjsjKgYpTVq
269PINgWSR0QvlTYeNE+Her8/ZDY/9y9Hux+LmIevE6iHUlQCeGByUmblKEn7edJ
s0FLPdS9srZjyruClrI1nIbuOpzCkNTOqfAmCtRuAcfJYbny5z7sggT5ED5zsqQA
HgwgcxmvJNQO5mzJequtGoVHTU2EnYu8TDgScKkb2WmC0fOZ8aIlEQrHgBjMbqB5
vQg97jb6rFqsJ6MTEU/Hx691Osmb2oH3B5lNDkG4ozuvE+EyKEFIgCFmhzSesW2H
xpkzwxZqdXF5Vl5OdSj4a4gxFp4HGBSvcpDW3Q1G+qFsXAHiOju1mpuPvWpeA08U
tBk9bZi8tIEjJ1fGmlh+PZbjJL6LkGxb0Wd7B1RB3dtFWHwNcL4U184zPV1sTszR
LibeMyrFh2362/Xg1NJh+Ksh+Vl/3nKaRgyTIeu7zjLd6H344R2/JN7VcN1CCXcP
81WzzaK1o3fPPsp7wI0FRagkM1byHVMEvbaaxQeqWDt3hsQbcfeek2+ujDJ/2Nud
8I04GLKq2SKmiaNQEst6bvX2zosy0JBwtNuJZk1LuVYWXwnAqZ4PliyC33zirEAU
fPzMroEjBYykhq3xefOf8uTaX9O7xGAfegIjyg+UUBZWMgeE+9wqSYYPlvsObg+3
FiHfHzaJWSC4K/hgktc7zlvB7OwlXorMk5OFXBscE1xlcDOIxkY/6QcniJtgXUb3
uOTRekj68EQgO9kwrd/l8TyldxCcllueCEFw3KDQZq3Pvdjm4cN22npgw05yGw3k
ETZfGklZ5twiEnkjwYqOcIkaJ4l1JX3DE+j0FdSqYayV70qn4DmkNG/PpXUT/Z0j
/zecvKYUpwSci/QGAant1fG9Em4fU07uSVXkw3UCsHVSar3IIX8qbvTsWV3kqSWt
5Sem8umv9AttzupJ8DcYGg2zabPcOB/CQ1iJfeoaOiu+M/Jwj+0n5pebUZJFl+fp
KQkXk9SsKJtf49jtvfa1GKGzhZcgifVqIojZlkYPp64n8vb8n5mjpMES4rmWxCSC
ofD4/k7uzBQQdrvuW6NazuRnTJ6x7zqmFvnAI0IQ2S6nBcLVET+RXqRf3vRPg+GC
Uimwz9rK4Z8LHU8XCm+X0dsVFrMNlEUWoD83/9ee6avMI3IOyEnmJeLphHHMZVua
5O+zg8Zrp7FGZORjS+j9WFX63UHs6FVgvf606g0V9U6b/CmjMF2egaWjshiw2MUj
sGw4ZRAIRXAVc3UomtXQ3/qqsVbUtb7OEtwyT5TqT9fy4yxrJhYHyPHrzkXAzRpY
FuxhGutpIeRWAQDjC5Jecf0rGOnv747f3Q10v0BszRC08/I1+JJeJB99ftu7BSfF
CYIDty9sGzPZx74O4GKG9PHJLnlvnMG08nefhLLsdPpQ36EIFIc2gHp8hSdbuvh7
`protect END_PROTECTED
