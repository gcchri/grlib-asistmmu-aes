`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U52XgHdFVoS0IWNRTIDhvqyB/Fr94s+9uXa9FXRtwNvBtJOGI4/zVaauyhmULHGU
ftM2E1lu7E03NHjc+GW7DqZJnfmH2kYko0yH6QIutSUiwWDMRa2Q/3rxe8SQailz
e6XaV9b7hMGQoJEd8uTVzJDCA3Anzfd65NrDqNmf6mnMNK8b7Aiui8LtQMTilFcZ
19P1WfByYOCD/Ippgj8c+u7Sk//NP0BbPufDZP+4zKlzdsl67IWyR/raxeRsZssr
E7ACHFXkHSsFTZHlQhwhTg==
`protect END_PROTECTED
