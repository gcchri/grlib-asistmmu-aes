`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JuPWIYjxaoszzPLst60laFZzg4gbbLnsF9BzBkJdtA6BOEprJ38C1XMInufchn1C
wywuVqovzYrrmh8DwV/TtGwvDsyQagqHY08uIAlK/Fk1AsNZnTDU7pxM/vbIBn7k
LfHR/Xy5rLDROtkrv4PyYm/yn7XpsmdXorqqen4S4RBdqcMgt3QXbGZkwstZli4t
m0o3hxvxdANx3cUC2y4c8hwBJse0bw8i8egxPhGRztXRB9mFbFy9eic9pxAZ1Kns
x7WAv3SC2eQQt0zhybrbbME+Oglm1xVVyRgM30p32whbpWp1NtrIX6HLioPEWlZH
dhx2rFnFT2Uqf86AmqcHL1Gt+aeRoK/+JhDGashaDWoF+60wsrLkXXDcZLNpgPqQ
0gwvZy1Ij7SPzwhjLlBlTVmBHICi3wdUn9VrSXpge4mngncn/5vhRw4s3sLImCtN
8MZYHDvcIIMiW50qSblWNWTJ2OBu/kKmMik3/w0nCjYWKTfC78VvEZY58CIrDi5A
4QK3br3NoEDLKzAUdR4gXohsc5T8iWTRNtUKgUcBicwB8wTs3Ebvkl4ZKB8elyTg
7vZWVX7e+2RkOW54FGpWDJ4UFkzmxT2sp368Z+RCPfjcRc+GXVX9YUXFRMcZb5PD
T2DGnhtvI9XYVraG68LEAvAW8UJOiGlwj6uV+iSgqyNkdiuoLs2jVRGyUuY2L5Ml
G/FbPZJjJ7+bGWMUjPz7yO5zPK50ZwJ3bGYJD08NyTsEc4/BLaudy0lHYafAAP06
KumFhDyAHV10xmtIHQ8CnOzE47katdxRY6jITU5xd8psWfBLZ3dNpJNcn9VXNK/g
uoCOqZCJLcdhzJlZLSVTvBD7iZTX//s1u7//hl4GOc9C77tC0jWUCmT2SHkws6HS
9VFfmE1hKQS0iu5hYY3Q7rAhH0Bmnooda1b9AaKAF56v6dcGDH61QfVJgIuZwTk3
If8o9nL318Ph2b9lq2D+FCx5bifI1Utts3/1nS07M4khHYjoS3yJqHWpX/bRBe3k
+c86Nb6RmlvjIVz0Egiu47VfcumTa91b4MKfL/njscA14zLM9RZwAqEL/iBBJVF/
hZd1778EYbyDr7bS3bL7c8QFdF7GwRsWYN7zuUxpxniM57qC7XGKvVrAFFiDQ4kA
+U/+3xolGmHSxP3phN0C4GsovB0yaQ+Aa30/+wg7cgJ8X+z72lGyT/NTSWQ7hooD
w54L/gczQmKZM3iEVe+XCdtd4FEjLd7eTl5lqafafMl0o6KAlK3VycvF9FqjN5UR
jhPIrLthaeluivGt7VVOK8y2RnTwjvzLaPLXLICHLzyyLBt12pCZ5jfm6kWKjE9M
pnueeLpkxL3z61f4+HJybw/6EXaFHXVC14rwku9l0rFwBpXjijoTyiDtUObQDAsp
ntGtOj0LI5Xz1syYSwB3dylLmQhPCf6siUFsCD0mE2Esveo+2308q6/62nY/Y4qt
OW9TeHoWOPtq6Rd/QQwpNjm+cAzy80ifVbsQ5o8soKBrssJgss+8/L9i07AgyZCv
XlxQhqXlr64aTWIkjtD4aASLxqt0289fzfxiU7PYkJB7GqAEu8vjj4k1N16WuzLj
3DyQheHjtWBBC80zNoMiyZg0zQMKL99UQ0edUwCy1ojTdGFQWAagRKW87rbBUQst
Uz7MI1QfRuPYlwo0CNbRRCuQwfQz0B9Zx5R/FNb74QUwBuzF+eoMaphCYi6dczZH
Ts4NHXrHDxeTWM1Caze4rSBZHiaFOEsWpQ9XrbXl9a5wUA16GgkNPGIcR2khA11N
6rYstD1GFBleOV1P5LH+K5wuEZoem6gPKQjSiQLR3+SV/v7eG88M4JNA3U+FXnNk
i+T0jW//MBgzgXcNQis35a2+vHu8G+NQEPC1QDQJNGG2Tevd6gSn5jHRvsXrdlVk
pRYUcc90iT1GBMrewsDTTjbVoc4E+kbWXAapBbmkHxrUhJ0HNFpGurB/ZAFoSK1+
rdgcpFY0pH7zKp03Sgn1KyQJUawAjDRJx28yOivvVpc/J7b6E1i9b11ksyNZ8ZSZ
oPPS8TOMth6h+6Ts/RtgO99qJNFq85L0DkG83UC7D6jk+X0mbDEXJS098AsiNC/Y
lWlHD9OCDQvpsvG5IwwiVcPlpg3CkC88Rz9zbkv8nSz1GxuFEokoSf0dqaTd8wiV
CmWLQaqjzcSiOxcyQJitKo3I4dAQIKq0fmBuyJOuh8vgejERtqnuygExCXWxwR/N
PjQxPU2zkjiB1d7ikTGbsG6pgA22K8fsXJfQZY2CZelEABXrBdRt/4Q2kUzArNoJ
Kl9rOYQvYgzqsGPsnTEA+krEIEWLmvZ9iTHQEt7cm8hLzhO/U4I28kI6E64gL/4i
Eo4hDZShuO7+FM1QMH1HdOTUvXKVajrh2XJhAypKAdxI2YwIgMaQx/kqvCimqyjh
5GDn2ZxQgFkIh6UJwxa59xzwMxABvGG5d+expQlxsIkKlPFoW2M/GEvsBPy2nE5v
Et3ijka2lx47OhXRVOL0AkLMEwSldEd0tz6tiQXX2wP3WMuvpecuu/icKklA3vqX
XF1/LJozVrW1NESUU9CNFaf+qGJQZu9xlwhFPJQVENvTqvJb3gETkgiHI8Av/peQ
QQ4xx5jYC+Ob3EUlptfmLkhXduypCMVGzuSUhpr6mbPsrRTin78yNlrJfM7wL83j
`protect END_PROTECTED
