`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XCgEbbC4IeKJ4MHpcqtAhaBlmHUh1ejAtVPlyaFtV7FZMDtNS+CL82yJVovgTl8
GNNTJ1iiXqGob3FSeHEt0h8dpxYBXxz+0vkG7t4T4gsPFbcPGAvGwVnvkNUAefFM
eCb0drPF2fWWHSHhy8ayiJIZeZ0ELAIU8MrSvlC2emoalAfPUa/7W+0iYH8eNksL
u6uZGt5vCK2gm7zeUC6aNA1SxCAfOqW8QNzD6U1V9Jt+90UvJe/oS2UcdjpsNJuA
2WCEP54yVVRFFRChInJD2aAiHrOt2jfzlb2N/93R9BUhl5YAcF13df1oSn1KVkkG
S74i4nWo46JJTya2ye76qZYQVzwvVv4fgjSwUYG4f2Z7ftj/kEiwh1VnEmTAkDE2
k1GXcIzwmFVlhwgSUhAlg1Uh433Kc4DS8I8/11i32IHq5w3v/Y/XNktTQNX/ZwTZ
+s0jGWQH5O5qq0c4SXzm2g+aRfZjQmoLTXFiNdtJW19PpXlMfTSL0LNWVwh8h3Zh
0hPUbwM/yAsLegmYZ612Hakcku6n9DRUcb/bws1JO1jGwF2TfvqTxi3nuYPFjX/j
iOHrKP+ARsVIyrw0DzwqxrhiJuETcB5i4RhsJpywaEYE7Gm+wk8RqmfFSqnqcKQD
leuNr1maYUMTL1GBP0bJt3ISUg1LLF+JLYbT7p615pokM4c23S8rLd2vTn/GihJV
0bvU5dB5sQlU7dOgYuLijf7ZoLPsnA0i4E+zNAEqZLRRNgs7LDYY5cP37RVDdm2E
n10fx8+z88KpxCMm/aH4DMPf6omqENst3w0+dPZz73FHDoM8WpTOUA+ohqj4LDHu
IFqSfi55VCtXVV0AOhI43CptB8IucaluMf69FcDKojeJbUzuLfX/pepNbZxFJdZc
aAGsD1lTPOzKzDHGoPWaJNexH5KtERs45kCcK37MX7P1uVGTpPdsz6a/Gm4zmj6S
r+k0FZP+VvYguGoxWsOGhdcDFcWg3nff1fo8+jDH/RxrgjwE4m8q/UZIiI37TsLQ
FG63lZ0CK7Fx7uq73NjWEbHKO66/5+Z754TTgvkV2YfhOjSRkvsfcuzE6DPs0LiV
iCTIOf1/IjineQF515Mq4FkXARn/EFQKRQc4pkROrvo+g7Up6AE4n1CVIlKkmxQD
8kv353LAGnsWteqkUtJ3Wktpi53kS1x4vGszWg9QsMCSvkaTrR+1W/0QWk8tHwhA
cjVF148xw4yolnGkuli+Ey/h2ZdMWub0/1cwhGob4VOnzzGcuC+a9wN5HnmdcDRT
kkWuAzDza1vsOQOcQiWtRjUzy9KWES/3TycbXKDVbxR1KgZMurZ8ejFMbmJkMK2r
HBMdppzLM6a3PC/hGonUFOz4T9AwiBljiq+yiY//PYaYGT0LnUvcmGabWrP5/ZLm
udXnsyTVA4j7OytUr6AMIxR8Z4QDSoe0K48XjuET19YQtb9Db2FfM368wWlytF1k
uC8C/9DmOkP1hYn2r9vU7bmm62UMu+90OisiGBi9NK2XLJqrTLvrJnCp8Kt8XSNw
tGCh3pXckevDyXYw/SxnZ36XZxqj/uAmtCRtA3OesREqPBrVnbgSB+hpQOr6xu4r
VlCBinjDofMYBD8XBvVRcJtKjBc34lSk6Symy6FbBxpPG14RbdruVjuPPU/7LY9O
7ZXklumKSa0wg7BjEKWxmgmiXohJHnkzIcA1famoBSpXDEwPasN2WtsH8oKbdcZm
ZSWYuoaWFfph95wGEr3uQsW5RBnHLkzmVw6qn2UFM5i8yPMkwwS6PHNOeeOVCqzc
W66Qw8g5agHJGDK5zmqX53kxaUJxhdvN53VAkkkpZwF8tq521Y3aUpps5cT8JKow
k8gvuELGI/68vunrq7n1QiNn6Ql46Ans29yGxoYrIhZzJSyOx+Y9x6LZTYEBoCFl
Q3JdgIDe93MPELEaGxirKon2bL3z8+DtJRYoloMWtPDt8d2ktxOmbZl0K1iouLY+
kxPI+iDjJRQZfZBhshPYiXn5dXYOrJR6QQA+qkcGDf1+p6eFAWTk9raDXtsIvB5E
QKsDtJY52cGuTjsdbD+7MN+ozh6C4b4KrRWd0w3yb0mjf64VNMyQ2ouWEMdqWqA1
wXqUtyaoSdftms+O3hkIgw6IajSLzIcMB2ALgPvFfbhT+Jqg9K+roXYABaoAc4Ox
03vWDVfqwOu9kLjzEqojYukvhTAXkXIKpDvlg2NVsLA65p5r9IoZNodBaoysxj3C
ku+OEA/37nQVQ8r3zwtoMDIEd/Dp+R1NgSyOm4qinAPzk8h++s51T/7ZNEun9rhS
EsiNIOPhZEUTjlLdWL4770lcGac+cFPx14IbwPrw10CRci22Dv/0yZz66M3mb3Jm
6zEjHK8Cx8/IBsc9UOBbsZstAaFR/W6yamm71C/dAbZB4lgL58CiKD3uAaEaeTS8
tCr6iLcAwcHEEpSf//o0iGw7DrF00gIwP2jeWxtoDApNdZ1OCErzeoddIhUs0zoI
ufcoPnj1tx+2lk9BrTl6tYQjnS7geph6wQCWbjqeaBkcu+fMYyBkK2gC0jMcup1V
v7JFA784OXmzrlDDcVsl6aFULVGYNOJSAbmPvsm1Neids974ZTRzilpJYNvEPt1j
VwgRznXNMbRtz6i/Tg0GgcQjHzQhI940tp2R7TGbVqPqf1xaWsHO8sBjj2VLVW7I
iEKCxXN7ncL1izvIFb7L/vDGs5ZQNS+0MwJDzeC/5w9hmaQ9AutwwT73BtwPhijX
ijHxTi3jEJwjsi3mCgWJQsBv5NeFmp6iXvelAIw/dOVLYfA85WPD87fKbPVFoC+N
CQFUD0vB944sQyZdcXcYmNRXh+8Ad+SrwIIunrEZKPyFMrs8lQfWm4kaRr75Xy5Z
ylVyWVzoPnOgLkzdOE03euchNXXBQe6X+c6uWOCpPdR9m4F9LsPm3ZpH+iBvQL9f
Z4hFMvHG3D6ZI9x6/5p8axq3vGOhV9EKXhsiLSY2r68MLzjcew3DMko8fRs9Jgns
mSur+E1NZjG9dPAO5OkyoERI+knQRh4DSYAi9fPXm+qpEGrPzy/jXfsni6R0FQmn
ertMw9AimsKhTuhJF2evXnbE4pqo9p4Qhto0yqtsZaCvHXaROn9m14yQjZduFxGT
IBhH8M5QS37w0R4pWNfHlpb9ec0DbYca1B5sef6go8N597I6jMLtz2/6Zx0TwEjD
y/Ngj0slI3tvWIMVzs9ZoBzZAfrwU+ysxJDuUS/X+pnkFA8igif1hlK6pLr0hOHO
/faybdvNx3nCab/FEBRrHGu1euWuc88BcI7r389yAUM0tw5VPN6Qd4n/iPEJMFkk
GiLToKDvqZ5S0toJxd45jbjWkdcSH1N6ejHZcACdQSswoN8cX+5e1aUGTI/+vH3i
/Cyb8BEoRvPKzHzFsFgBrAZgDh7muhEzX/G0ezEsZQRywnXiDojZBf69m3mo8MWt
HPQjWbU8ctmfQSc9vD7oSy58qjfPU9J9y/a6F8UlL0OvEZJBXny3uM/EER4Wlzy3
4VTrBpHl3yhhk2+01R8Hty5YXhs5KY6rVG5NQInvzHF239/Ojbcx2fW2xyiamvV0
+8/FxOa0Lu4Za/OYf4SM9Faxk+aKoaWvFfdmFbGa9SiA+3I5sBq3UK8KtVnxcUYg
rUrCI0NO+OYel4qrVC/stJgH8fVu9MQFd/VkCbiDHkTaJ5AmefbF+UIUREFupBVg
+j3tOp1h4aU7pONHu8CsG9XlyUS/9HSMWaWV1J/4+k/arWS+HUsmRY7crf6xWw4R
DvtGSiKpCsMptobiL3K3CgpDL1KlfoLVX/QoAANtwwxhtsy3pEGZdxNoIO16UOV7
UA41SPkWYB0O/Aj70h0Fv7vNQu26/KE3+ZTKg1NkGeTjH0fG/3ymuq7ABMUygL+R
mnUYdu1qqfoNhOCvO9Ed5mfD3WcHnOqlGJFbT3sK4nt7b8tOzuN1D10BTXm4ohXi
hMNQclH/a6XRKF8we+6k5l+g47Kj6SBVWlbazf8ftK1C++D5TuwkhPkwm/+JeJ1F
kh0WJNb7fbbVgnDiAZlFjDqbkmlY7ZEoxi2jEYcIjx6gDrbzMD8sH2W/3lSXjkz/
o6UdIUEjosQiUY6G5AqOEFYf/8oqxJFB/OzrphvVbTX/fqT9qh6nfjw+KgIxJu2+
uv4ei310pVtxrqo1nnkllRfX6NLlZEMC0NGQTgIIViOLLbw8m0rNeEZit9UuBLgq
9n7owN4sNWAnpHuGAlyJnNe5A8fUc9IRlY6rMbP5sq7wtu/d+VIRsKtRkgkA9I6X
wkgcmvU4CDCOcJz7QjaSazWPVN1TpodPuzoWDAPiS/4i/8dtN5SLuc+ybTFRfq7Q
WF1rImaPGj4ImoD7vaN8h990cfX2NI2rqlUm48W72Rj9367q/67F6ixRIH/gaIaB
xyAUSWJC6z88Jd0EMCTubU5Y7WXeXmKEA1+NgfNF+VH40cBc8OYC0kQ0BBKiZ+H6
jKsEtAmK3UTx0uFROiRnzg==
`protect END_PROTECTED
