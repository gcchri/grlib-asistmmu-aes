`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zth+Tarfgo8WFHaDg65KJBoe0jkWz9NIg8pr/cMNrfghs/acDQj6GNrQ1BDiaqwA
8fgtZpx4CaCTRv8JIcB0P+GrAeXPGk50V9FtIIvyWKYTIoI6LzEj+Rk4qOISWU6z
ackjnqWH1p7GXqaVhKYHd5m4PYP845+X5JvG4N/OgQSqFNtRFMIyvrZp0SAQ4jqT
OSA3mlnd60veSJ8kzDB7uJgWlXEYnt4bpo1mD0qjErdP81UDoqK0nR4gMd1PAJwL
3/zUcCKyl0/APGRAz4zC8W0RvW5Oda9rjYEeGI6PTOC06ET1wncK3xdnAj3QmSNi
ECDYQX8KrS8YbmBUio6OALMp7OW6I32fBOhoSVhJUtHeF6jI5f2YbVu/0WE+cAO7
JzBSrgCryse+WLVNLWH339loyKve8i4uw1VkjQCjsz5oSxnQPcr5kIvwxvRXmoSD
KQ/08sumXTcqWo6vZ69SxAK1WAGHfgoi18G2PFSPEuHIWU/ENmxXaWqKwVytgOEX
2qESDhIlg4MIi3N8pnetH7jKnPw2Oo+TY6zqPS1I8hP8X7VXFEyb3bh5+7swVHep
4EpqK/isNEPj7Kl2UvFmRLpTz3xmy9K3TPUHIqH0Musp9YQMy1eGwXRXDvMf46XG
aoQZSJRf+05ECM5ez0+WEBg7LtY/eEtRmVv5tu06Mz2elXO1cHIKu+zkrRSA53aJ
gp1XBSVn9ONtugs05RepyU8AoPhwtgXQztcb/fcl9Tc=
`protect END_PROTECTED
