`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iyVcnZJR+DCGYN4O/jYymPW5zIz8WItqQg+Z0dMPnGnH8fIwqSmd9H3P7+gJ0YPo
c4mTLWEwXNnIzkcSvDvU87lIICJlfqIByjdYlXgt8lvatSQP5997QkMg7DwIFfqe
uIwOMzu11U5GQ7I8aQWhqQ1jT3rVfbjZMC5p6gYvWarKwpPBZlEZa5YFboQYYdVc
ki7PB0z92mJUE00KcfCSlFH7SdYCgooVoKiY0IpZYC1bqlTjMfnSBKsLEKrEBirc
VzT9ikGz6lqYP9boKdCbLMEl/Yly3/hMCTAQiQ6W3XfZ2KqchmCyK5IsEuLgMqc6
esGeOppvqut/jDQBDN6Cop6LwKZJg/bC/ji4+w3P2qJkM8pXY1nGcylMoJCoZ+zN
9ODkhkEsbP1ltr3VrD74L/AP9+i+vX+ZvSw96jAiZn2j4EA7vAivnT0KdQmnBktt
CvYIYAuXTeZOBU45u0RJghGXZ17Rpl+ZdUFiWz5OY2gzYMd0KRGFTHxtjJ9igAi3
enz/wnSRBjZjKSR/5L9qEDkB5O2o7w9RXjch75ecTytrNBFP0HB2thq1MGAqeS0Z
`protect END_PROTECTED
