`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
adNg2p+kcblKL4YVqJEw1UarPYq9S932QHwkOPEyKAVqfQ4dV9HRA0NlC2eTIY0r
uLMmEd+O14IibBeYsQzHYdzXoKMbxTXkXjiZCeDHdH4ZKB09jU6EcM/heMo3+Hkc
yI1SHKhj+qJ/BahiLHnGpqLyJSdBgQN8myL19tPuAjyZUP3741uZpOVk041YSkZJ
INfQmXQfMhc+LKOTkO8kJcZc4tSNdxnMz6amUoap3DDJ1KeZCBXrJKdeNYu42K/6
nAGu448klRpchVjd9nbVpw==
`protect END_PROTECTED
