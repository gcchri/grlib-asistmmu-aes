`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4bnumKeMw0IHfufZnxp+m907L9YuMaczb01RTaXqBMsyqHlRNXQQhSUZGKjyabK
qkQiZSr/JgPfL9DtvJZVXpAglkwyNU3M2VcdQVYUgrJ/FbxGgbzr+00o54z8kb2V
JWijPW/UFQHomLOw8MTMAyGzxqJBGBGYgXzvXyTbGoPwCwWZnl3bQxzDTJUvZ9oL
yXEqTdXva7ulfBSJweIJNbpGvB6D8cWLvuRnwOLXY3BxA4uXBPVN88lqFSD0rYpB
yObB6NSTYQWpU+1+8DR+oa7KcrCxMLV1ikygINhE2UwlVjv47pu8VmzzdLJPftGW
t29wEk1pepS3lTXcUPq7Aj1eqM+kO9trhl52MUtY2a8nn8wzEJUwffm/2PKAczEl
VK5Q5BppgYPigBX2SqebE1VnMoYF+KmFdZMJk0eXWWBjxFGGYavkZywnuIfe99DJ
zCm4SF4zrdtesEDl4i78UrvNsrwuMy8jmDqw9Qrqq1VWsMm72PVLDAUAJ+SmovtG
xs1WdZ2FcirhQUUnSD79gfAJLpTZTGbDPKX4HMLN+6wDtEfhu6I41KKijxTO1n3W
WapyehP0LC6Ulf2A9HAJAKY+eVfj9jXUHFFacxk7qx1xl3ucIg6McM7pdeMdDUgq
3vHa9MvGgWbZHhnxJJz4nG8jzJTX4GjqZHN37xFff9A=
`protect END_PROTECTED
