`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Goby9WMd6NBkd+z029iC66dytCVD8nYvogpeqKh1nEs0PpukwRZK8+DbUa0Fupi0
rIAFO48B0/XhYipeyMNyiQdcJxpFGdIPNNSktPPYYnuvUkk9L+gh/y574TXhGEzI
0kUZCMSJItRZQCVO8EKLs1rDuwkn0gHy56sX2Frgy6GgdPAHXZO1gg1iwFeoI6a4
KWtHYG5BTQxTYKNGcDVayYg7/bj+QOlQUmxuZV8i/1v8tETotMJHSqq2y0ni6zlr
bA2xW1SmXPDeYDjGeZtYk3/PYWeaxCNQ8zwP3DoltTpc40n5UxyCi1EWk12LGdY1
NxYxGXCsHRoJfsCsqS6aUdopfZgmJO499Lq3Dlw8SnKsKzQimvvYS2AwOuH/XUc8
ntSPE+um+riypX3GuwnL/0jRDkYX92pzCWe/rfzWfYMZ7F5bl3ZNoZvebTb991MV
dx4tlyM9uvJthNg38fxEE2ILE3SR2ifRPBN/0+1qyVulNViBEd0jAx4TqZ9gP4jF
CYbUdgOP9EHGyCtPvXfzFwhvriML5eZtdf1HsOoFoFLzy1ZvWOTqB5Cw22BvAE9x
JRooSwAV5yQPZgyNxcFdKgcAskT5VFLV/MQ/dTMDJZptcKHWQqe1gNisLpwJPiVr
D+In3TUyZnK/CdttLPP5LCruge8ABvhKiaWzxcukR3yvXdaiEgsI+ZnBol1myeWC
v/XmzDbPiIn1xgX/Xg6hktIKUF2L/u+qa3DSLXQDeKzOtc8yQFvd8iNIFRS+FRyw
ocBjiBMUMfvWssGPS79kyqYY4z1Tx4W1ieTBuVNvWdPRR2A9wYOQgGgTSuZ4YwdM
Vs5wmgvYSoZPBM+h3eWPLyvtsmSUZ/KYM8fJyJDwSFII4JyZ6wTw+X+eIxZBaDcl
GA98t7X0DNPpBt7Jaf5zCZuONMvrq4v8pfPcF9NggrefVSyZXm+xDn4E1NdHyvXy
qVJlHuzoi9lS3T1R4ufhja12bMHziZmfJ+sPnrEvfv2Lcjh+BurVYfZwjsfO1rcJ
RUWTVae9x30NmQ0wIsUreRpXENS/RQmpP54fYOYlVLa6EHma68OMjCoet2U1altX
soxuGQijrmD8GSsk70swVJeI7uIBLdk+8FupfJxOpZKEoQk8EB36ZryW912nRF/B
lBYu0gp7ZcE46gs+1v+6Y9GpM3YEA2BhuOnLH/u/Gr8Nc+5bSBSBi6D/OZp02JDG
eOczgTVvT1NIb6C5kZm6a3sFady/h41r0e/ezl2R/VslFJmRAPfZ0i0pQlk9Rwee
s03mSk7GnoSIuAO3F7a/daMUpV0vzbabnzEqf66wkDTM0Yg4uZqT1KEPSdx+Hc0q
9PtqPBSyBLQLANgZe7VuRmjuX1/Mbfe35lYzrrw4Bf6WgCPKNiMoFlAarey4md0N
ou/0WCAT4iMObCi6aqdJwww9gvlVU81wtcXE+UhCcAF3Eh5HUOeZnm9+0dxHQm5Z
ohK9L4Dqnm+PTMReHrKtVyBR08UOjYQIR/NWVRYsJQCy+IQ4ypK81Wtu4EZ1eSfJ
8L224LiBnWXedtfhuddEqTYosJRy/KD4epRc3OANO1msPkUaknTFMVyLjGZzvtz0
1s8IEKMieHnuCfm6Oc2NZkFhtwqK1afjlrhmmTPHfXoBz+hQ+ObKO5RCq2BXmQjX
1MfRNKbDTe3mxGEdEH/w3U8T3KQ4mxMsi2WXph/U7fFKSS5UpTIiHUWlCnGJPXdH
GVVleBrvEznbZBpccweBAXgDgj8enVljCFyjmQmVXOMJywrJCKcoYdNCbKodw0J2
qEr7OpV1ahFU8DtUZZjuXpTyu8x+iVc1gNglzFOw1dQdGR2VwkYkBbA1EMuKzV6q
v6u37iuVhQVg+j1vpYAyH2Jkcfxz973qQVZ7NCm9buhbrXCqm+4HdnqjzhMvqpt6
ghm5jJu3yJkAk/tfCMKvF9ZoE2OUjp+3fn0fEEytRLosp4+fM7DeyAvyjAXYig3F
3d7CnWan2tpszPW8HtC7MOadHtescMXyESU7uveqbEBuhbh4/DFLl0RkrVB9DS7C
cur7JKiRjJ5C/rqZRUsZUToI9vrcIlhhPlHZh+4U8iic+bOn/Sy1B24aEWUqOO5F
+3sqzxbUFCCtxYXZb++UCuhVN+I4Nnu9OXybS4uhH4iBYPjAHP7C9TzY1uELw9r/
cvdrTlGfYgEzriFgv7/Z4bmoA02uaK5X9IDGhpKUvDw9n3eQyFFZPNrNvgz8wY71
TPBgwRyQlcrnUZ/IKERq+aUntBHs2Kv+/6Pg4ylI9hgYiugyhnWFDW7Ynkg9RNGx
LWANBtMvYjX+z3BApsjDuN8RsBQDyUI4LVRg0Vj4F21XPkvU9cbd/f7n1/wvDGEF
mg+Ax7vYvtonZPcF2Rt+DZiAvg4B2N9Dv0AK3IjFF+QMYMzQKjY44rVBfIsQPNF9
9ewsH07isdimu03jyHD1+v8OKC0SATYHi2yYB19R0tQbrV/fRICuUPNSDY9BKZtu
TO86dhK7Ih1mG/kWbBT/AeiYL+AOi96pk1TVIaLlyJKhJgkQ025rztGyjA26fMl0
56CuIAhtZLsaM8aQYEm1PveOC2v3eEH3MTaiIIxXts7zNHESo7gKhNsxPtfJ4uUQ
SfU+QdJqxdAiSh8XhLHubuNhTVwbqWzOCrXKYbiV9ZU=
`protect END_PROTECTED
