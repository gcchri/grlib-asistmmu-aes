`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5i6oFZZvgU8fP/JOjSo1g3pdrr+JclpgMVMsgyB9OuhpO8VXjzWhPHPp7CLkETx0
2yWl4eEZCrgu3ignyqLZcpMthGMIsNkmogisVxlej9SjFs/A0J4MXq9SBikYdUtP
g6NPQoHbaawntBncOZYguZuGELlReXcUftsaJGprm1TckPZcHEQTtMq+ymWmtFCO
Uwp56zR3N6h7wNW7v8Y3zi7OLuojIFNe9ImUNNqg4SaGl3emuSAV2hiBiTQ3eO/X
7OUB6K3QlngZjxuwnlZlvwFFGKcfF3Ch84q6QLaHgrN4lTrqZ/Sd1sFj6PhEaBGJ
oqyIn30iWEY2ejLURWQ8/DtVvMsZrwG8OicinfnhZXYy/+jC9TvBSxJ74AiUSke2
N0IN4MYYEeXDUHuCUrmQ4a1lgUJk8DmL9lhq1GUDPhxebShF4lQ0xO66pvkdzXNm
S8NE4+0D4u69y5en2aVjEeFx6I3VDCKBsW7WdZyZV4agnEG2b4sPyyQLX+84m96p
f0JvR7Jc9DUUYPM0RpIj3mKIY6i7RL2HAiaVsK+8limvDnGUDN54AX/Cn6hjnihh
r6CMuEHR7JZNITyEahiN7BMPyRzH1fnwpnrrvEY2cmDOJ4POuWHFW1yTBSTNbyqK
TXV8oewsefgAqcuL0ItNxCMnhWWf0P94UUg0ZAoMrMJq227Jk3BY5Qo+TFnC0Ie5
WznH1LOO2l7xOfAg657fKBiBoQUs80vQtdUkbkK+b0Ri7nIV9504jU/COxV7ZkO/
8UZ1Dl6BdvXgAtJCBjSYOO+8gQqk+gliiCHtEjnIgwnW6rnbScWqa/DGy4EXQSLG
QS5buWjVAXr1k+kEZ7AWnlympDWR64N+FQoyuiTPaCc=
`protect END_PROTECTED
