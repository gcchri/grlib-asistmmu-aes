`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0wJNanR2VQ7L88TfG2jwYs8f8D7sFJOTPYN9gKEHG4G07mjRpmlBYbEjUZ5iSMuV
HUgsTPrGW9Ry+bwVoN1aM0JWo3013Ifwj0VWDB+oLlIaiXpNYeOanrZ+svVbNkmj
H6xB5qHS4UzovF/4GNyDizjziDc26dJht8II4JqCSGBbVDErzZ0WCAspudUEzAHY
p0UZiOf58wRqzelZXvsxgvYKmTaEJ4kPRNNA9CdJO18VXssHFiEZEpuKp0zYPK8b
AqPhOxwgpfKwGcHRcseN/oErzr1XQrfEvydNPc2FhzFqynZ5J0C5/VuDMw2Us9WA
GWu3WB06wb84RAbRulHv86RjbVMKI/R7qh1oQQVoQP7wiS0nHl241zgorJzVVnEZ
EP3MpWx0d7atxPWvPOXpz8R0xvAGNefjvA9BRVyPCV5ptLoQBRjyByhvQoivNGdt
WQBEOrxhTDewMSMNW+6pYd+zKmVIRpoxpJdVTnRYgc94GU0IQoQZYs+vAJrsAbzU
uApPoeGtLZmgcnQ0kRO0B7b6qtxJIm+vZHQDL+gm+ClWyTbnBwNqokgtz8v5mcZu
z+OwJ01AcXoH7L3GNqPlkRxcQJDoqBejVyNmnrhaC88rOl7zBsbjano3gEt52Dg5
x2VR5QHkx/s0ZHVqXxALDZeFcXLLVWlf/iXgVcDN6+s3QRL2r53+2sWCvYzmWHi1
BQXYJUDbrRMfqpxZuhHAnMBKH87XiLZ3OeRxEzVsGes/cl5y5UaS0oAGS5rUIU1P
zxfAE2I7ZznqyhvtaHnqNCQDPJNjK43XifLNYl/WeiqER0LY5C2x2uzmx5iEfbn7
11L70/S/XYUS1RGDCp+Zk+iQ1nH5iINUpKdjboIU08T5zOFqD3h+E4jorMK02Mbh
vIn1Ipj4otrBdqbyLZK9vf7wZzJcIRlFSu2VJ85E0HZkbI9FCSBJEjFl7fuMXJB5
n7c3BlRXbO/9T9feP+6Kw+btBsM2SLG6YHDBfUQEM3xFHerOvvFvaydi5MXzvIq9
+azTyqLpZzL8g95M6eBF5TmLd7LhPfcsyK8pW2WqUkVQ9fTNJ6gNvgsWhItxfw4C
X6RZ+YdNC+Ak7stbqTAvD2s7kFWyE71C5kyPLvWeOOa3TosGDneNQNM2qtdsUCHr
F/HH3DKXEOa2SEL/Db3h7+u8jfsCy0poL/4CTDmSOyxWjl380vWkbvGUGmjawPoP
YdX/BSBzSHzmfyamGhEo1Bl1BEyb2g4pWxRlqFZIGrwKya6BLwp7B0diT7CwYR3a
dxpXnnsFQsWT3RHYzpS1i420MZlT3qbhia4mN/K/t8InNfQRIO75v5PDAwg4ccfR
AtDEVaQsIbNjlUYTL8HMW4EwZiVDTIgL1rZ3HugKKY9XsCHsHvK0HeZ6GYVKWG3U
RddSSTzuS5wojkUK0vVYlxZrb1L9TIbdT/DLSFHAsHJvJwII3CXCToDhJtAsugyQ
m7T2fCAFjEgsAfdhaBR4DBdViptB2ti/YFNCr7RimMrGZCN9dGTMTvXtiiFNOwYh
Ev6mDSh1850KuLTjI/QGtKOWPX+GZIidXB3P5Q03ufumyKodVGC54W0tnZOrURFv
0In3JuQ4m2Rxeuzejeo/uEOEpC9Xfmmw1UijdayvxI5E/7cJsgklkwbF80fgdr9B
bd/86PCLru888LrOjsKHT+ak764j6xKjVs4qgy7jI3/5jP98xKXEE/PHtGueJf/w
1OItfTr/nCGwDd29+Q07ZwSE/+cDhHyep7Xz07PKB9XLtd3sw4GWQkCTKA7tOxlg
+n9TvSwIEbcJGBw5d3EnY1tIsqBDR4oQUXJEQ0iXFn/WViWAbUYdqI7ZN3W4zxM4
7XWOLxFNwSrF88UWswUJNho0BQ+Y3ohWJkRoRszljO9YQ3rTcWq/R7GjiRdwyTsy
/BSolpuV5v73qMRvL8WfI0dTpkhNOCJzV3yvkeYN9tG91Wq3lzlxINbktZSgK8wr
jaQd2UsAhQowsiiFXuUiKhOOx8q+1hBQdErlNSoXxtS/BruO03SNSNp9OQy5WqQN
F/vj8j9Cs6WQYXNIv1bxQ1IAPcWqh2TLmZE2S1p6chcK3ob3EHLU5UNkjDOoTvpT
35EHjGRY7W41j8wmSdqmzL+hRzw2t6P+rCql/NaOSnPAfC6w8zkZWrivGP4q0ydb
3QEQnbOH8h0Cu60DtRyLuX+sTw6/SniUk9DuU3vukl9b/WBRThvsvPNHLNGWRI7Y
pHE+hnt316lN1cIH27HJlD2528daMqMEEMYgyaeN0lZk8MDP6ME5E1I3KW4CDa8F
/T/IZm1aO+E5QCR54Q9w8NDSwBQ5M7gVzK9ijjkVMbU1uUyIdctoiXlK+DvwEASK
d65MPab5LWS+FY1dmLwbC9uEJTXXHgnGwErurmwBrQT3g78hO7hp8K7Vo4H/V1E1
z+8rEV2Ibf9XgC0lKFnT0nTp4o2N5Rr0ZuIo2f6cSsoZem999eq7fB+gii2purTx
24WLDbFdJgRBGc/jUKUUVGyi5V9svlHExk1nUXCnsiLla6CSfLhGwvyve35IL7XE
Ry8cbhwG/Yptvdqsn6YypyUqmr8JohL7lsxE3RqVOpeFPdu7UrGtCww0QYMbLQD9
yX4VCI5yfyKDfW4FsclOGPbiI1HFwh8IImboPqEQBvS2wwnTZDFw+STtZ7bthXO5
m5g8tCcaWIs3q+M0d7gVlV4L5/ORyEZs833yBnYizMv3PsszyhnCTwb/1JP36TkK
u8RQjql+33QD0eLA0qIeM8z/l3OObpqtDPs82J9zPJoUVDNNcU1nNjf7q6NR9OBY
dUCFHEH7cBZQt0cxRah51e65bXKKVLI0ISOjrOR+oE4KaQVl/9yHe0b2KUkNCUVQ
yOCuvkehWkIbavBwFdggLaqrzVzrMsDN+WszsPjY2ZQTywJ6bcAivzmsO7yuD3n1
HzK1w8/tPdJ+TQHtjgU+1ujVyd/Zz1O1Fu14R154BL0su8sDitaKzhwfvTSOtz/U
XB36GUhc63VXuBP80vA70XG+HIkwUBndJ5fqkYB+rEjq6pT8+114gDW7NVtEp0Dx
HDjp6N0jqXc2pjGnM017OsgWPMXIwEBBJ5COuu37d18Q7oGKMVJskR6AAGdeEt+W
+y+5IDDsrheG32afXT0IhWVVtIB25xzyRl6xRi071JbSdOcZbBTKMX64A+nyxhEW
Rbnqy6jNcvAo/UlceML8v168KAYwrNSJGvMhOVtlpPt//pb0juXtg/UXbQXhbpNz
UaUp+Zvh7FDd4uWLUg4vc2E24vu9uUwll1NKvmTcBmgsadaAQRN5aacUlAhgSN3X
erzFJj7VakjtFeWsNBqm0xyUF1LEMpNOe071mSY6j598rzf919aoInQ7xWkhJIgE
/Tu+UGpGj3vE0yHMk0gOOxBHGzGlHigO5EjhODzqvIOXEt8zfy4uA2/VsIUAG/fB
dyMB+UkU17r1I6PVSCjssKEgzEFj0uzuor2YSSi20FaFDF9lbq1A0pP8iiBkEAsJ
Ei6K+732XBDrB5VJ6mNQ7RI45lYQ9uBgqwDO+PpkKb+lklQ0mJAt1GAHDEf38FjG
jrANI3LulSrtgEWXaJOj81gW75oeq+7njRBbAXH66Nrz5iF5aBQFjui/9nX3eq/s
ggV3NQ53slpegZP8GPDEZZ6atGN88E51HjFFdd8P4HkO7IcbIyw0kPTVlzAr7L7/
Ljb32WCnpQ05EArP+vdqlgOaTHN2QEzoNxmRpEajig/4BraR7VIWG7CSpIi8ELLf
Efj8LPS0+vOentBjXBOL1tSbYHEoNS9I+UFd76KMmjBJ3FjMXR6TFq6Cfn+LCu0Z
Hhg2ioojKfu74CCjbVEOWeQlM/Xi/V0hH6x8Y02uUPRoikJ5+mKbv15gaftRG4fK
u9sgMj6z2Bs74uAzZxxLw/3dBUltrcgDWyEzzxlCwSDByQtjxwAlG2ZTDwLXxyRO
cj8cT7B1qwwd2PLhhWukb4g1AuJYfZaLVmyij3hVT1mj2+7guF0AMjgPjK9oBJyK
7yALq1EHKSpEMAClDzD+nfnxvt8fkuhQO/aMwu3+6eQaOBA5sBPsxBxjxXDjS9oZ
OniTJjLvt2mlmEO4DvKYERRYxmsH/BfcQJszqENvom8Bd5KfURrZX+mGJEZQ2pzw
z5PDWZhWAv1kKt6hY9X9Wc2mgOF24JvTXqCjx85Ej7sDa3Etrp1Uo30Pn6j8q9pV
t4QGAtsIfmQ1mwzgQOu9JheI8bMjYaWngDbU9K+RFjNoFT91Nj1KoAt7X346R5KS
9wDTteeZkk5mLUxti7b8Jp0uZIi1pLImFekpecblZppJhfMVniWMlNOdHhf6RTcw
HRas9xzYgAjrUHY8axTSCK9wPmDZmJRrDpILgJaYLTUOrqJXgAzL0thGvJYWrGm0
8T5JvxSU4d1w0phIYrrlFQ==
`protect END_PROTECTED
