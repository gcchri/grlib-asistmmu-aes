`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
512JbFvk342JCz9mFkxZ6L4UVIUBQzI1cWQ/IqQuxW13peLjPy/n8ewC5toaCU2s
VmfBRDcLINBchP3LRegKZFeCG+19YbtXFlXp1xaBEHq5/BJos6TDVv7I1W5dX1NP
EsCN+Idcbkt9YVkYyCc67kUIu01sx9Al84ZTZgLyFdbudu0+XdWdaEMoVaf1J050
K87F0IsV9XVfJRDI2Eyguvl2G5QB4DqfCpQYhpVVs/HJVcJjNkGKXrusHP4AmPbz
4Wcps5kTUVRP4JHxrJpqYKtuKbGGXim3FMvvjvHrK3/n07dSokvfgl1TnxREy2eY
AK3EQhUV0JEMWZe6aCFxj0oZDrXvwlb97k9cF2pY5xjh/v4lqtrxHcJnwZvmZYm2
sjxt2ENf1ughcymfeezEwySfhd6ZQKwnlsPFkjzBPATDVt2nq7uXKMiWCH6+H3Mw
ODJgouDW0uN4+8nUX+I/fUov2jAZh+6Uz/YWmJWazxqvyMdxHzsk+AKtuP0NxMgx
YiWlKAyISgu1daJ/sBRRa6P5QBL2XYRtLogXV57feWk7jSph5SwQAn+aS0sM5ebm
0pK9zvB3xxsr8qDgEVPhefJIx3oAPn6JPUTgZ1Qpzj38cFMk20hz3RViraVtBII3
yk3IBL0PnbKZo+k0FL+Rpp7ENckjJY7H3fpI0pTff60ouqzBvboE3h0YWCosm2a1
FuXWs20JqZsyQqvSm7Wxr9X2ai3GztJbEo6hVqXuosqB7fbULCFIUd0B9OVTx0Er
47OAY65l4NlGs587TVRgCjdSwCeHFoWeZR+6PQJCI2T/HFBJpop1DXaV4bhOdfvs
094LefufzzSdXVhCQKdUt5xYNamwlE4eiPefrXJipmCmfCGfqj1t5q14VwvSORBs
3+rGxMoL5G68Eq+8kp1l1IjNdWfvk5wb7SWCOOypvBJJ1nI3aTzEvWFLFRkIrUsv
4myhn267LAbEOXP2jcuTMdQH5ssziEAmUmnS0pLhxQ0XAOt0y5EEPdDG1pVX3TbS
dDfUe6FF4gHvvZLHfK883oH68Ps78ZqtmVrljQMdYceaB9YTH/6u82r1Gv+tjHgz
yINlK9tmybUsCXQIHBSoIFuGVXuvqcYhJFR2LqUTwFc/QoR2xquOXOkJUhnJIFwj
jGm7iANCrdNk/q5ig54YHZMAErXnrKlaMa5QHlS6KmMVzEAIIWd9QiRCqiS2VhNN
/TwI1Ni+OBnPc9PE+DqQU6f+2QnV6r/i3d6l1wcND8ERYgGs9rhJunoFu4TP7ZJo
fKDGVCmQ9GUiVOt1AhERdnPt8T+hG5WNWxJIXYS0X5fHQ4nM5c3L5g+ximq3IPre
OkF5tmVVsfGkz36UG/NQmrEVYGBXM/vZHpOdNn23m20WeXvaa9shqPOJ8MTUtVCm
l767mImBEEfs+5njnEZJmuwGowtA+p8kWsm68UibchaqGDTXmnz/Wv7EZou69TK3
Z0+6BMw6p0agfTKMpQwa/s3lFBj9nX5hbwF96nq9toQaBib8Vs37UsZ4mavY0Hg+
fTlBUE/KqWnspYiSJ6CrL8p3EUymgJvEXyVyPPo6fRkbsrkbjtx/kHhixf0bvHSY
WjuyyYsjJcF4Je+/U1k9JHBbqIhoB0viKp1+HAoiYWH5elPbNXojp0zpeJ1oa44I
HR8bf9LIOihhZod7osdLFwl2yc8GiP9djNm0baxUZkyjPK6Nxksw65fdqjWi78D8
uP+1LKW8T1960qQ5F5r+z2KG+E9Jm4bcIbnhSe3HScDHfWd5VOZ/M9/NK+2b/yZX
VUzT09bCVccYpf9kDqct3MDJnp+mReYqmB0VGQwb/qedJfT7UA49S2od2k+ADUqI
MtSrezv8IZwPursQInOg3kN7HUkESVDVWIyn+6mNnCA0jYU98/VLUIs0GE3oiilb
9i30B7LtEz6BavOzB9lN9NK2q0Nc/FHAWTfSqz+zKXbNFQ8QmDNAPmj0Mh9hJoEp
+ulf/SAANHHgn2hOjij6o7fV+w1dC8aA0/jDPrKJWTJenZWjnkBFoczAcRLV+i5z
lIpZtmn/tNNyEndVtvdfwNFOfbKtZa9EkVSrElczSkIiZ2XGc/FnSGmpoC8aQEqW
KanRMNHg4SZ2V2zbpvx8NY0ZtVjtz2sOaon84gQvLZMXkLqSdEY7F8USFMfGbvll
jJUfxHkcAfo6QxB/lmMiRw==
`protect END_PROTECTED
