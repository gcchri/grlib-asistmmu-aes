`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VhkodomT4Sd27TwKfZm8lXqHccqn7oAwKP7VGOQHvvrKYeQYDRhca5dVFcleJ1sU
yROB68FrpLDCc1mHIQOcYT7Qvm+KRQuXYnXGs2SPN4ggnwPPjhr2ps8jvptQ1ck6
NrM5TNq8wM+QqBsVnFcnRXxA9Cd1PXRFskEpd98Ag+IoOiGPYhIyRr7wVu+NiKPs
O7t3ZN827+ynPk+CnZM4J4AW8NKyOE6O1LcSFOdhaxN1wsYssW9CVdkUvNwtKC3c
kOSXEPnb2k41tHRkFaYVa/0iSBfX7P8xwxgTfrgppgvwEk13hHfPXNT0UqOtlXm6
eCmV8Km0pGfyD1v+U/VYar3dlziTHHVAqVJjpX1k+zhuiSLFDNoB3YkN3a/5syND
UwmR3njQZmb8Q+CSt1Sv9PRLUrYBZTAAXEUM6XfTYavGGRGLhCQg6WrdtLhE+ZgX
zm3vGAVLpaDM871CfsVgY9Z4nE0Em9dOS4+MqFxFgvYt2KoB6YaewT6pwC/0B18a
MCTP0h3pZPxGgtwscoGgHOwPkyH6EdXDvzuRlzeTVfVoI2fyyisU7kp0oiYDOu7I
r/8HVh9R67LNLdl6aFRe7DYsrVG552aS9osmetaV2gC0WFlHyiGc2Ys8tKhODMCm
/byF3Jw4lhqN2/j+/sHJi0DkYdogwnkB97uqsXKf/EUxmHq6OOGZ0JPlN4WczTbR
zxxuEuhqMHtzp37UgTDiSxzaCLAx5EcOvZ3CO6Wjbwwrnp+wZ2jmmvjwjfbtfB+c
1sgdBo9NWPBpA79fL6+sm87TNzRIo8a1dF/JjJhAVjZhvfO1iuUG+JEwb0IwafKv
M72awOQXEpLgvAl+w969KyOIBy0hNGcN0kazqlEWv4et1QOO5krinAwkwQJl7Qwz
9yRO8oKcedAyIaUHo/okNKlm30yTNt2HSxfYgtcnNPF1jI7PEXjZTw/T2sTKHO7q
Z7S9drWMEnCVNs0N/7Gfk2SkQIQEGJSn7V0hDfl/JSyWuFPTzd6Ou05cBK5J3E5W
/1iq9xLXT10J/lSa7AIdGGPvXwFMSQ5aEEfMqNgce6qe/Cm+Br15VRrdiWydYXUs
ytyAELAehesyD4zEpNaSbJwzwkvvvcvc2MHDllA6daxn4XfUWrSRRIw89/0FEqy3
JFGdJLTu9eMbuTigJUcVx/ZhDIJhcY2L2TIfutCgoC/+iiKzFS0TjyQ6lcF8bpoV
hJUeLIbChggmNHTE9JNj1JkJLyXMvAjEd71H0A3SmPxaf9FIecQe24mOjJfiTCM9
9JxLbIABWnl5nIfzsyKeeJCVXiSiJdIqBCn4VsmU11wcxU8k93Hk+8WS1lNiO1NY
0iJRYLMApe5hKUzTSIliM0LklFlbsE7Z4n1aBT+i/AL2p2dQ0Ln0w6P6V+c/gXNC
w3JymdnV394AFk5EtJXB76mK1Q7oR8SgdY+ucZow7Nqlmwpvufn8fbdL3yJdOhiZ
MWOBvl16DAL8+cB9rmal1r9ll8+ueC4muhQvF3Mk0S9Mr0YOQN6ZQEilhrq8GCq2
8pVCDLAceuXQ5zq4Y/ARtcYnNo8fXflglwGdmfq+ucym6IQOzOChOytcxD1q6H1G
wpmcP14qrM7OmnwYgmH8+jTi1wU+BJBdVrbvnlaHdtdOkh1ZNMUt/43k49eU5Vfn
XDT7YHHKeXUAwuSESInI3PiIWmo87XPeSXJ0cVNdWkDhkqilVXYFd7AMD1yQhea5
CnnBcll4edSibYwaeLtmbVBa8HKvab/RA2DH1pCnGDICmHgkd+py4d+5MoKCxBd1
eMAgnVyB//xqypOeiqHHPV+++ugE4uD39VonG1lzSchYfR6KuHs7yfZQ9RcUmw2U
cV82O6cVVxYm8jmn9ZNKDZUyov39hICSNAat6ySY1bMUspeqcpj1s5sWQROfntkP
/vbVTK9XvZG+XhTPxepqMhAEV+aQ7oW3T6R8nZcxv+JwhUctmUftCcJxwbDORHRU
Tj7MKS/2XgiRF2M1kjq6CSC4UcGlDqmY5d7r80io1ick6g4P9z4dfnCL5d2Uqwil
N89MV2DYaN/WXlKQ8mhsIH55JWE5Plg5NbuJfcFnlyoOLmMlLgJkuqDKPdG/sRjw
J4GzenUaiePaXgf9H//LOztU36SpL0zLNzhTQPD8O4lymDpPq8m9B53o1xDnNDB0
jUpjU/Zo+QzfHdce+Wq2S2IQRpZJ3NpE+dbQIcUIbOQOTRUl8Tf6wN2qHUbKN2QA
XGwZz8dDbEnNH4eknK26cqcp8PhWZY9xEZ/vpvUPFb8IH27Jd/I4iWuCnEHE6Qch
lXPK+LtX8Jks4GsXa8Th98FIOgXjVkbxi7c9lHEoZ4TvRk/cYn2OnkMXZOOEClVt
0yFMykTOJ5d+8GLtO8hF/AA6AUWFwbdXDOdvUPAo8NLdkD2+iy5EzKnOlSv+ZJjJ
/7MuL6kuy3m7WjJayMFIIn6knzuF0Rwwh4xSnw6Yzqb44d6OsQ0dlOuRUZokIud2
Yo8tcLI3ma31tCs2orR7ChxW04v8X2GbnN6UX6p7vHLwF3MUVysTbcF1hT7OLv1H
vmId6UzBFfcB8ykjNYQPNAB9UTeBlIGWsvvkJzDvWyyvNmaYEvW2vR3usdSeWGLQ
a29yGERnyfOOGSlyYVUT+xu9yItggvqwGDe/ezGNjipxLgOAACeXm03BS1UHwuFJ
sR1S+/T+8l41YSr7vw1GnFniRTMItQeS8cHi7zLj/6sh65wt3oCaf+vGro0tC+/9
pzV+Ek29qHnuvsoaLizu/Fdlw85jXy1BVuvy3Hp4itvr2pSluvqgAJ+Uea9ddWew
CAaCMTPWz/9j+q1xephPdQpQjg6wYvVGbYd0Ju5+qdoqDIjs6H0LgXIWW0z4z5zB
9DI/XtGk4waLNg4mjTv1RM3dDTPEwrNCzbJOjDAkl8U/EgU+bkxsJjU0wy2mHolq
mIH2BBC8fzV13YYyfAADzWJOax2JOihtIfCUWSKf1LL2G+wUKkTblq9atOXzuasy
rOq0EeqohCO54Fa1mDyUzjPrE8bGVZY8RryJ+nAdCe2qRIjuRtMdIgpLlnx93tm9
NwpCG78uuNwKcVJx0IHzDp6tGNq8zXz5a5np6ncboi8wYQcFVep2BjLx8Pyb6X26
VMWtgws4iONMjM5Um4Wf3gxUIO/i36rVwr8408f3KzGowJs+ec63hyC2xZ85uq/Q
MOdl8XLETNuT+lCEozQ/JDfmKglElVq2iksPJOXOEysdmxLemnuWfQuk5gKvFchG
2rJo9MUPsUBC6QEfVrZBtY9ACwYBBfn421nCmAtwK6Rt/mSbpND29rAgGIimLHNL
Vv7PGJxdFa/rZUf+UoVNCBm+b8m8jU4ZQ9s/+1vMP3urtS8g0goCc4CvHtmcpvnE
w6tb7lmBNOSXO2o+uCJe0Q5Wh45TObGlXCPrsFU7a4w1yL9v0UocImFD+q8W2If0
pqsRsC3eL+3j6ecs+EM4EwLZyJu+UwVRq+7hwNqHNa5dXTgVgmnSbfQJX//0I7Y0
4mE2zklIXTlSh5rf0Ykl1+LqD+gVdJ2FDCPHxTQQc2hf0BFwwLr9nsIaUUrhNqXt
aox+CgSwmpL7n7ejfAg40KjtaMrDpCmI/phRTI+vk3fe/yS/Vis/H2IfEB+Nf01F
nbGqJsk2Wgyc7oL+pJ5Y09MF5m4nIN6AE1RUj+RLMXNDr4L2L0UWgvfr2Ttuta6V
I2p7zylChExTSP/Prl5YedKjRhYQ9c2ofX+jBu01us4PkRyRjdK/UfaFDf83sC4P
c96DI4+YP/svVy0Z52hof3LYgILrNuBFAmjhhpmfe1vEaH5GcEv+eZxyb0KJpzwh
3nHpRuOR7dPWBf884J6HlCPa6gr56/XuiklFbLZJ0I9STR2S519N4XHdA0mG2EPQ
ZW9Dn+QQKNoBp22zHjwxECaktR+fnOIEIR4WCa9Bpk0/OIUItyp6xVSucYWj+YbP
9h9rvFnRHmJuWTZj7NPznhKZ91xtaLtl9fZAWYMHVpT5MpOgSr6to1JlOe/qbBiO
jB+kd8QT4oSYn1Pn9zaFCAaFYTu/V3TUtzHVkfDQLgIDG2mwIMljBvD7qKza78DL
8tqtLGyW+EfVcsriFhpvk9Jw6xgF7BEeP4bOSIb4ovfx9Jyflmn9g7Pffw98UQOn
oQGIEXHBgeMIcLebz3FIHbBc0/5OnnCnywR7L309fTIfLMSqcP+QTFaNpjsjbwfP
+9O8ffA//6a8a9c3ZxDvatyYZ6YtZFgg7UOpb9OjRuTQPbQBkRDMIPECqG9bAGwe
FDb9tSNTOYA3OJ/vXtIkL+owYGrtCN7DwRYSZ0Dkkpn8i3eiNX2vKdbtprCevSbb
vsf8yzLYQ3MVDyNszliniMQXLAntVXBsEUfTrnLUxB2EgmqQR1oOENX/kMN7Nz+/
hOqEGccItDoXOKCKG7dm/eq+iI2HQFJ4v+FH7RgJw/To9vBdvAN8oIsvr/xahf3C
p2px/0+pJmWZDyZal7cR8tkA3zwB4ANSatmSRDEkpLc0Yr9qAkKyBhQnkLE7vA4i
uZhpMYwMta9jLrVWzDxg3q0ZHgdobWV97FLx3zbO4GyKBRWN4uScUUMhKGcf/t1i
+8MoSHLzLO9hbvTW/uE/ndVAH8dG7OWvoJPPeN8AziIuYdw6PF/GP9yesW6GVOvL
1QHCwXbNI2gka9flubAINhoqhSO3+a2Gmv6JuZgttsZi1/EfHENUaKFQQOb+ho+7
tLkJBXfK66EwMnDB1vJiLavvbQ9q368tF8g7k5aSfD8YyZfZZH1zkvQ1ElqLhCt/
rrtBOYxKVBz0XHoNxSLWoX/t6pI7gT07RhmlOV8KMPc9a5DbwdeHyb/WqwJgRstB
usc3vt9ukrF5VBApmrGH2UnFdapekQb6hH0TKzc+HOof/8cHaWG9z7jeVM+A9tCs
UIywXxNvUSa77+Zq3VT+5nM9z7tf1bqnXZClRetJtMDXMj6ByjXn8x8G3y6TwpZI
8BrOBdup+ejkPTJZ0yltMzn2di8qxpjSLvSZ7qaa8r2sY36dP9xdVFgaIA0zdiM7
f3d92kuh6rh3P1GFLPb6ELtbTOxodI9ZCwF7GmiJfgpsDHfNgbUJwsFbWOfQz6jG
Awo93RggN+b6k2VXU5kkkKRs3TLpTRVfPBBvnod73LQLapIs9pMCbYfJA097s2eY
khN5AvlDR2VvAs98iBQJXjD2lW8HizT0NOd/wLsqWcUJntmQszy8rxX7b35dExDT
h+1+Vgiaa2jDUu1d25uijn3QsNpnK3DSg9qDJOyr/SR8DeZRryzxHmcYGpQw2Fgk
55q1pzFhs7RymsbvSq1sjNly8HcII9ObM/7jd75zRts+IpoC4akCIw8Ar+GGaHh4
ZbwtcMwyaf1Rpv3iOUfwnv4Up/v5HCFteLKrCShJWh6ojXnBamNzCLYBOTMyh1OU
P70erlLCN8cBm0kE0MmA2fPA2hfvkta7ms5fktJ/8b5kzUN2OAs2UJ6oZQEIxvP6
oAW3Ob5AewS3puzkFZaVpZ60e2fotwHaRilKC38k1xQIKceZ7SLnLeeKdlF0SByz
qVH6dqZj3L/yQhAhzcHY93Cq8Hw4LZSvhhJcJj4JCua64lbv+vSPkucRv8vJfbOa
fDbTE7Thhr+hNGABrNKBbPYetmic8+w/P65MhBnqhMaDeFAduxD9euBszQ2qWwr7
bFWau8UfY/GsOp2TiopuXQH3WdHDBChyeMYgacDqOowyVuPTjdJpEaa6ADteOpw1
0b4Jflqm6QToRdw3DPKhj1JMqa1pRS79nOraFWbTNoNVmTXOJYmcs1pI9Kdyql/Q
VQ4XSgwsMoDADYgen6b0AmW35WE3d+t1C8lVqHl1vDOQyIMszMNJmMdzRbLszh0o
3ttlj+UwJEkVCGizGyiGzTOHMfdc8rC1rERqq3+BBs+zqn1AVaryGNJ6JtEhSgsr
uYy+gtkHP9MwIZjQrsZB86aq9J5YPXzj7N09cLlc5iK+OwOeAIeAFs+45gotoof+
QR1YpHryM1IIE81XgMtSUF+FPG5Z27o1shAOUD0riSHuP25OQNLCrxaRwySSJIYQ
EhD6jXvY8vg16x78SdCCXTVcrNSRRjlv7YYrGFcN6tcPLFaZbpFRyDCxIXD0OuLK
K+z6p9z8g597GdWGh5u9jYKWi0qqByD3QDiouAO3RV9BGuPGmdi+cBIu9IM+FI5b
m2/Jf5cxxKxm8/RVn8TNtsz8JemndFbxuVb8E8cfMoT+PY0raiPCLmDgRGxShvqR
8bEr1rMH6LMHIGg7XMdv58di/LaNfmEvIe68hBlmJwQ8hxXPtryGjJpmW8UtjsL+
v5OjrenDPmi+ZYJsxJUld1qSrtmisYVAuGhmBpkSn0jW+M+mJ8sFCK7hv7sSahKX
mns7yK2KaQflPgbdAJconVtRaj+Hg8Vtfzt0SmP6MP0qzbB6UZocnsnY3bQJwkzC
hzUNCpGufpWrYVQNhNbpQo05eUqTGVPzUnUIqS4v/fTEyIQQDyXzZ00Li5Zyvkqg
H1T3ZBvuaCHusfJ4iL/zuJyy4Om7EbdRFcUNfZTT87gI3vFn/gih+kKVdUfdCOjZ
Ci3ISOkKH3IGqAPdEWmQKzfpYFmHwG+x73fVBb2mozHoqupgPWTyxuLTmu7HALqA
z3pj5LERzC92C6TZHeQq8ShHauHsbfntnPj+LT3whTg/Nft8x/o3OyLyRAna+p1k
RHqcsZuh9N86p69IYkZguzu51U55vl07Fs6Je0MeWZ1Q/9Je0sebx37gO3RtTRnS
aPHMaCbjNWCNmfTMW7X854WKzCi602QTTrKMxq0/xkbye7UUC+SrsRa/gz3Oz6gS
r4+HXuSCBzRMHqSHwYD7akMRX4guZ9AxXu1gLq8SsFC4tspPGJyAoOLUpdzJrCj+
yRaBzRmxPGjwoMmVV1FR2uwPsjNGenywkEzaiHverA47IQmTWloLBLyurr6YKFnI
IIu34VsiElLiseQjtlzJECwcG6BJ+ZKXcVUh81Jwnandw584kssv5rf4o4UymWld
H7wuaYTPGJWC16Ic1fZrIkGxGrDxfNSDEyXDSiBGzx+tbzyO3iKhWlgOcJY4K0Iw
B0SNzeoYKK5C/FFfeXY/UoZGt/N1JDqFIKsnNZ8LISVmsIkjvn6YtMy9M6tB5bbB
K/8mbO+oQKZ3XIzX/fxbfS+v1Bh/pdKO88y/8ksOdkfxDz67qh4V7qIxEQ5xsha9
TThhFbPWAGB5Z+iigIBmE9OaKrzRXXjQFtyeI20nmXWM8sR+65zzBaD9XT5Er55s
GXegrtHt8ZI2icx0h6E1YxI8PInSP2vcQ0a/MqTW9nbHwmt8UBUuaO+cnou1XqSV
IHmbpgIfWPVDH5tyLj/5EVXGD3IxlVMNdC6Q8Op2iabrht2mXOhHZglJ2lNX8nWd
3vCjgpfMBt0jErLdFHqELGIiGpFjyMYDZgkdvUKOYCLAnXNc6x8MFaAFngzTnYaY
+qKi6GXLH0B2ap/R4O2HDdmobSIVXSL7nxhNeBr/op8kbo9FErm05vy6vopZ4HlR
Mp5SlODJCAwrZWY8n4LNiCL+qx76BdWt3kJ2Kl75pe3+d/nqD1ZGKgLpa2irVg8S
j+mZX7zNMh8c3MrmbrZA/ClCrO+cZqZUOBETHgr9IUmwdvuexF1UfXu9g9axhuM+
fN84BzcSzfICtA8Tvuy8aS7dM2wR55hJaqtBIlJLHzsPXumv8zNROvTvNIpHJLqB
z9TzuHiZ89n0tkpHXmlLSsMX7quaiu0kU2DkUKEv4gEkjJAIai/49oE4EpuS42Yj
AYhHqtXZ81mBSs7esHcu0LhwS8zb3XOL5icCey5EY6fYpdYg5D6syS2YhgCQKD0k
CxhdgXnM2rvBbtY3G4U6ptExORR2LL6yq5RHmbbi2zWpWHyrywg/YiyMS8fxC12A
IabJMRmkfjdUuzvWY7M0aP1q8rPIdQqLTfbOANRdMd4d+KgPgne2Td3XkiYli6HJ
0dcRNk11esLnuIdSwJ3N8QDfncuvzKaF4xVLdhNkOQ/k4n914nN3JiJwhApQ6WyE
hLDwroV3ZhfGqYOvjtsTezkAmzwXdc2D/Wh5C2h6dsgnbXnqyPv2uQocHcuSq/A1
i0uKrYoCRxzSMNrM/Y6zK3lH/3nhAtBspux1uFOizz2Ivs7K5neIsBV0oVEEXQMd
WljI7kQai5JwuOBeO/pDPh55L91HI4j1ycxl+6vhuK80p4e1+YLZsubxYrf5vkOO
8EeaPq0GylSGEPA9KTt2Y4aKWRkMVw8bB/tk+XfWb5/ZllKakeiQA8ubYw6u1Gv8
AB6JHOcHKunDa4fLhrRWSViiy/gOQ9deyG7wGEuHFl9yWfOFo1j+NQKvrGMT+7Z6
Czc5WBgg8cFcSDOC2oVooeBPGUPSBrD+EXl2AzIRxPkGMjifWR7JPT8d/rh5A2aD
rB42m2CsjgKRJRYWZR0Ge918UBZvf4SqfP/IVTDvgxhSxeHVlL9myY2oeZZd614O
vCOP4e3LXuJhf3k+CfG6j7HzAQvgwb8goeArgQH5Vb20RLHKAWw0uW/SUDLDj6js
hOluopySud+e3IvjnyuQzjgoR0IqHMEv9hVDmvjM+XYLXtkGN6Awu0YaCLv9Z8Pp
FsRwTrNuHxdfckjmw/7/XobybVkd0iXmlL1cBAj1gY0NCNm5zWGLM0238h9k4h4X
xSaG6ubmKImGleS95bFfsHRE61q86X+RZZSYj1+qjEJDurEpJK2CVgAEhuk/d08R
iEMV2XPxDiLsz81G4KgsyQRCBE8t7P1pOleLwsKLs8u8rLQrqR6u6UyIySAFhsa+
DKAUCVkqmNwxKq7i6SJNiAi8ynztn2zGVtam7fKH1SLdxa451bGT1q2CjTDvUHlQ
DFQhbISb26EC/fF4Fegf49JTsPWedMoQLssDWdTAoopT2nY7igr6yvJkTDsnDbb1
LhCH0fiZCl4aH6gX0d94cgxjtoQNXhidn3TlV0DarpOk4QDEuZLkM6mcXGhtcr9w
Imm2qUyQJO3S5LNtrDjQM1xU92T1fkhPgpAIMh8FfdGMnV0CbKKzjpYZbHWedtHd
pHVr5oXqTspGDb/NwX9Y3Ux6VKHD3EpxJn4O/mJljshIPDuFRvHmGnEi7yjA+HqW
KaH+DAZnzRBDbzQsTS4gGKo+t6ouakP316+mplSjspvKIpDHVQ8Kw8wgtHpR+cI0
2Wbnkt5Vxps4OEMBE67ZeEEb29VGxm397TKkP66VvDDBKMDC6LCqZZ6YBCaU6RW9
9qNJOP1ifnBjIqm89UW2D+oTbUfuWH2HST3W39BaPjnJ2mExpeNZi1KhthiGd7u0
d21oZ09sUjuA57Jn3T+ZklDhFS2zU3jLdf3rUZNfOOSPnKWtBz23tJzc8jAxGtl5
FeRxYiEgID1XmatsJNqCTs+OODPHauaRmbOxIJKuxVi9JF5eY9JmC3Ggeh2VI3iZ
cHO3meEtWc9Q1jzL47o2+GV3sEEGaQ8ABryz5fTiGxLM2FEGc3fgo8vSSmc5EjQD
+ksgW4+xr92TeLNdf1pKH7PbfKJMHA3RZPko3bzuGeXpcNt33TXA+I7ttqhln9qM
jvCNKSLvST5Mkf4U8zS9aeIeZf/sYinTzROIez6QgvSn6scDUTLFn/e6sA2aQ3UM
P3lHyhWRE9r3HcvjpYjfXcbUCwfGspwCKfodVYQQOD8sfk7z93VYPZLyneJNZZpX
cn1QMuzAcbPPReYv+PG2nyLC8UZ47atOBzEaKcJ8v5aYxO108Xkp0awtVUIEb0Pf
QZ9Zs96ehBMU8xSv3sUOBRvuvpZPMnjkRDBPc5l6eUHaQMRIbL5aDn+KkqfemnsR
v2ng0ktl9/3Ptay++GsaVRfRT5/RweJEL47xo/rxpeaDyuyNUKFpH2q1wBbViW+l
eMbaz0Rp2i0+T+Tp7evRc698BlCOj+4Ri7jMH0/8eMaTck+UTo2Ybg7AmxkEK3k3
WVGecKpxZ4wIezU5Gf9iaCLQ4O4MWm1Rqb1kFKl+7h4JkcoWiCX4YURyfyIw+MLP
y1m9Bi7g4DCGsGdNoMfENxu/JHs4BAaJ6XBIUiQ25VQZezVY3KqKJO63LsuIdt1n
KqcEpF46rlmQYv8vIIFSeCfHikLbIeBUEREK7hOBC8jLuVyUdgxMeOXSw+pPDunO
YyQFXI7FFjHnZYBNOWzsYfo9S40Abz8UwPRv46IWkVQc0TPUx27Cm1YO4JOpAMVH
NgcdqSEvVrZIixzyhQy6y3K3Z7UFGuhgllWD1EcbzvUfqONlfNuFUGEmmose/ltk
7SNA2VrdixrOMmfV9wWf/iv9AYDS+RrzLFJFPL3piMVteEhJfH82+6HCdsdu1et/
LTNEAqAkPxKlTEfFrqMJfsaN0Xkz9TXMkp+JKtJbyPMz6Q4VLFMhXifljBgD6fM8
Rc11i8UI6Rf3Gsa5Qpx2mWZ6a74+YbH/Ez6LDGqXdoFuHkyuEJ44moKGlQFY/pfV
cyo/LpcIFSOCMW9Xxb+fDfpivGiLuISTTWEJY8L90DUptTk0fes+0YR2/vgEGyWc
+r+qRjhC+I/nly2eN4/G6QwJ8Kku3/eMBv4oC/58XC7Y4zBLPjEnEo/NaIsf93oi
RG2+Zt5IfsN7np5ToxscqAgfOFxv5Tg+Zq+CnJoTQ3/6oJUwtSjmTpPR4BfdAfzA
nanbrWjP1p774NN0cUTJoDN1GMf3zhxoPrUIHD4mvIxtN2980Mt9Rg+IN+GbtP+d
76QP1/jCOhJnttwDJ+XM9hcAMpucLo3A7C/4GbL3RKcanlGbsdTEz8RUqv8iUOZy
mc2YonjdsGaw+VxF1mv7+eVdXX0qn4wxvzEMvMrNLxBSxCW0bw6GbAQGa29ApkGk
FYg3Li3gZKDrTCU9Qq90O6DI+zzK/Pat+jhsrmolYYAMAa90sS4b1p+n3D1HCD/k
7J+TqGWFZnxmrSngdnCPMqZOKM+bT6HX9AMZbCRxF3CXM+9xSPWAT850HM8aDXcj
xLuggyBIBLjlN7SA+9rqwPOv7J9udXpYOxn7oxKnrzx9Awz6tz4lwh9yHRmVvWOA
pnTi8/ivX9WNnT98keBo1UBCmrUAzE5P0ZidURIfPwkQI0nw49lWcOcnhQaeZ5p0
JXzBJ8r+htt6e71VcCz+Fuyv+f9EVXYg/ue4S/D6i5f/vSpB1x/tOr2Dw3QHrJ0t
boa9UtiR2D9eRB0Zzg9bQwBKSTFBaJ/q7rMI596lfgTk5mcYSowNNrRgRWE7DhWd
vBKdIUDOrV2Up2WJ3yT+d3wSFuRe7Izdy10huluQkjcLHOmrlR7ddhuAsA3KZRbD
XD88nyoCQ0nRK8YSR7femyVdve82b4unyYcSQDEPytR36SO/zOjyFRvWYejoSJsK
f4Varq/fBQ09f9SpdZ8IEr6qEO6RhZLpwDETovsS4cQtxO7O4KCxjQXC24zrQgQ+
cqMVdcMlcQCm5ZDjeJ79dGW1KVT1ylrZpM4GjkMVeTMmvQqkY5IyVE3jykFQL2uy
AdznxVbDoRt146QbhsrVuEtHnGWVA7eI3iWkOdLe79qKqn21+b0yKTvd6QFvzOtV
yIOVHswBNc87eBZ678wWzW6d1ZSgBzj0ga07q+uAcOMAFQQFxghlNKMosp77tq+n
StOMuN9K4FgLT8RQE4Catco8z+7mnOml9+0DIcHbRxS0PDuyFPvVXeU2x+O92trc
0S2a6aKGpvsvFOH6VVAC0BScXKh/sydFnea8zcc75Wo6XEar7+FPQbgbvzI1b3Tk
Ftt4bY6ODiOGu6G7ouNGwDVXJ/yWkfbb3wsTEDrezzBOYewd7wlMM7tccRBK3m3p
ZiM+KyR/Y5ClkxicLpCFxVwfxl1TM2X/dT8Lwa4Se87W49eHs/9YDO91D27d0VAl
DtrBXaAwHSkZF/QVf1YYFMYAFTxKj/XkBXuDz2m/9glDnX4wjL4Ajm/ITjAlJOyM
y4tLfsNYKJRcMwGyoNYwAGpYRWilYcalQs9bn/S4gUkK+hp35WLkl27smG5cgBvc
WScjCcbtWFMQ7rVV0/8sr0CpJ+uwxuYEbIvrsV1ujL7b3Tj92Ux+b7XHrctWVvGj
I3dWsNOI7+HP8hLyT9OABQxop0aTJKtCocvC1d6eyPqm4XqS0Um0+F9OBM5XLnzB
RB/jVI5T7IvbnQwjBB9E6QGrcC1LM8YVblnOnIaAbAOlOIPyE/TKEKDm2J66LTem
Q0mHeHqdHxeXLj9Moq13HSe8wZefZcX8WGk8tQRUhns/N/Knxaxrft/V/Hi/qjgP
Gt7KTHfFCU20Ri6d2cuY71qJqG7xrkP2rxQcJ4BHsU53I8XFumWf3l8aaEYDNcU3
6FvuCNoCfav17+6DE7FKIR3PD+MxUCsQfoLf9nSFPlDXKXiedNrAicwVqN9qnznp
L2iGXmiV0Z6x6l5C7vlNa2H4iqVHcGz9YD1Rk+29FkodTmopDbXnfl97TeEDklVQ
jbub5FllRDm+Qmcq4J+nuI/Zn+p45LmrnZVO1nXUUhJEoEK/leH+9kebzrbkSLqM
u3/s7n1HdVvdtblGnE4ct2p9lkHRQsyNyVpC1mU4wG9m9uR4rVy11Cr88MN+C3A3
Jv35tgBvAONoN5z3zbiPfkFyM0CbeAsqrlAAHQ1VKxUBH1VKWSEG7/2hPVIXLJyS
cpOOCB5BIWYS4wggix5OU+UcRvzIrk9NNcf4P1yMdUE88htwnPasAOMnEWb5B9VJ
ouM3uqdu54bs8GlOs2llP3qKFIbmO9A1FBXN7F4DusvOHaWgd6xz+TvvIK3Sus0I
vVHBiQ2ciWLjj0AZT9PbDome7sAIgPx55je5uy+Yp2OjgTJc+P/mFUIwhTP23ABC
OMAuKSJBgZp165T1P8HBtPiUywmWKCNZYNJEVT9k2F5AIVH91NmXaGZPNubTM4Lk
dZJ2l/n9J3vGbSVd/Vct4tVKiIKtwMurSGrlmr6QtMJh/YT49Enqbqp8qCC8Y9Y/
abxxqkIX7bNZ4dRIkeNhi0q8OlVAQccZybN0G1uAkTRDw/6CKIAoLr0ZmhRmQ/+K
pbm2QaV/BDofsy53GI3QVzsw0VpB4UIEQiDGB4pYHjOjr1QQh7dRpZBkGGT/ismy
kPai1uM933xi7h2RENtTgGz0QiBrizMhJVGdMi0DVqDEVjEDqupVHeDrMtc+quSP
9DRXtQDwEKPXLVz/lxDvAIFqX8sow8VMEfTvKo0jDmmW2sMqeLhotuJhjLGxQFAg
YAJyf+27iB9Ikh8GyBAl9QsWOd8Xe6zCOOsqkzxvwxDje14sBUSIcVM9Zd5giMjY
+KY7bjsarBkyjK/rWjfWAaQ8NKVpvgsG0T009VK3trHF/Zk9fWdQNTAoLVKlOCnb
0smazXWteUK3Jr9xVxqSy4aXfyA9iXbPfaiW5OhierAw+CF9L6WWGSBOHgysLwi+
u47OIVGlbCA6HgUd0Jt9QipFd2fymTGnr5d9qxL2MT6kDrS/FgY7oNpPCrnAntuH
GVztSW1LAKewM4hgVppClaPRgqty53PVN31Zi+rcdtrn7K0L8D4VbIC979Vzr3Jx
AEVAb5odOgyGCuv6G1/BKfDHD4J7yR7tvuEaw9K/Qf8qo/5EyK3lLyCEQrY1k0xr
EzSZCb9WhXy/DTactcMfX1lwI24J3e343QQAj1DrUI/rvUmGcaAS2MeeLCdWl9Su
peiukjQX3XyF/LVuMHwW4lioDhwaMyGjOGseT7mnuv6YsNZUgOaEhc2RRxG0ndHT
Io8DSPHRWjVeWnhH8mFo3q25PXWfddOqRh19/wt8aF4f34q3HnGU/+DcfiwDpXl5
XIg8wZ836sIOB6qX30LOXu7XSs6xlpwUkN3msjxCdDhlvhbBRJb4y91ME3PnYd+2
2rcjSATpnvuPd7jtfgjw3sIVhF7/FuVIvYEqvH4Y+rVJeCrP5UfKkLwld8J2Digd
q0ACgmWS6eNUuXOmnBSr5i6a7oZHM40kSBpeQJajsp2Q/VVk5Y8nOGUHUhtkTzMn
JpDOAPvtF+E5kgqrHIeVddXMMiT4E95JOBHI9OcCRTgIeRDBQj304ZsvaJ8bQ8q0
3nrZsZsIZA1ZY3a7kohxv4ZF6jNR8+di08w7pyR2d9Tx9B63LR2vTsFw7ZgD/Me0
zffR6dM4Ie2krzj9htlfi/FCRGC7cP1XZ3qt1Nfzddy0/0jVuSKGI3AUPev3GR0+
yzovZA+PbFxZNKA11NCvMsk7K25Acal2juMDIyDfc8WiiHY5RFKUQRTRhFwi7QBL
gwm9KtyQWxTZsXq4xxOu87n0dfCTLdAD67iLjq2mJCkiBqBttYyX1/q+Fv7GK2cn
v4pvgiIF3HW/DtE+Abst7ms+QQr+EZCKkX0RxIHTd+rCuOqoL70Te1Igv0mSxjpW
EnojV5wGhMi3PbpMWY14WmlmlVVY7u9x/2QHrhcN6O/1N6PFVnEoGHW83NibwdzU
yFzYsfrisEihyML/JKNYkoTrm5JwemUT+wFOj/y2s1FsOlHKbSVQ6i51SOh9kZy+
eBnPXKZyGA215hL0PkwS9+Q3MsdQSlya2L28YdW/OdZdHbpJFcfdZ2D2ZO2Z6su8
HI/IMqoUCIV8EB2VBsI0+9XjYMc2Z8Tm/jUKBkRElsJOhG7swqrSH3nUuNn7rDFx
YLZdtZ3I5Ke/XV8yv5I6yJ1aFuMa1L+ZKD+09AcPG1DZF/52cO1/NwJXeKKdCCLC
NmwqDUGvZWJYIbONu8jY+Tqylc8R9dPdsPkx4347w4HIfGkxrq7mOJ5xzScoGhrk
9sRFS67SAOjWusgb2MqU8vZ5RnaDf1D+snCRyIoVkd3sGAtoY6HpPod2XRRgGtf7
8x+AIhgw67ydi2vMtyR6UBqu45Mq8EjwePrhpLbKvCkUhGBXGmhTmkTZoz6Bb86W
vpWkxab9nU32o+XI2nDO4MWtIPyio3A5Jh4U6IOrvORafWxy2GPwiDS0kfE6HcPQ
gCqTNpBhuYQ7tUaPD98sQLsWoMUZrynFeA8q3pD1ljIN7KUa5WddvlyVrhZMWLC1
06vONeSUpY4SPnwHr6+X3FkIsoHmBGp6S4p3eqyzh7lPflXgIAJUQQIBxv8VXUQz
ZUxOkqnLRAzyBl3DSbVzjgR4C/Twm1lPHnEZaT/mhYkJCH1eBkr4+xWfT5KMpgp5
R0WqIUJN3EdhN7eAwldiFsfc//aZ4TnvFOPmJdBcf2bZQJ6u8av8Oqohvk+MayAA
9ozUIFUzQS3eF1fyvUokVKf30JNXiZuABI4TCnpumlCWaWlqhWNhwy4G+qxZ3+5p
BiMwWL/iBEBg9nstJl+S5Fb6spQ+8ntS+3myX7Hkc/ymrisG/6guEKRHXHl/kmnb
hF2NasAUBvjNjY0zX7zaD3WvQ6Uhf7SoqV5a9XRwJ74c+xwZhFrpfzoJ9/42kk3g
Vf0F29Wo9rYcZU3amhs/syKpe/7ePu2qaLQqOuX3ncZg+zAOh9syA0DFwAHuyogp
+lnQ+BUylcW8/fg2QgLSi7v3DKnKpoAfeK4C9CG4iZJPbR71zaEBa7e6F4rS4utl
UcSbrPv89YL5EbKqX9zGGIlQ11bw1ofjVOIYXyQljvJX8/BuBJ+lQynqa1ktMZKd
102JwKAMFX7D/lOYzFNbMsf8vg7NJ9oBEJATJ2HIzW0/HcEv3Rp3I8+n15TRUWAA
SRwjTEAeRxTyJYvna0EaRmyGeVE7CLnXD4gbue0C6SRYRbpj+A5ICR38i7gPnIsg
MI44YElMyBsyF4Q0gwq+bOC9sWm74mE46XNmjJuz+HMQnEXnJyWAH/QTMWDr5tpN
4CVtVXZ8ro5M6xjn0FWU+2RGT8NRrN+BwaBy0ucmOcGl9VFjKkYMjBct57gMsYwk
PV5sOIoOPzBel7+QqVVa5NsSp7G8JJ9QfFqD7qWGkXpe33uoCIMgi9jPticJFsH5
kES2/v9wND573G8L8SuyHzrgKaTQnToQvEzsFtL0tA6XQxUz2kSdqkr1njzVHLrs
U+XiNTVVPJ3mY0DsRmkbLXH2BE0Kkti3mRN17vlyDYYUEDZrt6eUoT9N6HsUVlRv
j+1B9QHLAjbCsoyX91NzfdvwgSOmD82to3FnQmtxpPumxl+V7Agm6Kia+Rl+wmTP
zQHlljTspLqjWgvLCXjY0j3cMapPprq1zOybfNNywSvx8SwnwCeuyxo98EChGGYM
9w5NMbUCeycJzpKn120HXl4f1cnF8iph45wAsH13XDuDOtzhRmUg+e9LW1btJCWd
8jYUKSyie4o+mK5ca+fYkkBaLRwKCsHjraGMPUR7GK6NnFuhSK+UHdYpsW6tpHGR
IxRzAkXMvzyFkVNVV6Qbq9kl6GZrF6AQ9AL8G7QtUGamhq0v4Lf6MoSBbLuZJ/8I
8P5TPmPsD980XcBwPsOg8aYvhsNBi+au1nIIpfyyeIKRWKybYqhh+VZu92cY2pKz
dslUy2lkldKiH/7fUw2/juTKOzZdEx6J70BLRnEARMLLkGfrsBvkKyjuqa09BVxN
WY+E1lm6AHQg2CZ7MkhguVREzXpyA8Q9SGp8Twdm48FJroTI0D+oIusCYib2xQYJ
jw0ion5CvI1ECfsuJjBnOIEn3s+vumPv0y0/JXjavJHbLNizOe0F3CYNEVWzyk/Q
B42urL/LWfl9bYEnTDoavcU4gIzo6bTgdgclMzXuDZGBI08f2MyQ1L/zwYA1Rv/Q
6/DYZwmJtXWSI+/3aksdx2Ofmn+DoM82bhpMsPGK4HGZVKeiYIuaM2/tN8WROZnA
/6kog339z5BMEbehiItUHHqEgQH97iGe125L3vnp8K1YcsOIb51PZlbaVcMv+agN
urzz1dgp5l1RKD24MuC3T6+C+VpngKcTSk0tEec541AiYGdzeiYfMZ6QBodJA5dn
Cih5TShf9FOpEZgY17umi4q/fEQyPWwtG5+min57+QLRQfE/ksCIUSBOg4NiUixS
+VZ71Yd8PaL0GY67wqQuMVV9JS+oyWqDHeScy128MwcC97snXqEEdjWTQrNtvexA
dBkn5SDD5qiuRsh/qQk0fX5WIfLs/3u0KEMWn4LnNrhhesGnzmbcToA6MMsHODlg
2GgUOTtlHbQLQHWf0yIR9TCmfCMhRqMxbXAGACDh7S3PA6J8huGRVPQj+hLiZaUS
HA2nO1Eo+VJwDAJbCO3NWcUa6egYW+oJk/lZlzjWXMRitx0tqrjq3l6KQzalg2u8
KPjs+/8Yf660YUWR0hnloar4gOXk15hTFJ6BDLvbcObBoihIDypIu5wP7qKJRE11
maqNGPTe+dhJnrOaNCaEV/kQMbIU54/TszEo+ImBA44/TQlH53gklQGUwApTk98H
3GhhxTA1TTM62LV0Yl+Wg0XOlAK6Bvs1UW+rypF6IXDYvKrhQwpR/GyRG3DhyRGC
D2/pKfezPxjIpHqojdWvbj8BM7eFT+viFOSiGSLEvFYovHJqRyEk7tb8hNA8MyD/
MH75HpWYA7kv2Ta62tigwnDH74DGJscBwZrKt79am3nkc+vA6IlmnuozaFZUWvsC
nMuUXQwpcgbpwxPQWva4W4lNUUtdgjSA+Fuf4SxKMSmdcXbztnLebLyfwU8JMhmC
VrJsxgCs/Yoz4+MWj5z8FMX4GTZXbSqiF6P6MXMn8Po11FMfrJph9/v7vJ3rLqNE
CJP35CUVu0FQmVTHNyouwbCK2nfavou1OGY55pO/vGSwZu+BR6igqKwTieZzU5iL
XphUbR9+1QIVxezIezWrZa9T2L6IJMeKp58lsMfnPKfTB1QHEYwDv3wP8i/s9R+4
kNaSBEAHcJGLLIBV7iIrWcV+jEnaygPaPNHHqTrnDBieJZcaw0ZuR8bE65qF6M+q
u/LZ5utF8HgWkT6fT3jfPgM1dBHXrzLEqzWN7aMJltPwtbPa+YDxpLYnEI+GsKLU
NRs+C57dANvvYG9e6UCoW3jKXceAePv0+QIiKB+QjNzdL/KmD5xSLZnQMG4AybcK
zTbPGzOviwI2qmy5+dsVzdqJ1QnGqkITzRjHzxp8XRYAGgyfWDg376C+BbLXnKhS
yzGMYOiY1QPIxvinz3/PXe+ioB/Ghqx87Q3GWhAnMKDvcnx0fBVEsMwCd0DtJxhu
uU39zE4QOVViwq4LkK7rkPDUGGCjDW9mIDgpvdZXjsTFkSPJxdR9R804IKJtXBL8
M9onnZ2kA/By1OHXOQZklHCZ6mAgpgE36bB9OZw/8oTGqE4jV0heTLTHFlJ/KV4S
PclRnohWoAexekuGym7JhFMOL5Al3ENMdyJLM4naEJwl7YI+piix1vuv5g+WuZgg
1bMlspFWscT9nbiIOJIewjW7szLmhz8vQXqpuAztlx8BtHHZmFmzJv4ZPLI4TkId
Z+Ko0cm4Ntucylt3tIWG6qw/V9ieH0Vx2LgAeCV7mAwxsnlyZVB3b+Ucpm5VZWq2
rUI+HzdxGfgeNpPuHE+m9vgDUFFi2dNoFviUvjP2vXyLSgyzx0kwxw9w7dm0m6wB
nGLm0cfTjN0nDoMb8G9gJP9/QhM6U1Fh5sxs+iGMXoizcne5r5rQ8QptaEbXGyFG
Q5FBkhreegjgd+01JdbKbMRYgwomCyINrvzqOoyAQEduJkbqYH/HALSByo22TUL+
2Y+Lo7N9S9bfDtCYwJ+JcP0F+YpxYHfJwXak3M+u7bD/MgSeAzNTMygQGiNBZf5n
a3jlpnLNsBztJoridc+b/i5ME/vDTsU90zjFzAw/TojSzowa9SDPDy5/uA1QUc6D
C+8X35Q/QX/jE7Jbprle1BdQXnjq1ce2gEd3T0NoUgjfEGZhHf6SmqjxTGVivKF0
jIndfeGoXcft64ziPX7zM283BE3RaHZb1h/FEayiBvF69gI1rt+uASE8sJ84XUQ7
fVD6Gzwr/k6Lm5JzYZ4uReLHotvMlE7F2qYi35gAtg6YWsurlPNYb22Q3yexW7NT
ZZfwCadLtYmIxsjBZO6AGb1AiASZiZzVQfzA8ISlDspctpcdov4HLj2OYoDlZFeg
uXKQ1hJqmYc1GvXCBIPAoQWv/nzs9VKGVDYuShf/+6t3rjmKso89UDvqBS4FbOLe
rhRo4gpiOcTD5XTVTX+NJA4jnngQiVT1TJSj4je18+3rS1IXCbyXnqIYn3fEqEu3
kKZtchFsWXrut5AVr/4OBWqyi2rElPzps/48WQSrVz55HQ+vrE+sWxwCmccZHB5h
TU9TqFA9nrpXH41+Kx4MpPUJYXNtajqwsGal9x1L5Iaz5qprXsXP79rYftUktafi
jLxk3di1gSj7disV6N5APxZkJ8RZ7sTqOcWprQCz3HHw++FbULzC0rcH/Q2Q3oaS
H3zNHB8Xx9uA1hdnnWNE7FxYS2nHUZjRYy0Rpqt33w1H1LdyyytOK+yNOUkqQCwE
gVheJfm2itPyRZSmSasq9VwVVewU/8imyBSnI07AGEUuOcMtweZMQkdYPhroXoaN
PYrtqQqhOYmk6hAbkdN50WivoGvfGtecYmcOWe0LTyYYVd42qVmPa79kD4a9Fxa4
gJvq+M2FdqRxb609F80P8C6d5MSc6ur4X8xGkXyKbOCs2DiUby30WzEhfSbasaVt
LJgOZqYaFQqMJOebDsF6CJ0BQI73/kZqj9rB83z/wjO+ixHltT/9jhlHuBp/WSCP
GLBfzEyqpdIOXGb4jWvgfzRRmK9FKONJ+v2CF+8hkBHpS099hPE5TAtGSzt8EmeV
HhSK503uRYb9ziWfXoQA4SI3g9Ny8A/gZdUWuwIyCQJMtqru73B14KGeCfoO+6s4
pi1SK4+FY0sz1Lak5MC+DJ3cvooipASC1h1VKgkx9KH+u8O/Rn4fbILd83dwUQRG
n70vKIMlJ06vlcJVaDezFFS7uZ3Y/ezi2ErjsPlTqJgiNLAzrMwbb65tCoqapPKC
oR5K0+Pe5/pQV5DUlXzgTrS4w7d769EkR4lP4ShGlJvFUxomWoDjtVRrHZoK5MTI
SXkyNxN/QrPIz2LKOcVrse/p0oVXvlipOX4kfxP46jTg4B2XZPYWoZ1ZaMojTDTc
vzs6au8F5T2DZKbCH1TpSWDhaAqwg/RirL3wdEBHlCH45xhr7IUjHTDfLIFloOyP
fQeEPW+3qpuUzkcixLobg7LNcoTrWzUPUEaCgWv0wffnvbuDTzV66T8QWnHUP98/
o1NnMYKYpt+ttm6Ht9V6JYIddybFpKmFB2IdRsj5l3vDK5UfmDY0UcK8WMwa4vrl
83CAbjFfXpnkGVV1Gew428uP+bY9lFdQPnkF8erZo7y2he2cjDbCITtvEAb4t5gh
BlhGOlJEiWdz5W5MVOndcU/REK5cVCrT+Kurd1ngXrbS5clJk2k4PVo272cnkS7K
nfnYql+9Rfy7RoNLYg/8QTcV9tkMWmVRxu7ztCpXwUTru5LC4g3hr35676zbSKN/
1CgnTOxvPl3twzYT4sXEW6Ski69TsMSgLiPrWJMWDsqn5AdjwV4UYsk0SZIlXUod
ZQrv6Xv5Mf8tDbALLmL9GEt9y/PlzLqro4YA93d6xSeu69PYkxJIc81AWdFDTIQs
wnw53axPZuZ7RfYkUbbMuWbrH3ARo2Y/GpqMGnbd4d2y2v/+nqDuXyUNInbrKj4B
35gaGPMpFng36vX3rxwImE2D9PoMRjLFPIYbCwDCB1Xk/m6oQBsomDi3LU9frZCp
coiW5fQGw7Y8vdkPiYYEP1rXDEpcrDMen/lPrJP+hG2F/XRMzNeJySrpHnMZjtQr
fZfG8QMyyJ774HjEqnbPbDN4JCmjYv8bDUzor4FJLwWjR5Z/W4OY0KiIczQBkTy5
V5wDrVLiQabordtmuDSFvgJmN/KV7e3NfOR1i/tMyeLv+dEkPZ0qkoi2bld1Kb5a
UIgf+1L07vco+aNmR/YEIEtVqypVXDXPMMLLt3bA8WPlnt9sHVwndoGui4u+fXEs
1IUU7jB/Q7nYBEA3ulj/twCfYkLJ4q4i91/yU8l68rlHNPfwqF7wgpKh+h9ANWBV
+aQAdua6tpuLfrnVV/iiFhzqgtIuaupRceNGosheqXObg2JKEdl3imqKh5jsbK4N
JtonVFQP0Z1UZETuz5pMrQK8T0clQm4Ztu4lXjIE7POEj1rhorq1q30SSZLddq3T
0eJ3ekUeY48+j6tUBtuGw6/K3mzH9MLyV/tbqqOAoBQLYwANdr9lVbQdllT5uvup
caVBdMQl9X++auMcgxGqFrTtwhscNO0DX1cDa6A3mzUMPGBsmTQ9CvR4pxNZSjTJ
+fnJJU+3n6Ggg3fVjf8xbhUnoSO2RAS33caePTf3hc+lR/EJTXF5a7QoqNFKT8sz
AXO7Sby+2TmdnykwceFcJ16fAw5flUCEOQ9/iIMxX6nBEqxA+fl9M+wfebCAEtkF
ELRDw38qGjToz+HBadoP1tYRTtlDCft8JRiooJqkYSTPd9vQ06oWBoE5icgrkTf0
5xcmuALPuXmmh+/lnE0ILahVSohSDsjw7zZxxK/p4tIrBAT0esD/jZvrStPLl4WU
I18RrsiGbK4lISQacJTBQlZUDqn3ijeu4KUM9DfbgvZTZAGH6q6kcVseIXixweNv
3PLEa/iU69/7Bd1Ex28H12OxQ1ci69aZ7V9PUsgMJpDCMeJ8XKgvcC6l0g4BwVIt
a1pmEaPIMdOTLpdbybUw6VR0KlKZLV3fEc79I7dzYIceoMMsGbEpiHA8/xYbUs4/
tZk10XJf7UpTLhf5uxzfr3Tez/pmCsQjs22p3il4nzjFWeAXjOxpVjqbsyouWipa
UYOttpuBWHek2YOtdURMhM5JQjr9goMM4DH0aRgWDbesMjYtDUy4UsW55/EJ5Zln
HPcrHkmu4Ib6VlFT5twfkCz+dW6ha/bqtztMjuyxJ+yvAnzpHaxJ82ppk5khpGze
S+y4nZHm1w1uea4V/98DGPwVdDwYGOvW8uGhbho+BvuJONcZ971iZwegE/hAn8nr
ftU0zfmtcxF1DpOUZPFTDPgZmIcs+6exY5hs4El6AHBhwP9BrjaO/1M4/3xVurv5
UWODhf1aT9P9S4Gkh6RKQCESvKkYLf64I7jdgfxt6Eg9ILUPRCC5mPSzNu89oSuJ
GPf0rz1UmQyBTEIe88+J5NIklsL7TNlsAJLx9816847CASOznXLsmSShB+E9jusE
x3FJQCE7nN9XOtknbj9kF9M/QJpHfcBN9bmpOzCRAZCkepWaoybQJxnSHvTFPnkR
mTkzLFBNKFkPcV9gf/8NdxtuMdmJKOyTfq7ssedwsMpx18zsaJ3jnhZYie0yQ/m9
1AwRSah9vC5Oh+AZ+w4fcBm6BnaIfdmMkVCVLBsw2IRDTUNJ9Ll7eDWMe73p3iQj
oWkDwBH6zTVVdY+vlv31zT2XV+f/dMBKIG7KHEb13pes7oinK/RuvV4QOU/uhgaL
i0J19OHYCaKW4+e+LZkwhE0+hNH0JD1Xvv+oHeDeyTGZGYE2OmGhFtcCG2TqABqb
O8WdLTf8IOoIG3wU2wI7lLpq4aDLswXoRCbfXXruzf7f5Gy6BecMvxXwcGKHbZL0
+0d2hy1NDLzxIRz81oT5JCizrl4W5WYss/GPrf4dGEEWm4ONUnDwCezX91Ll995c
eUIWS5+Kd1XpyqSouuGK9E6MnTvaQDNbow45mfNKIGgykK9XPA9xsTxg0IIbDsXE
7g4fXGT/rfzq++i4cnpvoSdl6DBH6mK9dkvSNPF4GHmZa+ySzWLxBm9TVv4sagEt
FYlP6B4wCjjFeVljecmdQ8xDXef8mRwYr1jIt/G/1URqxiRbKK9K2SwMO6H382uh
vkSEmbDpryDcEngettav+bNtwfmWNN+qsTgNcm457WSjvrI9cBHx+40uLjrLA0o5
proYx1ZAftj1QNRAqdwkFdjZo2uG77eieieICBK4idSBvNYP7YYqsQOTAa+h312D
3xu0TLmcngZX8nS9sAe/i5qT66BgFoW+WjPtQYQ8Y5qBkFeVG3GdBXUyalHutTyh
NgnvxTZqvub8jXhZvUheNvOBZKlWlFI7pfRpVTNEUIrTk4WN+DStVCzw4ovfz3W1
c6ZEFeEfj/JJ+HXJjiPFicZ70zzGJwtJFZXD2cuuupJh/MqprPMfwx0+NL0qUa/x
ftnPPoLdyglvES5NVBeJsTrbhzFEpXuZCYk37rh/oF4VQnn8TFnnAzrAbqut15jf
dKxOiP0uxNynORKcpifNSjuwx5yDIUlHE1syedGv6r66TRjj/ZHthUoTdGzs77jw
L1GvH3OoJ2xi/IuyQYdBh6y6jZQg6MWN6uph1HGtHmCJb/OE8v/oUxJzb2pvoYjR
b6aC9AsQCAbm2OdaYxVnO8eGLXrz7lpjPWIxCqZH9QnmT2KZWNG5wUPL7jn8BVYk
dG74k/HthvVKwJ7xe/NBQI4Y01jmHRoaT9A9TyOtdHKRBl0hX8OLoadnIuIO2DRf
VTh7SA/jVXs3GdE8xRymyKQ1xvb0G9sYgA315OMAUyedDysXLJ3qqbM60/qDsQwx
p11O1Yq3Gfhsh/4yHMU3LoVHyGIxt3IVAdMIvtTjN5Vc3ccS8Q/TUta55qkoX93L
fhcTo/nuKm5KApTA9YPFlhLuieYlf+0tbetT3P5eqhvpBgNQEV9jlgvODZoC7wup
sxqlaUdNeGFV6jfqNlkpzpMPYH5g5smRYRTKrWfr7iZchicATI0C8FD4DC3lz/Iz
65c6cbIPb9uECsRGKEBz+ijAMCY/OnqCxneAQJbEq/2qk0uUjzIo1M30U17rheW2
dRkR8mrGcbREZIkSeYO94KYd1awVZxzLumzbVyBI0bL/VH05vdA0iHhHbV6qy696
IUInWN870JpZ7gdd/6plwzYs5nIcmEZaeaSx/V4zeRDkBaNG5FUFN2XLXRNHhwok
X1ox8+JeNy2GO+aG5hXjkv1SJEgPz3i1GovsevdFRrPJQlw33kH40H+Xhdk6M3Gn
SjuJC5rsegEI9N46uZ6L4RDv5FU19zPV6zXzgmamUkUCAkm8FobTOJWx4ws4Jyp9
QqIT8kAkeq2nZmlJnjBxRZhnAlTx/ohRYtunGupSj/5VDoylGcO8ng1S95vHkoj+
Z+KzVWPSl3b9eZ5urkUKM/xVVHwZaSyaJLIyZaW/TxZ57M6KT4jN1+s/a7B9nlfJ
QaUe1Kgd08RBZmvN4WJxgT5qGfIrYop9HTW34mZK7JVYuSw55XYYHacDy1yI73xF
vNp8rrJmUCrJv/31vmGO7Zc1fyPos3gZFASLxnVIO1H4CmvHOdVHqyWdRAKtZhWo
rwWXDFo9YTiMV7qg0l5+exVVoxcQicilEY0RjVzmZEWU/3qU63WdkAuYnWFhOTG1
PvmtB1umZdoAhJlXRdavMt4G8IFNtcij/ky53FXIsKy9sl2gVCPmbaUqFcjqRRtU
rjgv2KhvY1cfzOLW2ys5smOE73PdwXbsuwRnzhIiUlOpDSCcMuAtOS8duiR/+qEH
71cu0vW4hcA8wT786WSBBIMjpwU3Fu8fTYheulhXAPJo6c4psr+ABI8rDCeUzwCe
e4UPcTa06X4+EXz/KgyJJsHyaqpJkaIgzgoU05gwuKBnxwKkEDuO/LviheRTkznI
d2ulrH8RrXbqEr6H339yr64J7VMrqJJhjSwLUX44oD6aoOob33HT/woL6jiNL8Fv
4SPsoTtxMUFT7Jgm0HjYi30papeRfgb8DsGT/BjsaCJhN3XfYcUpz3cFx7O+fWcL
Pw74OFEadDBtdK5ILhV50tfh3Ewlt17juOFZBwItXOAeOA4c1jwQTOyupZAlxrF4
TW+4rMbDOjP5P7dZoOSLt3P8240xaJGMb7HSBHPo3MeoDlEI2Mt2u7xYuqsqskRZ
gNstqzGoVdoDaIXjGZ6UAMzZL2ISgYW/n75H0HB3fa1wBgaPjPOlifpbNgOaudNL
2SLYY/YXi0LRz0gEseXJ6xoWZpl1iVk8zBAG6dBEnGfDTsf1XlVrBjcPLTGJGlqN
W8UikpxLtv1qmXjUifOhVNZy9ul3V9G7wC1RV5U9YnrfCxcUl8DBEnXmcnWHzDAY
LM4Pm0d+C8t9yVFh/Xzo8Tcm+GSOO9fwZRBoRel/Tw+OAgvzD9zEAV+udt6ZlGsN
viXkgjEyTRCDvw5GrQvMIJTVVQWvwBcI/D0XXycYhH0R6ZPDdJcVdRjR47+ZJYnZ
FTgqsSABHcFPVzfFqA4aYzp7P4eHJGGi6Fvp+RCTzwOxitVeMlvxFBpeJLccZW9A
pd55JLPJz1nD3dDOm1pFURa5/HTzvAtqER3sya055lhZHiE3xIZFgyHAyBT5S+rl
ze8JGyQ1MuFFIFamXSHE3esz7Ho5Y4yNWvcGxQUEoT11viCKndR8qf2sFJaLBfZB
uaDA2T47/bShP5ds2l+xisBYrt2vlizyVmTGUuhuNqMnZdOjCwWG8WgjVk2jn5mw
pZpnMzcT+CGESTgLPIpb+ehhLx3LgT+dt8TwEEs8lWInBu+PZxU/oQPXinZRva5l
SclvucNlxhk5t1EOXjd2LBhclfR1OLMwMt9fxsAVMK40ETk0MrA7ia557b+0qINP
MY8dKEq92fTXN24g1yP8zEJqiol3jYHPQo50mV70Ns6duF5VhYTj2tylMu+mYGwO
e5FNO2GtZTHdqK04R1FlIslE/a4jOxs41PrO3ZDgf0wv2X2oPGU4nelw5DbbUdfQ
VClA15zuPty2Y/HDdZNOBdbFtCnI4sAFEB4pEkuhg9OCUKpwG5/aWYcKLBCNHZ9d
HSwDkE/oO69KTQhLyFlGCvq5rtfGktRVMzhYtjJPHr59bmPIWN9A1r448eB0rRmK
1VdzrwWDby+mxoLh3njX0cKelAfIhKCxZA0cnj80X4pksIxna3hLS4DqzzfSFIZ4
b04JbKrSlqjqVx+mXOROFcyadbQIYARN71qYw9dxwK/3f4HzqqLNQFBioheM6u0P
fjFP0Wrg/o65s8VVASFh/ihqjOxGY4mTBUEdDlxaYnYByEppil/4nqVpZRW2TWYo
Kfurzbp/NShQr2Tp0MyNDIlPhqqDJQVGaktqHTBqUgXdHj29RXUsRpE7UVCCIC2f
7+a7ZN+VdEPITygaYOXDt7Lj/p6PezRk8zXga5jmOyo8Q87EpvYKC8k0h46TD011
IYZ9eFsitr+PD7WnQ07qFfJxi7I9L6uXvTAyVxHhG+7wEL5QtF1sV59wJOHnSwjs
lJPRUA2uONnaOEPXTdg7gttilGfQzZRaMkYSO78w3WRgb2SFhtOiDgmIymsHqVHT
1xiY8gee9zKjD5kEP7r0CO0UQxHdse3R4X1JQsh1SpNIEgrseETfLihKrr6osRYj
J+iSL2kvASik+LEBi2x9+AHIlNuSlDMo15CF58zRWNP78WeUX+hP2eMj0TVH1UWO
dKYhx5jpH4SYe3TFhP1jP5FbzIokB4isDqsoyDFsJBwHHvYZrCrEg6ybRpo7mdRM
Wc6syVyekGX9sxW46GvE48vlNWIHcnAgGvbPAAX7oyxbbCfIBghLS1m5qAv6IrRZ
5EsBK+DZyh97+bULrrNhO4PL8nJ5ePiNPYtmUWx7GGeZoM1tVkVdWO4S0LY+6EPi
Y6iahaOojsdoVV5emZ0cCjJKiiNIDa1VRG/vhrz8fwTl4aQQtIBw+/cDjX50hAOQ
zyvFUHHG0PLqvrYBdsnGOX98ZxsA5TVHAOmbSeZIuz0z5uAGeNtTTpCgigUQdp4O
cMZzquEpg8WYMiOqrG3OOj7qfkUy+dDDaX2cuDqkrpUrO9UCH1TXAY8xqkyr7Smc
pNjdKjC473yC9wYzpOuW9Du3R27Ah8jiy2Yt+C22NNNPFC3gXBBZQDl8c65ZMdge
68w8Lhe977lrREexQ4TPpqJESGqdUcbW9vXfSEwXABr62Te9wOcDvq3tN9MPCuKL
82onVkYPXU65BrEr2DjUnNnbCjWYbcPRK4wqQYFkf+N9Q2Qkid9UeKMAt5REBThH
GTu2bPnU1iKYzZnuPy1NrEyikQczzqvxvha5VULUoz9B2gckoVQ4vG7UGzyZOavE
i/O+qcpqjqLqp2IxXggC/YKTyJiG2ZjwlWTHRoPz+gFKBQQdTgn9YP50FUwKAqRz
RWStJPq+26ddtJ/ZyjipqXQ3TeXdM9vApTOaK7ne1Uq+h/2hWxROGRXEobSY1l2x
gBuLfMmgwZfM1m0Ikn6LTuWAtoTK14iCNrRaRvYUlrasxUXRo0DLsDSKTczR43st
Hj7WSEo0GQQ1mrLlmRooULIbMHN7PAG2TKw1runpSbuFNRk3/vKw2tVEMzL0rrvY
9wO6zMH8Y3xjlYE0QUW5jzpnBGFI//IGQu5ILBR7dvQqf8R/Sy581F4M0Bx3KPI3
DgwoCkF4llwPJGNlqMoTB2bK0UCZOZW1MM700dSH65KabIgqA1cD1Fe3Dc9NrGZY
NzybDfXSkbrHZ6w2NA8ifS1Krm88fkbSPdqfdcHcRHO90Npi7ZbtbtMW602eIoi3
FCKVJdq/XMchZyhZbjQAHg0ssv4k6L0AJUxqzGZECWGGoM+gkj8aipsxCxd6j2As
d2tZq7x4pk3ZSMFTyPFASL5BORGFMkgH9QTv+17yqQJCLIMqvWffZJB9TbB4R2IK
REpiqjif1Po48h1sbrHqBq6yks6T8gW9dcdONAgFLPg77wokwEnrK1AgoUf1OZBa
EEoQoT/IzlAQV+RI5zoFJSO+D6TExFqn4LdDDFiQlV8b+wiWDNyoWnhipQ2pcd0A
eYLTTTjNrLZ0gkECX9ugH+NKFHuUaPz/XT6JPcyvZXmJVjz+mv/slLgrFD2+AN/4
l+mQwq+7VAWBuW+0xjxWfHwa0STwbx356Bl6VAt8Z5ZH95Y+Gi90lsicGR55zo/7
S178/xqLprVY/BUWMJ+z//o/+7BMOVrwFw6HCD3Q5Zm1MOuaxLNVnQ9SEAKB/ApZ
0JRpAOv833cbU1HvtcegBZuNNqHvxaZ4XJFpzjhnfMlZBfQwO7ehWKziKrUrLYX4
hki0ojDA6cHOi3nNrFuDqaUOpel005FZgiI5TGw3fb7u8fyxy7D2Hsff9LSVgvgt
0xnvnErsyQSyKCda6Xzu8ZiWkgMMjbP5rkx46aTkp7hJj1Uou410uJDbxmj1pE4Y
V5CbvNrmcRcaBVdlj8b6zmRhlcMUypZaa/h8XSAo8utnSsYU+TH2cKUqeIbDu05f
0PDv8z+5tqkjipvCRQKqRpZ0N5H0b40bKg/hdkUGsuI57v9H9/pYt5Yq9o9fxTvo
+5gLyso7LhMG4nYWYseeMhi/6T9y30bxG7GGgvIkA1WlFQBxQgRVLxse9eelbD1j
zZnkc+ED5oeXX7LEzN4jOj/OpUKcnxKZTusQIooQ4NDUMwjtR5xUCKWwYkgnfgy/
ZGDK9hO+8Q4Oep/tPMl2ZBTF63pkQoDZAesTRNoqA+RCgt1QnIF6gPGC8jJuKh7p
v860b4RP390MFeeqs2XESA45p/lFlbvJFnbeUmPax8n/j75FD5e94NZ8B/JN4FM/
FullLK1SZRCORzp4Lp+u2vgrBJtZgXZrfl7hrtoCe7/1Oo3TE89KA3GGfeAvS8ev
+Agw5Ce4bOf8zkPOQBA1oJDH2hLahJfpXVHI7vlJekRjh9Bj/o6Vdl8hPAr2tazM
ngUBSxIb2ZbyVYIUfnNJROgzDLaOEVGqlRjZWv8FLb/kqesQip5OxscoNWiP2iAk
1/DrwB51o4/4XkLjfU8hvWXzXm3Iqi1y91bvlnn+crn6x0D81qwWRvYhiTvi6Ack
sTzKcatpuY286E1FoidI++zjy/o7azeTf8Ab08pLYd41/rw2pe2jEeNx0bEt5yNQ
FCqrVkIONtYw67MtXemHx23A/eWfPLQ9vfjqZegr8w5L0LCea2YHC5Qz+P7Jllb2
K2xSu7Qvy0e94mSml7JlJI/eBVxg2YvAgr9SFCDqppxwKgZ75/zb803SThPgxi5w
Hn0ve5r2FxlrusZEycMZvNKtiIuA29SXsRlXAe9rMWWTxcWdEdTvZQ4wx4LhpeGf
Z7K+z3Mkf0ZD7a8gU7VFENxXw/d0QUKxeew73g9pFLLAyhvIoW5YMBqQCQu69d/l
vTQdjbRush3woWR61UC51olEaN0xeOJPpvzIaaz97HLiim1HW9guWT/TUX0OB7IY
mlZbFr9lawgbMZ8F2L2u95kML2q2iF3DChsrcl5e36l24C22qojU741MH3D0Qd8g
Qf0fS+JVeQJmVAOyZ42kzeE7xkam0b7jk1XQoKVi/IB35KG+j9CJWMoPs+R7z+NZ
bWvMt4OJc0A07E/TLsKq72VjugUxUjHk/qN3VBuZyRGzhBAwEuHQsgn0QQAcnyWV
YwsgkkjlOeckzLcf+b3+ZU1XYz4iFd2KPnYsHtG5PNPMHKkThZh7TmlBP6QOyqNS
v17ooFYeLfJMD9ywPHXCJxQXWoZrd5aVa3LIdyqRCG6YElRPxhtNOQHC9weiG6Gn
39gw6YueMT6T9+TZNJ3x8DSQglVTtMJCUOaM9vc3ejpyJAM55GlDAy6oet78hRVd
S+Zn6ztonck3uQ83W3bJz8b5qHHf7bI82AYLNof8PkYvrH7lLcgEYNGRECmvgmH3
8RRO/GG5+iJia7NttPORp9nPtUjhZ1q18UljMsAcSyX7Dm0TRrddOfpMIZ7W+tj5
l6s8UX07X+kC2Un1ujDrsHy2pfRKeNFvriM1U9itilrduBrhdqgwjDMDjNVD8Swv
cRBE6nK8tQ+s/ApDta8//10jFiNmcSy0UvJ3jB3Olbd71dRhKWTSgai9BpV05zwD
rndniY581dAYRg3qWEuPdnmD8sJ94lBM+gfpu+22fBeLt2Yw7B3+KuMn/5EWx/HY
loVbciyAj1YBCMEMmqdukKoq5Y/ErQL92iPlg52/EKzf5cIzksoFK00MRJBcGtVi
cTHHcF7dqwjJZFwiEYY7zAlAIR+XdWbOxbb6ozYXaM01zJiK9v0pePeeg5JJs+hK
LczYk4ftLvY9bUt0sIWqZ+Dw9nTZacp2TcueMC86naJDxz/zxyMVDaGoRoiJfKYt
lcsocKCxuYTbGyslqZGFHw0+s3tWyz2hWILT5z2EC5dpLh93bZgHXIwvysAcTnFo
SYMwkv1dppu7iQncrZixqlgEKuIVmitasWC3BtwBto8QzRlkY0iA6VgnVnk3FspZ
PZ8sI6tBG2Yq+lCIlN/JB5oKoSOd4HrKHfjQgWTzvE3eG2dp4wt6nWtiFDDS/8Tm
4RWSxMfwkZsGGCeO2fR7A45Pg/jKpA7WDZ11ybCnxgeUQdB0DKYqH9YZhK5fPcPd
AGXuLajkTYTA0jFpA/DMbNanVKSoDPEflVA34Lk8PgGeW63XmYnD6guCE1gI3Ad/
bPR0mJY5kJdkFWidkkn4PHOEu1HaHaz3xsoq1SvwQFyS/Kd1yJ1ZhJxSq4XQay5R
a7e2GIKtGeHNUcV1TOakZfGt7mllnEGd7/QWdLt8kIzuj6EHqYsbAxuGX7SQeQes
NzFfqBDeKjgHC0S99JqpcgMmz07zWZh3V942d8K2OAYNrNQLEHF6P7hJqydoSqWT
GD9Zu+6w08H5ynw8rfRuEdp7fxidgmEhlp6fngfGh11vXwFpDDNk1mdSie2+16Ve
2ABJFvhSJgxTurAHMsNcD0GzEUphbL8taiBand4SX0Hv3HOHh/HKBY/5VbTYF8jg
qqPCjKBBX/HZLyX7XXhE48GTzLRUwEuUpHaIzfqpCk+c2SLffM02tfEJGEgXdWka
m93nMJtMCOe0ivsHCft40kG5IUflgYqgx5Xo5qEQR+3ZJVU4OZhAAD9/56S6W9tQ
L5AOjDvrUeAESgtxCJ6/n3bbymv6whpNYe02b/wsQoO/CzkKc3dEeHHG8/gPqpxX
Fsr/AuE5XK0SW4V+HjO09VhK612MhziVNUkOCRdNe9uWiCbV+xUmVjs8gkzIH4XJ
4tOHTDYrFBAzLMDHRnMH1jWQMExZBNqN0vl9OaToFADAzdX9E+fKttoaoRz4Jer7
UzFlTEWnqR8CIc0qq/KJ1iTJHTohZSHulhrJepqgJCX8p6vnV7pcc5/J6lRF+PTY
kVBA1TT2p99FUmnIm8iqzgiiGZZOZ+nPuCiiKGu2t9slKScXNdXbGSAiJxSeIMJA
8mBbufX+we56S0GwMY9suS9GjFpjEitdlY0Q2Z+GQz7ou3Kkb51mdKPFV9GcBpOF
wqpY93NhE65lT3hx4v94HwWBKQAY2Y0FPRiLhiZW27mmZaPkrod/2OgUdfKeCE1w
5/c2WUgnGctGNYJMZayP23EZMA1MqHPKamFVrUMSoZekJQtjXM73rJ5Menojd/JV
Rx4L3fNAl8hpMtGNxfoKHTqj/fdK92C/1ssiMeDP4QODbByCxGJgkQc2DZ1iEHaT
K9PzafalIXsxDjLEma/peyofOkhZv+hKSyB8Fl6wEXN8RWKoKkJYH5wxFur4Daan
fZkgtTYBGuRjY2MWZJqkseNnIVHlqXCu1H+3XL8xAPHo+841u46cw+B4xtvpp+ns
7ok2vBgOYDRpGr39Y17cYESACpP6SVZLl3y39Ez0gEsAa938nF50fTF582y5YJMo
lAJFu/HXBgAhH8qSpzAyh7Atw99OfzRiaQkTw8GhsF9JMqV4ZhdhUnmHM0ztGOat
AIm40mSZ7Apr5MXiWy0NRv5Ugam9OGiR7aTY+gUdZ4uQCh6dcVNbSL2AjlOmRv/S
DA3B5LPVrqATafeiJbMCPGCZ6CtLVOjmH2jHMdAbksNW9eoqNj4SBKn3H6wAPFLs
3ZrKTwifahQGJqsB7/mYiV164pvMCZJe7mgtC3lRW/GVsP21K3fHwVeAaCiZ36xM
OAFEI0fYIR3sNxNGtUT2ldNzjsSVIXhhiHrUUoeYPMlvaZ2cV5gPi5l0JGKyi/YS
bAZ3AuPfUzgcqWEIvn4aUsPdACQFIoLrp3pfrCBqJVmSDxVqpFkdklvBSQEIg8fs
yKr/xJPgb458rO03y/YW9aNxbchObs/1mCDAOOKy/n/jaVKi5UELt8M0ubUgwuNy
DhL76OSf0mwNm9zbp0JT7CGpS4S8xbrX6BtexvH+FHpsNgwySH5EWcVlEBipa89v
r9dZs/Np51jZ6cHhSrer/qRMoIjwA5hDw6wQ+qT8WdACOCxZbVjMTmBct5kbaoGv
O6wzcmK2b5WfSiiprH8REZzxFTehQE3LTSZXspm4lZLQBv9jchK38Bovg7He2j8J
dBFUa+8jWR6ysRacLVZv+Oxr5ImOfF3joiP04QaMA/8EqDMXjibzkCbTjCbOHwnE
x5v8CNrGhaEgSZvOcrLz+xgIWMK2PSijUodOEVceFZ9pfFchRmF7tib5feIQZ56p
JgHpzLp+vHKMLB+bM4flxlBvKyLJ+O1pML6THGdLP9fhFA+JF8SExw62UQLwig0m
3w9k0N6nYK7DvMjAqQIImkJ9TKk5CXAa/AaLBfyotndKvWfDSRgyG34Z3nmtlYOm
f9UZ/qCpENof932XnSRaqPuEf5yNBUEIWxZrq1TiiaImaEZz0zlv3WiVkSoehhw8
SvGILSvb2ar5bpYpGhjAX7i4vuGWADZi4wCtbBH/sgYrbOmI4+56mDiB0OGtha8z
01F22EWc4TR/XDWQjB7OIsfdI0AXFOFZcqyt7g5njMLK0RqdDxs7CNjS1Gcgkh0u
OhjmEj0dGzI+Jj3P2SON6npW/Yfz5+bGi7HWqy3hQ6L3bUAtxO4rliKgrKpCD7d6
ScGSrvFB20K5T9cXAXZDm9L3OI4mM+Q1iA2tHwoQRpTfbw5dj/UTAqWSm6vYsRSU
QI78zUnkFxpd7cDcVZyTlpODwQ/2HLraBSRUUAlBKxq0czGS9crsug3qV4hImKbQ
sofpO+gT6VcT8BYWXRK/wK5bNl5f0djTl0cQr0fD4Qn56jCI4Stj4XZzcI1Y02r6
gg5E7m1gKN6TpeXN/JLoT3ATPMmu2VtDZkFo+gmwslNQtuK0jJAI84CdqM2nlMPM
pGL9s/IdsHVpf8h1vFKzNpZqxzYidep9vaJwmO/92+tx3eaAtUVmmIAbIUaln3RF
fbScUwRFOuGHOq/lhk3WmMBGAVuwJ1mg1Yj5PBZBaqI+x+jB+J5Qfh2X0PYDJ4XI
hwxDJ9KYMWBF2CaHEB4ZuFDSWouMPBPvwyxwBcWobbCKWSNggvGMu1MgOaBfsbsP
gJCufPXC7kJRsDIUJa8eE1HMDTuIckBoa3Oe8d8HxhHhtAMTYuN1LS1kt+sxDEnA
BV6S+8axmAf+2njsPluxIw6F3a4Xo8Wcp3KJ+nBrbt93DX3qMs9NXwB8dMOrGqxx
3DzMwDSOrXT75axGkgSUU9L7qGL1Gy+vCHQEBiR7NxZxv3iR8WqTl+BvPQ0+kNZi
WbEUMhrSMvT5ISMWTsliJgPAUogCVTE3aO0oR01jv1K2gYi6CZ8CwqbpxO/hVEKg
GV5AeTpNSxi2UnRL2sRYTg/tzrJcWg15HLViibbronmmEP3AVxMaEp/S3f7egrQE
v6n/W+tkaHndHaCW3BNRWPG7VnQ1oLKZZhvZFJ3B03N+vZJZurO6w8TquWMwxs0A
xyCIIMkbPg68Y1FBCd+zdayGgfcs23FiUXQWDmovrcLiskqARXjmTzaEgPFYd/lp
oivgu854XTxmNDtnnBRJ8FTS8D/9ayMMERWW2uopnVJLSHjL11rzyBGoj6U0H9K3
I1bP3XibS46XdEFhQ0/Wjz3VTQs73N2L9dILt1mnAwoW/blJojIlKDikJ0j9TUiq
Z9tzhdxk/zD1xRLFgkTSNgvcdaJMw8ydZzS3zgFWQXeiqljmiAVQ/9Bq/HDpfWK1
PzRfZMv6JcXsGQB7aGk0UIzu3SlsmLPr/o5AB2FAAMgD5hOPdFP8wyVFHyODAxd7
YLqxDKzvNCKFs2l5qbk1Hz9AADTbhVZceW9dNiGWH0vm/9vXlUr7mBl/xYWopqQo
jYOAugPKORA/1eJsdtT/gZmO1mgBKA56zBa0eoUQa8mSZuVqRqk++y6G/SaScH0a
hq2in+3ztR9gGLSJkEcG5rrswPBZ3xuKqBrmFJu3RvZVGJScCUA8ibXBqdmmODq1
Fj6Ka9CHDTkQ1QKf655CM4B5AS8rQpJMQrjps4AkAhMjs+Ld2KGon/Odepp4PMTd
vWLe2hLJs4rr2SFL4x8LH17xQAFnufyzgSswKheP8qo6kpjzGQ6HVTowh9P2BMn8
qMMboL31Amcs4oMD+YqABVCJrT2HOpkvuEMMj4wJ5wRlBMTLxcn8YKROywQoVNaW
mv6nJv1zZgdpqiA4eQuwca0a5JLljAWQWUmtKuCRx4Opd0QIsjAT7PuDZ2by7S9s
weaql+oAGLsaxXLRWra2z0TSWKPL2+RJGUBRglettRBViSeTSR2s+1BdUTpB/laV
M+eG1MOr+YkW+9UrCfUmMjcU0+26xRvKOcBAYYWqDfNv7sAn6BRyvkB5AL7Mzie1
HK4MS9C3OBPoqEV3xjuW9MIr0Y8WovyOBwonRRQQeT5QnsjXUKQIBEPH2XjflXsR
mY54jwskOKKSonAZfgOpsZArjyUdPJRDl7j35kZrMTVGOqBkMhDgPNC1NTCwUJzB
oanffduIvUSNAwYJJhQ4zUSvYgv47VkVj9M9YJzqvrvgixnGoA2sJFV0Pl+AtN8v
gUWKazXI31nDqod7u0zA7h2e2p6lH5RIVnYfEO421f3pqQx0tbCpSi4nNslu5DdN
3y+Si0MeESxs+BdTB9iB6x3wYb02bns3xz8aV0MDfb8MNIUVaIrirnp2qkyh2r/h
xdydwbTFy2bFSTkByIjUVd5/pRUM6UKa2iADzViPGcs/OpTHoDkQWucUTr3/iI/m
OrUi8fYYyMvMBe56MHbK0KoCXEDFYd60BMKBs6h227sJVHroZFdzomHVirbJq7hB
qW+XkIMqswEUCp53qutI5eK4GoF+16zGGlKKyR0W9r7fTD1zTUQH1e8/obJcsIbn
vFruJlSfmqvoW3+rX0UylbZuTtCcUBRcBc9IE3vjMxzTe3wTJrsMasmQCM19PCC8
r8z35ehRKMQ7NrLcSws0ZLxR+xEXDjph8ZZ/3GlROn8/6yuGCF4iTDWLiUwCEXDG
UaoQIaaLNSrbzunkUO4o88Yj/vdKSFN6I2synEy/A4EIf30MWkTlNbr62aBw4L54
Xg5Fvoh90GaBYazFLbtWHvr5SjCBonDzHhmTZ7vpiqB5kMN+0NBq8a2H0Vsmxz9V
cD3hQAl5tJwMvi8cqaV3OH1EEkbdocxct7iDXYYF0waLX12tVa132PDUaBfNQdH6
IK5ZBBA7JQRmdsAdOOwAgjexzDheOXbuKXthyNI5jgtNlPS1kpbD4FdlkG7rIRrB
3W7Aohw3Aw4q+19M1C2XdUsCcHsIzQxon9LaLHpuFjB+h20dk2wMY62BP95UudKw
LO/chgAmkjYNR1CGkQtj0Gl2WPsOktavxlhPPdIpy8GzO/fVfhIxFaZ++gwI/PuG
HY54YO44HAEiapIOjr8x7vQC3usAGSWuoFI1CQuFq04L3duhVJIQa+GoXlYrXwRJ
nqZam7+FwTqy53SgIkqFxDqzT2/DJK27qnnw461kaQTzaTLqeO+8c9jB23zaVhEZ
a9qwhTJ8qabfTbPLEkrqkqP0u06Axe5PjvMi6E2PBKDfkfS9f09ksPjN9AePITG5
VPB8KN2UhwA+sMgR3B8SNaQpBTHKzKePKSCtKXAADMHHAKnE/6EInIJLOzGK7d2+
9Ix8Uf9MxzjXesxhOzao9ILhTvHbQks+8azDV8SD6AQsBG8W3jkL315/qO++K/Le
kM6s6XaEBz9l2qPDUFKEr0ICISQAmZIBaaQRQr5Xs1gVVlYyFl/zRMTPsZzNP/D3
YoIO9opXU76jOzpr0y4zYiZifImUmPWlo7HeDfTofvb3BivUooUvm3Z86aZVfv1x
sPuz8svNb/z6TgnXtmsWNWZ33iSrF3xb1j+TYDk8RfbpasHpQh3DCZAFq462x71d
mht0ZEu3RKrKn+RcbZ9F75LXuQsweEt47XlQhKJiz8JH58FbJHXpq0AVMWAnHQv9
YQ7xWWtl2TvfZ7aqpy5xnCpJ+6UiTVnrArchIBBuISzAQ25M/jp9tNvQdPNkFwvY
qRHzOIzLNAvUkV677dfm9g3hQ+wsX6is68iIPs6tjNKhFDSp643EP33I3RVdS+7L
CFkolHAJPLHQE3i1GSXK0dCaxwC+8Tktx6jPbqdwvoFgRzSvR9gge7YqqsiXQzOr
eHbwtNDTNeXUSGff4NmuemubzqpjdQRWo70AW2Lnhlyl1C88uwFbxkdR147Ih4p9
gtNYigvKSBJVAZ5o2zMH/5lpT0hgH6JPvHl+7QqbluR4hDhRUWVn+d8bYzVUx+PW
AKd8Q/9HbqC1y8eVZA6hn4n0N4EyTC8BjAEYjjO+qGoFCwuJwzxSAQHx/LVKQs5d
O7M5J2p1LLSmorKtNokxGtpbdvkKFrQR3jxVeEDcLVV4BcwEkmkzFvBg8HqdCqlS
huyfsxi/JOllYcHJwbXVWjZH9vq01FVmhow4yUJes5A/mlCt8hcaeiGzQ+3iFYO9
Anrz94TX0cBzM3qh6kXeZzrqB2j7NHuJeOZB/hZLCwjw2+XjrrEtBnv9M8vPm4H0
JjLsRtoke0/tb3KbRzdRQlqCITjyJUQIee4hA0phIRkz+wQQcd3AOTkWVhaySWAu
TxzOOlnjUzEXX2Uv7EA4J2CIxtHahJK98IefSCgw5dXCpztQaXz5+ix7nbvLJixs
H3jPGD6eSduJKGK6e8uPVVkHKUxRvsWbfszqxHj2mPbJ0H5Xb85cu4R4qDWohC7X
nNyv2n3HN5CgNBn69IbRdMh5mfjM0tnf+KbASvdh8KOycoUm8gDnCYXA7VhAV6C5
MwxjCCNDgZhReHXFni9a8XBAEy+wbwVLIfBgoSSodfVvOL1hkGcRLeOAkJ6BWk98
cgNHCQHvpSu3m9hjRmbpBO9zlOIKhu649gamDUISfofW8nckVFobs8BB4KJm7IRL
75Yt+aEgXe383i+jjrTUs40xJYvkJfFH5bJ3h2NDRjmEZr/jFcIZ8qKQszSFnnVK
Fc0UnA9wApIKpLYzE6TPocOAvBXOya75ILhakWAs++4KNiWRkRFvzz5MguzVqw81
U93hojK3nsc9DLzUEoojOOdpD2PeNTdLplyRrMnf6fL1X2SRyAWtGQhcetRyNG6y
/joQLyrVck2Xt8sk+nTr2gh1H5eZ6yomG5y2benhffkxScEERTvXrBiBwkHa3QKU
1tqJ9MxkNcPaOtKBrt8xqrREAES5ryF/Hx/KcoNWx/IAUyw63IaMHYh+J5wAUIxY
+aDarGkSabguw78hrsOyDVMcvOqjYKJ6dTPa6oGF1EJZQIlnVsweAnqAiD3rcjkP
mKiNNOIn38EoeihAHxfbDxLulj0dA+b9W292z5URBM/hnfCVx3xBy6ghr1BzAeWA
RfgCD7uZIUl0I05OL+JIQubFz5O1MGnCIdGZOAIZYo9R/rJkW5zQelSmof30L0Um
B3shbq/XE10NIwjj7SsYdJsDtG1KKpcQAsBTrw36GAlsZst04fLx9ojpWI/yBQ1S
6WXE3+9QHc9qlk/izNx4Ea5EY/sJ8g8teq2krexSLEb6XMx9ACaqHjhrXl8OYthL
rcpO8EwLCsoZyrBGUR7rps4dc7+H48CSRAkEblqBUl+AEoJLirLRprUo6tppv7vc
2CTRaQmff7ntLV1eelsOy2o9+Pp9PJl8I95c2f9JSyddeyNOgMLAEKpOYBITOl/I
Mvk/MOk1MJHG4iiJQsl29EkC4Z4w/nuqH/WQy+M9gAV/KT1YyzF4eKhJwvXGocO/
VZglL+kFv5oY8FbKbirQgD04vU7z+iO4+iFfan7ENC6hDn1Hxxv4/yBENmciOlOc
tX7Ai1lPkdOdKv5s+Y88vsomCVZxFQiL06qh1PjbQDL0jBKK3UIZkomX6CMckUHD
4i1FYYd6AQ+friAY0PlqpaUabzEAVwvtrEGH+qny6Z1Z3IHVxyEaC6NNKq3QNATS
amFRUEGQLLOU3iT81BdFULVRtFNWkK5jpGZRHkm9L9/SHLKqTk77PZCWVJY8jzqv
0f8Ob8wbxovSR+ya6Ex1MozL6LnfKmFB18PQY6/BQAEUte77RiAwbqYDFFAiOVOL
n1LVM3X5Vns5QzhnLgnrI1AuTy3T29V0/glRN96Bcqm5DGScdCq2xIDEtdkyXgbC
5Q5lL254+9xN9XptYL3r1U4QSVLqR8UargIWJya4GotywGSmbXurI4uJy6d8W6gb
zmLlMWNEPGGuOfBr9rizZzFxcqs6O/Uq6neNTYpYjCH79o5EVj7l1WmgB5sGuqSN
u2UsbclipGL5i7RlWf4ryEqVp0XjT4C3yp78YymGkKTGkBhBUOo2XJrikr8M8eaZ
69Cl+2nvyROGJd/QJdtxkyBnooNcVgnnoswN4dVmEPA7t25TEILrnqckHy/qUcr9
ROb/PTja4utICLLRVwfuMpsI7Dh3T5c1nGUWI/ZZSWDStKedny2uS7Uw5ugrKMJi
N/l7WRHzq/sqB63ckvDhX/ChHgXPzTFY452ALhTJqYybHrrJkMMucBQC0Sfo4lan
70nACHvN9EemfTs7MtKt9H5ktHMqNlS97jwt7lWnbUYEugQel1NgQx4Efob3QHsV
EZCV+nHbsJGijW4QUSHPvnQjllTH+csRQh1rEMkZ9iwllsu2Wu8/PG8U/kSp1B6v
Lo4URX50LrxQRLfTPZO9AZeVDzJR9cglZBRqeWekbjGPnT6zX1a/CXRxdK9BX84N
yr2jhyijC41qI0/sHc/rqMez2MyUsbdu/+tDLdUWB4aUk5pEHGwQCXjy0sgWpknU
a+2OmeuRwsJOIqVLB+5JxlW0naMGRv8YVbl+p47s1WcMXXluUsKZwQOo+BfkWgvH
kHUD8vQs2Z9nScpPBihM6dzB80dc0SbN06P/eHKhHWftBHZNZBk0UXKO+eqybrtD
l+gUFO9xnFwp4vQwyWUHaR+QUMl4q7sLkzS/6nEI3Nbpfqy6bFSxgLNpQwMZdAS2
m15zx4jr8j19s4oQ5SQVQCezpWXDiGI9takpdJi55Ene1oc2BQe1S1mAZe8KO03a
84SWItcVqfZR6qZ40ZQklVBZl2fHweuMGds0yKSnnLPOSwlTRkObZ2lt4dims6NE
PFZOjejoxr3i9S7D1Eg93JorpgujTW1jkZfTdIsmrFBuyk3DyM45GGYqE1/Woxrq
06nOwxnQr6Ubd8V2sFVUAHvsfebdJSTrbQKqmwq3oTxfmfrWVuyRItXtyxP1WIwR
jzLqwnWOF4AKcaW5N5w5D6YNktgeQlhH+YYNrMA/zw3iYAJbhZHStn4RQ/P1hbzG
Dh9uODUsUTrGb9EvGSS5zVoN5SXtRBLHk3rHfsWaJlRrPAadvaCnZrykj64tA++S
LJ67u8yoLx3UWPoRgakvX/zupu3GAMMmF+KJ+2sm7qAfNWZ2wuJm4TxMAFqR7trs
pYp0aloqF8fS5PfD25zBHWAT5ZuznBWFO2CwX+ARf9c3WgL+hLb11b3yA6b7ijD7
U+mH10Pauwa8pyhmeQk2qp8G6552hchw/u6+uKCgWQFD+I2xIKPUwjAtK7cAb7kI
ifdbRDB8SvTtdKWxLaL3FdEtRvEFf6lhF7otGL0BpuM8Ezimp2Hfr+8BqzAisEMZ
CBo/1G60b/PMyn+Quf70wGZquS3oEeeAT/7VnlNvoHbCRt4Q9OBt+MGmJxJNDMQF
Kyq+8TeJ20t4PIxZoUcTdZKDyuksnwAK50EY+FZhRP/eUPa/Z5o62p+1sZ5jmowO
u7XG+IXznmxRbSrei1SzfAfV1cAA6pLgtYz+qR5n0gOn7HWFtNaWkdNYoonb8TkA
SkZzj48PsDrRwSro6VsID/4X4JOwGjpz6/PqAzYBC4iHQ2Vr7TEVZ1+3T0qcTf0V
vXvcmyRTfGmbpXrW9Sz9vgxjTCDM31siRIgWLUPHW2ag2CVavKBtnCHaMp5nlqwK
e31gBV6qt+jfQ57A9FqL4zD+qw1vbq8AFlbKS+UwKW2NEBte0vod0dbs9dZEMGtt
45iIuZGOVbqaU1pRSjHCGN887+9UzmCqixI0n+vDLtOkuIS/2/EHJxJnQJjON8cQ
LyfBqrBFnxIXUXx6lspKiaqAG4SbhINomnAGTKWuUrGWYl7dbcFb39sf1kzEhvIB
c8aQu/YIsetV/jOHe4D4MwWITBMN1FzSwmc9L6ByM9W+De3Ul9E2Qk/s/Yswi081
D1OrVr/a7QUeU9acFmwEJJrZcAATtwehggB//mj5kKrVU56Xu2tBhlzUcD6q6rws
Fk648BlCYiCO+MarhP/JtJtLjWDxtynxo/++cpn74iDCpJXUcfkYqjnkCkyHCiMX
56xk1Kmvo0XvKc2JHkgcGXW9etQ9h4bAAJi2KppxLbOuAWdMCJu9opZx/zEW4Qt4
6/8VZxnIZ3xO3LwaSqVx7j31F6ZMgcuqPSQMAdci411ElILXO7XzVlb0/82OvVNA
/ukcbR81QAqtZoJ0n8c5O30/ipCXlFXbtab7AarEyKt/GvTbPsNIWjCR5qA912qR
Nv1mf7rSeWUCDpvq8L74sS4Mj5zrgHWhryhYb7EHiy7HE3Q8Mtf9xFEbKqtTnZNR
OM1Kr93HCA6U2eMbnJu70xG8+1EQUT2VxOaoISXfshxy9mBUq7vbP5rHOaca5O0S
xrvQdA0+XIt+JnKBtiQRwlM8GDONWusGOE6XGyc8NJgwuB0gWSnmaYi/Y/L6YWOe
hsxZvmcDNk58wS+4Lbdpdh1Q+64PY9U1HN17nqfRbeZM2muNgmbJrODzAzN3QUMX
KAgY18B3FZdbyTji4NpJMZrZsQ0OS0PlMpiOYb/swo/PmgrDiGP/67OeMFH0oEYx
/8WHWI7Jmml+5k3o/7UMV/keBA8nOqtOAACmWhcX7SYf+0c5HkbO7B3zhgB71FWT
IIDcun4O07UICXVZcQRCzc/Yqs7EXQgHg3TXSLuMR7ZVHrW9Sl37hCn25kkkc4d8
XcPxySqq7vGOgPYvvTxrl32kHhEyZYZLl6w8gIyk2fuyL8eZ6G6wQWrYc0ol20PI
M1HbZIbcOeXqsE+0Tpp5Ki3y7CtCZHdtp5ZmLXqBoLdXiNkqdYERD+d9nToekXL2
CQ2sRGV2wqXAWNKokQvm/ZxRpCbZA3hq0VlFhlzEmVCsgGJhEG+hlIj7/znijxPf
Ute5urpMvFZi2LPh7U57h2RKwfoTWYcX55++B0Dv6vAiBt+vUEfsILBtFDfhiXFI
VBvgbJd431A66l6Ltkr7VmOt9gXDoxmhO3APr3omUitaxu87TjFS3Jrd9+3pNPi5
HRqOFTFhErP+W90hBaxIrJFZrhXMpBOXTvnUWzgJQyoQJzhSB/3suDSC+8hXDJi5
kTfAMRAgEQYYstUSeSuWeivpjJ+gIk77hO7VWrb8z4CbcHjTXvl5uIqKDsdIRku0
xa96nDuPSDOYvFvzecnJGWHDGZrJZWkQxU7BmGFQ8zNP01p6BWdnTT9RI/IrGsEu
ERiRBJ51i1xGKACTBJlaVVjQC1ECxTY4LUfVFzZEk8T0wC+ghtr3whibJhOhbGyh
8Xm2IVfqV214wXBSxNYsB1PTO2It9rgA3Vb7eB1lZimxLRTAYBVb5uJCw0nOvW4J
RnaCSngTy+7koCs38nHBrV1YYvEkvpKaGB4/melvNJFK+qdqV4bCc92eRAOwjsc4
IJ2sxxR8UmszIbTxp2viTDOcO0Gi3BLNzn8hJWR1tRFcr1xPClFujctVZh7bmkwM
8CNVV8dDJJ1cswq3b1kQKTkILBUKffn+KpJafTYAdVMX91zbZKWjJiJJdpgezmFF
clYJtqwj3WrK7u7Oh4hqM7DNjeuoJJJYZcPyvU08wDqSh+U14OMPmvdlFSy2vq3E
RuzozszJ8x5mVi1Ryp7Iptum/IJ7aNv9lURWy9pUUbBsTRpQ1jnJwy4p+/MTB38N
xL/79985+oKU8OdplTlFW0kxq3OYreJEenjAZa75XObcc7BDgc5h69Ip65lq4JqB
SIqVUP9BB5OSHhxz2sQINi0h64Sq4mG3N8LYTC20+tDmvX3IAbRbpnALBQXfAisH
uuHLCaWIOJNpn3ZLwHNAlQJd37Coai/ECfwyPFzrXT4+B5ZfMibayp6JLbH8FVsp
C5D4okAgKiBXuk/L+fuxSxfDoXOCy5620Rmv9zrr4jM4yQY6xMvjc+rC+F2K+i+s
OBK485rmX8Xwdfflfhb2grtyAQP2oiGuvvqAqNkhzbeu0hk8hLrgivPQX1jlCE/6
nFhyu6PMGpLHYlnCtVMk6J8qaPnQKptlyIGVW1HhyFiNkBSgJJsKY9TFpgTuJhX1
CCG5vv9QRj55U6ElOXWPpsUdfQrKK/3mwZ5idtxRej5w1R8f9Zz2UVZ6gWzYC4CW
6tg1Z8Wdbat9bIurvZ2LT+zkCL1ESkFlH5lGYVsYABy73Za2xSbNQ9tmiZWrrymZ
eThK+Dbw82j90Sriy2Uy5cDi5J7xelJTkkOexwkTZ7vIRZPizhZ0X5nN3DKqzi7y
CB0xgKhvAsoCb+r1upyE6KSVCRKNk9n7K6c0gLc36GvTcApmfReHPpyv6O0TsXbs
uPFQbF4Ysi7OnJp7RQB0ZUrROeK41Cl8RSdqDJQ8c8lGjNy4isbt8dgkZoUwFnoN
5qEsPXBvzpyTVwvQxsyQ3rLTFUnVoAQcVEucXod4hhU/NHCpDB6k0Mr8r476M8gb
nOwjxvy4zl2Y/fjik1rVTPUkZTTC9M8+EgE1oscARp2jhT9qKzOv9nue4puEDjiq
/wjLxWJegy5FtNMsne+NMfMNlhXBja8h8AlGyb8wsb6eM8BpXAlzYaiCmP8P8K+k
m+eGYzNyZovtZY/W4OBdSEXfCoDWYvhEyMVa1wBogR2zXsvoLXyX5rd+wk7CH/ud
CLG3Keij0FJ20giPeTz+6Oi0SbboYnfzv6spW24oiZr1CnIJ52VhethsiQJR+cZe
XrnK3kmwYpcN6ae1WMvfarCOmz6Afol2ieZTVSQLLuFt6sWc2VA21+Exu+I7iUBG
VJS4l3FzPwmefcS8oG1rrW8nLnVv0HUrDnt6k70pOVaOFfrKZ8LOflAdaI/vgCgo
YA0Or4GNbPNPZNmNCEQ5JgRFIKSUkhMIWo/AUOU03f6HyQ31AQYjUlUkn19e3Kya
Ab9vE23a8TNPa+Q83FeZD6EDgeOozzWdF9R8dZy2UfXHQWypxKfzW0aRf2SCbw67
2hWD+5rh8rsdbA+PTdaGs3E/yO3BvLKfy7TQ2MKwStulNtBS6T14tQGy92N8VHME
51RT1gaA3wAzCB6qjOTXkrxRHYMKj73pgoyte1EVKDV5PuH3U+F9OxboEjJ6es4Q
D6wvKqn5/fXNRUth77y7DjRfniELrQQHsxPgE9Mj35KOEaoAKbTEhpU9iKVKfsqR
1BJUXOyPwKYbPQAMREC9gFhe7IexOQQinJclrgFI5wNfm4fCixmRT1fi3bEIIzqG
PnGRq7u9IP1/1Hp6duuUcv+IM+NI+ouvjcRrwOFhjCWpor7t1WvcF0VZ27OOX8ug
tmAY6ho5j8VjrsEZ8W76KZkjv0tUsawnw0DwEjNZ8NzglmlZG+lJwzroszYObEMU
XEwxM8oztlmw/3k9UQVZZ+VtSqN9Iz01C3OdgisP2x7oJ8T1T86yDZ6s+rl04SOP
Z/WUkDrsP5A4azga68J/+Ho4Xm2SFu4zIeQUcaOJ0HfWvczb0qt5XoFQ1fCe28rO
4j49cnmZC83siSvnCeXy8kk+otSquw3TfOfwI2KfQJ+KVWpeIBqTqDX4BDFxIYKW
oNDj7y8HVf9q1mHnMabXNQHUQaO7PgXIv2+GKevJibGGeHgt1vqh735vk8d6bGpJ
V5WOXWqbqiZHsAmyzZmsJ3wsspdAVfD4+xM8EYwRQ+L0fZwCq6Po34c0dCfC0YLc
YHWHaFIlBte1e5eCEPe3uaHVC4eT3bboDJGwrxPAuK1YIMXRjjp5Fg9dchpARZ49
+G/2vxjPQ80xiKOQ0E61Bi2NmqWW+JMgUhFER9xkU45GNChhAGmpwuqfn4ZCsAYU
YVZRUPu5DOVMhIUXKX1dlzrybn320H7unvy2rqjMKEH7NbqdajJMWKGPT6CITS4x
YGV0G+V8zaze8phWZ3x+7iEq2JyxCZewFCfR6SfTj7KK9uKb2qQoiIvwxCfKZ72j
jeyE4Ak2QXC4Uh7yvynRzntXaixn8Xf0x/NTZsdUJSf7uiGI3lt07XdyTPc6sABi
qVGO1vN++qDm+Fr7HlUPSy7PrDLRE+3PfrGiytXGNdCiWHgUYWmLUOi/hMhPbpjs
Pup5Zh90lCs15zEbhiQq/C09//7NrH1yBK8TQedBC9J6DodqSyHb7HDmItyDTlI5
qWG3Ui0Zuv12aBWBegQTAfnnSctPK9Ry79hUl/GzUV0mNRMdB6OFE2+ek0JXJuN2
JfrJWtU2YMz1zZYSUtv6wiy9bXIN/2iXT6zxMGQYJwXP0zedfvEe7O2s49Q9o4Aq
xXCni443EFPtTtTe6z1fjD0F9sit3NR2RcEQ+ooyqhMG4jh3D8UVXa/gF+ld3iSP
np03wrLXcvZravIAEe1CYkVXyPIlaxpM61UPuanJGnrsqM5KbU1LTsAUagnjEp0C
toopORK5uU/q3uCgGuk+FVh0ZTsnwPeK6GsY/lNTHeUj4oMA00RfRCp4HwQzcawx
LswWyaWz/rFmokRVg9WQRsUg5sKCPSVhG5XSpoY6EjQ+6AnHuPIfCmm87naCp6/d
XEKt+24JPwUjNbH3T4nT1JABdpy3jgwHtiBNKOBZ3K0p09QPPE+MFVPbF/PsmkjY
rjoWc8dKdncfTu1/r5wZfxVzWRIsHpueVUj7lP2sMudwWYDeV+4Gzo2uHQmBinGH
b0bc5ly7ekjDuHaTZ1+GbaYHgmFh3s8xPBlYxBq7AXGtCN2rCzkszH26GUQ6SQxC
BkptIi9OyY7dIzJtx99cKVC5D0XPeu55iKWm6lAwaYCoU12jhga4g9lDiS7wMs4l
ULWIAdULhkA1r5HFsyK03nOceCfFI1etrGDhyVvi9JyFe1H93LbDl5J9yeeoGL/H
Qae1WMVGDdoDQ9KnZQ49QfMOll6UXy5IJYWzv1Xq++bdJzi+aYavMoeZhbVAZaCY
5kJtkhqZ+OrSQuauPqn23HiduaEnTOmIWYlsGJRpHCi34Qa2BT2roTAlEwvucjMM
nVjbMOYt1b9Wp8VGUM6Zeyc/z2wLhzti1fQyV69SPaKtKVcZyUN1oIk56NTfPFP5
T98UkxgCZSV/MhSV/T3pKUAyfC1mmo6b0HuYR+VoZmDlrNBvJf+o3d8/pLA9zSBw
42h4BQJNF87mpmv3UxEq7fmdHZVwl4Zmp5gl9oragfrl6ClyY616OwH9J33Diz5A
mHnc/M6FZ705l6TVPnCDs442GipOMAqvOVxPpWl4ZfDDUZzMbQkS8zOmG8QfIzUv
eGIxE1uJq4ixd+DGPoGH42ykigkqOHC0Iz+MyPZun05Vkw75PhbS7rlPOJu79mnu
WI4lmHZhYzLSYLJIfb7o839szQxs+WSewCFgaACGU1vCcReLW4+4lrllKOPNP1Xc
tUXeQL4pfI+Q2XImh+qlgPQ5Yhs5fdmS8xtIi+MOKj3b70IfuyzneEcZBt68tJ5j
l0+51gb9BaobJnOnLV8deg0/TP45N5O01XW1xi44wk2CiXM6UZv6+3yBNrH4/jQW
Dgo91CrWO4WmxLJtHMIHgW93+V7qWMLm9yiqcBGELlukA1e4yBCmwaxKmNi1KNTa
B5LKkTR+g/3jfD9y+gzr2hd+QVDy697Rx9xJn3842dNuLNLUN51QPYaC8gQdtfGH
dIhb4HBjFYbIkSdaNA8FoMNyx3s/B63p61EvlmGgln6I0rgmpftUQgw9N4rCCuAn
x6EOect/lFNCHHnRCRs134OV3Rw98YhHSbW4G16jpRUU7zOYMdJr+PoITlN70lre
4qu1a8wDuxQ8FeIR5QihL5LqwpmAz5bW4VA/qKg36FJZ0+9XOOs2O4FgCNps4ous
HUZd8th703POhqccisgMRV35GibAH0HVyJoNQ+e3jwjaN3/diBOZPa8ATUt5HDAP
9urabZaH/jTL9lib0M8BCJqMglqBD8slVt72VY6kNyxSPZ85f9BPBAMF+ABdcO9m
585YU4DJeQe+6M29MKYa2gAxPFaQKMx7VSUyXqSOenPnJo76hb9Hah2R7lmizoT6
QWXzwD8MYapd1F+fbSSqq1CK8CVnUzndprZ3Vo8qb3LgAvg7QAzdRTyt1aqjukEl
0HX3B0+HfUPyTFGhNKRquM61TUS0A1Ps0BwxdUXI7A/eHGCqZZcIThcG9VxBI88f
b4uRH2jAdhJIeiaTxjabiOgiejwO+IT9dOTJeGc60+I5iGgoTY4yLPJRAAJVHYxP
v/3tfOKzdiNfW8PBFunX6Hy/6gv3meL7hBO5aqEQZ+FllZxNG3h5SyvTzcgMzoYy
0X0RY1uyz5zMg95Dtj9/qqi8280PCv2QU1wkYBhblHSDHnobI9Ms1BWLSpoULEnr
XVNJzmVIb814NfGPanodIEj22AZsuRAecOqgHTqgn3bjEWwuEUxqBDVZv9LhtqiQ
49B0qAxROLOghNawt1kH/VFM4ANubzA4n/x9j3Su+K43tbPdrqRK13B/LV+U17gv
qdRL8EnzE1dsBwSG4wJLCydhEvB9f+ICVlTUPuAd/Lh93Ah+Jaaxf/+UThmvPpLY
d6elo2gjJWxUEWDmYqNpB6m9OWs9Q+a7M+ahKTbcXoK6ppWJBNL9Xi7FnkmORQxE
mqYAOEdgFI5IX8taIfEPJMDBOspgkEXNx10/lISkRcFgCiI4CjGAauGfwsmFO1/4
E0Q9ziRLzjooM8VyNA0bDOQfgZOcK6rP36XMSKTvhDf5wm50zufDjBK+bV63LAjd
+v/x/a/0brKYzAE4b6vwhSZxWNXiAUCy8x+0tO3TUnpaSfwRAQqc6p6zMMX3LRsR
Pjb+GQavQnck85BSdYxL605qKAMbQ5DYnrBZ19qnacDDeVl64L9X1Kii2oUdvpzo
4/rLhPoRxrExgM0TtyGE6i/1A6sqR1HFXEoEqvRC3gLmkujIi4s7iBRMONTVuge4
TDvPyzWndha/C27fkwTxVpkY+SLpIUWWqxRsQUFaww67HzmlRAz7WJMmYuTLWZdv
eFL6u7WtjthiTAWeTn3hEqO6uNDAqs03490fWTddkSpPEcEg6K0WMAfwNYw07/oQ
QJjK5zYn6P1Qi3WpPYfgP0L0Ua9TWMAvtnCXfkxnrytJQqYK9CuBRjKdf2c0OKd+
AkYeicu2A2xcKi03DbTM8ovTZgzWmZMf0xZmhM6TMClpttheU5jNET4OWzkq2yHP
CCvPFbnvhP8KmPZXDatS//We0V+QFxQBZCHzazkaC1XVHTOt02eb3QO8FGIuXhNJ
A4UPQNEswNF1JZ7hSaf/KVgRbFOBTv41/MZiE3bBQthHSPPlxKk60npg0QYEcYpa
GexokmP9+w2f2D92QvvI8EWQ0gNAlDkgLaGI9ottwJzbh2sDX+7DHdhlvA23avTQ
P+p/HpWWfHQO7I2vmNjqMXBXMiE+JnOdYyitGkSXEDvrWkzaPuyGXzEYYhOKXOYs
PFWs8f0Tc4eps6oIz/iDbUA/jQOCO6IgXhBc/f0JrdAnQj2oIfEwHCxCpg7pxRlc
pWBGKVNR9KVLeh5sli+idXR4fRTGQakCCdvCDnN/1tujDQz+Vq1m4dCALp3fWAvl
yWTYFGsu+CzdVLP3HuxKb1OLCG1h6b1kFx5h1+mCTPlIhR+CY0YpZ6SRR0iCvxTR
55dquB52g0qBzBvh9ljz/56pCrrGur0KG2vH6I18k+yuPqcijvF+cOz5n2nht61+
ZJGcf+50sib9dn76g9xFZICveXjGT6l6EbpElDNVBvMWYOPTF7yi9rBQ/RNZn7L9
ZbOE87HGn2uaC6FTycVnLWwmLUumEN/zF0fLoGCb8b/9XmgfQYvlCtkqkxVvUhfE
lID/2EC6z2uMAB6FU75MbbNNP9Baq+l0ntXrh8P6lfkTfeo2RM+az71P1W0kioZo
akqpduQza9/ImbOUkTXXPfJtSLS7/HL3lIAq/vn8fFquvZPNOyAu2H88g22tsFZR
mhIl/m/EFNmvLMg9ZvSlf8bNaCBsep3/hO611XvnfG4pSAX+t6HGurdJl0bx/glJ
/AYQgNsbFUCWd1ZCv2gSjCMKG7GwCNAqkh09BTqq7zDdR8fu4xLkn9YK6U8meeqt
7jXJmrBHfij5Q+Bw8ipsXF/n/kc9VJvZWgUZiomdorlw+toTnX+fIqBhuzfd7bUC
QotaSoI5rv7jFqB2JNPF/AB6DtnAotUhsudaN/rfYoL47HEmsvx4TirdMPdO8Kbx
X1R/gUuLFoO707UY8WEsPEiXQDtwJ4ltJXykMWUGVrm4m9VSDXqlBY7NJZQMP6zk
NG7keKQkaWaFf22si0stCtZwa0Pck32DVUx88vuofyZtuBxTB657f7yRuqOcBvzl
+zfOaAB5guXfTzSMD32PauN5EUnA3C7KbWvaXzYANTcyWyXzwHQK8QU06zOwdBi1
TKDsFFRI6iRPg5Hha+eHf8ZiYaG2DA1k8VD354riBactCKbqFlB7kQkRH3GYlWWp
Ot4//DeUu0KlYgatLM2YTOhrxZEAZ3FGwXKZpV9WlwAfkDkqT3CUNnX+eJszRTno
IncXqdoUUQZkR+kcO/m/F5GqwAjTCFcnU1UxhhOs9VrKZ6y2I/vvur3fZuWKCx0v
rkKysX2u1pMVK/Q4Kv8igOarePUK1UhUY1VqbokGB8OrVMjVoKSnkbbzojdUjYXm
jn0RXbild7xRfdQzYP54cWujODRY2j1QipbWCxGWo130dY37naV9Vk6slqjO5CbV
TFw4+KUu6Ymw/4XMyFqz3GT9Ypyjy5YL+tdgM8zoHZTwzErbikdp12gjW7ZF7jyA
4ooU4KbolBCPh2MIs5t1zDGze+Iq2W6XPvsL3YSdQS8CozgKGlW/RMzJz47xATz6
a4MAhE2ncgxstDk06+Q3LoEselDqxCyjeN0ZWkeXEcYOEcZqvvQrHOAV5olnG2mm
FrUPPs7J2tbHFAVraATrX54RLwEH5EVOe5WomY9sztt94rUs23M2q07VZQ1WNd5o
MWezME4NAZab67F2RiAvsOHcI1e3SuUzZ+h4YTtv/THHiLhBlwPeJwwDux5tqdfT
PpiYty02LR9Ef4st12tKmocP9NSsYDTSo8oOxxwCTtcdE8xkY6W2WHJmmHb7jAKS
MeVdPx7owzryFaDpckXBjrwyC1DtGl34GAfrcooIZf7yDJH+C6JABhq7NWghUWLU
yKlPnLA5tkfKfBsWTId3yVNla6VZPEnKh/IfuLOgqDAn3CAzWK9cTWs2TJK9xmsn
s1MmBWrnpsP598XGgvZ9Y6BgymtWcQsLjOMA6YkP+nyMiSUkLOu3mTlvmgw6UYYN
WP1ESf0WZ7K82ZFxPTpH14eNBxWB6D5oBUpTrKesp6gSiepb/5TDF+CEVqTn3ali
IWGPI8tPHkmg1Nv+6tW1CMFU3EdarFfuDz6K0FbD+N28HYo86YhqmaiiK5GyVeym
5DsMhCL1Zla677uDQ0xckH90+wzRiWvHc0G0FfmhycQ0gn7B9OtxYb1uN8PZ7EXA
JzX84tA5P9Mn6/cpesLw3AL5BqI26Fn6URlAuFR3EhPBP0Os8oSfMwZH0GI1mCEQ
rfwfLo1dsz7FbXloK8inBGljVbCYLHrw39gupdZya2JanpEoVoATWRdQ2XkaYU0o
Ds1G/dvFE09aMEBdXy4zxysyGB0CCLuL3xWJGp955w/tPG+5u0SSF/XfoujFhgjH
P0usv+0vlXPUIyvvaI0BqtfdBGSqq4ybsnwCPYVF6o80Y3twbMjAEriKiXNUDBT8
gx4h3e7uzWdXymq6oMNrB7885BHUdRyeVysMqe4ba1gNdqOSiw6qjaRoN4gC6lou
ecNaZMSwSOAPTzapNNOGSxi+7Seu5mRF4j/I7zMJBE1YTRnjIe3qHr9GLQx+uDA8
OWEW4YaZ34+JRTvYWprtV3+WY4YGeSY/zZLx9Yj38ooSVnk+PTJ8R2IvXNQyBgso
grsokcqfwYxjEBk3Wymmad4ISwvtJBpOEKItPFRgLGPNruAnCqnYUpqqBZnq3hEk
vYWyguLvTUza2rXeHMEWZnPdBaXcsIRJ4yovO8YjjkZY3mkIQxmTP3H+ExYo5Rrj
tCyxq23jHACE+pm1IPN8V4JqMsgBlCHeoorv5hnkNTnlPezB6a78IQPk/twZ0eCt
FO99a2M/JBFKINESN2A3RdQAHMkx7J7OUEQ83kWImgMmtqaYeRikZxa8Jy2ezHh1
CY3SWoGvGbEW1EgRssyB4zrHWco6ThsG4qxVjor7C8t2j6BLdUuY7IFMudwezMz1
qngXtAX3z24coKf7fhqIo0Sn0GXgrPXmA1+ASxlHItVTE/N8WyOadcHUIzBhtlkY
StxHeWdd7rDmsRSpxueuPcf3slEClE4ghnA5Sot9c4oI8L2zXo0YW0o2rXVemOjR
F0urQAd55w8fQc1zOIlMztNSuir60eW1smyqzWGO9b31l3T8I84Tu8vRlswElXph
bXAHaKtxLZgkKsxblIfT4VmHfa/RE0q1d16AK083BdjP7AcRLXMvimQgpiEOE3UH
CTkLX+N7M9rrGlVk6nSoFYjAiinh3Tyuy09rCHmv1e7o8E5PtWHZelBVXuyMCSOY
005twyuucE+RvtM6Xi6HsS7ZAyjDZctAeDKs+ZbgI4weLWoH64amyu7nmKvVtVRW
xkAgOw3xDbnGUPFFDb0gG0S7ef5EVe6Ro0Nd/NURWV2/j8TVDvn/OUbi+4VU+I2J
31S+VU4oco0oqYkHhEJ8uCFlxDmLaufWvPAs0mgWPZLk3gF1hkBYdMdoxhdf1wvp
4r5L1t9HpJT8SzyhCwi3zWamAtvh23wObYxkZHX+lD96Ef/1HY90ZTN8O9lnXh3m
al2WcHCXpmuMJ4o5sV/9hgTxy7tvUC4EugkDR2tyDE995W2n1S12TkP8mnmYiJFz
nonX4DJUBTHsbbsaoeUmUVzE7ontNVCkr17k7TgDomGEhuap773F2YZoX5hiSF4r
qXaLo0XCfgUTOPtCPJd8kDGPAfq12hTqCfMdT/KktymkpeE+hh+Xng49CL32tWk1
5P5PzCq8Rb1pX7Q0B6fQq5eWvKW1PMH5P1xVKkjyo/MMZnQvNwN+REH1vTnLEzgr
pPwjnFNQxNRbJeuJiRRNGIcJMpg4ra8U1LTpXIJilyL5TNZwm4ZHgbMgFt1ht+GE
D1yYaojecF4+cJaXfdqdgHG0vdrje/M9HnvBLzr7dfIlW3ntJEM2Jw5wM8XwVezS
8q3Th8hKwCTLi63Auoj494MFtdpXVL/EeMSfztUpM9/J2gSeKsWk7x2iA9pPkp2A
iju4IqcDhB75qT6CzqCnaQ/3z+VxrtDPXiuAxOh0GbKttIx8QFS1qHpcHqp4x7AP
Sz/CfK1OEH0VL/wXQzRlvlz5bMM5HgdKtMRwv4yuyeUgNai6S4S0dgB/yVc0kgyf
e85l8fIpDNW98xs5HgPZjMdZUimxzo1gwdJIsQYbXE7wh8X6ueFUKWCG9+9bwdo1
CYpj7HKr9Sk4KXsWjV8e1+g+jTroNHgSLoOa4iuSb0nITZ50UGPSUaLd1nO06WEH
YsSD3GeTPIwU6DDbP9J+B1CXn+vOnN6eNZxzCXz+6MG7g+iubwyGSQCI+Pur5IVL
gEW8jx6Pm1D0SPuiw9Af40UbNEb9Sb/XhQuNk68Td8TSYRhYTczClF1x+lUxu7qe
NrlW5z+ls5XE3I0MkN2wT6o5+oWKlM+RLOlIVnhw+2xGqFjO2l2TqwAnNnhXH7Do
F9Ymb1Yjhw7XfVLOK6KfbNser6ioWMNT5sLDXnETfByi3Gk2qfK5XQ8DfAhhRBqL
DwDABoEv9tJBF4a0s9OlF8xqwZFKduBNgF3xG7SXCJ88S5H+W8hKBeenBdHN/C2l
dNOTaLNL4gBK4qwgkOSaFz7jorNc/m0PXaggZMIhwzbQIDjRzVVTslZyKPrg22xe
6ro2mtFhYrs46vgzuxqW6v7kubvbH2hvLahfwuKPrJ8qBQYWmRfDHUETmu8ty168
j4N1vMX/rrT+v9UxXyORvhool3IQzd1KTa7/28qWHLSJ6YRp8K2I+Vv05ONKRbaH
fUexlvnGvbOSYat1I7nfBUUaGo3FlheaJ1lvuKed9J5YIR0BrHFfx/jf+3TWOKUQ
Acszm8yB6mujLgIk/5t8/zzxum9Z3X7FvUpcNTTPUcHisVPZU3uvoK8gJTWsjANp
xSbcuKf3RYsUoKSloDqR7q7AX1twU89yr//ghuK4kSXLgVTbV8fE/2jTBSbB/QaE
DZj+IIQXn95XVqIIAKnd+KO363JGFyIh3S/1rjc+6jsiHpDUgdFpz7yviopJ++8v
rGYE/agD5sy/hmbLG/wa8vofhfwE7sDCY4Kmyu0lmjrFIZ3ByZXNV3X/JzGE78kJ
5ELpqbNh7g55nCaQs90r6Fqf+T1jNqqdDRdzMaL9rPvFQoyzi7PwCo+NGaVj5IPl
HBz42CIt7IbTH6oZnWUWKWctv8HkwEgfcZdsJW6VCpP0Kx+32l6uf1vMjCwd7kcT
rN9iV+bFm7Ib+27bn8z6Sj6exVVn+T55b4KvLY5uLp5bMASsztmXiSrpeux1rLdQ
lAk+EBX+fYzHf+aXtdP3/ijHFvvrqqNq9uqA6Ylcv2/TjXaHqMULKGE4ohAbRyse
X1dDDNPQ9Jfpn73uSK6PmG5HcPuPQlkvO73LkJaJuUA8PLqHXKJVMN7Gw2Jzxa2M
j6j0/3aJnIDheFDT+50rtPc5FLpMzOT1B3JC55eqcHSUt8Y9AAcx7wqByaQs2NqC
actEvNEWqH6myXyZjO6AHVI2hBUhq1xNrJxWV0i7FzpyuRevUdnL6WfmLCF4wxLM
Iz4NLxohcdM0e5/ZjZCJltrImnoDHKoW+DQG9hU46OV9FMYHMKXc/JlfsoMtSoaE
zTHf5IhwmOfZG+b7Bwy0LwlEtILjRrBXQlJaEogXTAf6w2G/SEn+poXhdYiqBUtH
Y5crhvel4/4+ZoM/tJ8C88sn0venIFeknh/ueOrImtZxgMSL/+tMc2nAonhxYQGQ
X3aYi+72xYsqHWWKYrj6fJ/trYoZo5s7WrsPjDucEwGIIO4cjrUop/5xVHs/5fjr
RF2ngO+zpIAaLlfHqKAsDV7pAC5P5X1giMb0/2kaVcczDv/tfqlcpmh/VasLo/vv
WQYRtZxS5Y04U9lgCaTJTjUY1gRa/vK1FGt4dcYXmbp+6JUHVXENQNcwrp3xFpHH
+ESFgyzusU4kR3n7eXTTLdyHQa+D6xObMy7CzfEUbrMlBPYfNeeC2JF/+PLRCrEz
v0ZpmLudV0bVzIoZurorfceLZ63Bxf8K1lk4krelS3gQSF4GwVc7WahnpN+Il7tF
YrQU2gK264pZP3hfjIF8q6sqZeveq3D/fihyYPTZGxUVaST7ORhCWTBwwCEP86tx
amplyv4fRjqSIea5fKGObplygio+RoU8AFUC9MYW9DdK/xZCOLUQKVUKzku5EtAx
bS0VIlpEcTlL0S9JtEeaxeTY6E938kdpuewyOWNmRMR0R+R92A1hVcdJEjfujwi0
3Q8/EYKRvfDLnp/p+zBrq8d0AoFArdnhNE6FYWb9vSHg7lZNp7+l3PMnXCbtwPd6
C55PYXx/mX/z6EDLvNRSK0TkXYw9ksCAWPQZ0fYm0loRSJGWjtGcyNeIQbKJp2Ls
NzK+WixCnnVZxaO3Zw4TakTXPxrZiytmMOxLdg7molGfcATh6k9+iWRCFVbiJwkJ
Ks0WPBG8xgvWbCSTtN6bJyxAL5VYYaTHYCYZ8ROd3Oi6XjRaNYPGZSep8y4QdfIr
QaCmHWEcnOlMb9yANKQdsLF6Pvj/QA203WwhbWgK7kYHpu4m7mCxKjZe/ueTdfJB
l6n9SXoe7IOSZi/bafTBKHdv9WXCwOGpVhROI25dGHW1UeW1NGZzsG5rBu9+09Te
XjNkjYQbkhAYY0PGnhTqng+gz7hG6r6CBtheBqDDWP9m7eSwQid4B1IkFwhJmU9r
LLnrTAMLv6o9NNXKpVWElst2BOYXgS1lgxLTEAAonwnYBmOdZ4929hv+BBOF1QuD
0qG2t3YKZPtsIirMUT/S9cKBWKbmwmrOZTH6KTK3g0sjz9sh1ibGn9l5j4qaXw5v
T0k7XEXPyOg9isL9Rk2X+2f4l0hjWtJxEglRlINFabvINpGYY8T5Tc0hjfUZxdAo
X3h2cTE8s9vTfyQdrmRCoX5YKb0yA3aAPXN/Fz1JMIKibTav2YsyIsZYT2kUNLfD
fd47HxjGToXI8xtTzyW4Sa+IJ4JZgZzDzsN+khQYN1hncMn8amAukFwAT1PTeVG5
8yQ5vi0StlsewBb8F2Pxaj2gd4uHReWEvyaLfjw2pmolU/fKQ8zFpxTKSSb+6wOW
L8VH3KwqXQFE6sdf6hdpTRd0t5W+Bn7ld6obrlFf/CUlQ5FmUcedZw09XTq2kkqP
xTXQqsrH4NYzXVHb1vua4Ujs2HEsCIesWtCv9khNH7qQCbqNckq6M2zHkDyjww2L
tMh4q+jKZF/Ud5sQUJRE0Y9NUsbPpCEGCrfmn3qblECn1ABigsgTokIojpkXG/pY
UA8d68jbhHTrOei395etWgl66KFt4JIORd6gXkiieH+72O3Y7dFYwfRJVkeJHaLR
TYtS/C21YxPkgqTFVsIGlUysK97fIcsDci4I7DH2wqwOyhmdwEqSJr54uJLQtHZo
sikGRvEXan/xATF2xcnez6Ls7w09dYS6U82Zud5qZMFsVNq1fNgmwNNKT/uk87V3
Ds9HIePK6ZydxH9JtPmJWnjxgt8DwkNl3+vKBcM/zm4LjSk3l7YRwvf7gVbKlqyu
CPhLMJNqpycvBH13iCWLwkPYWou7dJcf8nboQApwD8SvRQN+YFiU0NJv3RfHfAVY
G1lo+/VP9ElCnftUzY8E+5bOnyfy1sV3y+ytBaN+ntvKtXbY8BOoDvKEttyOAETq
XsdzFUVIl0ojYUtb/zzHH2dU67auuS7CwizcI3GjsvUkma9clT9J2/mE8MDZNiK5
oSig2ELTXPlSNPuuAgYI9ysj5eY/bf9jXlzPfiH3DHJSvbwOIzaBgyULf/fxfOZD
VITemL/QpcnoVIjBDGs5Ag6mF4WyEwnf1Vs77CqqTPwJkenHTjNaTUTBPavvAZIx
jbgl0Ngb3TlN+talPZlCHDma7l0FuDQ4GVyYxyvamOTUtWX4Ahyrvp7pg3e9MNvY
y53fb5DJZi1eVqeAoi7lcy74tYgN/acG+VeGCckp9GSEbHJ+U2XBIYTO56QinMdZ
qMTmE9IHWtvy7egn3/pZzq4b+7HBtgMMBcRD4wINd/HmT3BK/BkTO2JPvOwS1ves
Dl/eHnvuTZ/cw6t7CtxANZIA1iWuj5NvVIgYNsxbDlaEqiIJ4TImmMop3431VGkd
ngKUlOzQIoCg6NZihSOv8WjCENSkFUR66TqPSS+BZp5CBC7JgNuohyBEXh6hxxj8
ivd2xiApqVz9Bo8EKn/Q3C+EK7A0kKhuqbid2t3WAtU9CS62SRbChdTSilYWnIXi
j8L8JEWBz8tCD4c52coC6lYvwGPVvEqjaChnEQ0noSdYfyl+usD5FGBDnRNXrLJG
RtzYkVosAdlyMqv4LiaFJmGIjzMzbscEFps4bQqeVHNyWpSKhrp7WjVeOBv/jIRj
Ezj9VbSCYGKqLolE6lgcD+tI7kIgLNYOMIJrAPVFLlk1Zpej+yXiKckBHV7qGgJ4
E0OTNlEJoW4tqEXqMiKZIVBmnn9OoZ8zjH3IXRiOs1IX393TdfanfibEX8lbG7i8
9KmluIBlsXg6yxNdYEbcObMDw+CB1uBWgXHk04HZ5eGFmVMb5laPVZgv/QWsqpTu
raX4si2lBYbr7p2UbOFC6EnWetCWhY3QFFCbmoKep2+qn5OGryeU9hRcvGWeH55o
BSn2lceND8ewByUb7fFT6BfsYRe/nqgboteOs+tr3DfsAzn2t1OJ/2KOsAkWw0Wv
uimR2jKJNwUbfCGt+acop3Se8fz7AQylhIxnmnoivUgLFIIbWShiHrQ/RqAFovCy
MMYkpkmn4QHDywfONJMH+Bv6zVEWQj7enYuMOuHLaMKjK9wsrdrB9banshdQeRLS
NlyC5C3gszwhz+VSn3HHidAO4oOxNfghAQP/+nTC3reOuWem3qrtZXwN/1Gn9l5X
d2Xg1QUhB1X1q9viV9PTaYMPVrGydb/3rjEMeD5Xu8usxuBAFNE+UM22dvbs9BPm
G0+Y5HZ+cAT5Yq3LXar+ok0SiVecrsv+/Z8tDXrJ2Z1JeE4pCIhpobO5YEWC8d44
5UMIXEB/tQRjVxAGLxMlg4lQdsa8IAMVjwp7/rYAoH4gHlUo+1ZZrw7pGPP/BRT5
7w168Vs1ysecjVaS4ErelGARTtGQIRx4sLADIoxkd/b8hJXPgKEpn6+sVyvoaLEn
UlrBSgyIO8npN6Kmg+7tW8rDnwcQE0PuLFaLcAZnYajYLInA2cbDtscBO99cVh1I
O9I4JsfBjGDOSwbW2RA09+3lAzfmhyFxCoaf5CBWMBDpgw2A+jn4vcpvOavhAKBl
rfx1m5dfU8h9dgmWULFV9g1eddcg+GUsq+TXroSVe4YaWhGSa5sbpvAfvEzJkPlV
e+nWYcXUrmBKVctiw8pDkRzktMZMAD6HGzZSj4LauycafcrBvqIxhymTFiESHwFx
bkjWS4Hf2iLSiOaAsKVGdPR/CpMsdZPtmMNOJY9QUDeaNOKRHOhbdeYfghhXe5JO
mkTQfbAe+KZVtmhD7mebraKozCBoNby4CriY0KiIHc1ox+4x/f2tjYa+hO4N6Gzu
SSFgbiouOAplEP4bJ/Hz3leikYFDUm5+nLNC+9UWuhG5HPQuFwsNMqfeh50i8zOH
FxtNKKHPDs5xrxw3vGsUgX1FCHALaKGvwK4SseUQAfWlBk8jJ6GkTA+RhUL3SgBH
gdl/jDE5MlpiO0WQ09TgF51Hi7mBQ/OMEIRXp6krcJoep/3BqKwaPaUTI9M6kNgZ
qqPY3DRoOGtfZrZ1swlJ5OcxPhOqnAA1ZC03Qutedz08hmDxuUmkxrMJyrgMpu3F
Q4/P8N2HS/LcBm5+3oZurclvh91t8ZwtlJ34WlmFXeeD2/FZlVvHX+1OGfGNIoEt
bqhhs/x+D1QhpuFVt1RyPu67AvCOcK2nbyBIZxfFoLDW6J9mqI9Aasi1OUr+P5oO
ZQ99isiCIhhZTbqwK8fJZYws0cBTJ1/ODKJUkrHhbwfZQPTMapAd9Xu46HxdTDFk
7Hu+ehxXHCJmI+c9JoDAcPwFVxEO+JI7cwSTTU9DIVozrcSFet7EzkbgQLJk2CmB
ZQw5ILQnKC+iNEWUTT/hmMtIa40s+rauOB++WMsvSLrEoLQQ9JqJxQwWI35imNB2
aH9Yzdhu8bE5uodqtEGAfZYWIQKPKqP4OSufg0DqwT1Hm1bxIWkAzOaf7kkCIDxi
UX8ZVqYu/gSiQBGeS+VxOZB3RlpKm0oi71/TQ5L8zoNAnDW91tOQZ2Pwf6GL8gmF
BGytTC4fQ+9KPmGk2GvJS/CZ6yx4ui0okWc9GRPXE3kXNFkZ8b2y2gRQyqZhnK3o
NeNjj1TlyZTtcyyJf1jR6yWGaO+tVFLCUjqvRbRQBgjg+at3L1xbyCrunO0ru/Mk
XZFJxAlShkL4krG262XqDd5b8+hln4qUdcMlsSIVplVpsOcmYHGCn34Fe+7pKBxy
Z6jNLP+/R6u3/UMvTcEvcvH5Iuy1Hz8zUSW+8kLmSdFiMMjPqkxCMKgC3Q1ItbRD
wiLPnZRnlgJocvMXFgVHDQK37fewxJd4Lu44EqPxobb0EILc1Wc9b87zu1bcottk
jEdQOtTgZvmEZAgq+s/CDhzdaAnsvVrwympJ0bxTOli8Lid5rm3J5QQpg30hdtIZ
qnrib6KTunXuLelyIYUCxYZ4+6OmK8e9UBwmvYbWfAIFlyxCdabZK2+apq2MRvVO
seMWKlE3I5dfctg+oBEE53FA0FFDwsU48ChLIZHN8DDyZdQESKD94IaqF28m1PyX
L+Mow9qDsz2eoy+iQ/3U6aqjSkew2AIkHzpm8kJJhaToD9W0YGzmzeYkXp0mMiao
BX5XcPAMzoQIi7d2JESoViKmooYo4xAesACdTd4DIg0iTrTvBqLxdOS6dDdrEPY9
zL9NSV67dNYz+LMFaQUzOgrY0ePO0zS6SvVXXxM1RuKnsj+51plbLJIKeQzCCgHi
/OS3/IEY4nI3TH238EvG2W3EZH/hi0zT5QM/eoxYlQR+YSxWom52Vg2ugwerASEz
QIYyKPtc+HHjug5leFte2zp7jZ7ES53DE+m3dCBFKNethGfa+aLSThh/P6PJmbk+
jTA0b4PqrfTzLkcBv/AIW6yQVmH3pdI0ntu4Wwvfdt55Vpu8wmh2F3VyAK2Xov3U
aVGd4jv19D5t+J0MkdqdKvawbvf101wS7SVcJmKiokl3qAVfF+7YkfY/C45Wi1oF
sgadaNX8jwEaiveMxSyJ3ZDIzgxFlApDdAv1luAWrCpDXkEdT6nNUTlinBBDfnI9
j9bbN+wvXQjw7EitnrhS3JzovuZTRy+SfqWgKiQFDfd/wgN6pxltZReld4lHGrQD
P6O+PNMhhgNhsqCORDXaieLcT+TVunGeh+8t+I1sRSYi7rJ4UHhElcjJFtdUeLhP
ojCitXaG5WLwwrvxhfjgTZDLuKQqDxj1Ojjj2srT4FTLZsRsUN45CRGdjHlZRR++
HxMX271FapC/nuaPN/dlLmIbE1wDo+WPMxtHnfzmve8GQXCiBqssCIZYUshJZhmH
iHNec6wCSd4VqTo5Dj1DjnWqRLbA2Z16Fxv96YUATAKOWTVzPQsCrfWDmlregpQw
uxpVUTc/xuLIeiZrZJXquAOROYZbPqcrUcbwwGc3otKl2jazOTMbVPDp1h4QFzXa
ZLykTuqo+Gks/cZ4afj1B3gLl2N4Tp/fZFXEHQpqP7MjqhnCuVSJJLljNeQ28gqe
M/5lmzlif2iAboGvMJ0fM+rVu5QA3pdDsDiawhJfjs7oz/4B11md8aX0XE/1SIaS
vTagCIY95Lot0IHkjoF4Qw5cNmHNZmOJN7P4I2GvWj3qfbAsN+P+RCObgNcWYQC1
hLLMU9lQg1Bdye/R5vKkoAv6dGP+7Ebrscj/xzDK2Bxt3GzpnldM14VGoSPEYoKe
uPIJnQqXHLVpA/1jKxKUCi/bVp4bXr2naSkjU6z5Iu8hrrInug4t+QGI0hL3BY9f
6RwOx4vY+p2nQQOG8NaBjausOoW3+Ia1C7xsaL3Hks/4RLgjZ8cYfGzTT7BrLFrw
2sRrHgsSuI57L5G6eF2apmkOYDzNsd904sFHuIkS4ck9lABP3axCWZtQvncqyeXo
56Y5f1v5U5R8xQHOR1jaNNO1hKncUbIibHGZudYc1B1s1NMbEGFEAy160dbw97Te
lmxk5M4HFc64qg+0PU2YpF4sbxPpdXs3dtVF04tp/Ee6IOAhCDvL0hJP/QpMBBqf
zS7gXAg6FDlPcmTXs1uIr+/S2YhpGD6vqvrCaDBjmDHB5N3OMdSrG+h7/JI5/hgv
nz8xrcvWQvh5Xaxl84DUwvWP5ODy3lMXh5c+B6xgQEUMpMT5SLQ10VyB9NMLsKkb
6PDEbgEvFQ2Aues7Otxd4SjAX+VtoqEesmRJpYQqu4QksRnRZXe4fZeslsaKkU5u
p3knGU4WcrZnTaH04cWWA6jg+2c3ihKxLjTPPAsfF20NJPShvApCSbmH24OIqgGA
JfVVgO5z4N79nlQ+PqImO+jytZXgYLMZ05mgpgA5Y/Mcsl7BAyhikQ66fkssT8D9
nBJiFNEA7+ibwhS4jrdUy4+zyQ/svFqL9TBosQH3CSMAMCP0asSsmEwoX2TliUaz
P6lWk1PeUQvIsNpC8Pq5ERpmWtyP8Y8qeCP1qQlm9wY/6h5P7WoePjL4zAbmLbeq
o4+cWSiVce7jhNwqdNcW5iEsCw131cMU50DqqR6ct/XmVIAv4Im3z6yEnGlIPmPf
asSvbDohlJP32EfhnKIj4HySOjXRoFPuH5siFMA3ohomBVx2AbFi1wU9+naWNyMB
sVgn4zz4vGvAhVv/Ofz1zWRNSOxQbHiZloDj1PPOvihyPqgpMl4FTFDPtH34QdLo
o5yU6RJgZAUVSuUnCekusGL07jCCp/Jb6PQHTrN0xJFnXQPmEl35CEtxr3khUJAz
mCI9WK0mO5vH0UXD+RcpUcgFXiMDG4AUUgmD89Ra3Fzf1WIKinvvS8NIIf/xIPST
zKV50SPEuIJpEIFxJTOXLoOOUfIUs74Oc+gFadoIeHQp5UCgLP2IbWxQkMBjChYb
9hI+tJEWcwmybNwqIal/RPiq2s25p5cqcPA/1np43QvOpahQ3BZAMtGJlICTU5/J
zGAyT+3rOqkdSEd9HP8rGPBTWPZ/qb9Qf3bFCtWZBaDu0JafpK0/kJjQETMaC9n+
j2DzUxi3Qzbt0jzFFbEQGGuQu6vN6tCyFfl1gB1NmneP0GPKjkV0n/I5mL0/oqUu
wCk3c++phvrF5XX4JyxUblE2lO1zOhs3Gn5cXhv8xRV+NKHg5gHwKFwWQtEowc1i
Y5NOgh416CtbXT04CH1lkYMzsSMRcaT9Uz4OZeVjGv7/+8fCGzJryRPL6QvxHzF8
CvmLD2g/5mNZp3sao32wimzdGiWHEQM7q5FbJ9bT92gs/mDQHYMK8IklOfsCM3/A
91t3Pg7RTPCxEJ9cHJHdnGHHV6WB21tbtg7utcAKzfE2zowhvwPLNZy4qn7lT9DQ
/fZ/SSeHWIc/hK4nTy4eFWo7xSOwSb2wAcFcfnABsgrmVmC5X9oGKpPIn2OlcIL0
Nk4vLmXVwHElCsNfOXfED1qZHXpH28OSQD6OjbUewbV+7PbuXiatNPdpWBj3/9k/
A3sDd3xO8wICW3rmIruvVzxlyfc6sgkl0O4GeedckF42049JFCHy89lfzQt/gdOs
WTqUxnlmmmhyyk6zUt5K9bdi1eecaE2isPVnwVY2Z8Y6J2LYpPig7X1HprLFwikr
x5qUcTct/sc80hISz2aqPTCm+jAa1QA8swY84Ru1tQuMViXn3aHXjWRnLbzlOsN8
lJ6XxQffQM+tZXl6c5vEvI23F4q1MkBqYIf7CFZtPZg9uN1LrVpxtVIIiaiMw76T
CQi7jEHudFS2PYTOvwkZS0PRDB6aIOZeIxlriTMEIVY16bEQv6n99i0BTlKTLSzR
iulhMhNntbJ04SgB5nyo1ve+PgHhOSD1wjR2qidn8A4XkVbtU4nJq93zBfUEZL6v
OJ3aeF3RhTpyr9MyAqbOiCl+zrb4XFCzyVg4LtBjyHdkgkhY7yGbtb8paRZ96GL8
5f70886G6/DyfJ1bxpIKFCiVKL4eeU9NJNitKIm0w17PPTY5mtIAAZP+d3x7g5pu
syVk15oloCJ9Sjhf9664bZMa4sfMkl5qMRRkjxwbqQr+ifu3JWPoq7v1oBP+1kLP
DcvPezyps8ZVYYZ9jkrliTtIsnxGA08POAB+kZ0X7epb5onwodocZa/WLm8Cv7MJ
63aWOoshD5IXsPH3+qFRJ1KJ+eJ4iEglmVQu1GkOS6VPHD2FqBnKUo2iBXVtdCWY
+M5pJ28rsRvaIc2sz4qCnE+2CoweOmN5PC6RE9QqFTi4shkzhm03NI9yr3GOf8dB
TOYr8aaVAfwohmJ+fTMSs6weXfXY6UKrs5XYbtTNVTfOK8rK5bwAECqp7zBxHMQr
cv0CVUSPUknEkGYgmNlly+MkaGKLOBIxO5RdwW5XFpxL7J4/3GAFWB4WzqePvDD+
oMTN+9qSFWBN52/6Z/LA3DGEHwnSR0rysMwINK8PgP7jm7fY7z1CXDO1QbM49/bT
PcJiPCP0SBBI9ZuU2jFepsTXKx1vEB0J0c0WdvxFe7sUAcrnVI2IIJ6G8j6YWJXO
4Xuhtt7E9qz9jSXdme7n3Y+FGehMewBM5yohqp1ygRPpQ0p15satK6bTL2N3Fzgu
PpJ5mNnpSSwGZ2h90/YKNNFEpL+H0xzmf9ECXWTqRwxVpjlEFMpdISY19apJxFbX
xSVRdpa/IgMda9GM+lNBIi4s0icVSbOGmOYzCaaYnNx6oFRxpmBgvtJG/92nkoA0
ou/VHdLNkCc6H3iVyMhiLKICRXS+RtrPowBHimCI257dv3fnH5wnjUCivkK5Xjk9
wQsRICKwaLJ5rmTfDq/ajNwhP4bpi2BA35uumS1gSRKyh0pCKJW7yEbrCEbIJURr
hZlANYbOY5QVSuWe7Y0av6ZjX+QztdWWWvCgVu0DIll4IhBV9NQGGKLHBtyMozvd
kmQwKZuDUtakyBQ2hFZXpky8C51T+Iwj/vsx7anieEQ/BurZFsfqk3O4LXmEQUpj
9O25TJ+SyRSyzj3t5pW53JFrq9mzhXrjdj541zFR8DqNij4ezqvnDqm7bpKTqvD1
+PvDv0x1OA4ppEAr2/f2hfqUcvrInEX3+TyLUBhX4XFxA1vSKIJsI2eaQOMqJd2M
2BWYAan7/ijNjTP4Jx/agjVobg3Ah7nqKcUPdlf+b58v1jf+9IJa2o3y80Xyxl4i
V08Bck5oPsPv34oB05xPpuopcFmJCZEwSrqRremRDyCPG+35eQwoT86bczhO9h6A
xR3zqSAFWuZ8VqgK1RnXeDpnDqjHDwPV3nYcxoV9VwiJSBoxXQIp0CoP+SmWyqPJ
AKqqndGsWQePA8mfKr7e4GprqBsK31EbWQDSETt5vh1e7+83A058N6ZV08pYJCiS
xLGrOFl7HU3/BB0AScikZVRJGUrYZryQyCkMXkva+Evj5l8DcJBKKvBGXf2QVmyT
iI8ganqhlE9kXQ0de7+ZHsIkeKDl3I3bAQr5irgJDunu5XNn+cgNrQIMwqDTRw70
B7cexIu6OaocUymNLHZ+4YCbngW+qu00dwHhJjjygO/JDMxqCsDk4N62OGLhjJRY
8pKb+E7jwAmFVSB8d9D15fDChB9vu3fiaEJTelJzFtLe0RU67VMvjmxM9QI5D90p
+8y7P572670C84mtsjKqFKAjbdQc/d5GwZ5SWRuoWsJpq8TUDuTHwfpSZzX9ZUPh
oVh2pNuuhXJ2GzntiLYmmmY33HF3mIV+KSErtTGL4lJit7DbLOM5xkhR6vel6gXW
iBdWf76c8H+Bk1J29ya1XUZxtEVmy1HNklZ8CKEcDEMXHk0C5MnmYvPmK7RbfzMB
Hbn90r8+/y3w1bkVaumDl+zus8TQ9kXpDBe6K3P2K0uoDJhqSB048XBBRA/k5DNv
wymiBTLFeQqYZXsXwFZPLQk3YbV9HUOyJzpzGbmS3ETVhD6jCSVdLwtYAgcdNgWn
fq7jHdyK8RBFYz2zdQqKW7C0worGuyG3bvFAe4RExVsg94dL/cGmKNWwe40GbbPP
fLZcBVaQ8juzVRLydpDWL9+2cuiVtNbGYHHIkzFj+yHMEaOoN16M+bf1BTvnCjGb
LqxE7W4spgInYuim/XgUwnqzXGbPyTZbFYEeKJ2qs8kOAQkc8QmNxNMi2ZZ0lUda
VrwD0DeAav9SWRd6FYRgjTdRLLwbBbga/eRvMIujKWqcAPjj15g3VUMtgMJhkcTO
xp4PBDtofymEzU0f7cAm5WkDeyOu9hHX8VuhplIqWtQe+Ou8rp6H+MqBe//pXLEc
RQ/v597FAhUmJ3M3nDGrxIoOQkvVM/J5UcDFbRErIW8UitukWTDCn8sUxzLaqmgF
P3Ivxh7RlLFglRM20UpiSzUyVLNYnwm/PZCn0X/TfYo0/xUrUjE9NSyPIBXilAGy
ODuxPUxWS5C7XslZFbyCVcurBgjVF3KCDlioVHep38Cmw2kuN7MWTHCzhS6Qxovc
tnO3ZSAbGl7jbT9j5swbEnnBMqFgxAglZzolIfDn+NVC+1sI9l8bzeYGp4SdE+QW
x2HVhxYODRnaG2La5uXAyJwPIKEoPpO1pKIs6OPZvG2lwb6ntPLhCf6NOcGGnX+a
Wa3gYWWqYRbT3UCiJ7RxqDgxfNbYHZUS2b9C4rXCpZLYzYWDFbo85OILeDTJft2L
sAXrwjxUllJvySsZYAqx4OSehlvqZG3HpgI7WJgFARI/ARBM9D7eS3nHs4XZbmqL
tbXp6yIOF3BHedg/7Jl+//GtkKNei0++BNEPJMbO5H59si8oimNbUw/DoljIaGhb
Gy5jbyW/sq0FEAhy3dYOkulV2qTItwgDlexzJcu97YX8r8zhEMnMhzO7CaKf9voX
L4GIrCH7JMWhz0DPh96Bluy/RLphOnTyXibyf+tAJm/CG1lH4+2ofHJqXBhx9xoD
sEw5yKY3QtTk62bj5CfLm+D3thgSdGMKYWnrVAwVyZW7Tqeuoh0yIGAxhLbauhKl
x8hoXwAt+AT48lcpONLOau/QSwtVY5tlLqyMkFysrPcWM3V/xk98LEbztgiLKq0u
YDpmOGOcMCubZvEDKplXe21LFWxSz9eSuGZiiC2Fh+jTavjBX1SDQfMJci0JqiX4
9YAP0Xom+Qkurr29Wb4kKO26z9h70f4/G0yvBUTKKLjSM/3OCpuZEJ9e17xD0Nbf
nR18IoqUiYXdlGzQQjrLmV2W+b9WGh0oCCcIIRcjehj/ZydpJSMVvHkS2UD1J+p3
L7eMHDPSJSMKx7qVON5fQtxpzS5MwwzDNFr1DQ7dLawxTMWgw/MjeEAgCmvwS1IB
FebhXrWf7OLgxnWj9ChE4+pCgD9yz1i64gg2hfAUo7zbePUgmdtUCVJ002LMhClr
QxwRNlzWUvjDHezTXvrh2dUBu7GSpvXCIRWTOX3cjwluCFXved8yMzCzaZJGuG0D
bf89WjMKiFnHRhSS2do4F4Y4QmXDPgWg8PIulHmgARL3yf33F5PHdKl6hqAqc8Ng
j3fAV9LTEONt4Nz2KV0wbX+XcB/3BNy0yHYNEqXPJopwx+w+RJ+6SFt2VJjp8AkA
hsspe7Syr51t0t+yLDcQlxOE8S4/Ana7+e7OBmk8ChF6HjXu1Mfk4ToEYbS6nFxA
h2H/SAyzsGGK1L884Cx1ESxNWzqoA44PStI1GmDZkJFfRIF/7NnT5d26gryRRZ7b
hNSFN1xsDMaCAYfkyhdPi22YMRlfma7PWeeD9tDiitB4BZb+uIlnPT/rhOmKW34Q
2eQ84q7NE0GmFwXaGzxquLbnhsu9cSh69GnwvDY5LikSt5LTUMdUXcXuCzJGVQYi
4w4iasmgRAQfgDi3uPZOSXfdBhXQhjGD8se7Fvl0uig6ZBRad3lcqug9fK9FEd44
8+MwaZmLU4wF/+UMVoOIaoEUYOjbVzHCnK9ZTGrT43Y+H0V1+Q1Mly/oknwjareR
+mYGVxerMHx88z9sUy8oi9F7y5h1o4ozfD53Rl+KRkdnTSN2la5gF4XryGvnKvwK
UVQIvhG1v+OAlbI1WQEep3Le2Fjk409e8qmWx23RI1i6o8fSjZwqpftH3V3HDaDx
vo9Cqo0RyW9XdxdpQp67iyQA589pQmgFIOC5imf8cP5s3iWcAyyUzGKHpysXYrS0
LBAhHumPqWUcPHcq+d/vMVZzDmT9/g6MyRLORcNrPAwNrUYD77ETSO5di0v7CcIT
l8aeGcFZbFoZhwEvxTEkUNuu4JB91cJjHBJHSjo4V8G/Qw5vcw5ZshWTIvu1W2yS
45E9LSxMMbn6mc2Mc6qprhVkpzkNszwCfspYyCX5dx1izSL7IvLdGr3IbtSRXHwN
traWj+TmFR7jurgeNeLMlEG73VtfR6IrUjIkHOtwH2m7L8XAB55ubtceHg7I2S4w
nEtQxIcO94BKNVisg/aijuVijxmpIKHanJ8C865MFc68BXo9P97A87hnNgOYKp9E
myNjHjt2Z/uK+9zMBWmE3c69ZBJLPWSaPpQvY7R3cXnsNlWNTg96gpQPX84thvqw
alm4Ath+TzLrDQ3YrneQ37wR5ltXJM14l2QMyAvCjTGIXDtvz6hqsuoCHxKSZo2Z
yzTPJmc6W1XWlt1oKwwd89gjeZZEM347/wJPpbi+yRvHCUVZO6oRhclWibAHiZF1
cM/t4X+FRNU5sOeZC4a+pI/teMDJbaK/d69VTLa6EqupEnpNqxGPW3Huf2jSx3Ca
DIiMey0+WTmAczxHpMuDPvI4JLCL5nx9BDUAmokMJxLUJRZcYh/gWPtNWVO+Txpd
ilQOwowAJflVkJjf6fYzOyYY3bb4ScQCiYt89VlyzRisUKJ+hL7qdFI3wMSaDA5L
k1D1XDsgugrZ43pAY07kkfU5ZoJEDss0AyXRe1IOtKNTGI6AyHgOMh3ao/DjAh3s
jPJ0uvg3VkEYxY+60gTu0ZUEjPn47HbLq3+BLnI4AUSnhJqcJQo53iKGlHAx+hBy
/OKg4WOcLjzsQWYS6u49iZEW720nH4jhat3qcJPqqGjM6eqQnfItKEcDW/s73yHY
Ey31qChyNXn99Fwel86uJjnurNoI2NzkF+HT0PQt1/ZMj8+dS7TysttT7Ypsvjcb
q7R+x7vfUaB/WdCD8riJq8V43xMi2k4XRZeVlCgRcpRomebcQ8ZGw3jEI22/ppx6
yuIIy6JYrKMdSZhduGhFVLGiY2YwyE7rLFEBCubA8jM4Dey/wNuw9AZ6vlEOan8p
czF5cWZaCbgGtzbStJ7RqckwUQ5iFarbbOPtD6jGGKG7uZATXnILUxOSuPnKzF/B
hdsSMvPi7v4/iqp4ZQR4+2jeZZUlP2T3yNXLJ8JuFfciSwY7gxKVMcFXKlX88agK
aqvWMm9X16V4z/jAqHWgPcdxfQ38ZE+tRkFJ7E15xaHsGfL14O5XSLWREjrGbaGb
m8qnEbwJqQ9PvKoFkJGJ3KPyAcxJ9Z+1cwTPuI3K3Z9sVR5ULZAomjvT6CRgJ61F
OThqZeQaT1bzw6ttj8fhijnXXAio7G9jLLmkfPlQru/FI/pKRZ2FE5xB/xYgfJvz
tVM4ehPxmhPhA7OqCdtGCnAllZOeUSUdAK8BEI0wPaNd0p26HQNLM22C/F0SYk0F
qV1YvIKq2uM63yB1kj4fGn8duUj3OcJ4catkAwzOJ444GKPLrQuoRX41LHl9RmTB
Ma1+4IkbXHd2zMQ8SlK1hE8RtkgpckuQUi2CHo7ehKSnKExV4dOVTxQ/N6DTrHXS
4hSQff0Yu4Sz89xsnXmvZK/NBV7SC73gMhcfMrUG3xCDNXjD2464m/uKz4Uc+Gzl
N0CW8JHE8JjZwonIRDrLIvU61EceRWHZrlMGSY0SDPc7nLdvcFfm3p/oB4Fnbkdc
VeCLH6vBb7246VgTeNWOakhGzppXd/nunq6giII4RS0nk+OZNQ++h36qJMIIMN6b
XGslDGRUDOhCbzOrKlHxp702eryfvjnDk20gntnm2xiTFLikx7axn8BuKyvKY1xj
fpJKMP4t4MQmKE01IClpQJN5biy2DXxxeMJH72/C7CiZlqw/RvbCnjfBErbrqSln
rZ40e2scRZJuRceorPkLlhxLUIOM0EIqFfz/b4WXJJTphoIpf/k3R6Qixa1+8nXJ
jcNe0fQzl08dCrZxVgDOMO0tkIMx7dGP7ZV0nBt3X2YTii6XUDi8IGtW1l8w/VHV
l9BQsDOhvLYmXLlEpP8IG5BMZNhsGJjjgZ5sYutDZTnaZodpQkIwpjT6m5mtps2L
OFc/+N6Ditt2XCiJW/rObdUbYGGwqOwbGF1icTi1FJhAHlFVI9o9baJjRacnSkY0
LqEpd41lzLER6n/J3snZ+UyGK4X9YVZ3THHeqkjLXoT33qDe0OqcJxALP4aIWxit
KsFW/XTYGiBfZV53AFh0p3jA9e/HhcNioZFzk2JWbmTYMZ2KM0bZQQHhNTn/h2qF
E1LWALY1CXLhyWVIQZOAfmya1feW4++0KBNRB41YlALKQDL5eir6yS+5lG0MTvpI
QEVRJMrsmRBXIuO6IE2Bkepdnv0PDIWgKAdiAWL/+IcyUeW79+hD8/Rdz03RDubC
pHLyL3bohIs9QKLjVMSZM5CdKoWZtu4OB+6rw4y6MBNN3QbnucsTmrJBkKXW0wIg
XHB1n72N6pbhHKG01q5agrPjK5uQTdOezX8Pe1mxKktwzbD8NBZStk9qm27RCh0S
7B9jK4t0sjfCI8Z2rlsz3yL9S7QED8n2aEJrWmDPVWEMi7Wx+da2R1LIxcFyGr2/
0IKagvmAeLYIFYRhGw4Qmi4QADmkO8TDe7u+ANwiUZ/OlZtklTef/jU4YZvLL2i2
4MNupEMxa5zTMzjYmScI5rjfVc2M8uDZldPbkZDtWCP2tjZ0a3Oe5Fvx4xgU5Y9Z
hClR7LJg1H+vlt4GZyYwsrAsJrm74gQ5pxpxNA3/U2s=
`protect END_PROTECTED
