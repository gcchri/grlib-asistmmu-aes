`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvYET6DsRaUDrocAacLI11jdHsFWdzjC8ZRtbIxrZdpem2Xigl6nm0Ckfbi4luPa
C8nU+G+bTuv6BJSYvV4qaC+zIPuKeRBVimdJbaT8JSXmQoTlZQq293lpmSsriNzM
9qyj5UCC1UrttIbovWMPp8QNdNP9txOEkmb1LwJQFEHy3dBS16eZ3w/p9tDrcmtp
gUgPprR94QK1YmYK201Q4ry+u4RW8nK92AqVcun6/sX/qm1HS1k2TmvOM6Rk/9Ie
+1jXCzvLB1+jVL/b4yDTvJpHqPSSJcTgu4Wh00QSLBDlDxXs3kVBgTzAMlSl12+b
jtKuunOYaPna6c+ExFh0Ww==
`protect END_PROTECTED
