`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dfD3ehgTaq1stNNfWSLwpPrGXThRr4BiqV4mwFJSqceK8U0OnMTFiHfgo+8hK1Nk
s7FHpgtsVChN50St72MVf3dx+D9t0uwsGVzcVsT8ZYfaR/3TWVEnZbiaxpHMJ0Y6
mDbvtp5T26ZwOH6RPcuFB94r3IxdGa5okgjWQY5CJhB1qbTPUHJV2MOmDYY9RvME
0RAFpjdgHQFBAC3bC0meDzanhVTskKArf8UOkyGIC7akmSVB/Hw7gcMjNTumvlIV
CCgcvFV3mnyQDKJ1wFGnsiAM5IcO1Zt3IDuQDSnuuUHz9rDrb4DzZzmgGDnY2KLy
VR8LmEZPgTWHLKUdl6dqVu2vWujIAWnvt+7Rnoyb5DAswTR6U8Pnl+qLVguzURH6
mKRuB9B18yXXdoGR5ID5BQcQ+Q7OKR7JsL3furE0R7T8v0ga45iZb1AVsjYJU9ei
HnU64A9uJb2O4wFE5frwVjEhrIf8n+zqvaHzt9jyCSWg8bBg8A+eBjMErzah0Fvz
RV38mKyZoS01FBeQ7dKQuu3bwdCEttq/cxWOy3kGomwITgcDtyELiCr/LMTwvVYE
ERTdHLszKX7FrHI+GRIdL+vn5bRIy3SrCwdrVqGYzRf3yBSB7kaFt54BRaOLzEMb
AOAHg2P40cT6TWBFySqyi5dnM9QEKCmkvKWYSggMgvnFe6cSHt9D84ePu5HjRCTV
`protect END_PROTECTED
