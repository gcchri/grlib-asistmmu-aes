`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWAHhJ9hYhipK6K5CeE8d/kQvDFoyGWQjRemQmX2ldFhAXl4gQ08sQSukNwkvDdj
KMsUbCFJNDe1itd8oPu+PzMyEDq4+dVXs6QZu9jd6I1xd3O/lfSLVtdcV6ufcu01
AHs0zTCfrbdg0to3Ku3yY752HATkjs1puREam224+U2B1BKI8c7qfkQ2J7By26Q/
ZNwMrqKNx7b5MtIsujsu/CQLK259uEHJdftqxsdgVWhQHkJKa/c6U+Notfs3uvs6
TQ3zdksuUjWC1ddFG+Lf5YlDGFVTFzzNxpADRBjm6Mm8/usDu/xhiEK96JNupKoZ
`protect END_PROTECTED
