`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jytLajjsnTliGh+7Dpqw4fAZUO56Uk6QvhCNWaYnvag9eRKNMyFEWfL/hEpL3j2t
nxwQ/OALZMJEQyzBUb0/pgjlj2MYSrHFIKiF6rRDXJKd8YpuZjjuwK9lI8trv62y
eIOnvNIZuOaoETEi3rvKAMXgOteuwFwJVj73dROX7LD/GGL22xrCB9MWCcHomESA
GOalIyvoX51F/9Bt/F5Y/l7SMPdN39TF0bipp18ULas5mDOXB5UGqfjqiWWzO0PV
mTvUQsX+bnZgkBHSQRxwpDMyD/PmL1H162UpsSi6hHTO7T1bpkPafDVUm8f/28tB
YqVGQc5J3LdQXFmsxDRyp40o1cxQ3taSljWYqpWeGXFvpbpAbI1aGuI627CuqXLl
VPG+PHHK+f6bSTY5JaREb4831G33IytPqJy4zwPgEPFQ4zgOPki7QaAWgImPQNbE
lXE5AQyfOSa3h8ys+lSkU8cscyUjY1rtrHv6mPkW8n9KxTa+hIV2+kfOudOGPjA4
7xvT2oRdEtCCzoAlTOipnqFm1Ed1hLrX4sj+WktcSFP4cMtJ4JSwTtyMO71lxWvb
RMpzlInQU5Lwq3J6B8ftmZzLximkY9iyOmoKC1sg2O06ymHzNsQsgRBWcyVw8wGI
9Z3nrN97CV3JsE8uskoWlI8vtWWYPF/ncP80pY7Sr5Vr9XSgDADdgN/+bYxIdVaT
FthW2tDp0ibUnopvFCDXIE/V0e39yAtXx4VD+KBLLxfK8AkmnSmr4Oyy31dY1Ms1
DhbRrvESUmgy6jQE9dXicg==
`protect END_PROTECTED
