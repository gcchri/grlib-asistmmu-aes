`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFHkY+Fl/gFVJ7hoWsUhLd56hP0hcBnm4oBRDypM1LVEZ4hdhYrIHwSjun8tlE9s
EZTtX9RKZNVjY/v6gwW7hGDHTemYbyi7X2m7baLh0GsqSeongR9Q/nagfjnGKLiQ
Dl7zMfms6jCGiLH4xbU4KurjWm5xXc+msoIdD3TPdBAqGGY0u/PpTpX8L+q/a6S6
iuNWxjb6ZmJU2fiRSlN2xnAYPMab4IkJlMfhbvQqb9JBEICezP2If0YKQ+7OKPeX
bhO1cWNW+Y3TntEIrXsU5vTXxjbIXW8omWNCLi5JMUZaCgCS+/1yGut4xEiE6pTH
WIpe6TQFUzzV4pYBGCz5VqIEYOmsloDz52NJbkOSDiFBbSg3haKFEHvi0gW+/aPw
37ZMlT0GnPrD+rIx131Ykvw2EnEH1rmGDjXJsxUI4OMGy8Vk8x1BVOCEVgQBAcpW
bH5XSwdi1cQC27xK+14Zx9m3nL6Kv7INTokmaBnw3o+kmK1s4Y2Du93a36f5lrbJ
`protect END_PROTECTED
