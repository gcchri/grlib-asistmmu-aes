`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NnRNpoThT9iUgcH/yNn8WBjrGfnA0YLKfqdexrIRkp32mJcAZv1tkkpMzAuwskR
o7jNv88LxAPPOo8jVULpqtGqwqnxHsZUn2kTc42HjpT8lyq3OVip0QS5lnoqZHXj
ynw13BYdZmQydukGgAzulUz9/Pv8IYfuyrSCVi6rYQ+v9c1l03fHX9U89Rwh5zJP
sj5OhRBNq0SXL3Q16pL0dYMtHL/SckVfxh4k113Im7NSyzlAzP6gqHbg2dBNCDWS
UdPoOz0Cypp3QcC0atu/bj+jDnbg/h/oqlLJ7NiCzWOS9a2p+9+VOc7XcWREXb3N
1HRDICuVjfVZQpbmCHQghwVbp6/HYQ5icQVHt0Efht4TalEb22EDxewAdTMseBf8
rggOjjfJXnNrAScp6Ok9xeMoOdV1VOPMcSMXf9l+/9Yyrpk1JLICeKbNn+3cxas5
t1IbPXjEnUwV7yGU+cC/aJ6JYX4AAfZ/gQ6Ww3bsI0IRGqIJrxJtyNF0CUWU+Am5
SsLyihNInjX40wo0iiPdOz/vrD7MBh6mTIwQpQvRfi67j6dxuEp2Sx55QyZ5vtVx
kaC+F+wqlFC5wtr25iYxiSIYdiWqxa2GkL4jzrN4FVAhttM28XCnxAt0APwkqvyM
Xy+x3MQ0JysxERqVoNg4DA==
`protect END_PROTECTED
