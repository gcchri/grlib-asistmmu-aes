`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBMH31dr/zX/3YHQMpSiSIuaHpu/UP8Uh2UIxSCfxPbUupsxg3YRQbaNMJ0BGCPR
D7mRl+/N9V91WD4vpSDpZhRc92mzPA9JgX55qMdLN5oN5q/1XRU70rNUX1ziek/D
vXHRRT+mkbg4hmaqaNwFUJt2rdKKQxxsOI6Sri0qx/xXX+KywWlHW69rlvVhjxar
wgySzXFNgCK0O3LD4mI0ITke4LvL+pmIYaRCbtFx4UkH1gYwx/QOIsLHqZ13XCy+
91nbevn93nQ+nrSk4aKluyzGHhPgUb/UfDOFpmQ9DulDKW1L2ZnAKrbolp95aeoI
WK7QqhndwIMgxuUakhlEVj2RYm1MjJBC9Tl8TgemRM/xeKhV9gaGkXT1+OLoK8sb
pQnHrFLsOymobpZG6Y9i0qv2H39oxe2Br8l2dAjubQaoiC4JaNyCDM9RnCBpIb8e
l3qFcekmhhooLuKgpS1t0a+rm661uIy756tH/Cu4V9M=
`protect END_PROTECTED
