`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VRP9oSrxZLHrSYU+H3HvVYrP2OIbNP0fn/RLd0D6q8r7f7fVr3lqYnYUQKNHRhAn
aTwxo8hSpw/qHem+qsL+xcxuX/W+FdW+imJl749fYDdqlYyCKk/kz8Eagce1zIgy
WOGqzUDEz1lXD4/9e7iVz9kkrInF5NEpoai5SwJRBD61DOJlVOevWs7HuGaGCPgz
I6ii+lkh2Mgi06Qi2ot/kL/7wV18dQrz1dMY+b59ZIpUOy04E7R6KJEpRnWmiQWq
rzLbR2VRvZiREBl2mK4kXWvFlU3aE6ZHGArvakXQdJyhVyI66+D7WxtEipiKR6B2
+tJL5Fmz0K0PyKOknNotjXMOU5AZ09/aq468xyj/N4WjH2WvLHRhr60OrhgvvTh7
gtpYdEiULZozhPmqDTykPoMegmShuqY9SpUDCVlKZ5mRk0pQG4zGY49YdEFkQ7GR
M2ZJr25zhrxJuEHk/86wzDluO2XHdUTPR6T7fFUHZBLXxnKn1y+3dzr5Fd3PM43h
yOjjNybE+wqjBnx6IO9VQ/+D+XSNlXNfBe+o5K91dmD3CQiYnUENnuoD7NcXR1aH
1jMMV6jaAZiztMHvS5GD7aE+WxP1VeiR2K1dl8qeCTRg7wNXuMv9ORvUiPIwKs8W
I8ndrXXukoKlvWbQx9fnfqnSygYV5pTsp9HDomJXOUPVhS39ZFUXIPwZNeyyeW07
DhQ4hnoV7xlxGxf/Yc5QeB+IYhEf8skN7reM6C4Rx0AmcFDOHbZBLkToPyptLUz7
kg2y30HCUuZEk7HYjR+FuzwSokLwXnGc7rJvwrosVx4YsAtG64fLpbAlw/CTHAaR
awjl3XFjhAICGvsZ3vJKw718aJ5ZXT21ChbgyJ+3GeqvAzaE715EMtfnisaDPZzf
RTMr/K56jzDU4LphVP81xr6ahhRHCOuFF5TZQ4Hy6uWBPfHqEMF8CWuOoMW3nwVv
CdEtdZyRd+Ism3u12JWZEirToW+SoJ48TvW9sHVvKLOlcAKgBZp9TCH1fuGXVWX7
xBLIWX2QRee8nskkvihrzsexGGlAcjUb6h9Pyd8HDOVMgcgijUgWdyLDqkqLqTHl
mWy1SsVvRFq3csUBmjzdvecIPGHGHbmDa7g0Y6riNxhTwMyeZOIovvWtNc/wkAom
ruR1KRBqEf8Yb/vm0xQ8AprdDI8i0pW9aLmsNVdflEqUbcDjqlPXYIpvVxGsJzb0
NP4VDCVg4bUiI5/uiXKHi2nZ+zjbVwWPdszeXgH0A3Z08ty+RFNlIB9xfz4ROVLc
2STvJn/pvjjbxxco3Y6jWIdPrX7tRtblEIyw+eBOoHBXyF4lAji8Lre7lI5wUZAw
eWAH0B9PFPRH+/Xlg9yd2EO1SWQew48bZa3yMDhyxgiiVJUwFlr8NDmNi/zbjuX8
KHqY/i77tMOWiO7Lpm4wu1hcjx/A7kk5Z2Bmwcb1Yg3tAWGdR1C/7hUo65JJoE8Q
gPml2TXJ1ANSE1MPVKX8EuG7Q0UOhRW28r2Ym14nzOLx+ziRAs1xN9jQhjQcObA+
iVkgac8oJ/vH+HdkVZF5cradPytYdviiBr/S/t231ZB7/3njAg0wGQ9sEx1YlsiG
CjbBXqA4V0obkmfeJlWG4MCkidx7KxIwpe1zOg4a3tmrMYcvkQ7OHC/xnHPB2qqn
NfJU4+WGqEVj5D10NYtpc+CCV1JohfmUDIO6ituRSoSzK4o8U0W+abDpoC5QZuO7
zQkKKyK9WQgFzQHplGT1xF9d/gIoDPFh1/ZHbAcOCDwLlzsS69EX40WCAEKhJySj
bQlHvDQxZY6fsBm6MzzOvE2wsKyC++J1dovIixNba83aWLhHjnKmj2ru31EGM2wt
CQLiYszJ6whpwJwOIybQ+y6tdhWzzu7orb96+dy8J2nEtIVgjrLc5oegLr4FU7TP
Hrv6AT33NFcoFohiEa1dr1JgHdTzw1WqYLzWbKGd/rvZqYGXu8QCzh76BOY1zXl1
de0Ui7tSFIpRhbCTAsmUAMkbBZswibQjlorBPfpfvzJ8XRTeRqXdGj3wg2uyIJtr
YT2vxSPAv+LhmPOF/Z8j7/KgGtL+BWui8e+rT+6YAa+N+fpDMy5ODaU+CBYzKt2C
2p1tf/GKYqb5HqAuza5Z7Gqw0DkDHmTpmkbvuuygEmFgWZSn8bBD6vdVuslPzDM3
OsI4rnS25Iu7drvWc9+Dg3eAKS5UHkxZOA74yKHPXeQ1bNVDD3ZXOZwooOJjj8jr
nQkDftu1M8984naLwLoJOG77qEkYEvYK/VmnlLp7XgIlU57rAQTdUeAjtRuglKKI
dLcHriFauyaM07gJSOXZ+EnDP5JHGUkd0qYdmgSqA86y+OSOuU1JieDb9z9OYPMl
YTMtNmcpgIEuOgXxvGg5+grKwEJ4t5ABv8Yr3f1CJlJDovIZloYdqcFiHBB8Cw1/
OAZIaUHDyBs5dJjh/oG0fXU4YAy8tLgQkSAIQi7XPvzpErSyqktZJ1VoEFYEjbSp
9jpF57v3CguaUtN5KCbFUueHyrAonnOjJwtgzW2d8wjyF37DwBsnC2S+3AlJk72u
3CckyBgZAbdLPlbIPzNjoN/OSUDO9aQc/zkGJYsWINY0vSOGZMvGyJM/4q7oonXC
OItfwm0HF8A8NW7CyWRDtBNVI+s8YJaq5jPyvJ5fjUkJMEZsoheT+s4Dn52GCcEl
8+0sWGW6v2djNTuQ8rrtwXUml1OyEoxIcqNZdtBJvtdkptdy4zzrXHUmt4a/vVsQ
80nNLnkNFTJeF3QVzQwrnfMOT4oOLfqRyK1DTRyVXqM74KhCNnAN2dglLYpHT02J
hDZ5MRFkMwA2Q3FJlY8S/A==
`protect END_PROTECTED
