`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mf/pRb+wRqo4PAUCZHFueGgr+DQt9rVGkCn9ozN2npo7wc433XTs+ekcRUbEgBhd
4GbY/VihCgugszC6UbGolD0CebmIc0wpoXqDAYKRGwS012Y73gQ/LAyjHCWPm/VC
9/srftXko3V76QcQ/aOXesIsS8CY74V3ugF+vTF7Up2s9gmxBTXBnAmWTdwtL+by
bu5diiNxTvQlh6iG6cS0O1g6ObKf/zvU8xwhCCtL4yy/FDtR45yZY7WuWMkU3mrl
740i/e95JrolRSObsn+cG4WGYdoO8dut05tmjxhOdv8=
`protect END_PROTECTED
