`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rc2xelJSN4OuhbiFoadzWuWuL+GE/J2RfgHwHxb/8iOFEmFndwXCeFjDK/CLGxXZ
+xoiyxAu+yz8puMZOrqfZTEfN64zy2qRfTnpCFVjMPDJXNS2yQwXKOZbItYW2Hxi
I4XEx3QN4nBpNIwdwTyAM91xC36mbuztZM7SPB1Qm0jlG3AMvyny+kOPMdsGph6s
ldeLZQqj2WMekZ404gKTgz7GZjsm12FuqRnXCgoiPGntnm1uECZPJxpzGIN3nnpK
XAC/TwIhl/iAQdmvxq7/G4+zKrRve66xXxX3w4WkD0D51QITMgAVudMftUjq2a49
ZXlODm9Ok+CtUqBIvNDOGw==
`protect END_PROTECTED
