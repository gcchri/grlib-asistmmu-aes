`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tjbXrfN3UUG9nqbvSrwzG+m+BRnMIL9gSmxUOS16H8PT9sjkTcTKF7JScaZp+VWk
1zQILxuV3J8QRXbbK6Wr19IQn6JgWFRRtjmfojnTy8sMRoGxtX90oNyugudoIAhm
CJ626xyWKyh9QGJaz2ZRKiLBHPEU3SMY/J4qn2GSGd3C+u+diFUZFOPcGg0cJ24O
0XeFkhw73jgiHpagBcOMsAyzPrBMPLA2oKLKMRmLu87RCRd/QoeUJ7QT/aDcAajP
OykOoXCIXob2p6Ovjc9t5yjjJ2PYL1POsN4UPCsPTLZz+/KEy6CNdrJj6GEAuIez
j/MtNlSGVWLvyojrG5KCTcqbaD4JrlyH9zpE2pwNSP502TdTj5CcHL9Ly2dMYKxy
2BvlyucNJn7QrNralobRrs1Fv3Emlh/GwKjmZ82ng7FTgsuKSJy1McvlQzsS8YwT
vMfdNiG6wJRuWAubesIE1iiKW3cbosxUvrOguD57YSez/wbJ252fkh3bak//ejFX
8MrfFpB2jCKIcg5lydKq52/oBFCyaqKe61gPWYakMtl1BkaLmn1ay2DGyTFPbOGe
60M+QFqjkjBc6QKFxWHqpA==
`protect END_PROTECTED
