`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrLroPZl1vCPGoJZp8Aa7IVDhLwsIjDgcDLYsB18wrJ1HTMuMp1GiYCJejKo+TRR
yw2Yhw220diouQXMo2DHsxMkm6l9Vck2srpeC2sbq2JR+3orXVYaOkNat4uuXtPC
qX8AEV1dYD5N8TvURuZPhhgDkvrHUH4L7MHNx3F8t0Wimem75tPtVjxi5p+n2JO6
hpTYZ+N9Iz9Pfjimaut9b/RVkWbauFOHzPnLch7c/6NqesLLxmCSqQMOcJ1/yS/J
bK/tlggRhpYjpcHPd4lj81LTqGhTat3EFWQyPkuCevklj+0XNVQzyrF1bvq5it6Z
sLbpN8sCURoMeUOiZjS8mQ==
`protect END_PROTECTED
