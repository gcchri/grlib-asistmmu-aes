`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5AccVTVibW2Mxou45Olaun5m1A4C/J8kpANXJ9YizLJSOPTprz78xVau8wJ6ADD
mBBTD2usuEEtZc4LmbhZ+D5CxcLpZJD6xJHEZN8Lp/atLQMRSdglGgqw+8xhzaEj
n6f86+DvR1yMi1IjfEvFqCA+XgScbIbiiJtsuqfotuZ0aBSO/TjbvN62Zm39rENq
HIDR2pVm2Up9+qRgq+kXjSi3ukedwtuyzWPJ2qx46S+lWgKX6bTobydtCXXwM95f
ioSapacCo7Ddy/OrD4mxkAjAsWgvZFwr367YLrwf/B8N3n67KEjbCyJaWaPdWENS
aT6Rbm8aAd15OWyS4lIxvQC/MCjGP0GcCppOYUPN/i2q0WYeA4xypX2zkga7uJh2
6nvn/5yCWGPBbNrsBzSX2UZs3Xr1zZ0sG3iY5xqFgDAgi97m3MRhl52k9QI0iKL+
+qqARqnLzao+NpcDb3plvR8GqTk1h75oHutzRIzr9ChfQaYaaBqJ22+1/KOyn7oR
WRZl/XWNoufukNqo7xFVm2pBlmh7ewRpp7EcZh0MUg0k6c4CvRyq8SMDsmhJds/I
aYNp3AVfiVeuv7PWuG8t9zCSk435j7NuYFUKB2A+Bk24nXrF7Ddmddwn0rPd04o9
AtwwQA9sN/ytzkfEdKU1IzvCfbUzLKjcQZJ7RQ6hhB5k/m4SrNMkTGjF7cNBS+bA
csHzXiFNIFAz3ClWH7AG3g==
`protect END_PROTECTED
