`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ygQuLNIOJ/vhI4dyeChHTEMvjLlXe9F9BMGkZLbKDmmB6hQgmoZlVszCf8sMssJC
NHfhSYgBZE1d3S9l+SGSjZUtXmCvAqUHm0kBE5Amwc/lJRBmEJ12D/S5j8O20B4s
IMITIKYJjnZ3ng26HBZQ90k0RnY3i6pLEKTR16+20AwfYSAFZ/LV+tokCGJuUals
oO4BGQBOXSVqH6jQcTjmChbe3pFvlZHKK2u6wR36NG+OYLHXaAx03/1qLE2CfIYB
9ikeADQRhpvdUzUwAvTg02PBXnNon9VPXAS5+ozwmIBpYNspzvTijZFrV4n6bnf/
DkcVMVLUrsgs3MVigAx1yQhoF4HwDn7+/h2nVMCrASDSruADtRpU6xK5CRIB3bwg
l3XnivnvZzxrSVOJPB8GRglekZrNGZSejx1MFfo04FOxcWLjcXHeZB0noZAvlBUO
Xpzpe/tfxQ54nfRovAb9qwnBRh0n4t3CgM+UuOlnrTUk+LywH/twUneyHXINxq+M
vx5LnGnnxBQvxq7Jc3CamYROLOQ7GiWAhf68NkKBtlYaNEgAR32Y5ytcj7nBuBxK
DVuR4ijiG8W2r5Ob36e7hBaQVB1gU4RjG4/DLTwQdRX3HGO8+rRBAYqU4QOJtj1e
DyGbGayAh45Gaicagj7D5p7qxGcmcuD7z8cJNspCz5KpH5GObUXLuO2+O3/fXFgy
TD6VXSqQ5PqZsRSDw2AO/nH5zVIJVkk0Efrq1mCDdNntrieG7rSJWLfkxKYoXNB5
z2USepRXLKz+XrDNgKqcAYjrojBGN8toOyrQwUqMT/3WMttj0bk0pGBorW6tr2IA
k7fZoupqv1HV5U2UtaWsMw9OCI6R/iZMyVkRFjfLvFVs7yXQ2TBu4+JDpv97mhXn
bylfnoNFl3EQewjXPMl/IoI8d9kiYV9bLIGhehwd8CnW+V62/Fm4EiJDqgNEz9rK
`protect END_PROTECTED
