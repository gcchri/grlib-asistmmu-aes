`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpOREvgvqEXaaQ4tPF2OV6uvKv71BFah8/l1zDL/9IfFc+5b8ml1mgVT9nTIE1jQ
GEAW1j1KEpaQgdBv+3VLBB1x8Ma0QyICQmKKtT9DY61W99PQV8lHTCiLglshsJyz
vs9IQO+u2zkFWNv0zacgpTxAGR/mdn0jG5+oaJsX5o37N2rLr4eBM8YngtbCja7C
k/aL9cyseAXtHwh7M3+9ATxNPP/2shavlOyBwGV8EPMZyWzkhXx81BgYFRj4DwoG
Bn2Q+jKcXOYNiudUILawx5Af95UTf5UMI6UJtw0FdiROZr/JpTqFrVZPej8ssQ1M
bqbKY9yWjPb0IR3L4TzuEpZSpoIUbaILvlge5lZDB0fpv1cKHgO//HJ45uWFSIgQ
zK9vp3aNQJXdZilzoCNArhbDtvfqQSieO1OEUIyPMo51wQegsO2lkUHvZ7FMm/Gm
D6t+uhHztOUejLYNTvaryBYP30oVGk9lWhQWjN2L4rqUdO49X8bw3EE2g5dXx/pZ
GP3BRGlLZ+H2FsMwbPeWYMYIHJ4PGkPyr0M+Zqr4pMPpKWL6tuZy0bQp2ItpxRYo
DF0SSy3V+vdW9kmZmbQ3IxBMugUbDxYUkfGmd+ZX3pFYXSvLSsJ4pwmtnUVvyKiW
6IyWN0SCnQqJrPz+mG2lzmjWUfp8N4XcVd+u5O2cjnhfCI+xxcH54Der/ZmQh5TH
uwP7z4sxKhWcBzr2ugGpMjSPoLxTUkMDCYnhntjixcc=
`protect END_PROTECTED
