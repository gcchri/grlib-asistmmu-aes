`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUNVbH4zm9aXnXTvA4UvWL7rHcwsbA/bl9mWdRe3kQG14ta92QNydV7n9/1/yUj0
isWTqPhEIDtaFqMOozt55Yjn4JgoeX2Ww5KplFl7yTW6mfHh2YHxKzZvg03ps6NT
/7PayNAu9TsOzMnWi2ZYZuKoLqtrdE0A1kov9tNNUmkm4owKUwfs+yOcNk25yuZW
S+VLqEeCKT8IvmkhZ6hqmIf1cEdfikcQMHs3MNn7rCTsrwJiJxt9gHpZmewL1v8B
tvhzBOGcAoe2dWL4mlhj32W1tpgpuZvlKBZg5ATohOIrSg76JhK7/5W2Rm2mLxYW
NnUnuax7cUQ+3nfAy1hzxzrdhvhjBYbhRW4Qn3CF357AFMIgUB5drobGjL72AXBn
8TMDo3MAObNVyy5IaJHgqt2NOCVHr4pP8E+ZPK/Q5cjyHfu8kyEGaYzJyPY1GWme
R2JCUuysBfmLq0aoHQMPI2kGo/J8jXgsKQAxvtGS1VGofvafvsbKpIGDLSQ7Jgis
IKsZG+ShggUhcjaNrfmdvNaAvOItKrArXv6JhfTDt3dmD0Lwyx4DSVhpZDy0zK1L
1G5V/r6lDWPOe3WG+6PvdQ==
`protect END_PROTECTED
