`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTXmRLhdiIBAxRCsTmqL33oI3qFjWCsoJ817Jog+AcpLOje37fOl+Ir1Wa2Zw8iv
nfUkK/r9iJOUEQvEpr18Wti7ohMnRfrvuyFX03xGUNUq4tUGrtx8AphXwjT7sJfR
/R0hTDnaazhCLWrwMEE3NHO6MKf6fhtw/kEE4N/sG4UavT0TRr+GfzlALo2HHDMT
8R8oN1ZAKzqIjzzDSSeBN2/kLfDgcPmXBnq9j8o7zTztVCv4dYlaFJTQKh4BBl4u
GCDnesw5GsS/8r8mWyAGjuPOqoJODNwOJBJbiz6l1lHfIegcy4h7M3bNKBa0WANZ
P81/0edidgtGEsWsXRIKvLMXBACVyjvDN4+tMklZmkUfF0gUwDQ6E8pIb3Px0CNZ
idgtD54Bc0N8w8w7WPOVNAsbHGpeSef00oqIDkC0abLlvMTLLSciASGirY675Db/
fkNliSd3acqOBlrmPb73fmw9E8M/taCRXJnShx87gQXdOUIe13IOcFvumz+0cVR2
c534sRzzVJVMufazBhykLztT0DhI3qQT3SGv5Tx+NzF2xbKbSr5A7Suy8rUxV31v
keU4/PHa0f9BEo7YOjnVGnu9LaScy+q3DpSO9THQ+cA=
`protect END_PROTECTED
