`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
avYO3T6l82Mlxq/h0xLFe0B0Zcx/FfPYNbA2TqgHfxABzG6cHccEaUx7VhrMp54G
HPNpmUrMNFdK3bqc6EKZjp5TIhBwbcneed4NwguzA0IT3fuql0mYVyyBI9VwGPQ7
U7cxAnKDRhLJYe/PZLtOh6Oc9kcpCaDVezIEvD5f2fC4s8jVmDhopQTxr3BsFWnP
cJVFESPxzU7slgdAN9+YgNjej9TApsZ5aCsvk+9XHVAwIcjHisKavwDrkQqPwiAM
e1GUEjixsCKOOxhnN/fwhy1787mpNCtX9ka/tVAv//cv5SSmj1a8s3OSNdqXqOTO
uQjZR+n9r9KRSovNNW8qkvnhGXjotKHWDXMOgAoJ/rM4fOqCJq3CiiFXL3Ua2cXh
k2Dd2cdZI/F1j18jk2T/ND4hEzs3bO3CSdTNHPV2hpyCQ0WFcW7o27EfQnBTFeRj
/AF6GCj42Dwc4lmhTzyPidezg5e/JnInw9vxgVJKXK86o2oRt3pke7cG8gwZ3pF0
CDONm7LQ86C18bzRbTM5YX9tJByrzJlWPGM/SJuhy2qycVnKoWmqlqaG22zD8pNd
RHHTDus+J7qR30w0sZ6ICWxSgrfaa6uwQLR2RrLhqCguMNhDwoLBYFQdyMJm7Uc5
as253BSrg37UeQ2oQL+GtbaATljP8Do8d0vZ51UgJ2bn94vvZYRHrIvZ2KzEkg/h
2k4XnDIz/QjTheuUTANx+QNI6j9LPAisO/jykh6seiNbmGW8q72UkoW0TIdrCTUk
375fxxAewPVJGrFu1Jra7OfWJdOZKVnK163k0MrX2+QcuzzzxvwTqBb/YstliD02
SeCEOAlIvzrPxhp58d18Nh4xt1IGTGec0syrP1ro0xj00mubesNsugmkwr0Ecugo
DCAvRnOCESjQiLuyqfZ2cxYPelodoZPWgXiiA4ZYBsB0F1I0ZtcNNf2WJJ6cCOG1
ExbpEoUb6L/nv0VfZ5Z4mxKXW4VBzPSRCwFCj1plP9HWh3FSyqjbGWffxLH5Aibk
Qe/HoE+U8PfIYDr9Urs3nZVeZA8La2Ma222G44ARsl4vaLXXLhA/O4/QnRuer8mD
QtflQxDlfyJok1vFdLOz2ZvXJiLTVYcRML9MSzFogfKX06WjmKDVmf1OILBHspJe
gb5tfR36ZFqpaNI/aoXdXjxJwCNF3s8OiNMRu7hwpD8dH71zV7lUbqnavjRuZP+T
DGHKqKFn6uUFhILa3x4r7/muMowJ3DyL5gilf83a53E6Al9zmjJfw4tvp1kfUDfn
zkmllHJ/T8onUUueyvQ9MC2XDdVzrq+FsAp8Uq/iqB/Cuc+prBzzs2aqLIX+Pv+3
HHopx/pGvuxGZAelIgh552j83c3PIf0ffVUb8DQFKW8VTta800AZ95/X3yXlzlXW
Dcmbtav5KkTA5bdFbGTrZ0SXdIbYyL1jgAulMC8xjj9GjRJnNzR+QU8vfGLMS3GH
3tf6c0KyETsY7lmwbnaFDEfWeJxG+z2JbwgiZal57AkRJaIh2SVVN1+jSaWLUI5M
ZD3iAi2p7CDB9DK6j7AZPpxTMxa8Oe3QBtCUqHVctkxeglErjhV2Ah0IkssyDJHz
IYJs0bOpsQ88JgmRM5ZjDnnydpma1m78TfbCYPmkqEDOCFAWm6GMsAzmOE0EoPmI
GHW677NUoe1bCxnibMFMz86Tv1gHhitbOq/9C9B+ZBi0o0Q/UVpZhrAY9H1fas9c
kyNF8lgh+496UkWhzqPLOxcEbma2VmwgGWNrEpqWkv5U6X8MogceUi9Yp/ukNjlp
RkkW9ofYDDZuw0Ywj8u71LdZcKme8BrjVn4gLAFIPYecbPkoY4Kt0tFPTMEmRuUN
f2svya+eQ3bJ5bs9IiOE37dlP52oLVxp1J7WUrpXnfQxUibgTe6YyrPgARUp5M+Y
4T9TolpJXnFBoi0K5bw9IXBNVQ2+P83aLPrEQP6DRLB9Iv4yyXN/+s9FRyhUKGJ0
5/AC95q3bDMpxMA4Vj662vVJWkTw9oWfDeFrOOlsrgE2R8i8OZV5ry/lOKazr10S
J4jUrcsqSo4OcFbHIPc+g/qvZmQPAra68DwujU5q9UM12EaY+IJpD9fKVHAsHEhd
pVM5q6cF+9ecgKpgndX7DcwbDSVuLVCTFd1rFtzdKKxTdmybwNGG2s0LsqaUnudl
H/rxwLUuXVd4SGSPvsmRLgeTXOaUsZaLOzpB8MGydxL2bKVNJYeFk/zdwnGmn+6U
rpMWOUKHlKlFsFn7qxlvkr7Q3tCkr3j4D/S1LeEcXtQvqeUk5+9vCeoQl++/nxKZ
Mtb/TSiU8zJLcEbfvYXx3cMc84nO72xRaHnRb26GcyDiHb/d3unROmqrU9cC+YrR
c++WQyxVQLHEDGt41PAUWgBmxwbnUmPaoscyhXKW97bFXEYWwcy308TyxryOivpi
xsC/zh4Ir1tqlzIffbbZ1OM8Cj5VrtQd63FGG/PiZFLsOoEmMeJZy1skbJNfUqFi
ijhb9P/oEs71zyEJpdcn6pp+GCuVZZvXGgqyuGRBCf6b7TbigX6kTB93sTIsrC98
0Ek6muCRaLaUKDEwzVerUSosErRgMsFzqALBW0b/x+uf0V+RV0wKXZL1sF+I1KNv
8IDRVFz0tNqi/4qfIhGEqYWhvPAqzH9BPPRwfxLkqVHvjzh6g761XEWQgub6wm7R
fYwIXn8ZgspGQR9Q/oB4kcYmY6WoXK523t674w5DzY4OplLBm9zrkkc80BgvOAx+
RjnS7HGNl6ERtc9qAD5dGWfAAb8MV6FVGsnAz+tVFjo64x9ox3MDSqO0R2HIITrH
CiLoZdf2K7r3cbSgyD9nc3WBB+qal7TRtNCJACfA8dkKSSeVXe4xmMN6lHOBLjh5
oiBBEzlWkAKCHIEfMO5fmiko38BPUTuQUeWPfL3WnC0BfvXIbpUT5ua9YwrLiI24
MRHOXPSIRBCUEbKT2yAkk3tHQAJKTmSkFrVoj/xxnWOuOH9AnJGqBS6I7EZ4icSI
CGtt5BMt3J9oURoh319ngqEqYoTFRDYsrLtRQq4T3KbkdvAzwHs6hlMTsjVpEb0R
q6NikMIi4QSCPmo09wknxbB0yqfrLSX83ZSCLKQFLRIGGfBnDN66tc4k0Ubu3tgM
xLCUtmx+1UHB1MHDsKBu2SmD8qI79rxwFkgKL1ADTukI15pPr48Z9MCWfwiPER40
Dk6UpT4L85mGOxkHI4V+o9fFzyowCAh4Bue/TNhvLarQaXZqmYx7/51IbksBo61t
SI5VZ3nJ6wJAnynAZQSdI3Y3JmpdzBvdkhD4J9Y4r5wLUQulSnAAQ7muvYXgNF3O
zEHnukIHMrCIYZrQvy8S4Z7u3Xkt8TdPd2j09RldxX4myEHxftqCNnjALSHM1cmv
xwPmfvo/P2TEacx87rzvBofEucYwz5MAz2+Hb2elPJJkWZoKI140AwPW8Ouk+PVh
hnZ65S6Yx9W8afkyZCLRXv7EvjV/PQfjEQCDqjGIg6yBJemyHfSFzpUU2Ixaw66D
U4AhByFfSfuOpw7uREWOpey4xto70tF27y9vaHI6zJmy85F5l91vTdet8IjKc2vl
Ci/ODu6K1IlzSJ3qHH18sZaDdEuP+6FXJerGgkN3zAZbqsrCpqUPP9tO2sTAtnbb
ADYSy5Ht/7D8Pi2Dyg7kr+qUNHE3GEb0pno1TpCQ1k3H9gz8F4fSc7sh6aK6iJUP
YQrwZy/j1Vu2e4zuNt8yTsmTrcJiH0eu+XOKQTnaPQSIhQz7ZgVE/KMftr6mVE74
hazsPEFzmkj2XOcBUSyQiNFX2n2mUCNaZzphcIgiSES5ecqcyvG6uDqWvvae6Dlq
eAwoCWcCRseXnD23ELOnstpQuGtycc8grm8b3iKto+wJ2av5tXFlUQQLl9D3dbiQ
tCta0QIrb/vyRmeYw4e42W7798mL7lr7E2SqdiJPF38P3Cnu6/gJUu80PdxtR5Gy
RAM7fcUNMmWQep3ljtoJ1HfucoB4xNF7bHWlUJO/Zxuxo6Wl4KT7C16Azr8hbw/a
IIgHv5DuUn3QIFmo7h5JvEayd9/2Z0/na7U4+HU6IBs=
`protect END_PROTECTED
