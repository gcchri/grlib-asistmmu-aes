`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NbMEswf53NOIPByVcDwalpNT59jR8zl+Vap4FNwXVz/MjuKMzpDZhEvcKM0ozlFI
XYL0q6N9fi6W7thSKTBjtgL/n2yIYJ9GB7AywypJLS6HQOX2hxeFSD3VU4QmMCw4
tOd702a0ZW8w7I5RuQd09+IJhkBA0DM/It4hEiPAAeXClPlUZpBBa61GfsQ9MMG6
ScbhQyMbILSkMayGM8JfMGtroCJ+ZKPCxvA8FOooR0oGDUfXnf7WQ/WQ+tgh4QM3
F0pPudsS9gOmNmf2AJLqMlQ0pBJ+KyVEMRAR8yIEWHHOfJhACpTSTvZIh2U91tZe
DVhwTyXX7qiub0lWH627JJF5sVYoXTUuB/DQuqXVfOxIP93jxx/8MBe+jihQFMLN
JHV1AdhDLRlC8RebSm9vMqWTHf52k9OQgZOUjegChrIRzUdX3Yvy0tm0vxXx+UiK
VXdVjNnuK4tz8hzG0ImqqTtzn6sQmPCQhaTMDilcJy4=
`protect END_PROTECTED
