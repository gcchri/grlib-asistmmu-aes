`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LET7vQZyl9c+Bg8lWtPPTjvFiCnhXUuDFujnDKRAScnL1XB6BL7CrySAXLAV1CQC
TanSR3nHBLSLBX/VJiNQkl0HcPWygiZ060tKO2CQfMx2DtWvtCMkep0JUSN9/Vr2
h8IHnltcMBDGur+RJ+vRYOtZ1BWdA8RmjgcrkW75VLiDaBwZ/qVH56tDoVZKfoRw
wciGsPtwJYQUHoHqwBmqAdZOhmaEW9yfA5E5euwaQ07GNKURbotcT7sk8jGxBpy6
h/c0sAxt2Qvnn6B2fBpnVA==
`protect END_PROTECTED
