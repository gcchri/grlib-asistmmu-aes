`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GC/TgS6OFIJgvz8dfuLamC/KvALP5qUAYhZJoMvvj0eG4poEGQAzT6DPJZ/b28H8
mPT6Ht1nKksHPhitcqsMjqgaYy30viYUvvCU4gh8pqRZddgFwjlNSR+FyRdASUkX
3L4kKx8Lr9lHEdMhp0dm3O5mc4/l6g/2O1aV+3mdNQMBkp6dZnFF0f3YBA80Ks8G
ChYGmeUROk8N3Zcjys6RikUiX4nymmQ4vkDNgnHBhTYDKxGDs96Ywi62HfIOkIX6
ZKn00Dot4HeXxX944DXgAvShXzae6BfBRBI6yfTx2q05nsNqOjyTNzR+SZkUHFD4
IRsn33j6FaFJAAB1ApbWgbhE/gY2amik4DYc2OanQPYX7V0RFZNbQqA6szat5T22
+H1+NnqrWHFgV7H7yy06TnOjEJkD/WnczOM0eEL/pZGBwVfGWydMKqzqUQUcQ/tr
FwidxRh1vwroBXlRELrqCnDC/mmdHeIkLilPPJoQB2LzlSkCUmF4EM/ZJ66M8w8z
EMwg7apHwCxzgYRyiH216CKdgYyobviT8hKBs7iHfe49YZiiwb0xawvo4fceKRM7
hHFFn1MXsVOmJtSBo6hZlg==
`protect END_PROTECTED
