`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNERb+c/AfTj3m0341MvAHZ6iAl3ran4rkbe052lthCQMr7BkirTnVmv4kWKfKyo
ZLJZQlaaHfMUq/YgyiQOl0U3ePyDkE0G3cfzh9qo1DhU9v4nwDVXM9SLDYz1+AEy
YgvsxlFTXrMyQqI3VcmYwA1KLHe/ETiCH30XgUOFqT1hASbcGwoITa/bht3SIEr5
XzIUbfkYpncFvEvl2bQyQTRFlRULiYv0Qq63wZx+hO3FS59E5jEpH1guCFnTe/z3
ZNGkCUuEyNpBFzl9TriotN1rtcN7ADsqFfRY/ulP6Ia/6p3tAhJzjqlgu7y7xe2+
YYC8hwng7QYvcpTSvBWa6f/rUj01Ihm5cxDOVcBr+gWIZTUm7qLaS3QMOUgctJcN
g6tsiyEp76J/GrGePURgfB+kykxuo2xRbG8VFkgNypu954LcT4VzxO3BRmfMSPvl
`protect END_PROTECTED
