`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQHG2ANFaEvEzotJMNFuLSBV5XBUKkxedB6TaDD241FDrEf0m1V+yiP6cWJRwpfV
Oe1hIWzidvEbCoRFTZa+E0C9JKh3Q7Xn2ftq4asiKin+V5k0Yrho5SngPxP49arT
JT0ZLuaWMT9sFflyFgfA97zaAJWwfjlyTj9FcCP8l9z3ZqWtZhKgEfUJ/77/U6ib
5z8dq+o8ktRvNZ1MhnPjyVExZoTw6/B5rXlgHHyj6ueKi8NxSzW5ARPAWqBOHpXx
zob+imsQd6SioNC8YVMqtKyOLshPmvPBa798dVigoBgvVsWfroLrGHZ5CiB1ypj5
gOBs0oR1EQj9Jpt9AsgI+035L0Ba/I7ZiWL14uK65Ia9oiCFy2PzQJ9M+rHKCElp
ZsR/z7TSq+K8uMkVAXzSVZWnqu3HiSgZmbAj196l5OSy5r3Q2ChJtYDcpQHQ0zBy
`protect END_PROTECTED
