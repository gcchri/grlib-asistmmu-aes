`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y7Qv98QsYB/AO4fVcYiaZ40/HgBFBtnmWOf4IT6hgHJPWpj+68RJiFN3MjlZkRgQ
NZkJhpYOgoP/ZM8CfCA6ascL9540p96ZH2WBsZepLIRlLklF8CBM+W5iR5Eh2z3i
9ZZKaUDItyNFN5s7HArbUjVIIPGCbDRsNsR3xOSGNvs79b71uTI75g6BBq+sdP1x
MbO+L7E8c2vYSFxChmk5Jx68ouPNVEJsBl6eQ63YTxR3D67DVRhK8IBaBses6DLo
sM+hjjogHdyJGN4wz4Y3DcUSdBRagI2x1OSuNm8tYmp+wtHEWxZfWo8iF49vaiKs
o5vt9ss3u9xJ/AmpkhV6SkhWjmullEXMpK8L87999ORSYC46d1Nk+shEJShJq5gc
Q/hPgy1bRLA0Fhlfl72mp4ipmLMXr5eH1h5C4aggeWwopKfpnM1keG/OxcsNvyWN
z31hrEZSfOJ20CFhc78LEduCcT8w8JvuQWxUg+NWzriYpJDgIfpX/gHbYoFdjp9+
GonslBzZL/Gr4AvXwz405zChw1zJCSY3VpnZikT+6Cminw2NWAnGFM9CSzB2+xBk
ARpIdGcN+MKrGNOUGEagipjcIBmxzwz9wwkkzvRhIkNukDJu2QiP+ea8RWlIB32V
AAU2J20SDNofyghbYQtXCXX3va5AoaD/IKmUB46vIMcnqmBkFhcBLDdpxo7mWZ4I
MUjw8FGJZq2e7vVsYhMsQa2wJscVjuYiLgEtFhCw4hiym3D8wqEEw+fSFAvCbELS
cys+J1qnel9y8q2gBgqmVq+TTCtkUNA7Z1lm0qF4bm1CxsGs3GGvKS13TNfyhLBQ
O201LNf+Udf6BvJJki8V7Fs3FKHV3MGRsAsBTsoNyqkWZZiJW37yA3iUt7nHP77+
3F9ge24d7+fuyNLvPzNd3TII6wFc/GEP6BUCW0Luk+h1w+Bd4I/X8Xz7rJA0qQ9M
tUa5zL9gBc+FVXlmiL7WVOFiMaN1doFViOXiG56UEvBc0EVhQUSwep9PCSqU2V7O
IpQyPj4Ju+MwxFN9fs0tBQOLFpumE3xrV5l9cse73uIQZ5ec3fb3j4f3tvUp8wBa
37dJt46mBhZ3LgUg6fQUqrXBOP6rWz2B0FWhwc5uzgM9GqsD856tFPSC5FrBprRS
LylEYnsaWD6/fd/DcBZ+N9CzZj3/HBeCdKNkJ/ktNdRJrVcsLxsXFM38k3UgnK40
cEVyZCZ+M/Y9wi4R1h2G4aoxQuEvc24acpI9wOYlFoECEMBIctDM31vHUt+dbOTM
RY+IloL1YJ4NMPSAfw/0lHuJHVjy7G1fUXkCmGo07UeA8TKkcGU2RT1YY3I2wZVE
DYoXtrbjzyRgulz0x7koZrp7vVF4xRXSKD+i/lxWmUH6fyGrFUwcU3ez6bQtCgt1
OmfYoU0lxKWSERRXFWWJRikdHaVDoKBF80cC6TrvgEXsp0nZiJRNM0etig/ltqaR
Jjx1acVfZ38ERjsh2I/l95zPdgYcM+UdQFgkRV1bXeTcYjDB7awm8Aj/ANvk2Eby
E3QPMxOic/YXRwzf7XixAUZocKAs6+pvo6489rvtljra394Dyz8c/R37yCj/2LZY
VnKFvGzdtCy7L/VKL5N6iu1icmG88VRFvRTZTKe2+1KiXITZJz+XIVDjp1EYdi9h
UJ4ufTuY7rKWoT5QAyRP9DcwsJJ0DkId4haXGanN5NU6vvTqJwOlCJAVrJ8lCUPk
myMK+0cfcywtPOHlPz8L+k2xOIfA/KCcyyB0Bdq4QgbBDBbq3HDM8yajnDvvZX0l
1OP2j7sZYNKJYGaJwC1hepGgQ8/IwvttPhduSrIN/RbccbGPdnBNe/tBVgAXQMhd
T6Y9J8UIgXfAHqg7QVXq0Yj/8BjhYUwmPOzc8cRQZQjWqHm7PmvAC9C/AsT0Db/E
EFJ+cqsTI/y+HjoeOtFaVnJK0gkDvkVX4XCX2hQWzXb3uWUIlgq6cUvZud8/NITw
cqhFgVLMBS04g5hW17NXF3NjJxnvae2qVt2t18DHCvRWOZh14vdEKOKqdspVreom
DUINRdXWBVbRsf3rSkQ6pjAzT6Or6AcjTGpYrYNM6WYxdRsBqxASl+bxDC8VwDPS
TWhwb2QiQUG8KnYAiIgDU7DbFdOqkaAee5BrbMzdJvMvCklHdIxQlXCx1/5pOR2z
GDz+5WE4412n3Hb7KzBsBtisY2CVWa53Q86S8/Pu0MwDyZtrTCmaZJa/lKGnnwzz
UoZ/b965MZOiQJSMfJja8OnDkwd6aWhrGdcaILe1Vw5sqdYUIYke1yIMsVG1z5z6
EMxOw2zeePP3k1Gp1SQhLe1+hvtIsMxu9u+sN0v3gE1L+aW7eqLlxnA7ey1rFXb8
3OaVJKAbMxo+iRq/mA1cKtt/xZoY/vXZYBHa5WluXIkbJKHCkddaH9lZyrEpUJk/
ehh5vQ9Mwt8LMS420wJeQQ4fBw6qWocdhzN9CuziZrTU1INiluqKMf6eJ8rvUp0q
cx+sacDlHgAbq1iYaKqBiA==
`protect END_PROTECTED
