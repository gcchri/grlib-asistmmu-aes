`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDSRBbo2AX83FoTMQ87jPO3Blw1GJYQzOeD6oSaEDY3oWC2SXN6cwgsy/cbJ7VHf
LjFH8nbnk3Auqzk5ok3sTq688pVqi/qXFM6Eg49ikGJ3Jscqo95gDhiRhURly1kE
B2g+yM5ehUv9wgA/CtFINnIATkIbNblKKAlXRraUup7N6P24DQrAvLFJAHv0AJ9Z
uO8z8wlfw85pyFtVh9ww/EMJfi0855OftD7CAQGothGF8CrbOp+zmWgrkpsJNWfk
uleCL7XdR2+q/MN6jc2QrgSQ2iJhZSEbqt3CEaFdO9T6mpk7yViMP0vrHhyWJ0f8
GzynJGAewW8aPbyQ0C+cX9iSh6y6mPEms2LTMIqiPyXLGUnftlfHYqTVPGJwoQWi
ygEXO/cbAF7E152DDLCk3FOen2Y6bwOFlLcvxs8GOZoXwACxHQETd4F2QAQzVH4q
rhxkry6ckcyCBNGXJmhJE2lsoQJ8HlxykOQIzPrssJWjQATihV9gwnKzDNyY/vJq
7bEM1CDywNHTYAEORdQCsQ8lJlKIKRv+5rMw10ll1ClZRXqiD56zJgWcZY4ol3ZG
kLjTBoN3jcv7aAdN2yi1rrGQxj0Cv6tHIZ5W86dxLgSVt0RMJRhwvUepk85sddkx
sR0V6l2NOIEMy2Vlqua4D5ju/ELBEujLybiExYmFPlFAW5RAeyeS4oOTxrSXRIgK
yRkeI9gap2iC2uwEQBtewzECs9s0zh20OU25W7tO+bZErxM6TY+x7iBI5SulQJMW
og3FtadZnQXQEUahsRY8uH0UqA2tLWjRSUDswBoOj/S+pXMcksUhLMz+YcIIMgo+
D5wvA24Hl3cmBRXRjaM8Vg==
`protect END_PROTECTED
