`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2kMUxzd2y41BhpbV7dbo/jXjFvpEs/LC3XYKEkeq0/10EbfpQNGgVw/L3urtilA
SNmcd1O6vcJ/nyXbCNCHm7cWIHX3KMtBql+a3QCaIJ84rjRBxHSKf1R022olANUY
SysEOJ1ozAearkctev54SrAFtUjUilkxkmVX4r/8oIlPrGN8Fq6AHFZmvvUkVMpc
wK7yRwwD9fLvTG87JgtODrjOaV4Wn/0n/kKXV82CbsxmXz/TH2oXTgZGEQ1U0kLv
`protect END_PROTECTED
