`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ff2mrL7AzgdUoCBFE4Mo2DilkDHcAanpMRZssR6AQ1FMY6ureM/ga7R9egAmh2AC
puU3nNEz0qhuAcbtVq03cSzGsFnUhQoPbs/DOt9sPLNDLvcoL7N12msUpOn3jJ1z
8T2Vmznt97SbkP7AkifhJxKIdJXEb6jMFAjcTmNhgXcy0R+6nDl0L+pbBFDQWfLi
thUHJzeTweZ0Q2IHX/bd6zzF1qWcyMske0ZDibpLvenxTkuhYFJxGrZYEh84kCDx
p/pkf75C59AJFUwwvPMiEL9kxLcyagvZQ0e1ATIyxvOfj1tbsfKr/T0i9zaoIhSb
bXKdTHGjjnt7bN+wDIQxqw==
`protect END_PROTECTED
