`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1PTRf8T+l5DJI2gi6hcC7pdzymP8SRw7tYFB2RtcBUNF03vt4wDgZVZ4+jOCdfAV
oau4t4I/pvypfSdly9PjikytqhJTYZRkzbcwfIVQZNV7Dln7cmnl7yB0SvwQdKZ5
FDjq/ZjAxtI+OYw4rF8S66shS8yiAQ0cwsuTgnwtJYPAhTHZDFdO1BPax3M5G7D+
CL5eNTYtSY4hOhDWzfFbWFz6pgG4Yi826nA4RE4AY9/Yo2EhRgw34DwANM10M0+D
lPhc5uRzyOHDavYIVOy8Oei+s6JbqckcvdOLb7f2LcGrFMIwE15kz3WiG075yRFi
024W4664sdC0qbSPCSrvVhqf7hi/U82ei3KQCnro9OsfhvE4weHAO7XPBLc5hYB7
7EMy0NmkwfFnBbV5ExnEt3eh1qa3BdhoOjle/Q29CQ4aiI9WdFuCpCyucrIHMPRU
`protect END_PROTECTED
