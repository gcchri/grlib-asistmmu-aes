`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pgu6tG2mSm/jZwF6h5Y+9CN13rdB03VgM2eQ0YKfDNqtQbzrKvwaymcuOon3csOD
0XrxaQFL4sawovMx/bCTrg+zp7ZZrgjxQ4VKTiOIfqSFfoJt3ELPheQ9VIcD+Jn+
xL1SAtWFUYMUr4cUnFTWiZaiXK/2LQZ1tvj8BrbMtQkAjdUmI1bYj1c5uo0LGbJV
O8Ckvz4S2pVRKszGMxMoHSCwB1IWkqkh38/ELhgodLKT8qgesXED+z5BInO7Q70x
ENM8nsBSfkvw+SFlaGJb9GzudCchoJY0/A/gAtiyt09mQ0KuxmiKtLVVbn0gb9U/
syGdWHMUOMtEOHzbOh5H6r84t7ypV6kpN2RVbAvyF4R6XklexLXAft6Lv82IQfGI
B6WB38chR5FhtV3DKR/36rbrmabRF7uGxDWU7wT70LTxO7GZz3dNxurDnxIfkBOz
dCwBw2lm0XnAyvYtld4deXjt63PrRoDTRs57pFFixvp5HU/hJZilV1BVcSoFvb4m
9ipY4YmH+0mKdEewlzrK7IahnLY8zsoJ1BbRToF9kcU5kZCUsE8wJOsauXUNc2Qn
0IHG02h7v3IJ08OkF9ezxPKRyvkTPH/yCiTfwCIDeNG7OLLR3HNnl798mBVgQ9gc
gfffG6IdWbUYtWqOAoe3i2A0rgq8ADbsCDeNW4Ap6eAdnyicLTK9cSN4qF9PKs27
vFwXpSGdn8TowspoECSM94m8ZPGrZsyr+/yJSJRMBX3eOy7r+Iz9drGJKl1RBe1j
6r8aYF9VXuys94fxhKfaCT5dOnsSBLrCEFbT6bm5UaK8R1FVcDHk30KtokfPXj++
pp2IvVFVpwWYQm5gcH8CHM41Ie4qO4Tf0/G/BQTsPus+hVR5OrCLzqt5RgG/5Rns
7US1YsFzRiKho2KY+RGmYR21PIinyi6iqw4PYba+6vQmO0VnIPLj3Q2e/HYXJqxJ
4b1vDTYXdEqWiFksKCLQrHbLt8sVWXTWPDVTV6dV4TAEXj36Du3V3Od6XqXTRGqJ
QvvLf6HOEsiu9RmI494V3cobwasl+1+frdA6knSnrlHTxEU4O3c50w2Ee3r4x+e5
SdpOJq4o3zT3ewkiiGxqUMaFu8cDX1NVs6ediWhv1tQszs66x/6NpG2ogAhQShco
cdrBRc5MSwTYoR98783Z8zPMBpSwFqlZxR32ZSCUUvPfPxbTCxBbzh9zVVMIt7Gi
NZwBr2CRlRzCZ4vbX+Ctz/GamxkTZbUN5fRBROtO++pdyW86pb8Yj7Bu7QzqDh7L
fyWZgW+lItH6d8avPTcVoyfL+c/ndnqtlgb7oXPrD4uo9i+oQohzukzWXuGbAzNY
Vg11wh7tySL8L9PzFU6gWXxs+0x+9CJguYBFvkyk7KCtFgc1LPL0uHUz75QFO0yN
paE2x4rDKrw++ZLAFod3dA==
`protect END_PROTECTED
