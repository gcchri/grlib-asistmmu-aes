`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m9F7p2phMN6zVfT0dyEYJiGGbSU8xnx8SsQmsyaT8Y0OJU1KvZWarj8Z5O6IGkGR
eggzaqQzcjSve2ICv77jE6WimJv0QgKi6RcqUoP3bild/EkGZ9gBLgPoh1q4nFdX
Yc2wUK3SfY6RkVLj7cpMVrskkjCnM8O/49LwQW4Myzy+3AOnIAUztTCcFrMp1xvo
a2DpGVcOhoDDRq9NdZe4cw7AWy5BaWrFoQNTVPaPBjhJ1E42mt/24WTAvDKlZHs2
ltM/s1ce6YojSFqBqLzcFvEEp/FTrnDazKLaBdO13yUaaDZGv8qCRrj9G3QrZv1e
W+qZNA/Z4GaoxqDSlPd4kWjXh8EJz+xl+ITxKbznoDM0c/0The3sdWLWD6YS6S+s
aK4D1jUwTv1LZFqCMwII2k/Ad9jw9Zfqrp4THg2FoH4dU8tlD/EN4lBBHJ7zw1g+
sg2etwrUc2+PgGVfj9l8X08nslmr9eoFAGgpQoUFea7TfpabFUJiyS3gw0sATugI
2n2OXpJUObp3PJOIuWXRqm6ffLos2d0r/EmmPSZArDc=
`protect END_PROTECTED
