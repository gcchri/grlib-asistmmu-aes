`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJxDGxh7kle6GMcfRqXHtJphh54EhkADto/FoDBkpTZEkfA+6GwTnqPNe1UJXkjf
+fxJUl565q4j8pjCvPM4RXgEP/vpDLf/StyXw6NGE9Zcmj/AmUTJB3+iPrRxAWp9
B8CArk1xndFNQ6oSgvA29xDlfUAmWxsEIk7/BCM8yfwW7oHicnuMrdfiRUDUEKGc
BNfPTdn6OkiUz7mAO/+SVuc1TS8no+ol++f/1OZinA30HGfFCUhskM4KMYQgM9Ls
f4J484ksZLc/WyRSaDlqhKtgCczIA97jCh6ZYgJUUgSPe8xHQ3hCNja/P/JD2znA
alhW6EG454hBtr7mJ0gMu6cYKbVyeiNI30I4gCNS4V4hDbjAv0XZ6d+ZSu1cM6EZ
UhJfpsS4VhbGTwY88kQJb5Xt9YqMW3ly3CZW5cHgz1/003wWHNYunmB3HOA0vkwJ
T1JAwn3hswR7Yk1vcTiYe3hyu5aNJT26ZgUQWraSW55uBcm+vYZM0BXIS4E4DmDt
88zvVy3yLoMh4sYGqjgBZFsobghbZDEcEq+A+KcIBgBX/ikMdkwELmD8VO12SV8c
IusK9Mhm35MXS4oQvlg8Td1G0QnImZ9VsKrsxfRUK2Q=
`protect END_PROTECTED
