`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7095Db0yTYSYKkCbsvBzTyrbM/3YIpers2koHwedCnf/PLa3YH443L8spd1vJHjZ
pxfmtdz9xgghL0mfsf1GPBGGYFD37MpDuFwfa1+5Nipke5p14pxFsYKhYZTqLmpI
mqjTQl4+DX2rD24cZ1EF96YffAd9twIA945rbVz3GNOIrbnU+uECL6uG+c9bZ4aJ
eaA+6gcDqWQmH0CkoRR28vZeKWEnSmpsvgVV1Rz2kYteRb/qr9gAs9/Fzmw6PYtS
A3icgsnWK+FjLBx7VqC0IH4uCAQqeL15lq+mA0qkLkDbI8kvQ2yppSFYqUlsb2/1
UcJkQGTxWoXW3p3u6Dm+zc2xjVexJMStvOnjalhJWVeLR6rB729vd+TfmTRUXwZi
OdvYGGNoeYY+tCH4kwVC64GxUInn8NNXIqwsOKXytcYC8K2C+BT0MIQt21qMiWKX
KsCGW6UcPsL6MGX/JQkA5jUxSCaT2V2RvvQ80K0/bucMj2qZFaRk++XtHloq9p56
7BsHTlmzrZsf/tPGRjEsCna+U+GacoAUBqynhf+K0AUKDPioYnUqILPaAvhoMKuq
QnCv5/P4UQ5tEccW2lUbT/0UUQZqNveZkXlhmUd/d34/wJXLpInpkBcxEm6wvCji
yOODuRPi35OYrJnphXzd1khDS2yKhFX+B9t/4lb02pv/6/T4wzaboIFbLVAzswIq
AjionO1azegNJe1B8bMVDdB0tQpv0XzQv1IIxq1UnSU6VJNdRHSwO5RfU7QMxJMA
3JTW3AKSpWM2PmBUotNSmdDsKn/2EZXQChDZQ7LGx99RYAM4WUCJiLn3XGrI5vGt
RBO7DgPWZcCQ4QN8tBQKsefuL3+JO/SZt32tIA6DER+lJ0oDYS9PqqgnE5QR8Dk4
9PQr/uBlLmFx4uEeVcKW79w0UnzUnqKNm57YAlX+O96ds36gZehkX+jSfai2HQ6b
m0oj25w69M0jRJT1vz3+0+L+y9aOTFWMNJYqqG2T2v21Y9op8uaG7zS4bKU70Q5j
NR498vjSqGdPsC5LFeIDroiS0LZFuy6pTh2dV5eZ3H7Rvdw2LXilm3zELDbL3BGn
kTU0/gzVuM4U/OWQyOf3CNuwfwLNeU5xhRt20JU9ylBwwNlwnqPBPkqxciSbBWGF
gBl5QCEo+0wsoF0YSIGLQMmdJmsJquBT7uvsjsyW3sgaDFvVEviUgOthFt+g291o
o2aUUMavdS7gexCVVSusz/7UNuJ7b0LRoV5YkMmziBGsk9qOwt6z0iZJ9ZD0w9RC
Vco4lRMFWnfY4LlUh3WDKEDCEPe5NBBo4IxISotMiIE00WFhlHFO2Vjrh8MQtf6/
eR7pkUmhSoPzvEFx7CeD5ASFJkSBq6N6XFAnTwu2tdqg9Fad9iiPotCVbEzaXo6x
5LDnre6EnKiz+ScpqvqK7u5ek9saN40WhyT9om6U0RlIFRVT+0SyWndmmdW8j62p
OQ6tS4kNkjLg/jbbGDB4YiNQK6J3SmguaxeQ9IOrArtgfisTin7RJmn5LmAA+B9O
NqQGAnJxN03K0oHpClRci5PSm0Bag/+yd9T/QKk2v5B18HyiuX9kcmEfEB2gAK8Z
tC5gunTzn0UXKUkDseewkVb9SxN0Gbo401J8TCN1hlr8A29dtWJfVYQu4rWmKAFO
KqKEA8TqZZ+jSWD42/QPdlG0cW1H4PVYTanJZ3Z8eEFzLZbOj8cUKJ8tw4xnsRVZ
NjRq4/fp6rzpS9mC0djFachtSlp0q1pmrlg7hETMcH/lfDgBwKZJ/2L3n9lDMZ1I
JVyKv9rfW3Vz2Z0qA4WcRLlgR7mTfYJjZSGZxcmPTa23+lfTj8nedh6Ack0nu7DF
qwnPhGz9GcWMqzHzN6plFp8AS0/ww/fIJ/A7+YKSp5lL2QTT3y5tdJgPSTCO0BOX
8DZsCLXTjkM7KTCSj6MhZXmIvnl4PRawd3u58OzdUwQly6TfgROQjsUM2z0H960j
uaAXVFhiTpmxSbxQYrNhVmCM3aqtpqGu+6jiTNU933FfMy9ejCosMBvv5waPkdT4
XbwsTliJ/Sb/Dz4PWN9Q/gqvUgFTJxN3g3r+GV927TTqXrBiZks3gjWIThCnMvf5
oK7OFtXz51yh5e2nvymoh1TU1lXGfkFhaI79JUK2d0sJL8LxTRrsnzkv9vLnqDZz
frCKrvDacT3TsqWfKgxgoacVKdKUApxf0CHH9LZnEXlBerC/0B02iDniOfJ4JzjY
N/EoZQYagF3s9utNjbYUHuKgNXTR8uBft8yNrn6f1pFylmpHHaTIdLluV1cGAb2j
HPzZKHXZL2MrlaUODc8EAFOWmh7wC8E7QbuEg9st2BOY4fOcfs7qBBq4aztgFqa9
dv+1nUCdNfbN2JHTEpee9gOb844W6oy5l2jLejpO45bkLIQLkYLah90e/XQxmKmc
fjZgAa7ys42r5qmaJUOol8ag7S+ZzWKhxrv5FYAFZLfoT9J3TdrLmleiEDI15Act
GsBrRByUdxmzjSUAwEY6LDdX3fg+hW0/UbivwOn5EmAdgKD8lHs8Ncq1XY8FDFsL
QuN3njMgLdu7AbHrzu7rVFRy0ifHZl5kiLJrBbqYh0M6s1cAZWoR69Q/FXOnELej
XHLPZut74ZsqzUnFJCE0eBXQ3jaSEdM76nvPDlmOdKBNf72e4DxUORBa9Ud5D3+G
sBHJulJPUMIUKa7GXMAh4ZYF5jvAOiD8liOs7clWMWicLMMSsSc+TmD5afEcIiBq
gAU9v8Zf+Xyzkma6wfnMXA+KyzIOsIFUYUpKjRCLuSVPwcaEvSHqhju78lbDqk1n
fp6gUZJj3gH1ZCli0TLx7b+6DplDblshQA766iKnhfkCL9YqevpLzqdR6m7L5nGB
V1XfGhdWc8Blm7fdKCwamZ6jMuNEqDZMxHPB10f7EgT6LK+Uiz7bAsEPyy8vcQf7
8G3+jGiYhJBfzuehETjeuZu/laKAiQfWJ+NWlU9vS394JXW0P08uzfza2gixEC0j
KgCa4fdXn0uOK+ki20U+LHRL+Jq4zbRMP3sDCpKYM8semUCuYvxC2/SabQzaZqS/
HCVBvN4H3YrZsaGKiLcgMJ5Wj8nLndSqEG6QbZgExqLeE+SCd41qe9BiUI994lkY
NstJOB7nlTmFT2m4e9naWvRCtjmAtsfpDBeG0WjTwvdY7uNt5N3NCwwFbulLoYgM
ASKpE087FuUvwCjSnlEr+iizjxbEcqFbwtTVIVAXNDu3Wx7NvxgPAPSQeWHogbZy
jjlQnKr3p1C/PvJrSx8WcGaENeNIkXaVGDfdtaOxYIMYvqdk3IChmHad5sEYX+Sq
YoWu3W0qQq3um2WvfE76ocBBJhCH93pmZhA28zItgu/1Ma06cKpHOM/Fz3w6shbN
kvp/aI3t7WfpUx6cwWS83f4Uw761yxAbdwlGrAf62bzBMQD0LDnPi/NIUqXZmPY5
Dtba2xPxH/mznB22EtAwcKJPoR66XtgsekjS+gA6r7PYCpuNaBVA/x8LrE5dLkif
b0yjbmVfe5nuuf5GflukgjPWYwkfwiHMibuejyGKmYTidv8QZdnT9xUKIbwwx/LX
vKxFPm2P5KJgEfqBTDmQPkHoaawUHz1l0Cq1rD3LR7n05IZggkVDV4kqLe81MhyZ
zHjGKt9jk1O95jS9eUFvrA==
`protect END_PROTECTED
