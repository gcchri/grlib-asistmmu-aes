`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dquIOJOMJGENfbU9XL7p449FqY/T0mIA3jMWOovgzwDEMjokDnyD77DyJQHWatos
OlU8QYoh6CpwkKAO4pKy1C1v59YdJavILzWfDXUyK5eEV76Fu9LoD//+JgRxICp0
G8nXZkZ3qtxwcwFTYuqTEvlru8ki+wAfvFPb6LA95D7SAQar4z1YaE393+5uQ84d
N3pw5jwM7BTOkV4PQScXvim0oH86KCqM9SNwxClUq/5bRqm0tczZ8jHAz9661GXw
dxDJpHrjxkft2PXJTflbNt0vjeGcagbYXviL6jVvQDcAXnKFR9+HPpUqmzHZpnIM
Ds9GhetEiHJeK8wzvfhW3Jh0TccY+9rs8AS0TbDkyOir9F0Vd9Afat5buknCO3xr
w70FsNOxUgFytetkvcxjKMpAZAImfxkRzVg/S4XfZe2apj63G/ALQ19f9CVeZVpu
o/SYaFm5s431ZGh47dn65sIIIdyAvmT9NENKCIdHR3zfGAbOr8bQVj/mlS9T4V48
aw1y+RyvwRYhvzXS6LQVffdvZ3OaQhe1g2F2NgBbQHF0UAr9YnOt7cTESX0SNjDJ
+UQwVFbgCfqT4OpXM+n4wdzBeyxubWr/jMnXiKZT6C3j9eC6xdZ1+4yOmP0RXYgu
GeGWOttlsdNFVGVGf9rHC6tWpCpWMSx8EZDy1qES7Tw=
`protect END_PROTECTED
