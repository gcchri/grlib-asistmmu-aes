`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NyvRo5OuvW/4XZvM3ttjN4Mu1RWgNhjhC8L5vafr0i2QiPRB6PkrKAdmsH8myIlo
reCJXsYISOlf7siuipag1kPB560y9Y6fgUIFBTJUmo8uvy3vbZ3CUHfuNZOYkHvN
jCIphTJQlLPIg5vYtKn5Lgk6sgd3YG4wsYRjwYbWwY0mLC0DgFIsiep0kmN24jBY
CrBzOY7mj7NW+jeE1mmxnji1Vw76B6UzqcaItCpvsoQK5ZfAXDuRAAApI+ZD+VC3
g4TVp2pD/ETCYJ+T/OSZ8sqXX8pn8ZqZMow2OWU8nT6PfNjTUc/WRh4rQ77lZbER
c9I+BIa/91UbfYna1Rtme2ekMilMQjeowecQZIyna3Ekx5VsxAOtec+HwKNlhA/L
k/VnDBMUd8BA6GrNlyOKEtnYDnH8i1FQWndByywl2iqGnwokxvayonjLyWREofEu
jca/CwTGbL1s1jJEVwZOruZuECBsf37wp02NCb7lslk=
`protect END_PROTECTED
