`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9rqnIMYCY7a+sYfodOX3YR1ZFJI2JVoI7crxF0FIM3AZg/FLCommwnLT9ns2Uxvi
YiIjep2OylttowmYxf7tjCgH5S9WcZvw5HYjS6WVxDnsYUuL9V6xuD89aa7c+bsi
Bd0EE5zO/er7PZJtMG+oU6o+Z576ZZJD/oNdCwUyT5DV4TppQjR9QBmU4R3PJWl9
slrvmnkY/c1+KNB5oRYQyCPJq9hDO3M/yMDOuxRy/fBL1dkIXZ6tpT275X0ftbuM
LLx+Toei5mU5OhK6af2fKbLsCLEGNLKqV9JSD8gr43pBkZRH461/Fxmh1QUyESm0
SAPYEmjNyXBiTEeLMLYUEDq7pVDVgCbi+raMqp28+wvoZXU+9WXXQQeAFVw+1vnP
Fsb9UjUetCOllzO8ywJlvYHqPhinJWsLrl1rTlDXWnCFKy94bL8iwy4oAuNJl9xV
lXGlPR/eQu0BnEX1tmxUXG4S0jDT4d2NQnz0FdfIrvlQLDC8xInmxFHDqp8s9O2r
lFPxHIgAGNQoiF0/tyYh7fahbuvIXwIyCXIaS6LxWcJYQ/+C1w3J+r47XmhYyd/S
SYuya4zd5OzD26sX/WQbN7Pc2+OTH0Ke76wr0WdJzxvX9Kc0LFzNL3lvCvJ6yWeO
vl5duYkdsvh6rVy/AOanhjLA8479UqNfUGKXF3BgqJ46Vol1uTi5GPa66mKsA/V8
0ZVE+S5omNJ3Zy3gWnjYrojSbN67sqo9odkaMFjHVIHZonW02wVRxqoRxYnUZesU
lQLVXsHhkczmXD8C+l8wDrViML36hPuOUTyK8GmXZtW0tO9WGCqz4siADuqCg53i
MYhdwFAXz+2pZvMqhUr3SHAxpxuVMp0yzRi7nZ6sylccV1Ow6rZONBmYS1PYAeRe
N3YGnGxFYhJEaB0r5quk8N2O6HKT8S4UgX/kVZ1mxPbkcyQVrz0VQqSTL+ljvEft
5lv6D6l+S+gpymY4z8BR6dPn6ssJIahM8cb9YWyWJAZtUV02fJBifP6nu+rAjWE4
g4kKRXAoekVXdv4LLgiAs59Ej1nPi1zLC7ThQ/+TFfTEMuy6TtDzaeJWdV9hY/AE
xjOpuF1A1M9s9FiILPEjl6B0xE+fcgWISoAEkqOJhMFRvSPV85Nk1706GR5ruHk2
fTwhPrR8WU3oXIiT6GRuKG1dweufpHimNgW+STX+MCZoHB2LVmJKOw9ukI98GqAr
dk4iE5TXq/9roBV0hY7goLjbjwYNiSvYIy+5q1sI8MtQJTXPEuJBhvThPnrU4Tgv
9I/UZegrJLWuo3f+ThJcRugSokCIZuIDhKDKvbHlLmp4q0o5+HuDJjcBkcJQRect
QWX+E0diHiYS5p40Qrhp0QJax9+vLmkdvISFK09zRJ9d67P26IiWL09kmR8dALS+
ZLz2DREROqsR6v/TfeDL082UHNdCSPkbL/o4Vpp4VZUN/5+zUjiT1xARFfbIJTpd
/arxj+HHH/O9+//F/6xnAGu0UCekgdN8BVw5sBjWNU74TWnJDMTSdLnnBROz0i5p
DiJulFIg1FRFFBKLRcfjTMnJWi25Nhm6HSigd4fsosE6gKgxRaswJ13zyitcZB2c
VDys16ZDYMtcunHqpwgAqPo/HdeugmHQdpbdawraYdzmZJqZzLYFGWc3Y/kmHT10
IvSEFA7DQ0iJxvHMjDz7Vy9l25Um8ZAyDXO5ONHSMLGEDZpZ2q3VqzMKn1eXq0EH
THDkZQteX6Zhu6vZPqR8/ju+zQ1yqnbQeJ3J8JsIisuYgcoTXpA5WIxlkTfVeynD
l/KgRvMt3RAwHUVu1GUBJR4EHHQZl6n7XHDe2T9w+dRxi/3vHFCQeDDqg3eXFXC7
zobigziJeWh2ZTzqU+K3wRs5Urpo1eYiJXQ5K1uLIc6pyxvNDtRgogs3TuU5huxm
PFCD7PMqxs4eO+zUbkqEklX6tMq4r0Uldeg9dbFYquaLl3NbGKI5Y7KZTW2WrCiV
MRmlO+2JUwNWF6oskG32NfBaRtcSGWgIqPsKxwxA8LtzdP94DSvuNX/91NUW6gAf
sRozgsDEjTDg8uNuvsROuvk4+LcvREZpJ5o4cYQnA6idNnbzaHTDZOs6ufPgAhOP
Y79tlbsLTFZqvwq6jZFDr88Uas5w9YBJCUmM7z65wVLKIbW5AGBE8zmzdN97FUQv
aEDAlDnS4hBWWTozHd8vXEd1tFDqUk1Wl7ILZfK683cQq+iP1IZBild0TYHSggpL
NraOFXR1ahFMgEM3fbprXcHwvgqfLv8FyB/N1U2O7CSNBVTF0Kjzj3ORZzo5++r/
ChPuavyJrw2HhF2BM3f6ERZzISN+pdYCKLoTyx//HtUxaACLzVYQ3AXNRvJA9Fx+
0x39wZUXLkOIKh06dQShHyA6f7mNSqHiaYq8clej6yvNdLYyi0nWtAzIAUskErNq
P+fyRxLNUiviwlUZE8Xjol/07cKhDVUg8erJsVmYmAhSPf3aXFiiD/7yQVGifXcx
stTDxfTftrWUpnAMn/NAhL3aT51wVyPIYp5M/KPTCGd2L6VssuSnBOG4QX1sJGqF
urDOodKp781Noq+7TC2wPyAp9d053J4Od8E8JofMIIspC6NmHAvoTYBtzucmNnn0
`protect END_PROTECTED
