`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCN36gsmT2IoevdJmgVC/kSes+0cTW41w/C3VHRLw9juxikYkahVVdOfcIuBDy9W
fu2qqGw6p4L2f/rTxvhzmsUtaqvOAG6a77lklCl2msiCqQpigo+rCDLF456XhcVC
hnqG7ZshZX3wXCBX5z0Cp1xsTWMPxLOquXReui9ymwh0xBehG0ZzlLt+0/FBitoh
Hqv9PbSu9SGz9dTaB9S97eMjd6ndUQ7rhkpBPHuZ90r37ok8g+PZ0rA6ErrQaK7p
W6cB25Bkw/6e78+PttBBfJLqv/zny3m1jo2RZx8s7v47crIzswxVIdYHCLXXYWnb
NaN0NZTF8AJA78rUR8UfytX9xV8k2e/4frt+hOEBp6lc/aeZsExwaGjr3HJlfMcm
alwDgq5s2YBX1zQKvJJU2hM+JKiDiZ5vnPCo1YvomZ4eoR1i+f0mgMBSngCvk5Gb
z25K8ZBv+n+3daYCoWbrSfz0Q43y1CAqpSQ2Bf12S2tvCum96oO1n3inp10L4N+J
QZcl9xkUcpa1Fh7blH25Juc/ulbOV3r8dSBQK2eRzRcopckYIoptXNsnckbIQzhA
lxqBtI14FN7T/LSdcVK7wuoUbJQtegZpRvlCbVD2Z7CPX1G+dT6ccB7DbPJjskVR
9XSF7oXYNPIwX2kMZryooxZ144Grm6xYMS4FnMKKghM7MLDqrOmMFi+x6H9tbu3q
icP53NecyNJjII97obbB2ig/+pzZMr2KhwnpORCy6dhSQt5pSTCkDUPvoYq5WfzN
i9euZFlsQ6db3RO2FVNKw1YDr29SZnZ6sOmO5sqdyFUte4j9EPdDv3UeUfGz9SZP
QTXWo/+3+z5wR6HMYVS0xpCXypmMIlQjklV3f/1SdmAfbDx94MqaoZFNiODg5nrN
XUi5AQDady2ybIuivWvwraF7Q030xkaN8MS0YI0DauU=
`protect END_PROTECTED
