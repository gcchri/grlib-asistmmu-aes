`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8QSjsBzDFI2RIhBEdidvMMK9no9pw5XKITcl6wrtNSMbsSPiNeJhNZcuP50aHW7J
z9rno7Yjy+fAO6j66IfbxoiEClVojVWuSQms0B89Bag/KJhM+tTRNmlfIGSCkkdL
j+6oEBEPuvx09OXEs9cQzUZkMhJE8+he0MPHr8HHUbDkMvN3zDf7XwsI3P5KnzqB
yTD1YaMdf0qQQNg5MXODfG5bd+NVstQ66m8F1uLB53YhsE6KyDGfVh0TzEVbKiWa
D2qmeiA04PpAWAQW3jQn3IeEFs+IMqw3YPB53PSo6fdv6kwUv7d+8B2C7kwcR/S8
Gjd2J9w9hQgIbZklDOICBJJVAzcEtXgxOGpJeyHGVGTCT6tXOhGkeXij6pqTS9qz
r9wOqY8dEe2H7MsfizQ8Z3Kna5U/hubYQcOWeMPJhpZ3pO0Op7SY8HdttyosmVqJ
RKRp6mVUkkbqQp3sdYXpC9T/knyQpgNPJgMzfa5MOxPi3pJ6wQhB6XklzLZAuAyP
SBqxh6FkibtkZCLpSBYFkRbV9UZziQorvonxRziZL7HoVQ9ugVXmrVJy8XtPj2FJ
nWR2lABqm7x+ZQvbLuj8520KdiSCZEOJ9nSsakJHkcUcfWfBBuHyfQ2kTl/1BN0Z
KqDyMste2Xyv6LZl6PZzC2RxbgyBpkMAns4bWOFcKvgC9+MRefcV+YeLT4wJKOeL
1dnbI2+/K/TLw/HbYKOdO6mM0CamKQFvhYyTr9IsYqKtBWrRomlj4D4IXx00X9Jf
HYBFsAVCSWyeJNeCz77c4tw0AoflOoRSAeDr/QD7W660YyZt7LvnAJYhc5kq7kR9
94/df+DbUawhPI4qJ3/m1k13wHTc+c361Anv8hBxcstLJ+KGlhPhvJ8zixi8Mc9X
38NhdLpL58JvGWfi+95KajaYpUDLaQc0FoM25uEH5d6EYiRtCgCiJDLJ5iqtFkHf
saDgh1baKyGCyoHTIG8GfcT4vLKNTvHq4PthnIUu6UOzt3+pNDTiLTb0jJDXp0lt
fV7CdUgk2XxkIbclcdi5KpPnMky3MDT4vdAKAON7j1v6NhC3KVdQ1/VwqWlYRhvC
utecTj7ec1r4g5x6E8EaYOVfBi/NT6AZE+m82RYF33/OYs1UREJofVbKrGkKoLU5
xL9z/LVxrCmh2V13iWEHaukHm9zxFZ4BB9qhvxQOT0YAgfeW3eNCbMsOFKCsSfHw
3+9tC4Zdt/HBGS4AdgZHc96Pe+zY5MvC+K3g9ortaejDdvE4kBznyoBIJhkVhkYD
YUU288wY8UF1IBxefAWZKsi7xIrcMXaL5N1U0gRcRIY8+v4LnPkN9gyHw3WUOm7i
UXCV7N/e/cpvxX/osPWhBp7rrFW48l0M314hiBVuHuEh3PseyuHH++9Mfm0xWQE0
p+Jh6YhX7CwA3r3WN8+TJYkS5XUI2dKKpITkHmxWQoDoCeQUGthXpYpjABA0qtj5
ofi/bhTyQ+HZumYx6VjEq0obiJhEnXu3bHGwWI/xUsyLv8We273MxKO3clJOSmuA
o5W2TycKyoXEh0F8H+1x8m3UEdWm5R+lzJ4Kr+Kqvfw=
`protect END_PROTECTED
