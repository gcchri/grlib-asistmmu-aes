`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nnKMh9lyDvb64ovXlwhPgKFiUfr36R29h6w8WyW1yPeOqarAy4DYndbwnOc5AFnq
5NOT2sqB8PENZ9AY9LCln1beISOXEwv6TlQAQUlL7VhqsVICBIxWxrgpL6BDcSL0
BHDCC7GlT+viW9IbW2RV+clHZsnCSVzhyQ84TMEdUCD2owfP4myGVjxBDXo63jxs
BkU+E8xyxQOJwP5iiEgi3bn+xKR3OqPSxWHbhEq0LfuI7HUEdvcvxSgzZHaUKYZG
EOkjdsUWszIwx+LpL+sTd/KMO8fh3UYHGGiRIG7fbqO176toYuDXxRV3mwTS4oSn
T5u7327FVxfuaFBL87asuadQegnxaJKWJTJZtvj6rCgSobRK8Ps7cR7QCwHh7feb
X9KwGulV2Zl8uOL3pNrd7UdbCqfuS0l4+xZ6XJHB32AcdzEqUAJxorOLKY9JypfJ
izv4JFWnekDBUu0Wx0+S42Ldt0iAS0Qud+DuwZ5AgeqClPEb2JgK/xZhL7WAOgY9
8QUkzCiM5W8kakhW4lAZdg1ewXKHUkbsBNGenB1u3Q7eR6PE0/I89rxoTjxyuaYI
GhiwSU95nfx8S4SvTmrS5ahiAghGe95oBffoddqCtPQ=
`protect END_PROTECTED
