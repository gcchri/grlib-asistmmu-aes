`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5iUF7/U7Ysj2OLgIQrMbK5KMP73JuWmKco2oL76Kki7yrydo4cGdN4jfsZO1g0w
BYUeJjEZiQejGAD/gC5rVeOjNPAJP8S5wgJzXytGIyS/FuAuDtrPRe0hs0lEmgtD
Pr/i5FZxUUai+L3nFqh0PRk2KDf9t5zeEf2e1FSJFA/wcRMAYEvNcnsva/0yLkr/
2haJq/u7bXQkseAZNylL5DgJk+i/3tCMiRSRcrlns0WDsms66kMQnzaftAsHRhUq
G7UDn/1HWks653gj+/jG+4ktvioJexDoTGuuyDF6ok2yNn2RduOm1CTZAkHfdilw
bmbKV50p1vziaASfbMAftg==
`protect END_PROTECTED
