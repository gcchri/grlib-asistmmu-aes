`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wp1YBsvvDz+WEVsmEkFE6pojYdu4db1SvyyXIMEL05JfwbSKl8WHfZaFJsmKwuib
Y6Q2eF8g5VoTf/CNRRI/d8bR60FNPNn3nWbcDlfymjYsa4eiMJeo0BLh90Pi2v5P
tDDfMZR3es6LjoRdPWLGFunijWyKSj3OgDGO7NulXIexmPbfvSe+ib+JvNH/i+MK
he4gOkpvI7ootLz7chgKJuTgREwloKHCk8KCHTAH74ZjsIx/XDSHXG/zlVdP/pEb
RYquJs1gRGQg9INmHXNCqhFtx2cmaG/ZvYpwlYXyAsLCzb87Pxm5IlTUnpg52nRP
6QfCIHYJD+RzuSF16wFLTQ==
`protect END_PROTECTED
