`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EPUwkQGRv6A2LoLkFlHoe2C5/5nTuBIrzcNc3nOn7iNFBKn4GX1RDFcgV4q/F5xi
ttwLhowvSRviMtbDAESHaJbQuHy/poqY/90jrwHT8Cr6nfVgZ4cUyifFOoALSpsg
IWfbrUcm0RvfNo3o8epCvOyQn3vCnCMlFOZ/9K7X9a90KLJlCwVMgNkzXeZZyVct
/jm5dcKvM845ouOtCPOjjznwVdY0aduNM84r+LFM+GXusEFJnJMR0xb7rbs3s35J
mirIST1fijl1KRd9S25rxQ==
`protect END_PROTECTED
