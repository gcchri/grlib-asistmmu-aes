`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fyRUi8gDdS+NvIeC597GZRGEF+WEzLNoGuinBZ2cvqFafDPlBDdN1jas2jWhfFuY
H5gCmw/FnxtTOjbQ4I+LU/UQ9Q1l9vwqkqe34AWq9FLnrpX7vGq/4RmWnoHSOnN+
iTpRWhGKKxubN6D/BBM/vI3cMyjdfSnUHeekqK4QUA1343Ply6oPnDPwNg5Yu439
g5sAJ3rqJ2HG4lTarKyVaR8/ngVD0z4HrvkIKPooHGfSp86qeWKszItkUS8bj2dm
C2aRoEU2MON8psXkbcYSwIjJV+akfPuOWgyUytnaGEQFn9SOWtAqeoBdnfrrPgHJ
NT4uz+ZXXQgONriAhF43QOg40VlxUB6sinxDdgjZfb1qGquWLZkPOCy4VV/JwHUU
X/l0FND93yjm9UG/uHnXxV59U3q116n1/o4q39vwJmtl7n6X5EflFFdvMMqnJxhX
68Tu31rA9HF0N3JNCWMEru40Pmp6Ck1Wpf0zzKNGmaIZvnSsF3Zw9iUw3L3n2+Bh
`protect END_PROTECTED
