`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeyL3K3LoQULOBYiw8WHOY1l1rSrlHBPbHd/0Fv8PuamUfwsDm8eyneG07plDtyQ
4oVDCfADvbhVoZhYKKM0tQRb7hmtIFPoDXL2B5M5A70GEmIimM6isIfgf/8F89qN
vRR+IwR92JFsxjLVQ8CvobihkR+/WwjJUPM5d3+oSkUx+07c6/pbQ6DRUaL4lBjD
Hc+rdS1EI7L/jb+aOo1c1a/nL5w4JA95rUehVIq48yhKwc6UEFdo38UpxO87u0kD
mccBFIf282IY/AIM6lAWFI0/HuV9mGHr0MrXpo7yXM2ND0+YQGEyDGycktbJsZU3
ahoh2Pk/uE9MlyScQ2wWew==
`protect END_PROTECTED
