`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bFDHedxoHnF4Tf4rzZ6Jd28sGlDMlIS3giO07DozhWdJ1xF9aBawXdN41U71wV+4
dEX/Gr5SsG3Km3xjUCg5hsz1JW4W1YXSkDFTf7DBdtZUhSh7UQby6AVe+EczhSQt
tiIiVAok92/QPtnv9MIpTM/xwrEl2xnxEv7UoYSK6A8bPjXooT5WS7gB2V90LaP1
tjOnUFhmPGWCQNG7RAw/A4GHbRErqm09CWbrP+FzgyCSQPEEgANqjDUInWzcVp1n
vWmJ5az5GyFnmnMOs5M9DkpELHXzooe7E42xRyIogpJtVsvDTYTV9EqtG5MGlNqN
dFSiFWTubuTziuhEnmOuDNXRG6ziSoNuEXFl4X5wKoUa86yV00GMBurXWI+5pdzt
m2N694p6RzWgD3ZjceB+WQpqYQcbRrSMva5qszaJJ1Ryhfz+Xs25LkT+GN9sUnPq
Stgh2ugDScunpUHXDqdX9eEw98CW3dHQyh+ZRFBocBU1hsPwyfef2PpqjQKd7VGk
X2n8ApiPdxWzY4VwL8O5+J8uxkh9nkFKm+q8K10Mdw76lv+0dARD9rP7d3+1eZT2
dPrg1EmW6S2I5qRcKopHtGiEcEUtC/xgMPAUjbQ42mSQRTI8QFcfO0pYQQljIuX3
af7lxe+DvtHNIG8pHAIGEO/alPmFXcT7WAQ3dhTjye7QBpbP16S6W1t5Fnubqz7W
Sz5yOePeL3/cyvMm29FOnfZX3g0258dQ3hSnwsB29jmq/DZGu1HP7LvbQuE8W1hJ
Y4jgj5V2w/Si4Ir8j9NjivhFphqRqmXpwQz9MsN6I670Hjvyzhm37MQ/zkgLIFku
AjvLhL2XVzy+Tgu54H/LOW80CCHVMzga2xEIdDU2yHR7GBbSBL+BrPma19gV9/vb
9qYYMGbwoCSStXxikVJYgyZ49rdb/coScyDIUtvLmSIYsaFndd+HSNuLDsO4Jccz
e4Mor1AlLDGP18QvUdiw11FnOm2w9QxDltT3IYeyzrGFH98cz7VT4n00ExjESUk5
xEWiXFQxtRAxVuzn7RR7SxE4weroRltyLjHLN3gH/zfyAQQ4Unx2UvGBWKGJAJNW
xZ+oBpgLC5OEe9lsnl5oPPeUsbmNhb4R+szWXG1SDOwosZPK8AYfJ8VZ6su2B83w
dl/nGR8VZCZCmQHrZzUWPQMsZHEjq5ryWeUxsTghEDmQXGJLjKh18JoST/r4y9WF
1j0geOR9ZRZN9y914F7jJ0hDjH2OEg4QSX0rb+rPnIjItdOko120GbsKNZBif8jX
a8nTl1xdEzHk0yA8BqRmkzsueGd7pNAaR5i5TqwQRmI3a5aUXC/GfXaWocpL+shZ
3hhCU0Qc4Lc1v8fKz3l/mZQqTbap2d8Toq0GVQ16hR318mrM4pao425i2O4r2Vh/
cqDwOkyRtlzj5y667Vc6RTTxLnlTktT8yymH7u1ILykR7/cTwxsWO1wI8O+/Hyb2
o0af3sb062EQ00KHH033QOGMhTnNGP6vvV8zrbFArE1rB0/UATuxG/6fLA/b4XxL
sLFDw1Q93lvjFQVaQVrflg==
`protect END_PROTECTED
