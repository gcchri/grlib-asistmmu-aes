`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RIrZPI7gIpZ73EF7osBOalElOs96cuhDChqQPHABP4bj2DzVURYoaf1unlYf5dPC
g9DB+4/KEoRk7m4n/vrg6ngVbOcJ0FVcvO2XKitxyoLzbp4Vsf1Or4/2kXrziGWF
npZNjjoQc1lW8S/HzIM9L7g6NvV+Aey04cxJrK+e6bwcsObZh7DoFhEeAEr3ok0E
YqJkjkhPljY+BkZgM9CgoH+RFOw0Y2PV38ms1Rt2bilw+lHvjHWRFSfaaJ/Xf3dV
2/7JseCod3vLykSIko6hZO15I0QH/l1GWy2blm31Cy/tIM++GZBTeV0yK4L266NV
kqLWO5QRAE6jAc9zL8/JmYttI/BI3uO1Sb5s0hVrnP/XsC3yQi3TFBvGKmqO/OCe
7G1LCsmRa6q5yXr/Cxleew==
`protect END_PROTECTED
