`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PU1EjLRdUPcfd5qDtIBi/vNgZmNdsrT2PP4s18padwyQGFjK0jWVEcr1KFY7M9Wl
2sk0Gm5S4FnKOnaEJvECUIuw6JsiBAZ6cqEi4v50Qi8kIcWWI7Q2euafLfR212nB
5yzNXylQZLA9rFXd/rkWwZ2f+HRqmy41YR+yqqg97N/nv0RFQyq66fD8aqE+ytd8
CfxH1R8ZTY7eWahoMQAb+6hfZZhgXsh7h2lzU9SD0D+BfRPo4tjGelYseg6aWirN
mvwSJL/VUXp/REiXNKC0Vz4jHO9ZOZ/PAZLMW/vGiykw18lYJjwYc1V6G7HLvDFU
ZbT6PE44MwAdeLzZ0/9J3WTLmmoQ5XeDvVEx2l0bDUIx179pYkg5kdGaZOYSK1Zr
SUyf3K0mU7XQ8Ddb7P0tks7+DIKcxFnJZvpiiocYvqufIlNVGgGFqh26CgzesSmg
/4fM7/X6cl8sA2Pg76aqhhiZtdI1eMJPc90+hYeIWJmPFOS+2CzmJ2r23PU+1x8P
`protect END_PROTECTED
