`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JfYIQPdS6sRaqK95eBXYkD2Rft6ZfjxfXSA70VKUeVDbjjNzVXzchM1fK90sk39w
AOeTmCiFjd30KzfKUeMoGW0JuAu+EXpL2iYe/+mUQ6nnvyqywQ62VEgDutFlf8Ge
2fJZGFZCkt8F+N9nHtIER/uUPhn6JZpjhdOaoQohl+ZYGhv5cXn07AN6XURy/aq4
U9CDAjUNaHYsy59IQc3EPy6N7zzi9BkoKYgPaAoeu1+ZC06AxQu+9D16PbtXV68w
EJiB2C07G7+v4L2rF3mM/75UZ/h2/r2AOwttYE2PV53Mp7cHCAaeKtPnE+itD16z
3WUXb24mNHsPo8waJgYPeg==
`protect END_PROTECTED
