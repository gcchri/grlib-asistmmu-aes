`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ak1GWL2ckkUm2zyS7B5/Vv3T+fr98JzsNkhEACruYPR/0bf/PtdXHkYiYMR9XxVG
ZWotgkdD8/WhNpRcUT2JNE/oJIaA3zB9gjkoEroECuC0k3ccxzwYGA0+VSLuc9gj
MGzI76HzZaFqS6+AfBLpknndAu5LPg7djWmDIKKHad8I8qN1uRzpbeR80hOQgAFP
NFPXS4m0HBkoZ8Hun+mrLFJUBUWDNxnN3zhkyFX+zZPX4UqUmwrpU/wW+QR9BmLC
fCWn58mc3PFYf8M61y10n/k5haTk7BdeFFPS8mEVT9bQw7GGlgjejR8lOFZmqeQV
NFBebf8hV0JS3D8IB3+Tj2NxHCPqHhgCmxjitWUXVyTHZ8xZs4FiFzVB1md9sbxp
lcQd62iVENeis05Ll2St7zUL3XdaznWzNWHeO0eVvPq1WUPEWjDFAmh8KBwJf6sx
0USfcwVLyOtjd9J1ABSsjbVgG0H62zwuaZkmFJLnuRfWAfKqmXrKJ3ADfaNB/Zce
i/v/YfBkNCmzigW/CWdtrKC3zmpD76bp+GwNCSmjXOkmj/xTxW3p4FXTsW9BBapg
9eq8NEUPte8hj036U98EjbrII4+P6fD65XzB3CFP4bKur6eFYdmcVltldMRojl2k
bjt9Kjq/+xXWGsB9tGeD+n00JQ4+vWmFkA6DiGNGgkIFSvJ4OvKNTSQ8DTfvJdfH
IRPD7RSX02y/Edrc5R06GKf5vdu+uegXyuKa5j9ao3sPLHgPUYV1g7irR4X/VOqD
SqIh1ZXbn3hgx5SgoAgEjUHsMgj6SoV3/kXx7zhfThrerJa0HdKtgRkn0bT4Yw7I
WX/e/DD8/6yrh6dtUS8okN8UMnKhKjic9ClOl4LYDR5WWBNtujC15RBddTsLUh5Z
YFlLzYwM+NSqx5jp2nKKcpH0hRbsIjw6c0mMKHEyheNI8llA1pduNp/YUtdreyye
T8xM5TxXkNvYQYxgyAKku4EhkxaCZuwI40MW6DiTXVHKAMblg1yeA7wToPohmtml
4XQK5Egy3qJofpgY3BMyYk8NJSFpq4jzIYLveYke6kMwo1hOq9oUzCHNyuVYVc7G
S235NlkmoyNS1ov5Ev59yFRetuYpg+FEco/EfqN2VnJpT0UK1bhcqBz8iUCNlGVD
yUgsdPziX/NQvD3QRjE9f9JEToo1/Py0fz+yGKkyQJbFSZoScDIrXIC9iUdttNCb
mxQHRU5EBwDuYjHDzvOi+QrJpL0/d0nqAm7nBg3ALN75CXliPWXaCI6Rr3ZW0LAP
tDheS36TjQQae4t3NvlvCO4rTh+9VYdWDMARr8fTWuLS/nOpkuq+94qBBi4e+Bb9
/tQYldymcf6E45UnDT3H/5oPB9TYq/3aU6Y2lmMJzo6CZARXyynpQPmpwHR/igoM
iggmgbK/gP4ksqCq2g/kRAcM3/k9P78TA1HPYdp8xFQeSF6xgbKTpbs/C/IPyF6J
da/oax9SgQudgZnY6LjT16RioNektDDUJZClqMQxUThysZm4VW1vDAtf2ZWC5u6C
Qp+fY/VjspAiIrIgcds1nBpGjz1CKRNahdw3cIbxdiLbaR7SsgNt29AGTYlicn3Y
JuyCoUJi8FJ0HeiMLKEUmJnnSB7QSTZ3QYxhAel0axjQsSnDOqXO35bc7AkCzgW/
8wwk/L+gScbzm+HR7pwDm6IwRXfNDYJwPKjsh+p5CEOQ6A/dX24GtrMyD1hO51qy
ADZXiCrmlvucfDvYiVoLqlcFxXhmGPW37qGqna6nsXbE94TIJdd7OJCn7aF6qAy8
dPJiM2FZ7ajAeatmEt5M79hlRjvwXM96KZe2eT52ux1+1qAm07ZJo3cl2vlJoVsb
l47kIqRsge6iQSwbhy4nI2zouSvgVLly9yhRZ6ur4ls6t2AZ9vgCgTqlzrjGSbni
`protect END_PROTECTED
