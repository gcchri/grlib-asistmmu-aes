`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jiMqpUD2F5Qq98GzzVRYRR1u9B8F2I7TOJy4Cq4MdT7iwifm1/tbmcE2u4VibTD
lmE0rCCID0lpkNB4Rs5962rAnWX8XsVTS0/RleQecT/N6EFeuNTUBe7nis1uf/An
FbzgbeXHhY7JIssQU0sDUF4GtyQEdpdSmWP1RvlZVhWTHraOzfUxM4i7hF7WMmN/
GVQNZ74Vt4Dj6ym1AOacC6ld6gKfUk/u7p962o8KoBYPxm5+FYdy+bF0qbDjS+Ea
fm9OffZfx+kcQBTve63ZYvnI8U5hkYYAsqjZRcTU9iQqgclyhNI5agTT61KqMfem
ADlR5q3ibvpruJo3R66WxJRkoSI5m6Qffza3OodP6XC0YeCNz66gbSSu66H0R6hs
HseJPI3w5YHg0xEQSEk0A1WR1hPQlC4oWFzPdMVCfMIZzgaVLum+NcEknSVkxVG3
B0+G44gcfPIbKt3QQ25ApcakESf5T9YO4FkDrG9KSIEHfv8aCpZR9sO32MuggrxS
qWzrAvKdTo7BPFptJRrhJoMlMng69Dq7P5eJhrorBQQWvYbZIedDGLgRpyjiSZVp
38D2nxfPuZiF0aAVJaLEzzFX8o+CzJpaKoxtzXgNW9oBp6bLN5lrrm9ohGsyqMIm
GuISZzBVJsOVqfhxmmeCrMZnaA5u6d71KGc1ffTHmhK7N7hyldh0xkBwP7AFmwWo
`protect END_PROTECTED
