`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDTUU9RaJPiVzu90AnGnYfNfaPlGut/LPeBtbPx8kwecOCyrsbbEcwnFfRkWeTyc
GYfPrvYjedOxffdNU41akKlkYVSI+pCiW2T7rvSWLTWjysHKuECCHvmTZWKy4gFc
q/p8j3ewygJTB7MP+ZKNrFF4BnuYpFjp4FUym1ps1s9unh8F6RtdWHD7m6HJxo3w
b1nDGchBxBsmTOF0jNkXEJ5kbdYbEkajRcevbtSSB0CJ8+36PXyDevnxWIJ2fTkq
m8Lq+QHBDmgF9IbS1P47UQ==
`protect END_PROTECTED
