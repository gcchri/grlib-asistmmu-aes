`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z3sFF7X6UP3XXQVnBx4FS9iRMc4crbSVjtMoBaUXkHqnE1Qv9Mw7bHqlgmVd9oGR
bCTKZKdXFLSaC6EJpzLc9fEsTl/xGI6juEXPZMjHdD6/1248MekGvOJ5r20IfqCW
0pKKmK4FELkkyCN2+bkMSm8LSYFyf6SNVBq5CsUOq8KZVWiikGde5CzqQlBiAZFP
pTnKBEnWY9TFBTlG65I87c1RxwXITSVTUh+Noq5Fp95jsFMY9/cddmfqVrUYbybg
cd/eSDoAOmQnyVDp04FizQ==
`protect END_PROTECTED
