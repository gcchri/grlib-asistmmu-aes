`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6wkKJL4kM1uhfoJ/4Ap1p69GZf4l6QaYMCe90vy22zgc/tbTdh5fUjrXyt7LrLhv
7XwGqcFyp1JgDjUJolaIuYVGGvUfvWRS3geR25Cp0q49Z1CxKYKojJWSbtxhVCms
PHt6rfo5+1CECrC4TIb8uXid+wetxCEfP/G1zgPb5HnvsfVWNq4ZdlSmICs/nWFw
xfgK2z7Q4uBYWKUwOSHcXdEb7d4gw+B2orirQI8N8DFx4yTtqApK0aeRnuW/YkHj
HMkt01Hq61RpzU4BtQDZgkNRSpNdmQlPyIArc5lOVvRGiTeBckvEohHOGmmBagl6
9buCcjvfAg2VUrTMlOHvdQ8Hxiu43uODiRehQOGJMJyix2PjN+ImKwLFhvHwIIeE
cASdfH/aGWJdeb5zrrC7CwadLJCdXskS8XQdJ/gsqYhqJfrVD5k/ILHpPv06s7Xd
`protect END_PROTECTED
