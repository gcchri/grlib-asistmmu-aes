`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZYLFE7J29/T/HsSIjxWgnq43xW9jKGbk+Vi8npby8ydX3ernJtTtRcI2paNAQt+3
buTKuKACApflcPRnulTXYTHmVx06GWjsRFA80xO4G5bfyI7eRkT6lvvJxP0B+PzW
AyF1CcigCzltYrebPKFuncwGehk9kI0mlfqqpAlqG4/hQQgd49peba2SNT27gJ6U
qHXx9gTwMywi3Z73x0dacBM/CSQzN4WLvS0f6+8DxXv/vL0ZpGp9HF+qYGziLpF7
qkmyIQh5CGCUtOnCzrWuBa6DbmCx3CZM4b7/qxWg1QHETxcZP3eWPE1ieDq8smh5
KhV30TmUTk26OYOH/t/qLX3bXmbYQS2beIVyhMZfxlIbxL084IBS2dUe+scTqgKl
aj6I/gynYOjfoueR2mZTAgSxcdwfljBDEUttZoLMmy873H9OU9VIqVGw1+80Hjk0
w2B27cEJrZc5nuHZfqyjYaX3YWZtsLsC7uBgSlIHkeKbu8J18CxeW50weYZ0knYR
y/C+aNhBmNx/rkJP+eSDejACAwvt7z5Gzd/JgEnO40o=
`protect END_PROTECTED
