`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79FTHZ0vklW1xLb/WTD+Zvy1B3F7CxmjEX41iI4paZ0oHFTKow0MBUX1MbiU75fb
7+DxnGnWJFsAicqp0/j9e71Ty5+RTB/9ftQv/uRWpZvUKGe/dmZRNghCGtSSgpva
D3s2fUg3MhlBKZOR1E09+VEDe4C5k/7vcXux6/gjUcQ5vqzSUtO3gKuVRYkBd+Na
/JuC+7hPFp4NeyXRjxf7L3ULnMHlFuLPJcGP/eX7dZggIjEDiCCVBmTzUaBcTuhO
Fe2391ze5Fy3tT8yS1uE6LqktzvNXLhIHYsZPkvRjr1HWkA8be9fmwfQGcgQDMmG
Lnrp7f+nTMNBGGl6su5zDg==
`protect END_PROTECTED
