`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/CDYkPKePBV+R2E1xXMj0/OWRCfD8WJ9kir06t4vZg5aNvnYVVxSmzpI5Tro+0m
MBVjWfxbLqaxdlM8J+Q2yUny2fOaUdq4GmVroVsJ2t9yRQm5df5b8U53rVs26jS4
sru7k1swXHC4fAnIhjVYNk7jL1rH3VpYODJwUilan9GXqHBz0+ZnUcMLZctAC7de
5wY0aVK7n086X0Q2QFxPBU9k2Ev/voJ9N9RfeAllYClSQYMeYk35v/UxOfgFgc+W
GFSfhr/xQf0dnv/hy+SPIEG2wdsJx0Sf2JcLblsGHPHmlUdeC2gIShGnzaRkr65U
Kr9iOckSaxnypwq05dn645g1CpX3lfvhlk5QQSvYdRaCEGrvOSgm9SW/rZZxHB1N
dKY2BNvu+frrVM+zY7Fi7g==
`protect END_PROTECTED
