`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nw0yJHHaz6dJw8YeqEJtU0cfuTkWbU06bnoOoKoON9MBj6pe7/MXbmKtHbfIRGGQ
PC0BFcoGybBCnVH3RbvY7UdoNL+YOxADpiralc5Y7801ad1DooYLSdBv5jFkz/VD
/dTRV0X7OS8XCvj2NoofYQ+Ckx5zwjFve915u5Uf02h/Ysj0AIaMcR0h1DVp1kS0
k+KO8Fq6JwkOlKLB2w40NVrX1O3k6GyrOmqR4zUcvcg1fCwRuftIBZ/obLOyKbhx
R46dcl2BMaE6zbq6bPv3nF1TMcnxyHJKDX7vFL3hUvRdT78nrLhxSUI/3GoRa+l9
0Qo997Zg3w6PmFd6s2hUbd1KgOSkLtGHL3bsVdtGQAr4gxaZhDdq95w+XbBpCRay
mEIduavoFVPYti+YYoLAxWwZXoLhwdoYkDEtG+BAAnlFVkL9zitStJisM55SzhHs
yfk/scQaLhYT4aGuex97JMYLjG6LLPE1Vk7g7R4IInkN4w4I9eVRZ1BXABjWSvo/
6Q29FWyV8U5lF+85WXm/SrSJbp+BZLaS9eE/X3PES7gkVUM8CDiI/uEAKG7imVI/
pSpdq470RD65QzNQxoH7/jcGgV86paFpQTgtQdI468bfmFmmEmTLPK/rmH7F4FJs
jwAkeRa5fvvk2MIjXtGW71x5OqPPvmG6cWZJllLR53eukZ0i8wJib/F/1gVWsVSU
978FYgaBnh1viwjyLOVshEMDp5hmPNMzSXBrJw0AVKjUMbmGiC/7vItOz4QUejAm
n9qkWba6X+0w5i13yjtCLGreO96QgXGM0XGgCzCkkQKcsTvbqADmKh2xjuTkfo6T
c4WzD3ajK/Tq7qP5UpOCYg==
`protect END_PROTECTED
