`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9oe1X/nfGKgf/x96FuT4q2imXWEHWlKWDGMLaS5J/gfx5RuePHHSwMD1mDF759i
3VrCiq3z9djJUWOD27jcHNA9/fTPM7fFrUlASud0qHFwoZQL9aB6AojfGv99ymKT
ZSkWGkVgaOqiWYZLUUc/bMC7HzDWHTaw5KAW6FX7g9NCSIAGf7SdiinJ8Bgx2ZFb
2CAgx7zuQt8WBT93fYtzVEtYFvZSD3MZK7z0x5huf0yt0GEH7H70jbA4OhxeJGSk
dEJk/c3rCDEh6r/J9xDzk3/kAVqSTfCA47TaOf7PG7W58XREGjHbXnZQp22C/cEU
ys6dkshYl/9xdndh0Qn+HGpqREvjC/aQle/JK65XAlZ9Wakjo6il2MS7k2PLVDWz
Wri0T56snRqplAcv3NZfv3OmhnlHXeHBQC1VNB5PTJfBqZgqfvyVJqUzYBZbHEaa
jerdKJZgZFsVYxH8ZB+t3fF0cc/KQ1Sph7XQ/u2aspZQRvysDo8KUU95YO1aYpv2
guDzE8mEI0nFIhBV62fsPm16ZmLGCzQyOAylsi+Ox1Y358PXd6s9jt5j/xwr+CO9
09myYGe9aMj8X6iWBMmLupY/jJRwn9E9DKPolv8tFZWAF6pfD9q578tIwzpMiQel
cjHw6rLlvvqkaNgO43V71Q==
`protect END_PROTECTED
