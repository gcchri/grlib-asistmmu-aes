`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mDGXSgSkfLKteEnatTt2yaJ+rrhYJJVKV4fNkQNa1besW2/uLBusujH80Bms5hTn
WNSXYwkF/KIJk+d+WIe1F90fjBP44VnRDiUL6JS2yS80Dw/t2ZkuPYCkXNVIxV3r
Y6aqbsoQREaz92hrSt3qOZKlv5ziga8+P1/0HDVMb3prgPRP7MgDR8AMU6MGmVzM
Y38nC+iEZgWKMmjell1TRAoE9ptjaxvhLFznzUFYkr5vzlaS+ZAzhgjG0fyPVThe
Mzs6Q6+BYsQ3qEJRtluBp8mtl/BMRIkshKM62XIDuZ06t5v9U202zQlZ5WiunWzx
HWQMPea7G/nY//pXBqTTyDCRATzx0GaE08UNm/eqBemfO1F1WQMGD0lSh6/SC6za
aerrYSpiG9qvqOY1crORowo563bVYDNfyWUUmZhyuZo=
`protect END_PROTECTED
