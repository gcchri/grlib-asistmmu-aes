`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GiF1tDmKDgc/+m1f8toxvyk4vPYp4GRwKbHwqoedIOU4wX9ayOmVFeT9KBBd2CBN
GMFJ6Uw1Y3UFEf2NqpbIVhKSEmPL0tWuxssJ56RbI6PjmJk0Dj6Y/YQzL8zCAk9K
AHjxTeZcdB5clUKrREM1t1tYa6hVd200Zb7xvaJx6dCpVfQGQvg4G3ziSztWRC7O
hRE1pXYbFtB7Rq5CLefpJM9DKQfcr+bwIJVAzMk0+job9VQoZN0V5zPbLHZ6Q7Cu
+XuExFWbDpXmtiqMTX/MtSJ4nvuH63dm1N3uhgBSJ1iH6DtoS9F4vcRBzuwE+ETl
`protect END_PROTECTED
