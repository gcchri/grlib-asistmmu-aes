`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zOzXFtc1+0s3Dk4FD/2vgaPeQ4FmmukZJpGrjJuiLWsqdbH5UctDeuF1glbN7a0h
TCG/BhuNRaylacEeSChW4ksnzZuhSwFk/8XN7EiBgXGx31UNUtuFMDZqtZMywqA0
+mv7vBMiBZiIeZQQbmUWRyAI7Ffl0DHctoZSzlMqMtCt1C5JwpfPZV7/WByYFeha
qYM81TRZbd9s3uhpDNyCakmuBK94USr5xjXtXzg0pIx6Vh7DRfOB6HIsgaGxjhPC
wV/HJvEmAwgFHGXda78c5YbZ9gqrlNcoXRNNTaUFRlFVBAj7SPIKuS1XynZtClCg
o186UnQLuRz1MdsNI1MyMcF3jGL2++HIwPUg8vqrCFMFqGZRxxXXJ6lTkAShaVE7
k2MdjUT+kZ0Lk0baEZCYzA==
`protect END_PROTECTED
