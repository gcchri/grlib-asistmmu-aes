`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6fNNMdDbX6HK9yivbdWALUmEilQqz4f0VHPn6G8d3Se2XTF5UR496mwiglahIXg
NtwAJ9jZFQnyLmF/O9TfWkbIQt6eEH7ezQpaobN1C7RkWDAzcUCChim0oxkARnVZ
66OLrgKwCd7bvarl45oxAypOpNFhdnYYmTtfmg8xxWHZkfncQjl+7iyQNFAyFLZu
FLgqIREENCLMzP8GDTFsYHXkly7Sgg/LflZvkgMHFYNSGmfnxsOcHOAQJN3JfG7x
RbuNEjTsTLdGsWuEg5xknhp3Clu3oLofrT3a0qQQoj/W6LWt1uZJWJyzX57X48BX
AeRlIGMMWfsu2yovExs/jJ9KFTcBUC/PpIRZ3cKcxQJ4NhtzXLTKdVm7jjfiP4tO
`protect END_PROTECTED
