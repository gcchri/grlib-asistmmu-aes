`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTPZTpp0DEyn/65SqqIm7zmZDhA94U6Ds23Mj4tauNTYT16L75O05Qp0MQl04VI3
fNU6bhiV7ZcWvqD2CypsE1PImO13Gi72JWZCMOdVOnh3YPaopzcWSHvIHOw403BY
4p2pqByXfIbK0ek6VxOggoYhc1WMtQrMuTjKe3q5FeZNc83PHTONVTewUuDCkU0Z
2naS/cyGuX9saYFG0IUkuMzEvaMD++VGTuMnc41ao9EzvrDs913FEV9O1noPjenG
aBAK92a0qpFGdPDqNCIfLrQ9IVgQqvCnL9fNzK6Oy3YjI0ptb7QonbgNxDnIFjLg
xEOhwdKteyDQWgc+mSrb9d8Qtt8V6SZrf8JaOc0n45mJs9cf7ciuxpYqJsA8jbKW
8bW9rP/c1zW4yfz85oAYVcqHBx31PzgMNtf9P25Symn+px24ZvLv0GSdSbQuOnYj
D1C1CCMs2HS9Fdj9juYhBLKY88aGVIQKKA1pMBPJjsgGbDifCiKpmfKkLeVZXbCp
`protect END_PROTECTED
