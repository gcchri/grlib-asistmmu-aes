`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6pjv4B0AU0DmYZMqRHYZqpjEB3ilWtv3Eku/ePldQV4KR9zCLWqI8enKYEdNaZU
MhhRky04v4JtlyWe3tRFNHfA6ur6xF/XGRnTj7tVpdOoLPRypT2p3PBBaM5uO+sf
khRBinJhBPDh8wPo5mHMHQimI+75E6fFM7FQQUuKDinvSKVc70NS9XT+PamFTSfo
2K+xyP3cWrSWXRa20GquRepWG7ffQ9NlmT09n7AOhY1cu+N7xnnYmCr0N5faJJAq
Ioz9NVUdyFltchJLv7IvUTI0wKhuYwd4qnk/Wl9tFznEOcuUORNyMcYDlze9fumH
2JNV5z1/FfFD57lyvGQG4Hmg4AFohTzYsoXm1zUY8ERNpUxINuH2wwNPqj8Xc3/Q
PAGLSQFSdEvQoqmmHpfdSfHf0MePB70kI/0WFzoQvveJBCMPHyyKTfyPhgM5xY3z
QGxc1PviP/K9dlkDfbN6cM2JVGWO3jmmBAmE6IKa9p6HmlW6URhi5v5D8CcEBJHq
rP+TjYNTlsR2GLHy5NrwdtHGGnESaQKawVDJs5U79ESjK6YsfuJhUFZzJyW5S5tz
b9X2QqvhVo5IMtAqGz1nbN6XnPJEOiigc/5nBWxDicatKGzzUdI1iqd/87U7241+
xjl/8SeWB+wcfaRXHLn4NGbksWV7Nf2YoOcHVbi1iPqpXBvbG2n0gLz8gKwNoTj8
6PLTOuiWLyD3VwKHW9bn8k1t6ukUNeMZQFosr2I5Qa2fUmAZjUqHFlHlODj7B/Oi
mIPIdjauM9XIJd1DIUHO7xqLbJkUTYhmO74WCzzsBdiYdko+YdGJoj1oyZ3tT6N/
gl/VD2dAIDTNLTApUZjND2RQl85GoFICdSwTa5DJwRTZ64UPMXJOS5Kn5AtzGtp6
XeTtiiL/i0za7HOcdhRDu2Ox+aEnsekXnsrHjh+reRDaSnit+Ac3YR3SYiCJTigg
454WswbGyOrApUsoOF7RELsZbGi15yjgTwULXQ4zs+Q9N5htldxsezSLcNsjKzTz
xEReuvaU3R/o6vfDPL4YgaiSxRIWx9OvYCQ7GZA1K/c/XqGkjloSfescXD3Jr5S7
zq+8VvbBS8UDwNm/AjIVy7Lf7qBBiwj3CxuLShIeHCpyUE33z56zsJbUkL5sFImK
1cHc5Ob4TX9Y2GMEs02bvFwOtDzvsHSuAw/f0d2OExsCs7BK1LtPVrfIJdRFYZ8t
EP6dEPtV7zFR1KLi9EZjIOYACPmdlMmC11FfToMlxG/YZKbHAWrisCAqW9i4n75x
sTj5Y3spSlIzJIGkhLragGqksUyXw5hgHijT4AVUOD1Lu2GV++jlopbZWBEGtIUf
kxg+0jaB33sW0nKdq8zxMvYXcGA/8Sl1SyPrYuEE7fKtiINxhTFE5Xz3+ShBSjfU
stenJwsXCBvM0dLjxe0xBDuL0q+UybJC9/LxOSrYp5APNFCttVsK+5uoj3PcmqTN
YztZrwhqGEUePvv5HARNrksuS4JOhPslTj56LEZrE3s+5NFYDvKLPDQXiXvF5l7L
SCbFfGVp1GoNd4aExBxL5dmACEuE4l3wJ/eRafGXNZLz3w4J5iF3bAkf9FIfJUm4
GdJhfaU7VDdd7pCDIICNNV5JEH3NLY4LRIqsQN1LZ0FrlBVpVmola/rig+XrAui7
NDlkObyBiXTcLDvhTIE2qiIBnII4RHWzN8kTVaj/wnQShBUIbDsz+nO75aqbjUO7
2dvbM0GL4anQ7Lm1MsT73oOqmSLRHXJZ4Lvmw+h64OA+EYIUO1Xu0xVUnaSFcbpr
wyNIyn/zyeaIwoxtTS8w2kx9U8pZotJmrePrnjsNgHk33kfLetGuQ375sjeDLQdH
5NFJYJK5NoxOZHZiBFz+BMyJs8GKn4oMW1zEM4LminWF1csLSHJPgnpZsu5NUGny
py67tj3VTSijxeM/ZJAKD9+16BpScA5J6WnK/5hcpNgJLZkjZqy5jMqXKgmtrIvx
yxnHNz/fNatyjA7rtRTBN5uUZhabOKmORDAyZNBs2rjmxzcvmO51N15TWo4VLIrA
t2PVxCBl0B1cTdMEayu1vtdK39t9vfWCv39orHPp4N6d4ry42RteIFLDBgD0P1oW
zzYX4CUfa6wTJOoaCVvEQjZlAHqrP5eadmK9eGn+5w15g0JkSNVM2sqWzxcrRRvw
h1Q5hs+AePKhJggQEm2xJUEIb2DAvm4Xnft8c2DOuC+B2iXmniTyl8vSRTCzurtV
l3vjvs5gB4k6O+wj0JFU4Coyse0CNEgN4g/rPnQ8Uy3WSsdqze+P+opbL2JUo40C
fej2zZFVKfKBz/lBJtt1G3Tv6BDyZa1lt6ESEYNSdz86vlRLVCSbuAyGeJBsgbbu
3ErhHLOUsg6n4gXLZW+gqotjAPhKrS1DFcFEsjOwcc9x2cZb9vqNlHM07nUPrN1U
t5RX7wsrWIidv2GW4uBUgQZ7oL6mRmEB9am/ONHkZEf21nzBJZRVhXBwvdQBjARW
wT7Tp1GLI/nwAUYpuvuMWLczors9ODKRQ3+zIIyYTCzrVq2WxQ9gcOIttsZ3ajUX
fuMasQS28jr/AGnsALPghUamUQ+D3471hycUZAUG8yNIS1iKNOPbDtD1bRfGbkmL
CU6mJCBoy8g/tQuQZi9ENUb1LXuv8Ajojw6gdeoSfo2/lKnnLDzAcmhYLH+DpCBY
tCMKLeggw+WfOrkHggHQXWPL1B0JVpZv3vEe1daYJvqgx30XXCPGOISZLZkbn499
s/yP1A6yOmUGw4CWDl2cjAVxnl3mO6c6QFaaQMpd6OGYPdHhxADAf82hMAzZwPW9
SvoQ5yDFsy+iuDacsidP7AP80gKmPHXnURXp/TKo0gN3vQk4sDtq8uPIJUFMTl46
mB9RFj4dtRjiNgxJHfE4ycRk9DubYEX/iRMRgJqZq+A+QuXtIH4ApAEItx2xbS/5
ZbHqyG4zc9StLD08q9kMU3L2tcDN+f74OE6JTwcuPpNEPuC/fxW2j76cKhbrjWvW
2YjAIRHjvVynLeMz1y04pqRoiq1DmSfJJlrwsY5ImgtPydyoVt5KDp/menVtPnFi
IHqlbSzYvIXq9uz4dYK2OOBAfMrLHDa5IxZtqd2hLMdxSfEiJFDq2JGImMxFe6Px
pim9pGuNtou5Eg1DFEoWtINPRacUkqQHdGaacFKht8YPAXKWgTx3eeiFzuNnDvmr
M8LaV8Q4DGExbiQanAAJa9I8TQemEHpEU0Yv4UvXEpYKALcIhufTBZBKYmzvaYkH
QQFJhDqOFp6J4oCaEPFFzchF9+5sROu5Q2TvTm4s0lnsCdPMNiPIKpGEQW8+Uw6O
dZYCMRUuANeiEvYySd/jOy/fV8krdVOHBpZ6I2hKQhWPSPaTGRhnKy4+ZG4VMsnQ
lZkFwbAOOrr7WMSN6bMTlYIkpl2+D5RK3xTEIOTSwqOrWFynjvRJU6uaIZiINiIT
u6I6a5+zfi17t49wljBIHgRI0+jpFyCY9dTKhbPJo9CBSBjHbSkrNQggFSRCs3yp
EOHLdoybU9rm5aP4yGdYqmJz2vw2NEoTOGPCxW3odKODFKMErKHrIWcvUNWCiNN7
fBY9NVtVv96D4Dz+IVEOwO42W8t2U9GFwzcSEqdS1RD0e9hMTYsAqqx2opYtWIkm
0bF3Zgg3YRB32o4TwFo1CBZtmFy5g7lLTCan6Ehscf7soUfI/CHRHBXeucSvnUmL
NoeLh+YFaTgvJ5W8I+3pkyZvAg2dPj4Kb0slHzULAJxL1CBiICZrmZPUzs/6725Y
p8aT/ZfKbBnzDouoorqwvzoAkShpzrMRN221RbmcuKU9IZBiC9pYo3jv0NwdSgrc
sFREOEA+9bNsLm6T5D1z3RRkbOyROtkj3x4N/+Fc5w1SuOhDugNEf+PMw9emtIUj
i3bibOJc/w+M4RISnnKzdEgKpP2z9BE5QDRQwmGXnK+RSj7xBsaOt0c7naZ+K0dB
pKq+WAER18m7LTZ+vzF+iRbi2aqvIpZqWo94nJM9jFdAXQaoRdpfu6FheizYyKwT
r0BfD1sXv3Lz2MDPizGHti5foW6rdqimqUocNoF/Ge6/5Vbkc6Hu/Hd3vQh5udf8
O52ciqPqB0RsOkon4ZIEAhCfon+mMusonOFboHCvsUr6RoJGkGz7k1op/LRoSAqS
lbLam1QxMctPd8dYctn8tLMebUK/0V9TAoLjfQctWMHSzKHHdKFzCe19BpKJr9Mu
3VieAFAMQbiXEzl2f9fN5WEc3FzFDWqA3/Z50+fI0/A/nq82uWBH4n0G8JCm8IAx
lHPQG21NQRZ7PUr9KnspKShHmmQZKlOOrQ8JKruD8VuxCi/4wUssH2UFPZoKFuV1
JwREv9ySLj2fzezbLbbl0IHKCdm9KwnQx1auDy/OkQyNeGyXi3XtyqN9Frpysukh
fBI+yRg/8ZI+sB2l9dtxknshZp/Wf2y8315SeKk40ngln9uwZoPqynHhICf6i8eW
S5gF/ChklaGk/YfWec4BFPrpj8c0EtBhMmSLVL4+coFuA+DW8wkQChkKLgDRTOTX
DXFuzFxz7KN1/FjDUOfowL+QlAi5H66uXngylWSbYniP+UaOMNZFg2JlXDIifDPh
1ncqa5xGOCt6lk+xusEDRmnjzWVS1dDkfI/cY6RSGI8WGukNmsW/cTuXB0nL9B0Q
TKZN3TV5Q7DvCbK3LOpAuYbjQA8yMr2SyNhy4ZDAByUyg7XuUpRLdhgQDeOYvsad
pN4aQUVs/wZmeOVPaaopIaxZPLYsZs0J9JILAMbbzfLJ7ze24S/7SSw/gIcU18f9
`protect END_PROTECTED
