`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fkJw6NwMn04Skv+VYuLx2gSsTOn5EMC5+jhSgw971YTTOc2J6plKbXNE4NfQwEB
kJu73Znc3+zYWuTci3DWvD1IEUGLt3X4oajSbe9xGFVHTNynHAioTon0opi006pE
wWOQbEuqlt/nMHmTc7lcZOXPJgb8ObXqnRkRxDaSX0PhGrKDfaid4LsI22w9Wiag
f4g/CrfzfLJtiV0ffY3S9nbc7wHEtCTQ591UQN4IySwwYA1fQur38r3G2kuJkrZi
LaYS4iPj+YJWzj0BUaYhEqIWVUfuq8tRifv+oveP0LcDlyKOyPueTifcOOlkKdv3
J8QBcQExSRamjih/4TK4+0txvV6/LJ0JrgLsOr1pL5XGLFxXoqCnL/FP/WWfXz4y
c2jZ282PHiAfIGb/ZKIbebE6FveM3Gfqwho4bsenKr3XZOX/b+WXaYD7hHYX2eaA
4kVKZLFb4uqLFJoXo+SxoWDbFU27C+BaI8pg5wrY1Ocm9YlioX12ZUyBKxVnltVT
oPjHmTmbOCqTmk3wD3oV4Dcycg4AY+MY8iLOc6F78atm/LBRioOuaZq23qYQc5ve
2tEtzvNuBU/Lx7gcATWLHKjQLTTz902mFIYevAABZJyulnrrEKjKO9Y3bv7ZJlVO
TnFnCImqTeaAQkvqz8JcEmkZ5mMGHJSSJo83fG6c+oqrwkahQDlWlRylGBYyABdc
QsgcvsPrkEvRdjrVAuCj4q8tScWRRXTub962WJJMM245+sqBl998cMtj8R8EPfAa
mByUxs4qpb9oCdYHHe/3CQt+gjLr0hRMFXYiGgRfdt47R9p9nQ8MMGUvaVVFQwtb
nUUdDl2pa5pHPUo27tw8YvqBiwSc+xXs5kofiH9XU3RWIIKO/pNeOupsBzBCpqa5
FKXxXI95K+rdg3RiMgwB9BUo9gFdSebeD72m2j4Jp6M0fhCKgrb34BiBPo4ZewP6
xNVh4sf8qu22+DLSbndtrCAU4BbZ437KU/vMMQ7jurG15E4052v0PXUPkJO6B+8z
`protect END_PROTECTED
