`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MktgA0a/dGebBi9aJQFO7F7fih3z8USDEIzMM6jRER5WmkGWnypr3hFCS3q+r9Kv
GIxNp/ek3B2xYfWRNyPArcz1d0hoXZ5Gm5kEwr+g9IGKyZhmiD+fNzuizfecV1yz
YjPYhFyd6mSamK3IMEhEEGLB2bpo9yM8P/LCkIul5+w6atEx4XHFyxdm2Gt3MXXH
8pq0D+kAXW6LzI75P6r1gtiJvGkD6lOG69nHpNm0x4F3ZYswkL4FSLu+0sa3lPzR
ZH7jPQPymA33dL7dACG7b1ASiDFrhCZgKVq5fPzDIHCZgohH2Cb6ARF7ZDdKuHil
d/gKet/Eyy8qUN6KC69fM9k9U8KtjIzuL5cAX9mGT3Qj6O97N+3/lndFTFbD16uR
1fJoNbPPU+Cv0MbeijEoVyFT9R0apRyL3xD3w0lT9rlkISMhpmo/3znWiEQdfthS
IPx7727M/RI834Qx68RR5B1t57bpaJOvqnuMkwppUhXKdRtAL9eTgvyId9n2YcRM
IX7Q0rls7hw5wzBI5jpdwE6GgdpY02vMufmGYX59ZxV+GsxQvMqN15EG0M6V0Wy+
ZsHM2+thLusc1J4EPN4A6kc/WdLARKrdWqs1MhD6LxeAECQnov9CdKjP9iYwiJQW
ee0nf5KuJf3zj7/3Fptmog==
`protect END_PROTECTED
