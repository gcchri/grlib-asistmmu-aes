`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DuX1L8HbD/mOjyLX4Zofffd95AtKdCve/G32MOcLGddipk2LoQsZmDtx4sVlnDWn
IcyMmtItHPdz4/VVMKQBwtmC7PW14Oa56JDLSkrqNi28M5uMd1vzKwbef/NXRgd+
wxsK77oIThmOZt70XHmQAHUYH/1MXKFEYr8LtZ/34SRFoL6tWdStT67Hr3zfzF/e
g4wUxpy4VKdmcwLQEvgMvSqAGE3ycMm6xqYK/XKx7vGg2E09C4cX4rVBhrdnxzvc
BA5E+7mYiNEXa5CcIyoc9VyWDO13YLDMEilEXJnOVm6fZYuG6aIILQ/XOPLW5R6+
QELkak6MOGMgGikcYb6owZusR2IeqLHZzHiBH63CCFQ2XRsqJzSzaPgMAWGXiuvL
lvkmO0oD9ujZKd5GHTTDr5NOwBRAWg++qXk9cHafu1svygKTECKVeqDOr6iZEaO3
Gq6Fkn255qrp3Mmp8MjmiJA4fEA3bC1UpcHBYBKdbPa6RMLdlPNb8NKzG+rdNNUV
C6kCzSeSHpUbuUPJU6oDnFvWhmNDKSpzKRA7uTzFXI5ANJne3akk5tRkV8eDL59L
bXvFBzUVuOobTcLGjyEvWoI/p38XsxSVjKovxl7mzpJs/eAQbQAs5XCBxhzbthx5
CsK32LYYLcG7IX8preStDA==
`protect END_PROTECTED
