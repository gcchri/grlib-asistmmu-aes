`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2OvraPHTNqUD8hDA9v5bcNJkpfUrnok7U1u9e5arEe1iFtxpotspwP3DzIctg3D/
ucOxsgACbrtumZfwWc/0F26ugjaCcVmyKEzNWHVldsVI4JSVebyP+6lhgY14XVu3
qc5wxObaqD0I9IUPvnHiX59UVlAHJSCtBETjE2WUlGgVJl1Hsqm6qmc1Ily2Zm3C
ouZ2zVOZb3q2Y7mBbGt+bTDts+k7IZZu8x/ha1rI2SvAdNNVH5KOpDp8UxD3YzWW
MITz4SX4pHL14P9NAysPaRI7lejPcjVJQKudy7CZ7o/HQ/zuDhQeivlGkrrxp4Qj
Ihe8GzlIYxm7/jmGXyJSV6ywV8Y086iRMs8VDmzRc+PKs2ZrqczfSuXF7EqifB20
+nQrbMaNY+V6RDiqxL5LSbcziw3GmltDi9UEH5SWFS1TunUNAh6nL3HdYvSJRfPQ
ZS04m6ZNp5GSGaIoGGbe8Zx/HX0kl35QalNlL1FWrYiTmoVUjE1h5Uu90260UOzd
RRGigjBW63YiRYciK/1z58kdoEM9sC8aimsSMmlB8fseP6BzCGKTBiN4RYEnQll0
vhA1BcavREVq6HLOI9l13hmfn0cLABthDyXm8r3fVEZAKZM+1GkqvBO6jISanXHv
42XbwS4l0s+FagtV29kYqQ==
`protect END_PROTECTED
