`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hR7mH2wwCeAg+ceuKtUuLVrVfhzhOjV+1sz1OXY29gevV5V2NOJaF5jO8OolOPpU
YfbVFHwtcZks31GVA/GMjZAjMNXZJrNs7RdoiEVziMILL8E+TcApJyS4dwjCJwzw
aAEsd8c6mCLdQ8YHK4IQEn7ZHbnyr0u/pmEDN+jPnbLifaGgrDvNcT9Zq+4Jab2U
2SC+CUkpeohMEesOYvF8FqM3bbDfTtfCUb9r55Omhu+GWoESXxa1k/7JdmX50bru
pJo4sESrLiIvp+rAvHuzSwbnhLwZb3a3tRgifpANZnL6LufZsCKxEv6K70dOm6Np
wkIZSmq/8RDqIBnuvZSa/Gt2gwLdZzQ/rRl7PvVYP+quEVvYhwx0N3ZSai8BYOnR
kKdZEcugBdy3u/+/vfMBsYiCum82tTQkpCAGc0K0OeTmPwK970jt8G9aqTMQIxSO
UBpjkfzqmQUFa4PgBPftyh72miYpZiJIFN420B5vfzi8a5Fv1lpTxB9xpQWqy/xb
bGaUrTrFfbePklEB9+5fe/EJbfWu5zAoklf2OqpGjWVqda/q4O34Kfvv5duLYJ36
FDZqzpdmUNwcT/vwe79+1D8b+RTq0I1ZCmZpO5eNV2FsDjBbh/91E9yUehtLz/Q2
B24kGqiqQNNK7suXglzpZdnFxg/LVCHm9R13mBaDtiV2BNxBFdeiFTLDIKLwUVZz
zi0Azulq3QwQamKArpOd418BqfsvZX1OLz084sya65WPYv80b29IE0zZaUF/bvuM
o9xgNs/Lw3L/fcuxdxbJIM2Zb7NIwInL7qseUEayzGVmlLg357F/gmjpwq+6JF72
7w+8U2cQDN2CJGH9O073W8Re/u5LcTGX+Z/i3kCHNc8sjOhmHjFAzkPWMVfW38EW
JuelwNcpQnSFP1OyJhrVq9LvuwEf2EaxSrsUr7MTKeg=
`protect END_PROTECTED
