`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBoIlL78Tn3DXkiiyunMFX7RM5joQddbzhKbYULZWxHwNCChnwEOwQCTcKIzgSh4
kQtN8fam/zJ8c+2osUcMkWfv/A5gmOh4UIE51Tve7KKu2Q3yUaHhuMSnE85IfYDO
aHJy+ATlUzO4qRpHsJls3p6JbXEdAn8gQxBIhk2ow2jMBmJt785FzpkOk0EosHW3
CQsfnvkNN4ihHQJcs9ejdusto0OqGh0IuRhd8d8yb4TBso4DBz79YW2pgFWf+yHK
e/pM+XVcOzoEmKNimeRMdJPOaGkVXAdmSWAZs+KnVM6zmi47XlE6T/EK3yna+Ep3
+jbAUP4xLGcgqKckUsfmLHFNkIcbsYTScTcR+cws+rL2mDVXGTrvSNMASz2QI0tc
m2j5q3RvpWJdoHNyDQbAlwtnsZ3oNE/aNXQ51iQR99c/rHTM/YsdUqXRFUWsdGUg
pJAr3yJ4a0Wl3+r+LkhsBsNFb9u7ipRhLbxjN5yr2ciVExZwgPUl0x7aYO1/b4lf
Ssnl/sUr7TTqg2O3fugQYiDyv5cHcYg2NqzCOoWmpSL9Qt4TIRGgqqc8vFoj/Vde
qA1zRAJmvgDS7c9Axibj9Ku5H9vfBqtNmrkpu9n06U1cwcTqDJ4qkTrP2fC4Kxhb
3CZLST7qSlHjh/DUYXIAe6LhXTchnKavO1iMXrFD09iqui9ojiEVLZ0iJZd7947K
9hgrUnqziY9hCH0auZ3WZRtkcLBSy5QjgenCD4/DtV3iXDNfeZHXTSdPR36LMT21
KUW4t5mmlBIdyIU9vqud0WDHYsHVu1lLY6r7AVCmu7jy8QjLtTeXJbtAuevl/SAB
X0rnDprFEBxHeZkfBqfadrS0RYm3EUxVXj8cjTCr6dYFGTTA759WQzja09CkLOjc
`protect END_PROTECTED
