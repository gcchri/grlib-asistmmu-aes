`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7brWjPkQMnWTxtcc9oXQ3UvJuPgZb/mH1ILLdO50icopJikwga3Pwuef/Dl1975
Fz3B/1/YkRV5GGmqngZqk3cJtINFYnMHiLgpygTOVDOVPtXgnOIuvQUSO8Y1k+4U
bAiY44CfNFf5S90Omethok3p++8P9pyV53Z+otVQWsRbUQZkt52k9Vr0V97pqls9
T6ReiyiKNnOaGtCFHyEg1eRScgm7r8z7iXNLIWCO9r9MevSYFdPVpJaW6VXpDtkK
xMSdaPURvRJl1QhIvmshdfcOkwBIxM8JQf31rQO/eqplNIUE/3s4PwhDQvW5lopi
8rTC6AiNBEN5MzEUh+8aSD1axjKJf8N9oHfyBWbVm+mN89HdkS21lpolUo0/aoxm
4JfRoZNbXqHjKYqHBy0z24e2xjZ9Ykgm8sE2Yu2xf2YcNts6zZ2xsvFdXtl3mfFr
M5YCsFwijoRdkJlEl6D0jRC3xHmpL14jwOcsZodW1mOl+m+5avELQKlBXKSb+8ct
yYgGvi3Ce8/rRent3BN9edoxJStnIYSj02TOmyv1Bd9c2LQ9bVGktxVbAQ8X2Rga
iXjIiVkMrid1Wf5p1LTdT+IUCAmrqKHUJYpLKp4gW8bbJPlEjyBepowqgDytDVE7
qVc9gfm0jQKgNQFsLMEjXpa4YHthQnXjorbQ50oiuQp8jG0bnWMPjhahnCwTqZ0K
1o7/0PaNqpn7lr+rCo69YauM/irFgsUvsiCsvrDR1xy5lhhXOvZNYjKc/K3XLY7u
/kpbsd5pW1FQuGdz4hDm+SBnpvhbh/E1JJhh6lmTj44K1+QhJAemEDd4b1JUPZ9V
ScdHCOjjAQzwEYmFIsh6FDFksgrWjq6z2D2BfE/ODUO//V31tKYi00PKtDRp3KIy
TmVWd7DUAoS4qJDAD1ZLGFbqhnzgta8KQbM5jbw/NdAODBcaqhF7o50Zqz/+LCwD
zmb9wUzSRPArRXVKce7XgTpnqfzVByYmVYIC44zOLBm3hF2xzhUHYeTEz4FlcwGI
yHWDbLNXCf9Y+j/yHlTmbKt0WSZN7SfO0VadLsV6uM1hMHAs8m5ziisAmvkSSdYh
7gB0GB3Sm6GqmAvZeVzxi3ukv02vHF+dH32Ep8t5lICCVBa5v/xhOltY2pgyO3Cf
mKV//pCKvLDrMTADumqVpY8BgZyg3NnilY4mZW3lmBcl8ER2Ph5PP/M4ga+ON6QH
m7UK/I7YJHO/CUkLpvFKgHvZzxd+tkXl88pP5UjhisvC4tyqoBK2kPOuaM3iANbX
kNrYyTlp6A5wAjRwwHJM2LlYECznCZUuMYmbfrx5MwflXryKKfhFEoNFKbPbdEwL
uD/VVG2Aqv0pgaSxqEO0MbG5sIQuhhGTvQkatKkIVsHewpw37cr9Iq+veNsIO7FA
/9FdUA8JGDJ/kxiCkjWldgtyk71KmStGLWAX30Qp+aE=
`protect END_PROTECTED
