`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+FuoFu/gy8opSHDEUZ8CsKTL01it31WJzL3pBWKPU4DVE4uUAH2mGgHrmtk0WqPa
kCyPOxjUyWxD8f0eTmuRSkwnBBZA9NpQrCWBtvboHI8Sag30WVrv389OlAoV+cUK
P2+23uMj6zzIxj2kLOknbTmjdc2g6ytrJyW2UJAj8gOBproX3PZVFd6siBJLo/Ma
0K0B5edyaqQgR7zwHJMeAcQztIQ/VDiC4uhsBRa5aIUvvE5L3eowLBg6QTP+N3ul
Hy0/FmsAifIeWn5Lo3u4MuUW41ujYUC5GIbp2rYOY3a9NmsTInwwn5lf6mjKrJkE
2WCK7Wo5zVGmbLGKWRFV2ryKZvJU2NcYCiHQBuBmmd+awYEmsySM7GopAMFNJGc1
xG4KNoWkgrhS/CJ5fKk5tKLuxkPVb4G7CkKnc/y/DCcUDsMCe4/jiG6sv7L/uT7S
6YOEc+4fP0AetuTYpLdmVTjPSbau/X1BFasBzvnAKI8tlc2c9Hv2wRJYGRKgyTa3
I1+GUYFTNiNVP+A/4DtaR7Kkr8aN+biEwgVToG7MaNdKV03tSh9bV76xUTpvAW5Z
GbR4lGW6va9UpxLUK+7omL1PHPdESmm18EkR7avYZDJ8cRR9bWR0+BY9v4Lpk+I+
nITfE5+V8pI+LpUumJpgk9CW6QV1t+i6iABP4zRS3vjMqr/WI7av0MZ6/jv+kz/E
aZyoH9Y/Y8QnpE2pG8CYiQ2URpD8wKSJS3w0/Kx8IGm8AtMB9SBqm13hian5cUSb
5/qTD16AfrIJg3rdvyOBq7ffUCgHQpBqpwxVvzGoCzcrNKBu+GyAV2VZUl4OTkOb
xDp1SbGcQdNwhPLkRwhdQ94/4TPdo8QfoRcFatP8UsmtPX4MW87wfA5SfZ01390A
yeWxPDCpzLMD4TqiNP7AqycKSZgu78Ro2LDj7nvNEctZZKVF111XEcQy5pDg1ql4
BoM2/iMO5Scca/hctYkAlqHYbgZrWScgG3nNSlgBLqc3mheJULkMeSfcrxjoMVHg
yAATlyDitAy/tRR8j1kE788RKst6h8HpL+UED5K84wbaWkoE3FPV/FACyxD/RxGo
ryqAJ8XB5Arfkx5xeSHJwQ2C0pHR32OausoyVmOr0tr0KQIMnqaiuDy24AMGGwWQ
PyOJV8ixHbS1TloTYLzJnLc+K+ltOww0X9dXqeZ2eK7Lhvct3+v2/cqyRBomoy5E
mSyySN35HWuyCic2iXsBV4ibysBM8KdxjRY6zo186U9r+9t5GUxgGW0B9/OX23dj
SgQLVg9OEFueBmOY5WUBdpIF8NLQBnkcTm+fBYQzpzXUF8IPXRl8c3SsppIlLaZk
QrSjB70rop8r92KtsQt6JBQ7ywza1n1dOG0if8jpSbUvySopnNAtWMrvXH1+vl7h
CQFUnQYsmdwH0/JMgGaBFg==
`protect END_PROTECTED
