`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pigIQKq5NwM2qyodNm70ZEHTGav9n6lE4uopvrha1gC581TB1LFl5gJEVGLolrj6
HgQBuQ1/rCEmgFSP7GZa6ekjSjQub4OFW4c17GoiKyXewZz7+aBVgGbbg8g6vPAn
4ELWSGBOeKILj/KYaUijmlfwFaGtUnJnDdEOoaHU1RAjhTyl64DqbUE6y2BQdgFL
mWeGJzz+1tRLHPd8uyMQXq7tu4xtTVi9g+4Y9Sji6rtfMrbKQK2/SJDcV9M72m0+
GJRTcP53/OR8ipIg05zc6dasiRvEYphVKHstya0F7Yn7tx1rA3rXoSRsRr/ZmpVI
ohNJMhlPULUG8TuBJKY80w==
`protect END_PROTECTED
