`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CwKqKPyPcpCc3MHAT0fs/eanRZMXoi6RboR4Y936ugMlZtbfdHq6LLCY4u1TbEoS
0cgaLZZV2xf1BJ/PAaq17SFIrK+kSj/kTBh04suJCTnGJpI/tI7LMDDqZs0VTkH6
0tnJttVUQ40XTStUxuBnbw9GmIXBnHtVohmrDNQQx+GIc5dBqDnORemoTsS/+zNH
NP+ovA3NiVCfuj6TknWO+rK8azFoP7kMfTNNg81cmjU0qUOBoeWzQ6obO4nWFNmz
RRHeCxMsMYkBlL0VQWyF5BIfyUHM67ZZMgf2VE/iu0uZowdDeQcU7xif33IhD44R
mkHeWRmV+vJrR7M53QgjoiV/qAXLa1cccZ9hcpDQ7KcB3giZGieOfk2sPElh0vg2
5TU86O2ICxEQuHG4wTm5ip6bhhwumD2+Nww/K46B7uAf6CD4TGv1RrmbrHs32pKs
wLyYaG+VEtaj9OzoA/Bu0fywvQySmw+HpPRuBiXGFODlZfzEtZNqSW84NJLBu/eg
1dYsR/wxWpXRUepd4CYrO5r75UwwY7yi3QBNC4ZNP0N3j4ZtK14Owbu+TQKEuKrT
TX6ZhfVu1evmub1AIgOhVBxb0dBoHrYTiIcp1KqmqIFfdYPZ8oZRKzHR0JZbSr9A
LL2MHUl4rpceUcNXs+YKgi/Ony0zyiRsdzSpj3VJWrGkqDGWtFRIYY2O77NKIrLV
q9knR1/Nr9DcTyAsMb42PdWL9Bzqf480kkusI3qotNsi2GtF4CguRh534IwAHMyX
ojnT24zQf1M7Y+X1/VFza9CW7cbNrHRJEJzL180cW7CORAOhMUuJexHzv5P7D6mA
5JMpyare4kDnjfFuxhhgWPSN33pro+Lt9ZjeGjbxCVR/6eJWh00oMYyG5wQDh/I2
piJwyxo+hSzGSDRafDlmLPvsANdE4a96bam+5S3J7IFCvXnV+RJLuDTZun35sjm+
GqMvF++JyRkDDBcVzy/1Jl3Yh/4pkh9KwTn5x/VAgG8=
`protect END_PROTECTED
