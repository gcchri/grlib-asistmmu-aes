`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RdL9lOdJG72zG4Kki4HwLZU0UKymMGWiFdroLHX7oWieW534zm3aw/BYpT5wNfsB
hRTzl+0YcRVCpzypmCb+4AUvcmTrXrBTEBppz2zOsWCK8zdvf1VKit2x8+0nrzxo
bPq3ChalLL3Q4y528zVftv92PRoffGacCR5L/qF42vKwQvKijKDTEe7nSQcwiijj
XZUlHGhaARIGb1pCxjLnxp3AjYge8h6wiAl/tCDkXaoz6QkPrjtAdkF09piF/7WK
D60TBMQ0NkdPwtyrf0SK0EGW5cUJ7iLhcUOS/CeM4Yjui8tBRQQvsDr1OcBgCJ8h
bbSIgZ3j7QJMbRyU1FBRvfcWIqgTDhOwAROLgdMcZrhanYKVKURlhO83BaKHfvoA
suwb060P4WzhubxCLqy+4TTnphD1R2eEY8fHzc8b8GW5IdLWvZtaS3yPnz9tMmRa
W2vxlhkZl/gQvTU3fXf2LSq19mucae4/HLuTuOYirLiSjN+h+VhKno5LhYubECWu
zJYoNkm5uq4u69/WgehPlIZDABBhGrQS0U7TzMDly8A=
`protect END_PROTECTED
