`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aEFeuugnTbcubR1XnEOFPT/ixEd9EaCYZf0TijWwQokNJdrKkRIFrmlDCNidB27n
8I3i2L1mnpC0G57gJmdgM3A/WxpB2DRGrTzZE4DnSlPPQvfQcECWsEKQ6TEP+Cw5
PuOdC+HDsxu7HkwavOvIZHYl1os4xo2VFnwIcfWfYh4CYpM/ZPXkDWGDlqoLMbci
j6TcBuMXXEeFPy0VXGJkrSoSfTa6+kFGauoT5SJ2XVW9IZYTjb2TVt1U8pFC0akH
1DCvHPbyA7gdRQp9xY6jGCOfjZLSOOXXlqEk9vF2GrSTFGz0gbY0yHdgp1dn32Jc
3yIKette4LdtW3jgXsbbY0d3SJYH3yxtGmLLY1JHNtE+FmihNCL27dXgahDcOPUL
iMMUXSqabHtOp8aagQk2PfMPAxXCBSKYZrNYQ0BDSO8=
`protect END_PROTECTED
