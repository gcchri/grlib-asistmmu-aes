`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vy9pd1gww2FMKxIkbQW8yNlEVCRU9VR3lGl3DHiRsaT9BPY7JZEOfX3RiRHcQkG9
0J42uT+Iol/GyQBwrku+Wf/KDqKT78zgsnMquLaZV+TrnVr4SNPaQ4GK9ncpe1Vh
uB8gXeqk4ifbM/0YdPIV4C8jAHv4d9cayYVSvp1bbKUNUxrxo9M7Gr7+kbBVCl68
3pnanMnXKCWgcveHAaERAHXUyupo4LCQRkfVIAE9TgYdzJx9x+PKKoZn3qmMaLpP
1WBBDfxGVYGtfv2TjnCxAdAcn1tGDaodGKoV1mGYsRzz/5p84GA67nTYZUDYRego
Uhx4/+1pnPrYjHUgO1nzHg8QJLU1U0D7FUH4LkYfYBb2njhhvplkP9iHNWKUTiY7
1tdW9UJAx/jgixJ8cCMLcN+YnEPyZ0hh0APX/zuqxmTWhuFPUAc14S/8Nd2Gv8XM
VlyW94oxfdZbS089adMYgbEGYjuI4e2JVjzqFOvTsPvtM/KCwX2YrE19LqQnXtCJ
vZLLxp5iscXnmWYE85mQHeM2y1B9wOhHeDLALFUh7ElUYg7Dkff9O+mOY3/OPeq5
AxH3pW/p/ymsaa6FTVX7R7yeJ8KbnC1oA61vudJnkJYYTrf5fU8LwJCPJ6ByDD7R
6rm4NY8yug7r2QNVJ4oce1tHOus4NVX8a8W6C24WPv4qAo3fy7LpuOdpQJTCmmjE
rcl1V+dWI54v3jLVIlOD7DBquTy/ySwZUPomxLkrIbozgelDqKauUE1hgEOIExr8
OH1BAvinVlrz/N34oLNgelcIl4hxWxNgbX+ytmHRwHiWJuOxF7N/9MwqGqBMzuZv
A1UaMWTw3mbtjMIkw+Vo/AzeBD78+C6z6khLUMe1dW5LGkaEjTQ8HXeExCqHrUN3
N3PlAzXB6+C++DBcRhbpNxb5hYWCBiL/gdVJg9ct1buJ+in4a0JhpWSyTjKkA8FS
EHeVUAfRDC5ip4BrF1TCJnHmEOnsDkGOr2R2ksNk2/iY6y7lsiwDtepPvCC9tCEW
HGpohUKZAP3+Y/Lxv9oz9mPOC4O9BdR6T4mOuOWWV2DJz4duplQEfam5u2st/3+9
aeiB4nJ6kV6jHg/v+fk6NBvXU6gLWf1hwBVeJcjxQc2RBWOtRoZur2c7X2YZgzoD
M5RUmQq1dfu+fcp5tw9KDK/55ghTSVzGNXfEmAhcgD2AszlFs+YaoKAUi1JUPtyI
e1CXmQbYI2a2L9Eh51TLJS4VkgkkB+xqQn3BnAE/TZF6CGLuJWPtivkeyz9PjMBX
cVAxAC1luS7qrDzcp2OU7kc9dCa5joN9uIusEUNWj51STyG8pLgQcTBGx2TisPvh
TYw+BIPSd3mugscOq1l5651I662uNzXF7zdheNoxIBUEDvI2yhSaurcSJ0EsalG+
e2wnI0aeCLOO8iY6DkQY4389zc+JKm6sCvufy9fuB4YDDD3Mf6enAjOuqcg1k4x5
oki5Q9WihaWylYq/uYj2NysLwQ46tOvEwMURTfqPjSm+k1KfU+XaeLm5GOHmIF6n
/+xUOhyIsioTDZKkvdDz87otv+DniniOfvO3mJJHZxj8IVaxsjYR6+NTeaiIKTsm
aJ96RWCKweApMuOpdSZ5b3vQb/CoMxil9zNXF9zXiheUVZNaDniQkIbLVClp6e5r
t/94xhKMqrnGs487cbR4Cou6M3IXI6LyoRDwMWHM+Sd4i5OXRjj1FjAG1n0i5s6h
GtOebXJepyoJNpi0SwCUeJ00RJro9CQP2WICbTzqnrLbDj4R+QbfljXpYHwvviFF
UFHsNqThQ9XupgIjaeaprhwkaS62uAvWXta4SMc942ti1EUIK976cWvMquqNNKJh
VIePR4BBWHozwO6IIsV9X7R2k3BDSPq9VGw7+3/iUUO+GmMSMki3adgLibJ7Ak19
r7NuRWlAryo+DPA+3r7y+hDTkS/bnXV3n1iVLUIJCoDc8yzF9JDoEwj1YLRyuRQL
SxSXwYiz0rygqJ/CAigaEskUF4f68uKjZapG6DQ7R/L01KoTucwueR42YFHYbWCp
Ljm36eGZDOBWXlOhLuoJVihXApMblcfU7v/tNK4CtHfYMHZE9mHQEFqs8BuqPVqY
eoN/47MVvFfVTYZHQNMx9ZY9nzC0JRX/DOfsom3SYdAz3EaK5gwdOXqKlbpsrvdq
efHhYwCqQYRkbhW/laNCga0TR/V5ILYpJSW4qjJB+CjT5D5X018GURM/9blGZGtr
8mV+Ms6ZA0ti2LL6aDxdHKHzRnmhujXd4L+NEAMbXg+eeSs8n4mGeAlI/UuyHR/z
HC4HXeyr0QynBNKO6GzWo7Wm0NfsAA2/bqRzHrfLvKshdWeZa0J7niGSnPc3er64
6CMobtc/IS4J6BIrGpvGEgdXwQ2Fff4zjDDzBI6K9a6lO3/QiQdOqr7Y3+mBVVxe
Ho9LqbstWo2h3pOTUqYHqbSJXLTSURfj7GnGfB1KEyPhd4N5hv7JEfCCP2QnjwA/
fHk1AloHCkoH5Bdgd5xi25E0euuv5FUKJSagMkatbqUlJyE+fchKU3zyvYUquxYD
MDRnBVMf9CEoe+Oh2TWCx2jLBFxa7LyGwIo0hmh5Qm0yGyd7f5aQMzTNe+wTQVwN
n7+1ZemcocmKSdvvMs5ONojktLEwWT3Fk6cVM8yaaGPCbmI4fp79RAKr1bADRoWL
Sm49TYZbB3zDetJeplfAhQ==
`protect END_PROTECTED
