`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQji7go3QKr5u1KMrE1lbcJsEmZUSfhcczaOZyprm0xB/QPOZ4BNtMM3q6yLaQuK
BKAu4HTCwNavgHPx3TwtCIMyNxPanhkewUuzjCq64xB0EA6lxv796FeBdRHEQ8wr
VLi8R8OBeASqMOVhpwoZFTGWnYWbHYd2+Ywy+GT7s1sVVusu2TI5+4JVbIoGmLw9
9PO5lnDSLDmlL4n2rEd6hlLAs0UGEv9fphLwuZFC5f0wLswXFULLYd6vIVEOli9n
tSihi3l1KZMhdx67ho9Pny62JnW0wW/Rnjai9Y7U/P7hZ4bFdr6Q+xkeSTJktOH/
C/ZB9KXyW8OMCZavZ8dA2dtvj0bpbni0/+BoQEZagK1DLAUTkCpuGx3OR671IaHo
UHEqDO3yrnHR30BQRZ7GbYUtbExzY9f5CDrtxDqjyzWQk1SPKoym+SY3cSvQp4zH
z2SyovcnlWIyd+zUADSJbcSeozW1SKY71yIK/2YvKkgd2JIKhJsusqSnmFbN7Ewe
qhMwI2vkqFj71SsKyEe01DYzMazg+kbHypiZy1tvLKqiaqw5LCbmzOTmmIZMXOck
8h/dAXBG7fQB6/sOQZ4M/+cj9MwnSnxYqEKbHd+yLLLt8OWC1lhAGYQw5PKNnOPb
lIdQWSXrmCCZpruLR4ZWFBJY3IUoqgaYPsIqMLtVjsZLWk0mMeugb7dkPDEY5vbW
kK6vem5/8DMOJImGL3GX3aCSZPlrTaHlmwk5BL4EWxHZaGKxjqIdIYyuEc6A5MY/
A7a9Ml95B5BoRsRd4Et+S+5YFynaDbHA1WVZV6rpluRaPlXv2d6nM3DsUzUoIiyl
b4JyVYlpecX1BXBWswFDcOYgdfCI9KVHsEMbjW5/Z04+zjWlgp+Cc726nfwzWcmG
qZAAMhf+WlyACaAQHY190/GlZnt/5RYw20iL/G6CNMFB/voN+j5boXhz3XBJHTlC
MlHnU+pWJtA704FoYpWIc3zoZRW3N2vlIqHLyjjf3f8IPP65ixSKlG87NkVlzNUA
tR8WOV2ak49YkUVi4ms1LHXlkbVyCB76TsV0YCgSShosNaOPJh+IcU3dReMHjTSf
6tD1RJrA9h9EtijQybNQw5f7tSqyI3s1JoTiBvzNbWsqQCIyL4X2iVtLx1bZhwfF
iAsD7WrvA5hzRxT9d32LycrvIb1tWVyXAp4qKE/0ww8BVCn49dxqSMaCeMJDhz8Z
idmTllEn9aEvi3nKzkltfTXxVYji2no3huJIJ/uojidUdNv5Zy5DLx9MfVZ7Y9Nx
bZsfLFzrYGbzmyYnKjMVoCT16+ZGL/JnDjigNAuv3750VFh6XVxq8NQvJ6P+n2QM
7lvyfcQov9OlcUa3XfCF8w3UJBNrlKC/OZliccBqzRde01SFFXW/NvBx42lkVYod
9PXKvlKVCDZgzK/YcfNtiAmT3RCOd9IuHPtM/5+po9pskCvTHZlHG4V7l+MEW888
pCdHEsRuTqi/hXHbJQy+Rkw+qoPwSaYnTUg/8SBAjAIC51V6S64uH14oc3GtBhas
HYFgAdGrJCYymfRN+0dVemb+DT8gJAh4xX76f/KsFR1Yhn8MDBvOtC46wPbMNL1x
VD6JKuQmBUysY3x6v+jwvsGjRWplIW0bftUaWd1eBFdj9EIZ4X8kC6YI7ELGKmKy
IjSIiC5q8TnZ9iGcBZKlWTVcszl2t688inaLAAGdtMn3bTROPbGj8qoI2fGHI4x2
nlHoh0tmJ3L+82+dNrFLnvu0PaMVqTeRRg31mZtQn7TXLHQz1Nsjc1jzCBYWnFkx
pf6Y+U6bHhsKJcld6AnekoZxy38ijPpTJ0MkuRx0/c5dJ6pcT+DPDpFlq0eM5OnA
uu8iRWUqGvehocUtobcfRhsIa9WJTMHGpECC3WxJdBiEh3qEjCrlf5fyr3onbEji
Yv41Anef4EsymPB9DdF0zlwm2TXDb8BKplvLY9kqnrZP8uYCcHtDDfcYU52A/fKB
qtBCeUxkImADspnm86M0u7TNktc30Svhpy+k3kuYUUSd5ztY4K+KfuinokG8Xz/L
xEiEmTCgukRUrngyRuwU1vtoCp6FSUclSCSLLQ+jXNazbA+rNmSChXeone/1tl2l
lpM0JErxLQj3Sj65cMF4J3ETtdM+5d/G+IGdihBrDt7mJNEEXumoUQHY9d7ys2iQ
B3YB4R1G3p+XeVtKTSi8dMsdi5r1F9iYieY2g7pEJX8JUJt1zgvYRCj21ZBm3bSK
yUq21h/G5neR8lxXOU6ZoZ4R2mhbN3BfEUnkvoOZwq+z0e5CY/0oLt/4DayBQ2zg
psSmaKUTOcY4Mjhhs5RBKHcNYhsTjT/Hx/BcgPqyK/oBtgPIHfbyCdDCXE03pLj9
RxsTeKS2yXQdodn62FcRVTCA7ZdOiy9T9bfa1w6CGAvsZhn4D1nTX6XwezV3GyMF
w0eDu/Pb195uyMm90zBIWYh2igt8oQ/cc1Ns42Y8ZEMz+FtTINCiKNWaAyJgVEgN
Ssi8YK1qLai5zHHtmLlZsaSZvU5SxcUIGkobf0jb/T8C/cbdfCIq+TUPy0aypNMs
c7T8w1dsny9qXyjVNCKQy0pdXQ/5bPcOb+Zu5/GZrOmYXS4Urhf/YhITpHI13wFi
n7NTB3+290v5GX6HhFEx43au6BGoJ5aNBB4mWqz2k4xnpoUGQFPu/b7ExkVz7Zj8
LqkhI7sLFoaAAPAv51WCcTCZZk3LRXWy3mkpE58d9vNpMHsmqnh11X7235xL3jWA
12hSTbnrBastmcZ7nVS1YQP+IlLT1CG+pK3bq/sWwubuvtjvDMU84xt7JHyQmw2Y
sEuw5fMGuIv1ZVsHU/FaFf204JAtVz1XHW+9bXA/bp3hhU908kb0C5FjVMfTaxpi
hAiHUmzjECyPrFbpmPU7qtk95dHFJdHMYUmtY1/FdJvl3Gyp3BBfzuBduO6HrXe2
kqYUNff64RrNPSbvkmEc3fuXtAJnxN027FtYWzN0GPE+aE7tt1vNd/nMQftC6VIM
0lSIq+X3Nq4MlXPubO+7bXnTJe/kL7TVkhb83B1FMFgBEdh6B2y6uxmImtOnBUvl
QOg6AviZtFFFrzpvwwuHHizKZEUoRUwjzvoFF5ABK502YaIGsCY2WGGz5tXvg46e
hP6UyQH0Qhs/fmCIHsICmiwkqkO2Wf7KM4Q42YJBT3F7zPCeAHSAACjzg58AlQLT
pCjxr/rTph/IQmpHlUw2drXBRBt4NlsFE2LgNn4gYiURJToEnuNmnhCeMJ0RXKC2
Zx18NO1YzB4oM9361PDIn6Wt9x0DZWu/zRne4LNq1vb8ZZVxIc12jtVErj6fU/v2
+UXvFV8G628gLKug13CJ4xJ9GZqD4rwOSNc3jTbnKqJ1za3n7fX0l3hl9ZVB9TOC
vuZzJvbqn1yy0TPqKkVFo6aYcvxliwutnqqAFWZ/pYkshNAxj/lZBcCK3w2WWanZ
huH2+BRpIN9HvPRD7Nk5oLGD2JSoRBgG+W7wGG5+gJYw3MqQFq+rb6Ow36Wv0DkR
jEl53IgBkN6OxZNDZTTvDvVaD8LMMtiscIDnM+OkBo5uep2QTubIfSy6CusoIcK4
wmNWdUoYOKyTNJjfd5/YcmeZ32w5CrVFyuTx3VQ7dpD84u7jO2nY5uehweWtWO5b
tMnzMK151oCkWQQ8lUrhPduFPIFdB4jj1Sw7ztjG7e4TRtNFH2xiJGDSVXheGBtc
DO42g8zD8Q5f1SNlIfbf9iFo2b3QHTVofgFt3On1g+ZUmqjfEnPStGPIB0Rh2HQk
cN9q7k66hxYcn0eL0D4zbV465hSTFqTZALZb1XUr3MtTAFeA8WYfkz84e5GWp9IQ
9j32X3W/5Hr3m+m+4HOSEoRaS9FqSmuRD7bf7QRzV3yTh5qv6HjmPYzIe3TXk6NG
qknnaSI29VONdyVAJaJRNzREJAGCz8vUjAhAL0NyWTPvnC/dYzX/pgdeLaPs5Bmi
TH/jht2XML3CMwu6fnhdSZvBMwav8C71pPKvVs9tgeYd2sd6znB5sPD+otmIlizF
s107CgIycJByhyQZt3EgBRTAy3UpjEl7/TbD+fqO4rXcLZMRlUeq7zGMeXSnWFRP
NnJhljCtDA1j9OiLL+F+hQLAiEbNF0rFQEwMv7ZKhksdoPnEH7ONBnxuSD5bBCEG
PMjRVzvtSWUOJVlzRjgZTtwo/prN8LyrDdFwDbPQyY2sTNRtE8GJx2l/Yc7LXyny
9hIN9J1js22Xzcylm+9RvGuecYJJk00eIbdumPDI2Ox/fD8gp+2dq57x1Ig5KbC1
Bm4P9mY38if5XOsloU0TnozYrKl3ZP0qJHANt8BIcU89Rv4NUM4/Gqmu0uPTWfkE
pCfXh+wWRGT8V43YbSNVnjAUUZCJeIuMS4LvctuDnQbg2QEeN5HqplmYddysQzkT
jVMYuHNtFfyfCozMqBaTqv3J6mqVulu86HR9pyilpG86bi33r+fk0lD+F720VVbN
FSGBR3BEXOIIAneMV8PuNaLkLdEXGy/CVekQQRjow9+NtwqqMvMFBWKyVRZIUCit
Qeow8bUHTKPcZEjrgHjOK/mixENchmXF2r/fq3KnxSGLiNrSfioczqmnkL/sJZob
qi7JGGwZu11qMLiqBM7GwM4z+Z1koa1rYdhH6r0INBc0fACp/h4tfEhBtIPhGU/N
f41kSI1QA6mAFnZUcpOaQvxILv3AT+VJvXO4pHktugET80k9+LnASpYjXUDtFIwe
dy/yyCt08Fr86VP7X3HKZBZXcyXCEQxvDbVeSuN/RPfXTbBSEnP6tgRyBwlzmPel
hJ5mQhFgu6wPv+TiHei4ZU6dXir/NR6zFm6keEVUqsz7lNEjtsuuq7DEb0UnT23+
TqhSjLTAZWe59G6hExuCvxjEStmK8wHh5lduKElAuQTwYSjKR8BT5igPPd4u4dkF
yJ7xb9+YNYGj+8jUgy4PE2ADvV09qaUmUP+jm1H51GMH6UoSu80uFCGAd8vD7sxS
uMHCJc3pYOtZeIWPniLGnS3Vvr1ra73zWoH9Mdst+4JF+McnraNt/5o86EZwjiU7
Z1M8N3+6cLwzzShjWNbSl2i+fYqHHmR1pB8IjuTwIeqUmHQRAGJ9JKI/kPER/2Sa
gstsHNNTEkfPf+lomN2S/JysHm1sCGTIXvLS/sWEr1VHYmhZbHo4zHbZnfuz2qtV
3qcxSamYvsaf1WrJwrO01GKQxc/cgPM9DmvSRa9SbAXosS8hJuYfKn6lJiiSecCi
EqJAoREkTz8wJ1dlNpw96Oy3SMdOJ7LadWjyt6kN88iXS5loWEaYZx7lA+Gp22If
wnZ1zgKbt+QQlP3yn/riV2AHU5997OIkCnrnxxXl2xA2xUlVZNgxhnYVkKhFG/gW
VGZiHBZAjWzAKAuju6cc6eX/tBBjmobnmyxfhgZ9X/ErB1Ye/dHZ+Cn49ntn7/j1
xsJfVBOO0X8L7PdYPm5nIXiOuMj4qwNwBOwBggxcV4ooN/npiA/4KX4ifTbHI4GE
F7Otn+8KcYHNYzmQntsaHQKAmzoTXx7J6tgyoXDZBnGEaR7jApMds/qYrFD7/JJo
bIWo2ksbAk8k0GQj9nm5ZzpHyu46nUFFRisgGLCbThBrp8QrT9NAddcHGRjMLvUo
Ikw4/IOOd5lB9PqOXElF48uwHk5dnM4U0iZte91frObuTFAZBFugngC54WthVdtD
MsK17f1afaz7y0Ou5vIUBENrVhCYXEtDEv2+a9JdwLj0qqFl8SJzAbN55SXVFYgy
msJ4Zjtk66dknF/qddsORAph/RRG+dD+3ds6yvTeB2D9LgrdjXoV+QvhTvizvhY9
KYMoFjs46i3cldHHz4pS8fwyaF08247GZGcGYArBU8wIUSZntj2ml0ZYmincDlnu
1tOYim+qBp1d6LeDCqYDsiBHdgAO1yJXxubyellsRps=
`protect END_PROTECTED
