`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkPUZFDDZIVzG9V0R0jb+MfyiPYy8bZJjo1ZltGpgqzs6S29bbeaQiNUrck/33If
85nwp2+HDkEyxdiDqbOOd8WQneE4FosOcBE8UNVJlr6+W3no3gsDN6fOf/vxj51U
z1dL2NnhI/vDxzg0Eta4s57lThXRWWlYGPi8PmP9fWrEfNmEZYf/L+D21HIzROuz
F3AQxO876A2RuAHBjiH7NinUm7F/gbvKuAssN1LuMdIxnSwxngj9Fw2ahIV3t/Wy
EkeHRb0leiqdXrmwFoUKV4urJXuMfuTot+rW3ZgdXwU=
`protect END_PROTECTED
