`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Pg8dYIEK+Ojzf2QbIWOKfrbBdteh0B2TGZBtK8qoS9ObRVnsat8JVoVFbYF4xGM
bZMbbkf/tvuXcQv1Iv4AQ/HgjUvPa+GfV9oHxvnhBDnzejCDci0Dip5alij18gdL
S32S7qDbo0XtPQ021HVMfUAZhD6b5jh8uljbsy3T2IggwxVd7woXJlRrvjkZxeeH
x2bRJx+G0jy2XpjId4js8/b6l5mZ/SlXKb3f+UWsEyOFZeAhLOaNmEQjTDofY+9z
MvNkz/Nxk9w/KDX5H20tEHfhFHwz3RmwMbL71ldDwE7p72rvaM0LBVXIJacfT/6Y
QKUtGPILB5sIdVKO9B5Fzily2SUqdL4bEqCJVEwr24sCfwDZCSjfCv33prv223Bp
YPTzm0aq5ezp0+gUxcisBTxXZA/h92lphMRWfLqX9t166WGpNGMUW1WJdof5ngFl
jdzFHOp/8kYNCFlzDA48yzOoxw31mpcsZt0vXe4WOkjDpCAKdxiB0cdPEiN6xrIh
t+zf/hvMcHSPyppdq9+jtBeGjZdsbiL/jr7XzhyEGDl1/0zsmipzWOLpWtfgtttu
Mau+FK8XC5W1bI0feXdR7VeBBxTjD0gorGSyZ/1iJ8k=
`protect END_PROTECTED
