`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i1AcQQykpEsS3PkyAFwPjq9/yC9y4hUCI82BQ9V6fF1HsjTNCBImDAeJvJYO+2lb
5PWDZAQOXJJJGSAmvNrPZAMdElHCIayNeQfpQaZ/eqEKOE0M9VgYbq52TewhZMqq
Js2LJbdFoT5trEe3XjtFaVN3+jLMABT59LCi38cDSubvfoxTezVWW3nq51Rv5x3D
Vdo4TqXJo+Dd2VGutwi77womX7bZowGOGXI3N2VEXm5Hh7fW7DX4G/cGZ8qWI7wh
caClTpYmaF7RGHBennN90wTFVzVx/BqTIpMslC2iJ2rK8G5L2/axMVULrr34/v9Y
rTxuftDm/9m3H827u3d7uxed6+oZ5YnSCfkWu/DBIukA9nPIfwV25ntMvzgvw/6H
5XWgiWHDqRZmUAaaSdPwHsOF5wrJ3O6Z1KrXs0cBPi+1f1MHrYqVz3QpWd1Mqjkw
TiZ6WdfYRP2vYgzY5h7es/jnbQa6RxIbggjXk3++1evqGxi5hPiRX6kJgEQ4AflT
/N1ch3Q73l/oLCNeNiuD/MDl2aNK5qhpNj6jdFtZ1hZuJWkp+BNyNwGSPD0PivVe
IypdK3U38jCLXC4hN8zsxKTPiQOKs87zqGjR3bcUR1M=
`protect END_PROTECTED
