`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vb9F6nGYAmeHaDANvmGG2yJUfN0magCum8hBg0oBcMGaiYvfJkaCSfG899TQkEmK
AQTUbi0eXPiEbmsyTpXIiBzMfIOai6cOYmIQoCqXv/MD15wjjc5pxbbR8ZhPjjkA
/WcjJ8o00DBEF+aRX5ra3Td616qkSKRm0hBU/qx8YgXefWlPbXTHt8shCocPzFLD
3AsQjzOI4gzHL1xYIUzJiCFS/PLgwZ72vf+icQtx1+nSGNIRjUg4cQaGgkzl2Fa3
mBA4PwMRGvTUitRyyeY1H2uhYNvKiDd1nVnyyzcaqPBDsDXYGEbtbpy7UppfqggW
b/S0hwyAjNg/ZXQYz35hRcZIPkOsD9Qp9cxxhKVB0Z2zTZDc6jCZGsCxN9/qumdx
`protect END_PROTECTED
