`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGNeDvnPvxqMr+79PdfD4WmrjTN5qxI11yWno/l1y3W/bZTM3+ufDcnr3SIFBl53
sfFgFobkD9TQAZdn1zTOr+KCAyXmtXM18CT9tyulQy43lkUccx0aTSaC31GQwH+3
x+qZbMcKvb5baZbx24sR7p/GtTOfsfn7mGEaRd9+hTHBYycrJ1N4OrutV5xXmKBi
ETIPHKNvUpOLzLdBz64cMQSn3k3no2Wphn0lvsWHmEoflh/6LRoOTGtH/BihHfdQ
Fri/T84MgL6m2f/UKTuQ6Qtl7ljbK+YesM2Qqh3bnEyeOZAA4kRm1SdSRw5F4y7/
6UjIGM08nGUdjPYWLJkWtTaoenKThxtKLv52bFS3z42aOqFLvjk8tc1QKANX5edA
UFj3nkXXUDyP4Kis5xC3UHRDaJbQg2RrkKU/QJIeBWEywRjlzhTGEY0eLaTlYiKx
yz5c10DoH3pQmoIyG/vgUt6GFH/yqNkLULgB0VEmYzEtern2He3AOvjlIIofB3q4
azLHnyDBggySMzY82MgN4yfKsRAHzgagQk86w/2bvcUZ6z8RJ16s4KzCgQO5pJyF
0ZDQo9eA3xDgLWLihdSFQiBG4/3DJV4ojs9mxHB22js=
`protect END_PROTECTED
