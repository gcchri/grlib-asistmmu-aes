`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fs1jPwNWoVC4IQ683sdJtehGCQ36FK9su/cTxPKS0ReTgaIzOKy/3UDiW/G/ABJ8
lRKzjDavX/lz8omCzoaQnlH4YVxGfmDCq8TLNI9qRi40fbxhgKpguuTK4euh/kSi
o648JGc9bWWguGZc5bDcXssQs/D0jutUrY77wAP7OF5EvWkncvAsXdJ2zRnhIiVv
/7hZUkfc7SSEYcSbitQIhyYep1clwNeN6pAO9VmGJuLKCTg8vACh3x2WxquHc2tq
CWTkOTSZX7bMVEtos6nL+8rBSgqeH4Lcmhqw4o2Y62XsKLwxDWA/zC1kbWtlBaKV
x6ywME0NQomOHO3SComaWnCbC+b38JgfUJKAF58Yxwxh0M3IWBj7AZcXux9ezd80
vOtdwtnFDJLHZc4zmiAnDs9EBRb5ACLNWwAWcLhTftk=
`protect END_PROTECTED
