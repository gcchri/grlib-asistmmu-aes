`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ga+w1+qHlYbInq1TxtcMaqSGakFKxd1wGZ6NLfbK6wxi0KZGOukBJOb1OckAp7d
F/qDsWJQJQSRNEWEnNM0wDz7DT73PUvxZB6a9t6DroKo1mV9GSk7Yi5Ynu11Wpfo
Q8sFV1kJlSYBGqrgQtk33DPHUFYHYcwJ4kvcMJwsrLGDA7G9BkjQqxARgUXCVEFK
aqHCfB6cQg4lqJsLN1y3RSxWdd6MMq70SMEvt//ZBpqRRIB8nw7/jzANeKNx/BnG
Ic0SZF+iE/w/N/cakCf5777/l6eqlWyy9yYyfNcIU3Fz6e2N0AaIh8UQvTK9F2Eh
zXTOz3BLD0px4p9GvB2jhes092PfJavhx/OSMAsT+8pJJoBL4Ode1CkIday3BIQi
329OniporDNmAbbXOlvbITUm7Z5GRVuZiIWFdMpR1dN1alfJ/nx9XFUV0tOJ7Dg4
Ttpdsoeh0qJXrgY/2Fir2eptIMfqemqI677qk2YAQu+wQm9MmiTq09NC6OF8hJmz
BfOAUvwssc+bBTb9YcLDus13pVZiMpQXE4Bjoq9ZT3BDx7eZCLQdMoseanXByFzs
dskTzyAZUCYXZwD7VGb/M7tGnKB9pJKbbFHJXCz5gbkYvIAGYE+thJt20oNjBW/D
rIfeLs/dzrRV//IpxHuA014BARKBGkYzlpN7crnaY8mQyzAfEMPYLMrJwY9dKCSn
XM4q+5YAM5QyVcZ8RdpWGGipluF7ypdziCQIZW4rGcmpVpzXnakukF9o5NsdmFVN
eIEKpm0EHcENSviAUegjiUG2Yqaba/vuKlGCU0rV7Fv+1gAo/nYL6yxV4sZPodt9
Bz3gSVFwr3UMmv3SjeqLpl5jlMoy1oyTa9ZS5fX3EyVDuE6V/1k7Ab7ng13yf/bV
mHKRCIEReTdTOBDuGFUHr4Vn2tVAd5ZscQ+2ue5YjqHSQtI/w0/TTXbPCvkWpr6r
40dJWByi4xtuWeN/yaIjTE7SIgAz5YTPXhouYYkrLHpHxSYdJ+8JrkhcKp2PgZ91
SI2dwKwyP3HfL4bPNDCtEyMOCEDs1Tr9ZtRu9brwBl5jL7O9StwSr7PxMe67eWhN
ODtB4dKC/3Dr2m2kghP2FygNzthrnLm40p2yx429wWSvnzTHNKDHwiuPNYb6iDMH
w4ihNAlZwq2NXogTkMBrh56tJo1hTR/GJIs2tQBEiP6TO6J8Pg53DkCA2I6Bfcrh
EErr5ZZb1CdTmpiwV85CP/esXDjoFeL4noHEEyoTjeTjh2m+2tnqYSbxpV8y7A6E
90GDQ/oElsZ8hB+2S786pMhTs5M2L3F9pIzeBRVvZm1eqSvarpivaxiqJFBISBZo
qVFTKBPc/WcvNwwq3v90SvVtEM9zVLl2G9UgV+NDsFATKzt+XB+2+lbPHGp+80k4
VzuIZ0B9FD5cHWlYCP9ROPPIah24L7MkXKgKS5+C+lPc0L90IWNatyOSxLlDuMpp
3SfzVDJF5LIlhvS9/mYvbwq0QUiOkQly0NgDBoM2L9SVvkLZsV/3vQInzwXsZ/Rn
ZhYbxZlPBbivd2vLNAX3P6cArXOl7zsr4zzT9LbVLnacMvHX00iSQ0UuULgyEiFy
e87m/8G+oUrwlvLB/dzUHCyE7j2AqtzeClBbdL+eRgyW5Roq4jFQbfcW46+rlUdI
gyP9FsrIcnOgvazjEgFk/nopFa6+aA6FVpzF5YxWVzMTjqzdZFD7U8uyCuGTCSFQ
1k1lOo2vKekmI/c8E0AL2pfejh1kAe9tuCuoywdMrx6nY5FsXuqr5yAHOrDpcT1H
VOuvcQIcZWR2qVyzPec3LUs7AsDr7qY2Pgz94kG1yonO6q7dhvVYbhb9XtOX65bG
Udx5CI5sMh3uswpN/43OhDDiRS6jWQABVmyPbAUFQRJKSJWpZHJZx2rJ8r2oQxvk
b+t/5BBI6v67fbxvo3RZlFUTP58XftTDMPkvNTuTKG2qSkIaNMN+S6CXakBM9B6d
tYjp6NVs1nwHnIhJJb6utxoYMGBs/m8s2KIiyzWhqKwRfyFPPVUpja1iS+qK89PY
JTe4M4thzGg8eT1CLduok2zMQXZ8gpUk6uOzmt8bdS4NAwChVmBqfOM1BFJ3trFW
8kGBNPVPA6VOTmJvTV/EWZgHcQNcJs6itPS738qkXeFO63hLj1gXXcjwvF5MR2Xg
cW7qlqwNmQ/7GKS9+Tnda+1vXV9uFXOoML7ta1jYCr96hYk2We7RMdbsaRLoX4ID
5w1uz7hLowOvEGfJ7L6usQr8p61sMxli/J6+gNUhMyzoV0UVr1VP6RVCbPEDx82S
`protect END_PROTECTED
