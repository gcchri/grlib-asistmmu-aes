`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4cTCeOVxrPEuJfO/Q1rPQkOpKhUvPo5OBRgJHb5kOfGVldbGKKVr/mrbroi32j6e
Wvn8yfGTVCSBbV1YtsaI5Bvomni2XYg+29OC6RiBsS4bNj/fALxy4N5OHqc4ZaUV
CkqaGu8pVl7P/5b/tDUHw/ckZYCf4L8WiC6m2Qhfv35HKxm9vzRmQ8qk5ROyXSLH
1MB3RRSX2urSQbuOR3fnlXyDxGuljJSjSCsgLspVzqxl+rz2P3pozMMq+vEFF0/L
Jjx58vSc92nJR6ru2qoDTUvqV/l5d91RNGtZBICB8o1xgNU2++4NefGE8EJ08QCv
1V7VWtUrvj2PpgMc/k5S4dFEkDuCnE5h5DUdc2lXvIGEsJ3RSfXzbczKIQ/mtntE
w0iEHe40VLx0oItnFVQIf5oWYgTpq+XnR1Ryx2bYeIBZC4VcGFwSg9iQZKlb2mOQ
3L4EJ9GOfVcejvkb8FxMpaIIouGiUCRNWt1Fs6RjguldGo24bo6OW8hwkcWGSj5Q
/RDMCSIbzHLe8Pg+ZifNFAKZIghw+bd/NP/n7PvgQt3PkF71iIDXC1gFtILcBja3
EhJCyJ4x4XDqj818HZh1QJRvcpKNuYx+yLxM6AU8vUvt17KYhqx//oxlQYuj/Nbf
tsRxQKTtK6VQLJZAM8Gcgd5GlcInmYfmAXvRERi2Rnki00+IkC/J6s+YLKKxRhNY
DBMW1xtpW6kRQ3XcLTJZ07gYm3RsMVzaeNOerdTC/oJiWPgYMD67x/+YGTcgA3Rm
4FNlCSViZoiQyvUWJLlZ2Ire+eBWqdP3qhAZYN2lU2XVGb0xxtripMtsYGmj6dA8
8tIxF6PDZ32/f7c7OpO+CiNUOrRytxlekIKy3W7ITUj5IJP9rWnlqPEBIuDnPXC2
40j7+7KIHmv0SMHmZ+TD72AuFSvBlg6uORXbqI4XUdTe9CJREepgeSaBHgPQkoMq
bNoLkG78s/eWlyaiwWUiTme8QD3hD8vY8ULv+byc/F5+/0BuR28xkyx1LMflFTQg
MJx6A/sOlvR5upnqZbq3hClZHXIpq/pBOinOW1VytrvSTQTM7LTYsgM7++xeJ5Mb
AVm8d7lp2UsZNP2C+aYXP0AkcVlZkrB3lNFuWU70anzmWV7FwtI9r3ykNGvcUAKU
gNAbCrryaw9LTnErYglYQqaHdsMG3FxZVjJERodUTdhxkPGrPh0S//VBI6pArsFC
dvjHKdsQiCcG7qzqyNLH1LYxoHrpEoAdCIrFSVj0g1n8cg80RxNQLbNKUWGHufCj
gCyg8guLq2V34YNRYvOBWw1Ms2TeFwhAUpja/hB1OqfmcGODpBt7quSZkk1vK5w5
lbWJtNgNB9QMWljqIKPzMPsk8QMqVB4PMjtOQyyxNjDdNPFss19WifiCX6AQdx6G
prmIPd0DEtoV9amiy9KZ2hrLFpSxhv1838r872ywG/xcQiNW9l9xelmBEQUuWgG7
`protect END_PROTECTED
