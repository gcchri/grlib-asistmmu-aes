`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ngJKsb7neGQcKh9dwTOxOpcuqI2ncQPJp/NNgV+5ymSnQC72XVaNLtvLT8HJjjk
eCpMLmwsVvI3bvcjoSFPMrpwgUWVEDoMOyok4aKXxkq+Jc9K8wNP1wjodgRnLhs3
OLFMMPBWAz6dwMO1snCWi1zqjBNLZP6hBQM4ZT7LBAV839SHoLZub/4QS545hng5
38jkdryRvU6jJR9B2uerr2YGcOCla2DJT3ciWVnHCr8ZlaAfe1ant6h1gTRK99Ur
HuMcdiag3Er8bueHTc7s1nw4ScSwSiTAi+Pxsw03G5IinwMwuLUyphuS0r7RQQ4a
8phjjmMOCz483LrFNJE33WAxGdB9pRpJ9Oy+Bh0IDUw=
`protect END_PROTECTED
