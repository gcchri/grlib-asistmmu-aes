`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAZtQ8KGnBk8F1u0hRM3Yaf8y+uNUwbuufa0ieYUKuTeTR67JgZUaNOTuloQ9MvO
IZp2ED/fppAs+EyxcXzS+WmeCe36uTPR/8cl4ckwGaBDzOi6tN0hCBY3wH+rrHgB
G0KrN2YbNZpfMaXUlVPNQpqlULzM5sfJVdMGBKMZoCGcCgDeJxVkcEADfhR5jAa+
bC76/8dtCNrh7KmFJY2LtMUp+qPJNF6A8xcofSHi+8yuYFV5+5orjMsp4+j/CxJt
Ty9Ov6tsh61ZFcVfbVNBaP8RQfdi6oUO00x6yJFKYIScuHlJ6n3y4/xxNI97J0Aj
Pq+353hS9WvSjm05XMmbaEwS5PZj+GRfZ6Qgew5/LnjEMnXh/2SiGHa/4XVfSX54
oRAgT2mnN823JAz8cVRzxQ==
`protect END_PROTECTED
