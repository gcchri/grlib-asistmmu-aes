`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdArz5FTr4HMiqQPn8IvohbLTgievOwirsriSwuQj2HDDf/CVKtleY+rta0BW0Z0
4zoRCZBFLQlWUjyXUZlLTR1+egJcwx/jMGnThm1LbfxOe6+P6Z6yoOEMn4K1+LqL
ooVpAeVh+bBbqkvt8VguD4NdOZcdePPhlgEjSX7EKAZp0Z9En8zEljpUM70r8C21
JxJG/GuK+KpFUjuFKSnbfFNo4UJJ8R26H8LthGiz7HPf3NjD6CtONBg4r4+y8iOu
azBLLW/GGV2GCj+8NW1f+r+zYN/dRXQ25idHjp2MQzznyjL5NJpIJa8ApTQ5TMJg
pRwy566KixuJmOj5wprzWgqDAM5zTgFinlat/Ytnpdiw41p1g/3PS0of8HZirArj
ZLJqnc6i9M1WqyMSAF1TigSGZ8709G9a+BA/kZxnedpC+CQF5RklXZIptskZfXtL
M9ILuZbIViCSvU7jgmhQQE9qXWJ2GgPJoG8B/oDrpHsoMm8slYgWK5KUCAQNOlCt
nKeLNfXI5UX/URHbZBYnelCNabTfxjLeoRLOFcgCiPk0o6+Hvo8reMxwsgnUlgKS
TegB/1pIFLLrDhSVVm+GGL43d8byq64H29Td+RdDdOpfR9K6wK2+ER0KNiKW9ceZ
VE1YqNc3WUytqHk2Id0c1kjZaSJjzpvj22J/rebKEW6GNGesZ5EHQ1TcLGNiwFSL
FSTyk5IaqdtKvCHBhnrs79PBlNGVw0dV7NynbTYfGYT5SvzGYIliglLGtYzR+ycr
BvMtl6VhMegelz/VmtNKTZ2Sf0BS2E6dDf0LtbK0UuwaN01BZ2gN7FgJtu1L2ANo
KJkdCKdFCjP5QuyWlVKXgJ5/d/dfwGZ9MTMmS5szveYFl8zDztsEWX2S0oPVaTxa
4M+Igxt9psFeRHoGucwoLH7xk9+tDnw7TRRvSriZAAM35W9doqhHsjj2PttDnIum
6P0WWZPtq+Q/enyBPv6xGcmMCqt6P0icRDGFbRvjc7YxN3Yfpi8rkZRlW/xlJ30t
8AmQ6UlGUzj9PgmAYKuEWNCKL2679UuD/xh3mEBOgdyuwEMO09XDebcgJg+eXLiD
+wEvHalz5cuNCqauA4fiFw==
`protect END_PROTECTED
