`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zqis2lFeP5R1C2P+8WB6mwuityD1rtVqn7o3zANFR5yy+ZrzOP70jyonRFAMyJ99
z3B9uEWqRkbU+TPBhrXZNZ73ntsvIZwib2ljQSHSXMlCYgDc/pprBC3OfwpdfsPh
Pvky5keKaLrhCT4jMer945BYBrRdKjEG40u1JokMJDrz0BALhU/0qJKfLbXKvxzs
6rVMkRVM2rMXv8BnOKfMrvEINDwAr8fed0P92bYvvIYJwNdjQctmhO3Id18n1+ZW
X/qmFVKCF9bJKxIWD6kpK9MnBW2sc3Qx0aHbH5PgS2GDrjCgqwW39YuceJDufR9q
++FU2oA8WptQM0N9vQUTxAqM5CJu0rxMYnmko4ojFztsVHVdhm7aK2Ud13rNLaI5
DnMPHoWcJFuuYwU8s6G4EE8Nr0faqWFZQdlaXwx55sSH4fqgn2tBKVoTcGpnawWQ
EAMroh8q4c8q5BhbcuCACDDoY0xeLzD89M2L7cYEGyLxEnPfexLBG72ty8mnRAA1
5QLv82CnRDY3hYryMqSaVvmZgwwqZhn/AjTHrV4hFPDT0LeF6K2UDvyXD/BMXrzm
sjacdapYnui6UErrfFdO33sV5tIb5l8c+0f5XzbY5u6yA6PyIWhuYJ3Ixlq8CG4O
q8JRpVs+wAyc+lU4lZjNwYQQX1hxNr6mCVBlxVODjKqY8Yd/KD41eWUWYFG2GRaI
jkYiZZHOilP15SjYnOQ007KjWU9MSHYrtzZVNg4S4WlvdMLrfUv7QH0T7YG37WIA
fCU4sPdqoABQa7A+20mO04GDkEsVfPP04Q8WbPxcIJtutMYt1D+dbL10vI/NRVvJ
Wg3VN7qxXc83KYQ7XYjZoyTtFerSjA+s4YGu2NxKxVYyL0R/TgVWFwuRp08PYRrT
6lxZlCZNtYeziTfiEE7+nxICKmX6e4U+VJby8KEZkn51PBjmvLHwlSrwmVMjYGyG
VGS1QJNBi4tqoPDfg7qzzrP5prwuCox2L0sImEK87GowkepTIJa2HFsLxKM9GdVo
BG8fQLvJFWOJFC/fbP3YYu9VJs/kJHDQ3YhqWyjseWdDwcc0qxHSvFgaOS0Bc/4F
SQsJH7OBI15F1HTsPPpZFibb+KVBLzIGSIXLstHIP5VCJgzUX9cEsYfVRvtL1ys1
V2Iw3CwVfuHXxSLEilS58FruaRL+8xyjOjVJANRZdVcp6uWWe3zZfZZNhQPiTfjq
S6YgJ2IqPuntnrN1Z8ps+6D/U5AKM4vV+7eUXDsaTK/dzacKUS73kjpoq4uPsBes
4b3SRyJ/V86XbP3qjiOBZ2ePoZk8jwMPLozxFNN1+QplsvQtsecNHbgLjzQyIxn2
eVgJ6hP1JR7mkJ2tny7EFvshQU7vTZiCr5zYiVF10ZWRP9ndwyUijrVRp/xnDpMq
Ts3O8K3Fh/AL7K5P2VZSeusgxKHJiRXCwIT5N9u2XtYeLQpxyetpGzsus/Ob35oU
y7Mom+bcDz8XQ4PkJgSEFYFzrb4CJM8J0kTYenPVXkiy0eXbys6ESHHk/q2TP7Mc
Yey8e7nw0r5ga6/TciYTL3cZ3a078gH7ss53Ce8m5d3xbxKJiM7ZDkq8BWDWGmSN
PVTQ3AdGmwcx+9Hzu1wPbP7/HD/pasCXEL0qRCJbA9X6g6eQjInoUFmRNoh373DU
4xU61PLiMfQOQIG+yoWRjp8XB035XtA+oo+cMEgEmEfu22ArME1kGPaBrkZjLaUs
nu+sLNbKxNMOO3PlCKDpRP/0KUdt1AXG19EqOVoTYEkOMskrZf7iy1qRloR6mV7+
n7enBtWsBml7WwEVrbKriTLx90vKpEU8oiLvWbhIc8gBZwFhrOKaYBi3TE6j73/x
kdBTpeHJI+J8rktExdyWlj3d8preexqWfRek1tWHhjA3w4FST0kIHuqW9kM9I2Kc
rZxjeA5AjGkLPiNASoT30eyT/JCAUFuVN97wTqCTzJOk8Tx8LKHZw3DCfSFtcs4s
+IFtA8asH+4vos6tOBxbSEYzY/7dZIsZKA6etpOhsRtT4jGSc35qWKKR7vjvcwZT
v+feqGlWPUo9X0QjP51rDzA/48UsDCM6/MKZ/ku37fKNvFpg11/m3WAxRU/htIB1
DoBMslxIBRKr9gwlyIEATA3xiwZRvxSTn7Zl1AZYuVvsCxAx/wDGqmlCS3Q1JAXk
/NQACjm424qyeKQtkXoLQJ1E9zbLoUpplQKW8NFy0+liMeJ5y/Qj57a8/zj1ByCr
PpPxk+iQUUl0MRGELRLXxkVsT+/J+zSFN0O8Fr0q/O0ttoP1TmYZZC/K70K1430c
+qm3ascm5/I3lorv4iqOhCR72c+WCnXnYLMpfQz7xIXCmCV0iRXYxB7VNxb4hmUe
h097nQohKNPPG3UQr2v7P8OhmNw0DE6MVoJjNFT34cHiNQ9XeYMw+Cswahb2O8qR
PXkkPVB8rXHRI+3iUsXA7gS5YMcCFdJbOpFMkGQhApLZjvaM4MEKIQLNRDRVZ+0K
PUClDOImMP1RvYfx81ue0UUDId/43j65YPpHZwcH3zIrFRfq20127oGBoiv/NMOE
nb/LYF10hex8Vlit77pa9HNRxIG9quNvyd+15U2kTS4OHVlqtwdoaQs4V5v9Jzp/
UC69y0kAN1FcXAhrZ5aJKmD4zfsM7WkPhjXgnRIG373YmaUa7VkYN42wvmsrKw/3
8BfNXiYVKtljmWQpXOSODrYVOJzWh3CllFykH8TRcezclOUyDnXe3R01ZuFakhIf
rofb1Jp48HVZ9rqHHIAxPv1vy3swZNSP7clX1HBLTATaDXmtArMEDWQr2v5La45t
T2a4cdxGuFTvM+XhhBG/TwYGcMOPNCx4K+vWxdws8OfliPz3mkgPva1DEFjUx9pZ
0BK/qvVEYJbFynRzsyrfod9/JAsuirqKP98eDE6P25R7ymlHCdGB23UHWQG2QTFE
LPz+W/el0aXR/HtNENL9YjgF10c6alVeRXsTmzXSEwA/OnDG0+yWx2DmAUwb85Y0
YKYKvF58Yy1CKGzdO+2lkS517rU+hqfW9UCf6fUF+Mq/lfJqru3+xe5ipl5JZuCR
+SWCIO7ySvmlgRJLilywkbSY2dwJbXg1cYiVLeD+vYQNJjhPgMY119Kl8M6NuA48
g7uQUfIwwWG/sJ0Hy7okmu8epVfVI/53uQnpOJ7dqH+yz6jCWlPMSZZrODrjhW+B
3qxQNhNno51+CvSJTYxB1gusPytFvjQ2MnUMjRvjs0Q=
`protect END_PROTECTED
