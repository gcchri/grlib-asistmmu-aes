`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XsxUhBXC/qvcB+pejEz4p3uIEZtYE3d4SgD6PocYfXzEZZlLzv9slZQpklwk297W
ptHJKFP/tKjL8+ZqlHRmIpwJeZZgZ/VAaT85GLnsNm1API3jn6W6Pf0dNUMzs1A1
yDYuiYgr+xOePnmO285EkjcH8D07FCkf/u1h9V5UHWkV7zaH+Mh2nbTMy7sNEYVr
QcjT/3diIT+Vmq96WEZ3jxhYUnErCoMl39huCe8O3FvmFBEbMS6Y5HcK/Tp1MGru
lWgbzgtOGEItAEcKacwLah9/iwXKOCFgV31Ex1IzPOByd5CjCls64tQjW7P3mKOs
Utl4bmvq32SViaHWoHdtCyu+jsk78xxPWRppLtPyonPvtsrlFuFJPJs9ZvQZmPdh
q9GX5xk7HrylSHTjXrYVGg==
`protect END_PROTECTED
