`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+qasZEnONV8mCUv/wVQs3409f+IK2QZg982ZtSOC+RkIZEvMmSt7+ZRqchrFjiYp
Vjwp2K433kKfb+ZCv42ucvZLVDzgDSRL9uOb1kXLpWAkweyG9anmway7bmW35c5k
0Z56oFnFL3TgGqwwBsBGJFFKA28npigzWvn90y6eKGmcHVIWPAxvdVDX964eRfjr
VuoOw3JcEclOjhJfkezz7B64cwGfgtldPGwccSlT6y8UGoH6sgKIfPTMFoe/qtYZ
wzoV96lVQll6jecgi3lJaQ==
`protect END_PROTECTED
