`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qilUm/ufX0BgGZtbpY5zjNDwhiaD70/5wAmLeVbj34n0U6vdJUor7VwZHLKCHNw
Kulvtsf4cH2RvmZeJx1VW02wjXl7SNdSZWLyhGgdJgm4FJPGlrVqmv25RFcunkZA
poJAERi/owLym/yfT0r+9FGG7KHsfVkke6tAhi2rIJkBEz9vo1c/S5c0Hu2i9mEM
ZNgDPq+5nC3RcL3OHlZl15Fi4B4TJvJzxu/v0h1Ln2tKCBAv4PgkQ6YvYuz7yqqv
9/eilFgnL3bBgxD7/2HQg+gNwPVBLjhzVihED4K42iRWuJL2mZ3uipq5tkjXCvhn
JqfLQWMLkh+fX4AzwyQPqHcRG2+3AwbWjn22MDx+KEi2qY23rZu32bajrWsYh6kt
q9rl4/Z1GQEfiFxvzSd5cfUGP27tmheuVDRkYkE/G+KNwOX80IjUz4KOgkzGw21a
iExi4gUt3rYNzf97h/ywIBcLTV3VPP+BIhp+ckNM40V4xYydPnvXdKxAqcrMMJfp
KHUrXk94/CTnosd94gQOJgSZm3JO2fVDNgnMg9aUn2KOwN0KWaNVf4cGYKszRTbX
+kxOkQmnm1y+gTvgFXcVasoV14SD963Oga2eBpnLTlDJhxfhkJ+IG8BjI0Lplvbw
8onC6JuJbHqQeI3OE8R+1Ommsadp1CmADnT6ppEBiA6bciZqBmJTv9SXG3nm71tB
oJ3o3qJWaFTxaNoEv1TUpOFx6rWp3uu8nn+6RueswFakERrdwOAefujjFx85CGbO
2hzhEsv5R1vItWSdTyKmB/AoYdbJgtvNIMjhq1Jjp7ObtC8uRt0KAj5PkC6fNMAE
`protect END_PROTECTED
