`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vH7R+D+T0TLn6N8XOJXavzcYBNpj9gnWcHP3+QKpc+SPQYnF+1YgYX6PZ0eYESA
4GKV1Dq9uHjl4s/USB6kBosI6gOX2yg0mZaBm4wPvqA+4nrrc/5OtkINZQp52JWy
PC5lPlUGrNDYJOgV3d+RcZUdyg3A1NXNsU1VfrFWB8gdBNsxx40MfP+bvTVSSYGq
P0u/bqD598he0fQBzsbgE2aV8q7nNbK6aXWMSXwqAKJo5hCekhRMnQfD722K1GLK
V1wyvO0SU32gcVNU65kvTJnmddwyVDjFPo256XF2ffIROk9xV/yuErF0XWy1YHu5
lBKhb5L48Vmh1wba7t/aH2PH296IijWcbyZ9mQuSGhS8Ni7g7CPMBX++BAOi1bXN
gTCbl2H39ZhuHvDDvxyenKv6Ot+mioS72N1qOIaH8nyLDjepUV8zKTOj0P0xPM9X
v9l7efxtTxLxppIw91LuJSH3lNirpOq2YAtfxCZgOrsd//gSUagjKnqMlA0kqwbW
hX44DveHBm/G8by9ehRHKdPTa2eGyeYGemLAXebhd30YrOVqV8CYOkJquGJLDiS5
+2HPIFENNrqQkWFXDC0mwoJ2LfyBWp7+AFIRxoUxTgpB0U07ZyrGPVsvuk0XyqXQ
VsRUpyKwnnVoEfzDR6/KL/XaBOLQ0lSr5gb0d+gZvRWivE3W4m7CGVKAJ+SF3/c3
5ohS86czIkOjpP/ref4jpqPtI2/+8TQGSNlA1+YrrDamI2Loek1abPEZ//3KlXTi
JFBqA8RrzxSrG3TtCOiTe4BTa9R/8oX7Ol+U8008wbDHXsBHsxUTkhGL1/OEa500
s6LrzzZri9RCq5gulOM1LBU2qQ9sGYxhxSUx7/BfOlZ3pQ1LVLewBDPVCfwUBRcI
cZ9F/I8D1L+MAzFQQbXMo1R8Qgbwl96NICcfpZpiG31VERPGbjP1z8EZ1EWqzd4/
Uji/DgzSlauAndnZjPOA47wuv3dTGSuMpEglykzJ05hCe2wcqo8s8+3blPGUUwDi
twAKEAahKkL0IEfl3OnhBGihNx+nD/otriyDgp8elUVs2eAaelFvpfmfBT7hI3K4
BlhW95UwqQ03b6AMvnPDw92KC430huoRZiiGdCoXxtirsfIqOFd5KsTmj0sS4Rnt
oYCLNJnYUtBQkZ9PI/1pWYM2uZDuYS4V2lCWZ/dkhnz5DiXvxTNVK2hLxZbtrHsV
c538tZOv6yt38UFaLJzjDM0tSyEPx2lyXIDWs633gnFKRsE0I5TFgBU/igmRfutB
`protect END_PROTECTED
