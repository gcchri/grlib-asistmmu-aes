`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6ysKyziA3p9Dv4udF1+9gFk/U6F3NdTfmrbUqnNlk9fGUo0z+LDIYNHPGSdmheK
Rwp0AjqHNqfPXXtkkV215ltjDeYVhN99fcLzE9fHtPO6Ero5aFHPdW6Pas5p6SSp
DlVPoP42VCQr5FygxNHpMWXdEQ5EKgyf//c3JclvGjQgDnwzkULxhZ3bV8fceXSV
B6Qn9fvBbW5zq1oFbGBmXQaRrCcxpNpn2+aJYorLph/UEelZyQIkyebBDAKELUvj
Xx9bJPa3lOZSfhmtfs3idRzuL/X5YbW+mSiLVpuMre2xIpe6gLXL1r+umPXs/dwA
Jl8cAvsV/I0u+wN6W2Cl6MGambSpRIVq+TM1Wo9dfZZmu5KZXh984Q3y1eBi6Svs
w6cfNhvh4YbsC75X1vRcHVrviqij3nyFxso0YdW000mE7rPhDMtlpQL1VH/1CAnq
aBTTUttt4b0ts6fSd3oV3twGMRkR/V8rKcUZXUQVMMZCkTaTmkGCQ+8VSnXtvIa/
n/Y45FE7S4fOC0At45g2WoY6SZfksgdfxIfT8daj6CNIK3lICbqMJN4OxnYMyDKO
BZiLC6xvBnKilR/k8WBJ2Bbjsw5VYY6yAj7WYLJ+CQh2P8E/6BgYZlIqmzQ0saLt
h7emznt4r5zNYBx/NXKwoes3UIFeKsOvIHD9yPlR0C1drxh3zjAKvP1EA1PNb4nx
aQvCXl+K+VFnSd+/ns+sy0DU4vzqYRLdaw4OzcOHGwG0cu01xLmXi8mIW0o9KDJ8
lQSGt6gdQu8Oq60rJlRaXqV+vM9SzAAEZiGIlWa8Uayofzw0zGZ3jwsC8KPo6Q9c
lNkf3dowwNJFN9n5HwdAnoFwqSmbU08DOjlB1BQrLF6t0BzZ/yGFEfKq/Ri0AIv6
Xa9aj/FyyfJ5+UdIS+ySjFCL32CaGuMZyreKtN2t1aKbUJxlzVngh5ZgDuipBEBT
tRTIX4Ba5BLmTQouMziTso7H8DqZuM755WOdk3Fl94gVBAlwZ0QG0xi7itxE+fbT
HMIHJMRR0rvOpLQQuhmaGseb1GrjNI146GASwEYdGbIFUqEKS3whqxjal52QPpwk
aQC216deNrz16J6KegGfEOTVID3zL6GAzW3YwhetMIagGoH/Md1pov5n8gXp0HE4
gzaqv/O+yOmcaSj6kVEurbV3cSETrK00llJ7nn9B+RM9iutsX4+TfOOXbR+F4WnK
VpN8vqnORaI4wXsomn1kQ52Z+i9Lu0heTErTZUOimPtDOZWFtCkiamP2XJOejid7
`protect END_PROTECTED
