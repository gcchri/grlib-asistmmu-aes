`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NvxUapojKyozb+UYUSPoqtov7XNdLng5YWEfbu951E+f3TlUaPj+/rcgxLsmlMfN
Ukn7+5UZaL2Opva2wWQMgnDSjAdcqXcfv2D9V3LtH/LKmC01lDE6R8UBJkn5spNR
ymDYxJywwWCwmix9Hdccq+Ne2uXzynsPamgN/CzlpLv7YALLxU2KO/1fPwPp91cS
STTZOOVsw4rDnQSEC2L66LS+mYSOwPw9OLa6j0uMW+EwOzpCqM5oN1FQZR71A8yK
MoFvN+VLduj87K8qv04fjqq17DaZSDzDt1nDoxkckB4WCeAhAFMG2pmL8HxF3Aev
keES+rtBRdvE86QadR9pRb93sY3IGwB1jJMyPUUQYkxkrRYX/WU/TcjgStgJxORF
J6xczku7znSK2wgKR1jhaBPrywQyUA6rPzFgYwFLJ0wdS4XfeULRWRRZeokgtTaI
`protect END_PROTECTED
