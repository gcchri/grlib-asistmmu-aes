`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HTKxuzPKqNbgP0l8atHLDoSfl28D88eSDdayyvYQOn2GTUx4etxk1dWErgweuPA0
WIBds58dPVSzGJEg+KaNWQiQOjMaPSwW+EFldq53aZR5BJ6G4OJhUt72Qn3DwN/T
MewAtiJAXY/lBqPRPzH2uhYuKuALFaFwF5w+yg+72T3Pe5fRLXdqKJxffkpOAPxa
yKCuq1lFn2oDlhjS310Y5chNPQCQJRjumEw3de9PDvELPU+gbNOKeUZErpaHO5Rn
XG1iESuFF9TubFvqa6VL6hbzA0cUkvlOFhu1K1Vj1DQzzFb/rmBPvfoEt3nnlYNq
cToz1iTnCNbRgm97h2NGidrnVqmwU7Vs8/uvO+/s7G8/GpRTP4QVFoFBPFJA7aBy
i7dIGdd6l/7FcaypXgpG0w==
`protect END_PROTECTED
