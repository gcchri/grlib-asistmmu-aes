`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SzKU8Mvp2KqKbQwWL6JyqOjDvpAUXSsydcPQrAmUsR/b/ylCRq+HfYqWZtiZDiFJ
TbiXWvoFbZ/f35ZApvYJraCOuhf033mFCUYevyzS27BdZgRTzSPcBIqI1ycGtMIM
oNFrH4psQLUcLyos4Pr/Ei6n353r4D6J/8A8/GHZNaxDjC0fb5SpXawlgfkfsgT7
D8zL6J6msPcPYuikhNeb9s8IF4kBCHVUdidXd3Nrzjt4VzOp4Ae7Rk9ko7nOZ92p
PbIgl17yMXIP71GCj4DLZoN/Np+kdTtYp4QswzZYgQQ3fExtYcWQ8nI06/0nr7Db
EWRqstmxEQuXczKXokJR5ateqdP2g7lQ84Qwa0f1Ll78TX0PQAd/iemyttGrNCBb
qlJ0O/4gKp4yOyApYNP1AxkV4ggAw4H6anfyyjz7yPcVlqoZhhAw2dJ7zDCtjMaa
rNMVt6IwqICvaJaSA05LFiMJgA8tIzIQgZ7ptESnlQgs1BwMovRFteLAtW7wxdLP
gQu3SLaPdCdZ/l1J1Aqf3g==
`protect END_PROTECTED
