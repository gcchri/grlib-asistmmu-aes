`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+0QTY/9B55N3ESqiCXeHA0XtwQpfLRB2X9gUatYYRmp3WHqUbX3s9bGbLg+Xt6Kn
uJ1GS+VjpAW23xiuwTZLrTb+bj00PNVNBQ2pVzK4pA46GzS2r4s3661C2fF7bzmg
wtZ35zbIy2BOXWmWEAcv5rSZLwplXY4BSQA9kxGBe61ePkIq6fVotntba4r+jiFp
Dyc2EY8XK6goVnmRDp+RDOFfsN1Bx0YWzJG8+Hg/Tr5sdJ1NqARpAuQkq15i+puQ
UaK0+yHTruwV+mr5ZWdd4ObkBDacwvEQwCGDkSXIjiPwAZWbgjXNV3XqXgZCcX2E
oUyC1ow4juvAT61dx1xL9yR4K+O9zrrLn8zJTxB+sWctkRX9bkc5HeZmKT+hXaJI
LyV66oNxhd9OBlbiCmrVUgQ6Mc8KJSaHcLYIAkZR/pgOVy88G7assTvuZ2du5qYD
WyxwyT698+gJpXqPXO93UsVTs6tLpNj+UoV81q83TUzMZkSvlgX6/i/NyY0jPiCH
`protect END_PROTECTED
