`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1h+JSVkaf0cMCKh9A3hNxv7BB/3HU/mqw+Hnz8RwI0Pgu99NbvePMoFO2mcuO6oy
9maRZZBBIKcnn7Qti+LWVbhnCQ900O7gj0wQyWPTd4pvkHhlMbblytYvE31ph8KB
yn/Bkpdnd4oyKCV18jX+rsfT2XLf4NtlR94fEJPtAxwiNEJ/zgZ5DuAUT7bv3CCN
LgtEGcflgf9gp6YMSg076aWnXbDmT2Z+YyStyiF8BPtv7Q6jP8wRmDHhuB/IGrgl
fyewMow50y9JlXQeEBgUhhCp3l7GmJUNTM/Y4orjV8eFKI+8SvAsc7c0kWTF+Vhe
PqYl/uLcvJLfVrgqTIh0X8It2oJLX3wmBhkHor+dIw4N6mR609QM4DPThLBR87Sz
AKwaSHqbbrPlvympgS187HAg0Z47gVmX/3WRlkFgvu5s8U5tH7q9wWZ3UxGDRbgb
brDVby7ZyyEqqVWFf1kVo+oQuArixcpwohE1vMjTS3ce7tWFzEI8TKLWPGucIqjZ
svwBweiEzMWFRlnXYuLFAkit7zNXyQ5gSG61b50N4ebhfA13SrBE55XQWvhFD4gK
DTeQHSJlgfjm5uvQUDU+4pqFKGuoknWdfHkmnF7vSY4xTiIiPYdD2BvQfjSylqBI
Cj2cfedkG5QB3KmjFl5t/1Nwk+1sfVe5P3ywsgCeMTVtW0qD+JM8MlLkMlAwNndq
ST34J8uiUotdI38zlLb0UFa/6+gh/VXIR47GunqgCnZ8nrQjkvzani9Dh3W6BO3b
1geC30Km7AOQ/QCB6I/LUKmvBpPcSt9m/CdweQLVQ+JMvwgJKwvY0qxD2LRDmRyi
5mMVhXcLJWjjSXUKEuqk0aujtVur7OdbSktT/teuhJfBmJzdZoCIlt48Iy0QjegJ
FQfphZB63ZoawN2QtUe73pP9xn+l3O9yoYqsUE4CBObiqfAOqf/wkoojfjUsldYy
F4REB+u6FU+EXofAuVjybROcazZiocyEK0RLbx7uidU1f+YOZhHNoX8XZDTfOesc
t4LXOgLUE9DXSPNkTyW8/FDsBdayOr5DFA/dWgYpIisC6EG7+k+JiPGUMkwyf2t3
k/74iCX+K2gW7gVaMBvr1cKUlQCzKAUr/cz1CC6qOgofisTkTvSTLeClVNlDYftf
Y9V3aRXi9hyOyF18MwxbhZGQ/LkojwFBhRRTI5NVX6Tf2Fai0ICil6iuKndI5bUL
2LENhvFQSeQtLGc5fQ3WzFDNXt1iKl0f6vNduAnlfMKjSXTqR3a4g+Lbs3W87fLI
SiCFnBRju7O7XHjpSIs3bTzHddeawTLdujPqcuoh64Ql2eowKrmP36sJ/xa/9rXy
ZSpjpWEkuywmnfhCqYZBIxcYOjrBNKSYrAJ0m77JumGrBP9fkalrEJeEbqpuhXwN
+T01WwGdsLp6zjj6ySUlDkd10UqT5kR7qxe7He8/7hdFIQawGmWL1nQtLswBidNu
GvNwvdDZ07Iu8CFY+3dWwU+olLGpzXbltyW1FeuvRUfKSqni7scur9kxci1TwH1f
gGtkQL5+p8MrnEtG42Jhtxbn+ikTWKfSbMnNH49E0oDZ9zDuaMbP3R2c3knv9a0h
zjEM9ri/S1d9ewZXKsRIRJRmC06jlIjcOBwMHhCqtqTbfTqjR4lwd+P/udPNRWsR
YpROCR5PaU9/UgP4Atbzo/pf56JyP9yVyv/nxUDmsU1qWAxKIILQ3cfliF/+z8Sz
UMHNXoGK3b6N9bd14UG3GlZC+IVJF8fUGRx0Qo8GQWiulpB+SXN546gOID9xr6AY
v5J13rGktM3GkeDYlNwb3i2B+WExQfVvFd1WxSM46FDwHSePUupLLauGeFmFTAQp
T5KLTLD6dGNpmvE5Vgw2FYggH7Bew04ua18rbA96kNtoB/RJyNKWEIxR1temuiQD
KHE0/J8EIR6f3bSja2SpW/9xp9B36C7CQOyVjq4/IVYfqU5kJx13FSawG6abXprA
DEmBtzTtncDOaHxOWfRpXzoN7FF+z+lBQ0Gh/1AoRt94fkI92mKufFUutp1d1LRD
v8/G2ZtU4B7YRv5ludKK25o+pX2jXWBgwWpxvkaV2m+4Z7B9hNpxJDVEYaCNjm1n
wb/rLJHZr+mB+Nd247JcuWd+RiHsG4fWKeG4eOy48KCqAzyEZXkh2RARDwl2Ayqp
qQ98Js2KBKmSek8Wjs2S6ZEB2ITjkHqokgppHUdSWi0rQkiw2fRmzUQXEXvYZyN6
uARimXGbCwWqyKDdcI9H6Vp65SQ2DqNorqGd8Eq+aGh0KJbFksPdbFVPFXqf7nDx
xGSx62vT93h2XSUuIzSDEbNyHRJ2EEYtP66Uq4/trs2kXSAO2qklkfPZzAjY7dhz
m33BhPUGoKETbL7f9g65yvaPaKBO52nik0xw6S3bZJxXYd4hQT2zK51XFOHU3gC9
vSOUSQscorAW9PVHxLs17LvTEJ+zr5raQUry7fXuZsBrzYQKb621Ry9Xqfgw7iyN
EulcFcyOi/GIIz47swWRcMe0Tfi2LhLrb2HelrApyMNfXF8vXQU3y3PjtNkoS0sp
2BoHQoD8iNsZsQIPDuorvaGNQkIDyiVAQWSFN8I7R870n2e8PG0DNxh9gLnHjYSE
z3y3qE0lO/SB2o2+vPcTDOTcdDVOz/mkh5qQllU6sj/GGNigCMsql98T7HVJYSq9
PCd934JeAQDDXzxYcTwwRFRUErvNOl4SaXYPYh6b21wL0ZG+V+lPhPUz6yEa1NI6
ryrpTRPZsO5TzrY8sd8r/qT9LRtSyPr7aT6NlMLWrLO3lx3KgWXnJ12JalwgBA/p
cLr55OZTPbUHfDHqL6mCpjXV8clHQ7vM36lc4+tOmu0TV2s+mY2kVhBS9DWL3Cg9
3y6F2oOAy2u5RPXZw6TQR5tVjiMFl8BW3CbqlHA1jx01tA+SSvbKYank308LX17+
rlyBooyHdL6+bLgmNEeXjcaYV5qIwOApNwJDC15enBpuYxI1tBVpCkJPwmqoZ4pm
`protect END_PROTECTED
