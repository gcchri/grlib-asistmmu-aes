`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9dIUPn5/zsHO2HTPA3whqqgjypwz3yf+/qN1SqvON7FAj1ub9lZMmDspaBd717iV
1wpLDp5lPNNM5sxoY4bLG1TOJKvsOKzdkKzcjUZAMg0zltjw4zqJA0cdq2DglnYp
U8J4T6n+UE0XzYfkxH6dbgZSaXfgZW+iX0JKRwtl2WDwbun+aEaUdvCW8WkxpQGs
FuFD0TCdMGf71YtR6nqcOE22+dUL/ttYmdnEe23JEQXHpIjcgdb/lsSV7DRoAjQC
T550ptjrhdzg7I7RIQDp0Yy2IRd2QEG5En4tW+xKbaHLuXsZzSDC3QU91cfAKEVb
ByeHMdGxFAUL4udGDPkST9qigF17+6eq7S5PTG/8dM5bKbmmETsW29p7zMFuHV0R
4e0iYUvi+NkB+wf0jHyQ+Z3Qv+4CpNET9F7Rpx1Y1m1aNqwXFg9YS7Yvsvf1iTeO
qRsyYhL/Nw0PwB8SIn9MMNEQkF4FfoCvJF+gE1fe0/jTP4DqVGiSQUoeonu6N08C
LxuQ9cuYtEe1v2nt6ylM145WEoy5ipypw15P58CguMpGfqbimAsIpnR1nW0arYrU
6EAeE+kvn9W5TUieXIf2YPWqpjC5t+S78K/5BqbdA/1Ufs8+6cvGrYfrYPT6J+cb
Kn/3IfIPNftBBprjdpiAQg==
`protect END_PROTECTED
