`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohkq/7UVHPh9PXvKBwkadxN6Fog/pU16xaj03Gje47JCUCVgWQQOPdtml1Rm2kfh
TvF6w3isgj52zXWN2J4hUCPDizHBZgZoICuXAL0nSK67J8X+EtGAk3q0d9ZHxQcb
cf/NcE9TshFgCG174d26U6YuGGJm8L/ntwuSP+xJaP8/sloMfS8wQuhuJRMV32Zy
bhwI4acvBS1XPH+pF7Lw3TinnxZ5wlhQJO1K+sNOpQ9Rt/YWIpRY8qJeWyj9tfON
VKtG5AyqNOwqCx/6G4vkOg==
`protect END_PROTECTED
