`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hAEUPKD3FWmqdzn9/sSE6485y+tuORoXw+mjbmQv/Bwm+wMuUEo6EXgoQ3uBIjrF
YBHi8KXkvCxS6NOJldhWc+NOaHhb3RpzoHLYSGGWsX0OfvzQO40Et9yMSqBMijxJ
WNARs3IXhyJY8DjFjjxW34TIVRo4pV+Me+hJUdTDAPaUso5DyU6ICKNFPxlnm8bX
dSrNxRlazPniEqZiuLcEcu3gj6aaKokMs/uA5rDRUUCgMpf0OuZNwukqyS83dN/t
nZCdAQRHCJmS8kj62jENTGuftyHZVH17gGCds2bayu/46ReT1VLmzTpp5n9feJCx
cDZ8w9pAZioD6RfkDZJ/VqXMmWaMmOszGv8/O6rs9li0N9M6Lh/GDws0A9Pd5ZS4
OZ57xk0TihSVnFmOZs8FBnwACaSU1wf839grm94SdPd7sjCgJrWoBQelgLjEqkOJ
lnmQqKuzb2qSN81ljIWhODzBNz5OqK0PQv9Q+a9rDw2qJ3x8bv2VBJiFz+GYssNP
qaTrMrvm28+UYnTK2TmQJrqlOfu90/ZU/r9mxDr0pG6JHddJwsGjB7H629MdAoJh
Uf2kcYq3/dUenejPF3Fs6U7PgFAsGWDQwUoUCv9JPa/Jx8hRFYXbrUrD9bJHh0+Y
endElfPHn/jmA+Y4+lnTmQ==
`protect END_PROTECTED
