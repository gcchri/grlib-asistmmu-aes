`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oqb47xNhczXcAgBYhJaTsOLxbHvd5t4ohl1WwUm7umg/2AoEU/McpFMFFuEw0/0+
vwYLD3Cw1ZOqLnt03OdN5hHhSw5wZ3nKYw/dd/7WcCVYsFzZ8pu/zpQR2FxFqfYs
kf3RTW6iA88FG8iOoub64N4coBYsL5SfjBPb+AEwbz0BYLwP0W4MAb66QiykwzFQ
osAoDH90YUb0WdBuLgRlVxQROcxlkJA+CLV+5j8fIIgdtfzUTXzkma3kSOO0Fxf6
AcDFJ3SGANd7VOImyVUJO01sOUimUzrRtMw54rPk24X2ylbcoutMMK0YB39RIcVK
zg9/1pnzXeB6fwCgrW690/j+stQUoa1JOGFkHlMZxXZBJu+jM39awk8d6LUVnHh2
LdE/z8LWcJY2EPWeQmi5kTZIjGhwPsnoVziYWX05IgU/v1atfXzb7/gXQsTopWEt
FR0ZzOlG9+siym/buUeOTphAe/Zdi7oaBjtI7lizAt8CG21tGGuTGod2G7ShlxjF
D8mLcM2pKZTM14vQ22z2n1wXoa8+HWj+CDVdRxAL99SCR8mMAHh5bv+JqZ26LSJh
Ob1Lyk51NVP1Sc16/eh8MTK4yaywRxUCqoa2iGcNpeCk052BodtuVqklcyRxUtne
rkC78OdUNYebUutQajpp57170lvBqqck0SPZf2Nm9qTiPnm9Xon7jUNSS6laQAZG
+M2IFxeEtHVrnAi5cIvYuNkVWSuSPdMnzL2qP1BoJ4zM8qI813mD1awskbzCOSm4
x5L9tUbnA0TgOnCuQj54hX5AoCJfiNR9PgACXPxwBsaLuEyHJ29NAoDKUhm0SC3+
E0deOOiirI7/TlC6WL8Pp5oZ0YrvYZ1Y7IaeOZppw/XoBpXnpy+42oKeyzeCErLl
+ipWpc4XcY190QsS6iPX4VSQbZZYlOPjdsUyIrA0NbAordeMu5sFWZ7Q7ty/cPgz
mgIMAx/Fgduk6wBrArF/PyZWCQq7luyvWXfv3TEJZxt66UOUgQT3S71m9XdMGov9
44k49eBbENcyWFwsimPc0qSLMvpJKTo1fUc2MuwNKd7Grontk/4b25WW4wa701N5
UQrm03naQjFKwgChm95CPPLsMCfiLp1EjZp4ViJTc9gEH0i59tuI6mhSUk94USkF
cLPPGLjvJzSVdEmV8TFD/6Tb168WyL6Rc1XR4MOqr0DZ17y5gV0uW+lbufhVAaBK
ecXwI0Lz6Yg/XNWBiJeuQmM04lii4X79w1nriH3Ol99/nIh2Jm7rT4XB+jt6Cnmw
LdkEvgN6WgTrOqkY7uXn+LQA1xpaZuUMkP/2I4A8RfqOzz4VPc5B4z16S6tzEJet
6tbo6givB495Xjzwuuha3wYOSffNA5Tp66shvsIXT1lHdNcVfphwfrv0YWC0Nx55
Q9RL2HWO8dwVPZTHBEYd02/0sVo6/5FpRt92nhq9GAGMZx1MVIS071GgRhoGbpHR
/WyzT8A/RZG+zHp8PPs2oaePMV0UbyFmyEBDPMGCds4pzrhbPPvpSvs0pSvfElTR
mvWUY3Z9b1VBd52ppUG3AaDqxlPjMv20Q/PtdDtHAkMHW9zC77pFAv2RYCxzA6LY
q36DTg4LbqYXMBjFyXJokQWBb7xpZnhTuSr7sqjM5VdsYPewEpymszrB6jiKG+li
YcBI1rpZfHLdhrmaBVCgTY/SHbSujm1YCiiaht5Ub4/blyPrR4bR6oELT7EKM1UR
pIGWZu4L0LPfhY2OqtbHYsUf1UsOM1wohFM+pU6+E8ruIvxZgvdB/e7JcNsS3Fa/
r0vQxkJFH7swQTL9DBvQ1bfcUy770qdwHo5jHjXU8vwIw1QeAzWVIoz3DAX9Vw4a
/dbRzIZz+yVG+ZFPnu1p32GVlf6dW/VnOkapAhz0E7netM5+LDV5mJkT0EWVYt+s
l/6LiNHYt6pxucbZBxR67VqFLfgySFYHSgt2hAOZb9t1dkWzsp4KdmxG0/slPXTI
+Njnx5hUmjqymbmqcBdYaYaaMSWQQukp7MbNhHbzAYPNm+9pzM4a/FZM03L+czXn
NL6YCGd+oqRldwo4cf8USGVl9Ls3w06K1wxwOgwjYqrV1tQxDOCzZKY+kJqH6+fJ
c31XVLaum64vB+zymzo4+bAJVPmMOTtQ0urBA2sR3oECNhVtTODydo5oD0j2k5Sb
mT8fo2+4ZqPJ8+tswF7XWv2ESssnQULcnuaApKDzqzs7YCNxCZQqzIN0HJRzGOmV
uQgCOUcgaPur+pKSkKqB0Gb2nCmSsU6dCbLkPU8Sq/9WI/oVMJAUNeFdvOkpVyKf
kn1tUmB1d4nYe4xwj+4wMq1+L/0RmVHuJySrxfjsiT0Vr3TBOnusip/w7++4nTXG
NxIdwoHQndJ0VhWRqEgLEOd/RAUuI8BwXjFZI4FTKCPYYSJo9ayc6n8G/pa9jhFF
lQNof5Dqb+Hj1S4T5poPY4hbkyv0QY79tw8fxnk2R/4Xl1k2/LNofiAd8wE0rjWv
FqdZF0i+poDHExA45n8/Oo0Lb2UWd3zsYLUfow16OOXrcC8J4Fv1ux+7nRLqLco/
fLqCY1MNCflAavBVrKGHYCRczeWz+vC1kbzz0r13egydvEdAjba7SdV7O68gf245
jfnQiO65OLvfzqPR2I+/cM8MUYbQe9lN5InWvXMw+f11o8oYpuPyQTbLCS06CZXs
AshDBu+ZecjUCsK8++TQm+v/qCcepzB5SH1Q922UxNgV1wxqom64x5tUqgaPnYCo
4pGjeud/Kgu1qF9pwc7Xaj0SBhMP6EIcPgHJ5reRCpegT35/iBtIGmDhoQpvS27+
+AArDoQWMm5hNNWz++dyZnqZqprIN3jicvGrTQiFSnuyVGeHM7NdWZC/mfkpnJCc
+k8d+cmYpZb1eX1gei95YcezMikJsiwQvhlGrB41LoSAv34lW2NQSsPdlVU0FWZn
nLP6Ysc0w66KK+2Fos3wGkyZlZxj+tWsXhRhqTaPPgYo3oTDDCht61syYUaUQUrl
eu5OcRH9U0tOwj0W5gX1TLMQeImfcsWddbqm86wEh28Kl0XgiZaw+Ph5xSbdfAI3
Ji/9x07ZygIQbQrFSmYL3SSJSmBjmN23sKmPeg9Dw6FCFWxdOkpsZ6qkt6rf9H9Q
s5arGpN3Q+p0tgmxHecczAp6LhrTSJJRKe+JX4eCShhjynSSs1Kxkly/k+UdeGg3
yeDW1+QzYcCIW+9HFcy+7ScqerWcMEvZW7YOlWDbepv4aH/Iu1K4HHHDCvJgqonV
KCUi223MSualE6Vj9pq5LODBkJELx4h0lPF7n9PyxERChRmwpL9CH50U9mNT2nju
3GwfVknezsxtVmjbmYOeX22UGpW24SN3ZI5NF0EAo4gqq0FcQIq0gGxxiAbY6Z9P
ZxrEUilzY9qmiCIToVK/DawpyYnAhW0rRwGz76iSIJUJmfx1TRQKPAj3kKUwOXwM
oPJl9XSLsy4+LOjX46U9C02nrLBRGsB7ZaoUY1e1wsosnNi/bGJ7nEFYMvi+xwt/
Gj55S+w65NUjWFRpHM8Jdyj4Xcoj97uiyxzkSqyoAyw0itNjVToOpJbnpzqAI0gc
re+yOOqMoU1c75EPCCVctInXyq+EYFy71ut0eA1nbu7dDYJwPgT0ZQ+IOhn36Wf5
Swp7IjcWEv85afP1XclrWhnXDTR/dnH6xSdDmDAQSTF+gFFulI890szAEzk3wjM4
079T6oCQMYFU41a8iCsS84e9FMI/dnECXLpi92Z9vS7Mm5BQxakQzA+OkyiDC4ER
LSXv7QiW6KkYlL6jvXq7q5UUBb/2T0suheQ+QTrbgvIjOUQrElpXQqFwujAsacHH
xH3ukV6ydMWxDljO0p2474aQb5MHhHYx2pYmPck4yialpyGt5D9rOjCqBLJRD6dF
dJIfp6Tfrn+tO8LXpXA7AJMuZRjRIBH1LJpO9ZtyidNmxVD4vCgX8bX6kczdX2YA
b6x9E4M/5XIkRzb2YZcTQ+954V5u/k6CZ7k7NTHfaU+OP9N7iIWM7t9aituEQ45P
OVYYx8sYzXiQwxBs/kFcnH2pl602FGwqQBY1AJ+1/0cKLITde/cIiQ8MazxpuYc5
oAMhF6NRmswuqXB8VWeoNkU7LU2pjbxDWfgQEKIKSaQOsb5LsFOO73tZuPoDMrMC
ioSyBXSOKlhS0UaZZY6hYRjYU0ZQpQbFBnTN9qLtJdELFyYEodqHZ5wthIYQyBuN
1RbkcIV1s6y1aPqcWaWUNy7yF53cgP3XqXqnso/YEhM0v2OrEj2A+PlcpTkrjdBM
zOAX5q+w1efq8qJqbue8N8iiNrcL2n82XAcDD07ktA5EB8sts/X1xJQ3Bu1oOl1h
5+BbENvjJlTb7fWf/gf1BXqIcS5FhXAFotaCkQ84Ttd4i6Z5La8J+HTpn2W9s+SY
mFXHSWQ5XLaC+cgRU9Rjs7USi3QN4DcOyCsVzg/m8apKZb1xQDYjFsupOmjfalDP
0H+rZAylZxsKIgFBQn1CAY5BFgvLv3H2JbrrLH98AEa/ropegXL93dlgoayb/vmu
bAicWC8MwNx8W//zU9S0r1vedlsLgK/KkhVRlre98BXb8hHCxIH5T+k2Tf7dsjbc
Rq39PYKh4+7nqVRgUe771cG76su0OCbIr/LJzSC8vWtVi8R9NSTOsha2KarUk0cn
6gqUR5ebOvI1xNWZsylhcnLaL7DB33h/rT1XByapTmRV90sSDGjkh0AMwwmjdoLH
zZaMOVtmrcr8Wq67r7H9PKtnDzpag6CWNcXM8jxkwM8Kcmi8sS0SFMIr93Z1jHqx
QAn7ZV24eHXTaHkvhL76SD+rapXYDDPo9AkNkH0CqK9SozQfSvCK/85fHZMqzCwr
fXLDleDFh+Ieb2x19+TKbclnUvQ8DMCA4+PncCOyA/w7nM3M/BVJ2kyYf+qg8gdV
nEIzu8cmIrsSCZ4dqK8eg20EZ2UAnjCqTcnvwEJLwmf+HA88Hz9njcqRBJaFJQ9j
qTP+pmi8POwu+EF1D5AM58smrtPYg752YdVlxmyxk02Vogj8nzysStTxtghJ8UDr
XOCD2dPgaEB2t1ZNzrz4pbjqAv6DB6Rvy0QOeCKOgTnHSrjx47aNBJkzphn4pMVi
hQaBJcZKdIf+wIyj06valZxDAv+Ou4dXue9XPMpcsU01lv6yLM/nVuK8F63SaBNy
EuVjyZWDol1fz2XV9LySEVs483PnpfOlICWyPVOjgwhPBAgh40dfuIn18+gHBIxY
y0fGaClIZ8RcWbggzETF6giySrORj/RuX2Q9GmHvN90I6ZJotcvX2kD9GpU1GWtU
wbDpvJgD9cxKRiq/ljBqMo8DsqobdavMeriZFwkuAf0eap3LO19Pb/IhN00v+dla
Hgd5tC/kzpuBCYnCojL41WNDYmlGiKmRcJuhJknC6nVWbQRdXq3HTeteDF7CZJWl
VtubnLmg35MH5h7PSAPpneC4/a+TasglUoCU6Qr5TPBzSZcMB4TkiG3QWs8q+vM4
/mh7xCjaRF1BgBPqUqCNDbhrt88N7kWzL0i4itSbiiHOQhfpazZ67/BvxKBr8+Iy
xkJxVx6m/g4BkyPhR6E+5mx/UYHejRgPV60ZQkFUeONW1hegUnuLbA/RAML/R7F6
I7zUM8R21Ho40d28usD//ZEDKTR693Uxmu5XZdtDT8vWUDicx7tqruTcSrQy2HJD
6jdn39AZtPLQJedGFtotlC//3fuaiOCZ3cB+/LERRDbn9ktbfJW5pCfb1I/wm8dF
sGguLW1W9ifgdQqDahKfqTKQuUucP7o/zZdBoLyKoMy7qJbxTptEOQsehEQ8fbH8
ea2ebFq4niJmmxJIl/48gOfj7my5FSk+k21UazYF9NQWvqU1MeM2Zykr61RTdc4y
tdtj7fyUdOz7jG+85pu9k0yMveOigwySKowapIflAOxqaN3zJ1uKmbQ2Z5dlQlLs
snAePV90PaTJuK7RqY/uAS+PiKfh5f89uZ/65qx1xZS/nIfR1mRGeyN8qxP/eFBs
NCGxWJ7r5Dqh1OpS9WgoGktlCL4MR1EPCA+A7Xv54PkrBCgaRGoxgPysKyx0EuaA
guZYOiTw1UidwbD9ir9xFvlkCurk9PTchylC3xEma2cjW1ultW0/mH+T0zBCtuse
bR7sTvdtM63UHwXB8VMaqSBHCqxH+4oTDSgfSKnTcbgEA17slNUlgcz7orcGnUE4
zfaCq39QoPsaTJ2+Z2u9qx79nIokl4R/Z9QPaqPXx4sl6SLM3U2cIVKgKXQ4ykn6
Dn2Acw1b6dRqgWm9NYyMuItFUkgSqnYIJ7UPKzaZGXVHAKgcXd574ubM3HlFw/sN
W2FSF5bFPNCI5OH1NkYZgQzIKsfuHX004rPKwKq6wRCmKFsnp3Ur2sdhJshzKUUU
J58De277clcyYm1oZYpiDcUowqPzaXSsPWtVHDPDAuIp5P/rGgplS/EvMP3ZPgsF
l9t5gj3QcCL0kOtI2XJ64nr+oLkXMZ9kmhVvykDEUHxPvoYHu3bTLgotQuZC7Fts
zwGo79Au1iYCyAD9CbbeNPYjMmyIGteZInVw//AKBgs77zYDlVaVA0uOvEsxj1C3
4rknLuxu/N1KfZrmg4rz3AqOtu/4DamOfNYC6+57XOn4uPb0b5nRiFMaMq5zNav/
BC1WOstlbNNMlCYNbRGNRqFU2m9bSAGujv0GO5PUIBAY5i8F2943p2TyXnBASsOV
AkxYIpvTcDBVH+O7ctUdKL62nvsXoUFo7sFb7/NBAXN4yq7AlTFnHj+lozqQ+JFw
pLvQ3rZ/AF39dMyr2HFwDzbou/whBKeYo+305scki8Cb9n0ibnvqasL02ycjEwqu
+ICxKnIEtJEIZns7Jwk7OnfbqgnNRCs9Ao+4hITHtUkfqp91OSz0nKEAL/pbCGxH
T/BH4B/eMB2PC6BkQrQ0TAg2q4T86pdcjKF/pYig+IgmCNEy4Kd5CCJ0+scUvCOS
XWF99yqyXj22QVVLdbh4MFnbU12OktEKtHQH/BQIpXZcANkH0yqGow1hf74SjBXu
qgpujtw4LoY4V1WAELkwu+tu8nryh11dI6+pxP+hV1TN1zE0UkRlryuZsYg+iULI
66AVpJOoFOq5UNr3WLohR0O2VmFMH5iPShAWB1Cc3JmK3KHsF6K7UwN81Mda+UyD
+EiDKqVvJGVqhk1o46RGwnsg40oBOEFktfKiUzdlZ0SJ8fE3r6B8TTMbNVb8ab/6
jBJ4NkCwIpaIkH8y/kilp1EQ3dx+kt472fu0j3BTBIwd5aJehVcsEgbja8geoNdS
z2iaeCZR3aGgAx21PCL//ix7X7Ai2nzLR3ogl07Z4BixRPiYB5RxQKe1lH0wY9KE
n3S7ek28prdN1aXbpqVjXo/QUmhaaMe0casj2BGBxikw1Jdmbc2S+9n0FF9HndcH
tL1xRYsLX6YW67Bv7ii52szfCS6TZuUv28Bb31uBa65OP0Fu3qmg3UNumD4gvkVO
LdAhVyWBbq+2ScsfFDJM/A0f13eJ7gkTaXRuuw5C8PPWFzL37uCIO4KLu4q0+RLE
zt/ufb692JCXBh+i9ZO6FSLyteav0IGlbMHbwHjfexN9jKXa1NukntFxMMvI/IlW
9mSUClDuFjdhB8EAZ0tBby9s5lBcw8QiQcHGb+Od71E+24Ls2KFPPYF5QuMNZljL
Z3dfA1ufOTB9KwFfkaSD/JWcwJCBKqu85TY/Cxitj2zh11noGyousW0RHNHOo8aK
D9hO7zwX7FCzYLgd6vjRBYt0/uoCbLrSq2wQZAz/4np7HX1J8y/8dRV97rKt2TR4
phZQcKTEN8YzKNO/IP6cWCAORL83DIdRx8bSeIU7sqracc7PFMq5AzZmJi0rWk4e
+hv2UxVgMzVjONj3jMByvEZoTgCZKN4tfUWTpe58o/lEnV4oN/DTVAfCJUdczUvm
tNO5LK4mJoOXGN794329Rc368RqN8GCUjIsntgIVzXiwJM5ZGLWvF9Xz13soTtwH
sghpX2cI5z46rpRfjPUmzLRGiwvBbAqOVxFXVtNTZBVhC3+XSB/IH/k2hcn+ofig
DZZZNop/y0cn3RAJBngTHkeiq3zrwcHvNHfOJFbOFb5Nvh8dR6M5UPrLu9aXwRsv
7F9PniwWohMwTYSbJrwOhqFlrE3Ek7KPZ9r9Z8ay4DZ+bV71sFLK7BwKY8nHS7S0
Ez/O41S6RxbV78bUMfSm1r5hVs0GGIeKjdC4ZMpzME2wxqyPJjI72DrtVu5tOu2n
lrjIRqnK8dE0hGRMzzkW254V3Q0Q+5Y3a2Ex9gzWMO/IdO/nIIpCBhVyXWJvXNpp
ZcGs1yy7XXj+BnZXZnBrDbyUT5PJRovKlqA5co63b6y88JlvZ0cmofPTv4Inuwfw
O8qmwoSzs5pbj23V51j56VPJb5OKOs9S8PQGUHFZfslhG9T+cEhKelBDIkUz0U2j
P+WoP/zELb1qMHKMEnckpdPCwS4c5dbladL2KvekPObmbb2s+7idqLc5xsvoJWwN
tn3pBirKFexfhw88xeC7Re1uTuUUyzNdiz9++jSux/AUzZ7KKGcHFrufEmMsgJY2
pDyInfFlDfS4LBFjhkySKwGGzT4t1EBvkVWKKfPsdpUllhBPkaD9NmTwCE4WYJKA
doSmLFk+GAEFkslP5/LHzlCSASL71mudAMfw/dZhry2mmvKG+XCOxPlN5hofQnVN
C+E36wXVU7NUEJqBgo8Noym4qpTxPEFw7k24/ztp4AxKGYaypb6E0iILXaS6vFir
IT6Pn7eteWYjKK4zxQdBLBlXbZ209hazI6/s76zEkjacmuxAML2EiPxKSCMnYp0L
+t9q3awIuQ2Swa+bR/xvPKSIwCd/YoOYukaUfG13XIeQ6EWxR6vy092HGj1GrhMQ
PI3ywUG2c0cv3kJW0GPvJuzVEY+D7x3j9RBrYK+jbqa69eXItmy6ZcY3N3KAPmW9
Voex2kHzao4y5w6uUFvyxKp+4TYKPIgq8PL42LD0vGCE4oJBfRXc6PK0Mu4JEiiP
GF/utROxo71IsNObDm0hLspBumc+rzWeguTxPfBOAXOOsaxXsYMu2Tv4Y0JOJOx0
GPlC0AoMvZVXKaTVoXLvU2davDN41nrA1OJgxPF+ZYNEO9Wj1YyWSbtNOS3btpQp
+ZmBZg06cJCTmnmw6VV7YdmzyQKsR6Y9vyM/pkG6Q5jqhiegNjR1ML0r1cqgzJiL
5SUIltbdo7l/wRn0BM1AX/nW54zQXLpQ3HTL5dWu1jurOea1s8uEX2rDbl0i6eHB
T4QRr1AkJ/as+KdHsOCrC24KOYBDYrwYb/Tu75A22dMWXI/nhNiNn5rY3V0spUGS
QaJ5uzsewULup9tiLALmel9bKA5iI4ZnGYJlwSFIbtJMFg8j8gMBMRqQYgtsxy5h
lG7AzNdCZANmEgVC6goPHF2cornpByK89u0zwag4eRcKi032DxW8IkG/TZsnpcS2
Wa+WoMOV8tAOEyA2TmJJQAuJptrmms1gzyES5NR34tCcyWRR9T6y6wD0JSBhloPC
JzTsC4TsbSA/2zUSJgUYY6RhOvsx1Y/j8FIfZFyfvfMM3lMgZ4/7q+79A+wWEpp4
4ZxCoD8oQAgWjBOQXxA6bcmDvy3+1hwS67/oxmvgxShrBAltWM2qknlhD4uvwD0v
Ybc72Z+BHQH5KNdWtm6TThz2mX7gy8CjkXb3xNi8JsWPgGVD3ugDiRHH+XFGtwVk
ZQaxBrr/JKzgVDvEhlHXbGX3MjNu7NrDZ42FB/sTd4xDDJd8WRzf/NPf/KwUFMaS
+z8jcWXTssMoaH+wZIGWZA5Aiswzb8fRf00bQaZwm2bGbp2mTM9bFwfW1yE0MI3t
hHybpHxvilMZyEfQK/v/x0cXAk5IEY/AVAAkSOBMwAWIoUpuykppcdwGdd7MipKP
bY8y/QAahAsisEanL/Vsk7RY93F/RWltuq+BCvdSZLm/Mqn3bJM2d2Yf9opkG6xx
bDbabLiyJa7Kh/cjd+Ob7kbtm/RVDy88juO4a18xXgyiEcHYBPSSKtPpjiGO1MVb
lrDPNgTBCGZbGjs6gUbXgJpQ/4VhlS24g4N7tustiwJ86gjAoaExr8ZLDbxP8eoe
4W2udR425GeiXfzF0oLnQg==
`protect END_PROTECTED
