`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
159B2nk8CvDV0PwN5sOG+DsLztvbKAkz+M1jm7dOXdZS6FtnwuBva62Fum+PRxGc
+X2b+gelKoBnozoqpOE6UOyJVCR4fbn3WxfFblvIHZjrCPkM0guB13NFS+uqdkdn
j+OHMztByKjIRRWiDCAfB1buKtey0751O79shIZDI3Sd1oN0OWzSFiiJWyqsi2X5
qG6taeFVFwku72DjNaFybVn57sA41vINoa7gqIVTqm0JUTBPCkwv6S1dmodaoGCr
MhleQtyZH/FmQjDZF21lprM5eZkXtZttBwToeT8kYft/sxU2oVXIjZ4IXO3i0xmE
mkXZ2qRLFrTkZTPIhTl8ptsQxTUJBZCpv3I/pBhvbOtimDuhfsTlhlVz8inW7uSv
xzXbP/57BOF6e6vDnfbWjmLE2cBRIkSB2bm2wUvj4CubFCghOsOthv3kjvjmPHNe
fIwu7m/8WVeh0P92JVL7DHEvvjDNJRkwAYccDBmPtcem6Ky53AWvGOUeWd8ghSxR
Cr+KyNhDFtCopLrG3IQTXO3b473DyB4pFY1ElY8on3RYXZkSs+YuFSvcIdZ2fCzX
tkP4RK1hmwpCwP76mFCAjD0hR86g+qeboiEaCzfChJMWgs4fjF9mWdqZlM1pJbde
BXJk8mHIHjCtOUd5krtTYlphNIQT2nBn2qiXpXqgRYkhWiHcjutmju0fV7lrf12k
z1O6+lMl8z1jn2hDWkjOkcm49j63Z+Mx/H/qBvsCvUWWCRJSim0ED+VPCtYrCyud
Jt1mC8yATEP2ZvIl5REG7x34Y5w+oY43/5Q5u9+/44coql3PUEzv2S7wkvo1ZYA4
ergKaVDw7hPC9gB2PbXvfczCA1p1+HztnD/gufN8R/2qc4R6bdB191hstuCPlBCf
3AyHnf0YZHqFxja3Lf35er2YcSJ+yvQ9GI6lueVNR4SCIgZtXHPvOFmC/FOtGKW7
KYCWKdoVIhl5MrP3tmlAC3KV01xe73qFWiN5jRFaueBQThszQKdGTt2yEYsdQ5V1
OXyBwvTUE6LbzzIlUypObX61Ctog6lHVjcfO7o45y7o5qCo0bpp0HSRcjhwsq3zl
w2u1oXWqGkrLjQiPnhtjvCcUF2SCqeQM85fruMnBl0DoyM0rzM0r9Nle9G386Our
4cm4aoXmWfWom0ntom4Vaejudfw7QD5jaIJ9ijC2+0sxkvwqnbCD8MqvRSZQFav1
cCu59MVeIvhv+MGtkdpdsdh56KhjYv6/YRwJKALS4guyz/2j95IhCIDxRKlWQMWt
fuBK1f3zqMnRxqegOAxjuYnUsX8JaS49UmwbV7srt/x+Kahw9qaNINw2MB+ExFln
cT8O25z22fEohgRIcpdNSA8lmZz2gachVHznlDkZ15rczZAAhU0DCrZcG3YZOC0q
RAnq/8gmBvqXBcawVKIhovwgVhNiiwPPOO2uPDflxbRUb6+mk8OCnjZ9B9UHSqv7
+xbu+q2D/1H2UDlwgYAw21QJVUMg5417Zqkl7dMwD9OMh7gfcfAZN+U8RhoWdCeB
YEAymuaGny4qEsCD0ezcu85aUxwRNjnqbHI0P3jPejalQnW7di1/xd/cmZt3hPKU
BZbX6NWSHaILKnZMCcy89ikJwP/JvvJlfrbQZ+11aERauFLWfX8aFfdDD9sPIGPP
aItVh/4mSTwnA0NmAqeWkdNbgKxwymVC2KAEoHtzdgJnJElkUpmtgOFrnwxhwXUr
Z5AAfeDJkNlos8PijDnZG/GSo5eDWv5lPn2tftlPGBf+DTzNREsqmm7Nid7nolCb
ppJ7GNdF0fVYHFp8gGGkmzlScXk6T4C3eyYdUGQn1wjBb8rZ7tMD8J/yCXNEhp8x
434Wt+xgh9mqTTdk5rpl830oivNijA8B+YDkAh3ev8humXl9KacgdQfZSXQd7VRP
ND6PeAPgrY/vZIpa/T+Ubuys0vQr8BOy0PM3PEWrLUhxV88Az8u158i5IbnZlv5O
imZIjTmc9qvDhEuN2RzdT2mUTkKBbjNee1TeI2lkToqfYjQxiSzwJ9JtrIDq1GB1
9q1ajN6D0U55voUxHYpeniXusYz8kB/iIJjoNgsG69W3CNqQT2tYOTeg9mrfWZXa
xSv2nVppWwyJPYV7vo77mMBf2rjx4HlDTabOLndPgBM2ldpjCr+oAbisGr6SYMu+
iCvzdiqGkYwlEZ6fb2vtBbLCH+dJCeYMCsdAh2KNdC9M0hcZzh9iHtrI5GykJATq
oUxJ7hmoedUJ9EuI6epaoQfrLI889f66S6WXAplHosoilUUBzwm4Hdk2ROc7NaEn
JqBpEKIBpgY2rJKUl1aKn6wBzc4iQcsZu1nnFRfINVJ0SfFdoG8u5nyRicUPsXfl
kImis8v0d+YemvPv5a2f77S+YPllnmEdfHDrqC1KdcsVykEtbZ+y8uzsVv4hlaMS
XylxbP7vEOVeFlotwbukbrk2AqyL1pwDtUdEfyPAl4P4c5VPRy1ME/QbmTzm/HmM
pY6XIdcl6sp95LoKLlv0hwgqitvJFMQe9pxIYftOaz6JbJyBpsDP+AfPCaHuNXSa
N/Ni+2/ZofoaoRAV7rCasbZymqMBvEIbmV8A+4eEROsELSNa2/Ms/8eePEe5AE1c
YItVn4nkubysdN93yCH00Ni4CtElZnWiGYYZ4u0cpXowKTjic7eU7hYyI669F/gA
bjQV+dd1ukLEALjzPHY4fNuAn7X20iyf4VViXDEDUCBP0wxPSfpO4U7CPItBk4BH
mY1soRKoAgRGKX4OhwlIs1mznQBwHzTV9Y8Y5hp9Kh+PEyL9zkMkVqAVof2MPq7E
kU7zZh5OoAK0gR5KoInOjSwBcBQ+evkVom9P/6FV/ulJ6Ts9cSgHO9DOwHCF63Be
65FAUYRfLt87d6Sb1l8TP6QGvlavziQwxU7fSQx0RfEPw0ANcO6KPmC55Gm70asH
wDHOnU+Z8uaLg3s5J2+3QmKdTSge3+aZ+xpzpdQmKjL8HxjIfEM8GGzBNwZQl6w0
NRD6P8Gqpm+/hCyuW7BP6di28iOR/lsh0CAp5yVDw8Y7a+awBS/F/VxVbQSzP4K/
XU/UKhBIjGlPPymo32PH0KeaVP/12iLh12ecAy0BeY4SqQ57R2OtGrQl6FW6kEKA
26O673AVnkVibqo6rfEMulNboNGeRORXP5ilZs11UXdovYGPQRN+ui4h+opu/dlt
hE2xZ452GdWpp4v9JuAScj65aJyUYlDzc2y75n/Q5h/nu+gOmLySS76KoLtxxcCV
Jeg2/EyCO1a0Z91dPNd+gINZ7Z9ITD+PJlI9/BpbBwlwxsJOABYh4iZIn/ImTYsV
079yKDa9sxOWTGWzpQCzWWDAXVr95XnPQan1elDfEL3dspIHjKFJBmIIyXbq5bHE
XzPn+VGv2lmBEOGXAxK1CRyoLMKUAdED2bCqFLYg0kK8qhdJZE4GhPWKxRIj6JHg
ktuzH0nhVTyNEKhP7lYVXNMrsiZku7tJ2ioErJebujGiGFtIErZKqSP0WYH8841w
CGAMm0jrdnU1z/8ZH5NwgxGKOQM7ULuPAORAtLuGdUZVv2fAl4+aOOOJcvh/+qpQ
3ugyViE1rGTjBF3/wgz1s4dtk4KpHg/qwWE4Zld4hVs+e9aCEZz4lKh3gclLz03v
C7sG0kxmFfrIE3vDrN4P7pAZae3hxW/Ifub3RlxQtQSgwEcAFxci3Iw53eoJRaEy
KjVvNgpVI8GBlyM/ImEPxwQVd/MA+/PyggbyCqyI7UcO/Xc18j7iyeexjHHwDtNX
WKEylCHCKfc0lEAmy08HSQ==
`protect END_PROTECTED
