`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzZrdtojuofgseEQwtCtQ/NodXrMqwreXMpOsUf9ZMwyzqamAyXhTmsuBWXYYQ19
1CeYcoj/11rS7y+1hNw6Ty2xw2n8PRwGDV126JRJq8+hkdD0E2If79yxXwJBywa7
BTHNiVxbHYyyH4R+n1tUJFX/k9+IVYcCvrbfxnsouafMJKrZzGqUZ6fJGNAP+Xc5
tze3y+6mAhqy1M33kfihZKa26ykb6xQeJ4EbtdBfV50il/PHiWA3l8ev2J8W29hT
9ZM7lJl0gi/+5jFYNVPZE9TW5McBwPqOnSoLikZsMqUVwrI6Cy4aeBjU3OSJLq44
GFDqQeSSwhc7vCPu7TVpArek9h7dMjjL/wZVXmt8XlnJ+jUdF7JbYj4Im63hpfUX
x+bOfdPJpsaaGpc2D3mawGP6vLRczjtE6dEkX5UPaGynqDleplrdJYYk1SHAHLen
efVKYNqey5CD34NDUmWUx9qdr8JXaEQIOzHxL3v48mxuttOwY+eRSuXtJjfYq7BA
twZuvwwy8rahnk53jcRs/X97x6+YgLtRUmLcik4+PJvubkx4vCOf/ZJF1MbJAUo+
HKTPVFjxStrVeB4jjbrm3WD0PQeqi31USC8C3akYMHIQwAm3xXyIhnCPu6SVzeR6
tOE88eORmaPa0aG51GRk5vnjZ1jpfPANpbK5RJPAwSYlpboNO+Kg3KgBy9/mcmD6
JMAqz5FEFy7qqxrJgfTcMBqqWcJFg2nv7YbQ0VQqAoKowOIlbbGzYekdYUvlJYXB
BNsvkD8fd4n3pHU9hisp2a5mBMy9YAz4tVyesgnZPofrZommjVifyfXvcgo0Gt/J
SNg0TAlGEBaPYm0dGRU3PJtT9oDx/8v8Hx5nfhS0zxCCAB+bBMQ/GIwSQGbuVbOm
oNfeHq3nll7zOsG8RA/Fs5s56t851LJC/OfhE2dJuFXTnMxYoDOheAGKag2sVHXo
`protect END_PROTECTED
