`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vcV6ljvwoCl4lPHiwutviy8Xcqo477dmfbQ6sgsCm80Uy/9XRVuYyOMbD2OWiCOK
DKml8MGNNiarpUY1TjU6ceS/yhSvXHfjYXYcwG8Y20ZjMjsXMTBIL8cbf7tvV/iA
NJz6IhSPQUUzznHpnXUbv+v7GeJe44OepsV6ieHlk6w/BzYZ0RupCrCZg5ygsT52
wdahnKwojTzRwfUW6TO2TGaV4SkbBQDHXVHx4TX0wGTb2i8eYfphBTsu3YHl2v9v
hNNK3DQvgil5YI/LXvNQG7mmSOQd62N8yfWvWyQ73uFllhC6fudnkZpJGa8JzQcA
`protect END_PROTECTED
