`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ux3+O5klYqqFOb47orto1bX/epaL1yT7z5zRLWuO/f9BWHN6vw8pkN0RVfgcV92R
ZiyqqwFjUEZ5TebML8ND3NNyvUG4DzkHmGhiwuyjJ7b0ggfdDW6OMxMxVbodhMhD
HF2Up3oU0NCcqyPLL2yvTLg5iH7DGPptDkylwugZN8/LtmzzV30AnjGs8mkNA3Dz
IpkOa9j1inOt16Ghfn+Y/CWvVQolDf8JnmA18EGGe/pm2uTd1+/zZcJYeg1ORHGf
U/67U5L9YMk5tdTQ+OvzcA/Yr0Vgv2es4LRK1rK0Ol4lf4rct3O6uKyl+cgeDeZ6
6NE6Tks/KL7DUVq+3Qc2yQ==
`protect END_PROTECTED
