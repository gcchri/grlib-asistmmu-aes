`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZh2WR2xbwVmeIiqSi9OPRbzQi1p2lCCk6dms2aERi3vVqoK98m+9XBlSB7oqHlB
QO3NVk6RccMXu6Qg7PnWi/lVTj8V/3YHBFfcKd5NcH2Cf5tROeODXSjzVr5rqXpb
yfzWRtmGtbWXd47NgwVCFjk/XvdzAt8pq1oj9BOGYTnww+B5FPnqeucjidv2qXB0
U6U+4WMeJdTIdJ0gTio5hjNgQXHkGxf+oCUQZw3m+1S4j85hG62Rk7VOAi10algS
aByYgROLrBV9pHywlX/W9wfm/rXEah0/6o1mnw4uT0jt9XHcO7oQLDV8nWoll1u7
mhYPC+vzhgQWxeQO+E1HykyF94j3xBP5TOO1HKyQ1PRZhdThlCN9OhX2OgCX5KVC
diEaOwoSYm4F3TpR9JINhcc/OK7gNv3fM9Y0wRGUB2UX5tZPUWKlJb+9TEPADL3p
ZHmoD5ZdFDfwlr0/UYMmA5K9tavOintBcanqwYzH7UaBbSgaFDgEBRGMuQVZYurD
wnJiKClPji5y8dRvUyEc7zKYcZC5iA7BRjwg2cB9hOD4ugYI3o/+PDibFWjfMV9n
mvgjuc2+ZkAbILkFuixDoQ==
`protect END_PROTECTED
