`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tTd/uUlcEOSFy6MxVakmACM3o8zU9P1n40+4u9T9utbn5GeQv314YxbGnD+CTke2
uZJ8tj2jITwtVdaHcWBQfXOE+st9nawh8uQ05y0oWGNxGuz0QZRFlePfBgFZCODT
CuG2qJxBP+KYO+GfOsyvz6Bru+HlhDfbAy9VozivgVQy0JcriVM+M5kELalGwl8s
/8oI1VRY44b0nGgR84UCujIQj5BklMM+ksidEIG0l5u43LU4PbtLOn1uJhiBkYSB
cORrCSrSBGUHxYYCZP0Vyob8GoqiJZKuWXMXYbdWwAg=
`protect END_PROTECTED
