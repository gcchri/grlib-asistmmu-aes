`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4jnuBvgKNnKkF1r0Z3cu6yIy/i5DhFW8SBi3/iakxFoYZDepS54gKr0NFzC5SrY
Gtxno/Hy8OqgnoFXgXXQuxSSvez/hppABnWPHQzsIS/0IWsajyXFxXmhjoIA1TBn
q8a61pmuBbB/UsOpvj8kVt4e5m4N9KyvMVv3GJ4Q0ptnKtKq3ShFyTeIN7bIqDnS
sOH0HnU5T3W3/ucBYTVFI06/WoPK6bHeYwDR9cmtmFsYSz988fN5hp8Bhp/ZM7rD
3slZHkJEbd66Pd2uwX1fg2zJiuG5rBqOMft0psJQSnOHe0argusuhu00gjGfh/Nt
8SWhpEQZE+6MxA2YdMPvz+rRkhPzD5tO3GO0GJkBSwVN8lmYBdqmijrCzVUZnxf4
SCsjFiS82uF6CMHcJgCziR/u8D5VylnNGseEN1p5l87Ori+uWY5cuvtkQgH+XzyS
eZpf/ho0ad3xF5uSvuIn6w==
`protect END_PROTECTED
