`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q7pyxPZJbSBMMMKTMuIsbsBTwDk+pWkYwLtKUgDoFTFnsCv05++k/iSn1OnGKmr3
LKgfqlo/VB+DN6ytP3cj59swktDgN4ov8kDZ4qDhCJlIkLT4CxFmPgZgGulndvzq
iWBfTI+OxttU4ts5M/lr2FzwHwy31rRKzraVCe3Yzw1pkYj/pkn9ytYG3/9bVJ5S
YfVtOPIInGsq6f2qh8CYVm9SWuh+ELV10uQNab8KoaKs8TeY7i6Mqj7GMTQJit3R
YME5ick7QMrHt1tGVnrG5Ibj0aZCX3YUTrskVLnpvS7nETENW3eLYpbUIxYnLqw/
8gr7SRgAxdcApgUHeu4RCMCT6hiFVuicdP2/pYs+R1TwptmXcRGv4tCkDSfLcq9a
HV9gg1J8WALH0TJIesOTGUwxSMhonUUiScpqJWvfV+Xx7JyI8gMkNiqP7ICuR9FI
rwOKeYWviQfmuwT/PzIIzPGI5v1piHM2AIPi++EFmq5vWka8SCLuhy55vD8sf0Lp
654AWjT5gtCKRKFPWNDdfv8pVEdhKbWycdxwlHzN1Fx9Fn5Z5EAZvzQaYcNCBK+g
xa4+7AHqQFk6hCTZH9kSgSlC8DAimmqXb63YNWgwhIjHub+HMjBmDXgTdbyTYrSl
1C/NI3yEEcGFNxaJcpRDyVnYqiE5lWa72wWS1uZ2ozMjt5nyroJg52V9SjjAjoZH
tCd92Evfg4V3W88FJBYch+MPcpktk1DZTT5KUPbdkW0upM6iO83jdXomSHsnphxS
39CS0OxdK6kW2QxHIWv3UrAV1x/OWNW5tob2NvGxTjiYch1yPGdzeUkEVk/NEG9A
N7e1ng6RunBCfMjWO04e8U8ugk5dBwmZ6Te7VnkVqW7a7z7KbCr3quOOeQzuSEgF
+mReq05kRJXxYI88o/+KQfIySv2AvCEljUgJ5qK67auwMPodpey3B9aZz7SfgesJ
ChfdDdewLd6EE2uDtCfuBQ==
`protect END_PROTECTED
