`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCIYqiD4/H8kgTQp5x1Ic0s5mmVBMhFrxcodwSAdW4mmAyT7IyKEoJIiff+FYTsZ
/o+tmru5xnHizF5o4/3R4WScM3iC7Vosx7tgVJhrwn0zEp73sNViL2Po3TedeQtL
5Sriq3rYKgcZDOnpfa/mtyhTZb8wXcPX7Q49yz2WjdudpKQo3w6kPJWDyNvmvZg7
lSY4kky6ItjudcvPHU5hu+AlZ+Xc5wlD1SwjkZVP71pjaFbxHANxd9DWAFXtMnWx
irk64wJtFS+7da5+G39AkyMi3kHoEoaCH7TkUI1cxzKlM9vOmf3Y+aWMMs0ST4VR
IHI0tIZEZy/l4ID7Pne4eYGpSaH549oqImzIjGr3tzJ1rdaOeALcOGpd7gZWwGBQ
NQ1MNM2TIebjZqnCAkMspU2TXHWfcpXOB9Hc2gjumJw=
`protect END_PROTECTED
