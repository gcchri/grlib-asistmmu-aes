`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbLnBQnYrY1Mcy4q1EUBkjgMqexlZCLUTOqYhJnQp8AI9+J7ExgwJSWZACHIaLI0
8OmaG/kXqe0RPmdMBXQCk0IR7krmQJB3zPG6bWj//5BHfhHYszpJWpLWsZ0OMrH0
b5yWT6Qz/Wzz9Q/bGcjnfC1JVoH99BiWAQ27nQlmbWJwGCnKTb6ot0Iu2jQd4jmO
wjvXis0kk1nUFpT6giKQmpVsyz86h08nA6GOZQpn7Wq1UUJVlmKUjCwVpTbzojMM
1ugNYo9rHiiM+/5YU9KNs2yDkGIAmmGy0q8Dt1zOFOVmuIeEOb4FueZaiPqH8sPh
wOGsbd4ThgeW43FVmTCRaDBG39MKp3i2C9eHdUTKFEttuKZHZozPWwWUPPRfv1Ss
PYlaPmXDljlIyzFLF9PlD0FxY7wjzofuYvIb+M/axrZc7il+7xV/HvLceRK2QTvW
WuJhxMtCR429WOkcLqXWBVVDLIKpj8A9f4NsaKDye7KdTTDg8hd8JtCKdtkFZRbu
6+soIXtldpIKB+DS8Elephi8wUNgYHHwxVKXWF5QRz3An/EdHSHgdZPm7c2sxTWY
wqfpwWahpkIECdsaA+xIrMAZbjX6F3PgYYzJrmQJRtv2YNETEL+tVqX3JncPn1ow
wSo1bMnZTEFLoe3iciVJVg==
`protect END_PROTECTED
