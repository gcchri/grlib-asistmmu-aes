`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHhv/BGVTD3Q7w1L/RFxCv5OEbetiaybq12wEP+jIaK7dVO7hvW4DO+em1yYE/Gf
pMmn/LzOeFy/BRybRurt1qGFXZ7giQi9HRz4feC7Bca8n79oYJx+WTjvgCH3ewuq
1AMt6bVAeLC9MJKU2yD2OTE8JWwbk2nLHuFvOU9mL70pTqCk4SWvR+Q0iZeL7NRm
kJiyYpWSwoyg0lIUnXKKQKK26YWrYySnko4EhYw5re5EcelDNIrKVxvK2lhmMujM
qLVxwJd7KqORsU7aFXaPysfUh6UAEGqJE7NlbM2uymxDtjAlowCeeHio7dOScsOe
XteYQkEPJ9y6muQN2qot8OgchkBMcDWDLaixkYHpOhi1azrg8KQ9CPb2WJCoqmDh
smfnF1+6WHzTdVgdt4D91ktUby9D3um9dbeoaUyH/Rdg8BPTMtLrZR6FL5zWEEKP
`protect END_PROTECTED
