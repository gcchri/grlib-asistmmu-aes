`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Auj+W6ss2IGoBJB75nFFcTR1pcO+lWir8rRr+RosrJOGwE6bVwBVZW1jDPCfCmHC
ZMVJ6PqEw5qXFYDteFDqpEnoe6BXvg1BheW1T7fEtTT4gTza4TZiD9cw5BNmu1dh
SxblyE0+LiQgYC0jw4NYAufG/JE2YkgOc17ph36TQ/X64KlqM+J/OOdnhu4iWAol
mmA+UpWupLClmrfou1frmPI2B5aiQ62Fqs2ysc+YwkhlYm2Md/zl/wONu4d3A73G
t4dvAcI0mV5T/xMppqlUhQ==
`protect END_PROTECTED
