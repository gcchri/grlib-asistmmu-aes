`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDWRbw7uq9gFffP9k3lI3XwD+ip0vMUf+iIMs5flX8vms1ez1yPW8EseJIYV7lWc
RXgigStSSIT++q87hCXSNwd+5l5xWKkIn7RD+bzg+WkM0pOw+PXMIHz8qkN6hy6M
MA+0ObKpDpvW4KQltYQiPPu0Gw7ITk2GbI/BH42S6L1OR3UmrFiF5fCjEysSsevC
gkJqRuX7O0H6wMyuC4Gzfpw1xI/ZMW16JV46CVoZZpNUofTTT6yo0cJiXD89wX5l
U+bAHFDxB0FVHZTzME8soYfxvF6Zrm1TfmH1sGmGsM6GWI7w9hFkSd5wehCgjyB8
gqzTO8ybn4I1u1GwFiER2nmvNLk8ikG6VJNT/d3i9p4=
`protect END_PROTECTED
