`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QqmtXBE3HnA0EGaHforJgs0oFOFZXxeDgFTE9j5SD7LF70FBVDmW74FT+YW167N6
zO+7si5wxSeNhdw3Z8aKT8WDM1U84dfrla0uOyPESXpoPgkZWdfS+wqD5rbOZmjx
EPtxfft4eU/CGri0XMlVftLB3JLqBz9vPLMJoMRlOVN21ojN/itm76SxxPcmRdNL
BNcvZpsD7wdsLGoFjMvLX8q5ThID8eaoKE6brvvLorpluI8Hs5n83jrBMWgX7+ye
S5FUpqAMTHzRNgzmaf2ALzZx5Qu/hVwyHwuCYBX+IC4c3HZHw8YmfdiP4GEbSnKC
QJZnfM/JTs6kxOrF91afJxRcfPmyKsmrc/siE91hrjrVXPv74ybrW8pnu2MGd5Yx
5tNRjfFxwDe7KGi2lBuRPGmbfqN3FAQJvyJWwkKHFD3PJ/ersATOoMnHjnB8Z3hg
MtRET/HZdRrrIbmTPujcjK2kKgsR3BuRULtubvJdYkk8edYizbCET/i9mnUepw7L
06o96ZKLbn4CJqnKTR27i2+GVgrUCnqhC043k4T9jN9enTrv1i8GYMxKedFxJWfT
Km6TL5LGCfl0bIJv6KCWj/grmwAeoRNAvZC6RtW/Xu2v9pAgStCMF2Wc0xjdfToI
BsuX69/Bb6bJR3Hhb8JzVCpEiMS42Zac472XL9LKdPUpHNQJLlOTykYsueqTDd0w
dksZwjnnzS/Lgd0NIN2C2/468bExDRuVuj4CYQoAc6rsRkcmvCwHTAJGZqvbRIyW
0lxwcL5CGQ5RvUex9Bfaw0Iv7E1dh4ANArVZ76PycrAWtvxIdy9vxqqQ9Xh0dZss
D689AtTOPnWG4sryGKuDCigviafLit7sgpa3tcpTvWPANVmjhdWCvzCiSoM3xvb5
tIZ6/8hakAjJwnzpB8+POQCn8Q7iNBKh+j7q+5jsPaukbNqI5hHeybx1iZBSbgrL
4NTBB0TX62euNVW3H09FtKpP1AyQRbOeejkeXLhz61eTUxfiVD4evRd/pxgwNBFM
nTw63fIc1alYOP9DBoV4Xj/p+tytC0rf3WMoXDSHX6s=
`protect END_PROTECTED
