`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUdSj7+F21eUzDPoI64yf84NYx6zzloIvVS27SuDw8dxYmsfpHSL7YeUmJ0/LaSd
W4b2UEeDweozQ530M+5NuC0BxqHIroHUODdTs112i/GLY/pyroUWbTltHNdMGN09
PpQziFraFz1CosmrsnzpIgG712O/x41gnwIgmFIUyR7zo3w31ZOaJnqSazFPhFnD
JksffvcWarnO3ir1bOJqC0c4bGv3NhGh+vt7zUMNni9delGaz1UHj2h34qfk8SKy
SGE9JJR5I21tZ6kwEHI3QywDHxmroonFZKt42Wd0bPznvSnLxukrp9s+KlwI3XGF
B/C0HuWgT0YTHcdZR/6r4A==
`protect END_PROTECTED
