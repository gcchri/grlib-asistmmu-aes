`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qt8znmZwFklWOq+N1sOfJRo2rG7QatLEc1IUW9KbtiSta7JgTBXiNxl9hw+J28aC
xn/LgPstzv0OnZvNYfax0vP/FtxfcMOOOvfZmpKgWrqe5kzwccCoGbaOm77XuPvV
y+ougc9QVy9pN9SMnpuaMo/JtResht9WupKf0aE+77/+2AFzGhKp4eKy3gByT6PO
7E+QwB9+fYGBUpLEjM9wJRCWGqHMU1utT7/HMOi903qmV296g4S2po9dXpKTN7A0
vrPWz2sWO4NicS2G8491Q6UsSHRKWroxOLlIUuS7YnJI8DxSNCRPGdC89HGXwkjZ
NLshYMpCjn4PUEZkMfxuuyZC1v3cxiYzVMAI5bf3uJvYzYJb4kEPJ39RlGfMma/2
xJB0YpOtAnbggQNM5SgGpjvA+2UyeOhGkMHyBMm6l2Jp/SxWZPPH07pY2cUC0w4X
q1Z6huesxy7RsdNj0/TVQP5Y58JNYLP1jMVXsW7J4wZLFO0gQOOZE67UKpeEjIJJ
j36hgRuVaxr5k5jSvwwkq4nZBIgJK7QncwNsOUp+SQ6fjUkvRH24++GCwi1HnOjv
hibmrjs8mfI8vIvAAtokxUtGgaIJejEILgD4FwfhydyCPdqm18y+ndYRBoSLppIO
1vzLkXB6/3dEKxt/eSXSQ4OLV1jxKtYTv0oU8xVyZxSNfEYKNOXazWPBt8xHNp3d
kN2Gdvtxf69lR1fHI3Ew9eLJHxZrPJuhCB396jb6FXFJsf+y17XWlx3TFuZvjwUP
zbwSrl9aCWUEJyrii3mnILCSfuFa4XD7R2zXMMI2dAt/sDjPhqIfji6kGlGM0w7B
l2HSzct0kaF6nPelAijBgCOTV2ll8BP7yGluEQcV65y3cdbwp4sLrnR7jP6ixBGB
iiL/54Zs72LciWat2YJcfSukyYOMiugqOHFzqF6MVUiIes4Qp55kvhiUHTmdjslX
4mJyVnigCD/csNhRmrWPTJvZ+lt/J1MiKBYt84frWaPdvvWC6DXdA1Jbw6r2SKpC
IJf3+Is0fC5jMx530NcMmbPAhqiVSKYK7As6ChYZTJCap58jgHjk45UDwBWIX+TA
zHD6KACEZI60hMXAiFhOAm4xFgvmHcZ3MYz54S7btYkHkRRoSzyzsX/JB6ASziEa
0xKtaQW4Q9lBZYJiyvos4w8WvGkgWztpMkp2Yqwa8SOVE7s/t8F3htQ+gWztwNdu
UTRcqNvp91Q5w1S8W9RHjVE7xm9lCRZ1GSRV2Dx54lP+GUWZfokh4ggXVWzdrryK
HKoCsjW15WWOawF/ofGJcPocVNA9/FoEMNfNQHzxA5DdOBxO+PtyeVVCBOwt9QSm
bExNoNgnszo0LVdBzaqUjfs/3enNn2TKYKdJT9u8oVec0SVOi7b+QgIKN2aRZgfV
77C5FxxMHdJHVJ5mPeyWvAmEdiPcSxRQaKZkDjnuBxtIwVrUKS69Rc9+Yd9dP4vI
krBULug/v0CgPD3fDKpRZ0xmA2VuIozQRH1g8pCce8ajt69lvzptIvdkk0z2e212
WX0zjRkXhshUyVq2b9ojUMAe3x/0mzQxSkpmLQJXFggoYVzpeDma8Ook/+3D4C0c
ZUofC5OPh7Czdno4fWE343rIC9wRTQsitPCNmwOU2V7ENx/ZUE2Ju//UPc1y/3/o
KuxacKmjJNpo+vTUzkfymkxnq2LO1nX0ppm5EadQLyUYu6w5xkP6trlQHEyEIdwk
W6kyxRzB/EWEZsgvt1mSlkPuPTOfnUE4FSYx4CVu9MXH1EA4etseDuTA547su6aT
mJCKAriFNpB24a0om5np7h81dfHK3x7GZtADcggalWQaXlwzVl9eZu5qLhA8ZzDW
ArWvV8lJrbF+Yk5FL4swbWP16vYDSdXVGsMcO7b5QV7Pq0GV2wBJ7rFhTcPujl8T
6AcTKmFyHaiWjpP1mZTty1bzmxgjMcf57FQGnp12KU321OF3jniPsm4IJxQVryns
0l1coILRPYHPXjDe6ZTR/dPWLT9LIiEOcvkB7fQ8Q9L+fSuUy4kDaZ1sPcusygb2
WPRdyEkvLMBz8CXkMfHHry0l0JfjszS+I+kHMJttJEDtUL/+Nu54BuhndikF6awC
`protect END_PROTECTED
