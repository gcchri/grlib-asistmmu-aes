`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvJpMQssabkN8GrhRYP6xfyaeY/DSsU2H1Yx9g5wb9ApCRhmQF1BacmV7yG9cUUD
N7G1Z73KSpmgDY5cnPUaW+hhgjfk2zTApUphC4lIjUo7pNclDqH/q8yjplCm2KdZ
ui0wagb+HTcddLxRpxkOh821xcxjFNGoRO+QL8QkfrEPXwxa/2fJ2UfH4DEURU0O
dk5SuaV6xvrJrNY/pH6QpMmGOswnaqecj624mh9lf8BmukoKUVHsrhXHf5iIeIH9
a6R4bNRnU7OEuYtrit7sc+P4AmiP35ZuXmC8KQ7NI3/gwM7PHGALkfh3mlQ17JjD
ts//+SCLmi0rh6JIRqZb9Z42+BNZk1LgQypISaPZKea1ctpy1zFXd2AtW5FN+yvq
Zpnu223c5e/dFl5cUNsODCGQ6jCa3MCz5dZyWEzDnPRcjNhSRpI+wqT2TkDmCWrW
9vOW+GuUSigmab0jie6wPPNy6CTWvHkzG2B4TQqmR56iR45t5mg294raL8RP18lc
SciytrY88b8xKbB66PlVYczi/jG7Cw6w406uAiixvtiqIC3sQ1qwLlyNtrPASnd5
5Y7cgJkVKz9g6jr1vjVCViF48bfDEBO6hkqbdjSI5CRXvVb2pKiQYzN+rTigybGg
oN4TXoWyssIGR9gKODgGx060N+YL/Yz89ONbgZ/DKcGogBoIDUwY2sd+4BoQEteQ
PojVh3U6VhivnDe8Zh6egYNo2KQMAwSurROlL+J278ZEke1es/JgNuM74yS9qYqI
fmTu5ZKhFKTj9miojYmpTPZ5gCHbYUpMR8A/e4uBNHReuOuagxCajchDJ+P6edXW
d46vQMzVnebLE0EXXlC3Y0Qus4Wwd0QhCcOTKtbeSacf1/w+jHQdfGx2P57A0Dgs
GNvQROKfnBmTny1r5tjkrT/0Mcul57Rk01Q2Mlp3jcgc+yusqk+mX/4mpOUgfbgB
9kHHa5Rr5f6j/QJBRfosAPRle7qXhSIDxCtp3mj6kpk=
`protect END_PROTECTED
