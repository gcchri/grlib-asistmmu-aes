`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Niq9LiFc4mHHQcbHnIU4tl8uLMbAMikA3ldBknaaz5AgDu0Ax5OShH6Q4yGOIqB
/7rmZt5omVQaBdSy5LvVxJ+xn2ZkJP5CnWewnd2qDxzBlwMyYL6w2tAQR64v5JPO
ocME9HWbvNPczix/Tf1Z0RSbS6e8JvcDee388xpuhrjwn65fYdtQmvWgH1H2Ed4l
VbfR/t/ORH1+JDkup+tRhEFFdXFPDn5QFPnsxTn3nsD/HibtaSGnrCMbT61OryNU
TKvDwrpoq0+9DqnVH8fROQ==
`protect END_PROTECTED
