`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQTqoWZgzzzwoeTq42WTQrJB2uQU4RusrtVR5kE24EN6L1Mjsf7G8pIPwVmO7HiM
Pvh0Si28P9bY7/PH2m1UfCFxab/HF6gW0lU5I1kQRrmdMktPlyQRjPet+fkYi+CV
tCGfKe86+zj7jnEFgT1tJkyoXLlpPR2yY/FPGyRbXRWhQVCMuSXNxx3E7LWuhW6d
cznxetzRrN22FExvUEwNTT0Y0s6wSGrjgqP9/gldqnbRlLTTOj4KGJQk3wh38Vds
FTu0leHlOFOcyQv5o6fmG6KFVGFyDlDawUigA8uf+j9cyUMv4L3vjajogU0VHuFQ
i2mjrd28RGQMFnlDGN63GFpwkCibZQZb9A8EDuodxEIoCdXEcFyrr5LjeGqJfYXS
KcxOvX9iqLdQUviV4Ao/y7t8yzMpwoMkOeCe9TbZOGIMmg0HcWPTdFcs0XYC3MQU
olOKSydb+njPE+hnJskxxdFPlgsAi2HAOMvZQztKmdaKsvt2QWw1HWg3jpIM8C/S
0y8zmjgohoNFnaVcHDE2F8J2+SZyMno6UGj/es7YX0EkmidbxI1aR7HhF4lb6/J9
9yDZVkIj6zi15fB8pTdaDBkPylwfa+210jH6X7wTNCp7DdOUwewgBcWtdxwaMHEm
ZuqUCUOblMMhCCFtQwkICwFtyD1Zr1TDgdyQlsKHwuva1ZI4XDvuz7W5Y7AuYDys
Z0s02ger9V4W+XSsnX1LdlKM0b3Wsfzx/IMszp8Ty1t3xoedL/qsYfdOC9hsGQDk
3ipLKwAGSx80UsqaQFjs2bEVDlwEiEBGrvxiTRYgDUyUBnUUh/5XU84eYXKb9pav
ny4Yv2zvkM+ws9w/6Gx9rw+Jqgd/Bj2Qp1Dg3For8//xAUsJfGm8f4xibZVbjN4l
N+RIJqUv0RHHSj+hXzpOQt4BteOb+vHTqCUS/3qlD/m8/4xmFXNvdu1DMAQ5mYXl
j7+3DK0d5AZeBJqYqJ/kBcCXiczw1FQh7SP+MXlQskKVxRE+LfQM52UOCxmCP4VQ
`protect END_PROTECTED
