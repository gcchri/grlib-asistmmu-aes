`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+BEGuVC9yY8SCz8RxUjK09N2Z0BTxDfbnUFU8leHSHsHLX6mUcqj18s5Z+AUEDAb
1l75LLdllSMaGu/NvWhIrL6AMi5pIl2HNpMOEyOIigC1NHR+iOVU6LZABQPtsE11
rnbNRLfYqIxP8I2Vx4+ye4IifSv06qVFVOgVS0gANCZwEGpEEHsv4ZtfzmOxLq3W
EUVv12hmK1P6zeWeaaYmXmdN3RkDAUnRMomHfeuoFHc1tqvEFx6+nZfpJMEHQNY5
pTcFagFcKShP9M62Nzj8vZP9yM4B6KS66t9uhTgTNoyQfc1VaXNt5gRTQieEbe9G
H7XleAyfYAKBuJr6BbGn4/4VJ2T0InhtQ3kCW9sh3wxsvh/rE3DZSYm2LUF3HIhZ
uhnUwMoHEDn/2WyEKr0Fk7zDIw/OHagp9Yl5I4FnZHy9mjwH1CmIBMUNTWisd70Y
VATYPaQ2oGgfUNp+srOp1y6gsaLJCYbY5kUBDVh9U/w2QIikg19jnZNlJJTDVd0o
t+OFfk+QjY1lTvJ3Bn9AV77VadFUo4gXLiiapDdc62Nw7kMqiNIkkXag8fTlpvNc
P/EKs5waHI9+FbzGuojb1tAzpcPWz76NAhsTFUONir7hmlm02C+Z/RPVej+6RZ5M
bngQLZeMCFBcpUlqOeSBEQ==
`protect END_PROTECTED
