`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMIis6fRWbdf1GxhjTw5ZbzCHMXilxtLkrKKhsOyuPDg2tYi9XKAeM8HPHXzAZvG
GTBeJ3XhLsvEd9U9XillvrtIP13bHY+je8TVQFFfVfSuY86ePCRbAO4eV9zCy87y
zz6TbhlC3LiP2DoIvz7k5yXONmL9zREzQLEGkjTXUKMvNOP1VzTh4t5QIIdjCghQ
HbIssWpupRQOOjEljHiKE0A93fWo/0W6ZC+ZIkraG57vQ1e9t2jPWF61+Iaf3d9D
8Doi0h85hscCvRDUrRz2YKGdzjyGu2qSLVjB0ibwwe0p4U+Pwws8eNOKa83PK4fq
sTPfisUiAkUxCAAsWGyYpnxgisMx1LjGECE/FXhah3SDdLcwSIo359VKgkg5/hfX
aU9sM69qixX6TG0MRm5z29m4Ef2naYT2eRSS+EbVBlz40Df4Hk7rRyyLRcP9ljlc
Xk73H2BgD1a9Sh+Orosr+QBOZLWrWtIYj1TQNAlEsC0=
`protect END_PROTECTED
