`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETMrhcyQkCw7FkkUUZU0S5sgTwqPiLctXW/Jre9zaHoNm0Ovw7JQiK5h7w36q4CB
qouqVIGPebRzE4eULBoOrx5Jq3p7q0SBwVeYEOGGhORFGsUvQVCUNG/aTl96KBi4
CVFuKyCrG8euHJrtzRhNy+T7odoLkqkZZXFfAHeoTX0+M0W4jsDw45MR/6KfEb5I
oqfg+bJ9qT8mCmFcwjtbVnj70xJ4IN0aF8KBdY6Y9ldjf+p5MTfJmawov0e9Ih4l
UMFt3J7OJd4ZAzaaoNDp6YwKP844HkFA5CN7iqmboty4bFdSrgJ1tcga95Obr45S
k5aNXhwXoxwiSTkHHZ1VCsWuYVIS5cWT5Dw0l1HK7H/L5NViAJs5F9PLMLxC3gBQ
rzQ+xuu3/ApQKHPLfKXDDrnQ90A5/T0/rdPO6sA1DlIGntB3x6pbt/+Jqp3DpIy9
yhbVCmO19GH9RJw7bG8ZH1PC+nG51QW2JKAi/2yvVF1T/Q+GKYa3VWTSF0PSmAgR
wzus5VMsvnu16M9RBLqSgUrk6JyrNDHpWG9c/VoOgtZa5yRMOxPQrQpVhB36DitK
DjoA7GxAUOXIHBV3AGjxxmcL7cV1S7rM4tKMXMCuW0WRST9wk+1zmAJ10On4Jclu
RdlGXd9btvjAHpTfbmoac93lZsr+ytVnvjZHxr12b+Od128LXS+ktGJ9k1WbjUwG
QidCMuLjjnjljFA7fx+nZHkwVeF0BLROMKzkPf5Y9JUeWskeoqT9h+owsruw+t4E
lHa9g2q2Nto2HSGiSpG/QL64GgbWT9XMyCUyuIOSoeRYfQ/LUvRhjaqFVPdbEcQU
fkcgiNrcbnJRwc8+p4eUnzPg/5unIExI0RQh2VQddj7EihSOYRR+b34dZdLyKLfu
mrdhN4Q6OK0qH/3HrZeBKMnRjTdlyHXqMieCH9atkKblwxZkGuyC4uhXRn6EshoS
0VHPLe3hiveofS7cRqM8ZN2zJN51CNYeYVm6RGAOD2F6LUw76k1vUJyJX8Zi4uUy
+73LS0UmHX4NzL0QAd8+c2gyUG0Psb7C+m/V3vmBADKdGEsLSt1na08+29KQA5oB
KlAbX0MCW/C8T5nGBOzLuYHjYoCdZUlognwgBzsDFAoIc4YztzPmncFBzVXF+HHI
L5HHs7sXBVWdyQLFpffnoFLYRXP+7aet0srvYh+OFPzEAnqS/sCm7GJZgoYSEWpo
Sd3vzvTuzYN+0olgAjQEANX/8nbH5tLbAZPyeDlbpCxJ+DJmhRiCxo9K4lvJtRQx
HE0TjawJxrnCLxhitWEYR/yQH6ancmctXu3diAeM7JOFAgP5B8iLWbmePzELjNfP
/n/aHcNoUBmbQynE9bUWfRq6moTQkMi6CfCp36qqzMLcuveVCyCV2N7Iok7DPiN0
8W4CnGo6F3fP9YSQE78kmlq97Go48adlPH2MJAmoxYb8eXH8QADYIAaU4FeL/RR6
ZoBrIfqTWyv62e40SIEHViBdoA8hSj+Oiqk4MeSAqyyvOZT5lF/1UFsxbuebs16s
7mCHa+bz9EyDfCavY2bnAVQQLWBND7a1xMxxO1XiEruTBQ0JefJydQu3nejMLjpa
hqY8I7oqspeqilzWBsCSLjtdl7iigjgMSGHpsQpm5cxqCbM0EOOxXUnn7e3tcyjt
XT/3yJmBQKNCeG3+tEC0XYmCA+agqUxBBrEe1mKEDvngceR7xp4N7V3vaGdi+i91
n7AK9/rmydS85nArlyB3vJQvGKpxvECoIcUYw80tJfN+8B508BVwbHfuUPeDAWhD
acKwTOowWzwCJPAqlZOVVhNIN2CxWUk21rL5ffxgt/RjOQGeG5pJvaCMIy+LMoIp
gDEeTQ9/okDYeaOWFKCJxBuCjw7hNz5rlaIW1OkIo7n3ETHEglK5vWNiLK3UJOdV
lfqHWmdewezHIIJOXBarrwhvOFyksyt5UgvplD1ETi1cbl4fkUkN55SS5Oq2C12/
IqyecjuznHuovgPjW9YYP/CX28xGxUsIbD2HJWZhRWTS6XtqzlpD5yWi027cqDUQ
2va5UPzEfU4mx8XSrw6Sb+RNmPhCadaB38nvgCfGO5Db/Er9vP6fzm4WRBgHlIZi
mFlUENxQXwC9yhrivvJIRpIvF6y+th28uHe5bjCksb33OQZob89EYzyoSw8poUzL
A06eNRI1ujGIAfPbpCGq3iI+/H+eE1uiX54qsOxsXSq6PXclpxOapP2xbiBYM5t5
OIhvWAzioVRG3QGN90nxqyPUzOVbZDBctbct2aDaf1LWy35ZLEiZck7Lr/e0mWTC
oXd7K5w4OshUypBUlmWEBTI3BFNXDVvBkBhDfKVaUDPvR0TE4n7+p1kJfxFLFENZ
NmnnEMevrSdwfZWLzciDjM238zLzokyXT31QgOpy8aF9YKIGF05NIlLI1+6aCHq8
eE54jCCpMFFLvdjaLe92DbLEYh8Vdng6uRyTVa6iXACqvU3l+iurbxypQPcbxp+v
4Cl6PzP4Q4GFTDhWpJDvSXHjpYtlTrVMZeqpLchdsv9swljo86EXkHsGtNzeY9J+
bUKMz2JoAPdi2Cb4NmlBcj50Ad5xu0zSZxzhV4EGuO+F2DNuA5IbpuJdRWWMEDJk
DNCdDSuiijKB91E01QS5mdHMohmB1X17IT9ALdydypQU69yTITPtAV67Fe/Fx73m
Mty42OBuD9W/J9Fg5P7nu2z9TtjN8Pdsu75N4QysiL7vSy7OrcaVhI7ZLEX7pdnl
XtOL5ebUb190V4zaomURSuiwZwpzU9opz5u9vLKUcrlz7hdw1PpF0W7MEPCa2U80
E/TOMBVGD9DLh5cF1sJyo2W2IFaHQLWU7Fa3agVeUwyXL/iKkEXYcRTf6sBnkLVF
d9U6idXfKEQyZxU8yE+tOBzT6UIi/ZSiVBdC2ostUEyiXlcOERABBApGsnTOe7aC
96FObTdHXc7VKWmZnHNQYiZRWcE1XOTPteciYqINH6rlupVw6cgfMcD6d1oPOFZR
NdvY8+RzzVqANT+0/Z4Nh0WNbPdvg2N+U3rfL1iZ4a6Ya4ScOiyvpg+s4kWgjDDl
4o1loAYuO+IEPAgOEbeGP/DahB/9R0ZoW/kUbjh2E6ey8zwfpM2HWQSuojt1nJ47
XRK+jIEFDJ1xEM7XyfLBewFDRLvB86M/fDg9rt25g7ODtYySZds8PgEX64tI159h
MH2ww7XEG0WOMo+v9I+PFbajUdBDjuaQyaHaGuyyNdJqZvO8fsMvQiboCaEWqvuc
SzjeDnSvQ5Wg+L5RLPV4cA5eFees9lwOypz7aaQi347dy/ZyLnvLUvAMywtjSQmw
OIJ42xru7CL4YYOGrjQ6ZeKqKhzQlykibvuAOhVZH2R4rbrAXeKPiZUohQ8mPTL+
G9jpEGcOv/jFosLLoMVaDLfATYoUGvi5YfvliJg+VdBiRKqdTeh75ZkaAS3Frdih
MKGfURGOV8UlZnXj+wzKP/iRhr/42rqWOe5MNgTHRolu+5EsRsh/MLdnTEXImeU1
G2i2v/ycWe7q3kzHaSbvVTmgDaeiViKepu+0zx5eP1hkTcOLTze/jm3jSR9OWpIE
8V2//6aKTL0i/Ky70aadbp0G6V3b2nVaox+rPPHH6Bx1QVNSsD+bR6glFXF7vJrr
3acLJyGneN7lRjbz2GNV9sVWJUFO5/2f/lMUgELhJDo=
`protect END_PROTECTED
