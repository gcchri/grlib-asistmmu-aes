`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
71GK+OlIRpVKS2s17sF8SPkyGVbLksJEigPMFCfK1gnLBsck83AsVnJ3VGDJuONG
PmEeEuk8uP/aCvLGeLtG7Mk/Jelsz5esYi/GQlGG+YiUyfGm4UqkPLEhTJbx/5Hr
Ra5nShbcv0Jse0jHQcxyuFZJCLrcYAtqFhaGs/g8pvzs2Z03Wgqu9oXhqgGvqUfZ
i5IfNn+ZXi0RXg5OVhNu34/4swhrNgmcGLkxft6Kpu1p668hotIhG7CwtTLYu3ce
3Mt6aPkRfMkXVc33j4Rdlgg3nUW/FUOQ5y/fBZdPBZImPFgGPaWa+2OhfYOqMnGV
VOWmXGFpSSq25GFgGtI5BG4IOAtV8efCLE8wj1ZkSFVYrgktqpgLBP2AH0kaAtky
OlNE14kgvDBtorNhze3U/8Qrf1m+M1fSn+AU5Ebcu6YLajFFxoHVY43hUsfShp0Z
WWpO7Ax+ex2V/AAoLbVvepXDPGMiWYVzIG6NrnlgoH66fo7wtVxwfqF2re7tF2F0
6lZ4GOfZWUv2k8EVypegmqHFwQiWhyd4ykD1x0mw3+QcK7USDkpgcdcScsPfikLC
6ECkUem0Y8dmWM3NQAmz/ORIbsGFiZBk6/QA+ECQB7gEqJ1odvuy/Casx0BeHYzM
96ch0kfKerdqcy36XRYGecnYP7uhxIEIHx+HjG77qE9TNlTYNKp50IG3afsJ1beF
5Fco+XRnEsgB0swsnTbELlokST2la1bgCMIarIwjE0rL8pvZQlY2k4aGgcdnqzo8
fTm14eo0coLq9f1KDKkC3q8yTj7FYDduIg9V6vr/d1srQfuV9HKrAfEIjblNP7in
rPfewyJTzae94XvGQQ2mtyGznL4o7w0vsS9ku/Rv4RPaOXf37LtnUkk6zZ9DGUxP
OIjoMjXQ3Zp7+WWpxcf8iEKS6ezjSCHyqHKEzYFX/h7S0/ugc/1DNwG7sTo+lznT
d3scKz73z6VzpY6rloTLO2IauFPd/I9wz35VpoTFskZEwXi4waxhYpwSt4EsB8Gp
5rjbAzo3zn5BWjuqTqFxwSdQso/NBcUoC1Fh25wsPVLH1XUptq8BGsZYj/GbBORd
0P/2GfUa8Rt7zlCOFKzbr6ve6LGkS10UTb6to4L9jQry1XRtcJ9RUgBVhgxcAsD7
oeWSiiN72TAE2g1qNvX+O0GWBGGEdoVAUbJY51I1Sx4+59RowOz4kUhb67/Cdquu
cjM1JCA5X7SBNp5iic4538eoWXaoTlnBII6zGZqCBBdp14XGHbXKTHhY4CelL4eQ
0YXSmw17705v5U02Cvfe+g==
`protect END_PROTECTED
