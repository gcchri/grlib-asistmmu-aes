`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OXpyx3Ipmv1OVyGG15hbwf3CKjqY2XYN/579An0A9nVFJbWiUObxluMfnaMjJlUf
snmnASg3VZwubwtD1VszT2p229Q5SdqzqWWGqY7vKVkHIPbEHXNsIYkifJwdX4WP
yB7G1hhPUTCg9aq1qjWmlfIQOmODcPeWNqn/n5ciMbR7U9t19woe3DP3w0TJRMMS
qex4z12O6g0oYm1u/Ix/ANAUkE8aqWnlxbMMJBK1gULiiySx8Zxwfi2uOWEEKMmN
qjbF5wft48hjnKJKNAOSxx5zGsDT9ALm+W4Y51MdTWw=
`protect END_PROTECTED
