`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHd/mGMYYtIPf9muMCJmwWbJx2aDyiDy5pPsxEaDvsveYNVBC8fZc+1Iy0FhrFc2
0f3lYWljhw8DktnHmQe8Ds2uqA+ebQ8lsujaeGmk0XxREEnjpjL+4i80P7oEivkv
1i+Git1Gi61w7ZSkMTBRKCw2ZMafSs5JLsjaPN4iSbnygcw0E9TLC9g/ySqZsHek
LQHd82isuZNMO7GSiI8sJQZBOEq6cY/EC+nQ6LVpVnwF4mKLE1uRXz9+Ql3gDul+
h3WXDVwFyZk0t+zLps6si7lwiMprW1yD5dWoa5yZCgyeHuBLmnAVuj1dCMhLB8dc
CelFkTOJ66nxtM6jZ/+YF/Sm31TK+pudm3G2NLY13YGM0V0VJfDHeJP3ZBnU1SfX
nlVUaxCoscLumiLfuk8E/A==
`protect END_PROTECTED
