`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X8rX/RGj7++JNkieHIF853ht8XnP0MnGa4F5YOxCV/xbj5z2va3uxJ4FOiIZT3Rs
srMXeBV+56suFihDG2oETnn3E4oq4iHwiJdq17Cl8Vr49MoxBw1SlR/0fEG1rHtP
mE3p/CDa5PhSF8EztZUGppFTjH/5PXbNWeHDwCM339egynB24bwMJyDyWb3J7PZ4
VAxybCZ5QlkDqoZNkBrf8e/bDLMfQ6W5D2UiDf8XzyOcb+QteUoayJyIKO7EOTze
yXqD2XcoM1m09t5xm/nESXoPPZRxUNfXme3GnQxXN552v9T4MkFyFGDrpx6QwQUz
sWtQ/d1kmvXWCiGWL/ALNVhDRnNhBxxAQTJ6oKpa0MpzJ9/J97ViYLcMgDOCmngf
/GwYYhle5SJFSywSD3vshYzf7WiOa1GfWnDYMvZJwv3fj56x5uqpIWNs98B4H1T4
WhInEudGc8QMmEuD+jZjkLqXsCPb66VRLNXJG1+rNvJL1lzhBEkGxQGSf/hwYGmb
PdsCRholhZu+wOiCmfcCVlqRGQxAr3bV2pooHSvWASR22t+E00AbdN07tCc+y1ro
P3xAkrg+YAIPw4d+FoaMbT2V1DossncKh8oOwt58+nXck5lucMsqIcg0UQBeb9fo
aQ7GUa04PXUHi/h5KCOF0kuqX8vuJ/wefvo1ouEtllpciwjSIIrxu5fpbTYG+4H8
goDUSIns75deWa55gzqsqSY3kxRU/pHGa1kwXnBYe9ygtWS/NBlIP+Pf/a0uYrXM
eATk6VDyP5v8Q6jZ3GPa17B2GMUsMYRGzyMWvTwq4RsiNaV9GG1YLq9Te4m98Dlw
vSMymX42spq61Cw5l3fvOzfwyR1gIuU6Rh1EvB6nRP4EYT4gCxmfYNinkovdtZ9h
XrGX79n54EQqAumErYbkphscGaBeTVkE7XPZJSytMTC4HvwWowO4mG5h/1pqw2JM
rTiSxFvrl2NnpAVbLPp+r2MZ9eaT88CUHpc7tn1XWsHujEpH3IJhWhqnMB91mHZW
iLpRk/IY1TFeO11aVvpop8pSBWaXK2cNnOr0KLxXIekkrlZR1wT5rqxteDp8CpM2
NF6XZO0AHuef3WZ/3O91BQNFfxamEGmnE9xCAiaRfQwNbjbAqYr86rTMEBt0U5BW
Hiz5vR8yxjjtHVs/nlGbks9k3dbyhZhxzqaTEe6nx1w4omubqm33JmVadMekTkcP
Ke2g45EQUtHfzS5ljHv4gqhLPejaMFWM4Kq5IGfrW30YA0LVglkXvcUChkx8FNDi
OxUOMebNxyn1wgNmYGmiJ24PNtQgSqE1267k07Bv03M5WUoOhfzK5M6xsSJyefmu
0P66A490cE4CIBBC7zzFDfRCLQgTsZe+6YA4lq9eDZ2MGGHo3cfmK23XJLQ55VHb
WaUvIipiV39QgGzJrj6iJiQHEsi5tX21QeP02YPYL56UprjnQE82hfRRHXm98Zdl
ljOHQqUdpL5pmsS1i9OPY2bQhaCqCl9dY+NbJXJtnTM1+rhJ3HxU+6u3ty5nQw0X
RmYo0eQHv5cL7p+eVy0tlnIJ21s/2+D9U60BZoRjSPUO0ZlZVvSIXzi1/WAqa4gI
/hi74r+QOMejxBEpREbTMa8zUYHRMw+xX64jWpalAc5i3hIwOZ9tENBm2+a/mCOe
5KyS2Exds8YFoQ+BKPI7qfSVIyDCir+wJ4nQZEED4gl0Png5QC2Oh/q4GdYKMUBQ
vGTU6ftR0f0ZDJzi1xTfv+YaXRbe1C+SAU6/0xLmiSavvL1nuhWLFWzNMAB8T5SJ
nhkW0cozgKhF6/ENsYgaIk6ZHEpkhuW+wd6J8wlpUhE7UNATB2gW2B9ZWw1upD/g
sWDlwXD1S6vbP77bAesXsjq2R0hYmrys0jIArY1XRUob/A6j2CpbOvaKHTtErn6K
2zvAoGjPf1AeCC/CRq4FheT1bcWqs6J4H209XQBQZu9TnGrLHUlRskDEEK9VaGQg
aIxp75w2a4vS1/5kWhP8Ji1TDUjZ3ovkw2e7VekkPL0mKJxlWyYNq1h7fF+vnaVZ
4si2jyakJlUfwFhhcBFCL2RXjDnM18y4wQnfGgD2ne4zXC52UBc+B39XCFmvNPbr
Qfglobc+zPot6JQ7EP/f6Eva9MS5sUn7k3KEHSvqa7RED8YCfu081sPh2VXNASM/
tG4hlu0BojOQetHq0dbFVuXsl1PNsj2KSF2m1zqzCIUMciKrmnZZQD8CK6EM78lU
WljWqo2LbjZTTEIzsOzkumvth/8a9xRSzwEBs1jTnEJpXdFIRjzscAU5rUfEE5Fb
0uzcUUV96fKAyS0Od17KHtt6st3OUdJX07lwvjtY5xyrQV+zpvvCxEnD0KCBkYwp
sBjFDWHtM0hKPSdOXAUlPIZ9eYF0WJJ7i67Vqi7Nl2rOJ+VJ9KtbYfcEcB0iuQv8
tP5SqmIQFDv1V+nJiAaYrjA58bOiDiaWmu2tKUMeGU54cYQxBFW5GFV8oGR+LtAu
aLzAYPRewVLsUUWAWelcbbpALTUEIiFoPLeFNo58TMWm00wA+aErBujFNYMT5qf6
s+YJDIhB3hVqmz4q4DjSHAX3f6Z5a19ZhRp/ghdLD1T45Lo9e/nG2nP6rWMHX4lH
TPPrgSlCZF8JUwOB4KuaPWdLMWJyhtLpHTI3Ev6aKpolwi/+U+7B1/ubAKKoKeCu
rbYNFBvjmNKpjTY/CvQrTQ+WTX5ytjuFERRFM6dGslLsIlQmw4DXvbxontOS3hNn
t+o3wPu4j0RqwOKlW9A2wtlAeSceDfdveSTSCaXA4Sl8Kht+5rjItvrTPOW9Ncje
pQgxBZcy9h+xTts+3RKlyQTVBJ9cldCHV+kpFVNeoFoYIiMqO72pxWu8Ms2uazzL
Uo4W9iDmaigmp4EHljCA3rtHIzJNuY40zH8XicXrU2G5yUj2K/7K95GxOXxq3q1p
Q4zZ8Ew0hH/7DZWPZOtNWJSIjumzDsVw0ASmqvCVxKbzLPDAVvlxPFgB4Rjbyp5x
ySjgA+hQ12dvciFgnvJzTq3ZSQrR3mDpsGu14LU4dHvi3j4M6obXtLQ81rYzpKzV
QeNHU6KK/TIXBIU635FhBU83dPzQ3KSgSKz6N5R+FZMkhRdQ+5AXmjG0RGt8aIJO
bO6iBGxAmR/DXIW0z1wz1ecKUR3cObvuHK8GlR5O0OPh5Spx9ZHLgLgRYZE9HdZN
bgLb/YJnCMZ3I/o80USgyrLbpTSKzBfsL3kNssaIerqkDS1FYJq0xHLoGScLKrmo
FMPGoBDCNIcMMVi3w0Byz3KPwKsf4h1mrtPrmiE/zU57aMr5Rrjn6f3EQdM0IGWI
+afsELvY1T5zNJdqzpFI6Aht8Yb1HnsbyjnpnXrheUprjr1F6oAjdUOzwMzxeIcn
Guo/vYx3C7wKl8tfEkJ0sYseCFsrSn8Cx1OixGrSla2ReOYIBERCXwtld8WC0f1S
347MfZBzKO4AGy1NPCJKqFJBMG9PTzWc7KWSVkZlc5ZR/fgBCxRoRV/F2pCXLZI+
PQ+hnA1PpFdLeBDDJKBDOiUkGE3kN2CXab5y64xeWlG+B9lkJjWM7mDzPUc7K/b2
wCWoA44XX1YUnvViEe6l6juOChbg61rA4Nd1eMsGVv8w4lpUSfbFbnwYyXMMbJ+2
XqsKVQlEQZUEIw1F+A9T7RVEF+7uqjTganJQcYfDCOGl7uJze5SR/t+wLVzi5MTD
TRM/n88D9NMi2hi8HOHvZkyeQNwt6xbAVVldozYIhmM7E8gk9g73xWHg4a3Q6xSj
PJQ8uqA0EZ4AdS86Ay0OVjuoodPNj2v5fM8/NuHi6VRS9kRynvDFqFngoBYUZ7gZ
gbvrgTbfiEDLxK3Qq8TCE7A9/x9Rfizhg97UdahFZw2vKp7G749MGVyt3tYMiAUR
rmahmbO38oJ+Lwi5qXQn+YiL3LWtdtR0a53cB/1eiyqDDfPU+sNtS7FUfn14DPw0
WnymbPUVBoCrL16vWrwIFL96MrrZ5uzPr9j1aZiYFf5SPOaeLutgmLuXifEbzxqC
4aWnFqDu77CTkM7i4ZvDZjMvNBZv3D+FsWLBlEJlIgFz06xLEzz4LLh/1xSdZ6NG
FZCplCyh6J8pljtkCuKRUhT1Um6B5TluZOB82wM7MScOjpgqzLRBJ1rBYRqDurLT
1+0q53vi4mNTzuk3EuKg5sI8rov9f8kK0bgxUplMJ2dYYOQ6jDCee42F+ih2QC8w
SX/SnPL1TRX9OutVU5umS0k1GK9+qTsf38sF2VkGp6kvceI+lz2fvsnlyYUch21L
pZsEnwUV8A8FEzLUHDtGDsz23I+P6u86VufJTZU7wajRVGvY5E3O02mQK4jcPyxI
4ltPOZYBY1oWYx3xIo2WpWAa+OPSoRTUo+7SbmoS3cV6sHtm4zZDEtudbFFxiKkK
MZE5PgMGKdiPv+2JUDc2Xv/JtzRrvaN8asstKPM0HjW+OpeKAG3pD4VEew6qYWRo
HoHQxlaH99mOivJvywNytKdUcZsEZV4LpKeEWT1azgtLCKYL1RnxXA5BOq9wvyd1
UL150XAckBE2XQ9p5T5Z8xb+yNvBPLv5/nF4MOovUQJfrSWVgRSSTed+z6QaeoTe
Ys+MjXnRIvw4yRvaSwtpB2/ordXu5YikW5zt4fghbWPLZ2qSQudCvsQKlX1qI/4e
1S5ly167ZmrR8WrTZ6b/cGPTd7dLC1RCd7xHI8RQKTFMc7w9vZNOiCQasURAd12/
cTIv3neDg8T45VCJGry3YAA1NZ+BwfNbI0WF8wpTXeXjiMWztjn/6qHObJ4Vrsyx
noQfh/xv1a9wCYB22yFCV2/KA+G39MSIzldsx+CHvyZT3p40YI8YS0WkdXys1Gw8
balCd1PdHbl2nMTT8pP7Ecf9Uvke4CcvqTt6N9EYaPBi44G565HALtbGYG7WrkzS
Gwv1gBkKTCn+jOrp5EBTwToti9z2Fz9qmpgJ5P3puhtxETvxNo4/n6Az3zKp4ULs
fGT1bD2xrEUVT7L2XpluqxspFM6c3Q8O1QC12ebNsc4dwbefxrS5bZNRoEwaUEwy
mZQnCLmsbrox8h3h24DgyvXimQqjp2NvU0AMW0rVUJIwVX4IuhlGeI7Q54XnK0Yf
i+6dI6hJxVoWM1RSVrm38OP+pXisy58P2lU3fydAte5ei8vX5wp/hDHaKOBZc+jT
fTy4g5TvAAvFezXZtphb/OIQpnIWKbze98PJfJzf06lyp+Kho6dLwU3Bh46L055N
NHboTRCHLHS92UH2QY6Tt6TlaBMHH92xWcRvnv26VkMcmACs3g6x/wWVjrhdO95C
y3aSbZXDruSshP623NuXVvbc2vxuGS0G0YFxLOa6yZyvt/C3wfCU1eFVdZ99ypjW
B7BPIKFErHWtC4Jhf5wCJ7gj3/O2XlvygPTTIuoYxpdisb/LjJxwWQrr+6AuL5eQ
Av6m2xUb8kBPIXZRGDDR+gdhq68QsdWas0ZiJY3+cpbBx1RjgwDt35v6N7ksb5PA
MfN1RXegJLrBok51uSwJbDQF7s/FipV6BBiraaHJxCi3QM2JQq1wwS3qUb3Dqaqo
hkHLQ03CXqkbFnm2oyGw5SS7hY1QiDJCsVfljhRfM6egR0J6zfuvdOZh1NK+IP10
pG9onQI50Us539x8KLd2xYWtPeZzlpdpq2nJiyr5WfrTe3PMb1obiUzvlykS2YZ0
XPH6E/NfzNPgcuCpAAVXzQY2I7LnpnLEu156l2mFOPwtF6pkoaLrGMqNDszq0zIF
+urkCvwIOHCPIx4c4+V4+tt8EgFbQOf4B8SYV9DxjZvyqQsZuAgSnXBxWljWd2XZ
emXmYqNiIxVcHGzpP3gwez7PB7XkFvAhSiQn383eTkyKMl1ASE6moNLqhJiMtxMz
IWTZ3UDqeunTLakTFuIDAz5ocYt8uAUtOvBR2ktzBNs+++BC28Lo8WjExrEzdUTf
7fKXNfQUPQrFOuo3JI33q1HAs+yba9rDy5enyqtK/oQ1z6Y2Zh7aH39azS0WMxHb
L0V+uFjKnL3GAr4ybMGzXHdYFzAkmFwP62JjhIN6wsQwukCpnP/j6Ec7p8SS+W8s
gv8ACGubpLdGpKuiz89by0WJedO7MFgiU7Taw+I1Xjgj5fTULvJn+dLueJkYgE9q
RGyxrTnbkcNZKzIbCopHC0bbCMyOq64RViaXvb/UkNURdJAAfNgarSPH4VU6hirE
znGi6hSp1oOcAU1kJCiIoMbTXIBz/0CkNFWcqr3GmIk1As/dXrl5WNis5HWWNDDb
kYCe5D/aXqZ3udpPNiJFKb94DF/FoG3mxSl0MQW/6Z7yT4/8jU9hh3Zxg1xSrqTM
lgF4hcqX9P9SmxJWnhmoIZo/IOHmbVLa+IAr9CrlL+ZkR7XZ5R7Ss/FOLRDvlhev
JbCW9VmphFcB9P/ICu6zuQD4p6Ctu6ks42l8YwjhHQU5JViw4HjaOpHstJv/qAME
f0IstG0qVAptFlyL+E1y5MqMESn5VY1HUlPckc+j6wZ7v8rNNiDNB0UTSRTFmixt
mCIk1gps5iE7X2TKJTB1SD/Y9DGOxCFUNBM+gZLnwbzFO7DGqLCIE0BYpdxifyl0
fwXk8tBXH+g5mf8eIxCFInlCCEI2J52KkyblYY91kjEljQ3fLxx6FT6oiZydHnXf
aDmAWjvYO1h1DprhHK2EgGYohVI0ZqsZ8dFIce0QjXplmtoG++jkret14abDK50b
yKBjBSdsEgKN/QcUoq4emt4ZORvL8MbnlsgBSfYvJB9ZiE84B2rPaxE7WnEnVQIw
LMmgOg2kcNYaotfseFK2tgZkeNi2U+h3q1ZT06AlQ8iLRz7GcVvfWTN64oYoYA69
AVilyzF3eTjeZsJpeoP/DcMTU0EMj+gr/9YN1fSWXD6Xx9Z8bCWDI2FmmcRy706D
6xJUtF2uJL8NxpQV/mWzhP15rbDN+eDuxR6dOU9nM05RtTaSdMliNu7/H0ZgNGJE
PHxgFvQTpHhGmAZ2pzU+3ArLJlMvUh4yRwOz9smR2NyJv06xyRe6ZjcVW/3DtN9A
g9d8i88P3mDlZGmuxhdfmXPz+quQIUByo2OgyCRYLT9zWh7WJWv2/W4q/p9HUtNQ
BqbUGpdB1SEogF7hPjQBKl05bIICFvT48h9AwbDeI4ZU4c7Iv3MOS8qN3DjKm7dH
w/jLfQLjZnM/sIAe/By/RB+Ez5gAfYWzHXLMvNEv3ESGs2lDzOfaJiSz9MXsRPit
iSR0EUySX2by0czfv9CUj/ap7Nl9I/IHagsXW4XUz5q8I2w8W6gosQPy558YxpOP
YdKXmOc8tfgBK6CqO/sp6Hg0mRPwaPhESyuzbosggo89nuOBdKYpk42bNR0sFeG8
UdCoX6iei/QLHtkSJKqBvrzhS9llwlbwrgbhzzdPmUNN2NmhrgUG/3M2x18ld+MG
ry4Dnb9Omzx/wLQIBU14lhbev4X9tCG71DvlSs1SLoPzAnHiQr4zQOnvmUuF/GAQ
iYlJAN80QZZCwHPcSHPsEeVSGgyzlr4NiFgfPPUIzSW/aAyC9iC1Rlh1xPbvkDSi
ishZNfYM/Ef2h4K+iMC7eYTxtPZrhs69/MHtK/pKbeLNBzSY92H/vz96LHQy+VHZ
lQpoEHDTYbMt2pz9n63RpDhKUf39plmUxwgLXHerMlOOgq0WJzA5Qafui2P68v92
IzbHNNxrAJmA2lXnUTjGJIkeIkzr8ZcnvQ3b0a/5b2wq7cHXpir9L3cee3qLuFoV
JA4tTjs5yNAN4s+3YLrFralH+xztURiRvw2MlzSr95deLFb1by0P37YTL20LWAzl
NE28a3WaqXy9Uq5iotVjcsABdrqFm1aWk916k0z1SvuqQzf/PBp8noRGVpykxOAs
3A66VaCDt1AXoIRdj+EmWGWdpuLCohzUl+OvSAAspDOmrlkahazJYnDvc9BvKV9A
X5HCJLB7Of89zZ+asAesuzPXu96+5p26jliz/wF/4mSLEWwj8ozCQIsJiDcq4UnT
+IPpYl59teFW9hC0CV6Vh9496VacQ6IYyoji6tFXtj14usoTtF+riwnU+esasvWo
guWtUM9ySvH2x2WzwfqCudlvfbv7VXivfbU4AyyeK/RTVgYQ9b73MUnf12zjwOWs
7WWMe0vlDxWyxLHeVfESXE9QQ5tuQQMxuTCcx8ucZWK+TrOEHcH964s/790at/7O
Y2y9fYWQ0VdqoRBS8zYWNcVrMc+oUPww90JXvkNdzkc2WCJeRKygJD6SvfXjICNc
aOQcxPwKiw2nBKMgdMjVt99XiCvHR9GFDwwLOOnzTNkC2udM+ydgupS7wewdDaPT
SNhBRzmNIRCP8uL2KmdRmVSnJRdhbYcD4g7e6luS0m3IU3LmBvo4JoXkLZp4Jlfe
mrtlo5hffhixEKgfuWRCFgVdjG9+42Mwo6Ix979fWMSu40If0LawjmoXpTSXs4kB
JjUQ0aehmM0iEmjsgT8pBzjIUpjdrlCiY+HlHkxdSyqOr1p8pZ3NGywsvRJSjtnc
oWmpM4sAESei4NY1TjCQe3ZVnPwv2dGoIt5K7LUkuR9jVGZuzIDyNPw7PgN/KaHq
nJvFVD6sSQszWErBsKluY+Elq7vIQScMH2DjqZ3uT8E6G7UGVFC0bYTrX7wdKHNH
i0DWAsgbScMpHFZx6vhrqh39pxqb0KKAKmeFeQdMnMWKKptzYmwB2c/86zIfZtrf
HMI9Kj5qlXZQ0RAbxHEIIr8phGDceV27ScYiTcbP+ASROfBSQAvkWGPB8P96fbu7
B5frvKsQyypJY2USm5KPo517nXRaCzfMewBq6oj9TNVwQLQ1HhQ70uHEDNXXB+Oo
zaqS4b0StGE2SZprHbRyBt8tdacSB3DCVcQFqNHfELi+wmQs0GrjgIi9oK2JcArn
HT0/rceQuspbJROlshcumA==
`protect END_PROTECTED
