`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhhJumhsz8mWMOVC/ELMdcgwml6gN7e7vlLcI2gwsJGwcGuA5QBR7/ycgVGzjvlu
g5t47w1xny6novtRCEE+WApsX8MZrftdB3b4ICgZNk5bxe+PWNaElb2yojkh24x0
DnVkrGL9eOI+46SjpdEQIYU+pDECCcydNcanPFBpI+uAKaQQtOVuwmzyzhAjUaoF
3xy1VaJgKvCPHqzGz18k87IKcvodYYHEaPNrcYtLiilylVCRqKk0+hlNe4f19oxO
51aJQRUayJMmu8Zt0a3jGHoLbtvW6KPUbNpqCclQI/lU2KEtlluoHMxiBDE+Th2c
tfpHqnO2Lc73vSU8QbbZnHlEeG58y7JQaNqHj31jMCRCU6zhS+AWYuXANSPInCI5
DANIZ/0uqphSwF7ma7YPHEq4uLoL29cL7qFCb/amd5zwuT+xdu6mKiJkcBHWD7JO
XRiHZqxR12i/eZQw6FfdupdBCRHxiQClhv54gaT279erk5QQG/6GwPsUN+cNihoF
4Wx6JnNAzFxpUOVKgUB5Y+dfYwdxYGRXkV4mxshDI86iMIz0pyVFBhDu3o2YHsqd
R4Q49SLti6cEetjWn8+96DHBE51xdb8A/C5bgcgsMVZlYzSegkdklb3B67HE5WhH
toVMtNieF5CekB6P2LRIeQxXtv05qbDe3ZP1breWlON5gZn0+/reM3rMcqbVXzOY
C26E3m55EEDxozdg8s3DuUQFd+SPnE6eO/tVF2oAMlVcnyPLVwGJRZoRXBC4K0YL
/7lMjlDLR8Fy1ZCqWgvbYNqfyKpdwboOiNgdAytAGTgLqCYoPefTE2V99T2pOPX8
zSh2bqcHcrWS0h0dAEOnMULxJGhSMWVfxPj+jMy/y/AhH19J1ZYopW5eQshxJ4k3
PwS0S8L4V6wfmDZSieEnnJg4Mxv5bsvAKH6QvtpVJba83WVHblYsmXkYrc4mb1Vj
ingOlCQzzWmoJKJMliS3wIeayUi7eoJq+1Ff2MyCkfa3jIhi+Myt91P+HphdFtgq
/b4+9GpWa/pgjXI3ivnj+OtyvyZdnZ1fCNnHN7P80IF3ETqv7/AwXdidYXOi5l9U
F6NweBY03GPuotnhUB6vAPOm22E2AwZRfNk/AfRRsjXvSTjmbvXGN5lbdw2yODGs
jGwUsD/frxZkYibIKz+VRaYMGx3+u6GP3oxUssFPJaxDdTKWmrc9hkr4cbAAouuF
IGH9moomYUEpTd41Swn5l4zNyEyCnD6kMq4uj5v5RGt2/GgCcDSV6M7+Xlkw9DPb
LV9kmOuaoyKOPREgLExQ/gnolbhVLK4F1ZBHcujRcbulesipea5c7UI9o7M7Kv0s
D8zJQ58rZDnoGres/HOxIe3vXBYPWe69bwHf64Idc3RKkH4BMJoctz4qXEoz3VF7
4z1Y5iMI2V5rXBka36vAnP8NoyHCexrc8Bof9N9sO7b/Ow/6mazJhrJIQhurd+Yn
761MNJBBLjZ6xQcY361qzdxG7QLn3EoNCoujjMv1OjIfFC/5kDTq5s5vUvxIh8Sg
YdgMdt9i226JEiZPzOLkYuIpfWWTztCPpgPunY4O4EiNyxzPBO2YPST7iosgkthq
jb7jbUNiKGfnOhcF8y+k2GOEQ5mAcJOR+TG9gkftMeoY9LlN2Sh1Rs7+OmfOsH0y
YggrA8my98eiv3qOgePKau0lbOChSngG+OwoRUolCB0EZcbp0dGQdXwv8TdCPmWo
cdN0pICZVDzUpD+q7rAPsr/jqmc4s1tuVLG3gu+lbo3Sw2rGhVMTiTPyvGluBmkO
NYzChtsiWdFn0xH2kVesdI4hHWQyb8meiGWWDkwawp5/5VcPCFCPp/5QcQru5a7z
1R9X1zZ7l5+QEjcxMRJPC57MIe1W5vS0yD3586uXxjN+ZHGFV8ctJvs39r72O3rs
iI/dhF2+ekBo1PUBJ6oP0BKY4UmGjbMcyBJC59VSufNZLiMrbUu9vbnKpYkGFVbP
LDyilaehintIS1pb6mbTI7rUImNPMC4Vk8LJcz1OxWPN55LRvto6YJW+sUW3SgqZ
XS5HP74ryUuvSvZojsEdkhTgWEhdufRL5oBHr/iKJ+Lb6reJdg2J3ua3JzyBGp/z
Be8sgk/aUvKD4jq9PIApXuJZW6ZcIBNiMW4jILlWeGkDCopaKjvyseKRn+jBuTSv
mnw2MyRdFNeuNTm1x1KUpv6lae/gMt5hWkJWQ7bDRhsoKxcc9Q+wNOF2oLpW7fgh
`protect END_PROTECTED
