`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LGVp+c56IAOwsZQGZJ58/Jtj9DiDTwgemeZlkVXUWO1xSSoGJ09PLG0vAFFnPxg1
Nahhao/Ep6Qhsu9dcIDyQGJet6U1QkpxVjeCO4KPvHE66CuBVzjDrKr4rgNZv1hx
M5ZHr75Ri1STVIxcHJnvuEkKHu/yi0yR3L0zWRFARgAtFwiB0u/uPCYX77l2kXLf
6LXawxO4WPfeEmcmJwtoLLWORADx7RxzCy7sAZCO7QgCkMV4SFioD2b6EZr8lTou
nmcH3br5XeucJZmL6EaOp51b7pQaySaD9cHRpB7gN4om+DxzgWYqVpz0LMxo5MCT
Nm/P4HlgV9az8Eo88+0H0w==
`protect END_PROTECTED
