`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Upgp3+J85gXyYJqDyM9WQMmSdaKjYIlmTUMmiHQjZLBjEfaDWSN2la4WajwA9g8O
UXJXDHzW1NfR15vX2oMkKBMHo0bjSXauxHfeKwuyEO9PcLs/2GO5M3Toy46INHBs
Dvj58wg0iM7enSmZIW64uUyy/wOwdgf5esnaRh1d6xFhgCDgaw33nOyCtSaG4QAz
Mtd1nAM8hawLwPX5eFcKTl66c+lUR6wNXoai7pHJSz2SBwJjwYsSoX77BoogH2QY
8O+5cbsrHkv4N9pvmZRFfL7CHSpvdCp6Y1JOFngqJ0Rw8ZPXRd3kwr2uNyltf40Z
fUVuvcTdSr9GiV6KFI3XNo6EKLPMDcjJOdRBPPqEpqX7dtfxI30jlknot2FCWOgf
`protect END_PROTECTED
