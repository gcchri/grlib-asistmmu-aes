`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/f16ZU/FsjR/c2TUHY190jZGCbs2tEHGoMisUCU8tKRpT1u0fkHJQxFUM7eyZryu
+bgIqXCsSuyADZZuewwezBkSbjVb8x3zpuCruUkGoB/ntDnLvoMPid52PuJZgA5c
k2eH6kpnwiZ+PzhS/Lc/dpKx+ERNYDU+QUiQ2CYIVCHvb81UbhU7+ufdb+tLOCJf
cqGma2LNYsdw0/40wOFoAFwk9SyvowdCUuqv9R7gLQ5JQ7mj+MZS1FlMZpWCwrFA
gS76N7ndUtK0BPKYJFzvxpqqgmeLYZYbzSVTo1OBTa7LR1h12MNNPwigT/RdtkTt
lgZzMymZP50fS7+I/TcXXvsMbin2gXajr9qNnokfNqr+hI1XoOKkhRBUGFAt4qsH
1x2PP9uZqrpsCxRx8jCAI8M8IyABPYTQcWIEqZ2RhX0=
`protect END_PROTECTED
