`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VYP+Gz1uh7zSgTWCLmvs4yDiFBF+a85rlsI58vazXlqSKuQVBguy0e2ZEclBCeSJ
yC9iHyHtF6pMJUgNNwP6bwDXMab+kaBgzq2FwwaNIBUB12y4O8GzPiXg5wTSqO9A
yPb6Ph0qlnckShMGwe6gzlDZ57KjgT0kTQSIrX47Eot4B095XAkQR0LQCeDeWWt6
22JbtgVlfLYsvQNdeguRzaLpY9LuUgBnjsVM4JByKZBWKAIbQ5vDEq6nprugYhfA
YYDQy8/8VXb5bEQyRZSL4g==
`protect END_PROTECTED
