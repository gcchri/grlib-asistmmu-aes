`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9WASmfmIgl0qItQZLVAd3kiEt46zyowhgcQ5GZm3fCylac7a4q/wDYD+dWc/aIvY
J3p90F3UquezK25iQQht1oSa0MTCFLBYd1U+WLfZKynq6fwKAaCgyYN82QzvULXP
rAhFxU0DhLYx7XOMGnby8m9O1jX+KuSjzeJ6PJ6Tly46yvM0FM8BFgCFCOQqSiQI
3PWxtX/QhSC79I6gMEK3dnBmOj8l2aW1n9vmu+0oiicGR8+7Rd6YEAg6yjNyfxN4
atF9jRC/EoqRV/XC7lK+zYbBV9Dzh7UXjhgWfV+Z6RI5SuhNnzTvf0S3ubm58DP7
mHnwH25QdExepsbyuRi+Bzl92HgAo4fZW+XjG/CRcyEfjozK5Pj9n83oQDR+6C4e
UFwhso7lLBc2yeco71WBE9NuiDfBCI7g+J/6Hp3vGZT6lU9JekIk3wqQfE8FfxQH
29cCRifG+ipMNysqD8GcCGN++YKKrt3FaM+0lvxPoyh85gHokoHUtiC7F9t/1Ekv
zvDyKnkcGjx6enzZmI60wfdRzGLN421lOZd3vIjB8nZmBJhoeZvxyrdEkwnMC5Ao
2tHzBzzzyNa2+2OqzkYSzZ7VRQpfDma7h8Q7ZpiNqi6nFX4XWL62UlXo71qxT7+M
O65pQIGMAtXMiI02sfHLrO9c9/qqkUKl6gNEkhVt6QH2zTNZLDHUxZ7qGWfc7UwB
OfYgQ39tacWDv44w7vAUZe9yGSZyUySCMl3AJLuyje01AT1tldBLRA+7IMovRKim
0WT/5/HSYaBd1WlhFZJHEU+mqq7YUGUVeAY91XJPM4uCkd0EHsjQtORuaHWVM/wu
gXNQDn81k8b4y92ks8MDZz69VaaqWwpOyqOS5AwG+tFIpTajqIln4CCSs0HSQYve
Q2WbFIxP9mePjZfRZNmbGw==
`protect END_PROTECTED
