`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzLWt1bGBPa/1FNysZ/KBbeYxaPyQwacT+zRg2ut3OqnOc1/6ZqLU0t3ov/Ltj2A
Pf2ZRKmTwc9uQVFujWDrojFoj9eJRCwjICnTNKKFSHNkcVWnIY56X2voXM5FC6YW
zev/JTbv8FICAJ+zwLdIwH0OpGBaJESyPnK87je6OJww75ntWPCVm9uaTYsLHbT0
We8ud6tQg+zLj4DLvUigN1qkq6gGTQaiPahK3+aOeCL8J9+pd/xAnt8prRx6pqRA
Ky5UVXCBctAHeYLoKr4PHqW0jq2NxDo+fIq1QH5s7Orl6eTdU7ZyF9sbxAUSrqLB
DePJ/d8ytoW3La0tnx+7pL9nqn6G5PnjnduPhg6HOoZbghmk1Wq3I41ieKyE4o/j
KINtCch32AUvfeGBJSMppU7LTKWh4ysorV0Hol2wHVtxOmFoOxkVSTvP7urBNOGj
fMUaeDPybKOjFCu3vUShcFtJuLkqRuaEKmQF9wgqEAU=
`protect END_PROTECTED
