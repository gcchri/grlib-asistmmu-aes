`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HHv353yDKSnATnna5vGrZh3Dt1jkpLxnjCgvWNgJzL02c6XvUJydwoDVOp5aUKQh
ZNFctrYhjFWz7SHNroZ9FSuF8eC4wcau58Tz7/YGA9hXu2S/LXx9zZ24mVRO5VfT
3YE7AqmnCSR0U8KC+lrvG1ygp3kakrX8m3lzWF/T8Au7Ay3p2Bleh3QKkO4yHaVj
5ZPYOtBxmxW3y5rOG5jLKFgvCwWNHv7xkv9o7/0o1RBUUl/h5fUCnfyEbBiteqBQ
SSXnaZZ8Eu7DxZ9feeQQ2rTPB60P8ODIMZ4zuwcNnlI9ePiirW5d0TeOlXqyylSc
7dGAaDiZM46S9kw7c7Owk4/z5X3mZjhmYGxdHqJg5jyJjWqye1dQxN4G6JWj0IiY
u+S+ahaOzqVpm4PJPQ4Mrn9ZgmSdMUljFpj3UKf6KUXClR+jGvlPrWCDoWUAwc6y
YR3HDPe3n1yZFGTYvtOjSXoHpNXck4p0oQVo/jp/v55LcE+cDRgjuqBML9F0WJ5y
`protect END_PROTECTED
