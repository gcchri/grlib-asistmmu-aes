`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
04CJImbsvRk73+QcvjcU5JcathJgP9kX7ZERuJmoLWU0WfgSU11wfoiCf3y65UTq
UwJtlSUc50hFsWVn2XLMibAGFHrKtAWgkJZHqjSKYe+amj45SCwb+j9E+1JRTVxJ
Z13M/92YE/aaZT3JGgydUxVCXuU5Ih0qgUTssOp2aP1G+dgQ9areK14//U7+IimQ
C45taKzyT88sjjzLdnVJp5B4lM4Y5D6rVBVamNwGNvEw2rRotQaLL/e40iGEtkKZ
xZ9HozkNTtZGuIdH7ub/d8UxQekXb1G0QyptGEeMlhn+r/TOQ8Y7oV8YLPBmPhwY
gn6BwxVT4ukMGIgBWEeyk0cyRwH8ucLH0tGt/GV8HkLmX5dx2ODHefshBwIcvJwU
4WzURkn85qb22MGKtMHz7sg3zD8Ulu2fa0Jk+DiJp3jHktOTE75kPvUOoAtyxPvI
ePIuJq01tdXkpwmqezp2OrltyvKE6mQLL0pK49rw21jZjwAWbXP4Nx1d8s4Z+Kor
th8aJYkkTnEQ1+v8QzGge/1iB/8KvCLvgcWNa4ah4GH58KsIpZMPftRZAVF5OCIX
dGi0Qete1kfOTytb4AS9i8kR/n9I/N1n99a6dpqb4i86h3OaGbqaCJDJ7/NHMsLc
SiD6PP8FfcUVdV2spGCyfucjqJyz5k3LJ4imhTOH9q6Ywzf5rmra3BERX3pERRJ8
aH0yEqNqDHVsnIGOsDHPU63T3WmxfEaI5/yZsH0+hMxRfeSJxZMiDFRVZmnvw/D1
HU4ncux1xaeefsGix8Ps2pdLd5AUSMyfcqtMvUvKO1OKRhHwWkJM7Ly40n8oDxJN
RGNpauFEojXD0Wx1fCXfN7bbdVnU+rG71+PYnpTS/DktLDxnaz1qEkDcduWo1+ka
nF7R3aZd/FQ6XYnf+Mne5Tz+aisxLH7t4wOaXhUkIjPwSNVBwLMF/x6VWWLyVU2f
`protect END_PROTECTED
