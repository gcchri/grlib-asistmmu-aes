`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljnBu/tGKgJxsGp67Gcxr8ZeHpfkYyLBqaFj2o+xwOI1JvvXBTIZckhAfo9MkKvF
fRdhzlh9+lCbVL/qa5vwwcSrLyPc2ISmw4foByw9Q6Tcp7WuM/KIsN2BaDuNemVc
v+pXhc3/NqU1eYObOKG2DUj+n1+Fmtrn5Gsg/Nx/uQh8kkLlsL2kt4oJBLHRNsYQ
o6cWpE5mgQ3ShMA46OYl9wG+UjiDADaTEuyGfMNU3etNLEN7TNXFt73CfDS9afUr
jxvJln+QEt6MWkn3vUys3F+OsK1AryQox0qFl6aR79KdDvEZlI4bx4cuEFYP1A2f
`protect END_PROTECTED
