`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FhXxlr+vrcX1pcuJwlKPC5BCFclEpPrFJ0L8dJh0Q56EdopsDIdnEd242d1yjptN
3zc7S0l9ByVduuFNxCgRduhUemZrdpyxlxmLapejlYy3HCTYHTOWPNAOXBgVAtI2
8uLwaJDcdn+fq9zL2QZgR+NiIkiqJu8GicCzPT8RYNAlt2Op0DK0OxyfuVoVgn1h
R9Cdh+foS/UVRoeuMYORLesCbnGNN7FfhvIN4+b4+D5cEwJ+IKv17rsdSomVeTGK
4uwYNC1cPzRevM56W1aCWuFANuTFZDNuAgJr/h5S4/btlLaPnGkocP484npODGpI
nocxYxCU5HkQ9StSZqWigci2ydlOcJxRRgyCiG08hRLilWbbrho9wSow/JvKx9+v
lXVzapZRBBLexAiPIJlNO0JLbOnDAozWKg+thGINTUmip6XgjofAR4Jz6E9XurKq
1mxPbA7xStFQ2JL+NQRH/QmboY8Axt8tGLXnCPPlpZKxkSxwAqPI9ZMOHcHAdnC2
dW95JRgYNCxcTFtvUpGP5CzWeRkztUSKiwVSbo3dO5U9ttFSxmWjD6n+kG+Vz0l6
H35Poc4kQpTT9u6h2fES0cz8dA9CWPWMPD/KzljVG6Xwpy/bcU+Clj8kGeVYsNRV
pcXosyq3YVV3OWX+L/forAR3S+65SvSGuIpDf6wNCBcKg8SSzv5R8JsjjNOE/Gvg
lJ4Y7cF9fWHA9bCq+aCbCeTrtTMUs81/oZPpWD65GNlCDsXn1CfWpwGV2+gLthFW
+/mU7fbe3rn2YHK+XgFdUKTXJayO+ixyf7LtPNvx/x80FX8Ou5xF+ZS72Mv1EFAd
mitLxs5LTwWo0Z3l6HOnWR/A2IYyl+oufn61gR/vo4Y7HsJCgEl8ROHWHrgnlJ7D
3S6vPbD306/RBmWwsHx01GrJ2++QqTNXXGbsYYU/Q9uoROw06umVJ1ftqk4fGMuH
MYbpD32TdCk/vvGA8wD1wrxOMGuV1j4bPM0y3AJzE97RFjun+5pu2L863JxH0f8m
7O3E6MkXipa7k9ZOS1wgjVfWJwor5+jcrETBSC0sNxDsXQsHip63NaTMwjLd8jgr
VaJhbT5m9fdsz0sZ0qT7tHK9M6Vqhx8zRPX8LfghlHfowe3M8hIHpD4iUVYnQNck
ROFelImDoIuYwBn89kZtfOtUfIiy1Mz4pRb+cRljj8b1UIXV8dc5mf5lDyLQzpvO
qY+tONimgyFkA1mWm07wRW1dHzjZv4T/wcjVoR8Z8zHbE7yrPEQhLwCpnXHcT5jU
9OowiU2ATcGKFElfZdWIPUG7eXN/tlX8czPv2pgTv2D5YeeNa2g+pptxhnbJTJ8v
IMF6DbTDExvFuTNWP7XodC6ZGsVGd9XwKOv6e4u92nd389P1R7VZkptYi9D+SOnZ
IqQblrV/ERry17jplduEveMsE+M9kaRZZvUxbEV2akHnz5bAmzCWrjPU9fx74Dui
tUafanXf1sNoIN9TZ7LaeFA5b087BaCe0teJ+3QfqaPjas+GR25MxZvHvmZtIoer
qpQ86y11EudaAGWnuLwp2CifbaVs/xcPrg5Ju0m1+ahEr3BLT39OdnwXsTFQSCgO
/NGoY7BVn/QPbopiHCedYs+wv4oLGEtMhmb3LVeHf1OQYRIGpMonyOa1XwgRRaLo
4AswPygcks0lMYBsGg3l3Z9aSDRGC8NOZ315DnHk04EZVPs6EolSm+Cz74w3A4vA
HbWkmabaaEPhnVK3i4DdrCs/orKVhx9KBZJPwx1wAsXkjR1Twvjvrh0qSLQW/NpL
R+SrOyHx3UyhrEQeq8GI0RvYF+cGDFOOfd7af2RlkPKuxzAsov1pHUvTvDpUbKZD
OnM14iE9vq1bngpgvCgVSHGQyK0hUgngGFQHD+uXueFAvVEbwAWxBTK1mSPyKANG
7PA+aRKcAMA3eXNCTHU05y2qhw/GUUNemVjPDddodKjhtstc2vn0hcaeQD7Xdn2v
e7JA8A0DkMtBTMuHJET8S45ah+j6TcKM22M+dZad2h8+oL4bV0vWiSBRDvjvcK+P
k28Hs8CfGDhGRsrTgLFHwndzXx151cmWQazoujFatRYGaJROvqTN7QenRj8JvNc9
+RdXeY3+ltN7DoHXV1UjLLqp4xCuZG3Ts83Lho6gO+fw4XwDXrOh9zAQp1W6X+GV
`protect END_PROTECTED
