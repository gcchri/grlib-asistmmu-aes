`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61Z6HqBNz9STaLoBbRBO8FvysJslkiYnoYVoN5ib8yZb8bQGjuJwZ2hBnJQU3q1z
5Eob1Y4yvtegkTEpCkoBWIRw426eIryy57MNLFlU5PQBYG1iWQ/R/wTocs7rRmQx
eVySpwYr5ndbkRk5XmAqQxBC6ImEdjLYA0JumaZOntQrVum9PBqUIdAle6bF1Vtq
rFSBa43hXOMlIaWrDVH0SWH4MQ8FAjW3fuQ9TH7gf1tYMFoZCMlW22/hO19nJKEn
XbpHH/KzssXL9fS0GuRRngOom8ThkPMXwiSSgpIffKZ3gpmJbzBBhefFFkVWBNbw
5DiMrFkSxxlLAf7J224DTJDq02bcITjQZocBFy+vbOuNyyFrta+yrJMWx9wloCqd
n9WHeUUS72JBEES2b2VsQ+r4NlUGK9mb50fau4kvczUhqsQcglb3jKX4VUjXqqKG
SvyaT96Ta5JWM0xFCI9Ww7lmRj6fHcrZfXzpy38Ni0HZPD3eYWalbotRdG3ArvTe
sz1HJV+GxE18t5vOICUJfJkerrk+mk6DOKZqZnYyDPzhuKA7j9FccgUckQaFHSMM
T6xvZaXIennstd8eBiPEUEcZzbmfyjwx+yKUUpK2frZGa8SE/o5nf9jiJLfIo9u7
Qwitm/A6Aevtkxm+8hIRjO9Px+2+zn1O+vRyKBB4gbJCCMBAvbX//MOwFxwD0u2p
u5WsbaAC7RFwoeNwfX1r42u3GXykXaBSWEPvY1t5qxfaLhX3ZwdjFHKTSx//RIMn
yI4w1g+VKMAuTVY3HgpQIgNg8lGyBzfImYobCO0pejekGl6ijAtIMceEW4JkiT2u
yeAYF1xEgnYRzyrJDDGGJMDqprBgo0BHOLBEorZ5cA5eOpBUvBg1MBHHaKgbN+HZ
OSWirV4f4nT3jmJ4EiOH9Vq+rHqLY/1OGtUBx3hUvP4q6Tp9yF2FYAI+Niq/xgbW
AsfAyaJFvedbmN+OV6EhIG+qYyG+TmktbqAsBQhsJYPtwQbsTTbyu5kYWe/pRwJ7
v7qOJJ509iA0zlFmekZb4mJ2uiig7ddO31X4h1vph0BGxdYBrppXejkR7c3MvMqB
4UtEvGP2uRD1rzReA6SSW0D2LMMFWmbAGjoOfcGXGckHIwTlla8MLAFJ8zWmkOXk
dgkaKnoKcXXnfQe/rZEIi/Pzsm3sbZzfQvt4Aaq0OK6+l0yIfWP3e70LVdkpV45i
Yo498cgVsN4c0T2qRdU4BZ98gw7KetossH4fLagPGKS81BXapvcxJ1rb0q9WfJwK
hAZ9Td6O+onjwqY8NAbFPv4BJgDCVj6sB8WCTzCKQMRKVqEIGFZBXnfEUw6CwPDa
2kUgOm8ZFsPsnpWx/CGglNuyeCJhN7xmBxBo2xmTiWTe/g2FraTWCm4Xm0q8CAMp
Wk6522Ghiy8hgOFXUCaDRiUV3gc4lFfh5zdc/o0Or9teAh6iI1jiTUf6Z7+odRrE
dI2jy5SkEDQ9LslqLJ4hRe4mbV7eifA7vUTE65y6JOZ2fQSjQotHwsd9iGZacLrP
SXhmrKGuc7yagrWxIrhR/NXKEVEodk/XXwE4w03d52PhIH34xf2IEQCjd+JiMWW9
ArDnf2kZfdtgC3lCfdXgq0cAoUFnuLX37peJdRVpT+uAPI+Vm3/K40YYP4hZ4ZSF
eXJ1UVu/s1Ih2cZoN5TixA6IC0ANFexq1aOLD0UcvZotXd16fR33NUSQsPerV3JI
XBZby3A344patMmueeNUQ2WwdpmN4WDZMpvSDpcmDcv98drge9UTB0/Mr5WWot6r
nQoNLNnTMovXdgFGGHlFz3YlTX5uqCiTymC7t8h+LfJ2ilQhTwyveo7HHsq4Tt7n
PQg9bn6uP3GE6LBeAtw89A==
`protect END_PROTECTED
