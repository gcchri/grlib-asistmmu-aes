`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOGEkFwOAT5U5Ln5GfQNzJ99ngbhcqjoSgvAmjkiyBoTYeHGL5oHdxo9bOREM+zk
/g6omlYFS2LuK7SLEdbwN7ZwoBB9cOWIClThi9dUgqSsZc4c77nERFcxU6IylcUd
qGGYlD+TYZQR/xwyh1XEse1uSHuytFZGjL0hpOx8eTWKMv5ZkJv3ir/HtrPBBK5P
qyRmDgOAiwdbmwHI7msqZLfUsvwDalQ9xZ2BTbDbbiRRCzZuHBzQh8cyXpqis+tr
zuO8eBRlo5ATsPCaP8kCYlHQw2Fu8NcnOGPjhFhZLf4=
`protect END_PROTECTED
