`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LbXGO+kftXhAcVenjv4d3MlCLX4o4cGCdDNgZdQ6WMA82JC4k+RnfEAp1x4gxIuL
Au7ll5HLUAaARG5eYPwRFd9tLUxrGP9OKTMVMfZrWvgKkEKSICvFQ8ccQODiqcXB
lH/lGYKRAeT0J9vK7nWiuuhh0qNCC0agC4ZUkJCjdPcZiKIEh2FkvKOkU5zq3MHn
fBGTwtROOcIXguPQZW7peNeCoKmcQsZYBNI765hxrtdraCo0IUWsDcZrejV/EcVo
/yrg/MsI5HhkLEZeErndU+gZypmsr+Z+1NziHus0eJUhrCFoFSmIyItSVhf94RLy
L0Z2j4K5GETfVLlXvlRh9dKOREX0HGWS59wVOuSHiPu5ka1CYbd0gPQgmU6l/hKH
dVAfVnLtYOXpJG5eqpyZfPNbgwZ3zd83UTfn/AQAGaUoTpDiUnFdkn42VQLhH0BA
MTugEw+OKZaPekMKOCota/xpTZMKIz3W5H9A34JKQtNO/dozCU+l1a0GNEXJV72S
`protect END_PROTECTED
