`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OL15q3/SHVclZVoqLFqdv9Vb1SAymd0wS3E5RmjoY+dybeKeyS9DCPuP4Q2IGCxM
311JrEGNq90L39eo2F8gpVz9u4oqGkZqJU66Vbmj1bS5RlrPXr/qndiy9Ysm+DWW
6ONWcO0KaWUNlBTbsvGTuawTMQLqUCx4TZch2nVohZSXjK4uvgRl9BKMm//ucycz
BQejcPKqWVa082AIKynA2ka0cLGVIHvJfI6tYScG6qXUEDrUsicB/ox3pxy8Rxnq
lzLFcE3UyIRqqVwiy1Tb7XdiodbVMgeiUlngOL72NyTJZmnZj1mMg7jVYWw4QqW8
8efbV/Ok0GtC95IKaBc2rEIQB5imecayNxbL6LFGWeLPjMQfXINQ1s+zMn8g3GDg
oacWn29j3ikBkPvLBJAxMePeeAXx+IiMahH3luLetIqekeMT2yc34cwSGKCdYMka
lLL/cJQtFzIOPbAmQTZ2YhtYxZG3Kem/moKnAbcmu3tPnwEW6FxzZltLLUh5t3Br
aKLSpXxNwmKi5JMh4Gtf+y5Acrzqbl3dMa6yPUzPDalOhNXi7xQznbf2K/JcS2fa
hhqtvU/yH9TxoeFmTKqQl6u1gk5O1CpE9Xrq5hWZZ9+AO8HeZrYUfwVEOeN1sZNo
Pn/hlE5sx2BYt5NELMKmEZc1rcNWFxZr4qVZ3qcdh7KZRT7ka7xCcZ8MZuKIcCDT
3JYkf6zaY1MyWlLlj4rF/9UlFtzgsSYFwrhLJaRlX7k0PptHkndbEF2HWY2PBk9W
2hwnpnEZ3SKCVxeXS4Tcf/8YObfE2PXGMpRO2iVNGg/DBuAYpV5Rp0eMRmIuvRyP
l7Go2baGabhToB737WKexWc0TC+nrn7g59ZQyoP/R3622HAp0s+TAYlwiBhOmSdN
j7HtyfFjiTYUZ4831SLkYXie68EfD+0LZQyDj9BReg5kWPaHu9TJXyzzWbC+e71y
sGpnYEPzMvW+rLyslHb7MuPFBO63avFFwU0BnLK6xOZyyDmiHZQuiQxzMYZb2BYq
7cuATBj2GgvuCGop3PYAXhdo+xq+BnqpjHU+WH3ZK6kEuGbHKBeZrgkVx2G2PHyH
gWpThqC2LNkkZo/g6Ld+Xwq2PUHRrt2EfuDOk8hXsiYqG+fLvbC1qyFv5nqizojR
7ttev6fQGLWcqJJuV7vkF0SyHvsswodyyA/y5s+N+vf275KMcksEk76q12he2vtZ
odVmntgc08ZSd4K/lxa/UfQleyGztbINno/G9RyR0M8C60zGlq/wILHCyDHjoHXS
5Cgv8tSQ+z6fJ7vLaN9iFXkmjJbWgf8NNoVWa4AiDYWFPNt0htWJfMPwb5RlX2Vm
/4Fa2WYYTdgu5WBdeW+O6LBKqvukldkTyB8iKetfCQx3NfSi9TeipLitw4/0geu2
pzrFSM6ePky2xQmQx/GJP4nPfMDYHIrjoX2ZgrLNlKRG9hi/Ad7cguPpR3Bjkg5L
Fn33nidXBcxqi3impdOTQweV/jo5RLxu5GB8wsIsx3SUB4C+EC9nsj9ObP2dixpl
wMd02xrDbSdq2KOFyomzSK7x9Dkhr+8HQjH+zVROO7nfEPVTLnp+sZ0MfuV9W8mi
j6yGT+hloIS8o2hzatHNvKoUvsvm8wLgMejSN+0sI3FOQBfkAYWRJlyqE8UKRXfw
t+78p/4xniI+uY3fqgevjpxJoYgGl8guczpoQRH+63uATwk4oorqxKVRo3SJXkrC
KERovMY9nDgFNzJ6+laXw0yZ0AMMEMomMu32+PbFf99mspBVGmFg9nROiuG0GeuS
9eOy4Din5ahPQo37JDnOkM+pIyat3l/vqOIacH++8IfXwZcNBijgvDpzK4acPJYL
xRFObEaK1hn2rPVDS8a4n8TkivsnGhBFjx1a2bO58IRpAwdpzqv8xE37ZAutaQvM
FZnZs3HLheq6cKqdQMMywfDUXtt8kh3l45M3pRTT8l3PBzCXxWWWntqp/gVOOHro
wi97G8R1O6uJdwxAuGfhcLG/iRILl5+USziacJ+mN62BvDp3qelQAAAGmMBYhVTD
uGfCFyUDODoLPq5Ew+50DeiGai1Vk4uEHC3+u/PzmA8T4pY7Ntp+5aeUbN+d4jN8
FZt7hhkZAajAGEVeqogVVGgganhbA/yPmEzz29LkxrqfQenQb7YGg7dqguu6R/ya
iLcXBjaO4kIWg/13H0j/W4FhKiUsai8a7F58M1dCuEA1IkWCcGwWQXxBJvDv7dVJ
DHGfGhJ91uPnd3nN3IHt9d765inHLoHKe2VWXQpKe/JnGw/tXoDnSRCm2WMOQ54t
+WMKhg5zCDmpyOFrxP2SDYpLAcuZVlHrVTwqmeR2vtk7nAgWgSYivq9cdMlaKarZ
UELAAInyPyt/Ia0wt7CBOb0xe71Lrv8c86qwS+fdtUCJyim3iu6WwDabhBxRm1nd
yc3lrArmZPvxnMJV92XydUNatU4UwUcCOGOlFsRgFMv3T71ptKdEvUGrZPluwDkR
MBUql6/asE0aiBCq0Y0yOckX2Ofc+f5I1U83MwemeA9JGu0I21K5JQPSxYszXxC3
zNjSGbqMtsLkg+MsM9/Yz/i0fVjirdIB9TocmvvwzgqmRHLe8hxIkkYuaT19aYWP
+Ml0nIV/LTfoKbfPuKiLLyX5ZvL18JSPOeUeaiki94iFLxNMPKDxfz6fCKYSQ/1k
CtTNRZ8Gj9h2N15Fd7gmZYMKdnx/mW2fKrUSm7FMePrljoRfM/Jtkbdu5DLtr26p
DtNDuVgCPQS8RoMYZ+l6/mADuA66QcNWba4a+1WaWxvb4vBqvmRGt/R2budt+xWL
eVnFDNThUy9jarlloQKwtYq1yt/c0MW+LauFAMyMIKjXYzk92yDRsx5WwhKmPV6k
f14wHiTrB4xcIzfrzz/mzYd8wPcfP8/+VUpsaRJjnDEArewPGsWrTNRA9cAhDON2
60zrM/R57eP20CiolXGmBAHH2+CyTmIhc3OzEZnzbDPgRUxVHRKhRb89Mw7z9U8J
Xj62aM6fO8sF7+RPl+e8ERxe17ZsTg8slvBPKhAAmustyb+gnjxwRPy9FgqS3pm7
G68B5R/bOjpSJHYzhA8Y/tW4Vurkk0hpS+ti6h5AnkvkWPWD0LdFNuaZ/YdxRXdr
dIDU+Nb5k9N3v6S/iuGjn17J60lPDam6FjKtJclXVkDZScygr3vum8kEPJnp3ytQ
CtyulD0eCfaAOzR/aXPAyo8sX+o35b8mCTZhN2PHs5FTHow8ESFh/Rhc9EV+t2V6
Xc5PVHgssueTjnc7qDI9SNJ8k4u/2wlhv52vIpLpaFFnI5CBnKQQqubHNc9ar70+
+KHEcKFTQgNr/yenYoMFKRY7sP6Gb4J9r188wjJcOqRBfnlcRao8trjwva5NBx3k
A2ZK9eoBzVliJ9Dt6YaImfBmVIMUaQ8tEWqa55nxbBb9CaRv//CIc8Wy3pSvHAAa
33OOU7t806r9sPeeboED7mCpcIEjSjJi6H6JU+iu0pPN9ydwAzlXeftb5aSQAlBo
VaBe6RymIO3qbT9mLdXr5cPys3W0TdCfEfBPweAy7O7kpuLk0sJsuLZsJhKSUTuB
NJaxIdia/aw+E+EhEW/06Q==
`protect END_PROTECTED
