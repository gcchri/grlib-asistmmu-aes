`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3VCRvf7KLJON9jqBvkyKxWqVtbIm4/8VGmp62tmjZvDo7qt35BeYoutKG68DUtB3
0Bn99XJUUf2V9j/IXx2OLczhmr5Dpjkq/uFee0Tg5zAsWa++E9DH5S6T6obtFkCT
hfEZ0BkJUV1fg/j7+dBA9baciNLy7ENpHUuNo1yh+UEZol0npGwzhiaPJ4IQ7b7q
Fl33wjmdkIchfGc4nJAgfe0zDgxELeic6gxbNo08+Hqd4T0QlP2GaUEouAAFmTk6
gkK2mtzGuUjehIWrWEjV2100SnCQi81jEXDgfvb4DSIdUawuFFKRuinh4EZ63w6M
qLRglr09EnO1IInazHyOVZgFEJ/9NCdCQVEupRr54MU2M6xBF0Xpw0szdtUnzWTy
h+bTw8JtWRbM1+DRTvuEGS0vTrrPE4kFz/Y/NM6El8qSdiaZEwbRSqw8xvveqHCB
TkjR1KIDaSXWZvsCZCcxJ+zs6ADKlsRDs1itQcjyX9tly7Xo9BqPAcHtasE2QHag
LFEieJ4XN8nrqMAMjj1XqjD+hCO2Zi5OOWia2783hbaQJOIeZvwoyNQmNBupEGHU
`protect END_PROTECTED
