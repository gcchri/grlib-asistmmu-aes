`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ih2pRLo1h2NdhplV5bpxYJqvn8zR7dbH7qriwLOsbUxTfLEKkfzQbnICZNDYeoEt
OSdg6+budKpJ44ZvOhr7s1ZtoqePP2EPx7haj+DNiSfp6Ukm1mKK+EYHp6KZ88a4
/Ty0tlytMtVGg5aiGVd2oI28rFTPPvlwmcf9Y9uukt8p6Wpu6Pc22ET/3YGIkvpN
l8+pPbUwRxmU94cYSeLYH5Nz2l3LdZlCtAamzaO8PfJ3DmAhndm4qxBJuN4zswUx
2hv+fKQXl4y23H6cN+D2vpOQ3HKNIgH1o4IOEn8+hSH0bVUEtvDsCDFtY+Bh7HyG
/x2+D/MetFEdiZDWc8iFPxERI+yi/bkEjkHCIMOBu5Be90x9N3bJCCkSJ/CjyaeX
wVcn7VF2SqkgJkpW2qiwhjB5ZKaT6AZRGRlcwNktfCs=
`protect END_PROTECTED
