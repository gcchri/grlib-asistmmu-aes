`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rtlqyX+lOzs+aa7rH2psneWuizukqMuoTgyyqVwIheCBMDE8JQj3lT8rF66RQ7bc
EGgfkM8sGZvFH27vwyWOpnvsk8B0MvUj4N3qnkL/Zh8jkKbbrBSIvEV7o98B23w0
AJ5RmZy3Jm/AJHSv64tIH46pHNb9jwVfLqj2ZRyOwaNQvyAHs7KEvWYogDIS7ai/
ym2gtKNWSb+f4Pp7w70pGY1nmKJGAVKx3mUbeG3EYuGlJ8E1Xxx/zNiRqPKfODsT
jBrfNyEBFBGEw1t8DkFzWcgrzp6kouP5BA8YDWi9EbbKbWLRaGP+uhGLIkcORmYE
pNcD7EWgiEHpebKSNkzPEDWuBc5VuB/NXa8ISPt9QKIZQF7XxIKnWX+Ux4YoXJyY
`protect END_PROTECTED
