`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BaSr4xR8tiZcuixWTJ9JanUXffiY5EsQvZpetlTtBe5Zk/cxEecs1kYFOqqUO0h
E4XYEylCv6xYcTCzktIglzAub8y4gT5QayxU9Vc+LcT0ehx5HjjFk+9YfYeJidEF
Ik+vCu1nevcvLf9hAc8ba6w4BHXQhysoi3OLvrbSMX+lJ5wNqaV30vXZi9JdI1F8
jQ7zl9S3NpYPK+Bz0ENVfYU+wVuYzrKtoLS0n1RrP/Wk/i9eQG+3grmRWZb+6nPA
dqvYR9nSN75j69zcgwkT7ny1JJCU7stjU0cwOG1UJNk7FFwaEdpe8vG9E2dmE9lb
9ds4AkYDu47qY+OAJr1ePV3Glr3J1JfJbt2Pm3PIlxozBdyKRuzqlDucfiJzoh8b
`protect END_PROTECTED
