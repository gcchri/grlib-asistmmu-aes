`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPJ99dqyndavmkEditd1k6s7agRV6z23KCcBP5UpiiBedQQdx/T7R4apJ2Qc0YBm
9FXR1nOqkSpaVCQm90jo7NZYwsyaR5BA7R9gLRZQvOyYj3TNvBBZBNfiF77nTzc6
bdaQW8ZA3dn5SkHdE5KG8NPr/I05km4e49HRrFbO1Ut/ohDjl2EyEYgZmVyhbiOq
x0c9Gk6hj9fp5uQYM6EfRwQEYf/FWjDuhdMIa3Udu49lg56IiSWwo99AZLwfc6jn
uVm11Y1n3/EjBwn+CqdBe8gxaPvr2A3s/oct3T2E15JGUD9l0ra1CjM2M8jJ5Dn6
xP22h9EUCpKnAvD1u+AmRIFeW4WaUSI+9M2I8eW16ALGtUfarefLGDAyl/084A0Z
`protect END_PROTECTED
