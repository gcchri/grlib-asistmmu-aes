`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TqeQwlqRypyyk0+McVBeLqrPbwsTqXh8unyQLEKnfnPPHCY58ym7Rxyzo8HAyrzK
m9PfX+Al1V0cW3009dV7Daw8CWmsEF8YatFiTvKwSjRBr6NYySSp8lfwwF26+WBq
MlgXm0cBJttBDsQ2yOifD6ONwlYVLlYqVdftLFd3KX7ADRQx+t5wyEHuUhAd2WkX
vKyvmL70yygr47fCq1StzCg6k2nGXR+l352mqeXxe4cUuByYBFaNvH3WR9YxDnaB
xZfH5F2kCb/KO6Q7YsPk5/BZWLe+BxrWVk1VhhFnUk30QwT2LGRIY/ll3heJGSX+
y415uhU8t3SltESzVIFNgSOZj55X1r/Fb9M01V1wI5LePb4qfEPgA6/ymf/ZR/z2
0npwKSw00wFziAu7xJzMZj7A+4MGrIWWrHOpQO0Z3oA=
`protect END_PROTECTED
