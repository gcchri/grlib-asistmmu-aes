`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BY5jqnqIx+VF47x0QjYruz2qvInDy+CC5VKA9R7Y/6DT0GP9qWU9bRAjgIQ1VinO
LkFWppx9Hpvtv4JCC1YPIaW3sGZ3NL5KWLZPalvgPSfrqJ6qXDGPJhl7l2MQkg5N
YZXiZbbyKoZtnnX8rcWtnTm1ODgo9UC+bplqzR50Y7cgIlrIGk6ghSQ3QUvHuCVx
bKwifsLSako4QAQzxvep8ix9eWUR+xZAZxgIoDcm5zprhx0mPOcfsaZ2RSQcBnW0
JVsWIIrl322Uq+85mklJD3bQf/W4gAy84W6FN5ZtS0VoHC2APg2WfYPkZP8qC35y
WgSZ1gQwvoQYt/823OPYu1btzK4a86M/L6PGmUMdw4pU+CHO6r4be58zd4VDRFoc
45ikM2YsECpu754hfm6bTsX+ZRRtXh9iGEByWwF90jf3JhhedkOagReQfXInHKY6
QviIy/S1zCHYwCMFAAtPdilKvCSy+u16ruzZtHrSYx4A73p0+4C1t1GHx+Hhrhp/
MzLGhLv9Ml3Hg5VAB9FdMCHYNcvIotKN5CQ4cUp03ogI1PsGGF073TpRC+1S4Z4/
R/uHEcRVRW607f4yd+JbNxav0/2EPedHfgmvbNUMKRg=
`protect END_PROTECTED
