`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+S4jGDN8AuEYX6I1w3RxGW2SfW+HjyU27/Sow/rPHLSiv/1i/Te95KmUai/SWTeF
PYQwc+lnhXrPT/IWV9h18Dva9Ow4RkoWbw90VzQ3SWOKQtPLVgvpfS/0jWyopRss
2pDZAECVbsM4UBoqy1/L5bGDyPfEDOyMMTY1MLT5UOcQzid5jn+tuc5dLYiS1TPC
7nlvx7FS8zHbaSGeg2CGnZO8iv4CLd9/hkHjcc47mRTeE2Juq8KLlb/r7lDY+NOg
/0R9ACId1QqUXjUgH91ujpQ9bjgb5F5RVV4/Poey3Fi1X4s8Tw0MbjUQ9sDSxm7l
BJTm36gmxtyXPX5RssEWysZHgv9fnhpUM0fyoUH8GQa0X02pvTPj1F7WoSBuLbVi
ORUwnpLOANv47s7AzZlRnZJl72Dzxj0tULn9e4FWT8kEydJFmwy0ysvKo3AlQpoJ
HK1PsY7B7SwTeCv/YLymNrfFkwX4ZiX316E237HmCKJ2IKD9ZMEQVOtlDvuQlyXv
n3I/CqA/c/WyWQgECiGt2e3Q8iOrLexW6C/8AGe3lCD4nqwBOYIcIqH8Slyd41zz
7dEGxdkTTgo1N1UlG9pNmNwoG73W+6Zc4/48M+Ps7f3k0ctkS3JU3quMn065D3l6
/ZWmJXBsDl6kMfYYyhGmjQ==
`protect END_PROTECTED
