`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVY0HiPf91RuS1dzTFTXOQtZX7PWZnVW8jKJMV1ekYa8NTAz9MfuAMNcC98osaO2
OMMIBLVL/4lcg6DX+Q/ybYcvBK3+lMxHKNJgBtKiNB9IcB7UcrIGCptMqqyZoJYj
1JGDQ2nnDoTZ/v67KhBL9Qqutfxbsslh7FNZikDmuQE3kqTKH8wDs44OubV2bU++
xfG1BWE6np2vLd0d93qjdIICXsz1xS7z7fcwI0G6ONb85l2lrnJ/sFtiQ9svH6bu
hqnydO+j3uVFfya2uj4YTF3g7iUP8c4XdjV79RBO101rFnsOlE2SPi1w5355df0Q
ZbXKHmYfRdqAQuv1iT7MvmganjwbEAG/8gLQCWgSiQHsnjK4+KxSEkwh22xU2ejW
LGfjXlmHhDC3xf9g2IA00deKzV44IH673XPGaXJbFpefWOQfF7j6UCdmi71dDM4Q
eKCMKe4g4ltiQQyF2nFh8OnmfO3heXjlEjiLiv+Csm1VTqV1i5AlNjBPBD9gtQTn
bbl9ZQtHy3n4XpNT7YnCXaOLtSUoLZsGAuhwmWvc5TibyY1XWDPv6+I24Pursmlp
lwlKHf8WKrWYhFnly623Xc1S2nVD1lFzpAAx3T8XjA1lu+hwJ3jylG1DL0y/fzyd
MxomDZITapi26nqkdtxRZK1o3rhKD9FgQZnFvPCqvE40CBwm5EinJ7mOChmfut5w
FovjaKBf+V7iWpbOtx3OLp2DWkjLAQYmI3vdCd5i4PtoAhiYH1L3oOCvUHF/chii
lrhdAidiIUVA2I35oebjxNBTjIASRkpClmDeXC7KKRU6yAhrauTeIdwqDZznh36V
5MvgnCPR7GsFsGkmdxa1xyPMp1btFcIZG4ldCGCD1btHav6OZET1OgcxJF2bZrZB
wU0mNzJ4E4N5fL0onevtqxu79kVxlIcHMWeskUXFXLLCBqjoO5xWVQaCfE27WBlW
pezyTvIMV3a6sKnt3/i33sJ3rmK2uco4gfZWpb67Wn3ux81RSAOkcqLTZojenEpb
pMtxJFEieSz/e0zvJKW1mCpdW+x+F+RpkdsHUKdNJ3L00Nj6svYBoVaav8EjuhXZ
owUP4qmHoCCM36PGp1U6aeekoQVkPqG/J5rWpTZs7MNRC8V8B4ot0fHS0898Taam
HS3jIdZ4wKUp98p65BMi4FUBaSIlGc75E1A6DEwXWCsYA0lqUZNkMK/MlJSiPjT1
HSZcQNz+p+aRzPaREDoZWtohhI8mgmeu1SGl2mIXOI3xj407vkCHJaecuDoia2qi
ngCFXrm+lRUuIHnJgphoM+3crwSyAW08IOHcPXYwUYgBVmkheaxXRaPP7TdA8ZMq
kT+zOT62kJI/Nv3EFllnqskIx/X6j2FwegmKQIRoL47Uf6q7MT7KrdpYMQoSQ8+k
I/AQdOUjrPPeQ2SfBRF4S459fkiZUBGHvt6h+gp3fg7vtObjCJiV9ZXtBgoWKPxl
eKP/Fa+6mFIth/ZFI8LQwN3v2G8Gf96EsRQdQ6/GnN5WHKtvcp2+FeBBycKCW0La
4W3ZLmMVt1/85IDlOJ5/qjMxNVeg/zRIunEUZb46tqreSDEuEja3rOuMphhQHaEG
iAA62LK0OnceCbLKPavt+f+FH8RP+DSd5UfF2ojEnIOowzqX6eyJR0bkbiSGaLDH
R3c+rV2WvIzZUhUccoxEN111zhgu7vHa5VKRMaauiUeNDLtcSNpvwUCBI0TGe+mC
SsnPRqStF6wSr1XpTrNc4RdqcBx4g+ckkMtwsYNmnwR179atT70IQT/o8x9vViSB
b3UrdBYoU6sqTzJ7yuyAtVT8ddwYJ+8nsdQKuWvT30ysvRPG/YExVpPJLUk3kNq5
EffgOji4C4gBl1yU77+1YjvDz6ornjncfwsWoSajYWDd2JUkVrYvXwHzP+/4MtEL
dOe+bd8sGXh1eIFH69W0IObeF+pJosP5FBa1bv7dTuCscI3YIJYfVaVeZwLj2T4m
JLP3dkAgBXOe9dl3cpqlsURg/+u4HLmrRjuDHK4PAjy2c2rTFwRWW4EslEO1Yjkv
uKRJs8xfzbVRvahyqPI3W+itZkDUv2KjtdLbkc1wlqXaiOzu98M0aOXa3GXVuPRf
eAEBYKDTLqj2F+7+tzL3Gb9ZGnXJfkwD5zf4jbuR+cyC6OqiMV5iw8hKWn3F4BIc
QiY5arS7xSbVM6uajN2SqPlwsMoUkxfSuIlZlbJHEf58c0J13OBTP7yeOo1jBRmx
TUNzZ7BZyBENjCCzAY+rKqiHfJrdB0URd6pozghCQ00nFndxoqTlmmZk0Cd48e0a
h402uSeX2T1dih5fFaFegmmLkZDNeouN+jo/Pk60DA942EP2aatU+5h3u74Aw0nR
Ch3tNqaERdVTHBtLLQycAm8NftJSYHcc5X5DEHL2g5zV0eVfrN6FRM1poE/CNknC
UItI+I7m3Ql9hie7VAzXFS277v8md0TmxBDYqjdS2jVmHNS8c6uNy39kx6IfxqGK
tL8X5PYy58F8iE+6qAZztPzwLTdiN/3nDYXDjdavPgEXMMEf7m43TgLpfCy8hfol
qC2nbEl4DNrQxMwtRoPNryiH9TMHhmOZvANdclGUa64oy5panwKk9t6uZktJDtw+
e+BtoAUdHkS7rUt8TU2tX6l9WRbxKuVxOoAfkr7wkHYrE9Dnjt6i1mxfcAp9lXnT
M+R8i1W2Gki616iDnS2QzQOGiYkXBjUV2GEtVrAQv4jyTVCBHT6lXJNOQPhvmcwu
KTTIVwD6e+z8OudkvdeyYAZ9SW/Yx0IUmZ3c+Q8X0AGnJdnj+Nw9lH2zgyYkC23R
Nxk3R71tcYV7M5xZjzZ/Q7O+yC5GA+DLH2hD0mOvCxgHMv18kWABnvy6/tuETU65
4ZAz+KwK8JpZZetMhIA0Gzw9rwp2sz+iPEospM7akzQyoojAAwuzas5vgkxDpvZq
LqoSkSCeCJT/M/LaWS/uEQ7plguwsga1tUy0pi67bQf6AqbKclhxm+AgDEt6tDls
09K6G4g5fo9ImBpsTbmBlL/uevt6EStN6EtPFQIoFHToyme/tmhCoz0cQWgdLjog
YvTwztk/LyruEqyeD1wZP7BhfUMUmaXUCVSM9Opj2AVOx7fgWVILM9TDzX29xDqC
WHLigYqomQCTQtAN+ut2N2LvcsLJMrbMM69ZccsgYfSF+8ob5dSJl+zomgkjL+jg
9irbHFtRODGkwCQM657iBPMDWpbJQXSbvI3hSiJhEeVwj8ZrbtLuVjXnrJnDshc+
oBX0sICedE/qjasZz/THQIKMI0UfF60IITg+dQ9RLoyARzrqSayT5hhikrw025Nl
sKv0ixfrxgqKaswP1ygUQDakpkl34pXR40kW0+Vyu4EikUs0vHlwIrsgoMjnJol3
RR62zhcdOEw17p9rrzWqc2QoGJQz3vze4rNcJENl8qGGrrMomYji8C5D8jkUiKbS
p0gih1moV1sqKKy5EgvdS5QMkowTembhxcILJJ7t6TXRg/1apERfbzjb3NjdnTHp
iaFP7VaWRCBgfRNuWW4jJvpcIfNxK3ekygFrKxea8GOfczbCQkL+teAZYxtN6dcJ
NZWLEvQhjfnpsOjb3FwsBAqpEzuAj+x9TD9fb5Mtx5+YanLqRm1nx9kHQ05im1Su
ciRX065v83aK1O0HFFoRDYY+v5JucPUV5+PcJqv8EgJ2N69fWu6Z5cbxllCRAtRA
uOX7VCufh3ctOGwd/ZEoHNpgjuASzAj/G+/hjNU4eLTVBRfrubI3rtSj2qWQfGGe
p5CdP55xpNb2Mnw5ewTs2BxzG3Qc+FE5XawDThHWrH1SPDUiSwV3kTklcaLOvpT1
7B7cQ8d7lCP2McfBbxPRpbUgjTzcTaydpegDOuTKrIaArhmQtV8KhLF8bhr84Jb9
UhD0SR+6CJkfmrojA+PbpZ3YsKdp/SgZSw0l4FBEWFOpM3ikopIARFd+iGLsx4HV
eT/hA0Flh51kLbzHNzxfFJaVvSU0nM4Kn/rt+jE9OU+wLtXh2iO1brhsaiGqJ023
HSfj84JxffzqEbRuLgvffZ9Jt9ZU2wWKCEJ4tt5zT/x2r5LnrMV/KkzmevefHp2T
lwiIJgS7bV6SwCEwM5DkngGLhiIISwspqKpKI3iHQEU3OqlpeLBfji/EPsAYRykR
zKl3n9kOeAmrIWB1MqYyrBzJBeRWrEzBcIm6MIaoKVl73inW0TXA1ICndePeVavc
4t6BY35HKLog2e4ZXnVrt00Jjgv/cij3KMgZsn12CyHU+luXdiQOuSrgpxVVqmmC
xy+9Pi7A4IdxD/crQFEalaLhnOiYIuHHsyXD54SakmoexgrNfrzHXOAamBssBCv1
HKbjGUoiw9de5GgzDlmk/14iz8n/zferkx4afRQVYu3rg1ZSs4OalQTDP5jTgXXD
nHVpC0q6pBpoZgbabONyRTWJ45TZOnyFe9PQ1ECvzs33FAIXq3H8SmRamWIDL9CG
jH/bOpoCSA5XpJBFO30QkgTE59M2eyZkRUvWMhCTX/WskyvSfgQ3YJiV9V/bhqtd
pxeujVYqfR6288R+KyMJN5l9NZpDJuE+JpP2uxhUt0mNdMuGgHWI+U1mZNm5sUaE
GBhUEvC3VGJ53tcEopovbB4xtaGQQatPBynYr1N+sldo1m8vLaJ5jIn4EV5IPe81
pdprSSzHsJdU3THvwdszGVDJRnVh3CZq8w44OvcyqxM6CvDqacz3nAfLePl29z9z
xJKA+fCQQrWTV6FBiO+2XMN6n4pgI7NxrM/gjJzyW+8jamFh3Bx48e5rvmhhrIVv
1PwHG6Fjs099ufCpGRb8NuNbd2HCxx0P79e5ZISUeyIz1kKNrtOGv6ZDwGyoTJO8
ZuOdg6ahv4nLwTtYQksL/6N+WOJwseA/iV+g+Zw/QFJssG3j2lHcRT6W04u4FOLI
YxsZjuHUycNFuQPhFW9ruzj8aMwkHNCc8V2FTOjLRvfRECcuTk+Td8tjOlux2YXu
i5k3otKKMzW4yxFeG7+QGrd0X1KEa8Nzf9xqo4FvmosW5/wev/zLbTSnJm6eDRV4
iAMKVLRAfWf8VY87jF+ccxfUV1o78M4EG3M6/Xu/Ui/zt3vAGtK8PnBR77CU41ye
hHkeJiQIo0idxn7Fb0IcTxzV7nT9/WxmMwElO9gCkjQERb4Cxadh+Fs+8icNArT2
/fUkAat+YXd66d+xGW63YCpDTKFghQrf8tEBwks/A8qCr+eHzuNo6uXFiPeU2OLG
vp04KGzOg2DDz2eafeT+j8+uTPfR/NrqNMo7GRLOMEoEUY3jriyAY1NW+KL+ZVtn
+djk7BjpgDbBju34Pg+zg/ZVD8mASnUPwHnEwstOuES35B/DFUeYemLlcJOcXbHo
4w6UAR/kpu6M1/k0obAw+yacEea2rD/HpRKY4eNbPujJlapt7Ts/imrcXnuPN0U9
gFr7l71LSuTn71Y/v+TTLaCmk+Pj4Lxq9AB/iyOivJYsP06vQeLVZKqY48CYnVrB
RkhibpTN5VSotpyCzcW9XT9HxE+MGdTekCBO5LN3CzqMe2/Lxrr3+Nn/dknYjDac
VPUyUkoyrjNeV1CIDJvvuyZMyenjdqAI861gQlXktutbOqyyJOnSOetKMZzbCjlu
YW7f8P5JXHhMWXTaUp8tqbBl+QOqkST9Zt+Hbg4OmWaxIYSK5SLzU+WBLk1HUkZY
cQq16PcGqGIYvf8t8yOSuOp5gYCM9+tXakXKnCCkN5aj+rGq8KT2Ui77yDt4H++7
0mdSw3RmTLKHratTnbooygESb1j+A0NSo+9MDZflojnetJtnCh28dQ4mrsWmkp1d
KboP9mL9as6kxFBl8/10vqSuBxeeJ572sxoxmwPbwgT6iMSASNJZSBKzjtLHfvn9
FfLitJ9HCv37j/azjNcN8HjSuB4+5lcUt7FggoZLGjI4QqVg6CZ3MiQseJNZ8PrW
pdNdBQo50fr9VQ7t3mdUZ0eB3jdDsO6fIKz7zMWdh+SHr5y6dWG7GTgZAeucs6fO
3kvT9XFBTAKOTNYfRCpsaci4IL7nEVKn7EvqEteVJP06b361zMY9yv2A5zhq97kq
AGZ7CZ7Ee9E99K2i/PBH+Mxb6KNuv6Z919uzczNYwqKX1iyOUgZLMcRzEpn4y0KO
LbD2XJQZAbN1CaTyWHe2rSoSdiuRquW1koDx5YZDydrxsDC974vHp+wzbcDmIO39
KW++vlEaDhZKdu11ElBnDJAF6Wk1oL0JmJDqQiDyG70JKhp5Uu8e0mHHtS9uT6xD
MdNvJzBjtH8UkQstQ/9v1zdGCTbTxGlub9Fk9hd7boZ4IIJDl5MX9KbSGOv8BKS+
cuMhJvffCEzfCmoZp1IX8JKV/xl27Z2xTuC563Poh33IgT6lBX/ieGPrDid4u81v
Y3Z0UUKMgGxLOtLgA9pNG2ohbt9F4jguVW48kMaGZe43EkankZ3Z2qPIV7ru9wZD
Dp4SEkUNTLQZCVO5Tp2sKwL/DklogqETEwiIRtbKBeZyk4pHCFPJ2K+AgGHIVFfo
1p0k78831XPzKebH5JrM4GQmKRX3Hm+GuScAj89VvbXFOFbgx6WSzTYDkbBpMSIp
npq36Dq9ei+GJDklak1ydwGJbAYaLwh7T3RRRs5PcdSt8vWQ3OsiUcBHigkTr4qT
4PPqsTSxo9r7/3jO3FZB0Rq91FtwkIX9YorkZUILO6IVEltDoQOcoyu4AAFeT6OJ
wmx5yc+7r25SgzEy1B7d/G7UK43N0CHJWMbjYt9Wb5/VL9SXu6suGdF5bYGJPstj
JyZB4P7cfclV9VjWgu5PstSkZihB9VbwwNSM55mVIhQ8yhbtvJdwYlO55yFUYe5x
pjAJwVNOAOwFNoq2q39/VZktGmqes1K+2i9DNZKWjP99U8DbPqVVfoLliYLrbgm7
4deDtfPXBc+/J5xe1WrXBICFV1W1eIRrgLn3C01qfRyK99ohPdzM2FDApFmYumRS
O9SFOJtF9TzviSPPIf/+Ndh+LdUnkdqAD2h4B50Dtmb2N/LDqdX7xWWjq7gJ2Cpa
mTMa5ov/YjGo+h9mJ+wd7Ly3Tobd39YLShCYPzXj7WDaD5T7t9nW2pB8bP1ApYF0
hBkd5hlmIMQsFmhnYPNnab08nH1RviIs5s8bq1WpsAkaeIZCsrhI1Yhzzw1D5w5t
91dx+RkPyLfZDNUFqcPFBSP26ZVQS7gM2KhxAI3IPmncZKIQtYQWQrJZVgnDRTJj
+ZpLbvqGmy9pM9WurNFNumIIixOcICydGOnLRLHt7NBUyaywQuVhuHk+lc53y+K2
vDk/m9C4VO6Y744Yw4Mq/L1Fn9x7QRHedmxUzFK4UlOMmOCu7ytnBlNvDR0QEY67
z69IPogxF21fo9wEi8blC9Y0xhYGQTSr8SF8gL8uPR2KHnqivv9uHV2Cfh0C+Sjg
FOV8hwQHULdPmjYTQpLuplnYZ0IgsJPx/dOCEPDkWvWUqkK6TajAxrtogzdk5I2E
uoWXIDmjQVv1oHkE+YDogCvrRJ9cxK/f9Ri2r+b2om2vfdqyXYV1sUVqIjVI6PR0
c56f4eRxvuNR/5ZdH8x+dLsKMnNmsvg7dMaxT/mVDi3AvQCvpCJCRed9J37JI01W
0pLkbKbLzsIEpb5iRU1JW2gxjAMMAEJjaXElvx8jMdJWsnOEX9lmMRJTeRgw8BFJ
H/bsXpIlGobYCTuneeKtKd4SwfzJhxriR2PKg4zu3Ytbqa6ahuQHMmZ3WDg0OYSH
8v9lo5Tp7usSNdNwLHQ90jynePHaAOhvxkpK2aWm2P/sGfcom1/Q7JSrSYuEBQyS
7xeDsNRKZgjHrXherbL4sn90UqoR5osL0rsbiT7YJpIlGfIlHSHr83ryXftyRoWS
dF5I1VWW1bmw1pU/dwUsETibx8S1RMRPL/7kdKnDzmPiXuOaRyeKmJ8dpVr8gR00
o40DquUCDm3M1Ug+3ZZdv+2jI0KiybRIT3V587gi3dXaGS5fiYyGho+apn36bP9S
q+w04bATPHxMNgglwRPLwW9dTRiVAgYEbm3yWvK9ivN21GKgr/Iim+DtYMNR4Iwo
Dt0Fd4xs+wisNIU87SC7Ue4wY2ifLe6YYc+b1FMWAMtJ83RE9W8q2P1eplpxZoZx
xzyxvdo+L7gsbylS11J84t78OYsSMThyf+Fyg5ABOOwPDpj/A/yesY6Oo5+JrKnS
3bEWCnUPiDteismggB7ENqH8C1GXeMoDMfTrT97fo7M8kPuSiihn4Wsjx+aJ5gvx
eky2djAxwcGocQb8irUDkZdQon6XtOxtpWT5V5xXBRdi76CjbxzLW1VcnWrncl9I
eFJ7wVJxNONRGdrncc7RgUIwpqcjC1zQgZS7ykFceuwYVY5Odw65c7ZswrP4AuqT
CRMohcJhCjSK7caR25gs6x4HmKkox+wt35ovRnROPegBs8/Vv4SN5RrrpGYywSTN
ftE9joxDDU/V3KXAe3dhNrBx7tC1a8ucximy1taM4hm9NKsstFATQ3Hl1p9fwycC
eQRz4789+e0BBZUTZuQ02TyXC4o26JoRXTv6NGBV55C71rtXIkutAXsH73KY3iLK
ergbLVS6EZ5PI8p8JafyY1vGjUf21azhLuFEWun6/MHdTBF6xuidIOk0MlBm/5oV
aGUyWxS5h/3ZHG30yGIIhC4XINZdp0RgXdYdcBY96RCjKkj88uwzjV7XcodTLYZu
f1ZXxe03iLloQCJw2CMssAMBxUgdf5RCW8rb/J4uJQCU8HACSbs4c5aMwC68ZKlu
O0Ae1wRTboNr1wYqGyGEpW0mOtfNaZ6cYRpX9Y0sFQkQS5kdVHWeDUoQIPRonP+J
jhxzgrp3xRImbb14VxiPPBLswAnqL9FpKuamrEZT3pAMGD5kybW+AbJbxntppuDI
8Ls8ulYou3+8SmDbpQCEtcvk9okbPH5o+twZY3k9U2mUkVD1cFr6XCORPvbGoa16
BFuNRpVjJ2jtyVamCjrl6Sq+x6Ui3T76RhrQKH1E9QhHX5Du5MGh2ATM9ZzAtz7/
WltrS3VQK8/ObC1QuDUEhFHs6CX9NB3wyw6Vp7NtuvVTjpY6+fd9eSHBYWujUjjv
saFK5DJ07eUPb3KnDU6suzLVs83hUHNAuIGhwDyztrCyCDJLuEObbNs1Kakm6eHq
oCXg9oAlCD56roVTk1QKAJ7qvKyLEoM2co1Rq4npvMwR5ZUtxtezwdO2l245mRZf
3bTP8UaLCYMm4l5PSekVDhPuaqyl1sAbXCkwq+LW1EHY1SK+BWdblHkcoyepGUm0
tYi0OOJFel5C9l2av7NE4XgNvkuW72lNijOHHC+R0Duc6yVj3rKqcI/yeBhwx6Nc
yFkxHu77wOYpxj+iH8VgJ+ZzEbzAp1gLCCvDdOgRxRulOrYLJI+TF2XTQE7BoDvA
BIUPLmaFqfMEFydkdCeNkdcCAS2VTZpuYgTCtz4b13Ga6Wd+anMMRc+qBTP4TfkM
NV0Zwxu5GA0Hz77mCH012uR886MVMDtnNi5vqfXDu03kmHykEjRm7qsMP37Ud+z5
H5p74GzodEYkV7UlDECtlgeVtum+bVGY8Ee0IJDWOl56Ezr6vsQklUN7pujRNyB9
gvCJL58J9qU7z/YTPq9yRbnOY4rJr1/AWX9SFGUY2RLcDca2FHEvrqJwKl9iTFeo
ysakJMv/VyT8xU6d0VN8EqP/YLOiQKS87C/3PvvEZhW1cpR1jtQtS66v51H4RdE0
aZL00IR37Q8Lm3QKA2KBTfhlrUjL3UXGqtOeheSYwY9+fXoof1q0QsNDNjyQNOHV
YyxXACXElCV8Cik48/i2Krmgb3Mypodn5U3Ctqy/V4XtySFKcivaoF0uHSWdUuqx
fXZjb9rm+lrDEGnVITFetSMBaQOS8kiVxtcSPs6JFxxVtJ7SZElUhIiHmhEQYg/7
IhT9tbb3U10WMwjQtjWU6CeihVcnD3kuULmpM4g79aMiinPm4sJOUcZBCTw5Ogaz
6eqAMJvhC4y8Y4dHvvAz0d6qAjHo+cGA+3JrTJo9doUAISSqL+rOl4Dose4yqRJU
xgesQ9gvg1k9eSA5EYX5fxJ4gsCSUDKoa5JyRKvwz5KxbqAKSZ+DVG/dk2dCACot
z6B2tLP/5rHY2wdxva6+rpoEjGMCuIj+1jkkcKaZg+/XG5/eW+oV4GsEOoJBVA1P
bN5n0IeVFbq2/YqJFIF8mXJ924lvVdZQ0ePyo3VNZuuinP/gr8KoGjtVl5e5PJsr
eq4qLneWeXtRZQnNO9UF1ZVodC6zHvSlhhgF1mjVRbrjMu4yxzYJQHSg42FkHrm1
J5PG4qQbl7vZ/sNqIVjfQgkH75mC2LYDyHjgdBkBzZE5x++WSVl9BVsykl/oxbWH
qh/RGGK9R5Sr25OHgPBa1P3or+T1pWT6oXTJ+0ZZyUkRU4XVlGBdGhUhSI3aSm1m
jI2mowwWFf17AyzaJYpXT/FlQrTjxG+qmtSPiNFbUFKqJ6xgPOXkSCVHBBRLOH88
1gY9FvfHAJ5E2Yah1A3Te3x0RbJ+2tH4gT9abHXGQU/FTMkqWEI1HlccoBb0+ktS
ElqELcnUCl0TVWuZbiae0YqHzhWd6du3JWqVYfftlktLaACG+CX4/jwybOKyquZz
ACLRrxKAxW0l+Qi5bIMxwWafUPlQRlNjV3gHJlBrSLwaJLazj69lPn/Tu74zOF5w
NVurNnlvHBHbk5C0E5/Tk3l8ZLJCyDpuBxYP5/rAVZRA3vD3ejk/6XN/lqy38CZX
dazZuNRfkBRTDD4etxtphHzSQoHiFZDvDVhRshf1AxVbq2+Zzut5W2DvHspCxO4D
44jbNDCULsGgNG3A9HYDfwVlrwMQR873Ssbj5DCO1RQak51RRvX+dRFSmzKy/km/
QKaaQF4XYcJjbHeI4qfqW5LRPgyoQESgifL9NQqeSTdhojL0p09RLZUtWrCOxQBk
3xAPj2ffCwkMXNnIE7pEnjwJWyVqKC3iwKanwMZwagcf3/S80Wq+7QxVI0LRZ7gy
VTCIE5pXS1i7clL6CbG6eFnQrC8n3fRDG45Cv/26WOch0xWdL7JMcmyLW1wRF/8G
0cA38WTvf9gP3mes+xQ7OVlySikxQ/rDM9XvD4Wb6lniTWYB+KMWSpgR75j6sxp2
glgwxmErWEwNpnqAvxejRclt+Zg5adWMCHmNAMhsbfxKp4XZ4aX6qXCu5tPOzUxQ
grHYmeBVcymh9bhIYXEfQ8B8tlVk5cNT6lsF5yy2EsGwMzuqzkd2pzUFgAJx2F+u
0/7D8P6YfvX1EvyiJKt3W1FCf68rRoui5/0usJINsnYDMpPVfLB/yEOieYj0YFrX
DxzjBl/eWfaMTnMaLHrgrrxdMtNOppcUEHUtHL0/Z3iiTBk5YiK1pTkYrrRIuP8S
TWZQJTnjNHm7HmGCNA9fLTEVjeqaJsTBwYzWtNejK6pc8edqwxAPGV7kj1vg9jeu
3g/FORLucjcVnHsEteks3cBvCWAc3NfHszKZtIsaH4SKOI4POTCIGFbmq2XOf6AB
OlyzoXJjxz4iZSUX8V2ZO70aT8/1xB5K2Lpd6s+8UMcMU6guDRQ1dSXscjMT5SYM
YlH+Nmx8MMcqBgkyfcP5GHkpLm5OzQRUmWWDoULjQBNUpxpwrY/qktYfac+31hg1
NfQb6AUNCCTCMa+B/e/+pOwwN7zip9d0mh886g1S0HWnt7rK0Udp0uRbuCvsLvCk
i4j8LpDsiNtWPyir4+dPnIVIOf/T9uR5/a7jYcvgidldkUNJsZ14Fo4+tERpyYdA
ISMGaPV8Z1Z8UcOuJjdUtCfLfRicgom9IjzJ1dz/S40NuMG33C6CTvH7sKjY317I
LY5xZvRtcQyH8T0TTj/acR+cUm78cMsZHf8Ma5fmNyPM4Px8WvtWYxZ1b95Jqdo3
io5nJTdt70FTR8Zsml68pa6cuB9i+Rn70wHGZoiBdSPtkCNz75N9mtTk2khlw/kR
h3+1VWR4Hn24MWetTZo6oc9TVmE7C1Qc3KkEwLZO6eKTRoq81bRx9bSkSfDgl8eR
ZR1iT14dZUBQeFRKgu4hWrA70SNASrpmitM8NF7mXPuzvtdJVEcrF0JzrYL4meYu
rUilPq807tr7Zh3roYcn+QhRTuJimtGAQHgpu2gOtSRkXf5aVAs4KNq/p3cwtqzN
3AitkiAxWOvvD6dREhG0u0+OxxKCehLEqzBhYp0g7LdGoY6Xo8iGozYkJpqZwKAN
Q8sSwM6Q488c3mMoypkJIBq6TKrTEY4qzES2ZZJrukBc9NxadkFct+Ww/eT3oh6b
rYunCDx7ezS2tUDkxWgdHi+F2Kdb9kyNWu6/s0ktR6OFhNzv+RNFGROXfeuOHqaa
xUL7lw/tQBd6wHDDrfPBael1TxiqFoSH2XLGMu+Ba8F7OL7hCYYuVRp/aw2R/MO+
tZJrkD+hFkuFigy/U9pOP+ROL7UUZQyIp/0EecQZX+c4G/rAKAM0vu3GjWcJ+guA
Kr8LkQiIYbc4PWhtPGukjLX07JXb8rZ7SJ8uiFgdJL1mPG5pgI1wdRqYW6qioaeY
1oc6gwuJVCDz6PPQMF22CnZpmt6lx/m5QMkPuj7/ZtaeXq4bep3ijCAQtv7AYNkM
Ni1T/xnw/8SnQJsqU5K2m0z4CPvm03jinGNr/aOqgEQLyqXeZCJ+wUwg4jYFmZlq
BTKvKLu+5mHrvijewOznsp0+PQDdqQckwjdJ1GjBxMs1ghr5xo6ydqVWnKsnPFe7
30p7BAgysQ+IdQesTcaFjIQAVHyfWpYlI8Jo3n6T5nW7hHzIodXfIEriHXJY/0cG
fhMwZ+rjrVIL8O4y4OrGlyVQgyhyZrpX8ZZ7+wUZfcYS6dnlf1sK4slRU3g9359v
uAjG8kFb0onVd/nfq9aXSDdcYrwsH1tN8B7yzp1P19veddYFgfjx1gacT0RfGM0E
GOehH/nuvoHlCNDJRyy0XrapWHqALt20W6Bvec2tuNITLk1Zr7icYathFu7dAkIb
1300O2EsnYvqOO1eos8B0XZGHgTjTxo2IVNWXStOTkYFUpq6SM8vJsgSA4g3U/Q9
IkgBzqEDIv70Nwrdp0J+6+i2j/q+GgpNxZPIAftYNde03CtSWA13DWjq0eK6gOyI
/1XDnhZ8brWLUS/OKMRVP5fR9UtgrVcUAfyly6lg775TZzfBucXGpcy+ekxNlgNN
cEVej6laE3EPfJiW1y2IijMLpxn1EWL8CyLd7FsfdVNrHodY7vE3wX+0KWsZVmvI
FpSHdZt3st6SR0ewcqwgeWZ67OwcpKbuUPGkB5NOcTchklk2qKZyTvJZuXD9ZJ7l
k9UxhRV3GoJsudNM1hMbddOKsIZizZJmBRmzY/26/ZP39/tv09yVoGI8/LU5GY0U
OyriiP6DoThDdjTKiPWbmIQhrz5qggybjURu8zzkymiE6i+xAY8WpSspvWi2m1EF
BTOJ1doTpcxXdmy/1J/jx6BYNQ9rKZGthiAIAW8xPu+2DTrXeK+xxEasMnt3TYQ0
Y3+2qIa28lRub+KU9mvBZlTlDT69mIVm1ToNEhDsJy79YWEDI70457AWDBPJQ67N
+PSvcpzmA+0ZfeKM3LhAUaB0d4kxl5B5CIk+FCUC5n0BsR38k8T6rh/AzBQDDDmo
rTL8KNMr7clymXbaU/fhRDYjvfrPMj6Scp3Yeb3oN8qImM25ueJ3hANOts2WJEQl
IQ2tsRF+pDloFV/YaEwCXZFeb5IgUVi6U3O06rpzNYR7kt6D0Q4gwnWWLBpWo/yl
7mUdP6gCMYvkUcTmKrXwnh23ejkKI6ZKQfCRjgY3urNzkxm/yO066SsC/9ZS9ZBV
TNXvxuiFH1xLBNFsb/A2kOLIavsSz98MyHuQyiPIhNQ=
`protect END_PROTECTED
