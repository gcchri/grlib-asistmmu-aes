`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cxkwqJX46GTvtMmc8oUkS/WXLShgm35nIRCT2rnxdps9AAJKkJaao/Vk/um0MBHJ
H49Cwwg1vGC5TFzFgAOVw1lin/+zeVbu5qB6qzOZd/eSxsscc47QtGsVG0PHhFo/
M7WT6GFfwTWyaFy6bs0aNUgzjGKXErulp+GgZorRNixfabzpQBPaTebx2m2PizBm
RF0w/8kjK4K5vj3Xf7z7ZHb0lCpLYm0JMMuWTV/XIXC9hVQNRVgHSFnauLXrUYzN
cGik4mPi/bztvB4PeJuAEGaRmuCgX+kFZ5GM0rgNUljCb++fyhFdBTQjHLqwKKS8
GQYCRqjYs4oP8YRCyIkkrmpuFlHFblsLWj7CXJ9C+FveDcr70ps7DRLtzwnNOvAM
seI6g4RNQqT/TC1bXSNJbQWpFstBi42O1zELo712mCg=
`protect END_PROTECTED
