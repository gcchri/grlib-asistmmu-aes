`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUc3Ne3yop6Y33ivs8a1zWSZbyphQm5667OxfdJ4vmwgJ+ZHdvUPYu6p/OuF4Qu3
c56Bz8c3V7dC7uHs0uX6TfXMYbTpynbSzo62brZCIeY76zJgTgRdv/IJQGmDdPmV
Qgr9Tk7i+JzbI3SPyqP9VitDRkCnaI34hu2/Izkzq+zBU7gj8cfo/37eqotzmNgW
2CRbgdj/UUxHzQ3MhlORwusm0zx41WJcyj9TMousCoY7pLOMoqS1fq7eANekTwDG
KiwYDPaQYCTRkNj0fIFtPnQ5Dq8IyOJOrmObOHZi6TkrfApOwHfS4Sc2s2YMn8n0
Df8LaEuITmqeWa7nAp7zlGJCKGuMth/wHZgJ1BPscZuI9TDvfZRJI7gXA1dpPa6u
reRz9jGMbaCLkzuL+A082V5nv6nV8zj8ZyWii379VaI=
`protect END_PROTECTED
