`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzIqMf1g1r7J5ekPV2LFlXhykpWSUo2K3ICxyl6EmsZHZS2WqjFRsivRKm4n1/s9
7ld6dR30N56VMGPFKqIpELkiVO/Cl5Q5AYsSbujqbLe6q9n1d8MmvGJE5YZv+wqW
FgK9ENL124WNyFYgv7fukieSlYb/82grovZiAMnuAmXF//Xkus+amISip9StRoIq
kiGzkU1tMZ5vaMCMcbtArRlyRnii/v0u0ujewSKed/jpTma9eaqNZvkc7SfAHsx3
1iIjGHiEFgKUxdUo7GjrHgoz8UOdkrYKIRWQZeoHttpaN0hZWInjv40Bq4k2hNm6
xUXg5if+ZN6XDxR1d/O4Ijnpa9IA4Lit7dFT7zlfPaj13wXesYTmV8sKtoADNAhy
49Gy/mPaWdjE75HoMx2KD0YrFhOClTUgKmpGrJ/aPkdEM8w8O9govYnJD7z39WcV
mYSXsbMfOeFa375UWk5mV0xKAaZtoNMNSejOt7BZiritYsRQTxomo7t22RHZTvDv
kGExFBAwWTFDC3OQ79gE7z/BneUlvoCt1uBWGH6uI3CWOoXSItpbSWncoUAbSHmx
YpXQMQC0dBAzHTlUHqeJhyj460OToKEU31szvwd0ILwkhFfNJmpu+Mf6L/ef+wve
7wL0/io80ZKqFixGzsmYA8IzChXEN3y+RwVvSwF2dOC0oh4q1OOckdaUiyReYT0t
m3u+/s+PgM9tVuOz2s8ihHNJGQZwJN44Bc/GlukQOT9zDigySyg3dwsf+cYgk9pi
5lH2U0ZZ1hoZCJXclzc/xbM65Jz+utclnpedNchoA5Uo6AGrSpuYt1Zq9KO+PWSx
L1jiW7s10yic9gnxqdpso9vhX+sAR7W12Nlpry3f8NIuOSdA8QTKZkeIDqNQo2G+
uysSaJ9orEJRvJeC1Re8ukdeoEl0C5Buj7yIs4FHqSrDGToES33fYmvQ2vy+NBxD
XRmk6rTrPqJHJ/zG13Kf01K6vEIQa8yWD9qiUl1AThCVOCEGGHGf2aiSAVjl6hq6
lPFHmL6fCUY4r8rFFfAng+vzCO/Y4aJda3m4U/JLY6y1iiAzriw9UNXnPsSRNW0J
MYBF+YfzVvI8I5PYR+hfFJx0oa21WVft2ByrT0jgBHPdAoNwFp3sO4nPBZZDsN6X
ZOoUXMi0+8Ac5Ll2JiOwgBeESc1AC4sSA1wuK/zFCxozTOopkUuuezIXZPJrrEmm
fWrsv8shbErlhcvUnEY4/p+yD2/WA7Gua6abFwIyhLg5T5+LtrlhJjkkIRfKRR75
6++J8b5Q9qW51S12U2Ke/qCtEh5afabhzEzLDh0aUoUx39Ke1lirwQnRtYoypNDO
5zo6WKrYac0ex0AHa1sAl2IsEierkv/EFianCtZKekSjmxAbOBOMPCrgnDLHlBEK
+zAVVn3xkHf3ZZvkyFhBLg5xQEs2mgw0UCd0K68n4zYGJ0/K2j3gaZHVjkGADqzE
7QCuOa3gxAgUP+7+6xYmswuG4z+tXBLI3WlFmNvK5a7Tuiz9N0srLbRzbW9B8V2u
PzUS1zx9HJTX/1/dPVewcH0tRQTwlho15wb23WGorgtw2MclcIZAcwCvHhLn7bdU
uh3cXEOyV8914/fZ5sUOtEl4KswFldYKyB4TkBl42jHh1JA1wgDFM6fH9xG7LUpb
r7BMRsVWGLbjKJPHadYNJNQe4v360FGMmQoElg7VX8kSH4sRJ/WYO4BuSI7HpVpR
0QXnzfYqJB4rbWa30Po+DF+OSoKBJU4wQGtkJ8e4w+KnSFZFhmUNcHGzESYrQrLU
pb8N9quqvoZp3R532xfzKldna93Lbz+JgxrX0X3wKWPrNtx7mypNN5q+8oNNeb3m
lPoD/RLOte/CY70PJeuvBmtZ+w+TaQWQEDfREhScnwwzzhZ2dyQRa9moH1uFK+xs
q2xUA5KD3IUKus0VtdE1+5UvLUUVSPDzB9wewgmHnMXrD3T3tFLJ/FU5tmQkni//
OguVOkRTIEG6MEz0RsG1qto8v3xOFALqypeZrjicciekXfjz9nJei+++mqR5Jpr+
F4lwmzDXNDwqog/snmnwIShlqGZx0/LXsrqbrmtCEDUjOmvJiz9ojSsbw9pHrjPE
RQibSJzR71BVfA8jStKrAMRAubc+G+0lHv90pfnS3BffSORYocs2cZYwfg6c7JMo
ebNTfgC+mZkF9Fi9EiOjMED4gI+cLObLx/Lb7S2HnzpthQSqtYfm5bmL6PKf/fzi
GMWySI2W+LCfHC3uMKDUlbBqvcIZM2FMKoYQ87qr2Q1t789eCaiB9trWZ0yCcksi
saapQpCl7GqnCulJ2J74LssAB5XMd/B1g64lTmzfZMpWwXA7mbgXczARg1cj9Z5e
chxPTO3A//SOhoCNc6hPfDiFFMc7F4DzF6jQ5qFli/pnsh0p/OTw2OHDQ3Mv3YtP
rvcbrIjtNE24B/bhgHNbNRkDX79RXbsyFvxH0CsT+a9c30X1X9PCvI4uEOQBwcWF
5Cq5HE0LrXa23s+RfKcrYcAqWbAqSuk37Tbj//ZtIpHHariVPePNlP1xT+hynHFM
vaU6dztOKlthY7zwbHzlkpFnC8PhCBO4HNYCUYWUWQJPx4thsSiAEvXl9zeGUo5A
HnPgjW6ZW21STykUXWoRaY+MOTaooSVxVO/NkAlrDh0JdKKMpIMAK+ije3SEWB3s
IKmjOEJ5VTKtJlMVcDw4/KuNc/aDAcnVHfcjrw94dSItp47NkS4dTX+ZTROT1TFf
pgRy51k6gEpIUWmlrGih+i5EvcZlzmFkwGU2wQcCcFfYkKyG7tmrrHPHi8/u4rdw
Kotqv9TUei13f77LjkBIaWdA4mtJUnLy46uB4aMrzBhh0azUvr8wr7W+JGqhBzoN
NNihesFvvLiEFTazlTsFSA/mGHP5b2FNr8S6Fqlw8tERArqT8VmSv5OF6EOl9Y1B
yBb7uGkbleJHMmL/lCEPrmsPBhD63GndRdCUAuSLT6hPeXRnC1KOWpsswADcmLD3
rIbSkWVhsdSFobC8EmZJzkOIdz/WOLGJXIDi203sv5IXJN7PnOOixxW8Ii9AUexq
I2pk5jUGLHbf59j6DGEknhO4UdEJOzOV6dxd9GkBc04Apyac31I7JPFY/2YCFq/t
z81Oc6XF1nqmnpeQ/OfSi+2wDhlGN6imV9/rkGdw1/zfRWv8L5WWRpTwR6YLy3QT
kpoZU3YzpMJMn9AKBfxidLYpQSwjK/Xl9HTNVn+yXSQRp5BtNTRHEThBjupGcRwW
4EwRZB8bP6BEaWshvnsbwsbWZ1teRCrclZSLT3g5OZOClB9pK7zM4c+Q1h8zDO9T
HZU/U8bExMRG+wzhUxfAjtmJ1Fn8kwTyQYMNawBWxUoXP0CGSOVz7LKy+EIOiTXH
x3ejCeJfldktlsm1A+RCP4hUMX5VJn+JuoEt7Ol5iwY=
`protect END_PROTECTED
