`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ei2pxhh0E9Rep0XDEq7wCDGk74VmFWe72eHWy9CPI6KJnjOh8Dgiqg3gu2NMSLxp
C14NSLexctGs0QXriniYjwyqEG7BmSx0+Ev2RWdHMSs3hf9vLHBGQV04+mb6srA4
JGoIOakwuAUeYrgU0Ic2GsW4tILLzlKRvshFg9C7j2C4YGm3LsP4zoD6xNOxhYPL
WtzUnw6faBiMikunVOjucwUciV7EaOi1IA2owMskeu7eke9HBq+Ty+gwuzB0Ao9p
snnxD6DkH0/lUmCdv6iPzOwk+dJEdwhaHa08gCUV3dXPk/jE9oDxpSuKb6heod3+
CPxaM9U6fp0eBi9aHvg9K6NoorWoPdxnjp+3BMr12cHl+V/IzrS9g7MqKvM2x0Ac
0je2gWGJ0flZaDMdEN+z8cc9NUmaekIOMJYiiNWWdX9VLxwMEXaNuSAfhT1fZCBB
LQlpRLDrbzYD3yFAY5Rw5AghOTz3fCQThk2L7CufibHrpWHntIjOPQykSCrBrVI0
eGofeVkGHAtjsmhuzyIX+o1e94s9RE6B1f5m+Qr1tWB8oTrMJKNx5Q7bZ6dd57kJ
/EeEM2oZlP5/Uue2Ol2OCFzaOaMAwtQpFdeTRqb0Cxo=
`protect END_PROTECTED
