`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hbrq3QVmf0UPoMiBUgT5CJg/i+QncGzGI1M6e6pXitkVowngXoJUtzy9ZEEYx0Po
zPcF5ryAL4KvSeItb/BuArJ1nLEs9WDfW6fmmzSYr/yBh0jAsjZmehLJrtFd1sWs
HvEgyYicGWLfAq6nRbyjYdY1sbHmGnhCKWLTqtEORDsW7JUr977L6SbhCPvpW7aW
/2nEd8P+l6y47N84V5TfWxeAPQ9cy2D4mA3KEsoZbjlhr4oihi0PA/xe9rd8MYw5
1DZViOtJ6QU9gRFE/N6Agk0AsxC+cjaRHtPDEDBaYivWT4cif4DvV9e03rfvZNcT
ZArO5msi7Ra+cpVenTfMcZKxlf551jHnrXggX+DHJ2R4XJoq5/8g/wM+ryOXtQCG
wh+0HbAHye0IC4JZH8KglbQZ6fkdn1RhCeQ4m6SeklEA1WktROMJCAST9F+P4xQS
sN1JNgVknbgjmChFEnNBdKdr7tAVQb64JsM7UriMknd7o52WbwuavoJhTQFtidWa
nlIlg8bEzZwDB4MO+Ig1K9mIKEVb5o+Ak0TjMsNXhLhL+Ic1bRfKmJUJi41qMoQM
Ij2SnOnRfnpzsFQZP0VBErmfIsKvCBNJpVzjEL562yW7mDw5tOeq0dzJ3ew6egno
seiiFqWYSRixSzEzBHtlBz5hN+hX+J0OEyuUsDMvg4BtyvAd5c7413VWxHP/q5Sc
5AbWscMyhF4SqDhGbUK8YAduqybFuF5xuiMRR4oa+SlKZEWbexQY9wtzPUGtaXkg
ZL5Gh5uhewv1knFk6q/XxMbou+51jaO5EPYRxpJSxzol3r0lV/0rpq7VQtyWmIfY
VOEh6k0Vz8csiu9qgiGbPpxZltHJDLUuDxOqG+mQM1Ph8WCH0t81QnBcdbMWNbiQ
XrwUoRD8vXbsR1pt6CyPmVqQ3z1IjvhLIuNeTttYkgNXWGWd6+OWf0Onkc0IWV79
`protect END_PROTECTED
