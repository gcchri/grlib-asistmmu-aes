`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wshzigF3+DDJIiE7jRhnSDeOY7L/bUzA49LWgGs+318UFeGJ5zaYVjwunGtUZwPg
nYmXRTgs7pw9IQZrpC2mLyUuTwtHbYVfPKokXCrT1Qs/I7MLYv7Z7DnY87CrtEa4
rE+KSMV+C9eyFnW+fk1cuGn9oN02h1eKLMSJu8vGlF3dXn9dFvt5PEGbsQu0WE+S
WoA7daWxsGoC7W5TBng6v+4JbuoyUqmah2ESNQ7FCzIljQwQBg09FM6mJCe+t/zN
BoGi5gPBy6mfT/XACUCzcXfTcE78vcT/Cd4SBnXJ+/AuRWprDBxjCByWu3UbvwUO
`protect END_PROTECTED
