`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGmu6ZFngxEODryFLqiRAu9+nIQ1gnJcD1DEnvi0Xoa+Sue7N4ebDzKzwg9ZqK7n
BQUhm0Q1fChLVAm0xrMcygy2mYW+BUm2vG3Y3a9PTN6MSVhoCNU6B/ztnw/fvtZ6
/iQn8wU3dJa5/eGyAbVVIBMbIUN8ePdtioQZG1GAoNxYeGWpI+zyaVEXtmBx8l1I
G6U5L/6H4W1W48bdRUtL0X4IHWuFsiLA4itTecOWgOfI4IDCFEsaVYw+iMb27Yoo
cTZOp2JArCfsqorqHQZV3ADERFlrZDCkiqeF3NszpSlr202ALtIPOwW9O5ZOMG2N
p7/LheraS6IsmCeT+ncuKr8BYkHanDmocIOCu0MFkd7GFecRqSbi2X200Tj35Mfg
wLn8cg6Ylk4kO9RBkLL9EJbMPhLkzjKaldzSP35qBHHkBOj5fK/ND5pLIPRq1tJA
6YZBTYs8siSauuE0vY/bF9gMLmD+dvYkARuRq+oxFHnX79NUAUNbeCrtChq9kink
8E9IyiYVTFgVyz0B73KNKVPqOpsTR4fqIxUxPwgzEYVi0qjA/z3wTkUBQ008Qg89
gFvicZe7x/EVylCsmXFEwZO5HhWYXFeQmo3LS//fA+wLmLfS3kFFBGWCD3LQgLZq
UeXHHgdnrQcPLbIKaTbAr3EGCMMTHKK0NHluDDGOhJv91BDgANM8A/5i+sPUM78v
nNEFkw5UeXJg1wPMaAN9SFmH8mc9tnSvnAKFyvTi8yA=
`protect END_PROTECTED
