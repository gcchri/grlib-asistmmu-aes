`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zodUz/sZHsBNlkroGZd/iGmK3r5G7LXgrVAMHoakO9q/ioFuk01WV/lGXC13aDnT
tbQHC+v9eX7iYsmBT202ELf5+0pVLd5uYYV0yEzbopR3QMU+gngLkY3DzDA9CNev
vVdvWSDPchBeE5Y4WZNYViz/6VaTqvkVVREZXu5UcDi+evOt3/ma9P+DwKsz9J7L
HqO+uwG39YIjSVKv2i6I6aI9zaUegx2nYlXzeqStHV2jwGjkfFjkB3gy4haQMQEn
Tu4dDF06EwNtmzhJrYug42K8vGTV6IcWTpoX1FzHri54/NbacJS3iTbGf4Ct0SgI
ue6uwzicTarE3lFmeNnaZgy84RD53ZGFKpXt9NQOMIaCvwnC8cjjdb6x0L/qZ8IH
GWWrOJAiSGIDvNH06lc+Xhvop27Fl9Vu7eh4YpO2lPqbJ/aukmVD2nIrITIszlot
GF34vG2zIHVvFdvJ5rmmw1hgePUO8f8JYGNQontk49wUghj8Uw94Bkp9EGO2QqXN
OYJR9oLrF/TrV9wxW0J/Z/KpiDujisF+lY/oWwyhRMDo+6DLn6Ng6PfRuFB80W91
TBv+N45XYwGsP7U5zyLMSrmw2u7k5kvv30oOhkPUIglS/7rM/IUxjb+MZkckTGB3
/Sd8kM12teFXyfsomP1FE5FzwHeL0Tzir2/3wDZiqxvbpf3Xr94SCietkE/AApcj
TQPc3W24bOpgGhESDVx5telBMgOrUA9outsM+aQe2ly3+uQT/0/NTk5SACDrk6WO
cOu6dE1aAQTc3Ue+OLX43PfxG83eVvA6FfBuvB/hlUpnXHExHraykl+CLpFkiSDE
1luFH/6InBlKdbJRiI8Qb8kepmeSl+i/HdLMfOl0pWGfhNScGHKh8rEIYc0Wd15G
fDp8bVKYDBiDIJV4yYmIlimAIUO+BMyaeFJX/Ehxm2LtYK6FqXBp0LZFQ8fnqq0C
Zg1FN5vBCQ5cM+hi6BcvfuPS3+v6UGiJZMBE8/qtW5waN2yy8+8TRVtoqVqETSSP
IXRpsu/8H+dURM6cuX33M0iDc8ceKizn3+rKcfrKSSGdrbY8F8FazJ6taPpdRUtU
zJplqTYrU/RIzFJlNh6BOy/LZvW7NOzVnBqgW2jeI4RejGlolvO8vB2O4tTIGrTC
a5itXMqPwF1Ohnl1nwIZtVlcKzELwGWhwa2j9UTSZTI/GKhxw065OrclAUVkcpsQ
E/QVHRO0jfYLxPzwCkj4KQXfNymRYODQYv8TW0dCfk3frtEBnSgRsadRuqqNVWg9
Xtdn3PjI5OGxDqL+iaVh2ZyUBzh32KJAZzmPT50h15uOoM5/1HydNkfgHl3egATf
db1mzgkKRCXJ0RtJ6j8stYMt3up+gyO2S766KvJ4MJoGvM1WWi5wEoTngA6ADKZo
WQE+Q4zijaI5XOZhtVOVfoduryxM3gGC4WQjCiyBagXEQ4+FWilDX8xY/8Rx9VOD
QjZf86GLbgj2enRgV+/ZtsNKX039K3BFO2mUAl9lKQNnDI2fVME1RfEm95SM6q4C
7AV/UtuwbdqdPhb7aoibTSHQO7QAFeAo5klcaw089OQhj1gJw3VZ11JTd1jkFdql
oXdgOjuj4CimNGmeR5/YgrxF0ujJXNbB/9pX7x5mLrVuiCgXtdZViMd2pwEw+GkO
LVId1vlqs4ylq7GSup/Bzb+dUgI951DgESRW1RCp38+U8GjHf0co5J3zA5twXk6Y
sO/sq45m5OvTaWEXFLYHWfLzRPJqhmXwsvLSVMRISi7MMXcwXkgX8C+X9RaN9VKb
88UcjaUsdAUXvP4+1pBIl086a0ahplvKC8c6EKCtfLSxlVfaq6RkC9A6qrWE+sC6
JICsaOkP8h/ow1Nx0g1oEhAuC3EQO3Z5g9ilVO0lMevljtnL8fVn4oXfVanDI9VU
xrbAL6VzsIGa45hKCacy9krtA9dWG259macAL9LICGXLStf1Oszx44xfl5OgChjx
yET9C6CN3UxT/IPvOZJvqxXYbr/0jjq8Eg5/O+q0yrHnaOA9fjsnXiuA9BMT816H
Tr9p+9N3qykh3yoP/pLUakP/q4lSMUR1Tbn0Qud/2GYju9DNvSTQtVbqrByGLtXq
llY8b6dQudn1Y2dX6mHCcWsEURRwPOHqnZtuyT2Lbb5IMj2qxO8BxKNz784r4RWa
XIBtjwZ0hl6bpcWdw7B0dLwDWPaRWLLgGCZW9pTv8+S0OSkayG4868qXv1iNVmxi
cCSoChIbVsqFg2+psSdKT9ipHzrA3TxoEv0IT3kNPkl9zK2rrc2a7dcAnzVj791f
kDKFLR7+Yxe3fAKM/kBuqDkktyl4Ae9JrJuVjBYLLvCmf+Us8NmDus/34Wtt+TQt
8sj5837+30E/mySmNowr3lTAjwK6HgLkWNbguzd/7lipMpkHvfdFpdzKaZaFcfgE
sEdLgLJL//eqeGUr9jrxiLPtpohoVmfrdoOmnEBo3BUEMygta5SFdoCM09cX1bR7
oSHhEZJkkaDi0UE0WmKFSSdltBIrv7/fzeipNRgoAJi24CmOyXcCJi1zbXmyn+Hj
6YW5yCRWuN4LDAVwLFOXkFXorQ5IICP/X2LAbFiPzJoO9z9JGaaaxDixV1pvAa4g
JNtXKTJHIDlhHN6Drj6wf+TSPrygWvU0x67Uklf5s/4ykHWV9rcuFeDcjzLyuILg
q453HO5g5aRHQ1PtOn6Ozaj5aZYLGiRzy8IzV8OOOtGpUOIFaaxC43xBATLStJb8
/t7JmyvwLr5LplQtAZ8Pm6o3rmUQIrt0p96ifctqrma9AqcxCqZSxnfS+aWycmav
BYMQ6nI2TtNRM6c6CpajJ7Y7YZJFruYX83+5dIjNNgPxHcD6aBCRZXnzTZJ8Y0XH
omboLtHu72fYH5cnibubNRNaIczVkMVxOsQjfffAMO2ZAnbqQD9PjdxYBxgIzL3D
wyWQH0gPPlyKCJfDj5ddvjIiu4R3VLNIID0AKNjVWfAiLTjAwjixy7nhcJIFeYPJ
AKb/OE4AIPZRpba8Lmk5iXbpzJICWkUn5Ae3nRKgZsTLbwsgyLtZGl+OVfR2ZD/i
mW+5mgEm9yPMtyLPB849h6e9/XkTLHTEmaxpvPxypLYdMG7RFxKXpa4lkC55Bqcw
HJA/DKibJFepAAY9Gy76J7YzwZjPuB2UPo3kT9epeTYLhTplSP/kFjacg3h5Ttg6
qOdIaeflrDr27Whc/tbwKUGKn5omKySYZmpWoabWaq24RX9Q2g0PC0eKJcPwHmFp
eA2tx/aRw/boQHW+KUvXDQuA5xi07KSRLMOAlRTmcB0l2Ad1B8ZDb7vrS5u916mr
MYFGdvlTdFBZq6fBBZQUaFeAkcFXCIKxdBM2qAW71JUWiBEqfk+feGljbhui50DY
r9pzhmF4CLaIxN9/NDAJ2qccahcau3KEv+lMr5avrkhTLE3h6OYCZcsTDyzUuoqh
8JDEwhEr8ToEoY3f5fLdNu8gOhnSAGk5nNv7A6Z1z72rby3lk812N7mKVp5Aa+Lr
+mZsP0fzKOauAKBPsqoXHdM/3TNm9WQ3jmiHHLDcIH0JxRYpEuX8PG4zAekxRSlq
KLvjIfqNJ42LsrhmwQd3hGB+xJvn/4hhutLr5f0DbAr1TCSi3/Ym2jElv9nqz2GF
S4OTd3jtbdBSZGaJtDRp8BA9KYyweoyBZf+0Iop7Ez/L2i5tA+Msu3J++Gf6TMNZ
f3OMrH3S/87cjdJHslUmpVU9Yb6dJlaDGnxmtDF13DorAgl+ckQ/ZUvYMfklq46A
6COI4jP6FkBMOCw5klhg+ehVQD5v8o+EHCHufxX8dmZO8lt0ZM1Y/PjfTabGde1F
P+BUPtgouXlvmr3y2o2Ti3MR1YRhEVVIguBdGKQk9QeRgSIItuViNboo7fez7Ddf
qqWBN5VUqQvkWhKNIclNNL0QJJxeN38OkeKEtl2fHtTcEc6Zh7C4Bb1n6XHBeL26
JgnSPUmvLB19X9qes3EMlacneg8E6Nq/POdtC7G3tpcC9ZTqUSvzwvSsIvX+l9RG
28y0KwH458utypI1WoQks5L8qxJxUzlhvP2DucNmGrXf/H043KvQ1xtsUKApWPf7
FrHA7NrXNALKgj1JqjAMtDnDzldBYyKaXN5dLCEyCVZ+ufe0h6/qB4DF/HHb1GXj
5q4uHIZt0uxsbqonG7AQbEKsZiWr1+hjWfEyQt6DOFeyhZQ8rUtQFztmnb2M8KC8
zXffg7xtfSsXubkVMbts9eqiLcHKmv87Q0CxeHonwpPhXH1kaLyiR2U8VVhktTuL
3xf0IXy1ZPGRVgjUCB4P1I6875ZvUsPCg2o9C5p2u0GTnIhyFK7JGQJ74BGB87EG
r4E4YVtQxp8pe2E/364EHyrXvJYkDb42CDZEr7yWt8U=
`protect END_PROTECTED
