`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yv+eD4hrI2S68jQ9yP2zuC9drGuhrE8V5rp17dshwtZriqO+3UZHm8a84cDC8IYe
O4CBdnSUzLeF2GFu9nqGo/F3KIY01LyXFvt3ZH0PhSwtwIAziV4tg6nrQFE3O2xQ
WagKpHxhlLBfjXQe9i5aNyjE0NnqudeI7codFOOcwnYS55Dseei0LdiUQwRzPVot
zZIyCj3zvgADxxvQY1sPf0bNgmIUbcsbt+kYu6SIq3SMsZqVHa62Zua4pvyciTlU
noeU+bgNl1hmtE9GYa3BnqbK8HK6dxCZYCX06AkLCSgxBZhgSpLN7Tmq3dzLFDvp
r51ZTQMVwg6EaBkJLvC7uOgJOdnBv6/nlYK+UnOloCBBXjdeUrW/LzWwnK5++IWZ
psm8oya1LZZjj4IXSP9juTH7YHy/4G176oOVdTvyKuRj70RRpgtNbENs12wuPPNQ
C+mW4X5Gxg6lG/5xgxMmE5Q4ZYeu4BXYC2hGSroPZCBRdBl2ObXKRx0TqesHKHf/
qivyit3sOKj4rpQgX6tYP6Z4xU5Lv9Q+U6+cWtrwHPaY5ZW5PbPCrvp8AgEvu/bO
mAtkp+SGUSymFb77DyLMY0jqAx3FnvQgTdVkH0sUlPE0Rab7yuf46eexJYxlCwdS
BxxFX//1pi2Q4T5yILq7BcuVcev8QMCvvpe7d6B+DMMrortsSEPl8rSphvAyjCxC
9er0FLGjRuUU/sqIFYy0FJ3T4dFfa87AoM3mXvzrreKPSunnxyf/ovoa975/h08I
zJzbaOfcJ903Z6jlUIWsIzgWGrwrJONV+8pzCNiAJUNSQBtVIsDTenOdv4Tlc+3F
p/XsNv9MXOWBPZ/iFCMk1vmYyxKnYnaUsSZABvBDT4zIeTaPBRCg9/u8mp5z63KU
eqZGbsz0A1eVqo4WLRinbsIpc8Qx2bwGd0OmYxPZkIvD7IMdmSA2iDQsDbEL/Y5o
5iZ9rsnTXq6hEgQXn3KLkmwYOjxqDKf0z3+izPoMqNeZUAQw8pski9zKHDeo99wW
qIqp6fKNZ54dKsB4qC/feBu5TU6+kkJv5EjUqfXTLmurMldvuwNB/jGIK5kJeK/t
Sdig+vdKKAosY0Q8OV8awT9rDRYUh4m6SSgFMKKcFManJQemKcwfdv+fU2ZtvmVf
d+rlQXkNsNkU1agnY6xsSiFOhkJ5xukYyKghRm+Zu2BgbUa2mbD69R1CY5MeObBy
a5tMVlyHMWBYr2gRscgxvkq1zZV9RD4rLOS5PUcF59c7938t37L+eNBCpcUCZE02
SXxX2lqDhznA8TU0njA7bDynizAtOnE2Y4HdFK3Kzs0nR8/M2EgVDUutJzknQ0iO
KEp81eUTDvcec8+M9ImcRN65h2pOLeCeNJ/KLTMHjTCGXQ62jz8mF/xMCqQkbk68
i+21Em107lQ9ajGTesAOnHm0XuUfFYwVYC84G9uT7BZrK1jreXe5a142/N0OiIPm
OZY0WckkuVpMur33tkZWr77rcZ09pObhiegwc7iN9ZZB8dcfwwNkSMWfvdnxblZe
ecqHRAd3g+pNkP+EfEWpBapekdlLTJfY8G2fnaT3Qy+VcTjiGORDGkOeL+QcvO89
3IeAoG4I96zI0FmL3MlXAI4t4KqeT3+YCkCeRCU0XABwA9oLLdB35LeD/54bVVk/
9jgc+UC3TzxjDNXqyP8qcr4PwLGqa/rHyLfKaqtU6fDRkc1kdCzAm21qovXobwrp
gr110x+qoG8kcgmhGpGbc9cKlVKfGwpBROL7I/obyjk+yUHSR0Dl/9GDq5B5j4r3
IGTfFAc2vK4sh29o/BwTYxIEnpAiIcOi2ier8ztlxGSwxah0d0l5y6ocg8RBU1vW
s28sEzRx6j9yucwv+E5Bsn08CIXf8QEdnE4UdWMe7p548/iB6tKifNjnl2gXym/H
I9ql2xcCKmDLUBW+2WsRdK+9c30QXvW8MEyrWWKqrSzq462CJsJgeJItwyfe7++/
mFCzVhk20u0ykP9lq8bMSB6wER4n7RRjcoY/tFjrJ5KvAE/ODh7MSCH6XsL6Qex7
eWzut9OB+I08UGkU8BC8ospxregB9VchuNOwg80dM0bsGeyNHY4ZzVtA89UGvY3g
L6w/xf/VRh2/pM4yLNN9BkmIy4s/EG0A12OeOoKhOLlv2NCxVQSnnLpxHXt7mnaV
rVgGHb+RRL9nlkoSq/Zn4QA+E68x8fLYRnFSMLgILmH/Re45IrssKvCtgXMt/2kw
/lCS53YHblJZvPmv21XgmD94fslWbAkdupwoSiGybNzmU/0q3dMw77V93JzRR4Sm
3NpGO4DEfc5/z8NefhpEWKT2XP+B4R6LH/gu4RgMi21ajoqsUYX5ooP/v95/4OqA
K9SZKWxvqogn544cDOPw+PuE/sz1fMXsx8CAJHz68kaHTBZmP39moV2EV6r7G3tP
33UpgaCZhi3kie6nxwe2XdfRz8HizxgZKVsXooIT6ucstZ10sf0Ab8lp56KX7vZt
3VVXHqqyAwljkzA7QgQOMCcSUMytCsVcR5IvMYGTtnNGnJut0rRq+1MlA2oDJ7s2
U6hCNKgJ82vBmuYR0vROy2tf6VrZZ1s4PkOqzVroUJXMiQ8KwStw5LyenYeb79NW
uzBG68r24w3BuIzFfPGoJrIcauE934ONG3qpRVINQvM1OaJv/puLI/gbThHCVT+0
mFPq3WZ0x/c5cw+h0FG8Mvf+Cau8B2tHdRL+hG9SgLlbgzhyAOGnfcwdui/sWDCj
9rh6zsbGFN1eDnHP+Ljt+gykxTPjFAbcSW5YtpP4RsAX5dPgiMRTTZ4TfKVQD6Cf
rtD+v0iPh5K81DjoqWua1OyxdLaccrG2E/fDXs03OjixSZuto++JR6xxobT7yX1r
RDE1x921LIV9ajbpqJVPT/poWUFCMfh63gMqO4fuW2EpimtvGtgaA4zL1IIBZ7+w
03TErE6zsR5/pcDgtbpBJ4KwZBmWTY0fk1qMIy85eGIi9jP61R0CZiH/Ad/kdoyd
qoVsioTnFyz5j7I1YFkGMzTsWRDOw0us83d4qM/9PuiTOwnAq/JcRZbndmpDYBtb
pEC3NFdLvajgMBcIZUhGJHbyR0tKM4OtlbRnhyTjNMqYoG9IbNEAF/0LBK7KdKCu
WREL2wbEhboo3Uiew+Tdq5Al//LHcRCAYFSNFfhg66YPzi5LflLUOwY8ZPhD2yek
h0NWElxlfIawyQpIby+KgWOMvZ8VQmhOwkdmwRmJ7NEelHayxchx6Mu2/8DLphxt
KbkB5b5K0BzjXxiQsGe0iaMiDJrgri1duyjkk7I4yHvkb7THnkaSMSIjHcAlIH2Q
70cSsbuVptxRV+kD1QIJAKcoTKpkDk9etg9MBdI0IbbA1ZCNqePYZWg0Bl2zOwPD
qDWi1RqMhIHhZ7t6jv7L06qy+vzoS00UHdPsNxVqn3OCzufDUGNe3+dv3XCvL1tk
F7YAUD4PdShxxlF/LFmc6Y8iezLBtrlZNj+4EIlP92RkK9FziNyJs7jmPIt5TTze
RfX1koaVwGKMh1jGadfIRaTzk6hAXB6H3fICNFMLs3RZhc43NtxYAhhFVv3bAAkX
ZTHcIHBH6w29V2HxH/Mi12NWniXXkSklSFKBDtGyjEb4jElQvie+MS8Df9/yAYwL
pqnp3Sd07AZsl4Cp22gpZu6GTxOeG+HxiuzqpnhbFduA0nian4I5Zomsi4v+0SbE
P1YDxaAbr3BHqRG1faeFdvczT2HiypnBKTY/MTC4Uu6XP+jhPGvrXHgmD5U0OR5h
hFZUM/GdCLKfCKNhkb/bL5r6ldniKNJt6xV0BLQ2xY+jMr3lL3jrhJ16LSbLr+0w
DD6to3XsH6L3hMrKJmcCn6Eg45PMfLjsfy+9Whie5ekp5G2f9V3rq2a9GuESzmFD
MSCyd6uTemzQmHkeR9vL+Q8g/jtf/EWuc9eTVx2t++GPS2vBlGXKIF/AhYj9xEB0
kUNQkzQwIXcRIJvOPDvOMIhFGROgOdV/F4IAq+r3jmSgbBOl93STi5zAhzazV6jP
FrGJdYNUU9v4h1tYt+qh6u/c2cFpadtBbITUNr3O6Ze/j921tHdvLb5Pbg3UcCKb
XpJdN8CPOKj5UunTeCVhI/0eGHOQBAaahVjI6n6dePwHJNTR7DeRPk4Abwfx3KVc
lTpa32CY3CiRTX0vXduRXU5ds0jBWK9qzgdQyRTejCQDx2kXqm9tcGHFcvEByhOm
UOrw2x/b9KyQ8H737XHmSP/YrpkCtXotM6O6OWhPX1Iq1hAUCVJcF8I5pWfnT1M8
lf/AZbbevuzcZMilm4iLt+OGHGqMptuQG94eARUZ2CcgeucQcyRFijLijlkDORxs
ymye6vzcWyAEbO4dRBN84zqhmKYjKLA21U05X2jO3sNFpL5m7d8pwIlInyFt2U+8
HrGlvZFUXW5G0fw/fnERqcwoPmvuWqSexdkrYwoTBVbDzCfT/XEfWHgle2FZ3azN
ZJTmYWx52+uFK+9Gk5bf2A==
`protect END_PROTECTED
