`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cWaYSn6aqNxEAD771kVCWRgx0MpI/ErX7nY9XyVzeUsUD3mxce2ZkrT/fQWTEm7Q
G9pEg5XAW2RmVLqCYWLfFwDz0KlpzOd0utK3W/Zf30CPFXCPwLRYrr3n6uT4VvOC
ZD7qfwaSJZo6kQ7RuwvoCdwm9b2FCcRzQ8Y6zUDNndf8MY4VBTVgl7RU6s3tOop/
CSNwjGg+l7p9UxRaRtn/5wpdVgJZwGvcCKnmv1XjS5JUUMHPXwS9lPfAPi89FMIt
DFWNCwUZPJsz7Fswjls5jrEdrZFsXN5NfusNhci/48WZ9930zqx3R2aQUwNdVed+
3dnHHXdnO0uxUMz2xhqw7tMqDhdoELChVqZH6atljchjLlgsSadLJVp9SqNDh+ry
WJB8FH9zHR18uBFbBuV5iduCNT5ORL261bMc1udgOBVeoinqrR48uMikDG84VeXO
`protect END_PROTECTED
