`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HKNYE2N20RBTtmBtuG03MGlsCThZ9Pyr/07DK1eRaaHWYzXmqLkKgHhoez9NhRLY
dRhpHujc3iVXYYSBk704fEKsyvA1rn2Qfamh1OXr4mayjCqBag6jouPOIfwbMCXt
k9qcfuRQOTXLLrVWQknN6zFhhXalVJ/r6AoPNA5WzV9KLSFW4gdHNJdJazJwydMQ
8OspSkQzyINcnNMVF8z+sghy/x+UzGfu8Xr1fmvm/ToQhopAuHam+OSobn7h1br8
JNIkdoqXqVtjpxy8GC8vfnE1CGAHuXxxM9fAl3Kwq5h5dKvLzo49rZMnldMoqBlm
XxvZnVyHlUla5UAcEjvDcNaBefTq7jMgW1sY1BYVPMVGf59jvlIwBKr/iexMBrbp
Nahp+OGOOH7wBZX+dMVQQ6x4/yVK/4zsvXZtaD6Pvbs=
`protect END_PROTECTED
