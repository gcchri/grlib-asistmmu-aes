`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/l1fPJ2upc15LcFl+AQ119i0kMKnG9nCSSgUjp7Y+HXGUlo9xij+FcQf+iQuFCUB
snCl4v5Uu5fyYDitpLfDCSRnv0EalDB6vXlb65Gy33oOVc47iUofhgR1SyQlE5fp
ugZX+lPqgyzNvSpcIb/tU5/tOFKMwebTkOZryTbCk8EX31j6Pg6HV6zx6n9DLCIf
oTAbDNnrRhurB70pt5WBL8TYMK9+a/R2BBsEzIyXHbb/rRXQQUDz5Hx/TPMoJggI
oKstoTO9PlHy/RAtnziBRmFcG7mQJDH8TNDY5gxrpFKyLxRJp9cB/1ggQwb7dYSJ
bZ2QQzUQ4PQ1aSpxbRaEs+8oG0/j2s69zfV1IEf/sez9xsxs6smCDcUlfcHCnSQc
0M5hXScSDS7uHgL50qxRk4JiGSi4y/d9+yDfUDKpXHl5s9OEtCRHuPXBu/JHVp3N
`protect END_PROTECTED
