`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L/DLfLZq7h7khrQL30s+e6xxWBVxA5vMP0HuMMGusnCQC9AwaCcRvn7cyVwnBGZi
2g6058MTCFKobmsZ4ZN24FkhYYfBL+MSN751BkAbd7lOonE19ki3PYVfaxoDSCoB
lsq1SJfDo1xeGDCk3LbfAQHLkoF3cFCIY3ahynxt9NzCEN0JIlYRC1lJ4CWXEEAu
Fdb7dAQMSt/qDRyBsH+qOzxeEej+v/joXeYXwqizP5zCglUgLpKF99X7Wha+YQAz
hdcfq99jOes9mgPDx5+HdHQT9OuggBJ7U1O/RfWcxIJHHkM+MfWRqzozI2IoBery
09V8+dXCuVbn0Kj47Fn7qVyZAyZQAvBGirNlJHPpoL7l46zVl23HIjUV/Kcj6+uy
IfQRSQ0w6EzCn6NQWaIBQTxl2uUOB6TWqe0xfHnrwF6Lu2iT/TSoFlelOAy0J0MQ
OTD1PearP+gaMOGOxUkAJP3GiyXFatbRr4MEOVsa1aVAWUVUbwBWTB4BJb2sAwhj
DFUmPUP43o8qcq4F+KUxjiyoSjafKRYpAuNhTdmsgQ6+vdPb19xHqErOSKplYZAb
ZbibJNc2+1QeqZzRmJf75WEjf9IIkRFjxkBeLpGTvt8fTPRGXRGePh7fUZ9NRPLk
Ww0iYY2TepnSQ0JE1e0AZqF9rMhnVHbJj5qmEFuf2rpt06xt3RSTof51MXVE8mEn
zCN17Jdkh3o1S6hyrrFLDlLqFvmCfS2wecc/uaC1ibKRcAZ+vzvuFZvu2eeSRwFl
MHz6Q/ckivlNPWO42PyUOj2uaKpKDku700XLji4oFrMO+uLbW2IzG9Y0Z1TeA4Ms
x4CqK1kBqQ/i2vttMrjdT87Mgc/2D3nclTqljuwoVibsQNAdzxifKvjGJKtAHP5a
5KFc+DWTCXmClJ0VIK8NcfVwwatCk5eb1Wp8LbdJ4NLYbYZAZ4FHJwZhjAa3AJbX
RLOH3nQLpaai9yXJS3RYfxj1ouZoIoBbsFV29YcKlAp7Bqzkzw+C7wTrXZHtAMT3
3VKxSrwwv5Af3vMRNPcmol2iCa4K89hQ62CbZ6AQmqDKti/7YjdozJJMmorz7vHx
mdCxQrbJL5WimRdoozAqMoPAL/Wc2PHdTuq8sRxgb84=
`protect END_PROTECTED
