`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GL5HC+iQSgiXL3uoKmANNzjPxWALm5NKoVJ3PKEqB7Oq47ymNZ1uJ1tGoVdwKYP1
l9y+AzYQNtct29phq+qZ2yDwTtRhXNlPrrERP/DdWnLU61UFIoPKCuR+1R+8k3du
JdSt0RZqfyIfgikkl/H2bf5WHt/WT/l5GNLe3I9+j63gIvAHIaVE2Wea1bBwaLjP
C8ZcKLNA8X59CIuG1hgaS6NkdRAAPBflc+9yJIpuGq90LA5jm3Nq/ofC2f5Oh/9N
iYDkJHLm2Affh/VsAPeDdhezhn29grkXwldALyxZX/e5LmC+/YoiEQwAf3QQxrTP
8ZDQK+R9sHH2A1MrvaJBS/6WJhsUcmEGCQkUulK5dhhaHW7dWYrktaioaond5iJv
kAgw86RQS/o+lCsI9wYR0YfpjFJduV2tiP6HlbAvDtX064hhQv+bU3gygXghhMzq
+75yFNg9RG+z4J0XM9RLjNBaf9gXsLM3GSVTKZOQbJXMm8edtVG9wPmWwvnqggWz
lFkuyzRgeKXO6kTChMRkzE2tIA/Jom52v1LLxqvlGgwffVZ+EZ25VQlIDf/8+Vpj
4wIXd9KppZlF/22e+1yVSFAlW2lE+o2aQ7arE06nfLQG9mCGdfKnmNH7Rx2SMltr
+61zGsv5v6w+b4zuo/gDDuVgWaZZcVr1V45DjuhcuVM0WptRQfNiNwBkrusLWqSF
yR4hX5UrgOvHanEvTZyS2gDBPubMguMBlnQBnUlCweYJzygWuPwKSFWkh8fMIwKJ
eZh3SLxNka/6+8FEAS6Wxw==
`protect END_PROTECTED
