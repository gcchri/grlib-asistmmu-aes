`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wk1vvq67Bo/bP76WKf9iisnLOECz2DxyBfAAPU7OmziqSo/ZI7vRIhDoSGC6aW8q
QsC88uBSfhJNrjYIJDSrs5+MK6Oh7ODjqQcocClnGmA1r7GMz00vVX4iHBXye2uY
8/ece01i2G0YvUBRk/4m6bYEhmVXcowNWo225q+HQUFz5HegOHu5K5adPs3NDtAN
ka5g6VITXqLSdxd/q1PP+LRcRgXgccupg94IPPzA4IX1v9TCFpdbAz/YRTuME5I/
nV8YZe/WtcnmFqymSEawLw==
`protect END_PROTECTED
