`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a69WySdrVCWzvDo7IQxouhMBICNsuBKhSztaOO96Yka3kYczTygEDn4KOHaHOJ5Z
tEAwBtB+j8eAG245XqDBK7p6Sc0snTzD37ekSkoShR5PEvTQRMuORVG1RGV6hrlJ
VDeqZrjuptY9DpBYWBpMmAc6S1AxGvXFPzxWjfaH1Fcr+xZ5Ulabn7xqr3vbD42h
EORlPxibGGzlX11gaeZnakyTxEenSgcy2YrbbjR3JFDCafTN14x2syU67aRjw1fH
4ggsuam5vdPMJHoaDwSWGmzqUS0Gzi+BHXGbSCI3r9QjhmOYwYXCjRGWK5rU8QXI
7ADk+NtzE0AHq2k4xEi4rU+h+AqlSX85o4sEpr6A91GXeSr6SoReJDi7l+yOi/ly
/S8V+acZ9Oht/g86a/pmLtRlzsDbfXzoWXV0DNWVnYEiknp09jU0OEqXHG/ExTB3
HsyzoMEzo3BZCsF72P7N13ycuN6f4YT0gGXJUpBpQ1MauOHO8tdsUyUe5z0x9f/y
`protect END_PROTECTED
