`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JBzPlnViM9B6IVqG7g0HIXdNqYHowwUQYvCx97+zAEQQX3d0HcPfhOHV0Wno/RFt
BVYjywtEetO/dgx3fsiO9++CofwnJv2Ah7gw8FSSQuZxXv0It0fLXaQStDAwZtFq
41nyRFotWhuz8KgrVMBWkgjPIQYlpEWDyotOrXoW3cjw0MHPqzrLvf6mBKqHu4Nh
wnaYOFQlBEEw/8Z0WgjkAX8LHlN2hXgZNoqX+kxgN464Og9PWtbxi89piymnqWHS
Tna3sHqHnnTytO4Rd3RljV9PlNg+dvZ4Vsx9weO5FVoSbQA0OY/qgB7M1+FCB6fu
GodpXiK/qTX/uGcwBjVwHE+zMHXG2gqLs1JQ8r1Wtof9raqZAF8Zqq4vuk1GN2EA
9l/KF6SCPnmfz++/nL/BG85/KchasEdpMnQ97FQsAIrnFdSNC48SQWZzpSWIZ2Bz
s20Coy1xdU5Ei1dQ7i7v9+zBLrgLlar6GQ7DU4Z6GPthZMA/AQVIjGFGHUEQg931
`protect END_PROTECTED
