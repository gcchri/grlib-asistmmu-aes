`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
isNEJRZVltFvykbdqa6r0paM79qWUz+jgv5x4kam3OD4KlEfVPr0Idyx1vA/0DPL
msiI7X7nQBh+CtAP/cGDaVCREZjKJxj49ktxn9qCBKSczUy5k3Dvidn7gZgTPx8p
hZEmoTRPVWWNL1zms1C8lKOm9ax/vnGHVAOjkSzcaPCc8rzqkAxSvY+HbkVDzg63
0qWn5S21R0c7c1Fon+c70TBmnh7c9MHP4f6OaIp4unQXSr7y8CE+RoIbYJ9NWcgy
mrBTS0ImMHGUKsc9EGVEhabldwI/WK2S7s96RtaF5NO3JPvCMFQ5hO5x799rig3p
wybcOxZCrG4m7jzXLNfu37mWZ/knALJSt4uCqFXmZC7AXlglSVpasc4w3fqZnXTd
Op7xmjGCh3tgVfPHLW6N7s09Fgg13pu4qb6WmoqBRIGVxWq5UFfMcAQn1aVdfr7l
UFHovEs3uhz5kL/0ouD2nwKHc9cp0OS9kIz57ggtgpmDhmBdPCdusheUVs3pbMRv
0jYdUdk/muQQweZy4zodqhLUbemB9TFsBEu5czryuay955H2boB6jGKSQpRscF/1
K6cH9eZFVLupRMKEdVOyKG95ApC0oIoDBcKX3LMVpiJPCARr0HCuuR9Hcx9yCiQR
yQQyi4828sVxKQPtkhwDaf6pQSEannJDhZ7TCvUsIWO4cLha5u8EAk3R3cMDVwg6
SJSMdeeP7bvVL5iI2iPV0dGOUbMaXw/VO/oAePOnZd+tEIrJ6111y18cNQxEMyEW
fa2VzT8qNpcNLPbGojUbu9++3gXuDgm8gs3DziOa8KcRjokdmd8T3ug6PJwFl3xL
P2Qea6fSj1a+9hsbv53NBF7lEOGEV2UX9FYhspsMDnWYQDSzOACMBjGjEiOLLxiB
tV+W5e1gfTZDksskFjzZI4S+39of9+HzbzQCsP+s1FMiOrhS0RE2eB2vDCAr8h4y
r2KuVfy99iPXKPn7xxPRqSVnMF0J6jB40+tuIWZfmU5Nm7gDPYMMhd2RI+tYFCIG
NtF/L0jT6/ShzOxX9TOF0uzQ+9QFfEg8T/s6DnbCVcg=
`protect END_PROTECTED
