`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U30+37O8Nq9aUvWOTR3fao8JVEVRzs1WBe/IZMcm3Mk5GtQDVOBnvElTFWN8ITpu
+gPnm1ZEVbzxt2rbR0mR7FMPI7lU5xDvoP16qtxUy7mGdn4RpyFuLLYd+7TI8p9h
lA1BMxXzxmLmOTn/hvfONUUj8i8eZQabYj21LZXmbqti5vEJjfRrzu071QcOE5yV
dAia83f43iEtQMqk1V/tYz8auGjGvkU1rBSoQZv2qB8MCeGh+qUWOogR66aagSAl
xSiBkqGP80VWStO1RHm1z59CXpUcBhyyQcPWHfJOhSF+rw7RoEXmh6CzcnrNOX5h
O4YAG5wS3PXV10uGnMlEtBp7MpHRp3goGIKSTMUMfldqhbC0EglYLAeFrnDAvj1b
xYUrz4COyzCT+5IQIc99mSsW07sPokDPtUv/+nLvmE++jCG68OF/gfne74PWl5Fj
lahm12JJXGos1xmKXw6MSz56dgUNMVmUep59gW/CPyvfVRJfCx8p7v3u2BjysqDH
h/1VtDATc5KWkUnzY8KBDMvM9wGvXqs/8D6A2ZFjNW6nWa8k0HICbN3l0kVF3Mdu
6DIw7AlC1WDxnuPqfEfEGB5ad3arWdgMRF9tJjQxxJmUxTIDKjGZn3d+Qk6691GP
0bj7q/toATioXd36B+Wo8P6tXp+FzOS5rn7P1zbA1nzp1HpAD322idh/rqYxrWBO
qYwD+pTyUH4UFpxaZIDtHlCQaFqszEdIZewbVaDVW4TfFJ56CYZ5TZEZpf6iK9/f
6zsxWL1CAzVLzx1Wj+Nelw==
`protect END_PROTECTED
