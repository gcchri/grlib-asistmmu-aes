`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILpoDG11oMfvPgc50s1/HDRYkn5W7/7S105tv68MTRM3tzVFB6hVhBNEC5dWBleU
fShiEmzhHmYd46c/YUtTPM44RxulMf8aCYpkt+Zwvc4R57Pe8jvEYYl6+i99+WSM
AacVbIw+kAHqwu4EYIk77hLe74lTZb5P7GW5OlvAIkdfYOhUf788QwHAuVvU4xmY
r622M72NjMtJu6sVXGub6QbKMLmsM48zcxNHwvYndCBz1leQH7KqDof+eaw3SjRz
Gayo+gL2ALsjyFur10yH1YW4FQeIs5B5mOXQcu641eJ9ZT2VNOaTzT2InVIY46PU
G27CPM1WBRtTft+w8Oi8QIO3rQw76XDH4WV/evKxipkNrqUbVxLIf8ZNUsWVWisa
/IRRhJWKdmGUS0R7tgwY+ERQLXtqQMj5iCS46n8Vt31NV/FfUzhdyW07OzYz6onP
j20Smst+DvYfyX2OMCdwuN+EeOoMeCuPwL2Ozk1nvoeo5cGrWC2dINWT9wTj7eDE
3AEY5i+jHmHjAb9E8HZAaQamPCk6JIN/dmd4Jlf8/ZI3eb47YfoYaKd7daQXzqnH
jZx2buv8XYZ97V7FbKDQ+m30FprDqO3XtLd033q7c+37CxoVHCoYvX5IM3UsGbLU
hmzsoRjWZJIruLAqji2w6d1pn0KLXgAvKCQSbTVoc468MsdX9a0O3lymTAbU1oKm
/m30zGHuWSkr6JSva29ao7qi8bz0GTVKy57C8Mu4hkYFOvKmh4Gk28dcWifSXcng
B7JuciAUvQrKTjsv3aufl1mVipB2TxLISd5nDjdmlYug+5Y+rs+OFgeDEpWhuMRs
+DNRBzMMORcWITQ7CglmGwXdQB5E1OWfEPbCrHuFtnF8TKPYghtcRcDwcaMw7Yct
G6v65auNquCf3iEI7aQFKbt0ItCl0DHMChKZ9FB1/t/jG9CgbrLLJ0b6NW0S9sKr
retebycbwDk9ax8VKA8+5OwE8eKGVnwWTzDqrnBhuhg=
`protect END_PROTECTED
