`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jXtl5vmI0frdxWyTUhXnxVzVbJKNCk6Z2sf1y3s0xaMWzDoUoJUDk5WPtigtinUK
uVmjRe5rLbBoaSufmYUv9SEm9vjP4oFoVoaSuZzA267d96tGMZq7UqOlSfK5AMv+
DrQtHi/XxqDGwa3aovYxqhS5wwxGtjDvIqZu2bOo1X/LpIacUXwjaA9t+7AcewLH
tqYGUz4PweH0yiXLwAKl2BNJu661FUMBvUx5uXcfPAAdZP4zZuuxzT53ASY4up0A
uQJ6xXqkI5GeM0suJLjr/bj8UgetfU5gu8XZjXdxes+IavTEK3/UWjiLMgft6/QI
fPZFLzmaZOgP/pEIuJhBjdtukm7feE11zfirUnfxCSx9A9/mXIr8h6pSiGc5sRuf
VQPVoT+HFMC38AKHjlZgKxLWdByUZpkMb7RgGObQH9y/rRloM6jEMV3T/dED+AKa
TlBgfB75b7ObUDjfJ21nnyhGd+AtQyWF+VPwjvwaiwmJdOOks2TOz0g+vNV8ceBy
ep/OmYgwM8hoBoSqLYMLVmQwblL533Hql+8dApXZuPDTmT4hD6ETZ25VtZFcaj1x
n5iEFifi/FtFB5YWK+FLOrofW3b3pLJWABbMp8Di1ZfQIJsX9DCTsKIEZ8m7z8cI
bqq5YjEYEkjg1eXFpO/ZIk71trKAQIcKD33UlMED2Yg5ICXcPLKOX2ojqu+Nfu6d
fIs8aTTVLSEHbOaDrZxrxRndxTzQb9LEam5yIrDNLxXSMJ/7m1ZepZglinj9SaYE
sWPTyuO+EFGDRlseAicc6nPRi0GA6OP7hfQZxWlmD5kk7l8FKC+8ELi9rHcFX/f7
ZUtlO1nKxwkBJkwt+hwumDh4eFJxRx6onN4Qe1TmQc18vb64lv+P3YKQmtJ7LXuv
2nP5IBpfOfZdjBUHKpbsKkton8BgZzPY2hWyTBo9AkjBFYfUuEQXkcPi+yQhjIYC
qmK7xK5llX/Pab/WPR3R1FZCOS0vtjdtauu7S5ciPm44cdC0JXvaW0QW7r+3NI8p
EaPef0Dk7yALwJ2eLD1Q1AfthYIlZE649iYjmzJ31vudDqAsG1wY5jncAoojnkyN
bY22ki2AmXPFLn7z7eUmZFSvsP7Uf1+k1lWCP1hMcq9YVaemiqB670Oz1iAZ77bO
U5AhYcG8Cub2fqX2+p5ZxU3xtZOpq/WyVires5dgbd2/kNEd4RbTlxAr65kCFUC4
4evGVWNJPvskbeWJRO+QM7mtmVjvDq+bT8DxB9UcOMENb72oGZ8tC1FAtySqu2qX
amk1doWcOK5sdCKWMF3fFGZUf7hAgKV6NJbptxAGzBchKeRkqZdUcjtZiyvDXK0C
GtXCIxHs/p+9wewPJEoG53IaHP2nrdIRA5FJz/gvUgI6GKFEd4iS+DKVmyJ1XU2Q
Z+hU8q4IetMUSMu+q0pga/wF2y/CjESvEWIK6qg3ggypZCdFgoNiNhqTnsoDBcSA
Uk88ULL/BdMP2pQfgfmg3HRqimyLBqOluRrQKh4lRxE=
`protect END_PROTECTED
