`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHsStD9zEUZEfjdqnddQn5/gBqvI+35McRNsoqEAIGEGLJR1CmdZuwg6Ihavz2Or
Nc3YrqPaaPsC+SVNH8PPmwGk/x8YR0AvfxG+2u1m7hXAlZSRJw4tG/Z3YcUQum5k
unraBnEmvajF5h4WyE0DR2u/1EtRSdauCJiS6+cFP7UtqP4UJ8vtYEwjy+kiyg2S
biR2KQyvmVY4+bwsTiZrNd7d+lJ3mx8JU1lMi7qTsP2z/2u9xJ0WOC8Jjcv4wFFn
Gc9Y/xMpBw3cdM3XS4Xk8yWhOFZwKRiCNonZeyt/Zfa9haRUPm1ttIKBKvz+cJGf
+qlTOyketKmPmFqk68Y+H54/L1RQ/pIH8GZiDtdy1/6u/kBHtiz3wRqXZCDq1xtf
9x/mAkaLzLJCY4/6ptkaguhAoqJGLqWC1+RuzeJk1sMLbTBXg0+5r4L7lrgymjOE
WyLBOZeHjSkgcMY7bVMbayHtIQtuF/5dJUguo6qrQdaGbL9TM7d0Wr7WTnGSuS2e
i/o6ypTz9v6kkZ4nku0RZ4RInLZbOHoSXH2ywKRwtff5ajyV2jySzPPTQZKZrR3l
nQGX5Mp6xIraZNOjFIrElZ4fgOB8shFrWDOORQjsar4iuxwqC+VEDCztE8c82F+V
u7jA5gsOzCXkaGTxARD/WOVyMKaRTs3rvnkham0Hz8suyMGuwCpFRVRazIlZEkQ6
VsMelPDFVrtMsdflYcQztuiOKzLBx5FS4ejXnQ2+tVPzIxLC/QqwDv95PtgDqv6z
cAZNOcH0QfGpqq8CO8nVa9/ycXV6PKOuQn/KXmD5T9U=
`protect END_PROTECTED
