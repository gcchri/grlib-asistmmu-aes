`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZWCfrix7fyVFC9i/LsFi7eU5Nxoc23KKKkKYK8Fq9NYCgq0WC/D6Bu5hFCmnZw+
DndrdfuddBdhnOGpXN5bQcl2s9+2gC7SMqm0DoLUgJim2EenSCPWowzDO780aD41
20gkQyhOJs3nuFxG7gTEgHy6GMH2a7oMlVeSlJxgxJjHOwqarDMsC8kcNoypjIBu
ofp7rOS+rccrZ8mgC40fUuycCL7NCb86/lvsr8wospHksE++p1d155+wafLvPjYF
UojVqkh5Fmb6cqbCR4JLWT0DjVaj4e3FnmMie+bPDPDHGw2FZF0fL8IS/okskIHo
qxNqyjsqIBExLdknRV/rOw==
`protect END_PROTECTED
