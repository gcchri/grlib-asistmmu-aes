`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+FRCg8rSfFaw6qDeByMD0D2dB8J2jTOAFX9Ac6ksPk3QP7T2KuitE3lguagfW0V
9PL52GLTHAcUH7DIxOSCLuLKCQx3I9SRo+JW+A37iQBpgII3rDpMV086IaRwKIrZ
fgh4U128YXxnCWkm7Eh9Ad2rtSToL6/PIhOHLRlb004a3T2JWWYRwH/rITbse+Le
GdYcuqU2h0zxZh7yiMyF109RznxazmV2JhtCyjmNtHtYVkyNrXZHll6j+mFi95Hh
LITXHyNod8zS8fBT3uDjkuWcTfff3bL22CNYUe5kSgo53jNxa2b2vEkjz7myz2Ac
GoQlmQLR3lsAMLcrFn1jFAD0Hh+IcyFdy0pMO7UpMtMq6MAWo423zVzhArExlsII
of9mxvNcSY4cwyGr3tFkrnr1JMSqV/A9fcfasOx5n1OjvWKsJb/8niA8luPsOoRZ
S6Nn7Q13kNSyiM7adVov78RnjrlBljTTT5TelnmHU9GwHWQaGjGF/GCWXfO7VlMc
y4EHFe2PC7ke28cQMzlIJwh4GKzWloaUR4eosgdn6Yk=
`protect END_PROTECTED
