`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XO8XVA2GxHdi7AiUhRbMbmAPXu09/ZUM9gfwPGWfcGijRo61VBFm/7jDATpGFZ/
MewAlJfc/leRp8P2XDyU87aR+xSXOslb0JIbPajVw4RJXgZyH45Th0+dqkUgaqrS
NtuRzy0SDD3IdsEIR6gf+KomG7PAbPI+o0iHuKAZiwS68C19Ih9rvD+MBwr39mi3
xjdoiYsJMXHbNpN+sjK0C/kRj6DOe47ZPuHZxP+PpiVSbBdxLmqx1wXnYd/aCcsR
pCL5K5bCakN/mZOVzo5Pn0FEDO5YTnet4mbYQUViXpZwDcITfesx6ywZ18px66H4
LOzr6k+qP7U+93Buo0Dfe/HayiXWi5sxYUA6iH4SJpKO9B6ZGX+PUaAE3T1IBPRp
qOFy3WCbk9AiGSyleDGzr0FeNRN1/eNoiS3S0JitvOQ=
`protect END_PROTECTED
