`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OUSYGKUC5B/wYxjq/NKy9lkQhagwNJb5UgR9dpr3moLomz/+sxVCJWaDIToaUCh7
DiRd6vSdSw+TFVUbrBMBDwamkI2RMs3dOFq4pRVuVEYvimgxsIG7k+0lOC2mQRfy
grqwfq8UtQw+QyEB6EDTGyDFKgPDKZMrerai50QaVlJYx9JPk3vb6BEPXFd0aTNf
vwahv7XKfTC1jCbOrmQWowdahx1CHlBSDlBY3px4QKOzR3jfwaI0v4f+QaJI7qap
oMDU5vtTqsNGpoXEfh5N98/4PmPKU3TNGguIa34ONBIqrDHBCynY3nZVr9k9xq3s
qwAsS07KB0slelalAlqUkgaELVPw4Mh3R9kZBObR5GRV4oWdsAkHXxTYWLvg7ZQq
uwC3P+uG1ezZIYUBpdvDJmqVrH0ZBQH9UVaMmsKXFq2ihxS8oAmxNnOY0bzzHlRD
qgs4Zgul1zAl+3MyzDx5K7tjROcQGE8Qwddd4BuSdF1v8aCqN2QJrM0t0TWIZ+lD
NPzmOzcPj21TcAAGLH8BWxWxjOO4Wd5KYf68IjWr8SS5qJelnxn4NQubj2plZ9Id
n7aZauMdJDt9iN1YBidWRQ==
`protect END_PROTECTED
