`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqZYBFU43Ngm/Ru7T3L9yGtbS7MCgLfKjd++Op7OFrK3QQUHkD48f8zpc2FD35jy
PNxCMU/vJjBO1+3Io+Wp1pSu2kTD6BZYUAB7p6ZWwiPdH5w/TrvFQIAUdvXt2uFB
MbTXmm4MkCpSZ2nZ+hGACvPEw+Ov1q5SCEpNASjmAX6mVv80wE09LgrRUK9FBRFv
kbmRpIM3CApiLDfSYT5SaoLCeH9BxTXRGjHHdK9yWzvpqCOiP3FEllq91v3CS/RW
i0Cb/yKWIFV46Qzy9fdISg==
`protect END_PROTECTED
