`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n9LxHnSl3kqo4M2vOeZtR5b1FUWwvn9c3DD5B0r0MH95+fB+MGbJII/9Ic//cLaC
+P0Ruab2PRUQ5QQ7n3ZLKJ5oU0yhAClpQ0iI1x9BzDHo1VNmWlOM3ka4oueHQPCI
AA5KSKuXr1/NtcpjICYq9iqE1kJrgglkNGlUjsarzalyF5sOx/y03NG18zA5udYA
9iaNVVBKhkzYJZFyS7BEaIiGuZYVY9bKwAisJBUWqP2X9stz9B3yTjO1ZJ+d7/PC
7Ha0rEH4L4Pb9tt6Wi/+iukxZFtIHkiMenoR3HXKM2Q1g2LZ+5ciORFVvqAOOGAi
Ut0TJtDYyMkxGIeGnMMTOTdO7R8vGWSFL7YPJolVI+u5s8sk/Sbr/lSTUNWfiZLl
eLFVpH1uW3+ivjIdc4nvubk+TwVCOzg/pW79KViATadQ2jcO3aMJhh+lUHQswklS
smqMQ2A33E2irX56zVDwHk8cX4KHFnSSIGc+5l6BwZJt9ujpb9n5Mt8QrZqW3TaN
JnLUbwMd3vBdneIwyBdPbqKgeVA4OmmzgtmZpY7FvEhyV7DWQS4Bi5VmpQobE2gr
QnjfnW6L3LawJWO6yLZ/CdCwq98FAfI8MS82bdCzdI+IHMr4ulW+CLtNNqTN8LUt
6GICEFYsCKoriPETVVFPjV1AztKI/rxBpgO5KvPbhShXesyQyh3xsE2JsYQndSrF
dEqS8QcAmuibW42IwMv8KgMuhUWDCpI6AE6XgKiF/OC4MR4+2q7wJ9CxrjuJ7uyH
72oaxf97hqY2MyYM5XLwO5iulkpLQm8QYPiIzBq0kRpCm4Buoy+aMLCW2m257yHO
8WHuiix5Wf0I1hBK+DU8VeKTiMajLR1KlBfGvt+7gSFz+QzyVyXj9fYGZtgV8oTI
J0b+5DPuq0oApH7Yh0mc+M3xHEM9lEuvCc7s/n4zTIQEOuahh+YAq6BGnlLwRhh/
gXSEoUz5BL7Mu2neitNdjKe9SMpVAk0u4vzjbeezieq/yy2tEBpAbZmef+w9z+Vt
ZE/5HZLzIGOwIzM1VaFjzmGgqytxWP8fP31DYfiM4lj7OQP6pDGnRcRavaZG02s1
8Rxd+kMNfHPcodL7IoPmqulD2hGw7KFBQtZsltj0d1obMvNXqWQ4iyFto11Fi8OX
qjCzRBkTi/Ap40k7W50WCyBgmCDlWVvkoUcQTw0o3SAoxZJp3QC/vtV2VTKgHHMc
istDlhQbCzh16zjRtxc9KQ8dUSHiE80383o+EcNNm1jIQboVS+Lytv+X8mfl4E6T
TMAAIM9kgT5fFIJzCxWPOTjjp8gndtxIcaXf+zyq46FIJ5Uw3TKC6utQUDbr8igY
/dlzPeUZwFaqvF1JGLl7tgWurQ151FmTLbALI6h2OBwgM3soS4TIkhD7S+pwIRef
Jec8JTC0PFw6zQfJlgkPDvOXWgSWXNq+TgrvhwrzFLpDdNZxCJ2cRJ5Sl+PTiyTH
fndB/YnzqMOPPkX5/mXb7+txKXJsnRV5EtT8QV3axFp7z/ZAtAffh6OhfVqGRY0W
`protect END_PROTECTED
