`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3KHGWTPQbgmngL1z3XWoxvqxBqRvuQDUtsQ4twfpRkCRLeocz+aFrjUNjTO5u3x
6S9bUXnlWY9EdUEJzB4PITTdJEquplVqPqQmj49c5yr461BX4oVwSqzFwN2y3WZ1
mczJCVu2HKAB0fKjn42Vesi9uId3kZaq/wnd0c4l3q50BMNMmBODlQ+mCAhxCH5i
TpRo4Y+9ExhcrWtGVsQyS6pqkTVhxjOshIK3AbqweMVepfrRdSK8FPBUzAC1HtaJ
cbREMn06Bafjwu6qbjx5doGf5x9wyHD6Q8l+wJXWSqSZnLBjN/qk7vhauQR/v112
HFXCqn6bRa4iGzmM6unpo/FKSzfR9AgD8Fpl4pYn2QKU5gXK1EUFu4nEeYUAdSem
ZtyBRdFv9Onb65iIHo3Sse2+6nKyrBVHT1IcW8p45vaY0QDOHDnVcdHIOjcXdD/3
0VhqvXLdz9/En7DoEsrrg9vSLVIto3T97/VCW+5HBjEYZ1EOTa+KV+LDmDkTCpwq
th2NCBdNGMEGaxog38TM6UVBpRxtwU3coIBDwO5N9aqKmSHvFTykYY6f4YnOk+jC
jG4quAWWmFqxCptkkKCKM3RjYVqKfA/T56i+mb4ebmkboRaTZLTSZEaEGRfKaPhN
2d9DXBLCY5H7uORtPVKXUJ8v0vyXOd+bN85Oz329lfgdPwcfJVZLBH919VBLwb42
ZsLVbnuLUKfwLFRHNqDJQ765DC52oNYPudkUQQ2ymFGYYbteLB1H1HjDysKnVPBC
ob3Zi5tGdBYQ7DPm/R+4keiC2KvjcnXDK57CkhOLnEGzh8gmxmKKbWiQ/LPbvynA
Zr1rdqkNEbq6lKUgMiHwsWFESNNft694Mm76bS9ypaBMgDTe7/aLY3IEqDD871jT
aGnfHIsrxZ32VuMW5eWAXpHCwPfgzPUcuJRaP551q3q3HDk02uCp1+1v/5r60z+Q
GIJdBLi+M9Ynpr9zuKes/mYKD0CeAoCgo3Q410loifQqvm7t28WjmcHSo/uG3ple
RfbG+icpK5rqK0O2gFI+rSkdTCY7h6WoCYPuGYbV6UMLcxWSrkdRg8lVAShbbfhf
w5L/JHRWGZMSVQzqVD5woY4XKQ2CW8A+0v03du/CUAZV55E+ubX3QuYakweOC1zP
CW6V8C9E9N3/2iAiQVYW7H7+C0HYjpDa78BCJJFRb2mfIIStCXnqJjVC04ASpBEr
r97eYJhE1XFM5eKyovNSAB13r7qAXNw5kIs69Ug2dItw2emSVJ8fxkjfuovOIPc6
ut6V34BsL+QDKZjjdpip35z87fMjjVfKBZJ92cQDyYv/FA+3gkYU/hRUcA3W1c5K
psWTllBHAVYLyOhDptgcjF0duzc3bikcQkH+jVjAeZr/3HZ1B49thrraITAmeC6l
uElJD8S15pA3O1GkW9WzvjbPYtej9ixxgCvTvahZcPEvm+BUes0QTx6AZ75F9BHf
nN8z6P7ZlLgNqGJCHduXHexGeRES2U7ZiVqqxNWfjT03ZLsKDUZiELG2/bjD35V1
BR7ScrFUaAyJqIwxLF8Zweurq3tJqhzj+necOrNuWDy2qOoBz2Pc5ShNuDyz0AP5
eYCoQftUz3lOmPPKCUzNz2hR3+UjkgZccll4Nl1LKxqbOXxo06UaB3a0Yf9L4sCa
yfNPHhUujXuPyQa8jBIl+ddYVhXKZ40L1zLOEucaY679FrUusLtOxvjiZ7WsDW0M
y5Qd4413yZ2BBXgnFNaSNdXaCkkkqiZ53MuDZCc3wR49lsNZfpE9Qy98Xca+yh//
PNYVL7xfdb6Uf+q4RXobweUyQOo//X4uiss1V+ZrtEVn18UzpRQ5YYGBSK9LzZAa
RJ0CTJobVJ14ghahGYn0wf6Xqgme1OY1CPCQpbM5E+cxb18YwKZw+ZIxK8NTlxmg
56HSPDUmleu4BfX3lEQxK+2L91CVWAODI9+eMOUON5Em90tnxIv+enaL2YAdP3nT
cn9vFPk0WyaT9py4H+C2iI8hCpGMeT0+2Ees3eK10CUVOpnA3YofpxgLpbsEOH0B
fIBEl9tGGVHeUAnf7ESp7iqNs4ZiWLHPHrS8WrFyqzGqwyzjpTM0kWH/kOnhXk3T
ZGCzCpeMsYhuSptkIeAaaieuBioI+YCq3IiXzpHSWyD1A+Ch0SQOMMP6cGXeWlrd
CKNxeF5hZ2mStOSyp8dPslw3wDF2b2mxo8fI25BBsuLnvv3xla6u8gyfh/THcc0K
dOZYzNfWfMS4ANgifPtsHjaQdyfuB4X72n714kfWag8ZlLWxJDm14ngH/58akshS
pvKrR/nBOcO9Fdxi9V8xs4U/BwEZD3QfjvlqlRi6JTXfjvTXd82YKLbfsaGWiglK
9es6IjRMqb/5J+Qxe9o7h8lHGgITXnKmsNNZsDTw+rzo5VH6cx2ZIxJrgsr2Zy31
YL2rFomxC/sFQRIrA4igN0rlTvNT6akpuAXl3Qi2s3+xC3QNmqLejSUYdNxJ3Vv9
e1nNgtV7nvtdVUpGLtbm1Z/e8D9Bc1501xU44ugH2xZOZpDgo/ipMz3JrrLNZwOr
UbUwBDV+Avi30tx0sPWJhAcjPmcedpHmvdV8Mx0XXZU=
`protect END_PROTECTED
