`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rbEgqGVJ5OP9biv+7sLe0Ph8KlRFj8zsf24fFMJkjSYZHSmyAj2sDMgN7n7Cp0n8
4qhcLqtLIe4Z/SQRyQJlYzYDNYZeHOfmp5N+4SCOan7L75y3OFlsbxyxaSUGFaoX
UvCHRoeqwy43Fio2yJnPEzckwIKVOKST7aHAXO83WSvX6EMIJNUjySWGHcJasKK3
FJwisGgCMLti0tiBPaC8VxwZWS4tiVIUVQeHlmv/SCBfRahDkOoGWJ2UNO52wRs4
IL1PysPLQdVpJZ0aUtg26g==
`protect END_PROTECTED
