`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hNNLA8+b0TjsgBCCVdX2lB9sM+u+qCk7LpIBpJDm5EzncC5mugaAgEdxGEp0TbST
eGrV9uT69vCXqf1F5PlBvY51ygLgUYz0JvAyVNu3irFOSgriLV8HADUS8AJl5pEu
rczR8siWpXAy+JgXcDNxGGUD49XJJxFApnwxfwz2LaICJFdaQRJS939FVqOKa7tg
sqf/2gwy4Tv47d22ms24OSYjuphoeY20gKXiMn5B+N85rlvi59i45UPm5x2hCfsJ
bq7E7F4o5gUo30jV61r4FyBq3JmByPKhbZ1Uj2ciQvQGmA/Hg3934wxiSNvlnrOV
aoK6v6+0WpReiEudvLx7+wARIYUi0mvnN0I2sU5ozgsMCZ4LKP1hSRJiTSEKm6iW
DkpBeX/dx8kqC3zJMzHX23NOh2k42/VJii1RDpLRrda6aKbVrKBqJkSQ1nQgbWuq
HMrkU5HF3pjv2GjhnGlstiUVi7Eos/upeq0cSADNRM8=
`protect END_PROTECTED
