`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3qP1cZj8m0dqebdZdgwbPKhwmwwujYtcacodt86qxz1GG43obXK/TIHgf0/L4QQ
WRDxyttycOGrUrpsXzuRx2u8njuuU5tlgX5uKVvkuIsCDiGgJoOD5QlcS1U7ORVr
jeGb+VlOYXzZGRNViho3zxwsLy2/gV6TJTRzaWneIlSls1+c6XNisEDNkl/OVLTg
X90HgtuSC1dtJPIQEms4l2y8ST3z5vbfxjYKmsMH/peLoJpzEc2S6kw3/dxM/8fo
tin4y/D2BX/RM3Q4Bdv6T+CZhVLUhTb9JT+axvGJjGkG4D2gOiA2ebXv3jDszV5H
vXZmHWuIZrPrdRRNbAGQdi0eSIa6TeTn6427g1ixhkTP9lBV/hFtASR0zYsOCyLh
wcVPo5cY7l8j6XWtDcYrV3X2luihNLaKWXCVw6RwiuTjaLUKJLgCv8/1+Ows18z/
slERNL6Aiagn2L3uEd8ykqJIgCSMzz9/vYOD6hboqYg=
`protect END_PROTECTED
