`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YdaDXKXCSsNpbwirE6WPs7DfIb40fK4TOS+aCGpeYhYu0f2sH151A+X551lIGebj
+ll6QYNCYnBiVj8xvjlvbP22QlfDaLw/pubY/uiaAJVWyDPLUbvhxrgY6G6cZNe2
kNpzys2bjYh/MTFa6T+kBT3xZHBQI062heB/hXbODzyuwDc2Rq9LwWRIiDKFRoX/
GyP+UF0XDu7ADTBwNSYPX9OcZvIfgsi0sjzwYV9g6BLRKZ3GXyYqSdvJgCcV8JFs
q8dYnTC7f1bpBWk13IQ002eEdSxR0ZLcKt2JnI/ZpDWNyP1BRoFtKASObWUTtrMX
ieoE489ybhYA0BUsroKiW6mtn78A0KDb4Dgy6Vnk+OGOOpXD7z/w+6Gux61Fwuhw
EpMB8aYlPDAu5DZOYN7w/QMRXgbrCDlP9ecZDSxHwhVKZm6NAM3c5UEfRWT49PID
`protect END_PROTECTED
