`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfntj+nJCjgSGHCavm3paHCxNYe0lqOY+w3uW1Dkt6TnzBclZdG0wMBhiHlCq1+m
lCq1fAEw9t9kpWXt8Mr8MbDnavGwI4NU3uSJvJyIcCxAMfUihJY3N9vZmw/Tvrfz
xX0MbGV6Wff/CAYGkuF0v8kfICSSj1Klc/FoeKUhM8LdCdPo/TDpbe/Fh/prpE7c
IbOlHL130eH/Ocjrl4KaYxA+IKidiemzMQIqXXD0UzWs504eT3p7PRC5Zyb0CrKu
FmH1o60WasjzjABi8tyEuiIxQMrNNCsWvurP8/YZ2e7Aox8E8HIaQYM9UbFsM0yh
X3Gt1gxh50XTo7qWpoMUndrF3FaKX2kULimbxAk3TiiURfPA0oNB6ozdLn7Y7z4i
XQTokv1orPnfsazNL3JAkSY80Pt+uIFes1qfXfPlas+EEezACctQtvF5z1eQ/vWn
tBy91qYocT/fYL69kx6L1OroUczejhp2ZoIumT1nxHHWP9svtz0WuvwdZETPYkNT
BytFKXj7B8huu+qlcpVc6MOZWttWxIkj9CKq4iMw8Eena/dyqTEqyZWSgcgt2AHQ
ajzWrh4FzsXY5s/I/faLAuF0vKpXfYoavIGvFG4gKY19foWakjsqPZnbsi587M5O
NozjUiB3Zs5WDcQjFYw3EB6Az2pqXyxRrwWca4diDiAP17OLNezROPUiCH0pWsR6
dstaLDNReGtOZLcgGA0fg/hagGbv/Rn0gjMqx1+/sDup8OC8uxUdgKSO//o529Og
/+J9CPZtTryy2Nvh1ZbhSiCGCLnb67WjfZPiW0qFpwtanHlgJg6DOYS9B+T+HPja
bzvHWjpSQlGxsq4AsTnIKzyEVHDhoaEpcVYMDlrIEt9jU/9eCWkF4tsci93e1C9u
Z7jNhfUrqw4j/FQGC0KQk3DiqpcVGvW64fu4SW2k535ngv9HHwR3GfaVAIpHgjn9
nJwMoOMV8gv3/BJ0DNwYXEnXSdTBi4Ej/ye4UK6++Qvn426/De7GtvOYThedqSsK
fSpqPXLn/dx4aN8jzW9Tbc5Kmx9WdtsmdSndx58E2Sj9efoGTDqjQCEAJSqZnROI
jQBpIzzHAWWDr84pNT2uqZ6ET5Dhge4XUQQVGH2tGSAIC9ED4wLdumUgpQjaLyIi
B8Jk2zhmWlF/364tCxvSSgJoxj34mLN1b4R3eS7co3JNVKH9fndQsa54aWpgXtqS
BrsSJqtcnuyBBHYXbHevm9muGvxEEdz6FsN9e3a38olXO62bqH31Ze41KqHFh/ka
NL5YrGAZlNt4OgP14twyVSfO/AL+8LuGRiwO2Q7qAv/fQ7DdyENMelAScODYDr5T
71L3qqO6YJpl08UvL2Fou21beonNiVVtlExGe0tmdnn7pMijQA+GPp+FM/CxTeXY
EF8DzpX/xXAhHiY8TfdvmFDAoVxFwVQM4wTnirkPP/yE3onAPWvS8XKP4P6e+86F
eJWUJt+fAW4FGqRGfEeAG9NPGiMxIafIw1PgfxeZcagr0npjleziz+k+D5tH4uJR
W7nxJRYqH/0M6dKo5O8Fzhv3h+DzU8BYRzE/c8trdiAvcL3vQ3M5MFuyQ+1sLg86
TRU9L1eq1cqZdXa0r2XL7M1HIxz/wdxNktSmo+tShqCznatxpr0cMRJejpVOp5uP
/Nkv74j4/2epkTB+eseXnVmb2MSg5NpO7RoOL3+jp8vfWF2e4Mtg+/mS2UDBqUKW
MczN9vytQLHlv0udR0QgBYujAOhtGSSizjJ5pFSfm5nm9zCRxcyQ/K8pVvve4yN+
TmuN49aE2Jyvep1jeCPOMNPnA8ujZZcGHoHvHJyhH+Ea0RQA792kAE6tf/TkqjdG
Go9U4FUqWSN4VCHdxb9gWF6toWZseRUzw0RAXoeM6rSWPWi7lVbg/cFg1O63dRgu
S1HlB9uKh08U91WY2Mj8FjcM2RqNxFHXgl54AIrgNRPi9gnlNlsMtYX7hlBJn8qZ
cPlCBpHkZMKlsQZpuI97gxxZxsVlbWsKtwz6A6lmH2EgzN3QX9p2NrhIe1hLG2Jt
8J0wDtUzeu6+HwEuW3DDljS68yFOkteI77lw3ut0etb/mJUDcots61D1Q3eS8nGp
LtXNeKi4yuXTM/CQCrYt7huK96JBHpkcJ2NCkGuf3gIlwnsrC8I6fR40ikiOlQ8B
rwxXXfvtnEyKL3Zvzi3iE+/o5BFffEpyTdh5+CLjZKhJVGIDyUsw4Q4tFpUUOT28
U45l1GQKG8bvmlGqAno1ApBWgBSI4GH15Y/CgJB/40hP9T/rDU1s0dwBYQGx7KDl
uz/714koWjkH9o5TFlXLhpx96y01x5nC0GPHSVAgQkEZPtrCX/UnoM5UKzjHTUAK
1dPULy06+QW3Tp9yZEpJcHFP0MfTatv9aHWR8uxYDYVSJZQ2tRp+aj02uL9CZSMx
w7JT6/lwEnPyT4Mmf/QuYoWg4GKSRm8ll0cv5ZRlvByBhvEwxSiBJZdxYAlKsyTx
F8iGk9Sf0OXUG2MCxovafjKbEjT0yq/PZVem3WCeVdCCXzcowe/cHJm0ftylwp+K
dy+MXCRegurjjbrALlYP2oIIiRk0jwSRNQyxnQVJgxrsNyUiBpXFhl3eKYJMfIVB
+G0AeuB1yNrgan76AIyvoSboVc69KKrhlQB3pdCOfowtKly6WGVtogmMrjlu+LjG
d5Vz0ontEy8jihagxnI9tXEUjkNxu+xzBV7iLOYO1eZv6G45K6qlAKH2ZoECc5vr
kpv99qfA0ROpAexN1T+h7RALccRqjUZF8W6lc3E9GwlOhvDb0wo16QGOkQZKlECX
OJdyhaeAStkrPg8XphzYv3HsYbmnh2mWHyLvQ2vgDN84qQZ8t+WGGpjldY9KWt02
kEf0P5hPbHO5al5yV4ih4c97h2VHjIbBPUYtPuf8iXPLxQyUfPVoLGyTg+5BPv6U
KkRO0gEEgsrg5C7nD5KEMljQWlpaWaqRG0uNnO74GhkNH8LlONySI74zVYvrANS3
vXr5XdVgY1pqqc5onfvK6fSEzlBde7D/TqU8S1fCEFXKI12UrU51RDY/FgwXOzi+
shOHENNNud+Ul90MaChY6iwgzxNqm79YyyZ7cYUeKknhZmMWaA69UMvjb/CtkNSv
jtZ85oPlvokb95tUexB+lLb4KzF53Qf986AqdrgM0Ysw/NpT/MKeQmLBOkpyash9
roOYyW6ji6NjvWm3Z8YPB90hIUAeXT6OfUvx3WI+OtYItCNkixDIxoY22YGr7aHc
bl2yU+8nYQINEgUI6jqz5bXbI2kJY/rXxUbxbD7j8VB6b6bH0E+Q6joAQuTYXRCZ
Zl3iBwLqDvwRBSeeLTDvgbO0aYCKdmL0293Jb19jpyYOjMr8qqf3r2A4FkLAq9cd
GLOntSDhy7i9nYYmr/bR/Zcbj7cku1L4aRUUJfKtZ8+oZPLKsUroqyaUs7XZjwJp
vML+HiZIxo1NVvbDeOM4e0O+pFyrtYmgaipKuGT49d1WPo+Udv4tIEzxCQ76472Q
UFW4ng8Oz86/Wo6zMckqc+LcjYVB50UtYK1QV3zAqayAhgLNLsRuA2NgnZRKS27G
vxzWAX8VkTGm3ivnywp0QHjwab7HI61jnV1U2/mAHNw2043Vq2uqhDYRs7MyvuvC
ODvpEwfFflGpdnwD1VL8DUP7rWA1sQ+P1HACD0DI+RlguwpqvwZ6w5kmHiTdvciL
DCXFnCd/0F6NUtoI5My2IjmXv6XcaIRnTuKUZOW0YgZrWAnX9G7Yct0YeTf1DlUF
9kjtvgaLUPoDQdfE2u56sY25PvoLiD1eoOsgPfsyRjUMHqs0ouDM0tkX7RMY1QaF
0yylSQKGuyRNiSrB/lg7H3zeaB8MbExLma0ZaymM5O8=
`protect END_PROTECTED
