`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHpng8rYxgvRI/KK9X0zMHGmQ4R0eSQNJXvwpy0IS4aC7RdVAtLP9g+YJIfoseCc
JjcGcgfjzK5JrBR/ZWSvrddRjku6FRlpI0SAdisyYkDELDD7W2EKiNLha27aaNyJ
xlSljra1LEbnu2JrTgr4J9jylOvZV3GyaszJGKewFcxXhnOZN+gAc70cOtQKEuQG
qyWwmpQj33CwlP/Sjs2o7Z67hEPZO6ea0ZNfZLv7dni/VsYwYB7dhH4smvXkSZJH
tCMzDIGH5jr1BMJRqWTzl6x0Iz3iusM4zcjmhSN2P23etKUhL9c8PzE+QuyRqX1/
TJVf8E5FwRGXzlUc2A5qf2sV/AqZbpiK0jPrpSVJKIh8NX7022d98QWRQp5erYPH
8WlHdRWCjOeFD6JO7Fo5tmuqXHucfCBxSAyU0yAKBkPZd9jma9CGhzbZs6/HKwX7
ilvLZnkVps5260VMu6/gaU7AasbLxFXnPg9xuoEFTuttOuZq5SBhpB6EaV5GlAHi
sIAnhtw+bBEOrfcPJfq2gC7IhO/FgqAFk0VsYCZjCZLc6Ci4QdO+/UaRbtqctIX3
2Qvx9P0Bzt1Ih90GaP9l6KHHuwk2Pi1579RAWPxXR7wg901TgxmFhHSVj97ZD4N5
vp72lHu5fqwZWHtlF7g9p4iZ+YBO9s9fUE7FppHIbK8duu3HCKB4yGzg/RfP5uDX
phPjaCYyBTl5pjAUrwFgpypIaHhbFNApucMJ7eZdAp6UwsgKhP5Tfiq3XdO89pzX
8QgV4oAX7TdwF5gztNrn9APOU9e0tMstBmJRNk1ToPRyLgHSAIdgvHM8IvYhyvWG
Wtmw9JxXOV26jh1yZykHsgQVm8DnQcV17Uk3lwBqhIq7vcVcDd1e783nCbm87Tm7
tOkYrPihxIZcAxps8PNuMWjPJPD6TP20FHjKo2qrExCYtDguyiZldpVPDkqmHvUl
cCLp/+MjHwPFP66VR59GGq9U2aR44ty2IQO7n9CPei9gggvqa4jqua/kYa0bSXha
pIJt7YNU021WniI/w64wmdn8pz4GruBXbSHNJXlc3cwuAofF/mwBDyKdq6CGQgxr
Ia9dyELUtCFJVcY1nGT81Qcs8KEMpbg10dNTAS21uvw+gTWBKoVSsFhrgqhlp9d6
p1vdK1n7QHAqD7dpxMpeYrqil33ji89AVmWQ2OZ5LjpvDODb3G8etam5QoKn8KWV
wCL6bYUnEuAOKbKevt9OtMaHqjt1E0ZglE9smYyojZtu5t6FOAluYCENNRwyNEKN
XDxfWp6OOfc1xFLzo3JiFoNPYSnVhy8TZHTpfBZgl0QUywTCJFEpK8l6PWl2NbE2
DBi5nHhCZVDNDro6QiZvaqyiTSNUjBF6r/IoYMLdl5Fs6TbufVJttZKZ/bccE5X0
5ceNOuhtsh0Dch1JnSiYkKG0NLo1fwPH1bbMgLVj2FLdI1nQ+k9vxv+GAecOU8Z/
h5DCRvGQ1f6Wrj6vTqIzJlKyf9pdezujFvLpGMPt9EQnwV9j3vIrYkgbgPyZAwFN
AVuAPMoDJy8HQCdwezx/PfFxHaOfyyKe26XcjCzjyH+tPHxpaT2wpys8w+cPOoFe
iL/gOWrOaeoeRAsbgmyKAXMBwptVC7Z8S6o+h64pcs5bw8d7+Kvc54Bq3xB0WfbY
t2NAqdJ2giqJUNNfXHfvNI2S2rsHcEBgyhPXSQfJq5XRKvjMwI/57fNa15JSh65O
Lu/rr7uOfNCDeGUWP6xV6PEBKWfXh9Eh3jq9LLlPGdamSCMBXTVUXPPFnxwQMrW+
ZNtn6S2nNefOljrs3XGtEARxQMW7ybu1M7yzk1XQzkiDk44fa6IEDqd0mHxQZJF3
xGuy+HfDtrdp6Alas4WVqDjWD5QbhvaAM2EDTF65ZeqgHgm2XZNGhCh7IkEq1OaB
l4sslROkZJbG9p35GMk7Lysm23UU8bJauPyZQoI/q10UPKAEHMrVnN+ZJ+p0VHbN
7QDewSEerp7eg2y6drrCxHRIy+bpqUrpBqJwlcl6LUB0nDjbqo6+7UlZ1Yqgc8tZ
5kFY/t5SJVKFipNmBdZLMbwdjy7B/IiAfFkVfnHmHwMYVZ3XlkfW16wH/wV5u+H1
jVJyjEIU1FW1x/3VbA0WnEuikPycDLnuULWr8nB/srSSf1+8W70UuOFIJByzXHbB
CXH2mATsm0BL2JhMIKGeWnAaGHcORf8QcuEUrdwe1bWiFUw+gPYOEWOGstH0jbRr
fYX87/65eAiNlmMP/y/7sfiTnwShpMmUfct0J2D3+9k5oH8Ge8PI4wBqqt7F7fzA
OXAPBupevu2jHwPUyCu2sFInoMFX3Qpx85DXIBKqXjaX992TFD9GF4+yU2JvIrv/
MZg57u2XowmZDvi6Eo1L57OGwtKpxtuxLWFCL8XK9N83U64W9hpJhEVY2YSW0k2c
whgOmHm3kTVvLeijUKc0MWbDUSz76FuessSM6wqP+UyLUs9V3yn5FpuFbcCazeqG
yf8iyGrGKShb2VfTsmkyWWYUDdjiG20mtyWtLRi6M0gLTG0aRVQP1ygacIzIwWSp
AIYFxczRamgUsSf3dKmuRExpkcr1u7jvs095YVCfBFoF+65BVwJBYYehmObtHyYn
gnNK8mrjCXyIMJ8hzjcKzaj0qmxHJxq7BbmbbM6tX9zMRFOPPr+sel/NP0UKAHnJ
VpjjTsEUZP9FN82XVVA4Dp8hfuyetdBMfc5uMLA4aHDmsXYR3rP5nrENmj6CZslk
LKZdhckpRhF+/SkKF9Xuo3a508TA8aq+ZP2X3pUKw2Fl0LQQdXPgQRcQ4BlCmOk+
ysBvNBL2tme6ppmvG2lpJYvMg88Cw5NWchkDq+Bt58dnos0k/7thtaobF4GTUifn
cZOjQ9bHztaHlpTrfM0N4xjk3yXf2/eDBigjn6rS58FSMJVz8+bpqnjK3EffjUUZ
EK1c8LDHH1P7b3flNl3DVJqNkwFdWTgonOxJ8U970F1CroasShdOiVWnhF/5g4qk
WX2zwu4OncJXxzz4tjzfDAppDQH6dKu597sd2mLLSqNlDmwteF+xPdow40/rg8gN
`protect END_PROTECTED
