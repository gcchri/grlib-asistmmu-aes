`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BuphlYDwK1KVwle4x1lL+0upEy7ydcQ7rOWdfAI8UgZCqiuiOxnxDeQ2/LZ+P5sI
yaDk56vsx63viSKyA49vKsy7nKuLj0CsMYXGQGvi8rQGGnjSYt8/FWhpdTFALUtT
6aX07uXsWk445zQ4u4g+r7LtLDOhD705iOySowC2Gx8BvsdCY3Aud8zxOWImq4cD
YIArudb/YZ/KpGndtHgl9HqslLAC9dxxPWbHWMEtLVSrJ98M3by9NEzp6msM8jO7
iMxvV3bo6rYCM/PfI4c8IhAEI1fXInPx47CE+icDf1HxfcLqxHtI/JlDbKsnnKDq
BbgqjaC95pe+UUZXl/P+iw61CXU+oqjXLyiwd4at6ryRFg+VHHyVvfYgo+MWFX34
qILZDm7vlQhJ/2kZCpFzQaR7uDxPSbG0SW0J/zZKf9ZwHRrfyqH96pi1CXcYFX+I
`protect END_PROTECTED
