`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RiZkb/35gSvC/AcP2eEVGeDN1D6AkibnMFrB1+XvpROC8KHCZre2yhIfM9afQREq
p7CRPwydmH8YJn9XyD3uLfvfuZAXdE7BZ3GujFKQI6TlDP5+xRJ3tITT+To8TShv
17jWCHUzk9+R79pEzsddRAYGRsQpA98hqKNCIQmvkNzR9D3PYfVX8xDuTckV/hOA
XwJs80cq1nEABmRXz/f9s9OMG/tpxA5o+Ubgvc1ots6uebDPYTUXhsOIWaiJ9nXV
xwwIvezurlrJgslH2bfgYnR+gy+jta8I3i/GtwTyzTcrfyxESmDyi/U1Po43XcHo
0jywfDXgV80abj6pikQEsBCt8tCUv+yKj8FonIzwO91GHFMyFgvAGyzLl3KXyxKx
0lLDvOxPF4eZL5huY8s3AZWbz+pmlgyOkIYsD4t1AdEuStCtG4xb3hRkZfV/hfQI
/3Pt6WHe7jN1tSa3R82rbjJU8GkT6bynHJSMbg+IfeDmxf7f9YpyUIjr01+ifnWK
xIKfa2cubwAbaV71uylG7/SWsNuVAD7w+j/ObbZDCxenyxFd2ErTwsFMgDHCp/iT
9Z5Xa5Tng3kTmZ3JTBNhpKAHJHEcfdvMBvA1TQN1nUcykx9rp3RodttnARHMPRWR
rISpYK3JmF8FL0vrKkIKUS1t1eiwh7RJbx/5eI8OoRXaHOFeYpik3OG6siKA42pJ
3PMIUyYXnLTNaZ8nqo33WYaees0AysXnTEpOwCP87GCtHl47kIp40OlRwU/URUx6
5imzG8o14ZFel95reKBoAQA+sBLo9Ph+m4Lak5OZc3BmMs0iK8PKu4WE1Iq3T95k
XtGBB5Wv8L6kPUXfPEMfdzwT/7AJdzFU/ZJFzEdVwLUuQV8hOPLxLNGgj5zYPj0Z
unAdcOvNwohT5N9PH+DBcVcyz/LAVBVfSSc6tRWjigV4cgT3rFePs6zoerJRGPv/
2Cep6jWsOrlPTL3H2/UqLeWf0TclZssVjxlS3q9Xc+6t7JaubD/Mc45QK/icblQP
DmjMrSCJfY/0kREMSvK+sQ6FIL+huiu5JygU2i3xSO8eBiJ562uLRz0+IUOvxnRy
RWsacfSjULVk0T0QSWwlkT842oJfjzDfJxUOWVxUnEG2gr4UpURbO+t2EMDzuZtO
RHgvuWLZDZ0mY2IA23zs2+p1abboKoi743mybAqLFr4E/i7GOE6lJja5qZZjG0PW
7sVIJAlLzMDCT7PfrjMLrXEHEEviy3cZjqYNAZ8/4KGza+SblSdMisFI55mMxY9w
IQTpXDLGnnUifFRbzrwyg5OzIC5j4O7y+kZ0BLXkoEZze1bQ1x1h6ObGFJ06M2Ye
fACyL07b/VkrZHymEgd06VzOrvNxZ1Bz8/OCjU0N6Cc2/a7vnORhZvQ3p/go1oi9
98+cKaxp67ycG0mJ5nBurAntHeSbSAiYZYVO8IZv3GncdjXOJLW+DNKehk6VNoao
NQ8TICp6Mm3bf6PCgKA2Z4Qz7xzbKtQYA0tIsDgjVSoVPZ13rN8Z2TEon3aJBwNk
hO9Sox4t8EwXxBUjUd4tvpS227Kz3M8SIOCv3WfYYUXZhOeGFuO+AqJA/kFXZGwS
71dRre1iyblIvqk6Fm0hgmXMzmMkygc8Vnxv9eMfSvjeno7S5YqAnQ5FSOA1+nbQ
uy2PbhbBoHC8OEv7GO4CPppdMrPPwFdvG7LJDDXFQX2lBTBogj5Ka9B+uODCdfqh
vpUVnuD+b+VPRtbiM5+2Xa25L1YRpBwjCnTx7pGzzvNuYfj7F+nM4CqJDhkvuEG3
`protect END_PROTECTED
