`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rpsbleh6DXH5k0Y8WiA751RSUQOMO+paXc4rLl5TLyxvcNl6iPz3HJEMAujJS+iN
xJ7kCOCECONfIBCNNvXcImD5nElyGj42qBQcbAgd3QmHALQq9cBj6Xa/2o4oLQ6X
LMktnQ6eCnxvRzOA14CFmqefQSZyokeHWe/QwyWnO4wrWIQvBAZ1548HMJe3dUal
uLyr3J2IZNcleBJZVn+UBSzE3jDpBIzP2N4OoC//isy+eMMZ8Byu5eORP4dCnXnx
v95QsehFIFcHcZBqiNWLY72PeNi3+oDxPiN8ZRDOci58A6hIBp9S9w83z+SRvIXn
7khEK77kEBAVFvKJ9TcP6mk9F7acmSAKaJmaXrd85XbjvQq4mkCwTIE+zXYY373H
C7WQp93NjfMFd2r/301rKRZRpweo/wA/U1ZHiZMuQuj9ia3JmFXnQb0DmmtVwJ3s
Ra4b1jJ8/UDH7wf+1DdzR6tvUOc1NWR+2YreeQvuvDQ=
`protect END_PROTECTED
