`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUB1G0cpW1C36LYz+CAt4H4yUpX0MUlIba3VLD7r63vV7q8aSFspCcM8JzcEkSEq
jDPrQz3/MiALlqX8c6Siybl1MV/IFcldPxTlGeRqmNNLGH2I1ErghPgnvenwYk0v
t5JfJoNmfNwaWSeoL1YIzT3w37F/eXqHamihmTkzIPfy9876MFmiQPWVq7SOYnSz
ZwsDVj7OuW6M36X8e2sAuHjcZKyMtXmiJB/qQMtVTZLNqM33rI7C8fyv1IIYJorK
YKUQgaw0mipNyE348gKcrmyoVDO8mBW0L6LR5670ySfAUFKiDrvN2Dl8vuFj3hUc
jgqfyO86c9RiVOVQVXOUoSSGKoNJy3eeDxbVw/VcMJlcoGr6TTxCk4GoBLnxcLin
HVo5riBlNluS6P1mfZ2wfaADoSaEDHWwKulAcHxZ06o=
`protect END_PROTECTED
