`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3mytfr3Go84a34jdbF+uTO0mh3VYwOOQAxTQMGR2nituRp909K4qDs+TVvFtT/I
qrv1pngEHLhoL95XTKhH3BnqpeuylLoNOeR3K7cO+ZAjyzRltO1ztRxZzTmm526C
WnFA7AWi3WPk5LZ6UoQY20rBOslJYWmJmeWhFXPSF+x9wn+iRJXMh0xjba22bMqf
nkNb7gMupTz2xOt9ErDe9gYbHx422p5ClI79nIJVDsys8HaTbWd82Lnv7TqKI4qc
QnE3qhdAbU3U5fo2+VuBV0He9HKVl8CZyQJfNDRbPhGLQys6S+/uusBQke8+zeHt
X+XBTTQZdMKwNfAntassYb11RJuljl8Qu7PvLcXvC8lTB82Z8FZFL/L/8GS7cA6d
iO1RQPk647C1/wLlxMcGv2ueMq7R6v4o/xGPbCh3BEJKiTJRmmcRCJI6Fk7ix3rv
dfuxs/Dk4xA3XkpR+vyfwjGuyBaWLHTKlZt8XXoh3oYQYxRdiMAEv6ubRDuLD1p7
Uw+zkMivFw0PpkDj8yCCycqaRHKoAymh6mKruWOG1nRnzqageXGStFiDKPtQjb6O
m52KbMfYV9e8xc43HXQ3GTxTCvfVrVr6MOid0icn5BOG79okR56HAs/DPrLFHNJ+
+bhJjjRTj8fjCZvdoDE6LHXYJEBo8efsUA5oK7wRgmjC8ymOdk+EM19sA1Er/jU0
`protect END_PROTECTED
