`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEwUHOx1vN5Llf3ngDD4MUsDkGVsfmO2NQ11RV6Es2wAR1tPBwl+bcQdcnhkfAt9
EMe0T+jbwoIPAAVQFKenoJvCmzNcLRwc6ApyYFbCfIl/W3Wk1pXABU5cfIY1gSZk
qXJKwLIpT+AWjHhFQHcP4gtTENg97PSx2JAyu/25wu7rPTDp5ktff53WZqV7t6QA
pqDVIyg12zli1OshnD5yHNz0Ynf38vs/AGFsxOZV2EFDO8JT9TI3WqQJsFny4FI9
Co7DnIldXGBGzSsBJey+l/VNwYf93VVtaUn8vBxpUEuDNST8v5qvAJxP2oo5NUr7
bnJZZvvaQmLqGd8Hqp0Vc8MiBvx4I8qpzy/GlMb8trD2K8R9iBOKUUPzxBAdcUbs
sps6fl9qqiU0lMBkaJQ9CG4mhXvOlbJh/POpha7tB4HPdyWpMqy1j3VrgiPoTk/Z
ITznTYaOMXnfmcGuOH2pDRSPGc61EgUmmmSVR+FaGh+cpljKkAawD328vLYWeI+i
9de/VzNKTyRF0atJ/A0Nhpj29+AqbTFBO/mCWNoN1rM=
`protect END_PROTECTED
