`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n49XDxmmjWPi8bFg5sHOBwulXPnmhDk8wzTZ60NFGUoSxTTQGNSW5ucjQ4FqVdZL
Fb+i7ERfZsFLeS/gQtPQ+5i31Ykn9NgTTtaB/jkI7SOSGoAWrrA4ngRfvo/G+FTq
Kl1vs4090Eq0rSVWqnZRg4DrOkWLihvxpexoeI2UARQipEdCVDblTkufeiR2nl5U
nCfE6SmmgVIkyHGRZR+CUSOekhboq42CZ3EokL64ZADQ9yh2n34kX/OkXRIyyn8m
iap03jMnsPJtpXSdzVeLm511oHY1LN2gxjreK7Z0b4dmb1jP6UWcBD8D8mEtigni
5UxIzIBuuPcZ/ah9eR32728AIqGRL0bGyHByiYNe9A/9E/BgGQgd3M0rlCPj1e4R
M67xm6hyedwZdsCJwriafF+RGrdVfwPD2dhJ7qcPI4onQnNNZpE7zPjEVs0oVlbf
RISAxQliLkjfo1mjQAHqb3nL1HhHWfaqMSkVNsXUpBakPs3FTgbCjJNCs5Cviy2j
tClWfok2vOqBhIcNgId8nUgNLAGp5auQWz1vQnZYtbimosFz2PHdKNmhuxSPCFvc
EmQwf2xS1oQ2AiWl/bt/FJFg3lmK6Kbc2CWN4dMkjWU=
`protect END_PROTECTED
