`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7a5v7xDzNzj3fu2fZbGgyMtwlObydCxjLyRIR5YBGxrPgvK+HfvO6JyfXAv0iGQ
cNYidP5Cb/r0oNisrYF/jjcy9h3JbTeA3ItAyRdIFgXTrBf6A1dQcKqbpIr3Y277
vDzFKIauZwqaQvK+8/bsbrUsm79X00//loui1su9VlSNeqRSbg9wmfrag4X6N3ty
sRpiliam/7M2a9pR73kZDoOI6EtnxuZYa5jvLqWtw1Oe9poH0GrnnKDBqjTSwX30
Z5NmVdnVef+fCxrsrPo1nr7K22c35NllYSjhY1ensJA6FxSblNgwYpUwxUxNs//g
a6Th9uSIWTsfI6yIT24yA6Vsg9fdNttVR391U5+Og/GlMe8g8IPIzF7zwjPuj/vx
xDxwPrq5gUH1Fey8kcJC6Dd6JvTUFtv7C0u+IFaQEI6OYLwQouNrWDNNMmZrALTh
j6zpKhUDvjGT5hRXM7fVug==
`protect END_PROTECTED
