`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGoo3yve60vyNn+0gXYbFDjFllucXKHDRf1LjugF1q8QKonsbfvqV6/VWchMkQZU
jtJNsQf5aZ1tJpQIlIG4I8tY+2qmKxllGlh77Wh693zOzEwC6qg7rPH20smKmeYm
y8lfvC1gG8L5AXR8fEMCyPwbm5AUgdHU+dgBXKh5RvyAdjVNRXS+17K5gdpWu0Eq
OBddvIRFKaK/MJrASRvDDyyvJqwH5GoQ4bf9B9F/OIE34AdlFYK21MRCmskmbLhI
+kUEja8+gRQzjvMR1VAtU/pffqenqwbSwJ5RroohI9XQMSW3C+Ou6em1kJqTXh1j
e8pxwaCjnl9oH/1WJ5ch7MXz9lDn4HU4coFp80VHxzIyFUnOsioECtolNEBFBo16
ZJuvtF8+LeMtJBnqYwHoTJwK6uG6iBI6hAJtdt29IUHGa29jpUk3Z1g7jJpl47HI
8IV3YG+gpBC2kTqveKxgEYjcgrKYGWXNT3KXZ1YMXaGKz7EAb7E+pjJZ8Pj+orVt
eWxiPlbPA/Ru/edFRfUngC2zEUPKnaetX686TUHTnZlvQiVlVjvrCaEWABORTazw
DSruzOO1G72gisHoNu9Bhbz1U0C6BgjVZ3OTC0cx7A6X3Eb3ZAm7G7t3Gpck0iwa
qQBjScV1ntgfMpq/qF2ZJ5xwWvJt6O9b99nVhoI0clkVVuV8+MucgIZsjKKXeagD
m/ETUYYMArL/+rCZ5CzZ86xE3E8e/k4DhCIFkwbcrEU=
`protect END_PROTECTED
