`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4lb03GswumwlOBd+481QfcZy9m0rt77oOZIn1JYKJY8ZWIIDKujC5odkE6QHELg
SQEjPADz15XHTYOELR2l4725qg3CPDoopWu9SWpw9jg8EQ7v48UcXPLs2HQoTII4
4/tRIpZqOypTSJxa1D6X+pNeAaEyoTCCNws1uAEnPLP3PMWmOa/3hZBXeCT3wdua
JH6oMB7/U6y+UhBSsBjZq0UDoRKLW7nXBaIIVUsE30K+vIDUxG+7M/d8r0iedEUV
/tQ3/Lg3nbuOPFoC4rcVdz5VbX5ks16UOGIzblI3pSWMOh7K/CPSuVKN0wXfa/Fc
hx7eeBPcLIxSmQC4fMUKJb/xZWhLCs7IWq3cMz3V0UmTr9+5TWt9iwGajjjlAZ2c
d39143PmblmSFbZQv7By0mOOJyNLmk4uoFRezQuN2nt+Q3b3C57wlUVwTwFyvW61
sxAMUv9xPDPIjs8lJQIZR9teBkk2q3P4vLPj7zaxbiL21fUThzNwh83RXABGUTxl
ZD63VqarP8VBOQNsTKrYLnWIE/MOn8zvID6ooV49SjJYW5b8GBN+kMSHpG25X6Yk
8vudRRfhofinao7RbQvBXpwYWa91RfJZdwk4+Ip/oMHBKcBpOe/cRSE42iGWn0AM
h3gqkVfUUUyw+WPTxuGDR8vNHRN5ID+Y0u117coXWeA=
`protect END_PROTECTED
