`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+nBFZQWXvJMflfAu3nV61ICRrUnXckGjvLAUjpVFmOvzOMsf6FQqm6aXAOvAdLm
t8v/Idn0bLtCaIvCUzVV/iPftQ+D9vBrhmSPyQ6/1KDQD76R40qPfVP7K6M/tzvT
XoIxepjoRwyGSzXXuGG3SKQlsDwGapRnm0OXNgu9voZxwRD3k9t5SAW8ohYuCuy2
/ySVKWq/LsCp8zx7ojfcR0O8vnR+DEGmK/21s9WuDL/Y6mn0WoIq236o0DdImLCa
m6JdTrwaF9zLV/4VTwtuZ87nzSxNmFBzAGpZhYjfQcVQ0qz8U5ORb57Qylbqhxgq
81/DOLtHD4/BGXJveKWtM4wTIM0WVhEg0YTvytenS4KU1FsPdLR/PYG8surjbNcO
K3+m7bhieB7YlnMUO4tUEGLusOY2Wbjxk3C0DKtxM0/Ca36AztNKjtW+A7Mu7e7o
MPKxpYP+OujPnr0jxNoAQYJJMsQ72FMIDXR9CgwcezQ09aOcGx6InHt+/c4RplkE
`protect END_PROTECTED
