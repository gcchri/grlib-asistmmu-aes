`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vy8H32fXyyohPaI5FWt+D5LRob7VV4FWjpyU4CunqY9Ynbpm53aXCMdJ+ZxIUe85
7nwP9hm0MyWLX3NMpzLIB9IL9ri88RUqxJ6WspOCxTdIgln/4S+Rf3LoKwUY1WP1
yTVfjCSGnlK3/uxei4R51JMllu/farZyVMtuCYP17viKh5rtFCVLu+Pwu1XYoNB0
2jI0IyyywYKg9ODG9HjlrbksIxpYpJVBsNitUMDM+N/lXawQSAcYlw1KVKWfteta
2ymTWDK3/2/mU/7K+cL44aOrLx1RhEn+UzVhuNC1NRkkrcXPOms0MTrTuKJIV7rl
6E/nlmM/p4d6Ez6+fP8QLlsgO4I5H/jewmmV9nYpgXiftx+GbFFYPA4U+8vqcZP/
PuT99NfZkI3BDtnLF//OO5LuZwsHgX1k7ljYnOXg4R1byYzpACx8YTr4odbYDqP8
fwjo3fn7s/mNroeYlGiTMsufP5xZCa1yWd2v7uxbxGE=
`protect END_PROTECTED
