`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eH9FFRkv0yt8x5WCQ7iJj+Fw4Bb/F7Sk+Bd3rXAvMmTyoKXvWw9bMQQE2PQK4OA5
8eCGz9peWr3lmXYJCRrNtEl8e704TOpI6zSqhhZz/EG/h7kgJ3rRjzWhfLXzHdxP
6nW2czEH15YhWNfKdgjaxw5xDFTfX1jyLO6R2B3IsU3adlfzc7x+HeOJ8W0whWoS
FUJDEKNGMO/viE1uXnLiWfyUtT2OLrFSWjrfZXw9GFwbt9LA0e/tfwti9FFrsIg2
5rkzEl/0dlDBGO2mi8vqso5khA9YFRin4DgEeaVz/5WJHZo980EhQU/9lW+jq04P
6CMS0PO3+WFcOpEVcTEwNV5nBMdnSLsP0pR4hjB/OEdIhVRPpaQA5iOr63f0N1m3
HQoaMF6u15MCmCC3/1i6k0hWvSVQevu39EVlKvmz7eruqflkPyKS2SNK9jCBI3Ej
C0NStLDZgFHrMy4yEiw2vj8Sx0N2V+mf1u2ij7phxOACf13qLkjNyY8K6/Rgs//Z
vWRWa2PFmX3sqTZy/vpvZLf15vHHF7qxchvOpCZ6g9NJo6aZ6Q5d7Gf6xvXaBJQl
VpwR4eTcIjP+mkKNDPm182TblDvWElgbC+KndFMwWSEdeHC31TSCc0Uw+G+rKchz
gEbEbgsJPi588r+qFiBtCA==
`protect END_PROTECTED
