`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKXxfvs5NRAIfpPc3fM72SbI0q0D8YTYXcrzyqsXHf+ChkBXq91m6UodW1gz8Vzw
UF8HaD3gyzPmVvAuzuRZ3GudOU95xUPnfJ2VdrklcBgv7IoSLFx9+djD/+sM9hrX
ya164soxGUEpC+uw/pOzJKMaA28WctiirKkECb2Z1qLrb60pT5HcHsoUMOL02SwU
TO1OBx3w7SR7Y8hVm3L/4lZhor3nm5hXkzG4nQou7C8bTSXdS+m6bvOE3whXZHxD
RXH+ffTWkJKZhK2aJOCOVNsRn/ehgEAR8MYyFzzhoqNGj9cgfSfnhIcMoqfdP6gt
`protect END_PROTECTED
