`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cfW9WSWfqg2RXF2U8SalMWAMqz4ev6N9GtWT00Ku4An+VUZLBmlFRvxyCacs0vUU
EveywZO159JeOX0MsYrwUWqzZCzVhEDCcqaXV0Muiq+zJwDf2C3rxPZwBwyatCX5
pz/28aolEW+5oMuzj7DlebnqNLIG7VPoDhxclq2g5ppijJrg3VDVzmcbRwOEVg7C
7uDcjGSnaS6lsWSmB3oUDC4hG/Ny8TqPHm2DcEyd+2HW6Zod8LDPm3UEvuuKe7lF
nOn1gQG3PaixzpPUj3rTvbkuZoPeHLiS/WTdXqgzFivu94XVInGgL/O2dbOa6gHF
Sxe91lDy5Kcyf9GI10vspMDuL+rjirz+8BVWsL82i03VS35dS2Dr7OANFBfz+EIp
CUUiXfPJmBL5JwJLNJZkS1kWax2ak1ieEP8zlHgNNbvbhgI4eQof6Tv6laRDWMf5
Rd/LN2vrv1tGjmM7T/GdMYSIwkumUAG1AM+a6VVCZy6B2/RSMS9c4VHaag4AY7gF
`protect END_PROTECTED
