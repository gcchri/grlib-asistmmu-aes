`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hmy/rDwdb5+G2F/Yo9fysvRfYigd12qFp1bvoeOYEr1NhonAnfkTrt7yXcNHBxAf
PQ9tNqn+BTLP4XDKP0EPA2Rjk15ix2/rrHQNQP3TKRFscU0l3vx237P175wX98oN
T5ybaecIvwZvPrlA4obdVo/K3nUoXdz5viAmnAzu34KbMX7ZeN19oSvQaSHH7TVH
Z04Y3WRaqNLy4JCtziqEMIJd6UPSeA/0Ph5UtrfIxtty1IUlY/3Qo1STKGgWkAR7
Hu6Bpe6Pn2FUDoftFS3KIyzrruGmb3ZQ/0TF6EUq9ks9kQVwI8dQo/9VQNY7KlRl
clt9O6xYxvRGZt8s8yMwNNZsyfYMIqEsdLPzkfP+LVth6mY4h3ai4z6cn1CaDKDT
xwCKOE/hi1mbJvN4r5hl6oZTOof8oCiHewZ6xsCykAha5vPxNsediFL7dqrZ/tlB
hULAqhP/sWy5rolxBwbSEqmJ9tnZF0F9GlG6FDKhHRCDys1OEJUGuyulSqLFSrEw
ogsP/AEju9zzrnP/SH0ob526OmwJDrgw+qSNzQJcylMKbw96qvBEwqMzpCcx5kUE
Pi8NOxtSionM4R/PXCNfuAu3mpf5qJlpn4KXvdl3aDjMBmQk6u8Z0KAnIt/rVz7j
H/Rs1/EtKFxuUO7q3wIsTCzBQ/NaDKbq98zx2YdBEoftE7Exj9OzEVOzPlPrEpvT
hml1x7nNcvDicbl6+2gLjrvaA6UNrDgCJMNj3t2m5vtfrzELgpdwMW5Gksygu0+T
c6o0v149NgfVNwHNyUp5Gw==
`protect END_PROTECTED
