`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2UTwLtxQm07Qxx0jtZOtguSBrRrugk0UCruiz2tug4YJqZKy1o90/QalpU9FjQR
gRGqszpOm/HP7ubpOMZpUUdBdn5MVUMPFm3EppYEr8i4k2xLLd3wwFRc4Lt/Hw53
fjmWYZS5P0k1+IUFyypKkwD5dfHCUZO3vQE6zh+usmPZZBRqzixF1iWaQ1VaTOIj
qjS5UyZQjHi9NFhOGy3V2SllI0kPrU8eDqoWuDLWzbEN26furRDUNA04GE0g57C8
oTVaOLCz/0KWtXZ3X3DP/g==
`protect END_PROTECTED
