`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nMZWt63fezkzms3BP94miJyT2XSlfpUhwEh4kh+5qBK+4TXQYxX05h+PEDNUWSIY
xAtkXRpJlE4JpdyLeOXn5Cx26ujSN94BGg+L+3Gs/k9g17d6O/6DZbRccsjswrPf
POPMVYaS39EK6kUUsUZiLuox2H8NjR8sUMkEePAoWY6sKuXMd3gNyt49rN7Jl1cL
xL9rE6dBHqUsUNsvN4gU45cKH2HviF6HC5auX6K0SGULkex3doEXx64jtZ2Dsnz9
R34VoxlvkOw/ybBeLsbBNuxiFxat9kO7AatkOH73XUNk1xdROTBd5DkS/4ekPI78
uCKa/sBDupa9XP1Q10Zrig1U80KeSYG6NtMo08N5SYqK0dqSVD+/fzLRtvyxF2xf
6D5NWWyaUgGuHn9pEUsbjQq2VJVa7xHWNHIxYNUgrfTgVRKQFGicpEuKTJfuQAyy
8pp15yW/vfbw1KgdGiGkcvyCoEosypxae6ddbcA7XsAY1UuiCtnexwiBQkzGiQBK
pFb1qC2mdHmShnqhoJiEnRxDKjW0u+IoOvgoL+LYbf6p6IPIQpfklk20Jn5OnbLD
0/R1BJtbfKRYnv6oRm8cbH37E48jbrBCphGJm4ns4NXZjfE4FmYvPVSXOmX6SaF7
XaF3bfLT6blvIMLcvfUv8HhUlMBNRFpsWy+kEFVxlBvcvOTa9ja3lvzCrUpn+FWE
G0KFzWYnwO+cfyF+UiOmrCtypxRVLhKh0ZVv3t4TT7UDfeHyGPy2D51DTwBMdRG5
0TgDWsp4kQeF4NhRzLWMASYsVBsbfgUONzv1n6PAwdLrWOE1H6C+9F2h3cJdoNVt
5TumbuS+ga0rrFQy+5nqob3oeOgwe/oBLlzp1Ag78pJ2I29oOd1pebfoC7xvxk5g
4ymuMFI6cDT58APQ1dOFJudxIjmdxNlwzQ/mO18CNHzaHYm7rIjjj5Ohe28nd7zV
0AjfyydwT8sURTegXClVop6iQHnD02yDxEHfx4BCvPZJ7b9zn5VaKWYcMQFSxdUm
W3Z3qAPfJBgIAhn0mIMx+bUN4YohMgo9s+cTMSw43chptvPSQBFAuftJA7EH8mB3
haWC+wBBNS7+Bwln/CsKDb3DXEZbP/1hILz79i2DNbIXEsMqeV3Ye7vd71zrG2fz
9JROqdX040Zd5jo1O5TcekOWAw2wWKv7TU1tmjpprwK9PEaSQRf1v8WwZMBWWlve
fimcLTdxF1VXhu44LsPRuhmuEVzQ3hnqplGEgpiHfsddwZaUuDQaLdyhs5+G9bev
RZ8NZ+4GXF+fVkDPxPqDwbN/2L3OHNm9AVVh2R7tpeq6+A/zFfzSlOrKGAXmio5x
9UdFp3xNySCinHjF1M+RX7vXSwu9Z5F7/Jfsfchc3wg3709QJxghDYxerq3KZ9Cv
Aou2h5DuWWghbjK4lBik9aWcCLPCtpjrs2JUjqCYkFCumbv24f3uwGcO5qTMlukr
GeibNhlzO2AOYG7dZh2tjFMMF13m7GJ5zaBpyvn9rqAwkLncBS8T9eE2BOP5eQ6J
obOS89gpwIzmn3McxUfRN+pBCbaw/MrN+dUn83CVbkxi9BXbToC50gDqx2MA0YtN
uMTWTFPt/nIRXCTVbjPo4KEZ8BBEcwdKuz9YOTe8TyfAYNax+Lg0TcyBR24ElDaI
2Kwz7ja90kjLWnaGO2V5xFqp3alefvSxfRdKHDDV9aC1EVFbwm19CYDsgESZJwO4
tQyPG8F7bCMIqJHXnWrT4ecLtxf5rTa9z0kWy18rO8SBJwDCKOgNX9Dq8GXlTl3y
GJwBB2PWbkWIain8qUu+Ki9v8VO2gkMX1vkQqHpMzxRnAa4HZ39oiaMwqoyjNux1
WWgBUOOMROZSYEEJH5GgTYsDC8iKG8LTU6lPX/suU9llsWEDq7qXg6DhoebBycgL
B55M210jsniJuH/EuZ2a8V9mWaHKc7SWbzQYCZBBQ3M2AaVT2u0aALUL8nvnYBiw
/YXvjGu4+PmHTwW/yN9HXd7I/SWvVgCIvqNeA+S+ThkgnWztzSppegwkuRWuwHDS
saGSpxqctyFCLZvw2B2DrHsJmxKy5u80XIaPyrYg1FJK0y25btaSrmd5+wRExFeX
1oHECqZtZvr3E7CN1E5PcMIJEC09u8N5ZoagYyswrXtXgoyWwiNu4tQsteqS/Xp2
MwTUQv++vW7nj9K455EhTZj2RICk+BhvWEbTSq/0jgQNtQ5Amlb/IQal5c7tqUEP
NhSmd/htwg4NsN4QNm3IPP7Ia/iePIaaUn0k1sDSSFOkHDHxkxHiIoROmcvLHKiQ
3TV/A0+Tah7VlKzschGtXHyrNT6kyg9lEND1j941rl3MyeHSN+rFkDv8rpidDL2U
8XJ4Cylj+t7kGvvdxfDH8rLrRmE9nYMn7YyiZmGIya/2vFaqNBXOH9LhVZd6avmM
dUev2q/+BGLiEvjEVIY62O+ODpxzMjcHK7pqEucQcyjHYUbGV+amie/PoljmIYGV
hW7mISPtXNxxgcLSU7AoSaL9o/hYZ8ZTYjp6A8JN6oRg3+P56tYoOBZf0H99nyvl
yhBO/H5VGFuvAnMJtCwxuyzwthIfg7nw1Fa8wdlT2WjwNKkrrwTeJWr6j6dGYapZ
IjwVhkyOv1rvQBqn+m1krcYpSucgmRPVf7Y6Qs8qzKowqJFzEgAqTV450Cm/7D53
Zlezl+A3LpWX/eGUJAd4VTTwtFB0hFYMihBJRgLPju5QH16k5L+1g0W162g0tr9j
n0+RmUSTg9oMXHqcVwatyS1y9ZWaxcPi3V3p9woZDCvVTQFOle0x5TF6e4lNdaLV
nX0HT5En/tsOQbkR6rT4N6O3wyK9mvNhlyjJhF/fNMJ0R4CL2IEYr47VBOks9sm0
FTc6dlAiaL+UNNPJgJ2hT93wvB8Pc5JTQS0b+tkKqoKCccjxcw26D5quoZ6CLKga
jA5Tlpm4+Qj51G2ls/eTnQ4sBSn4SKPelagzs4KO/olnp7o55g6vwFASl0CYC8HY
nb4eWUOk7axYkq+GynLi4CxMB78qpP690mg1aRqo1hYig8hCdTggXBCQ9HDgkpcb
ECpgMcykr1YBkQGLbZLNbxwJN7mJUV4p2nsRxbh2x2x4iEzusnQPIRzKmIo51uSn
c6LcQB6ZcGjr2scUeD6GhDavURcjk4tVteQHPFq24mGgl9+BLm3kz5RlZTRVWjqG
H64jmGdmsNh9dkQCJlsVxaaWz5/8u9lP2uZXMrxf9pTqgWCF82VV0eCwp6aVmfVS
EGoIZtKt3GtmF8y0jPD6EbD3AyV9CtcAz/8CUUwKvUV5IGoKWeuNTyjUIZp2F44K
prf6IL9S+OXwRrEldZtBmD8ra9hI0YiefIGxiGEFKAJ4bvkcXrCKpiKhwKOvA1D0
3QWA2st/XAPj9tkxokGX7RO1bU1ClTTlc4dOGy3SLmLokdLHg6MHNC0bKHP9MK/c
YXutYU2+LqdS67tflgGfTEuAPHb5a8eN1U4hhmuwq8w2BV2fLtytTuDhs0kYpQGb
GYhG0+m0mkkXNxQf9w2geryc2UXho1eQmQjrJ73DVzbDUXjnxZO9zju8q/cvFcjn
0XYIAXZ156A/fLwkYiVRa/D6p/SY7bNAKGNI+Xw7Fqf58dfoHVSUz/wHFE8j3qIo
+Kz+vtp8nh7+/dJaUK8ozCZCy9KP/NS8Kdxa89Rm2x8euawMSOgd7prgW1iiNFC5
Oc6e5j7ASg3xET3lq7N2lTBJ42n+SklvqdpAnSbE5EMvW1U07mrAcRPmHxVJ3wzT
4q8+KS4zbNI8FZ+gV7AdRYpMVcDlQ+KaejVMVFSJdmtOG++zWLe6U9qrwbAlY0Ty
uypJfvNLJQGAJPpQpwNtphR6yY715IPfthAyWpibyzbTppsdTax23Ee2PyPRMc2h
5170qd3qhQI1CtuZWiqHZPAhUlIB//5UdaG+Z01NtMnk/zQwt9KdoCvY8j4tfEGQ
8Jjm7D8YYVjr1z4bqHLiZJIHRvxvnGqNTvMvXwOlWox28jJUzXMwwiWtl1RIE6oQ
GGGG181P/zNydciULWs3GqeQSOggdX1ye1yIPAH7mpiui+dWMYWLy+SZufq8+IiH
6RQPtwd+/rZAAcP9cel2Lt//ijFzxjsd03QGf06GGIh245bBjb+Vx33ncZbygCgO
rKQEQjVMm5/eBvsigTghGL6C8Xds8UmOgROmkg+astZ1fNtFSEv/FRRRPRGbOMly
5/GKubTcnHitwH73wN3XLAgG953+CFEEi5Vxxzm225mWe0dkVp9Oqa/wS4nZIeeZ
he0AVeALZoVRrtgrVZy0lw==
`protect END_PROTECTED
