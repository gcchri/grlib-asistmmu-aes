`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
excw+j6CtRDggpdgoVBGvfSdebBsGuTh5N1L68xeoTACapEdrZUcCP8CcnwzPTrn
XAbNlwytqCM9EB6NJoLR/zLAvFw34prrz8jIdedKt/cyNFPzFpUczq4AMaVl2jnB
D+4QYhOck3K9vUk8EfdF729ppsHsRl6URFSK4deMdyp6UvYYTbY9LG+7rssraRLr
rxV9jlDq5uQl3KrXJ0zsY8g7la1JGI5K5qSwpVMNOXphwpMtcCSPwM3rLP3kaKGo
64cj/QoQ6917yVpAGtWiZGFmQ3EVRAOh1lgWu65TY7B7iU1PTl9AAIqB4bN4OkVM
hXvS5lNegDu0XP6aaGKEP+/fd/pdqhRrQszhinHaIi2KLWuTpH1Pl1iWVvYbgLmF
lEN6owj4iNTwKVUHJVhRlSLtVM2subsrp/iUCG8jVVjw1MbZUqGRvB4qVdz/B1S6
EHbfgo5LRGvp1TWWg3oFtpUw3qed02zushuUNyhpXCv4oXdA64Dm7PvFZkB8/d+h
DIOr6WCPcEL/l3OhJqe+s1Z03daZTIFvJ3doDYqJZBTfhbNJEJ10dPR3Qbz7ajkt
XoGgxPratV4jp4n4kxTU+hv2kY96hXnv0u0VQnvUstnS8qtkyh9fZ0NVBT2zHZ8l
wJUF/LrOwsx6Ao1JR6TZDNa0W3Ibr9BhEFDa44YWpVnPofqWm05mijIre7COf5P4
dOmEaqD7yTU2pVPy144h+s5K6EoXfsp1SjJkHIGaoPXkzmmDl9c3zfI5AiULvuC9
9pCgXwWGhY5nWUm3qqke4g==
`protect END_PROTECTED
