`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4eEVMUg/Xr6et5J7yz58eMVLAfV3ItsH0p8JarW1iey3IzWjoZZYyNxUsLuEbxmV
OqwSLC1p0A02VJ8gwiyvQyd8DYiZ/vmjOEnVajSB7lYr0uRAE0f8zx4Ppr1h0Jbq
foOzIaaAxs29sBPt5pCIPE3/r3RwJF0okvUaUCUqSgIVdtERz4Zw+Zj7JD2QJAiw
Uei5VO7qmT3k0f4/WymzSxXKG0HCL6Ulk/cWKQ9MklffZb5RJmUbZjijxab0SAYj
0k7OH87voeybS90FM06UOAeeqZZSSMaYSnd9US479NDloM+8qaUlN/E9CPXLg+Wc
ao12CyFSdzpruzUdQC2UN/ahKlh7fQ8tUYd7/t9I16/OwnW7xTfxYZgWzjUMt6Zj
HwWz7XLqTU6jIkSXeMARQ1FAVzMQ4CuuegIz+4reM6zDlZ/FHHEsHr8FCTe6MRB+
aJ/fXi3D06g2hbdpkvaLhXIUw1pjwVxE4uBjLvLJvP2t7QQTYB0uTb+S+USEhEwL
FOZu6GgRnpEb/P6fDDEVbb/iMa2uBC9SYX7cdd8Yyu9NkDDoGIRrIGERBYmAM1a/
jgnxXkPoCn82P7Iia3fjFw==
`protect END_PROTECTED
