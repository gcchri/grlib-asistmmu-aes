`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
acJ2sY40UFuRQMO+8NaGC0FFSFjhxIumtuwwGYtpFkCfOh1xKKG5PfzcyzuFSjHk
OFd/s9ZFTDqBp+rUMsAmB/Kj6m+mgjDD9H7vujLCgmY9PsxUv4IzoApUFvNewRUw
QrZqK/pBCogqH1hBES4F6fAM78gwTIh3e2hNAIgLQUrr6s8vWc7DBWI9bOHiIPVC
9wQUesbfWm0l639smXbUriuNywtsP2EhU8DfFQUuNdBRzwfCZdb/CP9EvcTWpXC2
BuYuBHPFyyOdypmThr0H9+TcCg9Y0XCLiWpKFNL3IG88DdQfJnVL27eGIFKZsbMd
K9LV8etJkWyOYp1vgWPHjjhCvYTpO8N/ldHfFED+2/YDyrs3vuQErM38zcwn3YGY
2AI4f+jwoSIYGQxLpVyx0+6mHOYkNazWKpIU/QjTBN2eMoJGVDwIBKGPcLzjfk6A
mnx54KetWB/2jQ7Bs1cMwAepjcrdxAkX0UegWsMnlh2lzfET5HiqDNwOHPKwBl2S
1Uh3Do9f+t5Ds3pONW0S7ZqOZ58sCCUW/Rurf2KzoqQSm3SRD+y4ILY8z6Hb1tn4
WzUKjnmt1JycMucGae+XGOr6x+Ml8z/Dq6gRmKtuJM8RpJMuDOO5xwd/mpJ0NXqi
f14i1s/t/8KLYFAdb2NThabMgfuxufGFCcv0QmEqHBCmMrCcRzjoZ53R3KrJSro7
ZHGER3Yq2wnQzRak4irnSPL93iC8vV78eVR4gY3hgWFLMZKLj9lDRvr6JGoPOYo/
//hFdg80nitUZGZE1u1RMw==
`protect END_PROTECTED
