`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9P9os91g4dF4h826FWHWFj9u1AAWvHheNyaHt22O+1XtF9BJo0cmxlYFhcYVAo7w
Fhng77TMezp2Gz2FnrXYwU+UtCGjMsPrL3pHwE3p/EP63ypeVsri7Jnfc4pAaQ0t
/LZMvcZJj+XMfHq1WX9ozcaqB2+lik8+VRG7/wFZyQ+cIWO+BfH1MiCU2NxyNAfo
Mh6MGk6QOvp4RAMs68cmP2bjsoHzXS5MAbHlLCiwXWWs37ttCu82zHfg53SIDsgJ
h4OdVHInVdECKJsyvvkNQdrnM0r8AjAQpXQ/TJU8zg/uBt3Yasj4DzQOd2cZvTkA
yGjzhEDwYi9OgHWql68UB627XcNympy6aRo26KFYVc0tRjezw0BUQKFvOaILf1To
2g+vT0Z+EHzff16v8qlF4NeNLRumek8wU5yfNpTOb78=
`protect END_PROTECTED
