`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jNw4fx0mNgD79msgqyXk2wVtyWJT/DCuSkiLFiKRJdGM0TiamUJ7nmPBb7/V82+p
wQWsMipm+E+CgZFR0v5o8TZqRIDzR8M468unHpZjMvXPaMGt/7a/QJLYS1MpDzqd
kF0ONJ0Oi+a0kWFyrdz6BrnoenBIt0LcF69wt0N2xN5Z/vtJF7cdVmN30JjBRb+N
3V/CiSOsVQ08PCefj3F1XWHuPKNMPec4BrwzfEEr9ErsP/jpwD2yJvBAGEK4rVqO
xWEdUtyth933YLS6GM0rT3Q4fWTOT5e99CLDdICfgCKpWdFrejbAiwS0bqkZfAih
P1vIatGjBjhAJ2dee+XYPgzK1r/sSJ0if83EVUw1nqxX1mWeF/+Ra4Cd83v2rIfW
C77t8Ft1CwYL4VGbdvhFqE3BzlyV3BBaqm9HkmD7BZwZBgvTkUKA4ydwlZORP083
ahbv52fHDUtawjWQ+WPA5NWUPPMGuFNRX8rxC24NDyBA7QthcdfcDSldFP9YiEWr
`protect END_PROTECTED
