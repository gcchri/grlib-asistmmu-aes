`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+fJ5U2loEi+Ip8eBS2I42hdcocLYOSzRQX3JvtVKQlIMBLULRaOoSi5vW/mH2+e
iJgakU6iovNbLb8XxnKBBwju/tIWH8HYtiC1kL69SR+XHImNuFXc6BFXy8dUNZDJ
fiyudZkZonmaoIkfSAdiX4sf+IKhV6wfdsn6gRDXdUzCOeLSKZyv2Lf0GxQ/d4vV
aRmXk9MtMXP7d3YVR+fov81/7nV5kvPxkBJQ2obF391cYfsiAhOyJsIaGady0zd2
bjWvxCaG4qF57X6hKEaj7BzY06GcmZPKv6E5qsFvsZwSsbb3ytPvzDQyusuKU6Lg
JlFQHIm2vPQxqbSv8ygPsOIk9uOFGiVUMA+Dqiv7g2P2zUrN4baGT1gSIngqZ0lE
htGTz8GEpBFmhkJv5AKfWsMuPii3ahZzuEBPkb8t+/746OMPS7aiLP7AK86erKWj
jRf4I8B5zZm1ZNPEbpQQ1Q==
`protect END_PROTECTED
