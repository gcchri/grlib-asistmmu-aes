`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
syi50VS17JUMd7Cmcy+UN5RP6NrX01SvWEucVBGTPPVlqfPJH96/6AvH4s+B8vu6
O4ProJfbcd0PS4Kq6RKEDVD5QbTA3b9F00GhQA8YFjBYCVaTOJ+C2klO81LZIePx
XmvAS6Ag01xzrRWqgHS/JW1/RmZC4xEPqQSOQCjzExEegQt+y9gPAY46gbXRGKH9
vozJuZOT3N1wVxWRexJiOks7Qh9bFNi/sFGv01RNG4/sNlXCZyNFtvCTNDb/p9Pp
KyExWL1gqPUCMc+BMJJcmHiu+U0mLXu0+3OqfeNnnNh7+/PDo43w8Wp++Epu9LN8
LlZ+doCfsCp0UNxXN14c0b48D5cHz1LHA2rLbxUHEBOH0slvMPcTnGsJhXPRQJoo
ViPlU4z+S682N2lZwzwtKDSyZTClcm/BovCu3r2A8MiUZ1hq7EUsxwcrazOdsDvO
8tha3CkEOf724TQD7i79F1mAcfLm8kVxkM8FbjuY4t25gHQ22ux66UpYda9O71GS
8bNZMWBWIi5CQ9mgVDLUaIn9crqmGermhQUHld3sK8DZ9eA0OaE0vXyKAlPMIQG3
YbQDr/DzfIydySa2Ei2rHaUFqva6yb8lBkNrEsqLq8fXHtfisZrXU4zjBHmVxeqT
Ylbi7NfxsSY5DxWKi5/LH9EaSfdiOnhXNMcVqQDUxN2Du3X6b3CfaBA2WrYzG6pc
OFl1jr4a9/pzdZLOvfgk3fAawLhsKmKL2PrSGxqPJMLJ1sVrq43OzEgsctVWpE+2
FsR5An5pU6lTgsKnMwnklD5/cEhX970TgqPRgmrlTywIaeznCELY04Dn9zEO+hi2
3WVXr3LKiqmpXuLHvFSEOE4oLBinG+2H64y+Z52NJ2b++wYPx+hDe7h8/ORTzRGN
4xir+Th8bXXu36zpOmwpb2uKIO7gjr0BMYU/4XP/hqyOjvlXAFIWjV4Lb2Dxv0Ow
pOfcuu87JNOoHprbFaVAF5o5CPzUORGFnGrLtPJ6Xe2EZ6TwWlXFW3JsPpRYzN1N
Nm6GEIvft5UvrjhWKwPYOL4DEwCvddXmNaLoz6Ua7FnfufKKSQ6h1rdgHfKZehGy
CpsRZp9UJH8qgzADoJFH5v6rI2TxaQPCm8nq/hanXAVxyJxMI7+Iv1w1IgfLXQvd
/TQ3L+VdKfmVJ64V9IIr4eZwqbc8+h4xXX21krZSFcZ4wSGRQdIiOUxuirwkSe2u
WTmVG6Etn2fuIe44zqVqjA==
`protect END_PROTECTED
