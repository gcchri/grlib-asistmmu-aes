`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kpf8iapxs0quxZuipxbq74DeU6S3FJ9h7dwcZObS/OfPMPt+71JQ1zqIjnIbHOHz
Y9hkbEbbYcXXJ2URj7w64KC1q+UvzhzZVgscRn5rhbNQhvh+Qckqt2XgR9idp76B
sSwMUTrOQi9KkMgBthpdogEOuRe/aPM0G6Y6bxKtlZIVwqKtWWRueGwJGVR3FTYy
3S7P+dIAU+Xg7nKcyY1T5VG107p5oPykn+WQpe108DYajQVs5l8NkFH7yfgtINte
1sBpRHK7QNxZ+b7Y8Qk6YvIKEmZUy3018NN5kfAcKRE0cBjclVYe3MGb0SGH9gkr
ftTDoV1MRXWZZlIOm6zy8iUsI4g4h4/mgGfNulMiJKiVWAg5TjW3huWKUdSG1SCQ
sZqt+qN+LVbq/bchbJmSb3WJju9jpSeMk/JaE1WfdfxfZaVMSmT1TdE09UoHY7tp
/bbqis7HzluDQFqH98GuFHC6SUaLIhuVNaup6TBdFhIBiUBtdGU1lUcqdawFvl8Y
wnA+F2bG9jUxsqkGH/hmvXxR3s6VI82w5PGomfUutcE=
`protect END_PROTECTED
