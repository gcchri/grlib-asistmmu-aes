`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j8vZEAnHqzd2MbxDniqX5h0d02fAPYHnKm/qFSGrQtpG/QWh6KxnVGuThYZUcSBr
SfZCr8UDVsfGxjgTbqOc6UPJAxK8/SyLxBu7HTD39TqhYLpGTrq/WH/NjsU7cUvO
16sDKYvbCwc1EeYB1VP/ZuHri0D/hBETat7rX1LQ49DHXaBZe32eWYgcCRdUx7wB
8NWuJuX9lvqqgBqN55shkR0HrDKYPt7YsD+a3OlxsVV52NaDduTP+ip9NmI/e5rG
J7p9BkBOzUuPip1UBwV69qpquAS77xVXnZGjgtI6NND2c7nrCvXHBOIczLV+NU16
J2wIM+UY865aO7erlgxepff6dA5BL4/Pk5Nl5bz6gLN6k61Nj+ytvwlLz5fRJ5r6
`protect END_PROTECTED
