`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDlHcAVh1PKU2xN6hQ3MJH/VZzEp1sCis8Bye3TzVT5+Ek0+NypEzytd7QybQDif
g0Er8NJZGUnwHtOd9FlOdPu0HR21MKDdPnqmxCNG3auLxnc1uqxOYyW6rvk+qQDi
KmUSpZflUg3e5D6Sr1IPVZJfQeWQccT/NyWgevRzD9yjcSml9ZYwL9VFveBRBxEn
2p9S+cTWxILiYeeip82QkEI5floNHGj2G2ocVAm9YMskLMMrf23y4dkjR0KS0U6B
6hzxihtXV6s3uOknxCNin/AlGXUjZw2zy5MNVaDAWJXVPmH7L7rrSbmAbj3ftgI3
9bDfw2a4reiV9N828YgjDxvrwkoqpS3xAUfCk7s/cH4Pmys2AeKOApu+RVSd3Zv5
85Y4d7wnEgccw7Q43SEBCW9+Msk/AN+TcDO8Q/jfOZrx4G+dUd1bhsfLmwQgSM4J
qgepEwlfMCQW94SKbZxbrX1NXb3jcss+hto8vgiJBBtpSeyQsBeqvfgvt3s0b13f
k7EdZabMSf2JuPVj38CeZZ44fck3vnUzyzrfpbo/qCtI1ZcL0i0IKLR1hqjvRF+w
i+SLD37tKdhnlPi2CyrVQJwFTF/Iz1HdxjXldEIUN0XybKkglepWCJyR5vlDnjqS
aTvveUMSqm5xymI+Brd9Mxtietj4aL5xtG+/PqQn2hcPM2og7sqfOYKJrIrIJuQT
7s7Kfw5P54+W2RVq0PS7aeFMrpRud5CH7j5Rvp4jLeZyPhC/GxFUIS4tIIZpFIEi
kjLMPtQOZg0kqczXzgNkUiOjUhNsHlUfJOji5UaY4F0bMY9cd/4dFSjDoDl2TlBq
bnemW2hhOkBOimG/BpLfS3MWe5pA/s3no4H60zIzhbbxFTZ2ZzS+ZRNvTh7+JRas
2+rVcEcttCD6yaM40tlGqw==
`protect END_PROTECTED
