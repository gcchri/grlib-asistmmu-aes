`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/hUXhuPNJUL6E9bZwqKASMBfZ+k4/AQE8+9O9uKCJow0XK1IDLHbK1YUpqMhMg38
T31rTznlFWF88esTxPrc/WiM8/EpsxFoilcGllPkP3dcRJksjv2XgUXNeHbF/yuW
M/YLBckJs48Oa2tAz92qZygLBPcLIYAB/7GnF4lEH0ihKAT/36OWeZsaSKcYUHlA
gBS4uc2aocf1M8yf3CJ57He+XgSN/N3iYYsvOIovoSBjNijaE75r4W7HqzVEXhPM
zgW7nrUovGOXqgk7x+jJ0qhyXuPda0lRmTvJQc3m5MsuIBJFElrG3nL8wNFUZvKE
E3i3gqgrumTI18P9lDQ2XX0mpGS0HVAGlv5Gfa6XT5a9QLYmTe34WOVqFmOy0a/D
q8bJbPwXC529aB8DXvrO2PtZ6OTR/LWmoCyWuyZjTOJwFrKbNrRQXWByf2H/StOY
`protect END_PROTECTED
