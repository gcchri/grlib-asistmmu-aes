`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8EjtKckHVcj2ExdOSoQ5ftrANEq9SiNUviICQL4z1XmEMGENLcmTXf8xWk7ZE8N
W/M41SjAP6u3Dyu0IVupi/SvE3AUXTrIC3MOPEzUFwUGrX6FO7zuM12L3UCO1PHl
/746D9yrcqP9YlZ6IYivaRk3e6dytY8vRFeJ36WwKoyNjwCwV3lv6TAtqDLwsxES
4Ykwfs+O40zjVujHBxS7/0+K/IhP3gxfJ5oyftjDS8h/8i3ywO7Sq9s859jHRZVN
LMhsQDoVqX6EVQdRgZXxZZlnYzP7iFgAoqRxMx1/a/iHAbECloOFuPlmtyw2Q7Dj
`protect END_PROTECTED
