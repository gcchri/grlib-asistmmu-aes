`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Psuwqpa6Q4mXzBXcrmCJlCrz5Yx0mvtm/gIkIza7w9naSZkxmgFKNVTyxLZ/fc8+
ifC5ybqhi19J70wSGw0G2/8+03NElBjA+GaVma0XFDrf8D72LEqfiqNf22bb/POx
IOszKeH8Ds2axMr9/EiZ8JTaVTmYiEmKYTWmMw6RD4VfGgVv00sTpDXf08ZuwwDw
NnVnB3z3SIq2UOvDhUaJykw8eOOfGEGkYQ0Nxtf2m9XpsbaeTyuwg5cLauaMA+0H
6QUzlCqRNNA4lvF2R12ZKwRRO33qY51ro+5fUZsgEqg1wUq9fw0YF5duxutmbmHS
xfNSuMXHNFUSkYZBZDmyMsxmwLiljALL8Ks9ts0SKuxuE8bVjkXfo3/UXQVyyW9Y
tDqzjlaGd3lnhE3KRf6mJwURZuXMiLQ1DyDalpa3sgEjuRWlHkGETCXM8bf7ne0B
JEYFzCNyQAhHJ88hKoRnihZk4BmfBKj7M9xW1tHF5b5xVQxNkKxjBMHdCtcUzfhl
wXChXq3ecg1gQsuiwLHa9G/YtyN5j9vOf/0jgmpciaYYlnYnEZ7mGc7S5emngj2X
7Rk1V5nSXXJUuq+lfw2bsIMo1TCDqjEba6gnSnL1f0mr9OKrlMKVFMbn3LkrsueF
dMWs6vNDqi3UK/IdV2GK0+EE5aeSAt0Trk9zpOhWPfUZ5B6/DfQn7bXY8mC+AtX+
jW3QT/cPhicloQAAZMvP8LE8l1K58+TbCe36rKvaUVIlzGrZ+YuC7a7PKLBbEndS
RnSJkHxtEb+cNge5P92LxKObp3KQPwuPWRgBNWyEzUmbg+wDN1Jy0IpegWNiiNW3
wPI9/f/5iYSDJ72iw+P1G4B5BmlIkgyK3v3o1PG+okUO39xGpWACJFQVcd2u5BSP
FBjLCIkwiu72YoDzc2uYJB6Dzgg4sd/OvZIMQqqoZKsZgiiF7hlynggzmNpVLd1g
26BAin5hvepJCivXR4HQ3tU5+gJrzdcg+2/QV/CAfKfaJ3jtrtkvB0DgsS2TTUZ3
TfY4cb/K4iiyY7+0dYJcXFnW1Uz2VViaEpp9YnzmMQH2A+7TTMazWj3921cuCZNw
Vpr5jovVGBMzOD+QasZbGPPI9vytZPBCBz3qzf7CZVPZflaG8xVqkOUVWiGS/ng1
XUBS+2LIGnZmDphGRX2+QkcKyKJVwumXmhMoSw3U4kPHxeyTM0H69OBATqBHhAYc
iYNOk1lC/iN3YqJtc3Pb3pA/Wj2rMraybw5iiy/sQ/LwK/LlKtf5yg6p5tOf4b6y
fLQOZ5j1ZPI/FQtdj/7RLyQJQCsDy+x3Jhn+dAasz8hp83h/CfVDzuh0LXx+ANLN
xtx6aHV3PtV4sWMNZHFjCjtFCzX3/7fcGAVVr1NN+vz73muLen8YqlxQefJVqodg
F4Gp75aJngtiOny0p2uMHK5Xcr8AQIL+ZZGU4h5ex9To5m7a7pAiqk+K1cZp2lmc
USY41J5rEQCtjiENF/n+gpksFU6huAzq3+U0mKkcliskiwhfxke+bceKOUuHBkZC
dy+qjYKdqhMvUXepEyr0n4mDShquShB3phj/h9DY/rrXxcfsB6QSHTHg92TpGffo
8RTmp7llqTSCdgzfAAyk7W6AbEsENxB/E7JAv/ow1HbJJdLlQ6KHrracEw3ZAnvu
HC2j5G89abjiptrygojPmswazzw+Rx/r22aygT6HqD3IBj+7AU2NA/t6OqdYi9AU
K9BZCc3NMouguMuk3TFiMmirbsEEGoDcatErjUyNzsbzJgfiQ2s9yITHVYJpZZg2
V9nQbdk8ZnLA7DiddAxiT6zYQpGlrmo9t3qI7fUB2mDEIHwBrh3zWbH0tyhY0ONZ
k3L7HsJAbMpwRKR+XouA4LlQRZTkoY5YA1phrf9InGo0FcQl2hsLD08O0Bp5MTMc
E79jBgszr01uN3VLxUzX2pRQFsfcFYs82aWb2fC/IQpXLWiKBCkAQOlRTUI4XCHx
EZBoS/RUzYuOa8xeT7c1Oa+FBiNxveDRGnYqelzan7XNnnFai+VfT4apneMeAh0d
k6/nbmxvx3THjTlsSw56aRS8cU8cts1BUW6pPSu89LKicQnNoYODZLgiYRa8dJU+
F85RMy49XkPHovuuC95TzCrzJ/2TMGR6bqawQa726peeQtnPYBrYgMLVVXUBf1LH
MWh8v+XYH+ochC9NSNPFXRa+rxq/QqgV+uQfC8cD9OPWMaLvKzx+gLodPUKkHa15
XCR6Styp9Zi/g9HC//jLZIHztBJA7F+yNVoMY6vNUAi97ZJJD3oV50bsW6zJKsga
ND19oHDYLq3AvoFh2Tq7VoW4780iIOPCYKmEzl/Agzeup0cWSlBBDzPJ8vlBrLPc
/8IGYBqBD/qZH3mIJGvFjlCWHDn4cyfQY55cXZ60YpO+PLcIwT48DJ+BD6mtISOb
q+fYfBj25wvAt52bt6XjbQ==
`protect END_PROTECTED
