`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ba/urk9k6JWf7fToWDTExwSCoQIeC3loMzd3fBNI2tdCCuJ2W7N21ogcOcE1S5jF
4C+SiDM1vsX5Vs8knWskE7T4vt8SUabg/sqDFKKM/iJuhi74fDMF94wxu3vR1m1l
dO3E3oPC929WBJR2Bh8kytLpUughs5qKg/VyVWCQC5dFgLmkAqMv9ci3+yqPDjbi
XTS4w1wFVPsiUqz9v7y442y8K8HgSZZ1TLQUbNumi2tZlDe+e1HZFwviz5vV29Pf
8kaO3wgEaF2L32fo6l6kxj3ggenAjn39PN5uqY3NV4RmmC3Jk342Et5KnxHed/Lp
RGnPIkbP1tSHY/IwH1clfDUFMDC8NbtraqDvnlGMI6D7jkgAe7OogXPh+qo6YOyb
jv7cjxRlghFiC0A0vx6rGkk/nPEmv0oYekP3Z5jHnmzOpxR+u67f48CDcctugkbm
7sOWHcIxhOnatlnqN+DvDErIa0tTU9J9HA03FkziLndXQSiSUqq2Qy7vP4G38GR3
QSiMR67Kun2vkN2eVG3X6gksENOPZR08KhJdCmVD4ascoQU5sUiNnh1sjqzgD44v
+2jtlijNg4ZnoRJIdWcsBVh6TZbZT2CUxA2Bx97n6KzDEsj107OC2Qvv96mOYiXa
olRTuZNG5BEcBPDs8PUqOjipoe5DW64nhgNkqUFHh8LqrPpAkL+/3glHJUfItxF0
xJRpD3xI+MvbZ2ZtWk68qjvBSjJJzRlCVR/iQwcivnaQ/xtxnigrSPpSDwaBKKtA
1WudNgFu1D360mn3LDL1SrhDAUX1hzPS6+4Jpel23eR1DmMxF1cqLVN3v/5b3Me7
pVNGdzjZXxjqNHhov3wNFrumVq4JEo52lfC+oOkZ7Fk2Mw3o8ZJPRRXs2+6GttcR
c98y6O1yy1rQVhW4dbDGv0p6gPOnCw0UmLEWIkplV7aKxporpPhHA6jqAYDGkZd0
yxsxEba2QhcZlQOGmS5iUG4wd9YtTGQq1g7aAy+g+qnBxPOIhyUaOjgB/ICzp/g+
h9FVy/4/ZsGYXdGrGLcH/gWBCM6/bvYcL1QenN9qjxNcPmZJUsljYND2Gi4Fgk+f
Kg8xrk9keIhQ9VT+0DMeZiHAJaj+KZG2V0wQB4sfzFye8J50FehsVv46udVkepvC
`protect END_PROTECTED
