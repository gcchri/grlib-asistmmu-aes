`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6nj8Olo8TGm/jLLenOuNz2SoIdlHJ6avduBd0TS8K7vhDInmXiz+ANY1BsodcNO
Y75SgkQi0lfF0Zq8f7rHPiF60gpLaFbSxuf8fYUze958sqrocvepHfDjWysT4+QW
kZVDkUT20MlskgMGsWZ+AJEKkd4NcNb2zS1zU8h5zF+quiIcDySlXpkLlng1oOqZ
dJ470AYF2oacGPuGK61xBhtyhTwQ3Ofg7m2awpqXjDWNWXxezsajxURbt4jssoS2
VXhazrL9aT+UKFsfLHgweA==
`protect END_PROTECTED
