`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGBKiVqQ5Xun0LCNhlQ0WhJLt8Oe9sIy4gFTWu5kRsITFIGYLRnsRfm59FlMxt3J
+l6fRhyHC3AkBU1U4ZkJXdvGIrcdQMBApfBca+Z6GRgExfMlhIZpfP6GYBmncCsD
dx5WvEv0dccBQ8sRs5Umbx8NolAQG525/rF4KgbeSUKLpiDPTtNCqYOz8JQriLeb
uP+zA1XUUHph/WSceCQlsUs0qaFetgv+wCtBNiJ3sRStlyz2uJIfH/UnrHeNk/Ri
pazmh/5IwWhLuZ2WLOS54un5GS4RdkCYjMI043MtzNqluP/YXmn1U/Vz80pxI6X6
2+bK7nPUR8mfQp7alqNjA0Hl8jEDXN/K6puhM3b11YxRYgYK+eHAbn2sQCcWo7S+
8LbY388ZOK2GIt4hlYmfaA6hQ4RloZlUmVHRpmZgeixCQ100/uFi0PsE0jOMTEeb
QFEsC8IarrvG877L88rULYPCSsIozraELqjkzPsb51w=
`protect END_PROTECTED
