`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4vWcY93CdVGQoLQhHVM33+Y7wznr+c4OhM5lQDpv3V63YhQ6WFUaS84cCfLLrWe
tab2AmceVWCOdvnV2Wv4MJSssAdVpbUJgFrTY/9x+V9xRwNcy7utC6+T8DwPrqFJ
h98Ck3K8qebmvurlSqd1XiBK8tOTuR/YoUzKrDi/Q9r31O0FsydolLy2VO2YLyWN
2cs19WEfW+K/Gc6j17jxMDGGI16Fy2O7tgoksaYVONdRaEolJFHr3VA8dYKb5eKx
3ekTTCZIMdmathmdfkqbgVMB4vIGQuWX65zcxrBjljeDzBfnOL+DqKeO0lBrx8Pz
jJ4bckV7Se+DDoRqj5gVcmcGcvPAKofWgAraquMo8PCwIiVomqr+FuvAw+7sNU/8
Hf1PpeM/lCNpyOTYRw7pDwP3SW5cpFqBLAagAI3SnPosq2ycobKYaUeChcvw+J8i
R51+slF9G7lhsZnXo3mpr2+AJuftS62U2fsHohN2A5zkOBqEFCwZxrdCdGsWIzCG
gdgPBkFN6w/nhG7fsOPMrrsVSzgwSH5q51umum9aU55QjSCbBAdocRmN5N5ys8cM
w8fz982pkU/QgJi3eC8vUM+9bEWfuAJV4l4xtFbl/dNpcz7869mDsHsnmF608YQ2
AyzB2+inM3dT0rT9KJEXYWVHB9CV6W+qV73T7MAMGJuk+2oLbj46EyiECC84+aNZ
x9wEAJgctL3j1PLvLz2Gq3VGhUBz4cFGmXMGn8as63/j0eg68gVHHaDrjezNoKNz
uXFfaGlmewZiH6lKteWnI6GNbScERz2rMMUQsfvSei2aZNaAWM4RGp8foyNJV8k0
lguL4qTCcj2DawTI6WwwcNkgbn8mOQPOBRiPo2JcaFxjRj7ujtA2HIVBERb4Jyz8
a7vFcvxXGsrbQW0VjRig7dE266wFbkDeN3SndAzLJOG+fb9EU9AxPd3vjcE6sj90
4OrDKectpOZMNHABgqe3N/cER12mDLzQZ5bFDwtTATCq7eYYkHUSnMZn0dJFKZB9
/60gU2VX4+TGRqIBugcNfUGp//HUHxXqm1QnNRFTY8iNSQSbgWs7H1x3WF9Qp1tR
MqXjHVaS72orKjh4eloo9Mttva4627BHJu38b1x0SBScBsu+cPWhHTw3ioa8uIAQ
MXvXThW99AOnsY5Iiy/0nTGlyK+wcExf4q1TsYojY8zIktpOIP1ZooiH9qYIH0eq
ppA0OV/K5nMkZLcIrtCBXZRRGa3jsuU5Bhc/He5HsT2Rv8qPoWjKFiAE+Rxd7mTO
GBKVE+Cnfx8Z6uVO6BrUBYOPbNBHSKSkvpRKj+YunTRYKfwdwiAK+eXfIp1VZ/5/
mZNdWE67VU/8qw3H8l8LP3oZLuqph87KqtAbsimOINVnXF+5LPKfa9Ud6AoWBxjM
x3NqkYGdazYTGIxA6y8IISrxU1PT0F/WjuPgm9KTF3PI0i1y8IRyeFMOyO4v+E3C
3MEMCdGyj1xjQ705Lz5s8m75w6Jxu77kZ+T94N13X0JmYQJS8h+/VEYI7VFTJKDZ
upIxc3LgBlggwiJw0Td3JgGKpLGh0sBOdYPn8lhJvb8=
`protect END_PROTECTED
