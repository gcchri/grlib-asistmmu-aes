`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r1UHynrp0WwzD+XdYAU+5AhUblgBruQdhSjlng5K49YOiUtjaVqVCbN8Xhv2q3nr
Ksp56yblS2XMuEp9MIN4L/gnIGoG/CoeqGLt2MjRDB/xGOWc7QmepGHL+u4zt8XX
bNdoo0xUM1jb3FfuMtyIPNT5f2sjjtCKbVYZ/M4mKA+/vcA/k+8Iz+IIia8Jp0Ns
XuE1d4qaJjQxgaI4M+SrItbKweeK1fN8sDxME/lN5Q67Qi5/7HAP8dts5PcJD5Rz
1L9YALStH6rtDi7clQcanpD3GDgocNJyZJlFnnzczs8Hrb7N4aVzw7WGzPs+f9MM
NKVZ88Pm7iFkfeLg7XU1Dh0s/EFAtpa7TSgT/Qo3fcppLCuJsQGksRKXSJPtUmLu
tN+b9kllgZC4Z+Z8axPW7h930RJx0LpiRCY6M9sPZ4XbHm0lSbJNaQWC5NPcia46
CwCjVoLaORh2t3l8R++/PBDBmnhEQvNsaAosFdy1ZgF+LqWc/RepOpLXzjq1x3mU
/asuILS8J/AG0d8K9SSi1SWIpz18dVgVFJ/RgEjy0qsjkArLqnf/lopvbVRoFsaq
qo36xKuIUsVDmB53wIHvArTsRTNaL66WZre4br6vXMegOmcFCa41aO0cF+0HWErK
T/4g5xS0apcUP7Be54zwkXVuHILuGTcCblLg6eZMp2jRZBZ2DbaWMgC1JrniN8rF
Nc/iVk1u2KDbSirCsdoQU2uAKic3hE6cHcoj0MqP3PD9tJMQfQYXIb4mf/O6FnBa
sOP8x6x7zpspn+YZiVyphmSpr5hdU51IsoFrb2yf9+b7FsNsEvECy8TdRDhU3z0f
fP+XXXHUIXDGOxgwjHd6WtW+/KYGlfNVdnyQY9pbN0lEkXZVDt9M0nV6oKwCCOql
mRv1AjBRt6qS6HBAnTkkE800u0C/+M3H0SebU0L+yvusaPOLNWX+YRTmX8FcEgDd
Lb+fPurQlJD7GMhZ9/onLWMiV4rmDTgIpmDUubpFyYKnwu3ckOTDXe6pgnrFQ8rA
Eg1lvhCFYVfQBDl2IuE1QRv5QH8jrEbsX/n4Cg2TMK+Hh5zyxLaro2UGrxaTNA1h
mQxN5/afWRm4pzCrZ7+lJ6RdXmscZRjexF7mgJYxXdkiLZKm1ZY4wAiXxwENZJTR
mWQYqg0cQXa6EAl72yeFMMh1V8id++izlNCd6JVlh55KgZsqSJs80LrJbWluXQ2b
YganCohn8rL632jseh/ocMiNGtVEanEVeygPD71OcU9ACJw6dBGcc/4NPDPfOPkU
LjEnIHD/or3YEM+fYJuL/w1WCChoPrxvrr9dakaT92zyqVgUvT9GcW8d0loiwr3r
P2Wv0lackvTuBwhFgT1Cowi327WnUoijCEKvVR5zqn/rT/TXCAwEiSjbhk9mcU08
0K8BjI1qe+moUBEPxN92dQ==
`protect END_PROTECTED
