`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTG8qDxWWZ8UY16+5kJ6Ljf5/XxN9u9wG94Kk/t8NbneHvl+iujKkNAsTUfj/d3o
hqi98do4MaZGYlnmRdGFNaHwYElYZyUFyX/D2KKFVj0ssS0nIdP5KPeJfDr2TLVE
uirPX8e4ADGIWkOejejqYbqVw2liq0/g4IbnC8+9+ZV+zzh7/045Uyyl2Fd416H2
gk7zcdrnoNuTLBfikZLE7YB01bJLQgn6M5Iak9tqUtXV/lTMrGoG3uAtjR4IiEZR
+IsekGnn6kUZJL30jERGgjsM4RWNE83UNtEsi2yhctgEhh6AdXxlNFsmnYcwPvXa
ovbaeJAo8vftg0yjdTkWGw==
`protect END_PROTECTED
