`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rv6iBjK8CdAxbESA5ZgbpsQ96ErJcXK8j6b0+qidv61DfAu+Vb3gswxRbYuNpj05
03j5hUtc/AeGxBBDqd3Xi61530sev2f8cy5XJsHIMV+92iCNo7TqNfjz2LW8ppVf
4z/wYZ+Y3GBq8Ee+cfdC42Dj/AycCbUCtPHI9v+R2ZPFXqE3Mjk7ZqXOkgiyu9yd
mbRmy9iiDJTB+MnGH6sGEfC8y/VYb+HPMP/vEkFntkWAiHvX8Mkg7MVN8cbQ6xhm
xVf6zQUHa0UpXGMOoRheuvqnKxypqfPb8k0/Wm9AjRqFQ8srCw+uJGmimwuoXQjW
Uo4wL5ch+ubrI4Sok4uAteTrC070p2d+htwDdA7VUVkE4NrhDvqU80EWrZMt+bwh
6PhPndE4KtSEyZiJ75jZ9fgb8Va28BvY7M15AeyJef+z0tlx9S6TKxEERl7Manzw
WWI5cQRSu5Z9rF8D3OwQukm0mBaGr2OI9jSFN/HaBBXT+J44FNAF9TUAI/vhZNrm
Dlv08AE62Mxlycf7fijczc+WTborvYtJrLw2pyABe9wxSScAIsM3Nrim01za3i7T
vVVigvzX6//M2vGofAjeDJDUhE/Kw/PfU2SB8awW0NNT2ezBzw9Zsna6EPWZ8iVH
NNLf2esvdWZkKE+7ojfGeF3wy+zTsBSQfPYX+epOPsuyz2JdSrdCTD8uYf+YJMRR
HrcDnPQ2i+oJWcK4SKSks+enVUN08/Pxsfbxs4FLezJANIOgTYv/i9uXKqctRzrK
Ff62Ukz3oJhBWGQesrRgIfvqJEzsvQoRUa5ABbn/zHo9708vNxodVp6JGI5k/HEc
qk6vg7fHb8KW+k88kunahuTOBFbFZio53o+jIY1bAI+AnjebNYNY0N/J02b7O72H
1Bey319i8+muzKsVgIWXMmP6HC+ZV/wQqU4qqe8uAOw8zSis1wkB8zeFDkLliIAY
axQ4sR+JSpE5LcW2y0gu+9YPyACGsScckQlgz75qoAtMKREgH+pIsz8x3qAjQIUQ
KxxeRed86UgL6Ypo2Ks3hqy8IjkD+053LhDfVX3vTfsvjhdetYAKitBpjTkbKucJ
hM64j6NxrgcWxu/qfygcwQHmxfvmBnPdXvQ88vn0IO2/7+VM/URYODnKLVY1sfEQ
cDKvNw0iODPUQKfF9olzEpE3gM+DDIk8WYLVhwZ+crcHFZonyJItxRBzdiYQnwuw
5NhRNE0kX7+lrHcyXetodqgnrRuFvecj0pDQFHxbcXg/uf1gxoh2TUJkujucH1KP
C8F7MwPV18n2NnXfKJrIjrkBTqKH1NdNSw0ObpKZTQ6mp8HPKxSIoyQdxnuK4QVl
zLuxe7NZGTTZ/SOskdDo7a3tCAKcCFAsgj3K7daTZtrfAnQCzECnOIDDU0xQkjqN
O91WUD8nIBp86tV5Rjc7VCvPgVEYXKLNZWZauVKhrHHgm4uVa1GeLYxqtfpM6N5Y
KD1v3YwZNkn6SDmS1on73GE3/Xgo5HHbwiIfr4cI11IfYVN+g2o2Gscj5HRc9OF7
CKerFLjEjtsucFoFT3zhZjUozqoaFlZAJ9VrKKc/mGwDb30392RseGhTqHt94eqk
alfL94FU2KNpTxqkLpQv13Nu5HSwvSYaSdVnFPf+uXXIEJUodxyPXWCl+ANNLcML
jKPpZA5lC7b3ROBHqbVlAPE0I0m40qYOuyWvdMsXaar1vYBTskiVLnfe2/trV+42
iaJEbEcmTVHxJWZNYo6B68U6VLc4I7dTvVUoO11nGtqS/xLnafB4hcx+5UJEwU6X
sBUqC98imY80FjCrU/xaNeFOLTdeDnLMWTyZFjVIdvPhAw7M3bzOH26/zdvtF+vX
Y0ob+bh+9+PK5lwi6k2nfxjJdE87jCRSjpLGIBqKMpIDl3D63aPliB5I2sfqEFDE
X0mM1qOsCRzLEvO+a3SAVcp6iyyMgVkl8NpupT/FD60wFXxOf34tYr7bVF0gXerb
a29MOh3L/W99fcB+KgzByP0IKjipx+AXh7xhw5kfhaVlezSt16nr+qI7k+lLdQ5Y
o1B9CS3rlAqC47uNAJEsOizuqwf9xYCBziS4F9q5DA/Qs456srsT162vfCOm22SV
6vq+2noSORvqJ4bNhRvT3/BdFu4XsQv5o6xO2l2h2C6NqPFeHVjI64Z+UoCjqojx
`protect END_PROTECTED
