`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yy6lNC9HGW7U3HzkFirPok3pMKuVDJKGco25KTcO7n848dqz6NGF11y7boyTzxwk
qCNQ9r9MPP9NgQeF11Wk1LztWAaW7bzXHShj64ZEs3q8Dn3by7yILJ5TK9k/ITR3
I/FgQGwkCmQoUZRBjHULEOwyFP0R7pLaEW/sBO5+4pkTcgSa7RPZzFrnybuVPW17
cSCgHRiPtyI39+8rqDZKX8XS8kQaR+J6rvszCc3AhcEPsR6KAurVnU56SbWQn3rp
hwvGywTMwUos2DNegDoaIr9KeTmklUO8CUDuE6ESKI/JEJTS3xtnn83uHO5zujEg
qqQehBPIZSSbofv6X8i/Wi7kdlSmRfgAlVXiE4zzNnSZs1fgQFlLcuI28zKnVh8T
QaTBkSdjDSUfZra8aF5vlXTURgSZ5lE+aEzpb/xb9NSEqf8GB/EfchNjtmXsonIX
D0TM3+mxnJ4e2yfHdywMe5EIJfg2WQ29Ov3ZrvdlDus=
`protect END_PROTECTED
