`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0HxCqOUBvKnTSAsAomFF7oLLCEDW1xUb6AdXJ0uEBJPI249qxPvFCfB+h/ZxEUm
5mMOw/Hw8O5dD3YeGMsoCd7fV8GFUxzde0Wd/rOG+XVdCRnFpKkEU7HgCO+IVu6x
lqqA0Pye/0ZxVThBzGNrFI+ge/CLg25VBAjpA3AQ3TyvQoh2vEDhdGAHKx1R3bou
sReTlaAqePvOMyh+zjkESQuMii/LoxitMe3J91x/5ImZys6Z3UxOZJKI4z/WFB5s
o076NWrqYRrUEyileukq2587NZpdD0SzktKv4nWR9VI=
`protect END_PROTECTED
