`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjnglA6iLuUdr26tvkU7oGpuMVbtj+3wKx6J9HktwkBWS1xx5fnZdgyi6e5OScSo
ByfzQysG9wcmLyPdAzONZ//TNepZBvTpbO9UYc0pt+SVSB1zbcg4lMVLkd7ZB9v7
xSdO7K/Tp58QktQK6RemIesHJHrj6GVcZ3Ad7So7wzxUashtLgLPqIjQM2XnxXEq
QLC5tnE0gaNbNRS3p1fEZ81TLcqbQ0u9yYzTX8gWGy4GJvM6ikBLPjCUXoP+QkZA
nEEC0lqHhRvzyw5DLQogD73DEloyAqhQd+PfA4Y1xuTJEGJZDIUU6HAUcem5ZFP+
ljXdQXWf6jiMCY7L6QVFJCFqgeiuAndOIF7RhIIn6VacsNXfTioCOL9CqIa8JxhZ
jAeOzZVnkvDQcT70EC1QAb60xtk/rt1cgssrBQiyNvu5j8TMEi0MIMhyWGOr24L9
9CyhUPEEEAwY6B2lsFAd50W+vejtCIJ0UVv79G2d9OGTRmKkRe/bTL72BMycKfV+
Orzvuq7w8hyv2lAjfeoLV37AclW62WszrVaVV2iJkMb3QsiN7qR2Rh89ZdGtG2aq
xPvT/7FXbVfwCOQq9Q3Qk5Xx9OlX0SD/QUavWeCz82a1IqAj2cwUbbd5HpJd7q2a
vRx07DjjoJwA2c+AFvc/lMrUjqXSReCQDc9bGLwNaaCg9riF572vOpqn/xPMLtFg
yINCOmwRdfFUlLLssv8bgA==
`protect END_PROTECTED
