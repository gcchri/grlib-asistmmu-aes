`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M5NL3Cxq0kitZQsVQro8vKeBIfTzPmy94yNKCBvloF+/aOegu4G67t/5sjtvihs9
gEW1gO15qlTIIOERgXDaHt4nLx4BPazkOyNDHA13mtG1g/cwiCDbPdUqcKN/MUKi
EW8A4sFt5E3Ey3J52ooBBAFj8dytD97shGbhPiG9r4qbCMNuUX1ObcXDk8zRHJtP
TI/0HoWdh210H7TvB1CcuZ1k4D1ww95kmydlxpAvqytESMCyoHtd9CP54RmUIRqo
ieD0nLLkx7qUxqt/QARiRUojiqHKQSF13kuWvOw7Zf1xFC7OMx2znZlDg21EcKkC
ZrsPW7Qxo7OK4qDKeXl7hXIRNjF6PZ8UJt67YQSc64Fv7L6isDAPf2J7AERxdaHh
NSxL3N60whf38l9RzxVmPiwm/W2wgHi+NsRM7Jx9fMCSxbYM7MWNWiXf9v6C31Fx
i6NKtYRvUbr/tmTlR4T63Mva9iidY9KKcvIZtO2h8kCKf2eATzFYJ2UtGp58cg4d
fVkxj1B7x1+5Yc5homcviTb/lllWuwMlLTlLSJ21RRVDgJdikiD3RDDoSFtEO6VN
HtYMb+Q91MZ0Y6uU/QWaD+OS5jvBkqc8DBK97m96/pFR0Od6mlDCzlvFTJhJalC0
hyGK2un/sfjJNrjgf2WkTg==
`protect END_PROTECTED
