`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPy4sHCTjSspa9QOIyZc20CQFNpfEb132a1p6BQHdxF/mRCP9saN+Ue1DqyB/Onf
fOHFhkY98x6HUgbU6gEiAgxCQAk7J03rupc3gb+akfQD7lPGNiQMcgHFOnUa9Cju
cNDxbPoYkj8GHoh1I8CucA5kf3PyBLLk5sERKTH6QQvw2Dsz/hLtbM5khDbPr4+a
MgV1DxRllkrVvBW9a/9pyqJ+d86hQNT8kQZwncGOfe+vH4eGTVof0dArJ4tMltF6
52pQQ9xqSPEwFL305oEg/+eHmczCFrvxigRh9AOoy5fGBICZo7aal4YqqPOHBDRL
2wlPE6NwVQVpYydXEA1pog==
`protect END_PROTECTED
