`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
csXkBw3++yuImZUu92zJuwWtu0l/++oIpUT1kZ7krU90BH7bNj6rzuQeMqitAXvr
UOlyE18cJ+EOABX472sMu3RCDMnOhGmRR8rqXDZT7tC8JzVt76CXdaMjHL6zNEl8
IvUtDQUGULaJiIDtz2A4Rbne+t8NLT65ezgtoOvNqLLgioWXwuysaDU0cZYCWKKO
mgq+o8dhLhszxTz+aV6CA8AK5tMRXfWw0ih2BePgwl2pki8KPIRkI8kX7O+GEeqG
8e2YXOiJQwDkRQ4QHOA9fiJW5Wucb+rLk2NfBm1dY+Fj15t8XV+Eq2Kye/0Ylj8S
I0FEif5bwPSZvkPMolNbnw0nXR7Kol33AoHRAW7VdpLkgKquRQwQ/xrYjKxdW9eW
UACxRZ6AZIezxs4KQbGnRkyMEhLtIgyKUsOgpFg0+KHs7aYmdEMkXsXmLohD/dzG
gjftCITwYlt5EMKAyPpb7/SaC1exHEqpH7QTh7rX0A+lQ5lsIEuxUmIw7mtl1ugq
0keI2MAPMadTHx0FvuWdvCP+r8PZL80oz/XmIajv4yMOVCZeTYH5is4Bpg7qrwFA
9CiUauG8pm5Q4XiLunlGG0fc+zgvfxINOyJcYjMdeT0zUolk2ASseQyRRu3wPCzS
Bl6kbE9kV9zTvSoevrLkyjIh+tv/IRWi6w3LRed0kyYppHFZLSmhv5ttM9Oz6lju
yxisRqFKBbaG+Xv5odMqN5ptNIpblwQGmoS7AlqTI3Xca+UpAueK5etH2P58JEV3
0XXzkT2iojrmBSXYbi4EuhZsHUyHaSqR8JSwjS3NQ0/nSY3K3aGAZB9oJdnqgCUZ
T8qYccG9WA0eWWLvox+6d2kbGgFRxJ/jtdqnea+QqRMf4zHpTF1no9bFbv9AAhiz
z+YEYh4wqLIbX+3TB6j0Zfzh2EgHs0SOPxracX+Nkipd8guf04KP5N7Hdlo5y491
LoJ2sYR5LNFClkpas1MjbUhjjGW6hmm8tpjpFM6y7lsHiJ36GXPEqNdg0WMFuqwi
QevwVZbLvDmA7HCCauJeyOOujYgnWNMtahWROvN2JhjWjiLJg6r1uRdrzzoBR9TL
paYCh4EApgE8w9/QBkxevn5RfGnhV2kRiYqVHVMgTXn3/99ovVpXd0CAR8jFrAM0
GCrFYseAyexCgE78nCOqThzCt+Qt7FxGsdqK/9E8mpqEP0hGXHGQ+RF+l17l5CB+
+dHxAWWwxF7pTPRKPx5ScIoxCHGlDldIn8a+d2CzbFsgqULuNx+RGYMv/L/8f8y5
2I5FQ0Mse2jp/vbx/SBDiGYaL1kCqmNUVGhTTUlW2cSb2XPBhSZYMHfgoPjQ/Z1b
IXVpvA8FxC/EQAVJV6peCkq8/RSQyKugWRLC6bfgfXtjvX5aWZM6AOjG1nqR0SFo
k1k/F83Qqr/9m5GKT6AeMWr4yKaMfKNCZ4I/ZmnzjsNZ08CNSbsbZmDn4zWsLdLg
c5elEU5wdHMg7svGESTHG5ZU2FJoj/IwRSamJ6V2phN02SYO8F/OsG66RoNwaQrL
QZh5sE4HNVzbTpPNSc4bLJeVLOFjLR2O43LMczMIoGyQvVAZmzA9hsmcXRs9il1l
xfmeeq6uEZUJAqPYVV/sQBwhR/YNzutP84MnTB0OlT3d5POCvG4o2GGdZ5SVSAeM
GB032LkiLXLrbPoaOOngEbAFlSIctwrawzy8ZmSgJea3PImy+i7Xmgc2MUsRXEE+
/MXUzpGfgmTINfPwdn8AqUwEmk+EHYwlMgGqv/hvsKnM0ngOuu21BQ6YsrXtkF85
59mUp08KifV18cRqyLEBzXdzcvY2v5g8hNit/pnb5QlEuwA1Ib7+wkca0kB9evUA
QzJVT379kogbZnBmka5vJl8XFByePTVrQQJI5oI5fOzD3GPxWNM7H6Ka6UFSyWyQ
yxgUWuRSDfXzwOQ+583H+RfwJknZU3z2SHWz+WoduYlThceIiz+Q76p1MblRnRvJ
s88dAmnfrkFZjcXbmucwC/x7aq27NTNRBoeuxSxIWEQJSH4/rUyGBpEAIbCMSiem
JaoL2xOuNWJf2TZYtAfVd3cqs5vNw8GZ4nmE7ZKww3E8A0Mb75gNDkZ+ofp1E4PQ
t9bZEVdnRCpPyCwrM+0Vrr2ok+I4+VcF2q1VU+1NaD7s9L1JPkWG5zJkig73r/fD
uIOT1DxlNsZMqXN0qlAlVkZLHvx09Bi0WmrPAhc5mJU1a0CitHbyMLod7PfdZZXX
Ea5zggJYfbDJPv1/FyIVLxuVt+d5aK/nib1kCOJKyuW5CVbRAKP4y04gTwUm+9vJ
+6nvinJNd/MmP8jzT7V7gNplc+s1rILi1bnn9xtZ64pNFJV6gly9jJszOYOW7w/W
wnm9pYtyYxbFPCvgBP13xGCCUXmeBtd8FGEE3ZS/7q2ohGG9+RaEndSngyRO3jHZ
fNj0ESeqtr3X8jkO1aePkyQf4tAKiJOTeNtPUx3QBPjvxjqh1e95ZtsmsJlcOW90
UqjXGLOFwDuwvLG6+tOP/KmcRk4aFKkU8i4swKjZCYIVzDH2Hyc3l3ZTB0Dfzpmy
DjTZH8Mh4Fwb3p6hlojjNJzw/EE2L+ioeagpJv881QxlLbAq4ejApBEzFREaW7G9
al3qKc9V8g2472NmqzlYAc0wbDCk8xqljusXnZqcDY4xvuHIL0FE5f1n6bgmQUUH
Bg5s1ZxvOmFsIEu1q9aA7ZcYFSBTE3egVfx84EvS1BdKIGXWrEh2zknCYRvnVxEa
ae2Vgg4q634iFxH4oOAXVRyTvfWa9VQ3FUxMgpDIImOUyeeJJ/5aijHDZL18gOSc
e+xJnAqjRJEDGbsGV8FAIkov1HbiK/3fUGiCGlYZ0Y7zmrpOEDwmZuxAyB8Tdthv
E65+LlBn7UhoFCG2kVQn2mXTXYjbKymSQcazjOe7+4YOYtf/gRA+UiyDDcO7SP7i
MiCPGFE7Eb+uQPqn+IcC4Z6KbWigLjOQwttvJZHGlP7tRcdcpn6GCI/GTgOtm7QC
HxueXW2bT3/2mJSqosIKHkHTtcY0Wdo1UJpa57KgpVaDVNfHAiklBf0rzDpn7hek
6/cZxd2sgzAb5B0jkbcfzt3lBrD3K1cGy0v0Pe6NS4oJ+C3UvJS9tcH82TeTv9uc
Zn9CeiIagZWu2d8w36pBkqM+bUEgQbA8ueT5NRCszAwVrbgxZ32Vd7je22zooEZZ
lyoo8cLmJC7UnOpt7V2MQkeHlIdK7zRJdw9HBOsE1nHrDzhYmJUy9SEEGXoCHJjZ
+r98MKbSjyKQqn3OYCT7VuCxfUwEB2hFSDXlA3+nx/axfOoC7yaE4eRDlbivMPPk
yIb/sPFhY0B7M1A14/qei6ViWDHpPEIJhts7UxAzvFG59sdcqgvG6bBJgxCozcki
h8jIPEEcxEJ0HbBNAdxZThs019SEemHCPvMKOWQ5R2IQLvcIZIkWBzDbUSRM2xwe
qrC7TMHEajWun0Hh6+oR1T7dHv92GJyPAIL5u5uAMzpNhokg72iAGT5EQO073U7D
YIcnJATsyR4htCIMsFNTyH7eSp/du9MsCNX2OqgN/3lM30Ecpws2L5e4TieVGzsI
7YYw+0tb53C6MKO9BGiqJmEy8BbmNQMkVNeEMmsTO3sVlgNer8caR9ZZJQHXX3dd
bhHFSpqSmRLD7h559gDRCCgTZTR+LlC2AhgBHnt8YR/+YdvzVd9iy0KZ4vueC5vB
37IeJNjWACAeleGieUvC9+n8Gfu+CMi7fgOBaH1EyMv55sH8XsL9ZGS8pLvUaeD4
mz7/+bWHnr2GFY2/GdFo7PgtSpgQh/dO+o9dqy3xQRseByvTmMeI8YSDWl9gxBaz
sSphYrWNFm27Iezm3cKok6JEgzgK9uAjJ851OooAGpCKfEywMfYF+llbay74vqI/
WzegEVTWEawn2/pL5vMNdxihXlOfAjuRLJeaRBs33Hjpknshb0LZ8GMDiPkld9ea
NNgcY/EeD5ngVPEY18CBWRwAQUqIRZgA0hR+ht82gVRh/RRKL5/pwwfBhPT3qCqh
Tb61lfQ+DybUCLycp8jcGelU3wIimSbUy855AlDrQAIDJEzS8eKklVim42CxcNcD
yWLVgF4nrgazUfDPkiU8xbdMTAnRuhAtfCtocB429f6FtJM41R9Yr4H3ozCuykMJ
LKGOzTwrMYT/95WqT7ZECn66ALmeZ0ogtbbboznDOWygaLAa2bFlWMgKFFggPmg5
0ZUUQSktwdgL3+MYyP1tHbXdyw3k/S0waXJ1DHM/ZpCZZTy22SS0PmVzdtHBlk6T
P5W8b7XUIRP2ejXRe5liQQCtZ9amB4DwefGgexxpgbaosg4IHQHNt6qa0izFMPRp
Kg5diryZSZ9jr0B1ueq/QJOMDhjeASAR9+2jMUpYdE9dDUsVAJnb/d5P8ysFdH6Z
LaS8EpWcabEMGLFRnydO+qcMECAal9gU2g87TEc1t0N2WhO1jLbHxH6kOAjPPtUa
yEOl8OIIIiKALGxzT4qpVe/dc/It7X7JSAvC7Ljt7GscVC5T5B4+Vc9kD60fj7lJ
v2MpK6yX24ZERoTREy6nsbrzAamxCy7B5Wn3hXIr1soMxlqfdL359wYUnTdHwALO
848YwsXZbO0lijbPJEZpTVr6TbIGfcTC9irUmUBwhjR70bfTNlOY0O4IV7bgftcc
DWwTrfmOUi0c1xUpZbk+xMqIhXlacCqYzVKpTbgYwHbAuzSqWeKINka70e+qIng/
BqZgPgYUB0C+ok8IBuuEwLDy0VGZ3DTGFjqzKVhnUehOR8jnIZziOcSQbcEwoGum
mh477jMh0YwNur4PWQEokaqFxRLkXDfzskPDhFVUMgzi0srnzS4y6gmYSr6vBbL/
ZDFeBHsQJMkjvsHCzSqpGUPr+0tSs2tFYg5ocLhOlp4fsexkqsNzNLS5U0/ftVpk
cetMFc6GOHmIYCNGZ94MKamZTciRjRprtEcscIMMZkDIign7Kem7f+BWTLXSwJD5
OGvj0MW9LRp+MPnDC4rP9ooTCsjUN2LSk57Z/m+QVZN6Zycv+fqvF4BV4xVMFPT+
5VMXWlpTQKez2Ika/Fj/mGYRmjZGqKhwkFQNhxwM07X2xJUbbqMqtw98Rp2sSsS4
fHtlIYaMeGG9UlauuLNR8SCjh6xPdEz0usaANVd+Zvxby/a89MsBzTmhEDkNotpn
2s8Uv48miH+HkwTJ1yteUzkokH+dmzB+oXIwxRW11VaIn6toqLouzgaWOo5VhM0q
PCtf5IGn6iEiovpq03N3y6xnby6hl1j1mlCRPvTQRYwC3OVNaXmd6Ndc/9OS0xeL
wGswuhmv5jEwn8y3cIAN/mreHsIu+uOuPw/bZ/045H/cDR1Ws9UoGhZd16W8SIXW
QKXzvS9z4yDMnaJFws68vBnx5X+8ydE7Ax9Utfw2FgP1BwfnbPDqptVEHdzs1uvO
0pKHme9S2YcgXPppqTIg7pZRi2SgeUKGNcs5pwIsfkT6+iAZZCn4a09g0QpO9WE0
WKFo1381i2gFNu+EZP+ypEOaCe7NZGu6yePMT1cQl0iHLSmNyyGkFjRtoj/h8asT
y1die5VVU5Y/xIZjmjSsxWsKisnkEg95K2j8iUo1AXuWx+G26Pu1HAwyHDVJCrK9
eAA85r0g6CgwvmCGoPKTEJJpPxVCfjzuejXQMahJPkk4epYhURblsL0jAnvVyqMs
x3iW3/KoL/YPXxuBfuZq3UWrMgYthYt+KoQJCvnfx1A4owCmjp7w4wS1E8SLS6Lc
CGU1WZ0c7dZfLlKP9rI7HEN2x+kyfc9niiH+OEZO8s5v2puRPh6D6K0Zkjv8XBtF
N+xEWnDzKSNvC9LNxvJeLKwYHgOwtlpwBs6RyYEZ4ANfDiOEgOHbjQsKVdxFe9mW
Zno7DzcT+bKcdOk3qoV+bGxYp9aADuwuB8l4lY0CKXn9nfSG2MbS5nfDcaBOPYWI
dP+O4t6GgLXi5F/gSBOw5xYTyXg6FG9chJ6TUnz78B5j3Y1AL4YxVL+f8phLQorU
rzcR9SJM6RrFtLkYp9xgisMxjvSJAgBG+YkM0Nz+XtT3nZ/OAgPiQ1er+phtfijX
ROcHTxxhkBjsrboLGMHo1g3Zo0b5CNAbN+i+OvS2CerfcOcG6J3WvWv+bIp8DwNE
JVQbIFXAjY1X+IPPs7aCHd1g8teD/1FBV9AeBh+SqUr5mKIUOFBUHGaYOKAbO0kd
1e7W6N3kH2jppk4NnfCykTB8gaPu2ALTIaXVDIfYAOo9YPkU5TNWgESUqI5ZiHhl
EBDtmEJg1S4gaNgKOLbHZYOdEz0sYba4jb7aNm85p88W7OZ02wSDo6oxc1U1s9AQ
7J6sqKDkPREhBY1CMCQ2t5pugEXA94COy3J5Z9yWDbpdFUcuWKQgTGJrDqqi87oe
M+d9X/X2YAWBBLtbFp4BTfCNKdQFgN3ydfDx62PitQUfUIACgmNk86RCv7IZN9K4
+uBIReKN568oFrB3bnJTJeaa9zulYKz9vtCo5UM6qgfLCLjaBOOAbhGaPtzkRSpC
1qRp9V/5a3aqaIQTMJYRwX2Qeb1GqxAZOWkq4w7XYW5HJN55wF2nsf+z7bAYupT5
TEAwzgpJWr35IB9VfiLqSAAqW2Uy5P18cmiLU/bO8aQAV26CbNlDTHd5/lm2S7u7
RseSeRvwMAtTH/7motFgft68m1EjTHpiWmt5kxzG8/tBOvdcxFsvcatAnqnlCdNc
v4i/rWMjarSYXJ7g+YfGuKAwZHnZfAju+BLr5AcG8M78RNB4Uq/IKKwsr5KTQGlW
XuOpBxrZYWWom2jnwGSJKDsyIkjtxCx2HZ82eqeCuQToW0kDFIR+DW0c6X7b9Bx/
ZKzJcbXvzIzCeHiRhjo78wRW8D1tHdOJc6KRo9SLoy25U+MpzAO/O9mcKPgpLuM9
YuLoJJVPp6azfC0SCQe5H2lXNyXBE2eIpEUVaBi7e+HralbuVc+udf3qqjFbXeLY
hnxqMBDkBECR/ra/lgnTtXIEXXHzBz0X3TYN74cJ3miIzH6an+fPxIWAKxwFYX0p
XXKtNRqpG3UTPYoRdRm7eliJN/ZfhM4GrTBd51raEU9TSlGbFS+6NW9bwgSXCFXN
kr3ZvbFiwJ8TQF5OVP+bMQQvcINGYl5Jqh/VBtSa2CFEWUPQ5YYQudmxBpOvfM0i
D7pd47bAc2vWoHtHMogk2Gx6MBaPaiskjwWbcqT3pGog9XNxDAlfiLM+jcaoj1lQ
Wk7g+UVqT4aTVlXcZ427/utPDVmWeYvmJlmICFnoKiVnOKtI9D2cyFnam8DGxVXE
mBiX/YnRsHF1F0DX2698vsuMcWa4pvW62OHdgu/4HHTaoQBw3K97oRhwTHxcE79b
VpcCEBJSg7/iRzlwOpJX9bvUcNvDTf77enHdoqUrhAWzbRcGekA4byIggNQanfxX
eK6EPb4R2MDClt29nNSA+vCssM9VZDyNJ8x68JcnoHpkshNCUXN+HlzvpmkIEdyn
fBJyZOpVG1ytWg5X5mVSU3T7hoYasUONcoZTYSEjH53+BwPFQLaz2f/HDgYxzzfK
nOms2IZvzSOhY0MEZN545MnRfAyTTdtQBiwRJCEzcNAs7DG7B8tS3ZAPSMIMzeYt
zFRLr7OOUCCWq7fWy4t3ZB7P2IffxMvdxtj+DfD69fMDLMC2HXQoj7K5sJi6cFoD
6gEDLUc5/YWyBf1H9Ljb9LDd5vOZx0z2Ej7rcPwMr/oRb4o2jUVNo3LLyDxu7BCI
yi1OxM+z0bzm5NsebhzLd6qj55dkwiGhRlVZpyl2i9z3TvtCB8FBaoY8TyyGG1sU
7I59MliNiQhQ7t9yFMhI3JuS3pN1vvSqhX0RLMw3ozBsujLqkvfXzHm8lq0yyd9q
JgoEi+Nbz6qGpqNL0fYssNwSSvBHj9wYuY6Spn7Za4pmxn9O1Z3wu/BZ0q1aBFtX
7p04LCqf5FUL9XrjYjoGehjbnVgyL+7QiP+G/3a07ksmB1o5dB7P7Ek79OtAh4UV
HehHQ7NTgHlShf/upkEaoNccKKJY5Y4IGK8wIr/qbG8/jIrkPLxxueTsr1tdD1Wp
zoGkv53sHPbpu827fYyf/Ue1Qiw8vY0h/z4gml+pw2EasONcWFoZ695d6FNiY7fA
1qJqtPy35uWFfifNxKz01ljeeJOZl1iqJhgB4uXcrmWltbVYxgbP1xVhdVJga91e
J+roa3yE7nfhgg2vCSDn6umLONkf7LYyiQW4V+xThiL5N7ZhTU6pjgWMizHnru6q
rGozN++uADXoDPG/zjOtnfRgWcCWfdot9f8Gs89SvwA1Pu+JJ9Lg8ASarOyxvaT7
UnIRwcu2VKkelgRpf6Zm4TDHhzEpn64c+XLrKKz9EsX/16rlt9JUFH8kjX2r/gFj
haxndgTVEomLp/n7Oa/66LAo9r7B3YNUeT5o05uufXEun2yA7iEDudVO7cgth9wd
8NPGomCEFcAGX9Q57wnqpi/ZFweOuWBdkuzpNW8aXzXRkZv11y9/gI6uKVyV/ZuR
yEet2K994+xq3771Xvlw66aVwhjo9AqwcZ8th6qhor0Ugtnkeh32tuv/2ZFvTlbq
JLtdH1y4zF9uo6hGhVxQo4yGXKmGfUEtqO1NbgDAhGESfroVpFnh6MQ2nQm9b8gV
UKrlmdom9jUcARw6IVKtJKeJ70ZobR40zt4byRxDQs2Yn+nagEb5h/rrURD6pcJb
nUay663kwrcejpEjj+EW5eMxUaEqDaC96d6d/IwQUkhkDClF+8OvV0zM8jpEyQDD
nPckUPg0E1i0r8nYciturQh6NNrRuaH2qzS9x5oJE1F7nR9jBxfk0SJcz5mAO6OI
uatZYMG/gEyWL1qx+4pFmGijR00rhB5Z/P0EpVoCxRI8JGxwQSYVU8WVASlbl5B6
S1/ZHU0YcSceOLstsWV5evOjliangxoGPyNknBqs0J/osAXF3ws/wF6yx3SGifUk
JO3B7Uq9NuHgveSTIBRxqh97ieSXhdOcThI5buH4FX1YliDFBgy4yPRhfB/eb9J2
r9GQKHVls1ybCr+ODEnmWAUKxLD4Cir3J/P3yd3jgMdOfgfdw7pacl0EP2dQZhUj
6k2/k64pXB9mikc/uxJBk7reSIH6JTIz9BSclYEScHo4SChEYYALM/sFbP2s762A
GqX1gmSe04vZdKofdz4T0MnYDzo4Z8sHr+Tq1Xuqkg33/FHNGQ8ebbG16oYqY0Gj
93MztNoWZb+o1K9ItIh10Q==
`protect END_PROTECTED
