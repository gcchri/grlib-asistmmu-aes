`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ro3tyVv92FPDpOrJgs3om3dpUjhwtS3SETfcaBTolj3zU5+lPfyJxVwM/WAXHi2C
/t+QH8l1G8oV35A/Xl2Dt6S9h4ez0AVGcBHkbcdmO7AoIYtf5aZdae1XTXE4EJxs
rMiDy81fzZAEFZ0RyiTM4N4EIFuy0wSFNt94Tc4IRHCTOQtk4q7fFKfQJ37OipDM
mN6++jWGCJiKuSFEtx0te5bgBxsDZQooKJOeG2qnkK/XgslMinAjUjzJORN17tGF
teDd1pPlfWw1c8Zxt5i/beF6nzEp3BkdXVi1lA6Rt4F0qMTCo57GGw6aMiGdYrao
II1VNt7dvC2R38Lv9xqpQIgLv5zheZxzuYkds+LAnILS1igKQ8XaWSzqXLfpZAFX
FJOHxsx26D5TFeH9QsyssfzRaaGkblNZRFIvK/+Eue1AGpMi2jfXVygmmz98bWWn
Ei2wf9m/xYwrVtevGyMjuR6V78+BlJlIn3iq+egjBiK1XwODAETo1/PSdFenaUxs
RSu8dMunSTkLEM8JeJeX32SvbdRJYgEX7gP6ucrxN8iHlmLEbsWlDjKR1WVynGqZ
/XAXcVnm8OOyHLMqQ2yjMOhNoXtDHPFd3vorNNI1LYrFoA3vpCYos3mbsZo31+y6
vcW4Y3Lwn1JK1kB3AHgu/wZSMXdLL6KKTrLMEAHsfx4NYHihDnHVLtyZIlpweUFl
wn7IcIUKxtoN82RTCe8dwLfqZ2zIn2+LBlJs9Nmdl3g+mJEEUFss7X7a/FeVBoja
F8pwCb5FkNfUHheKdSWWErqFs93A2dJUjzGL0hqf9tzDkgtedXAMPxBZ60O9Y3y8
j95/xOWXfxV1LmmyLsj9pTfIl9saj8HjZwQC/EKOg8R3HUrP+Am1zTKtgvQIwJnU
Zad0fMS8TKdWTWJ7szDbQThmx7ivdWj4y1f/1bL8XERJydAtbWFLocSSTxC2lrL6
lS969Ua1uhhahNy6RizW3WyW8AIdqQ69F3ssUGYQR1lnxaGrZwUEc2o2q6BEI1T6
j503PVit4KRbffifO/2FREY4RQncSv/NnfpCxHAge/+aLRTYgGvI8TZz1GLAZAWc
V+Fi4HOgi5eyYpob2xiy/li/XOLnjeS26cuKMETMHue8uQOv70BzCS6Bzy3VSWff
xL2GbpJCcsrXr81BVQXgqIWQba15d0f16v5w+1dLJMuUY+FRH2+Z440dRtndm2NJ
su77l1bu8rYwjxAX0wV5pfvRjyGz2ajJTvnaKNDD36xo8HxygPc7RAPaB9cwHe88
Nm4/jukxNExdyrnwSYUYKKVtfUzhdP6aGpz3J+OHAFd5pDUnUL4Q89TvfTe5POTs
gmksWYdDg4RQS6K4U88qd2SNiJpV3N8bWihfw4A9n51vor+Pq6EuQ4vhPSSNWjYj
vLWNhpueIQ4C6tTPz0f9oovPZHVV5fikjdaR8jAaTblGr1hVfCuqmcPCRjOmWIcV
uGQ3HlNL5m3R12QJhHZWMdHSNrlRO7RTATcvURRF3exOUdeL2oQIKBDVWTRQXeMZ
apohFN+YAOHLJ36ILnffkCddFC7QqiKBkf9jVQeIATsEulnCjO4Mjbdp9f8mEBZH
8cC6OhTafLWv8Os8S6QeQJnj0QShKgooUM8Ve/rVr0huVaUpiCuo3JMOjfPLNOMi
hTBLzTAQQpkmSiivTTt4++lNjJKv+sETMB/CRxdlKP5KAYnalMHZ+hN6F2iouHCu
PgqM3ISzWSd+z1bq7P/eGCzP/NynduoLT1MGxe05p1PLzoqDZxUFVHW5Gq3Pu2ji
tOCeYkekuEa6bbJ1pr8CldlfTrNLv5jfNsFPnR8GuDBTme5KBF+3Pzt8kDPiTPFl
SVkA8zpeVuhYAgKS5XTSi6ATTc4fqO3d/GnjINg1TaI6Lx1mVGXzmNdhlGntlH5m
D1lbosiMBdYO7UEsACPXZeNWmfzj2zHCF9vBOO8OvkLIfSWUQu4PGA56bWkc+8Zy
V0Aj59N4mbQkHsatoxsyetHEs/R62xMscqpwOci1i2fq32VGalK+92GspmS80KaC
8VUAUEY2eMUcMmatWI1aHS5aLjqt3JEquzwCySyE/k7QJRa4QT2A0RmErnE5g8Js
m/1ZhYgbLyGxjkugDgzG1zJDOw//Su5HxkArtihqtAS10XvtBN9KcmyDSTEf7N8L
kNJ8Q3OVhV43LIsU4o4PUNJ8LqfcPQVVFgs3g/iYMO378QgYpL2BHce88cf6vrK8
UZRVUVCtwOxa+mAh7/iIVkRy/H6FV/TSwP3UJkzrIbIgOHIIB+d5xPQ5i8MA/MqN
JrF9FqB69D+vYdZLfmST40iMZdVlJm/PlbzBndrRSlfdkc3pAs5w/s6Ia8IpXJj2
JTk9Fd+S+zT7FQ4AFqvLJZLrVvWZ15+xN/39nyvizLhFtNWYQcWgh5BlqmbTGDp6
HZaqSXxiLtgbQws4j2uoq74j4YRqWqOI9fCb7I/OQnpAeyxhz9mA1v1ZwHaehJSH
vHX2VSFRp381I6AZhoDtmzwFOxKUUBFT3EenI9IpCOMUwogo/DGRtY2Pc9Q+FeOu
RDU9UOs+ZhOPmwCy7iVYv7ujrQO2s7FMm8H3ze8okekoJElO1WdSrRLCQAPDWsFS
+06fqzKZDzHYwW0Y3HocJbKii4MyXogoc1vdoDSbTdG1peaApLrTLxWrsCj1S+X/
pHnany7rFc0VZDTJN0aO0dZn24SIguJxQqZ0SG0S8JBKZy/lMyfC040luT0e1ItI
5i7WzbdK6OyHnaFzuP0u6pxH1XTOXUMWzftGNsZWW1bTt+mrRF2vXaD5Bb1E+ltI
m+JBvW8Q6i3jJd6R7I7xXv+NzReU6OE19+1aeh6cTaLQkMafVqYErsUg09qmpPf1
VLW3W6GQD6AUKMI1iQNnldTepNzeycmQrugIrB1PGjgZCA3LPZqpn9j2xYDI4omo
9irrTPARdgTuFQCVqhtRG0PnnSE/zNFCrA4woTvBQT8JoThISnB2E4WQeqVEsIO6
MclTLMQwd2oo9F7baGSR2cxAr07OyhDtiMqtzXGrF8sT+5V0pIv3qdKv87X+9b45
5GIMTbBJigxw3MOmbCzZ23OuaowdzmM8L17C8FdRjOKHDo3cVzUI+7bdrrP8i9yJ
sXjmRNiVS9BmLArO94peiDt2ldH3RKuAwVoqwEAla74zLwinxZBzpa53GmcPgfc3
O5kots1DZlBSg38mRRmN9unkWTfpiLA1+8HJr2F9TgiWovhvLrJTnNEGXkcgS9TU
r9Dl4jilMHISEH6tyCoxjdONPBRDk4mmFdh79O0zgre0LdRUDq/K0zir9sWsqBm/
K5nsQ5/e3btVS+maNSdHaZy6IzHsb/zwnHJL0GuyrZ85hSnOPMfBBGWpPjcGJRZp
WvlRuWykp5MFkLFglTkNDci7VVH2vptfFPo2GV87CdJmlUzXhthmsjyARIl5c/ub
Oo91J3bQNlJFHdCQ8poeKqhC5ISW8j9a6rlmkOaOlIzB6Kj8d6LqW7/+8EE6xD3O
hasQah5bn+il6Jxp0O1n3imDrzEvf5CDiD7hZdp5ehhaDCyMFUIuYHSWgFka/IKX
HWAHBeqp2t8s/mnLFTLy6c6RuxBK7GUP7jdg+ghXejFo6FBPKAzwWWWBKj6I0Dq7
/Bupr7H2o/kRU68h4UqfjRI8hVKOmi0/MLyIQE4g/cGEhedPLvpfqeoWliO2AH1m
tENrH0C13kL/7WaENpJJyRFSLJyhy1LYN+k0CQK0b63CZ+2fsjL8tez1fUeGOnql
Ro3cnJW9Te5eDHJzdCyBfPzyleJD2sPXbavhta21klVdgGyOHtgM7IIdHPebIHvA
2maEsg9G7ykCQLKV4uJs+qP00JQmeAFOTz0F5JduSz/v91jbAIVeRKMtHlP45LXX
15gQvGPLfoTE7QZ14Is3MxrudcO/uQZplWMbdt8CgSniFrddX8/4cQPk+tWw9TGv
cg39600KRhZNMRMbTdCVCSx2EffDB1TKNvlpC0X5CFXzRAGoxyPQlxjSDKtWEslB
2ANvtjJDthxJuWHkVHSL0L2yXes0jXG+v8KSekTN2Sga4gV9S+xfvqtIdgSsI762
yOHCWABHAQrDVi3X1tFY+FcPmZKKlxIL3nQSKXRvY/McsRqEdnGbXUeEsz93x1yy
cuI7k7QNy3QVHlWlnPf4S88g1ie3gP8rpEaPK7C2+WvBpl091av6cJzrdVVOzZc+
AxVgfckCBPl/N+0ksUmz34yd8CfJfhAb5IqkX7bgNVizbIP8gkICHZ89dZ7rgnp4
8GJLi/M7ZFpe1V0gwPyf8tFh/8BHOseWJAn8DQwyBGmiNxIRzOCGCU/+QZRzMXL3
0igRgIghP8MhTWOu3PX4o+s4fkdRVZKsFHHUs+iop1YYiN81+TIpj7cswzm3dHov
mLNlfZxJ0/3L6MktUei6ugXX26mEGMtHbQd7ClnTa1zvD4lWKEKZr3MMSAR7JlQG
2lIjDAXgzvD2vDJOuz5t5RvJXHwDk9cGQ0/mGKEgiEP8QqsrKz89YieJGTk2TWe/
HNTf11pOlX9xZKgVuEAXmjGliPLyvq96C7L6Q5LBlVVIeAaiqH4mPUq5/tVhFt0n
u+y2IclGdsFGRyLk9ixI9xQTdwtN9Z28vZxv3wqCR178D7vDeJ8VJ8MT1+b6vg8h
p6LzhSEXpbfswDl3zuXu//q7a9qsyq/+g3Qtqhxhimsn7NyMYicE2Do2YlFrxJ8i
iBWh4F25lJYwoqR4U9rDwt2yAc/cLq7xF5FvN94npqupYwhI/Myr7w+hQg9mhCAQ
2jHmxuFemCtuyb/ETMs8sMva7gmVlkuc9kFgK82kSTH8m1yOZIyD9vSrPHhF6RcE
XsEMsOf1vbWHSEZ+UrCR2mD0wkvbbURamyQdF07JZCToj1tyMOQD94pheiD6k7QE
/+EFZUexUmOs8F14DO26uxOj3zLmH4gHpNGoS/zfDIFv1OR38My/q7BZvJ4SmltY
IkPhacl08WQhZ8LOKL4KOFpdO7P077qkp7zjJDFkZORCkHZ/M1efqfA/YvYzBEin
CPvp0+lkD8q5g5EnNlpBnPZzFDT5LOv1nVGv6ShZWq6pLwyao5TNykk1c3Z2mr5V
ltM2iv4IKDxnNDoF0XYToo4dy7JP1uLRChn2XDBVTkph0EZeWPN4mf4P3+F9u/e6
hn+ie1J0yvW/bCNy5nX1Uu3XYVGQ7RctE6ZAlg8xHghyyaeEgeR7pKaCovMIMbGe
3/oKXWKQ2eK2eJXI5Dajo1g//tCWO055RyB8Hl0e0JBAkbjSr+MBXSAZNpeMBvDV
YRboU/0d42ihdR0WS+IC9YObrfz3BeByb4DePki2GNaFF/fYx/0iOw51g8vuRfhx
JT43WRKckb6nRsW+9zy0bLIzbIr/wBhltXv4/9nbQgDi9D/khZIYmXDdwk9CXYrd
j7icIdyIJgFfNNFaWSMj0fDhXwPEfT6sgTchbUsTWA6rOdIUHyQqbKqis0pFHCgE
/VU57UM2B9QfVnCEocXZe9d/m57EEsr6MzGMXRH11FxhIjr65Y9M2fztL521TJxD
qllgIW3GkVJ38fZerYx+qFxyYuv4R2Bq7wkTMLPWvoWRuuDaJsJVxYu4eD6lwn5k
fUib/ipUHBobFMprdFnIoizj0hgABEYaafRmnISH7dn7fdN9TP8nPg8sxGR7eGNf
`protect END_PROTECTED
