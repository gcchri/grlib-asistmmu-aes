`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dSfZMtJA6GXlK8Qf2oZNCzu7kb//PkuNOzJOAMGRpa/aEmqOOrWCpcXzaRwL4CYe
4zx2aEKzpgcjCJxI5MCKX4ymBSMuGa+tIei7WfxYBMUyiIDOkukG4EiRMsap4nXl
1A4405gJYb9uet18vaUIeUZSjl01c3hSRlb8ZIrdzKMUhEHUq/qFgYzUMm5jEmOc
6miAzVNovDa4Jw4zogaY5H2Raoi9yJ3AdBtCIQ5V2TAnSyR9cRYLB3Dt2yknanYV
UFW39fDJYEOyBtWIYZ7wYdR2J2v8mu8aHl+KSmOvLx3RHEtPGqQk8X4NbhZBq9Fb
lo5V8NTRNwF3CBVUytlw8qi+U43sFaEMiRHYO20gMF3ts2d9Ap9HNDJe+ePWYykL
FIJTgl7Y/HnNKUhbFMAprA==
`protect END_PROTECTED
