`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/GK3r3cD+SGzr2K+jLVLCLMk/Zc4RAwkkb8cyBmGRKWQvNpl6bfTkuEfExk/a1HP
O2sy+IFBZ1L0WT3JpVgKAt8STnw9pCFdYIJ+mHPfixDoQA65jK5i2gQvE6lR7BEN
Tel+Ad5FOgJKkLWeaTDBXLbyutkND0AcUaX9AW+GujsPPAyBZbIgtb51+rUwuny6
gG3UT9vb7u4391Nma7BZQAfXZ+L4ibzdYuGSGrJU8f4gvriysthKFNVTlOxZxOaO
2Is0ebi0ByKL+Efdmuv/WxRKyS2NjewUjiI76NfoqGc=
`protect END_PROTECTED
