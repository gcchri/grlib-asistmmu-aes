`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGyiuEbjsheKZj0OlIFvWtSL04pj2IcslZ8L/JzxqwMHy5GgGvgMAie0B53vAFIp
W71D5b8Nd9edRrbvYKlJGX6bUvyfG0ly0iQ5gbwh0XaK5fLqb/w/++H2oMkUtI7A
HONaT5b4QQGixBtdIDUULHJiu9TkFL37JP41/jxh9BmiB4yWz4oDcp9D8fhrV7v6
dX0APxrfy0a/Yf4/Rr7F4HPvpSX9Yshso06Fi/TDvUwRFihHi/QTpgpVbcvXSLlT
F08tW6FXX7s82woaqqxbTWOHFbyzqUrzlxUc3yCD/m8QhDKhU/S/5i275PwLQnbf
Mq/JJqk1jHsApCN+A/ZaUom1nLnJ7qTL7YZ05Kyg3lL5Tix5y3JjYOxnOfBJg5qJ
eIKxgT1h2CXlQ2S5YPPrHuBj8TTh9uYhrxrm3vs6ZkQT62hrv4ulH4IhTf0mMiuC
`protect END_PROTECTED
