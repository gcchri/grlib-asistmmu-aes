`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yyp/uWbh58lJGvq0ETjgGW5hmr64i2R24pJRMXDf5dUWzEqNyV3DbwoihvH+HUNC
aoFIj2eLKfbCIcgEngE7fj8zQMPxximBdPlVJgzfkUlJBmV9Ovo3grtqkf1CwP3F
GGf8Al7sOb3Ga7Bv5+wxMmZdpqY/s2Pb6SGV5HWRgirD3ZT/Te2P6a02c2wgMaaC
L+ExXZUUp9cbVZs2n9xYhDgkQaptjhSuUaU+kd66rjAjoJI78CuVuILyno76VMbm
yDlSQrbt46H8fS79E0bZs2C2/wjfYxpEkKhZtcfxjX/W+DS6SIOQ1xlcOLOjeYSS
hMh99lPaFEPB18Dm66SlS5dm6cZ6f8tOGwOTry2W1UImYmiXBnvVpGmkzJxHNcyB
u8199c6F+dVbH6NNXjCf8g6SQn+eas+UZ1lT0uh/2z//24mb5cW7/4JP2wgUSeN0
z0s20lszyd6w4t1vndxozeXh1IirIILYngGP6980qtFeR24cQQQpcbm3a4FeNHrf
H9chyjLcFxXpElbJxurxMIOe6Zhd9MLUG27DoKFw+QstTF/xIrrBhimRNIl89REX
eXsxmZ3dFh04YvkhZMFAdHLlbeYge+9pyzRTDhA8ivHRU/N6pXhqjcZ7+RR0wWUf
`protect END_PROTECTED
