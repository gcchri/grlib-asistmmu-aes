`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5uX7Gi8FbX+Fx/LvL/K2FOmQX6QFpKC2lnZScQTwCHFH1IY/rOmQE84/xQ4fsYOx
SpH8nMAGu3sR0hylULtLlH42LpufaVet+0KCl60baBLpqFtnw+rxDgqaG7N3GyuB
O7z485VhMAJHPjioLCQhOva1/g177KXmIyUy7WVIbVyWZ5LKOc7nlVPgtEdjKTOY
UQMcklDzKvMOnbw4NtoCt5/OMpP1c4Z/cuz5f7nZhm8TUbHXqsqTbKEvKqigF89/
D/zexLAd/VX6WseuEqA7atRXvRyknLZwUZpCxj1v3x4U2JVBYOXukMn3V6ORaFXj
xeQHa6HEIoeTDu8DAvKOyQ==
`protect END_PROTECTED
