`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1bmdrvvUt/qb7QiaRgPRl18rke4GV0fVCsfCMUZNTqhRVJhJhRbu58zk5nL1mty
69HKkGZZs06fa2ULPOr8PlRjszranZDzRlpM9HaHmMGHrEx9XREK9rE4uI8z1gg8
WE0G6tFlVI8+AjCpvl7esL9+unIKz4l7W6g5uVL5AS0Bo3/5Dd6ZAFXhjSO8pyHT
Juy2nMwx5SOeQBmC7G8JfhyRbcoawrZxSwGZgAHTxkN5HO5bYvbPLnLZ8JumfPhj
ehTj4X2P10PmfFF9/gnMCqbvejh0AWagLQC15QehC2a4vWcD9+1EP4W8mV5omUuH
2uFb/qG106hAEwCgnGEkXorGYMLZF7S9NBUN5Wfx7O+BvX12/e+ks22EvMtq/1LL
6D8Rr9KQ9Q4qnuPCW0lVgpS5o1fLN5We4/xkDJDBbIwksbUmFCMxTA16IDTZFvSQ
`protect END_PROTECTED
