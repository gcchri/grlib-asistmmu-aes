`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t956PuPZpKEYIDWzzaD9c3wYA7i0gWYLyUaoqqJWbjVuLtxNcPsm+DjTXIU9gzmJ
zNUvkc81ER2RSDGHeCroUp+9UOaOtPvY1nLnqtgaloyMkRmWjZ6BIuCDB+jWpqbS
gUIwp+tZeWE9Y08Iqb59Xis3hRYvf5dHJxPWNAt3st8nzD0XfKKbNq6BB1jBwKPo
EhkN6iUrG9HqhCOvq4UPHfvqrh5xawVTJNFWQw+REoHqTbcAhNqro2ii1rsTckIc
sI8bLCaBc2+b40Gw17gx/QEqDie0wiw2iHQLwb1KRvfitzlKxJQwL1XPHYLQuub8
MAFisLYdbPLGYyT/O8IhyQsJDpqtSHOs3mdVJ9hgcRpyLOUoLPxzhyKMrVmfhywL
+vu2i5NhxVhEq3SNgzY3WqGrX3MPVe2jn5HlpPPHZ/oQV4hlCwnuIw9PNvBDpuHb
R3NjyIugAwvhQGm0BlR8ZOerJ8TjPS16KPYsWQtwHXOwvqQbgWB06BrYmpMOvHR6
fofJ9QvcoK4vJoumcXCJ1GYHuPWMsx8pp+1rv5YKOtfNIMXSvtTR0cCsnTu3u5EP
BMOoqnSP2xJPj+/qlMDzuTu03NReOVWRpvTglGZ3L3b7k75e2iQU1M6OHlBP3L77
anZ6ske1WBytnDYk6Gou9FzjVjna0UeyPTv2axUbo1IZPwMXMSORoDjcwaSH7TFR
Xh/gnz0w3Ja9jMCVYOEkQjBv6MnfxrfG32R1wFU+3phuuqiKmJV2cYSwdmdiE/ax
XFnn12ikJy3pJFWz9eZzSmdeGSRzLC9Qf7pw1+eSz/O/ZRfEgLcAocIUjnyg8/hA
`protect END_PROTECTED
