`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDfLZae2yGpIf9vFYAxGMYJE/9vbTk262kYfqQtsTjy0u5UvjIXfOBo4PpgTyIrQ
iWsxGaPxt6oOztxiFThfGQCKlRfn6/w5s/Prs1pZe2rTQaP9xhZPIkX2klROIVyr
CKdVrriyICEzDxQDa/eGE5lxf8UUn+bhSQV4UMTE8rK9in0oC/X0/JYXcDwV7ZCJ
u89bHaQ974ENshw99t9NQ0UlpKHjCS+N8FRGM5knHWepzivtrGqo7H4Add+LUJvz
VeHPUEnIXGgj9+xsKfl1wWAN3ArlDTbquDn9flCTuRsr6RiaWGUBAsiqccROqlnL
cCbonX23BEfMev3S4IDiu8FWSZEs68oSNArpBjqPUUiQrH2FF2n8ue9LzMNT0CEd
hiZmMM4LzNXKQQe/5Ej0vlB3G+TZMjKNvKA++kfwJRKZmNCu6XteKWDGL8uumjlh
OsE/6c1oky8fnPz2ksSD/psYByGxxATcqJu2rWOyrefPFN84LfMid3dyEnygMose
mKh9iEYKpVTOFBa7/XOmO+TXlgzBqlDyniE8yJznmKwp2vGlJ+l68FB6eovN52Rt
xYoUkqgdTaaBGuTmKTZzOo4roo+MaYwXnUc9fZRP4loARRSWVXUSDHwwe+0aRXac
4flKjsttD92q9uJwqjs8ZcQscL+w//FHhq2irPLrTJLRCWuR8QrRwBhFzK2bNQB/
bZQBPi+L4ipiWYU9egjClVU9+2bjlI3pFFVQqhQBzfOaYkdsDyBMB8QTiWd/egL7
HnltwBeGzUx44faOzRjXVBfB27ozrKv2F33vhSHqi0fT+PqWNxQGUpAZQYZ/xuvK
VJlPxRpEZiol+MwLiwgdYQ==
`protect END_PROTECTED
