`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ecq3ElKu598+EpU9JNthz0CSC44lfNiAl/5OQagZ+FQo7gaZiI5c7y0WoOIwZ8/F
bedAUS+94U6kG/uNU3Xj7WDsac2FmAZbK2MOn4zdHdQVRTYu6dKNZRnXPx8KRIgp
yx6L5dScIzNLF8ahN3vuTY4kroXiCmblilL/qaQ6CxaZknqwo6GPq2YQqstTzja8
YHn3hrz9twBdrfesUq9qxJwNVVUo8Wlmci3/UA7xXrm2cGaJ1TFs30WRBv+HeZrL
yQriXsowoGHeqjknr2DK6UGqFC9dVzgx4twMGBEDWXqp2U7ikWYEoIj+9WIw5dla
iZUFzSoU0w8+hzpjHzbqqPfZGn5h4+VdiiNIYNVQ/C3dmr0Y/ycJk9v9MLMCshq0
T4XI45Mfgbiht7cD//C4AyeGAikm5AArvL5+UZduDPj7/fuOPGVQqQ4KQxVNGkVN
KEWGEU52KScPtLVpmyV5J/4e6KnbmRd/paTmvYR5WHgmawTLR3AXrgvEam19arTC
lH2PVFRfs9F5qRWEwDUL+j0L9d8/1cJL0/RR1MFDCMBBuzSgkvaAyP4koUVAHyHp
IDMaVTw7KCYr24ahc+hz188ZhMo1ErRDivnyGebrl4hRozmPqHSzSiOYO0MC5+n5
iDxHHGL8nNmlO/67YMFHRRZ4vSudcHSgxl/3YA5KMYnjrbqw6hlVtdQ7U5E30YJN
FatstPsHfx1RG44/Qf8bR5aJ9YDsj4d/Z0K7bc2R7GcVo/prhr+xAPCqSw6pdrFk
n4daHvHSR44vmSybLs4icu6NMiAhICr2IUv+7eisyP4JK25yt+mBB2W5nPakLyrd
Owko6Hr0Ex9yj+uZ/7rv065GL+ut1NQ6PNeNnTepvheqH28Ug0g/Jr1wqP2VxFFg
3M2/9gj+2Fy0RGZX4o/RZjAHGg/DLZRaTW9qZwxUJLn7bLCiTd9eioKm362h8aEM
pDF9UrGuAcnBCu4UIOlyaESnoLrtM6w56OE2/T8BX3Vor6M3p3djwLyLNM81CBiv
L+nXHtRdxZjOIEPRKcBSs2Cfkd/+DuXw0vr5B4Bff+KfEja9EKt+ioUtwi5dW85b
PGfWXYmJZ6TKvx9igdGjfVyxxE40P/9qTGhHadW2tKR/7hK5dc4KeLXnsz0v7y3v
6eOYmz5JiLi0+vc5Fm5hPsRoWMuH97R3Em5hosFCFuCjsRxL30jDrnw/ERvzHEzz
sfbVApGChHes9nPiD4tuQZ1BBTdejr2BlcPQ+2hOdbjIG/vmZPCoJWWY2Tv2givy
AXps572YUot3EMQ3PxqsKrfN9l4u+SUqF7oiFXNCgCPA4+U7axM2bO3ToxMIQGn4
khWwmF9pwUOj7gzz0vwVMpf1pzUoOrzsg0WVmPiB0ZG9DDGXDEm+WgKjOYcQEkHO
zpAsujxAQWg564zOjvWzPHt53U8o51vgTHn53Dg5WYgH3EAJnt/1lmK4PAfuOT6m
`protect END_PROTECTED
