`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7W9Mf7xpVGhE5ZlWyQ8AlFMa3mLPp7XRau48kqG4LyhzUtbh751xtP4KXWCYbDm
vooDfdyfX6Vtj8/62hunxzUhrKPTTnftns+36LvKWrlWddj4cSoU1kaYVQW5Ligy
uEYw13SlPn4jRHjqZcM/oFrbpcMcmy2bWFl8QwaeMIJf+vkjmawJPI8dXSfEz0nc
0GPXIZvdygaxZ/LAyOAaRyMy3xxShjlg0X2UvFCW1hcAgBBx+Isn04JB6uuH0dx0
LY2uwtNlc7QLfSYqVhqQd/X1kinbsfZh/YXQ6TfADutDkkBiiic8sDT2Mn59wx4F
skTyoc1/HG820LjgeJ6CnWS5AdiSy7lbr9ZDNTouqVSNH1ACsSHHhqBAnNxNxYD8
exSGl+xSLFVRJQmovCNoqDZ6cL/lm8We1Gy0Ce7DdnpDR0OBoSzagsg6QhPWvVhw
VYzxhQKlbr2r7rX4i7ZJS+dVMtwS52M4HNeZRROVFBk=
`protect END_PROTECTED
