`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y0915awdHH0MbWq6txdMSAz6FUq98nkhBvTfbjoQaE9Nxl3rjuQZvRXMnJSrpIQ0
AvUj6XFhgrA2/RNFyRjc31KhTXaEt1/Oh0yIPsu6h0li3rWj5NYkpUz/GO7qrbwn
yioc1nf8JM25ceuQId0zooF0rlcwTzAPDlUax090Rw5+kIwppmNZueCE2ov73fsp
rde4jYpBvhcLsZyf6cFY+lVMhVRcEQVYcRfrmhKe6+PSQ+LmSgFuwRTt6z+rqjJx
yZnl8q60FoW1aDevA6bVh1foyMl6GHXEuNyvCXjNATFq3NnLIb4p4tChFhATMKBn
yzvbvYr2Hmo9HjAoSlfaEnFZtxrZnlDAar9rUKs+i/ROG/9/FLH+/Jdq5cC4G3tt
AJ8sPhza55A58MW4qN6dsyibScOD2C5fWLHpVLTeI76A0Ciy5DpioL5ehUVMKUT8
vejVEmtdqfsYCETh7iqu3YOV1wx7Zhg2E4Njw6QqCSo63kBqwvBmKfWplPV27xKe
wTGP/cv2N5Qsk5xIJMgWjofoYoNiXjwLO1TfKJsJKeQ=
`protect END_PROTECTED
