`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cK5eacVkXAX8PXXnhP++65GgrcMJZWETP65UJ9bROBTw25R+6Ix3yijVO2daAS2P
gbtv8eSQl1dsq7fPraDUG/CoqSL0G6JaXHF7rDG+t3PLZG2zB5ZMlv/JQ0bd6Kmy
2HCgyidNov/eaa9A+T1rrGnYPVJ6iJLMxYM6fi3aEV+lgnzv0Rz1sRnfhCUu9mv+
ETMEeXLsHHuwPCt002LYD6Ot2MNyabg2yVC/T4zDFvPN6SNEwWeqKgH5VgHTIjQZ
xIC/5/B2l/yWgqLDfzz7jsMEwhHewJiKZsxlOaPNWFwqiQ/TnsplIoTIT7WeKyXk
B+eYVBlugObb5FWM/sudpidaStFpN5vdDjyYr0e01KwnLcCloLnJJBjLUB3tYCbb
v2QrkZMvwK9vkAUhbQ3eAheNVdjaveJfKePVYsiK8II5fF6NrIg693wiFk7vubN/
SjOgBNtbv+AO1wlij16IiXX8FTvDoUWmU+kpD19lEe5Wgcsk66yt82JOPR09iKpi
sS57RZaPwkbvXuEqta/6aZRTIbn+OPt2YjP9OcC4gcE=
`protect END_PROTECTED
