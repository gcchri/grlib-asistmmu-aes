`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frb2qUwEmMTPmvSJYar6QfEM9dR4R4fcR+nhdTxJOisVW8k9iZVoP/hMWoYKu9Hc
XFtyfIH1UmqdgV9VxcAyE9b6xpsWYatjqD1j+nZ+Us564Qig7XF2j0ZFbij4t5uJ
094UJUa4BkiTVEMixpzpTFxBd5vBGKC/VTLJ8B7JvoLukf2pufIz5IWiGcaxtAIx
G1HiEt/sIPOyh+C3mkDhSUNPkd4fyBwsyFlG3wpWfqOhA+F+t8QU/fp9UQip1jN7
PdP7pd2aLyaSGeVQgcFVs1IqzwS1N7R7r+l/qtPF3WIx5ozGqNeZpr5m/dy2h5jU
qKwaxCBCRdy03DAZn1mUHpS2O2PJtTMcIaEBoGCp3XXB4OE3HDBguXY870dhwwAI
wOSqS16Fa44WtBbF9++b9jaLhxUMRUKHw7HiKftZ/jAORSNUgHoEgZUTqK7jP9so
hFZq4dA3RY8wQZ6hOVPaxdPm0u8zoFjIQe6sNz7a84c=
`protect END_PROTECTED
