`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GtDepCYocISENqL2wo70Aep5ITB56vqo6EccnsOSWIgJzJa+58Q6yAkJPagXw4ds
DiIMMEXHvG7oew3vsR+7eWD1hX19y6NeZCGr48OK41c0jk3lz1OaEhCXDIVl9YHM
dg1jYvSG3ZyHEkciTH7c0uMhdU5FT1j6Uj/gOFH8Vz0cz7+0Ee4naiwukm3pI9Eg
ztkdLt+DOrn2fX3Xg6Qk/xizEMEbKb7zz+kX/CAbgUefR6oHSMCfu61LJCiyz22P
`protect END_PROTECTED
