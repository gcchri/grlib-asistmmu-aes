`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NpjU3NTL23aVS57fXrZSYpXfq6wu4F+XaB1J++oNJQwSGJ6XR+2cibTwIMbV7hjX
q63smPIsH3KDWoQxnRcJ+LjKjBu5KGAxcE6cAwZKKiqhBi8As2PeMSVMZe24INIx
Xv0H0OSXlq21CUaMAMFOsWv0+fv1nV2FNIvlZ1hLH/o4tIzZDwmAcoAbUuVVWOvc
niskbVlHwAu910gbMkHgeMeGbew+yA6PqfVO5jggMnHqMSjlC2ZyZqc8UCGAcZFb
+l2/92DRNEvuSiXlyvolZthhvHGf6TcyvkgxamG1VS0wZ64DAg6fzc8f0TB3W3Ji
sff4Su7MpoKyUHSi6f7L3oB2LI1bQqc9arLL4AliIAVxsO/dFILrPj+cka1ArTVP
rAIPc0pHxdmPJ4SqLoT7IhL9+1TZcL1QfnQWrw83QD51bHFKXUYYOq2ls7hTrGCj
6yCfvO97Zn4rYYwL/j9SPA==
`protect END_PROTECTED
