`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IdpRszIK/VQ/mcrYngc5FLdOt1G9WEHjWipCS9oTtOPT9sXsBOZUC4jLmBJ84WsY
HdtyhdohstKJS9K1f3uEVU1wOiWSmSifheq4GmsbkG8h/UJcPPjBNk5/ar6d5fCI
eDsrvvNsywTWGlek5t1vnkEm6e41bnzRvKp6bmi3xVdYpOwMKaT56tZuYqehpczV
t6crRpuI7xMeLZJdvwa+JfSSzmwKlW6KEqrXF+2Upn6k803pzqlyyhGBooR1+NmW
rShNwfrA53mIKnpHScC79MonQCqtlbToFuSKK2Ab2/DKWHPewn4PbhX923tRFOUJ
e/2aw5yMlV4xXACd1ELGE20GTQuJjzk4gu3rnZHqqD4j9cW1k61m43fKlkBAPoBl
gl6hip2IaVsOuvmqmpbm6PDyufBNewqgDLxUyxVgI4vSVZF8JY+pxpaIOHIg5g71
u0KvRzV2Yhrpoc4pqeoGAx03tidRTmdegSKch8qR5nttLU/SrF61McrFzE3bBAUU
NoHlprxFBItEY/Grqfxfc/adDarlHwgLAJtwHt2m79HC2gEAzlCZ+x2ic0EQsdwc
`protect END_PROTECTED
