`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bkeb2dRPzpiVouYiJ/oIPKht4p+RIgZ4hImRgsK0pbZRgFucL0k5qHgdC9lHS8uI
7YAKABaeVgGEuOMwq2L1ZobGA2y7DfgAvK+y4MjAKuxtqBN1cl7TS+7OJhW1ZdNJ
F+QcWM4LCqLmUQUKMnvfAeE5UWqT7gPiqCn2kWz+/Vd998lF75n+tWGnvJcfyqwl
3xIzI/TxTasz2r7aKdCsQKzCM/gU91C/FpQrqkoIai/yQ2CqtK5dBf526u5/9jyT
P1+Uv2ADlB6riEsjA6rhtzrgkmr94fCKRi6+3sjcP91s8yMFPw72W9c7JK1iR2kQ
0jWD1YiaNTIbZppCE9aOlqeSvFxEilPO7kLC9V/t18UNUOGKxIDl63BETqzM49xd
zlwzshiUFqy2ucm2Ox+teotaH9LjGfGz5uWmKPlDEin6mkyJJtlwVNZE08PoYig0
GxyZ57liNc7f2ZmSrCb3eWeH0ScbxUOvY5KLSJaebYmmH5WPcFwYcW3U+Lzf1NL0
eDMNH6adwX8eRywO+T3Yx2o0j3JrLCQgY5Ze5z0mlg1m7cd43oNTB04UGPx+XYwt
yj3X1hEMK5IaargGV8qA9O/48OT0yFXky7AQJtQu1+84YggJy1gginZABPNNmzbe
dfiLbQ+hCaWReeD34GGf7JkuoeYJR4xayO5ODos+ncqeiQe24qEWbr0xI9FHtZ8a
UpUAhgRbx9H/gBa6IrazlMT/PkJvSaj3Y8Ta8pXsmP24x8J7lWuKCH9IhmVtO9v/
810HiL+RMvglfMqJPlPibzMVbTxSGIQykC9wmUCACtkIhgKZfi0aT8Zms7zS1Kh7
SHMuLt7GFrzb+LIJUF7w0YMf7XtfXVaJK/hq/zSTJhQxFs89xZN0KH3FHZh62o7c
/nySnixVB3Yh+4OyxPjTjZJXoJ5yNq33SlfDc3exLZTQ/2F9HhXCapuPjWagYJY4
QZ16p9qBIN1l+3BNWRwIUt7oSR75JLOjUL/7HaxFIfLjS/XtKeVHcHV+p571fB2X
YjZFtd35YVVwI97UWs9+jicmFO+tPGWZz+Ays3czGFCH/T83eKMH1f6GyY43fT3m
tzvA+TONDu/3qkUjDBbhIM++Vzkf3yU20d/dHVYNhPS2b4tzKmYOTdP01zYV7F6D
UbmxGWhxhTeJZ8QmS4MVSB5VwlMRRHvoYZhLiPuWvOm2QvOykhb4M4z+9Jy4xJFD
kUhANRYzyFHBMslEcvnvUej5oH7Oy7QoFu1bDxMX4izVGOxGpA7+lGIguJ6f196F
ly1EBxwykRtMeTeyM7SGmP8lgYP/pyEBUpfZSPZS44xme/sRx9P/j+hqZVdZVakD
XfmulciTyDPxVdhoNbitepAa0w+R26gat2t6SiP+MRavl0mMuapTV8RFAanFPxml
jZLIiplJXb/pHsMnButrPYITEuegCB6FvjdkYSeUqczxXAZzl2m+uJ2x4HyyaIln
DeIEX5xfAlqZH8ykTbpJ9Vrh+jHLyjpDpkI2/zwkjfKZ/pnAfF9Wo8dQftVZrWSq
KKggANttCHKFHNt2LVy4H+F4q2uzUA7VwE1xDrxITJYbg9VbOx9iyUAsOAIePZ+J
h3TWDE4+O8NDM5pKzdP5Vp5Af7OHBtg2IIkSaov9sSLbf6Io4qT4LzLJs6GWvh0f
ASu0v67WdHKK71RarRxOwlVd1L4rY4FrBde2T21tE95ByCXWeQKdjo4n4NrXIE5C
+mXLAFUNUDiSpjrHhvRwkBpY/4xsoFzBJwZjv0uE2HLTmRYHoppHokH83Adkj4Rt
KdU+qlrzsU+u/+KlsCrXCVulpL9RVJ0U2hxAoTKuKkhbOJFRXeybpsseCcTCEcok
761+SrMADbQoRS+A0mqW+LQrf6MG+1kOvNL5FPd/ymeRHMJDrgi9qswvVRt/mMAA
g7JsLFuHWLtTWMYcB/KA4rpACCz2prUiYatXjVQJQ1IHe1wTzOI423D2FMxAKyoe
NoC9EJ8EfLBcz0m1MLQw5R7/OPhZ7bviIQoYXk2FfRuFTmojB8I5e7BLdSwqRXnV
9CgYg3q0TccZQil0dOl7jMbXhqPsvQwplJP2bc0cXKWU8PyrLoliOQiQPQZ22Qw0
YEKAXA7rim+y6LsWaO7GlxypOSUcVFIpAe42B6IhrA1U6Osmvv1ZHXJdQgadkW31
8D6xQBDwSr2x4w6FAXarJsdhh7ATnvbIfMVnAmoW2Y3hcaebCbKDq38oD9aBWbJP
F+8bNx/oqK7jKuLTgy/OJwY4WE9DCm2FC6T8eCYfjAS91/e593meoBFTo+2XPQAx
SnLhBqT4VLnkKjP4SYvzWaVjloyZfRIwFgHrSkRPDOqhDwxk5b1Yhs/3SOWnpevg
CmRyMA/u3nPSoHzYgDpQ1YYGtELMhzHrpnD7lGQQcndQLgQ38HPUxPcGV/NmAuRf
LgJ9NMN5YH/QlJAgD8LEfq3B+/ZHbeOGMDtuJRVRmp5ElRrhSd8dW1FOVgaxs0Pw
Uwt5FdFSqLdJ3l/5TVnR9CgB0+KcLLwqwNSOM11GnFtPPF1T421+wUHlxQxEaIpb
36Di7C9e8rNBStPpZVGBlNIFKKI/LTCyL1mIPCuAkby4Ne8H2dTXAu7ccmMLVF//
V/vU5fTcatKALHq18L8IetQIZ2WmPFzXe20qdoKYr4UgsSlUv2T48d7UYKXmLLvb
tTBIad/ePdS2GvaveMoIwBDWP9A6yikdTxOBPM4vUBOmVEDTnRsDOXeDvY0/nI+z
kx+2qmeZYNR5aIbnEebIlIhXtBzlhy+ga1z68smENGDM8r/0VUFSp67m64+qD6m0
lstQ7K6licBw7rTVDM5m2JwBEdES3p9gre4hNSDRRSaY6AduDdY712DE8Rh5XoBI
XoyHFHqtKClhc0OsJ4ZQnVX3uF16O5SKUM/D9dljtf07iMSGPlR8ym2ydsnnzzTx
mUvP6kuPIY1nx1ZL0yhdStJf5dsbjCKXN8QT2XfnuCtwDo8cpL7gSWbg/LQbuKHB
A0MysrfftqcKU4D/uoOcegp/NarbEAcioKH7/855FKhUvv6fvsSz5HlYyWIR7i/l
9TjyDC5EZ5/WzHDKjBXdnx3qWZE+PdWez4+OeDLFlvrGr/ZhYwUWt0QyXK+/zjVt
j2ZV4LmumBfeaZnapio89kpNG6wGzoD44h0lQDJaAJUYPKJGn/QljAvOGy9rX7Cr
Ww8b1eqfMiQux4zF3uKIxYBJyjjVBZ05oY0N5cd41QUhgl4Lng9c+4qSN9Dypbvr
aAvHPvQbyE5KhqEAiBtpAf++EBZWXW0JeOzVnE08dWpZSg24uYnqTS/hHOEn8S6Z
btAuQHMsMNgiMto6Mb0oLZZShMFviQx4p1wS5qdrqFh8pzWWaqiicWGPZzFWEOuS
zhlDYfJS37cJDprB2plm+aYBslqRZ9ssBq6d6BQ8L4xO4rknhg+RmYkzcMuYYV59
PW/T+WmYxP2cYNVCoe+Fm1srN/n2NMdSk0BTN+2CSpBDmZlVmBQrjVdAoShw1jV0
IuinNolxaZG0xO1bgBiBgjxDSf8pcz/BJhvChwuuqPpq1VCPtYHZW5H84tG7HP0i
SjEnEq32zrP4iSrWLP/zQOe9UC2zUaU9aDumkVQgk72/azD8gSsUsyzdasjI5TxJ
yauJrcP5N/A3WxFSC9YCgQMJs4RIhv91T7ZTc+ZD6nrXvW7ylfhjCoAQrZ/fStYd
XJn2fFeE4Bo9J6u+bbWNieReHnGpZ90I21qdPV52Yd+UgkewO+IlDAqAvtp8bRn3
QVXxspR4hWy8hAu3pZXGwFFC+Z+HynZgR90crNW5GoY=
`protect END_PROTECTED
