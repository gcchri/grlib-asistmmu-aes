`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SzS5bt/Gq4EYk6O2WRJ8Tru+b6Zw3zSBrzUifHT7EtCH9KnU+8QKlpa3ESmZ7j1S
dhMkvfcr1+hElVL8ydGwjqRHFC1vSzam+xXPB9H695Y/TG4QAstOiPiImBy7JUwk
aX7bfJqHCpQnLda6S5V1EG+ZYAL9Yjle+0CXjWxvHEwOQ1mChQyba7KFneKGG/8O
lYW6DVpc0pGNmxMTX5T+u+aTraP0L0YUQz9gLAnx2p3leZ8V6VYzLta9g6tlknxV
8UK3OFioeuDGSz+90GhdrAuVHyioM8/maX9geHfZSa/gbUbKZcPLeglBbYcxE4ms
x5eSXa/f0bWFZObFBfEqC+VVYZFQTcYhPzb0repxT1Gl1kdFhC5kz4X4SsjYvr+u
w1ahEMMR00QqnXS1/gHMC7mGWub70HEz8sZZTE49+KnoifwlEl8dLOWiX28Ra7QD
HV1BcjTXIHopNSQP9AU2nLOKWkq4CR2Ieo6lUM623uUCsXo3m8wvYfo/4Kdgfgze
nCPlrOqx/W/Nvcw15bngvx+GtjF1aZX0BweoPnBMEvm8YyiYVBLuIe60mf2uEkH2
4wUm3rKvuAcbOAIXYMGuxswBA8VdfDUB8k74yMtVS1mDsZZ11UXnRDPVMt0x/aVu
Wpqe6Aq39k2dbE9AM1ig3ezS2w+oqbrH5ZuFLSBGDXhS7n8cOBeOXUA2GoYLA2kG
qZo9j82M+v+xrrMgK8CQevyIlh7crXlSFmX5DYYzoDnrnfP9k73whCvUCu0hZ8vo
N5CuM5bzuUvvNrFdIIFuZpJbP8q+hdNHUUxHu61TewnHV/OYhgfduAptw+OGUhek
fytEWeBh81vnpVCZzsHj+U49/6i2FhpADEpPC03XxIkbZpOo/ehNfykatInvNLBk
MgRWI+t3qqvAr63mUYt7fB7BAb/gPzNkmB1EAt0CNlR/e4CnXhZWbVBbcNOI9421
KvjTs4i8pUPYdwUeaQqTkWKGItDW2GkOvPl4S7MOklUlJZXOS7Tq/JIDJUQr2e21
YTPBDhWOYBuzRtP8nZdgLz+046F3ktHfKznf4MBvYWsxaSXqE2yH5ZRpxhkVXw71
14jaz0GyAkFsKFVbL/1Yg8edz42REm0Lo+gfm+KO6hYm7rCKRrnOc6fEA4HPx9cE
IvI9yO4U39C2Y9I1pjAd4juY2OQhMH13TizPPklFZeMoMacYPoB2Gsmc4fGQuC1K
/drQXPWNu4QMn4vC2/PduuK/Cow4ILc8n22N8pPmGdWh20AoSaAmiRjVhBBeOMs4
G1KOrIeF6fVKyKooYGK5AdnoDMAmlQhL1v84eCfV7/JS6D91vM6nSSbmZtQFehZX
oQ09Ux6tei2oTfY/zHf0RQWbuF1VT+bw3c0z5zEFrZE/8jWMTSakUqPH7gFwdULT
jd1BOffxZ2VBTXW05HLYotmuoUnHug+k8jy/XLMJL61qn71iXmCndktlhjMChqYK
5bELuSIVYOiQtUO8gTNANYCnSHqWT8zhYJ4bWESivYSdHIbemUNIr4mRkP3LQFG/
ZxOQnOgwI0DijxNWra2cpRbFYl6pLTi02SzKGEXqsz6Dt55NfO/tt1Z04hifef6T
injU9bIToOaVC8GzFbdL0NEhdHz/qgqyrzsARIZ3fuPwFu0jH6AKo6TTgKe43kku
cBbjcElNG6O2CXtlXdLgCFp1uUwXaWvP1zyIosi4klCoVymJZb+dkALvyxLFtIK1
vnmJAdtpwMzlpD9iCkz+iZPaOlkXtneTkVE0UCLc0LpiYCxZwSfVAo1OHnupvBuA
Rg7aEL/qUMEXIzZT8e+Ev4jwghtL/wDxNtS9oFB3v4Yzfx8i7yh01ScElLNrOkoi
pU4Jt1dCeXSwrpdt19tbgaII447c3lNXpKXjDea8O8V8A7uuiIcZPFpzHhQ3YcpW
jzCDPqKClT5EUtBt8UJw7C2h2XYE/3OYRqAO5qIK5dT2JX2+dw7QfZjyysJSH0s8
6qw6a/CvrMZUcU/UCx8kwcibLdDnZJpBnk908sWIh289eoH1R3oiXrol5ZSf6uaj
MXTPQ77XbaAf4ak/0tpvSzlfiw6pqbuK2w9mBw2z/vt+QwzBGcwVNpHxQgRIFtU1
jXjrlIgPs5q7AymigKPpSEXgoB+zFId0CSnx2thEmX4fPefqVhEdAlKXx8sljPLe
4bF15lVz/YDFdc+6y2f8c+8FmABAlUbbHckYILOqjzzNSXBJmT5MeUT3OKUQTaAV
4UpXKYB+XQa+6j0jQT3VMTpayVjVINLyjWP52Lgyxh4hWAefZAILLNnKojQpLIRS
6lMCK9tPCl5LfFJe1iEn9emRcvm+Mo8EdIBbdipUL9lNay4kHv0lJdYbxkCgLHhx
QFuQDWGwP8KrbtIrBtR94hmSrSTLKble9L69CZ7IlUui1p7ZTM+Czv/tiJSbfyiQ
dBgrD8kkRJU9hFgZm4BEskv4Cct1C93XN7I5XZFXSnqrLNcgPHzFUVgKol0W6Ycv
Obwo67+b3/j46H0OqxNBhbFknhZhm1oi1nwq7+J7HQfUxOnmqaj0pkTV+bqhr8OD
o3nGlpvc6UGnZLXr6XQjq6W6KxguF2apLOEBCj+0OrtPDTLUUgrfMCd0Lt9FXtJQ
Z2iMNvhqBrQqWbeuq7tY3KlhUY59NLmQ/GLJofqU3quOC4uJtnAt5qkBc5z72zn0
sk9peC8OIxtI3p8NdVfscR8cetGI4N/3MGQoHuUAmzQDJUs0r+VMuOhrjhAU4mCr
YcfxrB4tb8cybP0sm2yfg916zbClmszrJC40ssvX36xIE+RRc7+MNTYZ60R/Q79B
Fu6oCyt484753Fk2I/3vyaKa6Jk1fS6h5XViC+sSxOLDqu47sfPFspY9tPpEh90A
tKN91ZasAk1Zh+Pmm2slUM9xfX+Zyv3jdWW0yiwCbX72bhBOK4MwLh106h+R1Z5H
SttEErjaDGIDyV/41dyRF3kpgRQnCPzwDLe/G/B7oX7hTzvKHjUgU8EyWG1DOSJP
FlvtjhmjgbMgty/d6pSYAXFPOwj+MA98sVc0r55ztNJOu6jrMcUKKuFJBd827tqf
W6EHkdvttGWzkxlMXyFXw9EJO4IRXO1mJaPC/7PhmqR3xsZxGhe2BMO2U3bjVzZ3
Fo1Nz3BnrXd9/6x8gXtYH+ppNRYJI81t5Ew/K5XvOxc9kHBKLvANbgUm/F1Gz30s
jyhyclsTHIhP4jGNriGy28voDgu1bwtBSIahRXRlpZqtAxvw/ytszEWKqNZx55Vd
CFebVgx4Kl5rrMRdnTumUQfCyP0MKANQWCutnIJ+us2sKijN89Zptrr3y82D62Jd
eZv1ldhY9ZYqPY+theHhQLcFG1qk9o8qmiJrRLsxv7SGqDAkQh2IYBIApZdY0Dub
nE2ENS3g98VHBU9KoTKx4PLLnP66q64cP0r0O6uFf9Qlaac4siXKRyLy2L65z6wp
v0vxuYpug5RjsFcKts/LcItouJhbSY33K0LhBvBZ37INpyzpBn/E9o80dByoCpZE
0XMGBqVwpdmZKTaH33rmVoMnshDSiXl7mH3fXILNPUNH6w/RjHyIqHc8FPZpN+3K
P0P/L+VBFFy9ELlHjXnF4T6JQo6uCmN8h5Z9nzZ71yOLFmQxf3K8XTcajTx8GWwj
fz5+93BT2jd3+6itdmeQt7iJaBPjYZs9UxwVbp2XQVa9+qtzUZLKQb1R4aGtf+iS
qEbJeLCe8RY+Cj6POHW50bBRoY0wrMGhbBu71X4dDKBsQv5Tzhxwpad2Mg5ROWwj
vo9xYMF0TlaRoIdI5veLhe2Fl0inabG+EUK8TxAAkmSCbt2XGLr+ak1hddTHyyCI
+NDl2OuUMxbqwxoL78d3MfOq61TRYol6dzq/qux3KCZl26lC/J251cc+5PO3zytL
Jq1KVHK8Mpgan1T7IU0nkpMvXa2EuGBRCX9YopJjED5RxEWE3yexBOl5U7hap8xg
dGEZh6ZqoRT3ZIRL24piljp6vugadBaXguiiRoB8NNhiYZDsEmowyWaoCq2GkFmo
DksmlUQuf61pZ3rcsF2Gfnq2Hja8DdB5/9u4RQxpomT+/6D13ivt8i/5/cP2YKZf
cjomT7At96oGUlWR3T7Rzo2XwGlsCR2fNF5HGIFmiym9c9ObKMk3i8rV91DIP81X
RACfIcYRz+vT29GvP77lc5j+3jxqhWLHBdDO1bk4mSxqsmTloR08AuDn506bLca2
IklVEqh84qUKUlmjNnpS9LHbbqojB3mDKBlhFNnrl6nf+kD+xzGM1a45NR0oqkIf
yci8c/RCjV6tPnM6MQZ++1DghIuibpV6Gpy0ocSfvXi44JySl/YABgOZ0Q2wBQlv
i4kzxqRSTZfTRJ6W7WOEWLOrfS+Uzh3Rt99rWKiWvKSvXLQUSuOAI0rxJ4u+EdjG
NwcvpZHjX8LafqEiCTJsmRZ1R6C0gqDnu1NJB3g2yr8ktN/FXpUr47bRydSK9BpW
gTImWs8DZOt9+6KUssxjCpNM/9tZEVAhCSPPBlCtyTWvlyO91CFxk//IuqkoqwK0
r3jPhTh3tE+oc9Rz8nfzMAYbvvGZIuFInCxM7pRsFAaVc2ZzVyQyBdolFNlIH56Y
GWhd2CQka/fzqTQv5KwuTH6eiO1CP0dRpq6oTRfMYwk/jiN8IRskbUWoAu0Fld/r
xyTaDgKtZx0AR6KgmujCrB6ekR91bika8DUrgpNwKUk=
`protect END_PROTECTED
