`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83Va7Dt9+bVIX0t4hLH6KFTnoYJo9bQB7cm2tpfurKSIoRf3ipBkPSZLT2EzFZAE
aM2RnI/NB2qoH/VwOI04zrEQajyTub8E9GXps1evfjYH0mBn1/uEtV0dQ2zOZ5ZD
Q3L2gAskJ6/2lJWgQK2rxJFIY2HJjdrcF31RFHmsQrUMUgYvdTJyNb+Lb3iMTPIu
jw55QXgK5p2YsvsmiRTgcN9EVJ6x/1xHdQ2fD7POijqCTBZo5qFLWpVpwRbPC0Q6
kAZfGG3IiV56Z97uKLwhk0LK7lpS4RfZhg69WzX5QVxhuvKP7aAqljGg0ufh4rf2
wzRVZhpouhUGtIl1YLgjttaA9cP/bMOAnVtntBQwWXnzvtEQUp9PS5/amHkS9udA
13FmJdMHp1xn0a43ybqeklN1T+3BOYfMGK18RB2pL+2Y9f4QwXGkONMaTp9UFyyn
Cx27YvdQUBiG3P0mhCOr4dh6QRKDO3x3URInGNGPURZogRrbP2JAOZIR9LR+b8+S
BMzEAeSXCRGiURAYVnBtVTOFB2lNHuxW9NYHVZWZD9on3IXAGEneweizlCjMYc1U
v3HfC8x33OuFY+if5d6m/KKXYD4UOrGIQ4fo1Sz4Ck1utYxqvRmc/2hDP//5n4af
gn5ybyWizPeXbUxCu06oeg==
`protect END_PROTECTED
