`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0EI24mWfHNI7iWtUTK2S8C7K+snnkc+bKfL/MOSMoBn3eaD/iUY2TDrxM2626D63
bZT6Whb8vmq5Kj5iRqY7P/KcYE+zbNSZi11SbFziV3wf1bieN27WDQoXOrZMts5S
ZxsReXv4mZZUnxKoXgXS35DihyiGmvP9saXmHu1BNoDQ/5G9g8LhKS4SuzCGmZb4
kw7m3TzFi/S+VavNwuvpfGDeZAKaVehbb0X4JJ7Yrr6ZEhxwsIH01drliu0PQG4P
6V3dQF5WQTLXMa+IszQtZ7T7rehEDccWkbxhmeTsAbAHONIBvuqEipkDPaN0gBYp
aOht3+Sv4DLOYBXMKtaRcPZ8YoLb8HlgDVqL/xdDfcdI/ZpJptp+1Ay7NCu0rSvm
AXMtZjRpa/SRHo/2xzB4hMVOk5WD+2eNpoF5ioBU/oXzHSZvsAiypfoNjNK9Jh2W
eh5prLKDS43/gO/tLcraEZBXaGStjI+Eg45rX4Jb4DLTXAY9Sy30GT2PMeku41V4
ByVJDleq91OA+EAtPSKh7SDJn4yAmdECLjNaTLOD0S6F9Jc0UlrrfRW0/Ev+LOdQ
mFdXaywLsZejmL0+h9g624mUEsoD1cIGDdbeYT3xhwU3CD/Pggpv0FcUDfUQSB7n
MtQT0XboofCybaTriX886JmH1sDS3gy4KFaXZa8LQ4wK6v14+UUSSOJY6gbjxj82
BL+J4oXf8z1dwRrtlR8Crl6MeXRYQLwg/Mb7a0l9GAtGQvUJZJSZ044TY+o6zU3z
AQBIntCQY4SwS66hE53EjzfHEKlvpzCIq7ISngehXyItJJQLIFKGU5m7rG7T6FnG
GtCR65oFj2YbgdwDqBuLic4J3o+c0MkjYzf1Tyzck8Q=
`protect END_PROTECTED
