`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMqkFWIxZjFTcS4j6QK41dZ5A8TxvVtlKH1mCZsOlY1E/40vIeXUz6zI0j5XPWo2
nvdwscr18VgJe3Uk/NtLtUVHsR7CP5lV74D+oYBGvRVOYvVE7yR5E/RPFjJz2FgC
frJ1B/phnK5fkq02O4HyVVtyiED8j/GY73f6/rUPruGp0RcXjq5WcnLZhjbWX+Ym
q5vyqrfeu4+FrEeLYINli88YHMDy8HXge5QjZH+IUhMoWkeEYR5ytetJlt26htjm
40m3H2VpggXv6dZUYUeEA3eFNCDJu+NkinF2FdFkN7FUAajwABJNxH8/kwm9fGar
T5rXgEw4sykhOH+81d3hFQ==
`protect END_PROTECTED
