`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuny7Ht1QfPXHIV23scLwPQEB/dQiLVi4q7kH0q8gVIH+1Sexno49pj/IbWX1Vry
2LnczEcUY+OOXDNZqdS+VfX+IuM/Rv1rmGuTdG1Brhun+I5UXKJCbz2CmDEwIUpw
TJXXyghZKiIasP3C9tcJh0+QuMe26L7ot9CDR8Joi8IqdXJpWDvjIw8tZahGZnPG
nHQ5nzOVadvwF4BUonnr5xMTzCN11RJ02gaEss3vdgZ6o9ooEXZRHPSOnDG0QX/F
cK+BFNMhiebVXyPMutFltmD+SFzSqoISdNtT0tjUe/NItDWOmID47VBtcARu9mo0
0kJKscP9velj5f7ny2XCMM2ek1WkW6gsiwHTldqbWI4KXkImdpgdSnyoNXmqR34G
pFdqrBoCTUmRR/hzNfT9RcmufCnjagBu3oOahya9BV0yyjFc26UeNqSWNMdgnf37
PxnS/zILLFwRvlLEW61UZHKiDh6CaAUuQGO9Pd3vTPadOpx8ycxnqbosVE6gOiR4
yE1MX/DP11Q7en0sICBwcJv+xexMJI+rqI9hOyhMG/bCxu/Eu93ifMaVv1qTWbbU
+Sr1tXj5orvnOSfFRsjP9Cpu9rNeDTCU8qhfI1/lxMk1+XFKbsMebZEjksZri7cQ
tJ6NF5Q0tj6n7Wd0CpTYIg==
`protect END_PROTECTED
