`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
usPDfZ4zUT9F4o287shUwJrAlJtVcADKE23LD/xH+kUGs50Rc96ybm5I1Rc3VAnA
1rKmsQVOmm+mMDr3FS5HQR8kcYfF5YeTNethOSdOGbG+ROo/JF1ERY/3ERiqskcb
a6dj+CTzU3XzVthUAzXCfZn+HYj4VjqJYOuB+rZez5ddfl2aOONX4ikhOCHIMgtT
R4VCqGt17CsgmLJpMnyrSz6zIYmspEke1FbsryWt0irRwqZlCJd2tvElhW+oYQEJ
I0jYgYnQse0vzoD2/5IX/JXfRRBxYCIb8ZdnogYpm7OWFHdSbOOPsdRKejDZuDMt
xeRGm6E3Awsn31cYsjVOom2NjFOWZqEDYbOhpd9mGwVVXWb+UwFl1rDHY11QOSIm
Dov9r9RZr3enGIlGIj4FmOogkGXrg7e5O/ZjmgtierYbNqiq+5A7dkfoBHGOAvfd
90io3zVKkLITGjBAMmSQ3x5eHSIRj3BKFkdD3jpZo2EtqWusEx3IKlKrd7Dm77b6
NYi6Ut9csRN3uAmRZF7KkWDDzWyUatyQ5dP6gQhM9u4u/Q0Q8kVKqN9fTRG0jor1
zcR6NmdKEer9RyezlRwGDs5ep2KsXCrPy1XiqjUIuc/qZRNHJvrHBJRUeBb45NTg
fTw44b/dyNimTI3MiMFxAt3ebyw5uscZVDd1srVtE8iyaEfEV6d7Soc2GNkFee61
hkA50KslNDrOmkPKaiVv+e8YUOJ2YI9zwXKWdFzOAP0IdPyfStoJNaAQR/k5+i8g
0YDoevTZkHQCEzm4S1GuIY0AjfZgQFT6TXx5z1wPSYYjaObnmPdoYJDhO7lN4Paq
CaVKLjxueiCVDvyT+ei4zBBnDvvAg8QGyn8sonJ3StTjf8Dcnm1j4GmJqV0O34Or
Z2lJYsV6Ru1MtdmG/VbQN/vRup8VGv23DbcnGdCBxMI9223XJESxu0xISprFJMAu
3DBZEdzIHjaCN0MG8lfnHIX+aPTkjO/PQ6SPfKykxxhlghxOsA0bzMwa0gHdqk1q
jMzg5L+UGp4rgDRptJN7egRgJgRPyVooeR/BYTkTCUwGKVm6eWO63fr+LxIv2acL
LeOTXlhFAuV7HWYukVpqIeBziGswk4Qu09+Vj2VvL9unjy67Q5h8hxWrrNmFDayG
17AfI+e+6Qif7ilCyZ6rvTBuj5Agw8yeHEdrvpCf9wdBv0cQ/BpAlW5LORXjOfDS
3XPIB7ORzDzJAKcEVVCn5ho9kr4oBN9OktqJ+uR6XLTaL4iw9Ba2rED+gO4DryKr
CUsEhyh2NsYKEANJoAKR2l7eNvvaKkP3YC0kgkcFRzBOGQ10icWTPKRs6BjqKdko
Pmn9Hb79sfpV+xcZHpTwOFwM14k9+wiY1NfzrEgWJcTYKBQ5TEGpezoWbVqBIjv1
tx7HLS070XEOVMVGMm6OYwEr9psGOrQJw8pnqiYXBM2qk0/cN4jNXufZQCQEE0S5
PGd0NJEwWBpCaadRCEm08hhzEFlZbKyh1EPxBLOWp3vrLaphIGiIwPLjbJ5x8JNy
GIr/skEueBzYksy8tbYVOl0Uzw+yyhF0NBKkzbdmPzM=
`protect END_PROTECTED
