`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vEWiE/255bKXVf7YtZv6TxOrfWnyCJk5HwPUp89/bBfWmSs39Y2MnvL2mjQKZo7b
kGF7WdvM0OO3IIpmwYHU0M8uLF+BVenA/rUJgiZ9MBYbdLFvQrKlJ8+GKYykcEoJ
2Do90wg1JZ/yGB68BRueVsSz4c/OJqpDc2cQgBwGoecxfE7xmGGIyBgyMSjJUEqB
PpYHjjIykwdBgppz6nLfamaBdQGWjGMAK6rJzLGfW64LFgAMsXWj3npDop2uJaB9
ZnTlxs0IjtQHl+Kt4pEoTQ2pCGY8upzFlSafqQkjmPsDmCQxMpXQgpNU/hqjjpUG
GvBKoUnp7bb+ze48eE49stJ5YENSStkpbttgWMIAmKb75ku7h9FpzKZAokbC4M1s
UtAB+T7yIpfudMUQ7dbdYom6HVwbXFhIf3tsGPVdRkDwHrcmVeFDRV9wSnVu0Pi2
qfmfJ9HFouY4j1Vw8ummK6isXyl4dxSAVTT1wLwLR18=
`protect END_PROTECTED
