`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMoiq0G54CF2fdTErXFLaetOoKlisf6Wz4uykBjvjs8TiBu7qtynUR14QmM4LEGO
LtEar5A9+v9H43ZktYS/3f6mGORkxqmNPtQ+4ob4LGqC8V5jMxugbSjNjrvVrUaI
p7lhZwEfl2yHXlzJSnkCxnQrkP/oaeGLpqlKX85u2p7xjw/A6yoxr6TjU6BkCV2j
EHNKxAT9uoNCQ/Z/QIGFUhWn4ICzyO+xVqOwjQy1yqw4nw6Yrwc3e8dmZkH2ahJx
pxPoUii1epGPQm/K9rAlgoeqsxj9ttfnEG9ALoeSxOpKnlT2UmwjB9bcGEJreTLQ
LPas3wMmt9R/giOaWabQRBbfezd3AHz1MddOAFKkOvrP+j5Ai05Bu7MzwvVU+bPM
+fWiUs4a3UD7yi7uAZmlhoYWqkyQrj4J86HJUBeDneBX4nPtu0VoW/tzfnsSCGjo
ZQHr716zd8rPAkgRLAi44V7ltZ5n5bGb9F8Ac6f3XQALXZt7ZLi201y+yEJwwjW7
GWyaNFBjzySxXh0/ySJcaIGiZ4clBNtuqUvbRy22UbxGZZMSKEVbPUZSuwsWjGPo
vVLEpuhArHhcZ32aFUwyLCj9lRD3/leLJF82KvW1LYyoQA9cAcii7uXqA4+0oLHM
m5EFgpc6Erb28rDkO3PDLmSRNyCQa6N1Y07jUfjg5EbVLKNbzcRI92/dQ3UtJlvV
3ek28Rxm1gUQYGSkRv4TYekb9z+nlWvdJ2xRuGTFo6yxaKstsSSuyYo6KN73JNYu
qJxJ+DOoK8vZmvK/MaqxQqqEoCTJaG3bHrS1HacBXSPURj4ka//Ap0Hbk89vdG9j
YGytfbKpzBhy4Ro161rAG3VATMa3eYsDFEM0jzmNmdynSuWRRT8apC+fTpZv0+YM
/UfmS8WY2Z5onrGNsUsWh5YiVWbEbnJ4WG+sY4LKf6NBfOTOYMzHrheuDScOiCJC
8zgfaFzyy12DC+/WKyPUhMSkttTpXuUPGAWC8QGCQ1T0XuWryLm3M6LoXRhPejpR
Sp7hur1jjkUOoovzgfTCIgaZYNpjKnVR6ctiCI8oT4wk6EqcbwJEtQRNuWletzM6
GN7n89IieuaEogiHXfWxaKkk5TuUhEgngKwQbkgAoLclPemt0iP+Bzk3T6TLpODJ
QR0hx6w4Rgyj0wmNlIHfx8OAnhNiNCzkAhepNkW2qO6S/duuLH5l27AOTwANGC1Z
qmgXwnCa7/MmCqh8DtiQXZQk2m2BCLb+uiANmOVs8hl16y2+vkwL59yS+PW6KFEt
5gix7YX66nduCq3/babs23m53X9iALNhk5Ud2XVqxcMfYnhrwLKkqrvRdRltfBSr
RoB1v0MxpwysAo66gZKjZQ==
`protect END_PROTECTED
