`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6v29HDjfwF6hmIarCdfSTUluKgvpSO8Wa3fLtT4b2mEAiBfQBNGjuT0yiGvgJnda
xM4SMg1DVj+mescbPkaykQuFfJxyXD5AAZp1OxwzKVTrN8Kp5b1bTB3ewSrETE7M
tiQ/0IvBzu6fqlYBrPWzRPCbxpo8gnExa6CDGZT4eSrZJqIJHlcL1jlwZey9JbTx
zwgQeGb817FLqPuGsWZhfOeLogatW1Hp7VU6Zaoa+47P7WZI/XOzu9P8/g6opksv
rajZx6lwctVGMWAKgZ39FdPZSwHFXxtQuy7VtxONWThRw7Jn5i5bxlle3BFnEXEy
heaJg+skF7kwF2ok31WvRCBUcyQX8DZiaTybIZxwqVU78daXiY7Di+FTb1HVZaD1
Ql0kawBzhG+l4eJCwfVqgbAk3sS3F+gaBxGqaQ7j5vZE+ShR3FZjU66pTimOuF3Z
MRdcgP/XI4p4S8dTN8+RawPXP/VYwdQ4yFHKjrTO+WNkm1In0pxSf3lWHwY9iBOy
I6yL4EJfNvR0GEvC6faIThn9SOKytmHeQpnYvpmex038WhZTZwHR4kPW8neokg1c
`protect END_PROTECTED
