`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npeMjcI0y06CImgG00ESYQZ+iUvSDbDA/O763HZN0v2xdnLBaGAJZQvLHL8XMi6K
ulYIJMoizTmIkVEIfZFMUnqQbXWxRPYOZAM03F3NgyUgtWg6AgPWgJAxJ5XJ02hE
1O7ObzOu2CkvvuNwoRV/nPdoXb5WHN0KwLjv1vrEkprg8v1YFJZq1vpcdOjMo59x
iLk6K4cVdAW9TMGXm/Nk5yX5U8pIStKdkFg3KOacUEYIvqIsd2bZcYUXRLGJChGR
fd/Py1ZmPKsW56r6M1vv4618LydQoeniCoYIBmftIGOOZp0SdlwnQggXw/zKohXS
xMQaIp/yjrwxMdYBBIER3+yyu5Wo6URdbvxq7y2NXpOUKpRDqqyZ52xvOB0Tw1uq
8gXrn4iuzsZDhcIMJLOUW78oF06GWFCw3NCFtvbgYLMN+wI+L01XmxXJ+O9mwYEb
+Vue7+Jy0neuovQprZ4UCV0DvhKxunzRB1aNidgs/C4axOqe8oo7kpEhX1Agr71v
6C6FIRDqdMYiOfR8Vb5smShus8szV941QJpMDj8V+e5wXhpwL8jdHkZWTixZlQ9G
oY+1zv0++wSyck0ByOKXYoDOC7mqpLAaB6H1x9QWxt2w24kye7VubMxolu/iAron
zdMgIzAHoOOIm8HU7VlgFzWSOtTB2rhrXSqYBavGVa/27ObIRoPGFxmGFyYoW87y
fwnL/Tw5Tx+L7jKL7aFVfXe1kEwNvmZxVxflqor+ibrWflDi4fp2yVAvUKgFWMvl
NvtzeB4C1RiEHy2B/f5CtnGYxj/02Ht3gSqbLn5EBI6a/tAkubWgY4VAPVqxjt5U
gUyWElRVnVB6TdYEr3QBiTNM6r0W302JihxcUt8YFsml9oJMKvDLvd+VS6mGnqwi
dxXuhzArg7O80skPzdmj1kMfeRyJgjoClz82P6qQmG3yKdtRE47mYzGTCz8Y5Pb1
zPbD+TVpwkarq2ykoP92J4kfJ8ZSllBEDaGd+Obm2C3aAtXbZ6iPqYHqlK/r9M05
lWPoZUD635qPbQpn72BhUfSuTEg7i1D+3HjhYZh4/XQEa9lnVCIlzP6jCFQGYloA
aRa/eXbgfh4BBFD9HWHaNBfoh6puFa+jnrvf2PKVHTG/9PKmrbqK+Z3CbhKaPyCL
4RJ/CHg3by2uosRMHUd2Yr+UJO7n0DLP2MbR++iM8r0PsZ5v8RDiokIdBzqF7m1P
gEJf1Azq7rBl+ZrkxWwZmA==
`protect END_PROTECTED
