`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vYitAQ/SErbIFsHKrffkirNEmEWvZ9mF52Va2BiHp66877Hm4YfCkhIHmWorou3E
WqNFvJPKTL/KoqM0pK7vMkgvyZ6EJChalNksIx6dEtn+ZLRt0dsNoxkJs+2XJc8b
fmtaDjlT+r/GstfAYrD7X8uFFtusSubEPvWkKBDqTj09blL4tFhA5Wxx7gl2U9m/
V3DbAtEtp7Z5/MC2YGh3D5X98hRsIBvIyD/qOW61+eeohRIRQDZZddi/amMRIgsv
7QCPhvPHU3nZnn2CLKgMP+qgjS5Cn4ByXTE98+YqD4u5UMnyuKyXKVdzexm0jcFJ
xG27Yr1/tIzcouugx0rItYth5/O/8vHgZ7ZYmXHKHtuDBgEaA183rvRK9YlMqWNO
M0s2e6w/kfhl09ob9irlRg==
`protect END_PROTECTED
