`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v+51EBuGwKdiiClKouzy/rf3GCApHRJW3O3DQJjgCBUB29VZQbThpDQS+/XlNJeQ
MGju+AmF//GKMTBgSE2e19go6A1i1wHHm1zZLiGK0B6q+G6XerqfnM0qAl0PB5wO
Rfo+fPSbnz8Hp/bZKsTAPPXcSaqYHTJu8OEt9jx5aHZLhwtR50/+25E1bozAhAY8
RNEKPMmaCExOv7hiTYO2r4mYspS/3pEc6PpLinTzRpwiYGlyMvZ+lbtommmQ0ajX
d62SYytwlY+j5KqLgufyMw4cZ/iRy4rcGOSO5ith3HZQBm8GnOdi6yVbYbqa8hVt
W3/siaswNkl9yr+mDfX0MhX3IU0ObOAUlic+r/1T+6xr+6JgWMKyy+H3lR2ZEnN+
P7J4gRh0Jra686OqRvLe7mMflUrHViochcsulplbeRe9sfSpRvBEHm7wVgeL9RXB
goJVMtwlBJAtZgiXrBcyaWuIefhPIlultfOxisoQkLM=
`protect END_PROTECTED
