`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fJ5ld7YdL350XMNVX421KKp1M1lyQ2ctJS1TtWmVIoQw3wJf/S4PqELE63DqS2Q/
/zknlH01MxcqYZEU3IqRyrOD+dGzEnIrPS9GUokWIQCmsHyPxR16Sb8soXl8MsND
m5KMPcqBnb76k4N6dh7XKINEaoF2ExZbMKvGKaUH+OPxL0QHGgCYFPtC/Lg1XSRs
a/rCeI3wTTYKsVewRe749Q/8fU8CpEs7ZWoNRTbcCg8DbF7veK/KDuAbxhI15jnI
rBUMZMcnHPVfn8yzRaYf9cN5n7PRyxZlUCarBXLqqt/F6mUCIM0HIhwTmDb8uVOa
vXWOzXgR+e+vf9cvzgtSJdezY52+kjhE1VIvznlLjsKKI/2q8vwfJg+DMQrZY6+D
DQtSkca11Aj3TKxmoCeWWdQmeMzRBh0gdmbD65+OuWKzNsSbRkWFBjAdQZWJ3cv7
0FZzvZXOF4TGb/ANXaS0mnTfFicoLyBJTvQ+51LUN7eea87sGVBC6WSI6MSPo4e0
sAURg7zbZtg+2zZ4jRfMwKioHr/eYiXKcRkyweeV22te9v1k3sdaKdrJ3ALkDyZU
IWULvFnC+7qM5ZTOG7Ebekmcg+tjR9LtK9f3mFdiGP3hdwzBs0tSUhZMXMRedVCj
t/2AG2pEoZzZP7tLUDUdp5H981js354RzLaJqfk0RDUDeL5bkfEWJg5+AflwqusU
/zfTgP0uJ6FDlgeVk78gB8PdFLPMNryBqNXBm6CKgyiIX2Jbo9hvqPtrZdGeLsHS
2dCczASoIWCePvY/5sUfrdAs0FDLih2AdhGEHAiuvZd/91j6830KaqczL3sEFevG
kBVUHCKxcm8EWlzkrLafSZ7V4NZrDjriHnckXjbXG6qej0N1A84G1QOxWh8POjqF
PSqIFSskebK5b1iqJ6ltHdztPpxDrTKzTt5aAkkkPvmUv/dFPWMqFAckLHXPz7tU
OamJ7sPqp3ScuJSiP1G9gfCIYO6RbjYqV9pIoqX0+JHniNH56KTJd0Ih4mBtAz0+
OAFPVZTDAOIltU67qe/N5sRJ6zoY0Djz34jMToaVnSS4mLVHzs+PeUp66kVp4H07
mQBi5pPHsirbwWISfNlQHFN756X28utjkEqSFQa90TWZgs7mQnjFfLa1RIdkeM3j
RC7uScOeuD1ElsNI4vFp5TV9i+v2EAyvJwxUnvIuU2pYpA9bNvxyxUZQGhZkl1aP
C6GMEBrXc0mO1wxt7M10wc7qtfp4BY2GvVeFpo6LQzA3Qpd4+iPotR9ahBuxsRf7
7C9bAI0Kza55YQ404vfTVqh1IbdthVElgsItIVL2YBxzAFxpuPpdGZMxktYuLCxv
a/XqeKAOjynSTeifcx+s91UWkkaNoW57kuhn3/AgfIkq7d98jIbQfPYg1I4rSbPq
cJ7Cc98cDLmaLQGEEjh0/0btDKBr9mJqhmOlPwJ3n6hIbYyIuPTw+i4h3GIIf7/4
l6SwjJG3K5Xhzei7I3erBsNaa4Zrqv8jCsPLAuCLynYl2qtOKPmnrqKyJTffk2m2
awEISwmodhHwvloziKytC+EGWKHTFNypGNCjaL7yBVZFLeZRB3ezaHV9eA+0hDVJ
4EjtfMKsbgo2Uvwt6A7wiVHD9IX/Q6fUrJjZnVS5FyjHQObwzWJl91qgQHBx/tVC
8wRyj2yownDr4Zs6DERWsvkXeB8hiuaFarR7/5XVeDjIfInDjyZcKMNwY4PDg7TL
983ACM3EUiNFIPxuYtyotulOVMwfrBS+C3bHUEi41Ic6x27UInvFGNHKGld/jOdq
+WkNdkhGsRSY/olKEMVeqvH1/hMMXC40RhTf4YCnYdKP63QkyuCbMheHantRJFn2
wzwvDui4YQyvlQMHxj+4CxW8hmk9XZwTYkhucO7iRSemKn3nWU64q64/dCWLv0Ji
5F51MbP2fL/8y/eEkU3vuRKgx1iJ6rRCJEY0eWdAgwHd5Ibimx8uvrzxBcTMInsN
dCSNpWe+Wjhxhk0huMcTA+pn/PUHw3nkAQYFUhGh4XwbFfBu8Jb4gn0Vjy6nW3Kh
ld1tixArv1bMkkKeW/PQHGpAWP91Qy7D1RBmsb0gFLLoF+AF2RCWNSsOTV2JtL4K
7/KapOi1q48lr0TOu7rP22v3AjPQYFeYnUF7ozUQfVCtBzOFykdlwA+pgciYiSh4
dcZ1M8OVqfyMgpvPboRbVORdELUxWrLWGT2I7v+pQ0tGje+uGU0DudBZf5a+KiRM
uQ8CMUzSUISCQ6OquSf9SXYrApgJgMz/pJpSUJ/l+04Gy5bcw5N/HMpaFP4nCEDd
8VpeuhwDA1el5pYRcbw9m0fpOzIt0PJwP2izEBDd0HeJiPq6IkNiDjATa6pTVK4w
Fqdj9eFEd5dZrpLzBoYmYRcZa5LureFzy2KSfngOD242t9rDr1gu6mG8M4WBT7Vz
mnDaabdn0i6ztZNzCxi7KyCa5oji5LicnS1Tn9Y7BwLQCqkTtOJBSgWMQEbHdwnq
4I1oBvszqFsW+YijfGVY2hDdyjDlUPaYxchORQYX+LjiKSOdXkg7A4r/PuoBvndL
Z2oJ+haNGZcUvrcCnPQGfN+aqGqazKY4P3tkOsixLBsFSKibefquPcxc3hOfrdDP
me61CrktAApSkvSe8DwoIp7Y/aFM2ymVRmJfJvV0reAt5Ac83iyGH8EJwOfkCUwg
Ht5aV+Mw9IJEBX9dQyN5om3c6Smzq3f2Ot5qoz09kiqjrZ8zSldjjXmLaHrzBdsx
dVCiO37hjzUv2J983a0NYAC6XLffEtAHJOXtPZfLWOacpeyX1Bifr9jn5vnfL81L
4H8es+O1+Uzi3j4Ie7WPury1GqXdrMhZ1H/QLauUlKto43L0zVt77yEB9f3J+9z/
KLa3LN1kAElc4tF+upaTvTNgwWa4pk5HoTk3YoQK+Oq09eJKGuEhyzw1kIGMMFWI
BQLbW3cR54ES1tw1zDiCTI8JJpaWSRH7zFNqeDf5D/PBSmkekZ9Hw1wQ/nLzTdj7
2gtMkp8l9SIxfOZkbi+3bHcWJzri2dUoHMiTWkpeBCFFuyXY1Zjlln7o/zEE0B3D
/zj/pnPNhSRFPpGHJ+qRR7l5ZfhSh9WsDUiMndH9S+AQLpZUkoG/H6C1KSAF+ZOM
3LsPz6H1oS/Zr9ymoHAxa2v5FhNalNzAvyHPLYxaEGTP6Q3D2/tcHrm5JfgCoFO5
FP2RIvh2XtiBoOA6SiwQ4bwvC9w7+kwvm4Vm3Q1tPNE8X3IVNswplyIda6a2MH7L
FHGQSEHi8ImoUFMu7ocuXs4mvAqZvlMGs7xB1OXhZ+1jZnHpUiG9yWmffhDDMukp
FL4HnPCHXm+mSvw6NGbWat2vm0LvS4lUQ6Py38Jsryye8QadsYyBXaBT+mdRTD5A
aU5zZ8yfmSvcyHhWYpQaItieWYBwmBHMWs2wMDJIEkZqbs36Yy5LWHasBMCw5EMA
1X1i5PwFk75+RRMe+GWt8o5mQijCOzpMtHuvTLLpcy/KPVLF/EQu4akmp7mnsDF4
fhleNrieKveyjWS2+F+yBj3mBRKd7sA5yNN71W3iu4lEmHAX8vQSWzUleGPbABzm
xp03hP04W8gmOAm6vNHJWdjFWiAnJjIKxzWAz4r0MqowD7jopI1121p79pmIMCMe
bXe6bvMRFoVDHF5dSR+rXcTratisp+CgVJ4t4m9q8iq/qypxB0+nZ1c2dxpZcmqc
2tvjntWDWQFZotfSReXwqm9D+YZ2SnL9sy2sWFf6zskSqeHUmcl08mzDGZ3p13nX
pc37oQ7X7W/AIyV5V45TLiobf1A1efrTTSUHD/B9F96MRehBeofxY5GaKhUMJYMz
a2YP9dqRns3+1mjQD1etJSNqYtfDDrS4rhXE+9vie8RPFm/AXmTrHBQhq14XCHbM
nFS52pd7AQS2vo2WAuMLOehq1usjfCJx3eYKGxskDIar3dLp5YY3/8KxNZqJf6rE
eQ8jyeD4llW6fo4IDtCn8qNkpn8Yf8UR3i4+RYz25XfmX6FcetHQNQaQsjuSOiAe
EnBf1lWZtBslrDByztbyeQILsg9ImNb66r0+uCHCMV/kzplkdCBmSD9PifcffHGj
B8sAKpO021sYdm2b0VgZyZiSV+xIzpG/PFtaQjmiRCuajfol/nERlkS5TB4CEPba
Iux+zDMwpdqdUPRUXfQfmrs2Hf5vpaM9YyS585v/1PX/JobHT5QpLQAay2uAI1A4
pzHlQwT12/wKpR+l665ExZrS6jZtXfzXjwtPwC1yY/GuLysq5ykMEoT2EaBoFfv/
R4+0c+rZrCtLP0WmITpONQuIOvn3teoCwGvmMkprvcZKGq0Rwd8DplEZ7yPRh6Rx
oHEmolDgvvIcHIvcicFYceqbiBPgNrM732jH1Q5ayb65u3toAUrq0Ws1R+U42EjQ
s4N5sk1KRBd6bPc9uUgcafFc9MdzCn3E7cwtXwiRyQKX9rpmLRanG/Xz9wsOzetD
1blqk2JyjlHgwMnTlKfgfpohKCYxztA6HzkO6SZ1tCc1WPeHVq9DlVaPzfdZHD5u
KP09hr/fsWhD1onAoRX4vHhbQILu8PZB6/4lv26RMzhbCpLbj+ERhRWqKlREsdr7
yFjoeoYRhXzUzNcNJXGZfrGZw9AvizSDi8PArqybnLelBsUeHNFyZ7iiElVXhlrx
LM83cd2/BL6YdXhNah4Zj112WqxKvwuMIGPxAMlWPEPsJPsBmoIKSEd0EYmw7v5G
4qH9bM8CShKkxPuyS+9I3zKoEwZYFvujkQWxT8yGFEzkyFhqsUXWHWEiBzXD33SL
1lpjlUR9H9lhac8SndQ8bbm7ak7gM0/LHpaY/8l4w4G7fNXhdS1W/dSeRBT4jTep
jclVzZ4GvgFLgqJQb634zsGLztDDAh7lrOx6bK0cM44oOSZVoI0mSGRzKuNt7S3B
JZ4g/m6ixyJoW6XkHZSitQ84g9gjJGhgZ4qOv+4jG7iykN+vypytuzdLRW562GbD
WBWAuunEV301/7kB/pUKv3zgPPbQB/aROVOpxgCnbv0BiB9zAVocap3T55olJbf/
H6ZDM1HkQM8kcnj4s2tG86sho0BPC/DPC8emCyUXkrMliwGF8IBriwMBNu9y/doS
Kml8Q/hWue8D822Gs6qPdluNvHQ29NOdWuXbJf0CALX4KHI03SgqZhlbUO1uEtKA
zvK7QEm/qdXWzpGFzyLUhIEFDLCZvqYEmET+uS2ZBFBnZyW62EAmElY3PPm3Nhcx
SwjRP/2XNNxuk7UHmJVzwB81DtV5RnaJVu9qdCmmeg9lyW72fSG3KemMEzNIGnRZ
LXovmZW1dsbndbbf4XVDaors6u7NoZTv9OsuVknjGC7z6r02Y0dS7ctzTkq5yF5E
pPjJH34Exc3Vlh4xLOUzthAJpgtGYSdzSM+bJYEt3SJd+Km+79rEU3JkNxxQVOrZ
KuYqfvRMEQkXQAEIrhlzsE9UG7o1JGNGOe1+0bEzug0XXI9tIpF3YHqIMrAxb5CJ
gbQYPJqB8h3ZyOFxfP3cwywZw0y6Ixea1MNyqKOqwbu27oQX4Z967YMIPUN4j6yP
EQIVFX0hgqT4ZcexEszaa8UUAWIBd/TT73sX3B5sCW2nJyV4/7H9f6RJsjrnrHrn
HarXrr/E5BecNJz3P7QOaAgdgQKMi7M+cU+UxvWVeG798znCVDxny7WvzFhBFtI7
Eq31TuE03c6hkkv9I98O70CT/CMM4jcEpRgW8kVoWQculnLODTLvJ0UJ/hR9oOi2
jhixYWsZ91mbjB75P3XZH1XkynoSo5UMuu6g2YH+6f1As9AaR1wESI6HfcwG9hlw
i+gObt1W+O0GBWmSqUsN1QjpO2EOyBH734uoZHRsTXpMsXyadytOMJVxTmeAmEan
xwUR89kmbVzb4Rx6JTFSvTkXlFtouHrPzYQWEzxuuZnxcIzghWQOGa+jc/5QE4HK
TKBKewF97hXm+IFFBZ5x51NIFAW5rDu0R/zAISGiCnc/rdvmVOQmQt2uc0LX/aUv
bJOLm3MnyTm8ZVrWEiKmjj1NqErq7ilZc5BQ9KhXMnHlHhrf9JJoGcMOzC2IgOnc
gtIU+lZstJMdyQyO5Tr5Wu8y3i0AxC39NfHSbiuCEDPiCZrco2nRc4vhglFiRZmF
PD+Q0aaDnv+clFAFEdkwdZ3br4ggLSfxvMoBAB5FDEQArBKx68aLU2ADgkrsuL6H
KmgUw4UPDYHJV4k0J+lEGssQqWIIZW880bH8Q4YM2MiSpBVSPlSdyHXVaOflUufe
WVG/+A/rjnP0IRMOAkaHI82otQX5FhAw1aK9nhKZl7pfEegBjVLi4oGB3FXNnuol
1Hu3BJkLCB7qaYR1a/5abChGeqW0Gl076gzDDUtEeUWSXt95znium5CBb9CtKnqZ
dnuKkwsJYyGlPuAzPRNK/zRWl78IjgM2Gzqkf0JgN06oCwUkxMQxSK/gNVEBLBe4
/2jnHC4Wt53TwugIJKt8DMjaCUjq2HbUkVKXz2bw76WG++VPF+5mkx9xgJMKKN4R
1d6TKzm6NOjn6VM3adwn/7eHykU3EoZpNKXe+nbOTEfXoQ2fOW10rrQcprHbKUdQ
i+iIIiwpVo9NwnIWJusETIiEBKVVfv2379788eK+QHE3EMDhbjv3OmzbHAmV7tPC
qB5NNFglpdghCwPMBqzfqCfmQSnTmqQZMKTucSfcxnTlAbOI721e+3zFwmjB4oDK
hjnvKAEqeRysY5PyKywNcAiqeeu/m+y5dRNBVdQQ+0PfcPAiSzU6OZONWplFW69M
7YuLd95IiUW3OVoedkBIM5+LYa1iKNj1Q1itwBr4P9yqqAmDNbDQsalZunm/fyXD
cPYXm2n2Pav/tiLhPEEa7OYCjrefQMLZefGNtTjOYKXOmTyOrSO4HIoVJwzCxdYF
ImJWMwR/hztvX216RflM4eZht9q556/tRahp2vqlWUNqf0q4PrmVh8yoLqLLAekd
LVGf6IokoLFAeDxec3/4XFnFcwpeumdjPtemaxokKmLwxOdgXEYIRMJbbQUC7a7o
pr89z5+a6VJAjFFZFsVPmGVsqbuv2xORUrUaoMnYcC1ntW3lXCxEUNowi1nCiB5n
qdu+FFeRB5zZyGLlMPT0rIaQrwuHPdfwo+2mkA8BVxY0RTFobGk1FlGjT6oQI7Hq
GxFsqi3ybksjTggEn6WqdS5S4uuL5jg6tWnwYl3hHwNed8CqjZWyBoUVNqF8HhG7
z85gAdxQCx/V1a+NId2eTI5VRApqtYrxJHbKxpaydYEFuVEIqFrXdq7QbTw6l8XQ
xUt/3NP+6iQjYg7OW/3nl61uj4QkXhy+BDpDgzdgYrbG+C5BlDRBTeIBQy76jZVJ
6RXc7DBGifCn28SeCR8gDxogDp5ypzV6KNgwSLf2smC5EHdYt/Wmyru56mquNaxh
ciPAIa6hwt8P67s7HfxJjEh0sMiryqbyNUca1HDiQ2+8Tv1Oxxmphw8ZG5bymov/
YvPMYYEdBoSR2PwRX1WwLPWMqwXATIq/bRhf3ohfgtErcD70CiCcENv/leeEBDbp
dln/1jaedO06u5UoqeVI0R+tNpdFXnXxuzDIPqWAOGnMPDakhEx9PTqnVvn9rE+O
ElHAu7kVj0aUb+DrFTr6q3x47QTcXKOQVBWOrQEFfPT1C+CldLIv0RyXZNcwjrpn
i/67aCF7CU4ZBLuSthQw7NPYfNbwXBQUlFY3GDeAkPithsEhwdi3l5srziUubPie
qr8Eyy2Fja6CXuf5NTxiRUGTTXzrZQse99HRfiNQ1KKPB4qo+3xy0SG1w5Ny4bhu
M10ckkSVuRUJ7dNGxDEpCckoz8jr9Ful8L40buoBeKH+iRhA+Q8dqIMjZE0TVuhG
ff6XBFkgk/9RezN/+J61eiFDHYRGC+2i3wAJrGjsKVHUNwEHTfnAyu484kOiIBF7
3crPL5BDaITptsdGiFkpdJmk2cTiUsLxTKq613RCUhfJ3BwM35Ur8e1FADfYu88a
cupmmklEwLGqgePKWwBH6hLRsm9iJRTbE9HWgjH0APN8et9ATIcStOqPlFogmG9D
BLt2uS7QXnuX196qAdxR9JEYnqH3d6fKzY6NMGs6jhzGWXbbGH+DANkV5BUDq7/e
KgUqLZWwkn3GP81V113ENiUxeFY9xNVebadQQAt+NZoi+H31A8e0QqBuXXAZ0i3v
L5ieEHJa/tBh13hcnlWW11+zhGSVFfLUjRBDKglSNKWgDY0njtZp2LdnlQUqqms2
p8LCC3nmu4/tVntet52YGCz+2nGqjw8hfemDJkWAcOGwIuMRbWnNSZR7ti2JHjNh
lT6ZpiW4LGzUHmCIrsIeiWUx4cWbXgDjyRhN/iH+dPoInm56enQirSLtM4wLTb7v
kyCP3kRcUnmnURQYxq0YIgZni9t7cszigs6TqlwH/k5xH05T7f3xOhE2p5Jut4V+
2XPq86Zgh8qI6i00o7HHEMEjmCNFqZy9V8LaQo87BLkyB7Qmk+2hSSQZJDff34S9
V3EABeiz2tF3vNmj2k1mJ+PaM5mAeB6iDm41tf6rqtGxzwWwSDlJdHSsXiw5iGUe
GPBmhfRi6Y8/8uo4KYfoBSClvsNoiIw/CE+NwpMIkaiVnMimiaaPz95FmrQt5reK
GqNAQ3CtXW7KmkkO47c1bJrEr6tbcnB08Aw9mzAFupArYneaLshyb3Y719w27nP0
k6k1FziIqMN8yZ2IBMBwuoUYrkxEUZIEyJRLBHMRaYktQ6X6batDw9HN7MNPBboH
cZFrsVlPSy7dnIfAgCLrRaM8Seo62AjCTLe8MVSmJij/j0ps3ASKCctu1gPGbb6u
o5M62ac6j9bFPaEoboGMZ2cZ8Icn6ZxdAdv1Z6zrkXqcE1HM30qg04CQk0QN+71S
SftXwfWnCWbXl1NkwVOfsX9Vr35OpNQu5buw0dGkPF5NVzS4jPqF/H5jqnNNZD3P
ludc8HVqnfpE4tEUDUWGwat8zarir0y0CyXoqlooDf3h6uf7rHzVQohsvUN4o3Ti
nGmiYkF+lv08DnRH+mt9JhwbMwHelDgBNrhVnE+hMT0cw8Lbi/AcWzDcgnuhca7n
llHRQvOrBN9/lWw7r2Cxcy8MotRnQNlpm5jOoqNSTstPcgcBsFu2cuetkMdoHGxd
KNnB6ly44xNftsE0I3no35qPvtLoxiHJ1+yKPd8eN0iflo+r24aDrLXNcpjDwY3k
5tbIlnDiCdE43cfOEA10K70NGQaq5TTQyfBsxKwyeRHyK+9XLdB3O6V6w4nkKkiD
2ZTiozqVE5TxjhmIFAv+8t/4VpuCzzVAM2w3YibqRlEV+O3S5EgOWDE6bSbGlFCL
aUteR0qquZXVrVFAhbV00t/x1l8WpNO3s2C0DLt9A1zOVMwPGwmVdhPrC61J2kZD
m5BeDEMci5yl7vAupomlWp6wYb9ZPW86nwhQZuSeMzR5im727XFRHrvaQg74zUU8
2gwhKGvLrI2w1AFZBq83+GUO7PQjOpQ8lC12Z8s8nccOE2t0CHJBHKNxV95ZsnND
VOyZxYWhvlD/AtXBCtOt7zDUkubUw3VT9I+jbu765EyyTR1y6FyKi4HemrN2yDMx
+VQy2Q7FMSgH5nsq0FPpnxG70xiEA9jIoPuYVN6Uhv5GekVj5VphxrAuwHKx7cYN
6CPsDjU4MgWSD5bsxLe01QVj1hTHVbrlVf/gxZ5O7g1WQ2lfzlDeoN9561+DOe1c
ZO7sYnBXt84i+wWmJqqxLuDBJ7rnM/GCpECCjNzYA024hwAPfEv331rxz6OJ+7WQ
Ipe/0IHNSgLrFmWNyYOGiSFasDHLK95pLypPrLP7h9Z4nPD9Ml0HRjcq62NTimQc
aPotTlNfMOwL2wk8e+MrcmEz+C6zKs9l09AHgP5JLTlUFVYbDgcj8NtOrr4t2MI5
KK8RWRmd16NmslCh26xutubwG4VIjmd4zuCHye27vZKDkSVYn4cmhwRfwJfTMJVf
gGL6NibBuH6n9Xq701mVX39aWUbSmvzVfkfBo3wLLsKvDdl41kgr2131oWax2yMC
E7uLGeQiBCkyzBkvdG74iENaGRbji0LueUXsVnlQJ5+E87giqd+DLTeJ7wOBX+Vd
xyKVDlRLtV2QKrRiwHR3W0vUL+JWKAyJrBTQsu4LiZhWPFbmFpO/n4y9eQERJfHm
5NIMjwf18FKAtwL43yd0TG713OsQIqBlN5bzgPq0TWcy2ECPLCIMOcUsRs4/ywWV
N+kBiyNoXqX2km1vOWnNUNAHetdQUvicFJ/D7t0/1sEmNI8e6oBQQEKg/QLqG+DO
Ao0FmZf2CzhePgtTCB1CuZhYjzb7Tm4w5L2vLritWgEXk1wqNBNbKoJ4rkRmD9kn
KJPu8QbqjPiX3B1Pny9N4qhb+46u5xg7vTypWGc82x9BB0eFjIMQmMye2h0DjKjm
pKnck1Ia+7vA4qDFmaSz1983vcK9pfmh+iCwHqfHCHTaRSTNFDs5n0psag4Fqfw6
tAcqVvsJQph7fSbf5H05Pll+qFyp/Hj+H/Gva5T3n2qTkGawAgLcyR/uRqTt9Ctx
z2X/ZEGM5Gj+EA4/cuKX0JfWz4H1Q7N+TUtYQiU1AZqU0kjxM89Oqdj0M6WWh4DT
qvYMoWbuw8V0Z9//JFeisYQRgQn/xRmHo4UkxIPcMfYo7moK6il7c/jmrkh/7PJf
j4HXCzETlwuZeFg+C36Ha6VjhpRRGlmg09ASACNoKKfEtfOOt/e51rTZ2PrUlC69
LrBj5uA8L3kwJn2htGeb4vf+4OjqxbjXKJ5vXTaMA2tMJrCugGkhoPcUlZx6xe3Z
7gCh5ii5XOY8MPgguEGGKSYKEpKwHk8SIJl8RGJ/Q7aR8wxl87eB59dTJH4P+eQU
PBgvvoK88RkKCyBKM4w78+C2OIBk9vvKJ17eiLlTE4VweUfKFz0yiB5xDQR58+vq
gO8C7UA2zlxDAemVlgPgyVohSKSpYhQum2jgP4f87w7QQDewnncrqnV7fD/9UdlV
sWVstvt7MAM44v6jcT3YtJlwAIAwwgGEABAws6QRtUc3FCQK9tsJ7n/0v4TqQIZq
ybecRkFyExq4wJ4WPrvURjs5FUyWkbtcnAEebteqNyGUn3U8aW61lECugdd/h2O3
/tPJ7Ars3j+j0EyCTIe37dPSQZ28ucdsEwMs6EXrma7mhjRZda5hRoDixApHPVh7
cLSJz55N6ZeddIft/36vvVvhvYZBktg2LSEllLC7RLVjr8OqVPl8O7qVeV4bgJu5
A5LVP+CHRiFTY9zKBaSY1ruMDncMt7p7BHJhwNqsp1J98bks3Ud5rTTzlPusKIgI
PcrWkh6EMZLhIdqmj2n6L0EgSpLBNQjbCTRurN+JZgyK6JpguDJFzWB1Y9/aaH8a
ZaAbfUs4bG0OcL7wikiX8FMnUW0Gh6lpCjYNe7ptslMSERnF+qMxV4uwnBqqNACe
cZAgJUVbg1iJo4XCN2Zwtr5Q7erH4f4tm2HmKvXxXHgTx4CWz2nyTFAxmHjJsCeS
JPHSe3mfj461PkSKUJu620SB6+p8cTIXBs0VVj8+F8usZirB3oMgaAsr+iyXNx1v
0AHIqcc77CzWnINwvjPUNrF64RRJMvJK4ZRx6bk/nXsyNL5b4KbmqtQEb7a2zxmx
W0LyQ4nr4+1OXZyt8dvMJBWbF0EV74rU0o7+JIPPEM2gfSdYTWr5Zva954wMpW5K
oY2k6IdTrwDFADs9/hproZI77tAZmbLB1GYePEkDUUrKKrAdExJ8D7cWiHVnWXo7
NTsPk7yi7XAFEggDKV84/SI1cyeCi8Ev5KR6dNW0Nin/uZuzRPkEAZLJoEiQaMGa
HCe9KGBJHshifA6pfLLMFR0ME3GO7dH5IiYA60OYXfnT3lcZUW8p5XZ4bBwarJ1G
geR4miDZvzbFjAP3Lv2MAD2RTeAVBxleYk+cGTvB5xT7yi88OEN7fZiDnBS9YlHb
a7kGdJbFyEU2ha92gPJU5SGe6Nmk0eg6Ul1KHOg4E28+jUS23+oQLC19yKjMJBbr
LnNkWk6D7FI8AbKkhk4x9nVnUbRASTq81Sf20LZxfw3U1tT98V6UeVVjto45UoN8
7EOL/OMyaItAABR1Y6xImT/GnH1U6PwSa6bqNpX8DJtpx42oLhMdsP2OdpLRZEMn
JdL13K0qfEQnhhyO810m9n0gJton7tkRznRj4jU5REKh+kUT37hi2xA6YoxbOpw8
urTovP07p0vhosaEgUU5JdOGIsELWgRV0bzEzuahtuGyxrsH9T7oFH13ChsAeTYQ
CVOgYOzkpwDOpYYyIWheNXdKT6rJOlEAcHR1ysX0f13GJwAFDWveZs3jYT+N+GMk
06yGc6AkqmZptnejJRw2BQPPz9FhBA2jdLqgQMvDX+wFdYoX2cWCKJh3MU5ajtjp
q8ftqbimwPyb+Cb+enLTPjr2Lca4NvahfT7ubMxGI5SzkkMQ3ocFlFxR194GMJRT
92dKLSmRD8wlzpcFUjqfVCvFP8i4qK74g/LL3RwL8dG5IyHjwoELsOz+I9K3RCpl
sKvvEZkCec4tOepYq4E2aijtFWCI1t0RP2FH1r+abBgp2179C6AupSCIECNwIlcM
8mrll3Wzh1RB6Om3MhcBIc15hpA6/RXEpTAKqNyq0ENMoYvg4ssDs346OKGZey8f
WpSDZ38lC3OACwFPTsKaeO01YJUNw+ZHVoWKyerMX1fUPJkseZuBtJXdd6bktrBb
w6SzYh7RnNRKAicQE0MYRvY73CoER0Pq+HOeaDDeTmNUFrU4l2g8tXsH0HBUl+GL
TYQeFUmF/Zar1WR51HxDfn6ba4D9tEGYZeM6T4UcFHTkfGOAtMewlG3oEE3cOPg0
8ORuoBJwTrN07XGKR1cutkfw8aiAIEd4HctMyOafcgtqJ6UQOsN1QVCrMMk5GVv0
ym9JpUmo8Gp4SsCXPwO/NoaOSwxVMREvuFL4qKEln4EAL61702blPWuo1k2ashtt
PHIYFJVVKgN0/mrIo/U0bZaqMjpngH4781vhox9mkCUHci7VNsxtXgm6HoYRJ7jb
Vb+Db/J59gojFgvVFgfhZw3g2oU5TPXHiYCgPrC4WvkqEx72zmyDhOjG7ymw2OcZ
jxyQdryGGZ3q8WVdcHocFdBCxjebhRDXszQ4pJhbfHPtTcLnfX6deIs9l2YYK5Iu
rtD18q67GBpGxxwI8om8RkaH8M2aJ1hNZ5hjzuydObgCOJJckqzsota7vkr0Z+Vi
aOm21TQPuUY5awlExSZvF+xIxs6q74wJAW4AiIWSfOn1Y8OzwcPqA1+wQBGke36y
O26aDwFTwU7JMd7wZJx7sFd7K5ypr9JT6lHzqBxxE7IjwyLCx69VlsPZ0Ii8YTjy
XLHP4JbrzlWuxuT4TG34wvoKUXf9rAkMcodGpN8WZXvI3q8HgW0rzIF8T5Xcnk7B
rJwvQe65pJQQWEJ8++mW0wwK4kJbEZtvlQ1sxOdnK4oFKaOB/qLLvKv4DOvw8+Hb
g0Fk3d5ONA7DINTVBTZMbBwR/rvPr9HXabIeJrxAnx03zMaRbEhOOEmkuLIua+Cp
uQXWZAACcVkjk2hbsMRYquyG8Ndzc1MNgCyJlMBAVnDLsjg7t2fYW2eB4hmL4gkN
/xun4k33REJaR+GlbbB6owDm2Rm0l9jXT4ACA2C2ulW+tg4hjaAIYBt2+4Dc3gQh
V9ovGGea38DhDv+IcBDIpC2TJpFnWX956xzzBTU2pMdMZ/zOgDv85turTp+BTIw0
TVhw9oibLUHByR11xlOsXGMowX0vXuaOLg39FjLneszp0UHoJ1siOlfV0XcWZHb/
g5qgWJDdReQpuYHoZ1GDT8s+PEqAHg/ZpV+jQEHb0PmA52j6qZy4hYeNpIVH1Kjl
s9Y/qEkKWjB5dFY6l54SOp9jnCPpBF7PTLq3L2LOhf62Kf2MzgwZDKL/wERp/MK7
EaGZ+Z46scvtJGMMTq45DbuCzYFDIS0LMwACcM0f8gHZhZO/cXUS2atkUF3pwxQL
b3PgNgvQo/f8a4nLSFDMIyD5kQMYBwROo06MQh73+TlZyZqjBNhder8ruh8xIIh6
oyrKAdN0E+rTiwDPBgXegh4CrRoeENdihncdK7JDepsGkggg3wR04I/w45+3hv2E
7cgDXNmXSd4z6WHscP7GsykZBmkUq5Sh9cdBf+iVKkIlI3Gy4HZ0x84SPHGgSS/j
/IVINNJ4/L3XY6ZL9islWAFBhyWOBq+GmpdRNqr/Dh7zegBahRko35cBVeHB0P2f
vtIjb4QJN8QdZlGqNellfzMiDBxRCK1R9ivMw0UF34he8YEx5uwckmx1oqPIhKPO
vi3rAm4zmmkwOO0FYjlZPC0314bN0nZvYdaEfZSTe4eKiOP1DIMaqRoieqkBx+Wb
Lw7NPJMjKjtgvWDLFLCt+CcU9e8qB136nmHS5iLJaxLEEmfN6z1w1h986wFgqgPd
L0XlD29dakFj0sNOa1xLh04fJzLVZrDEZV3gqfVonzFCpTtxAR7C5V6gLsF9ui+Y
4npuSMMh3hmsfqZw/r8tCt4m2E7R41W1RIeVCKgDy0qaoWkcb/GIWSntBI5duD8m
Avh5+krvZzRpR+eOC46MLF4x8PO9W6g8K9xxBaukxaerLXeG/QKpNSI5eQdkWWqb
XoTIy/I3TklCJKR4GmPYXOe3apzZ2GMQa6F5cmxsod+PZdRSZtKSmyLZ5xVWtdaw
iWNY8uU8fM/NGngkkyYTFGnsSucrN5VK6dljQRQcpne5Wks8gIALCgBfK5SFudjk
WgD+nfK0tg9gR7ay9kzEWOqiVz4uGwh3PP1jeOLOoneyMAr00n0qCXSGfU2m6bcK
g35oqnX0EYRgbTy/X4T1HlOTgP0qEXLUo56limPis6Wwlfh4FhCfjkvjbPj+mzg5
1N+fMTxADfJae1rzSyHMMZKFJieoHdAjKFnQRxs5r1LC2U1gvnWTbuUOse0toLMd
NJG8nKBLKi/Z9FA26o85N+s1gj4yO3QTfu6M9r4JfoL7oq56RpovoAgSc/TjOoU3
+XytrVqoGlz+a4PfR5TBlSJCkIs3o8Q+Y9kkY07oLNuO19ccDOEYyXjUkFviIO+o
YqMInlmu9ZK1nr71990goYVvwMqJrtc/FOFY2kWDpUgvh64cb6X6kOwvgDGGZ4lH
/QUKrgdmJwqA4qY78wGn0LWuAKPMptB/I6Z9iFCmZcwtLm/OykLSqg258U/y7yIA
zsuXZcwcQCmAQdqUBhI0ldy5w+gNqThaUMIOGdjxCapyUin05XsQhaCUMdxfCqVu
eJLDEO9iay34uz0mvrk4ZmJbAN7Jyahq4cKEReOsA/AgvHpUU1lGEpFF0z17myUY
5wiSldIMDUuYvB6UrwegfS8isvl9FgSe9lL+UJbHqoPNmHrzvGv9bhsntTtz0qWq
qbniXh8jufMKSRUs2Q4WmrWFxdGWIhPjnSo29j069B4BcCj3pgpbgTGh2mSL53aw
1HOG9DUZ6cJ26x38G7wyKOK5Jz57ZQ1uyHjMIsXj8ayppMGbLG/+HRzJtAOY1V3c
I9osRy1huoxnJ9B1/nwZ6JeTkLdZc7+QYfn7SiF0L9lQm3coL9Ck7m7HvA6pixhA
r0eYJFRpYM9QQ9kBlXnBve2ag2Y+eChW8LBcZ5PccUzBXF6h2Yl+FK4BocxYvahe
92JNk5fOOawCia+ejR15ntSakTq0HN5JGx58NOOZLITHCLqeHX0gS7gwPYmxFePN
3P5E4qxqwzM5fijMpnQQ8NvX5aCNvjbAiX+m9LLxXBrB1aieVe5U7vaokkSit3zN
esln6x7WIwhqNPDNHipIWYy7WEAM6UwIQbAR7W+6+oga9TzrofQYOFTV8K8K3C0o
PgxXXhWIi0FPoVKRs/ObPG2EOPf3vpQX7/kpcscc9/eLcv1D1pVx9iXel+wbLcVA
RN2hH0bUlxxK5qLO+jkYDVAW99FJoBYT/vf1q9TiJ0PyB8kiUzQyoPN/M8y/63gW
KLQslCk6yW86rH8cMm5Ejsilwc8TWK1tHCAilpiAnkDoscEw9cxrdMeUDvS7sphQ
3NWf11bdAKPb99EJ7dGFBPQu43Rh2ptiWXbrHGVu/S/cujU0cFNZyw5STa0+QoZo
QfKKveWa2dVri2DgH3fLwpe8975+UZ1nubrKSaxyl4ARtN7gvjoTeB1wHkh6IyDh
5JBeDsf8T995pa1Kk3QQhmTl5WgoPmLMPQG9Oupza3lf4HRPWY7j+DG83yI4uvdZ
XtK48BKvHzRxfXffHaigy9JosEPExUFcedsSbTQ+ek2ux0UFRAfJnl3I+rWtUwsN
XKJr2awuZd0T7xGEPcqMXn9hZJ0+FREJTpLo4o2ska7W3txNrJ4PhatkjOANTChH
Nd+7foSa/Q6jSEQvr1iKxGGBB928eZe53F++aUhDKtU+TXy3MpIMGHS8sIFj6OMx
mxbXeiea8sZ0j18/cwqDGe6fdYzaZm3Ks5+vhfnoFPijgTlumFDZ9XKrIv7rHG1W
YCYj08et749fDlKlGfRioo2MpfhPpRlio3sOLft2HZIdGwRLibNLsSmWgWavI7x0
67/5VxXlwU2nDkprzQgRbldMZB6V1E9ZlVtj/w15yRuzNHDfixWwuLcfWPafTTTT
+f8KuiUPsamEstCsUgfE/NS9RYslBXrbgnL+oS8j36g5ouO2GVCm8NrfDFGZMZKs
wH79YyycuVbXL7/c2RqKKvR37A+brwHZMlYLBPnZQfbf02AOWyeYMgqkWrj/I3Fu
djbgxzT/h0ZKcoVP7Lwkf0NMFZhc42pNZ0nW9szAys7CgtqhQS02COpJ7e8xfMkC
JvIDC+YaC8oth8+pr/t8X2LAona5Px/mXKNjKr373W7u5FtP/Z3GrVX0gTyiGT4C
GGQFMggtOUlXZ85R6DV/4guLkSlDowDnFSdoBGH4TZ50MkkeXaA7nyAFMJexuRlE
533qdlxez6wsRPi8wpZixJZD5BzvDD53gHj51E8av2KxRnbQW6UhNChldirsj9Tw
gY84ssK4DgZoPHhVwYYndC4pyfsPGuRUOz+oedGPB4kUhghYosTAPhNybexQY/jZ
/7gFVsdU6UD8zyIXbF/Du7R2UakZvsEQBes/v2Qt1b4r/T+hS2vA385iiZS91UF3
kcinaOp2l/P1AnO3DosRxMOWaylfQE2sEDcSCU0OQnBiQ3/kbizemSydynt2Bwpc
rWNQC718ddBFdnejSrEVJ8vrK6PbL+WQFpXCJPDr9gIkNp1YehZ55nbxvzRknGH7
1gbFQf3sXtyIPaolJaa5YNQCcjByOSjf5Oy4Lkk2hTnBfTrYzYQCYMloBED53n98
pGmFwhfqgMcBDNv3GbpCA78naM6+77HCPaKN0ELr4fZZ0pVKuMAtO7PPNKg4hOh7
1AWTCJMB2ud3uSDjMuOQRKc7m9rZFzARMjwXl7VyaRrIn44SSmCUMlPP/2RWjHpz
ZvzoZ7KfGmxW8kFth9aT5jl/evyocVzna4FQtu9+NFr32S4Ml7jdKFd3sIBfO5v7
7VoRuPPuqsQDYNs+7xkEZKYEOLw9PDMzUHPunfPUgepNA7HHlBb6Kw7YRtx852ym
cSGB5bD+wL3Gwvgat9DDzcxti9za+aHHw8qczf5dfmG7sbHBgI5NfmmyVPpvcylw
XPvVvUR3qwNDJaopUWHRxE6xKvr5yfk7ynV+MBadaPHgpoGL1MpsZkYI20u2Mrd9
7Jh6bfM0n+Q3VcigtxhECMGFIskbVgASCNZVMnV4ACg8RVjiRvnb6rWMURinbaf/
lmhN+ctYAKNVn6omVAVKNZ3KnMOAM7HeDwmaB3WMowPXDMXGGQ0j9yJzDqalVv3K
4+q08fLXNBHJ+xLp97Y70W1HsDhqYXsgvTYvHT2557s0oG1nlr/C9hAnCsW5ggmQ
Gc4Go41OUBTEmWkUyvbdpA==
`protect END_PROTECTED
