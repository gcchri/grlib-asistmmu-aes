`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iE6TysqyI2rQ1CR0P/3kCVjeffsM/Jn1I9vwG4QrEiZrR5kfsQTPP+VcqzGKAK4o
jg4FhxTAaHMtD+APDwTQL4P1tX+Ocp8aOQwOYo5/HX0918oOUP/hwTZWd8z7D0gE
DXBUvyyQl35Ftf508Kh5MHnClGeEFt3nOw5pVQMdqtzarZePC1j0KPx1HRc/nTMc
tO0ou9LkwCxPHRVG1xTYy/v010Q0d1MvPeIOkO2UdNkBtt1leo4KA2cpQMqsgzmn
J/QVz81DI7A3tbRSDYGxjG2o7YXrcCARPzf/rUK53HCU/j5ZomxmOYQg3dn6pDz9
lvpD5cS9xe+q0/rcSXf8/7DEW72oDrLJGunl+Xm5e4RtSzOLRqEktc+KsI7xgK4t
ektbxq4nlItDZxePmTvejaRZ+C17vvQJZBNjoDPYNNNS0r9ly0tSGZlpqsYlT8R9
RJSkYj94/62+H9QucN9QYRcx8FihPc0iagqpqG48hizP6wvqnrgXdFhiKPKtgLZD
N50VqHwjliC3C3wI/QT/x8mgSLYxTMrTozM09qDKufJbcexNggWEx9AOINaEpQWG
wo3c+g+qcYMzGh1v/cElMv4s2vD4aWAqfljH0jM6Y8B2Vu3W+An0kdg8AlOwu/Zt
sTLjemv6mDYAFN8UN+A4oGzAvrvOrpIOnryrq5N/vvvXs4Qjzd9NwtG+6aqGv+0h
6GgjaGeh+TidHG8aljARr05Nfq2498TGATDx9ZSmV6n7mL2ae3KPE/tfa4gJF4gN
vQbSSUGx3PKHPefgnSPfCIkhStWP8QDTX2enhOCx2QzZufsyjv/s1oy+m5wCmXqg
KMjpS9xoQkkNPZBSJUJYj1aJQvvkaI2vTYekZokYGU6UfrGs5u1jFVky3ERbL+sc
breWJcjGKxHb2xuJpJobTy1AV3IoWv5fq9Fgvl4lwbOOQlxwipcmanFEv/a/h+2h
opTvc+D8TfRTnHN1OzVseKM2KCjVYJ+PuKDHvPlyMHgDcXVDrZcb4+pUKSy2HRrG
QBQ98P8L50SI4gTRKFzmMHAIdKDFUwv7xLboILprOwz0oyiV8BrGGgfD+IaMEk23
+j1/ZiZONEnStI/F74p9t7bMM8TiHwgCmrwFpV3vTRMJy/Xrg+TVPrjcHztNUGAI
fCwZq+KBeDxLU/itacAhoyAxrr/LpNh7h5QxdIc7pykqqGJX6WUDpIw3pYpMmPF/
V5R1k1dq1BGfxGk4jE3Q1j14s84+wGom/AV9alx9eeY506tyUrqWIKx3rqz0Zn2+
y0ZCwuRLxIcuBEZxQ3D+9+V7Z634Q7HhupKu1tOyamM/YPXqjaHUWiCEEuK1y6B8
VMv4kLRbcYK78ekNS92gq3YoyBv0n2mUqxF3PkNrGTVGSQ1mJ5knreqQ2rlO7gk1
mYHKESkMK31YfHQH3f7EgxQS0Xxygr4BU5y23uwjINQk4zz8+nY8INqWnFAJH9Op
tPLGWbzn2v7dhJZu1DopLmrAzhTmTvXb2HzoI2FhsnTLEqIB088Mi0sYAN+0CltR
NVlwLHavmToO9FuY1/eSO+1IOk+s5JTH79bTqzlVsrtJdWZ0lrRaSKUOIB0WLzr0
t99VlXCxUGgJA7EZp3K7VMHnPxlK9BHAPo4rml6/jkMZq274h3cJTmQ87G6RrusG
Zcb1hddP/fCgwSblzNRXdTnaXgvxCUd/LpYKuPD1Kto33LMcyUPgvPGJhjXaCYGm
E/Wp0J1q9kS/rVx2Ti3TfhrV8ffXFucHaSkBdkLxFZRe25iy3Hs8A3FNav7qDqso
NVvJC8UoaF65UDGkCFZ9aozYQvXjwWQL06zLmVbmU4Kz/t9+hkBLreVcKx+VuHmE
ViG1NXvzHxykdDq9iHHVcrOJLuMkrWRCXUMMZ1p47Wr3qmQq2CPEsikFICAjjbBc
EI7F1nzMqAou0ZucaGeG8RB0h9g9NQ8Awhyj0InrvSNCFuFQE0dWkWkKr6Z3J2O2
lub+7bSrv8RGe4ZQ/YlcVu9KjzTkfz7aSWOZVi+goPQ0bWCG4hYreJPdprwD6JR2
9rYYtjPw5PE5Gfok9vPgcF6Vkl+nOPDEzXzQlCqjkNWNk40XidkhHQgHdaSUx91S
HYoU8A2dVwlfiAn2fQnEOGuNPhgspKlBfwqC6lcw5a6tmjuQ3KXL4T4Y+sKnDyGN
iQfqCPVpBWH1ZAdDdVq458cJXMrya7n7zgA9MkiUW3fGle5ZpUm85XycTDpPsXUZ
fcuuslKCSlWukDggNvGMqKH+YEwbj8BW4PFR68Ir90d4qvEttPOFfQYyTc7MOmPr
gDPeT8uzOgY5Gp7KWzOLg6RZ9s5sf6DBEiNSnXc0S+NYBXO6YEdN8gvGbAeBZx6F
7y68OteGCXoA6xuGRsi3PLXiYyT+h3JfexLIZ0jA3gis9rIgV9APZFu+Ik7BujmM
ONiAmiCREhTyFQ91+WD5vkwhI/f/vQDa/9Lf1K6Q1QIaBqsgSH98dZbl1TgY/wIr
SUDh6R/EBWG5+e+F3/y8eCgUnMOrq7Eo7ocJx1fZGK84BquhKL0h68fFZhrSwZPY
HfZsSotZ0uo9nuX5AxVB7d+VcqOa/lBjjZRsaqNGNMjfwxUnHhM/uLlHaUQIdS6B
Lowwx8AyPmyG1ClOcbC+9f+Q6an12OQvYpX5mkVZZ9HqEjbAc2VVZ24LIU95SpeL
hmwiNm6M7uW4vj2IifV/Yc/+KsU7RwPq0fHGSvP0F0Ic6H2Aj3mSIzqeVjuaQ70W
E6zdmJc0Xg1nx72HwKxyIQ==
`protect END_PROTECTED
