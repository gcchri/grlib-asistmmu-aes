`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A03hChcmWvUXAXQv7NQ1JMt/rX7bPXgPxjCmuszRlpdcrOk5SRMDPhYg6/4GUgyZ
WkKRCl6F/dB2w54PZ92ROyXLnsrBENOX1ZIigWijtEJDxTX/GFtxJLdU2lojmcz4
B10uHrG1lNkOKjvhboJjFwFDc2wvtNeLHLGX7rqSTqOmaOrWXyf/W0jeY/5uudKx
RfbTt+DTCIznz+9JsAa3WJBUZ7VujjjXxd90T1KrR4jqCbrBrBEvMCBv3zx39/pc
MZTPguEQA8SKDjKe4VbFgKEt+91S+HOkL5SvwkDqNlMl1jonoygIM/QWDK4F6I0w
SNJscf3QoRjGuKHsO8ZFy9P0xXnYjD2FMg1tFN60iOgLFr8ANrSU57i98nGRiArW
2pan6UTT1G/cnaWfiVr54O/XKp0MHwBVRH+rSrvmReJDmf3nBzkUremPEOMzD5XV
SWwpAp+QQrTs6Lhmd2TlJwSVjJv/P0o6C37XDdzWC+cADuBro+NvbU7wyvr6fg2x
aBm7oagEcsk53JcHUCB+8wmYiNV2rwccMeUm0n+Y9Ha3UV8slNRrP/miBfUXFFyC
OIv8HosB8X3SY4xC1ZJ5q0osQK3CxKslhLNTJhYa9r9zJQ2S47gnzbNRej5kOU8i
I62n6qUdmRAq0DbDnuLiH3EsKK+nnbzzkYOhlc2CzkdQBQv+uzYUqX67gDMh6ECV
77HCPClNoovkNh/wTCkzgL0n7VYm1AdizLbRDadEcJvhuwOXXXuGfUOAKiRUvoeO
FKSlAXbkkCbwr8XXkK+xOQ==
`protect END_PROTECTED
