`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtyYdzRFEyGbNhdaUF+0WSOxlXTic1JdD1NZ5QmMnSD4/yFz8oIzsUv7Srg1attN
VZmgPkC2VGnubqJEV7lYGy2N5SznqbmP8LXosg2mzgqAjfxWy90KdbOeMydo4Oq2
ii9iHIMvxGT80YbxsVviHvsmJegp5S209Xh7xNybl9XBCsglgaczlCdp7w1/Wfdx
Lni+aS25XH21XcJ1GrTO++9G7E/ESdoMJaGl5Tkr+eHZBIorZ3nC6dHI+Y6zpVay
mgEHIN/9d9x16dsIiQmTSVsEy/TPH14WfXvsc3uTnM4Gkrcw6dZ7O30jXcCes2MB
+kI4FkWxFmv50jkZMX5LLgMeZ2fUmqv4MdE7FrRQqlT7VXGeqhc0VUyO555tbyko
6G2Gks91wN18JjSnrIRImiJdpLtHCbxGbgUbX4cfatjNe2/X4P+mMRg6qMbIzxv5
R53ah5D5yqYme5UMHHGeSiVWu0UGf2sKWFkbP8ik+5Vze7wev0x8QWiBVWlssvsj
`protect END_PROTECTED
