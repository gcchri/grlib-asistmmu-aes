`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qujbf5WuzKKQ/tAltwA7xt51sya4wX52RphKK/lUK2aZzmO/l7mLiojqkj+LkLK7
y2LQ4CORNlER89xIIxG+z4IqGfvnntpvAaUUl/y5yzJgSCdEuCwWKv9am16tyTdV
xskumDJXKJBn6mLxb+dnkLAAPn/N71gKCi6GPF9rs07P9yTqLCM3KFP+6+2bJc0u
fTJwF/eQ80ounn+bLr3bbiH+X/UvpFu71zs0CZ6Sy7Jgey++DQ+md5DkSCdYRReb
rLdOCudydpiF0ImxcIJWTJs4fzQMLjL8KnmUyFbZuzyUGHrrI2v5jX0Zj57WiTV2
dSiLrdYleHsVAydMK5QilA==
`protect END_PROTECTED
