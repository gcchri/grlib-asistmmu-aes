`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPgmaOpPafpFKFGoqcCnFtuasQ1GpMUrc5ZNSVfjZFDUYuFTS12WkNoMt4LME+ps
tAb535E1FmIS6EexRNtO8ib4UNcndF1Yjyr0ULNhLcqNPMqbSJptT5BuoEOgkoOM
GWU83dd5/A3ZNzBd2zezEb6IFB9Dy5fr24KckE7c7yVhuM0/gwUkHnIoUPfEc7EB
9x4WY98sd0fg8zt7autqrqIhyWmQtjmRrTC6BBta1h4BLTZmT72f4iTO65MVUmnB
vfBTeGwsr/MWsM2zB+F9nA==
`protect END_PROTECTED
