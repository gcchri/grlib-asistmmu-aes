`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJlnHSAUIoWHNaHtqi3biubsRtbIOHWhCMi0VTgabY0b4F08ZqZW6vRzl506ypL+
VpqmTJJ/CvQKvK1MEFeWfrM9eET22oTkDcJogLKLiWAOLshJomXaXuRy5YyFsxgw
BGGohoOGkmlQpRMSHirSurMQaI1IN+dwt0jtoMRkJ0CUwHMMqvmCzccBzltsEZkT
RVx9+cBkOK/2yW4iE46r3vIYpWcFMvUitIdCe5XzXAssn2ZNRLpdck8/yLEbfh+V
vmflP1dqk9XKHIZ7oThaS8MsrJUKBEdWBFv4GpG4gyhs4gINPuhPDJf6CZtWp2F9
xDt/3vxxnrY8k/pD5H7FXhRuL5ImQks4gFBet7kwDE5OVPUbG3FchB/98crMvTZV
eWfbcw4r2WODUggt7DcqW/2Pfb/Mwg14RDpBaBYrARlHkf4J3Jy9I7wdkjNw3TtC
PS6mRLtHju9OQUEv2n2K/oW+ijKjjr/yS8FZd8VOBeuZV94nGa7HJ52MWk9AQSO/
nHTBbfRq4AO67zVdFjBSqaG0hea1+vNGKIwjBs7i1bU=
`protect END_PROTECTED
