`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCj7XJWglDd7ugY+JHUfCgs1NbMeV9g8HD4QZgHPqWoIPYnSFuwq3cfi6R7WBkrt
hDaqQgt5vgKGhIhE51mEr+3WwNFg2cFMN93XrDNVP+DftXKdiIhJ/TBqC6Bz32fE
ldedzG/JXQeR/3Q14mAL3rYPiQQIwIcxCSxJcEXhIoQCJll/Kvoo/YwQyp9idvo1
ni7OCQvyoo7lkVC41EBFNckFx1KkzNgM3EYVxQmLJztcE1MUuR0sBrpIVpWUqmu7
F0Sp7ohW3VyOUY+DKqC17n6dN43igO6/vat5LfB60GVkDlHZTjhsmvp5uqbr3Pzb
UPeyW9m9lRvy9jn0HjhvNyx6bXw/oWmnGrg2DCn01cRLBRG9vwvOMqxEv0BvyBHF
1PWI3VWLfJUwHFsuD1BJgk4ncomruUCR4piypgUFLLix1xmHO/mRZ6DUSsY2ZSqK
2qH+lPkWoSaCUANNub/3+vKlKwpwXjvGAGUBWjmwFgiQpI3oT3ypVT607HyT1MxL
sLSx+L4+g/kyHjYahb6YoVgEEn4GqVHYkDuGeEYKyDU4xJqLbba0Nzvx1UjY1z7+
8wtTOSN1mazcGytlJAa2eEsQmuy0bmWPmEOBk1/BI3p+Ijq7jFMQrOFItJmuPgzi
Q5OUcNN1T9o8Hj5jV/XLwvU7wU5CqPafEus4K3GUrYmddR3/3j73J7K7vNNqV/hq
kutTpf6bOpd2QIPahV94YvRPTkME4d6N/LGbUtnjpSeJIVnSU5+RL+VXQwyy1auN
q1MIOhEWO6FuzePTRQzWcwlWQoKzfB1jrfeIRkl69/Ih//6mlyK5REGvyB1p3bDa
6Ghu9P/BegXxwxR8Gj1AQk25OPfZhTMViMLXZeuLo3Y6o16Wtp2PPkr5iXgtDud4
6Mm6JILutF+Arbz8gUWg1w==
`protect END_PROTECTED
