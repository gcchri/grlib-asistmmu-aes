`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vM9wUJ6zF1mUSEq27ZBi9/F95rPRW04wVJ3kIHkf9ibIwiYsr3Cd4ztNcd/yWoQG
nUCd046RRA041YD53KFhS54iJ6zy+CdFgJeB4BrMlyOBJXVxzDsQRph7JbXU6cIm
3BfPtBvuMF22beToNyUqrCeQNfsat7i8vShQ+Ibstx7QJBGWIQDoe3itxv4XcApZ
PxBecgRp+BZg5vyPi0+IYc8LxGkUvcEVgsa3Tn3lz29dmyU1EcAcaltKl7EBSCKJ
kz5QDoG7HdjodaPqkT3+ao3hkIEGzyMXz/h85BLdSjGRLaapugnuKKwatv3Fd7Y1
CI+lO1/7xDzHODFqo+2iFwJACcCF+2gFq8xCq7tCAr9c6SdT6SJgAvUakTO0dY1V
AyZYfbS17B/V9nDQLFc9CXMc4ExURXt0lDzvnrxAfpGNbqwB8bnyc8ZdDFt0+qob
W8DfwbDiPKczoNf9ExJpX70+EJnRTnw8ctarf3WuNR6WpnG6zhvW4MTFO4wDcIV2
dnbyVkdIhBAxKL5rygBV9DK3p+6fCpTV8vfZ/9NKKyXY1rkUcjo+r9KAheWVit+p
3oQQhOKGXy9LsS3YsMttjhDYvoT/rMFVEuzJsT9yvakj671Bk3lQ8x56ZNxqnDqw
YhlLxr29FUpCQDTjWEiCjLR49vWvBjSO/Xq+XoQwhB9wIMJHYWKxiI6r9jvt8hb7
Th/eQSC5gYmCs61052vLJdFVvuPmRz62LdLFGQ0k8dVzIw8Z+4Fp/KPUHBv6CJo6
C8usczFKi93KGtr8L3AnKHLkEHiB5o9it5a+r1b++9B3CxwLJS03fsvWUe8fSqhE
MvmygSOhiR6jfi9t5bFGKn8d7WVnRYsbQl3xXfZrURG3yJWrzydWSHPbO+vOpeMz
u+03DX58wWHMWeAsFAtD/upkauluhNTeIG8+3O62qwmsjTCtJ9Cp5jxRGG6R174X
eVJ79HjvF6U5/lpUMYBVyC5Gk7mdcC9FLDXSmUeUzhLc4hHr9NfjEZk6br2+FqFs
YKUytYn4BmiYRAqhm/XmTJ0oiiAHtDqCQezxufY9yR5eNx8sdzPclr4ValOFdAhD
OCjR1FnsgWf7atbJgeFUzr6VCs8TVnBQT0oRH4F9OiY=
`protect END_PROTECTED
