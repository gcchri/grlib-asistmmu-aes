`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7/Q2m5s4Ew3AxqXEkrAOqUxJAfcZj/pQuRzWUBGtKcYTKiBEUfVixDmU3JEUpMa
2SZ40iUWjQaJh0RhZl548Rkp34XGR0n8cvMkM6VSAK1SJ9CXI1mNMsmp7eDkRyOT
dnbrxtJW6V1gKMzTeAKujxh+C0CXqPwe4kfAaNHucWL4N0XxF5BPJK99vRGO5iYi
Rik8rO02qXxRpUQAHgEG/Xt7V9Sc5thVX0s8lj7y7hP2d2VtwyY96g60ZVU10nD8
2XmTnq83+UegDbTA8WDXJBAmzZejUwtMixrghE8W5z2Hvw7U3hW22eGZxBw3F191
xRoyLczuQjY64ItEpl4RyYVlfJ+gbAD7w3P3e6SxzwpzVL9FZtNaPdwhO6p9fKnu
`protect END_PROTECTED
