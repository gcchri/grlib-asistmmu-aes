`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+8XSRZ+15MmDQujx/xRM6CPhWcwFJmv942Elkpta6F5eKAchpqn8cgLp7VLMkIt
k0H62BytchuMHmaVg8RunTHyIn72Xa0CEcAcVy0e8Dp5znr3V3wxCLDGJ7rckKSG
954wmG6rBOhwBW993SPcue5UpUeeQwUfsfYYPSpMgyYaKd10x/g35e1ZPVRMOOu5
zzB+GSeFBRB8o9khTMAhlRhOfd5rOOAis6XKvscvCdVvKRZtPVl8pP1K9Xc3TZJh
72ZR3OudMEZrVxwEIYelnTTnwXJgpmods+qiLz2u7Upsyj6HUWJeI21losdzBLMj
xVFD5USijk+SeHOdXVPeLj4Sj0RtI/KRcDXlAGZOuQHIdNka+fvPgBcA7RwY30pX
/gt/cjwaBtFOnyGy/+jDJOw2LZ5Vji2YAFt9GfqwVBYb3sDtdWjya8cBqRaHMmpo
yiUY+2cTTQNZMunXlFVyYhDZGns9Vya0qd9jbkE9dmez3eDG35TRreOPXKhdZuey
nwtITz4ckhELCm5P50hCw9PYbluDxuMuG5zHAFQSUKp1QyjsVjT4AS7nT5a6zlbd
WNL135y5xWM+7LXfE1mUM6cmlhKXI0sBEulXx5MJnCc=
`protect END_PROTECTED
