`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+mNSy2WF16c+u4ZmUr6VYp/EJwXEy2tB2EP9Q26VTWlGAbR4QCv6ebZpncjHswO
jYqaCLEhY1KvhrQWQOos4c8vgSjbjAoaoB1aLHFypf/irKsihGOfKL/sNxeF9na5
5GXk2WX7OeXwIXaORqIOZh9eIq2Z6I7DsJtybRi3J9mcvYc6MRig8oO+01aV32L3
dFgXLPu6u3VNJzVeMT/7UI/hHS35Bwbwn+oKDY+SqlaCUHDjOGcve25lPRknqgHk
ImwM4L5FB9buFnj2U4hXduj9eFJFfmbfElwR9dXeygmGsY0viD3Tshfir7EBw+fg
x3w/yOXK3QZpDrmkqXb7do0prKfaEis2VKE0kGDmmgZxZ3vhnod3Pm+NsJKEvG6+
OIGk4EKhz9Mv7S7gNMFYiWFLQiwfiXbzQC0ienZzhGjhkB1p8yNVoPrGb4TdRaF1
cq1y4drBEUbmZKe+xO/6XFZ5RPTdDvM0CuPLyZT5sPsdtbIR7S3G5trBQnNWCpfN
8KuLhVYPktJLCLBZuV2pOJpso7YD77dW5lBmjkn54/AzLWzK2sockPZY7mLy9Zih
ZsUUxHBlAr7gX4BEY+NoDLj6talj2rnrouC/08At+/eakP4iVMg7yTlUp3+q9Y6N
`protect END_PROTECTED
