`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RBNGbSjyXm2MhxR+3rcR039Zs12YATX8Dpz10u0q4KfUF+QFqYbSdzl8g/+Hg8B1
/rD9JB3wpbXxxFGvxmNft7v1spyeQ7J04fXg1CkPdAHQp1WUBks64LGvWKLBblEa
dfdwLGDT0wNgTYjPmOVC05zF2pIQt+jV+HW56HkMhprbQOTcEuzJoMBTr8M+gd6R
t2E3hCcSUeYHWuLDcKWebZO4o92t4bhNzmqNzDvfQDylcauEFxzr5BsqJruPL10s
W+Te6lEdm6flhYNi1LW/hg==
`protect END_PROTECTED
