`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nt/WQaaTrfTy9PXFkIoeBq30PLlw84XzWSQaeqjd1dyvLsZ08sXovRLFTDQfmwe4
KE8/jH2AHgJU/Va1HkzYi+TKLvJPj0eyBEkd7nm38oEY3VUCMpAF5DXatt7BrKdq
jO9D5QXEuLaHMpGCU4FxNNZF04HGPFiwOWVa/5ug0r76j7liA4uXrkFjzFZiyxXa
iwgBdxtmr+eli5Y19LB9q41cuJxdq3kzVD58rpvdNlrzRwzf7z/2I0rA/1U28u4s
ZgWlAcPx4b9M8tKFLuf/TU6QrQ9TFSoOVP/mEe9bhlDoqrrqb47zEIyAzjf2tc4O
4cr7Vgen+h9e9jFiX5mD5qN3LsCTSi5VxbhinsFnwf1TeMmqANiYX0/BqDB9E/fO
ynawj4BG1gPBIxBi5BP7bIuilurdIuBckpqWz8QN3SFGNDIFmBm4hv+biaSGEbUS
JNgay8uDT3u3hXMEdgVKyy78fDq0zpLjFvJXtQ4pvpMS8HOIdk2kNVOVjLwp/skV
Y38XBzKNpp5plg5b94WutHHWBrJAElKGHG7dNqhFO0bMvwMH7WtfZdXX6vNfONri
c/vMX3YhaKCdhQSTEximE5J55mJ3SqF+zVGG3mPZhkBYlH+zrPLuIyHz2/XoX0p5
NYNbqXk6YqYkAbX8Ni/T8nujacakAWRWIBi3gWM630GGdwCQ3n6zwCKw3Fr1UMZX
LjC/t7McYets/xLK0SncjVrskDF9gAyFQyC2lhZPtdoGZ6JqHKfIzjcemyeBj5Iw
v9kWRWCWVUoD7ct+XP7SumxMSrWDUCHhbr+9l3biD1/7FSij/eFMvObLBzutRQEJ
GA88gTk9u5nvjR2anLOcmbT75EZV8rR0PNcht46DJvCTVZ6RZpc6ogkAhxeyyGjS
R4LuyD24m+WDJejS+ziOV8dydxdhM8xRXC9BPhdn4NQo8ByPROscMQTWPO5fdqYo
afEVw9NVXAmCW+ry2lxQ3vIJ5Ejctl8ttfMiYreorllP28GaNSyI5befb0AwyVpD
Mz/xTVSlQuPNWz8NilVFCj3BYOqM9S5t52C+DgF19ewTSYLBdZ7ofnk/I+srKH0B
yDS6HCEUpmZR4PAHnNbkIGApuNsW1jNnig56LS9jXs/TT2DEi4xM5vfZB5C5jpzB
Y4ZoYoVj+h3my8baQy3PahrFakyw0sd2u9H1ZqJqt9q1wwrAqr+gtg8SFydNGKYD
Zlxmxotn2aGoj1/g4qrVtFTheZcOkxm16CNtAnF1HySfm+67wEybBY6pr6piJFTh
2Tpqr5ju9Y1X+FYeaH92wDJ+5NLfU3hwy0q2SFP8q4LSSojlleUbB3YFmujuG3hB
3LiD+mMVFso/AHbxxPCv2KDXWr3j4J8xoaFm3ND9d9YyLRiZOGyedwCadoU/1eql
xUVxAbnszB1vCHwLFAxxNNLnjGKVXsgcfLo8P2LGdXaVKIRlCsWVpcvnj1i1uOgi
D68ChQZ73Xld+SvLXrQ+IG0mnnsKitfBJiGklBjgriNuC79NjPiWPcf24SBxRbT4
2BkgLCed4vlfoiq84NmsDp6+Sonze3tAitl2p1oh+F/a1yY/8E8HB/XSYLw9J9EL
1WdCEkL6REtpqhR/Kvfquh2/7BIAKZPXUIqYySnpGJP5HVpPq9j4tJvXIVwXsL/g
yBnuce40TKxipV2hB8ONhCuGAFquoW1iGtEzakK87pIA4zb1eDfZD64PXa2xet5n
3vZU4zjS95O0kQx3KD+pkEbe81MPLZgMUa8SiAbj0Y8a7SsljPvNCoSLSpWCvkZn
3I1UFm87Yi5GoIdlAaQS0GaMxQfwHGu7hyFirS4ueW5l/pZwhU5V1GbH422Tj93i
mOQwksIr6S1E+WgBxGCGZFpjuRFhCeX45GNxK4ErfeRNUQ+0kNo7TK+eCDSpYttA
0LVcgbH+nX8oxQ88Qg1ja1/xuD/OTqkvicjIlFngfYRQ6NP7aUrWxx/U0b8pbEAP
to9DXbjq7c3uv/9dqVGwUsrumxCY9q1JlyzO0TedZKdlpRQrYNk4fvl3iFKQJyzs
RxiPgUT7EU+qYvas2Qjn3ccHeTdUQYS8QuNKHFPAWwCQgcAkuC1MxIlCKtSyzP0G
SYZnk2t2pdRm7XD/A5o/pmHrGyhe1EChY1eGXjg1YQrCWwXjscjXhZ4pVxmGlh8p
7cPT1xk+7S0NEZp+US9qY/x8113bNPKtcI3DSkk4JhM9LtfTth7sV6r8Hbx9YdxV
zzOw/rlPoGjPcwLWgldyT2dequKT53K20J5NDxw/pmkAsEiWJCIhg3moABbNWa+d
pQS2dWZeqozjiaGug0oblaXC+Wc8kFcjLb99uxVT/LjYhfdojNXVZ+/TlnAZsFS8
ndfVYejA9elZrO96xr2ZuPq+l5VqBr4ZU1kl83x/JRS7yu595AdBkBkfm8CoI7C3
tliml+RD6Vdjb4NsoX2a78uac+y/nOQcv66HhROw1Ud/i1mF2fxitmIMsE9SNLdY
kNbalaRA0Myk03B60uT7nF69xp5PvE0d2yWHK4GIl1oDbppx7WTqpjd94vTIQQ7p
MyWBONbZfLFvvB0Aq8FFOxKq8fjJ0VKTyg2TGDLgYLaMqXbAYiBwVTU9IjXYkq2p
GCZLCpn6TzRcCCkSm9I4xHC7NrAJu3aIMs4EecB9P6h4ON6KTEgO2pzoqCoUrVID
SFOAShVnYEyn/q9aejMSG1JmcF8A7Gj0cPoL0abgSuvKe6QN7s1utHNWRcjCLfr5
Da3kEM6ij75z4iIBCA0Mwkpof3mSm+XRFcnmIdzzKmX0vpsYrXhYHX3bkpX9DCuk
ZBKNb4JWuBWbGNLj5/SmBFzBggXMP1cRd3uqMsQDBiwHGfj65S2eGjqIawiVWAUK
lxkypPSn5bm/TRE73RzxXNDfrFP26U/gpsnvFsd/uKLkLIgB0YGfNuPRVLtJOw8i
FUb4KY26WxaMyAiH44j5+8ao+4nngoYjvRgeeOEf8aiknYbMERyA2fhXbKJjJ8c5
JypGtAsvdtE4kX+0Eq7pSngwhRfoMjS4x92fWl7kXZFBl+5tx1K+y0GRoP+QRo5F
JJJZtrdyC4U9ahQxI6tWpBtAGt8KxdMlnJAziC11Pos=
`protect END_PROTECTED
