`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MK+mM36n3WN4EQqL/SrDo72N3Ywv70oZKBHhgvpfjtvFdHVCOxWCMDaBHODdwoZB
mbzpEl4OLWRolGjNFNIe+nrDolGkVuBQo7kIoHxZOXp+Zvy2iVRyYryU43bW0JAk
csR3D2JGP+j1w48jGi330wLMgDfkUs07bCWmy47pQBOOpb1I9QTR1ZesfxtADC50
k8VcXUfyIutzRnceGdPMWtzMe8UgBpYEPJ2Xar6I97/BOB8v6hO+Hp4XUzB+fRjQ
UI9MSYMuB/ktSBBkMP3JdnMH2Kr4dh4YjTNP6rC5FeWylxuxsy3OTHRUz/o0Lb8q
AIsvUHjR+Dfo7U7eQrbcZDLuGrULPdSsSHraosE582X1xSPlIz3qzyUtYQA1Mu3j
PQq7bGWtKmlHrzB6jasZgQ==
`protect END_PROTECTED
