`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
666iza5TlK7w6mTvnmhiUYA0REktGJNar2mObTmhrsx1mFa9d7ZO+nl8m+XC1GSs
FZepSwGGvrrfF3gNNKhFKf9tIUs4niJHr8kWKmGN/CAF6MACqxkZgzfQscXW/eM9
AQxWfoxfyruwkK1UO1vXuZc2OneNfLCa712kDmk9uXb0rrmOMe/qcEhR/QIdaQL/
negtRUDULegR+AVQg8KOO3EoEOpWaPPqFfXTadF9JHp37fwDjkgpQ99olFtXTDF/
NLYIoCw/lQhb6rXOy4OxkMinfn1IkXibWOrkGL6VcOuTqJEF2fcoDh1ALHjj6coQ
TBxso/aYqEPfh/jJet0+T2AYK7jha0jC9Nsw0BY5cr9X0tMWa8HWldMVfbTqAm+i
3PliSFLZMFdmDr2CbOo5GRujK2GXsrVgCBSU/9t8mIUVYm0+C2hpcrbSLlqvdCXx
w/Ux0YnRKZuKf/vJzTVvOrZ1cdGS19mN7dcp2VVMC6e+3l6VLSMM5EOUXCbe92PO
ZcMqJX1NSIHzyvwKf8bQNPsjQy65oNlbQOdY00HkldvdVrokU5ssD9F5ftlVWAd+
3GSDnXOfmgHgUrqJaZ8MForP+Ar6exw2lwUCPpp/J92J+0+jwCNuA6G3fQ7nhH/L
wUlv00bsp5HNVPQUwlfRviM1HSZM2C2Mu0k9wnHM1WzpWeFGoSzLvE31gmc5AvEH
9c2YrT8MMdZG/ZA+bQquMzcNMdIojDsI+BDV7L1wnPA=
`protect END_PROTECTED
