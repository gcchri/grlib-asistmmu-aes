`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3gIFzX3ojmYGnR4D7+CzJ8oPW0hkoWi598WiZ0JGPq0UtBM5F2p+WEA/WXo+Jt6e
Tc/ARGe77DGKaMmOMuUyG3VQcBwZTaCd2FzT2NmHdBOtAFjuU7WBiVJFc76bYLnQ
C9ilSnZgat+hD1p/pgOnfwntSypnX6RtGOBP1ZmQNgM3z5Li+0RCuQNtsjc/b5a2
NVXmMQrkx4NvaSmpqtKwpbr1tij6jBzCpTWa2ggIwbCkO6kxbfGp7Al81cMl8crd
tX3iwsbDCY8g+qWD5LSprD4OMF8xnSRwJijMHMX+CqpxLHKUu/A76ouYbK271sV2
skycS4e5gzhRvDIX7eaajrKMsVEfNpSjhctvC5Vcp2x7kFDr/YbfZxyxHtBmOnvo
fIB1Xp0nlNKo4kbHP/aMi7O5lVe9HlPGwg2YeJ7HXcfRuSXyg0/uZ2cT5gcmlCho
`protect END_PROTECTED
