`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNlCW2Z643ZcHg/Ak81WyfMjPVbvuzLl8W3A0SlDFOAkLp+AUZbRYrYscagOuC1V
HvaoHXaG1dtX2GbQojcy6mhZsU7rs0Qtj5GXgxdt4QbtRlnwBg5CihnfegWoK6pI
RW9KtHLR5I5X2TMVj3wrVw+JZousE100aqQm70omw8EeUHZPcV1qcyzG7/I7MW/w
3/TH0EuWcdJVDcadkhrf68cn3G33J7S7Hautcve00Q7ZONdForNJ+qlSoXMm8+Gi
HLFiGGCztsv+u2HLxG7hcOOX4gDi20xQk6kTLnZqLgGj8YWLni1RCZ6GL3B5ODXQ
4XmaCQWbj29LHxdlIMLpc3ZTpjRYjrruJH/HSefFdCpYMPVtovTpUpwq/grEMlOy
lpRxmVNuZuoYPB6JHTuqjU1/SmvvFbf4iQKojSESOcODRNvJ6B+PBXEBAifPUAAi
cHT0RCQarLvFis4EsjL0sWapbkuvs0Xj10tZBu2hONQ=
`protect END_PROTECTED
