`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TU2TPRVDvhkrRd30eCD2//Bcfr2YVyQLgXfo13nd2JPIIyYwvXCKevV0byfVYYSr
zqFpZZzSCt12YQbdDV4rDFUZgII7ZUqZ06OeCj4jqeZWV+c0SNQw27ycUapC8F4j
ZskMSQY+QSRHYurFrwZK4vTEVHRwjHTBvBAthcwyGd4R764mMGzEG1p9GZ4rSkqa
//iwVnyL0qN3N4FexEWi54YBdY/I4Zk1D0WHEd3ncSUHB9XHnviz44TQ41Sa5USu
HoVcOL+JJ5cRcrE90AEluvaFO/hK+h9rfRmcd7d4KgH/6Y2+pGOQRQWrD7XqUwla
RFlBVoK2q6YQh+rILdXZax8BSZIH9FDJ7CTTqDJ35d4kuDIpY5ZAR/jpVby8Sqgu
zqFfTYCDN61MAdhqIMKrLORi2HBK/ldLvuOyfxeadRaTp1l1CznNlvaVrdV+K+ut
CFe6Ploc//ntOhsodw6l8GeJdqySMQ2PqNU3lN5J1fnuL9B2PPEMpoxGwnkEtyfm
3FcVN/OkfUwvVDKoXKAnsj3HO7K3qDU/fw2ldfnW03g3UgtPqY39Ja2ejFrGuSGO
U8Lv0d8SMFTtuAyKkhNJvtBKRlR/ZTkaMmFYB+F7ZKWHrANZP/2LzmFmGpVndDqm
d0X55TwEVPSdy0RT/KwOWI2FR7PoIi8AdkIy9BIn2J9eE9fV0rbB1paLS0xkkfIe
OP3kcUNe9VpnmnUGDwCI3Q==
`protect END_PROTECTED
