`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BF34WAqIZ+NCF1uDogsXKr/TVQvoRXJKNrf5mQ0U0xch9hkvgBeS3YEh2lExz+pS
GahIPYKF1HIFsiw1eoUGwc1o4BPCkDRWu5Ymk5XUqVBSiyrzifitGpSPb6Rw4UPO
dTdtXEZ4HMTNkc5o5MagjPLWHnKcws1mayR/c4Tg7orzTm1Nubjrp6w7ndTcKzzK
9EkMArR1d1wSPXPK4LePjCNPAncXB3GsmqMe7iJumMRug9d1BScY80EASCjTgaS0
t4kGO5WpV/wyKqqXzyMBWOuPungl0trXvSglOD0yq1Y=
`protect END_PROTECTED
