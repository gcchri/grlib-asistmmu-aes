`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpetWmPZ2ax2oG1iU+JwAw4GkV6tqJF6KVm+q5JZLyD4lODubYFTqGhAIag1dPZk
+8SCuU/sEonOq0wtDZmKssTaBqfm8+TuTT/4rEZR8+qQWgJqmALju6WHLUNmuePo
RCc9PFTGD8CNJPb2SLGGvxfb4s7I5eLl55bVOil2z+HwVadF+StYcUjkK6p8VlBG
dke/2K2ZRgjxWvwZT0U6gY1Fa8IKtNONxV8OpyRzfGuUxbjRxMnMyQZ3uN5fWFsl
gKd3V3MKNc6zOqbpg3llh+z+RR9ymgnQfDilu684cPPdDiICQ7PPiWSd4h94eNUm
H7dZV0xmNKIZXJltKDUwTvWAi2D67ED9LohKzzRHRyCwD3uBf3RWyqN1P3/N9F5o
5BMgaEF1lU76P27j2JDrbvNayQPjz32uP3jfrJneTeWgTwINhN2n2dwLc9b8pnwe
tEp9D5+W/sXs8cP0xVPtZ0yjFTXQDCjIhdjAoG2XMXGhX80hdNo2rDZTcdLIVEN0
4HQPMOXqMZ235BDRUI+k2njQ2YFhKAGtxMw18gXtr4F/+fclVVCR+SgaChCYJAcB
`protect END_PROTECTED
