`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wBQy+jTQj0S+iV5MNF3L/tZcM6GLRlGPPNm5OJ/z874vAZCnk/7iKHssFnk4vO8i
Qr9ONW/qeF6481wilaLt4OsU3lvBclsXJpGfCmnKoo/s9BBsuPO/eLh8rFUju/xr
8RWbLwag2cXFw6+P8fwP0BBGmBPmLmxOmCThR08P+7ek/qFvZ+1nnmQA7/QQoDoE
GCUVa2qnmFIRr94R+j3lc9UAeazfk5GzDHmciPhVJ2xeJtnDvB534nbHV2a7zExH
rde8d4C2VfDhL5hLdnTtptgNhSxL3TDKVhizXTCJyWfnofPF+r2lwY1D4yyRulEF
VP2YXrsbNIrhTlwL8lLJXsxY+qONB1fSvTnZFV27g9wAU9Vx/TNNKvWGcGO8gMSA
lSShntlBjQ25TVpPsEkHpoUEa3uIgf+aVfzJibCvBr3/kwLbVruBLGb/gr8orc/D
6cLZWrdkkXjhcA1GXMzCVfwGb9XwSQw8ZM26GtcFna+MoMU/SEeD33EMq2Fujvk1
HMMUKMbOjpSEtZKJus0kNbL337pzqMYfoXSd9248VAUGj6lg6LM98/K2Gsuv4HiR
z3e0amaYg4GveM7M4kebosLOIBp/IP8HRjf+EQBKvf2esjMdRWAg67VKzcUWXNI2
xJIgqCfAVvoB3ebEgL5JMToP2EtKuLpCInBRJLYrwm1pek2EfAj9inqErI4tO5/V
Gxw6BISnVve1RUxksCuvnBVnutjDd/J9k2+b2x1MlpB026CzsBnwc/gn3Mg1qrq6
GtCZsLmCJAzgt7F3+LE7aw==
`protect END_PROTECTED
