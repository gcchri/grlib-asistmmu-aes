`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p0Gw8vgMyiyBX1bfgnMjguxFxCanEsFtN9GO2I1Y+cOc5tZksWC0yesrjRJ7FblF
H9D7hmGsGkIPUsLK2dTG66Vet7cXQG0c2ewzSajW8sApqznbLjDDgU15/Egdmyu2
5fvlloL2Pi9W7D6i6B7SqwfKOTTF9P9A6t2/V+bFuS0AWF4JaW2PBO+vOOuplqGF
o8zuim2N5drBgWysMcQPL/Ot0U5pA3ESAQl31ubC8pM+8xyrDD0T0PaIMNH+0iLw
AdeFg+k5PpVbpd4I3UtqF9FfXFYMQaCkEJO2/dZbPT8wqyz+nV26ttwMTuVIYkH9
PPSReZKakH/NAi5e0qaVwVIB85Wz4HH61vVHKQEoryhQvwRdv97QYutVhifFP3ww
V75EaLVFKPYzU0A6TTwa0s7LWDQR9spKFAiMZzGNoZWsZKwR+pClH76TgA92IAjS
uYV19PcuBi6Cau4257FRCg+vN/0Fv9tx3FASyOneZtMvf/4mYiqC/3v3iDjGMblD
`protect END_PROTECTED
