`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uz7xOyGO/T6bFo1ure1tSIHXRDFg1HsVne8FGRMS10YGQKPOG2SAntIwNhZmLNTF
k8C5lIEDJZnAwRKGto+CzgFHf24k56dH0jBOmBWZL6AABYf/gSaavzkcI/IzzXvA
mKJQbuR012PSX5wDCohE193R0+S7Y3XnPKoFOBWo1j6wha9cJRVVWLE9Cpc3zfgx
sYS88wbPsCW1REdAZEj58PJJfsu2Ny0OcwPZkNkO9aVvJloXvjUNBEJNWslJnXgB
qZDGDSCnmNf+LkdxyhyLa0h3VPaPAh8VomiOVBjVEu1t0v2mv0VLF5vC0AzWzf47
GEeWYdtLdH/kzef2T1r6XGWyELjznlnCCcE8+C7//P/fMWCgFZr2SOm1jXjJpPFV
YZE7hnAW7XB1DrmIvh7MaGPgyaVKPvWoOgCduTLbpW+qaSP1cyeQ9lTC9ldf2eir
ZmfEkwcoilomNFBQM+1TCBKXNOVHiVr4PeR1oQzpyQgAOwAOt2ZnQHOV6Eme07x2
mDhNnKteRl+LljmNLLun5ftys2zKWIMm94AsTp2a6ZoLfHcSyZFhPTGimOSJenM+
xP3xdrQ8tAkQia5ZKbwh6tWFilffJwR0Etn6pi2lYYSyNFvW5R4SBJyV7demVurM
4MSaVz9dA6AoV+R+5gZoDovB6RRJP7bXlfLiK5i+Msocjs21cIWRAb/9FouiY6lL
y5zZnR+s7lTUsBRheY2r6wWX0pUSraLHSwQCK0SlNFuqonC+kWUP7Y3zNjKj4xYc
6kA+NIhLeDlGCEAzVYRmK6n6vulkeO0hw3DYe43cU423HYdGRiilSVH4w9KykXpz
3wouUqzCaGEJVYbHWGu95uDY6vOJMG3T5bMJB85aeTQy7SuMJlfdrC0ly9Kk/DX9
OXnjC16cXnaitQw0Gqr/u6X1nb5zPUxdMRQLqYlgIo5yW2Js1dFlnTr1lha3NCC+
`protect END_PROTECTED
