`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xk5V2xEQR1M0/lpAa6TMCbEMFDhwB1htK9CCFNu1vmyac08EYfMfZfoE3eCoouc4
ARK9pJXgtdiq/kYsMgyWoqe6Wntji4Y2x8pnCHp/NPMeIo3kNLnWISRgRuJ8LSvP
vC4gw2A9z3nh0nWGn5T5OLhZnBEgqLbmZeogRLcYPU8zz7YDJMoQzcKWhudj48By
0wlBQBFwWf8ICao2Bgc4EYz7b6K3EGLW4p9Lwy2uMPSl7LcE/F05xPOLxEaygZVs
zzuL8w3qH46Oklwn1sX48MfFSLXV32ZPjU1zMD53pUY=
`protect END_PROTECTED
