`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
znsp+p37mvrKVLWDJ7cR5g4UaYzFJhuwHYZB2eA2paOlO9Lc/HUSYDQFhR4Y/bvB
OETnhgLxfRvYlA5UwZiPiF7hZhjd+PfI30wwKos3gqTi7Z90VBDXEcjKsy/QujFx
mnDhlyhlrsVCaPq32ZLK58gb/NBjqlMeJCToQnuKh7ahVJthUrLoUn5rfuNhWyb8
mSy8cUAGt8TyiKcwVxsEiXsLUaUau11KwTuJ1OzFPogs4cCugY3nEi4bAGG+S2Ba
1AR4jKqdr4Ol8Sfe25VGUpylzr6UF+S6xUVNvMfcz+kN+GxDGEhn785MNyvR2Dul
hPGhXRQ30a776y4Jygll9AuwzuJC+GJ5Pdejs80rbHIC60zcNXS+h7TGuGQATB1E
0sRw0IJpqWtm1xp7/JsSfRXbi5yFeJkoak3s2I7ixU4d6ffyLxAMM4eHkGsTR3C0
CAlzN1EGmFgB2l4Y4/bnqhLVnVCsGsDpTK56P41AjyDRlZj2z61Sr1bun8dICQWj
mpWLtM8KjiEkFGYzLIVcYI6LySwB91vaqKN3phpXqjd+CkLkNEjcRssclPZkK/nd
yWBDgBgPnmVkC8q5lulwnck8xFfXf7SG1//OK/9nulj8GVGNJxH90gZPhq+gZ41x
1cDvgXtiahn/jD8aIyxu4k14OYk7sfKeVhHqgboe56HGIsVE3Ha9wmEe1vM4SD9k
lrfYbf3Jf+H8AsNVoR0njkmbhoandxm1HO1vOQUXDaBfHYS2JkZ3nla3AW3ikpiB
y3sD9ErXjX/9AmBzxy/dQm6FwGLt+Uj7GonSkjKPLeVogtnFuHUUYeQ6EdUC1XwG
Rhip0HnUGygsPHeWNa1H+kHgLbhV3pnrrgWr6wutcB21zbMytziXT1/fF6Tq2wU4
EttS60aMjQRtcUsL9F58Wr1DSvfxgh2s9C9zMpaBWp9rZB8YTTYH01frqaE5PUO6
KtzCAy8gKf+x8Z/KrDFaCz9zPUMh4F2ssceLwHsvYyeDkJaFxzCxQyJmaONda7ln
6+Q9s3zUqKqkgZOgR7RsBaQQEyx0uhklcrMS1oMe/xVrSh//j0s2XJ8A9/ScSp3r
Ui8V2bPeQrLfFFehE+V6rRRz33l60VOF6bVL9GdhsqbDaxtCgP922DZJ3Y6k3RY+
oleQ53BjZ0hEzCt9ugtwmVMFO8mgtUFS4uqAJwUoP7qVczjkBdySSX/m2j/hP1DJ
79TJ3+Qo6tU9aq2WmJ136DNRVxYKWIm1S8uAl0MQMxY9l7/jDT8JojSVYaEwB0pl
OANSXTFlMGcyDHccHh9ORMfjTJCJdEvE66TCnpuZMyI+IqsHsmj8NsF1iyfkV6OG
xayrW6q4df/0q15om0VLGouHiboXo85Mk3yc2q7DiGB/lQ+Db78fR2ikjIdDb8+1
vQpEAcq3HooAzed5+YIX9MPxOLFsEZwvLjIGKino2OEyoAWr3fzEJqqGxRsc5ddS
8hEtl2+jW0zc1wcxvkJvaZvZVyipFtw89FIbJ79rWu3gOF9XignUU7wGNNEh88fF
31Ug3q37ojaqRr1v+btr4RRewQxZxGzP7/TPjfe2fnkpJgINSd17PFTVhxY3VoyI
l3/oEMlrYfTSmp106HifGm4vPHfcFaqROTwdw+gf7Ilv9T1SLUNl3SokiBdhyKU/
3ozo9Lfh/sa0NX/gzmKWLIbzqDgaGo1X0EZ7tFXTx861YKGAEz/9RV7n5uqgSQll
BSB4xqcOUoMCt7jBK2F/Qe0G2NlnJzeA9eMRNMQoApYcmxJ59cTrASAAIPS5MpxL
32rbOpz8zAZ6/6fpvvr2G+B3J9Pj98Qux2ACvPLCL3gzki/gyo6kiSa5JLF9WB/2
wTbauHhLAFZNwkAsneNG5InHsfOKEG1/L44bEdVyXTyeAD5DvNoFOfhdFOJ4O4Bs
hTr6/Ord/m5wLAqJkSu6EytxSHThp6rPJhWT5p65geEnf/fivF3lMX5U6E21cy2V
RrKV4DsIw/wJmpCPD2foLrdsAtG87ZDcztVUku10J81UJup+QDVZhmDmXQq3SraY
cZi+26E9qu5HbD0WMKGfE4PolxH3RqWSPmGm29uoQujqa3XkOVPWtfGrTZL6pRFl
+L20hlKUXdd9DElNxh7RkwJsSqkDeAXzLflfb+zbsgLv1aiSK2GUWlzR9kIV1dRh
7SSrAcPPsgh3flR3LZzQnHQNdGsDLSgQgYmzJtT4JrkArvghlK7m3c+p0Nh7TmTf
P3PVKbK1PxTlFl0Gvajl56OHQcCVjsx2LKPC7U5WD0JbhI3CRBhopS0qUg3X9Htz
swhea8fEoomUIIxvBIwV20QJo1jqcz4qORzS7h4If4M8905LmQob4RHsyuBgUx5r
6pB1jhFrynyuU4BXwmT2y/G4WzFSAMovl/9GREbfT+8/Y6HzeCKcrgJ56xSqi9dH
3327/unrhXKTRApugqpOSKWX6hgK9QYrHawLNppUvN5cYGqGcsVlmL69HNANryeD
BryaGwu2HlXh4HzhYpOQHobKYR4Cestd8iUoTAirefbnsTSSFAesnxnGx+Cznjti
r1VYVUQQcMfntm9mogOpRw94rDx1IrgKakLDB46Wnj9cW3qGmtAlJfkvLYSls0Z3
w9TDllUbeyCsdyqRFOusMh0sdJOEPEZKAFiNaA7EinV0jIWwVQtP026o8rGxSTog
W7gRJfSfPwkrgntDhmkwAsNZIEmLi3I8ivJD+UrqhfxcVphwXsoG454TXp7c4lQC
`protect END_PROTECTED
