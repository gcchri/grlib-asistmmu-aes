`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ns7HNeZJOEG9aLrDkszJCzeorAqKIUngxcWWA4nZlK9TFysh8pljoyIPHAJ3G7Km
0EfpzPFzKftZ9PkxyKFCyshBjLDk1lG6jHPABMB6qvLpqCPE+l1QX0M7/1tfYnkm
luOaRrgT2wfSNdvKBlwyynS3yFV/xq2H2EBPnRNTGWBLuE21WTzWO4YWC56Ou1R5
18IIELxeueKzWzzGRxJGc/ZSFa+lwUE8eWJUqYp5fz5rl0TCtLYg3nJlknCNR/Jh
ci+0r1jtDHhJOPXi8Lg/h2p7kWv/0dSHIgzFD20ew60TXnoFyf0o2YABcFoDEffs
vjhBqMR4P5IJhSGeVJxXiGiEu4L3FxD4PyaQb9tEx1+jqEIYfDOulBeXbuh9YQuv
9+9ppGry3PZump4jz0JnI873h7fdj8BG1R9vJgZk6DxpogbQv5vcPZtdso4vgOPk
ijc21VK90vX1AVzPEsHGKBzJfDNxTcupBK7hbk+T+BusYb+ZLpugPu2ZUG6U77PM
6rJPVy4LRlXY3Db0kcbZsZWMupmvN0k+hU10w6eeU2BZHAB8UbbGzqeWjv/p91Rb
4khrnlkGxWAwyJXuhoJuZ459gNeg3G3CoF9/KedgxlJOmMPYhdI7FKXnpO6us87A
h92s70Ygc98cs079x2AjE64NOdocsHarx6VdyxB4lwZ0QNtAebxZFN8RqVL8fxEK
H/xXKK6AYpvDhoqxKLnZrm6WDvhLJN6N1mNA6YGi+ECE17Oo7wAu9jO2XEDVA4oZ
BXYeEVYxakNFKNhtItT9exx8OSqUPnF0M5HPqRX7rY1Mxsr5QqmTg80tfepOtrCZ
1uTYg1oxrxz1VXewhgyIOTu6Gd6EPk5ihalqdrkwII+AsvoOkjb8+5iWxs3UZ9bM
OIi1Fef6o4jtgiYWYp2oxlX5rtpSdUB7nF0fcN5RdA7gSrTGIRi5QoWPOr6aHnw5
NYFcGwpGCn3bTczWsWcFOAZDtLDoogMQIw1li2csfwI2hrWPnHUFYuR7HgUGU1wG
vMgh8OgkIoze+7Zu8uGDghLeGH3z4UZPmCmGZKxR7xeVEtVmzyV3zDzE/jjUNgak
Ibr0g5i1Ov6icfaxdQbai5VrjatBlMU1vDUaKuHqIfSOgrfxV+wSY1jhJCizvx6t
b/CnzxWg9NGi1ne7TbhiKh6VSU7G8TcAEJ9ZFjpX3G/BSwXEn7ntdoesMbiVvMu2
+HGhsIYQ3knkFnXJ8jJ0y14DLugc5U0GS6TTF5kSkG2hBAaUj55Ox/lPY53KTE/H
4P8l/jxuqLA7VbHdnZsGwrou54UKPplRulwQnO+gtjPDIhMNSOxATEH9hi3S0V4i
7hJSo7jarUg9YeZHnybFq6ew+o3DX1xKDlya/95J1ql04HQObs7KJbGTjgMDAfj2
giQyrg//J03wlcXEoUstBKmAtup8qVw4ZWvOh0/M1SOuWrfcElEuofTk8kGPjrXW
VulSCZIbctviqFkGkyzkenM0dh+E4vUassAP6tU1tyJ+an1O/7+cnjGTsAE6fYP6
EzTYS4AaTug/+29Ai8WAXRdoebgu7QnGXxf3B8qto6zo8le29BaD+eUnsVbxvZzQ
an33V9+oPsoE155H2clXuH/RVTH+StU1/hkMeiC94DYf47jKP3YtmPLetLJOsB57
qiJqQn9L7d66vlfaHcxyWA9AKQBmFBNb4dyLmGjJrLn7tEP0l6cuivcFcuD5tlWI
1Yy4IbmfGif4OjLteQDU+ngWb9tnvnH72PUR7yi+li4Z01x3rYDoi+3vuGkoy7PA
nzTc/ThkpHW366/Yk6JoGVjxj84FTZwGKYITFlNByAPmkbBwbcaVKR2DGVEvaYHY
xuuxsJuEtzAq6vSEtQRYgi0MCUkSjWLfR+/pxLWexJmoHMOvksGE+26jPNMTzjB4
KCDRaD3U4qgIILyt/Cgn0Jjj0hIDdtcgKfIRVX2Zokq6j8snd7pk6G28e3h7OBJP
qJPSeRfuupHbshEao1XOrd+Pe2bOjM8Lbt0LaPzfgee83w6Qu/yNNslUbkzZ4aFp
fwhR6313EEEP99LiTHB/b6K3embDIbPf96gH6SqlXt2Kh5yt8Trt+nem7QwiL18R
ty4SVyNgQoQdkS7UOAtdlFgBjPy8VgjYoFh7pvAO1mvCf5Pm7nuusotsk81oR4qP
+C1Hwe137tyU1yEqMdALlTHonCKxENq9wV5Qg83D8XwbL+O6oU6ev+5acKozHyS1
P8CydTVpf1976Wu4nyMbhatl98Y686KFHJG2oXnfulFW1G3B1NMoO3iWktYeS1j8
zy8vgMjUuPovnJYNAU+JckjBSABOuJzqlhSzFsM4wzDemE3hQhw9fGGWKxmcc683
05zZK4jGD0K+D7btPjkw9ut9FLNnpxBupvxizNsEQDBPhh7r6FAsD2isw4DretrK
AoXpzGqxx5+Tgie6mtJM1iW9u24zdIKZhUAnYYJfQ5BwEzeNf11x3cZizHh/EPWc
/X3G+3lk0PAL0MxUzUIpmaWUbyTKUYL0dNe6f+gre8urq7YGzr7SGJIzo90nK+st
Sc9Kk3wGY5n1UL86sKTs5wDJaMhpmNA7tVNMmoFkE6uaKGE1pLhDD8/xwvWugSMs
iXqKj+22ebBX8FLGSUjQfaabbNQDQG1PSPT35U6eQ/EcdyjbwNHslha5w6kEB0LX
vxIkRgB9JKo30YZPBxl66KI+rRH2b+aUfgpv9tmYwLxPheTOa//UkCQg0LV8yigF
DI3poRQlX4FttkvkbDk6bOlNiSQl2cVDPeptY2jODDyzbQykP1LnBVZnnCGEA2hq
EzPOnCtEEL4bYmmMpZwD5u/E4u5k+jLSeHg82MLPDswvg1MwHbmEPa/Pox+Z3u4I
aTomXEgWQaHTsAviplAlIOWl/CMmdYCpqEor28m0PlfQlmjuJYM4uru9JCBPkBr/
ReupeREa5uI8RpsG5k/BXDEqbqx/7350fCx4OHIzC5V/8tq4ZExNi81B9tvRjviQ
FCwNr1coVu3pMUbX6aTTJ+H6tQU/Qu8aVK7zDUS5VCHE1jnFYxShif0nyn80wtgN
7GjPWqenG2q1VkreY7SBoHdCAkjuwyFu0CfWCqKHE04x81DrxV+kV2zzS1iZRs//
SknawZQNWLsVBJvqVTMA9VbTemajCn+Px59yYEHXlJb3gApmuWB+Kxt/4+nJBNfj
gB0pG1V1Akz42Nh56eTSWhksNm/SJjEyjYkZaJjvfDD88tRrs54wVd1fhd/fFuWX
l8nU429y515aUbc8+yOIuNH1w9VF6i135ayGNPqke/7NgUa23wsw4yzgjjNmPWvN
sQ0lEdvuhf/IP08SPN6BKDDzeS51E58nd4lSjmMo1sUNNMO0UBhtqm3J/q6MGfTX
tixZc+F6GEyu9ovF8A5QKmTBc8CUvRIu6Qs3Jdb8JIp0wVY/M4WSwJIvkD8QkyPg
I/Oha1SJDp73g7G8yvea8id5fuIj3oD0TmeG0ABPkv+0jtsJZCGTtgVQLx7pmPL4
iunYbK9tvnQ5nF08M+f/jw0RkMtBToB5V9FbLheERa/u9QBhpB9iuWvO/KTtRb+m
x6mCqKAulVX/41H0d/qe4r/pV8txdouMVdCq3U9FKlufFDCw2+uvXuBbVGSHv+ez
/F6PYM5pZQe+28ozo3E+ekT03wdS5cPO7cJ6osywZB+iLaUXYGdxhHRvTSUGdym+
E6mbyDsZhpiS/311F8hYbn9A7LEdK6lLFhLYfE+yjMisvZIatWpZ9PmWKY0HTdpr
g+P7mPEtKWh4p0MEFJ0HSCnuv6+AIpXVI2FReTLtJZdBGpc5Z2tpV/RNn8DOluS1
oNp/h/NyI/V+GLoWVrwQL1Q2c9eauVUUlxIY4y4WGf6mDq2i+R27qwVozox+nrNi
OqbiszbT1MMwO3QwEGgigAXiZ6c3bb78FzXX7E7KqgtG64xEBkI9yhHlm2s1yC+o
0NJgberaC3nHvRy4z1k1TGPHDSv8LYCt4CnnrDGmWww0jHseFSZgMYRR8eHVlppl
VgMrs/wSSwoVd5Pty/mS+dn9YGVyACrGNHosH+bgZCOeKQq8A3XLpmA/CqAdFkRk
zpLgVjzpgZi+ss1WpwJ7B43w8HFYalxhxC2YrZobicqa/LqtWQCsxHEW+W4nkYnm
nKnlvu7wixzKeaCKnPX5a/gzPpMo2P1jeM69ImgtxZYEWZLvd91FVaB6IAmqcuwp
/9lYzw+j6Whzd/bzjq86BHY4OkG2JSwb87lqpT21qRdJW/g3hz+DlpNgXxLjUcvF
Iu++FRNGkAPchByT4A3Da+h3gvwb+2Nm/DhKUzUypWUuvbmmCY5tqb5zdIbbtyoI
ZIju6cu8s6iLRPYrB1zcIg==
`protect END_PROTECTED
