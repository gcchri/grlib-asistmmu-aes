`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LiyuDqAINfZfNeQKveLfx58GVJ3Y7F6HPkKAKPfQp7lvyc3AJ4SoSZ+m0e9a2dT1
mp+Qe+d7aemEqSCxn8pG6TIujoZeFG9Gs47qNpvd8IYrgb7wenKC58v2RPRfabzv
xOvDiEfuJFppRL3mE2/z0aTSn7zl2B4J9mit7OuqzJuC9WREf5/OMzJlwbiZ+1ff
08BiRqJpOKFaYQ3LVs2ELE4sXVKEunq8pw+OkUkfGZoFNOn8l2F89fR6kgCs30gT
9UhHvY10vcuGbxEtvssVRFAkYEeGCPyG1P31DCIBJz/MrUH3IHnsN2WMPrRIromo
OueQ4RlTjN2nAvG7kRRrYYgCV1ZBeXAbCmwxH1JO7bQunGnRxINN4RzmL0lQ3kxE
U/HXzGbcNK1YVQWpVER5raM7WCTT4H37lsM7KT5uGMOy7IV+gaDtUxk+wj+gLd1e
UruvHSPPmM6HyBSxEL5SPe77cY2RSwFdd5CqK30q1WiWeJ0mQDh2hmrpYV6Rm024
xQh2Uv2DjWIRLWd4ZTlyotWA9Ei23OguMoA6Vk0UJweZv0wT6KQC9np/eUgz8YgZ
49/l+dj7DZP9nb1fJd1O0JOMH8cglaPSVHrqQ2l72Hs2weoiGezVp2V/lIK/I8Cf
Z213I44E6krnQOM4j02kXw==
`protect END_PROTECTED
