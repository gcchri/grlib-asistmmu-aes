`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J82+mfCe+OcgqstzKqjfw4dEfBN5Ph52vSOr1iQWS4r4TM7srufNmbxC4YxWKFH4
NVFTG08ezXV2RRLHR7KZlcRNwXfAE55/UNBMvpCqrZH+Q69Z6WF5aFoSxo4bc5ye
tMrDyGLXHdJCFvZwk5CpbB4raps+hkTSpoFz/BSk4cCgqQLyksCczNrBtqHBHGaI
bc2vR1D0L64i1AD0Ck0+g99MS5khSVzUS3E9963NhF08LIWjofl6srnHloAPopHr
t6ol734Lz1DUOXijQCRiHKbiLukh+fAuBSpnFngzWje1yJkeApZ8YA5vQcxEnj4s
OR4YpIDcXOvEpRAtLtT/vp+9iEO1l87vWmCA0BHPRkTQmVcW/u7cwl64KV5zJsMa
UzX4IyakHmYI2seX/KxXgDSnMDhjgHho268b2FjpU4cVuWb7qC/7vF6zUlGIEkWT
+B29dXGwS1K/yHcnYpUTMC3ebI7+LQ2mGb0BARZXdQrsxRUPeM4bK+47tT6BnuBo
CGRmO+tJHgWL6Q0sGIVbhx2C3jvK5ioeIK14JOQ4q/XG7HKzxBuC7pJEBPNIn28H
QgtsGHsarRMS9/MsUmQzNWx+FVdMAk5zMUE7OKxoywZS8xldaWxAKkAzDqdRZmeO
5SWOBNkPMwk2aD8iJQZRKR7TwjTwse5AtSfzlqVMwTzGlElOg4KkVF3gyhL2nFwg
PUJbb7wUMAVfc5Y3eEdIqTQpa5NMcu3HdMKtPH4YT+jZ4HMdWbE402Z5Yjl8sFSF
HEajCGzt4WCuUpVgofI3VKs3J7N15QV/EewkY7aPzQMJV4i3DNJqTGF/WJTZzj3R
28v9dHtChhUUzpIqrEsqNhTyyg6R8HWjGXBzifAcARo8SBP3nskSr8meD6dok6cf
bunw7+1AD2TtyNWvfuTbeK/jLtGTPzSGgwBfx2RMezHGLz3/CkGogQQS100K+u6S
t8TbbBcAKsxwKDOqxNs8UUBtl5okuuqFxVTralOYUyEO7jvMEG56xYbgieYXXn/z
M5lb4qNbGMs7SndhvecGT5kWY44d+QO3hfIaahxi6pJPSXpTIffLBT5TXEn3ja/L
sYVzzUwbRd+7K7VFHfrcQdBMtZvkywndPoxnnZvBmZgPkP5lrme8yuJV9vCrtGS+
Uyn2sbcjlWRv2GR8Jv48XuEZvl2kGB78J/KuKN2Lr5nUFehylz9+7Y//5PPbI7pe
TJQ+mXOTqHxM9cJjWzbbArA2n17WITHw8WZHw0Vb+LXEAZeoNtk4YPcCDPaiq3Ut
CXb7H6XzGl/fxmq6N3LQKImp+VxCrCz0MUm/F83viwPTOzQdLww6OT4F88ss/5uJ
0oi3YX9ttFX/0KBGB68wCgyXkfAEQHooseGQ2Gh8/TkYfed/WokCnmo/XPVCWN4d
EhoMZJ7F1vlyjl4ARyHTrABGgidbg7mxf69Mkclx9MRKDbSqwovi+IkAdE8HrnUZ
C8iFTNvUC6MGeEQUb0czQ+By+XUVKoWqPoaeU3e+x22tIUfDlHXrAPEWn+p+JBl6
RQo8Tfv6QyTJLbNS6JXbuEk9uIwXrkAC8e3Mqp2rIQTT35jYi28TgyIWeen7upFJ
SlT++yRba6PTdOViwDzMXPJAqluhXbd/KbmQ8G7daTwigDBRvyO54Gi9HDg2Rv6H
LFGUcHTPESXo/5OpdCcw9niezSc+Tvgth3/bUVEnNOWVKxxL57/SWl8zb0+67N/y
BRW7KUDfC6krUTZvRJ5x/OhSOLotUXOHa2bvXYhJWvDYeEfnWfK1FCU2KIkMsQZN
UlK0VvPT44bY507kOZaiDyr5zq+9xewJcZfD/5X1TXU7W4w9ZMThzUq+ogN5rmAf
duhcHTSG0jZTxlmW5BN2CiPytt1Z99ki/9HUQ7GvHLvKqZ7tpfWKHGD2eb9DJy9z
c9BXAmdhU0bMqIK4Dsf8vl0AwKZYt85hAD6RolYhUbQrOFcswEnEZ7jAvRRx1nCx
PKt7FpBnCYJenXvXvBBpWwUhql5EIHVYwUA5cx9t4eiicAs+Wbq8UsPZVCG+Hv1X
M5KLuF5WWx0pbbSgKdNSIFgQM2abhFKkiAfwoYiKURUBu8Qpl+/s3KNUpeUIlbse
MLEQc45VzdFSoJdpc3CYNHUej/IVWMEh+3xwMl7zDg6Qb0WDBR7rDubhI5+iAN0A
vC3eU5WHzkBGEaLtVb48u6kkmTuK/bBgiuqYesvj9V49yZamRJEAlS6bIarhEhQF
tPfJYzsQkqtnytF7UJcdQuX73TVizR0nLRSUVBgpT2ceBZ7N6sbOugYDOaeAesJd
3EGhv9c8156z5i00tHvz1X1akw0cAHj9dXEAcjRt6a8oPrLWPDpfCmjOGGmApb1Y
LHEDHi6DGViX/QjfB6r4Yw7KfK6vGhLq8+X4L2jegts3eo3zfoRjCawoUSZkFPVq
4u36euSFXbz37yI77nkDZ+tYY4fp92+o0jB3cYR/yncZlRTuSexdMr1zeq3X59Z8
`protect END_PROTECTED
