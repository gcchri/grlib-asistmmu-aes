`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zO++IQhXPa4i39SE6bDY43bRcuSDXW0RPyWS5XFtVwp3fHhV47gWcdIck8QmmU1z
1u5GdgY59Ugbx88HfnqKFX7MAL4WTyBASCgi0cEh7H/mBLckY5j0CPueLrHIeiEG
SLlVay/dsCvR0uZ0+iTUVJsOMgJGaKOM5swXVBoFfgZJxKaEFQt8EY7YX7ss9Qu3
pq6ArHPvJwO+iFUef4YPdCH3PKcjcK+kOF3WI5MSRE/wdYwUdeEwu0jidH+Y9dsl
sMghkYCz+Dlt0S1bQWBz0DavNw5srEhmcapOto4pXrZ0jJ90Sa/zPaD40/o7GoyI
OMIS4uhfTdIb2uY/U0/yfRwN/5hV9drlvEKf3d8F9z77Lqs14B6PYPPk68zgt4IL
9/Zl876S12cnmFKdnSb7n22S/NeGHTIwK4H1kBD43wc5pVWZUigfuiwjWwKzykm3
Ke5YxVmHfLJkUel2M67R0hpLZBDBZVcuXQllMTRw1hq2nfSRLVA7TcbWB7yP8jDL
v8VjZEW4LqK0wBSmol3drbYJqNfreT071hyuUHMJBGK/V5VizhJS5XfbpcAwv9/d
+EHrxes+wolbTRgNd4rEiyEXzyys8dfiFFCuX4nmLFoAtybA6UEyLzP5m1sh4x9z
LgAyJ0Ok0/64VxYhey1EHngRyxpn3naLn8wD9cWSTDStLDhDkc/nsx5RJnQ9+4R1
RNG/lVP1JbTB8NfgNV/zsuvi47Hx7wEwHo2YBrhNGMqajcKNukx5W+FQZ0H6UNJl
LuTbzbGMuIlDWpCHEC/PKwTCVKtgoQEAhpoHWijonbaK88fYh5z/EdMxZDBk/68x
0fmWmI68J+RFUy0suRSCCBAIgAjxKg74N99gTQhB9yYsfCfpAXkKCg2ddZpnSQpL
e552Sw1Kt8Ve1yT8SuLwSsDdnxH5i6c3WzsyTzF1S97IYlIY0JZaqQucJRTTocWh
TMCD4suYS83Bf/28LXp6d9QOSOvWxhAyHPnQir8a/CVT7LB6ZOxI/2pHmyELY0Zd
P1bm6p6+oXn2ShPEp3KIzDBc6Ay/9RcwZe4adECmeFfywFJGvgfdlKkvPC22uVZk
pwYQQU7bFdQzBkQK+QAk58tq6n9nCpu8F5n0H3s/DZMFaqIL97nmuvBo2fIlcT/P
0y3o0lCPcQTneg8i9D5sY3wvcPqwzrFp83iS/23oa6WyGmJGZuBeStGOBrX/F6Uw
z54xN6md9OEDgtkW9uuhynOSDSQkU7uzfNB5m22q234R4WyYorQgovB8m+e3+QoA
NotxN0ByL7IOZeojGZQ1kA==
`protect END_PROTECTED
