`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hzmjRYzoS3JoUJ7B3R+JESczkdedBdRg8aQ9JEhHi6cpE4rEfYIf97ZsfE+KN2z1
gwqM6askRuKi1/lbk1JeiuOpMRtDCMrw732+2QPwvRZJq573KP5VFTQT+tBUQt6J
UWiZLpAeYnBuCCwmbMmMuSfA4w2Vt9ZHVQLhiB+CN4gEQ9nfdMB6x66xE41wYEtZ
j2NF2dhG1imIUxUt3NzfGemZ23FiBiAtIU9yrKq/Z98SHG8HOeyE/lldnakLENmF
41STlNEhwxS6WwPXUUVvPEm6xA7unRSgU9Fc+cnTCIc5o2L3Z/Dv5SFQvFUfeOnF
f4XdaG1Ygh6sF89Nsym4kRON678FEN9bXZBt3111baQS4/OupANhuVuDatdwaBzy
`protect END_PROTECTED
