`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIiQ8Eno2+lMztOnsAr8EBJf0lNE9y0UMjB8n81nCKeGLT/Ry3Ztc6ExgQAupSFX
NvihG/+hQZRHi4MfY8fAPQTLIEs6XfeBy+P2cNurhlgkXMb4QhxVqblv5ls307Rd
i5SeHRfMXP5A/NDZgnKrNf9BBubstMY7xkAGZoXaYQi1EhwBS+AA4mSdh2MviVJy
JKJ5lC5h/TkUz2MAKvFvU3zoA5FlgYDXRlvtQD6ZrNldVqPqTv/DNb4nyNjizykF
dn4WMDDVSD/vjgc9urmJou1/U0GW2RgJY8muHz9jWr1KX1uHpNINuQSiyLrZW7A8
6EZ6BWK6LEAHdRJZUbsqWJ08T7cg2Wn3Q/4NxbO4GvDM/wZemlTcaQRV318mCopb
rRRUWiflGq3ZCHWbQQ+5wys+i5CSz+DySpYI+lkyiBmuVxVt9j+KgPe63jTf5Zr4
+OByguaA9uke7GfXRDXOM+2KmCOIJDK5b7SHguPrb4m0e1ja6GNnbZCqrLM+0I6z
Jzg188y9KGp6qEpxw2f/n2X8HV+5GHKsK8Ev52aifHSPpc5n0SrIVfuubg5CcO0z
FN+6XpCzmWz+RJwDWbrIM2MpSgJBOikZnjwSCgYT7SdQAWpubVrZjsmjQYcrFlt4
zlwAKTSqlgskyC/KO6niAWXRKlqQFPo1t/pacVUbLdE3vn/yEhKOCDMUsau0hwUa
xRg5LTlwZWLs8fpEQsqmMzfX5dXkcIkJSPbdNXz4jx7hsip+SAC68/fztAPWyvrJ
3X3dl6F6pfshEtUGHbeE0fyxYR81KoddmyGQ8O97ZSinBv45hYOzgC+xkYZitTXf
r3D1B3Ejxgu1IgqPKvDgO/a8MkcebIRTjMRe7750Y7KKc0+UkT6DUe59ma5PNvSm
KpKWqc4qz1cVGVH2dh/t//I1VOD8XiCwBS1smTNnnUawV57lJtfsJfXoQVVASdIB
lu4XrmJhbPM//U+2cBDKV8lnuSQOqEOpZj6MG893EEG3BfrDbCohyWqf/XjZj6bE
QoOdCOY4cPVifCe9Ve6A3aSnmwEObzGK7BjfZEj476FwZy0nxQlw7zLQVJYYNNqj
JzOVi4jXwR5UvzKpMQd4FroOWRE8QhbGPgMLRKscUFbotws+PQGmHBMF5jnDQam3
VtYgLaBySbhqo8BlKRYAx++8P4/YlNRTXnspIMwgJCoxKOQmIwvukY7AlHPrPPv6
5hpSvLLKL0ugYU7gxE+qXsCiEHu+UpR7Xh3otx0EUDrUylw1bpAOAW6P+bcVYL1C
oTwSWxsZw8LiKF/S1VOrdUbN8yHJQcXJvRryS1mZIRcqyJsYtDJVJkJ4dDAFvkZ0
Lb5BqUtVtFZwc5Kxs6ASi5QAbx8EQE4DAfZEmlU26Y0o1plI4xZksdH6KCxsDaW0
EDFZLi0B0DEjk4dSxIwLX7pXaRV4f+Tij8bBUoHE14gTXyMEOhkqyMsjuCcAkjUx
1P68On5/xdLyIxf4jeroQYlFt9dAyWI2ggQ8WDCyopCsK4OKgZ2qn/H3rYoR6B/1
11K8DD6TCGG+A01tv64DfrLxGclM0Kusd5jQQt4ubipr0d9wpcU8w1WawDmd2QCK
5v2vLlaU+2H/hvFvknEqGMBQW9KtJlzG6IMnOPUXa0SAWUr/7cCXeKZv0Fj1mAUz
+eyh0BRJBhS8lnXjKAouIS1KM2Bh5c+rE/8jkctb7kyZ+COaG1QO2RacWEC8P8rc
tuO1H1TX4afmGBQDv0RXgABHREJx2+IbQLrdCQKgp/uShC/NjZbo24K2R9n0F9fd
`protect END_PROTECTED
