`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YrnjdG80nvk+hiumwHrYRLeDhRoI5L92gY1f8kR8VhpXkNN5B4BruYgbI0isjJxw
Ak6Oy1hrk73poQGPOqkeQez7SJbcsXeOjYO8Gl/lhTqhLwzpuOY6UdokNhm27a2B
jqn9eb8wuFrJDgAq1r9mJJktwAEZ/s9cCBX0BtqNEyhOrvnWZzDj2eMZKwp02VbC
4I516bu5nAfe68cv/B+R0hQRa4aE5IAsZWh2DIQyAD+gDh2yrOEfL1lmcdnm1qsm
MnKqmVbnNjfnntWeoDuzfuhMLilgQGHNfADxVRuDCpO7LNIi4XLFNwGVYVTn//Kd
g/2n2mZneGrpNGvTAJf7AdDgr4NgoEmSSDt4wHJI+It6nZ8dEsFuDdEwYyM3x302
eEfmfRnjoRr7tuyHun68oYMjKvAzJWCWMybyrCE5iRax5NKmirUiuzZMueytqY4L
b+hvdnTQASa1mlipPnJU7ILCGO8FaGCFe9BMIZBoDJIjfi9FjlF5WYZEhoo/4/7m
qW9UqRuGr8vWg/w0ulDbWj8MmmRFyQeQfWWAzVoOn32ies8m7x+mR7i6uwa+0QYe
+g+JNqSRl6igEMrUbu4Aquszyn2+xFg8819L7F9T1Tiz7ic75HUT4kRHhUHYzm45
w6gkVK5C3rVg+X5SI7u+UI2cF2qsUmTSC1Kj1p9JCH4EmET0Sym76ryQa1hxguYD
J0SSLszJUi34u2biFp8v0yyqUtj8wB8OSvjzHe/DAW9ocpx3xFlVmZLiZJkE8zPH
IQIsXN6SeT1aJH3CRVg5W9sFIW8CnwvF7DSHWnjcCsZCLMJG2IIe99oYCT+/KASD
IZLmTaCqJWhSpwH48e+vx5kmgIc+77+PIyqEOe2nVgaWZYSOPb5LJpOvKXVBZm6E
6sQkef0VInGMFJQfP7cgf+k2Wj0hyzTpfvwKCUXIcAFOFYDj/m8F1tZFdgs2ZuKq
oMqL7kJItXRRb7Kf/gDzE0CAe0enx4d1FfvfSvEksp5ODTnSyXFUGnyNcishxEMe
PJbzMmuZ5wCtO207I2WXlRPfPx9CsUzbrUv6cdi8TwB2lzu2xCLaTQoff8cNwE2n
A4yRfmPO14jANBmtBY/g5mW709wLrxtBs0ykNjukOTOoxDvllJIAy/o7vgnjfuyd
W/QLWn8ZhptAuQ9urvz/v1XSz+tu6cvjR0/ft200yHbg0aZsVuTLJfP78RubGIJJ
rNHiotWMP2aL8lxWVMBLnurHGi+9WJmsAWQyvX0EujibCCAq2OO9lf20TECHrBhJ
R5d8vfvsRFnSU9Oqhx6j1WITYaaJi+9f24tqdSUU/6Nz6PGOm+Xt+K4Qkba6xBSo
YhLDd7AbPj+eBKtsqEdF3Omzg0rJyUQ455eWyEpZN/eZb/V/8rXfJEAXMPCEAdck
fuUw+3/zqn/ZuhR1JfjmWFSd4l+BQ5Xss5THdmNHaUlLTc9sPloArk5JsZMmKTsE
sDV+pijparRhyX0CKlUtZKjEFPEuFUmxHpjYubs9Dvwnt0OV3pwliJ5OXOiYQHKT
5Z8l38j3WfetrX//MMQHzxmE1lfHed9fnAzRBKreUdYulrTsvKIesOGE1xjxoJe9
AsLHfAcEm2dL2qcOgUosfKv7XmKnJ8bvdSdRFYBg3Xvdt3sji1kLDl2C+oym8HfO
XanBAi32mZYh1YxA1UQQPzZtwEuuJPTBUi9iOjiZuxeIx9vPer7TuPfCPX76WGVx
rCNiguZiPG+j61IUOIjBzZwzTgXad83e0zid8DyeddCpv17XB/SG3f+M5BBYqNCa
hvahIbJ4A5EOxyPUAC+3uL77/A5TRnGiL7nGs0f6w5HLz5WFHeKpPwl8OunSrxpj
wMc745cSDRLn2UiKSZtL3TVh+iEaHgNgLj4/SFZOxOPqqNviWZEr99cTGyQ3yO1n
5JWErrYxLQKrfqJioNcXrfqVuUuirtqI8HpFP0ixknmxE/sJYzaRyph47ceGqmyi
mM5etttIqhbX3yyHFV6o68HZ1HN0iiX6EY0T5ljLRT6HURZ06cjoM2Dc4MqPh9gN
d0dtERzB+hHqURnldGO7jU8aBjBvq+Nyfgfx/RiJuMKPTcYbMrCSQVtrBqOFg1Dj
qNcxIHSYdDgi6NonUDDwM/d8pVtN+jFQIN8EekGPAu0uT/duXsbA+ESRfxYUkGhD
eRKJ9nr8f2fV53rECk4z8VNxCYKY/Yj1qxIBNftdgCdPS6oWpS2FdlTw6HPP7ZHe
4+LgiSz9aQwP2E9cz5BVzdkkowxHOef0ClZu0QfPGm9Y7pemdDBYP2oko4y/jb2V
WpiMdfmAh2V6D+5Yf6cWZexrEM2Q3Zt3IkKgGjwtK335QgZPHilX6qzB2lh3u06R
OHeHDKXjun7hFXx5C+cQhFLlEw/S1KGCimQmqjzEkay349EBQFKpLOK6guzbxpFc
QBVkcpjW4y7iI4nABcpJ4NeO1rNStNeOQ3Wi4fuACh7taLwKKORguQZJVHIeJi97
2y1amK1iDpm5Edqo7VvnyGszMXbkPqhjSXbBFCWqrJwkDkPrKwq7urwaTn6uaNQh
bbHY+7aMrrow5kp+NLH/fHllbGVPZUDsD2svQwYCwUKh/Tyq8y7lT3PdJEFpyrwL
rzUB52xDa6YItWoU3kkcAaasm3i5NNvCQNzdVhSbDk6VnKQ/rCOvvRrb1k+qOBUg
MDxmt9f2aVd4xiijJdmdidq/81EnxcV+Kh8J3XOS+fMq19jMTophKnW3ELrby4Lj
sV6Gs4Vg390sBqmNAyj089hiP2NiKueNNSRBU1wlO3d0cfKKpBYchbBu1XAf/3DZ
OKsGy0CJlmhdKyhXJCnz+fBKkbH2e8Ldj0E/XsHmPJDFwR/VMeLMdV6vo5Y0Wwyl
cA6RABHWbFX57LgBIo5Fo8LU2Io1eYiBDYjAAvxKHqYZ5ohu5NRkjbpOd4vBmmMQ
nGHP0JV6GhKVZTiAtQWUqNoI0cjOrWDVvHqAewRugEP8hVJweK3IwxXlGdTES/NE
StnerjfLWwT44c4PyUlKY59yqafXrNRXbxnDmqRxHzYZQq0+jnK6Fqcf3eDdBSOZ
ZnmsTjHRC+uZgYBq1z1gqt3OwJzPlZBZoBcIV2Islwd5b7U8+vFMXUfX/BKSE92U
tf6/YHMMrBhw4k0k9nZEUP+TxfSffLs8U+UGM90ADjK0/cSUtRC8trgL6lsGj0+O
QEN7qlPyfMIMezh+CESzsRTfwsgLe9ZxnriwI6oEFn/1niaIMLdmaUxPfFDapcJw
GV//1jX6EF9hGAWciNNA8rnPK+NO7rW/+/R4l8abhOp43pUd+NgPympGJPj9c8mq
x8UNGT1CThKxFysobeI4N2mBgmkc6SOx5IbANC7uxfauVthTWsBzuyCL3xzwmeX4
VIzIF8xzPREwhe7tAS6epMR1i0cjlhr+FrZZf7TQKu2glJDRRWvk2QeyEMhh6IXa
/Tp0MbfWoB+2Sns3AUHlCwZR+Sf/AMsxaOOLczZNSIQhDnCkZmLVW+gozHRs2+A/
1qidNf/Rh7ON5JnB7cQbV9mqIEg1VONDEVc7XTBd+pQHi9YoH0wnCLIEoX8QiLtH
5ORJHeE9y85KRkkPRStq+wMqOe24Sma1LVv5Xk5TVCKSG5nSqL1UzivGRggERVqk
1hP6R2ALW4f6eX/Y5schtkTyJyDu0VPp8gZJRYmftRB5HgPFeLIERz0c8JR7xkux
5a1cQ9oOZh8rBzIBTZB1sO0TDsCLaqSZrXoJbNbAS2oR3rz0cAEX6yrjAc/5QumG
3udQoE9PYkYHETXzwpPQpTRcLICir+mTAFLWN0ZW0xY4T9ym2HOz1qIg6uil3REJ
+7cfusJV1o2FM6fyMh67yAJKZ6fyQcqLK/5VifBcZYgw2RbcKdHhWo7Fb3aVuNCn
eZv7jU4JjSgpCPrOi7a6sANEWgZLMCBrIPsZW1IokPh1PmtKLsnH08QSvkJfqeus
lSSRoRAJ4RmmXXC44GTng/et+lR3uQoEuefmcTXEXmbVyspbzTK6pZLeQURTT3iR
Fyzch9HH8fvOswKn80onBZ7sRM/x0rRhcSdmJnmmWafjrH2ksDyyo8zUCfwKaObm
DCq9gpJlCTF1obXg9YvY4Fac6gXmAhUenwSWxaM01UOBPdK8REVXS6eBSNv5YfF2
r7xDfl6v1RteMw1u1VPmm9dtpu2kMJEfYT7xQ0AHNDTSYfMV3fOJzWuaZff1se1+
io2KYlhXmi1T0DxkkffIIMVXIrnige9jkGg2XWuaBfz1zelxHv9eqeyEF3hBMpMf
Sf34pgeSd3o6w1HetNZrkh3jNSSbreDUPR08jcyVVuwVCUdQdjw6lfUqrXcMGMXB
ejSF9hLeSvn+cmTMrGDc9HXa1RuznVQ0S1RvFtDLaRDrnOMWqGwbn4HbQ/DTBk96
7wXRL9qnCFhwXx1awHe8063z488kZS+7hITsElT8LuIvYaUkaS6KLPgYQ34T5hrp
yKDJ+pxyoKYZs0/bqyvhUTX6vrkx+WFjVsPjnU23PZ1anKyVpHv2IqFbJTxIUj/C
BdPnR83XcgbwmeG5zQcYk3vIBEj7iykYuAVOq48+CdwAb/wJOLDKubSfBniyORJq
ZZrijDB+F0zT7A9sp2uH/A==
`protect END_PROTECTED
