`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ogSCuH/l0JhoRzLP17TsvTO7ZiRUNAI0cdxr7svMajS/YF75pfSt4LZSOCACdLB
ROkVVSO+7BTSJHqPd39gxN4wCAhVjnsThfn8Jr/VQ0gcRcFGxiMAiHk6uioLtULe
kQvIDloIW4e8dDaFiNCjdLTwtp3AviTpXhwDg3+cTov01h+kY20VoTVVlpnefWeo
kWsAhrbiUiveh0zEfv6LbmSXxBhpd+NvgeDm113W3aMJ+zZJioUB5rcVvQyeIeFy
z1zyHA0n+9qBURAumgofWRA/3t4pz7qsYlEHcjYEj0EQ0xOM/p5iLMBuIaBww6S2
BjgYosqblFX8IP9hCm8TK65iUTe/GGKbTYnB+ysWU1h6s+GswsuD3/7kW6iVf61m
dXVYkuv1tNmxN+R8jFQi72LVU9OPMLsMujERzjnoY4HQpiEuydTr76HluUGl6WBV
`protect END_PROTECTED
