`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j0HANlDKfbwruwpdsDkxsFSQCWVVRM/h6To6JBUQl32Q0Xryl2+wVVwteYypq9aB
umh0MKBVq9XtxYshn13lYfa/pUuv7skfSvC2PoNRd63QpB9J8ydszzxe9KOUAecr
Zb9lWNkVod1fI6IPXgkh2vxkLhVkVUJ9TQjnz7BIowjtDcvwp7myzDJdn/2z1fS/
es92Lt9exuf0825X/zAEUI2eF27TinQshnVYHD/X1uCKr5ubcMdeFw01N/yEOUc7
daKRui3HSmUgr2Ys9vAugVrTkupZJjgkWwXZ8g+YSL0=
`protect END_PROTECTED
