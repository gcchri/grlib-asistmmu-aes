`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A21R2B2TyAGhYuA9Wl/8XkbKc7RQ6/eztS0YwP2aoLi47AaqtQIVu6zDvecbbJoO
sjohHh0NjeZij4f5M8W06th5We04xtCAQ60nnvReyC6NKKDayHWmXKb924DFVI2N
V1s4tUaUaXXlht6K2pBhTdUdS8yvZX73z38X8Yi/enWT7xeDebJHYTjtamnj0nc0
kNDvTB08ZBjwfsE2QZ4yGe593FWUj7DTEj3369OohXSH2LZ2e+L9+w4rkevwCqyU
e3Qf7o4eaocYCyal/ImdpoqVJrh7Et5yiXJkHky92s8+Y6lim0eav8hrHZLHanDU
ukBZkUpnMn2Reosp5ZnJmQ==
`protect END_PROTECTED
