`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
capUr29byQlss+xr3M7jrmVfYQI9Hm6m6knvh/g9oUU5hys68j9ogQhnIBl1C3a1
vP2njMGK4lkdnLC2zdnHlYesAlZTFHiaASeHCMiiPCIqd6fmwpyJAhRHKxzZMbu3
5Tutg7sezT+rtQ6j0LN0hDSazOx1vqHjmDq78XluNurgqoDtVRbpUwb3oHKRJoSC
YSVQgAV8S6hk2EjA1hlDQlYMr4yl2wlPpL1JGGax1zfEzPfn9RZkebN7Fz7u0VYm
59iwotiG8iCCViSHHCr0XNUG2d3ZQTS+94+gtmwQhCd9/RIP9m6jNlrkPgTd8DjZ
aMjnYWUauXuR71Yd3+16lCAs+/N0NXBSwauN+Jn/8hjFWd+xzj0oq5swqDgYtG1u
g1pydqrgXjEpPvdt5LC4+yL/tDJcRHWemrdprXDs+U/MQuxJMCcOomhJz13TzKRQ
hRPcseJaOMOrhHtnGQp/ldv2TT3eu5njRT6OFDMcOtSMyrv/AqwDruyp3eoN7vdl
6dNEtgV4Q9kfyNnbDvp4FaJNuPhUwWc73OY3PM/mFaFbihkwGXwEiwxoi7rnY+vY
6PXK1Tp1HRXOH62c28aBvWs+liQgtTEMWwRob8CMI5lp7WT9mAP5VFhqEYFrsEhN
06nXipcIPUbM7vNALTG0w1xQutbYcVcxFQlWJVjABP+CzFO52mX3vm3OO6YPhHcB
M0XmJsOgsqeWE7CuC34ijAvs44aJx+g4cakS/bi0kOCxvUBw7McehcfGFgcDqyh/
PX9DSaMjuTOoPVWQKXJ8S8y+QGh0JqZUrjt+UfwYBc7EnFXbS9Z2cKUTytWJbbTg
rfgCSLTsZ0s42iD0yZXaiP25bOi8Q85d6YjKmfD49nZ2V959wyS8uDTbERUhh0T9
z3oAe6lO2NyjpMUT297D8V3V9+otpxqp0InBwIHV1i/LMKWIioyAAoYfxfoA+DUB
2gbHNCuUR2660MsaB1M67wW6wazdsm0CXzYUQRQDWRPmZrG3RqlYVqFWTatKBkre
2+qyoSjABYw5zckRrRbgWPzv7SkgnRf6V+sBwD4RD7/Bpf6Mibxmt/0cqQ+S4vo0
/1M+C9ZM2qpxBtFPio0/oLrb2Ce3AoNNPZCMBvnkauGfkL+7TRE0N6QN3BivCYz6
3oAXqzeRD/ZnzeieJKZd4kxnsmOqpRKKxpxu/7Q7oyTINnaqDRC9o5xGJbGJWH7z
vKebCgkYuoY5nVBTPwaf65i/+M0fspRtQQE5RoNmCV/GLE8XagxkAQwW9KX31Kbz
K5lE7BNsIXRe+X2cJn5Ru1vd7Bde0zUp1ZDWlmbq8hQ2IMgnZuPh6JzRJuQ2xSDi
MSpHTXLDn9Btjzr/g5SOV9nxjKe9zs78HFpkA17GOu3lEaO0YOLO8GP7is0Yg9Qu
9gJ1tuslRGmLR74zQ493xWZjqgi3x2n4Vk75LBqTiNCBdqWHZ6w80pi++gxrhhQ8
IRM3JGOoKlR3Im3rgWMEuIWehDvFo6wANkmNdbSr/xWAFqwhH1H4T/hTmObL+vf8
EaCRQ5SYUlsQXSuT3sJuICQoN9WomMn4V+AALYxzSjcTY5GIyu2V03QV0cxWrp8F
7eHTUqf1GVoSc84a/7nOsjBWr3iDUon84HEN4XlDM9Ho+R3gFf6ihAvx7SQ+AJtq
6wRnIfK77/rCXUKmdvfklAO3gfRpizM88ZsMo5UJDEJ0zEzaj6JMhQI3AVymi8o+
8GpGeqKtdhQSRCpbUfreJ5kRtPDAOUxGNIY/6Z0ZPMBo7Ys1oxOwzHRnR/m+Bom/
hxfen4QHHRaus56t1+R2cWXjc7TVr5g4xz0M6SDiCLMw7+zbpJP5B1I/elRNqn32
QQcbjaK0cVAoJ/SDCANeVGR1urz4m9L4q3+viOvgHOLNBOMBF5XuuE/6fNjTWwxy
yCD0epnWI3+7S1dctibrpqaqC9sXC8yTg9azAD5qIpybmxzhqJpK3I05Mz/Qb/yy
IHmz1J304RYaz51RoOsXHzIEcnvDw6SuGhMgTrcp1jsP3cFCCl7yLldzWbUiAEqc
XUnSZMrj6dSHrNZQjo5qf9Zvkn7/veyoaIaKrPTtRPza5LotjRJP02Nuo16eVos4
GFfyU38UQZMmo1ufV1CfbibA2b6GI6+uVYuB4ylp9m2zv1y9fTFPOAJTRzzQ7H07
/Yzm504lHjfSAj147JunbtwDXNySPmHB6yzqund13kzahqYgfHuQThVWFovOFF+J
s6BX99tZ/M+rYcfiHZW9lPghEa47a8SNZYZdKz98qdz+KpyqhBeZlyWraX02WnhT
ioJton1Nge8SpSReZQY0ORjsEW0HszdlisQ4PVSUCC/D/3tt09H01DXdZc1aMCaS
ZWcpMeAqI3RSPLzYGBJyv7AAMyM12k5BUo12FpTerRlBmQzVGBNWLRRIySL7AoEJ
2Tw8J/Y7geqLqD2aNJ2n67HpQQ5n5hM04BEO+spcOsMcUFcLF7l96P34g7c+xek8
M/kYElmknsb3XN68ihwcMlBvSuA8WpQoJ0z18pdbC2QivKfJBjHy4yv9riWqIz/N
VqFWHJXdwzFCB3tGpdfG7WAOV74cDefUqcSY14dNOy7r9l5WyusfnLhMW0OSq2o0
4drmKPPv9dCgf//63IoypcKpv0GqOz7T/UWHU/nCHIu12vFk7zTdBznenWn3YNVP
0c8q1QoZeM64U72ro8HQgajLFaWzotr/r6Xpz19UKifYanwxWCy6GehEMy0n/UXq
DY2SdwkGubG1nhpYfwjPHn5ZJ9mekwhxKc3JLJXaCJMiBJqXYd+OiR+4GcXucLWn
fUKCqO3OVYP9gZMeuaBTifpTs3ir+jtgknx4d/hCYSrHofEBvf5hqMfhp9oBjK3k
x/cGnDZhUcF2LfGHhWqXrNFQlMgFAIvEUNVt20szYnw+E91o9o4xo3PWbdRkzZAC
Uiz5YhF6MPoF0MmaG39CiMJQAD+DbXW/ojDDAFPs3MwPRtsASbZkfKifex/bf2MO
VIp1mZ66TX2qOk1YNxMJN+grorx/WLbsNdkKH/lgD86+8znzxbS2vZAwGRCAkZ0t
UEF+zQCXCVdmXfSx6GIEkkr6618ftRjjZ/ztvLRmPu+Mv+Nb94jGm1SaenelOfeu
Xia0vZCA52U3f+94St4bVEtRgjCUZy7KdEQoetoHiRcaJ/4+Pw2GfxE36d3hmqIM
vr6Yvs8TvjNbHrfVfeZej8KEA3pC7s9aNq3g4T/qsS3aO/bOPkjx5vlwYvIhgLTw
p1Ryq+K/Gvay6NAoGs0UkjoT1CAeY+WKac0TFZKXk3wDx11eIctF/zXSX/+7SGcv
p1FtCjz7inHCY/KWIa0YFSnPNkoO4DxbXQVLU8i35znoHqaPpP/9nTA9xQA6PlUk
9v/EfGyT1vafQklr8oCZcQ8+gNZpjOqeTxYqnhY4nYU/9sCWGCfapqZm50XjkBkx
9eqBXoApvo1ChL7a1MVVKNgq5WufN/hzFsvnS34+WB5WlmznzofCbfYZ5ST+avJU
aNNRG5NgNFyAZ66cfwviyXzNTBjUp8UkyN88ctLQYnLgjxGd2TEkACMgDMUiaJKA
z/siyg+N/fZYn6hsAL1Om2JGfRUx2w2oimZc77M4bN9zAtsTjbHwjH2utyoAH3jO
I7JcAfARPzIXu4BwuAR3628LQUjGf9C4AT/H1I3q2/1chlb/6qXXLi9FwxChxFhY
4DyW3xSTNfBdMJjRVgrohybn9A4cjIqboDQrQ9J6HEgqBTlR9UN/fo38gH1ffR9e
+YDhWMSWx9TE0/UsibRuZoVCe2xre9G6jis46CMkOvWR5ZGjOqVmhdu/QVHE+T7Q
UorMlKc5DH+MUZ7q819aVpmtA04hnFEZkLYHxtZVo7k=
`protect END_PROTECTED
