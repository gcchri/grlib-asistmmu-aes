`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dyVJo98x8hYr8ljVsNaJH2UQ7Gz8SbLET0mJjlqB/JJbojdzrPEyt4/43xqHa697
KdKai/cNm9qfIt+qm9tRdqMKVlU7QF9WDBJciJFIJaQ3vhl3tm/0cavaLXhcfdpU
ucxHdmB5EfAZBwkYKJHw5P7iH3wfV4OaR4ZHfkyaUEEMlOknU7Cw6hy2r3HtMCC+
tnzhtpEpJ1A06E3m9WjraPlLr6bdpjTpLJm/jvhp6CfdE6NVFhh/9/F5OvA/gRKY
/mOv+8bLKF9Lld11ohhKtu7PJC+IdqSGiJMYZP07J6LBe1ZfYrKZ0CsAcM2Gm8y3
w2rGGbWAt/yGmXGC560ZafFM8S0+gwZpurtZ/LuJSCajv474LbjwGS7YBaJazC9O
7wdj0R5mNhXAnUJltwdjp/eoCvnOHQE1GqOy5I5bypo=
`protect END_PROTECTED
