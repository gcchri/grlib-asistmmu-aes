`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tjEjTx8N9env2enLH08+pecI710RKUjUadcYS2qv5jwAqRgvmop22G1ZNmJMX/+
b88lCqvGHO4XTwmN+EsmW2rC/E3aauNLSzhadxTdzcM8Eakhjr9KGKWX0e4XpQqi
rXpbtMichZFrWvt0Rajm8eO1XZL4iWc3NUqa5k5+Ue1ERNgezksK28qgzwGr2nQ/
0H3KKGX/JJ1po6MNNNQLwUT4/p5y0ODfe1j1R+fZP/c2vO86n7WX0oudsbK3PPAU
T7vXivOwfnYCXd/5crVGrGFvSGPRS2FjVkef57aaMQVfS9yVL7zGJz+gHkrPnMY5
kpPNkSH21ezM71pAhiHvgOiEFZiWfgsY73ZELEflSEOa9fjS2UWEOpHz7I2V9x6Y
IlvxhKydTgvG8tMaQ6IMHq/BUnzgtrgLzO1kRJE6FgKbYgasghvZhLl+DLJgmdwa
5Do/CLBchL1/CasMV5T51EUJ5aeCjWn4qb79XNnFi7fjfYbIMKmYpHl9v2IxW0Ni
RZLUJHy7lYJ9optFC/yMd1pHNldVgPzB+0Ek18Y9KMRk7QIKYj5dpDEJVMCPEjzB
Er57ziPFIY7BmZHKOGeqpdMdGkFE4yagZw5z3/3TbG0oWTUcHUhEoFOWEdm3yQz9
R+yIg/lypjBWPH6ciqiOMqgE643jZ5iuRGpJvlI1ELg4no9FRQ6t5e9zzOXMRPD6
jPtETjfO+pIxaMnBk1gIGU9Z+JGyIm0PZwNgODY7wq3PsOZEZ4cojD32liUXSRpK
2/Xv4H3wCN+mhxjuHRxZPQISfQKp9A7rd8x4fU51R3LhGca/IV3h/+EpGYEkj4RC
AWNVH/1sfzckfQzsIGHzH2XMDuUSaHueOUckcXUgsLUqeAY7wU793EvBlj5ThWof
TD4vQpwRV1fMIHJ2WqycQIMPkANaWMsJd0kQ8KigIw3E6GVutj39KcaJoygSRtML
6564fybe09HZ+q6oBU9ubc3HcmSKsTrWR1tzNTZfa1waH5a/h4LVaO0bcIW1njth
ZGfKPSxBLF0WAWdVcZz/VY1Lp7gS4B/iknj1Lhb4b0IuAS96Qh988592awPIFlQ5
JTOqWUEAdtcs8zYt5KfPx781MxGMo0WmNeHvUL7lb5eL3jhzy+Ct+PstQXIL+4Bb
9NFzWdZXkQunotXxdQqgnMQ95IKybc0giO5yGcvbhz8O4HUFQcXlyssFfIMJRVX6
OxgoPBjjt2jAFPfNNIQydj8vEEfu4318WOxzYqxHnDSh8D6kgKAGMCpxjaCW2db3
DM7YQnvf8ZJWcW7vgUtBYzqT5ifW88BsrgW536hjY2n4aplt0Rrs1p6UdJ+yt4IO
0+Y5V2wutwp1YOicSBDif8HdOrk5DiNsw8g5NXtr/5ndpq5wI2n5NSrLDZHSD0FX
uJz+hDz+nI4yJjVJkUwi6+JeDVTi7ND1/AWxCUdRf6p/BTeLmndyR78dXiVjTwzm
`protect END_PROTECTED
