`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHL1PVOpBCrnXJxusgcazzdrN3fd/YPF1V/MfiABH8z9Q/hkvWTSuA1tS2bRtaNx
KV61lbA9fT9mOaEMzd/3IXXHyP6P6zz+Ob6kr0N2O/Sc/iJIi+3O5jrqOGvmXKXj
wz1o09uFgZwLiYFLAQ0jtumFwEnBDAvoWBQmf/yYhi6C3VIs7HJzbrDiGcrpdF0J
J94ExrXI059vwbF5rrUhBuxwBm/Sz1JteHcSVDYfbgy2wvxYyV8mHIB9q1cTmxm2
wfGh2FRCL7JeEMXiig1facMrRsMarWv0V/FhyqmeTySMgpcWWujm4dWxwLvp21EN
ZM2pG11mN1fpTnvHpgMpDnn+J2D6Y+M8KOSov82Qf9qLlAILgqn/4Pbu413yGYTV
Jtz5VnXVOkrNbRHqs4qy2iPqMIc7JpeeO3jNjqFDiIhOzflCa7CL9Qi8Z7V/fcjs
IT0RFd+CIu/I0fFzzjv6LVT6bhd+n56hwqv5rl8jrmw8N1/1dMecm5enW1hXMLsJ
Oqf/TlMU0xmQZVQc4nbq7Gak3vZzbm/XyQWA1XaH6GUf5icYYuewpgLo4zXeAHJh
`protect END_PROTECTED
