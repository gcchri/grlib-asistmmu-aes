`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJDiY0I4sBihGabcAdO9wY8KhqITw0reiPwZDL/9B5adg3z0JXJGIiHJWeDAAn5F
MKP2wuAh+QKp9xf0Zwa/FOx60UaEYIsMA4fHNRcx9/GavBZ5HbaQV0zrlruiW6um
YDdYPBKmQmMHKsPpWmjksd78Fa7JWlWc1nNC1VrlxJrF7mVjmrtlfcIKUrwvCGUn
uU/znGAgkVOU75CP4ro/TiNyHrwyJS+xIRKaawF7NbpvfpIkpzzigfOODKfidiQU
+vp9eyph8voe8Rvhnu6LBgmk/8U/5RdBM5vKTrn9e3xnVQFREnQyAzD8cXSXHuav
eGqxzVpSK/pVl1LTHd0HptpMhZp8mUZcTHoNGBsvxZpbDI61tSV3E9+bSPCVv5Fc
PGoOnxvv3JPcnCl125ldxs0ha1ah5zhiEDMMefYnsam3tDpKg1rfVEdd+Zu2zRKo
1QwErddcZa0aYo1UAe+y/VgXEXf+GbkTrvKa4dRhAw2sCDz0wz0B/WeezsEGBFQ1
`protect END_PROTECTED
