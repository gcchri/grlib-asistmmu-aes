`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4ni0bPRrS0sT+QuVKfLNs/ErdgNnwGjyRmx0BjgXV5G4gA4eidCsuW3Tn/HXhYc
OJPIKEpVd2Nm5bl64OhdDNvaA7GPYJz59eAc98fRnPKjDPV8kaUC4gVxBTCOSi8q
xs+W5uVDKq4JOxgr9e769M8pQT/S7m18xH48/qa05VuSD2fLI9q9QDADPUz2R91y
hnPOxKkBL10V71Byz4pRC5qbL4gg7rjZ6vIRMBIpfPukUIrqNeHP9kuxvQj8BHbm
53CKOI5gWRt3mOwHsrZiU8OQTBU09SbAHhUor//69TZJ/Avp/oj/5Vzo6Wz7oZC1
3GvM9wV8WxhzptN5M1QIKCR3QXJ2X3BCrrf/RORHyN9ZMtGBcnmXJEbYZm6+zUmC
UZbflZeiI0SgHdrxxQMw+BmjY7LkN0GGGYD207BmA3EQygx8s0Dfv8SEyvXdXhCi
sTo8OU/2B0iTNshkU8fwOEfBCktLuLLT4bpAVWzy6UDLlC+5s+7lWvXnJaG6VzbO
IeY9tsGKwAYaO6G8syMvdDKZk9WvdgcdG4FaSl/GfupPi+IG5BuagJlVpv8Ke2bZ
F3MhQXDENT6zxz7rWnpC74zkrY8EYOyndBnG2wGS+SoMxMW4g4LFnuVCwPFNWq5f
XLlOgBiNGFJgzVou0TUjFm/Y7it2jHxsLrUI/BZIn4B7AuktrUZXdW+p+GCE7+O3
ErBv9dLYxZ9VtMjuXk7/S0i0N6vy4VpEEdH53eRQj44ZFTyr9KAKFweo+kY0VU61
`protect END_PROTECTED
