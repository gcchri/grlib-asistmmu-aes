`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nKAD7dHHYmPMvSbFunMeiUaq0TOmjXiO64IcpaImMTdK/ZNDBHlVs2oiHoBnVwai
lMsXMUh2p3E9RZspivvJlMhQuoJ8ghCej5zslpjah6PCapEfW42gbspj+6EN98+A
ZNaPLEkrXVwtCYj92K4aF9CM3Ajsm4c+1nnl1kRcvAuLxC89QD25t/iC2Yj4zO+b
tFkQ86W6wvbUQIw/VW3n8TLZsemVBcGL3iWqCnj1U5jVCv+72r9uklZtKOSzmJ8m
ZL1EUBDHoq5jxlM33Cnaq/lwj/hJzkXLZqbacdJRkOB1tkZn05PNnVONF338ofc1
bpRtFcUgGWcWWCtO91R1CvoNIK2MH/x93Z0TW7mkmMlkbtzt0YpsK+2GIPdG2niT
fVrNZINPrNZ8WfGh4nH9dT2Gy/rdk2HqVAiW+Ma9MzYtjGAky+SHE8liaBzSKVb4
zgo4xQORZ830i2zCjzJUebK86/S29qxkVI5aXAHT6RsuYz8ii/4A0hKwQJIHnxER
apedf6EF8pfL3+eKrtFILVd8QLBH7TGFfMCKv/GyeC5dmUwVnUGkRflOwdVKI9DK
0wy26bS+LYPd7Q64MUehk7NqRDQ092K90N+3+xIUD4n1L3DR3PSHtX2HahI5P0Hz
zT3MHVZmho+4OXUISV6Vwl3C8wX/EvuGh7HbGC3FXVKdnoFFt5ID9hDKuhsGJNf6
cuFbPzBOMBlA22FmczlgL72OTShIuF80YUhs5tRJAb3hsxSUzyL62rMyVGnF5g75
ezUBfYExQRJeJHKy9KpU2g==
`protect END_PROTECTED
