`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhAWW2EJvrNM08aubbbQAeNvaFPi0iOOD5rRqCCAnHQWmYy4OrwS64PZgjfKk6u7
i3fkNFw3cI60WqzHVWiF6nGayD/zVXqDfBLhx3D0ci+6TP8+jc5ZdDX+jzNcJD9F
0Yt/+8Gz1A7NdO7hwpE7XQBexusT7+pyTF3ZGUgRS/+aP95dYa/tNl3nGTHke+M3
jIIeY7WTI7L21WddsGJwo9LM5pTcrPXrx3gX7zIfRYoob055pI3S46GwdFXtCFN+
CUz31fdW2LvmRw0DYahotWFy9JRuPr0J6BPZaXr2SAWAE5wskCVjMki1MNAGu1/5
IpuyOHLZqqcOU5SJcGgPmelRdiBUNdRlN4hDhI6az58qiKtAvQ8/z/xzQLamOiMV
cjire73ZMJUIgwSkvnUY91anx/ral6eOieZHCPQ1iYqUsitYg39Ch8YzSVuukayh
YRZSsvVpBm00OMTlNx0/ZuCK0RrXHpEqE+bhDstpfPMT9L1q7RhTBwJ/l8i7Dn8N
oPbwTOTXIRWQ0wYP3XWbrJRyDe+L5OX65SD3RaVjfOv41xyOkVtr8edV1XkHYBJy
KHSZc91utlSoHAo9sDv9PxnHMwH5yHh+pW81rDgp5PIPeHk9s8w2eFzmc8HOYCwS
8GRFWFnfwepRtlqx5FbcLA==
`protect END_PROTECTED
