`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g9tFA68X6jZ6A56O6P9XRjD1CXMctHI/iJgcCULSji1Tmndr/nvTHzXEnICsnjMf
rlF+uQ4Neyff5qD+Hk1z4nSB5UqURznm5pqE7PuNOLefQF3imG+7jos4ZQQWUK8P
Ki+J+z8Cuz89mPa8yYrWQcUbhYbxNVDDDzBliFJs9onB/B5+WGDoUk4X87EVRPs0
0cuLXZg02wFnFj03k42Vb/Kuxt5pgnu4/KUkrktTY+7gdwBP/ORcP2silf+ZmjaE
`protect END_PROTECTED
