`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnX35Fiwfn0CEMYr1PF3gVF/9B6UeN+Hk28TTWlsAO9z9lMmJoFjsM+2G0ck3YT0
8pvXI8LDggrEns3v9TYJODPOZml39pKD0GqGpc6Beranqo1BOMUdqhjqTGsXMOtC
H91A7npuvCIrfVU+av2Cx/3p2ClwsMg4Ol0IOLBfUHygsd4y7x2bzb7c2cchf2Nh
pBueuHyDsUpgHRGykLtEdSUAA6QpcYbIUwDI4Raf5+xlt0pfNmoCNG2gePPFWeQg
5CzSEjQr7ScZf/rCGkWuLB4KwdkBew9IMYiKrMB8ViWRfBJdwGzmsunRB6h3VRui
v3mE/DV7aNJWrapHUTrgOTMn4akg0tZZfu0gn/vtRFEMoYFJwB4pKBJpklINdjcY
YBqGht7HMGfxudZlgzUxCpdz3ZX+7ilADKMKGs4V0dmwq16r8GcJPQa7wiGWXvEv
zrCn8f3tdI3KUFmFXaX7qdPqd9KmoS8Z1bUga28mqWYFKdI1EKheCdPfqYdwOnCw
cxxV8t+/waIY+VCmsrE+BPwnjSfKSk8J4L0fbczn6GCq+K7pNf0E/xaTNRvYU+bV
6ZiDp9Yewwuv3ExpmaNYeQhDj5FeazKdDKVl7Wxh+/TCRkltjlA3HBwzGjAzJICd
wOE4RSTVDaGDTO0H585axf22vrVR+6sdztvYzGapDGL+48LLjHyUqDASsE5K0Uak
vt692UZBOg6n34EZ2NVDah4CygCVcq/pO43tMci8DMsUn7GxxKG8ypr91JTQycLp
MGmBUbNrN8Qb05GeoI+iptsd6ZRq/X2JQDpQIKZW/uQKPjCZBHG+W9JKIy0LJayj
gFrSbRN/Dwxl1ZC8dQYkCQ==
`protect END_PROTECTED
