`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZiyzX47HxvmyFU7If+uzy/ciGr+GF2SRcmdhKQ3LgEeJGI9uL+2oFXymrj+EBxF
IiHiLBPFq8r44NgJF6UfOKVRSCOBfLdzNTkNPin9ru2OiQJnUw5sTER/jMqUDViz
j+KTFCtLOdsZWhcVa8RPNCAglPF1o7sRX2hfyNlJHKVa6UGdvu6VhLpxhu4Ku94x
/KT4RuznXJf6YqkNU/M4+ddQRIPgjr+MTzxvdZsGDdFYIRnbv7EIeQAVX/b7dMyM
JqeY+P970MFFTeXIJsvgKZysq/u5JOr5cSSWkqkBg/HHOc+LI36u/+HSDJhsHLST
U98Lsz+WRiDBC2SecybMS/OxirBJ65bl6xryi4+K7gMEpflEmXUjQtUE0ozhJ863
p8VLhCLBNJ+e7XxHQxQo+h+1tE+l6gRAIfmvwtzqHCDJHkVhF/+A8kGzMH7xInx3
nUvcIsE5Gxrw8mxHAOXELywULVws/r3O+Bc+lNjH6OnLHKFjIciKJwtkpgoCYvS2
KJDYoADW6TDQHX0P8HZIRKWw1EsADcQ+I4hrb0TokLoW5SctOGNEqBoHs8w2jvkd
WuUX8qmfxdi3mFMKlb4DCAY6IdwuBpJMI+R9GBVfCqdBMnZV8UVYIwuK+4hNnezh
24B7J41weq9mv3uSP4cjew==
`protect END_PROTECTED
