`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZlxVB2FYum1dXVRkYNREKdehh5TY7mVjQesdX2ZzP196d3sy/+s47QVmr2kUNpy
BzCAzLJuxZKLYLfqa+3wPmJNJZw8L+3DkqdR6g56zkKFhJWRzEqqzeWasmz6ZM/s
s3X3XylE1dZqyl5skxB4rzr3L7pRUWamd6ikss32jn9wXrGZMmr1PIf4gHmBm6T4
y1CBTikSuB6uBpr5gsMipQLLXRWb5+uBjiqzLsjMS3IclSXCVPhr6CqRmNPbS8O2
W+Z6hivKtrS5ewVbLyTiYou41p4ORhJavQm759u1IK6TP3JSZlfFCXKIQQg6bZDx
5lKVCtssZkl5ST0b6nf3rX3RTjosmnHdRiJ1zoqmRMC8cg32ZdC7LfmNt9plIs35
jMINLXIVEuhtqSh6k4j8Ao73/xSf4sO9b4s/hPl5FnqrEdvLfw4CQHKnWhnp8h9y
sRZX5ULmLNuVyaeBXYPwlcRrHT/t1mHuGtaf8rqP2mFq/9JCTWFqyuYnjz6QvGvG
bA2Ogg/L+fmlvNgrzAvt5N53m5DmrioGmtBVc/ZnFTUVh72yOVtVhJOgGxS4UVLU
7HZz/K6kIlnNFefQ7nQhEmCRNepudiSRDNMqtp+Fx7s5Su4OvPK44YHNSrxObsez
vQOPHlfJ7crNF4ZlWAzgip72KDpWfw5vpxsudbo8NlWGQ8pwmbZ260W0oXnJx1wj
U208amP9m9UlJ3ZxP0RzCE+7xUZGlDq9fu8dsddJgAazMzNIk6PIT5AKlFQJ6oL6
o4njgPM7QGJjoyFDKKibZvjy3vaHorh3rMTjqyNMA9ugXbfiFTKfi+6nyV6ECiVm
h4U8HLP0uodEjFVrBitOyKNp2KCwLWKtQNGNXp0sfxD9z4aq2dAFQpA2f6jT8DHb
zEeYI7C0VxR6CyW576rO7904hdTwsLfNPYeQ3NxUDw8fstqpiDDoB1hpJID7lUDr
Xvwzr39ReNuuglIzvQa5wRSCRiFBAk7iYn1K2PkT05BQ8mZe8ugmtMZsps/hiQHU
UfPVU3L8hIrZwNOIpGtuBgCQbB828Q2ow9bWH1suwJ8yxn/4ryg/nItEAhN2eAes
/ArSNqTe5Lv1JvOh/5CSlnSO1qtDRd+Eel56C2hdAi+R6Cr+VRTJ//uwMRFxjDPt
yn2U/YErfSukel2bx6u8gwRd4Hmz6pLphC5KI29eEiWJmNN0LLKqZWCM6HJgk1Vp
IWY+MDWyRSDxcaLfLllENG26AXlE+etkb4od8PkrxorDGjNfuXz/GglP9T67SCtE
BNKI9OiDRFLvOGWQEKgdbaIgNf7QehZnWWMQ31amIPINhXX+jtXWnPt/MYsywgBt
ealzLX6Uga6GSQdMtu0uTZJigFBxvqbQAYIR9wPTCvzsQVrS0w1Sx/o5hLqyltml
WxhnDCWG+z7i8czT4f+XncbipW461q/PFYsIO5FEsLBtil3xCbQtxjtFF+jBL03x
fcxUofun9n8RZToA+QUF0SnRmYNO13ccNQuOTkBtx7wPxsKYknoeNrofR3V3cURf
K1S7EqEJPUFy3Fw6RcQFjoHlKWj1csDxDGsJFrPuFoULm7u3LFiZIp4KTgXjrSTA
vq+tlbhhPKDFVnuPg2lhpU/0iVdRaaD5pQ9YdrC0vWnTO8VKSjY9B72nEPC8a4EW
Ah4v2O8lYfwflFyehlxeIJ0RmXRB7F0Uw8VvZG4tf4ioYnJaGt21zuUqbhuNk9y2
DDl2fMU/1TN2/PWsJgH6GuOQKfxNT+JnI4qdCVqODz8tTcahrpTyIK99lYnfzIo2
Bkxk/Y2kbLjhmUr5opf47PORUerKebrbpLbc9wjIk3xukW+LwjqSLeB52uGT+gr0
zrp3FK1caVrEVjdPOizdh9d/zOHA++BM+D2bINYJCAG+kw/EXNzYUi8VnG2xpyPI
4clCxzA4yr50/y/0uF1/A0LN+1Mdtg/T3+I5zRNkNzmidi3YS83TrSW2xOza9lb4
wtxEkJ8Q6tlGZo1jbIZwj5Rzn/SCuEZngJHg9nQX7PmWLLRDzTcm+6Lt2RBOTaUq
5jtXoNnWAS6PuUxSCUNNinivbmUMvau6abs31bJqtkaV0nGL73XhuoRNytlhgiwI
JVV50xrF4q10PMcMicxMjrcsrcUfjKQJbaugLv0RWRWsqGorc9EhO+MxlF+WQlPA
fqCp8Q07qPN/tRDDDQ/ns5XVqV1cASH/ljxWNNiu0am0ETIUvGMwjZFXC1XfVgGi
MCUwuFpKwDDLHgjED5XM/XouLjeSW7kjObkIXDeC9hUUyAtRy73YCvIifwnk4oxn
9RR6KnlvGMYJ5RB1WK1+7BnSoLtOp9xcqMqYEnza5IIuq5xMnoPvhosQ5lB33uP7
8UUIdELUri7xULlNRLC8DMvw+Ldg7B7Erc+Q5CYiEpJBK26QDgTMwdkp/F4YZ/U+
nIfqIxLSFI4+fSy7JvGKCluHTMCIzhsY87F6EdZ9p+/OG3Y+fHXc9lkeeBTf3ifs
kNcRbLoHhiReAjoCcxIeE8soraH9p44eVr7n9ePwgv8dGH8CKWzVVPGs++YHZrtL
HqlAFG2EdKUxbXZiysUyD4s6j4I/my9FxLvF3rsYGQ0pcPE8VAf1ehVnbcfoTyYK
16iW6WDOY3cjBCW5xRiIwlmL1PlwUwDdgkSvl9DdHx2URXQLXhAAxbhN155CKJbV
AcZ0elHyGq1Hu3Dze3xUtPT0Gp58D5lc4l/yeGKu1Fe5E5ALXyjEqSPj/IwmWcBi
OsPXG8tcqNAV6gIsLiVSx26MmZq1KmiKdHCRhjwGV4nrE8eW11/4riLPJ2KZbGax
bxry46HJit8FxoNFaibI7KPuxYPv064qEpbKa0QnFMc3MQkjQPJXackKiYGb62Zy
YB1VMmMN3aeYwNW1OubsP0kKJNY4s+iqAD6VHl8ZlABAxGb5K8UfGC0JKh/pJOXb
tgXmktfvNwvQr6DMW2ahF/Ont+7QyprfEMf3fZRoNlBDqh3KH7QkPM59nzMAX3OT
jQk06zNjEgIf9jD0zVOvbqz/4S/sojGKUpvdX9JgISjUmLt6NTx3IcJOBr/vgQrd
4QfB0PIXwjS85HaNKHjGLAeZJ8vBVvbrNDn4rsr2vHVkmwJ2aqOKssfzGTQiwmG/
2YK6xC4s6vTGUsQ3XMrt1FgQIQCH4oqJUNnQt2c8rF2FlTnvZ4TmQgiKOK4M0cfU
LLS2OGizafzgSw3UfjQE9jNedN+zzvHwFWm47243Dx40WOmO1LuA2sSGG/iYeT5y
/Fs0BYUMRDzvvbopJlrMJrLRUO323oh6NVUt3frmTuGywK/CfT+owDT+7wMx/iAa
DfRV3ub2YmuJY41DUQCRo8/93A3m7Z7KP4umnjgAjhge3JlW0Ov6RbIqypIzly6q
UTY6E7ofpsnO4LRnSUk7Efo9Q2FnYndcfPQivqltlhhNnjNp1X62OaexBWW8TFlQ
hrWv9Fxkg5QEa7S/50gjtGiRSIonrLkpbAw7fT6ym+fGP5lGgpBgxa2ztVeMc7mo
xNBNsT6X1f6/v7LOMnbFlMTKVTYCLfhW2VLk4v4oaSZh9TscPryBSRnUWFT59vnf
VeXhIMjRREBpAHnIwLsObuNRVtNuHZ2jSbFRkzuY2fcVB1BebNyYwJi+j3x6cHj0
jSX+3GZqS3hBwo95q3zKnjm0evKlJlS8SYFNM9aDD6xzgtuh8eR9VtHa21CVyL7i
RnWbeChQ+nxrUOQ95zBopEbUXt/u1/fs4FEPWFS1FZ6q08WaXvWuTdcUi9kJkroy
EN9fiz6I3klixzQ8u9XIGfLtuw2pzJPA5div5qSbQepesJgTqFV0riy5AgTH8nF+
s2++iDMugmRAX+yX1XRxUmG4+BkvQXejAxPaLPiZJgSMOZj4xMOStZg7gfituMfY
E5V2dAol5rP93CtJkk+NxT2E4OBPRoRtmMK7Wh0Gf7fiNf4pVDINtQE6Ct39crj5
m6V4LlAHUXOQKXhbjt3r0h1lvCkF6Wk+qtkiHFEetvf/GMHsFh5l2yY651jPcRoN
IhcKWwK/qPIBvW2bBMKOQ+iNMeU/xQ7hpQmORwy7flAdLDu8X9jIJbvIqqvR0x6Y
hoqrOms4JRmcRt59PvHlpypydjTG007GBcaqNOCWSHmXZDi8NYfKp0E/lzh+7lIw
HKdAdibKnIXJcxTovjtGVSWzYr9JoapeEkGT3Yx1K+R6bWT4GUekQJYj+x21G3tN
qq+pqWG1wQ8R56lnwWd7OJrKaiWPBtoZlNxrgkZa7alOcOJXGkvubQg/PEOAEqgP
UBaHlAtKO0gjTeBpfOS7zQAe7liOFqBIgfyyjkvs4OQedIqJMmWIXX8iPLXfPFdz
Ml/Sa0nCWTVC+MHBZS4X+O+JX7lNRcku3wh/sLee6Q/poUvBC2eHGwc3M0Fzuruj
VoLRJePOwI932pw0GQUoILI/Xcd8yK8eOgnUQSUfKI/doa+GaqMm4nPTABUCW+h6
NDjA1AwCC0VxY++lbfifRAtwqbC6g50hX3daXymEuH0000VY3dUJMEWtwoaULShx
Z5kHOT4Z7l7UueL1KdycH+g3+k76V3Q/c1L4f7HsuEzgQxhc0pCx67d277eVL+0N
2i3HdZsOYG7NMBz8Li6UA16MxjO/ocwr+tXrZFrO7GNseUggO5EsoL2IfgMiJWDs
m/WpzzBzBgTqOrKLMkS4AqhuAon8iY4VULx4IKT8E8fhcR/0SF1kRYcWBrwfHlpc
A55jYVPmc0hZauWfrb89l6siPGvI/eeR+m3UidXsMyMHBJ6AV01T8LPjNifRshQx
VWeLZsG6AmMUpkPmz+yTqOZ+A7ry+zJ7r6hqr+rQDFFd4wyrJLxf3En8VeSbJXX4
AmN6bFWVDSNPHIt1z9kvwCNB6nSzdPYURpALebfBb+kih3hyd/0YeIGp0dzWtkAv
bwAKYN3MRN1VAL1P6oSTMgW66d4HUWCurT2kN/Wy2jU58GoerqHrG+FdnV7g9lbC
pi6AHAXQvtUVdPmnTlKL4uHbOifPlFyHxRMBVjLGet44cFlbcZRsD1xePr9abujD
6B7XVJWYRA4O4l7p36rP38Plk4ke2NdF9QrJB4zs1k6rPehgEAOrkIeaFLdu4kCq
2wI78w/PnoaMXMrhPfctk12iFymZLK+xmFDDiqdqkjUnBBfByTCS1yXLJQMkXoPS
wFvL+MxIOJtkEqmByerHQV5SDglPH5gxSKD+z32Ws5MNdhzfc3Mmrq9F2D+rQ0QH
i9smfFvjKvFFx5cnxBLXy/JeR605u7vD3iruUXHqrFi8DGP6QcixclAYKu17z1Mq
RRLwKogzJGdJpGvIPUafskdAuDTZRkVdsV91m9UjLl6MpHRUllxATEMWFTduQHY7
9GA4w1DcY1BnlPMrmdyP+pG4lmjxpxo1bdeT2aP5YG4N+54n0PEIpv6haXsc1xTo
JqZYZK4IDqcpoDfJlczhcPMhyiBpTrH+/yBomU6oZypc4l+KGCIY/LeGgq2sE3VS
BHIcWAm+J4T7bgJcVvZVxHb4XoKr6WIG57wpLdLlxSQ5f7nnXQWP+ZBz9WX42c/c
lN9n4V3srxo+EkuoudcLGVfj4b68Yx3SYG91Lb2KOm5DZPZkNl8j86MxKgjIrSge
gr5c6eKT82KaWOZSsB/NhQU4Lby/XZwpC/1oNlKzSFVt9bCZluHJdEHqbC9Ose2u
LILBKYHxHexqjenUxc4SHxCK1jVzHc/vYUDxAjPYH3MekAmn5By0BRn3+SZ3PkU/
C0piq8g3WMQurgBk2Wi8MOrPcbUQboger8hSB3Q4ZMzwnLznh2qabuZIwObOIlPD
vyq/WuvxOeSJfXKFsaYKzAzFNT/A/L3LQAfi7bqebPLcTLgimNngpWic+KbGyTlf
/RGBf1+tSiz3vbQ6lntizIGk0RdpvrriFe8drtCXeTctj50WNrvwWa0UlDkzgke7
BTzz3SyKMWgc6AKj974rTKPZ/929ye+RpiroUSLuCZsvAk7lJaWTD2vYo+NDgVFY
0shD4KmDplFn96uBesgWwhxz/nAv2E1gF2mIGE4DSDclxSi4ppLQIuOWpN6F304B
9UvRiomnEWs4OM7FctKxKtxa2h3IQpPRerF2SqQiLXrJSg+6Z9b1Nxw39SUm43OD
uMnf/DOQK2znqPf7zF4waxlsadeSYZppxlm++7LF4LKKECmqdIRBL8dySE4mVhXE
l+WeMvNcO3zGARQ4w0yeMrXKU67RywgKRveOaqvsjDhN5GZoMC68uXOvly5u4Q/C
7t0Nvg1KZmBHKi0PX7Jhu4f7P2iP1/evqenOPuAAf9mI7Qf24znFYSIvmWXu9C5D
RPx+p/g9MltDrMyzPZSapgmd3BfCdpvHXxgPcfvzYKh4xCuywGgeFnRaPCxXehVE
V1vlOSRf97EW8jqIpGo2LqzRcjPAAOG9INpF+5vrMXf+zW0bGd3G1E3xnjVcztIb
3pnRU7wHFK9qMZd0zwY62UK1lpJz5dQXMiT241lKDYkaPmI9vYgcenNwdQLdPe+c
TfLhoXDAEJKf86FYusbaCKiWA66AA064jf+nYj0EEVz7Rrb5Kdrvo2HPp4/VksNu
JEHUqe7bitYvq3s8ppFTaBo08L2HLo93fr39l+bvG/HPCSS1bJrN8zcDs7aCRzrN
VwbUC0OM4KkObQQsT/E4alDn5qPKlkvuym3tcRPuGbaNhN2Wu8SDkzUZViC4L+Ay
6IeuPZNoynir+Tel2nx/TdsjPK9I9B7xbe6PpCFsF/UUMw6aT9BUAy3d/l23e9dX
aMo651eyF1lJMHmrluc0LJYnPqx5olb2MfUVsKn14MCwFyAfYBQePIiTdsyqoDAL
WemKsXdqZRwS0YujQ8AVjwaMYROzYz0gvlJisySZabjLyUfnE6iFHgJxcpV1bfBs
suu4uaKYwF33yImf0qxBFTvh9XIwknXgH31C9o7ZDMkEiOHyf6+V7lvF9Z2wpUmI
r5Y8Q5z4WEqyzwvMk/sH1zmPbawUWMTQV3iPRNk+pUX6AfR1/6VhJkeIhuPD4toE
uTCIAVa2Re05kJSAPt8lErk/RSbk36ZsoEcM7Ok6qD56g9Dojci8PWmh+SHmbV65
bzbJ3jerzW55KqIHjeBIvsa78eqfhhZIsB3h+muzQwdBCt6P3Qo6SnrqR16cLZBm
OoQOBwVz3ZO4C6LLf6iLnsyGUugYc801FdJvN8SHhz3TyjneD0MFLQbNNQ+HbHMk
6gUphF+bs5dlKBKcvEahLivtnRmdDtBKH3AmrubgaC/yloTacEAWuWWu8gKPGwcw
dJ8BuURMTJML/2WxoukB76Xpk2ZXjAoG6FmMPqbiLqs9S4CO4RO2OUQn2AE65cxx
rPdNHceEOJ8doYvxsKMrb0pc/Pl9UYwisdSU2wJcPtoFmV8tlI5OauIPkjs5rXtH
iNF+jgXhr+ZfhRXX8EyhulV9zmUiWpn0fU37WJVnYAYG2YX2qgvcwVIcJnNkJ9na
AS+wxl5/n61SkzLDMXvA+LY01M7zLt7RS8zoX0nmHSuC1IDKNt2D6Mp6HHjDUi1X
zQa7/qDJZkapIX5MXfOdOBKzVRw5H4kRSn6X3nvOFZKgDiZAjljxoucxtDTmer7e
FHkN17HKFepjeIbB0BxoU/4L9IrvKePc9Pn3PDz+jOjD3s8/H83NH7wIfGmA7Krx
I/J1s+RqyKRoS6bDh3t2sMdXFNDSxL62EYlqJq4rysBs1df6yMdtHGBynl68xkoJ
jbJbFyQYZdHVSbxCworf+VbwIhwLn07Mypwj7WoV2VyNecynqDXPldEUXxjZocXz
L2iz7DKCwmwkZrfwTyYNWAIrFZEPflriaLawuMuoSxcP3pyWJguHkWiwREndJq+s
Lc6u+KTioJoODw8lOX9He7tZwQlJ8j3CR7OeaULfmldgQB7eDsnWF0VqQpTpUzuJ
n6YgNteQ8kdJimHZJc6DVSyD24Vgdh6i47JFvE+IVUnn6rhyMIQ/GNVt8TGNnyxT
9nFmQ7VDfiNysu9kMTgCahQZazPN5LF+yORI9HK2xkVcc7lgCCkWlOwXxMouz7aT
4HAQ6Z7b9Jp1rxxr0bpaYITzw+zyZ6cmtJu5bLaplXtI3BOEdSpCxTf/A8HUA2FB
TRruA6kapxpuv9588YnGXpuIbaRAbeay3ADA02UZhmcdK6AiN8iVBVvnpVvAOArx
zDYDrQhf15EZIHBJQAZ6TSVWbbQ5MsqggTfEHd+rhdh16A+afMiWWR9WZO+G85sp
ISd9zuYipElfnrs7/BcYJdRgYLPmOCzPqL4D7I7vC0G883qyRyYUFEReftRlq3in
annbJbE7CwxBQmUdLQbxGVdbbV/hY6tIvJXNVsNcen6nHGK+kOxEnuZTYuw9tVgG
YA1esvn/z+b2Dw5WC2uLe37LXg6Ty+uPLV4kwPLSjfarSF15XZSLh8X9/pEMH88Q
sbX8rT5c6ABusAve3hJwNXNO9JjAA/R017tpU3x7zE0LjzSoQm9dnQ9pkeF0TbbL
aN+J3UTbJXn85U5EM/eas8tJsUyct3p4eO/93GtJtqfKjn6ZIPTokKKZ8GvBESfX
QU92xth72UKyR5oSaBTtwhzRWWyd/+0Olq/771Irhrd8+3AYj0LKSs2YkW/ZoVxw
tAw7p67TGouuTG0lPGjT+7iT2ILk42MFYK2px/e8j6Ww2lyJ2R3J5vf4q+435UrM
DmLaVe29pq8J2DpiDpYmkHyNqFgXoFiF5eWit8bm46p9f5BtXgFG2DDCxzAgsdkf
yOGAwT7uH1PKTYT3vgIzyv+q1OpG0kq4TswGKnOtYvtkaB+W9Mew+2w1kC4zrraF
YZhNAHhXDrh/GSQG/+Un2uKn13exzigWT5keszdlBp8LKm8M+ZOBsdpg/iveE2UE
Ji9hRIJYNapE/K/vG9FMxLZu3WeWphZDILyiCwz7H4EIQefj2Ze+yiwGmMLHSjkX
PcUrpD6zVsKpWeT30cP7o8tdx8WOoDGuHAbB8wJIrcaIaldUZK8dgPmBMOeTG6M6
nHWBFirPzIvLoYfxyt5LgMYmNyMxbGVMtKwsWSfKPy7OHmGXYww1x6izMKalZisr
idjqzVfnlm2/+J3Bt+SsWV8UMI+8v3AE1n1gwn/V3DIjlxvLT9dhnFfyJdFo4P4L
yLTIsBzpMHo2L5A3pSsQze3AmNlarS/nxWI7T4irfuI645WUxLZ+uyaloQdfftoi
8xcMAC9ezhXZbvtQzae/mP82y/eDAQvO/fMPfwMW/OvbhokO0ni+HIIfXS8rCj0w
o8oZ/YHR6smisQDK4w4FEmN8mtML7d2fN4K9WqT71grKZXq0Gji0ID46KRwzQLB+
236tew+pDWa3tS3eVrb4XV9XxFZqy1FXSKAf78JfyY9/V1nAWARvAfvbMGx60/EK
s9SxeaycieKkztMCB96QKSpMa/TnbwV2jFpARFRmb2JK/AAC7XS1CE9fBDJIz1Rh
+GgufDXXScgyYoU97648hxEO0MtiXTgEK4yrkEEwPqOE958Beh/QyVv3tREomxwO
iXSiuokdkIfRAGBMCzQCKh/G5+EVlKpL8NH/fek4Cg1nhqJa4b8WU4KoPKuIleTJ
DLOxJ/i+1D1nIjU7X+4KE6ErrffwI0dIwD3g/Cybm65Etnd/gX2C0IwA8Y7GGeYU
QToDFbUSDAY6+B2r2tvVitwtUwO/NqhsoAznCmmzD1vNpBdsBcS16UzejVAInpFJ
n32T/KC+MF1dHyGVyQ+JzPTPYwsPvx7QNQONIM66abNEOG9gicMqOFiePn9AF6R/
uhTai0zfMWS470L1o04BqpX48/xHW2xWU4wES1CwZeAlBqUSFMteUhMHVjiZsdsd
RW3YunxzDQBJprEWC2mOW4T4ljmByqEIyWg3xZJE/GXNX5R3DMKRZog1of+jD9nI
H/GbtX4dtGu/2H5OsWe/HxOU+CU9r50z0u78PV+a7sZzqoHEjkiRXp35eP2YYRbM
XKdZIBU91gV/6NvNowC4Omam/9T/ESezjgqoHA7qXAuaSHw7jB3KVdzH/BaGTK8d
JAm3N7UShKR5QNT3V0vvnIOci+2rck+/TfuVWAmIW51I5QS8wd42iQ/8jx6BJPgo
OWsE6baOlhqm5G9vQr8c8o83ud0COtLvp/XxA7bICwS1uzUYTiI3b/WjgqFf/qOo
5A31pceEwxFYwu5TqZnKsh7DVhVDtJi87tQPNMrf29/ncDdXZHdPlqoBTEf1EPnY
bxjYTqH/vIBjUW/uN8ROgoD563pulezxwsVhhjPm5FB0xQqodKswxNUhjiMgijyZ
nE5/EDnx8ooc1He5vPfQlSDd9g9yX0zpEpBqNr2O0T6vDep5Uhj73+qXoyBZzasl
uIxqFGjZHqE4oHIhOO83dRZOwuTDdKHLEiW5ivAdMGIVZk/Z+Jvyz+6A0m6Lt2ic
SGnoE65ZmznBpDV3XrV1VOmDqy38c6FM6FkJwNZnZhaUwAtkyIEq5uhdBli8G+0N
3ssMy5RusJfGFzvgcXsUH/Lav/sf0WGDiKZqzRm5TdA4r7cPHbLTU9umpPllVRPh
XDv3mHzDpqmsf0+YoTtQQxZT2xXTEffEl7dwzfFubOhcwKgTqOMsqnoZEEBPFi/3
5rTgp4KAxMBiEPcKiFedt4TcSQDWTqLhYW7MH92u5ynV94Sr0VrerilyQxwmWXnm
PT9yOXWVOzSiebuyt5kC+YiBiyVvFWPMhEhpJM3ETeRlWBRVPPMJQ81xU+Q15mdm
ZyPisntHFyPn4Vu8ZMjv9Hr6sP9pLYf9iqIbyeTJlPEDVQ671V3CTzY3fPPYqYDv
bIuRk5RSiKOXYX4l0eAHPqJbmZAdCfBZlACf/Oyf7wCMlw4VUDPwGAwCZnpBhDHY
9rrbzz/p6/VLy21sqRt7LlJF3oQ4euVSb09fslPQPsbj9UIKklW7ppz+fnlTaS/6
0NkQy1aJd40XS2ZB58GEcKhRFzPDjdScsuzfsL06YZ9qLbNc9F7EpQFRag5+Vu+W
RyGWjMdExMrK6f9oYHZ2+7kxug6m4+/W+FTOnE2PQBTQshOPq+MAywaqz8YoxGCW
G3bhIxLU7ICkuxm8tMs4XhsggESWxgy8bp3RHN6djxi3pHshUfOOVmTMBu0j0KDc
13hwJgC109ta/RSI93KU4Ar6wIgaphbBdIR+5CbXP4YLLdxhCGQ9x0J9Z0GgQhuK
cwdLeVbcSfTEFhiRiFDVMYOSjQdMZsl70hdlevoOp5iYskREJaXkn6zmHcn6TurZ
smO7JtAgjOJAp050mwQlw+Snc2kKM8zBODQhZZXah1iayFyVJxRCOFxWh7GW+TtU
S1PED4alSkMKNkqqBTbWr9+Qe2ToM5bhy0m1wNNcgMEQNHx9nHBEH+jGIJl10p6O
ud9hb+tz5UlqcbogaYwcWAglGwUx+vjmqTkj7VmE0bH/9VVEsvhluluei6kMINZC
NxhVsH9Zg/ObpTECooCjqktZ4JT2sfE1JdZbFQy9jkfUBlt3SIG4PUAUKb607Kmy
/A39g+RxZ6TclGAXLjZ48UfIhQz9+y/YzI3zxO8kcs8bjXPwvrwPWT2eEdxcEAsu
8a33y/DMsNe/9jy2VdtSqKPhJs/NPbK26FpBVtsuTEUd9Pi18mjNjypynMCVmBld
6vrmK5qj2hQFktoN33huep70wb3M2NDZ8BTmW5Gk7ypTCB/LVvyDPYncJOJuq9mI
2g8l9G6r15AXLAm+LLX27v+FFqpLT7MB9nmmPxMZxRh4gkoTdmUjXXhFIFca1RWP
pn2NkUfy6BqYmMaejZW2oINvxzk0J4BBM+z4iPMyfdKxMPPF9Ha70tMmeqHm7Joa
WyUmddRWUPHRCVMpM7tMcz+JDXG3W0gag2DdVliEL8XWEjSVcaJs8T8r8Fui8yFA
dz+nV0242832tMWUgqa1mGz3x/pSVG7ktDHOhBCdR3D/0WfYIC4/2IOMUMr5IvKd
EatZ4+8PcU/C6LPaiK1vtM9foLFCmWP51hA0xuYMv2/ZW4SUu5agbwM5Gggo9wwA
gxnDW3eNeOv9HyRrKHgWZBz6oXjHa1VCnB0MOEShwHmkRRmhwmO/QrVOzJ2+BxNG
1BIK8ya/k9BmSt9YTfPsjEKmFBE0Luq6edyNcb8tmgyJnBPa4jlhlf5+sDclE1zH
eeeRagZIUeWhS+aj1086UpkfHmCBzp2epymXua7FmlGeuJ2tS0M30Z11Dsh+7D3v
2SlFVpXUrgcRPRJJoEmR5un9I8Srh7hhTViPBOUdlMk6495ctl1xNfUepVT5o5TC
h95N05H3yiRCuqj6N7/aa4hHlholgmvuFwP1MVmIXcfrixjF1KIUDaxaUOZreCrw
bh1/gtZuqxG//AhrkQ5g4QpK3EjQpmp+QbJajFIp3mPePduGyGzmP1C+NYdOajxl
du7hnyBGpqKFEWVGsIfh767JCqEHJMqo9t9st7D5mvitD/TLqG9jqkXTOjFUYshx
EQYRnyM1vv6FcRMhn8c4pizpKayvIpX+N4a94DK8nSkSxfqzXELrN9IbDQUirUBh
67Q6r7l+d0pMwOV0hTFSbqIm3HLMGXDoXCWWQWChLU1EOHhvp/smuXdYivwRNQEN
2KorsQm0YjbkJZKRTDrAMgF/RCpgq7kQpd1KYUPlpQMVYaIWzeNJd/Vw0EGK6pa7
Aju18h2SR/RxXk3J4VizDA5VaSJqq9C/m1Soq2Qpq6tOOuyujMc9NYniG0FFcV7u
Qt2pk40sA006Bbw9vyHyyGvJSIHnJRrpR/sjdss4X4W656+HfMMcgdNLB+PD2YkW
HmHLFFDLtTU1jkE9uvnA9GWPKVRRp5is4nkQ7BAlPBr4dbLbuVSy3LqxN3IPyN2P
t2iASXfGZ07UB4261sAanv/Bg1ceHI2VpfjkXVdfYZL8FXj1HoDOzW0WujKe5aa7
`protect END_PROTECTED
