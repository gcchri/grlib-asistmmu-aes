`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CeS+vbMyQ66q6hgcXGWiE0eASdnloZS6qW7NzC+teKqxj/EXDZU950s289/PMBH6
i7QZdsNdpo+nH44/Pjg/nZJ56YIxsO47HpUZowHltdQ2RPWME7S2UR90LAdogIT0
RBEGxdJ6MaI1e/EkFWA5IDAT26hyo2BDEcvtG+hr+WkyHmxwsLVNg/o0wEkKEVfC
JKvJKiIv97hQ6F3gKtNZY203sXC07tzPrxTcw07tk0acMGmcV9vXeee+u5XIomLU
O9jusbn4XrJWanTZIL+NZBYs2rNh42lUZDEEMsE57ZXDxYj5818CDVzsh3Xm8exV
TuYSLI0y3D09aDJfD/4K9vjZj85+lAvZNDakmkUlGVmYBzDBkPBhMjRClheQGGpA
bfFlntfLCGdC0U7S6RSiDWNpifnVZCBEEJ27hatkZQKjQgPca65c2tcDZFtzJWrh
R6LkrgF/rrLORCpYUQe2lNbpoeG/ETpThNIr/TSQ2Ak=
`protect END_PROTECTED
