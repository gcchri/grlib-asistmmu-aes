`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HmlOUG9kKqzYf80p4PdUrqQ91uKYA1+qxxRhHI6LGKBgtaVPuosk1hj93O/klkus
JXfRS6e936ffr3/zXib+VhX5HmJc3jMo+H8Tt6Ulkee9Cxbkj9g0bb6rWwEY+pmk
eQM6bvXCrsF0K6PtBYq5oKWt0DDjhArAt5J1tXDzkh6qbXEvfjB+JdbtuvZYsZEA
mhlZlJpFS++KfKtvGm6hFr/fVm4wSRwx7X65Hxcc9HOPyr77WmkvCGPlQHMSm1g/
9IriuNaso6HhKIrORRtiTsmbJ+IakJhlqRVHSnYlOQD1+BfzX0MwrYfJDskwzjkH
FxYkQuod5qlbB5YMOv+mwbrX3sKHKhlXNS4eZxkgdCLub3VzdTvuwtGBz7WBwMFC
uKZo8nU/jDfqPcttou2dmbwyigujgk2PUEHqHrOF2Bm3C6+PGupyzRZyWW/U5fZ9
O7Hf8UNrhQoxz19K/rFUkbV1kER2RvF9cSIKMGavdQivJIEUVYvJqtRYE4y/CCMU
8T6TZnwQuxqIJHcAQ4FjYn+Uk0a8fEWZfhyrW+1qeYsWPz5q71pUGQd07JQM0Reb
Aj1O7eIZUmzN3I6ebmLf7TERopaPLgvnSqUWYiE1hgqz5D2wung7qzQHYFiRj/cB
tHRNUF6fx9ppv3WBrNXg9OIabkm30Xsg+n6iaRj4ds5NPTVO8XHWNY3Cxrl6rCb3
Dw+dsm3+MyILCfcrbwuYIKgpcogcRmcDrZNhBMD34WAmvn1+IBF5VOrVPIbQYJ4Z
crNn8ZOMCERPKStPOJMAc9ctTf/n7Tz001xg3xqCYgT4F12zPL9gq6hZMi4zvKNU
Re8ziDv9IOr/cyJs8vTH4K07tq0MGadpiO5HX8jLlapffBbChdtemM148L8eZ3Cr
07yWUkb7fkRtWz5k7AEGgVZP3+2awTHUoLLTs9UXxMaNtqto8JXP5qB0XNxlpLGk
5Y3QHouRaCun2HSe6PXMkHgFYLdidC+fEV86cjGB0CmFeZQyTEjxBsl8FppXR1oY
tEF3OjTXKcuC5NsVoTPrARCAcNLyqrdTva30W9joGwoTAxbTrnZDVEslVh841kLQ
Do8hBCRiMSjZNTR3AgsYP4GTOCOQKgnaTdImvz1PGxGVgRHJT7nX2+SFMOPcyvTz
SY6hMU8hBh/E6P1q/EW/UC7c1PFaIeZ7YyuRv7pbfUg3XteY8vn7zo+eTkxLcX9X
pW7yiIhB34NF4NgQkpyOfOO9X6iY9E9a+2DqGKS2uo9d4aRXZ/eLMJiqA/3HB7Pz
6rzVl/iygCJux8ZZNj3rcT4EjKfcr3QL2SuSW+45eXiEDNwPVwniD4J85pNp7hT+
crfRxmlllQ7F7cTWu+e+1AObFk1ZmWUGhFwQLqUai0K3yy5FkLFU2/tggaZ6VfAK
XxHrh0/AsWftMI3gLWync4bXmqDT2XJuWh96e6RbwyVKX/XfjJHU8/7lzn4nJTWF
O/0R22grbuBg/+PgFNk5wWw63aj3sZqhFNpjVhkz3rZThvgpxr1dPAgIx7TXU4mW
nFcStgq9Pl1v7tAESUyuoXJuvMqPE13Bo6RohP7SX+CWu5WYviMkmGLz4kWWRI8g
reRCwqtlXa8o7OVbadC4Y8G2gWKMWNGF4bjK3zeEkl6MqirMJCfBjra/RAdWW//Z
sVCbdbqQolsk1c6qz0iDQ345LBJAmspPSxw6n+Y68ebNCJvusMoVBdewBau0cv3k
VNMW0W9TSOteVC1vIVxsH8T7HLzh9LgVH1zfNMXJCoox1l5M26pUEJI7NxAzj1TK
cMtwBtHEjAjahKLtaZ5CxxXhRk9i3gSWGB+B0mzsUmtVDhdNMlabB+5l/G9xSCdY
/6P9SjURsXkvRfIh9znTeRgZKKM151uoZkKyuewofj16GOX+LTSwyBetkV7nuBym
vBhNEM1w5jv8568h48sex8kgvg8QPnLI5+oZchw0tfWuvN6TaaRFsrtgFrlPFs+m
sNly8RW7kjwoEubqUanfIWTboPlfaL6ZPJseZobsD4c7nkcccSKLcmZy31mC4k3y
29g7bmskMksMYkNL7xkzHPQw+T5sAEcl7hLUvcLC8fM4OH2bEp/adVue8pCVUY5t
zUcx/i+T066ME0doC8FhbNGxp2V4MaJ+5newh1BDAzWUsRprsO8ygnytiF1lRHvk
`protect END_PROTECTED
