`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAdmbxq97dr8l2LGOTau7+LWyS88DtJxQNs3lvlVbISCeR0zl62A5w//8yJU1CRo
C8uKhXqp8snlm5C6A+JXMpzU5jiJz88W46F5lG7ywELDcf4+NQQzprvDAzQg7QPh
36sW7+fYBnT4Mdt4eaY8J0PkdeIy/Af+cYU+UztdKPeTNjdU0cdieveufJS2OEBY
dAo7/I9uHX3gV2MJRPNCGPS1109vu97ePG12TBtzarKnKzVHV85u11UVVHDpUsTX
eQtS+aN9YfkPfcVMDroYu4vZm7FHtuHNlJyq5yW5DNMqudV/O+rHNMxGtPdM3Ufx
jONGwMnFP3s2+bcVtN1SjY52Kzfd4bm4w6eiL8M5QYhL58oHuRWUMjdTzGgOhWyi
bpukIHS9RA9qFagcSF5rJyzvpo6C1wneQwMVR/wthVG4alU7DHDNdoQtwGuIpX4r
qAl6XI36u+fM6eb+/wQBVR7LXzlVluNxdrEyxEBKttjF1yiqlHSjzBChsmSxJg5h
1MXK5ZxkbTQtEEIQfnKvTBudINrVpvpKmBkvsq7xO3JqJf0F551HhFwLn6ENKPIY
8usHY2wVKvRbQ0TLz9QGH+t9L7FnYzl/MidAy399PpZlrbBnoroUr8YtGRdTzjG1
n43Ezo9Wwp/0r4iqaeM72bpHqx5amzFpcbdgxIc7qoX1FVjGA6Of2NUSvC0hc0rw
NZzZjJe/Y31ZhLvTrpvFiyNFswfCCWGjNzQqTACTLwARpuXr160YXsOh7BlSFQ49
GpxP5kxy6BxyYRgRm9Z8K+ok+c/PqzcE1sbD4JZic2hDsKcROW10xSXozXliU2CY
z+NM/yP8+ayIO9+4luNSB8vLPXFP6p7BY1FRQ44pgfrOfeWSWrbxDWpKmqsV4pur
vhtZ6tPF98kVq0gPE/9EfZGGSsKjo7Il0QgH1pwAGPBzxhQYlHsBySEet2OVxY58
OC9ROGDiwblk6rlNvkoPP8b0NcPhuOVQbhy/RD+Q5GfbyI7WBwLEWw9Q7qIZiddW
qv4pEp/ebd9eUrserKzxSsamkFd31wcHDnx9gt79/ocI5TQotjB+ZktdbQOenmAY
G7/QeY+lIBwAPMNXjWRKmaAn1llnh73jOzOQd9rRp72kw88O4Dn4vRqPYi3BB7l7
dhbGALKGZphFT3SxDIcG+1Hfr2wccgl8ayt4f+/APRbz9bDo0JeLs25rRDdyfLJQ
SjiYqzbwhV04Pu3ot3l09k1dNwpFozXw5pmht4KjYuiyCW1XY4bvoz9/ubaYIhc6
UL6aSLT1ogjWhMh00w906ugYHntdGvCarGrbrpB2+TnqGMRF9OPzviD8ZPqck9+s
ZUWCCjMcSU4vGNYaqvV4knamI3OkIrcNPKEqUPptUxYGcycQ/BcX5eb/2oSZPT8G
p4R9y3mCWV7hIBt23upJspadUZybxADZ3X/GaXMTPEU29KsBzahKjayTqGw+WqlU
mPVxuJ77nMufdilu3r2AqboFPiB33yzjMQ/lWAcgLzmERaLFbU6jUukE5oorTNKf
Qbu7ASGBqt6wHHcMfhEiwkd47Q+rpKAieKlIaThUTbSV/xLIXVQJIZj0KsPVYN4d
NhOYtUFoi2WrldSwUWkKYaWR0ZzDr6IU5aUCo450jC8gsjyfLzLsZVKyGeTemSuM
hs2Ji7/N6LXe12aRt8XknK1C+a5ENWbU2mET+48amRiJlEqNztIJNnNjQpt161GE
UMn9k7p6ntxIa4+sfyPQV6he09ap8XuluFOa6SEzJnPdEwZSd11r1hFBVv35Ui9m
SXaZh6fwPQbI7o79Ii9YdMIscQrSImA4E1KX/oS2kuZZ3mPWvfaoR3e7FpYg/5Vn
Ye2duWfXeBA3hxP09DrNXqH+4MUQOjBKNgnzDEqG79YYOiEYb9n5nl7NpmXCgl8o
EZ1pq/zloty3B0Jh6cWl2K1FZJ37GWYkGRR8y0KW1P2fq7c6avXdoly4rNibkspe
Ef2COn7OUPqRrd5GX9NvIJPg3lAy8XC9Yf1+Stkxe5TwgnxN5+1/tEVGOM6cDvkB
eALb/EDbmQMk9De5aKcG8mmqxHQTulDEQA4EmxZ2ja5GPn1x+donxLFadTmlwA0h
hq3VvaSe6fW9rzIQeO6HxqLVHKlDttoWSXA1RWHY3u30/iCudOwYEak0Gopbsg9K
zHxfUWAT4MbzV7bDqhKozdRH0lSIhFIGklpjgMY6urHzn8BZu9vA2e0WEFcF4YBN
KPZgItgdyGMFizPH8gCo6HJw0lAIT76/Yy60D1O49APGiOAfqj4AZsSA1XO24saw
9dsjCvHfc/LtiM1AR3R7XVcNit2SfpBRIeul7QMlbsQ3VBkad/uMpPHj9Rz3NoWA
+IwYl/MGghyT3lHjITlmyIapocu3j/YFJJYh8Ab9x9oj5fj3+3O1Cen+lfti0NJj
C4ETnbODIKd7EArzpmpwSMYW0AE4T4gVjm4FR46eaUxn9X8SN++LlEMqCm2lqhEz
GDnlImQYU11kNZqilpg5rMldmKjbMv96Yek/Dkgd8v9/cnTOLbv/JiV7D0KuDM58
dirG8XdlDV8aa4hsYfjTmI7kurakysp5wBgMeQxY/h0vGWAFLsgjpbnslLNvRyd8
ImxJ6VP+jeZ0hIE0bZMSauxaYy7xejymLvqfUR2O6B2t3KNvwH9vnch5uNlaIgjJ
SevXS5ys4bwfztgyrGXo7z4MkL94Baghee238XicKPxVi3pzYiSVrJkCzSha8Mi8
HSTZAE95FfwL+NKWi0leV+77aAj755Ru11+Aaf5PQpP+Fo+ia3oWrUFzkzcktS+p
jtuHKLp/mEZEsoQmlE3Tqdua/akOA2qHgg7GZKF/jHqo0QQMR503R/AlFXBsn06s
idQFjFNpMqJfaNrPzbHlPfB7hVpG2evFAq0kalZEOageMboqdKLiJBGic09XtOe8
cafhK+E/zG7vfNMAoByjY1ghpqzQX9Q+zqvxdUTgOxX2xHv6owZwznTIWsln1g+O
ciemx1M/g2Db6glTab0JmtuHT7058DCl0/MA34HpksnPAqtcJq/Fcf3B0WH93fkG
uT8sB1tK8F1Au3BQqkYWSmRZyyJBR2LUKnTryFrADhC8bY8Qfp0L7Fzb9pkDIMaJ
Ol7s9lA2i84ADew0H/8e/9xJMc1plRyEQGXJZtMGY+KuUFVw21Fj6HQs2mPAAj39
b4dfNoY6y4F5lTHFy94b2knHDHBA/kj8jSgIxhS0DmWAtxiZyygqsZughh+LUWfR
Jk+++22CA7Z9dxHSe9hgB4sAs64WjYpdGSq/AjJ9/r6cWoSsFVRcptJBYb9xoOzK
tpEVp1BN9ui1Qyaz6K8xcnHr5p7wvbeFFlxNrrgfrRjp4vYsBI+CUOT+NUea3LTy
cuQjx4WjLy2SYk8uIb0PCJSVtW1H5lGgOrD39SAN0GN3Dbs/opNcWA+gzFvAKFaP
0+lOgbn2HOtTy05mq2aTJ5a8R2kcTG2k5a9hubDLTw1RRShEk/NLjcDFWsuFRO73
pqxSDH3KnXZ09UJUnWFcxqdgFyXD0b6enNKPSBetNmvNOJJRd1HnyDfEm2/3SdLk
ZHw3LDuj8TJbsRLzpVZXdd1EJbKZ3AFxrHE/tu3Z/zcfCHSy7Cu5s8j6h5hH7ULu
pED9W+poHb4ghwtx1afNaoEoMVZ4MXEkAi2pXzSTKdvMK23MGf9gHJOI6nq0Pr5T
w0pBRikepEkLKb27lGzWqpf9TMmHzUhXcY2H/4I1ZvW381/Az/ZcGfsGdPwe52Oa
lnKuPsQr1EvvdZ0MXaqw0vCQQx8x4LTRh7w6JjUXrqFx1bxbGoYzA7TML9mAuDtJ
xXSyUqCm/lyRnedFtCv/Jt6lL/efx+a3Lupd6lNevM8SnqhLYpSpoXCSOYbLKECm
E2BgwWKlFA7CG1gQYoXOBYkA5ng3cByJf0KvqD5fkNOGNBXYbwDrOh+2Ehfq7sRB
6Noubi0F77vbMe1ggHCj3NiqDAG7sslhRdoF/1WZIhSKvdQAe6QQ9ly8gLS7CXfU
pC9qVOE+lDRMQgpj65c8b7iZ3+94IcB0f0pQKnSSt9m+D5VcOoCutONkj+kECO0M
P52VjQth6i+3ZEu3IHvBaRkatejiZ1mgB7eAjgfc172NjZ3KtH9q4HYUQe3sJml9
`protect END_PROTECTED
