`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kd6juA5u+nOl36Z3mG2tmm4lZsALQhw5GAJi6KUioSPHR2YyBf/yO1qhY5OAFr4m
4VbsApsmPh0RmhLw6FqSHQcy72+2/Ept9tRWejbgKGO6uVKK7tuDkMChJ34fS0HR
2sbo3AXlAc4EdcMEdglqT+sCe0pN/CeweUZ1Y3z9RyPdEHEA5olLqptJ7jVSdii0
ahmnj3mcMdioVVet9dr1wGY7CK8rZgo5qVEbpuj90odfnb0aoD8+7y7zWiobRM+y
zGFWHA2eq6W/1Jm1AX73goa/ecVBrJfALe0Zy3sr69wkNrcWOtZOeftiPv2KpXLc
fd3fdcqffh9CHiJhlkQUguui+XrHhfhq3IaEVJtXxhNcJi9606bdc0SsRV2N1sgT
dBLzhM8+EOuwzzOhLnJOuQ==
`protect END_PROTECTED
