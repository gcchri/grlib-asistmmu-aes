`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VJh7/RhwxJr2UguPEpN3/j1z+BaoNCEjpd4mJLyLVGeuEm5p0Koliz2A9FaQ1wO
PCT5QIxauJkMkI4D04bymkaFaB2Ve7ZDG03USIvgYEHwY4bW37OCR6S1U2hGo/j/
6ZlbDfcREtUXv/iWl940XS7LhZMXPQAMVrlbHxhATFllT9fY5TGEJqgZGlh1Z15/
WxSYGU01G2abAoTmwAGiIVEumHZUsHne8CjRa+X+IGNr2pqG9s5iYUiKxtnBRFgl
YNEHVwUgpT6VXGdSimOGkHSaghcEeM7rSsFyK8+bDVjZymrtHb+MeRyWi5luTzC5
zdwrvqJjXp1R4LNSPn2cT0PE86inwCdxak/fLvk7wf6ahC4josC7GoH7iEh89vHW
pUJsTGbbWTc6AH7dMxgUFtEYjXbHGPL1eXSlzLHHOhMAd1rIpQ1c3WM5CkYPTkMV
TILFUFbNc86fDcvkiAJpjTZXXAfMx67BYHinVRnD0STRgjlQ5LKAS23NpcBKQcyN
fptT9eCbR5deOOwjewlnQoNDiAU9c3W8Xzjw0O9VQGTcdqXBqtox6kmGdVyI0QLq
McwBi14bacONmxWgbSNDfYv7TDwH3ZkofIH3kMzO+U6qmBkVGdI4y2cp55bvyBV/
YNBUjUUf64po6hDtGxtcIzpb7j1PPrYG6yAs6W9V6n9KDKy8miK5VCqMyJQkREg8
xf180q6K6CFN8jw5jWC6UUBwU6ouZiSP+8apbwE2cXinvkf21wWuDI2lPyBv0EpK
WL2Z8T/yu/EfNHLLne5ZiWpsxI3JtsA0J8NdX/DUY5fUxajmI5rKPEmxisaHR9r/
DUU/0XNyulvorEVAb+DhwhvqQWthODfcjt5OWXcXh+8bw+bfPNrdAVA/dgCld0Ur
qPjgErF9sKXcgmvkCfuD43VtrKRC1EY68me3e3mVIBuETk5d3HtpibQnDjXvwIXv
+EV8lKMKWdRuVA53015TnC2zE0ScTwVR3o05X+ufiqc/1/of5QGlOMmTl0AFKqN0
unQdRVMccRblw18e6pYh0O3ZXnxvpn4DM+6FylGOc3cvDUuddRO02+7l7wyMwhCI
h8xXzJmPa1d2i3v8vHJl4o1q1FbdazeNh5oZVuuEjXeBRLGTrgpa74S5Y3LWthbs
E2RtdX+w4sg5UgOLKxQINjZAMtzFkuZrsm7k6tOJYUj5R07D2EqCzwFhY54iuLL/
Ud0+xagKEpONuUNkKrks0nNawJcZnnXC57cKT1o3pyVkKbNS2MMeFKTfnSZzJS5H
dmotBuNMsYMsyH6iBqmzYp28egNJqajIJ6fHo9qYfZD5eVEUpNtsb1yQ14ivRb+D
wQWAXDxxRa6RugAXx/wvSUlybXjrBsTFAvdv0X0vDVtqiPxgu9cJpMmRqyFCVdF1
oQLunQiu/weOT8zx138vFyXFFbjhiBPgDYP3cwo6ntQbYCrJk/eeHH6X0EC+0z8F
4+eUioo83DeKNsBuMaZ18hiHL4uVc4SA/ah1pW8S2jtwattQBoGHH8Mt5n6m2xdQ
TNHpGVN9ACedFGH6CwpnmgEfBa/rr1g4wK9jKmdXzYf/ENDmzinq3s8xxJSBv8pa
EpWT5W02ttPEdiDf1YPUUn6/BZp433oAc0xHrgYrb98MGDtnD8L3WId8uBr/SeiN
kFzy3jSF1iO4QT8iiRoERJ7h2q152LgtQrjsNta3q1oZjZdDJW5ai397R+b3piAd
8v+EGMX53ykVuR7/AMCFdkcH8AQ54q8kksX8wNbhzo+zC7E3D3fxD2oO/dioZx0y
njIploozosSa5qIBxCKb1L0qFznoR4g7RbBiqYsx8Pbdu/y6vFK2WMR0AuQQADNX
kwZantn/hfk2IdM7GmLGB0cTqkEfu+PAhbj0ecYN/z9puOZAZQdtLaC4rH+6S3pD
k7yisZUDTh4QWY0FWts5ZiCHq+qvj+aW1Tx10/Tn3ghqtrz+CK/JrOzAkEE+wlnO
W4bqK3totsXmoVBjGDgSEFC0lbVYw9x035Bv6sZmWp5fO3JNd6Ibd6vY2WaVW4O5
YsSILobjfrAdeZP+hIIC3IIeC0yF6FoeHZXzY0AsHg2xPqS3PY/RxG9CBzBxM9HV
q+pAXTwVZaB8kOCw1IJActsJSAXr5Vlf6lRDW3qRdwCwKMTPndVWUu6AHXMcMBGL
s99e8k+ZQ75B2i0TdMKS44R3LcQYdEO8EbanTBfJnRFJZ5s9XjI8x7o5xC23y91I
HGrSC9OeNIRmZDtF5tYI8d0LARKq9f7Opg11+FAh+nzV/mbdjxQsGY03fhHoFKWr
km3ls/iolXtUPtWCqU4u3haKCVPATba9MUGpZj1oWkVuWwYEoJcNRQhMQbUlZN0Z
rb7Zn5rLeofiNLx/t+NoGyj3WlebPMOsUyHCswIwpGuxDHKuTyXYPXDzhOdZkkHq
hOHfLnLovn4538p1aNs8v/v0VoAfuY6Ho0iqFQ+hVNaozYB6GGJI7Muh9NuQDwqx
x6q0GmbB+TDnkdSwJwclulYVpm7sgrLGOxZSUhs5khw5iLv4CjG4qIDuq6WH8TAV
EdWorcweSqYjbxYwHZU+lTZQHK9vocks/0EJLhHsDRy/4FU1sWnydvSi0NR53HzT
ZBslyyfZ3PtFee9kNSEKQREXeEh4bSPuGjv8R19hdGRyYPdnMnUflBiFJBYxOplF
YMyvTk82+cZDSBiJDXTqnu9edSbeVesHHMFOSrLEiqx5uQBCCYathsLlVlpjnl2K
0LlSadAyxFiVnPV99bWqIN76ESiygWRKEk1vw6ZSsg2XPwSDi8gAQhtllCl6C7ST
+UNw2O9uaNffcy9P0tQaXF7PoxeiVCajBI56eGfCn23rX0kFv7yV3jXUC70HPrb+
XjKMqtHG52ITGd4cZoXnBJLZC6ynxEDH3qd4V7wXpSY0GhKwIP7D5qY20fM+/3BF
OkOzsdq75v4/WsvLKNLSI1HIyj2wFUY9l1rHKkTRK4omzhQ5zftjmkV2N6HckSnu
JL9a07Bb33C/Jr0amX8wrFO6uQ2bq/Z80vd2TRpao/KEgC5AE+P4NVl9UEVK2Ybg
mpGI+FA67oXUM61z4XhZ6m+B3/+mvADJUSZlh3NJWIXoT2iADKtZnWgL90TNvR7B
LgCE3gepShW3w/E0DY1pfHCiHcWL+wMAQ1Hbg3cxk6O6VAp1eb9lz9lo5QBEmtIZ
TAO6nmOZ0QK0fThBRmpFdq6BZIfznSSC9BTT7n8eKdM6YdO2nSDmgDap3kf28M3K
JtCMLWKZajq9TsuPlzePQt3QsSKEsLg+sVjY+CWzxIIZSkFSoWBiI/zMXMyPLXfX
OYKd32KXOAmcJm47XW6pdVZvxJaZCTccsKwj8Y0Js6czBQ+wSUiyWtxeucajWezn
WQbPbfud1VEBmyAFOdZRzNL7Iy1CbKH3Y1xNbUj1vgFAmxtzX06s0D1/Uc1Hra20
8oqDLodhM0blZnhSxOWplrBsSXSmI+kH2jecI1q/m7tgIK9boG5Us3DlOUffDU/G
Keb/tim4/cGav+mHkle24ZJtLhejoFmOPxuA2fZUTXNMMx5G2u9ES903MpFECZPY
h+qAWZ9lBoK4RQsjKicunt1lwIp3ZUuad3Fz0I8sHYPAXRrsH0/MVPHDhCiC+tja
ytUm3Q7uAS8Jsq3C7qhdUNkpJ87ev/5RHnJecNVmHMEG2TcDJh3fc1xBKlGmnfXR
onAZ7bX0k72twanq1LiuOU1uZBBKBfQAtx5SuX5Y0G+X1lGsJD87OZvV1NCxbH9Y
pTugDNjg20hj0WAF3nOFGoMqZhp97uhgom8flMX8yBwBCInw5V+n5SPw+PxG5tn5
OAJiQMjbTowABpw0QcFvPA1YEK4dpcCiS2pgTdYBEWwFT/N3bmnR3RYqrcSLeCFl
ulkETXz/DLuCmvV9TEzZ/Emymipx2McchQcbtdF181swTJjC0u0ew5exZGZ2iLvb
C6IlK0wzHf2Wt61yRxo86nPk00WjW/wIBvJKwhKBLDlqa4JSGyrlkpqbPqSjDs5E
OfbyDAspyNG6aEDa3j4+Zv6j/8Gb8XpX7hzRTzKv9cIV3SX2JXw35smlzQrcdg5p
AcqOzqhY8ChkuFXqtiYBQ6J+SsJfHK0KLWBgZyFCMYX2WfdLsDrlzV8Ad08e1tHR
8ffxBvFBz2IZ9Al+KAChG8RUyfB3BKkus6iwdrGOnUbpwbGLu5rcbxEV33/T/73h
qDHI9e2/GbcQH63jOkKGRraLQrnTyqQ4gJi1c9DKzJby15EXGqGWDTU6CmHY7VAH
25VXLj/5NE0YXNufVCr+tR7k2n2G/uSGAb0k3Y2ec2Zc2Kexb1LP2d1QpRCqlbmy
dlJUEH0Qqqun6hySkNTYQewMaTIua5zcAUnfo8EhuVJUhbEEy+fOIHnwsbBD9SZh
6PhQ7m91lmf374kr+Cot4fOgkuAAIvUayJmglEsex2bW2SuLczVYpkvwbwjysDA0
iDLlU39hXPiz4eIUR7TcNCxAmqmgndJF88QAbt5tJ/e8oDB8TOwMARryG5GfoYU+
NIm72AxW2Z0upELdSjNyHPc1jl2IE9rj6gy9L8TAYap1/a4eINtUyY4DpC/en67A
TnSUM7XmqUcH/hSjPOhQ8MLUD570ttPB/mtySTD5xsj/TDJNyyuBuZneId4/4+wI
P9hnr0dTC93bJ3E4C8MgDD4yRf70XP0v/0A5+JS4f0HKpXrn+kcp0sdvfXatz0wm
kZyUg3vHmYGKbkBjBpjRuGufRVMmo0xyn+x8JAlcA0qGe+RvshI9qMOkT6KkWoEr
IyD6lmtEgR8LNI+xEuRUd4d8Yo/IyEJ4Nclimh2R4zTp74xuE40f1Zhs7LavgrsW
/EgCExVsv879WCfkOm1xbW3CkKRAwABkDWB96cU0qIn456esVhhpuI9VXBSY5EPE
iQ+Z9wja0Yb7BnrvqQWvyD0ACdpiZmmSiUruOHHu3fQg1zWvcOtDDlK9rCJRo2rS
HFT4ipUCNqfnDbHHZKYzKGXXht1+9r9RNFHcZUzdcLeeP7Ljy3336iVVuh7Jd/jP
Lv9Lsw4uae8b/PDiZAsNSWBNSMHeHTUjZunFOy7LTnEp/S8faiGtpNRP0vgo0D6A
OHPcwVxtajWYXcfmbFTimtoD/Ggk66rZnlOAWSUibWdvT6PO9WhyyZiNptdvH4rQ
VBDIlNgMTHpwy/9S9IPoMwQfouHhTxxm2//JD81e+NOcyLc/jN7oMrA+NNh9f5MK
9gDdnIluFQXvtKXawiE0Qq7yNJq6Tjvb+BYIrj/yYxpuzAdQPNMeIX6NDwhLBfI5
AF/8EgcF9KhLw2ZRMwyCKrs1PSqGD2ho2cVYAhemDkssTIMhubtlWSwWgmnal/wY
dCsh4RsafWea1ILfCdpTZ6SMAqXpZ+McCMO9dkGaaHHR4KMPA9MpnnkJHd6PzKFp
CNIjgPkY8huttxXMssOUZ0b/Lkc0csi+0A+FO5BmyKkSP3CMKv1sFUzlM2lC99Yn
QD3tYVRjEkgkRfXKktVB6DfxQ1pe5rHKgHe9prID+vraEiF4St9lTY6AHgkP4Czi
Ez6iQ4fNMUBevp/L3vTI+BZaDFRaLGke8hti5OKYMwBiPRTqKrzlOPocRE19GkAG
GplKfI88wKGFnxfLOeTnwGMTRVDHfPDt8S6fAOWZaKjf6CQsGevT0ricFzxfZpuX
aubcEpKtcsZ/9QaELk8YUW/ADI732LDQ5QP/S1VnXxd8PxqT6lCDIdaHZPCLem+w
88CryxWCOMMyzmGsKfFGlzav+FVx3L0fnB4cQMri33QUEIpz9a2nvVVDum6NZ5cm
0GsVtyPkeztHPqLLwqvBXmPCi2v75sSMXArA6CT7SWtMAjkJhWoOMiyJCFam/RfQ
iB1Tskhs+E+2ke60HcQnD4CPV5YTjB0Ey6YmlLQbfVej3O2rjiTCQgHJah0n5FA9
bXmjh9ixBMwrwIyhhcykGGXAAycqxElUQptDotf6sDSl/kUNpy3q4k3uQr3Qr7ci
8ynvYbzKfDUxaLh8xOC8+/9zMrAD0uakcHEqMDoVHXUQ1iWbrFAeDgLq16vSc8MT
KBe15Eka2DlFstYwn2RYY5Jd5ygKdqCF+CEPIEVm0drzCAPE4MRt31AXU7J/Mht3
jP1TN/9jW27aPTcVSjNZUoh/SzWRHgfN4YXryclNgh9+DO+Ybca9lWlxDg34HN7w
by/INbE/5UqmiLrJ08osw8hbACZdqMgYYCcxEr4YjpLCvvN4HmtvbWLOkMiSbYAi
Nwzl40Tcv3jGoW5W6XqMdA==
`protect END_PROTECTED
