`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DVIcaKArDb41y5kk5dObp8tiPDQ/d7Js8Ub7/UKKOdRBgvb+f6PxTeY7d+CeP6mn
Qp9wg6ArYJGAGAj/ab8R6SDsO03jJwFKRazr80Lqap8C//onTh4Fs4YN7FmtbA40
ZjbKZABq2M87Kp13Wl8k2O/15spgewFysvhLoLuzZ3BC64xTTUQdhluVxZqmaSeS
mGfFbL/dmsBCyxkf6hrv01/BvxzxMp6ez9qNRAbncrSpygKmYpivP3ospzKQFME9
6DWzSOEt3ImfG8A7dePMroBnfaA3wHifpJwimQDjSjY=
`protect END_PROTECTED
