`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O24KBu+Ep/BF30xpTrUBCJ3jEu3hbdrQc7QdOpImzsUOeXg+rHI+xPOqVMgj/pMX
XDgcgOTCxW1ItxjCvgQRqXOWFaEIFm8gq9bUU+egniDBrkzgu9IvDRmgW5V4tjLX
71ntxqtymMXrpHMaofP8lOsKzIXbC4M0j1claxPtBxk2gwlH/d9raw5iDLO7hHM5
CMirkLFz9YsHn2mmA9an4z47JdvHI4FghNoWqPMkP3QFDqSB7ix7dLQunOzN5Zyv
d7gzaMCEgxty/UuE5o3Re0L04oUWdfYGusWhmlYmTF/Gd1uPo97rrBKO72jPgxyy
0oxEFajvH5jNkaQCq0xhMmm1wuA4RCmYi/JkNhhcrt/vfozUiN+Fwjc0SmbHe6Dl
VxGW4ptiiJOoktbe/lkDwGSmLX3GKr3cIxAkmtGP/1lUn25OycgCU57uIXonc1ee
ecYlpyCyaCTnzChPSqYycPJ8p4OU+p5CuE3BCEgl/rexXmSTAmfy/YzJBZUOgLcZ
RrzwMgL+qw9uZ0YnmHXEQ/208gY+PHOQZHMN3bizJH0=
`protect END_PROTECTED
