`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PEmVN5n8snNtstTpDABYz3qj0m5RfhN1ro+eFedmOyKpihurPtXMuTYHfhvPV3QA
kkc/hZM86viXX7OkWYH/jPou5uQYVSBTRI+Ojl2MEZqlBNEs6SOsO5HQ4X2JkfOm
UC3JxYJDagaBWVqYl56RCIRwkfV3givID0flfyH6Lk0zfqCRfbkpKuLVFE4Kic0M
u0nASCpb0zAVeBc8rcMrnO8nDgVdH/HAMiHPb3r3UZgIh+9+kNs5vwHfEZboE6gb
7YLYGcD2/SMzfkRswtJmAX5i61dHlG3IYFUzDUbiefSwV2lvIbjYImiKzMKpbnFt
94sn9wg0pxCV3TUxukeoMjx7TKtUC4WPMKrgpOaXnJpeQMRN+7sUvh/9+3gNrdQw
vk41udbuIYsmcnIXk/C1D4fuZ6lAraDX/EEEkAfebnVBjy7mxfpRCILF3qzy1Abe
`protect END_PROTECTED
