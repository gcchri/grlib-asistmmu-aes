`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zvRjOqnHPwpINJVNbUoz/CBlhipPyWXcDv7phAyu6kns5Zs7VCfu7zXVb4hhgzgf
iDvCzi4xrXCrOYGwmX1p530pNGuVG1KC0a8FM4x1XT0lyChNLJT7HWh+LyyZYPRK
i7M6MpB2ohI+kFJD83eYtmfDtyx72R31wEDjqhcKaa9FmOMrvL1YGDgWjqdr+q0D
IMi7SA7GeC3qvqWrZGWEqc7kZz8npDWLPCVUe5TIBYYFuQfnXpqVqzT3lZ9QOgsR
eRX1w2bnjT/uWdHdNbLrBkTDVJY9y+BW4WdwqOsaEPETR3h+ME/7xslOq65lgYIc
x5Fxpf5Y4BV0CjP5v+qB/KnVY7P+Y6lJa8j6AotU+VrLc5VriR0+OrE+up4o6/1A
U+W5P1o/siIxV5HjB92Khg==
`protect END_PROTECTED
