`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W9o1oLLRNuO5+OxsHkv4ln64t+I6+tg/CQhVTpuQgWzIQE2IVbBKus4ZC/myDRjN
Gv3GpbYf0kU/B7zq30tWvSZvCmdPW/Xi/RZB76kwfftzpP8GHSm7Tn3xsyGzru6M
I3wEKfu2RFpfyui0R+C2TVHW+CsxGDb6Q1tNzNYnG+Iz1D/su6vqJmE7jqAkELF1
MT48pPoK5rAJ7aQiWW6Z9ZvLGU9G5cvSajPqSbDGCmerqm0P4gaU5RKoUxtXO3IB
z019XAwsoSI/VQEwWE3jAO/4CfKRsw0I4Qp2kPWigNwaSkpV1l81Enc4dGrX7Cue
3dxXjeiv/Pjpuk+rGe4aXiXjWZypgz6cFItyQ2FUbhBEKBSSkkdP2oRqvXr9xw9y
Auu4SQwIMOXvJO0z/1pn/Q==
`protect END_PROTECTED
