`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QE24d+4tblASBmH+C0wh5Gz4SMp2Rx1qSwZHYm7pzIZOF/Ps20axudW75I+ToTce
4IkapPSP8y00uh1HWGjm+A1a26v6ZrCREsu3t78rniYVxZLe/7Zka5bAekpQTC/2
cwqQQK2t4Qs5OgS9/JYVZLugRxz+XLSmGMpqabHcK+DUWnZSls5qFqgMpm4SqRyK
x3uiqBJlpwmkp/+X6rlX3n97/tBUH6hWK4OZ9hli8jAKn49hYahx0hTIiIAPBiSs
Fe7jQrTgHAxGVh4oDXCNZTFHMjJcFEsfvdwKcuKYf6Cm37Bke6hCCW659pXlI3ak
DsbE+mXnIKXk643HhBTbAX7j2L6ud8swNm/fJyNyxV1vUwLJFf7qbjqTytZhDRFQ
65IP2jXsGVtIaPQAHE3kk0uS+CL7hPJg3fF77CO2gB7aaRH8BxRGTO0ph4bkprsH
yBSQk9zqHB7tDpTMo8RQk9+MMMyw8il2amqxYTlSbzr7XSKWJbbtYVmpr1MBUT6h
QvZK++VfwyvAP4V8GTK5f7sxb6ZEk+NUjNH+qwt64AsEVGDSKPzSjNeNVRyEjNpl
0YII0Lg13Tq2QGu9vHMDDjTNe7gEiFme922+DFCrwKkMGDvUYjYf8E5s+6RTn3HK
a/0k4i5L52qO4Xy3LqbBjoA+W71PB/ycOgBScqxLV2S0ADibK4YQpeQpIrY4/tfF
rkbmX6yguHD5UYV6+D1GD0N1QXD7hVfwguzte7gyNp8UzKPohBUODJ3EzIsUTEdX
fXLU/MtmoHQscfH8NCKKWB5mZ/yi9ElsRX080BvygVomCLwPeHg3ETg1BIvLgIjA
Gb7oeU1ubs0LKRYkAq9M0zQrgKlMHzKWPbMymQh6l0PwXkP1SYsM5CO5gs7tTEVR
HNG2j6XflOyCvJmqAxy/RN/dSW9tetBKe0ri640o1b+Q8UL4U0ak3Vg3nou3Vz0D
lNZLy5fJv2xfxcccrGzRn0g+qC5WJAlIBOi+9ea5qZWgv1R+8CL0LR+bDhELdZ6v
V3qB5msn7U9+/Ksq1XOSrZTojVmGEha8+em3kBBJN3QHNImm6YEhiB9IzI34VT6q
UhdCM0CVq/WXtE39zDCX0nBDGWzEb9S/C+EE5EnLsKNHy7aZufUO/mhHA2RM6qdl
sPgUVB8RYNAxij+UZZhTh+5K/H9Ep15f4KBpTUHeHH25ZSHlBUuqUGfNJ6zYg/M2
Xa+hpnsxklOMqVSnYRGGsC25O2C0xbzq9O/dP1URc+ng2AdcJs8qY4hTHIKgzCGh
eaFvK8z5Hzyc9hoMcpuYUFUc+sPRJxzG/ov+FKI3b8cxNU2SY9zKv+VZm9tHxxJS
m1DCg2h1wsNFqpbvAKhaRFRFI/LqvzvFZYrK41rHmAS5hHbGFsMU6/Y3HxcAq0kJ
LgdEaKNnwGosxsFJTDuibVFZTRwufjhZ9khmgtDa/vK0P8c0MeyztitccEO8/EdK
ie4EZR6zaQs55fZgrmXGDZHamg2sHq2AIMy4lCQAlBIcc6XxouMkFHDuAdCo2tIQ
2cg5lPn4IcgUa2NGYfg/V4ho8AQ2E3OfGJHm4NOBdqGgXVYlGfigENSQhRnLOsPD
S9eyZzaGaswG9FXQlF5faKdJwajIuAaDw4HpzmrZHOc+vCkemzqTWoVDyXwY+5h+
RiitHZ0kPv3UZoGNtrQVZajbAU3QuoeSq/3sLuSptJxVLTVviJetzjCdLaN/7URK
lCIsWZqTdVi6/psxFpIe0qwuD08vg8pQufm1wf9xCpUaml4i5BneKMM9AFxk7s53
4RzuxyyWj8rgYyqo4V5MQZmNcZ9Ez4ZhosmE1wBf0otD5X3KfXLbp8RZKJrTyMaU
aIXMdDrT4ny5+xLZHlMdMDAHI/j9N6lzCgX0IUiz0X7rmIbCVwuFg/jMva04cBFf
w47HCyIdlaIHZJ5F1sryTLF7GT26MynfasZ5R16YAccE8K9JN3/qpCn5/wecJnEH
sYRDgMlKh1EalZ/yMi5cbMZJDzjnI6rLoGdNbeW2B0/kPLNlIVQprLIBsm67Cxt/
CQiO/jX4OrBnhxXmGDz2rukdcfcgh9phCG+Gf96j4mYHeISs9437r0GJKG9MHurx
wkvwkyRVV3y2Wb52TH9w7gGBB9iUPdmQsvbanxn66nDeadhsnfqNVy025cUuMunK
y0czTe//IMQi0SzL6A8LYFABGh1e5fiNu86msNaBGZwPSSapKsf/KReA9Olylwjx
bg3zQPzpuIvPBgSHKo3Ng7suJJpqfqU0NetOc5zidya4/Hk51GiKc9KFqGzO8qI3
zp5LzxcjyGhpVg4Zn9zVzUUdpdm6xmyj+Ocylw9Mt+ZVNH6BoY4b3F7fndOcRb8B
2HC5HF22ChlSDJ2HBtU1cWLbKvf0VJmXB6nEtYykFEQ=
`protect END_PROTECTED
