`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKWJD6DwWs2mroXhwWrMlTuCAjSifI4LLZuWPMwcQkr2iXpMXqh8Q5/Fw+DQ5yYi
OBOnN6R+fjbdR027V2vGypwfbFRF6oftWlv6GWnCcMnH/BEazqXmbVYvkGuewBAI
GnK/bAnRbEn1DSfnQqc62we4uvNfXwmZXNMD4JYDjvOifkS3A4cODGaVPbluJCm7
R8sMvKnU0e/ZaIT/lrSHumqDJkVdcw7qnyXQufe3nfOmTWx80H9n2qF7JCp+a31+
uyyOYPLQKxqE50IH4Ijlj+BH/nO/CwVRwYL08q2teTGC4YbKezXs57D7QGnipP2i
yZoMJGsZBRM27ayjozwsbdsty77mLs7aRCmOhGPt+SnrS44TK9zhBich6YvaJk1U
7TBT1g+ciVW19b3xW92wVdUr1cTNhVybRr6FBYaxNCKiXpXr37WrbdfnseAHTUBI
C03J6sj0+jfEUVBBnKk0TfDAarucVV/ZBcmjeHtb68R5G8pQWvulF42mSXyFrVGO
rt0e7XDzZyhvLRJizBBy3myOjLmIoD2iS6lvqhl6qsjtyfz/S/ht5fkV6PVT76Mz
77ln79+wfO4HV8oUrjLQOA==
`protect END_PROTECTED
