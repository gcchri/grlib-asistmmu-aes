`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OcdncrlRQGAvMHfAm0lU2+WpUz0Dq8uh0EvtE5EzK3qszNWt3lbPTiExz4nzFElX
qs+lA0cWoVQzfqmF/yS+3EXD8skykUzhRff9KwFRQOA9iLPkFDWVApafCOzYO/LS
e6lfw7uP2utW2PxDbmWsJVFMqcBYpNPm/HJoG4ZeDQh7BTv3KEwHxOYrjtYuCw/7
btsrO5ISewiHY63alXHzTo6G9S9cv8Ck0psVVZfAbc4NMFXpwJDssZS/jvmiq4ma
9qmsghUj5vFn8g3a4RAK3MD04G5QoLuE+SG21PpxD28xOO+LB4NnmECuI4VJp0fR
FNsdXJ9fI/k8LmGpqyOvrxaluWxSBOQNhJn30d3sX1/AGu2vTYkD4QKMdbmrF7fe
oM/Ny5zuJQUrsN771AeyI/fz6WhfYyQQDApAqre731aDLs/F/baCG1KYJpBWzQuo
kAvCwaNyZGpA8+lBZK7Vb6gLlt+gUA8X1KKi2qskrXTHYLJ9kAZt3JzSlb4VHj8q
qD5rsgupgpqTB+6iEkzvuhJ6gwLXafY//PLlF4TSBibdZdfGG/ueYa4utPkEcIL9
l6GyLfPtZVfy98mdLClL1uoPqnF2VVjUe81AMARr0y9VcRQR1f9eIujZTwejsOHh
s7lZv8o7vHIJZZDi3yDWYyFDBwSMJr1VgThmydIjfVWuYKr4q11Eeviwo1Rnvk1i
9he12OZDX4jejt4Ly/Dlxd40O4XPckuHEjMZxpAv8E0=
`protect END_PROTECTED
