`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9xBKsF2Q21q2offtAFvdMRMGFHnNkhVIKmxY1/Yf/EIT+9Sk8n2QvQZ0DJ8FZS/S
Wkdkc2+OH+9d4k0JhqBIfJhoc5k6WiaN8heE3W/uPeS8oiu9w6QLRwKD9X8eN2sd
obSxRh26mhHvl/aY2aA1Dqlm3XCVvONAlw1E3Keuza6r5OmKXAxvBAfTRm6DjyHl
fYpLqyGwOIhqIwnErmAqmjoYtj+BHNKxcHOIeAO+iZRKrHBlCjceiUcDOEbyMF8C
999AnfCzscz0cL10b/ljxH6oOZTHlLiv+a5efjuvTH26EYdNf2POi4yR0XDtbRH8
gPDbp9HgNzCCV02l3ID2Go5J0Y9nA+BdOSt18m8fegGO7p4flh5AZhw5p5iOO+Ly
pG2V1bWDaMycbDVvRrQV3CXOddtI0zPDe92M+Wa2dt1p/ntbZxw6dY9WK+vQf79Q
+b8yFq6ouSC+ZqmUPfe8kGupt2gGgjQzFfDjMXG8ELnMEVGsFBTG2YdOuDmABG2f
LJjIS7s/66XpKem1VcwL2wtx4ze1kum+cipbXyitbi//NURh6voCFpU8n56tFTmt
RKBzWY1SNY2MPsJBCg+f73gaGV2qPMbVLQEDlDiN7s9PiKpdtOhUXdIA4XV2V5fP
l+ccBI9vUWNuqvdF0gn5R7AlM5Q4glDaw1P2fQeTWzxMJz4khhYbnla3xyyhtgXU
`protect END_PROTECTED
