`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lNyc9LgCrqWFYEPRzt/6wW+0H/AOsFdpn7rziHku7n6BXKZZ7kFG8G1nyuOvYxJK
ya4tHtW0fOmDLRYlxBEOWL/zN5PxEMOayryfUQF27pS3z03BPREgCbaCPxtxQ3qB
o52fevSmG0DQRKr4O+1BM5naFTHrcTO3mN8M6xvzxuemYICWZUas7ubcISxFWC+O
G4l/IV3LdYXX2hYX/ipuqEd02j4lT9Wu+35JGE71n1orWkmdmxdiwFlYLY/JEdg5
o6yQCCuXeClfwTVIN2GhlqdGC6elKz9VHtv6TK+WqJSpJ8DBr6nFDMkxX1aziV+2
Ry3WsP+kmftCYk/2Z6AcodinupSpiDJaOstOOPUKDljzK/w1qF2EGaj8b8TAtCdB
rXdDW7/3AZ/VDq6In3nwU9GcmvLvepSvhl9aEQDYMyUq+eLZxbNdcHHCDcrKqjt3
wm153+dUCGF+PAQpcHhNZkYbU7aZ9M62qTGwun6BCgsd9Z/oxscAPU+8eLPG8qlM
bPc14QMq3KpHrWIiHx4AhgXyq5T5LqtuZyQiflEC+cJAP3uS1UXeNXqaY63Z87HP
S0hSNQLjvBvOPcjpvCnWmGCVfZt+W2Hj8O5yA4w4sGfOHroKZ1+SQe2TnmRk152y
Nhb8t7tW3L0uRid5cvoFiNCXN2fnbWTgTEi1mjEmvFjPYWlzBVQsum+IaDoIUzPH
aAnk8mhUfftnjk8HvU4SbDK8RahH6W6QNnzA0X++Pcbxaa1NePT7Se7SEs0hM1oT
aVwxTlmzyu43UanCHQ2Eo2LxQWjSaZf6HaOmfiXkJ24SCznUkCjiH9UDGR5P1+ZT
yBcMvQkVgEQTjOTF4IQUL6ApJeaJoMvf2TNnNnicV+6MT2LyaKmYooxUxZv3Cbqa
S/cr4OqR0lzRGpDAdR3nfMCFnk5XoZkwNPZg0trKGRSHDhFRMD6yQv7tOvhivNYL
0F4xHNHMjSQMSijj4GtDItKLE+eRgGyt7AYo8SjTxx8+WoDEXBjLo6/PzbCHLjzv
zG30V5sxsRXHWfpOLAEU0jQqXpVn7WC3VIXYRUMerb4=
`protect END_PROTECTED
