`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QfJkWAwVrhLQskmXhVeiQBdB9pbL0zEe+SYZcJjdfaIhrKWaRPG2CJ+ZYRIF2yJp
/8jKqNWqBhk84EAjbfKdwq2lXYRVzox+/DWOzX7M1Ud3zm7nccmxfZYSnmv03yWD
jXNrpAWe5q/6TcIY95JmgDOkImWPhyeE3Yiar+NKUGNR21LQ8SKidDy9YORnvPvE
z2Mk0BAvPO0SKazMSQFcuwpRpEvzzJoTg0IUjKps0jKoJxh6k29J0yz0UWtMdja7
ULMVN86jQJUu4ZOKSuzSYv5KtcOFYsI/j9y3mZQW/2vdSp5PyC/C/d+KA+8hv5FK
jrbpSSvNoATpjistvMdBMpyNhxui1JkhU/ZcRSqvR62aM8alZDMElswRlxbGqWOg
vTl1tsdGugmHZWrp9fg/rI2TbVxYISP7OSOc5MHdfJlFxEegFbRfFcgeFNe557sb
8LiccBTyp9tdE0SrxCLT67bHpIVwriSvFdIRGQrNbVXowAnvg2qGwmB/rJzsYONc
/Su7NqGlVOHZntJyHn+PkajtHbSFbwQn07a2K1s7t8YDsgW81014UsDat4gT5QrB
x51W+b42QCV8qkbz38XttJWLCmpHmeWiWppy2RDwT3dyn4+X2ffpVtE005TJbByd
iW4jA5JTxkJaP86bfmBC2ERnGswjVW1F+3iYgzXRwAjkT/zIoJBqyy4bFVbSR1Ez
QlMVH7jG4UiAthI0xu6bhLvEIGbnfo2m3wE728IQPUzH+ZAzjLzkO6bSUr7AHWPu
p8aR6Afj10+eCIsLlRpCAaGqlv46SNQvZIilQqy7VVjosMr9D/72D70w/PhkPmlP
vEU4i6B+ITWNJYCaMJI8sw5BGDs12bpZr5GSlJwA8Z7AJvZMHoLgA8P81DPsJJIb
lj/m3vwg5XLaBh4nNaW8L4RkXnjuGXpC0jdQ36rD0Xy+7jnkx2MoszRTYet3+WI5
7veiJZPM6bBBGdb+KfC/GvcEz/upU85mLnL9ZDpm7kMpn6BYyKpC1exJcs3AjuJQ
hc2J7Vq9xz6bCwM0bjifqR/6aoqe3TzF6TQD9EvYWn6fAfRupdXg0yr8kLED5/9y
3HCaKNADsKC2lx8/hiKGWmKtAI54ejYkpmKuyBSLnWKBuJ/8MSRmTAWjgafa2nGi
iVICrYghddg6dB5rytAqz+w9IfIlP0NlwzXvQK/xxJI9WKIqrc/YflOnEoTq6nLW
ERN6rf6gnxCLcesPJ2yhgjq8NTwfrvJV8PFvV4/DPZo5CK+gF8Tl6h7AErPyOm9D
Or2rsq4qeXFYufr7Zi6+7QqCYi9fB+AV6dnZJ2upIMAKevQi2KwGJSktZCSnc0bS
ia97ZQmAaT63m7LmvLok+nec5tFnFvW85e44rUb3Ak8sNvcyutOiUxa/zcUFcOh9
tqgdFc0KUfJOPKALxHqD4cBx/Lsy6gV+BrWVCOiZBnVW+uSbYqc/64bvbPyYTF6Z
QRbPir6wqb4pnRn2KF0FFf/Rnw4YP5g7zqyz1RwzxgH5/lwXT0PBwQ0vx+G9Bfgo
e/rC9xSZWBnvjp9cZ2Tj2lMozIEQADiul8lxwOPfYNmuZ7kZv+Hxb79/VUfl4pIs
Y0bZYNgDiyVzQun54zp/GZ2VfBrgIuDHij67w+h90O/LJ6p6fdvG9TF1MXXVz+3T
R+4tnjTD/G/cnYwvFMsenCve65Xk97Jm4NDRzk9sWgk2z1cp3ssVwzXn86cmdMKG
bTrgTFQjhxca8CGON/UqopZ+sFvIaI4QcwvIjXZynrgww9tSuRWaQMrKo53w71le
1T6HLn0dHrYbZjtLnLc+o55nFE7/0WQLvpB5WCr1rpBuPs/7CtNtvkKlEy7nPGMM
h6h7uClRx/Yd4mITjfPoyUb2Umw51BVrWv6BtCNjcP54larg/Fd0ULNB8slRkDzz
VCFsWBI6fSobEig8Dfhjut3n5VDIx1TFZhjCNFFH1faaGNc6te1Ckbo1E8Oby9WW
ugTihuBlUV7TV7MM5hPa80jPhx47gaMV5DtXmwBeMwkY1En3n/nDrrl0wRDifnz1
fRx8eOxCVyNLUSuFJVfw/fTYHI9ok7bQw+aPtQFspaRU5U/n9NiTnCBL5VQjFXHX
GF8sc5nKZQzxreVLStFwKA6yBNESR0qCGF9G5iZBLAvEEkFAnctuQHALR0NFwycN
WBO7MU6z9kNNRB56UHTUxeenLnyrOUef5zRYFIkm/kLFcdiUKQaqpYotEusRY4Cn
q8pse1643lKIvnlJ7Rv4bdTqE2xTl9W+L9khlQQN9s7SRg/vr0/4UAxwxzQsbapP
R/0aXLm+IZ96Lfsv7BsD5gQ9b71i7z6Nc1+XB06XAxM3TBS8vQdgSF9UoIM9ekW9
92PKKWHYWYTTJho7v7BwTuWGwMsBUljMG8WtlKmc1Vz7IZv8IMNlWyVWIW0IfeZb
RQheLvo62xPf1El13J8pXCpXAomBcKK+LNSi5/ZxGFRvS59tielyeZKEuOoWZ1K8
vrjOZ40ZVq6NAkFMkE9p+rbIZwqAE3n/ZkpFblgS5/4FEULJMmrcHUnDfD9bF5nJ
IWinRPnoxqb9gAIJ4NFAXN9MHqyFcTRAsx5BWX1McDyzU/I/aNw3F5LABYCqocmE
QDVPQSril0INls26Nkk5/vGk7RUUsDKQN8DhXSIGfdcYesZcpTxF3Lx/Hj0lpkgW
Uf6jXgx6dkNunpIXRoHj7lJQcWtvtSsH6y+StIBQk10bCTfC7qv0FNxap2P2bksg
PG15D7EravDnON2DLqNF9rxVhJDt0lLnMm7eYf8dENGWWGAKgKpcghvukrzrNg1B
ORf5jDaZ6x9U+9ZfZizsBNe58XVfzz2o7RCFEeT/YPcE1IdF89T6uQMZ391SAhJ5
08tFQbKKai0Nf5vKksosBF8S0a/M9sK+r4GpO6eh++XIwD60WeObiubg/qWyVpE/
o2h6N6B1sm2AeoglFmcOdtlzZyQcc5QxNbk/TtND+g2SpQe2EISEOvHPqQmQoO3X
KoU0bxNxlUqB0LX78W8GGxF6Lw2R+exxI26h5HGXeORIVmKxxBCcyp5uzF0smnnV
YWbVhFoc+5jCpnaOkHAIIRQdjSjFMLsHmif4Bqru8B13JiyJabVePArHxmxjV0Pr
6O1Ba0A6qJa+3W/63VvaPmazxEA3RCOxATK+qdALGtkgg3cqP8pND/Eh7786I+yt
LpYLqoxXzj3Fwa86liN81mFLlE18ucoeMsuIBIhnAVn0M9POBh1ZSn71lbpTO53o
DJCDmSySKckoCu4WsH6aCCmI0C1yf2OokKeWCx0zciprp94oUrHRWMTTzmW9jQX+
i7RgeQiDfFv3NPXSaDfUn1ZlmW+WT/ml8DMsUqdOOQ0mtgAMd9tMZu9p24bk9AH2
k0ETBmAdsxc0Dt1N9P/bKpXj9zIc1crr2td9oAR7BFw=
`protect END_PROTECTED
