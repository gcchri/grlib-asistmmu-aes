`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rGkFH4zkxD6VD1piJAzvwhlkRfuNshf6grJZlMp1S429YMVOfwCEHcSXFCgAgUJT
WHxGSoWZmIcmvG/rejMVZR6osXSLAx9o/+giEpCB0nxyRm0is15KsfCoL3GDD2PS
fe3i5RRdisXIpJnIVFRjhu+VjL0YimoV0KgGdb4fqNuE2FHCMdzbuyJ0+/mFIlVm
ULH88owIZCMP8ZvC8Itq5nhv5AeYRhEp1waCzgjEAxicJdDPtAJ8ivPppVAhE7Fu
t/nRFVqb5rmT61wqbR+7ySPKHxpOGpT25Iy54LHu4742QYgnc6X8xX7pWVun5Pdr
ItBawsWcEJie9NOYNYMqVyKhlAx3XQH5cAsklb9mCUIHoSUZl2+zvIOWkIyBTTW/
qCI3SwCzqXngrUtV70wDnZ8W7uH/LOMpWUNIQVtoy17Aqf/Vih181oLfJgZyC9qZ
YJTMQ4FGPWXh4P+FqDQMsobDBvtQgq7tcHZLpt42HDIaJaAey71wDFrtKZln0NK4
kGeXWCqKXx5Dkqv6J0UgE4/PMCuIPxpfzKhYZvdmQe/LIrbmGb8WKsdnUxmaOBNT
eJyXj1lsjMkHmtSAgcy4TqJ74DfVFPyggKem371Nqto9HycwDwx/DNtwEstF3BX/
RF9sQx4nPaqp6tQ+4domUgLxILtHPWBCVDXQ/YNf6FujtZPz+h8WLBBxTJD5mOxN
ArGYfNKgoBa1A0XDSmKhIttW9NcqVPyqwNyhzMLBHIQOiPLMDZdA8+P35diNEHFu
+VluDThf0eKHJK/kd/i8UfgSQYiZIpSoDfSsXSmXf54zv8fR27XpWpgwSd8rWg17
aNc2fTGeZVHRa0gXSprBH1o+hR59sz1ieZrwq2K/wQRlf2kgKTyjV+tQQ/5fXEy7
zDbqunEYPKsZJPesk+QGT8iZwX1wmc2vwQGmKt3jFM8=
`protect END_PROTECTED
