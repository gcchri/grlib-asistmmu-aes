`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RKNuKButn8eolR8+UpHgUiD6IO0DAgwn33rjv0mdehbX72kqjp3SLPIZKbQ2BCF2
mmoTqF98KmvW9tYulSc/djr4uzHN3ng+7vLci9+TbRraP4Pd0ulyLdsHdG8ybngJ
jFnM1vJ6CgGhuI+WpOB1NopukPvy+fMFAc5Conus0D/a5dmK2aC6QZMz7Ds7+niP
PD85jkhwB4Fs1vBTsfpAX/+c2lVABtB+IJrfsAFk8OdtRK4aVO3nn//4TUwwBXc6
Brt9Sn8qje7G2K/k+J4UBKekTtFdI2mnO6etVL41dwPUZHI7isBsc/GnKRqT68xV
VdzvQJArmc6f+YrlAUv5jiHnVE8k3HFB4k1WrR4G9Tl+YIYoJC8J3XAzkE/qT7pD
qKsWqrqI+6zEEiYZh+RYGJFV7T6EZJEx5SJJ3U73lcrRIQBVfhLKSKUgIL5+dmH6
0leo0I2Zle3acQ4pchs+vs/woJe9j3k1kLqEVN/qQ8yFPY0sBdC4YYfzj3GTjCeH
O4BcTBCTvrHIC8q/0e3On3pDE9bI5qsxC9MWTjEE9whfRbrcaM3dg6Ndsxcf8Ox8
c6UiEu8UQlQPYlv9zs+GUsus9yorY8q2NC9ZRUx722bFnlAHDlx573THD69XEgN0
5FByFF1QDsbq8zw6UNZqobP+CeoeTKRNXqqdiWKL9ywCpdvRVLNgC4j9ZSHTGmQ6
BzV6TgRK0zfp8IZnvMJn4o/KPG/XqhFulbV0e8mR+lueB21/r+QrH4glc65yLe5F
PeJPHOAy7aaJTTjv5tnDZeLh7q1cM6W2rKjk33F4ymGjfjJuOH2YcdBSvv6z+mYx
Z7x0utx1bk3cXsXiudd+IQrPJLb8lblGOCTT7WOSyEIPWZfUGf8e+TDJL2Bzd3C5
tk6AgbVDRTzCMH+84U/16doCvxjlWIwG+xZ8z7V3Wn2p2pWRwd6Z4a/lzLb+gjmA
PGvk1uSNLVvehvrNVAzEwBRozlZCZsRvA6zrjTVSsoJH533mf4zR8EKjaZaWFFkk
aCq2UB4MPKXYUt94eRDAdfJAN5sZaMi3wJ3HH88/fWU9xPp38xVK8+6XDwN/AJny
0uQahRQVb8zhgJFsAq2/wMcp42ZumDt7CQiBIZjzOMahmkH5HQbNRYo3T0MgBwyf
sUkI++kY4fedQLjMj6jr4XEIx5Itazm+ksxodjueUCNz43K1ZAsVocz7slVEQTek
KO8vPpUKkqbWI7S06Fv4qWxvXKuQ9d8uH/Vy+3oxlsdEDw7T4hrMew7A4o0JvDEP
32oRLRk3UDVoD9H+uCKfl6emxfL6PSKj52DxCSsMLaQUvfr3DqxQRhNc+wRO7ntn
Pwmh4C9qLM7G80JxBAWcqMmTs8ggOymnfRT71LI5vVouqwtgpOQ+2UQyf2VcEDk6
F26pmgyxCKtPARF3Px84fwB0UX1DKdVlyA5gVJAELzWA1zxKn0yoScf9B3Ptc6W9
oy0kBeZEvRhr18A1ao1zJgsCy0zleIoaxh2beLT5yHBoZF+MHvAxvChV3Ef3LejX
1V/viLZMWknICgNQ9IDyFuqwMfflYSHsw9QIwdGVqbJvKF7Zyz/toq7DAVllCViZ
4qDokjCC8fpWDoCt870S2mv9zuFQ6qHQowH9yApRHf7Hcqxa+GpT2qron/s9FVvr
y4bE6eR6FAEZ/q4YshptemFHXr82XrOgO/3ysi9q2RUHQkw+xB8ANmXinP317+gN
38LWxQ5hMiRCI6FSAcMBdXbIDB2ZReHwvU/IbXm6nH0vE1p+QGUCxOpGYHG+udlL
zf0g8UqkRBH8PK/rZbAN/KX3mZYfjv3dLIHcLelEio2H9R7o8jNt0Epxltfqjnsf
9dMix60K4d3X2BZcCUGA/NdkEGdxbuyeMX04u8/jNyRUhRkZDS5PrE9EqZJ/AoEN
9U6q4BAM2kJ1DfqQ5McT+p2fDVFnMT/taZOyPbl5mwhHX1npC63jpQPW+thGyjRu
QkTA/QF2mXwmZUjb1tJTmuAIKwYvMOeGFu6sq2eLj09KONV/jPdGAvkBrN6TUqJj
iamzezjhM3xa/j7Qd5KBMwSS7tYv0CtP0USSoLvr/evQAZOIOb5UlXCpi2IIZR7e
gNotZHKXRGI35LjNqG+qGz8tQAyiSX8jNRv9DMUkVveO8xvKe6grbPUxLX/f66Zb
XpEcwQcgQwwHA+QqVNB08QCcAfXPe3lVxEkcxk4XSdqjRhxCotro3/lZM1b8lH5M
Hz6GPdrUoeIbG4KVLzJxzJn+0bGhCBxrKBazeIg4MqPz1chOg+MRuwu6q+s9pkAS
jcAM/MNzCxowtRBGhlAxmcQRWL3AMrdgLW3tYXAOlfks5rlY948s9fpafssUusgP
AxH3vQOl8GBkM2I7srbgEg77f2g/ItTstdubRIijzMZdXaxj9tejTWrDciLP3aWi
D/u8ABPtgRtXwnxXxgPyfl37s3xHTUz+o7eVPC3fpso=
`protect END_PROTECTED
