`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAzsSWHlgdQFjKqXwm7t6MdJ8TRBUfCeTRtmMCg6gp/GjRc5QYalfkXR2uxq8ldY
yVwV1Nw1wWpnGYCIwsNXquNbwpoF+gAWwnvvmVeJmKkDNq2W5UiDJm0Q33kfAiZu
E9YZqHztdYpO1D7272/zHZiaHohUepYHZx/XBSbkSDzGiyXii05tmZ7s2doygWpU
W8kTzcQc3cWeVv6LlDTdhiZ1mQZSj4gI5VSC2JKekPXE6RauRqGTlfRrOVtwAGbc
lW2wr/p7RTH6t+cDhzIE2mphVOJe/bZW3trQseMD+ej/1mERsoSJ+hGjbLFKDKKy
hYKxcPKWgoGpNeky6Xb851RdRz7/3ufZ0ysJUUZd/BjWJP0kE7zhcqayifHC1YqF
9NxbmuP1zRUiv6TaS/xap18EruZQnQTepmPKD4jKeQzNyJwWe9a8zRsAYtFBZk8V
QC7z7OEr03vEANdcmBubEujqdllVjzxvpqAsnUclVVqBY3BCqKqntW2KXGJ8SS6z
`protect END_PROTECTED
