`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ciaI0O/HrTj6/bMBeF6H1/b5J0k58j4+6V7B+lP7oqpOgI6JtlXt7PjFwqUEddvc
4ecfcdXlH2uSbLOU8c0pf/Qg5nwA8MGi2/LJ/GWlrF9cAM9ghwp78rPKVR+PZjmH
CLunbjAnimbtbWic8hq6J7J51fGun7XKANgwvbfCSrwkdpLFWb/ivSa8gq/qy0B6
z+yQgK7TxeQzLoJOO72i/3yEyxIQKirUzY09HOUtzJ4BqrHaqK3IgTUJmnzLVlCm
MI+tB7nuVR4DUxNUCmzfVt6eUYon7Ebv2M/KabCLcnQvnbz5/DbdUZFa2Eq3PeZP
AbpP4anbCO/N6jK03i/EyS1UbpuGvbY1Sy3s0Vk7I6km25NcevLeEwLr1Ku63Eky
lZ4jiRws6yzddw4Gxk4aqjb1E0yKR0JnvPj9cwrRGnNJpv/55YMMfPf6Xq129ZYV
afTgGcwDgZZjJaQhFi8ZkG7lmegYXTiVI5TmNuCB+aYZpxGCotBm48Y+HqwADOrt
OKmD7UZvEfbyNpF2hCvEBy4bGZ3u3SakyGQMosBHPZMOjsicB3B8A6pkRjq+kQKC
o6qK8sEv3lw2evl8lkH8NinBK1b8t/YRGL2L1xyiKEQVMRKEAo1uK+VpB7cAja6Y
qgf7YDP2BcGTtOoJYDmnrMSb1bXoOjipzjlCVuUk+ReMO4ncNPAlQxH/MT8VLTCU
0I8xk35HNn89ZLTa9vi/5FILb8eclLHRR7qsxREIMMZ4M8e/y/pbIE6pqG2x83dm
xqApiGx3BmR5e3Pfce+J0u8+Ql2ZgHoq0mxgEzRKZfaj/BOYJOSWGd6UE+envRqi
7rK+J2Sqm9aZjXjuS5BYpzWz9b9RZ2d4SFSXhtoBjiH1WQj4/sM479LRtvK6hn94
tmNPSIpsR8Pk7cHgbpPp1g1kJQgATDxHL58fyCTMMOumFrI4yxFQ8YpeRGcWN5jc
TeutWiTOktoWhBqwWia9LBHjRVKfsVbIeItuiaCgdOBni48j/fx3eMnLIyF2Oocg
xvmPie4yVs6AfOIqV7nE/dW02M5fi56CxqnUR0HTmCRwtDuC5t73IWNWSxkdXP65
f9oX6n5aOV1guQRaurXWk3/sYXOubqi6a6MJwelUSNL0XxVwywHpmRGjTpHTazwy
yB6Qrqb29+qYHXSbrkGN11XKZaJzNpdv9coyBNPnf3MyZXovjByyBLlJ/murtInF
c5WZwPNW3XOm4fdsC/BVzqWFNl1n32fzv8ZuMbhFyfrhRTt4PinfApRyxUDvQJCQ
scj2SaenOQ4HwNBqfIlSclVijmsz/90mhd1lPifoWifwnwLq5HitrBT+8rcjclvE
ZBFA9M74r0oE+DyjuNkNM7lScii+0+MC0Lekxss1+ic3rN4s+iynU1iuLAFsvqO1
+GiXMI1TjWUTT/eo/0MFFsjCL1N+xzqWI++ueETqZUrwQxxrIqfWOcX6Kmd6i04n
p6JbJM5+tJMngvY3KhsiWMrlvvUvOQzbY5efJjpF8lvFPt6SBvSbIK7MscdnM68I
Md8mYrR62S0HqwV1IjEYv5TpUlDw+o2RZhcphKCAX89KmO+QYZd7wzXI7SKiKtl4
vcC6yQYolwmvNyh9MJvZgVKb3tQNVUpOmFXK28kj9hW2KUIavX3afROxclmlcREH
olywGZHkRh8wQr704aiuvA==
`protect END_PROTECTED
