`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kuGNYc3FOEh03fH6QLwNsKkik4Ds0/Y8gkeZ/OB+PYZz4YpmKqWxwMSPWXY36mQ+
v04J//OfUD6sC/1F3HvQ2NDgw/hgnoojv4QaLhCctkHrjHhmsF8bJaPtrMBrehU7
O5tv1zDmFba3sVfpoHPCgupDTPILapwdbhN27yh4qXy4loLoBDnQ+72fduB1j8ot
d0hb4zcMLbgnadFQtmqdkUgIxGl+bLQnQCcEQ44RDltrc03h4COwCNVdvhyO0KS6
W1/LSWm8VC+htUKhO+x/PWhS7gCigk7CntzJk+sUqmtl4M/tssM4h24TDt6ZCAKS
5sRaW07/sKbixVJJR4isU7BLIn6VnNKsT1Xmb69BZ34Wm1a6wt4tP8FJDVcsM5sD
klo1Ga0fX0DleHaZ8YdmuO3xhC+86CtPYjX9Z8beuE9Rzh2ByPp54IbFylOiVZbz
`protect END_PROTECTED
