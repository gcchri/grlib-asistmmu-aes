`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yeV2G+swtyp0Kq/Zbb+8OpXS9ELYDm5a6l4RruFD6UV84GsLgv+ugYD9zuTwt3hM
vqJpQYP06Oc83EvYFoWmarangF10nb/Qv9fcwCWplf3MBt1S2/rWAIc4q7RgaA/e
Ba0ijxIYTBLwbSwM3N2arvcPJgBppG4u8LnBrKpHIuWqpDZB/5Ock4/x06uGPvYZ
ZYy5YbjZ/TPTf4fDvosxFTWtpI6vMDJVEoWIDr9Nf1eCxUiy0RvVnd+98qkETcul
+c9IrZZ6QBnPhxbmz04ohZxrHCgujWTGR3Cl/aXAgOGLtVbqItV3Wt0TMueQUsyT
VxnGF5q3XHE6LBexEsNO8A==
`protect END_PROTECTED
