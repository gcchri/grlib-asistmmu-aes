`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+K/VXRubCqsUFOHBt0KOn4do7wcsVS8Tr0Yic7KIl7wh2C9DaDxSg2m1QrMFux84
yQox0ntxdawuMqftyo2y7h/Fq87+d6dmCZsjZXZLdVdSBcMAWikF5ZRmIxBoQtZ1
T9UMoyReJsRFEf0TDUWdouJAfm4ZYfURIftH1MfkjILWfwHTJn3aKwx99+f5AaIh
g6NUgP1JZOCS/EOdZO64BHwn6hEWS7cKj0DJFgelc9/Lo18sU4R0kyU4f1hZ2dro
D5cpfPgZsUKClKjyDhMPKR04U+bAemGx1QtCDFG5d6Z+5JSkoZh+A6boSLzy52dI
q7H+uIpodOR2RY72ihtCixOfL7yHVEUNH4L6UdmCtK2NWdl60qnQYjFoKvLWk34V
DiUViBD/epztw2Ngx1CftA4LzYgvTK0CTsnmisOpz7omHGd5Y1HsHeIwfntzAQPY
w3BySkNrW41VQAfNhIv3mVHZ1rgg5nCuRQ5NtMAHsA8wZk4B1QzPijDeRcH9iaWd
nkxlGumCHwOOGSZsRKtv/ArKH+9PCJqLG9PYqhn/NgCpEMZI5JE6qyP0FmdQgdgd
g+0PHqaHQRyxsAW+BqTB0F2erB4R3Td20E2FiVNb7s67AUi7ZE3UQXerdc4e9ukD
YhcX+kuBC37Yw5uUxIOl1qfCedGHSbypjaCuxT65bzw9iBgEU9wOQ+JlbbwnGqKd
oQGiQ0TAutu+kO0oI7Gf2mOYBB8q2d7URTnpb99tIUNB4QXYCssl/1zrVo4mRzgp
FJ/pchPzb9TQ0Ata13PfLhEQn5iBJnhZAOP7syf73i2jMnsrrOGUnFOGGuoVkIuY
`protect END_PROTECTED
