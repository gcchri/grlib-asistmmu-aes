`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dW0H/6Z6XlunjPn6PMVA45SwpgPx4yFh/TKd2QNh0lApw7H/QMs9XZq0o/1bv/qG
O7nNTJPApa4iIxCAATgdPx9jDkcRNkA0GxxqKUHAraTpgqHu4y13xXRUaNYfxQHA
cAC+TSRVWcqp/OaWtdOJ6Miv8qgu2ylRAMAE1pq+lT2qAGAIvgVj2FMtqcye+qix
gnSQTcCtMwnw4qmCLD960LfsxIUvrBYq3nPWVM+GsidlTdh31YKn+HkPsd80zbM1
Hnn0G87E6cdHlgcnm2Y05mmPFz7OK08tTR3pn7uZJKzCgKgKczn9u4nNkpX6RQI2
s6Sj1tS3+sooMMQUew/kE/DgMrvwvGZUcGQQSWRHucm41iBWpziBF8nk7Ellael9
4d/ciIyOkvI9MbGytAKXUsVCqjrTSN4S/6NKcNGFVDxSaK894CMGk0NxeNkcylWT
JlvYuliVKziXjYEzPGYe79X5ysqVkmVo/HoU44DbQh9nYa6ONVQGhu6h+gWVEsSP
`protect END_PROTECTED
