`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+9y1JDp4Q5cpYT4xR9pupw9swihqRSsG/bmcg2Llv2SgejHBc0HQTo7GVFUBXjf
JaDHPn9T+hGWX6luIbOKZwQ8noPq165LLNCys1qoE6tGWDYy2nr7304ZlD88kLUm
ZD/do1M3mSUne+7VSSfWZmikz56utpvgNR5enh80UHPgaYDGrCD2ht6UiaGCxumI
weo2gfXQ2NF8bAvpYJt5HDXqQNdygC3ldyP0uhyQJxAIXg0HLCgB3e7rirLx0yh7
suz2KVacUk0iKaBrj4Ja6WD1cqGkO2h1OLFfyiGTVgEZfuRYq6zaBBhmhEAtRwhn
pbyQAGOMK325ESarpUZz/RF5dVPr7SbU3tNXsZJW5G80hLvIxc7yghJm7RRjO0TJ
I9n0Fo3j/417D6OO6oePeUJJmAlHcpfgNTfal4UcH69SIa9MH9OsQ/4IXQWdVH00
`protect END_PROTECTED
