`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jdBqyRqoLxcAvzEX0L++7mTCIu8NcnKMaCgYiJ6s/k2KaU9677DOPMylDphxoD/D
ELtGmQM6uSDeEknGttwusKwennkwtBSWVhny0qe9NG0cyCdhk140tXww4IDRSMX/
/Jsc655pvABOitE98DX8yhPjokRHBMtPQPVHQXFpBA0mCFe/BGR3eEuRTvyOQhmt
gQpIlRjS5Ed0L1SbjlseZOWeJHyvsEByJOw7nh6AueN/YajgU5sEIjfIFTHDBXdH
OP4gMPOYNyza8c3OHkoXua6yx2YUQC0iKzkaq2AR0uPG5pjaygG2liqAD2sihHNx
M+3DJOajpqQQ0RUEpuAvBQyw5f/yafiqbuIrBiUy+OVTZnACvv6yV2vzygYrHMvO
JnDWszWKdLl6qpD1DNZn6A==
`protect END_PROTECTED
