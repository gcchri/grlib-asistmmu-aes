`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8QYEtMTxwPMkyrXsgvZk1ibd3Hg9KMRr5t2wfX3KN/pH8ESQNxnX8ToeU3dvosn+
W0rfGdraj6sGMfLsk8jGXo+Xd26AOKKGFtf/MpNYwP1lyFqk3uL1Dl1Il1c/VA4t
GYavcTYFskrVMMBdOOetmDmhlnhR/iq0VtYejH2PWqRDKRQUCHx4fj8sBQg/nuLk
HBJWEYXtVr8+gp5Xzyx0OSYvBmROI4bXjzIG+IVKZxv28oNLuu7LDYpJSxheRY8T
E8PmPkEbFo5KPNW/M6Epi/Q3rLD6yqrJPogaueWgaqQW0IP/ThqfSgZnHAw2JUNb
WYnD5BhYbz5Wb7rIU44SYcPiK/YRJ9BJpCZfa9qBVBX62N+2We6HoR9vVNyjmaEj
YmwBHvuPoonG/LW3LSn4rv0AwaLrDLE/mP3coAWedmbwTKs+fxfUGKFqHNLFnecs
8RWKRgv0UNMxcwn8one27Uc5Jh5hzghdua4J9NarHVR9MGH9SDDxMkGlp8QrB3Pt
kaz4OkiTN+6UDmfYBIZe28w1/bs+b6Zw3BjYlbdqP1aGC7JynLPe+B9mpfteTTRC
OTbvzBJ6b+AwwGc5B6UAPjTWRfl9XwPsn4oz5Ce7pBZFKzpwsx0zV7v5ZgtF38rT
U3PXV0x1eOoDs21lGj+lvfM1W8jVpONEzq6+WvfczfpYAzu1s/MmtN5JK3gzdULV
X9kbuDzTBK6eBYjCi/PEvQ==
`protect END_PROTECTED
