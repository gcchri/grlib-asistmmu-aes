`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqapVN6TGDcXQtQn7KXSsMd/Yp3QKYaEfQy8/aSBEgh2GtaHQsloedz7GZclUBl2
CMFA4MRD6BdD8qmzQytMAfEe0LbcLLOiVRpN1y0NOib3T/xgk2gFya6Ld9Hvz5XW
jGbnluNzkmwLO6uo96Y4ncUDV0xWC5xXRmIy1nxzI+0QCEYkq91hdlmj8W2t3z64
Sw2ACL8jv2eJY2Kr3eU5HwszFNCN3XRxV4hVNteHSeSJ7HE9nN62M6B7N3d5qkTp
4n1tblsOcVAf94gmCzh7SZ39YnHh4aK8zc09eixZ4rRg+t5EnchIGwMXGrzFV2IO
KvN0GPFOc/Vv63rz075EeBtbwUwvpE90ID7JRUb603Ugwdr9CPlOGabY1hkSv/pB
gl/+MdtBRrN8mieL2IH7zFUhel00LmKXy1u41JHFA5j2tAb5iWvgvrUuu3xtXhnP
0j+yZHXxIs6gXdFANJRFV5vMCFHL49N7UmF5Jp026/1ZJ0RYzT0tOmCXvM3zD7QJ
lW0OSVDtN7YoJFRb8ih4XyBJkzUpec71czKYHAOIKpmSDWJIVqjvTsWYHPWJt+w5
`protect END_PROTECTED
