`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yKP3wolBCCOusbbW8wiVN2PkVMx0hi/30T6hVdNh8wl1jKoWBNe8hhPc3FUzs0Bh
PIKP6zt2aJT8475i7hhEgMFTu2i9oNPzhRdXiTxtcFH+UZpdA+Zbwf1WemupdB50
bO9ZaBHHKvH+ezLytrTpmoBGKofCuW2Tq7hkNK6xACpAillm7F9njQB746kgKREL
Z4sgHGatv5hcg7q5sdiCrJGneM9Gy7F3ryttGh0F4BVrFlZGLcCh1rtFqy8S7N9E
D6WAgJsmkg05aDz0ko0HSSKYWYSA/Pey+2GACD5WMFHx/Xvn80HOlhNT3Gkar9yV
DdxYs9sA8SMCKc1Nvc/NJ7T0vcUg+XGmQX+HrTDOLvZUXL4kszcMwyMbmz4MzQCO
FlB3u9o+BTzDCooDhSrR9HPifTjDp9yoovsR379Vpg+Gza0jH/qT2O3Q98n1YNc2
ihjUmt8n0ED0RVA5ijP9ZOXA7tk1Fs1hZTwTNytQ3rgaOHQnmrkO+X+Gg3Nle3Zd
pqsXwieJTajJA3ObiCuGGn9l0fZ760PGzV6Hk+MSi/7yxfxVU5Ihtaiiz3k37U2j
tWKxKleIuq/FBhcQP3ZvLfjBZ44kPMFZjIJQ7tzOgyLRWD4il7CxQOcKCyaCvxDf
PsLNG7ngwyRQzBhQ6kuKog==
`protect END_PROTECTED
