`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jvy935M5Zls6/L3KqQPeKROCIex393iCr87uuTUh2vZ/lj78YRcAh5cmg3KoNgCx
MPQplhEeIPxFxl3WPbn+zdcFct5W1sOl4eDcwrO+KT+mt634DZBiDr2NRifJ34Oy
YUpGNRLalG06Sa8oE001JzUEpSKH4ZONQcBq+VZ/Ocq+ADQeuB/nhOLGpnvBKYY1
0pLt/eHEqofkBAX6gv976qCo1vSg4ow85SmTBE6RUsLJUs+DWfyTi2tA7SufQNJ/
jweKi2iwR4X7z2sD1rz160ry0Cci9/hgzhSCaCSmFs68s+D1hKqKXvfF3YjHgLao
+vyOJFUD5Y03VBa4FJp4mEX+gZ9WXgs9RaLwJf9MEq6DZU5VFKycJtRpFvEmtABj
bNVgpea+RJUBezALcv1EZSSaLt3+2BrRo+5ykqnHC/jOtMpSZcUbKGfl40QaGDAq
pk9rUpVi9rW1Y7Anp9jK12BewPZ6CUhbl3Q2rCJe9049PbA4F5K1u58feuGnxQq5
sNkNghWZgm0hYHwGrjiU/FpmhMT0UMCrm7RZM5DgA4PfYHhjTprM7W6eV16gFL0L
2xWlduzGPXgoqUPUsIG+rxAL0tsT6ph2NBVK21+N54A3HXyB5l/eE08KMTnzV3XZ
h+Dmh2czl1COczOpAwYAKsEC++tegHs7tiMm2G8e6euL8kvOT8BcLnYp7HNQDE8e
De6hnHqEIXBGu1H3abmIIo8+Y1Afp6C03CbqCBA7+E60ahBfvMa45xLcKHGki0hO
bCrKdWFqH38Qx7p0ATYxHqbbl2lwGygDSuu8QmPCDVGiTL0XRmqk1zHdh8nu0hDW
d0R5IWZU7rDr7bG3vpTSzdsxFP2TvJg5qy4SdM1Y/46P4ZDPmTx5Py+SaTgOIr5U
dxMQ3Tm7TNSNfmGBCYhlfOKefw/8a17YWZkljglw34+48+crFErMU9ufj6g1tSO8
a31msT0pGO4sooAbOMfc7iiyMvZ/3I2KB1bKmuFJ/n6kG4plHVN/q6u7StEvYSXC
L9mUfHAJAcCF0Ec2pEqECO8wU2DVfae3W/TakxOmPNrB7uTT2TA76Dugo1iXiljm
sGIPiTa+scXT07wUsMDY8+/Bkp5/cttRoxTy6w/HcjUZJEFN/FyYfqLkWnnHA48D
hErSwkgUrhD5PpVYU20xquGqkwNtdGoQc20G7pw4VfqNQmON7ZrF4PzDRa98Gsur
905V5dl10+qdhY5znCIQXwRjQcj/bgufL0lHz0RZuN2e/Ma+3tLQAeXxznQeI4n4
31M8INDwV/TuLgZ19Lu5RzAy+fkruDsbhFtz1Pnk+QIf4YntYSPa0qyVJZxJwMlK
C6K6BE+qeCXokwXg8itojrVD/Q3Itb9VscLpOR3SOJEfkCH3uckirlyy7zWnpDWz
tLqDk8p6lljELoFj5UorbTetFh8Y+hT5JLil1BBBJypbr7eoXBzzYl9QvU1dDgSA
8uhd1vQkPFu10arH31V9iz+biasBus/O4GvyekjS+/wG4uUIPmbqR5BiivyzIuPP
LzWLKaWnvaBSHgh8DqN+wOngpx9I9VlkyvwrjOWO9/hBikSQ3MShdTEOyQmD1GKx
Pc+XR2uAHh7VKtidjZOUmm5hHSG8VJ0z6T5PEz1dOke5+UU39jyLMJlQVwkAEx1g
XdW/vYgbMoDcaMbh5rUDXyAU0ByX52ZIJdJ5yHwA7vIEiOstsmdDRmmxJJR1k3KU
brD301CnDAhK6DZp8DYNI6ABJBHevWyfM6CbsRl5801P0hy8AVZVX6bAzudgHPSd
P7+yd4Nwi9NiGBWTMxfygES8P2nGEr3eP61IY0u+5gAG9pJuAS0hkc3aC70hnvY9
KRXa+/pjyfCaxXGjKerXWRj2zM126iL152xCsvo7HesI84xaNV3KF4RazF2Rjffq
W/JC17+Gow/VOE7inJJmVSmnF9s6AiTmDrPqDLMqtWsW6PLLPuf2JS8/FJpz5gJq
MT2FHwRlWoRJA1bh0ZIewiIqLyJ9akqncA6mgXa0KtTcpTghz7CAbuxsL2025LmC
NN5QHok57etmfxfAGw1s6/z2NgFSs0dV+B4nlAL5sJL0GxDM+hc+RlYuUaLM2dgE
R1jV4NBzTvcUQ3WNb58ub+1jad6ZBCTHD+UdZ6tm7VlKYg4dUEFdsOetPIuyjvw+
CLnJ1qUjOO1gOFjq9dp4ieR0MyF4v90F4zo52ko33ujBi5NW0D9fUmH+hlIkcaW5
JNuhMAKfypsvoHZhOx0mt/4uZFrGhCsOBbg2iTM1acGZMKW3ujI6A4Tt9n9e9CTq
MFo44JbrPAJMMu6A4PcIGwXeKeuZqMtdTo33FIZOi0xzVZxTgm1A5kqCPBNDEaON
SRZCNf63dtG5TALm7hu3HWsZW2f6nRKjjzLW1JV+5U4BNU7PtNzOj5lg/tF66gDh
Uoa3tLlUbvwtPPixc93TdivE2w9eadC40u9dMZc2/Xp7R71NrO2tJj41yvaQ0nmz
NDnpwI1tcqMKTUOmmgK4874hz+Nc0JMvwy6+eNaXIoLlv2E5Wvc25EHjzRs9euSw
7CME6cEv1hoS1UUm4jpr8Glm6fkT9XdCwrQI7u3AhN9GpJMvQUNls9OQaFB+JJCa
H4lRBpCx3ZZFznzSICLRrYo1mZwt+1jBfUL+L9r6MGSxG3Zk4MHYzt1T8FTSHk4X
L7bIe2ISYHQSjMmIlo5Z/vBCsjTnBPjsZefC7Hyb8M9mpaqyGkInFFo22Kc3Y3EG
4LMnrcM2kqwQVvqRkYQ5ggoUymugYpSqqbEabcv0csgmjU/fed49cVP304dgLzmy
vDhE6RKU+uzBt1N6a4gXel8o60GOTjJYp8Sc2BGdaQhGWm1HbyAMjI1vfanG1uDi
+9UKaItBlPFDLyP0ryBtz9vPHja2MIxIUEa7msC9FLma8xJCZmvnFMoBut8PJuJ5
C6iOemssXxhxpyaiYFOpuetIn3A6sgbYK56qYnvVfRaTwPshcGGfWQAaD17gU7WH
h46JZThMwg6/Ez9zs1KoYLHbhFo9BBPLqu0tM3NCnKNb4kS1U3v0hJuomObStqFM
yMGl4nQT37ukQR+7MngFY6y/JU2vnDf42z3SXVX6MPaHxVtWilQNm38jKgFlomZb
u+S7hs+3ji/EHWp2vOw0HQdCHb5jMi/TX7WNSACGQrTuDku8azmOKmEuXhfLpKpV
ympstYfS+G9tp+/hr5vTU7/qZFXpT7U+fa3uBblhkW0bwvixqhK8wcLDJRVmetvx
AyjRxcjfOw6ywiH7UCmwKDpgc4KgwJMC6t6Nh5EMxAbgvY6/eMC4tcO1CvSDcfvQ
0QuVEjKwjI/F7+1HOIkpDgRdVy0Isq4SIVJh75WgJdKstem3NBjDt3yESbaX1h/s
OBx4wOTaU6S0L//NjgfRm/BJTUBv5g4sntfCvp90t1jpPhTXbkUvYvh4ozDWciQP
upQkeCutnhlnMgo/NI1fMDcFW15lPQ/j+l10RQYcyCYF+hVornVLjp/wopcunCzF
zjE9VPMJjtGrKYNi8HcEi5G8ZUXGEZRxgpjjh0/yKvE10l63kNlfTLt6XFFIiyep
cC2oii/HAtGg7hJpHQoquhghIDH6EY4RYATlehQXNF2gGLKbnJHJjzlcW7qQWiqv
kKTPrXrG1nCrxdF4tvA3c6gtXuwaBPOTSkNSxj5IaWEtKtRb76PZhxZzRaQizQ4A
LxniL4ATMFKjAVfZQc7+qzTJy8kd7G//PbFH/jaE11dHgH6iDgF63amp75FVvd/V
vuvBi2W9Djg1g5ox618Fbh7OI0S5Q0aumU7sJ3hUZOnYL2BJlADCD4QM2cz2+g3e
Cotgx15wCYlChAPWVH/7DrMmZVUuliqKl0eu4zQO685ZoI7BEOKP0ez6OdzdhJou
xO++Nbf4mqSCUlEL2e7vWd31d5KpuMeOv2O9+aLebdrUC5WUidP3GyNZvuttVq3k
xxj/xNf7psn4h91kttpwcewYH2Wqm3Nz6do9eNWTIviY/eww9zP72tYSzc6v63Hu
4p5rsl0YS8cMNPwaeYS4s/JIVWlbgNMbUDNRwe4GLevkq2RDhXX5xyrjoJRtHPm7
TaWgHhc7HvJji64MXqS0z0g2t5DKm5P2JrnQAVNncIY2k04/kpQCzSIsAZzsmETv
a7Og36DT4FM4WXU3Ka+1Hbc4mH949vI5t/WTrTCv95/K12XtNRKWPDz26GnTqo58
II8WlzIt+bSeoO42/UCRTHcgZb8VySRk1IZotBcwr1bAg87x9KIx2NnKWUW0NQgp
EJWH0tohKOSu0GKAE+wjPrdp4Q/3OwSF3GT5PoSYy3wK2E0YItKreFp4R3YkKd57
CGVMIGIy+lrZqgm65Gf4pn1LZPPgE6Vr2oEB5o+7TVSyyO78b5NbYTVmK+Q5ctDD
sFGG+Pa7SFxtCMPshD2P8VSwvuFjRLbWTyt5QFetAwusP1VGmyC87dsfm6Qx96Yd
6bHE94noTE5smvW4h5KiIOO/YgMt1iuhsHNyrAWnv1wI3oi65tOA8MC1oHbkWV8L
ixR0NM8cz6VFKus6M+Ngp2gzg8RDlkg0iYNv7+Ct9AdneN2rWK0wk0i473ZnXHBz
y6pNq4AQZh2/k8XJkqDItRDUHxFdI6TcqZlnpTlNsOnOL+SmQj4eZUwzKuQnv1F9
uAY2tXtrKfPdPDhopnueybqabpsyUqiw1u0/9zouir4by+un23xiZxEwmLhpiwJ+
rz5X8kz0a9hSRsUFotbCojc0iq1Mn1NjtxPNjp01TY3cqwt2Ofu49jeVvdVztxYO
9BJu2WB0UjfiC9b0qcGgY+BFMY2Wm0+nBETBUv+MaGuUJQvUZsF4TubrBqDlLedB
MwB60hfgC1IC4SIS8U/xD2zVgJj8tdCy1RH0b7xqvBGnKoPPNVJ8Yz38tY24cWSc
83NCOZg7CP6Rv5sJAoo9xTjDBF/oShTyE9+ueVe/RCmWonO3a6rh9pQoz/ng4u8Q
Jt14lseDtmY/Qn2q7opqgInMynLEX0QjuCjv6bSWRo6y9CQjdZLxYAvGtKgYoD81
/PjtmUL0JhfxcWZHUX0d3CmBEHmm/RABGMHOiEBHND0n0TZXMsL3BwDt6PfcQBPF
SaGB4SVdr7YkADp5ycpCQ/pOmbYgD2tgUqCwoYZH/2CFdKzbhFuDoyychtpzf73N
REVjVzk3Zlna+mZQrGBqnkGHwIxYuT5IR5tVycXk0xckU7mrVFyyzvrCNB7/E7UF
9a+50hFVr0sfg0ed+34vEpnww55jRCCedA5glgopZCH2NbpzY9lA0fgzvjugP3dH
lJSROFNrf7fcN+m+vHrEHjrg5ud7mTDFq2iXqPQt472j+dDL4zdVKwLahelZYKjx
/zcp6+jg2vrSPnDHQAknxEHjYb+ouim74jFgXVmsIOs354aBE6rDEeI0/xBQ02sq
wro9Mc2jkRzOXvwVXjBYZ527coFt/PbQDJLYTetTtAtRNtUS8u4e5zQcqZ3mn/zy
yi6tHW/xhCyGOvzKhs+GSukejjTZ8JqZ+qUJKiq+IeXMcgl/2mfnjnTluQ19gF49
gRTEMsWbIPTwUPt48fjk7dXhzi03zXosiHQMS4Wku4NcEUoFJwxaaX6wOZFluO0H
CLj/BQ0nmVTpvb1z5oS93H1EIsil2IUqqB220TjWOBx9cG04uQwYji5cTJiI12DW
+JFL3gZmJ+wFRWr51O7w6ssIv3kspvWvmzctrSbOyILy46DHyzv/T4CoKgZNwAnH
Qwaa42/qKQ5BPdAju4wvU54aDkqQ/yDQ4Sh9SRAN7rwAGpzjwA5IWs9Wkp50GA6X
ytlhMkDccqjn1Ad8jrSTePddUtqeE1wlahkqXPfmfIKcWMw2yy6Z7uN97fpnDeNi
tNJzHLpZo6jc1xkGopEoFX3OkwJIsWwO7ORXo5paQBhUgu13UKvVkeXiDKijo5kH
eHzHdHZd4Kzt5jkRVckpeySlnzh20GlFIyCmbZIegj6nbhzbRzWdagb/r5Xfv121
sODJ7e9yJQtTLlOjzxN9AIuOWbkLU8/SxITIYTXe/suItFZsO6T9KYkrHgNMjyGm
9bcem0rgRJ6zkjg69lQcdCiisFwaMYIHYimuEUqA627CgY8sWaeS7V8IQ40fsQq5
aSrKJiVYMecLe8CvxgSDIjxpNNhqG691aNPzKojZhi3FBNUPWMAS2o36Yg4mXbhD
MPADDGqs9Ugto1XNWx1EPjuK1hkzg+epuU691IcLWrmHk8JT6j6H9b6QyuTMu6no
n56jta98yyxuuzHRRfJr3FsteBi6lKZ+kae5yYXtV+xYwypO0ve7Vo6k6K/449M5
HOzfL1m+Lk9Vp8Gackya7zUxgJ5WJG25Pmqg7U/LNAeYl7H5vwrwhIL8R5j520Ac
sxFo/kPZhgrP3zeaQwFx16qKtYTZ9GpaBZqlHRMLMFDZCcUJWbzGWIKa0LQHst5h
bnfzwSrJQPjE3UbX6xYG+J8GUu8Nh093o+6rmPRq/eE0ibgu0atHV6y3mTWb2nMC
NBC4xmZUUilClNrrwh7mjODGLo/FhzO0s254JqE4YH52iWHoH0wc3P4qoqZ8o4oy
NNLtuluiaJqcOwWLkpG5r9NwPAZ8FaqpxNYPr7hFzbOlbdLSDmJMNMlXh7ZE9sM7
WOQCc0YUEfzVLXAP5Ysrx8r9aGju3LDL/2gO1VK2ma9gGEalbjHymFNM1pQcJas0
upU1eWAO7Se94y/+dpbMpnqQEHd09BjQY1NThfUDxr6QwbpCHEUEN+OZC3fggHqT
BhMjUtoJprlxnrGRdHQ+9musBl9QZAtVRa37rkkokI0ehVFFc7lvdzJJd5NlvzTw
0t9idZT7KfuyP9zrUPOpIsQYfllPR07W8TXEulh7UnbsIffyyNNLlFewo0mjHD/d
0NpYPMuVsmNKjpyBV7W33oMgo+IkNqn+E5gatqRx1CihTzuVnh2fSOFH3s32goBz
MnEa+mVheYxF/msgSmbwjpC5kTubnv1VEEonwPk+2M0YCMPf/q7MbZe4KjXIWgca
dg+VeoKnLPHIFIHmG31dNX9+LO2wKxql1+ALaIv7mf5QK2gGXCj69Q/uQ/f1xb18
ZrERkkE9LaHENzyjCFhBOeLtVIliCTWLj8c5vHBPwFSBGuDsVQjkFiOPWtI9JgGZ
DPH+p+IV/+2zlMtuE7CyWW8BU9zFLzMbkdedluSx/vUqunZU389E/LHwA3OR6x0/
uTR0w3bFbiBxOHWQdaEAHw==
`protect END_PROTECTED
