`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSWOZyw9PZGBHC0A/Jpfpy5oOy4O8BHX723GyWU8g29T4ukzHQS+1cT9+8klQSYu
RrIi4uusMiRyduvZ0uo5W2Pj/m32BuGH3synteTzdIjQ4RxADWbcbB9B+2tVRMlF
6nDJfGNcSwQXBnonDApb/om3nWb2DhR54DYKZlP72PeV2WwAebXkPs5JxtmFmnod
V0gHxgaNXJFel+iDcVT0BZnrbDX5xlBiVYGRxfKO3GTsl7T6cQFIdyeRNg9Lomgg
WCDATt/JLNhT4Sul/xyw4X3JwtDZxrUisnr2BYxQ6dOjQwKAZ8DjSRpqmqbx4xCJ
Qe9+R2W0BsY4dDQOLnVEaw82t+F7dXNApXdQh7HcEA4bsUQnsXaCyvIpfx1s77Co
+sqUed+n1eRxW63/IfkzmSnF+Le6r+EQwjtxXJa9rhAV0DqRyYIdGhsmKegcNF8w
D4/dh1BzHr24NKHG++4L0d2YOAfOr06vaInYZmiF3jcXaHLPFjvfiwLhThoF1wfk
R+9d8l2Igrp9jbR7JC0XP5keIyMJ2H5zeQQ9IhIuif79gtiB8kASkt/XZzrv4CHT
G3Z11Ae37UDQ6ejX9YtS0SDSFUUPB6Ln9QPL5vRp/6wK8wkBXuE9LFL9BbMljBVj
44IKf/ahs6tw5LEOhQvvXayPRNk16d8S3oW4tBRifArARHFUa+vg8DKgS8jbhv6r
wnnzEoBEQ7ndq8Z6ONDx7msTF8KZh2WHymB7XP6Qg4Gr0QcvFD3yQJe7uBaJEomp
RKL8YagQdjKykmkdD9LPSdckJgv3tAfZAfX4MXl5mWqlJL4qIAS7RaqzzFvzmjHd
KZO8k9qNW7T2jXudOJaEBqw7OZ3FTu36BKD3VPZOxDg1EmoAg+Kt+K9FDAd6v3iv
eaNzXDEXg7Twpf5zrNQuI2EGtPVzAK2bgmQwdRAZJ4i3hBzBZxZ4muizBjGd/VsT
5iampVcvoydIaa9InX5+7hNt1Ac++6/UHCF2y1PceZ3TCzhDBOg0i8Fc58K+9bM8
I/6A/OY+hiq7hAvc+cmxL2FtTMxcwqTTDu6Ktx+YlKX6Z76snp56P+0Nn5IGWwbv
XXTGUFXXxVWZXZdv1ysrUWtWaxz8ktVQmQBBfKWPzKrb2TZA7oD+leMNYCoWZwrG
98FvLJThzEdtgUIe3z693gvz6me8fNRgfBaDgX9u6kK7kTPz4nGD4EdeiBYn4N5t
fSI37t9pNd08v9FF9YuywJPSvIKPpCUHwUISy0D4DxS2NtHrJ0CuxZkA4QbVXL0s
ByDQHTzm6FgsC0t+IFvtzjEp7rOYvltAmfs6cP5Ab4X27kw2ZfDMvjmOj6MKeBL7
rLIRrhUbnx4wwDOfpcFIHvmwqC03a5nKBHUx337/8mAifI4XDOmGPIDyPrsi6Tgl
KdB2ypOdK2enL1XiFN5OaUhK6IR0P1RjuDVcdWYpM0fmXDQ4xS835orGfFs6suox
hMRYLPFl/mQvgi4axnrjCsB0NScPZ3cFWb5oCqy+i+peWnF6VHEWV+MG0iiFrTWa
wZ8KtI+qQ21T/SWoJn7xGQSFNz6l6lFMUuaZPvkEyOk60wt5fcx+CoxIvY6lymjC
Pxrkp0SYF+XcYpkAAr3KGcLEpekGUo9dRhINsmEMQOveitP0WIjhq0a14hztZck9
eYmtQg8sA1kBr2kEHBd9hVP6bzIC1IyMAlJ2iT3PZkRy924Pi7Y/TdXjaFMoCtz1
0eVlGN6Fnj/LQr4ti7LA+I9DngJAX5Z3jC1BWEvpvTjSy7kl5YdafVXnYKy6xNVC
gT3LHzNJocpbI95A+psVgidyPUg97iet5mhZ6Q+E5INHiHK/j8xXtmygLEWN/7Nt
lA6YSX4mQJ3qr32hOvzBfqbBFsTU5w/MoKlfML9TZEJrJuUkw1DmulpXmfiqvqkK
R0fenBrNFj+AKUoXUu9wV7mbdBSbUJ0g10Bqm//eNrhQ0+221Hg/5iW4qj/4JzNW
eNt1tJ4vUEbuHEzd0CyVBXg93f9ISFqn2DmTC21L+axPl8in3vmYIM+rSjBnzZVQ
HcxzI3krwu4Y5ZWCuQmhBHWEZdbqK8AB5GufGu7D7ga2U5c/3gZP/0TyA0jCT89v
q5YlgG+Agd7UiRhwV2jwgZYIcYRVLAjcn2EGApBxGKT6OjM0ZYlTpJXY+s0d29vB
7DgBfYVm9BmeYtmoVPrmN0gQX/efnhjKDoyND6KbaTxnJgj1BVfw408qXP+mnata
Zze/BPK53QJUk0GXVdh/DA==
`protect END_PROTECTED
