`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgWDxozrsXBvFLgUU39fG0gksK+ibyQOKuskjtZUem4W1l0Wv4YTkFEABNI/RwMo
OEEo157dst91IhiRJw4oWK7eVNEFLkysAi1wru8yQ5nbRtIIxRYOtvTnKAjIH7/h
2bolnCLzB93kyR9zT6Mf0YXpGtevz35vAEhwy8ctE2DBdobMYwrAgTDPqvLybw+K
LSLa0dxUm02nPYyWJiXT+BR86tpuvX6rA88tGMnL13GgbsihDxgQKeV41IOcfg0K
2sbjcgvAnQUuLJC89smUJPz8mqRW478tB2WwG9RgpwlYIDek2O5y3oPYqb9PwYbu
F7+flAy/r9rQtWq7JMhE1n1XpW9gEmJuKOzNBT5xI++Ndgjs1+2Og6nXOWqRRbuK
OXHOSHp9cBfW/C5j4UIHL21jC7vO5INuDYTFQCoe5ZtfWjERj4HJa1iXvbyDQq3v
wsKLCcRfRxDKDoycgzn1PA==
`protect END_PROTECTED
