`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ntya7v8bEvm3pGDzVPvIWY/no2yCuSJjER4qKxJfirsMArKxtBUmHwMprMS96N2k
c2/7v20rby5owk+U+3qKeyRYADJVHIKD3LkbunoOv5qOzgQ6FxPJW9ELKEYag+MZ
bxhA7c4mLAV0vanBJTJIcQ82q46fd23saKDpLfhdu96iFFIqZkyZor4Zh0GyKzbV
C/mP5fkCgBv3n+kMtL0OzctUeahjFv4B9FkODTzNlNf7VUf1pv2lohVdx1Awio7X
wcEms9myRWfaTnNd/DUAbKyQ7fwm04HehtSlR8ndkRtQHAFYArPyWzo7Ebb0JAoX
EkcOFEOSsidYPoQ2JMHDAWsUUsW7eiDnPqbKSTQ7+0lBgEsuR53Te0wG3IpecDdN
ZCUtc6YVtMBUL+t27uDI6/rqtKykf0lECdQqZgBBvqPc+rXwvP2UCK2/PFzFPDfr
jgK48rsrs8P3PpORlTBBqu69slpvG7Uv+QVSM9zveGJYyhfr5+9jVadKeo4nqw2o
`protect END_PROTECTED
