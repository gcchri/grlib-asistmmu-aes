`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOGauqcxtzwTuTAbFXzm1I488wKGnGOzCE4kEy3iYKsJfMkBnQnVQIyT8GRMSD3H
cd0ZD/zKh0hDXsAef8Zcm587zqUk/cXjOLvBIgOVLFYtRwkLRCHoXD7aayxvi0vj
gO2sj4jDnEey8YPFSq69YBy2yUq394b25CscTL4tGbSqf1AHpDUupHKS4F1Wqs2x
PmDnZzei4kDP79rN1zxCO2n5mux/Qcx0nPsYhT3JQFIgViJNgzq6FKP3z6V+qUzM
H93WkTHAziqaSgfsLDmE4pcIRSYpn+iFxZfyfSqkHFsZAQ8n5+cSuLf/SJf2qqRg
Wnifk1acQNj82/9Pk8DMT8dv0FcbEFUwD7dEzieiJhJjCo+CRNWXrr/C0xb5Xl+b
rtUKQU8WJOu2K8zuvOc+4g==
`protect END_PROTECTED
