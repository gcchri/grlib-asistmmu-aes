`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QA0L4rg/Ix5tVEaYBuTBDdvnxfdBNDmu94u/5laDASoLXylxARaqcat5d2oUpZW
o6FzhugE/4QpriLaRGA2ou1jD+UxoP3pdbxZquT88AW3Gwrs1waDBTonYJ6A4mo6
5oaYIEJDJ++fHQ+aeFSF4iu4IUJBAfkF/rjmcvkhPQYXd38+fioB1GUTVkCj104f
E159X1xbBV7ZjvBS+chCvShUoGwhctFWzXx/AiGuY8bfqzLVS4rS8h6acn87tXgd
Wa9FPWt5frAcw/Hpz+HUymMXfCHnvsLuzn8Du4Wf4OFy7vKgtZnpWPXChk/ZKQLU
C16VdWcG/aP/sVe5E3oQS8ywgwSiL6U1Tg8YInsPGPpiUHpeZcjn5wpx/zUpMOal
J/mbBdP9qXtvcY/OVC6rEgPLX8SlR2U0pgJTWnaWNHo5mbdCQxPjL606eUVu1UlF
/Ge1FrvHNTZmvqqDLzPc0Xhj4z0NrIWWToteRyW9mCSgJMl10/1ewMmH+T357WVv
xhFZt9ItTZ2Ye9LVwa1040joO11rdSuIYKuhSzzifqBWVdKYGyIYJtQZ3h5otMP7
5/ng3gdwnFcr4To/QJox6S1+SIojoHONIAI+oZQWutSGibG3sv1P22ZOnM3kM3JN
iLvVkQTDbT6VRdHDLhmRfHHwexfBn6r6Trrazj7tNliVw8XmP1kMsbnchml0ZuLe
AyQ6FS+aFYkDN7puSGnD6PAGmWD/lzMvteelaxDxUlE=
`protect END_PROTECTED
