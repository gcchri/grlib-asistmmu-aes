`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/Y/+pLPBRPaX3sDeUDVtdqRHPN0aI+rSlbKdFs/ahN7atQaAomuX5Ze2ckEJ5Lc
YG1RlmI2sHUIXzvVXiS7zH9fFVpbT1tlh5rJxecNrtp5rGUHDzqgFF6dleO5+8OB
CyHw99hocUSvPDsYhPWqJ5IgNoGug6yse4FD72DdVkNN1JMZ/zfM4rpQSNnGu9mG
fP/RjRUSgjUu++pT/gpriA==
`protect END_PROTECTED
