`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sY8lRmqvQHSjOwDrlj2u0r121bg+kPVg9WklRMuRkr4KBFzhUfb0iiqyeSpRIWjM
f3mPyRV+SgVwE6VUgFWpGzIcRyO1xpdgEPPkdcMoQKdpDg9nx17qRkLj+GeaRcPn
B1fps9CxmwbAJCVZ5Vcpb0pCFpy0jQYIyhi3K9HphEPIOdBVsvzDj5+X/TIeMn9C
XEu+0I6UNXcltJmjbZCmRjY4d9m/enukJmcFNV1uVrTBF139bx5csVRauZ4uUaj9
X6y+D/M3ceV+47ygJSIJ7AZRqA2YoPkfnDsQ7sCkWIM=
`protect END_PROTECTED
