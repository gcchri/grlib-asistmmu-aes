`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vUvjXe4ulNhQ+ziJ7JyndiuhpI6dT0F9Z0uDsH7YB7WwWTvMARQUQKB8gb3Dk2qj
MFJGjNhP9011yJQ5ljrzo4Er6h1fLV14iYXWo1AszA8nVEPxZYNyWFjzllzQdtSB
ppaoI/3hv+Q4qU/MvZeJzk7DkS9E1Xh1yaeM2HtswvRYl2LPIJNDT26/1qVS3nw3
An8Xfo/3CQv0/LISVl3ns/ABaPeKUDfzyt7Vx9JpXP+W5WGb3naF1O4CVAMOunH6
GqsTgaq29YPldYKOBCikS5HBate88evTy4fkKh7y1TfAJtl4jI9+LiZkh01Xd3rt
e6UfFWt9wX9eoqbMy105cbqPE2yEUmfvlU9QqQIZkoemS/uG/a2PQGmbRpBv/qxS
SkRpmZTbpULAx6WhPzPteU4O16zWMvsN9DOcNEScu7C9vXwZc4A9hlTL75VPbIKv
pCeO9zF4+Rx3dSRcB4wi43Bbx45M6CflRmyKVgyKqVAkCny/pShVwvnleA7Dv/VA
xOFSOvEr6m3i1PHcBWYKRs3l0i9l37ruy/T6W9f/UBUyNDpQcipO+QNhVrSnYQ2d
PfRBN1pHzP/VlhSoEgn/Pt19juvwUbk7qKFgHEJ3CFQPlZkP9G/E8JVOGg3bTr+4
yBlvsyH+RnsIRd+Fu++GD5MWkv1Q721UJ8UnaZdSYhrJZIO7keGIq0QLO0Ex8ihr
5M1BOcdQL/y0Pj5xMTmBaMIj3w+7/I0W8g54bCa4+dEUYgOMavHVnUO5ZqLChqNj
a1fuaZk+sj5pZ+IRl3MvNw7VZSViNZMyIwjsvod8t8i+VKKyJ/RiR3kb7QeZYove
HG9ZAEYqmISY4VhXcbxlYLIfL9YmBs/9+VD9MmdI1Uz5o4d4nsEFDqjDjG1jeO9Q
bundev0L5zuS8IYW1fdgkxZElMCanin7uuNLuukHk+G4sAZ0vgMPsTtP+J2stNqP
i2XlcX9cV3pf737AzKvHm0uU1z7tolZD+lqJRknRkDH4XjQzDBREfJiqIhRto2qd
grdr7xCQbyGyvLqGqZ/M+Tvp0kDC3/Y2kyvdGWJdgVSKnBTcP/oqLn3u9tE5m/P7
3jGBM7M5Y8FDG/XEcpSINNp3m5sSuWc7We1ysTLPFJJ2nInyv8wHmcC36f+OrMt+
3DS+jCRMRuHcRlzgMm5K99cYBsTx0F1cZIRMTh9R/ZVLlxYBZHCrDEdJhg7F7cXS
Ki8NTw+XksohHBGgXMqz8KvrVZedEkholcvG7PSkxcg=
`protect END_PROTECTED
