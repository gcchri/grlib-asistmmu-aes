`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbXisnCQX6a6zTj+ZbqbygJh6C1wu4e6MI++F8wi3mTkeLFh1je8F9WAk6yHOu2R
sDcvhwpihYadsOkPOQOjk6CSyZ83Sd/vfmD67GL078ZsjtTel236VvQmdC6W2Ie8
bHUU8OXw/kTy3kpUOkH0TUK6XjRoj6Zorw7Kidwu3KfKc44T43O+V+Y+NpTZRvJ0
sX0Ow46PksUnoXjjPPu9BCo5iPhHEypIhJC1ICXQCjRrhf4dE/i1I2ud8ICvZYxA
u3OfN6QTYsvRQtmqMVX5irutl55HUgmXxvV2IzcUCu3Y3IUjprfO9R1vmqdswR/w
DwfYWmb4xdp/9p9LTbkp23K/KlsWDuIV0ef4z+TylM1rXarumde0ANnVSJg0dp+s
tHuvp1yUH97bPVvRYS+KrQ==
`protect END_PROTECTED
