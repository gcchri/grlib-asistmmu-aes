`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NDFTAiN/MZzgfr1UKZBGuZYPaP7U/QdGQJ9FpgP9TTxDmVzqeYiDVIv6d90PXRhY
dvK1Q2tI9quAXAq3E7cSO38VWLYyWczf3wQX7GJW5QIWz5Yv3IGIJjnyupUjCTSI
OoNw/SkIN59vX/JY4mh83UxVZ6APvPYv5x8RPUx4Hi7AWyzq7bvGM29pFIsrFuHk
Z+C2WkYBeMGo+DE/zrZeQofx/0tWN62uHhcvsIYVMkjoL+qLqBlNiKFiQyDIuuV1
ls8M5aD4gY4OSQY/oOpbWXTBzFbSG/O2umY1FEKvEpjFu1oDHne8y90mjMJdlPYd
1XtTsfmPb7vck1gCEExkDjBkdXjfR4gmLWRvYbsNgWlcuMn8HF4k1MSCBg4B8b6O
CIz5I2nPiEZDmoziNUSELkKuzeyxf4DQPajup4HnsbhmAQizH8RPKggFMhfvoLcV
s35JM48XNU81/LKYlUdOAW1Z1o15U79V/EqQUtB5bBBU8Tdvh5yJmEjx7zSRysrU
2CwcYpxE0A1xocK5hLakkjPc82G3FV+FKGucXX8T4UG1Zu5O73LfKP32arnN6Dii
pXFUfm5V/UD05INO/Tbo0cLYfWUrCqrebIN3WIfFCw0Y69D9V+Fye+u3ETteVeGy
`protect END_PROTECTED
