`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mogXTTiZUi1Gj9v6sZ+xAnNMns9SZBBjz5XGF57dmiFVE0rpKW/v3Hh/SUh5rzOG
7eA4tsPrmeTHfOv/e8GamHIi2EFQ/Dw3g5by74fOg/yI6kzmNulCvHfT76NZWTnM
0nyMR1rFxTUw4LqcUskxsefE+bR0VXUq9AE7OJ2myD8wMVv2QzxEN5CiRXeKaJHf
U3IJWV1qivyuQbQv6ZHBnfSUIhnITspIQf+qSvnBosFJkljqw2qVBXJJoGU7T5CY
BG3Z3DMxAWnEVfe8I/Yu6wPlUy5gr7inSgK0ekarY/t4tt+pYL4BFIyD3WvvbSl1
/cM/ddh7DoHk1VenAxDS7HxEp+5BawI2FN9waGyDHvi0vgO33MUWG4YT0euEChd0
TV4xF0/B9jTfp9y/mk1H2ULfp4QFMX8R8mfv3/pITj9hx0LJbCXSYhgSSwRBAnFX
`protect END_PROTECTED
