`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4QJmCgLjpnSWdbQaSXpZcIETuMr3QYSCIf8Jpxx0RHnyVpHU/BsLyeVuepWcWEZ
kwouL8WYUG3bowkatt5Q+d9rxhGe3uio9RknBClG5ThF9Y68aYsUUrGwVFgodPQx
Ko0oheIUUPwnvsXdTtW06Pb/T/I9fEgaGJNukfJ+a/reGtg0G1R0IH0V8pc/JWOz
K3t1PNZgJZTMnx4Lob59GzcWc9N37yCr+NVYjzpMHmdJ4y8D9iss9jeG+Ua1Gp4M
IbJw2xjfyxPX0FHPaYCWDXp2XA5aUSz65MJPof7Ayhwwoq+zdLdpdgug+/OtSapO
mZcHc65eEXcikcIxaEgtm7RDnW3AUN59pDuqKRDq5MMF4aN7g1UwH1lt9uAs9Roy
`protect END_PROTECTED
