`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsjMdD0i5FXx/2m9sJOgV//kpqFqUXu/D/DQ/K8VxYqU3JpPzkSvKU/1Aou/Fq2G
gC8lzQIl6JKyRkRpsByYlUhwmMljQBF6giALH0pzyZkwjoEXoQxcAYs3LFaj3YaV
CXdjT7t5qSBJPImars33yZeBn4EedfHCvUqhmo3EN2WOy/o9e6mOPrTbmsJw1rMP
4AAHkxZfEf3vg3DWR39wYGf4KkT/QmWvF8HY+M/k9hvTZj/DwE8WG1flXkl3odVu
qD1oxzIbB30ZxG0Y1jOKcPGeiLOwVmbEw5XfmI8f0nE=
`protect END_PROTECTED
