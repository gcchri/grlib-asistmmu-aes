`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1b4gX5oJA+6AHcSLLpYf7CJH9oburF1ahGZzW/rM4375y4iE8bupb8gaaCmO/Ud
re5MTO9KhoA3xoBkpxrSIHD6Yq/FouMCbNnjf7zk+6xhohbs22XomTeJ7JyQSRae
Kq0NjserEv1IE9Z+ZxpzhBgafV8uhnYA7ht47JciDSggqfCUCsKf6rMcwUN3Of/C
150ia+u40tuh8G6ZtgMXIC3rIAgm7O+VBUesVN69V2TMlMMmwFfU5fr7qzAUHlgQ
HwKDAGovqgwsxWocsRuHC6v441CzJbG1qOssBNY3hSuDB1GmhqFUb2UvVaiQ8HxO
oZ7Y3/lX7gYT6JwoN7wxjYG9WCFwIdEN7Xi317uYbgmf/p5vYe+MjX0osA/bPk9d
86v+HV6Qw6YNrEi3v8bgTI9ibTQZFOwZeVjoDs8WH750ETTDHvoDHKGEl4sAwVqr
fh8HnDmPqWW/hKd4nhMHx3WnebLumlcr6v9JH5EdcGCihvmqP9z3sZaWmZzaQ0FF
Li853znpOZEmMc5Vh+KS+DzrxsOTBP+AM2ABOYpsnU5qp9wyeI54GOIOgi6ZQFdK
LeyEMoRez5Sx4WuSnFQ5zyDgbJU+nbGuMYoLc3xui0EaaiTzJRADmb1fWwwI2o61
pEo1spej7a6xXmaU2e6J7ghOCsfkacXROScunFfBIOCPW+tgsV9dpUuwgY2NtNnb
Yk3/dK2nP/50PiPiB+nu04JprHZYp/B7LJ9dW84Ij1B1e+a6lHJ6HkgEH1fusX6x
/BXW1R3lZpi2XoLMQhF7Ojurx4yqs58B0MXn5sTohmyHOfK/YWvHyb4aHZRM4oF+
wkebfebIFjVzVqWn5MBc7Vz5nfH6iQPSqSoYVmGLx9KRhNV/BLPupwBw0ywfXqGy
HSLDnHSexJFov7g7HjCqodRn2RBp+oGtUYpTK455USbiuxLUpu2VBTdSKa/dsQkC
Op3HsB1epZDqvGC2RMzDEuABqinA4apPfzQq++gwCS+NsazrY5Q4zLNusXX1+SmM
ZSJj0eT/TDYTObPD3asZeySJqKy5EgL4TSpUH93ncKIH015zzbQ/CWmYg1NPFidX
Pa2++bEzxHwuzTODXwWSb89sdWJaDAxcuvEfWIYr4kE5t8+hPJZrqPpkRRmsDW4F
KWqPQepdhFIGNmqft78CIOBpeCK5O3SpZJ+5LZ2Z7+lhPXEJ6IDKVYdq+LHv3sZM
wzsGcKXiakK5Ixc3vDhBqc/qHBWGlmnG7Z0EXhQ33ZO42Vd3Z8k/92j1QoXlIOb+
prr1Er7t5LYPN2gyiGNexkqle4AQhCIXbS0Z2SDnyarMD4nvKNCZxzgAMqj+YdNz
9emNx9oXomwwa1BFc6M4K9IoQGtH2WDn7QfkJ3BPhB7a4aAX3zzG4n2wkpcCeHI6
0/4MtjDwRE12TZG/5n/I5xWODGfhkf63iZj6k/Js2glbTZMcZBHIn0aSK2Ccm7eh
qe12zttiuKI+tobcrCn6BZfMLFkSIn9nXDbxxbc77qtOETwpwVpoI9JHy4n0rN2P
tU9W6c5nQSm7BaqxE74YQERvK8g7P8R1h8uGkDDmlT0=
`protect END_PROTECTED
