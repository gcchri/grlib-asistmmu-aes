`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WcNB+A5eLfGnY0ulNrEkjzUTDPJOjDeTxkCgNZASqi2uvYpLC7SON/g2jT+vwcP/
igtIGzLeONvhMCV1VuskZhR83quCFkMnziwNu+otMdDygCyCvRtGzA7IFexvfCZj
fllYGaWXsj5iwZGlKRQvhMH3P2z+J9A7Mb3rK3noANgvx3OSgPfYrsR3kVv0/Yl3
wRtAcHEBUCxAKY/7OYkdYhxJtfVMVtI9xbc5dWik+myjWCi2bURE2y/GIwWA4Umm
8QX4a334iNR+j7c5GzfUUPhShgGIxLHdyLH0HKJ9YYNaTKXehyy0QJ+3UyhmzEB/
ewWi/8FxnANeIDCfuZPG5uSyO8h6BxHXhyZLpac9RIOpdPeUjVuqcGh37xzUstEX
kyRx4pRsVzfi45sxkoAF0Q==
`protect END_PROTECTED
