`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mlKTJ5N5CbU5oRgmKlTRmG+ikY3IOJganmwetkM09xndBrtgUxzAx3WGWVtA1jkz
I6Y3s4ArAPTe0JDSF+iuD2i7wFsu24NDvas5FIe2HvnAk8ZoHZmShf2Eid9I+MMu
7sO3utvEnWbDZnEqM5m6+b7ANWZgUn6s1vRyJcJcStUMmmQAQmsbw+dWMa+7R1+i
jwPKhI9OPBIhMMT1s/piHvrCVVt1kyUoOPfvf095jvO9sfWcG5l+/vq5ZRwmlAUV
wxb5EQgm2KVTYfR25/Sz1rHE8JRFKyFGphTIUqBgz2Pe9PsppOTv7e8i7N41HhwC
OvGzDbntAyJJ+s+KOMvG/X+dYnvZa4w2S0keD9YJJ6zVVh9lBJ/hJ3VaAvJaWQx/
kQWQ8PzBIoWsS5KqZhQRjnGS1j8HZx12g9Re+UvvXEBFlM6RXSPxXd06+adC9vn7
8wZAIi5IdCM69zUs3PJC7Efwwd35kB3p43QaSWVxW6yyEOjDGu+KAujkhFpk/Umf
`protect END_PROTECTED
