`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LVTFZddcRJVEo83w3ljjYOFTzQ+GsFyVFF8Y6xVUPg0KTER6sPZFS/7BPBgK+2vA
aC9yzMNLLk1d71wltxSn3x6rAcNWEG1w+NWkXnfGEPGqyilsEUKUTR+H+/kSJFa1
U+yRv00NIWGEMPQGYw0qVOngP9pKOI0uSFS1ELP5xJZT0tujk7dNLWS4xzP1uxuh
kCtqc6b8KAJsSbI+ECx/Ka8OlUQSl5y7P835Eoti5F+dWdf1p+NRemS0cvl3fFr7
3xeu/O6eH1l3RW68CMSu6f4pIwaWShummVtIfneNl4RG6+C0pFhUi77AqHPGrGmO
s18rWuTGQgdlPFQIyFxQju8E7yX4mvtdDtIJeYMl3p5evBf7cYCXORaPTRlde+SM
guDZguh95CYdhCdsG1fpzNMt1HS3rFBU3PWb/kQPOxGXqlVzdx7+MnxBCUc4AiRs
kdniEPHFH+Pyb5Z2n8faW1P+f2WYB6+ZpnwC47hkb4bmTDm2vqWgbFiTynyiiEfp
36iB8vYhWLuQRojS9Zp5TBZElC+NZX4mC8YHDqai6nY=
`protect END_PROTECTED
