`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A+Pj4dDhNSLXno78iA2rv/78PTNqDc+s12YnefvpJa/+8d4LCfJliMSk1a7wSXDi
6eM8myEv+N0PlyniDe86lus4nIWT2L3Vn/E950f2QGWB3jjamvl3R7rqDHNN0CsF
2fcLpz8zOxT5fzjuilbd8k6/lCRi9wEY1fmwYvySUQWWSdqf4v2C0quCrW9q0IDn
pbVPPHyytwMVhpJjA13jG5DZ3g/snD3Fa0s/vZ+XHXtnimzCXW7Knmn70QxwDbyZ
D9loLyuWZgFL2YhC+Sc2OPjGvFMq2HjxQ9thf9i/TKRYEt2F/g58MqZzWFKVLCey
pnrJD+JDvyEpmpW9SDd9uCgYlQMUYNdIS19AlPUdsNu/I7ujxX+pO+yYrJ+Mg+T8
frcCDv67UiXTKnyRLVGUYzUxA+S+ljBtiTICCLl2mBdPq9myupHrtjUfH2MplgdT
`protect END_PROTECTED
