`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WkfzFJhO1zNyp7V/Z/vc3YwxuX4PQAzHA/cJSCTl2MvSTDZIfS+6lDnILn875T40
OMQ3IiGIjKljaZD7ISsOnJweVIjugIyF0DJt+nLIZ97sVUHnAhs5Gi6vr22tctRX
hOjI6DFSsOt/ZBT1GL/3RXqS9V14I/YRfCXZEPqMKVhsijpqSFcA4XnqaRHc5kk1
gUWelGKVOLamr7AzDtgSwJyiSgbfWWO1OT5zcZ9KDSx9Yp/1fEOortxBCign6dA1
BTrjPzDx05z02M99Wh6TQ1mWI+jYVHOENQYvrMjlh/ExqxbRkMntYXlxPLZBjsTE
lAYZsRmxC8oc/M2OGA/1s9KbjSNsWAWbsG+DvtL1vFi5R6Ocl+VRZM7GIuuWCMfU
ktqg2F/ZKJm+ytC5/A6Qynd0RjhGnU6JR9iN7sUzmwBhA/RJGXIO4xLe3JmJUW/5
SYzURj1RyYQTQKxinl6nqiWu0rT2c5jGnpa3yNrVLBmoIksHkdEQsW1BNtLyhpM2
delBCEVQF2xKIFKXibivXESJjJbnynQe+wkFAj+HTNXHFlzt2uRQYV1L1Jv8i7Tv
nUXB7UqdXXSEjomO5ovhuC4h2hQ6UM8k+YMINW07rCYUGmWKTna9b4hzNtxvIMuD
lN19ukNLXlnB9WSECx47wEuEKUaYkPMN+UNTo+onM9JNK+n13Z+jarz7UD7Muwah
L4/QtYtlnn90kXHd+9tWpTfOMY9mR/RmPTD1WW7Z27LElu9JUFSB4g/uoOU9o5fm
m5VOD9wYiWZaMY44MEZzgfzjDV0z/x0ZxZy4apYArWpkd5PtSD74iPdgv7xQq0PC
zHlMZxGVD2O0oKIDbjT414UAYhvKHxUip34hd0/3ODzFxz0gcm5N8797qR5iuT7A
lKwjJATOvNRgTHkKna5eBLyhtwuA8BMUUv5My150Pu/yGB8M3FQtSkxHCoIQ4UAp
WEhoKwr2SLDjAKO++E63JFt/cFQwAZfVZ6NakjteLzhbFbDJTA+IO3PalYt5Bz3V
hIYuLVI7sKvffZ//VWUQ87zNDTarOGRqMWtCY9fV+RQ=
`protect END_PROTECTED
