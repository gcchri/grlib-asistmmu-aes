`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+AJ5Q82cWKEPVAKMlvLUIVTYjmwPHw7zKN432so1uznkOFE6z2u4ShSv2jL0dunw
0EbvmV6smAVmODtTjNosKtYECji9/BRA74EmfO+91lCs5qj6FZoIGws7nmwAT/2N
eyr3/GplIYobVIihV4OqLK/p0XjIHvFD3d6HVRTL5vzZgjzzlpOyaBc1xYOLmbSa
cXj9XTEUyYzN8yrzulcQVqwiBkIRgV8FtUlz8mbUb2WlFuabIXohEK8nXJYMoR+U
1g8MzvEbENOnhfX4UBdBc2hSEQkGd++c5SZi8mA6/uX60oPrYpb6tYZeeihZptiW
tq9fXcL04I5CSrVGT2Thxg==
`protect END_PROTECTED
