`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/LXVBVcu1M/sjxjrA7pk8oxukS2246UMZCkcYFafXtF4S5k2rZftBeL2leHuwwe2
b3LuET+OGuGnkeHSW11he95pjg+CZCidW6di+jBO0AxPLcWue3AxNXeR5eKd4bH1
Wdvf/EfB717NJkS+Nca811ZnxIf9s8McyCFOpWLcO/oavydhTddqJIij9Y8ifPaF
peOuo+PGbw8YPs2jeRTzPwgdnoqgo9Eh8EKotY4zngRXuWKsUip/bqCLqwpxBJvi
It4BjVD3HJ3ptG5D5zuOdJNFG2rXg0/EXRzNOtvcpLnI/pQTyCfNeI4N4+d2d4c0
sVBL7o2ktL0tCqVwUakr0MqyTD+3qc4ZXc/TkaCMdZJj9DRl91sZchynsxjOAedA
T2I3xyLaOm31KPEX7OcQS1P4JBe/1mAPi32i2A+zpIt0Js72XrFkW2mLk0h7W+m0
GqEC67yuE01OuckHOxZi23frKMIegTU9bQRuY6yAgJkXjmUigQ8aWycNFb1zyjNo
RO9XDbDFFT+YEL+u7p+ip605mzifCiM8dVmtWzTncf98LWyrgajypkJTeP7wzTxH
169kKSuC1H6Rs0e3hfg+ZjuW6sPQd38HWW7yMguwl+WweqQP55v4Z69EGy1Qj73X
U7qW2pvEHvljCPHGEM0SdOfvk/MOrF7K+CyLrlMCUCCahyWjEWAncuGFjB3lwVh8
iydhh4HQjwza9TlmWbQP6G4aZGRCgeaethN3Rlu8R42WgwpyleYj3OpLbk8C3q7o
9QimrMTbuQZKaDHLBwhEyXsbjaty1W9UhJlf5gPRIYEJrcg/lpRzKbrSkbKd7lpe
oQt5ccrVK14BJjBGH08huqmyMu2lO/ssw4nA94cTMPiBkzObGBWk0g7dx5LnZoZb
vJxXWBrJq7SxAty1ocQ1ShrAnB8oROqcPOJcd9I1jNY/8ddHC1zdtnln2RfzT5Fh
LCIRU2Y+sIAs8BAbgfilUjH4eEpH7gugG9SNWXXz5uUY4LQoE17ACqlNE8Dfyy7y
8NZPv1pBnmhBeMVWA22s6rTdLo2tq7VhkFrVjknkBJFHgtP7/rAJoRI8F1ncPIHX
JKOITLTBaBgD8er4r0iFDBZXxBTIIYC9Q5FSYF4kQF/Tj/siz29zbKH+h2oK5dik
zkjTI2jQY5LP0dZgc7bq/o2dd98BftqHce5iiFI2DOeZHk0k0ZGrV6V6zd8fO5Of
0SYxsYUq0jN+KdOLfRSv511YFvFjQTyb+Nyx169sWNfE/0WNil1pQYhxfa5E9ApY
7eQZHAy54KBR0dF/QPx7J8aW6wAEfQ2zCYuubaspnpI++QzObQYAQJIr07qtYsyG
p4ytiJVFS0xAGAUuzwoNogBvDij5jWuNW4EvVMYOTioN9PMLcZF/nQjKhyY2d7zY
hS+b78ReAEaFhxcgQe4475SmXywkxzDxjJ2gjURai0IcdDEz7y0Shom/G0xboJ9F
qEr1healN9qsSgTKtGvaWPB/ShpxPNtIhk/j1o+0wB3v+uqI8I6JKCR+1Lkt9mZg
NSn8FUQoSZ5T2poICenmkxJlM0pFsrvLCBNuTqXKkfKpArRrHL/MPYRB5g7keFx/
7Azr/GX198ABtBJR+cNfRPKbo3Z8cJXNgKsgbO7jULb8VKTOUViQY8wMuZBcJnAi
QFs/mWSvv7XY+pnVJ3k8wieadBMC+wcQQ2F82Ujx8iu4rDDFUYCOLqgp21Q5TrIB
tYASPJgRA6xAClUMI1Og0YpVDZX6fNQCLd3cepkD90nuydf0/gmyMA602xzkMOfJ
D04vFqIiKTsWUVQFz9N7BBVPGha2ZMgBfTpA0HG/DyJO23SzNb5p/0/C2eMRvCyw
3otSfqcytDXdNhIH/Y5RTUwj0bh2xuSNWb72UXABLFvMeJXCkvaLGYUBOyxuNw/H
h8lWKcBkauCZqZJVuEquVyz0tw+Q+CXBIojPX5Aa/ald/3pt1Bq8xNDF6GwDh99g
+wO8BM+tYXlZZ49YxO1EgL8U6WFwKTUZuXRBWfSxPnuLEJ6ykUJDIMbtvWBvynhJ
SS/Gi4p2MN1wckrhoTcplOi8ougba2H7eWIIrdiGg8VmKaCu7KTSMbd3hXNsSXfr
BdsovzLN/YerQnAwfLfo4J0wFDhpX9RFWTN5hIbTU0Izo4DdgNW8Em6BBWFHMxUZ
jo/sJaLzRLC3FikMwmfqzlx903QNpMLQUD3LymLjQw34PhfWiOWrJmBZNj9T6svT
EVKdZuFoFwf3e6KwV2ZbZTCP3iKp9PFE5+KfDg35l8UlhiulrziN99voFTU8Rop2
4PrWqdYE64msbehB4fOGYEIi9EITwVaAkeuh9N4v5abgVb7nNCGH0+Yfb7KNBAVq
C3QAzviBWnpfWgxyNfESfPTw+v7v2XSNjQv/qCQwgRl9D+9zka+CWGgwUAQWdMck
bl2qSaaCY/bvzyCaVh1NxsAui6ZcVmqQyYSzXZZr7iI9FE/8yex9+f/xXL3oaEaa
8QZsMXIaA3BVytC5S7KrD381BDuVPvsg39fIZKH7MB6QVizcjvDZCG3TJkt3p9ws
zE31k6CNWYp7h4Z7frqtfeng1zoaoC/FQOjdovODvikkneBXD/WNR6F3g2y6pgdc
AHR6Wee2ouLWznKMt21KgB1CaSsgxPFG10zNMtt7lJZaJ+SvC2zPVbkTfEaZskZE
Swy6k4cEqKySF89wZtVwE+EIZ4C027+bf8/SPnQmjcWU6vE91jJ+SFazUiFwPwHd
8xJVY4NjLE8SNGDF6pF50bSUcb+gdjsble+oiYIzkFGGbqusvVeaZLBMBygbyKcp
jXJJQG2JR4aoHKNVHWdtXpbuwNtZxQLbhZHGtWejKEF181BWqIqWkh9pLR/NpVeo
h66Y4zyYQVaJ5cRd6dHIi0Cma5mkbcShWYYHXjc8FW2iT3ZjpCmWCKVo+cUltYbZ
5x21+Hy9LSlJxlxRjcFZ9gDmMCPRzo6cCZFImTrZ+YGTpwv1GXkSCVPUzZuLtrAw
91xPRidDx3g4DJNxgOR0XMsSPEyxEUV9jRzYWsyvsrj9svj8HxToXVJUGS9E6JR6
c+E6jpkAOCID1eVRWjVnuo00kHx82YnLTNS1wZM/GAeCETnyA24xlonx0shuigmG
DdIxjok7KzpMFkiDTKzcQxoLG6r1dOIn7ZAlTSixG2Q1EN7oXfERoAwJryKlVLXA
foclBmY3BRQCHeiyvo5O0r+gvhuGmaoIoOS+miE0Ju0HsQKpS7Vpjr/yJF7Imu6d
7LjrmqzIdI1VSKsdEXzufgPnxHUoSMZQFfwulcs9EW2aJwpzgYZ1QNr/dSvOIKcN
T2a6G4JBE+mD4xWFugOt9wtqSZC0nGW4G8/05XuO5kCO4gbJVtCTxGkvHN7T9LgP
rd31HEY+7a4gUgYGLikweRxaOhb/+a4RpQNZgS2OGoPLn7ARrEo/ou668Y9AJV8S
Osiq+Mj8PbT86qlTnoB5y/qTbOgFFSeinmei72shnouE3GHfRKicB6EXzsz0YgT0
1GOxZPdsUQ2NSDc/w85oGKV3pIGLfjtTbInfHXSjRI6sV+soIs18OAQ8OyyCk3w/
m2VxaLRzqSFaOdzV+JDkaZEO7dgl7ker5gZDYAkPN/HVq+YJGkUjLteRquQsQzOK
72taVgjlStlFXS4L5hOrxXPKaqGVH7IPs65uhvg+VhqP/5MW7Yie4qYvJrCFPdrg
griBmor3qdoktnLmKm1hDFdVKkGhLHmsHJQPmxVa/RXkMX8kagzJWXyGJxzwu/iv
yjFaOobO2eYNNTRY2wYbc6PFQ7eAmIrM37Xn/aX431X+/2lPFRw0uTRrjcjv9ARP
pIUKXqsApZePoURRTAjjs6t8oC1D42sBH08Qh4NPvno54SQd3EqUXglVkmeEgP3p
rQDjFxegfOaM5nWQvP/FG0n02zinqP0YwKXWP+hoGrGBHzjz4BfMlmErNzr/rDZ1
s9jNVq5UT5KKvW31fQcdkMwz+39+S5i+Fmy5OST+k5u9KYtRiGb95HMhTsYH6FoD
APLADD5iLeISuV6HfWAEgR6cqrAYsfXXlsOyp1rtQAte4c8ChxX5v4d/4mS82DVe
Nzq+bwkThPq7ydu/tVgkHAlxPmN5q4enPt2wYfkkQQMvYKSPubm8lt/6BUV+hiGt
AEkPDq9zshu6GctWUoYMTnxv1nPCFI94xnHsDPezC9lOHEQicxKQlse9ybibCAzO
22bzRjp9anT48gBy5YxjhVuDE4XDTKm+Ew3vzuS007tMHoyRTuRbn0SyiL/DPYgt
Hw+Awgawk1x3q/hLig6wRHx851nGgf/sbbCyeqYXI4Y6MH4eJHqA+s6ce0LVJic1
q+lYj8qyNFwJqotZiqA6gUdX+O9G+RMWkhEbUCN3ldP7imaVaT500gLtZ3BHvFRB
5/u4kMj5edsTsYg94SZKywM20wsJ6SghQ6lsef8pKljisEzQWJvqd9l2etMxzLSD
/2oRHL1j7qIKBWXxx0sm3/GTuFV4WBcCv5AO+ua3ZRT1g6CnARz0Uxx3uXezDGFF
nfxnn4GuO14o9W2irizW4T3hL5d6Z0GcadjpBH+3aJuiCmf4eUJnQ+5m9FDAx5kJ
X1yrobyb95kJKoIOeXXrYOwxcPJlpcjiegt2Ydx6awt7KYzrXbXJe27YUTzEFD9R
//cemQj4WnhQTn95It0/SsDQ8R1tPFHu3Uug/I2ikRnpDoSVvFW+bNVgsXDAhrNR
GP0Mn3JrKlL3jroHTWlOLhBO2taXtHcvOcn9n5TyaGh55NkAvkIxzN7jV30lUiBd
I8zs7PP5Xh0asSMRKsGLi6vJWTrha8KIpF3YcD14j41QcFMui9FPhASsjUljWbLK
jhwB93MtVMNT0ziEjGtd/bjTKR2nGbiFEHQTXFEBf/xMveLwHdkD3EWXW/xfIr6Z
FatHaI2vwYuELdGnLhJEaTWtv3wTwlekB4L9TyZGVohCboSyiXA2i3APbQgIT1Rt
Tplazs4Piq3uDIiR9MpqPhbaBS1IhZR9OA36dgH7c9ExqyM0oVSuDeV6cN2nzJUC
LEPqSDAiYUPqg5GeaatiumDPz3Yg8qjrY1ksLTemRO1c2B+enmproOyvrJk91oI8
3t/2fC2kOPAnrQcOAr4IJU7boUG5usFWkcEEQNv0zMO/1Wuu2aZWXgNcZwXedPx3
055HLDA5y1fHlVNOe8BlqIys7W994VypjJ89gCCUs5YNMrLdcsleWJUqHPxk2vP/
vCo0v+crk1RieM0Za3iNJr3i1j6lpuZJbhUb2MCnxLGAHRGLsMWS0d1yINHrtC20
3hyRjc48jxMv+rOTjbEvWu+IrRRBzQzkhmkqDnERSIG6dsq3eM3bk4lPkEXFqfel
zMWNoGEZR6oRFnMhi08DffINDgstrWN9BAYFfgiwia6P0wnjQOLTJRJo622Pv1M1
uV0AMNlKOyrnQVlHyyn7eeSsFEoIazsel8Ly+Ru7cR1Owwyz9JXEI5CW7gdqcjcl
4d765tCP8m9H0gBVNouWouomP/zjU5w48meSlu2O4PoM0U2CSORFGcr6aanh0loR
QN//Vnv3ER/wxpBX6Xb0lsIcSNHwgNkO8/GkxzeOPdHlNpTNBL7uqg4pwgld5l7r
ZS1UpZDzQb5FVJ4mECO5rwaEJFjH6Sdv4MvFTBOw5xZRA7AXhS87SLk3tKLJjYc5
qlRTrWM7sKJC0De6tcu5trSvTsnh+s+v+gXlbLZ1P+8JzypMC2zcWKVCbXA8DwFY
fw6a3JPv4BTgDfOfyXjs25MCTTKfnB3/B5Ix1zHo2KWiwv7wUAhzVQal3IxwBAxW
rpPXqk/Jy9DelNYdWvF3xCvSe0czuABoFAKiwheTigJ9GMWL7aFyEUpJw+HfQOg8
ddzoX1UKrkKkxeYx4V9f2L5mzTC4e4P/LlGz43blycG+6JyIj4Rg4tO2sXL/6yrk
eCSIPKEwbulKeYKwlFvBJjCu6EumV7cHiBvNxmPtHi7L9fr0llDJTmUkx7rbBlkK
kLOQgJEgpwlrw/rE2d0Bfk5hrXcPc+gbiRL4GaaV0rGrIwQGwsViQPTdaAdmIFK2
SVEr06SWf3VRiSYz65wOlzHtqqx/c4DnrrLcBzWJmDnE6XYi0fd1SBGCbq3zQOuh
iVjSRSpH8TGYwD8cZVq/xwykjLNJeF9jLGFWfk3EwYzrhotDbmoMU3ciUfgFdPlh
8DFvgNPVHjGMbz+xEhV97JFsq72sg3LWu8NE2H21E9cTx3MHoDjyn5kvFbl0ZYf+
OyqwK/RESX0OIrOEXDnCI4Y9h3ifU0EXIPNqv5ba8pYM4Cc3QpCXol0KJ6RoU7lZ
7kFNejK+DYL/oA+B20vX8LfjDCJ9WalnGDKeDSYqajc+iA/H+010WZEtCPWuNY4W
TJkoVPz7tCpttNp9/hm7IDbkGrCBl9hfc7WmGITXYfkSKNyJG9GeKB76V1poafqo
PSeHTOw9CJzY4WYnjL5XJ9a7nOJetlpwMuzhWoeFup4FsGxtjFmRc0WfAkKx+Osh
6ofDA7DJJ1MwnlkYk57DiDMuINPUS7tKc8uxgme5oBL9ksGHTCtIxWMPYdhGqeQH
wuAH0jbshyLQejqe9zgkqHGupMe+94c2v/t8EL5BBGRtKTbaa77khw/EmumASAF1
Z9wprLE9kHoZZdhGaE0ipTsxb2xQGvFKCOyxLMTJn+KG+gVBGUXHZgZZVWS0yB4u
UuK2exnTlHXvi2+x3vCuqvuTRhFwuB4FW1Jws/5PzEznM356KfsJh0AVRSkUdko9
vZcPusYx/lT37HEPPpY+NisMfj/xRXSdETLe7QwMdrqofpG3be0gA3JGa8Rst5/t
8ZDFnoW50kjrgMmq9ikYEPNK32rUlg1zjm1uTOR6JDoUDlIqt5Z+kRxfeOWGyWJl
FaY73aF5EBaDRSlwY5jPfqNIX7rVIaS7FWGJ+bqwuRkkaolmqV9VS4mPP/MwDp0V
fcErH9DRts/7Vis4c0eEQ+Et4IdpDEVEM76PBxU8iPcOyU+IHIrvqDu+tdLtHWfh
SOcjicCW8w+l3Is+xPOarmBTU2ng8YJ6+bQAWXV7pxDAaGeM6qNBzWq4OyqftxLR
mvT19DSfcMXOgozCzlzVb+Ydwo4YEQ9Dl/ocg5a0X0yBLDp2QtcTYVkLYBJXgsi/
9kHn6ltNNN3km2Dwhco3WMwBSLWa2iWMzj+521LygGiZ9NhxFvjI907u8164TDdx
J/MArj4kCgdV8CFTh033Dxp6dwQ5za0LQhZQ6xwjY/i3L9StL3ouB+DgL9lv+PQy
3OjmJu5C5tQPQfpYUwF0FvNIBKONWXWzg5Qw8kHDN8omszVnW5aGVBzIBylahsl1
9BfHpG0o+7opNM3GNFXIvciHL7G72uKvpkbWrHJIu6WBiJQFFHPiJmEHrnciNc/U
iRvUVukAPAB8/aQA2WEshe2jjMo7JGpkhi/xxhmOsUi05jb3AxG8qgcfuSHEhlqx
AXrsY8ZAeNWup2w/aHDrT9ZPJqFjVTS53lIsE3DhXT6RQcb9fhSwB9MK4JA6V2EM
6s+yjeT3vefEN9dQzuFIuP9SH24vU1ZnZqhK5s3OEcE6IKmci7P/Rt/lmH0ApdOS
C4T9L5stxxlygl7wJvBvBcuGd8hUubflzjME8Rl/0FuIiYFyEDM0ywheEQw50nif
qXIbqPv6NmBeUNa8Vg7oIVA0o4ZfnWEzj7+FuuKgZRksG7f5/FA5yvuBViP1hpw4
1C7hwU17hsrhrmrjkz4adJZGDaDF8a4xCUvDu1d6WqFLAslgMgBLMdoY4CB9Xtu4
vBWasUCwpyo1iE8w/QqQxMg1mWXFgJ3vC8WrwD5KB2iSg0Q/AwXyE/tDyvcR+s6F
SftcBzjUgSjb0VMtfeIQon3BSpZzSU38BHA4WRypBHr7k7F+3Oc71q6+O3wHBdoI
GCOOG5DwO94PpA3qg+6YHN5R/TnBGXLyv0VtuAwORpBqN2nCYRljDkTUEDt98ya6
xPEL59wpr1tw4Qse0LCQrdUK3JRSVaEHwNLi5RvQM/3s7xZrKzWR6/vlirJNNOI6
FqERD1UoovKKGvUNUB90rAPgZzfa5EBZkNL1mj6aft4DNUUXYB4vO6KkUBxHx7X3
HgQUE1eUXY24FSLgJPkNONwH8kpRJgRwC8n+hQ9mqb9qv9dTpMCx4cKomi8cQzfv
Zs3RpsLb8kQwEFE+S2xsZjDu7aZwvDT4xJxQifLfA3UJYqlS5xhtvPrm0RiTb88V
tggjfi8VqE8UaTXX5lCD5Uxcr+Vj5nMdUIppCqD9uYJI+5s03Tb4qGqc00YZgBOm
za7vO2hLFHfxT62y2f308n4hlBlvizwn2Nul+fJFaHLRysrPXSmA9OJaJt6r+2Jb
uKXXTV11vpkr9Dhc+nS1Ylve3KmbUsGdBn0WUraMpeQElzFof0VYeumyhI/Cqt1e
DQHivziWFOYfWrAWFS3+DjnIOLen/d4NUZc9Wt2sORFU7KmNkMvbQXQQBIQbKPcX
mxNJP5VxwBzIlkyBpkpKkQAnIFVTCFtJ/Fb8aeNkMIm62xeva9dIxaqlnRTX4yLv
l3XAP44qg+k7qirrd8ERM/3LaKl6gA5yGH8/gwLvcLfD/UYPWk/y4/aZYi9fSIuF
IhzX9TsOV3jCqfPOuNIG6a2JhWs5BSiLTUkgRSY27W+wOCvp0JN1tDtqRiumxQVo
aBXSinTPrZi3JAXrlsJdJhMtKAml52299vmB5FQqWZCtiIlaRl6PxmC2wj9wrOlU
djlWnM6uOLhIvbsrg5/dszPGeSd+zAMQns7SNchAUv3tXv9dFXhhNYbWLzL1TsUe
aqWHVGs8tnY0vAGsZ8ycaMGbcpo9XPJc4lOfDe0dKsvdsvsgSMwacVpNchLCSWwt
k+WMLeV5kOZSDg/rWKTi+D0Ur8bU9SsZ13oz/R9waIfATIoLnwFvDyEnlDys/qwk
tXCcLPlI9Pbz6NDwHyT1OBW/7p0vclhC0aRG1MlT6WbuogeIZ2ivqYZgZAGcLn63
TsBHrZ65of9aFl06cV/l833ZQSTJ4iKdVtRKAWD5e2hg3hvQAwy9zzpZvBjw2Nui
4XeOPYlozIwFEopjodShF3jfffCz5cX3BgYHUYqY3j2Q7UEHzOomQ4vocitACgvS
2rd/YQLCqM+UtE/cbXKKwjpC7ROLZ6koVd8ju+OLSPnbNZ/mG6MMrS3NhGHTvjJ2
R30Q/M/5069MSrK4s8aXcD+nkq+e2CKLjc8U9u6S51+DF+frXxEKU2Eh5YcufaS0
IWCkz0UH7lbagL8ROOlJITbchMrDJRzY/N8AyuoLyyIanJFxbZ+hbna3S+8vIMWs
8SQt0NfcK7aTMt9vjrRIcRRgywyvHzAYlLUA68HlPFERYo41IPbEND7OyMEkM2YG
o2JuurxTg7DHWbgq/D0ZpBIEnNjGCRM6Fwx8T7leksOq3gQ1vEtGodxK+26ssTx8
GVMML/IeiyzxHAx9iT1S0xWOUkOGt91FvDT6FkZ40v8JujhXYgfFNwccwHtQPn8d
hkmli4bt7reRPD2ImH8fV4xS7qiopsUhkji1WF5FITxvTPI2uHNona5QT1Vl6BS5
b6ZzqBwOYJltU1flZ48XVVSJWaiTgKq3sZpMWLaUNcJOe+Q3hbsrOaTzEv0CtAqH
ZOdXlyent3tCv5JOiEW+xaVxVAPLGy3n6FGvTd8/gGyiGXRbe4SbArxUFQUTtGGH
DM4Fz9rVAUPP+hA3pcoz7aaKxPPu/CQUyfOc3Pf/3UFVPY0gb+yWMkOGBxb4DDS0
q7oIFe3ONDQUmyKuhRJ3hc24v6VqIKb5PmVpgaj00bkskrdFLrJgx0M4Yc9pVPLU
kjToy1A1s1Jgc7EXhZc9EHmuw+i0w7v6ZnqVxKXBam6042ThRFU3geTYaoOfWVkJ
OiuRP1/S1fa0RTc9pGPJxhVQPEtL1uHIji81j2XOLOr9Ad9vGWY2/9btmpCWrKm9
qqHH4EQwQPGI9XV8gVjN3410VZKqwPtGCeu4gpGS9lFQrRy35x27Xe7IuXbG7kV4
5AysJxNCmMQoefLYTVD49TP1VQbqa5kALazBDOxDiXJyeRgotjGKfugtKstsuq3x
uS7PTlARvKcR5hXJal+rxKnYz8dDFI2syqO9rdOy3RtH2Elyvqn+eBEw767m+Bgo
i7ya/CDuOLRRfyGRIClnT0da2/nr33mvDMUvvULIfhHcO5U8Pp92f4n0hB9s+3yv
LFMy75X6Xzg2nQnjONHX5Teassii1SCWL38S5wIH5Mp8XTHBwdTYwQQU5ON1qo3c
wVCz5224VAK00Oxy3okDthfe7I1Iq0xkX8PI0aq1hVyCPiMM/urpCKYDO1o2TqtU
KW3jABFbNn0KwByzepdKA+h6WWDZPLFctYGlstLS6Z98T25NzyDIFYm5lBdaBCwG
Xmj1nTUhZYUTrrkTGNmTPS7Z3SQZWh9SwByjCYht3y89UOem3CSZuMX1rFQ8shTA
crdPruuF39DHn0URGUJYt86XStEDxB3IOqgZosGQV5Hxgu8w7bhO+89RvYHdGWKT
fpFJHmOUyL90z5g6rvRilYrA+YzOPaHmAEYPGax/BNc5PQwHeOGQq/g2G/1Fqtrq
+0GHMaPnUgP2WB8ovttfoLeGSknjPUKvSMEQxxvZx1zL+loegQEsUMzZyerJzBxm
zNRTgIVNO2sR6jGnjXXIqEsu9DSNsOJJ3ktnBlfWq/b8ayvcJyEA4miM/1aBxWXt
OwW/Hqp0e2LMP0SNnWLW9s7ybNBlN7ew4TWzP5Eh2EeIUChNau23esEKfzYQ/ldI
ZA1Rwp1MywAgAbLUMEn7a0caA9/qE9pH8hoR33JPNO86y82QBJ8rpsu16o1gsMix
2bchffBqnKGToDdmH2Vqqp4O32jcukojZvyzGI3NxrEE3nKjI73Rqfb7pncMka8F
Mo+gy9+zjXLh1zBK7BIWI1LwKqD5khCBHDdnoXBdFW0vk4MGZ+zq0vuc7pe8CnAW
T/YIBQl5n3m99f40Ca+x66o/Lw6QpFbb7M7R9zP0iQ7JJ9DfR4WDIkxGwNLA8RY7
uYcDccCWM9Z8aatf+teInbWyS7kWdJAOaLOkIVSWEVDWYycSTbSbmKhZ3EnCxVM8
wJxbasKAubZVdzyL54SegMEh4voQIvhb/VBot+f/Qqrb8EVoqNy6sfAJbu4cqVya
GUD81jMUMO1WKUanunKTfJKD19HjkgRUiinSqW/I++4sigsvX+PYdQKnmZcVhAqv
e22r/gjwF+wsmzpDsDY3bhQdI0tZ4Z6WEWmRn+0lQyC3Yi5vgj4U3CVvJd9G3n4a
DuaoD6CRplWdD/IXb0hlYWrwYS5ZeVoEFJxItlb9OpqWg8tl+irxa0roUX5idqiv
EOZeOgeV7gUbU3G6VHikDwCF2dAuJFHq/JxWtL0kxODo5Esl+UsKNy7PN0nBvbMV
/HarNtXeJUvHUnKVbWDNpftU94T+mTzIobNuBl5CqXi77d1IjpR4lwTtQPQfoTxJ
Jvv0/44suaFN3MjT+9ibtFK7IgdDo59ieTZDWByiXNNhwtm0nAMRm6NAzSBbP973
honJobFqVCXizSRkIekhqSucbB2YK0KqgusBMbDWzYaY+/oZB9bhlj+f0Ht/19Bd
pNedV7BLx8TIrRTU9jWBwldDBeaIoUW1UicqvuaXrOuC3LqAlNQiyzRndcRi4edU
M+hL/H4ud8n60xQzrHxaXihEefT2slok8S/leQkb7dXerBRVX/IdVaOeg0GFCrjL
na5QDsCpZ3VLSAQbSLI0QqD7cWmuBITtQGh3zAd5UmMN6agxl4W4tcpYowOXxJLQ
xKDH0hyQ0iTOyScesxJv7kY7E8ctGeUbREp+yMWykSwh/BIPS3c97tl7IYwZgKl4
xsQJ0fXyGb63aFNGn0Xmjl+501krukcHTuIY95QkievXxuoN8s06Hx/6uc3FCmWV
E9l5JZ9Vofiq4a0ZVHOmBs4AZqMBNGLtg5Dd47lXDyBpEUHFkt2J/HHX/zlz9snA
wsBPCpAL7Y8wwDena91IjGBujqPdiTVLX7mDKpcfzZM132848ZEeloaABejf8tg5
EjSR6Etza9Se8EOhdly0jaOVABuSe53gDwKo7CtlbWGXJXoeypE5ngJpNR+K1TzJ
cY8nbuj4fPmny83Fa80xRYg4aPxO8QqAf7bkYZcWnaafeiVGVEqejgvs8RBdtvu1
iGqq29CpsaL1zAJVVGCkO0zTiKjEMacUSZrhtJ/cUt6b43J9f6SX/dFNV1FwrJne
U7uK3E4WH4Rg837yCbmKJAw76X5bg//6j9fj8VYRJW4fOcGYiZwWwT7gF43YkTaL
pD3LpDUYJ75qz/900S/oBQemPKAjmHHIlLczLp0RZGCRgZyA8+ji95vjgWntj9e3
6+gMEJnpIwT0Fk8btk5ia6enS7ITsXyloDvnG/9JsL2I+NON/J926eYJkSY8ZKRZ
YXb8c8v+LrmPxV0sokJ890rgoblUVVSAVBniwLDWn+Cmb63Rb1v3BLbB4o2iTyXn
wM3VGeKgECGxNlLdO37aDdsj2McbF714BtLCQDjTS1I+NEI4+JcpFMlKjskHg01u
UKhIziN8HTaC10DUFaiZBm73tb/3S9L0A9ao/IccSR8C8WuGXVM+Bs7VAmDGju9N
rfm6EL0cJ8XeIBhr2zGPhhY2BBdf8QLyywly83KXfPxwse3DiyvBoaf0i6uQwpcq
DJ1xTUPpwGLC0KAJ4fkYUnavwJBjpHyIBblknG+h5Cd4pFLSiUJtViGHVHYXQO/h
s66HF14POFwtU0Z0PoeWmcND7uTtVt5FzyI3fmyYHAtyPlDJ6+z28qhEMkWJJGdq
7Z81FjBHol4mSgFYO9I0t6dnDw5EohQWI58hKa/EueNWq08ByZoEtbbcfijotb/R
vQRtBaYaVXsP5Jw38lXUNDxdGC986Faw4ORujX0xlsFETfgXLUABMujDTS/oSaHM
Z2ysAvFFOdUUI6J2xH9LahMgeDqiAtC7EqLZf9JII4G3lJna0MIc/18c8XWMPHmr
4jv9Rc8j9gSWJtpt4h9TFLMZ0eLWREw0aFi4lb1AmJ+JZHQrsMbRqzlKyXf5HO1w
IJDHDQGJcq0I04PtMDrzTRwdiX3ykXQuisL2BFNcwfEQzT/5SamzsqFbq87oqTP6
D/ANVhbHOSPBEaud1W2Z8CCH/JSBwDd2u5G7b941zLKA1NtPBtpWMZ/KbwTp47IJ
MU2zmJOfzKV9hnJFHs8Isk/60/tL2aqNGsZkjdeB69lEIMb+BpTMiXDJBP0Pgynj
Q0NHXvaJuC9+ZixIm2nzb4n8TgpK/ZiXa7SM9OAxiOqrb+hjqUO17HGSqHIk6HOs
ED/TE+8F5Ndz7lkPGYBRcSRiSKPJ9aTatWvWLaMhnq6nIgn4aQ7cI+S+I6xgMSrP
ASuJWMHBR42LBsLP3vTeCOkMBvBgEltw/hKV411kohiuz4026eMRjGcLoQEhFaHj
iGUfHHCDKqdEjIb5oyFbsGb6ULxQSZR41gOhElPEk4Cr3N54TTweipIqKME9c981
EKcddshWVH+NXWelssI0zVTdIzzyzSnKa91Te4fd0Pim87StnEMQ4yWcx0C+8MCa
uFbUMuDH8+53CizmURQ/kt9Lw4iR55zUaXUDVAklw66NzZeZubtWo60TkHuUPRd0
Obl495Tr7Qn9RdgE3JwdmOSCRs9WXdnXOyATEOEmNBtj7RXBrOUwg219OKQMYPSl
6D4yJvEPkzdpfKKDalS/O4Fnf/UYGJ4GHTmuBsXbdhpfwGC68YX94aJFL1z/9MaG
min4A+m4xmbsSgRbQNFow66UyJRyzuyQZGnDbkXcGVYUEhWiegQLooBiGKBed5VO
i/o58pKoMaOIhpfnwya0paKyFRLaXvnvbWp8bRebN7X14M6NdNTXNGwZWYLuY1KP
kEKqgONpRzKzVQOiNx6mTOnonLGE7ItC/tdHtq3fg9zkR+odqloY+HGBHu7J8d5/
RoB/WDPwKeJxLAO4pZR/qL0kuR8yrN9L9TvmCQ33EO78s83iRcBIUFxs2eYCG9+u
kwa2BHEB0I2/yLucqtgbbSMcj8b9ShDSQ81Pn4kDi4nqH+HIy1ZFdWJeNR7LaXyZ
51QANecfWmtlIGs2WVcAhP3Vy79y1fLWpbEdTWEsbO+u64XZ640srdSFvdkC6aeE
r4T66GIpqoYafq8sfFvz4YGHqTxIylCbK8OhhJNpI8sf1yi3M+7q48+vlepnQK02
8QjrC3WDyS43osl6ZTY2RgP9LYfxuBZ3icIxNf20GhHAAbODOVkJhsKkSJMgFjbB
KiS93km5k4LEfn2nvfYJeDkCJDd3RIi/DDdMcMMHpu08Wxgno4qh4QPbJc1CO1OU
bRYC96ZjXBk2onah0v5dXUtAMDSLkHcnCbabXpalLlPzfO5ukuHhYdvY9fDSV4WU
up2gswdQ9KD3S4yaj4Go8LcwrF3g1g0z2vR+wpOFTKXAldss6Fs8f23n3AQWbRrS
V3wTHPqe67CfyWJCekKvsCqQ16iYKGKlXfXOBlow0hU7/7xwcmc+8DRb4skDOEqD
oSVmOLIRkwo3h9ZcfpOtt8J598GVE2NsjN+fnpSfScWQ2UIZcjEpHiZX60RjO1Ut
jdJwKKRutg5+5lsxEl/6mjOpSyDFdO2qj5k0OgIF9sCqvRm1JAQciH0/iKwthoH2
XIbPtfurtsK9Ej8W0FNv0mBLxnT7TIYj42r1u+vHwWkSq91WQcyN++1VCFKqBg1v
eiOnxaRdnZseqbPyqnWYNk77jI7gZyUfpNYzd2jcvThu15m+FOi3tBsGoFOEhjSR
jxHuBsaXGC5He8UQ1u7cl7MfrlRoEt2qcVZMZVHR2+owQWvWuhUK2/UKKBLZN6mw
cZi6Ej6P97y8otd1i4VxGZYrJplqgvzCRGfF6fmohunfpc0aZPNzH+02FSTRxt62
hCvM/w+fbHysCXFPNniGsL5rvoJYHKx2eYUbaLErrTLpaDdeCMuXEXa+AmVGJtuI
hRCwDiH29aJikYuMHDfwbYkLO2Z/AZy8AyucwBmufoSXHVEl/I6V2kah/BxfefIX
wTwDQ6FmqQUSr0jYbDmxiFSHtH9Rpy6aWhtIQ3sf6XvVLxffPc1CQidMSzJi5trF
6odyJ1S4N7hfwj8rz7r45RxEuoOr8TAfTzajLELuVu5GwQoRP0BB5KPdJH7L3Faw
re8HOB5R+E6quiuK134j2V5vC9suQlMbG78EkhU8RSumbLWfXXACZym3sLLiv8g9
ptdpd48NyyoO7kV9+yvzPIfEYIyN4LlOS8wSiJT/LbkD/rgC5yVDLvEZt4RKlqM4
OWeWwCD5afWlsmuXMPx7nDPWmPeQvy8tOQcx9f6bOXujMAHYxH7Lej7gE4aeNrTO
AtqJBy+K55HA+G8YD2Q7zy0jKTbW1B2L27mEQzoJdNX2VaTyxC0FW6L+vc8XoJw+
RjUGSM8X9VVMEb7wNuZakueozw8/pNAb/HJe0UpJHfT8iwhRihr0fugD0BHoAkzn
VmeRI0FfNPyZvb/rtFQNi8th6lXVoVqF1hsuVOJt59v82A2Gyn4BpE7V86BK0LJr
YFvKL9b2q4Mql2l9k35SHKarV6Zi/97zmW5osS56+/wOShAHeXvpZQfvmHM0yj7r
T/jfv/3THBl048LAn8IqgtnzwIr36Fhi8bo4bozQcBJz1qfCiQj59FgCEm729XXi
GQGc7vXwzm1ymLJXsH5QDY1rnNsztPLjKRCoSX+KM5zLFVv4m5Z6NObnCGg04FHi
+CntoPIDoY36ZfcOJ9Mrr/DuXcpXyX4r1VitMUTsIdn7/D2/HjlhnnD36yzsBkYA
xnrDHMQjFWz22V7FeU7FQ5lUK7Hr3+upSFvfhPHivC34L0/iOLeak0kpx4D4Q7Df
2QZjviFddMCuSEf50tt84CbjtSkBEYjn/7izuUT7YJ96hw3sqdoJmEv6Evx96tJ1
hEdQ64+2Gf0xWCHHaI5VmVesjx8PxyTLYlLh7MHCsqGznUqATtmwV0nRO1rKF2Gc
XALJCaMT6ieYA8jfJiZ7TLh02uOJBQsCUBgoZwBozXPFCz3Gqz1E/ju1ova1ThUa
yc73wwvMaNeVsZ3x2w2As3VynW9lIj/FQ0XnA3BIkF0gEqp9xqI4tymIPX6kfSi3
TXBuOKm0e8to5/eTn6GhgOC4UIWPue6hOK9IXg/022y6WenvtYuQ8J+Io4JULELu
HiC+SgcBA6mF2JWYCFKKqDejAjKHQ7jTY4CZhLA9fvC+KDVeapO1mdFz+FARoBiK
Flp1WD1T7e70TP1mmQxKVfKCWrbUKt5MQasin3A8sOguQHunkswf+ti6aS5D34s4
sOfCHGiB9rsAHTDaepp6P+4hHmjICgL+DbcGfTre+1ozhB86y1hjBnKMHqApPHje
bpf77x/KZT7A2K29bsrUAmxSj6viJUY7C0pUk2hdcjTTAM/kQ1CDaomilszGyebu
ITd5n6YQsC74ybOVmkyqwtVQPG7cMNgEidwpNT7ME9OnO75xTvZkm+VM9cCglSzE
a9vU/QE42sAXIHapRclCVRspnoWC0iifpdsMDwIOeg270ldt/8YP4WxO49CSpEw6
oRDW4kXmIZwl74UjhcJc+wHV42CmrYBsqOxbvTsH1Lg7ncvhVcKMvdBOxiphABnb
pJ4jEX+8P21WAeRpnP6KexG+2a5CHBTLXG0ef+RCLKZmbRJJSMTJUVCb2FkfEt/3
XcZzRVIbSye/oQAA21+tO5+53sHGr/0iDvEbehEZ+plAeKOaer0jutO/xbITpmc2
PSbB/Zg/wx/zIt9c2vxigKmxQ9DMtobqaLMWLmMGXtrxuFW3j17clQMZPR0d8aZe
5PAUznqdXNmwG+ihNZ6U+ZSC51co60AbIJ++FL7W3v/B/odNbWe3NEU1Ju4DMDNX
gMj5NCf3ZlsQgNrPMsazWqznqumRHytCEcicIDn5ERmIFCBbjXIQqaFfemt3pY2z
twabw1IXKmOxPOOYAxOUcBf5q8+bmvzRGDk4rWzlz4lNdB6mlVAnOWYiGk6eUxGW
5L81Jd3C4v2fEPztWJ8RWjvm22dswnk9zlg+t9Y06qx3UMQgzDi17R2w2Qks8/n1
OReM3Wj2XBfUTW32nWRulAS0MgOr5mAfrNinUm8O0H/yJ4rCHf2Zu+zcvAfBEcxh
OFpERDi4gYYuOlPzSB+LAo3e0iHu38SqRdhNwZYZavPtuyJ75muVOrl0dv7DyTDw
qpM8xNhtNrXw7922R3aoBAa0nHUw5DDWDiljUillkwYAPYAHKLtGPVe+pL8Qxitd
d8w7D0SyckLhd2mLyiYIZ6Cmod5vhISpK2RvZdKInUZa1SIerj5xsy8dY3kQCoa8
502VerxV2HefrLq5cABtCARmt1hyEpB7EA+mqmff9YaHyfYjNzDIAQFpQSsopZL4
XznG+QbeSnDZBtMkK5u/9ntHhTUczG1XhY23aMgZV5zndmk/ehndEXGmylCj/Fx6
uhOSSVt5eo+B8+SwRVxjWJdv3hLP2XRXRjiu/pxLHs+WMZgH4TmPg4RzPswqKcd7
GoVSnHw2oRwBjDnQoWI0Br+K6doKx5eeWdIKTE10uvnbrNCON2FDa+m7mkfH2Nz3
ipVVFpdbzLMlpp+a1b/+TXC0P4c7G7aOOgqRF+jjWgg2xevZhs49iPua+Czk3BKE
zqibVmRTmWLxByhyb0XZMA==
`protect END_PROTECTED
