`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abVM0tEOujw0Yx2xGhdrAcmghrM3EJeG1DhZGhfWpRnzrxAs2NQ5Ev66maMKe5kB
bAIAJS8G1q2PvU+Rtfj3cXc5YHoiAeMQzbAiWqM96gRO/hD4+F0MqDHqG3YDO/PY
DbXWHpZLpm5DwimhEa28zg/MKUmgRKk19N8hj1TWB26/4dOZV1om3crFWHlFYJRh
3nGcNJTC1iEN/ngl4oMcc5IFuWofWRTRgW8j5XaRjPkgdpc4lsKvU2r3cb8g5s33
10dZJhshhbtySEDDzfLzZuF3Pq5I1smC1jY1FABYEtD+3R3WABVL6sfKtJ4he51q
0VIH4+P4RPhPOL+0LT+1vC78HIy0G8MTOKFRmCSlkR4D7BYcd9qUlRx6MePj2uwV
X34mb6aXJCDfrnMUZcN9Ti8mF/ZfynHLZrvtdCbVsgygEtB6vZPvEz5GqRUqbg4U
A89ufsaL8KRQjwYLaUelN3JLT0esF+kwvbDi8Iw/VYlLCAFNUPtNDOrxhGfnZBBW
SOtqev0WeWatUSx5AvQNkz7vN9smqGFNI6V8Q4mMQNhaw2AnITsSpuFymzhOZ/Oe
QiCzlLX3EarVSggwWvnCYf5HiguCdbQ1Tg9OLhIhIPYfPjxJGH53/IneKs4ifimV
3yiEgli9mvCRNuQpJNkF0eHrsN3Sxpd36wFW1Xl9v7NrCtqcQ3klEskwQQEyuu3c
DFB1OMqkLD0hOgs2tx/XR1xCZOCfbOedYAorhCUKI2QDkJAVj4ato5+/OsUrVqy9
2aYGd1xtxspaytQHRPpNsnIcCMWXympseW/BmMitWRVzfgWOMysQSWkWSRbIEBL+
jTgTIEZcgh818whmRQYniWR8ro4r5fPqz/5B0S/kCmPAjNjJSSD3zs+e8j4pHvn9
VRkKqk+zhOzc9I1TtQn8fuD/N68KpFnaQA5uGj7v6S33fkbBWzXs6nWZ5Ih3ge8X
9xSGZtBOB7rh6O/9ZRG4JIr8O85z4u4wy/tBZpALlu2ygOASo1R6+JUXjel1yFDn
ZaNiCsZYadYydEhH1MBCKDwnOI9I74xDHhfhNx4cvakLPEfPuqZSn/blXEFE2AhA
PPaMkUPvRhtePGd0dYGduzHSZishBdxtYwt/xqBE7SQeXLHooKcG66mXdzgG+Vjk
Mm8wAe/Ms/PB9HbMP7gxjzoU1qx/BAfRhqhx50qjLc7hPri18KbAtWE4Gz2GXEvy
Gl7C+Wi5Q6oGnxusyd4Or2dAqIXEw2FiySlZ7eRQHJuX5F6ZsLKnkJQDXqnF3k1p
7fVW0ryTXgLmKCX2qKQbUyCYsOGFt8lsU+AuYONXNTkBNyKYPJLv6AyTnSGBXtiN
QtkjZYpCgADml7D/aKHlL+UIq3idqTzfG3Wtp4NC+MhbZDZMjtH3tc6QoN+lTIVF
HUWK/tWp8NaY8tw5Tho0rw==
`protect END_PROTECTED
