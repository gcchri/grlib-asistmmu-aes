`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLh3n07Qxbarv5OfdQJ0x4HiSXhRGti7GF4bEG63vyLqfojB9l59H1nntngwFWex
1A4YHbHiiiUDmKEHqE6z1MF43X+giOQWoPN9dO31FskL0xCyWr/pWJ9PYMyCsKeN
95PZKvMvSX1yiiK0F6L7L9K8UgRoO69LCZBU9zzZ80IaElQWGmkUSJeGjjTw0uSS
IJz1RQxs+hLYP2msiuOYTerwTKtfgA0yeZo12LLSUYHdHjQWILH8iLYQTTrCfaha
`protect END_PROTECTED
