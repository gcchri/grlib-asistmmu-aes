`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XA7qw9b+xTu2DOcBmwfavmxZylWu/VEdvURiNlBz/QcyeQl+RAHN/mkjE1q7vSA
uNQxTxnEBgmC3PADgwwNRhKGWfmM41mcg+kV6erV3zW/2U8RhwlGrp8lkmPY+iqR
ZIR5w+tsFkn7mPDrKaCxEme0hMh5+Gt1FVs9pGDygxhns5oGrUgKC+xOpsx9shFj
eadQLdEUhbLLLIcOYpa908t2fMMZUnmKPuE3tPB+tVmO7HftiIH1OLpE5dp9uds3
FnjTM2j7PbiKzyqgmW91wiXtNHcoQaOSJkWc/hiwnTu8TIT1Ma+Kr3mMpPYjoMZm
V/hvza+SDWEy0o2W2tYsvw==
`protect END_PROTECTED
