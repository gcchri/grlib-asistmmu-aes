`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wMgIQYGuOs7+JXTxcEBNvAs8purn2mFNeOj2ZaM5zGDX1u2rN64uKLNeDDzgHTn
Zkptb3Xom5BmUQ6a0/CYi/tCOIhYmM2Lj84irjnUEhYSMQ+Y+MKQmXED27/spOfH
N1LCs/08gxYIMBfCeb9IsgDcdIE8E1V81s1KVhbbUnyRjUIh/uAiZGGlO507jOy+
lSX3kc3vzuTNa63pF9L+H6bDPEullsBNMNcBtd7RoW90kRJLuVnzF1Kg0hk5qw6E
aFnr8pkbtEv6WN48Ckd786BhwgwSIAaACG5G2hZ/jS+WpdDDcxKuniMAVvBGLqXj
FW6P87lBfhW5xVaFkpcpeTDp84N1iCy6TRPYw2Y9330zkA4eNhcEJYaZabxicrQw
5Lpnezic5cL3cnWPmm5YpMB6RlTK0tASc8Aym16M0TsqjIlBy5xgp3ApZuNtgE3d
J45doHlBdR+PqBHzZwJCFw==
`protect END_PROTECTED
