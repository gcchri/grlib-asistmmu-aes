`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbllYFdALSw/U7McIxXKf1sTD94n7qLlItiqnfAfBB0yz49bBO+eO22iwx/YzeGw
6NC0U599CDOUQlVsfLyKazRzjy7LYg9du35FiO6CveH2gk6nBmd+nWqgbuPKCJfA
Q1IbPMQZ6TegqgZ4HcugBoZHo0jwYP9YTYjUcTYuTSuWdUQpEYIHuit/otimRlfa
MYaUVq2giVAGDKSuwZQOOeWaDaY7Ntcr5o1dwTNaFTPEXEiKcDCftx4fS+ZPzqHD
+GIZN4o9qFlASaz+jUBFFAb8ASkPb3mzsgVA8k8eQMHHe98tvHo8hwGaFdxEvgF3
gp9NbIbBNsxz+AtZsnKSSv0/mualisP1LYZYJX4i56sDhNipDyLL24s8TxAdyTn+
uPIBfngck+6PlbskHTEgpQ==
`protect END_PROTECTED
