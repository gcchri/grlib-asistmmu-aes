`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLA6u3oB9JtGTFnDAVB0iGfNxAo2ojwiv2jOrbofrTB2lTHgivGugou5iVT378tC
7lPx8h2a+bmLbeMji9gPbg/PmYee+03y/NSHQENDqosOuecgkvGvwJ3M/01B8OIJ
w2diT0Ie/fmKtoAJftH3obP1rkQDD58wTFX13q0HEHqXObPIOkO6kN7cJmZUlI8W
4Q3jFjl+1qouv1N1GllHRHMdM2FiVlBTPvoNRhoVGxOR+EXgcQllfQNqbh5YLHab
IuxoiheHor1yQm0E6iCMPzDEGSdtrbTCto9VGr7MhTQu86YTssf3PSX6OFACsT2b
c5J61lz/a2sZAZGQmIyBP+EfyYpYJCmPjcVEs7JPvCQz8LxC/fbw7h+vupTg3Tky
0JxlhX1g3pPCX0F+PDRm/w==
`protect END_PROTECTED
