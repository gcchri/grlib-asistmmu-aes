`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ApXKrdfynH7Xkrjq9bzEyZuuQ4G3Odv5gqiADeuHmky1QQPoYloC5N6U2iitLcPj
+Ykl148ePsHdpbFw0mPktPgIitir+o8iErnVmALUgSHC/iSItawumf/ZM18KsFWA
1gfHWS20ZGnkuNUSVSVQlSqK//w4OMiw6AWDPiO4lKq1odHgda3uKsXcTu5c1+T2
9YMWpzq5a/Wfj8mwlsFz0qLXokyCuxdFt8bXUyFMizHIcyX1oGo7CwX2SjGT//OS
BlB09E+8YYBl6J2CDsZNphkMwsW5AqAahkC82v6IMplGHPGwlobfCi94XmWsIX0Z
sMwKZljHULwLXEcHY9q3ZcoKNKC4wvyz3GlG4Oo7kMAsjNlUAo+vPKJ2V6Zp7e6a
ofX/UZnC2JWidiELV5+zpgy6Jd2WHrYtqgDDnyAJYLX8FcNmvNrcvMs+tSE7a2cL
8koUFBPxyNPzEvWtcRD/0DTTc1oYXrhbBj6Pa45yZCVmErWhOTP3gAFfJl5upAsG
yjbKouzLbXkz84fn3u0AulttDaMX503HguBTJC6PsOxasZTGX08wmJGminlVXxDT
SfkgejOsdSQMqKFGknrVJ8I165fekYz3Ztyp9p/RhVVrcpfk8tUWTtVsZFV7lJ0d
E6XM+scO45oyCPhcvaogNA==
`protect END_PROTECTED
