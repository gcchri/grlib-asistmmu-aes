`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qKUyVX1BmxdKmiEBjfvPiw7gUl75dD7PrSw6GRvcMKfjrr6ui59XB6yoIvzlVbPw
saYZkN59KJZhUNvUgMDd1zOLT6n+TpCV8N5LupNGOUF7FNFU5NKSkslsqtklQbVM
s+jwI9n88RB2mtCIXmgKSw1k8xphpREKI2QFTN5cKomkBOL/9S3Qp3bXv2+JdUSy
oLJ4AbGfLafkhDLoCjLTzrBcmNBFSV6K3Apzkf2P9lE5wD4M7cJkb992zyXYu7d3
2XnPLcD1OFY4zLmtZgEdGJ1K+1SNrjAb0Lb+kUo86ba+cMlykezXuC4eqtOHR+pz
YwxSDyE5UlCxiQbdhntmhyY+KSLYd2DrzA71EkICNpw/eNgUWExSmhV6AaJn5Tx2
vMKd/n9RLw7CFkD+SiR0BShD0NSTRngOnY+330glWf/FPVh3qNERrXFkPTcJqXvz
0BwpaiuaLGz6UaY1R9rF3tyqTvVdWobmJd+wYbP9fPNLHwyR35faPcopjDrqPFNA
pqoTDgIIBLQ5MBvwz7EomLx8VItNEkTiyW/M7O0uOhdnpZOEGyJqkNRqn+l+dzxO
phn7GZc7JkntOyH2heGFlb2/Qr8MES623Ovgh87dmgdr7U9gnCa5roH0Qr5+dbX8
ATpIbLufm6vGUwNouwmAbXqZ5pFindZ6kDs01vfwHFapkTDBPA4N+R7DRA45HfyW
9A+169lx7KeDlIysVlSG9YB68S2AJdjeGsu+vnm+jhIITKiSy1Sj29PsdA1i44zo
FjWP8FChA355hEIrEaxhOKQtpWfu77oypbh3x6diy40JgPcke1RmpoaSUklz1b5V
A99Rt175Zo5QdUkTC/eCA6OBUlYJayAxiX52XuS7tzs/wqZtCn8ys2wflH0UGiRN
cBCUNbyNdul78pAneX12/VY9DW9XcD56rSALyd/8QplvLOOgS3ns6pWH3wF/L+fh
4TS0M+fVnNmVlQTV7hTGe1U3gDSR/FAGRuS15QVDuXJGmzt5wzf/rKjd8sHWOdCk
0gFp9SmN2RMMH0rNttYoJOwFBT4Ah5tQ3DkPJACb6RtALA0U5Rklipndvn215wiA
ty2xX1pVhhNTMB/qKgqXgJl4zfw2KJuAIll82gHWVamMxzosKzexMdkOBcGq04sK
T8/pI8+z0AV9v3rZSuX10eZLp4IF6ckjiYXH7e6vEhGgO/lB+ZSYI7Ob3l5yDEyw
JHIJZOn4DvpY+CjcVzMDxyWytnc0mkZBDELkSdJOUmdo9aGjyc8wv2KfDt2kHmO9
0Idj428w2D2wl7hv+2Mfug==
`protect END_PROTECTED
