`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7EUkFIux+apnu+xIJSP0rdXPUlo+8c0GIOgbbucb3/AgdB6LwaD8SwhwCDmR6wpi
zehnbFajDxRfw0CPTkj4v1sIvIl0iXPYmClMe57S2pEw8EURjc+4At8jU+f2DwgW
GoO0k8ZTTleGAs/oJcWWD/khbTdcaW3lHGpogwt1cJCjID/tUBVjBAsKHsR7nMKs
SI6OK/EBLuxfB9y6Kn78nd9NbA3PRrMVKKcZAs+h9jRRIHjIbIfynvN98/J8Ihix
u/8Gig4/eyL0r0HktJaOXurue5oD2gWrElHzqjU9CiHtWgRJo7/hub4sJiQQuFI8
s3oB79xDzI7rTsd/IVADnCT2gTKPzDgXTfVFXrfj1PP6zlpx+oDFKAdi1DOAx9bU
pqrZhw7vODqGWJTSyLLUrCgNg2ASIYqYYO0GL9+UVs1U0KLyVcYAHYc8PidUndkn
vtQ5bru1ARBvc8q5Nn/GuwRrxdO+anHR5BdrDlx9nxItbwkKVfTCSP+l9k0JzOTC
u2ixlI6dqHp9kXce1tyC+GuDRQg1sFwQe9433GKN1UbHvrxB1WxFC5QklbhB0UDm
CGhFBSkXTfq+sajiVHTzwLtuIziqso7U0Wv4NgGLRN0b10E1R6y24i7EozKJOGik
YRWWlaxomLRdshyffXoWTncEPJYTwJqxdmEF62h7kkF9JrlJhDaFOEP7r3N8j+4+
elyVS7EyDYmLaOa7S8D1DWd0C6c3ODWfVoEkPIVQ2kub/eU6Q8t7VlT1p/s7cKx5
NPmXRP7x5eE4pPyyd3TVO3iL9TgOEt8BRy6hGO4SQwovOZYpZ4SSYA7a5cKOcqpK
zIWHgDsE048tPHUT32p1LKU2zuKDw5murI4veQYL3KDTORrG+JGWVWsY1Srn3vih
HHjWP8ebWBx8i9BVl6WXJzBE59DlheaFNCJ66KNo7TLP2rNs7W06MHmXHH9covSC
4KxH7UxO3QqW4ImmyUoXKyZy5hI7N7iIzG+UIvok4seSKNwcb+pNAB+3pFwumNeO
5SFgq24ZAfSle+u4iaZ0ElC8i42HEj3lNxW11QcrTUcDeYbtSwO6eQ95ML8f8XBN
/Q1wSZMirb4hh3k4MryHUeeLZVePu8G9oW/s1Jy+jnBfAYmhXeqUdonsTbLUOEra
oz6tN12QJQvS2pls0ih6ct+TP0ShW/DpIF7FwTAK58SNGVRyQWqqr2QIplPEIU6Q
c2YAyu59gpY04t4DKlmCpiZX3ZHMAAQD3994HsiuohU/qcSSnhtjXdvfm3R7ZApD
eIgGk9J+O5W+r9oA8CqS6aPX+gEDYThLzhklBQsgYVWmn4SkWchiipNo40Fk3jz+
wVKECrgdZ4aRVb3CGImZtoaVQxS5XSk1mZmSM0AL7Gnlvlk/vS0q30RBtrNBOQl7
2Ka3rOg6+/2XlA2SEUmHxCP1iEjWxnbSjOVDuZbP0GGpmvki3Eb7DdR7go1IAoSz
7iJ//iRDfQpdj6NchRdtnNcT4OaUzIy7EgQOuHJ2xIy8Jg7/kPRoalrAFHvAvrLF
+e988VHVonusZIS1zqCHupupfn44o5dP9KNrPG2rV3xbzVDiU2UPu46bg65oIROc
nHhCI5qN7uIxxGQD8AoYpS39pr5EghwoX3kYuhlHx73azFIseWrr67OR5cJsheLx
1ABYZ9EE36QnPpEDMnELKigqpKfBUqWDaQ7Ym7lhBlOk61beOpejst2h+MFIuLn3
+9Hb0Sb8BZZqNKTeB8GMXa/byhQBToOOdmVFsbhcu1FHlVxTsx0yGjHKq+S97XBd
ZtmCOFN2Ffi6Mne3lXDG5AjeitzLxrm0QFJNPbqJ0sKlpnHr7cIX9WOx0oSs2iyL
jPvSiMfnaYs9rR5LEtcSIZzUTcuWm6ptFiyCtkCeXhKqXd8VZDr1nGPq1cWLWeAv
l6sBwRPH3iEE7K8NNKugrdvHecj+7V6LuonrpcxiwbGCG09XHXb4Svlm3tO+7dCY
6WVE5RM6knCVwVw8NvVvFM8t+g01TwBVqZNU1a5/DxIpmr2CtXis/gf63b7tCT4d
NyR3/yhF7tp9IC0mzoJ7OS9lD9BfuZybdmO/RP6znrt9mk7O5Jr7232uJx0mczLb
3UYtk1yy5uyirhvJlm0M4CauXLDw4OOdQnMlQKnYT449S4QSUFDVsDJMpGyNiGj5
gTcraPpT9ta/A543VqVmTWDpMOR4vbHMu7k+ddh5Wd6/Qo2r0YQ0Mzawhrdo3dTV
dPt0WRlr0ozhhE7UQZDZ7NNuhg/dfYAoHl+wc1aTRWQUBZrR3h5svyG14bNJ7K9t
nhfGYs+INPYGMNjn30zYvA==
`protect END_PROTECTED
