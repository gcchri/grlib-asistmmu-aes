`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZNSq2SVBbl1+x/ulqJn2piNC/kATkKRUfXvUCjnEDEWon78pQnmy+bgjMfnyq3ii
6pPBihhbu9+m/nI+mMH+nIbfZpODFH0vPhgy+enGNr222MZ5ol36LtK4xlWTghN1
Dh5CWiAM4wdLQtjf//MQWIDxzfzm69lNdLrNyPglWYMA4lYACOhXrEL3B8/hX9tU
K3Ye9K3VhB3npqqJONriG4/IFdIkq6rrkMS958ovJEDfi7ha4YDKbSOoc/JjEVTW
wzsl3ncBrHjOSdcp87iZSnt9bmiE/Ck+dgv8CMxQJRNQMsNl0TUwP27XWkaSzEgu
edcpKwvw3Dx6kQpTIk07o8t6zt3xKS9i5qVLIuD6mSmwVsPQRtP8OcJfP65yHGLJ
yAIW/D7RTdw+gnmhIuIFN9Ng1SJ8kL1CWFfw/WXyrzdWb7oM1TPE6Epg9tex+OaN
Fite5RPtpy7x5ZGgNbdzWnYqnuZjRnkOU0bWoYS+yMvdL/uzhulDqIJ1tDphjxly
s2frm/DinWvn+lXkgce0GQuCnve1yvQWZyhdZUqhHOr7r/2xSnW+KRYP8opRi+xj
02EzdejWOerVP9AZzLHsRQb9wZPvFQBgLEiZ5i23w0ssJGb8lbfIbW0q8N1piDGe
0CWua/gVv6obnMnmhCqhs9sYx6BtuSBGMbGN9l313whk93EjjMyMbGpU+Pl+TX+Y
dcLf+RazfA2MPYvvjZlw60gQkUDGXZPQzbmb4SIm6JZGdSosofCYyZEennxQ5/92
fc6X5hc9MjDkN4ou/U4uSyof+4r66gfYb/jazuak1M2sQoY8gJPXaeA4CGfULxak
+P4ZXcyDDaH8J4CCY05Ig6lbQ/1TXfFLuPhx+qYp5DAQY+ewqq6Ibzyp5vZiuNg8
PNRJi4watNUUwkTpxhqqj8Xss3/hHI7rgoUYdTVS1UnhFsSqb/T5rg0A+uD8eI/W
6UWDJIiDTGEAAQVGFatFxUREBnLufjI/3/8EuBx77+EBCyt9Vs45VtdxrqtOd2F0
`protect END_PROTECTED
