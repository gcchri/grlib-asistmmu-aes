`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4C5YCCM7nylK0bO2k9GRXZ94Wkk1h98YJhMKcXrFVxpMjhQLGHweZO+/Yc0zNo0F
2JVIqsBZNsHsQavrcMaPsHlkjfG9+se5BU1MCIDmsZcro2yHRDZKaS3d9OAou/z4
9YPGebTat56c1LOQlk7LzjsxxsaVR2vsBy3bV7nxsd64mdQjZLINsO3KvwCcaBp3
nFqCNCvZcSs5JSbf29Ga6gbnDBF6nBpWFBCw5NBHEG9ptlNVvQpy5MYqmUTKJY8W
WEVh0f2KpqhXR3v2DSJfVA==
`protect END_PROTECTED
