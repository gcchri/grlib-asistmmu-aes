`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9qGLwvvIEp/DsH3eJdPfqxVsaevddlFkWIrgMjeeoUcP1FJsW+SX3orp7tbMKTP1
Qn99WaMMTRP+gsnzecby24zswZw/OH34mDjxPtWJ8xDWHuzN6AxmwQHCpswUgvjp
FNoylkyAuVYF31wObNVzp6ex8ve5FdXUY1miIFN9V20PTr03OiaE9Ps4HO3VgfMP
FBIXnEtUKiLS4kRMnr2dRr5I5JdMoVKRKeXutl5p9I2J/fiHDu4jU6HZOXGFUyCt
q2N9ZJ9RX8uw4LcKkWNMcliRNnZagDURETznXYZDyCYRv84OuF4m2tt1OhAwYvRX
tlhiGdT6SIRKT0Nc2Ng45eJfpfJPwJSzgI033Eicf4mD+CJtISuwERo2EcDZCwR0
AmHr8cN1mnQNXVKuLfDkHRd5wrN57hQdSLRdHMCLX0s=
`protect END_PROTECTED
