`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6QzXFswdWLFagDlFRMqxL3oR7yMUpIRQAtyN2aEIexpn4qWMpc74Yf4eaMbZT1Cm
fyaVtSKiWj5Lguuo4Tdk2tuaYAU38ue8xGis/mlip862UqG8cg5hsFbzXGYeh/I+
SRQGBjMTwCwKhGFcvY5gJz+LeQX4fGoUng+21N0gkdHEr5sKRPjO7KmURii81RqI
TfmdxCh7Oij/eye92H3lS7cUaDeWcn4JxBgWLRQvUtaAxMMqiBEj6rLq5TmbWB5k
4SSmOfoBmwFSl7D5OuduCTvCBH/XVGVbYlLdxDl2I/pCv+/3RALHJS8IXaeU6ANE
ykEHXPhoMf+fxo/vpgraIbNV+WIPsBaoS5c3ZLg+/HCUcG4FusXxlQ6GMNFA7pKF
fFh5Qm7yAiHtq0K7I3Fid3bIqfmPPxmhYlAmxXQLHLHzd5pUaQOYp9YQRbft154y
f8W+g0wijbm80oKOv7gILGrSHKjp/mBYkoLUfIRME7Uj8Ft5kNUXl35477onMKPg
Df0aTYVV3qXAbv4qh/TlZjzRXlpo/AOSpKeIJQmhZ8o=
`protect END_PROTECTED
