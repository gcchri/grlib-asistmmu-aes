`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulKjvkOro/6f6J1wDJRyyVxg8q35+lmrlCTGqzuHRmh4QgjTp+KBRS12mt8arXPn
5sS3zxtaCnBl8l4KR6k+REVRIbplENr1tmiSotIn8sWtMlqtXrig3PdB4RxgSZ41
gY2+rVNhVClxuOZE5VRUe4OdMIVVRA59AhmiJvtS90gaKPk6vsaj4cj+aQazexO4
D81RMkGxYXv64A/g/l2fy2vpkEwHXIzBKbCM8oJnV9Ld9oic2imxjmC0iwRiS/VV
n/b6+kvJDCDzf/mLJnjgD/caYt6XS7RBNHy0spPylI//SgsupM0Q8zIrum5FnJ9w
bCsoKW0LbcYXUZq4mo4HwlWqOR//U0QtkxkBYw4VnmzoDlfyf8tLFNnEtk3hP1xz
`protect END_PROTECTED
