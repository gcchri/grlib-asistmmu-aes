`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMWvTMB5ukzBClpWCmrHbZO/0GPHGHY/EKL7230xRd3N/g/8uYk1Ute7q1E9rcws
CZ/HfW+2cTe4lWgJNocU/CG5EAuQKr02w2+2Q4GEfZrVFuBpPuFbmxB9jq3Rfm0a
Y1TTa8cPLd+77lxb8UgIV5Qr4TE2f3v3brC2d7rPZ4/d9DBxpJHp2pHq7WQxcpdL
PY3oztKPi4bPFZce+BQ759v8ZQ9B1PpM50syTjQXR5rFlzxvl2HTBUmmKFwcTzae
JHskylRymiPWDnsOdU3NC4HC2fNKx/30JjIyly8O1gUqWOmenhoLQluwsMp6/NTK
E7FB3Bc25YjpoxETfQg/k7YnJgv0hWFph5s98XU+TsE7BClFHHzuzdlDH7yERJbM
DxCrf+6SMX3PUJpTtfbYKdySK+xsjsJu5ARn/xOkAcw=
`protect END_PROTECTED
