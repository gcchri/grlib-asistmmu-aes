`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0fdcI9gbpn8Ry7Cwft2sJQp3iC9RxLIg8DXhOCcsAGc55+x0tPcByGZKZfIDWKbh
Q8gy7rDcU0CFHBadHMNwqRZIr3XGlCPmk5h1jm2qjbmgwAFzc4ydiUW8I73dTTQj
B7TDJsBPR/b6B3cG7eJWw1ds//ba6pEbiZP14ObOwtawQCJVzhV/Bszqb1Qyk1az
swGjQMuHcfuBrDGYxzJKaBiacTVhb1K+C8kLqWPn7QQ1+0enlrZChuTrW0uMqZj4
NuSVi4bchgDbHAK8EqPD1nmYAMfTlfGjnzhSYtgKECsP36zyW68gi2quKU1qGC3Y
Eoo5RmfjMrK1r//3dlMxPCms+dJZ3HqDaDVZ2biUQd1y0NKhi7pQK/ve3ynsNLNr
6oBtAOoSdmokeTF8Z5ga1Alskw2bqEwBNeIwDHzZyYtarrt6iur3yD++k+XDeW8D
has26TAPuGpYxSc5SGVe+0AMpgSUK10m0iCyyksEw1emtXaBiyx0J7AvYHlx5lnz
E2SoJf9RLiLl9GbilL8336/N8Kzj+2gJzvU0uZF+VX6gUzgflCszAMaH6+Ovmy/x
v118koA6LsCAW0oM86OVNsfrjNCdMleJw1L/rncC4Uof6JyQdftHNObbBbSfJhqa
0etCfE3SX4pNt5lGKGnBWMnKp9V5SMd4EhgX9ZJx4GNZ+3PhILkH7cr5VdY/cYLE
Fbmysi4eh/7KxqBcaR809HUrLD3CLBKoJ/SwHLujGT/SwfSCIUiDLW0KHrmM8vZ9
HKfpXXx/zZedELdyaVZMdTn5jI5uUT8KAvKYHo3JbhY=
`protect END_PROTECTED
