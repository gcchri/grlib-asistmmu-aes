`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3cEKAujCQ6Bn4hiQsfY1M4k8r14xjErbf40RnifNCdOc/ElchDLjWeu+s4kxb3jT
Fi+jvCc3H1ikM6zUFF5+qxHI52kspYIOZ9T5/1z0KVdvK05RzvP7mC04eHzbSXtE
yhLDR12FJ+bFRm1DWuAQG84uERZ9jfFKVKoobVZ9wIcyJ3Qj7gpXnNGzcQrpZDsg
AXBXjnMCvfBwaxYSo5MhBZfiklh+SE6I+gR0fupvw2NYvhtDKzI9cPa3pfSXg9Wy
4ISCfWCGrxlqfaicMCUBc2Qge4SQ4VhhEoniradS0fA=
`protect END_PROTECTED
