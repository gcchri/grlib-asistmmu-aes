`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZyjX+h7HcGegGsDrAjwng7cTCCB6iIEfFlFRP9/9PlQ1XKbBdMwyea2iSTPuD5R
kXOEKhURLlADJ/KmVUETXSL+0qZw5A3Lvi0yjdNBpGpi0fl2zc5hyYtgKDNZwDd3
Hh0Iy03m5yxZdqDzQJrw1A8gLYJI4EmfxW+COnLoL9DunhtKsTlZ9Oe0PZ+mYqLK
SU6ja+DDlj7MZ4MRg74ors45DPH2UnthCiYCIPgTm4A4bJ8a2LIvyDl44rMVzwlJ
J0oFvkQczzgpvIpB72u/Y0szdolhruk+P4v1wTpBFm5UgidefbZV67v1mtwBJHaz
1iUznly5fB6xYsR86NFBdVG8fZEEsccDkj8/YauaEttdptkrtvp2ISO7Qqx3tO6A
Ad1KVE06/HC70d9k3LTUbjDVziHAIbvNaPuR5eFUcQ7NZOfIoOXANpYBAkGP622u
3G3laVXxnN8bjIF1aofDXazFcVr5Ud7CIdhgr+BX+G78ae6xUgjhR3vdFY1audCC
ySq6Ez6JN9c9hzu+Bw6pKFqH8o9r+vsiladu9yggyd+Wflm4Ik4ibE0zBUNvpZWK
9XciytS1+smuqxPcaaQTSX7p1Bp/t9zXHCNGQKkPxwJPfyXykm2CClPa0zONkdJZ
YRBNZEMRJO3Fw3//p0M1qsYWNwfR1XFcxleosxgKC2mMw3WaQBZBPdBzC8kkbSoq
6OXJPuHkycSkFjYkL9b05W9e/hKXUVzoLt6DkhrX3u2C2O3cyYP+Skjtmbo1kNiQ
jffo0QdI5WIuWuCcKbdm9HgYh/MF/WXYetYpT9XdTbQ+WKEDTfFUaLugx9ki2ZfJ
4LOxH6/uiqA7+uMTpon8i+FO+kYtDaWZkybWpSmCwF8+rxRjxAQzY1KWSejAQLz9
Bk8g8P4+tXdB9xY3sVpcuJXmJxTUwdnmeBd4ECzqaGApLmSbe1LhBdyrkKfMUIeV
neQtU72jgVHGWtuBjTpYKbCqVKZeHLPb5Fvpnncy5Vw/QZykGWpd53JSYahu7NbV
vHWyG4uvdg7wiAvt3hLSTYoeq4jvB3kc13JEWHB1zuFqO83n169YVWO/W1nQGVn2
IKNwc1+LHfE3mnFNxnT168VpHANakDxuefqXKeFz7fLcBH2M+vgFL4bqr73GQMdh
DEULJdCeFLHuiTc0lwk5A+afSiiwRZJeG9FqrLf+WKKsVOAZZ34YHcCygf2eWE1W
ghiwfC/F8adnOQpq9mWQaHQs9YKwpnzFXqXn4/NnoF1RKvTStphvXuHFlT2DLU3P
AHOy1w5P3wu61zaUDNwUuizCFYNu+HwPZTd+nMSYQ5+dM7Ftr0yKjYUoNj71eEpn
ycSrmURPnBHXD3Qpp0wnoRJ5Sx+W3z5LbbArBD6tSK9etge748cGNKpQUtZx/uHk
qiO64dISdbicz5+DPB8aILciTKL2u/39JgQ9Yke8jLHX2t1mOyniLu4ouqtV3yT9
ZEuhJNOx956bWa6eL6RbB+XU7NtkxWTB5YsOuZ14Kd+5mjJC7wO842e4FgM3h55k
79NAX+60I6FEkgPZp4RArbPDwZasdgklBifN7moVU4glSjjTBfdlURnVHJuejfXs
bwY1JD+T7Ch9Q8UrfBQdUj6MBSkOBbDmZtDmCbrJlW6z3p4Us6RWhvo1ULNgeRMe
G4cvbB/dSnS7Bo7TNTI9G4luQfOxf4gB12cCgz+RX2/3Fw5DIbtQWdkUWNbkB6zQ
8XWMjl0ieZf8k7Vj4rNQ3rc5pNPh98CBQqAzl/VKRqAvWhXc2V7osnNNRWnpG8us
Vm85DJgRWCyGTyMiO/a9Tg8k77xzr3C+QuIv9nRQ4N9nKACzGlCA77U2J/SH+C9Q
I65M8ZNAATokTPnNxsCrqy0pcgnmqB70hDtugsCJBqZ1OLK6OSOsdks6ETtb8/3r
Gl84bygk3U4+yaUTQlu1gGER6vg7aN/eI1Pi8+JANfMILl3tW6ya88m2ouEDq4bj
RH1SEoAwycSlzPmB9z24t2lLJSTBFnt9fhpi1pulybCmnGhxia5tOcVimtIHOaBJ
Ti3Hh5LZq3fiQL8cpVtUWciw+YeNIKASQO/DCqU7Te925p9EvhKgaUY2s0tw2ELD
KZVmAr99Yq4h5ay+cYNEdIqTjC9aGjiA+RV24nE2M9CDnH+jTK3fGFnoPDT10cSP
aRueWSPL8DqAEyHSCy5s2d/oIWUyxeodOE/t+vJ7ms/jMP9uVOXB2rxR3No7u8Qg
nNJUyG7pAxtGeSzr9qx0Jt1svgINQI/4pCy3B/J/Gvwn+dPb78WXzc8HCvjPHTfO
7VCOThFs/KcyHrdwiEhdezwmy5Vzkj8n27SYt+aNLugDDDIL6IFreLxgHIUZsyp1
VgN8/gkxAwIXXqi6EnqGJ3E2TjxZ7GlvFK3I9SfmK7N3UOPFtB2Fobusp+2IEuht
03ewDMw4+YDgixwOLAl0aOsbyWnpm6Tb7Mfu78Nvt3xYJlu9WT1hK/S/V7hy9EfU
hb4R0DiCiVtpKKqBYFhRyPdB787Gi45MRokXTcST7mZXZvU+lFcSsIYXSHT25Kii
1BFQWtiN7hZERrJJ/E9jrVxCp5tXYff4/dfJ15FJsIyUtuyF0xFDvbLm39B8W9b0
itcqQgkznPEya1tetTd/dyvnn7CwOosSpNVpzaYRQFmOpsY2f7gj1w8NYd79tiPJ
NBZIH5RD7ZWu3691iiLowyIxLv7V04pIz0RRjYhVJPCMe9RdIWnaU7a5/HS40tfN
vaD52IseOrbVMkAD0lR2Mt0vNDXwoxONpFu8Hmb+/Xg0/fthwZDVm3itKExDPZfp
iXyeR89hAumZp33R9z4Ua4lZkHbB+wEUQibkbVOQ7OT7vP6tJeoNMOMPFq2K78vG
tBiaivAO/L28e7Cc5cuHKlvGJCWr1X5WteU+PisiQimlf8HhA9Lozqfg9IzE9iaA
qE4QKjG7GHst+DGmsChHgezesUnuI1LAi//SVJR9WmdGJ7ibicot9ceBxrCHfAir
iBfX/fLjUYAXi4XL5HociZFElNFYAmaC2GeHvgL4KzbLaF0YSBTPHvL2L5hsjdYT
60vIMS9Wmi9GNYOX3LMw0CTfsoMS1XwIIX2u4F9ZblLafEhiao7Ya3OwEfIYcd+m
6o5KpxvJZ/j5iwiyePe6OBuyXjHxo+QJLtIy03I+F7AAVuLa0h2ToktPIL7oMmmm
I3mc38MGd05DYL7B2m6PYeO3IKiBAG68uZLiEHGB8NaI9/P/q5bliRT3bEJrBBAV
FBmtksHdk2poPvXbGcvX/INwTVLHFDLRhoRfBF799Go=
`protect END_PROTECTED
