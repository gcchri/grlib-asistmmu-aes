`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FlvDDB/EecwDrYl/VekE0jem3S8bUvlfJP9szLiT+/F6xk/WMf3JbqFfSMjiNthL
w17+jQ/qFrCyuiUW1YU/KTW3/5SbGgQdfHUhlVryyA6WghBMn4UGfVqFPXZGnCWS
OPuQeTywFyIrxbK5PYH2q5JoIL/9b3YnXxsosZ/A65viwMScgieJOpfbDl5zt0dU
e7KjHV0HCDbOSEEntaczK7VYfQQVa2SCBzjj0XJPMJsRBMdxRPrMZnFNXPBjwYBt
I7vSL0X7/v8Y5wEjIUiOySmFjRyd5Kpd1lg+L1x3gXnLFNeHFan7D3VUjeoe+HrG
uJ4AquKsuNdABlbWrsJsUEO4Fl+C6mLRgCxJ9Aso1OrR2ZuaOVnsIBuwhkiFmiw8
sbQRx48s91xkqAskXfDd3RWv7GReglej/qQX+paq+5JAJzHcKznJunbI2yx+oNRN
w3WWsRWt3NzeQP4Qcc2/WpfjzcGWeyr+Xj8h7q6xHnMYmV42Ph9OisYYnhk/3TeV
LT0hE+ajrE9qtyMDcd2zsWywnRmuu/nAx/18a1HaMghZBzznr+Vr8zrMlOmGiiY2
BEF921FkLSk/WbpLB9mMN8m3KadF1Sm8ckEGxkCFcqZyPIvj/C9kAnTJxj98tFde
RZHjVAaTNGIh09FZ0Z6292JVqX9eoEiKgab7y7TRUb+tKtAnXxIIY6OD0+XJAv6V
q2oCvmiNC/NEIM97/IY7Nzclmulk5brc4rPhdEYLQMT2NNl97bmhzXbS/0Oy0nMH
XpT25mLzeoK8K01OV4/8CJCTIpm/EGlsGRFqhvHtJsU4vwxI0JdnreXcqgHFxW/v
oXLmRoOz5rWRcySkub4xRxviP08hGvbPsOC/kvqr6OCYhMUZyEdmwYYUyYv+5lWk
1VUL3+4Qv6l+AHOjoosthG3fhFlgXS12JH8qcOAgzFJuKXPAJN4mOeRY2ZV2hi8d
AE8aDZjqgCL2U9f08kg2tysTPymoyivH4TUxt0VO+PVLhrDKBkoqDWWrfmjwIz4z
XqBp/6DUDzeL9eJr7ck1EVedzHhWwLXN1KQneri22IDISfDoofUJJd0+hL+PbtIV
2mFEevYByqv1nJZgkq0yuAi126N3JpFQU1FxMJFtyb61sXAkPz+Lb+5iZ4E+yYdY
HxSsDiRDlGzRJMoXEjAYTA/WgG24UxOq+K+dKzG0LmasEmT/SSBzmBJfeafZeuEu
lVfhNqwsVguhMmb0Ztivo8JazCejpK0qLF5eQLEsGab+C+uLiLVNN1qklZkP9qZr
5+YwLoNE9btP3Gx2kvfMQQBxbiJ/mgeTZf0LzwZQwdgUxZqht1b0K/Hxnl0VCziJ
pQsqxVREk0yG4EbJbsjNHmlRjrjz5L1w0D6qIt4vRlS8HWRp22Zt8HBenxbS2hgy
lrePVRegCYRIZsDpvVKjZo90B/nKvx1W46/ia9ohpFlI000D4Z8DyCgU+o+nUcBH
+2plrWdsU7dAw8YnuixGctdF97Uyg/KuwMZmWzKOCSS+xc0F4n3Gd8LcS/ywexFJ
N+6m4pCCkpAypiLiDH8UFoevAkCSr0K/bPfiMp3uT3JM4PJJv+fi1sY0OMv1kJk0
m//i3tupINPOQyB0gG48hHgsS7tE6TqxYP8pPPAZLJOmXXns40NVg1T7YaE2tXET
twKthgFEC73+WwCMyYLB2OmpQMDU1eVhchZMXlzI8DqRq9HRKdLT57FtF1zt8pIw
B466wMmBGe0GthOwWCiZ9HsCqXHFp048mRpGPpCpkN2evNW7pyTccXLfFuweORlB
ivObrKsTF9B8G0nMHxhoxPLdTCxfBxx+CxKFmXc/wTxtPRS8WIykjgnk1C3BmYea
3RgJJ4Q76v9ojZYtFUstK+LoAhz5poVjGJDs0J9IJT1cfV5TYfoUVEph1J82yhxm
mbCL3UIPh2pe1e4PzzoM8NvL3vUn+zRgEDdsJleMMk9h8dEE6XL2ChDgrB1cKLuh
Fj+UddM4kYRvETkM9ibXhUPyS6ZgQf/WrWm8y7qsHC5PpTDe735bFTm09nURXwog
h1rWqxrYaX+KSBtKAkY5FTH0e6jjaFJGjriLa98hn8dfnrgOlGKSu9EMkPrso2I9
jaI0/BLICXQHTXvtm6a/eKeV+sgAX2E35xhrDQzh3WOBTfMl0zkwFCREaGu57KAz
BRZ4yZmfoNexmcvS4Kvy1+0o23YMferY5v3D2JwO6tnukFF0xf7EP92KJ3gMzZ3u
6IjH8xQmeEOj28qdnUaIzhAnpr21fAvdZwJyn4xBvxLWPuSJ4ffPvN08JK5bSieN
OKqjOZAXWfltdRToPtnDKT4lte41Od/ZoHAmFzdq7D2YGCAoPioGmtaRyGId9sad
rY9baCP5TaAbmZDh8PDSZzVTF+RP/psfjoEK2/mc+cc604jVgy/oMeO+Om8vBWjG
u/MU+1AtBfLNvN+Nkyjy0MqgDwEKhYJDyDBoo8FO2DxHvOJNKISxiNnX5OtoZHgy
P0CobmFGKLnuNjIYTeRcfu+sLK6ypWfptBi4ouoYSGGbYJkEV3lWy13Cu5SaX2nA
4g/adZIB4BPjTpFpmvWL+NDdTPryPaBQXuEr2FIHKfSeBjiaBBi1LpShqDNLBmSu
T/BmArI1upY8jRUKXHcdg6lA6bzqQ5LmaxtHskRKu1/G6t6ILh+I0ucY4PmJldfr
gDgRJojCvHSofDqL29g4avUXx4gaSkaWOUn8hAu0UPz0I+2Uipe+F9Er/2M9oJti
+8i5lPqA2GJ6oFZuISdet48MgMgpNQpD9Mi037J13D5v0In40mR3hpVnKjLsA+t+
kN/Z/zmka8u2KpC8AJE9sMC8aRY5Mm9ETWatJSihZgs31X/jHdkwsU9BB2XL2YMb
kV+e2/01C0W1j9Oo28BSsMroPnO4emK6P1SNUcc9Bv+ELzGccYtbA5ViE/GkWbDH
VSy+7HhxdV/nQDVYNjVDNZCpwPtZes5J83tN+sBuPfyTx/Z/I6xEEvh3aSGA9ylI
/HMXv+DomE1OnbrGOQHDrsKK+Pttgd7rW6M5wOgPed449e7klGzXo3rAGa6XuQSo
VyOdBrXUt+eKy/41T90U9QBY71JOmK4hYSinaFr6Q1lHLs8bbNgXcfrLND39+LX6
VseHnZ/9g0clFFIrjGqyzAnjfOSPpjPUQEQ5BGeCcoQzkfi3L5s4720HMX04wzxc
/8QpvZyqH083iYoSq7YnCaejGdhCrD1ajLSjINiQEf6qmMk+8E3vaNO4oUyZ780+
Zvrsl2c102ZepY/L/Fs+ncTtWyhCv16UpnI8zkeiy5wNgu5dG8lIsyVESuIum8Xr
i8OuEXl5tel3P/Wi0v0rgJPwSPrgqe2rpI+fciHGfXkbu8DqieX4xfqsiUKsDpMo
Gq/XbmG1iqhG0sUuS+EmZwpACBq2FZ9vq+IEZY0SphP3Y4kRIAPyZNcbDzMHNONQ
tBEQkChoLZntZ4FmLpN+ssLr4km/nPnM4yYK1XGnBFITJVcQe+Mnw0l1GYwPwkwI
/Hgsdg4p8PSrln4nQ/E+0s31XA6P2VhiWJkKw/q79OI9VIFbdx4cjtuPd2diLZgX
yX1cQCfUse40+CK8in2vozDOSq14Bm4aMq0ACNVTWQveQ599zcYwE2DQPaq4awqU
6f8A+MoHfkCdo4dMqh+0K7PCH6g2oBHHo+52UaPY2UYItk14M75f/WsEQprryh7b
ux12zRNXeJEJsKHZGG4LtZaFcS0RF1pDlx9IpQA8HCEiR0f1NxoRcb7GdOhCeKLK
yfepT/xj/amx203PbmYsVdUAg20W2LchLEfPZX6jiPMOVDMD/3jeGnQ+cicB3EJq
igBfGxobzU0+KCIpd9nD5zmcRfloxBB7qo2pMYquBcLGPJgXpA89zdj0yOCd45+2
vyxbOoQZgO5SKGJj15SAfJlyz7V9/nK/J3BU4TmyoUunxSxkpwHYTkSZ1R3l1m6b
qnjNTbTt52iYWWdaHLhBzASvtzFES36QCe98TPJXNiVk2watoPw3qCjqDK4WYJHB
rjzwvJTu8ZGCi/aro5aXb4H+JD+KL6tq0Aq5LAxQrP1ZPQEUWyFApgcza0xj1m4X
LArc5MnCKCAuEHt1Dh9HPQ7GDLVuO075khAkrgy5qA23hbSjHkBzidvB/qZWAZ62
PJznhuEw0qF63SdLvY9Rt62sdDcg2BiaQ8ImExK0REJkERJNg26xrr5eSNP/2Bsz
8DApSd5+YV//qX6A0buIAp0cLC+YiHZCxkNSbIMg10/l5qw7jiKDu2FThsENgTqm
G0rfAKGe3kJKvpTf5+3YO6xjQnVNL3irjbpU7N6NOUMCzY2gyo7gpeRh+mta3zVD
2q8G4rITagoNXcqB5/T3h6JKpMX93peSmNK1Tt1FgaqedG29fkWWmdirzJujxIjp
0BB0uwLA+Eo9I7C9zwrixRsZ+ljy4U58evCSdbQ5uEOug62pJ44knT/3KLwySHYn
GUP7nu1ELrUHIwyuR88Ef6WC926P8e/DTQyDInqNcUEQs/rleeFCcKDBSbsrCNhu
kCw3R/5LbykTr8P61CORDgihcn7cvf3k/QxIy7fIsdZdTO2JEaTTyqMzfbQFBkj3
yzeE7SdflguiHQqt68oVhN1qQedw1iD5uFnf2F1In0xzEdNv3u6zTr1UsrRA/ObH
M+2LxN59hCkY5BHNQdRpfssRljXh1GcSVTZAVuQEsigsdGbt+YbnRdJX+iu0qs4T
tJFCCFTfVH3alc9avM9kmSMw3mVDYxBNqxD6LDsVuH8ii9ErOHcUd/uTH+5Etrrc
QEAlbQbJr8gD20pr3U9gROetPvpMLHm4fTrjR2gfh8jPs5GvuOMQoZcjbl9buxII
kUMvBUHDYwCU0iZ79bhdl8sysSRyJ3kXGisszMMMTDFjp2M32fUE9UTZ0RhWBsav
sV3tV03ES4RQuzMjSZc5Dzh8NU2+aN8MBFY7vR9RUT7LM3bJyRa2LjRW/SNeD5iY
s1STxIy+tqPSRHTzfSqlvxkMc/gPflkySTEJ2LZP6i6GoWySN8710EfwrIuSlSa0
j2BmxUs/oVi5m7zU/yc3y7vMlILJ1nxdsO0ROK1Ju+Fx7ZxHbpXydrkC0nnTTVi1
kFFka5pGuXDN9ugq71N3riPd9pXd5cyhsO1TDm/imvkB3gYCA2V3O9x2m/t1izfr
IoXULo1NnhDobltpz0CDX/LtUhKn2ikrUF4mbvsd+aes8FjcErqjAdXZILgefkuC
sKVjaAdaUonbEO0hyJtEut5OHYspTFqECioQrfIBvuUeqJ8mbryMaC6s1C1hhjpu
JEbFMrNWXGCHosXuZcfVEPnAbvndlv2FTsSS4JNr02Qv+TD4SudFw5D//GhSOwmW
xTmTI6TekN9Cle6YJMNG4qY6ItyWdQZZv5dKoLTxU+XGjWvvPmVwz4OX1Pd6hPE1
X0I276J3TP1KGTtOztBn5qD6xAFz8WcbubD15CQiFfq+wQdPgASH32EipGnvTp/r
dn5BDWhsocbVmgoqxewW3R4N3ogeXdnSG1P4qbbn0WMnQseNq3G1IbUxzWDCRm62
TfZjsNI7q5QyFE/+vfi7CRUTrFueUIaMzoIeqsCHmRxuMhr1JTB3ywUXTh5dlVSI
ZyhOSi+mhATPbajn95QSTXrAI0rEeTKIGLOmjtjHqHZ17enidc1wtuWrGLYjidbj
O4+ERniJdIwy8Bxk+7BpLYN699xQOkoA/0rAVZWilXS+fM2MXfNLef8fC5e+nRRp
fY54cc9HCJzvEYypso1k+IZdi2vdZDpUZDdPWZahq+mW9OgET5qtg+ac6/1fObVJ
Qrt3K6Csq2BH9NYQi5hhIA++whweEY/3JHgqL3kHZ6qT6iO2vkFrEqOsKkcCXv2p
ekqiG6OiNAjOoKoj5ohapyFh7lO6sKLCfCRr0UGOK31xH5rg/e+edeO4T0ytQ8ns
HKT9v+O6KI99gLmgaNDfoNaYRFv9pj2RJwWU7M2e6TQR0qb6HFdt+zu4edpsvRaV
voOmGIKAbL5ee9Pq3aLLTNeOgKUDr6pi06MwYjKqgZsnZDQLWDy/ENcXveNEeNGO
1IVuwga2c6Eh+auD+rQ7ZmofCL3iPFxkbLEzW6Gx+T3jUdoDE8TJ7GqYk47ARrUy
9rlttvRf4NoXCctTpmMpIEMyOQFBTYJvgQhSBf2yonJvHiSdN6/lRhFCtC+BwmkU
3RVmABJx8IJAyppDtlvmxxQgMJt/nOawkQ6DBfvqcjReg5qsiGArpMmWGKpZ3FJE
4nhNiO4TdXZuCaneGhQp7cn2uLQIM8c1LDd/+FuTy2WUwHDrM08rztCgj2I811NC
5+mE+UdVFEV8RRfKagzqCZXWDPajQXS3zN9dRgH7M7tVBm3dCTzPI4T5aBpVD4tA
Rho64VO4ZKQxv8uxDD+Cyap12XfeJ1MGmwzpLDk/EoUjC4tvMDas3DbeB1rUHoOz
+zVibI9f2m1zF6u9Z2PXsbvrUioC8b7qGtcpHPu9sqxnUJuz83yrPbqns7L/Qxql
VE8E49v8/My0IEsxB3DtITK0OpPupKbH5n/ravuBi1EmFDuEJKsCA7wvbCSJ8PcH
uXbDFYbV3o2EdEDOeiK593spHnWQwBp5RwDI90l+tdXvmUc/cjxUT2Doz4Lbaajl
tI31SacNqmqATQkoROBlHKJ030oSgRbkmhSPY2Q63BwN3dSLlrKH3bCfMESaNKuT
NBvtZPcd38vrttv51eA8NeLH1MxiSYwBw6DOKCvQeoX57YH9gsqjJkShwyske3FK
vbSnwLDBi73w4xqNzveN6J7sKsAiR/RlaA+t4EqT64T3IM4VbGcjwQSc52dA92WD
+A3VG3pc4YX3DMFSa9wM8diE29nq7aR5JdwsL/1I6wZTJo0aEZGjtlHRYyFbWZU+
qiA6kYOx9xS5MSq4tK2ipORBGzyi4A7ykqnkWIKPHMOceeBrnybX+wZ6xBtPTH4H
gMAW/VwxzBW2o59yZ4NxXAETn2l67R84YNhOFwFICMVer2siHkuu4JyfcyZF7VzS
PNVR4lWVnpcRM94pYSf342h1iztgNDbm7GPPw8h7JuAzowrwUm7URKqfBk9qoRDl
+B76/qmGIKgCYiEF/GBeMi9JIemrjzkGFNuq6iHzWYHSdQTXDb8ZUiLnwhegSd/t
NCVqdmIMAkn5iXTkuNA+siu2ua3Ea3bz47Ad8DpDeGTlMFE6OGjuf9kUQhtYig57
Wb6CcTZWm3hX2o+ewxWjaYdKr+iOJ0tAkhcO80wd35FM9SRES4TNSMOgxG09b26Y
PYneElMqv8Xy4Uu+Q2DKNWjYztqm6ECJ+VScMfEB8DlpuQhcNZvkJQOuDbR4L0/t
y9QKsLm4LwgurEBf9+DvCSJZBVPLqtenIHoRGMRnmC7s7eSVwlScNhH9qn/COl9Z
n78rIBXCxdcdT05nKAthRDC4z+UrBg7pk5V3avLS/HAhK1qSS5fOJBs0JhuoRrc9
VCMVnLkJ/xtLT+t3jiWE3jawp0zOCihyJdLDAumT0CJlc/6Jg1jgD1a+qzNJk5L8
rnq2QMn2iN7rgCM43LLEAUGTN9joB31SbpGD81awmw+xk1y1FTlR7WfZ8arxT6iZ
96jqh9ENKXbV68CNzGEGk8i5OsfM2uVCXGWh4vvTedaV48SxYL1p/wskrd0O/nii
3gc8qooGYXhMEnn/Z24C+QKeOwKhISsct986T0B9jtUUA7TaHM9jLzqcxWC0+H+N
iUtIY0VQX7T+8v5l2CxTfvbVnEnEHKrTt3CwWPRdaEN/jCwLCA1NwJoRGPpGl3tt
Z3o1jYGg3XlwXaDj/MSdt63RNXKJXJP+T0dDoLK1ukPY4Ew445x9RxBgBGCZYXyn
B/8r+Nz+vnwyBsgkaLo0f0UE0SpwbCHBpd0z9Uu1NhYWB2SLkyLbWCmmmOdnDXWP
wHIgLJFsrBLGvJZVbTMV94QjXOMR67M51su3eH9ND/gjLPDdyGEIDfsciSkraAM4
VZ6Z8P7v3LqJwlEJSQKu0XDRNnvBJEjq1Hcbwm4rWxDPZGlraYzUyfTkIxMG7Wav
+0mVbcZ+Aj0kI2qPxUNlBcOC5+BpyCq6lXGs4OBogO3pi1NHLj/+aETEosj1YBUO
RWQkYEBxyTSDFcEKZIEYMHrUB1upqnF0dRcjAGeLXuwdqM60qAUZwZYH+JrucaGV
nIpREXonAkQKFnAl1KckLlTmJbP4uP/YI3LFdCWtnAN91VQI1q5LeL6vz39Endq6
4FK2PmG8oYmy1xPYKiCl1lHyOtzZBDEN02mSazbMowGqfa/TUs9JqnPFTdhrM4f+
vy0oDUzQGQGf6RwNjYIy3nD6p+j0/6j8mU3i9zFYQhe+/JZgBT3rAKGXvs6MXzjs
SS2PjeeZx1AuboQTwqliobkattHV5FNfZb+GCmy5nZK1B0oCFdEs3LGMxCgrOqnI
vo/mml862yMxNUa5TOgBBdTUP1+mIa1F53C7zdK6pqKwMc9/f6nNmEUdj3tS/XD0
QrffYrHKvXlFXyRWxVPmRL4WLZ/uwgUuHGvFQIiLyUFuW5mcqO1M+XMxaBLOZEro
15yiWbczrH313h4GLmix2I7jlmbDknvOneBRWi8mH70JbIeoY/I7dijC6+ZBhSLX
NEViqK786rqFXBx52R89aw3Nx4sr4680BCHKIVuPXed5iWw87tiM8juMpu9mloF9
Bi3KbSZnTXRaRHbhUj+O5kzfB1mw36TNRuDuXPoXeIRc08P5Ht9owwaOYAp/+QSb
iVbqop1LSdGVEExQ3TWNYxAmOoUcxfp+StiVWGiC/DTuQy6V9rQ/w4oSQNpON/Rp
osqbvTchmbM7QnS7gNCi2dkVkNOq4uzQ9+t1+37LZL6NcEPWZIqX1NGnItmRymNz
PvxCaqeqi8fssegRnOfkG51y8cODNXkBK7gyJRR/mqlGucN18S61thRUfZXD4KB1
pdzmRWx7RTQR0QrBIiHH0co/pSA4aBgLx3azMI0o6ZXjbMG4RZgm1+RNmjDtO6Fh
8loiSDvqNQcvr6uFPQcyrciEfYIWwVkkJLoc1OSCraTp9Mq/EZ35VVw4jr5J0P76
owOTU7O3+h63avOn8ZI8E5iD9HgcuM/54ZZChasgFH8d8JUxNTODuRt65amvODpN
asozZYzidnWPk6ToUDn+ZjVD3906y9ZUClu4kEpqWhMANDOQy4rZNRnq4BJGtM3M
PsVOeY/2KLEIjURqINbbj/fI8xDcQkahyJOOZmeix4horyNldJN9K0ziYskEvUnT
Mdq59FS00NnVqfSJ3V1JwExmU59XYMslZwMLIhgOw0X9tPowqTb7kkzMSrtfgC5i
Z2udtTw3ThW7K2ueKaa+k/BKJsErvTADJMD831UA36sYPjU++BdLs5FYS+ob+BuX
4QVug9QHP3wVzpzNIAwYptsYki3/eLgcs5lKlZNd8OCKkH8TKLboW5CK781G5yL0
qJFedOPWGzT+wsQa5ZTmBCbz30sytO4chHqdF24RWa+M2Nf05s/1dO2PPXUfvzRY
FmNi4p+1Rhv/+sGF4cjLL+SqsdQQbjgnAEwDRI+sfWV5l6C68uSTtizSwd2naGDA
rNZtZTcAxIHaGkwH9yJx1Hs6bURe7WoTJtFX+NDvHar9sWXhSgKtwqhGygzhnBD/
Vl81SK3JRTMIOcfwxM2gRIBiNoE2x2URbDsjblUA2ms2hogw1RqIw2cNp/HWW+CR
2TXK+ZAX6a2lWwn7a9FONEDeFN8anr9gXOB+/nZlqBHuT5RPC3ZpaBDOGO5yxx38
cG/lJ4e9cshsKi8NCq+kYXVVknXGEI1L9vRBkxW42r+g4U/xo9DljBHgWkXeCz3N
Gu9M9LyUshnMhXI5dfHlpuAJpNdQZktuzcq/4JG+VE95CkN+pH60+GPw6Z5pUgg6
Hn2c20Lsendc2LpYoUFfbNEcqw/ueKZ0ILHHtFae+HjHXQimmavPd3LP0c3/BEZz
JmuCPcGH57PA91185mLDn5aD/lY6B2Vcm2sNBC+Pt7zRupgVw9S4xPTkLfdQDLSe
nBV+RvLfmltPv4SAVK7VUyEXj7e5k1VpvHlmGdoIVe3Ix4ygUSvZRYu1jaSQcqKl
Eygk6mmCd65oO+xok4+CLwj4NfbGYYjqrBS9aJ/CkVopmqSkxCC0TsOZid3aZFha
83BX8nLHTbQholaLXI21WeYrfHir4RAZphLn20dHOt9T+NRZZd5J6ot0ArhMIGN4
4nPvSbx5ddxFtwkKes+8NQZi0VGGPJHkuV+MKbHq+nHfu2mZ/xSSgMAO4XLZZZPx
v1UKDF0FsktB42RhZexaq4WFU/V3APcgNcM/KHriTprgDf/7UlsQ4t5WAT3h9h0c
p4RacfNnSLEAX3PFa/LOxxRT4sh0dIfSm3vcnNh7tc7MVpo1dOoZfP+ic/W7gTig
XNtiOmRZxiMFNynm9U7Jk6akKlc3d0Bh/Kyxe568mGWSeDREpvAbcn8L/hozlNJ/
ahaTqZWJh/Hh/OVFEssqhXOsJgGaiXZ4OrnIRGcEQbMpZR3oSbrZqeZVZ/oQE1Sh
T0OIAdaIOMMDvg6AOsVkEriCO8KBu40c4bnOylmZjG292WnRUnIX7PGp1JMEGuze
z1kuiwLirtpvEA26QlpXX6sJkxpl/o/K5qrKwDCMCHmN7RE8oMlRlDCIHWrZQUz9
xoUXH8snkryJVmsfZ7T71rmg9hYX1WwdbOvpA+YP+4j6PbKzUwEDyRVuJQ9eLK3S
uF2PEMq9KuJuoeZLYSTmCSPYfJsW47atIe42SUKrYvDGogf05b2QxvXLemwLJkuu
6JRD0XGb/q4MVcVsNeeWo3bdfXZl2KJd75LXOLhjqOO9NPKr0/9IXLWIBRnPUHi9
bBJCBXFMhMfgVSO8IFsmK/pkXr3crE8UFR8ODkeL+MRe8XUNokHNV6j311fByrLt
1d5T0F1IPKAulm3ChnqASokPt14b112bQFY8UIwZ5BbOwkmq4Hm4xzssrHZzWQzt
8PATn4fkIhIAtUaFlzIdfe52sp8myM8q/UeNsEqQjEM1wl9FDsVzGam96AOPMEUQ
9M3XdmpHDEhUL2E98Rcu+4tZXGrPHqZUk3dTlsYWMXHkiXTmTEnGQUtVtYUVG9o4
Xxg4RKRTJ+wo8RNvrBekIZ7QVSjJBiJbqrqh72SJmBSMo2gos0JXEygsJcGGi/TQ
RhfnnMsR5TeJSxssrx8Sr3VSdbRjaPr1FonrtVZKkR93uzE2le2Kv3wEVcYOJ9mI
Ihu+bkB++JvrF1vaCq+61rDKDMxlMEHo+qC6xCrI6hQUvCAjkJOm3mDDWNSLDNTT
bquDiuir5ktpqIkUp0jwn93pSfSGZ6mcGeNvjc71kSFMUZUHDhuisSxrGqU+Tbep
6oPhFRbjXnMuQ+4xPXW0/PqpNdBS9dv2iA5RulkRpwSCnW7/GttMoTPxUGmMjsLC
5atPfn2r1uqMDPiz6msF06NY7GAGLS7OmiMYHDSSt6iwrTbuUObvqt/jlVmaDPUI
Kj6aS6D/PaGaTg8MrAU5htmI++aIlZX7e1Yech3Gjy3nAJBUYAwUY6DptIOA8EEI
xstY+Uo/76iYHsT3GgIGEXsKKltUH39RUf7v1PSWpDHSeBYK5R0NKLnYeuEyCrc1
3kU8tYBBze3AmPtewJCJrwhvsNfts+Cy6zODWvefJx9kOqWGzcT7+s+Qpy181nSA
OG8TtFpm2hwrkINjC+sEIe/iDX1L33xl+UTs6wNiLd66IcQS8z/WeXvSh/zO2rIG
Ez94SLExLW/83FGotbd0oCWgJRJYvXfMYQ/s10etBp+7Af/tKOJWUSdWLqE+wTyc
PPSzOdA4GW2Dx1LGTXL9xt2S8v+YZvqterl0ScuasBeagL389RLRoIaE0w7lkqzq
2fDIgx+LBCo5nX4Bvf+Q29L9FBZ0RDk1jgDVKzxtZtaSDcPloDtFLM0i8BCJtxyM
KDbbr+S0x1328Q/6jbpqz8efRFr0nfI6ps7FEMZgzVkK3+qNY3hMNX6i28bdmO1W
wxchO1XD+pkgjTiSF7OnmcbDr8jc5RU3JMs2+Joh3rnYMqBkOS1h2VVkHUGv4TG7
2q+DD2bWHNxwT/tircHPn3s/XVybniWV2P/3idj1e/bWWsLrtcSIM+yjOMFHAUEZ
Z/NOcT9631CuzclVW0bdsVu67d/HO7L9KnSw2SLSiKFmGMkgEo7nnNtRp2+xJcTC
RYGvED+6PThKB9lom8Q2s2tE9CzXLCYcTmhQMln/XRB6LZBdC+LvcI450di1cW+L
K0nUAwPEqUQWreocd8D3WWzxLmhqmXAl5wNqY8F+B8p7KBFMKQ5PUe65VIP/Y2sY
xjvV2y49KD/EfyPplGAnsa1PTKNjEMbanRwmYqwJnxd+119tKet61QE1qG+UHGT9
oziMe34MXEgUYyMmj+q4HlnZ+DBi3wF+Nf3/2Pw5pjYuZH7jqgi/Rlk3xOcYGXhp
RiBq4Dn4FJYgUt+dZGCPTU++k7Ha5Fg9LelwKLYnYKyCs8NgkAa7BYYsWwioHWo4
SnITf8UqwmxmNPFv+0l0b+XY4wR9LPMX20cBGpBzVjByuZivyB/Icr2XFDqTk73F
JOdTcWUd1IF67rfSBi0dBrXYyuzGi3yzqmnJWuNbnP8Qg/JVYAVoefcesipdFtt+
yGbIDTrO2SPuERjnabdYUYBcvqT/xgHrKQCdHWrz8pa0gLKsyiYNW4vObGq7D9ja
NtE4RTENmDVc6aAi8BO3Y+0xS6eMSWjmmBisdZPcMjWt0WI35mPvzXutCsyTZAJg
gPJUgkH/BxWpwND3cWFnn17oRRXpQ1qfbFgPoJaWjP7uIQbRt0rU6BIbX/P2fqmH
QSnYtrPOonPalYt4MEW43bd2nc9R7t1YeI1kmMeio6artwqaFjkxKam+RaHv/iZw
uPHQ6WgVDJhLyl3/nfF7xzbpnXF9SKL6BjNvP+H85bmz7rA5pQA6pVBEYuuuQ9G2
dpF6f/QrHidEC0tDWpe/KRCgziVfyIlVqan+AzTMDmQfxwKhBdx0lYMMvaZlHEbR
HkCXKauqz/6v25AP5R4ekJVPr2Zdn+MOdtOL6/KkdKRfZ+jVK/y1HCFbdnD6wGGa
pv7gFrd3+5xdFHp+9Q6I9TYnv6Vpg98Oo18hmnk+GkKjjOrmhHOPAoovSgxIQ/RU
I55fMZ9559XPHYEym0XaYwdAB8zXpXFuoMOZ5wH3BLAGFunITSIrgs/zlRKyUU+5
m/1MOkNNttC0pX4pgltoS82kDYWBaes1RUZ8RY//xarFQV5NouT1itJb1AjYaE9x
tn9kU6KH6rquRs1T9Q6mMFLEey/QkoN22WdPAbjh0RO03oqCYMBj3bfpVS+GfEbM
RSVDetPxpp6X3Hv1ENP57TWFVkPLd7JD6CrQ0z4ftqJoEhPW/Vtb0bMZyJrQ2gbW
PMuzF8vxnDkaUX1o2VB2OVLZriugsxRCKuq/1+V/Y6oFpLjkEcBkbmB9I5pdt5h/
+NsTdytuNxyuIHgJaQYIeOwdVC9DAG5zQLxyeLhJFz248oRr8bWKDi+e7APRP7LR
Q8LmTm0BagktJysSq772PdOdZNkSGOsG3523c31tBWt1HcdOSFNzQ2hNikrGT3Ax
8YgHWvciZfvb4NIjVGssxm9jjRfMppEsjt31ViRG+lX7FNQ3S2ErhbrmNSVH8pGc
dgX/lRm6wakeMGObt/3VMA==
`protect END_PROTECTED
