`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gv+e9FjEM7eHxtvKbrKukQyChjwFzNyIJOXM0CDbK4tqvHXrAZZ4FYehzTMfGo+y
SvBiSlLYUZKK1Xxi/2/LNMShKPnJhaPB2pZY+Dc18AZOQKDpcJnCC0KhaJRKIuDJ
IO4mUd2KCYQDcS1x4ZFxgmVQNr5JSEdtpFzutPOm/T+ENnGdr+wI2XKv5n6CfSP4
o+XOSclcGLo0jypt0w1/lH9ndqV3W6YvK+3Mj80h3NZCK/1G4RJr1cjdZSs4JGaN
1HZgxkdVxS/dBZOZ1/8wFdkPa2Jas4eg/LSe5YNw+do0hpaQIHH1YllS8TcedB51
+K1P+MllQsr8WxYQrNQdPQfsfQ2hffyOhlhjWDczNCZaORixQwEQz5OMq2KQiL9N
Q7sGLv8nuLu0d7jWdybNWwdVtAXoWd7mviAYg0J4ztUplRAGprNMnulm/xjVaEGY
BvszVbdiy6k8t478b14D738LfyQkHFRoEebFxkL8jh22Y/5ukSlJ7LB1cYWOG/tL
dsGWiUBD/K5cHCwHc8PGb3xWW4GvHYJekRv0+IZhACzJOEJA1pElFesXJWDUgK2H
D3/+rHH0PwMTN9AH14YOj6MegCkpodc1dOnGtjdiLrdlvsROWo2CiRLKouXccM//
E35AuIR6BIG3poTIwIoZt556QW6UyCk3Shtj5AczXbE=
`protect END_PROTECTED
