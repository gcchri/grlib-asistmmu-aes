`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjFEvPfNPW4SwCpNB+vfkmhG7GnlKSEwp9RcQvSscS4NYZ/3lVNktgBWj1vvkT3Z
J+ytUeQ2t5GArdTUA8fqFGgc/21/DLJptctO2TH0Le1EDhV4vZ8JMWDAMkGiSA6e
cRsPr03qVALVFztEpaDxlSRzks4w2yGNBf82xy6XozQeMCzWgZd/4MU/SHy2W4jk
ST3qiSQl3QtLLdDjXb233FeWQMeG30F5lm+mHfHXXwgaypOUIdemaij08I5BGvIc
WB0qbDo6gvsceahDgWxFMHNR9tiYEYpFFlhMjwGCv2qJDfQcAXjMeXzaoEmHHdxJ
WDCy9C7fIAukkxQ6vUag6M9tqmoa6+oZ/PKFw8pFnW34xyDHgFETiLRo8Vh0XM75
8xcOQzoc0b1Gb0zpfEUu6/TUMaXslQRdmZ4k2booiuKn4HMCAwZKaCndsgsC8zdJ
wRLtASZQSShXY9wOORdhNNHl3MCQrr6s/Fx8lcq9VX59prtShphtz/uZ2BktMPC9
ZqxDuXd4A++3TFUK0MbqG1Dtky29POTXgSMJuLj7cgV68w1dLlPfc3FwItkoSiwP
J97jrx+WZO/Q9ac8wL9Y6G7/77dmwT0p+wVLiw5tGDAXfoQx7C4npHh73nAJvExM
j2z36+V2lbKqARZ0FwvwAlZxCkTqNVbQ/gLdlXBp7x1rpcAViHfndl9q4oqg68pJ
Gtpx/QsoBlLlNH0TCaD+pf968HodVshesxAPzdU2UAv33Yd9IAI0VLPTIMbbLQYa
7aP/BzLIyKDKfbIeiu/ysEmXT9bATyUZVQHotQ0KMGNzP1cO33l5lcsjjLrrHpwr
4xktmI4PDCnQqsHJkV5jBDO1JFsjKPyq6/zCo8Oar60BCdoDvgj4HTf/TxtCbZW1
ur5AwRWaVrpWnU8KHFNHi36CZ/OxiN4wGcodCf2EyPgIVBQ3a/WPLhyoiRh4h14K
zjNuQcToOE/XIWVBXgMjfJCxr+vqBR+Ijjij+1tGzgY3N5QD8EDN3jS1C+oPhvPX
he++epu3nG5hpLiGZAOYzhxIkZQdCNmeIEY8XXy+ID68WSnRBiw/ILGW1H151jLB
9IixQ/zsAbhOyk+Vsb5HhLe4nQqxfMaiIMXdTW+9btyn9Sv5hEhKCii4O6BvcMLI
CYDe3aQBHz9iPG0fGE6hquGyNkBpkIMF8kGCTfZrZYbFQQSqt+L+Sqow7xynCVLZ
pv+hmsFcrRRdyMNPWJ46QjAMDXSMFv1rQlNjyHGFVtDIQ5gtwD/oUR5RXn8hU3G4
cz/HDRaxd0UG3yaluYBbzZqRLJ/Je6iy2GMS+WZ37XFbcfGQ3KQqFy8riRLP9v4z
P0vVuoICEjISa60ChzYqj+Zja8lTRorsMi7QrgPlJ0P37YnZRqmbOORAK/ogHmw9
NIivv7lBc0CgwcC4MEelDmw7OugEDhCsGRRA4KuoCJpSGq37yMhwY46PSlxkCZi8
V2xBjHTvRHX3D2dWtXmSwSMcIuw6aYh20tkESSZ5CQW1XEfo+Qjq9Ozrl9j4CnMQ
6CBf0MkwY7pbLXLWyc1Hi5uC5fqSlDGbRRwU/B6I7pUPOvkd4vARKwURSYPn+H19
AHcvl+aO6U+NMPt/GXo0nnB4JJyeNzcbcoyiZl6zGIkSSBxs8yd4RhshBBGIQP4z
3ja9t4USbMjYI6Z0bfZurxzNp2fHUnVsqb2n/N44LS5J/kQ8PAj6SyNb/LKj7cG0
O0jZQ8F0OCo0l0XVQznvhCrEtCIcFh8x5qaBMzN/Alc=
`protect END_PROTECTED
