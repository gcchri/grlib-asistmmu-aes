`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZnkt7esW5amG7HNOwKV861EW/PPdriJ5sRnsv+WBYpqTJ2n4Th4vnvLMWcWBi8a
kLsWjPgVZGwLzwngiBvo6zZcJGdm4za+G2Y4xn/lC/pSUQK7Te0sKUFJ6AaEEGw0
bYoSih95o8MYzWf3BV4L6RaJRulcgooDyvg2cE2xyV2K02QDf/WtCBCK9Cqd8CPY
WWfnmvY+tqYZ2/vcMoEtTESt5/nQEqtNcccJkqf/dlVhMhFerAGmi9bx5kwoGO40
fruNNFcsDLF3VbwxSeFzUmvqL9mt0GTcOS01B6n8c0cO3eaec37HHnKDYoiHmFuN
ZaVJOQV/NR5qQ7p/KQY0KGXtMpsXri6vOlQ+xFibedDniDzUQmtXJoWYLxfpa3Uf
cS6/750M92myuT1Pgn+IM5ViHN9BjeLWx48a7I9O6BcYKu7Ah4juPMP0JuBnKKBp
PteL9cEA+vJSkHPIqUaBklAX5IgdcGKQMfiPEXMk0Z7xJT+Vn+doyoTZewV6eXWe
/jdA26u+5yANsZ6vQcW5131O5kOze6t7cARrW5p3cj+DALs2Bfl4n1dSHco4Q8OG
TagTPLHeJ7SSvqwrfXQ21i2qfcqAsbv/mmSGze3MDN4KHfW/lSBjg7+Ka3zC/Chk
L/bOYSffCYAw3FUmYIQz2Q==
`protect END_PROTECTED
