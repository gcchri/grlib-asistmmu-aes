`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yi+OLm+NjBpKqkjM+n8qI58TzXCfmaFzu4ELE1ut6jh3gvJy1EIH9k0XQzILsNog
SegKmtZ13O7abb8OWOgEDgMWgZJ8rhCmJ8clgFkt0b71aoQPvq4yEwoty56xddSv
TrtvNL+MHI9Qg2RRnFANJqXhw5SsLkZKlDgvN+aJ2KeWmwAMIaniR4ejwcmM6aSP
2oOAtff5B8d7OldkZ1YMyhCvK2cx1nrYAJ+U9gjFwmheTsSCrbt6MqWBq0oaG6O1
fKpeHu5Hke9PkBts8KZrO/QPUFPfbhrtc4dXfhi/0W3yXU42Nw2bBLKGslXntRNq
RiZ5cp2Js7eIIBtvILTDFUuD4lvgsYVvgSLOWtEIfJP1RnrVx8JUXRbn3cd5E0fW
TcU9zfpyQTe9uF6u19RdDj4xnGULY0hLAp8p78nykoH9RE96Nje5zlYQ+aek0irn
FQDdI+XYVO2UxB9HFC2RhT7cMJIsF7NnJmDmYEaJbmwS0y/vybsR0N5dZbTnyFba
bJgOwsT95z8VFUKGzzfdXSoYGawWeL8O+/XPnGIKU2BT53MHQvXu297NddwANHqk
0x90UyQVsmI3/Tn3pAP7Zquc0Upl8dnQekpCwAunDYhpaCZBVNDLDIquH48/B+34
kszPEge7DaNdmke23s/f+JeumhHGy4tSRyLgr1rsufXo/FNERBxbW++Fko2B9eke
rxus6vqQZyagaicY4DdY8MjUwKr5LOXbYqhtiC+Vshw=
`protect END_PROTECTED
