`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
shWO7G4t8d8igCS14bJUP61LazrAj3v0VR/8hjWca9tRkCsTAWW8tOmBnAbWcee2
wQhIM0WQaboLwPd+Z1UzKLYeyzHfO32Pa8ItnjKqMZVaE8cv2nZLzijVaNEkVnPr
TKAkcG7l2ndrcIkpJ2FhHi7ujHA6Cjcr+1aL5v3py3YnAg0n++8Xrdeq1uXY1m8N
h9vkAiAuuSNxRltoMIa2FQJSm4cTKuciXVL4AekpHFFf7Tf0XdhTklD3krcN08AT
w3gO6uplkhfkanQbNypP7eDZpJ2J0WaRjaXmdbMJgqg=
`protect END_PROTECTED
