`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JEa5hBW9SBu03bSxovSIm/Yp/5yUWdXXm+SgU/SO7mF4xuDu22WRcq6S+5+sygA3
rAdDFcyw/XcfTiD09puf5Sk0ppcv59f3sYEmOeW96jXdCvuB9iUvrKmr/IkqazpF
gxSodueVl89Dv7KIYxFEJCYvTyj6WFlneRKZqhmS5JIcXCwR+H3zsUZr3I+H0e9V
zoukDsB3qNS3+OwckZixptavyr8qFr8/4MyMgnOIyx6HGzZPiVgpE5gdcnqnpgZy
vbF8mK8qUn5v0MrXuX9mjQ8EwKSUPeBnHat7VWhP4AhWf8rWTc+eEIiQCXU7swWs
pOffipIrBJR8SkV9ly0bG5lzD2wKSd6OcUIL9DAZvCe94cVcfbjU6eMlwtP+4niB
RTtvSYDLpzPkyKrMFsde9UfOA0okGI1U9t53D1VkL0g=
`protect END_PROTECTED
