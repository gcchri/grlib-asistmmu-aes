`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+jmCujQ4YXyr/mNVRvNEyGIjLpDLJzixRwtKx9tgcJ7NHuzx9RiYT7Wy5eCSkrJZ
Tpr6L/Xc9MtxEfsU6bu5i1mtrB8YXdx4FRxs0Ug4KoGUQ3r3X/lrFR2XI5Mirvyo
x2DJPD78r7qBStftAIUnTXDhVcW/OtmLyiv6IKkY8CKjrfGvj8Lm7u04k4yzHp+J
35h2hP5xVLqmziB+YSTYxX0GvYLBGOGf/8UiuBO+IC9qozJsD8UyJ6EmU8O/2/DD
JjtGmJ8wqEBnsknROEulid+XEVefGipOFIn10+YZo3/puEtxjkvjRrNAk5DOnRFY
GCeAQ1dc6aaCG/TNkdYfyxyonsfSteZDfRCS1fWhnEkkYSyiQ44vCTTuAjp9UIW6
USEUTrNIWpZRCi8Diubh4k+RH8KQwbRd1r+/oNb9YwN87dDkkPRQw75vsjy7Xu4/
0ZVpSi6eAewNje1tcK703h4N5E5qcOq0ILKCWIG2FdRJsiv9pi4p/0GjaIvdn4A4
`protect END_PROTECTED
