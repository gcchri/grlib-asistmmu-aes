`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwCMaSnKotqNxNZWoEegk0I1V8iGjzkfK8JRHXqtdKDDsJwoz5qaN+HolxkgFI8I
r1d+3OMVFWXpiNHxnhvp7suu6Umrr0g1gH/CGIXoealqN9t1JJEL7VtgWDkxk/h0
SwqcvwX8rbqd3PrwAimGdsfJ+4FAn9n2Rz3DfKF4eqT51qJMkWGQ2cz8SW8dj6OG
YfZGEyt4ojb1LVcTUNyHWIJcxlXW8zJp+M7J/0o8qMmIV/kg8RpWWkbo7Oo6tI0U
LVZQ2YcRNik/GnVixGIbj4yPg2LP/Mlr8OeeohTnuZ2BClrujsWyiMSY2cNjgslz
0lEu/WnfrN5iKIvZyfpGQboeAsx98ii3asPY/54vfe5UlC62ykeSfUVt8qRKhIYk
4GjyeORQr4m2BSW4B0qIN6Z0loZ9wwjyN/mMVp8gNE9/ca7nSbgqNmi9xhFabMDW
q/w9uLLNnCeHClUioUqI9nIRXbVO3EYesQ0G4WnbpEQB92NrskDKnXdRIR2aWNU1
WkjZKUSTz715SfmYtxz1XJF6pQpu725G744RbGdYCaYSCT2DgqOrrupEc0nQwDbx
DU2N6cBABV2MGx2qAzqx9qqO9ZVSaPG/ym4tWq/iNKCQzY6QMNWMx2EORK+JBzsl
6MvCzsoeh+obDg3X7HTLnlLFJX4rKKr1n+DaTKYEeAblfsudL1cY6B/9p1FnmiE8
8OvZz1G07Ay7yxBZ87rXiexoSZvdaZvePqXG4BC1EAgYHKtIAcVz1YGp42JQCQub
k5v815ZlA4IsyZEKuwGt0Q==
`protect END_PROTECTED
