`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ws68DnvclfvJDStDH0OnweM/5nPpFehfGi1YbJRtUEyohClbWhS4xZE5vQ2luW+t
juDMLasz7gZrcqn4YZQUW1BupHzD+EOT69m8oZ8+P1r/ByIfoAHCs/JMLyvtdhEo
kzStkQX9gMSeMtr9ntG5rOJE3s2ngz/be9xnCcGEC+k/Z9erk+v6xBTM4Mly0VN3
Y+Fr6cS8iCoR5SnhTnCoGNA3vZHvdaYVyvrBxfSOUIUtNKaWVnLOAu/LN3PnB5Ec
Tkd/AiVWJtxZvxt9FSy6jY88ZdrqBfMWYKGiK495xBzsXCJoLfcgTFHONJ2W1tWo
dTX7rEnPhm6TRr7f/E4YB9+dRmZ9KXgsAP9GuACQiiHQjTxlMgA6yUEHPaYfl6dm
lGLVZay+E/3m0/zTUmJw4Q32MJsHeh0UFl+4tpUQFak/JNkoNw+/p2ibP9QPnh79
gWTWq6ZOaj5xYILzLA/AFvD35A4fqzgLuh4pekgjUCzm6oTDMqls9pFVyg0x0H3R
Nxg9HxlVMFHVEqyK2AtR1Q==
`protect END_PROTECTED
