`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jda+Ps00KUV1YHSjR3M8mWmpSQSOQSWHNgBiuyPkBRz2b9OTIiOu81ZN94Ch3koj
2e5O6xEBqu7YfqCRrOs9ih3N5PSqvn5B16pMK6eBeedezNlBPtl46J3Bn4g+ISxZ
c530teii1zw+p98s0kThjeAmm+z42UcGUXaORgGz+X/E8QqYQyUGBBpi8rUp70pM
U6b+YSVDt2HRaLRsbCbED5fTO9bv2MJjS4gmRn6fWRGhZ171sz88awF5ym7/WIRD
AkQ1CKLW6PcJOZGWZAdBx2advVYLWhneHCnnWLl00u79qLV3af0faaLWXYUq++Fh
baGTy4k2hdoczX3pfAIXvtkYNy9Be2PaxQCjxKScd2SLjMeHOSRQ+p9Vy88XhtwU
SDuh9yQK8+uB675Ml1/P1+K5o2+qX2O6sm35EyuAEnaed3ebfJHkdWRXMQ/ECPH6
z3glcXx3YljP1T23eSU2UCl5rDDHwyemk/GC/qVyBbW27cbyiz2nJSnaPUybgjtV
FXyNzpeXfnva9VPXtxXU/CWi3GDY5WkjZxkVzSF4sVt8ESUGfyk2wzU2g1pQNRrX
r1IguMdwsIQLyRqq0Su2yKNiCN9bRG3z6yh52aEvyF8Jn2nimNa4u8GnYcjiY9Ws
uuA+y1By8G+ZVGspIMCna82WCRqnVA7PgcJdJFJ73pUk3xcNSJ+Jnrv6TpeH0Mbb
tUyKYqH6M0RbUdfqkOXmEAXJ+q/cFkrTJSnEVIHHoZj8X+H54TThAIzuEeTvrncj
aBaJgHIjxb5Dm84hz2SA83gpbcQlARt/EVPNspNfgam6dT63LBmQl8qo7Wfut00o
0Z4QhE5w/wUu/lV1kvtAeHBggGz8uK4+7uNRj01NBFZIkm5CETfAZuICfBHKE0OK
IK9vJ6wdlMwX0u8XPEYvZg==
`protect END_PROTECTED
