`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZSKn+ETDe1+cARC9M0vQ3JFuXf3N0iRK1VmXfV+/bLOfibDiDgNv9NRLIWofMho
Gh0plJBs3FdWDjIj86kAPjgp+5kQx8mr970Pjmqyx5xCVPzooQgdJVjTSRuERdJA
hO0t6zqe7Z3vmM4Rj+yWjygfaYDiQ1m12PyPwLqCQdI6qe3HGdLvABe8r3mHVHG4
OxoAinG96X0b7fx/AOKznFVUk3k+3re/o5k/B15sNOwtTDkN7fjd8dYFRzF5q3mP
SbQpVLig/lUgxIzub/zh9z6acX9FKKaoNiac/EzZPMTMs/wbz1f2fY03Rcbv5X7F
eQh9wgIDrwUdiRNDCTBtO6/SvlR2wsGs0pycnB7SSh9jJYPehzHZvFn6/LX1BaDt
HPeo/YTh2Hph6v9J6q7vAQHaFgrbLEYJLwY3kTy9NbGRhECvX/ypx9F4maqpMVMS
MctODC0lZg4sxOhkwqjFFoysiE6Fdx7G2X+ne+CxpR56FBbpe3Loy+7qTDeFQBzr
7XHIGzygBw40LVyQqldK4nA5OLJjLnwATTWnjVXEn8wVLT2x0skdFb68k4V8x17O
gkpBIRo1+2dxsXU6tbNCHQ==
`protect END_PROTECTED
