`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p09TbldwYznIAUrUqMsZ2BfQQnfQvOLOcqc2npcY0ugGojORA2gfCgqMJInHtnb0
yOKb2NHZNYbNhuP+2yXsxzWgoUzjV2CpGEde1udG2tI+qhk79LO/PYX62rMmytc+
JcLQEVjveV1FjImT2xIg4PH9bYHAPrh2S9hG7XHtjmUn0DDo/ODbiRUMVmQv8cG2
Ti1/GinB0eWbO6RZcqOekUhB+d3Tt62H8Is+am7HFhEoZ8JpXbLnXDCJJ8Xls43B
xGGB30AyfLjU99RWOqlHW8w08Qh10i89vmSBnmG0f5k6Q5jpX9SjzgWJWAnQUleA
pCWkvtL7azHV3fojEWMstg==
`protect END_PROTECTED
