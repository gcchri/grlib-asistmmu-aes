`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bAO/BMo1a5X2E8f5aKW4kj2zshehmeLNeZHeSJ/a2yTEFmHqY8dry8Vx5pwIXJDO
vUOB3MUqwiWiqdjiFFk06ca/pBmwCo2yTO15y/kNpQPvnLJprqpGgFDB7v7Zcv/X
JzjzbpPvlsJF5WPcQpiK7Zo8MVKROu0u5Bm1vBYT+Ehjc2R0qws5Nnro1yQpI3Qh
4v+tl4hgYqvGVj1G62XcWR2xIUwZvY9A8AjikgbFLplh3FVzCRKjdCnoUy4sGgHw
1jVtjjLsj20MS/iFZtDy8lTFjPSVEbeWGOGHECcT4EX3s3TXVMgr4YubeGsEiW/5
mRf1PyiBf/RCJM/1A4TZBUXjjx7y2/NwiTMQNiUjHF7/kYyFn5VgnmTOfRM1V4ax
/K1hNjYq9AIwwbhPxIQahXGUIisz3U8HoeI6STqaS4HERglr+39kAITzH7ixf7K1
Kr38kJIW74deXwzDt4NkTiMNFvQUiCGgmpHGUK2u5HLgYTsr71crSsBqG42fm6mm
KAmKbOAfU332pOvb6GyClzBnO+Oudbd+EeV22fOT83OcUDPFVsyqgILC64PRJ0pH
uKW35BOXLKg3XnZr8tp+uS0BTKxJPdjGPqFR33r4sqigLeC0lUBGbeMC8jqmuEFU
kI0GgEWpwcHG7VDwGiVp7GeeHNQ6yXcNJUEYSGAmDpW7CtKgPQcyo+GPyQsEpzxr
S1u9JxOe6n2LICH78Nec5sjHfdw+92Gbav+2LOCtSATJ1FgjSdc5uFoi0+AS6bPp
QiV6V+ndIbk4Jvna1kPyVyLqmjjh1W8i2QTV9V8yBE6RWr6zwapyLL4bR9W+0+zZ
LrEaDn2aAB0WBY/phDJDzARVhnkIxc7ZHXNqRtYbWVViemG6J77Za84rfCgeEpql
hSvYu3RgCRaOdTDNMbdyHHzkYwpzUH40HuqzfyUHVx6Gr/eIazqhAPx7wL5RmB9v
8XsizOp1aToQPWkrtevwhJQ6RFgboteF9v/MY7H+3dJUXMBR4Az6x4MHjCioVdCV
h4QDSoN5CyA2EQYmvVMztW5zBMFwRjCXkQNd1kS3Zuct1jsbTZspjqdDAvKMWeKk
Ihb981CzjT+UP3YbR3uMenMN2yGJ2tiQgivcfRjlKtd4kR99ty2XFsxEvtQ8dl98
eCnurIhDQowv7jjfl/8nIBDxzvyngHg+/a0Z3RO1l5Hpvnem6uvx5KPYsCh07V4h
DvvtD6uZSETIW15wr6gvOgnqiLdFfn9HqY6ZkiOEudEPU4H6rSJt2ZKIjS9FTD2T
XKFLJaeU5Oe0ZSef12j77CvkqeB6dif2c6WBn6UPiQJ4Lc74xFaImhTHA06NNMb0
2O2IyhVR8qwJk0QgivPAefgNynCadZjQQZlsecS9h3omnRk9ASG9lbFvZEQFM0PF
9Jno8X+yMNthHArHK8Btpewa2QPlAfCDdLe4oK/gPoZo2hZjCms08Dq14xxprWNN
B8RUzvChmqQopNcaTqqCaurDlA2ddzhFMUrgfzPSFVMmDyLokdALIUnDsb7/nDS+
ciexOI+oWuUzDGZkmZhmsy3XqiCxPjSqp8TkYBHUfbdeI2bJR28khf4HjR0nZqL/
l8emu8mUgwRyE6sdbsThNm6J94E6hsTI5oYU68K7Jh6vUy9NxQt1HWu+oSoaZbtT
qvhfU/DDmnonb2AWUK8kfJ7d8xSxWmHeJTJ1TOCPlK8v2oB5hhhAtCrLuNny0nSa
qsZxu35l7L91XlZbN90zx11IPd5KsaL+cJUjm111eCsvND/8QlGBZ1VnfP+ngzFy
8xTu5q50zPCw89Z/Z9z25ZuLpwhv5ekDX0w1jDND4X6f+sASj5FO4co2J0N2P3FM
Oy2rtuGNU365Mf+SJrjENhthDnypKqS2MIX6+cJbIjZWbI6hCsmcIPcxoeW1K0Iw
cQS4SC7pw+IKPQjOJGPvulWcfSW/BMFEw0fOm60w94+NyN9zjK5sAV4w6VIpQUxu
UvhPAgL4Rw+wRso7D3vgzQ9MdWGLKAcV58g0PttlcolOirQ3YeVaLT2cg2yWi5dd
IUO1Hz+5eczzeqIbg86zzKRvBs/YqwQcB/OGJCs6Z5HM+3Qooi32Ta2Q3je7tthl
xp3eSaydgH7h54hlFbfOH8OLWEioknbPCP7GwH6JZTkwWOXv9gnkLFjYGy5pksCq
mEqhJmEYZ7HAy7+GVNxoXHqj08JCT9hjd8d7BB07WysoC5GmZa+23ol0yhFgubPc
GthP90P6j7HkvLY7b5eXZeoQjpO367//+/9Tuc0QSdwSr02gnYqS1HowGV9RBa0g
z7mQ+0Q7mwAHzMXe7VoA6Cc8enHhfAmrfL/FnjlTHbdY4AG+a/9rmnJlhahqkGNe
qdDl1eXjxgiZrM8D3Tf9huGcptYQuXRHadF76T5FevCk1BmWYsa00DMnkdo43MGY
kHCPbGkzFPa0tUN+y71bL6IUtNhtH+L0SKlSsHn3cR5bMfG2Of1geOW7xodwiv6e
AcWd+Cfm+LFbgsaaV0XrVHNK2hNFrv81cKHjWtshYRDRY52xetYR3Ga4cRuQOwY/
s/Jww7hK+uUgO6QeXxNZcfItgaPKRgdoRERyIaty9w7Q3Ha+UANMDSQyoUtJoBTN
NsOoEv35Oqi8W0uw45O77uz/PEk2VFhRzlB5rZ0mq9u0l9/MT3L3s8SMKo96yU9R
9uWbJw78+OFSoISWHLbEYdoNK7OdtsaUzVKZyL9WpAnryQZmK43r9BC6bSBnKBEG
61xzZvhmB8vUpRia5zVuuQTAtbRXjMeARt4x8SZJ4VPhRfrBYMmsuOpYGt7q1ZUN
M4oaQVeRo81CU93uBSc7V9A0z+ZaguU2jkyaZmpkOWbdx3OuzFRuq8L2eqRB02kR
+QFrBT7fQNBOlmFB5Z1zu7WVmuBeOy1BeXLJ9xEH1ZUh9RQgJt3D5BrzlZHEJesq
i1UntoG2WqZCmICOUcLVhVNKZdFUPvkMYmzUc2ipoHI0A3VhpaJnv0FKmINjcu6G
LwzLn8ZBGzRgIzcQuwvJskX+22r/Dn2022aWGzeyW6egpDvk7rW+L2ScL3dGT9n4
rKah0ng/ccvavZTg6QFL5l8/uY7whzrm47rczcTX1cjBL0dGyxY4GOXdyaQrExIR
jP5/cIO+Mxn+Vyrv4DPC1XyU5e3cxjzAAzNT5hviJXwihc57KVbTbr+XisNptQ4U
K77gE7733GduxPSWLHDZ24uEHk+yQT/Og8Fd+4pIXKe639BbTSucBrYY7XADv0M4
//AxIyDQnsfoXEkYiuInu7JP8X1k1JC6CZF+KokwFDvo1LIRTI+TLtXh1ptcikMv
elFcPUYnSEHJ15JN9FpN9jYxJ2+shwKQ9eeOVlHToHT83w4aFdYbdfHqykW+XwBp
4jrkWWpgxjJtGdb/7tBQJO+ftZeTWh2xFc2Imc8mm+9EZKI/54ofoVwV4aQIqc05
Iihw2haiqO6p/CH7NIN/fEH9H6tVAnFSAE+Z4PzC2diBLKFWNVDi28yXpV2ig+zo
B/nQYYwiT+slRO0eNZWUQN4tTj9uDc1VJp8+bivh3VdN8Q69juo8HzwILfYBS8bc
3Ldq4GY/bb53NQzrL9cMnz3rr09HVVfYWKX610krO/mPi4/1hjazrAq4XC9EKqmq
k31sHRDICy5X5B1apFQ4fV50GPPKM2DbYGc36EU+ohlAGIuNK5xJtQ6gUKEj5TZx
m55ZPUAbgPhtDXc5XUFWWpMTPnVANXSI9Zcn/M04qxwUBw6Wqw1pWSMeK6u3W81B
pfnQBxAxy8fjk1GmSceVyWoSWpDHzFwuAvDDLQ7ALp2UCbPPEmGDKffqsdAtKCwW
c9fFo5oa4RFdZ3PRlkipFVddYz/k5nW0YtD+07wmaKakv4dvs/1kQyKWw+Xdids5
KZrvPssyPQxbTNz78HTmeL/Tg1jF44YwdPwxfI1ZQDZcdxegTbtTm4TShe8Cwwbh
nAbNX8PryEfj7doaq5Aw2VmnAN2DJ7WzVMqAOKaZ4u9sej/hUy4atMb/GLADJDoW
57jXTOZ9Q0RqfoXT3L9W7mekD1QRsNR3XPEdcz4+6BtDjO/yYFcqZfbpEbjaUR4C
dE03t5hE2Kh3QPaCiE1fI0pwKEGZKQjeA04RGEhTufd1zljy+Iumvwjaq/yuhVWL
dt40pF6WbjYLxpeqfEkGFpMFZXKcwqmsDG1zemekvrJjrZ+71J3p0E2z2HaJ7yEs
3gYeyGN1gyq3quRnz90a+tvQZruvVVb1iYa2Z2+rK3fs9/kYTxY6sr2hgGARChvy
L4ZCAWNBxpYEl2CzbCtbKvD9EG/ceQvviDajY2DrDt7SZRN7HMkV/Rs4gg0T7VfJ
0IRdUxVsanxDQZjKqq6MqcuDxUvQSWDW/YIrqJYFHveHqSG5r3TqT7c0fYgVYBaJ
jTyXlP+8Z47zb19wZBUY64QcLPCfJIbLiz7rbKjUwRRQlUuyCSeg0uBrEar0xtEd
tl42oIkH88fSa4YS3co1i3HEtwEs3Il56Q89UIItTqS+D/4HhQDn5cujcSjQ4S4u
y6C4Cik2kHhjTQgKzzdXivJSpsZ1M3xsXxy/+AU8wmv5PW9RAfh3p7+xEys7QP3T
YX7CE7jR5tjvPkoxfoJzn0eiEkX5Y2MroLG9rgiOhw5JuFPDrzQdg2Gm7xphFB4K
tRoS2nucsjQvXrmUgjlv26mTec0JHg0hBrto0YST2IqNllOYIc64D4gDVHHsiaya
kYejO5fS+MFw04gd8BVNC235O5LS074Q/wt5Yu+TZGnDBqAjjA7SNWToAHBJYgfd
2ndE0la2b/r3OVDHExYLsOnXSs+xBilgPjhBQO8khc2EBLsOviCix9pgUXzc8nNJ
LRcwpqGoB19MPbNzfZPC/uu0zbXNmxnTqKtH8fkAUFYG0m0yAQT7aNYnIlrN3SSU
FVakjQ5XbVJ9GeqYU5kVh6gyWOQxnAKe0bMlTZmeSALnfDEgHHAnsUM11hSovVKW
5+lsikgNURu8SN8jySLHuXmDaMuH/mg2FRyWJEnXDKxMN4AYcWBbFfPp9sfZUZ/m
xhp8JlvH/Q197PZHA0D+L7tWCLR5xa5QMUHNR/W7WUcXza5UpRTMAvWv4AgVWlIa
bCq5PdJ7cnJbHU2KvxzXAA+trP5Cd7lnj+XSJgAbpANxfAi3HTYozbQ1931CW2bP
0pZzal+iX37D6jAh4d90UJ2RHeSBbbUHmQmC1+YjLZ8HF3hxkEVbBYWoqFKQvwQj
lxVv+Ru4Cl6VcjemqrpWAD0aG5UaJCX6ljsxteuiH/F3d68X8Jjhq+g4SXX8A2wZ
VIymg7krYbncXeP52sfewRm255MRV4mOuRtMKfDeFNcSvi9Bow4guifTZuR8ngs5
s3T6ebPKGkUFNL9d16ulB1EAZYFMsOHLhE/tlxbWMbrLYCd3VAabgiR5Ob+YUumh
qSIzFcrg+HUEB+1CcbsNxNyN2N94HHsrLd3GF6VqRL1upoFXzU0a8TQcdVQI5C6p
Cf/7gKc64Yz5DkZOwwe57pRBQa37yD6nAmlo2OnYh6iuV7eIp9FLp+yCooYO4YNf
z4q4Kt1zbrupb1/Oj2r+uLrGrMQSzFZjFH4lCMR18nQpI5qsSQf9rF8bAoBNyAbq
q/+D+7EjypZizP2AtQ5hNnJlzrfai/VKz7n5ap8GnhVcFs58miqGfic5Y+2CHiBx
661tdXV+PdJ8bI2KZEDyqwU805s5FJ6kYMvQUpFIR1cu7VcfVMNEYyeFYvotDBCo
YWjFt5ya3XVtLFE0Efbew/cZKhF7ep1LOvRg6Q7jwciLutrhPmD3mkgFIgiT70y8
6DWj/7VOuejjscneXcAaqRnEdds2sNgAGgTYTE1W+RBNzOOxaN4EqcDygt6unkW7
EgmnRYnnRjSB6OlsJd8K5Wg5n6mCy2SfO8Yo2nxoga0Sas4OYPGy+DMHgqB6Wxen
21izWyQm/6lsq6w859HOjbIBBYLtwl68CteFIuZn0MWFd274SdGvYAtHTgMW8yUJ
P+BrvVsdu0kNr/om2lWLLNZ819ETLIQrEDJoQomzL2OYQzxLJleVMy5oZHpE7oD2
Ehixv9EvPHO5OlYGj25NwnCwA0g8tUC7pI5FlnjbFbCR2MOP8jt/pp6mCEAoHFGn
AEqJFRd95eMGNPPp7GFkjBi5Rlf9nR+fRdmuex0CIFpKu7binBTQxhJ93UpBUlmN
ObbakJkCCf5WKV1nw3CkzdrMJ2H9c08cT6/0HiIiSuKXsgf/iPZYRgLBZATsRJpT
Krk4K9bvSw4yhRUnruJ6Kg8ONficoI+GcAh32LX7q6pjAjYwLlgC5OEHLHV0naCT
4PmKbZ2zgcsqukbenXabZ2/XDE7XX9X4G7StdzXwdhC5jHFdj3uD3x5hD05SUMYz
IiGK8TTy/B+y/m4W7gC37r2QbWCIA6udiZh5/twjoeU=
`protect END_PROTECTED
