`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7/4bvySw9X3PZcGQLWUIcBtOcnK3Rrn95fRmA57rFfqRyyzs7eoHAXO/96cocK0
WlzZ5qJ73tJO8N/gQkDrUUCXfD3JTx03oUUP8E9w+jVq+zm88v9roIWVWZIZ+krW
nZH4+SL3yjWN2WwIrb/snIEDLA3lf+kyE4uH6+0GAVYjxiMlUaRTJh5ebPNLKlpV
gODe76zkpuLpmX7kcIhw3pojpRgYCAJZlqQ1KY9D1RL8GC7y7B+73PvxFVofqppJ
NRqY0CdIiPoIiQt6goaINSJ4i88Gl/1cMwg0P2HBg4K90ZILpaS6jwpabU94mcZg
zF4db0Qok6VsW3JE52+4kkfTf0nCpWK3zZiLtJncLUfjefWXEpD1aClOanvRsh6m
7fBb5VSdM9K3eMSi7zyhWrTXDNgBQHpRykIyeqnK1W9thliO/oJwHKuHx6EHAMu+
vcgi4LgGWydIcfx6QLwN+tkdsjjY4GNTch3A97Ef34iRfvvfWfDeS9I4cCdYg97v
+UtXackMmTmLxhEnOAAqdd/CygpBk9DZ9d3j2VRY4byMIcIU3gJhtIuZFg9TKm6H
`protect END_PROTECTED
