`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vKvDga+HCo3P/D23Px3+/xbpCpg6PTzShWFlIu/Xw9Sd4ILs08eTFuklyuUccBzX
H0/DlSm6VKhI/6qD94c7QRLZvpRanOkSiJT6+6kVUOo4owI+lKkafElhj0/aOxDs
3F7lCbaBS7qmj13FFFuAlsbzob8EvEz2E2azXBgS2KjPBylFWjWgq7ItH7zlldTj
XiTjs84RciRo/wiDK6cHRPPEdwZYsq45FK8Jw+Ml0zG9NdLxGUqTeSk5kKCLTicx
zz5W+b2ARMRc/McxYm9A9v+b9dqgzHQRRDHbRYpuiqYhI3Ew7FUrAoAfMz1JMt5o
Jzg4gi/ZWeMMu6YTY0A3BQ5ZVVMmB4NcD9kZd+7QBufuu9mtcCSASGDwav1xLaxu
7uAogaap8Fc1Pe17BLBn8odv5IaPxcSc27hBohs/sU/Y/BuJlwCu1B9vR63ivrsZ
5+XBbktWBRiCI0D6YhcK08458KG5C/Bx9+TI9jjyuzS6FFtl7dP1Co9zk1lDX3It
7bnuy028WCAFuRKjhP4xaDO5G55v3WRDWiz6V/lHNrDaZWlepVyb+DFdOPNqwWFQ
O741++JKO6ieTBMbl7xIHJhSHSETU+lJfqj5OJkrANg=
`protect END_PROTECTED
