`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgmRisvp0hD06DotIRFl/5FOxz+mFS8QkgI45B4F3MWe3Hj2eMwpRx19w6C6zlCz
btc2SA37UB+9LtX1gyMPzsV+7X/Ks3g86uzGK2WPd8zuv9/Xqf4sephjGR+Iu6rZ
OqwkPxeH7VYrEW/LT+uPf94gP/3LsBjxdonWf4nzSWwc8nnmX2M/1hcggKdT/p8S
4sqAOKwcfnYOc5u7KDpwjsAmwmG15KQQcNgv2/LL4+PHV94brlqAo3qykpWAgapU
HcEYEQ2aP7zuLiwioy2dpQ==
`protect END_PROTECTED
