`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gKno3dt9qwX6m5fxvNVYF5HstHbW0DlozSPDScrEib4H4ZbAEyOB09hXUyQ+lNoi
eQSg2Mg9zttQj/V69J3ldaytfURNBojodJNv0z5F7YuSqjs9FTsEvhnc8b7qst1Z
G8eSVblRfyMdpjOT7lnP7ZiDiaQJRHORt88BjWxPCEPlfmOS26Ks0+3yvnmCdE+c
bQ49aptlc+Ld+qLmfm/JSxp2Dal7EZrJl769K8gWPuihGAgTyZjANfNadrQ0DrA+
5kDDb12+Y1fYKm05FhVkGV+cIhNz0a2oyxaroMVSOTMdVG2PT2RmLRP1x04YTbn7
`protect END_PROTECTED
