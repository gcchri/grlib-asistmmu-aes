`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2VYHgDeiNAD9zTS6Ptrgk9ylbRjc4DeBKH0M3kShy1havM2cTZ0hlXmk4CnMt3l
qZDH8F/Ol6fp/d2pBTrgsCP2vWn9EW8nNboh+hobBSj0B4TnQC1+tADaYnFsV6qm
p8/pC28A8NZqHBAHHgpawy5/ARVEwX7reEm0Q72A8EkIAtP0qdg02oztnsyWQs9P
km6GgPT8BQ/nr9KeDutWat7EJgCC5mJZ9IpNCa1eRqFWsIMsKpWoxIGNgH2rx9mT
axW2/1BUUruz9saWzKfpx4TzizWDOaYGrQwDZPZ2FRoB1UyY8OspvEZ6QXL1qscY
oANEDMFLM8kxwVwmTk3D8wpBhzKr1c0AVZVDHqVZ4H4VS7KsFGcxZrHvlRAu961z
iXii/XZz2jWgTP6ma48+sKnQ3eph8NbVIjs9jtYSO0OhvGQbkHFHfhC5hjxn0e3Q
tU0UEOLYMQzqeOECKgJaomUGBL0KVotbDO1PTggYsxCGp0ia8jEpob0O3dh8ogPV
GL+Odw+PlbTMvCOti03y2vE1ijVdkz1aZrVpjL6Voa0gyg3mGqYh8Cx6ZMbwDmL6
sggR0jNMauGGCv5N8Hv/xjnzyzFL6/bMjrwh9dnNfk6JeeOKdJFMFNHQNr1o4NX1
c6mFQt1uw7AkBOSgqTUEPcxrMSQEAoQIkYdj0GbxGDe9DreEaYf+lLSZxHTRjOFX
19RO/ID1OTz968RkC1gB4msFPfJgnDfgktqAgflLBCa0jCV2Xqw17DIzG0Est8tV
tH1MoR9Pk+D3x4mvoBbqnupneaakuJa8nYbboH1U3eZZ9gjOg4sS0gXBGMeSN9iE
I8j++woXjrqHfcWqAo6ZnJVBSsYTxz534tpAQpXAnfhR95JEnBD/TUrkJe6MXLc1
3RIlU22Ct0P9XkBfhIIbq6LBvBozGG17nQ+sB1Bnaz0pFiu3ViYqGGJoyZdeaaMa
s/oQOj+r+SUYDOlDdYvII2A/Z5z9sckeF/I2OmyUUkLMf8LdzaQ9skshVdFPsZqz
eUbk0Ha1zWvm2z132O+7fKoxVIgIzXOvDLI2OgcLxdDundFTr7aHY55ehGtN/ZX/
Q6lQwNT1xbqhtZSW+Amw+Zo9rL8WF14oFRpLDlKALXSw++IPDk5UTyc6Vl4xqftl
0stwGE4BlvIM1/771+cZows8QHzlZH8wNXeMVgSTSctXlXTbSZwyGhOIqUeOsHle
2Hg1YpOj9OwYVi2Fwmtu4IA3Nx5mzRHkTpGLevoqLEOxkMzhfyFYm+mY5m+bi1Ui
rqz4UhgvRXy778ICAMGpeA==
`protect END_PROTECTED
