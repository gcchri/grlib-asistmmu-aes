`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWb90CjC33fc5K6xNivDaf90LIoJpThCwYN1CYBIsBnP/iqmn/6GdKqq+52OrzHb
yXvNWU68y+5A2MzCnZIlW+fhlwtCVOKKMIP5yYYNfM9gyGePGwXVt9x0qewEcGlc
SNvkaPgsp5IsV31yxg4Ojy2ft2FbA5zpc3sCxZBGE83jgcH9G0PD+2KtCK/HIioV
gNAOtzJbjXNShlCDZQTCmE5FxY7lJsEIK5QF5AeDgFh3oFfhEVAa/7NuAFf3p3os
yXxl3gTN5AD4grSMANWJSzoqSmVho59nkoWf3zwXUzE=
`protect END_PROTECTED
