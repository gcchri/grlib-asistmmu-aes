`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTig2dd4Vzl4fsbObUrzNjmXg/z+qzG/CSvy97lP1PVem+YPMyIEn90pd1rf+bqm
wj2QO8SMikNRypxH+zzTgUHWI+ztciut4zvYha3unCmngSAwYrEb2ioo+rC0KiUL
TUM1B2rqtq6H8snhudxXUvfM5Z817U3RqBosZgnuJrRbr4BB+cYSvHXQgCQUC8Wc
Gm4Tf79BtiJVcvLja3i0Mbn2HsZDhoWkdW3ITAbQ6c9zvcluhArBkn5mHYD2Y+pc
smkO6kUQmVPgpi0KvTqdhsiv+aVU8RvHbFj8wspsseRBrhwTOiA1l7y+ju5Zm7oK
hf5KdE+8YGSkKW7z8g5CpUDxz93VGCoHs6KXmwCr0W+vXn3g/0wQkMuznSGn68Rj
`protect END_PROTECTED
