`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jtY6ryrGpP3fzn/dMTjWmf+0Mgq/L5+SKQXqjYVeCyi0jieFZd88qigPO0aK+MOS
5yFFfEfXlgxQEdFWL1PlrlXSMN28/ifl/p24uqPMYY8Eri+cANIvBsS0IDZ9acG9
Amm9TzMd3+thOjy0HkYihLFmZiJEcLkchmlCxiTliLxampteXZshk5hIQnKFSRzq
ZcflamvUEtjp3224V8/QOUG8fYLgQ4ApIdDzJAkf4AvQPu748Blvwitk11RK1qAU
fkzwTtfF7C5fJXWP7dIPzubALANTllQpGUCL2cXqo2akyM+ptS+BbDQOAqDfUjIm
QC9S0VTKkjZCJiq8tsezlBAllrcSV08IKNZePaTFdeOlqjxU3+jxATvGCZ8Eqs7R
zVxOWgXCovVzGL1/uutcAhNbRUyU2V5c9jCfqTVTv5DEaLehH+J7rCRq/6RaCBpP
uUTCLV2pMFLw/+nXXEtZOZI85g40gLNrFiaeJFPx6RSizCLCvHHDDZR9V47Qoq06
4d9qSd3IB8Jkgxw13axYBa17WKRD3eeCil0bX79rPb/3bZaHVGd1H5B4lEgM6wvM
O4l8dxkjPjpdSaBdXTnFTHLuSP0unYjmdT3Qe6CinmkUk0cFn4NulVj0F2ipBG6f
NJ+zKJQwDAJC3YQ/0ZhSfuABiSOT9FrNgBVZA0JCCm+iUm4X9aObaR1ktzh6l+3G
zpzL9YvSh7/uacCbNsSaTmTQYOfZz8O7z19jGc/YMZ1bCFkHCRHUwcnUS53iB3i+
rbvk9fVxEnHUrrGgqVmhSWl/jYqUC5z8T2ZoStcKlyZ8YLJfsZfTW3H7qmyNk9zr
yvkfIJLg8284wQgfV77gVB1KzJynyYbaNv0/IKGgDvk8+W3YMblsYX80vJEGemmY
0oPG2soljjZCKrO7e6IxW8CzaH+jW3z0rPoIMjmrHgvxU8V94AUA4YvH9CuwBO1p
pUV0FhGt39kXX811G2e0izrnUHsoeZ9RhQebA2mCY3FlnYEupNxIbnHv984AEsgl
Te3Mq029xsBukwnXfK9jGP8PApARWFBsAu2mNhLuN9dDlxf0F1NSvyLLaVqyrdoQ
tDDxyu4p6HaW09PXz2oZdl8qiogcA203Vt8Hxuk166fAjEggXh6KiSD8KU/fpg0r
mHEXfwoU+RLG6MUc+IP37rWtaf1Nol1D5XVYILLSsNc8U4HdaA+f8e3//1/3jnxE
KkWriIJB0uK4xLTPnUVKSk3hl9GUdU46QjvGyjM7Gvnxi3VH11mRzJcmu96igBW4
8sDFMTifY+kcUcrP5/8YEIRm7i+3ySz9OHwguCvx9KziW0R8aqkxIn07OMUFU+GJ
PxVV6sBQW7GrUdt/GM4hIjFXvIDjzMVWH+7cBvTeNRSHoiCYDPv4lKMBewMoeRTJ
mdzbXgBERaiQ/2t5V3e6l4yiDjV/0JPJ1QQWCuDhNkrO5dlSv5TRdVEtF4zuo3ag
XhE40sN+SKUctg5USoXs2AVFoF8yiFrJMwMrX92CNg0hF+9BJACSTwOZpdzRKgkA
qNiaTJ/E85aXmFZ8R1td4W7ZRNuo/oXAC8kIdZbCw5FR9x6atdTXfar3sK3OZHJU
TYDMjZo4m//IkFqkSic1z9rabGo8xD6sCjddVjUTCC8OtKW7y75QABYPCWu7KvzD
87fmZ7oqEt8lMfKHYtdkAEHZ0RrE9JMkruVkwGfiJHcRDjGhEIDvDH3ec5YO6o3E
BNggZ3gaoqWm21hIAEhkiByod9FtMe1K2trRBLZDr5Vy1c6bS1W4OGDq2DO49M4a
55jo14DPQHmr+FB2W9HZSCSsyGdg1w5423loD9xIjxAt7qLBXfoUg6oPyhSp0n2m
RR6Kwfepow7FgsZ8ZvVqBMRVmOPgafFgKPya7LZbYui6jRQYbRhRY5OmOxEl+k5d
7OCnq0Ovrv6SpyFmvMdHv7uG0BSLLNxEYqS2TZi1NAXnhF8OQb/l8N8HjJqNQ6u7
lLbPn8UroA4gowHsPq+ss1Wwe7Vze2hGlvWOMhKwWK9wEsPxUQ39xzedq9cD7mne
FcALmIDkD2v9K61ZTHQHea/6b2XlU5OycFO/bsjaFbVtXq/aXmW9LaYxFM/tyZD9
qMRZAgC/EGfvphtKqxWfqVCBEYf8kt0sbsqcagQwVXf4+JGr3h2xKvHjFn9oBw+B
z4uDmj6jyF80jeqKaH44UCSeYZ3BiTaVvWE6oKFB+taE4R01hh0CjETO7LjR+ijg
MOkdx+8WpJYMIESBFkGB0/TcM/HtZ+jzluCIuG2w7j41CkOGbot53BWJbVPr+Vmb
efYLawXZMYwpkURg+dH2EXi2wqhumjnV81MLOG+XdMbaxpdzQ2WJ0wJVnjeITE0c
ZyrR1chTN55P917YF05vXRgqZOFMVkdI8aNmZ99pGxSFg0ULgiPdw/WlLGtfIPTa
6RYWdLCIjYwj7OlzTaWoLdNHWziX51yhAALFwKhQXcz7ydSjEOGaM4+BUzcjrkn1
vrJMf6nYJpZtLmGmpO15tppMcYr8/l5mAIxfxK7MGhvQL+Kh0ey4YQYu8gAHyXsA
7OLhza0x0OQQRMwcEMkTJ8RYLgiwvg6ymrhmjr9BEsDYQ6+uIqOM1f1aUKabYmtl
sjPtdYTTZx4HexpzzmqggA==
`protect END_PROTECTED
