`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9DLdPtO5Hsi49YzX7FOSm0DIv/7o+ct24Dx7zI6Sj+Wce4NSQ/BpqEpOV93TVpaZ
Hty5j6119auqXGWVxitlJQXWAgVXYt+kJTVcj81S41fbTynYyRMbE27uzSgK6odr
zQd/5BE5vOSM1QamYcNfNhuLgMTFdUfPfkHo1MoplKG3YPCRn+UZAY9wPo/rbMeX
nV9wPlKcM/QY4bgaRykkP+Kgb1soAsto/HuK3l1pY7uT2yBsLegpgVxeRS78E3jA
g5x61F3sfp3FRYbNrDW85s6pv4HERIUcqp/IxShwHxN9+HHwNhbqMkC9+ONntWju
kuMpVFfJVH0MvT2Wl0ddc0CGkR9cYYXgRiXX+akkRpVQta3Va2IKDcHDBPgyO+Ix
zu+djkXw2vzYV+A6y1KcEjhZ5K9eEpfV0hiszWOBBJ4=
`protect END_PROTECTED
