`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EFORVBHNqepn2qxToB/dCFjgLjwvoWtpAFnIIu3a3SJhBr5j1LqozDLgvheIP5Z4
Xg8yHg33bhNdW7ZgjJd3nYcEItKfGxsrayqApyd0Bf+PkmnLHGs8ZMnEy56hA/98
wCAfnwbVHlg8U30nFzxMLYzRg0kSOzPhNZKLNLq+YFavk9SfLhgxSPne0b/UZ4sa
AJXQeuDY3khWWxNnoRKUcqhFTNisfOU/eVArWyth+5JaDxnyIHLmwzhAZP7Ju3WM
0iXgD7oD+DCme0VYkU2wlFngQhUBwS/u/cVmstp1pzC86i3aUbT4wbZ26J6yrvnD
1Hm2E8bq+sFEeoshT52CIa3I4UBueZGuJRNp89l2bJ35pL9CBA7pjpxD2kVZTyhW
rSG0P90mqtLKjTpBxIBTIoSPnCkMUQjwoucie+5NHGF9zmxgQk8VWcxPj/TGijW5
grXRQP8+9ORqQRrof1d0ZzelB2UNkYZiHnabp1FPrJASnpVloBmFutYc3WkBfyRy
nPsANpDqmbF3z1U39ENLhvgTmQKABxCburXFY3i0BSk=
`protect END_PROTECTED
