`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rrrk6crsy9g3B6ls2ZV/h2aJoiVekLVbpLtoeTmViXIStv2pR+8gmdDyZGC1P417
ynajLpKlLKa8h3WRtTVNrY+8+DvCCKotohh1Pa6m1JI5ATqSg5JUvrf0nCeF8Xe2
ud6GFeQF8k/zpwEcYCbal1El2rPUB5C3VXksIxQWBLURbXxULzUfho/jlU4onkMg
DHREK5g36+c59WCBO66tWvDuUJhVifglIoDVWC05ldIiOHhGASeRM2wCO/kbMvJg
CVybazQGxD/SQoK5Ze/mFaw7SFf1M/q6yCARkCuuSHhTEexO8tB5VvYZUWVivYfw
qHlBunlJ95ocnMlFEtexV/YkYt+FHPqIWZFYPg4OME5lZIE42ZdY0fIUp0+D+Oi/
YMwvY29frmpttK4D/YFsjjPdHYa6xIhTjYcF+wws6THtF2pvy1LCqJRfTmUhJz1I
eF9IPURnZRUEygaMsd6vkPKFv5rbqA5sloZFI6r9jU1Zn7GM6TN07nfnXjiDTZvC
MQVsSLW0EFiftnfYEo+SYgaXJ5fgLXZB632VVdDSqntodKtPm7NMPDSXRhyULBcE
ChtbPPVhHijeptH9O0O9Lkx0XDdaSWEQSo4Nn+NU4tA=
`protect END_PROTECTED
