`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDyteiQUjdePIjCfRIovv+UnnV2hTNFAd2Aa7KcAZxXdIEjcSX6YVjQVqTF+NjJk
7wa8NlKc8AR83NRL/QwQyHUE6AY+VKIYS4knLgH8YWXHzIa4+1ywY5UMMUyBt+KG
TVbqc7KRjqWYn3l6WzRG9PxN0iM2GDtmz3p6vT+0y5fjOHxXeVWncStG7si9KNGi
Ccxx71yTbBU3kDW1cYTlN1JGZspFT8kifhCj0AV/7UzLOxUdrwhPsNhSG01nyrYA
pYDRa6dFcwTXALfb30mnfEaUBLmAzcbB0WXas56uP8ZO3r6+7mVDB4kRh4c6FGle
pZLLdOYF2XSOkwdXX368kmeweTOFEUA0iCcxAF21VAUo37AugKeTWy0o1fnUT6zC
9v09X1ZzQBsCQrmeBSXx4+OY1hhNTXm/bre6Hqxs8SlJCu2vSvcZaoIFB2+k4qmA
CR7jqHCgv1AtuThRMB9levu+6DN3EAt1qWIAzrJg57/rgN3lOAGVXzbJkq3ABPXf
GJj/eUelDLbI2Ij5oqxn6GPm0oXdyOZbPBTmuqRHbSPtPehNqOyQwqbG7v4Z/j5W
U9X3OP5uRaKOiFxWo52MxuoLqH/SWxvFA65OqvpfMha/JANKRMOuR7Kyje8/lv6o
lLRoCE2UstWOSgSFgAMrLnj4v9KDDLTloQQOA1s6q4MuahHsdQo5jRDEoLPnFOmq
vw2JQIED3x5t12eZlQZ476KfXgN4gTvstr5zOniW9j+Pn9IE0yJuAOVLpZOIOEOX
/nhTtTd4FFOvdTWOk3PHNOY/jrtahjxNVIdhAyAQH2n2J+MO8r3OVXLQ1iNHCiZQ
4X+WyangDtjXoLoZuk0TBx3eIUIsB5vD3mHe3xYAA7c/KYEY/LyHLOcX9RfgUa2g
RdlZ+lyYaI0xWgtiKaNfGNymI9HwPuywtgzthYwod2yFmeCJezZpVWxDo6tJAv+Y
Ldw9KlAmhcIpFdhlkgxcyHFtqKygz6cSkcZtfwyRTcnHxYG6zz/vKHK3r+o7c8bV
AVsCkaTX5U96QM2fbmJNiR0Gtv2Hqc3pI7vBilDLgaofcsNluhftWD8BQBrSIi3+
4klM4eMzF8uwAgXDoSRk8pPo15rVgmYAoPs95opNVuTEr+SjfKz6dOfXf+DX1T77
sUNCXLWdzDmD3uENW7zgqbKx2hA0dHpyt26GKWXPLenye/QzPrVOmVBNN9DXbkPd
+dXnBqfL3F6v8H4s9dYb/QQ6rcMnbVEvdGSQKN1YMA35vzA7yEBZQ48QSMGPf/li
F7JGMDT7XZxUyEPEtotLLvUWPK5BrNu5c+VEC8hHc1+l42XXG4MUA8uBuNu1phUx
lkPC5tClzmhu51Sx3R6k+LPa/jrR8C4E1LwyjI1Jyq/GvDN2S3hckhbAK0r+To0a
eiozSKZN5wvzzBe+g1I4iki6hwmcERs7ZosG6wjeCWqrPRPIMsYPCtGYLDo49Yaf
6FdlAc22vOAZJtRehLXlcdgPQiarN4A01GQNqtlhOYW44etc5immmkSFNzlmUQnZ
qnFeb3LfhdNMb3yYLJY3XOca2WR7LrLSHD8OP3e8EuEE13th8IKFB5xe1k0VxxqJ
mi5eYw7BLxOq5VzYTYhhJbnvkkcZ31ldDvQWbTsTZOv7OvpQmzqZrx4FnhdMZxZj
0krUy0uA+ES40vcyYSqR10/N9+4f2T6Xur6RyQK389a/YzKryecAGLz5J0Vn9a3K
64ZWJJp+/h9B5U/qUDltcC0pzyCvnt8EU9pedBdMbINwIxW4gMDP5L1zP+dR+3li
av12zyYLSZbpPI1W2KKGo80doyyL0jHO36jmR0W3PsMeD3ivspRXSTH9V6uTgxBD
26zo8QfNwqNYJrM6788Gtl07ybahIC1XUB0zYajwYS7v0Par8aeTC8mUbDRVsOEJ
uW3SOMgymUDP9nf6S75dmcsS4E3z1BF0OCDNxV1RWerfRjSjByzZ3XKFYIMd+qH7
ArhIrzpDM22RDsPB9LMjplPxBCRkbvo1Ba9QIKR5uEut3LfJKuppMH43Xr90zrcP
u8cirnUe9QdtxofYGnrhwMwyFhGrVY727ha9doCvEIabYfzGwuMIbG3omjGu3OIk
RhNvgEbsa9W6psNT+LjXvHxeVbwiwS6MYXkLzEjm8mn5y5HFORXKDv5M1FkTQTb2
uqcUjgPZKAqX1n0zmj3sq7ScSdu2y7GGfR11PSRwDh5XXRN90pagv5/h5OmCCF1Z
ULog1JFricen0nhYBywey5WtUgYrUeGHJARG8/mUtTuLxmMcTNLt5/6rqhuzkriz
c5LuPzBwULmsYsYhctUfXidzn9UYgqSR5+cr498JSKzRZAXt3Y78B3/Brx++T4/V
xEp6ce8+3dm8PRTSK/b9rvyHf+lHppM0TFSA6f8nYrwIrXTiQGWHELBGXrlCiiek
wlcRAwPSKH2QMces0sYOCN2dXexF8J4oM9j4i9+Kpo0E3vAdUdpQR2Zcfw3Cslfl
hoEKwIiKFHcRnwi/yDbTUc14/cEpN5MR/JqWEdTILFxOLYXHLgDuZ7T9pCoxp1Gs
bjmjs8TzqJ7xc/zNiQVLveVv6MtDUH5YaAH7+WbQhfJC79ZXtp3IWoGqLVVcf6rU
MxEqD4cuhUt+mJB0fDMZ94Qra2b/FCec+hQXJiPx1DR/pUK1Fu1UbWufu8kmZHD1
xoJzQryBDwfcpWJuBbRtk7lH34srzTghbji9VNYDsW7Rbd3dikSO5j42OORiCvbf
0svN+Ll4e3CRfBbvMCTSfaQdGLRIphQOGyiie0Oi9LuH480ExyBKyo3fubJtcG28
AcMUszjyMv8TztoEcyyuzWsTAobbrnSjSx0Lf18bKzo+BuxueODP5Ot06SreCyeO
FRHL7fAOVMcK1ZAG3WX48T08aL/B2LHgWSQSlqkriqbr84ao5vWy392XYEbPiqRc
dVZeJpZuDbHF8icFfi3v09GUtLYXAR4JoYdCNw0LGAA4f/YPhuMvplVEGBAY8Bso
7dzbuHo46/0dDeSryQKoQyIq76RkyQgcDHLKnWDmcqK7iFQby9UjYJYpGCLPpibt
q2T0QKSvpHbtByEhRw84SSnGghBvYQzktaCDnCn6uKpLMLeHTpONoTR9NT/fEbzx
HMskI7AirArd6NQiDf9rLDEHpfpnGE3Lo9MEe59mP+Bu8wqYp59lrDprzLv3svGd
wqhrf7Yn5KkAWQF2z4CUqtiAV/DIoS9nrlU7PUa673Ht2RsJUPJbmt3ul8c6KgG7
ieJFnyvE6bq7byF3ujQKJ+YffuQ0lm6vIZiSmVLLiahCStdqPIoz6939jkUuzTx5
4ViPLvhzCcQ5wkvVJReW6T0E9g4kIqmq8O2wbIT/zv0jfUjklwc0a480M7RCqSU3
LZu9WUdpV/Y18HweCdl/r6kzMbYhQL1i/v/wUppFB/UqdUwVhQY3cjWDeLTlAS3U
AoOdW0wHZ5hsm1gr0QZSnRhgI6B2zXcMrM8oOytfbQGbsvDNmws1yykLjSMjXQmS
DOo0nyPNVdo5OjlRk8Q9/L0ySSgpYq2oBt2CRNDT0p2kvlNawHrwK3D4sdEChsCt
i+F5MWpUhQW7KDHNErl81di9aOH6nmKVAKGVMLLi6Dw2aRcWS9p47/wWtj5PD/bD
Pc3aJ9Xhqg117y8c2R0ZgpZRhAwYufl6Vh8tfGqoctU3yPALRK/+SxbWXIgYtujJ
f+Blo6McljRb9povbe3AI9mEq/FB25zhN+Co7Sz9ekZpANZmkRVNbp53Cktgrcsn
aKGHieVW1ZME3rMdnPkfrmgzsE2Vq41xjHMaw5SwvDSG53vsF280WVJCshAF6prN
UZ/L4Ji+nUN/pTvIpUALK+sn/rVjcSHeQkiLVdPOtsCK3CHuXl297UG3V5biqcSZ
5rvSJU/eRKw4/bXDUMyFaK+T3TxeApW2GoTPzHobIIeodYmxMs0OkOulXr4UjT6b
/u9ZPHPJu0d0waNULhWxMcMWQt9+i8Zdw0QFWsHdUjLlEzRZqx7bOkEMKoJPyk5O
IpaE/6VJvuszt2IsW8aYizRCRRHwlVknrejDGbjZWLAS76QSeEYso8O38GE3uCaz
8sBH3Ia9Hd/1Hg+EOaF0cok5wIE7D0E2FVTd1m+PaKyvxiSQA+3phoGnKlKT3hvG
H8g17LPiqLzHLYajK1sNCkXbrmB8Xk2XQTCBV200oljlSOrO99+wRb1utZ02BAY+
XN2tartXoiEgAfNWsoTTPGOuWe+Dn2AJ5MD9L+OKSTiXDNdtXe5nzjbGmVcmSq4A
mX9kfUS7MEuYuCj3CXQITzBe8qtxSvNUwHY0QviXmZaODDcW+pAJqyAywnkg7SmT
7BQZL14R3Z1DBR897BL1J6rQJt6AZz0RFJnjXGDG4UJ7pVodfEKL2mgWkkfOpXQ0
EG/3kGEgykJSHP/ZJGNkjQ3V1PJsOBhM3PzpQ69Zf10MGTQO8CiPsmyM3ThC9htl
uUirJkvKsb30stLiiLy12Uq6OtxOachweFBWutqc6bBxhN8HKdLcl7V2TD094vxI
Sgzz8ieqD3Hp24TD3cihhL/XPZxSfOkQTrATmO/i5VWgvLc0TWytBciZ1zKHZ9LZ
pfW/6UKY4spWrqczXnvaQQc9NxEj429NhptPJOmY0lyDMg+jEUcWL7HwI8iLV9Ya
8e87nxd0sVN618XubkS6NV3glL7GmUUzcqbh+zJt9mgglQapL6TOJHsVargy5+e8
8wRcHswqz8gnV5Fedgu0ZgN5HLZjgwWJe8yPvZ3Ew4NXagbknQb2CK7+o8EvfQNr
umJvLT1Mha9MsD4Gx4/dUsaTDkRFetoCDCX7YyCDTlNro4Vn52qqP8xV8CK5rp4B
Yc/H7YLBOUMxiqr4LZEQKH5ZWhKqtIOa9Sx5JF6ejegI5W/bY7Ni4CbXbX7DhHAS
ErWPP0Gd9so6OTanSgTVu+ZxXAowxeaO0RRMzRmrwJLCKknEzUoM3D8H0ti2xJ3l
tCBmN8v75mlnwUL1nOyHyLqpnxMkx4wF/1weaaAK8sKS8+cTQ+dDTSVXRp4fcI06
R1cCyB9dtsKURuXG4gAoOWDmdUu+Ehq2REnrw/mUiU+6bVcq4G6a8lOkahMvthe4
Q4Oo6Rlysb090Rw7y9AVJK/WasAdaH6T6W2wnvIjtsEDr62qN8Y6RI9JPt6/NEHa
IOWZR4wJUcccP+fyikhvHhDR+Ph/StU3sN8Ys+qrCa0Mufn3zK6adhKywZS+Tm3M
1RB06CeDksnfDm8PVC5FqCVWUwuqPqWHaZBmzA0XlP/GY+ftNif6DR1fXvXo3iUu
CY9hOSn7QW7hsS3wMl4vmI6/IbeFkAE5Pvh9JLnclFKpZg9QpwexPWn6RaIwmp7O
XmUa+ndqEer1/zwrRREIDz3qLU0BWPAHrIMzZdahjdeLqmT1euxuH7cdp+6ios9K
PKc567Yh5JdGUt0DERG83Sg9DWwSgw1bNeBt+8sQt/b+tCuYq8sLwlq1betTLAgi
4hfbEit6l9gyrylWkXMHvCtGmjNDUidJ2OqtDlfjGKr/xGCZppSykSkLH4Y1Zg01
xu0XZubFEV0sQ/XAFyDrG+rGLFMJou+ZSs5IIIaPByE=
`protect END_PROTECTED
