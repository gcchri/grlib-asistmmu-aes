`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
22vps+DBIETWMW9ccfB5LctkiaIWKN9ECbEoO5vQQyzlOJLApo2Pm04RMlZrK9Ap
ckWVwYMjmIAqhcRAKRMQ0MvKxqakjL95i26zsaRijW1UhACjYrJ/i5A1DhG3QEfq
JfsM4KpXXdG+hn6yYTHYlZxZFU935g9YDp1pz93km++qMpDGbe7lvehyYf8rQcYG
fXTA0fgpyH7Cv8s1SAV6J+F2mmTmXx24ecS8JSFFZBPAL1sEnvZ+pXFcC2VBRcqi
aF+vKfDMpYZGMQD8Ohau0KRzwD++C04ONOEgVyUENPsu54KUwuh/A4eJiPOquFO7
RPOWbaGOVglXfa7RwEI8bJ2wz1FFWXVmExrb8Bo5WkY=
`protect END_PROTECTED
