`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9x0znPBkdjhGweASsadybIK+0zD5lQUmepVOsYeKobr3x0EhKZrNE/ZAHpXFTvZ
FykzQERI/UTNoH5Pp7qlaQNoplmCkiE2TWdHeFOvWvxG3LBMAqGOWzS9d8ZweZoF
1sd8BMRYOzH0h9DRvPCcxfSmGakW8/cm2UVRBAWgyWqUw/PPywmGECVfDaYuX8Gs
QzOzt1KFZuh5l8R9k7iiqzRFSMI7U4ciESzGB6NpuLWsDsog5VrI7WGDiXDvfpBP
LJBpRgR0Fqd7zZEjg26XDg==
`protect END_PROTECTED
