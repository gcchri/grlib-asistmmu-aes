`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mW33dcIH/xxWqFKEduAE3M/WCk3YXqzUCH/qhuSprVtsUCAYM6gvZHqgT19hSMTu
evo0AXdJRwNgUBzGaF6dk12ApitsHSy9aPy+1DioYikjYPf+lECwisCUAwi2dLBO
EQJCBntNMruPt/9Xc1OVJfCK8QIGenQIpdvvjELBtfNb4B/Ui1HUYqsiMrXX/t34
5kfpBTRDts5xKL0O5MZpspP0qKPUAcwcOOkcre4QhxXjNkaXR/KYOH4U/Tssb20i
bYQ0O3Cbx1lFliwUygesMTboOHalKGUTQ0gcHhdywBQHZyMSRQbAw/R4r4aB6PhS
0eaSk9GV0cpTeVIRgu7NApAOwQjU0IRaDy8u32uHyYCYQHtcEfX8Mnz4w9frZQFx
b7L2hiljhvNUuFr193QfstJpE2mUO1r2o+9S6e0pS70=
`protect END_PROTECTED
