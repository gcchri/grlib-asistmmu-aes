`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yi7r/7fhYZVfF6P5Y4RqfdqzE7+vdcUkfAMMedOcjJKiFuvfAeVLWs5QK70kObUk
dunzSnsQPR5hKqMocvi1p9Yc3ZZJGWEjsTO9ngTuvDwIn5UP2JmSC+PEnQx6GOKc
BTtoRofxQQ6Hbo7YE2juyWP1S/r5qq5o116e4ECP6VAdl/UmLjOOKFXvkseCVB0y
UVh3HqeLYuVspic+x3NsCJWWTbcNFW/lOCqyAVeJQ58hbymyQBxzPldFqd4yGbzX
Jp4PcTVoBmI8BNMcapVl5viifWckYgfmHderkoUZoGKe1h15sRupHD91aZuShfOh
`protect END_PROTECTED
