`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BdTA2BjpfcBE7fMc7dkc7JLEiY//UANg/6NWTSiOgS4wzQCTi2smMzIB9zgQkcym
+FY0v+3af2nTCLnycpLaz36SLqZKK5ccFU0EiFLLBZyxsrHmB7MP4tdXRTcniYEE
oA9KnvpCgMGbcwry0M4hqM5tT5ukj5j/0hDxsdbp0F7kQy21uP4E/GNIY6/Pzu7P
q6g4fD1EoiEvMiGxHbUbOEnIxkoyFHH8qqnJh/SiaEAYZ3pBX7etqfR0dxTOmxw6
ncGC5TC1QOY8ixbBwCUJmx7VfsIaBK+OWmHA9gEL2oD+1wafTB4gZ4AzKrIzysUR
wgVGij5blWjAdQ6+6NlsRpGaq9yos40cI9rg4qP0NgpmOCJxV9VeMpw0eZNtInxY
+VrxYyAbNX3A0Ji9dYua7a9ttlV9VVbADkuK2et6MWk=
`protect END_PROTECTED
