`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n8eEqDWRoaYFkYMMyOryzShloTKEjd2CKfLBsZ8dJJZ+HrtezVCap8ir1AtfX+Q7
dAZkxJahX92L53rebrJkHu0rExjnMlADjqm3LKZ3CqDbGqylEaMMfqCyihP8ym75
j7pqSxa66Gy3ZE7NuQyF23OW7BWKI3jlEMkRzRgdvPzfY38FdK2JY5h9ooArJNc3
6ccz3rHq17YGnmUipabvEIhzfT7sEpBAYYFvcoNgELfMxNNAh0H6PRGJdsiwAFoJ
oSEOxLTv6F2/EdO7zBEVc82z1/Yhi+66k02rKR9sCHn6vggqlATCDzhCPcd91XRI
ujucLUgVVQ6AY1u9dcipltQ+Exc+5NRD05xuOQEUKeYWier/CEJG5e0G2+wKEToA
h8Vi/dJ4bjOuPN+VNSjshWiPjrWFCSCgFW/4QMBA2co6CoXxvwcFRqOJQFBQ03lc
MBB5yaaHs883g0jcVR20851iF4wLlv3s5nBA+omCUv9Y4Pa4vi8ZNSBccjE3ZOh5
qeaIOQ/3tc+Rg1MAb5IeDpQl91S3EhqNL89ognjFlXeiFWuQQM7mksUS+guu8Fk7
CyTVg0PfSkC49Ak6ZRn78Kz0DLNPyhC3OtDPWh+0piVAo7W2DM0+2YAtPC2gdpfw
Xkh1kTZ9aQ/eJJDzy0nWMb0PJ/ELTB2ZOPALlrMderx48hamogbuRQdWiQkgNKnm
a2+HtkoRdNFBj0326BMuYci2UKpbrJyA0A5cKdG47ZI=
`protect END_PROTECTED
