`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ux6ejB/FSd6c/LRdhLVEb4Ogt6TOw/xCQHKCfetEWJLj2B7JYuDgEkTAyxmZz22L
/ihNbN6dotd8E1O+0ELdT5IYAhnUwfyg8UdjL7Q3I67AkSYORKoiH56ewqiQthfz
T1s8qoIqvPf2isO1grKU2CiXcoVhHKaiAvcXshRdfQLbi82HVQ3KR6hPJubs0eO0
IgUg58SGXOrvyZCpE/XY+RShnVezhs/Obd1n9Hd8tDn45fSRjsYllMcR1iri64UQ
yz921AKox78jKZ1rlGg2BbS+KU9SxW8h2U4eFNh+gDmWu3SFAh8cDrsMfwtgePWZ
`protect END_PROTECTED
