`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vAdZaABhGRfm/akNGyXbnjbb5CggZzAuaizD8JQZ+Tp/pJKx91Wq6pdVfO/VkgZz
ydeaaq0LkPFggZEnO1vY1UeJxIY8nmMjiACXlRlioNmm+dneC7TOzlcRAI/6q+Vx
XCQYDfF+32MuO4VFNUvlrEKdroEObH6oS/KvvfzcS89AyKiP/BKRemFQMBeGPLMt
Jt6b3HizC0I5jgrFoDEg/UBbvlqxc4bwsGoJMA5gp9G+VjLxAaJ0ZQUm8++mvtNs
v5b/RjXraqChRKEnaPFPGV0OSKqc/hkWkc6osveorC195cjGelgmdxSCoLdp9M1B
tcvxnqCPxm5hGme2/qPtSka5DsSFjivb0DbuqAxsp2oFYlYLHRAq1zdimMMzca62
p5CLWhN8tYg3NFS+E02mYM9REuBSnyEM3wdvPh4RliwNMsAE7WrI9Zw6lULWKq5E
rfPv+AIkPbtsQCCC2qRlZEbQ7LfZuNFgpNC49q2PGlkq7/lBxpPs/QYEQAf7libw
2lsWpr8hXqEeVufF3QRgAvPjfqhBFYptO5fxngKGqAGK3dormaj8+zmASObwgOyD
88D6W/rl8IIHgbZ6X6Etbvp6gwS3zOQwRx7QAA5bWrI4HMhxSfpT6W19PkWr1BRK
Zg4613+biiHCGekEb1gYO0ZgBpkq5IhLt52WAudH25I=
`protect END_PROTECTED
