`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euzkSqNeyyau9lMnpoLecBQhLPnH8Ny9/aEC4OMwOaS8ZBuTSNHSye/GdsCRTbHz
AxVPI00T85tbkc7vy8Vqr5792chL5TI+pU9q7wWvuB66jiHPCOE5bhV+5AmMNNre
iLSARpkZa1H43TKB/8NyO2wy9Qm/Lt08xgYq/7kxiW83jwBCkAM8gNAZZx9Z8hXv
/AvhpeC2f7P3Dhl5UTwiImkWpDuarU+bEoIcTFbzYec/F6x5Fr33bmPSMpqn5oS0
pUCupnpcS7pDu/LNKsJM4bAQBRYripr9nizSySPWRd84sinIPRC0VdkWClTolHyb
HkTugX/ZSnSo191i2sxR01QjSzL/3QPbT6iul8ZnZhuk4OzSPkOlzj/+BHR4RnOW
TszoBsAQvex31zRszGDBp6doz9ilTq/RTK7d87QS4f0abHSvXLhvdus/7RLdHFf8
YIVxqbh1M7VQGarlfHWFOkLJo5lmo0YYYTemRhzeWezdefTekLU74bB8N3AMQjLE
PH4ZyfOu7ArK4+zfq+duwaer6u7mamePvd1WMBPuhT42z2OgYY7L9tXX3cCuSqnd
BqeAkZeeJfyPCLD50GyUHvwrXym2G6THJaHavTD96VaLSN4hPdKXz4OyN1A/mh8F
0N4x46kU4Yj6BMBdwwh+f5RmtD0ex4+DJH0KMc0arlBp/BrY+ZYi91BWM1MGnpri
YCpCDgT6TGob4nM5NdoKCEaSH25ihym14cAZms0EGWVgA6iqhhE+r1s5qA9usoCz
Ots0uGee8kkhFo5ry9typMZcwsNppT6iFpRl2wFsEvZrttzGsl28faulyxQPLHVp
M3r4jL2ece5NJIgP+1C0kwzVovxP2/PKI7ckER0yJ1GujAHVQueL5uGQL/SrxH/4
Ao/nj2mfyGilK651DrctblRubNRRbOwOv2ckhaq+6NTHN7ld647ueQ5ntJ3caAOM
gSeXC8t63HiDjbQTXu+TX8Tz7k7V7DwdWa6QnY/MzeQHwA/H06ar1FyLBQhIBSX3
vTxSTJ0lTRCh82lyn0N8oEBio9pQWItnXH66Q0QJGF9oKuPu1QnCgFawQzD9OFyd
mA/vZs9OiTF7pgUwljkoHpmz6EQNihJYiv3Luvklr0/pbh9yk7YDVpLv29PoJT2+
YRlKoxqcB+SkShIzhHdOX1gg2bDHdsrwkr1JGJsb6xGzQDNUj78JQUnBbDi3pLjr
Q6f1vN5xsAmSkR5jHbQ3ZHuikdCjYRmNqysCRKDxHdLOmi60oJZCMt15d5ieysfF
8ATuzv2cwjJ4LijNtfZRTTAvebl0B/S2BbyUiI0VxrVwItBVYDlMyX3iACEArGcC
Ur4Y0CLylAbDkNXS4HLK7Az0+F8Wlw7erHy547aZyHbFzhYyoAr5FcAUoWrqjQ/U
SoSkQH/WfsJ+6UhSTTAw96uNE0R1AXa0FtTkKeCKj/80Id1TD6DatSO1sXycRECt
G0HZr1WitctqCyAc+d1xA4Vs4Wwp30vOdW6gZI5C6txClJV4tM3BdCbRoXfR0xbd
6HIHwPpU7ThYUcu09NBtWeYqlwlh34Qp6l8OwoXSReX0qk+KTLkCBBUFR9srnvba
0dr0611dCuHn90Qi1e+zTA5eMKwrIm8LFbxeKUCcIYRx8S9WjwwFNMY52R9ECT6M
GJmj0X4u5s1ruoPbgLsfxFvWJmrQMmMXzMdUeTsShzc3gaUx0xpmXrrWmpFxZvKW
wbf2r2pt5gxA7A3tFEZtbG0TXqY/QmPW5+17MBMOG87Gbiq6+dvxehpp+sRJkGDT
qPHjD9RuzxdbJqdEGBZWLiWQKw+JwfB9VDo8FZVDsaXNvV6NiV8Jn3Tunx4jkL1h
BtQe+QgwdISaYRPTzLThQuEMnkyz3yH37yc9lFOsQQZZwuKObExihQKnX9o9TJgY
Z7PdjdiUAJhRyAIxxl4/TUuQ6xr17LQ/aRucgvT7q2T7ZgGjaNWAeFhfoMqkPjcT
LDW0Jo1Y7Oi0Js3REykuqUvoU+/ajcMxLHukaQ0LQ5T4I8SqFYaY+a4vKN8U54QK
f+74wfYiImPlOxvVcUFhAmA0/gGHTzwsb0VyIaUHwJn//tPwk7o0Q6hQc0/vjdSG
S3ny2Rx8Kv3LEOLIjxm2DlUpOcQlIUapdt2T42ryBbeUvJ+HRhotgTz/nF3cKByb
k4CJ9F7d+0Yg3thkXQRkCAZny8MVILSBDngys4g+sVq4vgGxjna1P2aPJTcrnGJ7
zvlLrHZRE000SCVyFAx+x7+lziCTaycE446Kkaby5LhoIc86MBFO5MipigZopDp0
/QBzfc3GnPUzYV5xMNcYxfU3Bd1jrC3YJUEtMs1irV0QmivfXXK6IDclzX27Et93
h+tI25KBpBNw6tP9Bkp7bwWXnn/P4d119DVWaHrwZQfnj3jKT1TlZ2iVmFhcyTgo
/20QLgnVOW//6Zf7JadYLnYN4bXqD7QFgkgvR5wKMKBLhNDHjBahhnKY22oixeMv
uk+JUPRhRBN7VrtnYMc5buh+A9iaBnheQ/qhs/szN/0wV4it7U+/umBhgSLcGP5P
dIEhkSkt9gUlYxhWX/18iJPOdaxkIiB6nFI7bnqUEaes0BJn5TumQ4TSDuwmGN9q
uo6AYAWUnprVw33W+VJ4qKvA2e+i5Oy1I+qzmg5FdCsWwFGVQX+r2pSK9lTJkryq
NJJSBIVd90w1K0o7VPmquBWCQijfbNqNoj1fxWFAns4TC5UfDhHwzL4QEi9XxTwO
UC9RkxqRoJgNbl1sjXIngYhOQdT7Nbc6MH7PFqzC8mOAjJ0nmIM+IhGVtSorvlfK
fxnxrVYBbWYly+Qp/4EyNnjYbD6Ued1OoC8C+Q4f3pH/vuVHK4+E+I9Qhe5X7uaY
eENTuFyC0Pq8oV5vge5d1w==
`protect END_PROTECTED
