`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cwelV0IAwaEopGBoYAwTaSt6K5moC4p9QX45OFFKuArebpAoSi4KNLnwFi2ZxeVA
ixfmMFDkcztnPqixaGbVNU3qKQJCRMYXLQYg807JOTaOTOHRtZHpJ5oxj7zV1mx3
ZWW3lnxM+ESQrMAhu920UdEwdkrek4g3XTRTw3/LPszblv42zWE/GXBQL0nYokJu
fK3994JnArUTrwPjX9QhgGGqhYfue6A1n3QlWybAjx6a9ksw9kYpa/kGTrC6ZNrl
nMWp/kglg7+cR09AvADuth8a4bwU0mFLOTT/NSet60ny+5P2eS1afJ5ytuRO3Ixe
CEox88YrYgteBhsbrzKnvZ1qzhF0cjrPf/R0iME7p0T09c6NHLCRbxx4pWAoLdzT
LDJGlVjmG9j4xdQzbOoAh/fiCg5AZvyTaZYG97E4XhRUDfs7cWNkbSC6ggeGEx7k
4vjog71hpP/f/QzAF5FC2Dq3yto9HMCF/RCZYpR7itAerF/h19186CXFWICjcMb4
GRrl0KUJ08ENmZ1prDFkGFwFUteRTKfsL9+44QPaiu+Hkxq4hMcQSJTkS/bOXcLt
gYQPOwOfJEdYe7JCYNL1EZLsvSsCK4xOQrwtk3+FclRudcLau2Pr5ioan66AIKu+
jImMbULT/QCl2cOWVFwl5Jn8dPxlmESDcHgD24os5g4=
`protect END_PROTECTED
