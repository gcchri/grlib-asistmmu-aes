`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMGxkHR9s1zr3udc179bxxvQjK0I6TKjmAJ/WzUYsYpdxMQNntIJ05t5OA82UrLY
u9jsIH4+va5gMtJLVgGck58ciBowL2hJDi0CxVgnri5StCaT3QoLzDI9JTcaLMo6
bBuYc+ahf+D1A4NKKgNLoDmAQ41PLi25qjGJLrgNYQitP9fpDcH/rJ7XdpLPnXR8
qA836quTEuKDG/zqU9l7Y98r02mdQxnzJgNkrAyKlwpSp5yIaQDgG9vhiZ9eEqFA
tXOCPIp05bkHKpWQFugjA2Oll0GkjXLjeMnwsMDkvAABEav6DuKk8tANxTMIDv5x
tSz5ZhVjTax0GO4TPoDjsg==
`protect END_PROTECTED
