`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLXpSkV3JCs8zAacn85kvg/mA0kIdf/sLWDJvF9xHrkDh9sDVWn0zL5T2PdKHTNw
jhfOPk4nSkUE26nxoDT09svDZvaF0ZYAFjyZJ/mA0f8xKvyXdROit8SwdKfazFB8
lQ8K+T9IlZSgJGsTINqRkl8reOwC5S38GjHLGqqcFKs7Sefby41wqru73W+bE1wx
YAa3LbK6GzD4XhLvUpS4eRC35a94iPPxWpUs2Wqzbn7pNz+ACTsUHwcL7berCLdS
JDckF9orMvwfFKq8nUB2r3irinvPliqpgdcfj19uQnlO2TgAchYmG8dHra7fXG0E
JuFo61tVjM9rfYyGmgse3mTTFmght6lA+cXLzUK0dY8TU9tJDKTcKbLe6QwWcmiP
EmNkyZYQ5ovfVCNY48tqiKmt6ogU/jTI8tUOC3gQKj3DL99DCNoqLOwfsfXw5TKt
`protect END_PROTECTED
