`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9nJRN3UWYnU+q2x+tkK4aej8Hd5Pa9Mi2J/7dpCXhIcIxb0BZqPi+gRdvstybJCF
8IMKqUfI2LM9r6RI/TPMEgtUT4bzyi3NtNsOYz9UcJtWv/MFpKB6bix0YYkFeEnI
mOrDmMilYXJf5ooFAJr65tV8/+uu5uw+Dz7Wc6tTfiY0Q5TTRLBqXdEn9Eb+WoeM
dTE8wGBw/2DeVFPpAp0EzDzlEjvNwCR5txiqjw2nGRcS5o1haWcaU7Cdui5rMoE+
aigJ4l6CDKBkVH2nXh4gFgECA0fDDMpQ4U1sd5qGSAL9dK+iDIU9M2TtCd6vf2Hv
/KayaiMb4qzCLZ6PNOodPqQWvhJZX4Vu8foDXZqxWeY69hb8bGGcQMQtjedVYxnX
oAYyjJazzaFsi3uXYfBTcX8jG8ABF4agAE3tmQxozujYg1vghPjLLHkqQsysVMAZ
FDYizGsTKcewTNKp7DkSRAbxFulkrtIzj1jGSmHYZ2o+Z87ZVs51uldpsud1QAH7
vf8qRD2X/fCkANkAbi0BPVnG/fT5naN5rTCP543EFjXYmbAiVnf+L4s59w+1xPRe
WXu0dpoF+7ajt4WK8wYYy7Jw+QhWLER+zKQhgBcq6JTQeYnD0nrptF2B++5GotP/
wr7XN0/koiZe6OV/Lt94TY5cY3Yvp7VNm65B8p0hZ9p3LQVRUcHa8P40GjftGWqr
nLrkmpc7j2Cfm30FcI5ZEcuW3Zzb7iz1L3FIyW/Sa72u5kDHJ6t6bXYacMxKWaev
j6CBD2GoWyOt3eMjCL99irLigMXn0Jku4A+yUQP6KKnR06o6XnaeRbY4+o/0rAiV
RzOMK2VZHoM76xURtub/Z/1b7fxOpwVQsJ6vr9BcNt8rgfTG8P1gcPnGHn45wIdn
0GJK+59+wdxxcUZsDh+GXxLFoPxegK29b8KZmSqDq7CISNJ2furjuCN1E7PRKz/z
kv1qWZe5LNnrtmjMClzABghDeMtdzGDDkzYGl7+Nij5Re/5rmoA7Y0fImE3KAmVz
AjZJZ2QqOFeiA9ADPO8UIrfS9A4Z0imRiNb2GIslfJtQoJDB0C9h5Rq8axK1CQ1i
sYrsZwFX0EMqTw9wZZkRqKUixM45fjZV86BDbYhVyk505Lmk2blsnvYrvwxjv0FJ
QNezU1BPXvDKohJ/gMhIzGhWsr1h3bkxYgy7SCrn651u6GKUe047SzV2BflsxQJS
to7kbcEkba7rVP4Aa/K2ubdykRW3Fu3UKgJIybeW+Zqdb/hYqdosNgIocaW7uWOW
bSxzOERKspIGiTtUnOkmmAV3aKJzHq5mrIRRXjuJU+I/78doP00tUmyo5vkCsRoO
No8exW0BKufnK0lviVu3rU9htNvJ/8DkqZUQ5iqlpDN9MuQhqGMMFbwUBtr0NZLX
9eJRmd0MEnVqQd4+nAAx6A7akMNgytlHjQaNGBA3I25zaoEkJnWXdU1hCXqLCRYY
hxNPukJUVfPKu+qfDBw65acqEWf7OhjEmxAjTz4oreo8iciWtQ2nkx5p5NhIAEM8
H1C/WHXmVzmo8ABnL6BBBVXcIJj6cQbObWOrcxQfl9hUjL5ug93S0PhEtUPVii2W
kGOmkuO5z+iNM4sCf4D8xx7M0mT5j5xOX8OaSPrESJ25/RC9CEXITc7+5FHZI4uF
WMbHjQqpol3tTkqitTkl5b4yfshkiw8wlPH+PVMve+NLdVUEpzngCdbBkOxEr3n8
z3pMm6S/nsgWvt5HRcGHAIej27iXBlAEaT8T4QV/RPzaxYhmmvzTil56O9tOBIhb
TRD04XbwHi1IgNgi7TWeEuvag2mk4Gmyqd7caZUZ1YI+316ZPvmktipKGu5oBDJ6
WaHdyAv9BB9jveh3FM/WLOTK2h6nSwMpT8Hveqix8o3y6chKnL0YKHu1gjg/1AcV
`protect END_PROTECTED
