`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vcDSgfQ/Me83brrbvGu4pKsAuBkot6M4wvTUsY1uCXNe6vYekVD88cctlmjAlJza
BmCilTI7HoW1FzK0VUo678kbvXwSd/Z2QLyEtkED+1JWOKV49J24C+MRHd9m8jNf
znhWLZajh/D9LnoawVyDW6x1hmdkXvbpg15HHS9YKwtOQPzR8zPtlRdy9s+LSoJm
9PHwplA586OOst/PIhIqaF7Uu+zH+hG3j4w4DfIpZ8Iorh2amOkqOOQ5Ts5NaED/
SxhugWNKlXLmxTEb/SWhBsSoXWruWZr8tscjQSVEFX1RBTnJNvjkBY7ANmXReRV9
I8Ffw5oXWEj2qt3Y9Bnp/uzHy9Z7CXOC2515WohpknOztR6FN+c7rbioz9IH5gZO
3zPidrCfj9KOwPIiR+QNVNWq2HSLCP2xe9lZYwI1YyM93ixcJTASTaEaz/Tsgv7c
KAWhFFr9uP5AvwYwyKqGGPWrXD4NZy2Tl8gvBt8UxkkPqtiYgyx5xB4TPLAdepld
pKh+ADY/OD9PIoL456527pWGtLELLY8K0+znnII8N2fCjHFkFR9OkoU6CVfJj+Wn
0rR56wd2V2JfoUkAibKoQJ2c8gYA7vpTmq890wD946d/K6CncWQueukhmsjFQuhM
+5QCcH87Ri7GsBvmD6mCjchPueYDTn1UXXv3J6uk8IB/9MOAAaYYKUKBJWOgqqK+
YQzNPRaxniaCHD4te8XMa9qL04dk42rEQGYBEczpBuD6ABlSnw1g5fxPUN0dScRQ
fWvRkWgpDGgb4hhd0Tiba37ej4f5kglS8dAu6eAhrZ0dfL0MRrsbARGZMGV9+Wkp
FeyNftKB0NH88AZefMPFDgfHN92mwTPFvnqloyhYxAqR67JxWpdOphTs51AhsR+5
z9nTzSRa9KdZ/4Lh0Ra38pznape+LFzOyc6CWnJZm8u6OlyRaMhxbY0ZbfcLErEV
VL/edO7dqSkoaLSD65Um+A==
`protect END_PROTECTED
