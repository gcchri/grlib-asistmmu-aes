`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBXHWVv1r1bxIEfwm+ZV5XNUX6CvtsVvoWOO4HBXR+QceaEzMgO+727b31aawE4j
+PBW+g+VPSqqvo8I29wawrrGN8fBbEX4JNKBiaGmACGkjHGfikE8sgz6C3yPieLn
/J0sSwQDWEA0Wwj0aIt6cTOYu4bYb086y0Cc/5qHdiRK30/rn9AouEpUmKYb6keH
bTp49z4qQoeY25kToy1ubz09EcbTSmXNALHDs9+3c+TipKph0uZumFhkOV9/f7EH
ym4YMhHHSBSqDy3ne/C/AuFAphpVEzFkalX2WaLjcBbPSFifJcA2z7qpaoUZB23K
FbI7xIVYhJTdfYaKoKgFeRSravc2lw40HFGY7KdASNI=
`protect END_PROTECTED
