`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nBGDy5bhb0JRQ9lGrneKvspHClvWePIteQKs3t0MQWFv5JzM2z3KZ/rAomesIH4s
XqbKLb5TL4DoSgw2s4/gqTIa6N848wfyFbN9lAhp+hS5RMaVCJYYyDWxhDX0zIaV
LSN4VNBBCRsOQ+Np+zHoD9tFmlmcG84paBhowPjAP6I1ViwunmMA3HwC1cRl7G4b
jiAJ9zxpggeY/cDQPOhgr2sq1y2jZkItnXgFoay5JrsIom+DtY2IBoeD2IGyuS3d
Gr1C4CPsm4KhpUe64HrKuv8D1G1qfG+FkiQM8VDanWHWu89csVetIiSrlBAJ9xlA
OmaqUCDdhW3NznzWbg6/KT5KBBmLThrp99y0ghnVy8CNuxrjbrevvWqrpUhzL6jO
+IiCjkWLdzKP5rpE/GAYsZZAcCl+LOvZjE1cHp12vmDessL+BBjnmprH0gY17Dje
qDqstloLf8zQJ2CLjuXHoFF6esBcuJHlGkPzHo+XHro0S/6moxUqpCIGx8pQsm90
`protect END_PROTECTED
