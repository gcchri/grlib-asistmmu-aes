`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhG9lb4Z+sdMLJeX4pono67Aln9ysexeQjldHsl3/rHjKVdKUGKLa3MFjT/0z1In
wbcD9up1SoX+CnGG70JE0AIRPEU5QrV485PwxlKN6eVu04TtRe2YPA23dhLpZLXC
dEUATIzxMa6p4QDQlVWBvzNglHKpGQIwLHr7L2RBl7k7vIahSHyFbU1PSBoQSdrM
jPVsGQ5P3uNzRu+1TuP2/P6SONDVDfUoBAIUztuK7GyXIhxTJCNesKl3mtPwXxE5
c1JmNi2DFHQ69fMnS53rbzl5yh7vitWVK0HDH7yq50taNA9Uz22I/3TIuXVpFpyk
omgSsJ6boR+fJZ66TSdRjjE+6xS7ly1khBS2TiR7KrM9BqwEnTQkxIwc6OB/+gBd
fw8L6+PzITUfUki3DosX9vdzPejba6GH7H47n/u5NkBqRk6zc8I9T4IwQMpfHB/j
b55+zqc8JnINcul9Wr8tGNU/zIquoGiOxK32vrsuSGkFdaDj3KA8doca3WwresPv
wMD4NuGpQHo4oZv+tRHvx4lm6dev86P5CYIGbrvMC/r65kL2eNQaQVo7yBQtV7WM
ej2nZET31ays7tmBWra0nfaGqxk5z1ta+tEIU6Dl3Xq7AR7J4Ply1QTFvtRx3gDW
88e3i9zHJy6FFx59PDCvEkFLJEE7JSdoZHNfqOxRCr0Ym/myPHeumezKqUKefJAL
/bkTHw33l3ImdevlF6x6ZwdwicLMrLIdqdaRejQXPUeA0SbTMVH8bf73Vz0qJJYK
Akeuf4/AD4wVpVk41UZapv80RDKcr+tQDUYwGjXB5EjNOPvFlv6Q1nIrdY+Hqrxh
5slB1OLPONclol/TZFfYpV0N02aqAogoqxTuRO4vo2krRN4qe5xUpiyVN63KErr2
lNzL/78eKEGTQROWhH75yjQTMmTLaMfsVkDk+mSNNxtgtHbVu3MrYNw7MUhQSJBc
whRtV6RHdPLmnBZA8mOomc5x3ajh6rsifPkCMLbLXDPG+LHNjb0jAvOFbzPKplPX
wbRUAr5JlGaVTa6stsRDmqgWbC8xWDwM117jdwCTLVYYN1RtSBKHLx3/KTkZSUgY
cuf5mtmD6SvfmcSVwThEsk2zO6IRJUu7+0P2TrTu7JGJp32siQR7TNXl/np5/AG9
8w0bLrMCEydX7/YxS0SGiuwA7xxY6SgrzaGYohXfU0Q4VKOa5FU4DPnuGqW6MS2O
S8vzsKpH5gEKk9TwmQgnscKgjInvQC/gvUC2MUf9cwlVYD9Jc5/6I/s0rQSg0awC
qJPSpQTWzCQYZV9PZakG9ieYh73TmPMxGrJ6otzIlOFiv6ouaqM4GrNp+7iNNUFh
7Q/p3LUxd/ZvNHV7SVbMlf4snR/JOvrnzy7LyQFKuXeRiVJRt8CCw5AlWBk2aAxI
ddz+5eC/6MAqqgEHG3OqlEBBWg/2rkIMUMbaLRWr/0W/OXWVbJeoYA4Vniy7euJT
`protect END_PROTECTED
