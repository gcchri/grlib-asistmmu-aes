`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ag/cSfwGNlFh6KAsGDbwjBIEimi+RBA2+4At8NKMIeFvdsNuMxOZBKupaOAD1jfB
an5DFwaMe3SSB0NU//SY/yEJ2tEZqCjCsk/1q0l0LLVds+5hJ4rUVqqNkxN0zzmy
yS0TZYZILW7GmPZKTiBsJQHWNWXymZ+EQY1+y6oeqkMQ/xq0ei7Au2JJHFlP0ey6
SrciShmi1vqWehobN7sGgGXD1GmHEFh8oyrnxPvYHuH9/b0Y+mMHribe5Yhk58HH
IGRZ1LLoe+bG8Zdo07HcTq7efuq+FSCgVosw4EhloAr6EEv/bZv4sBkufLqStEgW
ZgJuCcDYOI6s7urdvggTYRGVXb/vKH7x/xxj8C1eJKSHfkmy/re7kAGvJuBww2m/
PCfyordyp2no5TkJR/UUuPgahuXqT/R4sTr9gZTkA77BXtXF+mrgMAU4qR+KOCbw
`protect END_PROTECTED
