`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BtR7IDP9bKiLLtugCk90wGQFpoBUt81x938Grsd2FHp0P1/SmxwsfwfZo+GwT0q3
i3glgsU+ZbMulsuyXJNwsWlNOfjCUHBlZV2nvRgYyICxrmbDRcOdKQRTa+3Tnvol
E73zrZteSZYAIHzppXXlInl7GvD3bknd95IA+9hgZTdCncApcYOLZinDa9ikRgQw
2CAUHbBNet9JIZqI9YeAM86KOI6bZTNKJ/iACTFBDI5S94+srnvf5yfl09i1mikw
QRo1Lpop01iHZTEWrT6KvxURj192D+Ho2Ph1h67/b0eZCbiBvwhMF/YIj+hFTc+4
4OGYAULfjEw0H4nABwy4oqBlDDvOEW2Rt8IHmJooerYI78aBnJuC2TQDrppQIe6H
pazF8q6PEgb/lFj6ZXS7nssL7RHxLcgKmk+Xk0zAMKg=
`protect END_PROTECTED
