`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pz3Bl4ohWT3pMfotzSnUuLs7oqQkzJcI9251cCBwXnt1AitWGG+h8pKm5qjuNzhn
BW69uv5sxKL9qVXpOi8S88N1AS1x9WHPe2BwSXUek2iuVafzUWSdPlE87fX9dHru
IQRtIL2aKItJdEtt+2h58I2ST/aM75Sin1Dqrdb6uqX1AyG1ciHrrnT4Q8mvWIJI
PNbXwYrrMORSCkIhXlaKEQle7SrZUKpn+vhdTJ8Wj6YC0Uo57UdSHiLqMlNjaihx
4k2AfUMRIybnh059087kmDnyFju3SAoHDz8tlvYDVhlsi8WjBNxXLFSXDxopVNGx
f43koByblumdA+sDZ7G/tHnTUN9/1u9DcAjkZlyQbk/AcvIZ02eIg4jTyy9PBcJD
O5LPfEgqYRHNm4CHnvlPI35wT2MsDV3MbHosi95e45rSC+2fRYPEk5fME90JaBtz
+bvb9P3WtyurZuwBwqGyhCGgkQN0UFFOLjNA0AXU6tBsFgYkX7h5gpy9XADQqHsc
`protect END_PROTECTED
