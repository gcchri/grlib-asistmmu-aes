`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bZOHoHB68GCul+YmW5t+swPLm+PgZC9tZIXz4QlPIEMKNfwFSYeywQiVUdk1en9
v+9wtLxs5uTzPJIYC9N8IQD29bzOXwsfhgxeLJtXMup5482sCvW6fAZuKsit540l
JxgPh7yEI8693jB/UFumPT8JuL5E9iLmRCpCHBhDhDKdpVpr7GpS2KLOscdJa9RP
FwSM7Tfoyk6LF5RS8t0Kei88dWITbX4R5hZ7sQYH2HTjyOrhtcdFNcih5gpoUhUI
8fMeRtcJ8ywvw24D1zn9dPv/Fm2N7TvOBIDAJoK+11jb+uOzgAcMr9k4laUEarVd
5jm9sczmzLFZxCIxuihm8mJcTaBpIM+J2ZMARifZ+Aw2ZD+c5ALmtcr01d0D4TMX
y1XqsNRfvNgtQ+VNxSzMWY4Kv3Xbymbd3OhnqdKDgPoOvTuYjHtKcWz7QOUHCDD4
5gTbXP+WZS2vaoygXEDUIvfBfJQDSLKCZ5OHpuz8yDyJXtk1SuH6lZidj/dEDmmj
7wKOMmVGeQuVSEd86dxOTAQ/JHK1+9xqZy04F6z6XiRtegG7efXNXOQc74br1TjM
gdlWPdZKCb19zGVqQ0IEK4SXN6cuiGg9BT9jvZp8Egw0SKAZA1o8JkPdKhKCelzr
vbhDkSvQYrTckFUMv7c8uiKYfizBAvqQDVSqnDrSUS/910HQ4I5vDgbTB4GifU6w
9MGIiLyJUu5kcx6p3pvChBvJOGOK4SoRyvsZnwWgMFk4ZcuIIP0wmPLoqSvKB24J
VlWSugubxQKsI8u67szq9jX2gx3pKztkcPIRRbAfMGyDsp7OV0ffiCI9mvaOGAOd
m9R3ZxWuhrf4SrhzFSttuAMQqbWLCbHm8qICmZl2HswRSLeh1CoFjpNF/6fEXzXJ
LNL+oT3s5jyIoQezJfkar2Pcg7JCdQ0ftUvvvJXLoRpJ9m5blXLmoHSYHtCN8jOp
bnJTpxeKCPhblcKypAAzHscIQKyI8NRj7TZfm8OBfemn7e+dC1Ms3cDFqh7L9Gtv
AGGnEANZbZZUSK4OXSXQpUjTse21XOEDmis0Q1J7ZjzD2pzB4fmV1HnlxTES5AHJ
dzQIYHdbW1zLNCPcAwQpSszoo5aiF6rUlxWQSC2A1lVidrvz2kpNn4W6BK7iBQZj
R+LA72DZ8b60wYZX78Z7M8bP0wQsfYNwxsD18+DlAOCUk0IqImAjj7LRPVvQnfeN
LhbOOK2Lif7M6iB36mtJ6nCzAKmo9BG6YUlpxZT8CbxWqI9dkyB5V33Fevz3YCtF
sfO1k+a8nSmWAP05C1AK/KtHxoML+AZm1NlMg1JDq+0udCIvgCmiSsqy4SEzEdJ9
MOXWf53uZkUIvc6hUbxnjEpM/2rtBl/ggmO2Gvd5tLKzMFCBsFkA2ZwphUUUgDUW
N1wTAx9+esS4OxZlQPAjVZAt05lmiZfSWah8ReN6GSJ6IVjfhM1RXjhxojrRPevw
wE0fVcSw1JXT2TUKmLXTPH1lbVexdLWuHG8CEfof5RyaCy68M9xblL4/oxgNXk9r
Rmvdt1V3kpvqxwWyEbXinASAAtHTHHWQO2lfJS3mQrRj1q3oBIauF2u42j/1P/X4
4mjBzm9KsHB1hFEP2taZZ6NhEenDUv09mghBIngZpeons4VJ4HULVBqCG/ix3ALq
yfy/NG59bVaWw6GkV38pgENnOSraG1NnK16zPDUK1CIm89e4fB8nfdjjS0gjqc7c
J1k84ZW6z/e5fYjQ3Uyou9Eg6gRCQnF8myOaujMrrvokFxtRS2wW+IyxjewD6j4L
ocpbGivo57bHOrpBQJGKX1BAsw46aClhw16A4lva5kxiHc1jy8hmXA8m0tzge1Kn
zZEtGZtoQEFNyAxhh19ReruC++HH6e2brMnoEi5tcJ72iecrizbTmp2iLU+dow9k
XHdH8rHdVLQFYgNoiVi+lne5WCXWqy0kbTyYWWNr6YXE4Y0p7RBVTJ7ccUFxKfcO
04H97RjRJ7YqNyEmrTbeI84/a7U9J+CimX9wO0i/FzRb3u4Uj1o3NJR33fIPUPZ7
zRulse0RUdrBw3yygeD/7JDp+7KpfUbCuhf9wREdkWZpe96VS6rehPEGoiJuozBh
XWcBCJRNaOsBo6mjs4mxAyRFxiaoqj/sGyju+lQTDMkZicnxD9bYRaErlSlEgx77
4+mD4A+WING9tvISoJ5ecJOcJt9O+QcP3cx3GkHwADyoLXwzqEYF50lXRdiGGFJd
ShfJZPiDM7Qyf/NUoeXr/FlSDL1xKbdIgAxqMdttOFgxozFCfS77RfLKiIaf7aTL
zyHnDaEMaqZ7XfPXyV5ZKA8Izi4tJZMTiXWDZYz4bVtTjtHFbIeLjdXiMvyyQpeN
2HZhSlCUhDxHhTleeEga9LXNENrYrlQNPwXFMoKlKnioWtK5HojhrXKy6WlUCgXY
Xf2sYT3Rkcp31OGs/ru1vZvd7C1U1BvkEcvjeREI7xtBkKQb+FDofb9Z0cMx0FwG
dlYMbZ1bw1jicqaz8z5so/GQwgzt5Th9MTxRawZ31eCQNjeRdYJ63QcwbN0oG5rt
d9n6xQckVQzviTDfPsSMc0ha8cKzQAw+yQXOnHEMxGZqq82MmxsxXr9dJSo2tXgi
CoQ0h/jGBCoLqR3zB2cZPGJ8q3qoNfe6d8SO13wHlNL6O2FKm5B4o4Ou9gGjjA1b
2KphlqBMrZXTg21jMgCPwlBbOPZRSkztzDu2eI3gZ5E/gUzkMdnVYm5j9ywnvXoR
e2nv3n9q1bopMnY+oeZqGkacQQz7GCfh1W16cdP8jrbLXGOMGrijKBeiCy+UFVOd
D1mOi/NQ2DiGLAyijl9CEC9qO9v9fjSwooOGMnKisNbB6BFaNjrhME+ndiWR1Lrl
x9L0t+snbbescZYl7YgifRYhJhept1GfnrTKFGDjNqdTTLzpxpLqxLevLymt14Qg
oDkHelks0Gha5VPER2+sUf1u6M/TLpeGlcq2m2Hbc41iPA5gvNGhDiYK0VPx8o5/
5DG62TBmzlmqLxDn6Al7z0X2ZBFxsl4BS+ex/tEJXpIct2aNuIm6rB11IMu/+7RG
R4r39gr80l9i+D4SeFmZcgxNhaYVR5MP1XjD+qcWjKYmqJ95QjuTZRbYjM0OdO8o
LNKwpBojVJRVUzXxi3UKNkbvq4wFUlc7Qg9znBHUHs4j6hpR7t8cuLDD097jfPEq
th66tmpx8GUuuNNHteuGh+oKWwWjxbIqISxW3CxMZNKRPDwAL8ry8VlFcSWV2YJi
jI5SuzftClFRrdKLxfjCb7eh9Uarnr7NeM0bZjBJZjjaLOQ9fwJ0r7KpbjXFdPrb
kkffFaIDtMCe8rWsmGjOHgzUkILnShZ3+1AVZ74bhhvXRM309vckqCvuQLa5B7kX
gB936gedAIQ0F6fQUDrFXE0Y9SocYFcixtAUpfcx6kqP/D0Dh5NHVxpPpQ3fb3e6
pGas1pg+H9QZowIBVe0l0+UZAPH3nTU54QNHCMfnC+Jech2OAgQ+abaIP3MDzYFp
deoas8qvbZA7tdB3rzX8y+h33kjpyGUEFgB6MxOj/kqC9I6uFwwAsMoT7sun8TaR
9FBvrAkS2y1NT+pCqiu4las1LTCGbeaauWs2I3E2GND38aDMvMg83aL1r6MaREOK
J2NXaOYmnDi8f8670sJz8zhhJcQVX/k+RykImjCks3vTTYAkeHZRdlvxFiH1XNkU
geQruXCO4p4NdOz9Vygt0IBIP55O70JXY+rMCpVZAqha3CMLuy1mFAUS8mlqY4Zh
cz/VKnbviImjf94863sUhYBly/x3rnrldj2EwJ4E7/MvEXvQi3XH5m3qeEzc4ULr
QbagMhxFFDyDZvYGX2Vai7mzTia1MkAfvWACrLFo5rrCm9j9b1sKswzyjA0vCzt4
8gRyxL2crPMoS3SfFfVIklMaQVTtfSp44dazAJlwcafstBIgDp1Rhw7u5b0RIPAf
OUb/xudG5uvkGGeO1gH+Fzl8xU1TwyCTTXlXSwIXvgGa5mB2YsNUzS/Waa/68FWx
Xt65Gw7GcO2SHOA2gZi1e16x+MbLk2gnpArBGvEAPiq72MKY1uCxfZRIESMuAWhZ
Kbu2fAmaGYhrEwT/xnOKzEfJlxi5ZzxAwY+aZfh20o+Bm2R9KV8smsawHFGUBfpg
mVws3jJiQujQXRejY149DrD0GCOSeVxMZwEdrFbNgmby4wHoHr9URK0ULU2P5cHJ
y23cddGXXk+AazH0RNodAkTt+klKV07ka/Z7SdpnLr8v7Fqy4Gif4U42uaYXGb5V
okamRWFx/1iGOWTN8IgOSVON0ygjPNnPkgKZo+BrJ8TFpr69hnk+UDDy3wvTvvLY
oeZofe11qyhVU39HAJeEb84GGz7GBUtS7vM3+V2IAuj82ykkGuCTBpi/ZEnyqlv8
uOubb1bOPgn+OZr2imTS5bTolHMD8BJDQkRZh+7LpwgE1t4TnNdO3RjjI4Zclrfc
tNnvGgok8FfKJAifFWbEImtYezlLJ+u0Axy6kD5WGpF68G9rDZMUidym6P2rjwKG
y9Im6CnbxJL2jwBxaJFCmbj21T7mMFXh5E7jKcG9Kjkc98KY4vbuUxfrkyxEATdF
9hxOkvTuvTd4xr20lA2azbxT7kxXIn4HuKN+fBPN2ULPrw8HHTxW+lQPbdTL3K1n
fIelVpnogGZ6spX6i1ZkQLe+tEKzYPUa6XjF5Jd1sQFit08X2HyttmfLf80u4wxJ
sZgfzgJlu9kP4Z/pT+A31uVPyeF6030WJcUwUQ9/a8zo0B21NwEFDVnmBVH52PlV
4BcpCETlwqqqc3lhxZQjN2NcxKta+1n5/ALlDcJSNZa6tlSTnUUM9Ak8QXORUQmm
TOPYv6UWju4BfPk5xdoa6m5HXKjfHMBuj6bl/VhO7yaAM5y8sLfY3IJ7QAvIj4C+
1xPT0ZRadgrfh4q1ZAjm6pDKeQoYrdrxles6uDLFgBBjjv0xSh1oG+n7ifjcrlBR
M49f7lU8NAJf+mwp5KqZ/q2GvqeuYW8ucfPGw0qUUE+B9XPK/z/ziruNEb2ZPUSm
nKQG7FHwGxAWt+e3iGuqUTrXnj/qCaoMWydmwSXend8ZKTpVOBa8nlY5tKpIHAK+
D0b6refjIBS3QOHtLa3r8Ej8qZzelqoFuvkjErRm9oCJcuJ73bWB1U5myCxP+Owl
TeSZzd6yrvWUDS4uaksqBvKN3zun5WgIQ3qUexzpb/pC/Zeufzt+SZ03/a0xRcF2
lIZmzQTwN0ePKXmUzO0vSwgvSLrNKAG2aTQsCueki9gLHkz6/xQmcnwFNGxpoih5
1nhPHD2JwnsOf1e8eQHGGjmLovUIKPLcvMl15f9lPf+o/cE2NkMpC3bF0wGEZVIj
ov8TdmtVgbUDYAC5x6rWlSsK00fbjVK0VmiWUyVqPNdd/MQYmaPbM1d442VAmZg3
XJdrBrdth3+12UKulCoupZhcIsLYIchnVtvl6IMIF2D8B5zq90XizxHZX9I1wjJF
bOjyoQFowYx4yNA2NG7dHDAMrPviaD5Aq3vBNAnKefgpvFkMKRlYQHzlbe2QLfYb
Y4NdJkq+J9uYYtWpFz4liTCpGQROHzsmNpvMqdj+uNul/VTi1ZklCaVuJE6NNgSm
Yqy38fD/kOoAVj6CdxkR17orciHh8ZCccPj1Lv9xDGmZJf9LEdCh3JNQXrBow0PL
pVfghCGjoBMYUX01L0Tofjqd1v9392KW2I/87K1MFyWUph7H8JNR0EjvZP3uHx77
mABWIq9+WmzaIv1Ta7We7WiCGi0oM2N1cNYyScOayerpxgpduIiuhbk9k6ur9G23
U/gkW2ReUmYkf5+ahsdoavyBkfny/ncQtCaB4HS7Q1adojoNMWRYfR6rpg0Jzf4p
4UffJxVUMiWt7diS9mzWaWttOK/ix8dR057q/qWEvo3qNgjYZCxgYJANhMgVGlpf
nqxx0fHEKYaiebH+eug9BA4K9vEfXP51lR8kqBLENAvCdMwuwSqtp//fiUSsxWl+
5CgSdGH2RGKxm0nAmm513vGeUT7YVhoxEAq+PDR/DBiYTrJiNiYiuId1MATxoVBT
Ls+2yftcy+67wBcZ4NxLTUwGAVT4rz0+gnP31g+kzEkZ8RPR8+TFGN8Xc47pt5KL
u+BAFCZpgt6nvgSbei7B1PlFbvT5iR2hZWAfaDOC2K6mWUHPdlGepNRUmELvpxj2
5aZ5RsOAscyfMlk9vvgbZbkPU6Y3fQD+2jpaxe8FdLOBNUmBCItPmqd6Daz21W1t
Z32oxu8Cc2m69QoswySUaUftfdXNyFgIgav6TmRVNecD1mr6g5zbzDd1WSDTaYgC
wLqICU5QWty8WKU7u+9w8w+QisoxjgYyl7u7jrIukutkrR3bM7i3kORs51hO1s1I
suPNXF/SvVFasUn2ikfcyXzN3VgQQLmoufX8ci4uxSQ/fHjDdLBvXubmLz3FBs7K
jYkXUM8MBcsTC/jdILunSlK3Uw5fqjWD35xzTwq7S0MiZ5cSAxb4osoxVTPXeFu7
sgMJcD9B0iva7JTjdkSC3Te8vxaANxg6hT9weCD9QBmzUqCuZs8sN4CXRjMEGVxi
x0uM5DnzVi56wn/x13T3E6ZMv/2iXSs/XcywjscLNLr0uaer5Ee2P7pZPQL+2QAP
GLlz5UFE0C8l7Q0QVcD0DkhNan7KTLZREWQ0KsnY7lC0biSljWUxsQ1YEaNNbnbp
kwrNcPM1Ma8j3M+PXDnUfWcFAo1Itq7wqybBfNKoB/8K7kWICasf9MeAiXl3PNNb
TMWaRn+kgNZGMpPmUdplKNut8/7hAZTKKnHBuLDqvjPF/8Fr+VusgmewhW5H6nFc
RR+kY0X4ZE8Ob4JEsVLS+o9iGwT7pK8G55VWzByIIQBZnjYyYrfs0tI0G+gEj5+H
YZAm8OUNKu3Q0vsi6wbfakuMoMFEVwdgSCeJ6ZV1HzWzo6ixVf3SAFHvCCG/nL6g
+T95zBbwtQiwQiVZdRzgXA4yZQuJeHXFGdPDC27vSZ/xQuOCo0/7RZU1GgMbHXvh
f8sit5Wunto73/FaTlDD8Gm228hBk0BsTXWKMkS4K0y9dIb4Q/6Xa3KzEUQ2HLoc
vT2aMtqXYk0WKAZzzhVu++4L6QBwcgemi6NsrByEFpwzFC0/WSK2MIjh2aZGiAdL
NpBVgMzV8W6cK1Ur7vkVLyy965hiD9Y53Ge437wu58j7PF0RS4C3b+jlscl7Kn72
I/iW2iytIgQOxLA9T6ud/frc1Pg5FSIG1LiEgPGGg1s6zAJyDWi9KpIzUBDvO6Yw
U5j6MKToi4ZOaULu2BU0Q69jRcBxmRuOH2U5gSZenJf2RJMCG1dD/AQz1Odv9zX3
ShVhiR9xuzMqhN6zTwsoIR7/58+pQuz2eUJ4FIbYpNn67k+pDXdJLRN6q5pthNHO
Xr2nazqQvw5/4zEluCFV4wgr0tJHM64r3sqhwgVCmPzRHNK3j24f18pRaBhHUZyU
h1mthMNp5e5HoRpDCyUuhWHmUGmeRrLSYhEehHbOedXr5wx9p5Uzw+yYqduyZsVy
AGK4VQRGGjE2ilGuAa+MiDE8524y8OmcMUfks89Yx/kh+gjgpbxGYmgqnoGF3uvL
X6kce7J1QtVz6D5+BrOxYK5BO64dAa/9vtr8RPSlEuGYnPiSK5TyMIFrXtLwI9sa
Wgb6OAw6M/CVIYhrRNM/+sKg0JQ9Vyp77zdczsRSZrj1N7ZlW1yPFW5Y0xGfdpAk
gaLF/IcPfIG+ST6wXPpuBsbCUdVdHErkysWMykbzqOoIW49ozjNhpwrxSKDOlgxW
sHlaRmEMklcU1qVyXxJb87Rqhu5jFBtQaB38pdCDs+OC0+vDPfcukOd3NZaDdDni
C2++5ck43wvwQeBIFB59TcIX1/hC68i5kxj7ifgXr/sOjkbq6z3Xjwn5t9RRlMtm
xm1tMfCDVV+NgqUHqAZuw+Pl+0jujrgBEUoLIPCPjYHPNSP/G5n2C9M3ZBEalAfJ
/1LuS2Ys17xuzhLa7CevNWUK+/U8MGCHEr466ZXX8gzsImWVeVmvm4/Tg5+aKRhc
6/9LI38c0rj2CnoZ+gbABlfh6wHTwOFbx1/APOd1XbHbJXm2S7Vp0i1TIHVY2kxF
T8Cf1zgg5NfdBSPovUVLxwQLYUhWJy5xonf3WQf+uS7CiiS3XpUot8WcvSDAhgT1
WdFO0CvRmMv7Rp2RcZ3Jr6wuL2vyBxeTVVb+N1a3uKVjH6egh1HNYt0sKtWHAvEs
mpu/B796EUDRtjhZ/8vQXXhFrejy/JU7GJlwLCSMsDHXINIyUexAiY2HGEo0MzOJ
eCpkNUcI+e+YKWP86tY9Ylt/GO0bVHG0YQzjDVdIQ+TAstmqyisouwTzC+t/KOUF
nDa5w868uqDwjJP47owyO49NB8OIWcz91l3IgCHTkUXNYi0X+RDvVeC3xVn6SXiY
XwPN50ORZ7Tebhpjk6LsBF7o2EtYdAPh2lXQJY44OHmR2VqAGirmniplN/haX//A
4kaZDaUFK7xFTyNitN3/pwUnw5i/bQgn+kS1hjZow+5oHuYbUetpQHLweUoGDCOy
3VMflExHoIX6TV/mHLiNQyvTPMRr6PoHftdVPNQk29ZBsLb4kOPnrYqfNTZxzFA3
kN3iYrW0muLOQ9pdnr8TdKUcCsyVWQAbvTtm3wPlCInLOfRA6N+NTIp8OK01li81
WuHqlkOQiChHIae+IfGHTi3uK+Fqd8fbApjSNsjuVFfxy2LQJjMjEmFpb95KR5V5
tufiK2H15bqYIWJRBj3/Dn36qsCxz29z7LG4KyUGpT0thoKEsQHA8lXRZAsBwTFz
ajwrU17+sPNfUNlRNtzCBQDAp9szsUld2XgC9U5P2juvnWIl8qT+9G3R2r+cRTGj
2XV+HK5ONkHPjKGH5Opk9OV4DLQGpsZDcv76DYXCl2GTul9Ef8jUTSOxswGeqogV
IYZRJNH4ZbTPd0i31d4wgTb3XdKDZok5iNCAIfDU1zLMZywR9AEu9na07p2rv2pP
BmaudkYzQQYED2+FKrQFsFwlqHviKABhF8RxBe2fsacvas20u4YrRPit+9PnPEHT
I4geHT1Z8sgX99P6iYQ0uLAXcRML1/4pdQiRz04ctUSisS9jZAjTjG5S1qZeSx1g
ogVbx5Wu7hG53t8ynItPH9NpeaQIuTEtqOqzWSDm86BDRugWI/TpftRWe25Tv6vW
U1LxljuRTqnwT9EypKDc1wZ8k2pM0qFsK9ytlb6bzWRNGigUeY6a3JhCKVd8uWwv
xy36QlNffQfTRQeQ+U03BL/5FXQE5hNBMODUiZeg0JE3TAYDV0YMxNRt6sgtZp4L
qLwzq+yERfYS3pQ7k38e78omjB+OZPW4DMZOGCpeg1lSiNnGLcCe6CfCxyjRFw6a
LVZxf1KIdzR32U468DcN+eNFEjtFg5AeirEDoAC6RZQUWUCnuTdLDe9rsEsMpzD/
oqT3/5yu9PaOzuDdAWUk5SRnbztONcXSHLKZHhR16jTc8IqlB8kcFwzct6K55IGg
bsG1KlDQMi3TMhBmxwyffLG3um78gJ3GxRSk0e0y7M7BCbkgDfjmvso4WYHzYz/K
YdtAtXnuIqQBAAM0bgH/uVA86qHkZPV7GIr6tiRLQfjFBMl8m36TMfq664EKYHTB
pbjEdmUaESkOZuAjOLSUcs0U7/yAq6CGRIq/pJGOB/JauHXFOKUWhOAu/PKIOCiJ
+soOGb9VQZbieNsDkMxPnrkc9VGsY9hFphCnJnRMvOalC4nmh4ErQM1ZZxD6xFf4
8OPnjuU9JvLJPqk03rPqV65hijB/HC0dnMw+xLThCAQRNMhSD11ElWZq60VMXwed
/yc38Tx25uZ6hLhi6QEoAswWRM9zUdSm9+uU+c379SmSjUVRCpO2E657k+XMOYlm
LRPp7JOBvQ8R8h1SJ5LUYJjx5f2cVFQyEGqdJEOq9OWX09aXYgOalGK8NhTv6QPR
3VrnRGtkcNOu+oGszhiixfQpgCS38tj6ga49YhkJbqXlgMH1NhDR7caPUyVaXhsn
TkE1f+m94TrPY2xqpL507BOmHzB/YZeIRhH9opH1KDIWwBcmvfavf+ZKJoDXy0PS
ai+zI8tGCVdQlvoeKnpLqlY/RT++tPEdLPQFjq2UHlbOSzxEYoRoR5hxf+mrktQn
h33jQ7xJwOjMNUqx7uoAXiDrQ3sT2or2qtF251Eujgz8H6/MDgMSNe914SVzI7vS
PXZbCzQ5VOLy6X7af41n05hX3sTt1/riImTKYCGS6vosiMZS8PUdoZobYzswXBX/
k6oWav8fuV04dbdwXZ9ReBwYXLjk67fCpZ4sO/xwRIUmBq27JEdlF9d26u62WDAK
ixGyqkxLQopdIuJqFGSAdpnYQEEY0ywEMypxhUmHMDh+52VAa/vsgz91fZn360CK
eQ/yhlknAzRQ0IMoxe+airjCT1oKxLAEqlFrZvShNqeF/nsTHxM4KY5xR5illPHI
rSBTzeL0AeQAnUvSlLFocpUGTpjiZkJrQorFwwId2mT4F0z8qxHEkUzMt+v+2cWA
MlBFkhbxIkMUah7z1huhoBs84OjYlRlPdZdrlQbWtpkS9wPB02Yf1L94Ksnx1UtA
mmL19xqHhOi2CP5YMjopqjfsd7sJPq9VVcueoP7DA1Qp6t2v1S9SFDKXaSzMhhXQ
ZoKpagwhazWxidsdb/REVGnY8txTLlzyPjjxRD8mnrLzmkxbfFSgmuImGILBSiYX
PLhYk3fxi/mHeJDgPhhtigNcQKLMtlUzjeC2Owt4BICBS/Ed/zXfgPXDxGmB9Z1u
z9dT9HpQ55OAXZgCCaGlz/cpUYfd3G6kkcI+izsdnFTybdBiPuaqL1tsUMaQSNab
HpwKcPSc7LjfscH/vsql5O5UTcKFww5t97F+WGTOFCORStR+dki/1UHpWxRgD7C6
hGDiRydSL1kZtiRdgKAFVKMNx1x3xxyWlp8LpmujF8a7ZByG4NuXsEKAx6cQC/+C
I3om+dPOLWHsvFZEiLYkOQbbC9V6xbHEzVApB98g4OaGiRqubJ8XdmliJgqx4lGq
nKD5Al72NT5PFp5803tda7tI0uzK1ooFBnSkcSUbtSuLXz7OIcuwvZMxPEyy0nPS
MHofCC2I39c97Z9j3uRgbhYqchGp/jPhOWC8d5Idw+KPPOddJ0HRFBuBfHFkLbjD
3SnA0fKPWJMUI5aGwspdtNDQBj6o9d18Wdzolq9ija3AbVd+N5Zu/BfIpPi3AVs+
v7INcROMebkaQpWnARh93n1uXhV/oDVvOSK3KtdmUtYLw1+0XbneawGfQsurvUtL
+IjOJsTUq/Yb6shM0g1Z1jruMJeWUHp3R28EL1Ymzv6H7iYMBXbrGsCl9/cxNfcO
isiha16AkvY4MNMwZAXlsgsluDWbqZuLUiweE1SNkdUudaXJq/t8GztIs+O9AGjh
ESNVxPFNdG5zvhburkqJ3TCXOucnst4sGAKzmNgPpAucdpYRlvCVoDQEP52xePs0
XbbakOxtVvLH73LnDqM9QkM3fTrgO2CutbCMcuzhPEtwwzVproPEIXcup4IxpPiO
m+TL2xG48VUYo0jhKalsCrdf7L9+LZOgusqknqrs394i2eZNpTX/tPvp1pbAb2Uq
1TrbE6D46boYubrgn64bFr10rmgs9KfkEfpIRp/z4M/QzTezbsMrEVelZr7nfp0S
34gcsS+xsCqiV8G1PTShiUiDyJTqFsEba7aBy0BE1epSB8fgnH7xYCxdG5KP6vcY
Ri9SLU5u5B6sxkEsHqUFM2Z3W7c6MHRqLGX7KCrNi4XhKyxapZhfxL5usdi+0a5v
reKjFWZQQe0fSIDLvaRGDE8ixW1HKAxKF3Vlh0FLMDmG+x5KBY0PsMLQh4ix6xpl
F+cMDPpMTDoNx+qwtvYpjJcI5ZzvZ5/x20sW7IcM7NCf1vHrcyh3I8M7a5Q+5kqb
1i1K777H/fQRq7i8/UMnGNmXxOiz+2soRqtDr5ibtv6bkM7ycfoMRJT4gizMWN39
MDu5jZ3rA5YAol77GCLRzTjLUf4rI4pyzafIjY/LiKl2y1LHAa2Q1VXZcZvnZ+PU
HgvSTZtqd+9LewSNWz+kgL3mRwsQN68exT++7TvDYzzrxKhooiO//w6sVf5bFTLV
VEYr0m0+z9qHEWhVqII9UHkWjqJrO4M6p3hNkV2/Bd01CU3X3AcawE5Q47EgTVMg
TuuRB/kLkfmksG6iqA7DIVpt4IVyAt97OzwwT366k6saTKOEe42nxMoZU2H0qbkJ
xWRakfIdH8u1gXgTZ94iGKQ2Uk91UJw8q3C7E2cVBR/8n2LxsZEBW4PvkN17VUz/
L4cD39jhAcktKQuY++6LxlOxj93ihuUbMJh2DXIyETfgruBSQnOE1ErBHKoH2y8P
cmHbiXwgJWCkqZ1M6owi/S4BNhpt4r0crjmQ55wV/Ne+8g6SBiAB3wNaDHmjTKaK
PEpQtpT4RTI/mVCtDhaYpZNyS45EJTzpUGLmNwvqBORjeJUSOpoUkK+Rp7SKUBuC
79fU3NmGaOSzvUH8YgbUAWhdNROTNBiQ+KuPdPYubkPIdwv660DlGkK0lzuyLKzL
UNvEhV2zECyH4+oDyNchZi+/0sSwKXdwqK/nz/tt0eE3+94eEDfnsYwWMRWuSglH
UwStxQeBc4eSkL+B9KVCvlk8JqRD05ERociFkHqrT5Cedz5jAotrHlNvzVi+68+m
ANlEVrOUJnQWo8xKzuNlAc/MrW7avVtmYDqSXyZ0Yk4oYoZELBJBoYanMbBUjXTs
NTYTkM9v/X5Opqba1p9EZ+WuVga9BI30Skc/cCa345VKfMsiEfV3Jwl5rd5jbRLe
W9uFK0zgcDFfHotsgz7+H6utHK/W22hUBq8vu/WEElEU9UKngto+xeMsgDBTNbT4
38lrSc/9dnf6glY4M+dB7wQOdTnJrq8QlzhtBhcjqTuDdWK+W5q6IUC0fAPJySV3
xTyr8auMsldHJWoq+zh0G+rOm1ce5mowGiNiC7XgKxsNPErNulebnGJhlhJKc2m7
O87rF35G0VSMaYKPq3dhy6fbZqCqF6OYYbwPRvLIQCiJ9DQ6BwO2DrwzrXs4qnTI
nI0igusRX2IiIGyN9jO97/i4M+yWY5UO0234IcUM9l/rwGmlPrscPtNA6pE6W7FW
E6Gy4H4ukvfQHN9ws73AnRVPO/lK07aD0aUvzoVmsI/JsVVv2oYlOr7Nd2Bx/9M9
amiG/ZX6UMJ1SF6CaOB+gVXQJqmcKiDGCUuj7NXX0nOIx7CV0w9CTDxUiTL6ZyG+
bMUEl3DnZ7N4Kscc7/yJNnoOvEAimhU6FL4Qlp/ptkOPCytg77Bk++eLNcnEsJaK
bngYqlvonO4K1J790Suuq2YKjGPvshV6aBtWJ6cB+5ZchxQxUzyH4EnTJ5uG9Umg
Pmu2AmCyECmua2OXhkQPLPiKkQlvuWtNYVycC3NPtitA5s+F9BPMVRrfm1RlLn0g
Ofh0fv6DXD+efI1ERh3fyJ06rt9AbjVBbCFiR+3fQ3Mm44Ca702i2fQ91XX7ONA8
ZdvCicJfyuEeqKl7lsSBDjR/fvR2fveuVMiAACfgyj+kXVBTCFrDP2uB4ROC9bQC
t3jG2cO4MgDQ5PQ6zC5y1eHHj2PAi+v/XjY+LW67Y+pNNOeRYdCRQNsudhC5097W
v6xfPSx6amhZH/EkOHXmtMc8bP89fTeqtJMF6vtZdZOFmyjtL6WFJ3201BJdQD3h
P/Eyreyv+W1DC6F+6DuJ3l4bXPHvPSG7lm9MPE4uAduJ2QHWbODQ0d5yuOQJMLlJ
OtL4IE6d6cqgK33HyNEEMiRac2MX2zCG7Xf4GvKHf+9K3FeKGfuN5hfNnl6xbQ7q
THZgX3eg9tQseJQONB0l9Y7awGNVrCL48qqTquFhpXyKR89xuQz0MHfoqQ5zfAaz
j6fhWeYQdwRDT2fUULv14s+MS4EGyAgs3C7yTtNdTQ55Vvctr8dt3qt3T/Aidwox
iiK6PcdV5vF4hUuXzwhUtxqlRQUxvtrFY9arVbNQn0TZEYxm5ZD3npg/qTIW6sxw
EtpHdbuq0s3tlk1QUTB8xzJLEZhnl2ZCkK8rhmeHqmcFxNFhZzxKts2btQzWEMhN
KGRWyAxDq/qq4jAQZgbPgln16g4l/g7nRLYbOVenHfdKZEXuM0WEj/WtFok5A8XW
0ymSaNNt/5HXuu4w3ArvQtXNZYJLAV2ndCTqeanO/2727X3nUmxH1sBPRfiRbNPo
2dNseHMIiCQtH9GbiFf2w0Wd8o9lRnLMltm50JFYusc7K5jSZhSrFnAMYFg7S5Mm
i8c+d1SnQMN8ufDm0KDZTXJEahZI/Dj7YIsj7IuifV/okVhRTIUpG/KdUkqzC2Do
LfEOmEntUTYcTPQiprRe1/yMaiIe+UDF75DuVT+Mgzv8kxjYmqbqxLU4YrdgTbm+
wLI+cELGjDHri6S9sJ5xOQCz8Q7FjH1R8fJIAXXGCZTcVssguNyW1YGQ1veihkxr
yA+xg0fAlUKYE82Q7k8FXXtNJ9lgbeIoijHHRy4/RNBnSiS4W0EuOKFjx+5kK8Gx
Ku00drMTdk/cizymp+kDUHwbIujw8hp6qmGNdrbUSf8hGbvlb/J7pO5AVNNhEkM2
B+ZSYEZXlUaIQZeb4tCwt7rAazmOJvX+VRiRaUqSYnLPUn3Hb8URhe4+t0wW5CHR
gKUQlE38XbTAzAdMzO2KD5TAnC+eOuuzPGKa+GW7icFCYfX7tVXcMsPEYOX/ENh6
Fs1l6WXZ/uKDK/JPBc8aTTI0Ea3jri/9DxA4PgxH66Lk01gpJUPdsywpeoFKTw3B
ko1evXOJXkc4nbcyTy07luRv+DSMfZ5M8KqDExPDqyeDDrqf5yYCrMezkbGYnV/u
4KmX/Na8kfLWsMyOaKfM51KlhKDTEKbWGmmzhtZTqyOXpuEFoogkV9R1ot/9jj6P
lpF4ur48GgwJiPl3p/stbTjOJPZeMyci5cgnXxQFx2xHrcuhraHOTtQMVJiH3V+9
aGwgLM0heS7Tx7JcwfK5R7umFrM+KTSnEUY95rVm5ybC/CgNUNNLIxVK6u0GYVdk
Igm2yBIfx5irZEXdun6k+nZKLat4zObuyvp8ksA5BpZlA49OvmPAacGuZZ02uQKn
hkwGvuVjUR9GtKBO7Ro39G4s83aYFjf8xaDrqIqtYVAxyQDqfYTOFEMwa+Bk9XIn
e18T0KbM7HF8OUHAR8uQoGyZDo8wOBVl1LVsi/vxgHF9wu6A4IzgDYRQR5dcVN7G
D+siEYjy4ImBm8AXN3Imp4USSLZZ0Czg9nJtEqQviFqcMsrkmZgtPniikYFmGZVH
VBZMXg8DM0yQF6a/oJckDc+aEIQW6UVQV6rxQnrxTt4CBLXKZRIul2ymxFm2+fj6
qhEb7GFr5Rpp5SioZJeNpWqmBOZ6fNKEPPA7FQyBIgfaZ1KyUXWJBjpiNAL8ODlA
T++c9X32X1pnGVnQjVcJ1PtE/pkcwvkLd0LOquowXFXF4SpyM14d93TcYn5BhvCF
RiIp1nX6BgpNUN/KRhGGElXAt3NoJvkGCcgsjrCqPfBkowROiN3i9SeTb2nCMVsH
b9PKUigYRj/nH2Xcz2hw2IC7uPg8P6r8S4fNvILlslQPRzucGY5TwONn5V/z3vmR
s6CpP0axJvKWIeboiPe5wVabwQL2AsXCIB896HVpQIU5ZMNpkfFMn0FdVdW5cYx2
PjOz+xCvxkxQ6XWLIro2f75v13z1cOHIMvbheS9TOD3r0TKCJNuLat5RWtYS2k+Z
iqpYt2i72bDu890fGmGgmawO8HFOiASAA/tS8lgnmkO9OAZ5Ome41w7TCfQwy4oJ
hHmz5APHhCfMNV+bZM37VD37glZHbrPJsWYn3Y6t9+ymoHWvGW/2nSbv5lbOqje/
cOtXEfkQnNkNMI8TJOUfhpK8VCGYaQa1aJiG7GmF0enOeuR8oFWyYakHrO9YpGA9
cogZq5IRJkXLXhvOH70xbtYsy32oGoBDiNgq7Y9yEheC/7SKIFL94sokvfgZtRD7
0a3/5tHt0KTPOoObg3Q8diYkHjpZIPTJml+58E5u5mmvdwvVtoz4Egd8GCBbUnr4
cCSvlOf1q9MRbD0ho5N2iuD0gNqm4I8hmwBgUgEIX9/eZatsC0DHbyjhNAEQuGh7
1ujkxlT/ZB6K4LaTfzEVPTVDrpD7ZAtPwuYruPs6sRmqJAr4awA6QCTtwkOMwKPX
0BOrJfOexpeKm0RkaF3FK0oJJ+Q3BNZ12fPr9f8mZPMEWarWoUIexCDgt7GJ1SYA
qFPaEu6Dne95EwM74U3pXYLfsXxiO73d42D7kCg6yVZKBucMhO9cFLfh8m0xMTvq
IRi1hsBaqTU48xG8ix8mMw1xBXPlSL6ZoWWsHEfBZt/Wm6HPf/Ii2B/gYGFm9zL4
njQSetwN+OR3M+I6ojJRU0jWCUz542jkER8F/2Z5lmrX5sdLmx7+Y93hX0OGxHJT
jKhunxjjhBxeXuuhiHZmmUe1MAgAumW+DqgcQ+q5CyIWda4NOwpy/d0NsloiU+qz
NakA+uNrk8ZFVlezy801x+gK5CZ/dQN73GeB24mVkbILrjC0fMgp592NyqWWohih
F1Om1jCvy8nlmu5XGux3R7yQ7neVsekj5XkaMlsZJppe/jEVndVo0MP2UazWBKHO
zMSPslwjWwkPjKp9Vw5+to05j290Q6UjRswZcaa+CNp97t4xpkBBJ6TbEnoG3mi+
SVXPzxxJphdai0Rx26zZANy9QsPO7Vx/A6VeElHEuZcWbYP/k9gu9itY5l67o94M
aVUOMndZclfkM+MieztNsAfj8yp5lnF8iFyLd6hc5OUiDflFVcxlKx4GKyoEgJ7M
HXQ/3Z1Ns4qv6MaBNr7keE+3HRcdyWnTSrrFxP1UWo6+UcQujTEhiy4aBwvDMBYt
+p/5fXjogurwr6rzp1vqyZTWhGMsCt+ZEcwzDLHEH+LaIVefA/wmlYQjtntewavD
xZTZa56loH0yPY9PbwEcci9D+jzzWK5tgNIn1HC6bZcg6nIFWsDrOzjw4Gx5Fsci
CUW85OOcMHGPU6samGwX42KMEmaY/DhIKaqo408802L9qdFtRdcFRoZZ1p45zWzA
44/96pz1LVu823doAYjXLAwKJdAqcFnu+MCGsyQyedvBuXzfhZaqDGiViZkfA65j
6c/S6E9K+ccq88NaT6xp9xr6LyEX02aDSfuVkKQDP8xJeWl1sOCqZmB3gqeqa+x0
vUBUyyDhriHZvo6YWnJ345/E73brxar5vqdyjTMWUSGRyZf6GUQ/I3CbNHe5YkrV
QjsQVvfrHBorU/8zguhAkd7tqPWNmulAD98fuLPoFc4PbIHszwoS0UZANFc+3pAK
XR44WM3OBC32eJ30yqyNM9ERZGyI21sL9r8tdEu0p6I+fnJLqoseOzKu98juCJ15
810Wsf8Lxrw9W3UHXw5UcNCLVU8u4j32wrVDiF/cHdQvxr4+mz7zLD2gPRzh61nL
pcgSgyKnXiTqeKeB5tPgSLssH+Mzs5r09MI4fGKrlt+5y2JcElDTAFHNpkCWTXaq
bgceq5Qvwx1sNxRzjxeWdAEtu2B8/Rt1T51sDzXh5qU/gNnOTo1S8U5KGL/bq18F
J+Yh0G+4rDNDPRx856Z2mutpmOphD2NyY2oigcQTSBoyL7DuQdNK4C8+MTr6bkEp
WYeRkp9/xx2Z9gUDs+h0Mf5kw6ccXrxgZA+mDwbo84yiCRtOntUdcLzdrxk5yUDq
S5oe/mlOe84qxxW9tquG2nqzV/N1Cf6dkQ9myX1ZWOI5NJZsMQc5+fqIQU0JxtiY
5DB220GqzXrjy5RKw+uh2zCjghPtrs0DLUQ+SVYuUhOHtXFHNrvxJDVMxxgLA2ot
1o/ZZT1MvQZIW/bmKlsoBycm0KSK6nrIrjsNShHOOoW76RjX4VNkScIUSW/jTaOG
XqmkDv/ne6yQ1hB/bOUi5oz77fXwKcR9cZz9KNiIBpBVTV/IyiAjbHo1cWhoCUxI
QGSWCdRSsCodK1nfD3Q0fLc8quxQUoKA2ADwduNwolpxcA4bZvizlpCoV/Nw+8K2
5UozR5WcOhafFK1wBx4ftXpzLKbTTBYej7Azl3iyg9qPFp946fdoOsR1AINqP15Q
l1yhv4VqzE7aSxm+OyaEl++kavq2ut1OP0vb5Ty5rHZHAAUW2b9IL/2lQDxkmKiN
YQNx8DHaHLGg0JWlyGmFB1VmCU+RqnHBDR3TmeYRS3IO8L8gL2zqOXD0Sgm+saoo
240+U42RThxmlzU+/9G76ANsDL9Dqgutkb/EVZoQkoqorPLiIO33GUafnIZ3qRCF
Q08oUGUm33fDedJN0rWc2n4OFImYTFkFfr86cmGHvbUKio4NmKeUYgfOtpYA+3Yx
BiQ9iReg8LyF5blaS3cojMaHuk+taI2b1KohvhXb401sTGkIH7OV5yIWZDPbhFzB
5tMeVEZJ6kfrttuVECHh2+uNGH5U4J1e3MtZtxBj/cTL5n6q1cTQy9R9pDA4G/yf
b3nk65YU6dOonnQjZBiDiZzY4RWE2wDxyrn/2W1p+ZoNdM/It7OPcTB3oDqO9mhP
AMBK6ODdyuLk++ZIkjzIFQ0hK2WKwhhS3FZddgbLSUNFCfQDfHFFU0B3S4jvcI7q
3NdvVbdRipcFDWWam3/ctXoNH4Qr/IDhgKUlUuPxY9u55r8je/LeUAt1RUVDlIMP
vXIFIFO4CqQH/+JpJSQMNDxQ29H2mPHJY9eEtayBmxemQl6iUFFUWrhst9JxgMIz
5UWe4uWD0HXhR+VFca2M2RDOw0hOCk1ejMEfFagxjcgYoAz5PjUZlzCWmubjhF9b
A7RHkVhlBAEulX69BwrBgYlWEbAX3lAE6QKpm8b2MpogzLMaiYGs0+fbpSYGSF56
+/nt176z93OnzqFYmX5zoJrMqlqUGq9UOQr40ALQMEUsD6DWAGkJ0rvUb8B1Mldl
tn7rvcDh9WaZcFkPsoenMv7Q3w01LXJWBOq/cQZgo0CYoO8J52Qg9uMgKQgmsPPW
uW73v6W/n6wElH0N+QRaVKs0boObTECrFhTtCk4U3pUDPocE6vx43NnV+7ytfi2N
p5pSErWGJLVOfqDDzGEpujQtqyA1Fgg+xnEO5czZw8+ZJ5/KyvP46uJCr3FkV6IC
0bf9sCFaycCUJ/oQZ5rd0NdS9pdGwAmpLhZ5HddI+W5akN2pltvsmvD6tF3dPx15
bUbT40dTwZQZXzx+JTHxbm3BytmtPvCyAy9jgiV3/+OX2+KZyZaBm5em3n4a9VnR
SXNzdeSbiBbH75hhYikWzBF5H7+sZycWJBqFV1KsH5X0+Asoqke7c3XlXu72I8UC
8w1Nc6POVkOcOMxaWtKcwpDQRtPiCDYnwqZrZQg7pyqmy5MQ6rX0eMifI2+GyB6e
PVv+yUOcN5is3D46QG7uxtRM6F3Oqo1i0Ywchor0XDX9BTuTLL1VhQfc/T4XEwiJ
mtEyRAezS70+DFzRSBlBumM8WhFmw0odL9hGuuWumMeeBt1/7Wd3uYigFl1Zh5m1
/8jZWdG6IAgYVFYUTlnIv2l5OJLQ9vqsjPZjoqaFIzPOm5O9tvtir8o98u9jga6Q
ZxcNhiTnQ+kzd9jFctWLl8nx7sAGf7e5zRjeH7fTONaBNivU3sb6x2o43bBACcA+
VN64nq/S0CMj+IVU68+vJuq8I3MnsvavLdbmaL4HrmK+N1hPBPVGxSCkNxm2Aqwr
CwmlM7fNxsPhjrFM5EONmoa4XhxSCA/7r/DxEIEXaVIPgqnjag//6GEVGU5PCfQH
XFKe+ThBPbAb2QoHuwIK6vjhtILnD5Wp24Lb9OCcDMMGEC3TLed5XG3YiTtz2IrY
BZITMftc1z3lnltTuMu75kBEDn0B9L4sjPbzILZ1RoI1zgfFgIlki2E3eJDO/ech
NRjgdfKnU1Su/yIc/BOXNZlksdtpeTOI22P7JfhcPVCevn1pBYcr/FIe28XNFfXI
rWIqweAx7kQoPmf47Xp5ONtGZxJFNZzvgU3ygCM7GSBcItXESLJzq0TIgomOed8t
VV2KdFIKKIx+VhSSRtCGxuVJJBN7qEeBwzc46nnr4okxMwK7VUxnLfLK0CrUj5gj
MfgugTKId58AknYVu+CQSu0UbvTGt+eVZmx401+DRXLnIgV51QPBtHZ/DlIhi7FN
+8lDOVEcuTDosmWlOfit6ttLo4fo+dbw/OOBGJU0qsAU0StIH6OPmvvHhkuXaly7
BaYCdleD3D7SloyiFB/wDhsH7bKU88TLIw1+4MoTmUoNK2QoZK4qTnc32sw3WxA+
eAyS+oYakkJKjuegVc95b+CmSZioS85ahsGJAxCeaQVYOOs40rl5r2M7oJaGQoMm
PT8D3Oo+bcfs6UcPhYz5t6lTF3ddcVfNNU3XFrpenI3DuqmcsoWLphMbWPa6O/mk
2PQUhNWCoCtyDslbyLJRZtSMDO9OLuLasGeE7itpnQeDgRKunnHt34Dge0bWvc3f
LaXHfnCYr1Vy2plruWWSumuFy5EIEHY6jQF83ksQCuQfL2eo4oeV9v3hQQaQ+BmK
/LLLCqs8CHscGNIz1yvjgjUpj4oCMZJTHXXhvBMrnN3EEesRwhjPjsEGtPcJGvXp
U3IYrmH8leKI1Ddpbo64XjV1kI+BL6U2BLtysfrP4fnr+EvYGpi5CKR5aTCj8ey9
WpYLb06Xs5uWsFOmAORx14IwiZehcMvAZiEuRtBzwdYLMHPtf9cCm70o0zrWjDmx
KoUUyz2WLK88vUx14Dx9mFFnbfwhimvXjRm2ex0VQx5VP1cjp/vdZLtEcys5qNNp
Pfs0M+IR/IbzrGzdXhXT1VHd0A5flPERu3dBnrlBoe7jIZZfHeZSQVTAh99Sbb6O
YQATYWjwasUG/pyRs3hGyNGFRTKOGeQi5FSjmgaVcsBhnuy891AM3xXfO/VQjtyT
NGvZGtnCNgoHyKQsJCuEZj22QrOF2/LhI9M+bTCtDQRgrx5w3NUlvd0qvErG0UdK
wrqYYz/05YpjUOnVo49H7IvXE9GFfkU94odEfAR737lTjrtKLrrodoOQAkk4X7Nf
czNvCL21dZZ5BCrk7KsXlH86S7x8zuKDuRB98c9O2qQID1oWMeIh/oSZ+4+VaX9H
0A/6pqI1Hw0KcL5YvsibqwlpzKhMm39KDg4G7LucL/h0nWihxKoRURk94Emng8UE
9bQeoupLcWBp4aNEn4ZcPFiSFnKscWlufl5QAHUBJRGUqM6d3lop2DMDMWmgeyd8
oqeQ7BQeGWCNpWwo5NLOVp/uDm6IFG3Uz+6WxA9fWmGvY3T+fdBlF7yaG/QYOwrH
c0tAcUISi5O9xxYTgpNvVGRt5AA6o5A+GtkLBPb7jXpm8rvb8QwiWTTxX5F6Ghk+
+qFgPm1lCvOVB8Wh6z8ijRw7fFadydOaOevNR98HiBsuriKnTlyyXnG+FVXaiXYR
F07CxJzMDdFD1WVLNSvAoRn55/nm0pckHiS4tQbSpGJS1SDluooWKrSp3DM+49I5
GhiyoOlywylxa9esXTEKyJO9jn5A+o5OOYFsWGlMXQXqa3gC/CR4ikKpVdhmykTG
L5WknhDaq7ysZQHOj/TvpkMiXP0E8WPiV+n9JLO2o7XZpQl+TyShyWL/Gk5q1Hdu
uuu7HnF1MXKNwPk9Glk6qXocr5CkF6o2MgVt+1Ua6nP19BeJsAilV1oe4d2SPZbz
VmX2rnFc9g9LfUktvpiE6sbjOI9cqGRVpkymSE45irMQGl7i/0wC+TQJ6HZFeTEb
NTAIZuVcVUs1ER15HiEw6fPumqZ4mpf68YF5o7lUOf556HDww9F6YexQRYeiQdpW
5lkFRBDzdkXGKjZDVescUwvHCD9TPdgoY4r8us01vmEke8Zic9R/3TlpujRzbDvT
y6siutVAo/Uw4ALcSJ9T9+f6q5RgH524obZR38IT291rThdzRs609BDdwizakHMi
J1A1bDMNCmcrc272nsoXYg0yHptrcfFYWfLZN7qUmYkEJHqOuzSA5N0xHHW3ZJ0n
1aF3SpOu0Qo1DuAqRRalzl8OlRDzNg2r5VVR6AY5vYv4rE5Zd0GFITrDbKstM4S9
f/jQJY5a89VGc/nUZRoc7bjvY9oQKbuoxFXsEmr7wBDyzyqIK9ymIwxJoYf9eJ59
D92eBG9PHOnfZpbea/rj1Q9VXKho7xAO5qOxrSZ1Eg1IDwAJjItRy/cVXwomQ/nP
DPs9MdxJKl+CarvDAiyxOBf8ndBkwmrFMaNdW3g2Oc/qNoaWatSRdjpSsPqo4boj
eUE2g9vTwqmBiPVniBDGrnJE4svdfY6KlUT1qNoS9FpxC3ey2JRWTkNtou3Mpu5O
59dQPi2DYnHrU9LI9sHz1A6ZR9WMqNpfIRhCxzAl4vKy4TAbr9aCkRlFywl5RnHQ
zupn3a+XuRkiatYRatbmgtknUXRgmgjdiSBudby736FobOAfFaaE1hLbzKW7KGdb
DbiHpNonrlD/tW3Fy42sARUDM81x0kmRCZe2U3J9a6e/T/aPacbEqc0Pg7W/YR06
W88z/Swm6lVpbLP6aGT5a1cZTx1cykEnjMvZmfqPBAn/SURJ2VogTOGu1rPK3T0v
KR/xdQw19JVVBFk0o8HxbwvyIrKXoVEHpdnBjOiLgS7+5iIuTxpubfRNnKLiwjtg
zqZ3c7m9sz43t52Ppkj/DQEaUyYsdi6NKM8fa6Ej6XDc26MBinLlpbLL3CqXmPy0
PJvZ72BevdfQVWQrk6X+w+v48ZKU3HEDZMUM2Uu8PLILor8tSgt7jpvqgcGnuL6M
N4u9o8OJC1rGWn/cUdTEJzbmlvU5SpK56bRHMe5NBqOPPUQjZFAScVv91hiJ37Ql
44rJQ3K+KvIY2Uub/COnuxJSaxPuCMgjLRyazlFv67Pft0Hu45ihTfQWfoxkoDFk
RKynhFpDAa+bKqkeX0u3+v3VgGQA7zdqpHAIUmlhI/m76lkpubAw6j0J+8dwQ9SZ
NHnEpP1e6udM6FJIKVrsDYLyGwBmdoZ8PJ5iTWyr4uVKq3l6aV3Ov9ejDg3hgcLj
p3FH7TRgHS+EdPJriph2U/ux7v0u8tjln4diN9jp9WVbDfQMKJAdy+5cP1atPjew
gu3LR98ANTbWmR9P71yHYLqj1REQGSmtH601wvmF3bL5kU0TjnuB8arwILrz+Lir
LnQ0hwMTkvc7nmcRQsh/YhgdoptLEyhy++PlxQq9U33B8Ku0DVwBBK6yOr+34e1E
2ZDIk4CNZ4H/YrQlqIlxjrg26DE2iMNwctF+2DuMyvgFCN79DdgZKxk2e3/wKFO1
2oZf+C3amaroyS5AdCENcHFFvfzrW5V5vecHV6dvXvv9xkbrD7HHt+yFNoMuxZ7Z
QGNcFZPhgVAs98IVqnxeDMe8MTHcsb34TLbR+fRosUnsPAKsZWIm6x65WzJzJF0q
r6RrhTf5cTSFi5zMlpg+oStwS2cEKFlipW7X/BAMlXKZUtqXTZfSWX62oh3KyYWy
+7Zd7w608cHcYU3m6Do4UzJ6c0OFDCepnn3QJ9beKBAGAbcMb4F4ENl/F5xx4WG/
mseWxkOBZm+C2NbZOSfRbaRUUDsjJQXNXwOQmV6Qb+ehM/Q455/9uMmCA4GsXenE
LvxoNkJN2cdxTYJ4lBmXZfYwJUqFkh3eWERjGJOQ6CWKm3ypnBHQ06YGV4uvIJM4
c50Mo3x2T3blrazVKsBTs5jbTZJ9XXXZgApPx59ItSiZHnSxhPDHE6cVivUhbtvG
d/OcXjs4WQzPmj+sxYz0RdVagVb8NteHsMcfjJztwZWVRocfB8fyKLbumrWeEosJ
zk6x26/4NzKvoC1+kkV+L4JuyLcuWhqmQufEvjZFXXaInH6mee0UuidSJDtwe3BN
k4+S0Y+pn+H5HJh3qeDj0lMVivayrRD203lMe1DSiQVbiBkgfumWHchUwUvxUBs8
VoYsSnsHnpJ38UxtkaCm8hNP9WneBTybbvJhtqgtzCiyfGB0OqfCUDpSMwmRGgtU
zALsK21wPURpXokNj3wZ77K24BRjMmYhvU7MwVeCv2v4frwHHoBaX49WZG4eMMtk
sKZDs/rT3ys2bn1KKqenJyAJsDRi5WQfFE7qjg5Pe+wmWpOVuacVyrvvH4up7bVW
pXfRS/yJuknZu5W1FgG9OhqxD1gfmFL8TK+/cnRhL4VZ2vUorSV+bGfljGIR1iyo
Me8/I9+BmuP2TyadbE6s5nzHcApiZfY0FAT6siMWHxqoA4lz1TaYpB/D9U/g3FMw
b+qZGG2GrIgce7GVAdbpdhvbYr9+6j3WSytqVPeEd/9zJvoNKH6gi+5YP7uOEJLr
dpgpiOjhFQLkPh/G1woVbjkZvb9VSZSuQv/jorKslXjRVJ5kxRtQ0Kns9P5F7QRD
sjc+cskQIbChBjELp0ER2Guq4DPE6Rg7EXSkCGavgTVw/Vq8C02NIdvoHKCJCMyG
cagQaJW4+qp4vQW9FxPjRaYTXuoMWghyXe6bibbRrBn03W0iUzokOdSPbVAb0+0V
ZCQe8dsT7aVnSusvGaElkvwEg18aYjUgXdceGNhyoV7CjI0l4QCkx+Pjzk31bX2R
Gyt/EOnTnEr/xTjVQU23Oiv9hW2YbyqWxwwr3l0wnO2Ota9dGLuzEjq8OVFy4NIa
OBEmnnkGG4jYiVlvGEmzLbwH77IYjYAxnN0MReZWNfkMHSL4/qnutPGaeL6y43ME
tSYPtagHyJKd1OWE6JZSTOBOzwZDy5BE1+IwcO3OQ2xPKa0k2eFzZh72JAKCo2NF
24Se5HuB11XdvQ1IT5UqNlN9/+JInnx6eUTKqCJQuu2VxAbA/0ph2rK0uQOhlHVa
iH8Hzkm5/TXOw1EQYK4jVl0N0ny7KNPIElv3/XrJylQZjw/Uj3m3ToBndjgm6Rop
ViWt2vOQE3H36o3MhSIzpxc7VqZNCzYxxijvIP/y3DpxTBMxBHQEq6YYaoePBMdH
998peNuiZgDB26rFbTn+RFbx49Mtu33CY2wZJkcS+vJJ5DfqRv4jvZbEubKaB3FB
KbFoFHX+DYQVxZZ14oYIEcX5YB8XPhv+1dRb2FBgr0F5nvhRP9RkRMa3yr7k5eQR
pNKrL2oJ3bLJLnpjHCvZxs3eI8rbHBU+kAJBcUWu5EsTeARtZvgYXWajSS3JQG/6
pG1h49Z60vX0Za+ofs4sLLnabiwZCC7tszgt+GpFYWFhGgeRy6A6XugVbrhLKaoH
NjEZOmerQ2NNFxmBzE9VIg3yB3eUJ0Z7Nru2O/mzEGWsitZodIiEqnnJ9/re/t+o
RkrXl7fR0eb/TCPGjndAKW4d+BZ0xG7UAHg6WYVajpe3TG9o4XQeyNzqOTQPxfMq
CI88mVV5eadZ1D3WHXxhbTGhWW0KFGf2el9FZmsb4ikf0YSpJsA3rO7GqWN8S1Bo
sO92sJmrS+MZtCBDcAxZM7MDrn7hPl6N9NtqIO31BYGATycd8O/qzSfHDF4tALDZ
mXZ2H7dVtkMTg7H7BQRqXpgPng2FiUp54zlvYNnLE8KgPo2aWleeYv6QgcCQPuCY
BGbQ+Aj1RKkkSuff19MIv2XpcBnDsk/XA0qPB8uu9O9ZlA12RdWMPA9Q5diaiR9D
DgFsZi9fu7HaCTcch69Ao1UY8M9v6C9YOEfe70M04zKGenNX5lgf1Y1bC8Eku4Pl
v8AETfjiVsL3mzplyXx6RLGIqMUSP48xJUfeWh4FORNP2qs839SYwfLdXU1fw/WB
hN45d/E94KL5/d2W7gjoUPQYtf84D6sHPKaTILDiqPi7ejP4gcf57afE6LRYaUuL
EVMiwWXLxJc/7l4bgC9blzEDseUt1lTrlEDCi5YCivsFESySN2La8dd9cmaJPkOZ
SaWANjd5gefG+u0IS3wxxjidW28Qg87r3aTyA4YvYtEaZ2R2Q02bSy9QB2W9lwfE
f7oX1W94GWuflMxEHK61gDq2O1bxOTHdDy1yzyFUqTcIh3Bp6arUXyfOhjLhluuN
/qMssHhWjk/kSy3xaQ0CNj/pXpD7RvT24ZVZ0l1WX01OY/idV/7mKtsQlhR/P+gF
aKb6o3O7ka3H1AU0IKESJwtkn/S1nP7bK/+Hjltb5rPZosstAg8JcyzkCpd3Iync
T+W5rx1ADPqFo8xS02qw25Eugbv4LOWXu9/0tQDk1fA6SqzPBdWuFNQbBFg7Y8so
8bCwt/nPy8X6uIMcHtl82E546THSeAk4q9FHP6Y0LNIcQYGEe02lOz7useL1gIkq
R6BxYdeplSKBwNzpuA/SOf7WTOacrmLBMCbMh4xvu2YljPXvfwT5Z1932hvX6W5s
bUOW1Z4rktJseuxj3quopSmIjpbGVjZAjrGTcpgsOgDP3iWcDk3d+IL3oxGiqT+z
4TY5iLZngm7QJojZbBJ8MykPlTzHUkZ99sijfb2BcvmUcz2vK9/G1EQmVn5FDIzp
X018QRMHVpIGjTzmI9y+ytE0Iag+nDzfcyOxXwBLOXbz1dc3bSnJFMUyK9zuofqk
yJFDFclllx88k4f/t7UxMo75p+9LVJePuW8xqJNHqq1KyzR3UL5u4uYE5wLwajO8
SHHEekEyAoW0+Kbz3RgYsUyigUfr4BRrbAbiqFaSMKLvfvTIBCO4ekh5pD3h+bcQ
EuH/uJfOUTACk4OmnlBKXz3lXE/xdZwyXiVbIuGGENcL/0pZnGJVgA+aewPlF4wN
Uzg7RlXl81/0nudw427RDYV36oz3nj/UWLoTBdcnFmGbSm8sgbxBoMLqlkS7HNJN
28Y+E3FBWemvI9NLHtNzqLTMS+K8lVzOf3GAfS8yxTwAvaVfzjIZmbmxwWG+1/5m
K9dr4NBFFXyixLCSX+6IO3BZY28T0hMho9OrUjqxzZmIO0hXqzIiKrFYICVmOrpD
pOsyVWjLjEI+Tn6dXny48ihPJWklKu6y696AOsYqcblIPj7fWhxnkjnZYeEQ6r8v
SDHqcEULGgTDMh7vj2oYgjaZywXUeNeAnnmhY3t9GL6uBAaTf4glD8qsoPBN0Ubx
8dV6DAWeeGXr5pYAxnjbNjaSDB7TzaXB6Bn26IeXU41FQEdZceaaQZro2tYD+3ei
a6UKH15ISkDUKVemHp6sF4rgUnyjTCoVzOfpE4BI/gYvdWUxlp29rytNakTT201k
qyOaW7OsU9qygGFjCMd9lbVl+qPG2g7USjb0i8+6JlSv5gksVjEg1A1cC7PR4+om
V/kFJd8zqSU8cU5Dyn1zeGkGW5evw4QOzJEv8bQlvQFfmBAbKwwZs8t1CJblu0By
wY3J7QPgwpmRhdKCbIxr9fpO+AWdxG6IuzwfdibxdUTkj7eBXo3sLSeuXs2n1UdI
7rhJYa1J4I30vm2UUS6QcJpvrgVbIbslwvkEqMGwd+5QrZ2KgE4EiIJMGtclFY1w
qr3HoN+oZpzWShZsS9o1t0O/IxynlrNqcEOljHx0acklJpdExUlmEezauuiId4i7
7Cw08laIVcHx/WKFIue7Qz4Cg82HdC+s/BiswF3nXWQOLtpha1TATG9xkli5pk/e
VZ+mDfdctl2pACd7NrbUYDuyR3Ee2rzU1CltG/LaTz2CBPD6pQP88btYcDbAY/qy
kfwDfonzsErtmjVWHRufmPj7TAoffOVU2lYpI6yDxIyMpYbMD1bUH19ZnotBezK8
/vzaVbJlvSW0eQx93R8AnhYtpje2ccXaFojEO3aBe/wxShPC1hUF+hQDJtwegDTV
FwDoTXySmhyunqZEn0/VpwlyUTwCMC1ymUuBLJW+QD3d7Rhk7Id4wxBEGxm6eB1r
4W4Z+ixm6O1LlHMHg5tp1+s332cu9biLnlhLpwvXDZ+1DXI5EiDjTLDF2gOYd1GL
taq6tfLgcFrQTntz663DAnBnUeT4i218Jyt9nON0AZU/wk/p5sLmUJ43lgcPT/8w
cfFecQW0r/D+V1/qNhvJOMQ6Czvs0IxFsgualVrOuMSM3KMpV6/jm99qnEGb8j0o
FqWP+XWSGu4OgvlUpOwQhrY0oHPDQkmozxaxkKe70QI7WgmaFpBjeHvnr/iY85WA
4neHp23HWeN8KeqS7J0fzGOEfr2B2lBHlytq3DBRTu4T2McXDAU3WB1iVZrVbUuQ
IZgoS3k2JGOD141qyk74Kl4pFR9RpptEew/5coDi2erJArVS01tek3tQWGFtbgmx
sfI+o79zxMbrFRfhI3EkuloUO4JUVQwcb49rXd62fL7GP2OggGETQ8u97psALvlf
6qOhfvGtgTkMez48VUbMs5jJTednGjZl+KPzNKsFYeTEdMmUAuqycrLrA/fCuIHn
hkz+0td1qAJ5p9P0Re1NrL5Wcq23AA0xnuYtibWV2vL9VlxaWcmn5EorgpZvZkzO
U7MnkB6izmHXJhFtYPp0REBA3zTduBtj7qsYgCT94Eg=
`protect END_PROTECTED
