`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uvIQQDJO1Q8/JCqOC33nCY1gYoHrc3yW/60Qk1189a1w0XQ8gVuder4voL8gpVe4
pLPQBeL2Rt8V2fkeJz5QXoTQAF/lxNCHyQ98kEAiSpK3PIq5rArUYXNuqp+ImdkY
bP6H9KIWhR4Raf9p+Ry5Uehd02yqLvk63wRU8iOydTwe9PrhCsu4TMqv/xkdXFeN
o2/L/WKoBtqe1XkZzqT8curxHEAy3v+72+a+SVNfGEHrW4XBTKvmaQ/gRxdKAlvv
om77RKTYW47aN1yOhT39mxXVS003/dqhgPy7gajfad2e5U+66e5gSPCag8Bp5tME
PdCaBEBqeK8lyd28FNZ2wCiJg0UBeez3jQb1LABCDdJro8xqbrw2nZjl4F4uKinH
S0048+dgByNRr6sf9ZBczzHv5gx0Fpmr5y2uHyhKGslFROO+SJYKML4WvxLcPj0u
EikIMAgYHg/V9JpI2UUIhseIreBgXqpaDH1VlnqTzhB9XUtU8V83ctocNFDNMQg4
V0sTErpTR/ZuV8KYmjY3kHMbr2HInsgqWcSAx+HGYllbVGRDeGWhDsX/Aj0c8VwT
4lQYptjeu1qnBn3BAvD1xsAPK/3lIa1ODr462ETR4TXw0v1SeRepPaMVumW5UskS
8MocE5i9lEB2AMkmdudQYWWhNtCSqo6yp1pSwcwWU88q22BynMbg+zTdmNf4UrCr
QMMEkaJe39DXZNzaAyU6qh4JbGP9aqPO4825VKDL2Bg/lMjWBMzQKTnEIeQph96+
CIO5AfuWCOczGLU3FfLlZvtcHgSNirGFFD4zovrOPDxkLXChNPaEfwWnLyIwJCu9
ETGIfDyszEC28pwknnZTNPKi21fKESP2APO3/je6eIiHLYCUdgB5nEpo1d9LFo1Q
+InvowKb4WKzaesQB6eHdI4x4i1d4rKITqqIzgeIZRqKQsY2FwBfe3VKqclWbllz
NbN4x/Mr8nm9WXmq1Ou81XCcqlbwEd8nz0fAuPBXbDCUcSRu2ktKcRtHF5SxndOV
iZWDfDJ0D8fq94z/Z7cRbQrKysa8ON+nT2LH6kaUrNr1ei3/uX5TSEzi8iJSzH5e
Jj9p9YBaQ3azlBnb8xLVP9X5XJ9NC+nQrd9RIwr6yMoyoG1uyrWT+hcz+GBEuSbY
13Ivw+5H9T9A1oRRd3YDpnDgFOgfG4clpBsGP3S5UGI4Rfh36uXT4HsD87XkuNkO
GPEIvqRM7WzYKuK2r/04XNzcd4oU9ISzAfTAFPOYQY5pO+G3ZSVNiG4gzQ1cQLL7
OqcnW3JW0g3dZwI/5UxXW34Gu/auIsKdsRDUEu9Www31Og2kxPKmPRwjw3lTHmhF
K/+ei9/w1UtMGKRudHFe8L5CLMfHDXNJ4RP9RlIb+/exOMZUP/vRCVKZmiy4AYE8
atH5l22itY3d7HOf/w9m/Eh4sfNJWPfwOPIwKZP1EaElYbxzn3E+SME15dajZeIg
oXZHg9SaIZw9ofYPK+1qhTT4zrAFAmRuSEczjZ+nJDYkAxMootdVIRG937lYpiJz
k3Buq0P/c23vKTMybFQsHf/EG/1ibsUismlpFWZ1iGnMvBLmWfIeiyj7Qi/wBY3y
x4L0oQlRYRM/k0WNgiPva8r0K3pssi5cSMZpOEW4cEZCqhbG+eo/WKP+QIJq09i8
m00gbmfxSzSdXRPQhLxBs5CQxb73Y8ndnPEduSqkLEcNUANuyVGVi4JTd3aU4r1E
UVQSfuih2sOiUofSkxLYF7Zq+ySHjvEwRAefbJnAR+DsEjXwPwM8roJ/tEg3t/CL
/1KCaDq2HeT51HA+Z50vf/Jh21tLZTr+jRnQUQMH5/XAY6UTRUKQcVBQH4q9l+ZF
a1/baEX6VKoUw1OonxqCT34ZG9eFZs+h6Ix4X3Y2QdhxrmUMkPzQM2R5vdOpbGUE
gLRdCEItYdzRbAetr3KY80ssvk7Y7Ut19sJ4OUT5Nr0PEhQ50WPhCO4aRHJv8YRx
BXDl1ATrJrGjR2bF4cVeJ/RTvxNQxBjPC8uQn9ENMViHG5zub9uKVU0vaYItFFJ7
xivzPXaqlnyOE7cMLhh+S4LOh3QZvaUWJvK9Oe56PEz0FTyTWqtbIJDJRpmsMDNJ
cum3SyQGMib1jNmcJIYHgcHtmbcr0lrDmbofs5dEQ6rX+V2u/5dawkxSxWoHstID
Iwy0aS0b0p1KTSFCq9Px9N6vKWGXEwObNBvfYJE7ViOuOgURErOAsHk7o08egOqK
vMO6/FAqI4iiD06WJt8tEu/1hnJD/QVsh31TBs+lUVkv6mfwUTrBgYMcri/JsTg8
pjcjACHw9p+xlRoB+25djDfqw2SC5xqC2ND2fdKqWGOOFZvd4gcy0qrWol5wyBFX
MjBGqSbaW7LII5RSPgSLDuTifNTP+XxnsJiflXvIsrjxTBcmI0mb4nf/VoIV4QzH
sHNE79KCQEpYUDGud3YtC8QL7I72k1jOm2sTPrYhRJNvEqD1GY8bWGveUBxoh8Kf
yrTdfLkkvJiA8Mm5FjwTWQ60n1+mF17gXvY+x9L/RnJkLnA2AtiizLfoOSDK1ffZ
Bn3ny7+BR3h98FisxS+nh5zRLVT3D2H4wkpwa1dWDVgw1vEWReUFMTrqiBbCTCNR
8m/kdgtVPR5Xu46TfjOIC4AweiwzjzkZ3NcRdgaaUHhacnb/PoP8C6dK4uBCBZg3
y4YK1y5oM7WxpptrbZIzZ6ec4wmjONr8jIWVgL3ALeblRl1jaWWK7NPVul1BXpWJ
f6Iy0QQnfgM/yBGOmImOdDxftcl/cUr09F2T7aksqUdKyiBwaU2c5WfmxkjVN2zK
peZORSzJL1kyhk5RRVLlRm91A7G7/FkGPnKTnKfoDV3KskmXRptuY/xuVstnjNqu
2chUjA0G3FMf1ndjkBmx2NMMB2PcE56bxnXjmZgDOZ9u71t9u+mlhNmXoH/7SiKK
NiNOviHqqaIYf5I+xOq46NpRFw29y7XovlWZuyJvCyd2KxQtRfqcxU8Sl716F1Kx
NGmbgbPzVuL34sLKhB3aOTlIpMLHGxgvuvaYPKTf2bQO4lX8XS68E7nw3fVLjc8f
zyp7vcloplJ4iAVGGbbsZuS9kUEbm9akX6o5BQbSGVqwKheyTmNFHYu3AH6HYOfV
/sjALwHqlkWEnV7Knr+5KPcPP9ZLls6R2s1/FJX59xADeIQ3Uft6vHpCGAk57eaz
Jymj/5JRzNC7smb2gaBrhALQcsGy4c5Qnmm804jC57zNCMwLeR230RpraTznmILu
l6kFM2xwjlaa/E5lEbNbsduOzgSqSbIgxTQ3nDKQntHsaZSsMVDrLxzEm/B5Kx0i
mWnK1Uzj6lgq6TesXXLFT2g1DQOHrtW6wzq1qm5RF0bya3Gp4SW+m51O/nL/9BmV
yrS4uSSfo7vhdtb7RFsD43H5Y16uGJipj3l8SZmtyT31ckZpq8WdMvcLuDNxQI9w
J4NGx6ELaZnMoQ2nOTP4ihK3zb5BHHpJvfh2Kp310L8uCGvF8k+CwQPG9HDqcLbq
meZ4jtSii5z1gy1GqYRhsYrcfD6gohASPCrfPAwQ25cSDaTCDHxuCGRD6yxPMfRx
aZHZ7PYYUKRpNUZY9OCr1kXe55gg52K57EAns0LxtOqS9XWR66LrBrAjpUe85fJ1
3BspfcK/85P/gQ2lSSG3rpVP4hQ0R/TuL8H2l8Pzpgr31/iSXG/f7L4R/up+sSgO
/ev7C/CYHQEBrUcChSxEyZXAHN9EGErt49creJpGonoIvbQipSTd4t1Ke/kBOtcC
N7szYCC0fLNG6HkWFPQXr3lVhHBHcsjBs6WYr5qhGICpxrfhC2a8JBd6FQpt/j9K
UDJeks5/uKAobIT/eNBaOStlbBzec8WIOq2sLUYqEOkG64/500nHhmnu+fkibwyf
sGaJyO90LSFYYMHlX2GBMGKk0HQl6Jr7RfZ+pOJm213pu4+x9UWrcHXDvv2oOqlJ
HaZ+qLr3PVh9zGsC4hO/TmYt1tMHE+CYo5iSDLVjZkq7T3qSefA5Vj9dJ1Ztz6xh
FaxJT/o+0uTW3Q1jIji/OzwPsRK9WgBRygLYyoOaw4xbKg4m5Rmdm5l0jkz9rZUb
WtJ+msfvyDNQ2OchXfG1qpW+9o5lY6BU841IWZXm0yRdLRmrmZkwBUoLgCIb5jp8
GWJOfmNZn4tLQ/DBgiI1u6ZoVSt4LKFQ2NGp8zBIJ+RmjL0xOvUCBDDZM4UdZL0M
bJ/jgdh81dXw7J//5xA+44zwTPBj3SJ+lXw793K/a8adMp4MEDHQDrDlFxkiwvQC
GwJEGiaxHmInkn72a28fF6SnsVwtfVgaQPZmalYWwHDV8J7+e5Bb1xrWUeVht1pj
FOqY3CqLV5/Z6CVmVnFMvAHs3thu2jMV9fD37p2T/oMJFgPrIEKIu6psnefW1UBL
JBrfO9Ey2vQuIEzplffRoUG6Wz/HoswuYDqMhipDXlFpESXJZHk2TdtbRCtuQRGF
pvUcUpZE8VYvx6u9ekGizKHwcfNsetvjhNiPv00EHnNUP0502lTtva7rI6ZZ51bM
Zdhyn1xPBmWjaLfIw14XgaIp7ZZkKbEwECrltv0sNsO3XFM6EAidM4W72mhSNsHe
pvSPOhhsZYkXpSwa0EynhnyPpaWxaHeHJ7VXl7cQAhA1QYO7pu3vz38IjsmJDUEj
sUeslUcETLvSvtYrKrnrDYGsT9GOOWwkG+s4I9lE8kHkuSVyv1GUAwld8N7TyXfq
27+mNlcwJxJDinUXyGpzVAEtf0UnCCP3pYa7oM61LTjKfZTwfRRzThCdjPoawH9Q
If9tAv7suwe8k0oM2aL9aBVanTpDarnD+n7nkMUJIMiPmFHUlxItkaKD97/KRAlF
A0Ebc8HXa+ktuQCXmLyVn8YU36GHv+jjal7Y8ugTUWPpgYqQ4ad/ASeCfeb3qxg+
okN1uCuxtaqyrlfHD3BqvgyPdFggGfri7IvjHozrZp3GJg8OviifsZklUEDaNcbr
mferVq50z3wXALNPyFMueaiRsp1wlLIeASwX2EA30qyKhhxd9QHR58PE1AC81JJa
36bycfZRn+CwUnp7A2B5R2sncEd4diOzQDN0JHlGw68lCo2gd+YW1NjrkkzK3YW9
9yNHdxxBHjxCU2LaJnWXsiKQXGYXOXiqDa9HVCuG/lXmrkzq9LKElSk7RJEM5Rd8
cGu9L+nDOHO/4zfRBRhgdWecDIkNJDTnmlKqBaux9ficRplAV+T2OhQIlCluVEJj
HSz6u8U28O2MeMWPC0UUM+Nk19Z7dWhO+qroA4bH0QtTou5v1Zu1KDOjw35qJKYd
Tw9UklLJfhIx/JPBnLdQglQhbIVhA3qoiq/AVXAqxsSOb8SJ/Dvl8PpSfRPUHQcO
dCZ/nxaKSTUW3CAC7daJbUBKfdpBEdkIJs2JtV60xpCc9H3tkPN5c5T/VCFywe1R
SzWSWldudu4bWKCMMhNJ7HAKIrEeaHUOTiWWqQStimMiGTO6XLNPoV2Fi/To4YB6
Xv0j97IJK1PU0aAUePQq4Jp87T7kpcR1JPfxmaaTLxOQzSQKEwfye+NyUSKHxo/u
6u4NJLMnr1fZUWg82LGwaCxi5DTvDfGI931jq3ZNviNLh4+1Rq5PsvPNNC7Sf5/8
yWJj6eDQ0pu5i2OkOT4mJ9tpnq3h2i4jOWN0tC8guQl/3OXsCbodazCvwPoyVXvx
v051/ze8pUS/dKiteJJ8yZavQ2Qtb/82DRlP6k6ZlhwIxJAGqyyvXiw0tXGXCIQe
9km0uAqWyVOxTL6vuBBECrPTL9o7Svh69u8muhwhYaHT00k0/mqd17ztSrmPhT3o
DDJpf9b9mHqnxzySciu9H0lHyeWCvYOG1uAuGNbWIonxbvfyuGuBIgTCwlk6pKDv
TCs6ead44mBgsNbr40CxpVDdYPzpErHa+1QsZDKzMSA/kWly08qvZX6Z2NBEMVMx
8B9QSbcKPn8Ecb7+A3JNOMC9eZdoiffBgQw5RJ88iCjIbnGEF1dGnEz2n2JJPLuH
q5Ea2ghVodYGRp9HV+VVJ1sNgOQ5ZMnxcGClxjU2dnvTV5LWAxusMhthYIzPBZAJ
HPGs4MqOrPf5YE9HdFQmF9bOe3/U8rdXUBlEY1FF5bFXMO0KhbrENnceF9rND57I
nrs1LpBS4gr8hrVS0aUk41c3iKTCuhHzo5mhKfi+NqLu7wQrwuHDNVw1ZBlueoxE
1lj+FYYAMHr7DCVUCF6+7fYxqV6VvsvLn0LMqUcX3szLcNQh3rW6fypNxZIdgtCg
FUgVQVSInSpk3uVukOXLKtQwmd/5IKY9zZaCIr8CsJ+ZKpq2MF7mGh1oJ2INV+aP
KzvkmDnc41Fb8Jhosr0L2mLmOLZ1hyiBvIuC1K0k7aA3HOpTnHnZ2BtV9caFIO/L
okGLQGl/0QiZBlmqbqZZ6cVkXEBMXNpdn3B/+FPuMw12PJXvc1Igci5XaD3I1whO
uHkgNSQ2KLE2XlkgLe2BvwStqlWEwoNZDIV+wmw7oYdXXmw5OSIAy/+5E+4trA4A
ErF2s/EYD8ehW03XDI3wY+X7zGJCkGErwTFlIrwRILdJTzOKrJoF1kL57RdI6rcR
VUlwhVFHJnJs18yBIZlMszj+T78ti+4Y/mkHAqxRJBoFFSrY2Gi++YUYDQtphKz7
k5QKWy7S/3PnX6tTeuPYTYwVGTMojduvPsefG6NfA932MvatJI1X03pBnV+LNWiM
Ri+Bx9Tzic8FM9zRnIJmlB0DfSU1YBIyYCPWEaSkUVpZsRtfHlkZF6OoCOhDkRZg
MHS4x0JYg1Q2RXMdGyWgKk7iM1gDRllt2otpGzGwligmlpr8wAudV/6SGqjcuaTX
wtNtIqtShMgwwkK1TBCtncYo9iOTClchBUkucL3Wbflvg5LymD2g5q8GqlTleHNA
yuGM2gv+MdsftKWF28KQUIJK5+opbMCiKcwCR/U0OBF4/NcDKoefZZeA2CI+k+/5
v0tSMtby1uzpLijN6VMkoQxKi2OlrZ8CNOJTrdlAHdzURyh17ezm5YLUjvTnExYT
Pzv5U+gjpDufQlSkcqoktXucSkMFm4L3qXlc4ZTZFF0+FOG38lIhXk54lcCaJ/kx
58KlskqyCPn/bgdn5VCHIYnFhFuWz8KIHESpDhPy23hN9uD98D7maZVAIxTi6kQP
xOwQYU31YtsgARyZuGU4F/TD5jiIYh81l2X5DnqoQkzlFj8kYeu+yCy5PwhSleZU
YCwFxsTmoYGGc3Hpt+u6Ggq9uxH9bhIFCgycITB9RB9BTGppCz7bZZKGh6K8SVIx
bNPTZ/UhMgJXzZCofCYh5mAuXX1ooCayuQ9CNpP3WC9obOXQMBozj5vYyvF/9rJN
K3pC3vk0FopXKTcbDfDjJktAxn5qGYWVS4I16ZFlaOGJ/Mp/6ZXFPbdXCJ+V2GbE
2vjeQnracg+MX8MYweAzWULK1haB4/GI2Y+T5Fgz0C1/Up6q60DGPc8O095TEwtt
w7XEn09EYUl1wUXnuepFf8wOEzRKPLnZiupNKUSvMPXhlZ8den1GyJg2CvxxO2Xa
WdmrxKQ5jQ4ciCaVgYoLvSfBSK8aWKiYA5hpk/mK1fWUWKzGP+PVYzYJKAiDXGsH
1/NySLsq3xh1GaIP/d2mJFNHSF9wY9380AFwF9BthpIHD1LH1OSRl2lHzjPMJs1o
Z1slGuuLIFfU/hFK7yFvGLnvCfNhegnXGvjG8059E6GnfIdrHGSI6ApneToedf+g
/AA+2N4rBfYTQU1setLTWeHsK37a8Pts1wVgqEkAqCZ68RFerzrZHgZnQiryKKB1
evkXvL59/QeSlB12tbJ45SeFVKznlOyTo6FJOPrNel3qXH+0C478A0HdcqApRffS
G3x8NKU7+1T8F5iRAUtehIrCTpQUmQLTS9RUOZMG5+e+S4O/R66f6GgtypBiRkmx
NFnsgzjT9Kv6cOb3tYdIO/GHevPFT1lJN8JEaByKLEAfQ+1FRxJiP884cF+hsOcL
N7WDn0SIiSxMsmIqOJ0RKJBIVwIrKRNiz0LtsviI958tnduCyytl6ZlXBYVHu+I/
GJpKPqlRwf11J1cldpZtH7vfjHS2COOWh45tsZRnjkz2oww4kUDysDRkZ3sMEeS+
3jZKBuYUxNT6xTo0KRc0Fk0kK8bCiWyC84BTebuc/tiJI93b9r5o8p2YLHX0EAjd
qZoDLqXtYkArf4xDs2MDn3/EiMZhWVmhR4Czuiaaw1fxcqLoMdNy44Qg6BVVr3b5
y3N2gaegMbbAAyahQda4BFE8KOZIXK8b89skqvEPzjEzgbJQWpNOx7m93mCCgGJx
ILlBNIPgwSgn6jOB6Ignyustq+1n5hUW0rUSECpsZHdFZiePohNXAAihB1mXEx1H
hpQDyjJVLpoMbVz/beVNCJGQq/wvBf4VL0IntfDVSOJ0G6WLhSFXEP12ybsc6ITU
EPI9cMDqu/zG9XizaKnJQQI9bGRgaiGMrsi8U0jW9pHdMmk71bZZazc+H9w6CcLb
jyvwI1X20WPKptLXgui/gYmgoRRjDuzMecEF3STYWuQufJQEdtKTjuGVL4BSKnnQ
85D7A9iiEUYJGTbw75WzokaQ4WojYyycA5PMHuEN6jMGunt3GkXiz73WKoN9EYnP
P9gOjKOxvrpB4I9WP5Pn6vbQCxmbBkFQEBlA4r/FKaD3KmtDx1bFLHgX4y2nqElG
GEeiIQA30HzOsBih5UBJDaFB/E1uY1Mb3BaHVtvH9xv7AirLpXUFej0WjMfBku+1
+iajV+rjlNSoJJEDkmw9bKxgrt2X2q6RyWoN1B61LIDjIfX/VzPjpCokjuaJDv4f
U/ZAWXvZqkPb+dJM37v0s419/ADcE5QRRFqDAj+V3X1GPIF/w/mLXhqAPA3Kc1FH
xsWXZrQww2z93rDq8d1l2mVycsn69UzOgIVg4FL31kFzo28szQEiBCu9A+sVF234
9IkObRyds4UwP5QMkdX+mUBSyEL1K6HTsr/UW4goTVrW5BQmMnSftasuRk1Mj8F8
tB44ek2XIPrCZll9KCMd12pVecOURWkWqHbIQC4dLUUHc9wAgUpbnVLV81sF84JV
JY8JH4bY2zNzHDwXzcDP/pZZEt2778eB7x9eppBwGLCcht+GN9akEQOaSnj0yO2K
IP/2es3v6TGZM+ACoUjHoZqv4ci9ZEOIA12b8efpBRy5CQ/tL4xg5FWtigX9xmIp
OZpsQoq9B1JxV0N/9s0smql2Jr2nJipgvX4ljgtnScL+OUP8qEDFPhD16A6ugMvT
WLFG3UH3VA+V0ciNIQykvsTzCHDziot+C6zyFcNrI6ISyVahW1AaYvMRsOpHVBG4
gyrxxxrV/Cv5HHcSyfyJMRiZY8QQa83hyLYfpBEbVHRFmvSoYmxV9iUaBGDGwYb/
2EwfiPkMlR0z4MPq5B68bFTbKwvE1wzuKerddniR1J9UObm/J3M0qr8B1aMHJzdf
TzMJxRRnSLaL1bKqxH9VJx+eWFH5mDYLCR08ysfu0AGLKqwNUoFIM5PINvHzaxJF
hl+nITAFe7ioAa7Ya0QhkFiWYoH9iNmtliB9n0tjTnjRMRu8oc43Zo+joo57Xu8L
HOUV5yxDJgWosy5Mz0NgrFJ/aNNj5vpl9/I4QjzPGSE9l0LuRpH5+euCHWqcxCK/
R6OEclyY5rPhG0Mzttnup8lxSTiltewpPEKGSIAPR5Cd9NwF/Dob2p0DNkRUF+1C
ZYRT+id/z4oFmffg4FYH45Ud103VCFqtOodXCKdxAi0MwD58nwSXh2iL0PVpa4FW
JWbtjZ4z5uK2tPIi0Fy65GjOd/YR5hmF1EGmgFq3O5f/uAjDwsK4Jezv7hOXd8cV
DrEyVjKerGhnaoXlky8oQtZSdiolcSy5xR4aJIpb7s61ey1ClAJRkQ/7yGk3rRDX
b+SNHw07KywFaEKbqZxMVV+mXC+DDNFPOSKzNKybdZ8TSmpQ0z/R3zvG3zGzOpSi
X3icGbQa3p8kgKeDiyKezBmDLxvllkP5YS3ESZlUYUtfJv6BVhdDFEpq1QJ5uBHq
DocpM0SIQz+KHA0bGIb1ZsVf7Ou05B4uV4Q/SxA7LYbaRiexgrZDvtPdj5GKmOZi
riXM778nax3ONGvy/NqQcbePQbTetw2scHbq6mMj0+WDeVMz7jdswupIT0mpLbiN
l889bdwdp0F4VmsbGKkjjJSea68nmjMxDTNV9rc44PYUX+ay9PBnOdvdKJsB37jj
qZyjHByvRq5W2BqPCVndafAbeLVZuDfkVPMUoBeH92YnPpHA2rfDJfxapCeS14yN
vAvwK38G2PhyyMrUkdNq/g+fOQp6HnFaWHxbwGa42TvOXIAgt9UiRQT4Cocaz6aJ
yOhT5kPs+JPUc8QRG2r50EO9kXPM9HoGsr+2HmOzvKFEnP1MAsMZQJCgWjBhujBe
b7IGUTdM35/kj91EHeEwlCxIfOZ19J2NSTW/9hzbyHAXqJPJZ7BlB55ubO1fqxaS
ViEmSeBlIT1MEqkU1yxkEYLNwK2kMHBcyUHmIBQ4nsJq2PcsDMXPV4cnyWESt7Y9
o9BBrwflKhPIcB3UYMmnZ6Fd/L2WqL5/HeVjtMzTteFKqHU6vlJko1WzOwGO2ysB
68MnVEzAN5DUHm8rWA8xKCv9jpxtbnZ3n8/N7O9xKqtZGIyeVarm8QKAqiua9OKZ
SlkuI9Xl0Qv97SwB19hpJ0LTc0sd6yLaizYfpDpTvwcdXzbrpAc5RUmlT8/3JQx9
1iChvl1a9oZhfkouWmh0sUPIx9CGxOLi0iGB//LNL6u147rKhOgkwSStsAhbXZvW
iGKwnPwYxuEwUrKPJdzKM7osvNlSAlAKSWzIkIRMTo/qczyAPEiMY3dEYfML+1Ry
/8V0SfIpLK/S7mpa4y7cmZKh7kkM4J145AeJAadaZDAu7mUsR2FR4/FnEK/X51/L
f9oTwX91daHztKvr988HJS3je/t8A4XGIeaXVhU7sEhmeKwZOzKjREaMiyMoRmog
NRrsZx+CdOpb1Slld0diRFidFa93jSSZuwPWZnJr1wXV9PkTx1PgW2podtQZTpK3
evedDSv0jI1w7Gf0pjz3hK+3fc89u334WzayvA3VySfooXQATw0imTstYf5WQlQh
8Hj0CGdYluVkP2SsN2ypJlUZHqMaSfxen/Xl9Cup3zQapX+Q/3AEUF7FYuULFz94
NN6C+fMgqxAapBBUWeo1tz7oPGu8caj05lgdDxfMjGG/N55+l1kU18gkV/bV5RO1
L+Tj/KisctoqI75IvNESz2GAVAI726cn9qbcIZHRk3UJ6NX68lsgTyDWkVgU56BD
h4wrv4ymGQsdIVB1COIbb4fphrqjvwG1ZGLF1maxaIiP+iURKHnoI5CL8k2h2K7c
aY5wLE/OReslgKwcD7nIab6egqFjBGimKVJgDYFffASQvnzB3ayzVRGdWKlJevSy
bLQYnDW4xtzLYQw7PmwwaPxpjadrL8nOLC2CjutUZtpf4RRBQ6t+sPdMPdu8ZugK
VMjbR1IP38DkrB+V+e3kffllbL4qoW2Aj1hgupmwGiyiyt2XWf1oWddAyNbduE+a
ixe4kCEVccd4GQ/rqdmV4Z8ZyjerN8qmEo6BLbiOxw5xjxS98ysyv+rHrqhvpGUw
7WmqzJFQKQuK2Tqyi3JuaoH0Icdss/Hknav5Bq5GVD7SYDqr3cgCob+JSkR2zKDC
nXREglQGnq46HQxkqb9vnXusyRjlrdLcCk1BldvDs1mlySL+twMC6IvCSrir0j/7
NYU5ne/+SjfEfmeMO6DNp3KzQ0zfJCB6euuv26edcc22Fs3kI3QFSoFkzvN09lbv
nKcdVH0L/87oo1E9ts+oWmSeS4INL4oHlV2+5gMMKr68eC+UQekbQOCjVYxF328S
b7b+2+JYUyIxoiG8+mBdLwxPyzh6qbrdeX9TxrqXiJLaDkBpUhe4CamcJIRv8lCG
ZHy4ZBKlvDxduMLudg0lnHBj0mgDHVOa8idvdH49KcP0/pXRe1zFJqmr94x7G/Ey
TJYym4Y7orXvBB+7lnKeTfgTzwnPPMg0rPVYHE+Jykl8aBHj/GM8AmKtPhd/YcfU
T310kPpsLnrDePzzTx2qjCdyXQUpOwuB7hNycxRe2mkOknHojqvTJ8tIJdEczYn6
heKhzwnohK0W8yvqGTmspc1bIp01qNnOJZGI/XeRmu4f7pGJ7fKKEt6QoFJNI4oj
XnTmhAXDohiR6tPSUTJ8g+IvIbRxee9FNrkMGs/ZuzwbIQR1AoAwl62Y1vwwM4UP
Jkb/Gc0XrIBz5qahQg3ax8mgy4P9fG83ZmAoCzHJeVPlOuBc+ThlyyGWrs6m1FBS
jl4LHwX9pTv+yFMNJY5foscl3BahObIU+QpxIWvt/oSuu+27yXz/mJ7YAR0g3lW5
c6BujfHjNIh4RdKKxAbwBhD+6TfCtGG1Q8MEgnBIJc9O5hDnMHitMsOAEzAIjRUL
+bbS++Kk9vk5a3o0hVf7XLvVY9cREmvfnpKPtEgwh3XFKFn/OUg11enuLaoItSYG
ta7Amq3QYeMuuYT0su8yI9P2IAN9BsmCodJH/fo70ABxOkPnAZC2zvbUC9W0u3y0
vwSG/yUuHjOQACQlidr7NNZXOfO14JDJDZjlNf00sZ0U8OqGKhD12MNjqEmMrDbw
zRUXWlq4gdws2XqJF+WLwTc0G19zgsWxzJyxVCbikXnkpBPsZrOXnlOb/mlMbhPQ
SblsgoXi32V8U5GfUlr+DtpfgDHgTEfwTQiMF+/FsK0pWAloKDDHZp+Pk6ZA8tx5
TA1aGIG1yaU9ptoGA96Hrp38aVTs1wiGzz6T6+hbSwKeF9bsy1PCLW4IhGIkvv22
l2NtCxC5CbQAjEGW+JfcAppPpTB9ymEvyts+o7yAtP7gLBCu5FpB0mEt9zpnryrC
WM9vsGXRGpd6FpWIctkkDZGjAdN3R67F20YO0rh5F+66433kv06hXt8TJ+E1JZVx
ucMueETGBx9uGt0BEl1wCWjChk7vgmGl9F93ySFSE5Tt62JobcmGaykTWMMmGObc
Jbj338eGpE3G+vjHxOnL67qPmcsHHZL6CT09YC77c0/bquK4PeaB0dki+SR8rBFe
sSOr7k94qyC+Iwt/JjIv4A/RRE0B69A2poaFa1oLPY8fpmiCrLxzvC9jYeHiTN6z
gV4nz5pmdxl39fIswOtOKs2j+iuShq+U7ZWioz2gnnQ512W7r0oi0oPGQiWDbiPd
iISa6ZH2yF20UX7LftHVbJs6PESqYWI15Ih4fGw0zT8SPwmwSJF21N6rOsL2qqoS
LKcCTyzkBDarUatj3FuOdbOrQ2OiGhuCCyfi77hTMSTvTamrbvXbwIfmtnl6zjFc
MbFSoZ9b/d387E1U89Tpqwlje+2e3v6CMpGGYAzO9GRcTj9k4v5ujtHY98J/khvU
FSSHcSnPjw5ZKU2TkBR15teWtJuNU0osI7lL01zHXgnXz8hvr8u/aQAWU8b6QosH
RF1bcGB02c7AJZLWPCr3UDUD1epUWYswK6HEBoM7CERb2+7W7Zwqcr05tofObLto
8Fgm0uwpVJjc2sjZuf4PPGpOwNGedXlZzJeQ6138gsDm1o3lbo2+GWFyxeIPCoAx
83qxKSjkbm0b61IWiaYK70aIyG+elcVrmw7UO6zBW+L6+/ovaxiLHRi57kniLlyJ
O2K2hy15uM/l8h7hEW6oifMjW8gb+Bdi/f/DGnwuPIHLtesgJTPiwlPiGcXlNt+Q
1YQbhVZnB+lvPc7PpWTjmH8Up/fimcByvyAsI08xdC4Y3PB6yY7JBtulv9vPltGP
oRwyeh2TtSiOnh+qYxrOuUB5qIE5M87u8br6TqIY4zs6FcvISp7v7VPJ/cuYFFWv
67F3FfMSuyw+AM+sJ65U5dlNgrSPiChH0HnYR2jH8LfF30A4LyQ5lFK9/3hXKJ8P
Q36keivA07jeTSgHYw5UuVBMilSAKl7DjSYS7LJ5W5OsoSwRyLdKtl60RQvEXrWD
JzYWMeJRhwQtq/JwaSLNbvtQDpn0RM4ZJr/gTsOYncwMCUyAkwkrDngnTEXKQLfH
+cnupOkPbo/SBx3DroTCuVYARftmhcjQok0m4dkA5ywejNKjGtuYwQNuTT39UTEx
f1giGycQ8ClIw7M7f7ZV0r1DRrACAgp0Lp2W/XmXl88mHI1q9jipvk8wyM8BmEMu
EjpXnG+4wuSfpD2d4n86PHGmW6Z+sfpyymfY0zTO4Fba2rDN6CLodqldXjtxP8M7
Yi7HaBhw994Nu4o7btrjgJ+9l2s9nAoSxFiIjf39xxSYY3dmz+xlSbdaaYQUthW/
eI4LICPhuaAagdtU1zkiFv695RSPYBRLD2iB4cZaeOffMW04MwD73aXMbHkcbC90
5vFxKNnruwjFNdf5RuGALO4AMH4cqC1mjzAOwur59DVWMCGf1iGGGorT8pUXzD0C
14vAFFLJaaPKOjTIkuEmAeJ57eh1Kcoj2LzFBeYL6OKt1t2avnjUhoIKpSAyEfJr
xoyda3oNpizWNZirncDJxOCR3K2Mb5UMr0ura4TS7BtoLtY0bUqi7QpVlMescakc
kxOndD9SArQXN40/NLYhhAy2ID32Iv+D6ksKyZjCt3V4Je+GMbMKVdcORe9bMA9j
0WAwGSrfSksP/7/eVnP3eP3j9HjP2tYNJdfmaT/7pnYAKR7BO+aIp40UqyadzPmj
5uE2+/tBIPVdkanr0q2MuCJ/SpJcFZTd1EFxZwRq3DyqFwSoqMLMRR0w439dFhJl
5F45OTovecBeSsuPJstzhxXmwOrfg6lDOnZy9oU/cO7TlvsRBLi8CEJWkku20Ik0
9j4zkQ7M1HU6UC5TEU9f6lNu/xHXD5GDkn7sT8Uh5FHMiluo24idtPHw5jsFtAcN
T//Tx0xX69WJK8AQ9PEuQcaAFD2SZArqoie2Ge6xIOULlpt3fIXMmJlTSricBLtd
XYgAF+lCp81bRa5V4/ycZpFSmFY46Mh8VIPANEKzjZlchXTlt2ZRxKQFTJE/9D69
wcsZC8TT/0LY3xN+qnbSbIcUzjswNlfZgsK2jXOpnFhyDDMj3FKOnszTA6piFGli
+vcocw0w972SBDWNY+i77ZO8UUm6leoqFOSTi40rrvudJgoKnPOspSKfvrTPzZbk
49vxinGsr0Xy8Ap77fKuYq1M6B+5gM+MRHr9MCYwSD7DIsqOZ7eg5HudM9NZDvuY
oK156xA6AJimQgdytTKKg70ZWIzHv92QW50aE6LBe2iiAJZaFYBPBZIdPazpRUUE
2tbU/rQgvLvH9nlJrkZxmngyLsjcCY8lTSZV1DO1zbUr7i+WSRrJo1kMX60tjVCQ
8XXPUeije9ZZLeaNMJ9AL7/rlAPwnl4ED+SYPzl26To6VkrXjGDkep9+R2O+uqNt
7mtGUdVsQSbc6FLRlL3kavDy0xOIUAPjVL3Oz6xsjJoNYeN9Sx+Lk373chb4zzUj
ED822WqDgOYLSX53Hs1JyoNRTYgyAAvYH/M7PLsU3/ejS2bqH0Ro4n1pvV2yAgiz
nN53oQc5xZ5YUOAB1kmPoraSoj1NuKjEouUA8z/Y51+6uffJUzf1/wjJd6gqZVnR
JmeOtvPdw1eSLJzzJdCBo2hfilurFUmwvb+rSG506WgHjIovAWjd44yBNRAyXUHW
g+mqq8liYcB+CH6xDkPvC3rYSIO0n7FQj1qLTkThkZJBlSNFIqKzckUDPsWfLRkc
CPckkFA1g5ho50gkxP9M+QSu/O1bGVIdffZKx+YiHUZSgyiZHi7TAw5OY2jpFkiJ
jDGpPYx2l8VQjCRyhHT3L3wcDesZ6bGyjXfuO/zJVpSel3S4XzIWrdaI6hkduoca
z1xne1eAFlByafsCIH1Kd5LYrSEeK8ZrGebBg8gtnKTCNxuHilGZ+KB2KQEy/cDW
D/Pt4iSS31I/xsECSHD4RGynQ1r+u1Rer+Td5pa4J+HE2WrEqiHCFE98P30H5t8y
/rOAEviZmqj/MxuP1hw5/tH4v0mK1Z4ckUAwhLC3Kpty45O0mdPH1vbod+i+o9bm
SKJz0HEp0z99Ri1dIIcqgSF5wMjFybKvmL3biKX2UqtaxurfxpJN+G9AGPD5PaIB
zmkcdchWheXhtuMGMaUngggfhPmMM8E4DoR3/gubE+uLfmUknFEGQz0CuaUXCWXl
lbnkrZrwW28MrnUpz2YqkVdCpqi5ct8lztrD4hJjM6Xn89NB7aS1pCZZRR1jX3MU
oG7h9y0uyOS8Dr+rTe8D7Jnp9JlYi/bT4RpLsAM7JQhkq1hCx0b8C3QR0EmelqB1
zszxVV4TucoRb3Ds5hs62eyR1mY6nv3o2ryBV/DllarmXsyDHY7BRLQDTSqby4Iv
WufL6NmSdIzyf08GixXq3b4LRGij2b08WvHlDuIuy6ZfGrpy3gwuNlRwJ7vwiW8v
WDBbiT1DNP+IJBZXB30PXLBuLksxWdU3qxAaTDhkVHn5ip1xVooYhQkNpHTj55DC
zZRolLjkWsevP4AzIQtoSicg0J8UqK+w0211lw0c2irOfXugRlNLJXOhR49iS5oO
snjIzY+1bmTLuxzogNxS32f3J2QakDjZKJ0AfT+g0Ai00z7HQSVlEupoV57NVHx0
R8f10i9lnX0EyFYhMWYDWnV5TohCgc6bxGirjiCeEEIrEmQJ34SH2tq68VlAYaGu
cvTI0tXCeNhyNPf+apVQkY6jkgae3EB68Cx0v2GV7uI=
`protect END_PROTECTED
