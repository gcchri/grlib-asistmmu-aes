`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sui9x8ZkxZIuavWweoDsmiKZv6ow8zVklwhb0IHM7wJRpSf4u1xYbSjAbJh+Neua
2ntvedHVxDAVyoFgZT6AOrXA+W+I5xcgDc4yTTvzjLsKcowArVtyBt/G4IfkWGZe
KN369xQ6/Rk+VsbSziytFsy4c7rv/qcWcntwDZd0X7pz7/XbclMB1zy3Q9unjKE2
Alt7s9gcWvm1uszg8q7iZyqBXLH4NC/VYzIMGdkp6lAa5w6dV8iSiRrTNRj/QzXg
D+7nmMk/VNbJOYtdLBhnseaM9wUfIqW8asxNRbcgh+pFrWCc13q2dG83oSVqrWc4
JcdIi2+zp0PtNFMrZk8+LNPo9O40p9i/jMD/dOkQKJ4CcO4Sq3bKML48xTRleKo+
1r0lfFoHtYhGVXm3Yj1Fb0eWM5s0e40E9Yn7hhSqd32hL4y89mVNRkIB+Q6MGgQ+
eCUuVTZdTj5AvS9vjC4ShN+X+ITiC5tEkYH6Zu6H2VOLiD+LtRjn1MZIe14lORwL
Pw2JQVFafAxGAvkyalZMrabN+dn/gwz9Q82TEz4GPguceJE7iphRxUa3fxGsY/Rc
0CnogMkLJbHWSvDnSTv1HNeF/bPFYzts/Yj3AWdkdyFFovmNXB60y23dIMd9FfQt
db59jZ+eME3s+cOwdnRq5wMXRhRG8fWd3ySeg8f3Dg7uq4FCz032zfi6UbUkHOcn
6BNaAEKiY76xbdHhd9RaGJk+7AJYTrpVlSIkdwtZLk5ZYSjArBe+5QYf0WlgVI9L
ZnhSBb6YWhy/875+2qCCunUsGjFBTdoeriAuzoqVeY4sZHovj3Cgvb8Zj02/dtA8
olQLYIdeQWd33qrDj1u5NucOxJlhcGquwQUp3urXQ1QJLbcN0NqG75Y9Suuyg5or
GMxdFiRoH7X3ud4JWo2s3YG0XKpUHhKUFmYMm+5Mc/kJihGoTvypQTgmSMUi2Tj1
ZerXrGYzZZqCYip/4QMurPpqFGmNTHCKTFDC2wzu/HKXle8q1o6SLGumFHiv1ImA
0sNxccBL/0OThANxeRk+2PI9IkG3DLLmy7sqS8NL61rgBRuNjBNIsLDRoaorCi7E
+mHnIlcmH6EIbjA/dkpfMhiFarfuJsjJM9D7oFpnx24N+PIm1JR7Edh5XKLCkS/u
BaE4k/EHyWtirHro83juNv74B6rVj7hsnAT4xXVu2KcOaa8K+E6SJr0NbMX2fhT1
Ff0jaYV8AU+4MjC6/dxxdBS2uTDllTCWOhCF2j+8SvoctkL6V5XZn7AIGJv/Ikyq
tDQXuYK4/HnjKot1NClz6o5P3RSHVKTuy74DfP+hnuCISavbA3DJFSs+36zaATsC
SPetWwQACR394uyAUTeafMYreZbFIK6ODrECrXoDrJrc5NdtdFWM2E9jihIArxtR
mGeRIG677r1fitY+iwj4Q0Ts9VCwLqmRLvVgjnOcrUKC+g86zJu435d7qw0EK0Wg
BRhsJ6Hl/hc8G2dwaaukzfrDeSAI5dm9M1MoAJUXyg0K/hDz8lWKI1sR5018Zyup
oapyLo1Cq2PycnTfrrKQaH3MdrEV12wd+3wY9oW1Wn7i07VoACqE3FwsMRVqbvb2
9k8q8rWnlOx5mRrKMEejjF/aZvDtnKyC3jqst6wZGjacN1DLf6ACsuKGbI9Xzk0+
BRlRTu6yAHmsJrC8jcSflUrKimvhAStMBjmEfmyMHoE9OT3fneyUNzqxTVazOnc/
uW+TTMF4UK8jiaHTk8kMbl1fWQ7xDqwjr2XQlixdhQeBNDTyb18Tbys2LNU1CKLW
DgQAqEiCQg7k1XzEbThFoMwr0xo3Ae7laBQjO9WYvH4/4iucGujcV6tLnW+u3B9A
0xuuTnQd8kHgGBh4MeiTlJs0I4hFYsXWCAK4H3rkG3L1s8aeuqMqXfXv21HUW0dC
q7/Ggx9kk4HALrg61oKU/4nTKtpKYZn4kZjMBVqKa5QSVLMFl4tB27Q/DcxjSDtO
Aii3VaLWp/GxQZji7q1En/lLrbTNiJiJZbZxcCSsnaUqj/OxE9JzNrywRLPZouwg
LhAYqo0yW2WrIlujmE2qTtL3HUyBZyS25g0bru2DjZaGpo+CEYDqa3uv8FXCDVfY
TtWxncFf88abZrF/lYGoJyWWVbH0cdaTl0A5GsFV64xau2dune7sz+szZkZUqmOW
tGWLLWxvO4i62aERapP98bKGdDu+bPR/5QQI5LxyN8Wknnbh0Jw52xaOKsUsMCz/
qs4Nlo1g0TJklxlCgqtcrWCJdn6zxVY2+BRqaJkKbqJ/VliI8N1Qi6Vdq7j061g1
YNh65rZUm97dbMcR3+AMCz4Xojua9sk7bOEJTPnO4jcpwyNnY9hgF0dL//ZGhQ0a
`protect END_PROTECTED
