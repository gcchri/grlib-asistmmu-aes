`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GVMPooGl8LD1y/ItMfp6V+hT1mxDrD1JJyh5fX+3+WOnJivzj0gOM6Jvidjtcpq
RofRh8NZyk4iK0/xZrkJK3GV7RlKerGL9x+3bM4a/ovUQ7ZzR/eGOrmjnFoLGX5u
rcEwEbM5Nr19ewYjSmfGLH9t3ex45yEb4HyEULHgE8JXx5wRIrXdHyzhcPqcm8YU
j8bvMefW+Fee5nUMn8Y4fh0pNT/7VSXNy++QeY/04jxJZGbUBbQ62vQlLu4tr0hg
KZbIbQpVp5Alm4u3G6OfBv2Vmhg01Pp5cQC8eLfcMZ99bdo3MjlFrebU47fA+KJ3
+E6llVXpU7sDo4aO3VF6pb6NzbRdMHop/mdAmVEEYtAF7NKvuGmbxe93k99OmfOc
8nsUFl5/aCLkMLjbY2y7uf+Bg6MqYfLP1Gl79VdTOXM=
`protect END_PROTECTED
