`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4eqzFHmsgVwjLOoMr9vv3CS0jy46VkMMgGi0UudA/Kpod1vluYfO+eNjECeeD4Ch
TkdzWqLz8X6YljlFYACsZKVWfC0Db1dL9MPoA8FeH4p62Bxpz8zzhgc7JY/OAXtR
72gIzKwUHwETzYCyu4YNqR0Uj5k96hvnsAlzaX1B+YDHvOhkOC6HZAbbzsObq5F0
MvANPupnWYPvnM0xL6yY/65Of9s5O5svo4M0IHEAkgNoIsub7OdS0+/lkZIU4DFy
wDQH3rIwIt1BvnWjzGkAEtog3UyA3MHMCFmxyAQPhFfxU1od8EdI76P7lg3Gr10r
TMlUv5TNt8YPlDiqDh89M9shdWSDMbF4wjQdOB9HOkeejVHwiA90I5MBWIa4gpjV
oZNWXIAwn157ykjfn8Ek6/Vgwi6paakaUNRqZ0RnzBuYSCKOWrKgBC2o8oK9jrsF
7KFIVuxkSw1yIMxcP3Ko2yCQ5fpmdT4lRSyZmPExv57ZoHzqpKBP6K67QKkafKHw
GZKGlrZycrOpo5XGJdcVizZSCxqSUgzi/r6awHjPZ/zyo3y7yv2cVUip1wfm2nRf
8L45Ip4j+iQY3HDh4mw/fBBodra3TC9UJot+lftpbNmYYyGk9NT7W6RhsSdOz1M8
SsTcTwGPHGjZ1tzIypJJLv2XX+l/LVKQPO7/zjqsEYsvKAt8LDuTi+YKPtvWNKVX
dqQ5+t7OKo6lu/wt2hJPhdADDTHMYrITCnmDRHFXA1R29cC9izEBDY/GiFG4Rpnz
XV9a+G2grNuvSEE6vxA3k3IydYtBgyZj5+Zf8Wd5eMdEJzHSmlZM+sgpUJjLvL80
O1todsTWIQjc4I0AKC00pVuiBb3CEtx8rDB2BuW5m8NwWV8AS3Gc/2sNMGKUMcbi
4ckCXfXMJ9lVDnWnzXpWu6F2FsNC4cJyRmNldwR6T/cJL81WZe6jmaXHHoQycSLj
edbdzSEHimGn9SAjb/TfGCjo3oDnY/cUn2+ofIkI2TJMZPR8eq6axNB4wNDKXB7E
8wxgi5aP6m2CH0tn4UTV0qCawQ35L7SJISP5mOR2A2WPCmmC7hlylv7MOARFYT3c
rui6eieVbSZ4jHtN+WEdUzRUmdt2soRz6yvBx8WL4ZCo+iBQwx0+ObZ16VIqwFcz
3+iVjJIjHpZLv93fJkVhi9rc3/Rwe0EoZrNx4oC5OHdRb0k7zuZ9RaKCa/ZP8omR
MJaFxK9vsMW3r/xqMTp/o1c4/YTtROp0mgqOtE/ITzzHY5hKh4sYEZ5a4PgMWjNv
5OzWeS6zFr4wdJt9KaAtSnez58WUfYBFBeRls+PQSO12/kCILSrXANFipZe8gLlb
P2JoucEwKXx9miK8+TS9f5qA4isfUKnGH/DFZy3qXYhDJIQBaQIah90N3JITLsgK
cM9YdrAsQ5abppR/nJ2looLYrqRcVGGACGZx7DAF4/FP42PHqouvSXn6FzuiBki0
K5hVyZQrL5xypbebcn40dniKFhc3LRDGSJN6prbe2wlDDV+TQ+XSEqeW69T1Egfu
KWtyaaqK8ooVkcZafb/2fwbNm1EFiV3PuTFY+4bTW+iHEnjABHB3HEo+X6Q3znzO
BEsxuKvORKzhyovgCvXLgB3Ym/Nzvk0nkWBQlTAd8fDjq4qfGAsB5ftPEPRrp3Np
tvurOQyW3xUwHR7u/MObMGQTN4ZXNb0ZvOijaqE/77LfXqdo5U1JiUo6voZiYukv
Rf+ib0flOfMZuFi5s+AVb9mt/x6iXAfU1AW7Ryw1DXWgtzyRRIY/lfuKCJxL9ghN
HtFN7GBDSLFuwJhC0FtwxLU7Iwvk7aPnnUQO9YWJuBUC3uT8yxLDQAob13YLLZRP
3dkrdP8R3nYrwQp5ABh+iKTCfil8rm5TuXISthIaDc6fZYrgWtptJqd5m75DmI+9
`protect END_PROTECTED
