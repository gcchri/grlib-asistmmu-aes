`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0OeMKTMExMttyInVOEhYkF0/5a1A9DSVZqNN8UfFocAbFj9MvEsFEt76OQ05/cnb
HZRm6HrW67kuumZx362H16ZKET0+xgMoea7eApf1oZYnoq87oKFqLv2PO/Cd5Y+8
Hv2KctpbfqP/EYkDZ5wWXtEod/ELPItQYYuVuESR3t4aIPDhYkA1X7rrRlSEDPTb
9rMiedIePddQczYmC8LhH9BF9VFdR3teNGwi6L8XK4OlSL0XX/ZB9aAe8K/jTtIO
qM4x4MdQtu3XbAgg0xpyyw==
`protect END_PROTECTED
