`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PuiS3DIIc/QGbT3TrAp66ffL/5Z8pzs55Jl05X95q9pk/2mfUBsw57jnL/neR2/A
2FwJhaTIZsXop3sSjNG2cEwZ+k74kchVsdKDUQl2Gtizeh6CU3Wo5jdT7L8qiXEa
fvJeuiAf+e8iQAhMRSMpMP/sikdxCwCe6BS/cN5ldZLP97mH19mUI+zlT/Zgx6WV
pwrEWtuldx4lfHtFxSw4n4+WpA6n0qJ6Vs8UiEd/KNLXi78S2T2lT20KzVFbEJqG
A4gSUbRvIJQDOIAZKj/MaGYI/u6sL92AVu+ZhZRXo8yVmp1vNXx77Lk8ZIDDxt45
g2jFQxRwpPWMO5nKic+9XtqS688p4AXr9mgXEJvkJFQ1d/CfukMARUAdLMB/Pby7
95VivnP6vZKv2ISawYyMTpI85f+aYRgpdgKQCA+s4boq7iP5VbNnRTjDK2eLHsvh
4hqpPFc+wpMHXybSUWXoYxQ0G1QFJpPg4AamNUNMMs3GMwKkFXcOcW3QLohVtY18
k5pqeqIoAf0ZNi0yiYs2YwmX4nwlT8BF1u05mgVeGDdm6cz9k3gEVzgRtUbBq6Ow
UEEhuSs0OD3Lxm7QoiUrkVPf/eQHTbXu1bp0xb2T566Jush1/1eVDboVgocgnxET
vCPFQHhg4c7NM9RlgD79syiYod1Pil0tC3gUOEqPV/3NjQPPXRFV2p9x02ewMDhl
1RnadnMeOtIoZD0KQkDUcRP5TgYzF0zY5HRxDguMmZRTjXbfKsJtok+X8FyZEdap
176E/fOBdL/1F7P93Ouu8xvAdh9DI9a5GJQ26bKqb7wiinUI0o9+JCMpcdqiK9p/
QqZIN4L+QbbdHG1+6TVJlzQ9mGCfJ4w5Mrb6AoUWzN9TuCwWZsZcyjqoE/cm4mI5
uY8xoWNUIX/eD7KhPyVUKVBgnaLeACHQxNKCajnvAzY6laimd+MriG1rT8uWyxSE
4fyMzzTJ/PlaBotRGLMrV7DklnlJ1LDlkfiE6lrtRsiJo2J2RYZOTpam10GT6vmd
pUcANQmScnoSxIBO7tH03KuiPrZWW8Ithpit2AwUaeGS64XGSqEdIRP+6rYvqnmM
e1Tt0lF2AETSGJtmKKXxesDzbbmGckAOQfwMd/Ms5tLHxHLSgAX7tS2OkLSgEGLF
JlURHS+sJT+KPwfnnK4VJQjbW40GbBd6oIAESgBGllujnr77em5YLknjYwDUn36V
6i5maDfoDdMcSjtto4SLmrkEi3UZ0ZPcwIx1Npcr8llkJBauyvazQ6inNNPLPKHJ
2RKlFzIH7M3uoY9N0y12W9/20rN6ZfQrrYTOLjB2h1PwBkqImDhydqqG9ltezTS7
hJiHrLgGDNq6kBYVPGrBlR/WZNgNtp9w0OuDGK8xf9Y=
`protect END_PROTECTED
