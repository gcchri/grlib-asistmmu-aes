`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKQdVY7V0/eLQEuJz3zDAMsqxJV+NaHkIFmj2QSfNBpKNKwg1xCcpBkEH9qm7V1h
KTNeqDE/bkl2e+vdQh1YGRJSkcH5vFD8dBILwJ/FgEuksaE4Pu7yi0dJHse5P8o7
s2B8zWsek94UrgCMViZgtvY1xYZxqe1jueJJ3Ek/6CfPYnk7ErcSPEow0xdcbHWO
5B/2uuy8LG5ctRG6OXBsQc1uiJAQuDfvnANI6DnnWmU/mA6soZCa3gx/x+/BCMz7
Z5Njzlbdp5mM3FR38r5Z2AIZEIshlQ8fe3EzGrYcNkk/vke1yhvO74hjLfpr0axr
D0RCjQyJ5HoQX81gJXPUNg==
`protect END_PROTECTED
