`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wivq1ZsbXA6vOa42CQq+mm0073aA9xFQuytgnfzb0/nYpk3EuPRI4zXf/NktO8qu
U4qun87RslifnHvgbzVcTRi7teRYnMXBLu/uDWOwAog732N/YXnao14s5SeOeJ+u
djeBrnU439qaUR/bcsZMK2Vcdhm3A/9/nRKhz2wTeWZPGG+e63wONECCM48xgBBc
MOsSMQtEylI8azqasZGi5JLJT7jM5Iwutyb3Qa9YaUR3+sVFlbninLO2vBJ6uOTQ
SM1KzcyLdRotgVodpUTN1PLEy+MrMwLBcWHrlYWTzK3r2hHfhfuqXFOjZQF9fGpg
VBbtNT9zZs8n/O/01wQKVz8kBrb3V+hosOLgW0sYxBCVX+pi+XcAyi4uf9RxLqVz
q1P4MFSbQgyQCJRV3fmD3g==
`protect END_PROTECTED
