`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXMr3+MKFzpx2x9PynQE8jQN4AORMBHuZYS8usK9ZAXo2NNSyIp2qIOg01OHYrjr
gPegcI1IkZnhllhf7t+oepZvHYzscI9saw4OEqtkh6L2gSOdl/0f79HF0FC8Slly
WIpSLM3MPQSQqVj/m1Iin6UdMjhO6k6rIr8URM+SuXkfb8tB2fWcxGTgHwRWl8wP
ALjl0v9PdlvjHWR4SXoVvLAJxoiIQd/7rOTqngv6jxZaA+aj+7h+ilq25mjJUUa3
F5pUrTRQ+jXNZO5Jg1e4VQ==
`protect END_PROTECTED
