`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ojWyWqYuxJUQ+Th7GRv3XEroQclx2Hr/Jipl9o6wFfEzpNwajYlfrfr+wTFd4qgp
1mPcitpwRXaPn8gompxAn8LtJRHL3pGQbSbUYvLgV0I0zPJuQG+cnVH5t/qdKNO2
4dxKIIVOs4iVmMVWqAWzigM6VB07QKxdbHXNZN1tuGO1K7/NLS1fsNKn4fYyulIL
00r3nbhmlT4/+WwkFBUcy9GUAnN5thiSpwOgmJJ2wVsuKTK5i1jRswrdwHnzLFsi
mQojJ2H3JdpICvcpk2RNENQ1bMDgdgYPAJTTgOmnffto3ivD9GWuMOkqfHT0mByV
GocPY/vUYw+2rl7LW3lEQDXBxOsG4ESdlaPhEGsCcjvVwjLUBHOYJz94BOsdUr4H
kMKmUbpbceaDf4WMAi6u5w==
`protect END_PROTECTED
