`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1FKwbEMv/vnAPfm59VMq8mQi/4eEFqOokDbRASV8pKdQ8Zd4lzzEdgQgwMcbJHW
HN1Fl31N+r5olLQIQMF3PLobHRPG/NV4RPA1cp0Edu7WeAs3fJGDickN449hA5Ry
+huR3qKpLE0lfLRAGNOVz4oy4hm5jaqBMYr5Svrosfwr840/VPl6wkiKKk0+yMkV
3RTX385PkSBC7JWzVDMuz0v1Ljn1oNs+I1eEeRtMZRm9DlIeSj7ChlX3Ovi/0XOG
+c4ML4OIQTsEJykTFl4qkb7Jcct9Ze1pX+Liuhap4clR5tcIJVBPxxUCNn+NOCgU
uAWCgJpvaKci08zu9Gw2YvxSwVfGnP39rDY3vNOAaxxPqzOkI3qy0bQcHBlI6llk
oNC3OLOv2pSMcJEOlGqYkpmO2epomMSs95fBc7CmD8FTl711cziUH0MkRqxqorij
`protect END_PROTECTED
