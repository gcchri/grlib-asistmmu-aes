`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSq6CIAyOn4nQyi8eV2lsq+KzeCqgLH2xBoWrh25kf3a/vH4qG0NEE0PzjIyuX0T
KtiW2Zhp2ry9f1zMnZa2sfyxe1P30hPXtIRPRzJFn34w7yMNo0sq0lteeoq+q6yA
rRZMS1B/R42Od5YdLdIdmHqlrtFA1dAHVO7cr4lVmk3J6EEc1NirL323fEtrKGEA
2ezkluUbvMqBKnDGmRVJbNUPeMBbI2ylAeZMaKLw1xVFTlID7GzBuWdMI9zFTCZV
QUvNA8r5LupV8BSdMcJOvUtJfrVklZ3tu9ht3EbZUXXE7zTJ7RjXVITV8hvnYDrj
0j7ENnzQtQyqIDNWriUHsp9gBNv8I1aLBnkzK/2KmqWlxHmrpDUrgbiVGP5Lwky/
F91SKRKx/l4/rP9R5XAXoJ7jzyyNeUmoGmV9McGvXZnFCFI7mW47bhITYqsbnvfy
RSuBT0v2c7VlBTNPhNA0E43bhjphHtosPIXXl9LSgoLsCe3ageP01PWRYm3wt4Sv
CouMhevoTUz+c6QzDbIwTTqViWPgirAMxxJfAe23Nmau5byo3T2r5aONFDHzzZDJ
3vGzrtVc2BE2z3bMErygJFf4eXc1cvvOBlJRw8zCC+vRy4VtqXwOz5w5ER0MqwGJ
cMZygTsjQFbdj2uR2w6udeZ5z1TAOiIsWY4c1v1vDzDRvwcqcbcBnXnyz3u/LHRZ
tYq5LHYJIyCtkyOcCII6gbjwSzGTQ+NQSblmjeq/eDCHabkBB/cW62P7iNgrZ1Eq
AHxGS5B9V4lrwCFKHS4thCfiATe2y6dzjWxFRtvXXjW3HRcXWq83cMHKwf+3Y+cz
/QDfTawzVne2GaaQvnCcVGRyP8icOvDIIiKxxHU+0tfRPuG3z8tJdYSPy7tb16Px
U6FEh+NRJGWG11/zTG8fkngvbLaXYjnHWLohWaN3Sz89kmYgcb7FqILkvcbNl9Fr
Ib5VZQKbgGN/fe4KWtKyLXlZz1nZdW/6q91xfj0gP0ZqLnBuUSxqCGPkQilg8ZiK
7EuCVOgOmnu2NZpMMduH5pnW6yKC412L+BO2GsEvGCpUWdXeCFm6HVkzFZJlKsD4
eAD6FcnxwAV4IJ7d1sYeEY5i597eXhb4vwIIxY9PcNHxXbDS8vBECUpTtYPIU+vq
+kbRmuKk12jrP/G+zOXvFWhCS0fJdk/pgwApgGmhrx9SWaag3NvBe9n3BBmzni1r
oWGJTpa+VaT57FmXIMNV0ifJw1XgFN04gJrpalmrpPIwObBh120QlGmcrSgJOT2N
EOnw+B1YnK0dV4p4OqQsJMf+4Cl8iD6aBW07GlhTI7PB7o0CW5v1IlkdriNkC653
Geos5iW2V2nvcL6xfmyvBGNvTmLmqd/XIrAgRIXRXO5Eyegbmz++jTxtuhIZ0KKm
fk4z8c8T7z1i1OIjHK31hxZBCjqHDq9J8075L+6kuhUZbFr4RJhFDHuVu37k8YB6
CBb/uC50f2GWcSjbMweUQVXp1/iWJJikm9B5RyfHiGFxgr+q/KbF0SRbchJrncpa
0oBt0eU5Q7gjyoc0A/mwswpdY+fh6RcAb6sOY6zHyANdBd5Ko4boCoVUvRzMgaIE
ePsP5SuDKjWm3J9GnUSo2lH/RaVHeIhP6mMaqeXEhocThTAIADcZGNdS8iK3ApBe
LaOYkNiP/r9b4/6/2+vpSOoxgzE+t2ByNPAEapTVE9xetL08aMvq7ZFA4PKoeef0
LY6v5+dJfUaX0p1oXaexmVT10Wcq3ScwK7SU+y16j8+7l3aNDlBSdAIjFA7N/MOD
I4n6gAcbs9wqvlwaUKvzFKCpKwZ6i59GAGTi8tqGlZwfJE556+EQfOi3J7GQNW9U
PuxGwSuhSJZNwo1KdgeKZnp9/WD29kRMkeota77euWCKEcjWKf5njdrG3aPuQQLN
vhMnEk5cxskdFhDPOw01daITajzL3xcY88JT025v02Td/gDZcdm3F+jImGv649FE
GfPcTE7HwLf/+ldJcxRTS5QlQQd6QRWSsCevwRXDU2axYLLS1Hnum7KvmYEo07Xz
lIT+mU6xopyS7/lme3ExbpoaKHUm5pmkwxpeRCHSe60+pC3KInt6fEF0/cjbRMzI
zv3BDyTVV+BoTB0n0EfLy9NatlrsDoktiniamRtzW9nGh1n87vL4DZGx3TF0UcoN
DhQ4zq8o2GjorVaeaFCzhNce7rE6BtKXUZIM2kY4i8MA2Yy2lkNgUVzLiGruq8zQ
I+hvdzwInXVX+0zprgq3LN4Ab397czROtbomyKnnUnuHS+NGUCdeWOj94mdO3FD0
RKR4vwfC33yqHuKiWi6+OaYPUZGQxVxvjJ2cKhGONrmh7mfuGpTQ7hqmBfMaTPcf
`protect END_PROTECTED
