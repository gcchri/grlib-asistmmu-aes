`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmJ9xdWuSU1MAvyNOqcQQrtD3zHeT9LkvC5cutRMY7ZsKvhtkbLb0cfKNvXNnFFz
C/KcIesZBBpLYfBYMCG7FE9o5tu6mjSh+5jzvgN+Lnt4ggyT4GJ/LTo2g6BCOMW+
DZtPJ40cHmLmA7qVmiMD+S0aPPCdDN+FzvIRgpUqSzNiPgszkCctdrbIkNvhMk2Z
Kn5dxX15kkLW4iOQqp2swjJMwoUvkDqfx6YoADtaSJtzmxaS9HxfB0KuxhX/Hetv
nF9WocJg6zNxvjh2TUslzTmIy6EJov+fKx7hEAn65y3YGlHWutn6zLQPzzTiZr26
r2iGQe5/0VaYn/XPoCgThP2xfYtVeEmw92/OI8Uq8dOfdaYqn/L7vdVNxNlwY7lk
AZlqMuPwRjfXo09LIx1uELcEOfzw+1dEQn3V9dEpLfM=
`protect END_PROTECTED
