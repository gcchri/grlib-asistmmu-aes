`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xt/+loCwZ97vJ1UUR4dh0MHjjLPHYxoPT67ByMWqSOAuJ53x6Ey/Sbt+QeY7z01r
YNgOEn1ZrJj+bs0PIkXAUnD6PK5B6RRx8rxlbpEz7DMgnrVA2/m57jSt67mFaFRL
DVBaTigKan6PmsyvbKGn0V5TxVi747BdlHE/ufSWBOPbhiEpd8m2t8odHO4wFx4P
Q7nm6vEma6UofK18kRrgbRCpHkF+xGUF1nfwuykWHo2K2lsSF9lBzpvGK6efy9M9
QxJ94cIC0i5A6p+9WTxCVn2UHsIbv2Ui922dwqbc2dhAwLblXFjEvdrIaM9wWAT0
9ZxM898HmYU58TdJCSZ4fYndYtp4tSX7wS8X+y40nzzxU4BVgmjWhkIRkrmfDbnv
/sz4V/A4um1AIwKXZJxowlUkyV7JJp3ucRW7A+BFTl6i+ml5x8fSTeRG+btCE7qI
`protect END_PROTECTED
