`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N1Lrm+4Yhzmc6fxCMMLsQwhSaZLSqHm+dSQswj881ejaX8yhYNRMzZ3dKaM0FsoB
V8dH9tNGbPt9iEN4/6wY5TI7MagBU2PhDQT4PnQNnERdAPAHjsXFnnnz7734OazS
3FDGzvz6uspDgNjErEhCqnssiNgl0de8BvDqwc1f38MG3E6Feo9NKyI04JXyRfVd
eh+udAJ2t6NMwa/MoSWKJHSr3CcmkCGzNrOpCe6+c7+V4ycAYqOvlYTsHUIxgwEB
FgkIeDHuYpOTU6lnvqCs0Bu/82NgYW9rBiG242vWM17PDtSkKYXsjFJEFrw8dROO
WwKFBU/x/isRuYDnZ5KPHwLr7TUDeNMMSwzuLzsV50B/NlDwfSOGIAtX59jloGSf
4IWf4S2X+o2z2aKMjdFfPJorLZ3Lkv+yQUxw6BWnouQBmhf6x8Yu6w6bQ/voXgik
JicETux74TjbC4K9hLhTt/wQgEY9RWvbRy5PfIb3DqV1fB3kIfXCVYhzeYfGgSW6
rVKXf5C8Jt32V4KNv+g+vpqeJUVp6Q3JjNuzsGkrhlUurJASXksZ3Thqk05hQVzx
zyA3h9nE9JJ/F6vsyqelgfPM85BH2pd0hHCcMAL2z2t/+pdzd2G7JiVZpcNz8TCM
BBBc9fhgIOXcb9PSQfrp5n9i4Qt9uGOkZHVCHeW3tWGC+yV9urZf+N/2QfmAWNPI
3mG1pziyNMi3XVull/iKkmCW1S2+T5vH3eBWEqsa7T6Co5B7XOd1dVUtOqJVgf0e
7Xtm5t8JQlptEmQc71Sq4meX6Csf81/pQUs7YqX3hB7Vcw6uUIYnYaxv37YAGeL5
FzmFyp/O+GR2/nUex5WtAkl9IfZwsbOcSaLHKzoyHL9VLZUgYtK2L4tIhBC++5LH
Pic+qoxzqW8vxvRISKAVNYN0JM+QTYKMg4BiadH2iOmUOKTB+j5+tikX4HgKJ7yS
Fy7d5ZnaL+MifrSDPXWW/t1c4ychgM0nD7JJSnCYF9GnpVy/I6+2tmVykD0sIAoz
FUaiZg1Hr7BO9a/bbwAAWGKpsPnFVRfqoghEsMDHRVQLMS6c6IljgjbypmrQ4ufr
5z8ckFF7plh5fLq4Tf6d0svaxGJLZLkZaP8zaEW7IGC8QZ2xg2yluzRCHxabw1MN
JXt3sKewLyWreq9vn+daEM6bie220FT5aB+KdduHnFKK4PcEdNTaTKBc3aSl3d3h
m37v93b8SmFvcTgVYBPjJ7hhz1JZCNqAGHga1moSK8tRPdOJ1JGcic+EYEWiXXZ0
F6xtqNZRpbdaK7fIIL2kmF+I5tPpO9do3mJU4yhYu55gDrEgOPVy3M5bgU/ldqKS
wk9EeaN+9M1WeEcpt7kyfUKo8GBSOm4eFTplCAgOulOOdSLSRdbEvK/IaBw6NU7k
ws3uSEZiMcsjC+p0vnAjhNgmvddDsdwZ/nibTIDP4v87rYUJaCoSkUkTsRVSDgbH
EzOJaSpF+srhN+21PJO2p9eQgmdvYd1jws7keTJ4tFvEemjhK/DAHsfEuo+ofHw2
iD33M2c/8uadHHAVGGPcMldlqWFg8xkQ2g++VQLGj43K3NXaHNiaJgi8lwAEf3Yz
W1GFnaXNlf9bUt7E9cQfEE0nIbiDTfMWFTUNmmawWNY2NgD0C9KhVqqMM4qIu4xh
WIL74bNSWvsRRu1OgUGxMlGUkmlL02Mc/zSagN9V4pYabhKbmIQsty8exvb2i/Pt
dMdU7SasKTNLs5YN30U9KWMkGVCvmcKLs9E95tTkptwu+i5In7o5EFJSB2FrmCey
FhlY4SGB5pNmGWDdve+DTN0/V0LC3nvq5woR7JlgH8nrVUuMFPQlK22QXwmV0imM
24pIGqWgmvXIR1sRim1L1gpelHwBdF3RiErfe2xwvEeVhumufXLe7Mv1xTX6B0cn
EqKmavSbk3Dm449uzTv5ERbr2uPU27bFJG+0xK9U6Hr/BSAdhbbyAUwnp6hGqxY2
bDHBbDPp8cwJsI/myQ7nmDkUfIdGj0SOSVxShvGgBWD+nBITcJr6A6c9Wcsuinwv
Bbd/VtP6PcU71fp2JRwdtPKPAv+fwc6e9UWc5MIA4LZhQdQq6MOJo/u0s/5Siv2D
zRcWsLrC/B9tlqXgwZYOpxBnadAum6km9iXR5aU+ufg=
`protect END_PROTECTED
