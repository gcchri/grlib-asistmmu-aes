`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EeNMXHzbztLNYip4SBDeCEpk5Nqn09ZA1ncPa2mtLkqWkOoE7LEaB6qWw7+g4yxa
l6KErJkW1CMPixcEeQc7xdQ5tdx+wdURTZeyM2Qs2bARBYa8ClC2y+ldjxQqBXhH
RdZHLfPMs+H/+fGmoLfZn3+L64kQp5jfNj9NnGWD4yEe2OV7B7VUUMHyTd1U7mt0
V3SZDd+BE76t5p8JTiTNu7QVzplP1OeT/lr4yUBlXGA/k0sorztzNa0jH3y6kaMY
k/XDSSUAL/Fs4uccFIbsOjYCvnohkSrwnUmHJkGrbHeL8veSl4WQPgr424OKJfNY
tdRaQeV8Znxra1XkWXkVZ2lMFWjP9qRraxKsiOlUBxypqfjk2nYQUQ/85sCMMfs7
MLCpkmP9uwclt/SG3p5h1mi8HZxScVluYTjCSzzOHqp87EzYKwhdC9EP8zc4R8VT
yDoYtzR3NuXlR67VZvNqHGZOPBV0oiiYjvAQ70J810Z5dZnyt3BZAmeeEXRvNT4S
lN8icniZvQ0tN1Ovbb0FSsG1tezHqhn5S+8eLmqLhayu+uy3Gy8G91cPHu2/lKL3
+KmLh07JRWp7sg3Zs1qHjcqRJUbG6sTlzJqja6XWNFCdY1c8YNS9HvdDCr6ZUjon
hQKpklYm0ZFyEwkmqUPf6E8b3Mz9S3vW17H96uKGIpEB4gjGpYMz6ofXWc0YkFpR
c37ASnu3uJNzfvj6gw2I20BWww58PjXNnx43hSkB1a5UcMxM2oNlYEEjwBdhxr5G
2puGPeNkBkFQV367PH/EEB6d0rbadVpw6loLjvN9evyi1AQWPejU14zXu2K4mj4F
WImf5yRrm8XxwMWjpKociwrfJwxec0ZEiUQyqr5EATFp7TwqOSMOLVWah9hUxqOj
H6qlMZ2l90qbR+XJYpMJRnkONKCekFrFE6xkEQWYZ9TWmLnO50gXslUTmJZdLEGk
ozo9xBdBZYQobTaXWnZrflVFaZfUUbcnkfsDnXZplbN0oHetJnrggPtu3MhqkPTy
/FAqiH9gEYjUsbCyYkamE0SpROZgNP2N6pDnPO7J7EVCm/QiISyZkgSsSj+Qz0Oz
VQUJLEtIcn2O2lmGBgKmdp0jqhy0ycoBGL0RyEcO8qCQUzi7lFhY1CE0Rf59p0SB
DCJV1xyguuUP724Ts9xqLxB3VduHdD3wdlIDH6Zu9zrN9EyoU3kS74k+2d0o3P7E
zvLMSpO6Z0fh/SrnkMhE0ywIw24IOINr1CH+vJDgsBFrC2jG/oM253rOSrwp5+4m
/ckbTEgZwDte0UgxCe3WU3/gjy/GB3IAaVX2LiZ7C7SfBOQFQJLtdpxyMu2uM7Wl
efM+opje4MlzZX7EwGNV015ki76uTKFx5PseHopXZ89KsZyRcAosfhIVlnG2FG6E
HHvYnfuNXMKRsXRWh7MNkSkusCqYXAEQU/jlM/6igN/xkkodKA5k5ZfWaaiTO8as
8xTG/5iMFzfQ3HMi0vekS0GoAeco6NyQyRsRGrFXCeuHEEXqoAP8Qpp3iW7uxfsm
XX4ZM1XAouVpl0irKSU53nNYszsp7I7lBBtpSIKpKbXwayoZ5E/o3nR/QWNyLUyt
hAkIaiTIURwswTuHi4MIB4Vc0MObafGvUytFINGfjd8u6gyle6BOCIt/DGVSOlQR
DZWd+Fl+GHp3t6gP1vtisiG2C0RsDaHRRew5x18h35CGRSh7Upo+o792BFmRV6PJ
PdZoAMxl9+CkT3K7olhBaT1KfdgFPt5I8GzjuK8zKHSsYIDZcRVBjTcrV1+MT+Fs
mPSTnW0brBADp7uCX0IqeA8BgQG8pEK/37BXSiMUNiLgz0OQ8bZCrF1KYBO6q3or
OcnxEwd6S/ezsv0c2kJUtVG3waOJCRcePxcyqvmzZsgxAQ4dLqTJU4Bn0oP9UsHZ
jLfTx5961+qV47X48wM3y39QCQBN8mzkjLFMaX8nnn2U4OJMPExOcvL7FWysVJia
9SS6FTUF3eapizBIDdfSxlHLl+EEP9ZHm/KyH9j0ZPeZqnggl4QxjcBqbiUlY7P5
e52UbiIDlY7ropoGYal7Pj3CKAAdpZtp7cNMEVEwfYFXdncMrbom07A/T5VMblIT
BHOGiwI46A2gM1v7jozO8YkyVYpThgqQdQFNJorplaBb8Qi1jZFI93T2ptZwrd6Z
RVAt4mu1XpXSeG7GaCVFAg+RLBOwJjOOklnXgS9zbjKa05X62DijBTMARK3BoklP
avt0xpNyxAFWN+fSO02Ic4vMjwGzErn7GqW4b7usSKtj5snkmWZg44Qp83s50qHt
5YNg7keB7tnUyKTXMznL3B4BBtkyBNDcqgCpF1bVgy/zj6kc8z9kG0/hTbz5Sjkf
GohbiO2afUFqhIWuGGCcKGn5XUIOyE0JhHGw7QLOtirRvlkVUCdy8JFiUlgWU6Wn
Ua9JLsSfSF/oUnJTG5A/NrLhdTNvBnPh/oBQniSvdaXAKDdE2T0zbIb/PPtK2HH9
KzZM2DbvkQhiApr030QPH/8S7zWwXqQRmfnPV8gl6SGVXrJmc24AKTvpvO6um3HE
sVxyeaDbkc3vaNb8RgDRVXqJ0iFfeqJM/U8vwfnGtlCEg9qULc0512/V9wFXVoJG
op7srXun1CJHt4SKKe3iU4VPVHRiiY2wcgbfkhsUIVgxpp8NPK1FauM6k4XGXUw/
DpVc1gpK6PN9Nf1hvFYWIlr3Q6t6Ro2yYWse1LDOioxOuhag1y4mcAvaM4xyP4dY
YfHT92p9hi1e4uGV6zJBV4eKXH9EftvmPsc1LKblYpUpxa5G/Q9Ou9rMhztIWYzJ
kTNWdd0gCZwEzVmmogaFZcQg93zuk1/QiDzqcp9n9sJai7AdWJZeU+rCsyjSyhgJ
oIB4JylnvJokT1X/3Co47acCGweaFa2SLEnyOfLYGq0zPJtCMGS68a0Ri+YIUpOa
59SC5y5Ca+ygwdVyO9YIfMj5G9WBV9wW4GPAZGtQlw0hIHqj/SePdLJX4n0cm8NF
zGvzhfO5N7O1h5Z3TSWWZ5R9A3WevkWQOjq9HZtBcmuytz9UPnUX8iyYP9k00vH9
/9Ve20kM7yMyf9KvFF283Fl4sf6DFibAGECm5dDS+4Mpl0EWh31cKZYfsNiojYfe
2o9B9p5j23zfumI+Mtew2A+wIZdILLjDwhsCcskUJ3RXh6yJich9PTsaoMEKbStf
5xYsEDHbZATrM9taUAMfbzb4Vd4OhuAo3592H14ev9w5+QddFcwnJqwpBxgSZWav
53crMJ3exB6HDIZ3g1S3FR2QWdCZyZ5SXf15GacJcGaOLOLCbOtEH6g1wDgduQy0
OmB0XyvV3cnEjp99XP/pjbL4T0/2T/kxS/ulqz6VUoEtdRw4NSXhx6rUP3btWRbo
wTdAaMEDkhs2Dlm7wl3Cbqdivs/yrgV07TFbKYwvBHB0o3nP6NMn+UQ0/2tHZRXa
s35CnSYUzoGOANspADTN/5vn2jCUZn5Ti9eFqL5545DO+bN9TrfWuNZ/KbhrTZlB
JUwbfOJSvVkRC9YGnl+UgM9hXMJ5qWbuGRRA/NHAcfFhXrvVbSNwQPmwQ+xo3Uqo
GcZ1J5Og+2391QWIz+P2aFpaUHyterf8HQTSuuhmdxesYzwAsvUTvEO9Wgaixcdb
Lfo244rBFLlhAhQes404riGyQKdlfUdGPTS1HNsLpM/V04XJ73i7t0wq1NZq4hLF
YGOsRNC6Fu+lWnrti/r/t5midwA+ltPTJRgmp2RvonO+8VWJxYArkJj2MeIisgXm
mYyvcnaTGZfz+py5Eho8D+6Okn7ztNEhFh9cG59GgNpB3uNHXaOA84CJH8Pk1ZpO
6fXeC63BUfvCCZfIfUqQ6WhBdJjZuHk6PGcT7Ci73MC2zLIXRwpW/CkOlNlp0PPi
0LTXjGH40ZIrOWb4WAspi09BRm4o1Lg981ORPiyzluYrtCxY2rRv/SAVPScNBLXZ
vFwpyoEgyJGAXlLyUQR76Sgi/EVIi3fVrYGrA0T5sgNNaLFy9IeUw7YiE0ciP7TC
rATDS4X8EqePxisJ3jOb3b4sTa5Yv9O/lVoeH2SyROO4wBAH8g8Cl4dz2W+zKIxu
4/D/UGsjb2MZvfLhzav6pqrw1njsXiAkrDlr7KmqrrkX8LhWbnEDWoKuyMI40BAZ
52CL+YD3KDiE0TEeCDmoEdlO35FYO2q9AAylmwh3T7p2Fr/YQRD1VZblHrp7PwlW
eafekWeBvocRlf2isvsLIxzy1m3Sqvrr2uikzz5Oz7C51VtM+GQeTwCQOBNvKPP5
Kb6Jr2ZMymI8zNdiLbx/wm4TFs6Q5zf+QA0jPg90dDPrt1LU7ZMn/F0radCkyIRb
JTEuDHo2LWuPp/NfD20lHTOhIj9XDjEgFt6OgkepwuO1DDNPfHWXo0m8XaiauMPj
n53sVI1OCwgSlVKYr+c+v3NzKvfeH79ewGePJSVbPHAj3RE0SNWygFj6ALZBtaDo
K6W4Z+PMkTte52YGqcbrz5nJ6EjOHgsT/xX4DNT9uBvt5pq2kXc5d5VEj84rQ/rt
P3L4hxV8bBbhBn04TsQiV7mRNhw3D3YmWmkFZXDrgpnsWPiYOotX7w+rhh93zgKD
ubc77SPlroPTlNupXS6joFy0m1fFOQ8PxdXmRvjeR6gmNRSFoN+VZQH9/4FIYatw
bT0rw/c6GNzr4fCqRzPWII6+tR9cjXL1j84yOZeLQMWfj0AWV5yKipD2hQiJNEWr
UBV3GC6FSTRmBmgn+sIPs0p7xF7M0h225lUAQCg8tqEDPyb979DcOWLX96Cj5Rv/
gtSqBiRZpSsTMCBM3YrbNPWmFJgwIJV7EHGFlefn6hrjPOBXxEi1jeEsi9aG1LHw
TedMNxI4+4fZbFVuWWrO25iyKwuzUfsrzQJSggldfxXR+HhRyb/aRMlbE2864ClF
tfcONsUsjMJ/3Vl/ZSc7ROGoHq9fNOTJy2dUmGQc9gyHR4IDz/ffBVYsq3wvv9xt
LFs4rES6eNB6jck3OrP/nmS7BTIkVPG4v6gRRWCI+xe4DhffYefOaJFsgmpNNyqT
1jDeJpl9n5KIiL07n5mb4AH8HXSTlZjCuakaDKA1gRwyZBERx+B+0k5u2tRacMCr
ooWc8FTntizYHwWWXlh/i+q0k6xnUIm0XibIIQ0Fi+/OGDWysgXjJLRBA3FEJzss
4rZZnVe97wXv3bSY3kFqepBhhH0Fa3Pg8WwFrxUoxLlJTDlw6ohBN6wsMpCDgB6O
wdB93gl+9BhT/dV5gJsaDPsVP1swKfpz8wwFFVJO4iWWd4PzMidho8p1r0E/DGuP
CuDBaXs3IzcFRLznuzoCywDPMKwpyNuaA38AukTwf97qc8D96t9bYG2yc1PYUT/h
h3AVWdMoH1135WTP8MTkB8eYbA7d2vBRvLxijT8Q1N0YhwbRHa8ocgCZMAXeLewq
43gAZ6ERdJs+baCsjv5fDr+nWJ8qVMt3EjRuqGb0OQHwPpRN/DxeJoGm9hIjd3ih
Ef2SIOf6mvEhropldWhocolwTbQV5E9JFbV8gqXecvhKBIkth6+6UbKppYTzcz/C
gS0M+n9ly2bM/tPNT/YiiW3ewIEWsqeXxuAyEJr6S+U445WbxJTY3zv8+4r/pkiK
vk4tXFfTebPt1r6U1ReShmchc9KvjEI+Q540iw6pSYINhXETM3DWniUlBvfsDGpI
md1i9SUZe9c69LnFqWLuwy8oWPVq9rqK0ScKfg3uWqUv5uOdx7zE8jZHxpc8nkVA
FtIJ3InoVjhIdki0HTQgTzcFo7Yxep3TKosN8FapijY7RzXpIXuDGfwd951GJsug
KqAzZTzdldcVPw0zwO3JgFlZe2BxT9Ukf/OuiGoBjWxeozyCdwTh+jmZkWZTsvV9
3Ulvsmtg9ELgwbTAWhzKEJGP6vNTCZda6JOvjjVe2FnNzmNofofD+3jsqF/Fo5UE
/G+yWXi0ZMDz28CZab7SL+K6IgnrkXu3Yp17xJgRgfvqUoAJ0WipxZ5Ci7/tSmA9
qQ9KQXJsNNPNVaYeUmWasYMs43Ar+qEqivg2dHSsP4L6Zf8p6IdUv2yjNZ0sufWq
eLVfdIfPgeLdcK2bbWmLt9ZeMDD5XvqPgCojnsEipa9KfnJWHfz1G1RfUH/J1r1U
J2MT4BuLOZoCyOOrW83IMjNwNjnV3gGj1vhpqxjGAOt7anfOavSIBkJi6ma15njj
t4U3b0SXr8fN2txSN9Qqyzp5Pj72sqkraw+DgpD4ZjmSana7bo/BdknejPY5Tcof
HYO3QmXnpY33t7eKoRjrvAOqqMjqI+OQSDGKu0QkqYcB3lpdftzMwmVPFMjTXoy7
zcZglhWS57bNcTD/ImCFfTzbzb51jOcHiigsFCuv7QvUZVImPDxdtAwPyJRyuEqf
uq2hVz2mJXBeu65zH4vYfqAxlMqni0DdGPaYXt5CLMKVB4q3fTfRhjspnmNnjjcB
osqsB4nTSRItty1k1DBKDhgAvaFOI2dplUnlw0k47M602+JbWFNkjpl+QFa87fDy
cw7HINeVvxxEYJj0l5qY2IruAELx+HOcnKJBccJdLWqN1kKKnKZc3UpfTXrme3AT
M5kdKNigNZrnBC2fABhXD0rdRUWGEfBEa4Ln2DD3uCJlwwEvi8We0DfmxfUeKXoH
Q6yVLJd/6jnPGDibMJyDaFiYHl3SiKxmoTb53Tqr2I/FKOBOsz/X4Cpct/oYpikS
jcPT1lg2CW3bdh4BUhV369Ho1Qk6N6OKiZQlmPTxTnwOO8Z8Prx7YYR2U21DSeBT
3ooIi2oUVqRPzlt93R3XgVVeKgndO26uw8SSO/3HRvt3L2kKi6VL5mK5lgtsd/hF
d4n4n+aIMdlvvLJSTIUaQTHkRpTwjkSKPDae3CBUHqztUTF8XfrIiXGBYAoMbwdC
aNGhbUkdFWxogF3RsUO98AZ7dbGnSMdFPyx6Q/5i7dBWgXE9+8skXRDsBk8pKozA
eIkiSOr/NWrmO5xRx9iVV6R2ziLjn+RgzIoKKTCy210TaqpG2isX7wmMsjgEXdVp
n8ATQBbJqcVwLoc8pOGZJG4QSuVCLOyRVWfqTRYORrRgZx2XJDsPdRbCt3QQvhQX
6hqr4f03+qvCtvGqVnNYQXalcJptybSYM5noAVPpnONY9Tyz/KDAoomKyDqwHRri
g8Td+4xh0Vq3/H5TLrM1tAAkP6hYhaAW96IdqMhLqObWeF1gimkVIc52t8aBy7BI
t8UW2+LImTTGfUoh0V77cmeGrJc9NO+N9f4Pi92PvEPKZFq9DZtWOUnGIhz4yi4E
ZxIgZYnYw+FneC6mv+RPyBvd8q6c2J6HEHd09MdC6cQtp8kWQtwObpm9bup+zpGT
NYHWVFaN7FkRBn4TZsR76K3P+mBhiWM7Qrs9sq2kvGjqIynLOXzdkYtL5IfT1vsa
dFsvQMRaCs+WFetspJcKQQfkVwK0uTUBtK7miOsSE7Mw6FXkBzR554HxEokNhddh
zIBMp7qpon1KivQ3TAU7p1hBmeWONu8wfqnlW8KhymOgeYL+YNRSLHaMIfNAapI7
Hot+DUPRxCfLOaFwFCvKN7zbnwPgE9hHj0S2dgiGkS0zr3XgLtNT44S8KOUe1cBG
VkgT34TAAEyc8EhrNViBQy0RGkNL7dfABsIze2yTJn4kTfgL2wkytqle9/tYeCIL
P8Mhb1ULjip5bM2GCPnbjjjlUu41nEqsj1J1YqaqbzYhTn9RmCmLEMHSRY1tjMM4
iCVHcVLWTF/QPNfeTIlMzZ4cgVdGrj/Q5h9XJtzrE4fB24GjpjBoPiDlvx+WltdL
9RjrGHizEMS/8H1nAkxtihxE98ltmtyk0nXVEu9qzb7guDJqJNS+dZ/0JM8ZDkn6
afIGuEtHPJKzmiz+v+Vl7rWuGyUXLxic0SZDMR1Gcw1nt/2f0+zNfTnJkQic6jti
d5LGCwEzO0lH1Y0qw72R4D7thNhrBAq0ntOtrInFch1aZkoFl6a9bp/4sdE/kstG
VzKYOPnT/Wir4GXHXxHw3Jpf3C3wBpGDo3Qh2jsYL2UFeWxnhrjXntubQqqE+xaP
/v6Jb7RH7LlwJER0TFBSAGWThuiW6JvOMJ/f6NAmvLoYCC9In5rdDGMKNeU+5dmX
YSKTsRhnM2hQj6IBTtMLnSTLjzIPNHT2cmjwJmFDBUedPzsBQkyRc8j7zYLi2SHL
rX/cohRkCFU4GtI3d/5exiTbWaczuYGXeDTaENUE9hgU+cWGQO80MEJYYFdW76hz
1ChRRh8yLgpnGOGPMdqN3y1gwd4twCFlbIJ/KY+Rnq+r0jXx0+5HL2ZEkKpMKshg
ttLsSkJ+aKYlHxJrTQ8Hv5t2N+/PZB5a6vLtp+iTGGUFVgY2q0nGTaQEWqxgLSYI
MSautEAWTDfVZCR1Ywo16atrcApes2+LfuxKeg/VFQScRCOikTrNYiTMMeHY14WO
6djR5rWxWQvYnSIMgHdQxrOKcMNNCKkYNdvCqLU3HoGHQL1pTXzkTlUfy1SZcO6e
GAgPud0Q31iK9ku+OlB5GsdmxpZj7CTGuCOM1AJF1uFXcVpTzPy4iWVghPM9y6V7
1Z6V1jBSGj+iQby1lQusnXPgQJIEwm1dSaO47VpXqQDMXvDHwGqlsvS3B4tNZ7iG
1CpJLXKrTWxAY54VNGvqtRJG6CnPTHW1J3j8Hxy0HVHoYjRz0jqGu7+OWwt1BpnW
Q6sP1cJChnzGA5yRYH2+c6v7GvyusCDvV8KqHXM6mZrvY16TtbXnQ3M4IgjhXpro
3Ls1xzcSDeAK0yxZTuAqQfiHTxtNDXQCOifTsQC2E3F3LOXOo+EjSspGJxDPPPs8
EPldVKb3Eeq74gbnN5T6UICDBfSdDJVZt1x02VGY3XLS1udbA+rIf0wmuOKcE1Jq
Yh5T1MZbLcCc8ItrZQGUBADeeMKFFUdDmLqd5iGyjomXYUiYz6J2pabuq4r1QW0B
MTbj1rwTrHf1VpSSFugdlSVuH7Pnyo6jGM+yPREH+MoOnP1bAbfx4HVW/OhPRyl3
X6vMpL/24loLsIbsLbcWCvf/escUbpuFm4mmbG2WC1roPM9kN5QOhBEu5874nEQY
wuzhfo577oJtXeV+PP63hUgF4shFL2ZpFiE7FMZjtkNUu3iI3LV0FuHAvp0HK2IS
KjM40A2w7NmfUDxWYLDc1bX7V+fImJOilruKtjc4KqJSfa0vG4baJOps+KUme0/i
Bgf6HRmZ//hejQIqNIpYW4/c+5u6qS67j72/2otePx0ksTbQ6XeVx8k9NKx+PImE
S1xEDviNVR04jpGQVIOlgIEt5wpcVjBDDdMZcdiyARu7CKg7kEt/jgiRWAGOxjp8
YrGSUFV0V8WXasTvX5oofXxw8DBlBvBMrsMsNkHz19cEu8tX1Gjgv/cMFCfIBL0q
DbQvVRLhbvoCjAmBjBCQWR3a7QZSszOdag19pX+PkMfkDtzEge3FI61bGgo43xxb
0U9TJYWMadJK472n8zO09zpMQbH4VaSpCjCowdZAbZmkAePtMFwmgHW3IV5zsWeW
9ApII1l4gXsIrcWD6paRaBk92sRJQrtJ//Y4IYy24jF9BY9Hk8Y4h+kP0/LNghTb
wdUm2HC8EXOSnr1zbcOU9890dUx/YDXOTY9YDe003lYROtJjrYUHaE8RbjBVnXq4
NDQQeufCDmkTG//RtmT+VaD9FXjKlvNtCUhIL4IYvmjw0LOlBXAKjxy1HPHq7FVH
rS5zJ0lbFq/i/hj4xHhHZSHEJwfMrpQUMqcBD9InihPdgpyR/F1M9HTd3oEsEI7C
2sOtVkgX/T4nHJukwqXAWMIInUfsB6HRg0kSDu5lbsO/I8MMbgjG3s6Mfn5zVmKE
YcRvzYgbFzLhw+y6mRef044Nyz41OfUUkmWxq8xDZpCQc3GaWeYEMI1AVTUmBJYq
xtIwu++YBPWI2qbWQLSkCPp1hqMp2cXM504zU0ZnfZwfMDpNNjbqDrdZAm3qoVJj
aLDJnYLmVdbU3OeDTH81FssrROFXLjhB6w8pPUVrVeTtKxtRTrTEuHazXK8Bequ1
HbtglArne7CXN0nfRuS38l0Po76ezlAYiPDbpm2b8muc/Vanvv24jHDgBY1+jLdW
5rMoEbhfrN5iY4mpca4AKNDc/X+e4dfSKlYAEnEQVxj8+3gzIdV3cRydlS5q8jcM
UD51zJX6J3CHzA/x6cZ5+OoQ+wr1gwmrDWapqCXtDPrTaefjn0twNaqanzKFR8DW
M4NfVOzGtJpaMq/AYKOhvpdYG27nHlPg7TdsWLCxMl31FEYbirQ0qQ01rJkxN24Z
rgfJ0tWPlY062EEKNzBxzHRdCoTW75fSHmIE/e/aKCpBYsBF+LCJ9ZBNUfhsMfqd
Njo1Y4UMoo1ars86wGvXqziWz4pzqiS8vCbVm5yBhzMtSPimkpgqndIgrLn1Aq/x
gqHPdbV89wLIXvZP8R3iw7IyZ3PYDVyEXrxWvX+mZPBAzxCTLeIhzLhbplEmLAgI
fZ8nX5NYiXbajQB9awetTagJU4daJ1DgMZg2FJbiBpunvz/Gf4+gY4I9Ds8ww9JP
9RcwkVQJUa0XBEQZ2Lf8+wtBxr4GmaykrDvHFF6BXZ3Wouuwq+exdLGB4AuFHVoF
az2eQIJmuDi/8xzvcpPgk1zcYvjotAnsu3w1FOrxcms5xOjf3vrnlL08H7s2zP/Z
9FqcJof3x4FMsalGKKcupKbmXrIY60Jt3L4bczy00JMCKNxxoWBw5GPqOrXYbuV/
RQ2t+wlkcHqCsrWOg4MSgGI92MGQc5XFZtk8+1wCXlz+3TDirIC6gKEk+kBtvmEX
qIpLP0yvn4ZXDj5JL3dx8E3WG9a3LhEiUUTVXd52u9aGDWpuAuw1DlSBVUB8qns2
1ZZD3gltir4VKK/lOnCFjv04eZLWaKqdIKICgqgoujoSu11W73uO/e6EgBx2UJ8M
8Yy95xq+6HrcUJH6kW6whmndwU2sBrzilVXGH6Gs5lFzNOIOiaSKW7mBvT4+O7Cf
rze3JAA7sQBjNfZ25LLHWOE5HcLCctK43Cd7J5XpTUZmWKthK1bxXLITLVcPBSpi
RG9w1HQzvsJWfwp6d6BANYYuRX/VpurVOkGuTlC25YfQMru6X9fzyvHZnbSl4SKc
q56N729yyWykojwluqbBElEq0i7gmrmIb+SR3g9dQTV9W4WYP3PbllW0YJLAVozV
KQ71/Gl9FsqGI37H4+JPkWyZRcqxoqAOhDvN4haUs38ivo46kHySd53sGpNcsZ/1
mw1Mbz5PApzJk0r5X9eBgEbgj1tgVU76MKmIOVhdoanlJj4ubIKKhGzUSVk+M18w
JSN0EHuc3mrZ49Bwz7qm0QEp56JDtw97IjwVUI4pnr9TLux7Q03mfzR4vcbNeJN1
rSleBu12e+uUtemSMFBILLLXriwfD/jo2UYi1EWnrf1CovHU1ougGFpjj7FwKv+b
UE93yYZllP4YWPjAJ+tXJ73ZUqp3EZ13+8oqqQQw0SWNF0loIbXNjdHZfDH8dK1w
dovbvzFRcNHWAo0EOqPaaCR0ttrPtTehUGz1UqMd+fQOskoRlWGT8BHKrB4ryeow
kruYNskUJQHmBTlhzTo/J/dR2HhxzOgDiOpfQpp1IgGQPgAF/iORxX2ZmUPXsdl1
EsJaYOa4N7gr+uF6FORMCSCazyrcsapRHjoR5ZzEcWiwuqX0MLusaNUUPRYlFSOv
d/gM2cu2X7ngfFirHAmxrsXtfMFJokR7Bs+FsmjvLWyb46kUnXGRusXD46UkH5Pr
5LE6Tb+BwvcQNO5sKXG+VMts4z6vCCTCBaPjNzq5touh1W0G66EFapl8xg3xQbmz
0BDchBJRrwuGCPF5YC268o4rjqhJiJ7yOA8UCZmfN4cBZcx725MTY7zwyozvZko0
sQcwV5uHiwXAbygiIm6ytAROLlH0t0OerLEGREMMgEQ/Pm7l+8rLbvF3W2YB7au8
5OAZZoXzs1C06ZlK3xTsPt6ylK3uMFiWcWejD/awRl/eiNorfXl8+ot2jMBNdxxZ
2otgsCiWbpA1tjdUVxnZY8Glc36lpTuZIoyUBnHzZTJ0936tZ0zX4F/ttvteTbpT
81aVWauZgncsus9NHMsF8K+rGA1kjxBAI97QGMKs2BGk4Og9hmM7PCxbj4kVBmlU
xiSFx2ReiaKpxiVgfVY18HmqZ47iEReBPkX+I0FYsqSJTgxrn8azPxyNEBD7YV10
qh08jVGAL4NTr5S08Jyb59Vyk1KNT1GprG+Usmdv9+1TtFzJ2oo+xHbAo61ecMtl
k5FRuuFLw+9cWRWag8BW4blb9LRl4Rrb4KLhoXCv0OpqmgEhnMiOAsmWmCeDNfjJ
BOi0LbtGLi+r6h+KaXmi/p6TblMzzVYIzLovEztgxe7HU/wA2Mbvo5a4Rp1DZBtc
pGIO+rIb9PsMvtWMJSRaVKP9uaOotykcGJy62xfSYfU+JPJ5XPKwrybS2vbuwrMM
i+b0WTOWVSlyf2fb+3dq9ZxeaCpgdD5zqkJZw5Gr22iIXZlIg6FGUI32LNgavbth
pHET46hp5uT7oaVDZutuvwfvR3H+mh9bHHmS1CwQWpifTVkj43hdthESr4Qt8nIU
MNBSXMxI6RRyWofSx7gCtIeUoYLBQv+VVJ24PAi1nxz+GzojSmzGLeJDfet0awRK
kYMbZTI0DmBDQqdjO4/VW8KOk9bTg34G5DVjNcEoTuSkEI5C/W2LK3Y6SWqhx/JT
e8Gjk4qK0qz4KD8ZxChrlfqQorHHHkUBh9HfKzs77P+h0TkUBhobxyTYqx+ftXUE
HyW4fq/BSbPc0sxiXIPHz0cJu9ujp2zrak2yOYYnVCtQfZE98Zck6jKkCLMSyPab
4ACJABbQfI2O0ntPopjO3phwE5K+YvMbn7MgGSGzE6xNd4P7VWajniZ5UlRQUzLy
D3rohV1EOoXfufL48g21LWGbEKonyX1bHLsymufuePHwQppCCrV7nqAZJX+UPM8V
fef6zPi/yelFFEhYXXuiIA56pMX5fPn22zzzeIGI0TvEv1SdJPkWmJphz7uNN6si
YQaRXan9ESbThmz2WyH4Q0RLenlfse9ZjxVtIlAT3frAUk8bmduMVZGMayhqKWzQ
r9BX0AgQw7LutA9lFGnanqZMtTLvYs7VMh241XUz9liB88G7t3Zo8eCkGHZUoRtS
DSObqZTrRRZKE2vK/2dLaqhCFUH18Jn6gojZTBFLq3tQ04asPrHcm+HeGM00/szN
c4BDpwYG52gsf7DSXyWNq3LkMPloBKnTWMLJMeWGPnh+3CEVYSePl9A86yns6+rA
LCrYlG6o/PQPw5P+0JILnEOjw1VMHgtK6Cur67YNWY6rELrLntfnCAE74hLnVMQb
Vr8Q6SuJFI8PWJH1FfY9ifg7/gMVnBnh0/dI5d76cTsVx1BgE7OC9DjcNzJL9ICi
zUdghc8s0rTR1BbQGyzKxLdkwadbcS7ogDeEWEuYzR7CWWUGOBL4vfqlxVWav1QA
npYKvMbjvfUcfLSByASS7ySVGHJHbYfFYgmFNMS3lNSersxdkxj9lxETtThMPj4S
2CaCBGi8WEcsg58HezOdpv3RMqQBzqHg8kX6kUL0/GZJHjA/WlDaA47bZXC8Grs3
6FdolkG2Oc85kAtqzLX3lR9WDcOKRdh2p9HURd8wZC30IDfxEN0eNEEDat+noNgh
K56+eZj/zj7UMuHpdy0uZa/CZLIh44RRAMZkYp1YNZNbNZbBdT1TsqAgMfm+gJEp
wFbBmm7MxoX6xYNFCcvuDa/nryIRdQ56rk08WiNk8aLRz5IQDvHrjDoo/EduFX7Z
qJvF6bToKRGNeXsMNEmj0aswm9XkTq0FTddh5sWklr4/D0TQCaJ/vmhEqqxAaq7+
nCVO0bdz2S9g3T41pQXjtuLX0p6I0giXfLGyflRovZ//MXcUEiTefk5KVneadBq/
lzVieZ+Ap+ZmHu0dlfbJEYWsictgFVlQvYxTINzEp1A5jjKwd8MWQ258Hxg7PI3L
8O5QJAmg7eIyY/dNhSQtmTMHLbyT47oxxnFQuj7zpTUFLbas/o0tTdAg7EOyYQFK
gAmscsWgZ6czM2tGdQgl/hPKvFlXJeuzsGt0zAgUtmhoc37uulm/bZo2xIadi4sn
5wbf3151TvZj5KNacSeDuF8o9R9GQCXz6U9jZebfAP5CUaspzEHTmRjo1c27gWjH
IQvtdGS2Nv4LFSGycCsbFjAw+DP81nF4olOoaTh3L8w3ui9tm5yMJjurg0vTtXoX
pxrZTcZjAutcIdaGwKbkWXBUVcVhVOYZsCoTFq3CH4OCSjPDj0KIdklYtdfGriu8
/6X57Tb6iOVuK9u3xLpGZD9ze6ceVF+1WWUWks3lDc+2uDP/FQqO7O2bC16P6E7s
/9oX7E3bt6uET6XPbnmrjgJki50dv+ZxDF5/zzLQHLpvCz/qjTbo87mId48vqtOL
ppS3z60t3ljx6vlu0pYBnLFul8YkRE8VLVGpCQADG/713IidafbDCI2rPoYAngrp
tO0NJ90VFwFUSzZATnHuCRIo7PRiCMm5QgtOojywDGMFryxcLKLderpMx1ysCc27
4/eByX3d9R/Q6BVtZ1SbZcr3ljnQzLpRyGQjKoSUXjM5gpoSOgNg51EUbe2SjzmU
h5O0t9PnGOU93VnaOOvZN5fpinPkMrdQ8/SVmsK9FrlAeTys3JSMFGPR/NpupnD8
gZcWrWvxWEaLAHOElC4C9qcN7bx0SuhuSlA1FdEBqMmaI+cVRzOg1epmcflcz74a
pxY1vhfnlkpCQ/SM/DGCL+78mu9sTAjZsD9ikLzyLQv+rqrReBp1IrgVnRzljwI4
0SVYZt53PtFedRIM6euoKO2lH0oY/O+v1MA9P6vUMWm6TXr4ZOjvCczkD9+KtHSi
fDkRFs+iqinL5efTwFCP3oYA8kXOggKNvNosnfXS7772Z4GJZy03MqmXUZgL99oP
yWMuXZsmfY10jwZAROOxZN3Cjx4+YKDY/dneCWPMqca5e5FKiI7s3KJ1Dg9iwaT3
DwEla/vBmb2pfekfAl0+Q6wyDp8qqMgPQvujEw6fqRea7DNG1nSYFhoqcGggSEW4
gR3/9dco/yTXAFlxA/nbkvRSZf8yAMVP5i6wwCbKEHpJfPtVXRD4+1i2szCWGiYn
4DgbNiiBhJ/AXvcQH3kFDmL0taxsQBheMaEaQfZ9nHyQBacUyhh3LDn3qsX7W1BG
jtFIgHquFo1MzjMpoQPWuaJuozNPkPyEUVqRLsJ45gJ+TpiulxPFeEm5cPxH2AEn
PVnGZFddv29gNTh5Z8EWb1ZKS2MVxulXq3RiXTk3+Nwwo47RSvjdnv8DZ+4DooE8
oWyQ4w4LS+SICFQNMJHfPePxShFoz56DcCyBPzYHgz6oDjkVOaYffj1BiiLITWtW
2RsebW2Dz5cBv3QMkt/wNgKB/mebYJTiDVlPhUTXdW9Eib1LqSRZYbC81/RXPmpl
RotSv828ybruQdPiCakPGM7QXsYnrv55JCnL0/NHYYkrBtUdzqAIr/Nw0PF2ODwr
wZ1xFctLcktk/ttUPT/zO5mOQq1eEyXbMdndOoSgKNc9jIOGDqDw9iOOWqP57qD0
bosOWMDa38BVvp36wmm+WM+kECKNQKViMsMnbCDl9KzWlT1180GtEg9eC/gWF3oW
gn1RHov8kDc6g8NseE+FUr4+zlb31W2X/EDn4NG1xaVRyIvrukYMLQzqQae34dfJ
3vnV8vRXqTPkJk+tshQK9fZD46oE5AD5AglwZLBJG9KhKczTwm8sgftilIuF2Ycn
qK62mFAivXpuEMCiS6LGD6WbTahe/I7L8krQLiORCBQGGczOHt8ocrdJV87KxZ03
ERz1YvgHqAeTS+seolwnGzVcF9zDTiW0ldZbH7zb/G9f/JdhzR1i6zgJ+Cyms8S3
0fYMHQkTMxOXFFsjTd+ZIbIO0F3r5mC/HBe0llxg1UeGrdRszcphbFCnOB5kvKtw
s9pZtXRZmlob1ltbdRmOItuuvm9JBWiWcuvtmb30/BzJKIKybJewHEYlEIhxTtvp
CrmRm0GW/f8Rq3Q6QeSTlgMg/lkEG7KssX/hswCh8veHGk2aP4Oa3UAMOcIEZ7+f
M+k3VfLtLzuBHPY9PSaLSRSEj2aZzC0ApoMpe2zGGzekd1uRyaTVPfTKtI44+IjF
qVSKgEBmPa7LuxnzdG5FnG1bvSlbgMNB/SQzJhHmjgRgMCUxwkQPtwMrzywa15Id
i2jyRxKYa+xWfw8DQZjoLtrlfqGnV5T0wK/3X+NXTqEMKzAwzX2rokyqwaoDAUvz
FFFfdNsErf3+M4+e0NhO7n8UFKU8d82/BH7QoMtHD2P67DnEkH5+mdBkMlfq7wuS
sBfAocB5D55ANOoUxWG05nk9kB1HhJIsDlL2pSAB0POJSZBBN3MfyFLVl8v7n35A
9ntylmIP/ccnEi/gzrcVO90mQmYLgjJv5kMSKKsxOEaS4FBj9PLQVUl09Eu5Bjpk
GIV66xOOWIJgOapaiwHua13GIBfwWWKqub1SxQqUn2YawY6xz6rXuYsa9fwAQn8B
crihdp157ltAhWAxc3ETZLTI/TgDiz4Z0lmH5LSpGZ7Iy5IRYNu2oMkxSl0sE4pq
OuNFzONQtYOk9NQFkvTzn/TT8ZP2hKYEondT5f/6WdO7oXBWbraMxNZM+82mb76h
lfj7jYKocGYyDgYyNF4VFboNGQul+7k1ZaufHazsrq8i5e8LJcgEAxYWTtiRsWIG
aepwxSG0XKUjfV5zb8QOD562vK0lbItsUx80OytgNicPuAtMPayIGisuida7p8vS
kVeclTRbvDtQgE/1hTGF570adTsl3XnmMMjCzqaaIf578VNkgLPt3vZEuLnoWwyv
0PWqjpFToAYyCxSeb7sbEiZl2Tad0698W1IAQzWTiWmQ8rVeaUEtvLBPGiFqcM8s
TKD7xap/FYYBhD3HY4Vyo34iqy1ZUbkkK7gY7dsE8En26YxrieLAwwxrtUTN/lYx
r9Dl4f8l8ET6Vqse6XXZJQSgt+Jyc4paA/BZcUEYORGouzKbojsIaeVZ65gqglTG
xQ6MJxFdCUhskaWKjtuYra007oN1OmC2pvmvN3WDeNOYLfUgbGDXCh19OfY23fVJ
hap2KNPqOHGCBzdrvsHu29hk6F1HqEnw6hqj9RHVnFrf9zmWzFPRiU4FKk0ehSKN
DdLQ+fRn9FX9iLCsb4pYbgvI6lcpfTEOI/XLmVmuIbltp/HMPt/RG1l4Vcr2PkZb
FQdIQ399r3I9L51p9aN2xuT/57UcdpuDtoYukGhfz6ofhbFCt+Ocon7Sq+bhXeqS
vvI56KbKxWOKI5bvaUGrkM4MXBPaMfBPmma2uUAo975OYc8AVVE6zxrlEcuVQ38u
shf+m0uYjaV+G/I+OsZzRMGKyalPg55a1+36r9LLpOZNIp+ooiv2W9rhfxJtGWCR
GIT0AyK+sCl5DlDWz9KqkjuXQgmcEcuMfrA1WRWRqycZ8pLAoAXvKqGlDWV8E1Ne
O8JQiEUz2mhrsdBiz2US5TS2vLAnU680grz2iGns2QZZt0//MZHZWO0Zf9kjHJLX
8cgHUngZEx8JbfvvZSVCeOJccs0GNdmv8IvttEY4y4Fb4Odh1sCIxQKJQ1CoCdJL
XJEnaMAPNLMYbachCdmnbxcNc7omwHZ/Qkp1EczGq6uE1u87N+IadP+x570oDzK+
gvme2ePXwD49fQ0HJyeKWP4zxWfJ7elQg/CYx9l0UqWcAFdiMhBTXBpbX620dyVl
97ImQODi2yZHVanvRKDWy6zkzj6ehj0R6wP8mCdzY7705b4RlC/tfFk2wof9dYEm
9vtawz8Ed1DiqDZlhRab/YOVtmozW5MXgpGuZ0Osaf74YkM/0tpByxI+G23c8UtZ
MVXZ0vlK7XLME95NpdxhKbuWpkYxA4uFUucSCvmbHh03xr3UorotuuGbucHEOd8f
kWGWI9I8Z1lTLKVHNI9nM24lMhLQUQwdDvLb0q23lBth7fL6S7WTTmIA/Wmp+3Y1
eq5ohLDnbDWjI4aiksPmlLzh9ArrGZ/6b6MGrJ1kSGyomeBJC5uuMYm8C5fAivGB
UTdq9w0MZvwbszU1JgyefyiyABoD6fIvjEGadMKrsiFLdRboiXXhPQTU9l741z32
o9PVavVQwSBL5oL0UhbJECPoUE97zoQ2f6L6Z5CXUAtvFBL4v+y/oyB33vknfeZM
XymXdxw+6K0uef3dxhrzOau9PgIR5NelZyUHzvqRG/cDbL9bViu0oLTN/5HcfH0K
Zxj7HPId1zEKw7B78WRMdlwOYY9ExgzGRTY3MYV4cP/7FcbUdvAfXZpHIR9yWxJD
YzGf5otDgio/SaTpcRHcrkb26xZtN/fav9H/In2V10HQ7YnglH0RNg6AuSlfF/+4
HbGkAmKN/r3n2UGAyNG6re/dhCZac9bnCJPfu5PTpANqKob/Hno3EYdCuRFVE8W/
IZk35tKSp3j4sS3cdsZ1HHm7ddfNEphWYFncMesf0B4kj4V3cUO8jVdlEKjkboTy
5vfxWi6keU8c6V8i/XXeW/4b/aludcR7zUm57PYRAWl321lmS2UJsMQ8HriGHGvX
vuInNKwbu3O8g3yj+WdiE6O9y8LsfdVE4zWp/fI8m5pnV/IzQcorCxMEbDU7K0Lz
VmwIyaFJHjfTs9h9501jkhGkLPR4ca4pa75R3H/97OTtjdqNB1qq5xCr1/enq0zh
g+Vmvv6c4PAMLoYQpxJHi4pqWFHA6MJYpY37cfO6glilsMbpDogO3RyjFTBLD23f
jRLdhGF7i/VGNWgYitueFD8oLI/acJOjNJ5+A3G0l1vjgPPjYIjIIPt3zdrkTRq8
dAb7YhvF65/ywJCmt+L1tjCd8hV6RodFdqxXieLv/tPGFGeXOEn4WK4lYwH4X6H/
8r3Q3qSmrmFOBOXBwde7lgAPRa+0WtweuegsmG+5+2BinpoNTiKdeGCzS3Fr60ad
5PLLwmv9iqhdi69VfBMz5lXkq7towccR3JKl7wWZ16CEgLrECXoUC+ygc18M+zYQ
w6vFYB07wU45FR2st4XaRtPqCCk6i4IL+AIU3arNLplL07kJ4ii6jEg+YR2RiXww
97nHSXTYGgl0Zxf6vdJufzD/koxQZ2yc3GGRm+sxZx9uhaMcVdAWl21cZY/UZMr7
610n5th8/UJFwuoj4GVr23TSamFPiHnzZwbbgKl6kn3NTlrA2zPadF++pypu2vQg
fDRrEDl95nSP2fM9toNj3p4zefE4wLwkJF+VAUH0I+okm2sJGdWNLyZ0Rj28UlKv
wAUHV1EdLAQHZjuPRJ/BLjclPZo2fUwRZ5Zqm8x/Iy26dcdlRfE6T58NMjhkQP8T
0bbQFHkMcx70zaMKeClm4rqaa9IrnjF8oL7SfFBvBZvEaMQ9+SNcl9gBpMg8vhFY
bHZXYIQjjO+PtaLFncQkX7ApfD4D4EOerjmf5v5LKBZsceHLq8TVPejFDFk18acf
moK9PRU2wt3ZNqxRXit5r246bBFW51Jyt1nEOi0bosbqE/ooWbLBDxA06tNffERE
h6FIlxJZz+JRNeXMuzZrDzh+in5Sk3w0ERUPRMYNXGPtwgmPuAlrl96VdHmIxY8l
eYxFPcAm0oxuvB1VY0MbnHjeuUnYQIGFQl1pTme0yBXJf0OhXVE+wOz2G5GdB0Km
Vmv9+NrZ3bBWe89R87TaU+nfF7vJklwNQEbYDvhYNBg3e5PvwJ45n1I9dY9RgyyY
lMW1kvKYYz0SB5PAMhBMW/ctJ6GcQC0qWgGYTp2fSJivTaCXazG88ivSkXZ014Nq
zzt47i6J5LMuAYDclwG8H6woDsCdAlx6sCi1h1fQ19Stt0La4rZ5KDZoOizhL2YO
loLSKfUpb3DSshIOzsdtJArjMaQ/OfxyuunMTUpVY5dhn3mp3/WaeF3df01jueUx
/JmVLg4uyphx+GFbXW9Er1OdC98KNzbNPlOIBltTOeqq8th/FdC6d5uPpsm3VHwg
sZzvkA0dKiwutPjltgdCFBWX6uGKVupKRTVdiXzXLN7/nHnLP7jC24xRm1JNcATx
AJEnft32CV1NqivJeq7x93sEtdTOYenGE6Vfe8Zx8BK+DdjTUI3nj/IAH+tO/hl9
4FA4JIy4QDLoq5mHTPtckaWb1hK++uc8JfB/qFBcqHzYaRSVjg+cxA8NlqTc8Dea
PecsNg9xW+v2PYoKhKPdnIVvCLzsg65UZ/lrz6ikyb+P5JUIHnJjEwZxOAujjgXh
hmtlgAXlT2aRfzM7qpmwFh0A7ko0QmtUTrQzFKXH3BAK6VuAXb0qegnbyIMVgIdf
tAXKg+nrTmIM/EKK99cGHSbF7cijpP8ENKdFCz9cLw9v0fbLEPRg3/MfhwJD98n0
CL5fHXzpEjWfHCZk1C0k8rNSgqXYJ4gMjsbh1VuEfJI1DJO0KQvgGJPrKVQAFDXY
grqeo6F5CxyZA1iWlD4e0+9KCSpAifNlcgJ9k7ESXy2J0hEDb+O+9lCM7YVsFvJ7
5qhJPgBkqzZLCCidw8Hjpnjj0799ptF9EtrDe8VIUA7MaGF5zVXk8LNjIpb3UN8e
mgxa+I1xbQmKIN35ooLvN6XkztzfTdtKyaYwmO5h0RDYfN0IStSddW8rUGvu23V1
NU9CdXHvDkC14HJ4SnLUyRMn0ntg5iBY9+U1e+LyPLa2taiM7Fmi4Pv1H4YFKtlr
W7XWtaNPvmiobTdCIjSRUwYXISAOhnpujazyqX2+b6bzfAvMYKJvjGrogGTiSEkE
nQOp9cCRT5pA2VRXMix6yAHH1c3oa5nUD/CRoC/xVKYj0/cw8FcBgWlxeiDri73U
q3VHlFrOHCDLhrp5XCRYiSt9w2ABLIp/jY7zIVVFjYiq3FIatpVfNclk7dKzxzYr
Bhp5IGx9U7IdP7lx0So+tGW1QJHR1aNnyihaeS7AQ9JYl7xQgD1dC97HVb5oFGKg
uxnLqrTEwgZ/wbr9G06Ubm5ubCH6sq0vhChQ6u9BSVmCHQjbtqj8/gehHTfcLHRw
WjdVQ4T1Ip0YBhRhrVSvNvIuPz96pAsP3Yd94Htb7PsYKlezn1mn2QGiDMBOIGbu
thP5ZFQi5qKn31kW/MjpXs7K2V3ZJyFZR42hTsr1abCTrYU7/Jlmeadu8oiVR397
3gh9EOzkHky3yYmDjw7uswjRVr1ApkGVmmiQiv7mLHNPGUN8mMtuilGR2NgG7qUM
td6FWcum7ovvcRjcGfgnW32KilxHMcxYU57TjlDqJue4uGlHlJ1g46v2fSkUhG3+
AIbt0V9lusS0NaQQK9R/GZ0jdprGI/jpXRRA7qj2xGdIJnA+N89qRBgZ1syofpqG
1iRswWtIMLSDa2AyckXn/bFcso1tm6ac44DAnSJl/64j+OdkfgofxXbNEjdBi+el
FymRqz1ekB6uchIoR48OHz+X/4XhexuXYdeD9RkhtZzbHvaXXm6NsQ9uoOxTmrU7
brBrVcRkO9JMJ2j9lWtM29eYULlAZzFVp3tRjtUs2+4XoKiuMu25iUHyxuy0i6aD
UEkru0i84zzTMVAgiXXrbsMzatyVOdaikh99bxvf8c4H2PoeRV70pRAphGbBOjiF
vxBqM6aV9ayPT3uW2JBfHXPZK0M7/pIbr8Fipkxv5zOzCxswpml71RN0DjmoUNic
xfxSap1CFL0LEk51eqVPR140RUslzqH0OhBY7l8p/Yl/et9aoAZYIHTDkDgr6I7A
IG8O/uZSD3WAHAGfGR+5mQAtyODnDRyyZx36/XSt0irjrzObifynQnTKIWiak5d4
vqTs0UCq+yXpIqjQcLfl+H5GCea4Fk3TTY3UWXsEmUzqPX2FE7rEtKm4bDBzyxvY
4jou6gKTFoU4PNapbSdl5TyezopMus+61hrss1hDsiAsWmrGBnX+z9iXvTzNMY1t
LrS6bB/XlpHiQBEyxoK06Zdzlnj8sS4ETab88GncutXKia007dG64B3+8DivyFfr
W/rh5o6l695oaj+hxaxbKdjZvkS+3xFykjcQ3eWB4Wl4JBLUFkYTtK8tZK0fYVOC
74tv12BIMav1CdnJ9g7hd5S1pi2IYy7eNZ05pVMrBjzeHV0TEwijot9eBncGGpEQ
x1QfGnc7e6Nj1CQjX1r7G5U/eRpyXcEAQHFV0oj5CgW0AARpYQ5yn/4uQsQjxUdU
r44b3POKHcKmMGNqgLsDEb28KYZ9o7poQ1u/qOO9dCnUoXinFvzzvlX7dv1zn07I
5ZA4Fe55BDe+at4HC179y2a9xm/YvhnQ047hcPkxOV12jlE2Ll02TpF9DWjghfXv
pU8iHkJWNSyV18vrygEmo3cJRycVX1bvknWDCiUQeJqVQyMTXcm/ryBAxNZpfZhZ
4oqqoWJdLVmza20YPM/M8lcDjFwvlXM7vNpC+YjO7fCWdsKTj4l8ISFARMzT6kyv
yVEuTOyoM/S3X7nqBSeeM45T9jHEBmS7/pFcN5JHJfdbC0qoMFH5Qf2NWTmCxYfq
4bSWMdReSKb1ooBeLHt2K6C+nfA9ImUP+34n97V8wrsOo+EX6v8L4pyGAZeNATil
ngF7PDZaRCeJ3lD63y85xkJ8Dwwx+MqFsHdyMaLuCH8ZNp6R+0t5D/Kr9ib6g2tJ
JY3YOd2yBCO/JyL/O7tMDeJDc0CgubSbNmG2fEF6rAn/X9jfhXgGULtn3bRvYRiw
tEuueDsRomUSxbsVo1PZciZV9xlHD+u5mRzVKl6Zr9zQw9CNcyzIieoahkWyx822
x6kvOs+TVyCd1v7yXyZfuXrV8Upxt/epYzuAMah2QdhVmwbThLqfhflnPEqK0ojW
FQ2LNZfOLMAeKsH714NStq6hcNbPx643kCrRNPM6mIHmvvPqBopjgie22ytcigCD
UNufV4qG1ay7wUJ6jCL4p4rsPPaUY/6/vfwbh0i2AJKENw8JHuXa2nwkvovtZb1+
Cijgl9yiGtpkSps0hOPNbLEveAARGGaS5R/+3fKBLJYI//QOUisGkRuqqNqN46jj
MzzCYZXtQC1qMqiLRvlpYsl+QodPKqHXyHzNj/HViuOCH2/lha7ZASokRvlL73GC
C9g82hpt/5sQm9wmQ0gGA8YDWp9x88WW60WVgLWWAaJIBLo1zSIcRUtiMwlXd9th
xpOkbbrPm2qiiIsldEue4QxkSuLuQTKwqfm2ZD/5465NA68WQAzwN96yFfQNYBwQ
HIA2cfpZVuARW/IFeNlWxVUi/6Ex0RnYeXM4BC3tZg8WQq73ScakD+4f5GOUBwFI
WbtiHMB6qbDx2eEmKEF6WX00qMqDjq3kiZcI4RUfh5YA+Bz/s3YEPiQClPmPL9DC
14aNdWkzfqyRAgwmppo84U+HlKHsnU8w/yfw2CPzQezho1po2Fv7J3qkRdUvcIJ1
1bHyzW+S4OvkoibWdQHmT5NH4EVzCyFcwfihESM0zDmMTSI5i8Lkw98dHEk23oUJ
CTqJK6mWa813acpLC4UVzAds6OA1uMixCVc4xR/1vvySBTxFEHVFU3AFo37u++EQ
CQ+KQA7oeNY9Jyd1vMXmHVz8psecaCXtyh8OLQBtZ2L+AJELwiuRLLVqhi6wJ+Cc
Udkb6fTfqQsr8Nkh/4PT2Ex8GvI8cCmVaUWLgzj2nIw6sBIr8aVdfzWJIpbliwuu
YJRPVhjleG1NWFXYyOgr8EsUPYq6vfDsl6Keb08DkWiH8GP7fiOtoxBI3E3zuktQ
tOPBUYnUOwJQ1o6XCqGbtzAwm1uqJXewOW6Mal2OfuATXcyqNMtMqmzKWogPcS6e
CFBNG5H9xFQxhkSOL/R+pmRdT6gBuE5G8hhIeIYUTpqmy4s59sEidN/JZGgXRnKY
3WoqiTDV4xOTuUbwMafTsQpwpO1Km5OrnhdtzZ/rGvEcB68hf4Ii/BnxQWoCzp7C
Fm0hdZ/WCpl9py2wIkmCImJTw/LUqoXUkRW3c0EWOvMX4ktxBQ/0/TcfYy4R+N/S
i3PSpYjgqVfNcdh0jFIv24tPGmOQm/hVn5av3qr3EtrWXF/vlogjkPFSaHdWCz8u
NdqNPFxujvuTtCBV62WuEDHYubmmU2DiW4GWHcHJAaTTl9wuEfq4hjj3St+BMT43
el7qaHcwpLPKQLW8uFgvZtjcf9vWYabh+vUzywJ7rImvo2yjd2DP3nYoFRAYvTeL
ZBBcW68MtZw71hjgkRt/4lDvTjLaJzCyz1Kz7Acq0J8F63EkIi0gQyRcQjAgD+vS
AECaA6grL2acZlr1hCwFd1rfwyeX8opuhxyVzsnKOF3Pdsfpd/a3Q6UadyOw6RYa
JOwLCdprZguUYqx52EvoCQf0M/5icd3hF3ZPHcUSb+WC/WfwLAzzgo4UORPY6AbV
84PT3zXg6QNBtGRO8UOoRPc6o9LxWpsuAWRxaZDH4TElZ377R/978MLzKpBMPQNZ
eWDpRn70SFnOSxLRiPj0bHlSU15Q+1NWmwNERHYGEbfpy1gqnu0APHDXWFeaLXvV
IX0ESg+VoTbOMMfdZ6/+K47tB/oiUiKaDIJLa6rQSigW/hNXghL40DXXVJDsDjXi
7vv1NVszPMDQGMrfru8r9+k+cdFv7JurBWY91IxTD3thbuLDzktIxLMgZq/aiHrB
DwK+xHdnKt5t4HVdHRDPBdoM3mHNH0tNtUKu6jash1XOhfFeTf964kwmxRTQCb6T
8s9zNPfYq35Ubd272s6n5qi7o4qBOx0mvITWNHekN4WbKgIX4RIEpdfBGjCHrNhl
Cd02V/rB4YML66xovcnHAET1vuFm41ZithFbOyTBxQ62SgXd4iY4Gw0Aegc2ox0i
0A2ehqpuxEgXVKe7lTn/2xmBfvoDRPS5X+mhCF9bRXI7dIWOYIwDAPfybljPF/DB
0oZ2C/fnTppS8uFx37ZGeDDUu0LUWtyaL5cbLyGk0Gd1/4UFIQWl2EBJfSdptjxb
o/97mikIWKWigzYzVzk80sAmocQ3yISCubLi5ibchayRea40NEdlJmkA7w89olgU
YaLp55SqznJG68RmCGqSdDTodb9MdPzII+Az/80ImE8hXmY7kP91d8RFXzoZpRr/
pwgun0mLEYT3w6Mfp8emjHORrRFrPRDhiRB2DSC2GMBxVEe4dOUMKRjnbFuV5iWX
rz5BvyCq51BhHziJAdndRP2SPX0aMr8If4rMd3UTcRtpDx+RC45bS3J7gzePQYRo
EF7Iq3Xi62S4fLzk5FGYQTvqcdxzFH9ijE/GyqEhYKjzfpAMCbNRgxmZpwFtB4ye
jZefduTFEhokqI9icESrXNEd0va+bsnC1VQ+uDCts+RfchE9ECmKFVERsr4B2/H2
LCQ0DwXWlK6SpuH2RYtY23LYRkvxCXBZ232VvGOVCBGGD0piR8fO+ZwAFW0GoPqG
Xg7ASXK+/D/S1+BB8Bnvd6r7JgwA8Jis4XZH1lb4k+mD+aHkLqluYqrEuQnypCHm
hNxNwTe+XcrEP45qiu4Uojx6LFmIe033TCgIO2+npV2q5QXHo1rL9h6Up9kZjaYL
zcM+BG+iplV2FD8K1Hn210bCZdOXLhVoH0crFR/Moeh/scinioGEhF7TET55fFE0
rjGZzxCWo7T8WZqbu9+8e68rnm7qL35DhVUCXeFQndVANWTf250GPEOVcxq8RXd9
4emqJVGKCH4+ovCLPOF6uc04Lk8SfhTBjgpcZPK0AK+nlFwZUbVTmGRI6hkh2z6+
t5Ghr7AAKju7jRYlADa+qJxrLMfL1fTTYZEY1FnjrRTr9JT9xT94rCpuM7+P+ljq
3ebdaU7j5DPb6JACqTHhgL4El35bP5bVXJyd8BigtfYHAK+Dx3pYEEV256q7K4+h
eKnLaPi5jFlLU2vESLIa0Yeuoi8EBL/VuglqIBTWYpOzWqAj3kHw0s4xtE7mfsEm
U9qRH9YZDKtVUDgx0wfIw5Nf0E/aM6xuTZMw9ED4tM9XCnHxtuRz5IcXnO6VH3uQ
F6ZyZqNCiRbSChpONL7YPn62g/C3jMa00lzUPer9hHWoSyI768jP6YYMLALpXwmT
KAJqC3B/TakHF690ZkTiQWYQNdMDm/1uESbZLsqr6YjN3ZFw7yV5l2+X1/g8RjiA
V7kt3caSVVtDYMKDYyXi02RnoEwdC0218Nrb5vlGheUuvrbnNLZf6b7bgvcigr3n
N8Dx5BNINOJau5mc2cSaGv1jsnoY3ascfuIVB/uhnD9F99cPCkI6T6y8LrXdLIk/
c35IkKU9AA2BafbIRtPvwV0GZDCmeUF3eUgoo8UEj0UGvm7OeeeHAwp4gruA2e8e
bS/UC3yVXyOR4mwoFWaXQKil8RqNLsytp49sVDCCB9BnEbZ2ycacVxlu1zkDqbt6
rTHgsMbzLAu6j+EeJ7gA3Y6sfkzZNasqcYIyKkHHwaH4ZgT9h+9bMWw43sx++65d
LwKqkAgKh1RMoa8N9G1xkiQpLXlRLHFHqh9A2hZt5/Lgh5xOZ4pvGRJwCBWlWiGT
kwEVandvBbKpeC0mNoz3qDQ6qFNCoMLJVF/EoaaUl9+D7lDsV83pPczrMFbEcF4u
nvM1GE8Bj9Vgd0z5lGR6yyjllxW0QF/y+NjAoI7nDaQhVul5MednQc25DNI7dQ+t
+eCP70JDN+9S4Bl7sCVUnTNRN8ORuUPXBoczz0TM5rnciovbRC8t3k7ZbtQ5dWKa
sIadtKVHc42ZXxw2ChORR2ctOsmRW9QINvS9yFkB3QtB9T4gTBWj/VuB904IvKXq
kaAPawuDCSEPUvgyDYgijk6m0wc2l4miUnDWBjiaddEXNaJBZKj1h9qAJkZK7WGs
FXLP2Cn54yjqC1aJZFKH6B4LpzqfHBrwQhPWVfKg+I+0aNXTFIpXWZH6onj4kn5/
YVCw/FFPU3Ksdf8vAlWrj150rc7CLkFOEuRnNd/E41OwNVz3ZWmndsQOGskESOZY
ouqy8tC0s4JT+b/sth/154H7kXah6XLOj5nOHWohGjrWMOFo51uLqtYGZD3idld3
wR6lwy609P0FD6L+8DAfDDCg3L8XD9M3yDi3+2iB0v6lWTXaxZQa7Sg7DkQ9Uk7f
ErwLzuf5EneGe1x4xbtKaG/TeTyqwCmfJzdoot8q/lTxy4N6/f6WpEdTumajvOa9
AXXm5k8jdaC2Q6Ch/qrzXvtFNY70d2jPJOhVRyNnW96KfeIHKvJVx1m0K03vmV2t
8OUqanW4vg5AWjJd/uulNSOO/nOeVdgsZgsTGF7Nas/ssQrfSWOXJnRZihz3zj6r
EHb9bbHmN8yCXqoCZ1q/ckoN6N72RsO2nBMIWfJlmhz0GeXbZVdgf89Fy05LvcZC
3qg5dgsiSW4xUr6rm93YxUtmDd4ShRVv23n/JdqtXhuAOSMzPSN5VXej/FpdKwK5
96ds6Oi2ILyNL1db+hWwHlF1D+AhQTfojaCbLgRkBECZl37nZ5t406ZuzKVGEI2d
12TjyuiqtplccZUGVAgAzLBpzKstSmZnSnEMc4hRsvoyKLT3Hk79QKwynSchtkgS
IsUo7MczDO0Nyfy640nlzHaaisHpPPfWrJab48SdRxLuFX1w8e7P0XJQNhC3HHsW
zcaGYN/RJN+4r8n4bNpEVhQyWVD4+QAh/su8RCHXfh9S/+J8b/li6V5QxZfuIcIu
gutLGGuk8vyO2zUoxB1W+VP+TEcXwbfepmlFTBkM5JJkqifZ9qDqgrgJLnhtBJ/+
nYGE37LZeS490e8J/PRTCv6gu3I0PQFu3IQ9lBj7sErgFUkI6xX+PG60csuxPdGs
/arFSjyeAszUsftt49ARu+WHyfxcct23uBOaSW4DPutpW+44fWtCki2gjrsnjnhN
jGh3h8Xbdwafqxe1UmOo4uF0snizH+GfgimMlahdl5rbAO0zWobyk0bHqPgjw0Nz
GyZbgExF8f8WTRgLhSrgPv+R2TamHcUtit86XeNJ70TNMYO0RovRvtknigdnH1oJ
NRbYl7pXo1iATx4s+mX0UUu+IvdwSgmqqc9upaxMJYASZBvsaFlpxaNJ91BfIFz0
v7Md2ZxVtZagSHrtKczJWQwZoCX0xlw3rWWsWGeysFbF5Z+IGEpp7OjeWUOs+zBI
DPSa7K44GazEJR0Js10pypbPC7sv7NOuNygq68Wy1BEiq4f/KZyuZlrEj++Yjkps
d+QQOP3HW/WTpAByR34WdttHuxHK2yIINVC7eOTqsf1GMTFbomyfICzZMAwGwc4H
Ls/WhqYz6UNDRhSQfXj0pENgnJYzTTaIAiZ5rXYPjwklbpFZB163MYXfMz24vrRv
1UlMVV+rEFCBheMy22HXCrSV+t5sDAvKTn4jlIZChCRxfH/31LLl+EENZEa3EE6f
93Ezfd8dA36OckCcyoqIZADQK5A0iZmMgfWSmVOHzkXwa/bpV5dHfRICdxEL2PAv
CEzIPAGEdbGu5zNqLbjoAEgV/JHdlaeeoWVanFRr/1BW1OA3W4XEtndCu7Kz3s+t
rwk9A7TIy6Y7nkXp+sx2GOFWUTqXYUqc7C5IqrMdkVfPKGEzBrw1Gy2pJHIbEx2U
x7FIHiqehQ/2JFcnGninlNiJHz2TBgzx9vYxxtrEe4OnzT+pm/IObXAUSV4st/qG
EBUFvO1yDJxJZ6QrvdxTxbVw/0sFga2tqNLDBcqMh1s/BSfw2EPUFGwECugKvcfd
R+m16sU0bF5EveNfqeGe7s9v+WzIzjfO9+//eVagt/vHwqIop3UuCdHoSbMDBhBO
PNMGmrgS+FVdsCLOw0MwZdrFbzMIg54MotwJ3JR80cbvzXjFt7EmzdclNCk92fsC
HmGNR8vYtXmL9gmcluvIOr4E1qEoOGqRLZnHako0/Krl5nGKFoJhB/MedqwFREf9
39DFUuCM3uXyX2Igv+yIj9SXNV1txrOB85+A7Wn1YfH14ctEUbrCG5HECt4rNXZT
hkKsE9MtRK/OTjtUEIY0RgsgTqzGCrFywTm1VrwUCblAwlXAcRDxInJnMryjYQ++
mtvQ9/bxbPY78B5PRtRleMlYmIGZ4/oBQp7kG0Eq8FxuRNM0y6l1f6w0peZDVerW
vPjdvqa3pSIeHCfpjUSgsWS8iPvIC+H5daN82k+Q4gtE+qKdFRWR9/MX7eDYWrJe
9Wle7LFKk/64RsxoTPwq9vIrC8XpSE4N6eOM8sQNnbqzaA1Gf665qMuzRgfZSZey
TaMNMh+lPrPrs6amiQNMlt1jyjgaolgT4+U32S+bCKb7nLaz2V4V3Lquz6SVDNVX
z5wXiG0OUW3Oo2GeTSgRcn16y5U/XfSery4gRpIpvf9ikBW1Xpcf1qrWOIXHUB2x
V1hVmBasHbbNtK1uaO4uq7bx5LJhOu9VTYe5g+P2kI8iO1hSO7Rn+D8NYc9MuAsp
VB+W58FZrHK+YOd03Tew2U3wF4Cdeipg8b1F9XH9dLjpuwZazDY/vmOjmVmmZxDz
8g5kNBP89YSaAH2EOU6VVFKFRaviVPhO+4wZ7Lr/+dPGWj2oCOZ5j1Xzt2CJbwZb
/ph5q7G4KLFQKZBSwHdnX/2QwEhPbdiqrdcrpc0nF78lhRsxKQpCx43gsUeEM7+1
1EUEJMS1M4k8sSNHstU9yF3gNF2LhWOtqhjrWd2Hd6z0PeYFX2WL3nvgs2Ti7luF
fN19XcCrMDHVr9vF0ZTYJHsWsx3yOlR1oRnmElDBJ1dO6mLenUlNCS/xxxPVTkFG
igvZXr0Wk5bn/6kwvZdMKp9EOnzHs9BjCJfXapAv1UKJU/rjwa2Y9P5Dq8+wMDBC
aMCOLZ1q0XTM1NZ1Yzudyz4OYtvkOLCSdesAKDkZnERqiQcum9/d8EzhHHE8DSmC
PyG/Yef0ots5DuL1ejH9ndMmC8haO1dDPADW+5pPAthaqXdbBDUMIdBkqJMzJUr9
g5/ifYcq7Yl4gD3kXgQxve5+S8I3n8nZ8BFUVHmovTUIm9Ys0kfhozBvioTtfT/t
rfthY6UlcyMZqanUw0GFQCtE5A4+pFmT0tlSXoM9CQMkRI78Shn0cCihYHRctf3s
W2BXPBB5360fxtEuHBxDQtIuEsT39oH2jFZiOdTBwSCO8d3pQAutFO1Ue+HgSp5T
GLjI2e6tYBG7KxLTK7/lnTeSrRLSvvmQCF0Ow7LKmiAqCBj3TevNHwNA/emZvY9v
FMmT9LlSjWXJkkgwL9CayVvw522oddK+yYR5jDPz9Yu3k1GqC8baiCrZMZ/b5zmO
wLuMajd48faaFQJpHZmwWWUCizJaKtqAwijKrEJVSbjV9NilRV7ztrRGTXdkK7aj
tniY88BKK6wurbLOtJ9Mg6YEmy5ZTnl42ruAVPZBie6cTmeKA9BT3N6H9C+Unto7
BIal7Sku4QFacayOMEteUKufrAyDrCheC0JQERk1QtqqoO1J8a0FM0vrGX4Vkj3b
tV7KyxFonO8hiiNvz/4sZjE/z7Goe8K1sRCXBuXWlpal6QEwz0zqMYGCKSIYZKuX
kteSezibaXthZW0xixOVTHifnNIxo+49HOjC/zA+N/urK6u6cZORCRBEG8kKQtoU
Nq/fltvBIb7dlmMPogz36nY6HtClllB92GRek+n7fT6LNWXLvCaMKi9kwpg89iVn
06xtKMedXOWhu9zgAFH+ZlPRbwP4MHlNeh7B6nGYCKA3Of1Es/TGeLyWehXmwa0O
TAWfOsY3rcQ8IsaJtPmJsSd0vglfZ3PbzrA0Lv1Bn6DFgbihC8HCdaMps6qTyfoI
aFRKV4s9Yj9ziQ59yUIeVIK2mqheftcXFKbzcGLQ6rgJxMGiJw8U1rMTFOTIjToe
HeT3wUCxZnoo18tjY49tz2rrN70TTvY+WfvyhaSH+UljYN3/DO+m+kaR12SwdE/3
78hSag+zlCRxjU82ge3BlxUP+ViuP/J7DnwAECfXS4Gw8WwC5iZMVb5RrS7ijCqr
rit+NpdXpNUW6eceR18wBSFN8GSsbRvbQFWUPQAU0DtCP0ETBNZRJUn83BES07nR
mc75PZnTrMUbCY8EnNPHEcFRSjmOBzQFaVC6jGCoPSgEde1mdsVMUHgo0fyDdUzl
SbbHTsJX8+QQnetfJJugWIpbPr36+FbOI1wJl/Qb4I+CDciw+3zdP47uG3Xw6kBO
47TPK37c5484Ia+2U+wlXDX17GpJjPQsPyNWNlmaBVvRxGaBOsGe1d4JMAgWMTnR
F+hDCv80b0SJU3HYmIwZS5xxSuU073rl2j9ZQIDEgEoc9+sfDCvRvgfEfH/42oYc
K86u2J3k6jRau5g49qv2LUnk4dtssShyuSxardeFGYq7EUUYJtKH5ljW5ms09JvU
/Dwqh/ynPW2eFkVfL+uUEn9OHQGtwE+z7oSG40drq6E8mS3Mpoxc2JcAB+jKVcTg
Xw/Q0Nux8vroO29SAE5rHWLMjUh5p9gngzC9Xpb3LdS0W9OaRB4PirGE5Qh3J1kC
mIbSvx7A9cDcQd8u0AGxxx4roSZ8BdoaNHbO7q1omzrpDRk6wIoN7pRx8LqTRMOE
72cQdtAisjaFzFMwqIsM4AzXUV+ziOTj2ETm6ysVmVi2RwbFti8gwioAjs1+TiEt
ZdWj0KS9+YryQGxCgN9FzAxE14dq1mM7SOEVSwS0snazDDkLSoM++pLMC1VDqrzK
0jIpMGI2vWXoQ81MUvcgXuX5wS+qvIE9JZ+9yw/YVQ6M1iw/p1GM25+RqYGIMa/n
zDip1VwzlWH/sXdjbY4tEl8EF1w0QlEXPbp1/ig549NPjjC2gss4K/ACkIaQKNaz
0/WoCXHlqSYm/PmKnFxXgZmOuwWb6zRYv3HvcN0I0wog33RYVyIBwvvOmCWtbYrg
rwN4bWeZKOvNmTfqVXFO3hgoApooJH3SXIEnuCOoytnyP7gPM3QPXG3bg4S8DNB6
F6uiA+9BfktboNqKt+T3OHhwrtCpUHgqUh8K4O2RGI+b07w+JCQNZEFz87pioESs
Ze5eYxUiynwTmO6el9feg7GZQlbRqwt1zMNaddg3fOAjZ1yRhE584cWJXH6PpQw9
OC8jMZ7blicMulzUdGT42VDLcF4QfPktYWFG7zK7dOc0KfWrLBqxOmk0YLBfj+vu
HV1znTNJ7ZCXW5N2Wbr6Rl2xec8ATLlGWzqz3P1sk8keAAZI3nhUAL4fAAOllbSG
7sqL6kaTS+WpeulchsbRH+YUWmBMG98OiIb+dXeyuztOJb2nuWCm5V1hFWryIVHx
C6nCimV1cxQLHrudhhS3SjH5B+AUJolb8ZG9cFT6aScPKp3zdJGJqLr4X718Nf8B
wjg337KypDSROhfYG5mSMFYsVidElHSsIf/jcC9RGzW/Jk3VTAdx7guhRXEjcBIM
5EeO7hlOoQCCTWeE8aeV+rMdgjsiZTyVV83N0/0CT3rV/Gv5+rXl5aX0UsMCgGl3
1Gq3gnBvoBxn1DyFQwPVIDB0Rc+ZJ0jFTS2veM/lqCvKw6YTiltpgyhD6soKiQmb
kP5W52R86fbCz5i7X4DqNKKGu9Ka+Ao2GadLZpGgmVExKgrKmFdTBDlbCe4ZXJSc
hu46OhjneIXRok4utwMBNm0IRANZ5z2vm5CFNvfg+LR7t3N8G3Lwx45FUXxP39tr
QEv68rVq5Nh9fNrRkSEE1wcuQSR5go1RjG2Mve6kIqxqIUJt+hi70aSbCdRrJ4Lr
zvg9kyPJdHWQSRbPZXXjaeC8s2xlVq3n8NwLvfRLcFq1IOEPkeGBim8BIVarIUJf
BsDM8HOCIANZRwDC7keiYrWABzkgVkXOFU5RlPANQGWVUN1KfurGZ+JtclP06Jyg
GVJ6XQzjGMSc6bNmlWsXukVrSCQM00buuQKLWPxBnPU2S4qYOF/ocJh67r1XTRs8
qxfNlaFmhyi1MGyUkGFPJ1JBOhGRRw/uiHwJ5hRcbuNAWtO90mBvnaDDTgKii8T8
ztYxbtNKpcmTQTuudj3nQ/9WY6+AE6dHPLvcF8vcbCJXPqMf2njJP4Xq6HmIThJR
Yj2TgrmDysjs3IuRfqZUPUYQ7BJnvTzps8b/vCzn+9bEHmCVu5pJUo9JgpHlGYBh
ksEtJeSmUV/mTgoijQtxYEBDm6G+lS9NG4I/vM177eikxwQEQOCWq9uv8+EV+H3t
LwZQ7xm14ItQtIDgGiQjzzm6CgdUJI5RjDC5l5osWcAm3P4kngr3eMzhPDbmNanw
MM1ZV2d16yY3ZRb9tNATICzVbmDlSEITpM9VlLY3JtfYSA/p1I3dHcIDZO1DL8UJ
6L9cBNIaqEGOqPxNPwE6Kn4msiXDv0yytF2LpLxOvKLGJ4y233qAaPairHDOxp0C
aFps71LFeqMXNK9R2GHdSKWnLYUeLQKm/DBNnNqKbalWFRgLNdRr4PPfb5CNRlKW
yjZreHT7N0LGCErcc2NVoBtrLUCBbR18p4pJyzHTs1QbJ5rKl67qtuYzi+qUYLZ4
vPMisS84ucwJbyFvY/g+DPT9FGw15HtZfuz5VogX1fTCHV12lLlqDtKZZ4WPJUAw
FsIqzZxtv3T1opq4Nh7Ot56l9wqTiomQDaTBTKvFwYU0AEX/5mmYz8GPpXyLDtct
ul54XX4xiswUxRwgllktFFbuP/LHmzQgKTw8HJtvUBo+KQxvynSIOYMN4nFMkrm3
bTnInysUkSrJ6vSfZRobeT+u2cM/wUjZTMyhIA17iH/AtMT+FIoWUF793he2HfjR
n97Brru9KhSAw71A2YejrsuuLKs6nNn2XCDkPDgZZJN9+k4aNZQiHO0gztX8YJJE
Az3y29wc4sywRFXPmFO9YcBCAp0CoCvxoiy6ZrWIP4ltbvCyIaNjg8R2zBMHLDJ+
bpiKp0KvSZL/OTYb7cJPC9I6wn5SvYqYNPBwwvmhWQUdhI5913bLyguoexKzInkD
+xXfJ+tmWl0ANJOH54oaI+M2lK9BOQr8r8edf9lw7XCc2BQY9Izesl4eOo0YqOCJ
O19SQ4Itj2jLP0hnHF5Y2SPX2Sjsfi/OoN9Uto6y0gHlczg8ghPRo6bj4bv3VMFR
ww8o98OJ9GrpYZYB0Cy8kYRi8av3DKfZSWozuNxArT86G45Zoi+MvXTTlDbFSrJi
B/QeMhv6HwMElQrPcn38l7XbR57ja6tVbYzRYsAlrWf3RL0IxldvpPSGih16u8Zo
S9HjYYmYa01/hEIug8XukLJmDhnb/F+K+kt3irgrkgZwfi7kDsmxRHSh+Jof8cU0
rmEBCa6jBNnGKdG3LH/+1YpUHwOTijUGrcdat0tT44D/y9pifnFNvaT/NZPxxB0J
j18LAJBOLD/h1EGob7bxLHhwlqdGrhj7eUtObL/mMQJEBCtRVS3BxvniimsWA8Ji
mBVXGNQatTh4fA6gZBvSpCHuWhLn06wkStT8cUpzzr+O5dCTeYCd4ZHlzPps9d11
XhkvhBnbUqN/VBD0+dGaPVSDjvkP12GeC0WmxsPEP0fgOhzj8vtzXE5NRWnzdNSl
bcNMq9bzXUTWuomtjlmgOyVfeA1JBv0maIjbKGwWew0y76ohryrWh6USSCcm99Vy
UKPrprWjEz13FslvwuA2X1EfHJk4EdvIGxG14Nl8j2LqtlFpeOCl1fR5UGcMP3zG
atQJzQJE4dQSxxVt09gsbuXpDkk+W1aeDh/D9crknLwAX4fNPExm5+CbF/l/02rK
ajUuoWQvXAJ8Sj3NjmNO8m9QhTQyZ07jM6fvD7Q2PGCZSKgwx7N+rBPU+woXarpu
FD/VrtYyU4Pr5+Ud0E93nVor7KeUE3yFZbfi+5VTDE2njyiY+eVxZbkX1I6te4Es
5je2rJJFzO/evPuX/sH2Np+Z4WfyUqeUABP05VSx0tXY0iF0dhyDYeD0w1hG3Qis
YY6kxbU+QgWUhk3xE/xcwmokN9VUmyPnI99btHg1mcBzGbCiXHUfZiEILXcXS0K5
XLSVrf9nAqTn2qO+h2skFQSvXm/8HiLKZUljc1W0oLDCpPt4yRpiz7J0PvEG7kOW
qG4JA5DDo3/+D+ZCuIDq5vF81L8gSIj5Aoz1+TpeBNBKl6Nf6OR5LX/jyTnWWvF+
a3K7cgZLWnPTboDsezrIMPtApaUMybZ2MjD2T+/B/y3zGH+RsNTOoo5dyb+oP1YV
yGIlg7HUfYAtW7/eAZ8bf7axhVuQ4P/6hQ6l9sHBsba02H0eN7U2p8iNngUXbpX8
0p06Ax3dVJx0wVKzRHzy4f6a+QglsdXTXa5basBoXi81XlgKCA7K/lhz2qQ4Uk8s
UBu9dqoxHfLHq7QX5xnNzBUL5EmW8RX7utFFzQ6AVFMaN7NLVd+cxoO95pgQt2RB
zFTJDnOouXXxkyMYdm3Hc0YB1iWRd40IvT9kTn6LQ9jDWqxbBqiNbzVpftxkYEx/
I/EUgG0FT34e89aYExl10Wld+5Hqkh2npMEv7K4EgPxpwu4rg1ax1nOjtwXdPyWK
GWKhKT9e5AdUaEuwBi3l87pRpMOPyck6hovvCcWM51ZYxCbG7gfZ6DF2hyB6Rzcg
csW6otQxcZYvcGXyA4MCapwo/sPN9Ua7LH4v143Kkxz2FXxQw+LePcW1bxbzcDBE
awTFfqTHOjiHYiZpJ1fUgzU8B7ODWI6tTcaJk4ZnTwSbKMBmu+P4KmFDgafffLG7
ekY7bPuuzj/mewYee/i/q8oLPmtLOyDqebGSFAIjnkaDu/TF2avFrxyPeeNHTRqa
1nkEnAwJGJZlHgAO2WJAUJpNYmQCVFgqXQ1mn4xK1c9EJJGYG9GC7j6LGYoeqgVC
2L1pGrQTLk9NcswBUx1zOfzUIOruJuIqwzWNgeET8jwJHC+zE42L++J/6jolFtAl
/vvKGhFgpt/xklMKT14CRern3rDHCgAvQcYlw4rk+ISv4eRJCxFHrCmFVRR8mPtb
+DA9yAiZSdY/RBNIBom/sC7+fgDSZTTARktj8Hr9V8OER8rOlUgR0ftm+e7572MU
ItyqGDqgWAtticUeUAp0QzKkUnhOkA3Q1w6GxeKtOdXwjMQA16vTjAKIWQC60pnE
d43wbWB8L2HZgQjhhh6PXp7WLtG8voBoj96e2i3bQrA8u4+9iYmH1OsniAS9DY0u
SvQ06pzjdKXIwA7XPO5NJs04bdLNxMihl/jhSZFO8NLORyQHvOAI7jM+0RzpaVlk
PPpHupd7rS1T02MdM4FJsfams6ZLMHzinHY2FsRIQ9st7FxVtp0DCsNW5Luii569
WW+iXLum9OwHq0XlHxvqMiriFykwaDCwyIt/PoCrHsZ57r5+Humpr7oNEE1/XuOd
wLQ9fYqQIRYdJ7ngUh5ZInrfns6OLlD1dxFZ2k+jEQpMqbtuFVKWArve3t9q9MjF
x/b+ZBXzyAidrMktgmX4XfyWLWs/NSX6PVg4VHfORtcoVQob0Carht1Z7eQ+V17g
LMb6xTd0X4FsmvI0uKhkp944YA9ijGlhF9j8nQkG6Rv9a0LteGz7mj0ECpMcgZRQ
KQRhH/F6uydb/Rsxt76cfsbaQwmHtXtqNaIXbxsDIH8Gb5Dd//u6Uu58sS0nYygY
I8daPYWiS1Uwnbs2wQztHQjnxvQ5a5C82rViUDhgWnVHDwagEIf6+iYWwytNq3Hp
FbhGPSYuJ8Z10bpJV0+wtHIe+oAu0ZSPApm4DN7kg9nuKTS7ZFkw9HpEfGtULcXc
cw54K3COyXlVz5qFP2l4uVfWGul5/YkXsdKbfl/FyM6sdWBEOGq28PXABMo5wi/w
8mJAHEofkPHu9qjrk6u6HDKMaMMtoQY5QCxo/HHjo6Gc3YZR3fBT0+z2fYUoptP2
yVZa+JTNcoCgAOX2lCk4OYUYtSPYxcbfDHE3A2oGqBwbEqsTpOmN9dxjHHbIBXZ7
/WlhAJTUy2Wd8hnWxOVWglQYLwlqoQzVyJqYVQbvk2VuZ/Qu6eBBtsDvylMYgyuT
+rNxwRaCBeF9goJyk5dYxvvJnaBkA0mP2G4NzkmCBwK53WoIBMIzS+3d6hH4eONQ
FFXTeFooVYsCg3HEHEuNOhKL5JKkW5T9FYyKWyJvCPJa5owUKIcl3yfMIs1ukVwF
Iy/f2jfw27XgGqzTmzphL28ibS6013G7cGnD6VG5F95GhNfOjKbBcfVQdVQX5hi+
nxWY70pElpd6zoFMuwY0SjTFxMjlrfYwxXxJWXL4dYiRFlyIfydyDZ9J39V0OI0K
OYTvhrjdizWh5oTv23W4fZApWF9VNkQ0E7VzspmaxRfGGpsTqkXbZKpJz2K0/72F
txsOv6XU2dsRT8eZV41CumO9VgDwpl7g9M934d4UnZ5mb4GJO1zuMpU7Gbn9Rjz4
PlhSi5YHebNSWlwm8HAB9w5Qs9bIOPz++U3iKEV1BB1ucfiO2luvcbZMND9CsPBj
Is2hHscWZ5L0hJzb6x/ZLEuxcX1MkIjHTZPFChxPlzC9hZAGuAvcWKXzXAYumUmG
CV4Rw20lMX5TnabIRhLHwK34KG+44iijz9XvjLAjDSuNgA1xk5li8U096X9GSExm
M8a4AVTKY98GgxiUMiSN8MLRtyf7MLZ3fuIb2iF/qJGKXBxpcpScaj0coujXC5Mj
4HvcuNka9bltOrGj0PP9yhV5SYgkimRCQUSt8AavxSTdAjsBMx5nmSRODSJaFqlz
SvTxWbxRe6ioef7jioiuD32/KFX8tV+/HlVSNImA22P2M9fQuT2q+bU8uJM30ILq
SW5q0/M8t2ys8V+o0j1TLNg459z+5v8YADi/whxJZqCiak28NNnIfDVhRppAcFYo
ZkXVRfe3mPARZlkNQwclwKaE9vaNoAPgw/XWbObefrun2M6pejbuhJcXtNecc05G
vUr+C03mlA3Jx5tUY0wraK++qy9ooq12yj9hGQgV6Rw9omWG/Qd1YTZnJJafg1Xf
c/qY/8Y/1gXw37xfsv3Hw7YimgudUi2TLV1RbB6BhxrZdqjJZ52eQ47PVam+VMiw
W6WmxHGB3ZSqxvpHlexN/FDEZU6JBU/82LNfpIj6wpkmNX/OpxFysQmIDaYtic7Q
0NfCvE3evT9R/YtJ4oRsbvS4fhH6+IbKIE1op4Q+k1pOg6CU9e8jFa+ji52rk/ZM
Dbufvrxf+YNIGjGNaeLo3YoSYk6gA44zSyJDr4DO55q0FtzJR7RgImhT9kJorpmu
9NccEAX37YsQFq+4yD7ASY4GtXla+imZlXfW/4d/fg6Wjf0SF1/9RFODZi+szN0i
/H/1AI0XxOLpOgVXNJdSqWQ++AaiNunywWzD1gsYDww9cB7enh5bU7BkKC9H7JNC
+n5zjFa6Omg9gpcpMkWy3Lw+wweZn8GPXn6CWsZvkglZo8Gmg3xhQ/LcegD0BFOz
Tmb6PPY7zldDflYmlVSgVbhf0yLwmRaQEbSv3vzl1ll9yhYRnycj9sSQZAfqArp4
UT+u8nYWhoE48UAz492ACx9gIW4KrWtBd14+jthtXSVsivVR2mCdkOzw7rcnJQTU
CNwUDH6UowePHSwvRpeHmk1N4km6irQc61iIVu3zAoCJn7yh/R+fP2aCgF4PMhge
/REFdsjJsIwaIesmUhrJoD/mLou5EHS7D8NDplQHlHlOEtAKgFlnYNwyYcbj+oEZ
H9fmRbFYZeH2yzoYsC69kENDSlC/atgKuLYDIdWWDWMb88UkH8FOhRS69GCcbs/W
PMAfXXfGNGb2eWUn8pI2LdX+eyIRzCDxF97YvkVtlMycUbjq3TU4Umd8Zq/aCMUC
hE28HjkQgJnBeDqG7qFhLwObVxS824sOpxzQogqkCtY5kbnnprRPbsFm2XEbaLIl
hUO6MY1IGGzACGzUuPt+/4V9hI39ROeiqvgKhwnl6/gxmmDk1of5e2OZ2yncnklV
KcRBOkoJzaQRoWHhygOK5rGVZBsKQhRUPhhbABBLji6z06bekNIGK+NY0QHVu4F3
oy3Yl3j0OulQyCB1aA7tmNuL+eugikmCHV/Ii93O2W5WypoNCliNTewOEVNGpIr1
XZU53kEaaM6SWfMkPjrRL8z0oCbflqD84ZIAn+253e0bEjKdcR/Z8TObf/vqiGBR
RJEVNWRLrBH5co28sWIGmRe+eFsqMMP2onWoAODbV6AiB5bjqaN1PSTI4sSrA7t+
Vq0vRua4xL8tdl7nYPEmzaA9geD+9xcf85LLAS8q9o3GPdlgzbWVKaKAjippjqRC
t4Eyv6YD9FYlD+RT6YKfg678NWoRt/LkMwG3D/NBRz0SM4c+a+VE5YubfZ8rNg4X
2Cs7puT2z854mdC2xxPc8cvrQW5cWA5lFncQgZvhcmQ767ui0zuvG7O3mXSGmgzV
JZSDMLlk19QUX+n2Kd/QSonsMJqkcg8QKvASuTiA5scwdGn8ivWZLb9/Lt8rYrx8
IlPUvQ+EBxzFYPKuegivKd0J3OukJmGYtRBdTStAm3ifyx6Lqeo+rUHq+D9yE8dF
YcGXSUVsN+RpnraeCL8iR7h+g7EsC6ApAT45ZHluKmLDAtTjfFH7xOjdwZ3LPsoS
c7nawZUa38MONboXEVbbuK4M+6DLFHU9dkFwfctpy+2Z90sCYVBAlVmipFo3BNE2
fUjiAX5xHfwjiuXDK6NyAOLxUPGjZXxWx4ju+AQ8HGgue16IBKg+EI4aUbwgigYU
A5mEH+oE+aOXFp3K35GWEaT3VvjLjaH0oTmJkEUD6RMiC2GHmdr25B+lTNVtw6/Q
lZ4PRQ3azb5M0/83+SGTV4FVJp0RY1s7LQuclmH7LxNO67CPcPgVUpfOpGo9p7Mi
IeioLTsXMInuE5AtRRCWGCyEqsFmxCKlGjGcvNWuU84YwcjDco+Xp1pyl782SUhc
JIjBSJMwYUoPxE0+/7n2nbMVrl1KfiQsu5X1R3Gqzth68DfYorLDlKZxyOqSAzr3
r2W/qTzZT69/evpTxwI3vOnisCuHOS7EKddmlqtiKC4/YUg+mo4W8b8CrQblABWh
MUIgNhQaI5uXni9/wlfo3V7iqjie0XKvvGcItRAXniIgwJQDD8UJpslE86C9ZI84
4VCih9H+XupQSXccVwiObq3TDWtllOtkIm+TbMtC5ECXUrONpqTSytVOV+o+2v9k
9NwFr+yxb8RCk8oZ1Z83fh1FUK7oBc9/NX+CFAklgGTdMCqUjNdM6AMJgr4ZEeGb
+ey/MvPJc+ONatVJeJoR9OVjivkiBLqnUooTTgTacZC0u0bLi7GjBg3ZXircyBCb
KCAzTPgqnDga5L95GY1iL6Nd5ICeXnmAHFEd9ltWq65CeL3DR2mhshErOmKvcsxv
vvZ/SQ6+MKwn4TeIEQCcBfDsscT0aKF8dSSkPlz5ol6rXcmRycQ0OF9ihBSAQ+2v
1cgKdnztV+9NkajC1XblT34RkJkZrxRLCFsfmZ2JnlQDfiRDnoQrp2L/99Oan0CX
752+DrhYFn0u/0U4ZHy4/5jktq9nx2js1nS787P0HDKEFJeyOSK90BXwZCJrcz23
LBHMtS/rRg/1NBz8yHyhkK1+UUwdZaIzbPQuX/Dya4SrkuiiegscEP1o62746P5l
Qe5Sy5VV07KXrYmo33QwyzUojhv5J0TD6CeWLykNbrNhTzgtsJ0HqEgmQr9R8aji
XKffaoQudeyqZXrRvDGPjYlNdDX+iMHJj381Dt5CKQl9Z0PxeJaQeKQ1kMbxvdRa
heNvD7epv2I4+LZ/v31ksgIVe6mFApkVskSLEe4DL6G7UueQTj3nZ43TrIvSWOG9
D/fDnPLk1D4b7VOgVpQPD9XaPl9loaYAekOuiuAW133LU3Fcch3+QeZ6lxRuIp4a
CsoKFH7T7+O3AQ47fWKujDX2jkuVojIZn3LVZKvLM3pDtE4+ZlLRWaKKColkwRSq
LJi1GuCAuBv1YbdCZNOh3Yx2O3KpQ6/HtDT3UKlWKV36me4ih/qgkZqRl91TuSc7
2wmX80scpEEWqak/CWEz5L9vqtXRZPvbeT4sccUrqyU6pVHb59flkRjCvaXoXWOQ
12eNyRWmjrPp9/S7CIXAZdAcwPRjJx0YHnRQdXoiB6u9lFQiqrpt5pxdWiplgdtg
cw12SSMQn1eePjx7m0qpZy1YHR8/I1mDX5Km+Cpfddqp3iuWPj/4KK/EdRx6HbbF
xcOf0ago+6x515zqU/g/p7+o1SLRsH6O0Uvfthkz8/09TukVBSTGgSP1GLiXAtgf
5Lcqwp5fmpKORaYw/zZCO0VVeZVtcpZpppXOV1OSO+oj7LAK94mTtSVyGOchE4nf
8frs/k3ASxCItqlwzj/A7X0PNAUmGoH1OfoozV9cf9XSp1J+wO0mFT8tQKfSQP00
dGr3WOFP20rdT/9o5Nd5v8CTVeoAZk+Q1fvyfNnBqxnJoe2uKyCMIUrmYhV5Uqsf
JCI5jYaR1AQO4dKT0alQqdbZXHmB7brdi4Dn6/OA2qYQGympkouzXUBO0cv1Df40
d90Dgq6AhMR5YfCN+lQeG5LENe1jZSBFf1dQEYlhauVpF1rLHJBpi+E8c5X+niiP
TN4xudAzEw5erRC9nlwVLbrzqf9gBwN896jSzwy3qclD9HvRw02Oqc4pmYwjnVbe
XnE/ZZjZ+rNEsSxoFqkM3Bu5mrFTyqvhMpcZC8c42r5D9mXLTeGq01Dc/FOwf/AZ
3UDYjBKxvlR17IcfzhtaO8hXIUpbFQ4OXIdWQ7IP7KI/bSmjVvYpqJD+TkiHV9mw
x84Qj/8mg2oajQhNS7vF7+p+jDa3T6KLCHqmkDPRAVWwsoSQcmlJLZhOxTDN/wQP
S6LnUArpdSjCwQBhhePYP4q2HqIAB9BbdmAi4K5bPpzOohmWvYh227vZ/UiSd8JQ
CT1bnnCDgAmDZtBXkqzBP3npxBzzzMx5pLj9pmk0aJX+oKCNJTj87URrqzUiw5fk
PgqExET2tXUkbKnHrPTQ0TNkR4gK8xanah/OXos6kf5oXUTt8ymjZONptzZoYwpS
9/Bz6lvEtbFs46SD1DjnSwzVD5xi75lpUuodubWsWePN0TLJxde6EkX1ClBXzU68
ZMQhh6ox9wVamK4F8CrDtGWaUTCxDpBbZfuRRBxBmLpqhMezUHM8HdZhZsQ/jkYq
U3ikDKQ1i8mq0eAROhp9q4zT0JxgtBYYCN3lQoF4koFDJWNR9owOjztNrKkDaG5Y
rfriu9Ap1mROOOaY3czNSfguU3vW9Qn4mkpKi9XCIChFQIigMEXkdZHUeOHgFYWs
TXAy3F44plc0wpbGR5byhQ9MZoVfON2yAFA4xOkxjFJe5R5LkEnkN7VnqtwheN79
vtiIHJsUdoevgxpo4/OhjfPtz7V8DY02gSIqenJCuDNgxzZs+xlkXc1O02TF7oeD
R+3Itr3ArPr6/FOEk01Zx4y7Hn8n24WjQrIov0qLvXb7Axr0RiPmrN8yp9Ez8zqZ
ZH/qqTyEQQEbzdhLMUwhAwoT3P3U3D3LHuyV3ITKFEUaLqnELwhKHVaLrQlM517s
ruOACtXErdGSMrC20LSSJoWGdf5HUjuV8NfesmN3ZZaVRBWPdJgnvSBFjrfsiwvF
cVNHEnqnakame3fUh4blKGSyPhJQ8kH8GzpGAwhPBHwZ8l2100eMDDb8nCYrrLhS
IcCNu7nLOHpcOvocWaoMRpBricRtxkp4HkInWkwVtUi8kVxbTlIW5O7U0IXvaRL2
xZmpDEiKKAjnJ6SibjI9PHbnDr1SpRDe3K+OPVdim8EJt34Z8ghgln/OvXRRmVrU
DNSIuwcsPwE5fuJbHxNi5NlD1wSqzeP7xsJ3kj77jRv8xmbUr88qsgfkX5jh8AQ7
78xRTZK1WDnALkWUXlQZk+aWXGKd0CW1/hNgyE+0zTR15BzppuA3dYX4BJEbxVYP
fIy7geTez4dL9hhX89WTLfRm5fTqQF9U+OUEX6NVRqGV7izc5PTTstOSFj41a9P4
4DQ8qh2h16DWDRg5g50lO+CQFi2VC5HfpXZf8rLBlaM6bUIcJOyb1u9W0UcLdmDL
Uq1RYxDUVUU7koVumMMeFrOa1aFqhaa6Nh3DId0XlFRlYi4tU9evODXObN1xAG8x
2Qh7lrLicdN/51pT1sSnVYUa5lQ4+NaCvrObVOT24ajTxCNPbw8M/n0eNHKhQeC/
EMJMKnYM1tHqVITrxzN1sOqhjJZSLnrLicMsZ05b12NdnHqkH50rOjRhJJjO95/L
knj47cFG02PZHuxgg2fUyfGK8D6dtZi+fkOarw8+tmhCpk7nhFyL7zBTgfPpqrmc
ccMZ+wKwJrR+2huQVrPyEm2F7Su7JTlI0KlJx1TmvPz0sRnlUVaAbRFPEj2HCCdF
eCwRnuF69Xjyjp/uMNnz9pzcJax2rSl50j+UHJlHHFFsh3uh4VwYyIFHcfVaPRvq
zkjqIdVA7Ya2csSQ4r30i928FSi4+izjrXXYZA7jpxZiSNuIbU5WgLODsMNTTYFh
CV1yOzTrcPoTMDkMgioVcZhi4smKxwg1Ox/kznMN13ij79KaQ1EOxA3M9J7hDFzM
Zv9pFMrJbIa1n6MCWVcpDxdyxkT3Xvzt4CIQwYdxNq/kiepZq+o/P8jZhs004VCN
wcPPCIpQWqQ6hTjfppwNEMe5F8J1guFbRE64ndrU/qFPsT43mtzJV7NX1hgwYzdE
zQfJz8F55ncE1qaf5pHZ0a5bqaTHP5iA7ulMDG4HAIx8wo4s0Igykyq/89KJ5DAr
jrPuCDFmK4BS9w5qdY142mTX16e8RrnhjzZe9Z/4BTFvopw4oxg1yHI87BDo1cXj
puWprGP8gcvrErb+Pgs/d7pIAUwP/gsCYtSxvIOxtmgldj0TON1eUZbPAxWUD5r+
03dnr99dkZ7u7d3iBLjCJDwmCdnBX3RRO2+YVoAQSylFJchXDcGFmexDSwAWuUe8
nllsOXa6RQNrJs1D1u0YzGHwYWmALtZUSLs4Cm39DhxsNE4BbXNytYod1Bb1dLyJ
dXUxG0VVOCONKxPTg9i2gNtlaQqQPjG6x5PXADexp9iIdqMpaOlpyyinbpDkOL5J
aNvscmfnEhVhBDNfORniSw9PEXDWEjvQjXyeaX+UWcOlaaXZ68LcMC7Caj+07aGT
6CxTHecSAzPNwiA+pkC6gLF22xiQOg/Nf1YwxuarNzizlSoYBuvcZ4JX8knph+sc
W28nAuIb9W1y180fzoWGEPbBMcOVBeChltqChcsWpc0mmOx5esl1m/h5dWhkpEEB
NnGL7c1415AqWjqSSsfH4Wy/UvTcrR02R+DAS/Mkd9L84ZpROvOTPAHZKGCzhLYl
5VJKQ9iUYkpcWRnD51wNOm4pIx+4zY2WeBii/HoT8b+TcHz3M6Yudkt30fCFO354
6Rskm1H5lJaYgS+1iU65O+Yih+AUqtWdlStFvML3twfjS4yvYlqPtK5RHAuSRrSL
D/+Jge5jnvV5jgf8BxoldR8P7MbUMSoEy16vQyHUNwGSRU9jUfXoj7YUDP1hP092
TY+lkbNCJmnu0JsQeVMRwNY3uAAlRdvOJIrSQLaxVSoHk2uzeYPVOQEF8LrLqTuI
Pl+XYGj0dLhaCwgWTnYdWWTs9lyAuXrk88aOseytjy5M0nFJLKhYWn5PiDbDKGw/
7rHzW3wrvv0crhyJba66HQ7GSnRNm2KGmZPV7tZtNCqHqpZCCa/5o8LXyJPqeKyc
gTFyFl1ct2w1IaLK0IjDCVnrmzmvTLqtJo9dC6He4GTb3ReFqKRzN3Ebo/gUbrca
vljJZksOFD1fOp8gM3uoxpTXeq19uSuqKU8LCZLfAuPsyOC7NAH1Taek4tVUJ7mP
A1kb3KO35IOKVkzGysvRdybbVFa+9tLI+iifBn2RglMbPwu4yYpa04V+BXWvfRxw
GFiV51jEEd+5J4/X6UH3bzLVHGu7UnG1VU3sIrxVGLiWmIrtgAw6bW2Xj82bDCC7
ENAj1Y+PzwfAA4t7HliGNuYClt4O3zz+rrdbLpn9rH5GGdGOYEgUXfy+Z2Sd6sAP
tMVx4oa3Bv8hj6CTlqyCtK4E8F7eCodKK2G4B0v8v34rGf7lk/SBRJQSLhc8lfhu
wHZSajgr6LowAsZS4WORGVjlMdht+5764KuTRq4N2h27CX2zsCMLJwzqz8wb3cAh
1yZua1+OOSLnNV1xCokVBNHzG3TGHCzZoHBXyoAxwOGiTdJl5i6/H65q5C1D/V5t
eESdQp0s8BmLEFhO9oSafJPVtKw5ygw2dX/L0Yjyb4RRP2WiwZ4Zx/L6ldheQgq2
OLES24zFakzHImYhILnqwDV5YIZka5E0NKsaokQm8K6uBujmNm9uJZ18QbQLi+Gn
5t+lhk8gPrs1SCb3VUkO1og7So2OwAnjh521xnVgXuxoR/viP9y1xWOtF4kn/uLx
IfmIhECz+lIgAMvWyH13H4ifD1BwoY5467QnDaE68DKVQr5xScWjIXrIX86er/wU
j3QmIFjKHlzys51mciiZFPoKqTDaudRFHc/q7oqiYduxBFUHN68cYS67GJapEei9
OuIjStr5KJOSpVl5uXFDwcwO0XvdDSEh3IQPY8gZ3AuAJlJwyDKu9oPgzVvmrYRm
br/Q+BsFYYen9EmH3bYpBFXBdmdf9c8WswhXtFa1ml+RcnHUMcIXLTtTNwKWBRup
XEKEoreH08npfN02mN0KC4ioRTymg3PGOz3QtVcmLTIeWsCoIwj/MuJEok1mi6Rn
SKCi2IeqeB7czF5YSISkhieXrwWdQ+bZEq6zdW0lKAiNSyIxzidxgpAQptEuf6+P
2SaRbFHdxCWg+DtjweWK/WIuTdWJWLbfPYdzsiErRf9Z/oPqyzlS6TaEXifK+IRa
2atxeQrLSvBzdVb9OX18PXecY20FHd7hWzbwgm4pFZfe2BKQSH8aT+0v3R4guHyM
CCznGaBL7n0U3ReUlNaEYPW81R2LfA/zGpxMl7gt0C7ep58dyobTgFaHgdrVLAYh
9HzfMrtLtQQlBAPanL70G6aydN9JBHHS3fA7ICHS2pyyNg+gbUI6aXg1Ir6mf8Fw
4Yeu5gfedCknf4bXeFbBXfgFfM1AMgZCy9xHniPVcllfTz8WQDmyiPUfT0DVOKAZ
YT6mmlarS6f322jtKWZ9BwOoQRf7WON6F5sWyW8HjegiuzErH51AXt5Sv8o+a58F
AFA2gVRalTqu5pIjfU1mjghX8Ye/dGygJ+LAzbhQ3gRFnc7gUbyuSRTMeiB1XcDE
hfb10r4II6nEWLTLMbqQVfUJ+z4FBeUw+yhETeB3AQCdcL1gqWzxRciHpLCGzY9w
blLR/TZNmhwwAc8K6Xbe9XD1ZRHO/8DhCGZKD+xnAoZFrJyzQjRCcjlDu3M3znKg
+a4etra8oEDIyJDuZaj81JH7n3gK7oB85MwvG59IvSE/KFSqR6Q2jyv+FlZ+VfDd
Bhfa2SZOkHbLNDtSt8Sn+Oa/jC9VvfJ+cIclTPz/DQTD2iDKNmCmcBJB+Y4+fyYs
8tAHUZVry2zKnGYQVg4xjtUpKNYgiiw1pRCFyTozsPVQWLjPsUwQnIsEaKp7lmBq
dPIVX4B/UlY5zcT8noXq90iVatAnR9W1X/VQWu9x4YblTc/ZbgWbXhs05IthI8xx
B6mUQ28ub+qEy/MZjP+psQnAaiirgyo03E3+nVq43+QNnlskQADFAd6ga2ph7YIa
JFJze79wSveF8NGuO3JkaTX8GVJwP6n4z1UEAnzNrOiOmjdwOJJeVJlA9RMC7ulb
eLKo6qnMmHicPNCRRugPxfDdwvezXjdRouYHYjaPDRXa9hF/i4mEIZ+6YO7GD8s/
IqBHO5mIBu3aFGKGWpC6BC6EYYHuTUWTP3iDajgv5yJ2F330J2qClIPxvlKq6HTs
Ti5f+HJLKgsy3yYTR7999cxVCfMl5oqBeNJRaNrekgk2t/uhS3BZvSIHJgWlXAb9
gGrd+BYiMusp17y0CsxUNYhKK4+/dQcrgZUGhKrtopy8/CPcHbALxdab47DziJWW
ray0CoWxhYDU7xKB8YNNJJ/HAte1F5paFurXX6Y77BekfQGYlGk+vBe0KiXk8aqv
S7hwU75OXHjfJvBPLyEovdb0awTJeGiqu9y6L9n/AGA3RYKInNfS2HY/cduSLDSz
zu6VzKbtQA8l5+X1ZviGb8NZEHpty7ppye9wFHtXu/nq/D6QuxCsxgTP36l3wTCt
Y22ETcTDRfXtoL0is+k1TLuOCY+dbmQBvDd9tRKKFv1lQxios6KAxSOwrADQZPdI
P95PE0Ee2thcfIl1OQ34JHTkks2BsZ53kM/nlKX6ME56lTgQwVpnLRssePuPEHYf
LHc6LkYmB9E3M16A39TyPjqh2VQgnVb4WQSIs5gdegruLxGWU4VMaROQcDQNV7vQ
hxo2v8LeYCXNS2tUyfsEYla0ciiuvsMUNm5HdS0zPDfAKUxutArxJ7UYF8v8fnZ9
2CnmZOcHxo4UesjPasNUx/GymmfBBHRhfbtCKEdWOsUYxfYmUG5cfrntGpo28t1i
Qp1l+GOfPu9JhQvne5qDeejrKjdeuStqFzNUAgFAsY5j7bq3YMg613qEO3xfVBPd
C2KsGuTRDRl+1PQ30YpFoeVsFKc69LmllNC8PCN0x6XZP5Mi06mJPSf0icIm34MI
/10egGwC1zLz9CQVuWVAClOOtvpoCje9u0MgsNvW3/bqkzGbJXl0JVCDBhcQeXxF
E/8dvDjwgIP74Ux8YijF8JamUdsBA+8CmEE63YxPgN8dQMFoXAVI0jO6SUCZ+VXW
G0sfGQ2ekYJLrQZWJoDsW5wPCfze7KWKUcU95VnUvSDe9VHxsqoL8lCI1X8KraRU
P2KarcgyEuUWNckXK4yezXomeWvtf3/dX9MjsGT9K5Z9bhmXaNQXwFPZfmHPcSoP
TVtANPo1IHMST30f+uM/pTNJBzkAWweNGyvtrkM2LpsoIjFVdUPVuWMHZZq+0CmM
OhJTqGGfM9DSuja9Exl6+5Ao6P857XrmXP99jLQxapkZq0PVPUJW7gWlIVlAdePJ
mlJF2yANp/yAW1y/GHX7P8DUUoO2Es3WyF47Ml9FLDq6BVshWSWp8Y3k+8L1oko8
EBwmfe4WwIezwE+R/WFjTWRE9BTcimE8yvw6Nz38dK2pGlHd06ZsZqTBg7zm/tgY
9GL8zNU82b9GWlsepDcMS5dbCYpiNps7XAYkv+O1ffbY2+ZtsU4qv13/p63l1De4
cD2Rs4d8kH8feDFb/lnKEKrv8wjpeyhEkhJSlbtcgjcu4FOGWcePQxbXu9rCE/El
C5JfbT8P3voLbVhR5z9tIrDzO1+k/xkOFszJJ2VldlqpsCTh6m07RjxrJZkO67we
qtwlWkyyoXnx5BNXeMoMWKofGZznfnIXYMi9DsIa3tWyYbwHr76OfYD4RrcLgZV0
CN5fHcne3rwIuzKwsna+jTiO+66iBXZ++FeoTsoW70K7go7O4KMRUrNBUoIDMg8P
dfEWxBCkWQmA0gnpq5w5qfA4w+i+5Rb5ua+VI310Hf4sw3Bzv0X1tHzgMYiqVY25
4qhZYyqL8KBwU4b+jP4UAVfBJ+eHtUW65vJQmSnLFJx4vUly1Jg7DWSly/QIbDBn
/tazE71MvUDs54M3jq0NFTcYI+ZSSl3iz9jwCANbmBS2mxEH5ut0xnwqmTN7XNQX
0HDBozLqUUHrYo+VjNkqFJ3ZOt1TtxTMxpVZ7Tuwli+Pd/ZRM86C2GdQd+7BmNCg
jzJFOOssQBBkrNmfh6bsMY9TEEA2GJBI11QA3tUuZDW+fl/EsdWchNwIS/dcyaNP
LaGrUyVYPQ4ZoAnsadqbCknlEUtvYU+sSn4GmJiK6ux5Eo/qUsqWXMmKncJ4ofKc
MW/4mSuiprRXikWa+guN3CDp8z7QB5/KuFN8rICP88tQLEYumIymV1OEiFDy36U1
6rfEj6LAQGsRwZ7+I2xqYfk+ZTqseuiIc9ixNs0Yh5npaFqJtxd/kBwgJ0IsMAbM
4YBiRmE7dU5AapYpLgoFNI966RJ4STiu7MBo3IPKL0KT/UAp5qRWdXA2BzwlaoDM
R3Bjzw858pBPb/ZNzFGoVH99zpAJpyPEhkUPr6yCQOS6UwxpSBvApCtWARPTETc3
gFjwZ0ECd6nbnJaaytba8LQm+e1SHFtp3Qcj8fA6TnO1ADLKYy6/UQHA8aCIS/es
fWm8yMlJAjTDC1QdR9tRBx54kyF/JlIr1FpcXNGSDTI/ud9i9v7fBRQTUfjv3CFl
UILc9TvvaRGf/q7PmM0/BZA0dlYwCRc11iRUEFhwi56moyaeCc0O1T2ij0CsPbl3
0pBErLwWLTwyLce3d+ylsfCp6ey/jT6Q5joqJyhYL2xxYk9buqe4oTebEfydDNO4
8Oc4bIOI+/w66FLmLFj3yQMbWvGO/QRms75jrFpNUAWNweAk01aNZaTos6+svtCZ
Fd0udMJadBAQ9Ojly6Q0uNVqEPCLfpdYMluCTLsb8p1lZbwUmJYIot2M14eKZXqA
Tsym+zy7jdqoDi3hz4bFpaDWBoRQsPOWQe9SVUsChACVEL0pZSOkrqMHbMM0RFYu
nRtcX5+z8nCmzb1g8X6sQ4mL5OLvAIS3ETfyXARhZdP5wg+/HzYsGIEdj7ELyeX/
A7hn65NH8nTudjqpjJuK6ADGWNUZkK2x9BMG1iLzYSM9X8xv6Czap8zYJVS+Faox
VGwEFQ93fkx476zBxGRhSMMagzRC27R/PjTl9T4cWdRkL97HkuPVDEh3Msa89/vr
pj+kAsvmavrGc0AGJQz5h/DOa3pNCOMel4DRdqzL3gU3bPQx/L/Bi8VXCiPc44bw
fD21Jaf/Gfg9914B+LFZ/nB9taHFrLpAAvb118InSw/LRNONy1iqZXMeuGB6Q8e5
igfzEV2GrGBK/U8nFH7ygBQiTB3YznsJnufPoqZQ++DEh3nWP6StBZp0HyScIWOo
j4YpYbsAYdXbsj5tcVqEqA4G5Ph12j2KGuJNVAw6K2M2HKLqDyrPjG1VJlJDQFbJ
yQZt+DbtQnxLVfyARPd5q7JrXekRYYzFC1XpaR/XQBbKJWF5UqHGLWgc0cDLpjSA
Og2BucEGqDcW9GrE/A5Y304w3ZZvZuQNU+w5Bp0tYHp+bZmcGfVbR5X0AHM/aHLd
8oFfSkhSnCdnWF1eymzfr1D/GqsIiPhyd79c6tl5vI6gelP8HtrFHljyr1B/X2b3
dGzvdlaNa3XV+FPeGwTt5koCIPv2Ocr/yy+i1ujwqE760C3fiM2FfeUrt5X9PhLB
nUYQ99ltbtKVOEfU+OiWd2Jw9KMcSyPWWNIsG2nlrZSORbTnvfyCebVu8DM28vCn
3tcmzwChRu2JojqMh+jjnh57DVif/TjmMkS5cJrcgum7Q65Ge08QCCREOwgc6q3s
4naxI2g4Qk8IgkJcXsQ6SZhg7SrTMaZtwUNogXl8fkvtJ2J85mpGpBcdkL3T6D7Y
pRpUi7XI0UB45GgbbY1xkgfZF0pN+gPSQwRUyNjz7b03gVVOlTQVdH4ulFGzbhkp
UMcweVchgi1DvLZ5jS8r/hupb1kbVpaRC2hnSD4o/tdaBmY+m2H6BEDI6ghpKXeo
yCJpqUMk9HWXweaa45aArd16f2qsZ/c39Vhr+4Q3i0AyYQbSUWmMvabDAGJ3pJ0H
fGo6Gt18T/qj/VoD6dUIOpjGGipNiQvx40eKvsz1a25lTVfyXZZzqW3eFFGUXQMK
WmqolN2x7T6Zcol/pA1HsmkFxjHWEC8egu+IGZSF0ZEfC2hlrd9RCNYnfKoHBTXd
ydFZhzRVHvi/KH/LSOYeXj9LF/8k0zbHrHE/mlZjdntGD0oNwQIwiYa28cf3B9I4
x+B/QfOHFCAIqNEEGHrOhg3eGf+rvXaMSACMNOeVidpYji9iUY48SGUlTpM7bKca
a4YYFo+1tQUB62sgqW2Q78r8/1LblqgP5wnIzKrrFrdlW3Cp9XYmUTRYg0zSkJeN
N4rooxng2l+HAo4o0qrqxOqJbRS7GrNcgHENgTMgG81kywfPjaPbCfQ8MfUyfZy0
o9ggmKCn/eCTWCIdWSeWiTWUJCbt1lNXLILeqgcFfy/eaEdNIIMbR7SSZv0rW475
6ZNGYnmBYyAdVQVgLWDG2pdcfLXdPXbEiD9bgINEhCu47W6sWtDMUvIW5qu1qkJI
MnbzxQ8zwNJn3/fRBZVWGIeH9M5Pf7qdYadRGZmbZOPqsnIvJiSDveoOEt+fD+lj
B3gcgnzfegBOQCHtFWEsqzO0gyqXrJglt4bRzKEaPgTVdQEYVZ6jJBp6PfYJ5kWV
rGA3MTKZnojtVu9LS1BDqgRlVPBxuaP1CPvRChwTAyJmFObbKMkWh1G48XqqnldJ
MboEtkl5nrPfYEOerNIpLi5jQfPMJgqYVzmNfelE/CTmvywrdnkO1ufFRU7sRYlo
qpMNWZWZ4h6AiX2M+oX2GW3bLbVrOOQxybXTQDkaig6gBzDE/hSAmH51bmcd3sJW
XlRc/iOAcq1qElPL/Tgx5muGoRrYXrXzQX+fSWVHVKIJ5PpUlLZzj/tN/4HyVzU1
szL3WAOzkNHHy8Q+vTl/XmOVZidvrz79wqYL1bEKzgiEuW6vKEBxSQ5c7f+XFdkV
pFuLAXdFb5zQ/szEpcUD57k6Ak70X+HxAYjo3M5bJCvoNIx2ZT8hYbJmOhL8OPNG
kcRPWpfFsQscKl4/3d9FgMYy5dWyaSOrK3Du9n6sI9OMlKTCqws4p5aKhu4EEDl+
LEdUwF6QaziaURK1Q74hUkc8k649AW3+CoX/TC5CaTSNWjVVNcG7Z63l0e/dqBR8
hlcjVHEwTWk0ugplAJytTfjo3hbd6/T1rUAMISozk0MAW4HqQVWrItHmoF4aUMKl
WuvJhmEZiiwY72Ay0W1lmnKeTrBEJ2h9FW9ch1TfNRTweBw87kazLdGLP5nLcExj
xXJVSio4oYtkPW8UJn1u+CTAV0zfv/2+5qsnXKz1WJVr26NKkl+t9to6McGr1DpW
C5oJpBt82qb3Pu3jOE5NnZuFaSetpIgKvWKwDVnsnHh8fIkJ0+mVH60EKtsFu3ty
8eEoAqQhqvkYahwbtglnvgfczCIvmwDrH7tZqk58zoC4cM0GiMzzhm8GBYoRtKue
7Y/c4JUrCecFXQU1uaN1swkFF8iyjjABLRG5P9RCFxr5wUGs9toF1WJ7rjz7fMlV
tVTs1OSn6bxd/827SF9wBoO+c2VRZl8XJYqQ5zFKLC66keFCnczPgIixSVDhRvS6
SfBwdqOZxmdQ+fUDvmMVSuk4HcZZmfK9VVOSJ+V3gfDwMKUhXtER2hTAvsiw4zqb
lofvKxOqe3yvRIgdp3vJjcDpsABQQUmbZ0+TEv1LA0rRCQkQYzDlb/ZbSyQmMSyd
wt4RGcUc6pWXI2qQ+kxLFSkopa/DV1XSgNKJ4GRcli/W/Wvkm4Wf73TcPFS4gpIX
7sfQF5PDx1JOV4aGdKt++otueaBr+c4ill2f9ODNSPYhA+6WGSQCSrS9ja1RU8X1
UwuTk++hJ+Gf2nh/tHTPCnPuoglcPii1wh+AX1e0/QQT/mff9fmWnkBG4yC7Qxwg
bgtci///cI25xbTgZGPk+Qr9dbH1TuiXU5yYbXnDJHaHy79lTgavFURJNPLnVQ5c
zVaoK0AZFe7nZlXOHr1r/vBCbDvBrQcr7yHJrEV/ID58drHXzheZF4g0BoCV8Gjj
FX+pP4z8DO31dr9qdTKxOjkZKC4DMw2H9nTB8EuxuPjgF83weoyOfOJ6a64X2i1v
kTBrU81E/tQCNru6QmH3hlkc6SlFhZyw4aPpRrzpr7ICnl3gL/WQFPJK3V8DsF5z
8nurHt5FST+dx5Ig6JVS/H4ZcVdQr2uWAYTTiw1fnWL24bQZ9BX19UubAgDIpqnz
a68MY5/4hf440nWGZAuTM6lMe8KoVxG6jikFsv/tCikLSapArnokyB0J0e2g0SBR
OAxIC9nnaDHnpIglVxFAqscwGYMaMBILlaAVWsxM5+BJ9TYcUCs4dSCcAFJwWX77
IBI/ZiOm/rnirmcKpkRPcf3TzBZZZfgb5ufL9TlE3ImTtFP6MOuo/BtMBxoVSc17
vGyl2wjwjqF8M1QlzRxpTmvmNhWWYFwcsdsoNa9X2rFu/5q6JPRbHZHJFEAaxNHN
vN382AEp8EfAvriVXFUGc9nE6OY9gb464i1saDvmvj/Fcm3liPzBf9qrPcmtRURQ
k7gKMOrhifpoKOtho854NOOO5MRdvxDpi7q1msj1N/xWrNEqr+Mx1B+SBz/cbHrO
mZBdmCPP0NIBxdaRxIKIR39csW/nCYGJt0ZfAzcdvIeLlC3wDk4ijMWIxafLrMSI
0mS5yv3dE1EaNnHnub0bJzNnG/9+0ud9UbpD1HOdou6jRLR9hxyKuekajMGQCiOU
diW420VWgOwqGDf46P4e9mQandQ/4IgRmfuzY8tW0HHog4Sht4u4s9DlMc0a+Fal
uXk1syH58Lo1pJHTP0kr0881TiPsQyuoUoLlEDXt4iCQPfoQzgu0haKmGTAng4RN
kNld7tYj9lX1UuZ0zDv2p3QgROJFD9FsNKVY5znxS3oFaNd5pD8MqlAVFF2+YG2f
xXQ8h8e6aKJxGn3pPenxMnycWgFQwXcZ88EJ2DAJPRy8yxpwdwjoPKTSv/bFhGT1
WIymZDu3FNt4cEihJWKLlmHBFb9XT04MlPuPehxvHTRWDTDUCgyJhLSnLc//5a5z
xybUfOavHQvQrA5hyRjBbJ2PLXpUL1tu9BomvzzsAuVPikZeHlNLrX6V7RyPC0Nm
4FplXgkmyV5SMytEfpbwtyk+PMxChNtoKzE06CBCf6u7/xLIvwVRUBnfyL0/duHF
ynaUd/nTAW1RqyXgBtZpGAtgIiQijxMRIgWsqTJ69TyBSsc2thFNtXcbVSBFzjQN
yaUKaj+w7cenBgImJGY0X75LyC7yaV+NLJ79bGjogBzVikPOcTAv1VDOOIE4fOYb
nqn4VFLWU3UieuArTtLiAKzC3RufbAooZflnhR0xhjvtDs9BixZR8mrVCehGJGvz
o5VnIgcjfFzPn4bwkEXhq+dHNUOn4hnjHCG66dniRE9O/kWCkzMOkAnh6FsY6BkA
Xapn6XFJofONmR3KfJcRzrZPs6RlmzxArfj/oiDcJq14UOu5BQbdGI8iDxz22Ha1
vT4hYQnbB+OMN0fPm4808cgXvdwDms3mmMD90JDdj3HWqvyjNO0+Z9HsBsQKwsAt
ayOVsy8gtinWBMV6OSS3qoSyooY+qh5/mT1H6NFyCqK5IRS57yAhZx5abpoCL4M2
aX4UdKPZDLCZKkuZx1Y+aUezKfHUSQOinX2vejkW/YDeKQIcBG3a2ogCi6FDQ776
rORNuC1okxfjJUlXdE0Hj78quPWGwUeUgzSUMajObyHB7caeIzgjlidq0W8q1Zlb
BY6Y5Ay43BHCg5bL2RCDDbOWc/r8/femmXaI8EtzMv2lFHSumFs0AR80AEh7BZvI
yOEVFDKKjfJWAvbWUwOP0V+uzqKwb6L1/UsaVvnOvPex/EBHaqLV2b9szbCzhoTW
08wlxUjDSPlj+n2b415bohpMD379QViAyuvyuyH9DgtNBoUXWB8RKrAtXG62POXU
R2bb/ofDyKtYz2xI3mFRWTc8UjNW2BmNSO5hjaqCicRXf5LnSRJmUkJ5ZZv+sPOn
yEUY0ZFMoX7GltXQGYxXGeqV4xq5Bnk83jisgFgWGzgi8Qt/XvNw0uc4I0Up6e7a
0iMHZJSWf6gwqM652LuFOahMUigF9r9Xetg27uo17j+jFjgCchSuBkRITzcI5877
t+6LEgMHIcuBCghQGUorrO4V2fC/a0SG0lltOPgWn9v9oHOCSVoqSKPcm7zlm/2w
NvbVC12G+Nq3w+Y16RE+NTAiYvAxhskQKmoMJ1ItchHtum4T271m9mgl4ZzS34Y1
IAeomVgh5YHsSoHVW+t5YDoCwkVKcjUIpwlf2FluGX2Ve25z+BBSNUhAUlvDG2CD
47PRH5Gp4J8oj443Ag7phAMn2pJ+08k+pF6FQ0L36nEJOCKB1YydKD9sThXDJJPm
eaHMM0XFmw0CnXl+pHz1tc5wSglxwu+Fdf/ik8T/L9voXQkERr6QSI7GN3lqFRc1
Yu3ZAJiuoH+ZOYYg7GpTlaJ4+T6arK2NPB43PslVn5AmZpooy46OdA1wy9wBhTAQ
34DOl6dRVoGeEbXoVkR9A/0pq2amnsq/Wik2A+5uOlAVY+b52gPqtjd+Lin9lp9I
Tm6SjxvfggOo+ESEdu/H3pbfNRLawkqBegiLq8pB2XgCI9zUgUYtc5WaIi1TRObx
K6M84UosbkYVj4X267ugvp90jy7we+s7eaD/JvB10Qs8wrJ55t3LDPieERS0/9om
VnzWokz5Hl5Yo+NntNRysPdRHlGvjXkxslyBC67iY9ptugQi0ygSfydvwrD92Ta2
dd9uJM2HFRpL4+IGsrkI9HYy5qnPS/gi6ytzFBLGxjY=
`protect END_PROTECTED
