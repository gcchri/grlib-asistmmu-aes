`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6yd/V6uFviDRCvgIoO5qimJAHCVKelpR1rxz+g0dqPWhwnXVj5mwJTjOKF8pyYq
sWvBOz1M5gbRs/6iID/T9uVibJY2X4yud+kBTBB0AklFcGkyfr9KqV0L//tzJFjh
2EadrZ/Pv6HzFAv0tR3hjlVNkOaZ+QAcl/mclJw1j5GC6wOkLfdif2NFPq/xf2SH
s8tNOebB+Im8hsebcY/8jJJ0R8/ksCJ3SF8fMA0OgaA81NifJgnKtVf+HSCmbhhc
4V4vSWFh3dDiBlEURq9eFhnXGlLFeEIqr4QZ+OgcYH3NT/4enpk8qALzx4GgqvLn
xVG9f94IgqhN4uRZl/UrmgbaQfnLy5fuIsZ6vn6Y5gcrUiwNBx4GLGtIDVmhhovZ
wWWhHcux0fs6YGZ4nIlPSk+mQ8gShYqYCoTLREnVspi4o6kI8X5WZuyAYGRkd3dD
RLXjfREoe7SMyK1hRedXETSJPljJ0/6F1h5bqtGleVbtE35TA0C6dQc12sINj1Id
aKsNLANJ7VmnwicQ0rjleEyPi/yiozsh+QZn0HXy2Fe1TV1B6sxna87OzclWWE7C
eTxBQJ7W2HK4SbP862Fc0sfYI9ddHZM9yOCFcUpbq3Bhf1zh6Tg7yY6Ng8y7/9x9
mjNclBwjVb+dsn/Fg7nYL5Lz3x7YtwILNnCNKv2qIjYQhNE+CF1QFC4p413YU6wo
2WcFWhTkklzAzhyglS47fmb00NZHfC32rZesLQQkJ709OoR2q8FGK/N2/9oOQ4cI
OTyVdxVJL9SCRkj1cr8V+SzpCE4Y0pKfgiHR9/Y2gevdnAHxJSg0HX7x3ofdrRI2
2ZYV9FcmmldSKoDaw9XbmPJ2HUQWKAWiwiw5l50P5xgDIJb/6Yk5xGwY213/S7tB
ea2hd58Ex3mQmpiY7JAjhv7ViiOSC3KAfdY05rd9W9oq1aPyx3W6/nZI9DQQThpA
9MWxBC7n0Tkn4JfrMxMhCWJJnZCvCxm6CM6T6VUu62J+/BkWYOWYBIkPAgh/E4PX
sdpJ+EkETZqcpOCWMEOLl9frcAEFTkZ797L8CN5atyTa+YQNP6tYFfCKGTK7Mav4
4fCY8oy3XMFg3zg28BS5vNhagtGCnrXsiC6VV77lUoIDaWB9MU1Js9DXTiE901Qw
dSYeW/FEUWVhP4WZa8SRNmtWDtGP74c8p648ey8TMrSxL9I1KHluOImD/VdlxS7I
XdZDIGQkanx/mrmiwAPgpjOjJMW1Gnt0Lmm6VmOCNh+rT1PptrvwncHlY1gftn4s
rt8DdBzAvC5AcSYFv8VX/MQBLbBmWNIvwD9rpgjXL3FRMkF/mnB9C0jxjnemc+JH
3hVQfke18LgRsxTxFAP8XlyoVKRl0aZ8wpdr3nVf566AtycfsGZVaqx7fNKOhR75
4d0iE7VnyM3NhHFE75ODVnZGDLyX/vmob9GmhncQmyJpLs8xDRExejmbBW4GzOZ0
EBO7G5qc5ozWpMeHz01TQK1nIe+3VtIJRQenjbZTs8IAfG/NCtxGhAwu92JZqecb
iloPicAW3x2WZVP+23MFEAGAzxCMAb6Hf5SsfdlT3nANvENGo8gnuUxsypznpi6q
zAVXEnUs71J5fbzSCKbSuAVftqnodCZnHQNb6rg+g5LbWWzQ3QPiIo7lEKS0DuF2
K9idpAX/d0FCqg9UyV+xf4RfZ8+T1DlP47UNkV+izrXSpSuEeAjTH8vKCYdU2X2R
0a2pzMx9aVBDkoxaUfnejY2DyXQl2dlq17u71zxmZKoDHtxqRIde1Z/o+DxupZfm
6HVvREXI2jLUm7DMBPGS651wAr9Qq0FwET4+SErZERcCjIobunnL3KE9c6Pk+8Pr
z/GShhcQ+xRs5LIDlzyxyfRxFTJ5RLhEszWu3VqF366r+x0gmm7HO2wxj48nGUuB
iH2cFVmY45jV6Ao3VdpoUSBCRsCG4F+Wj8pvByHySkddCdhRttq1QMQ+uIX/Xtu0
uJkJRdioAbpCW5y92dIJRq67Lmc2xzh6cyjt+RDW3oVRdW6fvDaPYnd3xbb+DA9F
m4NlSoPxhgoquQ71llZFu3N+m9JC+u/MBaPCSL/M8fDiWFODFfjLu93sBirTF+Cg
0kiLvUOaZSrOgbfwG6Gz/EjFV4f+6RHZWTSv68aqs7GB8Z7fCd//NTAuWU49N6Ig
H2Hx0lZq+6Y0ljINagqVoIPvVbnTTL4xikQrWvS7vMsfywPwjkOkGjCYXJtBgU4x
j6lnS0KB/VEEvmj3EcLDS50vtl3RbM0awE//NwM+e2f+px/ZO0bK7IKMFYmjOq49
ZWRVelI5iQG9LAt0w9V9RlDRJADUHuCeEh0ypf5rPVd1a2oaRQxw3tblSzuTYZA6
C53ZuuJ0VwUZbqBj+y231pupbeqr9jgAvbOBHnRSNeBG/vOByObLs6c6/zwIneON
M7dOu26JGw8cHMW948F7JOQVQ7V1Rww6syJ71U+beLvIdZnZXcit2SMCZcNH/77K
xl7+X68O/jcmEptBX3eiKljRYlljISXuARyO4EdQ9JOg2e+0fo72pT3P5OqPwyD8
KExkjeV6TPwadf2V5G1ci/FpwypMFMwET3yYTAPA/ku3vbB+4v5g48pE69kUV+VW
ISr9JZxnLUabVi2uMA/xrO67D1lEbW82PLL6QbQFegVo7nms+lhwQpchkWm4IrAe
zW28wOUQ4xZkuA7nXJ17mF45BWS9PKi70q0q87XYiHOmVQBZl4cOG6gE5wYkEjZ2
NW6Y6jK65z5jzSZKAAFcoGSdzSEA2Ll+blck2QnZe1R7TG8jPg09QYiTp9J6aXZ9
8ipZVvMHf6/i0fbbc1lGRpyROiXZFz7Pl0UMfxnl1kzz2QPm6KENX2YRX6HNKFDw
Bs8yL/UMkAzL+2PgCRfiEH2Fv4DDeahr6NP0AE0g4LCMDCij0G6JItDUt5d9bhUr
/OcfqWevUnYxPsGAcFqAPTybi7eowMHcxpE6bMsWP5VZsMdUhYO1Gj5oyTv86+Ez
bLoVlTIx0j0/BZAT9ZE3rryMYSODlpBmPRKuFHcgU0uB0eyoM9JxNVKLGCEvn0dM
8NTCfna+t7YCPtl3beTUz59b6xOAWuj+amQBXXLcnCPKJoRxySfrlqr1wWDSbYOV
nJLLiI6MlAxvZinrysy/46c6xemC9l+b3icVNy/1gqQKnrt65J/YcAMWAtJvPYh0
aNGYNac2AczAFrS1BSsjgejCauUHT3SZiTJA224qVKAjopmF7JIWhynoPuuSvZcE
JY+RfVz2RNYylwE1XO1IDDaoY85zKxaopsV0VhcZz8vviJihYmP7dPz8f7VqHxly
wMOgmeITobpvPoStNYBwd3Sfz4slNhJWpDRpygBoXz5ThVSrMoq7b2dQWDrn63s+
D+KilyMs16G0JWRqhArqslHUm9bQLWGFH+XHz3SYUoCG0fjXtF9kbTeHcYLHVA8M
aaMBpSBJjzWlHw9vugkLOriElLJDiyKmlSWC6WgeSaKJSrszLUPBxDERyS5Cig0z
+Bv4WikSJBcT9t4R0nYzuNB4wDDHurTdE0215Peq/x8Jt2zNXRRu9w+vYIfkL5KN
TMfyXpt66awHcS1wKXpT69kqYm9UVABOa6ec/71vQedoZCcS0qyIrVbazu4aDtX4
dqDcwdoTW9nx111dP3f+slVs2xr8XwvFFySMpi2Qff/fup+NxQVuSS5zgK2o6xmh
sJ+CXKSLwJi1f1hKM56nkjN0EORbZoh/IL8SFTFRpS7E67gdy3n5F6NJpPGGIWEs
dR6zJm1taRx0k6vjZWTWN3G3/E+ctN1WDCK5AMihWVIqe1XVV7yqWs+TPvBsIlIp
teaB4RMwn3aTF6Nq9WA5XH3yEpFb0NNvTQnWEcILXtt05P7UmFpoBC9feJG7ufw5
pOy/zmeLmyurv+/3Ef4TlmtwM+e9AoW0vaW4xS56VC0Y7TbIph4mwl0qZOHL1B38
sbWmMe22v9Y1mTG+dvkfG3+7xcXil9CAVCuVMejYRxk27Aau0xFNKAPUy+JeWRPe
fv9cCTcaP6qN724g+7jh9tGpywRLJsvfNZP8fMWv9FbgXn2lrahWkdmZ8i00lpWa
vAbTgc1BgmAux+qg1jtqX6RjeMPGnG0PgjR2M+9EfX6b1/Sti7keVC6pc1yXNELp
QAr5hq2yY2GjqjjkBQhJKOBly3yx5tAHS7cWXfV8nOX6SMlAnovBmj7Ko311Gnjf
gVL+EuRlRYmsW5ye01C/m8n8zMq68Dz3LOdKH/SbCwpBaJmQMGKbDtmchU16oe2c
AEZDYrEcZaujsNvXC4bLV9rfRcHGW3Qlu17WBhVgTROSabPhCdWJYih5zq/UH8uT
0d7pIXgtog0TLHp4ouMmel1c6I76J/nqCyV3qNR5dZ0YwGcEVNgL4cO3/SW3cech
ar7pF0zgQPepGycX6gmS1p0iL7KhGppr5sSKqFe4LqQnKnlUR+X0TngnDdz9W/Vx
3RVut1RS8DCNQN5Gwli87HW4BMXwDhObqzucYYOE/8y0zNBp40x4wPx1yEO97d8B
wKE1c5mRWb/CgPJTc9DngMFUxTJfArUidoDkgh1CtYtKEQ7zjCt8Lnbh6YT563TT
JQ9qHkKK0zfVtbAol2YqjrofqZhpFncOW3fSMdQk0VxAC0Oz73heH3+c2ElVp9dq
MIr722qt8Kwl6smeZEMjODhsmKLMCvFQ4Kr8MHWPCsFYLZfvApTY8/RX4Mwtlr8n
6OtsvEGLyLqtkyMw/aVPfA==
`protect END_PROTECTED
