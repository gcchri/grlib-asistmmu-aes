`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6xs0JF9iXQ7/eq787/XUP1c8ybTeWxA92MOLfLK34t5yXCBtxLkaRR3AiS7gQGQw
fYBJNJTkl+YsX099Rt7WlQSytitsEJBnrL/pzi+LNEr7jDf2np29u8P4tJtT2xXp
7MQJEsMPsa5wMXO0AoiAsZKON6sUgd5L5ZLjKnYB2KNS5hsZ4H2A3V/Inhg/DGL/
vD1UFbOQR4f9wswm4VeWWBfYGrP86cIMHJpFTzzayNECG9no7qMYqk2rVDveW067
LOwiwqjslwkJgCG841ki58bgk63tsiqBUrMTbnXFPRoMqNqhSwVzKqrrRjIJb8ta
jpQAjOhPdkRZctcvRoMBicTs13eh/Sk3N1vENOeh4QE6Jk7RmbFh5WLopPvFLHeP
yRX6zDLrDFShLRFHECUfbbIGy44wNlEy2bvPeOH/Ito9DAVrq684brynJ5/mVBcz
Ig8rbpC4FbvwPNiwKS4n4ovrHMQ9tWDCDndgIE6PHsMccu1NdieFiB/8XWhpoNUD
ll85H0Fcb+VjlhrxwwESCUWBHpm21ZLx5cGBZqRy98t8Xm+B2Foxv18GlHp2c3Qc
psHM8UXs9E9aD5X6FBjURnoj+8cTmIrdukFphiuiwM6Vb3rbXppYk8MLXHdbI+yj
pGYbG6W/ZtADsyjPyEUgTbhesAHWwk1Ap7oIo/SlxxE=
`protect END_PROTECTED
