`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
04UnPcz62Ht0jvvpUVMJmCNNwPOETt2vd+ro4poguhDVEp1TPzTfwpcfo/86Gxhb
KKXvlHGSpoe/wAQ5nOgK2tPpuZv9dfQWHFDyA+zexG5E94vlua3hAHzdVltvgZJS
BOCq9ILxLq7+Fb6NTQMy7k/gqyoPqzaShb3H60HE2/NJSPUQFZlDyeZk3/JkkAM6
3ts97+doowjExExfsvqkDvUggW2h7QWQn/k8uoSka6CaWZKPmsLMJy4bMoqzezav
0kZThaOu2Oa5BcjkW6sWK1mXMDc+IPQznxt56KmVnOmGfBlY85votAzfpNDtm+cK
8HFEHuyk6SayyvygiMNWW93slp7y7L28YQrnjmVoTlnSrSE5Zt43QDlsTUD4CFpe
OU/E2Ny3vJsRH2aWk4w9fWoGfsEk/5JkbsPeESL3ZguSmn2MpGgiCxMyAVZZwYpB
YsIXoC8SBb8WhfRptPHAMMC9DQbeXvOxDnK0eV6yyHoxCaXj98h5eAZeytbheZBs
8OhA6zUg0ZZZEy7l/hy1maeMCLFGOge1ZRL3WFV3RRDtljjhOan9K5CEgOVgGTqm
9LsrqsgVOll06SCzIWoRPVPTVkoi8fpnGqRedqgaLdtvV7pSgnSHqj1+6eB3LUAf
KWsfhZoUfjrXXkbjiVDO3hLkKM+roSJ7lHGvJLqwOmK/bwFBOaU8DagsFXw6q8gT
ATsNSfgmA+BeljfbFx0Zc1cpk0CUxyCp+luVFipim50mTM5SL3UMk3fRmBCcO9Ag
5i2EfQoq7OSA67GcS72u/mkhssML65HXKELwZN5tJCwJLTwFPZMxGMmnsR+Bkw6x
l9lbCTHRy6mhO6O2C9JGYZtbKRqUQDhY/YJUHn2+6RdVHHvaEPqtEfEwWSLPRGmj
6QIiFVbAEDB/MQ8V6TaW1Hn+624mpZSaIvCo04Y6tc8ZhIS/gwrwQM950iWWsM8p
Rhpch2ewaGVeJ7ClJQOX6h9uNo8FeeQ2YjliMs0quxX6V60+2RTZvGi5wSfBc1VU
2oESCKpQXUyH5zaR1EUUnH4aj0if3ndhJUO3NifS1JXHFksVqwL0mTwViqgQgMxM
F8YWaGKgYl/ljFKV2z855kolpp2mXcDOyWpYug8iSDWl7RHe6yFQfI+Ud3L4XcCY
`protect END_PROTECTED
