`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q236JMpT7Ye+grcMy+On22b9aE4y26RhQKm6TDhv9i+wmx38rwEk8QH3dxps9d7v
CdwZzKhzYFxEroHcAnFrJ/1JhpQP7ll8+MEWBwh+A3PTVb8W03BoEUTXxXFYJQGN
fAS17hsT5mhFYUq6g6Fhz1CgWyw9sMa2m4X/13hmExqttkwGheh6OR2k4dVlY6L5
Z3dmTHEtGUTd2tO82BSq19nkbed1kPb4RKuWhrr8sbT9Qh3yleUVwkabYvp+jiDm
W/fqjV3y4I1uOZTYPEOAyYurEZPg5EYKfEzZhpQYUKJrSJ9E9pXIb3hQRv/BiIMV
0IQPZQadpPuEwETHIVhw2tjCC38xY+/Qy5UNAHZztsc7dHf0hYUVAJlVA0WO7YLK
8LkzmFmrVTExMCrifm9j4yIc+lAFJe30ojwkiGPt5POYKnYuAqvRJhD51RJRWqTM
1XLJ1AV26p7TtCB7YYpQIXGq69Lt5a5FtMGzrbWFjQNY5+wrBzb+vgcSTSMSXfnC
+eyyZFDbez0YZi6wmXSgjbPIjNgZRLh+K0Gg/U+S4LHQWDlRWORVmWlXE9+hoYfl
3liIMqwOJ+R8Spo6sONL9zrzKbvckrr31putleyUX3xSNkmYNYaCIhA3EFIzxXV9
MxLXIVM0qszVtrStUEe167ydsX9ks7MITtjkjFIz+17V0/3ouZIqqVJBn+jyVv8l
5tFeaUZLP1scLd93zrZ5Joq43Owa3E9qXSlMTtek58CclgQJ7rry6IOi3ERHHxaC
GYGCtWNYL9LVDHUtp5vsv+cLnWk+8SqonbNnZfkJwPxZg2gf0qq8N4VNJEfrdXs7
R75Jp8F7f01yhufWHICshD4qUWIjOgNWyqVQ65iBi/oJqzneT9mBqCsNGlZ8yGJC
cJdgYNNxo5xVK4J+tPSe8JrcnZT+xRVndKmjdrgFgDWDRO8gc2EafDJ7D63iZ729
+JRNoz/hyIqCK8c9CpKgcFUw4CS5NGMC4qX2476BMEoX+BshYnlwrGpOSB2gkugo
F/AGm751aXfN621ceTxXmqS85FbB8/mzG/bP8PuzmFAumdTxtYsZeDke98CO/Wn/
5zZ0PG6OUxp+bhaXQbAaf5R9hlW9Tcz4adt/63NjG0drD95QoTEc8NK1LIN0jOHn
pkdYrFGaRr/LwRFRKEBAk4BwdlYqcY0DdoTWvCKAMB7uEMgN9e0AxrfWj2F0nlzN
/E/1VIOIBNWFGtH0981vRoyYsRljWw6lx5S4J0NKMD8AeCiVBFuwMF/VnkKmai5P
`protect END_PROTECTED
