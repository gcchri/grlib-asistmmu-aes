`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cE1nHbqBp5RTb6BdihR66GozLDP2I5H8uzZ72n7PwO3YtxcPebw2P6lJ9B3pP/AF
kIX8yGCQp8+MarZEOTQ7OFLPxvid9z9hCNaq7qtHa6wMVoZN4TpBNNve8xLB6gUR
MKzh/u9HVCyp7iM7NRP5xeAMksTBAsRlv4NWSS9Q9KhJS5B6wsSvEtV0XAcVI7mi
EllYIj8FMxdydbKrNiRqq1qM1ZvLpCzDxO7AknmY6seDIVNak8wAl0SZwBUZ45H+
bwtdaI4p5c4ltfe8o3ZbFt41UdNW3VCwXXSZl4gtcYdENzbdEW75Mfrz27VhEDUc
pkT2/eOiRJDgdmlgdmoz4A==
`protect END_PROTECTED
