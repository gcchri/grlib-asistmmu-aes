`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sp3JfSSL44IZnjngp0ZNhTzMbkOZmCihRb5z/tUcJzgmoRReo1XKdeSx1X9FrQXS
oU8NMoAWGnPt3ocHyMcONWMWWzNQJQMqGJwmCDcE+iCBj7So6CdS2iHAClc8Li3w
DMfFxcc8L4AJoBGvTDTNRgQCMuzJunnSAno1r2I/QXTOA3dOzNNJr511N/r8q71j
fPs+cqXOHbZznDjiSrdVsSn/a7mXXTXG9o5zO86yFW1VXuwYvSJo1Zs7/6Z/hVdl
tKbBAEpXDt4gni5Cf7ObSIVOcqKzlE9mBIctgu4XU2VxPC44U0xm3lCek3l5gpQJ
aKb1Pu33IKUA8UW6ngzrV0fIruXNPKQT4ZUvMFaA8uF2A2bR6HfRBXPSeGOHCSdd
YPzz367l4rbIRb8P8sShTu+ZChW1PE5l0w8xxBl0zmeEbQ4uLE4OSuev9HDz216m
v5f1tGo5nkrOeDZCOSXwf5/QWYd+lmExT4N7ILi/qqYaJBg4bw2gb+P7+MAkr5+O
vj3SySXDdoQ05jTXCUfEfrv5IGnID4lVTqLbF1an4BfLmKLbImkhgKrBzbXmLyAn
RYXYHaKYEkNAhBmsUAwKpSxU/iBOwtrlkpNEjQfv9Hz7GFQ0N2anzJ+fMWoD5Eue
gcL70stFNAtjB34/5KU9ajUwxHjUzMXJhC+95zLj1jkyG+ayb8wr9Dp6hafiLOUn
xnK5EZE/63bk2Pv0zYfOoa+7f/7KwJ4Yg/IaL41qt5As4xnQS42PqwsINe3memkD
9iLCCPEkXXAYqiaj3ZN2YVxKSbgS2EKoQ8oXi2OualYtoVdaKGqYNwAOnJn2frX1
TBHydSJ9vBl0CLUoTckAvE3lRB6CCUmaL1tWhDqy3iKZ/wnX3Si28p09x6t/dbcb
Ws18HGm3tEuwPNMrSbdgIqDxKhN3sRO/uA8JnjLwSyv4kBCIAPmaJPhnSp+ApR3V
jKZQLtFirbq0s5DPTVWsnWUnnINbB/spsjjOqYNmvO4cq7raUiACn1PRkr+Znjyg
bd2eCwgo3AV0hoaBjhfsrWcu623EVwMJeLq2pOtdNW1B5yAto1EKoKzsw5+raNZl
rq1y7ynoe7h3UpqKPlMbQLVMOZZ/EhceDrE/1wegwa/VXRRYhloJJ4Cz0wQFeOOb
LFtA0uzWAyZjqQkZoxa0Gr2ilZTGD7iQQ9lwe/9B2BcXZgCwjEC7hFZDKL0FIhLj
51JicoVrjyR7P2gksM4MPF4RFQqEsVUKYPImMiwgEWc66sHO1M1pvewCHqqh5Pqv
KZE045BsGSXpJncDvl+bptbnWHFRjldHeqvYy/uEvWppx5JYV+p9OD5lBBQoLaB8
r3uVdTWhujlE9Fa+x0TsOi+mFlx73MzBLeo3E6Q1Hi8EUJYsy+nPpDgU9dxeGkuA
VFYSejxT9bX3qkttFBkZJ0ZoRcRVPZ7GT/ef+ARf77c8DMaDSP92XC6vM/qIwb0X
ItokW9fWtUDwVPi3OfkX2tjTU8no4mukeW34fQYQtL7HjzMPElL3lqvhCZsUfFqH
L8UMXKD0cvseDU3/HZDDRYlcfgiRP6s7ngV4jYYVWbbqj6sRNxin/CcDQxyCPfDt
n7EPG2aXvG7LGgPTiTEYNPausfMd38TdF29tVpMrjaNisKee7qtmSOQnfVsaoDTX
RXaJskaUE8yF08WAuZcRdot9fz/RFy5sWUaRJfHN0JWdimzZOXuZwoSOpK/SZ53K
PMyzKg9oc1BSrBOsoh+6TiBcfuoEGzbBGNBYvAGSxLo0/2LuWNG2183CookgJ4a1
VCSLnU0J/ztkNKX0mcm4LzSXEOYLh8onyCJfICBjhpZNfBVBcM+59SWjPs4Q7MN6
74RqoXEKZtB5sWp3P6wASuf8xckzcFyteKr3TfIa+LxyorjUiMYu3qlvXLzdLAdg
Sr8wClto2Kr/R/UIHDASCG70lAGKZ8O2Z1QPfS4CB5Q4n1PRe5YbtrKzgSJ5FqPa
WMFa6TLp6OqU11Dx/aMRpdsSWiRM4pZVx+jKfYphW5wzzAJnXRB2NuLB4RJtfot9
3RG5qbYjg9ay3hBedKxopwAcQAcQmtnrSz2MqcQ4kn2oSQE1s3e5rV06vrstVFPE
JnzdBr2zRld5PBvNLNOLtcj0xAlhK5puRCru4w17eI18XuhKDLkgkDLb2p6hd/N2
ZnqHvjKXXDzSR+II6IMOd7U+CU6KoHfIgvU8ayvhoXVpUsf04v4HaK2hnAYt14Kz
14SYIR0njhey5IU2+zXsmLn5gVdj4FKSi5akPgV9j+CV26glkmA4BYlqGftPq7Av
0jkhqWRsX/cj8HuRopbFCr9QyNqXnS75fEyy+7dtbCoV+q8+p9w9s5q+x7S/0M5a
eOuKTwwW/qBDbHkvenYYROWpr3jDLd2ErysyNEFry6CNooBJyrpCc2qE+GRvQ7u6
woZqrRE6swEWfxm8xizKXbSN09mShWhD/+wCfTCRDazGgDBZPM7xiknGlQlSD0CM
s4wpXOSI5P6pQUlTjjL+gLBri85G7Qs4P/pjYL0+KJXtjJ2k02moZ1Z55x+9oHYK
QlQStIcaDFwZsqzieRa4Ieqg736GLIcQRuITdpiRi8qKIdHY2snUK1pIEkWMrrm7
q4zbJu3D+4f+DcdAWxi2fs9ZcO0bkkSPEQdp5Xwwo5v4+s/eLOLC7gG4GlgHlumc
GbJg5dUETcHkFVSPmELwdCLDj09BqYDwdBlKI5Yru2dog5JDHRyclVcX5vPRCl5j
/djN8C6DLz0+MvP7aMOZhfI6ccxDWdjzDuo3z1dML6pumtnuSjmycHK7MGNMq8Pj
7nW+xcEy9F/r7dClMEQN818EoZEnbuahPUMGwN2n64yUDb29v3OO9O5qF7EnBRv5
tp8dxj5qQ3VjWDgpx2JEbOMAVu6Arrr55DJObQdaBE+r18ytHsTBi/6MJzEr3OdH
OSjhFVg7rUpboAg7tjOqWbDG3Bw92GCkHL8ib7dYvLh+SXzhNTpnsZVjI9vdyHNm
zqGA/VHUK0fgpRgBZjhR+eoPwsQJIila9AKzjw6872B5LCTTTSt2IBBXG2Tjke3x
Y9gQOJZC70bK3Dn9U3DK5G1OsKg+h4mTL7yOrzhFb7m82saE3Ov+viDbt6s+/LYv
Y/5uBf8EmSZzyk/0x6YzQXVtXxPSWjj3uHBpI7fucR62PQWkeHtUn/XhqiQ6Ch5g
42E603g31MAolu1QMSPKXcQtUh7oxa02Vs1Gdp1RtwpJBfsM6uekwP3LxAr7xeX7
`protect END_PROTECTED
