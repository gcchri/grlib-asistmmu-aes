`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fcHj5tp3MGSHe/xwce4mF/8+c59fNF4+/J8FAlIOt3ikWxojzajc9D8zjbqwUzYJ
V/gb+4irpN45EZe5VmsVakjgQo0OqdJ8i+iLzER+etzctuRvIE7ExQ+1jq69KIoA
G9UH7s9S52rg4hN46RKIUwR6mjCxRspZKrDCWM2X5vUmG2zIDXre9EtwMlifP5KQ
TMXUqK9lm1bmGFBq6Eral+hEzVZEOY6UACitiqSNx5SQTnn8eI8XMckGMOw868NU
6IIjRDGZSgpiAB0ILmt6w+zgKJERtBenbjTOcZrxFm5NQ7z4hH8xkVijO59U3JAk
4CGtbsgigCwZplAjPiepXTCTkGgihENvEn9jZpEVqHzIRq721ooaiYl9RHw6PkFq
xEiw3fkbVVJ5pukgyvDTQt67gKZwG0TkGlJnaaDjeOcyKCFDZrMFKQC9jYhuHqZ1
wsmiN77p8sAvO6lXdpHwI7YcTSLcQwcdOAWdIpSXHPLW584shHFoPeIGd1cPb5fB
ek9ZBmskpzp2wFN/nnatMG650g2MOD5Am7mDVSQe10g4bpA+PR3uRSIxqC5AK4vJ
MvomFsFzRWmT2+B7CcjA8Q==
`protect END_PROTECTED
