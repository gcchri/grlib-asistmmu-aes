`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GiSduWQOI2DNTRK0/v+S+ltVvhDl1zoeDXwWs9zKMnMWHOo6Yw2uIPKYoC7L3PFw
DLNI8c6tXbqEqK0SuaywMcoPCwcJCNilgyGO1mDC5WIPEsX5FpRpfDk1MClTPvl1
ltke1gSI+/rN6pQNW1Uy0osDmoMT9IvUyQdFHDqkqLN1MizGmETHxUZfuoV+I8sc
R7/EnKEvSISNI+fPfrb8jsKmHI5ONWxsdBF3zT0s75SngpZhRzi/FBeymuUnA3Q9
DifdgMoDfgmDdjmK5hFbGMv1DjBZWjU3qlV7Xbrpsfzmfx8xCouM3v+1U1fDxAln
vtoC9XNAdvxWUsrtqyYLNk0CHKBwyLmnutyvRkoQJ5vnz06bBnxXDC+VOcSjeWrt
UODKdFKTKBGCFsrZhn6SFb9EnJsdqDbOPaMZl6k8Pnu7xvscXjsJikbmLX0/VWJ6
5DQdA2ukiA8vwwWYqnwe7OC6T/aUGx5TSoqGb5I1kU5mKbXF5Ezx3DFC/rfrLzn4
`protect END_PROTECTED
