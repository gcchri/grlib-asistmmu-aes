`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BDEmbVlOLqsvTEB915P9DW/DLy76BrTkhFClgb5uqLpgw4Z9PQHum5CQL/V01ZC
JgOk97lm+lmGKzPvkWX+MCJvA2Fd0oK+QCOP5LPleu0JXVgzFgaOLKvo2M2w9Ehb
pGtscDxskRsYZ2Gne8gprzhOHYKc9v9UCPQHXXwIyfgfa1xOYX/ussQcidvl8R4z
tohsnDtrXn0aRIEZ5DLXMhuLhC8aPSjvRx3DNV/YeFDBs7GECFheTlWRXbrqsAen
njLTRiZW13hedivw99vCTwUUfBJaR0fFdcG9+2qjbOYpQIa3023ERmwu0vl5mpc5
whpxg4CsjSRL4isnoMtqtA==
`protect END_PROTECTED
