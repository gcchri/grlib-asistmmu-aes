`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hs3vXxlMc0yx0bmDPYmm3iyIvaXodNu9AUHRrTkyan2MRScd3N4XwaxqOqTSzDu7
opQZAultzKvor1ek/f7aZ9QFxzyWp2zb0GiPrNb2TTA64loe5jGPaKH3wGi9HzJF
+krVqUHROb9BMb1NhzwegZSpYM7thbPh0XvVHzyJW0Uw3PfuD/T7bAko0NZe/EOS
OjfNNUBZA7Ehf6ZpDyHNNJChBYdeJu0ukC2fumAe4F3tTvm9C27ITv9vO+6553+g
nfQpY9VKbMF3Xsfu9knayQ2oprZ/X9Ltb6QCG1cTXi/kkKrf2Y/VWhFpyhNZ5iNe
3kxGSBu3wPZdSmyn1ncx1WzMNyJZ2iuPgQNYVB0dDW7/9uEFm22WmBMEZ8BAFOut
QMD1P20P9qJkyuI4ne8qgzLVT3eqSE3Y69LRAKrwPl9GFYLmjShhsJVKC1jvJjbJ
1W6jMQa18MI0e3aThYcLJeEKTNC3+tm9SWze9TSYXqEV8Ot3Afq8LecVOkVDXAYu
sjtUPHoMW2L2nSxcICiomswtmoTmTLFIpIi2HAgd8YnpueypqM+ysCAVsKb0ZWal
taZAy6m0M8GLMa+q3H7qXXtdu67plk6ejltwPdRhHKxcynpt4GzCFKxYeuFEqkTQ
hDjkOpxZIm+pcI7aC62yj8CsqTdErU5KtzLhrBuQTWtoqH3wS7m8gEa+geJ0le1V
OCShTtir7aZs4GXFEl2/PrmOH2kOh3StZyUYwpek5w+nlzp54p1s9H0MC/TaprEt
JTAZQiGUWGtgGLvgvEHQ+RbfCFWXyCX0C8fyDUdvvLKtW9D0x1G6uzjJftHxrAch
ZGIFW4VwO/N29ZCV2Gn3qMFbnK5ukwjo11g50K+T8iI3mgYtdL8HU1bYWrqJuh4a
g+z6cE/CwTLVmiZCpPAeR0DYrYB6Q9Ce/ViIKRO5UKZY5jT86vgoVB6TdFflcYYO
`protect END_PROTECTED
