`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R7A2IHQfdEI32fEfN1h9/JMsPruO6tIIBjPSFuK1JJopx3pXxF7CYOolDc/z6n1i
JbzxHG9Q+mo+nKC+fsTIpnuk6np1uQpHDUvIujv4piPM53sM06BosaGJIITYK76V
tzdYRTLhv6pN2J6y6FtLsi7J+9IgZrvnuTWkNWKrVBdZS3UvyoXzjl8F9fLrRlQb
6wjWPXPgg7GOj3xRiSSGAb0DTNKBbyggImUIRtZsPEB5WmyZy/vivepO0CAmoaK8
XCV1yviAr8GYYkF1Ch4xHHW/pnoiy1M5gC+NfwUsjgkTfOIVPsAf71I28V+dJN7c
+PF6/W4IfnMthO6CNzYT9+Jouq+GOvGqGPWKyVv5dAyBb8FmyBYLui3evWZyF+bK
Zyj14mSRkay2rfBa+XI7pMBjnUxcWbLYCSMwSXUj8eqEWN5xrsueRZfdZ0PdONm8
sUmBJrGTCZ/LWqXKs9fim0tNetREDJIw4XvEbTyUvywKu1N76vN+xbl+m6hi1ktE
lHc7xObE/0dOq3LbIeEQFu7oEgbEgAtmw+F26SuX0igiDhJSETpOuiIY7zJqmwp0
UFaa3snIB0NZDezYg+R3/VQoDh+WbvDoJJQb/QhU8UP7jtqMFi8TaJL5lCDxVtx0
HshWYtoBMFhuEFgNuwAV+O7pZXYbFbC2xA+eplvPepNRmJCAAAyi4LakJZBl50lR
OGLDE8BAMS+EjSrfwxIlKA==
`protect END_PROTECTED
