`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X4C9V4cKqOyBicUBIR5BtEGdy1FMktXPLM29CemJzvvXD6ODhFwal6on8PufjVn2
5AmAos5S/r3GnaXO5zuguR2MCTr8yQMxQ2Mcg0qN86leNxR5/j/jlxUSZSivo4ll
DDWBoKLW7PNH72Ki/OPwds0G1WEh2HLhRcU/yuL4SviZeBf0ryZe0aAhFKmwG73K
1NKO+dD1Wo0BOfJKRHkIsS/XP4Rqr8ptOQ7H6pM33xwkCYXChy9Ab3R1f90Qak+U
a3sGCMUiOSKTWEB5yu8LBn/f0JP12lLfVi6s9skRnsolP4+p4ZBs3hEg3PFEBatE
NSXMbvbtwhclnMa0QPOpdMKTrnn7YUcU0e5D28/UAege14/inYeRUw745G0nGva0
lcAxuuRRT0qtLTsf3HfGYXHcvor+FvDAIumbrgiXm3zkBhfylpAOZG7+8ME8GZLh
B4ocmymp9vl4RvzDVwtpF+1GjZUMwNTh40oXYNu/PvN+YVY0i0C8cxkV0svrzKO/
`protect END_PROTECTED
