`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kk7Q99BHQsCdks0BNkRXCKT5zQYCS6NMSn5bRK+XasM+I8jg9BsLVxqm0wYrSrxy
FeDS54a6g1jPa0FfH+LO6o4zmlDkQhRhQijAHaNHqequxuKR/sHrHB8E6M8r6SbU
PHFli2+FwdCTRrJKVIFVWZ2wJN3vVlL2XWqWPhCBlv1TYJLgUxdaoyu//AHIdRk7
KZDDZpDVcwud0CZ+QClRNoLAp5A72h7G616sMmh98O/qA9JWkwamppm9r2bXZD6e
RSvHdlhJLO54TYsQcltqlNxprkBLe9QcMYQxbqBMdvFhq6YGjhqN4NDpRsX4Jmci
hxfEjW/jR5u8BvFGGdefa6Cr95BpyrFa6nIjPE2PUXz7a1RYMRJL/TLqgi1tCRTV
j940YcrjUzKXFxsiAwCJI8q+LBlEWWLTfRYD96ojgNk5yoOlyH7gSVBvHuM83C79
OLqIHtxGEjLPUaH56kElyEL0bKJy+6d0Y735WguNWauy5HgD+2XtWax3/R5NXqno
6U9W9BmSbs8W4Pfw7ZZLag==
`protect END_PROTECTED
