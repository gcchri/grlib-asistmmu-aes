`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MOAmjNaCkfd0SRcSP4KTLGiKebCtGthSX8iMoiOfwL0nV5OSoQdoVqu3wcnxHSqy
vIwZkubZQpp6Oie4gwVGgXt2P5Umg9ed/pRtKVXnX+p0ZzRZ3ltNHie+sSv6/Qhb
Gn/97JxMejrM5I0ZPBBqpxqk8CcwMZxOa0F/SnikNXIJOTJSy4rclRWD53eSs+Xn
cH52D3wceAVoJUVpM/KOYrNIHIWTe3RBxpDoVhJXt2bCVFjOsS32uDk6GnqjhPqI
0C1ICYbaNlNZ7kM6wgQ7S93pLKgr5OAiC14T1DzNdr69QjS51/EeHcu8e1+AOxw2
7io1XRUBWc7rKLLReiGQmw==
`protect END_PROTECTED
