`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YRZUmjtsNRq3cvuxS2omtK8v5WexC0xIwRAU+fek7XSENXmkrVXTlQ5rf7va660J
S1QOGr5RZNULmiwABZ2gPwpezuZXw11NraViAwLjbGFb1AMo77nFzHqtibrGX5yo
+pWlF2yDtJyE8I+ESkfk7U/tzlChUxh6/4V0Hdl2hCnkj0lnO/xRm5qndyel9pKt
RZgRUv4mdRs7mFBpet7USYEYYnPLKcyP7dNeCkvllRH5eUrTauahlUgLGY4DKcYn
1kIf6P9IwXkkXc79wYvTTFbMVYsKW3t9aHWbOHgWCcqD3xdnE70vxB16teQgGfAM
C9ceplqyjwNIUwXl/uH0m5WQ4NQiEM+RrL9Ik8sprW0=
`protect END_PROTECTED
