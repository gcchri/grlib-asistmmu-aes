`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yntrEufgKrAK7MafzqryHajxHmXtQig0uEWTwDDNFDIYzb/WBRJtdYKW+eJdYrmC
unoSktOtAR+n1DQe7KD2hqGrPFhNGle2VJj0XSjcwR/vpsrQIXoohUL4HzyHZFLY
/CWYB22S3QH4iFZZS8gc38x/HpLqrkNW97KujIKGMXsI8h5zwEEhGjO90oPA9vFk
mzlQjmcNFwh/VpvqRhJ5KYsERE+R2Pn1iL//xwJNn3gSj+mLm5FXZQIpp14XDY61
A9jagXMWqYmqL/z/5VdrRtXIp/ihTf7Us/SXzV74xzsjln8Ugg+Vetvs/zvwcFzH
x3bYFT+GOtJ+jJhK/EQwO2qi3xDfUa6SPS0jzkk5mz7e7uV8TvzqU4nn3fhQ3rlE
uR4p4OsNjRX0NSZ1WEPcoghAVPBRP3dlkotKwIjXK1W1Hliy40Q/xbs8rRRjhad9
Kqg22pp75/8andR1pWd7ygaG2lq8gid8JZpoIOuNCZQhkjJZmnhEDm/kRXc72EwL
5+IYluUjK0irJQkyW2VM3tOeqOekZW7SKWU6e1hqW9oCdqWTCIQ9NJ3eKEuzYbjc
ntqmPRMnQ/M97FVwsUQbp3Mi12ruh2jl9tB3lNe2DTql64fV/5qW+46BjZ3lnPb9
dOA4YPRVnsUbmAqbHMBKOWsyClbRL6by6agGmMz/xXNW/aLCGvU+jzgEZvjTI/J3
f7mHcls1a58BV3rTvsrkvhwF+nivRfpUDp4lWJiuRKMKgUHYL3inMnJ+NNi0n1e3
NkhKtI26SVu7IG6AsJxhkJ6Bdd8CU0nHJRZ14iTsx82Y1R+2W3luC7EI0HsiFggk
feZmUaL0Izsxyimlqu0OHSm/4ER0KyXSPakpXfoZ814+m9gEd8eHBulPXKtjsul7
Tl2NTSiLlQhdT2md2JY4lQ4Mk7EpB3a3vASDP1mTYKL6fueL8hDhWLevHEKqBbTX
p9SmeBxecA4PEZbI65ec1MH1NdYNLg7qfkTE9Lzry8GpANXcNhP6fgPJbmnc+ax4
RLDtw7OPwpdxuRwyaFuyFIYLT4llsYPZVUOEthYWa1O2Gj1ubt2WhMLNUndh9Wca
GCt/JJwILINCuRXNvl0+hdQBvC1BdK5aycvvFzAng/pfvxmNM+a0zhnkJgwGgn3u
sFQY+eVoWBX8TCStqxp34jItd+tjL1gOMNpU6rW3e4ih4iDHRnMTi431KUrT46k7
f04Yzn3eIwmzj1cF9/gJ28b2GIjQKvuuy1MVjFauoqpVeUiwaQT23YQJUicPgquZ
iFHIMclFo+paROcjKzo1y1a1FQCqFWg5KPBd4A5VPiO+MUSSLwGtdUYmyNSGsjRL
U/5eQsmr6eQla+yXFTAa6Q==
`protect END_PROTECTED
