`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y7j2hXpzIScmoaYFTY0lJIZe6aaQny8mbLPOoSsYbAztjg2gcOUljQ3PlYx4Zlww
jyKviJqhEP7QIv2mmxjRJD20YOyEwXHKn28g8PB/no4zKkyOQm7oPm8Zjvi2HnUn
WllPUm2JHoFjNap5pFvbtLgQTOd9+RHLKSxfhEbqnpDBz3bDCiqarun2T6KU5kqn
4ZD/DbCbgtAM+dAyLzcNGkr3mP6N67XbIJBCrtHhDZpiZ4I184fsjp5OtISeAdtT
Ql/hrMlytmjIVtjDP0jDuAiD5lODZ2oleoxrcnwzQ3l3ZB9vENW5Njzcxvsaj0k1
Jvn1C8TZH7IMcQbTlO5+oa1JyYlPo7rkHpM79WcOvNRSCW3Ju/BGppD8drzhkmUn
rXN9SfaOVEt71+noBiAbeD0WbxNP0Qz9BCtPMbLKqCfMk21HeOxKIqUushcXilEd
fsHFd9HsF7pn1XL8zYw18Mzh6l5y/cFe7OlYDbiZ27ZYsvWSPx/4ouL2Sb3jiMWK
6uhsHnfOrRgGNJDXD+G4RVZlDWLe5FDOhuhaN8BxEQ19JMEWXB6Guui796DZygBr
k3pDED5dOuHWew8aPuiHn8Fap6yc5OA0lwLEmIweygySO50QoqHYdGSOiXHMHkoA
bH5VdJ8/DeFgyrbSl4VdAujFxIuLv0XyUFzS3LTfGh0IGyPRSWmy8IjUNwiqheb8
cEtd+UBfmRPGVvPDOqtD6XHOmlMUJt7BZFtjk6b0bzP9/eMCW+ZmFxsUh/kjvTB1
jkTOisaos02bkb9oD6YlAIMX1qiNaiq1Di949LCZSqC7SAKs5qKn2K9b7gq5CNYr
FGHKWStkmfiKMi9eykryO/tWfT6moPGg1zR3WIFqEyIb6tHSlcBH4i4aTf4pcQTP
+Uidy+LpZHYjDx1jAfm7LRCTr0T6zMac9RZ37ElN7t6MjqMro232SR1PUQCKXj9S
SIVLO/xwg5ldb9i9T0irza1/arjMEvHcD4cMfHR/rVFDxBoM9TAN9xlBq6l7LuTX
PsjbXKRTPC/ircE7T7RtHAw2XUBxB0Txsl3oAveWUBdSJyk6cxOBVGsYsbOWCCfa
REFvWfKvRsLV6RjRTclOQzES9XZHyX+P+C+l8uETzyj5uxLpTWJv7TiIGH91rlE8
1nf8Og5BfHvY/yyuCQZCFF8wRP8eyQEnMVLOjbBtqg3KsXc8PPWvd+PNXrc+p2UP
cSviXK5KzRNSjUEWCdIKV99k7kl3PRC69wMita8fVJgHMoDnvWAvvicFI9hgXZmV
73IgcZ24KyXzhR6tqzihrTGkZNa+vPaqYtImDyTbp5zv65SUb49OwRsIcSAQixjU
EjalE5U14fuoKDrs1ei9sFCmIPwvcKLjolSWuI718JnhvUhoRALcxphs1gfg52hk
f/E4gmor+Mr7cX3d2EGO9Gdfin9WQiNBU/EUU1JJslXUXC54C/AuMzOWNP50XkMn
JkrYyw2fZLXb8g3OdzLoK23aXJu3B65p+27igN/ZTz2VelBewoQagxdxAeVK3bnR
cMG1MXzZMvX5JXU868V1DSa+wC29jqnM34I+E5V8Fr/RkBQE+Krh4GEW2bS2JAdK
GookUs3Lu0/GH9F5C3KnecULgfDLXaOIONgqF1LE9cjhpF7lnE6bZl9LBgD89pVU
clbgdZyDe8r0B3NNzXIjlH5iGdhGKQSTQLYpEFqI1XQFBjnsQ5hNtaediErTLUA+
5AumkTse+44ym5TzEDikxdKL3767W5QIsrkPZAJhqJz2YSO1UUj88wPMRShHey2i
UH1ZF7YDxsxuBumog/qpUDu/nMtDhWj+BwgXAIYgWyfqRiF85G/nBk6xNVA54tKd
3vZ8K5accWQXrzvTK5MyfOiRK4KWsncmTDv9wJBgjevAe5IuPIFh9zECaovnhfy1
R4la871Evp/m3wNBwcwSke/kM46Mvohk7SSy9BWdhRE=
`protect END_PROTECTED
