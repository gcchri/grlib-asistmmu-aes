`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVz0oyLA01llLvhjKc+8S+MYBS7ClF38Q/whfDwT0pYjXQ5MwLocFH6OBvDvL4LX
jYARJWlo5x+W0ISy73eWpGOFpGb8kmIqkC72Djk1Do5aiodiY0/wtPftivLiA6jV
FCIhhZa0ymw1eEVN+ezxdxduv0rcN0ghy1AaiIedz4+RnHCPhS3uTO3y9JfjIVhe
8fLaI2zKH2onyGT7QFc6oOeDvGR/p/2JEtZW/NmZSUDie7/teHKWF1Llu7jA9WbL
4GdYqg5i7ty45Zt9oVhyev5bfqtTGkni3Mrc3hOsl2yxqnVkpDQOe/67txQ6ZlDM
2DuhtufQ3wukRWM6RC6r9WcKsvHtoMDAv6lSfbYvyQ1jT/NeyUFqyWicz45UIdDB
I0kywyjhr20BKvTsvQTxjyfuHCzM/pCE1/Z7BXPaFLAqqBuv1kaCU0nGuombtZ5K
fnAuvwBL14OUfJywUUelG+ormMXeWBy4h/v6vlzYm57XehE2PRjsYXoTbc+5fFA/
DbVGeEvm/qLnvPxtZffMso3cL+8Km6JLfSCCp0gXp9Cf3VzbsgqM9HT0EIrtTUdS
cu4Ad/tbsTuWX6zcYtkXtS2pYB8f+w1NHgBs6Su/ddz9JeHpQgPOVNUXXO/GP1r2
0XQYe6pji9Z8HvpKym+jnRhU0yzlQcTTIpxoDubMWxp27yk4+zvslJbZZru8/jr2
LiStGYCijp/IICXlOdxYeg==
`protect END_PROTECTED
