`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDV8q4jsOZMQuEG3JEUqK2YKwlQXJafPHA7W43OWridqy5J3vDXpPDauJCfhzmH/
k5c5ru2VYpy4BT9SylIpPGDMXuoawDxypdpHgiDkHU4MhDLFNhb3AQO2hoD3P9fW
k6HGVr3H0dGpdSPHovPFJ2Vi+j0Y1SNrDlIfCE0jDN3yyE1s1eK9/pW+WEdIth+e
XzZ2lUKTtr/F+0yZflxMqR7rJq8y6Vl3Qkh+mP1heZAR/ghkV/TChTZvSdUbb0t3
EK6V9/gncoVnvDrRRcVeavB+BzRaUzHgZ2RsB7RnzdBYKjfAbu3hR+BBqOcQFk5m
97uRUzONPISZ5A7oyDV1Y5e1bENQaPuPaZVTIzIdJWVdJ6zddCpIDwy19UNEo4xR
Lxpmn0jhZQZxrnN77omoaEwudhneLBJz1c9Sibo8uTq3BDqr3rvfCXCUpB+FZMNV
tQVv9lMj/aTVvPFoErD6/yG/PhMInmhHctfrptGR16wV2DuIzyqSLQ3QSrzNxich
CiJaV0OLUH1VXkFa9JZ6bEoLJdq+VTJkF/kl8/ZgciNgONl6nUbGvoMEkIfIq6BJ
NaHlTAS/6g4DMMPED/VJiOk+e+RGxGcgmywrVkdCc9y128qggxmAZGKsaK+rCqKR
Z+VJyU3WEFBbBuI41lUYI8ACDnizK1bx+K7C2tn8l4EZmEKriNlWqdMLDX8cOwff
ASoiMhS6urfAkWrG7qeuQduFy3pR7wShmWU0dGMGwZnYkz9GoX4E6VkUzXuPJUUo
IJA6IfacyZNyC89qMqc0RvYwXnb2ejDPkx5DeTtpBoqTbRToxBz01bnkwrxHpIGn
3p0omh2ZRVzIafhZtyYsFDzdJ+PnqP9aOwdzJ0fRnvg=
`protect END_PROTECTED
