`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDlWaE/FJWbjJNnSFdQtj0KQ2EEVizVaKvwvwU2bxQ27HvHgF0PT1Ef2vmxmGBeS
vRbYXzavcTaSMGre8+sYCPFPhBZ4tMAfawMivKBRFjjcGz+9c2Pj0EutCEBe5CCr
0xuSyP25hXH135f42DtJSW6TJl1iuOWvaPUVmjar8WfA3xOKsItvkFv8Jy6czN52
aJ39clnZPEsDryXovBQvDjkDZu6WZGjj0J5gl4ANmJyXDa1Bsx38JNp6mmkB3MDI
FiZ5F/kH2ch8/XifCkt9PFKDc8T31Dpb5EVo2oWO6Dkxcs4oZD8hQ26mjvWbgEPy
m7RC5lqFA4NKUw4WwKp1Wg0md1/catyFIDEETUFd+QSXBQT6Lc7VHx/S3SpHJ5Gv
63n0WDDCfzrVNgbUxLvIwfEJVj14N/mdGPbFFvU6QIGDrX7lM23NJtvyJnqMcxOp
XA4IGiC2pdlYuz5r7c4tIFL6bcf2Jrzj/nn1/6ccS+mCyShFlxNlFbmj8p+daxed
wP7eT5L7wG+ts+CJDgbTcBaWGcrhXJPwBtzW4jDADH7pV/6cQ348fPepqVWf3kHr
cFqEcU+8eOvUKm3WwUaPQfGBTP4RoHztTxtiE0ssZU0=
`protect END_PROTECTED
