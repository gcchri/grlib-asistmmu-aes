`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gRxhb62P2JbQm3MolTX4CLSILUa7tQQbQkZJkMVJOGKdl1FjJ4HzgdjVMj4yPwna
R+5kRyKA2gm3d4rIbqbJ8DJweswMuPl7S8Qgn7lzefeCHPPIoIZ6v4FWqabCz7JK
PVxisJqUsX9tRXHXDkk+8fG7jFo/RbqhzC5u4yHWYv51Gtk1aPXDZ3HV3diWeKIw
BcVRAxWvDOn7J4gzwfOdGwJZDpiqb9nZFXrDZFFjZwPtX1x7JCwSfQw6kd+Tzwm2
+Jy9T1Zk1P9w93OTz07gMLNHTweTLFf9hphJT1GZ1IYuYrT+MKH83zIAbNkEytRN
iD1SUPGA3PxGo05W5mfDXhZtzwhwmPxsvnODxEjbH7JLSXB00T0M0icj0Cx+VeK7
2twtb2Tl0KWl8TfL7afFlRZ006RX/lmp1TFud2dUlJW7rn7jtsARdso48aBX8cnv
s+x6hNkY2dxpAQUb/VZWIc2t1Wycji0NvJdZpR2L9DSU0zy4JZdJDQwDovH4Jh1v
CeFPdyVgdTHrnMnSKpuWs0HuLgKpRu4GytMvBMvER1kjZ9+yfWvL03BlOrLOmmyp
f6BZSZ359gfFjUekSm8Aue/DqeMIrmL72kgOPKT3DULWdj8FiKBPIWrcKusWQmhR
Y6ymGgg5DqHVpcXRHQAehFuVEm2g5rO5ZE4jVVXdozcXvHl8f7wd9EyhQJ9/uLoR
Tl9o1wL4NNBe0M3SUjuxQHZVSCpkkpPkEvTm/sStm9CMnGR3Mo7D0uxJ46KMH8Gw
tWuf8FxD71fx6tlL+uEq+IViJyV7C8Xkmm2VuHq3/j+6EMIq3zzlwRxko0NePbjn
huN2EVODLveWVEKlO4JE3p2XRDhCLHXlYnPMISFAfn27+ihs4ar02rHRxn3i8kC2
Cew9lNghJSevcsJfQF2GZzOrz4bKDdbd/GtdTS3LjhYB7HcVdMIeZymo9y+lE77S
SZPjLcDp3Hw0c/NuB0NVzLtoiSlYSyX8Nk0s8J8CRWk38To/6ryUY1Gc4pjG4BS/
KQxugfEwQGFRPaMvqFjymTb895IpyIgsxSanW6VVeEqJUri0Fl860gJ7dJ+18eea
6fRbTdHTz2CrCJM7DGzN9twxAlyqwSQlderWPHBZwX+nd/Q1KOnoM1d9NxftjJVW
sBY7SUmtaEZ6Pa75ADT0ft4M/l4NcbuOhE6x5jXVW7WGYaI2mxWx4JoMWxIH6PuT
ip6wPcDcMbldViGFpu+1uFjUOgiPQ1ft8LvEbxmjSSP87lRwd3TJ/2w2TCHbfb0A
8rei5HPDgmIIkoeQoMTtz63q72fzrs3eF4uFAlhKsE+9gM/kbssVfKR3KbvbvwMf
Y1NUAkFQkV05/N5qLNYjAuugC/iR9EuJM/BjONa5ok8ixovUzKBlMiXE5UNHrfDT
Qh8SpZoCJlTFA3OberoERcvFpJFm3/BvoLCcNxWFJdip4gqyDRMUx8c+xp3Vx6no
ihrlo1TQt4A5lFTruaC89rBXZowFIB9zwAptsQ9iCXdswl7i6PHsQm38tJfXiIuA
NVDDSGo8wpO717sFioZf6RF3eb76bQhnHl2ceC7hBlyWifsR6in1S2pucqHoILw1
sDVnHxdcgoCo9kdL4eMSx9PxOyEy0+QOzdRzStnrsZDSYiotj1Vc4nPCn06U72G9
tQo1LdJZf7sKGgv2U/Xh7ac42eCpMx3/9CoTg78/jnMFjsaasSvulNaaJ71b9sPe
4dFinJ6EMhr4Hoc1UMRcriUmh28cZMYc5nBjwZu/M6Y89FH+VGaFWym+PL9/cd+J
uqQidn3Ov2nSb5VWjvHd/zQoX4UtIbP3LrkelktrjDAA6U1eKfVpuqgO9b7orCxf
NPXZ5Wh3EE1HJHdrB4S1ta2dMQY7fLgMmC88JAy4e+oxtulnO91h3aezbZTZab0s
gxWn1nGvwjh2kvpcDSjtLQhsmLRhNyYZKE0FHvKf3FPIvC+qrU79xgDWS6qTIbQ2
Tte2eSnlQgPE/Ab2e6yDtLsbSBF/eWq0R0gwf8h2DqzzW7cLJU0nEhlCIv9KYz6P
6h61GRFbjvek7AepuAhRmJzAvSznScY+I8qXW1RyLRccI6wk8QJPsB2WQZ8QGGoX
/zdQyzBr0fFAOQYBVgUgLNBCdWhLiVrEoG3XBbbUlW73euQ/+Zvuw3nGGD3CwsSc
eTWzid9hnQa3XowdeSf2Jlv8bv6MDdC0sRGuvkDeOD/RB4b+PGALcUYLrg2z0nLG
AxU4hC+iJiNgM2VGg876x2AiBFJ4zy+cslbnVTXn8DktqzLYcBoVrRJ/Wc1+KeoQ
5WquNNIUbNXzmcFOEylhqhCt7TqWW+tUrBEjSd3u7k+7ip3YF1Gw1G21UUfr8DKB
5TGXloYtFOt/GDDPrfaHYuXSZJ3ZQhwMPY2bncOFUCgb6UwetFBua7+BC+hx2N1f
AQDrDJtmgSDZoIuNWoZ7ijBDSmAYCkE6nW8KPAVX94A7MJQ1Ayq0xYDHlRDsdG6O
6rW2/6G+mpHod4aPH+S1GlHn7V+3pSoQ35k1FFgK9YEJ53OIlrJudPechKMsX51F
yV25w4jU/xNqC1ByTYZ2niZbFnfbBlw5AtdnxzFRB1oZk1Y7WpDDs25OxEFgf/Y+
IcCsribC7Vi213veFlLuLhkhemMz0EYt/8hk464pwHyJp8B2LRdIq2e6+quKrW3P
b1Nk6U7L8jiYjQJvlBEKLWdzXFOkT/pFqQXbA+6lal3/cBHP/dWDONpb5+oE7KFP
Sm2UZ5wFYL/r0HtOhpVt7z2NW4wFstg9ab7fqN0OwgvRN/Ld+oF5Gb0mgHVTR8BM
l4Q2pbHHR0xKvnHe1QxgVrY6flGwPYHWwGbOS9HNCIVhKAcQhZeOvD1t8U8swHaB
7Daguanxy/rqCbb0MBsK7VWO8GyxH7f7Yg2DjzYLxWvP8hHszPhHp7YXnSREWvUY
9DwnM42raIwK0GaotsjyrGEWmFyaPkXMEbb7zXuD/GIBDJGzJwbfbogK/eMhgFyh
m4rqAbgqG97QXNR9KwDW5HVbyij9/UTY7TpzE/iTGsvqdeM48/PmDWeL8Xt2OFXH
HS+YJq/BTiktmxXCxjWOSuBPQQU5h/XATx/OSWL+/aG43CISJERAPxF4bBM4qiEK
TvLMeGV7e/06vEV10CZlXn/EgwiXPEsMnXfi7qt9etNN6Gh0WtL2HDqXsF+mWeH+
4YVpGN2Dk4Xh1Wi5dyusGrOz7e5LbeZCI6UYdPkkSNGYj12jI0DtKAxB3EzHSPac
sJA0+DWNHdDz8IFIgzpfS8xGRj8kPfq2CcEEnYhEplhky2dKxNqkINr2M2bqjOk4
6kS5+FROj6+GImLUcb4VpQEfhvNOw3OBt6SFTYTID7cdrR8u/1cCKWE8P1pOQG79
pOhjdkIw2eNMU7X/3OYPC2vvNN6s+zbKsMpNqhl2GV8CaB2oDkyTsZBK9TQJfCUL
sa3pKiiD/ePrpiYzdzsqyZGkncgis7RWNTtZFpN4aInHSmbt/CaHWVRVRp4SU49t
6eX5z7j04YSa+Wf+0BKiyb14E7gVgGsg17mhsI2fbeZvp5+aJebugGhjb8NvFKFG
FLGnlhF3Va+JYEdH//Zb7kWD/KnVjPn8ST2T+IAlsfW7fzF9YdgTuJxS6zeGGyNV
u83RivBPRxnAhEnCgsGppbjkUZOvESdJW1wNIL32DBrRGhKj7JPVI8LX98rp6XKa
Q1C35UAFWwbDn+83LRouEO0pA9s9O3yXCd3wquiRY1Lr/jolIcBbAHG795qpyTZ0
FYm21lRF9jB6kJuPz8FxpVn5iivAC+ArF69G8xHZFhVx+9G2Tv3ujlmwQZ5G9G8B
AuiJgRRvOqJcl1j+136c9xy1T1OoNoQ8USy6z8w1zE7MBpOfowfFF0UYIllRMtYM
R3dvRLHEESx4QqPHLL90ZUVCAx9vvENvQvpPdfLncCnnx+facGSqkgLK/QZ+4KtO
VmJURfb7bPaz6myekd2XlXAtKpTJ+dwLnA3G085gxXiCFg6G5c6XW6pMvoBUFuT0
CWkBAkKCyU4oVDvIK5hZDmiGf20ER2vJaLyQ/9M5bnKLlFuelhP1yAT6WGfOyCLm
kzn3YXTdBYa0yI/sibPxt0AlPsK3RJe5dw9iRx1U7+IgrKjtIArMpPo3zUMF+1TN
6UI1t3/WWayFPuCyRJKvfLvkVizWkcJgwk897BaX0b2qINl4+Ai9BrQ/unJCdypj
WbFHfpG2yqPRMDM/jgLmXpSPQlL+reDoy48GTk63MVNO2Vhz0uYxQ48UlwBkPexj
gKWIiEqgIDhi+r1IdoIvrkjGMW/9Kp5nL1qa+s0zwwYrZl/M2pIPKyl3HvSjZHDU
GWhFHe9gfeOHQ/j22gUQEQQG4syQHuQPS0+k1aYiIH14Z5qc+USRtt+xOSuWRaJx
DPtgCTIIxpQrD7j7w6JiOtkLNWgRCGzWSvsqpHevOsNnCl6ifD+oZzjCVGqE71vJ
AIJoZS/9HI7pH5DzK8OXSFRdGdKkE8Mx9WL0CJvX6qQ8rh7E06SrsBS/sOB5kTcV
l6DPNxhQygkcJsy0Ssi/JgkVQoCgq0sPjmlAE70+tE3iN0U5Kk9yI+DdZoDCyX81
BPAbrnUv01n06XbbZrXUN5IkWcn0UaXj6odJ17EPF4xBxmlSlRK4rpVWB3k6ahIr
ydUa6yCcOEiVBXHFuraflJcMGYIrP4RF7Ta6uGWkZMrTSdCBxj5miTOqtUwKLJ8y
iGA7e0222WDcq7VspGIukywLF+hPVIBeA3cQwkivQNsW76O93UnzzAf58XQPp8T8
QcVTABGh5tWA6GP/3UW18758PyoL65/7jMpoGtsmsKNlWBEwoVVng2aj3nwy0lgk
ZcGbpiSHAS9TiGTOIjAArgKqK7uKrIzO16miTAvEP0L5lpI2XowK5d62Xlhub3yF
aIUIBszu621tY0avjwsg8LBr55//Prkg10ukAu/l6MGpO+tdwRQghYQbh7M7zPde
NsJLIkum8LAr2LtLLRWOjNcFG75TTnBqNIMb9aJqsl8Zf4El1bWgVfcS9PLctdte
PcF9wbJ++ILmlaswjZdrge47+NX1tBqFgssAiHsT8WAgXIoPj54V8RFaRWm+e+v+
ZaeWfMvKPC9OJDatSs2dN94O9l0URQKb+YZA/sMZ5BegNBK8YPWBvjx+z+1KTOE2
kQTufq3/WNeQJi7hwaqSZPCPKx1kCbdwE6rqjoruHdixLOlw+b8cd0QYYq7Duei+
+yT5E3BUzPnH2Tv5ztzcE63OGQnVMSN9HtsBGmKPTEJHKn6gTCTfm01AQKD5zd4y
hsvOs8MSf3/KcFde4dTFyPO42LW2SMxwvNWXV7eBipa962VxRqeYws3qHo9LQF9M
u9ImHrc2GQA9DmPL7bE/AfYL3PKv4cUnrH2HOZBZlDIACCNjiYLd5pxZPj7z0Orq
kupiUj6y3NfRLX2P7Uh7NS3WXC1YrltbMosFJabJuUUKYy8RR7NpQCXhOEU5YY50
u/EkMjHhYudInYFvhYfnJ70tNvvee3aam/XeDlGHjjm7CtfzNiG8w3ScU/qh/6kB
5edF6X2PDRi+++q56H0hRkrWs/dqWYeDQl85MyEpT+ZcyNAkH96UDGvrfB9X5RaI
YcOaGrfPqnJTsP7f9f24lrcITbB9ia1uTcpfWsoDToAC7QdsGu7eulhPjkzl4QkF
GV1poXA79Bu0o9ASLvhCO71/Y5HpAP0OV8ncB3OXyleldgiRsdNa2Umuu9lsgyCW
JYaV/lUekh7d168ZkLnNI6F0H2I4wupRY/aMVhOSi7S024dXs7xwHNDsWBGMNqoM
wcXEQtF1yyGtNgAKwiL3JE/3XMQNSt8lImPfvBAgmgXObPef/nQhWihQKn1/gRnp
rFZMujHfxR52nj2EF0hTcL2xTaAVpezZp7RI4157AG9gatKlvcj7p/gjCqTI6Z3q
qTHi3h6pyNZMTW6QgiU2TYDdB47TC5eMYab+n3Z6KQiA/z07ovoCShm2WKhHNPp7
MniF0wzxUo3s65VTtZVTFATd55/zr7nSVBvYF4wn4qc9DkQNzD02sfRZrGbS8K7E
DPP6cBLZEbFhnfpxq4dBZ5NoabfYUvBuKQ1+0uPWQAXW1tfKxBVaIcIoI0CPOxnO
4dI2qcmkslmYnN0iceZaNWVXneVv+xzWDNO/wZuhdaOx3TZn3XE21HALrhohhH4f
IiR2udouUfNO5mctrTiVusiXgykZMb37SFGYxEQGiD5bq+VvTBhOQWHCmUB4GpiT
ipBqYx1T3sV0QFCnj5KLNhZ5AoBfvLc4etcJpPGrWw6dKDIyOju0uqncWrsb05k+
/DF3cV8sp3FQFIox8Qz29naB8omYuWEEua2OyH2kwhS+wH4v8ZazdGpGQ6vlbvR+
8G19cIQXeFPfP8Y9LkISUjZDmo8HDj4lYfqhG3eAARfKsEV7Co+Mihu+3lY5ikJl
dgRM5zfyh0fXsZ4ANY09XLpvFG4Xviwamrz248vwYTxhfWbe1NMjFgV1lCubsHCK
qdYsHK+n7W2sHfP9YL3NLvm/BVa+BJjIlSOy7id4ChjgXqCkZNo+aNNGQjyq8rW7
Kn2B3wj+xoZw3n1XsRldxBP7ZmAXLNevkhG/n/x35MFs+Suyy+Wl6WgbzbkPgt++
olgZ8AzElCgyljw/agp10Q==
`protect END_PROTECTED
