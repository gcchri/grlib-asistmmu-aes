`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGXJ31ixmsFkh9bSZBKb4JqmnFoqcOk7YJKCVhHto+bS6QfCtzDs6nezWseDKA6A
V2SBULibtBxca9jiTLeTzJgAaIeoDdxGKSPwRgYGyYd8VNKnruqEW5W8Ht42Bgft
+ZiZHzefHYdwljDV5NukauSrhTPIUQvxHRVZzGhdR41NTao3XFqTPXINjPNSVcUY
6BUJEKd3JsrFh+ulA7mGC2ROpuhmLmKCnKVX5CORaoG1PrAupctKu6OrQAUbqb3T
lbmN38ATnKne30CQpRrD5A==
`protect END_PROTECTED
