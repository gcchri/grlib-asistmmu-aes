`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGdbp0FjBbOJ/KYXlFs53//Cz61FubEgjnLyZcmoLiK9Ps2EOtD84lFpmx22RpCb
ilNLdSDJHrVblD8Devy3UAuMlYGA7NQylG24HNJKJI1RQ7DMiEPc32vbJMgJBWMD
Tlgoj1AWptcW4xmwzwQ9v9gLqh0x2OkAlN1ggtg85ID5w4kagT7xG06J3p4IWpsq
EIW2Yr01B1XE/dul8iMrhjDHw6p/tY4j7WL1IgNbhvq5QSsqq8idf1FegTqQGjm6
/erz0IYIQcjhejeFnZ6Men4Px3uXjf1d07NBtliEwftB3qtNSm+TbDWh7gye1cjz
BNMr4VdoQIMPmT5YYgrB0wTMwRt4MygSABeykmUrs/EO9gRrPsEzr90TcVqaU4FR
beumxUbx0wGjVO/JC7KqsYgu77tYZKtmOSO4XlZk0CE=
`protect END_PROTECTED
