`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4k0NDOfcMf2UrEncG5PtMX/6h9zZohkMIJof/TFRWgiTrvBE06GgCCjnvcIgXaw
IwZqxVA1KvszoKbcGkLB/Nft6ADyq3LXbvYiWkxHbGG0TFmZZU7qsyHY3petiO0/
BSM0T6qtR5yxXGUNc3dTdQk/QG5SBK2dRc1V+AV66w/4fuVTE5V4ZCg5o/Pyhdz9
8Z7N9+C9+S0qnMqzWVpOAIld2xg91KPRLlVyUZGyFnCyQzUha3h1jgEJTmb/6KVO
0ixUzDQ+ntVUeVNUlhfKMQ+4Rd2JeXuaVv7xcU/WNCvdF0Z9cClEewooNMU3CXA6
Qp77uer5EHOBKcrCGS9Rj8MZIf8esy5FdzRvPxGzCILm0IfOz1lUsTlyww6x+dQ9
mm5jbtxLiluIEqTB+xxjRGfSMi8ysJoD25Gs9zg9K1Kh3Vp93VUNfimTrkKfem4c
hjDpAIj0Q24zJ8dGPlTnp/hnizKV+V+Gw5MjsO0pi9jHpSYlzYHfgl7VQQBtPMpP
2HjijeGvYqN2KsglthqXGvOtUVHaWDy8aUxLHqLCtxxgjSuUKCfUFbNdpMUssbq7
TJOHIvuymYrVwJIIXJlCjg==
`protect END_PROTECTED
