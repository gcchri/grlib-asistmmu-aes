`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OrSSxgLBinuW+qM1/dOnoL8L7pxY1NnQ2ZsUnPmagjktywxtTmmIsSYChsOVEygB
nELsrsuIPI8gY2QIQG1Qbepj4ol/Harn22YSYHpqdJHogdG4ftdEd4Qs5YuJQYZe
/bi3ouabc7dkAyPnLhhShQvhjVRru4605cLISWSii8FXzqCMYXeyTX4bguOE5DbG
IhuWyYN5k2xZThkKWqlYbn1+6A3uKnMVQTqBCQphY231QC8TaJT7CKLcRHg21Sfa
hTukfrY2sJ5p3KWlwf8PgnjEjG/igqZbzBdtcRESZTREEt3jEsauTV779/ifvQK1
OBegKPiCA0t5lOfO3DTm6C0tYdP2a30+4bh65lgOYzr55LVobsa47JJjmf0PPkbM
7eR7SyIWtgQ+dpPGmw6M1Qk9+Crv9z4r6LGEoonnYrzRp29WTRQ0zgB+kvMJPTrD
0xA7WR0qi7reiOIF5AGA/wmvBA1PjyP1Qi1ZkMmB/FTt5gGu4SGoYTkGe2hV4PCE
b5nu6sy/Az7LoA8wP1YSrOB1nhD1O1QhFXN4NTge+pU1/li0QgwbBmcEeADRmxgB
hjmM76GV/6UvebCfsds90ZbA/cnpQfKM8fRKqAOMFtJQId6PmhaJQpce3g3PIM0K
lnQ6Q9p/0MBvRqGDD/oTZPEvH5/LJsM8uDt6kdvC/T7hv+ltJpEnaYYYmVSIxazF
Co/Zjd4eg0mgzaLbvmLvVU1UOJBZRK7PytTEaTLDfjsVPznsjZX1VDx+U0ge1sva
o6UGVB9WHeh4Xhi1deyWMXC7XSjKN+p+TwaRVJ7mZErJeeTRe0b/XkmGsTksIpPm
uiu43aesZ0+TNweRQEem9xWpO8lJyDBryEiDJfhhFeP1jmVYnS1kgN5+HDTDGV+f
YgmWrIPu15OxAYwgN2L5ptATc7J9MjEqMzQqRrldECA=
`protect END_PROTECTED
