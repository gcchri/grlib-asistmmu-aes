`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYnT2C2aB1v3gqb3x8mbR41tG8qy69qV/Wj1b+wXwUng4OC3GwTvOoKw7Vds26r8
kx0B3TP1DJ4Kxdqq4CnZdyXzBQ6QUoHQgsYHr0VvBjah1tPJTi6uH1DNwVppZkYI
udSXHvfFAvrLadzm0VI/+XmwUT/4hhS7pFB1EalwTcN4x3EDJDQghB4R3xL1VqfW
mZJK5EjiqIHYJM0y2K5ofRr051vMStHtJ0JJSro2k9i4xTA+igimwmj84LUqPa4B
tP7k31dKJR8PS5eWXW7Gxr5AkD5ttXuc3zOMslzPnCzVYj1SwOm8DLL2XGbijBAJ
UJQ82KzI0ny1Pku1yFd9DS0qH3+t7xqyIGtVPwWswGyDzKTIKYKSl4aemQv0/4eu
ryAThdeQfU3x1d/dUFVA1oJbGG5wt+Pfqx9RYefaA7RFLgQR7rvsgW8O28Z2WoQb
8sqk7EmBX3fZ0VMVo4kyP6WKIaTm1mLewwJBGx8kFfCTscdBIOKhPWYnK2n3JX5t
Z6RVZxkIjamQF7Q5DGMzgbdFcNKRwIk0O8mmb9hKg2uTGW7261gUeGThldccFaNv
fYSE5Hklwypr8EEcXpVoAuigtpnJ0nKWzC+f+fSYtuueQ4sE6bUvwG8QWNxUsZ3g
hY29Rg1UvH0M9bCjP9YKIcfsRQNPaQNw3YbK14Q9Z8WyfTA9oMz167Fw5qtTCnKy
PCSXOlArkldIUlB+rWGwDUUUcqtuZGM6pSYa0wwHuR8=
`protect END_PROTECTED
