`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XaC9lckHy9q70ulfZBA7IzNh/atD006Fj+ZSNjN0fPG4rPCBmJlg7wQDRRwPyHcJ
zC0/Z/09m0hxIjt+tidKga1bbSmAMUV40tRnLS82sZ0SDsKjlO6CBp/2BKxiMUjx
VFGTcar0grgrez4PgNVqDq4MWN6Y0zN9VJj3TNbHCiScyHclll9Jrp5+L/oWhJTw
Q4PeogG0EpJ5U1ixNmvIBYYWp3n4utKx+5BGS/R9fNVmoqHaTHq71TKL7DWOAQDU
3GrLyfp5FqwNYllJAvJj45IcXnhKurTKfgNJm56zBC/to3FSiHN5JL+HnZvUcXIq
1w0+DnwANMz2r+jKCvA0HMbdZb9FGStiZhoBfCz82eq5GE0jv9q7F2E/cNo7e5JP
zVUp39hdAq3KWVUthGmZ7O9X3M26FiLCnBIYL/gsVL945Yt55sqrs0HeIOk+7smP
oXCbch2f57B1vUBn6PVP2f1XN6XyXX6Bfad+wCCpli7lcLxGUQOuA8NOXaBYG5dw
hUe8PcKDZxicaJCGDJmWcl1Vo36TmLNa9gtAVzr+a1NcoHC8PD6pU7dQDWRKFZgU
`protect END_PROTECTED
