`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EugxrdExHPMN6KU6DbMqF0qIh8tPPzybkXtYcO162099vdFOcn4DmNmUTwOERLaI
Gxxzyz/KAjKHRdD1ul+OEe9DDTVtT78/DQ1Xp/NY6k1pHu/LPjGFETYkmYefxwCw
m9oIJKlNWdY0d8GRT91RSbufGkRduFU3XSdD4u3vv4ol5Vohni8g+DH4cnVGwMSB
Buwj+PU+9ULUB97BlKbIQVcBfCwrbylij8FNa5+gpvmEmcjGNmwDPHpindrY5Dzw
YlUoCNmv5vafNQ8DNAXUf+jHO2dXvXQRrGkLhZF1dXd0X608aPjNDu/H4z/N24Ri
Pqlt19ITOWVXPGk3pmQxK2+aJHvvPsd6hmw9EL/9AIlZDfFCwPZB5KM1vLQGCVMj
iiL9Poe1Z6EFj3C3ml8hK4VHYE/Yyr3FUjNchI+tmDI3a1OUIyfw/+3OydMiSJKr
QEXtE/eNg1hTJvDTdFAgctyplh9tw9EZDBNLXPzzNJRXos5hbdES+b2t0Tm0l8Zn
0wiFf01kyViUcfWXIV43VL3OnQD27A2eTJF+DI6Ws7R0zBFNgatyOiBjcVC85G3s
31X6CCgwZu4X4dZB4O+kn0nRoJKfjx9vQorIovHffs1NDEyX9H9ev8FM8sXUomzg
+O6UNpCKrXT0c0ynIuOSxa82uDUVr8FmXzNFjMZc/etAJ3REsbmH8ctaw+wAiTS3
kXVCHeV1Td9Dnwu6zJZEMb3r5R1wBeFnZxxsxGfM3j3ya6zOH/AluOG5sYxRtqok
lNSfmcj1huWh++2YvjdQJtzGWy0O4kpN/5+TZYYYti27N2OyCnIPMRho97JeHINy
+Gdpbw1r2OYLZCQdRfz7HZbhHqh+DkeqF1vfyozYqsfhEVzDTYAFO5fV+oQiBi2y
cC7/fJoL3S68wp40lPnyC9PGehxxBd83/U2hm6EoIGma3xSq0dKpdmU9d/8x27x0
LOWQK6PFWePDOBl96PzQKnfqo3sMGZkfCHcOU6Fq6Gaxl5IT8ubmN3+mjOdtsJlG
wVFLGvCQspaneCzB0iIDUUaweLxSWm0mkD2GIw2E7E4G9RwojBqyChIBbEbdLws9
xrofWXgFK0cljrCn21DihJclhcPnA3mhvRqxtZM5l0XxE8Od2ZyUFc54xwLTE7Kz
4GQEcvvw58T5DLhqZV3w+o4y2qrUsU7qJOdkyndQtdDNboaTRWWS+x+19XbUOBwf
d37QYatFkI0+1QN85o/QW8w45NAxj8BRqW6SLgbqPkuVs3x9sbAOj323e0DkHVYk
Pv5aVXUQKHzKv0n6LVmLXIFoJnC+oij0vIvfAxdjpCOZvigfi3V8HkR1aGdX/K4g
OWdE5Y8VynTniQOMz1qlrLMHPf5MNzJgS1rdoh/+XamHS3+ex32cMcNAUhe0XrIp
ec6Z1L18PuUdrbvgi7v3WdG57J9Jp4PIirWvzpD1Kf1T5vyYw2LmLVcuL5l9fD24
9g61zcGDFJNZ0uixeWWEK+RJHM7EWyVvkVOzoAdzr5mss1R23RgX3QfT3zdoPcVh
8GZa0rjao2QsEs+x+gA1+ydgr6GF5X1cJakMq7yEmXVTE0CUTA/ZRsYlQs6OQkl8
usTooMrzwGBceFoWnDG4OLanrJNE0//tu7Hjbnr1pGhupCtccF1aoy39ZRHWN7/s
SUnRCIh3Miq4WNiKRWg1ZdHLUZ8/icNiX3CKus+ZToNki12U65WUiYwLt63hKoip
mdwij+L97CdMgJ4vTIzheU99DvjKm+C3m0hK24x13n31w6xx9k5M71RHtOotmywo
qKFMMN45O3u8Mq1f0lAxjkUofL7hCQ8n4NCzW4Q3VQcA8U4Wh3hC2BV8Jq4B6gSE
iXuid2CoWUy4edQEL755a8z25Fka/p1ko2hJn5nb485xQ3nwhgXen5xPC84ov3t5
ESkC6z8sq2ZHzCHZxPheGjY3N68NCE68ev/0yP53pwkXfhBH7gfumQBEdUKTWVH5
IRVgOwAOtxMpL3pRSOZuS4ryFrfVxxZ/O5pQUMruicT2UFlLRlGNb6gJ8L7y1pz4
gwAPikmjR3eM/yi7Xk4Wb6njgbmxFgh95II2iyhB1jloDKvUTNOssMDjY6B6rlbJ
b4DbcgmEMlqubI0FoAsXVor0SanUZ7bVdwW+LgwrBs5gCO565TQsHH4cbyiEMfaE
VEimXfzMWRFKOw7Intr0Uc8fUurvGlVDu6szwzCdECkW/HcQKBKMSe+lPq/JoUuT
JjacbjLsNyN/+xWwjIdZD6sYvoTU9YCnDP657XsoGv/x6DBoLr8fyvWkDyePbTi+
IFjD4x+O70PguM6jQDrMqitOvaiJMC9YW7FJxFUcRVQFLYvgLqtBU455sEZcK9Ob
1lN4+P9P9V9nE2qEjohfTgKGCI1NVWQ7LpLBMgv3HlSzrVtlD0ylVACyc2G/5LM5
JbvRyTe0MVuGQPL9v9cRYwj290D4Hy6+xCSmXWUHgRGLAKE1bCWTAVT5rRewr9Gy
TZvZAQjXlz+3Fj/zxVHVtNDTAn8AlD35YV+ddS6kAMn7uFNFkzRY1Y9/obicWjop
XjDFP7OQR+ngNUdfDSRAyko7NDH/hY5kqBj583NcOwLSj2aB0/PynIA49ghEh+Ot
81uEvBNvFtiXBxORLHWSmqjzTqRfxA6J2savzDIZULxCHuY8ywaeLgix9HaVgSsK
uFZL46Om3ukEmJe0mXXYiTMaiR4koseIZndO2YtsNm6laY49uA3oYcrq7JpkEi8Q
gH6zG1E4IJIV3KtT2wLvDuqvfAiXvuTN7tFRP7+sSLClSpYgcNnqWXF7zCBgRal6
y58+Gq0GidcSavpwOky4pdrKnyKl0mvd5SgmGOpLVjW3ZyFCwLEErELkbxNUn90l
T+rCjCZtOaNfULq2AcDKAVe1ruqZtIT0I+euQrPtulTGXIbUS+6AsPd4KOhFa7+w
C6x6twS/WP0+UASwo+SXw8FkzkD4czBz2dk5gvKnoYyzooWExTCuutXaT49qfq5V
Ta0NqSj/t48fN7cM72JX5oC4/wZgDkGXeoA2ENryDNfsyROk/hjlmp1NSMESW4rc
6aUgN/UWRPtqXTCpmsjnKcm7GShol8gxs+NOghUxMw/5Lv7jXYj6Oi5HdkjfZd+z
rZOCJADD9Hl17fBdH3vUYHoJFxuZnWbUYLKN1L2KMgAzywT+xONKglH1Vk+mjq2a
KduN9tAmvY5E5WCI14RZZ7eTd+VxvN3fUdsrDqI6L83qpXoIQN4qNWJGCx+OGyzj
kemqF/GkdG09qu/e3r3mNyof7Ixsn9PxHZVQCegQ9kdH0RUi9I3qx4i0zUMSqeYB
sGLyLSWnDT+p5ZfxEGGHiaZODc3D9FBKaREf7VRLu/2pF9lLLxzx3WFwNv5Oav9I
u1ilWcDtXV6PI0LqCccfr07xOPJTQKrXuH3bHg0ky35LcLRxJ6+NKgIg0XwpUBP6
/+94guLlJws4qwAJHsSPT+uMEuZVMIj6fRpkLayluPzzqsMaWvbqqChu/O+h/F+b
z6WtuPWeOxcV3Wjw0fEslx/uFRGxMYyU/X91OnylgPULwXQebfmR17zBPx0m+gwk
zcEXqNbPAU+xEdoBkNfOKfooOVqp6oHz3NvXPl6meS+RKFuvT55rHRYSQ8NMSb+E
/mT9NUDZ+riBUTt/KS1kdXkBva5f/3bkXNXricyuqAzLqpsAQasmARsmh5My/kqg
nPePdXdM+Eef54tTPF8ahZjKysHBnywfF30dGbtOttbVanfZuszE7JARwQdPt5Qo
e8lvVFIAEkS2OF/rN0JXhUsMXXlduT6gDBXGmUKc+iV6cRM8jM6b6uVwiwargcdx
HPn5KqvH8JSVoD/Z+qPDxeNuN4CHCPjGIa0Ke/Losz+kD4CMJXMapcbsLbe9QsD2
8IFjCEQxEujwiZxU7LEwTxqn1zTSj2i0BGVpd2q8Sot+e6O+0TQjN1JtoHpgq5FA
F0cRGEYJosePugrQLGAnULNwzS70MhjeVMu6O/stibDzhVKGVf+ZzGKA9anjiT6T
D9AT0QHaVpBevf2cg7xLIYlj4I9Q2two51gAKQrKgRTT8NxX7DU5YbZzBbxhMdNF
x+D0byXdwmjPKdwDCiz1Jedgcbni+2Ub140L0hr/3OEjFNqskLx6xGx9uWD4mbwA
Gya3XsWypBPfK8AqnxQYxYGJxUm0+D4goslKEM7Vtcmorvj/l91XwTBhDmrCDpFu
fg+u6PiLhceho7aUsgpL+LGFmjUnEl7T4+Pdl8kqlFel2fRhv2uKiVCTWcge2I1p
Fcn7pjmsFYYHp0bcGE4L+e8cACJsWb1z42ZtitQcZrHIRX2euMaOZ1yJM7rzWRsZ
1rv5A8NkGYO49cDR7KnquPVnWEbKqlZEjod0fLGumIm03oyOBkU1TM2K7bd4fQmH
SsGGJO63VSwQntmubjrCdC9Tb/J48CLZr6VRn4cjx849amBVLOGtH8uuOp17QK9u
oq8WUhJhmt0YfWLjpoN4chDap2pblHuGqQGUCrd0MtG/+K2suaWcDSQqdGG6+cnZ
j0rPRozKglBlFH/l15FiFVHA/3mgDQRf4VJX9sPtWKEyXeJPFU0pWPY+/aMkCGd7
/gaYBfYUM9QyaWydKJDCa3ALVVjSwLkzOk6xRV+vibq27irYUzb3bWBIltMvi+t1
JEe642zVhBLlN+L4YFaFJhy/yPXYPghBa73YWoEbgg/3U2EP8tMoy+IhB5x7COBR
LraYuvIguzkWRN0A720C/lj4bv0lYKdgjNtKFCgwMp+eh7l0ZEmNVDd7MO1t7nvg
2M6kk6MfPDRveBnlbmvtQN4ry2UHE1c5GjNHdlyMDLcbMYSApv7zQpEy2WeRTnfd
1xnnMNrVsUESahPtKLRKQKcj6cPMn5UHrvvowjPe2uiK99yMQW6LQ8ITBWUCWqxk
+q8kwiQOSp+LgJ5ljtBVcDHbxLf03UuX3g5EeDW3xvFZl/mjaJ6zbPwPtV0DqKKj
1vts2qfv7sTNZtXIndT830zh7aNvqVjVux0PXRQt3uO2b0gbv28Su9+uw0LQZF1r
Omjm/27oJAHnlRFfrAaFX4vHRZAa5le/DWwJTTNLwkrGVNhKk9MxBicY55Spk0Dm
aMBFfLDduznXS3Mmbj56PyzNRsHPgJ/3XhTNNw0l2MkEScKOJ8SBf+KnOeQ73kqE
AO5jXqggfOf64uYlg9tkF57D9eH0qRQ/VaxdQEPCxGoanVr5sPKQtiSUNQBJCm/E
wsgTA+lXI+OCKokpbTO2gM7HroiCr/BcYtF956uB078j4bXhhAwpCdyA4q9C0ru2
IEe+HzEVsSEIi61cl9wehUxtC0+hjVTH2UOcKG+9bIjXFbEugCFKXurmuo274aGA
GZENfa/PNfFx1c11nGrV2KZml6mx0MvpzDbFAV9YubA=
`protect END_PROTECTED
