`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GB8kOIKJWciex3JwtuFPi63PHSeh2zNDHyIdpYepV/BwAOB0+C3JHMQBAQB75gCG
fFuHq9I3nQLYDjXVWOEf2LX8ie+uhoYAPvTU+i6a/gEfnVXGGesS4KjgqKh1/AeA
usxRmJRqnbyhxYFRrUslBbyJ/60g+jQeEeR9Mf4d8fFZ2R1KEjO1ZSGAzmLXOWuo
AnVF84o7oWJ0UtQE8xTxoxaRhTWdEQuvK7JwiFp2bU+2dmsk6oKIeukWeVvSFXtX
6Zg9NhKX9Z+LMD7i+ufBvgJqnWWYC40ne//jjOc2412HXWSsO3hM/mrsUdt7Vark
xnFuOlgArBJf8UyvBPT/A1e+NL81Vj/pcDFSFYVArwcQCsE1kd0+TZfXTEpM89Vh
XMHHZZY0b/ULEMP8wRiJ66k04HrjwB+znpCCcaYIkyWz1Hsot0ie9gID04Yo6uvs
`protect END_PROTECTED
