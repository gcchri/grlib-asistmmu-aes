`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ngS3Zet/luQBdG7+yKdGO2717bLHaLG6yt5mzxeIgIIiGDxKhKSqGpZt+d7dkPmw
dazahyBwCKYLtH3bSNRrJ4kG+sXl+Nf+JA2q2UqcT1iMRhsAvUJUnd+23Nbf8YZW
4tnDcUKVj/HKaveDiZ0rBSxc4DSs+VtSQF6Sn1BhzEa6F7qvqSQwVfgQWXdF7T6c
3e+jZe3+Smo1btvpSCDP/NqSMrR0lCLhxBSohD3XloBEkqNRD/AP2460E4/u2k2t
ysxS2SF4GIDSSP0kHICepX1nvQF3BX3tU0Vct2G+KsowWSNq0ofGQB75s6xBKSgJ
k2XnmQ3Ibvy7OtQiJpAATeuwruxp+lbr+5VuU66F4BiyDCTZfL0LUBIlVnR0ZVzk
4ZVHTztiVNnv9RKQEn96pzxDbzvNSviRd78AIVkv2X3qZXIps91LoBd53AiX5sya
VnBuhARhvy74GNJ1rfBTtcznPYe7HarMfCs2BmVflHKC4ne40NOHBsKj6I8Lj9Ea
khQ9+Bpeafu0YT9uobb+Q8XDoM8LwVfuFpehQ8zif/5+k90MRfvXdJQUFyzVk821
p9P+7kxks1jzOR5caQgtaiIylff9DdZPXjBYKm380lckFZq7YSUA4xSvmKdCe8ld
29JUNCSF46/Oi7Qlxiiyng==
`protect END_PROTECTED
