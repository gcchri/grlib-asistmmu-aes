`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iSXGqNME+qH+1jDbeZJhGgEKLqO4+TOj/ya6X4qdVBz/7zpteK3LnirSYdMNsJGb
4wEjEAIOLboRzKcTtGXWczTHK0nLIO74hUIsS+kgJMFtu1CLfRtjFGNAzlOk43X1
yU78S09NTkW5xH+phDjPwEdnQZo/5fhoQ1sqKR8WQPjT/Xia4cspFlSYBOOQGCfi
lD/ROn7jyZ1kiatHVL6Ai4MeFSKkwqfgsPvtNEddPeolgUsULsxwybIsd0KXCwVY
GDZuXA9XnGn4L5dWw51l112VbpIpcckdL1NCaJcPwdk=
`protect END_PROTECTED
