`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ou4zpkllarMVjUsgUhUCz+YdUli56oqUpTsygCSlvHW8vixv9/M0eoaGmBFQTbMo
Xc45aRhvSRjpwg8lbgVjLjyWyPxMVoIHb5o9nwatZo2PAXSVa553eO0UvGIPai6e
0f1gRyLhb1iFJ7SdMFDXA1xMOBbMz8i5SoZcpP1noPjXRB+Mbzj5Cii1jA1weCHH
lkXUMsC6BpoDBPCgQZPuvYRxIrVy83pX7myfbp7lfDR0eKGxKxc3sMTvAtJoXyYY
dPO+9h5scEs3CFCcNWs//DYvA4NsRE0itfElQYB1aRSLPwc/LBkSlvi/Y5UyD+z2
MfVM0mV4GhLEU2JdwFreFtwXpxirrJFQNWVoOVLwu9T+aMTkg7i6lBu6veiYcFQs
Y3BwFQcLuOMS6YKk1MbzO8Z0S4ytEQYaXH6p7r6p6VtD0lmFcih+utOI1oeh+s0L
/2TtbfcitOB90htOMt4YOns4LD91quuVEidecP7OXI+BaSpTETnwXMF1vpOoaJbK
+cXTHcb9W5X14gRfThFTmS9988he2w5yDwqyPpwn82BCwaSg7ustVOefUPlERnwr
6gZNoT8plfuOnih7up5xZnBw05se/8B54wRClADe1+E=
`protect END_PROTECTED
