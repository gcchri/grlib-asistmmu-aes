`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0j71dqwXWESVGgpR21f6ufwWNNADbgJGFb5MhmKjCtMl9IbrGn7NmLxHLP44nZcE
2DTjQAlxSye3TO66ZyrnuSzEgam6hNWX1TPLvjp+UURc364cUlEpKtHAqec/G8wL
QVsTtm5fc6zvW/+qOvFPdV5gYH2ZlyqDAHwQ46mIlqxkOqNxLuahU+sN7PheGs7b
4wDgg8QGo8PPN3UVpKVYQ2j8ea4QLarAWpdHElXJ7N6rJr7HSwSW9DXkuEljkyaY
GnbA0wJNkbYIdzxi4GnbbJ8I9TDukBDBBeEdYdqY1+RCVWBJTcKK4vKoUhu6uicK
ny7yYbkhug35TzqflrjarZ1NDfJi+gxTntTXCprCWNZnsqbaQDqlBI/pECh7dtiY
2TirOeoIS8d3N8jMwunYNidVVbtqJ5P7yuARdTL92CvL62bMyY06ElETjp9wcwZv
HGWveU1IKHOKlFoA9xlLZjU7IHtuIpmksFpZdTgOeCkOzCtaVlvel+3aVNSOChUd
sV03M6WecjwJI3trUpHWPNnHhSVwWg1koZprnLNO9zJanl9V/eDsDiBEtGOBcxRF
2IrtMvbJ7EEDR7XH3vwvALNF/jkBlFp79a6yd9iPCUNU5tRyg66GenqHsv+x0m0U
ew3SFDtAt+KSe9sW23ZXsKK8HccDceGc68/FLqAtOswLAK/I2VA34YF6GNNUg7ro
H4GQfp3vfu9T5DyktdaproGRHBwGwbAqAHJbNnqR7UmD+2xhsejKP3hXfWpGHnvW
i13AY5rI/XDOSSdAE+QX9oumIU3uNnEHNSqm4MYOvz5uxhr3d7/Oj+sT+GZJNrmi
hl5dgSA8uJ6JJyoHKvzQa3uDoXFLbMVQLXk56JXxqn+iD27NIk5mOx2893bB+Iu4
ru86e2oukQxXKo1vUCgvg/wGW7I4dX9wNZjiLUEwRiYmgokpkHZJYYiIUK9l6GwH
qkEmZaqlpevejjjlJQRa2ZJ6/VMgPQOQqYej++UKl0qmqOmUp6FuSEee0yZU+qhP
X26gdZvKVuooksErbpdix4Q2J2Jw0qoIaObPARHqEEADX00ebAi5SqdFDBUnm++g
kf6N64OzVHmS2TR/H+ZdMkCL+nwSnEquAJLU/r0WRrGn/KPgFjY/YRA3ltBaAdnK
iGec2gTm8Zy4v2o6MKl+4IdhO3XDMTzQ3tNB/slBcC8=
`protect END_PROTECTED
