`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nz5D+rEKuqu18sqgAGUmKxJJqn3jrO3v55qfDmQzR/U+6CfQkVDoJciH6x+W1DnR
3dRT3AxSBawez12bDfsZnJCXuIYX9aN4s/nlqhJuX+8LDDA+HhPhzR4zguZlkg8x
2R6s4i1nSEpw6rlnL61Kfg0aHD0YG2xdZl2J56NmtMMqq59TAL518f1kygk8HH0e
iWBx7KYkRzRWFhMcTKo70RVtt5x+RN1VpGfArhXytYo32lCbwFdFpniGU6wEo+w5
FP+gNuSPwYj8roeLAYH7KZwDWDetRDEPv86ppeslCG9Q8C8A36wPiLGD9/6s7Dp3
4kFA9xpOPQf8zx+4Wywt7g==
`protect END_PROTECTED
