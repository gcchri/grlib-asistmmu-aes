`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qG9zZ77pM/OOnZvTF6jP33Ha0mM3t/FQNbpz4GesOfQHtP3DFDRxSZmbpyji0oqp
7N3gnaoX93erTHWA8pNq1Xx1JFus6yB3nu9144E7akj0mnSgH+uZMAXZbuiniHjG
1PvK7Y7qmFV5tafsPz58LzzGGBkH29ZEGdrXWsa/JCZe+4FOeJAk0FUu43mRq1S+
KR9ADtmJHNqe8eAo95IIov9R0yd+5ufHUnKNVVZOA52L/QYcBxUZ8IO0NJYiax38
cFcW0wllW8lt3rIvbe9injfZ6fUROPsChEaIDoSSnh8uQEcWtoFKS5mEvYjqERFE
fHFXNJflfqkq+A1yhdzNatjZeNpl0NN6msjkW6Yld5ALWCLMMeKXGQ+G2Wi4K/dh
hBq3D/iWkN/JyrTBzN2M5sXKSprmN43MG9TFSm8qyStR3ysQJ8iREdIcXd9qo3NJ
6e0k06opI12kEJrCpBP4Miqm4wMVDGvKJrOfofH/7Uv9AxFiDv+YU5m3ODQDmWz8
eHPD8/I4bef2fAvEqxQ00OLPQXeVrv7PVMaeQkMxur8jhlQ6EijTAoW9Cnu1gLUM
ueeJclaKXfPuTuRigKZpANe0gvs7Fc9eESotiB1VwEI8+lk0a2McBXJ5nfbmRJyF
91zfXJXyILl5Kit5BbAMHo7fD8r9tDiXKfMGBwBySAdGv4RgDRsC9zmIClmyD9hq
`protect END_PROTECTED
