`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RYhWero0uHqZ+0lC7LmimN3dkGeEq7K+aJNwZ3AK/8N6nz+QR4TSz8PIhp7ic/UY
7QT2Dt7nnsAtW2nCFjf0BaajTBZBHKClNwfjtuS7sDggvfjU1pFLBsDRKgVBXpyJ
v7uIAy0BZ4Y/akzoFVcGYHp/C5p45YyzTsHVs0MDEysi0nqasM3nsEBzSEL7ILrN
2Tz5nGBBRUMB/9QSbAkBqe0tIG7chIuYHu1MKffkfzZdOXwaMPwBtrKSZ9TfJ8dl
DLig1wYSNOSfafSLrZxzq6BntUKcvPsKQK3rIT+k4Q6/pLer9YsB2Uji6sngM77l
nZNmJylLKj79sMkWh2Mz/zdCurew4OflpTHZTjXTuKBekyZBJc/IoCI3xW/BcH+R
Iuw/PYbZL469YwpmNo8kEbtwys5wkV5Ui/E0Pw4jgrBux/rhfWypLiAQ5EmnR+qi
YV4UoApoAia/P4JFrNQ8JtPHt8r+JFgY8hxdojexv7MG+hdkY0x8mmqv5TRIVrcO
bXfICLxcuso+CYISUCf2Wj1wV7cfnKoLqaacbyWBGO0Buc4Rp/e0jvC0JbN9mbFI
htwOewXN1CJFjQxrtygey4LgYFuiDjysj/VhhOXj5alZaVM4fhLSQVctvolqUsHd
aQpciQ0yWEfilI2YUZE3Kw==
`protect END_PROTECTED
