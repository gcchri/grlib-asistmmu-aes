`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FVa9aNe3I1OuEkfLnkmf2A67zxMPyOOTIEEJphC9hYwS5zIaioROLQjHtOzK4yxf
FlttirNEdVNSeX3Ut0YAt4B9klefa9uy2/1TglcGFv+WOvXjX6Ne0W8RyISo8aIr
U7MmHJCJsMAjXvkI3fTsLRdjH8zJYOyRyVn7mwzichomDcJY7ONpsF+XvM3hdAu5
DYegRHP4SCe0CFC3nnkbM2Dy4AEjAvPjsjjoc4XvHxd+UGS/XnCUjOssNXCshc9K
xjAt7cR1eykBaiCsl/xfluPFGmYTesp0DAzPFDaHXn37TyjlX3O7NYGkgbk4Afww
5tH1mMr72cBf5pVaqFoFZ0smOeeA8w9AqmEeyQfrNAyn5/z1j+m+ecEA8OHN358g
ZncuUMvD0fBmgw8hwYYVjui98dD6VasXalUhN2ldCAI=
`protect END_PROTECTED
