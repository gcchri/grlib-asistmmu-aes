`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vxtrJas1FrzW4Nvev9r1BroAobdvI3Y2njSf+R1FTciSiEi9pWcV8zF2eIVEyu9D
6t43oamyAfM1OKrMwPDTYGkI70NPox2B1Wm/OhPBchBrOSB53eosJE3pGeNbpaUV
HuF760oBozUoQMdG+ogFSCFuEpC3XsQcPIS1nh5lgcDc2R1Lt/wzJG7o8h6SPaV2
zAza6XFj3362jtmTvDU+KgQkkD0Pr/l61KDhyOq9BKxhMmgb8x/6U3Tn/34wIICl
iBFFT3+4fVOW5tBI+KC9sexmHx3NN5ggtvnprmeiwd6+FQjfo6IvITs9V2YgHVMw
v99Fx8PE3l8KQmHuakTt5cVIH7OLcCe3uDj4jC1+qPsBX7sXDcQ1E7FgxRnsrfaF
z/+m1jX+XOHbFLlLhM/XADwGwNhODU5xK2ObwwNSTYUSFca6ppkH5dOYsQwVuN0N
E0gfBDbxkMuiqFz88EYuuSP3hhhnFbw6Yxdq0DaE6V4XzWmu0Ze8PJgufsgpe0OP
FRqhqpAECni1ikgLpLkuzccg3D/FUiz68JL8hpTr32iT6b4+eLXpLF/bCR+cSTd2
M+utNwEVkWnnF/CCn1pO44bUYpvSG5ayLfIRj1Ndt4VUgcInNxlINIXZRaQ0jQEq
QbPuxB5zOfoZv5MS5z5zu+dTUYT6+ZVSr6wSOL6k1KHy6e62gaMGSPBKCO5CrVUu
ws6aDjEg3VcTgjCy4sJnTmprmwHbUmJOcj8v/xsmwQbnOMHkD6Z/66l5dSAPERVE
W6fl3M3xN0W7bNo5zmt8TMdBGTH3LJiaIVPerbfvN7wPrj540Ny0jS+6krzjpOQN
dHZBdmcwFe7w44sJn3Y5z2xfT8mgy9/diTHw3WURa75yMFW0HmjLpsLf7Jv4W+GA
+PQAaWw9p2uzuINZCzdc/fFvOEfjNrh5J0niOI2J6AzcZpd/jplKC8cqZ+LfLJ4c
blMN1g6wvthwcxKU79akbnhqUONAWttviNyGWK8kTYXfdPo7zzktVMAW/5nyUt1N
YNoAAz4o4LcthdU1igko3rTTTmFnL9V62HJXgOQ9TzZvtymekCiEhXrCBwsJZ5MU
B6EsIMMZniydJiWhIp/eTw==
`protect END_PROTECTED
