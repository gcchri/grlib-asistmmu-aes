`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpAnGcwQt/Gx1az3bYRn8AD2Or71xjj+zh8IpoJxd9uYSJLNdLtyr6j2UD/8qIJZ
Xcig7V6K6L2+XP8TRc0em6AVdMLJS+SjQuscenxldUgwuTCs7MCVKJAm67wPLAlY
zyRJlHGaYNT57Klp2VJiNmwhmaV9SGPIs+BuGdGmBkgfBpnCpPNbthAqkQpXx6Q4
XqgM4XWeKG5RWotkvE88FfjoxImmRuckj1YvhHFkN7xwJJd/z9KciDNiiM2/oH8p
QnXKw7P0j60JYsuZmYs6yzhguixGK0zGQ3FL/hv5byv/MORNlHV8j8huODaf+Dcj
bw/HN91h3XE3CgCiL4K3rhu+G84sdDD+eG9/f/VT4T9E6SOcUTNG1E1jmU17M2j3
UEJoK5fkEhlYBTzvig0zPC55PNXvuHNB5xvw7AZtIOQ=
`protect END_PROTECTED
