`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Z0h68SE1bsdCuOujNsMX7BKuqmvVQc7ob4XPsiCvfK/AVMcB0/j+GxGby0uxHu9
QQLqHQz4sXzihBS9XlCkpM61whGqxw4YtOLLOPHrtZ68vmZH0x9XmfjVJY1UAvE4
TWKXuEUpfcxvq4nXWewTxmVWAY1nIj3TJIoyTnbU+IgLiXKQK9ZScBo4gPwmMSib
wG8DMO9mYE5j80lMOCHKZpJHYS4FyYOe1MQDQU05kMM6REh6CTUWHEK7J+2Rgu/X
TK/ejDZWj79a2yXn8ZcluEux0eb1JwXGJNAJ3oobpbticCkCgryLS+n8uSYXYIqe
oMQbwFEJgrkmLcth1skRNBRx5n+9+vCsMhD69C0/UIffEGyUBmYN0+7G8frZOFQS
GmSFM4ancGiRh3d20jMi8EOeBXguqoiDHYylUUdqsluRejp5VEEaG5SXQS47KK67
MR31DRkvRkV4bosTHkHwKQ==
`protect END_PROTECTED
