`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dZDdBPxl9UbXBDKC72XjI59QnQUGGv9832FVbIMtRogZaR/k24qtgUOVK1uT2m3H
MSkTD3I+7K64yLQpbpuVfJqFyvVkUvkCQowbRYXF1ht+/PDkSwFJMGk4CrjPlGQ7
UDiMKRDBF99L58bJzacoj8UdriHJeEBLjYEkSzTuh2eIxO1WavBBTntM6Ty2u5bh
shOsou2d1k7duTjQxQYjHb0KY/8tML9OqljWetThukhfXViqt46/6aD+tku1bBoc
RaBBkSFLQ1m4tQUs6dgBcqxULgdgchKW93uqvsqPtJUGcTL5GatGIsaJxxbaYRc0
Gp/ZHoSia0RhjwwPtU73nE5arUDiXp4oaTwHPjBrrn395W9arQlkSiKa8aGTqaJh
ZFnLCnBmb7RFPCBvr1uFvet+JoivtQBUHGb9nuMg5IPh9McDIt2drm5kSf7cV8s4
fyI9qUB+tty6rkreRT0Zc8F7qm3/VRX4xMsHiMRDyl7PmKGpftCypwQp/9kb5m97
WAR9bY0TZyKrtTKtMuFroprIG5otxjrj2CdNj4HSpDmmmAw1yKpS7mVcHTv6CNoX
q41sBCRWe+MPnB2pBsW0Ag==
`protect END_PROTECTED
