`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fnLsZvdotqOlMelbk9LwxLbMu42u8IWbh3eWx3Fr9Cj8JOF2gMxIF7bD/5SiOxSr
9b1xMKLK7ovUm63FX/bBq5JkKkhg8TrIdFZZ8TCIxWHV3m9wV3A8pPnIVr1NUo0v
+XOHuB1H5eYscpzPTImgtdAWE7sPffRK0pzkbenUf32fyenttGgAuclznK+5NtQI
ApXaBp4NefZHAzbmkgkuo0uiNo1+cBCx+HlPI8iqf4/7RMhsWxwhKF+EQyHCTay5
SkFAkqVziDMdj+r+wzkB0x20tKkqQRdUavMjkg5Cm9XAGm8IwsPRVLeDVOFRIrCG
8vfMhpYWOQSxiiZe89Qx6gyNqYzHg40GXZBKSjJJd8XQUgeUIhT2peJ6gBLN0iGK
PPDotF30wzTikqyTHfe+sOjSStEoVR6830us4uCjl/QmHkm0UxxYJkvoC6d8oJ7X
O0Mon0JlGpfx6gaiQsOEHIGAPAPpCXanTxMV29MG4dyDLGneAufdczBW+q48X4AM
F7cuecdvSb1AjOLqOZqhTzaIKt5lnHxvsjwtG7hPvHEbIgV3nV7F8NpRU5n85NfF
v9YeartPw1NDctDRrNRFe3j9sipAqgv157M8lNA155bZMZ/cHcD5UaiX4TaVgNP8
FhmY7Y6oyGg+bbk1NNTzhyYwbuM/8JirB8lxW76+pXOVJ6VaL22ThJyMpno19NRW
Cs1N8IV2Vd/fe1RpoljDBsYiPoCvZhI1oiDC2PxH9xsQIK21a++T/3/KefmbTZru
qS1zsE9hXCm336mqYsiyoiEMfu7Z8nzavojePXiSo5Ado6FwLbWHdAOLi+8Gfy2f
bswCLdnIW6rlDiLaP/7t/CRoTzCz16yQ8R4fAjKtDS2tuOZVSfO6tu2ToYywQlWw
c+1UBdV0KwKywoZzVqGM4SUG0U1qGCCkbX+Pj0ABimmkL30S1AIpeCTey4B53Zde
OgyJ1OPXl6uE+GWIXGn9N7GrUvW8UWLJpC3TGqSUzKHh77sJXNrnApG5h8GW3cH9
SV8H2JM+cCq04/4JHPjLcQcUVzJYKuUBNIwVF/1zKuLMdUhf0DaTz1UW0nHXry7x
Yqa+cIPaOtDjXoMAOJEF0g7DIE5VX0OMHWnNevsE7AcK8tRwywAuBohvD/+jOOVH
NBbTYH3EpfvwbU9STdAIEcrU8nl+eerH8HgPS6a7BG8DMezgYOwCW0iiBtoEwn+Q
+7GjLj2UZvBIS4ABKX9naFlHH/mUpmpq8/7mWjJHqOoRJwjQLg7rp9bOIJG5kfWi
IIYJixDeVcDZN2Lvpy6PizRoHhae8Y7+EGkmd8A+jJ7ulVqoDolSLlYmy3WVveOu
xR4n3TumgB4kTvIqa+31Q3FklzlqICh7J56Kze3Y4S5iAcNnqNiMqUPnhMaRi4IE
G/77hDpu+9mJpzbuzHrhpJkDQCpCnRPjC/i/UuWHFV/CFOuStdshobTOBbcRHqzy
6FZld8B0BHXeV/4zTz3qsRfH7wdgaNNf3TTkE9WogjPuUdxZJ6ViVbc4nhalD6oB
5orUydNQLj9/PXwtbXgdpCaYE1vpC4qK9oS2j2wbeff8sKA6YxUaoK4wvGTRSxBh
CDvzNillVyYHF/l9A5C1os+ucHPM4xUAkuysEq8bqNa8pwmGY0FZhNjaAgUAtai6
93utTzV0NQp0HzPf2I7hP0ernNGtRaQCeINa9L9GYTTAEaFqyelyZX02s1GobxQt
EXd6RswS9twj3ieVcOUZPvtd4LWYbvTtTAvAfZE16/4JtKvJFzSRCDXBz6SNq180
79CzWn9E0v51v57Itb5yv+DpYRgUCz60Whnq2oIEQWpqygjNjgkTfK7zb8f0JNub
PQTkhoIwXEmi916JWqIsTlTAwGmBUgDe409ISrhk5qDN0U2Kz72aK7EE1ofsgsLy
kzkfhgaHksN3z7CkG1dtDS0QLnwAi9BoakVuiGShwaoxR+gGHcYd76tpDWa9hWvp
NE7nECbCKMei+u4hBGqVU6vgIwbqR0HtPC5NIpbfVFutRkik15vAufPFpSA35Zik
VqZYiqiJDQTtCsgrS88dvGTexH0w6hiFtk3IGr29P9AwKTPncb5wIJRJy7QkTmhx
al/Ko/pBIaRbjytEv81EKAj7Jcphu/meYM0W/4VUoi1eAOOqqtwYYluqjy/k5YQr
BIJAn2Qe8dJbGi+chqMVTz2Kyvq+c6pqMpdsrxri52QadCzcx87sVpkq8SQsN2UU
`protect END_PROTECTED
