`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j3eeo4jKSXrQCGXUnxSQM1aPEjOr3Hv9gsnp6m7flvZnPCDEUDZGjk4RBfyLReba
7hHvUL70td6cjufNQtrUsB5ao737GL2c4b/Uu1EscPnMzZxzyOXQhYws0yjsZxYS
4+sarBpgIu7irZ8wRyAR7eVgZN9GLq22QFpdxqmjJaE7dZn7VOAMG2Ms+L7E3jaE
dV3nxHoya3HOUAs0A9fKX5nr06KPAeEcOahJUxJNZYG9slk+8gQpvaV8OfdIuIiG
7BM/a1FBScp1YsP4qcFmyKSqbMcdZ21WGOtswkAIPOVmJse3V+UaXJBjMsGikMJv
VR+86Q3c8XzWE6D/8qgJ0JDLkzwF16vTdODUxLHCynR+zfcB5vF1DtFFKCwrU2nU
0pwSsBlJ3hXVlolIxjNonOylx/gXnRDNFJYL6fqD1UA=
`protect END_PROTECTED
