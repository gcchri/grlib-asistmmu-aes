`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zomuyOFSGsnoL7zq5wuzhZpTTgG1m+t59LL4C/+IjwL1ofhQ0mjP8I191QzLtPz
EGRVLxcsr4i06IYeNL+npYZgfzkCwuW34LBuI3g4VXGER32s9QoqEJRW8e1XI5wp
jM0eN+w74Lgst1D8iqUIO06Lekt0/I9Qnx+KMi5GwLoAWvjZmkJ8i8uRK8gQxpBN
52o8TYpP0Y1I0HvkVq4dl8j5snd4LTysNRB+nT9v6C0wbI8zI/lZZ6lQwrA2SL2i
kle4OxywHcscb/Orsm6i/BUVNJFcGkM8ya9mvPS45/C/HkKFtDqTMWjh3PERx8hU
HK3+GVAg1GBkqKZjMP1oM9+vD39HLRqPDUPjBPXAtpEDXvmGDsowCQWC5QcF78IY
nUleiGVRyHe7wxoQfdTcq6MuIernEx8cq/fx5JMEOww3gFtIo8mjRygVjFY23RCF
`protect END_PROTECTED
