`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Azj7/ldDZKDBmqE568eJIY9ll/cR/dwfkV2wlCEdj7hBG9yLdcyBy7UIih12gWqC
po2NtEKEntV4sCLf4LIhS3loUc6fIzKZVcE2w+jEC+ky9dsZ7FqH5X+VQXrNdgiX
+zrEuUxN2N/dVRmTdrlaJMSjind8dxdEvgMO21EBQ1A8E2OyY4SIUYGo90WPWHQo
JokvRcHM97jOqGeeAO1vnWZutIMqNxQ9qbxuMYPA2JamP7mTbMyvDmHV+pYEDNW5
HTnKbs3XSBkXpTCUR4BH+vtFFOBDiv4Th6aU+hegvH4PT5GOW+IUJRYZZS8z7t5y
KHWgXTRT9nMOIZC+HY4ZC81Kfjjrou5UAGxPJd+W25PpL7EuttoycHCifM//Umvp
BxOK23HioXvkM08bJtFFEQ==
`protect END_PROTECTED
