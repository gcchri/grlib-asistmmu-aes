`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7oO/boUa9+kqqopPFr+I+Id0pLXSK0CdIflhffOIHUKxZSOugmLqmjLLl6GY3I3c
D7qoMLhFIlT2lBydPDiIvt1wrPBgq+n8mgGcyBZGa/zxSbk4MkzxqudF1pUm8sDn
NOrhjkJk5K1oP1ce9MMFk5nqzBntOUmqgW+a/80P58dsPfGAHfmMtlAKrpObcT1F
yWQHhc7/DFe8MhvT3d6sAKnwCo89h7QxLp4oxInJSkIe4V7HKnM33TgeLb2rNsZn
2N+6nnezb2tfkc8U2WHCT0SztC9Z4z7nee//REknd+p0STCfbvdTvznAvmcK3z2A
eP5sNMavedjlzPfngqts9UOQ8BOgDGjaNE10ZnQnoFs=
`protect END_PROTECTED
