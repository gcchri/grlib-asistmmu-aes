`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
az2wSuVe0Scs/CA1hw+O5FTWKxn6GKkW6l9snQWKYC8sAkx7g3M/QfvoYzB1niXD
gu56htNT18h8XjH2p7cb4suw+/Tgf8IwAJGxWCOZJVFZBHFmxCdHG0JRs4DQc1vN
W72yxYQEKKp4G1mNk3/Z+OsaZWIUWSPYLk7Qs5ORFMVerW906sxdm+3h7cWJ1jkc
7rBvlPGKRSADimmdNW/msvfg7EhJORXrXgDnF3OC5r753Agm/QAm6C7j36Iax+w2
URhuQFDfxdhw1VduGL+QhGRBrDyLnc5qpC0Ju3mzpQWhW1Rrt/+0gBh4ZPGkFtkd
fS+VJdbGM7HbPHHTIEiNYxbCG4JFegoxZy+qcBWzXxIzUdCLQgKqq8pv+LRun2sb
71FkFBHoPbt9jxarIeJ8wNhcrBHhgcRdIJMaEf81l+6idsy3BSN1WWckaavZSFNG
rdv8bYZfjJsCKwTqkB4e6iI+omW1X7okHmReZABNXVMfEhAwSDwM3ExS2N6yRAZq
FwmbqlwjWmEvk5vGJnOisSUGT3I69DN3h04pbitUQJQ=
`protect END_PROTECTED
