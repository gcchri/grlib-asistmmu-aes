`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vW63T73vb6QfIlHqzwRYTp3V0QyvoYMYYkVRqb4s9anRMzYX8qTMErTantAL5s7c
YpHMlfHmxESKOW2n75PlK1sY3v4fTGl6SZIYjTGk3GC8s7qGEEzi8MX9/T6WOxZm
IopcBLziFvh4UfuGYl5YyinHFK497X+xpeNc3xAVJEW4irn357crKWcJFaDOrvnk
MglE1yNF4kUNjy3XLS7cK6Ex0CGI6haOwzy5V7wqIOwfvPeDREd6adfdsyTGNBW5
fOnq0rGYaB1r8Zroa/k2nJEZrAQYdoz7BUFPzGcpUqYedFFaf7HiytmT70Lji5qK
AaoqGWYalOtvcXfjYaK1Eza+f47gKp6WIkvm1Flh5+n6++jh5X8SyV1oxyQWIY7l
4uC1eLEJ6nDsd6p6pio13FUwTVC076uVaPxc4dQbJtpqa+Aaux5z0mfpKggGqAhn
eY8/p8kgRxNnZehOzrNO+a5pXToAYHFIKKYeR6f1dLo=
`protect END_PROTECTED
