`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzNK+t8wVyrEC6gX1GDqCGME+B53j/+XVo1BfFbJXa4/JLIQ4Ps8b7i3cUnznhG2
egd2EZANSBteMgPNTO2E7YJTxpW9G8t8JpWJ6a/9rZzYB8a3Ni+kAfSa3889pSgm
WtW06QxnLX5nYAzROtjM32ZHwpQayHMrSwsGrKqSIa0+V/CUJdUyt63CKb9BX+5l
AGN7b0I758yRnL4i79dWUJGwsGAwDBjYTwFdbm5Nyw8HgGy3L60go/4oJWnTiTUu
CtbS9kBCNvhvL6wMTAg2XsvCKthn7BGIyxvK6yRaVr7QqdPtBqRns/YCUgkw58rq
wUT9oVbFe5+7j4dSSk8gIp4/9hs/w46M2vx4BduNMwRFnZgvgAonq6WxBVY4xWc7
vE0q2p67KTzqwBbPs6L2LkfwbwdXsjoWmS0cdZ0VIfdYmYHHF3z3mHnuTMdNYarW
H6CzA2wvjW+C+XCcsfrtqqPUYUV0RZrnMeC+wfBRsy7e/EGSk/5+7xMrf/zfbF0Y
iPYyizT8/soWQBf3+4yPeIVcuiFX6bxh8dd340ff2H8HxZTcP41jrfbeZp/TFgr9
1J8avqE1IoWAnENqvRbuBnfItMPeU+6Tpo4PcxBGp7dCEwVNPS05JNPfNiK8IndR
C+9c3pSRlN6W5mOyufwIjw==
`protect END_PROTECTED
