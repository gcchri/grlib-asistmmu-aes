`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E6+Zrl6ygEJLDTMJwRaVfAHMCVYQQCR+pYwLJnywAbPouAyUUE2c6G2sm6njR8Cy
kUtT7FYdbMSGoPHVFFbib9pLFRWBKSxTS3SaR04DP9hHm6Q8BIeiFHb9Y7Torafk
l2UFQ3YiH5G4c8cBPtZjNbTGiMZMU+t2oGxKegt2Z1oXGY7eA8D2CXxe7C4zWf2A
c+lsUhRSys7t94ZScg275iQ8XwDK4kvFxBWrUsQYNC1EEk8M6XFJDYBiAiWecpid
vjQ0AyYUKN98Sy/r2PhsQRtqyihbFL53/iT5G49BDGO7wh2pDmntQbO4SMPvgWSh
Wu6WBHk9j19b/Q0Hbq78UXzRaZ7/IQuot2hUChEyhLRXoNe7deGfkQUiD/qTW7r8
AKy8nZVk5xjh1+AGAeqwRmlQAGfA1FzdW2gl1dssG1mDpBn8GNrdKptTp5at+ExW
ChuHh5p39JpUqZO72eGYZIflym3J00MNJklKfb6UR5KzjnNqNopr4Slk4a+t7/Gx
8Npg/soKB1ZuZZFHLo51Zf2Ig7WClF/JoBdsLv1ftdOR+DqVh6WIKgzCeZc2sghR
fybFzVsHfKFU4Sg+LZVB6+nGfizJTjFtNMtMkgmggk2QhyCba/5Cy2KQ1W/7wPod
`protect END_PROTECTED
