`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
grqMMuBsbMWO2KhMrXMtWYferHUwQKfKw5NcTwLJeX+u8jqEoZvYZvznHnP1WTDJ
gGaQbM2mKvkS4xVnc+EcDHgyMQxswOA5B0e2iQijKARsrhbHi6kWne+pirIf9f53
SFA+E6LVc2XWPtD4IKL6VB2sRcT/ZlLbE1/5rYbgWbRf5qx37PbiXzj15CGk+1rL
Fsi14QxOH+/hyf3eH+HgdSMpvKZ0qaIYUxtLQQh3hyzN5FLfCmHlvvBbkp2StpCZ
BJxpRtFVrp8071F5NmXiechgimDW32vTuP31e4tJCYSAHWHSnJBmbVriO1f7XXWf
G2zNfnbOcN79SIP/0R/czQJ4oH+5sSRrzQei9o7o7Zu0lncKG76AWystb7bmmew6
6OM3xv0vhwAQwC59I3p8RxFmak9xSIJ6lPQXLtzpICVVOs0MdBFx+iZ81fMpAtz8
2KF3yBEFOGKx4v94EyN2QdQquJ4t6rOdVhAtufzt7OyexRe178uqX1xdzzWEgwv1
lbEX45VLFwesxLifDc3m3MuaWH3xD/WPCnzTJOyQh5PhplxN/926IcH7sWw+8MRV
FjTmaWCKpzCIHzy+s0YhxyYU5GyunMvCtvVL0vMqNM4=
`protect END_PROTECTED
