`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zRa2vuDA9PTT0yA31Ddw6vN1K42rWCBe85g46dNDmY0tXASS/Rf3CwGpjkC4fDT6
Npxu7numDzq6FMoVKRIAtDBSfQIv8GwYgxU+WSrnDArg5Yc6hwUqOjGzW8PVw2X+
itQUYGdDwKGSsE9TmMq1eYGm20JfOB4mdBOo7qgYRE7iwtP6eYiy6W+P2v5EZ3Lk
K+m/PFgQadCURMzcYMnmoSVTqSjMzRbAD4ZpVEUy5Lpya78WlN7lS5rrcGqiHiUz
E40joXo6rjCCKR3GQwk9MnD94gSOrwm3yaglyN/j4MDudQubU4hlzUpa3tC0t/1s
2BaW+Bsyen+93XcvEZ2ByLlPaKmuvq2s29XGul8BIMgcgcXoQRS2AZu3zBPOrc0F
2zHfen0qw2zyQ0DhV6Sv5tOvBAfVWdh0YkfD70qCobJj1sTrSwLEUI0nFq4XP0Q5
dsKj5P5XuV9O1CSCKcODKhFJRdWSyp9hSlEvXoopR8s=
`protect END_PROTECTED
