`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODdYUgioFouW8qLjrQVk28bDo+PJT+8vOhqMOWePyvKEDnpxRQBpvx4HNid/g6N7
mA7b6tUC3hmNFepwUS4C7jZenBghm1CTHFTKaNq2GY/BK+gz97VSOGXl/6mQwKf/
fqhM2hQFjJMUjQyZIYUAlK+CT+W+fCRUmKePNRXFmaxvL9COxGILyI0pghM+yF3J
my//YT7etXgJyprBKYVk+3eul3BPYZf5qfH60CbL3y2G8QOHzkYbYPBba2t63/RK
gnOL6vbcxC14enMI8E+PxcgMvBL/su59F2tScaDk7dYvziAXv0MKaWYrwDDywbt6
CT194z5YJuD3G5+aauIMGbOivXisiUFQpvngCc66NoC7+Y+P8mI96xhNQmUHgbrw
8U0EStPFweuYfyqJ6l3lz2JNGN1yUWPdwfsbJ2BdZfQ=
`protect END_PROTECTED
