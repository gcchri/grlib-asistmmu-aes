`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bk9yWe7aa3YfGTVgYKafPrMSDazsOykab+lFsWU9o+QU93tMbR5UooSMMt3xgOaU
Ggju/oOMt0hdxHsA5/qrM5DDE83v6RGpFJda+SXqyPkqi9vqJdS4cttPZD9KHbJu
XiXnFB8CRhHJbioUv1WXr1kYKy0fsXej7ZW0f2d/mq+5zrt1gauWL5S5kOE+nHA5
cguE8KD+pG/P+j+QkaV8sZxnFK7o/Jrbzgzyej7Oa7EHYOTUllBRGq73ImhlTuwI
hNux4id6cZlAm/pBiBKPJEhVI3TyuPu82GIpNcfw/VwjjqSpSoUGG07gZeVuDCIS
HgT2TC54o+SKxxqDSEfy6JZ5qyQ0QKaTqKqzt8tnzaHVH4S2vjcOM6p4uWqLOGKU
Rkf9YIG5dwCzoNfG0d/gw6z5CrHhJ7iEEc+VTZ8lyMhWJmZp/foqKIRLlHyni8zg
BCxAWgVzOrAUF9l2L7AZugBCXkxE8YX5pY2NavpFIBY=
`protect END_PROTECTED
