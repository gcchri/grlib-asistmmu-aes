`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P5NW3vhP3EZuj4H/S0uHdyAZ3OQ+JGTuYkc5iAVOjOKFXBwg6YxQh4WyroLBDIrI
65kW4yAMohDFQ89mLgFaC7+YJ/wYF+1Nk+AnAfvyngHWebMIopAL5EnN/cfOfZge
DeHhifNkL8HbH22pX+8uTvUed0u6+nAVEPDippwFP3gVkhxCIOHn69KBYJTkqlZS
hyzSF2Fv/hSLUjtwcs2+HDWAaFHHgG3f9tYP5QzU7p9Kt/vYlm/TpYKmJ8dFQDhJ
pT8RtCQFl02Ywvn8dxNn4gvsTEaQH30G0j2jrVA+ou0vjA0OC4QLRoBUKKDpGtKF
ov+HSKZTeoscnO6I46DfgAKkBQbsiPIPoUkbKC7BzRPRKxkqYtsA6L5oIifwK2bq
Komnvde3OctSsQKGi8gaJjRJNxO9C6tP0ywk3sGVkPk/kYhWXiU8AH9oOi1x92Ch
ENcgsfJULkjYjvJtoGutVLL8+AAUP8xHPJMiimpKKKKljIEhuhzMTNQ9/TUd6uvR
ZR9wzEhcXCc2+LwgbQgfreFZ9mrYnbDgq0i1YU/u7hkywLBNPQd2mSSxFtym5nNJ
pcATbAVq64KXdX/xtZT6ym9H/x1hjA9ROxfrN3uwsT+Qf8ER6wPIFc4LC6IaDkSh
H1jOCnT+ynXFyLrrNhtcsBsijgM52+eH3q6ZIj0On+KltytenKHpcm5fI5kr1ykB
staBui4L5UuG+Ogz7IxOzwte4c4KGxYKsjKf3piYnDrbdLwj+WNwwFKyOi3xSxmw
bDzT4SmBQHeymDfMy8ZC/unYrbEQvbvInIknNmcbzyateufqV7UWlGB2TrBxm6OH
rpqeM1l8rYxUUj6sDE/TZ5323iA0o51erkqIKQ3ekHkzlJJ99PDZQLimeRNXeaIV
IL7TLYkQ7YlbiCLkYNm1XQThtPo9FOsUTtdfuwjLOQLC+dXCotrZE8IAk5TBHIVJ
5WjCpHtCnKMNZtUP4leasij9zSgptSHvC9iexxDie3wqLFU9ZLyDT2TgtQ56bjRA
MTWORm1SNBvPRrfiA5L/2zLZ4ulRyr0G3k7RgkuhtddtbmECQbmVEbWWhI6WAldp
7oJMhm+492B9klL4k1N9C7x1mt0JlAgcn0Bwz9fhgROCGMlirBP8kv31UMw2qcWY
Yr9CMhPFD9n+ql+ZN905HuwpJGlCYVp/BdOEFrmiLlpFmBkGJjPmfVfrfUqdZa03
+e4LtCc4iqoX6kCCZz+j9sAwn6tDQ+A/du9DEwqKHqgfMBKSbV//O5wYWVCMY+2b
sjkpzU+7OVS9nIvKGez2goOSqAL2fD1mlI1aZQQ1nKZLyMRP2K0WkBy5F5rYzDpP
Ghq7SwSp0OqUVJVYLsHQ/fcR3HUfcuA2feBi3aCdGgAa8Tcml+p5bvBbZn11OFbm
zywwOIlEM7FBCKVHT+p305n1qGTkozUEyuC8oNfYlS79clXnka9fusF/3q5rAUA4
nBLPPTfMwn2hePnjQ015XQ2eAaAHz7tt67TsnWD87g3K1HXA+TclbZ8t/ZxV+Buo
igD8rm8Ktk60xsRq2DY8ZmFOROjT4ACwe6UiD4OczJa/+vIupP68gJAVoniJf1X/
rtomv7i3ydjWFwyM/Uq5lQ7C0fg5XPXwLxY72rRvSOPLyf7P+YY6DlzCGXT2Gwe5
wTv2Yow3RaiG+ATbBb4Vz1wg37OOWLmmq4AD9DbgrHC/tNu8LmaOsMMck1hH8vya
4/bZRnZ39qqVn1gEUl40xg5QFUpJonlMUbjdt5Uu/s0bVI5COml8Gz7tUnaWKvbM
8eJ+mR8YBPqz0RY2Q1lZXfNfjFTih3V41KUFFRb8aUqCnc/CCl91QvVVW9Y2TmkX
ckqU5W+D7HqshqN/CSEfZVkzCN6Jn0e13GQGt6qidw02YuTMsojburuTplCIDMFX
LjlkxofUueUkpbzwRB7EKDAJZD7QR6XYECAlWkPi98yN3Os28hULza2QI6b4p7Kt
O1PfjRlJ0d9TvIC4cbMNAMr1bipvayYlWWaG/ErvTHewXyudn8KREOncJ6VIAvOH
TG0iIf5+irms6K2+ypUNb27S5swFK7rvWpQPE8eK7jTcv030mFdluduRQdhZcKgO
yS2zNXvknjO4zbHZRbM2QS7MJTypMVi6X/eOE+LiFTk1+1ROansnE8sL1+4u3QHo
7QsKMIRGRjR3fHlsB+yAwoQwgIbCrVBw0ARkqz3B/jpHSIQWrmtZv4NOZTeXRiXS
DGr0l8amofzhMjRBaen4PZUUCs7r9kIXheTnCF75woJSkp4EYXOjsj450E5FQbmD
oK9J1JI9YGk+1PAMk1sE2oFmLjPhgF6IT+phFEgPX7m4htqb2UywdOYggF8uzF7B
DS4a1CNR+Vz8hrddcHPkJCqBqZ+jwRkWlckgTeyeNLlsrfl5xMTvp7G5lA+BlmP0
Kr1iL3Ylf7GT0kH8QDXdUrquV+VrK3S9P42937HHGk6WA5Sh0kcEKb6bdO6eAfsV
HQA/Iofvu4RrdzAnKymSqSLo7srQMoFTk4Xio54uYNWJ3p3BxeeiFLYIku5QKj1D
pcVNA4YL6/G167SUotMQhMYxn2+5hcKPfK+Up85PKOejpVQnw8N7NkLUK+qoNSGo
WQJcY4yb7hlQs14l9HtZ6aCat104Z9F7vRX+T/Zhy3z/RgEfd38epXqPZXr0nJ65
NRDzeewITtXpidf1f1afGbfYZt+TWUQbwuyPUSCuacK6bpYsGb8JsZJb3Z2pVxin
TQ1FS/FbIDJVbdLLbvtcpuO0hlu8IaBXL2wi+XVeDc08j6jytZRXjoBdbPM4O9po
d4LB3yEYyrUNJmiwH8oRCKsxD9fZrE60Dg+jiRvqa5l4LY/epvK3QmBHXmasofNv
AxRNfCpJ4C4SU5UOEeoXF+V1/oGVpcGdLSc0EG4HPccC0TAAwY16U2+spJBno0+d
kX8+wjCzLN7o03xeoeRZMRNjENKWI4WrDbCKCKzlHdjEeM/E+ro7mOoYtzdYAtAa
QhDoU6p3L60+jX3eIvHP7Q==
`protect END_PROTECTED
