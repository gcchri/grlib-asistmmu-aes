`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Mnk3Ioedw8RRH7RdxxP7FKwjqSjRfHJSY7nHZIlzu9Z8WFJnvPYe/sIsXfcCerL
yuPc4+1iRiZmejFl7ngPjnnWVaqbR0T4C2nmqm3EbN97oKfdLr13JtwoyFK9TqEk
pRHlcyXTss8IoRoe92wWM8d24xWA/JLjdopSdQ7/HRUIdbZtcCizpgn7bwLsf1Wk
dGTabTQai8Q8v5TzGB4xLak+OwyrWhPszJCDoUMaBPwUzTUpmfg3yoLBOFKqkBOh
puQVJBr4QTAoTs4/NPkz6Lw+zmR0OW8m2Dsg2TqP4dGfqsddeBF48BOeGSeccRuP
pHH2gBFF+0k4g5AdzUujD9VnibuFD9LAUaB91vp44ObrYh3KxuhYO2sPBV8ZH4za
fEjeUS35CvHEpa8+WK8yPF9o2CIi2biychNJ7S3GV/KcdDUk1wf491QKs/rY+iJF
yw7Q99Jm+o7BtL/L8x4ImkJF3NLHNSAvBHiZO6oG+Jo70BWDZXQsUUyE7divWVGO
IVqF2XtqWieChIZpOTuimsxQneo/vPmCfXldMyIKtgrMchB/TZ7P2niuye5/dVNm
mZwj9wG7ZCYBRcmC+Tnba2PqHuiO5Yx0e0QmtXfr0Dmz25h/XL7b4eIjXtV8ZyJO
Zh1kWywO1cgwdNMpxaXvPpk6EFs2cEatxiurJW7zrcIm3NUWCs+DEBuPhR+uUn2k
USFHTV0tuPoL2EgpCUepBtX4sEZz/pdHIs8yRbixHTuIqYcp9zNKLov1Hx6RHqCy
gincptM5ju+plUNSsA1pCblPm4bo15Q4uLLSHNV75UbYr1mQU+fH0V3jdnIebIdN
WIxXV++3iRFOSQO8rfhd6tpeBd1S0J/N7QaTsPyCbJbIIEavpsjSxyR0mppL6Y16
1xOPdPOqlh7aWHgLb4KhxmcTuK/cZkQ9bFCRv/ovfAePqSaFreY2K5RQxqpDBz5l
`protect END_PROTECTED
