`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5s6BJy5NLCzyfQw6lDXRKwT8TJ+6X2nyN/McTk/1hEEGGgouuMBoLV5WAfCzimVA
eYj+vNdMP8y0M26LlDgjOWOmDgVmc5TAFdfr+G6D1eRbkPlAHWdZZwsF7jht7BQJ
jvuChqqzYoDh/X/zHKSThycV3dD4zOjyW8bhDPO6icWwE9L4hOLOREKYEhmldHCG
1t3oTEy5iwqoRBNEobnj7OlAvIWAzGSbeK93BLw0+aoVFDwcGdETxUFqPnQSQPlz
Qr/MReyFdgSAQXoKPmpTIwpm1uDASwAF41KriOaP22PYpZyqjnw+8NY5A9vKzW5y
XDkj+wJNmFrBoFs90MzS/SuOH62PwNOAeB3R5p2Me4LN+1CHZV7+tID1VrkH0kJJ
s8Du6tOsCKnxvX7dPvQz0FmqQsMCeXAHHyb6hFCxB7AZvqja6d25D2rFnh+1VqxE
TRQJV8IqCbyAyXn8/8KMoi650lK9/6GvLu5Aab3F+XvxI88hYMkXVoGxaLUDVjIX
0UjJJHhofgQXCV4CKe7GnvkSH5cUtK3AdBoDcM7acfTfL0/YVYmRnskIUcx6MTwc
uVxZ+TZ8Ungt370bdCD18YOJLOzgr8ST/2GRptOzFCp+Hoq68mLumAXDf1nimKTV
7x1jYaTosmvGKV5MGn/UnuowlmGBu192s3dt+BYDc9sFBbdio3GdukZEmal277xG
9DNH92WVnEJbZqvYmE7u1mEk1SbvPK6GOXzX5BoFnKZP9bBrsHria4+1ANAmqBgj
huB5BEMjtWl0ipwXP636pb8GFZAcaKAPjHPYLNyjhIG7/uyahov6lBXlLdWxhW9c
mM6weCWumt32mTJR0XIiITw6QYFJkIijqtrk8svo4TnOQNp/q4//fWvIBhT/coPK
XWg54qKtWU+uJEIRqwYvPUDppfM/r4VAoJdtG9wnbwSIKeuqCe7q6u8CttmTpqOb
oxdjuyzt6euKyyQ4veN24g==
`protect END_PROTECTED
