`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ohfl37oCi0TrLQkzcYg9GcuEwGaNo47iV8OQCDQK1oDlT1z/Tq8SAEjtpkUagWiT
6J8LChqxZ5gw5o0jmLvrClEFy05NnUBeKpH+VSJlwbGUapAX4tYpB+SClhS5fZ+H
ul1hClRwCIhfyZtHUtlcm4z+RqvpxFhA3AuaRtC4Zi44EOpRbZiyoIpxFaj9gEZv
LYM9y9FgFAmaXQxVszv6zmTtl/lcV2JunqC7ke3XCRgk++kY7Y+gj6H+j9cXlPEQ
9IY7iFXQG1E8qhUfC7aKZO/zzjkgvc20kivJTEPHUVLaGuIrJs+6J0puvn1Qn7o7
TaFpBPFc1eIvY9QnXfqkaHM0Foc+knLCcoF23AHyxOy6SUxeOZ73HAfTQa/IqvJT
eH2qDAr4w++0h89W/wqQKgp8sWHuEJV64AMiG8I97Y0=
`protect END_PROTECTED
