`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TdkpCt31lmsFJR2QfQg686a24udzYY6wY8C1CwOBSsgMGPgEqRL4FWEBrn/ShrSo
a/GyiMQCV9XRRlTOMehBxgedzRDvie7C+Ye60kihuqLk4eQ6eDOF5dzbildU46ZR
sho5O986qtYdCbKYzlrLRG0BW8cvx/ZtfBWpcFPFtYCKmcHOziTd/oQ14FyaOmpS
BsS5kVtdaO1SbP7V2gi7jKjHB6dt2Uz1oTmKM/rLA1Cr2EEBxlVJ41ZF1ckphyle
q/IJ5dG4gHl4Rmm9DJ9FBWxGmQUGaDOp6r0wF1Ll2ay/ZyjW+0Ecz6NZpEImRiUE
K3ikAIFQ0ZF8knbGbeEEFbPggYRib+30BOZ+ZjHC7bDXCn71y26e6y/DkmeEMEFG
ydp6KeN3cVftW9t2XwBjLko4+P+70Cit66YKmGr/Gn10rgwTS0gpgkfc0QH6/Wsb
cQLoTMEqEgnsyNlXhCVBTJXSIG17hqvKMwRKxZzwjqOC6OwAySAr6eYbJI6R17AW
`protect END_PROTECTED
