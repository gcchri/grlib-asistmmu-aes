`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ENXHxMAtNmAktDaecCJy5YZkfQE9nZuSr6pn2IYQvl6hk4fljlqOebLVShmewOlC
iPSK4ML8Y4nYyZDrxl5cuRvOHztUNNrr+vND4rLZrJIbSiPkz/Pifhc1v6t+3D/J
vLXEjteo+H+OtoIznHUCug3tY9sBoGeaaRbC0V1vg+JbvvIpY9wLeulbJwyWlnkj
73EXr3H6tpgQKkMlGhOnb0aH/OfQyuGPU+T3uc15UHK1AbZODaBGDoY07VZGEtrY
YE+TlYQ07HCvwyhyz2r/EnTJ1+/wZsr0BjtfgzH1/j7X0VmSWZ15ydXhjyijf2Ml
3lqIpesKrkjJ9yu4i+kyvnJ485w5Q3ocx3fq2O2z+54=
`protect END_PROTECTED
