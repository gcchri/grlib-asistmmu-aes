`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
40G2wPrR9OkZHOzjfVfmZaFfdB+PB7cAdT6FxqBMGIWyficgqWTlf56Dy3PvGTRa
NDDgk0UUBxF59785hJbTvCeynoxzIJkFgatjztNY0Ds1ylDHQTmGtUYzzKv2USzT
AJNFbNxTSreEiERpnikz6YTfWvowyj+5CBVU26YA0ebJz2r5LKAMR9AaoiiUjKvr
tlA+0NDF/SLKx9/476cn9nLlZfxDY2Yx7AqZDZhD+zEIOfs6oFXu4rgsbjleMRDk
6gSbxPs0mhvPmt9/z3U59dBrWKVcoeFwRvUF/f0DUMb4v+uJ1JP3+CrWf5NWdTyb
H0ofltazjq4WQDDuk7IFBBdrDxMMDpFBEixbq3jcamWEUMYxMV8kAZUJb3i263jI
0OYJOQREf4fM/AsxDwz0tu/iDjsWRRnkIGakIjy3tbI=
`protect END_PROTECTED
