`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9ZTzImLCI0d45AOv4Tb54v81e+WrN8Z1tIi56JFMBD07pH+16Yiq6rsvK+BiGzQ
jbXYCrxJoLCeaMFDQ3X7IRCdTwpSk0Gid0pgJVQdlev8ukex8d6hAWYM0ZkKz1kC
CPgPnJU4EecYnfhF/25VYUCPiybeLEIfZG5mNhUaZml+rsNl7JAc/r94Pobpwj5l
5MpZm+AshTOjwPEiDatCwIqxhSuzUDrraJrBoROwAuqwFUAyFVE+o6gI3YWlO/oF
//5gaQ4GLwFnJnvD6g2NqtxSYZKG6UjhH5194LqVe8+sK8/M6Fd1nSwhTf/zis96
mYw8pRn05vuLjbVlf2Q9nxr4ogLYnYWB1N5aTK83abNoejURZF1VzCbnQdCi0yQZ
krIBPhTid2THZqAudouZ6nIOd8W0rCd9f+2dBWFFpY4MRDrRdBWQsha0lx20Tt7W
`protect END_PROTECTED
