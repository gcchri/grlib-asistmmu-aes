`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkPNp1EIsd8szFupxqRp5gjTrPYzkgpNGZYuRO8bo3fRCM1i5Cp5UnvhE5iif4Aa
Ovb+66iZiZwymUuTbE5KCYDuKNr68N7noKzl7syCj3t6nvCytayQ2q/2ginpk7Ck
NNIqy9Jqwr5ytEw+zrCVhYD8t6QnTcb3901nXI33HRDTU504qTm8RLxGczBrdkD5
baTUJhFyynBGLWtmHPZlNM0cZMAUJaMgrFs3JHCbaywYY8dQ0UTCqdntWWWQf9fb
UcPBBc+li3U67T2Qnn4Kap6qMG5x+f8f41tEcZF6BvwuHJ/hTsxsWj6XgPffvs+0
vCSNYLJnHDwk/I3PRazw45CtoOeeNvi8+EyaFaLsrg6fxzA2ZLlSr9vk8oLPpIaH
VawX/cyUyoVZlk66fe9zJ2+sGAy07LGVxzTX7MC0bDjgXqDDaj5SO4oIB2cKDFuE
VElYUl8HSmxzq5tGWUruY9Sexy6VXLcoWBMDxmCJPZQ0ZDGcSF84AC3iAmWZItF4
MZ7008hVGUrg/wdc1tQcaZTsBr5XxMzQj/oyOxKzwz+DFRbSGRGQtJ9OF1BMOckY
7isfN78OFXafCuownnJ5o5IO0TROz6P6OoNnjSomXxuzSpH/XqNS/eACltblF9Qv
gVHQrki5KPjUf8uwdikbN7kUPkrnn03OCriwPDM93p+D98AMgGCzGMcDrFApKG4P
E5wQNi3xg1+gUvXTTwfCuwXzkmB1AWwM/HLG8qReKhhRhjKYdDRcYYwMDyK4nv/B
hM5xkwpUyY60Ncvy+r/MUN56amXE4Zzh4N+3dTNY466s+7M374I1fcgqYasQKnUR
/OOj3zwjXEVhMjLbXMXlTlmP1QaYGuNF40vdSX76JOBgNhIrB/LfYvh2ojfoeytF
cNy3M+CQS95CmXyR6V5lyQl3+/US07dry7hu7WgSWlwq5ouPMxwK0S32XRcEYvrp
kQ2nGxEameAYP9GrlHSQelwPnrJxVrZQB32sE9nnuFRg+kdlZffJHo0oPXTokuYk
P6KjTdimPB5nlxoxD4R3LbO8q5zNuv03mdx02wYEyONeLDfM/hLoEjVOro3JRx7o
yh+4ZXvQPpaNvwHp2JmPg8ZGJRLIg1Tt/qC0yRLjSBf4rb4+qxk9/m/KhlMi8liw
PiUaEFd4aH9+mxfs0ORcXbBMmwXK1D9pZlJ+aUVvGTlr2Hoi1XTf4Kf7KHt+Rjor
6WUEGUVnRr8HkB61X64xGR5wO9HjJD/b6GERXMcBKeZVNfW4cm0UsvliRUz7thsk
D/uxcHtV2MaeIKsfTEboNvTxFaj0bIVEdwAM4fXL2BSZ5PIJRSYPMoAwNc15MKj/
qsOqlBfdNYM0YteSPqRkoQdTec4wCSHNnVPMw9cOhgWq8uDaYD62Dy9WITfYIFLQ
jSdot6mngPzdo/GwQ8vOM0RrToOg9TvvS0CvHLeQ760YEUmn1FgGuxPV+6fHNH71
ApjiyQRJ92livEgF7elz1gouBrxAchw99bSBE4xgJnd7emFFa57/1lmCXJHxekjJ
Td7w7SOWHDsZGwoRkFoPqVJPDTeqkzVbkjXJi0LG+MvuxwT/VpSFo2369bvC2/qV
xKzEGIVFkUMxUTkZjvMO3OyKLacecN25NO3mNlXZ9w27AMgS/10nfJE3PbN8xkxJ
zTF6e6+TX0FPIA7FIwrCBxJicRhH192qPOWaitB1vMJ3oIGXOyvXQJF80p4gUMwW
y/grAiRiUiMLohqelY4NX0lWLDFpH7GTAtHAnzamiYh32Ihg6sMpLnRECIaPFfZz
VZPeGlLX7WJVgMythjzrQ9tf4F+ILXsUGic9//Ob6zQJ8NfN6xCm5m6znzqR9oVb
sictc8xPpfYV6LgAbTtfr71GayxZnkp0cQcouX0iJxVNe2I3SaXNWze9DGy4nM5x
MuTq3Le9O83oNbT1hXELmyOR0OWdLmP9LsRmAtwoEaUPVN4oT2oPGNVytbU3YzZB
wlCpF9407A9GfvaiTbhMadvzaRk6Jtqco/gGE+4tEqGIlIofoZW3zrymkw473nhD
B1YRO3hOPTIFxUYAfpLeJzmmwvvXhNVVSVxEkWnx0RNg8wsw51nm6jULcRKBpAgK
gkx2trJuV0gT+dMYnOeAFg==
`protect END_PROTECTED
