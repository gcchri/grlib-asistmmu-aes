`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i38MLF2oqEptte6u66/x/NX4rXoU0fR5W6yJ6Hcp8eDPX/VNpPCHeP1tPgw1/ier
fMmQTQjYYT7NiJDaYqN99lmyVTRucx2H2HB6Uyq8757vYO7O3ZwaYAXQdovuAUSA
nphLkMRcDqsvPbv7IbcqduFo5YnrkdJjqXMBAqqmI57kh6Z2t2MsdxQJN8COGsXm
4R0aYLfLZ5SkHfMHH8j1Meg6VUt3SL7ae9HnUaE/la9xceDe6sFc7BwjPllTXpcV
a1bwaromEOTVauYAw/3NFKTzlIhRR89RqakWl5KwPg4=
`protect END_PROTECTED
