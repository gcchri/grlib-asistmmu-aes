`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ywkStIh0PC3yYJS4zphcvd7xHTK2NhvY82hyuEATqQAYLZxLlZKf1xbxAoHjSmm
5su3lUGsqHk5TuWhPHa4/iimPkYtejBJSR8E3o6/IYcIob0M/8nuVtedQ8L/iUE2
rKBNZARjA04N67WQyATzDdoDodUKp1s7HhdJnCDZt8/JZhHhYDPxfAuKH3UKqlV9
Kj9YrengPOpbhXfh0qwvv9V72LWxgeWvuN62InxcRIWlIVq01HqxJmsFfyc7D1Bm
gOshT3Ix5xP1140RwkRMdAfuSb2y5nKa73H0CpUSkXGi3vUQXCl79xp2dEalWpfF
kEn4n4Mc8ZguAMpO+Vws1qAgJXOInvCk0Ik3g8ACmblC9QL50q1iJxs29U627AOL
RtsK01MM+ATkSye7Y+aXRFGPRNHAAGmNRC5Ej1LY699sa+fb1EYvszQr8/t9M7UE
GZrk9AEBcpIkfhKgJZNFCsMbL5hY7jsrK62IijN5JpS4o9fA4JMaKqo982oey0JL
Ab8EVyeZy5uXCqy0EV+tCU8ihF/E1fata2VEok2YGkXFlUB5uF6w2r8W1i9HUfLW
FODpj3OSBAw4u1acI4ooHcatMskgdyOQrr8aftk9LPkW6dEnB1EimKw5V+vb2j8/
We7+IzThfDss1BbrR5U3t9QcOyY45o0bf3hDcM6kFDoJdaHXEWhY2SuGfI7iIybE
`protect END_PROTECTED
