`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6Y3z+9heOgvbQM8kw4YUBVqL36KIjhC49yWw3Hbg1P69OFsVSnxsGk28BnsExaM
HozQQgUqPxwjPOburmg2jovIN0hchdZPX+Uhkyc+iBOMxc/OoP4Z4AAPGIUZg71J
dzWxRvBiNnOY9/FJPuOVbHVQ8FTF0SoR2Wmn+XAzuLBVxgKhmGpFdCGvp3a+0R3j
c7LCNlLJkC3VJWIhFTDUjifnrT4HYUcHwFE7sTDkE/ZznG502CJBWSeBQ1pF82uc
c1GaHKX/LyGfiLgX0OQBheZuIi+64+N1noUFjFEAmBzGBIwQ+yeTTX0Gb+KAJWYg
CTtbV1fv6XzmThaKIjTCcOL62iIRyds58VcPBDGqBdtO3UkFTa46LA/rB5866sJk
RsfklJiYnXwCFXJWdq1cKg166tIF4e7Dsl9XtUO0ALM=
`protect END_PROTECTED
