`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rc1QW1LfbVaO/ALZ2+zsW4DzKCRJZI+Ri1zXzbc5PqfVL3LUj+42QzwqTLBpEo6f
quLoba1Nrqd87frcBTa/jeA5hDyUMTiv7Jh3qXdallw5htkNotdPJAcVRAHkbfZB
0C4mMgOYaPbDQHPPChO2qVZ8sBVH0wdykIf5CiDvmdz1V4rzXUUGtLTXR5mjPokY
787oi+nfZamkjv5kHCawCyXdPkFgMccFEPfpjIlp2hTX+lbWLJ4vKkgDWkp6oGtC
e8xP7nyxuSjDWru+I1i9av136qLnkaNb3x1LbaadsMkipgMJ6MOEku8BRpPfsCyD
oyxL/h69Lviz47+KSQ9SQKq1pF0pE4Y/UcOeh0jyRgcWV6UuBjfaDX1mk50FvsgN
C+D2H5R2vQaoS+y2ebq7hgX3+NyYpxhSbOWWXZ1IXesO+QHGk+MIZOuHr37e/raS
KqdtpaY397RqUH3jsElnHjqlIsbls+T4LqYxJlit+XaGfdLxOexCWzPTzlCbPS2E
`protect END_PROTECTED
