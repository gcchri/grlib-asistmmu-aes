`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bAD+3D/YDikEiFnatBjxNy47IADRAP54UY7DSIzggmkveF96A6oCQJm0C/5gqHU/
PN1AS8KkMK9iVyyKvCRVHPkVtCCwUKr1iWm5DgYTEYsqxLSOY89iQacsPAkTZO0S
qG14q4BUJBvZp8eIhiCIurhNEZmpyV0qJtOrF++T9MDUMDkjNuO2WXE8ymZZjYZz
/EkNEBRS8rD/x25FowdtbLkgVh2ngSnp7AbueURAElxQpTJg+/N9zLSUrwdfC0GP
QZt8obfT93i5ImNQYPo4ayi87uhkif5boeehtNd11G2dfdEC/rPi380evVBoLYed
ON492RuiGR0CyNC2FtjQBfP2uOActxTsOnm2kDBbCVB3sufXNghGHlONvHlXUXvJ
bG+EXjKiitIdCfoH5sxRaQqgdZSN8BbE9JhNOqrRfpjNhTPNmdC2lzaz5HveWuKC
AxpHgpg2eIWE8tc6fbRFQ2HPdPAka+I/sNr7dIN2Ol45VpqAK0V65YeshCrbWWZD
Td4pOWeZ5N25v8ny2CWzAPcCMvt+GJZF5IHzEBW3RYMdF6oJG3T59jsyuaucPyn0
UBgciGjpqJFeIp8xoIEk5LCsfY6eW0F3B+/HxcDkBVbQ1AcjeOZy4aPtt3jKuXfX
O2Fjdm/tcvWTk//LDzFM6X7aT78z7DKe6BUuO/y46cTCgc7/Vy7rI4vXmCOZoIEH
vj+MZtSQypf0waQmAnwIGNAs7GHPnkv2XhBWA98vCE9M4BZmfksO4f5kfsweHc8d
hPAKbjz2sVXXuEhzW3pUTa+1OObG8j0pLqwdqIGtKQJQOfuEnhaZ7+IHS2k3uRwx
84TVN8B05850xO4acdvCn3b68A34qiD3aldxwRa24rjBMYs7JUkOi/2/hPHp+03s
J+Qbs1lZluTcDZQojXgs02LIQA4aphqbpyoAuSthqJFYkOOSSWFDwmyE805/Hco9
sFe7r9JY5SJIGiLGPU1jXjZph7ksgynzb00/4kL4DidNPUsPslhViUvlWOVlKPIh
wafsdj2SIlPyToW5mPAHAaSDGjJ+NGUHxX5+KPXTfYBBoB+BcqlJqGvSLv0JSAEO
746k6Wpr74nnMXTpBHITfz5hShZMaZb4RjlTLygPyc6xcVahxYdmywOlqHS15alI
fKLvNgEqyPADptyilZE1Fm+5cUvF3aZd1wWLOS+GLyYF8sb7EHhQozAJDSgo+xgE
ujycRXYcLoPLmy7I4H4xeMgKVE5ym7T1xxnSU5qRszT01j13LdUicBX7dLscL+47
nnwvPynvVG3uQmjZFhK2NWP0GluXKY3RPwjxM0PoqCYmw4ZIaW/iwIlWbLW7BVUq
muTkdY0F91hoKL0Gu5oMQyGHwgfbaSQcJh5ibzTFckRVvVL29AbgdT2yft3sP6eo
r2DBGm8q2pQhVBiw3pt0rIZhY4aYlh7aeAC8An/h3nhT8R7WHPZFwkhk6V98W6PT
Os4S4QUctE+VFaO2edbre4Wx/Gv3H5QXJwX10TFzItEBQvucmtFCgoSu4t0QsE5/
oHu7uZg+9EdITG/V94WK9uYxmr/6WEQZQuSaC658VpmAJoxb05xLhi2aKurjpomg
jwuaRWIsGK9+HrhjT9QyfVcvL/Qz3xwlLHJkcCuDORqSIf2rGBXxqNb8bglCTe/6
N8tG8njtmXNaDcg60LbjcQOEloNP1rRsuUWcFCjjbWnFYJwuMPbpn3hSteNFZuhH
CPdso5MBhK6wBrgtTzbWSNHWA9XCw4eBVtzhOxg/TwS/lCgY5zBlDNZCmo1zPQeJ
8hQ3fmwXrCio8LemQwmMLZRRSmhMLX8oFrKMt7pL2+dGIQTIQwoMuCEyyyN+4chJ
3rm3IcYYBKiQUR+DupkDZYg/mou4KH+HYUw0u5jNzodPk/sPonVTEbk9pWN6+St0
O1TdBvQ7J86y4uZTKirYI38QjSisLqoBOLzsZmqLPcfxH6vbHNiFQnjIWjm2EgvD
sHYe6obi+TYQFwMmd9mNYmC3n2wiQ8hFd3tXOXnbIMDhK2MC5KidYZsV9tW3DYvB
VfkGkTPhxzUaElh8kvJ6I5lS0M7YIu4y18eTwurNk6G5dhXTTKSylrXdnBd9pDPG
3fMtxLYuS2tE+9Z1kht5aNSLyAqo4Gc1on51xotQoNI770jT4G8o+pxiJ4qmK8fd
r0bPN8X0v9NE0gVSFcbrz+hNmfX6CmLfrvf8ty7yLe71uBOLA4G8lz9mPLeRrPpt
ojQWMKlquYgUcakxiIVd+3XelbewjUf2+EKwoOIBpHVz12T7MEMxILZscBy9DlIS
hWtI/nSZfIpM44aGXEvzipYKSKn2dpB2ZA4QVlCm6hncQiUyAbnuPjQ+/Q19HF3v
`protect END_PROTECTED
