`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qJC8yrqcpa+VKQtKk+HpzIMBRyVoceBXM0AQjB0BlIizF38+lISwqogMOHgRpyUF
q9YJWROxslSI+1zSWhfYap2nFJnnoxKRECFo2SE4gQkjoHSCCWePEaGJdieS8Ixy
68dTHU5sWO//dum/YVGyUppK8bdcMYwiN4fptOsjOQNePafkED+X/wGaeEnVplh5
62+Vxv26ELMWuUYRqREQneeOcgC5BNFRb7C+Qt1sb4n1DOcJ6bWG6YdHc/VsKT27
2/9TswH3BCNjPBAclIOX8VwI7RpS6tEAOfDPTQeejqnOVt7u19AKC3Ir9M2Ppvt3
riPgk7JUlX7paVtnl3q0pihZ3uVbo4lSnLq9KxbNLdp+2pepz4uimcOdTDlc1Uhu
CYgw6SwWx4l+ZZ1suVTTiSnHaxTbgrqAnE2PNicNgljCXmn2cki+FYwCtQgrZ7V+
U+DyilRbCC5+zAzUA/23wa//8Lg6cUcPmkYCSREgFdYIzghmexdyjp6XA12FjDMk
2PYKMDbebavQUbB98V1us6rhS23dLsrcEBwMqsrRPm2OXPTdyqBMv3IkqPrV8zo7
s4V0rHGARxzWv9+5QuTef8wqY+8/tAmgrBdPiVEEqgUx9iuvKciMCX8bwd3ARDAK
FtqzQnjCVcWeCWE2L1i/ylPCfwtKEvNxi/7JOCpLpQoQVft78x4mM+a1ovgJFtx/
uzo5o7zq0OlJwXr6+gz7MlAkpsRoiPSMPGiqTL1AwFbuRraVCfDOo8Cz9uGj7kGT
bHuWCgXUhLCAuu3rtvZt5689TVGCTID6jvKTgv1moMchQ8RXWamh+TbNOBY88iPZ
NCa3MYD84nVtJPFgLxz+3LpZWgFoOjqCemQ7BKpnUXEPvy9ZB1lqh0AtmjjPilcB
rHJaV6QkWQVtHvD65246e2gmFF8Mh3gGauznI6I9zdmDHr7FJlslx2PJf6qXvqgo
8mgmI7RISU0Qmz5OCpm57/Dz69R1ogzRISBTn16r94zVveajj4SHvBstb/lIiBig
6M//oej6jCPmDfHrfkOOrKD16N0TCP5ZDyB36EFoNw3vnEG8tMDJ/C905eT3pJEe
0nCAEwC9tlBeopr75h14L0tC8VdXwO8wiQ25jfsZvPaLLJgY3K/CVWe3w0benz7o
lv2EpN5Izdpn/IXJhUwQqJYruVwsowkjrEveSVnAb9ZDhy3frhNdvPAwbv8jciZg
rjKh5VoI+2GdhvCr7gRyp4OamvURMRV5g2daO3UXvpXhgpJKRp9pRd1o/HfaF9FZ
5C49dCAFRDoIQ0L4bQTWqayVudG6hyWtyLs1k76vtxR0uHcaaqy7YWMYM5/5ZDXY
ExTa+rtRYedNxOCPk4lqNTpvyGnib6wl/ePVLKoGZ+rWGY4BToans2xGA+lmte4D
RwWDH0NoZ5Wt/nkyIxbQ9JzjmTBPUkL1ZvzM4uz2NX+3lLn6+ORyKrB0YKUl0xlt
5PaZI+eLTSRRTMH/v3/ra+qsGaEmnEBlwTmCYJnvGKBYhw5miBaoNTSKZQ/SOtr7
fz9QhFeChyr++i5eGBjY5QQaFCei+Cgpi+wIlojUeVEoBs1NUOxO7ot61n766zyr
zwUSxuXQIPXh2JNgtkAx9VanD9TQewjlERV/CuwsRGpKCt1HXM+Ak4mVKPStEQI/
yhV00ExBalGS7xmw5dr8g+O/4LunjRlTs3PSpIp3RIbieJx8bv9t3cHYdzTuzGfE
vg/cIFG8LcG6VrjdxFDTfbvqx4boliaPH7LRg6RykBZYaBBeCzj3t/Xkf5cmV/dN
zGDXJ9jQYT0rlq9bqUleQeKnpI7DF+ea/jgnuqdjpwVcCiTE7N0W+1QlgL14NdRP
bnP5oBIIZqlHHVmZ9FrXybhpM3yIz19FlIt2H+GJnkFGAwZ82DQenJPJzFyS0Yha
ux63/6Nftbs/d2AiaZtJVnNb4XMsD18xqWdYWT29iCakrWvKUDK0FjXhpw/Muy/k
W6YbQkJobAi1p9RWFRgtkX4SXb/KvvAbICE8kaiJy+CeNXWksivDMzPni+kxPwU8
hI1/qUlo2r69STu9BZxx2DaoZf+cyc8xGcYirHEvvWoUYg6F/WBi0VFK/294tqWa
kd1rBUH1xZu7Oik1IJHFlmODrJQYWHn0gIQjaBIR7b9CqdayRnU5yp0VAO+FieK3
9Jwmo3sAE4faT3mszZ9wOhJlhF3MIMODMwPJx2dMJ8RHLXH2zcas+EVNmiZOxNS0
dr5QKp6f7SitT7eoIwCCRsIdzH8suqCdGq3ClvDdB4UIi8HMydr8+XoPxBFBkb6U
NwmvWbTzwIJcg7Iziu5iEUjjtv2dRjz3bsSzuUdsL83+wBBRjWuTg+M64Tteonur
7lu181P13fbHyaZiyX6nyOzIN51z0cHJD3l3Er7l4ZenWVlxZVJripeeSUdyiCED
IqucU29nUCEdkKXObgn5arW5r7jfJzDQymvqx3Iz28dVaUkCimWa9qD6jVIjWOnu
dUvWAP+WicNLoDnTi9S/XG42m2rn8mJjuGo/TIBzJyvxsDYJxcKEwqId9UGvSXvv
X70TtS9NveXR6GHo9YJbc+336wBkid3MVl11hZoMqEjca7dkPWHemvJ5413pvVfh
jLhxTXXdnmC0K09jmE8TDx4fEzQnDNGwqq5m0fo2AWr63XfLGcuLiHjr2uECxNxr
6I2VmRnaoa/dmIckSm25bJzKwSmwVT+HqA8TAOBJdxLNe3Vxyr3XBlsk64Zl7Fg5
PF8tlfBMCoiOGTkeIL/dsPSwdcqmFR1noTqAhxz1w4z3Fs7g+AaxKL07FRHy34T/
oOXWKdmi8tBC5+YSEpY5mc/0U5FIFCKkYngkoi58JRaSfOEers9RRsyKnuldsyTZ
B6MFqMaGIX9VygaOBLlaaMrFPPBsxBPgZhMcfwAKz37DmOEhz3MkNqI/vsfKCNV0
ciiBUVk5MjGyXm/85/5kdeTiNYrZDta60CY5TtrdafbW2A9xQ3zi1cljhtIYrHti
i6afxol6+qc/OSpUHiqTgMYi1TvacMWqfYlaWFeoVaV9y2oLjrO2wmtNzYixBnzw
7xOfYhFcXYU99wp3ZNEPXEN7BKA4g1GJSvwqfwL22XVA6v/1YdU+z4zprPf+It1o
psAyeyKX3FCNSJQr0nc51v9wpqAlUSsEYcX4dMRTd+IhyJY8OXZ226UrKmYjZ3X/
xt6VUBNg0NjYs1keh+6XLdudfCEKfnDUIdwTm82l3gARNNIDH9VgwhT+jzOmTZCu
4ESDSX8F+YfZFyaZHksAzrW3SvO9fdwLmO1F9YZZ8TpBomYFGwusDlVrFo9y49WT
BKPITQsHyf69v/MzvBBQJV8A5O+3QAcQ7Fxp3R9u9vP9U0D5mjFbw15CEJCvox1B
bkvcP4H/8MBkt0sM4lBRASiWLI6T6x/IJ82Tnp7ESvMQoNAzHrBrLR03ez+PhF8v
kwZvRTsLCaTb/FvwZYGNrTNnG/JBqaI8gffw+ANZ2pwvSwyzxGD/vSutBlYq25h5
5noc9nEdktloAwUS/0doJgwWPugJdbdmuA1oTgHx6eKJHGBWC+NdU+IVogNBkvnN
nUJAQ4nJvCsVEx7O9c+rcOJsHPorciO1FLnm1Q0bRodvrIqy5GisS+wxFEnBCoLd
k63tmBV3o+XJ8e6QGf73nXaDgw7RM/3IuoQ0+2+I7Ywc5cYrs8S9ICT21avRtGis
GfgIYT/qraWe/slK/JTV7o/QSkSDkxtJbVMg/9Myo9iYoUnF3ukskUu0/L4rwg0h
E11EWKo/XnkyibdLCmTL5oOTM0ACNbMjtDqdy0UJwNe7sqojyidFFPQqOSlmQwHQ
U6vdNYOKBfI0isWL56QYZMjbNBEvx7XJqs9eXtFKN5B+IE4xxvO/vgVXNbQ2CrAj
RCcZjNlmop0qiP7iDCDpG7dxHUvEM11FEeW7SzZuxMQ6Ngmk6fGknU/wVZfJAQ0o
O8X04jsN3fBmjh4BL7gVQRtTiXWtRf31MjdbhLg2PB2FyWJ60qCqJqdgUa74d3cH
9H7S4wmAbsNr6vBuJH/jcRyVzBwSKbn90gM3Y0abZxtPtwPHw2EVvr+bDvYv3G6H
DNNODLxOIzbUDScrj9wSjRhmF/NGZzC7yb+Y3Zl2E5owqsao0YUZ8e/ZPkDnqupZ
s9sf/H+lr2HoOItHdQUJzBCK99I45LLxdP+Mj5ABq6KjO3edRbzLR6wX36AjoCzw
+MiiuOPURZ2ju6fEwtDEkKbpfwsNObfEKTE6Cj7a8PoOh43oOLcAOqbREyMjI8AE
k85NmByeIfGa5T6djflHMfH6dOKwDFiRqQWuhK7KMJza+F6zzAl0rRdJTuSVxFZj
RkFGLyzXZdjJMXREzP8JzaeniA2Y1TU8cvPogAGxO+F1fROAEe1jDaIA4rIPVQZ3
C6PHHd6QM0w/R+s119Ve9xrCFPmHpH3KjXWfvGBGei1ZuNncFPSjUGDKS7fYsReH
yKG3mL6ScCnL5xVvFfCcZqfq+jllcxyy+rRMuVUT0vWvW9U84DTGgnIvtNj4VGbp
iqA5rVSDhJBO76no7b7aIQNIz6mbvKCmfCpyS7xN2MNotNudHmjBxA1/4hfxvaj7
yhZvqv7xuqhrKkoKHs10Ie2Jw4GenFroyvH1lnPjK4XaEKnJ0QyccTPeyRz5M8zB
8OYGKV7y2ZiZ87ClSDbHqzieORlOPhkyltQjU+40/gep2vrQWZmkXpxH3gxltFqB
ncrooHWihSkoHxBG2mO9oUc1Z87M+r5axYNR2Wema7InFMUubMiAyEf8EiplGTfn
vA5Z9+I0+qHkNhYo2tAFJ1taxJzPvcYd0lx/YgeajsD8kdxuVn49GzaZOu6bq0OD
om8lnHc+L80PaG2Eo4st0NEpjeaT/YwDIXq5ToprIjHPR9lgzzwZG2Juumefn/d9
CxA1iN6+L62ECh+It+U+UU6sRhV85dfwS0ZxWGSx1pz9+Ev9wSA5rvmZpRw+t1d0
RSGzId5NjiIHPPNGP+0wY1XmJq+hFQjn2wjfyr8xkkvSHJpjcCb4hgHpVMKT4DEt
J2Z3E9DYIWWL0P1KBq7wZdMqYKyUAHx3/BIcPYpunrySe6hVekePQOA05gF5EnPw
C8PYjymnXT4qE2X+HcOK9yzQIElAcANgWaH8+WEEr272RCebmFu6H9tDl8gDph3D
meW4T64KNkHSFhux3KPGeOhMx0c25ctBL9A3xJ0n3mqNV16TqVwfrRTnIBXYk+nY
RQ5DHEeVaxycc0RwOYjEzcWm8DWTZNlTeVYdNET9PQb9kjh3WA50bilWm3NdBMnL
6lXGn8J56H0zQObLwo3QiIfdvx+yYIwEc934O/Vp71xgEtUWArMFJPIEE0Gnnw9n
8aCPZgF51QyqxPut9poUKExQBMRmAQsuitaFhuKTyv4WVP1MeIM0v/Rbj0ys5KdI
D7mKn6uZ+uJ7zovMYfx6xliadrSqhBky/4P8/urgP0GQMNg9q6xmBrAWUmLW80ao
kEzguEzksngWdA/OAF+U5VMGcMBTPGmRHoTTBxDXSzOaPW3x1idwkljNP1wYqVQF
TLxC95ecyLpItN+hS9spDCFW3rX0SwufFWxQ6M3+XI3K52o4XmgwmSna3sz7hKt4
mt3jRPemIjdlroiiKFzVI8KefbjCMCpO21+R8xeC5aFD003njee8qujGvydT/34H
LR6LL0kjR0wqv77Axu9/otdipZB8IxtWQh1lfgoQB8iI2eZorI/0Yeu36ksrEioG
2Q/7FOMoX9y/3XGISQBBQzyZlvVOoUlAhR/VN5cHnwSDQi2NM/6kBXu/SO/Y5p9G
E10jplE5E8rnQeLhkA0AmHmBK+o5rA8U1AVdVriUDtQtg0XT+7uwGY+mQM8H0AyF
0VCMA3LztFb24HDFwjQdHd9NSHABHjs41hI/mwIY3lP0CRQh5zf9FPhS4hDukyPt
geKLrDq38AaIdIJYI4m9JhNuvbCCGxNMjeekhvc/voZo1/UYcJDAgZFiVwHkJcf3
QA7CgrmoW+FkeVZ6ohwAAmGVaKAaFVo8qfhDfppAVm43dT/qHiF+yN9qHHoJN5un
Imab6SI8Utlumj4I23nypobbJE+mavdAdoZXFO43iGyYrsQ839yCU3hINBx2n1+2
XNYNCdkXEkB1qOH8KH16m3lT4a6BQj1C234QbTIVFHmD6C7oBkVas75cE5cn3CZa
Zr1p8BoCV7uvw4BKR41jvbTC58VFJPFJCZTLUle55KfW+kDWfGu/xKfPmgT2bvt1
yLlKwOA47wZWcXmJrzcmbIOr79pff0e2yk9La0QLYlIFhLKROHbETjpI45IbMN60
NbnfuzO61LfwXcELheieppXhVLzFb736M4IV1+zfuAUPmFttqcsd5H4F4qNqy6b8
w9DTJ6zReg5Hom9FF+oCQb/EE3xKRD2qv85CBCTmEPD1LAlze28PxHJJ/+6wghuS
8LDERwEG1d8A06y816WL7+LeA1/AIBU3S3uw88g/YK8UnGCpAl0jAD8wQnEC6afX
iQniN3NFby+gCFGkLxOO2IE25F47ZiUDRC89nhCB8YbvrY5xgsZjNbBhcVGSzIJs
13LtODpwDO7+WfsUcl/Y/qKe7mKyEuazetjZj+YvXQvJQ0BNXmcVLiVup9boTWrY
dN7apKpxU/R1HdngPfAk56iL9G2QV09frNx6FsKnCJBt0lwqarq6cVDrv4cRUEP9
NNjNXqGN0pKCeTlLDg2KO/2ic4rI0rRn9d2XnzMzf8irvPXhtldtzOnYUXMEd9uW
eyydxpkCIu/FzC9ZYR/pBVyg86pH2xQ3byez3VU8im2yW9iBQO5jPTBjIDCJHCrx
yoi0wTasjJzjirYRXb02/MLZuCYz7lTiZon4F7t8ujD+G7ZIT4jDw6mfYPzDuG3x
m6iMwwGOV+vqLLhPkR1E9lE0XQFcZCb00rX2LL2UmNvwerObO/rF/wl/t/0v1Dsz
30egrlK/qGacnZLhwxo8+2mx51onGuk9dZzVa6UlJpRl0vCpviKcNvlBMnDKIkCQ
HB/C6QMbKRZoe1drg2TE8EtFtXxAxgTn7T4tNcTGXhvqMvdq906yAR2b70z0cZZ3
NQSbWghPE66+2CTVwLrwzAm3xatfGj6RRT2cfmVHUBvk3TTVHgAssWF5eIU66NfJ
uD8UoKwA/kMjdyxF+xSg7T0w1fz60XIHMVfk39RnsFo9+FIy3HKf6m9QS2Q4G4N1
lQ2eaoRFHJJqJ33YYKZvkosZsXGGY4VbDI36rMASVgsxv5xpS4UGGzdbfrx6BCoy
01dALYnZ5qu+NyVvG0JZDACqJ1MMeUGWJL7lSIiGlMl6DVz/3CEWB5ym2vN9S0wW
OMUSwYXhDM2CVh6WvCtAaWXdnTuul8YSyvqFTkHpKa1G/LlEC0FEiWi3bR1qP3YI
Jz0T5N72f1NcZrcQqGF74iz7PwqHb1+d9liRgt6pTHwEM2t7DmoqTAwXGrstEhD8
lstyXtLR98hvvOFg2bv7JLRXRza113K2JDYiVQq3t1LDm917QepYLcISo+wNPzKl
/eZ/WKH0VFJjvphgWFCUP/N0LmahB0KbT4aUKyW+IcUL0BeNH2RzYRkpOQSlE6Gk
Kzxnr2IQnrCtL9bo29qDIPQnXShFgIAWVMH8Y2aXuUw2eWpzq8uIE64bviXz5int
pEyLfipm0oh6IkmsM88mW/6B6y5rbFr/H2onyM9X4b5fSYNSWe9QQOCT1rm7SN4o
s8COL/J5ExJtT5CC6V6ej2vcWTmLBR4P886NH9bXKz3hJPOjfWebz0kAHLOcNe5T
ed8e2A14PvmvaHOCv4uuaGFQWnCxsF358ZhtuDodQWs+D/9zMEj7uJPjfSvnZUpj
78vUxcxkRAwZw/0M5B62146md7RmXzjz7YbFhgb0intiUsfM8vmi0kvsH/kzMaP7
EK8hjcwjFoPcb8TsWN15UoeL41tayLYZhmgnMtuYSMAaDX2QuRf8KRNBfUuL5Cem
zRR8/aNXFgAoO1RnkBHIJRXpRrAczVc+3edSVIdWBt9gzxXap7pLxWI0JbFAUEGD
HOUZBSWS3urwTKLFgwJaavjRQ8d7K6To9w65i3DMP7hRIH0I6wDPrFEZZHN0AwEp
jW7DNuwXwOODq3jzTh5wmFzDXT/xeUkKYOUPPpQlrF4Hlf8AsSsEtAvAbExl55eU
SZrJ+kv/BVIREBkEr3DgLg4vCJ0Pj5RGyIqJbfg3puZ5yU1P/o9w79cBjQUJS0XV
pu1KHBVHnEJuHESX8hnyFbvNtTXwrpXBoU5VGdbYzPMfVPffKY751CU7w4eEa6wy
bOKjaAbwlJzPKAXW2ejd4TYHvegyvH8fS9I4Fb02kYZ8kUaSP1pG5Ir15Qi1+DLW
XP8VTGY9/JroqovETM5GFf5p42QQtQmPD4FxkSUEnaUissDY1nEnIdtgoQY34Nnv
gYTIHedTKEpaA5vzd/2GY/PS1EduJjCk9SWqWY4K9Ld+P3NlEVCSeqiuusTqrMhw
xGctvRWGVq+Pth+tJxxWhQLPOnJZX+smf3oNVjB9bfV0t+czzeE+C5Nm5+nwpzB/
bXzjtHYrPW1NYBiqtT70alzLi0PeAqlHXQHjA4GR+PKSo9dN5H5B6K0bnn9L5PnZ
N4UkPZPlUuumJqNK41uOVtWXuuveJ2yi/uH4mNZ9wbuHNaP65a1gyMGhxgYGxMdN
uTF+byIpetjyYxNr6Lmqzi3yqmuEmuHlYb/11knZshkLeuq0681ShbX+JKf2p2LJ
Q5y4+Mjjzp4bbEGWMZPWraNNVD+ijF/S7zWf57gH2G3J2CgnokHc06lOhg4WNMw0
rh0BEgc3O6vUgOqTEJoIKT9hsZoh6IKxyBEXikEp6+6ltPWBwpwckNRFZjI3WcMC
fC7BJa0yd4DXu0fwBKj515YhCRoVgydNrxQECf3IPo9I06uU3Bl13qsALpKr5JqD
DR254BFg/AAlFGqxu4E9nuj2Cq1ZF/sT5MaltMPOl6hCGwYKgexbtHib/05ohY9k
2vj9uPUCUYQ9ByjQmoj7CwWLsePFcclro9FY0PX2HfUC9awNScBZ1Txv/MfRmHld
0gQGGKJVbjdh7xewTjxTEIGaOszzBsfdQm9XpTymRlCqPhSIenzfCAzQJOm5dc3I
ghBhf0C9rKwZ1X9B7tBBdbyeAhIGgyRt8Pm7f1uUfAIRLaE6uFejbd8fRvif/ih/
/NiloGQfVT9o68XsA9S+v3fcH18WW5RiwLaalMDpi78ilud/Iatmc88u9RS/XP59
/dv019EPTbzAccwix4dZ2WVwzC+JysTUyRq1nC1B3Q7OaSnObIn5Ddbm4ClJyuQc
gUFJxEzsghsEeVwQ4FWGHCJFMsJkTkoCXfAXISjFbtO/wB7VhV1U2jIkmlAivMsJ
hjbrV0WB5lGWHPcR9qhoY7iMg6iJIT0VeYFINLXE6TCA00d6DPllgTtpVe7gA4cZ
IyYJRk4V8G4ce06EhKzrHVyRuHiaZLGHlenGu5+1owwN+ROefvQ090DQmnGUMp+s
mTZBk/9vGaBmAkBmckhcnm5gjmyx7yj5TvS5a+KputkI72ZSpNwR22efu9et9Phu
0SP6OoBNqNV1pyAmq2p0hI0MbPYcOgWWJNFhHw8BonPpS7wnuMWFSI/kFxiPU7Gw
bA97zqAQpkfdlqvPXT17pejUGy8CKHQ6frAnD+L83NLQ/zfhvP/5SLg5IdXtEoC4
0sAg09YaLxTqFW62UJRyFVLlDgBt1oB4doC6BiUeHGq7cIBk4xXaVfnNc6gZytQj
tr202hdvtMBH1YQuTyGrTqGRWtgNxVVLGeJAICvVbVvDrISNwX7G+E91laEXEgiq
x+iqrSs2yNrN8tVYDwR9sqK2JA2BHNDKTgWBxhGiUVq3WAQSiLsxVCLpreceWA8u
62aA1fBEb/PDV3RLwj7gIMpBhxxhS2RKE4hFECthBvDHFweEZlJeoqZBHgh8SZPy
AH68qYh16lzMQZmeQhPIVbAquTzRLFXFXjYKVaUMMJgj1oOkmdXIKaNawo5yaPgv
QLWz5xWf9POoZn86YXR7koQLqDgnj96kNjoVdm5ia/xULsbDfoYfHk1IQMbPb0nG
7TAva9wBK/v6pkT3zEHVsAmKYB0Atqb7EsrQn0nYuAt/vkyoLtS0uKqloRIWFqrI
yrUiNzoiY+lnSv4EhnAEaUQ6hEvP7JYgJWa/jvF1NomhX2mPhDKGk/NwibNRNreH
FwIO1HqV5avNLrDj4Lt6Zyb1xjj0Z0P418pZyLRVydepUf394tA+F543Q1P8CfQI
pdk+W56NmsobrCA5EqAaue94ld1cklo/1Bw347WEF2u5nGR1bFxrdcpk10asrFm7
tBSBhCp+KX2jtQv3n/WSRN8JS6EGJqH6jPtfjm0LaqJ4dupW8TgIsMc8Uuh59bkG
S6BkqLbaWi6PlEn5hEhL2IqvcBP4zqwiJYibj8snNE9PXh6z7uXMcIi3iqNAA82P
JOsWPrd1rRN49gA2iR8LnWIJOCyvDVqvXjPHvowMDY5hsu73PtYqHGYpJADCw5M+
bDU/cfSMzzQEdQEoZzBvelziFOF3wv28mANWMzPOyVGfM4X7t3si/JuNp/EsNgz3
LyIqmK9JL28OEJLEgYiQK5IphZU0ehbf0/OA7l2N7AdVnR2NNk2UbNlYZd2Jyk4g
xdghaIG7a/731fbh8oKCr0r/JQMXUF3yTxqpKiC0Ssm5L89Spzl754uBJcVGC/sw
HXy3Fpw9bczqP8A9ivNLTON6cxr5tmPmX2G2GaPt+o5o9Nkio7Pvq1RHlj0xdaYx
TjqW3TocUcrYneUOvPFFxqaT3lJiIbBwOd599qDDVwYDvZfZ3Ef7IXzKQNADGctG
U7EgdvJOfjnbY4KikhiIa7P9DQJU8mhy4D5NOW7+eJfa5DFPv6faLDLDe9p9Eh2+
/OOONUIptUXSfRWthhMO/L+bCTkD2gE2VrAfGMagzl16udDnD+I0Ko+C2Y9NvZO+
QSOLrK/upNPkkBKanocb8CAPgcgFfB/c+OYcIKM3D/LTMFcKXWte9d20ZVLXlvAZ
iF9OIxC4mBJRJ8MPTtFCJ1fCKjQL5cPcstUAMm3hRinuSYkIf8KCugZrIsy8r/CX
iKnRkx/WvwLxUan8i6IQwGDSgRaGHeI/6kxPJxEqyZZVcdG8amC6J/rrsfOtSbd3
Apf9902/ynW6Md4p7UOurM1CGzTSAB9Gvt9ZF6QYL5J1DnnbxFWq68unwx3a0Vo8
+9Ch5ODJOhHVdwspZNbhqtAORe5NmYspWK2JqzsUnxn4lpSbRXsa7vhIJCu/aJx0
MlBkelHYiarTlka/wzbuPjbpvV1T7fCFsW5l6dgM6VKQLAgBmOrIEzcisWLFzFC8
0hGtetmO/4wtr8hrrHS4chcJVUQl08KsL20+iPuueAxF/pRUE7ixXfsXjToXHlAO
mwp0Ca8SpNcAdSqzGjL6ojLGRgV7Is0peZRFq8n+hxFLULJxL7Ci3J2EFOLVI69+
JfEz4b7SMX5IDgnbjysrOetJRiJ+7anWlAgBdYZ6G8Sqi1zfJ+NzcxFmQobO7S1q
XFcn+5mCq0Acpc+N+o/anR9gicbFajGee0N9cJEkStCggWTZsZrmuxA6fSujgh9n
3rsK+w4sSUxnN/WIU1NZpxa1Ds+YfGfdgOmzU2Sfkys8I1GWOICiElpyRYiOF+5x
98ea70oHdC1zJTsTfTlH339jK17MKODOGwoA/Tao+4zyOkydkhJC6y/PfO6+78Qj
xIoS8Ie5bNZnv9+15nmYl3OfCub/EJI6R31XhU/ZJcoJvVOpPAcDPJ/n3FvoJIvo
82FTpHZk8YCCuH3Mx7RiYVVvju6DZqj0Vdb5loYSWtkDqJxcje4WuTFNXJ4Ai6wW
ZE/68g0Fqv05/Zla5SW5gpvdoSPbFzfXuqUPPm1ePRteLcChgVt/yOAAvwz0aLWo
gKLqEfd3wBapiLywkqTbXw7TpTQfgkO2kx6YL08iJHpcGOiT/uCHeou/BGmLVZDs
u/+nd5Jdx4OBOjRh5S9cjxNKHV3x6sETXYVipJaMbXPpJAWtxbB5YUtgajnC8Mfy
Mrq+Ah12FTQs+Di1JHJ4hFX2Lb1gOYlS95d+lDwezfQwpkypDgWKBrWnPnjn6w/q
E3ugcI6MC2Qxc1TIE4Bl/K78uWTJ9uFxykINejZCyN0bUwih25EYzueACE+Ul3T8
L431YYiyVGFNK3xQF7PntsrvPZ6aJbUp/UKMJ4vU3hJHrnDuerPH1I1uzC0l6P51
I9P7dj00FdeLQeoQOWo9y96kfrbgQbZu64GyLw1pR6NtkL+GwQCTj2hutKx4Yq6b
mx09JWGAJxt8+asKobNBmd8yFkkPnnuXT3AITyqRQ8USkSm7bByKGjec7IFNJ83Y
YvnhLBMa7a5FaiokB74MNk/0h0GM1oKYwgLslC7tJvdO3DXAEqdqW0gbLwascGrm
wcv0MZk4tRqOyKysCyGAulULO+yIH9Pa/hExqmhn6LVuetx6b04uFNeLTz/o0yeo
sBATVITGoiarZEu293Fh6ja9fdXm6IDZEfcz4aF7lVKl6nHmFzQ7tjLFbxEtIPId
yQyHlcnEJKYV5ck5xrOuKotPWYTKJI9e0hjZU9DU1JdlxRl1IfbEiGThQxCoSUmO
iRykaLbLALxVUrtrZ6nlZzplV//5cN4oKGIMbKvB3hLbLBOkS/Y518bt8HZwDxGH
yIdB2GGLhQEfaJdNyTZ3E6lwPfBUxQeAlE01ek1guYTjkhgTDyEOd2jpXV8/a2+7
V2FjF6SSJbj9IJQ5AsdEMoDlbOKYpPGcrzVc0ZBRfpwhgRuRVs+48h8j2bkOmnfq
BbVq4bOSncRRgq9olNpTJiRxeaQcr7DnI6BDK8ZAiyxu5az9KxfQEOYdljQkhjYe
RbmWowOEy63HVdirNaXg3+/S6QgGU9eLOJYA2epE6cO3WWjFDduAJOovXgEnihrm
LqYA/1lqjKh2rqUW/Jqh/pjBTgrOOUeImXAP6Qcn0vfdx5vrcx01PaOtp45L4bNX
ZcapmIPic5azYJZxoqz6A2jk2BlAJHce4GKwrtJVE7omESG35zHOuXj2j2OO3pOc
l2uT409le+U6ynZizuDS1mDcgaz75vgnNsfhYxybojfdVXYWrc/e5msJCB4anqdm
S4OORg3XlNUp4QdoirUYzuxaIiQ2AymfjitHcwSSSw1oge4z6mNtrAfZJYJhKSxV
2LRfS+j5X/pVExeUUWGm6adkAOpTynV4U6CAlX4iymtHz0l6Y17M1M7Ntn/ytkCK
jxdB1HW/GGWUz8pm1Pn8Kqg0snx3+WunFzA+0vSiVUKzBUS4FBfIHMYIwFbq1ELj
MLCs8uiK5fof6FsfKZR3Tg3zKXc0Hw2PgQn9h/q83CuodAW3KJZ8QiylqTGar3VU
O5LiK6giaDzUQ9Lwj+u1WCHgdwflDxplawqkAK9UON0wOnqY46Mjm9DDUnPVkK56
XIBsnZxIhEBlxnMiUF0RTpHldmiDSsAJ6f23crBid0iMjoSc3YnBBJYGPUI1sPUP
w14wG0jgfsZo3qWsKNng74HpNsh4tdozih7EvSbYjkngnigXdfdGcUsJ+H9i/Mm3
ddIE78CC+XQ1Qin58z/o78bsDw+qqjm+L90O0XT1t6y2WewmZ3/Vf7nWAqCv1ZMw
GkpHu5AJsiJfAe+q1X6Fc4eiM2pqm/NfGQFBUgpBpvot4LAnRySXNyX6ps+6Go+C
BNUTUqajJhqszOL8QLmtnV8SClKCbqMu2J6/Nv4QzKa/BRdABjRRxRZZtEBQyKeU
4kRRDEm/6DsraUgt/i6Qc+hIlKl44PSsOLkisK/Fb5ptdBLBoLPQ3dNZGx+o7Ie7
05WPBzECKI2tcCAbxOsdw2sUeIr50FEeSejtY5LLMlkIThSy+H8UPvDu00e9mpKA
1pWaN5EPMDh3octBWvJrD2yamqYIUDvPPJfJGj1pIqaVb40y3L/C26SbZOyYx9iK
Np+Kvq+uMOUs/TENnpWZ2rRRCWk7m524HFYAExaqVxG4vWqN0PsSDfc1Qtc8Te9n
RPxyIDPb04SApsq+nL/lcEDdIeVwAlDAmVciKkgEQzjXyqiT5AU0u1TK769pZlnK
kdsmnGDJyy9w6Y9W90OndFshoyZYZjzBRAGEdIMzWlB1f4EUpHdOToKalBwNYP9P
HdQJ9WciM3M1mTf/kTgzx2oxEySloQVjtdndEQCFs8geaZ8IBJgosr6gQc9aCR4w
8Mpwqji0sQWHSZuuoWRrbmn/riuR/Eh81Z2aibXePXxyJtuGIGYUfYBT0FccuUM9
KAKPqCzRvIUgmYcOsSEX0I78Mm32CPAQly8oGATvQ4GJCMaA94XCTPHNEPP8verl
QokMJS3Y2E9wi59JejavwO9v33QvEXfDW0hV1hCQ1NS8UVXBU1cQgcxoM2khG0Tb
mxHfa/PCdL46vUJ4UP412dff7W9EtuxDOlTsc+5DBP+GRQ1iBvL02pOSoteXwJ2G
UNOQVeCMJbFXeSMwMCKH6gYkZKIsPkmP0uHCHGNOhkodYsZalObINCaZ/ANNsql9
OD4Pv6yLrKL4QH+XGZJokwKA2FmpKNq7KMzJp2QFtRU/ozRX/oolbU96VurzkMZZ
wptNUhMxv9Nev6/Brlql4BffKW/4BIpqnHu3filduMbADlUXQYYlc1XRqqmp6MtL
K7T/h3pCSU3KMb1Sj1fy43ZzfB0PybKWz0JURTmIMhYllOrVis+6cFWuRAtOJ8Ew
fOliioYb2IuLYhwCQDdtu84VhqifWcVdrIBitsINvV9gTuRwpx1OsL9NtufRTxU5
RoDkErMgoOrfMtQBY+JxGquFQ6Vq0kUvHRpba07UAdZfItZIWWnK+FLkqb8qGvXF
qQGJx+GD2h+Yx9PILHR3irTgFCHRh9KsBoGr/rQ8Jaid56weB6TQ0DCBeA8KvWIk
kx1QyW2zPsmzqgR7PS3YN1D+p+oKUh14AYVZ5veD04C40cqpJ/C2HC4DtuBCcuSL
o2QyYHfeoMTWGskI+4agRetmRlBwN6ViRSk3TmZWwGxmr/aOeQsib7zT3WSR4mfP
SmFZ+SBpTwgfrM91qXXpwEohKFUTpj36f7hL4SFpn0qaILKnSIP51A73r6jGIDWA
THJhe9GlEOkB9iIJyUEPoePpOrk5wjf8szmzi75BSKJV/QvwuHrUCISLUiq4yIeZ
tqkpi/Lg+ZEw5EN3WmmKvpOZ/5OteSK+YJ4vOqJsEi1cl6+9oSPiNsSwFiOTVFnN
2A5wLgVpGwkGmn9/ThhxkhVvVjuh+a1xuTUu3KoxWjEgoROjy+T7xJ5C6KtHuT/g
TlO5mLU8CxLTlfqOf16A+NiTT6hgohDjJR0rfvkNo8TEP/A7RbLXsEv2eUNuo9HH
9/uQM91Hyb5UMCMmlxHJt4p8vgQD8Dp8cnxP1SVXIf8n8K4X2m664KY4t5lhhxsm
19LZ5DwwKVnAIx53Ryg+OYKvxXCMwz42or5vOFCQpX6EZzqjAJTy6f3tw6H4698K
dSxEdgpdKCri/w7OT8HOeUqVJVQu3oPz8GjzSlawnZpkaizS8JB/ErJgbEfZhvar
1eQgPfUWjfssdZ3/XYz2lr+PFr3hv4IMqTXwKaimAFRFEuFvtBeAVWHt3PWCYAoZ
TjE0hMbCybFX5LCe2228vJMEHIVrPRGIUOo8IaKgLpHZCxrCoWpr+d+PKonW/7FI
pOS2hLF6DnUknkmU5Ea/Zq4EBPcdSiUUpIFIP1N1/A86mrJj3f5rmTImY/eXXhca
Spw/+DKaBcB+Nt8KVbYYUkDcXM0bJbP632IYZqrFVCAung5mU+6j2BRYefGuOC6Q
r5DCQjQa3t2qUQGQN6OgtmCEFNeCTgTOmz/Rya3fr/EfvOb62kkJNAWHBCEVs/2N
QOHBxd33OYOTtrNr9I576+Onzt/HFwliUzAy0uRfMM/W8C+NmsDgKNR2wd1sBnb2
K01GpoFjUdW41GcVZ4/GzGHrhzECeDa0iuSbJYbYcAOZJz26RfwcR9xZ6wWOEt4t
IQeY+YkVP8ovYEjLuI3I78/xKbC7cUwvwPjH1B6rwyobGY68sSExpCgeOXUmm4+h
yGTe3AgwOd8Up1yURtmGeZgc9HHn8PEwelGGLix5nSKaEEownBRQv6klgwbW/kYE
hQzfug9/kIHArDx3QmMG2Pi6e8fQPJ0YESKoXrI5w62wn9AdfIcniYW1bTHphNqh
aF5R/gqPnH5CgSe/Ly3EsFR+/ZKzOoYFyPJeG/JwAlK9XqdYo6AXD8gT8nHhGYz0
mTCEk5UxJ072FXGDl/I2lAZ2vOb/GQD/0VTpsUHQ4G8jZvMB1jmWWNrMUxVEH5Vg
XFUxoYaZICHiNIeQ/uiodYIoOq4s198TyDnEGJ6Ism1FklPJBelq8YuHyvkXHAA9
8otMAJQeFxWGweg/QNrw17oL14LW5SPHFuKnCOytIAvnGTB4NhGhMMzp8A5Bp8ot
WpNTQuxZfP8ye0fm95Gy1NYiTcw4K+MI8qY+jebxEk88wVxNnVbLljHuzV6PSvms
Gij92XLRu6hOWditN9iUpxuUon9jfjpx9+6f6tRtnmKUKTzXsmZMNaCJHbVRIPyk
V/nOfBfqdJXU4um8VEADghPM6YSX9mT+bCxKNvPc/lPUjZTrMC9G/zhj6ewNahNT
M2ZgiK8rd0jRkL1jy/+V7sMuh/kOrAg/fKIOYZuOzyWQB0EtolCpw5FmTgWJLVIz
mHuAbkj55ooZZ2SvrkmgezJQFjS9DpiHRkDmW57Sq1NQgWj7LS3j5ipiQ2LqImRO
/KKiJR8Hboy76COqquRgx37AR8MTIW1ywEWiKaUjRGoqn0eA+rzYgmzDotbshI3r
FgFU4wEM6nFiKh4TxKDj1S+I57S7iM10l6fbZtLUCTV8ZxAtoxTrY2gkj8Ww7rNC
VUOwL3gHhHfsN1N4EfH01KW5vcxAeAvbyTZh7D5F1jPDn/xVFzEzgmlxYVhA7LSY
qYLOSGRbaa5Y6i/Va5o/honAzvK9GnVANRHI4DTedM28WzaGPgiPz1YEELypSikv
/D4I7XI86VHcfR0VTUODIyChcymMGw01fhEGJV6lC8YRSyN+lIfZlYlwOrZNN844
/PbbU1HEafV/vkAXoNOZ2NkRKFwc5tgClA34GKlloe/a2oXrOz7uFgajjOUG28dv
XXFlcp8sNjmEGfX/7Mc7SpjLwP06Z3muhcw67NjBW26Uv5kb3AMVG+QZnRj53X2p
O+XtChtH90j9yBnajhirnArjPxoXRFhpdxTEGORJpRgfEIOV9UOQgx0YnW7DtiGs
glRDPT9CtukZJXEJ7iN5Y39kwvAHYV2DRHa7OxmzOSpWP9BaWN9yTr5dKJOwBFyi
ehNido4CMuM5DzUd0sIuEF0t9Jutc3uUkjPUPsX/r8Ky7p3K0pqkRhtTbFW+d/gf
hDlQX0cjCKJ10yhg+bURNhavBiVxWqFb/NDvueoO8A5idR4Vl/UuTUhstmO5Wc0c
PhdlkUoJJrlGEHKPYzJxHxgWfso13Abf5F3sXBoa490K6rZDPDFJYBuphJjBxCPp
z5Tvz5IBQNSrSj1SoY6Du02Xn/PuXzNBoKxhxhh/Gtcv7YF9BkAP4MB1DB+IEbfa
Gy/3pTJfclNjixI0E4N/fZZ/HYBGXzzZmFKXkjAz8AYQjHZMMtQFXSd3a+whMPh/
2Qa/u1Dhvqvof9A7m8C5QLRVq9MA9SpVdekz+KLux3MK8mAySKosFrDtJ1/OZnC/
iQAe6ydJnZbfhx1XupiFHTAj9hTDdUZUdvrXPUnu8ftpDq0uHzoLAsZdrq6N22uG
CKD+c25mTmuGuhpd/LzyG2jLu4+Yxi/W6BNUaZQYIp5AAWELpmr3muJL8P9YRHRT
wxVul4/zSUmzxTLDG73JceW6fQIP0wA+7gz9RsDRkfLtP4VBX9baYyCgffiuVSIV
VHW7B0r9zq2Q5/U736rk1YfC0fvAHhEmg9KCDJp1UMhHgr62PTf/CmmdhRcXbF2A
iNWa8cVyRBJ7wB13UnGoMxYuE9+S6rvdHFU0TM53fYaLvsGTWo7vgq2zI+Qk/rBV
WFYw33e3DI46GfJaY2G1/zcFryVbqmqmstFmd+ifbLiBjKponrfpc21f+yg4s7ku
QVXFBkieX/4rZYMrSjCh13SC27SLqSLmyPncKQ9IJMk=
`protect END_PROTECTED
