`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UjzO2sNa4hHgiikNHVODbZVHS9kuPIRsJkXG9cWr3gFL1XYw2mRq9epWJv8s0uZc
xDINeA7aWYbv7yZY2WpHiTTtUZZ0HDVYeBa/6km7/IUzwbCiEx7aFdxY7/2wlDlS
sFAbUuZisPK6vQjNtAxCT5MdJnDxCmTMkSOaOkOv9nx2dgAY3Agnm7keponkDHmt
B8S9OL526cIHS31RcRxArzVLOBtig7e2LD1Fiz/9VnB/tqQG8m4vZqYL8/Pn2mPE
TYgsHfwHaOoXrzDxi4Klg3K9G20AB3pa2H/R+nLfYfRelIKMZq9yTKYFfxOBBrOp
cdMKte3TwCZNbia+h8qjMeHlLlAiZw0rK5pQbh6t6HJ5dtcxBPrP7CnUCjARfEjh
FK4vk4ZUwuAB4afoghBB76TObqBMjmLVSYtJ3Ql8xKOMyObKSvpQIdVPZQe3fRCQ
uP9Mpm9k2GlQJWYdLef7ILcwmvwvADNWXG+tZJ/OLcjhq2tVqqnfWoU3EdWIMLDv
kdmabDCs3G2xe1PA3So0dudsR/QU9bwrEd4hIe54QzuSvgXiYLunztBpmfGulBde
dNOndeSDoA//WDlY2Ue520eL0wJ4d0kMWhD4qwgrqVQKBAvHbxY0zfsRewNO/6Y5
Yh3bce7oSXNO9AenWOG0pZdy4NNXaOwFs8Bl+GQxUCAu+va3w2yjMYrBJkkI+uAn
qEXi8VLsbWOb1/sUuWinpcTPTe1xfuBYZiL/jydt7G39Z+zC5gOAufqvoGRc7X+Q
dFYaoG0SX13stuhcPFolsHW2L3pu7yt8HtyfQYXKNuUc6RbgnolVkRchei0GdoRp
vNSa0jZPp3NpyGaCxJTnCzEk5C7yXWonO2zgLBLOY2PSDeoxQntnRir+2W9qlbFS
d9o47OEsDBMOT+cGxrIsGs+c9WJSxjDiTdCSnHSjzIc5hT8aUY4u7zVz+tSi6zxU
C8/GHzs+0F10+TBBZWC9ct13uVHmJ6NHcKTV1ka00Qn6nuJ4f5A4RbJUrCZgxcq8
HPX6Fv4PYFYipgr3OXS3BRqGe9NLWpDmbnSIAAhIlwcSIyqJJ5GkrhE82cY8bL7K
iblcJrjthQx0FFhV173hjQdJLSm+gfkF0TrO08Vr4Vnx36f0rW606swc1JUh0Zn2
qT4KJRdwj6N7FdsFxxUPUgfrYQFs0Pk5x+W9bmAlaQ0G/BnUccA/R9+Yrd7NZH6C
HTqsUID8BMB+IZgK7onyVGbp548ALdEnnsqm4LcdSYPuHhkretP3pjx+hqiNsUHa
jwcCKDXASlGeNJjgd58jk1i7DU+E9UiNCWx7gbgzwQers8rxVqn1dai4wKHwMUH2
1jnZE2q2ocQCdGepqj3HBfG8RjoNUVbBcWHb4rktp8NWf+z1Lih0t4WT0aVzs6Wu
xnH5SclhkRfwZESfZ+ysna9Niv5oTvvx/fqoyqC3vuMFp0i0rP8tiHVPW+T0SJne
uXBNtDBRH6reNb6eF4tSY7/7qCiFHZKIRRCCHw5cf56SyF0BDO5R0JhdVwqhDtBO
R4aTbKoFrFTGGiM0+kOUP+ORdJ17Mws9lKLWFhQwW9wqvGtsZOlQuDswZPNWe3RS
Q8q0jetQwQHYBfwqYQM5dYvhfgCj3KnZFYGW+cTdZZ6sIVPl2pTIRM+0KPWaqGSe
uSyX2oUTCcDCqrGO8BnSXPT9hhv2ka+Z9e3Xmgt79ODAX4ihPB4pVS1u/YLRzANT
HhlAJyTBjQpKGHb0RSx7/D63LaoihW/M0BHBd5/ve7se+D7nHS5/axfXq+ex2l5a
9rXMBzOMeVlyf9aJ3g+2zLFtBi03+9q1VxCFhXP6fadegYfhvdqLkSUmewRp5ifz
0DKtk/pg+L/3EG899MubxbtOzGomaJ9yo1euCPOKyjJvOB3TukdN+Rgx2x/k+ICW
B6a9ATYe2SaOpogdDZS7Anc7mZUQN7rn8VYKPJdKTQ35QrcOEZ8yd6MAdqJVMXX3
cgt1jAU7gtZkX5lVZqWQ7bmVXogPGVOOqfsxXw87W7JHV7zI8mrXlqgj/ljm+SQ9
pdPSC+gEv3SlKVzzugTglgtMuv3LPgrToDe+AW0MBHFSX7VChB+/YeI8rioEhjJe
3a65PSu4/3dy4vlRHpQju/SYGcuDhy5QAaQIcpO3MWBmxkfso33OipA36wBjZ7/T
eYjMyUI6UGYZrTdySe1VteKbBrJKESZzXpLuRsgKyeYHs/1gNNB4lUEvuYoXDlJt
GQugzl60hqMtRRRHEgn2YBDuucbdOV+sOgQamf0YRtNUDSwLtUFU1V+aolb+sy+/
JBpBAyCwoi+3q/wP/siGUP+btY75QrH17DTOQeQ0kM5OBaSdsvUK6WZxi06VQ/x+
Zvp98faNwdJIWByDGlWkCvo+F5ae+6crZSZ0/9EdZLacA7qlAWTgavA5XaWYpcvW
9Ndhh4kGTnHpNTK/vq/7eSKK5DIZSJG5Aoiba32GVANmco1CIn0mF1azs3JZWX7q
1lx83eQhhbRMDAwgSNp9M5CnkuD+yL7he/hz3gjzwKqCoWPGQsUR8CO4691c6CWR
xFzVjySzYRZbwlbz26jKV6nK+zhkGmldBNW8rPLp9pE49XIv0RlV2yecPep90uGg
0zOxrfhwCNeLKFyI0KnsBOP/wRfHfDVxrfp6p8zhrtyf9lGI1XTgUsJOPURJFQFB
GbzSjndl/5rYx+H9fj73JyeBXrmQ/TUBvz7S0KUYJ/SyQhpwEiKn5u+lb7YUOChp
G62dOABCIVUlt/GJzzCXIA==
`protect END_PROTECTED
