`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sR78ptQnj5RBYol6f6X0uqsdm7aisoF7piLHfIqGu1c2Azn51+V2y4ox64aW1FQn
hv39iIrMAOZp9K9/OQIBRYsf6hDcQ7PX/n44PrUKTVDcARcjq1ur1X8TZ8ce6EwY
F3/A64pLsReyqDvVxX3ygqzr6KeIGW3+RdXUKxeBn7CNMkqpOivPA4RqJprmfkwr
XqEzS1xrG7dt3CKIqam635kClWFLZH2AGN6inlwggAVSwHiA1XGQGf6zMqR2CBQV
ywqls81zLlNVWsgqshcfUz0bEeaxeCFsVvJi/TeVMv8=
`protect END_PROTECTED
