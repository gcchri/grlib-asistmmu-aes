`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tp7WlSsEVnhpl8tVPKQF8hFyi3/2/X8Kl2wMp3clWZP8R34T4yxVrmbNIfz1PjcY
Pj5vemtalD9sKbC7rXTY0A6U42T6y3Xwl/6wIW1/rBIZxRw/LoFmT4OOwxIRK4eS
h992aOJ3Er2FkX8P6ef1aX41jwd8FgvlOjaQkBP/33zu+FZVS4f3/Uj3W/JtdF7m
6g5rlQvLdhlCgKSmzUVP848InvnfmARsCRsMbJyihqjYggJY6fIhB6a4Ye3MiMUz
af3gb9mpFl1Q6xe1oNNRTSrTs03a3n2HBLRaHMUws9YIYnLJpzHjeim6kmMeSpQs
fjMghP49Bfj5b0emO28MYPzYHQIf+2b+bsCHwI7KNJCOoC/remgk/zVwaO5rXlHQ
3bwUPC/OqoUd2/7aXDDxWfV1WVnWVYrbUMrSwYTxljF4xMkmcO8IjFI+qE66fzCr
QxoaZOiN8flCGAcdNsYMkjvZU+ZjjfQbCkGK9wEZ5FbvS1bOyi+yGu8/hbpC51iT
/AccoEE+k4jVd1JsiECRs9hDS7mbei6B+TdZt50aVaQKtWMMH//KAo4q5ELbk312
mqTL6l7wk/QiGEWE9G05NO+LqyYnUSC+z/eI9hDnQ5YQRL86gTRLmY8dOMKTh4e7
y8YP3uUky+jAODTdl6RhbeZkMrvZq0upLw7nCzZlECGsvRLsDYxXFAuBpaVcOq/m
RQwWMtZdgp0DV9jSkEc+9NrVlxTFj9jmwi/IBmInwWWUKUBYzwOq6D9Io2mLZrJC
UHG34a6nqMYN86VbuTx51fKZSho6MyQA3x9ytb45KmrhBQ0DkvmJ65Hrdpe7Cpag
G5XljRUr/UshAjeQsRvigonq+BR0+us+tBrSgYtuQUeNB97xv1oqvUjlB+u6y1dO
GpfGQ1EyKrBmUiXo7faLxIU9dI5s4OzYx4sU3/waEm7BHngCXpcdfyzH5wdTvCo2
2UpmQO3xOx/CQbrejGEO6ZxRnMucD/eAo6oaW0QawDptFXAas4ECVgM/O+SZBHO6
kPg3mytvB8Wg/3WOSX2DKIKOQa504f0CKYjccoeplyt/2jMhWd3IX4/YM5UpVM1W
eWzim7RFC1IfFi/vEZblNE+ht8KFGflk8KLS2Ooj5geG07662SRntgLQ39NeBj5l
KxjHJcHLzdMIvi/jgtVtPw==
`protect END_PROTECTED
