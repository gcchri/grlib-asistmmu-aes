`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pu8ULaUzoWn8z76TZDk8d8JtgrzP+q0a2C2w8Q04Dc4sx1eEpbIrCg2LKSo5LEZj
VCsfTM3+tMrmFsP2fyy2ThK/hxA8UXhSfaZmtJzepMpMvcWf1CvnOj5zaxpBVG6x
KWSYDdhB6weNIpIGoEU5jddRauBrx21QNZJfgQLIdZbigrAZZQWUU89AC7upv9wp
v6m+1RcSnj/j2RdfYQU5I/YX3MrPpyHt+Y6351Dc2z/56kJJBzbQWjup5Dg8oIc3
S3Fg+ntFHNVJJIvZisjmBthy8Fq/0jINg0cgC5SASpCSqotfe8DMzQWykyZyb1B4
SSPSyNqjN9JccNbO9jbfPP5+if7t9qrZPUv8P3IkeWYYSaGtr6i7ArPaC6Jv1rXD
`protect END_PROTECTED
