`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XET+ps6FHm/gXQ40TX26FfcbqloYmJC2SBJbuusHBzB5TS+jw3Fh8BkIkLSWNBB
/pvOkDZ3QT5TxX7k7Y8ieU4NSzmurR13X7lIecjxTjMuKGnWT0MktQkSQQzWhxoF
Z/6nNtW/JuMMGWcmUI0iHCamkM+IIpjPCB3HBCz/NBT/LlDufZkmHz3ESP0Zw+tK
o5buOAEJ+SrZjdYdGWy1wtiROV3gXkGW4iE+G9ss4WyZiOlTW8cNU/hL0qCtWC1Z
9lBuzRP2j9ckbvZQS6b0EeW4bIPKAk75ZrCqa3JFRXN/nlUrkteRqE2Tf6WotO69
VBokXoCf9hdWfQFGtJVCCg==
`protect END_PROTECTED
