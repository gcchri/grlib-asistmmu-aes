`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YgID5ivmIeyTohHh507waiT+NhGXyzj7oeE+2GaCmQf/oPHk3Ii6GOubKNMO41be
JXn1lQG/Dqi6vdblmUaRnkrdVOqmmKRgku9seWZtjjQesqni7FzvR07VATUzzkfE
yvOGS7mhV6QWEL3ddnPkQrWGnNyf6nyCtZ0yKCbmQ5XE2kBqppZm1TExT8Gklvrd
rDP00c8Y01ZE29iCUtHq4P6mLH7Y5pVKFwzQI6I5DP2T5x8hKzDG5CayuMsKuuPe
Yu6ojnoNbqdM1O6hwnhhujxiWGDh3cEWOTxoT2czlI5N4hw5DGHLBsp6bi+MxvFC
SfZR7khmQidcO7/BGSccxVWuKA00CfOSLIxs85NbzQ2j5ePrt8tGEV0xWKJ6LlPZ
Qk2MiZXKU7XtugVyRYEiTaupJTvJBeY8lKKQvPk9rmtWPXkV4yxuZlwYHEhEM5Oh
IDD5AiAps6m1KvNpco0Kev3EAhpyGfnKr810cw4cB+WYQMEkb31CHqGOa9G6Sqp7
YMdn8sDNnHFk7wD/1m+yuq46ekp82g2kOq9eL9wO0/heuUHtZT2n8hfZhZSg1kOx
Vn5tS3NY+3QC5Dc7DZfKqWY5NyaVadUwf9tTSIt/N8dXkO/tQVDhSwv1yGtpvaU4
+lBmMt+YBBG/EZn0HuCEiE2kJfFtcPUX2sfzPJXljet0UX5CX09lGDf4iYQijj1c
vUxKGOiLjXdB1JKyxufLDyVC4RRJUAJkdaXOLrfZ+/iYfNxIuV8H1xL1hNHs+5uM
ZD+tnwsNuQNHq7J/wh2IES5BHsnxr5I5DbLFUOUaMoHp3q4HMZBwb7700Ao17xix
wVcq/aCVK9zG38CIu+9XzQ==
`protect END_PROTECTED
