`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZfGUH9/d0TsMnnzgezas7cHVWN1g5J45EespRr/WHHrlPtvas/aQfwviRj5xkrrs
VZORycYQZ2eb/5F6x6iGKztcT+ydgfrYcoKx/n5Cj1BC6AehMg/5J64Z+OloXuWB
mlW8LSMrWR03ucPfh4sGEnx5OUEgBGwBhPBY2BW6fqaTqTkFD/gYR9jvL47EX4Le
TzMwj4Mml91PCfnfvT5Z+POmjDvVUltrhkV8PV1IW12DH747lallo9kifPpaAiiT
DPI7IjPc8RjRLYxXH2ya4NP13Xq9gtp/FBAEPt6rnD5wMY/jS9oNmsAUMrnQ83OB
rcnyPQIK7V5a+4faj8gDasBhZiZiwtJs3EMvU2cbNE5qMLBqDT/r2HFg1f3nx1jk
fUZdn+G80WOtaNxR+SHQpKP8UzAbbCd2FkPRLlXPsA5/HWrF6wIIm669UgABgJXE
j8FHimnvq8+L72pTBCx9jjcEJwf/XPiMZbvMVTTLLNfGpYgpN7kpnKJZA4SS7pDf
`protect END_PROTECTED
