`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M8QthVolmrDYutt/8BTCAvhVuLSaSQ2+PFWe9RKTUTYYFxO0fWQytw93VqYedv6/
bDsOn/s29BNg6QWVfCN7enxly0kHZO3xhnvxmt+vWKYXR7jry8gBIHtEmOBbR5IR
/bIKrLZoSUjUViz7rBrQoagi2N13Py3ADMW/zsKwwYYS4bO0TwGfO7dROlqyAS06
SEZ5nmaFATpnwGBM07LTleDnU9GrmBZWKsEtK2Wx/WEfEfk0KCf+pVTSzMM+6+ns
o7SDHn9invqxwDr96byoYEhKFk4Fge1d+RbRWicXzUHRLnmaECWv54nBWfvbLtqT
Dc9BK7dbpNfNFQdN/hAiAK4KDJEvgTrVvM2OqH4Fs1raSA+D8MUMB5A1QdZTj8kN
NIxk2FjrZP06+IHzoXbm0pTxFdCeffrnuKFf0r3dZ2Awrf03maIZTNlk+52c17kr
WUTy8MwaZmW9Hw9eRf2l55kGx/2v/D6NtSFh0rrdD/Y=
`protect END_PROTECTED
