`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
flTQUqvhK4wXaz5tpDcK69Ct5tUd9lrMs/0/+L+pp8ze2Vy/XBaU10JvKzBghUb5
7vRsZSDQkjyZAUhJ+SvntXZ+NS0QPJZiSQcEaFTGHouVX6yTJnE8KCva1YIwxyW2
shw/LXtO3dFiXS9e6/MSqRDzATSbdMeCPwLQnLJj88g/e53wAww5JhFn6NloURcZ
0qjSzCv94ZTwtWIs6XaDydNlCwAH+t66MFIYlJCgqRhAZ/NlAXa+woU5uJr3fVVA
i94WF0MJ8UOf7a3hRyiAep7Fu+w88Ljoabpy7ei4Wy3E2rD52DEJiNw/pS3BkoKE
J85JRYevnRtyE4NNQeBqjRwfZnCAa8JYljB3iDjtvijedZIsuUs6mjgFE5Nelvkf
J3nqnlQEuvK/Tm5fgw6pbhZ9/ZmJc8J730HfAw1QmnGITBWFzFJmeCxfsy78siKm
q6XbxoghrfX9NXHI9ucI7Z6hO1LYSmW9F2he8bi0p0WItA5K6LgvA3A4W8YClzM3
Y3/OOU6ZEriuTt2ArhpDsdUn2vjsgZoTxs7cyUIt3/iH/bYpeZlkzLThQVjSE0AQ
TXqqw1o38O0fdi784Caxbe+ATT+QvW1VT1hmiPqxsAWEtymc5zfv1wi6Qi0Ou8qm
b5H6VfVqQ6GI3soBUvpbVIG53L6v4qb82N/kShNY5yeWolyv9xe8VqOiOU6Ve6Hc
pCnEXFiJWeoOvVtGDIc2naBJ9KdknJl3Ahg494ikKIRz4TxvLCG28gSrS4woxRQd
o+QP7bHDX/WGmWZrfZvgxxebkn0sZlsOG2/SmM5jwkDfjzaCicxBhmyBLQGMzZU+
lz28F8WM+c/E8yfYgKG5ul2larqbpsPmq1WO1UuCiDcAaL2bJJEBU7glOMnhqmnt
UHv2XDzj51aK1tAD9MLvEAx08O8v/HEjOhv2ERypplejJBU8TXtY8iH9VhheU5aq
BvTfz6vmYD498iasv04+wkcDNH6fMPVu1B3zHQz5aapH3E206TfHIz6eGrS4Q94i
OYJsH4fP4fpvAzbmfhaYEqwhMyyPIt9y9UiVyT+RnkBlDwUfYvd5+WPylu+MU8g4
SazxaPCPO10a/qpodFzoQb/QbGJwzQLTm3pTPAOR0uDum6Tg5QeiKI0gXCUbw9gS
vkx+n21ZHs61irOrRnw2zOyRehztJgKYRxYbkwJQ7qBAXdW9nSLbiBxa7VKaeXSn
PHh1pPTrTLIo5AD7o6+mPUWwkgzUvA/Tj31toE0GGtLrU60qcIsmp9iQ7sn964W9
dcrlNvoylA5LCU44Z2Rk5Tysq0rdPxDfUHzg0chYpqVtOUZb08lQD32RRY7IM5CX
1tN35zrTEHomxWN+lv/p9yL7mtH5Ahrqdtai0l+s94YRxZeLay1k9vWGrNUQqz7C
E3r+JtUDzETvgQ1BcpZqMhz+XK7UV54KWLMhDS2tYpzFPepKpXDfu70jdMoZ4wyI
ayLPH7ufm4/s/6xox/l8Hwp+BskRmrwEg4rI20f7M0agGS/nBAZHcxot+DXdszmK
6ACSTsml+O6Mf8iLIFsU1rfG9V1vaATDMDSGIomum6RYat8+ymE09Sr2MX/QSGMK
Wnrhf6YX4QCZF77v7EF4ayrwVNhLxMa3OZWnLoHz1WkVyEU3OO27Iax8PUrT4c0+
hX/72AOcPbHlW6+aJwzt4kVFFFv3UJa40A9sXY/Iwi61OMS3SOKEhzhAWHsOA1Oo
tGLu/z0mRksvBLYwVbpkmVRk/vwrp1gMZF66zfjTIVWqnXMcgYiD70VfOvvWNSVk
0uahYQE6ZJAE9t/nBpvEaUj5bMT+qKmzEXfTVRXYzPmL8yd042uDvcszOYeOcevM
ZVbdi+hiQJfOXSUmOHQ4ESSAu/Job82keHWKIekabnPqw+wENUFbq159mGOUPHaX
AeCmwywmjUsu7wZ0H5R4ZWGJlfO/TZ+yoAjRCT3Mo5K5Lmhtzy5jb2dRXlbkG1YX
CJ66bVD5AFGeL/I1TcYFTGLDtLpHJoVj8jiP0ggTmlF4FLzPJRiv5yLjDMJfxdlD
rcw04HBTihFGJPmssON3i4zbT0oviwKSQJEJ7Kgg//QxblHr9oqOkHiYd55/ev0u
Agq0sB2cgOmvcVInMusVv4gLQ3xwmPwRBvq4XZ+/BErM0Vur/DvWsCigeQNg6Wzr
XjbNHzmQOQQO4+sYv9AiTv0/lLeD29p+3ptlmb0bwTdFjyPQKsPxQD0joY5wrWyN
lK/7WfRsfHWkpI8Dpv85Jnm44I7cKouQg6Sdq8Pf1F40xt65oJjmKmTgc+RIvXbO
xKaml6Vas86J5abGQsSTigmqqy/NSPAeZbxejrcSDaz1bxePGWh07czXExR3whRr
DiVf/8wX47usm1PwH5egVjpmz8TX9YSTQa4qnhAGrk88sxmrdySbUREKfODfNZ2Z
uEv+IHkxSDUg64go5nwIyzfo/hbU9fYFyfMcoE9c85e7LcSS8lLdQitaRSLgKndD
oV4gveT5xWl72flcxeHJnGwqKEArjGsdhP9kfGaQ6OX59n8N9moal+o9wjByllQ4
ZuJpmc4tFnmCbTrezlZiXzsZj6voBB16WfRcjioODl+2Ow/kU72fXkAHIaUWsqWw
YtMKtF2mOadV4Laol5VhExPnE9dKg7NP24BZZ7nXc7iX5/eOXbVlz/yH7Y6JUHLu
gt/L45zav1bXSUGc+o2F7mVqGSRY8LbyLxakdrIguWlNNo2a+bRCs96WRWnJc5Ku
qeuJKDs2KJ5Wd0y+mhkYee68YZ0DpiYeHCleYMP2yEUwVBIVGj4loAR+ZChfLf3J
H7yMOYZOhzPRjVe8K02cH/fdniWY46JXt4QvALRqW5Tdu4LOBMaqj5wzWBTkKUQ6
J8aBNw9athOj9U2Dmc5hITlK59bx/j+bS1VXYzc93VUQr5ekz5pqYY440jljFu1X
So+XlBNsN8RjH9TJCnHNCVyQXD+rboYJVAbap6kTYvBj6NNTb0Nj7LnVzQem0GVa
Ik+8OfWimcO2V5pjTVBcJbQ/MjV7E02X0d6vduBalBgZQeHcrCSKh3aPDujqBzHN
lLtZe2+uel9UaCcXOdRoygKzlEAtjF/XwcJ3mIgZBwkflpOHbKjl3woxb9FHEsc9
gLsIzU000x4627dCc2mj3arC8o8bHJdFgmqvhzfklhZeh/djDeLKXyEnUI/tVjIX
+5+LXQgzNTyWELPSv24EEmT/mWy2MmpGEKpCzsY29/bBQXvA0bQJUEl7eogjBhOM
zasxPRaS9ZCCYqkER9zLnU8mMkE9UjUJobLIeGaeM+V4B//krmAfvahKlgmftX8q
bH/Xt/l2CnGXMHkxnldOMj5cshzMR4c2wGaFDMYWHMW157UnGRtdCyGToOunCcmo
L0gJyMw0BUfKhY4JHhHoEuKtfynJVm31rN27o7hjze4zJX1Kr+yOGT6R03rdMHq2
9OWs6GCuryNkwWJ3IPruTk/5LnS0SqA2AT2Ozbvi9EIm6qp1v/ZHZ11D+1PUIXA8
Qm8ZZaVL+lCpt0DYG+0+jxEdb5MYzkU8FqmlePOa8sEcwLZdEmzv84b1MbiGFpDi
OrgvIcQJ07daH6pqwqPYvAauwLkDqQwL8s0NljcUGYZENapGxMlFXtsxnOoeBpOj
2B2PUcXs2Mv+aQuXHHOG7hFQR0WXzOlaq0dpSi5XEWBVEp9CMJNgIdvZazoGhIGi
avLw6e0ZzsIFomAoUyZOJFaJ5toP3zh+a94qTt+ywhlTKqMbmyji9oeSDBuAV3Xq
VDRN27Xzw7WW/dK/CjSUr88mp3te+It/woZ5y1I2dpUDHr8zs3+UtdJ95KKKWu/+
tKOwvHpLORXIxGivO/rbNuc5UW3olvp2oV4pMlHlRqZJvV9iuR4iTIdo5ev0IpQ/
gdRnzKjf5HdS8svFtzgQlAu3Z05GxzFlETuJ+8nbVKs=
`protect END_PROTECTED
