`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2kiKneeQswGb6ul2FFn/u3ZkFWGEAVUoMlMEBMbTBxLzrRTyhfvAjUQBEOQW6Zj
IoXcNo3l1VAdeYmyN4mVNy/HytSR77lBvMA1yfGMioOQO9svXWBabe/6O2wApWbY
3qYVU/L7HNNpiuymhsU1vomd7kWZEZCnCIaDDelyNDLdD2LVOJBMLFzmdhjCXd/b
5nJjqY6bAPT71+N7AG7quethAWec65WzG25RPlQBbScd+Azr+TC1r+6upTKZDYzE
nbA4poFKQG4dnp+SX02vKvfPpCh119lScieVMg8Q4mYW4MZCF3S1WzYQn51cDOSF
kvplQltnX8Cylycei3U/NokepE4ycRzziMEOB6e5EtJPRagGEVvNPwFJb2IWGPKP
V7weIWymXD/PeHi1ikV2SKlMRtglWirFTFj+SnnxLlx/WE8q99tCDIo+9NHxOoFC
N6jVhtiHmeR+fU+pu/PMC9yJBp30+CDQVxd1qrOCcDatxs2zp41/NYwOUCs2EWt1
ARXh0copK8Z9chkkXSCCR7Zx9Spv6NrM7Kz/EHRkGnoELzOVk4YQJbX2yvlIcME2
HKpIdLXqG3mKq92/MHJZAzgrpevV0dvT2ql27c5iqHFSOB7AkjjipJ/5tl6lZEwc
ml3RhIrDpSozoUI2MEthWHwEM0qTV15SxQT/vNyGYpMkaqlJg3V64aMLBBgWpjqm
jkW5XIK6jn9vd5tdWfVZTHw1QOTZPdz7WvQmXN5ie+m6evbUwRm9QotFQpJUwvq0
dB1DuEov2Pl17wtGIfVicQ==
`protect END_PROTECTED
