`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EP7+Y8hRaX469chovvxYl/aoTFwmi13ysc+36AiJSeDllKnZloEl3OXg6PVp7nT4
NjiKQzd+0WbJTpEJxUHoBLsOdXrltoPzxxBtjqBgGS5HGaOsb3zd6/tlfUxr/XP4
XZeBRy/yJX4oL0w1Iz/mNoHmp+ktK3pvprEBpinLzl63IXmoogahWzMwEvhrV+Ly
oxYzP73YXN6K0n+qy0b2TLPfOwZyPLNEPdRqyVDnun6DbF9y92NqwekUDEERO7v5
iw6hriJQt7GarvD2lzye/pE6B2R57cU2lDshoGBNPIkuecaW1bFtbOKS6HshlDqe
H0Zn0PSiCZx4knTT9kjO7B72efvTCmPtciQmfZDhdq7Ymu96EV/AaW25TBwHH8m1
zK77m+5MQpG/dfL5OPALEGQxSDggOlhfl1EIOgO2q5/cEuGhWrrKcQfGt4Tioqqt
/atrqaycnqw1lIgGAgyYT6e9u5cDG14ATu4jVxhR/ULTvWF1yx7mU8f/+PU1tQX1
JbMBWzoVqW5Pgu/W+vp1E2BKhoZgRo03TdBVfTURiUbVBKwwMrwHSok8kIAJrh45
OBm8yK+QJZNLjUYvWz3juxJDxaQs7KI99FUE7jNW9VCmC80l5gZuagVoDAopBPtM
MGBkiKlx4HCU2/HSsoXqt7A2j10tZt//7vaWjV+2S8Hz5zv7iqe6tKwypA3Gptbq
R5bgfkvasRtPu5uN80XV2RIAI+3vLeY5dPU/Yn0oSnt0l9vdObgY333cdS/+MR+3
BvqynbzUM+tBLUfqxMPW6q88btl4uqTWGe0A05stgFC81mPZPgYMIKsd2aDnBYba
iZXDCQd0QBsB/ZDOLrANMC9JXmU2yvFNyplm8GD9M7MK4TbITNfvhmBWSG1X3NQO
nnB9qXqG2qlXQA28bauDhwr+wR6NsV+g//43hph194fukzWkVrXQx4dHK5jQEtnV
k0d5NvKWyrEXE3RN7RkRjzi89A+lQMI0+DLbyzC8KcY0wGfenTw2o1bFzOWAg3zq
uL1dqa9ruffJ976I8gNDlzHpCU/Mr0jLGF3PBDxawGu9oRrt7qdIqLBU2Amxe3QL
`protect END_PROTECTED
