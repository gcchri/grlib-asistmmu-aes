`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cwoRupO5+MXf9Y3eQsqMN3H3P3t4zm2ngIQQBHksG8E58CeclgujEApLFkyJcg9y
soqc/anpDSeieGZ901rC2CrfhdAw6PFFGloFgJG7sh87JCn/b4b/r9XLFnWhcpl/
W5yOEn6lUTcKXN4ctC/Xgr0tzx9raiksJhQFG2Z+TQn2/B37AAs2PGoeMSKV538C
zik1615jXb2aFRqGsr4x3IPOGOLnND59HIGiTAU5dtQqmnNR0kPBXhErZJctMwxi
XXBkwZ98Yf1hrX04/dTEnFKf6+VSxO4BcFd2XNdLn53pGGrwpIoB4MXgH2AU/xgK
lv33yNKG0xojbQUea1mrdGgbsX6by9YidSRD8VQDN8hDL/i1JsVjvhcJQiZc0Lk/
`protect END_PROTECTED
