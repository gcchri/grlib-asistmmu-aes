`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L9GqWqLTgDTLNC7MphaxjWXdrehJ0o9LPyEVKqAOjaml/o7+177lqLYmRbiGm38T
9J0v3a+QsECoSl3hZ6pNouyaE58SmBGwiTlXj52PVNLcryP449kr1f+h1ojHrE8K
jGk/bidPDZQ0AGvRd9o2sM7YgHoZk/C6xYWhSHfkHhnZEtGOfRmehrVR8HiS1kLQ
JvXFgn3/ezkhje4TPNkT0Gcpv94yzllA61G+dmMgQTYPIcJi3s11ajevFrQ3E94b
WldTqVaYjBm+WbceuM4kRD7LkmwvARqqpYir2qofibkc0M/4wfDsqm5A9kxFB1ZG
J4MAwOFwuous6ivWTbHG1btH2tDZ5uZb0cQXgc8gkubl3Wdet/Phdlp9HQIdgKlY
4nXbqxOII6dzjlYIUp2nSrQnlTP7qEhPD1Q8QPW3lYI=
`protect END_PROTECTED
