`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lJnoLObvpFRdUrpD4Y3YmpoTCSqwa67Xqm9AUobvz2d+LsWUDUoOF+PnQrZrRg6J
cBrDjktHT6mew0rBXqwSGig9g34/HViwFq7t3i843QRdvGvDRBZkDpNP9B/4Tuul
awjcGWfC1c2EKvJ+ssLdzflZVD+XDbKj/AjzDUwYtZ9X66evdM75leGvcnrMg2m/
HaP+BUMqH0j3wOh4Sg2/aU4+x3XrVPGQXIBf2ZfviEFpr5gVLQgosqZwW7OvgvJb
NB9eBpAP8fVGA3nEswpDl/5+h7mkbuIC7/XG8nhc0Rd3nL7sn3MpvsnFyZWHtvi+
8EUECFrmdIrnA8dBqP0ZsusiePsxKTitLbez6d8OAZq46lCwHuRWPBblV6uyN9Vz
1kni6ZIZY3hSZHLBiHAUWvTHpTGLeBI0K19E3mbftmV5oK92xFKFN/lL9IxIdU/c
bv2z4VEnnxELINTVcpTtop/jYpUfted8R6OwFnzEawE=
`protect END_PROTECTED
