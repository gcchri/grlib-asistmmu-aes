`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bAoHmytKcm1w1Yeaz0MroFfqB/biplFpI//yfsAgkVSIueuqeIrUpJYIXEvCXL1Y
U933K3sGr0y0WPtTgz/5uBH0NlNoq1UG/kiLIu9NUaVN1vVB5hxFPOuQhrD2tgJ7
CFK2TjSjYp60IBt32OgsXULYSNGOZVK1c6HMz9LWOe9nL4V3kbuZziQNDAUiOe+O
ygWxQxm24yehICSG4lgwZVEPX5g0p50A6No56OlpDqjKtKrNgIxyot9WfSpoXGEz
EPkwYwY0EI0BTa3tCGvCxdN1wbyE5reG1GnEhR23KY/7pQMWCouoT6+Ud2kSJ8X8
/QbmkUkbs0hypKcx9U2SAnkWVCCzWKb0yU2CMUmtV4QLIAY77XVECbLi99nsFo7U
Ootu/TvD27iKXd1HR4paEA==
`protect END_PROTECTED
