`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pBqWqewkCnXQ0SFk2wC6Mon/X5f0vH5hthHi7sulk7PzwoCsrp21CnbRzN2UPqT
XSiNHVKtUzE9GQCQwig76wJlquFtVaPo95136ALAaujHVU1IaXs2uB6k7z8gsxfa
Juf+M70NNgVPwr+DI8mE+tHJUImsNZbPD5IIwQZ3UFGDxObJ8vh+od99oJwIjyYr
2JVcayeOTlb34AkyMxYAVoVysFwDJGeQTmTRlbz6VB+TI7m6OOUZ1aG1YcfyZwJr
q7b/np9Grw+MubPS43SoEoGFZSQ1F5SOithdZkd60fjK22UefU7TCmuA+w0OP59q
ChhNYt7ptREH3CLXjGjaAxgHEplWPCrGmNT2/EHR+gXHYSIvAanJp7M2DdndZ2lG
XdvcHS+KtuErTi+BjTZrGi//vCJD5ZT9I6K030Vc5wkCUXWkmNfPoDW7rnk+WRIz
IeqXLidkWwSwO0jWGpzXlPbepOgBk9NukYcjf9zDuJg=
`protect END_PROTECTED
