`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMQ4MqqLsA1N2MMR0sUUAzlypPZmSHlj9Amy1PSqyTRSdjKLfiTZUPItK6/V3+8u
EvUuLlotDYZvhVkKnwZPk2nGkOUlJr3rodgpTQABMP4g1Qk6TEa5NwaoAzuh9XAN
dDVnot3Uy/9rcvnXVDHsk+GmIN7K252rshwtZukhsLccNRu+RM/S5/dYbxD4Cwwg
3N1b2F4ZExvYgL1CB8cGvNEk4q7BAR7k/CavzKTJV5MZzJu9RiEk1xYgabQKA9SQ
T3NkVliAgxmm3cOUdwXrmX7o3gKSLY29VMqnS+lzSRE6TqqS6qFS8SxA4/XzFfX/
tvgGQWsjs6fB9EcKIBNL1cbzoxlq7p8uovcOEXRuMt2xxxBdKaWhNXlpKKQRD7JP
EpnT7pS8MQeIK7ikzz91RYN+Mege4rGWXanBfri4WCLfE1aViSjYPetED2DiLVmU
9/juNiMXhJby/aH8qYa2WMWSetAUvSjRaJEnzOpHaC9qpKiIF7dU2Yvp17Rddgv6
9ITd4KzRRD1sCqYhOarEcfwGNZyUzvOTnLg7CN/TlbJdkZuG1cmPZhmFQVKawpj/
GQg0YpjfWN0jfosxZdXXCg==
`protect END_PROTECTED
