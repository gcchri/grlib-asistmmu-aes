`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2MXmB02Vw9bT2jx8ZvCBpqBc15rO1uHpVsoTA+KNUNEzqh9oLtzEnxB6umXS4IA
lSkOyCssLNfu9U9CSfn3s66BYk8oJPiiAKtHwSFZVurWmbfDJ56lcnkVMGNBviLB
VKRGke+c+JmmAhkCjOJyzgRkZUncmhjxG1aGi6N2O1ZH2ITDf/X6DfNODb9m9BxE
sem9IOZDIXRalZO+JetmDhsVB/bn9bXVc4pXYNL6a39wqYnsQ+vv/tralsJq0hY4
Exg7o3vHVqfL/mmIBIBKnro85DopbZVEGFMPmf7YWrJ1ue9JdnKIphgS27mD5RIU
IwJ9CoTF3d3xSsMIzuDcZvLZg/U2G6OG0+M8N5Pj1RBBHvNt1Y7bm4oSn2R2O2aS
RgkoyfW/xdrFA3FdXAW8dsO5JfImTwfvuEa3DXt1xgGVxIUWdEI0ZH5A28RLzR1H
cpxksM7gtCXpCjSQfAw2YhkzwDk9r+xOFLZFrFm4SWX4gPp59s6YgwJEQBvrlxEi
RYZVWDKyejM37cEUOsQ4o9dVLwipZ/au8rt04Lo6BthGFxQ/SYu7BUG1j9pUW+Cz
MIyJWEYoLlOKw6CbfCLiVBEpvHvWjj7cZwP5zsvur0vgHtE8cNhkaKnAWX3xkIl6
EhGUYi5IIk3uidJMBddvwcOlBdUFYJorOig/pRAb8zlB14C/7mvWm99jwVm6eVzP
nTMsUIR2/78Uuw9BE9t3txlSL/OEDMWyNwCo/wVx8zkWPgMVWKz42wT4gG96aO04
E6byaXEWRpNNaOZvfqyLjZ5kY8M1G4MAMAf2iu7Bvhn/hACDtPJoPhJhC6TFdQcC
vU02kllau9JZsReEm7MoaRXi4tSQeahNoPGQ+PDZZYAkTHUoHkMJ12F3XK5gahZX
QFBxVm1yCIa+hE1g93Fm5RJtWXnc8eXSphphW5muHhFwaCCFPFMR7XjkFCjZ0CHo
V2r0HQzngvr+LHmy4nhhInLNjS9ZVsCIMVWjrEQ9Yn8GBV656zkOsZEVgQRldEZj
uYaBK9p2tl41O3YFDfZfkD4FjY4aXASV97m0794VejUex0b8Nue9tiSR5muDi0FI
T+SDToculMlGRhbkrY4RfV88oNCWn3Ngw7ddqWYXrlR6yoCWHt3zAtwdzSpBSPWI
mbDpyH1Q3pbkckTLbY1FNfJmq/vJ0Pfzmtn0UY8cfEmhmmdkptv03NlUJQC133KY
Fva9KUTeAvjf3Foy71WkkmRtzJWN+Zd8d14F28fudlWHbxjcRYHF9yY4rLm/VVr3
aDR76Jehr4MiD+W+6lrTkpdi7/n/K66iLkIl9N7mFSGWRnfKlBnNo/xfEe2abAIA
xi0XlNHqy5UIztCvp+FC3WlC8vc/X1EeBrcCNf72KVoBghWdMzMopddY5S0IVxHP
Cy6FCUoDx8v8Of3UWIMz3cH6mDxTuTcs4a4SNrjqKM1R8fdBqMt0tIZPXiIGWdYX
C670xtqF5sVUaa4iYRY+nV8XrPDL/JiV7TCvwVNnb12ssax308A3RnWiq8IL2c77
pRCtqzlR0iCauQkvWrZvsVoBDQivNBO6viAqBLcNIiYNPrFr4+L8LPr1OQpbntCa
PMIKDyRuE3o5FmdmDCDfxWehfiMY9QdB5/gjWFpJGI5d3dVbSHKvl27rdnbMENPS
ySSVO+KtTeYTLQ0um0jifKcjM+bjUDAMGIq/uF0sFj51I2Pfoi/Ph3BnaDl+fzD+
voFgzDcH2Sg0QmFcKrIs4BwRzTyBXEjh6Ulw3VNhJAEydZE36oomfuS3dPLbseDp
hUiqPXxTQUt3zqiwTsK7Q0sIyJ2Aju1djWOW+YIcepj3mK0bkUQ0btNyMXiL7WJp
a/Ncke1+ELdhfl3XYgDcXuIbGvJSb3Mvi+LwIsPN2tbOxkHYaJjjSpTQzli2Bc0U
jrnv2FKfUiFqqCh8xEiX5b55sXxjee52OEsPm3+yoVLq0ZRTWs4kAe9LvucmItyn
HkReHy5FjZ/q1KdTXcMMIOadtT1SxFu2+WlUCUuH4FmnIgolQqf7ETR7pnC2O9Gr
OKNwFIFaCjgLV5sLs3EW9c6hucG7bWX3P+oB5h68s6o=
`protect END_PROTECTED
