`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QpHnBJUk0OnCg7V1BwrdTYxjRv8KkXJNxp6xd85hUEFRsj5TXg1rrXFs8eslf+Cq
U1wDNIXoM9o9tDJQTC6LjYJPkcAV5XmGeikmmJ1IfW/RHsFopqEluffmu9N67uHE
bTUoCTjPyKt75zkspkSNRTO6sqNhotpbUdP3sI8IdclNMGvPPAB7uDtPSGVuSWek
sUUZ/CELzEOnXHz67CTdEmnK1F1eW6SdCiypbdN5twtsrl2nZ/J6ExGO9e5BjDuW
JdYjf2Y04D49y5KJKnpUCEVWKCQz91KB5q5cRNsZuRPldXhk7VJlphGM4Y4ve4IX
oQcjaBWF99bku9wlrbeLCayQspmkB/7ch4tQRWiieyh0zS5Ebc5ZViQekKnNQjpE
H5/+C/8CsAqdib4sDs31eikuxIUpkzixvy0abRi6555O+OwJhzXMm3LXno5nwQux
j154XF2Gd1wp2jd3upRcHnXPeieXV3zXOCGgg2045mx/WE5bCzSHdTa3RJqh+C3m
p1soLA6MFVwNsOxfBjeHh0fpSAOtDpGw3QJDpVV9No02MaWc0Bh7Fh+Su1l2FjOC
qsr4arqFuyTKbtl/EWb+ZqhkaTodJ0jeBQA5QcVP2jYyltWFtpec9h4qxh+EBGXb
eFoT9Z9N1+yKOxbMTScRYm0uCsYAPCKNTx9X9i7tu0BjYyzKVeHCFf/SsGafTGEo
KeoHxnASlVX9jniBbt8U5PQO6Ui+wTFLaO9qk//mTnEsugkjci7C6ejVU1g78+Gf
QAua87ZJLkHTRfVVExscjIh6HLUb0yHUN25gZu3+b8Me1xsaj3ZGEM4zIEyrd95b
tp+1ytGhBYxcuU0+R8BDQd5wLhCr+h/tc+H9ycd+tW36zA3pmt4c/b4TqIO2+7ms
7qgMfR4IPOuIz4XdXpGo4dqKBTzbI5ofWtUjQ9VG1+Wm29ihLuXhxQEhh7X5imSz
41JjrUlsJE6BdEWaP/FRSzuaJp+QDOQWGo0SEgfnujzcNyiME19rusWabwIWH6im
KRtiAfb3v4GSj/+V94PN5xiwirkbB6b8ApLrGKtJSEk720aSQfRpdrpEol2pLuD9
ccAAEJD5lngkHOfRT2GO1E1zn6yYHjW7rpdIgICzom1AXPn+bzut3qSHhwWnjmhY
iPcBZDd7a+y8odD8sthbFCPJNp9g/MBpEHmnDWk3PB6wup8wV9pRRfLNY+oCTnrK
l7pzmL/1PfD8xTj5Z/bitQ3Wm9BraWGTBkVvbNxWaFv86bHsrgdhQFo2ObrOkDjH
PxfOiYd9I19Rnab7jRqxNYLpL79v0MjNe7Ei23Yf+pCmKAfO5DZxTSgRXIzCJvRO
1t1JYAPI1bB/iAOaFzZ+Tpy83D/8C1b3pSQ7ss+DyDLFGxDFPw456Yu6uVmM48Qb
Sil0Ijfj2lvEpOJoa9LUy/F4C24YnxhweIRThP2D6mkXL3aep6siR+8jgFScIW3g
B6k9bgXdQZfzy/SiJSFA7wG9e/CEh9Uqxh0E8i2uHJO4dv8wOilZlbd3YnlaJJn9
y5BfzFCviUO1M06M6jQxp8jd+IWaj7gU8b4bT0jnR+dZ73uF7rzRMAF+xrBBbI+l
NTmYQ5Lu+01bPQ3kEtTNu3KTgHb/kXfTBdosgfDWVe+2s9QRfYQXnxYEfTxaONz7
TFyYAO1M0kLQFb+Jz9vN0n4wWdpo//L2zQC4wl5fQbbr6OD/PernMvjNZmJ2Co6b
+r036hV2wfRTHJk0MDb84W8APOagMtHM7T6GW81tLfSaIG/DnmqTmsTH16I7nVHr
L0JHGjjrRNr1znkK/bxAtjHlaZ36AN8mf/gLlcfLw8CTDcj6S39fGb0A/FkllZvj
eorTKfYWZ/jICRExVafCIX2eFCTvvW9owtfB+/3MSRgwhxTItlD7MW5VrtQcQeaP
3706i4v4PDv+/bvWU/Z0AZRkTU72WLWN0x8oea+TbcfCwOq0fbgOopp2FmXHL9Cj
0d6i8KXpIfotNt7AwCsKiD3SMi6U0jc8rgpCQzfVxStON9NAz4L3JxFGayxgTI7p
rUKHA/JApEU65OG9ZVJ6+uIc1RwXmaL1C02jXR819oMZApW60kAnzfkeKjPmiuVC
ZxEBuT541ZrJm8NOApIaNKrWiPhx4r8ahWq1CtPG7q1iZjOy59+xVSv6Ckkrudl1
Iyb/42jX4w4N08fWnDyTJXIIpQEkxdI2bVAQZsFMxCNsz2XP5sNL/6jLMomj03h4
/LSRhbETkf8CP1n1oAB3uqowXhNSCGp72WRrXyhQhjoapIg2RKQarR/aHx9ms4EG
zrJTkqtKbCTTJrBHTcLh2jn3Oo34IQTzLqCPuMwQ7JtcUD4Zei9OpwuU1P0u5mOl
i2NIKHu9m1Fd3jXizqbA6Y0tV5+XmsaOlI7Br/S96UzDSznZMrrREprEmv63+aio
xWcO6Pq3+iTgHWnpwDoYPUtfsId4cFBXJ4M8TzNUO+6pmtvQ0Gd1BbFakLDVjWk3
D/Y/2AGN7Xn505bkS8Tb1lMbnqBqiQCg27f9e5wd8RyQeSkVCunDnW56LVm0Uo8m
BwXu/Knb9jYeaPklWuf7TTtx4nS+UdeqhNK57iYD7s125Col5N1RaZ4wPRjwDxLD
JX1DoFmb3LkZHCg78Vd0ErHrrOQsnjH2L/aY5PxsYQ7NHefbYL7cWD9x2TkeWqz8
zTnP002ljtq9tW1qH0bGDCceo0A+0TEUlXLWccA5NPb2OaoCh0osBw/raODg54dC
XnK5CJSyvrnVhdCTXDBcHjFHfVWiHT4FVqKFkGE3jTiO92/BH1fLHgUpqHnQiKbD
5GMJK23MFvnVzBsN4CQeSVIApJWdJcqYcGu8gyqdMbaEJCLLQYgcdGICwgdeWRtu
NmKTfLD5I10wK/MI/3UzicMzDX7Ez26yIySEB0ByMTfa8o78h+k5K3iJSP1SSI9o
K7PKnhOANv4WPlXZkt62nfCMg5EpHCdOm4cgBmrWH1ktdgHh8QeAOoYQ564smHqC
o3JzpU5mt3TbhpxnFWNlEvVcUWXTjoCZn8gJGrgGGBP+dJQMtN9zXhknxGDxZsla
AyZIUHRHnuMpkqtUN6+LDnKUmtHOf/bX+i9MiAd98oxjL396SIkmmJ6uRJolNKQH
tv3nLC2inoSh55EJiWyUvwArifpgqJ1kwm0rEEY95FpBp6nphCEz56jf0lBoA8Id
sK8VExkM2hLuIzisy/KJhQ6ICjEqoV1X61TuvvsxcOuyYvofvu50LHi+nZP54scp
exA4mUd1txJ/+7b6phePokwhWdMGVaJhgjuSjjG69589ky1MPuRbIyLRAczCyrw9
S21Jcsk8KJHsxP3W1HEKvfQTkaYfuES46dxkzxBeqXLA2P43HxtIpavr6z4NmA4j
TYxy40lXSvec9qfWwdv6/MGOr9zWWW1eykR7S35w5x3vzYkhj5aIs3E5VXuDlQVn
il3N7yaWVda2miECPKz2Ftydz+NZ2QfTYM5F+a2aj7Pp+l8ZFmcp+RTCOstY2+gQ
CO1EPSnK9N1qk+Q4QLutpIDQP5Eolqyxn+cjW6WUyA1SLDEFSn7xPOcBep1APdAI
/LHgBG/Qwa8s2kWw/YbeBGXP1vqVYNmtSSfFXjrxiQCRv1zF0z4B5xOqwxXQqnop
GheocTlzQ6cqwOLU/f3i5rqQ71u6p+16OEVZeuCKTh0oalH8p1ONBI9e38bR739L
Kf6llGlCoyHP54mzuwUfSJ/8a/lwuAJNUl4gKDV1H2jNBAlYt+sfypja1k1kGexM
+yytN3/qclBcMZALZtxRNAwnagiPunUJs2zuxfjc4gRUTDqqvyxKGLMaZJpttPQy
uOhyfOhNXkzID7nyZTaduD3D4fCoD98F+PvDJBwbarNdRZ+sk8qieuBwIWGY7PXi
ROvAqRyGVlM5/EgtlkcKHDSqVz7EBFe5jdw/uZySx1K+9+cM2tE8V54RPvZYfRFh
So0EH9WRanHFYPb+yqoOkXGNgR6jPs6ufNhm4U+m5sJtUB1XdUuOKxObqHNi+AqZ
TUNYDLU9gWxEGjVzJEhNDFVQFBMOWuzqgHFDafzgimZhkv/EWnaOpA8qzS6nIwK3
HkyPg8lL+qTpHyESpankMtd3igobXQd/IIdLkEo2Vr7Z299rLekwKfJmibXzY4zv
yCfsHtK6xrAc7ZIeo33ZEyFMAG6LWSbUEt1jmxr2DVU52QNka84EhKMRZTL0683L
CAgVXz+G+AUicF+N0RzmM2lf0rfslZbc/i4fTrpwW+aC2gu34lF+JU7NF4urAyTR
8cjWppVLyV6+OCxPYOa1Usgi8Mhg83cRazXYG/jTnlIj/jKllCYTTFhF2aS6sCDN
/lEyTEnQHPXBgRYE0A1TxzIa3MVRyzeJQzDLazhI7j6nSqRpT4XwK4/BMhFP26vz
UKjvxv7CS/pCn+QGcQ7XMz5FnKMpQvTmj4z4VBqaq1/gqW7N3ttQ9XP1WpxN/BKD
NA3LMBJy+zljSQccxhvuS+6hSAP/lK9D3zIYwa8OTOngPzCE1EWTJ4AvzmD2korN
0jo0LSGJLN7uP/9YbAm2G6NYcKzqSh/CR3KNAtsKnDwVxbfWw2MsmukXGT/Vk5HW
G7sssPJKQmW67aqSfr1nfO8/RZlAqvtAiP0MZw/tGBsoCr+GECRHjXX7b7mmXoo8
07CH84Mi/JbO8VBwAM6oD2q+Yx5VUywGCXILYsaGrgzRbVs4efPRZC73vpACS511
766P3SNH2ZF5HBFMwfGu+vyaGs61hasiCL8a4D2IWx1zI6+l/1V2+50v+w5l00+J
BkcySYQvLtFMpP86r82JzKNGXkGSzEPyvJWIlfhpQWoaW+Z62phKUT3OSZsPHLjZ
rAWSyZLFaQzhRFpY2eOcKaNDB+fwOzbRBdHF7ABamyDPvHsASnzRgLOrMK3iXUn2
wOt1wBjpLtj4nEcsN1IC3AGKVvMBobM/ZNnzg1gdQ8XqxPVDP8Q4N26sJnqE/iX5
oApdx7oIov+JkOKGfgJK9Wv4FXgUXZiNC/YKO14hESO840Zd+CkBpx4YzD08+LHc
x0OUjXLd4a6yxS0UNpM8Lc4PoXLVpcOKDazCX9cjrWNDFaeX4/FFysE8v/8CaxD1
X40h3foPq9+csTOh/nmTarLbIGeXjgpxRnM0Trn0bFBITd/hOc5AAJ3fjqTSTqF5
7Ouy8UMmtjFWfzwcRHDni84qF/4NuncH8cEH/olUD2M5ohFN6MqZKdPkOUt5gJ0L
eB90HFbWcoXX2ZvcPoEgQ5TR4MScl4jr8Yb7C8ySgbadzXaQHE9wFKNhYNNp4MHk
zltyJ7B2l/buG4/rdO2QV+/jN0BhjIY7EP2/bRTJtzTXIAiVjHUNnITBCmOpGHe0
TdZZoUbuF1QTeDAdVLmGQTfKQN0dbe3C6k6dTYMj4yGfkb3qQdO9VR3i2ZCOMQ+m
x0wVvdyfPAnyMk6I4RQ6pj0ZNu7PCbYjDa/TAD4kdJJYpAqtdxE8wgQ3j390GgEd
ATGAdxWR4wD2c3V4RlkSlvGLijoMmDc8vMDmk2woec4t9NJRmsESW9jaC+I3JQ9W
anuD3kEjlQg7LPxssWx33aNSrEMs1y3Q5DVw0lmMyXftbNImsPxAe8ZYD/lavsyW
CbGD+6f3Es6ydLIrAeSuEmJPUcqI9/VwM8Gv8M6zJo6lkmF2pUQISNIo1jjJ3uXg
/Ew9uIbUQIieA/KEzaQMIwMxzhQ+Hdk2UPGhcp8dBx1a6QmNPU2B70b0WGm0G1we
0oQOBk3CDqVO7fjeLIJmymx2p93yEwYylVS75q7OGOdxncMIbUOsyyJpmnERILU9
m5YnqG0cwOeEOWpzjx/P77NkwfW6PppuZC376yqXSFPyqY9vuv+X3USIaYEdAYxh
rHGhylMxvCQKepJ+7WjyjGCG//VpHI0QNgw8BmZgNwfxn6Tkm289sLhaxA5JHXTh
qLF5QTgWsZkZKlkpQow86BoOweaKFce+5s6Suzbg6LZjYDPxKaf2g5gIe4wxhNQx
8jo+FCiv0JgPBjUwu930n7lvwISmQdctW4LNMoxgo0B9jlQWhCOfPcmP4TwQCPr1
o0bRYe+NKVQ2ktPbV3jqL+0DfXgd/IPiZv/1+B7u3gVPOScTAhoMN2UZdB7U3cgy
aD6P1g8WtJViroBZexos6FgRkJZmibqCuja/TeTPetYc1TXN4ISeBy9SzHuBhk90
T9j5xJcYRFewe39xgvJisX7/OzwZf7S2iRJktWz3VGWRzhjAI0SsRqVJVRNIWy81
cmpxegPEL8a8nx6SKMvkwJE+VuuwKpRNhuUjG1xECnlAPj2/Y90k9Amki9eRo6lm
DP2+x2RBSuHaX2BSkhn7WMZRlci9K3LhFcZQkF5LdbSQzq1y8Bo78ImLDjY+shbe
pFNrDgXKVjkqSzz7zpvShgodAGUDfqRHoCY+gIDVh8iFtxATO0MqAGuhf7ZHuu0T
CcVQ8MP0JBF/nazbEtrMCI8gLccjQEb6JP4jF3ymflXvF3l++OLKuDgVQLBv7nYY
ylEcPxc2AXbp3i5n9qVGiRAzUARrUQxa/I8TXSHwK3dmT7RUyNrO0VCgZH2tIBhU
BUbTHVismq862x7oo4KBat0t0KYtFc605O8erYMU/uWnXrE5lVqkGHV4+LXHysiN
CZ+YqjPNAjhkkYCKBcZqofxyYZr1EiSQmILY2aT3ZUJalo1kuak/SYLY6l7v9wuD
bziAeVhj/vVo3BKNvjAvXQvErr8d4KfPYzTuK+DOc7Qq5u4L/ihED1M2RID+cKif
L5Q6P252X7YoBsaus4cf3xBb+iIKMbVKX03SDD3ktXneGDFsKJFYr+cGoG52wdLA
yZIBpURzIohBV9d15Dnaf+QC//KswK7HmIZWRRr+pMhy8IPWhX71/v4fA5BYbmBs
KSiIUdthDlux1cAJcsVPOSrZwmcDXKOqckiJ85z/B2kfrgCkG9CRnQ6/bgp0A15j
ZCCSDGluwjYnwy5GDnYdQH/KgOPF1MBt/Y1rr8rkQo2cAfZ00sabEFT4X1GamdQ1
WeuXsWlX3qlxYevd/fQ20y3d3bRZoI5rhHwSrXBZmdqMYewS2QmUKOzvhcB5W+0z
d2oGeAL0APFIUWynl2aOS/TZMySdkzcJB9dr89Q2AUE+bpWH7QjzW35z/pOOpFgZ
0HafC5HtfJlCNjhfel96pHKndyKTl3/VJXo94u5boXBHjmYw3pcWjTUqJvSgaVNG
21kGJJO7HiBlU5hs1F93EhGVUB46x+an8XXzDjb8jme2ukl8pVUHRwoeRqqUj35U
/pgtRUn6tAdcDi5BxeeUFI32FEPeYSlYmUFpLiulzxMR1zK4EIo9tJLnkORGzRPt
4YQVDnQglOHjHcypeEnEfmVN3idpzKpRaJsbWa64jKU099I6FsNzp3VZjvpinMTM
/MTqMZrlmFCT3L38tmtzXjWA64ixg58TvRCUz+ulRje5bkqDJRD43Ym/lr9MU4eZ
m0gCrU49IgtcMp7HeVlbRgSNYuoOy5k8IMuoamK5WQM/fU+nTaMQ7IZcQ3H8vRy+
Uido+3IFUi1SxYYamhsQAqPU/tjGGexDYjVWbWyeVEpqItO/PsZyprKmWFHKvVTB
RqXBAh6rp9yTl4qRfEmEMsYPLCQmCYv8j9fEqUcSAtn5PsMD8me77xcOrP+5jqe9
4WHsx+s33iPeHzWPKdk9bhhcWkDL4yPcP6nxdyV7EAwHOGJ8rEY5kYFimwkP+wAD
3GHrtnKSjzsAQxhTx0UtQ346xt1k17r0XXA4nIfqzkeJD9nJBf2LCBHo4+VNSiEc
dVPLE7SgMqOYFWFAgXsarriCjLvrKNpdmsfZiIICUDU+8wPGJN1HQ7rLvDFhZdoZ
P18gkC8tKg1eAdetGlgwMKOZtYiPDOQsru/54kI13UdKHEXT2xbA4iQwzDkya6iy
MbR0p3WH8IyrAYO3h7oXOzJ5+14vVf+o1Qj3mQ4RfqpAme6vHn8RpRD+ThfJtxnV
sDc6zcd7dyUI0QQQqEuNZZpl/13UIivxJ0AytQqpL+AwhKBvqItuolx+d5+gcSgS
w1fg6ceUci8Mq3SKbR4iA5y9d5kNXpQBRPJ8AWSGZ74tzDJahBp8ZwXYhffvZTvk
nb1qphnmWKOiZPdJpVJLK7XLgSdaMr7yqs87uFQc2foseqpm/IcGD4PdVeEFajgy
QfPSgqdL4UrIxkcLNYpn1fUxaz9Bh+c7PPEnqBttUHQbKIMeA85ky8rdDp0uNDyd
bcM7nTy88BhvLXjZbZtVHb7VnRz0mi2xNAHhAi5hyIJDyBN8K91J4+KRX/4Q4wBU
Ij1pXt7cFZZDtGSgyNnN+ECnirn3u5Mty0N9MZDOGmFDI7sA33KaTF5CFM2tJ+zc
`protect END_PROTECTED
