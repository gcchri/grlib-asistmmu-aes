`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOWTTU3JDVT454W6dFMjqkn3cvB06u3s3K4rCAjsn3/8hp++GRTFRy91X0JCysOk
cNY07aon0EqyJTMVuDimbKMv4ePR/oPH7CaQD3ZskMjKA+JOhn9SRIBtmVuMDlzw
uzR0mJAfXwiEIM54Sz8zKWXCLF/fbw4oDhR4igx9NsTlfwYSIGfJOqOgYMrJeofz
G/Bf91AO33dlUorla1BXQZnEymswYICVQ/wUG8JGWjr29xWJcNQa8NLf0sAoSIY9
vVVdv2n9P7mpR0k8EpFVg2PCv4+RQl7VuUMvXfnEefg2J9mgAGVurfVqT5RUpaAt
GHdzrXnJqNJL65VnDWQzF9QbxjPE/YGl+wSeEBEMETHdGjaAmmnUosVUw+I+2VLs
lqpMowxTTiqBH5oZybXd/RQtC0PyV2ytDvrexO8fhHE87AZ+Gnzb0o10d+x1a3Oe
hHOa0Kg4gm21Sk8goYVyOr4Xgn4Kb1z+9xBS5JdEEAA=
`protect END_PROTECTED
