`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SfPJCxLBu5ds6/pGf8atRg/lCPV1RP9n6RioBIJ8W8OX+Pk1zdq42yoUAIHAZNSS
Y7QR0fRDT1+bEvqmxrXsuvpxL3ZND2fRqmVtQe/ybKPCJH+OEKzRXkpsPPNRxbgl
DyS0P8JZo3+7MXsV+QUgMvPgudyl2kfvFku4jlMSCrAkhB0i18TymZMPqHhEVluR
zTAakCJFTqdQw+tTzDazoWLGq4wYZaWBX7GrfVnEMIphsuVP/CPF/PxcGX4kurMy
WrCAHfIUFy8xvi5lv28EQ/RZeKCSNLxWVusxEE7epPQ=
`protect END_PROTECTED
