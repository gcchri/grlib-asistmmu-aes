`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IkU04qeeNuZ8rNXgjDbZ8KphTvpPtTsHg78l256KXT+2jbPkQPf6r0FIimQjiPuP
0Sv/ybiRb78fk2ECEa353gTCNMYmIXqcOGp2o8oH3Tdk77/ieojP4MFJdQixo0FZ
qVEV9PaDFo8cTWKMqbH/+ISSLx3KaRBN7Hu93CpLoNL7toug9k3yzZU6JUIixd8w
2PuvrT6//em4taHQEGv3eRy1T+ANkNYla6XPcVAkCiTZ6BtSa0aVk4cUOu8S0MBW
zrtUd5+/whNbQ+YzeT4E1/NuYjZagv/vTx5C2QpTNlJt2Li0BXI4DzLMqz4INp/4
a5hbWzU0PWjipG+iYDUU6lPHVg6YLmOTNcDkHbrfMz+VWadVO126vvF8Q1Wgxbvt
ZMqTlLT65lFb1swd1etKiYcUVdG4PQzm4xwhLfyAA0nMdGb7esehTeJZIyULEdUL
FsDv+JMkCkPwXNUBwG1wvzDlEjQRYLmmehsRBCJn1lqHfMkhOLtGSl0WY858r7hS
0id68IP5Q60zrxFt/kY1jiMoYE7HTnCcYHay6oFJ6+fc2yOm4ztjo4iN+5OF3SQP
`protect END_PROTECTED
