`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VMtlffZyGo4PTkuyWDqNiuGQF9H7qYGKM7txKOqAGJx/LihYCw7z7hXZjfVTMDJj
va4WZtI57DvUoGnUSBuTfrsl1IKbR6tATEczUDcDVZNY+wVUXPoKZaY05f5U+Z9O
4JCmZT/o+E9FvPenxV8CA3nAczQwTIW3qItYFIHf3k6e1WDDzgFeJfxjfjsvB3VG
So8hkFClaNoLUGXi/fv0S8JqBvBqUAjL6McSWcnjILktdlT0bmbUUHkm8J+J8T29
qDE1icK4JMkIlEavEk+Mld/OdkAtvHajZ7RDEDwAI3yivL94DF0AEpli0RnRlZnJ
rz4GxmV1UZAcsl5uIJSwAyLdth+ne2s1StVN1R6Vvp4WqK5n44ZxGphIePN3wrA7
SpDJn2T0GyGCEhVFpBrO8ZH3xQnADqgl08sr/EAUS4nJmeydOehalM4FAninC+NK
SbYamAqBaWDTdGUr8AaJZn9GUwOO4qoOwwzEeOb/BbUkXzyNq3av4hEhQ/rduaLH
JHjGHq9d/0cBNxJg0vJ9SdAgUkTeSAn+QPEITHnxr4CX+m+fpIl6OXWEqU8l6VM3
CTItTbwC1GcGknsRZBrj+0C+sPkO/crx9A8Urjp8lkKAWNUtjSITqUHQLaN96SgY
RgVld+LTCiIxUubxx56sa2e73YSYmY3Su62yaHP3sAzVkftJDjtLMN4i0FaoQKVE
O28XYZ/VX2CIv4bIOTAEAXkUZ+UCchrn39JbZKQRuTdVjy3KByVz1CPgw90Jro/R
y5VXJCePYTxXD5d+PLwuMF5+R1BsZE7k9hYX0YL6jN8=
`protect END_PROTECTED
