`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPipNHD2NmoSkS3B9ih/tMRiH9+wtQdK2EFBCGyNlH++2o//RLb3CnJqzoyyBixk
qHibYsyAGGmedkWmPMFkCXG16IaB1THnYzU/QFP5VxKwERbJw/sxU3OEV/8Xy5nT
1xlkDEBm85/KxkmC9ZobdcrXeh58gHDdPS9nnrIRVmmbS2rLsy/VO/hMwvxO+/WL
ZLFlaJwOYQo42fVb/E2aAh8oVuVIJ/yIvqgHhw0sjyXzm2POg6HBBZKF9uhYtJEe
P/NYl5Ggf4Pry65TOg6GcRHMj7aop1A/QK1GIsw5sYwJN+zYbN4MY1TkCVdONEOH
+/PndeUsQjBymd/w6tjGSpk6XyjmyDqUWw/qkRYub/LbwCtUWpffZkMPx3CcPiVG
bVnBG5Ae411gKrxD3jxI0WOGU4TVtHRY8A1d38wIBhwnrOXzSg4aPnQV9TnHh/9d
lw0SHQej8+1bHsMoArSAz1bbcCN9EsPOAW+8aH2lPGMug7RTwpQ7d97wIQLU4Crk
ZEgqsQM7jG28LPSpQ3zX5itzKPrI0o+4iEJyLX+15C44EBlZ+V0/EXBXGMPnoa/1
0khZ4wEPIk4vCJkksuaUe+8CttNWVkMwBlXfI1kE4HZ8kYHI3FZiSeUpgpkDYjC9
fOQlZdrhDE8OS3xpBmoRnhrrsLYa4+Hy+OgIQfEF03kuBgK4q/KNOkFo7QZ7I2aF
xAxaYrPZTQrqk4lMvAc6Sd6XhhFxr73umX2Pb4x1lx4M/rELlWMWWqu/6nRmyZ3m
iL4IPKdLhO3xDxi6gwczvpIWXnzZw1Crp+yIVa9Q9V0oLlRndTmajsu3kOK3nBYg
kb44qaF2kgHRXs/7h9kypIvlbLRCpQaeauqYAkRWPQGfF44Ri1gU51/R+bOPMCvV
SRw4A2WhEsZosD/D6zH+uMJRscCd2N7/yzlAMkZxFvQycF3LSbiUknKRc/CXAz8v
9uP9EMXOg+q12D0ux662Vey8XkD46bljJVKbEVFoFUO9wdSF6uWTaJqzdRA8wuA0
Kc8Z12PY++R1GjCqrAbwbUACPXfnkIk2I8fD+vHn7vLKzFdnNBUIGtOmHqeW6BPY
VoWe/LJC6Upl37jmM1vRAZ7mz+QSGZjLVwXWtSvsQu1bo0jROwMgFBAJ/9faLSGa
CEShvFarWnxw3MayQtw1ITtJGRhWyWAWYiKyV3RyMlczr0P/QORIGZH7eqBSmYrW
Zg2VacR8MrtZbgL0IClGvORDh/tjM38g1PZxoaGxQJntIHWr2oXeVBSVM5OKTTE/
QnxW5Dyaw4Zb00KSQtTDWlJuHIPdD0N4hWc31o/K+mnUBVUZDeNh9Ev3TeKgpDPV
B05m7dEKh54EcDobMvIBUrHj+OtjxI+uBVJ8axKdhtOz4CRuGh+ZJ7HLk9Djmj/s
vWrK/PJ1pTnHpuwxN5R5uScBZm2dK0PFtVC83r56I7AbauBs8PqYvuiLpYtUTb9i
LZjr0Ggb9UW07RQMVpKkuQvwCCND1bPcwBKdRI8eVpIT4AOtEHW9IZY76cpPS6mm
OZn/XNBaiLify5UyaoYWNFuMRkWCiS7AWT4f7wRf2SMklmdYLmvDD1Cdw8TRHQt8
EFGQye0E/MLMAaDxBOAuwqiA1Vty1DWrODn/iNX8S+6dZ/i5l/EnApeIz9eQNsCY
CzRamrbB46wY+jAV545C9MzH63GXwzxA7gQmUodcsV4/MINF4GHm6mqwNFZ+kPhq
ZmsGkT8HhRvrDjClO64Jvoykv25BGRu0uxqAKP5e+BhmOBJtCGuulVJH7/7CjGfE
URAOSUovbWLCQV6lhw6ARTnZd7jLzIv/T5p0SSa2vlMrNvlPJR2QnUtWN458R4wY
5L3fvx0cuH/HQrGbqfLKVDeKe8nr/dpDbhZ8QZP7KoxEDK6+gfvKh1E9MDSs7A65
0+T3HmfU5F0XXlkDqv8nKQgZDC5OJ5vrL+dRmgS6TSAjoXf6GD7Adt/Lzpc868TE
RboiD84JYE1QuoVMSEYQ19BbS60rx1AYGjN3WmBomv7S0cO9IIUgNuFEI6atvb84
6+WFCOr1qioHKPkeF8GIodd8CybIu0+Ajw5pCKWiuGGaA7+QRSml4HXpgXWDRHYJ
AUQ8hy+Rb+UjXw+kqt/lT3bu94EcJkbTlF5axOz7pO8aqwiY/qin3Vl92LvpeRlm
0HSCUkK6GxmVHfKQvhO140TUnPHCSo5FRAonACbO8R+AHTBYETD/XRfkjBmPrGcS
iuxrrpVUaDKn33lUzfrzvypD4OBt9eeJBFMrenmVPMOMtzhDSB8QJMNGpBmkt+BF
MZ2fPthYQYVddvQ83fLzPs1R6rmOFqiqwQ0558a8FghC1vBGkSLeHXAXwPTzGKRN
cTwlz4x90ATDxiyN0T05/PIQOv1+N8RtSXbncY9YDp9ciLBS2n7Rs6KCv5PmyO0k
IWmZuUPYuRiLRVBep3IG3A11ZbTrg+EfDBGfQQa6rN7TE8U8vU49Ri6GDsSCLivc
GFOoB4I0Jx6bvAVO8TTqRgUXgOvZI9Cz6VmHAgnAFpCljpjPhb+VmyxEU93erA+r
b6h0n6xOS97h8BgNu81Tbtj4WcQY0zkt6slNnKyxXx4eZEk0mX9nStnNlr612Y8K
dO6rRfPvCo5Pi0nYPxH/BDS3KgUtpzL3nIiJ8ZRu3G2IZtl6mKVPRRQp5IFGGUoY
cbPK7gsqjmwy8LYQUUN5A+YM2cphj7IBP2YmrI0G0chzLB89t+oKjGVsIH9WhCEy
9YdHaXVZWzyn/h9P088KnAzRDywDItU5pZWgUeukaRXlDktayVzNVfLLlF4XOZg7
d8IWqwD4kzg2tChN/uR29biaimAXmlRpxCngOb1/HHpaMMsL6Lvzu8nxCGSa7ofF
ohRqc8AgEgf3QKi+jC9mo/27PoxnX4pbKEEjd462h0TCaxqXzEePtWsWF43bWFGi
sxpKJp/EH6mqlfUJqYPd6w==
`protect END_PROTECTED
