`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KR85CUaQ6xlLCoHRA/wXBkgrUTiUp2f4Ftczudyhtj0Ih35ANhQDI0WkOnlzj8VQ
tFH+ri3DqiLYy4qX219GViOp8Ed/yLFJaPbY4zBerYczVFypmSejQfK/4NGvqK8h
Pnq/voh3GSNrKJewvHxuXz9eZgPw1qCdb+V0MpQRXmP4+0tgUrRMvsgMgImWXQA0
alMzss02DuAb3QoBrGqJUYGCPVjTg6p6ENt+LAEJpr80kUeW8uANXC8lyIuzVtpo
GCUcTUl4MCLQrmFeL/Pdid2qZOGhZ8EddU7K1B1Yvu+OHb4lIyslkx82Iby60Lo/
hCY+70NU19DlihjldhAm/KhKUtGtiIqNfd9+N7OS3LCO/s18Ivy7225I6A3UYSa0
Ow60VadkE2kTYKuLif1Mgg0gZBquLnX6k74ALPBv4IK7LyYE2RdlotSV1NRKkZ/T
T2xYXiw80ejEjpMasQX2KlMYuXDWMg2fXTZop7158jefH/rHfJOC745MYZ/8ybUG
uuEaP8YKS0dW48gSzKh6EsCRNDR+HG55KAEU19y8bz/D1iIE8kl6tP8xNXS0edLl
Pwi13A4i2Y9g1LPu5kaH6PGh9MZPRojtNtzqWxJQUEfOhpdBPKyaxcyjJqqK/0SM
0zYJVeOqIYaq7yQpvT2dzPBpsOx4LWy3B6WhaHcE2YBO6BP3+ltElShx+bOdKPXF
6FHH7uyPt0IVI1kY8zgMU6BkNKG81v5Tr4MFnXyKA0EKrW1tEgn2JWEm8+iSN4Fz
n+reAyrRnLZZxiosgcP31CO71oeVy65nFzR8JlG/2TcQPhbqFjNenxtMrlyZqvaK
VmXvxOW5a7HCI0u0qJQbUsF+EENlVePWjQqKU0AbgGZmcB20jmNMoHWPt8G0SNQa
AFMUHATSAqfKfjok5wUIdB/4Dyo17GewbYGioEfxBq8/VKI2FVd3Bejga6MZKR9P
eXfv9c4Z2MHy8c75rZOpcyXax7p1KsBYFJYN5WJnSOvx5IG7pnbDIO89TVissYQD
16Dbp3F76PDStq7AHn5XHQ==
`protect END_PROTECTED
