`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gg3KP/W7tVyxgJCEdF0ysMekHEazTHmIZfXrKHug7jo24i6PUVJXjyuRh4ywXlxE
tSwz92Gcl7/YvdZUjz8XyjCCFQIsanlc0BsKs8kdmL6B6duz4AYO1nE8+O9Ru3mn
MjHx0UQfNA8HJ5XFal1lE4ybKvDqU6OB+vhcA7GCSbXe9+1rgrLqGm7l6pQzE+kO
/xuAuG4Op+R7mjwptu/08GEQ5R4/AehLlixUrb/osLUWM6JEHYi0AlrjKDwYInfA
WO92Vw1L1quFmxXVVEQWCKgg2wepXAEQWan44UxW8ZO/gUQbY3JndTNL743h6ZHa
9g5sTGoKNHUc33VmwtROk+z+IIhOOOlaIIFbt78ZNhtwtsR+3IGfP+pwKsnpfU7k
Jb6Nz0b4k8revEW8h1LBfcDL9bHyQ11hFrSAsW6JKYAEGUyWDzSDTk0hyx72cX23
BXmRe+pef8kP9NC2098RGW4jQPV3AqV/XTuXs5xiAa+hOe1WrADfzR007+oDK80R
`protect END_PROTECTED
