`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DakhQ4vrGzKefYP8L/ttUEO703t3TmvSu96vCrtw2EU/iRibX7KvnmRPcQyNu5FK
JRkjkmqyKSPJPR0ADhf1XedcMhxTUeV4hAJhdlRV9o+QntTSli1bricgddDZoI9W
t6EdNKkC0RFpBNrprBpd2PvEIfbI2MSR4+zfyx1xLhj4lnh/iyd5RrVfoyayITMu
8eh8/seIyTQGFNHipEuM3wS0vnKo+zqMyIUTKTUM6hNZToelXH0m2V86/Uf09vfY
u1ed63YK88FbIhwtXPmxRvkbsJeQDL1ftDcnPIaabME2hnlecZHbycZKCpaNOd1L
cxQuVUIKbzCYYNDd6puR8vd3lkrH00XSKaj+pH+L9TWR9lTH4Fk2tPJW2W+78xK8
2mljR49haeRvd+nje0XoqyB8+KP9jcn9vjtmY32+d447B7M/me7sKjJu/3+TO0yy
dMdXwxMFJuCTlBjOwHP3b5/w9Wf5qbAFusjRkXR8xm6BH1nkwaS2uNO5515jec4u
f0VjvAI3cWOSGpNcOt6ZvM6fEBZ3hUYuM07CHYozskqalrXnIraCvt8AmFsyAl2P
jEKXhYszM9J4gmeRLKzH+q3va7TbUu4Mr/j4k2qTC+WqEivveboPgRLZoeYzZBcI
5JhMivRTQrACnpFZ8c6wQmp/PC1d1pTsFuPs1Mv9VWkodADCZb3/Cr+VVFy8hosN
CqyMXeALTu5toBqc+4OPNCAm/AP2JJGwS4ZzwJ6zXZfvpnR0hQ8hYnVlFC9DLFAT
sieFH1PvpUg2bSWwkG2sdWqJyxupHjl6kTdfnZpDbtMhEkYf+khXEfxoI3jzNGmB
NEJm1112Q7GS+4LS5BF2YJD4S5oGMHt7uFEqrm4Mo14MFU3HeuCOMebQOJJ7X7Eu
DM4vmg2USCb3ffTmtakX8A==
`protect END_PROTECTED
