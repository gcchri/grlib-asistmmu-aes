`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+U5XT3eSpj3jUbGLimpNF51EdfOWH7LlhkHaGJexRmfjhMfgPyOSKoFyLjnJ4RE
S+7BO25ekX+m72OG2QtrhrW8jls0XWibFkvgI/keCobbv/31omb1J/2J4fm7sDpI
w2l6zdOXNfyP1Ji7+QflJhjIxTOIjPtJMm/X2FAU2+pzHmWmT+l61wLxwJUsoKwK
FO7vOPJXBogg7OVAPpAl3AVkaw3blfkB6GFZB4tYfDA0fRP6+BfpX5UH+v4y3IHd
PM8oEhvAsd94rmBlrA1+L1iDtFUMJDvxLPBsogaVGjvQaUSm7I8PBQhBU6mQO1EH
pj0hZcEcB5iQgxVsbFKxCtj9leXNfsQetMvL6PcOQO+CTWb3kiYzklfV1cC0Hn+P
NLX6QQTp5ipD9k0YMI9O8DOp+8u1IytF3YB28iaSWzb4IfRZiCv3o7/2aLk1qhkD
WNTFAW/KjPm0H43NMfpDZKVDQdgco8EE6OtmDU5vPgwNfq2HWWf+c1uLi99sr5eR
aLqZ/fJ4T8PEe348dGALRaAKyjsq2OWOp6MOntAsIkW5cEY+kQVW5S5hsX6S27NT
pwDOXVEKFDHOPmyBy3EYD3lBwF6PaVWPBqGR7/qwfTiDm3Jsbm0rX56PUzWB6uYy
0da4oiI9g443ZLjYsZmrp9WmlDmzivmO/ledUh7YK5aYQ6tFDvDvjMlm8+oPsdCD
va81RVUd9DL7NB6iN17URMwzGee7poKksSBUPqRK74alrfRroDU+kHYgd+ciYAx4
hxe1tsTVqs91NYDFAax3q3+3ySBgWzI1OsRh8G/rmGZHc4A6fAyN/F266w8mOuYa
DWVPZvAJ/g2HZQNwBancWGFuLCqJcklkS6YQ3cyHYmoBoyD/VKzrwZ1Nuq8CxDf8
S3wX2lW35TVTDN14M/qeqCtkkEZRGYgrEaiqeTm1yGUe5gEUYw/0LohXKcaYYnf6
WBg9oZmttcvn8qG850DOA1Gf8MNEhCz5eudeTn/TMXNbCCixkvFWtyVh59YLKSTh
RuSLL/0qjvtp7nhQzpJqySD4R3VxALqVBBweJ+Kjygto7ALhyC615z0DySFmQCzg
hgKqeHQZLSAqvSSVihuJ8qd7VP/hxX6GEAh0DJPNnXC9yOwLWZLbFk3yYi89ivgS
VKApnf8h/UEwUzGIyVt28sE+HDQqQDTNq1lXnTX/OmBUaWGP7noQ9Wi6MpISTDPT
8cWw9t56HP/nRiBXhLunVemTYFHX7R3klzyeU9+H7Dh0gy+2BndgHUR5Lcu+g+qu
3aw2EIcZzFYsQVLr5kGhSrwseIcOlwbI6xXYkTadrxOnuFnNJaHxEzFHjLdojsxj
Pdawb6FnzUJowZWNN8065iS9Cz2kw38Kf/0Ky0GyZk7tPfC+nBy9urEdG1KP9Kok
//txZvWdzEg+ivntneiaKqH+ivBgUQ67xZLbR15+lOGP84FnS4CWW99+TRqU1bYv
WHt+4zgifDTXRP28fTb+ZJ/u9+ncdfb6ViwKh02INnL9ct9qJz2pD4xsBpiYRy2T
yFL7EcoePDiePgikCJQB9XAm7ieV0kIKMn/zd8MRqEC+yVSINdCuZh94GeWfzBfL
LtwaVWHd1F4qDmbpKBwnWdjVHEVpOBWBaa8Z7pAbhFOXhWbEr9w2AtJp2mC4wMvu
UFHOBDfCX/A0QjkutwsetNStagWVHr1KokUYzb/31NgDkmoG+htshAZUPbgWfFO6
5ma70O6ff5HZuRTC5Lc7wcZJn7VNUCxurNiuzaKWGkCPU9dN+InAvlNGuLLSfFFU
lRcxq9dCMd6fo7qSiF7+H/zeSsBycx/pJqIcjDtYNtm1Jhje5HfCjWMN3k1pyJ/0
YTM4dn+747A0u/C7JrjcQGEYmWq2kKEKyH17DYC6TDlZIA5e8iW6n20RPsELYhfy
/VS5Kxe2vTduzccp3DZKHFiDWTFmaM8lFxZQfSF+hgMkXcmqsj/ZvUsIlMmCHet0
PGY+nf0WWsxidNAq13JsdV/Jti0uBb4I8bE7+3ML9etiQwctzLy3BrBzU7RxkEys
E8s2omvch6WG3j39szM2H4tBMaP23ZpR7ZRL9kCto2Hsdt7n6SvRPoa4/Fuwl/f/
sauhWufRlDxbkHh9vg3xFnF4mNe5UQf7ZvW115GcWSG7O3ys/zrcP9RO3pnkb5m8
BNnsHw79OgQ8yZ5f26zqHMUJHFwxcEbI/K5S/oM6Rsky4MZzALoujitwA5VpJmIY
GFZVzfzHaD7Ji19dv3m6uZ8WcDdSzRM2YLYqLhdWkJwCI476N4I+wmp1s11iBUlX
GwHtDOVdccu0nB051zkL4yAjYBdmnuW0roApwthu9pJ/3zpeJ0TjPmBnqlt8TYOD
BfyOaBwQRR6t+HgnPO0IPxEYc3FBn/n6Jm4DaJApybt3JjwFCOXDbSdZYfFBJIlS
wPp2Bq9Vs8DRDAw9uXKeCfm84YHam/hZ00fZ2y6PIYoo+NotEckO5f7IcRI64Qz2
rlVWg18EYhowU/00B4Xq4UzXEofJVQgMjKFQYOfAM68ZFP5fnB9f+UIv1J8id0py
DtqdDGz2mQXPFOITKY3mKeDw5evA0+I2H0Lex2j6QNvipxfm0qPyFpIb1i5d1/3z
4zoN4WcxKovjqHtSQZTzd6LjloK/MkYkahpGiDaHZIm5ScgGtqBbBCeknKG7uccY
VKqB2Amw5jTtqPdTsoxnrS4uLwe4uak5tg182us0BVQclqHy3R1G1uni3oaFmxi0
olSSorIgLXX5WvY8yGNOrF1we3DGiHwyfu4Esd2RNJun4aWOoS7ZrYWCX8FUqDyT
BtJ1U0amKpYlXEb+s8RZhC82zIoRLfTKO4UX5MyPoR2OKq+ATS1qeiKiI0MDin9U
t3zpEh5h2WvLISHyvzgPJVtyv2DQrxq/OzvODVV1uxp41VRTVHHZ7OO1RtBVQTrj
eM42PuQcZhCvIsxmmcJYjxakNPsSEjPXDTVut3wPRw6hU10ZOqDgsZxj2YrKXEtC
kUbqesb/suVkQOLwG1f/RWYaA6JjWIO8C5Mlj0UEQ1fjZDJsFEPQeeY2RO4vwszL
gPtSga83JIIMdj8EwBT9gYkPhxSfIyicsu0N9zScJPCvZ6LJyIw7/6K1rYXfKEPM
XQiDMqeDnjl/IaDwXckfaCCJru1ojdpKiaGseDfuu6sD2jby65DNTWg0y+S9Wt0i
IyhIFQS2iwWB/H37qrbcM8SN5QqV7E82Tv7TJNK+Ga6nKxifFYC71PFHXdT49mML
Y8RwDpFv/527vAH3N0JM6ki5KELXCcqjtj/Dojdja3Z9vbqOnOdjQwwJE57QbXMb
/DVEHhkHt515fIk+oSmOYX9zdQLwKNuy+lPv4SJB9v5H4Yjq7yvv3ahwGG0w2CIR
QCgGvDIi9b05TMJpxeyac40H7e8f+eJzUZFHlxrxzOYSNTfbt4Egacnu8YpSVkxj
dxEnk2Uw8rM/pNs6u2WDRdka0v2LPDjCfcHUZp8RqAv/RmVkrIdaoE92kjsX8Hag
CmnqnRo1FHFtPZMk5uEq8zhlyAwJozDGzqAHW7dtelkfs51bu3zlveOx7QIld1Ql
6u2oV9DuRKeHKpBgbSJYsCW7sKVKgY5vUm+1pBDu1Oa6Rp5tT0RP7g9JwbOGDXL3
5Ck+t556yt/nU+vYkUZzZTWvrc5d1EbI83CK/YGr/pCeWMdtDLSGGuubxQgP2WH5
Ifc6t7n3H4g5n4I1uEd9Ru6SQjAGau933iq56jtMqmJFGt0wnWKfA3M5zkcZ7u94
Wy0/ccSbuyovJwdkEGt+MvjbT1AO+6Rxmez5uqM4dJEfw/pCmzkaDrSj/ur53UqN
Jp6RZIzMuowGk+PVRODEM7UASb4psdKcVl229Oof2DvC3SO8rj4PsNiv3BmmUpqM
JRL7Q/lM4RxNEVlpK/p3jgELeBkDGvB+ABiIPC46vJx5GHP1zJygUl79odbau6GD
GFSg2+YRqPWezzred4DXucymMxAtnx6/Ibnb/J1t5iiuTVlD7so1rlGe0OBltZkT
9r0JuvQ6rooBofLk5sBfeS2mTVWWgNVazKVs+ABixG6m5ODhki1d+aIIyGCW/WQl
QtnL4yGqXM4xuf5m0Cy+M89zTqqNvKYVz5PpOsh5zUI3oE8tO7VPPzPaQfcTaAU9
hwxznVhsXiCZ1bzbwztVgP0+No6Wf/aHKTcceFWQwEAxmE8VrWFt8Zy7GJnPs1fh
BpiWCO69rdQdZrMo/PNHHwPE7zS8vI/ELWNLqzDd4Z3DfqpFNYpEx605VDOSknbe
XoSI5AKV9xg9XVcuDip4v4g6Z6JpZo4fZAAOrTfE3i/Nv26PIf+U0+KwMVeKhguv
vQcjcBNFQ5O4B2BAAEmRzeAeOKiZbZkqaCP5SMHSIKE23n0EmK0hxCX+8njEGArr
6PLtJNKI979iX+3ETapLmLO/o0pMoV9MNwSP9FCOV2zAayaBpqaZyyVrcnemvNTX
U8pCFdyTOP4Ew9Q/PcEzEp9V4kusEwt33AtqI7LT+yeYHwj4RDrly+VfHAlttRsm
I/o9VuHQPVyYYzq2FmIn5NwpZXVE847YqaBMuqRon3itI+6hlJsfuFDoHd3K5eb1
q/oPytb250izK3fSEPj7Q9/gZeiZkLE5d29dPlPmmT+kqIDSjj26ayIleB5cgtgG
hrzhzVQ48THdi8D4FXGsJkLcrshOfaa2maqcc2UMk56/TPSYr4wFWCy5CII+7a8J
PikUiOK/vECXex5QiZhsg44tUbPttPuex3TIHLF/AEOUSUxuFX1R/BCcS36PUc1f
CpehbiwNEEzVjnfi2LZ4mW040++Wg3jsOmkS3BKlULrH3Cb8Y7c4OjVMiyeUB4me
Ch9rSE/emYfRy4BEGEsHkcsOAdfHZ5RuKZ2A9CQtL0IFG3Osg98qlBZ/hLyQNHWo
kzVGLXH7NhMjeepkJGXUaptfvab+87Vzu2pAKf2rKCt3DZrCMTX0kFgQQ5yhWAZW
CJ3xEYlkj1VPEOJKDhX2R0v3EUsS1009yVnMhUV8y4rtMcHa102REnT8mEkhypJI
BZO1Lu4en4AukPHoKaYsvLCpwRdlKgPvlJz82Fbz7BLC0tqCPTYAP2RZKHi1xcu1
9evPId0LWFWpMPasOsf/+UlrpaFM+lgMGE+LkxEMLGgPUMfK8HkKQwQ5HwBej/s0
wc8j17WnrMgtzlQGwF54SetHx4fgZJeJaGSNEWmSWlitfjizxRf5+4N0oQX1abOD
H6epQZl6YrAkgZiFnhsfeuhJBBoknET+yIZ8bkPHuR28dwjYQOVjsGI8wNgTdnUK
jj5G3sWum/llEC/rh7CZtdbwlcNCzAX0oVY2bjP9HBXM4M6HJhr2Qnbz4J82wiUN
oZw8JQoo4/ClZx0VBPZCj5vrz9YIn5N/naBvNR5D2LHuSjwwA+dkEuN3sPjMF1LJ
DrykUzhmqJOXDvQXCA8//gYak/k9Dv0rFGfnchciQjs+mJWwTsYC5WcC58bm5Sp1
fRoXhUx48Em4s8vd4YtlxvpST2146P+PPZfRpiVQKkHQyjgv35Lj3Z+E1NSIr9d0
9hoSZJXnd1ONmUL8go7+ocevjqbngIuP5PnhPAzEfrL3+51aGtGt763BEPCgYzIt
1Ucjq61ACpMRSVvtnV4tToVWG+fKyotz7s6Barh4tL6mk0uC+E2Zbq+qAX4S9pVb
DXDGwS/kMnqXiMKnai5IT0EpPVB89svKclyLTD3aRy7iyMPyOa5mMy/y5dAUFzZV
M6ZDOlhEP9tOhO7JetU5g4Ui8QCH45MkJ7NrRWIIIFfmYWGmZG2nOBABKtlg+zlr
KxUnuDdRz+6brFBDGUl3IHtf2mq4GyKVbsHCOmnL4b9qCnxqPtzdvHpt7lGmKZ1P
UpUnDvJ7TyFUudkYu5LfDmZ7L8wCuM79byzIZBeBOE6fFrgrnaEK8dgoS1L3g3tF
snP8z1KWYzwizCf91KihIB+AHlxzBRmcBRRKRHCxb40HWfdEFrZfwSAFTaFVvRwp
jEQyboaaTedxuzgwlu/+rsQw3yNzZM41s7Ciw24scr5PjuSBYOEEeV47Z7P+TNCd
9BhRcIGc8PILVUXE3PI8A+6gFUjE/wLnykdUnmSfIS7gSYNumDSygwsE+ld3Luxf
xl59WzMDdk5td2B+PoTmXLzxW3T4ci7lj8BZxKmXrPrxvlCnB6geZ7B8vQLDx4/h
rKIOXow5HvY/z9UDU4vzzyieT7Ne6q6XxSIo7YWwnx8CDkFYiopkNge2uOlEXku3
93cFCQ4K+j1w+KSBjvwEky8wAbuJuXIZPFfmWora7FKSD9m1sPY/SS8vMLqwtoJK
tjQEVAyWFQA4VeRdQIhgZl9wW4RwyI9627gk5wS60+rZqLEtRdajqa4ptG2jX7dL
llZ5jsacaHntiZa8la8CPzhYcWXr0/qKiQBUObKAeJ5NrFULL1p56nSnNxjyyukO
MxObaDzqDFf4wphhMdrZahLOsxpyKnEhiRM6M0I1qH//ovbE52TO7XVMYnrg7as8
NTkxnRKgdkLdV7rkO+dPp63C5qSZEJN+kqlG4OxwIJbw0KOD4KXVxsF/RWj2cYEA
Z1Mjy6PVkteFQNTVfFTSLziEizRKYYN14jpMM8MB8VDa0MZYyE4DICcPKDoxzctf
GsLr8NMzmYgHvQuTPPZASvIoyEzDDSRNHs3nwSPvX8ak0p7b/TalqASitoyhdmQl
jzneBRmrlYv6GxtNmEgakHBCqVtPmraEUKvlDASMAXhTztDmaA4U9qTpsSl7XDF2
gnyvbMIXuNRLbLTSmXIY0QvRMPMIMTD2kb58Mr5vQKLXujFwyCyo5r7JJqSaJCf1
LOnUAQniGjMQr4Kh/R2u/VMFrbfae2IQYYoMeIgxGbp43r7BSYXpOZoWl7RYOl2o
maFxuzlzL5DQQqi1yhFkQGOwQbSyVKLtD39Q9Phaar9t/pvjVVFj5szhOzum+tD7
tWNWcincrc+QkSVncIZGck+fsdv2v0pUGt01r2+DI8uPjQyPKHYQi55hjDbBTPf4
MZ77dE0Vt9pkYkweWyZo0Dshsh1tCcFqFphwxfrke8ZoqSP0qW46/loB3mCN7llV
0leuvU9TN/PxGJwPn2U7EVPNtFLEp3s4wcv/EQyCOPz/dE2AeSzV/BFvOYeDTeE4
+coCrAZhjihg+ISdPHaP1vLCx9GZRtmvGNYJKK03PgQVzv2sId9hgSXwuVDVd1II
IsIJ6iy+sPQpIlyhPcz+rfUeXAI3zL6e95kWfQUwLi7zfcsqTSj5m5NBpa1GzqXt
S9iRtEmFF8iEPRCuzEoPqUeifLuUlrxpml/VdWi0Thg9q/+magCYArktKnid3/X3
W0CCE2WNBZRSK6blC2yNLWkngkw1aC3lhrYSmu1w8ivNlc/yDiRXCQQa4ww4V/TZ
TpFyRAw/SCOPM8jWw+4OSHowRkQEEWGZlTRnC9E1fGd2TOF1Pk2AzRbRvE8o3+Df
1FAxlpJwvPyV9yxCf0xpsg5DasVvRBM+FVQwULoDm1LFMB8EOSKHqcZro78tGQfc
FXdXuxDseiBqig4w7MN/sIuZstkt5J8vjWxMK9PJb7+QzwXiZwR4kxTRhIYnu05B
G8gBuIBGFlOVXIjFCyBrtGHZLd7o3JGeMHhzd6crYpJvAORgQX1iW/dpPZDe+sT6
J2roTi4356K2w/4Hpa2UCMs3URDHP3z/aOCSkUCP0FZuwn0WFNfZx/aE8GR1UgCw
41oL6C3feufdAnKzi2+Oc6btnqNfPa14kc+Z6+lMVJlTMjS2QBEF9bfqjmuUPbjl
2fp4PIcZIJC5AFxKA+lUeVYEyk/w3cErlcDa+99n5WsPpx8cGZFlmCo6KFh2ZSwH
dUsfQAqhx8FDU99VGMqfflVNewSQqe49bB5KaSemPvR9tkX++kl0hwBSkFQSIQM9
BbhA1Gy6eSHb6q/g22ivNprguRPWDvjIuuwvUkNGG1tlouU5oESkXOsH0Zn7cLXF
SMLiswDYjUOIZ4WE+umsthbxmQ44+xeaITIWsfWRqx6sjOOXvx71ypw2PWrWWzTI
TnixMx868zBM7l78urOpYqy04B3rr92Ok6YfQSIUtt8cooi7VHFGSp+rZaBGEXHH
3iILGFhGCyS+Fik2CWxAzbCDDdtqWxjG9U9EJi+7Qf3y8xRzo63dnmEH3j23XRKS
ylC5UXm+UBQWMY8LbYgUcfTYXt5QuNH2/wckCQbjMWmiP6J7kKuKQOBXWAFlsJqK
NQkn1wHZrx1jqRqyOkqx0qtrOiU52M+GvxHYiQWyvXa8W0EX8racXU6/iEgEWaQb
jQnYqigHcWWvrTH3EG8I4CoCioCooVO3HTYM3Gy1QyEUN197A1t2pJB8DGiWtofH
Zq6+RAmRkPCJh1ZyNqbsw77ex/jWMYTv7f0L5rB77EJrQXXYeX0esQdI47pA+s9V
XTVuTuSrqX+7P8bz1e1xT76ngCA+9UDEM2kX85v+4qIvpyWG+turH3YH4B/KaiQr
U5RRB1ZOcTaFC9Pm5dB7zfq567Sm1BKWVJVg8qwLtk3zZWLZy4ZDrwiaSYKryi0R
ctbemcWkvL7ountKkWghAjxlvxkcYqULjexl2djmv9N0DuIgZJGAKsFUv29NCJCh
TNZGYEqSu/ru6HVpJwk9IgliSPmbHxEajGQbxiBULpTS84W1BPVrJtSeqL3cLTvE
sPKHuBs/HAuv0Lp77kwU5GDUdC62GJrjs57yzrWTz8Kw3oxNir1HdGZkWUqg/9Z8
v4wVkYUaLdceTZBYpwJe2d9raJiXLjxl3VSg+9zW6DMExO40JmRVQ9KncPAXQcNb
ks8ttS7KW8lMnw8FusDVrITisf1zM7fKX8nBDF262P2sxsTFJd7l6XifbxdNqcrF
W5TmJp2zPIX8a6xHS1/ztpazODI7bHyFqp4eXFTi2sERalWspOsUn2w3Zx5t26aW
7Se+lpthyhEN4I0vRpPfNjb31nwDRNZgjni3inFvRaIP0+QRBLbOBftS8LZpItNU
81+QIo5kXaSKMJtwXwtUQKeOC1LIBX/f9owGBnnzE65tOl5ZrT9FZEAbJL9LnO1T
pNKw5f7p5Ol9BFGyFRcxU3Vbc+NZFRZcL1qJLZbf+OlHNG16/Rlo/LvGvrkvpp6w
B0wqyI5bFa7rMvEZ1q6Z30uQsxqAAAFtsVGDRk7FgBcNVe+oAN7D7ZhkCfhkhUOs
G0NmGklt5zwMpbhB79glIKMnD1O6DDzLtXyO/Dq7rY3nccj4XURcF4ZX/q3A07GT
c1ycF++RygBFcOTaIh22VzmH+9ZZhg6+CxLBYE/XiTWRsd0N9rwYCojE5jfauvQ5
JL7pXemkXwJ99g5Dv5EtEY/qIt+tPPvDz/a3lJLA1h+riq5y6UJRSx3l1IyfxkX3
AERiJFjTgvqRQSiQ+yBq0J5Q5iffzA5Z5ibF8f+VVF2zeQAQJW1P6Z/6BfpGonVA
pgduBvrr8/oeqOnYvJ4KKKpaJvlXRaL6bK7hQ6aYcQRuSh1GVdHMQ2PPTL159b3x
wa2dttmmqXT/fFqK9VpYO2sPg8LQ07DJ4ssHUwkp112AASX3bOSVyfrxDfXy0oXX
vewznc/5GAzFNi974p/LV8un3T5jdVBb4CZFtX25SrJsfywN6RSQbD4/FlHi180s
8S7lQvNrrPBQIWrUBjuNZP+f82dQPuLyfZsh4CChCspmjwtWFgiEtTwaDVqpjSS+
VMSCt/Gu4D9y96u2X8Y9lXkkc3NkexuE4XLtM9HcnU2Im23/QRkmkyNGtp6asMwK
MCoL5O6phKbv4Wcq4yk/vDR1bvg4Lk3zQIA0Po07SbFjwGd15Xf3SbF/rTKCx2yo
mBQ9e01pVTCfgobJ6jBv4gSXoHTCSW0BXQ8+FEgR4ZtZW485E9O7Mqd0CalbabdJ
CsXo2mOrBMULFHfPh2LNOfiSYTbs1WARQdNncg3biPFBwls5tZ5v7XNm8pNsV4Hd
HMWnJ6jlncYrfVpB5vC+HPeblUFB3qBwcbHjbLzVnexqoijW8drO3gwicf4E7SSC
rP1AvLMv9k4MhYCRptb/RNyjUemCX3AVhdwPB/C9AsgvSuM1sOmnYcfvLUe9RSq7
RexU536IzDvfflQd+Vt6bDk/z0pid3YRG47T4xGIS/PHbpjOtqKunCwqhqfM6Tki
sSnfq8fH00XLLj60xV6REYXbHwsxvGDd+BBWNZ2zXyw2bUQ658532TtyzhSqgu1o
QE4231Gt61trLtzx39kOcyr9GRUDlbullan5A+EJAnJai9LMamBQP8jPa6hHESGS
1rHcar55ru/HRHEYQFQlLqR/NSKWOJ1OQzA8sgvFIfQoZEAxfNaLglWHQ2TECMoE
+TgQGYj7m+ieCTQARxP8eb8Q/GKcfJG6/ycA6WHZrek5RkMHQzsLvlEt041SbWNJ
a0h2Huzt5u6y14n6eIR9gdyZEGliF0JnH1dyWIJGs4ZDGsy27KMSOqGcwa8UUMTA
9fxfPA/2tL9uaZPKJRCjpOf3r587RyevEtFPT4ELC9/RmUENgLDArGCRKdt3IOJO
opZ23HVxChJSbHSe3mt/IW3+6rYbshORDEE7qc7IWbc0I5MBvL14BYnXK7y1mFq5
BosZb+QIB5j2yX91w+2x+wbsAv1dp1k/xClCeYvroXUlKRvKp8cc7hBIdchakvlv
po/vhT+ity97OANKMQFpa49ojXYIHtF956Pa9evqouOgNjqJOZUMKmqwBdmDR038
5KgOQrwaKtc1X/PLHudrfrzOp1OJ+6z6+Vc4L6JGNEKetfW0DQRJOc/bWaebtu9+
ZUPHTwhcMKd5P8sVDdOnQuPIKPQndexzcMaQsiN1uMA1ZprXEWnu3LWuWIliqrRy
6gbIyvh2ACsa5PUHldkN7Fdy30UdqOJyViRMyT43uyMeTdVd5R2ncutTH3etjdBi
jUQVcqlmZ6S4lSAShoIQgGMqMcO1VmmLnyQYQZQaZYv0uy2XFns0VNnOmFpCkmLa
9UcvCsuCbNPvu/g6uw0Pmjhl+9SkFZYpDmkCdCvIfFW85Ko6IlKJCPYgR+esCYo3
dmmFttYEjSKnCPZm5KyCAJQT2RTvYHr2sQOwqwnunxzd9qpTBkGLVkXZnix6J+Xg
0DezP6+DeDwRFz0IFHvuSkGYyaV2NWUgHLRNEGWaBibQh5sZmscDf9Hc3uCw6fGw
cqtlKbmSLHgr8TTusqnUIatDCxykJYGPhFmJvl22xm1SRtdzXG6BZvkJNVbCrFwp
z5E3nORr792CslMo6OGx7TlN8RbYajf9fIPUPkCSxDeRx7lYpwv+RhLIBTmigDuO
xIas8/4JobL/kz21szcI+0a0gepgCj9b00Q0uXp4S/fSv6W/+6KBJyQgpaP7pdE3
EdJm1WXiY2Y64aJYVJoozniRWTiAzC3s6bQqqDYR6dlZKWYEM1jjK8nz6/KTos0V
4VV7XYMRTmnyNaCaxPA2iUK0Fp22iicM3RCxA8liA4FU+402Fkc9WjHHugZ/eC4H
8gMRZWc0yQ1MEwDqj5TvRD/6KxPC4zNDPm0NuD5Z1GwoyN28M6sQAReKG2+h6k0A
+fxKrW2JpPblJAJCUiGNWhHYMtMK1bOwlrCfmqRXbq0u2IdE1Ku1iGmzYj0KyEyf
o7IPz6/BdIsfVINc0oiVbo9vOdxo1e0nv1AoRAxGVSbX4+HfZwlX4DdcSdk+RSaZ
epjbKqmxkCEok872ENnRuod3STRrmEf4bbk1zQE4jza1D9xqKojHJc+ifITh4Zk2
u5kw8Mu44pUEuok0nt/K3xBYE94Td38gy/jUCpXMzn0dbXHfSySgR6UJ3v4BSu+c
na2NFcBEr4U4vDsiyj9VNXTRXAFkTOux4JJ7F1htgJjo7QozCdnA5MS3qQQ5Agd4
MBDhe1jlE9sw1j7JZ5GQ2SjJEJLS9L/2ivKuWYU9A4+pUyP7O1fwlRdn+EH5VZuc
rHs/7NHWCvqk7N/1lM7ndSY2ed+mVmZfQrS7xOr0Owir7BzzKDXOnSJ+wLBMUcGY
J5Ojh5ZSl1w14udpgdjLGKtRJhAtjDLwTOvcm6qcslKolfRLekcVDDjCwU5mtv0S
DkuN5Xqye2a7Z9/ShTHfDPnFUaqVD65FixQyq5QI3tT1zO/PCMHXeWJudEq3smKj
+5S1M2w1OEP6E5MZ5V+WszEKLhQv2MhYTdoGf+7Hh/F2vujq1lRqIFJdxcEoMEhg
qBXm2wBsZtKdFJA3l1o1PdLqUWmcXVutaJwIJNhnJiyYfQmwKclERBFp1XzsiX+M
+Ifuk/oHCcVcaF/4VSmIBM9UURVtEhVv4sPE1yr/c67sApDns40e7sIDcOgoL2pS
SEhdiomo2lXb54avi6Vhww==
`protect END_PROTECTED
