`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p7n2Gl1I7DtTFlgQTClbw6JZVflTpTFXB6PMKht3Swok23Z+CPjQZIoYT0tLdd88
OEwHxrwmY8jtK47aLErVwbZY6UYcA1ya3aDMxgkxPOHO+e9xIVznUmOm1kGQQx9r
d+FIpem1VHX+s3RZ8lRfHt0k8CMlTbg8DQetTFgVb/UInnLSMRDluhcj+UMPzWh6
McAHsUeevXnzBKqFLkeqCEJ53WgGoEq8KAnKO9mhUryBrR8KYaH1Hn8IkNCp5dd+
PPyLTGf6lLr+jBLpa1vBSit04b3FOVeV2dEsC0Mgp8DIqnmxmGdQher09NX7Rqne
`protect END_PROTECTED
