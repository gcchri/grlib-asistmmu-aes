`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tx+YRprtMDFCijoCw88+jtdmvdJv9CuXIrd8qN6l+Uya4yhMCFEPy8YQaO6F9b2T
1uC2P50tjA5YWHTvGXdtgCJg+yzhRVWC+XfDxbMyK2DeLjLXcPklQDj/gL/MNjzZ
L5n4+7hrh1+0Pf2RfXUJetTyPwk2aKWo2/nDtpZzW5RJeYtP7iIPp3MgvHCyRbJZ
HLc9qg/FuP8dpX/IYaJgSJXh1O3mfAUYr+YsAVUqPA7ycBJCW7RT/mv7TWXeOWYJ
PtBzydFDvRO/ik/tyXZgRdExBlYSqEPWK/r3zQLw0kf73Gs6Bf9HOQTZA98yx6Wt
ghcYY2Zape3BMGKj0i4Ufv3u2NXdg3UzZ7hCg0973UXjbw+LNBYuWVmzkwuGKAyZ
kWGhz8avHV67K2+xdqFjjbm+srlnPmzTtx3gvJ+kbH+kOfxlLEZ/I3k1PHW5dbjD
ecbDWjckip6+dFR0FlMNQK7kWFKa/tm4H7svePnWbhvUVBkU7u2N5/12zjz10PvK
anPKsIrCVh1VYbOMSHmpBY71zupMQEaWoeRRgDbqnnvmNKLKJUZgHjdf8tb4V5un
1ZOxb0cf4WxKvgX5ULqxfnNiShj6Vb7yP4iznnh1Aya9eO2WwTGsjBwwYeYCWoRI
qmbmaGia40mvinQJV/hAyp+i6bYwqiYlbfSLJZ3uHOXXmQZAw+RZxCc32W+v6BTM
ZBAf+eVTvpDmV2zQMleaZvAcfRoCxxfoH8Zjdtlfvx4rG4nP5TmKFR5+FISJMp3m
nuJ+vDrBtBPq5G7TNmwioA==
`protect END_PROTECTED
