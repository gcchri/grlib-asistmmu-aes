`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/wWblpWtfE4fj4r0V7j6pmhTsp5lwsj9tLK80wgXrthzfuq13FfZVvh20H04MPAt
oYR8QjFW4mTXo3Tu/S+fUyqNWGpKYM8CxRMIxZcaVtyo6bVdJ4Vn2IhKHhggen0Q
V7JSBrn/t8cQYkmik96Do5BLC0R8pAAOOyEH3RkBEZDI7080SMDA2wVy5otfB8U+
uN9Z32pTON95u0ZfbMifdWPBX1SaiVbuJtcNLrANyGT2f0PRXKAB7sMGxOUFX/Z0
vQXCvo7mritkzwNr74pZLYK0HoCFTpm19QKJ8RWwHyZcp5S3HF56oCB3zQmMSqii
`protect END_PROTECTED
