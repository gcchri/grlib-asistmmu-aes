`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gInSNp/xvX4Mpmurjb283Fwhd/6bA57OQ6g6bD3V5D/q3ta51B8orfzT0CaSqQAP
YUqRxtQ709dmuHVkTjsp2JOVPfqeyumj6SZBr3T45oc+oDDhSqAYeIchvSs8g1+v
smh2AiR+5FEd+6vZW1FfsqF2Kdght3xwMHFikkKQ6kBEDgzibmo8/7G4wywyVce5
Z0uoNVvNb7YQy6LWLqYb4W8FpeQjWLWkpTMNbRrNaC4o1oQb2pSvAlEOHfRW0im2
r9sSMq4wK4/GK3mQG6EdNw==
`protect END_PROTECTED
