`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2m3SrG+YrxtrcLFNqkjQsKJpED9TU54nEMugkugUQdO/XvmLixeNtJW6Ea3aUeR
6hIMmdvfitjU18M/zm3ncdvrVPp7RyOBgMPUu26IJf20L8d4rhUNyjqFumTTnV6F
oxAmZofbjavLIx+ClqI5VNFeNvwX+au/4jxsrlISTS6S+IZSl9tIGtMBDvzysjoz
KAuib43pBYjG0MhneOLKFngiPfscKakfZ3F4hfYEt6Ud46Rjx3t0WhKJNXV5Fagn
CYfB5lh5JEmsji8Aaspa1pP9i3khlcu45nAPhhMJkiDS27lggpQqdUJtQyawkV/9
ejgbwN9XjMXjPx8OKb9WqvfeoZXD2POiCKg02eR0o/ofnf0zdf6dqKyo7Z3tA24C
Bofd4Y+NkKOpHnOFslq6B36qfL8Y2NnB/c+4SViTX0vp3G0JUSgfvlWyNP2NXGE4
VBE8+AwPGGm3wPQ4B6D2vu9bnhLAGc4a/KP9EzOfA9FhqxO8zKdSbTZiytzVdY56
Lh5y15WLZ3wBfCVVCgFzKGffsijJzhXNLAgd76p6REC9XO/3ekw4GaqvpyHbD56q
N8ad54LS8bExdGqMCv32zaGfj2WJvnFizgpxC1cVwnh/KF5nuqUOTv7dE3Rxbcsm
ZLaqYA6d9VOWB7aVAGwPhWnfvbaDpGodHQVsnLDq9c3tNGQ6Ubak0KDY43RwdCKF
hHOeALoHQ1Z3dba9B48VcJ4hU79INKD3npvEcW1O1TuY7vAqyGuxPdki8hO6YqtW
r1Gzda0S4Fm2464vZietwVY2WmYfFolz2iy3ey8PaBo=
`protect END_PROTECTED
