`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ms8bq8DDdfLcBzd3nJmc4Lg7238hjtt1Ys++mSlucPWxVe3ZZ6NQ2IPzQg8Ojpbr
vEQH/PWBqlXsXo0/7VTWZ5UNyoQsg3ZiezLdGbt8n13iJEOVFFdTONR6RyYN02lI
7L6VNY8yOAPVFuWE5tw+I7OgNcDdP2EInJfVFThVcqT4gZ7862+SjO1dzQfo7lx9
9p3Q8mh5xupcqUAe6WNlgbIM9rfyCycnVjMIm/6POfnXCVCZAgmOXhfA6XLedKqr
a9LM9g+WL1v2aSJf8VwiyfiYYBhclXPceomvUDJVojrn6348BC3X7durIMCFJYiH
LxaTKg1umKHu4v+EnpzFI8eiglFx2OF8GsQs6+XjBh6iRtsbso9z0Urf783bdxYV
jzTdlJxrt9WWn5PgW6Vx1nhS99LyLshSqVY0C4ZhpWLVe9EgoYoZwTxVmw7BvqKu
4QuRXV7jMaDEK4/zFiQxOV2QyvnH7Sshd6IVplTlnms=
`protect END_PROTECTED
