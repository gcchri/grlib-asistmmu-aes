`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6GKALTG8B7rjGNB412sXy0yzjwpuUtWlNhtpbsAcxxCp/xrI9Ga25+2YsOWXT4wo
vztrKxZ7BEE0qTAdD6gwTmewAH4Nfs6FbHGk2eN23oJljKekUMLlu48yvLnMY2A1
46YOX+3PAO7mT88oKRGlUNgahdVQxIXUr4mnWPggklNl2IRfkN64mZsJDpuQoI0B
52CwFZW19smhDHz/vjpoA1aryuyiP6GNbaP5sulkVup07xaJTLvvSBIGlqIik80N
vLut769AaIgQ8rNvDyCfd2rGRRpN7OcmhTR04Y+OFHFJTbt43c+YEvyfoF77dgyM
iOxCbFQkMWnx8fmpdbZIj75eHrbISdJx1szRizUPR8MzZaF+WtGJRHb8tsbsMStu
3AK4TUZ2e6VuFqHrhpUo7cbvkedCwAxhiIS+v6B1RH3mt8DqhzTTQpmws2crRWV1
rHUL86jfhUhEfPlBzvfQO77EEzOD032jov5WGuc+ssVLsmfeFl1J3Je1gFXwHEjs
oh7wmG4l6/SMy8VqpcnHEtW7d08PTjLtXoAL5tB4+x6BP4uLdUKVmjurGpz6WciG
FYCQK+1+9XEkjJpkDkrVmrjiAEUMdQmd7LfHIFwFldb9a7Ip/4JYcjA79ufaTk5r
5sepLwIbTqLuBx13kH41V7vFxrs99ea//vKN5acWdTHeygbRck56oRLFJqk2mDcw
/Mmuefcz96/AkLspURigVcesy3SsOHgbGhR7qSJTcUnxguNnH254bn1Z70RrXNj/
AoNmb5RJm9hZKqSkYaXpoxXSo3rpae1TtRSm3wMvc1+nrPOhOERBPATBRdoFOL4l
8zQwUI1BCYs2FQgRlWPXEnsRdRCDyC/Wp2Od837Mjc2Z+EHnN15PV60DKjY97T3+
f5+XcsK/B/tXJPoaAWGm52Aylzwt7edZQ+6QMTHnaqzH/zKe0xwICgbWszCrvjjO
ZWpVQTvnBUDlZ1KcYsVsCtRvV9KIR6q8gjpzQ0Yk7//sR9RtQ+bo0rRe/UM4fHXo
2kMvhF5QJMATMb+rVf/XtMaOYpjf3us4Tbpf2bBEs9GL5yRgKHFROAxttEi+5IzO
gkHjQ5qxjNYrLAjviPsHv1oSH2nSlmsI518W1Ur8JEI78q7gCHPADZYXg1S0K+PP
MWI0SW0QZ8XyTdL4EObZZ7x2VWMbs1X6QrQoIvGPs7JzmXsxydbB9lwyxkMV+39N
vbQ9Nk1vOE13CVbBv53kskebbQTEGIXftQNbKjD+X1LxGsuKM8MNvIbez8HDv4WY
I4TVhnfFbsryzgJ5pWVhtfJm7sT2gLjJEXuPvVJNgBYXKr1XEFDlt0j/MgtQAdrZ
jJ/RErfgw/Wh5XXN3OPm1te4S4Ozc9XcbYDudeYJy1na3OVtiYI7EbuuRMSG7SL1
yhv9Q8GjDh4IWRnpZj61eVUSwxEqjjzwf4B0FkNjEGoa5w5Css5BSMe6RDc5GCUA
bByBAyzGnFGV8GcDS4kMOMUHmdzrHIupQGdrnwJDztZwlmu1SFlEhaOzaSetgEOF
kQ5xtgSWCIO7hyAcSfTaKQxmi8VvbnEuZZmepdPW+Nk8UBW9Tgpfh7deM9pRqq7P
cBvniA9NccLzsFQp/+a1uclneKSrWW/gGGO/dDSZM9ug91B9FnwquHdkyFZd1ttB
aX9KnAe6mnFqu/aFI43aXvbGPEWGoVOuDuvrs2cfg5uQVot1cif0i5H4KsSNN7iK
2wwAC4tx8JKg6oPf/yOmOQX1+bnbyLBMJZLWEZYJoMssylSYxKFeSuN/8zU0PqtL
n6wNsNMZnkMRkQfUhTD6pp1MAtHcLOXQ9LhlaaDmGRu+Nk4VdqGEG9Q07/s1qdno
WhqV+cZusr98kFCi18GyxRnnFSpsxrwpN8omkzzrDnKl6/sQ5UMXP76jJyLSznmJ
l91Ak0C2et7V9pNhAH4oAsSIaYuVdLpDQP+Xe5BAtlEZfUaAonV1uJtnm+vSNYQ6
Q+OxcM8SUiUV+zMUtXRdgmf34Ot0jBfYc8MEqQFO20AqtNEiQ3gx8ljDoFsEWilQ
10nSieocOAiXapcfyvKmVTNpPYH/GTn202wlIdRQyupbN7fUaCTSYMUUt71YBHm/
KJxMzwFTN0eyM8rIMZAvAQFNAh/wAQiqvcHFUdDQQnUM1lHUy1dq6y6OQP+j97xe
K1Eg3zLiwDtkUYVGdjCYe4wlh59FLx4JuWCJ/H6zbkKAV2ldiTAtMR01WW0MGfoy
3Ld5mtW0aQEpK5yihTLedAHd+1JDPEe5CzBFslZjj9aXAoC2a6mCk5us52G/Zow0
w+sD3bLH4W6PlYnIlQxVVO0lckj/Voy3CeRsQPqetnNebv9fqU9+NpC03DoYVg7A
UvrFhchjYOI1pZAO8NzkNNgsIup7m4+oU/POH8KD1n4rkXfXILHWLexLDDQCpCRK
4ErLOsp5Z6llcX6lgmFGD4QFqDr+9DpOcPaZ1zlIE0n0WhpgrNWmfRdKzVFvqu/Q
oXy6jgCk00s2sfnvrlWy0b/aMGLOV9TEJuw8MQyB4Jy/AaHh5VqmAEbw9hOlTv2m
XygicV828570F0ws/rzbkpN9fCJIvxjIr6ewI63IYmGPyJvWWD+jX1MYp3nya/t+
K3SPPXqkl6EZZIktpCZL9Y4+RM0UQc+mUP5IeLttwThTzMzsrBsK2f04LOkV6//G
i37R9kczBVOw2MpQ9kXBjqWmSq4neGUZe0IlnespaHDaa4u/MRnfPV6C/0tYUOyx
rv7AFTa6UAzCN7o504dyoqFrQ3ZdstGAB5JzfA7fq/SsOvL1fLAE/lG/N6FqUgro
DSU+cZ9IYb1YrYyUOrS0BF7+/MkhaTE73URo2FTWzvQ=
`protect END_PROTECTED
