`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wszg0U+2VzGyIlOrgi/gCEd0DRTM0SOgM5FatN5w2DRdQm4zuvzP8173WlIFRyMq
MzX6/YgkOH+oaIpmNAZ+oCSnNHPhvpXwZn+eb26uj7c91ocV+HBe42/qdgxX+RNs
ZUAy5uqn0Nt0geuuc7Hm48/w/2Ar0DJISYxRGNl6heI6oyDwAF2NfLpbUNsWUoRl
dyFJmkV8dJ+tNsZC6y3btGWHYG16TxKskj8aR1j9nBfw7rXMY0wYxW+j60J7TYSp
Mi3vnYljVpgbQcvPLk1J+ktVgNSoVOWbsFveutK+vFLDaak3FtJH6I7x0MREi7Y7
xP8uIQmMOyUQu0EXQXxLZpogy+p0154rTGyE2Zb1WATUbpSNOYJEJS7SoIVQII8w
w6m9d+TrXljKTAMyKW7dayZz6q93K4U6dQL0R/05WooZ+Z1NPBPVjTx2+fXBkkRY
cIUvbiXrIV+EUVhmheoKQbX6vaYl58CJ968TV/5YfT54GxRi2wjCre/VUDL2LExm
CmN+HvXejaLCcksUisqGhhUK/O67KwqoLxxB072iV+NAoXvlyHN9qhIdzJUu0+2n
wkjMLTQU1XNa9Pg2gCbHhwjOhpj6SpuCHLH/n0AYiP0xmgYM4s4RRZP8D7t0A7Cm
qfAF0odmhpbP0s404hufnWdv5QjW45x1Gch+wlOFVWysWtV4+/1gM3YfqwkICd4n
ehOKp29Tju8XwkXC9GDJQ24XOq4zaTQa4HeKhP7FVcAnuJpSyeNAazsImE1WCHU6
xr6vOnL8EJETzNoHpuFKtyZw7L1CYKV383DrykYtAc2dduLt3QwF2BaKXuDqJhqp
SKP0hLsLVEBOMiL5vdlSUApQNf5AJgAVz41/8QC2YhhUmazwuwTDg7b/5og7D8V3
hdBhzVO6RgyCHOtHlsNvQ2eVpMYlVq9ewOrLJXWxWhcSD9V8X1CpzGzpxXY3/WdT
ypgecuimGVFEQThm+f+/cWI0L0FtmDbRJdcb+3byu3p1en13neqtMESN0jyvmF9b
Vkv7KaUwaornvOqTgF1Jhp9TuAKXSaiwAcW1C6j6CanmzjiqQLZreH63cgxW5Wbt
jWMbs/0L4VINg6Kt4AvcmTGgHAnYHUhRb7q6sYRHD3gfpa60RkBYBccXH2bmhrl1
AjNecu1+BOgLlnlCp5BY5AvRAks+lyhmsZrmMCF0UgMgbxLq3+FmSogktCJtMFCv
M/M40ImMjF/dbzonSjozq1ut4Y8lzX5ylPQJNab3cHcHdMXHZIEgXR6B89gu+T3O
Cw01gdZmDO37+GDUum4jyniQwpdEXwvkbOe3/qaOtPNC1C7mYlusfDBpGdp6h8lK
4HsKRW1cSVdZQUY2Q9s0pXDejglF40E1y3iCcVpPEAkrYh15XX8oxqQk1gJwW0hf
cvymPuURCiRrnYuZycbPu7w0oA/MEVO5N9znKqyiKBsZcqBrejPgj+WlBjaYV+KO
LoQDgLdkXwDxOgB+90oevxZUpilsw4xMSr3EOp3WdskmYpbVQNeIZkMFXsEOrVNC
t2BXpPahm/lDCL4CEFdRf+hTJQwLcIJAKhMV0a/vF0TUnqYLVKCXzskjcgzPxCAH
SxmDFf8rt5WGkXBEUVeIbItZng2oE+Ce5fRYJBHR/U/mSQlVpkjCBLyTOA/yF1JP
QZ3CCoGI6PeWT3SrGNCAmn6ffZ7sehTL88/cDLln6Qvgw8oHVEEn12nwGbiNvf+7
DzaaIw6mmYYgOpL5o6rWGoq800ZpEbb1bo3ttYO3QSf3P7nraS1oIcmKDHpome1I
y4MtBoPsCCHexgjfX9xajXxEO+azxNw9uIgDn97FjKvl6hljTqe3doqjJLpcc218
laspIzfHEnh+Tj/0G3pCVNcZAYMP3uabXY68HIaIs7w/Z00zKxCJrwWJuJqjA0XH
csqP8TiJwgZ6SfO1oIQZ38VOmU/loXPz5WtP4gdelLuTyEyL54MfC0ziY90Tgj7Y
gooWN5QGBbeL4CVHZZM+AD32ENDjGfT/yQi61cCujtLdn8nT7Vkxk+WHpuar6vH8
oBFcrDoo/egFeRjiUZe2WV85N0MHtHbovenwOmYROPQexJu0cz63yoBp6SrdM1ur
w59LixqJYiuPN8+utGqYLViVkT+pvR58qTzW/noSGCzSO9CVtkyJUAavjnfS6xTQ
BFotZqoBV9DOtc2PrmmKY6OKtgIlS991nrwwN76OIaebRMppqZE9Fo+XXfswQZ1h
rU4W+uVru7kOcM7hbsw8hSumjp2ZUjKAOvwiglVY6Cx9FkPrOPXgj36OrzgPr/9E
M9LPcLPQqrTqxZv7HtkIzBw6yX3UGObPX+gaRG+/zg8KdiK5yhRh+z0939iLDJQY
hTlNmJoalFDi4OrMsp50Nn/qinQHbr0KI1HdqqdTbpwR9pA4mYgdtI5JHVbTHcz2
1OvUOdUjQuUV1Jgtak7an1hrFPTrcm9BYV+p2H1kvSp/KzOkLIQcbGKn2kUFUl6z
I1y8FUlE7mipalEckDoL0qmAKinwkX7i5cDIU+m4CtL8EeXcW4PePUm4m6K8TpTY
p0Co98JY1bR/CnKIqX0yANNYhMOcAXq1cQfiz3fZde6aknzsFUA2WPGEQdkgKCAe
GVclyBh7BPi9hBUGRAwWH3j85XGVmsKyq6ERH/1Dfdd9vr/jUvDnn8fZx7kW3Ki+
ViBagpw8UdUnLZzUySPlCZv884SzIQqBgukD8KiJJEwV3qEAxaRB2lLxfv8c2dZm
taz6tOAsvasBwslV7fh2/LH5zSuVwW+u7quvxnyg2XwRyTvLA9pGyQzwrGnPIxUp
2IX1FQvEu82bbc6HNFHJnIGxW0I2UVsOtUaMbENQu7zikHyACD8MPzlb6RboHM2a
SFyxPyXtlS5UhSfo3Tj34jAhmPLHXOZeJQKZH+5ynqCFSHVXVlcEHs7Il6ISbfuF
IWAPknG1SC815i6UIP6cPL/LQdbFjNABaOsdaOx4NonoUdYA5Y9lemUd7IIZEZxQ
KeURdbncjbQGksRhkp2iRxiRk7xcsaOeV1nHfnZvLuY8SeHG1m8tU002vDsQe3tC
r8cX18s6b+ZIK310DuBMhuj2df8P0Wv3/DgstOs3ayOLnSaAztzgqHjwgTgVrpXp
z6m2e+pBdy10p8QO77SPVigYe2sf8ry3fwpC8tbAjgdDrjewiQBqunohcaJF/6/+
+c86syHkytdGkNO4i7Jn501QahhrG60398if3jMXVFbT4q+K3F9Ppitq+41mYhzT
xfmsEyXHBFEoYoWOqK4gDMcZZG6D94M4ez0AvSCfo2Peqb33kGGa3qwAfYbgY/xc
u6J4B/xk93nglC/5P3Ia7jQa44ewuW6ufhIKJ1s4zrmy3S+QDONpt6olP8msDp8O
LxehP62dOy3L0shKpgb7ZPJ8+/2GzXNc+xW7AMK5qd4KNJBgbTLoIbMpiVBZ8xbq
cMtpLjHCw6ZlKBYX7YSKlRB9k9SBpNJLfQfx3HiEVKTDXycVYtxJQTAnCmtajeIE
Nx5l2gRZ767KFTFzldiC5ZzFtvPGIxpsvgp+3TcD3veUUolvJp7vfKJSj6SBHBV+
M/pY84x4lHQysIBBD86fDUDITgjYpwOUemuMDcMFq625DB4GlF8wYmM07qCMF3Zt
up7i7hFR/nW38XFPvfVaj1IxOtc1mxZXiNEtsBq0S3/vMHRTZaYtOZux6Cw4wVmJ
r1OoAj121sBltz04dP70mKOXrN/voErnccz3zE5AQ84UHnW5Q1uFcYxxfM+XWJ2r
/ACObsTFjI+reO6xgGWAsQ==
`protect END_PROTECTED
