`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNE340D0+FyCP9dlYqjeJ6/iGi0CGgV1vI5m97ZMoLd3sKARl1aAJo+0pvh3I1O6
otYunstPShb3ESJ5XTCYGZOtvpkfetjmAXmcIl8yNVnOEk6y1ycjltaTk6h8VLPD
2PRREVTckbxCP0j3Fhw+zRoJwGpIP6kcKFod1kRrg9hZEbUxjFGWyrBK7cmMBAln
9TDoDDJ2saUNF5ruCXEETo8qotJLXZkFgCENaxW0aCMJ4ImnI+IHY+36xEpUxqn5
RAOuBZX2MpAJ3W2Nv/KD5LisdiqIoZ4ArnGBebtNPghtiB+qcoXr03i4j/HHpTMA
dgtj4050KmJj0Zwe/spUM9Bwp6O5oxJxkqfITBHTsqBMjj3sKoqDxQf1Fey43FXq
eLJcyHeaKg8sEoDql+1+446edw8v3puvWSWG+9Ih73E/xzoar56TLyO25L0Ovq6G
Y2nTDevicQUKGKjEOqQDG0JGLOFt0t5aAOPUHFOq+bU=
`protect END_PROTECTED
