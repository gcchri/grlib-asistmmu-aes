`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6djfTEKv1oQZfhFAGCMuX/kZuPryukCg5mQnwjEOlMsDOD09NUxnb4qaxjrFtBO
9ZclDCZPIatuJ71NClNlQSpind3maOtR969JRi/oBiHBiKfuVA1dJt8CqdfDEae6
NdhfJPtitcHLSAVjDRnOOi2MavHvGhTN18NG8ZzCwVn6PO7jGjyB0ojs7ZZsFjYU
45Bbt7Imk12WuN3OFD2+NLLcyOWEEH6AH04zUMtxvZKFD7dEXM69UXj8r2QUD56Q
JU8Em0tq/7rRxzeIydm7ziB08scZ3iLZzpZcurQFyJ3ojyspoectPVjItJgVLZjk
QjmYRTEf2AqTlqSDssnRDlYpB+16b7UO8NfEOm+7AH7jS4UEgPpAe/EgTlTo6AK1
G1Nhky9LKYne5oJHyQ92hcoJzbe4mt1/HdiWFm7fYqmKt/9mK1jtr8NzZE72X78u
+CEKoT5RIvefLtRb4UBQk4Qx6+GmimQxdYobGSF3Geg=
`protect END_PROTECTED
