`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SqSmswXtvRaES1fY5hg+ZQXrBarYXhq6SXrZCxoh2Jwbd4dBXHZyV9f1Iuxk5IAR
bOQLor9QsfmddlEbNTU5TihFqb/XxlgrzgynrIHA35Sh7Qi7PIkm5vQo1N4WY4U5
KoiPPVfspNGzb7ZBHBdZ29JQINKwRvH9w7qvFb9mSVqfz80Xo0bgm8KAm+Vga8Rh
QDiwHOXQwxXQnqBDLnvfB1OfSFG734qtpAjYCylq83PTctPEbPvx+tOKh1jH5Hxy
mvJ0SRi7gAB3GuU0WFQ4K/ly7BNe3CrOEQlvN3v5eenm89sV3IE/pO8GIAt0/Kk4
Wn519TVSK/u+/d3RlEVrXOIKsb55Sqru36MocvYlt/ef8M/JyMnNRNue9Ksan+Yq
4R9Lz9PDA6bCYLaSCFSNy3BWSQSftsDlRCYh/Gp4cY8hNeSWHuSjf1HMTv74A2bq
gNqNUl7ZwIFNLc1s3atT5IlNJzrGqT/wJ9g2vLO/JQYKwym+fZK88g2URYFo44EB
F5hUJfNpAx2ZrAjVDF7mbMfseiTdY6RnJxRUrxD+qegko5rMn+gX45Xc+7kUyPc+
TXgEOYiUWIxAvszPuD0t47plxjw9ILeYSFZa/0lKovO6tTKN2PWl6bZdZBU+mrT5
ykc7teLF1gherSrYccaw9wyQyh/hYF0HZ/Hb1Wh9GHrKK9DLxmVrXtuK3WV6TRJK
1Ito2E+kr6kYDJktLxQUO+zoc427+kiBtWSqoJT1AYj+O1cwZilYvutp9gYjHmcT
IYNEb0vO+2ifbbertFSdUOr1AFr4dqE20HKvYlNFlIsq+611POLZLSOrJ97JlPfQ
/+SILZE1ijCOnDc4FJuZ1TJiKLRGxJKN+A1yLVzUd4XvbxvgXljuGqxunmSNHRP4
A1SPF3GtrUwd3XM04RbRTkgMa7L3ccirNjJNVEoDQTBxL1zcrYY5LyQsi06TIagc
lSh5/bzK5Na1dEr6aJy3wWRi1ekY9FtiYIeiYkh0P984iNk5lFEJhGbeREUash40
dI6rT9b9PWNlRxqgPPbaChXKA37H2h8ECh5hCGgqQobsOrl6WzlVtz6ythMfsKd5
sF09pFqFd1Ttsu4bzK73JwZcJykYZNHYQmPhUXdQXZXBs6k0y/kqaLYu3BEJeYWo
6lzg1QU3afSq4fXEfRRBXjFI5cu2+PSCAO2Kcf+AFR+wQseEp/1kcG/EprdVz6MD
gu/UlcVJV2USd0CbkGDDheA/yu1CYE2hyGdC8whxD5jPuAPR0lsr/wwyIPNRE8ey
Wv2uKQPz6KOSOa3zrFxfe2xpvSJ9fGEDaD+TSKcRhsPgZ+k6enL/9Lzl3Kyi3Hjg
Y3+TbUzldc9vZNt6eg06nUPnG/yWnVfyNVeqMtsHsFS54n5m806Wq+9J3o0eXs3x
eWpWCrph3MJ1vHVH4sx9eHTvyzCYmmhH+/t7CnGMpx5k1IeNVh7T7q8mzg2+WVwb
wuBaIn9VsLoONETHe8gHb63Kva1syuglKydUwYDUoORQTAmFcnhjuEJ4PU5qEDvZ
SeZmg4SDKhvf2qSJZG/X4p17sNUxNRVhfjnO1VcUvMQtm2G46f1Tzuyn1s06dpNb
TFCg24XSPTyDcv7KWqgAe1/GgMMI6A/JKMs5NwH8OTQlOovoPbMOgyUp357UJ5Zp
dy5J7ZO391pU1guWrM8REgede9uCvkJEsXm//GoR6HIM5zD2As7JLu5y/CJAA77y
wMvb/qGeRadTUVKTPwnCmKXbvFhs0WL/ZgcDwM6P1YJwtmtmUOUSAZkGXUE+DAUq
lPGozx4MtPg5KIZTvO0Pctnr8TLiWJvwbKBSlxQllPeSnY8wfvT9/Ln56APRCkeo
j9lFbev1ZAhdeJ1++vY5r2rjAb3tbuDCo0k7oHjgcKdjD5bgAyUApKsJXuagQsAy
d/9vzSF3XUp4mCLxyXhRbbIUOkVcl0ami0M6u1moTmoKNEMhyAg2cH8vyZtUE16v
Be64Husj3t81f3ZEYaekmbGATvbf3Lt/u88AW2LedOIwBT9WjhBTbLzsr9nL9qTy
uzkYn013cZKSJBPifjeusntrLy/vbfn0UAHd4Iy/trx2QaUOLS2PRwzBV/4M0EP/
ntyCGjU+atpnRajRlF12RGnt8awNQL40VegdYD/kAKuEARvy2z5ZSVz7ZmREJ+Jk
qCq7p1Ndx3IwXh/gR6gP01BcOQAc4Vxzxp/EWGxACUHdMjlLbZEFTyNFk+ruUP/1
TgNZAgL+BgpX9z8dYd+04DZhPsKPHW0BG8+fctsuKaAnKCGzuODmVeloKowntYZ9
jWmqsW3Ej0SP/0lLfQPd1HKiJsMUzh2kj/HXX4vvRDKVK/iNg0p21tSmUp4airTV
66A0fs4rzahk1jxv/Of5Wj2gbfmyKkHuSI09E+6f7IlzH5lhhF1TYrntHreJSxdF
XwZz0flfZJY8cFa/0nWr4OnnYITJHe7hEZrY9o2u4U12cl0+mF74jQRrJLl9idz8
yQOqKmdeGmbhsM74qdNQojxUkMJig3gIf4hlFWvJFKcfpVci+ZXDzy078g79WODI
lACwNIsSdm699iUXdJN3WcxMDdQKKF0aYGyZstbd+bB6nGW7FSkfPagyN4+wWJ+z
IgZc1QtTCrF/TWu1ylFk4480RrOBe583/NE4LX8CsvnvH9GBxhc83vETxbShqpQI
S2mzHn4bxXmTbxqPMJgXOsKOpqPexNKwp8w93flRRO8rbveOQsYgtZLhYHiYvGcx
Lrv1bmbqDCSgUq427cAj7iH78F0dw5+FgxYSNIVLG0zvYlr9BRP9LdSXLCsY388J
oZ9vPhkup5ldM1ucGvM7Rxs9BCOkHKRiYjVhImJXfvvpCWvusQph6h3q/NPy1CUH
kLLz1lSIv7Xrd2F3Mn4WD2+3bRaNG9jHV1Y3S4Je0FEqWHfmxilxM/eW87dAnhnf
QFWKeYx/beWnUIbe/eXpnasaPzGMEbRlaOMfWjpNd2rUU75G14XF6JgvzS/2mrIx
Pu+D4Zr6VgeIPbVsPac2n3d8hU9fUzu/pGG17U/cSYMT2BImA2P0s9COJAc22cJu
b1MiVHP4077zmZRVlNmLWsByyVbcJtb8HKJ47FIqS7fjxpBH2ObxHSr8u1KaRwhw
73LklGhixiR6Enxdgp1RFR6q6O9Q4OEzm87vqgZRJMgdKLmHxiEQU5a6iGObvCIV
hqnOSKKbZ6dvqflhz/gJQa+SY7dC8abyqlCrXEfrokbwLXjc6hon1n3ROTuepFFa
JcWA5LRSCMj1F1b2iREOJhcr6iFsQDnwZkBmUE3qK94lYYyKpeWTMcl039jETsaq
ahJMyGe+u/3ZU3VYauXizSxLNm73IxNSvqXujrd9jZ+EziiScPTKKqZF+1dAfFfI
edwNIZxBME+bcc+9IM7Xa1EU1A1ItHYvhv2IWBntB+wxYj7lUQXPlYhRIhulYz69
AMaICUYsSZ9iZPPVb8jjFGRd+ciXm3O0MPWkAHGoRsdTHCo0TZSb5aV7kxdRMRRc
3wrLbHB8+FVGPmMPy4B/uupHTI2j1ssVauIxcFM/1U1EMZLb7ATUHRMmcWvf6JPp
T4nelaTFYO8qDrnebAKuT9Bhv/zvpChdqDh1qNYXByoQR9z0SMXIFePWvpEYoc5g
TNdIz9s71DlycsOCRi07R+OgSuCblujuTEFP5XASsydL9uB5tvseqkhVDhNX6euf
vS7woaB1DmJE3J0l61gyaBDQMX39ofo41YdfsxwPx3jUivDWOoxB1qMVS1+rB+D5
Pz5WxBVaYKj/YFMDRXGIYvp+QE91Zzrp4JedIuVnzJn4oRFeBtsiR2fgLXOawzsb
ZsciKgJwtrAZwuVVt7PjPS+jEKSMEyvgVOW+J/ubbW0kZ3vhToh6+sIVj1f1Sz5v
Yo581D8fDW7eeTSI4HaOYx5lTBgjn1DJcylQczQIpLrrmLqvrE+MPV5nDv+ueB8Z
UYAws0jsXBruBKzfCl5I391fSz50jHr7DXagbIutUxv7g2xrG0eHHakywuz7Dmz4
k6LiS2RN7Cb59NIRYL8GcNUeqiQoEXgQGKc193qQr6qAHrYDgDN2UKgWm0PN/3oi
Y0FRFJNmwWxFL6tWnplqpnBqA4B9AuO0U5XmqqaVNPZK52AM5npBWeCl01fk73os
ZlsnY47DsvZwJLHZHyi9DOYjCviu1Dx8FphYsPbGqKZmnZi1TWXRhvA0ouWsX1Mp
NbMSmHON3vwJjTz9QplIeEHF3+sEsyfeW5I+H+mykq3wIvzqAY7EPCA3/NAj3dFF
k0eXWgmAbN9JOUMPlxC92+r7yrzDh0tW2Huc9Vbshm6sDkKX6uxTIi4KJQ/ZTdeF
oJ2Wi4S4vRBHZ1vh5u+De8be1CwmL/8GoCyJq3UW0CoOYk5OLXns5Over3BxvIEM
oFFloh/rzJksAec4jH0ZmuCIecSOiQefaAC6WDyTW5wX4mVgMgCJCUYLig5IxELd
4TZ8mMxOz4kpMWVE/fpb+E64zDW+flMymq+5DiFwxvBTjTXaUWbuXJl5VsTyMWMX
Roc8XJRQ+KR0XJAAVgei0PtT3qzyOYVRRrEVZSNz77BMACpWu/lFiBJAFz/D2Wox
ymztCX4l1AoRR4HfKMOmPhbxjpC5ih+nzfvNNyzuBZX4XXb4SeSQA0HjUBZwKvhq
avaKzquwQ7xSsuZjPEtmZSs8cE0rzdyzP43qFmO6qqi5230sJDFa+xMHZ8yX3erO
veXWIoj0xXmbDuNoUMCLYRhGqv+cOaZtAWxB3nNkH7SbOVtrUn61/jjvVWbHAC8i
hqIOGMj75SB2g3Rr0NNahpsJHdydUnQm5SDuO9HyEELL+ASk55s3FDBFqZ5Ai//Z
5LOwQarqtoclxF/LtVOWfzl97diEPJxF29yF6kjTC3BOXms2H6qmOeCsyAzYN62N
HWRa/BckWlaWsNUmAK6agdYEFJ9OQY3PKq6Zctfc2+tO5ke18LI886i1dCrPeuQ1
H7SZPo6Cxl3VoAL4G/TmUj1+siCHun+K6SbCGgfvdLoaribxQuGiYehBbMKWh8IU
XByWtXXmbWeHBSYl6oQa8jElgWlQlzxriyVG1gLU/kkwnh5WK81uWj74q0mEus60
Un4A6SCoZyr11e6NqU9f0LvK7mYWTx/uJjRTzCdl++YptR6eab/eqbvnVr8KL7z+
KPzVeRfNscY5tJCP8baNSY7vL4eTfkkEY9ehmVVYm6/y9WRVBlzvxYSQBEj/7aRi
p+Yug7u8Uk0mkMCjOnkOKB97JWk03bXnNvtTtY/zfzWrZEz8SERKW0PhmBqA4wTl
MAQQhNMKdBilnGZLs8BL8IE+Z4GQUTVeMGJw+kwn9k3B1cv6uFkZFQc+48lfzkiT
iyEPEFIPL6pK+ax8UT2NZOg7szmoqV+WWLtDPlG4tq+fiYk0jbw2FMhuNMwfyPAY
Yr7DO9Nr87jrb8noqrKK8td4GJX73BUYu+tR8s6urn3x4s4LIJFfuF2mZZLsOWVV
WI/mTU5+eU4upFJX0Z2ZUMAUaGeQn2kiyZy+wtNEmhkelIBb8Fh4sSEYuWk1gCpX
6h9UnaNvZ0S8jPaFZwMbPuXsIavWTde/Ol816zQAz0nSCJrDg7x6659EZoiFA8jE
UQd3a1g5uXvtIWkXG0G4bAI4AxzW0q3k9ae45f99Rikx7cvw4eRyRxIvAuVMbJN/
+WQQvTZy4AKoXbnSRUJyWeUnj3XZaTb6j500oP9YOPZqS+ZWRqzyn9HTMXDR0Liz
Lb26Hak53vnywvAhNBYmUM1CAib/nDrBmANux8ePzeLUcHAgdlyK4pcNHT5lbWoh
kAibUXEi06LLiykcQulcST/B50iqPORizTIjiO8Onz19Fwds8yJkwhPKTXWhtLQ1
cMVx/4Oprm8nZcve0PbSR/nj5VjsLI1OqZNDE15iGtw3s9+pwvIMks/yJRTAZldI
S0D3BXup1K80+0CNsO1wieDc78IJVwcCGa3LfuaEwX8BAIAYkNoY/IZT7DJWxnZn
jFtwb80t+PGNQIRsI/QfefMtA+sb4ysiVjsY0812jH4ncJ1/WJse3zB6j71J/J0g
5besFkXZiz2/IcXy9z8oT5YSCZmCqzwZorxvaRDpfSX5tv9kTtojbOuR62PCaZJ2
Z70owit04y5amiV2scoC3kDHBeE7NA2QX9stgHuLZOGf5wI+n4dVMHUXTWPUtCtw
A8jPZR4q+CseLFyaPFvgHPvgSnSkni7t2wZdyj6xxdH64Z01AlOb7hK4cI8krVMz
QG5K8FjXxxZjnewTf4791l4hbeKwSLKvgf4hzw82nqaqgxA5JUdcMgoh+5dD7sGU
Z/qtlB406mmCSlux+RSVczg9p+TxMtKM2Q5tZPsLi6ajYpWU+GmkyYYZBBBXriQP
UBS1G/hQYOOhy1LuIYlcoJYVuULDnTKEAAF1u0Tdc/RvGouqXl8m80EaZZqUVv4D
bbn4N8GRI7fTyw913bAsY//Sw4HZpQKmTXLU7ZPx9d/hekGS3/+RdDSD2Vhi483u
cgSOGIob/ky+PjfTRW/H8ryfYG+i/a8enE/ACzKLymle05HI8XesF6YN4u0HUUCc
rOZV+BkIzsDsF0rUqjRi21SBpPKAPT6/HogoXJ1XMD3bif/KtfPx2V6JERn9y0NG
kjRkeDRWh6i5za0T1VILPOZoenvITqaOJQ7MYpiOtPKbLxm1wehJIrIzxdb/xjUl
AWmHpDHkQ0PLDQtAhR8ScEdrhA/F7HPoRW5QWsj0D9xgTtCJCYzpC9NODRKJdDor
0zlQETKy2/MgFaeoYV5GcC4LO/eVPHplHh9r6KV8DbUI/tvNcEloNNqheANC1VWx
Kf8nVfC0YU2E+Cqwgf7ZuY+yPjndKN7s9VaZ8N0tze5/cdkSxmhKFqqN1YaoejIC
t+d1KJ+1m5AbzptpaYD6HSZ/iNib9SiFzdDkkd2Yqmqgoh8UojSyyjEaU08Qd/mT
hde7GyEChcVOLCfVNO17IRvwCcpW6U4ItR5DHUjwUUr5p0yKpmEsevNx3FuayNzn
Jnbjn1jjFVWbXCgnPe1TVNEUt20Fb0YkXRhl6C4slb0ep8s8SpnxU5K8bt1iod8F
4BGg+Nuk3LhNuKF30ven94fLqGNqo23FvoQ2dOQ3a88Lk6W9CsEE81aBSHZ+oSBD
aSJ6+NyWCeKxwZ14f8cp4S92E+by5jj1P5MRQV6DC7r5cc+XKK7CwmldKhOsErWo
cV0OhjgwBdjI1MalvIE8Ie4EHK8KGXzuZvyXxdn+O4U5r0K1hBWHHF/EvJTGJtXM
BVvkpUWcVc2a6Pfi/rpUel0C2dKAaH6hAw5n3Gt0QM4f2F2bf9OdiFkknH1AJKof
9VJIC2KkJD4gsO2KiBeryYqHceVB/cf6MMWKrw9ChsKScPMSqkYM2ulrjxLBc2iO
wFFHJCltIvBD+9BQAvvGjeexeVBgTYyLRDnkoDPelPXHklAcQJR8Xkzqnifo8hFF
ji2SuvEr/ioBKiBsnXfIfVeeXWRu5C5S4dGFeWlR0J69eOHfeM7+frvHQq5SYFdj
7EwogLt4mw2weqVrvCXpXSWY52cjzydRKV6LQECGHdIODD7LQzT78pfndFcO+U1U
iA2/uutNrrh6vccqEwNrms7LpOnvHVSVJWgsvfu3Bdiep1Vs92N/D/p18Kkmnbpx
+SE+n6R+o20UyrQ+KTPoTTHIpq3+nsWqOyNLpeiCXuk1pJsqmKx/J0PsnL/rOEtD
9h+0XNBoCo3n+XKXs3A1liVpAA3U70eQrz9EIgLrXCh+WqHYCA2XqPnHgN+dBaC9
QiLYvHm87oTx2g4nRQA+jN76WwfpEdNRERzTHzsV9KB6vGeJSUq+7sEXxc6uvKrw
F6hCTZwZSTp2LHtItr5jGegzKTlJyZwBRlOMAmZ7dUbyRLMekVm99imYTphWYkD7
vT0yNwHErlQyw1wfzOlZ0jwcNlC/tChbCo6ITg8YBFacW2oY8kwU1131fcO409oa
0xMs/dBrfGs2u4HjjJTBxZuKFOMg/489IPrTqtmQaygF2FTW2DOPn958WYU6MA5x
jAuhvdOivGrrBnENiC6Ij6F7kn2jGcadF3kP2XsSq8eZb+pFB1sB4Qt9D/tXb0yl
t6iDcHMKc0T0/6kxKnbOurwwfd4TSxIPiLywf2iVmb3O7jW70oOYYGqXoWwZFu+M
VkmavXF8oPRLGUY3ZH+o3YRFCQz0s790dvz8eMbWeqkONqIUf+GJz8YZVUHAvZyW
VoPACPdhEeHYXPAQ9/sScHu+O9BfyXt7pxrHDDaEQNafkxh4nyhulmenSZtDPD9Q
wNemkavqca706jfuxS1PW+5L8sm4cmcWLaoCD0Ru/cpdFjre+M/R8p4e5y5UB+wr
k0k6wD2NU6FYN8JhvVT9mEYOTHW4olVvTquTgQwfESUrg/rTu5IFyPA+6kD/+SzT
a9xaiRFK+deRxpAClDCRKUgHpYsmG/jfeBmvLpI4lesIr3I+WA/ZUrNmEphjcVya
sgSiaPWdlcA2MlFwpGD2ikwT9Zr/nKnZiYXNQHV34oqi1bID2NOpY1EUXSn3pv3t
OZojlqQI0A/2KIj7fVU/W6tUmH4ioygx4eXlZU0kdx1+9OsuwxLhFmgh4de+9sBj
MSELmHmOXBMns+QX1bRkZda2dqYIUifaNcvyFhWHdEvpyaL8hXxIh4dYPPQi3NI6
NrJr3AsyPOHuvoP5elfo7rPwryO6VAZbigU6IdYZYhVAADEpQckcc1IejkilPEcA
vH5d4IZpsR3N5Y7CKa6yVgRGkHJpaSPHfEmB3lQ2ALu08lfiI8XuDiMSdPyxS8WY
Xdhygr6F7/4QuzCIdNpCZex3qyKnXJGzY0gu9AB7osMAEqj8udq0Q8u6ZZ+zYpwH
9MWioEtuljGRdl8PnWQNoAdT/NHmU/5pTOGzRPOpLrivELNH5FvjDNC0JO0Pz+Vp
G02AwS4WByZbEANOMm5PC9FVPtk6YqI+E4NId3DRwMe3kSA4/67LRpmO6nj99UNx
cUDMLBMZVf+OJD5vmpUkN+bU8YL3k1CKnc0V77jI8nDkJDX3891EfaL8EwbIRM3M
B+llpjLCfaNxIzGMh+G1MZlge6xNJm+12HXyU1H77hwAv9/cjosZob27bj6KQnUZ
55HEM9uEPTD1isQ+PzVacvWGehSuR8PNAzdhCSEPbE3NsHkwlEqgV7dL03SwIPI+
QUmAEicl6Pju7RyjWSCHoo23KHFYMOTFd4vmZ8swtQhwhCTcbrXWEdKNT+wDAuWf
kli+0rMAAlpPQSS6QkPAAPtkLcfmE3qFOj6YQlbELf2z5k1nEwAYOfqwAliGr8BB
LtQD6zGEWdPLqZMf17NNkECufDXYpHuqqndp+TguIBYJxkwtxlYM7qkZxpOiLdpv
77vXW5WYslUXlDJJjn3jOLaDh6N1ZZR66w8vBd1bwqz9K0FlU87sXLW3FmhvBZJ4
+zC0mQ2P4JGvB79ZGsanaLI0M3UXR5MiguI2FR2Q4E48iAqXqNg/jTEd31MCJUGy
7oskVRbyRM2aGAEEB5FTZiK4ObZpNsi0yD5USVr9KZVtsQkcogpUT1OpQMe8/Kkn
5rWFx2ONQgBio+vMuJT8spzZA/t3K8ddUv/R/nsxBfbscOOJg5eDZOpytfamnZX1
/k3vJoeVK3YYF0awH8XnljDNYlzEkNwYOWhCH8fwhejWTm/m2qiTjcZU4gNBSRhq
/d0rY3Y60WwfvUSSRGY2+i2ZJ2HTBUfMWjCB315AiJTlZNn3KCBUQDTpQG8Lalt8
vC6jlRnbcFmqU7FpoXKX/GbZuhbo6vN7Tm0/ra4nE0UHo4OvnL17stOtreJ01K5x
uXLBxpsFMFbT9mCrzUl4qMmnXx2I3r5e5txP0FdMEujlsn6KtdoJu5Y/jQj5numQ
FXj6K5H7CZFtQLvjX8inDnu8jqnhkCt3angRfYfbNg62zfXIoc5EFOnqEzc9O/Tc
vJlHxK937a9WwKSuur+ZmAfnZeyhWFU3rZmwKMpY0nrTDcLAwUGj5SKvQDSFnInZ
AbyVP5i45PqACP0BSIXydsFL3gHwABXB26RIL7gYEnwYvJszs2+Zjoqv7dq9wyO6
FtcphBGvZyxIyCE05ZS2ndMSauIUUIrKmXzjLCxqW92jgWlgAvwWOveyY2QmUJqa
mN5M6G1D6aUQXgwxQr/FC7EVgoDixtbUWhww0DLvL3qDaiIUAMKzldXART7PEshJ
1gYxfyn/tuFb3rPaCekihx9TSP9nKQ83MjW+79BFv6mtuPAdmgHtnSlH0gmvs+Uy
uALmJNzdJnyY13+hjl6CyJsPLGKeKqY4/JP5YelaKc+aJQWcNaOzOsAbdMxXnehv
Uuk+MdLLRaUnOxQorm5A3EARprLtvUdHcexROQZG5EI0wGsAAFFY3Zf38OIcznHo
SbWG+AMo9NSAyC2qfMr3Ib+e+/Lr8yohU2aeBi/7y17oCqyi5vBh1Z0Nd3aP0Cxq
LCUlFq9aQP1ZvXRgN/YYiScwFW4XJTNHHHOg0f4VlMfWte04+Rl5sN9gPggI7SSq
ElWgqJek5JmxYeKSs/PNqpFev18h8tiSpjt1McyLY1MXiMonJEfykbPNRueLa+qj
CwzMw+izAjz3VNL0m4hvjyw9KOc1jX2u3GVavQ7kCYnZUUx48M64q3ysyy8mEL26
qZMrU8wzDc2Yv7ojSe2vbwjm9k5GAij9+L6ARXXCvULfdV4PdwRay75DlkJ6v8OP
Ev9aoSotsxeB5UB6+wockOmjulQIluVJPIOeg1VTgffRsLvZrb3ybJkmklhr/kzY
smRISIsdxbEMqZAKRikEkDqO5TxtAzQ//kyAqhsDNFGfL5/R/0i/TB7ltgN0qKzk
tfP6OhXqJyUJytVT+1P+bzcXSTsA3itcPxDTtS3maudcubV7lSLa+OErxcNb0cgo
03ItpM1Yb0ii9AnQfVQJjQ==
`protect END_PROTECTED
