`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1FvaDszYFmwahY53Z5/LqO+elmZNvxm9nVQ+g+yiP9j/H6IpKv+zlUONlhq95xzS
1V5EWeRK8NoIuVgJc8cCeb4c0s/mNDuj2FjEvB+/zD4zMhwbgw6wctYYIX8hdIQq
5G88GoZ91D+fjuKZ6gihwbkvkKDiLU3N/weiZxjf1BQXqaArhXNg0pTIXsC0+T/2
qVEtFCqPKdBNrnefypdo3w6EwJwlPMTyshJLivMaTRCzLaM1L5S3oYwQO9/k6Qlx
ld9Fh5htxzgF7HiRKDb9udA5Dp5rnNLrMgyFSU/SC9jVlnO7UdFeIATluiAy1aEJ
JBRxcGvdfsykccbGU79skSbgFkcgHTbhLCdDT1+RNs6aikA/XiqdjLRrUHCO9/SL
vvbB2+zVjLk8BRtXWcswW6+liWPFB8H/Gt6hWf3oXnvGOdPozZgIiqHfkSAgjgnf
o/tU5k88moGuFxGD7vdT0hyv/ep5hMFX3iYZku16cJpLjb0OW7qm1kk01PnLGhdZ
bDW6eLnt2RpdJoqqLWH74qZkG8XZjcyVoWRV74ril3UrqjMZYH4yyfCXve9UmSfz
g78Kz2jbdVmsT5cn655/yqbr9SF5uOXYPmVGtwVpa3ZoYf4i1+x975qqQoGietWe
VQjAJpO6M4010KTdD2dOll0K6UpfpC9/R+EwdfvFtZmnuGsJyJWHzKrFEyQYdEba
I0euRj2vKbwx98eYBNncJr5m4S1g3z+5UXNlgXu2BEVgOmTaUJlEqIrTcwSXELtB
s3Nzs4l/JmpI6We61FzSI1mFziDk/8PSN2+P/Go8hTyU2PEwPzswV8DbRa1feLUC
mVz6N2I2fnDdIVgoKC0OWW4+1ZG14eUhlKdunKswpLYwOtrJqK2vjW8UUAA6FT3o
vfSRihL8sQXdokpRE5lPhY+p0AyGnebd22Wn5In4BqXonrkgIoAd7E5sjJQ8GsEB
jfz84U84xygJq+8oT8kco/J/K5UYZ/VVLNFUuWrTSZbhm5vmMYsdxA2f1Q9D5jlu
PI2Tl3O0yUUQxBvHiGXbyfRJHlkd5CGtWOU9gNYW4uYKrebTdTZmR7iFDXOmcnQs
aRITCmC2eWVwVvj/rooz4UMPrjgdwC2V9H9UEylcXXqvMGiryP+XzeTg3vYzhqHB
8xBRcqAk/dBvwxZ73OWE1X6bqCWJAYlCLLFIM8sRSmWrx24RWZhKRVoYPXY2370t
8xKRKg9RSw+CqFP6wIqMYmvBuCyfYZ71Yw6CS8aGmKRhsuPtSCFC82qTR13lSpeU
93Z0M85wmrIXKX1vqLM9WTfbTOPjIikEeoMn1DtLPxCUPx2eFnahFE30gi/SmNF+
Jh10Qo/HekooOEy/9ksKV80LxyMvTdk2lSfh5e8sxOqX0Pabrf/qrcgYqvzFACeU
SWzpgP/Dm+1ATBaIWPkw+cLACkUSBu3Y9uLS/lLfFaPdfwYU+dUrxj8wlMzmyg/1
lvw7+fz7B/t4ZgeRRWfxtgISJTrmvUwXF4/6CWRgWrKV1TY+UfQ2LmIz+zzzkA+y
Me4syETLYS36lw00OsiB0nnz5qVjKJaZWh1GRFQYGk1OMCWuJk2eIvCI4raZpwqk
lx8gfYNDUEzP3ACfuUbWv7Mp8A8M/99EtRB2qQdHTclsD3J9JL+5e8xEXdskCHqp
6vuGOwpU+MMD81geJySZUT/hg9Q9akHXoa3Ga3/yrPX7XKMsDdb6IVf+AhzdRp3j
LtiXc6urr0lpqmgvwyl22vkeaMMSFfTDbRzx0NguKmkfsT9QgB/cQ5rdgsSc3Cm4
p3T1365A3qpK8Gj6z74wyEKNWBrYmEws+5I17YPWdas8GAsPHRvhrWDRhAURpQf5
pYt7+HkMrObLMh5qLnv8rg==
`protect END_PROTECTED
