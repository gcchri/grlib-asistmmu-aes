`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aU9uZZ9mkVR7zTK12gtSjNVX7oRMpG9qPYCQgAAKdV/hbrsJiPz+44FP2E9Ugvqz
x4tR0WkZoPXYw4L1zcYf2wSHLGXcn35zbwhlJT7r3lNID+AY48kq+5uVmH2yLbYS
N3XukNCmZJCqwgE1QDQc1BMl4yXrhigRKDjZoaX0/6eqeI5MTfyB4gErWAZIXAM6
8qfq26m96HKVAY5cIoMNiyYtaX+p4Y1ZW8dL1rFtWrgW6wpy/rW66vZeAeiahfye
7snwvwBzQZ9zHbo92XGOl30mBhx+ODtLyAVzEhOcfxZ1EHeFYCU/0tpLTjvvby2K
/KPdHYg5gfUCWsphZUzlaKFFwbnAqZixxRkF7bgRkIScXrS8ndkGcNv9v+oYL58M
RtZiII1a2G6oh1ZssMzkbFKRYLmU0/uiCDfWZuE7PqDihrL0RtT7QKay27Ogm8Oi
VZuuibNO3SynIBZtr8bP2PSRKhVCOZTQvsuUsh/ON1iVI4esriknReayb5YNP45F
toLrWRim51NOjss8x3SHbHdrLm24nITrkc0iIQWa13fapnLVngPqC7frFEDCYih+
o3kzzcFdr3/kKZ492oFMGuFzexmT2p52LRrHx4MjFJYftXM3/hRcz6Z/xhvaAIZ0
c4m5YigoIBfCtwFyqHdNwEOHHkFiAOUQM5uYnZZNdJnZqG/GMgS8mxX7mJ8/bsJi
tVOljxy8XGC9W0Tdl5f08rjgoDFGpfDPxKV68ssD69AeFxQ2OcRM32MO/9ghncHy
XFSQz4sfuHYoPt3A+fWt7GoWgOsK+cmqcDHdq2GOpDdxhoApUGRHX4dXJGJ+/jB0
frnktg/9xteIiy+MU7mi2Ho+HhJAx51Rill4MiYV2dxvZFfANDOXSvTXPs99OnQ8
ff6W03t43h+8fjHlLIeetiyR7xgQX1k2UgmcVyaXdy53bkCzehoyZPX4AsaCjKjJ
dGtnqPGTS1t+jAxoJqFSeHEcH5zbd67MvGsrK9/D4OkrQ5aqD06vvB11/zduLW4d
m4bnx0NEQNDWhRAvQfJm8E95zGkYFSbBPDNIY79tNdB4xhZE8bLC5XIxDh+G1BsI
K8pO6IU6fYPDkNfzizVcnbhuadv4c7QuctfekopByjKlRVmmvHfkIncxjNK39gl8
J8l7U7sU2Q//6pV2g+pzS+Kewk2ZH/Wk0gBZKBBhiZIvXwf/+23ZCrVOgGcsnJDh
en8/nm/xCi9iY5bd6I0RrUp7ebZwvkdEr1T5v0zqDxF/o6YeKyXrExBdCbJrSrX8
VltXD+68LTDcsahkG76qx1RgIkeOvElR5UtgtKPmXYBILMOar4OdrEHuTewImG3S
EXBc/3Ihg8LX8B7PtH4SkdmuwPU3Y3A7F05Z6kemlZ/ssVzjY6VHGkxJJAABcO3T
IjsMYNfAxoWZwnjStVKWQoABC0CWvDAUzSwRUNKWSN/k7CPzd/g29mxlbzuOqELm
F9UbYu8+PruVbBBFQrgYO1+JaOKwwVjHASAgu/qNBWiigtpMklM4eN06pIYmtX7P
iUokoR1Pe20Rxd9PzZD1Rj11gOioaOX6h58YNTP5v5CBh6+b4V1Gc9vNBu0kMPNT
fA0813a6R3qLdwxuT8NMxhPupqWLLoRC6YML5lAYRcMH8XvZ6p2lALDmEVsCeWsR
WMdGVT/TJkYNN+HLAKwxYa1CskHFbOPd8mUS39JQmJwfO90Ca0Y6VU6yKijawGn9
dQegncSdZw9m8VIejYwvUVb1ikzApH8C3wxgQJVsnDVmuFIlrusbi//66CXoPwjm
zXwk2ckw3DFjkrUks59HJncvN39clj8FfgAwwn4Gc4LsTvhzTQzh7geUpa25z9p+
ori4D3yX+JGVAzAyCQvvuo6sN7R6/qmaSXkU9CdejikFSl/mG8OmB62Adr+pqqyh
UIV4Fn4wUkMSmaDaVESpmzLGj6W5ZjyYQU64MjgnRLIo9g/SWLDNh6KvlyjvmGKg
S7qCowLSyEGOBbNDcI7P2Jc/nOn9SURhHQDyuy399y6OCuYEN9fJjkFFdq31lcyf
fGdCzCMurOz03fvG1I7lD7ab0bJV0qbKGuJg2sI9vcVKDTsacwtfqrgmpM82Ao2Y
vA1iXBGrYMGxxAYyS/7V1rfR3/pw7AyzpbO3Kla2cLecihScVjBZ/1T/P319aqEK
q2hSUokjuapz3h1eK8bXl2C1isee5M4kJ4RA/LYH0fczkW9StPpIMM18I5kZPeCa
uOv0dIVPuZgYdXNxhKtkFIOIDVsW+iR19ARqe9P80lieps37vWZT2HcoRAH8TE0Y
C+DKkKOCaNDHGy6bKJU0iqYypSCjUeoit9N/bnL3FSgzB7qbJBSxUi1xIBMxCLnF
8GnVc1oppleT0+G+lEHY3uzJDYB90Z/NtoIyErqVs6+cEpsQpFSwfSaE0q2wUsy6
XXVx9ZoucWHqb+1TAryYXaJhC3k5QM/MPiYDG1vrDaxISQE8YwJ/XeQt7Zy8f7ph
pK5HquG457wjH9C27827ailyF6XW3LSJdYFm9fzJPcjzkwSbz00GAdppF4oX3ji8
yiHrI62M4P3tHublj0RA6DpBITh179SgtHqhyqqfErcT5egt1FXmUlavZ8BL7yvh
hvKpJj9ob2iVkdSORUz/quEAOc5qsntjxCC277nQUP3ul8SBMf2EoBX3OvutgzBy
GPHW9EWJAQajDWLixymGopZTBtGEI/SAMzuCNP7n/COL+JugA6CbCFUs9jnE2tBx
Or+TlvzOWOJrRW2bt2B4RHIqtoDa7AX94Wt5JTMMfjAOYVKQfeXo3bB/yvwH0qoZ
9Ul3q31yEz85d9IZCIuaEGdzbKCb8prM3Ljgm8eGiMUtLkNAGXTeevN8wyFjeSPX
SaIy1uRg6fiY47HX1TVmgH4hfwTkeCUmERkuVgG5kbx8j81yFeFdWkOK85qDgiUE
NboSTlK4uPwtd8CSv18CCtxiBUPhoVLHHRic0Pg0ZqIOLElYIhuOZ/VbB0EV0vWC
CQNiivml7AlRpbu2S0T6gpzHIDPIcms+KwXqqsldp1vj2DYxn2UE1k5tWZtOBbPM
tQcnP4UPDC8ILMkAXjHRkIapNimWLJxo+XH3euwiFzkeFqlNLdvA5RC/GaN4NV1n
g4wMeGRz69Zcgj4aqOdRdDyN4U45XhT6ZDRkh3nM2Hhfw+W6uV+75g/fE5unxIro
I1ZmoxKT/42zKnWWiefXWnprfxpWr2LaXNJrMHtbHe0NbGXlYEFypurlmTerCyn1
wcBWvHFG3ym2RXeZjeoXOhuJ1RmTLD/VoUlMm1eOv2o8oM3522Z78ag8L0w+M7mD
Uoj+tswXtWycldNF9y/7RiSE1t5//OoMl1ge/zI70ARnAippG2cUq95FpXDgNfWV
lxVaOB0uGs6tpvcVuWVZjFP2dqUAl+oBua7Fr9wwVqybIaWYYDCpVk9nz+zn52fd
yujNPl791TlAmLRsSa5f86KjKbOO+cMttxDXrdjacymkkAavf6IjlYmmouGSzSBB
9dQOK+r7vz977q3Xk3fsdbC+WBQCBCAFoJ2TmQURN8ODFlxDlXl88ZVLF2AxmxT7
dbM7lmbhHkryOGZDHgthxvowmg68NNeNgHi9Z5fjZgh7FDHEXy3FxBOyBIH2UhXB
aCIOM+U2Mdi4sodGx1fE0cOyONYO+eKmdBzxsRFeUlwXaWH+Nh8tphBl0YqTMy4b
ABgqIV1EQuxUvH00VhmN7Epqo4ePRWJyle/8wPpcsEbfxBUWror9Zcshw4FyKHMQ
2dI75iVK96Jc2nX/Sx/6WkmmdNI2ROkrAGt8cEZq8eZHGaUF9sczz/7VIMitlVLa
cWY16bAOIoDewBkF2qpm90IybqM0GETvbJKywpPx+yQmjHN8K9Twhc7IczF80lN2
VlYuwbWj9tG4i7GMTHVSEl9lKoZV6oUSa56E9oryMKPcqRGC6B/ncK6gaVk3LZzG
uNXnrTlp6pD9u903UKRdRNBBAkZu4hdxTkfNlZY4IeoQwLAGbwSU9Wuy903iiJR9
Hcy17S9S+EzJZXN5i5n6gd6n8jFi9ilS3yP3k8g9wDLk6TkIdj6kUsJmDOpmlP+M
bBu+F+d2qBo56XqHSbqlROfSy9TZRC5ZPI1nWl7D2WdX6+v3wLFIckOHVP0jAkjt
iyDWPIUe34E88wmS8JS6OUm1lJB4wLOtZT2rjRG/jJ7cexCYD3mM3SEXfhM9DZI1
3fAre8jZQiEmoKP3qXFCIG6QluhGbXSggYWBBrcC0Sfa+jAxYwI0uINxsTsxs9+k
VmUKWS4n+zg1qd8VUGZfb2yLEoZ16Jk1MM7M10n0y5tAY1Vq2THA98hUSnfBH+L9
aUPSk5vN3O4ONqaSaTeyOZ4HTXID79y3590Pmm0f3x2p8QYo3QNbX+TqXBN/TmNf
IIWT9sFQW1E6mO/JMV3e+dZrp5bEnEp4npW6LrH5ZTJdUik02UH79JPlYBolcNzA
04GidBDbrQpq0Pyk4rniRda8Yrec0Qkpou1O1U/JCtBIYLdaZBwD2WJHzzFdyKuh
i2IEQhNZspEV+BkIv8mJBw4CyNh6Ngfh/lzv/81YXwvXcSLJa3qk9582Tb23faI8
+9oqRX0a+vHjXL4ui5ND/Y+HNA01HHZaxupwajPkD+iUpxCNBOAOoWRk4mIj2phM
mwVEf4maPYUrn1RcN7V64ppsqbAhPd6csscwkvEenEukJU5N9Zwp98sJc/vsE+Vh
xENWWUzGJzTOByTQQOjedwugAjOXhASMf7CHSlGt7GV83YIz8QWMHNOMwXcmbqMe
x+abjmrgLzLyzy54HyOyOTRO5hIBwhlj/2iHSNl2/cj1bfreRfLYgLOcJ3imF753
aCK/Gtb1RDaGoLotc5jgFNSdiJ4YkNzWfRhetWtBmWcfmBOQ2dWr4/c/JiimR+Rj
tX3n0e6SEn5onl4+1M3LLirDnkIPk1bHVJr4kONsd41cZGuNR1sYklgQ4mXr+3PD
ETuJWYqKU01sMA/vZyjVYnsFNpXNLFMKP85ukg2SOppNJ4izLNjPEaasBeuE4c0q
xYnP0Wa4NerS8rwzH65im5eimvWvq/V9aXYnYZXAg3VG5BE0GePtTY9gc3qeCnHd
pkAhsWKCgn+/DwEZ8ZSS9vtqbyZLTm1ZpiJ0//tQMNnhy1ARpWzz6EGWknor2Rxc
QKgMQ1gDS0vKvRhMbMJ0I3eKUCQTCb75e6kByxcz9J96shmTUNeGQv1aW0qNp09s
IuD2RnGXFg3iCHIqjesSBQrZZzMT8QUNRk0T0K1Z4HreV+oaDFgNqhvzgkajy92O
gylXED20ITDqI32EPTDiyd2j0DwQ+VCka2ZpxQ7raT6brhhjUejCF/EWESZ2amp9
Dl6cZYL37J4vOzXk6WKkSeKkYgFahO5qTM/PBNXFZ06Bx0s+8m4EOIeQGgR1HoHy
clvdZ986C7vex7WX1eCR93VmvFy9OF83do6BZ05EP3Rjnbn+m9RXcZzCOQTfIVSn
VUafS+pUYgG3o4pQjWSRuV6ZJoKp/xyV8DJ/hP7Ri1w5dKV2iAkT4gy1GZ9liz0D
Rzjnjr8MlB39qBlNOQyoPcjHfNvZQm9hgcf86NUcgXFOH3Gy6IPpuNGhT490NjLA
gzgiDIqokF5h9Jds6uFpNK7z/Vjhh1oTG5dwFDGkwwGzj/YT8oXbfgVkVJxwkAps
genRvyQ5RuOFgayKcM+dMeOTaVifRa5FHR5LEBjXxbt5ffOzjHAM+lYgjpierI7w
o5+TUW9QuVVfn4+LBd/y07wq1djavS1s0390ipV0HqeqKvI68Mi9RecvoVrIw7aH
NgYeuotN2w7wDzJD7yWSYisUVTUtWTSqQ1Rrvhzj8zKUqkAd4ZLMLvrgLa5TcGp0
PJkn7ua6a4zVLRDuULU+bhpwQV+sOcnWxTP6g6khir0xWuYLCtw9jQub1fVWxi0S
+5CPGwQO06vjO4Trqkc1G3KBdOMtPPCwjjtOtn0y0fva1y0ESLYn0HAvdGvPXkYc
/4dSkAGtmM7CnO0KYH5s5fm6tM/SeBVPCjI+zV0BRKBQ8pNTfgcbq1WyW3eMZMaQ
GqWxClKWpR6K//+0MS6ifpK+MTjc903MmAsSxTt5EhV5kthpEv63xtqbx/ycDscL
kDVEmcTraVQd4VX6EupeqLwPYyCwxiQY9lhqyDRDWv7sM34wvEtb9m70AOregmWe
MBW75okdi13paWvaraBgObXfXrNv4c6lcy2yyB2EA4Y5b1eXaQ4D3Ia2MwOM9GbG
4I5C+Wk9GnsT93+5GgtMY6dqtJSlqbl4CTWmMItqXldjy36bUIbJmHFH+aCc0Vtz
iZk9O0fv1+xs75DvF/Gnh0pGUIaA2hHa5p5XTLo6j8UZ7WGYGTYUzZpT0mGv0fkM
yFD7sqttcuBhy6kqLSzMz1UwYdV5vFNokvLFMf2MKCK4i4L8wQobDd1fEM3QmBwX
kTo+xpbMu2P0ilslkQE01vwVVgjuWvf1SghXvviaSORFQjfEXSSIezHr/rf64r1K
verKhlFHaZnQYiRrgmJLMBU6e8DuuTZL/lHHD5breUvwxhIk4zFi3oTFYKxrabMt
RDF/W6eHtz68uz3WbJM5/kS4j7Yr3yN/r2wqjJpSnsVD9ah5DnMqNXNbgc+FFTQm
RxB4+5/iYNp07oLthj0QKVqBz/J+BD8uKk0op5iLgDxkdVL95rrerUX1bQ1DhXjT
clj4dH7WAY+CLHGR5Jc7Jel/yligvnSlGGGgpQXfSHFvR0UMi2R1NEA0dQXm5Wf0
lLNydCe1tHXmXBMGEsa+VauJEZBjTIVKEmS0mJXghXWQ+S+MNTsn7r87At/zovcu
g3pQmpa3+zpq8ESthb3tguXVNe/xpzXOGWvOYGfYDrT7CZs6bYH+QX+NaQnjB/BI
nWt0pt0QO1dEguxFKGgZK5EcEt/CFEG6jh20WJtL3yw6zWiF0OYg1GwOiKAnIegF
E++X3G++gGaFAoPmYtX4N6dJV7gP8BvoagCWr4aUDpaXXU3VdniMzuGGrPrE4V+b
N+mW8POKFxvEoWkmDUZilobpZYBNLki6PHNiXrqXufpuDscdLVTBUJWL0JGWhN1C
j+haNn2CvVNSH/eYvZrbEizrJRi0+W093jsfqX0DGpzQ0G2l4Cvyk1Pxy284Vv4i
WzcElAg5KUqukJ76jGeJHk324Uqx2Gr9XfO9xPxn1ee6vAnt10laBX1gxbSZMjle
OL/U+D/iwll57dgsz5GONYa+Z4FQJRtnbUKNPh1N83/wlh4EBRDa+Swk/JLJ3l5Y
fK+SgNCbTi6JnYESNHB/yKIN3PPQEqpDphAQtKySbsHUzJRsCaVVqMyp6eSNiQsn
ncNClV0/hIDFIu/9RaLCAdReHT1ZDpvKMDs264Qc1J67P9EXDWiSACzdajo1Tgm8
9ZjJbmicoPjyICT8pQXnXXua+d/mSL+qzpRfTbXlZO9LPZctVXh76e5Jf7jkCqr1
pzLpOvHqgzQRw9krVpFIdBn0tPQpInIETrk2DkMKg4psnOCf2Ca93J6fz70dnmhW
fUOG6FDs3ziwhKMpbYXZGrwyW49JZ1hwMDA4DTKt4gXfLK9dJI8B0WUI3c1kXU5j
cK0S0Ln9wndU4/C1P8vBTTmg6OsKn1m1fmyst/r/lwxem4EG1DPBEX0dGkkfpLlz
gxFx3K1LJc19imXLLDqBVAQtuWP1BIFiHUCxHuHkcQZRGs8wcVLxRlnltfbnLmzm
90x7u3CYifiD7OpkhNYuUfNr9OhyCW4oCDpSY5vQLKIuVbY+LFgGSDf4qTo6OgUj
346Gs2tFWDbAJwG3wzDCy2oogV4HspJhArQUKKsII4USWr/10x/TBZ4JOsnFcOdx
w2LpQDhVPS/tJD1V/X6bZDe1YbdIbhebxB6hbjmatMzMdYodk9Pz8s5jXOwNSx4h
UbwwY5IJr/S2fcHiGqNUt/rBKGdKfXvNSF86Jb3OD5j3/EhBlXlV/HhDMgR5q0Gr
FEJAKnBA2QBLCklO4T3GdQOt182lqxF4Vwm1YvCN4b9EVksrFeA1XSLV/AUAvJD0
0k+WO8nvqasWVPluqBK3r2m8uJckGLFxnHeSL7LUFueVvmEaLZXXPURGh8azg3k8
HvFHLsMnm0As+PgGin22m8jk46xQTHJdyDrdsOYCayoIN87MlyNBk5lXCq19VoST
02gMTGsyMDzuBRcyLZ8QkyFjfYx5EAYAWk8jfHbq4bjK6D081uqCvm5u83i3z5cW
s36GtX/LM+0Hm1K9AeTMnaaFqACJnnkVCBTR/jcH9X6duJjO3Qp+r3HNWkSyqGya
gT5eCI21uXSTUcBUBDrzheNdatwzQwOpnuFOBzbgzG1jllzqOjCkgJGeaicvQVzn
MnXS/fV9aoz8Z+e1AqQ74YVmN4rWOFYaR9eKTKzXdByR7ghQRS8zF8BL/Q1c3F+A
d12uAsf1t8evOTNt6xhLATnuvu69bbp5g8h3G+6Nw9bq7n/cQG8b/8+kP7TkHuS8
mStkBMkBbeaPMRMSmI1aqgYMHhnvhYDfBLCUCt//DeRJlc5KvxxwquRZ/DztZXYu
AtqSjcidluhf+R9R1xwQn8SwAzC4LnyKrg89yJEiwLxFK1h2Ngli2rGwYmVL4uvG
bOXE6W2XviI5bi6RdmGzUtH+SMScJncLnmoKkt0Am1WVwuoZdJbzLt1sSg7snVbV
I/veM5Xpj/96EZD0x4zZmGXKR2BFmP4vuTaGD+danbvWGAQXnvx3aYiIKQMSZVRC
Hw80cFeg8NuvQBLTJOR++0HT4QFAbk1xs0hUyQa8/sn/hdC2kROsnPr3LEQ1XgVK
hyqrkecto6TGx1t6da8y+n3x0VznI6zW+ij22NpJp6IBGrKivdpBmcWJ9sZuhDMW
eZYHp2HDJ2mcUiUI3fiW6K1qOak1FMBLpIudvnWlsxYKDMH2EavFuaCK/1nuzcGs
I6zrOfhD6Dx82zcxEWE8teawo+nmgnrD8sbKUpOqr5GxYTBFWj0MeqteaVdUUtKK
vGArvueZ+Ows1TeUyyiuqDSVhPMK8jJzgjxit4LC0BlNEOGybY5KwO2CMsMD0+1V
371F6tY2ye/JzvdXVsIgE81SVz3YgioDxBZkR9OWVz7WiZCkxBjsNuEtYCEFpi66
K3Kdx/f+YU2wEfHeAwZpZGqHbWPRh3dOynq0jaB1vhOBtJyawubJRx5I9lwdgWv8
vS9vrFyV0wrtSROKcrDezVV9vf1BcDwnN+Db6Z46JAA3stW6zMPxqOT8EEdrqVRU
gkvNCEL1LMrpWaCmn4K5mFI6V24Mh77R5s1w3KW1YS/qFxUACKVqFrWJplxPKqJE
Fri8SXW9vC4oKS5blS14B3dnkPhR6ENUtpMv0dg3yr57L1TKV5xFt9vwGsA0lgWe
9cn5XOH8AjOZWiUf38StQpFubh9T9zsrW+py3zCHjKKKBsP9eN7t2lNawWRUG7Nj
LjztCeqPF2qsIJOAIndOsy3Ya9o38wLIuKLx/8JhCjp5zoHmSi6ef3xtjNSr8ymM
e4gcXuPate95icwvO8HqqDIBXkDwH+KCWf0/EntV25jL1qbj3P7kDkBX0UrU5X/j
Qw8HCcHqhSKKuJEvFg2YbfzisRsaZlZRxWnmoJvZnOA7o04Osp2aP/knIeA7oerG
csHxhuZTFk8otlyLwCZAypKoDOM5gJkzpSNQpHJBG+BAMpCebsju1V0tIQw+j3hX
YWQXwD4QHV+3cUnOZ4aihn7+8p1sLmrzvgfZjfsFnEHqMuIbUr85OXYrnEXcyEaj
BtJ4wLh4EIh0AC3TrwMMtdYEzntdJVD0uTgg9l4CGghb99QoflMV1xzUG60Hvy4/
kwPiFkzYV4hXNKZVCMb7YlS6wVkheux6ny+MgxmtQgzjAwhOEGm+mZq38/yZqWgX
A3nHDoH7bowyePvwJ+tvFDafEi9RmVDkIaTQ7t4UofVrDzBEVUJGZ6TB2Nec4uQH
RJjunFbLwXao740yWA9IK8+UyVJ9IcI/mNmIK4AWVWCz2YVK4X+8qOmc2NFsBiZQ
37GpRRw+XGv+iQZX1PI17b6MwBktOZlRwB7HyGxqfX+Cvr5tkZW6pVFa7HHo3iS2
IKVsLCVULeJzYIiSKkYSdGs2StMCweyfz6p4EYM7M8BjE0W0Etl1nYXTT7r6QZh4
nUhOqgS106zNUgnBDyBeeWtYcuLN/bxGpKXxORJ3B7UeXXK6AvH5iK9fW/ZrobWC
Cu6Of6KzmQ7QtxHAxjdirNYTrl6uDa2+2zpIfOs+qteziUcshPREc4H2C/0NlsYz
Ad2bD4L4qYCrXZR6HKv5VP9THwafP2waF2lL6HiDxz8YdR0nFOE0G+fyv5G4AQnW
A0kQbcjxLXSHYxBgwBRj+JT/FnqR9Shok61nqDA6h9YMP3wbuSruux6hjxnXMfEa
HOTaawPITYEG4P8tqZRhEMfKBUuTtxTlSwH1pHwKvIdXCNwOhdBOscrQyOvJljTL
4GSMh11JU3e0zOgEDqBdqWcwWmOZ50ouOVUUjcSFDOxQCMxUWQ2tmHk/HLjmmeA7
UslXoDF8zwxX+D/SW1mxl21BZHwe3nb+c0O6bDawpSo5FhZFi6sBeXM+nXcXjul+
WbwM8oj50lfi9kHA69ij/YBgtYwj8jQvwsqHVgioLdMgRaEf9O1sz9PbjfzO+WPp
RDenYDtlXm+hkIi88JhWidXgWPykXpxG71RkaWmTFrqanhDfB6zYD9wpBx4bvr1N
5Ded8ojhvO5EIcCmX9mRib3kikDVxc1w2DjVA+cRfCrzgjUk5PYkSfYK4+kpL/r+
wAus8phQxZqk/hZ+yE8SzKku5Z1FZBMq/iiY72gbq15weFlG+Mlg3rL1BdCfiEDG
pvwOWlV4H/Y0uZC5Ax25xLRTPbuy72UH/ZCM49nDURSrte4u8inpkFck0XLOoad4
hsxiXmcf5PvssjuRD+QAB2acxVtykV5XZ1+0wRiGi1WOdgOBe1bzFNWuJET6+1Ys
RGkHK8As89Fk2v0X+IADFfWDYt9hpZB+ybHTOqiHfA+WcFxUaWzlqSn27tkwwWCr
qS0N9SL6bdf6P4xvoVOYOIZ0sTw0150g0XioDqsjBBAPNop4njXSFwGZB+JcjWUG
uRaubBLua554nddMUyNVpWzA6+wAMLaN/xp+6PyUFvIrbms2hzLPCFQVgNkRZkXY
Pjew/pjiUdc4g71moZOu84AmWh6Rp/KD60193BAI8MRMiw5+GlyMfR9YKS54uQEv
RmlIeBSRHyIrHevb3k3Z4VrSZVUhnl+d6vZB/7xmcQSkcM8dqRB9PQbAdj46dqxX
+nmK7N7jtvkwHz9EJrsy46/MYVh+YOBzUQ04WIQjW5umDMaYX7XAuLFPZWAxLJsN
pDUsKOTHLe3wKJl2+hZtJgCuxY/GKy6zA8Q5nN49NvD8jEKtTjAj97M36eBxChx0
0pugxDTlhISp8BrX4A9YN4Hfj7P15iNHbeEZGIBAsc358mX2poq3B1nQs6ITWCO7
l7u5KxkXofnPE8xOO7f8z50DqAEAtbhxnL7gkFVTradyIEYSbX0JXjLNdgF0+OlZ
4+eYl+zjahJ07RSpRODUKG7kIsGNzmVmqS2zZAQeIFAicdiD72bWTD9bdNLWoia4
RGTu/Hl0aRKIsjpofk6Z7iYdwTD8hn5cy7elgKmXOi5abQGNAbPSvw6JklgzeLfq
CWl/w2UTMvZO3nB1KqvwILJVN6ikg4CzBlCViVItUslCWHXYr0P8DNOWcgsDJURN
fsYWQy7vW5YF+8FjGDG7GY6wuqtl44pPBx/oauLwMpCQU3xyqbVV5yGj8i2lNk7z
5QT/31SGO5WZimKEuXY3xWr1o/4nc8rbxKlPKAveteatJJv7HCAVYxKT0uaLRie+
6xm6AACWDugHvrehTn22eJHFtWL4gyyzhUAb6F1+zv3TlCGebm+ah+rtMsdBbG48
NqUoxNEjm5cG8BAe2P59LJz1KwnqP2hUhBcicT/+hJw0Phh6+zaqVdd4GMw+Oz0N
QBvj40YROSpO9PPGSBWUPIJ2Epp5rHezUHYeQ2vMI00OqBHoWSadi6nGKU4LBO56
i+eLScF4Z7/6WCTxDP6/KlsPJxsTqsB4tzcry/rfx1eL2jsQUiKByErn/YEK6oVj
mhCj/vVgDYodnwcK+31ZpDd2bRrEHDpOJzDWCda1U9p1rF3Ys7cXCQ1nz0iXEjNl
y6zx+uXRNChV1vvc+5y2/n37qsLdo1uFAJWsQHkQ1D1OxCBOpoBmU1PFWMSlTUje
CDM6tXQvHnpMQ1v1tKb+agScHzb5+b0F5pQwohQ2tYTdjiT7ySSHOIzNm542gRCj
w2SVtMzdBPg2F3nKQ060HxbJPvkFityq/kZkoJzynjqTQTbnL9ITFitZdMVph9ik
7IB3hvDHkBgSlv9M3yTlGLLekDBvVLMPJ1kZdfDvhO3rwRM3hBmKWLZN7AZ9nW4X
MSNkAgOYZIQQyaE+cN8utN+tJnmCdwXwhRPpYgDblXI0M1iK2jGQOL5a0cIqdjBv
ThvTLElbAibQu689DuYB1dOrTOY9SmrmP7cDPCZeBsNEKNOeiWQOYlPSD1SWyyMQ
H5moUEruQKnrmXhHVJJJtfK8elVi2foSe79SyWrlQgD+5x33uRPCw0rXwgNfMSrB
Do1ye8M+Izd/PzGWeGIzw0qGpgUqPf7IlfIyUcWKjnIRmT6FV4qO56zr7Ma5s8p4
qJfpSr3AJM05ZEql7TDU/qSBuhnjeYLRHY+7OgWIgWDimHLbzIrjUkF+oocmj6sV
C70iIBJtQLLzmcqgeKZfosnvVt7ATLktBqAwZe/QiAhZhnZlrUaO2r+E2CZizgWa
TRngo3lfjIyvRDDI2opeFAYI8PthjJRKbRxDnfBwPDiRQnZGUcI6Ie8LRMV4TnTP
Quv1Z9G3BMwMY/xcqM7c19lAD6FIlMAY6/JD5tNZVbvFRSUopYok3t3qKi+pxcBr
FrEOLxsHorNTVEM04LnxUOpiZ1YlwtYLHX6kZXeG7xQEb1x4vEo0q/mXe+h88PLc
C4kvdroyRuPEA4M4dVhlA46IMmtamcB3J3MfdDDHFsklcPca/ShXBXciDAug/rnT
tBzqR4veQ5ULZJXSq6dqyK0RT6WVvEZSkjCWybWLOnvinQT4IJDLvZ5nQxw9YbIA
KB0Ju9Y8tDlZtCjzTZcaAHmKbn3yG8GAZKU2BFS/0ABpKq2aRUO3e7ITtgcVJDlj
S/ZoQKEgaS0GNzAg0SOoQlNMzXqCqJbXGVzhW5mcIZT7stR7geXv0+OXW3oM+sLR
2Fnac/n89ROomEg+9aSuXAuAebD6UPwcbgSpttK2hRfLcNkkI3v74CsbeIKXqIaC
/1w0SsQHfTXZBPcJaFhPp9mQ5YeGJTcqapcH48Fi+FC9Qyp2RcqhpED1JC5ll0ZZ
3LeJqp+B/WMuBtrQP7KBVKHUCjG+gsZx8GcpEUd9WarGERfZ2Y4JZsC6K9QUsBrS
b6VOrU+5yEa4IkADH8svT7eWf15DZVVOnOQY4sxZw6XhvFICltNKuRx2v43heLV6
oZu8nbynIpvBZiiepcbtS2uO+rkjgOTp4t3bOB4+euCdE0L22rp4+SNzlsKG45sx
D+f/glnaMrfAjSF4H9tc/+AgWDlIJYTabub7/RD8XfgsJNQK+BOuK0Or3u7BsiHv
nHiTx5eHhCc/2iOoDrb826/wmDp9h+usfn7bbmspwA+62/uiylYIi2xAK/BvS+Wm
lPFlUNSSQWB/xOH8SSD9/WyPP4PXt4NdfgjVIet+y9FYSpp4S7ChIGlkCHw2+Loo
v++6S8BCaD4NewWWBH87rIoiMSXRU2WHB5KETfl9dhiLZ9AdlpMgGIIPmDX3tm0+
twStN6mA/EtCkUpKTuUOZwjFg9bBiDToXJc0g2fUsEVIo+WT0Lixxd/6+M+NRBO0
Qtaw5EXgl9GucRyMr8Kqin7RLnZaFIRqBohp/wDWyJLDjidcopbV94IRkg9+rfd5
Jwg6tV70UMrpyV76fBuCKa+PqvYbMnmCSBWPjVOyardmt8sqiGdp1LUzGVf6R+E5
we7k0vlPkXG4GC2SWVBoBvcYvJSnzJs35VbbuP8Yj/Hx2YpYuUbbxH13iMqBP8vy
j3MQdBRSjztKU5RmuA4wVbSSQr/PO5S5IWWlJfZ69N3jClkxWpOwvFMfomY5kT6w
UkTkzNS/XuCrB5db1Ri5WjxaYfRPib0ISm+S4EVciUBmFKmdzwn1Qc/PJe6NLBQE
fNhLdhqHWIZ7ePH/+LXytC/hd4GpnN8jY1R8mJI1tiOTu+9t8WbQ2UIsko5Q65Wn
p1UOqYIzMfsYDaU6ccr+sHnDCRulqI/KMbEagpJFsVh8jUGU328FVsdKXMvgROxF
imS/ayB0brGW0QbNjVQSkzchI28bMkI/LbGCLp0dFIXPExvr3YRAkT83ybHK8qc1
QzHzS0BSrteGmw3SBRAWWiNgB2rckQK38huKWByR9oG86IItJCXGH04TfBs8HkO/
P9/yDDuv6xN25gM9sONDVKUPj3BWnOLptQhrvQOQ3ahzi7jSjVlKrjGJKDcLu0C2
F5+zq8e752iuyoHPo/ln/7Fd97o97K5iy/tXAJkxYWA/WmdKqQpBfo4XaogxVET3
lKTnh6tWtiHLopX4AFfUEdN5ZCSTjQt3Q9HYz+cvfIXMIE5wFgy/rbcUHAAhhw0U
wOjK4QEDAKnukqRDgL/HnUQkVh71njoSB/8dSbCz5c9yJjqFlc12oLWiJI1HgaHV
NPP5L7PnjAGt+ZJU4GJgJWJfvlqaEXCJQLb3XYxMoviac2t6kWCWHoZKFc1Yo3du
ec/3FUTTErOEAA2lbzwkfIvXRzhk6hgf5i3uGW2XzW4J4W1wr9inlAhGR5wiHVkQ
W4M9nILyOvV/H98fg180fhZqleVVb/yld4TLXLZcRTjTvdKfjex8xHlNZMouTdVZ
2f0Jp6UMko4C/JSaDQz82BGs22jKZBCQ410GdMZlK/2dP9v1X8PXCIgXlBIiwUcb
foML2ooDfINMbschrGbivZmRJspCSKRbmd2TZA15jNfy2N9KECyhsmd70Zgei9DY
E3bEV1hXBmfTNWxpdkPGBPBkIcKp1/rLvwu+h9pLpQIbvJoCbjG9dQeW9bNdZOkM
vaZ06I6twaEU9AVilEBNmi2V458xlo+g+2Rbqw087I2AWDkLY6RooHy9FhemhoDr
hb0T9kzkVbCxW34X0UwnHvZlPfoE6PW+Q1UwKTdJHWr4Y2oTBuM12ANWE2a6BUnl
It71Ead1zxqH/3UPEx8joJv0KKC+NOzydDy2ZV74sRmRj0upaKumnikvW/g1jYiF
7J28wXSmHpVLOEUP7WgDAT9HeRwyl7ToyEpGPOHNOqZTs59IlieYxTbzqnAuxoCN
QQrkpLspv0uLpSqO7jif+11KenNkhZqvHrsLUojxf/WqbcKNSB6DWNQJvagK/jJ0
d/lUtBswV+7+xRfBgCrrDlOMCgfOgBJy3txguv5YfRZBH/f+w6A/wPaxFyq/dddK
XUxjKq8ptDkjpuep3Olr/wuBB/yek5VytJ+zeCP4lRkr5TtL1dLCv2F8fid7xP2E
Qapm/Hzd9F3p/YS1cCIQSQfsYz5nrY5extel9GPG7Hk8rVUSj2Ivzb4ZFqxYetSO
vHLYObdNKRmzvGOEai8wwlt2LptEgYb7Xr40z6aqkWLRsPqcPuUjv8/l6AZv1Z82
R4um6Dzecs6yzbgie1/Dq9KxWkfP0iPCvfkAkgZoo6jtgpo/WfiEDO+LjCzhsqEl
3/bKwvKnrF28L9ZHajmmtuoOCPSmcPSghOETowooVvrVA4H01FPUa08Q7G+GlgsP
C04VvWOAkX6wf+i+E8DGOgdXq5DSCzEfsXMZ/vZ8qxVqm0efT1MxTl64WNeW+/Lh
sNRKEwTP7Fli9Zpqz9VgxIFFY1E9R6cIAcllb+qr2jNy/1TaCuwjha2FRWvG176R
PY+2hwVYPe1xVNNYTzcqi5Tu728vC9+og023tGSDifSwHMcoKFVU6TqXX9AlCnlZ
Qd7lj2nj88aaxQIwTG2JTA/kKue8BFlPcifE8CqImw5ZdRdb6y2EPRF3R1o5hJv2
e0qkl0CqXmltnZbSJiA0TYI1xO0uRasa43KWgRkcDsgxXxr2f5itbrLaEfWxIqZ4
b3wv63TLS96lG3bvzfo0aKMeuP88i6Op6IKHQ8o4EaR2WQjLA1s6qafnV9XmaqVH
CxTFEZk7NoVxHLLcZZYFEP3L8EEruXuBrQuldsMLwBowFi4vUKSD6OlhLQrbHmbz
g1BSUw0/YZKURTRiGkJByDAAmpqBXQ8PIiFlrkBOmFH8NyYjuqBfWzXL/axlmH1X
lmNBOh7hmWXG6ZgSAX3VyFd4a0fPUcQUeimhCL+Dzy/v81IdSbnVNE4Z9bzWkWx0
LLIX/k+lkYLASayOaqZu3EyFeW7Yr8/Tpfj+0hIY9T4fl5lkyLmSFERSDX75KP97
M6xgtFfUayKx2xy9sr8yBtZTGwHcnCj/B4iAuABFEFpEo30UCl1lfWaf0/hF8YN2
yVgFDLrCFs0EeFkizlqeXrWHLmWg32RLuJi9UKdI8aD8FbKaPLEE9gQEVMC7vASa
l1beaxt7nvZcsV/lmgUoxQxm9G1I8gpWtZpQZbIfEdB+S2b8nap+ljl+iqcPJFpG
AH9Xb0wINV6r8V5d5foCl4EfuNmfF1KWkuiqhQDixxAcin/wZb7Pq93mEwU4seHh
tSHckTZ5FQGoJVXAr6oyi8cqKPcI6F4pqQmCpu/rz4DU/cX1Jx+K/B2bQ3DtiyNv
ERsL2bDclkUB4g0rjq/lYLRjTZMjFtLC6A+xjjaEBvFNEgkVkCqY8LJhdjd4rN5S
f/67skHN/LODMAGKj5/4zlOyg8hYJuDpFRRsl1sArg/nStulgaOzIl1HCkvtGfZK
3ViRWqNkoWcP/o2gKMsmh9GDc8ue5pkJmYdkVF3ssfCOuRLg39I8Y6MNagfCmGKN
P/15Gb3CXPtvKoWDauOiHDhvTK0tmQxXNbttr/tcrYZvKxitLT2kGcSvwbKAAQhf
j8MtU7m3Kd12jTKW7wAN/3uRJV5riDT02Z4R6AgfljNRlTNlxnXc7YNn333X5Anq
26T8AqZaavBLykzJzddy8sE6fWM/LuhAnqscsnbTtjiqCcrnyEJkNukH/P+izyvP
ey8Fpwzdmh3ZNMRbApMfR6OHFYzz90xLAvmVROBc9ujySI+BNiN2h1RWJIVhW1ES
/oWbMCRn4Y1nBUfxh/GMg6V2njIJ8FzyWptz+V6hQCe/sSryt4b9O/lPGbyzlDyJ
QgClzAo9NG3GZmbvNYR9uaZxAGdQXrfou4EQjorx58ou+EOu1gwgfxul5iDK+uDT
axKxGNhfvE7D8XHX7HuwM4m2l4wGnDVTVlL0QnBv8feH7ZNnzs5QD6ICFxIyVpkk
KLdydlaymQAd4KY5woPp9ZHHp4B81Ql6t2myF3wb9InRP+cNvd/NaTw/5wVcKTf2
9miDG8qE+oidwXKQcRJxN77k52mThVyK048GFIQ0EqofuyQmQcvrSawmPiLjJ9gZ
9NTXgKqoMnat1XzJi4VPrDo+TrFnnre2+B/ei98woEK0u3XQtg+FZLpmqZ/ZNcdZ
jkATGqCY9sHfU1q+q/XxhmBAA1f7GUpHetS3n+E73sSBegBQn79Uil64H61RR+NN
35WNdUnl3e5gmt/hFaXSpcmfmH6Xh2i1In5AO9MTcJnU8mtWELVcEUGMF7wJToZS
QgugQUPCxf/4TUoi8tjl8i5a+ij88WKe2neY6fu2cVSYY3m87dLnxBqBu0rROlAn
AVz15sD1jmyU8H5+69QdsvOEqga8x6YfkejCC+VzEumHL9T9aDTcBhgt+Vm4C4Zx
o2b24bg95E8FZygbJaPL7zQIsQYk0reAzNJ+kMqI1Y2y5GpEZ/cACVrEieuK7263
H1EbjDnlmQrJJ3B+5q7SGam9ky7BQOOwfbN3VFVUZmjFTXinHQ9Q6pRI3j125EHg
MsUEf+mhlsKcH6eqOCrEPqaBgt73dwc0ic81BpxXQyzJa22qMcJgwXhcVscDzuNw
9sb+aKab1kMYiKNyQJF1d9/Yy838LDwIV7HseOmzSHjksWjRIDqC27DPjBKxo8pv
tELHWLIcTbkeAZDqIZyXrFjSVtl7A+uyM9YEEgywaZt7IcBI4OwgXq2BM/xV4IcL
GnxRHz373re2WA1z707UPOx4LYUjzfDzm8hcfCyopEh/VARzvIqG0oRpjt8fqIrq
LWl0JXM7vXdnJrinIKmKI5qBnFcWc+i1hIt7fl0nuzDLBf+qZS4fX3rYRkEc+Nyy
7lsgIVNqz/OHTCQnNSMpAohfJrkKZlr0EsS67yJUc2uiSexoF1g1SMEP1iL1di+B
Cpe8f4fRmEbkun0SefRVSf7YZY/g0RgFZ+yiQETu8IiyXOcLlNAQdmyzRv29kQ95
OCs6gSdoY208yFMcJAKipz9vzb/Z/NnkB0K1sh6BB66b9Pu10RRxBPFT2kp8uXeY
hJKlyAsWUCU89ElJAsH4bnGxNkFvyoDaOKkXzb1G82Vnts7X5Sgh2TReFDxfsJbA
DNXY850mJ3CFCUoGxbriIh3sWBkXB0hg1rD6R7CeTLCgVZSwwjF/tA0h2DXBOCFe
ZFP2c1EP6Czci127EPif0kWzJgRF29wqkqnVeV3cRzlRuTysv6awQOInGUpl5hUT
VtRp2zvmOcyla2yxNy4vSNhdr6nKIJafQWIUWkcMaa5nLJQUts0KUy34CRCb41eP
Iyo+uGgr9zc3ytCLz0qHEmW1QZH4T4zyT/7UqmBlgO+fjgNUPBBfkNr44L0im8FH
1ZjQH0ijqCGjikm9H5BBLpWFhKZY9ItFTPmzJOZsHG1fuHvlv+YCNuP6NezYlqkg
oZRpz07Qpi+eTNXi0bEDlgHrGcwFdnqPkxjGKHcyRn+NIXcxbnbvjCs7cPBbnzca
XtnrWp30ai7BByygFMiRvcDbBJIP8xteSSKAGom+RPm4CvCAos4K2Ldyi67uekCM
+mF4c0mEnR0p0CLiF8fgcFfRECoRIdmXfY3sc2IHpyCjtgYSsv75oIPZxSRZiQ/g
hjc1TsJtQqrs7/g1GuhphHrxt9kcOUUAEqB+Lsc0TIEKX0m9mZQEx0ECPzkzFjRr
nx1/gRW2vA0KeI2bO9SCQKnAz12DcD6N6hxowhgguEAqOxBd2OTWhs2HRC7RnQHa
yma1K3aYhn+pxesOVpfTmfTzWrcPGltyhdZM5/ZQhueeyLh9jtCyoq1mb6Ivsqdj
QzIPEKU1h/cg9nSrDqamW3ceKrjLaUly7M/fSjUJHYCQmFOQz4RAkWta5OnYizkK
G5H2+7VPTUpuojaBVzLkd1JdJW/ZhJBX3gDz5Nxw0+HEhAYcWSHkH/m7qXV32+uJ
dE/M2OmjjRnq5s/QWBy9z41Dn2AxrewBUge1uKBjOYqMwneMQHuyiDBPrYaGU6q9
l1i3l9GYBNPR55l4AFoYclIZZEdoY2IW6WJQTB2nVZNNZCi2JTmSoufxGFPsTcpV
JPuxKpYa6J5CdcnMbB+FNQm3PEui1yugGZhAPB1AHmI5+n3DvykYqR8Q/gIg1QSS
afDJ19aWOGYycL3ZkUi2hta4LFAsNLnIKUlmAZacUBR19ZO0DNEFoviGuKldnHZC
nShFPT8DzDVKkjc4f0djF7DH6f2HEYiKOM3QNaO8gZzuDXz7fG5YpbMO+4M200X5
5XSKxf8y+NMXW06UfIC66vdRW/4IqFWcNWu7zWD1fisZ2Aii3pvPBntn6INuC/SB
GY+iitrd/KlBACtn3sQk7PdZ9bCTOCMddj4y0uHHAc9bjOus7z5nvlCMfSCqzSNE
BH1Ji9ROatVacIGnqs1aXQxCXcWLQ7mZcNxMTltH1kxfMiMo1JB1owBCSMTGg8m1
+HQgvvyg01H3dVFxAsLiEGrysBlMoH9tnRjllJ0bWPJtHycrjEtlE5fFbpX3duUe
P2Hzvp/VBJyctR/LZtCEZq1bjjwD90jTAR4S064Lx3OoBmxobtfga+M2WPcBc3zu
dhBD2tbfSYJaAatmHiG3CL3TGK8N1LPX7nZZejImaHXZaugQToIPS+0ef+iSP4WT
S1NDEdGqoxp3XetOiDPwIiC9rZV2qx/RnOjajmXEUdOpQCfHXr2GdM6jyt7xnZFX
kn7fLGSsNkx36rPWHrUVdz+pa96kKfQekAItVgwwfBWb9fiZQ8EK209FK0+UstY+
GKuDYKCB3ZtchYJwFkhmWTZodfAb7/PwuCaTeFCyiXp7B/U8qOJn6qpn0ZJIWUrj
i6ZbEOF57kLFf097Z+zRXMDMDWkc7GZai5PUJ4go8If3wEiIcFYoSXAYV0t018pR
qtqz2ceyKUpOzswHF2fMDFNtG7gfL88rO9380qUvBpAVWazAEMP86LYIXoiLLxwo
0Cnd9b920gRzobX+vZpq5b9WdkGg4xsWl0Ni85Z1ToiUVt+qjxoFu+rsNztGBujP
bqKVb/6peTU9+cZCuGr5QCXQlNQeMYUdTbaPQayjOLMilFgOcQ2+OOWLdpfDei2s
92Jjs2HcVsxG4Rc4XyRJZYlZZ2DFcfbpNu8HTvJNULM2L+CmWuJSQszDH1nCwqXk
eaUAqP0rrIyu4WJI44QHqJ++7Fk7gxs3htQPcf4F6hdLITPYCfCaBDBBVkWaBE9t
h3OwJEgWcd4HLTC16abh/6ylv6ZV8uvHhGxE52Lc0cYrzsUY2C6rBVPX+h/bY4Wu
6ZVcJcXXNssCx/7MzHc6ydJ9rQV2z59ICPW/6nWB/zgN3gEmqlRp3qII3OYRa9Pw
NrcL3HVHivfssg9Tr/X6CzN/HmGV5Jb/R3jn6uozingOvvyZ5/dAls7JjSmdXWcU
vo/Dg0V08N8M/uj1w9phlyhQ34B9f147Sy+O9MKfUL1glBVjBQTiInwi7Shcbp2i
DHcEbseXIy2Ea5DZLmLPdH12NhZDr9SFJZQa5s2J5qJMdTOgmMRumi4AJVNL3KB7
Bmh6EoammYpFkTkHCgbEu2VHzXQW77/gFvlNPmnT2u87cpy+yc32To5zcu/9zzMs
u/S4PXt1ivWufr0YQT4LnGdMTlPpBOB129lHZh27coJqrGaCA8WbPSedmlZm065T
Qh3d9VYrg9sfN8O3VniPYYNIXqZoOp2o+QsLPLUe2TToilvMyNVh1s+TkjgHpmiV
8m/KQpU1bfKpRQVjYEmyLrtNByEIl4wxYsBTq6nl8Lh1NHpn0xJJMlkPhWP8lA2v
4U2uXOOOT4CaNmqp0WEO5c9BU74bqgl6Q3YdGTHnbB3jljJKLheYZIDsNA9v/f0i
rlnxlzROhZl+5idEIafedzD856ae5vbXci7JnKLo/7oN519ti8V02aBs1Xligtqh
iNYCh1fPHC6oShvqP5YVVM3MBri1gVOyyjuvVDAIqC5uiujdcROYdfyPHBRJ9Ir3
u2j5z2uI1rWI+QGoJSQLkyty6O4RLjKmP9X71z3z7w+oVCp7lhxo5X29sqxRtQ9F
h1c65FAPkg1IYcjNAJcnJedVZ+BMj8HKJz8hkwT0/foYRJBBtN2+41fi9vJs+aXI
+P5q4Uqxf5b5JrF4TFrRN1m9Uf233lKj/7YmkgAF3KZ1i0eUemabjF0pLnsLAM5S
OZFSSjVyG8zM9ZMwWa4yyvHxbFqYzeR8JDKCsljKrI2E7D5vK82/+OOJFDZ8uUA2
a0km3kmUpK0l4KFh8DqPqMs5fFjN6jp0dtUq+RHOTAnxy4OpgJj4MXFATeD/fVsd
VE6/nu0XGH32cvU1Iu0BhauJ373XsFmhVdoATXSVGCiI5mnAC/6JgbOMCMC1rKc4
g0NhZjAjnBzE0wa6KHvasGuGGsoxgMuqVsQ6krTbRRPH0Zfh2cU1i1w1M3tRg/li
2JjA3FWWk8zVWzG1wzY5h+u2lD/NMamvCzKcpsqDzQbmou1BMs7T0TMeJllP+xVd
VuajSjlduONgYTH/QwOP2OEiN5bD09PteREfS0vWzomAMm5baWwqlUbK/MyOYvQp
ntx3MaqBLsW6d3wDZFewjmjFyzaIAI8LggWrH9ExcseiCCLxsUDavWOO6WD4EnLE
tBQM2iRVKDJxGJH4A7WCWM3MTbdf+0hfctkaWfwaET6NYGO+a+O9iKe6yaKrquA2
hK+5MpzAThwxO7HRiaxk3PzO+lp3N4XBVXI5x+oSa26fHQP7h5DK9bfGCto2Tk2g
hz2ogVhoqCVkTu++77adzPNYVJF+g11ZOTxksVkob0c6Lr1FhmEX1lfLhWhjAR21
d4aUs9iLS4FDzSrdfJ6LvGixtInvKK5BhOZuAEI+hZNW01t+MmY9WZUgahnJ1ClC
9sxjM6M3Xs4GsV67zVhBeke8xpKMzLwvQ5dcuLf7/nf3+OOo01nyCqvBJ9t5Qads
lcItA0oQhGnODAaceE8f6rAwVJJhPDChn2J71BP+y5RgqVGeLrv6n2/ErSma00uE
V+2pe9Sh/EfX4ZrmWWlpAciQts/QeuMhXdB9Sj58dvs9AZ5n9mOaWtPckOvXSURb
HyflmcJHnPcaXO5v5Sk85XRvl6i2MFd/10yM+s2e5I45aZgQblTYTXpRNKEabsWp
ZhaG65FpMaEZTc6VzedlQ3jFUbhd7F4ErytLAs6TB1OaUAIfhFgDIZ6cYU0pYW1y
EffxsVvD+J1yT6TwNeU7EAaQ/C7BBOREJvZ8C7+uEHB7UJTlUjPMy46V/yfScboO
/UXEth4XKq94ShOyl2FteHmvQ7mEggUODxkjoCGuEcXp++wpDltLif3mHCAvCDMh
2auWcgupACgF7ZRx9sTgEopR14OVtAFi30V5EAHgWT57FDyVOIugNj1pUu/vlZCx
78G08sn/rbuMt53f45eY0DhiYILJvpgWirPPVNJOdxMrgd3kW5/ES6YBB8yW+t5y
R0KMWB1vFeghBSy6ZWRlkO8qGqP/Mwrs34k5z+jFY74lz3XvxwOPwPPqbRQ5doyy
WE0KKbFpLiJboDS0bYs+pYkBxNQyvuUJF479hQHouiyHNg8GU8HEG9+2uLh7RhIY
JlXtMNnsNkwXeEedbl8modeouZ4NzIGcyzozFELb4i8mN5vajFsqRNA/2dgKQUbk
iW+oJRr6H749ZZ7hFMtAXBtKOiGT2bMOnACSE3P03yV44yC5ZGftKNrkfhq6EIA1
HAZwVV8ULm0dpsobVP6tIwYigUoRRzlRExcVbQeGN1SpJa3U8YqCNfzexenPDPP/
TaITN4uaBPGREAbpAzk1rbmTsVHCK99JLVmC7th8MaW31/pQVQa8zA46Zkdx1T05
GICM0fYskZti2alZHxZqHC+/LJFgX9J0gUuYRD2B/W8wjzX7jidxkMTiRKi0u48h
ngD4+3jsAQOMljDv2krahIikwjOnMimYPXss0Wd92q/TUs8MiqoLFpVd1DwCuhtq
Ne6QLpxpyXqV4Hf24Uoy2/2eESNRW2+AhBzRv4mXda39QHPo6kRwRkcEHwSG2FbB
fdVzb0yoxwMczQzIiVI+N5OMmq8vNVhOEULD7jxSeEIu3p/ftVdT5cUGLFiFOKN+
zcsnp6IFRjat+jZdxuaRad7SP5afJF7DGdOYhNpIcCXROzv3C5Ax8/xe2myGl5R9
ifZctX0tHDX6nsy3x1VwFGgFg/8UfAVTT6NqdunSnco2BwKWz028isWdIioYmC5k
0KJzjE5p73m2at4FmPg4qIFSLbiuRAGMZbxh2R0A4W4wZsGZtQpmLP3M3gYqAcgl
gQwhnBw3nbhE8JXTfAxsNRTnDQ0lP7CjTGFEbqL0eKz8g6Ttw3qKOlhtACFiaX1A
7Elo22qHlcdMS6QTzbeNK3S+yBZ2hvVRl1gDDnAUjKZnVxzrrUxfeboIhKSWP+s7
b3V2Bzjw47TdwrVTQDL3XoYLyFMIQMF93HwT5yvvL4cLQdeM6RShlyy/BkkT700o
+fpYkHoNdPOhMvYEEC857lq9hVxsVgzXTIRx3Ys4/HisH20d7LPVehu4IJmWCkc8
ycGbwFYRfLTSMno4tgiHG4hR8LXbrzEhrbPqSwKd4vll/LDxT28JIlpfxD3PE0Qr
jtpXAYvWFP1ythJ4kNipxlnOsy3P+R2nFhcwvwwyY2tJp4olsKUMZtl6AxoOw+YP
+jbFJ/Eh2mJWxrVrIyb+Wx/qhjAEjbgagXJJnWjQykKYOGnopSRCtAV8dyRsyzdH
rF5POO9UC1kXK5YT6wkz9OHoh7MjVKdklVXu/xmjlQI9ITxFzkkwDk611MNg5ito
eySkUmYepUeNAl3F81wEC7k5845GHn4TxV1jmwE8rI4IAq2Bbd41o1XO7dvyTK77
8EsElNwcnl2AGK4UiloXRrn4n+EnQcPLKYudeYKjMGaOQsGxSWnpZl54292DblJC
6yOtzc74v2P8+qMm4M0QpvqGkIgapvAEmEa9d1blRHw5G7jWieeO4grEh2Z/bqJc
C4RgYIdjQW/dOIIDS5MDWZw/pjRIoHe/7+7THez3Avqf+u6OZnA2xAHHCDtexspo
o0NPbtNqC+8pWNmas6NE+ZoPJmEJ8QTgqXKF9su020TxCIN2Np3bGnWnDceqEDw1
rzmbrTYFxPF9L46Dx7zXJ+XIrK3fAPGB6QaLLg/Jrr5/xIm8As+deINxuzBsyfno
JhvqSnj8AtUUZpVBkuK8RlTyCyxj6Ua2rLc+kZdHVRBx+zjW6xCOIthfBcJTNT/n
ezvcAeYnN4JCGW2npnTJO3YFVWcXp0g2Itu9tcf/6x7rL2TrvG1aPMZ8YKN9cATZ
kTrXnVObzJqrDJPwTr9LQORI9FXR3j173oilg4pH/UkD2qaMomU0qjV7b9LCVa5Q
JES+8Q9n+PQ+86dMqcRxChx/Se5h63yz2KCYY5MKDEh+0dL7PEKL4Rr81BnuMALc
NM+CCDl0wGJmA+gnsQqFEMrvjKYj4CwuCNtFCdBuDKzPWLreee6dk5100QPG6EQs
kvsEHQsO/6XYNdmUiJvZsLvhm0jQlnp5yw+kncbrNQFs2t/iR2pNuUAYnebCtYkc
wvrd9TsQ5xBYxYPJkUQtCUvLw5Yig6sClCf86fUg4S0IRrTSqHCGsSKI6Pj5q22X
E+t4e0bulprsVMVxaDIG5QI+n3zE1vzCUcfNrB4QLoXCZYeQzoTPCID1YzFs6imE
BWx1pSu2/XCZadqpdwjn5ekSwV+Y7c21LeBQOdsxxh1tY20cYdmxLsaHCxzIvRdo
zNSvPX8S+1UL7l3hAcI7wwi5KAWRa3It5IICueYiG3rbIvLJ8+YT6ONYwfkWR2mH
sWGu0inBr5IjLdfZrCQQSWrjoIQQFPStUjsutJJPXTFFl0lxj+YFG0DhC3/k/FEr
2XCjYQ+86W6caKKFnfqT82y0F6dGixov+mfgIUPj0pvKSPAfiL+vdf/Qha1sKY9Q
4JA+CK3L5Zo337x0LWGko/Vee6fUqmH8HT/E7Dd/m/XN42E9V8khmT8EK28CS1y9
UGcEF+MHtRPNx/J8sfpGHoGeL5/i6QDFrO/8qP3TCqPTJ+CaMQ08VVAb5SAg5SY0
d0hWI68imDL3ixTlklNhNfDqyZp2283Rnx3TvjPMk3q+Tfpp7zGkhW/qzDIdyCn4
3jTOoMEM49Rt2k5qv5GIqOfcf8wh1ARwpzcxG0C1a83y5tX1uS3ekvA9uJ2lf8R1
OKVWXvuxdUuBZY/ijxxhlcjtnwoNG5GdErQ4GIpVpKn+Z02jePrlNWlsiDHLf4Wz
72pZLnX9inE2UOGX6k2MqWWrdhJVLZpTNzr94s1yBKtdNtXUL53KbH/HIYWmCuSt
xgc0zHVhIhbigCwPMUVsyAWRPDKLHdXNuxV+odAMYPkAO2dB3tpKxSqElIbx6ekl
aT0vqdESd9aLNMmQzLxIl2md6pbkTu8GdbomzA9c/J6PrmUP3PtVphP1Y0wfi2jc
uYIJuo4Egi7/ZTc9aE/lp9ba2vMFXbpy/Oe6nJkehYdXwcVsCoQN6nC6hwlbI1PC
ar4fJBcECtSEJiqP6YGmTeDDneAOWqJIriS1S3KKDNAFKbtJdnFqkXvH2BYgG9ZC
RkHcIQd7LhY2fVq43bYSViIjW20RWQfxwF+a2AHODyLl21SNg/qo+LC4TJzGfTL9
tFpF4DqkxC9yrg3nhwMgpuiUJ/p0X9pBjtk0OO0bn8yyvSq/el13DCVSCagI2xsS
oIH3f7sbC9KWmfCkWarMn4rwl4HSoIp4elthn6GJND8VoWT/3Fxn881qhIp+U6av
QKSmb2MhkPDXqC2O65CqkO/FuaibPD4F7vp2yhHc3mUoX9jF7VL4+g3c91lmjt5C
+L8DjBmxIGzcCjvXvWjmtecPdq8Ov5/MxRjasksNDa+7dG+kYwS2mUYLudoYHihJ
QojjR02JbOG/gdrUhPVmspeIsV6rg2+wTCqq9Xz4osS2tOIjbzEICvplUaiKDubJ
k3MDNIyes3mtq7ggwHIbfDR3Cpgk0ebIEr+/CujlwJH7QbpapY8q//BOmfqk/tSS
+aArw3BudQmsbM/j/3EJRzMI2GDA416ZGHndnd42xGpF6URHY8NBVpC1VO4DtYJ/
q3wVHTTP8NrSmiqo1jbwXz+yD6k+eJQsBmzXcXGUm+VT40ZW/aEdFqP/7GLs7/yX
ritzbbNXQp09U6gzrGUqLxjX8xpGW8OZYHcXNfByeDzFtYh2Qdp17/GKY/RaHFmU
MY7mJWuOlgxn7Om7MLif7rOFbUhgX3PK+iP+D07Y4DEnDzNgYwg6BmHzUOiu1QWe
x7mkKWa4tsPyPIBl+OhliYOi1vAkH2F55HY8vAS4XjhraYALzlKB1OInCUQkE/4R
Y09dyVLJb9RoKyaFsev4aT5JX64ka4ZhBwVYICEQ2uWxJbiV/cCfcd4pIpINaJAi
enh+76oc3p+o/DmEsYMCyEAYpiocCKYLCvVyUH7rQML7sVfiNAvRw+JCDP8nSwQO
EOiJUuoeci03GTmX33IjDjBw+I9ORM1eaqFfLGHs9vn1Vw00N5zk8b50YRCT/sBr
sncC78IAaARVo6JLgeYaOOWWnWxq7sSu2ZSF4t/CTZoU3JFGWx3IL5pfCP6FPH8m
PXjs0EivxDMN3YLzHxf0nJTEkbXrgT5c1D122SJsFXenuVKCCIJcVBSr98TacEmF
TPLr/5j6dAJvC8dNink3/upofE9QaOrgr5L8giug1aIk8IS1+Y+Bg30vCzvcjozZ
B451AnW6I7Fdzk4iupkMvRfb2E04glYJLlohgj30McFQE7bs490Rq3F4elgkAtzk
H0Dhusu9cgoDQqes0WoBKJYmZDPzBSEQlFfhQQgjHEKl/QyhyJgbXtEZqIxv52+X
N3OBZZOVEyQDosqey4kuHmcVTzuyZBc+R6ypV/I+Wf7wYq1kVzzVNRP414WvUagE
EicUuk4w409I1sXQ1me5C0EblgsmjLjmUTrpj6bXH2/EKYH1HwDb1o6wC9kKZ3WA
vWy4TASCQPb2ZRqf3zWEWYteQ3g6AS7qRBvs4HT1l7OIoSrkMOikhRQKPBrORj3T
wGawGQroPjwmKxQmWYrzXoHDeKD1sWINvP9sBryWKEPD1nsoafq1o9btClbKQTzE
q7m3B42DYPQhXBrja5EF/jvl9I5rwdN/AxQGtW2mCXFgdbLjuFbUInu4r5jta8gu
8qZsSD4NVpIp5SjGjgG2ZmyFwWbdFjXpYuAMiTChQUAB/NNwJnpiGpR5nTe1nsPY
airUOi/qNtiG9QWgtCLMiEByByAnP5xnPTHLqF8M3hjP+KiQcSEgJ7yTN2JTbkka
O22FY99QjsBofSrG3qvzeyWtmx9IXoELmaVwta9Lus/JsYn4nFNa3P3aAAJWSD6p
Qk88bgUFHYu7bwNImbrljnQVvCDOZk/GdA7MsONzMgrzDUzoQcDibzAC9m3GZ+T+
PpG+59GJjRQNmbHPR18N/Mko6BUjFg9U+YajhoH6Ll6jL/gwpla80UZ2EhJaA9/S
L0ZDDEeHWa+cQ8Tj6kmG6hbzTHVG5LMtvhgsUVG3dbKQnho8WetawPFvPYM5NbeY
5xMT/nU7xb9K0YRe+2iZGIgFNidsq9sPNrFV6RWrqvuwHbriyzqa29Fd5QuCqe3A
ozIPHOoj58BfnbytddvDS1q26qXPTfK+vPZRG7lIjzbjliElpljPU1rSCNoc6n0y
8oN25O5m2n+iEdWgoipINqNcHD51p8pK79QLpkCCSrR+vbkQ8ivUyu4q61AwbY1F
5TsIEwwJ/T5xcq4MHg9jIGB1RC8nDTYtIuIwhXQoot/DEBatJwvtdF16HJ2P/OfI
IPXzptALaw0GKxeP6auOJWBLgP1zcTCeJhRhcgC+CneoRtWLIWXiyEioKISOOldd
BJDqTI7jF0Q/kv0E5sYESJkJfSUPpGs8r7SdvuE0KYVywJtIMiTEPEqz7L7IP7aT
2Vnm+jVlh92kAeMPUHc0nkXF5lnHGTCKauXY/YzQwcTspqin+od0ynxX8A7ifkhh
evCGsoDgBP703OJVsEBOnHNvFVRo9oV6up7k0MBpe/d8nLxY4/3SZxlroFG5o804
nr8GurIQQxj8gdGToqaC+5mQED7wU6QZ2DrBzyU74diZD7FzfeHSdYoIW/WwwO15
BTyXxNPRhfhALmN5mBiD0zIWnOqNZpzdTJcUit7dWM5d3PoDaoc3REenciW40urx
8nAZ9j1mXSsoOsc/6uuxuUZ93CLCRdZjNqUJrEqPq+TEZBmcNHE/xds3xjH5Roa8
X0M8EidRQoRz2uWMPX4SI4EANzRRgjHuc8xjuMFsWqVcdLy5Wzrb0vU/qKM9OLlv
08o7VqNJKXC1G4J/s7uR/88CM8RIle5G1u2YMfeLvftjBJxbQ2Aas+rzmIsMZr/U
TUMl7EcASrBGLkhSlhiv/DaPZO6VpBGcyQGPZsqmTI+hNqt7f8VBgNsUT+li4x7b
I+pPWbvxk2FVgEdrv489YFdILOlrONZ26D1h4OkbPha7U4nrJQ5nOKq3iCbgzV9a
WO0hvKhSeDfHO7b9ggD5RoePrfIjMtqISIWcXSAaVZkoKi5pdhn08p1qehbLJTx/
SK6bnACxeboTvpUy/H0lTd8ks7uQfng4ijMf5GOewEqirl2SQzJmb5uZrz4yqSNN
g6E7y2SZ6Y0K+i6aZ05kr3mXvhZdB5y2nlN475FvgFM3a/gdDteUOlvOThCAT7/8
UgUw8+DGRp0yV+W6RO4Wp1h9MzEplQna7dxDyIiVXqe2RD+HR6hnMU2DpjrqBA1r
0CEyVF2enF5XAHWkwhlFhN29duJ3McIbMj/WaHYfcnH0xWs/ZpSeMjekMVhLS2vL
bk5zHSvLoiX8pqOw1EMyzPJY945hZHiCGg3CboKH0X1naN1fEaCXTEhxvYQtk2tE
GdIO0rsGxc7h5hh/ROTQDXb/MPv0okCqjcsL74O205aq7W9SYTdRW7yUEftHxpmb
dQWP5SYKm4TUx89IBh+uj2FZtFHOgAVANTjuwrsiiBoTLeV926Ia8265UOcPpDxC
Xj+zivAQ9dPwDguoItsiFN2PjuQpk4h1z8z7WZYuvMyJkpTWMJEZb1N8Gm9UB0Sy
5kw5Z0y23wTVcmYWJXTCEi/fLquaPq892pO3cucpxQ6pVRLh1eegbqb10huDSAJi
pU0vXhyxRcoqhalxXOG6nFnT94RnkEZ2EC4p8Tzbl5te/sEOco6km3tth1S80etk
3FnofwlVs3jB3OqZe72yFw==
`protect END_PROTECTED
