`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2EdfXGbbvej5p/G8DbFIcTQBGH1zahl8w8AUBgrexsUEjFrmbfHAUaVqcVSbsnHR
wCiSTdKeVgHw2yK9uhzpiNmzyK+941uD4VOhDnHfeBleLcLLU2YiupQP0Lobos+s
nNcXOT3ssmYqT4/xlxmV+91BnPpot4O5dU4O4BO2D0BWvE4Y9E2HHsjne1XD7qBh
+kmBGk8ddOvUQZqsxIVEPg==
`protect END_PROTECTED
