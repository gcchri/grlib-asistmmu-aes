`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7YIJYvDL4Eumgg1u1KWoxJl4Vn+l8RHkpxYD304hLuYDycxsHrhj6TD2ndqRFiB
AlhotezIPeBHr9eE9SGC+6cp8WMFZeMb8H0tGEi6hDOTVqOOgA5VhCHssU5GCCig
hpb0bqOXQgEkZd/nqLdUUWBuPLKUoaAMqu0N40SLWNP4Kcn4fA3nAe3H+Rjda4+E
2whcZTOQxMOzz2XWmb9skFFTb1+puGQ8NFy+53VEmHZNKP3XSUmr4AIweP1kK3j6
aEX984lSAqAu+mnNbUy/XStyvMWNKIzVLOjkEZM24u/FCI6HylggHsvAMXMROmZG
LMzzydtaoiqsQatzMvDm0Q==
`protect END_PROTECTED
