`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ek2DxRf9sHLUr/YFtaThd/82+n6jbr/TA1W9YWdcliuzbAvrqoB2dDtPOBmOxmWY
L9e3ABDUKOWfwcHaO0jG80nypjroz8E6jgGByO7jCz//Bq5bk0nUjTeV8sqT7Gth
fTF43+iComJGL5RCAHfwTChl97qUFSvbk2MH1CR91vgTxKSTi6XN3wxUbQOdtH+X
583/P9ESa0lT2YYL2TS5bgbEhLpDr38pnRf86QjtCJ0vCDoit5AC7aQatk5ILbVq
ESOvE7hif562H5CXCSufABmKfDSG67/WM/b+02knXl2nai6FXAH3EHahqIckq0Kq
2/kd3m5K9B//tSawL3NVZ5mgJbPXBLbEPPvzB6bj4pFQTV3Wkrel/+ygoP7HavuW
bYPrz4nekgDnHrsgTK7lMiyYjfIMS4CNLOoxYU8G1eW75j1SZ6ClEDjXoWRwSFW2
EAtoAgFoEM0tD4Xnn+X5k6MgnXIkXFt3eEFBeze6fTUJWKsHivOJ4VxuXIK7zZXa
Bv9opDsW6lTajRAvqkLEXkhNqfjf6CSTsl8LXKk6mNApbO0YqVAEXoYamOwA3V1w
ThJHKofydiBfCWMDJV4S/0sI+tmcpY3bs5VvGSKfjo5OCG+eqG/DdRhJxim3H9cb
o44poc8FlgXUL2IX0VSLcuHSzRLgfHP6ZZF6An1RSkGiVJDCZyyJ9LCwiy7VOH3d
`protect END_PROTECTED
