`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D9yF5BtpO4AeNbswxkR0B0fUnEXmJnxd/Zkz7mOYFqT9D0oYKEjiSzXcSE+taqXb
pkZ5qCCfp5G11pLvG5kRoftmnbpvOb05xP1tEDzOGpFSGOO17kUvyo/ty4KQdeJY
WYWM3L+fmkgc9L2VgBomD665hPcXZmqLnS8DdQdQGuL8PYjBB+EfRdepXooCGHK0
hc6CZI5e67dJYYj/NTBAAI6+pv9P7Bk4c+fy0PpoI4f8od0tbBMAnM40J3qx67Mv
zz+XeOjlm+rTx0CoXHe0p3qPZU4nIenlQttXMMbwGYGAg5B/AhrOMyxAL//N9eOp
qATSrDyfhAk3hnyhvdIJdmqxeFDaFYVzAI0AR3eBUHkCzNMcFb7SPz/skQTjwUw7
hXF5bsbEZYhFiknUbupTo9TkHJAUq/FsSn9Qo86gVWLhEpGEdoNlZwDZe9gzfTCw
HiA4oX7xV2A2a8sHIApQygKg+56ZfOZFhzYegRa0nZR6Vyv6bmcXSxq2+IICaV90
`protect END_PROTECTED
