`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqMypTDBuHvBySlrNM4qKRvKL9/U6iBCGum6aYN0xXG/rRjHGfyvTTBhiSLA95JN
Baue96fdkSv5d/cjR16LEgczhz8AS91UYYUT1XH0qC0jyVMgT83DMDV/ezi1JNjI
t+qYdDR6X4z/wqBbtUVvq/6OnvXE5wX0uZ07/0CYvp5Ikj0L2NKP8h+rGWipQ7Yy
C5jK8GAEBOTOeWzj32TuF71qGHnwOBJFEOZYNHRfNnH2Ja9qEfI0ty2liZ9gd9iH
UnKfdv073FTGwuY1u6Mkc1Stp+eulDh94/ZSLp/w3E3BncVlAQWozwIIwkPNiC70
5LnRvH1DzsmQOIq+CfAy6fRY5xcXXsA4pUJ/OkdxzRMzaTlaNrAf324nSvnmlHlz
M2XHZRElv5/hGQgjaQWJmU2k3ffiC2U0UBxtPhgo6xdu0MMYBzeB+ExB+AT+HAY3
ycu2/5oMwr+Hibit2Ot41RIWF9c21tPETZAjH7aNNVZ8BaP1+O34ELjanZRVns4X
HzOtVn0CkbmZJnYXnny0JyJOB2ZfOKtclATUymO8SFzT+YPg/zDzaVvca4oLD7mM
SWaevIXXSW79maOekpz65d7Yyj9bE2hVlPUvQxSxaPCiliU3q5kmGBI/d1qTZXbB
1yHGlKtI+vnBrdlmcfjF45xpVLwYbUORePHvjf+RyP+G0cORUnQWmj91WnR3nAO1
`protect END_PROTECTED
