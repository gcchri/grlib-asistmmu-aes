`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRybwWfCfdiCguA3cmIiaa9fgXjHyxfKimAUiWBNYFtdE0ow3EL0qKATIvVMZTae
IkgKpk/lf6TxcMEfRVot8NKMbUC5aSeJjjq+LHUwLU1SsskUS88BtRAUNaAd/ytI
sOToddOucUxt6vrIauIPvyroOy5ECjc8XjLDD+JbV+NVvT6UD2a94xRc/6Wd8VLx
ySRQqiwmUnwxqdsFCOdQULJDeB7yv9A4Kypaj0qqPqEnSqUAFZwYWnW9SEzczKrw
8hmR/IDxrffFsDWq8/wHqcVlyNegJzGk5p4BCPLxEgUwiGprlU+9AmnnMS/4hxov
qSixceHg4f5CQ4CaoXj3bJ1Y0IKe6B1PBMtpVEnv4Ln+mOVkLpkOBL7xlYzThVuk
CgmWBIIzU0RALnX/RQ+HXdFAXnO02PkjuzWqbyu6dR19GN0x4w0yReUioAmB4hQ0
mZzGrvrdD1HzsRl33sBZtoHFIPZ+I34CS/IsNkOMcXFW+AIv5iUYSxfmQ/S8K71o
GyzzSLCIKnUCrh1+6s2rQ/z0tSfOzPPEp+GuD53XpbuEw4nowvvo3dzWvIft9J3V
`protect END_PROTECTED
