`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KoEQKH3y83Fd9QmPEdbjJ7b1fB+xfPwjCJC6IRDo1A3eL4ha5dri6tNs6G+ns++b
of3noPNw3SHE/sX/9dxhJZt6T9ZPPwC/nGU7piWaq5L12Bjc0/JqkTVlsMjfX30y
Zag10uRud09MtIrod45JsSXJzZxRRZYosYqMGp5m74iAAKCjQSt7WhQosS+7sRT0
/RvKN41YrRaJEomasT9d3ZhzWroAop9Spi4EW5l+QlSky5MqRhyBSX2xtt16KfAq
i/dneNn7AFRaCb3aablYjG/CDnyKgePREYPQq4NrM6P4BxZlaJs4pq0qq7NqiRg/
YLObw118FxeWbtkXnbCKpw9HNdG+fqi2A3y6cp7+t6nSdetuWZfQMWUhK9hKVABG
ISz+kVK9O1tTwDiEZm+mj6hbzZtlB+ZEHIuZWoRoHE7zECWazVgiOsIiz1LUu5LY
B21MWGjRMpne7Axpm0+LAo8uC9gEMVFKaNkljjyGm6+zc9g3hDqH9kovLgrq1ZeD
ohMgkoHCoIbIkGbECC300w==
`protect END_PROTECTED
