`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMc5x7ipWXh0SzUA7uhpW33Fvn5MRJhlVB65iVRcf7LNvnUBXVzHcR8LfuOSK+Sl
FynSMWgBsrwbGV4qllQBJTsZKY/bblWs8URaPzc6y/QCbxWx54FdTNwVhganYV8v
sDU/FIGi9aeerxNFLGgdjsvPvHNIhdpKLGPtTIFZV5UqTGguG21PiBi/EF6g4t7o
O3dtKQgkfqQ+AE/jOQdEWu7ohaS8vT84MOx5xP7GwdkqfM6ABNFa0FDvvgETEBlr
qMy3ebfW5DaqAJhO8/1tJrPEg/nsFIlYcUFbnjVf/ITw2+0XavWYWj9FCal5eLw1
QGe1+Ch/qTnFWOqqF5fdDe5gfAv66Dzx932vGZEAL8hEbPEWrzgf8VOExoTuP5YB
GKIzEXchon0Vl7GxCNqupYhxajEwx9rwxAIa7fO/XY069bDqvFTWn+4iIg+5Hc1O
jkDSM9BmGa0x4dgVwO4ANemnJ7d4O+Px5fIn9AfMSVhjwkJAT8E3XGpmSFcOLv05
T6ngDTnorv5XhKZGuPbob+neE6H1tu9h6RX1gMgP2+QmXhYJe6NbTwa37T3wLMBw
J46JdedHfLpXgtqzahMsaOmBD/QxIfighy5xf0jk6Fp1W+8iujN9LXoK2XsoNOAF
c0wiJVg4mN/KxT/N1ACaxuNxbpTIj76qhhwuIWY10D2cE42iBXOFY7nGnfmz+BRm
oWNlPykiR5pv3zvRsdzhndPAca1GAI7JGRj3reb78gG8l1C1pLV83OO6N0LzvZMF
4TEG3JTM6s8rXLaasKO2hKoo98GhrzEqux3JNNnwpL6GsYWAwF0vPQDMJwM7Yo/F
jGnNvoyb9SFxoX6blrcU6kokXHhWbwgpqGGcdJ25+Z/+DjI9NEqa3niqgDgbLDHJ
JxPF1iux0109SWl69Z+RITPGEUWyO1lE2fvuGCsDhQNDPm8V5Y+q7C8Z7lQ4W3QW
0G14DgZ7+Ev5tLJTR1G/QIPkvgspjOfvKXY/njV6eJQh+BExVsQjhQtqenXIgrXv
a73iQOP9ACU7h1hptQ4KiW3x2i9x/Xlp6/cI57ZLaCIbAzH90AiXQabng+WsN0hs
0QaPZAdVagqbLEKpOSaXqzmwy3J0fGoLMG0ckOw5vIm2QG58vsDStw35HKGdWqSo
7XQ99g0KW9kdWVesiI+X62l837lI1yxDMjIQ5ZPWhDrjwdiFvxREHgnFE03bBqY5
7yGyiNPuXvUdkJP5vkgxu7pX8Z3b6s1/a945ndbkjOWMJOcp/fbo9jR2BAEy59wt
iC6DhkTYM6t+jBrf7SJeEKPQOntwKIx2lo40c+DEukRAeAg1a0cI1k8oSNqumXR1
x/Zngri5oxTKHpXfreUtkNAn0pFMmarcMqljlB15ZPr5w0tFHWNqSkhjyM0XqGoo
O2KRPSycCZNk4WXhNQ+eaStKbUiIwNbyJXe7Imrzie2J9vQHAuYFHIhjvUh/pIgb
VFzLYsxogJFzuAsiwcGTv3e9bNCv7b7KAOmutAJWeKZshG0BSnbhTytO9FRviteI
1dSzv+Z2c74talclFhXExnPD+cdOMggFhBPP7rnAkxFT5ovQj4oMEBioFLtnkV0f
a3hXL7XI15/mIRgOfojxfxwZXEqDgFFXVrw0CE7SkwBH/zdAA9mDCAISuasn6Ogk
9ZLKDb8wnVoxqAY1TDepirhILPWFaD6FFQdFj6BrDCycQoHo8eQl9xjBiShu7R6U
+vrtLoDvgcd25EMTh9GAz2WexJZju9JlTMjWXVRSukU+bkpyJI3av8oRopZqGvHv
Ruk2AjbtbW1r3+I8cLCySrcnRlqjCmQjP0tf+k8/DqMRIUfHZukiAuzEO7gQeJWU
1SyM8cn+6REc7JYZE1yt9IYgF4NQf6WS9XwGde2Kyg61CwA+mlNmEG0tIVPUvsOT
VrGOs7zG/TQVINwpM0PvF7F2PCv9A/UDsVhJlp+pMtf4MflkQ2zaT+rJrFA59wcq
rspYh6JJSIcm4Q8ZXpILiL0LpgqwW+PdTvtxPnCRfPFVNJ4l4anEC5u3ZRrKdJzw
P/OyrYrUDABvHgvDYyUDS6/7VAY//2X2TkN2C50EWi3jbdl5aFz+eo38INHttzZp
qI5/wuHkNuudhgkMmc1c8REbhFi3o8uhK5dPOlvLi9admoi87uByRrJGjNgATLtF
TYOMPDbpkKPDXEE/hORjy7OeWUXjcydFDbWLJ73fLoT8b+Zyjhk8auLfLdq37YDh
lCB6+WYFFIESEUC1hWJvLBE6YhTLWlE938thnMZ7xYmphdhi3RC7e9+j8ymSzaQf
FSciXLXm8UVww3ixvai6Om3oJRiHGKwPR8Fk7PVxM+v35DoemKZlAm9csn2nuIMM
PnOsif8KSPFEFeHwRdZwpTGG/NSLgaWFHXN2uv6AtN/DRTUx8EafWRgQEksDd679
WmePcq7QePW7j5XGGtTMlXKdS0uXLeSXSwv4u3yVYxBW1V053dAnPEmkdjZADwa8
+ZsPbfBw38rzd+D27BD1fxXIvDMqWs9vupf7CrdGlwHpjv/Sz3Pav1L1PwkSccdt
6wc7xDXnIXqSfpFsJCT6chvxpKT/Ugut0HuEK1NuTdzfiZy0CuC9sXBYU6fnbYXa
hXrpOpCM7TeCNCdS3K3CTjz8/EyK3FvwgMPNpoKHob9VGRsuOuRmpvC10RjvLIws
hUiKkq/0ykJXdTnGM/YyD8EHIQv2nboFAIWkdmBmY7X+3skscmKq/IMF+WzCQ/zM
pSo6U1RL87/f5uMCg2J/g0Op+636VBJXsJEMSCDHbjLuDLWBMcW7uaHbch0VY1PH
Za9HVpzsEYbqwI9E2xnVkg9488InoKoQlMrezCZC8/TEX+eCHKLTTctW8fWq1I/u
I8KA3DkLumt3KQZ1Ud4S8sZiYPOnf5eysc4HVM9e9nIqUhNkTJzpwAS0Odj8cEmt
DhefJnG39hYy2ZmBeeXdb3hSPDzd6XZgp2Vm1TF51K0cSw1gRN+zmhjaI0fDw3WS
iagYTxXME2mOUBguyQj8NhUKapaBd68DJ3w9yRYOTm476CbVrLTqJ78e1SAO9RIS
Uw3Z5UzDP+o2A+sCDtYANGBxoEF2jKhAFi5k8Evmv3c3be7oOedmsl2k4LEsVA0H
s6Mv6NynRwOtbhKABQiBTPDD1kcx0vdDCrD7MoWvYQttgZsHf2sClG0kWEeR/3s+
+rgMzWS/mZKc6clNoaei7KjLEK3Hnbgk0HEhWoAo9skJb45LMf+t4FAuvW+507I9
7cN9cStVNaYIxbp/oFZrtSMVtL/IDFyBEHo5bgmJAAaodon83aFasuQKt/d3AuM+
YtT8p7vyFyVgmCbLhaQ43i+W1PMmV6UpVw0dmRYXs0Tt8luU1sMeEju2QtiyOwAT
272AjwAnRZsf0DjcLMtIygfA9RitmuUbeRjUJpalFi5LKP1sIuoDgqBptEK77B1b
XC7N31lkzlmv4PbH755SpVl+WJ8SujpwW5Kil69+ouPCccx/g3wWhiGccZQyTbY+
VlDSAaUL04yHclKwYQ7Nj29Fe4RWq/IFjWVAF17ddAJD42nzXqv63+icfg6a05he
3LZnBqV2X9ypya6c1r/xX58rbmW91V9mFd5G8BEmq6KtPdNnsnaq1TaHtPRs1ADh
cC2MID7FYTCjaOwEhuPGN2X5vWwaj02ELzz4jGr3dBsf8gjT9wmCRsYiGetxowsu
XM+iE9APxoaXFNwBW9rT7xU2lsBze18/SsdGkGKcfDiaGaTreLbC8DBV/ervZbp3
L0xrVRs6Ad7ygweA7EIV/VIz4X2LeuBn7sb6PHA6sUs2Yhqf+/s7Sie2L7dXWcz6
YF2/y+pGRYrnv4f4sT83JcwiN5qNmdNlaedmp3ewz4MFty+g6MlXpyQAGlL32Ieo
yFAvB1YvCL7o4Gb74PCbVg6jY+btUMhQeUi8WxmJn1nUc28fDD424NHHd5OoL4Du
JCMSZuEZSrs7QpTt+U/lHUdqok8tLL+j3bb/20xctdw1SSytbyMgb4WsAqEEkJzL
xyWKhrGqtxsA8hsqGoP0E5OF6L20iddxamUuSIBSByZwTb+QlRIOp6zh6lxXOBns
/NCtd42alhsEIabTSwbtKwfMGoAO+WIwMkk0gsk1ykbXLo2GiKWdOTBJzfP9Af5m
xmgGyxAEUdUUICsVLh3AJrNDWRJwyYtiLHEQO9tmgXUJxUpz2Qx7Dh8HZnFtphBJ
Ij/G3EXi2/pOmdERSgJOaSoBFCD3OfYnSNt02yLQ32l+wN+F4pksJ7qsOBpFRT4G
GcZAUBOEFtfWOwvWgGgxt6vEaAQGzG8yUiVkF7fNjq2ji768Hbqq2L86q4/UVhCx
w0e/TmAcTPMkbWYR6vmAET/EdHfkjh3wVpc+VJJ/UMQXzJ36npB0zGPC7WORT+YP
LGnu/t2WG4CUa+ubqy3PrsSjO7IgP/x7PJKSwdR0giFBoJYHzMDGkj2rVwxAM7vm
8//7tRfLtflC10IlMrZhGZzjvbzbG9JHL8YKS9YgQ1q5DxVVngb4ncifFqMOYNUp
SU+9/7J6p0dI+vfxyi6g4JTWk9nlzYkPe9sz9fdY53OUh6aRBJkBrCtQRwm7FDFX
XClpTdwAS+WO5HflkGrwcGQEYxiMoUeqqgL8dxvggfL7BV6k6RQqEyTPms0h7Q8O
1a98kBmyMisDCNmxve25hcEgZ4dACGrDIAutzb15QTl4s0MCWOMWynN/kIXxv+Ms
oeSQoh0UbRqcViuJhhaKbgyXFTHK0AP/v3rnN4IQs0QUxpxjOmt8XqyawvS1ajLt
QK8ByBSYLNheNsJ9eMlNMp2RWZ/tRC4QUQAnft8dkfgJ3c8v0PTGb/I1zJsnpOEM
j0fXIk6ygvjsplhR79uuEJwbaErSU64yIt1We4ZMIUuosYVi2Dq++u9kjLbXeenQ
+W1DVyk+Y0nlrnReuxaLJQ==
`protect END_PROTECTED
