`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pqsxob3OurcgfV1IHwVHKjSslJGA6NTP4RkFj/dmVcPceg42eD1b+5/JT3u+zDnT
uiTrwtNxPFn5nIs0KRSNM/p+h0PXIdOu34a+ZgIfStBo6pabL39/sIIbz9jFcdS/
TrjitH3z8iLrunoYZGYPu4dtm+pVrqg7k/fyrzVaGscSXbo56SduuiBxLYemliQO
bB4/QGjgeXjAAgh9M4bb3/NlYY6yvDWuoey05tIl9INVE/Ovz6n9dtshV/4aLA+s
eaWCgl75y4jHkXyJSwjVti9j8HFrvwnF0c/aIxXZbshE+ualDwzkVo3N7jVkx6mb
uEd/sMgmNCjzy/9zDuRYFWRqVPO3Qz8XKc10MQxsyVZw7okgR/8ph2J9pMEWqtoL
gBJe9akES0zp38/0/PjuiPWWEmROcPuv4xbJ5kjPkZuqqwyyMUr/KytVxMnO1+vD
pGiua/hPJcXvTFxqGs7Hh0JrvIJN3brQbh1/eG+UmIMnuI58S6dXcNCENftuPpzk
V/nDsjgOb2ELMa8pRi4IOhZsDHJ7PDhq3iNnHdEsFuZ620afzFVB6yDVPnPxPuVd
09R3FC5mV0eSouPlbe5SFshtjpEZvHVVD+byepJIHHcastQ6R4K+e6KVdMQ/huvC
MZwn82MuZ4x1WLfUMAwdY1sZa4ZoYbuyOckp6eGWg1dUR7gBmp4jYiN7tT6d9blk
HP9srMf6/tDOnHy4jrnyDXXLPSi4m5XGzNifIK9MpnTyzoeIFT4WNRl3AFEmtjGd
g85ej2CKjb0kF7VjU9W7/SM/kM6w8unAYBz5htGhQU/5KPyXIXPx9gg6s8FbKeCE
RQHirgTrH+l9y/a27fQkQRZZJC60RHaI6KI1E9FgbYTrg/xNFzuYsSE1zmvCivRQ
R+V/5mm/hDmJYvewZ0POA4TtrWWKBAirRH1Yv+VBnownUIBo7ZcSi6BA0aqChBLn
KEKwwq9YgIVQnWkMOnX5BRvjQ/rXNxcXVLLicJvtLWbZEO8tcTBVQGECuNHn4Tpz
s4GLrZy31G833vnfVCRiddxKxkeBhS8Tgek8nHic9KJKm43st4BO6RQHrXs0C8fS
xzHhwlD/rB/Wu6EMqdew2q7Rzwuo/GSP3mrZXbCjQBL6ivHoXYh9XaQgC+p46evj
+S3dxtIA/aQ2IARmNps4szqOx5XQd2/hNLDmaXhjI9SGD4korxXqUcII8bH8mJ3G
WurYXVo8SvH3CEWIL4kYGfja1kteo3jfNP2fjMyAPRfSLnY8MPb3oyyNBAvPXV/3
fsGHn6rPDovyObyRxrTz+tB3GJeaOn8Yh5oDbfrzlet9SBAR95dTlmm99yjy1Geu
0hdaaHqMUoz4+LEbzZg9Qe8CUS3xdyhwzoE+s8s/pPPzZsysqMBrFXsFCz8pLtwF
+mJ5tSxEJo7y3oweiHAR2OE9XcCFemJMzatj+RXWUyvidySaNVqSFwiot9ZKMICy
N/U+rW1pGDn5XgU+/eKiUQ==
`protect END_PROTECTED
