`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RMPebAuVjlW6iyTXFV7ONO0g2mbUftQhwGQKn+veH42Eb8IBVGXctp4UCjQWFjO
OkgIimxuApyBgcYIMS/NPwr2BkWnZaPoaI9MCDTLxv4y+6bVSu8ILsypPy8WcFzd
rKNMjuJKJvBmeSazvdnvnu5W+hwWs1ZgjTIOCrcF4xlhnzniHytSj6fIpvSQ7JuU
FDNJS6283puNbR7vitS6Ao2NuDVhhQekLJKgTuQaDszneOfrbSUa3318SKiPz1Kh
kMPTdfda77WcnPBNtGGaiUtW1b5b8HoZk7k4hIVyvVF7QXosNWbPrSc9sPam84kD
Ebt5X7H4ohfxxz3Fd/O+QrHgGalonZUN2y7zFMhEW5JwU8hj2U83hmRN5QkWC1jm
j8WrQuncWFr6jcZsUOA8bm72co5S16sHr6tKXVioVJkOXGjJc5qu/s1iggb3dvch
+4E6wsIyxC2731WlCAog/XqGnKBenDCp5GOS6HaFnzlIaY2yWvIV8A6jprZpc8g8
6JFMkYVtIazgHQIh77uNRjJ39w+j9Xd68UH6+rJuhN35ZlQ2Ue8JzS2zjuZiCSZG
+bn81stluKeUxlKQqaIMWgES11CYyP0ak0SczUct9FA=
`protect END_PROTECTED
