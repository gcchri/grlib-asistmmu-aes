`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RjIRJJKJvE0kgVWvKUWpUgvl8hHnP0yAPoj5eAWqsopFwQ5rDhJaKWd0A7fNj78q
b6owbyKQRSq6F65+VclCOLyIb4U4xaBZ5KtTvgJ+4QtTWP3xHHpuNZ2CaudZNFUJ
LweC0/LOlBoP+zrSKxGLlZ692IYQEf2AS38N+ND43trqSnPGtsF8hi+ACVRfZIka
u7fEHBjNGrTMhPKWDVUGmbXxLm1y+mHutCQ0ch+CTdIHtGrqaosyJSpfQjm/rBAz
5WbICyCmPCdGGgCmbvDRSqLGBAp9cqSB3dlNTe0sh00ZFnDI0nHNWHUVleODbz3E
BmZYVRbZ+Z4SMVe8Zqai5oHGqAjBE44Gpcesh/+qoSI2ZU1WamEglOUJhb3qWBUO
uUyLUuI5YzDniqFc0VmurI1rI1rk56hXHrbg4doWFhzP5fUA3WZVa6k6OwBRPrZ6
Y3sTM9GI7ysnp/N3EXptagHsSUDtguntObbrWlxl8DBVcE5JDT8wctoashhYiXoL
6IHcNZyQXcOdQNfke7xYTFeq/N2gWc3Me/ACtTjLrf0=
`protect END_PROTECTED
