`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70eG5TbyWtrwI+cP/5WRzWfIEItNbpjIdhMXW3AzpDE6nJb/E+Fp8ECppihTsHzi
7OtcsxttrWW0Snljf2DwQyQdrkakZjMqfxx/2e5/ZXhFfCBE/GcUxSyss8WVEzlV
fVnvInxYcYt04Sn53eWXXrVVHsMYDDWtzNsdh7V9kPo/2/Hayl1WDXY0/0t5d8wx
HQY4c38KjEjrHc19+KpdoF+Cmmfa1iaymP7Ep9U6ZwHeb+SbOMmqQpK1pzn6bUTn
SvCGszAIZEt/wpTHBwc0T1HgfcBBedwj4WbreypTBWrL+/zGKiVUN2N7h725C3C8
jc0eUaG3VCObQzX/yu1kcpySGivJ1tjpqEbZlV0s1TZltjpHw3Sbhjr7NIvyvzaK
fDBtJv1piq8t65l0JEQ/fxOyXc3vz8gLK0OVZ1ZILPG9yiuiwPj4ZKuSt4BADxx4
`protect END_PROTECTED
