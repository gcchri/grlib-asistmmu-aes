`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oFk42jVGCubbtuXU8qyVgGugKEgvcz07CQ4TwjxEBcXG28xJi6zAoCSg8FqJ8DQm
/E3X7tm/QND28tgIg44Z1QkuOeqLQm+/5jqkLZGuhpEw046Ll1MvlZkVKuSzA/fR
ULhBqWABXlAjLsukCNQhsj3Cpl/L07REN7KnZF/MJrqasx2T0qVWGwp2VG6cfUUr
ibWsyiaRCeQNufIWCFm9y3wHTXkc9kd4Duc50h00MV6HlKFIljqLl3VG2GZssK2Q
8XA5/BTK88KnkOuEYkxAdI5NaI3NsPkEzjVdmBepPDkCnYfEi/nr8Hvnf4XyC8Gi
OFXWpYsWNaycGHexRkYHN9pXQtXJoa+PFJpxNHiF0r7xCJaRsjHmPTDYB8WzEJum
ZYmvYtQ0+oW74dGWfmwpGIX6wa6izaohibxpKnPfTF51DGkkBJHZuQ6V7xp50kph
jPNJQO0CCC/EtskcBAqWTD10BSEyMwrezux/F8or+FHybeGPKI7FTO2B3v/5QEd7
GLMxr6KWjcCe0hkSopNa1Exz+A/GIzS4xiJBznZ1hdD9jXDyF/Zl/9J7FSbqKeBD
5WXgmIQ3DY0BSG2Zo2s0d7OeSNvFrpgsuZMcw0ICZllLEoW4nt1W/2OpFzb1RWEE
oSIWXL8rO2WWpGRdOf7Tx3ww4f4BcFtDvK7HJ6qwB7koB5sZ5VZ6+nY5rO1L1z8j
7bA1ag5jnorwWu7ACk5KZNGfJ1p8834D24V59UACeQngpvek6kx+Mh7fQDHBCrlC
+22QsiIZuFoXOcRgrTzxeo8XS3Lf0VOrlP4N75Pjaosv+jdZ1jaiXBQl23xVkhU4
ugJxO2Ivjsjua6Sn6X0618CP2WJAXOkuvHcuFt8MdtyDWkztw/oJgxdfniVBuyRj
SqxW3oTF5Q7xUAMhFobyKD2ZgcPxQW7p4Nj+3eUggumKEUO3AWYRh0WonuLWuNwH
eE3dszCZ/S2X2nn6N1Sfc+KvYBBXp4UFxY6o6xO8XUsmui4yUYaNxkLz8ZKCyZ56
YhS1X0yfcKbDrYBBAN/PbrPRPIEaMaqg1y2CNO/71NrTxLhwEEgSL9nqKQIQknLn
48y0WKbJ1Pz/3BvwZtRpmhcE7PW1JAQshsUf4c6x+o+H61g2rr0Wp5W4oC9FCWTL
OkGPzu4tIKPXD9EWXZ1Y8YekoR+ZYT5EOn+SL74x/eWkD2DwUxA1DU6ead6KDuhZ
766yaMBSYVhzOypoyyNZf3eX3bEpOytGnb/lz1xNSX1pRpvVfoekWigKtfskdp1u
MkCyOAU04ACYg9kXKy058NdMRDreJCcgujEpLzyaVhfSnRZS1zOF2qxOZBO7npLS
u8kCWo3U00zyTcgc82hcHVtUQL+L3hBM/kiuGz6pmK+//uHyc1mVVU6vYSeud3EN
9qfMcjTDmLA4GEYLP8qBbARjn00e8j6XppAEqeM1MawjlKDntg99v9Uil8i5JJgA
tYsuS9nDEE+cWNr6VlOBPXkMToeQSSTgI7W9CxXfGMo/5B0tW9HfU1C96lO2IJcu
R+aY1xZWayI6Y2bzxMVbhSoAqVD602hMa0W5uR+N19bOyCV3ngtvBJxfNu9zg73v
HeC4ALzBN54kBTN1MgSNS9bb4COfiwOIrhNdfPjSo3XLV7hl7RVuz48LRn4H30AO
01Crs3oCcEe2q9mHZB8ghYNWWTLeScWNKrBh3hTSzMXoidHXTOfWKFo4b7AL8kK2
8ijus8ZvSl40CSvvPdga5i3/XWX61n67FLAqwGqTKs4xwRKcL/yJ0Ia+x2AdSrPM
CGmmPSnVmCyk5QvG7XJf3Y9Wx3ZiU8k6iB48ixzJWW+iqzE+m+0vLvkuW0p2Wojw
D3X0es8kb7p8O6w4w6tOaekBXl767mObfoAwneZ6zUa5IFx22PeC6eP+L74Gw+4K
XrRC/MtTXQeunFX0e9M+VIwtJwrV/vyIZt9S8Dn+mlS7w2g4SKtWBlHXU6fai/jg
kJs+nV6rC8uvVmnmAsred4ImSZ1zzKqNuL9Yk4138IXplxNWsIcEd7O+xPWCJttI
13bHx5X6BWoWVZZoSZZXYAwG3aKiD3XA/VB8D0rexITNQUwTbmDWVxCvWl9XFv9o
IWPyrSgkDYl0TzKzCW6wiRO2rwRKEJhFFGrZkxARuRCFhJKuBeJ+bSseqLFAO9iz
ubg/XTQEBcEJtDKP6so6AnKHrQnKMwgQ21XZN8FYWKsqnpButWFCN+fxFUGfBxC5
tTqPY/OEUrS4ndzFScl0awi9i8ZgNv2YeiygeQ87VwlP9WtsG+EgHS2J2zcporZI
o1TV8PH/hW1aXZRDFlYfyFTW0CA5h1QNeIx5mjZDFFdpMdqUMDmIzb2O7F+SmqSX
uuNWxMEiWW58U9G2aSK5K3ri/BVdD1nkmXPa/Ptlyyy+YB1ZtxOcdjs8P6a5xxP6
76MSbiTbuAZThMMDE7gpzxFJmHyOvL/ygzbw7zGjMTGnrxnU7a99iTxS8GruJBDp
sgfyeIE7SmZJJ4nkfhVEl4VWG2izEz+fQTO3YCM8fmZL6llF5wMyPyn8j3j1HTS9
Fzl+fSh/WobHM5JMJ3XT8cImTJGmdp+2ielN0pFKNwAt0IfjE1k49m7SSnhlBaTC
6TMPmSbaq/FrNeJAAPL4H6ip29IPD2Ssvr8Qk3olhEbPP9WOemMtQCwWITn7VRPl
m9Ps4I4Dmd79C88xRds/vyAiaWgPpuqiq1RxCt928Zft0CzIliZTdDQgm6D1Oi7H
LtiVJ1jqVWIclN6JLYotzXBJRZHkpoKp4xjsD5Cyv7VaZ1ahuM5A7W6myAONq/NL
VmcvSNDkK99QkdC5jd9Oy2/gf7XmcWutHAMr1u78uWxqoWJFMHNIG1Ypwa0DRtM8
+ti6lQtTyfSxKoPVqcol1Wv5Y4HHI+lqwMtPXD8DlN5J7+gISGvszYsrkfG4T4XK
WOFOg44R4AMwSzFWoBdYdxSJxr8NosEQQNiJr4Gnv7XLMsaXsbp9wrS6ZXJM1EQv
ew6WVVt8WWma5hHFGibN/GAVSRjwzWC/UXoKCgnPEjiX8sQJ2L7oEBdXl4B0Er4x
qpOXihmVy/qLWwHiVrz4Xeb6rcoks/6x8sHI5CXciVF+yUsJGHd1gdh9R5wwsFER
Q/bhOuw3mxBOctpGHJDqnj06QQ5WXIrGjjyk46d3gQgB0xacF0QKmzd+pAjg2Q1D
MXXJvo/7vdkJFpqxZ5DsBvfBKMCgBwsXhupTJAb3Vz/Ec6BDl/HfmMztt2L31F46
vfOwJqoFf2D+vdX/yQB6Jw7qsIsuJC5iFFj2XwWRZy3zJO3/VrgvtyHGfFAcPWR5
Ia0X6oE4hanJ4hlZ5XIGG1W0enbE0jcNzpZfqlBxXcp7JFED69/oaS8MdzqoGwMF
PMEcjU+6xH+aJM80wy4Mq7Z7htgAYxehdCQCwuEKrzkvrzJxgsoJizYFyMRCgaeQ
i7tAFoaLAgit1LQnhz/ooLyHxACAIxTM8FZbVZk/T17KJTIgnqumT9Z3EdrYD9Te
6ykPGJan7e5rhWcKeMrOIVqyExvhlhv9P92grnkDWWk4sye3KLWv2BQVGEtrqQMA
Ue06buM4LI9ZeXrVd1XReaw++uyzjOsgN4nzbfz9FxPhTMuDOBOZUI6ihmvvqokd
cNNIgFwO2WKo4qbYJOAbOMR4ugOPWHWU1a888gA9KRZJjVSMFs4fAYIl8gKSHESk
pxkjc4y9LrANulq5F3VunOqtlSvZpWgddkkbTCNl7vaO3Wv+X7Qg1aiTi8FnEdkB
70qcnFkFztnnD1TebrdjUfBuX+ZolTc8qPviOThC0D/j7IXGDAsD4kRe1hFd0jNz
Vd7TiuvXDLWexP3XrgA27q1FbvsaYfs1VZorP/gD75+bLSxQFz2DvdOuEPsj/4yv
HD8uIfk11fjzrReFtANsbAMgK96eKg+BX/Acn9nXWPHgckRoLMRBaMvQ0H2JTUxU
BWoVmISS/c2JQfRsKusNsyWX5NQItXaVs52gRGknLItqtjtnhBNLngKto4k6U1w4
EyqWocjq8D3efQOpnr0uMCCjEYgKkkE7IYdMFiQ84jiOgW3mTyXspSSZNuEGP75Q
o0FFezMX67N2VtKQ1R714Ajf9c+PvFsr+zaRfu5BHcAGbvdnbH+QKJ4iKZg5WCrV
SdSO3NJs9jqdcZ9J3a2VfXRYDj68Nmi+ux5vqjxjGZnGEMOZGn+lZSfjiw2lf8cs
ZsTHZGdQtByLRS+kCR3d9alueqDOoBzT6ha7UQ+lcoBwaiKuf3H7v+oe93+BR6bN
a6HY5OiV33MjlPdtMvcf5BWRi4LfDCkL7H3sC+mWSdUA2TDi3dfsFfz5yk+OGRkD
2DOsjkr9pCwNbZO4DEUiDbrBmRf1y5W34zccT5zbTp+YznWa455Exw32glTtVI5Y
WtVECuZ8Iuqy6NmXVatvM7pv9P5KgLP8WRfBdE8UJUO3zp+nK4vHBvpnM52UyjBM
VHNPmx2IRSPZwgTrERcQuy100LoMAejZ9nHslCamh2VkLbc62lB8OLE0IXHC1Eb0
XdGzX1K1R2JDRCj5ecTwaBI5kKHAMED3J6i+0kRFAyJc6452wsoUFSo2IayhxLHV
192rlJTOaDotmQe6udlK9Dsl1h+ej7SI87NMA846VZn/K9Mb2qRfMdns0POr6Lh7
uJvF89CINdcgFJFJxsmI4aA5mnKDivOXLErpAbHo0m42cX+UvBiy1XKUJ1qbUkDM
GtBRofr6uHShuWNkvOSTji2P3f4ARXDpwoiqqMMhEQg5yJveFJ4qFD5uxgKCQYiZ
M0Yay9hxUCxy1a6M2e5nyT4Hd21hPVGpMjwNfY1TBM7J48h+ZbRFHq2OZgPw0L0g
LYTV19eR5zsUN/c9+2j7BQEE0eNH5FRvi0EuWMb0GzkLZmvYX3mrxNQClFP5oDVI
mAR5M/VGJQglE9ZpxijcwZZaKHYZMZEnHcuodIkbQ+/JeG3rWySBoTh1VEGnDxNT
pzbV49wHoENeuYOElgJwmQ6VaYghnehKh2An8XdhEMQfPOTSZMWicP4dsH6DRepH
Qw3IOZQogV4WrFAvNN8gQKy1OxYP8qgcRld7UDUNvN6rNMCYqPeFLV8aOp9vjyUY
oQN5f4oHa7lUMH55qvewi2p8l7USdxDmQcF4+dfaaLrOFdH0PNxrlLZ3BiFeAYIL
3DtDsgPJNfTDkGrPwGJuWzSvdG/Dkncwtfn3mzamJIeNMus7mXZy7tn4/nfid4jA
ogeT3VDY70tgFtB2fCDqQC6jRlv7v+dWd3QMPqHpOqvLCYzUR1goqobmx75ZTNO3
jgaHgJRVkm8HUsvxR8JNJ1CR6ypz8osK1cSo6O8aZPt2FfeeKmkuw+k9UzEtF3Y+
gQA4xhjd2E+NL7ei+8zzcUexy46ha/he+/hqxqJ7BUSAWUp94IdHVss0ktsJJ/Gt
CYikLarKyavUUm/uqLWROpYChYb/Dp+Gc/ZkRt1dFuQhnRmm1SOfKwtuKXxzXsBv
P2M1bNv3VVKCk28+RQLyLo+cSpfBYqHtfaFm2yHiv2SBGc6yWfyGLBvJsPOLUUQ/
VdV1OUYC8G+4vQXrWUmN0UUkXfgSnO8SNjLnS8sFODjjzJSvip1K+/3QvMhiNnzU
/7HmBsdhy+cyLPe5LQ0B/12ZngjQiwefrpT5QtRFH7YENkgx8BXMuI1kAkKn7RH7
taZ6tt4jxnFdtQjduZrAYzYiDpEtlDr+SYTGVQyumfXLvqOxHxWj6p2iljO6CwxC
vzeFxTpV5LY0oLSf0YNQr6W81ntEPfwHG07Ku3qX2k/PXaZldccsEHgl5W1tohFt
AkTq9ri7vlrG+r+ssbMthcHdSR/rzYPGl/WG4Xrtc3p1DQBAp+o4Psw/UbNhLU7c
kV5jwO43AYgVnobsx9rwDliHBFK0HLbYD2zaqB6dE2o8Ybw4nQ2rVT/AFxBjJXQe
hX3vUtglMHPIW7dJvhZbS37/IfPQTdvl0mVRasQ8QEX9dh3dRS5waqUHkTAD50jU
7aUolnYv25fGDkcEa6nOJfR86g1UlPH9W06cvpSN1JHP1/Bed5jwWhQAOM2S0a86
hzPbZIYfANcBow9HI0KW05f9D/DEQCqfvXu/qaeGQuVuz3OBsie9xFVJ2jsFrNCd
dcptJrnG77zlHUEnZ4Csp/KVSfmqavNXRN0bDZMIHhA/Cyq3j1aT1fsYl9guV8JI
byKXd+15DjS5Zv2P+3Kp30285PqXGWlGqfcKfTQtvmW5Tir+OekAr3ytP/Pd8PUV
NZxMwPmcYOV8IoY5Dozlo/Mu6laj4zXvodk3LEMwMJgdGBie4TTgCz2sGf6cV3TS
Q1qzykY80jik6XNZ4tS3OgFtS78IbshSSaD+5FA7fHdN/wsTEOkB701G1QbKi7PJ
CgmDh0a37VxgTwMMuK8Umt/jyByJ2uIoaL4XChVhEu/XjktDT733NP8+ZTlBCF5H
WDqvO/yefkMsTstnD54Ad5iz9elsKvpiUiN4kqaNwvNb6T9rNaTW4OTF3tos19pL
qKeQqmpL0OHkEvrpCCQ0bzh2iv1s+DMBPDNcCX2pw8xdsM63jwocfoSt9Rd3bzUH
RYND2qcfCZXtwtoTYGTSnSR6WTFfH/IDqqb9zV3+tuat8F8McJINh6/lGapcRx/V
fevE7PwlmlOqvGGzTVwttNvNucI0FuQ7e9ucHpUiab9WUyrDEsSLGEhILGEh3e7o
LyaoyDIKErZJ3sSkqKUht2yDeF90Aig8TADXiYczbQFngg98xp703voj6aKelVeQ
GxrpcWMlE1Vic+Th45IJR9tdl/VU8NkYDprFJ/sIejfziJP+4u5vDjNoPvRUCPPA
7LC9KFJe8W1Mu3acsue6y0/2T2U9ujJxpew+p3x3s6hmGllXMsJxS2e5l3hDO7gN
77ULXNKeXMyfHN+Xh8EH4moMGYmSVwgM9fGiYdo/zVQTLwRkqmMqsM2eYwGDI9TP
ko7d3PESeGJm9uXZ7Jhx6T0/LW68epKQQ3IIK8FtCASKGU0PAvFJfpN9zYSiCOQv
2eL6mkI5VqhuJFNzJ/rlMQG13YZw4QyHMPu2L/0f8knPh6RjHdIiHgRerxcGlX6w
TczQRzo2SyL5y2UN3n10PneHQdF6rMU7qWxHB1BhR78vQIMpQXRmON40CVnbqOSg
ZZ462bWjreh8kjxJrQu4a/ccFBz/0hbm4/4Y1yXSrkO67jwDB0ggSdiBuZ/NyF4+
nZD55M1WzMvLh8LaoIJVIaFMhoonyUuxzcz130dtEnrXNmCnpVndD4PV5cVGsbtB
wFPCRWsQOvm+xHWW0dTAYcZGAUX6ElLUde53/v3F95ZNuDiYwVt9d6L6BVsrw4Da
kZEluDtEH87VYAJLYGxzdTV46VWxSK5WNFPpxAP37fxdae/t7JJkKnU/htFrcQHX
MUqpKIEQ6lydtTwIZ0odJ1bYI9IdB6d7M3TFMcDIH4VtUdbsbmT+dlvryutm5V6O
FnErX0FelhBkt+zDbvd+R9/Y8wj7uWzynGovQxJWmfLkm3udytn7S90vtzYMLu0x
MuplCLhBx/iqf2pZ2ijTwGcouc/dO1Uo9cqdDkF+I7OiI7N+0zmi6g5uZ6z7ME+v
Y3BFLRIHsUEYdDIUmrvi8/iNPI0a+6sbvmiESnVpMm7Xb11cfTW27o+y+fkBpeeU
ejMZL7OuQDtgtwm1pnYc02peTAouo1n810FPt93XuTXDWwUMAUGfHB7obaF9P7V1
HzN2Cm6F5SKX7hgUor+0tqB79dVsouhWD6TZkbDlj17w4srwu4iC9XPPaODDLR8a
/ZdxXDgVpDTKw8tr9qqN/e/4Ju2DfTWzuBTufebwVK9oGcLhq7TVDhAIaLOakeOL
gShOD1/YgAO2t2qGIxvRX/1lv7/BkuqiwpHs6r0Ph8yCX9JhWxZHQuEt1nJjfFKo
gY6CMFesHjj17nYeFMaS5BKxjkq2ueNDwwzZ2o3z5FfI4VJVjQ1QbdxEIkuEaUcg
dTTegfgzSoOwPemo1As2tggi+eJuc6VbLRg66gx98Do2UB2ktptfGJmcAUpuF+Tc
LDicpyXczNdGMRvVd0oRoAzhpAU5dDMK9Z2KSoYDO7jf9SJiOoLraW9uLYT+1ns9
/LjocLanis3/jzmMXhGDVDgc9rdvhJ2AhqNPykZe/S07P2v/DFqA9BGB8HaipE/N
Gw8TY/z4PIHkW49ufXwqk9tWYmBjn4X4iHH5a8vfDL59IIErKxeVz1lTf25f8G8C
ht+UAKhO8StdWmsLBdyABixOZ6gOKuK0cHHgV/eVUJ3OT+2BrPMgBIseyygK1qZz
khWbAe3m2ALEk1hKsrKZt1dDs77dd3BKdRBqAEJJ7Kv8Rxq9SunKvVIoK1bskv8o
YogDlzh7S0YdxFBHsAILUoA7KSJZxofcKIgA/smrulLjuO7lSLOLoVJTbh2WIPvo
lxscpMOp69o4Whn/ueXu/mDo9tJQugVkaXmFd8AIDvjvbBC6UUn2ZTRsRDFwFJch
3TTMsWDDGWCRVHafJHV9aKIortQvP6GdyNIjRFxQ6G56W2VljYxI7erU0AawmWrT
sKLp+qdHHKDVksaNvwuSoM+VMaBDvQb/u8+5zlod88p0u5WPGyR6VBIJyiUuECvg
9KLbCIvlq5tGZFY+G/RA1jGf/9qzmzZV2M6mqLIOahjQKksIGMGC0QFKU9WwRTYP
27m4ICK4EARtRNvfBX3mGuNzIuqdzL91wHFWegsOnglsKObcl8KlkqGwsYDosQNX
sNhqDlCC3LNTzvsGFpTGzVrBfRRjXD5pcctGqhtAXNNJDkx/9xfCNZlRVRyht8g6
XAoMvM5zXx+JTV37lJZSYcEFMbPdicR/O+EeE1g78JujAk/nB/92VxBzms8i895Y
/WIgg7pQFa/WsiQbMJ4ZjtoewxDQL/NBM69NMBHmzwza2ExP8PpbjXKJRMW9azyG
c8HCupi32n2pW34n1wZ0qIrs5E0mRodjPHGWGQ7nX8L4MaS0W+HJile4DM76Dow7
nvT8XRXGta9kyh41AV/VHwB2DF1nVl8Ibu7I6f51Pgy87aX6uPTovZhPWOOM5OAH
lqyT0ymAupJ/dQWTfhjTNolm4sJdDTdMnIjVUXPOiMwGzUkssk2Mk2AmfFTutYpE
pLVQrLK1JRUhrOqOGrsiBLHTfRqwteSkdCb5kIrREikQLeHvkUvaS6I2IN+nLVLi
b7cJyBusONrNgEVGfTCYjByB61v96D2qj3s6zG3GH8cwMc6aD4eSDuZIY8AM5TKB
G7PopeQPV7XalpCIQmtDEUo8wCBL4x6YAcrezxZjbGB6FIZuyI5XOPMC/euOmrSf
v8Mje3x6AeLPaxyED3fz6MikZT5RUJnYSP2FsIeDAvugk7nxpLRy+kgfkMjjo7Yp
w0PL1bcsQeVD6zS0zVADG+Te94MXTT1im16z/NJ1qKdg4Vv8yC+ok1q7g22/oTYD
51oMsEidkbWwv5eohaSr8TShS2tYpSKf0hs/TY7fuOtQVZUS3RVdW4dSnFBJE0N9
iR0Kj97MZPvN6TizhDP8tklwYqxukP+6FopzXVEASr5rMAnR2+YyhMfSQDrAxj0s
KTanLkkKVs6TNrdVcMJwEzpI8p4zh2OCe8NCpJJ0PERIOF47tP5yt9y+gTvunhbS
F35ax8XRxAj2xoZH+L0Mf9w0R1HzJZM7haKKB6AmJWmHjS7SguXx6S/IJaNLI9gv
737bJVvPNYNLTLnX+fB/tmTEeolF++Du+VZBUYRmz4arbpMhba6uPbHjOJdMxi0X
6bz+TKsl/Uw6Qhsa3zqqybrljVomeeFD3ogfQjJljPOZ+WVaWPGRKYaN9J5dwcq5
BYYn+j7gUBCZBqSwr/k7PVKT5pe2dBobFZn3Wtvs+dqWZ11FwdXMrHTpqW7RgW06
D1tnRSbahHXpxK5Eo+iMQroGkBmiV6+pSSYbPsISFO7/5AVoLmU1UUUx280png6Z
qtSECeyYyNFU+bbXBdD241Q4xK8+dJ0wEiU04yg20+C1lgvj9+/hfLkZAF7qk5k3
O1JlyUHxIEQdHmgzYpG/JndVdvZA6OjzJ4bhtX86F8CNjl+V2kAglMtJ9+BsH2KW
kjlwSFm5eCt8Nl0NjX/xCDlKIrDiSgRUhhCi7I3KBTEvHvxOMgV9NfN4KcZyQHk9
8Mot1GX2QLXXQaijcYZeR63E5lsVuFGTYBpCVkQnie4nA00EIff7dh9WPXzHuOJZ
mkVQ9Pykvnt7YW2+HLto3nSvZh/oIBHSyJ00aBpw3oyAtAIfKBvD9Fj4j3qHL0wU
A42U35OuHQNRm0iadyx+NiubMiAQFF8F0MgaMAotoZi8uUkJNgBcRJJJqJVUaXry
1oKl/1MMyRo/mAxe8qIfnHjH0B1LWM1mXR7r8YLzfV4BxxIosRC02W/anLgOcYf1
DMqmNY27lD3d81KJ72k3/E/5uKpgEoCvznunoaUll7AZoHqPzRK0AK1UpPdOHnip
9ve0vWeeKhQUIIxsZz2CnHBBlJBSexgIv7xcLo3ZJ63VwdxjQIYptEVdqyjDNJoV
cfI51IuAbDCtr6pxLuEQQ2yni1cljdQt2po7gP5HLE2OtyeEQoGM1gcNa8iethmo
LUEK192fxbadTNd03CDHK6TX3LIDkiIbr6YMSh31DvwWlDd+l6LMhPKVtrmSo8hl
gmb18kiFPC6U3KPnmCUHUG4aYlyZs8ZrGdpoCUN9suaQUVTiBVnauOO774lxzxWq
bZ1qrhQQMsHHL7VPGLePQiHCTdUAbF1bdW8CoSoIYumU5blvKYaNYwpwqPXvg8NY
WU4L/7RnE5c0wv0MWPTbsBrL85CHPB9wjB/VEdM8lIfuE4nzcCIhIEtS7p9AU++u
VeP+wLLhpvefKb9IPuy13rTrfKbkmJUDVaPlI6oT+yRNnZ4OqL33iuRVVYuzbOzg
brV3Tp8V+JRf1ccieq4/EhrolxcibI264YDI7TVXdq84ddLZUiG0wk/2cTk6F8S1
ZYe5N6gzrp9ktjUyHGAG9/n5BoLCsHXobQHKsSFcm8hv+xx4Rl+JmTV8IvyXGLw5
IJvkRSoHxIM+mIbSsMIu+fmksvkmpsuqB5Qa/pN+rL7LVyAfkrcrhl6kPUkVbl6C
LFql8vaXqMjB5WHECN30IqIq1kJukEjVJcCV4irH/oOBOFL3m6mZkQW/GyGPhxk+
Kz1YqLBen6WykKqvJD/8fqL+SiCwu46J67BYnQFaZHFO8B9ideaG0Fzldb6v+ZEI
gf1XKP2FXXn3N/2DHBUoohOkZRerJYAb3Ea6O5tlq8PruwDBQB8ITPILSvxHgVIH
Yds/HZBzaUUIiWpc5SXqcZZ4mGKBMMwoXcDwnp/F5MadAtVosJQjGnlcxd1WxBob
tcUiX3D8+qEhw/0Pqsgy/CL1jGLO30CwsAn6+acJswj3T5zS12jmC5+VDBAsRz3E
stSG6SwIVt7PJ4iRp7IZ4qP9AEFGd0xnTq+gOwQ+KWdypnhuEOCGDwEGqwO/7Vtr
NxlZuv0mQ3kGVKgdPKit5ooys5Af/UgIOVsA6oY3sgwFeiPh2imxsIdk4JaldIu1
83vf6YP8eu5KPBVJnSNM6I3qJBhsr4YDPSN5cAEKom7khrbrDkC3rV6zKf7Taaea
jKpG9ssw2HJvjwA9J0KisH6izTsCdx2EOZV39B+aRHVBbWjTmvDI0SgNyPxXRM6T
FguD9PJWUb+hDfHcRO6OHLiPXBzejOnM4PrTwEd+juv0TxFJnsCDtYhiRbR2z0tg
LaBOeqbIU+KW/Vwi94DJDIBLKX9nAt5E3tBAJ7beoOc7ErsJ0v9c14CsxlkVBxF5
Y53PV3L447yiX+kHYEcDJ+iWQl3p4Uhgq2EPdlxj4zSDiWiQqdz+ufSsMJdM/w1H
DvKkAXVZsJiZX+yecQ2FxD+DfJObKbEq8e+kCoqo7YIJfAqjOuv/TjbmGHp2joON
b3qisepD7SydngHsIiU3HJRJ7V/LAc4lgrAD3ZFn3UXeQjBrL4ahsi15PDcJqCqw
2TxTfreTy3sJWw4hNELXd78L9cPLjZ9gc4DCxKmCSlxHCEjI9D0/MoQEKRJrB4Ny
NJ8Z82BmSczq7qvRG9GiVMUR2bcMijgF7MeWuZGFKgNYDdDDApca0GrUTfwKWgH3
uqJB6XA32gMz7Ualx+AH0oLZ8aTvxLmfOXZI3WxnIIFDVpzvLHUFt30F2Q/IQmKK
gyCWd90B9BjNC0BvMaKguA0Sd/+1uWdAaU3EXH3V3DWAga1HsrmLuZBszaImTe+Y
ePHFBP7/EHg3srf9WysGfiY5s4YE1nVWT676UD+ghL6Ggcr9mItN1+8ha+YZVeyz
emlOvZVWwfJQsoYAzxDD/Lg3GkpYkTmgRpM+mcZOTU7dEO51xsYqs4NLUSNmaA7l
kUAqnR1/qjNJIuf7/CEJFnzuigfAEV6FKvY++jaIzfrXLyRO2+WemcIyXIyrJ/Om
U+ynL6PNL4NQqO+xBC8hONVWPkUhKh/L9JNftVskTfTLEreOe2qKG3bde3LpaimV
DGl1r6q4pY5Jsv1UxOBn+EaY0BvEAss6+dZE/jnzDrO+PAmO3VGAHb5XkZ81EchP
OA8s3McP8A1zDlCC2ivq2zW2QGDwBIZwpvKDfuStXK7c9z52Bp2g/A+UQC4Ic2+8
Qogoz+dphftvgXZlXUz8rS2L6g4QpaRUcGwj2VGn+EdShxhC5GarTwat7Ywjvvt8
FkogmohSWdxLgP6qht/5FlxM/24uw4oJIV21wOXNSvct6v7KO97PvKC+lqs9VN3d
yhZ1GHRsAtBV0ByYlMxN6LyVZcYyyVZj0oN+sKuerWqkP4vWDehnDh34DcEXxOKz
qMgrILwU3335oWSyKNCv4pWtFSo5+G0e569s3ZfdJkI8wPSjq4p+Y+VP031JiUEe
1L0PwEdlR0bRakLr5zdpVyf0uWy6unKcAczrXbpnfkC5Vni9Fu1phgheMxg3Iapu
FRSTZB9c3d+TnpUxSFXcyls+3p3OTuDN5NLGuM/xSjUcJE6G47g9w6QtXg9xEaMs
4sJSd7xBqetbBix3svL1vjlxTcRNYmm7QSt/HVmHP/nrc7WZVpvPELKW2wH0LBs+
Oda13FnVjl1125Y0sdqO9YndBsFDXl5taWWu5YT2MbgAoC3hzrHjGktmiwsxQN+L
6Kyzbeq3YqUAJgAfXuMPEMhrKbAtwLxoJZblrNJRjc1sJMAlj/PGNF7aNbNA249c
M1NZg0YoWjfGrB6lA7Ytz/y1mWtIDkS33F14P6vM2Z3cjyeFnu2xk2LXWdRhhB0B
6qwycnF2i0DXQvrL0WK2LOsAjNCOukGkF27JjRgor129GuWKftQqCwVHvSfpFbJN
tHdfJWuBJWYv6A9WUXLF4QXwfZQhJAkaYTGmUJxIS5tRCVGJVTtWsEOPM+10F2Qo
4FNd1QK1KSdPmsZXQdpqr6WvRCO1FYPDPibk7vxDDelJcTLeCZUz5RvbD1ITdVKt
XwKbZ2dZMBU6WbKIAiIsGB+zLXlgxH6z17QO+/WTn4U3q6o96TP3ciJVCr3yxeDp
xV4YDxuEYtj0/fez5gnqUYjgNJyI/r+mwU16l3EJNgG/x9OEoezBOCx4zgg1LSgb
HdP+vdbCWAalW7yzW+hvPvbNTP1TLy2zLpJZai+T9dfIuBXzMY3eP6W6mp9rINqD
ypodngJlz18deEXJWZ3OjGYX0RVHmujzmKw4kEQptWJN0Bhs36nbUnOtA47sujJR
Gq6/5VApg8GYKpk13iOAyW7IwnGTaw34QOTots81nfGA+ccMumfwvl0PM0DJ5psU
Bt18PoDlzd41WgARtm2+alkl7fD1D+tQYx9Eo53jronF5JWlcdxC8KCrQkg2vuTe
1YRIn4iKqYfiURRmGDeQmSRO9E3RzEQs4u0LLQm05ZW9O4vLf493Wjue7vXJdVHs
DN0Tn08r6cY1Lz2LUh4d9fJ0wTW2li3yF/NjddwUIHSkDHp4gRWuxGMLzN1Hf3iN
1bTXyOa5YbFWv1H1uKXqYTQRuSBzVDqX9LdzXVFo8SZ/gvpeb20Wx3GZ5mH0qkOB
kGR0y4JAz6nYDpz1dXN2ThKUB4YkXU4NeqnLwmjlmdOfvQ55wYQeKSTOXuNUYF6I
02i4IKTGrK6hk8iafRhe4p/wgelHnG8SubAbkJyaHAnz+1E7S+iXA9qNSZekU3HD
/WvgUt0wXJIQJ98/15r0JZuaAU+2m4y1OmrANAKX4RMG7a+V8Uq/JVUf+1TQMxKm
9jqsGlyXLaVwEx1zlrHFomV7opa5DdPIokT1yeO4RUZ8YmVZ4rM/tU7lqosnpcW0
ZTDEDj4yIiUaXL8k4WCsI569Sv8dwGDNA6olcTeksGVpgADhzcLPSDj2/8A91dS3
2P9H+9r3Nv8V+qWb+42dv2qV2jAk29CRSsRRD39kTWu4PMQ+fxcJg5TohsBj/IB4
IG0WKF4GvrsigM4Z/iyQNUB7NlhYt1GOJT/okX/2c9reHdWnYEV3FsEBzVGLp/DE
QQ0YskK3xI84nHfGTQ9P6UKRY2jQdK99g/8HBc/Bq2450U4U+aBuzCXF+ysSO3K8
9mK0/lsroKHfMoRIIXOkBHN7iqqvMglRZHEvxOnnsLhUPQjq843dvb2ZiWE40116
Jt3sfZpItoMBIj59iMsKj+5LkKK67k6PAoohx1bEcrQYUxW3AqpFxPF/CVGSBRfR
8lXEKOdmmRrPV2Vk8UJyrJr8O3SEehjBNi9ytr2JrFG+Hn781dboKnR541wvl/Ek
qWS4aHDC1TdNz1wr6YyMZ0ZVqkS5mfx/g6UKObmimIbmNg5o7/xAaLZ/newunfSd
9U0fqRNix+udqFqW64PcyU5aFHBQ/Q/QcBW3MnhNRdAY1jcmx3hemStgy9s0AiBB
yMLf+iKMZ133ERAUsGV16pY7AieMsVL9Ug8VbWW8Rxq8TMJPiq6QStCdCa4/CJVT
ZjTTYUUM2YNO3GjyiCjmKwAwmzZJ0THgoR5FBBhzvVt4t/rK7Sqo6ay3mvjNHW6o
lSOe5+GmrcS0QiQTzMa3LAaWDjzW1leemrxMFfnqSLkiQ0fyFtn6Ig3FNVeipQ4T
G3gsyRJiSsChHUfC7+enmSsuRIGJEoriRuaMq8qu91BXfHJVDTXYzjS28N1JpUYt
+N874lqj5lzx6mG5lXf7ZxB7wgpk5lY9MJiaON2jL5XSgR6QM4Va8EMNS8ECElxw
/BUOhz530sgP+CP1J6lV0f5z+OvyxoP4ZAeY4fbVqaO9f5dpBfLftPocwoIEACqw
T7unC0c6T8wGL5Nx7vEQ7OncPJMCjr94DvoJN4qwAFJPL7iI/glgrAdiA5IazNXM
tEu5ISli8wQKK65WUxUUZ+j7P2zyRb00PBG9Ch7+5e+Gbt6n0oRZKFl3CgWCWbUD
uDTSArV+I051MeP6BHQ2qLp7L3liD7sfGvv5Sb4myOoSPWmQGK+X+YmHmM2izZJr
jumNd9nxy4XsNrrzCwtw4sPgJU3h/+RKSRx4YBzzeK2h/q7ZZmdIJAYf9eBG4ojA
l1y0YzJbTkHD/tay0HAbCrwx4Z830GivI6QkwJMMebIIEpdLaqLDMjcxfl8fZ2Pk
AvCjCFWhnjNrX2lOMCsoxN1bDUhYsqA8dXcL/P0Z/YbR6qIkvvDPEguMBophkBca
dfhhJmIE6J+8mf4MKnlev7bfD3D5/pTHJ9s0txlUvvYeZA7j/emDOcYDd0x0QppY
QpLXjPBd3k9jFV69zbXHwxfRCcVrmEHIQo9kYyiqR/9pbv8AITCn+IhNQ+CX2GuB
7E9SFq0r92UOVQUSTTCapvjIBf8VDpq4vhzIZ6/HBOZPvHQsrG3UjTB7OXoRbfQJ
qgi9F3Nl2dtwqNh2FITqZGiPO8pVhqbpgbDwOidqlUotX7RyVNFECRlEvPT7mobL
6AZOku3mWi/z2W6f2Ky9a1ttkFNt0/+WToDu286EuBpIrQCN7bnf/9Mk8Sqxd5PI
r5XtjjULVi4IqdZ1pxQJewAkFfDBokE+y6WiyVOSM+dDHPTBh6t9RuR6VzFpmfu3
2o9vV1u1d4Ek9L/9OuPwbkIzS/o1Qw5peYHRu2xZReysRKh4M8TiU4ciC0Py4oHv
6GBFIxf38bbdpW99ENsreydJfjYf2EgJbROQBiYN3NV2jq98BvMtkUPLxI4KTJ6G
SYPv6jMsl/SUzxq+YF3HTIm54l7Nlf0uusbLMDbe2JN8Zv3FrAcF2iisX+290bzD
3sia+w4/w8efFvCDofNqXkU/TEtVzFqggibioh25H/8Vv+hOX8iYvZx50lY9JfAO
TU2nBIg/QdwFiOqQ5t6nALv++nLQaqJ5jNXDjHd5vYJrvolwHUpmn8lXFTKA81fn
KtSEFdqmrGex2cjFhSn8AXZCBM2o0PMuwmrkN2/Dw4+lLIfZwL/o/vgPZUkoECeA
n+jhYLsSWrRdckaPfWLXZ5KQI50xy7/NWxqbHeE2uJ3bJQ5HpqL+Qo0l+YT5iUC+
usntIjNrz+IuPQubdsE5bT8q9PuSew8+mmkyOcMA3Phg7W3RN0OUATTbZ1XNWe75
UYz4rmo50wFoSByPkIq5dtAHkUL5OygFc4F4hJLfV4zkY16IN8kROK6ThiIx9pmi
KAVr+9RYVnNtjW4YzOn7EmI/t6Kqrr+4zE7R1i1tj6s7RkCuCRsiyS6UMKuPuVfL
vfNJREF8+lKtj4bZgtEjl1mEfKm2J7xgLYn8KUmQUhQdYREq1VJtVZhCNrnp0p7L
fq58TPOrZEajoMrfHp3FLCDmutQJCZp1VwKBnwVkOJxfrB1SBHgAfCtMV/r6Vm3M
cZ4rB5JZ7AXAN87/jNcxEUCRq4hLx+gcR0k8w5sU/IxXLNrxt4PScmMJK6PrcS4G
R+JjaB1ozvR8xEZW+8eSCDTPAUZRwey6wysjvME67NtTaBfk9fTwgC2MbQ5Uw2Wi
dLReQHC2oTKXp48d8oKMaSutviv3m0RZ8tiMUpZDyFMHhZ/wYTdk0J6K2AXkg6D0
uc9/XxDlocRg5jFznERQgkWQJ1pB6AIJhl0drrROEpjxVNxhD/w0RwNMsHxI29gS
kgkT9JCxP1T7XEUib3AtdfznvFY9ix6u+AdyQHO5Itjj8eeDolgWVCfGKOlj273p
W1xP1OCHj8obQPhZ9170wS/tmj++hkXMH6wTcw2t6GqSwPVRX2aUo3iCpP7BIIP0
/UgFB/9nDofgttUzmjxwwjAMgmaTUwXmUOkvBsb2kzApAtYsUHFBQ+e7xYFyDzAe
gOYT51q25k0HlZXUmxx2S9tWX5p18tcBcjDZbavmjpw8G8pwAq8ZcJXUApJW4U6m
VP8u9T6ukpXIzPYE7jiGHq46ITVSYGlfVAc10sSmfZIUhtD2P6TKkdmIz3SEJMgd
qzS5PBEsl3h6RK029+zVnLqYFEvvdU/NJemkOh6pvgZAAJORDV7m+KzWlAR2e+Du
hRBVtEbmvbqQM3pCgw6kJdr976dVe7uqLwdnAMI2cYfFB/Ly6j2hbAiWL/2ih1TC
fYcYxlb5I2IUvMRUYtoda1QkOgctZpxQH0jstAzBqYQkuXpcpfi5oSbfNCkzKi9+
alksnOw83S9nPS3BLMxGfw8lN9BqIXftlUzJCzkvyZSxAknKzFZ1rppE9sGBKaox
oI7OnIax4HtB+8pNP3eMEuNzSdMYZgxJ0c8u2tWJNAgtTWQwUEvphLlG3TXhjTyQ
6nYOcVDOWU9tZrQsml01JWs07DPqGjXR3AG26sXRUEWVUQ1mWGJ34aDYl1bSYOYh
N2KOXetQrVvNV38gme2ynNGaLrLWIq+n/Yb274wQf57YZFfFMa+bYBulhgCbP34N
ofbOuGBGodicly9/qEwZb6dcjqUQVNVN+sJzsB3GK+ABbd8WQSHx3g2qmZSSATMb
Qm8kLGunacSxyHkimXNQBo04/Nrnnq+2QOvPdBVU+VJud58tsSQy2CO837jrCNnF
f09rPFQUzifOzXu3d+bwzr/U47fbB+ZynkUI6vNFoWeh06PFKCPSEVqUBGHrBggW
LoT9Vxr33IzPTT04bshcxadDTv4oTbUroOCinZ1CtSs12yGEY3Jeo3c+wSSCHj6B
sO7qv8HLvG0bDxYwvE3BaJ4l1YeMWiz/GBYPq0V37LA29Z0HX5WPczlbhVzbMqkL
MMzJyxVwaXqoSAGdPZtAKN7MxVu2QHME9eqN3tZikR1WqHhhEBSFzT+oBCzIPW2i
/LS4ToA9ooRmtDp713MfPCF8C7SnxlPnpi4uh5DPzXDj3FwrFEum5QnUXST1v8sT
6ekBFT+7V6oOzNeINjHFoCU4imtBjAPLucZG7Wvxy/OPOtGb9iQVzvKpG1oz9NPQ
+aZtmQgx1WMK9X1a6HJbISmtI6U40ppd183k6kH2DHIZ+7KgvBtzn7Wk4ndFFa/5
U78d5rReMr7/+2oCj0TswV1YsqX3H6uu5ziwhf073BpEe80pDXl2EBoDga0M0ZVM
2tzglxc40ID+0f8DO7yJQASX2OAIbhWQn48DbHdi23hlYfChNw6/8ReF6Ft4x7B6
Uyx/0uiQO9oXAf0mhUBDy1KmGVRNtwYchIcvJRTukaG0SrjVs0SholQrwxBIdNdX
zHgZYyns0dn0iD7scN095a4ioSGolTk/8n2x4mvK/8aTsmxWTcwz2oERbpI8wQPe
077M3eyZqPKL0aA1vMdzHSWT3l4mDD9gNFv8Nt7mVD9/op3X8FjEuHC7R3BqzsXB
yk8lE3jh43ZaCiFCm6zRNuVmhW8VvuAxCik7wXc8lcdvCLpePutADpWLZtRGgcFY
D/ni1PGw56FXIgz4pktc15jdf3gj/qmgVxLHICSNd4we/Km/AP7WEs1Hy3TFq6ni
VRIwOK/WbQrsYq7+O58MVWAw3BmHyrvo40ePbBn2dJVXIZv3E087gn+gA45QHDRo
4rJzk8knBYpeeKLUrcAAcxX+7Huu+NdjtjxfxzhSPL2FrdI7fMy8P1EmlrfYvoEy
MAa4p2VztUq1vWKOz+EQ6Ck74iNldh4aAxPVZB6wayKAagvdpedaEHp5UxBgI96X
uaDv+0I3WsJ3Oc9A7JRbwT/fenceGNlPWITyXTjxQVycUlhAZ/SlmkwMNauGcC+V
dft9FLAF7+TV2Elzc2C8QKlnM8YTebpDN5CHo2GhWsmnXdZNwVVGD4MW1ASMsPwQ
5AD9BgUcZ4FKEVlAHUTlYhjoNgkzJCTx76Z9JxZw9x29fd1qoDtRPgXVjewmIHw/
cZczTthQWRywxQvFgeTE881DH44B8Cc5QhtI+SuI5lCwfhilDOXiuP+HAF1q5I/g
eul1U19HnrGjwae1mflLc7pGPw4P9JCCiUqpbK3YnsVIl1RyeUFzt31ymuYxjPbw
wDXXU2mckkUzdj6iYYGEL/CYxHI3iS18he76PBTYk6VBjThrjGf4TbRqNdMd7IU8
cjWrM/gZmnHAjvHmQDGgXgVJHMYh7J1cTb7xb9GoTRL9nMgd3m6zoP8oPYcxeG4p
r4f+d6g6ilNqW3zPSu6MgxA5N0FZ8DFmpripbHujQ+sNHH3IdZXaZwLTl/eG+6HO
095Bq59RRkdG0n9uqmnyrONagC1CbkJWo3Qq3eLbUEoFJvZ/oA/5BAdgdgBAW4v6
RIFVq53ik05OLAkoYR4GxFbjsRaS2RDwadReTXCT50EdMwlpYEHQODTaRhjgknrX
atVeY78cHSWMyzmtg02iZQfdLH5SBmpXp1dnUTLJ/0Rbu8+7Bq1p2Ok8jMSJScY+
1a+fxJWKmnBkvTL1u5pUNNevwBbymSrSVkLwVgSZ1JFCGmWdXUkzLu9IldNtbz+M
abxMD86IMhmp4JX/u7j70Do5mn8+mGtYvuUBtu2CrGV2tvyvfQLdTnnGq97AQ/OA
7N77cdcWKCE/8Obv0p/CJAKhWpENnhowvuW0mQglkdpUmKJFE9znRb+IwuP5Ki72
ObnKhV3fMrGCHkO+TrnvMFhLZYmno/QdtE9wP+xG8wRx1ap7Hy8V5SkloqGL8RbN
2Dmy4ZGd6TLPqlBpmANP4ukTcVi5BBuJawVQzaXhpcuXFbR59eJHcOEIU9JITmoD
bJBHk/igb6DC7ib0wodakpjcauFUhVlsPCwdBh8VLkBBW5hvjQqeLFzInlQm57jo
pErFiB2Wbd3cHfVfVtNXaW3uvaz4p0eLzJ0KoCJb2bYsbscmUk8ItRwhXzLHvoor
iF8FuqkQoBRmNaKaI7UhTO/QsfXwGcKSg7tCrKJXgd0sDoZjihOkcY3IXQMH+S87
qnXxp0VqGkTxQNvbjBdes0kaW1f/glpq4YgFvNvAMM1WRWiYbqlJ+Pv3BJmceCCc
wRw+CSyY3QXWP+hSA+2R2J4W4kB99KQ3ji83VNJOwxMnht0qcxgf7BOrL1Vyj8iM
hWqoWPC+FBVCURtdmgwVzNApZYysocK47NQx7OnIkwJqCwVy90rfLkvz59G13Cpl
sNtQthXV8/Rx1XFemp/QTHoLF4S9u3gwFJM/zdZlPyW2kYh213nowuRpIc/HNBnI
0iWSRSaC684qLtmmKTodb4S9V0q9auICym76Ztwir4mF3bvCIQVxY+NXbOr/b4c5
KoynU67bPCxaTU3i62eHwiMMh7/E5jOdd6UzkHdtxXMcLqE3+tA+8SKqIjfaihZE
Cvruv8nkoJn0U/sMVpgFKP8OXgz4ZgYAcqwGQ/0xZXhcAZcs9ZxhyyD2LUZ1PDUh
WOe/YduT9GOsvLew92k3ZspVP/boBLc+wWq5l6sKFeV3w/k6bmpLPYQ5ehU/J90l
pfg4CRDg3HSYEf54/rXjpDCBaogo+Xj/MavtKDtZFJA7Q2CKr5YtkAopzFs6G/Hq
Tj/YRYUTxXiGtKTx7aKM6q5HgmcGRhRADo21OrbfYYxC2KPe+MBfgy850kdnE31L
AJEJQLb5xNLY7x2GnAsctE/crE41BMKHehWXyUf+Sz7sHvPPxFLX8l/7udxhqWlI
nnrgQPFYUfURmgQYsFwW/gKhB7Wz+CRgbX6hIpGqN8nUGSDrZNEcslS3PL8ITyl4
9vaKsl3e8wN/G/zeFgBxeXMsZd3FugwbkteSuEYdAKyjEESDwAGjjuO+Km4QPFlA
ukbCdGpZmwEX0izST7yLonwKE5zJPaies09zkWu6M6khPxB5acEa0WI4twq+SgYb
f+ILyikhCsefxI+HBvZIqmRqdjexxYwgn/LCRWn4XsXxSUuhIxC62++eSrHL07YU
z+lf3kbYFMZNWVycFzOhiOC5JW8jIVMY6mcI69c+5aV7nbnvBnq7ew9hsnqPSsCE
XvQT9Q6k57+h4/iqzaKqinwfgHPBunOjnBwLF2HfOxb+Bi2nm1fSWAaRIJTsxYR2
Ud1wL3shbRRePFkfQIKAyS+up68REbPWn6XpjzfodIWagiBmTBAfcFMI43APkRoW
5SXpQtu78cPybaVZcsLeREmdLiWNnNKi4LXR/EDekzZC8lZRr2EoIbJelERGiPPa
PWrLX9MAC/GwXMrzqDl56CEJeMj7XrVw3Lp6s8HsbGdIzCELB/h2YSggC8SljjnR
/1zXU6sgmFsLarAYLJyzUbaqFttDAw65HNOAW/SRw3FMvvoejwpJouv7ZPOpjbxT
oh+i/Jcz4dRiCtnCAj6urFqlfJ90Qr+qgRow6PN7pNhhs5z0DtWsJ2wd7T/7tS2+
3LDDTQZLirVFLsBQDtvHWdRqMAg6eRipZUlM1eT730RY/6Qf//MthJSPDslgKCQu
kbZ3o30NxHsgWnDuZ/na4/1qEfYa0/TxiXgtJZdhzOtvcfPsfEO5YCczchgcP/Rb
rBDnDqunEBYe01kc/DqCHApjbxgh267MW6L8Nmv9bG2yK7ux6OsyeGMI1gWPIKKO
tWxtX7sDPxhB6s9+43yTgmPtqTOKfm/wgd+gdMqwv1xQp9u892uM8nYMj1PUCC3m
GiRwOjGwOLiRBwHMofiGKN8epzvJj0uQW3OVFsZflhdu35EZay1vBA/MtvKSzsgJ
4k18Zn821ZuqZNF0nC6l8UW7359+b5WBoMaymrTtPcuQUWcal82mT7RA8c2WZDBR
cndA3cD7PqOTubtgu3HgOKCoPgQLLZ0JjyX+p6S9FndpoGe9t8+5LgfNqpQPWAFu
Wvsk6F7zfklYwVHTX2XKsVrDh0WpmGTV7glqP22m5w2jRG15AB4RpZuipApl36cF
zo9uG7OsWqCv1Q5gKbX4PvU8g1z3wZNHQxz1yOgiiC8d/augpscqyU/NnIKXtdzK
PsuHzNbavhGrn4XfkcN2hjXTMK3KJL4LX3jdqwi2ZhydIcNXcLnEt+UsFhLbbcT5
WC/NMv6IMVXCxdKaIC92jXs+uRC5X9DXZvFcGIs5uSh2CFn2K4YZmWwjqqrPedB3
IrUzMQkhJJwTdeWi6qCkntndF2OHoHQ+XNz6V36GWhnSPobqZvourzM7xAq9Jcna
4D/HP3by7bbnd52qV8KPdr/4gHlrDrF7MH0WTyin1H+Jhv7TVNwPZN7nehB6phQC
FMf9GfBxRFbgr5GddwU5uv31N9NGlNeXxdXLr+gH9wJiptWVdbDPzl/nVOTDmqdN
LmRRm/XrX0xsU8lfKlX3jylhuaBBnl7JlqBLCcdKZZf23Gcs4zmHP+TVIG7qYS/d
1K1uXGKOYfo3F1LfmOPZq6gN8Wlan2EqfEzt5oncVuKVZghDcBxE8QHlPSzd8XMU
fY9rUx+mTZmgrvGCK/oclYmc6USvkfHLEABLPv6bHAg8clIhEJ3e93fmrOfHG421
3A5H37ZVSg8w4eaNc5XiSOrjPk8z4KAW3XcQoyKkWNWGUHJME8bUsirFqU+yZ795
U31rOnfAek2yH693KIFuek6rjhx+pui2AeoVQPl3Rdxu/QtJf48wwsMaZy7ECQQ3
dM5+h8Oaqh81PcqStX0ZumgW/sJphYoncA9IUZkX+64TSfcwmLg5ewZAOvjpc3LK
UZh6OXNyaKQi1JfobJfhFpkCPJwodoRn/Q4MK1FomKW6Rt2JR89XfulJKPphNCC9
6XH+B8mi7VYstk3q5dZfl9RpioUQ5Aby4tm/y89orssvxCsN687/6YmC2jzlf+fa
P4pZijSKEm0qMgZ/aQyiKLY9mDPN6jnSYgUz3rTujMlxxrFP7WN9a8HreFw/yfTE
xN+qCXvhLgQSnqlJJFOdGbN0HlmnX7hnB/o0Rh+kFHSRSfqnyY5ADF7va1Q3layD
I74ZgwWvAeuTXmIdE1nSTgirhib1/oZxg34MK7NrnVIG5LiN5grtP6+k7urOC/id
rw6N6diV0h36+++9TCDWmCxuvJ54GX1GuG49tXrWTs2sh5U9XS67O2TcGijtD/Kd
7LZIN0vlR/0b615hqx19GebiT3R/b5QZGpvuMNB6D+oakdMgZMy9BGtdNMyPgPhL
vOAyqbl7hQunYMcJ0HLOQA4hlN5FP/l6YZ1ShAGXdP2I9UtmL+XEaLp6ju5ao2Uf
DbHbIsTQ7FNp2TwrbEVu11Vqkop+5pkG8tE8IHP05I4iCclt1XjMhHBO73WTDZQ+
Qq4xgsmUtWEf88eHY7A8czhhzoqgnsVhSrz3dWRhbyJnfFnDbLaoocYIKvH9owoA
muZkofwzAn+kxaWjfwouq0s9Iv7CkupFjN1vuU0RkicWYZ9gMt7bLadpJtDpzXOO
NaD3JSPXzqZKM2d8ftM5dXz4jjAswN5V+YP6HVkIn47C1FSt2bzBKNhfX2AWMNux
T1SKCVnFGuM04H6pn9Vw52ShkoxLhnBcDNz1yvtDUneoOCI1h9LXC50z2DAqN6lp
z0pcBqAi5lVU7kFkF8Da+QBqwjoqXCVm/NIzGbyHgJ0Sxbu1q4fYTjD0C293sdr7
kxDFfUQsc5nLZBTGI3JAlhyjhfo8vXzh5P0AuHJ3BDlCt8ktWE3E8yd5xhyfKfOT
UhEnf3t/USeftLiXyNxs3IIga+XnKD/Q4DmFWqMQ8TQNxW2fxcDzs2oBkV4HsJH8
1LeZwXkhVQ+dAgkzeWAJyTv1cmEssj3WvXR4lxWJltdf84Ztuug+pLk3ThyPNC7A
ax++sr0qjXlW5HHxUmFt9D3SH12Z5Dm6CuJ9PLl4h00hyoFq944o9SIfmm1kK/IA
PNYA03UMsfqhaCHWWgY9PH6yV46+fZ1skz4ypLKkmnNVdLomzHPT0syKg6odmCIk
l5nd+RxHIgGLA1RKT40SROUU0PfjQYF4M191sYI5k6yyHYHiIdEiMFlJ5EFO1d/g
NGDm8IUcTxgNa2w0G1BfiCPzo9TLxjyS6r1OVzZxpBs7Tu2/q3HoaY9lxe9N5W52
tcvSwbMuZUklcZP1gkPSCMjT3eNTeK8RBcHCqDAMQa2rkOOXMX30jsC9TKEN+oeL
zhuNypiE7AGfRC+Lhn8vUwzrU0I7Ic57YVtd5TMeoCWSNj2mTwl1ByD7EIxyO21j
nK+Bb5MaUqwzXONcKs1IFko/TCUHz+rKt3l5sDXW70I0dfIcjJriYyzv1Ni2pdpF
MsMx+FJydElLqt7MwKxWIEHtli4EC9cgjvVIbNcqvsoFzaqj/ns9FqaQGkKEb1IU
LwOkdf2lnO1I1esdyhJjgJSUS8lh95wmbEGAvTfhBm3MtrxEYtFyVUAohelBqlwV
vKrmEchfoGy+4n5POCjNm5TGD8yjRAp2KCEMhDCiw3ArWblz2DLRV94K05A9LfPR
JNbWFiPecPouR1EZEkLYPA9hLMO2yXoHTfq9ohD5tVnaobuu38y7B7U9pfntsI02
uUrnOdm6Wz93MnSeeiMoaBQMT2Fc2gfYyqQz8x1J39u/1MxUybhIbgD1ACLWMknj
6rrEZ6GkzjD+AxrH4VqVkL286aWrNcJRaQpE3A0EnkFBRt1ZyBAeHhIy/T3TtXaq
0YX5op1qqRIe33YiL7X0HwVdnV3Pg1iI6ow3j/Y2umXtppiROSZBYYPIJHMgBeKk
fo5vHo6gXq1NIkaQ4Nfof0H5iCOGmRIXkvI5AI6GgK1aOdn+SeKSEUPQDi5roFyT
VPf6WTHZfv+ZZWLSWSG9VADQpMAU7xya1zUiSsvtcIM+JXJHahJMr/mR/JaWr1Fa
4+zX64bF7yowPeDVwKW+M64x0Ul6n1iXUcqvB4zIVOrJ3j3IR2J7QuUQMira8dIE
xLCr1FcZqLRGt2NYCqnOl/70nhAcjY5ZpCO+9RiAHeW0KfaQ5TRjfxBp0DbQGBVw
qMhk8878fdWr8NUisvu1IJpkR/MgcxuYqFn8Leyep7mCW5GTNojR8nV6XZY/veTP
ITycowxCdnf5FHhbhNy1f34VclisCdxxSIwaHOUDye+baJ0lJ5MfbEU58SRDFZBJ
kqqHZlAIHCvPvOdvGUcHq7E+v7sMhlTygfHxrTutUjiu8zZGRxXM9S6CSF4Vz0Az
Zug9j+Iq0B7pkEm3A+GTbZzjUdyBYKUOkFMA6rR4aQoBemL8aQnCE9xJRfnrlhTB
ceXpTRjSl9IyWI5VF6lz7Gx4oP3aknvdPK1eKPoNy/9J1hjMlJBQ6LipjD6Dmrgs
y5DcyUL4ogQONt6JhCQUzF9/jGZfLXz0PCrP0myXt47FUfbJ6G+e/iM83wOPJBdZ
YpZvPT4Ri2yjByH6gwy/acI+L0ohDl/LdOHEOecC8sP6GPnajjNXuGWFWllPOADd
YXdRKBG2wmczdQZP7B7LtN2GYw4xzYgSv+MSYg62jjLYI5644ntA6Z07O7JIve3j
2IhZc+KD8EwQB7uBpYfi2Nd8TwecSTFG6HNOqiAhY1FgBKFF++7oMg4CrSE97GF0
W+rCECcudNR3Yg9YZYa7zXomAROf5iWWl0I2XArhJRuWnbjJNrKEX0FKOCD5c0ME
QkAVrYytEBfdX2i6DyZCLA1fEw67y9P9HxdfzjC0vQbdP7yN6kUEjr+6lOz2wSFu
S3vWZMd5WznMKs22ZSldiK3KsuSX4Vu+GxDOKpfTkLuZFH9onS1l7uW3j4lSfaYu
CqQBt+IyTIILuhW5FgFo5rgoD81KCEMy0e6MuQX7RNsO9ZpGUMNvN+Vekg+qC2Rb
PCjN0ia8jWWhWLnAHQJxVxBrQDXcUwo40pKvFT2hCYfm+DLMQEdPBMicxVMSoRjY
JAIZv+QSFJWcJ+6HZS6cHx28jNIvcKdr9YRUJALruJ6XiYOygZDbDNytruTy0B/d
TpeztbfJ3su44Aq+QVaSGhsVnu1GFl52YvW7WK1nnB+BjqCmWoC+sH3vgGJgOFii
qpNw5rbPgRQgndk6WmbmaF+8RrHIAXu7SHjMjUSSBvRHbk3WwU563gBbN5f0c/hy
bM13vC+TBgBVr3d1/C+d6bLcYzH0xZrKarxZmptVnZZNm8iP8McEFg1aB+pVeZ7r
1Sqx/VA+xcu1G/RpbauIQC8tn2JbVt+FxiJ1AoZX4hGdLdqlIEa7ALWmNcsXRWUi
Xs9rxISbhYciQtR0WwEP6ie9fXVYOdWsk1WMxBJo+SJSpzypqliKe5B0UUiJRF29
PL9tHGOAOwYlhTBlViVSU87J9yIUNcfYcttFsWO18XphjE3hVrPTUuvSHEka9ff6
g7vh+ZgvWsLffnGBm1MmAW/Oi77IiRSaB/xz9T3PC1zfoeZ+4znAuoSMFMlx/mFU
yhVpsnW8OwIWqIRipiR01lsj+R+GIfiPh42vtE7w7nE1IiLqHdIfgOEPktQbMSxU
BWD9ue9wEwceSRCzNiLGeof4mC2zW+ofhd54PBDo0eXYswHca5NO1lFTGWAnYhC5
+09DJL98yjt/NhXZddbD/NVcchym4em3ioQ3K9G/O+xM51/L6ViFBMWItxxqxqJo
q+skTJr4ja6XA1QCwNtfCrpUpE4SfqTwII/aaXDTGbYpggYzWKpuIo9dzAc3TGG5
ZdbixhOETR4GskG03PdYUuSTVvjgbbSuCgpq0WfWkL8tnLqZXSqIAUqKaoHFZf1I
HPlYLEqs9cdUTXDUsHCs7jYKd/0aMM72F41PKLq03uIK3J6Ge8BF1CixJE2T3R56
z0tTix7+lCSXxxscHoNxhkggAMBaAdzj/IpEJuyW7EN6SqL5JHaEmmlimlf9Om5o
JLERgIbGBQcTfgtbdjEa1HzNi3qEaaPSaNlEio1KU4tzwtj4Q9NmOWB7h0um4cgv
ucMJCimq33oC2vysM0jfb4wf/uNmd3ORAdBM5EOE+9s0y/HBbMhN/TsmEWd2spk4
vXNCkNL8JbbzLkHO5H050JkVUUC8cJhrVytcr8pfL0CVPGnVvueayFZzk4YYuxDi
UoNkgpkqhhyxcQQwA+AjdmHQhk59b9hzOqRmTbZtaK18YSItbJE1M5ts71CAPVuo
nEwbAGDfXKSfdA+N4Z8yO2E7JY0dTsHUIxLy/m0Iu50zNv8uWv8ym8YJwjYeJll1
GJVHhikwgjT6ms5Fivgr27aegBjyHNFqnLcTWi3Jvo3OTZshcUxx1c6XYF1NTIHA
kCHP8l2hzkMXTJOunjSvNrINYN3Yqe2CWgmzHBHVcYlQpzhsPgTDeGAC9rMa1qhn
RkcsZlDb9RtyIht7jA3IbNlFms5Shij96c/uk2EtmNi8W42LoGpWGnIVbSW+DLhm
Y13RcDEK9djQxgZF3aA7x8jE7TyaDWROByTdbKNGx90mWZiI8ib4KF1WpnPUuhis
KHg/HcE7CLVzct7GFJD7QCWiVrEHrhKdjoTCCgIwQ4aCghZNVWx14FyHw4cdZ6dm
DcXPegxEgeAy/2Lb3UKyr81HrCtsnaAFjPOVWI0TEiVvxQSULR1FoAN03dkY1Qzc
BO16VnRA5JcRmLdpRBt1gg3JIT+91/dsv+W7g6f29tVAcC+ejvsXcpX0wvNczvlN
YEKrhfNUiQIi3WR3R2g2TK7uhUYXxy31/L8+CSx675hIn0k+JKcKbJJqQ6NZ6dqH
3nRvj7NOtfScz7uR7OJRM5k5CpIw0KMjCVKzImLexI7YDWAxDto0750ii3EVczzc
9MV1wLWzksjNQ7v/U0gqAcQ3vwL7Tf2yy7aLV5H1VPcJCwof41DKPk3tfZZUdPwZ
5qPVpEpC3k7oNdp/t1nvG37KlmPkP1HFLHi9B4/l+C9JpqqET0xoul+B9Bb1EkFz
6JZ/r0PA5vEyvqWXwkxT8mz+Yho/9w4t0tHGfr9YnmmmSQquH9wNieKIXHwqP90d
nzzaHFSHTtozo4nFR7yhs5p21VtjfAs3o0+ox8vRbeNUKZuLjtq8ZjOReeBGIMU3
4a0Z9deltcVplhlT/WWtQ9d5+DjimIwyQm3eOmy9Dk4qhu/zlWiDqVH3tbdE64oP
n70E8TbxDID7aO6Jma7tyPoRD9WeDwctWCorTyUAShNBryfhGFaHGhuNVEPiOaQG
wWQB5aIgzw8DrE5O9eGvDeMHol30DBHv27Ji4RgnU81XPHTGUkPZtPdO36JoAw/i
AT7xoB/hVEKe1tTxj91aPYcapY5AY15jRbcoEE9eme0fJ/1Wk27P3wYrRiid7vaD
qNaQLUJqI2CnRfz9TqfmlDZBkR6ZW/Z40flIexpuJpNi0buTHGXDv8XqXbxBYpxC
4NhtEQ8O2LyIpSWR6bIuQrtkmkyrrScA+JyLhccwRbgOT05OdDgNeh/mtbzv28Id
dTidxfrcbs2V9tM9BlT4N467YLcavNe0QI1teSG/E2zWp29OlTgJhXBYVxFo9P2r
caIGyS+IyMcsSarJdWDuIIQycYCBPlg6fQaLPe2c/Ipkqkpv8SfsLeG9qfPwKWT2
i63jzkHUEoXnTjZmagqJMoEMV3hRAFYAcnY8ZYUkLDtrycmoPC4QBn91Z3fhQBDj
JxBYR9rVQFgaIIvLkQ3ngaT/vJzhVJ0z0jNXMp5VDSEbP3DU76E3z6HB4EuHaxMP
Ey6kywWHrFliQTIGG6Ir5eGpeKdkK5T/AHIspA/mCwItYSL61Jv+ZQCUynPUwps1
6j1LQ42/Pk0xiyB1etpudX1tyN2Bvfh++GywPOCxGHru4aS/HEOoElkc5ySVWg5l
bfInOXgL36ZKJpjihpuFzTatDQJLJdFltPgFpWQmKV6YlxlvY9Jx3cSBXcKWYYp1
Gwa3S/IZxMX8UPc2jtnGE5rLTY2D/Q+SvBaelY2+YBSZ0nZ590addXIf2MKysL/5
x6Q0O9HPXa4qUVDFll2MIIULoFiTiK7XCQobbEswMJPecmCukrBhsa/JRpZpoFiy
bR9tM2WCc0doEUFziJOG0rPeSY+1f2+KZeckhiY2eorKlSdP39zioONC9yE5PGc6
8VyfCnSahyjBNHwigiNEUHfoflMgf25/34XXz2pUJbgIp23E3LBFV73x4jsEZJp8
XaWmnOY0giZBW+IKXgL4+Qk3awiRQ9y0JIVJ4Mt2OQLrA9pKIJPsVj3NSMYZh0TZ
U2JinA3Z0NQy8JgqKEHzUpawV4ISy4fe7IpjCCtTdAq+qKHHUbUYTTnBRS+SRZE6
sDC3QN/fKeXOnnVl6Q8y4qzpis6zuM/i+BdgVlpSfnZTnAgpbezI3UvMxyK4yECC
K8UBvLzj549tvYE4H/iXK7s8TI5ihOwa3BnppPumzVuYac3xApVzz1GdI2zPY1zr
5EbB5ks0s+eDcPnBCXqJ0qPfySwSgeHdZa+XL0B1KfdghDzFrTAbKS51KVqoWSyT
2SWiTaX6hcopxfNyenz3fzaM8C/cFYiEOAjgwyWP6knc7MZGcyZrRGPMqhWbDNtO
cOFuGchDvBZMVZ78aLSodeOl+dAROby8ygBTsPpJltKgRZkrtLgGSVjAiO7SJOQL
EYOGrv1HHyvU5MMDvNvmvSKccIRbgRh5gQvzN31lmPjx5qT2qkQNhKXLVEnRwH3e
1CbbH2CRnLLmzN8M5r8OBwSwo5wxrp6fwby0MSaPCFdqq9pr2F3U4O+IeprCXWOI
pITm9xN4Z5vEN5Amb3RSbkOhEUVx4g6s7Q2642rkj+uGTbx6qMAaPZJoa+Fkcvsa
51sfPJA7Nx5MNYxeEgjbhrnYFc5tbyoWk3lc5pKdwZH/VIJ7cTQBmVdWbdSulMS0
Vd+j0nsdOwoeKTKyX+2a7SApZEwbnnAqdq+X8KdBDPZS23I82QXi2I2rwQa/UUD+
31Wvlg32hZ8da3cvTM62hT42uQ9v/DClaAznMY0X4MxPa+HrF7LuPwCSMotnnvEk
KLdTv3BVPRfIbfU23R0Solxd7PGGT/mYPnWuST4foeyS4HvSFp8gsAeMvnqtnfuj
8gJhXKzNAHnf9qH6gKT2U100tq/7logEvozmd4AOJVzqLVg8BTaqNK8bnguhjHmY
xeI2cpoVH8Fva2nvlVmOF8HUzNFSfbpWBf5MfInSL/bqqj4rkcXsoA2aeUn9xOcs
joIKoG/Hplkk51RUsBgatROFQel3UUjYx0S+dU44uqVzp3pcCBYVWRS+FC/X1vF+
YpSuc94RkHAaZgW3X/v0DwgInojPaT3Zb52Hlto9VQ4vkg6ZkMiBd47X75MGdDEd
Ph0U4W+uXurwmSfULabIW008xQkrUlm4RMf6ycCDlnmN/u75jMNOZe4CBu8EdU+d
ZGEahGlZ/TIWBm0J0r5AU4YIccsILdVM+eM0/TkelFsis6ZUgwSm8a5vYfHFuUOi
W5Gq6XUzMX36U++30wY7hR6XgnNi00a/k+jv0kLG4aXQVoUIQJohLyrdadwccWjm
o6+htByrFdHgeSKOFJ5JPEJBapgxxP+xqgccyvwLZywh8NAfT2FLWYdpbEr5GPbr
v9PA3CZSHV60OYbPOMB/HOB29m4vW63/4QfUm9aVo/wlNRDKp5LMYPEeIrMmC2h/
ceJrM+59+UyoTyMj0ngUj8tdYVZIjzw8iOWKm6hAIEERpaAyQa47ZiJGXClN5lM0
y/1Vz0bNS15dGE+3o2oQ4GwDe3qSt3fHBxNkAC8khj+xQaQnSHVZPPAb0VSTnFuF
Ama7zkhmS4CShPpDPcqnn1oMW4xoClMBacLXJtrdJejlPpPYuQdTyZ+GYRhWgSpP
eHeX5JkCHmuDDL+Wk3TpjZxRAIfqvXYz5WIBP9UswieVLSUGWikqe2QdnZJPqTuj
+2YZ+HTl+NRMuxO8urv5lLLvAuvDx6fSZ0xM7/zD6ZZyz9fBhtUKAXcs5vvnNpMq
CP/yHwO46f77h0wzXfz9tDP4ShezhuKN5wPNzTxEgIAh9SKaACxV60yAd2fFwzip
4U8uqINxk43Mb8umKLhLo/MdfNhYWWcFuUWBR6bDlIMW+4Ujm8yQR2VHc/LkpbRE
DNj+6H4a69afxxVKIDrvM8hKv3Hh7lrg8xqBGqwcqqNKuyJPVDTGft98E7vCvRCF
/M6O2HmiA9ZiN13vY/g3ze8/XYpKD81VLtNhuVUfssQwxnBgkPF9ZF93qhAW7s9q
Y2F98jAthFD2V3S2DmQhucLjFs6S+m8mIwvDvkSlbA5DFgWZBxzeYMKUb0NkAGJ4
dFg1QzYu3V/DReDjuuUkwwQvmZU7nznwH1Zez8U6PqykA/rCyvnHtfhUwi+kk9yP
SiUsJu+pNYz2xdbZHa9BJgvtt7aTinaFyZy68ftA1qoDYfbBJtK1ZlMuhW9bRoFs
0e9YjaOnfIDwbqtF4pPSvBh7T89JWlfjnpl+Q+yZpifXT1Y5Jr+6TJb3FdWJRGyC
DWe2PyKlw1cc1h2ZclMsEu9sTEGBJqilpZ0YWAF9RDw+c/6YTCtXvYzms/yWHL/F
/vlDJ5kUTPPI6/q1DVK0p+UGEs7NIIj1fkHhsujw6YCrheGz4AbEgomqWN/hEWxY
AhRcdv+s2e4PgI/Fe4QGOBZIj1sK9ju2lAi0GmLV1VlLBuYtQJSLjgVuix5/t5wV
piQyY7xKNuq4CgbW9r5LAQeTWWD3nfZyyIz57MkEF7YENYMs3LhBlVqBEDj7Tu2+
cu1hMz3B1EM09PDhKLb1JcmqDSJ/xnpRliAR8Q4k1uZ/opbp2sQR3P4uJhXTOclV
tsoUudoPxR8WWb2hb7bqp2AMSKVuI6g7OdoE33dioLl6zDj+BmgbWwyy18WK1V/L
j6FLAr8n7yYR4qYMNOanUNyWqEd96opVWtAUU7r16YLj9EpnfX+CSOwrGhxffZSs
kr2MYFaASoB3I6beTuy2vnxxP9xThc274vD0fJG+RhlaEurEr/S6ecZY09qmCTub
695ZM3tiqaSZ1weB19a/rgaUebOp2zukkf1UnDs3X8ZPHxqVXDsxcTxYE1KOqObv
GszJzFNIrjsXOYBtehHWnlWPueQKFS/50suRNbqlhyjZeXbV4F4DsLNZ8UDEZwBk
zBj1x3dcNF8YeDLfcqaJSP9+sR1EH5/n4u5tyfXRR7KmH3XGxpmI02RdH0cY8ln1
1bpWN1XfXOFPq6q0Ig3qKpO81jeQ+/bymcPcAS+iUEe65QIBz+h1o98g3yGN+hIT
bc1JM0hcPZlzh9MlHl04byn/C2x8OKXazXdPKo0RUD26f/nvNLaj/Sl7IDZNNeLa
jKrEXf4xMxPWCJymoGIa87iEZPKiXXTOEZqXqnxsdEkxMxvIfuae06OUghFEn5bg
qCPvORPlx4HMIa93uGTie0raECM1Jp/6Y0RTFahcIdQ5paZxNzuaPGNt6gG0BAYD
d2QKUGWIJUKP74u/MNq+uFkwArsPQgVIUlGrGA6OBIpwLNA/0kjeO1OGeAlmKsDN
Oje1AlCC2k3s5i3T4HSUogQ8pDH2M+n8RLcsGYgijd+tnhIyLuBfpWiodq49ujs8
0cEJBNQQ2tNSwEFYE1TaDzW/RrRHjkMQRm3CzpWWJDA4iGaK//6w+dPwrwa4qUjc
f1UGsEFnUFh8tUjnNXGYF1jSWI7H48fxJV3GduSqjrqMIJYITAL90D6DIHYZga5J
Q0DDV9xrxkrY0JVOrU7ciu2tz/6pDIz916esHN9OSUUGZMq+EVSQkis3Oo4tfQua
9E74ZYQwy9DaRx/ghoaCIffkwfwgJf5XJOGecWUwQEJEUfByw2N3ENU77wlg0zmI
GEw/p8I+B7ZguzMufOB1fwptuXka7eusK0GKrHHVf+JFDku6GmCwPBAUVWORXV3H
5Ql9RU+mSqP3Uv3DE+jY03cof+V6YgN2aktnN0zuy9i+lt7UC7XasQ2ZLRdSUxg4
oU2TpqqaH829Ci3pyYSPK84aPbJrO19nFibBfm2IT1tL6fhrT/up4r2qGrTG3Hf+
ZZsp4HXgtnE5II2zp3OvPJLN4GKyhfu/54BEKw/s5hkm4rA3bEHibygdlcj0LCAP
EGLRQRQQMCRTfOGi7sN573VWLHoCn82v1HyWeC1yHoqdN+a+ul1KBIevYCOxdGhK
WYAPzXkm+m+6kHAu7ieMxsU9TizhsR+bo3MYoiAiBTn9xL7KwdfrK/lSq1IqxVql
S41EJyypBnjXsVSZ6QVB0kI/AfwbJZhCkpS0RrheR9eigjxldaIg3ZCs8iDjXqhm
khcqRo+Jxc/h6WAq3B4mTgoD+tt0H943Ch3rkaOUtCBU4/D+at52TaS9zgji958h
s7EHID6Nxe2jJHTEW7DxEUzDsPvvq22iIpxc11QQpZPI1vS9TzxMX8HutpZYOfph
iRiXjDk9yowg0LM9kY6/jJAAVK+6r6P3QQIA+WvvnMP2bapSb5Ca1ZvpMEOhCIFq
PRBuuuhNbWaoLEgZG1oQaloSIu6wt0hsyclwqiZJCuT8IaL86kYNLMDtsUPDR0Al
yWFx3EjEfZ/6vf29PTCQMZbCcbWAYgocAlpOqZ/751Q5jAn+CjQg3eIVgy5b/auB
GTlsVQT5JuvLgoprjCTbDzRCl6a9jRLoRJeEuOFs2ljXhTS6NA+mjplWfTLsy8H7
Li96mCZXHwFVkFv7e6ukOA03yZO2AujmCG9BjLBZMZAotpGKZydDoB/J3M/mI9hP
2GjI1FTrTJWgk+l/grQzzYb/K5GFFUIah/Hl3qku5L5EoZNlW5mP+LNe9QDZ2VWE
YcG2UGzXSbs33aWhddGpaYHyQH4YsngstCF2O1mEAH+b8QZ0oMs5YDHGqxCN4uY+
c2BDAbaC3cplUYLTw2lrf/vCZ7b31sw47MZa681MgUwiit/MNXGmK8Ezm6/cVeNT
R0vUbzCW+yxfxlVQzFH6Xg36VniRrZBINkH2y53AoEaFSHjCN9rMTbuuuXGVKQrU
5KGV4za5xq4qIMg0mrnlgD3khoJfTnd3TSvUV/hCo522aab/aw1AfIblypTdOJed
ghPuwJNJ0FAQXIOvDU9Z5o/foinFj8AWVO1efINtiMAk23hi3I85w3hIViJ6c3v8
fF4Yr4+Q1Oj+QfDyDnpgGRvxVzqqgYRFcL+/DLiHFYzjgImQOSq9/cwQ1JyAQ14w
X836w9ayTwGyJZZN/kesNJM4Tm8HgPGt+KMrzpuwiml1eTDDCcz0qSR58C7nqxjl
wRFudDURoiHjXJoCEUAlaDb/2p0mp8S38K5FmOjOswxEIvdrPXsWS/SQd1jYAcrU
E+YHvwLtZtS6roQLs4M+3062DvaChTXtnPOZ3ePnAo+6Y6pJ8dQvrM/HDTb4ysmX
O6t2rBP/0ceMvynHGg6y0uQUJrOkUnepBwcgwy0HeAdimyjoh0cLaD8+JQivG24d
m1y/8HDuO42i3XxTzpSdrVto+48G+K8JRoy02IHS50P0ThVh5B9iYtFsRJ0SHxZh
N6GQfhTi5OpmKbhSZucQR+Z3vKYEcnI7ZRdfpLKT0pflj/EsSH/QU69Qx8AbkmPR
8PAIgbw53HDKW294C3g6xve89Fmjo+qNe6Eev9JE2vmbranqsJd7n+NvO525nD67
nFfuzBC1NaWKrR1eAQnMey4Q411MZf6VcZ48MOlG8juATSdICcCEKiVCFuo7OjY1
IIMzbRhD9N11Z+vErBr5Su2VInZoDH/d7xOusI6FuKHNcdmzgObcMe51WKn1QtHL
uNb70/ALL/w1gR2X12WRVMDiFJ6c1TUp6i6XTJ10musBO/qAPP/1vBTE4vzP87+Q
3wFXYhPG9VisvZ1WOMyrJp7Mvcrayv0hWLCtTNkAQPGRUpAOjOCrFrvuU4HMg5fb
5EKM43T/PHNJx08P2wPJPMos64xVKD7r9+sofdeKifaGycx7NBv71X8wh+S2gQ42
Jg59W/fBmzmXqmjUVoQXNdYcCS2yt9XouVCLYeTfrBxqkOnAI38B23qb7wvmuggM
01SeWpEQhvz7iyL+wCIy1uIxeI/f35Y5uQR0tmurSGBCVfeYqi2m2JP2aqhkwdTt
rrgkBHsY0z10fEx8wCdBaYbRASBhQ33W5m5NAaA7Tk53BuJbFeR+MmR04UVKyIsS
6EH6+5e3Wtyk7IE2AMeyGnPCraap6be3dumvSLSx4wRibkQys7MMFdTmc6kngC8M
OBDwveK2TbVGlKZWetyLzhoct5lWJtc1yqpFEV+Hm2AZePmCCKLhu69R6PKcYwrk
3+j1CtBE+7KLnhNe+Ym2xYPrZcALg9l3oUQ+1uHNz17lM6JSfwzNVs79e1mtZSlY
ZFud8wV1hrUYsK/jSnHi/vAmkP1Ss+uyuqkIsCtzVBnaByBxBavP55n0Oo/9jZrw
yQFFi4TKR992eZiSZZ6ute26v2LkO552wADA5G2U3gf3zYSCw0dq6Em56Aon+0cy
5HkKFCcc0f3mTLHE6HVO8A3f50tCuO0KNEkRKs+OZ1+K3UlxWh75VX9g76J76BGp
zwmprVrAyORhlwytnqgGNkWQiu4ozqtj81njilFXHHaPvmiSgBnZDU8vPLgbUp5x
6yFut51Sp4J/iWoEZ1JomzXV/YY9oYpYFJSh+9WkURGy7ufq7EMN++LMqVJClx2r
yYMSARdzoWV8z/zduI2xcnKwbklEVsgWuTSYAMPaDN25yUhePPMzXykZ/e//PIYO
j4xdtqt6++2L6zPAHHDMQmDoVa6WallMw4p9hnV+W0E58spV9V1dUXX/3FknEhV0
IoxQSmpp3Vmf+rDcevSXzg9YUh71CwFndTrmP2Gg7odVpI6SwFwPwE7j8hM0bFAq
QGiRY1H9EfFi0Kvhx4g4iITBX4C6WHOd3BRVTNCLC13ykbGPCMzi7qd2irA1v4hF
Ji1x8ahhj5FcscPFXrTTvFkQHFtEKstJhLerMCokG1T75Jlc50Pok9+HeoHDJ0xE
j5mZ3uj3V1SxvWcL/QUYD6hKoQmXnhwDodZU6NcDv8KgZtNPI8J+5dlOhMxUb1JF
nvwrHr7eKnlX3xF0swg3thNlHQEH0o92DFSOvPW7z//QypSQ+o2zNWG5fc07F9ls
8OoaZMPIprb1kdF6wgTYcVjdiaOWSbL3KqScCxiR5A8cxC5wtl3b+MWkZThS74Mn
QlliiS97AQPMmzA3Bb8tfxHxjrLW8kZpZZjPnO2PP4D0oD/YIKLrT8j84mReqpCG
ISk6OnHBCqsVm/XU1bKSjioOcsXg1fMiGYkbf5v+M4Noxb4CMoe09Q6a/HF+mQjy
YiVgCrRp8fRAeKkrTJVA6fNFBAj4iCpc6P38bYUy8OMcDqur67JsWFCEU+2TcyjJ
HnjmUd6Oxh9sxlTScd3d+XgSTKP/ZYC0q8grEZWwRwLnp/Ebmdz//bJzgCMlydy1
zmBqBIypxUslyaKjyyyHxS9HABb/bCWfRNdzPMg9l0E6I8vhp2HqN8w51OR8mRr6
vWcFqtWHcsx71Sc/I0i+ZvHLDK5FWn+nMP8YL3AfKAKhSt9yN2UTPfJpxiTQCYpo
ZpJx0/htUF8hZIs3eqHFwb2Ye/vCKTqqMSa51lh9w13XMoMLTColKktLzqfNW+TN
puK8w8Soxnk0J0qtDDBSYcYubFJ5NX3qgq8kS+/7kyP8HPVogzg+k5yxBgUYLrHf
IK/Pgy9Kg8rmelYHpEMtqxjdfAg2HZaywprTeOh8/6Xx5r3Q0kH/SH94Q9O/w58N
tb2FwYqkEYXy/XA6w4p3TyFUHepPBObmQCHzJF4eOgz34C9ZzUwkKBs+k//5sVJv
5uCrt38vVlaR/2YWTeQXJ+cDuhIyQXRjqpfBVW1Ri/prvUthzv5fTE9V8qIzmBRB
tjNRzcyVjXRNmChwVQHTKAS1YE//p1I8zENICP+q74liKsuvL5pxrUYnKkJ5ai0a
Ltw77XyumJMyLigcE053FV6UyeXfYQjCo1ih1PQPJiF5j6lq31ScXaZpN5FEmYCt
wN0r18rRYdZr01rcYeFqCDgr8bgIAHd2gEvza21BIDrDaoa8ZVI/Sj1TsDG36Oku
wcc7SxPniVq9rcrQN6dMDQwyJdwC1kLhS8Wp91Bs3mTk9omluEB6ujvRDXxJ+pWI
Tzv3UHpCtbSA9nP0d13SWacqGdMImqy4L2w3g5x4Spn2PEaWloFJFk59c0WNvUhr
1i9RCr3j7FkaxaGn6gPuUpjT5GZeq64BA2iWO9yHEfaS6NZEP8RIF5MKI/xlNjF0
rneV4mXKV8u+ulU/s2TpLpY7D95xasJ5sv78+HGA6H5s1WK9f7NOWJsWT1u0eWhs
T8QoNajwBGafLdjU/m0V7cwRS9o6yrQydrL/xJj0HuvHCfD+xxiniFvavxcl0LWG
mOYsF1yQ/7ioFHdpkTa+2YVdcs9qiiNAMWlA6x8Hn7ypUxpu+cliXCK5e/ChYm+6
nI4BtSl1pr/W0hl+0u+YAUUHSfqvCPoXKOMNl14yJmqKMvYT1TrcHPLEBzbU2e7z
1QFs8sQgpBkO8KsWM0ekM8ww/PU8eJVrqqfZl5zZuSWviatcczKrCf4k/41RiACH
vXYTsEretXVX1FU6dU8jqd+08ehrgsNLOh0a+KALivLhmbfnvdAqmwNAC0B/NG6Q
kZWIk/wgVa8h0CuAd6boVqXNbw2Xxd+pTsc8EqbOKU0gtAsupj0Hf2JkglKYHtgt
JkXp75jp6vpQ37r8dtPnmdYtL5zbYgNYHFO6Qpc+oJtUKB/7UzzRYJ7mn4otx8xm
waWoDFG8TvDAQ9sCn92XdjRql1sWIoFm2UNBwU40RuzSulO1YUQk3uWB7vDulEEj
z1fTbaGiCijarxiwyNfNWcwYLHD+nUrVSd72Fd/K6/ZiSEzq9KexkUFGX68vtUrV
LeX3+je8KLRpt+RbrvmIsyRef8C24canWI2bb2vHsOZAW0Uv8zt5w41exLqLv58F
vPt2GfJHr6IVUUtFyKNVbTAYZsgT5jrR2/Q1uaR0Qht2H3IwG2/quSWJNuJ9V0ra
zlzDsy5gnPBi3+cX3v2RVR4pT1LI9lkWVV3GQWXN3XjlQNz+Ft0v7krXTgxuk/XD
uklcI/0Fn9zEE/dpSTRVH3ynPw/27PlWKrkE+w2uAmjUwolZYht22w7KCPizFO4l
twjoCd0IFTigoVs8sZppV8Tbz6fihRuR5hiH8pLRS3KWq32zBQmDf6S+r9h//Swh
5BfoZZBdRVQ6pwD9ElGl7Gh3eFGQTSD9SkuTuF3/SFiUyKqlGSCdJtzG/ju+81Bu
RM0WmqDhq41g34MH1IG6dgsatl/8H5pDOqVWD5/RCrV63zIUoxjqTYKrwLUfO78S
OuxuE0oBAk39YWUO9AILeI2ar7wJhHiM2yCF34NMQ0WMk4k/fdvvwYVbQxqW6wyM
N6iLdBdHouHmlSXg5k1IqUiS4oyEeJU01dNkZEtWbs68vHw8FvBi5Ntl89lujVtQ
7+k0VLr270Lf+GDA4o5VWB6Vpv3Drh7vknpVhHIAozVke3oqUWUKmYKx5Kr3zpFS
TTpHoeYSIOgagcgDqJu00QAYjjOpJa7tXce6Iu5wXYhHJPjAhV67wPPdmEcjwMU5
8pjgnTLodByRRcBdQqI1aoQPWNxV8IJEDA6zIAxV8tPGJB5af0lh9hCeUuN6pQo4
CGdMcdfKdqO8QecEBisUktz+cbsjTFuZ0h+dbHOKZOaB7x2WcJrL1AgDpWiQa/eo
mVYkd7Y/jsMRsoNFNxE95xNUo5msbzEqxAP/g7920yJAYgZxNBUkyN+tsHbyXT29
TVqCFEH4xVUCPQm+qHcuTQ9RYIsCTso3I0+aj0Gz+da7RtFwO4RA4sw+SPigGiJY
BA1NNohWC1uWMyfUOWtV7MmCE/KCkMkuoF5mcFbJIqiIZYXFYwDMiH3OifLeCH9P
hITy0xub9k4kA2EYhyZSJrVY1nZZ2JNEe/u07XfeyMae8ARhbBtQgSD2nr3K1qFb
SSH125YnBoxNJBRupZOBySfTWyCyBZwMXDIpjWQi96A6uA48iG0l6wfpE7WNlRkr
vbS237tgDgI5xSiCfp0HuAEHbr0Gq0xHh1exvTUvt46QsDJAMp7YKx14jIzPlgAj
K7l9myDL5WQcuMsFIJ0UDAwAB+ePFwAq9xtgDYv3z/L7qhsCeYAwtZK74MN9iPlj
B6ay25Ey0ETgx4j38QDxI4nQoUqPbGJzoWOXTWiugVVoiTmxCn2+oOmRi7FylsX6
7IBqwAwSGxzflbdCBwqWV1E92Gl37xYLwmMQcBZjEPG501KrEPgXIJBBfhX4c4i0
f1h6QSYxaPf5nc8z14zGHJs5tU7F7qwesrfQeXMhJCBU3XAmPUnDKImcap+wS/2o
Gd1XyaFFMIkNvCNR83I3A0KEvekdP/IrkI/xOcysHyG3CBO5jmZEcKn4PZ2POLCa
624OYCfJq3Ionj1ZFPdzLg1jAGoDCGOKH1FXUGnvO0BaCwVVR3xzaAv5u2qc+7G2
lcFdZSEz93KdjxIcnl1KyXIFbXmsZc8A0L8UqZGVY6blFnpOsQHrJNRmUF1NiQcl
QZ2dlNVb2TgfzZyLTF6XpGbZV5bhqD5fcYMoKW4cH0LkDeYMkqK+T9eHPX12efTv
9OY3wfWW0ZmlhoEt9NcaDn6wcCIkJvkLjDvq0KdsI+uAqtvZL417LzW8aXU8rK0j
GsEk3/mqtyW7zvSoRHZrHSG1a1QHRvso1hPQKAV5XYqfxAOdkwSeyO7lXMV2FZBv
x18nT/8HqSHbSZFU3JjpcA430ZsDJWpp/g9zZXjom0Z/7ANJ+Em6YFeAzKfFGdWK
tB4HOFFrANkXQprbjb4Ms+IW6u7cGqDL/+eMJiHc0eUMHsfcINk5EGo3um3ZhIKH
mO97nlXvZugilV7D5i6WYm5KlRARBvUAo/WMrRP8yOWY36MgLIcA8zRLhParNQwH
le3SJ3m4o6nSQvrrn9nktTmyZBvxTO2ps5Q3YGrZ0ywfU6taPiu0Rl/H86QPUAcD
slOamw+I80wreUJZf/QLpmGmNxw/k89H5T5/OV4fc1pJTJl8ygEQDmAR1qXPWyL4
V9PZjgNsNvFMIEMXKL1FhlP/E/SdqhbhnsFI5Dlsel0IMzEPQ6sDv7La/2m+E5Zr
tIB/bUrf4U31YPbMAlXRfNruBT+aTDm59k65NVVve+hJVcuQ7Tt4lUBSKd4PjT2I
T1k+douwmYpNyTx0qPEI5s2ZOKR5To2cEw818eYInKWLADa1Xmkm+qFUK5pOqRGg
ASNx9KIKD5Z9ekhQt1el1uc8Vf2xOBumW+rO05fMzXIwWGW5vHAENjUZEPl8oYSB
GRtX57V//9m235wujxpQm2zL6Z7GMk45DipMk8EOpAoSi/FgvFsDF1tfqZRPB/yE
nsl488VrhkNZ8vXpZwAFGwut3Ip57QVQ3mXttq5U9v3XS11mFFQOhVg6LkulluEt
ggzyUM7A2cJ7ix7XT06mkFwI2VHxc5l3JT58jhjGdjkhi9Wt3SPXUpVbJc4W2LaU
ZqGeo5TAspaxrLVKrgvhqtowh3WVCsYCSs7XIBVsXcIgJDVe2h8em8mlS1OlkNdv
uBz7G1o6X3YJ7EdlFmTfWEtqh+4lThLtfBdS25eRIPniuzz28vfri+YxVboGzpZu
7hWWnan2UlLMbvx0WAfwWdMot0HIG0HIBbDaJVjt5o48LLGtRVWQIGSnSNdC0P9I
xIlzv0M9n1onorQNpCjXw8vQb5p6NqUtwal2aQ1jvZwtWYtvEc8mlhO/7V/alDwR
EunMYdlPLYpKwGOHQp+zCTwEhKnPmu7sttCACosAUIVixSMPmZ42uO7k0xiLoAsA
lMTEGyNHaTqgHMNXO7ZK44ELJQ5L/LKjm7Er7eX/rzipjvwHXYRAOg29oZcyqImX
CbfxHRD3pZby6/RzTo5lkSQFuYWu9Ca3leyzdmBtUYXdY0ensw9YRiK2hd2xp3Ei
Odi+SZ5hdWa/H9IG0iHGdtQvBoyUIcto8JLL4xtgYw5fyx0uo3bYTFXEu4tgX+mC
EXXzTVQJs/r130uk1c+KqvuPI7MSuTnzbci6C9Gz4BWa7muEwKpbEA76hVDYBD/i
GxFzOpQDx1MiUWMm39Edjr6Ugvl1rdhzyW3Y6+nSMGE1L2dJ2OtkA6WKW2XQwjgT
waQxFLTrvlTyovAE3HtTt/tkgeCcMqZTXiD9+0dDgVSNN2oK2jZY+RMym50BHzNz
2PGUGy6vCT1cvq6hEpTL8evl7MKjN80CAxZ5w74yPqlsT+fCBsF+Z4w7WPTQ0h4P
DbpLrYOlbvnWIBTk1gcSGS1ec8pDhC2yv8SdiTj/eD7WRK6vTK0g1j03SjeCn34b
xds2ZC+TUc8oeARQrTk7gVLLJPNkNRanRYxZYDj5yE4ZV+6fHvUrj9wRAu1UBjbK
cATtuU32w1mNP6ObBKTbgrpcoR2qO3iWVi7MPJgLA2gzAzJ6cDKyDPgcLgQodDA3
I8X66aCJ+Z4hFV+JV5V4mdpnXxqPX3P1BIZXJAPme5qtq2qOwPu8xMwulTWU2pxH
fXuORsh0Mno3O5Ix9+0F8CD1OnigXh1dv/CxPfvb5hUFN107EU4Pbof8/fC5XoZD
GSbJBSwYcv5UrgxjbFE7rtzV1SL2Y46gjEGtyZz9eoUoekm1bSW13kjEmBWJGKU4
HQfFCjKql/q0ch3R+r/TgoWWabvVl+vftSDgZKFMziwOrEDybRQLsQSYK2+6c2j5
55PrrP4bB6ayvRMPhuuFAzsYPgND/VbgULrUf/HKG1uv5T76JBjjKaWwuAKcoVHR
00Gr9moSxerw3Zapm5BG72mqQytjLdZJpXnkCC0oHCugs+XPTcFq4sDQphcDR9Vj
3mXjSbZPbw6ldT9g4zL0bfCslKgFupezvy8uITg8r4jyXT7A5Sgvn5+Sh/XojMVN
mGipnhNs/dpWkQ7ikh0A5cUWdU/VSRSfbEuHvb1ecq4HHjLPu1h0nGWXp9dI1otc
NwGxUTcpITNptUnomNjIawYa6mnmcqoukJIM61+oxuSkxrEyWKCHM6N/cyL8Q5mo
BxtqYCGi25AQL6oPE3M3ObCtcbUgYZVZafbj/1JlTRDipfgo3sn67O7SdxKG6M+a
1LUs0RhyFY9UE+G5T1J3568s6UInRENM9l2SfFdF6+XZiu1xILrmchaWRK5SfcJa
UGATRdsu1mkv43IU4xdZhj/Y5Bve17p/RAD9KFQQp7nD7Sh9uIiehs4xTw/rtrF9
2A/XxHk9O7cU8C9meRQ7fbBNrbW5wh7gGVV7Jw9OvdlPN5rhLLkXnXTdvb7sJDxp
mXSQrN8P0xSDOMgrVnGVG9vJP5nKhTTaQPViJPnhW8p1G0T+KdmDzOOfjifGEq5o
T0P11LGH5CH2i2uGiJ8tCr2LY+25PAQCNcGecxTaB52tCfLiEG0otMUcEPHufWkP
CeLiy02W53Y+3mw3qJQgdPIwz7mO+qN78h2+lCcK5GA4TK0n4rBQpxD0ikuIJ9Ah
kHuXZzyO86+G4e4gwyAJGNm9yps0KQEnIm2sIJ2aXvL4W3NglU5NrtOsbaxnyoaj
s9bIyGmh4gxZxsBatt/B0RVRSufNB0/RU0De8mnbb+lbB6qiMlHPIjGm0lJpli3y
7p/1PBEp0jFPQPbaCELNps2Ahah9LuWeeHMd+a+2YhudX+uf76aZTy0dMCK7IOFV
46Le3NYLNlU0qYSdrYBDrCdvhM8leCp0lE0Ig6ZWTSuECvbQdDn5jM9+Y0r18BoO
GUwavZjFsiEjxwPfDmJnqgOwiaY9r8T2VJ9C7kcjfSD1F0AbuJfL23+URqGhzPbK
w1yRQCBOaZKmdcF2Mf+LTzsuWkGYY1BC2JdInwChKhWL8eXfXvLKyCoCoiRh7UHH
aa1XwRlxEgCjyzHlehmJ2k8MJhHlnHF5oj4ucaF3VXiz2OkCi5SCGqPqLjtbo1y7
qvm+9kXS7ozoEjabjLZe7b7aK2JXWC6RfmdYP/B1c2tw/QY1QjEGJA9R7DtmNAsp
aAhLyl+PRuG++A4/YBrcbr75zT4qamUBqIkp3plHdS+vRFTjBSlNXxkPDMZj8Rei
ME3c2vTa4Lhqe6dcd0nCPwf6uUuaI5oHcXeOdrjV12W9bf2hykMVzhui6sdg/Zu/
3EtMuwV6uUYWKEm8Kta7aTfEr0FHq2sOzkBbt5qX/MUUlg/HmwVKE88l+fbT8zI6
krv2gXhkxB9J3zdAarXRODWPY04a22Em/YgicCooHC+aULdPNlAfoxKkNl17neW8
cgBVfxvaFdEVy0xVwKpPrNzqzcHinQRG4lrCNqNOpOuIQ8E/vT8nrMdfb6bCMJUO
FEvXLxTlTCYe1kO6mzDmi42fIYI0UKFWv0AqrASe7uv+BY+9rO0/t2Aq7FnTFSuR
PctEG3wW6Q+spWqLEyUAzbFKYqkrXTCM0Z97Tg7zvp6HwnyJsIvPtiqj2OgF+4c1
v1iCLS3ZpvFHmW2gm85E6aDQ9KZIi+k67LNsteaQ7Tjdj1qg6KBF3kNdz7fwFHEx
HNSCGWRVQncENgK0m6eMr0V5wGLZxMZLUUIVWICvgf3T7YZKLA9uet+vU7467w4J
ieEo+nkfvBDx5ACvkiIhiIRaOCIsj7Hqa+yccNkK1f13/ZYC+EDkNRvrhtcIatcE
z34zc4BvGpPwSHAUvlGJKPkyX3y5GM0Ppxz7Vj83gHaNmhjl7xKqLeeSUKL/Ko73
YtIeG+sXDQ+2M8v2WEjJk4Z+RE7BWhdSTJg0akptNnQePkG68olqT4KpaoW/pc6K
9unduw5RI7g+VtBO5hpQ1Rv1VRDZc+vd6F/7taM/q6js0xDLYLwteyrnb9i66+R8
vj6N3F1ZWBEB/WwwJ/F5bORbe1jRhNOnWVxjV0bH6afA+USWYBzhpVlLDc+ilmbw
Ym3dgaMZ9rOi9+o/csAJkuUdSKWXDS3QxzSMIOlR2UW6NNlsXtwB+mW9cDTvaJde
GFMFvGgwVq91LV+smYtSJbdS34LGid6dDIRliXqizwDaJDhixYW+72ffSLPQdgLY
cVHybsCVGhEgoCynAS9HiApDSinHL0mAW1M166OsxFmypNgkq85987iuDkp8pJso
POIJpJU9u3Tmb9w+/oJC043MFLErkgeHaSet1AeB48CRIJBV/DDI5XOG559B4lia
dQKq2HbqnE/OsAF+hSRJ2ZCBZ1VHir6h6N/MwZOdQSHVuKqOx6Yl9whD9enatUMU
Bv7GmRHhIaXmdqJyqpEexcADDP4ke66//BOdUlvrVjKevyPUwbQUy1hxkJ8kLz8+
wJOjAuMjEKLkf5bWuFzFoqThINnEXc8V5lOhB7DSCwJUn2SxUHgh4pcc2uBuffAp
cEuUJCf7+ctY4wQEMaW8yk6DF7UVl+RVBWRTDQ7ypdxjPF+8IxQXISrp/oR+kEDa
ue+9GZ+X6OtLl2QA3SJ4fwAhfXOTAFRvNRdRKTo06DUabe+1Y8M2lYFxnyUCtzO9
G/27Gn4JpwwDtNX6ZXiRI81xSHVTzS2Y3uZMOOASYJ2T/ySWkwanrxmLCGZwzEWN
fIMC9DdvOSLI9gGF5BnJEfNE9K50YQkzSA2ch1Ry3divnECzJgqNTW5GmmaJjlEV
MHri+TI5HN/+gfJZ+IgCvW46ShbGRgkh9wBdMpsY5veZjwSHUKhhfeobK2iYUHtU
nz+cPy6Orl1NpirI8TN87pS173iYs8CRgLW0CCCcBoeoDxM3vs3C78oSocE0cS7J
WFjJhTYXiA+sW0ZKc9THUSWvCOYWMY15svfwvo4W4v+oe7jO1T9AyHjdbrvlcMd1
q/k8RWa4Kx51Mgyw9TWP/5rRmboqpFcsbylXpUQpalmDCu9j7hjZ4Tq5k1i89And
B8ltzdMJfszL9Rg++P5WRPrepVEF/ztkAgTeLdcZox7wTUVEzXRm99X+91R2HpcH
8ofpweJoqerGEtD5CuJ9wOW/Dt9UTsYGvobzxJMDfVlUgJW+XXylIoSbgTzaB7FB
rUUzwQi9JhvIDAy9ePgrl9CiCIbndBbQR2RMhPn7iWX5P/Gp5vp2XqbSvFEkYOAW
GYJT0HATletGqtbImiVHo5M8Hd8xVcJHE9NZoGzf56DFfFnSwHMxDaX8V7VzYqt7
1pX5a0WzHvuAWmie4M+8mAqOoXJpI/PJFukky9sB9tu4wRKOWJHoRvxc+RA2iZsm
H90Q7hH62HLVhITid864nZsEoGYb9t7GK5dYX6MzgSqt5r2a/5xzIIFLK6ayjF0+
SaavsOw3hYNRSdbaAkUtKmhxe7ggef3qRI7esYSejuTH9cCBbSeFkGdPHCs5iRUD
9ym2n9Gt+0ABOIhZaCgt41IrPrM9Z27qKWN+oLuGZdy3l7gBw6Iv305f5Job95J+
1Rpn8D+nWqIi87yyuLcaiaXCz16YcmfL67EXibfhAcZzxRviZR40F7MAS1XYUfaI
e+wdG6f1Fr+vnZrttzEmWyEQ+ZEtkroK13+oUb7PSsN0ou3Uz59BBZqp6EL4cocB
l9P0HMrnyyWeaWz/jpXIAa7slqGYktFVCok7pUA1nmwLZr4ZGTCc/DtenWkjytGe
H1bdul2QY2qgs+qK1MiDCzXcEtwKTSzYQmRXszzW5NSofJegdWyEieL3I+pl6CJn
mTkwR9yVfSMqfQgwMufNhOD/NBVM4gWaRYaNsg4+ppbUgef3/sZ3DVSe6V915J64
TIcoIvicvIglnecalM3VOI0l0HB1yNLdDhBTJ5N/mJAFqPtpJ8gvBNff3VBI+RPE
/xlXKHjR0XCvfYyK8nI8sXrFwWtnENUqGuzlGtJyKx+SAmyH4dOxbV77HiLWXY/Z
u45EnTCTVQ0bh5DlkSjOGfNH6OvIEQinjwcLWkTuBc1rkzTvkM0kX5PQS1fODZ9E
esCOE7yTSuMvZeHLn90d2RvcX5Chm0NHszI+ceUCAZtHFeRFvxXV2jkgrJ2FPDLx
/58bYAphww5wCQsomvYdaTXuL+T2LHBhsa3a2Ve4RYRhSpzmj5c7edoxpE59YPRh
PKzREqt7doiw84E4jNz7SZRokNSr5rHdIj3cTtor71CBKfL4Ch5ZnXMok7Xq8vfZ
/EZFltEf5AZ+ihO7OrTJiHO0HowtqtwWyQrT/wX3DgHuzeClkBuaD69VYsp4tAsr
2BlEZz5sbocHi9x9FciOqd5jvAB09v3rjquXay3pHbKxGSd75Yn5IhOmsHtyzovl
hH6NYyamlYmlVd+H0iUOWDXn41CoL4USX0TWZ5bkWoFVKpcnuq9qk5s3aiN03B6M
ls9YEFt/aKYdRVwKdtuE6BrQmsy55r/Xe2Ap++EYyxzkARJYKZvQoDbPA2UduVKy
ONA0Aqqi9ltm/v4EnTdPY7A6qcTWEQjJFZce8iNv/UVZW1bISziUg8pRBa4v0tYO
T4rHS6qdP4nBH+aYpXde/57hJqu/GX8yn9CJWDUVYB8ujXcMjSZJaMhjFWuS8c/4
YR4YOv25II7dVinlr6tSgb0gvW03EnlnctoKTczQaYL6Uw/HbDME5F7HHy4P/mc8
X7AunVmOtLaKx3PsukMYzg==
`protect END_PROTECTED
