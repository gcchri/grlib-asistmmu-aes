`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8u2tyZeS5qNw85QzKMpeRQlE6jasyXLTX+FNKYh5vElCqJ59IrHj3NnaAuDmbEj
a2HAH8ObHeC+OYFxLqfVdVpXh5U8IuFJd9hL/TVpxF5fHX/Zl4cyVO+sjxUUedxQ
fs20nyKDCpfh2gf5YFCdH9AjEwmeR5054VgbkqWOLSwujuer8T5OjxVCW0gpH9r/
CGHAiz7YmoJWSPuAgl5zP/vRLzFGaS3EzmULvyNPdwAsCBWUlrp7w1upC05nigrW
CaScu4hY0rbZzyP253dkuvsKNo4TnUN8KgB8VlhYyr+Hv0aoErVf8v/njlreKpRV
q3nwd+ZajR1UIVL5ayEJugic/9zeeAaGM3AvYG693CbEYZeblQUzm3XbcptXFV6g
KSENlpnUy44uCF3IURhAPw==
`protect END_PROTECTED
