`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
25wGE0D6jmraMGGZxGvRdUNvyRQGFryhuGJyEQlHaEWjew43QJLLacs2woWLcqzo
lxXPsYjaSROaoCoG5ll26cc6SEGluU2tcwLIVyiABV/1MnfqrrvWo7uHLRQA6ysc
twP9STRPIQPshf8yCgsPEhILtEZJB6+tJ34GNAurUqRmwp+b6AhP4xaFxLJmSwBa
Rq63P0jtd9W6dS7OH4xXhOCw+3ozZak8CuLi+BQ8Un0HTOcwDisgLS2NUElXdZ1+
0dTQq0OSI+RlCGiw4O2ykpjBjWg9+gs3KKDj4E/esw/2zxmMMm3icf10PTaHaFO7
yytESyCYCJPfEdsg+Wzs/M//pO5vunkXDcvu1k8OjYCEfg3mFr/zT3mFvxIlA38H
U0XK7KJ163JZpFfJBxlbHHZUGE6SHo2mHSVT1kUBDUA=
`protect END_PROTECTED
