`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWJ1rPKXEiqUcylwjpDcw0b79b6SWk/dFQKtCHz8HZ8UVIev6TxBPLY/r0UvEkqH
nhqf9QcNK4+OrAuQW6JWmwOHUT+MjFsIXnSRJeaVuKDKixpzfmCdiS6gxGQmBbOt
Kf9nQ6aGS1xE0WfeANa/dvRKsXUbIQhjvmLIRRb9WO5kAuUtcJQlgkhFhA8hXQC8
/H8KNPjGTaCHc+hLljdYg2bUijZ1rL/T2Qav1L0aLMelmQo3PKMvMJzUD4z25ri+
ua9E1EtYZEmLeTl2WStHyWmtbDxyA1L2RBjuEPXs/iGiJQNGG5x3UY5xtjd+OQ/g
lPiU8zhfBZPR3i4rFZFn6a5CaNBQEZGeg1o6wbd7FHrloWFF2xZ9NCkZbZIcO0Ij
FbbEBirDZloXsaVVpzxwONuaDoEWT+bsXQxaq87TG4WNveT+8I0xs9EcrHh5gcpx
l6h9XRkuWW74T0xhA29MA5c9yEQweElOttDsVkphlLdZUjn3Fm8fr0SiyN8SrBcy
F5iqKNoKuXM1r2driDWOr34NhR5TA2orfi3+tB5Ea/hYxQDh33YdFjboip65NTUp
EhmDs7jZEnSi/ebEUjTHlVpjWk2XtKR0C5ZqQnG7PuRw9LjBLSQpdSbOfSThaItK
HgFkdbqP585MpibbYElzVV4+4TEJdNIWF31/rTl1zGT/fRWtjdcfrFYgFXbLaHKt
+TEl05CUQojzdXX1+HIIHwpzXex1EjSb2vTd+r5f86v79a7RyUyukBOiksAyPnIQ
bP9Vn5f2LWGdojseJRLYALc9+OEhWIui4zwwdFwnAqP25c6RMSs6k3Q4f0F4GKnh
7elR591x21v19x7NhPSe4/vmN9u7FeerHdLWziA3iLRGwbhvZXoSyLSD209sz+NA
cgximCLMS6FMVuQM0uqEW3zVWoCrqMpbBbZtYjzRSTH4N6/OqU+BVUAcWQIs3d+O
DWm8M4UkwwRhM/HWU3TOCH6d9tgdkl/2ZtFA5E8NyDeZaQF3O+NfS8O8CFTkw8x1
bcrE95F4ZKSkJRgh82r9/Hw8TnD+8UGhMQiz9g3+Kvs9i2x46+qbM5gN8FLYWOeE
ZVkteH9v7MDm0WtCJgJeRLBEb8SRrMI3CRpxq9fO24J17i8fD5Grwb+q/h7pnZ6o
/R7dsnUZx/d3kFgyJHBdFV6+nyQIU2knEcB0qVdXYHU9Xw81rFFvSjAXh08HL5KH
piE8qraLWHDcoxt2IUAU86bCicZV8ydLIyVrKXF8ki4GKAqst1YBOhKUq818fG+4
uYwdAFvoL2Dh3Z8AO9RGtYWW/fSPdt5RasZR8AX2rLwGObP7rSBsAduj504OLTdi
ufKiwIipGc7pAibiD2ziv32EeF4r/XWFY7DezpWLTQBKHNSfZvGcSip6NuDhuY2x
hntqbxzmYHZGK5+0SIXI5M8xUyaOa+aoW5h1H039V5rAtwdzboeb11HwlzQSTlff
MtOZXtXwlJG+nMXbU2DUXhDee2f5PaqHHxLuki9dV/7HfNFMYp9M4GM4mItIl9sw
5JtQ4vlPXxJbgLnxm/WlICfkM00W9iHwMFbhAckVBp70/tfcLKwDkIm/5LCKdn/t
d+MTTUI2J6J+ops30E5MIInX7Um/YFBcDJSR/jUmH/412JSMB/RwOijBnNu4e70Q
iTagsRjVF/QL7zAzkL4iC0WrEvvRO+ZJ9tHONSR4o2Yo499DVbhAywvTvpLr1Kfx
bcHpt118OXW9x4V8tCA4qRKFZzR6EWLuMgYFyXAJAtBxUCpOM9Ffb+c7tlNQPE2P
4snqDJ711nLOnBKpTpLkjmdewfHCLJuxSjNMgNpC4p8/ZbkAtgpY50J7J9H3eGnj
q8snjdBo7HCnqeackwOeMzrFNruI0BCgVMyN85AvBBc=
`protect END_PROTECTED
