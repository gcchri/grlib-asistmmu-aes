`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qB6M866DxL57GOPM0BC2FBYu5e98sUo+46ji+lJI0QqrcKT8ygkjthTUaprNfQhr
fO3AmdhvXSMj+NJfdqal+xnlxpb8hcgKsgEKxCrTLjO3iWlFANcxGeFj/AAheuoX
whI5KCqyRFr6e2htifemyksPk2SKf+hhWvAZtfv+jG5CY1O/Et0yLBn1KSsfQPQj
Eim0Kk1mTDkMOWaOXSs/IOOkQjctXdMJ+dIWCM7p5Gy2PNOAyKAM9VaxsRJqi4ER
op+aYcF/5QSo1zjqrvWs2IkehyFD2OlJKxH8NPAx11IUKvsH9O1vnsWn5T7aUWZU
+0ICT5iGFJYfH0JmnA8FvP70SCrm0L/mRMI+rQf+4S2hvclxRRcEAF5p1HjJRCSI
Ps5bqo4g53/G8eZCMnMNqV4tWXpW+uyusSlkH0Lf9j8U7gpV29jMmU3Uqfn/YdpI
7b+6GhcGiQEq5PTOufBWdWOzqiAKXl8QQha6/2xmdq71w9uoNO3tWFMyRD1p+0g/
gQymBqJJcHVtS/hq5mCyZcUFTAASZx2vDPOnSgRETdNO4taCMD6sIxtxFPNgGGRl
cKcTXLWuuXYmhQ85mVaE0uRPSPly9Fs4YRBVmpCaIrkLdTE9oiB+vOjrHwr94noR
lDJs91+1BbOV0WthrCdR418FAUexld1oDmjO9leglWdy32UMIsd8DnlQjIGiJIgn
FTfFW3Y6TtPf6UipoSPz9AbAcX8xDJz6F3PueZp6I3Rd427Ye9QSYQ2s5pc+Ig5p
I89/G92HmVypyICggLoZSpdgMj2yXQi5koGzfqlh+sD+sTvaa2pRIdbaJCs6aBHd
F5YwixWe8BNZ2xiEKP9iOcZHxXB+DdbrqERprA6V2B4yQS6EKefURhecVT9q1q+5
vP776nqOWiuFpcjOT4LPPoaSqGcbWDJn7kam+zpWgXSwl8KF+lp5J1vw6/6bMCqU
FXczigi+B+KVxYvQT7XHDzkoXptPWC/AVTlNkZNW2/dLmdupiDg8iCKM7S4yFojh
pvGi/jBzeVtcWEF3K6vxBsW+Zx61DqmKLS1eyi3lUxOw9DpWw4INbecoMKcRSBp4
S+3BFXx0jk+6N2aYsUPO9jvNl9OdtLOO0H338TW3iACvSqTgTtme/eqvA+tQJni0
ua/aNxSvLSQ2srHkR78y3wsQxnmfFyBT2AnQpLpjWBBBIBdhQCVK/B+ipChW2rKA
ctLCHzDIurccgpsFU3XnjplSjASPW9u8V9ePfPUFfA+7bxDkvUH2M+j+GRukgHCy
GBomdzsXZPkB2zSC/OxI/8SJusczHhUc8cZnbhY5CleMS6gC3hGPL1gdF1bBuHwv
GOP3Un1rvCqIJX54QDtpW6Dg0WoPCQkcKDNtun7Glp3NBmXHsDaQWCwVsAv3l4a9
VJ76paBAKIQsTuBlhScZEtfVUHGFkOJ8h2SHr+4UKRImceQrDgBWYkez4UEbGg2z
CBW4pQdwBXOkggLV4pkoylUAqPzrbDWV0Um9b/fIRf2QXPMUNEtaqHfDaeQA9m/b
H6bj2leFiE2rV+as3tG87yKSUJjYpcXCho24Gw4NzGIoXSf7kNV9KDCEPl7MZyf8
SrGalkH8JanO35Baw3skSrjvxk6E76rmQWyVhSVlLZZ3F9M1+IpfcvAZp8VCNwMO
G82lUIYoOLAdn6GzHjKfGqgWOHux8BIUTQI7P4lfzPYFTfw4bpwhR8fpvvy4x0xM
f1OXckZuLCL5Jvs8PfMJjANGbyr9Kab4bqaInzbx1dQltpoSaLAbROpE1sNiS47O
H2gzM+YDddDWdMSsBzfmT5DniiPzxmmcfcNJIe9elIayaVJ1PbtGgmhlhfxPRR5F
d9+FJxjcsLcacRoyZWv8XK9MggnJHJoRUpg5GZ33bdN7sbY9SHwdPWlM6Gvr32YR
K9B1a1yiR/6vQAyhk7S7LD/p6CmwI9A8eDa5TC7gHZ+G92dZKPSMNO2Fa6cxc544
CM7sFI2jrg7Lc5scdfOW3SY3aybQrYeqTA9MdVgJX2AT/SH3tSV0db09PP9jwtYD
QhN0+bNoQiFLMFrkXdDb6jQcvhj4t5I81oQayQ4cqmsfCJ6bigqFDtVLIaxeAF+G
I+rRolrx4obZ9Haf2VXo0A1WswkXRRjmN0I3ZkWRRNb/ExWtLNBRZ+CE210ErjV4
heXAP4lTB0wvGyRQ6Hn8/e6aTzop6Xr2xPbxGtzbnRy7DAo5WMi4G06N8jA0R7FV
4ymvGx8EP2HOcOcscCTBcZF8vj1w7xmEnmnrJ7en87c42L/7aMgDtCOR6HYD+E0q
PKN37b/ERmHb++TM9K81tqc99q7/50CHSvgH5XhaNfdBxLav7uYkCfRrB21G0SWd
xMiIcwYlkguOpzpg+0+yuKdtQ2UQYzZyeaLLKEnbQAb+erud6dTx/7hsrdNy2mgA
3uu9AerFjxBGpVmHHk5M9SrhN+GVJz35a+CZdNY5ydR/xneUvUAOB3vs5aKPhAIE
VUz/7TnK/8CoLDjRxqGvLiEZk1aKbvazba/IocYHNteJ6zrYYBvjar5HqkKsOtEH
s72lbX4B1FpDXjGL41EXYYmfiaoZxkZQWMMygCuy+HINHv1LaHjFKthJ3F59LLRZ
Q1p8jkhb3z1xao5UVaYt1xV1td/vq126MUiM0249XIqep9+dtIDJuNyiZa10pZF3
3K46YfODByNf/YAzNzply/8OU+p8YyEtLQ1S7+hLfBJqiPB2veOSy7dDkRlNUn+3
qbtExESNUUwSjNTm8YuzQ7xJ/L5kcHg/xYvPaVTgq1eC4/uIuwwCXQQlN6T7QAwV
hGDDQLemJ2ImVGSkBHhpHcm/lP1Yf8fc77Z+Q2MIPb1eVHbZ1o1Eca3cSKB85dw8
3RxmqgRG5UnBHsuiNxz/fiKk+QY9WYApuUrUkHgPkNCH3+R9vREsWDDmHkrIIrcd
yblvCbEiACVnco16fzx/UrwC6lC0aHl0XeTSI2J+Nwt2uK8PJtEM1xKGvuAMAk09
uWvIuIpALeZynNfTikXRpA1oY+LF+DXK68eM2irg9DKvrk9nFvhiU2KVbjWvQexU
wG85INdZ2rwc7bDrZj8jUKqts61lc9FCRF6C3g569wtpw+iSIN/9v2Y+1vNc0GNj
vuHfNlWnADmvCCgbUN2dML0hCGFSQRJY9yaXYt4eRp8Ms9EKk1S/clbgXiFf+lLt
gw2CJ5l+j9eQwrC0x5XrappSLokcJHuu+aWuqYB8VtSH8xA2M/8ENHnE5TSPjOwX
2xNj7JouWJtNXWeU+N9WBvozYOflL0q0MM1LJjkbudbMDf0kkDMUZ6neC5hxSjNd
ILubjY4OLV9Oq73DHMHkM1dJuFsIPQwt/lGx8llOGpx3I5eUQR0zIL7EixD2MBXV
jg57s+JVPQWGSTYKRrJ1r9awADpOlIKqZXnYIGHCY5hZbbvfI6uYQAqwA937+u+b
zkZT5+eTecwuQwhKkYZWR8SZLXLMFk8Lf8lYhl1a3cgsbsyN6ova/9Pxxf2gXzR/
sOhOmmVagHvrmotVqbNJH4o/PDUpBf1JMod0VrQp0hKP5TV0HMU41JBUxQldWIwo
6KurkhHfYYZIOM9xZsYmDdgWoCxWwWLp8KVFODln4UJg8yanIiTSC0Hu+D6XAVwL
/L+0WNSuyTjsUMmp/M1RJcsjJUp3tuw9bfSfAw1tMGO8KOYfsxV6fqOV22cDT69p
Z0S6TH3DFrHV5XQ6byEcPpEAaShlV1Ygqip1sTzvnY2Nsy0XRQZKI99d//6umWDu
oFJt3KSPY09VXgljyRUMXqXO4gMYJ7F2GfquxtGCvvJqduClsmrSJwUZ+7To0kVu
dGjq7jRvKZO0wvLEaHDW+pOgPqctLw83e3zfDdV++dF2Naz7VRh+96OgWCMgiuqA
HLVcNwWgVEZNBI0ORy+ikIbFgYbRCOWbhyy4iHFZPV3VQec5RknErdBYr/VrBQuQ
esLvX4DZn6VBR03MHtyoxQiKOUfE3dTW7XS4ZhlasBclIMUYSH+w3XIW+/qnCiFf
lPJP3vjqLHpkHRuHBvzL2JN4bL8Un8+0JcGuQVNcOVTj9U8Qu+aMBDKXqx2RLh+c
0qe+gJDvusYSIA0yp1xPoa9etUpPj/ItYPVJDRk5mLu9QOgZMu4K6q+QTLdvTPY/
lQXiDNOABnwzfDwa1wTFtsWJFXBgEUEXZXC7bsd8HFgaRnwj4TSrJ7sg2A2RpjtT
ZTW1ks4H+jwyHUbfhgBSfMP8+Se8B3Yq7l+W3IMF7mDC7HFGVVaOOpUEYaRR/Bhy
5mSr7e2eu9cLFsa6Y2V/rQ04BcAF4hEsZ4ytadyExbLvSLoluRMxy+a+7ef0qHhV
PUWEKClnEg/wyjly2ynV44c/WcOxqSDivor0i7gugAGwS328DXQZve64Nc+8uaYx
ddjRVxQ+G9j9uKCxkXb09lS3ittQBU2CNpU+CvQz8IM43IfMXGei/yyaTXsEHodR
jdGJw9VspQgFLPJpWmm3nP8NSGt0lKSeFnHxUD55HqF+kWa2zBjPURO7q3nlGFNc
O+9GnufrebOx3TpzvI717kIVShIBPxLmUICs4Q8YT9at9yImEIHrq/+CnLTK39sQ
w3ujLF1g7VVhpo2yqvbiHx4WW4yV6K9tNzyFgOJYwErDYM2RNw+r1+EmKqmJO+p+
TZjBP90scJiWU58htzHIkZWM4Zf418LV8rZFDEjb7FfWM2c7vU9dn3OccZBP/jXf
1PyizTYkDejFMrfgxQL1Yn0nUdoe27NClglNfL2gT68SP09Et6LHS9zmpXupyxbh
3pDYyP+Oir+3e3V1ORtOh99ZudsRAuA7EA92AZVyHM/F+aaPAYP8F5GSwFTgfqJD
fJtqfFMV5QzV9tRv9/OdYHClcIXIJvl1OkEbZ45NB/CtxNpGXkgjgmMqT8TUtP/I
Gb0AxDrdSfne+qu6tj/ygIwAG/ZedMUV6Ju7qdUKdpoJXPXb0mKZSi70wcxdSTws
QV+uh8JxwM5giJcErtLuXmwFc/s884Rw/tZ1a5qeFO8Z1+vwpakBLUKZVjSXD6YG
Qk0ELo1n5wtFMbYlzldpEKK7imtCVLBLVJcChvnXSo5uYaLfFn1g17hs10d1JviM
Y8rvQNVJkvODAW9lZIBxN9ChV0IKjI97EhR94s+8BMK4mWYCT8HqDfD1f22XJ4ip
GjELPAIstSGm117ftfdBJYxrv+qeZEkalHXyT/vk2/br3siKYX4hUpMJbbmO9qZI
75QRCx/kipH3EiRxIVXC4YisXI3qFWSayajBYTJU5RmaLy2J19p7bPIfjsA7hnp1
0xQABody3T8Sj8wyyeU/8gkgq6+pYWCDaR0UHitsivthqUYtPTftWnuH3GgSjeK1
JjMnXy/zvwFKrI95jag/2VAzlIi7D+ByN49OWMn2ZJlbMVmm7G2v68HDIgDmxt4H
QdI6FhOU/4A7eZiR8bNLzcSpxlIfJ+uZ22yPyTTwiCgZFLEtVcqMCGMx6eyPjB6a
bGpImGyOZIdTfgFwj4QWcHF7GzF5mxoAGUxhWx+Rlyd2ms4U5x0QfKWj1iIHb1XD
F+OnGrJWOCcyKqEsM62OIpUOUMnBuDI0FryYKQAwhNjZX/iDoM3dTUo+/eo5/X8p
AuMUmk8xYAqyyQgNfDLEwJSIDZwgJzAN/BJqjgN/rzx++/2JqoOL6MsOqHoZ/9Cm
Rbu0fF7+0pB7BtHG/wusiDUoGXhyOSYNub80Zpjx0x/YjPJ0t+tzkRx0sXo062f3
gBnHkGxju264dHtDPwUBkDI3/bC0WjSNJc7E269779n49ZJ6zyKgspjXufA4oeDV
5YgZq26/kMH17YN7iUBa3fPd7YXBnVfYBH0JBxrjVP6nf/CWQcpRCyIO8FmFGLVY
5lt5tKGMG34Y+Xxm21aPxWTBui1fy+hQ1JFvVwibjpM=
`protect END_PROTECTED
