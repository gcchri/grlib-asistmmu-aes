`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2xmpaV/W2Ihukgb2Pzaf0WkWrpIqO8ilYtxtcgz/dAybdNV/AioedggQRn4oHSM
kBL0f3QtrXgT6nvs6jXaFV/MHxV8uBJa4GrEI7l3mvdCynh/eu7VBr1GPG+HDFkj
wReRHiDvd9XdczXCJcXQ1+pyjpCCJVI1GqtuFGlW9JNrbCfYM8z1kL+hh9StHbnA
itik76oB2LyIxKrs2wm7FFgB9n3dAM7feOZze50/86al/zto/dHRPzWyb7edDELj
vlHco1hlMgXVouj2AMt8GPfsFJ/O+3m6doT/7A8Ln03/wwxLUVPb3+kyKLnOXumy
6WzUZPdLvbXq9H5tVQ2CT5JeogMbRQtfVD9CBkuvEZsm6jfQyWyRrRtVe3BqsZUO
xvZlFvURD2JADoEFG8YyEdJ1pnehJaGqJlhQay1+35AsdFOhHJTsv5OAbzvZJL4t
UkRW6w9CAg1eYggum9VDqRZbuCwROzBU5BgDrj2tqJPH0u0YqPcZ3kp39igR0uRM
PQYtgsYIqobgICPj/6B0WJFCgLUcqnEqGj9QZCH1mob8Sq/ztaOnsei2Gi1dXhHe
eXQYNzeZzIj3jSl/QgIdHscQcyZBKM3NtSmqvnCgFfZTXMK55wzG9yd/9a60Pbnv
pdEBRX+ypc7Y0NGfb0d8Ni5/xBuv9sjyEe3JKbN/uA2eNCKSR2oeeu9ISiFHGGJ/
2QB0hDTzox0oKQ63Ba2W//+WArdfpMd7E9MRS+M6N8Y=
`protect END_PROTECTED
