`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zfEpI1ZY+V6a4eUd3rXpFRUANIfsdyKCIQqO6ZwW4gCILNX+P5NWTaVAUFbFcFZc
ISatWHmousNOU6+hgc2hXm9cFgGMiMBxII5keRM7t+vJW92v9DZb4IKmfJbtHnZ8
6x2dMncBdm6NDJlv1voixjph1p55WgB+Qwbt4pvmGBNCHxtf0bFlBknZ5VnoPrF2
fstVYgACZP42WQLP152Mh+Z1YDE+adbksXoDE/1q1g15siycam0QQIAGhawJj3Nc
+qnOCalOugLDXM4yWIq0l1jacsL+eMoVpHMJ7qFmotISKsHM2vZ37qDvSBOOr289
uICrPLAolR4Hi07gQj7FAgfj69nSpGzBU1UU+ydclYKYOR/iOrow4Pe50T/EvYSX
fKNdgTYsicinENA2vxZOcoscoBMAhEuULRdNk3KM6YUgV12CfjyGsbuhq6Y4aSEj
OypWQTtjkOXWsRA0OMq6vxBuyI5Xkjaza0JXbniun78VY+FnuyDBPPlZ5vQlMoIv
TM9R+NBw85GU7ob9tv7CJKnxtqFUYXjeX8Kfldy1uyACepXOBSRbCgbSTOkt+NYp
G3Zv9Pzcgg3fOLFhi/cX63pAhEawAE+irBi8ws9IBTjBhBNTzQkKb6sfRD9YseWi
LukRE9luOkQdiBOeTvsTpjgys9JGj/c7hu43+xTxKFJNg2Pe9lpEBnsmvrqm5igD
pqRrsNCHnk1bp0NLUPsrEl/8XW4C7evqwxxEVj+2fMoZ0tjOcFt8MHg5OaZVmBF1
SFcn0qzgLzIZJcjq5F1q9tP6B30Oca7gIPY5LklAxcWuM0JstX2x61WYKvop5nAy
lICt+XoUz2BWRjylYvdNelXw8AVG2LrJDf9cpCp0H0ZHH3E4YNI/kdXWN4afSnbi
HZZoJFs4SM84ocsHSsyd2mf+bZQKr0T08NjrWtvA+Pfzbo3LGJu9oYBnNkdLclP3
35j3T7JcvUtLBXFTOPyuxHOQnH1TrKa8Ic0tUHyosVyO9+n1oPZYulGMQ0/vuOIt
/kCvK44UtstgGj00QtIHtUANAeGkebJXH8Je8ryl07SukKS3mPejbctEjuJN/SId
v2sYi5YMDgS+DPZFK0qCqBpb5YhdKBEgh+nujqIl0ak8inNJ5tcou+ZOqrciRalH
yRKZ0Si7rxKvylbK/nZIS7FwkNFHABmXUqW6vm6BCZlw815A2waQkBl2JbWwqaZr
Wnma8EqbqZnz3nc7a1+nHwQKk0pW+Erf8MVSHBUfVaACxLYGw8LezrkEGTB7A5K6
Dquqoy7o/aeEZ8r06FhQaiB6mmEANen1WQt0+h09ZOk8/zSiMwy9rfPiF8oMj8wj
kpMqRhduQJV+zwsjyYWeMZJCqXx76MYu75prELa0FGtI9lSXiCM3a0h5ugCSsOct
OQEoDXm67fbguWCOKJavAmQgi6g2V/0L1fQO32ZkaUrSZEJN/oOiZqw2R3pRkDGa
EFc8ziLLOJ8PQgCBIi4/ru8yRFcklUp48nhMfHqzDQL7MPQUiM4cfoNnOmPA1g9l
zwf0VHkKJdjr7D5cxjkcR64RJb4NSgIFymA/RtazpLDkj0uPten9Lm3xgsnDYIf5
gqinHmkKdZDbJ1/pmfRD7TwIppgUu3cr97UWcnRBQ/qIAFtbUEa0d4M5mRpkasR/
vWIwWtWzE9Otnn2SDZdRusmjKUUhb3U63Id87YGoXBNR0SS8jCOqEitfbWiogfT5
YjXjHfESBG8wh5ND1BPfWV0yvAZx4FW1HiMSP36yjOOAbMCdARP50SWbDBeXprUZ
JomMTLqdQNr++LNPp7G8ObElj5OiTL1NNQDHono8Gm1GB35cPa8GIur2FNEfLGWK
cprZXqGqtFu8WZaELOEXpbux8D7zOkIb9LehZ/TzcUVnVC2r1V/Z1n3stZ1yLTrW
GVwZYW0XCWruQU07FPC7hR4MjWlpY/tK9OlHxEaPLq9a2AaLw2H14U62Or4SEvQ6
fG1p6BGPvPlJLgIOLk6Dh2kAWYzeVHX9KW/aLwl1v2SfYYnx1semhiGwcZJoOIXp
ZrQt1vYnPDrM671y5kkWaMQehCNRExSB6ERYJJrcJqDKcNfaQ6Ap0cCiNKrtmeLX
jcfgAnAFVsGHwXngD1I/ZIygJzEGmZMMHWIE8Ht9AADlIeydAvXQdIO9+VR68u6B
12eg5A1+daC/SRX3N8yWssLPaGqth3RHLW2BOZrC8QHdGhs+fz5csQ/6jo34qdQ7
ZIduBCyw501C3aOyZU/tzRL/i50qh4hvuBF+d/T0SzR0r2A0c0MuvqsnkQF2acAQ
Ugbqukgq1n+HbNPFwYQNpsEASNU8j/8mn3p1Ma0L9RATYS38WNI+PZrzvsF4DYZZ
lQz4e7wIoI84HKxw5rv/HYFY6MUzKVyvvuBmCPS7O2J5we50hkF4/eDNSRZn/G9r
Xxlq5/pvFdbSXN8lVjSFbGFROce7KjyE5N1/CFQyZzkR17TSy4oe9nFtTLFS+hqs
xww1JhXEOyCAemknDZWEVhVtVWTNMiwxscfDoJrqNFmJrJ0XR/t2CBJM4lwtd74C
Xznc8pbH2+SzF9wij0KBcRWi42UEsBdNHqE7/dMWvOBzwAI+Bn+SBMQ7hjZFyjn5
0482Jurk/hTxn+4HJudXLjVRTfQDJm59zc8UmVe/hEeVbbQRvgnT1g+3aO/Zg6eX
fRh4g1GILO/8A3rEaxO7Qe1Adi9g+uRESCDQX1uYL5quQujjXd9iqyaj9Nb3z6k3
a98yBlEAwCxLRSi+ntBozczaMt6p2si4Jph/80e6qQ64LOjGCxSDUlurGHVfsmfN
7uybWqs3B1++hSMW9PRTMMkHUp+jDCmTT5Ud+vdVAKKqpOwxaAUUQvh1WjfuySRq
1GfnQMczZamUuo3fdIewXpcD6wmVKiQpcMKarT87E8NVjDfVx8zXoabecf8xkarr
Zwc6rPpfJdmtD+OMcjyhe2J6YLF57JG/LT7EKjCa1v0By2nZ3HWAGmMo8soeZ4ot
sIFpRJS4fuee/Ng6AoAP7lkTkznrWZWkWsqi6CK2bpeQIvxFk3tSE06GuOLBoyke
3eV8RGXn5AJ+N1ULfPxrVX2Arn6Nq1VJkLvYnoCRDW6dUZ2C1vWnvjL6jgRoqL1v
VTAeltRwN5/7JNtjhN+MHN8wbMcfQaZBGKNuMpgcwv6Qey9KzW0UqJAEkAfipF1H
Unrb0T3oX1tOeQKQM5JJxS4pcYyIGYPW+Ai4sSOy0XQc53vL9DH7phFyBZdlGVjh
IFnh2BgcTHALruWIJIPVQdfboCupOPtwFnlHmUoIR0xM4rpuM+ToWK3WZs7Vqyyg
0s8yTfcsq8byPcHsc9hXf+tQ6zr8btJGwdllG6B39VGpb683g8z6qrMTobreA1at
vHmNNq5Ree+N4DANV5PuC8lGZkfwJXmU9oE3Iqy2YBMkIW2tdS07WmX8m3vKY+Kr
DIX4u00nV/38BmyRmgIQkO9UOpFTJsyQ3QvXLpIe85FtQ7fCwKH/M83/a95B4+yK
xoqcAl2IMR88c5cNJTxCTdBieMR+hFr/tryycB5ngxLncw9DsAYVBwpWGF9jNBsu
2efDZ84qbwLXllhNJY1pQYgXt+gl0jxM58cZ4u8yzFatBX6STiJNji5QfNN8oDp2
O+tbbn1DQLFSyb725Qdaufvp8kd/adckW7IVjZdNscJ+rOKW0L4P4WMQp/Oz6o/J
pwUqlpBolta9QqIxkYTpkB/V4jdfYLuRTLvKh4i3hhzBZpYYGqDq2g+CpQwXLdcg
rRwcHUxAeKP2BwiKlr/F0kDJlRAgV/iqR4USnEX2Be9q3Z/7bcbszk7ic/+S3WRj
OIVJlepx4/1thk9DEkrY2uYK7MwlwL91iRIvGQ+85MbeClJ2FAfmWTVn8guCGrrK
nT+Rt98D6xjC8ruxRHKDaA3/mWHVMJsRhBkDFmqe7UmR4MmoGD+L3yXxnNlfHA2U
R2pFsDqWyMPilSrcQGER5287MpD0GnEDn+wYcmj267S8iR3Qh64qOwpE5lSleHXm
HSmZGzf8fTJTX/2zDIRFhdWYfhMbSq9U1I/uGQfK7OlrkRkJCt41HWPkLbHe1dZ+
Ym9eogS64psy2PCm/Djc+Q4PNFwf9i1tzuMpkFadveh0Ix6MBwO1zvDbvAZkXZmP
rJrQq21KdRsdAQI7cEIIvQ5d8QJlIlBupBsvoyCyROIRvSVs/+C4/IBjk6gWYziT
MFyM2No929qvb1HAj51Y1aJggHZYLIaCMoZ3LMcWdTlAcMR+7nj8uR9jVURTWrZ0
CUno3/3adqQ0i5cNKd4eR0OZX3GArYZoTd/PNHHWXm1hwMfHDQU/k53mnm4bD3Pz
UKP0XST8v5/CELELH/EMovxWICHlPV8iVQ4k/ACkceetRAhn8ydRM2VaNhyS+8KA
AZn8PWvkiZ5AvDVrecoakJ2AFTeElsnE8Sc/j06PcTaJiTZn65oAKMJ+EunpWOpR
YADkBCe3p3LKi7/TGxkN5Pf3fhup1fWZEcmMnBEOOd0/TEW3dufYkB43xxTqu9f1
unW0LNlsLAZICbGNuZ84AeIZQ+ZUxSA2DeQXrJTUxh/lhPUtVUJcq9ikHQTC+zRN
zvu45TPusCF6Egfio+GA2DqupvSiDHfWAvqHidjwfzg83xVwI2AQatFl3q1+Cwda
DKMjWYLAE9NdBtCBUAIKTGQmv2+kO102enzC3i82QLvKnu4nxVEWFdP35UBDpSfT
le3bFU8Pjiz7r0MRCFqYRq2z+9UprWerrv95Gp/eSxl8uLowCHMjrsbvQTB37IDk
mIoJhUUkySUu5dx0m3oqrvRqUWug8OvHrVvyrh5UOCmzSl+R0zDpCL9GVRoMNP03
ZrwqlN4eS1w1E7m4jiGXqyWFsq8jj6ItUkeFxO620rw0x4I/kYZ5ZMvXgtZzD8IA
Hg8fBnV1XgVoKMNgVcOYEKaxTNffbNhgyndgfJ5Cx1FRql7TB2UgHcFl4hjWgoAq
U1v3FZ7AF+17xOSrZ42OkveJCIDWXwNyVkxDAXLMXSEqPrg+xHq/6DxKvB3hvhjB
DUwJHLXQ8k+TO0Hu3z+VdPhthp5RScABh4vcB9Agb9GNoDVH/+whR+tBpQickRie
NxOWJb2pNanw2F2m1gSlWCbL1QS2GlnQU4PvhH5/khrRUCtcj2UhGjXE6+Z40wXy
A1QNHctDoRslVAiMlrd5NaESJCEdh8gb3EShCy/F+9TGLqF99ohIwshCuiO6NFUW
yGohZsDy/pr1Lfkwsrc0K/tmMFbobw/fmL78kafwu0EhHpz55IQzwdfKaQd1luaW
YpiS1HpYecvhTvSWtqUoFLDjmOuXrtUhmLvSyeheNG1o3h5z38b5ziipAp7sBCdl
oYIHO+Jl+JCeMLCzOzTdaq0gyH2dQN9nL3SRnUcWItDQWBqfn/goaC6BeDYi2TsB
/Wv97kC88jaKoe8FaGshn8/JgN32f3yXdMfs394nx8ZuOwWHthCd8Lb2HDK96C0S
owoD+gPiSrP69+9ntBBP9vzrGzXWgyouwp3Zxt1j0MKuelii/X6itAe3JaCL+ofu
FOPvzQCijWkBfy2mGLpfIMle7EqrqsQwODs4FejOpgy1iHC/vgTBfnE5ya/l3bT9
i9YA9I8iHhOhSHVixevMFqk5S/xNCKUbhYJLMLNMVNCxcUAaRsTLVK/ZDdhAZ7DE
9jz3ROtaCBcI1AsDRlojvXMNVEB5AG9gybDseYw0XCWj8Cz8PNFY0bsfqOhszAEk
6EJTTL3nBeqp9xi0pSbf6LAFtLG02Pp/UPrvXIwx3XuEGBwK4Q3wOSBY56DXp1ie
8hc0QXqUGoE68GqyAhdZter2J2/9mb0u5qDmNfGoc5pQNTOxnNiDH/t+ynDZq0dT
GTbB5P7fUb+mrCgaAkr7Ddcyk1NQrYgNIitKtY0mJtwDnw2nFGle797F6n4yviHh
yzKiw2ne0W/G3Y/ivgfNQDGTIGEVaEaagFhHBnFZJ0gpErcpoQn/Arm+2BGgpIBz
mF3n9+wLBq8UiSISwcRPHgMtqMTIKtA2UP4BAR1jn7h63Wza6LbKUkZsqu0eZgOO
rRD1iR7n6jmONi4evE11e8leqO2Nuok9hZjkTJUJLTIcmlBrAhriTYtUcPtrK6k+
WxPL3S0YC13L6pE4ogkyngfKVIhFsNhCcSAcBYT9y1dzGShLpXZdvZ/4fDG/wQHg
P4OjEjESjosEp+JlWcTt0+v6DrxPy45LjV8qIYUGvpfuRtuRo7DB8I1+M+Kj77BK
D0BhpEB2vcSnwImChnLoBc2ARwKTyExAZuGPUwDe+PN3L3nwVMMD4SK5M/LDtU2g
IrETtVNPxSWQIhIdT4TV2+kLh+EpeSFX5XJUcjXWNHr6y/JzPq4p0XsT6WOv8lYD
ppy/6LfdqKs4YyCuEaWKqzAqFAcE8Pt+33Q4ZWC33QhXP/+62QAHa/xN33FSlQTd
AM5MkQurdjq/fLCggy9K9vp+gSg0IGejBzYmDjGNdacC3wRt8NM32ni401FDqJnw
VlP8XLHOjD2h2kKDs/wsoIi+gk/mmT3jd6K4ENySgoxDxtOYKDatVa16Yuutpj/y
jG/kDdccy19krjiAMbDjQ+QBfDo7MxmD7zNfrh9gzWes3G3eAJdiTpoIDSHY3v5/
gxf2iLoxLsS5zfQnqWf8zQJaabarRXKuMsstFx1stGa0zi/DjORNNVZG1BCjcdGa
0GeA9JlM8gkaEH+wFY0YMNb7iOTlzDDz5Jj0VTzUuL5hDjZGaygyc/Evsga/oSaQ
iR9uJrHAoz7HbPCeSU0TKXTwDXriv4a6IR7sjPCiTrwoMZYXuT0WH5jdnR8KozDn
EMUyljvaGAORyybmIP9wwwj3zxmbc/2LRiMlXWpisnS7jSdnVmCPYlXASRWj2ioy
g2/6vN5ss7w8u+i3ePkQJ5F82Z+bKA8S1NRD4jmOlj2+Lxmk4sVEZY3hRblkIf6r
PU9qsKZ/7ddx4sffehLzEOy4W8Vbp697QONv5afQ0vMrGHCa7OY0KR+p1l9YWbNb
Vc38ANSiKIudAdVN62lIL3eKiH3DfMZmjAwtOpXBtaep5MSev/o5iXGLQFg4RZlB
x2f8EIG6sDoEMuDGe/+09yVRVH4g06lfrGqKmEbzwLL/0kg6AGi+bUNmHBJIbXtq
TIIAR5q6vlo1zMzXJRRx9HV2mIRPmea3NszDS6k+BFMM+IY9f/mkSFZS9LD5O8g2
Nddz5MXuMFIvxqRwXel+2DBPlRibnri/hhWmpV8LBj99o6Z9V9zkY3Oypvz6Wsk6
8KBwMc0ZctFdP7Pe64cOv4kD5fasyD+jcPDVpjdTgTFt42/dDAVxpbYC0F7o5lo5
`protect END_PROTECTED
