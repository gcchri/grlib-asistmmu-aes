`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hDmhczrz4LCdGCHA6j9roj1pXLb6ssdUSvGk9zPqAJDQ3iY9i52CNkxev82gOfaJ
Hfkl0FNO8PkYV0+Q45qLCUK9pUExrAwkz2BMqZ/1IqR6gnUGLKxrhvmt03WB2kWC
+c3y29c7HHfKTmKK+F/5+OTo0boEy22EXMafOQcA2ihnnoiYazn2q9E2/Mqqi7iC
nQsEWyXLUTNNKBEcjL5TzxlTEQiQylexUGgs4VibOrabuiHrlGcN8q6B7LB+ACmR
M/UKRDm1W83g0c0Pw2BQQqOtuprhYiTkvIRUvIUzzgb8Qs/TkOLP4RyrLJLo3plt
RgeUNTfKUVNIRv+N3PWvuKg9FMkBpk2C9i0c7lqaqpyWouwb0FtMgbEmgFIUAsl3
SSqkH5E6M9ao9uAArX6gZGchqe0iIHdXk4jgHbNYhe2fC+vOE3g8i17fVTmTBrNm
0iDbFyccL60esdEEhpth45RFao8m2k0RKqbqz0FNLbkb04zF8tNNDNn2MZR2LP0x
6l1/aHgVe/2StCdpoRyHzQnT/p5wrk1x/3d9rq0r10B0GHmRh15ce9+zWDa/r0Fz
Nv5R/om1X7HQqc9kqNR6qAfIP0ADedJZyAMY2rd7vV63nNfB9m8R0PiWqoIXuN2R
a4/8RoEsRvm9S2cgnJq35XaIGiS637TlEDT1CNH/gK+YAiby0oceYVgIRsBcpvI1
NaXSAvzsZrFu6Tyi/E3ULA==
`protect END_PROTECTED
