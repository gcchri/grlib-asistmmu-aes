`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
atVYHcvACpKseB6MOoymuGNkxRp508uFC75HgXQdqTLgiSXvxjtDfUwzGv+zCU8N
HZRzZATaqbWspqkEot9GCYmeQZLqbL2qDOuXubNcor3wXgnRW4sTjOp3pe9TccXH
hUYs/6jNZlNkBkXOYiTR4s0or0Rd8hdngG4xo+vA2fp3ICYqAgqoITkXRXUgUMvR
tK5VM22/EHK1bTnXZOFol4qD4kmcxOLif9/maKqYdZC7YQ1KscdsQSYakD9rqRc8
jKtSjagOXs36Kdo289K5Vl4cmWJLFUSGp9QwQGe50UAoK2Y7zS7SHmeHX3iJr5m7
XPuqp2LTf8zCnGPknN1FTZGLU78kF/KwIlqTxjKQP1e+f1CEJ9ZVqd4vUgTF6s+1
k/QXgGYSoBebiqa6hCeIAENZo68/BleHR9/v4DSZNt8H8Thi78AtC29NuLToEMbR
`protect END_PROTECTED
