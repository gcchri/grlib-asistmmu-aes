`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l6Gy8bsXXgFZ8Lt7GFdg3jeY6PZUHJLbOOFkA6i1qg0eV0KRsSWA9rWdCPOw8Xuf
MXqKeMz0fHlZXIu/1RJQ6CnrrxStThsKCkS9w6gCzCb6LFEDulQu7m7bqIco87ym
f7+A8S0/Vj37RRH3c2fK2ALmx38nGierH7DIfFQBMhGyI8jHtZNdYeG68mW/oVEu
SqwZqVMuEgmJv4xP3yBra0fK2d0TUnkpWklaXvmltJCJrMqwAF/wk8E2IY9rO96A
ne/siQo7OfiU5vn6TYzzHAll4FR9Be2tlGI68XqKqiIwSR00yjX2dNMWNSByG2A0
pRrBT/ypiQLkTFRNykMpkL47qTRQtDSFkxM12ndbYgBKvEofUGBUXyWnc5XE6uwy
0S1ZU7XhFloGE50vyldG+252pckUMMaryXCbEWjHuwGz3yaVQmX1HFGSpr/ImZF0
HIRD2YdTogckFMaT+2+eZKTrhO9VFhUxErnCobu+3lGUKMB/WeAj+ll1fT0zXxdh
O23x342vSn5+j/UDdAhlyBSngicqj1M84U2SeZJ+JV+YuZgD/kJRBvuZ54xP98kt
4/fHEwBHpEYsfLMiHgHuYd62qG2+X0kbbbiuusqyM6riM4hJdXKNob8+scNNCna7
NPbFIO+OkccWRTgCuKrKpOA6XGnBLoaI4UCOqryDw2CfJotKuvIEx0g9POTf8JyK
63v8+KF4miRsSceY1tP8Osto6FL2MqyXXgqWLmE0y0aLhGfuCxhT4ubuUnqMizWf
LYYLvAdKLTdoCnQmKvsb/HkpNKTcV6hep2JJRtSLQLUiu9eyEhdqbYOZbAPmrX/d
X6qMo6LuK3Z5tQsdQcGrv88YFIIIq6SeMXCGPCV/W30EkiXDE/aTd5oHsO6JfC9M
oAUpKlemSijtQFC9gumOQBWe/WTG5K+j+PV+71MvG759umuW+AJBySD/fbudwA0v
zaTukr+5mYG/qoB7/D0xpvkdZHNSyBFTGP3wdDQprV+GK99jq5Nw5BJ64gajH37h
0ArgzUmbrpKPwfy4UiBZZHucad0lR+5FAoG/+/Brr5Uebg4Qoq0P7FR/cfr3yt0w
6z+Yzb2Ex0CtcdmRtqO5MJecssryOuVV2WlL4atGNcFAB15PeIDfBRB00EzJNiQR
WTY/dVVhSvTN5r/Mbxj2MQfWRKnQ0EsflpQvtUMW+b39IuyJM8sYumtQXwZGdp4t
ygLci7agkVPCMmcBvLLDuDm3amMrBqE88a+ZNy0JZviDSyVpiqoglay9p7uYRGlb
sQGfELr5bPf7QkFHJRlPSELclRWzvgacEyj52ipFgr+igtenBoVqcSt80IxvKSpl
uRtYOQoBpRKTYYoA/ZV9Hk7K/QKRNHcs9pZxz8VLrlsejMl7bl6pAuwnfOlg9HNF
WBmGdjFEuSJtnO+x1z0JMb5w4T92XJx5yw2qmtDoRHlJhuVoC+KaJAAqNQn4Inye
SVPaNcR9V7O/6JDnU5v1S16PCUpnDC52I1FtSgWiC1stOpRLb3k5weJsG0Fxz+ix
Mn4Jgyhv9RqzGomqRVsloIvOVbM6tc4wplnqA3qVs6x6x8iWEKY6StNztmRNsmib
NBCVpfI7M94lcqBsONFhBUUMnkyWuH+ZlnePrQ3Ffu7fTlhmRGrld+5FrootZCoE
D93e+SqIeX0PRgJ1coQ+uwk0oh+tHuak9hbA/Jgw4Q5/WgUw1p9U37diBVa0zuWi
rpJ5oiWx9MdDcmcWouCSzt4zoV9YkZv600fzV3TfNSmpV5ZYsXzHbmh1a3tFOlA/
bLFgaDWoRYbU7ucNsz86qltrTkFP2yAhNA7FcTRltNyTZs6gJFDf9J7HYj7RlKuQ
qavQs30L0vYvsCwU287Q23aHO1M6SwR4ZDbIZu90mEulx4o5B/5oAjHGUICQb/cF
f4Xy8cCFB0o39XNzGhOgbavlcOxNWk0kJPCnJTSd+odEl7k3IYxOyo/vZiYaE4cm
kwtDJDg+qBkrSvFW1iY4BTzju9PkOwVhjiwW5NwIhE9oFVZcD+2GSs/Rg4L3Mk6R
ouASh5ZclMEABphQZ1aap5JRMl/BzRgXV6zAhV1H6PW3DsAG0N3R/ougxYoUguTU
eRifYLE3HjkQb8ULDFcCATinSHPAGdQE+ypW06TGdAxX4omSZ/up8jzl7Q0S0S7F
Xd0u/BN5rXoNuq0nJp5wfh9+nMzwTYIpoFXXj4x5ueruDHksBwmMRtlMG6Cdu9ad
w+mNA9FfnP5ovmjfwPL6Yic1fulfXutmbKcrqda/P0H0oo2/pKtDZFnwPnnGFAIW
JpJEQ+51v/7rlnIU2diYCe2i0Wq6vrRnWTZNxTbQBvzKgxyRCiZH5yHkCa3TE6Wl
UWHwBu9VrqrUwjiPv3uTZ25qk8lBY8FOf72Zx4gpUlYQ/OAyvcDM/tProJDL6Jst
qk54yMMzvS3pInXMOBkHiHDwzFpQ7UOu/bm9t/iTgPI2XT3KZjQx8q4feuquWIvL
YjWZp5BN55ToD54gqS/UtQZx/+jc993JqB/wi6vOr2a2yWIf7eLUy537SgpcDAfs
LirNe+M7RQ/UI/sJ+70fAvfqjA09gjop8agmp2rx7W7Y7+AT0QCFdAhxblqQnUY4
WVzGTeG0jZ1gxuevuysnG7T1Uo9rIfnLifSDau0rvRZ0Pv8IeFvLe4WTnKlXr006
hxfFsfKbEJ6WVgJPQfDOI/Z/JH5b8kLyymLd3wcC6loMPGOZBNi6FSnvkZV//d5D
bfs4W3KB9BCzo/eIKQdEGSnHBH4/ubEvt/77QwQ2Km51sKGYMsBGY9A0HqhWjJbX
cx32s3CWnDSHC5I66aYrGzwGs4Icl0ROlZSRkhzPbojanceVz8pXCGsyB345E8gZ
k8rbjdNee8sb0kw+/hRd+II7vW8KWQyc78FuvH14uQy0Rrc5PSyJ4toTfyIdTlrt
TNay4c16CO8PuNkDqrThihf4zUYRRYUGeoW5gV1jX5kd94SPAEbHSVLj3HHJ3FWB
Q7esFv0NCASlrpsEMGSnT0ezu8WllAuTB3+ufqZAVIek2q0OL0nAdTgT3Ik7CtAO
DBZTKvklg8V6gFuCflSt7rtvTHnS4iE2dpwbikCHdvWLJcM4QzI1/q63vIgl5h0Q
/aeJ0VqRtHU2DJSzIji6EL+msbw3/maVqMq6jOqOZc3EPwZ2Vw8EKB38MrReSkWp
9kbh3tRUZm83qwmixdgFwbBdVLcEo4CTGuKAmVwkVedg0TvT9mLGSc7zODhUpdyH
z2h989FT0JhoPWN9SMssJobCvb/y7PtMds+gfr/X0qtydzHlIOrVxLdJ4Ebmr+Ge
QeP9hXb+TBBQaRYUY2Raq38rmF1ht+Sdk1zyyaq442iJ7XcD0Xx1hX3C2z7FSAVO
IEONGxCVzKy8b14oxhx5809DR8s8NTxqYaKekXJuP70MQMekmo1s/VC36jjzeplZ
N3zB57gwDoykdf66Mu1/mB9zDAsUkVhNmNAPgkUsrsy+Zd1bLaf+RCb/sdz6Ew/s
fFUSklyuiTVOX/g7HyJPr4gEUUrImsSiyx9gjPRBK7pvxgpVcnSjZCU0TZWqEQAR
hLNyln1xEsiYysE6V2bGhP5ak0SNJardXsZjqXAUNOami1NU00pfVYdaiELLc/AH
MRhcguewxU380iMgBdRlfglvK2+FKhUC2LvbrLXMSSyE7sGsF0OVgz82e+/7D5Nd
XeGNIkDRlQ+i7tMvtr/PLGOvHu0J3fGgv5U6OnzjqrBQOoI0BLDVIqF80+kDnpPb
SaGqsMvwIBsy5OJLn6Rf6aS96i7UNWmEathFjK/IK7naiKFULqgjb+u9EbdWbrzR
Wy222gF43qXbItZoLMroup9QjbO31VRtEbV09l2+DXc/TN+MvD0i858w2vLeg0x3
PEtraMqllhBuoDjLbb/KtmtuLCXW6/vEZsLrg6otzEeUFRV9zSjM0Itcv3SpS8R7
uVOaHdOUImE8Y0hrZ6aVYwVrbSmQDZ5HuuVpSYeVLuTKWIwbNXt02olph+8Bw/h7
YYImpvf9SmTMh+yhfcNcr5KOkeP7kTAapRW6cPLJjIwLoSCfCM6pgo5JRSUiyRTQ
f3ljTSLpXg1clC6fgn8YPrwMjx71Bqlbe0SRuMyT01yB493b9i2wfxVyMTtXoXjp
v27fdXWeBaFMmI7YohprvUynfa4APgHtM8YQDChrrLR3cp+6gpHym3yMtAhyEMo6
Z/MGUNC7UyDETQiVEBWGqVktgYRpy2ZEm2fyYiAGQkJqvNLtHEYFNRBbpKqWHXis
GJa0m07+niRfuT7PoWGb6AJijbCuZyaHwGKbFUkmGOTxesmMnfpwzNu9eaA9tsK9
2i2xTPgEL+qA6uty+gBSSivfUF/QEem1/auIem/NLWdG4Sik7poRl1x7LibOLiu3
Lx9SuMRCp6ConfYztRtQ1q5hHnblNRjXRU4tLcV0TbNAjQTJc1EK9/h0ZoSdZPCd
ZX0RbDGPeCZ+ip9iEGUFkb7Fqy4P5HJ5VyIyAAh6reI8ltrEH87fNsKsGV9+AbgM
lhd/F3D5nxBRelKA+x8upzp4qVvvuGHV6bd6UXjHoEeA/ln4lPIy7AYNtmxn0OyZ
Mj7X1alqqtp0goFxDj4sWU6JDf2GxUc7NQEMBgUEktJQUywfWRTvSCAlPHzItjtl
pTkVCpHxju+yM1+jobAoCi83iqLCJahjM8ud7mUCnxib6Xjlng0KDUXFQDkYCehl
8fW3lsXsegF1RC5Ai7egp9tnOfJCDnZQu+rRpYqmdV4+JHp96Rsno6NKuVqTGYg+
D5LG6fpBrX+JzkyeXAi9oaJVyu8Bix3dycAPtloneDGtcAieDM8qCYqiZ6UmEyxC
68ES4nAQbhjJ1mRNgtx/gehXhsUKLRwM6CF90iUKXhSzSfm5Nr3luDK2e08xYxuO
FYW/AT4DeqBwmUP43J55LJjasBuiodV8AKWFl4qM962oF0d31t79plmg/RRhT1ZY
y4mMscNkPSWo5QS7Vphqw055/Xk4KQjrS+6rwgjoVkB5bpbZcINqMQporaCl+gms
zgxW3NA4kvMHQYfs0GKELauhL6/vinCur4wlBzDVzJv22zpo9LRat3SrFFYufN6U
oNM5MH2Wn7d3Aa0Pbu579hK0DP9YlX78J2h58vzTWt7t9abdiR8WGTJU3Wom4mSQ
WuP9CB7aRZ1kAjFNQQZ86gKHjpYkh/YlPeyTDkaKK18mFIWPUhXkQf4xzVc5mnJT
XbY4YwKL+FiGQGHbnWNIjx2R/8Wv41qxwsDeW4JjtDzYwrBy+6wt2Oivsn69Qgh6
2Bvl9UTkkbiAbJM86RRG65ComvMviPa1jSO2K3vCWVwhbpvGn99mH+A5geRxTs0X
kt0GOfPmTxIQ7q+jTJ5QgLE0a7UQjFfIvWPXLQaQ4rUB5+B5N9ViCOqAxuwJdf0f
sHeqRHih0VD/8mdMJZxl33qrB4YfbWPo5rHV719CiWzygbwKGrM9D7FAp3scQ/ts
jmuFfJWLWTYUlkJdHQ6onsJ7los+YSztJFG5bdhudy39PtIU1ImYHFl36e49oH9n
Yv657cB88c5QecmdjxxSom5YX6xxtwxPjdeZz+pkG0YbjflgwfOUCTGcTpThX/aV
N+xpwucZ0ZKPcWlBX0jo5o1WoHJuishwUlbIzJvr5q5GhxicZeXpE6kY2FyXAdqm
Zp1pK2soC4PYZobpfp90mgH+g3BvUJh2Oojk17W6nPJuQrJm2uAOxsHIQA80dQ1l
U0gEzPDC/3/kCP5bT1nTg+/xxihRCWQpE5occPAK7MvS5/v5lfmGNFJ11a1WHxEw
ddPoJgoVoAw7FJCavHzD0pbmTaHCgz+1e56jt/t+QlybhiRVgno8W8Rko975HE/w
aalVBBJoE0JkBgaYErgRxhD5oSVYct1NoY+dYllcnrIos6X3NlQ4ukcq9vvb9KWx
sOAsv9dsWwp8RjriDD918+UP2x1FqaUj8P29KTm6x1McqFFyBhyoxzB64xR8Lswl
EdzilmROwMi66iR7MZGkYvqD4cE/xIaDhXf9+WqCj7NE4MDDSLbujWqxoXUUy7wF
dxYct4Sh4M2646gix6/qboQYs6pTJqorGgHcM/WUDNUk83PJuVq+dq+s2ZpyKXfy
Q7ZKjS3MOy2nOfd/0jo90y0jHuk63kRJOCY2KvU3qmtNCcK6zlgRU7YgY0j+jNEM
sgmZS8YTCEjRyyFQdRwmCjvFSaWI7tWvJZbXBTUAvo5ROKrzByV7KS3zjq2t9J0S
DSHIQXB1mkF2D1k9K3iLZh79DbfRhR1FooO1yoMPSdMrYmut3FcJgUERjmbouWKP
GonLmZARbk46i1pca+v3JyOptXQgOeDk83B1qjv8N38AQwHjfyCStw/BiaISsg7Z
oHBTv7ThPwOkoBtMKBMmNmceUzu6B5B3ltTndu/vnP/zXW1KKQ8PWSB6+145Z4o8
o2nhNQM2kRkmUMbJQOmyyH7g5XNgoN9rJzDNJ6EeAYEO3ZWETQBLa3WUHEEIR/7N
6ZPNypu9OsF5kTGisNa5IJEDuZdOWX2NuxWfF2HSMTpn0nXpQXWXRVbxZU6j3ThN
cB8fH0+M7a9d8TE6vDo372Aby6CW4ye9Iql+weM/QhH1sme9ARzjiicvzUe21x3f
C/i4ve1ljWuKRzjI/I5feKNDQnfJCLgOqseKpcx0bwNEse01d6c1Uskvs9iv2rP+
zfmiOHNc8skZtV6SRWQ8NKiGHFKWN3UOQ5Qu4J5WWXIHz72To/MWn2buWNgFX+Ds
IgRuXFH3coZGlk9RsNdptvgtT/8VgG2Hvr1S18NH0q/7aUmZ2Ev4CepJ1ZAqrFJ4
5LBm8JhKfhA5liTPhnVH6ww01jDCvkWIbWIXaC9DAkI7cvjsz+uRMNQttW0H24Hk
1Iql5n8g1+QDVsWd68tlOZcPwTgbTO5ksPn17UgopQv8DLh1ne5bM/H0Txu3rFzv
WSawryKTTsCW2hdIMzEDxNc6HGgrptqBSCUTKImdCuuANn+WVwPOBLCJT+EtQqX6
enRUNtEPnnyVZabQ9h+Xy10Gz/SjxsuKYYKIEeIjWK7Sorhl3Xscr8sEtx6qvATG
YLVfdOQeUxlCAA3zz4Zrx2caMz3M9lFiWwArpLSffRssG3Dc4Fzq9QA5pUShFsk5
sBnqZNtKuFE0Qn0CFdwTkBjcSmoyv2xRfKwDFqgaW+1Djcq5j+S0fEIwzU46KwM2
fRB1qVSE0XgQpboAMvQ42wG0158eqf9psqWn1vO/3ByHAQLv7alnP8iFq67hWq7t
Eotg/27KVCXVjtEcc/Y7mZoGxk2DxaSw8rbZ7RKozapQ0MkFEwkyGsFytjFcC7T5
6SIim/fsQXPGUUqoz+xlPNbwUjd1ChKrU0hXsyXHhifUf4CwRGl1InfzoLA1vZjz
JHPG0kXVP7A7sPIdQ0KWOfWu91Kib47bOnIGC3UmOiJau3MESBnITeZuDKv1L4JX
E9yytTOnBxJOXxEOILVdYxC7J5bvXTFP2DRaWOG1qUwyC6E7Bu2Niy64Dg0KVaSH
OvjbhiuByCoIGO/AmQ9o8rWi/H6Ndox+51tdKHbw3TLAJCIcK9MwXXmbJor+9GkB
MOcmj/ev0anNy3PbdTv80WiF+Lf/2VqBFdnaIMpBx+8ZBEVpxzwZ2IPIWxhKyffR
0kWtoRIHiHsuyZ+sfpO7t52uyVcK+xhldCFymi8sfKe1kPT79goMG8iYjp3/n4d6
IUzB+I9Jq2lhEx/7HHdmpgjblIyEm3jtYgPXXCgkYPaUK8TjXGuH+D29pTSmQXdO
fqM3huex2lBiL9bYtIKMFIidiBpm1YgxBpN0pIJWNA87Bw+vmDmT08JlTrtWbTqw
1iwYda+O6jda4DNWGQkM+MZhCgBYh6l09+cuqG/GzR7n8tTGDy159bGg9XJUhtKh
+brZcKBZvko3s0XfWtJQNhdNnf/Y/iZDiwB9n69+U59atCxlYvYBk7tkdSe3CbVh
zfN6J12x/ugAmkrE4hYNUq6rd8sey0vjDcpgunPE+LhAxpJEdP4NYvLOjjCrjg7M
vMjzrw7CPB6RoWBnbwMxm4wDfZecl9bZvx38gkNATECOVY2GClOZ1OBae6xYgUmu
1pZaV+w3EuUPtc6e3LdXrNuqxmcdTNFBFM8G/afHAD4LCSwVfxkKqa1dzDQtXGEJ
Jo+oGV6AGZnZHG1QULSGhtYmU5G7+V4XC5kPZ/xP8KCPR5qErBOvLSRMb45FlBtC
Is7I0j5h009y/MdJapmQqVQZy25pLOojSsSriL217jz3oUb8J2Qd60Mvlp+VFsQY
FdX8TJxHjb2K6dxdIvpUP7jdmTiZAtv9nY9vTuwsYbDveuDfqwHoABNs3bw73V4D
73w0hHz3SAGPeqceiLg/qODU5nv82zU1Li+nG4dYBkSOJUCMgRg+vfa3CTFHGAyv
s/Pfe02aPuhqCe28Ph2gM0OCpPqfkKvtTtV0ljftdZ3RiNLPj9dmTbCfdyGS9xRn
G2iTMdWqfflC3iyf4GsSf9S2GolNZMhDcLh8d6YZLHmmZv9JimsYsWHYBy2zSKn2
FiogqKeukHeGyw1cLL582PNQ4Yr4U/o1K7EdDjuuDZLLv1x0mvN3Xqyoi6ttgokP
swhStERbq3yAs6ObNuh/I1uptVI5puqNWW5Aow5mNgs+9XYfSMFIrA/F6GZFhnPR
KvWzQWCIC72RcZsG4y/c5nGwJBZDjlwK2sczIT6391ANz005g//aAjN3InoBaEcY
jlh6/5kcYRZm8bMzT/FqH1vIs7kUwJzg6PHVl4f5rVQaLVR9YXOX0Wh2so9DiHie
9mGFitfACEHUktGTyvafos5HxESLUMYE57YUhkvNtpRamFlxfE3QUncSy6Qz7ouN
a6V7mao2c24YA23wtPGg2QBSuhrOfaARPQ7A2RJsDdc1NyBR2Nmd5VKCZtO0dd5W
6pZe/XgbffwKciV7GMaXj+FS9v53zUfqKI0HIY+TGsObJHEGPyfnV1sA81BX5iBK
7iO7P/ICxcrVEZ13M4Odb3fc0GgO91fStctKb6zS+zNf+IxDDzG5hTInOJiRyHGP
DmvoR4PC2QHjLgzozjKXjFKtzi5mfdl2PMI51rYupDW4GQwqCTMwYlYO7KecouBd
8n0kNK4dHAnKfsqkscFspYcldTgSGcK/pLgNkl/srLWo59V2ugt8iDbouAKCBGyX
fYx6OWLh6viJQWB6b8vaAXDYE5mnXYWEkzKQz2RnN/HsNqmerXVMsi8tl11+iA5R
wbTRBpaCzh/kN0fOccs7KUceNV+//OEYj31bQC8LF+SA1Nzmxy4FABHydHsq5MKr
PK55UkRNtzVqDq3jvbuS4EkzPSTKHOs8FdLOLMA4FkbDJ0XDHdR91Mi9csI9FF73
GbMbC8BjlTKicSpbBzxjONjR0yxkAK9ixKyoGECGVunFPI1C7DqUNroU6dvh2U01
aJCrGIqX8ydsytg4mOxxgl+ave7ZVBRFwh6biL5WJQ3b1zBsqwErroqqMMxBsnyt
Yw2sRvMPqEjJW4ptY6TOsVRP3aEhUyOzT/HYndzhdLtEKvg/nomvZcEbYi2uVBac
ksd3NjlFko0rS7sX2ljcCm/AzSf0PdjCZ7bZ7zpR4be9oGbhJIU2TkSE3nlLJSEy
6huQG4AX8ggLaDnG9R7MMrJ0FGZyEbgQ1ZrOYn6acgkq0fd8i1sO5a/s37QIZWOX
t5mbciTt/rw2yAWvi/eYBsF2gg4dM/u9OMOAx/3Toog6XpTj7wsjjJPDts8KR7+y
GPcNcXfsWo8H0rJBmaPWV6Kw2AGdB9TlKwmAXAbjRg71UYAoBYi+/iqI6XqSpXvn
IP8Y+sJcD/BRXx7RXf/+ReUoLeEHiX8vHlnYP0qK4MCOTw1IR1+uTXtAXjo/ho2I
GPdDUNH5B0tYw+TuEEdtdEuzXtgpYWpHvJUgoriLMEEojSkfMzCXPGppfVMJpxFI
VIvMv/SsT0pvkDW9+b9AM/VypATYUCY9R0D/0qgVIDVVdsQC96ytgq1UBYIe0pVx
ZIfukAttcuOnKooQnaG2XtIrWHW5H5JuEG3ghjXO/+PM9g0VUaPwm8/dDHPhegtK
nwkbktLgeYrLvDDPhNlQDOxZoiiihGZOJtay+4XM3emuOGIIaMyiaWrKXgkmspLZ
RTxayAv8ssS0KpPMldGGqX9/Nlw52fpBS6HkJfam0s/GmDSs97M4Ks0oyExLAOUK
j13oRCsRZKVLsSWhSQsHWMtJ42XRmz9O6soruBKZZX0R9j17SGoE5Cg36Dk7s3HN
c01C2g+tY/6UXRgp5dO2vTf0bd2B8dGkKny8rw0mJj2OgtHWY8xCtzgeHGQ2GeNT
gOBvQAKNXwrrfLivqyucpQETzkH8RQsVo4+1IKbzYEGN0drSt9e1aYvoZNR6Mn1t
Na0nSaAlPFls3QjUjLODujkSoM+pGgC48PqceUA3UwF6Owz22uoQ0xhhQ+uERlW9
p9yrkiPLCcsDJRwpERbOjF8Ul2gwgRvK/ssLvRu/sTuzKTlUvCVQ3sgAACzPtY3g
RLO0eUFhAWcswan1v+e1QGDbLZ8Z9WATBR3Qiw9cqqPC6PVfR9Dr6Ld59NmUqIPy
8Dr21CacfzYrs64j+W15mav4AnfqtPGWMC6OL0LobRqUP6b+3o9xXvWRkrNOWv6B
NX6gGLmm5Sp1efLsJJlOVCzD+hewhzFRrxzN6CdXZESMOe93bs4lPDyo967gp5hi
TMSwAjT4J9aIoxAVeF1v2E51nAg6Rff15nC8zAvvVKcnO07zQa9WJg5LC8FJBOUb
Wq3GJFnO7sFBjAngE2QHqw+kNyLFiQZUPSJu/JUTUKKUpr/Jvk15qGg9QJdMy8uY
PtLgsgK1zVZz4HdKvXc/pyS8Wn/fsXPuNK1xUw4ESrw/AKlq2xbH2AWy/XkTgBzN
59TmA0mY8kFt9Vc4CkOiNVpvd/NlLiZQXJcR3z5+IIFNN9n+ogEjOxUukHEK7cQC
gxZy61ta83GCXN3NE+7IC5Yc2KTPadnRXdjQcbwAgsTLNlo6H0Mzhb0LA5yulsm9
bR4mmfIVnlDs8YEDP3gYJcqBRYUiCGLqH8rNodM4bJ+YekTRmVf+MctuIUtMkx/7
3ynxja+chBt8CmOxSnee8WPQ81ujMMDNTRq1kgNKyeQ0rrUQ7DuKEyox0BnVRZH9
wwI8/QTugyPiEz7SVDuLqAaOR7RdCQ70Zr3cbgAjt0eXMqFba9G5Hhh8Vjc7zVmj
phQLt7DOvZTvr3ajz8I96zv1q/7U0RSOLLm5N3JuY+MpptPiJInxs16ZVACGHIUl
pQClqGXhmlPmXMafOQaDdLCsjl8xLmh3v5D3fxYSkJinXx7Fjlm9ijteketpuga4
wHlpyuN+Sa8y30mwc6T3c9bqu+VIYzrY4wGczgyHZkKN7CUu3EM1wHz7WaqL9us/
b+o/EZZkhcRS8NyuHv4KxS6R8mgUenlEBbP0JawSra2qu0pvE5SOXDIlKlOcTCjM
9v1i7yfVL28nRq1KHa4Ye7Bla2dA3oZ7sIseV6CicZCgV9vndkmQZWmKE5xoAI/w
0aHHSbQ1rkFQ/RE6RTC3UO5sbDrAo9bpIffOtkDduuCMgEynBtGO/oIKaKsvYFFP
wEC8RmIh1RmxC4gTLtfSsA2PtZCwUgWcf/8BBr4VfKBOTv8bqH//4Bo83Pa90l41
z79nSxfNg95M/iIQz9c1jWXI3idD3qQduJM8vST4Fq/uoPsKDHnq8HL+qSLsD+te
V2SjTdjJoxBNkoojkDQGNQHN3h1GFEUDm8BZfO6i5td1NiKWqIqoPNFeivJv6iEh
M2BD02th/ZqA3PXrzLuWRS2YiBQpV0nOl+mImxTD6u4ZH7S9dvsQrzLWz1qpcfic
FsScg9UwILRdMlTE/YSil9MX5UZnS7SlHGckxD/HVbOipf0zG3OA+3nNE2U+bjOg
iiHJwRwuFhIsLfdWHFfLIFjSzdlix+KoSPPuXuioT28V1UUQwEPQp2YrdWE741n/
z/hTtHdlbP7kE14sfhJnDFDhwmf+jgRM5hZNfHhcR4UP7xv0nVQmE2CX4lIZQH4V
R+ueexm10ZRHGxLSIIGAkxbRJOk6BcjF8FifrOtDgFLUkjMUkIA/584HNEOSHiZz
kEmHohwdYWQzqPnNdqOfKyvLjPNvAvQCTtk/SYhQNeTYYl/MKdaVyfoD8baAlXHh
Siht6w49UteGBg03an5NNmJ2JK2tR2n+TiEhvK5YEA38ojoBF3FBXkoY+S4RN/Y8
0IZWqaITYnJWz8mxI2kUDDsXnQM/HKX/gxLP41SSgshz9OLodyIiJHNWk7UDyWff
eYoy2+P9q1B11AjkMhGiaXidLogW0B0o/16eXOtQXw5wYgzZQG5ak6Q3iLlgkFHA
HUgYkUay4cqtKy5hikV69OD+N+QTPgmDLgH/gCg2yQCyYiJ0Nq6GcyllWkaiAj3Z
4ZQ7Rk9safucmr7ip0RtbKlP0RNRusD3lJfofxt1upg678NqEuD7vRk2K3+gFvEe
x+H7CL1HGtXVegZ29uQBvqZYXIeZxBu/rLaA+3Xd7BOI9y5/0pG+fYQDNJRs0hOg
k0pVbOdvYjG6tRl/7Ck8LOLTMCbfOa/6yu4uxIDFo7oAqAEAlTlTcIjRDEZ9sTy0
3D0at9TUDBLmDlcQ7guU9vJ4SE5L3lo5IdYPjUXr7VEadnAApiHlEJKSdNxUC2Do
xultBenv6E4z1DI7X/9sh1fxe7DswfGb3hmCOTNgTgtjh04/vRFXrkZ2EcmFHQ77
Ybj9THaEaVx4E32PqldkOI/V8z7tXZMSk0N5ft7gwTdd8WSiAoOYkXTEgXsLq5BI
e2KdwCoUwCGId6Y7McIfo1t4RMp+YOSYBPbG7NXXhk8jBXCaLC0iBw2IGTU9+nGz
jBUnCFs53z/JcGOzv1hJ3vmYha35zmBzNWH8rzTvsWSEMkzrd781cHi9Tai8/pI7
yUna0LiQfBQwWxmbBlf+81xyIlUiI6JL4TOewnE5AJIjEEWQQVSq5f/5OMsQrbQO
YL7HHnvf5FId2ySnWzfS0SSOBCpw3m51BH9Q2gb5Wg9yrTBI0zEZ6d+AApNOyP4P
k5e6H2NbfK231/Cn39iOcs+ExInsrDDN13WN21whd4eJq3n0Z62pk1b8Wxq9EKSe
SWJ53DgICXX25scUOikdLdIB4VjTfnwqu5Rx2ZIv1fo4UD6pADYIXIgb9lU7BPa4
M9MoQVCPqUzB0NkUm4xOELtfdFYeaEVvzY8LAIZ0A7ejsvfW9EQXmOm9DxX4Vf2e
4DPwxNAPFsMuVJGdxRzzTb3G4eGFlbxYnQ10ZAIEcvsFkT1pIQz2lQ8p9JT7cyIH
C5COwGrvO+JlRoUPpaDX++qFqv/3xWhpNRhzqa5197MyGo+PhGWVslEn8LnM+YxN
HrGznj8iUN/6wA/AtY+WC74D+snYQhC+Y6bhi/PZC5ly8LZXNIkm9vHdFj2A51V1
clsL5IIVvmR5lTjzyWFxGGfgaanPyu73i+nF6bcpyCTpmgI8btY6xSx7ho0O6h64
cv1Pzb37dtmC6BauOhYe+PLZ/fZ1J1bY1R7Q8D/yny4aS85CwqssStRysFlXdu4V
Q58F+2B4fIE8NeiEjXInebtr5zfwCEaOCRbwcQRIDgKcE/WTAf/zM3+CguHpqI1X
zrsMFATNg9ddLCvMkzmP1OX6w9NvNnIIbZY+ie7fsH6bOg1Oc6/XiHtJjqLfXjPL
V0q5WKl5FWwFJTjL57fN6/R7NtFkDQjNeUeABE60Rp68T8yg7YcUfYrxizv7YIzf
U6PWCSRXKhHIO0lJJh59qVzkl3mgdjfey8Qm+ZeO99g1qEmIBynhQh9S/2Wb8nPB
C0qU5JiwfY8nhWj51bonctE35wzfy4EQfhSJ5IPoPU2ZbSfmULO809l9XXagw2QX
u7SnOUi3ndlwJ9TjQhiLpCKozZ3nntITXlMn/bjlmmNeFBIY33xLG9E5l9OOfS0C
2QfsHjYJGtfkuu76VWt/02p11mXvgYJqiluQ1F4lb9Qj6JyJ63SibqVtSckht40B
mEoB3yCV1ot6ar9FtPJAvVXO3FKPqDQ1OME55vP4FSL17AgmXdHR2q+5AF++N4OR
lnLlqkgDZ5VzHV7SZIaBZ+9hIPQSoDOm97vPMA6AFJEL2/qWD/h8D6XhPeB1DR3v
xwsbI1Isy+elyLu0CEedGV0mNLeiml9R+NbEQnOipfflgRABqcA8SoUhfdd6PF0C
ZuZ5EXpXKNMxI9S8PEBENMwbIDr7bJ02fE1ATVm/ftfz1oL+WT5H+mK+QgEmagc3
9JDPoNCjF8ObMZ9l9suOdlo/bd/a1f2M6QreS3wu4cb9/9HBQXY9eCqfJJLKnvWG
G7Q5trwquPyxH5LnltnY3W/+NQhDj5SiyWzSXhXUoOYcU8xXl3irzq/JbuRV7uNW
XIPSDHQ8LfYgOploWeBITjizVQV6gkCin6r3ACQSTR2htC5n0OBJsx5lDRgq9GhK
cwnqko10BlSdvYP5PqxuI2r/wfL4A/QukDIFmpofTqIpHDOkAtoRp+1nvAGlo7c5
pyuQXIGy3Tn6OcOn9QWSsgivEwCa2vz+qYQO2/VsMtYWpgd5bfTQVNWqOSN7liGM
fo/S+8KPrlgVH3S6Of/2Sw7fcKUjd8drKkKwnOMVufiLR73LuyviztfvWmwAq6Ql
DIqPsnuJqTTtEJ79Mq0yAynB2gACM/eTmxGEjhVAAYrr45VjW6Kmb30PMfPzRfqb
RDa+nfQk6+aRI5AuDW49NJQCPQVN5a/SLgKxLva++7F6m7tYk/VdKX8lZ96K+Vzk
+oLuJC/uiXSIveIBg7d1jRvSdE4lds9BT9XQihZdLSs1/JgSqRM7o2DYTQRGD2Ch
LVfKh+z8hLUbv3k96YGiCxk3BOhd+lQI/zTxtBey0LKa9Gc66q1ar3P5ck1islnQ
mX91REWfNr0OcoEDDrViuy6GXIdQ6V9Y8TgowOOVWy1C+ZowkWf2PI/p3PZA3k7z
sf7nqUnpdIHoFgTGnMrZ+HHCuY303kYOt3I0U2zketU5MtvSsJNLd2OcRlpe8qI2
m00XsarDv5amQnyHbsz7y74cRZCNzK4rYXHHEncZTyjbCh85Rgf01G4tzPiIj8MR
KCBQZ8gAkaxgW+rQAKE71RY9EnZB/4YecrwORWMWCHk7oSzb8hm8eNg8XVR/raCp
8/5vSmMoTPyaa1Ip3Wyw7xEjztDE6m82Mxaee1eGrOLr9PByriZZYPwZ+uruAc99
GSCfad7xVDDqM8HnaonNN+eGn4fA/LatOuIb2mw2vZAp9qY8zXwg4Cf01pdbJN31
FAKCxKuxtc5IeHOdeFquXxGWYaZK/Lef1R2qS1lDEuUblIgewb6ZNkLDDNuVx5T9
YPXAAVRBfiEAKAd6Zaie0LNJ/QU5ZG2iaeB7wvCHHjoEb7RY0vK+qJUNj5hKjPVu
s00WCMdm20MJbcV3E9sjylNo5BsJFkj8E2lPijnusYVDWQN6crCbH4P3NRbGJ0Cb
DaVy4oT0DdogyB63+fzLo0Ss0ELhMNK5WkU3NhUubK7FcLMdnJ6SsGfgCYWbaWFC
pzkRpMzlITqSGyFGbzIymilJHcu9wFdzGUa5kqGMeAMT8sopX9eWE48Ax35hInLe
5KY6h9AzE4QJBtNANz1hZ6uxREHEUUPl5NiV1F/4Df7eCjD6ZipzUEMBCJMF3vGV
/9iuOibMp6Zn4w3+1w7OwfvlS4qPTOrk1ceFdJez3jiBdRd7eSrbWAc+TjqAq5na
0iI0c8qZMiO61DYbJI/wcNxRdgN+4NDT7v2UJisWYUJyfuQbYOQ4CNazSrBhEQzW
ha1I2bZEM92aik7sjz8Sth70cou0Z4dnKsS9SloITNQK8jev9OtL6JJedl4l2J3F
NVXNaPRIniBbMHlWHpqPTDH78FlkkRi5No31Olel0UpZhiA3ky9nauow2n5dz78a
mRXfDh+uKj5TD9JhNzNH3d+QJ1yOGSu4frHAV8Djyq0DjrRCTOGqqImieukZfbDL
LKjxzRyJlTg1fJYUxDo53A2fVKvrV6nnWGVAh8Z7hYOuHem3Zif59AveCTJqpS30
vdIyiYLbTQKIPHRAxlNpc86tG1jaUeQolW6cCMVVZTcLFSYTfFfADREanVjm+IsY
k6N/s7HnNNpmMD1Mk5gFX90jZ3WbONcY6kVf4gX/9PYYopoC8ntUHANWxybp2sy7
KuGiVfluLutQ/d/5CQ9I1c2pAbUvR7D02GnBmiBRE76fJ1w7yubAjvg3oOfkNAIc
vnGhZ7CrYGzTB0vc+mvWmEs3Z5O5chliW6pxVP1sbQBWUISzV3o47K9v78fZQqWM
h2aBgZIwb79BWkgWNa1OTKZk5tBmQ/zrjcr9YmlsR1vd6xvDODOHlqAs0lMpK/de
+dHMCEPMY7nU669BNo9BULHR/U5YSsNdO+JrpRaV+APdgb8AQ5D/TkNEZ9Be11sv
d/Fw83CIMyw/3Pdgjk7mNXuWbCczSI0spoixTgiMRQnTm3twdwUD52VN/+O8gYVD
nrXhR5EdSFuxQOOcQtXxrObSxeWzC4yKZUdlE5z2ZGHrOACCsybwYmgwkLWgzZSq
xPo3/QKWbHHHiRUwcFgXRMhNFtK5GQQBTlPaFrnRhybu7rfiejbv2MmdjYx+XuzF
oN1/+Xj/8sGRvi8E87NzrtY1bSJA8AaY+kGiOu+kSukzMohWQembx52IiBUxbkuU
Vbx7bYhFjImQ6+X5LPsV1qVCbyJ+6i5L+mUwauIzeFtf2Ehbv8b8omHc/Qjppn7t
RdqjBTVScTS2KqxwecwuSk+dbv4h9++d+6u2Lm8bBZCqiwEkvvhMhhoam2gbCv56
1IoVJlrEtSSvmhzNokksihnQGUaxOIv5o5o1F/GictVhu2S9YlXBNG3GYN7yiv7+
umXkQT5FaMAVTtiW461iUJdR8b0+bw0g6u5F5V9w9m5wOnKOQS6jUXKVFOZFSVNx
5CUaUxI0sW4xWPw5N5vcFs/9i0sRJplK1T7JTDqFQmNvyNFloUwWl638hNljfdPu
pE+t1SYwalLCjVJtm1ScRm0mTaE6Hi2i91yNn4mzX7n5XNODob3TDFh6DINoRH+9
IQa4+PMoykMI8kxk7Pqnrfe0AiSsWzgji2oz8qQerVzd6kn7ekM8LC6WTyFH4QK5
lAyWk6jvQwfIryaIxZaoTjupXzyEyttfmYBPtey/09apWhxLiMRU7DcrSvOh1HHI
0EMvZ1SGCAEAL5JNa5+d8X0aC/sF9n7QX59xjDlgwo9ILOxkvF4h8yIITwOD8otr
ypFC8s5iEunG4HjRCvwwE2qvheCiWGHm5oVfm6DQOk2kZUHR0uuQ8+7yqTzLH7eY
pwE1hunCt3tZfvt6OFTHs4B145QR91Mb6CdMIrpwodmlv7u4yEZVDMBSdRpN1CdW
0DzvvDsJmNwfuE5OSc+K/eBL7xIZnO3BYbvvyA/gT5gCZtAgZVIUwfE5Uv5Xpxk4
inbdW7/gOCiKwH35aeeJ9DxHkJQym2RovwQ07M2YLu1xdP0Xi3PcXPBIS4F85dEb
1izqMLHj1I/SJOyFjWn7hQJx38/A+Bc5JrfPowE+VTTUYlXaO7rNFK4AlW203wmP
oWwpKspRPgSQEenvkXSyBhYNZNg56KMJqJ8gH+9YeHbQkDjMoLvxOyS5/XSlHiBp
tPHOpjQR213vCkymsWevJenuCnu+2VZqYM/av4K8ly0vZHJfSs+JIhHQYXH99GKg
7eF/bwtp7Aq87vozbC6O9YgdP85ngbQuSQkZSnO8Zlm5eF3b4HGTyZPnyEgMaMJ5
p3R+Dcmr81wcWxe0YXNjBmq9oMQ16mxOMMNhTzG+5pehKxzcQWT83plC7zAWfVKN
fwJ8H2Pxn3U47ggDaEsEvJxJMKbmLL1TfcY0E4bZ3r3xw6T1krVNf0yeSgiiZrL6
lWgqY11sZa2rD3DMw9zu/aGofi6eaaji3SzyhmT5YSt7xF4FHDVsXdWG7HXPCYGE
MlA0wg9XAMVTuGZ65iMUzwv+HS7FxS8PbxqB/+1JkpgLaY9zIlatIQGKtaXRwAvc
3FXDsdPDMsKwDPBGRajtx9f8gQgnTdDSZpxRMA5ivtHIxc1PPt+e8SoKBztFxHBv
iEhuis31CClBvI9WOo4ZQOfUahtSpgEVBClsJJ59KYrg9fk7nC1L4FgjkNSG8EG0
Vo7ZkMsfr4XAYWnZ5h78xS4Bte8u/OAB/twAotU07ZnXmkxhhCJqQFRToru5TqY5
SqjsO3ph6qXVcQYO1WYyPd7VULNMkn4GYaEEZ4Pf0eIkXG8y6uuEprQaUXb9g0ag
+bYYvWepo+X5vYqq0eL4o1doR9MFK+deWSduBpKIzrjCkUOB+aXPhYdUV4zckjMy
avGKmd9k8bjJM9pKwoZqAQEpHonIG5VXeEInNtNYnhjgxwLCtaUKxK/0cE9GsX58
kQoJ0+x09wJt9fRXDOT1060erDy4bL4Mt9YYvVr4woF8L2ekYSoQJNpGpW9rzAqk
mInoqsFydieKvp/InM2ygGucb/HU/lPpFh5WI8uKHAJBqogQeyACoX6kSO5XW0k0
UVLdYYY6e/cNuTRcRSqyOJIvbBV+ybdkYKG5clTZD3ng+prsz52IBvDJenJYzqrI
hmy+gBFj46YsRreORBsyvx1CGby2BvDbGT019H+zEzyxzb1m8mFxNXe/59SC0Ass
wna/ZErKkV5aNlVIC/zmjRdAGlWdxhXgpLxaVM6u0A3GHX86xZ8VlCG6Hd9PuthV
wODVut19+XE50espW8ciVpI7Kf022nQspy0VCd1S/2v20OQsKWp/HHMnBldCapId
Vt3ZMQa05jN3n+iWfOVZ9iLKvWM64lbu2Io6CUHZfGQErO2JNCfEO6aydOWtoKxf
RO+p30aGwfjfKD8bd8PXYXbAEaysZdcrR/MF6xOaLXZBEEzZyWWYzZ/zsSDTUZ/g
kImNMKJtfC4Pq0+ZgaY1FrnhlbqMIySaI6Z85TX+fV5O++MA5IaqKj7YcHLpNBBR
vSciAb/GBFslDRbtdWppYVl/HH/pBcKWOkKX3sdK8TE575zJFoMMZ9CAQjkTZGzG
H7f+gLr2PHPshiVHaDipo/dbwi4efklJsp+8NHOiVUa+wr03aIotmjrXDA1oC8E+
5k9TJiBMLjHB8iuL/LQVcmEoV9J54o7QGK4shlCaBGEskuNAw7w2CUrWe89NgEzp
yjcd5kfHonFIDxhLxzpo1wR2T3rh18RgluYNU1gYWjRKv/G21k8dLUe6jRrtmxO0
iXaN95mJZXtjb1CjNyF3llVltA1kaYfvYoIZJ1eaF0n/CGoO4+yHklQnIEnulQeI
bnBjp29vr6wl0nHLxi8bUq8chMZTr33xVOIis/o5SH/a4DKQPTOz2CNv24XZZ+Tf
q76viFFGh/vHJEN8BdndjEZPQA8I9TmfMnzHaPhaYpadD3krAUA07PJsJjf0rOAD
xcOshVlVUtoB5ZqBe6EnxPVHFSxQm/sx9/6z86FFzNu6GySEVUUuctaXDBjEJkbS
vR9EYJSw29wn7fHqUT39zH5d+8XKs8LkE1Gy9WWgDzh391JiHRyeOv7iORI4dCJo
pzOWPdilkoRFkeGhAqsa45oGEHEfBwN3/PD15OkV/5kgTIjgSKGBH4cQyv0nEYpM
D7kUP9LvC0iSrWM6rUVDJgFVLacW9VSWKBinl1Gi18e613v2XQsxlCX0LsmbtNON
k8SpBxMfUoRsYX/NJQH5cHmIMnShOS4qp2ofbhux9V2TB3UIaVAw9FE7eYcLxhfc
KLfXfEVEFeex6i9SBSdMFwVH3zuISB7l/xM7Rjj2Td5TQRtaz3xHM4YdQOruJ1PY
m7QSKLtoHIo6lJDiWd17nW44l0j5Z32Ow4LgLbJBZvPjLxwoIHbysQBNH5vGuAyn
pCm0FTENUfBOW4ixwMv5TmR6fK9V2YdP84XLTShmHZgKYnV+n440RqUdS8doQGyJ
cEeajQJR2WwYWL7axHxl4Ky+Iy3fLAx+KGFpClLr5tOCFyCDd6BaAH+SEOXOR3tv
+7UL9lT0NM5Yi1aks/NjuuZOn+LaBlPinBsAd+3DVdZJX/3x2XzWdXyDFrYv34mJ
XzlzC/sF9RGm8dIMEWdcfF3fkRf/auYwjxSEOSJftvhkRhIc8OD/SDGBtLUCLvpN
Z5NOdG+Kc1+UwTAXf3BXkv52fkDnMbatWWfMhbwEQmLuket7G2W0gcG+Ipv24NQ+
NvEGCuX5SaYQjeboD8XgQ1B/8Y9AcqRaPjbTZ1+jBXUwzNkIZeMisqAKOkKh1pAc
W1aPYpFiwCmmfE90ZN0LQqoiaGdmZWg/o4YMc7AfYopuWkUGg25Y0MBAFKXIqR3f
6TmiAInbOlBzy/c566Fqc4setl46PKMfeBDjsenpa2xE07M1viPhzIjdthYkRtMH
8lV7VZzzueYndrYTQnD3nqvYU01SU53k9nh+ZaE26awzZ04FmXccNYE3Img2cnhj
cByoN3xWHqWCQhhQsrYoirb9AQS/WsbciufOteWrXZu2Yw3OeRC18W9gMwkCdU0Q
QQVBKPKSNevX1wAN5RakTuFrI5ugfH5E7ZdHUOAqTrDqO1gQnQTS37zz9KdY8fiL
RnC58jqRoEdR5cEdlUax8uzZu0Ov96ngy33naXFQ5DLMvv40kBkGhypaacFLeKtk
QajFqvA1PCX0IftM5Wp2/2uvWydQ6K/5ozkSuIyZ7pjQASBRj7qlXfKGuH2E+MVF
bnXRzZt0AFRAIhlWpMAMTHafO/EJc7+/NaQB8bp5FQH79GI02z4SQSjSh2XkO/ds
DgovSDTn6TsPd0sCDu0xfaNYSgpTj7aCk75wKkQY4qdcrHlkJqL5fRdLMgc5U/Ts
yxWiVPet8Z7q0w9g8Krj6XqDv3AXImaWuStjf/UyKX29DrTajHI3qnSsvSPAWi5S
hGa/Xha53x/8wcmq1ZMwtw2SI0pkfpe6Ea6cUrXQwOyz6hE08N66atZYXhgMf2O6
+eAlx/Rsl7HwwZqMciv7ut9JTTGyuc6zCYYaAjx2dv8yOXz1ScNy634X1S/dWadi
h1o/YIEAMn0lTa4Rm1VNxJ73LBfGRiQo9t0l+8OeUxCQ563ssm2QTqh63BQQHPHu
YI4/RClIIGsvajL3V8GAhg3AA3POu2wa9jqmHr7NzDtwAGB8McQdLK5Abs9buE0y
NJpABt54lNdem/DXXZ+paANUzE4rVjvxzboqpXeJPeaKBPUcT9SIaHrR941NZV3A
S+WMVEZ12bXLbRay2fEGlzzq16eRKcj1vUAhmMJ3nK4lClywA4O37K71qCmCsub3
boZF15rLz42NVTGvjzDGwyf/XIbHDBkE7I2SwB+xu5Bhad4kQWKjXWzkBQ6bQa/J
A61v34Jd7V/uW+02CUCq5jClC6u6mQ3qu3a9ZnOavbOadC2u7QUR143TkHbkS6Ul
ytPhzN37HvVCKxaw6xc06ImoqCBPvMJMeGJyCWSbKvSFJlK8uI1bLlp11XerYNYZ
COKc7n/jyPG0q+vjSP6hEc5UNALa3LDIGuY67FIffQ4ai9C6yzlpR28tJoBtbGqa
SyHI38GQxmrYllVfiiV7kbmb/Wow5JCBSKplnX61o+ZOKh7w4u7T/6LPF8NOaFKT
poRr2oD6wcdUxHMHSjqeF0YcPE3i+a+FEsU9Jl863YeX7pDjfa3XTPl7S/IpYU2W
NWcO9N2m8AKvFB8Ri8JvSej8zWrM6Su1tPerwKX4BcZJ57F9q8bdBbEsRc4TdeB7
khLZ+S+yR34W92mH+kZJpK8XefKqb7ytiR5htIlV7gpb/V1PTkyKS6bxf7jBLJwD
vMAD2C2/Pxh/ogMaDjgZgaBZQyCvO7WZWrZcyVu4WcB0W8YAPDTSPXagK1LvwbyI
g5HH23Z01lXY8aLOzcM5XllPzh/UoGq/NT42U85uYadmJhQurPd+B3dFRKzrKpZG
lFMEfNzPU6R4xNaYKD9kguu6QovqSt1LzV3woooyfTYm8i6PcowOmHrbL7cFoBun
RkTvm9EfF5N7tR55GCLmUNM5xY5Iw+Ce6DWpBxyACrnu6GGaZMMkIPq6QwIpa+VY
a6BJNDLeGVxaCRqEVbTUtzEESj6bCb/7t3tuj4ZuzIOTUszLTEp6fr3j+gFySBQy
mY+X+IMWFV4frpm9UOYEOdfC+HidlFkP98zqokQv4u0KGbDt+1M4fDd9zjKvwVaA
/9ktC5YumpI/irOgNiD/jZBr/61GyBR8b1uZdbh1T209IFotn+5BfKr8cUg/FPCm
hFYNNJV+YRuQJk3t6aB1vry/aY+BEdmsSwYFokLg+l4/IWBre/F/vuDxAnS6cPeL
AEzdd6mbbNpH/Mmecxvef3JjoKHfnuIoMJyI0h3Y6t0hGwnx8oOFBWIC2Lk+6I6b
umXgb3yN4gEWmY6SMyxFJtAEmqI32tvPbo6yr6ZlgLjtLXHBseMlTab8zXLFlIT8
wgiO2UndYIcqcfYFMKRGZNWqd15rXddQXVSEDyc74J0nlClqKRhuy5J1ur18DpUK
8MFKrg2aZ9emeuXnGP246JjLBrsOITPX6ZaDlHQLb+8Gdnh0qYP4xEVuIKWsG5+i
vXWLAMkuMYEoqhGKkRVzIfKuxdZ+FmetSZjQZfnJ0VNjrTSwB/35OHNmdObYfntz
lh3P8x9G39mmimq0QAvxEXn2xWQ9E0mlqQp4adTE32aDKGlhk11OAORTLmLb07qR
7UiLTVLmfYpWY3KqFpF2Md5nEeYuQIeuVKIaxUMmOjrGwdWUq68u4DO6hkyINLML
+0Sirz7FNYaeOWspA6ve4Pkvlz6UjF3ymL6GGIb9ysWD3KMP9CFy7NNUaLrH8CM6
c2LqLPltlhW9dC9jii813E7ItkPY4L2/awH0U3gJD5VHGUwlBi2M/2hOhC1xl5Ul
K3anI1OzOxHQ+YAkwAozxhCQ9c8/2XNO+cAVVemHL9OOMV5A3cYUpBqDtyLnPK4m
lo6rLzWT2Fj/lsB9EtgYYV8dgSdnabJF2XuH+Hxzx2DL1GwEUYOiu8jDFXLzQ0Ry
DuvaMRcQKKG2p9p1Ky/Qo+aeaspCnC0G5NfCcl8BIcQ+M8xFpKwU1kv39YTy6yGB
Gv/OsIvdhGiuijrY09lDcy2zAbJFsxzKt0qeL2dH7CvI0+pdSekA+GgN+o5tBuoo
n8lqdjIDf4nHyeW+OShpvg1ohpvydYW0iq2a22iSN2gda5z3hDGZAy32rRFDNVsq
3b03XI//nec0BoRfLVnHjK/uuozLogKFhbko1vUd80kf1bm/5EoekQ5gY84nssaD
qOpD2BCx7iUlh0CpH/vyNhlQCa5UynEV14yorZRut1JK1gfbwGbxwWs4c+sd7Y49
sBuZ1m/F1GjfV4pQbuAA/rlyPgUDWm+OnfZhAQTF2xQPah8+3TAiCkO+kgz7VwUD
CW26b7gdsmgXH4IZF7hSgIZkXWX7Tsdw5sTI5SsmxA3HCtKhJoDXjHzcioqx+Emq
PmDwmqfWlyvHXMA6iZIQFxhHdkbXa4Z0HIm+kdbARgO7gdAS4JaGRnuGJut7kKRW
7BB729WYc3HK7soegbqb/Lzc6sZ0SqE8nQb20WudBmLaprCQecinOqhitXAy3dae
9JcDG0eqCaGgc2SZ3UcdIQSuIKpwTk4u+dkv6Ns4X3O2dxvIAuP9iCPJ5jr8a3kO
1Q5/ydaYKUdPSc7IC3BmMlE7buqYonybTPTbJbyPtVZOyTn2XoTGtuhXm+jr9zUG
+XK38LupTRYNsNZQQBPAgzqFvSYYyr4sPURMGU1DHxX5dOL+MVa7PCeshOiRC3p4
+pjTQXkrPEFEueNuYb1Q7zlCn8gQNgBv4cc7JjK6D7k4PYCsDfSl2fF9OaJxOFc1
+gm1l0OjFMbbf85pvFlaSNKXsGbzFjzSCpSAhuOuIkbpM2KPxdDvtGWu6GvioUKI
3sUuzjV9ChsII0Notj8a4EV8JBnpGfFvWJuKWxCcApbxpnsr3Zds9mEeGszlxhIb
288BlI6HyAlaBBd4hkeWxRlfCVikxyZNrAPbvugQyqwJ/FZh2QcqO5oyJaiLVxZ1
ij80+d8ZiR7WEwxIEOglFj4vNceFrDh/VWS99swujkBy7wbLyqTZG+aihuzEU2LZ
lM69rehRKoGDsvTSADAy5qdw5H6BycjkjoRP9txcsoLhNsF1Of52vaz5CY8zrV0Y
EImoUlkNtNaLc3nJ/U+6sEz43Ysmb9D6cX8S3EkFSwRcOZo+kxDHtwDsR2rYOPeM
dd3fDMJcluzv2TnRBIJPwC1sFCafuEoh+Znh7YH5q9eIY5GymrC6oDJYy1KbfAqy
5a4RmFitxT0enV9bBSfv/R1/57fuFtdz33MOAoQZ9xEZ2d/3oOTGNnwYbVybsZf+
TcYqJualZPbemv05djIsDykd5hlIWIwjojqZtU8zeJOjFlqG23yiSnUzI5zUn7eh
ilUGonI/D3IJ/BMUvfnnCjTj5nNer/eCYuI+QsVVvE45PXxnDxxWK5U2p2vE2I9c
IbWwuRHpVoX8CpZqNMVpyoNmBd3cOZ+I4hmkC/ESxg/+RcQQW6jzGxxuumh9jxPq
/i6wCJdYHh8Okyb4z0qe5Af18SWlLlAWhyGh420YBCUbOr728XJaU+u1NaEYA5bH
Uo1koSCtnYtED2Ser1X5a28t+WacBJeQiDWYaSCza7csuuV2ghvjtppLIVj6+iIL
lSx/1u1iSbKcQrmdNlZks2ELn6mBD6VjkaAxjraW2Tfa3PIx8qtBWbdptQ0N9IWX
IoFkFWDBeebo+Uf3V6PD35ZOl6b9pCifj2n3rr4dO0ToQLdARZPHmxAx50a6PizO
6UOfvR7gKRfdIgn7a2ygjT+5Otw3IZeHYnwriKuFIFtdtrZV2RHwkZW753UG3j30
8z1pCO4XmcPUPP2y0s1d+SHHliUPNIvkIc+gccX08YBO1Dsly9rvnTLy6UHWJif4
6u0aGAQ6dCjeUxjGOo7mWFM/NlNN2sPzG6Vyq36+IozYdIdx4gHKngTUcXG2Rj7O
2IuDIWuOCjDEQpbdmmxLYTt8y/passlNXEcvra7GZSaROHG+78673B9sb9vXvZ9Z
zloD69VLLtfJV3s4OW+kYMP5CC6LnZESZbDfYN89ZHBG4zqgpzS910NoJwvFDlSs
KYLOf66dmn9oLo+47lLUfxgJX3nfA8gTmyz6uWqjkY88gaBhABXMdp3IgLIDIuPY
vo2X6qDlqjDrB62ab1BZjEroNQmhJcSU1/RIEs8aHDnHpaso+Rwqk0CH9508lj+q
KCQD0Sb1OpDvHWOf1Hmy8onMQImRf9F7LjFlr5sgVGHsxn74Xu/5Ql0IcpTT8uXa
jA5MPHorskor5oBa9ZCPSQlL+rjPIGN3w7k1jXI6kykIjUSA5PMJzA3mwjX2A+rq
s8ISP5PolQMCg0GhobFn5H0dpGTl/dbE25eVskdr/NcOgd8csXOxL8lNDPDCHSg+
4T7JB/t1Yza8twKueaQO42y+BVqqdBgvq9OAEgFdaEaB1x96h28ZOMq0Y0pc4Qoc
JRArwx4y0XgkMeJ3jRmRbw4lx4EwbfbsCtg6RmpyZpCckV46/VnxfVvDcue/Gi47
0D+QWr8pIKJWqhRYWPsFQ0Y/MGLMAG0aR4m/JRad0mJXRlQ6+j+q/QFcDBpago4I
tclxiREuZqrje73TrGAoAPGV1+kEUp7i/U7z9KHoUzSxHxAtf7P5Bi1qRMe2cRlH
CWYCCG3C7FKtNgDQaZ+/Eg9aJkDda2t4C7RmZrI2da7dr1X3q0wP5r4276Y33H4D
Dy8QoW2c0Mrxi47tvWFvtNEr4YVPOPSWMRC69LBuftW6lfUmdKwBLzjRaCKzWZwL
ENKyikYmspfrS6cc9a4ZT2meMIHxvhGzVkYZfPLALQ4NCbENGn4s2Ol4b0d+kXvk
r6uXSsohqmsSNXPIHgfrlcoWxUzOYg50lVC1+7pJvyemOwtu71VAzDtm0o80qLZf
K7pOVa2wUH9BaEIMYhjBlNDEZ7BswUd4wD7cPh7LXRfUvWMcpG+UTAf32Jb0zKIB
l6TB1MPvIXJK992tZK1i/MXrqYYZOLZs1HLA3tFOYMRBCb52AtZ1jqw2ecSbRyoa
j8xGECY1Os9TboNKehJ6Si2JrSSihZeSzvnwvwtXWhSfpRX8mx0mHgo6EUE/xjTY
FhD78/8vHN00LjqYsL0IYLw/CCSIfezhLuI7+tMVQQgMmFvJlhCsE61cWL7h3R6w
Gbwv3waA6MtSu/dP9A0w7YWpBnSCXRa0tVk8Oxe1VQdK9H1xPglknS5+u7Yv055l
fij/oQmd+W8uLhGSNq6wdhQKbsyzg4qEWRLl3KHiVFLXgaqJAUnzCNpfityCpmW7
7SKHpvkUhzRk2Jfnon6TMKCt7/1H9vzW0J8P07rz+5s//C4YVO2A25jbNfRVKOLh
P2zH7jeUutHFGuxJnT7wmK5SUajlnoo+wEWZa1ysqotLVevCc7P7qzt9zMAw48fa
6lRZPH+39aN0qyw5gerCEjPIU0AHM3suSspLlz8FX3gn2zamUb/rpnIUmLHpPsLV
VNj+SgY1/HebjVNyQZnuvLruJ6tnB9f42gXAfSI9YkmB9EM+YeZHLwz4k9yDaewl
AsIF7t+tLIDDkvD4yfsdDfymSJrbCaBKwnVJJNm7qyZklF/ortPFnq6nacBEFtP3
+gTkGoo9oApMJmEuPRm69+qDOB0U+gBw9Gnqc7gZg2hhgQ5xYcBrjPBEDfp2ivaG
kreAQSbWKbry7S5mzjchIvX0VBpMfPE58Maj6SyUYa3l41zHuDWWfAYjS4bb6FPK
EmTfCLf19RiYajXtFtpOJsnMP/Q3S1nok7yRL/K7Iyw6UQWUXKOsBd8pa4keCpl8
reiNc5g75Q+NqSCzGasg3sAU7pBxQvlEirBfBWXGKPXu+BrkJN64LgiH7kJTTpVH
NSNinsr0ahIfS5q1iPXHNrHiB3H0HMy2YUCQg1/UmwB35AvrVIiYWhNwkCQonS1o
qX61nGEj4i+T/H+drZ2NJRG64m5F5mndHvL/jwvcyqOVL+gHodyUkRnvzA1qnoA1
NdmLv/0o/BHLEWvYY3X8oLefYEbZ/RheXB9w661rlYc3CfOSahYseSOtkp1QAeRc
F8gn6nocws40GE/2hyYxZGEp6HAFjUpgcjJWYjOwkGdM7/PulzLKDaTGOAXMS8pF
n4I6AgSIUSjbjg3n33cD35W8RPqjQYRwllV7rAHOnkw8rW/qvBhSX5sTZg7g3O5+
zJZCCY8VWA09gIOSCG7m80RgsProYuZoFWQ2eJxHHYhJ7J3E7EU3WAIacRu4ouxX
VQsU4wjy2vfh+Eo36RVUeK7Hx4SzNbvPGjcof8Dgn6/KirJsEjMREurfDe6Rod9p
0o08Jaq44bC6zQt4AwxJ/YwUsYQHslHnVTyFcygDk9GqgnAWNZBI1kTQVWstdyL/
/prd0VAL5fQNBXNJIbDlo7epUIOsbOaV1IUpyuVILPjz4JdU1PYAv+pXY9PlXb8W
Rh7ad7M4rkH/5vW+8uP570ipHAzJ3AtGMhvBjJ2hANT4JcAHcD5+FR/L6lcpKq+/
8gcQwaKyiZJXO7sVfThuFyWKhOUwEk+jf81ustPvPcfJCKNcjRXkhi6+X8vg66TB
UH2hmE8tJVA/fbBuVExcnTdJWSDXDRSDHX8SmvqtLJV/U5W3WOHpcENUjaMQuoFa
Afz0uteYfC84Y1b00treZ1CmZJ+IiaY/CbhEVetrA0x+qK4cmrD1cILwkv5yPQCF
r6sptrQLQ95zJXCguHN/6uuMjOao6ec6dJizWo04zLfsGOTQ2e0t4PfnkuWoZiYi
W8AfwXwxZsGmi7Td7l0H6Rklt7rODD+4GuxJ1N8Or/Ryz6GDftlZ6jW9YzWBEMoJ
SeRkMkz4U1US52+rxQb2S9WhQ/8vkBVXKvRA3REEiSHZQi5dJwppAP+6y7jrgiho
KfOBSKFkcuyD9kPT9ND8T1qDAAXk34Td3SY3z81IROdmtjOXx1sG+EZmSiKG95Jm
aBUrqwn6qJe1Jc2AoEkaylLjGZya3wYkLejB1M5q+4X5M2TjzY+S2No1OuCoQnTE
KmLbggwyjCayYaqcbOwAOttZV90LBfgCWcz4ckQ3G2JKbV9xhetPz2zX9WNKD3Xi
O7E9jS5egiUoRBszIPF0ocENR8hqrjDoaLBQjnMkVuNckxcWz9GexSmH1ZGGQAWF
veEFiTV+8aAgJufRUx/jEEpJnaLi0ifXq9tefdPrR//Ajn2pcIx7NcAMxhZZKklG
N6aTh1DzR8Tvs08zmO7+eSKXJJiGE/KcWSMZdiaWW7Jpp5YeDGXZvCngh5JNu/yj
VNYe/jITssM93NYy1HecNlmBLf5alpl9Kr6zqCwIti3OIFGuBRvouy6l7QQcJFsI
s7PZE89fCemXxzClImb8a7jTqraMK7QpTFvJrRaQT4s1tXRlX3st73aWGXo7ZHUR
BrkK+NPbAk9X6NVbP66UH/u5YXV74HjtDrtIsVEoX1I+o8/fuBxfCGZqIqoUUfr2
XEQovexhZDhmiYgcwElot+zj90FQ2iSKbDotE2Pg2TOFKtMlv3jkYoocEu4RDZhj
tCf0Gr9MDLf8x1kmdFfVnU4BgenvoN+FAhn/nGoY4JzltZCXYGobifYB9NOKBW7p
9Oide/fsYeOmwAek7s2pZVVfEZ5aioDgyZFaH3vlhea0xRYOKnR+5DRloDls5uug
ebtsecI9HafKKP04XvT44Wlb9ZTsdONZ34Rnz1XLQnBhom2YU1ow2C6zLjHXITuB
yB7xS54lSmn4hgoqNogSY1eJ+dQQ4yApLCNFpBdIe9cICpd6WBBa52c6tKHKZzfm
aUJYEVjdqr8Dw18n0acow4k05lkE8YVi3mSTGkTUzU/QcKD1W7hS2Ug0Oi8UHssW
qiYhT/41CXPcugH64iZqqEadXUQlU8wwkmjwbx/lu2N8QThwND6KbTwCbu3gHRu/
kgkL/rLYkRxBiayO7DcMVPvW842tYUN3YU7CsY7pFWZ2+u3nCf0NP6sCD8e1kWnz
hElNcoMJyk2nOqmwQ3mVrcf/z+8cN2L8g221y/4pA/LxbYZofnJumZp9WQecPNoJ
x4V89wYLqLNpOfumqKr+p4NMOVsetQ0a8sXYqpijOtZAUZY22LdrrI31uFS1fKy8
90Qt9MJCJce8NCtP2tOGoijr9k7QiMImX1qQTz+bYyQfTGaeOgUjdvRJ/mSW4lXz
/hFvACiztT/s7iLaMaonUZ0CZzljzVzITOvGY28r2Iy/R4PI/pk2EPdL3CRB1ZQj
t5KTA2pzIrjYp2h6TiEioCtxDNNTP2//xgjB6248J4iHo0OjOo5NyvrPSQOw3SAV
XO2Pdl4mYsqbLSr2lqbJ8xAssezLFGNLbGhD/3+UUP+j9AKDm6R0uGGWPJDrVgV2
AUYgpIe+AZB1iK3T882zkUlYp3rWEwIidQdPr6Qg6hTle9O3blzQUhbQg7S47fJi
eSct1W/tyV/z8eQzANUWQunXISjRLlLm5ZbNYRQXi4+7whVjDRuziMiW5tRxlgCK
ppzRkAM5OBzX2TGyOC6S1j5MNUDwLQDlfuEcwsqJc1/OLZR+zuOdo4NLVevnPnYN
jdZpPeqGh8waycb9ftTN17W2S4skcWURQxJXYJw/BL84tB2otZxOcZhR5zsIecot
osR+j+yC4a33d77Nszilaz/CX0CPnhqPELS9jqbMwnTiDptixlQtL/D1q1IjvxLv
L9GtYFuCITRDdfBDQH7jjvUY69TGTGvh/XhEoPkHrnlNRiRooGDEvUjyCfFMdmnW
v/rkfuRMsOND3A/V3D6ye63+vG5zixtUBuC6DovPHiGy+UTsMDTUxp1tJGhPFSwR
ZV1wN0Yd2Am517bXpggzRsG5MrAdcHfAM7p0/VAZEcszbNa2zFd2dMnU0EbDiBZt
DtxrN1AGfldqbxHIs+pt59Q9t2ej6YEc96I/3sIgcAV/o4n8KEYr8kiWUXp1s5/E
F6auWGqoHZrpQnC8V/0LCUhOVshqIdPqcbSsxnAouNU1oaplXKHZkphijl58fhuC
Ry/cNXp116CWgFi4xy3yOMHLzpLeFesVwLnraJ1PvM80GTelpe5V/fSMcykZX+k8
+48MQMvGsrq8DMXsRI40QhEkB2P4Z+3jiMziJ/9bZ8g7zlUrkr4qnLf1eLq7iWCT
tvQoiovDuH4PZkv5aI7TYwjgDwvKQaRFmFTubCLDDmOBnJk+La9VZJG+dhFy7X0H
xjeUUZEHqA3daG5Y2ODQUy6HLAi6Xd0XS600Sm6Nhjn6erXBs10/iA5bVjM8bsdp
HaMCz2BD3hEmJOsgk5k1HDZSFaher5VXrwBb1JrUfzokGHnvSu7kxFu2UAqThYpU
089kKjWn59YIEvPHCtIbtNi2c8bLpIxX/1PkZq6CpmfBwkx15BOAgYgQDEhFn7tB
A0j93Nv5Jqpx+7ARBNtYYv/5aZfmShU0t4A4oMqwBqzxxirr5NhGORMfZ+QbvJwo
d/tKA2NeXPdPFlMDR/XaPkvq+f0E3wByGjcKY5Nk2wQaIRDDochAI/6BkW5hSM+R
lycpNgLLI5F8S+mp6CUURZsVhIN+XkkB+kNMOtYIDGiOpl0YdjHr3JppJlKFe73n
3U0FE6Jnq+fRqtehliywlKzSExuvICXAV2pVU/f6uNryhb7Qjb9YLLRoc8BEsWtm
vNA6khW2oaf/gWqfvde/6K3xa0E36LC3yFxUfWPPv7ot8ynCaxzsPokFJJWd9p+t
uyrje0ChjTPM1vD0Kfj4i3uOy+o5Rm57NwO/DGSCh6lh5XNvUA/874eY87SYV/c7
MjlzZZ4kddnD+hRu2HebujR1bvqeuLYSRFJDTWIwdJEpxNXM76XtBm93tUtl9iUM
ofjvPikue55fxu6SC63zn4MlZSEle/owbwtGUEwkV0yvEqFx+Q50Lr1l1jq6omsW
hvK1LTexGpFhWuDvcRJ/+aqy6fwu+HVct7I3XI1CEmaPnwXmXbaR/Gnofw+Kthmv
Lmfxd056MAb/u6ED+cJYhWMcQo6dDX7xHBZu6lzRLYRSMLZSaFdrQ5XovlW9Zda/
6EWhIrj56RxS0Yxa5YcAkuRhDigAtSrCrJcty8NHWN/eeV1uzkrQAhzMd7sCt/gD
5oTOfJSbsW7bzuSVGRLSvBu901CoZZAV9sLCtQKBOPILoxkrAvcUGtJqJyIxs2IB
LyCeu4T8jZp8EwkFl4ls9A7VjWZWWUFhShYj8baTyOBZ1pjXd988SZEsMBmoodYT
prxgy/DRR2bpRvLMuOeNeecY6jWKIYp82OQVem40V5hMUDAHg2KGOdfsvqjJF5Ct
hNKLcqwObNf/fM9+ZJNYTE+MvVX3O5eC600dT3driElFA4W2fZi4SXbtYnohMbjv
aWqokMJYOj2pnjKNvQea6fHsvD9xSIN5iJiZqI+EIVZyRgHxkBm1shTrvXj3I/P1
8rc/8XA3GvBMJzgO+R0YYPyOor2UZNvY0cMOaatcdnEXN790MXAtvFXVrCuwBzXE
8SJIrvkrnvZZi1qKEBl9F2FeZKcOre6pv83KVuaPI/H4Bqk0+AhOtvWFpOpAAQTg
NJZDvxSNkhiXzA7Xq32G3gA+bFmHgfMtiXxS0/x3E6IRDygZ8hfsjEhwgEIZIiEJ
glC84akIz6x3CVKa1zPI0+7+rGqqv75ACheAELe5QluCYQfh6XhbPqqsjEIjfXxy
IRrWlwUbu5QIZ0iqvSg0ryC16yaRVF7xikpXvEXhC6zLq7b6zVXhp6VQD2Zhz6xG
oJ8Sr6p53M9Z4fkb0IKq105SjtRJBerzpxYUBgUKSS4sHF/S0EIwWhEwpLg87sjy
mdU4yVtV4Sa2afMq1z9yXO6eOOm2YMSaaLwUcBiDlNiFAURBEytfWb19mZo6BsEV
cyK4Brhx2wGuAi1r48liQUj36F+hMRzz5JcVn7DEpZsBHsigT4GGkLR9sFEElMYQ
x5mQtnXJJ9slzTsYdR6ri5/KQiGBS/KaiZrsVOWe8Yj+xpwWVfPsLojzEyJlpZiN
DSNUhDE8i3PjKyOfeWOqFUqC4b+jn9bQ2bXM1clhdyvAcPl+G00+kA4tT/R1n7fh
L5ok0oxgHCWPa206tYvz4N4bWXA0A0nUABeAVxftQTEwvwVelS8q/gaXTczxkQhW
PjcmXIx3G2vSt6g3naB9juzWolaeSUmRpZsW1H+hjaTlyy9QDvwGtTw0foRYInkt
nVjWDNNOYh74QniS7AXEq8j9rJwes+B4b9yAk8AcidWz9wZDeMqxrs8IgLRriB5r
5+Ez20yPAjouTUKgUosOEU77+fv8FSxEuQfzt2YqV38O6rv8yFZpwQxsFpYH87D8
YXjEGYBEKOYKdcVuGtyHX3YV2NZw+hhlnmSW3XGWT0YJYt0ViGg2kJo/8l9BQafF
amqMdqvi4kEFKCLJJISrncr+J383K9lzEygCHwotyOzmD4Owsw1I5cB18fEGCJ1M
WFiAgEzokM34T8yVgHkFEKhAj1Cqls1+JR7Yxf6gCtOqqIteSQ0CFRDZOLcLDX29
cHIMKkt+9WV7tfbF7h49Dw+W78pJT3PtQWGbHLrhJX6Rsitc4Yjy0WfgJAkb/Q8B
WVSMbK+fZt58RtlGHebQldgG705FxIMKkZ+ccWR1eGtIzgE1+a+MEFGnZ0UboRN7
ce34zPonUaBtX84hjXccn8M9knqZdzDq5RVP2R+oAwvP9R259Y23bHj6p5+ZgDX/
KUxHa5uYKT+2H29pAm/+d1dTbq4JmDdN8bsgEx2AdPZYwYfZ6LLI2Wb0AghfYvbJ
76k8f7Qd0HfSLB7T4/YBswnkEAvhmyyfdUoekM8LInZ+SdXTx4o7OOQQ1EknlZgE
8ClHk9fLFjyBKWK2jsg3YhYJob5JRZmyrG/TjYLL9DLershThoQ3opI+d3+WQNvX
mO4Wyi8nCg/sWnE0h0hEhzxnr0aafdj6mOMcEWW/jEWr6iLVA42XgcT0/FAeR9nI
hAfZ0Qe/h/2PMgsoAe0hxtqHuQFJuQ1gJfBWJX0yZ0ofaHRDgTOtKEtYGpAou6Q2
T+yAqzSBSJE0wndrQmV0QdcTCokqUrCmDbIpPeuCPovWfm4juZtLGTNArxjd33mV
QSrqg+w3v6UyveutOeX4Rgy2wWE4qacqBPYJnhazwL9KMIvPZQQw7LRgudUts+WQ
/lJtcYyyjhOvAM22/kw+h0yfuRFZxmzHI8bjg2GuStRyjF68zcyBaBWrW2sDX5Hs
g70uTEI6nS7QR+7JK1ooJXpstm5fmjVa55sre1EC6Y/tg0tifvN/S6o5sP0o3kRx
RbRpKcJc9ZlwBzLjC8oRx7c9rFVtFak+FBW9Yn2as4HANT/2DzTqAISvjJgNWqC6
TAoqiJTJy/jxnCIiENAMQS8csw/n2gws/fCrhFMPAy7+Hq3TuEhJc5v2md4H0Qho
Y5mNn8Nqb8HjgmLLNfgu1rytArNfqDKCULi9vqvDXcfScqO+XdJxzTVXogYRbg17
i5+V59F733Paq9TfVQugjrZn2eBPWXIVUp7BDchGsb+ORg4tUC/x4haj799N1l95
hk4ffQe8UHDP55v1RieeTGFFFB8FLkohOIYrTptiL59SaHbi4bETomaFr/j5OGRi
i0yZoIK9IB8ykZzOy32eZa0oGCNgZQEnLUoxz98Kx2/+pn7MsLr8zUtCuJQoAm8b
tNumbzAexEehDFCDP+MevJ+BrhudmjPKsFdLt3BBesJ493Mkprda+y7+Yn+IzgYI
kM23DYKNVSZ2eqf4uC/cfoBBvQwcLf6CGMOZoc9+7nkXQxGFK3IkPUWpBaV87srT
XkIgxJUO7uneSfxnN0kXj4u9mRj7NCUODNhE4l2N6yEBuqH/KyWbbpprvpX3s9+K
Rh/kCEIW0nHLK2DHAZ7e7QMbI+a3Pogo3LXtlgs6jGOxCRunyo6EfW82PC2i5Ff6
6eftAvSdsFjrAnZoO+6XFRLTueijuV97sM9OoqJPuap7YzhO6Kra+6HGAZwxBMYZ
zkQPPxdyMh7S2UnXAihF86KGPurpC/OIu+9amxD7BClVgt5XAQfPCwILb+6w+Wsk
0hJlf/EEbGBvNEpnRAG1vuGTXS0kDihphoAntYWqhaibNI4c/TINBrHva/HOiZEj
zeIqBlbAlu2dIPxnGIg4U/dB7Yn3YI0XJmAIIEkPXJXpXtbkrot9HmhSFFm0XyQF
hGhGy36FjANHhZ4ptUHMEhFSwYvm7N3O1GKOIQJCbPgOI6cJU+nxhJXitXXk+Flg
beT9OeRDP0KaHu/kWe0tbnH39mT0rVoFMWvGj6IK6tVl7JMlXuw+A4HS13cbvHzE
RqCxfUPVv4aETYS8K7Mh6ZQVR5cPnu5avSZcxGHEQk4tmEceu7I4g2iiiV0XJAOA
Z3JNncKbT6gjr03BHHk/4SWYtvb6ZN7K7rXy0W7av+fgJ/4dynqxHiuLMFcZZINN
pqnYc5CcnHpP5//+cj3FrlkJh09qWDEJMwQfE8neqLysE4nygTDd+K/rRStjnRmY
dsau0KUZXnurEr1qnMoDoERhR7h4KSpel8XWi9YuVluPT6shslcQ0TNNPuQtEAck
+umip+VIXVd8h1Vu/mJmFK+sZCfwtLDI+BthhYBfKcyhy6pPxCp1qJgHgARoWUN8
FYYrsxq+0P1Ge/NMuc1zW58o6jc1SPWq3d/ITDW8Ukt6VuEentjygTPpST/OMw+I
qF3D+H0w7Xu0+pTn3wpJD8FSH46o7GdxKDbqa7gWWPWa9hloQywiWiXLKIXFfap9
qn1NcIUrGr6YoR6tY+CHaXcWb5HuIj4QA3q4e03XCiiGinQcwaE3MZmR6s5dI4VN
HwxOFT8HgN/DjmxtAkad4eQpEp8NpcNei/SIwTfahl0Bj4pt+O8XIDg1W/YWS/Zi
r4S0oNoDY1VZFPn6PL2VdfJ49YyDToH/vNBxr7xrd9MIJj/0Jzl2/JTXRE+p77bt
coTzltjABq74Vw3dUTy3EjFsdhfG2HmDLjRBWmtAwJlxXeDUD/c7BAa71llVP+DN
v2T4+cH9k9Qf0fYS+hZWOhZTUWN5YUnSLTIOjCyWFzrxo5Bvd4Qu4x17J+IVJiwN
H4H0oVCQt4SvPWHbTU8jmZvf+bJEHYDvTVnauIo/IStpI6pClH2RnN6gEl4c5epE
4wthWJk+zKTloY1eprvVo+RFum3Fk7pHKFYzPoIqlQvcAjzw203lq/1paMeyhvy4
aioCBMqItCl68Tb0OXySi4rzLCngSeLrTJMYfuuEwNUR81Tl2qWM6QqD393YgnYP
tWFp8KM3cxe8c3yhy7Y9Ozs4dKBgRn0QT8weh11ohqN8r3Bq1HOHFUYySS3j7GUL
et0trCFvj8++7O0R0rvkyYUXGWxhpfh4mnJwZ8BklZsZvC2lJBGY6LgbTTGll3V3
oSBgH3QDGcDuCslLhhfXOuK36WZWFTgi9Kn0NGTjQLYFBIm79vP4mshMXMbETITY
hh2xkvzLtEBB9UuUIlfVy7Of2LFzY+hVrptqPiBIIBkULG2LeawlVAoTWWKxjIlT
SJHRcHil/3pSROHyTrxJ6SylG0ZvnmF+cNu/RPe6tMONP2QMnCZggk+1e+Jt50tE
cEKY0V23M6T1fc45ga6MLTdCrsls+svAT76Si+0AFgkjgfIGArqGTmoPkVDkX+c2
orAf/ckiSoWdHCRm0pLxQ00vJrk8eCpngcxIKI9NhZAkK2lwBnxJ1PGJWM7pfFZN
WpY9SlLcn3FP/D0rRxtJudzMDb2MGSAU6RoQN7JQTz4JxqniGi93cJbgHdQCpJvW
IfMBRnP2VAi+tD7l6AeqV5FPmr6hy4GRUjyFJdwHoRcIKjojJUUotrqtEZuUN1V7
TQx9b6kN9YIwVqWNvt6XK8g/Q1t2vE8tyM7T8qZktPfoIAr9bP3jvS/Nzvd5NPo/
Rd7iQ+jUZWAzwTMGwdHTVPp8oLe2xEcbfAGd86aqnzA2ZVfM9oWMrKObkfKHhs5c
zN3uhAWfZLwfPmrSihhqBoVMTBT1Ro/C6vNqIOxSvgHu0XLv7dstNA5hOQwzY19w
UgAf3HuYk6H9P5c/bS4EQmZ7iC+FxNT/4eknIgSXDB0jJdVLoE6xv/9/JlTsrGj3
NloPP0ON/zcdP/6yzTUA9YXYp4W2J/pdEE7TQy9S7axuQYEksj+gIitAweZpuFZf
eOLR3/DlGYuN+KcMfQQjAI1DbukjtcJ18f8sTqFYgqrGOeszBvMu9866Q5nXbMPy
E/TMUThsX1rTBZY+TJ1dkgNvA3zuvXPS7KzYm7u3Fm4nH0iapDOjdrYYKIbzG1wf
F2yYl3tJY7zTjBLql1uvzdMmkHbYwPxTzJfdQUjfc1Hh6W4+FA97BixdmilH+BFr
25ppyBDygkhKvZtS+Z90K8C8tgR7jOYcjbcv7E+FIMzmZrHflRhMkYgiiO36FlZV
LvgzA0I571l60oQCrm2ICw0O1sYdYv/s1yTxYwbBDzIJREVAuJ0zs71Oc20wRitW
D0cbtNMd14fpPvdofoRKM929aqbcrgdfUlEgrDHX3d/lB0fX/vCFEQMHdZl9SFzm
u0IkSOpCRtI/mgyRKVcJu6jLbVfPDppUDDACqVoRBMDYVM1fL9JNT3v81Biz0aZZ
pka7c4z2Nh8UnMHSDi8/TirNra2XK783cO7yPTrZQwEkzO9rVRI6t5xH08Q/C5gX
kVZXmko9c34aLk8gpyDjB89n2Zd4xFiH0BIJB9wkoUYtGuV3oFf5YnD+1fsgdghw
kqgOk1p4xuoJ7tUCIRSDu960v85f9TWUb3Kw88nsxH8GQETrV7tiwO1Cp0jp2aTB
njVEFa8X7dh9oABbHa9Jn4JGb0KAatNxnSktbf1N3cz9F0oPsLzsx7tgzDPJ6dJ1
k7vdHp/ftJGoALPYqxHKXobp7OuGb6OeGo//cmCVVevpt/g7MtloNNcBfRqT1d1f
MR9GajSwOyHn6lBnKkuutH1lBO96tJTuXy2yP7s1AzC5SuuyIRqzpRO27bepE1O/
F+6z7ZiLLwgUCpil5/crKgSEqVax0FsTHci/NmTosUQbjxqzIlY9DEfoEBp1HEpA
0MysqfF5uJ9Kq7mpV8iU+/lSARiupjznr/L0Yd1+P6o7BVuA/tDcJhMAzB7VaC4V
4bZZz1LSzq2mF2f+PE/oSkX3MMnmWDDTRxMQr1rNIQ/g9FXqUOBAC2fYPKTjii03
eog1K7unknzMplJ4p8WtUV0bzFhsajQHGpdVq47xkJigfq6mkdeqH6fOzwoDOBuX
6d39RJ3Tg6Ix8GduYEnqNV9fhibnekQUBuK7R4zcXhjzgXUyhOBYmEX/NE9wjOQ5
3PqIeXZ1RW5fuqxlc6nCgeTo3OrU0pnaM2yOnoSOSstQDScTgsKPkoaEo38eEv/z
xEeLx/1z2S45TbZfFqT51WbDXFj0W41+wQXoURw2k5rKLTqe24OEoKp65lBKf5r/
Psd82byVXR9gi+eHm+n9JQbkLe/fCm2mCXubnh3VX+rD5E0EF9V4M+LuK4NmLml1
ZO6ADh7Ck07yyxVdkXPpqLnX/VlxJRI02rpgJmMF2Ur+5cOWWKfg1hY/5D+BvD07
sZCL18eJrJc+r33044pv3BvSKM6HR9sm9Zpeb8FX7UmqsryA+oaE8HJ/uW8H2BDC
Mx3DKxlERAJzSLwdvEq5q9aQ5ElniVTUiYCXuHkSYfjVas5aX6yY/NY1ZUKW6kU2
x07J/RCZD/jyJgfMEpl8oVwjaHqRGqlVQ8AmhEoaEa1W2c27O999nFHMW+p5irpG
XLVqoGGHkCJWYkoN+smTE1S/eg31dfOExzVZAsyUXWbtP1fZeuyfq0Hsbj0AQ81w
D5dkT3admENSLkJoVCom7hzLGr76PwfwQ9JG42FrzcVkJhrm9Hb7d5ytdldRGMfw
Gu/qmLB8smIFGQArNOj+Xu0mt3V+qg3JC6Yi4wRsNLxtR9Ql6eaDqGEcm4InRHfR
qqlQWtbir8OCOW/38PfXTA5ytiyAg9ueL/kUdD90WHEH2mm09P2s4DOpRGGxz9F5
NUzY3eJhMDFV6pZsjbKxdzogK7EKOGdWoOTcUC12m9FMBJCMAW4HgwqdgaBZip9g
l6kZfIpx6SxKdGtHNxT50KDG5zcJLOlBsiBLyj8xXY7zoclTW7GkkHQHnJ24dSZF
YQz4y89oAB3kagUwPlWNHcFjH9bHeLJygO2uLPk9RjVluJJSrWzAsmGonU2+Pl3S
6cGsVwGPQ+i/v8bg8M+Wv/RINppPPFp4GUVoCVzcW3d412K/AcWx1Zw3rFEucbeZ
kUDkScBGzOZKAghqomSA8r9V+2lKrZTeBNI1VhT31Rb3h8E/t9ug9xOOSz2WAaNj
6cIri/iDnXV/F6iAajo63z+DYHP9Pl5PBoTEQhPnFofwBtt+QxTsuhxeH8u/j5Y8
NWPuntLCpIFKI6BM2wMoJFqbPC0bOUIaS1mBTr4rCjbtn9btQ+GwH4fG4TUvPRDu
aEUuO8Xu9cjooWmtJjzWMhdLRR820DPKSsk+bOnCcjklD3RE08vZXP6HeI+rpWXY
xqAPsg7owT338TAde7xAFUIaHIaegbv8szdR4juCCA97b0J8nwOjQ8F6qw0UE3OC
rwn9SZyX1D6L66aezqGTWkGT7dKK+6NzQ62qZFwIi1HHiRDPdsQQg1X2I1VY465Q
d7q1VwnbkgjICX0o4AnkomZOAptb7jUhc0o0traWUcmtxsuHTB0lcBCbQQRg+73h
/NMfdu4rNWyu9noIK8+Qxe+VPUIBUjC2h/VKtBuT6elrkKq3f5b7GO3Qgagbh4xF
gRlblCUfl1UpCrJCz+P8AzibsYQZyCGXpd2xz+IQjabBuLfJkkKOhW9+yOWT+ksL
y8KPtLytscHGvepITJYlldf2UvNAWdG04CIEEj9NRLGLsDCNUxoQwK2+MD7FkBLy
jrt9S4+acUy6hygFNuPJrxidGaLdAlvgnND+TNXhOqkOBuIAeaZK6Yd9Gw+SHqWr
iL5exXL/guO8t1UDZWFaDQU23HteNhJC+tE4UdDjV89SweNIxLR8r7/KZJ1/81Ko
5+j1/7dsEDPSNFePg5wNPv2k0pTq5FT7mTufLNkeYaJMb6Ys8T9sTMyPJF9qjx/g
DMdF2i3do9zXuFYgrRs19KKbLqnxn/6pOD0LSeqOcNVODlO8BoH1aEh+gAcK2iqT
RzylhLdqbnU+y6zGzXUmWeWuLExh7QJfT5HAVk0rw/M/tB33tjqdIByS/gWnczXX
6sEphDuaB80vT6Ol0nVJjmMGl9Ypt5LbKwWu5cYZr2xadvXs4X8YZsWcIotEbfCJ
6orVVjsIRGG8GWWX9cRGmQ8IDgbuTOVCadmlkY0albmBdlagJi1RJBcYuTD+UsZY
wugcQ1/Zmkgd74340ov355X4Aj0yGPKI3PK8PSdQewCb0m2JXh6mah5JSazJbUYz
QLuAbs7FG4fVO8lx27P9NizvQ8t35HBqcu4FElq01x4rQY+5E3jLmAfITxQXofAQ
tdh6ByuDroViPqGpeUgsxvR3uwjBrvgUp2relIa0koVwTq4NSzfEU8yhIU97/1Wr
aDT27bdSCR7W4+uqZjjNfewFpKoiHAaugn46FWnVdUqh/dG5jq6ZqBIT4ksKoeKS
jIF1+cHixXmFbfjBe7FX7oki4mt8E6rwcUftfEf4/u8cTllk7hjGdo9QxvpLyoFi
qIxz5QjIg4QuDWzGUCPqzvAt544NWue7Ddah5rRL27rOnEagAj4j7UzP2FQTAVxT
sjaDT9TRuf25kOpEz9GnjRo9zu3p1q4ULwhZrv9rckP6FSRX0vOTakMQ5kATamS/
h0WiVgqDWl+3+qAO0PT2zNFUk7/pQQVYmZvkOY97tM1aFrekhNLCyhVmWuuzbIJ+
rzNZxcybm+v5Dm8CHowbm6jZL8IJViiBFdfT9cmsQ2+h8SHwq+YkcQh7dr/vtwMu
8uzVaK389l4sC7UmG9hHF97nluRf364HuBMIKV8qRDsDXriMofCqkpRerHgtGO5u
qeXTygTk7LrX1CpOGUzhoVQbak4ittBPrDS2slCklce8H4K8ePXWxKFtY8oE1+lp
BGv4xLDAuS4sI5hGo910DLyVziuN+/OneVzhx1ooNPxc2sb45oyJCWFKe+6U/c80
DK7SXfeGOQn43jMCTLP27yfEMM79z2uMOLqRe/wBIyuvO53+KD7lgfq+DZdBjfId
bqLRQ3E7AxeabTnVju2aSWlE0qGx49pbCBghiIu+vreETjXjUfzfmQz7dZFmp5ue
M2ankZW3x6zHmVPjhw+V34iVxww9/LbOmUkI2BctgY5yQE42iiDiIgwbA7CrBrzb
2nWPiS1KaRDGhXncGe9ZcLjO2KU+OFAktQj7a4Vkfzf3+0KXZZyn32tFbbWQ9DBG
0QYx4Fhs4bmAxLhVqcMUPbV2vSesmJ3yZAFxjYWTOME50bROWzfBTxJSC2gkx7JV
uoW4J3E2QkYbIByhVu7m9PBzphrj5Zp0tr577sr3rL3fiMuxkvd/YK6qxSXcBRRh
0WWqHYuyTSBWKCjyBDJargpsl1hRNr5R8kziaNO01j2h6ImL1x4Wte0zg9CHP+GZ
JQj4SpozsO1ur0WgSl2c1+FthG5Sp3gApMyehKqp4+v+3wS4dl2lzk4h/QH74afN
G2jx8ztg6IvwabftGxBObr6c05+EHuCcXPWtLKiFCbdL9w5PZawN3/TtO9RevB4u
gRCoCE7oFucPd/ZS0LYUToDjig8hqMCu6msDQ8H7Jqc+UOXkrOcv+GQVPbkpelOr
KOkTzpBMPfI2J3hFkgOE/8rInoJLL3AYKuCkBJ2cG/c1Mi4GBJlvJMy4Zm+y3oeT
DedBAgmtV/hjSP5y0WN61vJQQMT/TpcGbhYT73jRpS/n42TmxJa+V3C91VmdD0va
M3FILA7wEq4BdMTS5J1HEArm/RiYMfumd9W4JM9AmXVi2O3ovrurGMgchSPk2ikL
s2l2+IdqrHhYRREjKBur4lnklN4kaLgrUJ0nPkkQBA1mK8HKQ8T9g2NvW5CtiFVn
OWMy9TCt2FXI5jr14zvHliKm3PJXPxPYvhj3e/b/Dd90cDlFTkiqaAX5aeje4eKl
+X4AtrA3KoPlB8xayqSa/+xs6in55NJ6STb+Jps0cdOzESU+DLTFWKJhqIpfqymZ
mhcUwI73ayONwSiRBP/OMeDbLgK36sHeX4VwcB7ahHaufksU7W3rfRKE8zZuOB6d
JpKQefCvemE2bg5W1CrdV0C9VmySL7qMhYMlnB7NfGrH07NyJOkfH8ny87hRoVQ0
g+o0OV/mSquzF4sV7Ugfc69Q9Lh175WbZhx4BDAn4sMj7qvIeHcElJRedEjSpik9
AwUGoQZ6+1gprHiezC5e6hDYcC4RGMaHdvzTue0dIxIuc8/wqjgQi0dAfLdj3OCE
7kipiI8i+zXAEnCandyyFIhwDUxhlWpS4SsUN5bmUf/efJi9ws91fDETcX9Si0LM
oRPdVmbZ2jtPQMtdsB36qzgJ9pvdg/Prw6LpIiUnUZyoraJmV47yuVPYUtJqgyJE
HehPLOrUOYgffPSbINWUlFquFXah/fzpTTGXdmJExC2GlXWRhjjEu/C1tzK/I/JO
bmoN9qND9hwH1YccCbPQ6r6mtNAS6ZYSWRpkoNNh7Ue0zVa6DCznAMZiYrEthJdH
DvQXPwFWzjALFVolDa7oDOu1kXW2Lzb/xFn0musKfTNQFfALvYMXyk7gOH7vA7QU
vwhfbAiUpXGNg7mrvNYndt/0n+aNNtast5Lh8t8VUmJ9TH8h/LO9lQiXwS69zSQ1
QWC2K2dAMklE6Z/uD4yl5oPWaFZfZAEr/Erb2UnWk1wZ7vjqi3tHc4zVrSScoD6A
Ci3DtgbEtN4k65vTlvbhLiUNHLKjbgfKs78LVhknOC/Y5hS3ZwFBVV1ysuhcWy68
ZTVNnS7v+fzcmi6h/e68QE5ZkY0OaR6MT/3WS5zNKurtIA7351lUqVUs08T5MQvn
AWT81Dma2sYUvFn7g+V1J6HV3fL++gUkNOj6kFnNYgc7Y0iDPMy0MOY5iayAFjOG
+F/+RpaPGMoWFOZ4o0qlz/zS70UTjWB0GDpXGCaRhU4NutNyaFVG43bt0wXHwowH
+uE9N+VtILB5q9fHWNxeVanFtlxcPrqvpOwj47gTGCY0bSolzVxB/0CkMKTOvu//
J7UtTHXnunr97J9UxC0lYaSIHEfclcpM/EjUHy5fvoVzh0eFg5aGSAVmcK7T8kOH
pVE4O1aLCNk9lFup1zQrMZPaFq0/zgv0NqTwodXnynzMxERAfj9ANk9blsgaqSKz
np7xd21C+G8AheUnk5FdUNRejlNd84eeNNp/meaRP2w0pTyfHnj1+BGxJMVHBRZA
bWMEmpj9KtizuedInWUwNKZyGFFzUzq7JT49MtO0KytWSjpyZr5QQR4eTFG90W4u
cars+fqEXih4n60TLI5Nd3P8+IjrLZY4T1H4u/RBHE6igt+TZPacEN2QsuEu2pZH
K8DibPCITJXMc/Vue5SygFJE1XGelkxBvY4qCEEFPHpRuapbaGo72gmPL04BCDy0
s1SIO79QXewF+GxdYD69aLps+TE9bux0P+DsPjytUNxCnY1Bb57KqIIMiELzUrI/
zHq9jALIs5ADLNqbgV3wUb3S6GhwqYFsST4uZbkD7Gptrd3ln81bMeoGKypx8mT+
2Hdo010RN5apzEjevqQ2PkOoofxNdq5Q+yV6sDyQq3fGbUAFWcxwsPWktC1SE1t2
ph7rnqJd43osJnh4gAtwSLDMhQiLen6mx4PxygvAxUVr9CnFkk4Qg/zjzCJnS9W8
YueLiy0+uQ2UnaoDxVUfX+WnbYfyvxvDknTuHoy5c1p5p92QlD9iZvN3qs+HnybG
LhtmCtRpJ4qUiqfbYhJiWv7y3S0VEXbR/vEmOoPiAIVA8uoMhsgT0UaQCcYsOWL/
N86OznmkhpiCOx/mo4B5LjnL03CCohcVXjom6igK3iMdURPDqxBsCAnd00G3GgjH
oe20xPDzq4z6XJ4DdVQKu/Yto2+nG7E3uAlnt+2VuYZ+82qZnW1Owpzb7fZXasn5
Ope2ZPvYEc4fK+JUNL34qxDGUrnZhGkwC28eZZcl5/d6tl8Bt6qMB0Cc8k5fQVQ8
BYZRwzu6oc/DHR3gEuJD/dypWGyicCITs5TfzXkLAtlNqsehUem2T2YK3QVvyywq
IByktyaMqIZFMLPuF7jM15XsSkTC99IxucLPlQsBD05Pu+rFzPS9cjZiCICD3WHy
k2n2zBvrDw7sCSTs+pR2hgClXflBxmiWFNEWaJNMoK9ivTD5j1gE9ERGyH6KKjIv
rZGxxlqW8+GsvDkFYMG8mKSJX7y09R4xRw4giMJ0sZBBBdkBN2g5V/TG1dPmqAyH
1u+hvXK6xsF235isjl/jIV7nL+cZUM6rjqbe+ahWo6M8x6G/9yjvluM4NRh/zB4g
YRI+ti+njlnb8aZdlPvABt0LtSd+tfrT+vvCKclM/PN8/M6fAQhgsz9WQvLpDeW8
bjvqnGPDppe06d3Ti+4C18jilBmYLW7aKbakQG15sqvD6G09+JDB1uH1qVWEM+7V
FueSCkf4DI5mn4ttR0qSK4mqlzQPirCFMMQ5TylhdifwfxH/iayEWYpVG4xojY+4
L6BjAxj/peJDysrj4yz6XQi0mg7pEwN4ShNW30+EGEMgeSSMVghhNoPYSteIIv5s
3EmUnrj21DOETuJOnZ4tVUw7wGiAlm7UayRUlbrOJ57lJBYSloYXoQhb4QKNFIJR
IlghpHxpxu6SIXBAXTJRe/Xg8/nQb/W1FIDR8S+l+w7am2w1+RDzIE21DskdTXcw
lNVMSnsn6jvVASYbEGVLx2sW7EqAiCnk2E4ofXrqs4Gujv6LtUDtjrMBE5UPj8tX
gBYeydE0ZQJfZE97yj1odnYS7tMGen8aeJwVxoWlegibHy2wEZ5Zuc2X734WSRGN
jWfYyxt+qcIImBQBi1APFMIKNcCKKIwTl/5g0xI0ekndpdKrBiBkOxUBn20gYraP
uCHXRIQjozSK+lp2Arw2j+WM8v199FycQNEBXAUds+1gztpcWFsKvKAfPxHoq5oO
9spVzIJ2Xx6hhokfFpFP/fLZh+HwZE7RFoiTmNV77r3/MphNmICeHqBxkxMxuApQ
pBNIhhFCxfAVegFtwTEikPlzdl+F77jwSrkxYvt4SVEhCW1weF2OI1zveqaUBdcG
TUrc4Iag6AUH7TaY93meOYUHU2BdaFeW562zuSe0jvV6p1BDUkYLaJS6nJQLJBS+
eMUcEl2Sb/qTfCJGBxoFix4HqHHWzBx5QdPWphlYBa8gQPAO+IDpFhnylKDQ1FE+
nqM8iNdfEJA3MXMO9PSMcK6cqvdVnhxNBf25l/P/uM99U39BhdegAOgASp+zHt6p
QynxbziK/xQKpZU8bUAGSWverRVvwq+7OB2ax3jKSLXRWr+peUs55NN09rwoPXd2
IW92Pou/9IWwih+LJm+BpidQ0kU+z7pAzpDt2KtbjBakDoo57/IzUWC+wbcaIsEF
waofBeKMeUxDTVDoQlZjJSJC0k46QdOYmAJ9KxipVIOrVtI+pWVeNQQaj0sXya3x
oUARLWv+O2HlltCmtiCKZqnzMx1DvjCCqjLCay1c8NiKa5TNVzNJguGju39Xb7Pp
rZgMvn/n25ZaGukorgxO+J6LyllB0YhtCFpy8ubfqwwAQuQLeRdw+yoUsbve5ijw
0yrqSWQNnihk3fs2hDWNQjEaCXH3TZ6cM+5f71n63T0cp43eWVGCexwjD0bPfj5L
6XkuYL4Gw/ezJ4Slf9snt7JwoXuJ5g60Lc2WaW1BUYdcr/GV1wp1CjosqBkgT55L
vC+3VTcIjvtO2DkEwPSfjuzXVLhV6rHyzvTpGa5c+bGeWuZckW33MXhSMV2kXGIF
cKxE7ZabYvwQZzbPpHKpDA/lAxNDHT89QstTYD3PjdfIon1mbedmWLXNDNKMV21t
wn9PggvZGN3PKJ8pboK4Bts6n7DKm7YxJBqqvpYCUhLvYWz0q97im07R2s3THWwV
eVOxhyVqslxltBnTUtJULNRHJqA66cHBCV6y5/Nl4wrz/Ha6hbqGz5Zuy/efj40A
YwQOdKuJVLjHpDKU8gNi2Q8YdtDeotrgfo8P/sRzd8KKGO2Id88KUNb17VCWd56r
GDEbY5W36ymmWdzGnzdOtW2TXs67Ha5q2p0AzbyUB26we3UZfFZk3yPLiSIycSY7
zgroONgRb//HoazqsoiPzGjZiUlbHeW7I55yJukTMy4Rwr4nhLWxJvg/nFDE8d7O
iTP15THuZMsVx2/KsW8jW3/4Fz0b2ckkWReSW7KWjQGLmdCR72Tv7IfialdvNggR
LqFXHFqBRfsHRV0XxTGu9fkAjibGlmadTs4nfS+kY7q6fh2FCAUF68MHANZTbCMT
g0fbrD0J2iQyi4rUeTKQQawFmVxAsneWvnziylK9bScN4ac7/rYOTlBAyw41SwYO
lhPk3uBbo8ItLNzn1JBZouDsrEYCcLVEC/0yRVrBf+EpL0xJy4ni7qtYLY/H06gB
CML6lKmOsSp9MYXPBWUxbjVO5XplMni4DuBBd1JK5K1NXqSG73YYYVUp4UhnB4Ke
tRZ3YdBpKVLUigjWUKpdp69nZIcEcFVKgVr1q7o0hv5sB6NRf6YHCETU551BkbS+
uzgAnDhZq5PEoE/CJhxCtXturEbvZkdp5pqp0EJq1fzWpNEckrC/nnPxKkAQxDkf
XB65+GenkHi888/GsWOqgeUh8ccdZ8NPlQ1UGUTIiWMlyESybgTY8gW43LJnBI66
8Jvz+gi48sunJIHpSoO+mIFRjfGbCfEpyWMiiAaowhsuxcxU5JcsutyXce4x72Ch
kwdH1dtM+JRR8t+yyBiePH/PmKt2qI93zGUuCIP35g936YS4Te+DQZDWYRTQLHrU
4CyDOWlDM5Xu3Cfq+MpBpqR7HpRPKqXsKHdeAJJYyzUtWPqhv2d0GoqluVrGreDJ
f/L45mTHjQ1hPUmpr1z4eG5bVoRlO/GTtk1yD4YZxdKOcgGOGGuKLorflT0xCtYg
2C8Vvz0kJHvqdVVyslQWsryyCdb6yIm+iVr/L7Qvz++VpoRmAlB7NihfXenFiOd2
yqEnkcMyaSHHWW2PoEy7vDO2uwLItclBbD87WWzFD8fqbfT2sHRZMuoJvPlaUOj+
344qSwPj9z8ONNjIt0d1/nHVoU5IDu2b3+8xpYFt1HdSyR+KQZr281GyVc/Gl19m
kVWQSY2oUV6B+VUIGUF1xKWecHH9WVz9H/P4Paz+VxqR9eC1ziuXkJ/1QGgJOTmx
xbPB57nlIBT2o0sx/XEfx7GeIher0XILwmkJO3HM+2Ytf+Rih7iSBTAx958YGnez
3vdMYGIopa5QaWvfxcquogEqFD0/uV85mKDca2J4FsMbiaEo0I389SOOwgWH8Xjl
Sb+IgzbzKEKbP4V5eHiEsMcrC5LmeQ165t/X2j7tqm3Uh611jQdRVeMGEqD5/dVZ
l3WWIICYHs5M/Acazfnn9c842thOXfgliMDgIXABJo+aws0HjCCXaUZWoUomjzGy
vzUdv3A80gYpi8xShC4kj2Hm/FJFJCZafisLRJWazzMC+KELrpgyqIUWKDAl5gZu
pDwJr2QNgMjckLtOu0CEFiqYHFlQVcLls+vs9NWWjSA51UC8ItqGAKe9PyR94gT3
WTljWKpqFxGWMX/hSk9sPNByOIaCVvAyWWhygt0NDgEditUU7jRJohAe2CbBJPny
AXWXdx/a1qfxHwGyXLS5Y5m89xtn2W37ChBqc0fZ789RDD35gp87dqG1v3550U/U
a925KUlwTOsvExQSTinWGNZqi/vtb2eR6Vwvuk5Euer7vIQXU/iQRYFCcav5Xg7R
+jRBxub1LX1MHFtQaeUstR4T9iYlXpd0uNaNA+XcV6AHBTFJ46CQ/ikmvt9Gb4N2
Vyucq7HTiqCAGJ5LOKGM+UXy5Ua1U3/qa+TIOe3yzo8SfY17maRfgtupyuUkWJAO
knkmQQHnROnb+ceR7x+sAEtGXpuY+qU6jLMM5+/a2foa/WwA33hHt/NbWPEq0Va7
evC1yxN0o7CSXU5Zdo6Wn1IvmCJwmZv6DwHUxJ0BM/bz4i9oqkMELScu3P184PDP
f3BxXIPGXcoeVQv1qhQ0hbX5yGWH2kX5NmzRok8gGEh1T91LkKjthY3S6CwY7xlr
HZ7iZw8oplTvRji1hONoaBNhCbRfzWzGQWpsUF+r9uVFmf4fXdKoTjpN7UsOrDvv
8s1baS+INhmnjLtpf/8PwvvdQqM9tHBe16SSBn0/anc1KUCebbfv6nwevmpu74RX
eUgO59otm8yU+3kqMD3jOKACNLD42vP3A7y7WdsL9VlCjxIWBUE7ZyP6CAUVQ2ba
dgvTrxddvhOmuEilK/KuSC8U9ckLmXii6m6rdfN/MFHUyv2E348S3czeQ5LiHJS6
zkM+iNY/Q5ZhQBXSho2L2+EgGQ0+hLGgmpk6s8qR3TqZecNhFvkQf8rY62bgHCzm
NOOB5/5q43hiXtwyXhc1n6FmR6cw3p1m6dAdtIOeVH+BqlX+KF6ehLfHv0d7/VTe
Z6+Io8lIDkC9J1oO/vtiFP3ffsdZFxAIaBiTo73zmZT6+4EwbddJqsa/G2+PPbet
KYgJijGanDd+ueshNjnBmIfrOxIHtttmvaNuCGX+5clZccoygdnWRd7PuyKEeB5u
iiWy/lxoFtb2Ah2CTw3WrlvAjBaWVKm3SwTRThvBZk+XtfAgUrG/Y2hBcocUQKQB
aa3WCQse7+7wCjsT9BpZOCr8R31Lj0pwbTrwL3xNIj4i5cOIUCVKq+rD9sKQFnX6
WIJwPHL8oVxq6n1zqdpWdegYtJiIfrxnZAtC40UE6bcMk1nLrVdQ7MIyqEsiUt0v
4lNqLEFeUGocv+uhAgfTZoVzEAOOL0CGXXcmdf2z/iuYOErdEXAcLyjihQcc7Tlq
cmgd3fK+kayTkOpL8W9P9Exr8gVeWNUL6AaakW3JU2NrgGh8rHZfNTamxcRYvbo2
JaaXw3PrFPWfxEDBZ+A3J4yJd7MBgNIX7A/xg8poNJLoBT2HSyKsxmVvyZ77vsrK
ZFVLJcd+5PcaVCYSo7nZXeSkmhdspDj3WRt2XvKU6iWDMigDI8ZXR5XVmd6XjH2n
RHZyP06RWpXhzFR7emJe6d3bwwakVTa4Riyn/LC4lhcLGA54/hTd13UqwloYmfEB
ggTadeRhWG7nRS8Wk8Q/B0Uo0ktz6Mab4ERIwYcLKz07f4arywnP5dyermmdtGV2
6m0TmHFrwNpLd9WsHI+W+yaT0dwnIN4J2/9C9Jofu714d8sDlPM1IQn1iJoEZzRp
IRdDePvKKZpNwENxxjWjnQOhxzhurFzIjiqVDKVg2twKBpk0S+EyaA0nrMJm3x/z
RarPQm47uYEUbTE1gV/VA2FifM1j3wguS9RMHgrxqlK2FzindEpWL4tsVQhY09Kz
McqrWAgtB1XMTFnpPLZ3xI2kVfi5lSL7FbWb5i1ltRkBmxdXWcRE/RPHg2OBjckR
oOmUu5h+bB1zBznPPzQDY6CO7otBaaCw2MotxW5Vg19umAHPGCWUfLWLeuCdcNrx
eR6Wq8vir31FpvRKM0TM1WhOVm33Y3lNpIslqiEdU8hCIrSz/b/yrjG7DIHwuldr
QdbGoTx+Lx01Itt5TsxMO2pnmZJmo96PVNM3dbCuRWFBDmAH6OAJ6CsGo9PF05yx
b0gh0KwLUVsBhrAIajT/WY8riEAAC7W9HVgBVgEApg7Hh9r4XsYBNjdaNkFS3CZf
r4FSWbwfJKKbN8EUG26elFJt4M3kDigOfkxJ+0is1gjDPYzmInvyZoN8a99RjooO
NMpSJ6EazOIRKaZvyHFq6+7TNrBI3TyGk7jXqaN+2IihQQB11Qpuemjr0m7FVW8e
fl+18kCQ/PEwvT1l492ThvZZ77/SRsCYRB1Nb9XkL3Mu0yETWYmLrZQGjcG/zaqg
9pfDy+3YIwqDHEtysoZJxCwo3dzuDT4zWWCg0qyoIwBkkI0w0tdpRWAs21r1ykTM
Ar0WfICMFrNXD2cKLr1jE6j7+S9pZUyx4Dfuu72/TXkG5Gxp+p0esH4NUiQPZcMK
WnOZS1NbwHhpzuRv/SuGTYUrb72VHFQCtRmXv5QrPG8DLP8Ig2JE3A9uTo0oDLnu
ctujHHMdShKGzBebx2bW9Ou8yBvAeFT8wOzmAjyD73v4LZRI2x0x6K1+4KZTkM13
jBHUJF62vqEv6HlQq00HmKO41btqvw5RnQbtYAn2zgzrI0Gg5KEZhXUT10cYZ3nf
KRVQU1OFS117eVLJySZhhrK789eIU3UbJsPHjrQZeN6KP7TSUslw5UJ/e+IdHvHB
gPUxModc5qtsJOMiNoU59rSO2CTd3GfvjbcHDKy9g0ZFFQnvz8nJtvg3Wob2NePj
XPYdBDJBbSuIob/8Epo3Lj7+5HkjozPQQc/ColgwF4/wTMOheTryI/1sq3VZKbpJ
WdhdU1WC8Ig8Dbrz6PNCuD5nh6BL4Y9hxNNNnkItpZlnY61Wpe08Vm+BF7Y9e2eA
GvD3eCUQis+5emodgaWQsEphKhq2p2IQDaGvZk5kI/Eljys+lB8S1Gavpbi9EPz+
TRAoTfrZ2MZI5+PqMxNRvECMiM4oGnczfdBqtTZERzoEtrEBmhm1wK+lbZ/4iiru
U9vBnrIHdAKoZ20/JBjKCDwzB7MzkXxDtCba9zHYgRuYYP+pTcDMUi//+bCan5uI
1DteoLiLLU+mBx/tB/oY85mu6RvmPMck0bm+wipJiZx3x43la17KFf/zqu5nEsuz
xANxlxcr0EuQzRgDlYKR34+7eA+wE3HLufSBirfy2B7hmYoEo12oB7bHWEFNlNIp
MwzmX3w6p7FbA1iUVWDXMW4cI9eue/yLa8pB8GjKSPw3JueowjdNvRs3HSAsaJ6M
1jydLOZ5B44E7Dw756ZhQ9K+GSI/H/KPiajOiHdJEKKL7d/stEq9TPPO25QMAq5o
lgaQ6hXJCOJALMzmWc4vvnX3YDhc/HdG0Bvypq8o9wUWifOxw4veHDNBCQioSra8
efukfm3Kjzqgd246F7FunVgA/AYikeTHED+N5UNLG6PHBfNZm8vn2/OXjTiervv4
eG2/ZPsU6Vg+m9gIMmkWWVIiFh6Ff7kBu2TiwHr53A1AfVITa/K1CzSmAhZSwaQA
bJGOdAkOvoJlDKLsbx4arYkki5FngqZXqzRhEJhyJ407Cf/5dlgKXVS2GK6hKsVW
Ou9Cl29HwL57lvjXdgVvB1fFa4SbNAPbLl3eoTbtFt8GOstlLDAHM5CBpU4Imv61
jk/RPfKwWX+RP3EBd2MTvuvIck/Na/USiceE7q+K/LgS+NgKO7+8Q0TNbOY/hih8
xgMuNYDM/i+OgjnjMXcAYf8R8qGORtDhFd2/RDFIaePp3sKnXG7qE6ZyYWgMQjnv
paTyYcup0VHA6oi7jTw4lSpnwziWJ7uQ9VU7rBvDFRNnl/uWeJUjkjw0+hSuHBdp
Y6ZXX+Z8bkEUkobbEp7tLxtWBpi1VRFn8u2+0oKKajScINfRs4dHsPEzghioay9E
rNSjBLvFAMIHiO3MEN9iSNy8mFk+v+ISjwIfgFsDB1l+5WSf4Xh1djPuajJHzoTO
gW1tVeKGCt54WzD5bT9gzqQxEcpJbGHD6GUpoFujlL92r3XpRq/Ygq2e95CQf0Cr
nJzuxGgkr4ixmUdpMjFWBt/qXTRGZhqB4rKeKtysBcUD+uBj71jKIXr/vNRXUNOr
8Oy5UkN+Yp+AIvyWtCgScbLEm+ihg9COptHp26wyOs8NoIMOSH4y49Do96BH14kh
SAxDdwYbiOhLQDiGWTp1peqqDNE113REPMPO9hR9JrD5GGdIm5425CZIDgiq4erL
/pKPY+Acb0F17lDH7NkVZAbmqlLFWYMjNx8o2N2nTWb/iTXIucZdoQzLbX9uGlua
bE3KNyB/EQa9mpc4QvJlmUcY78QizN8l7J+LzQ+OH/jCANgbJ02HDwpJrmgFSNs7
QZWSPF06ocH8Xrb4l1cZMflCCK/voGPZqxaTiLnzLYs8JLmEM97AkWlPdodYSf5q
K26MGv8GbtxtPqF1Zvck0DbIwYWzLQJcAz80dbur1OzqwgFj4v6YKnaIjvpx9pkl
f3gIRbnreNIr6QOGzC7VXJJ134YcFXBaYxj0l4w1gMRZrSjRjJmDWsFK03NFJn/i
ZznoH1dEbYmRch1j0QNFgNlE8wtvF600yQWDd+X+5ty1QTX4EuOTDYnx8kVHT32g
HIDa6kN/+dCyW2/t2MUPV2eOeZvtJKI7rcNU9hK0ncrP/VOSUXh87HIi63fKHjRt
5jhyYYSGqE4KzXQbF4gWbpLhWA1DWOaEYAeiBjJyPmqROaCOyejBQbBXqAkijLhE
69H9yLngB3PIjxr+7VuEe2aemAN3ygUp7VKiqQhfYF6VCaqX/utnnP6cd8uRp8aj
EfPS2orQ0v4bHu3M8+kya6EbWrrdPogKCguZnbzqT0na3NgabMOa7ATZiAvtNw16
ffEgGWD42MgbJLNmhaxUasPT5MdGrYOQMKvVdKgy1DKOzfpyhXbcvdl2oHoX+46D
DgIUAfOILsQcOVBvyTEpzReG/p+mfmOFwOWanqSXRM1JlLzyxWTQ80wbJ1kCY3aM
unR05D4bnNDglsr9q0ihDsKvZlvwo5zhorb9aT1SvL+V/0Wd9qFYwZYI+YsmMuaQ
hCPmu8d/+MrliHw8jsz4EBTPlREjbY56B+C+HXTOWT3TTlb6hCnVwdP1CkALba/Y
vi/QhuxhGyHqtaGXJJmn2V9QWgtvmiVp0bXFT5YnFrWCJqD7+Lv1/XS/+JzHm6hk
oAbo3sluSpyAPuhgV//U3TQEKh32QhHiapGvwZqysNpHIQ4ltVepYKtPlnxEmln4
KZwNCTHGGEteJQHBq5Sx8AUFXkAj7MYpHkMP3UhlOi2rX5KZ3dbwU+2uB+fQZSAu
yStMcGlRTe6B/7EJS0TY/xXsDMxJT/2iDWL+iZHjsMzg5tfbnm/qkwJKiE/xrzLg
2o1sBTC+p3JT8vwU0LPdkgdKh3e79x2HNZjlp3csp4t+56iFwB0HWJWbdRw2KBgy
CnWRoDq9FIJkot4g0oqma/IvoJa0LUKClqjMHXD7dFfVTEwcpwUuAt4UlA15EszI
mK15Nmd2npgrTDihsdh/lddNkFrfJJHClvl3dtKRAg62k8oS5INDe3Hw8r3DOlOs
5gCRMs8WZw14PAExapFEu4HcdESu4FdP95FVw/h2PMvD8pgLYr7A+QEVpBU9DK7s
wJzi0CEB5Jc4+WPbXU1c8USh4XG/S21OFmATlJSVfyNlpmUrHjbKsBum6H7l/DZB
LlAx36oMYAT2jIT7BlYDZ/w9lrCPFuE2ENdflM4qKmFwM0CG8rycyi8D9wDMAdwL
iLRZdYR6eowFctZ5XfvqR7EV6Jz94gu++UFCZqHv0DxnjT9fQRnzsulusT0TQ/vx
fk1H6tI0B1trig7kQILBgA8YxsxsOpyKjqj0WFhtkWSajnb2mfnDxsMET67ubP76
SefKPJvy6gnfvd8/J0ViKOMXGTuFRLfApxKX2QRaRhfJp6pJNDP1vH1ertfQ0qq8
7OG0jtyeVVmrgoob4tKke29tX8UoyoJeRIvJw77lSLcvYXyDnxP58Hddy+eOlAq6
EKDKLPlZfs7ZBNGRDcwBCwKoHQACXmn+SSKCu6TD6m+SHsAen50zGw0KszFDZo6V
oas4iOv4bXycmgaSwooFyZzxl/GgdeF6fpUg6KBxpErXVJLfXpiGTq0Wph3D0IeQ
jLc1bDQy+MXDs85jjgEkv0kDtTYX+i2cWF/UdbqC+WPKJ3AlLKNoxBqN+Wb7a/N6
6ezGWEL0fCyvDEZHcfGrGSl+kz4caRGUjlGQ0KctiYQbaZjfMprEoyTDSgmX5NnU
3wLpIsoOPOIHZaySiULi5bNqdwODL73H24gaoO58sxsWJ/4ULSN7lqFkXaUZJo5f
UefRcGxptIRGLg4CtV71TNYFlQXSBTez3Sh1Zwun5g8H/zuckxZwku7WaK85ltP4
g8cAOOuAnqQZ8er7G7J9/MoGtWqO6hfYFGMJutBxLv7MzOMJGB6lgS75bBQ57i1W
CJxK9LEddt3qcB12jzRFpoLUQK5Du8tQv7TQ3xR5Ab79XPcNtkNO0YvmEW4uW8Lp
Gk7dAxLTzzHNe8qUKNk050LlywOaUKj+RqbnMM2KfIgMk8eFYgWkQtTnVVPzcexT
THflok5aAmbQIB37kYEqb2KSU9a0VqaKcD8gNWpDHiYZ7hMj9EE/Iv9q9/CrkgbQ
RSq8tBRoVhxNe/9YJhCFinnPjphPMZSZAJXEQZeKSipKk+RR3DobRhvkRENc/X1C
GReLE43+Ut0VLDVeknkYgTyIPuZTWGMAvQjkkOZ1YgXaVoH1+SqR68TWD78nZlv9
+orL195OZkqqoT38o4NXOC0frQBb0hXuIxK+WV3+gZytRoBSZQz4rRqdJjO7Vo4k
NkJzhxfRorkt9wo+h3hhuVv6h5cDm6l/toLLAyam7UFgSM70N+KNOzZU/h5kB3Cs
D9bQJo4FAC/6UT7A7Gh73oVQYsmyRInktXWitQ5naqZnK+k9GOHSWAhjvI1HpMGc
UuZmC3OhYsFf9yk4kJbKky8/HAOh/S6NA0+2OP5gndG0y7Zh8i/UAUUi63jFCmCQ
3RCVgW8bNRvpCiZ3CrappMH3Da7WZwECtUbWViPMhmSZgF464Yt2Pe/F7+N8fSWx
3qzHy8BWZhyacRthCs9/2WjXZ/+1ivOGmMUZZbOoXeA120Oa4wUIpXOHYLwEdlFA
OCvLgHhG4O2D4fQQ6ln1nICeAGdfD0KiYQVnSnj8Cwgb5/KxL3jLIgd13V6XCv5M
cVTbCcX3/qUu88q2usN92QAOtAd/eiyawqPNC0RJQv4Lm7z5yl0RR/ioyAgaTbv5
1WKwX/66tVc6nzir/whShCGIwGSWQW9rHaWJPIrs1q5XCObuxlCsXvzvIbTbDr11
DVMYA0NWs46aKT8mNQIOaN4acYSZhsfp89YyJQjTfQTMfjq56Caq4IhNp7mY8C7u
hJW783s9cj+hcvoo+H8U0Cp2fMbLgorfwr9PKlQtkzbawhBWNqYzkGmGdmNkOyvj
I4gcWGyjLG0x2MrbwPHCjuAPZw4JnjBkRA1KYRRElr5I/atwj13YI3pbU1rXFQ0q
7gmTxRxOgUyLlSuHsBPpLLlqr/fXLl2AvQ2aeeQ8fevlioyNLgztiLNJFL3lEaNW
CKZ/ydXYJ8CZ2OVb4FBN6Aa0I9Bmv0/V9yHkFeUxYgKhSUcCrVhYHiwUwH1H/N6x
t07xgumdAMqyBvoUSB5hjx7df0Osjcg6NTWIOLVtZlsGf2hGfhYp2OXf//w1Mhcq
+qUztw7Wewp7fKTHaKG4NO2q4z5oL0iwK3tLP9eGlMSgrpPFe9ZP0UNFPhX86FVa
+p620QX3SAi2xNDA2TmKuSKFTq3cbo6yDSEwUIrqGqUJh0HJl8kOONF3C/p8fEr6
Hee6FfafE+YoXzrAZP97Tei+kdY90+E67g1fl6PQGZSrIHI+MxminxGC57gk1EWa
XiP5BURnIdZw4h36MpqXb5RVm0LZFyRuqV3N+9aCS9Gw1mCDnWNt30kMrlyONa3h
LgwRfDxXpHiiLZSMuUCYXKWi6jqi8FpUoWh2qrEBnIJX3uOyz8YfGO5R2G1c4p7H
0DJaA6V9lPVimXkFsAj1cS5JYWW5GuyOB3XoW8gFZLKAVw81IAt1RlI9pWFIWm0/
1TSfyO0kzRwofI5oytupW/DLg5qD6d9T7KDBYMudTF8uEXFoiE3KH0CakaZgerZz
PMwqjh7PY2LeApbdIOrYpy02GE7Rj3AdNrBZ470rE7byJrZD0v78aQWA1aBIJpY7
kgqkeWffVxt8zRrMlHz2/fMaQASoLrG4Tfx5E1GqhSpUocU84NAGV3wJPdOI2qt9
6C9XY1jsVoIsd+1Eo10c4ae6vLPqT0LXgbtI0UrmLuTjyzt7RmBUm1yv8+wwsIHO
sNcl8pp88zVVuOs64cI3ixrltBXqLqjvTE+lD4yR5pfqFEO+F6Hs+4uzFzqeFgMa
bEpkPTP34tIpb0ZLDoORG15zMYpZyqaPFAQjFlgP9sxU1pLORPgZkQXtrTPz9Gu4
gUg76BX7vIBhU1U30/n7Dp7gA8W7J8/eD/pCO5K9ZjS9pCj/I3DsrBkYszNYS1hK
6f3J55Yxnq+TJGGkD1bH8ifghG3nXn5QygfoY3BwCWZPDrXzzyasG7SjNaPo3oks
nPJN3PLyGJyrEBLbu66cv5W9Fk+WfkuwvdRpwxdbprXc/gPHhp98Hx+ACgYSojJR
RU4Q3oeycL9BsDEM45Qjm3eC5pKQSEJ6G4SBF4wSkvPXRX2viiv8/hwrEV9XFnfo
KGp3UFpX53fLAosEktJKZ932iNkZSs4tKxWUT+4aTuJkS/SNmFHqBIx3UCjbXv/R
6/s9WvVVoy+trfyfVER6Im2dfzieuV7TtQ1bVKytoKP7WYH3SBca7kBnsyGekdcR
tgm+JLfpPHZHHXJBfBo3llvvNZSGDql/N/SjJoWDZjMS7SiZPWfXhzoz1lKkQ9ix
h5m+wQboPThuPzVxrv8pFBvFnRCT57YkY/gUnb2PDEsz8P3xcfpnJErCFVaoHNQM
L1hCs0dRTEc8kNHXG/FpI5T9FfyTbjR3w4FFTcAgd9h2yZFH2ozWQAeVrVE6v+uB
/Jd/4/v0FQB0UwA6NNq25Q9MNw1uY+J1WflDd71BR9lF21oootP7KOu4x3cdfiec
kCoN3sVWERYGLUN6ZmV0DIXivuLSQiHaYu8d6OFsw79owqF9pJBOCtheBBWaGuFG
fWmhhBGvK27WZyhmibfvElN3BdsLXLyLIPxZw+M/mfXaDi1VXhqAPl8XIAl0d6Wq
OnVPzN7YH7Bd6wL5qjBT/G9vZ1HhhauuvpKt2cMp9ENS5Nqo9OX9fEtNzYHx6O86
0N8UGnnzJ8XRrOhU/uZuN+sOZFQ1nLwAWrxY/PRZu1/kDyGvkk9pxeGNKEaa9rRD
o4E1aTWinw4R9+H3NvG852yIa5J1mh3fvaOVR87HPbKpzvpWabBBPKshnzTjUqvm
09XayvhMrUMJloN6ZD6ndLX3hLViUUtRHbn15RRY+E5VJrfYuOBgZYM4Ss+zr8gE
P9Do9Td3oKiorxBIApS/kRcuS+ewwTZZSsADNa+YXVL8wkYQR/i7Bx3TzW3LLsj+
gi6L8alWpoQ8C7u5uMQ32YM/gb8lR6GiJ99QIORVWgoIVOgKASClGJa3V2xC9/gd
+UY4aJP0eMuZ/fuUd4fw2BO2kzbBoKDs6qKXSRNx6dRPVff2vkgN0kwv6Fzry6Gu
lB2AFOKVgIRzHhnOqb3tiX2whqy4540OgfUSbveJUalTxMB+dLyo9wI325b6pQAG
OPyaUTHB44Z7Agl+7JXUZR7X+vxBCsKP4om6U/6s2ZLDfOZFswq+3VgdvVix3plT
CkakU1xj3hPOIKE4PZu+1OKUv2sGq9qZGw9+brJ/p7cktkl+bXe3GsgkxnbHyMfo
ZXIubevcuPDkhiqPEZfjBXTXttsmGmTCbZ/Tprg0m4uvuyouWZ/0p+6/YYhsaRpQ
VdeibFxElqpN1+0QG5er/nH6knQd+GWC/qSiy4aP5EWRhHdtBEM5gjxNM6+fRKs3
XQfEOu0QyvNbd4LWn4WH9haBq8eEp1MgHIYXGorxy3v8HaKmzKlSM1IFcTVd1IWG
WAoaW0693vXq1mdg1jS7yvumvowTzCuPiDjMy/cz2sKbvL08puvvEPMmuHnp+6V6
/J0zbJo91KvuGLRKowk1TSbV9C4SrTQsKNE7MsOC2Ok5kIJKwUio3WEPGIjWchRk
6r0zFGykrXl0I3MCFBJneDTTdERUAPZTcCGzQq03Wt57bGBSyao07Dc9rVBSxqmT
ACujKWFHydJucBntlnWtw3x1r+6WOkLeYBUEKsZb+5wt+gcVOCK+WQZychzs5MQf
FFGW1iFALIRVhlXxNBFfabCoYQ4XHkxUGhdQItVcU9FExD+IdJq3CvgWneWxOStr
rhv4k1TM4v2/wL3sxcLiJ3cWXL1eAsYUBRsZ4Ox29csFoMWRErwEoNbpfvXqekO6
c/XyqUbDhsWJ2z9uoqiqVJDlmjntpwWEIrQ+d3efH5SLsZlMCJQUnFSOEVlnS02c
rMrVrRePnSS5hkvI2NZtm5ZG3U67ybKrG4SP2dS0WfIZjyJzOJ8PUaL1ZG6d5uQf
P9fpvZyrQtgt9r2ows5kfzgAFZ5ll9cPKbnyQPhM4sI/6YQKRdckpL+SO71brNlf
GwdqAcuIDo0TN2e3VudRjoB4cB5uklLTE+w0qiuf08jd+/IHl0Z9MWZ8D+7elr1V
+OsTX4v5xQP7i+LXZv+TTnGttFwi4j3/TttAAp3Y9ZsWHMC+YPsw4sOH6Fb6iQ2w
yNfULro4RntOP4jMZEyG5VmwWmn7KikyiPsXCnfyxszhXJL1BKdmKAkHqI8KcGVi
nw3iuFOrUEA6nKx5ExctGKrBHr2NlIusgKslSWRViE1695dI9/zljdbK9jiF59VU
bV/u7HNbTzQLJOQgXJQjjbT5ImuQER5gUcVzTyYt+4u7Mo1J4FBnlQFi+xCxwxaX
pIf4cd+/t0mDkd62weA4Da1Un7yQ1JoJHglxyI8rx+NeBr5B0ubi8aiGX8exfQGh
9XlzgbfEBeiCIBW8fwZ5pz3t75a0fa/f9NJtGx2nvkeSuuMSl3itfH19dEh0ieJ9
95pFHcqgTZEI3HUop3f8M7WTr+mlYBF7YHJ4xXA2gHd11qN2l+0xVA1sPnA3n9VG
PEfJXbe5r12h7aNOJ82FEyZAEKHimY/GmftcWPYrPbKRZTMcQWjPXFvbE9fFRDE8
qnexPVIw/J34osi9PhuSWp7T2gHB9TyT5zQX3j9p7rnWhc01LiiiTLCvjtzmztt4
w94WnPOuCsAk1ecOd7Cih/AHinllYx5RYcmy4bEKzyhnjg3WDkAvgJtfGxb2vogH
BVppwhSyeZYoCI6dSnyITdVxWUUHe/ME6TEfd0SHFZr1Wk70VKlRrBLSUvY1ZNXj
cuQuU4cL7hXGgcGiHbRzXOGEc1OkTSu2YNyTBSwAE0Pa9OwQMpzNjW17L0CJuoOy
GeKxecfFZph1A06kNXwRgSLb5duLY7wSjzzAd3zZR17NTKn4AgtLsv6KKKpwyQwM
G3lr8yrL+AT++gzEAm5W5AgAp99iOlG3T0bDyLudbYD7Sj0r2RtOebd6wcXilwt2
qTxFNnTBukZH01GQYlGAPkUki90vH/hMVluDXYVt9GzL6GWtexmVVrzJCLyUyOFO
cgQKdDGowINQkCZNgiswnhxTdNqsxJZ3VtKOd3Z73wg0UAc+ci5I/d/rCas8utsC
8/4EDgPo+hkXB43arzhLLDFSbUyr33W6Yd8n0dHc49uy0rwEYM2eaodjDvtBOtvE
ZlLJLJhyPArbrTDESIEk331gl9267eFcb/wIQeA3hLa6dgcXamjC77AfF8FZrad9
zE1nMeWw+yfgxrIFjLOu5R3AfON9WicsbpwjcM3x66JKVDs6EyeIQ9j2fTAvbdeK
2Y6f/hL0O9LZylTUuWw7uT2T6VPtuI0IVB9G1EKAX+1AJ56K49gK5VJADyX+AOl0
rVaKaTHQaD/PVhqyW4P75lw05v9vwZYNc1oW++MmT16tqniZWqBbaWavkUug6xud
BVhQujHK2D5xupf6J4Hx3gCZQwhzDmLKymdSTO3xA/DJR95aNFHwi1v3IdRq3DM1
Tlxnn1Pzyec5E5TK6vMY2BBSD9DjB2g5rZX+OKKeACkjclCUIGgeDWBydijmSEcD
ihQHAsvD9pVDAvL5G4tMd6JMYJ4gok0DfFy4s0wBw87I1Zq5RUwlJjwI9PRHiCw7
maBVxlAslglhWa6MYbXTE+Xfm5GwA0EMsia+rt8/e6/mknLJ1v4o5ylSUj5MCtph
lVQGz0xsEY89+iVTbx6Ns/5kUHcTomab9jtAhE9yUaHfWYBzBOeTWa49oK5Ka7d8
eIdsIKBVV7dTRha5aNL4tthNzVmrjf0RNvF0MqgH2e9tR4lxBgxSDbHE2GVD7ue+
jyELBg5LlaSJm9fHKqcaXmTW5vFWh8HxJDgErQIzmh0W737nWGhglKMKqklXjdKq
WBwTyN4U/kK2WZJO8/x91gogqWY+9y39CXxIhANrTr2jx3Cm08+fngMJt5xuea5i
CbT/a0Ps2ldyhKnFnzhJEsbpWxwMHtkAaQDbK4I2iUgMs/kXpTHdqy61I6EuthBW
5jP6qVuhAv2Cilp9KZ6hLOB9ku2IIyOmpMpfXJ8HKhtmRjgcFAhvSl89BSKcrpwg
q20Sz0TqBNkyvS0L/xluf0SzF10ZAPwGSGSvSf1De+AGHMyJGFShDpAEVB+5aFKp
B7je2RYlya4/WrtPhRGQ2nUov1EPgvQP++m6G6Xn+HG4fbvJNQONBKsCboFdsUxZ
fprd0LuP6/2JxIlOTYt/kclurOf2DN2109Ucg1PfRN8K+dWCMhMVidOg8WbfMMBE
ocYhmhX7qcNIz29yZyGZEBYH51S74s9P42aLjYT3BB23RHgRz0o7I53uEguJKgdC
YbtBER9kGeoxVwmN2UAEv3WgzhoUphqfOMBYmNaBs9r+TIu8bL08tnVMiOgRQxzV
EuSzoj9VM7uGWq6mc2UWLdyVt/ZO7+XycR1TF3cmwqoNsN08SXLEuluD3pvz5gbE
FV272r79wjmd/NJhHnqZg3ts7Wq72IT9yp2xDWxYycx4n8XWH+QqiVGDzRi8Bpvs
yxntvzRG4XUYiqNYLZ6HkD75XBfRmd/XOnoxQok1tq9NJRBhzgGJXKXOcMdaSmlB
IQwuUDm3KO/bFm1GzUlzvtmnB7qYaluauZ/osHwvAr7SUzLvL4+FK0jcknm2WETo
8fzrQ549gTONB0hAMh2G6b/MtQbgBYd64PfM3SNgjePXS16r52SAaUg0kATXJm06
SWTh+aDXmBfbUGieLgRsuS8hMlBAnkyuTfunamM3q9emN6+ad338YfikgSsCgKxe
eY2c5M3j8LaEJbaAlalfBgMxlI0P61MI59HZeUDvn5WsOpA6uZld3XJh/OUfWiV1
a+ZKGFc/A+wwNR/m9kaPid5YUsMCt3M+pTgh6+4191b0VP4L19i1HJWJt2SCFIa1
O42bt8xI4RxdNHJElpkojbx9xEAVm3XmhMeoASNaWf7SnpKebWcKzAPf+sWkZbNM
xvJ7LI7uXtdAahDwqugQifv7G581vzSd0RSywcdji5pvemz3x0U1sQ/66WgH/WBA
XI1FeDruQnJd1a0gjfzrOZz6EiIx46RaL/A1KLdAwVvZ6Mjz8gEAh5lAHUfxcuxP
Qsy7fP/iwiEcxPz0ftiTdc8cK05yxtW+3NQlVVj0mcmntgjUfr88pD0lxKwpnUUe
yetdkQpf3mez0rT8AnXD1O7Y9tfxyVxDUpvSVjXi8t+MOqwaJIuUsUEnF9iA00Sl
FZgBZ2ZdLyXXAStuSX0KEIqLr2Nm50bnqbIynZsZ5J55DrgyBEp3Db0Af2gCesCs
pzNO1SgtzoeHfcQQngbU1G4m2mgHS3pqmyILi4eLiqUlovKsb7chdQup8DhRPy7L
wp+3fp/omzK4QTTFQsfz3Ha0szR0F6PWe2RGNx53DsMCzmgCD/8RsHQ74xqiwLIA
WUsigDI15dwtU6mXRaHJo5fwG3AqpMXRAWZ9QHVJfkgwZ9v5olcWC6/Y58QLqNEG
83W/jHmI6nj8b9fg2Dh+pi7SzxYgOOXYAKXdCS3t6KXr5ZzHFYSktvnhtJFnRwKU
3cdVllgWVkqnnYgxUkx6YeoF4EPlzi3xSBi8FM6ln06FToKb+zDQO6gPh/8Has6+
DY170t9LLYoHaHyDvvos3Ev1FpKxlBbG09tCUjAPtc6UGgY6qqHpx0yPXFPgkTda
+V9hAUw07ZTDhcfMPvvDXjWC9EcCo6BRxnIirp0wB+xayEX3v7Y4kICDKm0rby1N
hjGkYzIHXMOoM0jL349Efsrtb1TLNDyBBCfiHUvPhzp85JJXJvIyVfNaKQXCCrPP
MkszXyQ+39IH5kmHO+/Vx4XAtYaev3LxyO3f2y5I51t/ndKezdOWEgtBeEQEXr9A
/lK08McygbeA/EvtRhag/d4B1F+zIv+I/RkXwS1Ckvarfi+tmAb9k/w55igFrGtN
bXr1oRLiJiXa3IaGCtJTnMu98nnjAgLhfF4fNg7QZZU12uszBeglJZpG4Rmg1eKT
mfXfrDw7Xf5jittl43WuTmxAWhkIb4Qxc7qwQc0tibIVh7IWb+QElM57FpaHaVqo
BWWqf9H/Y9MRDMrwiPYVO+Q8+RHx6wI/lnTF0nYHWTuq61cWi0kS6pR9Kw0IQwN/
i+Z+TpstivaOu5mXJsqYfXEvuHVwqcNuKdqPJCpn39/BnaK7fr5TspA2mrdigySt
gx6xaaTMd2hg1GfXHZ8mscJh01acweBwFzC/8qRqwENZ/EVBz1F+xDuV/wQ33ozt
33Z32lPR66hrZt29GOEA4nfAzY6rnwhVFHwsVEqwYnvdnRNlrO3HbQ1HRbx7E+Y7
Dx9SAgP9MEyloF4I3jq3BRMzgST52XgKvruhwqUXZzVbJ5cWSuVD18a++LJsHRHp
DNlFcRRNa8hJj54g7x0ZCPjlDm7UbjoUgZ4OtyuVpukkT/8LRgesXEal6BB5CbRZ
fyYoiKH0Jra7kHL01WR0vBHgRTYJBLFHEpfoTEJvT4QEt+uloVlG2enVMscC+y9x
n/myp9gf3+qr71YVrJCyAZqDXP262hDQh2VmdIgOhjj7R2hRKhcrwhQNZ5skO8P5
1QRxapsVQJME+dRUzojXa/eUW0rUMEF9GIBAfJ8KHzqorvtZzyTRdtB1zOFDz3W8
vqSx1Rs3sFU94N3ZWpvcz4oCeZagBYfR5FNL63lLaTHxyxE0MEIabcMDmJQo0Pjf
3IeETUXKmaSCGMnVS5/VfF0ABkcgY22NYMHAxbjstoHNMkwjvHXMjYOM7e2mA+tf
XDZOiLOAfJ7x/2EOs/oO6+L0UyhyFF+BxS9iS/xSvT6AeQKUHGtPBa8TSGNV4OD2
WHwMIQpnbdxKdLI8A7FcUWokoRNmvE5S3QjMUuOwB+/TKRui/MCYTKmqrM7T3Dz3
0B2/q1MlT6+DHQJNd0YEgyoklhF3QwnodN/Ui+oKcPlbuifQU6zMCiw8wtE7zKdE
mqRUu5k2eLjR+uq1yNXnZ90hkiSd1xf0KB/WEN0W2+wSYgRVb/Nc1qifR+XMi1/h
6YfPTctRotExK2FwRl38WQOgGiiCK7yjsjEWhqjroyFs0V7+THj58gRcaA/1xb0C
b8+W9sSSzhjYsss0jO3B7MR1cMInOUtBLXTLAM6qnfo1l36ajO9jlGcegxLDieL/
fDxdLArOQlBLOYSvTkE3rgLTBUYXmEjb05qeV8beCLJf+6r7oibxyKo4GgCgt7Ns
IPud17083BNq0O5X/esQoh5BmRWmhlZDI5/YjV4QLrWb/onPUzPY7oXtfmfLEwjd
ufetHh+lngZN7wVV5FWS4EG9GO4bXzBqviz4jEZRF6Ja0lpAPlrXhcTASsOHpLce
c0N1oyrb4L6AGrl5zUBBXl6UxilfI+QDSVbPtcerukpKB5n8cJYMsZXfSlPEQEbI
7PznORQwqcnBEsG+VdN6AvdcXcvCvjHM7tJhYZiOSQmQxLm4RaCF9Q3kEWnfVlIL
djE4J1T2L4LNGwyXODkbU3wcZ7XQ8/Swz/Wn2nrHyPIXDYnYhasjISNgiuQ9R4CI
KZ945mEuQVh//oDg+hheowx0LmepJn6lmKestaPoPRgjqZ4JBL1st69J+ixDnVOX
LTuxZMD6JtPDZmiavuq1szPP1tid7GYMq1MOKkIyC/Am4cKN0BNvGMtfJcSYDNZV
OcBvPE2pvJLYWdlFCprr2UcbXw+QmosdmsoERWrc4oiCchhxivK5W8ixDa197S1v
ulhMtMoz+SY9fvG94M0+TmfwmVhyf/3zM01AyEPGSy8OtzjoIl/XuqeZeItXBweV
G87vAsiN+4LdrnkIv7+7nsNoJwug5WrHlEoIwQwBi1YqSJxs3r5uK1qQlKnfg5Ct
+bF750ixKce2TKO0bfDlO2+cfuOmjoxXzfeLNfF0p6ze1X8Eni+vkcqLXd76zFVk
ZihKH2gey3cqrkxPKohzwdntNp9ssmU2OEeX0svpDGTFKJGYR4RMnesEoUDnvhgY
QIzs9eFpkTEpYBnVakHyxewE+41Rmuv7bxennw0C8vIG804oDUdV+m/podTtnYco
FdWBG34cZGjYpXBoobN2Pyn+5NRzv+0jXFM2oBd+I1ALgc0cDUCaRXgI1rglYeGE
DdO+8Hxqm9EviRu8zXm82GZpbPbARQv+KoU3Eiru7LVZaGEiJOMAMEfNkpDgNO31
PbHJoVtgSqg1+rRwcnIcp0GCGFNCNT9rq9n0RPMqPYIdHCSO4WgQ7XNsIA9f4rft
DXOhGbWtS749AoAm2nULBggITG8D6a58X0Qgxae0RhXJPDCvKGUpkL+yPi2H3+WK
cleRAVVM5/YYW4m798IB1+5lXWVcKvwRDqhVUxpzNmnNLm69LC9qk9tjY+hqZaXR
wzJYq/GJYpTj141PgPoOWvn+TWj88DbQDVpRS6K2Nf8udyXcyr7nBmKEAiySiPHA
4Id5wRSOJUSikmA10aMi1iYgChcY6Jb8lE9C89AOiU45JKU2ktweqFPyqP03LzPO
OFbI0HLjPGIykeWFmbAmTFBSY0Hm9UjqLT8q+lbbghYAIr8ySVjxfrJ2iatpyi16
L60VQ97V3owW09CK6XRDI0HeD7PKm0pYCRgaWXaHdXWTfqUN8+iRy5pZg051RAki
MyJW6rgKWwmF/aIWV+WU2y3kOVs9h6Ao4x25yUFU586sD5FETyfKyP6Y/+e0rJaQ
v7XlsPyv1HffSgXAymsAwZB9FHCNQfnq4xYQ7D5++kAYmqopjBFmGIn5W33sqShg
NYJZ/l0eGOdlGNvt1M5IRdt5aP7WZ8tMtd6aFGdOGgTmGhDATWM48HbwnF5uvYDQ
RdsEepVtWDixjcM/Q0oP8JIY43Bcr8g9vAiBskVNL0RVEnBb4ffH+SuX4tvMDVsJ
tASaZbw41E09MogVqpqHc5Zhwu3YTy5GgkpVUnboFbJ2NqorwBLe7aym+pllVT0U
oqlSZoCJ6mHBMI6QtYw7OtYU1IHxFTs0+UwQ8zi3Q5iG7UmaaBNUoH/3+k9dzhTX
cx4HIxY7aMcjnjqicivD9dB0gScZynt1I98f/tVBtE3ZY7IUVkdA+sY4k5L9CV81
z+SyivXSzrydc7gBHuvEBFsXgr7j0uDrEoafUOI5rDDe9b5Cm8ekPDx8rSPJH2C5
Q5TBMbb4qieJAgTAAskoXDoVC8ga6EAOys5SaBcbML8DzZsXV4mML/VY3QwD+uad
ZYEeBb8mu1irLhu0a4I7cSBtsqtrNBV4dzGm3/NMuzsZFGNEqTEnO32t9632DGC8
nW8g4wo4wTa/bdZsxkCL3ID+a+3ejfftkIhJI3Lf4IO2BqrWSwJumVS/7c7uQ+sM
OIntF0IVd9roAbK+txkykKZy5KzapiLJ3HjuaXRK+Rt1jOO5FoI7Qk3YcVHwualL
8z9GzzndDv6BdnnM/C3E2KuYWsvd0D05gTvaxKsijLvAAAhFij+6kSVj2MVj7nij
C05CJqHouEUm4Mm87MCc2EpBCXsk7F9ExquUmAp5WHGKHsVCoHZRttdvDsaAH1hr
6xkoT5smWtI4om5/kuva0KDfuJBOG2YghFXiFaMg4oVhoejCrQcxgE31Y1dHiD+8
O/h9VmiW9krxQr32OEbvFbGQZYfYRI7sfAIqCj0oGlMy/Pr+ZIaH3/OJTP9MHUjs
4Lh65F6V80Lh3ZsyldZBRCY+/u8q+ZtxjY8Zid9YDrm+gcWlI82jYYnoi3aUy1m+
7HPTxOH4cHBaMoA2mNleiIXWT2Wzg9paNpIXh2rvW7gI3NtZTC2kPM8VDC6TgDSj
IpG6YPoj1NV5LxemC0Xxs6kicI2YicHSetTJkSN7S3FuQ35z+uB2kQ+BBe2MmlPB
fusG9KALJji/aw1wBHNEvBMb0D5WsSgEmeTWfDEdUQdwkjyDZF6BYqRtKi8lzEC6
V7Q6tmV0QcoQkLodnk038Z7b6l06ZpQW76ICpPh8Wkv1FV6TOGXkMQaEAjhZvUao
nL6sEAFwPnG2XezUHigssM5OBnkjdAqKhUSVMXqDPwZ7UePF3fI00Z1B4J6yew6D
DB9OyhXMO57TZdVLYtmGFZjQvXdoOwvQqByvpnEsUHmVl2rCaGgxzzCWEaBj8n5s
tnxooH18qV7p0R7pfAR/6nrINl+VylgrSDoXZYKcBXakXU9yeQFglLXPeT6uWd7o
OWdWmn3EvbgNeB9e3QWNqVPDNeZ2AUzWVJkY5bU/d6a2Lqjy6LeTBk74nJ6j6IsD
M7h3uqdR+DSR6FhFtzytgnvEHe5WaJkq402Bf4pk0nhKj1b7Kw/+/d1xgfBpxoRm
sLlrcaGZcLsi9c8haHMVPMerBw4PAUpBP7vS5zU2jOjVs05Of9rt26EhM2P39gIP
ovsbjJbzZlmzM9w+eb4lnhENWFxEG1A26yVKWjXkYC4OcGcrDcsNYEwo3Yi+e3zC
C3TfWFh80RyyRjsPjO+4SQdrBqeqFz1gLHaw8EhPn+XHgapspUYerHWJEZGjdBD9
03FBesLXAk6rH+eg7uUm6WkAO+DwCxFdzJgK4srBWf4HQUJcBr6RziBJZCyMGlgj
5UsUnOMSv2mU4bETipTnTWwuqQ328YLtR3+UlWdW/JU1GclOL3PUMb3VjGVM/NHO
OQfTCWBzHJEJvlTpre/wBx5Dw5HCpwqy3WTa1ozsVmV41fGxnpvWdyp6ALiXRMtb
C60Jg9eb8iHFi1w/Zpz+geMHCiS+tdeofx8H745zgOSmONAvPcwzM42YIe2MBVXp
4B22vcqaFD9taWGYwWyyDsx6ak715P4GU6gBvMSXFCwrakQYqD0TyR8JLOhYiF1h
W4hwnsR/JNJK5WA1dfCv28tyJOY0+EPcoYoPb91LGEVq9P0f2xClv048TnH2n9CX
4G63anmC9p2oSveMQm5dJyLO7y5r55SXW/1o6yldpE4Px4Kuw4565vfYrWgbVU7t
bcBsFglrFC0rDEO07RTKHChgUu5bOZAdLuPouwqp4DLKqc8UJb0QWZ7hckTIuJNS
ZBodSrixHXAaYRzCCYKrPMN0HUNfjZAqOi0SZhZb/XETYbIHHGMcdQdCVU5hMDY9
O2YMUVfRt3wHh5o9tHHENFwhsW9pDdASatanTUZvVy4MXJNavpsWQr2E90l3sdhM
6o+92nEpqHLh7Ui4zqbCn62J30+jyYTu+zCamvKBUsyyRaK4+st2GeumP8ecQrRa
SrguFw/AWHQwjVHBiX7qA7IRgaD/HAKjkNrf/5cxj+I1c/8DTeig9uEgINtCeqsu
kmJ3rm7BY0gQfBEfySEWVO0XNM3TJPRfIAggonJ8sHFG9srFLfJ2J4KovYznAqDk
Yx/OIQPh6Kjwl8C7QS5sGgG4bmA51/j926OWWvaPDxQwVYwVt/3VFdMXzZOlHS5I
9ZgXcDdg8OpPfEVnXJzjjgZUX0jahc1FFEI4dHipjNPyhjKQP8WEVk8RUfZ2qwCk
GEJzkXhZfFne2zoS0wCVXMt9KLTjLkpP2pOW9AoyBtRRgQC/14rOGmavnNBbSfWY
crSCAM7uJDD5KsYXFYJLUYS+5ir9GI8xb9SQ0FevuGajEUoBT9TxES1BBPxWiDdK
pQe5h7/ICRm9ERVA5eBsDQtuFW3/ljjZ/cRF7dbJpmmCpCs3vaOlfoAGnZm2T+YS
F+IO5Agu0QZLdA0MTmt54TLR3ZkVHGX743VSiRHrsu8R6qDwq+Wdh2Waj1bY0/G7
UMQ2zpUUqGUCB1XoiAxCEiePe09DI/z0BF9CdEfeHadDaeF4g6ustfVZYw1ny/sR
OzoGTP24EvOQ+HUfhvUYGyw1Qe2Pyc+bHoQCvc5B7TZOi3wqVYCmh+NWqxCw+nQq
85z5MMAjBvrXVRgsHNB2uLv9wiEIaSoWfsasOEaji8tUsul/qb1Ux1ZsNNRmhaQy
rDuXYn4hjcR7JFToLuXvxJ/j6KI6jas6Zy5Im2HXJ3JBskrc4cBaCm2JGak8JFpo
U2FK1a/3VQjve5bwn5hWFS2lnJx9CR9dFb2bD/4qPqRKJB6I+vpQGcji6DviDtRg
ntFKHPMu0/TBeBnXO3I0Y7sOyf/CtcB2UZk6CyyB42bHsHjZAspR+RzzNNvxBszT
XRq9wnV3zlEPp32yn5NMC2AZ55J2Jwy7HoOj2axwEQbLgn5DuVzRTz2/EwwyOSxB
x8R4KjiitNEQDHHr7/eN8G5GQ2aElENrI3mc3W/WXPQQGZ/50+ZM+lpMsZmkjCrc
PgovovuzxQP++Th+Az88n19wfDWODfgJ2P37uWCpkXU6Q+5wB8bPAnbKAw87yfNF
UALAFJ0f5ZJnK2MdDy4jFlNBozbUvxTCJ4x+VvtJN6GNKq+9EbYSF869Ikt9VD4q
Jbz4byyzwB2OduLq/1MN929j2Tw19waqXe6CPSTolL3QpwoN45VHFKj1BO/eqjpx
j/7z9W40/0FQFkpoCrGfS1VEdLpbOCWW9b2FBeaszNq5jwYBwskFiXuPAb6WplOJ
xMpRbkSmPXZek2taU5FfUoXoCtvEz4J+Z/YIxkeHy+c7pFZlULShQLxtO6aSjZrX
bnPeJwEzlmgGstgSxOXO4XOfO8aZSyn4g1nCv/NI5NOh0twq84f50FiYQdGQb/Zv
UVnMzqWcLUSVVek16NuZpk20TZbIaGJ00eILOoZ9Tbu3w9QImZ00E3fKhx5LOJV4
O/t63ATXUr550tFj9EAodTgpfNuu60qKAgLgfuzs7cQ7hcqIwotTzGIyuxw1Jo9U
ZylONPX854nX+hCbzlHrjIoL8VHTXrgURCUkm7+rbgxtSTQWSHHLE4mjIRUR9tgE
RxUclM2ttQF89YbfYCL+jKvLh8jQRbIG5LkDxSczogL5THZW1etQMYJ3fZeWRdVB
w0fs5CzOjU1KiYwU1PqlpHgyq9z4E/T6eqASRTSL26CaYMvTBOFQR30vxA9f4f0F
U2De28mkriIhGscrFk+La3py7x73yxWfuAude2a4G4qPn9/LhTYj0bL2ntROdWLA
WvmFlYKhctMcS/Q8JxSoPInHJM+WEvG2JL1NaES89OtzY9TSibpbcOJj5WAercYU
G99gZeOQiFgwkVsf6qVXMGjWmkd9g0UpcR25eepwTz0EdXaqPrsXWzGlBQttYqD7
zRfpNGtD2+inb9pVtJihT0SvuhDeb6Q1hCRzn5nuob0hlADo9Q+eYMVs+h1sI0MM
Rn4F6VGbMrgHSZF40yuY8yo00v1BPATTBK2+N+BufMRyRjQvT7w5zBh3onfHgXrR
YPIGvZaEz6j/YhotkX6gQB5oDrA2VtwVgoL+5SeJqvFVrk0zoRaTEVoLKB820kVA
d9Kvj132P7KBb+GaG0Al1Bq9Utduj1M8BBay6t7ksTmyy2kCArgt5EP5UpsnAjgU
VuzTEy2h2mThT6p/oM9aDMqjYJCkJiu2HOB4Q4H07b+LPGuazlkgHCka51R0p6Do
E8VScdl9IMQ3jmS8xaRRIAQNUv7DXkANHBOx0oK3H0TuYEwgbbsEzKgBDEnTKc5i
BSGMwq4DfKEchIfoRpNjS+dEdm4i2B7XS33fwFg2aXSXW54yRLxNviddMTIoCGq7
W2pZjHv2EtirupMLx1x5YLxiOvHQvyjVTRuO6A5b6swKy6mkgEygXElfId8/1QBj
6hrG+P1Skdh9EqXE34RE53+Hq4m/e+RyROywUumUBWiLp8+8fGVLX9rVC/6UvkHw
Nfqok8H775e6mCqNGP85W/K+Rus5+OE9ynE6j0Vqh7KRIQWpwHlxNSTHRlM/1QlY
yrAbdtz0PGUic6m6fdKf4cWQpTBeZ+OJhlJeeWSY1ZtPNXDQjY9TqR2APbmLzmN2
Gh5XD+KhYkmYMCtxvfsDLZHdhDxkb53PmRJw2mP+2lSt2NTJVgubO8SaEUWupzn6
9ifMiZ78LB91+GXwv+waPzNb/B1gP54jOKMJ9k+IeoRBG2sHeytWc5w1Horw28bY
CXqZVuUZDbIvZgRuRaCKEcnGkx4GqVLKqecuy1qpzJ9FnC3nVCTwNr6usBc2rhL/
ylEeV0KvfT8ARs7eDL/YDv70mcXzHZBynp7GA/gt0GceAI91gxaM7QEH7r3LhfmW
pYL/SlW/yGhm911cToRE9y3c/bn8mAVvHuQnG7ep9O8RR4F5osFK1iPZeRvZCVVg
pyBXF8DGAfbkKDkHRkH6bfGP78R30Y/8K8FJUZlhCOVqlD4HYCFylJd0LFWP1usG
esWSz6wmaWq622Fh6xsI2cVMjTD7OQrYpZzHtmCMlGnMb9s+gPxKfYsShH/sSM3j
uSaEAWI1H5/5o0nQylD+V4Ds2VMeFVA5YmlTJEtuCi+JpoLR3v00CmkyOm1fMd+u
JoviNdTTncjafyLItsdy+4bz2rTuPecxEjQwuV8s+Zf8bO+ddE7Z6JoP602qiQPu
GF+hqJVaKI/WLrUBOdRySqxcDeAlkq+Bd2ZLvCyTS7yjmF+oaAFkY0gOJtrzC1fQ
3759L8Vll/pRvAFMhwymHh8txnoTL60siTsdc4PtVoff1ja09uTTaQLk5rWo/Fh2
/I0d3VN+mjvTR9FwXztPM4EOrvC2yLJt9nVc5wchMYVTUmeqG8DGLWT1FCMlVuyp
/m8WSnspgDnRYf2BMIFCJcwQzdtleaEDjBM4jdwQNXpeMeAvQSj3D2ud+h0mY8Sf
jKDghOuw7lv7XTRh6eX26WAvjx5P48SQeQVchAe57u2TkRXCswJuLKbkEHRe6GT1
ywbDz9MDz8fP4psjDnj8+xNvzqESJQ5/U0VDevs2mIZZpV52UbGtkrf8QUeP6RGR
1+e4JKlI2TrKFgmKdynd+7FTriX8Dm4YIrEO+CuWRUNN0lJCWyp20pBQDcqQrAlo
3yC86AIbSWneJFoVNlmQH3wDpJzlNww1d/pNMyptgohLqE9KQXKE0IyaldFmBBpZ
skpwMF42AsuMMNV4/4tS9LX+bJRYjGLwGQmrTAgHPCeM87bqkyyzW+kOk6gkqVti
NctH6/+uy/YXCNuta7Y/9hz/gPPKXcvc6T3krld+MsFLDB3L2djBVb217PPRaTX/
uRmWxsa+eAswf06dsH5nrMCxit785vMl8Rc8WPVZWEKC1JTD4MD82fHJC2orHtKR
fY1/QB3iHvWUBsOVS6XcG2Y74bAXmXdEZ6/bgGkDw218dl+NIenP2X1wXlUQ9iq0
1uZOVGy2gc9cTwwA+qhuYO7Tt8GxT0fFtOLyy3GbXBYboia5QqBPR2RlGNfNJ2DD
EomOo4KtqjU6caab96FHxCvAkgYFCu/snPrtmXNS9kKJFEFC2+s2m5bZJ2seNDgz
F9eT/JvYo/n/B7pqKTwLFrer+oQqKs8WFUXDkDr2LA2a8C7QOhzePHb9VELdrFLe
jPDZ54JOGXOqxj9XWKVhVconqKAgsLNON0aorbmiMH4CPT7xiMITMQpFoqh+GyCI
MxjgpP78tWtfmF/XtawL9ZBxHi9OoLYiGcwm37N+CcV5duUFWyEsnXoZhxuYlkwg
C2N9vp3JtBx1dhC/UaRLeHv5nzeVTXwS7HSb3risbWr0CkNaJPzC6gKVbh3wknPS
OyE8/7MOuTfA1LC7RcrtT8N2tB0qvdTI/EnP/kOW9+9xcQPsmoBWwd371L4njN4f
/+yISZicEKxhXXWFVHRQvZb4Q+NcWFczwyvw1Ah1rVULcO3exHiaQncpwk0zDJkM
TndU9MIx9sWNJtKAoiFDQHHh4LkPgK5dfUQw+mEWSxquCnQIS7Km9C8GhaKkaClX
P7GQfAVSN33QgGCm2hQ1gaFvA82t3Mo8UoP0MuLCVxNyu+bCNxwQ76c3oE+EQt8a
+P8hvcAbU48YbA4/1rbjWSEvnMt2+Swnqf1GdCUwNNjhHulUND8dvEwwBmfEqN39
4HEmgolubAoGxD7K/kifHG8i9S55ehMqSfOli1qarePrR7QS3Ws72CTR2IEoH1Ma
cb88gmaeVKxMwOG0LeCFqsUR03rMGAr3mn4hvRHQfnISonegMnLTtWi47d7JKhUW
CLL5Meyo4+r+K00AhLyivzQq0ew5HuSbdq9UPEscJgSxYPLOaAogo3dOU2j8tTyt
lVY4dV9ZV7LTbwqVJwFTm6tQMyfREg5C2VZP6GKDBsybNv6tlkgJlHHv7T8+4Ybq
C4grE/wh7WrW6u/8x3wHB8Bsvvu/TFRkLoBfK/QL8JF6fKs98dF1eHIb3Qlvvxog
EeyMlaMssv4xggEf0J4OZLBs2Y5lFa+bNnlWcubDOuByOWpDbsyvazqPGYBDuQRF
aaUwQULyGbJNOcXmX5w+3Y2XEURWD7eWu9UN0QQUqHNwtvYmdGIO0HQiNo0Bfu4v
lwRWYJpoFoKZGzgifBvYkxo65RIt04iS/Rq7vfB3aodkb2hSO8oUA2QCBNy90+2O
O71Ol5V/5f6EavmQIddLXpSjlUmORB5OCkDkTIdkZ9g0ormI7TbGYEcT7KZOSgwR
uYYSliJOqNjmRFAFVAiMjLwy5YaTWJaypxgbFWrBDTCG7K4y8D+6dEPaVJcKvivH
h2E4OU/OuhMX+lLe4ljYAI/9XpMI1YqvdVozrGWQWk1XI96d0EsEP2Nd77bg8BLl
DlgE8jyfgdFi6Iy0fsajibLkXCdH+jnKBLmYH3cz95KExbtxe1hP9B2Ktcdlc5V7
727c/u0czzhU8Izw89C6ZjnKlvPjxsSnc8iAxlehzl5FUpXMJVmfgc+sXBqdzli0
CEzxSXv7EJgeGWwlXUnd5ssVJQwNxo42f55ffpU+Mil8j8rek1JgJyexPfOjqDDF
w5YlYFo9zDDhgFsswaFHWdiV/UAdHgaJhFNslkjgHXPreNR6K8FhzL0pMS8KpJxb
rWoQhQZo4FVQI4yXKYeOGLEJpVBs9THN3mSe/Fzfuvxy3UcRucrhmSYLpKuFc4KB
sNUvKRjbRJep8Vnv/PKDX0pGt/HQspyYdnwVT6J9pj3L4+iSAYm+y05tTBumcyvY
z6h9z5p8maC1Rad/VEeLtfmvEFl4YnBzNWL7M+b1MbEtGPJst8TsxvVlMa825K3H
kUO+w7uh3RQiQUT7C1X36hfgFZH8PHLgNBxRiP9rUlhj5eWzCEQfm8R51wApUQq7
EpWNkQkXr5i9w3/E31zbHwhm1yMn7DkpWKpz3EPuJePgFhudOoRMYtB9ZyO+xZVo
47JiDNC0EYKoaUacuIfOHkwSizse/2+T5PVCWaZwAq5mhTxDUnfmbmGbWbf2wvRj
BeI3akBAepdNIUnP73p7gGbZlVL+N7Fp2sE7Qmi0M7aKhpFa3lyigaNh3GVzwcme
H8CIyJUsrJ7tSP5sA0qTyBkueV2AxoZNQJl8ngAh7lrKeEGBjWtOQ0kqJ2wXlnJH
pcOBDkr/LBWf8vpSEyfqzTJuaKxSc6Bv/Cd3v5xO4fB5pAwUWEsraIrlrSlfMEJJ
w7+qseRaWTVzyMsgtc3ajHPw3eCm+q+d67H84V0f7ggzn9EeX8hRnVvRxUKbRyBx
oyQK8Nyr9ANvfXoMKVCWogVfbtcG20mqTmW7sey5SrkDxA+JJ1a4BV9PlTTZAZnx
p67ox5gXr9UCPbdGrywPmGknPfJoPPB0R+P+gHMJhyNyIe/iS54nZXAXYWwEMPan
JLpkmxhmbZOQJp5EPjzSmahyHsvMKHqWp0emlhh/06hLCX2PPlxyEnXFUpJWDNdt
2zwIZGzrY+mlb7WO6wvOd2IxTMn+Xv3UEZybIKg6Q5Fv10GVfowD2j8nQllb8m2q
ri0NCY8AhIRZkKyGfJNX1/HNJwi2V7TMy3KPzmGDuwKUO8he04mFmYj6d0BdSotn
cy0PAUfZZistIyUgOSt1hTmS/YCzKLh3CoD07oftV6HorpoKlmyzMuqETz/3ROJh
UGQL6flQJGpEXG6BZPYrqD5AEgd36FD9zL0hHvIn1nK5e4fTLmcYYZZSgRxV875q
KaGWhgT7fgZz5xbd8QmM03DgHsQuhmW661QIEnBeCjveSTV4et7zhnUx/giL4KSF
BW2YIzAwuJIaUNdT5DsOh9mqK2EdAUuFSR8BUqioFyTYvCFFwZl0An8vITltH34U
irdAQeGU7kl0XTqj1cm5W5nmdueYLOLngq/zlQR+GEyz9Ukw9LS8AoH8rRN6HhC+
2/80NyWTCkCuZ5L0q9WvktdtiCsQu+BaT71X4FNgiBD0caNlfZDE1PO7PCx3pZv5
bVFitAEpMzeTVp59sClXwF8XoA0J8z6BbkmcUs1v55fXaT1ECgT2gu5Xl7poYqR5
7V5SxGr0+majHyF3L0k3UkQIPCS2Ox5ta1r2Oy0E1AnjU31obczBUcMYTzMIAQ34
z+RqmhplakXAlNZLGXu6L/H9P8JPLCCUW6DFesb3noFjkViCv150WmQdogMSS84l
ePx/D666LJTsi3QumyKEp/WdvQKp9jTw14A+DkBTwLXQX0rn9SaXPhW68aB3MRSd
SoJJ8IYteUM0LSv3vE/is+RC6twbK9bHoCvvps35N2YrpRMue+XRzZ0vive88OdT
+q585LxvW7oErpNHiCAj8KSwLFSOnKWOXJMbkSyuSW+wYKtMY/PQoiwC7QS6XsPH
/Rnk8lqujXCq0OHIzMKlKbQGhtD/iqZ3i6xyDEaNTVm27j1mbq95GnC9yhF2OPCB
ESmLNVGQS8vi0NSq0yJLY99LfZ57XcQOm6F9IgERr/GnhcAT7Es575xkg8Ej3NxX
abygw1IytKMLxn5arj0ELdgbnF8gNdUQj0h32nbW2kkCBwv1Uk27iB8DvQjVNftc
x1h6JKCG1W4cWStfU1ME4Wi8mVJb3huExKB8FZV3THklg/86rFcCxAwp8xUeCBPV
7GIOaSUrYDoquTg9Zsm+PcbFCR1yjQxvgPEbfRaT8p1Vn1Jt/e+vcREQQLG0oZPC
M2TwyO0HKthjylZtpOtdQas4YPIADdfSUxijFPKTuQx8R3gL3twiHucLn6j7hJ8J
+OjNZUaLrTIfJz/mKQOvOwH24FfCvsXNYpLlEFMj2FOuIUB/Xt/3UjbWm2T964K7
goFPhxJQZN+Kr75GdbXSp1jSm3MZiJai4NGnsF/cEZx3BO+Mq3Zo5XdlmmgCPyov
Wu2DEzzcn06lmfKTHaq7uPEQBwfe0QPvYDjeK087gZTtjG+wLPZ5gvV/1TWjOKfR
txRBaB2xGdB2IAc2eTvNIpDClXRnMer8LZ9hb7imSUwncAQIbmeVlhanFY1ofzsX
2ObL2pW6f93kdSL55wMpqGb0Lmjy8zawj269C6wwZTpKviLn2uG4YlFiJF7vSg2R
WRCvcPPN86Iblq7QLlJn+L9psZjc/baMtKSuP9PIZ7P1qMF0/yQ4lItsBnNyMlCt
WYBuzGnWc0cvsk78tMy38MyiulwcgP7pbitPz9OJCsoBoyMFRWpCTq8ikOsJ645i
KM0mifYituENlugBUwTC49Iv6kTF7pHLuqEMS2i4wpotRbQwjNrLZuwpB/0V7Y7P
pguhrT5Y1u+1hw1u8Kiz36y5QibuY+FapFEg5ywryBzm9Dsv2q7d5Tx3AQiYlCQh
g1TAHty8SiVgui4vOgmUrtdAi1lPYXDpUQNE8sQSAW/AV5CVBuhBnDUz8hw/C6sa
os/b6FoBpLOo2HqkYPxk5uNAPvKyiEAacZM91OJlpeQrpFiyPK8d8wLW6dnX2fNN
qRNh5fYGwz8CL6u/BvGYmdgrIMhTE+f/bt1Jhh2/em2G/Pytj3Wo1eq6Jt4C47gi
h/f3pFP1CVBcBwm/t2m2iFE+9val9Rc2uPctOued7G1INnxUPG5/1xQ1oVzDg3hW
NYl40PDmJmI2oBJ15AOAD790i0OVaq/6cGyYla7+un3Qj5RgWyq7UL5pneHTL7Gk
eFQAvXmQPKDh6NVLMO1/pkzHo71S7IqinEXHP09s9TwJSgtZGPNLIXqMaaX4cJTU
oW3NbO/CyyhXKMc1an4vw0j5/JlulXIL/r6UMXMgpvkVpIXh5BYm7v4SIDOV+vEj
1zbrtO6r17F34DNMqgEVx62KB5vafxYwRkJEas3nSFULPQD60+HKyQqV5gEetDAB
L+HFNaKal1nbmQ0NqtX75pmKfGBXeP2Ls2V48z/O4sXE+waNbrRPDH9alhBGSA+d
CQ5aoTeJry50rxGAe+1eGprSHZ+silRVh8/0JC1mvPCDgoRVj9tTC03oYS1GPCSt
nB3TN3jgyReZ4dR0XzXomenXhgpLtgKgMKYqaxP6ewpvVkUefYxkTq/IqiITjPCF
igoaP5nsTsENbJhgmTRCeaXOmPUbmURWws5SNxSMrLI4d0FgCqnk9zWW3JAmUx1J
H5iSmx7Gug8/b/fKdPwalbhfdCuAJCwoE+pIfC8KvCIZ+9bpNvkYUiV4YeWu56F2
qIGSsx2TBJne1R1KaoGHMz0bWKb1UM2fHcBpNbDpYx80qhu6vlFbH+ztstAKpUxP
jaLcXAyYbVXrbxPzmp8wMnpPkC0aHMxXPHQZDo/UM/eF1NMbtwE9VBR4TV6Pxcbf
nASCXlA9wGr8ZjNJHI5IHWxVD8H+t96WAcZzGOKxJO6G2qJadrikcjdLcfactMjl
3rOf5e0Sz630qCHzsWFRLgGNHsdfVSG3mb0P7Q3FT88afaV6AghDfDrGmS6Oc+Ye
QaxJstdzhN1ehDPRmIE3x2Ch5kI5zieBCGpR6eO/wZYyx37FhmliZqn6vgcoLuEq
2ta0Gqkw42eqWP0kJK09bX1zNFi/ZexQZhkh79cvpDrSiIWzx0GvTEX1rU2l8/ZW
1bfPMxkux5Mv6JxNtqlCVtvg7oUhhTefnYpL3wZZ0i6Gni9E9b0ms7676azcRipw
cqM5GhCIxSD6EaSo15P0UgHD+WBiHJeKX4RrPQ6AFa8KcZqcKBTg5Od15vEtbGqM
98r1nPyWobtgPFwJIAIfCh5h9ynX3OTQCBczkgHMBijSdmeDJHdoZyApiVxfTnwc
51n4uV58CRgzH+Y1+aL08Fa4OMqdp9OxTWw4+JZ1AJpW1ZKUhFEXuBaReWD9ymrX
OvRlCOdIb14V3WY4wB71XIgXbnl303JCZ/rjvufhlXIobQ3hbgjJ3/N4W57JY+GE
FL5hUnwQ/y6y60GkxQenom19powwYpmVD+kD19xELJDvxRIHFQpE2TE+WelRQ88K
`protect END_PROTECTED
