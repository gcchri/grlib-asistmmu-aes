`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3MCrGJIs9Z7jmbV7hL6PoG1u0yD0kAKcMuyWWPdKkKple2S2abC1CJ3IilISO2T
kTWYJZWj+PUlImTzI+PwV7BxInmXOCkW9kR+8HlxGoz2y8ISbyBQDbKSqjoMn8Xd
2Hwb+lviMdDzO7Qu41SIJlHmR7g/mSBP2F0JRyeWoaS8d+UU0yE40vzUhg7xasOL
2qw0xscSD4fh06z9AQ7F7738qtKnZGtit07+PuLCwwmjjo10jzuE5a86hrft3s1F
nvmV0KCsVMtUaRQPbqZdVccsHwRtijBxttW3TcJzpSTTljn3vhTItZbY2dlsIDiL
+6lfceLMilG8XD2R+sWYZ1oGe7k9ZVOLJ8vFCX3gXFlEkXLXt8Mc8aD/TwnjRfj7
2GRL6bkYQztXOAKlnNxw6p9ehAHvfPh5NyHyWZn1R0oB1aFmDuO6v/UtlPwarOXT
Lgu6+QvoZdskrY7cm8tKx8RhFLmU5Vb/f6RQIKsZt/v8opVLaDdUkkHk/jV5lWcJ
TY0/f9LF5a1iTMzv/5LlwAx4am87fgr7JE66IlpaqnCWhHiyPgV0NAQQ8Y2b3QWe
UGhCaw3rYSNXLEL+FSVnbH5NUl3rUXxA6yVkY+x3heYcSRs1sOLR6B+b+xPDAhFs
LREDm3fP7r2BiNAbC8D85ZbSB5D3R7XQn58EzHKXXeg9fI5qof5jfGFamkZ0z+pe
E37ZVagcrZtA1oPGNUv+uKEmAstvzx/CkhRAZWIJ4M458Wt+em3ZO5miaGfn9Nsq
HJd0v8q08YU4i9jY85ssD8/pJqxvkI8Eaff9cI8MKQ1n9P1mR/iaCcZi4lky3YOv
ofshN7k+F48Ga+fo8x69L7Q/OV6sqNVxNazXI8blgOWYOBPwTmibjUPe5XUHKQVG
v0kNuPEnLmYkOOwb5tUjnz72RWTyrZRBvXT03b+NT/J9mCVztZc3CdN/QWXh/Spl
WEDdLVnC62cDeWP6h5/EaMSXSyA+c5vVMH9LiAilDBbqNp1WsnX4qsXnU8c5S0Cv
hF7uPBfk6u0+TG4x4vpdPk1mL/JBI/M+4FRvXXoxv+fA2/6DGXN8rDlQ2KoiOwxj
SJLGR6lo9t6iPLd6hf1RiGMqGhhNJgkt8id3+khqA+nzPyYAGMKhyV2g/NGeKvrQ
uhIpqcaND1Ylg1a31jGXddqHTblAuFZB3IG+WndpxZE6viLlZnqAxOLYWmBmQbcv
DIFZbWOecRxZaLLB5Q8DquxyEyEY44DWnEe1e9JmR6WqwlbQf4dQiYSLACk127aJ
l9bKtcVJ8GrEqLsipINQu09hM0hcmD48Of2bI4dHV7DkHQYg7QmYDWelfn8fVxue
SdrDa6vaXjb4hEdV+piJ9o9gThs5uO3csUv1td5LNzntwWHB7EikONhumj4djSYn
lo3uDPC49TuQ6oaR+XdzcMpOuBehL0i9JhVFzzzF2XqSQqSY2nUcWf7iezAC8s6g
cb7z7pNqI/hsSSRqbtFrnWy7aIqmkOXj+dzvmcraUlNpHU2LHwLudRm32By+EU+N
qD9eqxCL4lkjelaclhadxs4y6Hm+16TgipJXphr8k44iR0IdJLppne9OrCBsUqx+
72/BX79TyMlD65DR4g29FnDEH6q95EOkRJFFoL3qWYkVjzPCERKWZIsyhq8X9y/H
T3hsePwqt5wUjWQQ2LrIWOu3rD+qRkBovl4DASqByjPtUtvR8fZCK0STjZy24USE
ukl39chHml9oRiFOozjabWRRJLP9exRDEQEy+Q1uqskI1Vw1TAkwGCNJtLdtNN6J
RDtohk4gpQ8njMl1DSJ5q8khVGGPN9OzfAS1KGo+/ob1MZXvGvWCVwEwpsEKT3CX
Pj9VCh+m1Efhv1FELUSMBv2813HBBI1HdhEqqOWuOUf+pb6OSJRQlnM6jOrHar9Z
7w01Ci+IKvvGqZ2RAA8X9IPDZkopap/dE4hbfxrMrdLP0i8tUaBQ4bbZurhQ2r5X
a2HnM7eqExsHj3bX8yKagfsokN2MKwv7YGF5VBmfvEMtbJF0GwH4eSxztBFokAEV
eqVBQ75JQjYTGRKhO5M+QoYT9oe0VIggW/JjljfN2Fk28ZXNb6gYmd2Ov9sme2w6
qKz3upe+y3W4yOCURzyVRX+l/oeD7ImECnLhpbyipA56GIZ7FTdHEVvBduhHGoJI
ErZ1iSzKvWODo/7n2Tk8DQF9YkH/L6XNyGhAvEb+uQErcbzEc+YpaA81wWJI3i05
SHEMIJqvUP/Z9mbu5Jk1etjI0VccEvsVCTd1m/KtvfYdPJtwmnKjiu4zKO1hoZpr
W4ZxFN3BpqCNZqWheKV+h3LW3gyrwN/GjMo2D+tqgD4hrsUUxNi6phuWFo0UQhXc
vfgmWRRzZEpLntFwYSOH0vDNMgHFELiJtA4wPn/El1H3h8KlpkDD8O4tO59aTvni
8NAIDlIuEDjNSNDU//xkmEoJP9V1Ufjh5vBwtJL0ttaSOVKvKEEVGPFizRYAXoHW
cFmyjbns2A06G+3gY+Y2Mwde5hoNLp69v/YYl3uIqkLjNfBZ1UJrgQk7j4BoFxl6
C7c5SwACW5qRorB5ECxfIyWMPnQUlmTqW04/586lQZXiTwKGbo2yW+6jox+rsNfW
JOGyAYeEhmyq0XsO9HhlMD7+u5jfm1ZChFGPqq74iW8TQlFbqb1ia0MTdNmlvbeb
JdzGoJNmYr8V/qvql1UShNJZjx6rISVx+CGIwlWYAByIaBrz/rEus29QjFaTZqQY
LnlTjvJFJtGpq9QQQ+lQJ+dcW4FJm+NQuOlmgV/ospHK7cAZUJ9HVR9V9bR/4rLJ
sWFK1gCWZOPtGD/5AiEsf4OfIDuwHDTFx5Es1LwV5EsP9CpEEw8jCJwFe0A4bKF9
9IEvKktm13sjxbRBc3s0vRfoh0cG0/tcI0jwZD47BPI4NTB9AOPzZDSRRGzAh3hA
Yjo6MbZ/8gj9BAQXh55DfkgskuxgsKL03e60n5l9eouj2TwqCQr1y/M+hsxIuIiq
5Hs//7u3vbidspTaaeMx8WRvWOpoUjXGAbPjXsn8cgjPATIn8qpyPAgegLefk+l1
6Az3R97lQfQ9hVyzeyGK5AnsH9yeJ0cyTn6opUOZeSqbzArUn18vgZhWuLht8Hq2
6aN9sxvkIpjC6zqg5pLgmamcoTByYLbXuIktS58DmuszHYLG0ixgXM+1JhNoudjv
R1Isp92PlWkh/OP8KChodEPSRD2PKHKPyigUp/O4fm/XyXQihVaUwCv4uYg0phcN
ysI6IYXA8TIDKqGTgqPw4CO7rNIHhosN5dYom/g2Bp8CQ8uLICnjTpf0KgeQfqp9
Niq2fxwqurSEZh8+h6nrDy3XhMraBkU25KYxT1Xxc1iuHJe5KkRkJPqSYL/kgb2r
scSLQkafyCuFvjuHyZQGzacSLN6CJGSq0Cqq2UbO2zyJXKUas/gGSJt6oVZ4hDdx
n2KpiW8HYPw3kNxDaF3So3cfoi4J0iUQYH1IsByK2v9+2VXx+a4BBXGXaqRStg/8
RYOOsSdunCv0sDa5OMoU3N0uDp6RfXBhMQgQs8w8U6g6XY3pMbYc92Jx7IqequhA
L2fil0J1W+rVgwhAZej3TTO2jnlEN12QsV5xI3xl9wUuuTkmSxP3t4wQI0QETrf6
yV/vgZ3orPynpVE/8GXRQbF7rHv8fMtP4cisCSxX6D7CnQT7vrR8NaWscxs0n4gQ
cuH2n+coiT4CJ0x2M3mdn6UylZsDFGm5zpBP5StP+Z/XT5rptDzdOl3Brf1XP2/l
02Nli3YVQ7APLZgtoCNuWT0uiYgJ9pgDgjQtOA4wDF8pL7wx3/qWVafEK1JhBR3i
KAytb+xxd7KHupKP4TIYFCgClQd+h2qhCeKLbOiJ1fKJuPuA1VANeNgsBR/vp8eH
9i9NM3cg95nstKsnVMnWHWHXdWHzyFPP0/zZPik+RsthEiFiGt10nj229YrzDiIc
f+pg5He+p3zgSmYH3eNcYVHmizG3r0MVuOXaQEOygAy8ZyGsjP1CLhcXeig89x4w
+etWpxlqUByahiK6j9jMnCLucmVEdQLEvt+SDQdGyRXZOAMeDmXV0mDtw9vvm7TR
KbRG1MjomEiM1wb9hVrHf0W4hh1KpQ21SbAGg1ziv/1vNGDSaX7MzEoA8KMM4ORi
wPcG/Bl43wop7SiovCfbC9jJHx9/tK6Pmj70Tp1mlNgzF/wTPuFk2Ze0zTgFJE1G
9THSkqXvlCzXPnJ3Poygsr19Kcph33pTMvHoCou8RauZY2IFYZnjctNYnmjelH4J
VYA7Xhmpjd+TEdc/gVk1ZpRQEN+fVGmhrPTCabH2akDtZWFn7V0QzIUN3oAcYRE6
FaG7a1Y3/1nqGwRpEPH8Ns7UNFmYQG7Ckn27/qZ86i+TRcUhnVgtZd61fQOsfzs2
Z10WthtF3WODUdsp+JKLPKbAyVM1FwB7qYM3I0g5AAMGYiO/CJH8xQHM88Q3ONGV
HK1/NBay0Wm+e4c7KHSUQ+wZWxBjGPkF419ZJBqsnuLfQ4l6IqMENhmNqR7Lbjcq
y1H1z6Nv8QfW8IL+nrU1EitGCCu8PxBFZTQRogY+LecgWuKPWk5E93+vFNt2sD7u
0S9ejL3RAucg+BSYpnV0j/q4guj7HH10a68xL2MVFGPCk8JFMsWMTw4I7kZjTb2e
crkH+oDZQxT0rHXoExlpbTTYk6/9Xvb1GHOJeyaelXY1RMQ1GpmCx715hZOr16o4
8M/Xn4C72j5e8gI5pMyR6mTbqOQ+/hI/JXRnbrEth6iV86xufzZX3bxDpWt1KS0q
1ns5Yu3f1l4mGcYzTpOtCVUD8q5qvqV8VO6N79lanAnKDhzix23O4RwDz9aDVfoM
eFUdF3MUKBKECF8ESN+V6LUs7WciZUTZl04+x2a+hj7EHM4HLc67P/xIesntsCpZ
2zb1LTg2JmHvOaOvmpIYXZTtsLJOaqVg14FJ/K1jmP43H30AnV7oSnJXPnDEDObC
jXnNNCGpjSMA2jq8b903soptbCsWiHbEYJ4lwvDgZMquadgWGq0cPTmLrPhiCYmU
Z1IEob4za9BMudSUdrjYE4ggUClg9/6u39srzGC6HdLo2nwYmX6MBsPr0OW6qr71
zfY0vdlqA6O2mFnfKyf3Y5gT2S/W42eQzAfN7BiAQbhVitkkGJ7TtZ4W7CbxL11t
UON92B7i8p/GAopjXD2z/RBwcN813SL2tHFYWJYPSaFJZFI53jybYhiUgSLA8pXP
uRd9zFTv0s+4wfratrgQNvZvPGVMn1xsAegKh37rZ767XgPWTho2/iQF/I5NO2bF
GdtTIUWwNJBeuUc4p6h1TmSLplor1J9UVOkymtrBiZD5Oo9y4ePDTh+fre92n07B
pf4E7ad98PoMXrs8dzgKA8xiPnnC2hJo4R3zyZJ+vTU7kqR1Td707Vl2m5wpfT+t
8Td4mJRNb+v7nDuTvNEC13bDoGzQwzqGsqEImOb52w7v5C791T/Q+mQ5qQTBf9vV
7caSNR8AFKy5W4qyaR6q157UarNcZkKGSbjLHjj9WUDWQ29e8Htyr7zzebbCxn4j
ypT5Zcp6IygRgoyQgF0G4fbMaGyJ/LCB+LNXpOaWz5UaplitkVKWWjzCGTDOIDy1
vGvAVdG0saRRUmj4IdeW9D4sfjdMXk7y9IU6Dctf6tIWTU4fRbKP308xTiBWRRqU
vDgmRcyWEvHPcDi0rawVioT6QtAKNvPrzCtf/01dTQdNMr7Bh6xxKIZ6BvafExhb
sxLEPcrn3FJxf3nRMYgCcJbZh+8OVJQQp3hMLbCDeCAvU2+9k4lHbUrwdUGFymYF
Uq++4kCOpMjNDho+ImmR9AQo8U9aqM4Lkpt+51/PaTuTdkZSu4vHxjcwH2fZXyPn
RkVtA7luaFr5k2Dx/hYKD/awJyY7xD4gm+uOen/nLUTMIN3eazH0wOF/5H1tOpVX
BrJcmJvxaddwHQDD6+Kn+t1v7bSqXD1r7VsOgBdDKd0mTQS8JzJFV9GhdkbkK1kq
C+LjGvkj2R6VjsiDbdjU8h90JT3lIwe3KIT9Ps9O+XBsnaQIEqjgUTVfC9YayGE7
dWLEPnLprScP/4J/eSC2MsBGj1BETO2LhGqky/FqAYjZQCZGu8pztxekXTjam4Rp
3TIBHZdIyHXH/5zSYImx/009igtv8As8vjUbjlJE+ufkaL/A7h6aTB5EhXESdo/v
8Ug9hi6AN345FXif931f0HZlsqwOFzC4Rt+YI/VfQdDsE44m9LT77A8jBWRGWsdT
cAKhZQ/S0ZSQ35xu4zQRNxHUBqEIjhYVa6qULE3AqqePzBjtQnvbEQ8fx99EabOL
T/U3nJHd/qy3BE/fWSnbFgWmQnHiRzjk1acmE55JfMH8R6ga8n1H0Tk0Ts13vK8V
99NDEAMraB7x10BPzEDD36nSEWyAkaSz0WVmxWgmOmf10kJKSWyICKhmwvIkH5uz
En5JpdMkiceMt48xTT36B3uBznv7ngwBntMJBoLXxWZTbXgF9226ghTtW7C1LVK1
dI/+XtsuwBUm850s941Es+yyztI4n3QSPYWFqkd6/CoiCT8L0y/brE9Y84fT4Qyl
AkC6JRrEm3fiuwPQ2e/hX1Ii3lau9uFpHKaPov66q5WI8BkncVxYGuJMDcKjdG1D
5fbpP4ZdUkd7sEGsNTDeYLvoJiFZxB/AcAy+nNfgqyl5Ppyqvvq++rIeFNwHRRc5
t2TteQwFLqwmmxDRpG2JkRStgupViKFx+fN6N+53cLzqovoNtx58E/PVyXi88+mZ
KaNfO95pCTfA1A/xWvyhp4GSr8C+gdAbonNLRnNH7zl1CjsuA9BJFzrZbp+cZIZy
/oGM/3VUDKTuJIxSjGW5bHMAWx8LdBwLwBNSeS7j+HQCaChBmIQNZkxxM37uKtX6
i+FDe844lE4sZT2+g8Vk+LrFzoLCxgkvFTOBz+JK2D4zXjDrq3b16BPKSIdE4p/c
Qbk1nUP+RG4F4qfDRItD1l4c9feqRDTJI8nizd0WyX+Hrqs7mlFbixV4Axax9sM1
S2S+Pe9WdRD6lIch524EMHs71WbZxMpfg7meRYndeLpogq3UtjHqYt+NFyxUYZx/
E3XH1gW4zRwVQ8Wh5zV0fSbWvtOBUhUGmXQftV15pS7UkquXZ+c+eOGuJOUPmta2
R1g98voBbnsyreO9iJECkUoTkyYr3M8FTirD6LvhfJkb5UJcKiln3TeZ9h2teRFG
nad5KILFLqNE6AP5sY42FQV3kzL6C9uqbAtUur2yX9y92rXY0D0VA622S3Ozj9/h
IRUUgtcu7wRvtEh3NDE1q0pab+7+v0fTUsGr4npmmJSHL521vmZdjRlipWhB1UgC
uKkl4hm9cBRrV1yUHGQgYB61yo1eHLjkvEr+6uGeq62JAS70pXqs4YtLV2ZZ3k50
twsNQn8tsOSdHJDqAcaptvvhpe4IIsWr3cIXIQf2+FEsjus7pBJnZvWRHwzmKcmd
c5MN82TULgm+NgS70JpjD/G0gdAbPN3qveXcbsNeHl9fK/R6+mhAfkvpCD58DPdt
k5thlKw7yQ/UQZrfUvivgTiDc7hOJTL0EA5S8i85gcprPtGQ/biyQgHmElmZa5Rg
vJUTUlEMp+RQdcyBe4/82nMmfepw0e1RSffHuPUxwJHzQUuaxjjea0B7PJ1HMUHJ
sBNK3k9HYc/ZK/yOzoyxupOmwOtYzAarmcLl6vRjLzCQSO2wwlbk448mnG3hckDm
Sk5rh60FtSGFBogtN8Xf1dg4PXB8ng2Rg1Sgigie4t1PRc/5JmbE+AnmfkxWcPmJ
zugFNxi28M1I4EUErcWP51YSwdv106xneW6Ox6Vx9YH4KF5axBLcFNhLNFWOVpX4
+lmxRjiBV41bn0GovLl/rvm7xyBc8CgZRM+r5yWv66E=
`protect END_PROTECTED
