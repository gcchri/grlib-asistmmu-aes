`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Btw9us7oPYS7Byf74/mVq7NPxu75dCh6rr6HjMsIH2KRMh+KQktiD20hnpIgor4z
dFttMlnkUjW6XnxaZuV2fjdpYM6dZUFIKkE21JLJ1XF9PhAHR3P306Dye0a/2IPv
nwCZa1+Dj2gnH+80aIiJSWewNqjPKukiPxMlDcwWryCiB7qpbnk/meNicZ0pu1+Z
QQPOFs+8JTcOJKA2Qui2UD35eThJwGYxr44R2ZvEmKf6QhNsxJYnXqMVzZ4Hkanl
oDRYd5YFqkJ2AOKxcbGs4G8NIWn8Z8A4GX0bXl+Rz0fsvlM5HeRCCDh/Q5vXkE9y
rvg2u15u0kCzkSAj0UHBIipNFlDOQLjwEA6hPIKHaNrsWxDeDhO/7/7hW6SSgBxj
OipAMdVMzfGBPDiAKlq3ZaMnFTlcFFk24sRJ24gMDdywpGgKK7zNQgHZ6aoEr22x
YfZMqD1D60DhBvhBEZ1kmUgzvOyFrIoGFQITF94XecGmazs1T3YvdSWRDV2UrMiI
CfjIHDj6W/JfYOah4qCK/TStA55bTmkDpj3aoK+8yyWtFOrgIQg3XC7X3jmqaG0J
VxB8a+9JeFV/0jsizEvL4TsGMR39pkxPWVSIq6RpFunyxVeAJxxn8fpjBIyd3X16
jmS4XkAs7ihaLTuPjPCC1GimxNYvvK5D0bjx6yQqemYEB3i0EL6tv6cF6Fvnr8dd
+e09v6y1win3EdtUfxZJQFiFsBoj0ta1+6dYmpQjTq9YuODF+ugvcw1TkjVK3CK/
fV1wiT3OQexWzc9kdpp4wDSPxUu9wuDkO+rqWUq6Ecq0TFeY8pLdTHQJiNMQgRGE
Za20HY0lZU3B4SDmarEu1I/b8E6N1RIwUfleVez4+qFuAD9lUE/JrRRJjfL5xLTJ
bKLOteAE/SIMO9F5bgspbg==
`protect END_PROTECTED
