`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTKpAf+hh0Auma+sOFWtaB/NXBEpdzE3gFRhoa1UkYR8PXKexOjbuKWbhfsRT7et
7OdlDC4E9Rvnc7ijoWgjxoAEfWpEhl51Ui1yNPavgTex3hQUL5d/A+aVo0QtdRT+
6/2tTJv3WFE1CptDQ78cRbma6ndB+OFy22zG3e0GMqaEZYBx/NHwAg1bdcVzxRWF
HPhrU5tJQBFCgr9yGPeNbMvtYJD6RpAl7QgPJIZ2r41aaNNwai9fSreHhvYdHiO+
TuSoM8gYVZEU02Zddjk0bn5wp1jshJrdcYfyfMNylP1+3xXdnBhubZu/EY6WSqvz
QyIT5Ja+Ue/tzR0lV04lhPy1htYOmEj1JHKQv7HyfLZ9RwINf4vmf4xQOIoQmN4I
6ajFZu0cD+B4qnHEkMRr7mPiXNj9B4sMXKAol2mxdP2vhfAgTiEV7g1qAT4qxmWn
0czgcIYtg6y5YBl2qATVRyENfxH4q9rUdtzsrkTlUJKqCNt8VE6fVpjnLB3UXuwV
/zoUpqlHNIpEA+NwC9MtqA==
`protect END_PROTECTED
