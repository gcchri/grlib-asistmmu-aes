`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lvreq51OSN2mZclILk3lck/47Jhc1PU87+Rly+A6IL8OEefdm7TZvfkGMm8ZSEOr
hz/Ztij0r2ci7xAgyqeTbAqFokenkN1DHDvR5cqOHBsOeiaPJQs2wF+2IoquxkdX
9vEzBeiXwezu6uGsKLsXuTKZhJoCF+U1giJI1QZ1qDsW82emAZh5GjQy+9h5CpOR
XSI3Mff6EwyIJQT0NhZlhZ/MMHwD2lNU90kryQcXQIuVfUyHgZ8dqdFBs41qFLQz
EbxSYwAKn/U4Iq+eD9YzU751rg8LVZvu2PaQ+QNvO7CXJ3JCjci233SBTadWEmf2
QVUffM+KnEMht2zZSy/NwbWOyPUNUmPXpwPh3QFO45C0qHKXbEdMgvqeUtmHpkM5
8Id+2DCkaC+yt8w2tC8B5bfroFy5bV323sGRRIfJEJVnimH3hRtxRqda2SqzBp9Q
aWZ2dJpkXZrPRQZnKJ+bRP4TIJQLaEC9CtiC0c18SfEe5+5f8YH8Ru5sMyVwktIg
mP3/eSZV8khEq6oWYgbjhYIry7hKpn+gs5OniFIT3oz0Klj0dBYrVoM541IL9bDj
a9ZYW32Zo9rT5MSbotO8cgv9hET2wSFGO5/MKmloQ7DFxQezgtwbsNDnjP3hwE0N
RPRLzt/w1KvOSJVmU/U2TEQVyJ+5wf6OVwjhdLwOFiPBg+uvl8LoZz9gaHeILrmK
F1tuIy0mgxsLC8GAMa30BTuRp21yt9Z51KpXVXi2MP+Jzl2S/hEJUyDKCTEGBnz4
y7RoBtyU7rIugmCasYLoS94+MiHBjmPL2gB32m8Y6QoJM9h2aMkvsOgNYOAwj7Dg
DyfLjUZWDplKLaqNpiueZg3qdVqBmhwxns/8HNsScxCLKkUCBXjeihxe+Uw/ltz7
u+Q+5nzxZjxs6Z5Oht6Chgp68SqHAVZ95VWhybhBXFZ9+sR0BMyQnQ8AHUWOX7E7
AA8Wvf9rSM5D6RObLzWuxVdl5eYemiVGmTPjiIhhN/DAkhfgFQDqDEPOlNwOe30r
aZupSgV9xzHhLMotAws6uiFFL2MbrDz3Ic7iULADFD+JNnIN+ALzrX30no66xLqe
NZSjtzg+9XpvMcAghe/OtLC9tskkUnb5d9CZyWWCvdEMFsmIxRi2wLcgFQaysKXl
FKjXROrL+EG22iEe3Hrv7Psss0eEintpn2WaDsZe5OgzGQJIBol2w990EwQlORIR
yuCGPhWqu6YM+GHytraDMORqrecfkxZizYmBfAZJssZtcaKAUmmlQ7YN3SLAbml2
NZX+nd3re94SAmyccuLrNoAqFKw8+1Fdvun/LfxiMGSL/KRTAGwIHnvjSWWc9KBQ
6J5To2MbRR+7v00cf87cpC4Kmcz94HFySZIKlCrSB0UeQEUmhkcFdeA28GrmLMUy
51QCVgNRjJThABNQwFLlVkMIsjtWWnDHJtQ6+ZEf9rxZ7CLQpr3+QOUntybZpsbO
DZUPLu8RcE7XXTYT+BAUAmgBcjhlBmVTnfrIXZvN5yVGwEKAQ3YMIHyLIuIxy9zN
ZDduLTfmnan5IoT86bfl55SzvkOUwKzrkyd898URrSIMr8oG1Fki3etfREQDOkL8
yknN4Gk7x4S6pjXxdptL+z2giyQNkWTREUebArIkDHngc750Aqa5T45P7QCZgqDK
defdepPtsBxGINBWrOgP5Bnl8OmOt9+NW5nRTHL+J+RLTdC5gF/tmp1BikRO2hjV
BSC/Q7aq/64pjlZ+mtFSJoxpmnaj4AY9YxzjDML4PM/BB9M4wu96/JpbR6ZDrsZN
SjqVYm6aVAbCa0xyr/L32Rs0uH+3yVseQAqniubiyl/qC/X6sRTuZ83Dar7JrG8G
ofkFMxCTRMyJUXKL3Ly8k0k0swurUK0otJZSZbcMkvomT9gReZnzYHH0JMRf1KbP
3LkFaZxpW6ZeP3ftcFLML7yzvbBHdEKImEyp0O6kJW5JyqVTn9a+drCcXaa4XEt3
5+EIzbzLPpub5HEINsEwC3UEHDkckHpapeOQpInBGTlT08yu5r5uaRLxJvuzsRPM
dnzJqqSTtfOcLXBZY/6H0ffUtHn/ccxKvHx+otYXmbCI9txfRUdxtPrvWL0/oXxR
SvYpEy05nXQ4KiBgvxRcykbavNDyIG1A9kH1x0+Zf37IUIRQ4vMAt3njfK0JlWZU
crjMT7xoMBh4uP38Qc7SSVPa7337kOmImqCQWRs3XtV2/Eg6uUIgDRQgoUJnKlhV
X76Dd7njsl476zHIoG246A1pEgoMGiferWAGrhyYAfz6tN/8tstm+1FTZCO5twUz
erouG+ww49zsAMAc9GUujtM33wkIGMj62sSZBEk0AjTdCWSulXe1ro3AUnuiW5yJ
2nOLyyrXAB2kAVoMYVugcGlUnznhTjJ+5mJFyuzpvTGH9k8p2YZbVzw3ftxKJvhV
gT9y6YTym/Ru6sKCbfKnbfMoKgAE7MGPJYpO2rXobMwuGrwHtCfEQZ7B8yZEshTI
Qwb+CcA/e6azWAPQLRANUy42xoPwT1p7U9ShfKYEW6NEg9TObueHAU4pTxK2VAwB
3LHpzLp2PVEAzIYPy1hGxw5WIv4IUJJf3m2R1QLLGqzJtRqlHexRbVqDUSv/v1XI
tQ1kKz3Pmf8ymzrVQLnrWY82EDT/1iJf4a6761MAQ+AJeCpMPf+yNZ8Q+05OHNmf
jfqJnDu3j/+hT57h99Ib/FgcwFhBmAsyF4SqhIFEwpT4IvvrJNdDcLsVtqjHI7f3
alhPbl7jDk4G55VUUumepaqY7gfOeNQ2IQYHeiI97i5BBtMGdgu8xm83yUQ78MkM
FvG0h4cPWTwmUkcm2cLa767gj8fZxIvDgpuHpvwc3LSnFD0/EscqVAJ9FSYTgOS2
cy/i6BCOHgD40yiLu5Q7NGVqgi5bkO5GqdnNDl6DtQ94CcDK8nut1FvEswZZ7poL
Smwh3aW/92T+u4PkE99A1Ls26/RdshZ8maiZzq4pLoSG+fKs0LwQ3OvvwmrZqqpi
SOSUueSSGS70H2nG1/Yie63hUfWp2Sj+KeFpxUD42fvVJ+0/0qaMDvtUNx0uTY80
4P376xLlRPUxMxrdUW62kWukf2QiN6NpoWA8NaYDl1bCeIo+hCRNs+gpnvKZiSMM
UfME5x8+vIqsLN4JyEVzJTJlqHxkoWeN60JKyezHlIMvAthWhVXa3F2AQj12CDcl
BVTP7Bjr8UgxhIImPWsCpoNwyBjRVMEONdI0lCKr4b3hYsK4NHkSMGB5kuUVGrQr
/bhy44Xtaij5s83DgGI23oRmwh4exHGqcDaJciIlrgq9uqxR4yQBbOWLuvOVCW++
AUCyWZI3fPAcO0yrHvxFgs7+WyFarMW0/KDqNkRMl6VFDmwAQwdDxNYcMOwNb8l+
GBs6OcY68DU96BvlW45eE+Ig3kSAUGO7F5PDZl34J7xgQHK53Aw828Uo+GU7YK85
DijCyFVchF6FqST0+lJZeC7VyAWsLsr1EMU5Wft+azVfB35A6iI6N6XbMIt+GdDq
iixv0Yo+1FkaMRYhYb8ruHFbWGQ6dGJVCZl7rqalTB1uRjiOWgeHUYIEjt2xzG7Z
9zud4xtU1mDlFdNccNTAhJbn9dsXCW1EK6bshEKIoQTXlZkfIUWPRpMB3OEN8uwB
xDcqVS/LTYTMET4542h/Z3SUCi8swNh61DZ/zc83JSwyYUsqRNACCMnae4dmlNjF
8uqAo7SOVPQbhhlvwzwPzrti4hxiDTzQBdSl23sz/G3UUTGLW6FzPqQC6/TY0H0Q
jgj4kpoxEY4GIdh7s0QRxQ==
`protect END_PROTECTED
