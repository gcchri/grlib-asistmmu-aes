`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r87dtIKjyRdotEL+FTTnsc/QBSnHuqPsrtwHO0L7KRBAmGdKKyuMV3kdCm8XnJo7
lXse3Q7MXOVehWCcb87nxO0uwFcymOVBLpWsFDyOIgDYOC+7fp5JcT3bMa/2BY7w
wYtGU7FKBOkG7Fwk5YuR0OHCPvRIaugnhfnTxQH8s9jQZCDH9C9jyEeHZRsREXTD
uTqfnShHi8PkajHnn+XBTSZiGHce135A/Wj6V9U1g16xBxRG6XoHxEOfBkFLXacG
tH3O8/zmxruyMF/1OLuAs+nb3U+39ZkuRefuiFkFeNMbrElX7GBgpGYhWxqMXf4E
VQRklA1Hb4vTu6uDrFrp1L5CJ9nCbZcjKGUoDcGBGXJ8lOI+EUrgI3UX/MFMSMkb
uEWzCq5Fyn3HYoU1K0tBzmYkdCTgs/TGTuuGnwibaTf4rudsf+ztYBV4J7lE/kE3
8hEL6nduBmZ88somj9cM+YmKUmtEMR6VkNLOIMyZEnectSW3Q1rpskshflY9IEpv
GoMuTHsnWmTHp6a7AyyHikX4Nv8r7vRscj4BHWj4+ybZ6XvdpOTvdg+L1orpEToo
+1Suf3IJUxPfGmUPPXy4g72ve7BVE9AUp6ma7rf6IU8q+XHaUV8CvFFTCT9OrNJY
5Z2rDsqKVhY5C1l93FRqlfSbO5IR0m0NZ0ucPGpBXpB7y5KhX3wZpUIz+ttgk7rX
6okBmjuPm8f1No7bKkc6CEpZtsOJ/eQtRe3ukd9mHQBogWL2iZ5xatTGIIdlf/LI
n0L3hbu2eYPdk/W3R/BAfmkDc+bt6b1tVpNdbuOZ40dH/61JgtOqMxjRAdnbiCVb
yjwyTwEQulLDJCZMAHviJLSNDnI2Czwmgnz0n9oM5dtyRYRN/WKYlELSSbo4AuJW
CATOf41X0mfh/+1iLj4ofd5TEmx4D06/Qyar3CRDcxsaF8D0qvj3I2x0ZsgxAohI
2oQYdhuhhcHlFZtOSi7YVcFRIgesa15K/wLWzMBFARlGdRAUAeHS3suV+xFrApNn
xqZapf8rN5Ujry71WEzvo2C+LMiuOmOaNgI5VUerVAXldVepx+ddsfYofHzc/de0
79auLQVSDknQAiFkY7By8Q==
`protect END_PROTECTED
