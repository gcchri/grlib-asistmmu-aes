`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x0lWW4Gzvm9NwhPtj257ClirQGZFVW6HFpHR123EOxBy6EqP/Jspf4vaZO4aTz49
LCf1dV3TOY7DD3/QvMIclKvn0UDH1Az0gbtaHxYRGq//tBRVDs+em9nXa7ztW6uj
m7JQz9QPhK9qTRal2kU5bhakDz0YjZSWX3kAObhvR4mjwpPrkjCsaudgI11nF8z7
X4lg/8NvsDhnrTr+aysOWW0/3sOdtAeoEm1MbgwuUwjsI4lS57gs/BeyyRJPy0wV
VQvzoGMiB4bAx0GHbVA88A==
`protect END_PROTECTED
