`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJnmLe9uaY0mwMbiJg+CgWZ1b06CnS73xr1z84QUsOleYwNjsn64HL2bFQ0sZHgA
+cc1YXXd6O5eU52rHssrOPehN1Pl6iKSNw4SokfH3KX5z+bncqJxYSv2oe+drzoz
k8f+fanXw51GBW4gTuVmdniESSj0TLMIFBpr1p+QUDSj40u9U7vUvL5P1hQPUHxO
grFTCojaXEmcAMqrANMqUzae6cTOvlEsaoOpE3Luu4KuufOjOM97L1UbiVMOmlAL
`protect END_PROTECTED
