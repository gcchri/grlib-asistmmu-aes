`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+spBOHMuPDSeMZETF9tjwQx/wMdvKXZeuJguV7nRfyM36BRuCjZmLgNUNe0fN7bG
OrL+nmo/FXRU1VxAX5Qm234xU0IaTPd31abu2jJq2HEh9RkMXC4MUe4UxEnwfnzC
w516TkAUJTdMbnPT41/Jz5uQe1n80cSrEvTN/obsc6cks2D/zQqC7NxUgRzl7yf6
Ex4DhfTOM/ABXDuu7s8eiYkwgbM7FOsRIlp6NwajThgnpoiF+vL+czWIyQoHTfQD
9NDFx0PySRotm9RAz56jUyBZ9UkNURvVJUrkzSID5FFFMH+pgdD7bIP617ChE8Tt
rFTGamlJ4tOgUQOVT6nhjQ==
`protect END_PROTECTED
