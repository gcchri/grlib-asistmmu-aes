`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ij6lmZBjTWaDLY53W+kctiPL5jEoTq3vo1W3Ys8mYPPp9Ku2ZuJAQ/yOWHiocuIM
Dm9xl+aTK9AtqzMw7XWSJq4NddvRJJmu3rIWyfXvH7hBLPzcZidN5tCbkYDvye7D
0A88W6m0rItu/17ocNmVAtyxbHKZObjrM/U4NWagpLGVCFU2y1VHq2Z9DPPPjMy/
ylCdEMqNRlXp7yv88lTS3rhokXQMBrMwXfjyct7s+/gpzwCXgszrCI/ISzOXVy8d
AexcYK4hbTokiFG86x/DBMfu4PxLPM25Wh8m+zE8XwGgP6kAJd6RC7uuuYiWLKWi
N+PZ0OL3pl42iBG2cW7q+KePQEfPMl0C/rVH3xC9pQgMTzKvDZgnX3XzcNtGFEze
p4Y2j5aDxjmVIzQWBVh88YJJ9T8LmFx6X40m9L1YRk7IaGM2179nDfK6yI4StAEx
AfR0sjk1UaYyD3f4chqeXvkCnkGFwN5NHuJfkbaxu6HIOuCYwQj57wG8dX6A20wM
kHC/kVJaF23WMEEKgj24SCoKXwGe1h0rcx8sZ1Mzu/mIqstD4O4Oe8d3Du0S+JgP
Oiy0J1c6qUEgnB4mY92VM0FYsdfE8kMYQj09SpsHAkK6OjEJTsZ6llXSJxYUjRmb
BJVMqaZ9Pjmy6Ie7FgLJdABJ21bF4CqhmdHUovmEUIwDZfCYbkI4RNqhRDXZT6zE
abgM0UIl3sqHstTv0DR/urDphecEcCP5zDJG+4PDMoACsMGl6El8zvne1AckArNB
vfycilDtl07l3bqhkjj/VvVguKcIsWe1+SvddriZCOCBclNnUSsauShj6y4d9h5t
BzjGrZpdK+gbM7g4mqBZ7/MxMd18x6l5bxeDyy6msWqDy9wHqbGMYb8Bg1SF628+
PtXiyxwFBJ3ksx0U/7msPGUHU6kr8QWzjpl+hu1mQSPRRvtiSmROA/oVORaH0B/6
OJYL5ZmIFtnST6Htr58TWvjjnBTAyDGdfZ65WVhmhqlSH7UaeOQdnh6d+RTcKb29
kjBWOZ4jP23VAWlR6noQarnp0uspLczEUXzj+iuC0nuPHHYp+pnzVezkvkGeApSe
A93FSwPGkW7qcqczzfWac5Y8VRNBGi3kyfknWSj+jaqJnmLrnFKHy0VvqbemLGne
0Cz3pcLHgppcbO+GWlGMmjcd6J8nF6yMjmwyG/3GEhuC20EUirwMoISaJJf8J42G
CXKLSC6LsqaVtC5VxKQrbMWq0TSThhWOXWe2+UX7IdOgPXkJBVPhitf3DNZd9ZUq
8LDzyLCJsxTSzlIuM97OfT8zB4/Uiwyzo8IrMvNNWVRUifUBmrRNSwX/YMER2Kll
jjmIpTOgqPBVEcYmA5rI3Iugo24LogSBRB2GDGwVVJU7WOIYM2F1zPgLOWlFsitO
3ZZeRxY/2Ye8A+y/Z+hQAcRKjiB9Gei6CP0ZmSI2aVTSeiUSaLHshHtNBV47o0Vv
RaneXUCi/YOwAdgDsbZGoH3fP7E6wLNvCpctQ98ZrgnBgGkoHZ/q1BUJkwPJ0HiZ
z6ZCn+lohYzEJ5n9uy3XRGZMwgiXyskAYeoHI5Sehbw8PW9uk6Cp2xV/4cfPGGdF
+uWp5qdQqQjLJ7gXikhuSynEjch1Z6tReEKFbBTMG5fZG9y+HMKOMhLYdflgivFy
8oK9e3W0WPs8HKAkVvIaPw==
`protect END_PROTECTED
