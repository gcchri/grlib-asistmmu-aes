`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
st9Q9cyXk/y8K1CczSHmZ7eaRRSlvPnl3MslpAW90CiThk6KqkeUuQP+YNV7N0Qe
2fRXoObFVweBCFsNYoz568p/wjMrjQ+Voa+Xyb13zAWXu8JSEyJlRPoWsEz/YfYH
o3UNju9H2AD2Y9+iSgMrgqxVmFpKG/0oGSdrDN15LBvPesNW4534NYKRXgHhCQzw
RNNZOccqfkHcCgZtJ6ex76fFffblZcdtklNiATTGgU+Egt04D9c7jNm1/joQXrst
EPhPqSfkmGkqLh2sZeeb/kxHM6lfXZdULc7GE3hf/Lc7odSfZjl/A2eDVoZr9xpc
1mTioFA4fqSsCsZ8Jlo30OzjLp0JBJNVQCdkMGsjY5FAY5uxkGquFqj5drDRqyRW
eKlxTWzulaWO/wDBaxi6pA==
`protect END_PROTECTED
