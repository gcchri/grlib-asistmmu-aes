`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VY1jdmFr2cZX5O1NMZkrj2P2tzOELsQ1Cot7h69njFlzAtRtXVIiZmucCapZ9juq
MELNYtuzU8rGp2yz+yH06tdgikIhI0DLJiLaOBuEGh78tVqyCsSt9OEpjJnfCTK4
gqSoOG1rU5UGCVFcaka40EF4AcvHjPPqYE+Dh4IYiKgpzwArWmmovtFObxw6L8nf
UkRhLNKW1J1SMxYnyJ85e7/wqiWe8e2myIwLShbpHmn9bRYXKZ6KIB/X6X21gh6K
xJpmG92T2+PwTROow5420ICq2ERcTh8hl6UjPZJBqxx70XBzWLUh4hmEtCjBGQ2D
fkrl/W8n9KDD3yIfcG0iePvDsd+rXCr28kT0n/pJLekxe7aFf9nl0c0xL18ERF0T
vC5VjxuZKVyMG1hxb83jbw==
`protect END_PROTECTED
