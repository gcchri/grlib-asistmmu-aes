`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
obEP4otEqOspOR17/7UzaWklkXJqL6bmVTi8c2EdTDCSXSknbw5sWtyAeUUd6D6K
R1jiWnct3XQrD8e/NlEHVcpoc+33Y/EthcfsJyocG3GOMRWWa0prIy9h3/dKZVpo
ttiZvqdoncGyEDmV01CRNewcxLF27uW+aMbzw9upoyP4J52rtrd2WkpUGK7okrhI
rFfo82N4b/lCaQd3KoWjdmlJRgZDMwaF63DnviZLQ2cKjPUfSBTuAJdf1Z2gSbXP
k1O9aKVjVcV4+k/AaAMDmUOmk48TqFeEDMk8Ph3jwDWvhWSrPM+RwLZKPc3AEtHc
FTKG9j7WowYLWYiPGfIa9/HhYeGDdC3qbuQusHf+pUQEIbSOLk6csx3Osg81kIvL
DZsB4yKLhLk9H79BDrL2xi2WiFpWSMyprwtaDLj1ooUVUM5KZYGur2f2pu9/8Bb+
fzEorQIAgZPTTcwaoyQ9hEX20HQhWzxqhji6Y8MKzYwiq/HlCBF1itQL18hYK2o5
8g9Aoa5nxCTxkSJFJgEq6dgLGmABV0QjhuJ2lB7Nb9xeIv+j4mX1XMpZzib3d0uA
qLJiuHDf7SaDQD5Bixa6EnbuuDxP/HsR85LQOxKaNhr71c6Alu6DJ339lk00pZQp
znGp6+NJPmkcsBCNSaYjDjfUSwY8aNC8x8xzvvxbHXYJ6WxJztcMDj9IRy5bR7wf
Gy1dYeZ+DQg2s6VGtPt3xfQ48KJKe+MnCy5nQdxI0YNWyaAexrh5ZdRnuSCCE3Ne
R8XMAHMJI3NA9zNBUwlDJXn8m9soHOU9rDbtgre4gi8FrIpAn/r0yTzKcQ0HMoYY
`protect END_PROTECTED
