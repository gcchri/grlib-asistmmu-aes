`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5dWAmDHDwK3DIPkK/5DkzDtw2ogcW609jtSNiGeohS8xjCkWEfr4d9lcnFBdK1U
HeYObl0zD1WUlpx+Gx83QmJoTWp9uxNaDQZkh0cSSQ8W2MZiEvn9MBsb95SyKLzq
j64JXNcxBrMTmwHNBtj9sA81t2eE5Lfn/BOmy0aaf4lDk+qyrL5Dva4C0/AXry/f
TUIQ1F95D7AkbvvsmbTDg3ices8xLSY7LtqaMalZhomebqBtd/MeYPJbMRYwMMN9
0PNL8DC7JYNgq6D8+zRmxGuWQ5iOkgDNjnz6lP4CvTAn4rKZsSdajHQ2+2Ia+Qfn
x3u5ApSNVrDn0ifo5QDULpnyJpheKaSaXgTri65ttUiM81pX5bzreLfkeN5df7AB
P1uxFUtUJCp6WOFmI67l8evPRnLXOXxHlPI9CbzU1eTefzIDrJUAitMDxB9F+9DT
dAiKI7KDHOEvZr1Uw8d+/JhFcr41CZpwAX5Hx7c6J8R+3sPnFtSMyU1M16q4f4BJ
yFQBw9ZMFfU1uTm890PQzc2kmm6MFqHGk66uJQSz42r8idK78IGZX4bN67LIj6PJ
gHIR27tlHchI77K9pRoI5W0MJNszeJNw6ftvsMet5Apl07Hi/QlpPMPrV1qVAXLK
eXHJAPU2nmOjyJrk6q7KgO5zQhT6RzGy7HunXL/1uVAgi9KfLYeCklEO3jqmkzjS
WZzfNNayyYOCbhUv1k383bQW2ljy31w14IU1z+w/hxT40NHZpMYN4jBx9aNxuMSu
L7dp4woB0UyLkaoUwpSyURgwGfA5JaayJd2OeFfI0kV9+dqdEB/ZMnxefbob77nr
yxmj1WP9zXbbENLF63iPVypQjf2aXe6GAtrlS2coeDg305y0fFJaUoz2u2tCZw+h
9+iPo8AwYHwS03/tv+0vZt2sZ9l2Z60EFUj8XakS4Kc=
`protect END_PROTECTED
