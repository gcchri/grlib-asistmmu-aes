`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+4ZS1dw9W0kVwji8mCmxqM+JXie8HObXwfIyB3uFxxbSkP5I/M35e++nupz8Cwv
XUycO7wOuEE8diSRwha3T4v1SHBRW4wMCtL+wBiDRyp/qdW8NpvnmD+6pLgMQLMk
4QwsQhCQ8nzwX8U5b4nNmEwRwvZoosPd4EkHYomuDHg7Yx1szvdiGPAN6jpUS9v7
SZjsIkaIb7uiivad8cjnNxjdd4xDJHcgvZmirUWSeRLhxU6kjS7MRZKyJpJQAg9g
QrfzhU8I5E4rJIRyK2oACvKOxRlMj2KnXB9vH/MJrAM1eMrzicI5RJ/9a34yLh+8
bDZRziJ3pOrIqJF3qJ/IS3Io39F6iSxi92u7MzLRenUSFA0Dp0pyu+TNqclMOZcu
sYpHUPbfWGvgVf7WPvLOA9sWqt8hzED8vb3GW8BhA6UntexIb4JLzEgAaFkTUGar
/ZACVQsVt3iBglHYWrdWz1tsgZs2HCRdqp2Cq/0alOsh5bMJjKlH85MVWdvM9EQO
DoVob0yd31rH/t3alPKIrTVjGXaFdcNu2gtoE4PE3XQyp2+SqjslT1+hlIcJJnUH
vtWLR2Y23bfP/TNBIzsAb6QpTVjCW4lumUxf100WB1Ng6nKet3PzI9Xnp0CsV720
b9qdpplpWBg0R43BVfJrEIz6CxsCs5HYY5HkEzTqOgXVThP0hauTOcuLT/wgpgJL
JdezsYQk23nxdiAutUy6iFNdTzuAmFj1dohUEw0V70b8aksOqMiXjSP1H/AfikPp
3w0MdDBUhmdVi8GUM0mOM156Ea9HqteZBK6juWGMP2AwwnCsLEvj41TT+o1ClaDQ
d4FjKlVpCXyE28WhOjvIh59/qjHxFpJGh7XUCGM9QgfYEhdJ5s5YmoucQVGEEYL8
qfxkMQiysRtDOiU9KLCO3RF6BtWg6wUEUgqNEir4/mVZrjg2k5OhqNh1o02evQyn
2Bk2kp+RZjamhZhCOnLXxphqe5A/tjs2LLfQ7izsHYDWFCplS3nr010Sw7wiaZcs
svH+nOVR1FLXkHhlsNFCDLj78h2Ua9Psp4POTeynQFxIX1sn2/tyFv5b33lN/AFk
ZVWEmGLBmnAHvNANfReIK4kyTDj9qZFEDdJyg+SoglqvatGiup3j1u/AWJHe+vil
HBuxoSwa/CqRKMamCAwyqEXwC7idFyxDJoKTxcIC6AEdtVZMj2EFPflHt1SxiQpr
fgBgx6F9JlyHwZmxmT8O33zSNHGcHol8LMRF7rPKWdshNEXPWbIy+GES9n9EQ0Mg
gDByRIOA2j8MciJOaXQ3OJb9PPN/hZkW7udeKULjdZV/XFZA7HDVzTA9z0u7IZcG
3KBEqXGbJ4AScKZyin5o+xslhJQ56/ohe8acxTFd4frXTDqlxdfAtI3M57PnVGtc
hJ10qQoRrO2vayyq/NqbVxED64G+5yD0aZQBrNWk7P1rF+ElbRv41WgbmT5UEnFu
vOI7hEJha+mQxhMFKr0D5IwPAacznyu27/r2q1lWJcVOqf1b9XFqt5ZMbvJuLKaP
ijZdN2xplMntWgXPlo6XQW6NZyZWcIESnx4o8V6n1t2UAjy2YlLYuT/Ne05daKMc
V57V1zI4JzrJUfOQt33jz1nskvgk7bKNqy7ROsFZeqQmVKOI9RbE1RcKCDyDVBSo
QI7B+oQyh15PNagiCalOsUjSFq83rwcMYutOmD0FOG5eLsIIhTfz/WKAiUFeIqSP
FhtTU76sCXkB5KlwbqN3OL7ShNraYJPXM8QixUp6g3z8zXSXiU0ELsdhhjpuAlTS
dEzTTU/hdRIGLXbx5uMFLf68ARnOfe3k9+0tmHr8bppZL6z1BX2sXG+iH58yHfK/
KXVcqh9xB75Pc/uTdpiOUZYgcRbKny8G0PlMBAyiuA05NZpQogGqolCX4BhklUvw
en5EPRb3ZiT7tHe92SFbDfAQJR2X9gS4VOtA+byir+5j6rs+AK94gWPkdITCIsqF
g64sEKLh2L5MhgWaMtvv3adOXO4SbHhryOjXYvRjARgW4pfc4iX9ZoYM0UoQq1/Q
pJ83kJ6Cd/IchbygAb3DFcqeCojmxZlUcfpNduy+zNJ5P9jbSc7cxf6rKOkoEDfK
3zoF69PACC8aWCDnLLm1m62AUQ0PAlmxAidVuwRk3UE6gJRVLTJruGtVTU5Bb+hA
Se+EWNMbcDAzTt4f3YjrtiPyCJjei5ARgHD4C66kDBjHykMbq3FL62yQ09it7o2B
tT11Y5uYJJ9q0Fum21MPphbIqUGKlKDWjfkveBkgcYo=
`protect END_PROTECTED
