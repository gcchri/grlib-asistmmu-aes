`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifshTP38NAOc0B0h8+j8lIghyhIdncTqTZuuoMzHy6f0S1Om0cdZnSFYxcqR7KEU
p0cWL+tf4tKsLQN2nlUo1E73Fzccynt/Mss/11BOoNSZIWf44jsc6zhQXN38KgIQ
oZhkspRthI4VNnqGxsZkUT9zkyaYiJk4f5QxUS9o0b42Cwsh/pxOZQOr/MBsizsq
jjc9ZcqWdU7StuRZT9u4CrMt8SZr9XSTx1qxATxHa4ovEsvuM/Q9R2d8OgZQzsio
UKkoM216rV6+TgSbC6wAAFuTVU6AqnNqvR4fY5K8o2XX80qiD2BQymUz+bEUR+6+
w15lAFNiwELvQYVwsZww+Q==
`protect END_PROTECTED
