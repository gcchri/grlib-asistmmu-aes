`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ta2dyPr34kPg7y2qQ1LmO5rwyO8Bqc1SG+8iZ2TDoBPbpT9JV4Jhf/C113wggF3
jMUQF2gT3FRjvHjIE6NsX6rHVJSFm45I/wuEKhRQPc82pW+gLDmSCz994bRiXm4a
9Ikr9WNg2XStZtDd5DEAnsJ5laX0IFpcjrBoMNNWnpzIT5f9UVvfOpvBGlL9oIC0
WOj4Mq1PuGs5tchLnGjVe9dIW1YC4tRTgOGPUb3c0hEgKqTN7RIikc+9UQRQPkZL
vnSakZx1OgvRySC1/gKsNU+I1lAMhyMaNzidRIzagX/mBcdswpJ00xG37xZmLA+o
kFZPV0lhHOCVr1NFnfeKsRQE8OPVvmasV1PjF+4Sof9mQjWGE/6mlQ/biXxM0c0+
MY3aqJDSv8LjIERwr3NdyiN1RuAKm7rf5++FJT5V4VU7yiQthAemGu7ZHUz1306j
BoKnxk5YaFaqjuJ5Niz0leiNtAf1CE4j0v70+n/FZ5p2oXIHL0PQlwUIXpm4oHyO
n3hm/jXx/T+1ckkBygNDK8sDzkJzyhbBeDgwda6xTMfS0+xw9DtnkcKSr+tKSZJG
soHpaaLgXWPXUoqqr4I46ess/JoHY98DjwcApA14gT111eV5Py1F8xJxUFzBhGgD
DnfnoaCCfNunKVXoTPCkJXlHKi3s4eKPrL90XJx6trg=
`protect END_PROTECTED
