`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7/4ObnUXCSFGv6ZjMlCDsAewjaGwYhushwOlq6S3/m4F97G+oS4Zqba9q+D9AXZ
Gjt0vkYkk6v7Mfdqu0Y6X91XpVQBR5FnBxqxCwxsz3q8Wbi3RQD1M9xU4P0rUs5v
0WUQU9WgDCKZ+dQWwGoY84SoVlOTX8tSySklyZ1p24KjjAWx81LhVFti+K7QXWPJ
e31f6HNqKyJAyGosxiG9S7YMh8kjMhSHyPe+npfprh7xQuZr+mE9/5OvkB4jcfcV
bZldyRFGUJEo6GSuEV58zpOS0DAz0tjE0T/1vRyd83PSBaAC1LmU9yfIY4Vyk6eA
8un+AWI3mMkX8YbdlL82mOOJJvlHSoWtAWySxXvH/FgvLJAc6pxbmEJ58FLedvnC
85SWQlayJ9UQCUxTIym+vA==
`protect END_PROTECTED
