`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wu1dE/Dd61PIJT9oBboObNgmY69LEREoaC6NnkZ/Xc0Bl8aVqL6A5ECkQRfxGN/P
HV0Jq6fMaYRYB5N0CAxAeGpsIlwYMgs+qhz0cdQWU3mi2FgveT537CWz+fwNaKza
nXk299P4YR113y1xpmFyX1/6YK3GdRjyA5qikhkTAAhc56yB4uMxFNXApJ0i3y9s
oDVYLEGdNEdi3jw/C3f6AmDERfgRxjEAfUmQ4ZMk5HiLlk+VIRr1uT5KmIz0keOP
iaRmRj7so+7N4Jkh+ri89orMv0cC6pITPcJMddkICviLrEQ9t0n1CMrO9gnmQYuw
WqyyJr7jazUMaQ/1XFnLrlR6UYpcW6vhpjWyB7Xpcv+u//4b3MNMWPIaUKL8V9LI
TP269e3aMzix1RvpgwdvjPR0uEhSwaAPQ3yxCy4aUpGz7mGwV8NK2t5/iuyiJpIY
0456qxfM66BtEhJRmEN/ri11ESY9owd6uDOgt3XQoEzhCAtHMWL2NgJkFl1tNVU9
1lqOb737DofjwtB8GgPDRrJLhi01uSUw68/ypHe8c367I3D7qNa2NM1YLAs/fgLW
HRLDERnVVVGxs4tYhPJ0GYbY6DoMKMfhX4yvdKpFXWSv8CJpJtSn834QOe/wzHh3
+0VXvUxnkIj37+XPMTMIQeGFj4QydsarsFHYo7AUJIO2QqcJiBg/ctPkjX++4uES
yzIdL0ftsLUBHYdmR5lflSpIbA9QVo8LeaqZKS9jpsUA91CFbGHm6TDQcoe+0H9B
wxluKWGgk5c+I+tc/VkpF/UkUw5J4tbtOi3nWoAI0LZ1eMpp2owAwT4a+oUwKraV
edJHgDaQxetqI8mZKd0mLd7Kr72vGPt2H5J/d3XQ+rhCqsgTbOF8kSiUkgcNSxuO
XEXNU/1Gfqyg16Qbu2QTdmCP5T0g2qDUeSGvQHMphiUer1CviOsikWnbYRo2bHHu
desv5y/r7UapAcMbvbSVOr8Wz2ku+R22T0pvCcHi6KY5lrF2VDLdA08V+yicerka
23li/+SvF3WXyEjzjG03Itq8Pw+w1l4qNuePM9lHwLiQ9+WZqz+OsKyrdqVUwMyd
yyhR7jVBy6KkrSExKpTKRkYc+/Y0N8RwHJQwGb37VGrq7J9ienJ89PeOCd42oLy7
cCFF1tBNer4gdFrnF8M3BrLM7GmVWD+TfVs040BSgBNYIbWhfIMkdKjiMwFgMfdo
PDrW31qSBpv+JpLlYNiYUKZHY3C0tiX6TFA5jvlJzGwUW5CwYEXSK2TRai8VegHG
BAPKlV2AHPMRBexGuV1NwalSyA/H/aK+AukbTFvG2uOApnc9N2Rzz+2ZjIdiMH1Q
0MhPAym6XSpWTSZxcw0lrddpCVql/VqQBcJS93pDwMrrsN678o667zq2M6QRKC92
kMzLaHdLpTA17GRBIsqlDhckkVAVlEBqhotB2+YFOrXZDqGH7Jsd54fRuPBydGsA
IUNz6N2uO4YpDFZXGzyBrOq3yOZzLCVMJ0+TCkNrytIfFwKfihLm4iJ2vt8C4OhG
ecdfPnmAnliu6DoA7T4lzvkLrp3tpybcsXYG0WgNuIunCV88Xen1F9S1V5g9fzfv
iDeNWUKW0RwXMb/e3hqgOgJoJpd5SSVdlq4VtKnz5Z87JL7cpwTj9AV8BL4GZx2x
/cLAvVMgJ/TlT9N00viEqcrBPMWexnUWhWmCsK8z+AK0wTHqWcdZGNz7KASiaBn8
suLQ0Qw2mKA6pszuIdVBgu2qOWcy+frgq0kx5zjkHnCIouYeLVnp68y9xqin5jgL
ry2LoWLq1yRSKCAtqpw85a7SgVyr07zTjhgDtEHxarSaKuXE2uOlYxjacZT4XvHd
kU5sX6Ku185dILSNwwYZ1zoAWVKwOs4xjFTbsyzFuZsqd6ZQU5HDi73i3R5YyX7U
sJ1Py6BL5ZWsTzJsOgbUxg==
`protect END_PROTECTED
