`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lxjmt0q2PQJsggZ2UQzBdHL5z3IfIuHOQfG54ExMLV7baTPfvv+++4hAu2bjhrAJ
ihev/8ZrmrnE4pJmcCBpKM2vJiZncmrEQW82qUx2R39T9L1j8dutnMa0GCJOFrQ9
D620upUO/1pxFp5n6wsd+qYQp88IXTutSXZnVxuyb7htyDDlzGmA3LWb+bJNsZ88
x2cG7nft+XCMQQ9mzbp92CuBUxe6ycyaObeomQv5ymqmZed8+NbWV8S4y1E48I9y
UuB1GcfyImG8XQQTBFilJw==
`protect END_PROTECTED
