`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jCgpPNSqpdHIKlNfzDvoWjzAvwdJgHF1U/mra/YuqmZ/K2o0qx8QY0tFIRyQgNNp
UM/YXIQeqC2CUWBQ0fl2/+mrPgpFFKVfYHFQtDXfm4OhE1xM+VVToUG+x0bpzbFg
cSYWv1lcTmV+bluJjDligYGb1s+5IlYkCOCo7wCWhbTwx8dq89oUZbIOUu1m+7O3
zuxIP1cTXO8wFVt5yUNb9Rj7gTMXLs8NqmIPeo+N1OMex3A6OO9x88FMzX77eygl
kuJoZichdvNrr2QALGR06bbKkPdUHtgn8auy3VQrpBJC7uEAksm2zUUFvBiJv5wn
qjspFgm7x+u9cmPYymZme8/NDbrHqIxvXEp4MkHRrMsSOHkZBG9TJZ4fp6oPvQM3
RGVJ7J/7+KSr8TIqoCXWt4Zwgjee0CCFm9E64Ke0eW//kDRmcnHA4lBnyqS1o/HU
rHlSOu+UeivlbahdXv0rL0il7HoAFD89gCGLUi1DC7ywhEeYxhvZMoQvBlprRn/e
V/hh9A97huTes4l/FkE8aeM1gq6ssxnxFE7wVStpAAzjj0vaa4W4EDXPj+Rv1Fpg
eemS0iTFdJ4EFQv5FZoRmrvvseeSFGmg78eG9NUyqLG2zYn8ndfnEAQh7nnT0w0B
y756hiZ3BGlybLk/w567cOfK1M8KfQAg0nxnS+ZV1PqV1VAAVRvHjomN9r6rho+2
ze8CfdNoZ3ynNiYm3l9Lz3o1ArM+Vp98zvreffsYdLsX9Hjsl0A8yrxvL1cQRtV/
w4fXJQend5aOqNtVmq3p9REysy6EkaaQyrYeDq3ewN1Yw3oYUt5GGYVcMFAJ147O
ms+2Jz6PVGCsa3JZco8cw2OQAfftYNuEOoYf+gp15FYqPWBnMLuJhBFfciLDKtjO
1XrnNlAM0J20Wc8UxxUqIRDUgRKKDvJ1EjLm7V6yLM47dZPtRPwN65JAmPVkWYrU
jUAWo9O06G379tfxlx+UQOAl62Uz+iIs/9/Fj+9oFQytoaC+VvuPY2feACfHdF0X
RBpInqf2TjRtj9QsBq/YLnPwBrZUwmg6Uq8w36mxGTRsH7+23sOfflNCnazfZBeq
vPtevrYPgXKfNs754YhxJtR9cH2j44UjHCAtBXvcxvypvhMaAigjFKmXH+wnPFhy
hVglMMAAq+dmTc/FHBUo4uU1QvWD312+kku6r3PCCfHe6wyMn/4eWMKKnYmiUSGk
bElJbuOg68eyZy21qT/Oh+soMv0P6gIVOkIbfIT0y2yNaZ+i3JruWWEeCqTkVej4
`protect END_PROTECTED
