`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Op2MkHG6Z71H2/7XnvXaa/izRpiwgJpNIh4Y353k2gO2B90usTyyhqKgJtyh9i2b
paj/gQdfDEiDI3xsu82rcMseNgBgr+p5AKlixkdYkBlCnG5tz8iTiPpcAvssAf2r
YKBXAuqu9rtWE9ZvabLAVOI36HYS8ARrodnahtGTNjrB2EGs9vC53C51I8jze4uu
ZOxhUKZhCUFF9c7Qsta0Tx211w+Yq01QAb7us8xXHZ4l57be4JgsYtmOTJ7UL2U9
0LLgD1ebMe71wrjfvq6gASdf8b5QJenEUlRCH3s4/I2EYU1bPyUrPukpUKyw87cG
RdQVhqgdSI54xNIV79Yl7w==
`protect END_PROTECTED
