`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNp0a/AE1LGuLAA+yiAlf1yZetAHbQjNdGh+Gls1cWVy0V4ZwzLXIgfH7hiJ15cA
/FALoWiITuBqmdLu09qEsp6jWNrHe41Dh2Hf3HVYNlwWIP4WwDF3SS6jH82idvi/
xsBF/7ANH8FxedK0hdP9vlm53eICsG5cOom5fvMyK0zdKLCH1d29QSAt+DIEejqS
tonbY59T16MdmP9eoqmt76Att/aegVmYzlTXrOm67tIGcmSloGD00rg8/80EoxHz
ZcPf0hOY/mu+l8TYNuHRxfwfJqdXAYvOYwziy/RF0+Q8cHv5J450JdJvtoINJf6L
b7AoJDi5/aBNEgWbIr+5yRrXCHJF0PfA/Glxuhg/gt25UoMuyuuukhbciJnthxVE
T3FBsvSlv8HvfTVwcxUx7PZGeimR7V8shB5jftQmom/ioYsa38FS1eokU/YBUMB4
Gwqw14WjiMJu4P2CWVMXHbJXY+uL8dHupwGOcJFRzAWdrF4a3vHQCge5VjpXIbNp
NlpuK+xDmsDFmxSgtRWh0ZW27nQADFR1HOCWK55Tm7xZVzKY5hNP8rrvbSzma9zr
ETAP79dqs/HxVc02BqUn2Q44CeP+ikuQs8s/hO2zzvkCXfrpWrfTDGlgpSe2MCrP
oWRw12ZvuTGpU/tSoN6NRvPnWLqDQ230G1dgNX12KHIm3PWp59M++LXb9sidCRqR
5lECSSnP01JgdEn/1hGxHamEcvm9I88zI30QRKBE7CHwFvCGO5kZsJOwuWAio0cZ
2HZGwfcI6E0YG72i5RaJ2A8I5UvqTKRmQ55FA4ZBrwGvsjXWpBMTwi/WdWekPK32
2hPAX6k4P9gSGsMu2KLQmi+TA5CqruZgPagfysB0fZYe9sTcuxtplMZ2UmUmNYju
ObzyrVezRGqlctUBdgJq8ZyHhfW62ItGaAekCYHCIUaXR0rlnZVjIW37EFjEs5bO
iFMnetrqL0K+C6hNYOTqz2MtVGqidnbojpPjJg/ua/JBed2YXvnDtsPI75zRacaA
1G4SA9NzUq7oA5y3SavhZKlLLrxdqbKDBa/0X2sEvtPbUZT7Jlf9iufjJ55fOeB0
9/nRtWtCsu//PM7EWX9f10Id+dyUMh7C+9KzpKcIZV2pcsimGVmJE9qchxeCCSdO
ZtOgJblBJxBV+2y2yyCZ3Q==
`protect END_PROTECTED
