`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cd4OcS8l/FeAnp7D+DiKr36TuSRarePJU90srIk22fIprCbJ8lkAVyWe06CN39AW
f27+PpvqahtQYNF61vPtAwZrEhs5C4pYcPdbqGOkPD2GDM2D/fKktCSxJShq066C
WLjLIWWi3RPOvpJjONrJGaFYiZlHPpf6uZxa6jwSWJTSBVsNOl/+8EQ6EuIWVG0U
g45aQBBmSzrjdXz3hm5OjDqLEw2M9FHuBKFKFCUOJ5Nb94BFFRD1t0Yw3G9Nbo6o
FsMA4P1JW1hmhkR0Zt9WJX/kcJ4TII5q/ruJ4YX67AQdGEOCmJcT8CxylnZf8Ld/
ccSY8ejIa7d5mH7pgNxTbir1/c4JdOTeldOUU84bXqW3QPPPMxtyvXEe/6nQhUhF
1utCQ2LcDNtLyWOANMWFPA==
`protect END_PROTECTED
