`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Co/4svmH9A2HsExkxFFVHshnaDyv8giN6c9yXt9lhEjGi7raMIPocSz0FVEZJojl
MRd0w5CEyhWI8t6a6W5EffMl7Wu4V9zafUSSt8R+pmjUmoieC2gem3ZcNw9kTllD
BKDo7ZrZxXuxZNuCWxMsud+9yX7OIAatMVW4/2DTsv4F70JJYSKKv7eff8LGJEh4
Uc2iMX88UsGcUbPqyGCXiENvIIM0iA0gssjejrh+3HT/5CFm3CYCLuFV5BamIw1+
RpurUU5wyNdsc6qdkgjCt0qwzWo+qEfF4UzPfAf0sa2+OooFbVyCP8lBoa2hoJ1W
cdMcRzCXIx5vlrjFlkSCa0QfhnLLQoiVozipZvuwHikN6YBJLhxG9akFX0MDkat/
0wABsFV4sc0wVBbgQOKJB1AlwfaKOpnG5x+djUyE2t0HiZHGanCKgReFcIMysjQe
CpkQI7mWbdT3bSGtkEWiIsvrNTSiBK2K7x/Sy4fk4uA9B5lOM1eYQVpmbjXfEhvM
xTNQTn+fvtUXfZ9Td5f9PMbNh6GKoJC2MC9N2CRfEYGltpsBr97dgxdc1ir5VVgH
no0lmVS6orRMsruPDVqZQBelYccyk3/48I32dKXkkVZp64ROLeSWH0Zldo7YR5WK
4yTNKMDZwLN68VzjtycSwqpAmPP9agVwXtQ5ov1LtM1/KTAJCFqDlzwJCXnHklcB
1sTp89UCTohuyrIVC7yqzWkny3aEQ4a/9QbMAl+CKIUzgJhRG/y27hfwJmPxAa6L
9/wkd0zp3AUOy8Lx5U/AZ7bEcSYhl28rVs2m8Ea5PjQxEBNygVJekF/vRLCeNC4G
9AbFonR5KhG2DpgEI0FFjINDtvn1eNRFDyIx44iMMSl59N5GDqwSSE6pvNZ81vV3
lsHYFmLJ7tobXG5vuXyROuM5cPfkWmGgxG15fYmvsDA6FkWtoI2yb6NbOwKm0esR
oFOfEsTsR8UdT+57HoeltdKVqsmIaT7rLyPbk0XTvqonuVf0V2Lfv3vK0bQbmb6A
O+zhJdhglYVgb6y/A6uk5gWRmQw8eVPR+bv0inA+uTXKYMD3V49rjUBpeJEu9zmB
YUeP59hzUE6t0rPNLynzFsN5UiJV3NFh0LFp2ZhQUi33UHw8WhK1NwPndxztmGPS
YWf5PfqkPzI/4QcX837yNqYiHm8Bo8m1rIDU/j3bU8XDUD4rOeU+eetdJgSdh/GI
MfeABdpQfpMlBPM6Kz3kE0d62IU4DKlsbQckvrbABFolS43oKuxayi5IEdm7gTdu
TFIcPr5LkHCkyC/kWBMhgEZCZSJbEmlvyUZxK2l+jGXUiZ5R3FVjTUQeUtgQ6ghg
8FuIeO3jjuJ5Ir3NUNtlFUIE72wu0L6OmlIvoSNUtxcSuEmX0rzN2cDPNAbk/cRt
E+CVRW+yO8XCxnzNRN6ae0uSHmYZVgL0sljI4S9rlRgcUrCwBvc9ZcWIhxE3TGNP
3ak8VbZcx2XYW6ipJsWsyAjH+rQl5NuyS8pp2VlBG+NNyX8DdR0kYRsxqo5Iahwd
KLnr2RA22HY5lhSTG4RBWOWgS9Ctqlz8PHq/FhSmStDO+Qui2ioZhBW5UmEE+5Yo
`protect END_PROTECTED
