`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3GHfhhKF6VYX3oG9nEzcTpTznVk/q8uNFalyiSKyho0KhKGuwzdbYXqpCI0uT6nW
yv2ojM8NhYADLiIqixJMDw4AGyE/AOfNxzY2LVfH2c15BLvi5agSB1ZRR+0JSqJf
hr58IIOkzavOR/KwgxXHStLbTKEZjtET9FZlKO85YznlY/ntvM7cUZSjHNHxuyZJ
dVLbe/1LE7AI++3abRNphK8r3qqDbMa1Pg8uqOYCo+BbIN+AUBG0kVT3M2owMzYR
pcr+uQhLwiUR/edJKkYUfA==
`protect END_PROTECTED
