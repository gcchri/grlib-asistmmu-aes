`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DaVh4E2r+XiOcDuZR/x3w87unmQpll0itU4JW9osnFpZzBkStWlCxpIPN+LW3HtR
HAYuXr7vbl8jv8S8l3VJ+vDo55Y5WJIJtLx7+sxz8gtZJ6HMt7Nc0E0g/vaphw9E
pcHXQmpIVvMyWWvu0gGCRrKlBp0nChiUwsCktFQQyvyLee2hV7hBSZYClHJFlFFj
oPBr6OVZppyKo3Ni+MGNdcP9gDhrSjsfi+rGzj1ILDB6GktdCawFRs5IZrGHEK0I
AX37t8PFlpzZx4cOwodSEQ==
`protect END_PROTECTED
