`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eUFH1znKoPqz64nZ8FKHuxqdFEcWdsuWZEocwEKUoIBmn2pr2crQ3wtmPmvpaQrV
XWsbpnzu45fLRQnBVvc24YaW77yx2twUhWPbv4YXbkshIX6R6DXi2a/nHoaLDa8Z
vIlNlhw7eXF8+GWPc73U7rH4TjaYeM42ySksbzJSqB3GKeBI4JpiGgyY/dTbSemP
q1JXruDX31BUisVVYLIUdaJ3fLiToqSZE4cxZJD2itJqCxvdZ6M/3xkBFXeCe3uh
OaNGrh2v4vdPFQ58gmbMLT0QSJDab1GvjBGixJx4xCulDWR4cbjdCvmmMFgBAX/V
uUvv/b1xFlaO8XWtEDxhzQ==
`protect END_PROTECTED
