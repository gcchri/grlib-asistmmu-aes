`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cm5Fw9JS5MrPrmNDOtjtzTXKPp+qQBSEq050etFyPIhBc7KDuhd8CdcQ190fk/gz
k8j1qkjkoe7pIhmbuuvAej2Ohu+sEZeaTB0GlpeH5CitMC2V28hD/Msu+O2/ygW5
l4eMYw/mfYX+sVN56Ima2vccInJHJTeSsiBWSHegMFX1Fi0OFVSRzINnOl7gmQJT
1Q4+DUiJKPdSALzvYepQlUOjHCUd784R1rIUunuGMnZBElKjXu0KHF4eLTSQF/bO
+Aci7SbsraZQe7E4NMFxa/GvhJWdaw1j6kE7nM0xwOYhc2E6LNwElbxnbdBEXEQ2
wsYQ2vNKOVjvrb+0ttn0uHFpnni9dpu+PS0L1SpMDv9cIeGEUbX4uX9DSr4pI9gQ
GUEo2WqcXJExxd5WAxBjhjWd/fKIg8Ox9cnl7fRR3zKx2ePMSTkULzanboZUiVX3
Y9gaGfHHD9BHud1YNSqz2ZHtkiDmfQTRB1UtolwZsQvQMRnYsgIHpS0n0IDIuF7l
y0oYFBmKD1TCPLHBbAFc57Hk1vNIIIEVrP5167f6ZgrLcOXt96ScavgxjXs4qc0C
3ceI0s8ZF+p98oMchLJs46GGepFmBBWOiva1KR4UQYOY4s4up+cIngcayr8r9WFe
376jIN+eEbzRtcD5bR3w1A==
`protect END_PROTECTED
