`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q4rrhRXw3LCI2CR9OimX8ZNefJxmotC5sfkWkjeUern0qEezuIH+6OgkEiVUoPN9
ye2ZDmwYmAv8bzCgLUrGWSPRr8OHZO27ZPopo0FuSKvnbCCoNdmd8zPvbQFx5UUR
hgwHlCcxaZTlinp80FZi6NHbJmWfHab4psEEPCxySBrSEOCn7XEqF4kX7Ba+pVne
BDecMHKTYAOi2Jo7YjsYfBe1RPwG4KYCYXtRNREQwC617/0Ttm07YYPv0zfJ6vJf
CQAeQyk54/C1gclfJykXkCMXekMtjaXumG3XW/noQ6J9GGFLKZ+NWArrg9qDJzDg
EPMZVFdb/3W5sEJ5v0xFxwF8hrID5muiuVRjancdDK7Q1Xy+HoJs+Iy0biFAld7w
GPA1w+kd/ZZVITJr/pARYQjXrz0AoL2Y/VwaPcPlyL16dMLElqsIlqkJB2FBISuq
BTk4ojwifDKFtmFpd0S8R++eSQXa47H5Uvr87I5ixt/KN3EyaRzhErTmfdxvfQmO
upD3p0P/J0YsLyBvJt6RtSQNWiDziR79AXVB+cmawjoXRcGl3D8HGyy9ss8qleq3
g8W13+zw0r2te/zObm3iQI340SgAumBnjKunXgM/KMJICQtCie9+Pd2wSQfeHE2j
Cfn9eoHw/BJbmM1ODaS0LWHgnoer14ucBAo2l+32emdF6rdsOSLeM4aCd+oFjOBV
Jy8csFkuaHUj2SPzv8vnQmvxQ/oLXfu2NhbR0bvKSVizE38q8oiR6N0JuiKWdqEM
Pz1xb7c6FsHuhO6+xsNl4hlDUbyMWY4Gg5cLHIxnw3+IXg+gDk8SDKaEHHMqWlV2
vXjlwYuZvwrDEBEkvIuV3c2NBOBhatfOSgNc/KdSC5/EMh+BeWu4OjYMKLexcIRE
BAdfTl/Ik33Q+hddx6auRkv+0B5WRc5CHjEek8FkxI95j1AEzRYjxc/veU7DvvjF
ir4qTgadTzwSWf0uGOC6kItzJguVz7b+O2+bZ0QTHxUs/g3kbaaK0wIxjxZqxr0W
vat2FxAAo0OzAwSlB77sjwE3RiUVYAAhmhek1gJWf1iTz9WTGI5D2gXoC15JgG8k
9mt+KXHt3pgadxAkFjT8E1MaeLYCbzN5AabJKsT221xaNslADKPQ5BwUN1VJP4QO
l9K9F/3ebzRTRWGPUcXvwD6aXDvIKuc3zsaqVY17xTxOKUFhhGDEk1PGHOVFDYgp
y0DfMtkmHFNytaZwoZeJzt4RsMw24SQcJQmGpG9h8cVfzZqbL8I0xYIScz36wBrm
Ulc+elBa41Mty2KLWYwu4EorLZw8yURbYGojPmtOBmCGlAvrgqzYYdfslEtkDKYQ
WozRPqYo+hnB7oKZIQB5xW0Y/fFMuoT5OKRRHpnDyIaOZutD/kWjtpRqX9aFiE2g
nOg8s9Yl7pl5VVN7OrwkjK7bsKYV76VgSe2NxDddcZGx2QBvl1Mpk6W8UXodFwHy
U1CIh4Lh5HEemdt05YqHRsLstMwU1bQI7C3dUpg6BN2hWkem7Q8UonrUc9VLdouS
9p7t10z+yswY99USkuqB8p1KGl7DAt433IERYoY4weFpoaEP+TBAOJMoyWCucFMx
+WXLdy3HpHkPF5wkbduPC8NgXhGNKDuCVr6yZ3BF0wrLKEiMB/feWye+ku201+9J
amK3uPnqf3qrJDf7v9rVtn4OYu07o9oANAuG3C4gCOcYM/tqAbp2878KV/zjF9I1
CvCdLFMTwhtZvFhLBcQr30gfO+jLs+02o4Aq7XikcomaLhnwQPfk90dVCpHInRya
4R+qvZseY5IeTW5K8xDA+7lCIPr3NBoTCSqvTaStn50f5tJvQXlixqQ2/gHX2z1N
lxu6FxvjKzAS8n/4gPdloR2kimkX2a03Bw6EVHqW1EcdxF6NP9Rd6VM9hCx8wIfc
J7sm5ekleUwjM6aVz0XWkL1cpwaqhI/vXvhztXsVam7Bn66qh8CfVrHbhWRsW8A6
UoKzGIhlukBCWcEeiP6T2qcGY0rcSmYhk8BuBOHs6WawMwjaLX3qL03KMUUkr3BV
2cjOhjRnUS8ZqCjtNISeJDD+A8RA5WEO1tZrTsRNvT4MJhINFjA6VJootGqY1Zmc
kZDOfzvbANl09Fh7HgHjkx4GZePWpO1dgwoj/J/SFIPe4RXnzsOMPKJ90XJBRlpv
6TJNc45koKaVeQHWiDJAH3/b5mbbdDHsbX6qakFUyFRGhRWiFDP2zITnciVAtp4d
Q9LUkyDFsWYak9eHDlvboT16IMwxy0L2ahNnfXhqhjh6TCWbxoAtK+0SMS5NO48F
WMkqERid7K/AzJCNEhRkBCrmhzWiKjFQvQ8Ol4mmU2pCRwCvgF5o9ETdELbI49ul
clVeeAPsgFuSzT9brn7vW3JhjdnshVaSUQMvIHJsA1RWo0i7vsdKZEE23cBL9CJe
nF40LLTVN8HKfNP8rJAzB9YMoawRAK3W8SkGl1wBUF/5kfp7dzb8uKGWuQtQQ1nb
oEHjuhFAOfm+e8a+xrgXzPX9qkuHtt8F2BMjptjITftCYGWNFgRNgHEzPkKfZO/i
LC6Q/lDyYhXDaOA0P8Gy1LS72rT5VVA36UxOtKyAN+F2om46I/C5GjHyj88DKZdh
iYLnbLwStiQYaMXgWGBtBHDmdfVqQvneJLPg3e/qpBiwf1pJZKkvcL17nEyG0dt2
WnyJKuk1Nsv9IvGG1vCbL7xUnI4FBsSncsxQgtvgeQ7qxKe+NCOpjHd3sgme764b
oP+qhu2I3Q8vnRP+ANYcEy7mmCFF9V+CwF1YU2wCsJndu98V3hGgMfVtDsO5TxNQ
b1cW7ql13iMCkEeIF+jEo3MT0wfL7WF0KKBzuprNY0kgB1h9vWaiYhGZ2uYskai8
spXM0d8+KTLM4dQyTZgBBBpJt21OwpbGnzUvKFbBJc7zziUVfvvUqzpR+TubWrA/
`protect END_PROTECTED
