`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+fOeYJ1kGQ/l/PbEFrkVUM+PTkVJn6RmejYdYaqnX4IiIjvp4ZEfSfzlyySbiG8
qDUP8FqeeDvK+MNGF7q1mKEM92ggTo+XQKBdkfty23uV3Of10SYrxLUiTxBtGCgY
WdGJI3p4jiyyzjpT1vhNNKPYd4ZmobiCSlqNuSH7UTvogO+wdYL4ZjUZe4u6D7V/
szTkoxJ6LAJRt8GpcrXuYuDQ7yIGIdUGQlaDYK5e9t82ynEcZOnY1zNnFVXRLnCp
seLZIZDczrkqqEk43YKyqqUz/JryDdkKV4UA+v4Y3fs=
`protect END_PROTECTED
