`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHMlkHnfqobEEooFyeBGsqpVRPh54+PTo6eBXCt/phMhY4d0W8kXWGcA/9rvVj32
vaDz0LbqwN3/TOBBrrgsa9SWxU+p3hVeAMlevIUKrBu1u9vj+a/rNVTThd45c4+v
jVNNctBSTh09O5wBTjPQ3aT6eol6WeK3wmCZynv0OdRem/CheDkTDCuqOij5yyGA
I0m/9Mu+f8NdXOnERDEgH0HD4pk8AEt15KLN0W9UpYCFEyHn+Ja8pa2Vd8w6Z0EO
rbeEsVeKpEtPm2i86FYnUTz943Ej3U2zprIjAJLx7fJkahT5dw1pT09YFD55KQwZ
nd6Z9jQFtH+5Vda9UgUep3G3BwjPYeEx+bj6IZv7ntKts1CZCWyf8HOO4hyEql3m
tCxUNZ2yIoJboIocQJjxAw==
`protect END_PROTECTED
