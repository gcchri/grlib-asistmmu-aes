`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzweKY5ZsPOcUBpdY7LVxWVdRGbQyLxNW3p/vN42UEs+KEuv0IuXSdCe5bNxoDDn
PM+RNxjRGvL9dfDevdJBiCCN2y+awAFy92OEHLMuG8p0VabbYKxUDEaPjkVZFzZ6
G0APp8h1v/XH83ciFcXVZ21uCD0Da6j+S2judCRjg5jp7PccBUj45HJxx6Rps50T
W4QOnsMv3DkLo0HNcE1Z6NSqQUAzQlOO790c/8KTehrK9z2Ej+D3wEMWk9832X9J
yGGN+XV8BU5zcWY7w9Dohy3FYxfvTU0r+glO9sF8DSUEksmAMSV5TNurpJtoghwv
+tEmkPzkNAEpss2I0QP3gSvCQbdijwFlpRt6PywbTnvbN2enU0kIQdUoX2DLo6ZQ
5tvG2PPAolsArpo5z38kRbSopPn40qmqWr0N3yPs0yu1mTBRbC6BsJq+KCA18WqF
UZbt2BFTcPhkfa8xQ/syDA==
`protect END_PROTECTED
