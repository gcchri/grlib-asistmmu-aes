`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D3rQbzHxlVXwMyDGrH7B4gDts78D0uvSLdFbRfYHRPyWbh1jxNIIJ3LOQ9tdDGab
l2Ya+DBdKGwTGtovzTu4Aq3aPjX1y3IqclbDtEECFnLdK1rkmBjtJEnBTdcPcZqS
li+NwWfsoaMp8m7M870YHHBYG4iI/6ajeETRsbYWLxhOuZgKgEaGhSqDMN8OZ5J/
wF0znykqBU3mETn4aiYWDC16+hySKeWa1m0yPOCSS9s8qLUyXI8bt5gVrjWRvCmK
+TBxjP7CwH5+8ZhgMkn0Myusv1kqdmBWwGY8XBGG0XuYZ1aHjJpqH/QboCCUQvoo
wy0GS2mC/2C31aC5iwewW4mzU11y7IojgwP6oq4+K7amIoJRTIWU2F8UEQA+Mckh
JOlmLeDHQSmsXYQP8n8C8b1JavSWVB3CPXZ9WGe151w=
`protect END_PROTECTED
