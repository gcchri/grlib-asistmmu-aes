`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDd5gV/yCaC2nfL24KyFKHzKIFxmhknQEcMMlQyyZ271t+6hREYP18dIQ9qyHto5
j1zwbpmMeTUUqtqQblfjLug9avOimf6NFgRFNLmA9twMgmlJJpLMcbPKmQnA1D6w
2mZy/Tva3Gyu9ffAN1l8wXfxz4yaluopx/1IoFMIRE5P0Pkt+3Lkh2r+ycZMH1Nh
imdlwrAQ0bCIZ3uJPWSV0wb1ymqVHske+o5NPUtqd9r2wQlZQZscGNXhXDC/f2nw
KqqrCl7jD0uEMUgR8Fk3K3FEkF6H1+zvU86NVG2FHalj2tEHrqA3BY8Wjo+Ps5B5
uWE/EriMjhQerXLENak+khH3cNiNjKr9bZdYlZwQrRR74brFu95Ku0YHM8+x3snL
y9FnqG7ZauM0KcJhdH0B7+a9PtZFALx22crUZQKIe1Ptv6JbKIROatmCkwRb/fwy
pPU/qUCjvY9+u3B/nUGZ2YFPvUU+s0e6CRLTleuwNVzl/H8H3GrxhyTzrh54kl8n
xc9c9sIN5LJv1EBcVKf+fWSqtSI9vfCBprTqK8NZ+Qhat+9M3oJRDzUqZSIWRn5h
`protect END_PROTECTED
