`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Mk9WRNste/HGCyRZTubWYi/INvDqBMsYDtZcwV+yzqa8I5LQevd05SCkizdhuOC
4N7TX9olgDaR/CNS6R53S07ReBXuEvWNhmTso2q20eBANNvUJj6cAs1KM58eXt/N
suv/5kp/8kdHXnFUxk+Pygn9gZacY4h+Uwt5w0G26Qt+/RVfZvMi5XYWwlEBMlK6
+y6daYG6/qy51RDcWC88k+b9bmzOXzUT4B7DSshQTxFjrX08VD3p33V4sLGJjdT/
kzTLCHxQ+Lm8bBGG/9CNSKQ9tR147SBsMfMenAFzbB8=
`protect END_PROTECTED
