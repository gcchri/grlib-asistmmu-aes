`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqoVRUZdVxE0B6uS6yIyRNwdPkVbDFgmKcHeYT3Rm+I2wLsKZEsUWgANc6yiJLI4
GZLoSj/1Bh/EmpwnyMUB5k+11kFJ4s4gOfuIr4NcIcBEEwiqypoI7Pu66AjFWGiE
KjEeQdk4sguMZMpqhv0S/THTXXl8QsldtGehPqM594XiwpnD+d78BxGmx8VKHJh1
k3W8bgHHboYO5S0yXd3C3q2d6nemF1p1Om4gA5hf4bbmSTrOgG7uFmfvnGzuwZ+f
nQV7sF+vrLQ2Qy+BP1T5WfNtnVLJISGNWCHJw90g1CgUEYwblKts7yd8tIWe1xDg
92m76yGWbXnXUtXszXLBRWEz5BZ1xAqrnkSWgIuHH7KnrEQJi7Y7CFe8dPAVrv3t
vjCehqHxaGQ9T/iTaiZtIUUWD3MBOOmzC4chska51UMVW3jsxg9S63DJGhDdiGR5
GWLzNUaQS2wCnEcHigv/ioQxRSI26OD01Hs6g26CaD4fp+SCzqQfNKQC0A2XPDfT
ZyknK+QiMTQrBcpNMQs4VW150ukdvukK68xoj5XFOhUWazAMEMrxxGb7rhyVc/CV
4LS30YKJ8evCQB1I0VG0JFfYlSVOLGQdcXtVBANjKSKks8iLvr3fSjfkw6bFKajk
DNILhT3sVWdMIx1lekBG7Oo7oRHv5mRUmzQ81rkCu6I/SPND2sOpemEGiw5oM6sD
mN261ypbwpoTsyDkY06cpGk/2OiwMqZTDg72+4Vh6NZBNKZxPfw4IYKqTOcD8DSH
Br8G70KmSotm1wBG9OhW4o0dTHQpQCCiMu4TOggH/BmFcVPLa2jmo4OQeRHarpt9
C6+tI6ru/FovVAIrSlU+K0brQFGFNC8ZOVCJLmu6Sx6MVAd9FcmG86roMu1ZxvSy
DUi/hSmzIO5lTtaZL+fTwQ==
`protect END_PROTECTED
