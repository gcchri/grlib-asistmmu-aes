`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYRNZUE35CI6I/MOlkQBtXlmxtO2dkL5pARCI6CH3k9xUbt7XHk9wfi5vaBOFyGm
MX+3T6YM67MRcq6OZAOb4OHDB/3vdSfu1iPIVFjw2qgJOh8Mtt0Lg4wCwcFVB+SW
wLZJmiUrcGTEY+Yc3AXMDIaiOetrkddLBD0xZfhtp66CuGtO8CRUnWAnd9etk+Ap
YCYfbQiQ7ms6gF5rbMe8KZ30qxOZMD6hnETMkr738pijtSf9M1cmbslqdIYylMxt
/IpbzgabkL9NNQsq8tTun6Sxx2qnBsyNfTR4g63JpJ5yD7/+pd2jEoNgX36vl9Uz
FUwUNlNVfZhcfznXA+Sf1SxIJPLGCJcO0qD7ICkuz4jFm1PJ105MeAFQGKqn3yur
PXioPn5ozVE4Osd0kadY+7HNkswfqnQOi0FeYOuSo1drawfU+jR8I2/yJLFTl1jc
iSCYRjfGaqxhc7A0luNjJqq4tzMioFLvCsRC4wn2Hes=
`protect END_PROTECTED
