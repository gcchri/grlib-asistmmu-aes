`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ojUNj9DXxg8cRtLLxQmy4jxLkWiBSjaLW3s8TjrQXUJweBueRl3DqSOtFTuwtQLW
YZUa/uwHPozL5EoD+uPok0gim0tSQL6I9oFMNQH7sIgZbHWY1EGoreP4oTMKItSl
Br5Za4+C+aSklyQbeMP2DTCEDuOeLMRQ44lfQT7VGlRFvVLWkEQrczznzBi2xndr
T89hw7Ho72aYIwsLJO4VD/XVGw36SIQ+9tm4AzgcZ+csvx1qkSz5I+jsSeRQ6MLd
ntIdaTCJZrKiOfKOsgYe0qnajqovb7KvaeO8ioNobZmfclKbWeN+9GRMFBqJ5umM
yLkFm1GrRohv+J+fFf0k3rfW1OLQKwpBs+bXTaAWcr8TAx++4HfKYu+k+CWsl5eu
/M0ZgXUv7vOfQHA0+b47EfgA1T5HcihvYm5TQXKi0mpJApK+STOoTIisUN/Qv9UB
0jPsfK12TbqTCgJRTxcCw+UmCXD9/AvPIGBdXg+cPzIk5aEnY1Iim8liwLpWzpsr
8BGIleq6boEUb7sz4HizkesCrzsGM+yJByU9oaLh0rS05jVUiOwfW8QrcPoj5fR/
NNpF/21kPB/syD3WTjlq2t304mn6W/Vg2ldwRuecXfBExBnB6A8f4vCLyxi2BK0T
i2U0jYCx9vxQXdAbdHbn2jTbdNG81dpfy8jLdLMA56Q5aGbTUQISsJ4mLWln01MX
v5Jba+AKGzDHFxfIZ1BTLBCfPcYLgmri4vp+/ndY8JEGowcyAxGxEgr6MOmNoVOT
nA/sgMRo1ZygN1YD20ZnslOiGZC2hBkpJTOyFvlcKEc4KUcsxf81kvPWg3RC/7JU
VXXHQmJTb3Kptxdw1VmJhE2mef0HOgppXnojeQJRkIRDEU2+Esc3fFDtkoqDSGO5
dMyZ2XYzQFs9bJWHuckJF59nVBlVB4ClO8nEpwjo4AUAXWOZWfQMTjV27tMOMYXT
R+X/FTAr0Wq89beANjbHPGbtq2CRcE5yVrxc/5OpYVmoDchi9cbeQFLhsLci/zv7
9R9Xo3Q1QpQLgCDaEcRechKNkkE3miRMmco4E9XvCaG3aMEbPCyx9kwkrmfuJjWe
8C8uZzMufkWkOKVwWsTGItJcZzetwnN5IIw1PZhjLKUL3Vh3tup3rzQ4Q3fX2bsd
WDrrWqj1Ga89LVkDnGSjODAF30XWeGiEizyhIyovhgfseMVgrDczT2blSP796F7N
sS9yIGedUbkZedL3Nj3hfQW5Zt2r0gUMQFWvNQOSqRBZG7UEepOXCrwzWWAh0jb1
+Sx6VQ3frf41aOedFE5BTyHQ8FciddQSPD4aODcKZV0UKy8mnJ1xGFc15aAtDH4p
cY5hHrbJgAq1OLBWj9sLkbnbyZjms1xTxtyQ7RKbPIBaygkawcaqsaaFk+Svw2wI
sNqNiihMudzvfLboK+y7HEt0Xp5ze7ykWz8qhWRchUHvPcZSGMHFdC7DkXmCgHSK
qz7w/8z7Bnibl+b2bNVVLWp+7I32ZKG0HYFqUzsfem7xaR57IJiV8nomG8kesvEZ
`protect END_PROTECTED
