`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldEMzluR2yHhZFN4YsXuKzHExZ3GExv1OUmPHQx1gzm/pRbW1qZ5mloSYAtT7+sn
+FP2p0+i3k6kY0hwQzyOLHWFdYilxalcvfBXHZBi1dfhEWM5EebJ44XhG2TSmXJ8
HZzzhjOynPqd67QKN3bybguz0JVxS3eSXVIZvampmm5bCbM4mlHgM1DSHe0RROey
Aobx4sLqcCZY0Vz+Jnpwa0Z421aQGQ4nbRmLa7Viy2XiiWmjMAxhEnloz8fSgTLt
n/Ipim4pmkXBmlU7fyN/3MnEGPapWCyfOlkw1MrmKHvO9Ro1FtVtS087LEwnUiCd
haY7e87Fhn5s0nIl7XQmV74C00D3H7IwquR4nGek8D8rrJi+D3fARnirTYk+vF29
DVMKWzquHhdwCENWnICLLulPqPzAmq1MzK4NS7fzoWiMGrgI7PMjsb6qnGPr04lh
u46le2t/svJxjujb0dSB3bNrNKUXcUUqiBcqV5uWwhgFt0ChspwAxcjpgusSta49
WkJUywRVeGHJUKtmbjSnWc3MkPUmROfO8YdxFQXbrZZmpuyW4l/zVCh+SFcd+69t
qR859WlCzggEbBB0Yk5/z0LEaIo09eQTPyPmuniVrv6uP37t8iaUlPr+FK8EhZVR
z/3Gzx+zC8I2IKyCwcN76TN2M8R+KOTTBzlDv9TJzun1tRbb3udE/bBk6+qdMRdR
8rBRkRZAO5ZB62w05Bbvg80N4trhQ15XAx4607dNfAnd/dx/NhM4tfn07YtB7KZ7
s8ojRctGECsh5FOwIic04K3PJnmSqZv7adMMGV2jHkpNDU06z+hNyiWNLTPIt37M
u/wLi1mdHHIytgksajZ43mvW/P6rlUhnNdmuShZe005LTtHBAuoFowzvNADKzFXs
Qt4z6x0HrWAs5TVQue/0NEncT6/FbRRXSvoCuWcXYzBGWrV7T6eQBdeL0mklODvK
K5lDQoPRS1x0t6NFommvcqeCqjlYqhdJHchwn69V89oxqTsdjIdN7DCAOHW8rPkg
Xc8rsGDfqc8y6B38ofe+qsLJ7vdwUFo2EpHamFolnjfXu1/wjPT2eRkHqCy48UTE
GRLMSBU0+zbHicjcrawpQzCRPllChPT9+7xuehPul+SBMIR9DLWsG1W7/nujax9c
zV/39BnE47+Ld+VfT93ppq64m2G9B8Frl1PAlfi/aI6wTid59qGBxcQAKKAPj/0J
+Arzhj5ZA8+MfIMtCrF862w3ONuMteAnDUecginIAKpcpvHOcK5vRUtVnDYBJy+v
BGc/U65eiXQkaSTBdcbjAswuu5giUcePXzNyb/Q9rP7bauX/vpxsijMEVzaLJzfF
CUK28fHi4MHgSkMA45UTuxakWqdaPRH7wE+u9npdgx++4Mzn206ZSVYlHfFAkZ2h
992RJ5LeVPgMQJYZEkmbHg8t57DnoDUsbw2zLOt/iF1YW6S1TtegUtD+EnU5pQzX
fYtxOxQqyWhD0kR6ypBWF/ZKJpsFefLiGj+OF4KNeialsKdi+QSne7dOhLDpBKPF
`protect END_PROTECTED
