`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eezqYuOWN3bJdiuKimfKaGZXGu0ltVImSjE4WLKDqJh1M4IM0le3ghhkio+Gh4hZ
iKnQqx0YnDzg04usnsgbPWSlpJHzV5mdz291RwEKHEQBc4Ih/+Zt4zWFTWE4txPL
lLAs17lRja8EyA3i/4qRx110+njLwXVzJlqar6LCyVy/IBPQ9ZjbqpNqGA2F+aM/
kMm2L9KfzMGF1NO0tcrOLOqA7usBFG0QK97Mn1oEOM1zZWEPlCw43YTBn/6rfYm8
L74eHsiOylxCl2eTBWOIwSMpwjsWdiAM+v8908vaFKdJ5ho9ak66BPZLjOUwPBvz
h9DFGR3ed60bI3Dgln5ncJXPiDcPzQ8RoOSP4uAwhQQ657J9P9APnyzqM9aKpDr7
hjUHG2l21nybNfahqyOxX+5Mvj+oh3UMZCBWrCfqPkltC4l1KZWxYWToTzXXB0x8
`protect END_PROTECTED
