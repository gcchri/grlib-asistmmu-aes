`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MctJKkfx1sR+71ynuv+baoef3LUPJ6nZwha49+1LUOnZgTdb/ApA/CjXsO7wXAip
bJGckBPi9h0u8Lra4kI5JW53Ya5iGrAV/7z942O6mgPOi6VGRYVs3lkEQU/sJYp1
Domsd7+3bFLodsM6HKKNfVZhOq0OuHneObu+CRTQX5xI1v75DrjS8OodZhNIFtZp
H1Ixea1zmWG7lNompetoLLhzk+Llay0DFDtxxc6XWjhTY2n+Z9omHXL2eofj0npH
Vcs51XUkZIrDkCqNjfDLeNzQ9Z35DeL+x+k2eGVuyQqisdBKZu7ybTYIRWHxNSuB
/sbN78YgeMXUr8boxauoHbWfHZta0omkzLuL9bsTg2WkbmbaULz5RxGCWwA7dAlF
+VO6NWisZ/ZzDyuM0Zb4oTFBc7fYSHK5ig7zO4wEcSPcw0dpZb6kNkoKNHtUgru4
/e/TaE1fXBRpuM6K8GiB7hd06vrVyDdr38wJ1PKpy/9BDIq4NczbYYeeOwE76rLf
GLVUsUlMKe98jfB1OktsHW6mDgHaMiePG1rXGT0AEjK4DqxjjWyKcPB0Ig0ZLj8E
F4KX8qlxLxS++KxIwnRZTUhqdAbGzxcO1pIulDUdwuOmrDp+xFc/Zv8pTAaZ7QqB
AHY9rdCiLiBvRonzxtsb6TFvsBJoRJ5sSIO54v1198WUUQ7w/kvAOBNubCvnr3mv
i398j1Z2w+8cvcIQSM6ExJCqnuIcPiqROQ4OrqdwyPWWgCbAFrVDIWVRFDaHai8J
J/qOH99fw9hukoKv1cgVNFOEBhf6eS8LcH5JFtm3S6jfzTZGJ3GJfUfZMdMsSRIG
`protect END_PROTECTED
