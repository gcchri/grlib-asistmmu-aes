`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sc6FgPjtJqZUWfxvt2eSY/wOofZZQO1TxLsWOQYe6wrgZiR268moR8AWGceS6ZTl
sLrxOrSsXb4abuqHPhUaVpNBXU2UB5zDBSXYTRoLPqcslA/Rc0VGVejjSGjlwP4z
uiiD7jtd96Wukiy5pN4m7Gs/Bka0jqZ2njgxEr+r9CnsRdwn/UgmV2QWumVH9yv4
cMbF2MgofqYaaERfSS7Oy7efp/ceGeyZauWKKnlUAYevPuA9+8ClDH0e8kW1+s/+
RfFHp3Exx6Hsq3eNOg0x75RV57l8DRqZ5O2zfl041A4=
`protect END_PROTECTED
