`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olE6HgLROSlOfKi65asrCEoysoUwyVD9Kbk3Dkq9L8Hl/v8ep4vlJhM6LKzvKNZp
vCVEcSNmY9C1/Vu8E/j/+BkVY8dJy9sR8qTBNHLngIcvGmcg1x5QOzixTA0fDOyU
oxm0bgvHlzBukvZ8cL9pa5m9W1sLRqpvThy1EuAGg9BmE31BrkVx2DcuECkY0TMT
gm2kzY1yLG4lrUp9+iDi8PmPUAn1fPUEm5Zozf99vg+NRoXzCaUEQZLFu++IIqN/
3oYIzZPUr9V/3PH0tLlpGU82wdaifpY4nnHIr9L5PJOGD3qFzRfaokcQy6Mki6g6
gytqZcg7PYWvrDaQl5NgMQ==
`protect END_PROTECTED
