`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pT0kZxSmJzp6xNcJ9wGtb6Sr+x696CxKLslInlCqWcUMsMK85d5IwVtqZ8/9uS4z
7LfTv9TcHEI2/bXdIj7VgE68b4w3cuObwd+O2pW4KBelxgAWSrtg/kRbD2hSbaoS
AF9y1brlAdFBde7T/NWPfssKwbmBI/HSuws3ZZBzmv65l7fJIFBmMgm7J1qwMoLZ
DqipZfYFFd740H5XHYKwiY8yqyB2lWTH9GFbQggmZ7ig/cRte0kxdvE17bqsq4rY
w8AlxL8Ch/SVGZwi9a2D14DFdFWTj8BwjMHgAjz9q2iVltBHzCIjGDwAjtbZgfGB
f3BYxdZKKCCwo5JjpCxq0DP77d9YZY9LecLe+YTI7jvJbPxD+DGlq9RA2HcEIM5r
8GB9DJSXB2s0byOtuo69gj5yY7gkoeXKxK8zamG3glU=
`protect END_PROTECTED
