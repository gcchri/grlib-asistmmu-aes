`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eCaKqlIQT3YUd1s21VonHaSeHNrnZGES/ujNvRykRyVvgeh+yOGfBGYlyVv8bOHd
VbJG266YEZO8psgYImuQ1JjHmdpZEE9TrDWO6+WK0RikRUcLAnuRK+FZTBawSG8n
5F1AIbvfi2w97OPJbEPzFI4QJZDf9U9UhLI+clc938geJfwmjYd1cA6wj+jOo5bJ
HxyH1nvdtJQ9oDTtK0o5pg6XC3Bo7+JPWA7/+anlvEKjbye6TAWIc7bWLOK36iRv
UEtkDQhi81ceJQKUC6ghzBRJiiOtaF53AFya3JGBkO+I9J4ZEJRpsM1W50zkAl8M
RHbt+AF/CAUEDqSvZnQoDCL6Q+ibRpNZbEPShcV3jDcdvRyC4Uhj/hVsOGl4L+1C
wVEr17xUYCv1jT7yAm4JULd0QKgHbWRwFrWO09zdUt9eFsdKVAGqqjyGeI9epADs
Sssuz60UrJBHoFkLfkjV7K4qSyGa4mLomFOp5dQLdkx/3OykMB8VbK6xFN33OAT2
0y2H37Z98t6WVjxiTrCid6LN5IU326P/BtBhy7z2DYfdcUYg2T9Y/5ZWJD0pRnv7
FP6wQvbOw2of18or8Xuz9qwvr2W8QRSP4aRushj6OSIqEkZ2y4wf138/W6QoqrUr
ZmNQlBBxUZhzBnZ3gieZtyceK50rT0JhPXudRPCFl1AUuN3uXhs/9haS1GRjwrJN
0pV7Bu3XsEQGeidwhPNwo+CwGoj0ME8WNcpQOpyHSAfqdXMDIOKcudAcgpgc4hU6
cJVlJwHGCFgc+BvgGQsJ1BueHLIo+b1F2CAG4PMUqONIG41l7cjAG4GXY2B/03kJ
VE4tHZJ00WhOz6GEX6YjyWV2PFoR7Kqx4eWPeUxPx0iv5tn4+rGkb3dESfz/peWz
tdHC5nDU33Pq0ZFghqlo1KWUw+YCMkTvQFxdaV+RrRsU5dJ4RfyYjEknNWjlYLJ5
bJ/h8AtH7cRebtnW9TvSGQ==
`protect END_PROTECTED
