`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c/q2SzqM8vWcNa7cnBhZMVJ5I93wCCNw6RZ/XbvBggq/OoVOc/+oxvFd2gV3t0TQ
fo4ZW2/iVV1AS7Y3z9xsWdpjSRxo27lFqaFN/gAaJUR025gnOC10aRR9O7ZshrYa
KPTDuf+9q1cMcG9IGFrODppQFaQTmkqPI9vELlq2iTg3Skq13dM8eM6Xy74LI6rR
3HZYHo+t8WoMKK27El1FBvBwvTB5CLg90sFY1i+HXVvtIr/cIsz19UdFD2fEvxzF
IVwAVHdcEDE621cfOI+ufavHc2G+DV6GwImyce5gpQgPoRi0Pjp29nzbEpBSlopS
HAgSVRMCEj7D5lfTLOVf8w==
`protect END_PROTECTED
