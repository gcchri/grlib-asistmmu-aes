`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nkOc/acytMPUc2gZNf6e6ki9i9OHTjrzdDe5MlVwajSKMdGFWD/Zwk8Hq/M7tzAH
d5eZVKZlhnL3E+2M4y79fOfffuapjD4f/oipo4EHOX+NGJ3DrQ6+Df+2AZjDSM3y
IvllEAXOdWu69A0/IcRZozmBrvGWt1xWzC1TUR1Wzz61qbP9FOFbN4oO6zUC78N2
qPG7w5liGunWEWGaEZMjfng3iaXsX8fy9HwjQQ5ICG4QDSX9iMdCjCByFCzuqTQE
t+VVUnq9hoxR0nHVDpxzt1qzYRunwxZQDZ3cYyyRFGi/UdoAv4QqsZ974QUjhSh2
PTQoJsiBh+r9JVNsyNcgqKDwe5WSUaj9QrkqLea8uNxTzBzrxELevjJTQ0AS+FrO
BS6oK/NJDuWNgE91iUatMTd6QsRgaxQh0mtKpYF6OS/4WW7riZzvUUEnhgB3Pr5S
yP/hCoEQr2mMmn3jTf64b7A6/hHEFDyXzYFcepQaeLuuC64/8eBVyK6C4uMxTMok
VQ98wtpUfV9dM0Ew3d2BYQLB9/O6lERDD7YRKRvbwBKROtFtxJ2YSs4RK1efPnJo
iYUDVVRPMRDAFcp/Vyk6wFb9w0YeE1oRPgdXiO7YoLegRLKoi9puy1G4oxdYRxty
fKSItKUEvcqn4Vh0wJzaLVI75wNkMqNCK15LlvvEmH8ez1t3Xn28yGgB8ugNPzXP
GpcMJrGvya2bVdyukC9K2kjpDRsA63ERcyoPRtIiHq5fQzSL6rBBHE9/IHgDVMX2
OvaR/U0F6JJPUSOg39zfaCBsO+s5p60rOeWJoMOgnJB5TG5mZtjtl3BjAX4e1h2q
pIwLmw+N1GfUJPXT8zdUKAdZUGovn0KQz3ZKt70xQqxJJ2a22OkFNGsiM6dRsWEY
W0DlZ7qPBWupJVQ99TB1rw==
`protect END_PROTECTED
