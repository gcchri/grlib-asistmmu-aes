`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35v1dHDIV5aAysVnovTiadinq6LtoD3FthsVb3Zcd4GsUuHIOEWf4tXLkapiDjfK
Bc1peXg1dnwYbnxTERdTnr/7NsxpC3fLLzrxsOLPRfuktzbm7WEzzUTryjnT8eTz
otD5F0hiYnnl+TbCDrb4qvZH1rxdGDJtgzPk8zzk+P3EHNNhRXUDQtxP4+7rQemz
/Lqr4n53B+B6BJ8TJ31TkK8gO5yY/CfZRPi2pZ5ltshnEs1gt7YupfIzX9sZEVrN
IeTXPT1lI5fzLuzYtbNUtWfnuIwF5qeC4NIYEdg9LsdPTNeU59KcssFAierzjP56
eQ9rnyQLHbqunY87CCLVlN14Ji6wC37iPuly2IrmbfE7ClSSjWW3UK4MxokYd65j
Cg0nBs3LHEc88fqvnwaNGKX5XUXv26tOQ7sKi8i34n6MCI3FfCFL6lij3aK7F7r0
Wt5z9vZSLNCkzCA+5Uubxyt3K8saLvcmeeG9VO60KaRq85Gn2rFV4yQzEJEqw+2T
D1zM+wOiCqtNaLdAsmSwkewmmFS+0Ihsadr90X1s1nU1+tluSdl0mpQFhE82T6Y/
ITyAQEfq3mlCz3RFBW1CFPxVRqMgkc/FRWhcqHD2RoBjlKIMmTm/RaX+ptcocm6V
vZVT6kAqUH9C8nB+i0hsQG/7QVFbLPNBMsTkGcMPnHsYn7eHx0KP59KBEISF2tlF
jPpjzNMsJiIkvrFv7JG0a34o8ggEcGsfbDLSg20FXQWVoY/A66M1FnrSSyD735jZ
PC4/aLvhd2LzJ3NHJh456bJ2HDbfP2bz85RcUPr6caKs6yLCA3xdOb/V1+mssqzV
SXzn0LYBDJ+GNC3dlodGnMslc+frrD+w4phRj6g1P3jFb2urSENqYn64NbpqnT9B
ZycCN5/hT9q02t30eKH3PCpIiBBJTvnxzLjdhwsxkCiApbSBUljrVTsfDotjbf9g
rltMz4wUolb7UF2PW8IE1X34JsuxAyjER1cyoZoC6uvBhDmZjXNI/uPDh8APsKpD
h+/p9n7bf6+49GlZGUn06sQwwZzh9P3HQDtNCTlhadzsEfnRCeH2pSeAQgN+rW8+
JVN8dgtI6WRc/9Nh8lB9YcgQjfWp7Zdwu6AYfczfQ4fMUAbgulNzjAL9ZJvNNar6
XCXL+xWDx59wt26WDtqXmoQ4I4AL2jRMoQ0CSyNpFIWeM0YRq8TqJnzYX6ALRPDh
7V9s0cdePDMWDCqAdCl93UOVzNgo1yBGIC1OvKYsflLKrEu6PB9hZAUCEc8qrzb5
qoO4VdxhW46jAkzo3OmikF+L+olCB32LrxQ8zHDThlHK3lBOpNee04JaCmVtSpka
fy/k9EaS0h+OgCyizp6PiYtNsAuUTVtSppBwEI1lh8kVDytoWT2N3hw9TW+6cWjO
SIAWzCiSYXrUQb1R2No/u88TnB8I8Ff6i7WMyx/SGswzJNBkBc4awpy1xjgpKgry
x0Q/MTp0vVEC1/ovuz5cdwmqOBFNGYu17XcWQpHwzg+AahQM6YnBHuxNki+xb6LV
AUvIff+bdPYbwzHXKe8NhyfXtnFtMjI3uXg15mPX62ilChUwe1gnN/mHmEk/uq/p
J4OZDofCH45v7Pu3p7BF/Hu4TTYKPwFiPi+oZHtkCxyBnFutq1vrxeoJ6nBmb/a8
zkLd/uqPX4DiP/Kgn2i2s6Fx/ENWzksTiZL1NObgjPCZsvCrVMEgB4TZ7lylHy3/
7kroLH0/jtEJoODy/lAW9wgt4Ywdin7IWqSxs0shgvtfPOYYdX/X8e/smIg60N85
3Rw/N+vTR6ynZ87yOgKCIDiQxNons5bJkxscmJqnpDwauwWgwOKR0x7KhLchdKPg
WxGd3kfg4RBM+7MO4sBmtBZ/6XWNfTF1QDCAtGJMb+ZorBAJ0HW8oAVzuoyQSGBj
nl12rhz8y5VV0vuIbFulan3hd1zakoNyj8UHtJlXwF/yzOXSTdqdHkTMUV4ydeDR
47RZNPVWg4iHnEGsXKP5l0cngs2LKaH+BaOfTmr4cae+qb+bDBxWsrsgeKXvsgwd
tc+xJHtF2mQeJACfF7hAwumwKDgcbC1UpH/H6bek1pbBK8Jwk5gk0aet2iZ1fQ8g
a6c2b83VFChMEzgI3kAuB9Ml1OGY/urlmptUwb7iJvCGl2qRlQM9gFOAVRiQ88Dg
zw2gL/lwMMNk2AJd6dK2lIIrM5nBNpWBRhbiKEmmHuee/nhZAXNaoeFMCMXBuvBi
LnQWdy9Rfq8rWyBVdvJvMz8kzf52M9cqN2h56o4F3RrEuG1hmL4Pz/bTfdgTGwys
e80k4GOmOL9b9qE6XgdUoVvxigBJLGHwgao0Fi6dFXtzyNibcpD6laI1VS0Iue01
CPXJSRmbLCB4VEb1SttzWJpivJ91zLoHs2z1rTk8oK+q4SnEiYkpjGxOSPEpSqif
Q0Q0Lwu8fsVZqvxfDJoS1TwEsY7UYRJ90HFFAIqhGsNwpAqZS3FbpS3yTtSbDOt6
+aBDwN7nKoQsYogiaq4Ko32WJCzEZqHJ2be2C73Fqh+Xjdk/YwXsGNWkiJsydA3C
VliCHW6cBUdn27w9fYN76szLR86Z4nBSyZU9Gy2L7P+HOkM1yGomAuH5gVyeBuR3
`protect END_PROTECTED
