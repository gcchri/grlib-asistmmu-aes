`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Zi4UdH3fHrQXcxCM5WjL8JwkNxU892SW8lal1DsbEBHD13Owv0ujtEhdC6ZhTFs
bf24JaPkrGNANDKVxXad5NiQu559DbyElfg9bzZbPZe2FSybiRmuttY51Xv3t05k
tTCEw8M8xxCMHq/8hLgyg5JjpIuaacH4Q60FIctu+SEqZ/m0eXT3M1nFR0hE0bDd
gqiRvYFgBLemOcn6LvIQKsRhERPW/QNYtKKLahwX14/dK5i3cPR4B5IQYDh2Yw/s
UYDjm4UQdLaJjIE+wdL21LgyF6hEmuJPczGfMLFgGCS0Bth2gV23KApoNh9GLCej
9p9CI3nPhR9UIB9UufHIiQMxAPsdcdmzkqLXI8PlCohk4E+P4gD/GZgkeX1v3/6S
WsNL/f/Jys/XrzmK54SalbsatU8uZ8MNjBaI8gjzqRBbbe8uRWChiDbf6nGILS57
LlZzLvBySc0BKYZ0W7UcylGSktdHRsO0Upbl20FKukhgfXkeiLFMbbZTiI6UiMc/
J21nK5nOcdgF2rl0Lph60hAF4joBxk3rx3qSmFnGeNn1obaYgJPVH0vJSYKIAb1e
EfNe/ziUhFyW1jGSQyk1RfpKIs++J6Tossiz+LRb32MD7a/tS/GFlFXEZM+1HaOu
x7FDYIXAJnQSzjHAQXFpRGKK0UbBPAgd7d5UH0bUOwhmSLYlOXfI0BoA1mEFlY7V
Lm0ormuWHDCWxWTqWCGiNcEfdJ67rwFw9s41GbJZAP0MmC7883XOCrvhv+c6H30B
u1UtxTjiSHP6Qxtm5SJWQ44n/9QABIeS5LzkR1P0xJFh4WL2U9BK5/9I8T9YgLAW
D1kKvNcKjBYZyKF76Yo5cA==
`protect END_PROTECTED
