`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bdy+Tyxvn3Er8k1tY22ht9ytDRGfje3CHlki4u1PD+9Y+McIi2VZDW3rqbR8dPDE
notupG2JYM1FAilokXvMPETOxkFWxqCO3kK4PjBjBikV0BqtwPlv7AbgAKoxSuAZ
Ggy7E09gwKOHULrkO4r0pO3hyLRqO+KFav+kedvUJp/FEiPHNqdpYTBB3XM5Pe7Z
3omusEYkAFk4BRBrL8mxXiX4bHGxJYsw0rfKsTao5cO5JZZ0OvKNXBvEGR2xEGIn
ltKcATGCE4GOiYAEa37t2GEfUsv7p/LZEeBC8+AjDuc38aODjGl28aTM2a8MNamE
rbhdLIYztv8GVZ0Pu2Fef4QiXdTw+Xc92w5Kea5viynlPfO31hfBTvFDLdNGo36p
QAor9O/YsPV5yQCVSlszvg==
`protect END_PROTECTED
