`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uF7RrmvH4lUtBUlxbafbzgapbzggNi5G45A5bVPPXPf9i702V5nt6GTAXSzqa4Gc
7IGk/pdrRYnEXN50eOyNhsrnCgoBpuYVLaBI8HB/PhbVyB7j6jPADuJG2vfwtRjJ
4Q88uZ5WAzWROXvjbgoWthAREVODT9w3m2lyXSVIfgX8uqe194lr5PNVrmv2pse7
cDqRnLXLXcfI3ooSFUzOX2I/XAbAJ/YrHALbvjG5iPJnTVf+RHW0HNqfQy9qFAtJ
uRhjdi0UE29WkfBWKZjObWnjOWHTXgLOzjNf+PU061UTNZGZg9ehQ6+3rVrtckNz
8l8sL8SL9YIK3YZRfTzm3VjCt9JTPPiNGUovWRS5ZTXjT2PEBsmeNnD9RaEkq0hw
`protect END_PROTECTED
