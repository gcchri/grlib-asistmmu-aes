`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eclZEC8pYCAPV1zln1eh/mFC0f44xThH6tBsHmyOsGJ6vd7kW9dEv/igT1Qezq8W
pTIkKbBG/03KagxFI36I/ZoMQtfA7W0DNJrlSZyfr6E+Qo/2YZh9iVqdGwpvVhDe
xd6yUvOeFkmQkld3yFWtJi4/x21I44Wfdr1/z9qkuXQEO2t2hFBlD0u4Y1tt41qL
1pko0L9/dDce3zHNMIQ0u3qgD8vW2G6CKstoQsn7TGoWVDTUkKl2kGTpucHKfaut
TladpKjMOpVxTNNMsgLWgezqn2Km+jgGJ9uDAB3BbmJEHIRlkHbY0yAtrzoBybT7
CMO1Jv4gnnWAF1BvOy7FnQ==
`protect END_PROTECTED
