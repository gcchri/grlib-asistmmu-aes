`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JkG/b7VKGU5MKVAJLtz/IOi6BuSo9fHU1A9Vq8poE2ZfkVeBw+TP1rnX5Ep7rdN
6LJvMQpkhFh+jXSkynM0CVKYyVe8gjuIReYmQBbCRugRwrkyyrZdWy/BTnWO+7Iy
gpDxx/cNMuoPmZH+bz4yd4fQVtjfM9c4yXMcUkw3BxEUrFFrhoN1RH6jauzwWXcw
kc2jzYLHlHf7psi2lqKjyKlB8RjLW7aUURv1pfi68JrExE3dAq6STlEV2aCNNgOB
sp7Yu3fdJ9OtUnxu1tDZpdjKk3FfQ5a0pacTLuxflnEFTRiCcuRyOmfaq71nMNiS
zuahaBOmxWHYNmyHxLQ7rVztkSdOVAKIqG85XZrIqqFSquudoOmuxtgIaJPdf2C5
fottEKOeL0Zix2DJudYE70c5ftGPFgbHqyPRjvRZltrRhcv2nKXt7MoQZj+48LqY
1AyaJY/XLGO045RioOFNoKAjY/D9LjlvOu+tM+hjym0ZCKiULcX6GWP8ajrsKfZ6
3KwT+ivthZmKkKma81Bxk7K8zeCMWswrCo/htoqbvKfFaY0rgm25dcNPE599DT5W
m3NJM4LMt/nGDdU3fhtDOEl7ncVS777KnnVPEn2oBvSwgHH6FhqbV6zMKxKp8kbl
nJWZ8B8bx5lPCjnuw3bCmg3w+Tq856BJdmhqqQiJYuG2okORwFdvtLlFPGxJTi32
5TGpAa4boDJzUSSZ6HeMJlCe5b7xe1ivtU5eHM3jDQuAXgMwNOkGSTXGy3dIVIJT
86pjRvG43HL4WXqiX4LHiQ==
`protect END_PROTECTED
