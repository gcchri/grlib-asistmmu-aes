`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7tXaB8b0XTncBCn7rq/cdWttXk4LUYtsdXjewYP0OeGz/R9mB8gsU+Neplshxwh+
lm9AYW5vyLss0iBCt3sZtBJKcuwwdzb1a4dy9odw8E8eTGn8kGU1fg/AGt5CkAz1
u5OnT7KMv4EjGDGjdJJZw26smX03ylavLLlyZ3V/23WUmdBU8IDv360RPMWg7/as
1mTzQZjMh2FTTGwUC67B2WclX1SP8RAUwSPnalpkfjWwvS8Vs7M10B2hFw0XE7Au
1aQvkaCQGgajYrz6DKOnca33TCqtGKECQNro9vubFvnrm28fvx/5/3wFhMPZ7ZvU
W9osw1WXHXNh0BvoB/NKow==
`protect END_PROTECTED
