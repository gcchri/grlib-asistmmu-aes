`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SPZ6p4tbdi0d5uH+axTdYb4Zp4Q9YPoBopzXLVTDdFtphjXSx3dw0LvmD6wWhmwI
+o0oneHQXm/GOYHGO7cJN+edniSzsTaMFMvBDB9ly623SjC3euCnGM/0Ja4M8X2q
pGvhGe0si2siYQHbBIiCfR/LghFerg8t9gaZnYnXSF656atGwfg+KyeQqg4Tc93l
W4NoETNOBvQ4wbejiSb0ZOI4mxyhFLVWtV7B8YdWT7cEDypLXp7tjptxAbckoTGz
5w9MTJx3AhqFWh8X43XJKGUpcLyY3dgAbjN1qV7NTbcQ57Nolh4xGUpRwQnKhukF
sSFl5gsyrvYAjBIvfabVhGqj0DpbnzgrUXt0ng1WWb37Abs/dg0yVidaqUyB9+3S
9CiGsAaNNnDPX671R6GLLkysrkOd53d3gfbWJHUKR1lRjeHLWyJXjWBJzyhrQEnv
sXutWnZEObUPQvAJXq3SLW9HAh+BxdCgvXX3mC4Z8skcKgWUK9z9NviIQ40SZZRt
`protect END_PROTECTED
