`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eYbtA2qrJj+zbz0DvychckHBZ7FSaExXQWVOk1/ln7C7s3FAgT9MjO0E4UsyyPSN
+uhPY+IS4sVBIdXUMrA5MKbWX0+R3+LBr5OmFyGCDpG6Wn8CLp617xW7pYgs2F0C
t7Yg53qRgCwwbAXsKsPzaD5oY5hxC0A6WxXA6lBoJNSx2DumzJYRzX4VGHMnKvmy
cjlEAuc4wlAxjB8f+uGwK2iZGUsH+icOl4dFD8172cwMEYkgNk139NtwWx2J6HQ6
xyHGUafoB9V9gpvDHQmBfQpeeeiwF2V5FA4gEKAQ76YRN3NC0iWQXMTwcD35ArXc
8EwCiQea2avWXYh7dVt3krgZ5TXaILtIbVfpRCPnFeACGPu/HVWRdh48Io/m1+E8
BKac+FHPWb3qDhd0yMqJITOVSrwqWS3itQUcAFe8PUI=
`protect END_PROTECTED
