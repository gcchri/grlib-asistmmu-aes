`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uuj4VWVuel/0+Q0l5WR+jZxFKr2zPCBfyREQNtCNodkfD247jtglnCj17CyigMIO
Edr4qzKMJRXKgAIcrTAxubDlBikoV8Qpac9oKpWqrDw42bG45564dlmUL0KH2pCD
WkF5wqIlQgvnTzQn6iKJDrXGE8cQ6qvca7XVEg/TxncSZ3PHRa+Z92EzcNbI3PFk
TxKRf+1rJxqLeEcod3znD8DJp/QVJYAt+hEdFSybElL4pdCyoW9Ti8vLF+jUd1r4
Uj32NVEgviU0kGTELfvTih87dx00gv/jwkjKiyDHA8FLxcHsCvf9sl43/FDXbS1d
+TQkM8DIafg9UGq3lFQcGa458Kj1Ar8w92Pg86LBXDdBhdt0MrxQaKTZT6+tpGzh
DanIf4o0eRY3t3sd419B1gGlHZEaRGjVkk5/MxzeVvzRAcGnBiJduGcpF2LcrBlP
K3TSbTJjrvBjAlkW3+UGPiV2izqbHn1xCIisDsJQDhs0A/7qQ4yk9a9LwkIIuh7Q
fzYmNnzj07XAkA7Mw1EwGZg5ZPcVV86P9Kiqc/lwUfnHwjLnOXR3dn8d+ieZkjYC
vkDRCbOeLyCirl7FyFuCSJAQpX4PTDVYuYHuW/wVMPpDxG82pefMSUn2yJ38Pmhp
O84S5LYP5FvJLj0Q84lERAnMgRxyVlCemsNfBlACeLJoJNS3rBXEPJO9uzCEZQk5
5/nfYQHclw7buUni0+0vqG/JVkjioSi15tcyoU4hSnxn6s2m/9EG56wzrug58u9e
KfngWssJh5/OnVHjQJC0AnlPvqSXkCskqH/J98gsoUzu0YvbAh9c+2mKxfIA0uvy
Rp/aNRrnFFQdAaHQap2aRuaPXLAUDwjkSrx1sZzJTHwCSyFZrnL2qdbKhqxCIAg4
UtM8NTFPCPMiYE0h+BDktMPtCl6rZE9sSoxtBV26M3SRpanKQTR99hpY7D/zjsTT
dC5nnaS7l6O+XZFQm9WNKAm77jdxQb1UIG4igxXqQ6mphjBFWkcqKpYM3VtoqdHm
NE69OAhJS/MOfaCXUhhScap8u8zXZ3j0fJl1vr/MAAlGyBs7Uv6+OageSe3zD87Z
RjwlsOrjq3t7xpO+hBYgMpKT+GVl6MchR8UBH1uvoc05OHSAYnjNBuHjIMPINQSW
WTtCiX8fXs0KLs2i/wjZWUPs7uqu0kmUayvTO/eed1p0oLKwcZop4+sF/WzYdJbZ
Osb6zfwoSAW8tRsBhEoSwCVgRxoO6TjxVicWDf/PGWO4Fp1mQKCB3XqFECjd3Z4A
jqwftShICnZ+4CeGx+1w3i67THHb0A7EwA5bW2w10avHoHwvuU73IFmSr+I/o8rh
`protect END_PROTECTED
