`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4QuN6JoC1ZTcMAVfv64GXhe8MzSrDHi4JNU9ZzKElIsfvd4ZfbZiOvd1s22Pqurd
PZF3Km6ZJ0SKHsECXt6xP57MXoJnpvhMMfsoa1ycT7k+2NiFNrrEwpQZG9aGHZhB
1v94nPzAVQsMbhj6VySr2jalyMTxiCRKxQ17UuDU/LIrZGWKBg6oQ9KuhYiTJRNZ
rblJe8BBm5dzsJ3D3g+xIRo4t7js72rIvz9eC6GKdlui+zlwac+0jft4dIhIWdb8
qTEhBu/+DQM5sCWqUw2SdR5tnaiPcJXqweiGQWOEIYlNDiQVsXxqFMXMp0S7kSLp
YlUtoIdlcTaNrRrJALpqsXHVs6t6r8EA4br0sEMNIlwJDLlHaRsAL1Y1VNEsVKsA
LJG/UnlvV0Mdf0WJAOCMZdv+HqOk6JT48VfCVWsVDmcgfgu3bOTkxZO0RSyqHTA9
QSzwir6wTavXEn7RFs1wjdUFflK/r/sJr/2L8v0i74JurPzrOT1KOXpdXWBO2iTA
VJ8Uf8DLnMEeDhLr6z9b2agwTijZL4rwNR6D1pOsBNj+MWi3+xTJ6g4IwkHISFsV
HCoEgj/f7WbAlgU6VZIxtlf0XmQryS54Sm1z0n7/uNTn7w8yBA8CsPRQbRAm9njh
R/T+jnf0bGcirit58RuU8SDsaWP5FJRFTYTR1prj4JELF5vJuPfKUXM6oPV666+l
pVQ96+mZdioCvsmmpVQNOjLZPKBjg8fEhp90/NG8pfg7C6mlaqmaEwD8qLdjucye
0KgwBbr84YpoyHL5fo7vo0YPPCCMzkuQFQVyf23M+iMV3m3aOfM16sXHR7v/J6Fe
61mYxydWFSSjNpRHhkgkBUoC9Wdu95od6d6Jlf3YS0XNaIkamTFKzlGWsuZveKrc
hn72ZJXG0ul3KDLtWStH0BhlySqxWgitZLi1f8LvIgNk6uyC7wLxBCN+5+qaL4eI
4ExlNNuSDmofGF4IE5kQcz8dWqhvCRrTzfU1D7XtTrtsx3y04Jbq1Yf+eg5F2GQN
/18wenh2Up+Wl8ZoBa+sLFhUm7nC818nkOqtTZsmP4t/cXKHoqY/9d/p+hfELxry
vx0POhoanmD98CQ6uKhbGDfZqI5M3mC6Yj8Rp8CulJiQDCmWma226qxp734RC9Y1
HNECpqSarEQjpHhWbL78IvKT8TZZrizC2ARyoGg6dYoHeQpQFAwxbEwy3Jwe2+de
eiUorray34AJ56QC+ASLPyrVE5ZWg/GTTldf1hI2zd8d6dWuB7Unj+yQvTqxqb9A
+h/kZy0BQmBFrVfQ+F80pLDLmSxWq1GjRZNEWSBEN+Q=
`protect END_PROTECTED
