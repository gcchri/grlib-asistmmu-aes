`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDqFLfV/3afX9gDpywQurvEZ6R4Y9Mj+kLTBgyI600QyhZ3LM/Vwd0STwn22CFvi
nTSZAKSBrmeZ15XUNFNpFWtnw+2HNUzu8j66+DWp1SjeubIZPANE+YJwhTs60EcV
hNlMEgWIJdCqvO8mFnDLEAVWQnLkYqWBFYWpgT59LbrR82G6ZfyByctS4AeHo7m8
n/ij5Xj3wEbb3FeTh0kPSxL674ZPX5jdKJju1hDOv6599CqsXWZq6Q54Qtn3SwI6
vttl6Kq7qh6S0nDL2rl9fdrsVaBYMRtKXdtbDg8EUTs8i46sypGYnt9kepWJoXXY
hyoJzsxE0O/HrLwlmfLYx4zfV5K/yuvO4ITHgXGdk9ZjMGdt36gyYfxuTVuTxtwX
CXkCrjvp/JAM4hxyYQxiUAC/rkOQ7Qg83UtWW1vJa5Rh1p+ob1rNZ7V26n27419J
1xMdodsDRqMcP/tBBtsDedEVrMW3mJnZN10jYgwWQndIvF6T1e1in/hUz1yhJ5vu
SwcM4enwTliuHZrjjsRADxioG7F94dkV1DwiaFhBF85LeQNl4QzPHOzCUN5fYRE2
h0q5eDUMuzIH8B4Ihmdg0MH68g0MA4Pk+bwnPFitwBKtFRfxbFGN++GSELKcoxzC
KzXCmf15d8AStp2fvd3ynylu1T1MxUBsPNQ/FSeEisTK4C0kTqUnrIDUB/KeqB0Y
04aduiivIBePjwg9B6fVdEmW2Zf9mdnpBkv1YloeePWdnHEgpoaCNIABYvockrxy
DCtZuvzz1tIwI+xVc77QxYpaK8Welk4eyTlLO2N84jmzZVpzCIiFMvSwA3M7chZI
pgjIPyp3TRGpoA3l7gzsTRLha+wufVIbb3EN2hHuU0q9gWwFx4CgJctZJXFdsT/H
svnUG7QbWkVnAQPh1PKKW7FB6Keu0da61GlgoUTnMKc8yvOXKuHJkQVVOT2UgTB9
aYoa4IbOIpvWNaI8sujT9ib3LCBOceAumDSe9uFMnxvaeP8JIKz77AvdfwsQbTVt
x0dLckahipqRqnmv9HAYCZKUpoa2AKpL1l2UxvPCQUfDUaCgPcCpuzKrHP4CSxBe
oBiueSk+zhkXdS/I96ycTH21f3IeE/lSXBn6413Rf+SSLneNz0KrY90NqrMusMFq
mrfbu0Aavj6Ia9Uu/t/EYovnZhxvoieHCXuc6yhZUZpL5hjSrW7jpgirQITmb+XS
DXBpw9RwR5TR5rkPAQzjwHGGetAiUUFmTJ4OnbREsVB6DZb76VtKnPJ04JcMHKxU
V24edxwv72l/GcLoq0R9kdiAhjTuohEJRMtX9NNmM5DGPemZ0/4hR6JgwQAjX4Vr
u0vWkw8i6Iv5egQpbCg3m2wXGtPBDalIpjs/yEZ4MPM9VwLa3Z0FBTxgPgcDkKFn
A7wOuWoOjQHLSsW5xDXGhKgzbCYpaRv9Jyd0Tp51Jtx1uITYjn+hJd9pEjLUpZRs
6d/ylLAPY7iT2/WJd+gvSYk7NiLpJJrJDEDlZlOndMNhYSpRWUzf6eDFRvuOCXOQ
xB3ZbTWq+S0kU5SGVGnX6nR+6FHZCNo7AGmYa+GjcqjpDgpGvhqPT2i+o73mbLtc
EktkZk0Z5O0L5gmVK7x3WyGLgS6l+4BarX3PKa+C2tAfjo+FHQhB4VGKgQG2LKUF
2GuYO/zk3b5+Nv3BNHhoXsq0ANahmJslIRLg3bRQ+jwwygXIMGL/LI9W9ypq2k0u
F2Y1Ukz7lKyH7MgdatUdQQWHSy3DAZDCaKxHQeRxz/cN5Npj6SWWL38LIVm5Gaq8
BKoPdW3e+EAajuEiHYcVkmgcrYuVMpF1VfkF7oqEMVU=
`protect END_PROTECTED
