`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lk6PehgWekGVhz/gDi3seAUd1qdF6EaApGsGrTaE4H/FeVzOoBdeozlmbyf9b9Wx
BZ4j+qVxQtflBkGwW5zHZILnXf2nFyFNxHn3yGXDpLNInjOg37NIoE4WAzD8GJeo
RLcwO1MBJM9Qa4pZZAcmiWLSiWMWj/7gFjwzcQIilHNie6UGCI5DU4/bUcfWBCEY
zOoZTZGC0S381B38v016zbPAc57QSIJHIWKB2NnEJhxonp4KwEmXx4sO04/B/MQM
UvbLkF5BgftoX4B4ihu87aq4G+Vm6bdJ5fBdaOBJw2c9ZdfbKUcyWrQ0fiAo+uUe
PRErcNIxUkOMCuEp4ChnRRr5y2E5EkROCQT34vuSd6GZwNvWhWIGR8Mbhq1GPSir
vZVjAQmN77zP4PT8rPnQ/aXTJnBKLZk0fSKWd8uy02bt092zpTIPHeo7zEvmNl6i
R78u/QDSLvO9x4qRQb7geFFL/H0gRzgSeMza5ocN+sIPMeSRlqIFh7IDeHCLJVWt
O044NWyIj1SIxMh01NJKtimy4ftUBrTGPohSm5jkjvyc8ok2tO5hYUqV3eGIV4A0
lcKCRi51qZL2EdpzYZ8xa8PIsnozs7N7k0hDSF8wJ2f1uQXbjfp+YxjHv3yaKmdX
fwcO8CCJj4/RYyNWC40OiwRb+gs6oSKgws9NCBZQaMlZr2Q4lrBCuxLla357ndia
GwUbtMQqrYu2NFUJqqQB0Q==
`protect END_PROTECTED
