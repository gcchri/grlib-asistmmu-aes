`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3gy2PT+bAQatoenl1UEKp77bIKQgqSmnhRLq7i9+dNPCiRmluTaKsQMeusvan3QN
k7ENKy81i59ND7s0hv+Z0QcqrB44WDjgrP1RDPu6RDxtf3EfDD8OzGrKprQK9l8w
MmP4niXeOMcvOzTFIdXr+XL/H4ZF3CAusgdFx4p/dSzBr3wIfGBo7lfho7SjckjT
DXgcEIsa2kEkoV/rbEHZiYgYH55COl1erut0pSao9Gtj70L4EdDNnsMwegAuqarS
dW74qWis0yZnMebHt7W8GIMXcUlwCrZvgINVx+guXGZ7O2uKdIDguxAG5y3nyQXB
sexx8EmrgzSO7ANDlI1fCeO1lEEqXLlEvinnvRHtDj+g8+EatnWZcP21j5WCbB+p
22++M9Vo8F0PxAWPcOxzW7L+eKnLE77RvYHSjJcOGWAbauly0GfSyaeMG1A992EQ
LMtfuVGpV3hajX5XuvCf/gHXa+1/2NhD+IlI0MafjzQfrW9O0oOuWqyr2MvUUJ55
dLVjjOl4/XhozvI3apb8mKrqKTw+log6YfT+72lsrr5TadXx6LRJ21bdCKCmQsoH
RqycBPg0zYntGNEVfzU6zULb2TDl5Pq9nYBptIj3ZUOMZkgnf8PPjVDymfE2qg0U
K1d1E4LNJuyd+reCBoLbkR9xyq2eZTerkxZGLFmaGPDLsXhChbb/OJ/up7npHOkx
mDHMhM4VOik9+5ngf/7J2Wqhdr1kCc3CddX5yJ3UF+2httgVwTx7Gz3Iwb1WyTaE
Fuc6JCC0FCU3I0zQE/QVwtscpJKCKsNPPZucj1sY5dELF9ax+TbUqEmK0Kd4v6QI
Lt0thtbfN/hkuydbHKv94vk2Ood0bj+2bvRhinhS5W4v/bpWTS6vaw/KF15co2qE
C3S1KPhAXUISchGRC56FZp57lFoOTWhf2aGA8ofD+WdiKLZYSRjsuAjb6aj0+WkH
Nx4gcNQ8uaK69PfSkKmSmyEtfxtgBDh23TwlB+E7tUK8oO4XWGZzf1OfLu4ZfNyO
OqZ1tSgBPlTLQemxZKt2f1+bDSSsn+gfb43eBbLYXcBkvQZZ+8WUjSP5EPJ2mm6J
DYkwawXfAUapaSVRVEYQQiIf8xuOl/RvMymS2HMRXj61UzWL591vpz93M79rj17n
+LlbF3LZ7u68jw+J8aR0h7dqlao/DEoEKsLTVASb1W/KKh7ZS7pYhMpr4Un/3cS0
bg58Pz3eXIKaRw/A18av+6UrprdgZcgkUtweL2gB1ZYb+iM+zjyzU5nnNMoUUk7+
rV8RPb0s1aFeNzzCXNlkhU/d9iRIyIbNxffAysK2HIAioIbqWIzDSjc7niD2TIuI
epmCaYOL9/s/ItuAQEaP5ZjzScxXO6dh0ODMl3SK9b3q/r+8QCaDj4Mxakwgh0kX
7DmQAoCcRtSmdCFMHUqNXK6x9jK+k+WaNO1cj+JJ5vHlyvh3zzSRPNta5WeD0DJ3
RsZVs5uWWDeaotzc8KRYwuyzqqxeugoUfxKX/LHQMKE+IjO/t8GykrJAjM8lclmb
Qn42WB68G56wSjgnctOUMk2OBxKCGuFaTNo3Vq0deK1N4DM/ahdAWNfItpu2+q6E
iok2bilcImb55LCs1/TCJ1hKPCjv7PhL2Vp7PpalDQ7GnAuv/3dqsBAPbMwJ53O8
L6MOnGVNauFm2wX2oGUG2X7PtIdATNEHvX52WF1eDIcmA81CbLyXkmMouOG3ed4N
R+HnrC27nMCieMB++VWZVRYSscmnhSHqIoMorFqBhF8vmEmBH5T2coBlcEwvIj3V
8N03nnq1TY1zjJx1Ugxp9FXJlEdDqYoXmQgKUumny7uB9TuzT5IBm78l5OFn0yrF
s4fpMPayANuk0ULQwLsX4zgsZ+18qRFQ6aDFKk8lsEMWOzJRH96AeKgVFtlQvyII
YNaEU6YqbEgVj3UjJIcWmp6aIcflWR1bB/Mc/Sek8T7DVKU6PO5Dq1joVMKarUaj
cyRM885rhWc7YlXjsGg27ep/bSV/cLTm8AXKAH0Zqf9iARDtj6TpaIKVkDB9expq
fdz/bE1OSf7cxI1lFl/vBzbPXsKlveEz5gCImiljGc5WYbHOdzfiK5H1Xf0WO68X
Rj0Ng5WtVrxBdeBWTVKy49T9U9OrEGK/ZfU2nu+nhuR1TXWyFORMLKznjTXDx656
kVHau/sFb7ZkWmXMwJ+1vqkVjitwDQf9d9vcWnYNpH1Ok6gIOGF4ZWVfkpMRGOXK
TQI0i1Q2zcu3/7HJr3X3ICzFV2X+CzP1xJqOfyr6XtM=
`protect END_PROTECTED
