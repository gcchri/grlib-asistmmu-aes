`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hukt3Hrfko6QkHahiNFly43x7VQMehuzL4Ar0VfMoRV227R49MffyyE3ybudYJdo
HuW60KW1tDjx3+OCtXMNsSwB7mtXiyl7nQIB29wB2nKKxCS/b/++crxAwX4DICu7
0ExjT8QxSg7AATwMMxoemBS40FcC9vbG0EBWCB7MtD4fcxh/+uGMI8J+2FeQmM7w
B4CsnJqvVFmPtdjmJvJTho6vgZpNJVF7fC8mx+ZXekHWB7SXkxT4j1j4WosXvqvr
dV1vSAERB1LewpfIX0vCgOUrwpVweDVprAG02Qp/JuKpF52IOU8DfdIYXf6qZBGW
/d5VD7xHFeY15tLWhxkvIhWbKHqslAkw8di/YymVQLGb7xJ+q9AtP8Neh35GQyRo
JSea8cuWqx5X3R4Dx6K85AckZSsZFuj/a9xfG3CH09A93yp7nHUYj41iQC7Xk6DA
Z0rxVxZxyrGPFKnJxsSQ0cLCqT7L/UHge6Wr0qNvnJky9yDjNeM8WBnupCUYchv0
UhcwyoWKcQQgdFLZsckIZDVVm7u+RXP2SYOan7BKuWNl3FnStk+8X4YWnoLIJcyb
3coZD9QPNrXFRyvbVlFIwOHBCUkO0aA/K3jcoTDxJJdaf6+KYWSR8WOfiNaRUlYx
8AkurBwvsXp3EI8PvyjNq9+PNEw7gYhek2NpMz9KcuXNEKj8ZG1K465k927TTAlr
q854iXT+pQTPi47tFcmP2gQOH0sQmLkHzdKafDk3lQ3JuFij6msg8cfBYFlU1X9r
WqgnC8ZmTpsh80k2t5cYJw==
`protect END_PROTECTED
