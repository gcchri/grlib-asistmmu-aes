`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F8sTAs5SXdkHV7P5np+CBGoPOnucxOoASXqsiE3QbPqE7Ors3K0kdc7gGMVFTsYo
COqv+l9xteWCK/5XaNmuMrcL2xipcDC6I64Ur8l1Ua9buEWXzHECM/UJeI3CYLvl
ZfzW5yUDVwtR20QQYBO9nYdh7fRRolR9Z3IhFaDKtGFWcZJCCCyq65OHFndK0+3y
ugYVYrbviFfVa0HgPRw6ditRjlrzU/eEg8/CSwyFlcDAXISMRVJU27HzMDCu1tt3
bw7WrrhF2nIIgceioP5UAvy02bW35oRXaPk+TIMstSiPjXxarf7VS0Ln35nfli/m
ME1BrIRD1MpmK32oMtEBnld3jQZ5LINfK9yzl/DobbJxqDoIjqsa1e+2kH9iQlfE
wbDFJeQWRWIH+DeZ1AvkPAVqec04VADRv0JZXxmwzEPX8qVsptNsroX2075vrzv/
r+c+c8/oxHEIaAFzsQix7nrZ7d8YIbTwDeL/Lvme4cXsQEnEcsMc4UHMVjbCe6BD
GzzBynINzNUPMH/RDM5JGTBwAAFPUW2lHJBj0j+Z5ZgdX5gscFEm85mrHri4e13d
H0mDUvOiGsDzPc+MfON7ur5rsRCtigO0voyx+kxUQ27qicjFzZ2a9zWyadJ35VLk
USxymMGEM6jphI4utzkWCg==
`protect END_PROTECTED
