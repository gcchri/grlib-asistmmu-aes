`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkmXfv18+Pa9mhX9LsAzzmgQkF2qVYCQxBcwUSJc7kfCmO8orl2b1LHmrVuNyTw8
jdFYDZsjzcOJYEY8okm52/sEOVVePXKN/mV65O2InmG2ptijpYb/5b0Lc5mlboU5
DraIWn1d+a+IBro5rymjYS6ZY+f68jSaH+4w/D113pbcP4X1OJnvC+PwAtrpKUiE
UId0m6vD4Yv9+lGJFdveHCMvc5fMxjoIWLe4FaCmRTmUtNT6f76Ka+aoCryppG5I
2gnkwhn1TUUIlp0StWDkrHJYB9fGFn8UE+NRalqO3nYfDK0IcbxKYsxPGLtEsxO3
KCBMfQ2rHgaZxs91c/gYR26qm/daizurbTP+/Rz6/iezmQuNa1665NSkxAa/Ft6g
pQD9+rt/1JcS49AaGTW7o709M8gYFwskIZGnOVBHbJuIoyBhgWuvrP9uYwUBDeGr
L2U75TasiKXxEO4NrxOj1hS0aZY/NFu8x/5D2fAvFZGCVHECfngGhw1WXRy4DEyf
O0n1GObGOcfBEWb1zZuh1LBdkOx9XZenwnXpFaW4zdSXD1tHIM7deOQS+OERe6uz
MHiemyXLmWwkfFTfRXqaFkq5Vcdbp3mwxHUCX4D09h1CN+zq3Z+llz1vLCjVbHva
Bfs4oNTVEnhp9KB8teF6iQg+E8pFj8Ky2Z/4Yv0PHC89m7Ha2m/cTc5inOIICFGQ
RLS9ILoDKuA9XVYqZlyHZAgN/ME2oLKu264O1Wikf2N4ERF1UFkmnKpa7GFV/nvy
H3Pn4ISMXXkvGvlDpWnjbYX1qVaJymr51MLSCH5hDftp6Xp42G9VLSI1O+b1jVju
yc+wq92QRHk3516jC0M4Z11aXEdGX2jiGCGjMUAdEw63oVbkDJQUnxXBz2nacwMr
0EBIm9LK5dck4xrQmIOJLboL1YmJejS4vT/gq+Y5qQSGkRhCXWsMn0di7zdIyOJx
voWT65Xgw1tj6VEEO0l1stzyjjFeJvV33KbFAu4+KZw+t631o1D95ALKZbr58lOz
7oyl3OCSwP8k3SlEqbvbDBkKnuE6Z2mJd4QJXSMECKAL0DdrdKrtf4LRd2O2PtqH
A/zadSEXlM9OyJMQmy9lEndkwRRUjgaSYQR7oXg2N8D3gc1N7MP3ul57mBfpF0P6
9ZCygWJ5dQwriJzdI37faaQ8+runcZ7PRS8dB611v5EEvVTQyLuR6YskuKVx46Ql
lsJOk+/CVCz4PF4JzIDfvEQOUFODvN3h2uAW3HDEYp1G9z82x8hqYIx2nFPE97xw
hfClVVYm8gw0i/fFNIJO1mhNjEE1xxTLbukyZ0z1rFo1e8SalelAYCaLwUXMZdfZ
DPoFVdU0K8E1tgBROi55atYqfqyigL7m8i5EmIMMgJaJ1G6A39//CrkfljieMdgm
RXW/VobS2A+uW7UCVOEnayv90nXRUFlTY4yOlE54FJWLLoKYDsrF/ee4QbibrP3U
KdjmNHyqezxbOh3YpOg24iXnzqGP9O4MNGVyMcqlytEHH3kJo/8ACvBRkh0mFHeu
zI2rN9U4EYSA3tYrSusl8KMXgTKtO0lA/q/gnIBBH4cqGRHtr4cK2MaY7Lvnroz5
aXMWtNcSK97fVt3RHqd/8WdhA5lTgZvjx34bHY6jG13g6I0qodxVd8mMq5CJ6Vq6
CNKRaAv9z66mgGDrFRstOw==
`protect END_PROTECTED
