`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m4yuFyIRDSOgqUkr6bj8j7d/MOf74HIOAethVyHgbUTFX4GzuosIqLGF0MZ35xPM
6qF4DYMDWCVEMvGGAGTS1rPqKPyj76dcAEt65iEMDRQSBHW2+Tkh9mEVpWcUQAW0
AfTbKhJBspGGVNzEAMKnv5JOlGCLgHpI/WF6/bIyOmnb7yOon0Dp8rKlO9Fb5Exc
X0uUR0ZQOVZpUkLFm5mo1llZv5LnP6cRWiX1ptxv7wV22+jO1hNUnokkXJ4pPwqP
HJVaPkTtRh4GyLxU3woAVJbGf93CkuDIW4vvES3WPH3umigMwdI7AsTwB86qRNPB
injDAHHdS3x7uc5dhWR7p3+8pzeLcGGEu0w2kIcNkZr3jmvN9AhhBf5ircsNFRPf
i7sHjlZZUqrCdnTaSLCBNl1WY2GeTWOmFotmd8PH+bUNqInCVAEuqZJJ5kxYvh3u
sybZqDNvfSGCgHTmaX3Jqu5+WJyW4KPcZOzKhTgS0iS73tYMdFdhEGk94v5tlHNE
haSxbjCKXrXbHmKCvZmUS6OKU99ZyJRodw5SOHIEqeApiw45lhtNu80G8qxjQKhq
uYptXylr1fJNw6uzslxnQipYhhvPutYCwSTWamA1zX7KSE58dXlD4wUNJP/2Eaba
iO1ilsNhinGPwl/gVKH44JS3m19zN6tbMtQ5v/iFAsEfWJOqRs7q2d/7S7+GTkUI
ebfPUXlWYIdeRtHqma0DzgefUDTi483qyb9JRIjfCtbBgcg0AnRQ9hvTWjQoVwVc
2sBSGEVMJit0FsWKlA7A5k8CcEa9D4Lf/89NphzvFBWns00oaIj3e+s2LwyJldIW
01FVxq+uMUccv0hv78tX5cWedqwnLKWzznWvIv9b4FRtP96VIxDJ1VGBKLoy+Szf
3DojjdKQc3sNkQ4KqyJASQ==
`protect END_PROTECTED
