`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jC5FB4+erYRjwWOSqPt3rD5TFbz2RWoMekcI1J4exjw9Ah36diUuwqDjw22tbJhk
/W5asulG0MrpEihapKLiUWpTelv2Pv03UTGa9wQDp7iClOKfF+8JhUVytGIhn9aJ
U4RaZYnR1QGF0ceAB9w9i5cNTXh6J6UWCHYstlLraGNe49NJTRf2ZEWwqzqcmrTX
6eXo8NMG90KNN8pjijB9lX+s9Y01oMoJt5/yQSCVLaZrEe2H599oIRkaBPtLcEmJ
zC12vIt6DR99sTn7OJ+5bxk4DSU8L8fG4RU+QUw+f1QGHCgxrtrTOm6Hpi4ArNF1
VTWRUc48wVdAzLFFmTZcLhfIhOXha+sIW7z/ny+uzKu0bvVymEfQcVmYpDZSnSBU
9TEUf8pfoblQTrYiKPemWHpNfWn/Dti7f43Pj+88FSRXwDjBiYaRYm4dD9pBCImb
ojVgmsPyxX9OW+1RYHXl1P4sFXgmK84cESFslDUVs0gYEwCeZh0MgUX648g/j3NB
1YvP4IBlYqqjk00gNf3F+hpsYHsvG0jy/wbM117hvuSfGA6oM9RHWD6ejcMehlmb
qOAhRK/gIRSkAUrq54J9aQ==
`protect END_PROTECTED
