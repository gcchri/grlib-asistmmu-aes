`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UwRwC5YMpcBfRAEicq5i/tTgUJIErQMFEkcfIBNkHsyHqtOinjfcENLcQ6vMtfnA
gwq3m+skXdYir7XcU/mvwnXxHUUo/U4x9+3LdTy3ngLm8gm+w8hVqXiR7NPYSUTE
d2CbTTV5rpB+M7x77OggEjY2d+0dZHt7Uh4H8LRgPpiRzJH/qJEWEo1FdKGlCqK5
/ns7caKNwT1PCM9oLCb1EzQAUDifqpqFO7+L1jdS0HlkuySGNrFCsu+GXgQFw3DA
mP1nBMG/9f58pNGQOECsuYAy+MIzupZ6e/vu+ko517/ak7lxmut4Ox0nf8/+TKeH
csx2j5Z3ZnKu+PF8NgoDUYKns/hK0Aep+O/TV5+ZYqZeIAHUrock/MCN2pknxTLf
2v2ypFEeJ7MEisMUuW5A/XC/DqwW6PVMFJb5/aSywSdYopH/4W2J5vyM9O/rSp4O
gNLe5/GWLIUdFPh6F48JVPyb3x738KrS5qtzHZ2jOAc5ClZC9xxXCdxqd/8Pv0zS
pfQKJhK/cEadlFKw/eR32Xq04jWIrmxQhjyL9YoZNo9r3T+ElWAt65SFeV8o+V68
jn4CICrFly4eWCnqD5PWoVClPVT6O5MHjAIku+fVSDBagHDcAJsWqVhED/oyBV3E
vzwJO/PdKlUaA212UOTEt5nLF6GxRx91kCCOw2/VOQMVjv64z/WZtncEq28GFta9
xgXgTeYJ7RNbuHi0cTangUQicGbA3szLXqX8tRoTYgL0pfPBa0BBs/ULgZoaJGHY
8Mor3OlTVNfDl6RZOll/hA==
`protect END_PROTECTED
