`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnLijLG/Scf0CCtMia1aZNE2lMbrcwS5lSEc/eszJyLEeRu+2VUPEQ5KdQmxz0+X
fsX+MNnHQDQjZFl4NRsoZXNtq+ZshtApoJEnQnyN8DukYprQxlKBKu3FtRY1z538
+i03MaRmot9wNjMMTZtr9WPJ87FYKrouDJ9U7PyN/ySp1nZekRNR++mvt3ySa8bL
D4Gxy4aMK5E+XI879SFSkmicN8xeOvx4XTDXVR6hbrTEN4s3StM3lZENc+iPMJrk
G3xC/9JKsPWLsaC/UGY2NxzAOCU2iq7EP5ispT4rsfArz9upQ72P20+pqopOjY8N
`protect END_PROTECTED
