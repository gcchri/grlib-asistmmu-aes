`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ztSuy7xKPD0FA0pRDOxbOGE7vARMav2nVcL4N04tNTBsd+hX2jqxWOL+6Qu8oi12
sZQRaYKI56jZF5/uHJXBPa8zsjtNadQR9CjnGvvUd/dsoA413kHqbB6vivMG+iC0
Ux0Kdn1L84U2EyF4eyW6qZn4/Buok67fW0clZ0KuL9hZ3C5ZpaLMuO4r9IPHhUKp
aii5OB/TdRiab+k8kZXgAYSJNorJEo5xhDFAguY6EnFGwS2by659eaQXzfmCpg6n
hbFFZv6snWGzr4OAIBUCl4tur4NQJYt/Ep7m1SSxlR0eAww07y1fWP1IPjQOnINT
WPneX8g1cSiTs9Dp92qjOAfxjJHqth9FZ04sFpCyslL6ogJRwaPOZrJdCrWtdqG7
RUZNoz6ORFX+hPJG3JB6rTZ67fQKVsKNGWi9i+1zDAUsXg8CONFYKw9gRV9SMoAi
YAkX/9nRRGNwUSDkjCQKLvSlmTaP9J0jPrV6YPqskxgApr2dvt89ySGrFcc6S5D9
INuJeBW2LGNA3xAo6MfNVrVhIoo/yCKTdlwKbL0JCFkz0S8IrOqNfawBHbs9DqCc
`protect END_PROTECTED
