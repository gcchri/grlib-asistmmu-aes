`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
otV+GyRg+wR36OrV1umrqO+simQPKLTzEZNoU8lfxYEKxZ/aruMEF/9gdsyoZc9G
1tvMGTh1TgN2PWea/AWFrwApvEs3oQf1hqSuv/a7qNx44wBNZCRiNZriELU0LDIe
OAo5gJ7MP8OccmfQWtAuB94vcbuc3t+8viOyHaUJwKdMiWqe4hQVln2TrWxFLpCy
gkhLls8QIWZwPz8po+/TFNsW0f9SpfdHot1ObpZVLBKvuVcICn055Du/0WgXw5IG
5CiJLe5aKjkniHnmJlbhgqoT3OTwrfHbNA5LbnwrIxmUcA4g46RSbfBZFxt7xlrP
LhKXVbIqh9GkZjSQEcHAUw==
`protect END_PROTECTED
