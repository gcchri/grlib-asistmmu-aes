`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ck3jIoCDir1k2HkYJpglegUUmZhH6tllpxYMg9Ppa+Ezjj5p0XnEzeUQU0b7MA7f
Ks0E7Ta3XyWPJI8zJIC7LR7XI37IOFEEDUP9+AUiJ+ig65Pw2t6Z/BVy52ddg3N3
9qzVkoF4V54U61ooNTuV3HImWzhdbbfntJ6Ss8pGSnbLFotAQW6oZCFNFc99Y38F
R3qOcVCHYdfZk3zrG4fUT0tCbk2hEe27wurn0+gD/1a3BO2JMnaiuRDtOjUhbrj2
EkOvTCNXzYnPUljlq1FVBXkw3ZIlgqrsggBXkrYug3E78aLbxTqXrT7/E+AoJbEV
W1sg582i5S47gPgPKtFTva5fMTU3v8bqdWwvmkXw7+ysTWx7m0eUBxEGIjCS2JRK
qLzd0TGn/5tzCayDkET2j2ss9HT6T2Ak4c0hwW2WhhuKlsiCBP+m5p84j+/jdau+
WYFs56Xbp6ASJI4nalpcIQ==
`protect END_PROTECTED
