`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
say+Xgf+ZQgG6UxDrrxBFjjapNaJ3M0BXehjbxzWp4mZhQSL8jPUOztP/QLjc18B
vlHG/uFNQpk4n0WSqJl51z0xmyXGcWRlyOThuJq/MGHwDzzSwdzLBn7C6Q17+G/c
SYBzqCBMFPVxZPghvfhxAv0wE1yKRxcsmiNF++amnBgTkwyYz3SKKYPTtQmA4xJD
TD/87VfZkd+Iyj7WLF/53NuRyCIx16KEVjahcUsO45RuTmlEr6dwmV/H+xFsjc0L
ihUTAttRB4ge4JFheP8+TGSQyLHrHPS0EzTB0qbBbGv2BirES8IhRLkUlPTaU3pY
bkWOo+6aZzdyM8+G3kY1jZSuzoGKoM7SBqna2MoWm3D4gZePbzkskcu6eJQVDHhw
dNWzw8BQz61C/mNJkuFZwPVycPL57yL41jqpVm474f4=
`protect END_PROTECTED
