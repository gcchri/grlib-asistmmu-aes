`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cjAKRVe9NDbi5kFS3VUJUHptNj9KcQ3eqdYtVG596pEkWIbki3rhf81juyn3lBJP
4HJwTi4mCvVX3Mwrno8ADWoBRpWQmHFNHSbA84bvHoOItNJdwkRTlzlhU7NEN4fp
vq5Y3g2aopmXBE/40TqM5KODd23tPB5zM2MhUTegTHJ43ASd+Crq6f1bOrUoaJ85
QhcPvkY1BPEhhTG6e0iSOOnQ7vngbhIWJkWIcbnW/EFuLA2KY2x+H+gUkj739w/a
Zs5Pm5eBPCaA5Z6EojHWlsFr+00SFV1EaZ1h3LolOz47ShoBbhwvFq2j+Xo1pydi
cXWy6hSS4RnmqQ/P9MCLrQ==
`protect END_PROTECTED
