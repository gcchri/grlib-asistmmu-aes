`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDfafIlYxxMiutELiYOICwTtIkT2eV9VC8dvIZtfrTdNefPRjNDUNAptUivlk4ho
bjcNqdcWI0wdMnTZgpamcnuuWVtiKoYNvn44u7HfjRFUxA7r4kSd5EpklCIpjlyB
q681Ep99O69mKbqzHkc+n2865vaeckxtSlSzjf5B5Q64z8aHtZZp7HAvpV9Rom1Z
Jn1oIMkl8g3SaQpfXmEtw7lqye/FyIMRDppjWSBrYoTGx+15jx8mIfMLhM1Ebdks
rEZRXq+15fNXb9koUS09jYzuxUHuoWS3wFpMxIB0ojsNdxCi6/UpGLBvLOg9B1Aa
4kM3bev6JgpjGlIDKs0jiFxG5J/6A+TO2tSSDXHZ5Q5eksHkQRQ/rvpn5lvA0ART
znfxPdcsUZMxTZXDuvcF2Sgnge8TMnKrW7ej+3vSPhxXvDvNSNnhriBGZUhwVrq6
P8Yy2EQe04yN3zjeJZ+P2WGgeG7HlnSgk5PzgZhbY41kevcVFstShOhqpQBDG2cq
EPmrdROG/00fAczSYafNhMQOOadlXckTecTFFvn0M+xsJ6tHNdlNLp0NRCrhyV18
7esFd8uMZaGvfOFwP+LdUcTn1158ncShgVxLS+nfga00fZVhuk5FGMuFcl0dKUX6
ATRJowkT+n+7hrVoXC5EjyQ3vYimq6nKBQjfaI/0nbGCTHg7fxujhMTZ7dqUlN5X
Khl/kYYy+rq45jNgMbVKUkx5ANC7rHaMTYC6KPzqaupLlZYmyMlqn7X2vjbRGEAr
D5dtfoG4fEZqOk6iBrdJEwKmk9A809yF/6KuiD8gnywfYMTtXTTXiqC3EOgHheDI
2lDvEL+2N9hr+ymo6I2bPD2zhL0ZeQKlHuqSiCnO5gj+kcj3rE5oJMt0ef6xl+zB
XuRm1hAXi0L6xdJuGycFMGUyXG6KnwbuXwsa5cKpPyVOWDKgdEeLRB0clSIXGWdP
EoSP2PFV3iTqrfPLM5HwCbDJWkSv0DrDFnKUu/ueiteuQmPhFMNDCXmECY8NG9Fr
ZdKKAkMf5OoN2i2QrND0YFh6JkwAmd7lKziZAaHra7kaUxSD7eM8aV7Zfrk7o5FD
D29qpJJWNEOsDCfXWJ0wLBWKJz793xSoQzPIWHWKGKfLgoEx0CgLtX8Fivw2JmLJ
+XGP9Ujd7HbIRn6TOPndOfenStO5D7UCxJz/X4BPTb0dMt0C/2SSQqcjJMJPBXaB
yntoWIwOYkb22w5gEzXOwgbyXkskM7bE4keczlzk2TPCWLVRrjjzhLTs2uvGghBK
kUa6dtWQHOW6/Hks4GWjjt0I9+pMZg9LHsTGRDcbYawCEx1dd48L1dpByHIEXO92
`protect END_PROTECTED
