`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5sHITW+CzWrLTwBI5czHuw3zMsy0vqUGdnIWqksI1aarQP2a+RDT8g/mLlVYAm6C
Z3xdqRvW3JcQjfjImwffQp8aDb9bpVzBQRcM7PcDHw/azQWQGg3e0JZrL9dBnWpM
XScw21TTDMgAex42jziIJS3hDzTu6FLxu7xQnO5xQ8ZG6a2Ql8VOlz6jzGmRR09U
NF0NvNUmZjDDx3aqAUWJZsQ1dc5+8lNHGsyh3QCaIOuRG2hRYq0xInFxj1QLPSOT
Kd/qVt1mr0Ufq+7i6rp5D38wa+749jhLYWM0UehKqP/cy+jkrt0WsjoQbxjFISNm
HwidIjJHlcoWZwQ3FAA6BdJN8m/UpdIWU1VpL7sf+HcasJ6dzI3lY6txeKp94xVs
LjAtJvioxdeA6ErcWEmsr7Jf1Ln7yQUEshOXnqtXlEaqX+44/QlgajqV4jnXXi/p
BWfRq3lDfV0Hth6pZEKRsMDKIBpwcF71I46dWsKcf3VMCE0MAvxPCaz4qii7Isr3
RBn9m7j+RjwF32lm/FiK7eunSvTx2TFT7/eESiDny3Mkj/05LFRqp/6QgarZUSA6
I+BUf26q9OjJIdySAhDwIFk0XH400Qee42ghs5mGgh6b9pwBZ/K5RcK9zSXnYc/+
4UELt6SLtDAe+nc9ZYg4bacJBQNLlmIToyX9xDvBL4jE2EDljljFDwLwLTwwcCh8
Oq8kshQ270GX8XFKnLe8rmxM5iGw5e8+HHfLOg4iXg22y5AajEgLE1tq1nCc37GC
MczMxTU+PyYbKDEFyyvUfA5k+3LcDCZz3DDoN5kMNuo=
`protect END_PROTECTED
