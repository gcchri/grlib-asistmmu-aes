`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ycsq/NgQW/pA3Giz8f0VcGoYbxBysvM9Xg0T8+p6lfJIKw4+SEx7ishmtkj7gCSk
I9YfqrXsORX3c8NMjhtP0yzXFcO+qa5IGrrQcqinoUBGw8tSUhaa0xXW6Tnsnpyb
2fZ5hvWBmXaMchlVQlRIVAkBCYGVatk/j+h9UABGpWpSDxqnuTMUGrEB3QFtqKp3
oSaWsVFvLmz/gGW+OmNK4WSz+zbTTrJWUPhNuPHFJjdcjOlGEQMwaykbv4CLRBRS
jaIFD+N4CrL7IJ7z0jstX0Du4Q85lrJ7xMNNQSICAgFqgeVxdNo7ygwetwL05w9O
ybZK2cxt/Vk0LCo8hNfkluFDdcwvcEnolwJ4BHq2mfpDiMAsa53OhLggFDxC+P0b
V99GSsD6NFpLKe39sdoCGCutlCKiW57sUq+WWQYKsPjJX36ahPHg4rO2gaN6lLyF
HoY+FHImk1KOfJ2HhNPfohV978NGpK8crtP0CEl7K6M72igvFDvkt3Dt961X91Vp
BQMshHFPMF0RT+Ahx8JGLHvnCsDqZApaV+KGw5ZL4fs7XxqTCduDxlfIFYW8ydPb
xdgQ7njTQR8JhpsOPAA3PQSxVAsrUBtoZtXiCYIiJEiiwrgyyrVflktET7SXfaf9
aZsU5pzPFeFTjLbe+D5DpCSeqcwKV2nV5ilPZqtd2xiv9U/MySrZqU8+ajyQFRuh
GvjSVYKaQ1nH3cXyJA6U17tu7fsHOZF1LyGcTx3xJIfXnVC0FYD88aikSTWcibbH
0eX7mBd1LFGN58TtNKvG981VJHjuYXrdJsFAsG35v89tFDY2lAoXeRtACx5ALxhS
DFt9Y66x7JwIkL9bUJPo2zQ5sp+YC3SQ3nIvtm4QPnAr0srK3d/lAR/SU9JlJOtr
/IyIkYMHs01rL+b94lWyJlyGXM8F4YfFGozosfI2zHfebiVAlnNuO2cOM2v/rlJu
KP96jj/3vI0f0K1XX7OycG0NTrqoFPn2hdZgs7t8kXZ4NxX5lJGE0n7T7W48ywaF
ZRtzUXLX3oPYwR/uMYKRnnyOqE2KD3pkA603m8BShUzSoiPzqtAW82ivVlD+lEiP
lGwOrHH2Kw+jZn5e2SqKrJ4Sz8/Fs7Zmv31hT+7Mv8akMA692I/HqyPfIy+5s/rX
6Ja7PcCYTOW6y9Wb16jZEqyTAdfReMTjM3oSlTeFSYXawjJBgQHDCzbQtbghIg7G
DrMx0fB72ZUvctNokitfDJFcyn7xOIvQ2lSjCxl1GqwDYs4G4bxvmxUp7IUoAXzz
EqZFjEULqebqLxzdT8kXwZY/6+UlrM5KwEPAjVt4zdkLlYKIrLO8muH+2knNCZXg
tmIPqtA9EcfVZQ9+vC1OMkHc9VvgcE3ZaJdFoUZIuU/blV00DQmMHj1gLWhN9A0J
ds+2YL7QEX4s7OYcqk+LdcFHdQmYhyd1/zLHKcJU8YeTjLqZMwONTzrSjW5tHY8R
srY12MVxTyaAQGvriGX+znA//yPjlVpQql9ZEAASsHcMx8SV08yfvi7WTb64m5R5
i1N5nfiY/QZWYm+h3FZcXSSnb+xy8Mdckcn2Cm5kSRdZhcGQp0hpcZGBUjscmp9o
ep/vdlUM3So0cXYN7W++9YAjKXARp/gXE3eU5cf+gUD71oz5g25f7jxIflCJ/kg7
9I/UkCTsqwxIJ+qmTlA34fuZ6e89GVmBV8QQPnA0qD2VwYAPPawj//kI2dAkVMx7
CEzma6qeeocChmXhoumNTU7g4YNzd6Ve4ytKtebO4eJpVNk8x2pI9VoOaThUt++i
Pt7F4TLcb2mXvH2ncRSd5ATpeEkFQdtyJRfyMRzgWIB5ZmzkLrY/6GgFBoLLE6gW
fl+7MwAU7eNWFoewh2OWcJteABSR6WCVNr/Ppz+WgtHEXRCKZiAXlOgHctIlbeoj
`protect END_PROTECTED
