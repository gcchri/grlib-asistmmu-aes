`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YpQ9EW2CVVFdyO1Q6fuUVq5BJlsGPOXv++VCWmVXKFv5vgfQfbTBH3lFrSOSKG+o
Rq1ayvhrQv8+xaD413dtgg+k8BXvGg2RaUPWOgtwOwZIxAgqkm3+Stjy0q48XROl
oGojkuEiZKbdtJnVS6Wt2O7yoQw8uzbccNl7AngRkwpvgnVZOOUJHsYhYGuwoPFR
m41KIJ2GcqVw5++CQC94Cn7W9eSNdKE+ED+EgMqoENgz1kF4PD5+stuHJK55DAwe
E/p/6wgwiLslQLTy3dIJNhcNdtbEx7N/Bq8dj7AkPWvPCdF8f3OqOTs0XpDMzpyC
s+wmmv4cu05lioMY7T2z740fYkOXmP7iVdVItCdC2/L4gEUWK5Fwx8kEHPw10Fcc
89ix8Gjppr2PkxPbpAzrOwaZFpQ/J+V0kJsRQC7Zx90jtovRhEVugrabCRSLXA3Q
+W5E4oq1TQjHnJc5Mrx/tsZTQqmaJ2qxzFioD70dxi+QyXCE5E4nug292nvxNNx4
W0XbpT9qEezIOE3kQ2al8fpMbgWtztLZRsDUF/srcHBNTb2pba+pDzkJloaRegeh
YnhQF3PfNZWUAMANqwJl8UOWzb4VfhU9+d3CVMF1yJQRSO45MgmtgK2AfWKBsCoS
gn+sJDRGFaadPn+E7BE5INRNtof++sbAWw0X2UmsgmPzcr4O35HBsGbjVDvAvnOB
YDI9HMXLjhye7UI8g6YFJFa2B3BNSC6wj5nYecYoAY9rFkbDNjEdWzCwtAfxn3JM
`protect END_PROTECTED
