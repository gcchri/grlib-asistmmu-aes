`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mS/+UFL3ua021DxElib8+RmTVnRdnetUiKkFJitoBFT28ONa/4ehH6BXCu8mMySk
by4tX6EB9MNrDlX64wZxKmShtyX6MnrYk9MFRNPDRCu6Zm8/TeLIZeEnUppmV96T
zs6/LL6fHqgHBguDeEqnYSR2RerB8l8PSTdNaT2/Fw0pU7AHl6MdghzkuxcqByp6
pU3yo8oHnvidOcBVBzDpDSSdEQIj5Gw8qB7dKgDMxGZ1AZlyHdrqvjhGS2wmB4aE
AGKmi8+25MMqfdGov5hGw/PJTXV+tw6RwWIq+tRkIW5r2Bm8bvqv/RuIz7UvegW9
r9lav7e3mAzqwVYvK8X5Y4mie1TzCUw9Jxae25EXBKf+DWQxUugDQcGfqf8P/sE1
HuYz8aS3yFXMlYIGi98H5ywBFAeBB0Jd5mr8e0+bGE4=
`protect END_PROTECTED
