`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZSJz1VU1J8HdgI5R6q0taOT4yvLghvyR4DcJHH10/7cPB9Vbaj8ADgorVYzCTFu
48ktUpw5WP/ipm1PtBv4NeI9RIArLXrLRyV195Q09YS6POS+PvHz53CkWylmzuSp
iPNOVu7oIlwJJ4H9ajwDqIjJ2oHeRpInnBDf1dwt5RWla3EesogpegmBaZ7Hf+wX
MG447J9lUh/WyD2YypZoGFxbP4K1TYXEcfKFSkTxu+HVCIeKLHY9ldjZsZC1EeoV
tUON/aCQ9jGhwtI/qNbauLb5VqDFx5c2JiaOumDNsialOOUaWy2mB2ErDz/QAenV
j4dM1Va4sprcE7ZadZgIvSCUoYqb0K6NiSIp/7snHgRY3yQ9Njl77q0qb60KyUH/
fCaK+98xHca6Bx3GiRMhGm9ULl0TqW0NHNKhjuYG8CEF74svhBNZFcA6zbWy6Yv9
HCC/6tx28dGwoymfHapwKsbZV+iHQp/7IdG7tfJSCnGMEgMFOiCcjPoRdKZOglRv
kwFu7lm8CTWWRtvoIl25xrTBakHLOKuzliw+hBgMG1sR8C7GOspZMXT+zcbM9TnG
6KeT6CoLsfPkMRbQhmTvueO1QV5D5eO7QJuV3ELfR86eE5lpe7t2i1ry7Ic1ACJT
mi/ckd5MM+f9T7eWamfWFLujDjbcxmUhmBpBvRPAsJKFU+ZH0SkMpJgu9Zt7a13K
dn0JqKgOtgE42jyx+wjjxFrzjRn0RjbfV3hmOdMTAhg=
`protect END_PROTECTED
