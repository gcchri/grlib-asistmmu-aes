`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pHHAFgAN7yfo8z/H3NBbYX/+1Ei4aLOIirfiCk0nSmoO+5giGuEBTSMVa81CgBMW
p5uz5jW2XzLz/3+ieEtFC5JAG6V1Umeq/1QsRFUdbgdJJozByKBgXyGN5NFqi/P2
kCO1aQAt047LQXyiQofPcaCGtpmTLY4w1b6rZdBqkPyq/dMZYflViVFwmeHR27mW
jq3I5+mz25XvZ31Jh55xJszLZR2viT+PH5akDLjc8FCfwzZ0t2+JbtNH2yPz6mZM
vZBOf52UN3m8wVUg4wgrkplhnb0ktqNUPr6nMciMKpSul83rw7vbl8gARUUD5jhj
g2zG3V6F6tI9a4bl2SgPQTz5Fj1WTO2PNMuDcLB0OrtIpy0kWEPt9RQETmzUQM18
QxcYdpP2LfTjQYvZa78nsWhbVg0vG+haqGLls+jKGch6iA0ZDYX+GMclfFCrOosX
nnIksjOTaRYbGmXBrOUvqZ2WHJRiBQsdmGnAM17oPMPfHI8D1BWgGnD6cB822zOQ
VeSZ1Cirk113UPHGHvlypleI7D1ZGSdydmHEC2LEfTo0KLzEqHaweEk/BU3x61KY
vQ7mA6gJVr9RTLElPWn810U2XEisl5a0/H7DSC8I6zWHVl8sLSCRpcDhCT218b3H
`protect END_PROTECTED
