`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R8DHRviXXI/DEwin+LxBmnDn97u87jyzVZ0x2a+bmvwQJRXZBXcszL5HUOIgzzbg
po5Uao2b6sl9JGrW8vfS9sy7RgSwpYc9jbDPHVyhvuVfBSqkgFBeCV1AoP4GECRM
byZ0/eJw3bmpAaAV51c5a6NsVPA/PY1KVqMJwkbmYjJMYeZTgnA9gEGEQX1Kt7na
vOB9XPES0ghbrJXaTRZfVE6xWVI44g2NM+TsaV3drz+SCkNuVWC6AOSgOWN8qYPI
dagiqRpTYvNaRTYTrBG5miNL7bzObq69mc3yTdmKHZJ3h8c9W7nW2kvOfaMK5TWO
sqm9NmFgoJmRN7RyACuVrk8Mh/6beD/mZhqUjxEseVAj2n+ouhO6tAdhOGPF0vDn
xKreKaEdaRfI+Kue+AySYoMJUfWU9HNEYQIwhfbJzDiSAOAihcuVURCuN6m8n5Nk
sNipvWoxHs633lQvLAihm2EX6l/JBQe0jLYTuBCD3rtl/jlNNPS4ajDqHe/3L71j
xovgz7sHZ4/B1rFKH197JBfA/d4WgJGLP2BeHdattX85PKZTNWYzH9o2OFDw85Ds
EtiSB5zpfK+Odd6mUo6T/Tg5BG2SlHofA3EBJt1bDzd+V0/uYOdlJliJ/0fZKpgb
EKwbdZoX+VgEDOXguJf+0h8Y98yDvFMbfu6t/uYo/1kIHQgkwUNlZle8u6Q/Q6Wr
BrDUgwf70r0J5Gqn75iFG78jjIhZAkTJKSUGWUdxHbqEx5rIXh3x+MSWNYbHZebq
E/GkFSxjvLUeb0AKN5+0EnPwSYOqfnVi1t5Vivnk4qBW/71CuLNZ23MvvQRYMJbN
FfnFG5NS2PcpIbVp4trDESZSPKEO7wg5/BagJOFWQPdIiMovyeFnt4a7yM/uTgBH
557wxOPIuchip7Wo3l1IlJU1x7VAW4YbLo/yf89X1MhyidSMZM2buqc8YsCUxMc9
RerLXFScXrWRyKua9f6+wMnQ7ZKSUUPTAIrisT6SSwMogafZSEGE6y6oUgcPalN2
Wyp9rweenS8KsxY99Sy93WbYkHgv1TMQxtIF3FoPH/Usdazo0RudVE9sfGp26P6Q
m00kqJKVRoWvhFXT+XFa8vJHCnWt70Sm+qqD+agrJR939Er0HyVMLaCzuFEwGyRR
dXTgNkknkyjQk3D/eH1aZFzWOz0V4GkPK+TdlEalLoQ/1JVeujI5G9K7ekFNZ9Ak
EP5RvRfOCzKaheOx6b9CRWUlCGQZx7GTYJ8UyFSO/kpn0YA+Uzd9+YvOmCAXiFIV
48YjUuDZdz1l3zl7l4pVnbHEZoMOZeGh+ml1fCb0n0G8p1AsH0OMKTiqNZoeGFzL
GZbs1zlx1tpS/Ar/YDwvrcO46X6rJG6zHWEMVDqRGSZ/1wYm4MX163ea+5/vkx8x
Vk19jp3UB2klOAgIMIDM53nQuyOeMI8q3Xi6qpo4kaI576C1Vcnku5RmyENVT8m2
YIBzmODn3jF0RHBYTxNBca41UOP06WbpCzcs3vPCPmn8bbjdcHcf787b+i/gcscw
dUD/laqwRgqZzeqFoHdIdbnp/yhUCxyUkiGNkDMYumQ=
`protect END_PROTECTED
