`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kYdZB6TBDEt43SRwTVfTmJaFRT+4G76lGkf93t+8z0xz2UQP7LIgJrgsn45oGFdV
Sf6CFXkfC6uoXegBMuNk2Kdeb8JnswLpJeoGcL/ZGjIREeqT9N/ImJdx15anve3x
DHA2Rc+uDifJNeq1RDzB1tGxdfKi766m19VXVVrKgCKNPW7BHanY7tyM5yQqg2jK
/6mzojqNH3jRTmyaW8g7OGq/YNKm1VP9H6ygNYRz9G/5vEwpkNWcridL7ed3ivgp
zBseCsK16tK0ubzBuvXlpH6ni1+ZP7rGgGbJQ2qzpuJLDfBUU1NIXDK1D5aiFGv+
5JL7vr4k2UQQVbZCh0ZwMA1PfhasglCtKg7FW3MwoNjHisoz2mw1ajOcWg4UMi4O
eSAkX+C1/5WSn7Oee+KM/jUpVNiWxkv9eDo7WowK/91BQfYY6mg11y4W7F/daKPz
`protect END_PROTECTED
