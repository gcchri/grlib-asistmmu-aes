`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLrlM6DpFuL969+5+kx76rZ/KndBOTEis1RSIRXYM9330ZFkZNpKj1pQ4OZfn5XM
FcFFcyDCfGGfTDFpGc/LAkVCs2vOybuAwkaXTGYRMKPyYbJ5Q9pBUEZZec2tmR/q
LOmu2lE00I1miUjoXmWd0bd5vFICFXPflWe8ZbmQfXNgNbjr+ToVRZAHrbTctBEl
VDyuJhegCgXEQrD2liCPmlsC0sBLX+0IM5FpXn3S9xWS/+2IrOFPJ4KfSJRiqIRy
72lFt/GQ/Hpi7PyzF2hQlIxLjxv7q8bj79gMbtUbnk6kl6TXT0BpPsyiypYwv1GN
SCRCIlTNadqe38iqqqXl9rDFga0L3aboDLUAc5Bo3sVOu6Nr2EvOHwTypH9OG9A1
3mszfJVk3FNCSQ8Nv5sIQaGRkGtoLyQGFbXx5Zcu+x4kvQAuormMipOw+ZpVN77h
zo48JKO+lLvwX1mNpH6qHu5eXHPnxFMAARq6CS1Z4Jc=
`protect END_PROTECTED
