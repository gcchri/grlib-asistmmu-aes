`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
enOb6ypPjj/G1+KMRf8cxLF7ZrsSNWYFe+b3aKs5yyB6YyK47I1S+y6I4aSm+bWx
qpnuojPl4gzJmkE/cyBRVap3xyVvS4KzjI38/B7vsVKEQKqSaTHSbYjMV1cM6mFN
Ycnx61HVEJV04faEwKl62+tDRIAaQh0ygk4yt/rXfUC5uOyZMbBx233s1vLrYHhL
7I/Fnq3QswmXKe6D0mAcFVxI7tIWMNhJHix7Mf9Gn60JwPKhdeB501h6/C3vfch7
aEzPNg3dEby27JBLOkqXDLIMPdVj2w+uppaZfndIgCZ2P+/njT/2abcXZkUYTIFO
t64yHVq+OIzYhvJMARnW77tXcPBntRMgE7A0B4HpMyMep23FP5v4hzrQKublVGW8
xGIuJ4M/Tq99JAcmqlPA2eyQWzBLmpUpChzMqf6RSGtVlGlHoXUSnXftvZq/j/g2
Jl185Zs7LtbH0Cx0boLAbbyJeMkATW5SYKsrh1e0KyI=
`protect END_PROTECTED
