`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hMg7Lcw2pXVGguqQJTfjL2gbeEjZEaVpGdCVmEY4UuXzDoppt6zCwk75k23VTj5M
b+gUhYHuPbwKW1oWQEl95nq5pi1ed3LCSWCjyJ896zwjt2MQTwK+myY+CDBliW5r
rOiqKmOWbVOXOQP0F0ST7Z/4z4BVFHQfWAIAp8JHNhTp3+5J0niHXSNZbQb2bG3N
EEzrIHqD50ZEITD6stKWEy2c1+8EsW6gFBes24A/qYsNKaFbyVk3aGlIGT5Zr7yB
Y/AkWTarHPvSalydA6omXN6a3NbyTKjwP7wpylbXhiR4YUIItsbQKBxc7HmXMrxc
EsUCRjpS/iomFQCp1/+hj3lFz6x3x5ncdEJ80DVyupHTENKuRmoQW7zSjymTfe0t
CeY7mQJ3SKGqnmKaIxwGnwvp3A0c877Bd/CUilVwbX4wWbJranBhdSeqc6JBY8PK
PaBqwQ6IGPiFuV0UNPS0v0LOVecbs39iT0npISJJ+ltBRqjlv1R5Bb8cWSVDFMQt
wvBFbiUXF4wj33s2Op1ayXHW53zdZqDC7s8Is29qPUOqVSKTJwUoWoJvX5Lel+oC
kUnQ2qBAQ6QFrTl3vuUY6Is93HdNOcYBPj4yWYzVO2gqojCBf9UWDThxQVxAr3xx
dX4Ihb3CtprOjTKFozo/zE2D0orF+sTQUlLRRSYPsdyEZXeVWUkzjia58cMuMQ21
vJSX/bTLx/x9QPEGvCsssqJHkjEYM9t8gUw8WW5UyB+mq+B06+hstghw1F268+8I
HJ2c4m33yXD9ss6bcIh1zA==
`protect END_PROTECTED
