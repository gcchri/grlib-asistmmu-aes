`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CymW3b3eIX1Q7aeO3EYCPYYAW50TLc7HFZMvgBEEsK3NN4JwPXpagkQ90+Gkc9rw
4zDjqtOM6THkMVRC7b31XWTYttFHOkuZWVaTBGhsEkN86b5vWaxiEfHxwQFpD2E0
tVn2bRS0TSXcX+zn0OmGVSDcyQe+IFc40NEeykhy0fxF23K/x65ofBCAci3/0DQe
pXM22Hzi3zPZ3bh0htaZsz0D/STFQi3TW+rqD57KimovzmtQwgkEKlV59zLA6F1M
Qk4nB9RSbJZnmP5ZpjzLOWQ7bKozzDiMXOexB9penOIFGpI9sToDdQD77W49824W
gW6Y+5YGMLFt06QwX1ZxJV0J1sK4nzmwzl4R8ho3agPZD8JgJ4ljoC/uIdcwjhIf
ngWxobSUc3MdnbRWqq7XY24bMJa5tiM0v+Zsc/N8bEn5dvPr8GeUU2ge+nL70jnZ
GnOoSYIAh4lhiy3vxTkC6wuI1XtT5idD1nW833JEVlveeW+bs0sitXJMa1o17Kr7
nlxCIXJaMM4mbIO5U7jFzo4zkmlBfDjcQZaVchCcUX61eND8VK+OkNhw6+CCCyNK
CQ5alEx6Q4UvV34gIVDvk6rsZKBlhVeEFzuAYuYBeVU92cDbx2mI6vUBREC6XEVM
+qVeMeNe0FJSiJOa9a/8KbQsVztqYIHj4xsakojd2fDKaU3FXloQw29NWjqy4O3s
D5MaEROzwKmBPNSVYhIouomL2biKyMRgcQi/A+0MNdLq+1dhMVP7G/pBtisqKsNh
Qf1GEUKRIta+/i8E4oR4Cwb0wF7hKuZcuzQ+CTwgOWVVDL76TRUBDXFnfczok/4M
Hr/ClCocS0s+9sfRQn0SrTrg1DNGwLk67dquJZW+HzdBAuJ9Iu2jBZRLTQxhFJzb
2/D7g/K+nE0rRkTfSYgljqnXTglxu64yNWVsMHDnMIc+7WUL9eYDIxd3cXVLOxvO
+gpt80VBxmNJnraSERH/hSAtkpMGFZ4/oYzsehEQ6BNXoXUeAuOcTqCJ2WGfAfuD
0l8AU8CKRndoU9ODUbdsAMllFxY0WL/n2H9/KbM41dHlyntm2hubcalREnO6Vilp
LwkNrxYmLA6GHPkcmFLJB6kf5vP7b8mokVuaKQqFOJwdLizYe+4tl4ZDZOwkQrpQ
7gVecB0vEekd6ouAdRqPaqiyB1+zJrS/ugkGW19yMXTh3sbHrQwwJNbBn0e9FFTG
`protect END_PROTECTED
