`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tF6uUfx8mq7KIq0ueHL45mEuEbPuknPYeTZqqnMTBD0m+oIzRNAMSIGVtGL1+Uku
mhNvrkMS4UDB4D3CeEN+t517d1SvxtQIpgwK0u8NUvkFXLRcqE6A2fwFMjy8WyJG
SakMnOm9D3jWSfsPAEGtR2BBWJEb+keQ+rSpK/7dHs0mLBYUXkoP/qfcZrPJG6TT
hiDXi6fRCuPGaLwUcm97SVafJJzA3QcJrlPCpXMDLEEPIZO3d/XC+U3aPz30ox1h
2cjATY50IJQ6S74Fw0dS9yhDitlJ3rR3jZsUtpIfhNa1tuOJH87g9Rkdo908q0Qg
CiudASxbyvj4XKb5hWxe+z0RE0pD+t4OkyxCe3HnibcHZCznwtH7PTqtkMGH1tsi
P01qxta0oa4apiIcwl6OPK2RQmsu4Qw/PY3KD/M9emgssXS/AjLCJXyzGlyCK9W+
EwJFYqyQ6VClBObTPH6+WJFcXAxec+kUDWYd2i/rjV0sT0pIewOaxiGe01P5xaPg
pRHNJvkb+5e3w9oP5K+sJ+LwU6R4tSgrz7EJvLUKiueu+nJO8mNQtCmDPwAbpX8d
g3k4RNY7ZGiOXs4Mkj0GUtmARq68JoE/UJg2qazH5DFzHfsGdGvnzkyw540vz55R
JNPD18+PQZ/0wIsBWYmyJehND/jCorebRNIBrH7I/cyiWVxBURGiCNdRnC8c6IU0
nb8MgYDZkljNU3YSi4VYP6J+U09kBHAhWE/Uupd8ZorYrEyDSx5Zw1zptBDwh6u4
kQTHWtK4zUH6Bl+GCfcQqZa71eG+fKABpo+9Ghuzk3XJIS9b9UrNZ5oKIdmxlnDH
o0e4PK7axScHAjQzzcOVwue3j7oZabELxj+CsqrwRtCECb9OV6l+q4y2k8m8YkZp
K8PKvRGwJob2wveoxUN34R6NmQ+WwfIGmd14kZ8IXH0t3o38uM7efoCU+ZDJ1Fhg
MjnSI/0muFTMR2/2hnVbykIcfZu4R2nrwLw4mg/iUYr/1BAyq35zIET49m7BON5f
zcz24qYJL8Io8ITtCb9Vl4fVpwWj+Y0mhbqMXy/30T0E1yzmlQ1K5Yzm0i+AiiuU
DfMEAg9jqKO1TvgkEue2TmE/NqqNMLZvlr7Yxzvdo+5Y1l41jfYiA0+Nj5O0w8Gn
KIiab4AUIGJbx1OrpBJHQ5MF4xF/h/keJhoo+2X5Iq1ZVwJjBrUpoFqjGUK1q2Ey
PmK0qpIJWF5avpm28dbcFbUbgmr5rjc6RgOMRAsBonL89NeVC4a698YR6mzOvVZ1
/+GtnauBUnmnGLq9NpSNMmYkTIcJA3ngDhvMeJqAHIOkE2vftG5iVlmY8+pc2b99
VkfgZxicU25bGfs8ltrx60llzEDb6pxM/NCzYyDwsr7hXt9MVcKBfVBk39bHeT88
vaETJ/FDVz3H5Pu+Spofky4OZZh8iprPojsQi3FMvuwjd8x+OfxeGXA3DzyRyYCS
6vwsnVwgTlaYc9BwWp361oL5Nz89IgKMNUYrTK/hVoyaDurvbM0eT3sm2yaGYz27
3ko77ioY5jk57+6mv25NmUDsRVHkahyeX12OcK7uADIUDETDX8l5bpzz6+PHt2vM
dtaJeTqOA2j+qoE0+DgP5DCfirnos8m7IPbosI9dkMwe72D6RV28p/vKOe/UUsWK
BjvVEIv5rgSjYima+5EpqVaZeqXXLqXHYLM8EBnRJ+vGAogfmM3qIHqYDQh4/b5F
2LivctFGVpn1hQ/4+e77MQSnquCJmer2zcpbngYbAykRHgHJu+P2x4M55gG0tMd6
fWO36R1ROsMyuP9zieWk9fYSRpHvMmmR7K5jfbz9X3ijUOoPYI2o6c7KKS3YEsW/
22w0L9oBGtfhWhWFQ6UtkXFIk3F3FKSOrdweJZ9JAcon0KzCGUPqkA7k3p9E+Mpn
O2iKfrFW9TixSo6wWc61BSUicB7785oTyu4c7ay7F1okrnwh5blz2ahHMbNLV4jS
VFLwikOVErIVo0rUGEMEVgxTRuKcF/BoaMJLotoq68FZPS1l6+lHzNgKZvMSZjgD
LuruDyTqJUxr0qBdXI306g2N6gjx6Ux++rgzKv5hAXeRhB/fn91SmZyUVLcvY0oP
XWtrkvSp2qixgBRPGHUuV+l7DE1shHOEb+uGmjhoKBRVgMS61Cf1AZ5ZOzkrvx1S
LW7Datq3JT0jgozQ+EeCJR4NcouOHf5/Nsbq1msI5/ahqx1Y/ir1yYgNDAtlhnDu
f3oTwfllFpYHnapETgKNWXP5jYwm43XIhVxAgR4Vl2LWfkpgudtiVjcLy0Ov/DEk
c47RO6Vt8LJAWgATkdZFDp6dsTsclSv6gvZe+iQcCrty7JUNkjxz0V8xNhvDRS6N
T40n0cM//IoM1dw7NjDeMMDSoAVeb7sFXR2ML1NC4pIvPCvkJEBLyhpZciS+CQEV
2kqUXe65p0G3Zn2wILm4Oqf6dIPwrsQiQQrjy1QGG1wPGbG7Yhg5a2F7MuZZEvU2
M/dxVxiSZQP1EClssV+il1a/Vu3/TlvfOHtpos2nKedk7nTam+6GmdnKunp+EZOP
CR4LQndVa6TAdb0oUyKn1XquVwgvqqJPAFODlmZ/AmLytQ1DTbE0yivUJVcUNFXz
3UodFMLmizfzm6mvDM3EPYhWegKlf6ZM2PJTC3bAxnMdtxJnHdW4DbvMpUvhwumn
g+Sm+A7JpdW7EF0P9urOCaQisQfJJPByA2GPQLCYBt6vrE1wNYBFI2f75tF2BXc6
r399lMdfx5LgDP0W7qxZUFqudXcFrInTpbE8S84iTpck2bSUxTybU8noVZ6c8dbv
0aIMdDsJ8xsVCoVZxj/aH7lZFn8uarp8odVaXCFXwi+V/7F70xJnfJ/MQpH31Xhc
FNBu65KNl3O1wjU7596x9efN1I5QhVnp5MXqS1UXx7MbkRmlxE6KnPriZjfmZSgc
V/lXIv5C+Iq6J0mBvoVg7dEuBRpqbReuhFekhS6SE8dkQMIutjd9PGk5TC2jvcca
s9qIoOGvew7vyn+5ZWzLcrlqjVPmYJQt5VA9ZqhC4mBMNIVRc9+I69LzJFIyDZl+
TuZ6hdZwJhmDk/vj6zaswH2WFj7FyjydDxr6QoNw5a8Ere3uvelS4Zc6wdYG0yI1
QqrpP9NWNEnyG0N9Z8POwapxNN1x4IIg2yo8RpWqd4+zwruUKO1d7NrBDPPKhrju
wJZkEF214LfMEsO9pt2rHKzYH27xrr4DnR6sHf8vYxvgroi+2oWc6RKdWf/5Xofp
t+rvEgUXonuGZXoUqD8rOon6SWMAcHjnvjx2oxcgn2FQLVOD9TqGLD1pMV0WPWwG
PjS5mwN6+bwMVsQPj18A7NpvtXWz3tlokd1okcxGeO9ffx/cl9pDIhE+zeioBKe+
SjWPjKiOw6TSJjF0V9P3fgKiPSDNVQDoaUn6fBXipLlLN9YOPwA93YmAbo/g6/N7
qr1OH6vRheqEkeaGJBL8Kye89XV850GuwjpS/7B+DoPH88/JB/19WZKiS3LZM/Gz
vhoVEazwYpJ+vPoyXv1GLqt3HP5xEtMUPCgHRo3F5VM95vyLR4lL4H/FpAddqw2x
S4pOf9GRKrWzWv0Xsr0hsiNhuucUALIScAvJ9/Ibv5CEJcghZAuaK8FdlTcdLexo
xxA7UPTkDGr+WUGXJGnHU3CuphbRbm7/yQNofBAdh1RjuEDCArzxTcPpgRj3QiD+
IeHhrNHorE6im3nMO4Vd+lnQOvQpUrwHODYfgLpunS4YDQfN8oJvShelk9Q2Vmag
8p46qZu5jkbMoMFES1tZP+39uv0j0apuLGe2vD2n5hfNqju4Cl2F/9BkbJ77Y9Z5
7U8a4E6ffWVt9SpGWtafU4KVSF69bLQIpHtGuvwiVeJwtYmvjKSV3fMHfEWOrD1n
WR8Tn4YQawS7zNZat3dtethtcoS+BkRJZzBPt2YjcjVzwT6E46AbaS+rceKjK2lm
`protect END_PROTECTED
