`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+E7GjuCVfAWiFGUjn2v7pfGDDlP3FsjNQ5FqNYdQAnoEkfTyii0u1ZD8dEgTGPy
7p11gXl3OprZ/6xtG/dkMSPIIEhqv0av6u4iY8gWi9NC5W80WRoYfB84gsmQP1nx
jKLIvu32GqcGvGVeJCiAjZGmXW1VvkHEVbjVGHBgdAYgPPETUAYX6qYSYmCRE8Jb
mLzE17GNWhI6d2FsjWybEFQHJoYE2nIET8W0CAesZHQsXVgv/hpPTXXeO+42y6M3
mJpSJPmDJmCncWfJ7IlP9juQSynqvVzTaUTelU87ek9XSt4VOsKmIT+L97/cI6MC
WZ1+IHGVEG+PQBCP4g2J3g60JOQ2BxU6z5AJv9LrusvrrNLSbNl/zDptn6JShbdV
pfY/9+/UpdZRBVJmDvEQtg==
`protect END_PROTECTED
