`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1UDSRr1dw/3hhAeeU7ZxfDcDBndUUmhTiqYMJbhfdIez/gt9CM6IhbDT9gUHGB+e
PrjizVuFNyhENsA0mFJpH7CgHbep/kpw3bEk4MIbA6oJFTjuix0kTuWn94H7GPqu
XiEPpRzr/A3xv24LhbjFnG1raLd8nVs7/F7MulmvfaGSbf/5sTowI2w8I2sMy+gB
/NEQA8wgMZX/bI5m/xdhpNp3brXSTXqFaLoO8speb8nVbBv/rYMGfIysKJfGF/3S
UhCfAC6VXt6i+CD10cJAbvNgTNwQ/w4ZmcTy44js6ulTl9X+rx8faMcNgcUmGQWJ
C0pWedbD5//tx7jzZTk8AVkZeeerYwtSIdhnY2i4oN1xTLhxexRHJi2Wx2fvkasX
LnsZosDLrPoKZaP8VhZ3R7UEOO1YJWN9w+trVSsj3GoUwLspAkNgUeeZRsGF/j58
DEhHnty0DzX2CS0Qa66/o3qnGV07yDEuQ4cl9/Ss8T4zAejCmByhBwrpmoxSfgZn
q1zT24FtxyUdYJM+CEeQr/kPWjpqCEbDAUX/46694Xn1/2uelSioL/ud61Q0FmbX
0cXej5Okv8e68g0u5/Gk+aojOiptyDDnyZpVD7fJ0N1BDiVn1OrxgHKGCM88Exy3
TmgxwUqO/R9Ed3wZw3eN63eBkOsNWzroPAm3EAXlgvoDqzjcExujKGDtlEav6hh9
/Yx8zet8/SRRpAG/boD9vJE47V/KjhG3LmcVQIEoD1gQHZt1UAEGYZArkqO59s1Q
d6d1p+tNBeaWXPx/+4ptn6MEsx4AW+FSgQpT26I41g61HW3te9A3XwnXFAlBXfH4
Wj/aucV+d4rs0dSd50CxBlQPA7j4m36Tub5+Ldzq+FcOuw6exa403kpee9orIC3t
a5GXIKata/XY/bgHWpzUVxQKNN3spjC5keCq8Ls7bIyRz8f0jXSkCu+87QrJiXDY
w0EgxOnE8qT9Fe66jSWG2qnkSAPzkmIb9fyp3vzPo9//0I9Qy7qBFdFSo5cG0yls
`protect END_PROTECTED
