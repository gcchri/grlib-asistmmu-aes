`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sccQPolC9EJei9Z/RMWSLPpWO4ONIH0qALaocsgSYgaLrAH3HxKhcYjz7BP2gglV
bJTYP9NbALmHe+KgWFT+EHA1kZK/WLeRWgEgEcTr9b+zmEAZtvbW2LZ0nU+3JT+j
PstJFb0Jqq0sqzSgPS3+BI6BJbkDaaQkq3Gg9H5CXDPsSTnAtcovlLXdsBmWtwa8
rwadSwYctl1kvDwiN0oN3c6/8vf9YOSu0dhsE0GpYbrMcC4S4qZbst7RJrcUZGE+
RAaYE2s2gkXSUDe63Xbd1lkHBY5GT+88lB1pa4U5p3RLZ9Ay9VQnOdtNbALr45MH
k5fAPnDQnTDzh6JPvgf6vUbiA/hy0MxpCNVX44tqUM/g83uAhcow8MkCobQI/wWI
a2MQs786OfEzfOt9ffR1se6vfCjynfEwkhMeT7VqgfUZaxVHQv27O8Psy0lk4AEN
iS0miMn5e+gg8mTgslGDkwxBzYYg93fWjHqlV41gEm0iV5/+Z9CmPUejHOoM5zW1
O3qqYL2Yr1DqWTMM7VHayB1WTBp1MXrsiCDMEDfl5zKsE+fkCA4frPpqF8s5N/u3
UPDVeveUA3qJObDSh+oGh/kUGBeix5hUcrmCA6pVaOElbWp9xUxLRhzJ7LUiPoSO
SbVRqiEBohn3Bw4esx/aV2dNOH3ARXcBXQEqxV/PkhioB7G7TM6QN4o2iwpeEe4H
SMsSZkvouY+4Z9O+qZlsDzcdlpPwmn+wQ07TfhWk9Tk=
`protect END_PROTECTED
