`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eu+D3oF1kS/Czx7ZOJ4Gaer//OxBCi7kI1l4ORI68jfxMLiQUjUGxZoHn5sSB9kD
OjbIAMNDGKXyqvk2ftec3uUI3Ojq6nppzKAOe57agETTAaGwf3EKg/xaBAw84aIl
/FICvuiviXyWtRv287rvivwb7gTPXqU4A6Aw3531M3pFV8ACmnkwOR0Px3dRPEao
g/RihixRy0VzmZJIuPJz9q3sc5UQd5kQV3eGJVcexquT/DrHexpH8i79OCHomZFf
qfzsHJpn3/vDMAVwSte/NAuJ7tEj9YEeV5LodhtuV+I6dtSeWLe2GyT3t3AvNoPF
82fGPCxDDe9EiskNUmJJGLFHMlvsLkeOUMfLFQXnXB8zQ6s7Jb1SpOP+uwg5H2G4
jtRV2cRJXwlS160hY+6Af2R2IK2MT18MmdiQW6zwMbe31V7y0boqKnQkqb2HQShE
ROgepas4HJsundwhUUOLT0IeUbtcrmSlrW05AD1CjpAFKaH8sHDiA0ybssSSkRzm
QDpJ59QlThcvReKfjYQwGydVOGbKUqYMKu83CyoE0r74dtRvgcNCOGqzohOd96bB
cjpaRZeNOtBBZNtF62gzftN5Hvb5bFTazqL/F2yRoenQN3rknoJRf53/hseGXIq7
uH/2fzAjirqOKjT0nih2AxA4XVoGV5X9a61+ZHBwWoEoQ9LlseKZprtnsWfsa0tB
JUpq5iJQywW63RbP+j9AQVFNPyuM1E0w6ez5TJq/SnWjWtXo4pUUP+ynUpH8JLfd
UAemGx7og++akvW3WLgUmoSY1AX7buAJ7VM4XIfBEgdnRnHx300e4ARrXKUS6o+h
xUKYM/niP5nhxGIBbMIWOs5nG4FhFRYbVfUouODOnZohZGodCteQDnAsJGEnilnn
m3RNT9v00lwhUlHLJsqSnloFfi+DrNM0fs7P1Ef/0LJD6YStftz2HkGimZJrADQu
1mbBwGe3ywXTmxBq80CStc5k0rAEEyLIUrVQQ7F39JvCqVzRKniM6IBQgqYE43Xz
57hNBLvrn51xp0Z5lhwl09hWsvU3Ingesf5jEPIfMaZqdPbDbiInrFGbwJq6AwlD
oLcR4ByuwA3idXkYIU3deaE0ty33ogtaM8qn6A2Xx7iIQ+6lR6W1u7efpM2TlC9M
+QLJECSO3I9bpRBs88EW8U+yefNi2PpK+qkMiFtHl3k7pR9otdzB6i9+d4uziiaL
i1RmV+UYpl/tc9Ct37oxhHuZct4MNn51Seu30i6wFyChb44ddUzWHsHPDOMCfyuD
9d+oPXz0oFznAJSVWltlt8DSLHb0fSAXXCyTbgRkGhPDHu/4LTqBGro9J4MUMqbv
TjA7l+TGfu4DMdw4VUf5o5rBpTiBVkH3J6cmM7f7y64Hjd0Hg/7Frk2gtXecN7pB
UHqj1KBqr/l9zb8A9aoIXcHfPqRwXjb0ZmqQ2fJId3BPhP2O6uBFMUIhm9dwkckd
0ublrTCJroV/t9qQrv2zpaYyznXqETXbd9MCdHS6hnslBD2u1qd1VrBXDNkUO6g6
nhLH7JqTo/OtDbhjYGNuUk0BvVJtACbMsLvHlimnRZWZGRUCCwmSXiSZi7z/0E+Z
jo1tjpiAbW+5UNcKRa18NHVxnBbxLolui9bSgmyc3pWYNBks96gDRfIBirpoaqSA
zRJo7QL4TCJCmsSIzSEZtyFMovHvLPqQtmanENmMRipcGK77G5yrOGqDU09xIvCb
a2eIOKY/8sWClRjhbj4eBigx3uHjLKnxr9uYRJGqlk2Wh35Gg3jKSILvjyy+UVJR
ijPXpRAXTKsjkDna2v59jvnBwykefYPdtrjDBMqw8GtDYtV1cdrhtIbU+jIrPNaD
mp+uq5TGNeT9sn1ZVTHbH/NzwFrVWrqkvXMhJyqIrKeZIfEN9xXBZ532ExDb0GyF
dBioG7WSp46o0tnZzH6AN3lroKtHjOqQYXehiF5JkgzsBmjRYqUlXqiOfvK0yP/l
fPNS1r6lIYqy9iAB+gBIvbrBK1QTPv5HOQdgXsWobAQgROUxM0GIHFRkhfeZ/NNa
1Jm4jMXsrbA5sbCwfs5hT8LiVqpMXeD1XjrCxcBn3cU7g+M7601WsRWCqLdeKTBC
GzEDFVw5++tSmQy8cFq5ybZ8pN9mIrcKYH8m8G82X2pjYDmw2HhE0dDX/gdsc8XL
uF8pKI3koip9+932dvVuzCnizufeoA4G3Va2m3984bAMbbrgnMO3OCEesJ1BKYq9
rdiEj0GFoa4TR9cWuXKflnFMjq99GjWXXnHuJfaeurQawo6KmmIu+ilQ+wZ/RrMA
/c6H47ygrhSnmdP61iVwdC9AskEZcpDr+Ifzf/7QodJDEBr5PtfqOzSfvk59tLAU
58ysH5srg00NXPjxT56DaPJM6O788SxzwS/Lqo6jf1ZT0veT6TgkJAjDVv5LEs1I
pCfnqIeWaXnvPTWaKoGb7s4SXczdGGc0ztgPDN6X3YDFdcOtngifxhSmP4s+YxNu
tJJyFG/tAbU8xflp5F0BR2jKEEvMddyuktlkXOAR87GbqDxNuHbr4TgyMr3+0irk
RJ1qJDjcfb1qSi4OFr0eYtN4+BJ2t3v+qkJWSWxblekbkoZ3nbPN3k40JISkMQKK
BXNxmGPCQjXx/R/5sqM+yQl00h2AmHjBUXFWAk1/+H7OABqh8GhReLbdPREYPZMP
qrsiFPdUt02rI+S0TV3mN3VV8THgotAlrNLD90TZScOR1j4LaS8P64wtDz6XiTOc
WuMfLTLAOO8d0I7KhIBqLQyZO5KGKek1LWFgead5FyCkFz5rLlDcTKdJYdbtUXxJ
FTX+Je37yTEnwuVs1IPvSpQzmzGYft7rUqbRG9WEpI6tr7jLIQlQF7JvrZc3q749
qFZy6zt/hgLozQH3JelGZrIsYNUvqmAJMLq35OyY5nnAozC/Ev3rOaY1cdNPTuvL
pyoicaLgouV8QE8F4ugJxIYMfL2mit/Tf9BSDdTgybJUlPTJyCjm+bJ7+L0zLs8m
SXTQ+jXjscSg+R++70iOHRfvQg+vl6UydUbxTTyqEYvOVrPWZOvzte14bud+q4f/
ctir2700Zota0oeiaobJGjy3f3W8RFCZeQNpuf2XzM+G79I86tnVumPt196Jy+fK
rapgXkRr0WjAU00YMlYS5RMl/LDoLbuheagOmClt6S/iWhXJA4n2DQLo7rVHB1BJ
ZkDqB3ZOqFvfjeMm1DdYsTq3P8lgx/uiRfpTtsFCiIV2OmC2RnYjiqrIjfFONW0h
Qr87xrTiuNm8U8tlaPOVW2aLD8yQjLAgRIku0HkwalAMb0i3HR+Iq3zXm6mXoq7j
ZMsAw3RFDfL/meYcsZvvWzSBVYupXHkv/53ytCBbOf6ZB4vmx353+6wERTFKhUyt
p9aAwlnd+on7tt3UNFNbuYy2+gnKtcdOycmfq0jC2fPJazeGscpkuKo2798q8pqp
B//IpLclcaYHGko6myD9RXDLh+k3usrQsucxwQRqwRYmB6/paekKmmmMPQ6evR7d
C12QK7103gXM9Wla5g679Q5dEn4woXzgUlohLTYPiVA50i+rvzMw4h7Do3L4UlMx
D7b9FAz5B6Dx07de9ADdGGvIG8U5wxyjhvolCgvXfhcTLQjiEPSYEOVNmKFAKA47
mlHnCtantSKGyd4BtHJyRdnUwyanlNmMM87KbuMgggQL0Xwc0RrtCTyZohRAWQSq
bcVIuP4Z3cZ/sZX0bp0QHgVNqWxGU2B99b/CUfHI7+tNTawLUzzRJItYi/X7cF5d
dzFVSdv/pDr3J1EP9jd7hw7tkifOG63wZJ5CW+KVNY9lk6Oc08s+OLUmVINQt4tR
JI29v41zBpNLwA90+3tq68QmgVBJP70PbLmffsh4MB6sJu6q1tCyaGD3UxOe7K8y
ui4KOgxW6uZrkqKNE15Dx5bT7HtpZywq7UgSgLsNXX8cSXTeyYptzsS/wau//Yf3
ESJZ24VNlGEpSu3U645lpoNPz6zR1/Yiy7AsENKhhSKVCKqDmgS2AVJG3SnypO3R
7mU0EIDy293bbnFnUrhsEsBwis/DpeEP4QAxQrlDje+03MY/iP6qIK8YtLOCiQFZ
Dt8k5Krd4XI0753bT7de1D6ab5Abe81KHRt1d456wIhFnXvKFMp6yvy+QWJZIdum
TG4SIR4mgKiP2w6qMGJ0YmiJ0XYTvi3jnRzXs4oEG8j3zSIXcYAALhjM3ialZiKk
LDP3QWbqGY4IkFxi4L2nFNwmeA8Q2IQ9z7Gp1M4/wDue9oaeslyktqcSEsvhA4sN
Kf5ZEOHikaiQQrextRitzMygeCPRxOgP6NBAH2HUd2ajcGXTUJEzk+AcWZkCIuXr
63AYV75Be8mUzaY52bw8AImbwAH+/yMrFvVSzXnmRPjeTORBleEK/0oiGYvqZ8KD
7uYHej18ZSyUsB7zE0vXl2kt2soOo8qIsfVjSI6BHG3BwKNNK1afwf766w6KZ9LU
Bq05mgA+1y+viSAXOK8dbMdXCWnzwTTj69x54Ch9cFfFZV3OXYfVNECY/XqwlfiN
eEfeNMpTsEhcQTkTeymTKgC7x8II8Q7ECImQWAu/JWR0lqYmQP5DGIt0vRBaaeZy
o8MHT7npjA3Yv4vCYQPpW5DTGoe/9ztWYVRUTKBGk5YpBty4ybfHINox89n0D1nr
QYKb2JxmSBhuFP+FSTk9b/mdiYPixB6RVJY640XrHpOTmnm95aZ0qWK6wyLZ5gf5
Q7X0sMbXCt6ajg+dCgXztjifScJ9cUvlXzIOjLD4SzJULRClqZp590EX3YgVM7E8
o1Npy3GekUW/SlTw2U8xurUWKYAm1il/EuabOHAVgywRtEUgmfxU2vKU/oompqrO
YSP0JmNbn082vnQKRZ+St0v7spKmWgyqLgI/32DdOF7XnvmqWQFvV0sWWFuZx0iN
sxaPtjoqodsm577hcvjRI0Djao8G48rf+7Y7Drp4k50PiJzLICcM32VUek1QWE9T
4u+deXp2Tvs4Js48z0UATK42/O//RSgN3Iss/Je1B8586Iybtsuly2u5LNT1XCHZ
a3TuctjceM5Hzz7IaUexjzYLBc6+4qmEufqgLc1RQVIuWLpxOhuXKVsXa+KU7Pr2
TMjERH4XqadwI/ebB71krKkWpIN4ETMlGBGdeU82ffidpmOY06yNJNinE/5BtPPx
457timYUnn9PTaV75OTEwdarvZh1L8o9IHyRYJZkT9SvVJ79ZtjVCc357vDSNmM4
GkFZV3Z2kjHyb6DUsPIH7ZwN9j96Bseg/+8LJP4tgIzhF4x2QXwOWxgJLRbl/sas
NIPjrL4WdcmV2SkU4ufKrPz4xC3XW/QtK8ld0zgtWG+Chqb9EOEucEb4swyLNU/u
paOi8PFdg29Ooi1ExCrpFXgBjoiIzJmYQyl3Tt3pqR1O7Z+LMsz5F7/sZG5eU7bD
zGiycfrg4H8hMrtp5dMqem7NXtq1DDQ49x/xMotJSX7C+OIyMmnSsEPnCLE0Qapr
jvfqkNFdKPuszmByd0xFBaLN38WHAXTAUI0UszqbTsCptxXtBufqwB9ktHjP5sSO
AzrdoVs8J/HuACjJomuCuFrMPqQ3pFBPUo4nvNTDjpaLpXKMnvgL4y5LYAaTeMaz
/hc1wJJQDAXOKviXT8XQFNAhRa/NGfmdGtP0ayRIhUdOZ4SeAbTGFiNiAcPBV27o
DLhJE5Z179te0mjI2VkjGDAhVrMqTPMwXhLthLkzIcxgGhg9o9bcB+nuSFc0/jYc
ehuy+H3UD0oe/+dPqBkMUXOIyOorRpXxT79ncKyDNK0BH/tn/dVY8KCRXL7uhsHO
N6uqUuFFTe57c9kp+KAW9WwvHzPP7yn6JLKW62kbdN+BE1BvZpbsLVoFoMVNmcbr
gJbnD3QC/h+0RXUvTs5Da6PHDOOz3bxWOzL/swd8y5KC3sXAT4jAuLWbtJFqoiQd
a+zuA1tzRL1DWdnoxAYjX9SvSjDDHGy10CFl6pEF8m/rQSGKhdV3GTviagTEjvXK
xs2zSfSJIcJagi55TvQfBD75nPGBr2EjBJzU/I4Go/qn7IpSdAuNIXZfZq/onG+q
uykR9cNIpEri3Rb021oqmu5F2LLghpDsP10JbR8Y3L8a4xqec8FL7mqifhlwCU0M
HTsbqWE0L49stO3232cWxFUCtWobXryXLHcykhs+xA2ojPzUgwHqi8RuZi4rZ4Wj
Ogncin6dEyA1/1YhLacO0w1nLLGnWBO3cr47REoAIh4FSV8Bv+gwGJEYsKoRZcuC
KiOEl2Vp3ofbnDl8wb1Zjp0CDGVB6ZvfEtOuGKKTqfTh3XmuvcwQijgeGsoy7tF8
6LkDqndNc3Fhb4i2lh28AfybsC4rEiaDNk7keDItwF6QmpCpyxA4tyQ1A4p67DlZ
9IuhnP186bmvv33UuJx4O+j2+jblxP/tTS0FW8c/E9dd28GhTbbdIJ8DbjtRhMOu
3r25Jw/1HQAufY9cl90oNjNjCUv+BaPtZin5zGw6kRYX9LmWHENwdRdPyZzqi9Hd
9mJFw57vR3IYFybsMXBaRwlMqD1s6V05PXtNwEesfJiLbX3uAZ7gfE/SvHzlPMhD
zItEIRqg9b+GyQIXHbTB77vHwigd2VrsrhWJ/APKQJmQlf93DLPIcq7CPJ9oO8Kl
/rsqqFBB2RY/IwRP/JjOTqkNbAOVEsQURG/Wz4Dm5r8XK+JvR5efTDJwm+ZHJzHQ
bMet399zmIEBvMJT0hIaU5PwmxRfTs2QhN269LVPDJio7vv5MbpVv/suVkWH1Vp0
Gv9txM7PIIIftRDUN+0/Umh2gjgAE+nn066lfL+3qTmusrTOmAYga3PZdAiGPCm1
fWTX8uhH4HMYuB2Y2AA6otlBP2FWSJRG0+9O6VHt8mUg/yIMTH0iJAgBj+gJTAZQ
m98krjJbHxZafMTkl7mUcVdioSMMlosnnFZOT1dmrtT6r7O9S7h1EYPubDL/3SwC
iQhQN67ZcPnQplX3whadyHtaC8BZeFXOtArF7dWqDlqqE/srK08nI2FbqAW4mCkd
SCJ6xiY5yx4l79Zqys+j8FtVDoGA3ez7eRNyvzTYMYHhDBsvT+sjRfK0FUyisj/b
f/d9XV7Rbj7m4h1sS/+7EFYxd44+8G8q/jCXl776V0znF6ZQr9lkHN/tKkx7nB0E
T7Wen7fkHJT8spdF8TVHrK4p2zBpUgoii5lMjZw+eXxrh8G4jiJPQy3wgwlVVe/n
wc37dOhxtSr+e7cInyMdVsV2K8xjUSXmSfaiuvMRzMKDP/yn0PRCeq2dP4Yu/o/S
nrPvRtH3d7GKgcYm5IXEgCL5QmEmThzn1++BAjw+lfS5UwqUEtuhlDvgy71mFFfZ
HTU4RcedpN+qiVp5tS2ADRrQ2DviXumcSngm7otxIDWI4SL8E2OqrUABn/ApwoKR
J6ylyaI8uK3rr06a3P7rwzO3ygy7cr5oeAjIya2AhnkiONHYXQmBkX+mpO9t9G69
nwHmXZP5JD6eyOUOBMIdW8Rs8EFL7Q0e9obcw7pOM/+WliWvZhowhhrZJh4DC2Y6
fiHwzBKbEju1XZ0CUwMDTRwPUcC/2toAxhcmnWhve8T4zjTQvYji8j46py/q9Lxu
04/10L1WchHcCZzhJXIev28/HYPrG7ZsZ23HttdkMiN6HIO90f4/qDayP6kx2+2U
hw/qo9XWikCPExhwihmX6W21V3H63g5EtD3bi8KHz85gJP8B9BAVontaVM6I5Md3
Hb1tjzCKmUHxA9ahKbFKVI86rxehl9OBKV9Yoj5tNvOGJX7gcwBqv1X43hbb87lt
1mKc0tijLCoG1mnjuzTdOUeYbBPyljO3NtMGAQYvUKxgy/qfN7HYkKgjG36Y7yx/
lBVv0ifjIi8YNngHSlcbf90YOXrp9o/1H7/x4xor4Tv9lAZ/u/UYhHnEsNFWIFK8
+DiN5+y87zbMvD/xp9yCJqZkJQsPB4rRbgNRfhGYeucOPcy0zApmTT1k3b/yOXP2
mzoCA+Yz9mlREGOudf2ul1KZZA1Z9EnkFrouS4Jt8iAvtkn2Df8vUc+1TtHcYDm6
gBcVznTpt2iw6VBd0LXsMgaONGxFdiD05Kt1F7xXqdBrDYdPCaMLNZUzhrLJmXpv
UeBc7d2clE4xPqLWoEXBM56muxpYlJc+kNURGfduJCCEioc9qsuotw4qWg6SKQ/0
7GCOsD2mqwG6G0prUeHCLUQ62x5jysRw6KaPOYCkD+9uHD1G2Tghx5cbK93LHlfY
LR11TUWFrw/5lD0krnt9QnlaB+xktgAXD/xBgAizQaoCzduWNeKWhmzXHgG9PYB6
rlEFUM0LBwGpMM8QX8QP6bi/Rjy9sDrdrzTCSOEySbYM9IUkDhcPsYRwzemlhEvb
M5SoqS1xSd3WM/Gv73R+1l5jzpcJ55jc21P7G1XmEopy6fPJCW5P6NJgpuIojHRY
zCVM+zgob+4TRphrbBZ8mn2a1j4XL6/co2/on0JKIISOQRJGC21OxemAo8CCUzsR
aGHaJI1d0qN5iwVOP5Jw9i2IR3W4Rt3mfUsORwB26sGGPWNOMGTufBh8IKPSIhn3
C5jO0/5Kzu4zsvuT5FcwmXE9Ri1NYP1U6SpkUCAwGJ1iZx16HsaD/LB20G1xNPi4
XRDloY7GLHRd1yhcS/7Vl1ZrLx+JACcxQe3+t60bDFGLMD/KA/tnCAivekmkh1cD
UvVWeJyDemZ7HzaIzorjfbjgcmBIZ+HRxSGgfdKWIJdIiU+ZHS5WXBtRXN2VXDep
3VCBsWq5P/oF8iuvvQTHpsudqMkzLE51U2L4sLE7a6DMGq5tj3wT0a+e5g2KbuEF
kfEvrdGK09kaOHyfm3KyV2iIxeg2DwTSswJGivbU30e7rW8/8tTMi6FIMbXpIMew
tUP0G/1YmPbegGQk3Bn9Y6GhK+8pcs1iqQGDZkJ32upFT7gj5h4CK4Zgvn0gi4f4
haYzKa3za+Uu+umV8gSeaqh3wKBwlGvSLctpjVxZiUYOGw3qP8G7mNvz1Bsv5Sfw
LmIo+mGiVEOqghxJKntykz3WJE66EJm302wyUtlQ5vXPLYScAdO2uhfbEW4LIdTa
YUB0iZ3hD2jyAIZzDjNZLLV3PZ608XlZ/hAWr2jnUkAovOLm7SSgLLCbSnQC4gGD
qEToljiANq/mioTurH8Vrc6cIqqCk+Hcc+xdXBq+oP8rehk4/V6fOeVx7PL3e0gP
dLZu5S+2jmHu/7XsPJlXrJYTTQTPZIL+DVfKSJFxygSwMQ6f5NETfOqqFRuuuIIg
4aGsOnK4RO+dr84hEFfkKT+q3xvK4NLKIUWoMr/bOa+PgOxWwUb2+vnQMun78qPW
U3D4kzv2PptwsCW2FsyNL+islHViQYHHoPpkD8XbWFQ7vmk14O9TJJR33c0WUr0G
AVn+nRvDEil7fwFtNWJ2XjyKCnxt0oz8mACzPn3nzNssjkYlD5n8zv7tN0zdZcKy
91NaZwjLWkEZZslEZ4jXytTn7/RNkY6Q/ctfMXIPu1rQbebEphRDV0riknSGSudZ
GebfLveuEzVpDL9D3Z/Ya8ABGijePLbqtgc+ZFa/vN2rUUhiTyQ4zi1tfrZp0awp
x+ojPhGPjpplvDxU9MLsy2QYF8dn4dHabnike0qdBljPlvaM9E2TuJt6QxWwVUzf
HPES0N/Pg0E1+7JsDYjKbU5iI6+ygjvW4Kigzy10d+GLRBu6BcF/Ufia1zgnO8ad
vJwV69MYRoZvemLKC35ZHgUChcL8v9LENrRYr1jm4IHkBXSNAqLbyDF6Htnn1UP9
UXrYFxJusANy736a0rZsHMeKvhWck2CFawseGLVR7ADlqwp5VS7Ggj2RxyoDghfi
83o8dvaRsCZABcnI/mhYSHWqBqP5J1eiIMvhM6aNZkrFrwUktDEt38pp0VnHS8Pi
d7QsVYMetM53jjBPdBbgwS3khCqnV4yfoZmu1j2B4Rh3o6Jj88QIFVBF2oatmPaI
NufVRVhPDT5kS5HuHyphiGYZo2Ty5x0R248zk5vF0IhyGcer5VwddnyGLSWH1px6
BLFuuYA5Qf+JhupqPKoFf1irjw09HOZPRbt0bOL2yf/XfMGLz9tVmLG7isY1+zrY
pz+mS6jmRIhqlz6lZJ7/L/HtuzlFldE/L9xTufIm5OcRYc2H0olfyZujwyFXAYGk
Z0vkCmYC1vvcOuhc/lVeoBsltAKt2M5kff0leGCMs4C8UWgQCKfmqueYmerbdAgF
I+oSlmzSqv/EgYoMNzHQmQxFYOYxLHJeb8DhZP5O4dwKZsZRLZsg6hqZgI+XCUts
4+zuu8J88b3LO3WdH7SNvnWEtdxWpJ6usddMOxuGzxHrdU67AxKwd+55BsYTTxoX
8OiDIOX64dwPug0R7+0F3vU9BfN3FSru+a8ZoBOeEIXBCxiH/GUggSbefevFK0QB
GHEq8iTUR7/otFety7SGL4TuXn6NZT4qxPJL2NSEouMdYvsyGgmLviBOQs6nSbQp
pDJKCtIKwUmX0YVZEN3FEx8GRIm6H8Iq3Lf238G2CAFhWqIR94wYeDjbibKZzFaS
RjTQUk2eXoOSM4jEL5uzJw4gbk5htYpMUl/FeguEAu8qIGU6eL48ZWPBOlkkWwNM
EiySrk1KcjqxELlG68IWjZhZX58mq2p1L/okV5mIqSexzSR8wk4PZFZsc0wdGpIJ
CaJRwA6++CROY9jjyJf8kKvGaQ+L9I54QWSIwR8CbTQarguPyPYbmG47EAhEaty2
0LoJPHoL3f2kCY7u7RYwS0Kab07TxltSefLcpaBO9cDc4yCcxPU9byHaum/IHAis
8L0IV/zWQKkxFmQh1AqcpreYwW6t/JkPSHxbAtwVU5umddc4itWlECkepQ1wBBvp
slBQEtUoyyEOk2NsBmpVn63l6uD28amYP4XwKdGp9O/SHYfW7FqvhGApRZX4+LLX
y2XZyqreQO6Qu7Yk31NcI/2JllGZWediTFelsPA0WO5T+g7gAR4sVUuiW+KGAlJp
gVBN4r5ESu7T/DLPGnFOP1k0WkHLqHGPB2giuDMtXPH7vUyBf/DLTu8UkgiF+WJw
EjStLfImr7/K3hJO/8qG5HuCO5Sb26TWP8QgRbUuGqNAOazzJN+JAkxvJNW64yUN
WdDNPrBGiz0/rMaydMoOJzooGMmVOcn9L/fBHLMX0inANdBourWOqQn+q6HgdIh7
HhbZUjwVg3E/rlx+S0dBlvjYU38X5q5hfweJePS1yoIn1hLV/Y6bPMTbB1fS6dks
GdExDdgej+jtIbao+Zs7CunliPRBZU3OyoVfh/6xNRiuRWKskwI3Po7sk3wNTk0l
osdHhdonVavWdbeT/s7Xsq88+uFqklCWimWBRzHQEawYcUNG4nyAYbdzmFKmOt+O
7ozpCo+h9VxQOu3VBGfPjlbc9XUKFEybz4SJeqv0ztHjOwwRViK4XYoe3M2A09pI
6VA6ePX/R/ZVntPJVqvIdrL/DPNdvCV9jMFRxQc+YxMM9pPlLqg9GmG5LW8sirkY
sqOj0QKz8jPkhOv2/r64iDp9BERO9TTyX1QloxBF4pnW/jAJnfSWvtxu7U2/gMRv
d2UrWxTG/VOR5jbBJVaYorpsyHCXpWK+5Vnai3eHpTykIfEuu0jImwK1HSIFVVai
kZTGJ9TfzZDD0ovZz1gxN0nyhHq0GZRrmZEISXEd4iAH7ndfpOgzHTBpBHxBf6yk
y3xO4aTdxTt2vdTA8Hg0br2bmc02rsqx3BCMu/6aWHhhRUyvF16YGrShTUBuucT2
Z4kr7P2xjh3No/xtKS9KwnsOK2w9dR6O2N3RQ3rsLOxJ6NwbcQi62uGE+eYlVUOP
ajWuhWmOgxzXwmyHuW+A2fTKg6fN7uU5jLPKVnzfxFIOAgxKQjER+VdHsRYwqFhm
zKNngkCzZa+UU6OXPHbAsCXVlrv/9SSqoZFbsq0g1AFlIwwnadGItdFqJm8oHJsh
Q+/pxpch6N/uyWCDNR6WuTwHzhL1XCibdCCK3BTXd++RLHVFMtc8WSRzfR2WjhAO
Hd5zgDRnRtllnVhr6irCPeGpROuMPljyatPrZ+NDKEmN3Ch6OtgFejxX36nQoWxe
oYmd3n7OYayPWu3kAG/noDTec/YCwocuyGMratcYhOxBHrJskMk9Ux00THJ8hfhM
fv4ZX5ruO/+Za8i3iu3IXT9+Xeek07cy0UpkvC+eh5ScvCbXRph89uJ2uPASqqbk
o+O6NF8eqYdqNhHTglcghOQoLde7eRMpaS5ItF/5d6Nr3cWD853gwtErBBZic+Gj
3Ak7wFiuXxsaR2ELsI0TgbqgesPSYq3NHf8Ouj0MSNky8Wo+0RXgqk3xFPvs7877
SJCDVy/KP/yvwdNEgTV2wM770v4zghhN9FvW9MxfNKZSa0t7ojicWbC7MXA8tZwM
CuQw+31OkOY4PlmlxrsuMFioh3bNsj97tqm1y6ki3zJV8ilV3i/gbMV9h5/ahe7/
UR+emtgjsr92oKmXyz0SgrvgFJMRedrPogga+zz5EFzZusbDNO2CTaucOX+KfIvr
tQa/4M3bIcarEAB3LrmvlRPD1mAlT8Yspwuys2ff9PO0ih86FAU/pYflZTeUrE/m
eCjidA7ngGiLMVNsDun10fs2ukTwDUaqTftlZe/4yMtN0nRChreOil2ensJbPzts
87ikrBuvJwqVvgj0TBNSP0ngSGO9ryy8P9g/mn6WTVN/ikRBZcEIALQTgEr06wfI
/Bi6J2FaOmxH/kw1jDmLeVNdj3HXsTCVFt1tGgFXn6PK8d2knCtWuha8DVTUQa+D
ThuRwgX37Q8PZ4vFF67leszMGETxwc/ljizRPRhOClQPZfl6NHuqZRksmYnFWMF2
8uiHhlONr2hCn7V+OtiDNnGFc7kM4lkZK3tI0cSu7R1vG774731RFZcqh2bKLeg9
oxdXrfolYjyuHVwCIgyNQbe3TYpREY9W061UDinrRLUjz4aprWKh39phPb+JKivF
h8etqzfwqqH3ZvJ+pd72lKKTVHT+5wFcmg/DqJlT4rIhl8vL2UV0es7TnEwVzFHM
IpaauS1bPnEnuHN4nkT4Ok6Cf2aIVGvpOnOD88CUa3qCAS+Dl+ylUA2lz7BEiGhG
wZD/Kk4h58/H0wr41ENn2+M0tgHjhV5Y+DR/dwMF6q9JeLlckOBZxYJGVwS9SDtQ
rIBYeEbhr4G4W3M5ZCU0xp7t2AIuv1hgsO3YhNBIcmp+Idwx4kWzsfSc7qj6BhnV
z/CdHmQ/Nu+5RTW+vpC7WYGPJ6oBoq0LhPZ7pKFUgvKXvKJ3Cle6I6OrOFHojVQz
KFUu7LT9R7scuNecreBOlJPwqTMlT3WxehAQJqo6wxdSwadgIVLluACXK7v4ONmQ
P97l7tZmox0Ipg8oG7xnVudu8l6s0iSPe2nP4naTrTCmnzdj1bWvApsMlWXyxwWu
YQwDJhY5ZYhQKv1b3UuUs64hB/1ezlI+Ai1BxZui6ou/3qDxPBMjk3jq3jMO9f2J
bnUM08qqblhpMrDMOL/IQRmnEtg6sDBac2m2iK9AYwjaDpCaIsj9irlxhGNWrdU9
kTq6sg0ltOcFDv6WjmHNtbHQGHjgB+elPaq/AcbORCmQusT4ApO+hryMcQa21cAK
60fECmyo8o1azflejyoX4qM5wDrpvqzXZV4JN0eEhrffwrDz648Nk3JhdyrhSaLO
TQSCNb2pLymsGYYSXQ033eIpxKMKQF61a4p2cx5/wzyexWFjQ0T55C7o7CTMBAeJ
Vh+atJ2nTjQR0bxByhn9C5kiEaIZFyECgMqqB+7Vs3OZvUN70LuXxVV3eaeorOfM
Ft0w+ObfATkDxe8XajAgf4aras4IuybaJF2ufWvQc7dVObo/I2P5F5dKg1chekip
+8VP+lLkUovn9N/rP8UaQDBxk9nTH5VVI93V8c8kKSQBtTJ28qDCkuNr/SXG+AYh
9yXSpJbuMlzDFMFJwCtZ0nRW+DiSMVUnRFVqXGaEAvb7GKLuXf5xVdyWQJIB6qrO
Wve5vUf/eHuY01CN+Y87QbegeBnqG+6vBs7ia5fZiyG4M2OTZJ98c3u3YmMu3MKN
aDjt/TgfVKCvCqiJRl+4RMk+zxMCkAUKhsqT5t82c1/owsd4vGJrGMpvVCTFGeAn
Bs/hgn//pJx4GjJzhVwhWqgVPNXtnaHk8B/fNJMASCx/IQPVDLPkfgehS923bNLH
qpG2MxPwDlYvdRhYwp/N9LIBM3jhfL5FBnOZhAvLXar0Ln0QDjmL0PP7hO6SttsU
UQOOtUVR0kTP1A4p6mRTQ8Kf+lPP89mzx42FISZoZsHiWJ5EfQlyZoOGZv1OaWcw
28+N1LoMbzOBw9O8m6VDt3+1/B7/JaeNCzWagaHjam9+IWDMdtmlG30I1iD22Qe9
m8W/G+GBklafgtOz8MfPr7o1R3OyXvOZTAZz8jx2nx9hL+eA8P1wvr0HbxJQM9Ui
lmp/n9mX6g1XAbh1o8NlYKiKlUDFTqapGpRLe6xm6WN2JOh+gIRxz2S9T6rmMUqh
HNuA9i/z6pY7cqVyIESTgZUVXOP0ARazphRbUV9MRw+c86UQF8f8mWntGc0toxng
yhlJ8D+Ep3VtE++t/epMPNeOh6O3cn5Me9iF4Xv//ZlbMtkmfm5hqdwgAwuY1bC9
/az6zGSjxqN+erqXoIcQHmPlkZGAobom4qAY5N19TlO0xH8UPG9yblnZi8nvrX+W
cKhiiig94pkdyeJhdrXMmyjRoo/Y26/l9zOBw9jWl4xxoJss9qP8dN9EeRyUI180
YFfUAvYCqhhMxFne27qgyeNyA73Pv17H7YLqG1aiR3McRY6L9nYwqQttI61bVB8U
vjCuMYwnOUBvkdaOWPtgPojO3smkTHIYc7YOfQnci4zTmdtfbQYuTAUzxzEqdW4D
NEnB0DbNOe01Dcpd7TOGEk9o2ptChHLZ98BFBfun8CEcvc6K0JeGH7Dtt/SKPkgx
iPTSDTTORUe6PpO11KhgqtRTqKhHV7eV4nJPJIz5hZrk29ELEiSG/ilftDShtmbS
Wvq3+uPHiAeDbJbV7tzl7ukPIQa2KnN/wmuP8JRD722ise/cq1XhAvBBa5Pb/aDl
849LaZYgYTDB9EdNCenJY6FyG1IYW4bYW8sGcdvbI46L4FmP35TUGCcGPKV2fdca
V3O7RgF6a5AF9gH+L9tn/5AZiEqB1DTR4u7PwSW/zrOWd+ISvSbSEWT0ihRhPC3b
D96/s4jWCzhI1JQ4wvqDJatOmEqFQKv0I3BqtGGTIx97wffOR7b6sL7pFNpNbD5j
tLpSB5yDX8tFxRVRj5eiRE9CDUfP09zQa80ERFHZZsYkzUyLi/H0pne2e1q7+8Ym
yS7QgidlKq+kjwJTtAlXc/BlxkncD4v1H3bQDuSJPXw++baVph0id18T1H+vkhIo
Obq+l/TLVVTJ3llm7GTbJVjlJPQ8GA13yUe6stguN89DRwfiQvibHG2krjB1PpbR
WyrHHf1VQlSwoCygmTCmloJc2LD7yPwBw8XYMYLPeMF1LDDWCo36uYvoThpWdIRN
UAL9Vb+co5q98GV1PONEp+irkI+nQULejsVnHHFLi22fvHzlMmZDbS3r4aAzY44n
lBFT3gGUT5uGQBXNfJaALtRE5qx7aHJXM0+eKDphKcO5o9c+bzigBEjbPnF501fH
eIJL6H6coMM1CZtbatJ5UAuNCuaHjgT2yTAa+bj2u83quKUdOtUceOBQoNcBWktX
3ZX/h4C6D1ZH58lBLlkEtF7OP4B4hAnh49XSBndWAcj2yQ79juikGJBptvwudd7T
HnvS/fzKzG+ajtNpyWOzaAuOVFCpMNbTC86Qx1TlV6zpY7phgXYDJoXxrg4YZJXH
wWboCUb/VMd6sQTC64JrBFU+Iwm5A5mip9dthEB+qrAxY53hneDfi6uFfQ9BhGPa
x2Aqn5zeOMxgpcFwArZIbtPvDdXNB+ri0N1IEgFLU0PV0CMh7ZxOStKLnFv0q7SU
JAo63UyopLYkWc/9e1/+Sb/2q/YUffRFCdE5XNrgVmBpk2qxLdeO5C7BT/xYCDos
O5z7H3L6A/taKKMjdPJOg3HjQ7pneA6qwRt0eGKThVtC5j5REmYIeG2dzuhLSUxU
ZvHeS1j/h/xUuep49LrQFhir1wJQje6d2BG4bIVrob7hXkCNhfOd4UOp6ZgsSzLW
Wtf2iP1n6Aswtmesm4jbpSlLsryIfasVNnStXbP9jyTq2G/euLr1q6+JmY2xnlIH
Lt4Xfki4YPjAQlI5hQAY8NYT2EdlhmRo515zafkjcK1EG6mvXaIq117F/eS+PSZN
6aV7cmJJArZJMs1aLQwEHBdASbnWSzSMy5fQxZCjRzI6wbBARppzXJOycomGDcm9
qBUyQgsjZInShWZTAdAk59ZIYQObAWRH4xoG4+LlLBcxGmZX20OxWABXyy2qrXiW
9Q63AAwbwoSAu+RJyFNBfPYAUMPr8l2q/veFyVyyFb3AX3RfPdL/kFQ5bxN7eHD2
gPsI7VshSw1B8RLmOK/F0qIRcmbTwC03+MR4+zzZAIQWpUk7XxkBZeUXYdytzuVX
BjwuDHQ2ODHSnsBxufzJJqSOcWa3ZzIKP4WOrpscJ8L+YrU4m5YA0CoEp8RwNCuN
RaB3ydGC5kEKEuyEt1dqVe/usoQx9wS/gUlPCmg7PggpUj5C0KlxiQMyetjVAeC9
SYD7fcmMNaUm5zETwmc5UstNSJhsn0s6O3HihjiJrJzrjNeXQO8y6bdFXabPTfPs
fNStmDsf5PVyDbu4Mc/zaZVX11vxBAznvNa9nvTU0VNAtiiVW2z5dm1bUIjRkdXe
3VxmAsII9b6TmozFv/QdFpqfU1IDIlGAkqbS+DXwRCsipZEfJGYw7bAi2r1Igahm
/G5whh+WP+ewxTIMzdeKmPgUaMoEwqMhuT1C5v3cZ6gg2ycevRkp8dZ4biyxHDyA
53lK1l9g4d+w3nBsHa7Rjt61RZL1/aPMOoSPGqB3cLFxKTJaEV90lFxwXeoz80bg
J1E6m5NZ1ikoWcDFy8fxexstjdvlYiL6tJL4lgtoSbJh3cJW3iq+mPUIVOAcp4Rr
+WecZmVmmWQSoy1IQ8RZTLqnBp8N9mL0Gm2bItG5JR/+DF2INpca4KCzVkIRj4J3
Nx0qlOEVQCAqe6SaM3nNQCopPDt1ER/x5DbH/VkOoiFNqdN6CHrRygXJwhNHf5lT
kTfwl4133EeqG95kVTEJThE6NZAAfNEw+LOANRvUxb944j5HdIWgTeT0JDPCA7t0
pnLch2dUy1cFVX3MS/rCpjF46+w9F7P80AxcGq4xf3KaxgSVFcpuNR4Ehler5dmU
DBlChIwKYOTaJCo0axbxxkea2PHRmsOGLFr5jST7gE7ZZrH1ykG2olaUxuW9HsOH
JNyFgwjqLbbI7Au2IX5vCSXMTw38WN56ftKtwNQUoYPDCgN0MgDz5rPgsjMjUO0k
G7hXlVtBWV6RgQPIZuR5Jmz6jtPNPcSTR4q5IN06RVbyq1ftuiM0HR0xqvTMGN+x
XT0rYk/peLtTUr1Gizj7SrdLVzlQURydGu58m+L2F0AFPf6c5PmMSFOhMwhJgBNG
GySKTjEmwVXVaf5dktsJnXEnzhj6XfzsKLNP5fZvUv+fa/4J3cl12nlG6YpWYJWA
cC3Ijjk1CpmfKtPlEMsr6BkLyAQVbimAwnOpOyGSad6M3O2BubVTBTifnevIX8eR
ima2Pw18ufJgD7BKdbHdiMX3lBINechGQGKc4+9jwQPYEb76LXSWY4hBUWDl+Sz/
Xn4ipK1rW754cqniwcGQSgCBVArEr06GskE39MEV6rcPgeMsXlzTQ/Wf/P/QtWxz
IQ6hiiUR4Bc76DGvnOnI+46WdmtiF1PIE9NeuDLz7NMGgkK8JM9A+WNMPrcz2ln4
fTsSx9nHbMvo62kIbDearZAnHVubdCXBZl211ZExzh1fbH9FrmUcnW7ypHU0U8LK
76HHhA98Hfyy3EXcHPCOgorp3W1+fQbY1dBvGxMQsgWGBzEjhk0pl7n1RV+kIqDb
yeVRz5CHbmP6xfTF0sv7AV2EQxfnCc6+N0azrth6LnoOTiM/1/CMaGEgxFyMem5F
5rtFbcjTxVf/UvUGR7K1cy8GVhIDwqtSkxncROGmHQ1mZVE7wH/UdQB6f8Cq0AqF
dRGDLwGaNh53pQn+BUa7yEkEMvKmXxNPpc/12zLAxZNjs86GtFBiQSH3F+1sJqwJ
mYqT9EDMOwo/1ZV6RioqRU6mP1lvOVpyALttqHxvbAPM3yHqSM2TdfHHhfbcjCCR
+HCQ7hoZig6+t/AqJs+jPMU74ycqjTlucrQeRG8Or+we626LldVE+y7iHa0Bjlnm
zZ7y8n/JdD9bJhfu/bQjMKuYKu74fbOWJ7s8jOnVQCIMSMeSqTSF4pnCAM8VebVF
tdyQfDp54Mo5P1xZKefuV5VftOPAxMPtBlbub0GaWg+duq05FGm1oCgKKzqg3iS7
enKtu+hFI+S2fowKKjsv0NTt3EWCEEaAdX250rr54MoZpWfVkihqp0h7FmHESLhr
SyqvRQBuDdStPhOwijhFDgvSQwk3W3ssXTUtvgLndjgGQ1aGlsD8E4IjbVU1hJpo
GtM99VCR5n3PE7tuju56vRhIItYK24GsKcUYQs84K8xb4/o3IOBCuqc0VPR8wT/I
hf1c3WmjcELLF2veDpOHtuPcQMaTsjTUGEEKkzMOuhj5YFue+XTKXUajpAn5cnWf
fUe4WtzCdQdGFn/FY0kOfWKykbID/YC6od2alBI2c+ClgVZwSXl+40R9xdlRv6oO
4CWYEfeso1ssLCllEu/rF/cV4ltoZRRG9GFnUx+31aKLhA8+b2ESSQ6I33CsBAy4
pA61xZIhiihGWcPkA33W6kafLAqlp+N8s3iz8Xs+HzGpbVj36rGA7ZijZUlJ7XVk
mRF2Y4EVA2Lv5TS0kRgRon09qHsCiYR0ITfrGWKHXOCAiw8/ApT2VWB0dDc7pt/W
N8cTHJgPuqC+wfOsSNlSuVdYisqpixH5R/o3acGDzCNbDQmBGS3tCNSpEImOj8Zt
kAsP6Issq8PJFLXSRwD/1/Yl3o9r5qcTSrWGyo2j3iV63ZHSePICuc8B07L0YO9V
9nrjAoB+wvZ8et5E//GKUdgPTY0gYpeeigEc2KBLOkGqS1z/vZ4PhQj02kb+kVY+
74DmVLlTj0R6HNVVZPiRVSK1eFC7SPQ3yM5lQnqFkvU7WLOBMCeH4QOwQdtaIddf
qXLH7RofAp4z1J1VdAr4u2F6Rr1mLXJsRFCoIUA0pX2F8begTyvmGAs1DhquFpIj
1gPBO1pRJXFkhdbv5+MUovIjCP+/si9PsaosshGvgdIXSv7CmyJ3cfuPWlwXbyAO
Tal3xceiV0SChW+FZc+/57bg5XnF4BGKKxJO+go34NkAYKLr7vco6aHJO1ZYh0Rq
gamWkokfnCPBS1ZuyzOP3uBDOyayp8TCYuwJVd2Ef4zR/bfS+UzysoCdcqh4UNlw
ZAL/iiQef0hiE3JGcie3Aga4Fcr8bbbMS6IDQNAlfNTrRLyx1acsj11XdLlvAGpQ
N5dvr+96YP6p1WrsUFZaLZu2xqap04LsSBxY1Hh4TLdjpYEaqEZSECFsQSvkphPc
5cj1XVeZdzxuPTvK+PRct2dpBauITufxILHS7V/ceDdgDS5kQ/x1idp/jjRracYX
24iKkfrPt3NupLzLxIO6NAFdmgQ+Oxs3GYxct2Ke4KcArU6DDOAbpUFaEEGdnMfN
f4o8N7eaNa8cKiVFbZZFkMRcK5OGQdpP9BWEC65MdVOMSbFCrKlzO3u4Jxa2mwTG
1ODN0wZCFJ9oGCH+XognAKStBsWgQMMp+Tt8/y54iXiyM3EPvdBuc0tGJFNxOk83
akKvJi244tVbSEL3lQCf3vrvwf/spqOAu4eXxWwAR7ww8UwsQ8aURkgcNUbkN0yN
u6F0+Nyln4VQvTf56YW+D+VQ5VYSmePcDK65715PFtLBhuXqytpzfjt0y8dmMJH8
74WdipOWpjpUFwm/20Tdy8KbXw4G4xMZ7NltpFThokchMNCHrCnaJ8/Cb8FppTR1
TYBpupvI8Yg7US8plzl2nsOeYjwAlX7p5+anl8DejLkpiPBy2/jMEDd1SR2CZliF
qtm5UKdxJee2N9yS9n1ghsS+g5A0GEjhguupl0dr+Tt5AbzzIJ7iW5wZ2Z78omzC
XTOND01zIkyWkaceO3NXMjDeUlXF98ipwXgRzmB72Y2LO2Rso6IWDznMTXEJQ3Ud
RP2tOcLJL+ROlRLUZJenIYiXcYjLqyOkumriUa8WnDGP1zpZHR2mBtt2s0j6Hjr8
laWHU5iY5EyBK84U8L+XslPAGlti43bJe/4t5eZ+GVlfdAyws+Gmf4hhaEZpdQiw
wimpTHddT17PLQYOHTfNr/5tOes0CwG5yLsCJixkxpjeQDBmrVg2QN+FTYHggaXH
3/oyg22BREMmtZxU0tOvk/XzseohzbGA2UPgiRmvczCcFbxXGlKUNuVD+f43K1A/
rf53kIgSzuM8BPQJJl4l9Mp0UCqxTJ8pm7xwLqZpPNGIAWDkZMdW+D7VxCMxdXLR
C7zAKL3lxTGz0VlPzFepSiQQXA4SSangG+T+nga9pGh4wx7KJoO6YxkLkArK4ICt
0V7qkn6RRcgJwh4roCPLlbiz1j4RYamu9SzrYib6pZKD4cPLeatJeiarhJClGwEt
96xAYa4XSVWclI/LsJw07D58+zs+Fiz6hJMJAzI8A3LK71/YG4B+CiyT7kjD7ef1
+Sw7SWNqVEUqYWR9yydS/K7EZTsFAAF7AqOqKcwcwrYbxR98xxrrzrsNQK/jt/+o
SIjsA46ZFC3nOhwWMwtWwKTYIPNZR8bCHZ7yt3OzFXFZse+R6RjGmzvhQWOlJhsu
eehz0hlAFX8zAGFAXJ1JXILRYzioePMcRZzK9cBKsQlvV+9fwTp462zRzRhuqjhr
r73s2PWJ/qDnLSkeAriTVbWjhbzai3yK51BWHk580LSxjDDrDlu/ntJNvbcAoMvS
X1bI1qGtGd0VuVzdEqld25QJIKiqiYPxkWLa7bdAv2ZPGBTtzml045j+QKYnbxft
cN18rH29t4ku1UyFJcuiaovmBwzfiKs4QIVXrJlZ5Vf6ykJ0RgDdfQBD6gfyPcnB
VRMuqSVXLBzpKOHj8k4SOwkrV4u6tffIu69iZFHVxMdLsxyJDS6dLFgImGZ8KxqY
TJ+wrHME+Y0yKbkvP29Z+gZNXBGuXesNzXtHfW5fQwqiWLT2I2WLwt/1jEWhzyXM
rqw6lHIomKgzl9KXU1Vl9AKwn/Ci388lZm5EmztFQ/xUIBhJ7saWrEzhuQ3f8JQR
wbl71Ali3eg3yK8aRnw/CYAFq00Crcbt+7FsldI0EbcvcWjAzpzZ6lyBFcvpuF1V
Z3FzFjA5DxX5DI5bYex6SmCMcqz1aDai3zlz6r6yIRF6Q91vbriDqxGnx2+s76EU
`protect END_PROTECTED
