`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yswcyO/GQck1DdNhWHrWrfEkSbiK/nXHAzEIwPKYAliOnkVPv0+4KRJFMb+6Lwb+
IhvzRLr/Kp3UrvSNUISXKrEi9QdyXLTdoFHrLn0tunjXwtSHWGriFU7nw/R8al2B
jTXYNTLkZvPgRVw0eXbXWks2Q+9A5SmNO2+QCJS9Q1JreOs/z8R/XwYgbjfnh5Rb
mvTVsF+Mb/kbx8MdvcjR+eHzRffgkWi16xqcYbpeEAZegDxAJHEjV7x+4c+N5Ugc
Bc137a9buHYihtOJTdqVDmlEV8q/PyXDAB40iOvdtXv0qWBwPrFwZkdoudn/H9mR
nFav8Yr50PpWjixH8RrafXO0SlQaN90uYEMRJb5/WHBYBQAHVQALxQLd2LKcR+wW
f+M/DTgONyMHBIGBkv3WcFnX+8gFchFdAU4f5PBB3oeElpbvf9JOlYNOD2aJR3hm
3ZA1dKQqFz+8Ntt8Cc3HERpYMIC5sVI/ZRAb09rt5WvAeepmdfsiZo6CCK69yXaN
`protect END_PROTECTED
