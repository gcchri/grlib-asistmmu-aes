`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/kcdcNBF8y9RN3GElCYy6G1VNVJgGe8yxw1XFGxAaeoJ5Vwy/3OU2lwhlAnffji
FeIX9y0fL00Qu9HRTdBvTTy4RqcDNtR4g1IgWlGxetxx7rrgrszjqzofjQ6EzL3K
XGbQyhIvkml0XlsBx12LYrsI+UQ6XmuEzmzJpQJZIrKy7+V1S/ArCqgZSzEhvtPb
mon9GrnuZaVg7z5u7+B/idDGnUdNFSCxc+36xihTeiIPPlB4hRWJZrj1eUvuiOBT
H9twcy99MqAQzwas5jDDYefgeegAPsWabY+64w5RlYWumBY4B1Ue+p8STL7eZZ3n
EUIGgwCe8/5FgUT+qo6i6TLIgjuhlMpV2TvUvqwXJh8lgNgFC9yzmj8Phv5mvVwi
y/cj/51qY5hVY+grP+5KnmlwG6yxyqNdOGZJK9d8zBA5ydndd0iNvvzf6lXVgWH0
umLMHIp4cEnE5/y7bqx9xGN4G/YnffYGlbJtmp9trVlnqO8lm4b09VDAW9HoVWUb
8Yg3R6IHQU8J+NJ8oaLV9+jBoulfjT1Hqj33TPdwB4+moaNixdWf7AI37aVNNO3S
SCLfp5x2Jwrdf20SMz/5PIQgKGhVQy/JWAgvXOyojXZyFIyjIf7W9XvK4WFNX+pM
oUHXcxqStgxAhxdtFO0j6Tm9JCLNkECqV/W7M1zV3Xsafug0Q/TdrERaJQLXlsZC
fesCyon8qQ36mg9LSbegZleGV1iZXf+iBs63IblMACM=
`protect END_PROTECTED
