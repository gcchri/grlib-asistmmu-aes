`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7uVjuOR7o++wb9/PBFCDezMHWpYrCUknW8NZ0rApjxFZWGl7gIp7vixIn92s57L
+yLyIuK3ahE5T7axGYBUi/vZs252Z5mcS8SHO5RgPrT/i5ateX6jpa/UwSRw4GCW
MpRoq+S3cJ8faOk4QuJsS/dlicM/3sfbinBPqMZn76AxRQVJOlNy8RnMdnMB2Wtn
Hl8jbgrZTYHcIewqfgUJhZPJjTShnoBr8o6yeGH17dzX+yp3vqlYb0myuAag/9kW
NejFQwJSsrmVd9tc/VzceIhK6L7+1ujSwJJULHeUAvx5GaR0gYYGEDme2dUUzMDT
T8CVYpHDbm7mCvnhasmrNVExv/pzZrCECeaKTSDqJ6AAUJiAzgvUrJT16BCVUcW7
yeE1RRCNQ54Zqe0bgTOe5B01XbHkBCCB+lA1vkRxsRoQzxYOGnGRZotplhEAxkCs
QOnjoi31nqpyiDaMYPUi/iSyIFd96i4jn8L2YV7C4pDCzSo1nCA0mGdFhLS0RWlN
Yt7GEQCO73TDzbfNAz8kkk3qzqM6PPyMZLWxyuGtoItsY2ZzYkh8JWFuyNnIRaoe
Yf5aEqaSl3h5B7UMfvoWFxZLpdChqhd4iYXRsRcZnGSHSiN+pVofuq77c1TNXMMn
ShzDAc4YLp5ZCSETBJ+9LzBaS3FmS5dj5ouQBcY7b96I905wz58QTXL1wxKpUZQI
IfyXGT5yKpYwz5maJESnxQ3J+Zhqm0VzEJ2djlg6u81pxuRqFkysmy96ZCbLfleV
GNR70LeSlmPkjgUUnHEYaLc3JQC/T7MruqAKmTGZxpetSjMBVj5bmSc9kGrzz8k8
qVTEMvx9Tw2Nh99UYmgPgGogQECk2N8fL789hE41oYSEM/oebDoWhp2zmFePcu8x
/bI1eQnxvTRRshGkxA4EM5WRCoiiWx2GqhMXw94nEu8hogu7haONvOJBO+70jKMJ
6KCrBv3D+F1nomMKPTyGnelU7GuaF+NPY3Ob2oEe9plkHdqW2ybgj/f7Lbnzwu4Y
oQTh7ZXP/oYX5tkf7YaVvtazbINvWsVsO7jCO+ywVYVrNJGy6x9/5z1WHEeeThgL
Xk1ZRaiNd6b/T26Kz38EoaGpNckYKMPHJztBiC0m1X8LeODxatGGjoFmyz2ZSLZB
iN4+R4Lx4T57OynZr7+j5baCURnoc8nOpQ9PpVy2Xj8IJ1u2gWBy2N2cBIAkN4gB
PJCTiDH4SeMuik0h9hvWSikCJ4eYQ07JMgM95G6CeWmRV/qZS1pG6WnON572ot/V
WrJZKFEBKFmfANlsZrvqn3gJCZI4EIVXeCKpMdbnnTXrvygms9xikjflie4wL5LJ
AfkWyBWITjsT381Pzhwr3tn5jf+j+EWJ3n9OxwbGXf59/p62qLM5wByFu7SJZFYL
ra8k422GiBswZ6DYgxJljGuSoZ7Rf7zppawAXpd7ZWoWUMypatQU5l4dj7firex5
qHdI0Kh6ynWUyzg2ZC+6QvMMMTfBmpQL9kRXTmpdo3eVkvC5/l7EyLIoormRZkv3
ctE9/m6KEaiSjMHBIZzEdLWk1KP4rauRc2Jm5orQicqUQN9FxFaCzSQag/3ms6Ev
mZPdmpYesCBBMSbirGNRhfO0/6rbV5vEeyq7mgDKqaDmhN+TMv/WC8CLSDHvNLyY
viiFZgduyx/m9c7AjJrwdwymlRGrUjijtcgvpNhbJKzNdMEySxB4NLrZZv6MtIF9
SwmGto90vArSNuy6drVKaVc8l445C2YM7UZ5T+GpESjo5QTAFwC9jIAukNQ8fLLH
`protect END_PROTECTED
