`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmoIuc63YrHrKV8Rvr2S2ijKP43B4eplimRY0SkKMw8O6SgTVVWEIkqnc1gcAo1u
Urefe2AC1ZENJvauUnE6ejK0mrrT8OvK7lTxH9t8CaCxqdBVg1v8wchE280igtJK
pgCE/B5J811GmwMo7WZc3vYTM8daarJ084/zfgGNBlCYm6jlonR6h7NK37p4HR4r
mG07XNu7lBu3+xo90xW7gIMDhRdZVraeSVPz/JU9eSnqQXMBKCXxUcAheYtbigZe
VAOZPPNoPdpLmH46eUh1F3VNUSHVXqZUiiieJhLYEsAWriNF3B4fh47kxHpalKsx
int3/7/BvS8Zh7ZCsv5kv1/PVoFaE/ndkSzqEqB7Dq3b3+7OKJA0zkyB/vr9e0Bx
tE6AKclfc18iaSbsyWbQvLrYescMwUw4t5qePcT3IdPKfLe4ViGOw0YS+uW7QmC7
0sjly1oNYyfEqHtgIMqP8Q==
`protect END_PROTECTED
