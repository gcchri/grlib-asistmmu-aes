`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8F5vAHeCPYYchlj+1jtQeQO37tZvuLsmyOedF7qDdnUNOaZNWYpegtxjTB/Bt8ba
BOcXzl31ZQEr79VJ7fujn991yjbKa5HkmNxyt6B/RtePVpvVgO+owxxh3nS9T1/w
Kjnn4GzAjnSqbsYiU0IRYvtLwFksuJ9pGGBl1oCgbaSwTuiSsD6UUP8S/63bTo1g
pscAJ3KCjUfSSusz0sAUQ0AiwyZAzWJvamLH27nLC9g8z/5LwRD5uGKLT66JzKSq
xTSR6MoPxKvcrizCmZH/IxPhD+b2IlkhGgMMvZjEbmt2DXpX+ef5EQJ3Jm0L3/FV
orG+50IRot+LFnRFL7sIN26Ya5aTZyeyIGq8xOwgb1Mljc0H1ywKCNOTp8u2G9bI
/W7+Oi3CXxuN2+Cg08BMMowHwlzJFfTkCw8TbdZGTVEoSRsnGPSS81qnmfBb+lA0
AL8wzIlqlfMGY1plGjpyF2Lx+lsavV8He8LzUP7NCxtBRYHNZX/yycCBPzmWU52v
k40ciHBXt+fNBP5VnKYJ/3CuUL4+D4ZW8NpapvZn7ikTpI6gYLVAaOtlD8Z0ORYO
gd8hehvbdJjF6c/6GU85CXY3WKoMI797j3fqh/ZyLdDaaWd9dJpeDIyZvv7K78EX
NSYeSGnaYURFScvnyexDny2P7tF9uKSiEjF2HWZLPrng9fKe3kpMm11GhmN3f4C5
79R8RF1TTfGw0TdydG9abF7AO2iLKv9kKI5yO3VheenSWZ5GilaEDp48hl5a8U5+
QLTjTC4nvaEfiwzk7I+kAdWhNhDLN9cLxEhJ5aAasMqi1MRx3aoXkrkniglNRRIO
AogoOs/trDY0VWQaftRhD2tJTQKPzOP5Q1/iqEo0i0h9dm3fkduSogsLsNh3W0Ae
6ICupe15jBhTQjtdWnnaXKzMzZaJvyLDBGXIanFmAmEj/IwfqqGlu/rkBgG74IN7
Fi/YOJqhsWt/FkxKRTLkESfCPTkPdgt9/8IutElbZIVWZPGjH3j6RvPgFxu51bzX
`protect END_PROTECTED
