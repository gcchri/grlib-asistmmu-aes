`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/n3GdNQzMCDFshLrAt1ywnFhuRtrKcI6LRPrSExRJhwaZCX+26WFvpRt+6pAexK
T7DUkz+LM5iRsntbvZEnKqH5w69qk5kcr+a7WnwkjBNbjC8MQfSgT+g8x8DuWQsp
zhZQUHT1cnzUST97eE+SDKV1pTFhFZLxOT9jb56+Tg2JkQ2ufbdXspyGIe3ee/K1
uuaJ/5zzkHQuDtsENrwkPlPEgAxSVSUtw7f2MMpisBvkzo2W+kbjxhrc1pBjk/wI
2eKNEOL5H3jBEnhKIVzz14Qh193E80jZWt1bSZD8trqzXgWbfPlOREiDxWU/Snr1
PVO67aozvFzHr9hZJOntUouIwZOEtKCsp0A3N/NoncPKpw0L2+OXvsrOKF/1qkxC
wz3QGCKzxXA2cRVidcPyHyz2CEzlVrf1ORbVdDX1Tra8f9gkY4IYlmOazSzmrtnr
yJjSbIoQW61cZUpjxTYaTYnFjGfjYzM5GN/hInPl5BBSEwdJlpdk8+h3+8gh8DuQ
2LFDGzaUkFykdSwOe63WW4PQVzTk7XSBpqQzNiPISMvVERiR6DVpIX1e1HvE9JTs
y55z9sLTD4/6DPm+dZ7jLqhaUgZuJ0Y2tUCiIWxX93grHsNS38K9Y2iK6VJuvyTt
B4Hp429Iwh8Hm3/oPDoWeEuij8dKx4GkBDOQVJYfGw2rmLtlpUGuFGqh9EM87fc2
dtCYAXMTLxloSB8e7M9/x1r1EeZTEXwE5dHYhu1roYgCUkjoOVrrgKQKDfm5S1Rq
OUYgFWCjydqHtJum/1kffaAUvGmwHZWiA1LZXVVqSjZqVoc3r5HpwMyUpUAKA1W3
Rsg8pPurb3uesoG1HPj8jysx4VdTXzTYewV/IivTSimi59ZQVbusdD9QMHWO3AOi
vlsW25w/9Bc5aqfN+aESxoNZG3u9lK0xfv0xef3XDyEgH9phJ+RXJYPVjZq64pKz
xpP3P8ocVjP59EQqoQpNUQ8CYImeqJuR8TcfFJzPaMftS4FFxE/GQeYe+q4wJ4Dp
Pp3T/vI1l91WbqarMxsw0WGJ5cOn9bsuyIm83qKFpuaktO+yQkRMfuxT/ZB+HXwC
jNCaifzVzkzKp2YlOIKr4ccOTNMaFaVGktL0fR2XTK0Xz6rZ/J4tk7aPjXxCBwC+
WLsSMxx4bnpyPfcllHj9UhE9wjcF7NkcATQdjJsWIWyX3vfctG6dvUziXUSKe5tD
mjclo5dQpL1aIEK8oJHqYILtWPnywZ/jI9pi37vNb2cTrufbjLNU9ACiYfYKgM+S
sMclKy6sCI9v3no63e1F3ysjMmuhoCfzr+61xoiUXh7joHhlwraCKxKlMc5i2UdB
zL0gS9DzIIdlYIhbDvLoK+ilLYxZLtMIQ+OTiw/lzISWTnrhqnbfkPBR2dskvXBE
Q9HUKBo3iIya+ZTQThBR6smNBgmmgMI1g3h2XQtB6SzvzcBhgoz4UtGxP2t6V3Gh
qT/hyE2qbDmxYvF5HlbQb+O5DijZWY4qrr+I6UsH1BeqKa3aCNJYISAaVEMXO1Zw
x1Z2R9cEk7cyd305Ioh0TYlAS1xpB2oAomnX3/XrUZVKnVSfLMnpQUL/krR+MY8u
6CvPFPsBazWXZSQVJlmZ1+CvBxNNjy7AmZtaHviuqdbS74Cjk6/IojkOZF1OqbAl
DQsTTWQQgJIiC1iF1hQPBFG/f21jEveA7d4hL3YgIq/qCD9z0B8F+DukSOD70NMm
MQdwyRztdaWAtCFlpKScFonSgJHfbIdCrdznejEpbXzhIk0sm1Z8KgjpjoNx5LB4
+BL/IOq65SusN3ADUFPL1lucJS/6gxkcGQDtSWuRLWYTEhu5DjoiC+lrhoOM0zxX
JBO86sC0vKFwmIEcSe/JirY8Llb5Mqd51itQ0cg7JPnLiKYdVBZohENzNXqbUjQy
22A/A2Xc7XCkYBtUd9Pcd0IuXCJF3ouTKpH5atLiro8WGXGIC4s9NF36vWQ8U2oB
9uJxwsdUYVL0tMQY9b9xVq+oLRX5ml6cHvg3PA7+1wtpEDHcicPPg9CoxKRnshw5
ETyaoTdfe0tYe23DrLd0din4wxgwOvqsGeNAONfhSb4jgj8i+3u1sxV5KiXIHQE0
V19aV+ykkQU/jRNMhSlUFNO1jbdZLAvC5ArHSEAaxBjPH4+IZFzb7ab+t5pSVDts
KwvXPJfeq88m8CzLZcQEwvXKwOWU+NrZH4K52kYbkp5/JEJ25LRJw+rAY4YxHFVs
eLkbaJSdx6xiG3FBI4mM/Zw6VO//bneKmxmViorQis9WJUaYl0iET+XxTNFZX+6Y
KcCxk/b1E1BGxkcYcngGIE2EUpjtAU+xgjMcMKJZbDNYEPe0u5QcRNhpc4faLHNC
bjns2IE/6NRr0Fx8vNCiwtDb91EnDCB2rfWhS4XoGbRX/9ahKuZQjWdsaMzUFriO
EmYdfSGRMGsYumQwqYiM3HxP8etcAJBVagcQfMRa5nLRLpS4VcBBosgS/jRhbS7b
O0kV1ZxGjUOzwOmqfFfe7ooaozSu5e9xC2usw7qjuC5Fe0VNOA9bKF1Yqix9kXni
wt2+EfhXvELZzfR6WZbtnonixwI0ORVk4ZzjoZ0VCwawFLdHZ+l5a7oDf88o1l6d
2qKTq5z/3zTXx+ZYhGU34HUMzGmnHshDYEKyMressx3h5Sk+Qic80oxO+5emodsX
/hOZjtOGl7OSD7gVSXCxCGAVRI7+QoEi2c5v7bEAWoQSOpvk07BjIcxZDoH/zfIA
GG/nGUleEpOF88WSdv5UN9X5kl4cLSPd5c05tgVUP987PITFBY+ttpXcSqv5DQUi
LjFTxJfh+Mt/4I+Qja+459kF3zLp5QvDp4C+yyaNCaoZmm2sD2XDr9GUS1yyQs8n
BSK6UxATbDGoH1PyocWcACEc2rc6NqIRauHDgI0Bb6abD8MH/+F0++N5RXK83/+O
VCkgSxDMXXqyLnzykntRTvt7SQgKdHhHX2T/5d8iNJByvrHu7QucTGdGddm2ADGy
Uq0cUXt0yqQAI9Pzyh+0eyGIpl26K+dgUF1GwuIdXQvrw7HuVwj7spGHAyVdNeNi
W+nE4o6CsefHzJHYx8mBPMWZSLAJnXW9YS6gg47LbtHsDRvfzg9APSuQON/x8u+h
LN8V6HxHjxr4apeuOBSX5+FoWQVZFFfCARj3oW7Cy42geFt2rThc+ouGFXhuu/z/
dD7zv8mam9+6ffHVsqGfY60JH/yv9VEwEqTbyiNDxWqCIvv29P949HMR26Z+ZKKf
L068vvyJuFrb9fB56ynXl8MVlnRYwZMZdsXv4ra7Bf2wof7Rrmhq431bQCOb9i5W
o6kK6AUwDk3UmFn5cBBbpCvgneKvVexRl9QY4+T22kiuDzAGIIR80TspuaShzKD9
8MoNgsHBi/Ry07vGAVJk33XyOiiHctpnHyrO/iFTeLwAqEJGtht0jAbFNL3jlzeL
/05Q8BOKI+2IqjeA598HA9a6cht++r1Z7PuSpAxfRjBgnCX2l23BwNhqgjNbujSU
S8Lu6K1+s0gHeE4eAMy1O7P+WmODX+NNJHNLblZEhmZIyhJ//BQPh83EypFqdfUb
WP6Dh7HKuO1j5mFD1QRPY6hulSXOAKLQH6xppwozvONaselz7SD1udliiUvc3eya
jHLcRxJ2zJPGL1yFKHngKhW4zydQr9GdeLoVwLeLn49uaupv6DDSm9aVlTurnhq1
1YnxJsahaR1zuA6aB2hyWSDFrLa1nwoJalW/6brM6LlNN7pQtrzyFa3fBNhs4Jmo
cHDyBhL47NzMkkidUV0zgCIWoL0WRZOZcAqVoKDKdZmPYD1NtDYkhlTeBF97KepS
nC1gVmAJxwoXgW9lXU2wtsOSRJ1kDFvJGURZ5mgemxMDiNnGbYXfFA9VEDQIzdlm
qCrpjEB/nrJODQ1UZ6cO4OwVGUEMSWC3XZOojL7b9cYvRqh0b194mMpS5lvlp+Zk
XyvQ2EBWiUxWlGiE7UufjVwV3f5kpK1GI9S2bnYBzUKV0DOGKzR9V5nDtmZfSbKz
mrHF/JzTeYp0jTBUB837vkRCYKahQlues4QVHZUFZo/FmXUUzNqOKfznnmkhZFhm
ob8Sy8rtMiJwQ1JYDS+uItHY4G4z/clix2d7DTkFxYlK6o+lofPjKyUsaIxxyScn
UhpFbNsdglOVyPACLgZ2q4wyEmltvKZWjgDXt0M4/deTHD/WU8P/pX4s0Sp1gWDX
VAdjxHfCpHYz9YXeZoo0EkgoeoyzFLjuvcssHt9gIWyuXRC1TRwfP6kolpieqC25
2UT7/aE613LwMWUjqRL3sirM4zirM3rfxU9u3mGwF9LeIl+kPfEI04s9EEOuuTTw
YbcEzgQaXFkMXMfkQZHi02UTdnKrKmAFCmlMobZ6DtRHk7RPNsaQWu86i2HxBRKJ
d2eLNaj4rjnmvMrikh2/Ys0aFAmRMWcl4VUPuGMnlTi5uiguyJk4uxeM24j9tNQZ
PFpj5F1P/5o70KkwWe7iKCzPXvuZxJ/yp/jcfej5lwzwU6sG3Yoy3nWPFu73Fs3c
+lEQZ1AIUZdWxHmnf86UQvPWpEabH7Kd7ZHgU4CixRW3l8D4vdg6n7iID6Fpsijj
f/rD0/wFNZzHpUGwVJa3FTuMzX6u9uhqjan0kYoHVEleWdN03Ro0Rg/CLBC/g6GA
kplc02ttJkppV/0j1XmOKUDGdKrWIuHBcV/FXjfdPJc=
`protect END_PROTECTED
