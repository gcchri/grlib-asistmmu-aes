`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5leMRhInVEraGidT70sn1r1tkNRCOAvLFFgNz54XmeklBmdHbRucQLCMCugHp7eF
2dvY6y25hla7BCjxEwoyB/8Xla7nUDYvjDzvbzgABdvlsrp963/eeEJtCtByEuqZ
b+54ua3Vg0LxI/LEV0e9Afm9a4hmmBf91Jw5DkTINYE+9u2ijjafQNw3GKuJhbL0
s2EWDpng0T1CAmqdGg8enbl6wv5gP/PYD4fOjosLMIzxgHWXN2UlNMz+0ME63gL2
6tllJHh2Bc26IqouBhbp/Q9WBjZK63pf0n9DgTmZLc0=
`protect END_PROTECTED
