`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tKAdXm+7WJ5VG1iUAYES2EYGEie5gLuwq2PKGFNr4hwhr0kWpz/Wn1ZiGfp1F7r+
pnwZl7x3kaFmJQcqeiVOV6bS4N+jYZqJ74NidKwYVTXSD/G6ibFE2mpKKyw4aH6F
dvkzAHJVu9R6Zrh5ZaqNKyWuM1OOuhc0gKHt3IRqVSpxPyZ8TlXJhm51t2EQwUew
AzOSFZ0uYOuEgN8xS20Zj2J5pKnFsb2T2gz0yxK2Fg2a+T/VcQxuIm1tuGDwZEBU
lQ3yVqxdLwZpkncebBlUff2f64w4EI6cUQyLM3xhsTZzLg1vxnp05goKgD2pjYYZ
3PpoLSkVYfiUkFVhtB8ErmvJ8f93cEda075gm3k4/JBweH6eVjSEa4qESpErVusq
UWG2xqClJRQFZ44f0beJzmtI/zcAN59O5GRfR5zqOFORaBTzj4kvhWDVeCxQ/yr9
7MCs6QRHj3GbPT2uWCt8C4E4jrguhCCz3gY6oTcdqCjq6JGmAGXR1HYzzDcP92wm
`protect END_PROTECTED
