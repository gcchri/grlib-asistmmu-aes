`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3oHcymPt3G8TCQdPyADsPVID31JlgD76vj592t9awZMtEpbj4qk16pReALs5QClo
WXIVIGVAfTZnAGrOy+0pCO0CBKxf9XZI2IFWlCfYBlnNfdx/CSHjzMc4mnxjJj7m
jPpyh+sEfS8UumDp5l4urHAB/S0EF764akkoc4az5oAbPRNobZlDkdPBbn1XWNyD
9BpEhFjetV4oJb9Wt07FCa7yqwpNKM6rq20i3HRvb2D+8M+KjME4u1Rbzq4wQaw9
g6IJ2FNCTF9nsYAQWhvB+VkSJIzHXNigfjGW9e39ccqH4fN8MQBG1KsfNkJ05z10
t/+cTFx6yIlYEB6HfMD3FTdtNigCvDkaPFK0Riujjhgv5a9BTZTDUetSpOy6DUn7
lJDDqSQso2yf8/R54vObkp/Uf/++iWhHO3qhdmzN0sc=
`protect END_PROTECTED
