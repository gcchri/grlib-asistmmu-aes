`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zprhyjt/9iSHk9psbc7PxKPFNlSvmiyULZqf2G3e58FI3KC8n8vr9m6WQXvrkVzo
7QUgjiMiTcEfTzatCiqMp/rAQyIiRhFARrICMJViagoTIxV/py+hCmygO/8SoeNW
yas+SWh9KbTKqsGS5MylJ4J2VlBQnjcVLFSAj66CuZsIj87LyNIZKINsncYAVhNT
FYehBfL9cvuF1jrbr3IgE6byjYH6yFXzjFs7+xMp+Yy4isFAMAl+n/KWAn6xCujS
/blSN/Eur6LdMctYshIH6ieAN6PByMp1VfiVeTEEpN7kmcghedrGX3RT6aD/R2Wj
4DGTxOQnrkBEfKB5LIDOLA==
`protect END_PROTECTED
