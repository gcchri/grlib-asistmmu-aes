`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGNo6as8XTB+XGb2gpNb+5T9j8uzCfTdBvuSgsUwmmNHf6tQmz3lCYH0Z93pXA1O
2OnpVDs+YuD3QtIBPGNmGsOyExsm3VvW3GCHmvKQjJbhpOAOGqxBs4ia8leVJnYZ
0WASrrUniJBUMdEMxJIa/KXeH6PAlrjJfFgNKqzbYjM/IB7lcNbkuH32fyHERJYx
+aGAl+Ji42tRS9DoUkcQDTelZDCU33R/X8B4XCuKLTktl5ec9abopLkYeF2UO6zU
QMxeVjgI4esUQLEXuHHYmqbMFE2JeOZkC5w8rkaMYSD/QC1u/4kVqyueEAvisZM7
P26kq5XKTe518a90gdudcOR6TckVdjaHmLwCsR1Ut3orHILL3GiqgH7mSMEqe7Dj
0aUVJShTBR2TPj34e4Nc9YJXTwmH86e5KqFKZT9ARrNCCkAyJbrKD8ONYbtug/hE
AS68blL3tAnGu2yLNnFhIODm97eZqxfZgsnrn7ES7LX0PQxeoQhWqTT7T0wTwt8F
`protect END_PROTECTED
