`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YuAQM/ehiKGgSdypyLYastMY4y1EI5bUwsqcm/Zg8HOpjcctQ+LTya9RocHNLa0A
ZsQXbPGTgyH17xkjHPLtbdlGNwRJaSX3YHED6DO0AiNw+xGVJf0XPOt74U7eINx+
Gsa3VAsxMRDXrEPxN/FU+eAUQxS1HlxA4F17/t39GxkcqRQq5Xz+jKsW7d//hWSR
LMff3GDp7AHML4+h6tObXe+ZcbNZK/MavOq/J3PrJedr5YkHAOv2xZeTWVgkzV34
KB1eh9ju8ntD/SmsQ7QWek2AipIc86tYBNe8KnNzAXKiVSeqtFKu0plZMk6lmrwB
qLJiElSQf/9GVURdEJBXkfoNDHF44mgmpmn7oIY8i2TYataRKF0xIxApv5Y+3aEW
`protect END_PROTECTED
