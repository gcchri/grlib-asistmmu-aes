`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uj2HuFYgljvMNt8TtMj+bdDfmfY1sRABm1o78/eVYd81LTPTknjrQLIp/4BeTKBN
Blrgr2q7HQgmn1z5xaMXT+E7CZK+NSjaJwUhL1UQr3jKikVOQq24Sblkn0PZtY8t
GXMjeayyJPrnkAOUgOc6s/xH12FoueUHw01gOcbYMmCaO1R1lUg+aqqlqRR3HVQW
QgxWbXsqYVjNM2aFsC+gkYGllCUGrKN2bagNTi/LGHIP1VqpLhSTw919XEVf6Wvj
s/3OOmCOuoArY3iDikeoNWu+ENQxNUfOiIkj0kYp4V3LrzD4Jmr5CoROVDkpwgk8
vnyTm9y0PYkipRIW2/2hWn+Vwb3ufWR8NUaCX0f/AM5rT+t6ePpWtsd9N8EnSYXc
giKhdslk0kAJxx/CTVcleJpVeTpruHl/GTj71Pjq8UAq3pEl7PzctIddwq4V6NN0
E8cf++pzPEvwHi0e4M+kx+FV8gOfRzR7Zj12XZWO8dsW2hzDcaGUc+eTtqGrdol0
Th+GodD1jR4c0hKNJZLd7070qgH4sWPFhYJEE0AG03QwRHSBU8uqyAq+1fxyCgnh
30Ab3R4Rl0fYhIe/j3Rj132O7xuvftJP/RVBsucRk7irEuRBERNHj/qc/y4RrvM6
6sRbOpQk/d9Hngj7+8Nund99smdFX+KadjXYUcAuLOr6gjKVQFBpsAr1LeleGDzN
iEMVPSiU1iEnc3F3Psddt2/CEAe+h5LKUEVad0tCM3RZQRLMBSAOgnhNZmmdjB7i
tniKkeOV2sNaKktT0Y7D3f5JjGwIbcCbhB8STlkWMA349rBYQWVZAOvInugHxxwj
36aDhVSGVFgH77AmyL7oJSayhgb+V4Dt27LENpuqUwDYL3HZpNWmMvzfmQRS6O+E
7YybxLkwSZPOMT2tY99NPA==
`protect END_PROTECTED
