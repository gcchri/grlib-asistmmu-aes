`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBuGBXRAQqqSltIshVF8fpqFudDG0nh2VIS9D07U1gKhfhO5m5W+CRSfdOoEO+dW
ykg9gmJTmpzMKhkG8hLrvEfwr1MMdiBmt92M8rgts22okXMKiMUQuVf/fHgTyAQ2
6iKiv69IZLHBSICi6BZwsaRzTZdCBTIApXSA/gUYMijRTmTSpAn3dtYO1Cnka5rD
85PNjcyjDX9qUWyA6HaotV5OOcGudcacEIVvAk0Gy26FXbFUJIlkrgjJAJdeFXbO
ua0MkeFjxeaTXdZqmANPaXpPUwJfVrVKRJ/kN9gHkMVEHfM+IsLuQxr6Veuzoc0Y
HTgD5UqU4YTf6cj1nMTeH3dXHoAO9klLFXxmYDBpCE47h4bo/vQNx+upfmkmP6we
yP9GKS34wsuo1gcZ4zj4ySJn0erej9Un3ua5dNKkswOyk7TjJGKiSHTEQ2479YU9
pOjUoc0+zjkszAWAeb6bgA==
`protect END_PROTECTED
