`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
miaJJB+uvg0H0WmcWG8iQkZq0kcFMcewnQ1RSiForHkJ06ypuPfwJVztgLuyXGRL
Mwi/nrdClF0s2jDjROCLI/1Vcl83ju8hnEage5RsbmRX4M087cUhTpGJXNcl0Sqh
BhEYRy3dtwrEL5FOycMkya+yogrPUIDRzWsBLmcYKAbLZEeTM/6H+vuHAHu8XWau
OU3T3AKpS/Z2icN/L9UHEfCuUMPifLlsMu0/0VcDhTARCeN2zRxJF+SIoUO9xMkG
zxyptRDcwWFhWZuneaflFpUy1kf9DmrKGl3y8SNgKr0=
`protect END_PROTECTED
