`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OC2cP9+lK9iGrgQCkxIFM0IDf3+eSo4KcjhE+KfaBscp4s03g05iGdhX2TTXYFtr
TRqi7YryxkGc2mucF98MeWdXKEjj7M7oYG3TmG/hNPvrhS8FMAmVmHQleISTFvQF
9Fln6Z7ICZW8lbnieIkWvX0H6WLLL0k+Wi4Vu40bzdnSGqfjpZgZO6vY0wjBAi4f
HSCKLCt0giV8DZgYVEoXU+W/5Y98dxlsnRE1LNDlsZw6sugB3zoeIEjYFIxoy8HA
`protect END_PROTECTED
