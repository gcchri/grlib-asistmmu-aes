`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BaDShFDQXv/gjwzg2bHDkHiSVyhrSvYy2N0EihXnJS+5o6pe8xwlJCmWjyCzkrfj
dc/+ggMdlCOv4i6opwrle+V0qK0p2sG6ifJWzjuABaXw1te6T5MvcySXmu2XmAtj
dyxo5qIlKIYmhdNo25RcJ6AYgockAh6nEjGb1rtGCKQo6F7VzZCz9QTJpNa6xkgn
YihsxUics0//5wDInhkLRFt0tKfbCXmxlZlAYzvuIayvp+61g/aTFF1prj4VH5Il
UkT8uoD5FbLF1rc/Fool8KwrjNCj1WqGEwxsJrwsWaH7vrANBwfITnZMuZsipdX/
qO96H9gB6BtYwWi2LCIWdw==
`protect END_PROTECTED
