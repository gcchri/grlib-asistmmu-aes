`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FxvYFEObKmzgRUrff6REPEtDRUpOR9ox7KVNXAQFrghIlA1V+3Atc/RTFJG6eOUA
T9Kk7TwGEilj5hCyNAMUxRju5pvpe0EpMarxPcgkQTQ10J9uxyuSukGjmCmFquvW
jrMQOt5l6YvMiTp2cvLtbIj2B2SVljOlbLGAOxXOBS+NyQgtbaJPlLhM+gRz1ErM
/xPvlYNAWQnXRtHj7l0JmM3OEevxHO2BroEY9pr7gdXQG93L8L7cgtspQ0IAY9di
wnEpu0qtOH3HTQATY4MHlwk+NF2MjHV3LN4cmfU0C/45wnrPJL3MQmGYq1LpKJAs
58hYNtD6xAQU+d/j9f2VyPhwgSSz1XU/0iDHQaauBshgNOx91S3MxVmN3A0MwgAg
UBgXpBJErRTrY4IhQR6HlMD0KUCdiS8yt7iIIM1e76k=
`protect END_PROTECTED
