`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmPo+CHmrpWSX1N+K/vvMOk7CllfRg93DmjOWLacRH9hXg8JoHe+ciKrDibnRUZ4
Eotp/67MU/TcWgmmf06Q+kIpqG4hq6UFwjP+/TYcZbzu66q1/GPf54z++F30So63
hcl7zg538ubw7u1/JNsq/4u5qknUiIcUj/p8aXkSmtsxq9VyRmCkEJugRA28C1/4
xSGUeDnhF0+KOXPFK/N4RypiUT48okRT1YH6+qOzGUdB7xiSxj8YoOr8hNHP7MjQ
F8TCTFth4HCu8FD2AauDdb+STLV0WUBx4zvmvAUEpjLs2pExyctLDB75UqOU/ONS
ai7aBWehQASr5a0vH1aljg==
`protect END_PROTECTED
