`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y7FPLvqlu4N7R+zNp2AmQ0/dvPVZmo8qGNRS9m0CtMCqFG5Ki1ND5TBWH5xjJtMF
EKSbJDvXpP5TP5gQw3EK+DhHDgG7PTptMHC8rrLB1+TSdaKy+TjD291VbpqvFmGc
c5GtTzjdHCONIw5+p9ZGzHUeXGzVmdJK2ReoOavDf00UM7Iy7y7MHcUcKvkAQDRJ
GVC92uX65zQOma7z2kc5V8Sx5tlejC7S2H689R6XDTFTjrG2V4KORQZP8KLY9joo
qW/SgipunYij//YhtahnXWsiRjAG03g+VKDUVjoblLoYhqvkWw1BiuWnqa/QE8I+
Q1hGAK1KiF3ApEetCKFO4DWd1+32jMciYbCxmmY33yAhSz8To7iJ/+kJESdMaYGB
hz7PD9s7iJmidyOJA1ul0BXlIH0Ys3lE0wBs64IPoqvS1Tlja1oXA3n/DTJn82aL
/xT6X7xXC9PyeBwkYaiiKKbWO/fvwJSuudOgmKTpkES9hFkvCOhyD8SWQVINRIRM
xVY2671w4E+EzvQ2snj3+/NrScx8WmiWmZDgaPsEcquZHZFxOGMPWADqutk63Oe/
Srk8U42NUJQC0qZyJJfnB6WhiJw+WiFGUu9CknbQ1onops5NBLE/hYpcJdp3pxeK
mDyq924b4+HnPil6/vvsaldQ8HQOigYG3o51Hu43+4q7VYB26iJIRaHy9rr17H9l
JdhFwJA/Mw+3CE+xk8CDgEaH0y3LBMnn6gCp57GMLtknh/UWMU+Um48ScDAwlT3C
uB0WEWoUHlHCxdcULRfwsxsOOAc3TobZmHkbbGDcqlHR7/h6i1gEIfPIOVSfsNw0
4y1Zv6fOb50i9GWgtF3wCbvHTpV0Nwmgu6kuQnXu/CHDROMnjjtYhbN+xQl+8wf+
/3Oi8dnjrqRNU9lp9kKQSejXgpPu+HhUp6o4H7uZL/9Nq3zrluGh9eEIRKugr2gd
+uZ0LrqXaZxoxWcI28Np3j2k0dLQzgdn0Qod8xMZhkPyJB20N3ISNGV8EHGZ9ZSG
gF9yia7Zrilq7HvFxvol4QcZuW9DxeOCvKOyWd/sJjLUplvrx4Uq1fF9YM0ilM+L
TMl4tXWvdZbAhlqh2APOqqb/aPXFzpUdNODUnc8VGfZTIeLqjirgXRQa7MfnDZH9
LlD74VrycSXPqkAd972SY7FVbRIF3FmSekgdDMX1/jzK/67Qnjn+bG/GQz2iUJfh
0l1tGlLye/mjnKAOMoP6vnLIWyTbLgcI3dKPjqQcv+qYnkFG1ZNRVEP/qUFSOUK1
`protect END_PROTECTED
