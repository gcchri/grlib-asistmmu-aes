`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBQt1k3uJSMZ6yXmVuZVbqDnpwKgHAmWSwknPSuI8BuYyH0wAkV8tyTRQeBVlEki
uFqSCSBrrCnotXGFIofbWucMNe7f5vyBT0zR0quvcHYikhXLWy/ldGLULiTHsECh
W/WW9UTFQfKnEwJl5S0E5cKPJpSh+J6FF304F3eVdW1+pzWqBT58hRbD/Pzg65b2
zvRdR5SMrmIkYWc0BxqXQJQtyCm594ZNQN2VTgfuahY=
`protect END_PROTECTED
