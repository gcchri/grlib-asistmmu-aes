`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBTHKWTGt8pWu+VaO5FbdUDDpeS0Wgeo1NZz4qDF59vhI1BGr4pVjXEgcH8g+WOI
8emvOYGPp1EwfAtTXViQnh/Hk8woHdfR9lLGrF+txOI9w0qSuSWVOF4y7b03xC4K
XVNwYnX+r4T3iu5Nn7eVK/bxGSTVeqw5zB32fcvTOIhlekPiUXRIZLxranJh+Mcx
lA8zuY3XtBoNo5UOXeXQ0dK4edIEcqW4Lg5XaXPEOxayKo8e5pl3No5JrwsyJnf3
bAInpt+zzEu65UIRtONXO5reGe6LyTLbKjgR4+F1TJTN7tzyA+XN1bvxVjD4bGHJ
sWu3FyxjWySG6eChrybgn9D99rVkdC+Mvoyvn75+vUQfiFKVkM8m9N8BGnqw48rO
0E4/2YoGoaLvtP00RWNB1yqUXpe49Qd2COmjk2psIBcjDelj8TGcLfie48yDP/Q5
2EnPnGjakZc+DQqmonPL3rXMm0iORhKLB4mVmxvKiHWq6FYZ4TF6UJJ1Ja8r1FqK
NTX2VaHrkJD+TUeQgf2HKbMT6jOz3lqz/gTU93+PT0v/+H3V0Jg/F1QfaFUWBENC
AVq5KS1vfX+aJBYYUtC9hlNqGVoeAP/5aqe40Oc75YCrun9Rbo+ldqTwUv30QTzz
Vs9DaEpNJPlStWOdm15zEdJbMaogPxSTdimNBKtw/J83Hf3gsqJxEa4z365QgHee
/JZyOvH+fuudaxdJpawlECEV2T1n30HAOOKZg/j4si8rVm53dpox9AJuI3jFydA+
C8TdCtiEL4b9IVT85OFejH7NihF0hECBmMi0QZiPGaKC79pcfL1KUnUAileI4L+0
fnuUEiT6cuuLFLpz1LLTrjyfd1hWKTWYlacrkLmAY21clRpVD0vPg8WC9QJKiScH
TMKzTE1tj+KsrK7BAHLgLZtAv+pFhmj5gyQyYTOPhMyR7sjVJzvWYF+u9APO64Pm
ttQ9cNv3gpmaEjQiZbp1y5nRLRUXcqw9EWjGB+FUtNkF91WUDev9kn5ZLf1VVHNR
gNHG3dUnEwMcPKA69OjXLKLoLD58XtGwiqChBscNhgGgVbwtPWxGVWO/G+v1/pSd
V3S5HBv98LXineajv3Ype5xYql0DO4GbWPBzd3jURlwkYKDsCuqngnjL5SIefrnR
YPVUtMN/sQPvmvIFTkkSQvqc8nMe8qXg3TTYve7KT/o8fgjDVnPCR1iLumUJphVw
ZEf8WXiwi5Q+38MPCdQmpw4PCAEkfwas2+dbKcfPGNslmFDtWOERGUMwUTkF7A2r
QMDUONVcYlo6caBofT53CN9oCHjqWoE5E0GfK9QYvv0x/Pis7t3eSL7QOePAJNrL
Icu+1dJIvv3HKWapZaBgt2kEp6fdZC6rwnjkZobMhtH/fJmLzw6xDUFG1IyYCheF
DWBiNQffr47EevZiWfIjqfjPiEzpo9cZxzgjsi0Xjv8kUzijCJPUjdgVHBvB39D+
Y1WJ1ej0NjxEtQr3Ca8PHpizuF36gdxn1RD6LsDG/mLbbFQ1u8FdAvFXaOc0DJDw
cb6LP0TtB1ZdZohit422XfRG95XqXs1dm9Vm2OjU/WrONUrDulH2bBlgE1xZzsbA
8dHpEjyxOXmXbKaC30lAJ3wjlFgRgyF7e9ztHUSwbKzk/gmEq7NS3txktQ4Hmguz
fTervPrLN/AFWqUYiVQa5M8Ue6YWxn5Ij6t/l2ulANMrZh7HKCHM5o9WHuMXdFBH
te5C6fA8kevDnslBJgCct9UMiDq3tjV+e3F+cu+UFRITx78MYl3M8xNVS1EJypJG
dVkK9/NekXyv6j1jd8gH6xX1Az8RnmoHROI0+xAwjPJz0hH9EwzmFalzZDKpW0xV
Jqt8Oa6uMA/2kjaPZF7OkCL7dxaNidyVz0h+FKjExwleodi5osWlOJYuz/wYq8+h
epqIoHg/nO/PDEkey9OIzeD5foPyZlp+9qzLPfk4lxVfLxNv3JAdaDv/xk1glZyM
KTdQgHImiDkxe1q7lVxQWtm+HswwnTMlFK4ICiTYaQvUVDtJ110QgN49JcyvxanO
tmDjH2bTnfGIW7jBmST9021ufFWOwYk3GUjwmHyUQ1S07+ubA0odILYQ0PTNb17s
Zg2sANMx3YEuPgJ6+t7Z+4HK3evVJps3eCeh/K5tVAwSkDXVly62BsK5uMDNDwR2
NH2r8UvidS0q0czh3KQ6mx63k7LRzoyk8I1Sd9XRql6bVi2fCNGp/xLo79okjnnb
um6zKeaU467qen3ibEHLDHqPJTMZqLj0wFV+F27s1RAjAOK1VXkXkU8+0K7cN/F8
w/AVxV8AtzKcGFauTtDDyXqJscLbHAoERNiL0LoY+/TY0mT/gzKd4rjQ7E0GtB4q
rASZd+t15COD8VOEgNDDWhBQcnpHRFIc9D6GfDxgSHZWFX7i6Ja1+osGi+DGA/Wm
1VSpGiwTJR0mJ153+OzB5YWgo3my8LQWl1Y76mBM8gwF0BRi0qkcnSask9Rrmanm
brPymYF9RsuURWtvhtYFMh6bDfJC7agUCdnFCDp8bcI/IuMr/hkY15SqS0lISZGi
3kikKZ51X8JpqDvcpiFjv9bD4MZCEU4K6MkHb+qHtt4AWIUn2D5W3FKqXreU4JV6
GE6zqVDV5kkkU0P+a7pGxIE5ZCCiWAkf7XNUFgNMn8BDA5wuqq4Owa8mfvT5508I
dKJipyAOaui/GqfadrPdjBFELbk4W9LL6VilT9ZVQuwHXqZwXiwK2MGlGAnegoYX
0goE7R+OfbUSb8+NxpRsVXC1RATF3Bx82LzFq/7POR6SdXtKPeXpJLFXWPmy6Uf2
TKa/ZQwowZqyJjThQJF8oJWwiIlyka/yJ0uwuF+XHgMtztrdAd/869xJmnh2hlow
UYJ3RIq1CNhhiOMqAtUbujw9gpI327r0HmwXel7DL7jbZQ41ewCcqTvs/ZnOrEpZ
wzCDVx7j7Gy8LMrtjqk8/ckbTni+CrC2JOlZ3Qa16kWHLCBVRRtqIM2nk8oUOefU
6qC0QyvEMBYDhZSDYkGd/KkkTqwMwqbleFwAen9Hcq0mH4k41NlIFCQnxM+IgSsf
SvL/nqrd0bL1Lj+xcEKtiJF5w8bhnpGTdNT0wfmDIYRb/p1ER91X7v0wazyCz9Zg
rA7ByISSXTAm7DTsR4DFaUGocvqWfWh3nyiHmg3nFghokLc/hKEqmdb6RbTbIkKc
UmpAVxJvQ+IuXqjR78/jD7vgZHuVnkya6wLvZt4Vmjph98d+dJrE3GxH48xD5q2P
cgA4uK7AFVRFiY9OONGpXofY1nz68qyrpbYk4k6YAL4yC8C0gxsN/VzM+h/1L7OK
bvg0s6DiCST0mOX4Xqr5Qzrz3MccwgmYGfH4EEiPNfMBBDFIWtWaMjZkvk9ZQkQW
gIO8wTBDwC21TSQWmXvrbaBIrxhndME9aZZo0Pi6VrS0+pEl0Joe5oxT8GpWHFVl
K7YSN+zE42q+dRLbXdKvbJ+PrtLjsDLGFU1JRDigw/Bv2MlsnApIQSbLYDGMExa5
6Uv4wf8z0+TjZH0/w6kAcxO3r+b1FLaWU9GRQ1CkTiwVh7oh6kzMFo/rtGTXeNIF
LhL5XqqB0NWR3zAhVqCHPtjAuUxObv1rjh+veLOP6y+bkYZ8w3xzbFW/RtmINFvA
kflv//QKZvFoCrJZq/LOuIi9eEbL3FbYbioNmRgYzc3jgulQs9g+HaJRkOmPzlrG
tbaBPoxnSScIuVxLHzdf73lSSpsPERMsiq4pWjMU9vE1Xr9RgcfKNPf/rLEByXQT
Keb9pkpzABFysjYkBz6TqtCZu8lKyGRbaAMWbFGIryR9qKmHjwo9ZDPz1bYx8rPZ
XvQfhpXHWJkR3/i6kyAnji4CiK2BIAsPxqeyKGSGdXN9IXvndZ6ImTz75ZRV7TQS
jg9LIbz5uO1sgAlndEUQBYUHL20Oe3tWj9WHIsC85d1w7i72PlZdsk+uZEqD+9wD
iAhqe6EX24KT+qmAphRjlfvV3F3PY2L3DumdoeXfiENBZNMcErvaJt5Ou+dAxE4m
wp27W/2qfSiTwAXxojNLKNa9ylSnAQA5HFlG1CwWDLxDJloWzE3QRL5vQi38rHpC
7y+t7iwMWyx9RaunVw3ttMlyNnftYzv4MszRxeeM8eUufjKpaWpEvXaDQ/N8FymK
cOVLUpMULnv8kJsJSjJOhyB64WKaYemc8r6a9q+el/YUZXuYUusvB4WFv6FmEAuP
+zal0DpzD6fOqclnLswVGD8Hz2a9pq82XZGJsaMS7xqemU7Jse+MiwvDqpFkMiLl
D3LOjCICM84zy9q0UlN8jQ/IgtOGNORirM8g7kNKrwRQ9TYghYyfuAzieIwsHJEW
Q4bD1KsxdtJwcFBEsWrMkRBuy/xea3Te1PX6Q45C1p4IIgSJzBb2ZWhEefRYEuO7
5nTUAq41CtIRjp412if/Xe69rC2XxVoLs5QDj499JFmDjyHKesofd63IUjnrxiuz
bJkUFJl/ryjYgXwlcko6f0wfzwSCBq5LQjsc0Lgo7molw6kvxPrhgOXOEROjKqzq
P6JfgQGnMpzPiy15fUZama9eJ1P0945awTWUDrXeLq0LJThPnMvvrXxQw7+uAj+4
Cujx8xC8MEfmKbHz2qILKECLEgiebNr4aa+hSAWR0e8Qt+0xFGRadF3OCyfcPo/i
pLbbAEK4CPQ2fEAWLFXnyF303uxAz1QE/Rguy4gr2qLfkET1UZZqsrhfPlmkuND9
5g63Qmsc2lq+B+dSJ0We12VNqWl2NoXD9z8piEIDnNcVHN72bj4EO0jOQZvLTGHO
Xr1ZBlTqwwZmqpmju48+9VvGTaq7Odup52+f7zIRmNol5az0gVlAvDJZX6NaqOKq
VfOh7b5Dwl6is2bNKnCYHN9bNCUVimfJyxxcFDzoiX+QL0JHpd9EkwW7YmTWtr/X
TtYwlJ3qvBaq8us0kk1QiHzCI7/HMN3KC6RuDs3/vOxfM8Twjs6yTgdCcXDQ4+kS
b1m2AbYWIwER6/Xf+GmNwY6smVRZVRJ1CnHwe6PXGZAPyhMiy84yl2o9zIFByQgn
ARfl5KkG4reGhgBNxL3LhCOvR/Hwwkhx0bGECK0EE8YDDmBkP30824Wrz9J5Ptq6
Wx0mOMbEvFsG0PvmJX80qrw48tva9aMl58h/VlcZLOPVpk/iaV+x/w5S6Lug9eSI
bO0k+kERwqLrsrqOMFPXNfvLgZupzilGUDgDdfQRyyaPrTTRuc4Ugu8rFLCiWq9T
oNrRFaT9PU8O1m5X/Y74EUk/H1Dww3vKB/P4DvH6hSAKH4SOSouGSJ8WZEElw+YL
8btule8Y470lLPyJAPOgF9lDnKu54Q5H1h6axMjjVufqX8SMfqKFXSxPlwt+S62t
l5GmOgOJv3Ge9SR12YK1vYBcGS3yJJ0quVECERPJcpFJOSLCBzvqUG5hfH4KrzCc
c+CCRWM1vTQu19bkOwyh4WFMCZVqVRlKISZCu1BLYopXKdAQS6g05o7uArY2/mK8
0A5df+7Yk61LAadq0VX9ddPru5vVCytnq9DGogkSvXezuJnsqC3Zdt6cqK/08Pfa
1YjICupOKoObB56C+wyx41Ofb1Yy/1lP0HtFmbTo1Z9ZjOXoximfZAyrZwEyvMwp
eTqtxPPjkcnKZAUKuIItIUHZVlbXCpapwesUaoCa4QcVwGlDEE6L5cEz2FSCP5wL
Jioby+ovL0y7G4BV2mbeCTwRWYa63j4HyESAaYnE6rMc1PDyrqsh0b05NxotI53E
5QL+B+iG4q/ZFWzKymqKsvufbkmMy1RBSm/1XKjyrxaw7J17FcQ/NSY5NSDboEgW
UBti5gXutBx0+27hsk07lxLkhzlqbeD3awWDICRDwbdzrktCnqHWCLctQ+GEhfJx
59fXu80naK5B4iHkyh3j2pD/LdjS128lALH8J3TZcPmRWU+HX3xxyH6w67FlgiKV
G+XZrlepNyIKvYMaNBVrv2M2ApC3S5mQabKuoA3gQ/klE8iTtre6OpSnaKQ7pU3y
RXbDm4ncsfR5j9ieFlK5mijml8o3tfILNRKTHzFICKSzcE88uPLZ3rHTJVJwkM3i
sdfjwXbhGGaZyKQ9j6uQ35qoSPYoECyaKTeVj+kfjRkvISigNgkTXQ3t/IYqp5Qc
G5mHDMcPlCw0Eeqj+0s8r4P/pXdJNpbuaOwmW75qInlhSBp+Sg3mqRK3zlONhtSL
9x7j6WRsD5pyUcVfSrhdK9tKcfjJEC06njI9FUVfy/fNeDyaWElkDfot/oMmNBhS
0Xt67FIHgkqyUlKqpqeEIMguYwjD3Oa6A8DKYk3WUcLu8yppJ/pPEwl+fzZqoDav
CJAiKq7MgzKyPR6kowoBzC/agVzpe7mFSBjYrpV7iHwZqr13s+PqqM0uhTZex+fY
hAJUd/sDSBnU4HWPDEU3+rypHf+ZHgpP0GFY2yuRJ6Vvjmh9KRvq6r5UiVixNDO9
lGE024FASTjhLsT/od97XtrfvQypPKZPKRXtu5eJ5Am/xC+wPjiSBxrt+bYtL3nz
/22DJIjvDyRI+HYoAiXD8edFxoscToZqVIK6oiPx08uNsdzEvdlgqVw2u2S6+2Zf
DvGkBrhtaMqDMQMty9020SD63gXuPJQmn0I8Nw+Yy6S3K4TdPoucf6ofKv1VXg5E
vuw6kmWDbniMh4+XjfN7zquvrB3VLFbWPGiIfileATPkmfTLYsJ6r4QCOD9QLWGA
CFwcHQKON3YHAF38pNkAH3XDn5k2eDwctlw+x6Mg4GAW6ZKBZR2M5nqzuLtME/IE
oWYZyg+1yeOuPLnfLptY81X1cZN9QfMttAQfALpxVBp9Y+pggncsyD4GPguvylNq
dYUb9QwcNBUz9R9opGThbjT9gou1Ior4wWtjkK6StX/2qGhw3JCxUoaqirf15KSY
aXoWyNZtZ6OtCrkofFbdvRZEUVtEgTnXxHADdjk4qRQcWKYRJyHEIMWyeR4Fbx4C
d3QhDcBUIsKs91pnZgim9TCmQ2jes6mJMD313ihZn0uMF3BVwFmyT+8iFYfHbghN
OfS9neD6a+E+3qUCm/bAlnLFVu5vZJWStXyt+8I4zEdTyAug15Xyef22AHkv8tvu
94cQdR3yulieqVj8bc3L4Go7Abz+0VnBAhRUGCYS/a3KjeijAiLMKdFCxHfHhjOL
EmSyyXiSU5Sy5nMA54sFJj36MkDcbs1m8tBub/F0S5QAWgf6pyRUlyBAO2gPvKF0
8htR2tcZ4SlLZ4G9VWmmnOGLUiWVT0K9XtTtUEFjLW2rgKFIyRsYi9i2O+aHkLXg
IBRVBqvy36fmRBYi60DLOU3nZIuTrRjrJtBDXkMnsXt6zPz1nGmgRzP8SHLQXWWe
ZpId5dKNTu/h2E92OS56Ai8OwnIscPySyvrSfqS9evPURNDsyUj8pMGjnR7svV6/
KYR4JroecJELBIkRRxUhXII0sT1G0lhEqrxuITrsrtBA49Rz/P1IBiwaD6d6ZHsm
xhTtTxZ/2tDDdH0J76tqlisr2xVUy4rlebQk9S5nZ1/ti73Y8tDX6K7uxSZ3GIcF
C3CUC7ty/ikICV/5hMw3vYsDie7Y6eRb0GxNyEpYJ96cZrH6Qw2JNnCPdA6R6B2y
UFoTh4ehhPuL3rHaVraCWtB5yYC0MVpLIbxF1BQTHDklpSkL+drwbOXQ9FGYb56x
8+T7xDQWtqxzW4Mx9g3TznP15LhKKV9bDEqt/PrrRi1clQEw9P/+zJOkB0zr2a4l
b7YQB1P1cA/uiaK7ps+GBTbe/fdeYNQ82asesI5/DC+uk0BgOcuRR1ARinWiPgYb
Fcmd8a0J/JXTInJbfGAunCEN3TneKu/h3uaSRkg2W9EJb2hnLDFPUpyYTztyOZHf
E71zkHuOZ8D3ymgxvO7b6x+f1fR82pPLKQorHqA90e6CcMTZxCZR+uoghHnO+o+l
5bXBxlJzp60nYBlNFZYySB3s8Kjca9HJzxYIR6ktoBb0YGwfxq+ZXiGLHCamtyia
MugMOs2Mvjxb5lXuL0Eyss78Ql65VQnKijDMyPisC0vMZQNy2DE45uOa2fIw3dLz
gG7B3OG+QxIR75kosmRZnUNjjko3+8QgxPgrzvn0hlBrVKPwK36Pt0cLbJU4+6xL
w4ZvRVV4V98ehc5RhfD4yvWS1OykshV4LS+QcsEfuPAP9w3MIuvgAAUjEcg+C4ib
jB0bOw9OAkjeUkXhvEqSjPKDsrK815VWn2hb3BABQ/F0X+uFuqUMImxmR09k2xYf
k2wPiw48HSheS9AbRX7WfVuZngi8NYjsjkF9njMneuduFM8wQyPUmBe4+KO6ed9O
1op9OrshQciPurEPsKmuVxSDCKAQ7ZO0wYLruyHujxNvRHCcPtsdV2iwBEDXhs27
UkWY+lC5QLabuQugQT0SeHO7+gERL5QtvrUaKmQOVKCHCjsdAgfJbTuO36ZlmPbN
+qgdDrAt2nR9qJbsxdqje4uyOVHOYVWt3LIzIgMKHkqTIEEoydqUUPyOJ6QUHl8l
b1YTanHertvEKgij68WLMlMa79DNhvpubx9JqqtDW1cXHsGNw2qGYFpKP0wthqKD
b+R8XI/mVpLbbpKchw9mhfiNfw9gYicLkSWYa7RNsQDWbtr9arc7f2gp4RJYsn6y
Y+4OwaMbxDC20VOh2473nlpqWnELt/4YK4aJD5mJStG5v5DKHVN/la3rGRHSaa2i
M+fntO9ekCDKo/BqEaDvwNXF5A2U19co3GcIiQ2YFkUbyhZnYkxDSJgJKKqDEd6g
p7NLnjn1CnCrvUsIhuXWAn3iRyJCsaILCiFhDuySb7HdgcWzpjS7NQbBSCL6k8MG
4MAW3hX+DvN6VVzIF+HtgJXFYfRt+Qy80wVtTDkKOVJYcT+XaHRscU1aPapQ4Fne
WeGFMhxhh4FgRlTNa/XxgCLOeVuPbguVtlYW3WzX5FhYI1udw6Nixq+FgTD8bLOT
8asTxbCrIRZ45pCZ/rO9eiOBZ869b4IHh24s9LSpcdktNUmh7vSkJU6Stdtga/Ol
O2DSzJE2VKASRE8lsoEqeDGRj6jNNTOsgz4bd2bmu5xTAqV3DPaFfHcj7vp9u1O5
MVCGSUUSL7lAx1XcuZoJveTKwzR39CkxaEY3P0cEhRS6MycJzZe9aTBnw+36HWEh
oKNxHBsGkmDlawTzu2GtfNM3OB98g6xtnSnc/oZGX48Vt5NZqTSMKiNREoRACYeW
fTU01ah5bvrk8h280fJooGO8rActmRMn+U6p3OvA4HMyRzUrPHsAO9LI75zulhXk
MM5uPd22SYpyztTzZQbIoWi22IipNdFKDLodUnXq/BOpG4dGLynl8MV9w0VRz68b
nDBTY4USOgMZf7XdsioN2mNqhpd6EPOmDb9OCy4KCCjRXGkYauwxWKB8bixssbJ1
VgJjxv2JNeIQaYabm9z9/CsMaL2kEmsvdSYIC9YNSqYWi0WHaJEX7YOJfNVsj7V0
U9fvN437ngTMKiTGGHzCg6cFP6MkLTdybW91dbS+rrocaSCn9SeusoYbGDUHLOIx
CUOyIAs+K/2AYfoWOL8Vi9SvfverRZiHkAy/4MUibaetL9k2H32/H5MCAb+mB54i
W0FukfSpMZal7FdVdpBynrN0gzkG3Yw6plw5L6fFgh/Co0YZS+U7ptCdukQBipqq
bXaDtaUHMBTgNZFIKzUXXkVPsLG8t54gP3wbbcFm/yiSkqClzfm9r2WfzvheqHdg
07rBFyeyx8y8V/459tqQoqJOGQiNOsOU0aPapbET0WiQQPUtqvkHau+8Pjf91e4Q
JunWDpnhoUttp/ok0xTEd2ysoTDd4YalYn3EDU38+eVW1cIwZSVMkgF0fGzqFCJH
bhijAnAiVuBMbbOfg2bVR+wb2G2nxJmkxwsTA3m8Syk1td4k9F2qFWebgjCpe9tx
Lr1GGq7YdayKNALo6cUgvrA5jx2g8fIhbVVuGkSuiFHs0xB4rXBlwYzzXol27fSX
y3VoKXlD/T5i72fI6gMA0WDoP+foVi25OdezaPWi12QAfpZeme/0LPDi7X4ocRQD
O0xxIbndTMoR0oPmZ7JSamZxPnta5m+yyn+YDDZVnFlE4/mpxgGgShaRaJWGX0WA
05PpVrVwsNqhIEiHh+SNkO21VJEbIvGLlMX10IT7WQ41F7ccPbDPzQtONjqultYu
8+6qBXpR6Iu1m9ByCwSAhVrdF51J1E4+PtZPIu1lVXBpO4fd8JLNaxk4bgZNW85H
rKOmEeW4zpfJafn0gzbs4wvXxkJZmFhxqxXbSY3jRXCNdpLXrgfoT0CrYKjxEbRI
9Dw4ts8avXB9RtebkM6ihYlwysVMx/oULKCqTen5vxZrX8Iov9pj8MmgG1tKql0n
rOQA4RgrHNMcYdjnxpIsHxSE+1ui1SslW0dohqQeYsv4E0Mg3/jkcK25kXeOvo/M
ra3CYeujgU29ApRx6g6mi7jvIZnwwe1uIv48ihUVL5iun0hGptRuLQyzTdotI1tO
TFnZ3Pi0gIr8goyXOew9P/6hJFMAV6jXQb97cOeXiF5i+EIcCii609Yz25Rms+IG
3eQDzFbVHbqBH/1O7CPbqfgZhFBUTxdUzlfaCYsISEHOWKotdUvxaDYbH3L+TUu1
Ag+87BsA3OWeJTLc90x8N8IvaTvpX/og8KSq9sd28dw20x1lODN7pZN6cyB+Qv0A
VsaFjBxdNd9Iw2Z4UZKKZrgLP+D3nB0gNVKMN+oO5cSraJOzsFqF/7XwgVeoCu/8
og6vg6Xa2TXl/eo1B8IytBvmxiinXVjkp7k29tQBzc5j5O8LHKwnY95uB9O3HyX3
VRc4qXRzeyYvhzzZHlWDe/VQqquulNqnrjiP8nlmMbCJj5O+URvlMDaFSo33SwpH
mpZ1zwsaM5BgS6buKAoNc0a6mhpWcYWtqgCwauRlNWQJ0nlftgTXeNKywzyFgetu
X+hvB5Jt+VnajqUOkkKDnFPg/rBQmuW5CLG0MB05luFYYgI4UslvH2RuKRC3oVFI
6Y5kvLML8Y5mBknO8i3C1MWId7Q3G8b0PsEtf4efh2x7dTH1/AhZQFA5xsaycZJG
8DoWC3+PXkzOPH9A3PpbfWpfumAxg38TwQdLJrpxdKVJHPq8dsSHB6HYNxxMSGZE
1mmaJ58aRW+MPdgQolMb+nva81BBUrJxM0Ql9uVvQ5zLztGjzVDPRaB1Pl3lyof0
O1EKvAhA0hx467HiDr8tMNcLSfznVbz3serf058K2M405sWVOKnnUjCmoT536dQg
pNwDdD7UcV3TrvnziteZ186VTAkB/HGd6mY7RpmlGs9qL99AOcPqTtU7//5D1ZVH
plpYXi9J2bC5vxvkNzduDD1gSXB8trDwu+rB5p2jiqz7OVwaTg2zbZm9Tx4U9fAn
o3TjFb9Zrn0xgvVkmmtADZDUirDKzI+1Y1eyXv1WPmrR/IgT0Zci2Srn4HxD2hB1
ybr3m/xHZxI4O8Hb0zyCtfRAFJm9u5khV9vWsGIIDjovC/AkDjfHghsyFFKs4J+i
D28FHT8UU+DGrWsP6PWWZdpEQlVmO6gIjsDx6eTT0FNtAY796wJz2rCl5u+TIHYn
MSk6XzkptwMHF9VhTRLiZ9okR3n5KWkwuKDA1JZYzSxA7d8u5Y/OR9962r52YzBY
hQ8Ac4TcXZRG25eZc//d4ypqoHa8nYeay83O+BqOrwRjW6UBRDjC9HbrH6zN34Kg
NIt6bNqjYATWYpg04gASGaU/e5ZeLUQlnV6dVeUb5ufSwrzWRsgylNHTjya57NlN
5me1xnulp/KLLvfRfLW72OvN5GKCtT76PGeAE378p2DnLvklnxByo3E33K/5Q9A3
LnDK00q6DjdZ2ZYjoK+DNaFAzaYpHsfAJM8MISS+PRWMxkk58WA/J2rU9BeHXJxX
zB/pV28MxN/SOgX1xVLySbqOzAwkUMwnVF72vto7cy6M/9Ool9MLjz0mRYO0F4Y6
xRmll0pQCBQz85LjkqMiFOJHgT1Ol+BzlNWvH96hTh2yBMJT3PIxjLJ4mI/GqvTe
ij/vxOkm4qEHVfaWsEyy3HrltvxbMzCbaWhJE86AQhm6XO946vET/02vSVQf8XcT
aTLIF72JkysepxzNp9DR4qGAVkL7Kstvzhdic+5BlgBuA6zymDnzmGkeMkIWIzGJ
yd2McPTdBNo8sp5XuHEO7fQPqP6EMFQFKUDWIfO0hA7GbYXDfvY24Gv6ZwJz8njO
iIVfcUTwPvAd5xvcI1QdmBUbQu0MFU8knZN0Y5KKSMs6R8FvJ8aYuoX2mVIfkl86
OTvO4R8bFOAVCbLlGMXTID7FxMtQvZbhtE3pyQkbFBVuJxkLDsHgwCyYCm5AJb2W
XYY1Ej/i1TXeh2Nq/uie6CyyDvCFahT6y5RgR7wWT+/8R5oY91qhHoZkQrhlu5kp
NBGizj90ZdnojHE+8x6zYFnOelVdEI63xPzQKPC8Wk5fyewXFjfYgj6d9kq4NKFd
ZtwT/hBl1JQgP0GrYjyJ3LE4VEEjYOOVoCVeKeNAwoPp4ugOJrKjWZ6LyoEErU6M
Wa1KE7hfzBfNUoObrc3t4sREtoqL5UTIiX6HGxX8VK1Rs3bkv8mm5IgfbLsiE4fg
1oAtO66aK/8B67EHGGikKOkO80+J8HYKsjBNCZLVo6Kry/W+zlKAn/tDety07r4u
Ampwz6JgifIdYWi+ccEvI/FNMWm1GHZ6DxgHk9o9MqUF03u54hLbBy13XnUlLiHc
QQe01f2hFF4B1z0d6GbUj8GFlBaC1I1RzuVkOagXIkJa/xV/92h7zFXOx/Zwh8hm
Px7R6kqyR6byRS/h5N1mrLjBesfqcIdqfN3xniYxkiD7Jxi32wtgkaCE6xO+8bsq
Qnl1r3i3jZcmhFQrGpDhTO6Ci0QGz23sCiyxh7WojmC4Xc0S+uN9BTkW1Lg7g0P1
EKL8J6n8RilbfUtxeMQZLrZbLNpD3Tq7krH9Duf1rGokb+ix5Ef3ebvVhi3nI5UO
1xoGwQeBlCsPKXljqbRqCUKmi0e0iqYIspQLg8RSM5uBLIL1G07czeWd0VdoGEkN
PdGeabeXK2n2I/rEOeQmTso1vrJt6ms3P28T53B+WSbg3Kps3xm8Z2CfhNqW/IRk
uQDC1wzzL/6XHJSP4qP/PRMYWKpyY7+JeuOb7bhld1sPLi8YqKqDyWQWgemUVnub
AR7e4ZkrFIIx+TUL6XuxxEre6rV0KUFdZ+oXueVsaKOQTspV3eNFwyDq1pCWu9AM
Iqx4HkxcgME4D2CHvLoQpkDF6Ix+SSwm6splJ+5lJPVfOa71CyVpQPii0GVk8eVi
9FMXAGpBTv4Eih/EaHUKNYbktBKdi0FeL866I1ZExFYvyBAqkCg7U0St5q+MLtYu
MJlDeG7PlL5HzudIyrLMnXxgsLckLOvAP5eS3RalqqtqW5taHxsv5o1kxEDMn8Ab
VLvxRvLAmbH+uamkArEHDfZL6AMjGsv/oMPPPlcLbnuDZtYJz4HBKRvW5jVdFaDw
hb1Ti/2zwwTpFP2gSDbHhq5oKyGVJQL80wsI60CGRxHtvjI+ZHTIc1/os4cMyMQ0
qHt2/0dEa1u2GvnxI6az3f0vj71lugIIB8uzCepvXx5SvPjbx6AwlhyC+JNKq95w
gN/M2ypfYl8V1rj5ggDroMN/XIWBJN0j9iR6m+jJk9KxnX8ZLKBAe0uqsnjAttte
z21H3BxWeJJFbU8p7ZU4yHRHSiBPIS/wJpuEyrxg+YgGcnU5cC1FbfsadpG+7lMe
krLtt1zrCCUqRg24pJg7gjWcQnopUsQztwTyxG8TWY0XM7K6hJvTEU6KiKbMTVG5
IFKyrqHw+65tOK/hHQhoT7O9B2q9468xZo0cEZDTnmBSCFwwpOSiw7A6vnwf9r26
0eJLeGSYWvbeK0MCvXbvNTxyZr8+AAvtz1vThu91gnqVjsdTnVfVU+gT3NNvxYkr
l/uB6YJLJoBrAodp98WZ3gf54khg89CrmuvSNhsulI/aMmGxWrXeYwSbPjEJnYZp
0ZkLv2Uw6KIMNvM3WrmxOMepvTKsJJ89jKQKFD/9EgTlH1p+7pHVvUtywUeegqwK
5P756u8E3gGl7yGBmUge4nxmH2qy8m51RMObdPjD3/+lrWKri0CDbKAJ7jQ0n3xj
tmKtuWJFYmOOI9hvJr3oERzWTzRop30DKE/hiMniQj5m+biVyVbM36eoKmBSmelB
fdJsQEpX2JJ6j2Y+nIBctUQi4Wfqk/uVD/XjO4HAj7hu/qPaffu8Ttxp6w6l7Z4G
AWdQxcy8D+7ov5ErMSzFhw6VfOpVELPqzV0o4UcUqAaSOdFq/cKF0ZK4yQx6S0He
GicX+DQcKbS2/fyraaSgweVI4klZyBsKTyY2/xXOn6mebS96RlHRjN3ib4G7odjm
sCzLK/Ue/A9a1LomH94KMY2v8nB+u6VdewWN5MAUpAVHxLFlA1KsVHQPMYmjkPGT
DfC9Dck7VDDXamltuesXTOVdz6DzIDV2O3wuZH3s1Tg3Hi9Dw5IRGswGW8af+BzO
bMzjvB140x8aBbHkisqHiJJJioepRaljF6A+sW0KcZa5+adjuRWW7vXqNQS0pXS+
9ntcZvPlezhPOt57qIFzzNEko+W4M7GiTLg+On9hzdlcLe0q5od6MEbP8mhuieoU
DgZlnN6NYA81pR/OfUQBLSmnBLwkXAXM0+zjEMNqjNp9kbbXWNQyXFuqlrCJx91B
YYtjShXU2k72VyY3WyOrNcAYzTV6iDDqlt5XCUMhhm5mHFStTvN4lTEFGPyrF98g
LzAzPiJ3pdlidy48X3onN3Gln0+Y8q9MhvqTtRhp8nekV8jBX+SOE8jR0Zgy2I+R
h7YUJMae8YXd65Rl15zy2mHip/P6oO68TGinInTs4cscQBUr2RNoMjo/b/NGru8i
9w+fQxUINNR9D+X0Ax0zpH9Blg1zPy0yKf7uvcrv5Mt+acGPDkw7LLJ34zGgIHvY
ENzOIZ6KgqjhyRpLboBxZyBWZPnyo2tPZFuxiOtjcfSq5TDByS2AXVMiC1gQDDGC
R7SVB4JxGpq29JK5mX7ze4qvdMgzF75a5hMNumv/zQPOtbvQglA/kCRNxws6bRc9
6wi19Vx4LR0+nNiQJUkoWXVeUz/pfXzFHyIMW6KURlO0TXoJX54jhPnvek4rhFbL
JdavyuRByilYoAYWO3q3aOLPAB3K1bOfuV+JfW9Wz4VyvqI+w62ET7Q/8Z6SnT/y
3kv6yd+fhYyPLsiDxDc00s6iqM4l0ABQyd6uf1EbtJxpowfMNqmnaKqEIJpw0Osd
2tq2+BBeU54c7KrbTtVRK8CH2TQu6UTCSbqJ34SFuxQi4ApMtkaxddPDb0WfqX2y
SE2uKBWXwUjzAvT/Ja36oJfdoGgstoyohA4mYPoyogpfP9c14DeSYrcalqFl+agg
gfMV6YjpCDc/wT+598aZuyRcCGzCiGZILCsfia2mC61ndim61i1f4cgEAPlrcy2F
ub7KVCSNVU4IOPsk/GTOE0KihvAhkuaFWorhcsGOKQIz67DcJ6nAIW+r9N0Ft/aA
9ja7irs5aZtlyZGz4ozu1RKWfDi7pqOjrmx+TsYBN/ehy0+zC8i61maqI8nJl3nN
AjGMweWGdu7ePpl9v/UrqGzwkbrZvG+dAC+Hp2AuMCQu7HG6MhSa+vMFzKo4Kjl5
rkATwi5Qwwj1RaU+0eZqyGuAG6ackqv1H8gICMoum8GbaRSTdWyFqg4eS1oU82A5
WU4xacPh8vn7C5DNTSCD2OvqlEFxcvWjyOd3wInZyikFlHGqPWmqbINrpLUD5evh
rr6NznlZUI7LFuuEsIAN//eAwUqDUN++yulMnJuFvzWzCVGfI4BtqxQsfYYeW9MX
j9eRgUKyyGsZM7JUR8ZWCtUslT8rJZj7ITVbR/5eA/y9zAIrwGTakJhVNdJOim1p
GlWgtWf019nUmoQeDbfyYALnF/o5Mq4tsrKPna+W2ADw0lTKfaqzGcrm0gL5pn2h
ZZyaEuoEJe3smJ5pKvgPpOreqsv9nwb2Tfv3uNRuonXPaxspQv4zWJ7Glj7aaf04
8E8puFQv5NafmUTKlmVyioLHGFWoESyU4EoWJFsKnKy5a0cq46E3xPpNf4IkRFPb
V2roNjVGFblAdWAfp99aXCxF8LSqyZqKebd3VIzTw5mOX8WsD35I5JdL8UWZl7wZ
PI5XWRNvd8I09vrqrLehLIdT4tr7BDv7U0s5kwC7+IPRA6FjULq3babtMAcsaHGh
JQ5v6eMX2NjJWJOYWyMUBOkjA2VYV4aBcJpxA81C5O4MNsZGw/yRhY+ouo/fLy6s
C2MO+lB0kk3jzWzAfBWTTuw9b2U9eyNFp8QOiuFo4VfGztFzlOOd5zaB/gVvc+pB
0+y+WvhXDfzl/h34lKNpt8WAw+7PbJIQlfqtjHa/S9Pqq6Ayk2UpzAxTsxWv1jXY
bSOIBaAL1hSnf9mll39nx7QtuEZnX/Lc8mfw/V93hOo4stzzLXd5UX7raHj2k6rS
BZKkCHQZ1jED5HvI0nLu1Z6103oSE5zwaDZu0EUSKfffzuegqezF4vFxqUQ5VdGq
UtsqlMgh1HqaRHFLA2Q2WvB7aodjJofwNiHpJxpILXWYffvInzjLzLHjqcV2CKwY
OMHvjnfmvwzG56jQj1z6GhiOtij/pYPhph5GQxR3EPL0lCAxXoq8kl5xrtw6J19U
Mu6+GsnN92Gbc/Y9Is9sZvclJdk7mPO+2IKwW51wRB6wk4zoE3EXV8p67xFUJVNH
iHg747FM7EhBZzr28hH2Ns4ezPAOS2+gqCXtJf0aZOyNDSyOUqniSc662nS1/O+V
ufUuACufHp7r34XzO3j6ieun9N4S0aIoDnFD9QluQWADkpXD3w2JyIikWaZ12efs
oywgQB9Or8Fh8IAP83D/cg62oZYpZL7lmxcTX3aTqRc2zMUA3LfkpNGIxrRATla6
Ed2iFzWLSyYP0443wHqz2FBGQL2VsApSyOTMWWgASFQF5qIpX2sPak+ryRmfsLAO
9t8JeJkf6rvbK9gBgarhtN09kEEqiGccH5kJyHM4NvRd0ErC9d6dpEXYVe1Z138v
udYJzJ3s2JTAun4cXddp8eT+8mt0XovswqczBcxQsdb51phAa+E5ab2XQOkPkPKW
ZJjX2nQ3xaERDvpI296ACHHk1mAAqX7dvnKDo/txyxen4oKljFKn/xmdnMmdsx3W
ozyn/NVqhkiTFKeiGH6ZWmkbKlGdTBTX8jlfcbwaWcIUAZv7ua85RppM5ttPKYfB
TqA3EgvtOAt3G8vbi7mwq1cQQH1dZAXXHVh5NXT6yXT7pns3D11IXDQ3EH2c4/NQ
xqLbWomyGOv58thZtOL4DJDfxvW6AgKECRV6iuKwU3k81TN+8DWAJ38rgP2mh1JU
JxupjlIB/NloCFR8ia9W+6nf8C8a9Eno1Eaj6+fISvblc/vHIOP7vTsgMFpiWNaJ
OHZI9i7czz0mREQzdFvS4gXdfSjYk+jV5FCX4i/xmaQfcvMLPTVRsAq5+QeZ9p2Q
yEd8lxChLNd9cTVOmnrEJIy03YItkut8n9MuOBSb8lP84bX1GdxhDx+Y9ns2y3jR
kA+UXkv0bMsaZnNxdq1sMvD/H4WwENUNkrrplGcAyYDMBkIaJijY+Gtk3z0VPYwz
E83ywaYS3b4Gq9C00RmaFGCLFa9tSiVinvy7OymKI0I5ao8MdzjdAaPgmHQ6i49q
ipI/CFSc8taKKacrZb9sxsgphrhIQGbh+SO9XRmAzFzQSqbCsHSpNHVeDf6Hi1m/
xUEwKXaeGOs7f59WrUukSLhhgoJEK7vP99P5Tw2UAP5WH/eVcadKa4Hj5ka43A5Q
86lxURIc2GChs8O0LSkfmJ2xeBPMj/VGsv79DxBvHSPPBGrJmoKOqbEnAmG6Po7P
b4wNhAC8XgRBWhs64vAVy2X7uz7V8IJXqsAcKPi+7hgSt/obSQE0NepyFVOh3OUC
mOCm530Bf7AqKTdYzXLKwiouPmhJsBmNm+46g41+iNjCyUpfdaS18gKBM5OWszzZ
tDJWdw68BSj0IdVCqfFLHt3inUYij7dZ1WOP7Zj1O6tsLJYnZ04IQpjjBaRBWxqW
LQE3J6RBZUmXYY+jNiAaW7Pus69R82drwMbQq8zJVrFjSGFRmwpy7C1T7qWKiSBU
s/je5KLF4iYDdgPGHZDFafBwEB1OKVSkxbdffHP6z1tRHx+wlk+QX63WMQd+uan8
6cbjhcyF6nRdUpD4gfvA8X3qL4AZynGlfX0y2uqc6qYorZEiM339Mep/KbKKTX7H
CpDePI5FTsayEY1gUzBhPm/H0lbFKyEMTrGLdt+pB6jRZ01tVNEHnlFICz6ZeHz1
+o243CvQNkFp2BU78t/4IeYWv+YwYGSHHpX+WSD98Peg+3OZHfYMydi5m9aDWMwK
S0ZDMpQ3KDeZ43Lu1K81GO1vOfy5G1qunrzVXEbGYxXoRLsf9xoGb0zduI/mxXQg
p3Vp2qnnZdNYltiwbco0v0oeHudbZMFl+eHaFHOJeK4wGCi/Zw1rUX6gWrmKU6XU
zHDW3yV8WNEp/0KiiPsrjtMAQrd4ov24L6BuEhYvXEUdETuSCielf0/XNwoQA/NM
+s2G3r4/D2YH+nLaubvXkqbZNTsqQjsqU7IZktPwWnLEYe4NZ2U5hJ9zDS/pBAzA
3cP1TBSo9EjbhfJcTt3C/OitS8nJNobPrNokUpsWNG3S9ZosXuna4E4FPzV71SSQ
JmynYsEWiTRcdw50rUudkjQk4H1naTEBuakhHb7gS+ArS6CgsNSvJNpvVYihusEc
GW1U0NKhYCPF7upfD4T+a6zR12y0xEWaodC50rzhV7kBxNZR5WR+bGrM4S2r4KiM
femJQ4MjOTW3NEizkXtmGpYOPgjPbswnqNm25uigr88q2XZiF3tGYWGDmSFwqEv6
DOyKYsLoVstfP/cnnrc81uMDz2tA5GLOOq/hLFzWjtIiA4i2VLPmcKTaZRxCYF0J
9l9RP2ckjPbz/+tqU1vKmk9tWNfKxzN9p2+jjYTJFto8Q9fn0HPp8eRGYKAkqRB1
bj6djEqW7wpE2CzauvCTIDkASLLlECg/XP9DNlvEQJ9NMZImFFVpR7yKwv+78tQC
kxfG2atU5W7cnRUHwwDZYioGzwj4UMlRFo2MPfhlAAToazfEgrooexgM4YGqrfSi
Kj/43P2uEEn1bqVt9aaHTybC7u2n6156zteHparhnllGx8qhCrpl1PsEoZp4MaQ4
v3kxFLcGL+lTKE4HO2Jp1ApU5hOdcpU+LS8cqAgQLVUoYi3pwFaqNOfIx9mDKlhM
COhXxn2MdXVDPQ6dgxJqM/FFqItdXSaxkkMuxordOj+7lunctRz0+jUEHw38ao+L
XROVrSxXUuTz+6tldzXBwqEj5t3MFttcHKy7ykH2R4me3QFI5CH11KRzne+FjIDt
yqsX2dnQCuDg6iywAZntmmmWNDTxcuaWCmJ0NFLUIjvVKx9jgw9xQqe8sJj3/Il2
xVvQQLZpWKBqq3NFRc63Mr6nRwjT2vJFOh68yyL3kErsoiHrKA2bsX1liFkodAhN
olOIxPZqOFkfrxNHshvvK9NDYfq46dHMmpQsUuipGykqAYhAJGIrhjPyduT3YK2F
hh6KZBqQexynr8r4KD7qh6ksA5o2iawGML6N9/7QJlaqBBOiHVtTnO+FwaKEthgv
BcRBTLK5GrSezKGGAEn0d3rb56aD/fY1lSawrUrB/+11MFgCo0Sj5F4T5B87Xxl5
06R4XxkLAkqhc+LlZQq/827hZbcTQbly+iGMza2p1NyuK5asRX1m1TF4yky2CrOe
f6jrC+8VwL6NnxqaMNSIAmetEX6m+KXubWtsZ0tG3WLkJW8mjMA/KJPZscS2Mh6h
nXB1ecc64/RaGBeR5luPKejfOFbs9WAZQudny+qa5ku+VnHeASSfjttlZQrZc/vC
o8oNalfIBDHdz9S9pC7j+c7aIoeoWcqqizwCjYvexuc79b8jUlWzGaoZpLBRXiL7
3qg0sDvl13YNrvZG1ymbA9FpPaUCZEOzY3UIbgmioY18Ame1M+/9Ev+PrHJ3qyTD
NSUzePL9fjkemaRzSK3/Ju4L+CpPsRZnkNRos5qX/lcG/vo0qznH/S/xEC/znRpD
+Ya4Iwv4QOrjaTOmq5ksWm4bfwtO4okq29gB1MfcEe0ieeSs8Lawlfc2uRYcz9cW
XIVjtHKFig4vQiETxfKvWLFCynzi3Qb6A379o4/yHnXT4NFVZ+O1VoCpQW+Fwi2g
h6u0KuSZbb+TjXoIeOEuE/nF0iVgLBT3iBZbJ0qw+p0EgpCGT3I3MLb3vQ+paSfR
VPN9FuzMNiNGSMYDypPJoVxpTbOz21OO1+P24vg26q0+z1pWyggMMl+R0Lsw3QA4
k0SWjI9SL/SKsR5GL5DsCCQ8tS7mf/BVqDckDtOOI0iC5YgGj1brVGO1SzlXd08J
JzHHiB6Owm4VwjKPZ1fPOu/Ri9ZfKQX9Nef3DMbqHDN76IbS+8zo02aZ5nVCvgIX
KXVeo1H7dvZSWUyT5UZPBxjGPJt8zFsVuevXaL8/D/PxRDPzTHfxM4wL/o6dAoU9
MqMzzNqpXRF8i2k3dVf8YyWvPv4zRBFg4p4a1Rre16K1ora5NluFKk3Br8YUE+qs
0GqYKxc/jH6IhaKzcYoYkSp9+/jBJ7KD10hAG0K9vgqEqSZwdg+gvaCD4cJRwiXA
+cOWn05UmBJRGFdxiyGtlEK2FNW1KFSRDWZe7tBwnHSt6WED4GIZH9ViHW/FL/4X
YQm1oid96DKV/cJMXTrOOdwP744LqqQC890B1MyZOkVU0QFFOJ0WvebxTayRmwtb
VPbc8IohnOelQSOm6SyKImKREsjf/ukf84W4A2QySH6U5B4azjhLAlvUnRxANM3a
y5KZGypL12DnyEP1GYyn9xJo2x3nrFBj/E3HZ0pTQ11sGR1Tuq21AX8otBevZG8J
bHPmpEBgcjJv86P7URUgbSfjhu0726rD0yn3G1E9a2nH+x43I8R3Q+aUov9MOHFV
6AqjmHlJcPNz1VXQI7bMQTaW/y6g4zqN0AZxZ/J2X8Vy6qJ5TmVMguYsCh9X6Z5o
RiI8e4hy2ZSmMLNjHZKgz1b5fXztLdswNlaO/MtrUhUiLYY93jxEDhBMQwpi8rm0
1MEdzj/pRL+jZ3Z72hXeFM/wUrAruJzMNs2WmD4LqW1ARvC/EnCqWnDOUWNN//Pq
uWF/BKGy6pBj+6PjbVnhzbNcSr2WOE1g2Ns4TefNPCeORiWccc8YGFKORCcIm53a
f3ZepF6kxkj3SfsLtZFb3GVlmvGLApgclDXNfgr0B9WzLlNgCuGghH41G4rYt+UU
S5rsRfJ2+xutOK7NzN84Nwr42GxE9YV8NHutJF7n1vn+jt6pQbPQmH1YENDqUSm2
xLXfzhSwDaC3d9KzaV9bdHlbefLMQwYqHjPuXbrX/mr5jeA14H+jverRyl8XoLPp
5KAC8tSLuunH55Ade9QKgl7A/w+V810LVj0H5acuML7zrVgiPTYCkJl0lUBK84o3
1yF7Tjk3QqYH5fOVWDLAv3eC3HIUBS+eBzyWY4CbVkCsxMwMMLsgCwGKlFOjXb/a
6yNWBhwGqfcXFABhH0mISzkJYHedRpelzYwy2zwx3jlqj2bEWyn3lvgVABcqBCuD
hzStQc2sch7AiqYoarFuDM6puhj6vvuPQZbLbKqN8yDqbai2Ml2BfJTXigeaiq2K
slo8ihwQ6LXefQUUWG/SJz8bv1zyUYrileQi5Wo+8L3dWYRGjs8qEHn4g8PS9I6/
PAk1tfnlLbgTHlF2j8re15OoESPTM8+PsxoL/vNTzLMmrlURHOWjKr8MVjvDd2BU
tsnRZ6PthTgNgEpG7o4OZqdef361QU2Z6p2wimcrVs1UFryDUXocOQf6Klwn8kZ5
0N+hQ+StnXXTdUVKBDL+LaETBOfJdiNHfBd/HDiWHvwGVRXF4FUhnm/iOOtcMlLS
IcAnB8V+hFL5bwJtGcrDWnbYeLMr/+DSOBX86itEwRxeKRERoFdhqXM3DRbPVk8M
oibkEHfzpESIF6SCHjyplrC0Gi4/XY6GMQ5XVlHd+rm9oMJytPtk3c2hvkIKyZ2t
HedKILlnvqsSlcwOZ89ND9Z7AYNnW6QH9heb+2bOy3sPMp3DfdTZIF1zeCHWav3D
Bt1wswvpT7g3SgQL9YKm6CCd5aWgMUypyjnJY9Bj1yfslE+2rprGwByZ9jbNqher
kaiCmHgrUYm27pmLB3iPqa7uB2EIgwlotifbmwlsGbH7l+Si4PYD7U9KjbNYYJHY
UxBW1+ZUi1JMmAA243Kg7ewe+YiTzK8nCR0ft4EOy0E9oHIzpTZCQ7qlHSqKNcOQ
pBd014Pr2RM1jO/IzziknKKcqdDcxoHvT7sS4Iw1oUm7f1OdFz0eA+IYH68ArhR4
dZ6N1gCEUHoKnDAvL+Q2HY9jNhkenUOuPdOa/ZLHYwFWFj9R7vwjSLPruw6Wztum
C2fa+gZIWScxD1Tt6oMF8QL2vKPBsKva2Pdbh16rA+CBs2i3g64bL6yOG4W3MNbe
05P74p3BNJIa2cxIqRwv2kJ4vbj5Sh/5twgJeWQR5WeUNPXAobgcYv87VyCgAH1u
cPwSkjAE5N/TaaxhMNYOiSsfxwcksgogB2d7XnAneKQ8gnJ0rgmu+inkZtzcbxt4
QDKsVVFXuEojsD8kKI5yWCXv7ba3r4GLMXW1a06e3qFA8/SDiWGqqOUqRp4ujfV4
4PvBtdTsFV3X1u8h1jozpjA17L66ZAuuKLyVewK/ojxjxh7xPq32/8lzXr21fzuD
bCOKyqLJhRTH9ftBnevCCsgmD+6U9v45ym8QUO+Iea7YzxHytpAZvaVPsFwCH9KR
6qmZRoZ+xg3oQ/vtZI19vYTwmni21R5D9HHqM8zPKFxCwlLDjy5OmaDH178q41A4
o0UWCp7vsn8qgG/Zr81rpRZc4b0mB/PX2ocshrnm0kVoJU60qh8Y9eF2CXGNo08b
2HvIBAjIO1qX13pnymJ2Jtj+v69tWrds6zQO8GqNJ7Ywu0MsjFB3HerGDiJW999C
QsGEOOBSGlvKmFUYsleUgy33VT3ee6B0NpiVOSOYdRjbYroXlLRD1B+s1tKc3r7F
oWmFHce1Cd2yDD8x2f1YYSa96pu9g9JKCTrRl4JghHcpXC2YL5icLbBEFKtJ3teK
+rcxnMM8ZIY8gATbVYocNkVmcAz1GBSII6C6rsXbOjqWlEwaOowkBhArdGG2oH3S
JwTZE1ncVjDZMBO7Bm7oWzzEhSVGQepM71MowBb2EF/Iovpij0WXpCLgnd7cBn1l
dk1eoTuNJr4jGEcIG5mpdvcfm0IQ6X+J2QpDgu5TEhWTD1yZJ3CmHrDwJ9B/ozu/
A9kMs3cYVPdRZXj2Kj0WeRsc7Psfd6pIwWCOFHYZbq3QgrUWzrqcjzeIb5dbCpQS
ujJb+JQZuCYbpA21EgCpO33oOCxm8YhziT6UN8yXNM7U+n23JJkd2q38yXKnwh+r
rfF/atccRv3o+UhprIZ5H2UZzybE9c3WZitib9C6Ogb+THPf+jt295Pvpvb7uQSp
5fw2Eupf5VP/IZEmFEFNdz7d022xM1v6tqzOxEqiOcldcmzfJfMzje92cJTLUmVj
1uhI43oDCvfRAI/t6FkkxST9mkZuLMOvALG0LE+Ql+9y4EeGhoqEgvVyyUKRP+aS
G7EjoL6Zi2Qi7Hy8322F1ibKVuf0vU0pU8qbFhdN+eCIG4NyXPE9/yJx3VYGtc2B
dnUjoaKrKEXQ3lrbY4vEOo9ce1IFVuBOXdyFLs1uNxt4qbbbPAP6bE3CawpqL9nL
Kcm3ofD4dh7C2pX4LtqAxnDZICnhPPp4nROH4LxSsM2qWeEfNy+knPX6BWzxlQ9U
uo2DiQF/mtNC2Sn2rv0qLAVQU15HxIBYwzHXyedM4Jl7QCv7rl5xGYW/8qziC8EE
EEZAJuX2p0Lwp6GsapxNOhViH/hIRx1tWexyoYSJXljDYv2MAssv2oClAEE5IiMG
RUyjOMIFD5oR4ne612MwbOty/FnRQY2CWDFSDPfDiXhfmyUU/y7Ba9rFcumIQyZJ
P6Vae7L0nOdQhNZUDdKQKg4x8vw6EpfCaKPqifTEz2Wxx74VWDt51L/mz4hKiprx
ADGCDjbKJrw2I8G2O+RxwAucAapGsXMBp5uQ4w+pXUbc1nvFivJ+DTeQHEJY4Ffk
jyDtBB9SL9jNWwZfZYDKqT2t4NTNA0uDhdWzSx9zIRq2W2oN3gInk9nWRuwc8mxX
7V/9fRWNGJ5jdtAnnAmbqWOS4qee/PmHJJ6tK+ftcsX7Y3tH1cjEhkL2oKNCNt9T
MZHB50Wc++3QcP06WQIZn0aCUQryP9OKkzvp/sX/0gyXNuCvf6PhOOud3L02wtGE
zewRGpHxYJ1T5DFYTT2QYpwLs26i1ZGkDvBVkOPlYGZB9G5H9wIu4UONG3Cx2q5R
5CVY/tcO/ods4KgvYfWPUsiiacsrTq+OAXm9JFzsoJ3D9zlEB4Qc77dm9JfQKV7x
ZQsAjIgFaKTXTU1wlMA5tyqTq1v5bHOHnTbIz6nGhtXGeKkDN35pFP+2LahbmHbW
vQYzosdIJtrfp6TQHJd0DsLTwJwCu5OdFkG0KkHuLdYbh7LcFuz1At7GRSljgrCR
EXzxOFxwc2gVM5C9Qed48dk9+BCRUota9Id/RfT+b+ibOrkBkERj6hMJsg939kHm
qFHUL90WN9rTnE6WOHkoMNI5cOZp2qbpNPe314aGMcQ5/Ul1WDawP2R0ngUikde5
wF5Naw6bOyt6j9qHJfuDkBinYrdAt0Cf/DdjJsf8Vk0dR5oOp8NPUye3sSzDsz5X
neYI15yElIgypPy/qn7M8aQ33IXSWmNMxfQ+bSnLwlWGV2MXpDpNrd4dYdVjs66R
axlcBSrIjonipXiehduGRZJuE+TrK12UC7/wzohJGTDTAoWn8RkJfS4fiPrRNEEt
z1dCPpfOMx49r+jatNbNdElog4OcOaYYvQod/UG6kIpzE6ioK3r5d23HVz8fyiXK
uvhvJ4hdm8SjfuozTn59jzmtYqKI1XaASZ/dohn3k6tTLuHqjsPCmlz9NRp2WtyU
iqTnuRjSrG7ZCCEknN/HaPkiNseKfrGxpZg3aqH7sIs1Msbm9Xglfyrzk66jMXGu
ZYkUNPf4GKqBY8D4POi1Dx+B5ISgq3kbJ2FiotZYpVskzPgq2GNXDvgBDNdCb2iE
KWp7bJg2bBHHwKqPPVqHNHuPhaILfFaFGLjayEJ9EtAwumHTr0uUH6UbwppbNJCa
Lfawxy6y/p/sLvKCs77l5lQ1mcQueAh6XOo5jt57Pqns5n8y9bzQeb1D5EcXOI0+
n/7ilZbu2qVON98uErBRU8os8Mvg+pMr4vF9A2iCVTvlr5FPvotNU1zyqKWfhn2K
87axBKJOwBXHUHDHr8x86ZqVkn0niud7xNV/s2NeMcU/RXTEajr8ocgX6RlBcsBS
Qht752UZOji/yE+Fxsq51NOCrxGfW7u9onGfdZx4+L5sNHOlRbdAttm5sq3aGcTx
98vDNf2/3ucEFThPLHx9ssjMW0+e/2YTUicTNF5yaKG3EiYCKfTKuKgZzWIzU0H0
aT8u538aw0JPYo9yOuZinOZxDiuz6tF8PTwC6cjiblAFXwsghgb0yZVzjtaFqGAN
snNV1Bdgue8KMSbvHVf9oM0UP+dsqD+YXJs+bVbDjGJJOO0NXT3X8I50Zo+f5DCP
RMOTQjl4AemwMtTraWkpvIkKuufp5tINyHFv8Tf35XWAx/6I8zL9P+As7xkrK7Ig
0V2HfpXyDQSazdDbBo9HQRthol/Ip/HjLwlxdJv03vl2d+lXR9oYE00+PTCKyb2Q
Rx2lrityGePbWh43OZznnJILWVOcdxPot1H1HJ5kA4oseFMq0voH1uk0ZSdIBXbf
Psp9qzZLiRX9ftHB1hgJoS67Tw05dt1p9UtlT5Ap9FOSiToqjnX/aclMRLbSSzm2
pZYXq08GyDIEVStdIWX3yD/09hFF6rW2L0ZnRwxTiM+DfSBtYMoW8Re7Pl7GF7ag
Lxq9PZUw6Zm9kdAiyWvHVrSMvF3g2uUl52eYdVuSuqywDIo6wSvRjpqOM/ZYcJB6
zYRRF05jgHCM1IpNWlM0xlqnNyo+AesqnYpH+ywnCHZ3lfjV5fRQ+Fm0TEG+fD8k
WAFoFV/iMcUOozEiqso6i8OVDt3cmb60Qt03ZfhJlU8232QvzbPcY6OlCDqjQJIi
6dleX7JjOGr+p/qHJ7MNYHwWvBznVHhotrALgqDI5vdfHtDXFGCmHyLe3tQE3irk
M1E3Bj0j2cd3FMXdScMUDWLeiWOyIjeMwU903sW4sCF3aGjPTSW0kO9zd2C8a7VD
KytNeKXovuMU2W1+AS3lbz/XXNAcztEr7PvHlo5sahB+IIJCQgRbJ0F44+o2o1VF
Bl0gRtNY7l/wH1klaB3vNSgscPS3uxUJmorzcdmTnu1XXiI9473Pg4auHspRQ5gS
fh+IHnWTLBLhj1NXdCUgs0rj9CsaBEsa5OPMobVOQ2bO/YFTI6H5tOSajrtmr1ls
PZTrVjHMC34w5E+faknc/8w/IJs9913EkEWS1P7LSqMkSdneQ0TF3HUPXmLcfi5s
47OxXtmD93lygLGuoVUiiqpAHAlITw6QMO0LHcFkZuYtPP3bd/eXbYKxCvRETC2Z
nUmSEJXRPNlJ67rTDGGx//asovo+S8+k5xrQcx6UWLzx3X6nlqiD/+zqtHDhD8GK
OmOE5cdXWSidaLBptBQYfg6t6of9kJJSQIgVDRBrydWWf9ecVOGOsxD6iyhGllJP
PhrfkBvRfzIZB0TuZ+fQtK1j1hp6YLK23pKTKFq97tewU/I2wXSnqq31sM4HREhd
CCCRZk0fyqCYIvv/y04cBM09QrX3a6jlhFvALLtTf+CpKqvff2OA51GnqJipmL/q
ITNkjeEbK3b6bT2UDd8uw5NCoPXHcNHaHXHIumprefANL//hwRG+J3Zr5J93HPj7
9X+tV5k3/+ZlgtJfJ0it6jU87qpqlA14jbLgN8Gq7VRXUncThQEntMnotyacvoAD
c1+5POx1BFHcrgTSGJaz7TXaeAgUGzQew9cxbKvBC+2U30zzQfKwCzIqBngrBrWO
xnpDdoExZZrt0nzACKci1Ck8rdvaA2zIGKoepKKyoW7OejWryW/K70iHJ85sbv9i
k5BrWe2JvLY26D++rPJOKw3aCdYkU5+hGg+Jjw+MceZCCa6PLCStVYx85WpzDMbU
RpfXfp9oE67IDPq0D2xDZfVbbWqKmpeAvkdOwCJ1mEJrWckcA5PzPTShg5QaAG6u
zwJWpXc82gApUsLJmBAYJoVoPtgiPjg7/s+JdaGlBWRJzV2S1cgQgBZu5Mgr4yDX
XHNyXYOVgQstLO8RKnMRb72W4oFs6bu7Ok8aeinkD0p1yZR7GC3cRBzOHOexO1JH
0leCrje/atJHA4BuPoPuORqpCCiwJjRIkm2ukEJSKja8tPyr5trzalrvmSOwL4+F
lIP/jO9Ef+W6ENtbkvvP8SgxykyRQGnz+FMfkhb3szWIMTiJVVIDBpJ4QjC/9gm6
kAwnHCPAbKOJ3YKUe1MidIl/eI439Ua/7X1oMtGPPgk3b5YwhBJySXNGXLBsDZzA
FNAdD8Q+pzqQgTicKak+GxMnuRK6vidqqWX6NiWo+dpcSF7jhTbIG4fnHUX3q80H
8KZ5YPS6aLMS/WFkEua6rGM3Akf14wbaKXqjvAYZOQf5uCQNn8+mXD8dOZmdA8D3
k7q1fugUA7J5dSqe/Sb8MziCZ4vcmvCcVV3EdEll1saNOWl/UbT1Tf8banCxFidm
2d9WkKEfudMNRPQE1HP5DPLwRHnoYuHYmOVkRvntyZzKfgqZxpOSLhujqVQfWotg
hKKX54jtByJGDy+cqyxrNHLFfGIPHkgr3Tw6I2Z3PdIeQZKH0UkkgGTuM1EjH7wR
50z7NjZ4Cm3BQVM22v7H3a51G+r4oAs6QW3T/0R+4zbWvc07Z8z2LjJgogqbscQ2
/7wxcIq/+fTj+2pIpnfbyKnMOiQasT4L2WXT4ubmDpNttT9/A4Mw+ebPpmWJ69m/
Y3M/jWRL5P9Fi1QA/sAAx9XAcgVsA4S0EBQCtgCm6+gdFfifJCaaiwCRHX4TfVtb
jZRa9omS5mxRvZ60J3/+vVq9cwCxlY8ChBoIXzadOopH2sqw7Dpl5I5havxRgrox
5VsJ/uCUlBdtjnYxflYntd8bJ7dYUAUY8Pwwy6sto1cXqL3kZThkPFJFOiYnhZt4
SnimmYe/BMzub4gTWKWcOoLHqt9y9vA95FiboV5vBPYDhubxrAJkK2GhMlqR2KKM
D1vEAdJn9iSR1eyulkT2A0WTPYghCzoogKVSBZwOPPU+4qeKJK9eivIJzrnFVXuC
kA2icND211wHYfX2GOBLrut7apuRhyic5D72TkUOit5e5s4PjGmnix1HBGKCmfaW
6lxx4du+rzMuyjfeZ1E/6OBMqh2EWDXhfSDaFR7pdms9iv6DWg2BBAP+uN7Yy+g+
CU6r58IeusbDxLcnNHp8tKsAHktTjp1/4lDlt5CaM9i8A+YVYo6rGYSmbk5hHpf/
4p5gwiacmcyelCZhkC5RwcXYFLJWFUY7fRzAm2wYXl3OnN+I4uoenuSCy+7gNoaK
mUGSk3Cp7MjntxqoX20svDkrGWlyxXljbyD4PyWRCNxGGKcC5n4s96YmrrII+mYX
J1mj6D7CN5rPZrTdI/5ULUgmh3digwnRcFiDSdDIzLHcTTLgkyRkJrd793OUvWNb
OSHBTb17/0qAhcQbVEtaPV9d6UNC4scimKSv7/f7nZe+o4t6Y0ndqnWsrRFYeAVx
JFHOfsD/EIYzNZSFZb0hYhnj1gmW+JnEcmg3xCxOR8KpZ0n1IECy2xpozwaH+LGc
IZGlnPNnAtmmQNLI7d1tlh0Gv/zFKV+ngmXR7za2D8woc3MurWz5yAMLm81R1UVl
kAsw4JMVkC7jvdE/Uq5cl2oXQpB8IwPVkFwCYKGkra+28cXlztL47HwlaMhjNJ9k
rjUG3Lw0d8rxYp/MICVa21Olm6ULSKh0HEeJlvjLOJHiMt1yMmWlPvBVBlMkbs5G
TBoXrlqsnneYTGEGQYEDN5A3Bxlde4gj5Lln0ZmOWxbaGVpRBcCHO3fs44wnE6J6
mmtxDgecfb+BKHf/xy9zhqSi+v3pO+CFju7O8JBjLN6H6ByT9ucx/W61fnzl44tX
QTTHyEjL6uV6xc4B/GBjPFZ1bgnXX91StJyTPebrnqDFyuQy2fuzeqLKGRzVdfu+
AG03wT4PCNR0K5634zvTDj8K9WKix30/NKeEn2j7mdbYUyLEbt0Czs7ypYJxPysC
Z/W7BoduQgsicJg3H2EXB1fHr6lWNarcDf0qhvIawPQ0GRNC0e3eetsJAy+I+m/e
+MjTUPcAIh/eTUe0EEmEYqGe/4Wfafq1HdL6P1++H7TXbs38lLZ3L26Juje2uWSW
BAtnszgcXs1ud520fbHAiFTQRUcdnLQSA3XWR3Y7AcZPqIVF7T1Px228lx5PoX46
Q++4cTuCy8vHPi13yatZexCZ3pGgwIFQTHiPjrNXE3XSUiwi83UIvzPhpypPD0zq
Uco0Kj4qFcap4cGCwdNs4trRJIdNR0wuQ4q4PINuqCetpftkjcxZkTjBncoiRqrg
yhhBNwP/B2mNDP7fQmuiMKJnd1TGoV9gwmeNtnG/piSxNrBk/F0SIbXhRlW4jpKa
iBceBk3YRxijgW0jSYISCrqXXHqmm6zqQclVOdZZh8kF4c6RVDZMt43RH/SSW70o
K+UUGdwIMfecQvEy87tTZolXtrXHJPzJ/Uk+qLT/0guv/OzHzmvcmzThTBCQ8Dh2
OdxI8nPXIAng5PI5olGh1rPU2YDp5e+cElmAt5TkC/6Mm3AYKxnSeE474PL+NBp9
PKiH0JMVAeHxtwMMQwf40cjmNv0hHNqYZthg2Y3zaEfm+08nFojcb4nlPILMUQIo
xC8cUKUV/OQLJz+0ZAs9pfv92qU/kqEm7jCijzF81rRMCXEF0sJcruV1/bJJAR5l
X/wfilhqtLyXr3y+OEA3ef1YTUidqW1ZagDsfAkBI3ELYYenN3o39PCGoqWbh0cB
zdo9XhzNd6VQdU1bslDLnIGUDm9k6ZfSzPJx+2miFzCBOTeJ/Os4oO9a60p+z/17
+7P1YoW8Hh/1CypV2tQRqzPgjq3r0U7xqMAe843L1kj56VE14w+TkOvPXUabSrSH
Ze1nGvyoy8jKt9knyOCxb6d8jofNARJLE1iP12sW6hRyxAC/ujiOM4azZvGvx52n
MsyHrpaQwoufaBbWms8TGPKN2ViPW6+aGbW4se6TyCOspSVlQEsjgp4KwxZ83Zhx
xhFDWgiQlW7aMh6iaF3+k9bIPDqE9/qzHjMnl+toQ9T5voSEzzVDonznmWEmde1+
QcLlrIWTTNLPH72eLdWmOyYdonwnmq+3S+wxewmbjH4KRZSWo682IomfGuvCDi6K
S88JGi9wCHxw6l6gnvKXSM0RDowvkeJqC7AEyrLR++b0qZvOgwJfrMUfBgORE/wu
125Zvpeps9RK0ZQ78GnEP+TzsNMM0TG2UaDhySFadP41fiYgsBQQBsQvU7DLOyBe
O0/NDZOSbYvFsZaHNl7zk8y2fxbdNAV9pHP5xda1u5x/qghs0mZ3p2fM9btVhQ1a
LGI1rjrdO3bExZ+wNh5PGnTAzCuxP/6liDKriJ6i0KRlhEN5naEa1gpx+SdZRMez
XzeUPIqPfW46LlWF4Mb3nGbS054epSzBV7BBP2yBOhw8xPuv8/6J0GfmSM9MIu+E
aOd85kx8IS1SbfXKcWVFYIbcihSRdyPsthPeGQl+xZNGhM2rz+dMhG/hP8J3Gkk4
81M0VKcYwo5z3WqYd2hU76P5HNFQHG9OLTLuVeEtf7BAz5jm0FPPgKZ1Mq6s+9bo
hRjhYoU94WH5yuHr+AoXbJr5u47G0d+GjCcCEFmonH/BQkCxisrRDBPS+7Qlu++8
UkX1411nYnNk0a7vEl6pbgbcJKRA6beE9zQbc27kL41NzZlnW3j4AQnivcsQRA0W
9srZS6ATGmflZYp6c4itbqHnN+d5ZDjoRXjy5OQiqXMXqb9kIqI+14NM+AUxV9Xv
ba/PHfQnY6e6O2FKkWHSUUHdSsGgUh7j6qxdBeNKo4DN0xHoV/JK5e2o7PCDNDwt
6DAY6qIaWrVCFZ9V/RR45reDHUTrrGT967aXO5Cd5pK5pYrzwGNYZ9Cn4z+MtpNH
FgY+GZOB9+wQ5zOjOcIElQZtrHfi4d4h0iL4zo/Iw1E3Ht/0Bg+5lw7b6KG09y0J
ovrvrFkIiInsr5f2eCKT3QLBUzEvQ/U/TRLKfPAF1EF6BAWFEzhcNq7AfGlnMTS/
Sf82EB/Dmo2aJ9eNqxOgrair3I3gMxs6eAMgVseTIVfEz31ZZS2ewKThDdU8Glqy
9Vy+fw8RIuBwc5tQWbTwtnhNQ6SgZJp5fpAtvbz+/vMHk8GJjnzUYI6VkRmD7czv
TCCZW7J7sBczNvrcISZexADqzrRWAk/t3Ylw4Xf1PONMglTUMHD/PryRosdfU/ha
LXDRqno10e7OO5N0pb4xn+vGl53O2z+8mGEdpkVVmIpt21wyRnRLXHbyzcTOoLCc
UdbZ9AcLFJrmKoNGIzD3yH1aVu4eyn1dBkcGh5juyqj6BXdRoxar3wsrZ/B1+1FA
j2gTWw3aL2Jn2j9uS9e2EHRpkn2g4rSz/1vuQZUi9ABy1QQVkxLcQKUfDev3EcH6
chZdtQYQkVn9pmEEMK7qapQogOsBN6FYbj/uSqjrBowal7RLADxdYYYNn1058OO6
6nG85WTrqztDDdOEVOKyBXauFvrbbCDwkO1/fjCWYfKXXOm+OR+ALy+q7pYuq7yY
kUkRMuyQg/8V7uG9K8/VLU1WENotRp/tWvpfiYxkkbkZcky20Dc7L6KajQZDnriy
0rkpwV5uDto2iqYg2QCQz+mb2KwfemekjS1Y1HKHYwOxQdo2bUt1f/8Fs9IX+pwc
iqB9SwLdhEd/fncSrl6e1koHcNuzxWskotg96nTD1UdaZOcC+C2uLhRoQ/ZwXOGF
WetnhcjYsMfofXPR8r92SwIMxP3C5q83RH8EwYttwToq1SSOC6oKYefVsnH6+taa
IlduSRmrGZN3S5XSPkpJ0rFfMfYm7W61GrGpYHqb9d8Q1+6awH20yuwYHlOpBibq
Yt5uYhsRuETB1c4s2tQeYEiFUcgfXz9lKBP6MvxX38gMwYikiuSm3RIxQzoBEkLw
L0ZtcKTO0Z5zduCi/WTKjQ5Yt69p9Ndsvq6Rnr911K73Cj0zc9cgMDRox4DY+mNB
LUAUj478ew33RbTGg7yNJ4caCPx97n8Y7Ccnk3yAge6oVjcD68uN/nN6xRyd24of
HzjxXmPqEj+yOwmN7f4xIxGRcB9to6nbZrHMMnENBsMncExjnDxpeC0h7asdK3Ef
8QoAmGiL4f+3jCuA2MHdFQ7DaEplsTBf1J8jQx/QsxvpUSiI2uLkz1xzjijwFodE
T6jesl8zNg5TNUrd2DAUSkvmKi9KLhM7I0beiGpHfTbQZIyA8n+hyjIji/t1XHNK
vxZKSZdiAG+nIbTg8Vf6RaxghEcHXr70QcFOtwWs6yxF4FS6vOIQqT2bln67EggI
Gh48tOAGlCoDSoPvGBiSxYgHAtSe+JprB8UWeq/chIGa7OceneJN/7ViBR8xPxlN
uLLCH6rB/ezNOwGM9NhnRviSNeLJ5FAC3ysrkcMOMrbcANhn0hwbyApXbUs8Rg1a
KHhRp5YO5pIxB/KVVmqGK4KdX8yNDtRXzv2+U4Of7NkRl8EzGd719UxVvBfvMmrx
McHBliVFapNeJ4f9g/kBW+AIkqfMVQc9yHmT5YBuq9uAX2XiV+RsybUFH4iJfItj
fEAxHSEhtoGNxi0H0RcAwFeNE0cXzgGMgBkLXL81SEVt+Jy8Mt/PGqXIRlSxwL7T
a0Wg/aB7TkqR/LYpHFEhbUmrB00/8F8cjSFfZvD2Ro80Wq3t/bmWZlGABGiwG9p3
L5jbaN0zC/sfpqNMp21cwy/yIfgGad40GzyTE2GXqLSiBCV6V7jCZTVOmgVUJYXp
QrQVAfUCTQofP6sV9xZDaOV8/RX8jJlpc8wZ9ZKQoGs/EpcoyHz6Bg/aaoN/TF8l
kOrfkQTZloNlOmkjW3eRhWdmE5oOFftkRIGFSPZlF7lAKjGi49UjKe0M8gtePPyV
87Y9LHxHo0nBqwIZljgBFuIAiDYLK+lGaeujaxoyLcxDnVh6bAdoRsam0Rcbexln
a4xpmvEA+62851/pZJYBwL3uKwGvL1t8VZlYzmwO2v5OzyyrC3oxpnz4pQbiA9tl
SOtM+nRk653T79Qq+Io69tug9C72qXzqOLZBQCEas7MjtTCl+mhlF1fCgEtIBz+y
D1WiddfXpIMKV2Ic/riicfYhdjAiCjjLmDyv10m+Ij4jwfOS1yWDk60dylilZsfp
JYeDfi1FL5fvHj7PlDHhSAv8p7l3VKuxNyI9a3dwyKVlyRHD0/EvBpivTfIVZLzK
Bo+Z98oaJgADjBlOHaCYoRjUqwPnWrxsXwNBh1RuyZe45x3Cyoufwc8onK6/Jp5f
n2ohvlqDrt9XDaxkLAvCBSOq+Zmpi5ebQmOtEUnAXEWH8+j5Lf1m2ntwzFM+irpC
6p578l/C2uett7zLDEvZrLc0yBAWwZ7AUmpe31dR1Trwt3G4Oqh5U2tJtbPpcxE0
4Y9ec/tfgtx2jGc//axAvRCvL2wgFs9Fre9Po/FDDT0xwpDEOQVVlMEuMPB1uDqG
GIdOza8xGqyho5Z9y+ldRj8jcQIocfbdSt2Lx7HCFyan7AEIcEmKYUbHjJHk1nS+
S4NSUA68uLymW/PEJhvgzW2+r/l6NicUwE21nB2nJUFLOK9VKAyKV4u8UV7XAtj+
VuyujcPhJV0aIqnsoWY8qZbPiDvnUpylL3+g71yileKgNy/Mep700tW2FWsA5ppH
TgPr2EvG/6BWo9YUdY96c32mhrwucdJ7EhXGjEZLYeJ0p1/NJLk2M7yi+ljzCYSA
nuURe9GKxTISGhzxilM0kVPA/7QF9otlijSU12671c05hvcyZjQ0+QGeZDERs8kN
tS8XVpejzmxV4qCoh+NwGVJMqS37NANSR5RZ9xE+/KIJj7sZ1A/Nvv5t9FfwQcpG
R+9sSU12LDsReqy+OZjvW8hEGhVKa2nbF4kwESuVWeRBYlHl323ktx9Ym8AUcvf9
JZSL73kaoLzERY465kpyxJmEmzRD1e7tmIaMk5yfknTOevhfGroxdw80xOOQmdb4
uuqzEuNXHSByiZGRPnVwG8V3UK07319gVOEAoiGbEY2SlXOOVMOKAPEzbDL71p+o
Y0Vl170X8P1d+QnUG2SvlZjaTNVLugYf0rjxM0wVD69TR81OIC2jTSkMOkHRTWgn
yLt1+4ki/9K0W3qT7gnFoLZzpxKepLZDlzM87ilqUmxXLAdziqinAVMZFFj9se7j
QDXGJd6BLtOtiniHT8dM7Us45u5dNlS/Xxi4e5WJ3yOP5tluwHrha59+Zsy0SqFm
F8aeEEUGYAKh26r9KTX4NMRWHZscMItiT7dXjrWmMi3Yr/CEzwGLpUiJ+kzCBart
FakuzzJuKrgHQPWcj1TUot6bR3/xycBrLqVVZRsCXSZvNpjyyvHlbhvrK53S9QEy
JC6KRy8UR1KQNGYiB0g4+u+wtn5uRo4uFJ4PaUonNmKeu7bG/anKzPytbM97EUrF
+tqw6F1jguSAyL62q5uzwcNe9moSb6XeG6UImd2rSNGt1oxcFPeENI/Xd57un21K
Y7iM40YN3BWlrCqbvwJoXHNQJVzhXByHr06WLY5UXypsjO5QsqraqchEIJMAQGNF
VRCKAMzXR+G7+p49zme3zL0BU1CpF+uIv6VKSRAfiPmq8T7T9FqmRcdWiHTS3RJA
/VVw+xaDOzUPGuBQBoJ12SdO9ptTz5HFCpO4tm4ZDdzbSTeHNPtdTfQkAhTb+dX9
g+1sTXIGfYqy37ltifSRCPmDBRx7EL5xDfj9R2Sy5ahCqHH41FApFjIsuLpXyite
K1/WInX2Ull0M9K1oMAMqB4Gk1OMHsRSpG/8ZT4rI3/MazaiAeSQQ6GuoUtn3kcP
aWeowPUAPBL7jC4c3Cc/0ZFcyjlUiD7l3zm+WCIidEhPzoIyZjggA8tVvqozPtDn
jt6MU2m1d9WuOaNJRkZbSU7N3m8GDa7jv8ETXTKPXED9HHNrEnh0MVbDvSsv+p+S
rgqnpG2CB3upF6isWOFleMPlZkpy2eUi2OvYl7tVCfWbKlL6G6idLAVlGzgqeLTq
CRdlkrlR5TljizBTUFlL+9/fnsPomcEhu8DKZah1SIlFzhrjldyxQmxLKaRV014c
obqr/YAHISoeRmTFI5626UaGx+wwmXfxCOtBilOI+ptiXN77hJ9Lfmt+jAPVBnSt
qNcv+aFda77k9HDgFPi9CMdmBi6v/XrMATPm4/68DzNgv3MFDVygxOhl5cIZIvGF
Ua/rq7eP6N24mmmiu6HATqThgSD6b4jz7pm6kBHlBH86bVs1viTuoJZf2tTWE2q1
/zwA6LxIu7Qmyt9YuKKJ9iQP4/Pf2PIqKbe6/dujeOgN+sTFODbL4BtxlbdctO0x
Dx0pS9SkUUZMrZ4eB3HnwyEGfVtvr9w/tcVQ9Ty4+hwYY3xvf2PZchcWahJWk30k
xbbDVREiv2YhhDAO5awb9jNg4UcnGzghEg/wgjw+DF1hI7z/Zu3opYDwsYaEC615
rQYAkktdFjzu77scMs2aAUrLytr+uJUkDoTPBqsbwEUQmrJb1aI1Cb3N6No2hjXN
Aqe1qCnzYObQ4f1gDmug9XC86TZ3E34+eKFBjIlVcPSBXKNbdHzB1vekW6YQ4a/v
+xprMWyCpdtrxKd04XDPIvQTI2dpVBSdxG8yHoidsgnW5nL7sUDPHDsB7XmWVhM0
SsFm/K1uzhdCGQEWJGHyPeeJcTlPDCVRbiIWJCoSi44geD+y/BUjx7AIqdsdFJ86
lzW+b3wLWTnfYrQzkdNqe+dGVDH4H4jJ5ImZUFy6rVd3wIYTYsreR85z2okmnJZT
6TbhBM18HfePuWogQ9vg5572MSJoUm0MNsrBTODzLsQTrVjats/T2XzGGc5HGWFX
SoDatz1NbugtvE7UC3L/3cKFtDzueo4V2nkDkiKxf1ioQ47De0SLKZEvuuGRGrcN
DCvM/d5aUVYPzBvl8D8f0g0PWEuNGvSUNULK2Grz8znDG5x72gNFIFJVg04RYauh
De+CHs/qPpF6z9Flx3/MgbMBzy92+8yW6HHoiRgMwTuG1CfUwfTjlMcPbaOPNrRS
KJWC4qRsHn6F6CvaJS/66RoNm7qLgUYxlxBMXWQ78o/8TvVBgGDQh0Sx8iA9L10S
8ekEsX3jWMaDrrLt4lBnhJFJrgr5t8RIVhzQqBoknH2heywrf9c5Y3fve5eLZULQ
74h+dMaZ2cgzVNPS0GXqRM+I3/zN4kZPHnbFsbOISOscmXst97AzA6Fd8AexlPf/
l8sbLpVmh+YOlSgG/ZD81sWgyz9VfGmmbUdO8xMISl5f7QIIuAuLb3GYH1co+T6F
41zQAnSLPsZy/RkG0QOWGtPsth4dDOuzIUZdIEuCbsBXeyDADGF+mV6Ck9QtBx6e
Sy9fxJszbLFmIw5d1jizBfc8nHjJ6WEdAK2R6UB9bFGrdA0OyrGjlGbAQRDuE2tb
CrJEKPP8hPMgTQq8dULPnnNutIlJCCc0f3DukHHmD0/lYd/86+0yQJGP93tWD3Vc
FjJ5BL9jc1UbYnhg4mR0AKDw/WpC/k53RjL3cmgWKrFi3yftOlxhZUOHS/WnbTg1
myN9eA383+EMSuePUpgrrpi8Aot9d9fEVUj5GW9IyhzddAA2git5SQvegs2mujsI
KqAAqkgWXX8SDVx2/NyU5TEl5eT9Ujtl1r4q5KdNHMkCZS0MbNfI6DNbFDFr/eID
dScf575xLpl1UZxmxpUYoYOnNivg8JSOxe72UahRiXwo/QzMbhvi/fY5J70Q69cH
o00fOafI+41q5M4zHDT00Ay/WmsyjeW4Gyij0KLeXpwCJ98JMZF4j1Y2+tEu1hRm
Xb0Zb1bdyhE9P8WuaGkbaK1HC7GX38WolcM1xrWE75KmwrI18EToyrjIzXc+YPcA
EHPygrYzHgErMePUZKS8HA70sd/f/LBODZ9QLP4ryP1oj1aWW7DvpzGC0YYJv5nw
Vr8W2IuldO8d5FZBw6e5/wvrXj5NcmqA6j8/tcYzEjKKuRRqXccUfNfoakKQQ/nk
9pbmWV6ds3yH0bOMMQHPOCeO5y7CalAgKEeOgFA45D+4Jc49ZmKwtP7WGdEDWcg8
qrFYvkzQdq8jaegwZH8UgbUF9GKe+ZsP3X9zZza7xfgLE6FbXcubPaPW7ajAcUQi
54AlzBo4G+7//NF7RgJuuZIYSIOR8VYKAn26/U3gMfQVska/UXS1Y8+ZcrVTnFtH
dmhI+3A+rUARUdqaosMuVGJnu7PIDkF3xEV9ITlcxJ15kOdJ2E7T9lleHQOoiAbT
1PK4O0Mmqx5NH/mBNmAe3RXmX7/vq528HDMQ0sIiV/kiwVVgNURTKR7gL17SXMqC
taLB+EXN0A37/eQYAO7sUjF14Xv6kim4M47L8BCtmOj8tCPWG0fTScMt3aT3YSsh
mdUqr2BMLlVoHpkPT4ol6Ukc8wurI2QpudQNdi4Ylq5h0AA+o3kG+8RtANKXt3JE
nD6NKygRnT4c7JK0D6Y6GVduRE+CUxyET+Sj5kDUkKB8MkocLCsu0Zi4wTIu+gXP
yM3rVTyR0lPEXTnmfmOvlbGAPlDnpxs9cwM0obGOqEa9qSpx/fnYjBtngLA8z988
goucyfDq3F5BcWyuQIHiYQ0nCcXO/M0YEwu66WNzDY4lJoKtGY1XIf2StZNrwdqz
9foDvcQok5Ar617JA359sirXIIpyYMFyM/r32Oi0wTp++mYuIaGptOIbEXLciIDo
wSRXx5R85FqyeDwNiBkB6X+40zwgFdgsGYddD7wEXpOHz3fUmnzw0XVdFQkvfHQw
6h52HlslAxsT0GWrX9YUhFY8XOUvth3BPPP80OPIuPHsAdjZ9KfXa9t8iPHPnzuw
NSwjfP/yuI7wrjMhZ4X/dHNJIKPtp44L/n1yvWh+fgDR1RX/L6s2vcrLjGgwAZIS
ZaqX/7C0Z53t5OdFI8WfqEgCMdbso0lB/lil+oMc05JnsFfB7DLwlMQSJc6F9lva
zYjmZXM6TzSKFy8bBHEnIIrVw1BIzu5t/oVgZc1iy6Ahy7mqB3lyjilSn8Skxi90
XWllDAtkPZ/zL0YP47G3uYeb4r7SFXk/yDsZW2XTtPg+RkacYD9m6E/L8D+bO2N4
kKlduUjpasjqR7FbR8Il/QJekGqMdoUyyaEBDgDkAb2KPrHiaRCHyvCbYwRTFOdM
+QmrYJ9msAYElfw9OsymjKW3xfeW9AKPsnrOwDw4gl6DZxHfFlKdebB2cinoNUzp
FCt0EjabS2pS8k5zMi3WJ0bVr4mr8/hWXe1QMHneVKawBG1tb7ZhG/zxPbFGP/jy
yJ/GtG08LNGZg3otO8J/6FwQODdlvIQ1eGFpJC/3JnsDapcwe5IctiyCFM+RSzeC
SsOx2nJTeuvR10811gxs+GExzwaQiw+SEmKAj6q7aO60/0WYwZQfCccoVOhSgHPq
OJc6W0QHvmPUsRlyxGWnD+ZK+FwBriQuwHK1v9Rp1FiMyGaQYLqP6POB6b1Sfsmi
mHx9kieoCqIIC2Y4f7c/GzOO33PyhU4zkxaILd7uXireLPgItXRFZ3d++Yl5VIO4
yoRt4EFUioszXHUXZTpsrvF3GD84oF1fUq7QprBMVqHKSv9wB1FIdrU5fVr6+fjc
VjBeZpOjqLrCd4mR9/tbHVS40tU3vAdqU/Kd2QfvNUF9ZOGo5Ieg03luxJjOp7yz
xe5KDtz04kQNpz1pPd+ygWTLqqlDZgEbBt7IiLG05oS6YQj8JPAGgulCHnffb+0L
GM/Hzv4y2vshK26xGpqtbK/wyP6H3COmKhKd/Cpxj/r+RT9KH3glUbTX248jH1pf
LBXP5JbycXyWJOAKthnbNjF+QQ0AAzNrXMqNX/v+tqLWicYN7xv4JtNeNeIG/55W
tMQZjn2DG8NL2GwFrxXb24SjCLfoafiniKbLmXQCxw7gr2sqVJRGv9tZcFdMCOKT
3iemQNi54GpQZfF63g8Yf137h5hJ9qOu2KK4yJjMzObMqpQTJ7mfWt0ybhlO/f1w
U30PxtxeeNu0Wvf9CjX4DFubOYVVhu9kITPbcdUyVm90oVVfsRludyWal1mEPKaO
WxWnByUtvpQ0sgf67u30w7DlKbVb7F3x6nyiHCLa8uP4dkw7ibneCH0MXgaaSGT9
iLMGNXCLBiTZUKeEltEDFpz6BFuCpGC5wXMrb5JRNDubTEvAQ+jz18SJT4xtgvOX
4E9k+I7xkN0i8J92+oZ3LeSByB21zapdAMugFqoTQ1o9f8FVApTrg/uFTVy5qj19
fuhUdKG6HdPxMO3/JjiRk1qb83U8qRwSP9smkelW2Ybzge7coe4/IFUwH9BVIXE9
HQliOhlGNK1BW9QvThuAclDlxbuQPc7nTe9ee6Ca9MCatWn+pALDcmkwlp0h3k6x
5F+Mh4CCnFlXbpQxZTcOdCqkm5Wa18/Y9u/U1puM9B83aGJ/uXyKnTegyknIvkAn
SxUK3H9sWstGftip38QjBw3N86mr3rSiN79otkNOQFt2oIyb/lxO0lCCulxgMk1O
55dLTJ/DgMYpc+GfCrcGy/QHltBYX4R/icycMBZyYlwEg58M6Ik+aFHBoFHqduAb
mJiiHO7TH/j3VqC4eiCfhI74alEJQ2Vexwx9oTIfTOIV9IY64JWNTNd8N2PdjWx8
e74EUQikNQQZbmEZjPa/vrd4nFM4VO49d2/EKIdRhiBBDx4R3T9mveSeqWmLHAXo
82peHn6gNua34EnYmQB/mYofYeVLPyAYIeMfPEGi+yE7GtMKznKIRveyhCwlpVWG
6G5yCG3O9fTzATLFWVsj8Sy7pAHZkTGyizi5d5duAJlIil3OLs4Eai4hOibNclTc
S8+ZGjJiofQ330pbnN6mEndYQ9Ayf0Kxs/9SeLSCtDHjCVSOZQaDqt1krb0tYQyH
xI5wkVs6VAF7nKEM/1gpxVnL8K6AXHDsRYQINIqZZTNuWKU7OqHeW/hehf5d4cFw
uVfR6RPiNDUWaWkq7WXT1Vc/XzkiEW5N9osf4vujht5S0XoF1KFgjioad6Jn9oKR
0FKf1/J0wJ36s0bUw60WceShb0Sb3lIDlso9uXIW9TxM2nQDXkAFTXQ9mJF9NNNK
GKXpo0eBG/4EODZdKbpBmfHKYDNiry38JwfzUo0TnE9LNr7LQ8qtxi217hflKafA
5Ob70tgccuAXKmvxFj4e3nSh4aOrk6Bil6d0ou6n+8DsKsQ9xUQ7a8MTMOcTAYbN
pCPqy99/Z96bYaPZVz2avcUhz+EmnL1VIpC3qiB+Ibd4mHlI9Sx6/aCu28jHhtWD
LBFDSq8B63X8mi8G7inW8rWWGrhJ35/19OxuAXVbwZbCa5WqwJzyeuDEUxivi5kV
W3ppZnJSwsmk0wW1Tz4gilKcArBq7SAluTWZh9V+MkG2X5FzOhJT5/faK3bU5epl
JJtH51TLIzb1y4J9JIigUz5Vwy1GjikWe6MknsNZIgbs/1CFJovX1JKSPUSwHi+C
MK9NjuBfiFqLRNdpwDvTRptVk8prEsVcuSwk8d4RvodRAml4bD4dXhOkj8i9h4k2
cDhPnV2gxdOnEF62ancBEmRsy7hhcGRqn7StMpClAH4LPUzC/+IFeFLCxt/5DWtY
qEwuYrXdl/Y89Ic5yLU3VgVIKJTrqac+obenVpRc3JQPyN1Nl/rot73poZGg5dMo
5Z7NESb45D4VFdAv7JYW94HOaRun7OpeioKyYZcGHRfBqZN2R0Gb09W4Yn2oQv3S
rYO17T/Z17wsm359c7oZ98W9JIFrkH73F09hbBePIPxbBEGu1A1kuGl390/OlqC0
Z1JkduU7is6XGzcZBt774rf3HbIvd/xkih9iMQGymb1NEkmxvOWoyMEVmB0QeE3V
Y84febXE2E5BFmbZm4+s3n2Sdvsci5U0KdRIljEq9RQQQabM2OJZSlUVeCMoyfJq
R2gPV9NFgpwWJ06elzCi3H3X765GMOvlZx1ch2CEWT7LV6UwKZchO4DU+FVWQjUT
FdY+O3ZLj+eVUsiFAYNLees3hJCOMhDFMde2B3X9m1TKH7+truVXsjriMVVRLoGB
esLQ+yKROgp/OhhlI6qkoJLnDNApn7xjw8e4BUj8zkNhrxNNLIyoQIX5fLdpLcs+
dnDp+tYYRv0R6xDL69D8c0l0ggp5Vnc4C9VVH76rFkG7Wl6xxgfxvHF/D9Zuv+qP
wSS2ViGz/x0lRUgZ1hYKpBTREo3ZNCsYwNTeoPGuzF7XXrLB+zle/ptJl3wL7nZ8
etRht+g4NTQaWC9iD1NcsFas7NVFG93c8RnM96n/EmHaPNLaqUq9mbYavv90pGB0
9Bc2l1G3YrjXbD62q2JYD0+J8J11u3nc0ZRXry3VNBK9kpKWohP6Ke/CoKi7f8t8
t8VoR5qsJqQzjdBcTFrjPkPvCdIAuyOiRqXeQ/rbjXU/BbbVB6BdEsAQ1zJpH2Jm
a0rVdEusSmFo7bAye7opePb4Dai38Cn314HaAS/nCx1UWuYOBFUUUdC/z+cnNPje
JDJ2aOCLaiXNsb12SGqCjOQYj3uk4vs/7j+cVim0O350ARaOFneq69sYYyVykUwV
xNfro8Y5N78aY1Ynmqn1IlaV1XCmGmpUJlmDgzFIGuKfW7RIWzr7OTTe0UeT0rQU
U97ih7XWyStHIMnLgSILsLXS5X8vjn2owQi5a/HY55ByE1LY2O8Ut2Hf8tWTMLQP
YvcK0gB7gq+Re7VKn94hm0Z0VWUWRm9Y+Cl9W1Oe8q3FSlIF9erM7nVpwjJ5R3xp
SVB4Ivj8o6eCx4ZAvnLPKl4X/hDpT9JCNWKEYyZjziSpn3z+gYP9rtmXcWdygzgx
BPbchzdlWHYS8GUXge2DUqDsq5ujQ/YLj3pK8aZORbbWRyF+oN00emDceEB/n3cD
Du1SmrL70Sbzk44l1TSoR6WpIZ+SHCGWUFP5B0GvgtK+QmqLXNtPonuWWOp+nE1w
ALiE332sNfM/7eK+0I7ioQhi3zS+UT2/P/O6sIjOPlUBcqbaBq+ivzgcdEwb/R+2
EtTjRTkuQUn9ht5ATP4TWAq6oJ/1d1BmVdbxYbCb6V6hpFNEsim3gx4GWbWRpvTo
1xTvkl5p2EW9BGR+I2lWsIOzljbdfLCULfqVN3Z0ryT5IjMe6F/SFHseNabLROGH
d38n+CeeRuEj/sjfVnPxku7sv2UeK7etWDjoGYZcLdQTcaXVzfyckPeT5/r94CVJ
W7zabL2fSVG+SXn2ilqKVgcvJ5hqX/ObRjMHCKlL92V/0q9OFNhDP9h5s3xgSy3z
hxhYl2Xj9gPoUhwsiqOQdqJJA5AjbbjdBraUsy6h3NoRz+SZvPd6zk7SzhX3DXjJ
eETEPtWIghDGuJLYY+lnSgreN99BELsyK0mEnVtpueiQl07WrVjGMIj5y/AAFNhz
sRHE5+vgZSKlmw71+xcucO94S+e56n++zOWoXJbx/MGbsG5vQb7ElyiZ1OKvViFq
Ppy+64YteV8WV56cvPJpzs25NPZgJuyysvS9uLJIFEPm59iy7mKD5ph+al8Xjxcp
kIiGVKiluVOkp036Iib3N+YtmxvwEHZBpNe+argRLiRmTMpuPNlGF+Xkro7Rv+CB
xZCra/es2VNAUkZ4QlQeE0vIjJpHMvMIC+3noRqu6IIfyFVWmDCQfKujiosUoj0c
3Qnkj4Tk/5rKQ1f/DfmacjQpDe5cfq2vEwsI5C9wiMxK9yX2lQFA89FFbLuwOTc5
GpD5Icg85dJXfEiX144KyJsMVK/9XQ4oWPsPw1YVv/nrRt73DsZ7UGElF5UxjI9B
/8j/MNA2FVsjQ6Wbq9X3QAnBjYGUvs1dZy5gcFEdxX/+1PK/oxqbzYZIIrHG0YFv
czNknt0RVDU7pOWGjgbR5WvsT1pxLtgbTnyZwOeoIPEvS0YJkAMY9R/x79+JdLj4
wkdSDzh46s9al+BlZSq6ilWlECr16gLUJao7LG0pjO7e4pLB20cI4IT1fgStW7/t
yHHlbZ/C0QU/O+dAHr6/d/p33EXeStT/iiPrgKuDI1HC0dh1xtmdtiQUlK/IJl3B
q4XU3vptYoAlh/tF9YRc/2w3UmzLpI4d1C00WETRP/lnCOhORQjrsp7noKoO/rVe
KBcaHh5JqlBayJgnM70d8WrYN7D17f89L3OIgApi2M60ucnk732Z02D6MfY0o8dw
fPW2ZkKTU91IjkRjrqLRcJtf47d3PFRRPSsjr4psKDVNIyq1XoSXTOLRBYLeVN1W
ccmhqsyWL2/NgGfGAoXezsHTZVqRDODJt2XtSjqrCZnrCJwfods+4iF3jGkjuGM0
fVD9sLUyS/YjibLnhMIqSAT+/XLtjx053YJlVdPT7na/TqoarKJtXry9sEGkqyEv
1kNz0ABXbN/ueSyleq472HC2MAn95KVNxzi4th7ztrSVR/N11q7qFkLj0DJRBnNF
EFeeMAt/ZaOcjYov/70F9YR6LGIXpfPhtsSoBsVlpYAa8yeuphWgYuHyvZWupp1n
rQeclxX4UtGormY3fJKi3T3vmBCDeZJsqm+H1z46ZF2JVVUgsErr9L4Fl162qEz0
r8hGLNgnk1E4DZdLn+U+vtnPjWfb5SgXqIDnFebFMawc+NiuJTSqFedFXl1HB3jT
6GWMDwi2BE+8HYte0cTlRZE+fFFcyNTVyhk10tSlIBad/zTXKUsZ1F4dWBATBqyY
ynC7TeruFEfCOKZX0pPVA0JA5tpbEaNkKBtRtjhFQizdtDuNJNe+8pIbAEqqY3Zr
6J6RbdgsBkXRT9J4yVq9QQpwvHr7owWYRPbQCNknr89Q2ia9eH5vrim5SOZoimDs
0+RhOFrG2mGOZQvAyGpXcSfzn/+28SGTQldPQnqgjEW7TA1YFeesIQAdbtjbMDWu
btvEiL9piQym2a60vmfWEe79M6yn9W392NFPXQIeHqhA5KyZ87iZo02yKB6CQfxb
lWCkpl0jBGOGK1virO2KT1JUO8z4a4/pasiiTgeyD9v0nvY9UxaYWEE6dwlW+gje
AtssLAwitQUAUgLvL3fd4JJ6QdgM2JFSG6doDafVv3Jussk0f55Omatfu3sXIN0t
YmfG/v/B7FxP0V6sfi38ctZZxaLsUBsUTPGIkXE5nEsjtMOQXDAXGrlkqLlVRGTM
DAD8hkV5S5yTe9AduUmsKfjT6Mw/ckxx/WfpYOCayYH1VL5o9524MyMa/Zd7taWb
//JHNsUWUP0rXXFVtUllNs9Xy8T9rKro7dnPij7FYRqPF73TV80U9vYRNfERMjd+
lnwaVYFhEV+DjLHXlruZbZaOWfU+HOoDm6ryuhqdYrklfKWl7z86LJVt942orpGk
uRvuYzHpiacxQAtT/wnEp7YiTFVcF4UOOFNmoJCHubJankrPJp5nQ5kFfVAi5vX6
8D44T7btgysJfZy9Z41qQo5S6NkeqnYOJfwlc5RJ//k5KlWwqxz44RIgE0rMP3/M
oevEUgx09nASnm7zhp4/QOqxclSnyDmobQNbjS4T8SXoZL2SHeSVK8OmcIrIQxTX
2Tfayi+yVO+NTUUkRWspklUsZ6kKPZj82eTpC1tie2a+yknvEUVPkCPP4lB6pdxu
qEhrbqulqjPPCwg/0XHzoWNOPIFEa5xuW91nGHsaZEVEqkxRbWBdO0w9P2rbDSI4
acPRyYsleAJEsOZ+LmwBdRX7fQtLHI2UG1ptdhrTqvduwyFFSCHhRN0ug7JRE0XT
CYS+HIHAaL5WJhktm/oqzOhe3fNc3YfSayhfw0LIZ6IyT56KYWkwcKCKgXPqG6HA
7fO4XAizBieadEa7cPw7JrZ++3gCZsaoiyvOULRUNaYoG6oAQB4Gzjd+q8pR+va6
tzFwfUYf2vmf6DB4dv/lzwmApuciFFS2pzHFU12jDH1PFmblnloRArxi7onnLkdS
gjPBwcs9qCamniTn07KkfHjAmCwKIQqQKTEJCEhgmjVIjANDZXtaCJUCsFx8sXTo
bY5mTrgHeeRn+kKxPTN2/JwE1BDWMjJFi+dEmhUyP8SBmKN/oOCV7q6BPnNPmBUI
AfH36UKSgj2JWxnpl6wF68okiVObIBXwCYWv14+SsxCIwskumXPC+dffAQCb1a7S
gfQC4LzZXnAXn5aeD9TfsXxze4v+c+tdSZG+K2uY/RlxxrU18a79VppPkiIRoUFK
XwDrbx6uVBfMQjHqGIeSih13TclrvZNfrmqaFTo9q1A0bFDh81/SN6NOk30T1BJp
Oz81UIbNxDCsHfcyor2UpmBLN3LPqDBTYNoFkPjd9DfHkvR6pHalmd3DY5VlNzKZ
BqH/fES7lexV6odUOqH7ULuMY//hPbbR+dI8sbMdhQWLVYubPAUqV/PFRyjTPTfo
hsdD3P1PsLvyFUBm+XA86OG6qJEdLtWQXutDXp/KopyYXR8tQaoRWV6xWGOyN1Ye
aDi6AQYVvc4r/qgx7RMvsjzeVfCx9TzvFIMYm9waRyXKOs4tHBQTH0w4oS/DrMqX
NHD0WHcl+aAqGzr98PVQXMSJGa9UhQcLDgNS5f1/LiIaz5QWkUQ2OPNETDfzhVfa
AIHSRVcFkz/cF+xMoQy1Bp6hISGobiySJDuB83htHQszOoxkmfZ68VvTaOx871ea
FkySsB0zlbu/idUIDE+KI3X5DpO1PHuiYnay+pUPCLnAEwFFirrqCkYXPuzjIzPh
kwmVfZuSWN1v8ABwrYPpts4juKK1AeogCPbshfViRkoA2qtBzoKPa0tVHUgfhACd
Fsr6hczX+Cu+1MO4YTMwS6yzw4MHXEpFR4meH8AeSBmQNcb8hkFCC2EqlJyJKjff
3sL3Eud9Mkly7MQhidOhAg05+9+qOxqIcla7fHqv95vKrN15docR1PsSoL5HcK4B
lBwN4xdcblW30Sw5odm9Ayi6bddJ6dzZk2f+bfiTM+JuIX2pJ30hfRDjDnz8yn6W
UUEprTPZ1I44u78WxjMKfSFmUtkpzz1YdEhtlG76af19Di8Uz0PdpOTIPQzhIoOt
19dvasEOJ65YishAr5aZXgLMxAzGJ+557GnBla/zfc6q6JmsAwZj5HTpDgTFHmwp
qF06idNVgeKH3XoaoIFVgKYvUfP8FNAl62QA3mMRsGzBVuCXGt/kzJEug2Z7BBuy
+uZoUclV5wKWPo0kvkKzBLhQTTF6uyEKot6dB5cDAa7DheGP4+yhR4Q45bJbtKdD
iP4wo6tnXQiuYJCKJmPj95B3q4zsQ2EqAbwyJSvT9FjtorBWP3ufX5kDPf/OER0d
lb+aWT375gibQ+MkQW5JTbJwYpl3TezkT9CmfOMDLSQBPmtyjd/h1wCrHKWCWjvO
8A43ePf2Ku9/+a9pIwIei7VW2GX/vjuoB+nPCnH8aVA6BjRgHGzfRb1XaWTw4dXh
Q1gWpn4+16jVxe0XOnVfa+SaAsY97HRkGCzIZVUi7wXzDWjfw1MXqvborIgYb7aW
1POgl5d+g2d0oK1fe9CiC8G/EmpKeBTIRw+KV4bTrVpH9VFSI8A8wjkqnKwA4xKC
8n0WHcIg5y4BYE+2Zli2DzZFE6eK8XoYU5mNdBuTerIuCthgarNtDo3n+6Vmf55s
8b7W8jJpl6CDz+zuhHfh6F6B6UG0FZA0qKd8Onlsvg/yKC2lm1vJb/jZPy6z4lHF
3MqLHvQr+3Ar3FSZ2lqu1JpEorjNjkNdEnd4tf4et6BJ8Z3NpH3yv0e83O4F4iBl
aYwVsaJNl2oqtlUqZRhM+D26wOmfkiK6+78V4kPWRpfsLRARIwsPxIa1BqeGddIj
WGgwu5HA9WRFZUbbU9qZf0sMKdiEQeVcRAyG1w3Swgy4hu8tPiKQZgO4Qkt1wvVP
XoFqtOJgYhHvRrqkqOJ7fPwU0q2UH595GakHIdzJ61b67bpR2t0/k040w3+/2G0Z
xRyByFZWP+FgO9LAVJu0atwn66ttie0Xs4u/pS0+9T0LyU335UNe3isn70bUVh9O
LPprtCvdjlHWoa/LC6MBmYUJIYB1YIfdAOXvkkLFB/ZGTmeVHLHVUn++8kaUFGWV
/fOE8c8fmx9Mx9+itGsAK13PzWZprXCg4a/BiL1HoHNLz8mhi+yrbFIANKe8Cmg3
HEO5WzGlEhwGzpUV9SMJaLc5AgQBaKO3Jc36CdKvAZhBIukcXrRd8OAMJZ4z8m4+
KPr3RwQq3N4pOdDvLAfiQqJfYhwl8mTPTpQTQLw4siiQrsm+9q9N1Ledu3UbDvlv
hLH2Up0lBnJmcaFrY1rdJ+G9hIPaS+jVCT4fB9JKjj7E+QlcbPBnCbHL0MKatCC4
15BM49WKxt3C87Nd+NLyWqSYIDKzkWvMOt4UTdntVBHyV20Lw032Ic5n3xICPAoP
gFRtISdC2CPs+tqgrzDjeLfBurBtpI4KOtVcOjbdHd+4/T0VR6AwEZuzdhBMIkUQ
RPnFzJaLOoAJNpCC14xsZIvKujtottiuUQE6wVpWuPFQ9fzvFQ08+q1jneUQbzq0
aBKCaJWy4LaZ6P7snD96N0GbSOjoiM9kA7IAGSvfp0yC9g+WJDMusAR6rZWj6FA/
Q+WKzbfvjCJw1tj+Vcsxacheb8ioll3NlqxKgnH8yiQq5USTpo84kLTECg6faFg8
sNus9y5a/YXTDEGxE0RF5bjC5gOBeGUpQXDe4HsxVRuhRfYTf8LHwIjQvGMtXCrH
Nx5XOxET8aLAEGjRZiotQmYaus9EeQq2J/mV/jeBkfBAyv7T/if9bRZXaKWibsLH
wrJGNaL26x5E3XP3vRHPfWi9+SXqxxmEnNgxm7AB89sMHkFhiqInAE3W5ghEP3hW
vkmdIqnaHPAvfaxTO012MyCP98qKjXMoMT0gUsztvn5yk29ppJgwiwo0/xD/RVvY
CniVpMzSsm9F4mtiSThQCJ7urOQxHZ78j/Gzjtmi5+KmaMhvErECdGZ6mADyp/SQ
4Fc0NwwR+X/zpO/sQfBbfbRy015DqiAWwT84D0o5GJ7SOOmeH7GUGOVDSAQbQkrk
v5M7O0k+6JCcKOAkjfnCA4kj6AxqSaQ1tpUmDUYMVjRxhtS8DY/ITWLkFXjJ3cSG
dzYlk2nCFi2+rMrK7DPIag9b/AtQbygAeiMYsE1TaumUq4nRJnF1gsfudQ4T37NV
mXCQef7sD90WXCtta6ySyUheNri596/3uMF1Ig6eW8qnSNzaXK7Q0ELMLgGt/Vfs
itNEGnNjE0DjsN6zhwhHtJ94G5IfqPRFwXWMypxIWOtx7KVB7EGg1b92IjGwD/iW
LmV0T8+0ojAKRb7OUHzAjoLiTjKfYc5x3x6svHtqdpx3eWHvNJtjm/z/iDVfxHO/
3rLuI2ONEOFGxw1JyQWpajirs0NQN+04476oQPZQ5tJC06M/TOE9pgJJYhCbsw5V
A+BsTyzrHug6H9uoyF4nXvmDklm+LVRSibIqztgAQF0qfO5s1Pc6gXfsi+yZ6e6Y
k6WaL+cbU4JuMS8OrY2twNY9HniA9O/XD02SYeXB48bY+9j1SVw60lq6TKzbAKKz
M+NK5Ji1DrJLNpVXWFpV8b5EPSDdYjzooBwIQenAjXrwQRYkWcj5HSUItiwPuQcF
ZBoFJYlGUrAr6b9+z6UwmjcVVNvEo4ZijmF/ht2Po60X2D+k0MkXjxHjdNNRRfp7
V2Hzh2eW8fO39g2JIdlQe9lyuHYRMKbCq5OTgdYdhYro4of9uSqDQ51QebtibIbU
7z/jUxJrR78677hu5Mv5Gkb+Bkz/5DDb0PtTtKoh5C9OJAX7ji791nzSFPU9esoG
vAPuWEoJMeocM0Gn3Jc8F0mClUSOL1U0JghKWCvO4unAPm3V2VS9OMB/mia6vVSH
0qbCVfI1YHoraW+afFxSqnBNnu/ShtW+UE0n1ubg5PobZC0yYrgZoXS1Vb1+xbJ/
REFr36K9KO9613fprMZbVe5s7d0ziZBEerzS4PaxT5aFYdfB5BC4K/oousl4xQ2V
RToyVhrp3wMTWPvEQur36ylHR+9RGf/uExaPu360cWDUxEiQVvRHtQX/UMg6jXiU
9I5Fd5wVxe1NFrEf0jV7J9HVrevfCAsV3okBdXNs+LBvyOFG6uFwwzV0SHLNHDf2
xcqaBvUmIzicHs0B7Nq5rnYyi8VMgcnvK1Wgb/mZc+FNSkYFB7Cc/MnRyAdcgIgw
jnpXMNjz6fc5ZSLOtVh9EQIPiVR3ubd8T1kpVGja7prNDoJHyJheNhKLgzlpSGWV
9BnBFMtAViEUBSBOKc/PzEZBOe6xBke5s0USbvYBRNSUdlbDQXmLZUirxMWIHzOV
qliKIndhUp1x1QcoVZf3zOzGsruvI7ZViJBwuNthauqxhDQxX6mmXsHPhG4swIpu
+lIG2NXXPlqSNJrYOHeOp6dAbFm5u1DrI1/Y9DpBLD6XegOHK4T9xtbfjRGdX1j9
GZjKjVdnLtzrAyJO1Yb9XNwAreHkyGTL1ffbKcSYCGdmJgGXJnM8NcIhoE47Cu7l
UNjSD4WwwsBFJrrjrTrCIBXJU+eLgAkfY5NkkIQsPHo8ImwPdbpQ4z6YdCE++O8v
1u0imClD5gI9N6wC+EsCWEMzzas8gx87eKKgCYjbheck3ugSZ6ks1hD5OzDWdjcK
3+yrmHTEl8ByP3qpW6XhTKOY2TYQEuc0shf17sk4kHzvRZl6kHisvS/Cxw2FQqde
3u4Ia/GVh+hjzgV5mK+jEI8EbG/VoacbVOLQWEMbRji2ANQRmi8m1NUC+dth/I/I
z1J4Er/HTUBfeJSMz6sAngplTgmdUeR9Jj/XlUmr0S+hGsS8ZkX17EOJc7Qbxu1u
N/pX59thAX94Ea9glpPV/5oyCU5OZEfw97JosIsGsoByKgJUxAtWnZcyCcur3xtg
e8rKLgXD/U8scbqavGOFbUqt4EVlfvtDHro+MiJZqBccwOdRxnlLpU9uEvK4OFzW
uc9p8QG0lt7cn7FUCI/pMDTczbR2rUzKvY+8Q8CViFoGjWKmPSz+IrOCZsKDY/HI
6sZnt4GvTHn5LcJOc6VV/AgJgeUVLtN+351h0yOcRPmo1PP6lIoKnIdEPvzN/fwl
kF2VSeUY0KfpGMx/gqCx9QsYbF5Mge5Jc9W7J6S0ovRu7XLK6ovxVTs8WyycPS4x
JTXCM9vH+6+z5jmmeHs6NkH5l42A3TG46SVtaX12jsGGFRqE7KJEYDcvK5sww4Gw
TzYDQTmw3JxkPLZMWCy1Bi2kVKES0vm1WPKJCwMDSGaZ3gch32Xtya4/nwIUhUAO
J30rNfuTDDK6rjNyhq/3Xw8UDj2CimbqkRjt+nhRH8hxYdzWzLmwqvSqG8bh+I5P
80EOS+cfcQCa0Txwr5QjM82oZWrjRcRk1/BQNflSv+gGneS23pKetjkn4gudrZUb
eddF2rPUcHOUjPxl/AZcYpbaNgcMhLBx0bFUYkGx7Psho/5zEOKPoOWcPmhWw4gl
+NZSqT30NQaLLJJ171ClXSEZMHPUvqosor8S4zjSv4P+TSufOURvMCvgtxlEWEqt
XRkLS8+4UXXCOrxq16z1K5FhWjp6nk0q4I0dvDInNsqVPvFM5r9Fl8ll8Sx8kg+4
YJctOWsuc7SLd7CUuEUB/FkCmFy8O1SjaQacj8nz9c3pDzGmIMTdIONAg/sI/Njm
dqAybgqrID4NTI7e8UJJG7rN120/qHiolzaIE+QCvH45xfW/rK9DCc8piTLF/w5M
3GYrZbiA+JGtc7/VdfTTEjdQsO5PAxAOMc7MhxNRgsA56UgDDRyQRTSUOBxqZm8t
P5y+Wj3haCMmFR7lU5EyiDBax1G0W2x9GumVBISws3jxI/PEsEE5+smpZgwXbyfR
8tXKsuoOQFbKP/+U7PhML+ygxt2pasYkoFAZV5izg61V8z7lkB4Nlh+dDF83Z1OA
AnUT1njApuszViny+Qw9gZ94ekBZLBAXODiDknpRbR9LoQ2qrRMS2U1LaynC/LJI
TjsI8e3siFRBuqkIVxWJ5gLm3TNNPyky2kbWFbnUZJMV1wVzNRemIyHbk+USpdxw
PZoLZJzF41UFcXZqy82yaMN+HrISYcGcvZJWT4QCg+97YhPkNvc2iYkAQkyUUSj6
N8hThLXCJnxLOQoCk2uDJ+jVWNnjY26DbhMVi7yTPbpRM6M2IqLWokEmEupYF160
+Pch22/KMisqw9vDzpIgUafvOMguinYeHx7fQm2V4Ne0yELxQceYtCyqEW1SwYLn
eGWTcn6qq/lZmM8Ucj+lXPM/+SnO9V1viMrgilnRQyLjS0fXzDbVjWXIw5dByZPR
J1JmGm5kizbxjSQefphuMNdiSo3ntf8qjeqmIL6W5iy2wU2bW3U4EBYlFlXFbPB+
JT3g4dCBjuFj0kEMK7fzcu0RK4cJno0/rT8nX1rcLs/L53mY6uflnfda8EqjtAMv
eVzWK2nVMXt5iMetA8x8eECZHJGbGD/PeFZBZxpaC4XzAZQ2uIYlcRBmTQZ9sCPE
d+5XIFd6ivZzOm97rxdA3tcw7Th3YFDTH0pGgGcwSD3D5Ja95hI7Q+OsRvKAOYuv
iD9NH2w630FY9eiXIIBirPtAWrplIwXDyiagLMfRURugEI6hOavS3F3X6CL8JQE+
iJ1j0eAHs9uJ+YjSsr+D+8fHwERhyBAVaQSUHQrf5397MoKOxF8MQqbUDNpD1dAW
06xSJ/56hId6FGvTx7i9Pbr/9TdoBIzucDTaEoY7w4ZVsDrJs6oerBxfDm2gaWhz
8CqjwFSbU2ubD713gpDXmUfH+n2nDx/eJwnuWPwg1/QRN3AgTWXsIBLCPO/hp0Fx
W1Szrn/efll0Zzj/azmlh0Je+Iz9aSkohN0VTjG4pB1yO0h/jTtuRrku6Pjnkpq4
I4CW2yDJ2W+IFvfsS6MeTgZTGdLGOpvBvoHJR/swSPVd9GIwiff2TUPejGpmkIqj
57nv1EvFXFzzOjhFGwCyI8or+KKpuInvrGcmdzrqHAvU1LbbmliuRu4VUjFP+PpC
D63gUpedQdlocSUFk6mU7D/wHpw0F2FGCklHIe4wdr4YFpKZ0YAI2LuvQIDd5bUG
MGOCsOHQzWKzNcBw9UdJgdoT5QS6J8bZaRopJAWIFn5lt2hAGp+X+JJMKqbN+cTT
vjFek7ktQvOjUvcl66eW74BiXdJHvEP+eixmoZbUD9MLvGeUoVJn3o7FN/zjaD22
XW4jcOr1nyvxfhnLC4LQ1og5M28AfHFtf1NJ6hkw+iA+JydOlqg1Bdzd2GAPFQVQ
KBMY6U7PFJjAXtUT6P4pZC/JocOXJ1Ak4XI2iI/2vBG0PE7IjN26JiWoRSaGBueC
QQpk/4WL/zuUmrNcaezFIAst1SlvZtsjZGYq7c9w/P5O5K7z3iLAuK3P2oRtyzjJ
GoayogTx6mc+ZAWZbPf81OBzL/BAgGB0vlzkB8X8eS+kFuZZXir2UZhjft2LtoU5
SKcN72sEyXtk0YRK/uXyoVKTrRWB0ylx1P0eow9wV7w77ZNGCRF9UD0owDgY8a9m
VjmiHwElIUnDhJdyHiD/c6Z9md/guRKlXP6kiusaMfcLSrvg7kMhNRbUK5+3aQe2
i85UhGIkyEAU+a/Ju6SmHtxCpSrHxhGD9GNkWDmE2XSERUFVzpVQmhsdqvsUdN93
xE892ktw9j+BfpWg10q3Dv7OyETHjTFWBldadu9gjEc3szDIqzPNmDKYWxKHHPFN
/97P0/5/iniTy5j9gKxs+u2DBLzfD3adwhphujSQfuwPqErQbTotS5sa6I55+jR8
vqs4KyNwNrxEddBqGbdP4B37OKfDwoVqKl4bbKIoxcrd4kOu4CHIGkL5YFpj2ge1
rUSfBb/wje6RFYa9YFpnXYuES4G8ycTM+5h1XFlVV714Bd+cFjhw7PxCdcOLWVjy
A5ju8q3+V08dMIZdrYwUjgHZsZctIiSRtrd0GUa5EuF8f+1XkgKq391P4X04R1xA
CDjakimLDyVa07GkyojtrhvW3SNitnJXX59fZUMWTTppwroNScDveNgVpB69REGG
NSOcYDa/i4vk3rPlGKSJIAmLIEjs7lEpOpCNUHfqi3o2CrmWbEk/ZP1rDmQfSxDa
167zshP9PUq5+QcFPfGhyxEckGdytTKD9ehknP38R6AfV1QKPI5XVx8oqEzk80xc
+KnuA/btcmkHId68zA/wspOwXFaI1NfV1dfY5K0kJyd/06Iff+q5y6VWGpSmbNrf
9QwuIP4Ot1SxbS88IhFEq9pCYiJzFgrCU2yTWDxvD+dEr4+uxY+M5DkeqzD0ijBw
IOiJoLb47Nz2uYHzOwrY1q/Zs7bYOG8R+aF+YFMGIqkSuqC0z9YYIevmaaGse/Ht
TK/ot4RvDYqOOKPAkFB/Fj7vjnaSr4Dwy3qC+hdITJeJQspVOLTNT4q/rzbDSFTV
GAgwIVJynYIHuutSVx9ofDt9Yh6mgRHyRstd5lQ+Y6VNdeIKv56wYaSrzxE4B/R4
VtmDX5FKymnLy/0qGabU4gJLLvbS/yXUYEKqfRb83A8rd3M1azp+/VyVWp+1bE4D
zOpYwa5IA4yx6MZZ45S8akBZhz1EyUCNwHUCRQrGTp6v8zIpbUKCW87QQPcUXZOl
H5DGbPJwSJIo2Sel4vBoBc1sH7r7sYLZqs2Q/OSgVYNw9hg9zcYZ2RYPvyfxihJd
/0rIarmhhn8N4Qo1PGF+y1xszfQXVoWvh7DgeV2TXJlLxqyxUHbXAdlz2l+iO2/L
BQcgWOzc07e/yYTCoNPQNttpPdd334Oyw76fiuFsyb3Wt9Ztg1j9nD9F36hTV1Cr
10s49ptdyUZ/X0c9Bvr3vc44PRXpF/RlAhTBBzI4LcvYjQU/XDhGBFzpvwoc8Osa
FWcCNR34NKc675OCHAVJb0S9ZmO+B6zBnB7WMTNDyGuI1y0lagTl6Jhuvu66FFpd
BG3NqPy7R+ZPL0MtpbMHINo+Y1V1ukO90sVqMqcaOHDQiCNVrDJT+4jbeyf54Fz6
B/xzCr8QwEsjOQqIqW+N7HKTYSnVLyRGTo5jz+87vTdFRzJWAnL0C3zFQ960NYwp
YXScM0Yb80sTn3Sa2ofGr61E5Nn8T5INJjhv+2r+VCziQyJio0q7XkIw1EZO12W/
gA7hp3e1TQEry69UujCeKFsa4Iw1Z4MliKoYyg9DPhkn2okqPd320yD5DDUie4pV
YmlLV2FYG1sv2EE7lLpv3GDez12Wo/cbIgscNJcRFb2nK8bYJD41XgoUV5L58X9w
fJpHjHHC9fUpKvVWPmvnYsPecuiwVCtQPLEWn8ZR5igsSwM3u3O7q0lAEzmGPJVw
6VfND3qoPHtpeg9yCjObIQOXldmTE9ftuMpaCcRV1qhCTstdjzpXC3kf91ds21yk
GswVlRbBnraMaslbPdvGNPfdcdfHIS0uuewc6/Ub2xmqRoqumUhGeY0ARv6L51R6
hOojQPlMHbTMm6STag1JiGjfZ62aYqlX55S5zEMSbxTTeUX4gz28ndg2IC6OTOhY
ms/H/KsS7ud8pUhoYMVv3Vt9k/D0nxUXf/tuZmDpnm9+LzhMsjATIpGcVBy0WLLN
OzIUt6XNdMyv0s0vjHnp/1SRB9WzjF2kHfylyvyz8A8YcfZbUTicNZmIGwuVO25A
Jc4kacgmR9hjKGSqaT8UXCs3HBWAxSyGy1oTBXY8Hc5JpdOwbew6K3xvDVV5TsKL
sKVcjszrLTpLcjIwhLU1hthsTIIg3PhZn9arT00wsWGb8+SZeioCC1SEqcY4/ec6
SBzaBbo+LsbItkGa3uIIDO8mUm31Fla4arGdDzYLFYyv4j95LtxqJbqdzicXxd89
mTIZu3JV6GlXXRV33qIBsrmyZevkpbra15gy9AMRk5nMXJSJly335zbQ0PB4CICv
rVUYOINDxbkPYuxXYOI+sGDS93HIa7tnTQ/WpRwOMuDiU73OeFXg8XWiPaGoEZo/
vWRlscNlIWo18gX2AiifeAB8g/z7F3IeYlp1e4nilx1dL5cz8tvxL8tIE9IoCagv
yIeV3qfQvP0cwUbq7mYeB2/A36GhvDD+ZPVmkW6tQ41WRsv/YXcUa0noMqIMvuyJ
7pWarXoQLKkM3y+vSfFSVvfdXcipO/UbXtPFl9xJKjo1ofBfwsGK2AanRTQd9Fmj
a/1H/29aGKeF/BgQna9bEGWk9rzbC8i5Wd6ZIY0vVzZoXGR/QIV1eBxnbiaTvdXo
2lhvIY8HtQkeDRPLh1Yv8dsUka7KBhTEuwEEqYLodKRBdmIV2GQDWaV71Fy9QCWA
n2HEllaelFovtWjIrkVKDeXfuJBNf4DikBbjLqDP1GyyxXmcCTwOj6ElyHRgO3MU
bPlAZNCFk/KLEgzlhH76u8KUT7+cOP//af3muLi+NOPgRF644WgpnC432dAeKnPQ
SnuRvY/4sTLTnXq+EJh5pQHWB5ks0ge/cAfCtrXqvd2DsVvRchAlVK2WTlkkV66g
4equ3qW/QJERNADXBvAXQg5eWB1UAPv4o42logoxC1+srczal41S+1ZBgOch7rFx
THLWMLVEf0B54J7flopzIDowqPs2/i2UAcLUsd/yuDKbJ8VGCYWK3Hrrkb7rEDTB
EujkpBuX9wOwhufJdEjG5jmH7VUTY88upBeTdtGjfPFoo1Ra/Nbk4/hJHrniwYFE
xklvx/J4y8B+mDp/2nmDcDT86Pm688E6rbgcQES1nVZu/r6QzsVXT9+Br/T/Cwsx
KdBNfvn4hQzJhjWf/nkv5uKSEFNGhj2msaoURKvxK8mz/XB0za/qfk+Y1s6gG/jZ
ezp1oLyfvl1DmcK6b63cbazA/O8HNpBAoJACry9kBq/gMlzkIJ3+iZ3hqCJONbzS
MJcmUTv1uJ7vwJyzzCnHMlnoiEo9tyvbWBSTf98miHwF6mzs0NIR/bdHU5OaKP4N
Now4KyNojkp28xNIEjGzH0Horz4NoZXQ4ie9zfpTPIR2K2UmPRjHv6mDZx04nuhw
p/6IoCqR3/D5Z06yh59K4Oyo9TZd73+xG3IlTnAENId+V48OSfhBna1JDb7svKmy
fB8/g1jr68FGsmPhYStB9reyUJQ2bY0eliM1L0NHhHA4I3sx+gAegS7a06C5RWOC
0+tOeSD10idO41Yx3RkTTz0oHcQdZlVS0OeP9+n0a2i2XG5BobSfhnghg6CaHOhN
kXPaFnE2Cln/qO99RTDHTczz6D6/D35my+7KI0wQ+s7qDA/iWCOP634zs32KtjJI
LfQupMNSCxjG+scWFjt/0VmtddfDGfpb+qJadJ/RF7/INSb9XGqDdfapspfkcUy3
qQRxaphheAcCyAdZ7XaBf64VfcfCESUPSTREd8qiss2hIQi5Bb2L5dB+2sNvaQw+
YOdyxyrS8JN04BW+u3fxtOut5fBomPNyIqE9v6fzkp+8ekdhVXsqco38qqdQ/lBa
zX+FqtWmJuX4WLieqqJzgvsGGPM66NQMzM0Gf1ylyNSWKDStZeLMTlJr1l/zrO9a
6YSGbcnio/HDCF96nqXIT4ufzq76iSF9N1WjCGJtDy6uxWlEwOfslP9GEGISezo5
ExGGVzYLme+qFBRa6T+6gu7fojVtu8wPDMh0uil559aQQZ7TyrDxxIsDZ4yfU6/P
39hh0tIJmBHeajI1SPy76wLRrr3Cz9yDAVWQpYJcQdP2yD1I4XoO7Af9DaROJ3tk
dT1aDswzKHiEKk1+IdbwqkpUrjGUjnYjw1anT6Em6KwD7aNN4FgdXAsbpkcYpypk
IIMRB9mR6R0rEuy0YkGfPNGsdfESNg1svxMAY0OqNvcwYmjLapgHG/Otws5dp/qQ
IRCyqNYAGat3WEeHp8xQmTHG/iaYNXXfGBf2VmNZPmbkRjExceAVv3CdGvFjBo9y
La4rCecVZh0oIdNDPSGYDqXNBl1YrGICtqWJtrfJYsTKpbyZrBkpdeb+Iswd627e
e+oFmjvDC313y6vq0a2tWolVyIblynerK5OQBQhQGHMP09ZrTihZt3tzS44kWV4b
FYrkjTmUfISpKXKjYgDic2a8DyCCHpdMI1jH/ni+WFEkY0GGpTInfw97glHEhigd
EVrc0BQq9APZaczSLlI8B+LuwZUZxSeAoBgPUPAxhOqpG/EMyLuDeqcFzzkXWn6t
itFFYMgd6Xh2izatz5otxJDqLZ+WU+RFv7yoHg7F5R/sztZ8HCya6HYJ6iuYu+XJ
Uf8z7EnBvKRjCoYrYnslCHZDQDqSt+F/+v1xdb915Col968Kv113zqXKyTDr6o3j
ocXy9VVOrG0LafQk/6tDZpP7Aqkz7bWHe0WxA0zG5OYL/z7rGgwJFHBNvXAvDsIX
dpvFqb9Fz4taZQsRjSsPFjTDpgPl9Lp/ufW6rI07mhLFrdmmlsY2GLkPQXbbAmMI
azFcHQaErR/i41x04kV6Xz5W4/mpwh8fo1sUZU0OyvHCwKjkG2YFx4ZTlRQ9YWNv
S2a6903vIONXi4B522hXNL6S5rXsMZ2E1adrjxTwOniemmtkvrMa7VHHnqsdG5kM
E5AwTvnwM0WhlFl7RLZvuHS1St8zQSw/tbHv+M1B9R317rD/1ipCJvbVZZ63/wpR
MV73kmFjxniX8ZWdt6eK15AzBIq2XrdFwAu4bD9rhBOd5Dy06koDaUHft3XInqXW
bHpja8qZvJh4YrCIsBMP19/jFVHD62muILqD4JIKSVViPtUFAj3owCSVZQNpfeZj
V/N8d2NGUT1mfTiRnzyCXRJfTDFzD2vgbZOiPBEnx9X2hZY75BiHFClaOBIIV4Nx
dVnbqwwwWVq/O5FtCV3YT7q3zyxXvCWSBP3QIvbr80W4ESFeZQP4n6+1UWCYv57Y
TbaYphgAqj8OrJSg6ZpW3f1v1rMwb87NgltBL/4g4HMKWlkD4BacLKAzwYDVwKkl
Xz6ZtD1yJ43kCgTtU309Lcxm6hylHqq+QvV3QiA9IkQAITze3YZAYaim9UgEZTUe
VOkoLrid7t1CM7yC1VruYFtYzmWnREUkDXF2n0K49buZpb6+31u3ecACrsEDAwpM
+kt8GYKfdYkrVBdv1Zg2Epxff6LWD6DY3zwDdQ4tgQD4HDYkee9S7l71/8ANVTBX
lVwdq3T2dozvoB9iyuziXwWD60gmCnCWxBaydBl5Gef5TxZEbmHGwP3LFrvRuHUX
NWhpA35YmJmBnr6zJcDS28ar4mKHwODSnx6CDZyamJkVLwP6sjEpBVhc1yMBSthx
GKpZaMXfJA933KU++v1G1/CdmB6BF9UF2zBCAy8o+tDRxnq62IX/FJBGb2s/rz0+
Z+KyPWyrBWXZL1aliubpq9X0ey66GlfTkzv4cG4SgUd5bZ3yYoyo2J+thTl4kKxL
SDbAup9JNd30svnUqAJ8Y5dzAwmhV6I3LHWwzT6XNf/XOFGFc5cbkFJQHytA5YVo
v+BhAcOY9COkRVsGQR2lJ1+YBYJNl9rvBOIEfKJvqNfpS8ItajkdFUvQsIf22xho
yZuv3gX8zNJCFwN4uNnNv88h9VTc1L2XUbmoqm/tcbAwU8EGGnUYjIuM3MUWhhkR
A/cfs2t0FkCNJ5Dt8PjYQPyZn0hUWktnIBKme6sEZRnvHYoeGtIbrn9aeP+8kNwt
WRkUEopRxP6GagETfx7JwDDtRBOW38mwcKyvcmk3+nfATregZQY+Zh0Bd3Aoig7Z
gSmxumchWWTgGpHAY1qv6D4J4e7QcbwtudbYBucMG94HfxYjo4unZ9BQj5w5xuwc
UwgGBkxZOfqij/oy9N7XvyLlHBu8WSJQ8uEWukZUiSFd/I6X7Uob4YpT9mlC2/PD
Ca2JC96h+7UcU1KJkJyYSRVIg9IdoZB3erxnUBT17S4ayNN9xvHLZnnGnuZ2383Q
VzaJAjEhFDhZDQ1XgPay9/k1XgrU0NdyXwgzxCMNijumbW/Ekx1jP8koo4SQjHPD
oOrCT7toBxtdOBFzTCoWwW1m7/FDT1iNPBFzWjvEJOqGMIX3LZXtM+WTNZnit/TA
AZ252M72AYTiJjJbmJj2vQLl9nGfL0rvDTyDXHgaDEB9gOVIb8s0DWRkjbYR1JbY
k4iVDHXSFkowZfJfxj24Dlhx62aWurF0KXh5rjvfmzi/lxGyf0menJydQMW9EgJw
7ZvuH3Ath9debs6A+TmONXdwJ9EAwrYX6C4hhRePZ739EO6v4e73GuZNK2WeBNAi
DX8/UQQXz2ifY8v9Is4GdqB4ASZajD89TrhQo9lW5W7mlZ+izfYqFgQkHPtQrsZZ
a15m3r+NsHWWg5zA/rxKbK2Sf6KL51WndfIKbMyKLlcY0dxmCwWIsmZxnx07x/bV
ON0PoaSkNAXTEjlYzmbJa0Y9zjG3kugaXi2p63kcnncSVNu486urDCSXlohY1FXc
8FKNp6skvAwu8IY7C9vCE25GEWAhNIf07lzSmCUL3JpJ7jGzT46YISNSBJcA15mq
A/5LcIr5LkW0hcfdOitSBot5xzUxV0247QFFfdegG2/rVOm7pRcFlxcXi76zVd1V
XYHJv8jx1NEwYgKoHK2IlwBYdYmxjrHD5C2w1nV437yvmdBbarIB3Jq+4ZO/LqM1
nkSgBpook5NP3dVVKr0kxBAkb2aMJKonO7QR+ygW+wQQ/cQW9a1fYb+bxlg9qe+S
h4Ui2OgbhPeK/AMC8EOVIgUW/CbdMwKb9XJJDFZagKN55WAiIRR0DGLxPSKXobbm
WWgvOQMvXVN/BKkcgR6ane76qkWx3J5zDxDC2pNp3qHLFLOy/XenOlMrjgSpT6ao
rzf2GuTYpOUoo4U5GyhOGPOEJHk2Ob0ziCb1T7Q6qtlhdOAUI0ZDiCsx/yxRrOqa
kqwJYqGW793qTRWDnFYTTxHpwDgq2rKxA3oDQsAG7rd4pfSFf86Cjhx4efBqQAna
Marw4Ukgzrt9uLZHbKSmLehdaBh7AyHDBLdyS5PYwEy/VOEp7432X6Y0dWcL5D8i
xOBgWjoJeXD1sotq99uomY6ddz9UlyH3vN7X3mE/6WE8yJf5O7nFE0P9xD+8c9pT
1u51mpdxcAMnZTvreYx7gT20GzeMJ9i4gllNq3pPowSRF+9Vj2v35z5eqnttptGn
v01MzpmAF9RAUmeyDxea561KGg1qBn+JoDUKP9grTyhEHLKTWmlj2FLfItmwOY6/
+u0vTShqjb4xOt7XupvlNFWlr7UtWbg468DnLC16BqRyuh15Qpj4ivN7ytkDt8Mm
U+KQUKF8DkHukAahGnTcCKBGrZ+6cHpTL/Iorr7D9jcZr0KPE8sNBKGY7xD2HvU5
MSc9n2Ag2EsB5XbJoooQCGmyM8a9vAiJECrF2yv9D5PHwzPVMXfAqCRl/aWpqOwq
WFCubS/0teNmAU5LF348LYeRECfrMIw16cfxSjfEyHn0u+s1PCw0tEfyw20R2WHy
1dWxc4wB8lt/rW4YrA9qjRVNvMTL7mrGuwSEXdiJSdKtkYv3AMnF385DLHbwrXsY
pqYf+xGsJeG3JL3JL42Jw7ZjU7Fimg0CKthlTO8nbnX6Lxv2Gjxk7qwfgyda5A9h
gkgd0hCigU6VG9qUnEVrdm4dBsMNDa1FESQZDhKdn0yQcXmjsaiiP8WWkK/uXMXd
PackxFWYKTJTPp8uhb3FcCg9gkHRc7jXHb2CcfRaajot1f2/gn7CP40hGvWupEzA
/hQIbnoDVfxryuUsy7JOgc9yOgqdO4qSIdLfpfgVG9LF7mi//sO4O+5CFg+DAE+4
dkAt4hFST/vRJXS872flJJ7cwd7Ofhxor1HresqsiVpqrIy31tCqkDXvymvwaIgR
exkpl7bOXH4vVA9GRJ5cGm3nEIuqAtTg2ChyBNf3FVWh7taPZ9GSRotKhw1r0DA6
hcgRvMaqmEM2uUCRvSIycn/bZgrC+2VL1gh+rx7kbE3cTT0frC434wAXX0vAQ2F0
lvHgiHbxX+gkVQUFWeeeZpdysgd0w0G3dwBO7YreNIByFctGIwCmp8YvaSkOQuJQ
hhPUtdSbuq12ecpjuJ15iCNx1Dtp7lIP4lUYTdehPWPqRrZ2B//wioEmspN1/PQT
Xpk+RqDgntejtwSXD0PNwjezCRcXifgF3aSiRaXmqjG+kVxsE0f2YjIe3+SPD6DJ
5oGvh28irBrnxBBo+YKFBbBv7USiARlJ3DfeivTA1Rib+SvCCGLAnBMei/eNnJOJ
vnjvUMwOuxQgnJHQz5u1Et6En+OHx1HNJBXkfvzWbAYaem2sNLv/9u9KZ1+c/zJl
VCu88otFK/MwrRwnD7KPcQvUQYZ85aOSqVw+ElM+Pr5KS+cZd4zx6tMG76B60txH
0tGL7XLNq8vBzVSGWpgwAZXl7N/Al5mTyFesH4Gen6bIluDJ4rYIeQVXLPf9xTvx
H0sbeywHFUH03wmimUeqrKqN3tJlFBgGakJ+HeF2YTzsJwhxu0+GOw9O71nGyWph
wg+6zLrOSaQ7B94vOhnmr4JeeH0OnZKfGStiq0fQbsob+bsaQ8TpOPjpjkbAM2ky
T/ATafrRIsaCA5/QYXNL5b/nLl57omnbRbJqMlh0oU6jcO/ZDwygtaJuXfFQUULi
dSoiO2KjZz5kggkVe0XQKBIW0QSfjeQtZub6XQdATzV0LWgCQgJEDRWrDcfZxSbJ
OsF7bBSaFAItPu4ENtXq4mTTeyxWXnxpPztW3ca7caLrdyA+4lu4kGRAWEJHcgb+
6D6zVRK1ThgawPERkBSJBSAqRKL4PFHA6Wq4hAbkH1tdYuBScOLPjlkeglOPAAPf
2p6Vmi7RZ3GsPbmRARsDk77gq+MVQ6W8WgyqMB4NNp+GiNS7oXVqBfcIQpvBjHm7
VkizQwAG0s5olaBiqwlI/JVN9+99uHAd5X3bvgaFSeU2MDUxfjRJjfoztkujo6CD
52EORmo1rV7NUygjphf92yVF8wXEBrv0sIL4rFZ5EghXDGoxd2Xf7dnVf6iAKg3V
/Nzr4AB7UU1jwrHHkLNJt6wTAHqygJsWCdgBdbuCfgLZE7pRny9KUKY2MNp/W6+M
iOjM2K544s8Gcyd7zec08n8j5uJKTYWWoKZKHF9XeEyPUYDGdUGOGlcK6/Gnf8Ze
nXCnYdDhaIyrTeCI9cJKYfbF2tzuByQsJ5ylmQ7BpAapRDAljR8M32c5yhHgiOJN
jh4UCQlywTbDff5k+nQrAg3AN586Ipk88Gn9aGVDOpU3B8mxSQ2W5VQa/HVTA2rw
irk4pHpgvefXc0p95B+M+pC8pN3KWBZEAG+B/CuyBAaOCg82c9J2UikzDWB/huuD
UaUu73JzUalgWp3x4ENCbspB1ykX67FNlcFZaF6a97bi0NuLIr8BSeqv8nm1WHOi
CHLqhzxbXRRlu87GJV8jHFlJu4Slxbe6zQxVMW6b5kryW+LvOF0R7XQY8Mwtmbb+
5w4QHKqX8+pzX/l+dV+NQ8GfUU/ggjvY3L2t65BXs/5ORg+ri/MJOllZZuDOufs7
t5dUBINDSzWlKnQZmPZl9oxadbXRK3UGuWP1L4GQ7O5JnIwknyO51lJG9xOHQKor
78Po598cIvCO09H57gfj2jvwTeEbdbhkfnYuPnII0zUUXTFYEkxtn2+c4LkyuRjY
1S9kmP/izpI2SFgrE6e8TagBbyhEHrCCrgrcexzYA26kPJAG8godF4NcEzop2SGN
3C+hAe9A3ogn6qhUBqM29/DE344nij/ZreeSYZ+4+iihksjlmtXYhWtThMdZqr1H
//7JjC5iRr+rVPCAiyc6n2yj+RywzYgyNz5X1hnn5DSKuSy+SWJy26lNMk03yuwx
QcspHIdSCBKjdqEynx1Zq1hGtmntNWNdUDGKzklDkWNthBoI3XQSvrOrj3fzyJ8k
rXafnxus2ZYgvPxHCd7PUNi8gZ7tfFuKRDTBZHe6Kbx9SrrIe+G/8c/ts6U2KnA7
ci29X6lgjESFy0nL+SofzFYwof4FXJlIly+wgX5f2bTrQsU70fF8QlNdPrEAoEg/
HwrsC96QgCTh+zFIbjH505aYdcFxsqYU5s3OAOlx764LX3vPCxPR5T0Su3FHbXm+
gwAWEZepQicb7csjehmX3ksUCuF5Jlja7wMtLvIiYQxeJn3GlfZZU3sRU/qJM6Nx
BKwjJCr5nlEq5MJQStNtahEFaVZX2PbdHP2gtmE6SXOimt49xPgBe4dWeZvqn9xn
dMEi9bG6AP0/j79wz2Zb92Tjnjx9cW6ydEMU/z/A/HzSJ0+Vfwd6nk2PM6F6HRyH
65hK9p/VcgWq3OKOueJv7PWpQUbQxMPTYcns+VczehAWedhsleDMhGV/dDMh7nHW
NNFNQOY6DBEodhd7tO7L7xHvopZlrD6zlXWKNB6G2ab6OB5Qu6e/RPng4cO/qn2v
AkKtMcZXDLe4m9rUZYflB2W0sih04EAAckypXQ9mnxnVRv6B3coWbJ42sldGrpI0
6H0D2o4GAMiiF2DKO8tuqt6W/xHXFvWIeQPLoj0Eun+qfpp9jLW80Me8wl39LpSx
25qk+6yRS23pMykVRaDF2CAPMNvYRnPPf7pKg+P6keeGL8csrlkj7axa2Ely3fxF
emNsuFsF1jVEZAograw/mbBG1BG+Nl8tZiJMPk1xnOI3NYsTDyTy+unLM8AJtjUg
lY0uTaoOl7/AjfZCSP/I/1KPRN0i3qzA2sOtFUoodtscXumOD+LwMT/h/I11ERCI
szItlytS4Lvlo7bWzM6076C84jTY6RoBHwurypHp3s9i273IqbLx1x7YPTQOAjv/
e0WApsWMiAPp85p94aNou4yeBNQkCSqx77Em+p9XZssQY0DX6EOw885BJ0m3sVSH
FhHgj9QfT3Xl3thwUp/jfe0cZeNoq5dUnYY2S+Nce8CXNj2Qz0GAafeoeD+naRxN
arLL2U2vVyqh//MA934y+cgze7PaXyAAzqtCyDM5P4Onbm4UquVxEjbtiu5jFNpB
eebB6gddXJRE2HirbvQJ/vrUP1ZGM2Ysk7hXJJaHMxOaoqbh7vA7IX0ZWQ59Tlcv
8mmy1XndsZyrjHxvetlzbvpYmadxSCkg+mvG6sEc6WOndS4iXFTq80rxUfJ4BLeS
U6QCR73e9/ZGVybOVxUDV7aeJbwW1iA2zwxpkKkONdNa/cWEMHYQqgWMGBNJZhxv
oBmFxfO1lxLsSl8Bnu77TdBS5FyqDk8r9bmgikv84JqgI/y4Zd0YbEgGqqm6Y3Ey
jm+HbGzPP5MEfsaqk+0G374Xbt8jlXlou1qi0loyi7/tHWjE8GtQo5oEbefyieGC
4OgQ264CXPOHD9rad4bKz9m2RzuE1vWp0KYY8Qug/ZiN8H7SWTam9w3bvImY9R6R
gzabxPSyHa/f453b3dWWht1+WuHmIfDVkGA7x4NYe3a2deIfvHomctvtDJqiCA81
MmKOlpSCt2PWqBgVU1Oe3nr/C+qDEeiuujR1YqPuhKQOB+DIdy+D6CC8zvJ7FVUC
9YvLxABH7X78LUJT4WWAP8kOlHMW/f6vhiYfU7vJmW6SVKMQ2QRThZ1UP+jlUpXP
LH1/zMCAoh8aNLX+SHkr+RUWQoDDMD08FNJUrjgHOhPNEtoh3SK1Eq255o5+5Bu1
O+ZaVsO4InMrpdKg+wJQAvwFw2uUgN1t0nutjl8LdVFo2VmHBKuqzlqNZmPsb2KE
/eyzj7CwpLsYMLd7x5/tDpeJ6jUvI32X0nRt0FeXhgOfONPw2dN8pEOV3KxucTMP
SdQ3uTWdC01wekDYAbhTRHs6n8sbqlizO0eXyLYnzFvXjJjHWHdFX00E1MNV0l9S
qDANuPJ4y6ut5K+pHSECWjj/gJpmMlVKsOCk4OMQY5dS3IFDOg2EEE+yEht41foK
CV+zQOvxUxLgPz2AAwRCJyEjhalqZ7CyHkXR5I7aLY7SnE7EEgMVQP5PAlQFsCsA
8cl3Es5yFRYUbpDQI6sCkLi3mAjXohhz7WHyTMWSeBMu0RxeiEcu3od0ogJfry9S
XnL9MOTU2jy0sjen6tR5OXHAOqb+ammQIY9PJ9SJOouJP40gEGThsruoXXtsRIdo
udrFLWfy0ZUlLOEUd/aGCvwphOuyOU77XaMHq5MpL7b4xu1rwirGOKPXDYZUy4XZ
LBuL9Hb1yhNSDkjcUjugn0ubyEIbKYdstn/EzvRh3ZiLhhN84TUAEeEfaIgfswxo
5KZTarq+SO1NDg9IbM54g/GmDPVj00fINH6mbEhgsbGJ9SBnSCFfSjL8U08AASjv
YDocPfyTtNk0s2hoAqUA2RSsJDrb43vdXYSNGbWzaU8fi8rebaPb3bCiAl4OrhMj
qh6WGcmwKMhWPfPFlhzIsgvIFrOvQU1xjrlKFfNXG5fP4xJn+hdY4gAR0uNOswap
GeVcC2zYCvmiXwt8+1QoB/QYwoXO7LGfoycwBtQY1FSeZmjva73Y25kYjw8bbQRR
DUsKoSJWkIe2JL2/hcpijIxweRQ7p6o3BiX7MBKGIrozvUQGFg86d76iwanOBQrO
pHTy9xgBDqE8hRn/mNdefU2lkWvq8FzVkJrKRqakqJUJec8Hiq9fWXKbC/EjsOUo
/m66/8S5HuGp1e3CNEWHWpPNfG7WeSPo5CX4p8eiCcJZjZQA+jIVQvCE6SL0WJq0
IcHDGpGdB4KfmRJbyJX5m4XoPF8ClTbIoR0XL0cCWNfwYw65S3q4GbSX5CGZalNe
ucsxMBGj1h5ITefabhM97ebUAi5GMqOrAqMr9C1ws6BN3lQwzsWDtQy9ZSt3lcys
tNXzbjGQXfUo2Wlwlb0gqci6rOZC1qFyifgeBcdUy1nRB3UChOUR/7N5NGGh+4pz
0DUhD3YV9V+Gt8IMG06zwlegrmizhueK4ZbdWg6Uujm8SXVywx4/rjW1VUiAF8Vq
pfMNNzaB0zZ1b6bv71n1YXYn2PChPHTCTODLaYdfCOw+XjKd0d91sRe0S2D+xfD6
lhb3Scm4PoTcTOZv8DiCcrR8lEMMJnfT10VuJKobnV0FLydce6hLoGf09g/ypw3i
K25FGZEPqjqJSUyCVL5SrJdYGxb2mjav6X6SfiwDNFgDawemS+fom6aJqjx0Nwuf
A1vHmAnBINuaXvCef6waBIyZSM2Dm+AvJN6kHXdcYyp9zWvAtKrr/m7j9n4ZTwaB
a9/z1twPJ/DtCO3Mte+d6UhmfJm7dfEtmGYTeR29sJyl1kIYav0YVb2qBGRgB8Pe
B3vya688lzKFCTutV0VPa7FRoYuBIVYkwvJTyekbQyEmXJsiT+eDDwyNCbzNbugP
sfQ3/TZZsDr27Ylx4YixDZKZClZUv21dL1X+EdelPwlPlBHljJbmJSGMPWjujExi
OUgiRldp4InWc3xvhtP1fYlrgRpE9DG1gm19q30mCuUGPgQVOg86kefKZbIPpRpf
vaD9urhyjPvhHpXf6C6k84mrATApM1KzF0T3j6mQUsz+Ne3sgsdeDlcMrJqZfIFM
yDIZCQ/iz7POTmDAj7Tt1b1VSjG+tBBTDDtxv58EOjWXT0USBghBCPSy53VeFItH
BWqdIEC7FEED/7T/pNuR0jRDTMD4/QQ5m90YHju7Bm2qT0sBZuRwXFkSVQ5+HlB1
lNkafrbjmGoQ4e6vtlRaTHmcZlgKQUQluST7N0zE/LyWUivWkc8tnUe3fj/xcaRg
LEOOb7YNL2uuudiDNjVQ0LlHFk+ozm1alDEQNyOGz6yHc7S1qGuCAgFGCZiwPkuQ
E9+2TgU0k3badXrFksxnDCQJZFKG2X9TW93QpT1QbbAcKDLtjVSchMt0J5SDger+
FY5owue/bbBl1X59ScFllxCPl91U5o314h9YJ2+H9zRw/nN2eM47FSv9JmK7NVl9
5nP2rQU8JQX1F26SavC0MIdX2Rz4JyXscfwPTNMnjF90MzB5TtPazF6L1oq8Ybl/
T1Q9sZ7zrLztow0yKLtwQu4Wsk5rAhvJQ698AJryzV0/U0zRCT3Uod4AS44iPR4Q
pGCOicTIguHxEMjb+eV6D9mQO81NB27tOYWuU+Q5+212916vVuOJ45ywXraHDRD+
cHNV+iSRosMBNj5OjpqUD4Ot8vae9+6athv5jJMnuaGX1kdNJBmRAMur6nYaRGT1
q51p1VYi7/zLYGPrsuXtwGtCTr5n3NGjXZJ6lMF3v8FLmOvHHmTZ/OcI4bqvxW1i
W3yVJV4M/gUCuL0u6VEJG8xR43wlAOOqNicOnjLYG5xqjh9igTWG6aH67wzy/Ybt
GOV4CwY/PSnIKCGU0ZOGx4eBUU24tA1kUyybfOkiuPILETn5YUBh79nVLKCn6BaN
+VI0hrQ1HNHC4irZbo7jVtc44n7R2vd+49xoduQC9ja2+LO8FFuS7I0aZ3iPlEDK
3WjxFm10W3myeEOJYHRANQ+njgETGnYg0hHvMU4hZYde8sCpu5zApLJw8yEffVio
AY9PxgL0Jk+4QMf2Wqk17DnBfYLq1zEu6EvFOtTNbYsIdlu7mPEG7sTg4lG03BMo
C48ieT0T6d/dBhpnacvnvpfncy4baEqZxSARbq88N2ULQgivjd25Zdb9b69MY8bs
f7nzvDg5wEuKHRxtGYQj+Y1ExqgkHd9Zodn+AChvqB3eFTaMaW59uzwxSJpt6+4I
7IMzMWHpwDx6Hu3E2QCo1VQNdkX2NfBUndEVYHa6ws/xr4OoaePnSG6pkKzmxEES
/sU/aekYerkdISsTut/hpeiQQsR0RJTqV6h2x5N0TObnj61dbh7iQwSc/7CIQrlU
kpB0F5mM5xKQ4sZ1ETm76XRTC1ACyxKX7beIlYpPyNSvtccxexKhfnyalyyN8dTL
pu1+oywemeBu8mRBU4JhPLQvlkJmCcwk5fQryCkJKhZ0Z3EFg+kaH7QfPhOtFz1J
gyTRNpB6QYC3AM22yfasNUtiY8JvNXIEPaZauqGNe4y+1UzKNtNY6JVRnfARaYuo
20waK7a6FIjXQUoTan31Jn7HacO4UM9oREPsJJ7JY77otBd5yaQ4DwY4xHZsx2sh
XNDK32ZOG56EX7t3dZsCoko7E1TIJ/Qlkgvn0qPya4VqksVbfsjCRrb9cL3fQIvj
gnhA1PJazWwoSVze4vstX7kM7oPmIjuY2QjaIPUhEmRI8XEi83weypvPrP1gLC51
5AjcBKn0eshkV9XLXWUkQSQpwLoWpJ0hr1U8QakcJ/U3W4GJqyVEzo6zrZgU51vH
x7/31n6edXOxQwAVjCV4iBTZ5ObEnMse+cwZKJY6sHQOgasokIq5iqAZ3yhTzxuc
Cm7ymgirLoMwfhEIrzN3DwvGGXxgaM8VKzt81QdYa06GvZX1bVMPONjJX3Gay/rE
e8RABvr2ondEBdVfU7yCtPeqb0+zmMZZ8fmcP/RLjuDaNPA+4MXIjRrO+E4dokUS
cCzt1xkv5wdpWMqOTnT7rM1A4ZbJSpgDoFm8hYZ/Qf891iYcr8xHOxwGDronsGdf
ltuobayicPTNWp9W4G57w6RkRl+8B1Dc29hFs9feD/61lbIPZyKYYlJIl48uTLud
TmQynDwiqHBkdxskp1DDRXesVoHyFfUUBnnPwX1d5UC4UIQsIJ0lV+7cyTsE+SQD
iE0B5g4YDyDM3FaeSFDoMvA8219w1qWOSwb0TQvxz2O6bO4Z3+MfEd4zg2pRCe7q
UUXPPTC5dRlI1R4KXMQd8O0qU/22FI7bcv4T8baxC4f/pMzSsP7ZFBRBJ6Hmr+/a
+nOIj/TX6d0KhrJ4QJfo/xZ6Bla5EQPVTksvJqzSok933GIO+ubXpqiRJ8TwXvU1
qm6vNksF5RcB5RjpMQXQcmXzfAZ0K+WVI7XXLOjRFCW7hP9lXgTQcnrAkGyoRpr1
gQ6xuv5d5xNUQmfh/QsRMi2UTjyPNZRMft/VA87pi29xk2cNI4P6LAZDA64SNy6z
AfLDBuoYbZedtGI4NEE504pICq/wc/+HDqH+SBUv14jvv/h1o+It5XJLc56ZwK50
Xskdy0mCTqDQCFB/+pWn+3xCiGmnalJrxB8FsV1OUhEtw7ffbIXc7eYcqYmY4eVK
TK8jxZWee7Bw3tZmHyp9jYrWBNA1VcY6HmeQwu9ZjVTzvI+7kpAHjKnlaeFJHW55
IBdiZZfInOPaO9aAWuYhKjrSa8AzQ/pIV0HC0mVkqWNWecCc4NFMM7zitt77POx7
s/lmp2nxaNkjVHShfc5WIstcKKOh2tKRUcFEPZOTC5maq1z8WsEAdx3xBdqZXgwF
I5jFdfX8UMOAelUSGDK89XgF7DayoKrCAtAcWRv9TFEVLlqABn/Px+7y9KjUbyzR
6U2e2WWNaj+K/0N/LOtKZfFWCGzvHFS9+6saiXVDwNAZw+q/YO/ghW/GNi9BTSFn
2o6Wt5RfR8lKUXaAzUYNaLrBr79mKANcXNQO4FK+qftOQM48CI7kbqctu5IKhhpu
Lkp7y+HlIwItXk+niIGXZPPTZCn9Tal7/3vqUxxmWihhfjWhqTY+nVCu3XoDq3KV
OgiL3SKg0Az7JqvFnX4vS3lZVvtf2ZbO3ia977kSjorG/lOULcT9dCux8slIegbP
WBmL+xFX0fYwLcLevDO9ho1lfyJzhcDlzgSY/FEsTqro2Be6SCeAxPz4OuvrK34G
bWiOJne+WEhX8/6pCVF2pdSGtO1PN52jepAFWrnxZGxKC+KDSXTSOCfNV+91ZElI
0bx0E/RmVUxAwxhxHb9ATQeOy27NUE6FK6lQh+DM5IfkPvPyMRP/DtpXRgSgvDw3
GAfMHUZo7HJsQsSeZTXHQqIXEeaXhhXaLjl8g1IYk3NfkaEh2Rlr0a73PUVkbh8W
xkBBBFSIeMEsQvl/B2N+jEGMnUFxiQYdiJGe5PvmC6wcak4LjGwN+Qh7eTUj047F
SuHuhlbhXES+++EWh36v0Lq65O9zCvxWuupsziauWLZoPfnKpWP12EjD4tiNielX
7SrEHxUJLW4lZ2ebawKmjzBURcDMdmVOuWB1trtVbV8tkYgeJM8lN5IFkK4KViFv
5zViL0Dzamo594pYWqeHXqxMxehIjJiRGSIIBoisgYA59HclUyfUYb/L2B/hvH0Z
m6ZhyZ/EJkILA2SToOAxLtiLr1nOm0VpdYFNBoJZzf8TJEJTFsxkhUo3JsUFgjzY
q5+d3PhofIpA0d76AO7pBeWPmhJJd8FQfETmbjVvr282kGiSKBfW7WZ4SYpHNjCo
DrZRHri44crSte95oW/B5dJlJUgl0aKT9oMlbl/JN1frluT9ddzs5PIEsnmJ257U
W++h/R4bxi7cyi3iTbMJ6gM/ZqvvoDfr7wiDS81V5qd1Ovlb8ii21twfVRpEj2op
ZnMpvEfpAUSO83U5stH64ktl9+Cp4xEYy4fGDbOLGIa8wv3aNBAcZ1YU9O65Wxxm
mAu4crBUt0kOEFqVwJwxRoiHszHV7qAf7eRG2cP1gkpxxlOumqC0J8HgvzNVyTOx
RgpDlSqLFNBW78T7s5nWXCFdZH1xnby/xvk7uRbtoPUTEYwQvu7v3DtoaXQOkyVd
W95dl+MDO/3v+qTLDQxD/1DcBRZ4ebpvVqp9JiXtPFXd6jzK+KBP1ekpIMvLhZme
CErleUqYapkWZFnyuGo3RU0S5w5aCKKPrl4PjLdkdIWYD/ZyRL+/0P7NtBcHU+WT
sgR0cRjSbSxY9JPm8SKxt3TKZAxZJQeeVxFyM5ttIa2XM/kgfab8HEfvobWEQeke
ezSjjZLpaQQZTOjDoxCOOvXNc4j7ll8J7qS6Emg1v6VECxaY5Y4+GMvFZNe45Gf+
xyR1evH1qMv4p4aOKp43IKJps/P3lSLuFgO8wLsx16ereFFH78dvCfZvTPO/yKkk
/Pc8Akz5ndK2FtOhkPjV0t7OIlrrmYtamOMnds2FcYLGTDw04UMJGy4XZxI5W+Dc
axVi4jhLD9aSv948kJ0ybK3+UMq6H+MTt9iheZqDJY/Q9TwiCHbjeEC3X3IMbTW+
nJn/ZGVa+RwgduqvWJN61lZbbs3M6U+/Y7HuGP6Gv8GBHrEudGlM70LTQcfsSNJa
72aE/knLHwqYBR0Gyzn0VdRzSVKkWOBGDBTaX4T2/pGYUxc75yjWRwUhh6/K/HRW
1JWVQmuYnTgy9e0ovXCB2os8BpivVKeDVNvsmId2m97b3KH1UI8kkQRvr7qbvpx6
JsrM9yRUJmlt6mtStqUZTOQaCAckLK1BgUM5PJBPP6m35uoIWvYpDu4MrbESHw44
xJmw8s0bL3bN92taDOXgFQ5eACN3zsfZP2ujI/Vee6Y5hfZSbmGZXuMKsHBDOa1s
SsnUbXBHsCmUxxXybEHQ5Oq/tT6JQV+oaTV4JSD6axMffxMDHByaXqPAVcOEroaV
yL7/iPB0ZNDOynWr3DWGULaZHaKGhQD9ZHBjpJ/DSBjGU7tCZa3FI1WJxz0ut6wS
YxvdIn3axE/HThww/m2lVSBDfiQaMKnaPHG8FlwpB8t2ZDN/zhn38xDXRSYKml4H
SaCj9hon4O2er/dx6lVLlFDxIA6lNapoHzwbpny+jM6kabB3pADvhZ3N8vjDUugp
kDpOUcy0lbCxSO1T5oqoxuh7WOlNFgobJA6MgG2Swx5xlXVoQMZDLOSG4ePnZZcI
l28lPhJFgmw1lgeWqRbo2njmq1J12EIhTkwDlsunzTrBuyq9BT0SItKPvGpUWTll
iBWZdrwFQ0/Ur26nMGq81TDIgJt6N4Sb0qtZ4ON8aCICApbsN1v06Dmfhm2/l0/l
K9oh704LXIF4LoosntfX6Le8oMuf16ROlCCYyFUHSEQsPKgfaW5IP+u8Oe+g1plT
P8rsUukWr+mPj0XFKmrX4C/ThhyC7faeB+/OMvg3Vb8J9uo+K0ZcR6BJUpfSWPY+
PUK/AX31upTgP6qXGaUcvoHVc/vRk+OWbndeMosAfjtYcWwdYRtXAcOKdSFYFs6w
1ws8NZfe7nAfzUJ4prYXrnlj4O9uI7mDcREuSsimTul3WN5hDKlCI1psgexNlmbA
GpeldIJrb+oJety8w0Vbig+uQTDoGFlZx6avZKMdUsuvjLs8c5uTY3bNTEvFtVBL
Fj2I6DGpMLbH4HU5DI3tnwgIogCSmUyzwXpI9XX6BpNaUTsuUiH4EAPZtZuwqf8u
sMfesDSlIyfBCHS46uk+8okybEr8EmKcEjOUWc7q50w7n6d6melli6ul2mZNbFgU
J5QCZVzqOES/ZcQsmL+VV3Dud67DMP7ns/emnjPJekWGJu9TbpwH5I3g3MUPH4RW
35mNpD/xdYH6bNzU36GrCtSODtZ925y2S8MaQWTNw0PeHe6F5zP3bah5NHN1Cr89
mGbWU5BYUF2SnjD3Xrzfk6A22AoC8pcxV12+pi2vWZyGxzhQmDu0DjI5GHzXVb3j
pGsbYCKT7WGzPyrVrfous0m8GJcpQd6vlN63GyhXVOP8gffWa29MAwBYTBbZZAco
ioql92SFJWU7zNgqu6oeBIzipLN7pgJ9/lOU/NGZCIwuOn/x4catvBx6FdPHgYfp
1xM8P6MbGAu4BQUoPs0+pJJSqWlD3AukNElznr3yqu0F53mogk/cFWGNrrGdAo7+
d6oOK35cQXJrnEjub8ZgXPGZi/Pi6UIC9XVRFGZMBJwU0dFC4H/L4kjcQ9YXiRE7
DGZO7iVcAppKUrEQqF2tKGJ3j1PKPha3qVdIXWPjC6vprGY6yCpOw1PUohp+81S0
FA+BRDzsrw+mM5Z4SW6slBWN9RcWGBK07CjfoPiK2KfbmCreQWVXSOC2qBnLnQ9m
yYZjFxitnWC39wiibRAubYEuI8TFlz00lM46JqPWIgkrfkpa5gE9gwovzv+TkPO5
ucxVM4aCtcPrf4trZrvUC/lbt6bcl2ee273UngXe3UEXR3/PKwNHeNsZQz3Qh13F
JkCBQc8RLmi2IK67gAu+hyNiHd0j9pUBTJbKAjjLz6HUu7rO9OOn4S/E7lQseVP8
EqtP+x6tFgoM7TAB5ZrqwYAVo9Uq4AOJpFZxLQt+3tq85vuO4y1mJC+4fKEefSv+
CEjCRLCR65L0h4sZbUC1ERKGE/qxm6U5sFMkZgzbXQ8D9AmmOz5f+mkt/kg34+/U
r1r3HlwVWt7q3TWAEJgkuBtEHGeSvkLJXFX4yP0CjHe8gmLWAQ3cFVA3PYU302hn
CZbmkrvdh2lznLOsL2/xvgkV9bNF0oHKfg7v3DeTQpOcH5fDaLZey1NhTE07ewsh
Y9D23En8U9k7cqJQD2ifm746xXVjYXvfEV0h54pVh816eJy1s2/Ie9WGFPO6naDF
M9C+74jmBM0jweXBA6k+NKZA939X/uMkZLbIGHjBieDw73LoAPKItPR/rn4ODsXE
ccv8fZeVPJpu+Guox2E+ufHP4U1y7SZ95+EtmC7FuTau1kcmL6nX94YWP76Ah87N
lmIgHksWoHMl25fqhdasKHqsqv6mL9W6qfp3wkUgWjBWQdWcr1DmMWDeYfioT1yl
N2Mx1o8x26NouNpGbgxgCw9+eC7HwgtQ1QVpk+QX4h6qZZXEKC1mtC6hsBHFrQDf
oUougMjEo76zLjbAILTDewL6gNDJv0E5fvfSyqsYb83HzSQMWLMywUhMbzuvBaVd
Tdz/ctUGc8XF/xjcWCvFQG9JcGMcuoaEfStuWbmwdsbs5tV6JaITtd87WDTglHYG
WhzR3VYZ2rGlvI9k88l4xJAA9J620MFPEp+Xw9Cs9keeFkIk/BAINYvPc17+us8V
7Pq4y0qFB/xV9I+ozRrVUse2v2KMi5VPdMnfwoUDWgr9ulKFdj2jppNjHkTzmSoB
3/zhwOaX4FrJa2Ds8Ps7u2XcRd7R8/m89hjAxeD3mK6yIvY1eVrKkER1GY93l40x
qbK8TC7jiTOi4KHUXYyOotyyUFd3rRqHoDM+uR6sWNHCthLBhT95ZG/eC+4XaAt0
mCgAbHlVwf7hpvCffSsGfTOphVfL8AqulMorL1GAxi62q7d+dNf4GSZuzEE0Tom4
gMLxYiTwYYvZowNAGmmQ56z5vJZ2jLuGHDuDe/zK/wytQS3ce8ecuXef1OZeybSC
DVLOrh1Y6FmLEaNamU4NySeUYg3J1kLDExDWBHkuXCiZNJcghiOR2zblmA40lvNe
7E5/n9Raz+HX7SuSggaoP5VQvLZd0+z3xJAYCiMXjHevV2CYW5tukxeTodAe5sQ9
ZPR7UP8a7ww+KpnLeXtCJoG39fP1Vkq6yacFQ2FrNoTOp1Ie6tSU73+moRl6BL1m
w1OonZT74cpxZ3iCSVS8JEpcUkGNarH+MbhKOviPP2FY4JEXOkZWDnE7Kug93qsA
R2Bg/+GlKwTe74d5yDD+gfZI7sDCDud1vjKh1sa4ijbpAh65dYQx2hsOywF3Gh7e
H7AAUOyzQ4t41o7ewOkRjJOMG13BJlbkGeEfUC6quk8rsZUn754n7AboZeYh+h/i
i0OrWkq6E2zQWB38fr/hzMat5iVGEn+RyGr0joCabnXVY6xg+py9AX8wK2twHk9o
yyuuDA++ttnuAoP9P8F9U+cFyDImr6v6GvlruuoTQazsPo2twZPoXRlA3xT90wTk
Tv+Dtb4BnV7qVPSc/f+7R2GAp7orCsAwI30KQZmLWAaz4+/q0NQ60h+HAcfDcwlo
k0hcLhzj+nLASS4mgUt4gdN2CdtEWq2deeX16BETVeFuo9uF6TIWsCz7mKMRIV8E
X2xRMnhQVcabMRErFOoFIHtj+eNQvnnvH6Hq87j+bwm4v+j2OZRSVEkqT6UR+da3
rbY2rwE3LGyprNk6wERinB9C6tf01ZQ5R07Ibdt81ZIADKnScyvTlL0UrMDC01sH
Xf+vQAYPeRu/aSwvg6ojMUScgW0HsydyNbR4ODpd2mHHMtBzfQHNMKg5CyQVbtVh
V11biBTCpaEgvILbXRaQdW9fvFFCTG+/b7Btdv7KVoBlLA9ynyYyL8hShfLEXBE8
Owawo+4XXyP4Wr/gvx6uSF8MESf5bt9FUNLr0bU7bMofBmlVys93L3YcVi0UEGoH
0zjkyTjze5PhJTlvcXitm2phVlpHh9yVpv8jDCn9dAYVPr8bz1KG92rCMp7UoUlG
vV/k/aI5DD4ND8u2UUc2a80YLhaEAZR7vn/7VrnYLb6T+ALCei8Oyd/dTUIF4apx
mJOaHeJoasfinzzR2r/h7YiLLxBgX3/0x9Vp8Zc0cOy0NgIcEvsbkb74HfPOgx1F
jJm+YdHg+ntaCQv+MA8Kv/zeJbXoO9LrVJ3pHNTw5CPRKedZNVpU0B3Gm5wMM5r9
lU2619wW+EhLKaMILdSPAvwG5QM4NNEJE+IFGmxjljv+2OE0BX72PXbyuMH0zO4+
zjgfOAWwruySnu81tFFmDcGbaTv5H+PoteT6Xv2xlVAPVVVtgIKoZ9QRVAAEqFln
nryZprIrjVyCoyRnX5wWqA8ejKNHHX6c+Tm+wneQnkiVz8nDda8E+1J8DzrHBTSR
fB4vJH8tjJLfcjScNw0rOPZHrNB12bS+PLnVIETh6zFbO2tmq7ElXrcSSHE+eWqI
4B4cmvOsN+sZdeVLZGZAJNzZ0vUU3atXm/i7q22A4NBRPUkghmBYVNM3oPBDtkUw
tz63NT4RDtYquOjEirahymUneAMySXStUgVal9z7ZVVLeIDnIgdSXcDsZ6SPfIJp
81g/Y1JII9pKfkRmLwDvbUbEb8m18mfqwA5IcqxoFvzhuUbJR40pgegGnK8o8lJz
AsydQb0DpljTz0O/swAjTUJn32OiKRoN1N1M3TUQrEeFrAgWHAEBKsODwS7q/pye
kYtDEYmZmJG2tozb8cl6wzre4U9GemIZIjrlsuTvN6P5lt0mc+G/pEjxL7/4kjlx
XG4NGzfrhsxXrdzTr74EcA1VXklzUR7qMqqm/hPYwQJaBgYyQj8cD+zmjTqnxUCI
I5Vz3jlKPrQGstCITcUlvCs21a3EzRsTvIXrmPFf058Y7GuDM4bJtKz5Gbj9UZ4V
zOEwY1YACVJKX4bC6Q1yOF85rM7ntOqi5LGRN3goTqzlvaV8XUlwbJ8/NWWaxG6U
yXjW+UomGU/X9FKP3ftLzK0i11duTY9FF2cQoN5h3s2dt0wh5pQTVrvvLYCWRRlc
6fNOlIxWpu6u3gSuRDB6EmJq2stJyEjd529GFpu87Y8mPvUrMDK9IFH/ZlmXAEcB
eHKlN7T5XlzzTGHMzT4V70ftPskqyGMSXrBrpUp7olPVZe4XOqrSwBcbNPRM0b0e
mN2WImP2G6gnqzrfE42UgJNv/NaoQplNEpeuPOfQdWWkFJpbmv1i0O570sIK39JT
CUSHGgBF4OLkYX5rD1TdBox4HWCy1HDAUtUB7N47S59fM2Nes5akF1raTxGvoIQQ
HYftJe10e+5xiWHV2JOQ1O/+X9ZI6tVHoNnAjNhSY7iUgy3Rjs6Q2iRX53G+780W
qnKsxw/KTG2hzutcMUMwDg0ZT+pdJrGdtnjMeZdxCcViIm4tSnzWWQRFW7HZXJwF
hcMO+HDRUzXynk2isPSAIJZIRZ9iG/psHAW8xVozz+3ipAfH8LARQJoQu3CP90ev
rjpmUTvmUnv40ZNHAKLzBL40xHjoLbRFPWxxtP8JaGqDf+KSiLCqJ+gfLXjv+Ag1
7Hi85xrmWDaPFPP9JvWvMy3ejyWiDwYAjm8ofBPu7fBLLz+Opig28JxGHeBQPTKi
pKQg0UgkxOiWc8nLamAHPBwcxF3lHzL1b41OsCSQ9uZUTGSwyWnNmu7gqff3LWGX
lZGKEK2rlRcmC/IoqkPRhkuxF7KbjIPO++4o1Gi/xKE59jZqMEKdvnFZOfEBA+/I
ajgxjWYN1Hc5pajWHm+iQBZ3upStA/wLwh9MCyULTGPL71yb+YFVJcTHUX9MyPk9
GfKevsS94Td1JeOFj7T+iShOxyauVONbSdQNfzzGXx8cPpRBanpXy/yLqQ7KVJd2
krYrxH4nZchamaPFKMRsYbsdGvtc1+MR1cmkho1UuV5g+PlrKKYo+y9CISfTlkvZ
geprMjqi3s4uQaTH1SJSQHHslQF1/r1ATtzUdLQn+EDrj+h7PtT1U8KT5A0w8uiC
LFuYTj6VKk1A0GF4/FbKakAxPvOVjZQIqMLVPIPY4940xa28c4lQ678IHXiPbwK5
TBb7Xn/93C+AudlPkqMZTuvhm0wPUmytV3vg1JB1TmShb0tXv1ksrljtJ44Bb6hU
6W3fAdP/Otf72oqqn7x6ipkXdWWCG7Q/9xGa86sHyHoEw/js/4Yjc6Dt+Q2xOkBq
ox0Nti0Q0BoT2uNsCjay+RsyrZMAPXbnMM1SGSrseDYzEsbIya00YR/lYM0hLVM9
+m2zr+TzRnY/o2mOKpUJdNtLXcfa1KrMRWaVMMy3GbdwV01OMrBBegOHXDNZKa24
Xzwuq++qI6Q/rW4cSGJtTigmVmY1lDxZwo4fjP4ZBApcxWR1n914L6hOF6GvvHqy
/DHO/o2AHcJJo3wsdh95/SUOKH3myk7mGZ123VBpVmmwKQ9fQteKDlLidLHwFvl9
EDsl+5F9oI0NWqQEAW5ABsVRu7w9LJ8og4VN/ubbSKpi72y6QlhiBpSXpS6FZQi9
0d4WRgGUpYGXSogI1AZkbut0VpFyueLK/Vq1/V1dhIQxBmPWFY+Us5YG4ethuHlP
23SXjtYwJon0LzZ+7sM2FLEWFZ1pO/PKnhOFBMtBvwNF5DP3s44/EIax2xC+L8EW
6oUX7vlWxdqcBT+qb+FR2lGJw+rFGCBU7TenNKh5jT0qoDmccUE3aC/rl/aWGxBk
YhX1DrrhzhVVBaZr+Eu79EgiiKrWhMnDvCquCFrwNfKKN0LPeKkSVRo9m8I7byWZ
/q6IRZH89PgxRT5dSp7Ms5FkwdxD01sb+n7hAHl5YM3o3THuA9lF689XsIo9B8H/
7q2LMPzH7+prkilMBCXECVZZfl/htkxTvKmMQqx3aH68fqK5QzfacQ4gMBci8PDg
EyyMW53q8jZmE89dfA1cJrd6ZV3VlcKx7KvHc/DEoVL3BBukuICUsAdBVr1EXDIv
skq1Ml+PfH/P3nkVsS5nZuktC39qcr17eZPMHFb8b+aQ/peEyLfU6V6w5SolxvOO
CuydfXhWpHjG/L5Aolxi3esgaSEGwa7D6p0V+PYbr/NgVyo8Q/wgbELfzyEPT3MC
5XEhD4G79AhXqaZ9TX0OZ6nt2dBazrrBwo32UE9PplA8p32BDy42xkPz/uhEuDep
Op5sAmJsEjazUNYUCRSBKHCwKeA8ty8TbPrxWrsY+WLVuuzcu4MlUoUiiCpjhN5r
geMou1earDawgSufz/hbCqLvfRshx6USQ02RGoFEURpVKdvu0GkQh6EfJN7JSL3i
Z/BpXhbfndJa+fe1htIiqTnYQP9tbQNTx0zoW1bvM40Nl7GQYeV8xRNoG837LHa8
JZB1w9p0eZRhkRxf18VlRvDUoRpo53+0AR5tP74u30lLDShV7GD3TLDiuZuEI57H
rEzShPSVxujP245f5P+YTgUnZ5yYQ9Y1ZCfL+OQ+9TmyOHf1CGd4lMmocHhZLLZ2
NC1V6CzUXaXx8Is+6Tpxkgeikb7svsSjt++d7B/tv5954ywP8ALVaWjeAw0jSxx9
RabMLgMFO27kKdFBap9Kl73CZETWLSFN7kb9M5OvTjecAOo+t7LShyvLF8KfZ4Cr
MjuwAYSKhmR6P5pEFNk/O+EwveRK/g9znFVXwjxNlxCbEHtNLGAclRALLEMech00
fmXB2Gsvf5E6MX0Qno78uB8dz3wOYDMjEiFhZ3vSsLBfUfHBCLlRxsWFrp5AwLmz
fV6yz5n4Zc0DG4MtnNl7mZf8OJPtRbRtmmv3Q0635BhTRM3HupYQmBLMeUzJZcgN
AfoBJ0f+iLSrBz7iSoJUw60fDSdrFeVsud5HQnTUNnNjUMKdjekt3DShrjv7uc09
iTiZtmMh3UTGqM+2iAq8q5aPupGe1SSXWXi0dC87knyuyRbby0/F/mgnrWtAeJXJ
FrRSPkOuOcBGFTMS0/EF7QZLH0Je3kEm8Ta+oOHbCi8M8YVGzoGt1k6Bu9dMAHJm
KxGiQVLJZQmQEX7SPB9AnTP3oXeTRQVAG+3sjiS+WmGsx/dL0JrQPYrGSOsvWuVz
d2rfP+jxaA5xDH+9jP7HqczGabAaFo3/u585wjhSoyawYp4aYrsEWjSGcLqFjhU1
YQkBYan7VzxxE6zSdWqvIVB0oRy6JGyhkdWaIdn2TZfgBPq7b60BDz3PESoER0Jm
qv1dUee/4eSdzbnn7AcBhSG2qxiOQWE29dB9Bi+45AB8fil9HO+rKUk0fD2kQEml
CDDEUptrgYDw9WN6OB9sSNCKKBEu8aTCK5eib/dEU9vJAr/8GNfHU9x4gKLDI4Z3
/IfdxDdVkObjU3BGanHQ62BdRgEZarj6jQH5+qUJb6FXgTh5RzkhyvfDr0u11WhO
3H52BFgpGER6fTlRvzS1u9I5QDNR1FPp/UBp9kuHQdUlJyCVR1P74UhlEMBSCbl/
tttTqEEghSfhtaEuki8355LsWVMmWCiJbAbgYWNcS+VmAUolGZgSKIdO2g1H0Blk
ANtC6TO1lrqxVKD5LgvhbNH/q1OXOFxsqKfdgKK0Cb8RBYduJxVFVy/pJjTcTnaV
W759WDBMpFP+3QorUNbt2zbIEA+DFgg+SBPOPIEOdrGd0x/duxSFMoX7rqztX8Hs
UG409Eys+JPXL1qbIr4wxZM6bIQQoBoSKnjBsXKtY20tdKNUjTFx4LeJTrLOA6Gf
SsbRZ5Ow3AKObzvq8R9yS63aNYgfeY+wUc+oi9trTBUu4t+nXYdDHb1iNU433Bxu
xACD7S4pRNYt8Q4s3nc7LePIv3CYDjyJBxfUeOE/UZI5LqHvyHmL4QaUBMS8spjs
HXDY77fxxaRZVx1ekBFI8VXiQxFrg78T+PzQBBOf8+cyaAUvyaTl+6sKil2KugIk
lHl3GrIvuEHXFF6AzzLgdiF8vXeurTwZBfcrT6GLDmx3oyzRshYwpe0c43k02IKU
IGLpXNNn8mMIyo5PdbEo4S9HnoL3xcW1u49/dXqV/2bkSveSHwhV/KN1muAjMbge
322BipZ8VwhBS6zTwcveVfX7zhUwCP0F3dgsMTs7HJrXhBeoAczu17uWQMDCCshl
aWyuNbjRxzLdZMD+RA+xjJyBdWErvHz0kNLpFTnfn7vWJ7JOfDFfQwimMzgh56gN
LrI39TJSouUWDpnYz4kkuz70zD7aKE48CflwP7kE1g0PmegnHNjkjxnmAouondFJ
C4xG8eRNiLHOpivEurCUxovmB9X77tAu9lyCOoXd5ecUzFeetaDS4MNQPYGPXmVR
+R69DplpB4s6fF57BDIxL0SpbblXtRDsaCZ7kOetvaB56fFzPrfzKDNUmxVjsOYQ
siU+G3sEuRINM1QGQvnzGDcp4RsYxHZ2NIVHHlg4xuWo6buFm33u8KsySQx0rFHr
XKzSKBy/uzBcamO786oM37gQR1CAxFzMevuJhW//atVhlvwnhadG7LPpcpmaouN4
dO0jBuepGbuYxgq02vmWdY5/V0TA97RfLSVGlHugEiYzJY94IOc/eK4K+Wwpm8JS
8qTHetzcpqjRj04q6EBa00ucOJuZJFTopXd025oWETfAHSrmvPHffBUhLeNoaiyb
f7nOVxnnXQ5m4JnBuH+IEFCTrVuZQlbV+t2xbl41neGGNDbPWjp0+Gv8iOrjIQWo
PRb8PRbUxnXjTs/tET12d4rFZCHEwv0NUIySzXK55bKcR07Zss+v4TuNfnMG9mSo
0VgVqjMMKAWdZsqaFEsSLrWMKjCuXDx3n9DAlW0tYwMR7t0cQCG7iN0frnxprSSF
NE6EZU0MwzRKX3bGhDAsuyKoYSphuY4qH/kDCRCXlj7zh2bU4xUQzM+FLMQ22R6W
cjPPjrayxvKcqhLkZRIZjGD9SrUDwPjcpibkSvZ8P7mEwu7BpJwrd0ceCXRm9Hsy
6n/S9Mn6HrS/vmFByhM040Az/akIIKO6DRVdAWTIl3g0W/MGZpqdaaWZh9sntN1a
0fxQPxrQYDv5DiqlHZn8Dwu5LZA/RJSJOYJ6orba+qkCwTNcYWTL9NWU/ag1kU0p
fWRxphukUCqcqJddKmTyw597rUjVvu31o+vXqW/hH0HvoRM33TNB6icWRfXiQH3m
QJF5NZFwlAOuHKbbsT6rcgOuoJYwv4NybzbT3nWt0y2MQAWBXKt2LmZ93+3IXg70
u9FK9LCPrRk4aGACrBPw0GTJqOGfTWI0uW3xOpJOQcO6cKTGEoRYWn/Z1HPS02lu
oLwrT4TE0DUDqosvo9Z9xLXqxim4rcK21EtY2XrH2QIzxf4m5D0621NJ+iadEliM
IFwlEJ+fb9s1fjWi8pRz2NNgMT5GCKsqUkUYu1xs1XSeajOIVDEmdmOO0MDxGKoc
jeQ+6Oh8tyK2rouHP1CwzYe+s1rgY1QgSq5qoqM19Fuf/yCZunLA/+zEM8QfcOLh
x8H5UA32rrhNfXAQUrOuMewfY3AkamUxpzXfT8xk2gxQBlqdhDrtwJQ7Vr8KKN0W
aDp+03eBqxFCXLMJGdHogigc85COqc5xkzIfYbN58AjE0YON5CEUpduPeQnEBrj7
RbY4KJd59i8akcZoqI61e+KLlN/AZTtkEjGA1fC++EPoPZZM6Pr3f5eHk1QYNGLh
VDSDQCw4/47xjTyUaigakvClkWCrDYFUJUPWBoxqEiyndFLOvs0+kELWSiFLGb9M
FjpXFfDES44Vhg1IW17nY5FHU+3WfdyOFQ9UMSUM1TNayDCJQDIzaMHnojbG00zw
izNh+i9rPb+s4BzW9dICNPqkblGAofP+bP5gEx2fAzTiR1NXYPsCLG/YKWhNZT2r
QQS1xH3y4UAabJzJmTsC8ujnjro8vRm0jCLWpsxzDcTji1FvhGvSgm/WxvYPAAdR
DNoy1+BMVGhOY0t4IRcN5Tp58nGZicjY9T/w99nS07nqYFaALS90MY3fYBpLxVhF
iCh12ImOynPqi5/7vD2oV456OnbvliJ+3Qdnw4n1Ehiqh3TpZeM9pF75761Pj5f9
fkIGNsAxK1tBoHQO/BO1Yjv4z5j6cHsxB+c/2Bx5n1Kzn/pMct1RpZhVte+jW2eU
rS8ZEbEGUoYaDNenuJ+zy6CQrtXK+RwIiK+rSrck04IQlbye9Bhdwg0Lye69UiIV
0ml+s30hAJ21x31edQjdemjYeIV9He4JWERGSIbXxACy0qEDLZYTsauimQ+gvTws
pATybTwYm8r4mMFxAdwEwc+fx+rLGncEW+D8tLUg3IUUircOQoICTikdGPp2DLxz
dsEJnIe0WqtZicev0eVRouIWpAmwQqjiPs6kHMlt/c+jjGW7lmGXEAfplvfyjaWz
Z7tAwZQR18Ma4XvsGjRzjdQcUwno1H+es2QwKfdTMsukI/ZG3ZjrTHCZj0xJ+8ET
SueXvvvGNDjRrJNVKkA5zktNwjczlBZUmWTOgcl/xxXwEkMJaVOQBg/pfrSQB48S
O1jIazkgstWHHLhmAveRK9g+HcpXdRGppEx7/ZNavdXhuXG58LIPKEzrOBCHPNwh
/Rz3jFpPoycvdUUZxU9ye+X3Xp7H5l4B7IUHwlCFk+rWyoIF+Y4W9W4H9A8CheGv
jkEtyGO0KY2iDtO9jzwDq3zZav0IeB7RfL3GGGfrL+ibY6OXY8NHbLnKcb+HQUJj
mIIhkutkVHgtGHLsx3GSqt//wApZVGvFfGiGbAIxZpRjlptKpA4cl2qkgIKCxdtL
71c3zDY5O3v6qQASa/wjWVJ5lehJYmUIwHHR7Vrwu2Gdr4W4mvya6+Lt4uLNFlBr
Jx7xeqgPxRYROU2OOkvQxvsC2HSCFnfOP3jYo3TOkt7OZmnXGJ9/woFepMxfwK7K
Iol6ahpo3I9jnwohXPd7drqxSD35a40pnlftwXsjtXgRAOmDEghtQf+5osdV+TPz
FqEaD/06MilfEenxjz7f7W2Gm8gfLMjbxuFME+KTU08XZqgBvtAh4Oeh2mZNeLSd
JLQKhSQOmj2X6qPVligzTWkJh74s0PI0UwDi2ofLkaRgRvRPIihfwVBBul7Mtunu
owMQMC22ovNup7LSmdBYAxzwD6Ro6v77BccNmIs/F1FebptvI+cHtc0h2igHmc17
8tLXATgr5SUKGlcY85k9UqInrb7ZFBSeIrlZcriK1BAglf9XzLFnSc+NR7w0Av1j
6+RAMiu6Du74szK4mM8cxre2km6aNoVGqJcTe8D9mLlRVKF+Rvox0TUFGp4z+Iy/
5lPXpcNZcWkf4jSWNf4WZt+UQtkiPf0PXw5x4ubhR8a1ZUY85QuGugoMwazHQyqM
sb+ziPPMw/m7P5rWwY9IFFVJlWkztDTzyEULcV/RhHCJQtIRCFzoj7/taxM7v/7s
hQI5I6DK34nxy/9qh8LKx3Q4FDOeWkig9nr9xjxTcUE6ehk0EWXVptapJNCTVgUF
7Az4nFabAyfOo3B6/No9y6l1oRg4vx1XX+VF1JJs43viRAlyBMORbgZRUSH3Y4Da
MVpX2VJi7sjS78TlRg/xK8UZf8gGbQ440kX9iB7xFCKGQWJ+zzezwYh4XHJSf1Tw
Wsjdj7Hq0uAe6urLSs9v4oOsFALerH+0Pt6z4z7g0wy0YsUXS+84oLNCl07/UfJm
4vkg/HpOCCnhIq9Nf720GsBkt5phYry+G2fYM62+lNDlXjOS4Til4HavyztEEN41
Z6BPQIUhJJj9YWVZQYXI6ncJ9+WBLF0hx6Dogu/s40ojCIk9JxuSBjAFfaRdT6mb
2OwW7eiU3lS7IitLtJcwGBJN9ewYZcyk2OBvJueluxUo8oUP0JSCc3EGHFqYBFVM
uARgjE6SvR6GKHSU5NPtsb92tJ6vIGEatEelkQYF8E0T9FJxF4WWRYyx3lsPlE2n
3koR8AON0grMZ36MQ9g3n5DjRUUIVw54AsP+umO0A7Kg2G6wbvYCBd5JnHBT8Adf
kfNklm3YqyL/9qh9FL7XEm1h+vEjlsp1Krqy/0THlxBySsdXSqtDX7AGWkXPq0ir
8tIAuRAvt1cUOUKXuk3SnEFzzZ8wptyvrqWzjpMWOvXP/qRU1zb2F/+nax5P0rsw
p77oANxt5cKZzcKfyWThmLTCwm5EljHxYdhzGwRxyHQZjnt29SmO5RD4hcRT6Blx
e9UUBW2XesiNEuKY9D0bTHFSNxkDk6vFWMQBJjn/KDEG3lcj2zdcnzpJwIvhD8Qr
+ej85dfsFVy+JVPG65sLQ1lDuJm0oWPjyULuwpUgfEKNOAQC6wCLnGfFBRQtaihk
PKN4tyF/86sT1/MiruqlTSsW1L/JHKBmzJUW8nxDcznCHmBQYlJzAlCpIRhtHzU4
gbqJrFjx5OGjGbtFSyXQFROSVqlZSiylZC+BG8hzwLgUbO5AkCaAJIGVhHsdHJ1b
2kFLXuANW5YiVcnH4x7l1YagdgVxZ8QbpP6cU+atIPNNMMRFyjBiSyEVo03EJTrZ
/EELpYxbG1V16+jQXjQFddnjnLQ3D8p+U7WuB9HXXgSI7nZDdKGJrzfa5go0HzPu
9Kg6qxH8zkjKNySpDn8HHbRSnOghIzB00N8ry5L5PY4l3HbYSydQ6KKOJrEiW2YM
MkgSNACgXNNCgvUlXTEnIFE9IwowcBQRrsrlcirweXrBc7xgMicVUwPAGiuz0nko
4BdyxH59aSWRdZWwcTWDm7NmJ2p0YkMIcPzZCn5OcA7zOC83dnAks9pfNSCMNZYz
JGRkOyReqW3acjDWKeaQe1lwNHfEg0Ao73U35puTbo2I+cU5skgMWE2J/ksJub9W
Ji//PEZbimPq2vULFM9u9OO07El6cQXvREf0eYxb3dmZ4bMxWIgUqdiblXhd+e/Y
z98yC+3Jl8E0Oqp9lQ6sqSoNred/yRDDpTdqxxENGf1Tg3MG72YD/LRq9DGTOnOu
lOCbM76ubJaRtf7YpswsCz3Y10SPGwxEEbtYM5uIMrTFsGhsM2FgYFyadEGpB1g9
UU+J6PSZeuSK9Hjl4Mlhd7+BFqzYLc+7Y/lbEUAY0folfmB0d1RssjLzPMsuqrFh
dQgt+0qJKwRfuzQgaK5mio8gCkqNJRYlfZjtVQ8hsIed5b7NacXQkJBLpl5JJ3lW
BWTCiRDJQbcG0hdrUYDblxq25tUGg6K39oPbbbhQRDOsyYFPbmF95WAd1mwsU2NC
OgZIh8J+8NDm+tmzvimF9/GaFx8pNSKc9Se3vS5A0WR+u6zWQCjuOawT5dvC3RD3
e7h0GIukw16RSNH16lXbLwu4Vd1X90vCZgEgw8lcW8isk24VBXCwpa+v9dJVbq//
GjOBgpoB/7vPuguLfL3B4DMXOiH6TjhVed9D+jLuC0Mnl5hdb7SF2QYMeOTqLwMM
RnH/RgPKDKQM3yz4tY60VERJLotpwztjJuRxX7a//LyEgsCaPeoPxzC6wOyC5ozJ
Z7Szvd0VXovPgMUMILPt9C0FYmLAj4OQAqQk1x44ZbG62CQBNYqRg09GDZ98fRyr
QE6q4xMfuOnCoJYqaxdX8T/FmgXjYZ53taqZuKYo30GoUStbSAn8HNp/ycsycBZP
K+n6WF5xB5xyuVRYdiYQOvsxvu8hDlUlXPVEczftMsSqsXLaHMSR1N4IZfk8oWNi
Zj1KnSX40M4zsrJZ/gosPpBErDT21LNNPDRMJRYzh/FuWzMSYG1sckaCRsWcc2my
h5eEudaNdQWpnL7n1/6/NbglBYO9Xujrk/4PL6/lfLpj+3tbD5ycCEOXqZwtcmJE
V1lXiGUz3dN0mTzl8NoSKW7vj+ePEK7BKHL5UfOn7swTHqAi3B9RBAYCDaytJvYk
opnYAEsA2mexXbO9+zmorbLwE9D8TbtcgPSklJ0/nfMLgpafr08FXnRHzioj1+Pk
6vD8k2Em7OAQc2KoBFV/8tH6/0hbsP8bunmJpX5eyxezV9EkHbumf5vmccMHhhhc
lNkLM6tdgBW5hUVSlcHJcYCgGlsxoEl8UBYrP1BX5/ZCwtSIxzDBs9AyiOLWLxKE
h/6usCZW6xr7IoqWY6h9VTRBc3CMi4IDsXE2KUJxIWv2tz+wv1vcZs4wdVFTcUk5
osFidCZ2bzlLBYvkOhDyKU0UTwVA+KGnSFug7EGEutfXvYbE/9j5F1USHR5qzXKG
UUL3oMG5bTCpYL0LtkPHXjvXGBG2eULAIkMzS+PxGk2FCm0Or7A4BHsFc3l9t9BX
ZJXRuIeKmvLXWFDyPem108HyRTVogQWE+aLgGxUvcaMc5Y5+36d6ZWyJZ43g7PLm
QMBQN/0io6Zwi19XJSk9X5UQZq2m8fAMU2rmQuFIl4b2zRs0Dg7vA4Vf+ixZZn0K
ajnbCHyJ9QC4US7Z+3s0cp4HDpiD55TF4XLvVazWDhBId1Clkozhr8JwB8AwLcoF
jiidvll+oeNbYgOAF1Bo2VC31OmZfeMzRr1pYH26zltQrNqEAN5I+8oToGu1KLtb
LXEDnqvkO7KNcjpN6v6yqj9c17sM+JQLzaY5pBZTYVLt4FpfQ2JvQxt9Arwc2tjA
cL0dilqAeLX3Uvrn9h3e8JTNGQWDcwyer989YLl697ZBIpth/bO7otjx7xzDNoUO
3F5YFvaHVFQKFNWaIdzYIuCKWxB/y8XoO+fsjysevsXFEluhj8W9pZGwZPZvBf+M
cfxKwihQRP82KKA+CjbdaRTiTmdPTdQw+G71uoP7oY+4tcsQE33LvoUFvkRR6WUs
U34/vu3lkqtQmZKg8m9PExEnVD0rayAA90OBMzsFIoYYvdGiQNV8D2AKEKUXx0II
PBlHR+yKCgRRt8SKNEzSxksNwDOlsNMqOZ2vqN8+pJDIU05yJoZGuVRE5lHyF6Bx
L5akXoPQ0ogY2WrWGtOzwimzD8r8qFk77oeU34FPX3trcTuJOeRK2Vl8rrTgDHBc
u6cLcWojM8yq9sauLmxNH7EJO1JUawuCRGwYgC4E5GVh7JcYKfW3S4Ve2Yk99BMh
dXu7RxytJ9jG52MfR/0f4XVFjiBvo6rOMgNyOS5Y9Ig4IUuFWN7Yyo9gBPgfeMor
JJ9felcRompdfZSIpfk+5cy869ryQKmjJCiMA71KcDpWLlXvNjWz8MN5ga7C7yZ3
l2kGV8GMDtS1ML9eP4HoXSV6+Y7G7Ty8265KuXMQDoIZ+maSRD3b1MWv8o2HyYUk
I/pVuFpzYZN/k+lYQP6O9r/qOVky/keQu3fnt7lkN/H/BQZvRoWTpNRYou8n9Vp6
ikzgHVHfx13pgTna5eqjZsYzms96vzBgx5dGJMwYGAmPPbeZPajUUBptcvwM7Cq5
t0rHv3GPcX0qZEmtd1f5KaesHzCwXFROctxphrPwj0SeABSDLT9slfj6uf/GJh0y
Iojy1dSubfGevvIP5DyD+iuKyeuTqRtjNPKVs4vFjbgUqJ5NuC8N2Ukt5n/AKxX+
DBncYugkcE2YicTC9iax11bCsXv0lVHMla0XqfDn0HkOU8V0ki8Kk3vupx8vcqXE
nw2T5kIHZf0/5GJ3UwUOQaku4G/P1ZLeeHZXfJMXBHn0bmHq72F8XL8X57f7Xvel
kI9uNIDsCZQ3EilcGSDBvw45GxJguRgEkjXBdF6dioHkZrkABny5C7ABQaOsAv2e
uLMyArPh99vczeBUJ+OLfCb+67NWsUG+Jyfir2kWA13I7xHr5jDrFuvlT34KrpdP
tGtXZz5W2hdYcNSnNp0J0FhC4cnhpDZxd+f08ieUdyEK/aCjqPOh5MJJ+23zeCfn
JGK/wXjOjnAadyieb2juJW+6U42kMpQf2FrgoEltcS9mJ2T6ttUt+dpE3lFXS+jV
8sR7dYQrLCHFwzeSVhFO3oSiKuIUKCQqM0b8MTIL75sd0977mwI2QWPmW/eJ4vPu
7YYymGW0eQkL02O69bRduKshbbZ1JZ+5p9SRxKeWAFhT2CDZ5QxnCI68l10ZjpA3
vVQtSUkck9DeIvkUXrYrFNKVJs5s0iyuRjVXGYObTKwyUUHUPQq+dNikOqjeFrip
BaThP4rxuHHIb7qlI2qOb5BImLmYvOjWP31O+lAM539fCkLOA491zSGfguyQ51jI
cDhBVYqROUgsnhM6xTsLIIGwW0ZLvUKreO780DcDhEeUvI1U6USkB4KGQLFp0uBZ
vAE/4QBSRsplpuhBSt1y7AnBmHT1Pkq0hq1V1vS4T3Z5osvYRf4x4VKVGMv38XNt
YsOyMw8B8XZOMmCdyKFkVfSHqyW/3DmnsELiRkoc+Fq1q4zNwjXmoX1BaUuVd2i1
1HyVk/g8VU91EyP8rjlkTmYFCKhQzFQSXSjD/ly8bIEiwyCFDM79rKBvDdcRRYXr
5jcYaVG27RNwTZxrKOQufQW0B23ZlHjDBvt/ulEqXBLVU+L46fD6CR5DxPNclySL
U1yjXFf/2CqhB1SurOI/cFigbN7BkriLjwYa9JN0T7pL+4ceMydQWyHzUtvBsrdS
9BsTnz9GX0rO7akXWuC+qmKCe7yk5jLOSjGFzwcx/vkIlngDv4YO8fJPJBEQxuON
eg2GjeZVpPiKD4bNNH4sxqHqTkUEp4MTZwFKlKAyT0IfA+Qg3DhGA3JM+iSVNrcW
606SznOAkXNP54M1VIYUd2ytKEVWiUneouW6wUnMNbQKVd7Y/CgJsTWBiRy00Tm3
hntDZMHbA8YYjG6JQl0dqt7h2VQGfiqa8jws9r1EwhhdEvTbYn+7luPyTvAbHgvb
7fqsVm3Kz69cL1WFPRecFyIipAdP+CPgYuZoAr6G+XH3A7gCtkdvW3gHgZy3ds7X
cTo5MdbEqLbgnz9LG1xq7lcdus9llQQMH2sfQh6TtSyiO+jdlJGrPsYRfw5koKPo
y4OEuGJamB9nTxxaBIok2z45t2iPL8jtFyj0XVnLkDkgMG90fW6XngnBkrVgLIvi
ygKd7DiaaGD+IbMHc4KjrlbnUsxqn0KHAb9eWILWOU9Qx3TYPUQfTXc0fh5GrQbN
gR6cnnJOtaosJ0cC4YRoUvV06A/ENTLGZQCep2MHSSv80A39M3cw72oU/CRJGHiU
6LgKzTA5F2+2n5ShjrNcRcLKeIilCXgAGGZSC/06dF2+1tcpJ2Tpj4KZZ8PhOHjM
a9Rg1tiqKxjwGIYSts92jFF7kGn0NdGn7jzFffgU8gyePWk7EJvVz4U7WgvRwr1D
Vexk8oTp22vYeCCqx77imeiEyYg4JIzot4T03YxEPhJnrgPsE702yMSCZ5XVccfS
zJL+2mxR1Qv/ggt6V03unl/CtbJEYmB8ePT6utHJVFy8VmL7DSOPCxPd32Xerw0v
yxskMuvgjj7Ua4gVt4gHyJ6fQuztmVB4blZjhbQ5UfPg3NZ3Cdd+EF8JwxF3SYuP
3be8XnNS00N9VU9Po3z9AdGGjs4fez8/3iHgOHhHUmnsid8DHuC57XF7JpsfTwHI
BqO4DYQy9lLifntKiT5eh+RqraQF8AxOTX0rtfij8Bos5z7wxP/YImUQow46yliS
pECjzt26ZHep8tL5/njJc9cce8/SX6ppVDL1y33RUyclQVk2+H3GWh7XKo1RoTP4
4TZca23oaQMcuumKWIX9HgfZLirSXKP4KRZVVfb8wjzso7tZOnITs4pO+7Dc/U4j
Z7GNrGNJpL+QMWYxfWuvuEz3r2Le15bjKaDsKAH5prpIXbmraUC0kKNhT6EERPQl
/4ssdmvmjga8tfZPeFSpjNjhJSIeWkxe1BohcD8xaXy8qDAdaOMUwc8g6NPml6E6
AzcCr4nc/RA3eu3N91/hHIEfKbsfnrnFCqkMDS0eXc8jXQRfU2yj7eUM9BZMJaua
FBS1YZivJc6rEZc6afJtpuCTwH+lW1pgAMIm0ZIcDtKNwBJbjspC+LXCAJN81FzJ
7mIrCLuFWe0JtWj54M1QRR2UXPtgDZ+M9mWtRuNwqHI1G0VyVXyBR8oyKR7sZ/3h
hjX8weglJjFXFr3EogbiS3m2LofKBkoA/1oGFNuKIsM1MorQYFPzQgugHhveBCau
wiFgpPuTb/TIrHNSeChdPmZvN8nBTCPntxr1xYTn0C6Wv9gAe9UD+ZaW320A8+cO
WuhJnljf3LEOwlbXmIL6F6XgqKPo2DYX1GjN9BkuMhdY65jxCb41ANi0XA7LI9H8
nd8UFLhAD2Q8iNgbUNByaJ2/lLi5I535AFzf24XTPZzK/+hWMJqWtKmJZXZOjNpn
tNfYqm2Bq3Bujgv7pqsB+ghaQiU2emk04QPnTue62tbGXbr0RiVyCVQNrUfk9pVZ
83RbcTaxRPZWgU77Ab7eE7ym/vj60WmwXBakV/KAwqgbwT+1E3TTBjKo0nDr8BzI
03g7fSDrOT2RMGikRzyIuJdn3wUjrzHv73XXzjDroNcp+tKMfMLLkW/VQXK/HLyT
2LlmFCJuOc46SFLPHqmIpOHgC/+iC6BCW1cudG4AADoAsGOp7F/uYuy2aet6+ut/
BAQ1eNhxCbNVLt8jC2Wpv4x3dxld0J5g0CaH7mvCrueaOs+aN/mpygLvoRMQ3px3
DNp/yU7HVq7S0WL7E+xXfPmbTpKx4iktqdKqRpOty50EIm5ew4OMir5RlVfPtbI9
XA0UCUrVCh1UMBMUXbcJtQC824JtYH/dY5yBvIX46VIuEPyQ12JWf6L4KHfflpZ5
Qlv6KBzp1dnn6CLRvfAqtXqhyIE71chWgczu1+BShD41nIh8bEv+5r3cQYoLkElG
i6dtfIQbAcFPm/PSHd0xPzJUqq9KkpfVM6LMbDlQbnVx3codbrYHZPe7FvVQ0G/5
F1QWhg7DnV5JJk4/VyK5WM52+iep4gccazOQrZqKzLhCi6oSMI3SlaoJLREXbd0C
CqYnTZuqZxPRtkUW2rqLif/OqAgKJxclvr7K3PXPzltBToIKZ/b6my6L2T8ibM/o
x0M5ULPSI54iVCyCZGZAXGMtMJtSOqfnmhnCOBjluUBloWjozguHNkH81ZA1d+Hb
/lvJFFrJvnCXdP5hg7Qn4mh8kirQZHq/9e4rqTm2lXpqwCrcn4caDgUm0e4r/Hpg
wBEUC6pjvHPvVspeLd4zmYq6HQArBwo3gsDOvwbjOpIZJ66FD0VBv/VTlE0mTyQ1
LqEsAuZQAdZ3nYltKP6jtQT0AUdK2HfJXHysWUzWkSpQx5w8O5nF56YMAzYzSCjC
Og5kA+m7fslY38BjkZLVs+qohL3krGB1jxoarF1bNDfwRmbZmXKu0E1W/PllWWlP
2gF33JEfWmmWmQGEtFvBL1sC6AOmjlx8gzExG4OJ3qiFKuEFGdqhFVN1vgolux2D
usJzleDuGYqOl8BpeDK5Yf47kR9EeGmyM4h5WsNWLjLLwLMxAN9CrrvgbudBUrJ+
7cgBfIs7UXsK8N9Musuu89JSGc8zZiGQVOcpkrgTH3UT04q0EMxcZw3vA580piR3
NFx01sIzTEBDy8LJ0veN4Dw3zES/SxagnMH96TaxSLGD7Ck3XukBpbJAK+/axbRn
cutn81mohCNjM+uCS+bc1kfaC/4k0dJfzVy8zbPdNd61Hj1L++KVR41J/dGTEOQw
btX7gTjlhciPVyA4shw4cpkjgK8MW0rEJ2LczbQC57Ny95aPSri4bz8I7dyqYedN
eFnQ3gfJSLY/YcfN8CAulffI8BH8I93NJzP9+EhXt8YuPmURlFuTx595W7xiqIEY
Ko9rV+t8HJxRFYz1omjkEsEq8AvTC9SUiayFhDcF/XZvxkI+JDpQlQRVVtibEjvh
CiD3ZQW6RQGnTsSSM208i/aOOw/ZMu+CoHAd3uapfeXF9EN2fj4qST+jMsXSDXFE
N8pXrgsLfktYa9mmr+Sg73Qu9aUM7X4IQkQR1neTDMbjTs7tV+/yyWoyrGljvIsF
wGTjFRde2vkop34/2OA2HNb/HGs3Yz6c1TZLonvgCUwOxb2Xb7lrrfdQkXe1TTUQ
TyI6DB2N/myjMFgyNnXOAN99QY2XzQyRI2cGoKDYTpzK+x9PsndaAnzPv6xDq+qo
bjwsprR/MJEM9Jln7dfyxjQxo3nBZGvsRxSDnASdkZQyEvGMdE1fO+KaPZAJbss2
Hvfpdva8JWeba//1I1WzE0oexjW82qujBpNkosyM6063FjvJYUQgD/IVkYfJC6Zy
GfftjBTZmuoAPvLx3vjMSCp9PntQCCX2RPfo8sHhU0qIvd2dznc3v83ct2miL00E
4M4pYpvB0Ul48GUSNuMf5dcAp4jQQ8hD66PO4cQtXnpX0VXupWS3yxIaY0H+Hi73
1XpBeOB+24szHPLmV6sPTc/nX50VlzcsUu8N2112EoHmen9YdOaDA9i7pHtHCBXR
i+bNUNB9T2+AzcjGniysRl1y8qtf6iqiSBn2e6f0/ZNaX6cVactaokrBeenu91c3
c/aqG7ht09tPL93DVkACPVURC0CvbRB12KRPNl27E44fBlBWiTsMTEaN8lgCYJfq
l2Lh9mbiYzAlGhsWHcP0qNflfli2i22xF0NLTR2XK/Z3PsPi0cExtHtNZ/jblfyT
cyBU7h6k6UTYoflORYJdGLPahNqh6tXjFd4D3Uc+rNvJwHhsbJ8WUq5KG1I4TakV
J91cofDbHv130JPV+2rOa49xLKFGnxaYaY8gTcrK77cGu7oow9H8kFRhycNhFf1/
E0zmBgn9v3oNnoOM+dcSqLPspS/y85AUPrwsnvqi8Ae+QaVyt5buzTm0WtQNN8Cu
kI4VC40oKbwBkdAJyYx3D95xdw/lZh/UU6K9y6i6uy0Rnz+gnS+U3I3ibXvBajm+
XHqb7i6/MzQy5aGpxkeOJi2s6zwbkcKnJJo3/iisBNO8FhnIyuGHK6ehARMz2HcQ
q7PRX5y1d3Cc4Q7Qhx87SgARvicyUop889YtgGqzhT0B+LQmxPne7BgN6M94HieE
VXN1MDrurZfanOi91hsKMPr/dH8cNGbbTkdI/2F+aqkYVjDLs+7UDrjWX71y40H5
9SS0W8rgSzb6fJIITXP19Id2lBaMzEI+j0AMWaqCDHl6hgxxGTnHXZ80e+hmrWmU
l2ZVQbvrOIdU7pRjP/DnzowEjaFwAAdmzQZ+vY/yCRIWKd+Wa5IK8wcRjVukg8+9
Fqu3vH5dcSB/EKPhG7X5tZrX3q+CnzPJisThiL0ydFvmG0dFIFESkfmxF9W3Yxv5
ZGW6Os5pma4Ovhm2MB8GcIOvmzcU8hGOAY21EoXAYOr7I1TIXNHXWQn7VzGt7gmF
aIn8g1J7lBFOs0luewAgXdyKiumWr7N3lM883iceyhvSswpLPTublMmnbVSH0+3b
TI2+4gQNb1uvRDCpvd5FpZnwNThzzkSmvYoGJi4XTb/HmpoMO5GhF2waS5cVOBmN
goWMwly3C3LAsKO8i9YcyKleVrWuydK4vr1fY9EZEQJAAMSUAeEwynx2x36Dn51C
MqcWSPSXJSa4Y/OJW/CT45L1cMqdW2b4AmbX+BGd5HRhI/FhemLkma0Xz+iD47dN
kkvNTfTR/Op6+mqCuyNuaSKeFF2fvfir5CibnGUbO4uCkbkzqxH4nknUi5mD/LdL
Yhjd/F/tunPfLr3s5//stMXvN2FOF7YskhnT7W6TuvOlUoQ5QoZ36eztw0WZfEta
nAR27eRQgZdXbAxmBHUCW0gZll+UU6CAsTj57TASkP40fjh9HBm0dHCXhofgbMNC
0NvIYFiVIbWuKd5WXDQHrqf/loc8h8Ahw2Ecq0C26TrR/XEVgexZzjAtugxvOucO
5itba6+sqqls77YdKvsDe+QqTcmL6ctqwl+meCPS9ukRrwqZSn8YYGKlvGY7MVdz
zsTLSNSRq4iRPEkl7Ld2F/nhLv0u0tu5TB1buz4sbmTUAD8/eXjmtHikMxfr9Buj
za9Eh60q9QvP66Yzcgk7JXASNOqzQBRtAuQ4QvmJtGkZCw9EkE+TgNKlfNdnGvqu
Utn97Di88WmFT3iNGStpzOt5STBQWrJsiro9Bi4OqrmSB35N/S2hefmUji1kx17b
mVPZHQzpptUMNpQhq832tlmM3CtWoDRZN7SDL4QTDSOK1pE4uE495VQSHbAKjdX1
WgBM/KuLTxH3ec83d6iGmAE5YhR7drHAcRah2+yPJAqkHmrV2a82jJHKqdgXltY1
62OfTvwIVqXXowtvGBhhczUlFnh6sHviU75UyFoL0YeWznjCxLppwjPbTTEd4y9t
M0fBcDn8LwluYJFIz/1RZ4JC62AJwMKhCov47nfWX2djDd/XlDKCmJU4VXRGvSLV
aV6AIDF3porYpX5eRMFpP17dlOAWmJZZwccKcuwrqh+bOJ1LrxEh8KyYhWfv++2P
mB+rE9tZB++rn4DJOxJOohOZvFIu1cxf4A5PVG0gyFoUuhke7KnrZ00E+YM6U01h
TiPUhsPo9joLFjr8I18NL2Md9F4SB1Wc2K/UXeMNIbiyZlc7tNzM3EJRV+pHNJY1
GMa2EC6xrZnZaCHufdO2iXq2pBo03l6mHhz3OmBITMPVsuouQu2enOqYX4kpdFjc
GburnNqBXLZhCtBt2dTV1raXFQFZDgMFNzV+FLAqF5ITybs5irXUZHB69ht9Otil
mRNEXWAnHQIS9TD80rRfOQUa77Rtm+qfaKp/3QYhT9Us/l9fmokxmLLbbKlF2OXU
VVqjl+7IbfAr7efOBoMdh+HwZPDK6qKwBAB/lXFkmrFR60czZGVVgBvE4YCYNmdD
ifL9h7eqfJ4PyV49//f+no3lpHraQguph52+ClzdjwU9jheKfzoDY4Txh+yF34u5
wWUtsNIzK3OQWIIr5N17jjOJTC+se3USRpbD0evYjvrOEMYt6xnk5LLAR2NPoTcM
dHkg882q71LeftdGpJG5jhHVIRFOKLhah7Lpkgo/Jgilsum+h5//6oGAMfj87DPR
QnH8a5OKAcqXd6FH/6BeaHErqQsVS1qOihL5qITUgsydGQlrB/TbABscI5JWUSVR
Thsf1yhTPcm+tkPBIkezWZ79baHpqV1z3dMUPC5ppVCCVNokhrGRs3UwfSEuJd12
gVIYuoCyJAvVfjcFIvZ0eHFzS/lObnnW4VygeyxL/PLRnVKcsqP+uXymwmpRMPDG
l2oc2JNBG+FmkGdcSBKxb4wd1Vg8zAXu3ZZ1L1za6H0edvMdpWn73N3SLt9IGqDB
X6jrHs+YJT3m9Fin5Y6QI3QKU9pJL1RvYIzOkUX5o0hgLA4vKqjzz+c1Bnr7rgP8
Low2srnYI0nPxIQENqUv66amo+DXDYu4/IGwUgI3g9jJsvxmWHd1FkXfgI0Pd3bv
MSruDGcmOK1h4u7yb28sqWkNLSVMc2xuInwsQPoh+yPP/HbMsg+WdWjabzk8GjIC
t1PGk4cTX/6XigULvh86uvkzdSEkJJL0vw5OBabovBaCkxkY1Dm5jD7yHlXuN5ts
lntvEdNWJM3ejBfXqOKVixpR5Mxf4hAt2Bo+hOFSE8xOgEKxZWR6xXjK7U+b4f5H
0Mahvdbq0JAHtDfmJic2BpE3PPpqFl/EO77a35nmfVquTH+HWrTKJabhBT7empk+
3LQQMBv8TmSS6pQmAiz1epNShygcwvEWX6wcChT1HV/3rINL3dFWgSquFcFfcNDN
amzqHMrLcb+yVOKH4EzyLYpD7eq07onhoRsDIiWHPduCrfpEMxkJWdgQ2Xz2KQtP
Aa/eqqDgrpOtyfgRwsVTG6HsGPTL2cHP8uOzflYt5jHBO02EW2kW3x7WtmA8wj6i
6cBYXjfNVC1rhTL32sSHxEBe5hHc18WXfoL6fCaNbRjJO/9ZV+kDsU5QnLsGjdTj
Xr5Ehlu+s/c9zCWBrDvTJfr2RMCaGY3j6/uNIQ8s6Vfy24nVbA6TCrQmQvvKXxBQ
M44nJkCZywT3ynyrYxad7ZSowheyBk5xEA+MHHzkDV9qz//ymCUmaCWMUpK91QYk
bxzx4G26dmX2HZbKsE6NojeaqnEykgcpDGOy5cczmP1Uv9sl6vD5CmxWw5qGYcWt
1P7H7bSD3hOfsI16MCVo7FS8xJocAFh/04EPERHWD3AfhQ1UqakyQPjNLV9DnyR2
55fuYf/Eo/pdQseT31MBxKQ1CfRlmcbexWx0fCJUwT3bGyfWv0RgKzcSEN7ttB9q
KOGsIiRKX8aRVfc3Yq4AmITIVxbHXQkmz1bLqx+32Owrx7O/qCK/kr5k0IX4hJ3Y
6C7/ir6bC3FeslAqzZjcFN9hIsBTR7poo0AJHzBXpY/KBosTnc7WN7xmkbOkOK+O
vZC0QrB7wpOcrKSegxO4B65CT794MLCpkV9zIT7TZYunsYbREjyv3La9CETOdL+n
EIzrAjwOMlZsTd+oIXZPEuqGMlhW3E1+k4wX8enUCsthJNp/IHHEvqyIrf3XsdUg
SqgvyYLouluXEsfgDAjOECfWSz44Ce7lA0eDQo4Lg6CzCzTWR0Oke39yULted0R9
PngV5qAPCVZ9U6sHnuQLQLj+0HioDapvIkggIYxH+iMixYyBCkVRf+lxGgewe4f9
Lj8/D3aDi1s1qHw13zlTljGwWw11QyBeBV2d71iBkR2LKQ9gf3UKyYkEAbepqWHP
hSiX/L5jbM9DtPzF63LTT2ZcgRnNh+mjHn90qIahP1ZuNCSQ4N95KHllx0eSotgK
AMqb9opav6B6fpbCjFcy4ujsVnVjoanMa7MOtpXg7ywDrmL1Xeaj8oCz8uTm/3oN
L4LTxK0UAcuvhqhMi8XBVvr99fj3uX5HeSSycQYiRG9Wz7yMC0znXtLvmanCX/qu
85reGUlN5rA3gkbt1CMZiKkpYcOSX8dD5HTddz5G8o64v8uMpYFpSxkAJvEFiuc9
0ceS+AQVt5vGW5gWjkeMxsqs+w9W4Zghama2lbLN1lQFY6f+8GbtSefxH1NxjpX9
66PLqLNtbhAi76/PuHdWpFymmRPPB7nYf4i3oB9teh2EPs8LLNICt7JP7QOzDC9F
Pk7r11XaWVdOXgMc4Ej7geNxwWYSh80cWZMcZtb1yzt9oszCn6hRFiz/i2Sw9UYC
hsRtJf7bhG3E1poHtwUwctXGpm8hQAX5AtT5mtRXE9abIU6niftwJPwaOv/WEtWI
2+8pKD/j8mJA/WQ2aDaGBWng43Q2rv+RsNUJuZbRQCBsQF4d7OqBGEn+BOD6DAF/
jLNfVHDmiSNaQRnncgBmvTGdb8RgALIP8dremawV0zj88vy43KRBxHds3pSnjCWS
0Ib2iBpQqEvVbGV34Z2ho0/NezbrkpXzN819pvQLIshzW3D0qVVtYaZ8kbyAbKr8
4vRjDjgecBx/PEnQ4x2U2x63NG2joy7BZ98pue6jZMAyuQEAEFh9MDWovjr9ELm4
2D2xRrb0glNVkWlHlbZZgcMMjJS8ZF5yEppKZ3OmRrteJoDXjiJBkWZTqc++wofS
7fbdH65erAjmDNQt6AAPr5lsGsS6u98jKkeZK3I4tkr0WQvJSZaFS4qu5H7WaJo4
9U8h5f/Um8AEtMsUdzmiD0JV1BgQG3pehOfKz/XTBrVPDyaab7gw84UpLXQvtv6r
xKlEc2ncgBx6TbfcFdEU7fXJoH+SS/2taPqA8zEYHFrLg8ThBlsPhKrjY5Kv65VI
UAzwQU340G5sgqic6RZ9HUdBJJo+Ea8LZjWEilqJa6g4UoBB5X6WOXpzd/2ayWD0
0a6zQ3/05qDqe/HURYapCniU7zEHa4tYLSbU/JLTIs+WZR9TjpsTgRC/lyaVnbN5
9/ifHBlZ4Fnq/BGaXL5dHLXu7+ZoB0IMo0DRiSSUilfB5tABhlzUVejQPPbxUiej
ZNskAYJyOFGH6AtG8fz3HOFTJvlyC6XU1m7zidEdRk0NOMHmjR+TIPy4YsV2CcFd
toXcdzdajB+1A66nhcICbM7Y3HPrhzNhrLQTzefhte9+ib6DWqvB3YuyD0F5h1Xb
xVqpy+UJLDNpyCKWa1vc+7p6D4fleBo6bZENzEv1oe6iFIP7AzYAb7XX8fKUjdnI
a/3fMa2xb4ylmcV88dIouWJlNzdtplYXzL1EmBRS8j0Iad8XvagdGIwwQ1vTuWkC
Tio9qGvQDgRepm43JubdzfjkkcMS8+2O34KkC9rXvPA5ogSWwzGJG6trju/3yKHq
2FwPIadEocjGkp7+zO9qSu8J2thbOfIQtTq3m0bAg+4RSRNREIMThmdECrv2OIvx
jbLoa5TNcxR7wqBcNyD6aR/7GJKknm1X1/tDq9nZHhTGFBen5DbaIf5AUvLYIrR0
Jzohu5bZzFZGR/bMn7MYQx9RtNoQEnJzDv58UJMN+aLuXTHfi2hCUjsi7fPC5woX
bQr/x77f/1R+cQUg27v8o+e7FzoNVZUPJVRjX0r8tdOEozkyCaQ/sm4pnpBpPajr
CwhNtfWYkyGliQOfceULtoC1XEyBHyXJ8ub7hLEDB7w6KcNNrNzuyBPVeshsIMhw
HtJ+U5R7gKhjs3mioxdLhT1O5zu0houfBmV/tV02X3GBEpjdrxv96Q0YwzMla842
r1R2AvCGXojslhABHrH9UEL7w0OK0pnS4TOtBbnJwy7mOjRvO65QwL3FgFg73PeV
TJivIT7nlCV67f6wyiUM3Tltbg9otWCujHnWV7lMbzeIgYfstlzH9H0t4Sl38uhg
Q8oEZUotMkmcVStJIIgNe3jZ/5RPoO0BPU9CeSBrayAilVq8ZcpFcUpSa2ytflN9
GAqs2TXY0jly4yi1opDRrg0Ti2SEfwzd5zEzqZKuCpi1aISve0w93h2ozePj2Jxx
nh4m/k4/YIpm/F+lHxtk8j/qepAFIKCf6hdHPitYclB9bfrRAORQxoFiu5Wkq+Wx
vKbVVceSey5xkat0ioHjuAw/vmEACTYTCZwH541Vqpo1xBJ7MgRP0V0/TxGlxLjO
mTjY5uOh81Z7nWrnDXEg++0GzL+AY845vOq74u7vs5peJn33qifstxxGkO0TXwd0
lzwQwG+U8rxWZ9SYNGdgFFq+0bhJK1cZl6IMuDMcmvZAuFJWop8qPuoDeJrCk8Lv
YH13BKpF5i3F8+NYtmRW6enF4adh4fMlufttXO7+n5IzPZcVMyxd/aqTWYu8vP3h
TYAcJc87WlRFVUsYKbbp4f6P4KXzWqJaYc993l7dFehGjLoaD68AS4JgTHNSQuKs
KsEnghVgcChz3yHJdtKGuCwVDVRCvi0Ier+odB9snjiZr2Zt0QDBk6z2fzcmpgCO
6mV5Uhcbkx3TweePB2I8qyLahDUEi1/y0LdvF9Yis7Wlxgv7Ns24fj2LAZZpIkiR
t9lFXqQNFR9zkEQLX8EMe5e4XvrCN0ZKkYLi3dQdwxGF7u0ccJDDYIxznt3nDoB+
F/b07Z5LtFPFBhvnbN11TNCGCKTRmIaFI6/iK+NwEWlorf/TFoFx8NMVDxbpUs4q
SwEWpqz/sZpRlYqwDl/xG1qmBnGeVGCnmcKooUyo9HobCFeXI/TCqRcGpuIw2joQ
hI/z9ejovH0RAJpyK1jFIaqLES6URgQS4ZjxEg/QDRiydeIUVaXOz7XFaxA9yeqm
o2pVBx3GCOPh0yxItoptsJxsQxOKpB2QKzJl9n82dwlEpM+2NM2FfAElkhALBCgA
afwsIAmTvcEa1m+kP7y39xAVqfqsNvgbhHSr+zG1u3cDQPkyiBXeeywl18d5jraG
2dfF30qsnVHlyLX7EElhZkHeo3sUIk5wAo6GexTluZQ4/sVjQgExRboWLWd3EYkk
6PhdBkwmCvQQTbmnswv5cI//djfSduwN7eURPAo2pheySQAo7q4Nv/+hgvBiT3fw
eVsedKChoFDZsXjJgr2JJRpFS1vN3AzLGjw/+EFTV+6RkXDHiEkJvtkYdBYwtB0K
LLT2uqQ+W6vLzCMfj6klD+2CUfdlVtcwJvMYDoasMj+4BDJb+wNO0rJLkOtFPQNq
SJO3+vZk1AACvzt/633Vcc7Uy6JjYzj3xskKuEirsRy12HSDV+NrQa1YskC9wt4c
lrI+2XtkXX0on7E+5kpwD6iircg962nyec8g5YBHPmiJNKUEA7HOGolcYaeEnmx0
BpYYxyJq6CyTIxwTP5da9izgBR79szoR2JA5jCw5d0E+fRtW62visEW1/WCBrWbs
Xu4UdLzEb9rsnmsw8zhM6SV0qwiBFVHEJLabmXI03iLEU0WOfmMxXzHiIMhNER/W
8cYHfqvC3Qjt2KupCwIUHNwHbWcMnAq3KHYTnhcW4tvhauigA51VNcbNwpb20w9y
DBfPmphgiMDfNX9QALOtftLSav9EEbSM+tTkSLqyzouTYAwTOuMnqNYBEaT0KBvi
+BqL+B5hhyNxU6zpU6j3H49x2RuH0w1sIpI/PlO6sIeDPjByQqNYEW636jUh2Obd
60dfhYxFFeiyHF+cRR/Gq3eyXM1W0/VCe77q8E1DOAZ20AX32qDwE7+quMHCpd6K
KZkWfv92kGZaU4cj0fy48h4h14Z1OR+1s62RFdKbfhnYT4M0KjWonV1Nn8E9rpKv
fxnl9tJdIiMoVNgEMxMmUVf5NNVbGEUq2HpVAuQPiPtS1BGrltgF9ms1iNSjdw8I
njl7VhHpE7Y0WbSXMEHLR+C20L2khu4p34wTeaqnNjD4sd8/s1vO2vd8urVoQ2ye
Co5bI7pOMg7L1jObP3Bq++30I/atqAWFzEdPwCPpsk6XlKai2+eCSIyDgvFWx4tD
Jy1ZXgVWzxSaSRIeVJ6S8TbjJZrXpDwkOhPPwOvoE2VLibSLaBVDUtRbdj0Ni7Xc
KQYIpKM/sbE7lHLKEFQ5eVOWAf3J5MFvU4m2LjbEnSrZmnhe43a4lpkDJ8XWBSMe
PQDrGX1NUE3J4TikJ4RZGsgJ4Nq3WRQkwEzDgDsopcVPb2XeiMu762RQXDP4dEYD
fo/rtQCvxzzWfMlBHEoX0MAtbxZMRPTtfAEhun4Pi87NtL6rBTfzDG+UyoGIDx5Z
xNLran/kXTfTk19PFuIssbNVlg+lzGxXI9ZPnSUJT5hrg9QrO2Lj/u423ZGmIa3N
hGtpG8MV856EXwFsbNYKSw8f9Ha7FZSd+TCKCFPx/xL2xOCd49pl8ywXQ0oxSb1r
fqyIlxFWrZK6ygg6P3myNDkjJNHW/o7r8OAV4s/gBUPupmZYpcC1NRm8qvP5eSUQ
kfn9MsrrellL7T3QrjGApvdywOyAUlzzYB1d7cG1gv4UsyKKHDDrmuZunhQjGI2r
L01T6cPWVJEdybbElj/XNzgVmmOYzNGmCsZJeRSof+ZsBYEjT9+qpn0MhOH2VT4I
smrxv3cH7o6Ec5bVxR9rxBkV7bS8Ntx24Nnta1A0l3ZoVJZjvbiHYBxEBz9GhfSn
yBHd3xv6U3q9/mBgbBJOYwzkc5tMTq/snqtmJ+ieTHN6uqtsDSeKL/BbyL4a5PKw
mjJbJ3Bq/1401dEWmECLFt0hwCE9E96U61ZFMckKnboalkyTV6ebcWBGccR0qdFK
X9sYMCrtfxr0DJ0fDA9Kpyge7n/2bFX/tUofj/B9ukc0xc5pWPrhUglNfH43NwWN
k1tTtX0P8TtP6OwDq3vq/BGyU/zNfgc+ZrwregtPFuIpBP29Yb48DQE7kTwFLqZY
hMHJm3PY7/NUhyoPslpTDNo/1hngaAeAOLFmCvrnRJl1wb2A9OKCFl8SEnylTCW7
vCTwQiGkSluABDjxKoGFqsZsxxE+oUKkvv8f+1fmXbWD80s8rlS/ZV6VDxANSMUW
DUbfu/wYw4Eu9GqpKZRfkitF6iYWjmD0vLORGmRnvA41RHhCkl85TQgMEZQ0RQz2
k8saNKHQe2cvbSKYiOtoJSMpNj83RhM6Quy68sNr4rTmXWUl4ovBpH1Mz6/IJiEe
s6rcpcXbuFUJvftuiKFG9X+thoejq6pxjSGTLQlPvROslsLXhwFQK5NwyrGlpDfU
e6FWy+dcWk+sIdPzeqKSGmLROn5kE0wHBGasOMFORFgimfwgChwg+aiT1Cfgduwh
7ZgaFMu1Hgldrx9xhhu3mKN0gnMwis/pTyrlYGHPm2YQONYVTRBwZ6Zn6YVdOYwK
rr0H7X0H3Q6eFQsF54Ad5AG5lnL3s+dAGShCZdwae09St6/8C0cmzZcw12FIkhLW
gm0Gul1NhD6IHPQXXNzyFpc7P1gDV+U5izhtpMg/0iqgSZ7w8bTnBcbstUBZP6jk
Ii2macr3Ik3/JKd/jBUK/czdQxJ5J1YmXDDK8I46MMBbHwe2FGI7GtspkcwO3K8D
r3XPZZAUUbaUoJk+Ag9JmI+21LQoMtRzdKAxSTUgtVs8rZHkbq7Q5PGedi0XO4u6
8cCOjNAwsG60EA31+B3lSoQcll/Wm4wWRaZ8GQ7Z/5sP8h6GVC3GNfkNPYCQZ4p6
+ZRuMUo96Mmj4mTFz7Y4mneDcypXNhAoYCLVW766uJ5qBzfgtmUm+A8WlL5b0tiL
S0a0H9JCJfpQGjNjtNAwUJtT6muT/Ts7RDogpsX61GIaltAOGK2a0iLHq7L5kJ0V
eerzY/MmyvQUCa5sHpqx9Dq4EL35Rsych5kO6cqaLqJIHfRC0uNIOKiwHPdVKmWP
L9rlj0qIUN+WJ66gqXuGB1v7sKS7bujomrf95bFVaRZCZq2X8iG3mTGeWvnBBMeH
avIcX+Tj1FmctwMFzJXjYuMXiRlQmHkn8LsrfwKwIWmrg7Gk2l6TqMFIYjtbojVr
BQATQFqVtUJcc6bMqt4YbtJz7AV4Bva2U07fHvdlxhuGyjERducOCF9qMVdkQb9a
j2zxRK1U8GzxLNw3H37mq+/mQqnxll/DrtyCT+tKxP+8VUjFbZG7xo6J79/uxXh4
2+sytAW7dPj2KSAbGy7tQybrYxZsxh0NyhznrY2MCkIQbA4dYAg3pLVXWobjpyvI
1I09epLHukXIbMiY0W3wIauTdYByi+n03AFEnfIfHrxduknsfUPNynKojD1SgJMg
dfMJUd71E8gT5PH4BEkbzx2DdIhlGWmBE+OPK6A6MbS16XxIP1BN8EUabHkdEs1c
t64lsjj1m8ozo8GQ7yRCXR8Dvln1ffqX+aN3iER566epgun4j8cz6SYINesWaC7T
fh94StffmSbmtcWhzd6lALLCUusL+z2llaUyhTfWM7etntZ+LQcREKVZCsd/rbwj
1/KBiRPyca6bbd/JWqWCvQ5KyvdR8L6wVHM2y0LJ+pIQEErNzqP91Z0bv+oLBMG6
zvilhVKya96HKdoNDoHs8lEdulTjy0iVPy4XKsEwCmlbGrzdx+/Vvt9caFi+wFuw
zO7cXCamEv7CijisTbintEoOEqIAiS2uNbBi7SLItYCiqrwcldUP6vzW2mKp8w8l
RxBk/6ADANYzLFy2SXDZgaJ0bbtWtnPWI4KZv7kzes3wrqvDieT1VpRaFyaaIBnT
kkf3NH6pheii9ZDUWKGv9vyU95pMpR9wGA7jSaV6ice26mo98Gx634PGPOgYMbli
lTAYdyWt//aM15F5SetN7r0zzhuqM/tQDPvEsVxR98EKen2nYJh9G41gSDWhtxDQ
T7QxJG8/8y+W9JCwnCVl2H9oOs31iSPOcvSzJDB3HHV2fV+sSEApZqivUwx/5n/g
ZkBWglrSWH8EcxpJ+C3q0JrDj1qPJMklP7gCgzSkjKIiJjBy2+Cec3PWDChWRocp
CNnHJElvP4qZxv5fi2ELU1tfFnYUw7MzWX60snA8q7n/k2vnPPsHLwfB7A4lBkHY
XqgQtLb3yz1bDWT5RQxySB78uSZoR8XW5DY8bcc4oXtDIRM79kEBSUQJDWYCMglR
Cjixhw95kLREY5CGQh8Ho85EATZE/YvzAo4SnFWQmYn7gvtR0W569OIoDFtn9OSo
wVmdjmGRxhsAfkRHpDhuxpk/vN5q5ASafCyg5QxCYf4uZZ9SivKXrL8om6jI4pt3
FCJnGYDuiHvxaWRXdjkLyKuwMNtmacihMigZ6R8FDKUjPCOKZz0z9+vHk/w5puZ7
KvBSxsM+9JLGT36+jlBTTZ1DmOmI+rnJByeRddILSE9+XTuridJkS8uMpAJBwTRZ
UlqgP4/357IT5wvnVwqJQSFv77CLAqJFMMYJfn9jmrR1KanRzGZmaVFWDbruKBVW
Kr5HVX0z8g9wFmxNQKv8kAUkYcr3al9+cIzI0yRpSvtP/W7N5fzIKWJXYZYf+EhS
VtdkEynww6tCapsrKG3OKCyYK24bXC1O7LIY0I/k1pzvcNwnVbhsOmKNy9aB6PgH
3tlgoRT4l/K6DWCYlr3yVWW3WHaaQuBPvd5EZ1Rk9TpreLb7SErOh3XUp2ZlkSXW
+4gCvQRkD1tIngWEBkmIPt/cG4VYjI6ouDWmCCiQtLxuWAbBW79AFACcMIhaLI0I
Xhu1AVbXdnyrUpb6gjOvC1OFWGEjHVPnp3UhgfYG7ZrQUwRztbwYiCj2/zCjgCS8
fz+frJGMqlquACsFB+vttMqsSbtMJYQCorM/baxWgx4xvMdFd7ij6NUnBp6o53Ab
faVEZi4XrQT9eNcRC2mHKfj3HbZF9HIqrmrSdkri0UOh3j2qIZvYo8bV3pH4k4ps
RCNR/OVpeGnZZKxQspJt82frW2eSHIeRBLrZHZw7n+e1NdnOpzAdsPdGnzBfvLI6
qXZAhmJ++d70Hh7k1xF39T3jeuszVFiFuyQX8RxF75E34yK3AnKKbnPj/703WgCG
2BfeqdgVRNwX3xxEJ9KJpfBuvFnOtNWugl0uwCBDIKZccWpduGZQCU82xMgr/Bwx
WiE9lrzccQfKYu+5zkLBtfsWvVmN0klCH2cYAd5B7SRnVJr6MTWzr02eyEUrNO2/
1S/Yn+ce0O2qlnrXSjy6tpRCXxbw78uxEWX92t7qxyxtCm2gQiTVjlrH4KfKnv46
0yLqOAphSDA1yzH/lf7mY0w2UyPFrC6N3FUME4bENDnSsol7rh42UrJRWVkdijY2
CCZE1c+tJAHJrp+WHw2p5n9RUN00oBMOOQGoVC9ChCPxCEi0QWatNXhUlfZVxrRR
WKo1HccFMsAzyu9KDXDL9Tp/myqanJjjKmXl8B6V5N4yQdLZcUFE6CDnD7GYOI1n
/lZZc7lmgJsD0JQ4sV351/Ije+8gvREndnkpxpKJ6RKGbouRfLLsaC9JJaOXqe4l
E5bx3djhucVRvCjE6oVUOSTMu7I/7RJohLHJ/Ic/Xf7oSP74iLf6yFlKvcvAx7Yv
O1K7fYVrQvm1iPGUt7xnn1u9brMnNF2TH1YtLptdF1wGUETI1duR8pfXAEvSvC19
MtWyEJMXi1VbWpsFqnoD2PgH6snwop+x+qXklHNmoT8nRfooLqOJ7zGRBb9g9jhJ
XKIUbKXoYu8UU8xgkREedH2CuA+yV6xK3fE09Vm4xuV/iWV/QvjP+D2fBBxrRCdn
dTTcyA2ZrODOPPFF4L/cQV14F3vVLGNy7MTwo4DGjmP5X1ABEqBOllZM9QnlGGGa
wVIHVxvyy0fHm0NuhGY85FSsK9vK4wqWD9diWI2N2VOCrI3Kr71keTuXHzwtwi60
ZKCckPWgfjyk9tVLe9YcFSMxzjQoUaH952/TfIvdOmZ1ht0wL8eLtb1pORqNu6FD
pLQuMvZ0FxKxFmn/jSlbzFDFKxDVjTkU3F/v3D7zZV5pWzqrrY1miXQx1UWM5RBc
qfGgRxKtUGrpO1mJ+BXvm9vsTpTQwSKfnLVKJ+0jAHYWcRZUZ2hwS4F8qESvBAxE
ixpcLhz/kZ6mG+kNbDX9oChC8EMsp9UUNkFebUNOJXE3sg6clWpJp611HWud9ad9
argODOCWasPRq3b7eWcKhtn7i0+Kc4pHf0yUkQdw5R5w9jIWt3sp9Egn55kDYCqo
XGnnHUctK/ODw4wo7/4biP7h16xm1zgiLfz59K702KvrOPxIJGXMPW/RFldl/PGb
m35OB1j4lTILKcWJlxLb3vEXG13kUorXtLhy6m2LOKi+d9xsk3hTUJy3InS2BXsn
I4LidLO1zRGx4tHyzHYppD5NR6BG6de8kYOn34zbVgk+byGAS6vp0rTTWuapyMju
SIY5rMXzX1rkGsyQ/slSrTZ+N6+Kb11aKVAx+7Nj8GjSg+5lbPR/qPGofYLvw1+x
iWEVO/JAZYjKmTU5mZMsV5LTCVSv/Le6gXX0Wj2n8Isx1wLRW7Z2Lvv6FVJL7f4C
dWqog7T0yaNrwQnt97Uf2V1LAMBJRr/HSUxrwgm9XN0h9dWhTXnEq9S/jlJuf5hs
SUDvuyTWL/kpwGpuAearLGtoCe+1gjpTJZUQRT+yhEN8o3QEvWYZPiZ6w5ayg9t+
Xn8Y1XyFvnLQPhbogYEf2LsJnF+SrqutkPC2ieGqgyFirnbWgv4fEeU1o0RHpHtY
NT78FlEtIFZs/wg0Tn5cht9IL856TtVwKzcnSZLiOGUd1hl3Ngg8Way8h3UODjKO
QvzZEOo59tFzqcTk80ECEgUnVEC56O53RQvF344nPiTf6zOaVdYPPkFIM0fWjJ5B
gEpmgoPiudVHbIGHlZXInV0AI4LzsvH8hZHuthoUMoeCLXpkAll0xmK1nlstzzKM
OX9Ml7buRH+0yFUf8wAZraUTZ82RMBt7cwuOcxlrg6aX39hzMJ1rHit+zNWDCBRm
hsKuN+dLegxcQGxNRfFj+J2fiL5mpy05sSqok/yqoGH/VaVDnRrieiZ5dz0BkZKA
y0LF6QvnJ5tQCW/EpT8idmUgqVw0PJTg41c9f5nzLh+2SOA+xyOG30QwnJQTragf
Sn2n857LFO+7o1jkESc/Zgff3iFCqukTZ4idaXIFMHGzCl6Jynl2JVwKUL1vcriT
aOU0Y0bEdaR4iZ6VAzfdhtY8pldRuzL2YH1m0Fx1tY55lC4lbeVxOPgBvo2rsRl1
71CUzeLGrH2uBwCHW1qdO8AWUfu03/zLtupl6ccKYCmzDtx7Di7LgcKqbbCleBGG
FzUED5Dg/JDrsq7y/dAyIoadZXNg4KB2IAunMcX9ITREJ0ZzNgg4p0AOwHjPSXj6
jw2uNHLpVOMBXNmI80u8o8LI6YJFDYJehKJ1uu4OZ4zE/fRnC8VnvV/LNhiK3Bsj
7xbYJGbth3LJFwpH5xSvD9DWMFHc2YV+/l9wjKsBsgRT0AdRMxv650c/R2zu9dp5
LXrOorHrKshC0e5K2TolUpsMH6Im1NC/qsvEElMbPWPZLPmB0Xy6Y6SH4a++b0LG
gd1wc8X1RyHi5Jw/sFO7sWjmJJisY5QgY685R6PntemFBY6CWORUXQOat/HaFKjY
pdD5TJG7ZkR92aUw4bFalhZm6w7lV8WiPrhDwgyr8HUGcridK6Ln2dAXZmLDtcPO
iKUN82ZqODYwETkUlcyRwI4EcslzX7xewp2iN4/H93PWDTb7aVBxiGLHmmLfQsm3
MofTAnHi0ELrMlqLoBV3QvSJUnqD9QsnJUospUu+uFhOIuRd5BU8cLPl/JllC4nV
+kmbWcG+mIdw5Y+wJ8znmt9dh+I4JS1AVysuFhclxe9VVa2dvAugIDvuvTRm+vGR
/Y2WuBsfBgZ8xaf8+lWfr8jkWPf/RZ1X+Q6lipCKowCVF6OXSyzy/VNRDsl/Haow
YMEAQ0V45Y6ywTzb9JZDuRYaNP4pw4IK/W8mQjVtjL9oogm+YDrH8QbcE8A5z3nx
yamveYmwAv4+9KuLLa03L24h2GDTSyY+9WMvUfqez2kzGJ0AUFDdJSNAv20Cwg3u
B2TFQE+roHvwpMdHDfp0QtjNOXRjc8qByspDfGbNPtC+jDe7Qr4vJVVrpSVzpAJ2
d3GrH063I3PxZgzxi2HAhB2vH8eGdXaJfLpv4Ltm7zHybaxWZ68HmZXYkYu0najJ
AdiJoksSZ8Bjx/VaxeT8bnxeFtjSzodf8wG51+mpLiyw1YndqKpWwHEo6jbh1MVz
c9IRT9e+9oB5sIR7b3wN8IzvArTpLhOdnQ/7aXpSOHX9SrxGuRtgycHS1tLJRc0k
+e6+B4+ozw1/5prBg6n9HXtxZVKynHlKw31zwJDLiMy0wR7y5HdbcARI07tTieiQ
Ij7YLIFBLqC6gZ4sg3mddUhSvJCxN5PBDl24uF6t0wyDpnvay+E1TUqjJ0xQrznG
sRTMX9j/hcu84lU3c5fqX3SDT2PmmwQhllQjWApY10imgm+X5vGeNdvF6yYMzaLv
VBoled7zdpVHfXPPQNniBmDMxY5koL2NqBOskK/ly97BHAv8mFtn2loUWsHL+CkG
CJvQ/uyxsGiVL4Y2F3OW1N2sfcvfcpyEVgYvmRpPhTly0xaYzwTQfP5VtQ0qy91J
HGo9JXgLx7H6hcPSWQdA/yehFQS+hZ/LiuHfVPzltHuzYlZ9Ki6NaAo6ZH4dqWOd
/H+lliPs9nRZDgeo62UQNM7cgBEJjfXgjHKAJ1jYXKAHx/fZa7yJkj42wN5DWpny
bAvO2bIRBhpkcwCJaZBjkje7JRittLKwzESp7AFZB/iBbz0sijBwlm/yI3GiVUTh
Xn7KpjDa0OPAxD4As2pLtp4nQzbJMHLROT9tKi242K0VSHpig1fR/je5KgVIfxNj
4itgctGUq5/tTAmDVg1tjUaR23OMuUF4OrZBB2oRXnIiDspQYlvJReq7UBq/vemy
5GsODbbZu821Kf+SL5yuvgP/wFB2pskFQRFra2CMk8pbRFx3ApwYW9F+4MUuPzWk
M1mmfsUq4/C8+kdZtyRypyFp/IiHrpTZhxd89JY/wWCD1g71H+FMFT9Q9muR/km9
7IKkrYP7Hzq5YMh4lqZ7qF4GOhRbQ6jCMJhlw4skHiQl5L16MQDxVmkn0O4nuvgS
nAFJtRB0hYGYvyYQYk14FJbUcdy/wOKRPT6uCafhceMPG/9kzsJb+5tgXMGlPvPx
x6meZkEByKAAcWOEvLmIP7DxA2NDSWyLo1RrKnmpER5LebZ6YFdMuvxsTqc8F6RM
5heoWu2hh5STMXhFANeR2+rudu2UcTs2d2+hKDhTouDwYoIUE7orr+RsT5UEQEFw
/BNSBBCIeRiRLtCJeeW/6TTeeclHVlxg1+VlcWMMA+U4+QPcnfacQ8bfbf7IFHnr
hKlvKaa2iPl/4Z5cAjfSL+PAkWYngFktPXVRhVbrJRqhaC7e+LZiInljJnE1yIdj
4VRDm1e8Qi/gTLYhBWmfVmaIxYviRi/USwWoDsmmpYnS4x8Hy+gV7SiPQgk0ro+Z
9pXb+kDxZ6pZRW/mwQm7D+giZtCJ6zf0IhKwoDFbusnZRWoE4B4AG8aS+4A9fawZ
jBKXYtJmrZIjSmXro7z/W0hmx0UlEomM0OD5sOPxH+BIxEivZzv8NXc0YYBrMxWD
NGkM2N44ScSrPCHdEfjuldsTY3Wuw0ukdeM15bfIX3zB36WAqkZFaDJK/K8FeGzb
1qFxSOVwUVIqQcrKT2pipSu7gk+UAOo3HqvVyXpEpcOHd3LQICCy221x7/FAHD5I
0ERsf+QiAeiX6VdODUndDLIe2Cnqe3BmKtKq8Voi7/t8fflbIqlzdfhynliaXaMR
U/rl+p9znGIvJoZQr30H4iFs/GiLiFmEG7/nvIAWRPG2KI+uW88/uUpV4+jkWX9G
Acq4ri4eexempumtpITx3J6lUNu0RPdMq47iVfFqj6uD0rijwNCa8hpJFxiOBSjk
00e5lQm2gTJ5hHCj7pGbc3nPtC30LGWLwshBjLLfAQbJKvAtxjIlp0nCf1MTIGC7
JI+YjQwxKSH0B/fY2k59179X4pvqttcaQWoDqAa7/0pEpwaWuN5FaXY/2jZm0Lys
BaZdpqYoOUti9A5qGijMTl6A0HA7/1keza79/ROJ9mjkQHVnnNduyUB9xB/GiPyq
MdNLxiUo7VMO+PHX30UiBFpgx6YUiiBv/4HL2PsyQVj+twHZ9mdjCnebKo/FUY1/
jCE75SE4jcWd9UzRIgHxOphubNjknKGQwpbyyKtboK4VzEP9q45nRrFUlAVkCpvH
ywGmpyzbA+25re4/uoPp0+IUOaJ2dyybsn13aOnCRTeSa4ttW0mkmczyFeQ8/buw
2MpWfjUewnpR47tKrNm5tebVYlJPgTRGUh0txxXUM2KwnN/FmxjLbhB6PTgjAWQz
j8DZ3fMrug+Ub/jTJWRkLS0k4N+HNA+rHwF90ItOUJJBBQRoJ9sQO8u3swQ9yiKQ
j+xl7LGQypWsSfHROvWUPCI/EgtVT8CKv5ym5fEHMS/HLE1IdjgErNLA9pQ6/muQ
G7de4zeocCdERf2loEWMqpni3JwrtOqK7kf6DhR4s6uLm4iSZQnvWLJ+uVxtw39D
kmOVs0JQnbKpglx56mVoFgXuV/GFALjIgDmf/RR8rGO4h8fN+lHKQeY38y0Xr2Ef
JagNyBWso3epUkhYQBah/KtBbS059M1RDHXz7amXTE79pRyWXaVzJjuC47TmlNh2
7WgUXNea2yyz85cJBnUjYjYuZSQCJJL3RuPyo72SRsgh7z4HReEMO57Jbgerc1xo
FxMwURMQRJSFqj1hTCwOok/mHfSHpzonX1FD3mEjm7DAt3bZYHmpagB+nPrXdHl9
UkwELEW/z0WnONP/mQ1R68fRdXRYbQoUVXTtELF0yuupmom3l2qvkRPIE+myoEsk
V8CgFHipIpGedIznPUlPLeo2ICPnPvzewpO9BrrAf6oIfn3rXHpWRThhJ5LEbHY4
qFq+BdZastslH7UzktKEGyEdyo5m4RSt7YWzllvQF7aogZ686stD6R+E/80I4xYD
+WjTQqWuCBmQPtuxJTs1qYBtnM5Tt+/sxcJ2rVfthgrMTG0m9xF85x6PzpZ/I1rv
iGSPsIf2ML0lO15zHHlC+UFR9KwPP3Bdz4zKIHnd+hNORdWXKMPdkjEZam57qNBg
9ACFsvOcrP0m6eF8vjsz8qscT1/jgdiU662R8b6jANPTMp5zG2eqZTdzmaJxAvyU
0aiRfrUoCJhCOKR5L9qEVhj42kUYe76AvDaEg/YYeFK+qfNHQOCpgmfxZCeUMSIg
1U5tbDCHna+0LMv8xP5kL+79Ei75SZCWLTDedESgmKGEJ/urd4q5Rnx8bg22hN3+
OyYY4DTy5xIyrYHlwnyC6ugrGruh56pQlsEwTMHFGFBrUv6/8kmDfsT4X3/wDjp0
auHTIdSx8DEq4lwFTAMMk58xlTPjr6nlLdN1p0ZTI01YGHm3AWC2YZxTJh2DEc99
5IHoDTclPgXmurzLlswth/bUNEl3LLDPnZhUuwY7uMjR+OSacTwCTbq6dQRFoPBx
Lh+vjGFgnqS5mXhOzamKUMbxpik2Ck6r4qOaEMGdY9dkOZXWSml829b+ec/YpsmO
bW3hURTZfMtj2dp/y3kI2nrJPHBDFu44lq3sKsjLDLvw7LbBWw8S53Ug6xbea25M
X4JoTTbEToWbz5WLxeu34x430aH1hIeIvgILLbj7/wYLgzp7oVNA1s9WxuguhXYl
ijyMeDSklKhQD9ugnHZMeVjNW5xOnWfa6r4ZKcsRzptCrBNH6YBtj4Io4xW0oCsg
URRFqmSEB1DjXcMh3YVbD/V5Cn8vMmHQpbi/U4bdfLyFL4bGxKbmlZRQhPOkNlhD
4jsTCcoYoHg4PyGazr5mOttoIN4ESXO5Ord8qoVInv36lvBnvCMsavyM2JROs4cK
ZqnnSBtOqNnzBPGJQ3XCXl04A6iPgqz+vMU7bRRzj2XEEIlZXvJj8RZhadhpsGxB
518y+OAftUI/m4/gAY7hAgTuT5XQBMUQ+0m5T4uNkM0YPm1UmdRy03uLkTl/6TZc
iNngfOE5w+FelPxeRmCDl8Mgq72wDsClR7eJfZmJygKUNPq6ESiQyVpNnmuUkB+9
8rUMFfDRI+NsSOWo60NrHsOC4OfErlHGbx2c6Eo35XkUeg382FgZWI/Bl0gLGWZ+
KwIkhIVD+ixKUAWIwtVkzCHmlSCPuJmetRYpJyjer1fpitaME3AZnieTLyYNPxiP
akooJ2Km5Gch4UHzpqN5dI5vhzAev7T+EpaCNGjkhUQevwHhkyOGuz6bwk/QwfEl
U8di72wxqy1rAbrWPz7k3ukGITPGvMD/nhxVvX9NAJNFKWdMk+MvrLy5Gc+ihBQo
NJfYiCFNnaEoER6awvtDqbsQa8Qz71cQt3EWPlUeM0xVYsdfyJOFWpdSyYTrhAjo
m2RGXHFXft6RByJJOmu3FR5zfbsQ/dDvCpKuKCiY4kLDYpkPIq/4IsI1lUsYp+YL
P4OrxXx6p2AP7ceYRi9gQZwDPa074Ke9lng73hHwyzG/M13Xc+UPOki6j/yW77eI
nT/yBbZcMALSaCCAnXI23h4s2yG0a4kaK3oPDwE/lMh/w0foTKJW/DU0cQDVJSrT
WLZJgUuuah49tdUw0V1zuRskMag+xFF1Rgm4p2p+cdal1XyXWQ32pR7cUc02emPX
xPc1htpsVM/gLGG2TK5V08YAdbDGDG2NtaYnHtwP+xyICnx/n2x8HxOJuUNC5uJ2
R+p4qbFpErb1l5X0RYRKQpSLMTj4RLvC3n/wTOLGU6XNQ9GzTL4JN1at07Sw95fL
l87hnql2tgGwlY7pzOf73B7gneiNlzJO1RWQBHQocjJf0eucQDZOWcHo7S4UxQ22
sfUDcc7mVtT2mIp6tWJFLQXXqp/qt8agD1Jp39E9zA+37eTiiunUiTdWc3kXCEZb
++/CexyPrSbCjhBv8Kkm9+BNyYkPXAlNbgLPKAc5dupApaMMg8005SosA/9l5VjM
LC3mZxMyrNnzpFYGpbz83Mih7t0APZAbZYrbAxKziBXjp5xR6/iEnyWYLxGf2T9b
rQNuxV59/wdlV8ugU/9lzbyB/uOI01CyAMWOCzspTtP3Tt1XSBaOZzu70AUEDFhc
Ou2EeMP6TSgUC9vP4MOkuTRv78NhR/tF7a80hIbx0m2XsDTvTL0MRI0EM6WDsTzS
2BYj33ghb65ImYjFNtb1zvgxfWF0DVTFy3zujUxSPF4XuWRhUyiUfzrLGgJmIEe3
HP9qiJwLW1Y5/AGMV1CPKaGM5MnzLjMNYAdYKCDrHpO6yMxb2scyAOKuXCRl/5bq
JYOnHeUGzxuw2WQ8YsyvGJzdBZVY/MJkMueZtwlxKR0S+GmtGA7EJf/wPhLk7mQ6
J925m3oixKCVCmd8ecw2Fht94pHvfixsMf4xfdM6z7MLzyf/XQ45fod0cugR1uTx
r6otq3zMXHyEwa54luo48V/53wxGKb55eB9lOoiYmxQCUdVVCAM5Z2E8Q4dBk8QS
EQYrGkBRgRHJqyWCpc6m/GNttyMgdqZKLofxWs7coLVTv8IQNrQROCqdg7RkZ7MY
TezoGiKkACpi+2tLdCxKi28XQnB5ExGUkdZZ3kOVgOZTmr4tfe3PBSFEDJYqie8l
wDrqiWFoGy1lMVgJFaOwJ/QILZQhNw3TJchAxJTLlowhBbSdefIScBnxwqCXPPcP
Dy3zwCop5ImWGMbPmUhYmO56g8q8VAZ6l3CULwDD/I4PKksjvQ6iWtjQ6eYHY7I2
iG7vNMDLaHVCTQoluOub42EePQuB0H6GF6uL6WA66Lrn67lmfuN3c/CvLAVLxkHF
Ny2u1DVWlKkUUsX8qE6h6M+9yCJnUFhw60KT2C2uJp/Fw3CEw+Pq1MDB6EZu/Mc0
a7fBJJ+RCKKikTHf3XnHdYdrbAbF0jICA04wf7sVZ3RCKmNcSdaIWS4OLS/Fj3VU
WklmLMCilZ2Av5WwuyS+pHUehm4LEnlD5PAYT2fFLiXIgrohUcgB/bpiX6Lc5CDh
nJ38HRXoCYXQOT4E8cj39v5oUOk/nDQjXvT2xqGe/3aJxSXshxq0SU4slfU/Orw5
J8B/KzIM69hPCzJupkCvMAW0Q+yzB6UgYgZIvFLUBvvNe94PWJxe+fEA+MoOsjVa
iU0OWkcphk3qoBqOIETS28iMBXoU0U9xp2AuK6Nl4ECPpKEszCvd3AZG5Y5Jha5J
UbUlbSHTztIIEWMttdOXVm//TcEYTYkJ4D4COLE96FBDDic/88CEfZPjCeb32abK
FZWs0ZnuQeF7PsJ17hWsvbXUSR/Zw6eI0PIlIn1mz6OfrgR6rJiZyIp0ZO9VnMKr
klI5KvcmTyrLvzqYVftMB6e2HAb6UAqmBTLmoFmziEik8j5pQBaBp0RGfO1xro6y
G2gail8Y7hwwKszoCG6FCQcyqPgSEkP/IPe/6Pw3P15dEXil6QxT9ietnZIi+udz
fhz28EPejNZsfG585FnjigfLXRqW/aspz5H6N4TOgQxc7cxuP1ZrmCOfV/hEXTyX
7/3YywK9nQNTWePzExgO6GIA+9mqCxonzahdQBbPsHUmxVwVByD3ohoukqk6Yqvs
zijKjOmGjgiH/xJ4g9cGbkYuPF5KDsfJb4vrCSCKEPniKOcLjPHdE2PygtgK375F
yPxqHFz3STosuBxUCadRrLg+3InA6wAL4PCoBIKMQSUUp75HkxH1dO483FXFSdlX
alDIDlsLpEU+BoWFUpF/0B75PUIPaHNmdTq5EmFV9jdfxmJnetDpXwf6TaVbA2+p
RGrz7Ktn2Tzlf8sST4Er2c0nlZcXuu3Y0AohLBCzNYsdisVeOSZbym6PF8OaVDiy
Pa5ffnaYVaHP9NJUxE5doayHZrdwMgM5dyfixS8aVMYOnI/pdH4U/Sv4mgOJCiKg
0uoaDLcV3KNMgNn2lVw1mBxO3ce5/yGNtAQwwM8jA6MDCCXA01OQ/vkLiemI3pcX
n5bNeVNAhYjvaot8YdjwtRBhGqXtcsGlugWh1BcusiG1jO/lcT60ioYWnUvPGW6r
Oay5tMn4Ak5w5Gg1B/4znKC4NPKHKf4WQtIGk9ezY3f98SZClab2qkJ3U6fuWPbq
d2eiRq9fZVuuBbgea2dA2UaNsnvodJU35ElMuKRFyVVhABNb1W1RIYEVvVHuWMSt
YHdJ7RPr0pxIht249u6YvD18pYcGVK7yOvwmICt/JkHQeQ0crSB9utqLBN8Xgi8i
F287LKH41bMA3ycY8ANTjEaORvDJuN25A3ztF35Y6Xa5AiYcNEx/Wugo9jC6Sg/M
GgYM55JZZfW+DGrp/3+lPlkPniJX2O3oE2tOYse+Q6h5LkIICofsXvDuoAWrn0HF
jgJWBqXrW8qdIrmV0SmPM2Q229pE7cjjE0gHPgcU7wuDXrUcrBUAZD2w1zw7afVm
28+1FZCp+jTwgpG4V+a3ADZrq8ZIYM8iRkRX3xwLT1FtGLGj4lDdBUlRvIwosuju
yVziS6m/s3KN5X9gHv+7l1rAuEvUiPHKHXrlrUtv+wHKmvoZSstAXuMKRm0Xj4g5
wZpdn5qNRHJgC+fRt5cbxDHxcB0l0VNHyJrJHqpCn7XV9RQxmNutEb+aohEIHwSc
NhQQY0MzJyQxCH9dXhL9TJRp39kgCYw7wWrE4/FywvGNNhIOwKbBnXS95NgOXh70
SMgmDV+g0NqdOj8Kxw6C3ksHEB0dTJdDBh+i89Y218P7DRX36k4Yk5PFrwIrqEqb
l+xcho6/fHthgymsEXXJjxVVvIemgmmCd1Ibu8wSt3Tgwc/NjiUSnd6PPay4cLEM
Rio9pCNLNqadLt9cyNfoualAP50iTGi+mq4bj5QCPy8ABFSGMT++A6EGrGJYJMqx
Xgg1+DC3Wn9WjH1RKZpQrFFgV0IMpihds/Q6d9XTfU0f2011/HZcMbTrypVq3Q5J
A+FJEenSPGatmi2gte3leOeuH99V4PRTEbwu9bK+BRE4XMbt+7I2eCE8uVRM8CHy
NNnoDlpfJnnI9eT85KCCfRU7a9Ux9T5BT3u7mTrh6TIMoNPHvSzb2qclHwGCn9sU
11uWhR9NfiYnhAwlINLzbJYf2A6S4HIj0rlXgVUDRhyVGHn+E0RVAJ+qR+z+e0y4
uNL1d7rHdmBKJF1Py8dAmnN8cnjS4jLGeydEgiiwlvxW1rLULj8uXtkxJnHD5D36
vB3TXE3lkIx3FDGU9Q2XXXWFlyIUtLLSvLRtuWzcU1zvyACawSCxGwITuVkmQgUA
bgvjzomV/W8vQMukECYHNK5Zwe+havJYpbtdCLDC66O6LyMAm0r/j7ZVONrS7tOh
dWw904R54aRPouI2W+OF9mnhWbNxqcTDjbVGBHcDYZ7UMmAZc3KMVUPsraZqH60a
FrqZeYITudo4dZPWzJ5Nh0JdrQ41dMMy7gHRe8faey5KYJ5PZ7TnL08LPKuuFqJj
NG01k264p7yr6eABehsksBlfbpFapD4j1PTabJyPhWpgOqY/RLFcktF2xXbFWMRZ
fKKWjrnN4Uzk+aiqLu4X7MU/sj+FCJj4uG8H/wdkaxGUZtJBWbsvlK4G9BDz7PWN
3isQdN4nR2Z8wJ5gGImZk9FubDL2QWObRiZvNIqD8ZzEap+4u7F0gY3P8v+ZdcE8
N+q/1zgSpK5akOa6kD66Etq18olZ/TM/juzvH5DtnEx6qrRd6Uaid2UplUJ8fiCA
h2GNTizU+jjSuM/3GzZC61ZB9M+l9H24D4PWF7ZOUMkOPF2ggsuL84zXjKyJ1TQS
+aqIJCwtt9mhPPdJghTwf7wWH4Te0J1IbGRInvE1m89RWmypptaBoyWiTB3RUZC8
vmSK2h14iWbTEZanq3isOIo3kHKv9gvg6WHOdAGGlX0a/dACQX/UaH2ihDgnS3Sa
0DPGe65eITx4SEdOack/4NO6Vkf1S5UvjtUpi2LCluRY1eDhP1AcCPABjgWZriIV
VIhHC7L0q+GTvuVYI6iPPL2+2DQrK3jmD/Eyz6RlQFeCieqg5CV30h6Hwzxy+MUQ
DCp/5k+kgrCrLjRg4Nrg24t1cHQpNLwp/gXwHDwaBtuT7+LoGJvIc74vCYYKn19K
e5YXbicGZRtc6esTM1s2jnq1KUfc4cY4VQQaFT9j03B4NmBfMA0T4zKSKdY7mDha
hVXuDu1uQxRpJybFStMGEANrf4ELM/Nd+HpXWhhBLWKkP7TDkQigI7VFnCQ27Kbu
GatIkNCWB/1xynDv3pzAog07OcUeO9YZwZJwJy195cvolOSYEixZKXBVI5wnvPIF
EskIdaLWCwSpr0RfVOkuqAbW1CSrkPBPSdSYXkf+aQfDmTc4uv6KYTaA5lKuCywW
ywVeWDkKDtLP4jtb3eQz+oL0BzrDq8qKT4faDrjTlwDuqcRhuYmI51NwK3uJn/k8
BbzXuOdjW5T6igS47Jr0eIGAv2rPX2Xa2GJuxFNqsI5FjxelH7vl3klCrkmePquG
nuFaaKv3jidfRtLJrBLZmzZM0qrydVYXe0ANPct6GxNTWVJjmA1CirxHYF1Ak+3X
DuTo1Y8uvUQGqOXvECisZQnnXPjQiyZSGI8sWdDkDXozbj8Uyb0DkGeem+la4Zcp
R6PIcNEqWx+3cwAzN1b0L7DNjTfTXxGY9VnhKgtcMXFnjA3OGNFuq5m7VyZLrH0r
7pIOpL8nuFjjTaB1gh35xpoRQcEGPuGvHdNlSNArZD7DwiNzL5gMDxM863LVgNsP
VcEI70flpSEyQi5vjQJK8FwfZvYy7viw8xgMlEYldv5tlxTH3Xt8zlxP7QNqh7sd
8hcV1l4iQfjI9atJB40D32B+XejxBZGc6EbJ0uE/1HmUH/LKE2TaVzpjSrEe07AS
gF7ALqICWhtrsTQB1T/7U4orFYZFz+8hYAbzEECCy2v/jKyViSSaSskhbJGCbEuM
l5lR2n68arNgd+5iD4d0BYmpEmbb3Nc0ezqc1E9Lut5NJoKl8Wy/FjM/sF8mJ28C
R42R8hmNY0wazooxXopnAhE9svvuZzY8/j/1YHqlyNVcWmOPnCa/TKBwE/KCNp8s
fVhijqhKnrryemFrmudfJivqJE9RahFq1mBEcNiP6qcQGWNDOOqp7zDnmEp+Tsll
K/pQtNKOL/H5tmd0tRFr5Nma/r5JOL5IOFC/w52exhkHf0mdinqcqfJ4p7rpCk7i
cf6nagTMpPj80Rez6oZl0KPV9dRnj60WwlzA+q4yFQT1/ZvgtOi24mm/R9Z3qRuZ
0nIZ/Km5RURjQi4OddgWp96kW0ljVvimRQQJ0vjqOfepinTc/O4WJZ1sSXZACHWk
a5OtSf5AbWt97cNPDCmVPrzkwG4Y7NVjcq9Ji/MlIM0v/LI+NmPJRlXKWjZoe4kz
63n4s63vwZ8apT3+uR2wSHJ557CS2wEjp7yND9oPZTFPhf6uJvcvAmAIzKsLh6zG
oryEPm5iasrPcyrUNgSqwikmTZFtJvWZtZMSswb7pODvCYuDW9W9NA9U4SBD4riG
hO6BlkVm/jq8NkV2+sghAeGN6+8/RnTY7h4AEuGhgRj5FCHylTo+/Xi9VPjCgwTf
uCMeALo/72LSjgpaj2rvwzTwj5fXusiX86l9/h30C7EGMWJo4US4eC4a8TIEPwUk
Pg3xXh8Nt9yA174ppkxZ0BYLqYmiWLTMqEpYO/Hs+Wt3fnIYO9GASkyUTelEXtkb
HRcjJPtO8QH+P4BO7eeN4bCl3viVv2YIeoNYWRqxTU6PEDrsBe4d5Vy3PbehYcCo
jdccLkuhZ/viguGM7AkiB0slkcW6Ldy3nnQQ+Y6I/Y/YnjfH0TJnlgVu6UKOuZAu
upKqkl3Vhfh5cV6ZI7I7Zw3P+ckzvrnxHd199RSxpEj2ni5k5glvFFe4R5H1D/7o
rgfbWiTz2kij/CS2x2PqMGZ+PaYZJxA3RkEu0XbDcPiRjYfbinIV5MimA6mxoQpe
gwj2Anj/KKn86kV89abs00FxKJf5Zqn/mUgYGJYOvDu1TyhYz7nO1GGpSVNiuLRM
YeHT/ASczj/VR60iSugsjuSSmulAAKXDJ5r/CPLFSclS2cvXfyoc+ZA3fAg/UJ/2
RM13w0vbf+VbyrJhK7foLARNaBE/244y7EUBnNcPFnutHhlXUvd1GgkUcyZVyaOo
Uz+qgu3Ge1SS3+GwZlXFsawrLqX6V8yQZOmGK8HHDWyeuPCxS73+KIjrb+MNEIwW
Bf9IYcJdI1vk7NMaun3IhDJAH4T3tXWLTkUsq2QbkTzFnUERNng6UKvZB/HvOHAU
haBI4kCm8IYKJpldoIvnFoV+hAmUAqwl6mCW3Rad6YtHZam1Kay28g2BAKX1cv4j
JJzmyx+uKXXWD2KrCBymwgeIhl43ET0UaXH4bUk6gLHs3jwxIjcCTCGqZNpVet0r
GaDvVw+jxEhugVNGDhgRQbSU53x0OSneDlRmmkute/4ZqdsfUWFsdfuYYMGnOPjs
Zej05QqZoPZ5DLRcxxn5llzJwfSYu8Rsc1cSzD0B6Bycv8RvXB28F2kZy50lahE1
s6S9N1uQ1QaBWnOOjMoS3yTPdInuG5iyrSCbkOMj/Zt58I4IvkeDPTqqM7OMrHNp
JbpEn8dedkiA9iveoKXpN0SIyznOer8ZDUkvjkGMtNi/3dKuEzrB/7Q8RpWbi0Ac
Dw5zI/OqJDXyhxwbukMy02tb9IxwZk0Hxrw3/fqRq6vVXQjAV+gNRRHM2HrI5vtZ
dnodrnla/aJT9WG6NEVxFXH0l1RCmuYmA2InB9ggFcTztfivvOD+8hbdXVEyWnGJ
cvUrK9sboPut8PamyQWoFpR1tsNneTElbDfGLRovH96GKqIHtyyY7vttAgIGN9cT
wZirxh9uKoAg5grtHMQe4K9qoWjjXOF6ths2pKx98bo/3vVFM80yc3zVKfHiOWdn
MeIfnFOQkh2zfFUgVT3kS/jNKB3I1cRkICwy4TMsHsaaCwiZG/mJQTvKPvb58tGp
thxyNzIuI8LW9O7gOyxxhJJmDKz3Ws94P6nEo+Tt3bQSh27y+njqlENREugX+0UF
C9WdSviInEkn91fsEHdQ84AzVtOts7e8xHSmvNdeYFshpezDr+KUsvpmIa0WqL9K
pIgHKw3DOj2QLwaNNc/9W6dCSiRb8bFGrbNFqZyG/puBAXBgBCzKjSTHlqfECGeh
m7cWSwLC84BQOfDOs4ktfPAjfWE+SNhuYw5i2jv8di5c6knbDi9h8sbbhCIqk/qj
lU+riIR0dEn0icbO41EOVhwioArCaMb2TOIvTSAVnUrnijOrHuBVJfWsVIDEnDX+
MjIpKIYGBm5qpmZA6S9d7OjpADkpY6Y5z4lxbiPXgRk2QLeXuobT2rxpa3apUVC3
mrDeiPKTCm6I9mhpy/8ngIjje0du4wXJCFMkYAxLthWycvcw5+Kx2E2zZiv+I+T+
qY90ys+q3iS8QWExZtESJYHQf9F2Ma9gEE9wHAAFiDJRlAl4q3ks0JoKXqiwabuz
cGqN4A0eEATZsKtBnPwHol9DJCgfRWoz4BTmpAyD2O27jQeHI0iIx4WURj2RAMtS
BaN0GsrmmxLU1rSSxURGCJLXPDeVRwexsJIsU25by31PmzWITK2KG1XOR2M8Uv0O
yM07NJ0mpBjSjIfXU2au7o6YAYW8gOAQRKmX9rkOBWeXnZj8C2coBMEx1wIbtKDs
HkH2FLyWaKV4RGVxIgY6lHPJHSnIziVzh5b2IuvSWWQhGOb2NMosbIH4nFHPycpm
/Hh7yDCO2CB3BwFf9QAmemIL+d4jYQ74BxSMPfp+xevoHp47vRGXJ+u5ooam+VOy
tftyzTVhR+y/1cb+QDZZMiVlFKKB0QWSrxLXGdOdlZIYfOtKV1xfyvNF8r8OWJsD
2+/jmNWUB5E/Smt8UnAD1AdcjbNVJklIXJJJJhvx1QaI6HAS87zBptQNVbReRfkI
YaggYrZMz36HdOXy3LhTPmVKz7pSWoRBVGRELLyBzIefnseQ2gBKLnT1LZ/SSz8A
H4AbpT3WQWIstobDnQKFxIxME6X4f3u0cQqFsKOGJpePUullZv0f+lmVeYjLFZD6
uWIpWyUg4f9PbnXle1dIrOhsGC6wJupr9HOSMfIkjDZoSNYZyM8Bq8yOF5Xb8SBI
rPIrSrQQNsBw4FT7IpO6bj7HCqJAN/sxpXn2X7rfxhMpCyBXZoAn2VS3N2YsKoBh
7MiL0V2SulmL7qKIWBzxeXAuLKHImwTv/eHUg3XKg2gY1ta/xZlQSRgtQjqbl9hL
AFtjrnvtM9xptt71ffCcxgDYRgLtkyD47wlw7W0fGXE6DwnERfVMiSvTvyb6hiRT
vgcvrc/zbVcFH5VtOb1cbGRq0Y8H13opk42d+0VzVXiaBtKhrFYOv5rXH+Q1rfPN
XM4bY2iyhuMQILKGmltsDcfUqoq9v4H8T7AdCio+m0f8BRauJkS47dpe+Uw/iJw7
5qKjiJWH75dc6bKGsV0xcOhRKVj4txxO4EO5nlC3DhAsmRJWBrjBc5oKv3VExRWw
3krECjPdkH4sdKIBUK2dVdJ+gsCqxojrhafrM3bCuGUYrQeixovm+bF6S6KE7oAO
fg6riVsC/rqjpoap+4OdJlqldSPdIjKsdeZnmjERsfXWvZJC8Ob6qVdq1jlB49eX
T0sW+s54JB6KUsA7QnZZYq+1DGOO1lZYB0XZi1trh2e6rzdjOmWVOBWN/l5F/X8W
VRfdwOChHiGOwWZGeoVlnQGAFA205HaOk6AC2fxgBvf9j/5+LOuk0cwBCy2W5xut
gWFxR4HyxnsLQPKOGifMJ3nnirMqC7rlw1lM4QsmSS8FD1tkdFkR2Y2hTcRV6ih1
yHiXROlPVASfVNWDPx26NoOQIW0py7aVWdR54Ad0u/byUVHLiuWHlZkejqwWiLUC
Kpn1tfdpj+wEisaKNij93j+FUcj6E51rUwKy9a6IF8E9Ary6FEdqRZlGcJcdPVy1
T3V0e8oEaiGRbleKQp70zwiN3gQfPX2EZq6T79zf5gAl/175QA3VbAv+P9nYsshh
iJnl7h/x/hYIMyJFhAFm9QFTGpQPhd1tqcYVzGe457OyVUY8o1pvR74OJ7BfOoOM
kr4oEp+2U+4VBNKq5VVw5TyzlubPMN9iGuat3rO4ldHDCtE+59Yz3fKtVPCFQ8Hl
TFeaWtMIF1/Z52NRsonw1Sid4PGvT3AMbzbGiNCViSj1nTr1O/SwhDIoCv6dkJw1
jmnt9RYLcARdaHQcUQzDrX5jof4kQT74Iyq+Lk7d+CRCmgR6nZZaks7K7Ynb+hAM
TYynf/kgYugiPD2ElrRv9QFuSe7KZs32VAqyHu89sQRY59r04DTd7NxsS1/ll85k
KsHaBLli6VY4d1WVbwC3tyUpj2CH47VZR2rI/rVIhhBexZO5a2RB9EhMG5GE/loJ
DsuP5MKM3hChqchJpOcbkzoReiBVz+Jy+hzK+U+lnhJUZF6vw8/ASGMzWwUicWMG
Q3Xbx+Te1HCCKAePlAdE6De2ucqlTHzSDRuX2XLCYtvej/hPlh9jDlmqxRixS4un
EPYW5GdUrUQnU1+84PWuv297xRFKzmINSE9GMX3pgN492KvGU7ho2bzGsQY2NTcG
Da20b5QvkoNiYk7P/ZTQqUIEjgQJWosv6fu1/ydW7uKauu9jBkZFoTgYx9yvRiOK
tqz2/vW/6NjNMRGAtbTYqzoOj1jrslbjpac+nunOGLY4olSHWQu+HjX8Kfu48bZX
ZJaXSqPuzm9vttjm8EALp+rATLbewvPlY/peXn0iUTStEVvVI2ubtSOLAnpgCGVE
qpE/x+1fsy6Or0JoJGKyVIMijCr00GVVTKCeV8MF1nnD3K2yWCik330Lqg4neJP4
Ywuvf1bU1KbUQnY3Xvs7YMXo2LRPvXe1V9+LNneNrpv2QaYSAIYcTKqc0GCl9Ubq
B2i8dtVZk7pbCX/N8J5oyI1M/hH0V7NoLFNvQwNwJ07bWpdngoF7Yn5gjPJgm2xg
cmLBXseDgUDrgU+/hy729Lh6giDjVxBkRcFzDj+0jb7XqQEZ56F6yREehJtBrZuo
MrQQPVuOqKo3ICnu2HwOZz7eCKgwCaB+unh4+Mz0el1C+XERD4DsAE+Ig4UFrcMK
R3RodgaK7odPcfH5fOQbG4BcdcF23jCN9HCVHrCGR2G01EH1gKJ/r7UNY3dJ8dEq
RP5uBprwuNXg84a5etcUV0qPU1ONapITDyq6oK27Hwr8iC667w96zl5tVwpIz+LZ
WgqL1Ik1Vv8ZdJOJIGY/QZ97bFjek0yEJO87kMO6N5aXLXkZN/HIjA0Hf/GkgFm4
Yp9pubFl+TNPe62lzxqOSMz1rZWEtMpk6YBmn7uu2ZwIjdhfURL7Eby5lOrQ97I3
uCC8xPSXMov/eNU5txsFa8p2J51qbyvZDq1AeikOwWoLpGUsxOdIawzNJubCpSEh
/WG0of9dXqWCtNVEcK30iJ3103sldjg2QI1mEHQ6ZamT8wNY8RxXSqerDkshv7C+
bYVSTn7iOtQEfMZsYXpe7jjQ2jdmGiDe9nTY5B+AK5wkDk6spczshwWz6JFgY3vd
oYzA9lqAeaPdAp5CugiUa/8nFoSDNYxctCQ+K+HbhVO1L1awwWkJMOSiPeb44HCC
Y3sz+jGcLaDqL1geVoLNRLGuJlOfaFQ7fYI3IPvGJTxydlto8Hah2FWCE8IHn79m
2v5S0siSEl+0d7UAO2M3xHWSE2VaoiATBDOXoyieCP7/SuBhC91gddpNQnrmgKqa
16dcJOAelfe3iCePeX8e/K0Qpc6259pNlOc08iIjwtMNtqhrznaNBloGCfeG1e52
EPTtauUsPL+ya0fUsYKbXbkXgB/yBrEe3FYtJ9MQMW6DU7pCpWrBToqvIIkuArKx
0k8WIJGYHCosyJXSlbnUb0aoAId2tUFY9vn9tatq0fVNDacIE2S9zE/YBGSavS7v
atsWoy+92+ov1wSQ37ouTfm/NGIZrpe7KsHfl31yAlmn7na9EX1wG0EZftH3Tu4W
TFFzmar5MJAZkkbd7PVQ27aWtrjxQ1urJD7EitBciLDCRRKdRURjIiummKKlDkZD
gbzNsaTPYQ68dlcaL79sGHDIdTBriqYa/+L5BGKOhtDgdsH7FwjnktC+mbwTvOgu
7BjgXdOYncy+x+VLZ+k8uiJvD1g5Z22wIiMvBZTfBsrDo5AyER5H0auHh0kIvqOy
wVayie+3mWmKb/V5qVeZ+qSDfmhVbiR92zCxqHoXJaPvPBFEEmE9gS4aBWcAqnIv
CExsxDFSqg4DZRkImieurLfROdlKC8EUXwpm2TI0taWATK3GR7c2mnwYN7sI8+KU
1wW7X+XoKR5VYEQH62fsbDMkPSRXolUGO6XNfougTj1B2TAhkRVHAGccwkxEkfpj
nLrIYcj7v9l8VDEZFrdNevBH712/zVDD/WacQFRwfMC4SvJr5SS5n26BARWOgsHC
435xTLYZzcEwWvWinhLuHUQJRkQJ8YZYYwdAysPUdlUZe731ed+NFkopG2igr44Z
Kc69wRy6MQt8e2V9czOIw/AsI1bSeum2QQwHFyMJd4M/DlrpiqE01g7dfFiu1uPq
d7oD2dJvAznM1zJlcHG0O+O+C7dV06nbpVZYY4LAH4giIWuXPoInpa1PvzOoLydb
wKU+w9aZXhj3iKlbo5j/U9RAES5yl1L6xHsyHFnZ/n4fLuEaBrvV+Mjq5TVq6ZDX
RR3LwhPXkWbGbTcpjkMm/Rd5sWtuCeh+RVu1WBUFk9OAn4mdoZkRicugDsRAggG0
Ls8ODGJK/3OA685Pks/tboNRiIhXHaiMzSW875toZ+rxgF6IkLINb77JAtd7fi3M
OSV3neVJFqkqQeQWXUonT/xtq/+E+ZRNsi7KGlbxj+N9eBNeEYAOPbCf35wGaIba
y4lfEZLlqCdUqQ/SRstIjl3ZBdjU0w9ahE64vYsn5ZNtZkJ+43/vF0SgTjjymaaK
vpYXdR3fE+sQKA4dXtbfiBI8mUqecqsex1s+ubbfbKl4LTzmOqqaq22bld9Og67i
maRlJUCkrruVzluaKHin6crqRqkUOnAuT+zZNRQ6LBMrnE/mqutFCz5N21ujsSFY
2SRuz1XdrA6+cyuL292uPPIlwGpvIjeyU3QmaFnR7Z5Pg5faMGoO3weT1Eg3RmBj
QhygY3uNgTyEEDtIiWAeeHGWPgLfFSSwbL8qRBkMxGeDOLorCEi2NM1+DUtasrjg
UZ3pmqNxU9fDtR73paFv1lVxyS/duLCEnb/ZnUgxJQqxqsqPrzmt8qM3ciJ+FH9t
mn1hMYSEdsWdgX7af4x0HG3TS2sFU75GQQTVz9zurNViXjJyDrkV2xp+I2iP2/L1
/FQa63JX1OdE4ktf5ISVsX45s4mRssB+JI+D2WktAxEHUcr438cjuEzkRN0XFP9M
QbtfnteNETZKgC6wOjp03YiAwxeF+1+IDeka3uFyKfXtOJcboiqnrwxZVPfwkwn9
UttPE4jcY5/nlb/kkMc5L6igvyUlPtaOQV8GVS0v7SBQDRZNSZ2mWv5jd+6EyZaa
KBpNGtJ7MoMjhsomfhYgRPSOyeRjbbMySmRTvKzz+QQARjNfr4/81lQXPRa/R90u
fcMfZRev6e0R/po88aTgNaYxqaSQopSZKVBXxYIhEEhHsGfp0kXD1LRmfigo5zDx
iMoQ9puvztmZPBu/qL6U0wMvBccLh0BVyW28KqwkEuQZhOQ/Fr87ztltCW9Ney9N
IUiIGTwMK65oslnbPEL72HsCo4njhbQcF5HaAHIzAvwBpaoUILM7hvEudn2ypMY9
rVbnOwmw04DbGwlSLUusw/Wl45xJKdD2nYEmiWuejH9Y2d6oZXAJtZcR4gbo3S3f
y+33wbEjpPjLvu4Hmph8+mPk7RoWQA5GJ3gkbxdpzCSVizJM9d27wT0lHHHsWBAX
hA1M9ealIDy7kCdlnqNXXGhixmaVMZ0emmarIof4IzOGMUMz+dgs7MQUi+CTdQu9
bxuQjGEc2oH925fd6NvUq7cp3z83/UACB7WboH4hLsWIXwBN1oEoNh7dqJYOseoQ
lZGHEZQXRdj/3P2Byvy63Vant9ZwXM0VmHiueyPp1rcJJ+u44DGHdfRzcCKhIaJ/
uoK+NcgJWTqqgAiNlVDLJkwV9Dl4sL/cLUCxTBBvtgmjroWy9vFRiIs+JTNKxREW
o9DqH2I5AqS1H19u8E5OWvDQHwdhWumjC9iq+eevEBPVM4yZQ7UMd5liQKaxOuKp
1DNoATVObtCA9/7SVoMO+ZCEp29JtyaCBWikuPkvPW1vEN4Si+8EjTMFytCKcMP/
i4R85gUNRdMwFVqXZL1lAtUBGlJRAH62oZXx0AcN7c2wMr6jrut1gdS2AZ8VXPr5
w30aP76+BpbKeWKq/hJIKpqQOttt/HLEeMlu+L7xrVvjO/yqnkn2z/3+Cf/Q/zpV
mVXYO91cIjZ6cs//CJhBKAalqiM/BmAybloRBLQRm2cjrlJoFG+ho+SOsELjqPhn
vCzPH1jFrI9Zdr2fxQAnq6TDQWnk5HG7Sith3td1MKKhYF0fSiKfy5d1pdCBnGPm
0wTZ3VlOG6WJI5zpjEFZH2bWpr/kWJKFYLu0aFSqpIyfmZxr9vy+TUFA7n97uf3G
AQhOxjLZ0OZZA8+bEDIf4Tmn7zwKFJJ5vunMI39OEItgEV3HDBgxVJKiHdEE073G
erfBNdQ7bsHtABeSPhtOCY99vXkprSiKTAZMEbScVPVWKqnVfHybWgmfxGrcJmTH
EmLmoh43R2BCfEXuYoA/O+wHU8F6ZqIbn3NdQFedOOUqQ95IWGm5NBx8KUYpvyL2
BRJ/eTzNpkmdRtYwwaKqgzVhi63omD+8Y02UnqCp/Yh2jxzbtY9WCgjg7Tdyspai
OYHA/i9LAFDcA66XGFIExeOwhJaX09mO8AGoZycxSCHPdJQ7K5g62Co8BFM/5AMz
shN/E0pDlZwHhFQgjSd4L7ljwvw+gw0tKDTMihh9dkiCdpbivbCkTkzhyLYByXMT
XOlxXdNzqpqZqiLzQXC+ijfVTkgnan3yynMnbNvD9IntLTsMTpjaVlCHq4i7NY5x
pf7JJL0cxPjo6DuEovMyoVXmyyGOCcelMVn/S1cN1iL0IhsFryxI2TLmzrHIFQ0E
mzQAxKkZUhilYaZa+Zv56oJCehwr6awxIwmgWO60kOF5QZ1TbxGtFbpe3aWfzP3W
o+QZSmfGEylpz5m5iMWXnhCViZqqiqfKSQg1u8+BkH2xj5tK5zJR8JrDGiqKNWrR
C7phhYgyQM0S6vCGV+UVTqnsgr/gB+iIPtl4uM3fGhq0tW9KTjO3UjMoCESJ6TYw
wgfYxSfUuBfzCSEr06sSBmxrzfIhH6WdDVlXdAuBBE6B2aWuM/5F4aJdL+uDsRNY
lK9Dg198XFsbc3e8mVL4QsK1xah0lb8gKHIEnufXEKb7l3Myvm45tExA14/GWMt/
5ZiVkbnSEC7HZokzBxxOqDvcy20MSYftMkj9Ioue0EyWF4Vuw0nCZZJveOyWzR1W
KzJ4Qkrw9+UNRcrfWFdKjkkmDSq2XLJH1UW5lCpoLTiCpo4owjy6phlcK7+kP+gN
wn1w5MckTCWiR+lqLbHVu3TUXJGQrmbPdEuGxSkq5SWiXAR3ncyIQJ3zQHTVc5lR
lJf++rXEOKpYwbki/0Xb4XAi7jmYM6uEhwlC43IL3x+A0URQ3cVxNEKyEoQGE/tL
F3iIakr2BtcyXOS49azx+OMmHFk/w3X9l2k5pwBu1fH6aY16Zpb5t41KpetYOQmo
8Umho/7bZaKLebnMkfrHo1/vzmbVHiHnYtvCAsRJURjC3Cr9uUU3wu10tiwOxg/h
TcdV4WMoYApEgL2PpC5F3Ivy9Lz7FL7I+/WNncNceCcE1TwbhVnDiFEOpqvk2sw4
sCJNsna5MEflAakhtT6B/+VPEYA7IGYBGNSzSPpUmjQhZ7ZcQPCEvZlSrTO4fhW4
c9l4TgNX7Bgdan9O7InJwaHuSw6y7UTGERdEf5CU06dNEznqzWlHEMsVtlgFJXls
iCP+xwkmQQXBosB+b86mA63cz+uPANvXAhJa8ESPrzRdmt42EYEySSAUTdRCNYXE
iKRgFBlfS/dmnsbqWG1zBfUu4AjQ52Z822QC42+PLohqA9q/P0TzGRM49o6LWiSF
PTona4m3g7Ciud1+gFSF1R5rRW/M8/i4zH4u9B0EJgTmBZEiCSlu3D1Wdtz4lfQm
ldX7FH5+xorlPhCWxAo9nJZpVn6L+w5tfeKVjwBBsXEPMCnQxprU1fvb9s/w0/Kn
oEc5yTTK6MZu4HtZM18TnVzdZ/UsW705cDlBMaNmsG+Pk62yFQ44ig8E08m7Cn7q
mtxKgXWHyeXhkJiu0w0a2NEeuHiFrtenRV7rZHFXLRZPicj62V4ij3a/Qpck9luW
Bx/FZODMHnUPOeLBaLlOytBcqN3Qgl1aVWuxYU+tFvAixhqhJp+/Elgem0d0xin6
VbQETYfUW+h5JwwqMUsWHDCw0p/vSC7FlVTBJKKYGwUl4ozNEf3ebkthrpsfoRbq
h9ktuFmRFPWWD0UrYQ+mxz0E8XtegpQlwEZGOd8Q5nC8zs9KkVk/3jNvRPUH3uVA
w06Q3tYk9Z89AuZQa81uGXa3pER2X7gq+Q3jXfrwHy2ZtlGoToMNNSdDKhK4sEJ1
nmZ63d/NOvOIQari+6nLZgR18oe2mUCn9zxsG5Tpl32DTNUV55XhQsngJfv/hBWB
zMHXwVVm/KDH5dpnenWaoeHPSFI9aRbTLnGYUcLcrF0FDB7CgwIj7EvI14z8ZgnI
iyV1xaZV8WoFKEUNXVRWRGyCWjc7zDdS/jJB18guBkPdd5a1RNondfnnBq4/yNvm
ZYXxtAKn9fmXeu4467k/7vRKWYp6PhNjiSpVqJ3cp2AgAaB68gl454vAAJgKzbJr
/Yo8RTCopF9eBJnTfsSQjQsZR+3nRlqr/lhI9Ano01G1fugFAjLGckx4lrnj4INw
Gis7tDlmNHXLjFjCNv2jy9UtibTdrA1tEMXXhEQyqIkNCS9DJqRhvivQrEwJHSXf
ojEs1C70GTgJwIQGhk/wXxaytaocpEwRuQ2DuJkH9OOzpJdmlksOB8SidpRGz8EA
pFhRKNBZscPqoezgZw8kI9soL74C/hUi20L5pTwTBSEspzPyk2U1ICKp4/0B01JS
tJw3imJNaEd2zQN5g2cCI6bxFJ8v+eV1s6+xlKxXmCHFLt/E44vIlBlX5ukrTUI4
PkPuhIChUy9/+fRsL2/KMhrqemtRxWhiG+G4Cza+qpUSaeOo/yC2XpniuvW5iaVL
dghTgz1W2oGx3gqAewPWse9RFK4R2n0sM0a99tg0CLI0pxcrppcKumB3a/iRlpUE
uFSRaK3hFMinWwwxyQD9mUmWV3YKSTEKqvDKS3MZ42N/tcdZIUtAudJz1SLGiM8r
1PLIjC/LRQS/oMaky2R+d3EXHsCjKWOhpybsd3XmnJQyBGsnUhOsRxM3mk6wwB8i
pIwknBog9my2oWd87a45w7s04kx6qCSc7sKyJ2w3QToZ+YB+aCyz38o3zuT+nq25
kPAkyP0542J9OKN2UY4z/kbSHqYmIX0JeoG8AprUTwqvRePuggU7UsV1138jS68M
66kvcXzm4LjW+DKO3EmRiQwJJX+w4gXwV8bfO+g+i/Y/43l+dCGdKnpJsWzHbVOL
16OPHGr6XxjMklBDJT9r+X90ywbDw0vLi0k36fBhAVkjYrXjyAVs0zXB+pm4o0f4
UQQ5HdU6etpsmmKgwI5ADlOK5MvALwwft1eMgfJPr7qyYB58scSKpBIvMQHLf8M7
6g4IadS+9KpExYbZZaiejCw1FcNHQS1YEkmFgUId+bwL7YuSccgx9qcHuGWq+INY
rHweVa7UgyuANEys78oUHzoJKlO+9FJLH36c+jOJ+iZbCnCmr3w7iiFvWaCyPq0u
Why32gVIZZEHHLxiIbXeNHauEdQNedQAmkxaWrAEfjGqNy9kS7wDlDllcRPMs8GN
k2dDUi63hYpeC6OLxNJ1Hmq8cKiQVEqjGpB114eXYrzkn5GXmd89zItsD8HUPzln
tzH3gWa8ryPJC37aJCTsOqVKAnB2l26FIEHsNgmaw7foFQdSEA3KAyJa0GbiGdIv
sDL37puzXI9AeKWQyP2QVw+X0zDBgs9kwpGq+DbdnwUBq/3Yvuwpgnw8bn3u7l99
D9sgwVuUrYEwh+KKNY+5ngI5S62E6Qj25k8NrGpVnbT7oRImUKsHP9+ALfQQJ/M/
bkHHu6DYvtt2Yhh/n1GcSIIAM2bf9HAWSLV6mEYaD9F3h346fWmZmjoFWalN+DgQ
a7VYiX30i9vjPvA6W/Cwi3WQ5FEdqUX3FoFo2YDUUCsbj5prDT+1J17my2PhJdR/
idfTaVLo1kLbM66UPNz8DDeZilce1cbfFkZIuadX3Qmyn5LXb6EdViwH56mkA04/
xgBfijsB/GKHN3lMT7XqICs/xNQTkrKyJ6vwF9xNfKLcxWEww17DP/ZGDq7lv1rx
MKX1nvMEgnkU5ZK4Qb4K9w1XJn4clojw8R4OZpavCCVgdxeGN0ZCgc1tgrMlJ71b
BNxJFVrWalZg7B5XKKU3mguLEhXXmzqQOc54kwiwaX54C5CbsDTLFUwx3K2nX9y+
XHlvn4GgHoVnD0v0bmYeCFH91TRBNUzmZPmcSArmRQLDn0u68YfcWYoHUPc4xXfI
yA2JKaVmoBeVdGd5p6LA7cN7nyqT0dx57qksyZgFK7ByeaDjl0QNPeIbyH8kf175
q6YjH/oOLQS1j5uyFrBbl/ux4g5GQ5TESdjqRVkAWQroA5sU4bSPUFUnde1HdhYs
2I+IcqjiXSY9dmhWhiUrdQSSajOWpne25g/hGmpDYeHImEP6OfJrJ+N6fK1lm90J
CP6NIvrLsABm7TRbfLQwDHPIBb+ucmqrMwmjKW2+HpczCyd9g0ag0wUtA6Uw64qQ
mNx3yhognY6DvZ+trHb0ZkEZoo4rHHGXf5ga5oD9vtVCj+oYT9o2yR7YIbgABagc
rxmaySCv3pwRZ6A59LBjeND0V1OoF7Bhx+cyo9gL2J6qzZIX5l6lT68jggcnlYd3
fqp1ynNFIdLI8Vb+6IUayiMbesD6UIwZPtUlApyjBBLqGdf1X63ldmw9BHu68JhJ
jNZBCHlMHbUHXrnhGOi2Lok5ScuX4MERaT9t37Xugna5YjLdnke9RPTkb3Uzvgnt
UsdFO63ewuGm+KOIPk29cBYSQTS2bDEOvJm3JGy3uzNFUpDJ5Ubs+MqQTjX5hs3W
ebfmxtXn7fjbS2x1p2J8eRyN90e6yhYjMr/z5t40yYUGZ4AJc4m/7yvr9uJZHqTs
od0se6TPX1A/3akdoXZVdnNMdgU0+7cV7IlbTqDLlV+1SnJHPQTBmj5vcViifebl
TUKm4pNGT/4I/4/kn1elm9ssB8wnUkSGIv4IFW6KIgSVcmK1wR8zV5FFqkbhZ4ia
sYxUcFU0fz1JxXY+FMEykSaZImBnQbM5J+IsTi7IexAEAJuMi8QyJ+B4kx/g0uWm
H4xyTVPgKkvCwZBxdRiJtv7KAY/07Oqx/bTmNhph6FpAzgvGmvLjusp0kji8IUDe
xl2H/kQ15caRAZ8vFMPfnMAyzdwRntWjcJBTlGiyEkEk/KW/ZptRo9DSrKkmoG2g
87ErffUtbikyPK9z+3PitsAdHnWS5ddzLX9xpKC6/Ds3wMe7V9cpAGjNjTajK0me
tV+8hmLJWeDQUUQDR1HVrAtW2JneIPGQS0DTQpiQTmc10pm9/umPI8cbHNuvIs/6
Q02MKfngcAjNV6DhWLNwgBlZEriuhyL2ZVb8yS65p+dT3Pfa4eAY6LlmgJRi+cSt
xdkNjy+BBDys28siaeCDyjkEZDSadi5O3dvoItrmkNKHvx+ZzaAA7nvglS2s0q3s
DpAANH5A7x3q/antavao2nK+dbPij/mUI5Y5+F0BHT96/xi8jgIejPtZPqBOznf1
Qty2akrsK1JP9gdLTHUn11s1EEt6ecnxqeEg1Tyj9LGaW0MX5AoDV/UtJe/heMR4
qYzZ41DcfXWbg93toXWdXpmkM6Yth7gU+ekaC6HFla3hqWd1k07R33SJHincfbz2
eSPMezPBOfigJZautL0d3ZTKjrq9W4pYASdVdax4YXtXjTtL3Jo9O4O97S5P+fWH
Tv98VK8U5F15puWczSXJ19WIq0bobpdkDe2XwoqZp7C1DyZGYj2jPs/diWlTJEgr
G3JCKCHpEaUzimMDrRQ+MVGshggobDtOWCFT3HZS51Wyj6PeuuI4tNfYFmnVbXbO
vww2uohziaqk3DIYYOsL3kYjWrScVSzPwvvBnXmInToKSdC5wbBA0edG3emFxxam
nmsotgevGyaDzvcM7ejztEJGBij5Tx0EUlMnDXACYt5knaH9Gou4Re32tlbxtV0m
5fYcj74TwnUIlD2B/QrMbrdx+R5PEsVGfTQoP+Gf9NKIAWILDPOFUtRKdjaoPHwS
5bGWCX7vsF//y/Gdh5MoWLXZp3T3btmwZl0CwncF0N5OGJOxFNMNk5A2xvH/AqkD
urt9KMwglY9vmqoTns0Wdlqj1Ds/qlyDZkLYu0EBEEK7x8CKsL51B4S7nQgX3QJ6
N/ywjzXHmvCSqJWmqK9CvDS7Ybnf6mo5zovEAMFkMg7ocuGiLvzADbqY5hstqXFU
3WwGoEp+xu1a8z9SVhxyItIA7YXBvk+IkWITnPoHI2B7OtVvBEk0mu3S4k1DbqQm
EeH92vsnv1kK6EvgyPPre0u+ttDNaq2p5yozPq0WKSyjM9ZjYL5LrCKJ5ZeKt2+V
dHxm55SsHSCqWbgOZhLNVdagJOWna/ZIg9yFc2DYpx0Sv9V4R2W/1jmYfJrvzBs2
HseVobV1Rm5Rlt+Ow4vL/Dfk1Zw/a223TkPE8wDUWDrJBRJZQGKFyjqlcvTIXesj
kbLija5t33gJ/a7p1Ym/0ACC6ZVtQvndtDa7vmFoSHO1J+0JI53VJDyWGyFMFvRH
gLzbmh6BI6EfUyfqQHGbJQPMp8AA8/O+UFG8LLIl6TzW/jx/eEGJ2gJv6x82P0bd
frG6TPZXQ/KcAycPA4GFxK6z4RAGwPBrZfrHLcDSWKT0Vs48eN1l7vPdMC4wrUeW
YDzQWfJ0mMGmMuZTm8DNg4xjDB9sPPFGdZnJXfUJYxVQmwAaoZMrQH9rqs+ZpAUJ
9LdMcF0Y2NC5B+l/Xbi/bKx8fHQeHnOsQaeHNrdrWhr7C1iGmlZYywmDR+Bw4sXy
TfWyB54IoTz5jDugd5kULEFDT/psKpgHbwXsvfW6SLdiS3TDviryvyunBfHhvK88
tZm8rtktbVfexT9sM/++oGEuzfCPQ5oUC1UCzYirZIycqqPOX9Q+MT66yBwkVv4k
XdnpPwxOTMTQc5Dr+9Do+171IUwiLLk/PrZuMBd3mwlem96L/W7xjVjWuT9zmFrP
rqySW7CE5Kl9Lr/bdUGVz6wVgdeq+VtbFbCrLwiqUAVm8+j5xeSp22lm+hG4Vyf6
Wlw+HjLUkoBdyTzIudYVDyO06lg4RBAoL09qw5Z/WvD28XZC5VqKMt6oPyudbbdk
rzoTwbkwYGaU81s3nB9YDa7lQ1z+13dn/soxkDcq/eYhVQlnr19ECOsEDjdf6gb5
VbosF7YaOIia/0iNgoK9MLc/ehEJX3tZgm8jXW7fSZDLA17Jqda3vkQS4Zm8ee91
0xsd9N19vYkWsf8fXyS5fmqMtBLD2BhS4DEMvR1C9xxztBJDFfIKthpqFeWIjJtg
OOS+0YZPkLT0DamLdLmIesK7PS/7gdETFt2Up+hB4jYRzJc2Eo2/nW2O5BFw6UcV
2d7VxteJxIk0y2mdLcNDAlsmVipljR/ulr9vf5FMrSwJRgxsYrNQWyG7MNjqbGn4
jyKmTuYDxzuSuJtjFrUKqEPy2lKjTDA//tqye9TE/44sEnYJ4AeQRdZlB7o8AgTo
7+NWF9OBxykX6mGgEhCypTrvIToAiG6hwWDaGlXrz+VRwqWJd6VZ1AZs7PfHiuNa
3p4/e0AN4cHPF2p+e6y5eA4onlHFst2CcvB3zvFax6JYw1NSstR3ZUt+D/sFH11d
czkhAsTpX1xRXr/PXAwzFTPxVznlQqK827RxCAm9oaZ8VR2jw/rOBuONa53RhrRv
NtV3Tp9PdmvZJBxE1LXpchzo8pbIHpYsMq7V29c/bYvzb5mYqM8JttXY3lPTEi9k
MjdUYaBa+a0Qy1Slgl4laP0bpT/qH2FvBVNRgLLFy46vDOBOd74YjQy8ROCEe0eE
bD+1vx8cQ4QaxZUth6m/g1OI32fsdQ84ec2oZlOb8UrfjA2yly+XlxBi8BUWh/E0
CGcbLdge3dNMZuADIMV7qEPqIU3e/Kw5gzCJcHV9vjVw87z3Gcifl2W1ToMFVMX2
5lq8MTag6pw1izXEmfr5i1YZd51SdAAH+zZOcOzEgxAMqjovorxmtIB8vqTuwkmj
fCxtAPe5JpRbqcPWyEddmPBwoAiSpDYa8GBir1ebFEHuzN/lBCGglmzAjhf1ojkn
fjt5oe2i0i7fL/gxJURZw0rnJ7GBQ5pSjDkpElyJCgMVvWpjoMzu7sN2FFrihibD
tXAybeSKK06USARkFMMQtc6LktuRWIQXB4XHlVMaIwruyDIll+0Rmnu+KrCOgu/q
MOb/Dqhxwla9IfrqAT3XSql0hZ+i4u6dVMH+A4PIz51VJV0NKizdkgV2S0YJQV4Q
62ZJ5lvSv/Nv+eXWpMpupQLMaS97JFB2bFSt1cieC2mQ5RRXwSxUof/X5GUHMOPu
4EHBoy+NYRwP93jFlpRc84JSc+4fHHqkN5iwLERU7ZFuYIoPuJSgwrx0e1XvWOYW
a9GmZx2YYgTNvZMQNO9mt+szRAFTsx5rF2LSGXw8WOqb+OFk2JnYazjs3HCk6YrM
KR2YKw0Om/yEtc3LinvaAmX3FcWGk+VOTwo8Co0z16zDOWEdSaDUL7aBiwbSx2VA
+rdRYAGRQ24CUxirXzCFoamBLXTIjKF+OcwSvdKrM4hdHvAxh+9O3qi67RIUVQ0z
yclr3rRsz7zcvzVAcwC9ToniysLqUu6uswbTwEJtOx1t3eN2/p8jo0vS4+n27wId
MrrgmygGt0NqW/4y4VuDSJCnbfzAHlWJKwaYOcOKV9E0grAbgTWY+xl5dUk+VFbH
7t4V7IClkbO/AM2IbDVcFkbq/WWhj/2A+943VvmAKkFQqQSzrE+n/9o2zW9iZxYN
UsdXdf1VJPEipavbrEHHIjwAFpk897yW/8exW3Ko40OwEUdy/4GmpD61IdKLiMvZ
gud5qMONRy4PZ9F1VWO2oi903StVW+3BEVHKF+FncVYiz3/pJ+Em4c4tCk8WErZy
XADZUjbB+m6TSLC1Kbge8Nw9gN79e6hWOuwE/X+4BAZgc+nQ0qJUt0TkmWr0QSVX
c4KgeK98izQXm1pIpS+8LQwYrYvJC5gD+SlLin/PziA6LqNSDKJRwASaf8s4rw7l
QKEK4Vqvo4nPaNGPH4ifooIj86XimnATZVeNZSEdq+3f5FFfIo/FQpKChKpY41rB
rnOGFRn4YwZH28sU1GYERLCYpydOmNam5765enmmL/x9i0KVKPYfH6oXrT0d1XYJ
UEnyrIWobxPPqsP+LnQr4vYtVExVQoGv5PGHWxmRsPlkPsuKDdvRNlUR6sTMDql1
2G/RU8XfZQMGtmvVOdGpHU8VR8hXLyNF261kJ6A+LgfyJcfAQFLy8RoMpF3KGq8L
YqGh2gS9SiWDsC352XTTJJhlEMEpK0t6BqVXGQM4VPk4/Rcv7pYVDgDG851aPGj4
jXKfKDFgwCNrSBXhNGioF8S3K/ffGGNy7/ezxXrXK+4YSWSdybgTn/DuwyiM/ULM
IyVX4t3Q4H+YT9yxfSJdPwTxZe0rcVet07zJ1+qYy1L++P0izt/j9D8M/IVgx6i2
dKZCcr/IZfz2YE0sAfwjUUEReygyDK99XGFQvYjKeM0Bxidtt/1wL4TW2FykoIL1
3t0eIgUp+3b5o1hXpfu2GaXiwQIgI2rQiwfnwv9T3X9tQ4JXw6usuzL5QFgG1it6
nHMBQoZe5dZk34cnLsz0Oy10j7B7k1pbytmxh1WIqplsnD40SzVusqFG6gpBi9+M
1HWp3O0BasYbMP9OB/A8KL8bVraEYT68oCgAjxCrm9/EzF7J1KnMPQSLDrrPdCNx
UAkc9CQ1kQb3tPLJO67lvhSc83oxaaF9oDWAALG8lzZY4eXq1NM3vqPufO3emzBN
/eIz2iVuwO09g+lp/plky/kNjwO/97Xnq212hDYx+Cp8bBOdA++2ZOvJsr8TYyBW
bNqYQPIuEzo1X13ZROFCgVgfM+h2arfa1rLjEl+QKjV+DUf0Cc4d8T1j8qBYcBgt
XWiez+zVvZC6fGzBOLiiReX+Gt0ePl4cmMYZVSr1r64AJAkzy7DZq1RoTeL0Xe6Z
yP055NkYVVFyxKgvh+SVbx43HusiMw9coMfH4bYnzc4XEKnjztXmgRCbjC7w4QWC
6UK7E9UoL+YzE1diklA5//pnZ7A4KBB2iimkQQMPfN17Kk4DSjvq0+i5CsfoCyM2
dsLrMQcxS7WqZwgrIUovjXWg9Z0C+zyKyaVyofsUkRkndiTCvSWFJaNylOEEB6vr
kH9LmGJoiC8MGm5x5Af+wtkNKW9O+jCfkZebZ0ooDZeXBlx1xagQU+7cYKxe6YeE
jnPK2H5AEliVO0QStvyohjNfC+wFRRu+bgr4FB6PCnzWEEfIZs3ecS6iMFQrrXUZ
Um0fGRMWjCPCDtS2eVokhQvaaTpGQme71gKf4IZ3WO/Tz4JgtThdlg7mvtE6amgf
4+X0fi1bqB9xEVTdih4wjUxAgWDuhlU7DsxaNBZ4KavII/jMzd6EXobXWinMX+6p
D+mhAmr78/COUINtXJNO8I6Wt1EAmPFX2lu/Is90vH6QtP4KwnPQxUVhJbH2DQ/m
+jhhBrddWYoK/Byw38jtxtIw7ShfsS9bpJDeW6ps48xBJZdJJ4OUbAsyfLMveWeI
1f/0YtmuN9iA/TqX57CCEQ/hyqIzcZ4TjiDNmtV+/usOyo3CZmk2UQokBRP8ZHBh
0EFbpgOG5RViqUNy2o7RthNgPCeIno1lfP7Kh5odo0j0v1h6ZgR7CrbxTM/gUx80
BikLr+eLUm3CUtaLyd1iVxvG6tQpbnrG4k0OmaJpvIbAZqOzmUyVpTPVor77DDRh
bZnnvACGMWedyykKttpo3+pEEy2TPJgWfCWvavszGsVSenfabRv9aZaEH+ONIbnW
64/n/yfnAYlhSFRetf9pQCYbVTZsg/OcnSQYioPpCSwykKXuNpXqSH9sWavodXjO
TkuYW4YXSQOaoxePzzi4DHoNB1DxOV+qin3ObpBKlchfDORESKWKzhTx25WgitNS
3avX4h8OVtqGP4oqNRbKqJC+KlmFHOSUPMmcnDT9Gb99adLHUkcLXyC1puTW8yvw
QA0CkeIWJPNNPQ8PiCmkL4HO0USgwUn0Kk1NzBnTxy7ERXX0CCX69VETfz8RTuq+
5gE+Ov+4yg/GWiTGBdY3YVQERph405EeHzMejpCFNxLXbeUpPKWupBF39Llx5Sej
hN+dnVcva08YROZSUiLxNKZu3ey5aGoFAgxm9lJqBttAm40D36XqYPwaxucqhJlp
AsCV5yH0Q2N7h3sjdyzyXpl0a4QsPNUWT6bmgNy64scxSozYVi/bozQuqjuejCbv
dEgVxwjCER8a5SCZYGckTXjbvPWuzpHpSYJhxpPGS4aAl8BHlUNlmvFRtsXkfhe5
FdXA8kAaOFaVoRWm2uzSaebfCKISuasDpH3vVPjWMSF+JgTFgy+dk4HnHx1GrKns
yTyjCW0zVmf+bexwpiD3JHGqLLuw+sTgyGdKKY+bCkmr04AeOuGhm6PFu4hnGoUM
0ilVV1T+6/q6vKXssJuL81RAPhqUUFVrF0Z+zgjRvTkeR/6brXpomDsPJNkrhNDH
iNqlXaGZGW5ZJxf1ipBcZemxJZbv9sRDvYvr8fQL2TlJCWg1wewtnzp1YUlYypip
DuaOVOk4kxT2GEEQYGzsFyTQxPaUkLgqPm+hy8mb8K9hTbqmbUVLQi6aVLl1WE2K
Y7dEQmELfjMfdmG8ESfKDZOpj1sWoN9czQ5AwIH4Oc+uSBTXtWPvSpAJlHh1QxIa
FQIf9Ew6jnYDzr399WdUHEFuYWGHld8Jw1rveXTXU9novlq65tUEqpL1PxoxYPMO
W9AHorT2r0nOQOINzZKvEPMzHmBqAMq6bVHPe6sDeU/oTWzXDcUQpMr2Ig2bW7tZ
sdyMyWTWssmQ8B1Cs/Hdgz2Dgzu5DUDzyeKgrBedxJpPLMl6BUvLLaYOhIcpeY0F
pJkVtpbFXLvAleFC5JqGxYJBPzlohkdF8u6jwHPEFcYYe8ri9OhXd955MZRv/rjV
7EsO0eGMSRVeq4lYt3rsnO4ZDoj9cOOMZCj+R7BWxqP/I6BGMtwRBy3g2dMIX9Jx
xvm2ZukflJbo8Zg30aC10j/WdCawnI1cWOAciOSkx5Pwa7W9NfRJ7sSaa0zX309o
CnzIoe6qoJXx2XiAPeDHzRnpco5aZAF7wnaQhmozcPZUyCiHmc3zd6rN9Li1w48Q
WHUTqLIZ0vcsf0fqST3C/MstoXn0yRGuXHbNa05YReyTBAklzb+D8ISh7wGO2Ud6
DpFBJsg5Sx5+TpHLtiRU/Lx2U/+ADsuUyNUV9RF5vL4+rbTLs12YgNk7Rh2eEGRE
1SPv1JTRSs8f3qmjh1z80IIT4+4Sz1sc7iULfWS/Lx9OQ/FH9F4v891qHvwt55bW
M1D+wPEOJ+n5bKpvbKWDleY6unURlI9kyjzd767y7156NrbWcEYgChvEdtRY5m8L
AVYYP1nycwcc9G/nGGzsU8k1MxVD5129luz98nw6n20/se7Q4usS9nVJIMQTGRWv
+/ThJQ6X864isEnNC0Zxmo/t1DpsE0NJaaKzDargd39KabIt1bsicxikNc+ghojb
pB0bA0R9f4TwOMKvw/haxziIhBaKyLflntCljPj4fcPpdB/4qpf4hfO0RZkoDPKK
OilDn+5M1LRrAGYnYYwY3TFKNdglJKh4RZb86MDf9/bX+ikkBfmgdzuWPnmTZ/KX
dnsjwPmhVuLWq3XR99mnxJtDesARkkiFc6mmhgFBxQZeaSDU/GwSRKU0mD9kLwzG
iR5jR7It3udAygzrKnqXS00V8To4vvuQmY8vmpiBDQjSA2EzklFDTUsyrTcn4g4u
iuzoR93QxxCJCvbeRa5pn92GIfOe+gd3Zx5Aj2abIUiPx8JiioigD0QZXroOlx2y
km80ehhCEXtY79bDT0OmoVfeRcIZJUfuVqvWEgugCPgzvmgKU6/WcF9029fSUn3j
9xb5QLTASJAlNAKgPAXa5nln4BkgetRlOd6AZQq67UwzBfvX9lqKa9CnlgfhpaXn
XeRA3VyKL52C0HxunZXboZO1SxbeS5UA/8l/6x6rqNhwfS1vb5IfDzjapSDLi6UI
A4iCzuTKf2l8bh/l+9s3X4NIrN+NlpNq3Ub5kt4gdGLrGafeiuOoksgN9nZyy2gW
WvandqIHO1/5AKsYubGMFfHDaSbVlY+mTaiV55qS2mHzPQ2FuFp5EeWXG6REJ6oE
zq39mhSSXjh/S67In86Vbt8zSD0t7ZQHXBSe+XaNLh8vluQ4J4BVuhFHEudr2Mxc
qlUBnkndc4UJh0W6++cuwWLadRRzPr6tj3frB+wp3T+xSDsAWWgJycuOSIkSRfTm
qW6eVKwraEeNIoPr/axh+THodGxDC2aSFnrRu6IonilnLqku3ltRBlLh4XcqA6ug
EOtRlc5CN+rVpsp7l7V715USDgcYzf5Fr/6bFkYMLKcUMUiJV0WxJy51zNdSoZCo
WrHAzwoN/sIg+3xB0JgGK77DCi6i7KbUcfRIOT39D+DB+TEMKtkBc30Vqt+WIZb8
3e3jSu94b8ujscRXa2Q1K5esNqqt+UanhLeLKg8N9fFKuG9louwQscqqVtPzKZgN
ynHgxXr2476iQHGvn0RCkOKJ7VHGWWeeP+naUCYnE5hQ1N/W1ranhU1bRwG2EHzA
mN+lfe2y6Ucvsi9xWQfwavUyiN0G8UAtjBlz+P4cu5Ltl73stccNNVIMK0lKUO5v
H6bozQSeTUXCKo88R61qsDNMLhqKJ124swt8YynySVAtF2fnrPnSPwjHnHqVt5Rm
IGvGV1ETJv/OEYCNBfRDDssbETZ5oyp5m25XAH76PPtcInPwcdB276AV6mTRz1Qm
xkCaSzPUeUc6IfZ6AsDllCmHzY7xxyVD0G4Q9JPIILCP3ezr8CMOhtwxYDeQcLIw
nlxucXw+j2DBilurSMszF3h3Zb9s3iHPpp6rb8jLbnTz6TxisXGZjGfe+SNJ0y2+
wAe26WMy7hubc6WYhyJu+sR7AMEP7L2ZMdPJ9Je0h7hyP9O5ijMOfPHVje9roY5D
kFNA4VbAfYRvsx9uGjAPggYy9WRqpRg79zldPNpzqeIpZ2txD7yF7DKjOuFklDj/
5qXjrZ+0M1KCrV+Iqnyzp+a1gEbml26jz4Z4dYsP1I0fMbp2rb4LMEzlUWKk4OmL
Jb+wlturtOobZe5TV7hyvePkONfycU4E8evpWwgE0jGx97Va1IHmdRwJeH+OvWl7
lSmrou/gjdrKhjiZ8BzLt9fDc9dq6X4Uh1GF/XOWUsJQ3JdqmeGctnD/2UIoP+Ag
su9kN/PiQveT95WtNHLhctU93MRMDKkco2XA/Z32HRizD6IL4kdtcwJLCg7iL6eu
/Rifq3lq/yxZKptTHCTIkKiQunJbXORFVDRRalxYZNS8ME3VX8J+1OLofyiHVLTW
AG1aTZOFjIrQGUdFdS0kT8LbCunYZtapBQdmLmVbsVhHOuDv2Blkf0n6gBgzgTWm
a5yCpyvWIW6i0k+1zDS0yVTX8mgjSYX5VeG776ITb21OOgMM+7I5jYgNMOlXtOzU
oEmv2drKO6KOgAhC9FHV7n/fqfTyGQOJT00ZeA+nEJb0H786nvJuDKoLNsvJnNlx
P8tcjCoGI8nuI54Hlm2ng4cF1rga1HIqQXbzjEOFYj8gZi3rnVFnvrLzTeaczb2F
JZpY3hRZ2ARG8S1XyKGFAB2w3AA1Zfo0ymoij5zsz+fFTYdaAkYBe9/IlRd6LSR5
gAjhfQcCBFQ34+nERDtjqZKmVy7dY0X2lJ2fQwErT4paTfkrYcNVpD/brGC5YFHy
Ai8o2Zj/W2IbPhOfFtIsp4ahuqmTjggnM/dIq4GAtYiWYP4g1FFpvc3wjWm0oDyU
Rj8A9lzuD7Iyu68WBgk5uLltmnzKpCF6dzR4iLV0wb7IWLuV9yav+pYTE/ldsJdm
Cp0MEgc8ojlkFo+LHL4zrXT0hP6TlQL9msCyL0l5yZT+99GjL6zcSPXAe+O24gxI
I02WODsBt4fCoCkhDOIbufc1mtpeCeJwOVplCqynsmuys1u57lxF3VTX6bKtyDSN
tsmtjEMBMKxJI+DqmmMPb0uEdNooD6BSzpU2ZQi38ugR1Tm/zWg12mnsfxzXLHRW
+oxBUprI1tCQ4+AiknWe642N74rlSKmKr725MqCaCiOSWUV56RWLAc7uQsz1xu4E
M7ygNZMuy8l6h9tuVCGCkU1HIPaoTo/4IstVDoIyYhChVUlWyO1gWzlyS0npUT1i
zazjnvRZfP6i3iN0p6srDQ8cABpzqIaEeOeMTI9mkI/AJ3LwAINL3Lzt02kvVf7f
mzABIHbzZ6Op7rQkKBKyex80JuWczlymRx2AHq+x+/hRCNGXtjwfObpZGvazmqpW
6OYMIDYQxHbfAtizTbZbagi+16rhOaPXqJyT7DMaHLApHUvNlL/hUDuxsQAp9IAu
2AT2KSx2BS554n7PqHJNIfBIWgOWVWtR9AGza/sP1pW7U4MlQsMatUP067s6lzgK
ebaiI+0BaKlYakJGOsdAQerhbWfwwE+/2GCRmllLr1fAtLjR85wKPTQeTjN4y5WL
fw4ujtRIAHD31n8C8CJ54SB+vL1k7UWV2AnDXkohZ/+/qEkZEcLjrDc06/artcdk
LLphQ8WtEMx3jyC9XlXARTa+F6CRin1BejkKZLg4Y7/7+F/9buof8GLuloNErT5t
zjPjxvcvaB5q9GakjWy0F+R5C9Y8EJv3xF9+kIBRSM2ELOXqn5TMHjM6tEM/iDuj
L/3G1PsGyw76nkEMj3pOyBew/XI/ThCiFXFZ6Ko+jJWiMp2Am4Vea2z+iT4DCXYW
cahvg8LbV/BZHX9+p7rOwGGZfuJaMpyR11OT2fLT3hREbPPUIbuNRgi6+Jn7XSrw
oXvkKBsZz98yC2erqh2n7U1NeO1KDZe+L5Bi5IYOOJTudDkLn7AF8x8GHvuG92wh
6Odq9gE0TTYTas40sqEgWPbXAKdUlBMNqiTpUQ5VGMJIcSv5NYNyG0S5iMjg5tnN
okGiUgOeXNbbmod/FhgNYjsEMuwX2tkrR/pWuEJnGW+bdr9cKB14x+3OmiBJQnhE
s2DZTaBB1x+feKk7Csriyk5xSbja+sMfMvCWBVFAHowH/02jEe9/AOKNNLdVXBzl
MuXPeN0hCYJbjAtzkWLRmGkqG7hrywWEwucz4zZn/4u55rKT/JVZpX1K8qXnoCyc
QxSHsvgtuE6VcYeToZ/n8FcGnM/sWmE2dVWMakb4pr5mLx9xDUUjENa0GZn+2cWL
RGHzBupz2QHH3kEUOOWAbPzzOl0Evtpz0560mlVcvQ+5xAiyEphBbPOL2FPFsYdK
08Z10/omzmUaZYRxS8ukMXXwtivkfUmlS6XeOQyYpVAZX4WAqtJ6fumbL4WI/fZW
isiOEkDwCvFjv7IJX42wWTQKuJ/+/4Cpj74MzhNUec9ggwxqdwDMbZIJNOLYWeDZ
slze2HMYRmOA9NPUYpDiJJuMmY/2k0CogWcIRQFcrbMfiGaARErpDVoOqWO2HoZd
mrbmSix7SDv63yVupbaEw4H8cXqqdkfLhwkbLWwG7YGouRCAT98rIylqMXwtK8R7
wMnosbcOrdtH0VW99kTEX1x7+OEDQ6P8FeJYdTMzmIt7SS5JXQ+Kk6XzHP8JqI7u
Z35wxjEsPhBqq0FQA0zK1g/ERcljrSyzsyJ07S+5G35Mf8diHJ6vo3C5tQOCbLRH
R2nD2qjovmMh2mY+cSa7GLsC0sdwZcR83UJFaG5HEQfW5+FsBGlDDfnwAl3CTWTH
D6UUH6roKFx+jw1Zk2/W5OmXipXPzk1lXtkTL1dTyilFAFGjnM9tNODVS1h1yAkL
7wCor9zgQIhKiFF9e1pgHueibKjGyx29iVtKDplP1MqMd1txUlHIXt1NteizUNQj
+41l5H3qQfPwpXhERZ3WCiBEjKA4E55WE2PrH+BvuyTPT2M2/tTtY5zwz9AYjdXd
NyPfZuSMTY6FQ7bJl0nVzg+BQcFcagCUylcPNUNzwMJhCI7RIgMOlGhSqT5yddmR
UUD3R829m1K1V3VZW19LmGfkFPX5TJum1OAuw+ZKkBXdPo/LFKlJjuuLCOrcTchL
iXVyXquU0NHkaVXAyTDOujvYpqN1ZqE6NwxgP4Tu/YSbSjyV+ArZFqYlcRr7iyK4
DBjamWHMRqz7MtmsqM6QUOMy51FDJMqH1G0OTSc2OjqTdjh7DdnCDq4s2r9q+VMA
vDbooCaCI5yOjJ2kKr/DqdfdimQ8G8xWKCV/JAx2jUwo6StMz8QXaOE19CxFv4Qi
LhjEMGhJTcpFWSLzms6mWiFP+mI/+7SkGvNBQaLInM4nxI7obkGWdDpIO28l905I
KM8dhhJ8ycmqISPHdkok99sM2OvbDmadqxMrY8agQE9Xg/PhqU92vtEo3eJ8egbE
Mg7Ahwovky8f+xYYGCNlp1Q66TkELEwmpShv5x0A/YlWLUrVIr2bF/tjkWxqi/CI
mUsmMvCzyzN/o0WLH1I3APbt7X3jzwkrr5lF3/VqwTrmHaSPM9W7DqdX923NN1/H
D+qqoKEjQTZNLFXyC1l/NYIRN0uamH2T2jn/KzhHWgxDawoYZgNjb8/vspZJ1lBt
YPpleewLq4U0tYKkxj5z9Dm2a1azxFSFMMB+k+iJbErbEsb+05cW5VtOBbKkIPA2
/5VxlPT3XKH/H8Eo+B6cH9Del3Pyg0Y3VDDrogsHKdkBK1mhjSm9lKzcl42W940s
+7iQtxiP+Y7oNoGZR/H0rvoQ8gvCSA+Iq6UFYIjhtWg9uG/0aJJ0tsZ00XwTDO1u
4LOp9TMKwoTt7Tyi1gfamaU5D/Jhq7utWLeR6ukydD/F6/emspPAmKj6tbHaXH9w
B4VvcbXFSTk7mky10AL3tMT43DyH7XCWvkk0xmD822hPafmPmWEQNX3KU98+103o
vdNB6BnaxAJDjln+d7WL2ikPzm6tP2muiJbncMHiXJafQ3J2f2kPyAOsrwsUIN+H
ipFFRoSf1FhN/xk5gkiSMVffZWIqxCqc/B/zAtS+qGcv3hzooebR2iF/RPVTlFFV
0Kcx9fQzDc+VA22WQSiyFzUgCxKvezmqrgh6QHyIkPGAIIDAod7bcmBjqnMcCJu7
MRR1HH55jXA3cYguP5Oi/hfdrsY5SWjkP7Zc/nZmgK/OJSCfpuE2+vmKMwMNpfEc
f7HkWo4aHQDaCnCenpn2GjfhNIEtxViG/bqKtcAEHiYUpTIor+tZU4/o1DqAzpV8
OQzHBGkxpBltKXP9nxByh/MJn/ibP04NW3WovxgUQ6RGVkUUz/mnznp2pLLGCP2u
aZN6X6Nc+J/J020vFz0NCC21vQfrv0beeoUBSnvXPfSBrgNhV6vPHHco8r/NW4p8
Jb7JYxuzjkp7YJK5VJXi37wRKJQCVih2yuevCkF9r2+CKjcAwLdoTamvyM4bbAfv
jE2GoMmxExnpq4cHAZxfiFyUKEVlqKwPRBzZTbP+KyVDCmy29ArVVIJLWFPauiPI
wguaY0bTO9qMnimpdp9PDB/wldPRjvWbYSEOZXXwr8iZ99Q7Vf3yZELaqLk/7+4s
9DdxE1hVllR8rKU868kwHqdvIcBbHfrvRsB5IlVvA60fNPURivCoPlTHZIBPzIO3
eib68H2mUU6SxLj8aXfkm08nzFerQsJGLQnuEsJDsT7sCaWvCTmknEVOmp8F8bl0
EP9dS85kh83AqLbtTOzhm65I0utxAlIwqKTE4iB6VJrQiZXRF92OWNlKdNozEtRK
rfAPqaxyXQ0ZwaCDHieG4Uv55a90k9pKu/f7be2T1GBrQ9VC1QrhU0h4PQCuctQp
cnTSSHWh+u2za6vMBoRYaMGxbzRMLYp+mkFZEoyhwVwXXASFAfVpJHOracF/B3MO
/4Bo/UrcG+OBMBh9d6zZrG8d1Y4lnWXARu+4RJefSnWhBoctBxiZ5uphY0eth32X
DNiRcGUsHSRf+2vsceWU54L1Oq+5zSNtSg52XJXDtNWSjI0yGCinW+xRG1cR62Ir
5rjKrN+UFZCSw3lV4ImB622QXbIh7u/CEAY1j9qkMsEXUnK6VMuowsVeGRNznVNW
VvJqQDYZvwen/PtwZacTY4C8enc3Rx4qNW3RvGTwB4/+5hqIeurjIQBMrVSYzmXa
D+r5+8jIMxDBZrw34EWA31JXZeaFiTOEEZlW0JV0PVV4D2ANTmZ0dGGx0DVdHj//
Tbg7x9Hc1n6DauqK7Jk8TuG7aut8HkuY4jBx7kaS/biajfsXZnmblELgZIMtUDtI
d3fiUj2S7llLEQb5B6ovaShEzhBwXmG2ZS12xF/sAUI3gMpw2h4qNqPNpKl82kU5
TZQbtDMfIEtxECLz3GntKUlcdw3GAFYyzs4owJTO2A3R2/MTBHmVSPt1YJN0fu/6
yibosG+paxel6vir0cGyZNu18DzGkM7XZ1EHqLsj0I7kmMCBW0haHMCvlRvCuhBS
0kZdC7QY4nP1SkGnBtWTSGgvITZqFio8vAU8Bh8ZjwD5q9gANHUgJYz8uC3iN/dN
WKBL+KSN+51yGzQNwQqI0JEkY2wZhZmW5WvZf0xWlLPxtM1FlGH9W5laUfNNJtaw
LAiOVd+t4sWjmDeV0M2n0Bxe/Vt060/b0JU0VvMWy9QIF3v7sBZrK1PA/Yn97u1z
EL0+E7j9QiI154Yj8ZXTOBTCBgr92uVnJ6xGjHp2msE8ef/U/5G01wRSQFA2djon
FMyTH6NyAwWKTKZQdvoXKpvUxIycuTtJfOTprM115f5TYJmxlGAOuLhrJEgevlQZ
eR4mBQ32e1lZua6fwb0dDec8lk4qjsi6SPnWTgPh46mon+HaLU1Orh9a2hZgUlND
sQNIyv7IxBloV/+LqH6HaLmvxazK7LNIinfj11VJX39tBGvcuziRLo2nZeTsLHBg
OCzbJm5ETV6wi7aKnzbcm8teeDnw4bBtdWKW4MLDIAhnhuHOM171oca5B0AU8KBB
ucc8uyAj6T9upkQ5bbZwqiWbeC0im5ni9rQ7CoFMRtIW5UM/4rRGB22TubqvOkR9
UpDYK2VcARPFM7NXtNt98XUNtQc+DflMQpouk3+3C9EprfmtPG0PmlHvrW5IRtHo
HdzT8tiMn/DYkGQUwdt/tDCzM3PgFevtEVsMhQ7pfYDxXBXLiP5U/17z6V5CWQqB
IdX4/XtNj65e7BkbhlkGXKy2H8TGM0iFHHSHZnon4R3+XlJs6A5Rk3an6gaBLt08
5kATQDfxR6Tdnrgqwn+GDwJwgv8HQG6lzvkXsE5Ffz+tkibnUoYy2H/Hwwh4x0/O
zQ7xOdjcjGsR+y8u1uhngNk2GZ9m6rTTqPI7oB3xeUBv+H6HPAY8ZwsiCFzs8JYo
0D4cgIBiXzMSH8/RVv20dIx6FMJOEMyGAER0aMMG1L30qZr8VCCj+9l0wBALtGKt
5CagaPEjl6csmp+xgE76zhNlgf6G/aR/UobNg5FmTk6kIZO8qOmyGmDBNdzUcZVj
ISQcULRySLB0Jhwe7DNYCDpK4NrL8x+5x3ciUHiRKPEdnmAwFXu0Qp1GhyK7be7F
kP98VTTlIE45/D9+9FcfhD5rnz/9Vj1qXHwvyokPCNKYyZIZPhuEVnTDu7GxknoY
1huqVNRGafqD3s5jDhZaeAhkFOXqj5hAAQNkW/lJDkcOnzL6kLTkBDfOyfhDgjel
dg3YRtdEeLgdWON2u1neZmU/OwDExzrHsmHrfGJF0BpQEm+1tnfBKA80aMy6ZyLO
VWMedaAAsRWOToFQh0U1ZFTyAVxe77wdGzmPmJndQ4IcmPBjTowFE2ctcV/0IDeG
cvvrkwKSar+EqNWs6yAvau9OqaHLtSfrDUb94iDsZraZ97OE0j4yrPoEvrUzKXKA
VfU9RX047+SBUQc63HdalbpZCy1fuJE4l6LfgBs/jCczG0UqZcr8oZvYEje1ZvtK
QDG7eT9bfNLXrh/5h+ddcW/hWdml8Y9FvCdTMItgVsmoG007NRRyCWNEtdDZs/tJ
iTH53IjPqUEcEccBsYygQNTsesuJbnc7/kVSUaPW+c17fky+TNugz10w9hnxQqLV
IgjCVjHD/DVHSveKVwTKFumMT68VrQ9rqdSR9wbJBwBPIjRWWuyNYU+yChp2tlsV
VLiMqVRN77OxCrpNUVPAs/zHSk/Gg3ZgXYLRdn+Bxg45wl47GT3VLqFTAOpEM7kv
E8nHcz5GIPyWOrd2B7El7kuiuQ4uA+g38RC/IGDDq2GPrkgkeBYu5E7pU/p750hW
6MIKykVwEQLoiYwl0zwiuvLCtU81QtKpF8Nt6SAQhDoDBBE0rgnCJncc+f8dhj3H
pANf3Hiu46iZtCIdV6BLrW/V8j/re/xNpx2D0bZk81j3r9fqNgc4YTHB3FMs9TfY
nah8iLsi1rCEqzdOcUWazBnehOuJBWV2PQjo5KZAvmRVU5d08evbzNEZMAPZwIaa
sBtJKhBTGatQRyPZGT+3YFbvl4AVdebN3l8Cn5mGZsBjVfMd5eyvGyvcZNtND97i
6wybjdRoFqNg98yZvqvGDB5c1ymLNwY6octWtD0GPT9B+49Q/Cnt1+f4TrtxyK5p
+e65pURd5CspP65XVEaCZ9JOtMKQ7Cx26mHmA47JNuqxxGcJTK5Q6vy40kNp9Yxd
WOT4mxHL6THcwQaq4yI6lv9keh91qmbOwPvQfb2aEWJJlCgREMcRSu2MtCL+DjTj
bqn74S0Gy2shEBbzliiHLeiVKqzJLqFnIUsPjzSKWlQaeoQExrtnvHst9Ze5bFGm
YYG315kQ0ztFJm+1hYGPLitLs4cXoNSKJSO3X9XZ9coYlmPlu+hTlyZyaxHYu9iv
6zxPrLI5bg6/ja8IAGCI1MDh0I5wvMqQl8Jy/aYsnVG7DrRWOmpx+fvWPml+BiBR
q4c7w0wEEsckM4BkDjhcQ2piLIkbjuzTnGHfHkfKuCkGGWm2Dkx88s2dPn+FkDzE
ngsGxC3vu7SjIPVW8r1zCYHu81usR9kQG0WeTjVKJ8BGr+zQrIF/1BfeWcN9on5s
YpIAZtglv0+R6dOGmzC/Q/ERJEPrLNdONP4bMgmpupPMZZN/YXMRniziXUgPQHOd
Qin1wGNOor1JSuFDELCKwzCcK2c4pyYHwWoOVyhpuJYge2NnukJXLcFpCKZIXpQH
50+l3aVz3S0wo2TVaD2CGtTx30pRZy12L0t4Kg5wjiX6iTeKHIbCo1abtpip5XAx
G2KOZ5iCPYHcZmg2XRbgrljWpdi2z5Ra/MCEHyiqBFc42fyLDtkJpjtUKRmw4efu
z/x74+Bn48lggXyiNJu8jL9fSxIqZs12gtIr5l/jywCCu8bbjExv/zyUP84CQYG2
6PklK3njOmjybvcgKo5zkiCOQthlEbIaPzM9r9BWNr7LW+wxh+r9NlJjHf7Zxsqn
7VoRteobBhzjkNzTH3TH3t9XMgo2mfre+JIvd/ejVjKJqeeHjwyODCDFyn892fQg
0q7+EwC9ODiGeQkvLxvWW0GpqgFs2IHhNkPBStt3C9n7yhest1a7iIQdgT+TFD2Y
6GmULvtWrkHfHtCtGyr321Ol2Wd80bQqcHvlG+A3Abk/pmwybc0grZzcToMvlcm8
XCijINg0l1v7tqvJcKFTG7KeL7ot/udkjFV1C2d4ODx2f5m3fcFUO9Lv4wpPcvsA
pPkodoklJcVWKAyePep9feClB9pKrrxywiKQsKk/Q/PqnA5q4HH1WKptVCusCtMB
Px3pbxS0qF4BBYHFxHO3ecLIPiz3T80+voPRlKB29DI60+jjD3fUlxrVUfYlDavL
jVLgmB/+4WVWbxoUJ7eKwxxPuPo8Who/n5/LX+bz7NvhHBnp9FZ+0EPsPKgeaNWv
CcET9K/8mQhCKXr8BuX9bWOFAx4e5RcqQWrtp1sehU3Zt0vnrTXB2iFDZ6hA+IYl
f8cEIKBMrtL/5iG/isokTjZ3cmZ80bVR8bX7dm11AvHNt2PwFuHZbJ3/D6WFUgHK
CRowgQ76fVHfddKMHgNQdMmYKeCC1IaBGFwOfxSb0jWIvrRQqzF5hpEXs1yMntwY
3g4URj7qmg065jE+OMgajXA+NjudjFYRGQ4MHpmmPvZTRRZ1MEBwiSABqCcekeis
ML+24uYhTpm6OXuH8TNIvHry8fe99n/6bhOaEud2LI5RJpQVHZemnu30/UteByK0
asy90qTXyVaOVNKVVB8Yz4iEqkdRv4cZl8xlS5gXeeSZbLOvcAVb9VgHDdvqRIyc
SK4MJxqh/AaRFR+d4HFIUadxBTkGhwsKfp8peWPFIy9maLMIHBAXoYvtwP0fBt4g
Aw20837xEhR66C55Qgp2BZ1evotW3JCDkE8pGYyvwwrqdMujT9kahW3zkWRjkwHM
4e+o2rMMe4S43yvN1KGsA/CiHV1u5viamgEDxAQoTXahCXL/ILIhmElLyoZOkX3X
Z9t8A0O4bwEa7KoMMo9oUwc6WQMssQhfzEc/2iSv9PDeA+gPwAwRo/kZDKnI5h0a
WmCiDLQSjPDAiaQbWT39fnf+eTzFJF324OF2EGL8KsU5KrffOaZ42HzQLn3vGHkR
8zDcooxElQYXcaMaybEz6hV2Ja8lRa8aWPz9yod2/Pgij21AiqtSTLObITUtgD3O
0fr8zStwdI79Lz/UG+fZTm9jiitsp2/6RR6nPlMHt3skvjKrDmG31MmnNeCx/TvA
PXI82UochTa9n1qun3wW/KFSU5H3mRf+apRuY6a3ifRzwt7hBseDKXNy6B9fYMRC
7Spiq2xajW9NJ2x3zO+/pII/3KdJQ8nn/uUcgGrck58NdnoMwWkbMnXFBEFR4+OC
szfvx+DNjL0ssJL6X0m4j6XQ4d/2UU4IFu8WUKNscfjoapDI0AXdwGL9gnxZTOQD
KRFAi6VUuOqKFFK0GfiBzd2ltsoYUhRvH4NuQP/I6zP+z/gBfqVqkOcaKP492VvQ
bLkrTssFc+gPe5zHeNZ18eTBe/eAd/NR7XvVsmzzqhKKVn9XOqhqcnjZ49SAnmqR
PU0FfUWC0cCLSjPmlhza1wFD97SbkItD/ILJ/EkccvxELedkjaaOPY55EGXUdc0v
nSU3uAxhtgia1uERUkUyEW2/gAsoJ4o2W6ok1dBz7Zqp6YkTdBSCgftoCeK2R4u8
tiW+oykEI1cKCQd1C3x24zHCm6KmSR6MtoEGRa0TUWqFakud0htypvtVjCb+gk4s
ChpmIETf/GYr0UvaCM4rIehV21SXBzsj8Nf7Zm7A7R+jNxdpId4Or4AYeVguYedI
atJWau+agv8XyocOTYx7hMVVVztbIQiHG7oCYigrU3SWPxyKF82DmiCioSb30Jyo
3IkVzIkDlDyKRMcDtLEUbLztZESdJPoVPz7y8R8B86vCPSMCkp7sPMinNXRZSGcP
mswwID+qbfBh+mn7MTgE8htb2/RqXxe/YOi64vDOSdgk+EaRfaNsFk+gAn2y9Pv2
4kmWyODzRYvQT4CPumGHuNxQ/aC+tCCze+cEhLDvx6YiofFxBiVMZx6vNvmMX0U9
oN2PgzjgmmYSR2ce2taVN6i1GLV20nxtrYgDkBkHG4yEPYudKuezaR62nDYBkB7E
0v0ykVF3uTZgD7U2cHMfrT+c+hSBwmaoK9k2xDJ44DbY3RT47BU4Odu19Kx+weLD
OC658zZKnJaeNZJ9udGg+q3GDW6+xOh9y2qtpg1mClKIS/BHgJ6w10jOUwgVqKvz
8Nyz8l+zJxVfC4BN0gVTmxjyJvvzNZoxSqisptOu2T4nxmon7xk9VI8We4dcQfTV
n0gxbVJCF0bukBAwo6um5QDZYa1lz9vcPWb/B9cDHYJkZX0K5fbsjwsygnpSCqjN
fOa87MGXmnxzXPLLEWNgXj01OrwsVCxY0fph+4y/XQRV7HjH33M/MqQEOUMRjJ5k
K7TKgkX80pYWa7lBpH29zs3dnDOBFmwamBJoPFHUr0tUxamXAU/4HzcbY432rUZs
QLJDKJ8NjB1ThdeaFL2feSlzkSzDSFqjOkMFIXMlUKApN7J2th6oBHv4N3eBkXcz
KXfG5glX5bRHTb17gmm2qypl5BLut2KV3rse7iyac1G09dGMQuGMSMbedxUpv5BS
rRJbgv6YzZfUwSGdznwXRzh3vWIE6+DccO2lFO8afBf9GAHKZC+7X6AwmBWskDMN
2ka4b870z/O1HBx6Z/2BW5Y3uzgFcTAhENl2fOCFSpHXIft/e+p7KNez+yFVeF5O
GTnnswK7wvkyXcuUOcGn/BDSmxSaKaoTpJLUzVYxLtmBPabxEUjeJpO77wRUEVi0
FFsNg23+R+OZpIyOS8M7RwUhOoywUhM9YptrbzOehw3ZJFzfeLGViFeU6A6M/5Gi
wsizusLRD+agHzMBcyXP2TmZcqQia9FdTBvAFyL52sPKkgURpJFslawzNUOFxrdp
ua2/bOAoDUfkDdCV1xfVsztqy9dIX7HHrC92pfOhTdgkGR6NnnvcsWRFB+nKEb7b
W8QZAShDCR2m2HyN6zO6IxzzuE7G3O5XbV/bXITNbHdhgVd86Yj0foCyWnQ8H7B7
8RwQICvCLzf2K7C7Ez/8daX2UV76lrhQzcBCDVIcl+1MuemN/7PZmZIBa3U7kXQD
1Fovuaqo6XpzkViIx0a3geKJUiGxjtBzd6+aTMyGnTcbgoYOjeIjM8ZSkOplNe8A
KNw1hs6QtYDZsH9FLOVlc2Jxrw3ZZOedS9aRdmXJLyfgYiDz2lm+6b7DNIl6as/w
DZcqYDNsM8987R+Z+PraBubBPIdbzN5DmheDrOEqqduTtVWNcCFHOyP6/AzYHp4d
7FifAxemFgvV47nU+JDlMhh4Xwkzg55jgnZiaLvG+ITC7e43uQKx7rN93bzG5aKn
cP4KvBE8HwpiUHcZvgLmjuLakR1JY8OxqLQlfk56yOsbEaGGWo7k07/SJLuyJZyp
VjSsBwpm0OXCrOo6fBt6R3AvcYCuENmS3ygrQB+cQ1oBzCQ76qu26Pj2H3MgNK6H
2dQHfyxtVci/8Vc1dGFkixAcWf5o89EhgCs406BwIhHP71rLIJ/ujkexSsOx+9Ig
Fc60a0na2lh9QsI+mr+cQulizU+rMuaTWvYmt3D047LrIdaSqqwW9jLgPyuIsWbf
BcYOo22iXxp5fujvED2F6k3VLL7kID52/avO/oRyxgF27DOhIS5yfNC+Cw8gfq+C
m4Mb/j6Nhi4NcYxGcRpSKzAZMNPVCKORE5QC0Wd9wQY8LjvXtUXWFjHehtxWhM4a
xGX8gWPh4PyWaqSQUoBnzn2mCT9QkwwYj5S/7Gg95ESY8qhuv0JB4sad7fRELXA5
46cIAy6OJCRtOjTJ1BtpH3RgQ5wxyljAcufK7OKJXMulqaL26PlwcKFX1kSS99Of
nE7TSi8sF9IK5h5S+qjsnz3hg2KF0MBsgO49u2gwEnLRrAkBNBQ8LyAqj8bnKUcP
rK+70QC/mgm4FQ1iQDViLPqoPRcZsrQdaEqipKpY2Vm3sDXK0kgRJxEe9OsUCLyY
GWJGbLeNTz2KGVuA53aroTDBXq14xHWhMZKp/FcO1t3IrtKIHWVYek+FsW0VOIok
k5LfmsqBwVKiUWM5gyaO+LtvUQ//AmZLwCOMJD5moxvalQ04qD19qZr/CNT0ApgZ
NFYIB9j6iAXjhPJw2zQQ2nrxfpiXMuyjA6l0MCXpGTQ/KY2wOtFp3RSBNUgbP9wM
GfGoEkKIIkJzY4a+kFZLXXYCECjXkS0rRmU6GujlgwVVIXZ2kQL2rIkN1/RyQpdk
vbAqz2zPtbxPhxFaZFKIApSk54qZwFC9fjtHazJ6O8FGSLLbo9Be8TQJM8knEgjC
+3JDcMavbOjypYPtnGDKJ7lznZrfLAGg2CMs0bMl8TQEPT06D+IgfuP6oXWTZjzU
sYpQpc4rb0LeLK5Vh9zw/TpbMmtGqG5FiUi7kPMTOFS+oi1dviTXUu9NmKNUQdO6
C/1T+tHE72669JtpCyB8gp7Zt7MYJi35MJ96/KRjMssVlFq5bKH9Prapn1iMi1dP
a+oFHVBmhcSF//qK5NrcbLAPiYlKOPuVcDvNl7Xhmiy8R0tQkj0nIgpQMk3M6g1m
mmfSXJKrMi4f3v+d9YHd/n1Y/QmRIhzZwaSwob7XZ0khhjIAGikAxjHqnQd8xTvz
w0z+tipcY5mBgFr0Mmj5Yo4M+vF1ALNew4yCW+V8nKw8SkxAubK17oH0aP3x66z5
7n6jLNTqh05l/83n0zJSgTPfty6QGS2EyOvyXGU8rvyTH20g2AeU1oB9Noy48Agd
eYx/bQEwItHZcF2lJ7kuxqOhkLviWdtKn7izWsYod82dDjVoodMVfRpoun4DGrLH
nYgL3vZLS7vau8C5ALpg6VX+JaFniuZ4cXCwpbphZTGEsIqB7KRg+bYB8kxREIRj
Vw1+jDGvzxCq1yY0kvW43t+KreR71oR1ymdGy97tc3L0y1HlpZolm8yVZTbKU3DO
CYByP8SVKY/1/33pm89hK5tu8U8qhDyV5SfbIPEpUuAiNl5Kv+VTUHJZkkUDS+d0
dkT9ouU7Bb7kr9WHRxNk38TAl6K3nQpKhUFqg19vl/olEAo48yg2tQJwGfT/S49t
yZNNdAu4X1+T3Pg9uVo2oOX3ygKp2Lsmdwg8YvzqPHj1S2tXQELVf8+wY/prDcc9
5RqD2GDCp0gGWNQaR1idif0Ox66v/KWGtjxL+B3j+vQUr5dzvFtqad8ZXV0i35L9
jbjJkN8r/f87Syni+anh8pmF/046MwDaxfAnIAh0jxse50pyvL/jbCP7ZBXBpCfd
OtK3Eao30AprlBogPmJ9rp/R2yZvYCgtDMdR8XF0oyVnogSQhdV/Y54Rp4OmwmnI
tLBuW+QllMloVlfvxOjtBipVFMZ+Sm2nteiGQWE8EkUK2HpOlANIzTP3yaYXwCbx
VMLVOx7OpsesM+Wv8IwPpljmG8BTvugT9Ibbk7O7krKu3ZjZoEXCf0I3wveQUzU1
w9uFzcni5HBs3tYkCFGLn5dN3bhmANWG66SLfZJOcZDSIUX903gsxykPGeU1nJ3R
S3dJBsoNzgk3xNcTCg/n4S+cahykO7x3N+Pn5vTYsOLsc0VSU232FpDilY6H4n+z
aNTByzZwYPy0l4sLyMeRPe+XToxtA646apGvN/7V+N1LK1IUFdr0UhOPxO5RfpjW
bEaNAfPqVW2XVZqPLZ3QpmzeBiGtBMvLrO1g2RUGWntmdtB305N/GP7o7XgZ5GEF
ZDgz/Si6HW+JAekKzfcIPHT6utqqoGmb8rTfF11simseCFyf7iweM+blcqPZfRj9
hhDsnPuEDf0r3xK7NcHXM5at3h4OOKSZChz+bJe3P1axpUIHGVAISFMO2CS0RxET
UVQw7fpOK+mqcilCtNqJpBVw0yw2Dd5JVg8kudyv5g3CjRtgJVKEkUo/ckBNULUP
ZRSdu94/YealSkc4aT7aXYECq7cF/rHN+yetaYR1K8/WKK7JoDQee9KyZ3RzIHOn
qkU8sJp4Ml0FqstDz84AaD9RPY6j5H2bT7Pf/xsTzLOXoQ1gBPAcqe4u8iXUDJzS
Pl3Z6NWuoc+bEwwwcSAoKx1EOlrJqFQF5ni2IewCmiFSXO3hPtDZ32g6dL1JYkaC
R24xU7OqB0RwUv4Yk4G6D1Uhtq6t85+lKiUg/0qz+KQn00WNcDQ+8osTUOgZz1Js
I0aZKLPd2o+3Qo4VsSePDBEO+8BOlg6ysqFtw5F2969unWjqaH3n4XJXNjRmRRbf
HdTcNC3Dfoqw6CbuxI7xhXENxouBpuloignAz97T8d2Nkg4MpqNLOmtdJtE17ERt
EjLGcH0Lcb1h+2a8Zpxw3WlmWMOlZ96UtqIgVSoYXy214Knrq6H+yYwJtr9WgGk1
e2px/z40FN8eT17x7x5feRYa8SK/qtzXVmcqVRAlALLljYBf08S5YhR0uweoU88p
IxSgrZtHYh2RIvKH2Qo9fJYxOEObRu4Q6BNmTbCirkEXDLl6bzOuK6Ul8TW3DaLS
zthNzBNuN12MDzCX4YPdggpv/TddJVJZI5zhuo1vSpabZZZDqU+djoRzRotcGMDV
GImjBSwJRSkiNHFVegGjweOeG33kblpCYcn8G/E5mWq5hbTANpfECvySaQ/+iMAc
zCt+CztoSD6TKeObFUHWm6XsM3jpwIMFCFPGI2XpDCj2QPvVXpUwzdCopo6xBNt8
Ey1H9rjEZSe55x+8PXMWay0fcnz2zz03bPvUAlBwGeRe8O+g1r3NI/7jHWTFDTc4
WZWqkiV9Rz4g/8ebrKhK2I7cOjDhKLTfLW4pVWBnpjT7N8CQsNEQnJrcJDdfhRhy
mRI7Gsbmoa9uobvX5BHGntLN3ri3ftdJJ62vB3OxkZDALv+TWPky7i4bSgJykKsM
G+yxnk9N/5XKju6vw4KWC6osPmGPSkMv9NHnRmqwAATJ/4zc60DfwIEi9HHSzmra
baAFXrr3bYoq756FkQVLVXrYqdZxy/NQ5HBOMrPyN873sojhaFOyY8jWU2ZHr8pj
9We/7nCgUc/Yc2mkd5cMY+A1FIMn8OtFFeTsl+XbqzSDNLgFYyZaTMnB4Ce+UR4R
sODaIneAo1anV7OauS/AAS9qwIVhSCAmsuaqBO8ea82pOAZx/eggR3s9zBtTTbnO
V2bZSWNRnNcNcfnaFjiBR3BpgMC8bHcSRbC0BGNwA5335CaXi9RJE4TyRJvZi6Uj
qDTz+g0K7Y0Zm0fDWs0bzceBX+9ayyljsH8qcYI7cGPuYGNPh3zyfeOmjfv3DxYc
ttxWmF0pbXnIpsMUcMmuNR1mPeumEGeQb4jnLsBTV8t5kn8NhjNZRoaFX9Wn7X7u
9l/KjstD8AyW3JPrcNC1fUw1hKJBcsg47Elkuh8A3B2VbBzb8gNo9qtWwQae4RfR
z9jyHa6s1wEE3z7LWWdweiVuvUvcde6iKLRoHY9RsVzkx+EsjUEz6weKa8gGH0go
RxlivxLCFfOIUwcqO4nI2MHahV9z29KaibNZwKOIbjydb90sx8dXxHknz5BpgPYz
JZla83CjYB+EDZXSFnWNPXYbUviBI0pdvoDjrtb3J1U6CKVXl8HcK3tC7ekZrobn
pUohWixjeXK86KnkMF81RRedJpNH7BsT7c+4FyR4//BIVkPN9TjAaMnLrP2/5Aqv
ecCotEwIk+oxYRPjQLwKUT48Qke4vdjNcO+8YQErUnG1Lz9JVPo2YC8o6LUp6k5m
efkWvAk7xqizrzi26FXrArcnta1sryoHOr+TcyKSDDIP89hzxv0sL+zF1aNtMO5p
mOEI0eFbKMBj4iob0pLFYh5KB/FcEHxSTHwL/KZibzjjgB6JWNx4HB71ozkUcjrg
CFq7otBoMGT2QoYJJb7RFSPUJ4PNY67gZHNiwbjgSVlYBEBOkpbUG+P+E4AWFdif
ZRSPyleaBClhyd8A/XrxveJvDPG8NGV3aweEo0+zAOyhiqkllliZORJa8HQwfPXb
+u+xxad0qgNwL2z48QxJQEEt7wmDVSDrBCOCGBisuTH5qYVt9TOgDrcuVYxrMKRZ
O2x/KtXFLEL2x/EER7475jeFXY6GUuT9u6icQ0DIng2r+PzrpXRFUtj+Wc1cJMyt
fBHOt0SH0vWpxMfNBY4PvlFtAieAh8E6EjM7iyejfFQC/pko84523uVEQump2S1V
Io7/GxZ6ZkT/zutBuMehD5QqUOQDrRSuNk8ZbuVBguDVok6wsXAjh5Iv/6p9ATvF
SMJBqmPIRoKZl3TnqNfCk8aSQAq2IoaE00LitBw+j+PmZ+o6/2n7HKPMf2ARA5c3
uwpCJJQ2la0NrZkoIc9jEvE1zSQEPgnsFCu/DbMWf/gDipdot7p0AfHaerFlfT+V
SZwpI7GogeYAWhYPvzKxNXjCBRJBIfHSUTRBM5IWgeFXR6/uHQAjq306t9oucpB9
vPWR7QvHDH305SZFPNu4cIC0P/NoVNSZL1T/TcnoIY8XQpN/G+uJe0OdfTvGRgEF
6SG8qMfd27f9Qk1sw+fMmDUJnwKce4MzbuZu8iF6BmLybaSKR38jCML4e9Xvmz5k
LiBCqxbRWJEmmxaEmnQq7bX+DA+Q0p+wlzIiktQn17FO++TnJ5PfoNW5srOva5kT
C7p0+F97MtoGNZrJ2ktAdciK1KheloEhaDR//+MJj/tFwjzBJ9Ql+f5POiQR2vkd
9E+AzBK1AfJZA4K7iXgmldJVOhDD/bmvOCADMhbBNRL7drC1fagp3qrXZU0oUiPp
hamc3IXLbm1Srklps3MJ24Ri5/BHN3GHd63iNBVqktpmH1DWx1cdFt0sdNfuQbGZ
AHLNbsaTKYrbSLqHqJB/mZp6U4SqenE9qO90b2Q5eAC3P1ahLCvWews2/CHQSAKl
XRm4FN2oMW3sPQDcwtAc381x5AuJ26VakDyFhdBh6hbZLXUrpvLeK5UmNsjYXNYF
1aa4Up261eYLxg07MPuyv0a2ZLn2CcqgfmB36YNfY1BpyOuX8NvLdetJbGpbaM47
cjmP4128zZpR/DjlHPV71tjmHRXx7NP1RGoV5W18Te6Xmk/SbO2Sa72acZyBGiLP
OtKi9ebmaHZz0hQA3PqMu/P+qe8gLK1KP/QuwrpGwzRr0B1ktcEPDsF5PX9EWxM3
GbV44/AeoyuOEg4/TesPzc5AmVj5zS3BfPuZiujLSLNSqY2kHFsgC+6nDwnI/8Qp
NSbH/KoNoItqzBTvAK8jxdBaAwuhbeW0GszLNiqlcgAJwubKop5AasNwBf8xsQXH
HEw7Zs2jOLXZt7RFak2bJiHzMI6CvNTmjBvRAWX3JUKnrlSin9+8B4URaHhGxR2O
GrPWaDVqFISi/7ECM+UiZpD1D3ntYCWMSw8j2F68mEWHzQ77AybGXE1GauEHqf9h
cs+UvRr+XE0+CcUzwshMpSTtt4367SdGDaW+6rc0eddVNtzW6GpaKibNtZfkcFrq
CPl8A6qGBgrgcgH9Vs2IjfX4N0tbyfd6diXB+HDmZZNF9i0DDOy6Z9XUqkBnVnVc
ZM8vNjbyZxFZpDAz5DzgW6Y2Sr/GplRlD7Ta1/VfFjb11KMpZI/s8+DTL0wsAM3w
jdCV24rGTMAfCjb78KA1442O1ttrc7BWn3zloqMbBjTSlrwLoUshC5RIvrMms7/B
9CkvL9pdR0dMWEKJrLuPFSeShA44fhvAOx/uAljDXiOQ8/8JomfSGk6HC30SbzRx
ud50dG33ZAiusGhOy44DrUCe1Fw0DMaMHDnUYG4zXY0/qttaC+gnrcvnzt7MAOU7
PK88BNt1CvjB85gayyoXT6ZHiWCDicDwGbo1E3m1JeiRMdUglNp1VEN0CAi1bu6L
zZIr+6BwS6+zB/mK7j9FhWcanRPqdfWTEvcxNw/MmapuKCCLaShVhAM92YzMFsLR
8LTwdhXuDqVYkRCBdTbI8vDqNTzIUyAzGF35Th/dXZDPr6PCX6TzclBX/t13sNPM
f8rZ+vngarrQbxzXp6rr9s6nDV0SXjXUg61QTplusaSZcGCRyU8LJKXwkMqvuh/P
aBAFS5fvYo/RhpqtAPX7nxL18sEc8finoFGJDe7x6+uAgSa4/2XrulNnfOYmLrcp
Swu/aV3tHi8/NzUMaUuOdg1G5KWoH8BcQTuyN1rG82HAYhS0UEwiWfDqO+7zlvTZ
Iju/RBM12jFSOwOnniXdQKXN9I3aj3xXjWE/3yN4Bi1QQwhpCVNxy/V5mAbzVRqy
WW/t7xaO6zvHhYEcrWFvDv7D7mHzn/EscPaQEsxuC1mpKWLw6ZqwtWkFm2iYs6wB
kSguH1Gy4ilUmLIjCO4xPe/oC2e8iSrarZsmhP3lYtVRBqTZRUAJpSZAZ9TTE1YI
JK0r1yV2X8GgKGfcj8SwZZT9TBCr7oq5WNyTU/zl7dCO9ocMHSWXPOWivWpG/fPj
EWZIhUIZstXZLgmUbV+wCFWekiyRQlicGskRzLQIBtSH46MFxYnAX98QLQ2t7MwJ
+cgYlyAqJ8kK9Fv9/eVCPJv38fd5fM6LPMz/drHcwHSditsEB7z0Omcjxs2l1ItQ
xkNGMP+/nJUuHkCLd4PZhZk7jRCc+N1sjUbmYCbrZacl36t9t0yZ+NyNW+lZ83+g
Cr7ftAeLZtjI1Ot6kmn+gaKjtOP9nUfcKDSw4gslm7UV83QZ7jeJbM+VBPtNKCHa
XqCydmQWCVE+bI5JKXHIiXYFhS69eZdrjfLDEWHvqrj2Aij+1hUoPk+uNdqHwkwJ
6Stk5eT+GghujEjCvMOuVTUwFgBbDYow8Y+jfno0wIeOr6zleJyP5mPBR0OzLhsB
IbvRlskHZ6FM+6HzKiBT4W4fHQWY8aojwpUjptrm334gViqs0Uak1r89ipbH9+D3
u3dfb1FVcpb0dFXpBnqfbiBYwRgnkk8e6iAW6GCJ7ffYSiRJAxShY40ofYvZ0YxB
ZDRgrTq/O7rL1XhON5tV6PHL9IkNGazt0uhyeEyWwKkjOX6vpYbA7XyAY+p0cBEc
YI8YIdTS5AwDLjAG7DI+POI9Z5XKW8hNOjfb/zTn3gVpIo5XcGKUIP2j+x5LsYYG
q5iMoY5VQ9RFV1xlwBXXPER5qNH56/TAyZ+Neyb/f6t7zpN+BEZEXt6WY2dI/Wwm
gc08QeICym687xrd8jYKFrwqucV/fagRTdBe/CpODGU/sFZez3rOa7Y8SS5MTOBU
f4brZUhaycTRw13CdeP31VU7xpPoL6B99ujhwrEKSEf++psAlUcsA/mNWnjOf9Rs
r/EjSe+W13EjX7fFJ4KaneB+Z0Ut/fLM8lvjtJPJMVFu01KInfZu5SIunbK+OirI
bp3RLQ3T07ylohKrTUvINFDaPTrzxu4RESrlBJxdzsGvjIN0WxhGVY6CCYQW2Ebl
7wTm8kCuIYwUMUP3uqsdPwt66E/eBnaehHsbU8/i8cSpeHQh1uyS4q9rqGsEx1FB
iCOJvrhumqQwUWzEO9rHpKtXyZ6+Vq+5xjAjE0ywMSeA+ATVemhhgQbGprhqquPM
N3TUuAer+6/RaH/5R+euaH3XZueXyZlWPYIl5jHnoie/QeWpR22eDcQwfnfpZpbK
OGIU/XvW8cI9Ht15nSRsckFApwQcqGADADMPz3ywbhAfpKti83OONrqmH+JIZ7eM
iO1zKPlcDFyNRWS5nZwFyLlsD84OmN3hBVASzgdUl35G10cwRcpwak+fW//PJCTz
Jtn/GN9vytKz72+Q648+cbwkcYWlBmwtdrRRxLtElLsti+5txmznbt/q1vh1NT/y
/Mbfhrw6CRNufNFg4GDdSri3skIKnJjQBYsViDD1MYX73xXeU5VEraF8hZIpslOS
oqKLUKncqla9Z6NsoVODAtSXT0gg5p5XeQWMPiS80CVLli7ePJf26LC51prTJexQ
adGW1NYKjdxIJKzNDIelEfxtHLsTRQ1hl+WmYUzouORpLl+k/9m6ue2xtMvk1rvn
EIP9TUCmgG7V99bI0HEf5oXnoPg18acP++Tmoj4wO5qlm1ggX0wkJvhQ5da1isPx
SL9fWkcjX6UhRl+31o+5W6JyxUnJSNvgipLyH64s6EH6yxPJexQUakuo2D0MS7Am
CVhAutod1vluTAdBuX2wT/LDcxMd90HSBeAg5y3+kBHAg6zUQ48RTAyyMPm2qVM+
qd4xKt51rSRnBmhJmH88RFWL0k3c85h1xsTTU1OYSujKnDV2lgI79DngBGcqdp19
YgHBD5+6vMWP55n5uJHoCxLPkyFm9nMTVNs0CwhzX2hArnKnabHUqbHLPcU0019G
gFakPzaZ19BCNE7PXHTPNjQlqqNRl2dwEVSyHaUWabUu8a4UgtHqpcmqri62hHyl
1IZbsNTCezOZs/aiwCzu6X7cBFrRi26IOI04dPXkYBD9+ZGMrWuRphW7h0GuzPNV
yqVPfvwKwBZr4rSu1c/yRaB0eCAdhtaeYDzcTycowljqqx/n+Y76lhL1BBZJuCsF
Zg8xOdF44QjxFeh07EiCRMUzLrHfw62FgUQVIjhgCEqbS4i8krwFZyqSlFlrKjih
GF9ZoMShxfwq1l2HFwnIvQ4EpX9zeSEUFpWOZQqi5JLyVX3uMnlqF8TRT14JP50q
pNamidHQJvybZrZJlUzYg3tNckHnQ7o/lhSi3un+N0OWWf/SE9nK3uZLz3/nYdO2
KlC0tuLBB+8c/5CSUBRzRorjs+3LCU5I2uK/Nfq10QC49PcWUgGxiFU+LxJcBXHI
l9kg5a2VwGAQU88pj2g0hR/+k6u6UdoiKp8A08QGs0YuVdiGwgKTV9Jv2/CkJiYJ
l2rEV13vvnpRx9UwkPjFbnUMgeY11aRBS55UN+eSToMJJSRoL11DrY2OqJq3GaBb
ZamapccJEjADRe9xk1HSaZnVkoUjrJ64u4CMJWl11+UerzMC5utWziRVctflfwxV
xhWxnOiRUnRd9DEJ51MQwPRUq5+UCFziTgwhK9KqEngNckNF/6887otAptj2l9YC
ywMvFBVALgSvUf+qvQQBuHrRNa+Zof4pnc7LTd1VvC2ljq8lUAHKZopGkSvcBGJh
108AOdTLAydsEe2g+SuHgLNgthv8yCVcBCei+g6GfBxY1e2xBBUUx/t1ee1YZhLU
2CW1KD9aMZYOW0ODl5HO94iKssdebgbW2MgRdGMqYu+WmT6XVTBQ90cujZMwzMe9
3R7fLCBFKh/boafGr57FpBQoiFajMPVI2JFLoVd8+R0fN/4351jd2dCnqCUf6ij+
jSCvOjHSytQ7sDB/n1KP8eeteEbYKfbqsnkKzquy6QvjSk3HAojz0H3W4jReT8XQ
qPI9H4RcPmvEjfaVqwQfbmfJHFr8CcQYr+4xmkCQ+Xky2qT6QnK3yvD7zJIFdDAU
aVos85LJAnoCxptD1XEfpVErWE2838cCh9SL3beA2cYMFc2mti5AdHkhs+EXPqLx
5Ve1AXB4PrjwPlBrMt9fC6p8yWtx0Uiq406ZmTP6QmcvZ3uEfDhKztH8jv3Ai4rR
Z+OxIFVzIINimklYfISJ++rLJmKfuIYNzBcdb40LpxoX8cHT3M7+E3lL10x9Z2X+
8Ql+TbFjRFVG7WT9QTl3VwpIFSe131UmaOmHKfcKEcF2Yy2F3GdDqAcsXN3jvUn+
KYpcJv7yef1Orpw8WS+50L9HC7XvXN44nTEKzYmfJHfvhe51eZx8yl0FRWLnIF2L
j33zMe69GdEyQR8UaA59fFwEHKAbJU7cFoOYkJY36XG4pp0aKoyXNgidbsG1rVLB
N84gwshq9C0zJVEcg7MPmbNhnEa237TQ3uvMkS04mSkx4bwVVuYSqUc7VtQ9+CjC
MoqlrPsMh7nuYnhzQ3CiG15umRMQuPnv4A5EHGvfn2JoQXXwwgHUviFXqWr4gpKB
IyEsF8Ms3a6lCnpOwhrUwSnZ3HcTUzho+T6wUtI6cLizTzFD0/YuGAN5waPAHNvo
JR8fxvYVuyLKpQ3TVhGZKFZM4aJb94aEeHYWvbTTNRulC36jzs3xzhs0Nzb76xer
pFdeHxVA1jiFGr1s2GltRu2WV4TGSzmGiSf013NaqT99lbmflIFzaHDq8Yn/Eks/
H5N1d3aW6h/RnrnJ4buMcVxo9DaxqLwMqZChDFSQHyd9+QKAVdVLHI63c2BtQS8+
vQ3cFzSM7SM9f8jArUJu+W1IAn3C2EpivLOuJ0FEDrmlGS0VwOMlJsZCAxM2KViC
b1ORP9HTWPjDwwjXBPuKn1xePBCjduzLVN+TmPvL9JhgGSSBihskii2ikmhTgdxQ
q+aL0S6Eqkr36g50UsD6Al6KigILA/VnGSN7sD2p2tqPDe0PNuIV16Qi0HP3z5FL
xbtEvFOw94kKjK1pSYd6Bi1UUCu/2Jh5DS44c1LvGqTJ4T7qWOdkfJ1iil+pzu+R
q34FC3sUrMrEeSUeICTXxQkuAAVksI6gbPB6f1x8W0JsqodEgWuBm8RDWxthhCe1
ev+YWzP1ntDhlVqEwT8tkzJ4Xa5QtLMzP06nMTABEYIwJlhbyckiRfiFjPcJALdO
3UhT7qB92fq0PdZyauN0uSlAaTGVDtLQ0Pt45eBiNgfnBJOmY/55PVDILjMsPybJ
QMETOYMWQsW5CST+k0izp7erzplkVqqc5SB6i4UaBMunpF21oIsoLLlmaOAiWsYx
jHXsYtDk9grfGdPAY8MaIwaaMqSMHno/QEG0ARLffDX1dnC7RlhedsvTn/XehUnV
dnYEYQ5cACv+PnP/5bvg7iUUEgoN0MGJ9pnfewoBiNrplcdGYWLAqNMI7TpxSDxM
o52qW6OHbIa2txlpLDz0xtq9kCiuqvi97HxES+zhC9IuZY2/a0BgNUspXworKUyK
/voowmhyr+0J+bf51lisDw2EPfBYUdvG1jdsMO4UZT8hsXvmVPoy2XeYM7XfssFD
yT7iGJd5TN/+9Bm7GVjLkETltZVgm0wla+tdJ/d73Gpn+tTCPM/nSZSGXwmddeCA
7WnEKgDnFLM/VUmnCA4Svxuy4pX8hEQ09ihAZGp4jG4nfnokVCOEleCLjq0a//Mi
B6l/uniVXllZOdpjW7CWOAy63/mOBGNMk2cO/UHtikgFI2HqtBkqhClhmcNhMVPm
DT+vvl1J+hQ8fbZUX6D5/pJEtp+SZ+Az6r/y+DJm+Dufu3Z6TGj/Q6mULGyzbiz7
sGAJbEjSv5WtBS8TiFXMma4yQbSQRKGvC2y7LypfqpHJjdjHaNg89+jrvGd91B2K
SjlsfeYVNY14iQTifG33y5LWFXmuYxK6isfT4/GWTZ5ybeY8rHdTies38qvC4Qbl
wXF5BDQru5PcfFuIhil27/ffILCS6fGcTqX2qRgx6UgcTnKrVrdhMnDToD/iCTE1
qu7ZfyrdjtVBQGHquuJPO6VaFautaw2HM137qcRv+Z1Be2ai0jlUQVbFXAs9OUYY
LaqjSzwH3jdjE3WuZ2s5YnLf/KUoonpUaJXAHJeDpOTaNoGgwh7nLXytueQ2khi7
WXqHkLvwz5KvkA/VMxsoM1+zimiRLgfnj33lbaCeAkJzM3f7AYOveDybFbpAqEqd
20V9BPvXUxd2UBvQnWw/GBLhhLuh7fvKe8XbyeHkNPTQ0eiF5SVPNOKOcdXo7uIy
8zy0+JPCDybLCONgBMoYnOuK+rTqvLRSwYJ6qc7PcUsFZ+bRcKn6LPgw31A48UYr
Ox2ypKyjDB+NUNHPqmXVM2Aojm/ujBxSWdPCpR2P1xt59n7MtZryd9vqvfanbwje
GMBJDclsifLnChyr3N1Y5zFSPVu4g9oqVDn8rV7cZLKg2VMy5ujCSCvdDY1o2Plj
BtStJS1IAbNiNDEI6zepFNPKvN0mySLpXIQyCS/cC+BqB1NN0l3DisVgNH5ul6sP
J0Vnzv6eqygOXRkrirwToBkp7nKr3f5dQk/PRp5z/maWTuzHeMjc+QJMVQcYrp6N
IYBjXJ7GLw3FP6by+oFVLz40x0xLBbwur1YQ0YAeWh9DAIKjiEVpIeVufDf5Jaco
f70bkLiBWkJQM/W+2FfWSA2R43yd7yXRjXCHv1WDzY5B4O9vqjDNd/IPz73+pc1b
SEqerBm6D4elARcntWWXooKv5ZZZFlM5UnVM5x8WfnCJSvA2gFw2iHh9m2wNijsq
b/tIsgN72WS604G0KsxKyPljWOvkQT3vMjvcRItohxvqs0YA4EECCQErdpH2pzYJ
UJNNvqZBiQvtCItEBXqxDWx4QQ3u5uzkyzZqDy5o5FcCnDBOcsUdbi98F0pycqF5
n84tZHDegnbFUox4lFElTNiV+aJ5RuxDIB7XFgHqbftfIHAtbaq95mpPNYwECKhe
GaalA8NddCcPtsd7gXP5uD3hdEqZt5zi300W11wQ7wEwMHZjQJ9JC1LRQ/IT3SzQ
uYubRkv2/EEOLl8CB37yst81phyvTRP8TGfhrYSpiDbMLz29SIC3yV8L5N+W8a+z
D9k1kVae7Tq/b9gN5J1mF5K3RRhzsV96TkgX61753B0N5DOYbxUD/nySYszINP6D
H+KTZy3usqqVJyioPxXsMPaQqVnJo1Ke7spTl7R0xIGH8Mk9uxCBI183nShihgpT
tafc7rIqL9PyikToWPU6ECOawRF3/DgBjpcie7o0xMv8tAfqULzo6iWydFUGhagh
4MrYQJq8ff9aFu/KWoD3KJZpARjrehpd08m/6vcetwULuF7Xp+xN0MSatBLwVI5V
V/+l2epkRdcWCHbKsmxx1/Pu8sdyzGlk0ZNn8VsJIPOoOand3YrYr9IhRBDbbucK
++QtPzH4RhD6nPTiR7wI+z8ZA/Y5se/fhD5BEcKOe0tr82XrRLDls2aWjP4Hb2ik
i02JgrMbwxb7gPodwLae0M5KeJg8p+Ue+M79Rfsj+G0k9sNPskcjkY2o6dEIHqek
4VZNRPiFgLl3Ru6lMgzv7b3OYecyQorTI6bNp8ucKoMHqZezzEKJUV5k9IQzpq8p
J2bJSnyBcPKa+fD8zEZxFpH14JeDcB6i96dXv7QGKymZYlWjwou7dFEICrLlB/+j
XUQGNDBjF0asDrfvrY6AixBcMDoTQEOrIcdDdJjRY0SEdbzrHxdGIV0wRWtnm1AG
f9zLu09JRwXxXNtWOGu0uQlg8WhznZGzzEUDXpeTYhzIuo2bnFY5yZ1uk2wI/s9A
c3xE3skLrrJOt5/rQzkSs0FzF2vm4KaSPldi+j3srZV3hn064Vo7GPCbz+I+wAUw
Bwjel1jRH++rUKSy6jZar9cX00PFCZ3lJli+wYe9SVoXd1zmHd5PV7PUhe923ect
fPDyOhV7FuULtdfZmbXsYrkNQoFx7loSbVN0NpwrX5adysI3U6jBOZ73uTT58YPk
Sx4h5AY1L3pBWxcxJc7RR9wQTqfYyQ9Rvw+8UOv5YNDyInU4r2i+VSX0zuBM147L
vSNMTgp7sq6+A6zhcn+oOLiPkKDYQicxAcoX5EDu6r8a9uL8AxMO1wEL/xZelFby
lRfSuxWYZoa69NkfTGsl6jJ9+JTyfr/8R06wmrj0G5JnBFSwyjvOZNBZnHU+aEnp
NoEOjwwtz0Fsh8ItNBceRh1uD8nT2H5SBnwFGPlabr4hzxm7cfw0GEcP00YwaLMf
skCP7YsTj4anZn/yYbfpn5htTZpRP9yeeryRMFncR5mwHxhZOSTdStW4VUXmuY96
lQcVx4D7P/5jlLZCHs9nZFSjFR19fYHBm05uTYqDL9Kw5tr9awdoMcbFf2Sq8xRd
Ud2kXlR0Dp500lubRSch3PATVIfZXxjj1E/KUOEp03qs3aa2KkPZb+kGd6PoGti0
/SBj0d+wjHCcvHhrcNP6gcCQQ/pEL8wmP1pOdBvgfrKlCVpOOWl+dMTAUufrew1i
hm9HWEcKywnMT3MVoGQnm1ywS87IGTTUahv0c5WY9N9O/i+0gIiPF+XOo1MY5Ypw
XWNTahhydB0pDijobgd23lwjwZ1pt5+JWD5NzmSiGm9fvkPMxH4VWtjI5prvxOKR
FqocJWdIQOhos+IqUP+qc6fCRd8ugM0ckbSmm+23PEYS27Eais5ZHC3VNrIhVGkF
aRJ1tfXt2bpw6XlAsuF9fA2qH7Bl9uspUJ4ee086V6ZkpBO3YYmU4cCvEaEF9v/5
Pzxjoh4JIZS9CtySOmG8GUWz2BxgY93l8nl6j8WQ4StK1uWVZlFigbdB79uXii4u
Xn3eqo0u7wfpH38JU6EWZQwsQxqHijfslz9BN3TBHL3ibpXWCIcZAfZ0jJB/DqrX
tqV1I6d1GNEpgfsEPmaWkrO9dgY2vTPSing2TxFZG9mvJnqLibC52wAsikhHV5yz
yx4HFe+yycFNHNUtgCCjvHLqszPrektVeC5W3DEL5gbbXJpzCgX+DZF7MZnW4JK5
Uli/faHncuwrixOTYgMFrOz/5fBsFK1LkLa/QTmBf1wTY24dvORlmSCys1XSXrNc
diSrVNh/Qb4D2hIVq9b5wPmpE7jCkGScAH9HesV38JGV/jC2eTRKow+RnGrMmrwT
kiOJMT5lHrej0D9dFEZFOK7okLGM03bnt0JLOAswPNZV6jCc6M1+a/xUUJYD1HSZ
p9a+ugUmuco4b2uLyGwt3CJv/BemjlOkh98NSoOsq7y5Zw68gb71byu1cDNx6sJQ
lVr5gV7v5K0cMMeUkCOY1bt1wN+vSD3KtTa4UTsHS07LbHUfn0OwVeyTs+YkbAY4
djy762t9BhqokPMLxj1g65e+gIpQbpl+ex+LWayqma7obzO6GwJ0/ocgQkHQLEJM
TwqDRuhxVtx4jvXnbUFzXsEBl7Q+V1NEgCAkIfhzwyCLYHj3Txwv44RWpdRqSJyV
o+6ueHJJenxmvQpl7UpZHq5wGqaOFCCJ8a+dgGqq9KQrzgi3RpLe8FIw8Vmwme/g
akA54l6drqFbNaDUXLVNXFkvHflrlsGw8PAOkeGpCzUzKtr/p+0+7kCWD6Rq93ay
MFz00GUJt0tJrqYCw2GU0NkFB+ta7Gdf9TY5jX8HTevV6eJuDUUN8x58zTuuBNAG
zw8YagAmqnlSlv0dbVM7RNNs0qTq/1v7qy2y88okLsx15ckwgLXPGcTtN2zxzqfg
R4q3x9F9RMgrdX3x3FtMODepJ75VcihPgSPMeO7HkiJ6QJAsvhbPD+cbod4qaG7X
c1RyY9M0fJULkyL1lE2wQWj9E7a6/hf09V8fIZSeRAJ80S09TL+By14hEYbRlx9M
W0CAaIX7VZDzhbhaEnjnQmR7orvDz5Xx+bXVkEicxBcGNQOEvFvGGWcxngoqFaX2
+DT7Ay545FajTce2bDVAdpVbzi6WeVp8VH1ow2/L5JzA4VnROyL1vSq4ut3Oh2c1
dzQhFDrd9Zyfz0gD1fjdrgI9uT4U/f90Pto0QM8/bdIFtWYbUXJvsffUzuyp94qe
JM8PuecwI8OMJ/h8Zk948OdxVm+4BsgxsvDhit5FXC6Eb2IHikWtCDzBGT5kbVPA
LSxk8Pwky3AORJgRp6bjt97MJb20rWctI234xV5k1kcrwVV699p0CLkO5dlu30yZ
QEZRYdWWVjsfXkBF8rCNzRY1whFvfNWIKVkICPVajgi+elFdjQ3zYkVlXyJI4gEg
woiRttkj1NAZb3i5XO+/Ug9xZ+T9bjrNodZ8FjKp1loAq053qCL2GEGTtTipzbCM
WC5LP9naJGzg1vzdlXDaB+bJk4o34lcvP890/7we0uHwAkf5IQz1ZJu0+AvthRiR
uJVqUyjlLefVl083XPSO+kMXNLmDrh4hA8uc1LwdzXg+Z4z9wsPd9O1/9AvQyLb7
hjtlyxBDofPq0Sx3agZ5lu9xriGkI/dkjFZ6ToQBxGQI7sMYVNvMkoIjdWl4Y5bH
+WaRs6W3A0K88q/y0WCgjJKUAIv1K/Rg2BFl1VgUWaE79qPQbkoKixT6RWpU7hl7
IieNE+uK/Mo9zDRZY/cnXu/vwkOAgJb445Tbdt2hHKr/EcmdbXYvlAgNje65dghD
CI0EEVhVtbkWng0C23CSKu0QW+1N0u1eh/J7caTUFAoz/TwWwAp5YemjRYOx7ic2
JtJQNYkMxuJBnGryh4O/3+Lb6sHJyf4FYC0oXnM8MB5sUeNvMvn+fekuKfuzkjAx
qQ6M65vZUq84zSZ3rrHWrVdnIKR3zNv69fd4Es96uCJAk20C1I9Y5m3AAJBvlcJs
GIn9pPwN+H4/jxt3gTlP0mOp047Y7Cbrk4841/18XzyfoNonJX/IrXkVUoGe0ymb
ZvI4+SbazZv3VXSpV+wnHExAuoLnuroeClm4mJfWvuLQzDnNWihMHZDYFy3E26It
isgh5ryvyijGFhZJecMqtYyGmiB93mdOY/NJ998cUgmSQD1vXmPL1HV3UOstQbhB
A+V8kMCnq71YyY3gB/6N3y6r6cju/FWk8xHam6GPG6N1cwcEpDsuSo1ugukLZ86q
n6Oqj8Cqpt3jdGGfIgkUWPKfxqou6vHmTQ7Y8ox8KSg2ZRDW/0dR0RXzhUZTrE72
5eF5UfvDjX6oVubabQtfJMByQyDOB5Dskg5KJUooPHgb/lL6Y22u4F1mGJVnl6+E
/oBn7wsE8G6JgQn3WfPxnC/DlKfyzD4kYGpNf6cYvKphSPrAP5FghDmR3DX+4/wO
f5TN58XwuUNwpcBTMBMugyWH5kEtgcxIgr8ZifpB3LS0tomRcWbcxa9YTxY8lACk
i0Hd7K60Nh8O7mkO1dts0DFNV9eSgDbXZAD/lJtu8k14aBTti7tOI6OaJVOULR/s
TjpqMQBaDN4bDq19Qk6SEIQ9usEyprLNqGlHtPyUJ0IDgju9KIw8BZeUxbS5p4gB
m7V2Male2qLbYHJvwj5dk3OgJnWqh3yq6Z433QS0nGZTbfnR3Hu4r9cBIiKjgtmZ
qToGb74DKEr3Q/4UOb4nmuUQj1WeHlCyivPVtZcZlGKuqGMRkyThkVbE58TQjn+m
JFxPKh2uH6TajtXoUbSppFOjiFCqrh2DX04bLkhQe9+y4qigD65YiwYiZUVy8lUi
RnO3wEryCTu0oDOwxdnxAcFZeU7sId0y+/QxIIrmAgWf8VUwnIy/xfRhQuafSmNg
oO8DsZAjWPHA1sJ4YC2C5dQIzCqbzv/H5x0uNCfoNio2wwTYfTGH1VYT6PpKg3Ce
ftYe0r2k1tbd04z4FImbSXLfP+1A9pAC4YFTZmAvA6YGQ4WTjoN2CIJCAbn7eVzm
L+M/Tvi9FodIxYJlREesZ0+HlCauXjp+snGIHBzyZMyOD8LR89erbWYjA1OKHO2H
I/a9vqhDA5hWQ5E4jTmmtS7+RzrQOIWcj6xLnxAZ9q0TqPfw3iBpl5/VVQAR8oz8
SIugBTA105fcMktOA4L+rXOXlxv1ZNMpOi4eD33mtdAZ5N89IpkAbPMxJjO0Jglm
//sNo9UoLe803aN6Jl799NIb0ogvWjY6f+1NghzzIAQw/8AnpGUor+9Pb2JbKaeR
f+4CulFSWMft6MrXfPViBWUvd0txCpAiLZ5t40k0ccVIwH0L2bIrhkg+xIgnazbQ
B/RXVwtyzyapaVoNXJ8pdoXW4tQDmh7/o9CRm51TD9dBG/MPaORzRo/nkeLHVBFw
44ZIWk93PAyb9BkDKN3DOHYvVVcpNmHMoGZwWEcsi+6ggVg0A6ZDVWiVCDjcEZE2
tjBUo4h2FhDvjqDMuPLcLxcUovs2WYp5Q7BkXtnMQrfYyxUlSDkH1Yyytsbncdzc
UHvWIhHZ2b/suuas44Tw1VYcKI0fHrBX2lWf3IY3zo+pxvqplQZuw+jzP/JdiuXc
/urB1kBdkrbr3wQgKPUtZd5Lzyqj9a5M7MNc04fBzBQJ2Jd8snDv4bjx58+uFFI8
l5Bup6fLTb2Q5Z0i5fs8bDENPacYgyOpzDg7lCpGGQx1pyeL6rEz0wC4mmIzxzN4
s011hEIvPNrwIYPqbfXhATE8KTS7ZGYC1rW53+ugol89G1rxxQNWWIAnNya1b9bZ
dJgNYylN0KeySMhf9DC5W8ZcvWf3qMYS/adJJBBEVfhmlRBm5+Xn/zQycDiEdNA8
aXdzPRzA2ZNh/QZRsRg5/BiI2GipeD8fH1XESK/v0tKc4U791d0FL9Q+9vxbaOtP
MseWIAQTNaLevHvoIP0y1UzbRiSX6RXCCMfFX5hrXP7ZU6ZuN/NssM1C3VYvL1Ey
WgRnLkxja3Rk8elROYVFTZ+I5/fgZkcPhnhGh++Uu8O2dIu7CDUuhOl3o2bTIepE
F1Ui9zMO/PfRgOadGq6VyD3bXPe+jQM/meF6X+NBfZr88K5mjQ4sXPonNjFTYoO/
W7HdRCYTyXARnOdxcAfEtuI1D40Iqz0JRw6vYk9NUTuWlNk7atjE9OgOhHq+fvSV
3YVNDTHPd5Uw94ut5u+SxUQ2FDjAFYLEVNOqdkxiHpDP845hlkDhMuWcMUi6czQg
PZ1n6Z/J0vzWz0wGgz13Mpmb7Nbmsb5PmZK8VLUPj4CLSS7YW43/8Pf0l/M5xepv
ecwXYZcp0UYbAQ1dQisgquSFX4Vycf5tZ8bnvAJepdZrPFA08xlQ7EwMypP9Zql9
MJm9dJnSWT88fKQ70OEWuze5mUKPKCasTYGlT1GY/FcJOzT8fviDJbzjYn2tm5Sm
X6o5BhSvPdFUOSExMatSLPrDQKLB/NhcyZHlDW7nt1pSfGA77ru92JjrdmakknBK
mguQyVIhu1v472VjfTZnSrfcFSsrSSe3z/09taWUU4lnWg9q6cgnvNPzS+H62lF6
TKS3JpsXIrSgtO1Sz53RGwhBMem+MurF8FFW+kipE+lUAmjdgQsA9hc2pGPMabrH
8oCaaESWKzijWRN0REVAtWgDBFpFDEzhJpYUe97ap0M7g5CoynDxRbuva5/tSy3T
jG31oScyQHXNGbelaNAspdGUSxR94eeVzF2PmBHVMP0Ep0bDrQjnWmg7Ftc1IutM
J2K+8TM0iNUkj0d0IVWGad8rifSa6C9zF9qlh/ddAuRs6L+MSkkOVjGppxV8u7rA
RPMVrARfaAwPUbar5d/bkZszaiU73xulaK7LPpEIADIjKp0qaELaJJ+qJfS9DqWp
PtTJD50SjfbMtb2odtBqbr87k7U+VnPCzZOtQxsSM4Mx2l7JC9EgmoGxFGwlll9p
KL+s/NrZdY0KSR7sv7atPoQ8vskRYNGCeWTaqQ8ewVIPIore5JPbSV9WzqhZE86M
nDRIMDC+wg95+6S3+CgadOlnLEY6lVfFbS8ye59kxYuIEXl7a1V5IVAQrRAKHauK
ecK2mXfgbdkavGeT2f0gv+rsJ4kmy0f2420ifPDgAAHIzmWnzWPcRj4C0qco1JrT
AgVZe89P2xhTVw4CYnu8wtnY0goZ1PZsOBynxodNIboYo35cK1PpKlr30bJf46Wn
tofFMviK38hmQ6S3oIwzhjYmtHn5mYciCXRqknIm2kFeLQBXUenkqoWGUNr78Nx4
dmnN8wLJmHsTshGwNRte08i3SeUGgeT0H49C+kwqv3rb4km1ZSFHigijxola5ANY
LYaMraQuQXVyHJLo15Qo7YGEmJajD2Kn8hQuX5I1hsQenmD6H3gAMdrRl4USSVw9
CN2K+0Uft3iSckril8EtiClB3UjpXFtbZJCvr9ag/k+/rdefEwk6XjMrgZSOwpYB
AclIgCbA6OQ9bclj/p8sDd62BR5VHbPlJJ2AmAdyQEhOTO7Ijz2yObJEjyvi1Uf6
1alz0ei8MryhT7Xbo+pf7XomX4cqt+duPvBpfVn58MP3cObgATDVWRtUz++sCDUh
dfw2WTWS0rJaqEE3Rl8fmGsPEuMNjnFLeY4JkPZheEKkgAoygI1FaTuHnMEgovTc
jqMdDJtrEg8vRC3ifhpsRIs3Qmcu6nkDwOi9uQ1V3cCqRhPRsz3PcAT2xLEjPTIv
q1n/PwqMfeUWmeh260b9h1z93ykdGBLvCjJJVPeCJ+WzyumLWBs688HXPh25ho/1
WQaSNALr6Wxh9trqJSu+ZCRJ5DHtMcpneV2nUQZVmbBdNDrx2mq8JTmdMeNTntcK
+DxUKZV267c8eE4TewCSwfbi0XYi7X3Bh9FIzhW1t8kaO12famU0yQFa6Sbs9FQz
DfJbyg+J+/vUfN7r2jSWbLL/Gt8jhihvt16xNHK9r2Ceo9KsetVz0YX6DqRImsHO
fjEW9GGiVYJmJRqvijeoqCnrSKvtu7Lg4AW4f3TtpbSBrw/GJYjh+AR2WR5E5HRv
BpxMtC+5K4VqT6glLWSAe9DPF41yHULjqPnxfNeSmXx+IfYlvI/FpqR59SDNIp13
WWAuGmYDpkV6loIn1+RAoys3bq6zPL66MCzUGpWQ2oviYA82zw+p/eXwYyeivSxF
v6QPjA0Vz17efH8iK/hvpiKxmsWFwnbR8yq0N5fC0HnA0Rd7BZZ6VhcDmmkHvqJV
Q3HJYsi6tX0kb3wdUV2jfoU7VXPxIuM0Nc/MGGn3IDcna1BecvLhmjGJYOT583Xn
mxukCOjhRwx2FsE1Cn1HPd4a0BXHO0pfEQMjk/yQa8SJXgUi7LCtrsl//fSWowuP
BnzjpoA7tCU5lH98Um2Y95HeXxjzXsZHnhgLdFMn7oWepjJP6Hbbjatncrk7COTM
v+YSmB7ycJRuTxlfVUoPY+beq1MebmotSImy/Q3ckB+8MV4p9amUrdLpD2tcVtm9
pIIOdSj/2+oTiP3+yT61+FbfsjowD1esIvp0PhgRYO/wish7t0pzfLeXxu4VnXi+
7Rq6YBSiYbCA3/JLdP5IwNrQxG6ucH9E6zOcjRqkWRm68oqAvXtmSSuEEVgX0K3f
PXK7ooqE3Q5HvnbX+DV292sN4vC+xrrmFyAYUcnZs8+AG9bFidTfP2061piu6vfw
TMP91GggdIrZRMRmo0z5oqfgHAByiiDgHxX7/TczDS4SfhR/0T0BE7bgNNpjzVqO
8xZCtfySdc5zDcpug80r0nIpaw7J7IHWt6OF54CAmYQ9vupfJkzf4/g1c/Bejtxb
jMayXyG6u3MGWCj1QeD0YCsLhvWIJl9Fp7KkN4sxv/SwscyqfQlk0fUbaImXHrBQ
mSe16Kx4BN4/xxHaMqgM59rtTVeZAMNmcmsslj0fYVSvbl6MxE+Ho7wpi0QmtWNU
gmrvJr5XLre4PfPlnN+jBTngxN+ez+CXOXWXAsmFwmEXxSO0F2PPct50VuJrpxi0
LYnT0vJ19n51NBH8SFfVVsXbIDgy2fMgUEW/hV26mXvgn/LFFkbKNCCHNkOUbuCT
fqe6YULnaSuIAFDbrXK/2pruVfeOMLSGD4kGsbx9wmmHmCK0R9is6LMpaZZOIrt0
uObKgmuEPP0VXFbH27ugowBr4tUDaWx98TRJoiobZubeU5b1U8PGb3juu47U8UXH
UWEeGmmkHrAe/NLJmb1xf5OODcsOxh3O0vUrw4MCdbD3q9IPPLCC7h5ZMYVrgYw7
p6Pj64e9jn8TSJDwgOtOJKuy1way/UCD7WysM7iegvgsqdCO1z4Rcnh8ef75LEQo
rWurPxMf5Hms7P2x5euhQi+FbY+ts6KW60QXvoKEV4ZAEKV/j1CCgz/pjMbqB8+D
yIGo1nuVr1atI5Ed0KV3zgbyiFqQOxYxxO/gtm286Tdn6oKqqZiRel2AGo7fiQD+
nLQq5iNhnQjVW4J1pDJbiX5ffBmysDWd9baOdkoBJmVapUUFHuGvu/Sbodu0bQev
CHGOqmM+oigxSkSldeuZa7MZQTcCOeUz5wX/dvKMCLRA9JYmLDW9DA5mHZqMWA10
v6ClYIwbT0uPMu9zRvY+6KK88QICh+IrS5f3UwFlj9lscRvL9rP3b7b3FIsTgxpv
S+yQLep44P2sxN/7FBCVlv6h5ZBgmYqU/Wrx+q66/FxjDJkup5Fhd+S+LpeUmxY9
ylVi6Ps4Y34K3YdDJPi7wdJ+/hzbf2ZSZnOftnObgRDq77iuPStpPbnziSUgtf86
5tvPPnxFYbFN7lqle9IKToAPZnHXAiRG1m7XKDnJVInO6Bud/DvLeDeoS1CnP4rU
ftVDhxa4asReMQqx6+kHh1qhcp2OCNlCI/SgAgC8ulV6kRam5Bam3BgER0avRo9Q
44qAI+gOT0YaqKgRpGcn3p7dG8SPsYJwYaftKoA75FmOVmZER6n301TNXbPamHoa
cDu5rHPwQRK6Hflr1qs5G8WKxf+l0AIfRYbBuEyFm6UW67l0gS3YXGLrgCxEy5w0
JxWiWPFAetxlW8bZMCmdGdPgxLLDqRlrf6n6lspeNoOnA0FEnnTkWGn+MHXfYWMp
GdTKSe4/uCnQlAocUkGaL1p1OFD91UUfvpn+/anzeTPWRYvhKpi+fFf6BxzyEBVb
xZwzn5jzEzixjlWMr+QKdTVzwCexaxPyGY6HQ5lNJiaseblPzauK8l5BqoezfbkA
xePnlRLwu6r9XKvV4647gwhGtYxm2ERrulAsJjmeREn+mU2wrqYMA3EVQjGFqWo+
osGYXjntA5TtaXk4hIhtOeORaXSvKkRaNMkpElwrepXUhccOzitWNzjiJB/W2R9I
urz4EjkZYuhx7Os5j25EiCWqP0DiyC1KKVeqNG7bt3W/0g4aUvq+OlEeouuIKwfv
lWnsrRwj29oaTb1uqmSdD3b2YL1uRXJg9lPaI7LFErziCMld1UvwWRmkIPUxLMbK
/z6iOdod94L8xtM5XcPiVZ91sU/Z9MLGsDE/0wiV2sijBR9wpmRkj+bC8E6Q59Kf
SdWjHuNms5QxfYC/5TfL5u2whawpw67+v1Awi+QwTQhKlShiDxYy4/R9NxnCde6t
AP9r/dq913oAdoNbSgOu2SMHAzqCaXwBTaNiMbiaLHIXSHecfDas+3Xhegz2SNAg
5sMTNkuxNHtt4PtyDappdWi4ZZrtr66BmhNG2jhucojfqUPOUBhKIuM1lB111eYH
LTKzCsF2EA/yBtm4v0vgjQ5ryO82GUIhPaA6e5ML8/R94C7MEIYZmVxKsybrcIBF
5eBoWhv+tgF54mqilv09GTWxZvqygIFGTCtTPInVbqhipDWrPIaE6FLSKqhrA1yy
Y3+m2g93UD12pNA+tpDNhTXanKiB4zrxHokA7l+bxPpY4KA6FdtdX7yyezuzb9fn
PUt22KvGuf3s75Op78D8O2UuK+EOqP4lHE/NlCvaGYF48YihXKYyA/T+0OHShNnf
IGB34tkJOyblMBrQxEftPED5ip0JxQHDF5e1Cd8x5gkTRycsNbObok3yjWqBE1oG
ukPF+1I1CJoIe879D2ARuUamAzhJNLgmqrqgfV+2XC+CqNzCkKTSe/E5xO8bapw2
2laDKye0cWoFbRxgDIMnGzIMAN4E1lm6B4tDYguK8PJ0AHxfG7O7hgfBfRXx+khu
YiSIvcTogVp3zP+dM8fEpThukkytRgGXVJH9BXIm3FRGXCeVqT3xaiALVd/DAD0g
funcZQ/xRA/ilKam+MuaDgOHTMV3Tr9nI4wkYEOx2pIDP7gVKM4gV1vezo67IIq1
7wa8CWzuwAXMGdu2ojVK0zo6bm2Rmquwzo3/J/zfp/02D0QSot84RT1THJrY0OYV
Qwi81y/07ED8IQf4YzlMTQ1uUWjCWGlhaO2CvvxbT/UlvybC4FMeMWqIG2R1jbCj
hQfNhHN4qMWCknvugV5kuvqXKVoWs2POiH2hIvFHqjBOhNN4bi7q5f9b/BVKGpgc
SqM18BBp6esVO6BCR08FRiBE/5uTdnlKR9wJeUlh0runqB82XuVbJQ93GEmOkskB
moBOCO1botGW/m7r/+pSGkHwuPqCVoDbArY6d7WwXnhQuBbjPKpWIC4p4yR6sW7g
xgsZ4Hb4HME9iFMP3nI5ydpgjsadpr9Ht75nH8ysXFzIDD9MpyIdVct2wduXG/cM
N4yweomz52PbIc6udOAu5XJXq0H8KlJKAt4FV+Dv7aj6sFP3yjD4lLjs8wZ/a2XE
icBzVULE1C/CdO8e3OdX+nTmiZ5jYE+0z+fByNQFa2yelUa/ajlC7zWMf6WA4ApY
347sW7vd5BYnZdRPG8J3ccBIooYbrbSAbHlFnI2tmNmH8NjgpkY5rYFnb5PbK0lp
ka5EljUywoZ0dRN4DWP4PD955VA2PWaB+HN8PvTs1do1CL93wetTr4JcLfO3G73i
xMl9K2BdJC5rc83bkiOIOMWXEW9U57MCPQ4RNsQUxndBo1aQE+EmfmulerAztxaM
g0zRyWnQZF8evUIvDzhdBUGrW+OdpHx6jhdqkbQbD1CPluQ0qUzXbQt4wnNzpJdm
KqltMhy4oJBaevKuIRbSumR9L0QMhAGgB54vO6GumU9aVwW7yiP7QhAigPNz7MOU
ERX7CIDYBgmddcpOXiRlZvi/nKa/8+TcVqP2ROC3LVpwAT5Wrt3P0Mi3PqiCjjeZ
07KMNo0RxxrsNVx1wteLvFsxMuafKXYhLPA+2CxrTmjQVzgN/QkcxYYgVCHVsjO4
IZ3nbraNQj1vQH1gG5TrUOYC97CTzlDIZn2nMwebil5wIFyUQQUISt4fDztNYsdj
hmcvg532ZgznCATipeJxxxcFj0L+gf8TCmocZITSCcpXAbUeFVhh+5SOa83fN4Sg
WSHRA4tkkCKpYHCizD8ZFRmgiNXrCp+NdkuaA6EfsOBd9F6+uDHU7Y2NbFykerB7
+ZCSu5NfEkpfEMQnrvvC+mZ3t0NLXxJk64OmrQIhHX+KlW31TRJ2cGL/5g+kvOe7
6mTL6bmvsHUMVt9H4uF4lw29inu9kQwofJk9d3mLtgm6T8A6y8mAcjp1JDqf3bXz
3U5Fl4cOva77Ao5CsIc+6HnpvCTcLDPKQxtvCzjkC6qbB5up72kOb3UvwwTlCslk
hswLBtmpKWAG5Adw0uvY60WW3dvA06wxR/NxgS9J5BO3Hk4qab3NSHSLUdnF4k8B
2sj0kN4Bbk2yrPCtgkkEcSC1B+WVBr4kj/eBWI2iY7Wz5CS49+mnH+ChEbLBNz2o
OrjszqSBuX/ZkqvuZFxQaZ73QcpRyUXo32Zb0PQ2rQ9D8qVjGBo7dPftgM3zExaj
XheYGHWr3J2x/as/jOAG8e1C7ucCKIzsfzhnKoPCdghTY7Yqd977fJyM9M7RyI1t
IJJBiZaaQ2fjqHJlvHE6O683aHGweFVeY00xjBozG7TrOWTzwR27Qba2uBI7ygjg
M5LXrRAMQiOdli0YoPOYbjqlR523tpTQ7jFptHf+sZU2KeFAKMGrKYLF1yLyiDpm
zp0KTnLyutyM5cG5KhJymS+GKu280klXs7cl5i9c0jonL4PJptUjtKRxRqJPWHal
U9yag8otD5JATg7AYaYfCKNoMpg4GArSR0yv1CuHBM7TfL9GOyTHDUx8PHfZYY61
k4IsIL24YhNBpm6mTFQKWe6sA8hW4wyOeP+5458TxxZWeBNKxEdzYpc67/j22m2f
ZP9qs7+xl2yhW80n6c2PH1QB7cT8noI/mvFJhNTTNPSIK0OxdLW1xKfEETKFpJtl
unEj4MAAYrFhTAJhVpwBO2wbSjB2ogl4IDaxvIIV7crHU4oSWCDw+C9mhLB/Y9Se
vPs1SwkpEOFfRawyGbQIKjgCbx0+fHKOur8z7AB5Us/CTTIIlpDSrMxjtLDV5Zu4
ctBpxRe6JRD+lvG0l8y/mzRPZUicck9fx3zkmPsLw2gbd6jycHA5KFInrdkhlIra
E1X4H2E/yIRLEosq5vfOMOnkydQ0rcG7VFUZKW5Qly9tNcdTc56egvGYDtPumYp4
jcR2X99CYC2qw7LnpO283Ak9uTmB6ayKiRQebw2mWElsjXiZH6qqpYXQvR/Cb++p
tPB1Mfymkie3EqpF9U9Q7Scq2QkNMcVPIy4G7JGg7Ua3gQJSxzXk6N+GJMntt1/z
mMcHdBAMMYG1LS/r1r7IxzY1Hsfs31FQOSD4v1i84qnyPNEbmUJtwQ0CWY9aL340
5kVSMJxF3we5wWxQM3ekAc1mtwKLuskvet0cMTchntwspSFJ0okmi3d5/T6NF7FE
L6YQRfhm6hF7lm4kO5mejRIIUastSoTaBEynd5fFRMk6V45KXi5ZSAPhx708vPbO
iTpF7vJ23NDS84cy16wuANmZA60edRbLJM+IiI2eYoyPXSCSzhnASjWiE7L1uMQn
RajUkX82iJXO+vwGusQdBSva5I/S/g4cYVubJQKWM1vbvB3jhj7yODapzfprdN4+
mOxW66a11GW6t4G6H1YU7+RhJrohv9v9HChHMD/WqJkcRt/HvBTlV53e4JVkTniG
jfQjwAk2YemfubqnV1lU9KHV7VzkBcAhKbc+ckiof14Et9BuzX8GXIP+TdQ1r+r6
LzAd+Mj6/qNyGi6FVOnAweHoY1vOvYAuFjtmbwg20OIF4YqvHWYx4c6EeJ73PlAB
o4M6HhYrbw8g0+nyrxpazsOYmvneCHCvc+hlb/ndPBotjUaRMK3ibNsiraZogOEA
M0tLgJM+ZkhT5M4ZJf+RWp1pVqW8jq9OKfXZcZzZ3tvpTN9U7quAASiCW87jNUlh
hms4LzDu8pp6/OjvZW+In/DIBt6l8NB2VGzUnlghNOcqpF9ZruHWMJ+jJWhgayNP
j7vBsjhKR5Q2g+F7bSHVaZzfdSlbmNBmHWCUiDHiloCxCDzW1yYs9lcDq4clcokR
gTB23RBZb3qB6WMAWfrF4Sd+4miymeWz0yWJEjmfOKbHlXs9I6SJRW+Rrh3VuIBj
9PDEu7O5GctsYKUJ2aI8EzosouoFgpYfMNvWMPFNiWsoQa6H+6LL4vzhJ/nxgOlR
TIn42//Ae9/RdZmB4JzMBqG2ytMrlBioCbfxWPdEzZKpcAvkmOQy+FQsuVBAHkFw
mwlaZaKRa555xAx9XXFf3s5vfYydhsm/q9pSKHeogzYBqp2AKXugbhX6E7ywJbeV
AoGT5JReOt6QuQyQ3UHsdgNyO6dET+fZ2b0D1PpCfbhZGbET26xAjBfPr/k5FEHD
pnAoG35yReIDuyyA9gtTXEMbsuZ5vcaCiUhVWbyPWZDFkLTRQM6pGLt3eJhuIUAc
eTtF6QlHtufe5S18jFINDVe/lfpEsuQyCgdODVnYzuLrdnebl5T9MlxREZz92Flf
5LHWbzuIx/mC5vKU9KG/Y18HdwUT1GnwuDHmmV+MeNf1jcEp+pl2dKS4IJ8XwXYZ
A7QAPArsoWgiaLYpcYUMFPG7xy6ErvuLZHYDM72L57ZEaB136n68kR0KnK5d1wtX
FRF5axR29KhOZ3bYZmCPZ8YK2GNfJMoLyYKxYnpfkLHUetr8zj1eS8Oer4kR37AV
Tk4i65dyusXkKIxjEahWydsg6cGSSJkI8n/2ZwEfrRiKw94xY0Hejggz0xXU1Z9T
OmYjNYzV1IKGPZ7X1cfV/XUJWhtqLwmTmcSnGYXfNyQ5I/W98zy/ULUzHBQKL8gS
Dy91TsXb0mBspGajcK+rjCs/o4j9c/ivwFN/xattBs9Q28kWDwB53RMc+N/Eah8l
l4mpdg/imNdAZoKRtmoO+UkEYgI1XiyeTBNaSdR5M2iUj/4BReBJOs6vH7P3r1ev
oerqXv0xM1GPOsna151U5JpA7BbzhhUUsHZijzj7fda/xpsGbd3Rcn4TE/H9YZhH
ifP8CPbdXLs1U0lKiFTXp1rWelVdIxx5AcE0HYnwheLpDIAxXBSnW4DWaw9Z2YCP
h4Tio/QYlD3vDtL6YfyASPOxvt3RFXFd++kCPoqtBTMv5QiwrUGUpCjkV/Yum7IH
OL0EpX8/05S6OyiNIGOP9KhU8qqJfgBDx+ypoLpzmKZ8N9X2cOBoHbDITYXzoxPR
hSTEVd35+bCHkFe3DDsaXbJj79gYvDYpVMUaiYyZmSeQjJ7C4dO2wG9adyP8J4iJ
/IKin7jtEpXBHmQS9FWuo1GTYgAasnU8ooU6hzszQM3yKO5yDYwqPAz92PuS9MHj
0ZpyPe7g4FVoJix+M+oWPwWyQHz1dv9FypPo32gtCenuw/Gz+8xjvPe5myAghhNz
IAS3x1r3EeiWsgo1+CJpXYkXvRfnM1dGjt07oMSqi0XILJ8YzDqo2YRznSeABLVr
jEQNA2+3jWOnLUt8cJg9v1i2VOI70tl5R76JiYZ0yHRp3sFtShHz3wepw4mvSZ4w
2gOyoXzieEXnVpj+wvI8OHcS8EElPWAHshNt0foRc31uNoopm5+t8MkAuLlBl0DF
r0ys3hj6eXfw+uRSAxNegdCS6JfqOe+O/44mu0d4FMPkowYQnnmyndzFBtCRIUJ4
FgOH94ftfjAQd/a4t77kliAGY9WB2UcilkO/EpUyWi+j/7EEApbRSjbMZ3A1Vxq8
EGf20TWL5lfcsKdl4eHsI8sIBXuK8+V/BK3MX235/0KbEIvC6xzbaXRtwq6VlSXt
fmjgPy7qobR+Xt9e/cR2MApktYEItZacpcWsQ5nB+hTXKTswRgGWCKJJr9HQCKbr
5MsJqB4ff9ugFDejGu0cG34cvJKOUovkkG0IMgWrc+vxuj4wt1oXFXGc00J7MdbB
mSz91Zzce8CFF3QjqqbIdW3vYKGHJFdSqzE0jk3ZMpMi211Tij8gxhn52DyDTRRn
NRnGmYk4w5GdpJaET0rldDunC73kOpHlv/5lOfHRjJhdmMQp7brShZ/9bPcdIblM
7oQcdmDS/nvZ1XIWubhWL6+tGbBxEL5GK/WlhIDFV75th9oleo6IApbFx5yYABOH
z2sv7Kt89poHeL9Ny8XgBl6Es996+6e84Spik2EIfGb1lt0FB22VSdnKWnLEIQCd
ft+DEiTq3Q5+HA/xa3uHtVZydQe6okDi6uzrlUmNyfhxM2D3D/+V6NaQ2AakCmA7
rHWSUB9IULrMgzb1AM+SdEk6UW6k2MGXhVMcIGtvA7KZZkh2LgDGRYYGGSAgkSgy
WrRoOXTQ18/R0Kyq0b2gJzdbR+VzBGm7AF6BrMvRTvVdrmpVD3ea9uobvSZtHTT7
XmQwCsvQcl1LNYraRj3FbIfooo0MCUUJD3BTeQieYNO1IYEZdpniSmmA3T+Fw6M5
ScUSPX9AlXmiWb2Ka6r8ovwwizfkN5nHGTzL9rz73YbqlsqTXvAIH6gCNJPqI8CH
Y6AVbDJiUfZ+3I38NnS/+d9fZGKIwqcS5TjOys6/nBKNf9G+u7PbsDfMTUjSA26G
ZXNO6h1sZSRY3uy0e3/HmDUwtmi54+zMbBf8pWZgYJ1Bcyn1+n/B7HGYNYDAOeH5
Ai1BlLcIVL17N4n5UjYZJmze9VoQhASfeAfauuVHd9PNioG63LRnPH1H1KxXfJaT
zmJIOAuoWOuruj1zZRuohUZdDk1PLVsAcq6zBtNiKON0zfdp7CAU4po3nwYBgmHE
Gei4GRmsQhQdwmU2tOhcInSigmDSHGvO29MrDM0BkB1A/JbVoa1O7CgGCcX3I6h7
T6PO3pfiS5haaKT7dyOo4pC8YD7eP0DEdlZY4u8MmO2i4gVQQeEmTs3K02OAPsCe
imsahiFNvVKrs/TQKjKoRgpJheaEWnq9kx6bgPfCocuWuc/RgfxaF30LDv/VMEfY
iciytZpLXDXJlmCiIUj9rZ5Jn8aFeb7tOHEidblpm+oSw2uzB/lrfMsnWK2J7DL0
MEvTQsqUH3BAR5HwLqupfgXEEnu9u+coacGsLyvNFp3I8JmaeroQTAeR7s/NB0yV
rge7EFprRj8jByHRon8jPQsNidcEfQstnagc/okHQOVF+wR2DPPk07e99ulJ/ToK
p6nZav6/YeiNbNaxje2VoDqYxeWCW7yrRIM8cdeztWRvW03JmaZaBO0Qf9fNGbQv
CJiJdJAAkcUNAPth0W0agcV0v7Vw9SBnuuzNdd7PWed46+wJmPtObRN4DbkVaw8M
Ts+WPUY8mVdxwtEkiMUNqp+JZZAZ36jnrFll0/SudAAYHmzp//Rf8z9Og3UgHeqC
3s8VXl2F0xZsBSL+FKntcwVqJGx1XqdaDLzUtL2/pne5n+xDKCMZ0wrzP/HApAtw
0yPt92pgc5GurU1kTlfsqx61EtDxwunKoWN5aOSdAVaHtlQg3C8uZA2Bo2dphfqa
Ldm8N3uJQke/FmMtzxmqozT/h8EeQx6R+N234uuqFqlGHFQ3+ro/W+667erSFm1M
ZM6+fJAtUWjxBC8iI8DiV5d4L/q6CYPZjqGrcNbwEninSYAu9Q+XbTDoQfMbmdUs
xhIxjOs9I/0GW7CLEegZ8GZIdU0mT4weL1BRe0uADXCDA3CJdZLvrMGWBrZloNby
FOxD9IggBfxLqlkSNWas+x3brRvM9/EucUMWbq5LKQ5VJXJw8KMbYNdUyG4g7TXF
8TN9VgfMR7qu+OMMDnUI/sjhOYYMLs9GvZfNkILuFM5NLW+C4FQKwCg9yrihFh4P
VOS76ENA0PGEHiWrgmejLRPZmOVKIUFserTXwGNRSi3nHF/Dk0FAKIAgnlED6eO0
ihj0qSZyFEUhDPdqPIg0Re9FP3EiEtKlXCT7y3vdjRtdl404TQl7fWMB0LBegiD8
gQ4Fn20fLfSiHBB6Z3NnWsQb22WQr/WXRVgyzo6ZGfnOGTBpHKgeENRQYimZT3Be
fYho5da09SCxA/CANe8SSbcvcAqvxaCbtb2LoY9h3chi3fbp8QrxrjVPO60qr3SG
vBkEmkLyu9sdxttKC/Dzcw5Aup1Hlb8ciY7ypMh8A1f3mUO/850pCxLQZAtkfa53
p1fXKvGHUuALfFmLyDpep4VMK/wul9lfhbYboXTI9llKiEWvBQm2he9O+0YIWSua
tnyhLUyxRo2H+qKtP471WwX2fKcwHp8bBya/lkf6Ba+T7mLu5pFuNFc2/vc47nNK
NibM86dK2Qq5feCiWrReuj8cAiYifbFvw8Rgjc9vDyMBKBjnIq3tqISpnxgAKpOR
GgbjLjqBEVdZ2LZ4cUfxnaheYCoab58GVmFBE/GnvwMSDq9229Jioc0UiuO8O2p6
Y0aiMmeOhG8AGtEfGlLlFB79poNyH10Tuv/ODkQqQmoQnoQ7SgRjmPUgrbfbVB8q
tPDDbRAoDWijY3oG578MF5oN5I6iAhUupISzD+H7eSUYHF3rRFTNN2QUFxxc9a5j
RaI57mK9eY5l/Snv217AoAeK+OO/c1KNxWoRM/8OL+ypz+untu+pKRsycjzzkcTX
u5CHW1nEoxmD5YhwAAl8Uld4qTA+J5FH189NWhsTGHNaakXmtu7DR6YhGUnOKxW7
eiBVyTeIP2InqcJPQjcDKMRCJvdoekuf8P8oLnqF6qadb6IJa9S6VQNAN3ZibAJ2
96ukSY+bTFJBFCsgUgE2S+fAFbyeY1O+JcUsnI4/lSmAVnQZGnTQMhJHS6W8y04A
F3LBh5B0TDsNaXVzP4XvxD6yXaDCp/Y5tr2OwuuJ7YTtjuctu1WF3/9ptTTVXaIL
YmmVdv6wdwCTkXyKbb0myf2FeDJK8TmaDNwmyvif/v5f0NUsXVdHU/lAN8TkJxTG
Lo5PqBetc7UilWjjMTLAX9FluSAAFnE9kUVHRsiJj150oGfF9gL5KaAzsPXp/9UW
KT9vdO3VLLeJQ9buD3s/LMyJ/0Vh8j15Bmw9nmu16zVTMr9lNzUszvisIGyxRqaQ
kD7+E6nOHtpItV8u/r3wdmehFkhHXbz4szD2g+RYvfyw35n7J3byTQMkIECZNIt/
LPuXu2J1fpEiJ0Kc88BGtgxVvq7q7mtN8lwNtB+gvuHjWw98qAVg7FMNYbvsZolG
4K+nxFnOwpZeMcYlU4L1orDzA87B2TxAqhVBiQbp37sFfMKkBXFaYw7IiHVFT/h/
O0iPdRTLXblWuVfMWvRSw5ADQyL00X4fFT6RaIdgpdC1W/+XDB1kf3tDxWsyRCjl
sJjGS5HCf+Wm09McTKK91j66h/Il8hHwhmCIs6eTX/j1Il8hxRnK+9lxktwWGSLq
PrJoNPNH+evadIeQWRIJDoS5bZwfs4KauzNRbrfyCuC/xINMvD5jgs5rYxD6VILH
Qc3QSOg2/7ldvTX200H8K0kkhNhjv5oGld5KNbn3yhbb5E5apMZbJYbVxnenzcjY
k8OHPG68s/OEszkIxdkVmXoV/BSXI3Mm93kpc+j7t/vqcPXNCEJeUwiJUfBhRwnr
VxG/aYt05ZWzVgwfLIop+2aR73WKBZRY3MfL63hxeIn6fVDI7x+4Mc+13ZeNreCi
/RE8Esx6gNC0b1jGGfWCILt3LVkuzT3aSUkbeJSUbebrQSPclEXXzaH6Cwgb4oZo
0AwVFzsZQQEbjkbvBcQMZYnA1QfRFB8Wd/Ze5uezf4uXWNTgSARxO3pV0XNZdjFZ
ltjZe+WVyHOmyi7DdzOSRImf6h0vCjfHcpjVXpPsUAO6VYxGip79/2qqCed+UT3s
fSOyey5g6id9RGwFp3+OKnp7KXVqbmIFvtSW/JScLrmBvBXLw491sp4hEDNNlPzN
z9ztIipGsmf5ZAX57XvfccLw6Qo4ILC4hDTansUFlgJdFfsHjH9AlonKvjCpFJaG
uJZhXopbH4sDrRpU8Xc+ABFNW+Px4fUglti0oYAdMeophHzj117vQ0+D7vJlzh26
myDZKUAlF+VEeGvnMVzTrQT8jqBRaAjf7JTw9bOleJvxTGbZCUWZeo/v+c/xQHuP
5pHKOtS4/ZbEClQl1/RBlp6J85sVoeO/ocNiVA+kCtQnSls7ENv42R5Mxkbc/an+
bB6zrITjmj1SngujeUEhcZHG0KCXLvj6lZ42xZpsS8mzJLtMMzoOmvvqNWHvKQMY
grbX8bsrqPaZryPyo9BBFA04PBa0KpiIO3XwNzv3/yefj05wCFgY/JqTsIchBdcV
iMLaRUFg0gMdcd9qel2aLsxvgLenE+aTkIPQ3PxH7N4aAwrJbUfTammlh43MN3WL
kCIaFPhVuuQt2XZ/wPOYletcaL13LeiQA1aEX6qE8z0JaWHZaabAjQL2DkWdD/+9
NGYgvkwUlxOJ4LHt2q9yjPEAlPri3LO13bLkmP+Z0cASLV2bcrkot+TPj7c5MOJN
gh2buZlfEOiSyGJLFEGeg/fxd5EAtwiUFwzaDqyd+v1c+ydmiRbEfXvHXYxM9WOc
e9pRewBiJRyjQZ69X2WsPK1T/6hlEIfPI7JflG8EKd/rFpTtgIBEecjOrj2f5trH
QkTE8ulCOeDFuuxc8ddL5N9g1J387ZJtDZbEDsIRlnhUFUKZGNzdbF8FcyoA5IAx
F9kbXpzSK1BrWwTC7qbFqbK+0POLV6Dr8QvtlqgQGvDF4iZac7gnO02pRxOypxJ7
wNe4GzEguh/OdfbVxFeWZ+E5gN24RNi+rdwjHMkMITx6TvF4FVxR/EEU3d8uqjbG
97YarB5OJixEzdW/CVCyM7aPPRW4sHmZ/l0RpRufO/LqnjdJEdmMMhPLQGaqNgJN
Kr9f2ZZbIsUE+0fIOuC5GR+MWK7XzzOVN3ih7nLNddncLac9CM26BJiwCLmt+Te9
eW8Yc0NhvC/GEnIn4CFEb3tcwQHvsyfNQwE8bE/lB8yb/WGTcJF/W5lhR3mmG9cR
J/RnsKTuXE9yIOMJ4XgHneWOa2JsTYVxMrVcMPLbjVinqZjxrTbGwiAVp0rOE25t
PbaYVjVVxX9kLzGc3HdLCUjtKGCJLlqqQq/VmuseR/1gn0RZVflNNscymFt5ewzV
HIAeMnuJZgjBvK2FskmD9wc5I7XmdO7pKxDTBKgiI6ku1XVr/GHFBzQjdVMLovOb
67gKtrP1rIQd8nY5o1cnjHais2DrCnpVQXALoGOs7UQqxk+QNYUaV35nZa9aW052
zAVJwO1xdDeU4e9ZwU0R/3Uy4+gmlwg7H68eChin3nSqZ4bdBgP/9Xh7D8kppJDq
zbgQbJE45/mUb15YCIJUBHxgHy7bbQ8PVQKB2z6aVeBjDTy2HMr/s1FID1Xz+PIo
YOoX38uplw/HZVwVjm257mrMvrayzR//Pivz13/Bi81L6oCdhiErH6/s6bakEQjR
Qck9ZIRkAzWbwknNewf9Dx848NJ1V4ZMoty5vReq4zHyE+X+hL3LYEKC09yYGhW/
QLYZL91cmmOPuqjGL8VD+cA8hEcI7ZyKX+i/qla733IV/r3355DL1cznQthlXQGY
QhZ/9nKqmJnrXKXY/Yb1/ofHcWGkIJRBJwpRSpY+TQTFCg5OD53c/yPHhh3OxTqJ
AVKe4o1MGXWhpLBzdYs2kKIY86zwIU38t1yKaN0QRw6VNKSMj/zjZXOOb5DsY0SQ
MCPcElc4IStqzbEnX64616HDVDJIJswbwhhhiJLoiPUil4aAMcB0cWIqD6+cqGm8
QWrGQ6+ZpZh76K3tjYxdHM0A9xehCkI+cd4hVRVRIxZbqdEXhucuVQZ/U90TjawQ
CBlc85B4U8AUlpoZ5tMZcN0xCoK2DUDEgEiw1C49dvW6jns/8ubeyP60xAcFRkem
ibsQO7YzaK9Nyjcym/ryLnu2A8ZDMPjbFAM/iysPuqx/IXFMXll8XFDcGmBfyBGB
J8jQ7JbkZ1kYO8jZ2uZIz8OnMoTyyrG/OHbeTpOW8KrPtfCEUCkJL+J+Jk8F/iUl
vKXaygegZf1vLwyqCsskB/H0jzSuXzRKLTLhSiR/NIoHL+eee3hjIwAzesf7lzKT
Lww49d/nZGB9qS0kl/tZDqTq9QXrFh/UhJ9ouD9CsCTVeiym2RNoZBtX34jd+m8f
nIrNmFn937zvFr51sMkPnblNjnx+CpOGHP5Aa917M1y+kNBHlPCyiuD/94Ta+CWd
6qLU9g+EoWwNx5YUihs9xTPqgmHUQxGusL86EYUjImRyqh47sHAKql0qGCfZfbVe
xYHDc8ecogjEYuJmCcjuVAfdpLlinSr4JtDtvatnWaivUUpTrSmC+Ba6NGg2zSKD
V/+I9Sze5cC/q4YC5PE/yTO7J2821m0ZHG96uWNzDLW2KTybW0jS2s4vtzsEKavV
olm8skTlRd/8yKHoCAnDDKB5J+DhVfeF4aeM5c4+oVxBl9KPp23B07EYDuCDlIe8
O7HN1fAFMaGVVbMFQD7rU2+k8WWFPzvpXQYmhZPW8/WO2+AlysVX63CcaCiWyS2Y
ZeYC0t7PncwtM7rqe6meI3dD5F9LEj9/SDzgNE2PR7gF8qj5lQ6qpBMtsMLy45AQ
25ZvX/HHrZV3Pe/gpZSnAfBXIkSMzTj3vBJl6E6K/Mbr2VrV/ylO8+AhFB1y2J7e
zhjNPR8uyew+ESXYCsitUpAvo4u9BvXnUAisPH87RGKLv0sX/09JKkhN+U2ahkNn
+WN7msAWTQcui+1Z5NweqyoSSvG069ZEw3sXdpR4jYslN+BBLC/Uwrkp40BWQNZF
hvdzNO1Uo8bXcGBDiiqatHK9cKz4fQDTimQSkVlyxObqBymp1C2ZWeJesVeMjGiF
CTmGv7+fZBLKf/UvZCxdWTJ+kzLuNW40iB8vmNHYZhMV87KcqziWZSrgUIf8/8c/
dVT/3XCA0nTfGTFFVqLIa1VNfjZTh6efgXblnbm/8p+RwJAVaCfwYNDy+rwkax7y
TIXCt6+UL5/AM6x3sq4eyZyZpsrkHN646pSKXnn/vtsaD1CN1+YPyodfuOUKmQPn
mksjns1cEZLcwx8AHUAt4UGqUnaI08SWvgqvPBqI423zV2zTECIh9ncVI+ZBzHiI
NViP6o6x/e+stWowW0GKRYgcydNONwCUAt0Zbmt+l+g4j6Gu+c6Ri90Tq8wv8Yoo
fU5h86O9qPugmzFG/fO48GePMVzveUPYhtWYyD/ArHVCyYY+6BJx7qv/wKNZq4Rx
iVmAJqzgWS4VMKHX2oe3qlGnqmXG/kvd7gUAWPdB9gh+zkukItZKkrBD2mUzBz5a
w06zc2NZ9pVXmeh7slQ6xXqGobvqbezxtxOs2DFLLyfrxP2J+e05vlO9mWKSKIP6
UQjZy/vDw17+0cJ9MGZw+t2wzE5IKeVV1U+EqwVAtWKwBN+zc21CRHbfgGJSi2Ln
h4vcaEPOfZ5qvWELU6aZqTHdsU8Bt/7j5TUg+cJFn9NPWooC4pH7wG93T3fLX2od
wy+c4vyDDYC65tEwUPPIe5NFgNRGzLqkzakLBM2ojv0YQ8kU3fstBv4xKl8GUUpC
44jH2IU/8ICVzMrLcmfGL3N94NQNE35nRBxPsFF3e57uAzrrm/5HvFO6dbEisug+
uUGqb+ukj98R/AUtoiAp6W7Ld3iVc4+5tPQ/WMs1err7RCfIuvx4JUwoRx61MFRZ
/bwnesKdZzvU8b9hAxNm+W9wxq4o6fMRjjgrw8HBUkGw2zj9gqTWdnUKLKmW1dOX
P47lotJu+wbxI3NQqKB7Zyc7JvQO1DNEDNF9kHg1DLRxGH2tIDuC6PdeCDxDAWFI
og3/l+futYkXp7D+Fiw8EOoULwJrxmewnesANieRgQdNid/p62FS1VRNNbOV8T7F
yvLMeWTstQjgHktQQkXDCvI3qu+8YjGmyTIMypoADrcaM/LfDZfgvduV7pZMnJ0V
HLuh2CdBFhpzZ4Ef6wDd9yLbKI1tRsVGm8bMeD1/Ymqprm/LEPtNZWll2y40CCM2
hwwV1NgMohukeSMUlSP4nEMS/smOHmoelS2LTDUUNIEJoevQ/zGRdpcblpcEvEcx
ozPx5hyF6kLQFRp2scKaInPvzcMVUYwv51KtEtkz+Yjbp1Qcrf1h5FrbIlG2v0m0
pSjKOy9WAyZ3Jjg6AThqojDXAaKDu/t83kmveWNtRRs7+aandNmVaw1Jmj5ESNR3
ig9/lb+frjDSAGw88R9WR5Z4yyn0HfDvExrKZdGvJ533QNUDQQXXSOEjjXrQ06cK
c3yP88q6kuzeEyXsOOXy+0o5bhiNChQ7HK1Fb3Qy9FZu51dVjvv2Hv9Dyh4YYvor
ttQj+Rrvxl2tmq0vTdpW6tIos0qc18cKoxgBHidVfe+MTaAW04RNdb5QSMbXWUYh
NZqhxM0RZEJAmeHaps0rrkIcvJmqhPLZ/+ovnmxCKDAx5ELs3Gy3mJD5/xFd46b8
57wkC0y3yCU+yMdF49oOzxqeW2hnbl6heL/Vmlfecxw25yb5Fc8bOMiANxqA4maa
+M/2cpGnsJ8dqdck6s05XfAUJVVcRZRE0SccBUGlT5G5Q25vUO0lni0gBAd0LSKn
IiFGCazB5xMP7MBDCOd2o8A9m16py83sfvinttJXSjI75hfl4gEXj8v1B2jyX8fG
ni3wiX5FTuzm1E4kXJEnnmB5OSQysUbCRj5/D5ByFzcAFUkrh2a8DvbotaeCPIDr
Va5bdjWBsEn/2nqJhIHxpAy1SG2ohVXOLGCsvm0MFGPtVsvTYbEGPK4Aobu9xmlH
zTqUf9Z5zDpfUcytu3a7g2yuK0VY+Sc/hTkyj1K5h28II14EIfcmca85ayF+hjg0
FPrmnsgDTzFT/zNxpPr2ap9X2U3PY3tn7X+bYTDyy+GQT5XXlZzsroN0pWPBv+qU
j7Seu3H++G3xK2FBpVPQr5sKhmAjAS2DiwDvVu+P7CoYGXLEQp6LlgqpoWyfBr0a
bwL3rluI0H9vM//Cf3jIugPHcrGGdtv6tEE0RBQo3LkwuDzmOc+fOANkHiR0r37o
YKNkx6kiEOUPC1p3Sa3yYarvQ83FyJh3Ggi0Ut7mzP8doKTGChwXz0haNiQfma+i
IKDt8uyxWrcvRk+hhK9AhjRcQLhgECvU+Ta7FjtyOo33JtXe6REOjb4mXANFXu4T
amFm0Hg7wh9NMAOINgVTZI5zyGKwl5QAt5AQl7aeV+VAJiC/DFlVlqCSKS0AXlQP
PAj+yWL2gxAduHxnNt2gg2a1hOjrW75PNq62VfEYBbnJipweC0w8+v6/ZO0dDdjk
NFWGyObhfJ5eH25WnlA4je5X3eING5PZ5Mv5poMfYdZr8tOu0tetD5Yfht0rvjWi
Ic4WAMZSqEQ1sT1RDtHDRdo1q/vLWaQvCSu42WmTeXuc4JNHv00QiAD59aSwNscY
0e0I1bBEn5KC6CJDrTYxbWJablY5Vww/sEw1VYmRdmDsHv+VfRnpxzg1XJfxUiQo
foCm931xCLRWULR2fF8ER/jl4PxTIj3obK3cIjTmyPhB1ni+a/4gC4s74WOlM5Mp
Ch2ufuJt5X9lpKmxZK1fnJDxM3MjBcm6a9PRs6qITVCVz+3z1flhJ2JS7j6Z1rHF
AlXnS+tZArOtsdxG/RFxnJV+GFV14m3QfCWcIFHvDrkY7wqGcQb5M3UkO8/zAdP6
FPabj12LdW6D2yfyjWUi1l3c8AOn1XtZ/6yNB27SZTG9KQsguKcpyeJYtZpQ93+Q
Yi6Hym/1FCXPUt1yx0tL5dbeN0gAEURLhCK5wd2qYPTEMfovQCq0GL7FK7GfPGgM
YnvDWpI7RexlpOSnNecgKbTXYa2Xsy3i7QVthejE8kpf1BmazY2euB0teHhucO/j
eLOKNEu8Y9k28JV5+WNbgSJalvs4MZzFa1ZAUF0m8wokicvxTSDU7hvoA4JpZfr4
P7Rha2SbNuufiKfz6FB/oFFC31jWgseELdvaDAkD9LyYgRWs2PUwNCxDKodlC6hG
PaNEmQlxaMX0BvmHB8PtJMbSdBvqz0PRTuPVUv+dgx8I4yYSqU8np2lkouQ4nyL/
2pomobdgLcpHnbiK5AHM05j5+TEhRiu+n7yLsf0wy6oY1VOpnTa5xOzsWck7pJ5O
rXHj07+seUCxIihlsS1I6uP4b43/FMbm0ecyIF8Wc6xXa/UlhYpROQJdIgxF7odu
aXjCm1D5CwsFgCPnZq3bHpiJ8YJNhun94MsuleLbI5JIFN+NhoB7e3j8rCzCkh3b
d0Hy5H1rWfvOOyLf97aM0Ygem3A790ufx+MSHXzo2B9Hht4G+owpyCMzRajjd8yp
Iwd388TmygR5hf+TPJi4gtFpOp77s6pd8hT4XovMLiaAsdYDOkoGsRmvULsImbcD
DdGedWOQ2CcRkaXrqI0IKsoJ5xrSod/bBlfBcyusDRAqSCmyqplcvqbUGdaeizV6
WWedbyEY4zxcbmGUDRNeBZLkVLgs0hRXVN6iFyvbtkURZfIgLboisZffTv/v1pCR
5Xd6JwYd3s1NHP0oeTuQ2ahaJJbCNjtAp6B4Nf4nyIBbSUiPBW2U7r6Ng3+DKBQc
+r+66bbGO2XL0mmNx3HbUU7ZhqWXfQH27k1uJXgBRT/+ltsyfT3g1uut0l6HVO35
aDm2kEiMsQ3ZQlKtYA9lYrYbqujY5x+kFRAm3pQ6FQunOcwRYhdHxdOUgli3w9Q0
jfny8SdZS5u21gdEuH5CacUrMobP4IzJTl6/8mmZ4XyvpfzhCCjfwE/Bs+9/Aa8G
YHPIBmNdb9WWgzruhItxHHO1qeLpprloa99Ddp9JQ4itbwGVeEOBcWiT7c/9ZWXO
zmTT3x2URB9fKDdANWgAqAhARVNLRCLQ0H43Ma6L3i1nRZX3Dt238CseE44v/M3y
O0Ys1SDF6bj+TquwuYYl8Sw150zA43FUAWd2P8CXyWHbYf5OCLhM9/TNwFRW6o1n
DDPO/+Q2zjXU7Cu70MtTnjuqaOpaAuE3uMUTx/OH97MKBhaPkn7Q8BOu+qauJT1U
oAWwitCqtv46Uk9xXhkUUotpnQWNT999j129aJBjPbDQBlej4gG0QtmltSqzdPm9
zlQRw7hPNj4IfODXH1mF9k5WBGY36fFKExWmeQfLW/QrM2nv+ySaZUPYxFKWx9/D
rIa28BmVCD3OggPAwtu6IL+9WWp1qiqKIEfLYN/jbCQHdADD0I0JYfpQ4SsymeBi
g3psPhOeuf9joJpBF4Otmef6UYMIBq9ArIa2shGziw6an5B7kUeSdCsGhRMBS+wL
iWUNZf9HDF+mh0m2xQ8JKcrqdeSGf3D7eWOlA/Z0HVG3ZgiqtBQss8c9laZvCg76
cIFoGLqrclFBID4VX9PXelooEaOOQ/o/pUsAx8JR1lt3Dl6n06QHv8yL2Nix83rN
AVowKtTzqJOREvKkGKrXno2hO+5JUEEUufjqAgrhycO6bj2JRtZuLBR/ZS/q1xuc
E/Vkita8E8zy2+5i2ahdZYwJn3airrQawphJTGNoB5H30mZn4SxtTOMwmVKjpwG1
dnzkfbIlomcr+CoeRu+e2DEYsHYg5AQYtf3NUhKoVGWCAfrs3o/LoBQH7d7ZTZb6
mOE0TStPoROzA6Jz4p0KC6xcEJG4gEAbvaJ2wmMpxuCQH7depuaxQewKHrK3A8uj
ZGix2rNdzgx0Fwon36oYGYmoBZs5ehUhLcJwNPw48jwzufItXcemJnIbRl6Pda91
b1FkMwR8E4suybFRgoX8b8bZlqGTzhkTqUYS+4/kNxO7Aja70Ss/7b49kFL+/Mro
XNtGq1JdgKZVHAW0Gt5TwuDTc958WNq+qSMVWN0wNg5FUMcaRx1Yswjf0uOJAC9K
sDw7DV3FqtgoRptAF3qdINtBPbxiLSeSKzzArQXj50pFfGaZEn2Hs95/G1+MeCE4
41A7ZGxK+zRk9r7rK06ZFoKOZkSS4ml7xuVb0erZ9/anfO+VkYXFlnz93whEknz7
j2dQgQJw3j+xz0odfzHsNOSImihBWHhkisKhMtWmplOb/EhBUol5JFVDCdYowKqi
odySGe+wOkV0wzyZPMPe4Tpr2u0+KFq0SbvEzCZzrBG4I8hb/J+VX12zlvIrGb5p
j10bdeRL5tuJ0Y/0De1c3EJJ88dxnRInw+iqHvSdwUIQKmlVLZ+ss89cOvAOcJWQ
9i0mzHc7Og07Hxzt1ZJFf6ZTU3o6ak+GRjjaYf1rBtWrgOAbQOu1D2QS/kYRLhp8
kQNMpVrVuZGfkjbdRnmNHRSGnPkxytU06huy0FOCdYZOaf1TvIoLvqWzG+dmrqQV
7HzUdgBnmGZtemRE78smqCuAB2UxaneVFXld2CnGX33KYKp5Ff1xF+JRC3mhgLcW
WBndEeFXTR6FBno0XdtyR7YiGG6yEzoTmxE31PNMh7+nFmvkyR+BUmZd12eN6lbH
Xv+hpRyT/04GHUtjBxdgBMrnaF9Ej6TGf8DmgYJgkNmMlPvhhdrlfUy2nNlpVD8n
8xBhXHWRdpWpTsz4t8tQ14i1Dqg4JYgDuhCT6cmlmgAjCr4qx77khVr6Fqe00ddQ
dFdwFDbn9CU99rPvnMiRIdsTDfq6N6zWILoeMv3ZoTJls2tOFoX7JkCRUMQ9o/P9
Y7xu/uKS0pPpnSL8+bV7TvQXM9nw4cQRTR5Maf5207PRjG0RQGdr3FOegw+CACYo
3RHvK8eHxV5Z0rmah2BNZOz9SmvprpfMa92ZP6U8hz6z7xWLL6x0iJKOYZYaUe7U
Se8bTBb6uk21P9ES8+l42MC/F+McVdn6zHoPJq2G7nsDig7siUfFuUZ4zSIVn5Pu
aPfoaJVzKUa00ogb56D6EZAhQkDLS0aNvXIa7wOjUVwlDWrPZMSwCY5Zo8T8tuCZ
VYN5VdGWht7RwXnTK2zVp+1B071OILcRGleB59Hsn4PWYJ+L/R/zY1cMcZZsHL+V
A7jlBrI8m7iO1U4M3/QQ53mPY/dPvJULfpLh2yhRoYdtb+OzcYc9iMw+z09ocbBS
uE34SUGtJls/dXKI3oaayiiReCpzAdB+H0WKeHR1s8biCY2dyWxRNOlUhAPTUW42
m5R3EYkZGHYUwG224o5euC38U3IooDZxlQu3CtyycXcR8J79KciZ5VYTRtXZzlOq
/ISSdN3cNiHS1/oBp6hZLEEAi0XBe/7RPhHuMLbJzwNUgEh9lNX0nwDVKz79Q4kh
lW0VCWJ5rikY0to57a4BSeWDSnwT3SDbK+yPYs6wMkFAgoMRQ63jEpYr/ftV2XQ7
D1vqhmi6J23rl0VpidSxOax1roO7t3EjYcIS4zCm2ezWIufSWZ5Jv/G2hMAYj10f
2zmTBwpJ+FD/q5qk6djQUlGAGCeEbe5LAkrB5QLFGoEU/Wd/YLUZVPvnxP5g4cIf
hymUjc9cVLXr3H2PjvA39GuwB2Rh6MfEFpn1ISMcqUACdcc+keGiIlMR5O8mmMEp
zlxzH69UZSTnLjXFdkAKIvF1wD+L18PX8D0XRN3Kxw5l7wJuHyV7gNYFzJN7PD+U
aQ5aG6oLxXrAnGeEBD4BmyUPKs2cQyKifYqd8IAbdMOTj7GsZmFJnokyN0+6QPP5
yukNPaPLVJIS0MWO/LF1iQYgyTbjROdkYv5NjQcznCDefqIHrVGd8oqj4lV3RZdd
E5DwilVmIHzZy7msb3jqbe5avbfWG7TcMKVh+xdkTRM9ioaJlk0BjIAiLIzJ0Qv/
a/A6xN3Fe9KGIhF/o0oszqDNkxv5bJmReJX24w9ntZLxcgq7sXCS8WLJ0K3s0Oi8
b8IMbEI3CeWwICL7JG5+UiBq2daExz59ZED1gu4j4BpwFEqKQB3OEGKN1giYITT+
R+I2JD8IxokRiyapwmjj4KyJ196FTTAQ1OhAuZhszHRq3L37O9bA7JwKhHWecgZs
LRa1nGup7ZGlAH2N+D3nYe3zd91kQEY/KAjvA2pbMz+13uxy1g6N06sOOXr8x7Wr
oHZOcFE3P7YUkiNBSTxKgpd2ebYm/Oc+yXf77XI2AJcBMgZFTfqHIJHs7WNugj9a
g74j3av53u98geBIt5CsmyDtPssg7L+CriXYwcmq4HVhrNwSvYTmt5nuDnqbix/I
x2mw1LwpSD+rNXIwi9n+UKl0j6YOTelLnlo7CG49rkWhuQk1VUmHdgUdYA1M9GCV
wHNzy7RB+TMkFWSM+IU+kWFl9ltqgbqxAguTuQXY5ZSyjFgPUJneffqUSbpsv0s0
lk6I2ZDqEdHSzMbYVdGAYB5jEBb+KTIYTjMSeEgb86Wzg8E4AuiScHqdWZz2jZOo
qKqLjQtuRqzYU5MO7B+9YeGArsJm1WYMEQRDA1IsxcT0esdGpH5uzItSq6z5r4bP
UX+SMwdpZpyLa/j7YC5VtiUfNoi7d0dMzBgK4zO83eHGgwILlnVvL+5LIX7uhqDP
TQuoqj84Reifii3NnZz7O0kUl3OV5GtoDkeA3H184SOJ4cycWLL49aoZwia7wKq3
KITQRmir+ZLmO0jialgmB1x9zQSQOVVCUy/k4rAtC7ZLDzEH/gpby5rXatVnH2ci
f2CwdZHMjLyYrVIVgYjR+PewMbP+XZCjqArdOovWzt6GiDC/XAtm6RBvun6eKlHs
ntAzOsocIkCRsxw98A3tgoaWTX4qQbpsctAQFKprOjnKWlTAl2HBJFWxUQLSATr4
1In6uwRHWji5pHf2BNcOKr+gPrV0Ci74xmcHhgR+y9Mc/HBRXcF0EyQrrfRDJGnU
dmwB5Xyt5rNEW5M0LW7xwYDAr8tidJIQPnlD3YFlFW4UX+fQ7R82KnDeEWxR7RID
z4MmmVSmN8UACLZsH/lZyrppKt4UqH49zuQCvlgbaLWTfbYDLFLLZ9d6R0uRih0d
X0XV1r9hSjWF5fja4h6TNmkP56oYP653VJ+uaSDOVq7B1T5gYksUclKAqDJ/oD9d
bsRT9W5r8n16OxrEzpxF9tES0WC5UNaN6Ki2YVHgzQuZ35wH1R4rPvSmVJnMxMgH
x8NdtTflOqqx3MHyt5Voq1m5hX5atRrtZpWwGL9YQey6ksE5TWNsOPNcuhVTuJOB
EwMOuIzCF4kBv5CaLaeHA2HMRg1O7QzWWypbpeWdWCL6f8QhPwCQumM3kH4eDshi
ajfMdv0YfRcK/LTqeSBVABWOFhxCYmc7JgG3UNr6+rRWGHdECY48zdjGCbcXIRTJ
PX3pNb95voYqIBwSzzj+KAeYDnQ9opVUVwD2Ka0x3jsDAWvO8QajcKDatm3619U3
H3VcC71mxxZ1GRCPUdJIP/cZ2Nb3BC1h2yMvpHjpSRn+BAS5xwG7v7ireDdJCSCs
GtxzyLR+hrVAg+E1c/JL9SxjBesEwHfqnfieBpn9r1/jzgWhUYmnhcw/+4MREjtN
mgxaHiDEFdMzO1bKN+hDSHvyESWTSr7jRQeNGxzstrQKuuXEXS8Q4PgKtdqgCygU
6RIJ7R96E0IvqCw4x3nO5+eUCeyL9ArTKJL9UWG3QAbuYahYKGsf8CNLjFLv0c1K
gvHv73K4kdP6sYJhO6jbDdBoxheWphLubtQru94bqGfSKmmliW9DNgry+KWvemxh
EhQXoJfKLVBbJAV8UuOczH9IRBBIbI0LNGDFAHmNMZk8oiwL+01LgZ8B+z4j6tIn
BemFLJwac4HmzPzNMEtT5UWMo0NfoAHDwRD6FM5pgdqfk9gIxKVmIlL/LNavRqNI
ze642oRkGKgzqWJzmPK6/wynDqWDN7ft7enDapd1ZxNmlF3zwyPPApRzcm7LYIjJ
1WyZxE+3mo96/xbxIpPu+iTGpdmpK2jx7Ar5HnGheHv3Ab3PV+LlwCAUbN/Ad7/v
SueTwiFnFrmrY+uIdttMRrhtaaZFQNjWLzjGa3sqD7xB6RYmCQQiXEglXwVL5ij5
LvxbmT5qgULJZt0Y0I3G5aEKDlUjgZtdhL1KqOqrNbtUOvFRWGSOcrgMFmzY8RE0
v8L3gvctvyLbngmlm3I+plrOjdaspdfJAGEnmVh9bxbvWtDGlsG7KeaV5xSdIT/z
3Sx9xRPmvlpjVewJCMr6iL3z8Br7+bcNnaEHmdL2LK/F2l2xyZyJEF3br+mG7Zyn
JqKBQbhr/aLTaHV8BJurT8DNp0u0EcL5CHm4ZOReyH++wvWIOzVIJdoSlTrAdUXW
f+ItFX9VHo09cu5VF9VT5V0t2n04UfljfTmLG0M837Xa/+1qQ3yZobtRgqHRI+Fo
tneaOK7J8GVSAwARAZo6VNqNw6EE7qdads4EayB3fau1H7XBq379eEDpIlMi1Rez
ZsfP0L9bD4662E0WNlxZGGA6rhZuowwWQeLnJB/JCn+MUA5hSbnZV4BgjBxc7ieH
KvogSDv06gWuHE1PHqn8jnEz+6YeYmjyXuOAuRXs1BmtJdRQETVNhPR8UbxC8iCR
uFaf3WhzSuQT3XA2jzUO/KrWwuH4ES9ZyD704eHfWnK8n7m7tnyGk5qDJS+bNqTd
rTU//Z9sbHLyCB2yUTF91bXwmMSSxRLKcfXuOZ6ACEauHQelfPPJ9DkX3cEkcfpM
i1WzqmkM8B4u+AimI+qgUmKqEI8tvP2HswccqGpkqvXy5tYt6b22Jz7H2f8IY1mz
+Z1Kqaf02mpY4ziwoIi68c+Pan/gaSNPpk5jHxCgx/dATTuUn2EGIfxYsJ9PYgnu
TvxI1/Py9xVWJSDZ+QlqDFeZDgbn7oLWqPtvJALHArY1D3Zp7GWzm7zW0xMlu/9N
bzFxvkZ1smKRp5ij387dzPndspbudHEB0HhjK24pB1s+UWNl/EUmWLQBLpVBzhcf
IEDiwegDKw9RdRphcbRpaSz7QvmUQkzn1+9icxoFO3HlYeO6QTm4gLzznWmLjDU9
qKLMpgjrz0QG1JzZuStLXs6LZ3ffuLiUnZKULLkaC0zIrENKSftKiWUJJYklBUlc
C13sl+ZcJxeszY+8cbNPSe5M42lmsj+xcEpnSsoJGRb6CIjIKrXluTxDrU5r10Oh
+2nXBMpwdxw5wuzz9hnN89IxZnhB539X8IpPP+rq5/XvECoRz3OasRZUBGqHE+e+
HRsrtY3SDRHGSp31C9kZ5RJRGGywT3uMgC1GPOn2SkwSDuHvM+uM/ns3cNdjOFke
IcVwsjdhFWpIRCUUd8GrABhOPwsLdPOyLCTaZ+OiwcsYElAuduGYiFKnE+AvWbJT
YqS7meRh8769ZZgvrDWfDvjaleozcdclAEoFOIH8tf/Um14+SqMyjZ2lciWNjfGF
o0r74PpgRx+vS1kQA421iyqzRUCj3AWszsrb4bm/xKUwcN8pcDnV8GQ0eHcnyGbi
olfkCvnRQoL6c/JKscb83mdjR3dWhjrO3OOHfH9yPxr8s1QDrmYn8//sv2zMDt6K
GYgOlgCQj7nr7cljW8fzy1DzybnWtnFmxHrmXIbhnU3j4YPnb602dbx13+twfMmQ
/KLog5uRob/URDF+oPjlKlsurO0Z/HHgsQam8sE1r6+2ITaJtOuXHLNSKRKOQ5SR
ziyG7mdNkfr2GpK31B85ChD39CjbYuHz4OS7ZP2pYpu9bdj2eNOZ+8CJ9xUA09vx
wzDsonI5kvHqIbQTRDsj1oZCfqIn0bO03aWG0C1HdBSFRuA31h/T+8MqDb0xubpS
XyxIxNU7XK9rhZUaAIl1oZf3VSYj5zDx0oFZhDhvLcHA2DiCbaOkeOI0SKiuo45b
6eDa9QoeA+aBP/hEhJAHmBMLrZM0wznWzTO477hg1oYfre7cWxluDLFxgS9Y01w1
AC6lgz0q3bTTUpfwSmX22KQLmHv6M5dg1NT767Skhnmxpmmp2GrRTm9zl0Tu4/i0
w+TaEI+oklZm7s3dVf6XD8sWyrD8jhyR2dJhLRpDrTJENTWB6rIt0cNLZdSwRYhG
0kF0l7//2bSDX6iuw9yFX7ttSPqk+1lfVHkiupifq7/Pw33hkn51mzzZ4l+RZtYu
oMlT/dkwEc1V366Hoekvv8AeDnfa1cqf8dpIIO6/JIS2ftaYYURXpnckGD7Sxnsg
EafWNv/dWakfip/k1l+qYCtqxJBNhPwGPMpePApyEb2C6LP+bOhFz9ECVt6/9NUo
5tQM+PfDc6rJDLBL7aEeIE4M81UEyiY0z46nVfndCASANt5Hhy7DtEBQidpRsQoH
JqTlOM7OTtd/VvrcRi7z1nwzPatiNHlICV5czuJb4iLdJ2+qub0xcrXqb5cBXsqG
ytb30gC++OVuZCBsG8SgDo6D/5d/DDaYfabsKN6Y9TjmaRXVcKoBt1G0D8l+uqqd
tHyC3n75o08gvYNmgcY+hPkoIMG0cf2uYQC1AtLpqxkYVJtnZoLX4XualN52MLab
rJpvBCUUK6xZHahna9OlyhxFc6EqIAnSIrtQdOgMJa/b2s4qVbpXCGbYlQYUN5FS
nMEMdHWGDuvOw/AMBCinJkWLzFeLwzhYxvwC4OjRqTHmNgaMJpLqpkJxZ4P96q8G
lT5wyInF+HLETZ66kF6tVCzySB39XjpQAWMKfwkkFUpPbXpwhpFwnsFCHyJumi1k
88ckmyy2YAfC/vygT9yOLfYX4hHAK3Fwaw5EtJKGaQIqsQjqpQwyjcokX6sv3tWi
gJdIVLiD9pD9FVEwBkPlROcdvhXl1Buk6HV62oFDUoBYVovwm9Q8d6cg4qU9k77r
xMjLOMxcOGAEoYKwZLVwR7WZJGq1l8fglmS3zqSIia9mHpBiRSZRLGnjQNurVWH4
LT53ocie3g94HVgQf6FV71iKI27zUN0DwjQEAuSwlFT7OGh1qZCQdRhL5PnDx4MD
q6otY4qKa9nCSrvYUAJgxTnfno9BIF1HLUr8khBg4cx5Ch4IaJXl6hWohvaw6/LP
qycRTZbO0fovyJq+Wjliy/DVvEw4Vk2cSz1xNlHGJ/CtLm7y02NUIbWlBa6+tnA+
xXmhvVFOjNUKc/csBJNmEfgygekrW0U9lrEPtdwLpfFNN3pxIsD7672m0q2WmI3u
siC66RrU9WW8HRG+MMHoeSDNmdOrjPkYTEw6tHKc27BehlS0OKjkJYzrwa+2ks5A
0r3fUqIeEn016yt3ywRxdC/IX5f1mY1HgsI/JgMxkIM7ZApQBeBKjtMkTGD/ELxK
zowQb25kr6WoumhwLxefzbv7psUT2p+XP9KL/JWCEcYfy1ZKdnvOPQR7p10nZvzA
EsdRnkgbhYhrH0UjLMFEnp5TIW4ZjSt9V1ZyYs7FYnS/fZzD1d8JSq4sxfnMoaOj
+sTcLk1nHjYTG7W0hrPw7gOESYqyKtA49oI/K+NRZ+b0PN7JJ71GcuhDy2gkNfMV
y4lDhji+8U959LcfdZ4vfONjZHdbRgLaGWocW3fgSqRONrZJoLCGP8TQvS3MSoYl
nnaBafqA3s2Hn2Agnykx2BSROPlTo8x6LCncdBl5WOEwLTXEiLepecMjp1ZcccrA
UdhKBplCfs4Qayf1hmdgW6E1I9lMwjcY3AIWk2RdSkI5boRJlLxfMHaOlw95hNFZ
mhh5D110IHSgO9+lfS69+KzGZtJoVtdOoaGl+JvaLGV+tTUYZGjw8IQrKMymeNYo
lqeGltz1VrH+nNqvDfWoOcEHsXxUu/Z55x4TXdHoYZpOEpw+HLaHOpGMlD573Ue9
uyiJatxu5o6x2ftZcwXPJaNMOE7Jf8yxKHL1biN7B8qt/TASE4RaXqKx7yWtMbZY
7qRprhHzlNv0guvkdhPAvQokm1zlVH29I0DeFPEiC+3NftLfWwQ2lQathaEakcT2
vVfoFjvT2cWrSy3cOFyzO7tJGpbrLufc+mRBSHnmnzdDnRTcLsv/QibkxqM9HtCZ
8QwJOpSdMT8bjI5KgZUyLSGIMe8hI2n+uWmJNboMC55nh+prTCAeBSz66k3NYRTK
t6Iys3eJ4ylk/brvSEJ6TZmhM/PiJElJyR/cqsdkAJyMMbPpzBmpPNsYlhN+fq7u
YYyTpn+AtBW3sgdkCtUpabhgiLFWtCg5KaniORSUHsN+nafx3QrGF/2MkStaHaUX
7c503wlxz8vCcGIhe7qMhBVQkdUwaTcbQBO7zmox0T/Nql9l5tFIFswbszmgO7ac
9W1U7taw/h3OsDkDa+Ui2rkZGvHX5VXMdSUX4oKQHNjNr1w8LmmrjY7kOSeB0LSM
JOj6sr6RuaiH42+d3YCF7E95gM+6vyYew2AjQMsnnXJ6C/l9N3zntbhVNKjBDHcu
wbXsnFOYJY5jzuKnO7mogxOSzRvuX+tvACyIEFcRJum3uo2o4SGlzxDLbJDrcXoC
ToIYzanf2Ylefxh0tJnVkIL1OvL/Ylr0RAZIYEeuNSFfwJSj+I4QcHIlHcyzLhsj
4FnJNUzWe0AYnedLvRy7bENNSPO32ZbQ1rog6/BaWRE37xOEGxPZG3wyHeU48pmX
MzIGj2LYru7yu+03Kzd35ecAgaonY1uDW2+HaMdB/Ooa13SdbT8XyQoY1Z3Wh+TA
qoe0kUmWZjpxdsKfeqjoGI4p1pogtD5aQBbauOYtu7qnEzrZAoJSzZyHsBeCNTny
j+VxqvL0H09yJGsScrLbOrXRdXeMdbp07Ly4oKy8LgHvoAD7Ln01DdrModGPGjPE
cjzsg6dPuioC8zF+2cnFU+7sBDa8qZ/0Ov+v+ghKfuk2JJJxQFni9a2gNmnZtR5P
xMf1NhI+2l8Fmr6Vcgcq6sNTlVA3c8qp0spL6+uGXhLsdwhjqqrhYB4IKv3IrAw8
XyLUzmCYVXf88Cos80V8jimzH/PLbjt3x9UP7dQVQHll5vA/DrKqjecRNYDp/qbm
M19sAXviJuKStljAShHmxcJqtwtUCv/yp98O7VHZCGtM46ekn4BVjf6jWvSmti72
Dp3hk9SPeg1BswQ9IkJ1QwBHuZ3M36H3aMkF60DtslOa4rdscsRL+6VeADsZwUjG
9nRprsbpvhoreA0e7/dHSMJTkx+afyInqi7ZjajKoJWWkK8uFC74L3w1rEEwbDEC
oSXSfNCT2lgc33vpn6Yc3LL1h7rYUbFSj/Apxf8Rh4yP0m3GpUGQOSK8tWW6fsp6
A8MMs/wCrM6ddTI1pSpHjTXLoaktgc4eQgKobnVVm+AsRCVRI1TGwxgyiutzMxhr
IUB3KkV+TSPWVKqrVPhx2C5OiDYFIVUsnrBL++3skyVicx2CbDNxcJnH+cA8b6+E
avcaQey3otTxVJ12F0HRWMv0T68GTk+1EyCTTX3dRGMfN+VkE2Jssk8+BZAQR9Ny
njIDY6JguwNhAxmSSO9Kx770cdiVXIVlEAKs2rDr/btaHPUQZG8vQUMsHT+dRLd1
/PBRBYEHhcOeTAYFtZgZ4H6jSFQ4SGN8PWUlVREMgpnQNPZhbAnOqYju4ogyzf9X
3r3hDfFp4S9TyoVt9Br8QTa2pb+052uTt/asHavGrEOGLFWGEjn9qBKzGVZxTuXG
k1FDttkVxAJM44BFyqWed26S74677+Eumx/zOuJnyZf7BHmB4xMm833q4p/vk4ha
WdIXKMKNyTo+6AmU/yi+m3iF9DUF3jjzRyoKkZfar/+wjnxEUfQEvP5tPWlTSF0b
u+ocfzQ+XOW3yE2CNPuayVg8lGC/NeD2B+ayqWOT0RRwY6bfakfwWuLKf23T/n+g
6M7IPkAQ7p0WT4uiFyMM0eMLy55tcSsI9RggYA8L0nQl/yGnAWt08ET9ebSPHCLE
+iBaPvYKS/Ql7PHQ9zn4syg6Q575LzPWZPPE4+bMY+/4ML6NYnPRptN8BPw9Xxiw
E138fw95gapQWMUfVf82MBhtlRyeQGXAFF0VTzl7r00Shsb1NkeHlSUcu9FR9L/G
ttlYzLN0yr7XTotTeucLvLb3ogdMxbHSBuDxsB9H/hzAXeUFxRjwyFm3pYPerqZ3
A2nB/m71MsoRSeHyLgKIgEwSrRfACWw6ujxEhf9P6bl+9yFpOb1NBy6TKOE4bI4c
Nl3yhxKTTL25sd4PYdYITIZcSVmUfpMfwOE2/JPw52CKYcuKxhN89UmZp15cfPnv
05XeclCZwp3Nif/7DCdxKaH6kYRAULcDz5QMrwwj9RjXJWJ2w+r7xE9zwEMzic7N
KOZRGeu3ioaoWJXVl5lIGJ177KUcQ/Vczm1A1G0Iw/JbjI3S/oGHAj5j5M7bZ/Js
cysQ/zm2Md8M6T86Mri+apxJgka3e5Hwo1MyvnCD0iNQy/EwFOY1nbz7j0Dax1Ft
P3/aGNUBRUCwvgHg8U9CIA02H4Pm9oJQ4zQGXlD92knxIa4x/xnKwLiweKUgqecR
Xa8iG0EteP5XEp0ciIrN0YrmxTI3yRN8FWBnlSeUtRTKkJ695aEVXHD+pKvc4L/b
LxQTu7q4hKp5L+svhq72zNCmjgDHnq07xrUjCbdtB2KmaDIJMDKSpevd5DP/ZY25
gaRuxZs/ImeHSOe3Qm5bGdcHylxzh+z14Fv4Zuv6LvhobpBsrvRhwGKa+/zyaHW1
i4IIz3wofsh4FJKJyPK6mLkO2WgnCBMM54Y1uwwPNoZIL+Zy450s390cVOVoiy38
wGU/xirUyZWMtJuoZs8i1jGTMjgadZYwAb3MrqxfphpXQpEoyO2XJ3jmeVESSqcE
X8oyIS96wP3jVXRTW5WNB5Ye7BgY6c584Wr3FXcX5moWpy+SHhoX8loMY7xuewp5
owGqvYVyLv1RNra21A88kd+1VXnhXsM/InIt3d6mnyUgnj8Oy+63xqSaDjtGM8yq
mVxhMzcOQIJlKzCbRBULUsj1pypZ+D+1QfEEBVDAaBDsIM2o635zs95GFHs+heBO
DegwZZxKwYsA+Jn/YFPecok8oe/xNsfu/+to46odMX0FDD2l38NZ1GLnbMX44vF/
DKIuBs+SJkeYFukAWmlXTl/HqMIcTGrgHAbZO6lSPVvzWT+qmDvzj2S4oazkjugw
bRylvFwoOVbv32wk3Zxus7pzrXUaHapE4qfcNPHF6TjU7SYRsCwcTOvDJ8OVcAra
b4RkoqT/1uqejQHumqoY914kl1lzm3KH2TUsMaAsHC/5uqcyeZumJSsVCsQws7h4
HQrCjdgL28chont5XQSqHoIv5cgZCO1+BH6Z1dR/vdwtLypcJjvuNbvZECUDKFds
OjbWrePLTA+mQV+CjlL42zic7tvaZoHrXme7tUaMR6Wts6I31EOU1MryqNcuvbou
ZkyGBekEi6R362Xn+rSPlqNoFGUpXq4GhdAE8xaP9LCLHYn5Ukb0TwBXXncTLf/q
XWO+WekK3K+QTsb+l+ia/ka7l3bSOlPESQDLotCbcNkjuumP69oAgrYaCriT1wPI
UnCn5GttPoJPVIea9zvQwHuAD4GFk8LzXqbdqv3cx34//W31pjAgOD6W+tzRy+94
ws6T0Rqtw96Ha+PQpPvIAKMt43Kilweer1g5jKq1pRw9HaTgzLrPtgbFlA/rxU5x
DKXqqurtewykA6NLvsr9P0m0+0Z85wzUXQJ4Q4/mZOLRw94Oi8hPswbZZPxDMVMY
vRyiCc8pyub6PXBQenz5UWxlRV2L33urqOA7rP+UPl8uSfBGDqun0X89rH61Mga9
l36qYNTBlLoB+KIUOU7T/sMd5dyz2BTAyRXt3vDhIyWWqSbHCKyaoH/tCIdemLYr
9suVXYeLZ/IGxf0tzY/NFy7m5dp1L/D2/aCbkm2WuX2Q0SZvj5I43sMOGQW7iED9
lKR4C+l56iJmTAqw0EZJdpGGjHP9IkQvD8FE56wQ3frnte72To7C427SQkcZoFYT
q3f4PjAUX9t552m9RnpXnTwZHpT4ao5Y+XvyfR7Sw6kOEtkrQp6YWJpP8liDW3Bm
HLENGqU31wpmLOPZQY7pTqli0Mpg+rBgcHuPtLdRRs7lf3oQt/0dphP/gveDPiW2
qNorjUfZ/1kD9DCvQqfORKEbl3KQKz8wVjLOG98bP92Mcw7G3Y1fxSCOii6HBhzu
pchpY5Uxxgc8nXoG5krpBlRkE+oreYavxxuDaIIEJ1Kzfwz6D8WQCVaF6EGxU0F8
MTXFQ/qDHhkb8epl8U38cRCx6XqDKPJKvfMOix9CWUdtdNR2bXM7F1xc2vCZ/Juz
kt570OBe5AERxyOzF4SMn/Nlephzlso7Ds8cQ/xQO4iNbMAsV0Q1GMf3EkuC2qL8
pWFwtIBKRhxY9IZofWzjiSY/rJbEp61UOfdXRQEeB/VfOwEBwznLIs0UhtlbxE6m
/ubg3Kddz+ZTLZ8DLW0Cveb4Gy6f61HHMZZJEBvlQPmUzGoKZohUMfHmKtyUgvV9
eoGtBv9gAxOVxRAvXZ83D7YDpnKzeeXNX+aCJK9wDfIZZphJUzV5gGDPVJgxRObi
jKaGcn6SvpOgEr3e1dut6XWcdc/iibERUiK8kYAbmLVKYFvIVDUpnIYShBeqfkEV
SWUnixqpwB624fLRQX5fJK0vreKeXLyKfNUc7EYzwFHjrMdUbetok57ZRQuiDeE6
A/Vm5qDsB+iT9+p+N+gV+HSsmAbS3iXkTaJ8QWy9B1m8RzcbTCVfJYIuHpsxCuG4
yqRJPHWVW2/Hhk1hRP4qA00IKKocq2arG/WetXg7eAhIxAiTjWibe297rMgjwO67
1lOhC2msdY2yRqvVPsr0rUdLb7/kS8XTXJTOX4I142PaxacidlWdJhSiNwhBh+hj
siyHhKYGYH2nLn9kNMpaJcmWHk80UVzRTyKNy4fnmMUBqICJzx+d20ScBjFFcUwc
jN9UR08CO5EqxqBZGdi3z6ckHnrAJ0O0dJlucQey9IkngfpPJ2P5O/Tz5iq6LMjX
5OpM+aS9hQl1tgqlyKWuTgHxRWcEDku4t8cVNbt+45VQ3cnHaoTOH+BhBE3QoqD0
TQNe9Sq45/9Wlo+SdezLn2ZS1c5LpgbWhyYaFWkzDfi8a/P1cKyjYP78OqSt3gL8
kj5ny9OQZjd6ebGh2+nvj4LfbanCXq5ZqugszPmlvZkkYcUz9wBW7Im0kg7MFHMi
kL97Zhr8RW9Pun9Gq5NLmX1OyyuZQRfghumxsbb6C+OSAYXcWAEYmRPAh4SFhRCV
4exy6dHYtqlkjrPOCs+LvLKQKrrYNLJLc5j5Nm31pxySdKPhFWDLjkqxs/a+4m23
UbKCLp/73QzcyxHtJcyXzr+XRDQdSY7GK5MPl8jTJAfMbUsAn7lJQeph/VKmZA+t
XI34eqahA7+dryQ9XvGHUAsAQvjQ6wFvZm3J9fgLoXFGc5lhDIiWUgrvfKNNps9s
gv0OzwRVoLc9hOsqx1OZ27eMblX6d1cH+PI45kUy9VsZItHIxJJ5E3VXwPABTwHZ
xPYRTA4cbBf579W9qvQFniYjSJ4LvkfKmG+YaMKdjLhgg4/lRhchVKqCXaVWlN9+
1CbiFZPkMB/HCgAkxU+ah4ZkbXGi5U4mwTlkApdZdjzQ7Xul3+hK+0+nKaIyLPGA
l1hEpeuAKD5uwofjk8ujNH2OLfTJSPSjhc1WWNjy9+I5t1vY+kuPAA2jF9q6LHwM
aA16jMotWoQ42kntykDPpZ/Gq8b6iMAsmmuToqYdC4jf76fxHLSi2c6Rrk9JTinu
qdA5LOBt/K4x2GH/vqs9ARPe/quyk6mSYf8DqpQMhm70ugCMJG5GNPeprhq2u26n
MRe4qEqfabtCXasrKP4xljkCVd+KwwcxNvIMSqe2oefVFkBw1SC9HgtcclYv7BPh
u6F78FoKBhHtrWyMZMFiswk5vJGKT0vCTfbpfOkbnVNMozhpIFDiSvzSH/KtayyQ
BOQWMmAO2wYaI0FiAUCIwnopXSA6QC9AjYM0mmHSR8t36TcgJbduE4mvbM+xmgCy
tqWeqPy4R5annSTm2LDdhzuWsFYvtieBuEOCVtZRJ2G49Tjw1PsCyYVuGYbio81l
F4RCZE1xSD6JSn79N7NfTb/wZMg7UgDxhqChJDeL/QinINGROF7uzVj101uOdfLE
LDRRkYhckan2VI8APW1uGKueQL/F/qXs22YI3wWQ86C8yFtnSXihqFLs9jkWRi0G
Q8jO06uvt/qKvSvVzDUHJt18IMx4v+S2rtft9ZYG9Hjlp7hC+EUfH7PekY154qg7
e8FwcqhtSOB8jmSjGSEKBp/S7jfl5cl/PbKaRQhCjPdldL7/sTzJSHvJSRxkzoY3
TjgOYR7RBaBQO833pqiOfYNlYMFxXevRbgnCODaiiauGOhnU8AurloZGb7Mnm8T9
VmuaFnRy9KHUanbO3Vp3z6Pa4lSuYE6WC9C/d8CYGNGVKwOtieVzAmSohVj7drb0
U5o3/OnfRyb76QNQ/MGTyIq5AyoQ6LbNFSt7lobAJcp7kEXBhMWK4D8DiS858qZI
tR1b34ngTMxULNQRQOX84IB3UTPpLDh4G3voe9uShcgPrsXy5L36gr9P9jXiW6Wc
1jCIp8zrYvFUdrGH1nRNWV6AHx5KNQVZxo7etDanCLmiFEnbnIxvdTnr8ecb1+vz
ZaiSs+dUSAO5EQnge/2Y42qR6Ohd1WP/bUhfV5YSKU90W1t61v7WPYrVsPGA4NAj
TyABWUOzFqyhvtjlopIF+PmYEEo6ClgCY4dDpUzf/iC6cJT1XPjtuUBdL0a4o07Q
SHOPCl5BQ4tqrnDMB4cblSI38Pq9V4IEeXQuY0ZfHM/b9RJqzwBvAJug4iUriYrE
1HbgHEfqmHA1xlQNf+xhN3DOJWbP9otfwbTSs+UJCfUclopNtsUevKjithH7zdkV
mZwMGSTFJQLuqfwGAbpnVGOvYPpf5nA4t5O0Vy2ixcxaWwuKfSbH6Qq2ITJWmbNU
uKEdJqnO2nnJyVw4YDvJ0JljKAZFFdI9Qxdawts3tRbZdIlETvsgMK6XrAugpwZu
n2HFSovOxt9k0HiPrQ0JZoys0Rxkb1AwuktnPdJ7BdkSF5+8JjaPHK45hCJzSoDa
PLK0swIZqzOL8qIXQUsEhD1YPZRTuTZhCMsbY3MQIdR7vD/Xeu+DY9pQqwGsXXdx
PP5FtwCf7i68F8Es+hiGE2PFKkzv9WSpOmWecASyZUfWCYpCH9BZvh4ZGNDq5g0H
clIWA8F4U/GXQKExepexS2XRA+eDUwgFtI8DRlZhERcum99tVJA60sIrmPzPHG+w
BgVjJem9xPQ2q+0NC05QeAWOhmGrS/bezpQNQiK0anNXj75HC0eUGL1PXCmTA1mt
VBPS17Xm5oPFhOYPF2Np/Rub4KN8hbllixvCGhQBZ4mw+hJ3UURjZN+huZ4ylWPW
B0YUwN8kNz27NJn67IfH4YD8cYWM2OMkpFTTSeOz9bonU7csxRiXEzhzxBeQChRW
TK75g19k3EnbMbxlM68Vu5vNfBoU0w64W2I4HImrHV2l9EM88PJJOAh87NYoX+CA
4BQ3OBDPQncLBy7rSsxr8bCM0MAOkOg3yi57ZkK+jDb+YSzL7UsUlb0+rbZyDA/9
GLAx9sQvD/KHtgrYRNfrx6m4PWs/94/nZtFVohPIgesjKbYIeDkDfp5NrAsGdLNt
kwBiCZRUq1uoxRJLFt0lomAhpRiHaAtxOSCgqWS0aBbp0aJLi1qoX+OlLcdubxzi
/3wzsLf34kEh5Wtpyg69qgFtoiaaf3YF/6u3Ps6y6xSdML82QPqIAjDqkoF3LR/k
IXshCX5zJbXS+ugLA0S2GxZGMQPSiQQbi+iAcK4fMsE8bmlwSrVTNhYDNE5ohptD
D7NnWTqTUGmU47KUYQiWeV7XWLLosR0ykBmxEXm60/yIelrpM7LiuoBA33bW3OUR
Gi45C14vc7tmernRCTkbO33kL/vg1L+VlV8ZjjiMPtxbcTRVMdUVjVaZYlOPqtKO
eYvJvISYoyvH44AgpqAFIL91e3Rq949tJN2r3OqnaEgwSqqxEKtde9F5UlufOflh
zwz+odqSqMj+45/4DO7zmHW0iGWnFMgPbmdoXFnN1hXmG6vKyY+aSn2fEeJbKgC4
0a6ln0ri1JNe+X0Ue3/JSv8cSL8KHYA0h/4guCjSOwyn1mB/7BTk34BDgB3PSKh5
LQmUbZtYx5ySnWd3BJql4zQVAQyb+IeqCNNLMpTOuwvwC+PP0a+GTPmeYSTqgerq
g1ufnHqsuv3+1mqySvAzGQn5eo/Unfcjwau6x5rpzZJ89kCGJgqXl+w5iMgxRmzZ
QSrM6u9BxMk9BsjcHA1vC3JWH/EKw6+IQaDW6rKvTKZyGCo3T/iumn0Dz+T5hbNw
LCsiVayulzffur8EVmUFRJKbPksgad/68czuVLEC7oKl2LzsXYj5XTx2bXwL4qEl
pYc+c7x8EPR/O8EtuaVphL+lGb9Hj1E57YXHaIjkFIBK10fHurH0iwo9ZH0I8DOs
5I/BaXFuExPK7h74SRpuT6Ir38ybjoZydWA1LEjb2lk7ww/kCxKCIaxNOlmHdnJ9
bLwOEEX/IWz/b/+xkm5yqq84B7F+Kco+ZsshoWhRAZnivohrZBriq20mXcF64LBp
iIe3iI6ph3D7Y57aOaNroO2pdnoCenZhrZ+6jIjeCLTKmLKETGsXZewV8Unl+oC+
iX87lgKzl1pPNOgs6oSW7ZvI50c/hqPsXHYhFiJQih+6yYXWyM8n2FxjnPV640m1
LaEAcCnlvvLADduguokSgF/IMZxLYomVXbwWziE+AqAHBVaKcVPV0opsPwqE4By4
cAMMZB9/LuXAKRGOcgflX2ipsSLzeZ+1KcBcNDOugeMXrPAU9IDsN/2wf/4lmZ/q
+iWeL/qp9MQ6UPBDjQe+zSVukkftMPnYgXKVUDEaWfctgWc6/VQY05LiVR9q6r0e
LMgl3QAY2l3c9X9wqUuQJ6RcBvQPaVFi93pd2dawYQbvROKEI55xxJVmVICSacMP
B29Qa96DQ4PkG3C5aAxTTbSIPkEyid7aKk3U64a+6hFBezHN6xOuu/DI2D2mRcob
Ix3hDSQXgvM8sbwCa0s+0lR7DWNYS+IrZsE7a1F1k8mQDxoH2Ik/uF9F40jnGM6n
M1nnp/+fPaN4f2Kt2wVmilbG1RyKTgzgRAS0+AJjSbQ2R9yc7LcWfIkrcbhs7UnI
C1z0DdMqiLNcZN1QWfU8qF1oMRtocqSzFZCOgwJuf95XYYWEIvEuayxZ19FeE8ck
xIgahLUyTGvqS+2scsdl2GH779UX3dGSDWBjxwAcAGc0yLqgCQmQRMoDBpqxZTHg
XQhnpQeKnLumSkAPEda7W5/X3elXl61AZW+R4UvicBKUIfEj4qv7sqG047UV3hAb
v8VD6kIXqXfMKTB/hmNmLRapXchE96+GyLhIbyI5YwAj7tspgtiqChUEPNfxUdw+
Snss8n2Ymc7rJF4pG4ntCwmaXjp2ODX+QhQdvGeQi+Ck9zgclCfu8p1p0DCdeGiX
h5prMeIrE0aLJ/0P3Tpyyfd95O2Cm5C39mBMWZmI1GHhXkNZehwHjZgdeyqp8Gx7
2IT/G3Uma/ZXBS8ufn4MLXpivMGoiZbXpxVMSLqVM3BGU2+bNGXG64tqvMqJuJeQ
U7uLz7iUrbD0+VjoT5HUnzzo5hfYjJr4wAwvKFIoh5nfu5hJlg0w1w83PQMg8LyG
kWNeAe7U0zx/huueqiblP4DVA+vWJStoEi7NpeoeIH1JTnjgNnBqCGhoT171ouBD
nJhIz+TBD+5aNmwQNnFRbO7JFt7oN2rrrTAupGhbCXu7oipyJ+ggyWYXwss9skvm
6ql+0NKXpYg5fy8Z3t6EFRUaPLPWf1epIYvt+WcdBhjZ8XEx3dmJ34GtaTjjT6ae
pI0W0rRJxCooaG9GPS/2HAFViCcTaSud6ygKIQKj2LUcNOBmcoO8DeWL1IDOTTgO
Cb3HYNxKOyHjizgYzi8jYoW/FeB1gpigH4T6uvEJkg6dh0Xs/5MAbWXBJBroqyb6
u6sIgWSNfamb/r9oqTvNound3+IIrbfuoywJ/yqPdiLfBXnVqF29r8WLczvvTmBs
YIxzuZeB4++uR0UtYhIwWPxlxiSYl7ruqKlQd+fB42UReenVJFCzHYyJlRLCiwwF
pWtzL+WzlcgDM61vxvpc8k3W3ugFzDRQ/6IANw5wxhqO/ist39ybWmpz9ea6gZ2Q
6z3/Deafytz2BSHn9P4IYKJjmpBeIuJXeCLB5qCL1m/rlm4Jzdb3w4cQne1D8EWi
RHRvU0OTvIKtd2WVTNcVqSqD8eFP9TZYv3CJpSEyeoWk+hEg/QwQEnTP3mZxsTpg
kbxM7a3KT3gL8FtMNI4YtuplqtZf6Zfwq2dM5aQp/Jz0a8cwnWT732KXeHe+FM1Y
Jnh7dyKVJFT4hImdQJ3uCkUdWSDh5NS3uUkDg6V0S6EJGPu+h7+IyoA9rinrynGd
umHoAyZKERPuCbX9NPACG3hkys2soNNrdlP+j+rhAgIHLi6AFFrWcEn6tpOsTNe4
MoUexPoG8GU6dmypqtNrhc2JbPE4hmo0pLtuYpKb1xq/+RJ7Zz5A/NZ5BQw7ANJR
tXIZeRr8e6ckDGxOUxa4ZGneukQ6zCQWW2lJ+a4EmdozxJVRICz4y6ZETayX7c8t
j/suSlTlVk2Sj/YnazgGLsCJaj8pI1mKIwWC4DnaYRAQIOW++IfYILw0tBs8M5Sg
JGhN2XwL/8NzdvSPwnlPx2zayZ8TAgVGI1NUMxr+SLMDUoURv+uLdWqhEN9/7Ehb
UCWL+oi4vGNW/3AI47vi1obUbjdaZftTASU7FvWRugC4l89sROyxEql97yDh+dQT
Ag0exjxTtujknSFJx9AVa3wT0ZIZUvucjmkDo7dn1fZhCNeV8fN2vFJB/qfM69Dn
s82Z11mX9r4whfFxTnFv0c3YNeY4/fUZSuqeuNAXIehH56F1kD/LfTzxGoku7BPM
Jx3Abk24MkDjEUxoxKZ9b6r5p0YJy22xooUkZGmMcO54/O0dVld/kZVcVuyBjeW9
16w278j3Tox5pgecLqfMRcPriDCHEBwUtQYwhZTLIg18sO4tnf/oOLzPKxQ5jS+/
RJbxEXzN9fkg293iH4Nbvm0YjID5tk7QOa+cXgjlyL5sFS/63cXIXjWk7b0Zeuwx
Gs06JeugrTHFUuwpqpau8zgXDLrCwJWwS5UGTx1P49ASpNoukFKAfD7OQ+yszwbY
fCXLa/N71wgp14Y9rwLdV7LIGuoB8Rq5sP1VDIqlJ1fK/Zk4vdo+oKB+UFfHp7Ad
rOEleTiTqvC7KMOTnovI/UVOgdtKF0OROsQgbNZZ+R2icfCJ7tjQhvCMcZ3w24eW
ZL6nrxKWKzvl090ieFs5pbsnoZEj8HRY7nv7zcpAbb4eM/ALwpf3R+VLytTdvSuH
Um3yZNKK0fWV0qv4BYJAqIA7mkHjJyhQf98wvydT1PArJtsNiF5zQLql2PLNNS1U
RvX4SshjlTvk4LPAcWOWH4JGxGIQsWlPQDE9pGF4ne26+de/R4JHQHtU/nPttJfJ
IOvIeL/5kQIILxznBBl2yWs1fYHgoYRSP8lhfCdpn/hOUXVbDKlxxOi/IIoicC3S
PWLlIu1hntgwlkOudDN/CTVNyq9JAQfVAwm4ey+IBLc8VUoCFCjRNgSAulbVQqV5
ZPcYttHErz13mrrNcApfQWuGeDPoSNCC31hXP76WDJqTJCKO44W2q7SqhAJFavq8
I6/Gq3is8XBlWfvCWzhyfqg4RYbXcJnbuJB+dilBo8FBd0ty7sw1GOvsAJ81gxsj
0XBP/F+/LEm3Ru4asmCZYdDBsePwpcuPh/HwivNlh/QjG88+/6G2CJTk4dfg0eYF
ENVdDRHC3vKLUmdK2N7PrV2QG2M1ThbrLd0gkN/OldnEm4yaZ0EMnV6sptu3RL70
ng9uGQZG/LK8MwZL0OVQzKbjVt2hGQeKcN1hjdQQ4CR2ivH2KL3yWdVD/ujEMGst
z19H90jCv5CPVAwtwPgUUTJWwLi3S2MjGoQZwDhAJuQDLey89lR4mubgV7THMD68
jpyavogqEMlxiLptxLXGrHWoYMOUSVouvgtC10Kk4eEQ9T4c1SoYb8AIzv/3GX8V
pRpGVSSNmJkt9V7o9fNaHcD9daeu1+5l7jfkjfpOz2SpdygVoqVHW0jr6qpDKiYw
heoneC3LQNjRLjmiwhwJZiZPGOMUaAOMBjX24lNwCo3AVrSv6eQQTbAQpcJPLt4L
Swz7U5YZQqUslCzc/JZDjzU7NAvBD2FSgpeSV0PDGBJccrRmVfijI5Rp1Up8cGDa
P2rMIcT4KKkw/3PFnkdONjcYflD3r8HUsAdwPThSMgDCSc0rqFSn/YXuYLL/BSKI
H+yfMf5FZAYuz2GkcWcCreHbZzx/xZWrr6N2LI2D/8rbb1gYz6MT2qxVQ6nn9puW
J9sUhxNAk1YUkcR2eBzzITOBceDPsGYXxZrexcUn75VbF8dpOHOSF6eFweLFAfFY
JMJzmMgNPV93a/K9DbIi2jHyxbu5FASQ8zz/C0DE+vbqyUOyRJIbwi26tKaUsFOq
QmXY3wemHtNdYI7CpbPGCAQyWkpMfXIAMl09x4AWYHI9WUaVqULhTmbAjqiUp9sL
Z9zwylFrcX5D2rjJfiLRyJixkVtECXxlhq94X5uCssHxryWj+hdEhPBuBrc7K2Rh
zhpKgifT9owLYYC5du5271Vz0Oh+xSsLvv6HseqMfJdc8sYegQ5n3YtMgdeYO4o+
6NU+IDwb3vJale6Hy6Y6pTrF6mY2q7XJU89SM3OI6ozbuzm9eUs6ZF9yuvy4b4lI
z6dnzTpDhsM0BvvtDBpYYqW/HGezf1FwSgr6CRZVMwN7GDbeML2s5BG+qBZuph0q
AU10vqSwjGOAqpKE5YafdwkEV9D7+S9WIzjm9Ovr3ow9cIW77qP4uwW7GLuITLj4
yaIp53KIR8ZV4Ys0ROgyetu20V/Dj6PJ8Zp0lj1hBd9c+YWA1Wf+umqN4zmm2Y5q
CSszJcbxjVHgcWPU7VPPnLgOVyBPSDRByMDUEU5RHxKNgDZq1mh3Xz5lfjR179ty
s46yohR8WSh4Pw4GbGre0x5AleSkaiPfmJesqxVJhi3/5XDc3RMBSaaQOaunRb0C
qWKgTwBkwCjg3wYrMiRzJqvRyHpXFUcINw+Gu870K2K62R1rqWQjwH3OxCzCdS+f
mVOp2xhr1JGmzYitjuwiRHJon7IWuBcydiec95E61ZaZK+x6DOM7hxIbsNwDTmJe
ETiMWFwzEJtf45fPvti+WAiEoOSbGmVvYeANMl+g01guhCRVVKb5YDLHLwMaRi/v
dUujkCBqOBz690+ahhVatwIswZfs5blwCpNMlAFwRtE1YSaFLpWL7ypKauar5mSJ
7wMHnhjv7cWl6HWEwYrXyawzruFSXeOZZtAREiQzxgKEMykSEsizlM0ArpixolVw
lUJ+ieWrXpQDBKYWO4KRI9/PAH5dJMn0/7ylXQlZuQn40C3m4f4Bwt5c93YrZpsi
QpFdtEMWKCTEBcuwWce95BTi/HWY2/pJHIS+t22/q6clgu4stFAx6HgrTjZvDp71
7QP1GOoLIfECvd49jtY370cn7SV15RXglPknZh1Ijm0k1Cr5IjQZJovJh1y92NwN
A8me9CJCRMUad0I3k+8CS9WHHqK3K8w7I6s+t3d04nlrtOMURGxBXQ5TxVMk+lV0
RWRJlmN8VgbnSXjU4SBBh7arGOLyKsmMR4MOYcFH54Os+mYxY6HYi1uQOFaW8jg7
R3n5+cewk/DDTOqrOw5y/MuT68nGNPzk7yIcnHyIvyYW3dxOYglQlXH1WKLR3PIs
Gkof3MqNy7fUzxLyEpawtp1EJxM37XyW09yHLKEY/fu9XfMlPVsVD3T2x8Eyw/gy
NySYf1CHuFI0iF6dU96qhM83eAWkRlIh5hG2KEyLLH62rRFqBiGtFNiHaOhPrFcV
JOCd0f4KkfE0UQkP+xifIm+7hm6y8G9KD6sSWo+bTIPPEzJHfzzO7d3uZs2yt8HD
68GvEibfXnAws4D2jPO7b8MCmyuz6LRy4jXaQOC+AiBUb7DKIlTmxFvNS21fjl/C
B0EV8ImdI7rS9GH2S3rUjfZ0i/f27cj8OpZdSmwvh6At0WratxzQ3ZiEDqeA/j6R
lzlahDlMUCvHeA6i72S/V5L04YWKaCECCDd8ayW7JquQij2b6XWL0Jxvg1sUvgmw
wtD4E7gLhPik2LiVjAzhp0LBcCUXhiq4uCU/yqWQSvz4z27R4wUvZZWau6YWLOlQ
ewL5VzxborzhWvgCPRX5MB3akcrfi62RVBL3DtwXCYHbkv720aTZ0/OVnLSONUCO
FWfUtwUsmY+3FPcrxKspiejUoUvPehn9PrXnk5QP5SZW0CgemOHLgn+2JjwJfJpq
r97nraKabBSngElA/FeTX1sHOQX0tu94kF+AoTCljOvZYd3XRLP7fx494M9/OReu
CDefoqExrYPkLqbRoqntNB5prz/BreooFBGihwuUzEdEMPKwHUr/eV/Jo4kE+oPY
aHUcF942m2/MV0PK+WcAHh51NI/VbrWIr8iGzBf9erJY9PFxZ/EX6kCrHR/dmMiO
8hEDFUGf2AhlLY3dBKPrT9ClmZFvPyjvvS8JWI8PZ+b8JuKHVKNFYi8v8n3d7Hzm
ulkvJBlgTuHP42tpcp9EXfZyOkirDCjT7yWnvPRfUqqkVQQmVSOjsbRLkhIUeP6e
NjiDEADLVh57enHOzdPuIz/UmSe7j1GeB4mu9b03Tjzw0V7HLxX222fJe6AVfft1
NRTMjbx1ELPvsQnILPY9/Sj/qmtfI1qdC/I+MGQrKDMZNUogwEDY5KAHLjCTAYu+
I++GBZHyr815TOPrf4ETquI269+0iYeVPvGld/MEVdteVUUAiZjGdKzmVJwkc/ap
81STfRnAVMT9Ff31ffcQuQAkXwH7wgmTZH/COkm2A101DVUIFTAZUQLXfq5ExJ5N
fiw2C1p4X3ihYqJEXlYuOD9tDSUiNvPgePflYK3XNTEivft0zSIIQwPycGywGFv5
2najBqDYBZrKkvi3vZKTBt4OzAjOgNfbTIzb0dOoWV200TIPQhmz7fQnw9wBlkKQ
EmnX3KZO+hVb52JElQs3JibJA68pgCw78OopOQiIHksDfFeuMdlflR1CJc0ry/ry
ZzZMjXup7zvJrQguV6ftYgtJg5W24+uSx2pTAzIXQIl78wjaqF+3NkkGTerIwtlu
MHc4Vqv93kWdPODJkMTD/SmOuWitU7bDeGeJNLrNCHpt+zMwpNwTbw5jLV/3sb19
FzQpq5bQZMaOzFeUqI9oTO/XkC3JP+SYKiDE80LCmzAXrpe1wHLBUsl14boN/X2t
PuoGBl3T6+WKvxbiSqI/mMCEaqXEvydWUdaBjcKHfjRr4Y1EWnOy9ZVQrOLO+2YY
CkFKJ4Fa3nuYlkKQ3NVnho3o3Z/qyQx1hEBzuCJBA8R2okLKOyE1xJYtxZ7y2/p8
B3x9GrfADmE3iCjiOxGo6jJYkLUmcBQXyCy+d8leCOvc0xWo0Af3wFVt+JqDkezC
3skZ8URELZ0EqFg8KUTrcymxJqExABtgSrUdsn9hQDkSwjKT3im28Bae8jhth+O5
LU7l8s1rGgBslL47/ecyBL6e/euyohSMXrLnURzmEiH91pbRetOnN+nkZ5rg6lFH
FFWjZ/3H6cK/VQ5HIIqNecKydnCKDflrNhsnkzuVP5VXVOrJs1QVWlOxTzywzli2
v95JQm2J7GGLfY9sOFpN+m2/++5gd+P3ksMsJoqgwrQQ6fKcWfuBCyvk2KMMhe7v
ZJU6bjq+SsshaVvSotUj5RsoTdb2rAlp08gqUNnV0BbRXgKE6E7nrEPqyznZkYzO
JxQkBBLhkD5QuQeTqNOcRaTt8QH3jRAl8k453sG6fwt07kUuluDCszE1Mop8rSEw
78cNCg7tJoHTtEdDCCtjz8gJGrLufYNWQQwC84ZuFUuvEQKqTHHzbCQ/RHsCcRN4
dPIWh8aGHprcu3BKuzTtsyD01AMlu+yVioeH9AqyeuI6XIWwEtjo/s0xUaqxff0D
WM1S3cibXXIkRWZ/MZltSUD9YwbczLOdi4ZcoZjHZE85VgL0VsjUlVTXPJw/twiM
CdxuVyB3xU7KXwdSPmfm9n8IUDHiWK4ZucX398+bb1HuC5fh9HaoeR1aq0ry3PYD
+TSCrlhDXIEWvs9tUi6iHANyjWq2hay1wIfj/i2L7rv1fwvOMGyhFkyKD9djzHG9
SKqqt7lC+owyId21VCi83aLGUeEtNjAL2ypCrGpxNSfznW9jH7kTm0562/EMotDL
rdx/oO4dI1GXTSg74rA4l6vsEYOAouBTcBMqqj671lkFYYdnEgJiI304ANxo5ls2
8MXdgKmcOAbYXZ4ctQMSQoo6OvYpJdOyFFxThZlikEWQ0PU9Rk2NTZoOqM8tr6O5
5gVPZP8JF7iXAKVmBHGu8K74Qa3p9WyukiruVJXliE/3ls0rYgTraXLfV9Ncb5Nh
vxccmihAz3ZhWiDnbikTSJiWGyxqIAZ5FFGQwNJXqBUabd2rHJ3vB3QixvYJekxC
Rzk1zA56ZXB0+YgqnINo+QIF1xAUBbEo3mZ92cAGu5SEZMKcUHkpDX/vSfg/kVUi
ftJ47wc3CXObCpbEHGSS83zoDrifGxwHj2KOVKiMLxVSVVflfiYxd4K4qx+mCYks
0VpdtbojU+4jjrTwICqmUIj4fpynokwLSHv23Jgaw4zUpTjTBQIwq8l/wI2wzyGV
zT+dUvRQnoUJsCaCj3Qo+CUd5oT91WiGQI+deyZjC1Fl//4MAdCkBAdvZSUfgFgy
10T7900VFfodzsrrNFeouuJ6s+w53y1CeiahU89Hdo7/L1NNr9qExNfPytFuj4/4
WBuSEAOt/QWo16o5TupTeacQTw58kQXlXbvzUxZGRvTfbT41VPsENdHC7abj6W3L
mk5N0Q4sNWYxee66qcUjUS14kt6K2+m05Zir70uI/wSB3fErrO5Y4klWwO8WvCqO
cWMBgrqRmUJtu7eVcEbTRfFOeKQe2iw5VPUG23ysYaWQaE6TOXmG6TJPR7yRe+N5
Yli+BSK3B5Wo8ToNmHG97Gw4Wy2xEPh0G6JIN+7M2q9UpcjHOYR3qgqeyF0FAqJW
5ad4j2dEA8C8MdLq+/EImzjnSX7LYvZfOlcmR/s4351JBWR6Scul3QKTL6+7Y/kn
f+Qq2Y4SK7DzvPaV6o7Jc3TR5SH6ZMolFtTcQDIZ0PhAzaA7RQ9HKEGkFF7uOhM7
nZoW89TYQYnjVqpHCkltR/Eo0E5+LBRKBFsKGf6InMNBc0IT7hnfd0z/Yd8jYSiA
REPZgaZK9J1hIPdShy2fujImE8iRc8A14CLUYlsSlood5W+zFxCkiYnY4a9/oM95
gNoM6AHiKiACJJEPvsThAOycMb4WG5C8KiAhQFnRY+nL85QDaX8rbzL0S8nrlzvd
itINP3RO3/RCkRP0RGEzw1Fpm7oprayekmzf2C36uu+nhjfxPl7IP9/VjuND8nP8
9zGoIJJdpgSw4aVPN6wZmes4YKAFTC1sRwXX6N9/+huuDD3wrC9y4YWrKjmEq9du
pYaXBuW1kgFfzuub+rWRwnzl+CvCmO7X3hjO1yG2KsoDNsvA2xMuxRZORFD9Yzh8
kV6zT2RupBOfDvwXXNiqKqj3qQ3Y0trdgKL0Ess/TRRVSxz6/wnJDXJEMQKNB7ak
JCF2hkCwZndx+ilj8qsF6O7t4E3fHfCSgobSAXWKFAhJIL0KcQr5CS+yYYNrikqe
c5bn/V8RQ70tp+toGWVEDuwXSB+NuTX/h0FzBcYiLAxzXDPUneLSMPD0nOmsDEHF
pSv72VVmbbhNQQ41YAuEU9fPAkbSjyiCC/SZbWe+YFjHi7bEssIj3I57H/Dm/WlS
Zfa3EqSeEWnYGnhd8d2fIEtHYCBuMM4PPjoNw3h+uyZQcNIMqH6t4PG0hiA/k19h
pAgJNhTiqMfprnmQ5+fbMH4/hhWotkCnri4ZJ7lJOKEKdhOE+w5kHUBJcfi3aLU3
kMCsyNaEo+VOXHtTTHIIE+d09yYu+3lcWUS/8GpnHSqqYFd/eOx1WouwsfLeq6h/
Rp30Bd4wYadsxjCAVsmA6d40T2gxyUxFeCeEo6PsOYMEHK3lDL68dDBnuq6+g2Fb
DF+rkXcwceNdtNaRM0c1kcJv6lL3CX6KHQFDZs8+VuiL18sII9y5FsnIISoU7uYU
uvIP6apQrSPH+yYopN1RuHX4Hm/iSFLTPJZRt2YZTxjut7UKuVA0pEftYKbl0JaZ
ZK1+VSZVgtaNQz03vnYubqLVohpm4U8TI1L4DHioJyCi5KgAWjGpYfZ1BK8KGQVd
ymCrZzJVtJX5QKZABVYAgswfnm3SAChOGpKcn5FoEjhGPf2wPjYTLMIvvrcbxbhA
5yEbl7FdjtoIrvoshjQ4jlWtcF1NP9VbcEUOI7iEtNSVrI09WUXZU1ud8ehG/csQ
tO00mrLRhgQT34MU/FUQxrSP7osJEc/lTpJAEYZR8usqWKafmUubfvhnrsQp689+
nOyy4zOM6o73Gbh9Sqw5UXvGiEP9K3B9V9+KIT+uT20DU1FRQQ9gV02SsHVVgX3Z
KN64cyEKpg1sZImwuQYR9dBuIXRoTcXt79uJBputwUP3bvkQMmM1OQqvUum1VjKa
voB3wV7vg3nvX3S3N637Zidht1U3TJDIhonsQX9Ab7ztWm4dcV8wgI/bNbrN1MUK
Y+SeSTmSYPFwgqTLbAg5rMfwB5LEz61aFoqhUplpI+lwChslijisqKd/2OoPHM0b
9XkmiwG5U0lpA+EGffZbkvaeyqz/kdyUhq+XRL7fnEaLy2RcwYiVzobKYdE4T8fm
351SkWYsGNuyua7HfsKCGw1Q1JckB9P3rzH/gI2hg+fvEF6Gmzts127s+oGUxvKP
cxWo1UP7VkozLvW6HU5A8gbn7X1In5nGsSDzo2rlIKKwUmOOnjqFAETZ+mA1pJnk
k/YuPoevVX27HjrLsBgnDCtDg6GlpyfPVkjf4V0XegHu0xXa8GcP+xTvbTe0r33a
A2fTCfw1BJwJXjQVjiAW9tffv7nlMlOk0U3FXVm2Vyox4k8Dw/6olfNy17dZrZvw
MXKcQN5eeMM7+MfN9xYzlP9fwE3UbvkEJHIrdR4tMq/U5rkfjyIqGgWPSR4RHC3o
Yy6+iJVYydv0PidGOEOe/wkL89Zdfn5PAuKdB+C1K7hLxll1L0P54y7fAJu6ficI
tVc4tpUHrHKbBg1MaiZ2uqIthAh0RAqNzgHC0boamgQIKwDzujSF2bqTYjydQB0W
ZPxzoQ5sRG4k0UmFjtROKU49d3pu2U+jKZhPnBJFS22e6R/pGp6MW40FMNArZjN+
UkYoHZ+WoO8JLSgOr83xud/Kztt6fgevnyWO8H4/Duzg4qiy054BgAhvDuWsBM8B
0nlB3xyyyHSF5RNyOT5suKYCqtkAcxiDuYrs5WAE4s2Yl40+ZqpHZE3V2Y4R5Dek
vdVjPeLajcYspGjHI2bZBGWwzG60qREsN4b8qieCDL8fGODY6+1SNeGwPGSiXgew
QZRf8nRoIbXqoYYaNGHUIj/NJ4NCzhtYIptaIapRbgMar4US53HeBCDf4mtCr636
ci8hUkOEJaizM5FkCjfZDmhSsZqm5AbIw9aZOyXFwYRM+x6eoWn+SbB3K2CcrJgD
udwEy65c+M70U0FQ5TuD8lqW0SFJ7NRG4k1O09VLQNi3r4rxUjrCrToFAk/YgYDw
AR/9QN3w3ksvmUVOtUAKtALo77G0+0ul1s/I0NS2hMpI22cxEviNapLnOkvtV34Z
Nsc9KGAVcObnN19MG8QeeYW3oCKO8SwYnmsR3fUNjjTD1cu/odBP0x5sKISU07/D
7WOINB4RVedRV8YuGfMZuSaYppVuZuJpxH1RxX9t7vWzzupMz//KX+jeQImg4cNQ
dKpzxXJ1+UQqD3RLkvr/eeKdBNcLp0x1lMUFDE07UJcG/AyIe4G4twUv42ELoePt
YtijBPPqfs0D3CvVFgXEMIjNLI2XbD5U1xaqOUuzD8+acfo2AxZnA9+Bf7MHbFHH
tIrPDTGodBfnM0bRgEwiFA42juBiw1wy1m6vGoHT8q7Gs26eVuWg5Wv+AfU/qfMv
anYR/2StJ5beUTWMC0HkShoblIsGVwmSYWJvSVFzwrvFVj9NYJA2xaMkyjKpFbzF
tw17d0Yar3BGHhhIdV+LZpv1ErXygIBLRYiJNaLevxtL3Qh23Z/FzuwILNpxbWXA
XGC6aKBPeqEO14ECpRlUxtWEnvWkSJO4FaTZAWQDAFbQyCBL5GnO17Tr6BSD677f
7ZuVJlZzxsyF6uXo94H0N7A8UyFMJlacOZYH8AFjajh9mDybZcS6BLJ3PT0BFmKn
aS5uAcOvyRuC6sMf+YHOkEg/iBFDBdaao9yzBA7yGiaBYzc7tuUym0CRnt3FKRMf
s07TdkSD0HM7gJO3aJeXdao0MO7P81eO0kXglSKkWSuFqO3IqtF+DJ8rT8sYOx64
bBN3jVW6lejzqcyoLktVQIawfGBqfL+Svue5rQo3Vzk1VzZVKpIw3aKZB1BZlqMF
HsUOdFImi1lBsmtll41fZDNEdHE++3UQTrzV+iOOKBNjh91czvJbP0yU/A3XdSCb
3BrSqoHQpIMNR3v98Y4oxSmUhzQ3KcUXnGUgdED45FbPCxShjbQjNarUQgaydSkb
GTxnTGLfEpeHU8EJ0Yi3RjFl3uVwk4VTC8Ot8v3OYm/mPZGhK1RYgdZWzLzFfSdj
XKK4x/FYGumv/jGD0R/17sCdU+1XbePgxti7gekGfZJ8ynnxS5gjd0Ub9vor6nDp
7EHk5Neg+wgR1hn3gUJyptWBgztrAQaPq+2rMw6kzRV1m0TfXL+XxyFs9q5IEsn2
yx4RhAkMiuwP0NGiqmJUJDCH0CI9sEn16tUvETzbByu/tukVvx76YzLkRh9aV57J
UCtxrwCmJldLSzhfibrxdxjR+19wuX4o0XuaVeM+bWcPx8kMFIDZ5CdVRCR2Ok4f
ZlJBibtQ3j19TcO9uS8ou22uDCcEwzBDoZRVHlA4PfwkbpZjTLxWnWG0BETPeNij
7kSaCm8VWx+1f4Vd1epFiBCREwBjF+go3m46Up9OpLb6SaEg45sdYd0UUAo5Cocc
ueWoTNOK3cT/hHa9bDTvMk39EILRE5eFlB3ki8RWExafeE/u0Dc+T2Jh2Q/DOnLX
as0CGMyPhO9MG+yDNaKpcvtcJuKhUgDYhiAUknNNxxJ56H8ZxwpscQOmQA9xOEm+
1IvSOc5yu7YlF+RKWzSUlssouWSj5VYBCKb6+Z01EWtY+IQsiMT4scI09yNm6bGC
yFp4Mocn56gbgqfJ81auXNSqF8S+4SZZ+cmvH//Wc61xxmMFWc/G9ELDKvHCWbIs
ZPFgXuWkUiLZcF/+wRrDuNrBdnyCOvgVF5ANsRyvTfYQmggbhZf0jI2/v3wlz4C6
4Ob2Ak9D7HmZC8mfIM35tRVz0xXjPqJnkAp2Hb7++XerhkAFVhMyKHLOXrAxL4SQ
yVLD4oOqw/8fFoNvTx9awU1GICaHcemdQI4aG7AmBKCKSocgMiJPb3HnWOF3mmSU
JBVYpc4YPTof6nydQeNvKYiAaf6QKYPzpt5dCNJvzzWBCsF3D537NuAs1aU1vWhj
0uMAYr2t0lMkm5bdaOB16cFh6NUZu+tjcPdN2QPm0zSnDYTV7tdu6I8jjO9oM1Pq
8iEw9F83xWbqlKEvzhS4qQKHDIVL9OSlVzgWgjfebLOsaJalEGE5ixYRh3YbD8/H
wOg1xl9m7PtAdWcshF2K8AAVFUhauav/TmBsEjBZTT1RbGumA4QbpcFfYCGCVoHQ
69Syw0P1emctIAAyOiNN5EK28dsJkpsYrMsHfxD+dULMqDQx6axPWvS7oP72MgnJ
rJu3JmpSSiIkymKhk2PtXL6VIKjtficjunfFiGq+kM1u/u8DMKbc5GQQeLaVUkND
287gHnT0n9V2T7KMVGptO2/tuKBDEsUMrxtercPSFI6Cn9stSxBhijmiEdO+7WnN
t6+p6IIXbngEcqytoNFBrv6MbkqXtk8Jko1CS6DkrT5rueTiTL3af8ITOVkNwaOn
5G2v+aq5gYr6f5qlBbDhxDlMKbc5C26PWWXMHajQg/oS4s3YIQAAeETX0h1yeRuN
Tm03WWddBFe0KtxGmUH4mmn4FUG4KZZR8vB/UmiXEW6MmyhIeixJPxQ9kp1kN+tR
ctf+XLnoj2+YpWemn/twcZyxry8d75jKwCaH9Zah1n7DlDCW0775uXMa42/HhZvm
DdT2jyKIqaCqGIsWcgOv4Bi+ee+YnzIgKCpKifkl70e6JaPrjM+8NmLq5q+8GGB0
m43MOC3jdS/Ss8KZICSOy7XsM81+IBchnnXzJntpOZUefdL4KQ9NcYVpwNaX5E7Y
/vnT/TdicuRn5h/ifhiVLbHcewFl2UVUhuolrNhMXFnytxOOHPOie9vi4/PHBgpn
wTC+aFRPcnc/mCHKUdj/Y2vr/x52aZ6wQ2pJDM02hwE6RD7PZw1S3QEqPY4wMw6B
PFVH9A/aTdpcB12cqkqXjee2i3HK3A2I+/PE4G9ZG8SzWMhUWqjrqY0iwh39yy1T
ustkdJT9Tcli2360qURXUgvuyO5ERXN1tvDWZNPfRlV6SEcJYWQm5Ni4eBrSSW8r
kf+LNFRUDuwR7TGDgc4y1vpCzlOHzDDTfkImIJ9O+oQiQ/MT6Sf1SoR+O+Ttze6Q
UTCATCLQ/rjD0DXVvQNpSyLeDVfxIR6s/tW+IYmym5ybzwWtIUKhgMTvtbVmp3PZ
ALN3yuMHQImKrbRju5UGt8defBvppQhDmYLP42maOx/bM6Nijgp1WyHTYW2ogmYb
loGOoiHMUcnU6vITIBXmYWEZdVYc9yrytgJ+EiiQ4vsXDhdJdbXZIJPuYdGxHWHF
BzkIemFIvZvJ12ghNBRIBTQB3rUHxDVWDr9dPBokjp8I/17HCxUJ/U7OWAqPZYqS
Nxc8Utzb3B2+QnrYNlxvUFeuJ9edlgBuLUfEXdIlty5SYJbPL4t2/R1Rtnim41Qd
VrEBw76W/lXUpArNbM9mtGUKqvETMGTgauuZMyUit70WNgvVmoUlSi5dhaxF+vYf
Lqkkl1p7MiEumELI/hDRHtPy1xK7/ZByjtsoyMwrn54aEiItJpmNTBLH6Ciurt4m
O+LJLK6VDf8YR5g4gNmxJU6XmcbH6p7gI92fkw0n5NLoLSKUYYf0tSc/EKJxl0DV
/HGEcjs4rNkyqUE2zy3yV24flIBjPMe4ObWJsIlg5BkN1VpQW4CJ+Fbn1AN+9JYP
Vi1qxoK3L3R3y22H/vd3b2eCw5V3coOV+eg7/BDZAXzy2UyvIxZsZ3fLoipYIS2x
YArmoZ8Dr9Xu/qQD7OvEMWlbLPb4VeLA4cyv9JV1VuzNHc9ZkDNL4kUqLaEuuU/H
8L29tn3+EPNfZfUWc5Wi0K+ApHI81nP+h4WU7StnS6uqeqHiST8+ieX8DTBwyGOh
uQgCSO+MsClPt5dv37WWN4akY6JiWx1w7mt6/BqydmGJLuCF08HqOAWQ1vAgn6yC
Tx/5lQW2gMaalc63kX56FJTJFRrsoGEqoH6HjVEAKZqBfI+Oum8zAMeWggWG7FuR
Q0HROp+RqqRDsOXQnB+1EHdv5t5GPK0D5a+Kjo0wTeK+Iq9Rq9hntGICsfTTsPx9
PGmwqDZX0r5C90NdvX5NydroSmIgaK5Spz0BUUIrHBBo9QxRrRwrJ79n8WDla8JK
Hp4Pla+3ZFhjdgBIFQOOXwErZw7UUqF5hUpjWvO3aLbfMsRnbNPJERKBKGgCsRT9
+r7jVbZvtgZNzMDShy9INz1h3sgx6NFXw1KCVJXZV9Z8MpyumO5PAJh17S/PglHC
Ez5MgR5p/1Q2t4KNGLwl2HDbHHiaxXrfzKTKRh2QJu7IC1lCFctuZWu4bcwet+j2
Pn2QVYvxSaHa7/SvUd9QZ0NLwaevYQc5yO2qJMa6E82TZBX/ZUqSUDSirpjW1duu
QjvT6UyfYmebpkl6/EATDcmKpkfRf9V3VgXD4InPDfKz6aTXFFj5IpRynMs1Pjtv
vMspHudyqsjPn+d13OETMXrmlhBowmVLXcc7G0YIEOoXw8XXELm6sk6uvraEPkG1
7vPjI0/dkoZPxg3bOtbRxosHzYeaLa/Unz3ShBrJy4p6OO+UCYypWUu7mbxLELvg
7TEbtWNlGCdrktu+EW+sbGmiNEggbDhKwwiDGUhhitAs6ypfA+TxMII5YZVVmhxD
ELkfVSA95WPN5W33w/X8aVVIJYmVljB/AarVnIrGy/2dg+v9kSbrWiQ6kQt6QNQ+
MH/6e443SzqLcYLONfP8lfEI8z/wqYpLJzM7HWLIO1QcrOAU9wcmNyG97oOR4nbS
JoFGL7yVbdlFz3znLQAx86UZPD+yzQaeVzSUrOEu1EMqtjmQZLMiUy30/Ko2sY97
xEG8ljhwlP0N18b+OGVBETKHGrtOxwINx9F7BfX5dqo7f9765aq9AQXZ+YLhbPOD
/m1ZlR8BuJ+GLMQ6ltWcy6/A2LAgTZoTYN96KCwi73cegOjL5GHa7bLecc+K/BJG
Fj3/W8AkDXW/gB047PwIVbflXdsKiPHXLPMJX/c0FOezS2pfIwMyGJcHDjCCnyDy
03XfM3LNAk0UmyKTFtMl+BsX/+r/8vaIdTmhTNIkagQZ6ElzirZuoWYirx/iTdTF
XanqfUazNSitUvmqg0hIM1+z5xLrTCLqCE7CS7S7ofhf5GPwRgGztO6n85sP6nYy
cDckakwE3RSCU5uGAIldkIxcVKI9DBVyPqfgW1rQUGp42Ln7Eri8IBQ6NcFLDG4V
PDGdi1Ndv77ldKXVTPLUOuI/y4t+Jj/wLcMMjtzKiDU+24gUblN5YTZzRl6CLW0S
rNtfB9GkmDSEA+zNJ4F55aknBSK6cESXMV5dwkPzRcPKJSixlENg5hyhLaCXd9X4
Y8doXOPmie9j+yrEiaFKg3/4Gyi7T42DaQBw5RJQimFk7GaWat1igenJupELeyYD
FG2eb+W9GfjCsXuh/IAid2BhlMhb3uOWiibtNpuWIxaKiQU8VWGE0YYAZvsEv4kf
LFJ/ukFcD4KCme9Gwqz9u3jX6VkAhHLP49FAfgLz4s/w/TElIbDXzx03oU+T77XA
cEIDMU97+nMp2O7J6A6frjmKXC1t9FXYoR0UlUZlUQ5KxybWgVPK0xRg4P0U5SMp
dm8t1rFySe/qX3qnbep0CsaKe3Mst1UUTvh86dU/5SsYDuzm3nrJKzVdepCZ0J9F
F334vBfkdos06kro9P4KMEaOXWEjbI3keYfxnNrcKYHq2CtA0X233KYx2VW6l7wx
qeyIihisXuoviA+P54MG2uQ3ue05MhnxlgzRAt20rk1zrVJ2mSp2AC2tXbV9IGM4
9q/xCT6vmEe3UEGGUsOooRteBaVeJTQhqUAux5UBIZwV/7KCTn/XAzA3koCQWWWJ
n/FAWmsbtA3Iz9qt1yglSlnY8MeLrqJXSp2yGjntD6vDEYVFuluo0tcVK9D8Ck/+
LQTivl8v6mBQccIT79SLngQ8IRuOggCWbwE+DpbcNeZzCbMxsCRPj12J17Gthqi4
OiqNiBZaOHBOgenIuzQWJ72mrAEJSiXgKMTRZp1wY6nKSGfQU6EPsnD4czcZJ4Vf
tG7gxIHJGLKLWsdLMdegEf0ARQK5TyqsDHEGjvqjtJ3fWjOj2MNWvjGDM0zmqLbX
ei1HQEOXUrr1ACjds+M2NbQqE/QGi9PZVtOHdWkn9kXAkVlH3qx/f6eP95GUH/Gr
6lhJUHGt/liL/O9TJNcZkoSMl1UDofy3X+chM1SIjcmzfQWZqlSqACPuD+JpIi5a
RagDwrJ808XUJN5rvAzKRW+ql+ayDjSF+OUOFQp14kn4wjh1PVgzcgHwihCMjLZ6
R/lkRG3y++/OxRsODB1bSmRfgK5IpgcHJuWHbdSvbc9jlgKZKVCgMNQfo7CKJAjw
+a/3cYuRae9W/I5WywN9AAavtlgIvXYYrutQjfmxQKXn/xyq5cp6uUciBiZRPrwk
0nXijuGNasF8d6oCN/etl9aWR4MAD3mS78+RFlEdxQH84dcUStJXxFsSDe5Ve5g0
L8Kee5v+DsUGEvg5MSnNlXIysGH+pYrLfrC3Lz7Z+xlJxBqWsqlinN3iE8alSafk
e5wKC87VN+20MUTO+mcPtc4+mCmq25IQqlemWVv8dOMhplX8y6F1Xt0KEi935btj
hBOP/apOmOWKCPTkFnCM4OMHBK448D7XM50M2Kj9ASyawX6BXW+FrTCeGZ2CWHGT
qpXIBHRzxXGTh5Eie3NbLpsyqfpTtXF9sTU+Ke39XV9lCiw5ZdyNdGehbEhR3kgA
18GdIYD7QYNXWkEryb17K29ONRx6Y8WMSMbOqKp8joZs0HXFDQ+rIRznpfk8vh6w
WZx4qhMhtqcvLIDUfeB6PMOAgjYpku1YS8he+1/8Vx7b50SuzVv2rC3Y1tSakV5D
rILTSSgGrNv6VIkP4H8ROxnUcLz7OcW7UixjasoknCxnetT/R4mXhkx7slWg40Um
+2iRU8MoFtSR26r5eMLjQ7NC7y4D8K4W5MgR870ekoDjx6W+QFL5Y3pq79LOkwiP
EIf5HoAakC8Eaa/oHi57aTzEbeSxDYPEeP5RFLI+ZnYX8dfJ44eRroSKLxSzK64l
l228hqWW75mtUehQ+mui+YvltwFPl80L+60JIxZB+zuaBV32DXvRvhglHIuhNLEk
H+zKlbNC5P7CsEhQZ9rN7PyMcM/M2i5aP0R0K8SQ896vvk9Ms/GdBeW3+DoLBgBU
7TkuA2QOG03PA38KYUCMvzeES+/UD3nk66vgoaZWkaYX2+TWEVjQ+G9q9/U42qUG
UTKS1cUoTdJuQ/D9nIE5Qa0/d+RigktE3tP6SaxlX3dS9zKeEj9948EvJ5zeE8vp
4uVjf8vBrtswZQ82G4L0LX5Ce3vnlt6PLJVW1elIwNRcJsmvoNckNvU1/OToI/Cv
3g4dFhZIc32QbQ5cEcLhtQAwGX51YLQwL4LhWBTQPW0dxFDr9Kqde3X5EmOaVMFm
8kEnAt37+V+v5Ubdk8cTWopvkISADoIH4Jug8RIcdO6Nsj4aVw8bKsAedQrCTTXX
t6Fm3CubMQVRa3wLVoigN99/pe8uwqoi0bV3Qlwqd0bFOgW3WvdTCxmdkhYjC8ag
mH3bwiY5mHRkVx3X2sNjO6QI9OwoZppHNSr9d5sAs4EnFxrLbxsajTWBBbbzP7J6
035yZkGRhs7zMk15iscCYagNYF/aZ4xuznBmwvQeJf4LWBxoviapoK9FPwR0xA4d
Hj6E4fCKb6+pbj3RZG3VOdSwDQDWEDk4LLdXuDjnG+a+vpwo1UdlA9P0+IvJ2aRc
xLFPLt8UWtwWhS+ScaMs4k++FAKwQt4zwPG9s2PE+IrWn301Hm5ezQ2yOkzahdVW
SgqipVc0DbKXV3jfG2IaAhrzHLYS6SwQ0NJHPXKJSQjIAnUjAvUeeZxdF9sIny6x
z/Uc7n1mhJkDE8OD5zfjtdZG8Iq5Hj54WwdYmNw0nQVlj0pg/W2Y5Y/uoV3XAVMF
M68X2FzayDjQ64t1INeUC6LY7RBE2IrnY8kNk1ruWzZX25AWttcj1Yt/HlxBHvBe
jQxIrOIJE3RQ+2U0PVQfDXLiuSw49xrLrm2yl71l3TMI/OYJXQMuv1Up9Ml/RvgI
WgtPinlOI+z3u5eGFKcq5ZZqWBKwWGN57ZuvTobv9nK4zUlX8fEOEFzg3XXtvsLv
dNv+rSFYMB9bsCnVrFwzm54oz0WrIxQ6zwWyOmq7+xWga4E11EVtuL1anOk/oomV
JdGIifLkMIBRoJCGEPLPVAW521w9mhkhX3ajO1aHArXjLTDHUa6PRVGfY7uczEvy
tbYpPzF4SpfdcxEhWdaPPEBlq6lkC26uA7vybEJQ6tiKtkTKtoiI18I/UGH4Jlz9
Wfl+1OnwA4XRMyPSzKP4nWdHAIuYhSr7P1syhLa7aamU0XDUMYRjr9AJf4iXQZMU
iddY8tDbV7pN3udbYeEAdzkBWoXoAzcjteYRPQ61dXYySwFHJIiY6PJJt/q9OFvV
+y1DhoCUhowZeUXgK9c+0RvD0fVNQdXFgoaAIvzu3RdUEfS5/OcfNrhi3Sr3rWSv
wi61Ksad87nVSF46E4uiR2N8c6dUVzzW/IwZ1iFj+oyPDdxPiein5gDlzw9bAx77
3QGlcdzKrbWEk6MTXi/rti8qqiIyZuyJ436T9cRQprEeB3SMSuOiVyfQuxwh7OgJ
93wf/wpb2EtZ4Q5G0ynunqm7jRGVkh6aDi5Z7AquEFMzskhRvBOPInfhIfCX6u/O
6UPH+wHQ9cOd/LJGyRegWLazdXORyYtfamV03oPmfM8SDjhcg7J3y9RDqcQJmvfp
MMRLRduAMJBEDdGsWAZfREFrjHy3woQ8CZx2CzhWHO+gbpejYRvrQVFq289fMdHb
lIYgQYGp7I5gvIT5YrFFy14j2vRNVkY39jEmrZroHl6/wk9ZHcF2ndsd3Mp1vEpb
ZhO7m4l0Q/Cn6vT2xo3dSwR2UYKxeG4x4nUuyah1zFYgaI40Egxgd/AdOIQuMJ1q
i2eI8DuuccKf93yXbgDg5LCTdYug/uLj+aKS9MM30zWGqidT/TT84sW+6sTwEa5D
/GEaC81E221VS0hnXoaxZprkwUf3eOKiXNIQ06oBWLaNTTOUo12GZXXpafjb13zH
56RJ88bNqxq64qdo5o6O/QoSd2TxMkwQmItBkJlTthxUGW/AIcDff1nztxwv7a1d
re+nkc+fOLGy7FbjvCMKFjAR4t9XD8+8eFH8LFBI8K1olC4Tp8Dek69+1lDbuvV+
LWtd22yaPw6VoXBt11y2zAJXBET0Y4bMZk6lMErwc1tlTozi8rsqtMxD8aWuz/y1
DlhJITvpVCQrud2BXWFpBe4g8D1r9T4nxnYnqcBYWSF2Bbk5CD6xS09u3Wp9XX1K
+Gyi9Z5a0JzIQpwdPQIw65y0ROKfSecA6k0m2GRGTwPpMX/DHbCB+blynzbKc/f2
fxzQuUW0omyX+TiGtHYWESm9yJ7MEw2Sx0MZ1es6CftTMFxUB31zZmfad4H2vTsn
K2FPRhEcGFabWhVtQr99yTq4jwR6JHX6/n1fiZHlGsC5OjZ53xPXrKRgJ5g0A4xL
oh0BlYPV+GKyS7Qi3plnyJDu2Ksw08U3itNlY1sn15u9lzHnK9f3tfTYq8bjLT+J
7zHI51Fvq1jtfymIJ8jCevq02F6Xl3765CJ1CWWX3HXhrau8bwHranzz9svF9Z4z
gos3PuSHHhilwohDPk16vv7euztRJcSPQGF/E4TbESI9E71B6kLpdvnHA1+yO47s
t5OU88Lgva8XUqQcTN9ShPpVuI1qLeNcoGYJFDug58DyLwxihrbVd4T/FldwXeLF
ABzbxeip7BLTswargU+mu4/jUVRQO+30yqs7toXGlnVEhH/x9KZ490dlFbbliJO7
xxhNzNX56mkVerHpo+K3HD81YFvpA57ED9z3/vEtZTe2hn9ELe4rRfRlN5iQimo0
ZrF1Mmbg64QsnCcPWwaJbj5ZR1k2y7w/1Yz5ncHFxjmIAUd2t8XBp5dvmCCXiNJ4
nBNkbTtkIstFv+c22T+W9Lsri3B01jrPjVqJXsaZBKxbsQu4RE+c8FXINXuF/SiS
SSSUhEjvuGUfbsbbUZ3eQprcD+66e+iPB0kP6JtD0WaoBefBsGO0j11bfxV0ZYJF
FC9Ehy9Fa6+mGL+yp0Mb6OFgVuQSglItw9ptdqZVAi3OdEsXJ6UEyMb+qVrYumC2
e6SekAkJZanQQX5If8o5U4EEqiEI1C3cP2OBPGJLK1kifapFYsBUPyiVVUahraLS
5QM/eIfZWAgMv7UJ7hphixbLzAhyMgyGx0nIEYN/BS6zui/0xtDAku8yD/cP4wBu
OfGh06UWOiiuXgsJg9FaUF5oiKICmsUGk65+uSugpbNq4JoN+ylw/skFr+b+fCyB
2SM8giFbIkvcSx4S/UW3VNGXnW6VW2P+CPaI+SWLpQgx3gpTSM3u0yL8LFJ3G2l0
AvGfkey6PcM+zQe4zp/smoy07VoWKwJipp6OjHfdOFeqTEeE6CwAAmo4w3l6Tw2J
bUHPQV5opXKkrtqCrKWAjum6QE1Cm2xChZ3Eu44NSpr9lDmGGVEhbo8gf1FJDyvU
LdRZ9yYqnogny03NzVsdmGE4KDMBfY8jJWUW8tU4BUhib2+5V9kCu0vNLINI1zp6
WvCcFPmgK+qdPQN4aMJ+ohqbGSyVdD61G6DvrD/EQp0W0OB54HDmfpLFkgweDJRJ
GDsvFBdvVwns4hVEEInaDCTA5no0xYAvEJbc4uFTujOq/GAPV45jVpBkiPjw2LMm
wT2Y3L/mh/zMIZHruJCjijfzUw1BSu2vXBwAFZEBsq0iR6r4BRKZV8FW2PFy9mZW
54gnpRkBaDUw2jgO63OUB8izmAUMfsaeTgdJJvgBBn9RgbLB9WfcYR5dY2oVMW2F
IQ+xuzCcvFi0JovZUiUFaZqQ4DXEsHePEIy46eS+7Kldmn7SWWBET3L9lWtT54Ie
qsMW4r2nBmlbbwBk6zoKswDJTr/0PgUgZlXdF9H7h5nFaPUaHi4O4l5NH3S9o/FY
VPvuCYReQadtSr1bemqd1kfkgfoNT94FotxA4bZxuSH4wi7Zs1VxgTRC2WWojfcW
r9Se3tITRgrVfFPN4I//N4vi7PHpv7O9Dd/DlBwBAlpus7STfsOx0snjg4nE+OKu
0fz0aDnXuZxJQ6cYCaeqNAE+c8KVa4MKimvZheLUH19cxG1Dyh4yfQhBXnSxtcq+
F+AHvft3w3Hv7boF6WtkrxgiE5rPjywj6QfBenpmad043ZTToDY1h7TA9pDoLeSK
6jLAllxlCKaSxcBpNWQutx35vsSQmEWGon/eZG4r+9lHzO0999XDl3wT1Ru7g6Oi
CYa2v9CYJnB0TbyIqeWenudxu20xi9+Y7Sit8dY6p7TjZs12hHrLxXMA9o8fj+mY
VJkWTIcMasmZpeOLlj+mJ8KHmOAm33OPGK8QgGtsrqFrj0m5gqOEIwKgpfSyY/z5
dHXRb4ZfhELnEmocHNVoh0vKReRTD1Wo8zcTcujJl3L9hLxkjA8rYAsZ5DItEtKb
CJm4ALn4MzJPmylLYWk7ocVg8gQKu7rsXiNECuJv7knJEdINe9yF5/KsRFFUco/7
/C2p06vf4a9gqBXNgsgU/E0lYK2Fs4wS/gaTdxm0HDkX899WIkrEc7hqzL7xlbfz
pQxg6oSNW8ds+eQ4wOqRiUhfY/uUFc/n1gGlAA9iTjtxa+VGKRPd6dNLNjwkq+Zq
Dl8Ef2U4RI1D3bKrH/KHwZsIf9WetPHunbFg9NIiQM32ab4hiKhAdMawWlnAXCVU
16ipIBw70M2Ps69U+soUF4LzcvhiG3NbH0iE79wA+fYxe28fRw1EE+ARXubk0B/3
Z6Ju5JoEwY2ZosVE3iojjQR/BwITa3U+sqiT+SCZv90ArAN2MDO8CjYe4ec7Rjjq
EtX/26Q0bnEe1cBbbCYGzo1NnmoPKNgikYPIIqm8j5F1cMaCUx3DSUUdjGc23noS
RO+OFPIX4cqYiqxUlyTKUyNRur1/O6Q+Xt6QVAqVJIxUB7cffos/ea2vNFPBCnWV
BT0Sf6+DuutDoQT4eiNwYRaJcSd8cZS+HUj31XSLCJu0lVzJLrphIr38GUDH9cKs
EsXSaj9aLXZg78hHcR6h4jJ4z+TS+nffA6VrpiCj4XYM43PQ6L2UUoTB5zoYwdVy
bvw2ECplXqiYVquoOtA4sRnlYk7LWIWQc6TdLOzptQfqUN2qP7ZC70ka/L3HPREg
PfVpIUelUI09e3JLYu07DePty6AZC0Ekm72caZiBMDXKaDRje63oSaw64SP4P+xb
wPeYPZBzmVwKHv4iFmzmWjFDtMk4hGNJJTVNd0Gt15he8mL6wstZYLHvHyrc2KDO
XqJrZ9MCPzgkoLpXfiln+ixaCOEg3XD0axrrljQXGuHNFMPhZNAg0dl5tYQF84pH
kY8Pr/TXdqwSwkVXdF5HkwFYXXbhEsAY2ZV97ve2MtAeyrRED/JxSUZSELzwdBtE
GycdnSOHMHLRq1BxfE6A/TmXMxxs6975PHw3h1GcHXWyfhNIog8VtO82y1s3Q6cp
VAD16xn69PLVZxH036HJQ1mA3x/qDR1UHxlG/GBgHr+Cc9pD+M+SeDlSpdv4izKa
Zl2rKCTBOoeWKehordyXCSaP82X2aekZ5MlJGNS8avPbAUmx8WNebZK9xehnXwa7
+DZx25cZxMpLVkFIQNtkYUyNY4ihS/c8NNMrI20U6zfu961B7et7ygl3au/KJ7Ra
n4Kl9ryJIwAyuwj4JddvV0EBfQRv6A/jY2vIss5Ga2nEMZPmqbebHseX3525T8BL
62t3lEnEK3pwNLGFSFdPTScdLQpUnDWxEnnte2v5uxGSCIq4i6QggMYeR0q8u5Uw
H9UofbahoFG3R+3WXLbgkSdUeeULYJ4T0MKaawNAuo6km0UGBRK7EgR0NncY1Elo
7LPY+LDTcroVFh9JbtdvC5pUJYK8Yg/o9MrlliQ45b/f/7Hxr4g6D/fW7R5CWlgV
O8bg66qf0Xz6AkEYrfPJkmxQeYtVIxxaq/TzHqmUYpL3sy6o+6eDYCNPE8qDIF1q
/RiTSr5Q7zFq0/Z8+uOkHpJC3aoQmjCVs6jfCd+xZPxtai59aOiCFlZY6U843WUz
bmp8aWdOxVP6OdPOrMODEaqKd8izVAZ5VgHByYygEqOHCl5YSGi6JShZfpieiVL1
g3GdK2QxThgyNSc3nSW686hTItQW8n8OQcTkLw4HWkmuR4ENPLwXvEjw9tEH3tDM
XLCbNui43hYBhdlq4JDn6AsOivG42H5X4whON0xtg50sM8zsZiG05wcmH7MWvPvA
eifxiXFd7HT/GSwM6nQTOnY1w6mbIoGOpBiEn84RadY3w66kSv3sU4f2FCaMKEcK
LrGCA6OOayUr9GDCqLOPmAbI128QOXvy3alkxzhk2LRLmSwxQ+EgGwXukmuwx5Wl
RjslNVN8+9KL21rUM2GC2CtzaNSAd6ShrH1OEbl+BXLVJBHDfKY2tZwCgCOgq/hq
g1vDbwqXgS9rY0nNvt+lfePGmLFJv87yAEdffDNmBart04oxFTOzi20S7ehQFLoC
kBJ6QglwSOSmf4Wh2FYPVEuWXY4V9ge1+v+i5df3qRjQ7iO0ya130guiA44knN+B
9/9xbuUpeUkUBXXBPbPOPC8a5E3/Mgb5FH2zhlftPBoht0wuFBUoTcxlzzxOuy6F
60pC592ljdvdnGGFzLxALlIVNS3iGMQlr9N+lhibxSs5jQjTJU0famVfKjPKhclr
k0my9Q8pHeVRTcw6Mz6fFDsQL1ucsJiRT0A7s6mOCZTPFaV7/F8bcQzhHPqLiSh9
LMNJ7ZWci8cct9Tu17Ybb1QaizpgVII9UH9f7mRsZswJ7xWz/ovINI3coL5ebf8h
uV77XjUs/1z+ljk05dx90Mvv0181QCYBr0bgiH7s6NDwvmA8g1jFX5/xeddcKbjt
Yal5EEGx38KMSJlAP8vQaAM3snHr4iohLNS6Epre4AwRxM9BldeDhlN0qRtgVhOF
rUMyZ0fWhZqeWuGLZE9xWx4I5SjnG00FTSTeUkPN8daw/2VFapTC/xb5522Lr3PE
O692UzqXxzWIW1g5DML0TWZk0FgE7DtbSmqk0aV/r3GtzEhclEaqIeDpsji5ORMX
l37vuzu1NjFLQQJnXriwnqe5ImVKAnWKcObtpsNH/0atI9wcWWtBcTvOppjTugZM
/Vrc1zR+DjzWqOaMZfWafh0oGzbkless/20bLUWsNwvnolAcEL8SyIaa+dPIpm08
j26+MaQcmYeKwRP9sL+VjcT9j3oWbLE0ZRKzA8HHwrlzLX/QmSs5W4JDyTehqOT+
OvyYKZQkn+e9OEwsSXxn2MA4hGuUnDINGse7KTCIiCe5JkjOO9uLR5hWCKFktE1s
u3Fj8/EppI3Gdub2UpKng2d7p/y5avFsfMM3HgKgsZsf5tCz0sXgN2cG7rqKhEAx
CU0IoEC+7PNkIXd4Cp7J76rdtCD/h9TidLjrBQBt1MpNvVo9XXGT6PKfBjRuoGY2
/60caKNOfDJwJAYKz8Z+UeC43VUsGDZHtVPnl/PH3Kp+QleaHNOADDNdLkqQzRBz
9y/bhtfBWmzgzHPUBfcOSiqwdu8vMOIiVeoXlsOqr/7WSDu8JAcrvIc8ylVEbBG4
52Ic709IQP60YJSPFqc4ZYNTa9EzUugWs9Y68V3inZiLG4tLpkTuVAD67y75QNA6
BwtHFmoVl8C2j2XpQCIgMzjN0OI5miO3jGzSXlJLWnvZ238Dq+qZy5tV+5lQBLES
0NobhGbcivm+Zl4u9utqeBAjEtcQD5PHtIMKqrpXMwPN77pdZ5LC7wfWbg9Kc0cx
SmULCyKg7Z1m5YBpqTet+PQH/Xyfpup9S/M77jUhJVOV7/TkXtJ0J+/l2u4w4XvK
akwm/bZCiurSBOPIkquJXADvrqbfF0NmyHNoBOYOfiBkg0R4vLEHrVVUvmHA0qrT
+DhuT+RpMbvGRJyh1JHDXkD6PurJZ5c//8f2/44iq/Dr2QMczVhK+WvW1XhvYbGf
P26SEa4DxNzCqKzToZOpU1WpngD5SK93s7S0pVp/BTVVZwsaQGZfJNZGZ6IA0/PY
b2Y+m6ozuWbvWYaIajwY/ORtwsItc3qYq2UfYfXkZIeT9QykrlhbimFJYP/l2jRa
z41HRjX2sdtdYe5jUenhN5JfQru+N7hISVd4dgcsZ7G9kcAjBv75kRrr9sJXMyq/
1fKtLn+/gGQJR/y48pctcfnK2JbuxxO5CrujlDRAPBkdWD2NCzgxYn5qLPTnJ2K/
xwiQUboLe5JgG21WM39bzP17/R0MnkxndDXqc7kqFVvLhW72r9pZ7Tf/+W1hIxUJ
IytAxyrGvMOR6C3rEPFOpreyKOQDRLPHQPOQENk1XGA1F66GYXq1hQSSIiBK2T+S
JHZK8PA5+sIW1jctb0AHdmqQL6BfIVdr8d5LAxR+Nm9SRHdNTVpbXtibLgn+yNex
ghjdT3DLmOTfNiCfnqKt/8vOnAmvhvwb0nwHL70cT7JYW/EkF2py5fOiY5/5UZ0K
bCKlxK9tGuA4qvYT6SwCdvxEnyznuAS077+y76j6irLsJLEaXmtBvCnjEYIK1lq0
7yAC33C1h0rL6qurosFWUGOI6w9OU7KjUoL12kwVOHlPj8SuoPH70PJKAHLwrMFf
quBJiRxQibk9FN0ZKNbPpKekBvAP8fDjvSwFQBbv8tGddEA8T9kVGKKNN1BTtQ0+
gpibk6Ph7NdatqRPnl7ECXCL+ScHlJYlAfu+/F6bNhTT73R/faaT8PyKIA6llTMh
gpBUNhuGNSzPzGlyk5GTXZPAeUWYwkElgVMqh7CO42jIksDQqr/lrHGJk7eHtBlK
1O0FGCqgRyqdZ+F3QC2zLJ/W6jx/VJoeDcGfHtdNV3ECE5RvEAUORhca4zQ9pr2I
TLXEnm+jB2Rgc/UBS53ro3Zn3Yh4TVVdLqoXhSQoh176Y1RrcmcdKvdvScJ++G7F
8lnJ9chDMW74V6sd4nykXxmeU0hyX0RRoC0lYQMDv4mpNbyFf9owEtMGEgb3ih9U
OE3iP0cuhmWgrLF0/SDSOYe9m/DivvUmadzqaWTF4os14/HVdIZXmMLUwijQOkCC
vkxQ0Goi/i96vPT4Adi4RcWY8q7V2W27oqZLHp3VlBWnwEPxjXzHr/4mXoguou+L
bUwGmgE/NSk956ySomnewAmtM3dCcwXsEBlkRx/T6rSCVoR/a2Ay+Qr5ZQehG6Ul
qlSojzqjwJmZS2O+Xjk1BgzILZ4/dJ2/qkfg5V2PRigcywRK9ADMwF8tIvSiUfIb
w5Z7B8QOJvOnnkfat92A/zTC1RskWsy/QVMcbncb0tjc3ODceVBMdDpSepyOdHw8
xHht07O0NEy4S/rLZqgK4RSY+NzJ3oZtQEgZ7/1ig/QRRcx6TSCsTS2OwCmEW1up
7uegnXUzHlkymHN1Fh/6T468AL2jidu0hM4WpOd2D23SgtWVG/35jZjJ/ihLqaOr
SqBfY2MbiUNangEAWTop+RkdficZsNuA9Nvuod3AJzp/JYqbs9RHX7nXz1AZJJVI
lJm7zdY0s715KEk2/MQ7RtTUkiskOhOx4A/corcGcS8AyuhpeJP5UZRv5s4+/w5l
YmhE850d51zwnyTGbUgEF5momX+EejVt3qNQW2AXX1wIUwLAygh/KLGojGuP+2Sy
Sjq5iSKUKFQO4f1XbXvA5rjf/LzHeo+xoLks1ri2f9soc0rGpU6QWJw+pA+PpAmZ
Mp8YXUMaYIC0cxelXz3zKwEQEvIk2NlWT/WRu52lQ5OEmU0yc0uz7iLD/d4oFZ1m
jNOVWNykTZeceokuEPNuak/hoNWc89pE12vMSyCZmanlTK3DX23anyqS2423kryW
Ej73ouEJSbzm+dNitD6iIXzmDZjInmWw9R4h7J39btp36TA6Xb8EQgbnORSGJ4hv
JONqgsTsIzlwZZzpUDoGzXt69sF3gfcvzr8njdeepkf8i6b8dbQEkVLHjXD2iX9O
a3f6Mq6yUwPCruQBvrpHSfsvNJJjYxusT1BXRhyrA5nfbtXZhaS1mX4T1slluVKh
bIElMkp6JR1dCsID0ToXAlWtzJvsoIgkTrj9n4ZrRWU0dX4k50Hr8w5moRJXnido
m+LMzPC2AYfvA53v4gf6svhrHoJTpIdVqDVxJCrOtdqyPSCLv+Fmgy4RtvK/iJWE
On4M4I31blLDYPF0lASmhT5Wj1YCBRpvuPt0reo66c9tbqs8tMo4VAKdn74/oroR
y86ewZyCWJhHspn4ozwOSlA1zObyAXQvWL4KDy6WYwUxnlyBQhPtkheqaZWUju1x
NxuNyGKKt/NQ1/1Fv+phLPKDRvoQMPBKz2d/JorNXWjusMPVLt7AL/NaiRSYw/f3
HL9Kcn5rUd4qJr8B7Zrq3rsaCNwFtXzguY58k88SY58ARS8l+DJtZAenSBtL0tZU
5tP04Bz31VRXq7446TFYW+TQZhjPCdoQd1NoNWVvioi5q8VkA5x/zsRpfhxQnDp7
HF0UZ+R7KTqbtudjGXPUcjNIAPYvBLYlRjdBvYKVzOslfD2d5JmfHAi15THv1KNF
XEtGSensM9Jjcd85DhQRjvM02jgJW7Qo9ZqD0HCEdl4QAvTzTJhPgfUNsrd/ndh7
OFPIdb6P0RfMxxKD2NSs3CtTGsiQeUmFCoNhA/XnowaTTkBaSF8RovvLgMg1LWWz
hHkrZRE2pzCrPFk00puX3OO1M4DjBROZel2MLRP+hhabEpQxSnPe6jq/f+67CxYa
5sXqulOfee5JnJuH24QhTr4Jjr+ND2Ds/B810JbJ4ZFsTEwjVsbdkqOXpBDde+WE
SoK6U1OYBqbD8gAoRPLlVPy94sWLa3LBbP/mgKo9enJbmi1nXU+usRG1oi39APk1
2JfM+T/28Avy4qL4gTJUq8MEDFVkBFTojdjew7nK9khntNu8Pc7prC0pm9tE+q42
kWgZzPeIU8Lr+Ijpld8zwbMpjoy5zzCEnTNZXJp6/XB9sxX7WPhu6XCvVGgCv7IM
TuiDRkGIcYo9X6cLZDZswvkd46gL2gHumEPc4iQtYrTFmu6OfI0+jqGd7rU7t3lu
+2qZyQMKTUuRh+CtuTRCdmPo71i6XnoQsBu3SW7AIku1q/OywcMeiXLeaxKJQJHi
OhOO7pJbO0SV+91MfC7jWYeLc77UEYySV3JH4xcBG/NNLioZu/XMlTJ9hBruxQmn
hNF4ko+H5g1mOmsfobLUV5lIr5qFhUZBHfwhTxphk0PIbdUokGnHzcBuHr2XvwNY
yMD0ecautfS2xyrsInH0OP5wPBA8quLFzPPP1PaWwNPgtmX+WjzRmf3AbIvXDcA0
x8I7ks6cAe3RxY83LL/eHmfaRAdrCBM2HO222dKAb3CUmB5N65Ax5JAgjgd0ngwV
uhqfcUieBGEPhnZn2NessQsK2isjKagJ5afoZDTNNYN0T8ffcRDVK9h8fm/Cbb+o
Zi5T7NCE5H0jsgJwlwQL4nk76TvVeUenIawmU1D25mvjXW/OPfI1n8GQrRHMFshY
sUvaoASkJI+H02RPz3IEf7f3312yLHNu2U59aTs7amjjr+ICW5qYi4agEesIZ8h2
cyKKdoNQZZDl6oTF04tQZ7LRm+D3KBTA4OjkDkUAoRBT/sHwm47E3bekSOUaz8Zt
lxCWbXk35ttu2wH0Lhl5prtdilQqpHbWrpYX95dGFiN68hVzUBA/S1nqMcmrKTSC
wUw9GIllAhnoo2gLOthYL9lqudmiU9OGt+gLY68I+aZ2GdY7Zabq+FVGLA1KT55J
bwM5cs2/9QS2PNdb+92SVGbJKxSHoOEyUUXRqEitlvKitr6gf7mH0+XT1cpZNJpv
gzWCFJobVdJ+Tty7jLf7y2LSizJmck4n/n24hRi6fqsQtQehuyZoPYjUoqfARImI
giu9KUSQsew3A9CR0Ld9C+FG0bS5Y8rs0iGKL+wxV4XXmAF3hYzBowpl4FVNc40O
ODqG6qTURImMr7grmB2Tq1RNXxbUxrYOfgJVLy4ARpCyG1XPnYfXl/a9K3kBJtWt
JTetC4Nmk0tqKwkRbBe9MPv6YAaYjxXmEF2xVUJa+yrsK6OqG4b47BONiH1r03o2
F/BmLxUiqOD6z6KpnqcCvPr+dZ4RKJsX8C01D6yi45MwRhDrFUtpx9MfJbvK7IKo
nWgEGJMoAVRKk+/apgewu1PyUEo+nVUqrf1jhCyOshcHkXLd3A97TL71swPJ1mch
/1pnMeaZIWddEGByUHSr20K25UN7ctYuTDLivEcPcfOCfQC4gsdE/TgtrV4g63Gk
c21s6Bo6WKarQJ78i+lAy75YFJ/pk84ckHDwNc9p7gs9DKLe3WwE1aD2RRkLRaPv
LZdr2krla73f1NpVNQSeiYK7MWXhTCdGrrtvejtINl7NOT7TdlQEFRa7ih+hva4V
N2eYMaRZJDInrntY1K55ofGcIaAryT6U4MsXcXRRUoHgsl82K385jTwZn2evebZA
NFM39zP/hn3s+xjoEm5ieG5/7sLPi4iV/cWmoJgXEmT+a6rhE6FAw2h6XYT07Jjk
0nCsqbBlt5b6uMr81dbDdISUpbiHIRTaNaZMrThxuVNkFQUMfAOjWNzWztQ8SCpO
l+plMf0WDap560oYJ1dXD6ujcQiNhrMZe1L30jojaVSEcK8KB6EfsbvBuwYztKHu
ZoyI4Nt/ejEb7gDpv5VBio4Xb+KZi/Pcmhhd1ONUxlMQnF0feCE0lXzcSe21bnzj
pp3v8FEcZsylJFDqp0729yDSSlfoRxZ3U4j6FISbsAAmDe+lND/KIGHPgqcFMnnn
0kBnev+PQGLk+eajtg6mkmzMrH7qiBJUxzAeVzuljcAv+bqETR9FfZDXNVOYZyw4
sUM9sXg/4afIZZnGkN2IoOcI8NCnNcmwWbMCgNqXOVjG8imL9lyWThmlcEkqKBpa
AzMsmxLD9Nepio4OdP0B8eecyvApEQSvFh+yZrW7QC5Gf/h0Vob/OlXKbtC8cw8t
b6xAScn/G2OWcZcJUxcAtx6hvsyBitUQX3myJ8sSckn23Vu3lIaVar9uIBG0iSLh
XZwF5D4+UZPCvHo305rXRrgb2xK856SQVIPcuwG5+VnItJPjPU/PTHvjCdu8awy4
yqzvWNHeWj7Z2j0X6hn3qPwsdm9Mf2JE7namBz669CPWDMVRYtuDuIRQaue5BmXg
mL3P+Ey69+MANeF1tSbsmU1WgiPRejr3GB5WwacWyNaa2uuzJGG2WuwzPPtu//O4
zCxcvwtQBpXrM0fcfL6X24kNaIN4xYMlC3vBBdRwDTBwljONkTk76o3cSO3sTc0c
8/x1wJczAZQWvCWBQ2yAI5WN9LZZLqcYqu+lG/ocuQRssb+unXPyYNz20OnUwDIM
KnDORjIbB2KBTMVm4yA2SeopVnJG+jC5F2AtgMCRd52ZCOtRTI9A+wXznB7bQUPB
ZlV/lsz+lfMSLlrM3dxFnQikcuxOurXE8ELLtKjHAYm5CvXnTkI54Dt1+clRmusD
BcIu62cRUSMXeICTcdcqyQu3NrVcVqH60Jg60JcGb/mMLYnKZEtK23hSLYY3eJZ+
OgIK5pknaBZAUdxIGF0D3UZ/HGx6M0V6iAmU2l+hK3XXSxAovrY7vT8UwHoIfm9d
rCrjU3pfXogWduWWEebuR+14dVMeJqLRs0/u/ZQowX164XEa3e9Ux4cw1QcIWMOv
GX7tLFSI45ZZW5oLVT42NkwWZMQrW5tH/3fnredKSfAdV80zF82Iie8XqRdyjLcY
EAsa/RSOlqwIiTQMzrkwxFVQQzDOi9KUiRufjC1xenLxgd6eVqOCkDPNb6bOQeQI
SsrXWOrulKSZi0D+5WxD+8r4WCC77siUPU+xEf3MH7j2u92UBbI7vYFEzEHguA9j
zqfn6TISqsRZs0/+rEJeAphnaV77msRgeLo04uT6zVU+JlztwZh3Y9OeTTBzLPh7
nctdeTTL13MP+mze4/GQ6wqk2e0aPsTWzlJ7Dq4cjytjG2DA8zha76mCkKP9NKok
q2260q73w3eE8766H/Y9cowzh8sVO/1shLyd1LMCn83/kwSimLsKOSeEOqdEthtQ
ajEVOKXikiaO4mu7XSEzMGzZmgpe4Ymd2RHi9pOS+eIf7vHmhSdQmRKB3MchnLXR
s5oFjQd7LNP8g35GaDGHYieVJAfM73SN1sY+hGVlpDexPMFlt1A5uyMCJqkbKc+k
yodEcB9Iwk6QHSrhK8OfYLkgUpAsdb1sSTRovJxXyost7H2ruOa7OaypdsV/AS+V
sEySQRcT41awtrwS9Rh6Sskc6hJqPr1fSH8w3GterEYMw4ZPnTbVA3FLotRatIm6
7jT/isFwtfTskB0ms/m8S+S+4b/NNT4qUgPtTlH7s3zYxZF84qjgCBNXox4JQkq+
9mz/7RsdnmSKT10Z8cKS1po310+bqeF8VpPYdfYZvGiPPFBbokssilRNtBGz6nUH
GFPfy4yTqKe3b7hVMjpsa3epsSBXKHebh6z7Lcez23oZd8cXwC0R7mC/JvCiQsEp
NZpAMlugc7KRvTqJYh7SJ3ZUbeCvfNVwJ70ogx8bYBS0LzzRQxS7CUl0C0pnRHO+
hOP4kO8u5bwweD69j7d5Gg2fkh3st/CORPqv8yagmqLY2QIIJokmtXG9TkseoOWk
u37eDX1fMs6vRqXAdGuxClpWYAPtD1naEJy5/MKeoiiQEsNmidzpqwXL4ip+0++x
zpvLMfmjJp48J3S6Mc4nWvfeDf5LRe7vh6GjZAZTg5YCfUbGMg8mKAyNB2xHoof4
7Imah3XuQqlQzjK5g+KZJew7HcIJj3/+AzroaTAH/mN0fxNaZ0rTJw05u+41mRwo
E+VIlxzdAmLZtoiOjQsRvxyBeP8EKg6rks1Qm3wxZHx2PHkj0EV7QBGkMSitfsyK
B1zpYVXgVVQ+ZWE3Jjo2iSfcN3HAPudiok4PRsXMw/GYLzK1vkShT7j34mMcAo8K
pVO+Y699WBLUOU76CPdZaD1PgXtBA/x2EpcfDgc8lIRnZGe8CNVgACxe4VWxX+Dy
DeToe+pHTTzcCKBlplM3fSYeFtW5uTdAZmBYwVhIltw/VK72QPZyfElTJ52vcrf+
axE2BPKBpAY2+D0J0WbWmvF3Bp+GFMIpSYEN7qX9LjBRt71pUVRPm6Or/biF5993
SN2qEu3qDumtZiVgigC/G1pWS4wG7a6v37dnlP53PGFz0+68nsOWRwIM+R6VH5md
bXvODd5NR85GJNcmFdz8mHg2ISG/NmEK8t5YlX31SdZewULkVZoGqU1qhQTiujKO
sn9+puuGSuONBr4C/QMLlOAbEEr/JZQ44n53Ti9ssVd45MPuzdWs0faChWi+E0E6
VMBG+DEaFsrs/jFGhsjPcAgzH/KYI7l+oAkL2r7YvuFCkHEshDVlU6CwobDiaHOy
3/dTnCLAMxfgXnEch8bvyzUCCRraLqVhY8WYYLIwC91jZ48fMRziFKPybwYasj/M
uAByNY8aqqEXxWwsbhOGWJDCEO2OiYwIxaI1lk64D8Eyg++SpAxXCe65mdnP1khm
U4dFVGFo+MkU1EDQccsOB+cCnaC3SB9GimJB6ADbdXNDtbLwIf0JjESmjUYdnYmQ
i0e36UjKOVyxf2pTWukDxJgbVZEVPKUCVSSKfId6WtukER8nXNTUxLBaVIcxSyfA
idD9awzBUvOx/a16URXEHvSzH9g6+NBtXiSK+4EgsUxoPZWmhllXLU1c2urVc/G/
dWiR5QBKDbLjMRTuhOtXN01sMBkLJoL3DOOiadVtJ/u0Xi+r2a0pZzNnrhCgjxQE
hvteFIX9IIs86hdUadBIRLMO7WUtex9pzpJ0Hcvz5h7RbANAN5DV9p3y+I1Km0wv
ectBAV+EEbXpgazSG8G8+kaHoFTAFCyYBuMm19qP9jh7NBuLTIkg5GUnlFAhltqL
dG1ZVfriiYvI3G2SUc/OLAhll3jMhtBT/ZkC5uthVvj+DkTov3rDb4JZqH0t8iGq
81k54n1uzpNr8tKFdCdXz3kB8PqD89r36sPK/Hy0KRaPcyYA9nKujQKf+nobeSr+
U/nb+grbpfa1VnDxuoW2wvYcwpdloAyO6uJtoywWFnYg0gqJdSxMiko0YsM3OjJS
2PVmUPt/HCR1Dqll0qR06KNqcreZS+tOCXLNZlEKSfTaErGYZE8qZA3M9OPidjQu
9YNzEqtH9P1vTaBY9Dp67BABSxv/N4HKkTmdwZyl3vaLqxeVV65ixyytcDJSPyo9
zywAn95lFIURUECazLxzCw/r+MCaitLW7e9nWRIA6dzLLtCWy/mctviz0mfmCCJ8
STWp/EekECe8mjMBhcwvMGr9O6b9w4sQ/58U/ogHq9fky4nXqF+LypO6RHTiSxWH
TJfO3+Bo/XAavMRD0+rKd6jbqJlURKy5h8W/ydpGGFzNZKBaEHKgp/QdxMbQl9ie
hd5CcwLaZwhBYSuzVcFK0RcntTBiGefNcz1P7C5yfRbB2Q3jKZZJBvZS2pluLCj0
oYY/y/3nE08Bb+paMDsDajK8ei/AJE1xYC2CSIRdGyT76blDW9JjTvZ1qt8BZXMD
YLo7atV9pZHzJFpx5z5vJ56nraJhPlDpEaEIJePGK5TI/x/fyB1pZuL2IHmI8hPA
yceCRtIGllUH1vgQ8x7jdPOYyPB9xOYsWc14t5WmMbCeA3epGaTuO024xiQIQ/2e
xS33lcmN84gIp7UlBQALU76X4L9VkGchTm1/10E3TOqXE9mmqPC0Q95Amg5Rhlld
oB8GJbq4xLHo1C+uuUC2NXdi6LLUIl5iGTNykTnOSEH7X12I/05fbCZHa4PrbKNr
bpr+1GKoznRaFJInmN+8eXdf9Fje5isQjI9CGxwRkXl7q41PKc2xySWFrZRB1sVs
61dGNuMjR3mnDkTgKO3+Avh0a1fd7/K19A2u/7a5t6lncbSkXnm1VSnqZ2zVeFhN
xKYv6MhWAfaSkDadVXqGonieuBFekGPr3tKCkAzYes3DKxWhmXnCt5TjpCykJES3
xq1SFGm2BJ6p38muakZaXbTjkucv6mi9TqqdDXkxbXw6JgoMa8uWZcC8OMH4tryd
4zlLV3JHCEmnCh6i4BPvwc8VSAyCkPqKNFX2JxhiHl+yqq2miYHU4zj5aRb/SraX
xCcszqInWDirm0Dm+XntNu8hVac3iXOaWt3hZNQP+5524qL4krjLOf/nENnwUI2e
A95tsqFuI/JfF2QtGcptle5kzIPSo+DQEVomXqvuMDI+ISmtYMuMazPlnSuaJ0jB
6rpcQECX4kuF/7hF2QAL5HZ4RxmUUvnzBrmB60AH0tkISr4k59vTjWeqgh2E8ukN
tG01sBtsfcXB5Rv733XrnZBEc5yO6wBPPW6ybgKYgfcVPDGSh+pgZFHKo4JQLAzo
Ob4ZclTxFxlwkp91SpfPIuv7Tkxn8kPdM8/60XeQaz8jcLjRawqXHy4BcV8jkOY6
N8KiYneo+QiHMRtjn5rBEYeVOB6AffOtnU/kSABIc6GCUp4IfsBy9AM3Dnzrc84A
L8popJvufVUeaFFxK/MwpCB6cCtRv4AVJoqszxkSpxB++2ac7MEmEuB0A2otYwjR
Z5RBCj0fI6SaFWkRwxg8nFLjll9ORjDk43yG98oWILNddEV9o3XJ+1WRvbJ3fovw
opUHuS3filjSN4U8CD9D8pfZXWemRziCXidVwFTbvWB2fuyql80tn7zwekSKXu1d
tk+0KEkqgjL9ZlvmPtCYaIf8OREbvjy+lUvNDy06+gM6ZetHRmt/uXzcYPYEOQmz
GvjBe4o6ZsctMJelEjSS/pxXngWXWMCNl6XZgORN/j8CmJzCxoUpGlsCsdsUgY/m
DDoQjRLi2bmH9T6Eq+vf4slC5SgZ7hQ2q0MCv+Xj9D4h49d1CfAYu8e9Fv0IcNKm
8ftL6f/BfxCLX44U8NIp4z9h+dK09Vfia1bT7VwwTOFu0tYj/fOYW+hs440cFfvC
ShID6lFZ4Pu/fZxJNhwHkSGOsSab2Cbig6BNaeCxZ8+XvC4+rg6NeyNHjC2NSRVC
/5p4xd6JoTPyW7con6kVB3JcPY050/oJax7aOe94lR3ZJyNd7t4CRXXyVFkf0VSn
9fWRKPL72CJUegx/lSo4+cnfvwGsXXEx15tpCSAgRUMlZVZ+cp9E+rqx81GZmlJk
wSxdr5Ez63EJvpxr6vl00tYSpPItZmwkMT1i92k1kZz80VwrXhsRNAAowboeVrS+
CNOKTZza2kQBgFGcwTZFCN437sBlDs+DAw9n6tppKe2+47OH0dyX5prEDhznrtD6
FWF/Zs8Jd4f+ynK0hLM7NjX82aeXRhy6P7Q1UYcA8/ShG1rlGfhqQYJKa/mi/vOx
Y6i3XJILSYhO6ENIAjVjj1zQJskfj3dNqIPcfU8AuZ6yEtFkvCxfstojpZfjJBMp
He1lzhQPltDyzMI9pwIPFpKX3ia29HqVI90q7+vuxIJwjzuUXuVLNUaTNaLJPISl
6DIvk/qYpN+leltpM8UWcqVHGmF27mHYzym0SRAdwiDkgR/XH9vQsyUiYgGIjJIj
X+KqDDWZBJi/kc858pnpvPPEulDo08Jfd8iTZ1aHuG9eeGYcDn/CyRK5v5VSn6QT
fRNp0g+IkXP0/Rl3+AIAMY1HSD2XzTsDIb82CIg1nRqUjJ86/HEHCyC625FI6UfH
Y4/90SM17/Kfi070oRWm/Gej0+Iz4wug/4g2NaB1GeQ4BmjAJYastXf+LW2/y9YE
S3Yvkssfg8rvaf0jcRLNcZ6TtS7y8AzIVsLaKHVnoaDzg5YKAPqCdfjIloFV69oG
gAqxZHsamHSLjthJft2Cmxa8sV8iMHiDgHJIuNMCRRi6jeODSSqoJ7FyeUHb+5z3
bqn/5IK3ZUcRyIUwinzhVbOcRZeItGxl19bj3OgliJYnbnwSKUxT0H20uhdvQY/y
SsnvfBGEfXWMSH0iT+6mIZp+cvqOgPsuBuduv++xwgmrAPXGfZSXJNx3JkpXaxGr
sowD5wpu0W4KzE/oAw5GTQ7nRePa3AhIZZoZS29PuM9Eyeg1fGdLHMh+00OeUdNS
Fo6jQZBLIB1XV/rr4/xOrY5nudOXlrTOD/dZi1lN+m9iK/lxkywCK2KyXbTVlJSS
NN1CaME7k5z2nfj3VPjANkMI9uPc7woRXcJp1RK4e6vf1NRW3+nABWPvcQDbuRxQ
FqZKkI+ZbJT+9c/D7rOB5f93un07dfpnaEM04A9DLVEtYx948vcrr4lHDPhMWUrG
X3WfEbvyR0jZdxDZZ28tiFJKXY0OPzh95NFq0Ov4YONtlAIUBUunRB6y7d/FyZqG
ZsAoVYBZsd6NN9gXHinkU+8fqKz0Tm3ZGuykD36iMOFrusnAzFbaPZOg5/0n2QLc
kejP6gWubeAyZNrvN8FjVpb3kRT6+vH6sOlv4QATAV9RWgRMwrh6xtDxzTJNH5Tl
QLLAtLr5RE3JCH+lHpxGRKcAdx2+kb5IpnbZOK7FFH66+JHJTqTc5SKt0JvMcady
DliqtQxuwfA4/B+PVL8EIB7rPoh3Jw4d0ZkLTsqtu9ADhcGp7Qandm8i+K1obZqC
lqNyH/s+2UShBja/3Ab3z8P5yCXIPLtSYj6pBH31dM+Bop5NPZl5ujDLXQiK5DOF
GtiptHwnNXUDjzfxSpMR0dPCirhxsliFiLproUQ41x6kEbFLZ9WcpD6+01q+wk1t
l61h0lpLWj/xlOo7ME4hf9hCk2FUnMFW/xFt1yGgZu5YAyr+J6D5vypCtjbjzQej
72w1tLLrAySQKGzL4AWq2bAL0sy5PgJ9NpVq/FDyi5ULRwt9fanA1tdI/UKl3MY2
bjKI6ymZT5/0W7wV+APBtUk7X6VsFDZtWSPlskO7eVkVyLKvuCNLbz09ItHFeyCC
peNQSQwZ98h16PXvSzIPz/q44/XGed0+okWqHrl0KcqyjNtoU3K0gtymKMEtZXkB
y7WyuKMiGWePEiQlGfATbLgRCu71rZtugim9+XWtQH2RsSlBUBxxTreGbIePHO1e
kKM/TCQR9DteIGZJ0WLRfcjTcyc2jn375hBA4koKCGpw9PX9oSDRiOsoeqXiWEAu
osRj9wplhvON/7kG3T6CdpiQbz1Mot8BSh4W3jZ/Y17gJ6k/oGTvjaUB1WktwTrd
5CKZR0t9li+EScxCrHlMJP2une3RAExka/j2bDYgc1W9qltWNBAr4HA0y72zybVn
W3klnfNEd6fyG2+sZRZ8o9Qijwd0fhE5flO8mCmwQmX2qnxYa4Q7bmfURP9w6sAB
JQVc1egXmqTiso8ZdYvqgHM4oCRaEtiFIi4QjxAMvCT3zQbOcvPEOxeWac5pEMld
5OcluVAScAvCr5VJrsaz4hHneroQd1jnAWX5ec3jpIZDC4wFa3Lix0RAG5f6AICS
rG+0SpnD3UtVMTAe4kcYGJungL/rLQLxrnvxXhb0mvewsY89wgOw5J4X+pEOApXH
ZtRaeDpr6yGd+MDT7rtP1CSdhVMr3kDHz6qg6m0nqemATZh2hWlCq7KswJuGDECE
T900SSxJGv/xJlcLeRVXcB7MOCkFT48wLmqUUNGq/DJn8K8Fz6/hMR37jP66gZr+
CEh0XCMM1NCXn+Aa+D7RabwV2NSGY5tQ1vj4DD4gOljneJz7r2iwZyrOKN7okiwe
uBdgE/6Y3mflWzcXm5AXUjEK4ZzG0vHtbZPyHSrVYoebYOA6/aH20PTLRWeKjCZQ
04tLWIceAnAQivTmA449oCQUVxewIETDvrT3KBb+sBJVSbDCLgUJTH4otYPPJxnl
MyxvSyq840zi+wspYsJkfQHXaQkAx3Hb818NdG4nvm0T281TsTbbS/ociaHfqoJr
61rzLlkN+2z6pSUPioiyYRrSi9VP1ltMJxMVyXqpHbcKphdk+UbuCPojRYktoVum
mLAHzIhD3XPx0UsA8jNKOJvTX1mqozHDXs+i4FIR3WdoMdGq2ar5d8FouhAe+6lb
sVS0+dkzvSN6DMDc9UNFV7tinVnOBAZwgzVFMnrmJd5N/zxRxAyA3JNw2Mxw+SkP
cQXVgh+cMiOWnApUCr39hZELPYGkuLqBYJ3Q7yndhpAedPdzVTbUh5Jjd/vUETHi
FHsXhuQhDCMtVTENSLaNu9+gkuocWcx8AcRwKuSkTSt9lEnox96jJ6C0iCN+YbGB
Y7U2BBIOsesP39JIOe+FThzBXCBRnRmcaCUWxqxXGYH0A/tSdtJHoabrFveKfvob
G8tioGPed/j/idV35mXLU1lXJdr5wxRdkedyyA38BNXoIclP5H2CEXYXeZIwo/CM
BBxCWXqWawVFPV19Cbnb7td1KLfuWEfhnUrCOeF2VALBFKL3/cjoybOh5FkDB0lU
Lm0Q76jSGK/4FqAK2GENeAaSiUST4QwzMAcyw11ms3dp1fOZpO9ObGz3DqfCGAEy
VvM88FfYGB5tmbIdVLimTufUpzALLjgQUAmcHervT09omnWLMVx6j5TRx22O7coY
6oDRzhj3vC3tcys0yEqOALYfgLmB2DkdtLxQgW4lM9lSY1P19h4A1kRvjkcpnshn
URJOfzfxu5SGECM81PHbiCxtgsSNlUPsXdMYSWta9LJhJNTC0Tv6HBdVSOSnaXC5
m8g7pGAhPpuOzzeE6hsTLrMkmowH/ULhYY0F5NrQGa6HuOSWpPyLKG4FlhSa1M/K
Q3ApqFBY5P5ARiIvEk8CpDZdjPB6k4FFrGJnSCTu92cuxw5cPLXXQ4Gq7+qzlW6v
seC88HsgUT85G/Dm+xWfhrkuY7EJsxpjh5t9ME/UPJ055g30uAWpoYteLk1BoqHG
b5/41cXUQFasQ7kA35fpXyNa84iVqeYbcuWGTDC7QuPzODtvb+J3Gm+iCW3eYfH2
k0B3wHc44cLyEoR7sOrsO7j946T0b/vh77Nu2hm4hxFJy3bu1hpZDKo2nrc7Nc/i
FrHONcGqk+yjbIHnX6AJHC1W9WekjjhTCTd+ru4/zHGRimfEazN1CTjzbuWB0xLY
WJ/9N7Zw1VCsOsBsRcxio/ipIFI7gZRRNzPPv1XLD3JltNUp5xtN5R/7dolYI8l3
htcSaqwYM85vN0XVgQOrRs5mQgWyWVnhGDOJugZYpT57o5t9FqH2Xxpm+YPz+XRX
DmmWnaEkBO0iX3EokD30QcD+6DNIQQNwFb7dbus6PoIdjJYm7aSEFnsVlV4AUOj8
h0R09ET5qS1+dBagVJ11zUyOZQztuqtKiF9QizbVhOe36wLFASiWp6NxTlwbdBTk
WOiTElwEgYqRP8adxtDUWtokceuewqgQEsJ7YhiQE1c1NB96+ml3W+lsltHfFCj1
FqEy0b/+HF02hLD4oQLDWsdvb77uz85QPFkKR8n7uIm7ZHDt7r6yrIGRer31sJeL
yx98NDj9teA9qMKsCoN7fMaPI2j8lS0snw6FOvtOZSEB2MXE+tQCQaFxwLk0/4WT
rLE9w7RDksUVjLGEFQ+X1j3aRz6VIClBt64LwSyJ1eesbAddQNrE+Kst32nCkuV6
Clqa8jTilzeL0Q214HNmWayHQNV6HA1l0jKmE8Rv/gdw+l7S/ka73Pl70Imd741g
yFeiJ4Y2bqhcRwh/VmJSKfLpxz7jddscgAqu98p0mLCLPcbcXF9UrB4CoIX0WOiF
2zhkBMpusAte86lqu3yM+p01WzNu3ssdr6LtPJj3aQgUK+NrH/Oq3ujq32NvVcIM
Mu+zvvOrfavNPirv7ZGvM9LHrYtW7Ndqt9a6sPYECtJ5dBM+wSGxdC5iviiAEZjS
mPBo98nmVtZtc1sWDZM/o9mKZ3guUukU5d586AsBj5ANubMEQYAQNbDP8DGEX7KQ
gtLpZDTCbX4gU48UZvv+gI+RK64LXqQUibs6soYRxJ9YHcDttG7IHIa1IcR/7ROt
Yl6o4dVFxAFMXaGmC7g5tDHCtTjcjwjvmhSComLVSusQuNlVUJiNQ14L6znH13dA
pHeOPjV2U7ys13AAdbYMZyrbRvTkQB+xPNJRUwWH2AFsKtluHWLZnDGpqxBPjFTM
mqsJIYxb+DwlKE0WSHOV2cU0hZqyyskuGIKeGQdlISL/laO2C9UnidAjaByi5NDB
du5rrHzoAXk4yLrn3rm7deZODE06qfVqzac+gZNax/g4QheZIAsYTPrBEkReOVjg
1qLwL/Vh4PpdP497eRGEpQQpGJ2ya0iOzGEZdjmJuZX9GYV+kDv4EJeQzp3X8l3j
3FLBCLPjxBdNTx+iIFFwI60v2Goegk//MzHHu3yXvRPIk465mZjG5/W3j6EnifP0
btmGErwwphkxDodo0gx31CWGkKdUWOLGKCkKuXMy9FC3827bR4MrSXO1KP7Beh/g
DkPqpzh8BpdqVBBCnWiWKubvHSmhUocadJOaolWCszFfv7l4GJMkuNl9BlmsPAwF
uuy8uxuMzcqZc/wxrn4quWN7G/u9l0J7P9UH2DG5RFXYwyVoCPOsJwYnnbNO4EyO
7ngOMsnH/czSbaxuTu92XVf+ky+s2EKKw7dJjehtWCbtjUIDz5MfKzGihHI9z0Uo
v0L3nbRf2Totd2uSJ4mmexUfreSA8QmTnk45yuirfNZOvGtTDTVosYWE5lrNvShB
98M4IjGcU0shPEe47EnQocH8V23aiaib3YlS5xkHab5HPOrCqgDo0C2kznnsvqr9
BwvvYxoGg2Etbl93APkpxcx1PLwjd3YZL3daT1F0TsPczgUxx8Br9DRlVz4qTgdu
yJVQUa+jkr6LfTlnaC3DqQTzb8rpK0e+xF8tgDng4FSXM/s3ehbg8wCXy2NzIvoh
H5ACkYjaIbp4Z891xi7BgQSscrG0sDSsCod0SNuh3mLy54erYsEuIh3LAA5osiNb
u2VnRgO0YqsY1XEM8Ye1BJpedePTZk6d+gTnvfPgfg3tNUI55et2Xlgf+4dlULgR
KwgPW4O9c4aWBivTwySwWMYjPX5Zv67Oqd8xtf5+SJQqT0zRsHZUoXZyVT6Vq5qX
DxjWNqQePHOcAzSlTKxdDtZZOt4O4OcAf15a2gh81mjdgzqC/Pa4zJ6MHNO+gzRZ
PfQviw3WqU3gQEXcCvBDHib2Qkl8v5LBicLN/TgOTwtYWEpOjdGR/eFp7uBzzPW9
KsWpwRLDV6hG24x/T4yvno2PgN9fI2ibPijpt3KOt58LmIGymTN3NvGLkKrJjpbX
FB0OKFeS3/Ghb5NcIQYiYjHJhR/Ct9rP/B2+2mRHmWwiS+drnPQ2F7e08Y/hKiKG
FiDgJege5pjum9B/npjdFsGphdh7aqVnnhI5qq1AIrkdZmJTxUaVw0ShW8fZN8lq
WdknoyRjSHBZzjVHIpq5LoDmchek1UXR5SxBRrNLvqder0cSei5LwYFU+aZ6YoYe
I8Jk/sbBxKgBe3dVw23cuWjZhpavzxwfWjOiR7ZfbR3doBMf6Hx+tgl2Ixtb4wpN
kXQzKevw32bDEVhn7JIHIeoO5Yt1XZjr3JJKEQhW5TRhwQi0CKRTtvaMq7NMZTMB
FQAIE/NLcZY2zNLOxxjHtVHq4Qs+9Dw6w+fRUCKoufWzHbxPwxbfM5TgQXiu5Ldr
kx7iG+t9K/BuEvVB+yAKK8oE5qvMx2YcsiguNN91Wyu6t1bVGwxGxSa7llHy3y5A
MUjHZgQeBbm1///lcAKg/8JzwVALh+FirVnnBPP7Q5555FUeRSss+LrQC3Sr8v8G
VOL6Is3utQLv9Q43NKDnE8nQqfRIvK/J11TCGCPDHES3jaG5Cv6xpDBExalfdeOE
FdJDpM+NILvMrKzJVpzGpa23ibnDoX0aWgenaqFv7nG8I/u7BZJL1coPxYmNDpA2
Q4W6VeX/PBmXc6Wv0nnPzOkdi0li9mjemRG6dM6xK/c1XOt5UqAD6BDxOUXkoKwQ
RpxNJrHhnRSErdzQt/5/b0jfRuD8XhxNXJM2ZWSVc105q2q24kApzFqiprQIBuRs
6bc1HGHfK9a9Dv/JDKXWXbV+w8a9lI3eemHGLjDHFuVh9lj6J6n0o+1ceV2R1tzV
VkaXvDEXVvqoUJy/vv8wrQWty+wnJUMqOtuEe7fCUq+4E/DJsDPgV0+lOWNL8RH0
TppEnF0pLk6oRZKR/NpuKhHY3H33fYD6QbeCiDEWQmvTbPbjiDtywctTyJ86CofA
IS9X0wLDh6SAXuE9mNzPNtV79DvPpE2SDlkvVcu4K3OZ8u6yKrK20QNk08lM7xbV
mU5IGRqy3y2Kxxih8QE8IJI2bdqXvFp7JsRpmsf1JegvXiNMsh8aGAEVqdhBpXEq
kaN8ZG24HE3WnMv0do6tI2NK7wQ6Jby96QOzGABtEUIh5C+0n10g2ifWksnnCt+E
wzzjMoUHMr0PCA0FOsTIHS31OJp9yyKcsH67Fk9v14L5MPG25TLoyqoeXQaooK6s
6njKukYdRGLU1prDGCJGTKDAjkN1f8+4kKAFMaRKLTvdF16RQNdFeidjBcJasKRb
Dva6J3bfBmx2RMwz7ppzcn7IDmIRGpRro52FYN2Azl9kEDA+tAUrNc2lyyA3Fd9B
guErWYC+ZmgLwju7peFR709s1X8QytKWwd9mmUYiHQVzN2JeIeb0Dzq6Vkw6XFLe
FqCX3+l5f55EpsCPCeOKrMCquZQZ9Dq+pIAgSWr9cwpog1smj/u13LrQfOkXgTuq
vmW5FY1sDEJkPVHEWp50qCRBveG6SU0n1lLNkMOnpX1UuIn81UbM8J2Uy20zBzUR
5MF4O03SZFrD//O5GY7F7M/SUMqt8sNCImJRr3Xu8zOy2TaWCuhuTm5EQ91S7IR+
pC9M7CjYkLc71h9KQIwihldtdSuIz60VpiPlYRHfatonl8CT3qVJgDHRf+G90raS
brF1ptpJ3l3Bp9oOCVwqiJUi9OU5erMjVzr7j1ebgDpBdTELHe/4Hh7QPPQMsQMq
aTuSMypVUFsvaoosrtZhAXeyAVciMkUR5s0Z2KEQ82oQ27qUhfjizlTiyKjk3XCk
kNb6bcNi6H3oJcDAI9O/zR47qbABIlVcR9kMaqIRelZP4YjyfmlANTl8+fiKz6nb
4C135OKh72VoZOme2qoTFAaOOzMrHFmbsvbrZ80PbGwCbAjeDDmcHJgGT/2dRCcp
Xa2FqyIskhuaBwrRu9AKyoA/TmRm08MzRGxrnVSqfsd834poKXswRJYjykmQk379
kRfefxqhUqPq/uwCAT13sn5wdDy2G7RM2/t/K1Mua+tdKbg60Mj2YghIVsiQhQyT
dqAmiL81kxLcJfFxJjkS6mi/ILcPXBQQ6IwsHvw1hw4ozcqEMdGJxPPBUw9gYwBH
lzSrRzS6DyRAsjPqgMfky0zj7/ucH22zjVimOtoTNR7Ef10XDY4DZBpN8dKB3BCa
b0H+IXuFVRdc6laOSoOy6JHW+WOrSxKwOsQw/J+pkRoAQBLg2/jeg5Kz2qko9qJA
mSc34NxFlzXhDj6cafo4dm0FPF1H+ECmut3TjUAw87+kK5/g7nv4Xu674e3j/dPd
UYndZbndv7lPx60tLVgiBxBRglEWdektXvpvuD/9YzwMAHFaAuo05sD0Gy5VO/7r
Rsvo40YNZhoqneDouV+2QHPPpPtByhjaL1kMJUqXLjXQ8B8ynSEf6s8gv1MV45IM
BIrwa3su4F84rVI3GxbpcdYWCfcwtKi0TRFDDOKG9cC0JAkT5U1dEdIz7ubwtsIk
2CQ2jDBpcHKmTEwMIsN/hT51lAWvKI5PG8mGtufXBVqBng2k84oKjNBMyLKeFwuh
NbnFGvueNtoG3UxtUqHjBW4F8jGbTt3GpT+O6YkngMP0sR4sFlWuT0L/9HPlKwVe
IJ80gHSvqMMnxjKowmcG1CjORMeqXDLIJqUUM8C+VYBykpP9siqt1ZWGp3hOpYrM
jhOMPYOgPI8L3PQZ7OroZKz/vT3gghVOCRd9DLxf9hdnMVRieJj/spV6AAC1tS82
G4BUzu5oBZxyGSL08Q1q89AOUtxOi+IziBu3r3Kf5fGROnIBbe/JxQrhYsehIxrj
pre09GpqIjtm147TvZIZGcxT8vrcafDo4CSagxltLWGtRsAEIoWouIjOSC+dN9Oq
v7kkmvBe7ishDar5S5c2KY8hnlCQ9NkjJF666M6sebg+PSXjiOAZc7m1zdDmwD4T
lUBk9FikxFhRtqDYbiqAUijG3GtszvatU+v0QLatvmXvbWjTswppJpuz9403b/lP
efIDZxfJfr/1ZXd7F+lJbUJ/HnuNmAKMcnwfZ2Kg4OX+PGsaFAGKJwvtt6LFL60H
33hFmJ9MjKgOvBRdt/Y4WT6G2ISKYvgv1kC1/ArTjS/nlFwx+KlkQ7fGSwHwbinF
gwdRt/XLBT1CNLFSUM3/zoY6zL1o4x9cfA5k0OApK/J2hQ41inKPRk2/uqPjJ1ZY
R7GPFfxKDVbfA2VjJWKASlU5OvHl6U3OnCQSGPEovqc1BIVWEwEqS28T63x/U39g
+dTnU8Pzyt7zCC1m8JTZ+LWGklyFghtY7qStGNXRk6tzB1zRBpg8v2HxlQdDuqjC
AHJFxs8kfhgjUFxaWpPAuu+IdSRSex3lXJmuohyGiszTK2kg6ksla6aHI02iEtSf
j2OKx96+ZCEgCLkdnzwPHu1Swu5hVDewy5WjzTBMZ1sNw48d8W734OrPePUKUFcg
HlcjDU9jyH/bUDlGj8PO2APEDYmfb3XyGr/Mmyp0wLczhGxzYV0eUpdmgKFyiXRn
saysPbkNXOWR3asg1dBDdYpa9DvUHbhIjjEhhwOr4tuPhHqanKYeE086AH7KxdCV
2NHBzOIRLUd9Fsk5rNNSt8Rq+ZFsu/IA/2s/HO6gsGT97gpFROZ186YnYwrG+Asn
j4IWLtM8ash8hfuXbQrqyONQdVGpGG3z7/LqCaGcJ18qroAG+Kx0LA3kyNu2ilYm
mrir15QOvQLk5Dr9lXAMjV295OVhDm4b+olB33QbANdnNr01D7x1qcKQkUH1tkHu
LyWtPypMaUphVBLd5R8FK8WmeDI17nnUFFlU35skvMUprF41ppIiPQBQwl4Etwmh
x+cG3GfZ/mhD3e1cXdRjgacd6cl8fFfotEjxRk0VEvRJoCX+cDD+QXX0Sh93V6Xr
7Ng0fFlt1vTkaLZGi8MZKXtxFjpXuqX3HmAo3iRT0RYW9D110Z3jgmOD1aID3FlN
M8+Me2ZlFxZLiAWl7/mjqsz5HHp9GwNE/sOb4uo+q1zpZ4y8FLBce/ylUVNRUbHi
M2CD6pJihXB50/HMgAc4DTaa+6v4CKHnQBDxWivj5UgbhO9VFIWS1pC1TMxgoE58
EfY+kRalbqlw/Emcd26RwtTeimVSw5Bri37sNT8bOlFEYcCEYiKmhKJEmrQGXlEm
ewkk4VBEzID9Xrkbsqedrc61lE2C+64J2rCSC4WLREtRXk4O45o0fRoRs2NoldvZ
uT2STN6uX5M9peiddiwT64/YiUdVNCab6XtpkSemJ0oib/3EHXRhQf9N98CIlW9h
JQ7Nhsvcss45Kozpze8jLwqbXl8bO1MPHa0UNEYHuvbuaHv9GEmQfLcMDiTJa5Ig
xE9eqXbzsYQ/YQ3SWLLJVv+i3C4p43mWC++UfxuJ3FTIaV2smKk34ibzpXlGxWgG
m4jAcI32kXF0M0gNhBj98ZPKi5+yV3HHWrny7rdipcM3zx9AHpQOi+OLbS5uvGL5
L2Br2Q5DATaMWO+ZUnI6JWmMDlfvXg1WaXgXea4ObrAxBQVPN8V0RhLMOjcyBQXd
CJT2GKDClk2gGgey/xTt4UeURdcSTYHnpX6AIO3zMLEBSdnMCpcyGrd+0e+LsY0i
FHhT2j3KJuvn4xi4OU9G2wXAZM5d4i6prTAC971q75OWfW0h/L3hJVC8xYmsqUeN
lO8Jc/5R2a7tOS58jCgjlaBPskNFSVbgkxiL0xwyW67EGF7bFuRUtszEoCfvRtDL
1TjGo4PTLz/b4X9JxDYitYAePg7M7dODuH/Dxj4qnPO2CCCT8yXUvL7O/G97/sVI
XVZCfvsIE92soe9qr3NCX/FdChnvUgcDKWASL+iI8yj9vHxe9QLJQ3NtrdaCgBhu
9nYlFiHSnAf+OKFkAgjcV4de4/ArzPBfC++y4SJEAxtFuSTse6GfDna7Dsok4snP
Qh86sE628qseo8pwWgRfySExoAVhKAzDROVYESuN6XvkHOWN/MpeX+sCjFlk6pkP
UUv20ZAl7uZBs+ENdpL5vWVnO4+XOoB85MoWiPw/R9D2yUYhoKOM7iJt1UmW+XWs
noTiWE7sDLgqFcQgrD303LN6btCtCqEsigJoJPcJoQPYFFH93yYJAM/WnJUbpipZ
aW4iINnhcSOPz0aOxBAaWLo3Kht2hioSEJEAKxeSCxUwFrqfgfjg4kvqDOO7qD8S
fbemS8L2oE9xZdBOevCk8scSMHJSKb3rX8ogniiUzAoUfb0YfoKx6Lekkd7pvPmb
HLGbAk0muRNH9mbMnQEz19vodyFO+2OGsO4ygPF1EqG4EXU82jPIkSCalf8Rf6RV
IU2UiZCUOZ1QDX7lHOXoMOBsGT3+2cc9MVf5eSSYPpexZoItaw7D/2RRAieFNnyz
GV3ck6VUBeqg6BRhONEA6Zpe3uc/Ddn7oXmYDFv+Imy8dF5JthDuzspxP1kbqOU4
rN+9XalUb6YYWOBrLz544pCZMA/M4k1KcQB+gcX3zL9blKy0NBsv8ftehFsLui47
hQ2wugc23f9TKhx2/M1AY3oW/158gna5ooF8Sp4/CwfwDMl+pHyiwpWfm8y4Yceq
sSpnj/myZ2x6ueTl8goLcvKlPeEkv478UqfTSZh+HoJv+oANVfZwdh4xguEeDnmq
uphDZGYXV+q7x3Fhuha3n/NgyY+YnQXeTecOXZZdcgJEn4x7Mq2NXHgchoup6qxH
X5y8yOfjhtLue+y6VeTrBu84j4vMB5I4RsaygKxqqJIxGLSc5SH8qqLeXGnXApls
hRHI7U1FU5Vnux6zsKNfJAuJ4RPRClqjPi8PdU1RYs/vaJmW+mNd4TDYTjTeUAD7
MtnJxe2ZhR9qJyi0rRr0X4+jBdmiWMdq6fk5xJkNRDkvNmN1m2+k4qthiESJvA4t
T3WzTYd5ZGQ7CnpjVBZtbIpJQgkDQ2xwATHa4mkxC78FzS1nSoctYaPeBXyN7+hm
31ud0NgHFydJqMla/Qqu6mGY/0D+mXxd0lkQjDfktZSoLPHNUtNoqXb1WDJKcYUS
RwJLbFLeNMtQz/bLnOae0rxTTswQHp72lUsH15HCFZi7U2+7DqmL8MH3j4b2/q/q
okTk7mBNr7DYKLKDyB82dZ2WdNELE6YO4n4ZtX4ZQQ+ICwf/WdBC/id8EDgfLrdO
m76fmjGJxF7D5RoNec63UQm+AFrmndF0S18rrd/7svRl5CDNwc1S4PS4aOtNpoT1
KU/zPcqLQT0srKgiXu6TDyqU9oxtd9dxFI7obJnABP6NU689eQ2iPE4jYRA4Phi7
a9DecRUAtJpkvKsroPN3OR/RducElt42ir3My6l38qpiWH0TRJAvj0bVazc2vTBX
X6wnTrm2EpDCbSVWJSMtx8zcaD+N+bR8YevJXgNRE+vgqNAK0gPMl5aFbKJ0iElO
Q6nPyZG4GvAmoOjvcbnPFib196s6954Wk9dRv5PtGsUscIk/OI4SxAzn9WNl8LO5
9Z3iAoM18wlfdYp5xJbSO6AksxVniD8aMndxvhFTllREhMxu3BJktFpgrqPOmRqv
3fd18AAYaicJpVpvyAmqQ1/h2EjjJrYyaWKeYj3CkJmrt61xkeVebujewLggFY/O
E55vrxTOOHeWDbuXr78afG9BK9PO0QCr6jr1aqDwARJ3zrk1fL4UQcpzbF37Ay5C
wNJeEL5vepSOT5nz7Ia7tvFJ+BzHQ39Hm8JpVOX8/jvh/FbgMMtTXeevtVBuXwmz
6Im1wa5lWqtaOPUpDkcUkZbOnUbqddljmK8S1fMI2Qp6o92FF5bU1YFkfRrLmet8
cJcCuc2U6PUWShCcfoMgYzUwO7qdYFk4IpsO80m7+KXoWoKddTRxxTqeHgiSlb+T
+3F+IYhBoxi3QfkGaMKkSisHT/gkXdWoAjyor49aqPAOe44OBtFcJsbcjFmvBSjn
M+fy0HNAb+oMER6Fp3znVZCjou0gWAJ3Frh4zEA0y4ZLRWQJzwpthj2nc0DoROyw
iFpN7Xheaaz4rRHNW+PTODSh87QFeBQeGw1dfZsoUmzLPyNzBsHG4JOmK6bdZp1o
uiTJadol5LDjoqudCS7cdyA1W9MfxKy5zeTEQ0H2KoPeaRIXgFvl6YEJ+6npOJBs
hJlkUqlFdohaatC3FZFWrw0CLWBl+LunxxtzcrxUpVvEt7PmHp3CUhTdHKzEEAQW
HiVu1IID///+70cb6OSAYfWCFO9FNLubBj3RMhe66Ot+HXANGZd3JdH6++YQwi0/
4yArHJe4p++NZEmquB93M2oMUsmcPY6ADQ1NzPBGRJAEyjuE9Sj/cV/4cgTOWaEy
t4aLxzSIDDnaTw5KKPqlsY2qhSxbU3IhQvA3r9C2VncE5VKfCAYPoU7pKAzGRvya
AaTBkFE3hP4aD2epgGbaIsumIjpYRbZD1IobCPYl0YmCYZf3JnpNAkS3gHLL21Ua
yRt+Oqa6/3ASaSfWo4fkAudfJ5CoFRNRqWcc78j8NukVay4MukAmSDSjba3ViDXQ
O82qPi3dDXknGH60+Wzs1ey5lDc9F6XXXnggvyqVHom9pDcd9QG3HkUCmVDczBR2
a7wPCMH1/sFzE4rAIZ8hEV0K7gcczY+gkhZ2R2FXQV0YqGjFNoFn6C9a/VEmHqd0
7k6MUcV81nrcVhuOSLB5Tj9EZ4w5IHt/gQAQJhY1BRwlN7Y6wvpZUophbwqBtBtO
XWx8k9LVfn0goOyKGJwdiqG6ugBWQM47K1HwxXA0LJX6t8w2jv13XYfo/77+0hqU
rJqaIx3ISNMpqaWjoxImoojQjCyYubTm1iJNTIueI+2sk0OrhkBk83LeDsnU9rUW
GNAwR2unTs2jsQd2FBHvSZC8JqoSY6fk79fDw2tAizkpoGMWSqIjFBclebzDwY5D
KkNmrqXP97SLqUAMUT6ruKwIl9XsrVGPv/15su2E4vsyVOV6n/8W6CbcDwBCGtiE
j3dqYcyhq28Z3oxDKReXBPMHQ4TSUYV9G+w1MYEuPO472l+rLXRpalSIqahxBCxj
vdZVwWQ5UsNuHqOtw2AAAFszKfGmZC0EMm3VtES/bxK+Vrja8rNLxPeV3plpORSq
GqOqNpeW1wan1HOfbu6wvnASNMnyFq4zeZFvnYrzfuxXXv52IPqz059aku9aaU5g
aPvNtal4gWZu5/aieYn7UGLnB44KiOTK6ADSNkjzOzUskvgKaPMmRaewa6Gd4gdi
nBtbMqb5goFnztyytbfX/BDLLktsPjacF7IMhVpL2DSmjygPIHM1f3PN6JHUpj3M
I2xbpRoaXvB6nQoOxdFvneYrU/Nb19OADMkmAsbXXvee84NokGp3VflxKLg2Au+u
PA96c8hkZts+wdJwsxHAOwe1rgyS3+uUnOaJeEczDGxljrETu3WORbII0JgTsUvi
cyyLjzftqq08989/u7021yRo5cckHbxLM8qvHFbx9yJqtNxEyfa2+QGp+uPH8QDr
4SzJr6WnLJ1mJDVt69REnMaiuNNZPLM6bHHSRnkE4lliWCBP6aofLf3sNYmYtGnD
eGtm6i/kzJ3+55g6GRAV+CoGa6OVxJNG7ne2b9u9Ny1OyNgV2r5PfrasTXobIBJq
WGIReZKB+OKY6T+NApPF/hZlp7jgia7k+p2LnY/lJaz+NPlVE7QcpHLKXdA8/qIT
3lpvhbduOq+q/NOdoe2bjPBNIKihTkTbZBzw7/4aHE4ijjLR0xv8nwKHLIxihxv4
nQBfQ+tTyFp2JB7OfZodo1bfbqzjm+iZAF2XkfwoXfntITC7OjJIuK+F8c6OMdpU
vdB5UXQ6fmvWBI+17jo7iYo0GCxF1W6GLPOVx6q/61Cuv8nwwRCv34AvVk84NR2G
RUfA51x58ijuhz7+jauN9adjzTM7s3Igi7M2Mfh3Qn4/vUFmkgMs1FhQMlwoc+Ip
RVrsWqwPchiOsQN7Q3HzSmvnV5r6vklb/RWDIRW8dg5EfYtyqPbEPq6SGlNQJCrB
OVwovarVHcApLnJIj3DuX80V/QdzUCSvQ/ledWQ6ljlhgZaGdk57E/JzRCs119Iq
ETXcPQsODeZsHonJ/CO3Jl90lNkBvYreNZAz1vDOr1xhvJzJAZbXJO/CNCkaZek/
NgqDZ0vycDk8eYNsoSVXpNHkIzrGHR8ghZ5NnHPX4gdK1hOvfHkvqyufs9ksErjz
fmf9ESRzUNgkr0ylYStEFFBJBoCUxAuVZTboBgMSL5INqPEO+lcV0aCkoMvMt43g
KThSFVOY5bgADYViXvf4jp523W8J91L55bBmR4iw7mTgBhqq6sG509Zc97KwGiPh
OO9KCZ/QoxxgJK1I2tTSwmsJd7/moDAvb0wlYwX9UwPc9Zu/7GXzxhWQwmcpSeBq
SMi5ICw57nKJ9dBARPdch3GJ2u3+ZstdN3CUhBw6d3aInLoKQdVwXQWx899omkAJ
BSjYrOmNnlrIP03JLgiwNdHCcsmfXi27HgnrqMZ8+4uqro4d9thiZ+vcoUQ2ZgNY
Pe1ykrFXBKahLBfmnmJXHGMODEB7eNCXcvi9FVZ8fPLvEaOXDRvVWZDdB731yK4b
DUoD+Szq06JGuBc/LBbddNJX9ngFWwHPXp7KcUmY7VaxUuQ2OAtMnhq9sXMHZTS4
E14GgzjEk4Jm1jMR5HbIoT/zzyvoV5L1ylJ3DpfRiFIaQd/kpJMzdu224ozE83My
e3tFLeKBQH/AY3FW1GbOs3xnBT5LR9c020MM+3JRWLSBq+AieDbMocLfUyfHJX74
z3dDg0cwwet6EagyyRnYCDZTbJNyiv59aCLX3ZYJ5xEANUH5eyiP7p75TRJxRrs3
FaBnKdM9y7NdhuWEcz6P1HP9UV5It7/NLOCIZ4Bv6NNenIPC4YiVAFYbGvmQ/qsp
onjfuxGPYXD5fBYkhIGCqvzQlrXvJ8jBFl1etW+qRdfI2z0X/tEQ0sCGSB/CWTqY
fj9eKgZyUO0b6cr5QiOjqz3ZgwqUQjHs4eg3L6TrviLbhHhw2fSC2opeR2sgUB35
wORyh59Ui4CGA1B1EdN+7zSZkYkeQQHgUj/eeF/Uy++TiBv3Vs8uC12cv5w/zz/A
djvjHsd5hgFkYhcihKtynAxLTVx7B4C2LAKZr5lUuDygz6a/DnM+h1zneqUg7TUb
eICY8TQSe7vJBYSzsN8QF8rsAZNFLdy53/T5Ensffm74xlk8w/Ln2RY8LgAHJzrZ
pDvelyAFM1rI4+hq8QeOHZcBscgd3Ovq4JK5MmXaC68GuGT6rOjTv7SNqXu9S5c2
5gbx1bCd8AYiwkoiC7ki0RPD5F8cC7FIlWthWKfgy6gv7HSUZMBAMaRIaatKAsfA
yH+LPaT/IUVKhEvQIR6OLhwPhimtEkr6GiRouEjH7qGH5LOq/30HNmQKV1QBbzYl
YSFJo6DACjyaJvWJrBVS5Rw7E/JvTWDO9bC0s7PZClDvlMSOe/a8gBSn6q31Ygde
1AoDndnRdparQ5YjOvAvFpU9D4FI8PaMwyY8CxLcocb75b3WuhSk5x3vBXkuF+8f
jeUgN4rGFvEHAOWqQMlj+y7MtATuQ3C2cjn1GJ9EYxt7TAUM+Vmm1ljwaLFwt+WR
Osp966yEUtBjZep2vuBZxlRvBi3KgUWV8uA0kCiuHbe0Qv+9BHZdTckQGiAysu00
gvbTdNtTbx/e2laqZiBTr/CB4eDYRL28WFUQ5R8pkMae4CxwwvkCl+WwBEFt6wJL
JDcO4re2GHk+lQoMPrA+pqbrMwBbXhEV0WrERYg6UV//bO7aM656qxqnbSXhgyoz
2ilYoNV8gwFBEy15fKanWlrF0rZkpxavNKSlEEZILlVh3Yw1zh3iqJIWSdbNiA+q
2LNgqnOBD1N4BhS1HNi2d1KZdp+b6Qzvdctz79i6F4j6/xz2U7Mhm8Eu8ogKDPfo
mXLYUwYWgbrYmVeAkU0Kd/5zKM5hlwZg13qPwO6cXMAqfrlo4Snl8WYggob/Q5Oq
2gY4AiMg5/OMgduKVsotVO1s16OYzx4eKPqCxGLtPTVOXH2Ikp6QwzryjEyY6eUR
pW+i9Z2FwaXRLBWgD+tZQSrC8iCiuPyiTU8qedTRuh3T/iWwm1Elw5qaOrLc+C5B
hLL2BxoYa8KhVjntBgfESyZbSV5eTQ7GeUVh5RXF2Li7+5lOkIwCUNuzYl1C2sci
dkbMVmMbfdfR0N+VQNE37ndxTSAxkx2gsvJ6UtWlAq8rpTkBA6+rDNHYd6S8c6FT
AP47Rder+Yb+ttA+3yurZY/T9XxSpptMGE22aFGsK9RkzGqeMfNNZB7HiZo/+H0E
t7BLVy5DBQ9AAQoFU0+RAsR/bYh2z1UYrz6bO49WxVB5VMwtBL1n4blAfG6Drijm
yvji8BAghEonYMW0R7NjW1T5OqogbOa5E5Pcf/r0WDSFdiwn0tQmE9NlyPLUyhMx
jrQQK5BvpOzsG95krEGV4vUW1nOupkHQ8p00KjhQPz4h1UCL25YsGbVg2XAFJYgA
zoZSAoAmnV64sHAPGZ7M+1DIn4XWm6jBVfgwDp6BE3RIEQJ1Z6k2diCuNPcZKazi
d8o/1KNR9v6cbBDTLOZz4S2Mo85iNAyDOob5dCz2qYTnPBk1JZCkiSTvcTeTz7gS
BUl5yQQAlQ7a8mZ0Ix/xDPeytSlu109NXj3nKcMo7Vwh/G6JoGgwKDV+vSD2RklI
KBcKylXslzuhH/j+uU/LYv4YdUqO43ihLoBHO/TGzHkutoFlclgyV5Oj+Gq6K4/E
5t8yPMJaYrokgvXXYiNzKvWkKWElYSNDPNYUir9xf34op6bJvRScK4z3WsESYsDp
RDN9AeVQjjw5v490GqfE+16QFrL+9KKAWgLV9XqDUQfVPcOGi7AU0XNdQfcJsYnd
aeumdxDv3wOYuBIIbbeN1c9n2SfJsd9VatjtrI1alN9k4tKHTRHwDh+pxwLRUtj/
1/rebjDQfqDUeBIcK9DP5GhyWQZXhmnchEOM8BSkBiegpCU5umTW/iREkCOCwIqn
106/i9WT7RkPZPOVRUignBQ76436mUYjdbWYUURPT35SoA/STULpyBkfjOn4u3Ql
5OUWXlw3CRzeqZVWBqWAF65qf2Jo9guZueyqYp4ITh44nIy5a54wxjX3S7Tg8N+1
r8r2K6Z+syqPEUZGBTUYTPzoP+9lIrFeCoKDmhv5fIh8wn7lirzO1g3bHo+/Zk5p
PJhOC3gWG5lpbWduunfqZQw8Uz1g8cWN5+VSPDqY6qzgPvn0+FPo+BMK7qp/Q/3k
eLcx+N3L7YDor5QmiHX0ZvBZLPrTDhPKqxfXTmw1HOz6eH1QR6ObvlWCQhzOQsvq
an+ckv7zX6kXCvZxu6bgYIawS/1XXfENSpJ1qaChkmJWoH+CVzqRDvej4eQ8oPGd
VWo0RgihG+Eo5x96n/myWG5z9u8WJF201xcxy0BrhGPPeTQ+9LxXNSW344L4S43W
B6hfiYVP3Mt7krwFUn8ZgpNUmwlr22ay+1YtBlvtA5dHApzfyas7kX/SOlYWK8gt
y3WY691nfTaK/4mtEuzE6cBumP07jjHjcSfXeOWGacKZDsL2ivTV0snynhX8K70I
/Fn0ni68KO5UzCtPVlgCxhFtumUgnvsZO5rA2N7xT4qeoGg4W6YnG3Net3S3Pif0
VRR0JPU3jbtguNq9cXGDMazQ9Di26y9SicAK38E8v2WxpDB1muPpXnrfZVgErbHx
D85Blaag/FS9BrN8wbe3h+4dm1Y8ccZcWJqIAWSfl9bax79soXvXjl8NJ+IDtXDQ
a2OWsjI4DFB56INUHOTbyCvUHsa/Y/pJ0ebxyyirOUIdMW1MNzO5ZGd2B59YpN4L
ak/HIkzu6YnHsyOSjdIAKe8OoFT1meoYaAcOT+V0yza5sanXJoxNVsHYhVy/c2PL
emJMGu8hzdPWcJgi7swXXdDs682w504zYlOc9ah7c7EjqHY6DFzmnftJkAqQuKuh
mooqjc5s76LXkRambXABAxzL9mhi1KQ2xZLGQhjf2WeRHRsx6v5X3nyFcRb+Biym
kDx7mLa7ffY1SgDM4B2C6fzxGFLpUSWmFFBwPMbO0Ad7q34j/eQkh586bb+G8Z7a
BZ67QQ73VXENvuQgLexTaoY/dVnC1Yjmo7XbgkpmNoRqGBoCFh7yx6yliFDQtG9X
Fi8FNhZ9BJ2kdU4ejcx+wFPf+nKSt/D+gm33YNc+9gIJpykyJeE9fLMMhgpY/MdD
ts3OK6SE0Y0HFKqx2r/4v3Kbu7uQvwPdJnR1tB7adAYBd00RuBawN829SV9l/S+Y
CM4jGPwTjigcQkIeyJHh9aWrGLu81c5HDlx/ZVJTVAs4+G7aEBdhGp6cztu+Ic0z
UFKjEM3Rvm2/tQ2JmvTrbakyKwB4q8vEkv5caGxWjT/OD5s55MsYp3PsrkcD+TtZ
2UpBEVzqVUPaPHE6a/FMN+0R0x3zx+NMb50DzASjZkOqJPPNZfXGfwnFTImCbB4E
Blznb8wncjngD4QU3977PKRkP8CmQx+pcUQPZ71tbST6GYc5xsh9RPV/IMpS8ESE
jrEvUZAPxqs4fQPh2tM3BmT9YlS9oaRDsXfeJtr58wh3x0wdIh3hq2piMYNQs9KX
huIC3B1VfTUBthAuWzT+wHUM5W+lR6XTWhb37OwYH4PzZC671jhiVyu+tbyf52rq
wjdrQY0Sc896ztL2P6WTrI0EbtI7ON3Dgtmb8LQjpPjuO0LL+INmZdFEAyugGxnu
A0LGpfH94ySpNhwZXZNiuSNqDaGq/C5KMcDlnvlFxa8JQC9tyj5qiFp1Aw9+jZ0F
B1K8g+JvTbDz6AWrpdpXX98NFt6J4AXErDQ1hERfGmBIGb9hCIO8Njeu/UfETP0t
vt2tq71TEb2Cjhj4x452ZPqPAqY2TQIYY1Rl5mbEi5cEfoxIKWs7NKrcwO3QZDkk
Vs9Q2F07Dd9qAwQIIsz4IXe6+BF4dQKEohfM2iI+HKhDSv5IdQq/rADMii62Y0/M
KKtucsuUNQj/ZTqxq2MC7NEZ4XATpyye8C9AXR0FOKu+EjqAzONRjS7MrNIaauTd
2tpqdDU/grpvUstmG7zkqT2qEfGZjWR1YugYPXggbz7PnDu3n0tvwGBH39xxGHlD
0F7u6SzSEF2tHVukxdj88rWBL7jN2F53S9sZ1GUq1BF/mnRQDwn+xap4X4ljmIAn
8zP28fGkBPHL7PXZt/JHiY5ZPcUtV+l+tJzFjStev4nKEO9ZM0eGG+sqS5aX+7ze
rQ+QCW7ACxgNtjFpeNQyEtjSclZPiB+jJ9tscX+MCID2U0E6G+sxOAAcU998HdES
QcXLKhX+FmHISb/bvWOurIA8T6H5JlemabQJOm5rV6ImOqJSv4lgkdJe79t1K66l
rUnW6l+WF0qjuux5tyuFWrPo/5YAKn40AzbE9jNcBTFuAl9JkYLMutaxd+uwP0Nl
so0cR0SSzfR/i62u+hi84w7gH5G1rlg47DRO/u8vCDgdDKGmgn1VKdrrYrVXursB
C7RFuTiWJHxE3IzOUNA6fAcJXhxjE2Ph85U8NFGK041T9ZSSUrveITrqi9JPLAhg
3MZfeioS9iW0hqLNlwPUXEeLizFtjv558hx5fhAD+5Orj7ENvA9hbXf/mEBEj+28
8r5HE1oS/QyNuZdfSNgW1u3A5/1oTj33xoTaU4WSttvgy+Bs+xnrr9IJkSaL5HAV
VXX5Gr82/BVI9MUZ47tDooSX/C1WBokltvNbWvBaRS1BPjHGM528LiERV0wlsaxH
41RBMpF2Lg94V94YkIbVKnHVsjAnaOenGYLDykYdQszhbAgwYi4Is0BVTDSwYKDT
aD+KUSVkC/Vld/066e8R8WJJxFh4cfUHsvUo/aBoawqqQLVGQssX4BFjwPPT6yV9
bmYJ8Y3B8dPgJcvr13Y9WHHSlwb/w6DBu60MzVesAWV1vpNq6k4g9mhcDaQY0lSp
rvZFt7bBLMbwHmsuImKo/SmQY+l4Xi9z9jeozRjUq1DXKFWNQbpU4fQu7se7nZaE
2A3BO4NbjJEXEzyFPZYupcQ9SUOr8+z3lOTUncLMHv3skXPKOVt+xld2obNreCwL
XVBWFDleZkYYmbBq0GnxcclGzzRJIHvkxukYgCnn+jC1zRX9yRNE02jTluJ9/ull
leKwoFAsS3GerN8r4yppQa/DFLTEe06b57n0zkmfZndFG/uiNkDm1z6FY7NzcLLG
7gnuFecUO11jcrJqSBe7YMaF7NwPz2tiX/9Z1X+li8d6nh20whhn7r0jKzV0nc6J
rmCeqhRX3e5JI2wZcHuwtb7mRuRjFXthQh7h/74jCNK1IbaSjKdOtrX1ZsqRbHwN
h0RmhKd1kFdi37p/xUyM1iUY26Een+eFsM2pISm1BxvGpjoXWsiK/s7C/Goz3jqx
qdAZnEmCuNl796/0JFNb56MaIu2Bt4sSTL5I9/Rb3TKgG+iokKY4tYru7yrWcps9
xyo1j36dPjJyfxgUtK2AoQfa7r1wdc8Ic9Z973pFrPBOTRMA/ENFtsTAkvG03xa1
pc06iijCCw1t90bj2Tv9n7Hm7j4r+arvJ5Qv/sEvJy6TqvDQX4FTv2dRgqLbdRcP
RXf3QNDgSLpSxZ3Ud32MCqjCsygZLjb9P8/Iyt4px3lF90EX4YtWe1jhIxouLKWy
tyh3/09py+csowdPEpPEgs4hK+2rHRWGyXIlxRLqnLIx57TFEudU61EgeXIBofd2
XTRST5nBkSkQF9UPVLmYwyoxonxxz5dDTj72wW4d7l+gT74S+zKuWTbLNSJTVFK4
7zPr0sDhC3MAp6pkWPRbQUkt13rH5pZn3s01tsowykfzRzfsGP0AhNrbfrerx1i3
ENDI4A7iCQQpWzY//2Ael0WXI/bduHejvvwi9ryQWHlvgJKxeb+gADr8o0ECeaL3
tBbsTJO60Z6HtnX6598G8XH4f/wj2QXSjUL3T+XWDScIlNQ6MD25Pzplmqfso7v0
C/P91Mazb+woOtZm7IqXxroysUezpLjYJnZl5TNiJfDSMh/9SfFD5Jq0/wIAwbmm
KWrvirhcsGCDj0fryazWpo1tLF7qGP5KBXCww7agjtqU336BZ3BHZKjaEfrPJBjj
+pT4a8HQlNTQIKuw9FfKfVl22qWrLn/BchTeRLOOUzPh7Nuv6mXEsUJDzUbm8sLT
8aup9zlIaG5amP3f1W8JyA+5snyqqzTyYz3wGeWtxREIK16Rw2muC+AxGtExwG+4
eT4I8SGt+a42X/9wRsPfgBc2G1XreFor1oGCakdBJiO5lvTKREzMevt4RN/XNr3n
lyn6LcxdRC9M/lXk7vB/oe+rLMr4BDgVjoWZa9ACP0LtAInVkMG6Lbn97zdruSpR
kmtTRdCgM+f+JyMaSZpB7Efl7w+390lUWO+fGYuyvNhsXK55hV8LDP1zuZ4F8Ev7
i91PByhOhj4lyZvTQp01KvxBbWfLXAT358qK8LpMaIrd4gU7D4iGBoeyB2xwaKv/
aVU821SaWqxFhMCs4i9EXhCIWNG6Btg/KVaqZlXcDKZ1YfZS0S+bs9vVEIJusPiS
VLUXANdgkIXlSNnY4WcXO2chNdT8KjwEOLRe4u0ObGUBOmNCA/reWD6nV2j3e5W3
NrQxmz6b9r9imqRL2+MbGOAPnHsXPn3LWwIbxdgwOn+KU+jdbPMGdmPXuSirZgfw
eythKUneeXyHTa/1eEhxvwlY5BUVrwV1RWakIbQ8zTcbqPXGG+uj1CwjOOcH2nVG
NlcugerFjduN7gKNXM+Rvz7GlauBnZIQH0tDcS/IWfHuCzJp6X3hQvS+lM2EFxW9
W0RW5HG+Y1NfASCC4IxzNS4v6HVoDwF1iinsM0UI7rZFsrGYM+221qflC90ajC3q
/k/fF0FRyrDfIY0ApVs84ZhKzrp8n7vbHl6fREVzeDABayMSa4KN8oi67h1QRp9u
Us8xE98NFK0ReJ0NRGPqUxlEiMB7GQ48w5I6r/RiRuTzNBIsLMT/oPhFsUyatclD
nj0Yk1OJLfLCpsPzU512RAUo47HZUYkep4EvZIkcXrGq97TLukfTac/OFzWBrM43
GJsU1x0Mj7dZQFrCk51/Sle2hUe36eeMvIxkxalhEnnce54urqNFGhKnuEh4Y/qo
AkaGxWm4Udn6/VqqCPgcX9OOJ7Bmom/1flwvTSZ8ATHrIwqFNle3OepnzbnD9b7+
lisQ9wnQGLi+zHUFumxj8GvFt4GJYI3epEwGWJhAaAqZ/lVTnv7on6NO3YIAcl5O
vrJQmT7W4MN1hnBE9mk0JVc1U+rUHdrrNAFc5gyjrmBQaaN0FKro23n/4QL6jhay
2KbMhyUEPIuIMFLJVpKA9aJzbbcLJDkvj/r30pD62DNHOaWUpFmpi/0Ix5Tow8d9
hRlgXR0xWoBnbRq5aierVzMT+2xXN6t9Lc5HGcx++nOqNLAQeHIdQAlBSaKRicL6
tYFGL2BYHoZkwvE7D3yWnQcf9WLpx6fLKfB817HtJA5r+R6Y+R+x19c5Qv9WSix5
7AU3GlDk/PE/ul6qIFWqFCQhBUzSPlch5C2oZYmK6V4GTFGM7Z/EeFI6N1YHWoSQ
B6o0GY0AGksG+Xh2lvau2POHkbGleynY2XLxC425jdXAPx5c4qh+hORL8rSVvLGo
CucM6CNc2xwt0SrqHp8q+q9uQyp3pc4/p5WVA5j3E1/LB/ljUnmHrER+RvTnxyto
I/Ttj4x81yeZqhe87dZC5C1IhDeBTGgyYw/BkYRA9cEPiVZHUwB18I1YrjFe9zHf
BDmD4dfZbY2JXQhRNeB/ej/IFP293NubicE79xtjKZAiPIcnk/36u0PSUCmkmxPi
qmACpgdFC3H+0LSwK+coghFcR2XCet2FcNCqQ7lvajNK/C6gADPPPjSrz2RYQCOu
Qq19sUC2/P6uW+4glJvAWgXrwzskwuX5cGV1c9zCKYQtLl9G8cHjE9c/Bxe3mBQs
4m5dJtUsPsBLsab9LF12djRWbtDH77n3Yo9RV+g/68qKlZiLlIDROvviep5T5H4F
bJkR1XgBhIONpuOL+ZHy0dIzS49rzs2r6iNWO63cNQYWhzd41wu5ZDSfpTDTDHEu
Lz9btTlNWy4Yu9KiBdeIw6kqi2DmwjrNx7uTCSjuzVlcARMnHmtTbSmnxJ1jHYWZ
KCpL8Kni6C6zVwwOPxvLAvrbHhAXDfttTsH44xfeh/8kgppSyGqasnmxqBW2w4kM
MTcpsvl7R3HixXC2m8pcXfm7IYPnkmw/81MoJsgrZjwOHhBHZnt44SFDUZpkfRbD
z4T2HrDK+wvonlY/3hcvPPjBlItAW0/DdfxTlAviXqrYor/OTAvMsrAU1CBpbh93
dk9rF4cfNliLjqUlvNEo7jLgrlsWLOkddHe0bgtv+LGzKHeoTncngoMWyQ/HjJ1H
rLhPmwdFpQjQX0bsmCYPlRgba/mXIq2IW1DWv3rE7cyegg+GWyjooqolL3HJ8dZc
eexInUt7MkZHbEcP9Jo6RnReM/pskRXkkdYH2xmphQ8qJdC4j2htUKZdY8ojZZGE
bOgR1BASOFXXpfYguQooTQlhlYpfM4Cxi720PWA8oKEcFce86ZUMTuRCBp11nJPl
ybx1bkLZpoyQUPMg52jOovik9uPbmo0Q8Hi1CxNuXLlk06C9iXapIg5Zes0c/kcr
lEVwJvDMdCDFTeCyaJ3VnvfMyotBL15C/6xNIeSJq3d3jopOPsNlaTH/+LYU2fmu
gkOgjuzBmNfJNf0te3JiQ0M2M8A13a18DLAl/jN2sFCDSGl8fb4/P7K+ZhuA9lbB
LIrQ8cgpN6lOi1g9ak2vPC8fHoVvcjgQFe2vaCIXeAEFdRiIlPqDkOXwkkhMj42J
zGjZTXeAKQh/+zRjSIAIROy9iY9o0kbyHHAQi/FOiRdcG9KwVgD42pu8AIRa8pcf
hvS3mQ2ggYPlBKiakcyCGoeJoeyh+6JeISiaAXDYWbImIqq48hXcxOC3KkFGa7UA
Q1lE4PSXjPbeU/mhQ7d4rcdFLAWAvjVEdvl3IEY5Ra6tMQwDUSmTJkoMVLsRGYBg
3TZIN4QBym0/drULXPLF0zWMUHkzD+TglGL6kcdk3n373ivhzoDlJ7AwnopTxfbJ
t7+WsJAaC+2NqsQRCeWyO7fhYU3I1hBXu9AJwwNqgCJBCtjiknxyXgeurPXDa9mV
pF+monZ8FpMgxSw4R18z/JuoDb2IJT9RCaTlOtgX2mC/aV0aTtU/QA9t7hxBRVcx
du+P1oAipQT5vuBuuNNlfHPQN1/dK2OpU/nh7+Gcub2qtJY04CP/IhHE4Lirr7Qv
zSsB8uZ0sr4kSXZX+fT/LGpw4WI6J0FB68qEGHF8WY7ZExLGZodfP6sXoIkPWQXH
P0Ip7iJuXeFEKvqP55CK1WqCvsqpxCnp9w+fCGlPGSMaKwEjzO23h+qq/gvIaayJ
Xbhha2KwdDnqf3aJCSeE1kRZJL19a2pMajdd19WSzevXzU5AHMa11yKX8dykaKSW
RWW7KfUZDAV4FrtKVDlgMbYTXIMfAUdB1SPYe/38f1Jv0Os4QdNHy3+EzW3m6wBQ
BhRh8tiMLDcxYZre4tLk07lvIOU7YgfGJ/455DKenTs5ZymW9o6ifjP2yVSBc0E1
HpIMYRFlnXsqyWbeM45J7i/GWz/OmzU0frij7gomeKUqfy/E0+V+uggVu/gG/Vcy
OluIRwEKzn2380H8PwFp9CP+6u7Wr+QsFRwknbeZFdo0vZNotGtaa04VMIPAFPAk
z4ChOl4vODqIVjF8P5V89mVdwCKIVRyO8csKf8dRSfxMopSvB7BbovHAKuj2gcKB
tAWIjbr4/iQVXxK4AAd2wrL28BTguzknY4dIZi2CPPwemjqGBrbSH7eFZ8/5b5wx
B+/RGUz3fP/vjuRzhLmQNQ+TDesmfd1n23S738d2xQypW5P2yEbp2ysMutGaVsGf
DnJIkRe74LhV19ZuTpbn/cALsAWZDUwLV4173KffH9vtOU42RNP7Eb+oXcUS3KWw
N76j3CR+VcHenQa0KwRqIKB+H2w8dJFX425gIS/Vl2FTwUaU5abqNuqP12LC8l3t
uEcGEPulWBEGWLgQwM9hZOxroUOUoGkZkhNq+GUCNzx7XNWPvxNPQFfWyv/s70bj
GmQ6N9JMHhdNejttY9gdESjfSQAdimAFwcvPCcNpGHmLqLXVM9yTs9ud4M8BXjkX
lgaQZ3jHnK98a8pI6aTZbrF0Sx9N8yHXi3URYEbApkotM2BTSajpbWhdEXKD8mnz
mqWd2MpIzfsaVK3NA5d8F9+U0JPAH95u00Oi+4AxZyNbV0aQAUvPV4itk2Jn7k0g
c6ORt34EakDaGAQAOc8ceyWMHZPBklkE47ZsyCFmaJKd6caRnIFUyOO6HdC7QH/v
RM0O/Nk9Reyf8XSdTzmGy4LxAt/0UJ3YufINj6t0Xp1UWGm63Y/HkO8HArmSaguK
BBl7/VzCBu07c5H8PwGmH7glE9vmeT4UjEJBAVhgsS6J2HSxjocs/y5XrsyamTnp
Ik0NmfFeUGSGm/fJNvflzc/gzeJxcK7WyLa4ZaIpoSmCfByY9DPxs6wGnScYIui6
h1S0q3BzK42e8TSea6PWSTt5dbjykGWRr3uwrT+uPDDjbjuIGu99tY0K+dShmWHu
c5nDJ0S8nW+MZ6VpzvXUBmXLMCffpDZkhHy16JnlvfdBIUU6ekUDszIzzhL1AD4u
77hftG8Fz9kvv0bT4QdR/lv2bSSxl34+yr9fEZU9W4/sVd8IALCTR1IXMWn6yl/U
ny3QsPh94pa2K0o+dIG+tDOD+kaO18WHCXgJHrUEHbwhvLW2yl8fURcTDzMOGcIS
FbTi98AjSYJF5aB5Tmzo+SWosjt/9q8S3ubsuHgE6KLfYVjUWU4ge3//chtxC1L8
Zcj86Ss9wVwyumAW19oGc7EeMk1whhC2A1YhQDbRV4z2WogJqKkPTRF+qnGJ1pD5
uKvVvM/gOXNgeLQzBUKnHVOl1wOaCmvIg4mQCiSJblBA+FmRPFbH30blEg4z8rqP
zh6vKjcmYoYB+gAjg5XGTlwBL1Asjy0pklutvnTK6w8m44YaKYlu243N3inToTyu
KBjTM0jOB3A3n2gndoEwqISNJuPYyIMpnejiKTj5u9Yr031hefkJyfkWQgzE4ahl
FXCNhBoFibYODb4VG+kzNLbSfX8Gwf5EhQV2fSNXsO5kKMH/YQOIXjT2oJ0V3VMB
tloMnpUxxLtmIwY9YtRRQPTySgOgOC6voI0q+xgMXb/ICCdW481kyTcPL7kWgaR5
iaj9kriDBrWQhNxjAFgkwgWvp5PjsodgSeN8b7PjBe5vhnT8S1+XoS8+nVPs1qcM
wg4k95+oV9G/duwYxS7t/V6W0vLi3U6lIaWPy1T7mKaDsBznCEV74sPHphpxN5Df
gy54wQCVC7TsxVxMcw07Yu7YVQol4+rcudLmEKKPmvxz1XGQxKd5YcClJpJ7lPtc
smhSrp6c8xLQluFzxAo51of1TxucLSj+GrTkOqCXEVcVuMAReYVPmzUs8TRRSQN/
yoRLFagIPqQ4/FsOY+j34SR9jwyvdCrX/xRro8s47yYCXVmVIiVl9q2k9Wy87zaF
9jp66wtToCH5QxWVvaLWhnUZmSuMs5UDQybLnP7MFiR6rlHoWy9fZoZG+zTJ27bN
EI5My0cAZ6TdTREWqq1w6Kf6QivnAV4HwE2kUMxEi9ENPO90vn8S8jeu0kGCFO8S
dfDr7wSVPBck/RPiMZoL34jMcTelvAJp4danHaQq3cN0ia1Hn6cOlCX97rmRBhtC
QLsRNRJEa5sdGa7wUMpb3W8NJhYjCVFLWSdikspG6j+Nv20fQm7CN7vERK99ZawK
Uqsn1LooEF1V/BwT8US5kHcKAcunv+XDqXkPD22mFuFtNTrdgwLNmy2LmDJeWQmO
lAXrHJP5TqAZ9D9mD44FDoJgbpoYf9oADutKS2nTnYHCUzP8PaU9hRNExFB0XM/+
MkqqZ2n3Wt/VH8JZKoD4970WxC12qi2cT+NPWqEyX64DMWgrdPfk5rk7+9suquoU
bfqjC+JY/NpO68nMTbrWCvc+ZJUDBr6wREHQXDuwwzLS6PjAGbFuC6v2+n77K1Jw
FDMh/h8jIGKF4Z/W7IaOAeBE3I+8f2DitUtL14d7acf/yp7B+A3/TP4NY3L0zIUc
laJoQJ8VXd8Ak66rw+5Ax9gy5KcWGwB++NIZO8dNNjxW4dT/ExOnuJOza0a8mOzl
w5i+lB356ZRSiqZIoYCWlxoxBc2ew7XlahHJlqUubDgEQLjyZC8W7wwQci/N14EQ
Hodgun8cSaI5H3SXb7UxAZ9ps52LhNz5PElfjG/hdQH+Z/M+ocfV0hRyrVlNWnm7
nasQFHJ6C5HnSy02BPbLUGHSwIRA1My8gS4iu8cxVxlA3knUzw/239VnyYMVsidP
NT7Z6gsw02CntsJOqiyWGN86QZRG+NZxqZIQw1kM9ukbf2SQfnJqRy60EjtvkmNk
na1+0rNSM3VfOUWMI+VxZb4FjVnygQNJJ+ZeiUJto9/htkJO9FUYAegXiDyj71O1
f7O8vALHs/H+qtiIm6Ohkxz/E80NDfc53Rc6XbH5ir4nmYVJOmFfs+UJiVh+f/Vn
GHsm++DGEXWJlzUfL0DBAKo16qAVCvkHwFTuvnQNzZyQnpnaDkwo7oZpBjezmbvS
SEHswcpx8iFlQHsA3vFsdyD44V29Bg1zhhxxysCo0i+23K2p8wRn0dcgNhgGtpwz
2glMMyrUa7rQX9mvw1SpQ6k1OYU3OqN1D1ARspzlsuEj0K8i+Y98/HbLRIYtGJqO
2kdIohssF0aN/9L8FO/gJ1cIaVvGPNq9HX+oFNu4dOnEyXyyyWN6AXHO32/hbanM
Y2xt5pLod5mElWJ+MJ5eL6WINd+cKqmzq7MxB8YMYIvSGxCxf+YwTp4O6mir4uxd
hhAhuIDp7FPwuZlH7qVqT/n/1Lr6lgNbt4MW0sc3bt1Qg6JzdGdqKDBKRIPEF4dM
do7cYlMKeijiUQvlXqzBD5ETcTZQgpwUSraniFrhrB7CP8mtpzl3ZOjlkzF6vX10
tazUaH+eHZZd3yHrR0tOatNsaFrtMcCP7CJkFTgY864z/FNY7Cqrck4mq80v3n6j
SrqSnx0dUOMSudVyiUUgJXnZ0u1bDzB45Fo+8vigwaNhnmdxNmHA6uVT7/GwyhDN
a0CLMCLqL0TRCW7fC/lUgCHCB7UGthejq+5vW7lJhYpR7Tw6qrV8Z5sQsK9G4fxi
6N1dApEZ00s6iunpfrY5oeg3wjPl2/LE5TK1we0z9a3CjFCaNrQAMbMcsXwun8IG
1rpxwFcdYi2OL2jKH2saLnRYZkXNKQdm4RSuoLD+l79b14ifjcDew2qVBsC23owp
r6z2uqTguA5RqUJ6mdHnm1qS/NcX7rBK5RBqZXsudVXM2kBSWfC+kHd/zpOXqHIx
yIfoRqET1Q0ixKzAiG9VSrPg8UonsJHUEfKbJ/Ae3kI3UqcdE+iZtYOiZnzhKuFD
C0N9iXmOBqQOGutSlWwI2ipPfhdvrYC17N+jBE9NzH36zTvDDjaqRkGXwsVSjW9w
KTzXG5AgJqAEwMI8OpgylfcLPE1H2aXNEsETez8yiLAaB7o1EgpCTX3qzJz7xXa9
AYi9ctJC6LgmvUuojatWSo0uosEbilH4I9cmQBixXcp8i0Skpl2r9fSyb/AG3sSL
A77C9uDwbwsXZ4IP//Y8AlrYqpBxoBmUKWGMSFG5mOIVjH0H+SQk0a/wB9uRhmtp
4vGTrHGvujNULQFIiOfIeAUTunKBPEqtYyTPr+SfBbaQqojxTRt/q88RMiV61p4C
lSIs/QtyjYcCGqwv9sHr3jPsnLsYwUa7rCTOue/gNxAs/vveeZvm8ESdkwvFk4KM
nzSKAf+a9+lHwORmb5wX2ql8fOBo74jio9jvV6f1MPWCsa+Ts96WjMBJAbJtBvvR
h+fnIcTExmWd0yjz1eLdKZg00cAjwaVHtfPA4749ZyKQBzT2duTonCkMEhOEuOF8
PsaHySmra++6hEh1jdzJQCPTtQAaZdGZS9NIduC/jzDy8xVXSXPaX+N3Ic3VLUUd
xA1w4T1T3zTSn7L6SEesrGNaz+JArwlSXXbmqxjYgmlFuQR6l1vrmjgHZkbsBopT
prfWxwZV+mpeO0ybwXx7thfq7rzALbLXKKHX5iQS909ampnN+NRKPjCnhBmzLdvQ
fVF1mLeyQ2ZYb6G96LGOGqfGJd4PutBkrnhCq8zY9l1Ndujzx0noNuMfkcsy1I2M
M4plF8aBMgpSA7pXsAjCD6C+9p3+wSiDi0BNwBPafaIX8ey0tgWiX5t1TEPYGXvg
/2A0czID9RxqV8lDIeqz2dVSdXrCu7LfaPxYMCW4MlapYuEvBMpcxSbNh2vk/dXE
ba425w87cO5aFd8u4yYMfudrXYFLWsANmTmwSB5aK1WRZ+Zmy/5d1QqAzopGofWV
ut2IiCV51LF27rwmjrJJtOmBd7cPXsd0uI6z69pxv8prmqqkPBp02Xh1DhwjK+8R
aoIXAIiHLfJi14DL21Rf8440x2HlYaEmzm8thghymxN+s8iM7ung+zEr/0s0w7iH
LPUtvw4rarSbNJ4Bq/ej0n5+Cp8cePatYI6WRZg/HO+/mA/WfUQJsVyYDaSwmSMB
UKOuhReyua/ZnX9US9rqSP6tw/XyhPPMs2kG3dCskAM3u6Yq3O7M8Iy66Gl4b6p+
fnn6TESuiUY/gDPumkYxdzlu5tj3Qaj7/e7RB+xVTxJEfaLLHPjQ7ak7mzkitHZi
pPZpetOgL9zrCOlfhlsZgPRQqL5XoQNMyry35Wp/mDVyyd828DKotabWQa5q/nU0
KRGtqy0fJ2wshgsRAgANO7g5o4TsfXUOArGfON6Cqxx4d147C4dugJan1labrDvv
BQalX+U7DaHzfDlLE1JNuTeK6Pv0AxOxTnMCWA5oJfmexiO4HDHBPaUzh/hGwORW
Cr3rmz9daD++mYvxiIn6LlV1huvsprAAC9dmatTXC7MT66o1rJt7AHEkCb/Bmdfw
WAexozEjYTkWnpJR8wJZqSaXivyaxQVAX7XH6g704c5GV/2C0dms21ZrLjT1RsIk
DExkeIaM97+wIoSckUPsINWAQjWlbrS0YuwDLiMaevUcV1vRuyNmdygMqpo8symr
i9kuXZQjanXjMJnfr1TcyigBg5rs1CygVw6puUsqVhhkCTdzDLXZbaro7ftCHY3E
KDv8pC0YXC94lPDUzVPvTb4RwPdt/6+7x7sFoSXl/2Aid7YExUXa7OlyAr9G/Qwb
R2op46cY8CW47iU3evGf0Jl0k6ZNL2KCl/U1fxSUyBC91yROXeKpSQyvHhvhDKgO
577+Gpd2vCq/+Gmm21gPLRQ82tk9bvolbnrOyehbketxnWmVtMKnIqTiFDEJrJY+
RAupjwZvvAWdZtNRN5OE5vQZ1JGra/ou+QXBrwSeifuuZaBJ1/whrtrWwNBWJ+7X
f65P8HxHP8dDPkXw/eanv3iBM2JUD1budsu9mdTOcKlViQBu+Gl5B6tzEW1MgNCi
Fl8C7fIM0WEswGUlO0BfvykuK/DcFMgAe4LqwPFcNpPExkpKlkVuQ554tr3jaP+x
9bNRns2tO97Syf87LU95f6n6MA4fxv54vepAqgYAwukTxJTlF2A2dXB6iPnKJwu0
zLg8VRnAUdafiSioofrurz5g7Txdomqwq0c5cX6sXKGub4wCyJ3MzvH01hJupo4i
o5yvSbF76bHwKfKjTwYM1ukst5OBREWWQ/Q2XsbY8Q17Nivg5wsOHW5xcMQs7+mB
3XcrZ+9HGSMj+6XeT1RCIEubDi0DeiefPVh+xS3vtthaK7UqG+6PfgE2lD6VEIcM
mVcMDZg9r12Y48DEeEovpmTSDYMVgvnMj+hCRfLDS6rIm2q02FElojgyO+CgJyOo
1oyNzZYR9NcCtWq/pIw48oBHgTYUU/QIQi4knOHZ6d5uHSjk10Ptw1MS7AGPYTEd
GwIXodlqrUzYeDZogjkpW6AB54tjeldKbIKYicuxPK4cCLrq+nn+dUg/UOg64yn2
7Hz2ZCNWLE24zyMvvNHmcySbz2Lo0dHUIn0WWvYxGFpLFaifAwlnzUtVJdJ3SXrQ
U/F3AeHPX+2BMyG4+CjMJV6A8BYFHXgNQ/YcbD/QbE2ZQk335+hA1Su8+HC4704Q
EgJ0j/W5G/tEp0c/qjAtTT7nGB4EZH09zVThcm5MJGn7Lcgm4rl1I+Vgcb3/ST0E
e6f3yE24w9WUFGYKHyFZh92YPPdgKx4ldSbnMOv/AIHWMl95rX47NMSMixn2BON4
D1Y6/Cw9oVgg95WM7ClLh0l48FGMw2oo6SCDCcDvGgHaMaTvC6JzJnUgNUvdLqL5
N6NuZ4g+jzIt72FgVEJaLbAsjuK+1TItWM1As+4SDyv4c/nlpqGhobIPN/ciPgvw
CpN6D1d/FjvAUNLxhmuJdW3OGdZECg5K+6EeEgvMxC7qSqk9Al0G67ROxIU8F+g6
rPYhmqBFU+CCoxL1hcTed0FSYohq7f3RwKYlSplFLtTouu+15rzhrGVATRmlg4JO
GH2DI/nE+yrRe7DCQlkfGPhE9rqMHjugSwLwq+mzdSXjpneyqssZqkq+G35lOma1
fz4A136/IGlANpOuMZvxD6BTyQgVsvnxIL51YXFf/07uwOGDUJsmTn1vUvrOAYCQ
JBDHdH5sOR+9bPPD13wBriYoJhqWrYTaPw1kGOXU8ejDwmzJLWM8d6dUJ6GlcGkg
NFZfgtk5L/cKnHdUb7mbpkbq6EYysZ1Q4nOxhGkN261P2Y91urhcxJUZUEjOxlA3
YFooFaTASqDEJq1eq6MA9H94g3Lj30+dSdXYDYZE8QeWQN8AhFHzhopTJBIghR4J
LYLYTNIhpqV3o42FlGC7Ky5DTyXyk38moCHMYxtoPzWpJGvAPgmopC9Va65KvGtL
wKbuRYtJuhurdhnVVr+VuJhhodtnrQsG7W7aCjkCCsQ5H18pz70sNdSl25N5rURq
JJ0ujZvKf6BBG68unauSZEkJpW2+jd2k+XfE9XEjJsMjFRMSntKwxC9zk5BbWLoK
scfeC/Tkrlx33XyRYTfnaLv/ThmQ4xI/HafOIIzK16I6UbKWLqB0lvUlIRuKdzsl
x5+wb30+3H1nIaUuCDLtO5Ko3f37jfbDOOcVCsAQoJGM1a9SMvceWphxDjxDK3RT
tadzhNvcK6tl/KsmBkCSypKvv5y/z/s8Yupd8Nvn+ILixKnanXORNrhDHRB7JJcg
95lOu+xJkQUgJ5Da6GssuRJDuxyovlkTpKePgROAeiraG60QtT9HVIq3L5Ak7Hsx
tjwgvH0FMVygcFj+VZujPwfh5POsSA1fBL7mxwmqXpTNCq+0/G+E4nphfODRrvFA
Kh3QHGfv7y2t03wx8axXQEg5OVOuvn2znGOVGM15viuOUwi2+4fFOj+DC/deXOyL
s6Tt1lSGy9ZK6YsmSEw1rSFLqdPGeNOhUkH6nutK7NirCO6AEWTytqaNUkdLtiJg
RztNEtpvYv8zXT2W6wIdOJRsubc5epBSRfuVK41edzUFy1VpKcP4V1hPyfn+36Yd
uU/SaNTRRSxeXao5pKjd2NA7EC2JxtngSmmDWsDmrgF59Y/URUxlaVOiC/DWjYhv
mYdEmViAj1HaJXXX7nzmuI1XXjteAfEzHMDoQebmtGBP8nxkdfXE+1LBaS/usAhb
7p3Zzz4SaxAIpw2cd8iNCKt4VabceVlF1IvfdSm8h7PcaCFJ08DSSPFR3cp3Oysa
9aGl7T+eDPWToe3QNLWXF8dGDJTHZIsqzGwRMsSkIvKdbZcpxCRSg27uMaOXg610
NQkBez+7hB9RWs750N1Smm5/4caaOqRK5vDrHyfhxHFpiVJWHQLJUFhAAvnlUB2+
3qt1sUbNrgRyb6lC1w3rWN9TcJutCFX9lJTovOF5976g+bqvyiGjXc3uXZkJvWv7
8Wd7lev3Dr2w+bx2XVjWQ5FY8pJzI+sHPvkkWQn0EahYH/rCK29K9/7hva2T0O+/
XWCxby03FahOmzi1D+MZEtiyGMWOQa06rzIrq9azIvl5FNB6oaYjBvoj8H5mOwDX
VcqBWoSawWduHjTZFffOb2Kv+nG5E5rl9MLRW5nWow40zCN/CwHTXpChL75SluV7
LRHP3G37vLw5eFCNl9jd382fBx6916XI0NBWJ0bQQgMJbxNGTnG3b1xFNnDVUbu1
RjjvAMtyGtGHvHaJb5u+tgBBM884367jehjZPvTrUoBnn4cdeyd9weVHZkhJ56l+
7JCdx7dRQFex7AC+1O1/oeEmjeKNizHETyWAH6EDrPKM+hdYQRD0tgULBIeFS15L
A1P2TTcaDQkh/lbkUFn9auXyJpnDnBMcrz04Va8ZTVTWhIGiQbsHJdkIi++a0wSW
TpfG9l1da14/rc2ApJN+NP00rxaeRqQJ2pVkHKMS7TSyyiPI0C8TnUj/0eVNXeX9
nIA8j3fxaDW1issqd5vJuL5w5p9XiHQTL9wpK41Ltly2/s09UEGM04PfPujbmlIQ
L3xTdfBCuNbzbAc6cH13/7IyPdoTP94kRQmFUq6scQg85QuZhkadzjZpO1RhFwHc
N+1VBLl/xs2aCejeSC74Ncuz0yGai1U+bOGx3L12lrF83Ge4YRHMMD1IAoo1CVmF
6NjgKai1zo0L3oGennwvKDxKuP1d1Gg1MiQTS2bMmJLFueqtH1NU4DfVV++EZIuY
8CdPVYYMjQbgVietzvZ8Ir37noN5+lEmBIqMTRSwKSOW72wS+b/H+ZTKM82pBWZb
a4bDRBgl0nTzrGQgdAF+5VWhk1q651JvE/5tf5pYfVGvMIilXgq5F3LhzgL9l4bB
XaVqKcojWvsNUB9DI1TImkckVxSl8JfbP8T+xbhr1VUyraHCgLLIefkq6wglW35g
8TukkBFKOb/8dsxXYciLvS/qA3MQHhjflRkfmQRn/p8U1TyhM8B23dC4H02IX9D8
vPsSniz4KtzEUG/ztmT0fGjwYgS+brNW5v3DiuFmm0km/ncW+WOZ7geF/E4tWFxD
TKpGFsH6E3SyraecDb8x7A0A3hdim7Kar7tetTI1I+txYX+kxjXeq3yD8NG8mBSc
PDLd0kRWQUz2SBKjmeC4phb0yidDcMw93Pf3vF7RzD3YJRVOdG0+HUElxI4rbZfX
4OSXrm74cQyp2PLQ4OdeMA9OR9yBw7BvmndfTWR0XGoPfBRf1hDi8/aF4JLJT2iq
kXL5xxSVr2fvsY71P6TtpI6JkTowli6wSmHKUxPKBKF+/SI9+kSFo7mwClzSmIjc
au2C8sBD464JbrdsaA+unS9ar/cHE5nuWlTaTGAUWmkOQRjfP/D9NoPuTIxnORZT
5he+8JviIaK5HL6Rqj6fSk0gPz3MBk8UGnZoZH/qsvf/hOR7B7p48S0yAXUO7UNt
xO1pMKe5KTbPj8tyWsvNYOAbUuRKCD70A2IB3XTKP22enFsIVzcZsl/DbL4xMGEp
DNZg996bSATfePSZt0lNzkErMzxP4Q9QaZaJNpnTJl7n/ai9Y3g1lzYp6cJdkxhu
vZgS3z3RYwxPllpF2Tq0uJxnEey1rttGqBRLLtOUKSr7kX9uR9H8nBiWPYgFxHZD
FUbBHGLkZT6zj6AaKEVg3FWppcwOasGKPQ3nMPmx7gkpRYOVaXM9NubgTwTa6wxl
gj3E1d4xyoL54w/aZ3LO5hRFbQHqfCW4Prsh8EdX9HNclJHvGm/LBshltfA0sQsx
hewivHo21IsNicK9vhj/CgzDR71jNxTFZofIK1/KCJOWtDmJpPv1fW+n3W3eVkPD
zh1vrRqsG/hExKcOJ4ALOusL+l8wvn0e0gaVw2d2P+p2iKffr4WNPnHeA/0tM1tM
ybzadz+Hb7Z38Vjv2cD0a05Vi78gnXp1GfKCdCpdLd4C89zjXhUjGXbvSwM2UHyQ
0Sb13ZQ7l0fLgTtmff7KrIqX9FqYybOqv9PvJtllPZeFmWKlTeeEnxsDqyRNMFBm
/nHbR/uhW5jCFquC0nYfYnZUgqXOmhRRsdBBSnfeaqtJapjtUvFAn8MupEIFWbs9
nyvZ2avqkdD5m1mI9HZHcJE4e2h/JmVRM3YLKuD8985sCYsi3GNJTU26w2f9tPRf
IJOJvZ1/fPZz2viHWcavDlE9TKkeh2/thGqDDE/oQQS9J4mmxKVaxYffVh1WaF67
AKEYb8EpV9U7qVY5CB+oIPeGCyrcQgZKPiKikijIksRr1t+9zzV/AM8ZkVUKOypQ
exy5e0XXzY5IqnReyfSSlFVUmJwkcoSfJ2ThQ4QCnn0iSplFuXT7tLs9yBoptIoe
4FR1vx/2H4biNSykj2j+YVGYUKPDbA93jBW+6v13aCJCbHYASTJ0mH4wmGqocUSa
ljXu4yRI6atrZUcNfdB0d0dDxEK546c+C3NaYa8CwuTqcYAFBvucrUHc2WmP0yFx
u8yK6qy0LWbZLnp+85/yI/p4ofUHKVLFe9IYghOULC6ftcTJkNdA3yCVZEEmNAlw
s4UUYRYmSKzxaRxaQzs1YooTjoLOurepyeot26Qyp4ZhS0dgZ77//QuG1zEbu8A7
OmmfVgcai13/6Mf/cGBBQcoFXVdtTFIgRLZqmbHfiDR6YMtO1EFCZx63WCyaSMD3
N779eNYR+7H73TZdD0oBT+7dgs8lZ++3fz7dKgOLXjVW9HusA2Bie/AkbLa0rrsG
dlAqkfYBZagYPcceRcUkR7bRznewdkHDl/INdvivE841d4OY+BvRZtT+TRl0MIxU
1j31F9pAhODEGJMKLRQggmAGS3R448VGb5+bmU6LFARJF2oA2I6F2vleWI7KvoEk
1k9sSj1Fe252pQv82r4kgjFEPjqZBJwf5fa4ricoeZdSGxbOKwpF9pXeVtgkvag/
uY7XxKjpQfHWOpV2E4i5+Ha05K2wJrm/WYLpWVavYmvz3MVS/m/K7Nxr1P+uL/EB
oszcxJjeq013Go7eXnM6MgRJd2IZANtWIJE+aetu+e6KBMqcWcxiuG85ZBNtaxZj
5YTYeuGgcSoZZhOcSb8LYzffP+XB+ZjUH9r44kyS4MMwANeAOHIsQ3/gTfmcXNw0
smBUwTNzlE4f9OHWBTsFPi4IKCpi0atFjHxvLsCyRDxtaZzLnNhau2QtfPeGfDnp
QRfyrxpXX/WY1s6xoNAKLxBjMbMwMySeHLT4HBuLDVwhAtKsCREm6sVvCwiT9VN+
sq1C4rfD4GiVj+mE7asO5A8Sy06MIPvvBiY6R460OJhKLs5QQsYVNB1y4GwUeVcH
SQva+nJlzKdU6yguGBieuVa2xPiKt1OYCT0Q8YzeVe9rizc7KPpCenPEOgpcxjmE
8b3U5zBx5HeWl7XIzgGssYmHoZsQbmUbQjUo6/GDhvbr1s4/WyyFdBig0STTdAL4
BHBgDIndXN5KCrnEzVhN+GirKEQZ3Ijml73jxtbrtxWdN7MhGgan394tzaIjP94g
vaLR2VJkY23WvmiUMRVTn+ks0DrObpE/48MUl/BXDNPItjTVJVaXzM5Xei4Er6dZ
fzXqWOJ54FvETqjNQgZ93/s1NR+U/TljqoYvVN0/4jj1XY/VH0TUoEJl5VL153UH
2XKvHH8AZ2IzKRw/o9CpCrhSuNDxLowK68ETzabn4FfbPBB6Te+Ro/JAtVMwfSKq
K5wfNJXBnCQ9H3oKCvLLyyT8V7dgdYQSNxc8BeT8r+1JvtIKJ61t6pGjP1eRD3RF
r7PY4JybUvDbu+AOBRJ2UBKA7UWPuS63b75LhwbbgJ3HpaO8O0R7t7FPP+rgIL7d
OShG5WTNIVsv23FJV50zNkpKWl0b/Ou0uB37uC2U9aERAga6I5CGrHDlbfDc9a+K
FYCCVDNo+/h/3nywr4fp7UwCGLyGGUHPDD+N+YOKDGuplvaMlRgfI4gbLykQ6ZWN
KhCdJMuotOQgj4xPGepOGnVNMlL/wEevE0NOcqb9oWJ028NrUjkgmBvkDeHRdTNI
WiJiGusSnlB8ew/usLnPL17DpQjN/YI9B0KDyJIYtvIHwm7JVhmoFstXAstXHVJQ
LfzSc2SSGl2B/i6XO0IUdtO7W+4opA9RUJDelfhjGZNWs4JBxmIx1F3SIm49J9Gr
GIIPPnnD1r9wUkyDdHfZZ5Gq33+RI937HBxBnUUiXWbJEiOuLhHTKjmO7522fSls
oNglKTOsAVj+1Mqs1cO9zKSfSx0mkNpsvUE8+XgrQRh2pIW6XxNmycLo3NRwO/WQ
Zbf8iI/okUpK048Bg1ow2FufYqSbQxldzixbkQhLFvdszIE8iEYHPWlkCg+mz7Gx
b3oHZecYCtKfuUjTzxJ74BjWdj5V3zIrIi3Nc1WMniBKm5JbUSpnkslDLPGqzy86
2Aa3DMJk6Wl3cu3zlFpser/I2pgUDEpOu9Ppwen/B/FsEWNQ75JvpJdldubVBoLl
QfqK2pOuekyP/lB6fFhtvLYadqQyUp9vSRS62AfUsH70MV0JblaVGpM8h00dOnsr
uU/OW9gILK0I+jl4gKT3fHirlWJI6QSRROCauByR59uvZHW/Z20dw3wbsNHE1Ul9
IoaT2037g5fYiVHH0CNOtqlG4soSxFtxaLTxIsw9ZjpOeiiHa42vXM0FR9q23cX6
MUvhL5av0CsaIJYmYA+ogYD/kEulzjDOFZ2DpcexSSExJgLmUb4Vr2+Tb7Pujjgd
V+nny3/BlU5AlW4m8UqMZ84gTX/n+UGF4b1lCiFfpxh0N28V9sHACDhKSBvA3DaV
vkzCnAf9EzAxrHC5LWEDv0hoBSF1Kmona+Sb2MwfA0ofaw7Ljykdw/FVy+EiIJ4T
3yf16s5sWugTXubQh6Jwnzk9KfKxnQAa1043AEF/Y7hSJPWS01tKpRv7X/99oqly
4hIAyQMeUzUGaNuwWqZ4iMYLVLfoAf7w20ErUyT+YIzcSm29VF6KLgq2PPfIgls5
aiUygpe1gPyYNoPVSBojWt/ZILK3s7JYUmFcemPBhwyNDUQrRfSBZ6HuWpFCEDSs
fnxv+ds8e0/sQ27Lxq46aOw2puJ0sBS/mJVAMdf8a7r/l1LsK2y7Amfz9XFlrSdT
QfENO8oPouoY4qzamjAuHXXWIP9Wus9MYEruLR7OoSlwM1D1CjRi702XWjGK0nfM
IlUzcBRxfcwV7o2zIkBfTWYwfNPLkZbr6IhlfKt6R57j8cFM4SJyhzm29mBfCFcN
5Z06eBcoI/D4qlUP1ynsPkQJiQtJFr0UBGklOP4L7W/RtuWqNrAuElnTFofWdGh/
cPEDkY5dN4TYgQAya+7hncuj8wIpLAvBuYPpKbiTpLauQe6lhCr+ix1Epge/8iDd
W8XX7zoQHLnqigrl+OpRAaQSlgSUhGusfcE4qe89X2oTR7GgpGVOCSttUXyxno2/
2omB6MRUNFhFi2FH0w48c07tSTSwI+4M9Kj19r6BX1sSK6kQbOSWoAaqy2qfy4pv
BoZ1AB+wVR8wGkjIklORRsFbIE7M6kRWFcIt4sCgmtOtSusSmiRMqADcieOBLPRe
BegVxIFM6hjJ0/ib29b14wlo+uVMGSMX4OcEJCTeASNyW0qVNhskhak1zitJUXw5
gElJ7soCF3S4l+bhLdUVSuV0vcS75dCt5Zc+ytW33vAcZk2QivH805KXedMzsh9W
MH1UA3B7o7H8KWXZQqKD82RCOhzpVoS1YNM5nJK7jOkAM3PtyFHTuFEc8MS+svlX
tDh4NSarFM/dS68ylH+U94pOlbhRoE1VAk14hqfsOYhmrtOCXVpdMBtJVfbr3x+y
9FsFZh8u25uQYmkrNnwEEh+4ffU+LxsYo2Arf5fYseOejTt45xv4un02h/dRO/Z1
aOH84qxE8V3/gsYnyjBuePP/1CtA8NfdwjdLCRiOg+RxLq5CKBQtnfetcHgAd/+a
351V6vs+sIsFuK2wQ2OOJZ5RGyCz3JT5CmM34GXLB31UAl66H3BxEdqtQ74yeJEr
FE7+87OagTJwt3gEoVebMLqXgRqVwKPytITG0Phl4QoX3W/HtZ0j4HuKZDiK1PXO
MbJDCRumqqOAwD/7KI0xiFHvjiJiP9VHgSrkJNuTPL/2H+FmvAjW27QGelTiioV+
2bsckxOZNA+8/7Pd7Aqyn7d3+Xl/JCDsNQVUzdtA96rP5Rgfm6myvCQYfAYE/mpy
HLmhDvhnj0FLOT6Par2T1IfWk6ZxMO7owiCborWjrgVrPeL5gWmjg3bzQaqiGQ41
dIovL9ec+q2FsfuAjJyJ0EnxY7njgyumsVfBsL0KIRV3jJ/jK91PGqyEpmuaUXdJ
WR81Kc+DWiD/6YA5awBSSWy1Ec9PSB5NHXNXlxhuZCC29yjS6RUZzOjDopMyF6Ga
KucYybpCxK8fIe0m273/Iw04sgSZ3A2A75lxzoxGuMWalk/xav334WvcKrKnRmhB
N8X5+Z8JfrnivahiJQF/WTFb1DNEm9ZTrXxwMlUEe0YgV7hv8Uy5KRuO55sKtGfX
+TtfS6EXM8cfcyCafx5RKs9C9kw7dsRZJgZCH7RXwm55EJNMi2PE/O1VUqC7yJpI
Lm0qSsHc2ryI/sSnbx3XzIChKiGt4I9vebb/RTAhbB2Kv6DngJOWUfS1Nb0hr6ok
psgJC/LFxukUBzMTjD38YQekV7+p+82H7F7Of5vahiK+w7Xy+Tp8XRoPfUFkDf5z
mOFyC6hrYfUPN9vAAWE7jR+1QcwoBWs63OxBA7G3buD7AKQKzi6BYRCG/XHpv762
4+6OfOuINT7tcEZ8+s1B1gmXkvOKvMA5jDtckptU9XRi73j3pV63fOS8uPsFsyYE
Z3hkdbs5OKqxg21x63+T5w9Y54dzrsh9Ixv98FeiuYAlKjAbbLL61iVvxVykb33b
35TNYtMiRQdYwfkzR0CMkfoBPMScRVHCWOOEGf0MaRmg3z70fz9656OQbgX7AJe7
QrtZdJaF53PQyd7fp+X5tNQijPJL+PKTdysls0VuBmPW8ezmYQzzSWxeKdv6RB5v
aoChGoP3Z+UAvVE0Xo5A/4JYe8JpfKqAK9elIGVGpx7psOpRdRiMM7Cykv3c7KPL
KZM92MLMuNVVLAm2y6pzOX4zozlZvul4YcaOd5a/CscUlioECRr2kNFJwV05uBEM
MVFhqL5nM1ReVLDAPq/X4pIWaBlBigvXX+4Q02e4cusHoi9vHp6WB5+sz7h09LUQ
Haz5EqJNoONCVYhldSfPBU7hzKIk8BVcLZFkhkffH8cuUzscBpKWnbe/zguU7PS0
KZfvLFgnPrNjfSopaUiblIsLRsKfal+EzPZVjlazEDAzZHlggSORsyDXmweJyg9Q
KOWAYdQxz4sW7xUgKU3LIkm+MItlOH15cmEB47mRPNg9+9NErC1PmH/Oj1LnTjGI
CxM05zBIuayAGO7ow2znActG8Jx+On6DJQNZ/e8WZ2ZFu6QGTFEEDa9gL2JqRmbw
dFHHxX+UJCQpVSG6MkADwWOPxUK52O7kxdArTmnA+hhtglIQWCDXPn4fBLI/cNKe
GfKoaV6SqAjyw5xTJKVEjljBXy89M+V6KSA0/sM+vwPIrjQzVDRDv9zT5u8D4V4t
cWmRFHk9Sf83VdOyjLSaELfQC8fAcoZFYsUnYtGLDmjGZ2nY3iVfoz9nDU3Kk6el
+uNfg5fnxhXNYrczyp2FvuZYcM1N0IkJfZcI7MTSVL2ihmP7zzyzSYLz46dBPtI0
s8c+13BpbZM49uL7oCMKMKvDODT1n8ffgOK4fks49vaLeGVSzOmbESjQCkrKlUK2
eFb2j1awJnMq0UVbfMhri+T6OZjHybZ2UwmgHVYdninqI2BwNkgBlcDoo4EvNYsV
ZuTRayNa37ih/gzKStIej2EO4YSEyssUoCCmzt5R6ih5WpdSUcyIY0Ru3rS64/q8
L2UXVaQ1doV4sYW2M4BP+MBFx/GhIl61AD+bxnXvVhUmC19lktMPOuZY0WzIT5oG
73fizIxKckxG7nfigxW1HMZYOSOcF1mu0ShppTmvmJzEa19mF4Jpqz26bCWtB8nk
FR6kERxQptayMHMgQF0X4My70cZrW1kPMJsxEzs4wfDgi+g/ADPXjlGqhQMtRP4p
o4qidcrh28i9Oy46k66u6Gj06KXm75eBcxOFK7QL2bmMnxgP9c/C6PMVsNHDUGwn
lJ8VLPg6JGHlYjuYTa82tg/J1s40yrCGKqDH2GdseRZqlnK3fjK98D+v06QBOo+1
yJSPN0vSfiPC4dXfndrQ7IJhTF+WwXuWF0+b9pE91drqXGDnB0RULWQqzsSCi/a7
rN0lRKxzhiBsGs6kOMHpPTdd3FSRGp1OSlLpgqDY/RL5fxpQnlAJcbC1Mlun32VZ
yUcJziDL6O4wBbdy+4hCeFmmutaMF1pm/1rEY2JrQPhRXh/xnSqBNuK+TLD/sjRj
YSwc2EbhN0qOSQZdlKgwujq4y9pHY6ZHpGvCqYAuQhkFtBfEtW7YWL9ka4sUii2l
iBnCIo7cI87Pd2jDGkVme0I2hzYujxr7tHf3Y4sglDTLs6jyHKFESZz9lxhbzdo1
QMG/O73M8u1VHNycjhQsAl42qs/4Kbo51gGLrgLHTYC0HQyOsQH0JIesZd+Ji5wX
DddVSd4gF1WKjIYFCvPIUZUaQC9jwYwshdr3lP1ix2USvK8NEdftMoKFpTDahuLo
1JdRFiLg5vQfr4Ekuns62ZFC2HDLNOivyGArT8FisgRkRA17tTbivDRmXGFwMur4
1ucSNqb2lgKZsJimk3gc+OI1ROWf/VAtehxpy6TnKcj6BIClaI2DxHcZW2WG2Jkn
fEeSsKpfF9WaXM7Mt+l0xc5yWcp8E06cq9bnzvat4i1wggYMjuznp/Xwh5vJRziq
bVZzceBWz6RNRcP+FS5fKSbnpC0jHyeoEsY/x7lh/iId2gM3212QvGiBYfXwzMHE
5+ZDpOAis5kdUqdHRdCMW1nohMIqjBT/JRNE/0aEirzIlVQa8WAvjJ6ZZwgM0A+A
COumleb+qgW2mKi2Ikb19aYorTgSMUlG9tijckzgLBl46ivQlrHJM9PDJcp/YceO
eLe2Egsg1CBO2z6juVFfiURwPHfQAAxhOAUMSUVNEnhIF/PHJCwDJa/EdgFjoPxA
Gi2S/gasP9oWxUUR3fyOSQq8wXYeHQ7F0FNX9b2AWMjcE3mVOOBZkkgWDLr8s3yC
N1SIOvrB3w0aulufTdacjPMOcb3fgQh//UQc+83yWUe/tOfHPek+ZEOY/aLXn2qr
oaOJfkeymspdZkA6FO3zzb4WRBQ0pgSHiR24wfPQi1l9ZOuA4zKvcpbtkxqEP/Y3
YifpbEg1Gz7/bHpBBBxM0QSf1iL5GZgaaihC1sEiTngtEjGL17KpsZwzcxj5iFwm
3+0tlEIFzAbGpWuln+nkb3011wIeLVvHDDlvAmpZ9V/BigOiZNeszbuFlGPqjyFq
OHJc9Lnb6uVG8aDhf6fJ14vyTbQjWshtyyUpDPRhBcJdREM1bIWnkQIxh0F9Ctcz
WJBO0xNn26JFpX4IqP/x+9EReIWr2Ja1yPE5OmZxO8u0rruQx57A1xXQhmCmFlh7
V8q+aPijCDVMEBQOk2TvtRZVy/TMneEVnV9phfA72FwwU8qT1HqGkHgY3wxWpAOE
rFmASJWpFwJoc8hFR/Ti04jgq6YGiU2m81O+JPYXYIvoIHfrQyV8lAJ+WWAhsZZ0
AV0DnhAVM3+aLj+u1asG36Us/QyNAfohQTjHpX5SBqQbzi7vSeliDqjB2NUW08Q3
gA3RemqbRKBOWbc0oeF5/19Q/9TRoBzGhzJKX4a2417ofkpMX5VfjU0LNPmTK8r7
f/d42Qx3poGyCKrx1yvh4ZZvXCcajoFL/+fgU0CxHS6rxb13vXoZcLI2VEjslajn
3GahEFe4KV4G5o3XoqlnD/6me0Ct998B8Q4Jkwbnrf3HhB9a1ztUgK49XBYVYGyr
FMof06j2+i6lm68JP7h6Kb8PL+pVifVOAGKw4g506l5Fmb1dso3x+c7SFfT3wp0c
DCifvkzKCf64I++HD2lJ8CqhMfuglzeibPCVtrHkF5sSwtPlrdbKCyL6LnPcVNqE
O/c1PYdnUB7im7xazo1tWRKe6v4WcuRCgiGkkz081dLuneK5ARYddwSfoTY/f3Uw
IQt1MP4PtbPHCqfNjt98q3x65SgOfDQdN4rk2mP0GUYcXCQyjss0FJa3g5o+I3w0
jbS8zJtyZZbGCPQOG4IsH+PXyZCOn8ees3dHLfDc0og0U4rmsfhNnn4ilfHlSWnk
UR7us7T/ZFc/mPZTCPM0xf1WBTPn5Qq91fA0m8vtNDoMObYjvtU8NfVOvO/EHs/O
6VHnG6hrJKd7Mai/8eW7tCibyvIu70tiAjP+TbSpRzHDeZ2Kqkzo4PvO0+a8/Q1s
LCkndmVW/EyAqUVPodmUgXBrFgV4hAU4J2Q6n/EhOSzjzIicOd7UtX4X5iGB+Z+U
qlMgqwIYp+auct1LevDxmqqxUVp34nQ27DiYHVN2UD3MkMO0ivyKvImYn2gL/92D
473/FjCGJ9MD5C5rBPEENaOPgXv0JeNNlNg77wMtc8zxXHdAC+kmeqGshGPE1MSm
4OZxmlM2ocLUjkhEH+Rvw2O74AZXbV5/cQJVNui7k/fcf07sJt9NYGP9/ma8Po3n
K+nTCQGvvKZHDcrdibE8VUsa97EIuJgui5jyq9FOB/bryRrnxckZtOcYFrnOAKue
gQbFgncuqiMgO8POWtZEMTosYyP4UXZIS0RJyoKnyPEH6tkkPA2sPifh/m+QVTYt
BCXje+PgCVK91BFyZj9fovKBxX/bWc1E03RT4eUTSOx610VCmiKWWmiqr1+9jpzD
uOVbq8/qTEx1aK+4nE/a6onQt5BfNQ/+v2WW9mgj3gTQiPG80MNt94YvFm7BOpEr
nrYvzZ8KpxC0c48gjusrl1ajNprifxQL+khkoiBzTOXjksl5amb/3ksKGKOPZnxq
CV1Qr86J1HXq4h5WNTGhTg6QL47u0OJ2TG65+grZi52omcbonxp6Ek/6NJwTzG3J
iv7lUhqa04AV9GnRcc8IdP8p/Jb5qdCB+eSgzLEmOqYHof28fS3j++XeyOz9wfDH
S5s8A5KTo7YmmH8z7UnxA69raE9kVtBX6sjZdKSKAQw/SRuNoqt7E/s8D9s1EgJS
jk6U9KGRG7jlG2jm23HQ0R1irkihANyy+N9JsZtZZm5lBzimnRI5pJl+8Qj/aWPA
s7GSYE2D004MoDlHnK896la76QBP+jq5LqycsXd+HXTLa97/6HHQNCG5A0Nh3fVk
wPY7F3Z47Afb8jjhc1HisfxZEZfqfFviZ09ECpulVCNZoUij6Dyu0LFvoKZnerSo
MRnBTyqoY6arNW45fQ563mEai7rBUy9tP/NExizRJa3EiravhNyA0lRy3cBJnR53
/F9BAr1I6AXICd90bRN1BaxV7COYHS9e4TrEn+BEwSmKLvgZvMnX5l6WZevFEeec
AG69YfnlPK9582aVb38vFQMaVaM+AlJJahgcOC62E46vPgBSC1+XqZ3dqfa+bv24
bRXd1EkJlEpozSEaoDAT9soKXX6cEW7qMqZBQxLJePzu0JtaDj0UYE4jcGblL1Gs
Mg7cM2d/BWOvE5/EvhuD88cpFjhAM2mTONfTxT5Rznu9vYQcHwyZyI7Qjt+7VR5M
rjaam2RRTUUjIrPALd+1SnEoCfkO4ndoGJ6MjsGrJ3K6G8XrM0hhJG+Kc4v2zb4a
sZFGDUA4JGHoVA3oIPn5Mzu0jMpGBT1XwXcPFR7ONNjEoMit5gcuwejC3A4sYV/W
gdN0UJ7WmcHfI2M/gVcrv2/0uerjrOX25BOeC7iVRh7DLro5d81NR6obJyhSH1QN
fYuqsDhFrs6TqHJsIOwecXeEGAC4EhzJ+rDmkaDr9VhCRaQpqIJfOCVzIx3KU01U
+cN+MXd+3pUQhT2uML4nRhX3CQwpoaTZI5e83Zo+O8TzGslIRIhunqkG2scLhOV6
cluDM+4F6YTDl9tdw41EURxiopuCfSLlmUGo2Sk8tEW8qgTuJAqep64i86tsMa+B
bNAxW2Vh369QZwunBiSf1wE1vN3p3GbSIfznLl1EvH44TgVyZxM4cQmYXgmmjEoK
RVbQs6MyZVaXOJHs1hbgK9+2Lx/EhzG7yfY6WmspGyRo7I6iAlv8UPkeJtVQ2sQk
MsWDKl4bnTIf+pkMTRHXVlYRFWvsaZQocNDULlRcZ01TD2ZOGMeOLdK+MbKJyIl5
0DS/cZGntrE6sHh5zbgTM+l+O0NKF/Ro0eZcJPekR6yGB8UhMzatXvLMFRZXcjDD
Ty4V6gEPHD4twyBjNblyB8oPmJTrtQA8AU9W55h0TRkVqVGYC0byaraWHBojY1aQ
55+NR7+qzRUocE2/BFf4U56vOdb1BWN23J2dHN+9hn2nVGgbNNLoX3XvVyhNl3Wk
BBwt0LN2/euLwL1jETU9opIUV50/93atKbKyOWao5z4CSh9QBXKO8+/0PBpeJS8D
0CZMFez+Pcdc3HpjrgjJgHkOwazvnx1moEn9UtpO2bGUwuRu7+zsi3YqfV3AyDgk
9cv9QV/BTp3OkMsjFJhqA7eOiIQ6yk8OJZjWgrJ/uJcMtI9Q93oxeq1F6pq2PgPe
vpL07py17JYVkyDXLCoBpWQq3kZzfDZTS3d0YLo6K4cme22tVsFZTPEsGtwGQrn6
e5RTVGsqkrwrURuCY1jyjZ2MU8ct4vL4Od7u/wtq0RvYoU4x8P0NLrbA1tOxXIAw
sbbWWwN93IGmlXgCvJWQw2EPkr2nEVZIbqmkrVmB3SWeFsS9zMA2lYDuzbn/JTJe
7vxeOZ0nCnlWETXRrgM+WLen4Mx9LtG9hAtHRdxpAq0cdKrIrIrRDPOFiOXqKL3Y
eRkb4YMmKs8rQEvAshUrY7+ORBhUCYKvfaAiF107MqDFPUgQZs5Ulq8w0bZrVw8q
QMbIDX49R54gJg5DLqvuiP/9tAjcJoxy+8VaHL3WNwcm87k4LqmV+4NmwkQgYt/y
e1yLDLZGyjfF8zL05D+Cpm1YlesBorqwwkx7Toyq5eI1QAy/l7VEco+2+uZCobWi
Fgq5nwjLyaHLKnaimIhSIRdbgrnPJrVPYDXIRqRmfvMrxK2dOiIJu6BPLo1KOEFu
RwVAPmtSFN17A1b5CLer7qlcPBXQlb5+WmYpmZp8Cil9wbpeLpH4OtlCEkia+q/z
nPUUj8WxqbKdSAkyNHm5dGMx7Az2wfECDG8N6woOqgpsUjjScDIc/ZfDmixhqJDV
+d+qwTTS3fG0+uvPLT8qs0QZWTB35Mef3rsajo3xZ85fbVZdsyeZtU/wCP4VY1xO
e8EamstOG+YQjk9SPYrzPQck7biKC2vg76562BD7PZ1IjW4UTrqms0sFqNMMOpt6
JRdu6ZntJfp6BcBbydJgQ6+eA+nialzgrhvT9XqAN6U9pK7PKSVyB6NVIZZvWke4
6tO8Wpr/JKYIfy3gWRUvFM9fv58ihanEtzTwEvGwTn4vYBYudzbNfxoSkz66Fv5N
3rx02o0tEfn3CU7jquhbcFoV7YdFhmYl9i9mXhwnWBDi0L8ITbH/WLPuvB5X8M6D
x9h7W9PBYF/PXLFMZeLBepwFJixEo250M4jr7q2oIu5anPVAn0ia75wifF89M4oK
KJGIGvcc90nurvDUYuOiMwZWg+GDTY3b6JObVGlzQ7w8oZ3LxZi3qMwfOe+f25ih
qt5MtCMEge3AX2iIBQ7CqsPmZhO7DfIf64Z/W9zq5+gfC+SjvD77TjFyPrlM6kpl
02Dcv4jhh3CKEWHoTyYkm4XlyUhehYE8c9X8FRWsoA33qa+Pvp4lKZLZXpKW+i8G
vOW/gdOnf3xOfKu64zlqS4Y2YkGZDkbYfLZdzmMu4zin1Go74GLsHza1R3oKlPRB
VWm6Qq5o4C4BCPwASc+3KSraF/vG2JExfK1f+7/IkGa/RZyoaAk5qB3PZamCXZDf
cwYrQ0jP2Q/1KTkEhHWFuqIwu5zmWHaLKKqVdhpZ05ZbfHIyOArJwiVwQAuEXG3m
9Iu5xjNFzVOSYhwSIUYZyNRIKXfPqCa7GxOFJ/1Sz2ks8SJNuA/R+8CZnXfDbfi5
4r806ifzd4sskmttz1SqG4nSiYckTYXBbWHw5E4K8urCdZx3Mg8DGnJmPiZFQT/c
LKQV2qEC1KAUWWnroF03fdIImH6IMGAElVto2jvOlXsMPafwDasnIL7273eS0zpW
7FwedWQ0rJJwJzl99k2VbADQikPmXeBkfeimBUUshxPdhiCCoBpWBLi9m8KwvkLb
FBxMSbez7isxmQTQ2AlBmoS/uNSpwdvgo8uijGYGRqobzbBLVcUJ6xfqMSRUzMEo
8Lhb9BHYj/ixJOtT2weySibdoqbBpAtkDj81Gx9rEQUubL/1cfYqxPd1ZMOogfy4
IZMZeu1vsV2QAhOHSEPLsiOZNe/trLyGGUKXxH6nPca5eparPO35e6F82QN5VNRX
2/M0dkOW0GZsTZXZoqZdR2WctF/+b42xNEhKxs0HRp0ubZ4vVvweQExvOCUDw4Iv
10CI94k+DTagTJlh4dkjB60c57EY75ABWKZbBqdXw5JpqL8hKHc/TX2BJJzrqfLd
iAxcdBeSnLRQ5idZZTJsa3wEIruzgzK4WvWtbLeCzGVtzWaoRjNNBycICpxxWlk2
p8+qBnrRBAyjg3blg+nBN9lMPn4YJ1R+ek5FKDpK9vM2l91+VIEn+u76/GmcrMck
26rTo5QC74mr/FHjpH1H9itW2Hlzs8yXXQrkyJviUp7E5Y18O+/VNwCW9xaEe0AZ
T3370yNiHqH1d+W+14lvOrIUvxp7/nponc1L6sVpVDAC6OXAziBozhFc4aFT+ss6
fCZGGsTnLStl2XLsnD0wZ3TaqEJ7GTnIVkGTm1915HUR8HsUs8vuytRX1AOKLde0
GHjjSFdSH4AhLywGiPRVC2/I4+kglIhoZ6flgNIOcDALUPpUppwZ001YSCFQXQx/
5oJTHV5fE2bZgmxNDHikIqDnv7KbGeAyMlBEe7lDQydHJbZysK19xkuYni4I69nv
OAI4COgSVTdYBA8PszllWCVpnV4wo238rmfTu0DZ0wlTRHHAALf+sLrJhSOLWzhk
Pj3zr+ypO5zYac0sJut3LVBfcmqBcSgHZcDquYfH6kiKWv5eO1qsPSf5VywVpwjB
YkiEuZcXKNpvHVn2PkyvCbWI1I/N2PZZudorVZ0NQjo/wEVsn83tFe7Jl7+w8ntF
p2qBPCqsnrMJMNxhLfZWkMGJ3kkOcRfwApJfj1i+Z/fwxx6JLP3qSfJZ7VCQVdCY
W3edRY7yfdQk091MbaDw0iwThiVJerLP2bH/tigTd4SMzCGiRegPsBNVoMpnlwam
QFgHUWnfTj+OKEbr+zVfze6n/TC1/h6IHrV2mVXd8vhH2XHET2EbbFZ/lGHJh0Qx
ONdT+AYbBxjLuJEVHR+XABPflZq/e88lEMxtDeq5fShP06yY4js5uYPBEtXTy/CM
kGLU3yOvN6gAsqO4xaoWFzr5ZrLnntKq5xWlRK+qpCp5YBEjRDIqumZi/KXjijMt
xBzg53QtyqJb1sSHPFvjxkGWO5UHPVViuXINNK5PU/GsK0s0UtxngXdLa1eIBHm1
YH6cROuaHeAHEUwiGPXnexjObp1inI8vzVBC5rMaYD9C6mK3tmbbaKfyXAIec7HO
YJ1G+Oli2os/uBrVKESPA3Yem+QCDomN5EjEyYh3f/1nWd8QlezQor6xCEBM3N8y
7xnv64G+MxfuoBJQkl0Ag30MKjnKj5u/YG42tzehm31PSoe+fB/HQ797jfqJQhjq
nW1Wy0DkUIf/VrrQEmeg0N0wQKyoxO3Zwbc3XwtO2qaJm8HsAoUt3J6oTOppZ6TT
/e/NzX28lDEapEKIM9Y0PxT78pQpEc+KS7HcUIA6c6A5fIE8KXJdCiOmcbxapCnV
dCF1HNfyKH8EPZPM9BZ4xebhgDtxOqlurblE2HvBrLJ3SxXfTT+K5Ttem23rTqzG
m2vGTC7h+49rbs2pnnmR71W8xVwwXomcT36LeeKoUFlbi3xcIYITWURIuAP5DTF9
8+sMJ2flDbZ7lljU3ZaWw4S84xpN+kdemCxQ0Ia45d4h+gzFgJnzgnEZvtD+zccj
JiNrZ08DDGq+T/c8zX7fE0Dvc/zHnhje5MYmVjgZVnt6u8e8FyXvoAdDSrrSPo/4
NEqkEgQJdvkRN3WNYZ4BStUfluMF6zJKwiKqvfHj/Wt/o+NgUNxvVR1fGd0txVWZ
DLpxyHoilJiV1d4fNxjD4dShkufz6wjODEku1mwkR25QAaVY6Q82i10nXcaJyK7S
NWcUuqXYbbLqXCuhZ1uYOLPPfHnTAj90KOcz20HQeYG4xaxqWvYOCgOMW5pIqr+5
mDIGG3SS+F+VwkOi33yiPAGohvdfAIHAeeZ0iRyO4aFjdgrlPTCNMgqPY4ee86al
CMfsOVskpz7Ox8ROzOA8pryS1xcbFgPHpS2fKMqnQxdJYbFQyAogtwo2YOJyBqBU
BQd87JGcrjRfyxu1Lt1zNGtZ3vyf2lKEaSOuT0/GcWmhFSG6SICggiX8Xi5WE89Y
MhoMwSPOBhUXue3bjAxh0n1wo6lXTW0X26/msFNZUaaUQk6v6QOQuws0CGrK8w8C
AQhAlcTV4OaXivxi7Q/AtKFr2xzeuobMBONsVZPeaZ3czYLBAXTjMydfjjrGQ+vB
iLhO8kvS2OOlAKeOZQiXxMInpFyRwvw9q98aI500FbHweP2pWqmI2fMAR5JU/WfP
Bn7W8kFVt1KdppALBN7W4BsgsW+qDe9TG25I6anOjG3RDNi2X9mhN3gH1iYK0mDl
hWdGwL/CiFFuF8aACDehcuPhIdgMKE7xctDmVS3FfROAzHRqHjsyd6ujfQngvfJU
A1iR/9Rw8ukUwg9fDdZblpfPVylqpKEhZz5WxwWsC3T2hFX9d97zkflAmq89C//S
d4oW6ghPj8vp7HpvOjyJ7ugewetZ3Ts3kYenBdRBM/sNwSTCx6OiMlowH0Z8XWMK
4bhTPkz3Q9B3eMp7Jqdgh9a/Ms4AAduei2kXpcJ+oUzQ2IP5IQKDd5EtlRxC+E7H
F2or5SnbVr0IAO4/dRRm44yOObE5XVK2Bx+MhKYErotx+OxiwvK+CUyRW2z58/ce
C01p6eTFNj//kWp7FyvomFbg0g8z3zQY3CJ4TDKTSAQT/LU0PCllW1aUDau8Drz/
CtBRCAEHnAUi1i7Ef/+lzVdWMO4Iubv3m7IFTIEN4Ca2TdfifKFVBaYPzkyjGXWt
C/vo8NO2cqXgYZuPuPJxB6ES+MZMh1w9NsJP2xCuVqGhp17vUiEvHHxF+fcdPnfC
gfNpWYYswbKvkmZzCwoq0q/AZBIEa7WutfrTHE43fEu5bdZZFRvIbA0YNqoR1Udb
abMBg/mKh47UiCWPQvz3v8fvPPw6Lel5dKRfrlcf0TbSovamTXHTQRVEAhQ9OfRy
++XZGaAU1CHXWEbADe+EHOL5X7OYxvqVe1CFDyL27Eu7rW/IDnO6Fr9kdj5HDWk9
0aZkXhIhbQzUn6ATmZfzhAy/Kq89yxhWkMFuVp6LanFTUZMwlmk/rZt8//gtf9fq
2hX6DTAR6fwCVGBNKJnEGYo/SfHfHzRqFPQdbw3v2hdsqxDeNc+agy5g+TK4u2cr
c8eoNLRFyHihgOHCmLqwM4UqcQnN5ZP5RUT23vUPYXGGqxPcMxPeuQejza3xSQIO
OJ+aoOW7ZwXRaymMXxpEh4XzsBfgtv7jCJGTJsnerpZejP1+yCyAO3xYhZa97uSP
u8Sufyk6VL/98fF8a4ug/NfGiUmjojoyktkoXyQgsLGisTnsb6FXgiHWpsNyUyx+
F/Z1fSBeLaMDfvt00XFEYxSwvCQLKSpKILA+Tu1ENSAy8PGG8QJ0KOQjvz0zZiol
+5IK2WufNBO6QpljwypNONgX70JLGTb/3i96wH1urSrd4BkAPxOD33n7b698sYn7
rwnqdRCH8XzqGqDbfknXNXGMHS239hrRa+lFxyflPlWsGVafNZDcJOfOnXufdX48
UjAdMJ9nyviQboBspziyPwES6UlvesYOgB4f9cEoeZ9/6npQEgoH7TeU1dBnsAdv
am7bpLHXR6YuxyOHJSo93SOpWtN3S+cm0qhR8VcM5t15pu/dirkKUHSYXt5zXtU2
5SvjiYxjHCTyZ8RdZgdllPpEPS23Gw7KndsNnq3ftj+dzEk4EvVAJfhhzqc72DKy
0LvugP3QGJTxAuYebNQxNOmnm5RZiHdq6n0HEEQ6T1Lj+ul6Q4wiaWE8EzWlVIXp
49SIq7J9rqbFr1aeuc+Xcxov9bszDdkYmWxOpwoei6SDTOx1TeD2c0el8o7KQDra
rsIYjDxBdR1xz/+bHgb1X4Q/CpG8idIlXRWw/YEVqmC0rouPkQGFokTkONX269h9
n/rhLxvkzTDK+2J9Y8Cs3yivakIZSkNJcCY6LAxqSx4JrP7Z5uvwI0p0AoKqoXL7
5QbGPrp97uL9uc472MHYPvCOIJf2c7ksVsu0XGro/TxmKmFaGqLN6c7Sf2BJmV0z
qGqlmRORL5LdT8YBOqzgmWUxZorWfg7D6+A5PS2QHNUR273uGi8ChmOzJ+BIXzPX
M/N+56s1Fm4XJmAuZBXoL2CLfFSzLAWpHODwAMEKXlopOGkeRB1zi570OoDZreEI
2qEkfFi9pGUV4/qai+Q/bfeR6SzJ5tMdugqLeMIIkF7l6EF2WaP2yPj5MJ5LkYLX
XdbgKMkFJmYhM1ZOoypHn6mg0AURnO/vQiDeJipzHJswBzRpEHrsHYoD+VYMOaJZ
9VoW0yHKBywgsN7sVG7/aORaNCS9vUSzBCcopq5R5j0pics0PMBQN38Ds54BXiwC
/cOgy1PLFEfhUOT/Avi3o2pDtCnBWAN6U+3t3wB3B9mYUnRcjzXNaT7FvLaV5OXl
0ql6UVREAUGaY0x7G/3XV0UnTPx8Mo9uVBrNBdIZPDkAD/WRUe4lHqRN2xNfWl8t
J7XNcj+qGn5X31nHeU4JlsHqGha34O1shgJpKe38Qbt28kbVJRoLkdoAebmIV1BW
n0NLmlWglDAaex3CUkUsoaEn1f6eNfWkJwXtD8qedfPTSpOBecVZYNESiGCap08F
4cGB5I+tRneQqvSBrucYRv8flFdndJ6aRsCQo12CGWvOndhex10zk0EPMkEYtXiS
CHJT0Wj/vQZnYiyj/pLLr7YpxvmuHIAgXdOp19bgQV/0I1ejhZFUMtNlCkmZXVA9
b0LghedOSY3SLVGxqqgaDTAQFozP2ZZauYCaSaYTbUhStVZJtPQb5KD3s49mjYhp
5JQeph1PfOospD9L+M7/afRPKz8E7UDBFWZMTtwN2jEQWIiKBRJyaffTMPLiDOKx
Gh1da9l0HNlzttPNTewoA8X9RwoVmnugn5IRXtERgOtY12MExMUf1v8TAguZ6Q+Y
Cc9IGJ4U7mT5VJUpbXxP4I3KEgLAQp9LJzrz6875iP2N+2a5irbHOAs3l9J5y/eI
9qeho+n6sZ208CnBnBzZHGuDLTaX4E+7mrkyPSIlEhdxPu1FupwW5PBnaNuLG3jR
iJhSgZXyIHcn5QJBE5eh9wg4bc8Sgt7HHe6+VvOP0ylx58Sa3loHwSlsH5PQeC1Y
0eb5F2ML1bLE8HqdFt0ZGkdmzIS5bVEzPa8aDYC6sqYESpeu3SbGD26gtRaYg+ly
757adVcKXGy5YY6HAoePIco9xoyfP80sKam8Ymzxl7mvDIlx1XETbjRjQYgnO9Bt
LX0Bgrjdutz/kyztmyxb/GHSvjsYhen2mTk6sAcV90FQ/O1JIc4EqvvNqyTd1RxR
qEpVGxI+Vh8XLDTT6WoEh+LPy+creILWTtkhYeeGzSHYjMfcPaNmhV0st39pSX6M
YZuGDY4VP5/G/nhZMuZboB/TOD3miGh2bSH876hjlS6GQh4Tfr+w9Lv6T0oRK6mj
XuTM1fYvqwziZmgc3Io8glVrCUUz5Icvv7PAmMyc9peBZsnSwffjyWmYAi5jKWmE
r1pEyyKmBc9e41RUvgcCwd0L732mGIr4sJ+oEDrP19a6GFRXgdyYppGEy49MzNj1
txNy8RTe/VdXhIMsRVQvHCAYxpsA2bryGzFWqGMDcQJrGQvnhFwKPM/8n2wpgs0n
cLrvKDIMidZEkv8qXDaDVhF4jhCYOPkwOV8uxjZYVSfn+2/05o818n89at39LRUZ
wv+f/IdBli0pvO8FXSKr0Co6KhKz1Ww+MnLs3QGXBbiqk7HU2NG30n20yBGLr9Pv
9GYvFz3LBJIOolqJ9M8ydaL3yNrhvRfjLChR76xOhnzbRMOEY1XkdVPpdlgvU70s
d4u6g7bBEkFpD4SchL+cCyqzLHyf5cXHRgg+qHM3SU/MU7TgJaGcnXuF9xo5CXS/
kkGDo+MVK3W6A2/Tfnl/w27kqACxdQY73FQCYEXV2xuSxg6DhJpwsmX4y5jvF5Ko
Jucbu+vzRqMOepHQHEo2Uzco/LOy4mVRBT4ofRmQ8Q40eluPbfo2Axt/WM6RV6ZF
x6EZh4YNuKcWIRs3ZkMgPiT49KH3Z0X2y7AaP6VUPEPva7gNHatZERZNEgThpZ/5
SixCKpo9it5Mh/GuEsJkRlZaZk9ldbZkRQ5Q6Sf1lebTMcWx4Y1hcn67AzuQMokp
MELUDTbWoLh9sZRCy17fXDELt8bb+4epYeuKSvwoKPSXDw2aHx5mnDfFeYeN+BVv
BymClKOHpaV4Vf6BbEMZcRQAsDEleYSMROyruM+ZvN8N8qMQXAFnw+4EARJcW7lG
yaRMhG46AFlUspNpLW81qyWDI6bFHmCEymP/rUHkDPfGl19+1Y73G+aOK3qzhGQ1
KKeRHa4hSZdFxSHlz/txfIhnAVvnmbpCR+QhvP7MHJmWkP0Pp8pjBxXpAfr0lVfN
n3powJ8QTAxCJIm8e1pNhwKWKl4OkM1psed/maaUP9FqHYPH9kjE+Ub05FFIV9+2
Hl1glVxnGaVii0JIu53r8ZwVoazn7UbYWdJT5dTetp0GkkILbQbOVP0lYKRVZpX1
ZsdPym+4Ew5BjocjP1a8PTCEvaRw8vLanxufRlEwNgbONAnbS4nv2b44nLjHWpM9
IlN1d/fGEqrTmUYLinKYraVMO958qLph60s5B8tauWNVzukJX3l5Mni8QdETXp27
xMH34+e7GM6TPbFRSLG9zsQQmx5TCWWLuHx6iVOFa9I3dx4k/K4LXddn+NMOkLd3
uqBgK7yUZAFo5rlSvDMwqYoyx0JyeFQ/qM7B+WAAksl3T+5LWIxByXsRW2HfTefj
L0DBoLqElAsaOCwf4RW9z5bO/k9xuI1fYOoFU557sbm+0K7Y2GIVZM/R2WmXuOrq
oNSSFgHKqPihlj3coPaEvIxAMPmZBjThHGrymYGCR+3Hlve+pD/GTD1xHmqK5WeQ
F9BnhrZC+9p4s8dcIu2q8jrQyT27XCm2w5tP0bMemr1KxLjWSG4G/4Hb1oykQt9Y
KFdXOrqBaAQwzjKXDN8WZos4jvMtyOkBEEZG08TQ99YaaMYTQPq0+m2xCAQtJoXj
tGITVuFKuTmthw093/yH15KAVbr5Nx7iXJ9d4odGoOfnyIraTQ7lEwZ3/NI3K+3Q
7TImooBlUglm53GXrJw+zbJ/pwDOJf8fln//9NtlqGkY7f4QkiXFtWpbXXoAuQj5
TGUBUmJJdPOah72HZYfVCZ0l0Ck/4gUzUKLwChhS0QGJdZCcXRfVCVhOKwLpn6LD
Gkdvn/FZPyiGPA9pYiCM3w/BTHBAHGK/MSn+TH0xY2euWZm33FdwWuZcOFqluP/x
jTT2qwbEHuidqL+2RDVIyPXf/NTQmxqqdlIQqk01Fy0x2+giYwewkbUDX9mfgGXR
iuji4DoxzaMNd0e8gmcQb9/FZ0WJZk8Oljq/2wTvMZc/NbZwmWKOF73NKOgo+L/A
X1iUY+o2+aTxKooTokNJXB1L7fgMnG+fq6UBjn9J6DUBrCbp3kAUFeE23m286EAb
zB/IsKFNlT4AM31L4ynWc0EAh7+MlSmVuDeIe5t31ndth35N6QmXJnnOuS9mx40D
R0VIZWEWOx1GaFV/mHMyCXyhs0wzMAQmvlvjvHYROjttb7UaCKNrpj7EoEkRTHli
7gKncqok5KaVVs+RRyeVUkXXjBp4uqCElOeXIPIRaHQocSGoljTN08zvZakO5CKG
TY37wnGVjHU8t2fTaHyQqaRBoBf4aZtVh0fdhvHZ7e81yO7rG5y2UbqiasfwM7ij
zT5GeP8leBjkt5LowksAGbTc4HC9msrzp8nJ7lBOfvCO+f7li+FTeD3eC1hsoOPh
HRKynpoHI59RDo+JWvRkGQyDg9v9vaqVj3pvUTPXsW6hf2EBjLL0EoVI8lAk5kDD
H59wzWvZ/X/lC54qMb81AGeFUyMVJ0VIZtI+abShDG7BX13/cc5iZpJowO96vmcl
tAtykS3PfGs9ZbAu+2TQOpSxltPOV5urDDx6HcgK4oc5yo4pgJjFmLq9inMYTyWh
vVOzt6a5nORrFDHr1jjQUGpAqZXeJlYeDxfDJjKKjd63kialcjkIP0psUDKtY8Xg
AASwmr1zfE6MF5XGwmxkD2ASoEF6KQKyUWmWHKBvOsV2HJzEqlTFE+c9zveT5vxF
GZs8HETMZ4eJ5QnP9GOC8F3aVPCAdk+p0mWnd7oxQXlgl6AFQPNT9UN8+v/nd8UD
q2FGzy5oLC98IoX/jA8LMlzrDm6dIIhOjHjXocDtsz3OAAEsfGNwqaQt5LlsIUFR
bZ5Ybvw5QkUa7JcV31XDZbtOp0gSyB5o9e1yfoSQ89GVIYRnRzOOPJE8PCOZYKRi
g89q2Wu9XxtlmkQL/12arePcBUX6oKI9eaWcOw2XeBt4XqMtXFnnrOCyxOzJDj9o
02kWoA1SlriTmTb2Nn3VidVu2kvwgf3oTCwFcdepzq0eKq4gor/QIck03narPsg0
HOEUNIzm+exY2gOJf2aoy7tIA5pay7k5l7U5mcbHd7HyCa1x9kk2Pzu7LO0ztThm
JM6bcdD6ONU0++2okFgaGh5WmnzO+ti9FtY3o+4EqwhLxLf/uK0wtbbir0NP3C5A
6x/gABuki7tkVzZp0TqcNmAvecbY97Luzo/eBCCyy/tN0hcFyOxOXXZ4iWrXTgEG
rmgk56lMXnhrF1T5QtP7WJysHHMo+t1JWqddOFrnuDxShNgke6F5J43SkRl3YdZ6
WWKGiQa4eWc3uWBHhqy9LI1J16dlkJ4j8BgpW9ixbNPqjPVq1HAMRNqbRW5Gb9Ml
g15TcBnxGmyWHzild56UCpQR2xaN7CZfzduwmpk8pRawXD6EfGiH5dhW4oReGMx+
Qtf790wHfOJg+BClKljWEWgoh1efFpCcmmNGcbTU7iub30P5WQIaFPimTHJvgfXq
kSGeRgcoufbs963rMzD7WjjSuBlKvm8P9+ubj7tRpr8612q02vOwbKUFmB2TVXNG
FY+jHdzCHQr2MdppztxVJnpiqd18zUUMhlNwTU5X/NEPrkvsGLP5hJSYekoaw1sE
wXvO0sbxpUhhCX4iqb+53yj10Uu/BYaJtFf7HCY4TXvH6x1xIjWvINF/SjcV9txc
PWsV/Ryk9DUa8hOshDMUbC4tHEOwwWyIECRxhSiN6tw+03vk+kaQmvkBDmOVQwWi
3urt9+Psh+wYowFJ3VjjymaOW2zDeaTUH9wcv2lGoSQPwmKYtJmTJ8p/0eq6F2jR
7P9SsGT3x0VRK0g3VuVX165WJIDD7gzhfxQvV2/k+8huUfClor+F1H1u0JRWoRLz
fec16yLTGenETTKcTuh9CUvKLwZzAI2jJlyLR726tUap3+RScbCT1ISnTM9oJTgy
9HEHNOXziHCXICAfABEoVwBTv4HW4YeV6nbKOjAo+5I/SpSxy7/BKiMbKOEyPe9p
r5aa2wZUGIxt0Qr/Rt5V2LDCqgJS018QbEKvaXbYo8fbrS9qTg5fjwV5Oi8gni7s
bxaZJcxfpTLrCv+AfjamhAWvlXxhJZte3PUXG6xWSHfOOpX+60EKm258rrd7e4VL
J11EcjNqmYuTmt+lkeaQUujtuSHHGD1qeho6dS38+R3Wkpo//8a0hQpVM3GhX89l
vHTWtPWmpgmZygEKn1M6jlRkXwCUBA9Af4L9mezYRvtFYUyYAW3vw4pQFoTsrGy6
t0J6agiwKAHjhzfmnTKrW/cghy95EhAxKRnHgkziitAks4ETz/utUpLMhDwTTVai
B8KmqOO3wiWKNTFydERjXJ1xPNSekgdBnM2RdjCbulOLTOHAd7s8Q+OTUy7SSVZd
x1j5LG2hd/OpzJJF8d5VeF4c3f8OJ3y9sepmsF7RDrbTwv6ZoNsEe7OTHLZqq6We
5VuX652DGNZHNjYvXTvGOt0hOi5rZo39Y4ehHWugOk5VRWrl5K2Q/4ZfLU5aocWZ
XWS2T4LBUoS6You7Zd0XMlQy/q/jesQ1fDNeiTH9Vr1144EBtl5XQmnwIwpEkOzN
C7TGyBoY95goRbqY9/PK0PgzP9kSBjY7wPgp3QC8uz4zoFshvdo93+s4PZLdOgS+
GHEKl1UShYclvEEXrQE6OlVWAgzKToyFz7MygnQl8JV8YdJUC998kpIFa5CFN0k8
qRPV+Q3qRnxvS8+PiCwZByxa9grTBnf//6KViu8nZU4jbw0AO4cAYcNmgKFiScQZ
gGxJ5A+iyfLjHBFPQRtSxGLrlfOwfGEbz8cwS6CGtlpzZUrnO+2BDVYnBkUnvYtQ
KNKQHV82O7HYWLUfbZ1kreP/sfeKJ64GuilWPvTTEvoZ4c1bcwJZztCMYGj0yEco
ERG6vCapNHtiluctbtIxw/AUAlLXAON2mAm/FjE06nMansL6M3ZEezhFdzpMdIsJ
kv0IhPXcAne+xwUS5zsyj8RrQxqPLn8WtJmpYE2UPpaVg3WSlZVK67BRPYGecyBZ
5qMMxGeyOCBzbPzc+CPd2aJqh8JGndqvq9OP3+xDdM1plR7i8WT+G93F2UQguZMm
8a6vqbto1hhR8jsKwWPtovUVHIT6fCGhD9qDthDEsNyVlsvk51QGYzGE4icB7wnM
Rp2QzB4uDbYmoQ9ZWDxoOBDijECqZS5hlxmgRyZabtVYIInJjr58a0WQZHGlL//E
tCJojZojGZDlN3S+WkLlbMZwf0SDYOMO4PFkX2TU+L38boYF8EVD8az5xMJ5B3nb
AYZRMEEnxX4S5pplQxKvzTEJGIf5hxE2q0oBxSsXe0kkXuJ4p+qG4hfHMvxyYt1f
6OpQ7ZkuEQ3qcuIuwRfde5zrQ6omci+DpoZr/1lY8wWSw+QJmmTcA/ZFwnCIr5bC
awqxR6g342IaKyLGGdIiy0xU/i3Qy19Tw1UzxHxfOux5gYzfXZmomi49DuYCTEBV
c2f4sNTlVPkf5mTSKeQ6t/EbQ6AvC7Lwek7EpJ7amJzFgcCxMER6vSHXTIDdxofK
iUfnx4zO2juU602LAUopA/zUkkv1zHR8S2uR3/oIS2mHHwzTkfjCuAVpDH4GvRQg
mlgHZGF/7WF0XUajjxYwAKswh9A0REmrKNQ8XfGqbEEK8kB6wUh/RK8RKs7rTRcW
RIpIHsBLF7mVyUpkCMD1zBoDfRfdhB0uxVjTOw8DMAsMwlElUFo2MpQ2j3UFIiRe
llKCSs0LSfwnYdtDIZLlb5lUzT6t82cgONvA85EWYtXVGoXQR3eHe4O0c6c97mao
kjVUcIdVch1EetswhvPKVs6udO9EROt/FbylAicM1UB4pRZDRm9jXXTVnf0iBRso
OtoYAqXjDi0xY/5n1/xyNsXk5HuDArFfF4n3Uy+vQ0UUQikD7+5ZDniikMOJtrLr
kB5TUZwthEesarszSq0D4DHK8ZJJl0T5k6pu4G2QY1ZMVFxbJFZQklCdehwKRoEd
yh9A2Kc6ioeKQxW30lMm9mPeRjeC2NBOoCJt1gcuHDF0MuFSFOxXGVK2c2yeFarV
bTLsaOt4kom0EvIkxbI2SLGr8relnykij3NexpwibmPbzmytNP3Tsu1fM39fGq36
fI7Ah/G8J+MKdSD/0iGYnMQf173IUQWlNllC9QdDAoOs9tJz0hsIoai8btL+3G8w
t2+ZRwT9NiSOvGxlFj/eXYEpMxcsWUUcjYhw4DjpkjefaPME3ybygokChAuW7syf
vqHSMFmamVSInomaezLJrJ8ODv15Lpg1ZkHbMV3gpE7qn3yyhNsV0E2h8g78h/rz
sNrM/1p8hxfYcQ3M13TdJXvlrPhrQHqMDzY1p1+9DQp/vqq0jBJNVd87VuqKpG3E
cPC9I+5SGdUXtEA4g66lcKQhK9zgPYEPz0oe5yJZYFf1g82GbSjFonPD3HICg/3v
V/Wxc+oGbSTV+V4YGXjl87OTYHrzyMl+UhUNGnxSukeGwlqbOE468gdsFT8scwUu
4imToUhi/t+3TtHpx1/eyxNnGZvquGTghnRL809jDBrEJVXgOeUOgTQHusWI+YrM
KuEcXfygyjFI/tlWXIfJTcWTf1akpqFkgu+BZZgHFB3xQk/InI4DRZrgqX0kQEGG
oKZwXY9V1K17uXv84LcE1ZXsYMwaSrWRwS0LFC7aFhgi7tKpyIm0YDETUa7LsazY
/DM1ZtnaYlfr3fIuMdv3uozx9kYKyu/CDZwh7qsMgcrjHtowMtV0+cIDchEMElql
GWvVmisLVb6CGr6JLeI5HGY46GV3JsxDIrePwka8IhqOB4uEMVcI2BJMr5EFF7D7
alLcw+/M5qUtCz/JGLgb8Lm1X0VrFCRIpbCoSIu2nh6uY3AceM631ZJLQvGyl2zL
d36SjZsRyJ+O8Ix9NVJh/1sTJLzBtP4a1SkW1oH9zis/lnzl43jMZQgKoXxr2rVp
E/U/w+SMULUKILDCgvw50Oj3YBJvfl43pYQPRYz/V3eg3silVU7IiCYcO9hyeZoS
WgIBMwJ02yLnxI4YBLA2jZIYklDbPmBVA7uaFD14R2wj7cEaRawIsPKEwcQaPBcp
eXF/qiJbUzkarPoSV/5FQbbwDbbdH0dKpKYTDdwc/XPbSNaIihPNX7kBa+4IlumK
ke873I8HImmx4i7c6slx4Tyl/YA6Pzp3B6nF/DBNOkzARBmdgiDFdwJRpmguQDp3
6zf/lFK4+q5/vKmV2DHFtBn3th6d0SfQG2/sahMccQCgu0KKMM0F0O42vFaUlXaZ
Vr24Tu4MFUjC2ZEaW7NIEE+LMOn1tibkKiKfvzUJZ5JZMChOcZe/W6/eu7SKmmr6
OjxqiBTVwL+wO9pKK9rwlZqk5PvzdAoWX9C5Emre3Nu+xXW95+DwizpWgQawlmYK
uSSCDV+702zV6ZDl1lyqEtCihtGKdsPy0ZKxwyZiU1zdVdPQcV2vWZd6X53b5vI9
gt0Yz9zSoS+fSGvIaZsWtwsYFMZ8ki29Y6gCeFZbCLqcpNscosLBWimfDlMaK+vC
eG9nBQqHRuZmjIrtfG08VDpjgKu1jy2T6zL3hUlM/Xy74Vj5bXIeYs4XrPJ4Vyue
oUv1BjlaQqjYN9DuV94CCkHUjLwqAjllcckogntk0QxvCFSxJGIn+3QCvVtomRp8
3dixs+y1J+zUp3tDFtWTAC4orDt0KjlWaWE2JO/6pwScRp3mnip410Los+0tOBpB
oF8pdaiHjSvyaV+7P4pBL/R7eHXRTFej2YgnaeS4icuux2wPNKaG4KN05E+nNYw+
gShX16v4CMheYI/trTmO3srPQr0e+lg5Atm+7zIGFMp69b95mv+hHIGqUXMHKynU
8pPLeLCyqefTPYqlGG1K3MK/R5epaCPjqm5jTEKphRCSNAVhmy4mJlWrfZ2GU8Cq
dDrGyek/3QDqBbYcdB/YkQekpj9pGJ42qrm7I/Kc/MZKFBgatxtOvdAYWSGh82DR
3CUZmY2dzXDKXDZPy9p6GOPjPJq0SFjugTmHL0qwMmmk+X4C23YvsZsDZEHJ9q5i
0q1I7+GsDrb0xu13g4DY5b5m5D8nRNAwuz6zIYR+C6vYSDrVqzp+a4zpvu41GLIM
c/gp+/wylNq2OykN6F7XgasdUGkz6uzyVyVP0fw8dAr0FIFVesvMmW+QoQUNVGI/
auWydu6TghgQLs8wGg5J6jGSFIfNwvnPhxnED6rAdZhf8TvdkXLT7IOIFFd2at+k
lDCSvsuqeqI8mrqUPzAu5UTPVG84It0gfnmlRtYd/Vtu2QSdCCnc0lhfiud3THo6
V/wlRXVcN3kSalTu4CcgFWD6A6k8wsrBAringY2T44ltjp6SEny8JsP+SvjxQgOu
g1bAfXxi2xXsE2wm/GZgb6r2dXxolejCJ16869pVpwKlaHlL9VAIR6gpsTd6dIvM
m8JW4JaFeEVV/Hi9uewi0QdqpAXSYfzivm0kPkyfTR8/8ALG8Bwdhhepvss7MIRO
Wo4zL9qqo290vfth2daP2WW+6+C58x3AYZCOK/6BSu9wHQfVO9bOmgdmx0cMVtbf
QdNaKUceZgGJ4tq3uHeArfeeOR2tWrvW4USa9yDGDGPQONblaRdaYAlciZwpPTPY
Xdz8NYGiiK36GqcXAsc2GpylrlnT94FmUPXFfeKtzVg+vS7tWAGLHky397O3VYvj
b4J3nBxcViRDtr/vgsQf7RKnzPHS+WiNGc1XTh7b48vRll2yuJ++KmWNcEIcncaA
7+kIzq/RbtLR6RlMRwTzp9tCArcudTTFAfrkiJYGWuTj4eU2ZBOqXxc/hO2gqBnO
aT0wYeFnFwmhBuTL9+EZ+YVyWq5K8EPV2V2rpEAlpXCNgc2zpHsiFPEEmvXOeqO8
hJyENy9lqb3PtZ5OHZa9zloRbEKNFCl7FEHuP0pczd8QfUJnxsq0xJyTwmq1QInq
4aq4ofJ/yw0q4AQsC9ov1mlJ+4ujO0LG5EAU2NNxeKV+QSio4qHn4wFkLuAj7KNq
2Qt9ahBx3pTDfzNjkIUG8DH2VewGMmCCYL10KQBa8gjaS+irv4wkPtZYptuyGz7Z
0STSksEgJWyE9HXPts0yxzwR+oDcj1TkJyc9vVJM8LZYvHomvVCfS+BKqnZcVhCP
XPEaCJB+o/LpJS0xwMpncAdqqSSpK1B8ZVfUv2FjrzRTh4hi/9l7w9aeuX6lm59a
cldJJitRL1zkA/WAjGKUQ/FU7uCnFW8Fb4xZUZGlPHAFS/UrTik0cuW+uSQ1gj7H
CgXcURfsD3kmPimnMv2hFvAy3qse3zUAs2FcRXNMypba4sQLWQ2GD1Cp2VOAqfgF
ryJPdOBPubcd8BIwJ/dlufjuG2/sv0N0M4iQUTxHjK/Wnnpx2jNZZM+7j4zmVXcI
EXckJnQjOLt7xChTVRcrO/2iANQXYQCCOiSDOi41Oh75IqdxiP67aPW43IhZrCv0
P+2e64xF8Blz4EwVlGLSXkT3dj/W3QFN31eJPECKP78zOsPY05jIVtV97ILm/AXR
GfV0DBD7ODeXTBNvHek0ltqvkPDS61eSOovkWEGgaH1JAf+SkOzjACMEp8YDkiyq
hQ0A534EAzOMtT18dSIuIL28rWV8A9qD5TCB04TY4try6yYXsnwF+c5AXJ/aaWpQ
5Jf08JWR5FYJZV/cmQZ4WL97w0qv2kh7J9AtO2NklN2DH5LOoW1MPk/IDVhPM8B+
SXJxHLvITx/R2hj1aAlhPKLb4PvuSyC3V+1W9KMx8HBsgU33AqVqKAlZLqRozXtB
A/kqZ3uVhpqR3VVVegM7jLOFMS3KWdVA4BC36wVwgGTDZN6hSGPZllNekAxBC5DY
DZuyq3iUlJeVgq7Z9HYOWnrGxfg2hEoBm7dnvE1Ec1AJZw9QprwCWr1YVUN/fHVl
wI+ukma/grMNZ0LX+nVDZotbBa8r9m7MqmLz9YRJmRs/oxnwBHDWSauqEit0Lzo6
x4RDlQyJmJEwmSHEi3VWhXz7tFu1Kb+h6cuCrd3MDHuSuTOMnmkAVX9/Sfhm6fsh
nCsWeQdRcf+c9QVGMipojyA8GAmItUNruz1YeIg0oZcuMJ1+TIqVMhftj3PdkcUa
/jvnJl2iL3JrcQwfUJD1922r9/X0OVdiwxiOcoW18Jdkc4nMCXf+umuoj+e1r8Gk
mF0r/Reo/lqdL47vLEKFsSzHVqyL5JBdmldl04i6T1ahsk2NvKEuIV2pJE5eukSf
uLbbyqhVG9JsJckW2SvyUGUjh/dRysLZe6AzkiDFTop/J2sOeTrzB6EN4BL+SuDp
t5H8zbWPrhFDmZaXCWwZaXwE6zhF8vmVtdNRB8Lfvbfc43g8ffD7X2Xn2ZJ7lkqJ
TK8/mIhjNgz/ZhqsEVBeTjiJXcfhwAKWHb6Iys3wA3K4EjiI28Vj5KWOQRRn/ZIb
QN9c07+B94uiLjBi/IWTr/SWBv39nLqXAlZtINOoqfP1GiImSzR1LAdHHSE0xJGb
jwHJb33o66PDYvQT223a93exq3zwaI5IozpVJzLqMQcAra2RQp8o5cGTRKg1pDbm
MmxiYywt57Qrs8oDOCoojwhF0YJXNgVUuUH06ntexeMbxdGHx6vFNiR/1dV/0o15
EWcWwp/kUM7LSwpWupTVvvevTdmZoiW9cGJDSK0MfrtZ+To+xueoD981VB1xnV0F
B585iHi6CjA0Lm6JlKe5yPAENF8A3YMhlVi1ApWlg4BkU43TlTva52RGYLhiGdI4
Hs8+nBpSd04NkXg59zyTKe7iOi7Klx14hqPGa5oYuECO37lE1l0Nhov/+u8rGdQn
2EiGq8OEQwgnWg4r9kgWeRovF3uoYbpwcj0EgcWJz/P0Xk85DQHb6UoH0eGxPTtb
hwSqFTOvbe3VV15/Dp7xK2Ma0TAvdo3pOdc5cbMG0gsMZ2a+wIBldlZ/JHJx0zHo
iZCTPRzmoCEu4d3dlsBLkaSDzBQo3G7D7Y/Rv5GTYocfsJlGsDVXwuOqMLU4thCS
M+ynqY+EPMdJISQHy9JKvXMjD6o5SsZEHtdp7AUBl8FwE5GdYt5roIxXhL+0vC4n
3A/Dsu9tN5CSvW8Y+j5GhXebRL0E6LqLCaC/1Pvo80nN3fo5/wnXe0t9Qd0G8SUW
TlZ6nxeDBTH2ey2sXpoCIbQivH1Ep7tOFxB8dm5iqafRBmCxsUvrv2GPFpFjMKoc
pfM951XWoPfDnXNSyZqXfgVgqXwyjfb4ROUVA5p8J7B3OS1CvbTdV/YIci5dbKE4
4OOBAdYKjUnrBVJDGKUO7LTQwLvYOoLxIoxMu50lPUcA6za1OoUcU5vJBLVczzSl
fZU6MQUT/E2ElWrvWuldHMZTbiIbLRYJ5fllu6diz1KafCADqUPpiv5tlKUcHK+O
lqs6PiabWbA1QnjHEzrksndDqfotv/sbx3mN2yiie8CZqEzwymAR6iCG+SKbhfm7
/maKTxHPnRPXbDXiYAdEjICNdV0pt7XAHC/GaAKd0iVsAm51UK/nuyv2VzFQUFkc
ycy4+0JrwodT0BAMOO94dSUABIlSji7YvL/1O7pXWXuMwAXL9FIBXL2OfDn6GZd0
XKk92Z63dWPoaX7oggXk539HCYqAcylb1d1TVNB3RMTPDo5R1rk/9HUOSVf3rp5r
bWrrm3XOmQzhttUaPue/lmDBDGh3M0mpqbxISbuEsKqEjyRvTSfHBJDUtB0A3Zgh
hB61eEpZ+1Ynbcyy2RSY3Dsnio1Y9lHVzk9MDqeJCqy0X/a9MJsDO7JT/+ocJ56g
H8jeVCb7jzluvYznqNZWuQLwRx1SrpevlorNkfQdZuic/Pd8EOlkvoINl7BLvTLL
EiidnHYcEtRyk3ZcDMTv9yoXNKVhoLFyvSBdoIJ9E8uoNRNU63Nb05cYA4YdkKeB
moN68xiLQ0lDl0wEUbe2lsoOUesXWXx4NOHZ78GvofV7UKPyzDiXScZoFD36wC5g
+7SCyCJVswDnw7Ri+Zv5inlh1PE5hGjUHMt45zfrVZCl944X1FPXv6LhBeyKXXxY
Zc7qVZHaA+zIvw4jbswRSuY/Bx5BmYLoXuZBPjYDYNhGfhkQAyb+zLZvkIm6MakI
zxzJ5NjPqUzMkF9Mwawgdo4JsEKpbIGNd3DB2803LKgeaZBFslzca8hMDMnLrxFw
M33uhIFYdQmleEmjHzq3UuqzShiM0lnrCP1ka1Ym04ZsElAZl6W0A+3yqXSIyI/z
wneD/Am3C3lH6Y0Zyf57XFLc7XoJ+4wjECRNjJ7x1LpSfRO5DiGXxX8p7SmE5MP4
5dbQHYaC+LnOTXbEXGrB3Y8IhIACVYP6zH+kMTMeuLMneiSDoqBYJeWDtkthRKnH
cKOImOJgkqPsCzPBKxewU56hoGDBbcrHpcxHd+SocqYM5tx993oo22r+vgNm/7J/
03/bFwX1Pd/2Ie5iALzJsVN601dGOJHZrKNy1CGuUMVvMdAz3JP7VuanUGsgn+d8
akUFn9eFHZJ+HvQm6/YKK0TzB4DVc5V0WJlmZYgSGcxzkauPD0T1CSEjNMGBmR+U
CeheqFGPQKYC+n+/W4NmYbH/pOzuwAfPRFzeLlH+OZNqHzfOPQQhk+t+LfxMv+sQ
cPlzugw0o3eX1gCcxsH1m6dPVghXn9+uRykUT46UlaUgIqJsIpAjokN0DmqmXE7T
rEb+3CW8wiS3b/DqL1ZPcvE7XpV7H+YBXSXAyJr7irREbe0KZUsB2XU8M0lX6m7a
Ljwjf5hy35RTT3UEDWcrYRDrIHVL2DJdKSjEL7Lx0jQZeINA2Z+KWleTltVZMN5B
dZLfpbrC+LLkJoDBcYlmZBKCd+SSS/lqXUa/beg65mrLPeloTyWSlf6RVDSdiFWl
wxbYBJOryqo8Ou8ERCo2umlTZ1K2UMb8QOVLRhJMCI7jlGXMWT+nWIEsMVlxMpkH
NA9POKGfxYi01K1k5Eo7vuQA/etz3DxLEqoActCFLthhoepy6tM8lJ/qW+nySOeV
TIFxJOvtoVU2xR3KHtgs0MlsBlwxmlWrPdQgxMcx48WWSsNATYwrZNO9BhnRpW0+
CbGFySzhpmdVt0qN8y1zkHdgPry0fsbx4hloyLxtWXIXzDK8HMyCZiaAP3h+zaUx
VrwV1r9cy7lSZ+Vn/cjlEKZoj1cz5Oa2JZBlDS9LQpFEcgosFOGA+/ZtP6bUQTzj
8n7Jg7BzNouiumQCT8aYhkcWp5/ptwa6Smt2pYLk/GZ7RU2eH6BfEWsHuA8gM6tk
GwwDGL4gQWbwwQjZFesyCoh1BfDTfwQ7undAo859yxAkVeIC+r44LVJEpwjLD/mc
e/DxKc7jpBreghaBmvG/xdsZffMqDjHvYeK+z0o2604HpI4rbR4VTX0yzXahw5xr
VStXnVsAniQZXrZeulVgHXvHeJ7kAiqoAFHIf3hcJwuXjoQKRbxiIaN86f9b6koR
+OEmnojfUyScRK77pI8OuKbxO+LPM83rbkDTs1L+t+LZ6KCx/R12jjU1K/HTwkyB
E2oAa1ZEaV1DMzkWWRyl3MPIsU3wgrYL+QdcCcd8lYHxa0bDYSo1Pztu/4ECBvnI
K/2lL1pSI5ooXcY31KaO4J3GB/hXQ00Ex+yNnd3sWVvG7nh4lk/FbI9iAWTIymg4
DiNUgrnQTvJunyWK2N/RDs+MlamudkFWafpqDYVwIyOFI5MwZs34xhT7Y8NEorUv
0tYSTPOXPE3oy3a8d9nwCPbubU0+1J7QM2oVu1lihlnLChWnrTbJbac8HLlBG4/P
7fJ2QSJnUXKWhCuHshUa8U4A4lc7Q+mvVoXXTOyuNDLVbWqaT8P7OuKv51/aFHx8
f1iOBviBOVgIlSReEj87TJQACXFmVTXX6N86UEmsd5iOlRa7FGfE2fPSS9Pk19f7
K/jTv0hPRCDySYnke6qYG+InGK2sOVnt2da0gSKhF1ALcipDQyOwf0q/JJlJAVmv
dC0l9vzbzwh38OiUQPuqxgzLoHVyOgrm1GITTo9o52nWScSPMJ2XYKrdi9Pf8Vlv
5azkAzi9NyGoss6Pm1YsbgrYnkJF603IuBle7uo0RomAnEx/zOjkd3vP7+B55d+6
chPz7Y3BombX9NFMYu+50s4/ZnmG8vIhkCBA2dx9tA3Yzv1Ic1ATNSq4Klt4dcww
sN/iqvxeZWtSibAoyEgL7qsAmzzAiacMJznIjz76aHYyZxITaub0T2jbiNr9MJw8
WaXmFv7KJ1qtdYOyCiZZBfZ/aD5AOLlbbYmyzoRI3KbM/SU3vLMmqk48UoDRcf0G
OZXg42erHcRbC4FAvRRlhdYxzA8gS9rMPWFOR/rMj85GJ3Op4iSU+pbT23QKmAWY
RBOmZvJYKgLbjBFCtHQu/sCsn5+xg5ULoijKEzx8HtZUXEv6jZMb+UHWF9/xGZ4G
TJIeSVjKjvcZgNeMDFA0Bq518jxdaPlO9dGMLG8i7kgr/sG6uAe+WybNK2J81byC
weht8zOh+EMLoEz/ee8oXX3jV3X5vcdyarcrpHY1XtlhHl//BQEUohpzfXvoMeO0
gQl35UYLK5DXhVMaICKs6JIdMyRmmVEaBeGjdqck5cWyEKl5e2qy/uLyHZ/zVLxa
FQ8Rqq4vt3xVorEIRBZKZDJPrRSjF9BvrCLuaY0ij+Qtqs9RB7UmmarxqbIkJ2PZ
dcyo5eL0Jl5FfMt65j4+8omL0In8CMg1SOAWXMPl9SivadqSqiyZ6xqk5t3NQ0Lx
lLuwcWXWjtWA4wXyQcgE/a7GCKhLwcuLBaC5lmPG87aQjI6W2kJ1vSmvxbMNF95n
sYVpklnJdyZdXGEyewFwYbzmy/CR1ZsZHwFAU3JAYqIbwvnKrdh1XnyHqZUECng2
O4l8ukL32rbF12AQ8qkf6HZxtRdx27bzefTPf9ygUUrbxIr+s6+zCpjPfruZ1kTs
D1++amFFryb4ng0+MnELK19OBfLV0jeL3ETAZxgtx/12fYykUi+eH7cFySkhft5w
j0bOAs5Hn/UNqT2AHPdAybFLbY86w7Iroqqcriq7XOvYyacWR1zgJnTPXaFW2BYs
iG3pXkrXadFRMnmmGX86ND6holai6urCrCNk7zBftlRGjN3LxRFf7cKFde/kjwVJ
xr9JoIxxfdI8R7TdE7PW7DxdRdPONTwZVvENac7j4gY5aQhsz1Hw+1DBjNDfEjHU
LotZBsBuLzH4/iFh+G4j8qoD3m/nNDDpBRDPNU60ephQTYIjbK0s5/tvjJwakMx/
eRwNrdlo/0r95TU2MOyxZfRktOCoMk042Cpz/s66CZMSiMNpns8pptf64+3qbeg2
J+1bSQOXSYe30L7DSXJsuS4nKr31yUDXSgpwcoEaxbtfpJMtHRLOU4WXj9A9Hqtx
BeTTnJuDCvBViHLjX86KAuv6aFYbckqfYx0b1hrqvHCiwd0rmim1CU8AnXun1uFy
XtSnKrhbndxq2I+gyxg3iPqfXUmOWqYBxnYbf17fFn0g2R+i8kDaSMMqE7xwzsdd
Ky9g7xG6TIRwVFaPsfVBP6bA8NOcGQ3UXwBWjru3GGbvQwBKXdbj2tgBfhZfKvbV
sshLsqaPbSBLq5wCdI+eJM9/gXQ0iCuVH67kKyiLEUji89IuOrjwoTkSaRgmSGde
7Wh1/7AtHyF60OmW2HF2osboN2rD2yvC+7ApYUDjJViPHgQfUgrsnlEWPP5kKKU6
FIqqm/ENgzVoyo9Qqnk0jrzQj1Fm9L4PIXzRSMd4gyxOtoJIaNMGhvxMfBtV/hag
VBAgh1myEzB7VF2J8ZrS3gOtVMh+5z1qANguqnY3VOWJ20pqj6w60YwHKoH/HOFN
+1/fCca1e3C4F288iyPtt64/2w58aRf0RWvR3dMP2Q35GQWtoQvAxhN+7ZPDqgsR
yaH28u6acvsSRYKiW2LhOj9RWUu6PtlNyIQoy73AQtuHb/r2qyHZzpv9Cnn5tW0D
EV9mt/8XmQd4OK2aImSV8W1knE8ZNMngGMmQBFMy52+keGFSUaLn5aYALEmPCm3k
DRtgOi75LAhl/Lir5zupL5UAkcgYssREPZFEQFP4XAfYawuQBqJISu04gkg1sxaj
0w1jR5xFGXU/cULlitZWEJNopHWa1saHpniFOYyKEGO8zFLsRnTjv8EkrTKz6Icw
Gv5khzGl1mU/hv6wNvyzVdDVl+C9oI1yriD73QgMPw+9AHYNgYEtAZ8wRTewyBmJ
GNMARXiS6uYH2CqVwa4obNJK+NA3Meh9u0jWMrJ+WyhAJFOxahAOl1XpyxAn6d+G
3WjUbDnJfsuLO1TyzhsmgwcCc15JYQQjpLKerPw199ej6BxAXcJHvkY8/rPpLs/a
gGCPU5jgMaj9tJKCojcUcbFTs/1Vu7PRh4Dmd8vp0etVsKZrjcF26plBCp0prF0z
sxA6JHsfuEFYIlImrvcQFrhEogisBYAJ2C/ul//ZuLPHC2ABf7ZrGe2jHp7SBfYr
3Qqfm1IGcrkG3/Dnr0SI891AZEZgQbzOyqvAQPvPUa7ZB/AnFXtRrz8j+VKzNK03
pHjVnKjdZ/VULAFjK09O3VAAe6ZbbSOyKxNFoulYSLRxCYMuUNNBEJqvMQ05Qd7K
dR+Dit0JjxfQadmpkB+lnRqvtoKrWt3b1wjEiyOnursSCCRGy2k4tF8MYXbOga7O
zOceqGcrKtDia08CrAIWjIPLJyUmEeE3BLqx46Vce/XzVU/617cvmSj/1BNanfOX
bupbcjfvdF2jMAqID92jaGeeQeKjHKW9qsd4y+FesjH5Kbug/PdCDZQ5ChIcqH7h
KeXIahVpzBCG2Jg8oprxpA5mcf8CpmFGxUD+S1ryA9N/MFM4T7bcxFpWUOab6kda
bd8CNr2GmtKXIbc4XP6TVjvRuMqQ3TEsApbT0QS67VqjOtb69sGshQhH28Vr5l/T
4thGLMy23l/QTWQ9usPXY9OK/0J+GRaRJKR0cnlJSyk6jVHloLKeQsTiWiG3W7+U
4TJkPHDBNNod+rXWHnM4ilQH/aJtYNE4CY/12typ+KeXjkF8ZpLjpUGy92cOQIG8
SJMdOO8+dQ7kS+68IjgByXq7N2vW6xYQTvt0fOO0KsflemsCSL35Xf3CjszfQ8o6
WI1SNLRoNQQk1bTaHpR4pynzGmEjbMYMnm+jjJ94ttvAM4mw8VNfoQeZz3Ho8Z+h
XsrlCxv9kxu6NtSvqepKQfwyVAdJFtXZ5RdifW6AIrmu3ktT7DlzGZc2gdQTNh3E
2N63Fjpzf5uEXtc/gU/I2+45rjaWB4PoZBui8myoZ7oEpRVqAYWw1d9IR2OMpfi2
6S5QdLfNk//oo7PwprMbLOGaEBJaQ1yOT/cA/pnQ4cOVFh9xjiy5n2iC8axMaJN9
CZdXNfylgTbQoOek8AKeV5dgue36JTef6/1wNkq8xUeT+YkGr0BRG4aT2BzpSr/D
LPhd+4chiEoMgzo3IeBJOzE1P/LWl/zKP0Zz8+j49StMY3WH7XuyORDXl6oHnhDu
nzGiQ0gV2A8fDSU98UxNzjuKMZmwVgdfHbisgYvrg11d1Tyghf29IfE11EopBFvY
n7nL5sYl0uaFstM+ncn3NkkearJ6X1a54sbPK7wryds0qZWYbHs1w45L/3Nyac3H
VzO4ayPVt5PZY0InIeTeyKF50s87XEW2KL6/QQ0N/7QgVkf4GLlqluc0v87AZHTF
53SqFgJ66btyX0wpvJJTQwrr/tMwmzjBKrvPaHZUWGEyT+DssPy6KWj4v2jdBDbl
zhMREDEZmg+oerr7KxtnVDKJUKg8JZ4ttQaT1bq5JdpC0hTk6xLR+c/fvnqgmaEL
G2iZoT/1Ls/re+LuJMpxzPdmf8UQPbIdx8lmSm5/IES5EqirIFPJXwCinVaMudoi
Ni/vyPXI92eOmyafsyaBTLOFnztuEX25tUUKSHFxt3KZDgJ4TfjMpRNvjkt1v6ip
K8p8snpyuKNZa+NjcD4WbtIRemCAnNbcYlOOruvMGT0HOep4vyWw9/yTKhXVMx/p
K1bA5w8xx+w5hwI2rpXov6axdJHlyCNUnHNDHSfIN0a5d7bsxtfNZwFOJUJBCswH
YMfYOiiMN0pycPeea5wCYEOiNHRoX6RiBYALdpG2hZlw+vLG5Ij4keVtOVlWVPFt
anTzjNPqradb/qATajl1Y+Rf4CYhCaCTajqqmIM5Xj/MsnoFqdfH6DnY9Tin4wg/
d/Kdes4HiKcUhZaLDjtndJoXoics8I/XEf644A54G6MsDqrnKCBueuF50PE51DUS
gu3dQmUk/nth1vSMn7v9T5/crmrauokIWicoh8tZW8mCC2PIaXcntdtbI9ZfT2dZ
c7pETX/62pGmNJAs2lqkdsSvCBiVt4xXwWWwwsW6ZiwSCJ6V8NYfQUyNOqJgaNnl
fEPU48GG8ohONm5goitztldOL4c1oDR6FUzmCt/Ha0pp736hxfX9owQvyPV9FmO/
kYF30PxTW0fQAjWL6DsvruH5Sw0F6WEVRlJRHp9cxrruhmRR5Z/6Fygfu+hXrQkZ
8A4YXNg9FM84hFpxvKZB2Ah9eQq3Iq9OD5qg+OMpQmIYUveKzwV5tkyLhW1YeR9D
BmMuLDBf6O3iTBUtBZXk4V2hm16rqO71eVMYcgBbf2X+eCgyDpon8qqS/g0CIfMJ
SmM/tOxlWBAJ2qgrFQRonOKrtC3qphaLCySuBx+vaAxk2E+9InL/fSuumokIdsKx
5pZyA4YvJuWiMOa5OYepbn41R3tk1CuSTZWnvK3uKUnxEsBeZrS7NZtaWR2J1wPT
emLyLQjWst9KEH9wm2nyrIZDqVPcbhHtvGFXVr5RrkiLRptgShOX1CaLQgQ9J4mh
KUQpOgFuwliAK+P68mMk9D/j9B0VjFB0WNdQ7MoP3Y9FqaYZheabOdUyKdynxIcp
jKXdQwO/7xPQeJWPUOM1fH/faaEbfFtRX8SYyInmjwg8RA2NlywZFRwe2BgPy905
CHPbKA1g3xoOBvo13VV6CfJo7dU9n72wJ44JZD5NOrqUtIAyiD3Im3blJamFpxoi
d6VwuqawufAPQTo/4ZMOuyTt3TzKMpnIk9J49L0pdzzXgsADAEf2Nqd7ljsrFwcu
rBcvEb6j7uXBgtcXT+oIZrz2ugVY8fcv7cv7lZeqAR6Vr43GGfq+P4sLaGophy0c
PqYL+jVFdniE2Z/uQDeuPD3VyTDgxbQZTYWtSox6qCi19e9dwUiL78DwQCQTKMl+
YIb58bkmAlvfaA0IH9RMB1zhi2NH9zS4UDf/2cJ4mGPj0/Q8n0YGGk5nDXbjPYzz
Dh1fP4bkWs4DlH/EroIvZTZkBPmmCjGHy19FY/rmV6dEmDvGw8wH3e0dVtQKDGqJ
vDtnToM/By2s5I/t6JjTShYu1U5klibOpaes7Jxu03tp5Ib24DgZdRUjpKko61eP
dIEi8MYDStXG8aGkWxOQb0ahkWfYQI9yJzM7kZyWFtgUMv6UMN8e/NiLQa+FNqYN
WxustsICQhc9ZYA4Q23e/dClUAWE6RDs5DvOsGCtd1zrgE9Xselz/prO6+I5RoJW
HKcVALf2cYL5K/Qy7KqnVhLXuG5P7O/N8YE0eRBcLq9drcIZnuLu8DpIiC0qFs2I
SeoQVe+OwyM3Cu6W+TNjexcx/9DI0xIF+Tg2JAwtt1FveGiRhKb78bqjfZcXf2bG
m2pfgTzqPaFqes4u6IwHxnf+UDnzljF1WVQmWcBX3dHgGnCdlKUr0TY227rBfR8M
VxM8BeBmYnDo5MJK0Oi5PTXfkYOvIqEkv3TQlbwRp4r3/rS2Fkcw2wgFox5y24Cy
G5HkclQqSTNHwtcnZzKyFRZbZgsxxEEFiCk4YseDcMNdQCZ7h/+HHp3Y0MFiXLn+
VmCEHvqczjNYcw8COqII5yiak/twiMP9ZjIBSpigtlR82S13hLFZq3pI447jOjNA
E0VTDJz3bZm3hXdNEGbamYbWxWAFCRp5lqjaSg31iFSUI7kGT6ZZ8YOIfqovC3ac
iScGGheD85Gr4KhwnxElYQjmgn8PWZC8YQU1B6laDE2UZRs0OhIZAoaF8vIsSy74
sOnhTb22AdTix+aP/1A6NIQjmPMkKUUyEuDK7Jlpwg8xzPW0Vvj7mHk0GigYOGbD
Kvjz4QftVP7VmjIvxJOgzP81jZwlwwuG4Wr+2g6pCxo+HKVBc5c354Su94PRNZNQ
Jl6O85MS29ZR3RIjSxRK1xKjmu0uk/QpSUsDzAb6XLZu3fcEFai6Yo8GGajWxEO1
1kaKkNWdE0xJXcRi9+ZCdbwdFgaSIY8XZujxpeY9Zu2HPBJ/5YpXfu0eMt7ITJet
FDV4lgMj7gsH7E1Ygv+eSbApNb8htExhkMTv+xsf40KPWccEkh+8kQNA1SxkyfcP
OUo9lJusznKP71YwKhV/8fQq3i8+BXWBha9bwsEdewB4IjApxXaSBY4i19Knc0tv
RHo66MbuqwoOvq0/6uAeLGm0d7qfYb6npzCJyBwtleukWEuuAxmGj7TCZ/T/GwVw
8SDs1Wisi1MOeX2rcEI+FZ4OkaRCuThk1h5V4Yb+VQcOSGNWlUkQog8ADUC2PTwD
0H7zRlWYkCqKtFgu7MZAXcwe4qdF9OshDXFsDxnMirpUHin5xNyIGNTo1sW3IVeX
Zg/Xf+yJIeUj21owngMIvMlKo6W0cbJzz55jUtJkf+h8FAtlN3T4mjOfo7CS3HLv
QyashtLIkrVWrbHa4nqZiM8haIEOdkC3zao7pL8R/l+7EEcmYy8p0yVlUNL94bWJ
WtPCAWTbu6//IM83np4mJ6nkia1JZfK8rXlI7P9T3/mNWWMPP4Z0R2mzu0iPiQUK
5sydRnUx715+E4kCImqQvqNiovEyWgoe0nh47RrjCg4A0LTDwuzH28YrHKGdeNbP
XyyZLas3F25ByHa9LT1KTu7pC914jN8TSlmg2b+/TgaMnhvltJ7ifhSdYMqL0EEk
NEleAMv0mQdK9pU5YHidUY+sbTNaVBSroWlebhtz8U8dF3r99CpfFmuPnzubt0eB
D5J2WyLYFYTLLbMEeb3/xzIUWoHAQit40eACcHe4EO4oLQ6hVs5YLFR5gg03DFEN
BfDahdFl/P6nTPD0ueXeKXER3d1lvxRcvmAAiyuX4T7AmCzgC90rFPHZNvdvd7Ng
Po6QG7zTxBLtege2Hs/YWBy/sHeDG4Z5Ht3RExxPygy1Qv/yfuzf6N5xdJ5d9pO8
n21nA7Z+n2X4FoO1KP1p1lS5MzJmjdAW5I/E2Tpxq1FQZT40ORZCGPmHOSIQvbOK
gwk9x5dSmfn0MUAE6aSLqhaag7KGVsjp/4a6iXTSyJSKQWW68yCbzNisWpG7mwgJ
aeMJZ93MpygzJs9zbQWHxuISFkjZuE7n4cMJ3pIOGVhUVD/mfPXdDCmckaCgF4Fe
IO6V+wSUcwop/zxcSjd+00HzzPNgCuG6oo1QVPlxa1S4Q0ZyUD6GeUkP5tK1XxoA
CAT1LQx7CIi5K4O3Tp9qOHgFqAt3670aePICJaM4vLzsxhyvtnVIa0sl6PjT9nRk
/D1y0egmq5yEx/oV5tGxdQuOhkaE+5dxYtQvHSdpVZCNJtCQQKvcnjQ6tP3u6Edr
63KY49zvg1MSHR4lMC1ccaUYxL4UWkJ5EK3RT1ZZllyR0kUMPazZXLaRLXDwjZCL
h7/txUMe++UfA4kse7dGsMbLtL9TPmt3SX8d8bt4Dc5KNBsJSrYc5b55Sc2qW/NV
6y3PAcOqs2l28dKqtxT/vAnDHuO8pAwsXfWPdux2V5DVhwSmMnV6rHLToYBOYfdi
eCpvNRBlBuBoB/VTV24R9p669vD0GuVuwBg3O3R5DkV5Y5coKjez/4EshjKd927J
4huMtBNxM9scLjt11HNoJIfeA5vgD/Kw3Al0KDbNu10EQvYmMeowOmY7mtSWR9J2
QjL0mqN5oXwhEEW6/GfzJgyCTyxgPHeUb4ZVvnEOehODkim/LNLeynAOOwXhxwya
NDclxBJF0ISDOOokM0uliAi8rmq3nHOQdBtE+z9Epd3yVi4hsNQ+HBqx1psekGwn
ByOPqJKovG/ppjaqg+Dir54ELT8jYnU5RitOQeYtsfYNAp8Vtor3DAOsEqdaq8Hf
uA5qQD24CcY9LmZyIMy0/iXr7U0Mo5gb4FL4a7CcTF+7ROvMudYmXWbJRH/q6yks
HDDZHoUhuubJy5y0B1/JvzPiymlTy+HNJZQ/nFzk6TATcrEIdt0IfxBWafZ5Vyc0
WFiPanL2FtjhTc0BZ/fBEIiqAUgDkqp3+KtoPpC5E33ZnlLdHMvz5LwVFIAQWbk7
+/KmSmyX6PSbI8qJAJtohMX3Wd8xYYY4W175+y2FzjZ89zkKFW9vm1OP9NruZEid
uL71SBfw48U5R8RlCkaa7CgGhxoe0zZlSko4idobXDAT+yhL9nVMR1ZD+CjGvhN+
b+JR4lTeN7RiYscjofi9iG9cJQc3JE+/ttcqPf20mzuxjFUEzK4hkfiys8d6yZep
KBx1qmk7Wpuf91WF4R70bvp5zn35ZAf1XImNM/4yQUqbsp0Ip9A2RlV5inrHuOF/
z9ryLRWROVxFoFyqsha+0WSu59EKa+OU3PmDVkzej0W+lTpXG6TEXuY5cUuhP+m1
ptRXEuDbtpKf1PCActY+19cDn/IGkKiuK7bLIA3UKXrx/bKQNCnNL/79iE9GxTil
ynK34twtLbSSAmpECrtNiavxEPyRdw1Z4NVnNWtVdtpDd8PYe3IWbXB43e72suXm
wtzi03RAo8j8dvgaxivhg3xwKYcvsu97nkEBPe/sur303HkRYlxg8Z1j0Yy2Y9B6
BV//GWXlf5ZjG2g1ipCBhHE+GMGB9gKv1iCwmUbMv4AYWbc0iusVraL/Lr5PxKOj
TqwQDI/DDjESv3k2euQIqmMeZb2je+OKsIPQ2iAy1vBAYruAiEAULDzqn1SV54Wj
QuCD/pootwcVeQPAumc0+HzE4LzTmLz2GJyepe3yJ+5ceEwy25e2+jNwXSPJDHUf
3+pnMmg5Vclp8XPnfxBb3C83NvawP+Ljqkg71SQeld4+040f88XEQ+1yQCLm1L8v
OVfipwZHB85yub+ifopHGzPhI30hm9D0LedlVeQJ6YpGZrWGKgTAi2CLKl0/nxBf
KxebImniWEqtHqDpL7cYytCjvWw0VAu5JlgtkVDNrVwzVe90vSRovoUMW7FABk99
cMY5pknt07pgy16KsEFCGVdB+sU4lpdeAGdvT/3N/ayVChqBYpjD/dAjX2OW2mM1
mR66FtPIEuVIm5iG3id2O2LmcyH0ihO/2ybddS+JZw+7Z4NzdyS/Ch8WpMydKIiy
dGTDbVsoU3fsnE8Qu8S6vSqlqsjfswLIMoZ/DENTnWssGC03UsPCMuwy1Ni/LE4e
oqULVNBxfUMadICHHzHwaab4HvbYeWtOS5VN6j8Hs2aB2h+mJvwSZOooGssIbYnU
0q03L1MJTsnGvP82OJbvqEdPpoKXq5BPwe0ph+TtfB/m6WOstLEmqT8YXcXUhGYc
CCFo6hl++iOL/u/i3BHduLyIWdcEQb/nWHqEca2L92OonkIv7IA0VYlkTLSaXd5H
6RDcXMsnKLVDbQshLcWGErYCHjctH35v3rXFnLygg4scPut0oiPcCFXq4oYCp2io
NFTAjO4Kb3Oc/ps5EsAQgftDMYr2KAfWvKP4qZ3rP3I2vJ1MPYfHAvaTBtRCbIk+
5rn/BOtwhuB0QqRUtQ1h23vkRBOs7Axe5aY0gDU7aOJkHsbjyt+KLoKgz7CGekiS
pGpdZ/KnohJzmsgl3rT45n5k3emHJCtOsYHMs8G6/+2l4HFkZLWuuIeQwSpqPY+6
lXjZp3WTiO32Kbj2H9M3va51bxaEPXj9at7ZSYZE5uJG+sqt0bjGCyWCazehfsgA
RelHXFaSHXKeB3IL1aeZ9eEG1L9gEcvL9GKc36jcki2JDU1iTRrkPMFYVpRt2f4R
TM6AVIT42ltB+2P+yWpRTodZzE5EaAvH0UK5ea4W65WKCO560Cs2lnB5ks0Pu0wL
kRRfobdj3SUS0HewAC9GoDA6/Gek5SJ9+Xc/hYDVQji3augpuBGnpah7XzvuYtcV
KYAahCD17GSkrAI15Msnfqs65cUyfk1cQ6UAD5VVvHtU0jKm125pIjhBqjqk1wLB
KWzO8mqTMrmMSjiWbQ+rUDG9TD0NENje622w3iyKoxwj/Zj9AxmxTc2oH/S1jZYU
k6JUl3oN9jvWt3BZJrlX6zCKUAtm9URvhUNwidRBQVeCj9qbFT5qO4al4o53ZBFH
Ph2Znd302bc81g9UWDMwRb5dqFHMZauNhW8CdM4J62KltJ4VXm7870yNoFQgO5/h
DRFP3Yu2lmiFzj4S00FhKiP6WyKxR00LkyqneVxYjDG969/qd/+0FzVRIvfs1xdT
yTnrUSA68vC7RzvICZigcZvRNPwIvNljf3yjx646hDgVtFXNWFtpZLqhE+BF572N
bGmkuglEbsueAgQz+oDzAj7VAHSCNiZxeXn07z5IC0ysieJKP8OKI9aFf4RG6w+M
qeeZmsu1qAsuI9zf7oL6r87W80qUwIIk2c8MNET+ulwePrG0Fn8draISt/VGR8QL
POZndWWV1kjCkeN7ZfJOj7KYFO7QeBMKAmYbLiWwQMW0V0Ypl2t61c5b4SwxKQul
VZTABGXKgd7ovQ3cY3exNu0ip8oh295Ghc6yh2BBLJvpT3A+Rc7KrLf7GWbiPkgK
gDZmJY1y8nwl8V8zHkj5iN94T5u9hD3HM+WPH4NhwStrYWXuLmk//jjxpST8IUBN
hY6Oknj6V01T7L7dK6wFMPiAOWWU+1IYZt+89A6TYKS8MvqLB+5fFCdSe7zDf3Pa
06FOIHGw5XUV5GcL/Uv15Dek77FU+e00ye5IAEIiUsM7cHWxlwOIsQCszFWZLlIT
/iEJX7b9AmtkFEqgVksdOANAldDZghF2lwbFo+9rJ8NOfxotC9IKzeWT0lmbxieN
u+lvVSIRI6sqIYaB95t++hd7U0DXz1vZXf7IFL49Pa2Yd3OlyUfCKF3LZq3PJ47N
nElqaGS52mooM7LRyKO+aylASB3T7cV4zntivglx+Dn4heO9Swtm2zhmfbBYFPY2
Y5s9rqA03p1sUS9Ppshq14235ZqBvVXQH0egPV6BJAEop8XrO6Aq47Ff4YHfBF01
BrfEDepf3jf7UDcWwfj12oMNDuvhjrJVy4DRVVkE80SLgnzijLFsg1ZRGF2Ju293
Uu9z6ab7cf51LVRbBxxZGkepIPpRu4Oy/+uQzlIpnykpUjoc9WvT1lLO/DuHnPbd
Gikpyo9lLLxhv2bm9o1GWmOX6eQilncmZdSAD3hTSfVIVthThS/AmdODLY34OQ8Q
xUvWeESBYXUt+18bBcKjkmLujsHu2nN6Xs57mzrSbTiUftpyai2NhUh26Jw9DUim
Ny+Ej8vaEoiosGUEjh4VyOruEwP2BRM+A1dvScwozj0CblsL7wlMHhjNyz9eglo7
gA5yGbYvg+dSGzhiKg7F3HlwDELQsKisOHdfQgdLvF5o6CaFTcGXD4UnOaRgtSs2
uOg0Mj4jc5NllZYOkcZVIpCvU9YyS/8YIs2JVMtiUiYf7JGrglpGzhck6+y3VBbS
mSWXlnzWGh/S//JTQO/3jlf3ta5J52NAyNxAynNR2jRgmLFzLeiYxbxqiFEnjHg/
rE7yfjDLZgfNAJQOW/2TxTtRVKT5x3+tKUcCHk1Bk87E/IsufDBmYxnAE5r8sMOS
/TzOfECFuWLPRHeA6o8ipYyk1Rf+urgQ2WN053US2QGdPFD0FQENaWNzkNZ56gr9
w2oEBJfjIoHIWMKU6mpZsqVTIqs11GwMyT1eDYTdOebh54E5LkaUN7ihrFIVKC5H
TDlL2pIWd5TLD8N0t7lau2nE3aov6xyWzCagVMTeJpZ6aO9lkQZsrEVz2DBJ8rbA
kkb/f9ZlVcv/pvJKEwhsz3DNnmRgyftPFwk0IUH/y4IJSai/Y9ci15FFZMaxS2ot
zRCfin4TdH16ndo6w5LDtT+hwIJAaXO/+T5LiNmADhn4rDboQZkCaKp/TVYaZGMp
7+UkGE6atbiCFov3fBD2Cj0donV355IDzaA6xbNtZytpTW/azy6nNGYi0CdONbMb
fwIOfou2FbuqE03TonmGYo7qWi1CauxYnfLcfpwXjOtvSpvkcXfeNn+koCJqnMgA
RgHuEcD23zcfkN5O0IvfymhJB7aNSVV8+fskROWfDUIDQLVk7nFRIIiSkI8dA7PZ
1zQiB4INFj4g4YKLI4zcalIFAZXNS7lkQ29RVK4cvlofrF0yMz3epgjdL4IWsQqF
A6JaxXA9WaY1alkP64oM7UT+ABlVxYZ31eD+5IDcsSAs4AMQ47djq3O+gfD67Y47
UQxas8UAObQppDgsgSawxTg5QGPAWMqC2mCBo5z55hjvRuVGGn0Vztg55th1Yc1K
4wxT2gaWc8rY46NWHrEwlWyW6powCJ41ySAcs9n9/VbnvSFQ9pbc4hbFF1TdCvA6
Bm1h50LDQk9pFa+6wqCOHYZBraOVLpUf5Yb77drNW1O5McJApSOVhemwRsRemKb5
ggmKreGwcw3tsqfjH2nvdQ0XMP5wVszL8b3Gq2v712bFPRLN6VKrr1NSQ5EPxcSz
xC3f+YE/t10clOAPwXqVpqPi+YLWuREBY/tfEBftGUJe6qb24I8CzGljP/s/nlou
gQJT0BghnHA3pAaOAuzinW1KNiI1TY7US4Ofu1zQKW0rNMK+nkPewxYrCsHetSUV
2qoQL7M/O+nBXZOxN2sykK+yt5jzzT256kk9v+t1xXdgeFtTzc/QmmaCh5wJruat
JTItG7DT2OqumryigQ6AkyZrj09Az4uZ/8b34SGs8iIYkInh90k+JAb3EHDH/Khl
mB3GwofPAgF0fNJGjc/Ldl7RBY8XqYiqRHkfMl9MLmVjBd1K6YmNlA8MEpTHfwKc
03EXHHh6RUpNmlyYzSU/wKBm3eL/KOQuxs4Gbr+GQfmUK2P3KV9B5tMolXUPV2DM
aemHIpRK6wOygFi65pVASb2dBB2P/0rSmU26+jNQ84sUvehxRmChEitNqmIKWI1m
61K+vSbZUAMnFtUngSnXm0wE7TNt6KekFCqVGtHuUxjoTh69B9RUp3OileSFzfoM
DQxQhRFrtBKnaz2FpNllnW1QJLZkUqFBw8qFZocHzwWcZaKcd8VpeLXWqaSEtif0
ztU7h3jvw8GRTMusxC1jUIxYznznECuWd7K/tfxP45qDT7w4PgLGh0aS704zcDG1
H7HDNBGzQOFZPcsSdJvD+q/axKvLrSW5m3UJn0umuWFwQzemRCeL2GS4bwOOf8VW
LgMgAjhMQ4WsnJHI2eh+ZW0NcMGSQGgNJvapssrJhK5E7HkHfQQHvGtrPJc9dw0b
iH1VuC1rVLOGu3ghc5ouJliAfAQgFj2kT5rzNdfZIeVHgacMqJg2vHuEWuO5KVMR
pHbZ6bFswx9f9oAfm4EWUpITSgbiQZXuCzr7a6EMID5MgV9UKbd/jKxaJaQKyQor
RhQoSMhtEg8vXxXAmXHllZDb8+/iFnWV30ESXcuAGBDCtCKn5fTfP/n78gMAhdQb
tk5mpx9JuUHU5dn1pm7C7JWtQZm7y380mp8OXc9oziOURU7gJbQ/WQxpKQo+42L9
h9qm+sMul2Jc+zbR2nDn0jxR4DBrroGs2PY/U/pGXR5pH+jiuCmKeROCPxNgrYm/
U2hZHoEYaCHOa0IHFY2dI1T1XnXxAYhlgD/cm1ihmAUO1E+oUb8junz2T7gTHaqs
9pQ9pc67ZY+84HOqEs3hI6EHg3UktsO5anKwN6VpM0Mc7KiBk3Vel/M4Z3RgSWIs
tgCrmkuRXiQD21YJDlBd9TxNwxpQ0JrEDQVxbwN1b9BeYvwR9DglPuDC8q737Jwg
nYApFB2LEsNqPUbtyU6qyVhfKOxVcwfTYtspiLVLFEZY5gha3GvU0oVclrrVlvZU
rGxpU47i6655xVkWTE65CEzFL3tRrs/mSyrC/vKU+WsXAU+Qojt6/ZG76hqGPF31
WxwpCBDCPL51cmRyx+MukCJ8TvbSg6W3+Ey2jQ4ArEw9wTd/iPOHQ7eR7a8vboY6
PRt+vlymkk9we2J1WJaeFu6HzHJBqCE73GjCF6CaI5Aqram/f1AqqqDi2nIfZMmU
9ZpmYtSWZmLCpCf8N5K2zrLvO7Zw0NH0sr44aC70fD2bTrbcuZUZBUhtWXLhhuZG
nAIQKGMvESrv3A2Omz4PIPer8apiEtkBxJG5iXPp1ByEC/9a+FAK4g7pkK1BYpG6
Nq8uQKhcbEbZjyW4T0u0Ir4VY7y8zEBDlmg9TjBN2xcXtrCTznUFZDsQAApt7RFX
um7W4MUq2hOILIUodihH3Cs3g1ooazktZNPOaCpWDYiTN3SlhbUMKSZAoGzg3IFo
J6FEWdcb0Sy1VRKWVz06tJQQCpyqWhuH8gUjWK/sHrgfSVhZuQBToxM7SNWqJ2Zq
JhZFF3FQeXHfZD/z+yXVw7jD0in+qyCeYY/bRPJYbLMaiuKywtHIJ5G5SHf5K4om
3GY81qNTNyub0Q1yK5/Zcap4+hU+7HgwclUNZxxFPeDAjG82vEyGmBT8xPprhSNC
vTM1epYCadsIWLuWxQ+44zpP+IBglwHVJFrRJKXdJ8LAAc5TKAtCzLNI+B4//5h+
tMC8lQ6jTNdQsxNiEBwVwZ7vEGPW8Ec/8P1vb0plt7NHxX6DVX2pf1+hyIlDcANE
HZ3EouTaVDG3hDVM5sb4eOlhnZ24QXUe+BtmeN9qbGxW5KxPlBm01NiTu7EFlnmj
HDyEl9OZngqpGU1D//waNIT/egdum6Ii2mVzIcKPHFGfd/T8lIh40Inm+0jiqLv6
7IYrpZ85N5sdR4YSJyyKD8mq+AuXHVG9BXzQsKSlHsInr3oOpdXIu4sUE5cOWIaS
vHnPWG7637ruTjGh3En33tPbU0KEZCDZZLVK2gnIpB1AcKyAEEco1TPBKqxQkDFL
4+fwWClRv43kvdDCk3QkJhe3ShkW5g7DrMw7kzeBbdTtccb6htp3SnvCP4hUOewR
HFBho3q0vOkp5NbZDsod4pJnpacZmp4bw3Cv5zVfRn/6sIcEYOrHoOidSSVDWFpw
/33PXeirIfbX0bKzuPuT5jOwtHSBdjU9UzyLvVwe5EGVjLhmqW4kTEAQpaOq4+ym
BrDgUcbeJV64d9+zR3ZyvOjXX2RUrL2JWkBKBmLa24iNNP/AQKkmBXkm5A4xYIvi
mtOGb02hoO2QYBKbrtVYhpkpdwUnxpm36HCoSH7Hv41eTwCnoV8rmh3ee9vRxP2g
hV297qingQXAIvdWIpKKBPA5RHI+zoaioqM9rH7U2Sg7EDiEAV3SXdfM0/tMFmhj
RFSVqEVxJOcBXeaHrRui+s4l1KubhulKzqtpC0jyViE5VDllhYkTU76UvEWxNfJO
dLOgKPEtqN+uf0MtZl11Y47iT9j4pNBJQfKRMuZbaWP9cNp0sB19vBiIftxQdwt3
KNBKDm4yfWn9HJXPZFNPFD7j7307EKRVbSxasG+V/lb7oNIa6r3ZHkrbLK4+vyMR
Y+Jk1k+DyPJJfFaJxxgW5UslI0ICy87jK1MmkfSjqCCJYYCZqGd3pkpbwVyJ9INO
ak4oJahjyyPwtR8tLJDFAvUxrZiwRDrqZnwdaneRG8oeowxnxlOO5/kciFxOvMkG
iLvgTTwHEEzQVsknU/5Vp2tPC1HbvhqOIJrw9xmTrfhMP94lcamPDGVLHVzjhc7q
B9UHqnkZYdLYugrwCK4ro9v+ZPHrW8ZvOXUSLyWc85USfyTi/LGc6n8R90wLZQw9
ohur1T881kHODj8W7gf3hWj3/aSLmbVbh3Id0pHmWBPkQRL3NLA3hwFiVxKfXK3W
ivBD/xLCp5wPe48/whDrI2/YjxktnU0Vbx0T8WXv4dC6cjS1u1SrwILCLlUELCOD
dEbIno/LqZYRgX1ePx6mLpQbNiHYkaa2zcaGFtoiOsrA6Q3sNOkeBeJVYaV96Gmb
VdleWIWyAjXgvB0SCY3BWHm0Vb/zolufwLCI8xwRNIbWCgpp8GA4psSPwjlvApnD
DKKcTaazdxPZAY/XJWSwFsmTtjMEypwTF8CXu5I+bZNYt8vG1vILrPXM+nVV/TN/
c9cQUgBEiLOgMB0MRl4Dz8NtbZtGIKlq1ozzb3sTj4nUf/2Iclr3tUf4okPhCMvi
P2tyC5QvdV9+JWRTToLNorOI5rFh43WdWlBq2dZr+ShY+JALHVgsMXSmPqaOEZLg
dgSgMrwY88cMAW+2fkDsc9nYDhIqjRvCPKHPtZE+wBX7Udl30VTU8I4JYq7cNSt/
26lg/TUEH5rTImOepDfLafPx7OhLmyUhpZdMcP47S7xa4nipbWGvriY+BP16Vy/7
hYLfjkydZm1HW0vfFQTuiApHKR0/B3M+s34h2yx5a2L0rNt9RqkWw2JNScmWG80X
PWOWnsYzQVMle2k02EFiCF0vzqbCRzWL9MmT7YBSvjpJASFp8UYtLvzHAU4YBx3A
LGDbs+vYrc1/8UV9qO7N57nRgh+T0ImAqW3XaFNABdFO1wsqbGJFId6MFiWcLfvW
p/mzggk+7uHj45yyptLXtCRehRUcSdFgJ427sQrbaKS8mhq+pL28SlgH5MnrVtxf
OTd/xmgI6oQxtasCcHm5xSnBj/6SAFGTq0x/ek1nMN00jPPPYTUVyOAYzEWO8+ZO
SvoUTnsGyqgQEx3EDJYw3Sw8AGgFL8ob9Rz41RCXpUkLjQ6UVHTG+e512+B97j17
m3IDnboOB2fKRYzFdbVU80QmD/gpY2AkEEZD/ztiD6iT+wicMLQ+2Eg5Ij/G50TP
Hu0doZjl3VCBkvjCdlvqkflMI0LXuq+Us+B7qSBDOXf2aa+f7xE4pOlNE7kez2q+
2EAHmsPjNZZJBLRemj+F88hn4LaSpoeD/h0FhuiKqB+zjyqAEajxsxeBqskK2rvg
VyJJnytm9Z7g1L5OYI5r8OrhwtxSh3G2umo5sfVP9BCjOf9BoPwMBdQpiw4b3WMP
QDZyHJtmz9F8ovxpZWa8v50hbmwnkGawnm5ao+7usbkAB4H1IutQp9tFbtfp/ipr
iRJzUGPV2ioo9CC2wuJKKaeviloqhyeqnL4fRI42gocfRJUuqAiSuG+ZTXV2u2Vg
k4MUJU3HS7vO4Ctu2VfDWREzFYRv+mvtQjhLSqtZxPNH3BN9viFK4S7Sjrxh/Tm7
S8njNKvJTGMz16mFfLb8iz0BNBH6xnn0qe+Z2gT2Buc7v8rpTHEU1ZKBBD9dAlfM
EsXjEkj9ikkymO1L8ItIvvezf8m5vKG77kwUlW4YQ6UZMwIbZqpTsqVlHumwzY9m
0Sn45V19Sx+7QwBWiVa38KlIRDjWfVZ/XIATDph+nuYUOrW/z6qRJnpfoPVK/ixC
MXrnXxRgRWXpoS4/YMwHNqTVuLzl/cfkxmdD0Yz4tXo6YW/Z0ijJSHoRF2m71A9s
sS6D4DpoKhDxGwMmg8DqOsc3XtD+Oe9B1nGoXJ1MBjeWZFe+h3quPDOcQVdIko9o
YHZ1po+yOKhwE1rhODhJs5xnQbCbDNVgyTN0MH5W8xjKPRaXZqpugF/0ICtMThPV
sihU87fFd7ymb+3msssyIoNFHBVRbKloOL9v4jbYJinzCj81rWEIqQ26cPIn/l5i
zE0EZ4MQ05qWDfTgX8JC9o8RP/J4BXjiJE4Hk9QywJKXAtfDHcjqavEPBaSNevRm
ylUA3B/UPwwO0L2+ZhovZAGcW30Syto98J/aAlXKg08S1jxA6q2PlzGHZ5kxbaHC
AVmKh26xFm/0VUyUlV/zt/9yL9Uu0jAkn+43QtxdgUiEZ4m9vv3vYMK21AJZY6Xr
7O8w6ucK3N0SX4fdLQUwtnBhU23AqjXG3w/FHees2AjaEbopy070O75V0wSAjLVW
4x/YDZZrgKlMqE2Cfw1LslT5f/lfZHQ+OCP1VIIyoJyZGmCshkURQTw+i1TQhZtG
vh7MTnndgdLFIdnjKdx+f1dsAuEXtTapHLZ7Kmmldvn976kZ1thGIAzJdQ0VwcRJ
zj7m4ukiEADYr7AzsMMLPPe7v2e+H+NBajovcWoVLMNMtTIXDnBjWZdLFOn64NY9
3nxlCGoxChyFwJ2h2qOULwhvcil8qym26jN6SfjLbdCgNRMrO2Nm9Aa4R1nY8Xu3
4GWakJtfRQjMLJlbE0+RQfIsMkk2ic16rRWnCXAaYpNTaEqe4WEFNlb6M/OQsjY1
h2Un/cjhn5o5c8BdntM7K29iNia+P6rEFW6OA2vAC4aM7M81P43i+ThtXHXTfGTA
ILcUm9t3/e3W+rBMzJxUT3MD21Cv95RIahvrMtBlQLNuavxG/gI+h6L/pPAQYr57
jkOGoEwOO7q/jUDyQTHqdFgat4s9BAnkoZYQCKF/9gBSoMQJcY+PrJXPWbWwqstE
FnTgI3tMgvXoXBTcmpx7inf/p6+6zRWE/Ng1gkWMWOY/uLx9bXmwZma1Q3guXolO
TbU1D3Hii/jX/zotYExozk4PKIuF2jxS49jneg1B+sC8MmgJhtj9EVmopHjB3BwR
aq7JgijjYZdMxWoqeGQvmfCybKUnhtcMHclSwsvVJNV1H4EfAaJjr2Ie+rGb3tE9
LFEZhkA7QNNNjbb+Pjc2B/1bcXebRgTlDj0rrUd4Sr3LyPKle48gilB5OjsbqlI1
p8qCrd0wAwR5/ZMegmjq8Dn3ly3lKKhyfyrel+JRMhMqP9xlsvpeUdXzD0nLbMBN
wAQR/jMr7T9wtz1CRT1Z4EIWZziHeluE7Vdycca+aArNhfH/+PyQHWoLc0c4eKMf
pxXU0Ff4bZFglsVnS7mbEpUob/RQyd4B8Zhst6bHeZkRrKF4+3hJ+9RA+RMpfD8A
CALCtn4TRRJjbNV/h0y+i1+qn5qkENxX7PMrgkhif7ZR/NDyAGHIqTZhz0pzPiX9
nAA8p1j0NHPNE/9ukD8K8EzwYIju6U0LFIg5ovrD43r1s4NJMjc2nv9iuih7gdws
wtBTERSoBJcgJQtK7gp9Kc/XBpjOn7m2NoLCOZxqhhbONg1e82DS/gljbNHmr27s
L0/A4XbZ0c+CqKSPCteqKrwScMhZNoWqlj19MH5BsPbh16U0t6zqGOY9aOXDo+R1
e5NnPkjcDHk0HY0BaI+3MvK4SyrQypTXzQW5zhTsrb5HcHrtqqB1F6zBKDgRncYt
QUCa4IWjSDyQUCPmfj+J9Xe034P5f14bc71MT85AxMFQbV41jWGM7jJ2EaR5K4fC
7C4l82iu4mF1GBr0ata7q2voGWp4ecj46lTh+hCcUMwWnI4+p/3kHJU9AyJIIgcK
bKHxHAMLjo5pNreYUk+V/t+d7+eDbt6hjLPd9U2ayPyvWcoqEennlqM/ofpc5De+
OUmkTTEExXCGulvP8+ndUEuq+0WfWEQyInFvBj4oDKwP13oe43HRvEXzh/goF1VN
9+y/5yJeUXgjV4IevYhX7H2XQKbdR8WUln2rQVffBO3L/TtnJ1yjkKo+LSeERn34
cyL0b2I+PrGtiPCdnIHjP8J59l4D9+KbUGsUF7iHeQfatkuvJEMHESP5G+ARrPDU
D0AFrKbeVHQiOEEmMM1ef3KVibxR72efRWVB/mF8pST0Ntze2zzwdi+h5kLmc6hi
KJQkySSrL6BVqULuFo4sqy1eGwAcflvRb0hX+UC7OutvgMvnvu/5YivOciqeyUWS
N72Rtjsr7tGIYAmw/X8b/EIjrjgEbuJ28R2O81HSv2SmIQQh+7e0dUwLrwRW/p+B
r8WnNhTCKqBB21LKIpA0o1RaL4DXHKfe2yDVyR3Z0FzckDdBbpA92aov3K5gJkl7
NvGIbzkj8ScjRBDXGjSFR85DuYzYz5wzlLaw4jWKnHdA7mjM79ff4iFNlZ7VAOSG
hYOSr8WwLIxa4hJ0VMFZdVebYFIilSopR37UF5qudeh4HcCtFRiNcBpelelIoNcT
dT0/LOpTkdcIBytLnV34LlXlRts4AJrXS+mf8mp3yo09CAWP9zuWk64MlPi6CQLr
li+p38XPdxkugvuGLmjbW6fw91JaKNNCC4HL008m4YQM0Fds1j50PS9wMYWu8cAc
ulWqlcrxnEYRvdG74y5yqkqt9w6D+Qxepw/Gair02hAaoeOm9jUczwjr8p0WOaTl
GSb1JUYuomvyiGi6cSqMqQjMLNAuGSdUcAO4ZD5jRZQjekiNshhEhBQZrBSdCLAK
b8Cs25YIz4xWhVnHWdJL+Pct13D57v+rrqzbdHrAx5w/CPrNK8NwU4JUBCES2mBR
vvwiiKb6CothysOHNkobqfavAOmY+6P3RLB1hX/xO/m800ZOFemESNGJ4eY/zjlQ
LGT5Tc47SKBaoP7/kv74Wvix1UJ7a61H0mR4QcJsGybZLfFM0V6y0hY80FtmSilS
Uc/HLMiY3cSRnyqvESobZrEC2JRetELWZXUdWJXNSYyBZ5SFzYOV7pNI564VlS7m
7rejidnVMqEBrb3Qq8OfiQFvtqVtndAqlZ/3y5yq7gyEk/uH/FcByOc8W6G7MRDI
MeyTcgrIhiGsvcdd3lqmr/CH/R5j0pcwFzLqwznY7lWP/RCCrMKSOpPUs/kBdA78
fTt/R3SKzXGcB4eTnojHH9/0gXGIM1aqOogvJBkKOXP4wdhKck4CnukoSaWUsTYv
jtew12uLQwOrlh4m1SEcPL976VgLN9A0ShmkE5pMj9tClUkSTjKOFkHac8EG29Wl
qh/AffwWQMCc0OE64Cep9EBRiLq4m+qqMLpHEdQlc9PCew23hfC84IZfB+iYwpUT
btrRtKDhIMY/5G6FRIdBq3srYVApSnmt8XiDESMYdz5Vde/K5YplKV0I+rZi1rRJ
wrot81rYuqqiAGPuZmTtsUT1BjJwln2HArmT6L/muUtaHPIgpKPKwyfd7uCKFQMo
Ubwk6msk/wQjsydQSd58O6HTh0WiWB17nIQjz5P008tVxoH2r36qJcIDl5H7PlIJ
Oo5qocvu1rh7Krg+puPEYmalx4E2rBo5JHcZxYJBA3XYcY7YeLhgKUGCzd3ThOo8
Pzcw9wizx0hhmgIaGhYIuc4i89Sm8qOQvFtFwjTxUHXwXFLgdJtxzQ+HHSTC1lwz
6wxEoXI/BJAZ/uje/mL4f0dYVUE28np1mWyL9oW5ox5q+ES5A8AutM/FKSLKf0qh
u9sLZSiDdLnUeethqouNrgl+FMT+oS/MteCZrWjJS1c3dd3EMwzlzBY/RAAgoGRm
WlZS7G4pghA3rHja/c0+QXmO3KmGXpd3irQvCyoeJTL5PL3vep5/n+K6Bt8L2UJi
OHIpDZZ9g2UO194elXutrC1PDst9gB6d7Qt2FonUP61oEQgoUDkSmu5QmOONLRrd
D2pNg4E+c3Mmnf840U2Ek+tAvg31MAntS8PDzLSaetix9TnbLku70hgqtBPVj5BD
oFPuIKNsMS/CWEVHTv4TVuy4Ho0wmduJ8DYHYWS/QqLFPmiM7P6/opder4ca4Pfc
qeB5m815mPNoWL2zQt6h6SPpbjLBHVqiW9Id0YxYhvGK8F3syeIFk0crMH0GeEm9
FBRbK6dQnQtqM2gd3Fg4mJKi25dQgx6yQGs/dp20MyttTSYMRwE9YQcB6m9W9+yK
BYVNcmRTvPsaek6E27Im2Z8Gg2Tez9QClj2SVlE1bz3gsYb6IR0iu0Hsm9b3uNDt
S+lbdVx+azhMC+YwLATdyX4NOUwoVrmAg7mLmy4s27gLKtTtX+4991l31KShklyr
R9JGEPtyjW2vVZp8ePUPJSH34SAtdGdxdwW57v8OcSYFYZ7Uz83p1jvwO5vu1Rwq
mIv4cAO4XIWBLDWxannc7CLHhYp7UJTNBkK/YfEgWo3j7S0Nfy3Y2xqYyA5WYbl5
hVgeqb9PJfEBYiC0685OBwvbZ8lvC0XxTIWyfbptBhePwpn50FImiWBbDJ61PXPL
ul7LozlnuX1+MG19NiCK0hR8iWrwQg+/WQJ66ghB3t199y5OVnT4TUiTwQj6OZzK
Ag8TlQCrK/QyTmB+xopDi/8jxOYlzlwWPCKtHJdVEpBoYe+ek/ec73qs3CgmcInI
XGFHadHoQckxfL/N+csRUw1APQo4U+MiFtkv5tMjJZfjCdT1LZjt/2cuBqNSEn75
A7UVwVqHhRXYWCh8r2B+0/Ypl3a3bu7tPzBh91/RAsYdiJ2WSkT+h2cV+0WaisEq
420IdA/f6zDsrfCx4D7ldvg41yXcXhprQR5qu24OrA7LcKPjobn7AiQHLaVENJyK
nCWHmd2DAOJxpzn4F7ULarBXxQWu2IWKOThmwACqkNhT2OEmACYMWKWgkC3P0oXG
tkOQmfzbT4oyWTC5hMk1B3bSkjpxp6/8jYLoBRFe9PM0aYfW6ULPsBZTkkUr+KWF
re2pT2VOOSagc8D1bBESpdnHcMi9DXpP7Kpl/XP/nRMr6mW8czHDjk6wynKDk9nT
O7Nfc/nn5QKUPpg2JRZR9VONrWhOTzqP4EMJyqhy71wYHclYrh3iE9BW1fz49Eoy
PS4ZLqJ+CVed3G5s9Ru62FXumtkq7PF/NClrcC5UUiYmIOOR6xKCh0XKsfSWPlvq
5zD7IdSXUFtUJmtZc6p5riIXz3eTW96JlthJt/xAUiptkDMx8leXsjoG248qr0Br
YjEWzcYynIh6wYavItqtNFJ749iq3WgshsfHmB3zKrahTUh8/JKEOTkl02uScnad
ozH5iXaLk37QFkiOIgIJLPWrD3bB02I6+IuItZlXczS+HXuFWBnHfT+PuEv6Yeur
93Zu7YUCQtNNF+QYsudxPZDmDMMKAHDZ3MhxTUn1uhowW+u+/iur8lhThu+POQZt
CrapL/glFPOl2BrfRqI+vqubr4Nqcd/QeokA84+vTJ6aPzR1Cdhv3sCU6NrtGF9n
kjD4nkzbHrDH26OiBk33HLnZslb4H6tHULVy2Gyvyx7MIcusyaKF+mDXdO9AHyb8
OiUHBjdjbWBb3gxmOhWTIM6zJgyylLrGZnjI5HRhu5LSZnluHIUUr56ErgGCBmUO
7CjTC4ZQ33ub2P6JQfO/f+p2xq5WzH1zpMPMvXuKsqeWXF0JMzxPzAZ+T9r3h+it
m9rmscXVIwrbMIUlS7SLhbR/TCcs9ULzp54lR0fmJirlUPeDFmj2BPKBeyBQy2R1
vLOfgIzYZ2dzigckRcxlMnAzCuZnmuScUla8RUcq/xk5ftVPrKtDS4m6Yw6jrSNF
JA+FLuyns2M+BX6t1vGioCSP1M8SEePRYu4duMCuPQJvIjDfwEAQ79BZpIoMLS7c
IJmkn8Zh2gwZ7Iqtuz2PNuli6rnBJEmNob2t1sAxZH3vEkfqr+wIXthB0cH1EUdR
lsqbjL/gH5sIlgLn6WEYF9KgB07T2fIkA/dy701g2hEB6fvretBHF0OfNItB06Ks
+5tF6GO+P4YOWueEL1rXuNWoX6OEN5xt8LOkhw6+FTbgWsl1JKywL0LnmAcx1bJ8
K1rpQiePG3mfdQ0Kbq4Dh2nbIpNl+B/2H4GKx2V0xrAjQ3NNG/PO8VJYgF7qk5nY
ps3xCgp4gitKlOFu/HiwmZaNEkVRxi1A+86Rdd23YRFTjk0OylcQ0XhmPR64Z/gU
YKe0vr2Ua/PRZxTkCpvoHIgGRH9cs77AR92qLCk4O/6vwUvqE2O+JjfyTbPsXqjV
1VxbZ+JPxz6LQlpae768O06wiYuTmVweY44lN6xvJWb5RPov5Wnbt86R7FGfLu7s
dcKuPJ1z2XlY54W7/i07sl0GCrNTQIbiZheFvvfJif24Y++meC8/YI3lyZg53ZQS
HaHMlJj1wMTyZi0WoeScjuB6jEoK2Q6N9rSTiSP241AE3JuWB6snMITO8ED0YjwP
6vgqxvpv7U4PSelHCR6ydnwCoXfexYRAysncqcAbR1nlOCmGpKT59YzZqZtZykHu
deQsWyjIWevwOw4gmuLw+J5mEz7WDMEV8SNLbq0Y3W0nMfu/AxT5mtvhxd2/bX2Z
/QE2SXe8uFIDAqz0/Lx3f4ukRSiUdyZLCZvLaiZykML39ePGbUGFJX//wV1LvKpK
GunnduNR8zQNoxMJrQmxnfY2OUFzwXAkr76pHhd1bfBx7GUVnV2uYClPEFxnY8cN
lfuVqcaSijbz7dI6d2HmYQO/QXQ/Evt+a2ozu2wXYViHLh8mpYlr5Kv61xFoFBhy
L584nW0LXA+dO4c/zpx5qBGzOP/1Mi97dXmhKwzp0LOSON/6MxfLtaq/gGIpAiqY
7/pfgeRZ7AR2DnBDTa00LrGi+E8td9AyHQ6QF9brQZKulJ/pKfxTyPFwro9OcAzi
CSQmHmd4E3BtNUL+bUSD9MCdC01lMUPeRK7AK9hK0TdpUJc2WOJTPUk625PBPL/O
IzoPTOsL1I3LHP8JfxKmeEezDJW/lZQSkqDVaU8kUs/5MiOIxe9eXSJQGGWldIxy
XXDD2AbScQ5LbOOVNl44cTgEb/BLFySh1peE3PrTHRwAOGpqyLTFYn/C0vAnImkS
CeGh0s96jiYx3CKqfKtLSElN+qU9d7QaLgOeWNGrKZoL81YhdVFqPAFFamt8c0qq
yWX3Upa7nfo1BSaDxCmUnIFySOHEu+a623Cl4ZbxpULi79pYdGq2gpuCu+d7fpUV
U3i2mJ4XUwmoW7nEqZFUF8nHona5IUYjPLUgwN0POVsn09eHMGdpAmudk2bLo0sR
up7J+FckNJuEeZhInIK/Ftr26BSSO2v3yMO4eha8y7BP2ExXiVo8OZ8I20yDQLBs
wcGwpo7LfE29Zd+n5UsnVGn9PGpY0XFxHvahBDQ67FthLIwsbChYbuzCWvSbqipv
dgcEfxa59J8RhtG+UYC/roXTfkFptVdvqOSZKP9XPO+5j3qtRJKPl4YN2va/jzAF
Fwutfy6WK29fzhOZC0GuHkRZpHn7c0s4BjBdwp4SGLiwWV1W8POpZ8mJfNTftRVx
7as9uB7lKXYD3j9v5JCUmXul8UCMcIVplpdMUE3flwF4cyk5z4Pu9B5Vdlhz2RGo
lYkHcG3MgQArWNS8FvO4qdN5/59AlR/obt679W4gKMDDTBnV7vlfz+BlqDHjSygL
mcSxNhCU/8NWvM0J90yIfJ1Al0Gq+2D89bAM+JkBy74GxIgHGaFEH4vZSDMVJCF1
CjJaeFWZNFspYhtp2Szscgsd6C1+ss71sUhyXya+LqJ7bd7/xphLNWRjgDFAuj80
D3O0p9OAVfQ6P68XwyHcS/uOXXz8dDf+9D4IaQ9tvxfGihmJm62REfEn4L5qAa2e
kxbVI6Ff8U+A77gpu2VwtMuUFwhqKIoP0okmzDk2DIHb3tgqo0qlHMB13UWCQ0/u
hCZH88R9UrAxBP27Wss2TEoZcAeXD00gzEB7NgstK+xai4mUa03NpF1MXS/GknIg
RCUo/DocDJKdXR+maoCYeQs+nTBP1VfkNJuY2JiecDiSDVR95Rga1LuUSP3yOncW
TL4yp3Wf6DYtOJIO2dEYqsqqhjrwqHxUf8zTW5gMd3qo4InxS+JXK9vlu27USaWt
B+DSVylw2xpam8BABunfd9Soz71pDrqRhNwmwUd18LNWnI2GoBvfmSPXx08Q/5cu
lUuOQ1KiQ3yrPp/2F+ZlD+wtz4ASI4XqU6xNScvRAJ51d1M/cnCEWwzlxH5lN0Gy
MhvuFrC7tgkC4B67l561mAW7kN/TFR3ylRHQ/k8ebjCotN5Nxz1LDLtgtKWlVgaF
rU5Ypc15Qhiz6l6mEsMS5v9FQ8Q5qCI/K/71iLmxTDQTP3gSJvPYGsujbH8qhuXL
1nT/k05w3Ix9mrtV8mrPN6zQp+Nwa1xcWLbMrCd4Yy0QUkUMXNhiRrrwHRbKM9Eq
Uy4un/IDQx7yJwBhWdOfja/0SQIiyNuf0OBx1jgsTz8GspNvOL7AQ9s1BflJKWSo
WzRUajnZLVXsxNekCUWwhGsgNfOojgf3HfQZuJW8j5O3CYiKJzzdXVCEaIiq2sx/
yF60mZHmxC7wrltxrosNxSIgUfRGjzHVQP0lEMQZ6qlIVTP9wpvOkqogIY/JhFKu
tlEeFaBkzEnhNL1HUKnxuGInPeMum0YodYhZNdIhV/Vz66c8en18zyulyAi4voYm
mau5OYgWk/FrnA2PLk6xjhwwzMzrvyrKR/0YviXtSOGWz15ObqG5Yh9lOHilmSy+
mSlbv1V/Xc2dMV+uDhJ57LWexSEq4AFcXTq5Ya66jqbSqssneiba7mGQO1X4lg6H
sg5olzZQl4IyEH9NNB0Ql2jqQzKg7MQsEo9imQI0w3rsrFHW9OB0uXjRZREsTorp
jxpOmK3SZ1eyS3CR8RTiwGzGA57IKW4hG9XMl7Hk9hcDpReiV7rJ6PLqX5KVepAk
eE31S6EknebYBCYP7mNWzpZS0mfubZ5N/eGB7fljd26IWU2xBigV0jXLZAW05Vnv
YRFqyF2kP0rqnv7Rhw7kFuF3IxPo95Qqv7jEBkIV5dALOlRdjW51nl9UA6xxJxRa
n/l0mf5S0OPtt4SGj34BWkmsL8LbbXt4l5RpBHJrZhUr1dwdcmtos4U8Xjn+u2Hj
cDqrMbjfwjmhfkrW9QTxu4bJUfQdDtFGZ6en2vNzMYRZyIcU1CYPpLcJPye/NtqG
Mq8v3XtKkB2IlMlNQUO8J7jUPb14kXGqv09Uj5yv+09dO8o5WWx8gxVmUrsTtdh/
fKG1ShZLArChLFtVYiucw4Wq4MEsXhAvC+TPOa5IPs0rdtMEZllNESyMThCFfZxO
SqHpKQSa0/aQ/sIcc7dVD5cAHoyNNUIlk2XBgm6JtAsTI6jTa4xoswnhgvF+uLTq
2yk6FZJbmWhm1RFolK0GyJclf4t67pl8u2cqaV8j4z4mQGGvPeevNXuVVnDvhXCm
6dgAg7bTD76EL5AYfvz6u34kAvpyfswf3b7iVbNYJrEhn5teePQiDJZ3iAYwcEgP
JO2qUpNbr3FAjPCo3ndZRWzmQv9ALT3hxfjlHKkQuoPLCi5BnMUfes164mR6ZYHq
45G3+acGDAjL6tTKpnTCE1qf17AXU7bROZz2MnqnIAvNRkXE+vXyXCCgABI9F8oT
dw8+z9r6UFmv/Lx5J3d5VKWpX96vrEo4DSupdGO1rCWXgyhwrBzWvDsqFk3wgEVF
CiqZoLVcV+x2cT0mudlZ38YO0SHwyZKmzaojYaBBv8pguOQ8YNWmY7IxWOmo7IZ8
RwOul0T64LJ8cXYLqp2WDVwuHqZfOBn2LlkfrPhI7T/r7XJ9ojzyF4dQjHq4Z8sJ
Cajjg3QU0z4y2mVPAofxHXWEtH9ysIHlau6765QbS9TZNtoq7rAyX8Q8Scywodq3
/Tp+z/WMbymHhg9qDlvWKp4puT/taxu4vt01fiWaJsyyE0HoB8DN+Om/tDBVMDcx
OjTzwS55T0xW1MIrmTPYf8wxiz8rp9zokJVp9Y5VhY+pQMwYdy/eW9queE9mX1Vz
+h/RkwClxKH2q/2vV5OnosG6k6KcZ1MZfDrC3bZNjtzS2cKFvlQhG5467BPtOkgy
BVspW9S5oOZz4emhQTMSO9xotuXZinONJhwGw199tcWNQZ++p58NS5TFKThY2QoT
Y2cITNX+kfkfVRfagP60cIa1xzbA2LIQ1spdF73l3ROvjZtFupC3V0htYqJR8MNQ
Hp/3G3Q0+8clQu393Tdn5u1PIyAK8EHxKy3VQmqkbF2lkPmIZ0w1u1mrbGSSP07m
1OrY7lEO5QXMVAuYSdUUM7k861EluyfFNOsUhukZOVKCACzOVRtzSOe/uk5W8Qwe
umqH9Vur3f/VHQy/uAZdbXfip4MOFWW5b1ZqAOsdDg8dEBo/9jhFJYw2WTnZGxH9
w8AyWEkTTiQ297Zivzdu4B/byxInH3QNChZo3bUMGtACAhfjrNW9xoNhaa6WoL6E
lEHXmZkfKPM5TOxb870OhCiArrpUHif7qHbTKppCsVjMnWj9FXTF+vdfpZc3Ag6M
frPv1iu3tIlRi9vrFt7L5cG3vKPZ8wN/xwTKC4P6n4Ec3Tkh5+kty+akbKIjC57H
KNJioaV1mycNzsi/IfmZ5zAmzDg53ovqtbwuV2W+8VV6GhsXXjbo2jzroWpaSC/Q
ww5DrYp3Impt3IgfqLje9TDgfAoBGLNSgO2KkEHZXuI5JbL899+DS034jJn2U6B9
hQ/GViRoUfExnIl5RREpiWSd/ZTQe5kpckVFIj4V7MY8RnlgZm/bRW/qJ2/0T9vE
N1K6M7WZhCcGR2GXsoBLOtMig9NFspS6B3HwXcpxCBIbmte89/Jx7W3g2Kf4E42u
LMAUTm/CzJmwRiwF2/W/oT8LiBI1qL26o1qEy6bAVPubFrJcBtvUCEpKTZa4s1dz
RJV+CgtkGfmvSbQRxp43IpA9E3s0WSb0aYeH/EI9qJZyQZGm4BU2MlEN/V4oGh++
nFCnF/zuaBwL8uvyZQbXG+955yuZECau4uAx4uuYDZ/5EljaW31z8uKKnZC22tNV
wsSiaK2BAXvRdvB+s8dKH1LFQbJwTxyRRs/jb8/OtBcjDLvzFVd2ZTsbIIwQ/3xs
IVQycGZYiYc9N0r5c0PTqr2Tx+hHZFV6kgL0XtPjmtN4rph0bNzhi+ASDDHVmqlk
78Sg7HicXpPd3dfAo84D1UHSdCPI9fgLF6ZIE+mFXxUfCqdoo90Ap/ioJGTiw+sZ
O+Q9B6THOogUfjy7oOVnocU/kCMc8uZTDNDjDVoQiqRHeDjYAEtJldYPG+iAMbb0
pJyjGf5hW3RscKSb1lw7kkELpIoKp/UgKIBUQtNjPatjHNWwS81lwGJBVn0w0YV9
RtHcubDMM0qDe62zp91HA/2vvxQHhmCrvz5XMVyTYLaIdKC1AHc1FLShHaEx0fwE
HT+r5OKDT20L+XJbKrCuEmKsfGIeAt0aiWDwXrg3QhESB0JrxBgqPzQ7iT75XczA
Grd9d0Eh8IrQfYp2dBFVpcUQxaQe2IZnfFJY7KXPbJJa4+sv+YLxWIKdUrcUDs0d
96wLTnNqIlyy1VWhc8vMg9Z1IDvTq4TGA6Y8bnYVd4rg1r4f2gB0ctfCqovrj3TK
VchqmJ6/XtImH/kgZ5VWpRcXPd19xGiUScs4I86vGjEjgJ3yFrcd5x/+B7ZOSI/9
qXvQdmTFrcU7h3Ke1bzga0U0VWSPgMV47uNilWRtGNJhtBXIRdd8lc5B2LPoPk8g
S9FtWTJ2nyVF66YzthjznFikFJNPnIktvjxfXhSxlvx4YSVIgirC48DXRKgjyVb4
bOXi/lieDhXYlhByUldmG6hdrBQ5Og7ERu2EwL0h6F9i6EPnWIxJ44VNuvzAJ/s1
QNPhUgBYQmwtvZJgGG909H7MuHaN42L1LeG38XGlKeIxyIpg4YYJUSJ5SaW0oBXY
Yn01IVKfivXQgbHxqb/ZgRTiiCPT2jv0eFnNV0YVKJerPrc5ETEXUy7TrMXeCPcI
J+EUbrWgPuzOZrwhySEO2g18gGySliYDmqeK1pBN4bOBIJHkXXYF/xHw8CRY21/q
f/vtqr2hcCclUTj5Wh3AVbtE3sY2Qmv5lwy5Dbnyf8Vmgvz0yas3Vb36D7bapj4K
82saaUx2Ve5mmSLETX/ne3qtMIUMMV6zso6O9Uz6FfJ7Aznit00n+aykR2fUXmbp
aUW/cJ3qIY0Yu42RM6znX44XVh+ZtAx2a5GrdWhA8C9zF/TVTQPPYQwbhRmR/uok
/VXwZrwUDGmI2O/zfI84CwN7o3/8/xqdHwS452nsja47tV+TB/NCFD2u10+QhWio
O8OHIRmbfFUDau1uMmazZB3ra147JAhOSTaGOkVCdMKCAUv+bgfdFMcfMvkJ8vF9
JsrzLCzyWr2x82E68lvpZDLgPaD6SRvev9IUQGXQQsU1bPrnzKPzfWajamAwlaoX
JW4UUpzpFWfSTPfMqomVyU+2oLbXLDQg0sI0x+5m2aWS6goPdaVTHbz41IanBlo6
/1U0JaUbl6oRHqnXiG4hbLiDwhsYkzPTnnYp9Tg/qoF6RfRb+0NzCrPNbrBer6Z1
jv4lA/yBS3+4wMT1OcW1kFlWGM0MKFFbjtcCYtHQQHzObCveHnz969kW8rjr5Tts
LDYil4J297jAvlnnbLo9rnjN1MTnnHneiGat13VFtno97Vz//oPKBh8pfU9RkhFc
bG44ynAdhrybsqJ8jGd9hG3a0O7QDNsohWtFICDrIU7XQmkE97LfxS03oZP2aFW7
AdQgHEXXjc+QmsJ+YZtcJyJFNiHP6MFqPgtZKVwxQPJrbygi7ROdxq5KCOks10SR
KpPh+FZfM+VTWZOr7szvEPQlQgBsbRtqp9ECxibX/Skge5gbND3SPU85AHq79/b7
0d7FDlt+/U8Q6+trDoFKx7k5XIC0IQH6oEmn6/fdbdkaop7oJWPS1i22owF+1zQV
maO6qoqzMouEBqePGIBAou/htcmrHXUASea9uu1qpu7zylFcx35cnMl9UR+jsME8
Hw7c9brSOe1QxTBm5SZX2RiN0Cx8Q5394Dp4Sf9j5NFwEcDfx4AH+BeqVSaoOd0G
tP5cT/jDHiERJS//NxvE0GICiUkMUoCYhiky8yF+JY+5EESsc9wSYyzwyKkIxNQx
F1xAXx3/0Pu7KxlH5rlOpZipsefT3qZOENMb6MxlRXpX47Erzom8S5ZWW9mihz5v
/BszPLErMHmf5ZTAJd1aW3LP3ejEgMrwJp+PYx/TQiVtvfpSwWXilt/pCAfgjdsC
60pzyyumfJvJFfiefh6ckbks/8sW7GvbNV4Lxz0yZeyrXvbT3YXtROj5PU5XkcgT
rYW290GgtPanqZypCViUkPBxee3oR3518yv2qc08lkk4CdRJCNuNhAEtnQUUFsjl
tnabXRGH/eROrIwY9aSCCbwuYxLO7dJFczH0cNOcDhTh11u5XLAlPNgWXiYUAzdx
bSdRxt8yrJkJUSPGvr7HGh4X9lgup+fXVe+sgCbg+3xoOmT0DCsKk6wtuskUyiFG
ngIhKxvn1Kh9oG1SGO/URbUFAFFkJ8+jEZxAKMS17zefCD9wqBEUkmF274uLjEnv
EC4xxtqQRtowYuGg+PP4IKHbXT2qGwen46QY6jAIUjhVaJlp92rXLTF+R8W+YRz6
Jo7itxpeL9HZl7Kg9OwhmHCtWfK9+wIc2fXLlMOvJ5NGjn3bPCii+Qt8bub7UMOO
XPC5ndzRUjb+lytVmkmuShrBi8UuYt2lfAkFk/q8UaOYc0D0P14Ij3K0ZeUGngtv
jQEgysht+lBjBUu4EXrDsclj3TH3CednEwV8jk+7lBSTbsd6xdU7Wj2lESjNIyW+
JXBcoRIcIceQKugQI4tYfB1MC9eF0+x7RVaB/K5Lu6007W/sLn9ZseUECV1EnMIF
SeGX3wWTlJ1PYAvRIz08KVQW5wP4b3oI5oqyibezehwCM5uAaWMgKqWBzhUYp4aR
hHsh07lgRVU3zIkpNdBWoXH9qR07rFem/8KWQCXJiZJ+l1EELdEZme2SR1eOkYV2
tpzEkXwFZml9UfKE+nci0wO4ICzaZlAx+nMiOEerRdsuUhInPyNSuWcBEsAy3zDW
dErI6OcRghsraoDyIcG6RgW8bPJwuQRZzvoxw4YvmM+0HJtyKx+LWf+YDUvyi5ng
2SA5/N3udNa9WdTIf+7Sg+ZV8limwmPj5IYiyqAcY7L6JaAIEGhB3rgOSkMhdWwK
CaqZEG1pSCRxz/3m+IhcDIEOULUorrWAOmeLVdlW/I5XJhg8/GvL5dfbWCjR+2Rv
TPWOyRJFS4yOW6dYr1hFPFmQI6GOmWHebo5TQPj/7XBEUsqqvvPAVn59v2ZydUK2
cqDJ77qPaqIqkKfyqVqHsSZiIPHKYmBzYV/1dJGM75Lo5EzQ4RZFVOdNhNAjvlyd
0jHxUsYtEVHFa84zOpJcvQF+XI2XVGlmdm4bgDQekycpIq5zVstkfXRk4q/JuNLA
3wAH+TsT3qt/Ay6141/+rNs1CVx5sUlL7T4yeSz6pY2U0qSlME3O0I/PXWIDEf5R
hWn9eDTsILtAbI0URlDpM0GrZ3pC9qVf3PK9Cv/pZjihKRoF6GwMPItsW6f/OEh8
y2OavpM356SKlKbBpFGIiEWmNVVvXyZ3jHzHgWCEdzjFKMxqv6EAmhciIdYLVkw3
p6Ok/dQYTOeFQHI/cKbkyKeWS7TwsHNovQs1ETnyxeXcvV4EbpdPR0wH6P58hDfM
oUQaoA7yVL4LoO7HgcetHd8FBqhOAyFDA2IBFUN9sOA7n7TB74FQP9iYH2dIxCRt
Rv/9uqm5Rvn9gIx/ZhRekq3BYVh1KdREuJjbIa5X8m7Psx++3/XNf+efwfOrLTZJ
dXx7O4Np3+WxyZzuhu8BnEjJ8CdA7x4jGZbBMfvi+PafhSKrnvoixh4QKkzFl/hb
c+NkAUMWOwdPbVU4jVECbDBuoMhpP+vrEuZxkXFaIjNG9d/JF1CjpZlbE1OAMijE
s3Yhh2OB4L/hkoNyRLC//AO3DPowpdMiA2HGmrF9SyIWgbi3qpsNCm8UKUafjYAU
zV9Oip4rKMfc0y0NaC1T3BCOdJ+M3+HDvEf2VLOX0/O+G6UzhSxNmAuD2k2VbMPt
fx0qv9vFqBm2SELpYGJiL1vE1B0jh4JZwTMTyyyAGyTLR4P+brTaUpUCCBqRwAWC
x8D9sxv9/3OW6vivg/Tde7gDeNyGfupRaAoZPUH4zT1xjGt68T6KpmpN2CbC2j+u
hmDsCt7plNj3ZR1gC141YW1nh5w6GQE1cclW/n2hQxJOQjQV1JAMATGzTNKBEoAA
B+DaRtXFQDugndQEokgxD/0KieZXkhY6khPlM4nw2z92RQqbkQGm3ST+ho/ZpzlR
XrD+RviEyZ6kXFQoeLqG3ZpT5fHvnThdEhH+Bu92InxbueAYtWM1ZETJLtDB/vzS
DuhoW05znSF/0iEO47mxWp2dBdlqz3HWp47mxsMNiAnUdo7UGHN3hjixFVoM26Bn
pCniGbgoh7MDlt+9x4hPPKoJXMBCt2OCYLrfnCOfHscux0Bb5l7UVEYnka4/EkM8
yX1F8E7PTlvXZxvQGKsGAwvLBcArmRXbBs0hb50Qdzew8QcA4zS9/6SjSlm3FZ7W
RbKa71W5udcWWHjkTYFXifYi/j/pfgqUp6OzbmUZqjqkwiy4Hc/MN6OiHdtO1s50
UZKtCQrbxJiu/VTAWGdNUT1CqG9Mu/MltMbgqruy72GiEwGTGehsEzuiK2aV26yi
qStk2dZp9PEYoIQtrg0i3RdJHAMqNADmDvxch3mjz8pz1zYOSS7FLX1IJ6OP3mfM
ey5bkGNKPpcSIr6rC0VaVqkUb337cX/FU5nbKpilK0jSLAanzM7b3kSD46lmc3ap
ekwmzo2Afpg4zyLVvGeOkJxSNFR5LfZ9ojxWajct2oqP4FIFwikm5Ocsz9KpGF2s
A2pDfhOFufEuRHWBe2l1wujdSgrwMaBUBXyCOewQVDxLGDQvpi4UhXD56paOgul3
2nHzyDvEj8Kgm4SGDhXgk/H27q6ba5p2e13tP9bhGy0GeekRkj/wfdBXeFQEaTET
KQ8Q5XCRaBfs+FwvttbpY3v3ohKyyw0043XXUanbONP6H5aKf8rYLsVN493X4aRe
P6bybKHX3oW8y86CR3bcushVLIupVr5xIDlrsaqvmMYK/a9cjKmHLz2OseyoqbqC
GAx2cRA2kSM/3xwDkJylEiI2JSDi0HzHQTJio4xUXlAxKn/qkkpg5XFMyK2qXArN
6vOomTfUiOg8dDCWqY8hZZF5Uz1+IPJt5URohC57nesRD6xcChTzrIiSTBPJwDBe
6MW0Q9LdF9yd34sSRM/RNSFtI/1m6w8l47Yc45UP+/Dbheg11ZgxP42jTDNUt/ur
RrBaKoA2zFWgSW+95Sj+G9eqhLB5VL1FbRb5RtvnMyN9K5D+ycFWNbfNuF7qsWD8
ka3lqm/Ljha+mOBObekdF/Vi5zISflgzYH1hBY1xgxDbNowoCzXpgdcEIgqfsE/V
/QXiCrwNNMwXgh3hmRkhcwXcJxCGNAIY5l+I7QUE0xz+Px2kr47Vjt3mW/K/rCkV
2bx7+cG6uavJVLO076JMedf4sc8w4SrlowUO1V0jwteh3VNop42m8wspZ+DvPYBn
c/qk8z2fpxXoYCBADvSu8BUxQijojKpzQ+8LGSVexzdCBsGS+Sqdantcqf7qWCtm
6wJ2N/NybSo0+GAViguWlWMQlKDs3nyN2aYVY1s0RoTOneAwlBJpFBc+RsuMB4JG
vhMvuhMffW33OFyfaIPcQ0UJAxlrhqmcOiXxgStJ5t/lpuU2VKhfLU5HIMkscfaT
ElDZttsc58xfuuOdWYLRvsLlH+j+1kPDPwfLGiJMvorPks0/T4ElbTn623E5+04/
xY24Ncdpu0oOvzouOjtjizF6pPAcDLI4HodhMRCcxGEqu2FdGTbskIVz2+zunAEL
0ID2ou8k0YMn/3776gLqyPzz8Z3WkmmBWBaCPojmYF/oJr2Mw6STewo04fcfig/L
afkfSGD1ArpD9qBQkG0fEPN1pKPUkgcbCk4Ab+Ti64XOK8/ERatC7e/FroSobOn9
+XFPys73rS66TQsEB9TvxzcP/ueSLIRgsdR0LOqLFuZP/oPCOf02edAASfCgaqXL
Vbl//bd0gmfpTjU/SyFqJ14WZ2xcR/fM18Fb5wlg6gmZj6bOqJdpduSx/bepo77l
IdAmdcEx4rEwTd/WtJyrs4Pxlm0p2Kk2OubbOF5xsSTA/Vm3mf7f1oHPwWlpNjSV
SKzQxrE4pxUwBJMdzw80GFLpt7J6uxBznAlQS1rTjb/H8ETfL6JrxxSMr8JVra+K
AggfaVKuRlTywBYT0j3Qpod3TAcs8H2vlF5ldVcRZ+Sks9mZeZGgVOsfuZaFq/Z8
ZCyaF9csbBi4Y3krmAa8yHqYq/CmpRqT6/V6Ioi9ZsnQUbpVfB3RKuYpS6xlMdlR
OdGP0VMVQAoOHe34X43Yiuj8F/Gm/mVIWwXKCMgILEKdQdld4s6q31PBPF4XI/7O
F+XxBHU3YdPXwsxXQBZXaoYCT49oIpsbq3dZkI34+ZXuwsVQy5QORxQ1wvE6Uhaq
nS1qcr4zgRt/20R15DCdb5qTRG3pBUHecfPGDfWDZC0PMh81rGso5pWVZHlWB51l
6GGInIa89EdPKqQw4Um7+CTAPyIu8eKhNtoyz7b7tZ8OdUNaUaVYtADSjy4GzaXm
zoyhhJefwm/us/P87GQ1C+utK3gUL34sMnRXSFMgPt388AEBL13ET7aTugafToI5
E1RcIP+xTgGmf61N2emWjbai+gtluQk1oVcwls6OQ2lquAEJr/63J1/4XSJt7MQG
e8UyqSCapWpkAsZuFOM3+4zplDpdB04R6MyuN4MrcZMNAz8ImqxTQ32pQ/D76lpy
g5fWe0iGkbS2vqYKeu7uFrBMNFpiW4kA4Dbn4Cq0BY4Bf4H85c0/TvklQS23wLBg
zhBgWa8O4DpSZSr8oB82BL+mxTlEjBGGQoQCrHPOpR5dwtQK5qinPjsI22VQoqUz
ghs2reXkXc8reruIOdYA0xAeReKlb9xyKRx/W3jqXgvifqPJcIx8WRxzIA0vWv6g
HFpqN0mdkfVMrouya6WItj7Qs7ctBNJEa1Quehostf1NN2eQpJ0JUf8M/0YJQaHr
DyvnjJR4VkmV9GPwUvBWW6wdMG0ajB1JR//0dMLRf7Ds1pkLjSDy6G0OL5EbpvH1
4sPrRwb1nADMnRyDn/bW28Qc2YFlsUdftnRfrKxTt4so9qjLaX9ZDjN3eZw12Wlp
d2brVWlPRU9ssWlAwy05HZba2pT9KL0NErvWDWt6J5ampCHSGuy+x2wpfuguqDzk
QPxuy4xEOQLvTcyZHoLXJkjrd3EM+jE9a099AuNcBTgQuhFPvpMMLzkAcudF3mnU
zqJtHQaXqqIe+39uSD4nmLx/A2tgPu2/bjkcb+P2gJ5o4/fbr8pCxtCEPglmJq8S
2NC01NYbe7euuxsRyLqA4xKnJLxu70O5tNGr9TLqKqfeZ7k1CMb7+cyK1Y0kPONF
vV0k64oHl5g1+ATMSsaOLN6JGSzKkInHypifKwxHeBA9iB8wk6A+9R7fj4ijC7XA
1OhFv0ZDSZAFAyMXAl7eKCedD77Gzlog9DGvaBPd51uoSEJk7C7J9ZFOt1mC8unj
AUGtf2WlGv7DxYJtXsPAbxPKc1i+idUC0swcGca62IA/qshp8XXDesMB8GwFXhYH
mSdoJsOi4o4Et+kCX+W8QujMjf4lHKU9lpNLJeslsvTd+kNEyGYiePkYk9sYK/ac
c19tW6DXNjwSFQs7xV1mHr59k2s4Rb3Pz4aimrjHUf2dZvM7qu2sdyiW0I6NDZa2
boj4tnhU41TTh8p2ZX0bCoGJ7mjUehyF/madFiVuKi1iLtQbPDdMEL9twscDd2dH
/cGxdTrWIpfKm9p6EsKyPgAIAFAXpCh4INJO/Z5Cn557WHH+OX0kVIE93+Flb9in
rqOON/hgnk9al7hfGIGJ/iaLMN1H/sGxN8y0tC6jFZpKhqvV4HjLNjHx/kBtkKaM
OV3EOnIs1hOQNKTeTrkUb2hf0PEQq0a+R6yZJWHbsTTwiD9iPZyVhb1D/NI7a8MW
9COIRHkDIA8SimE3ppjuF4iI/a5B2Rx/aZG5UDCtlFaVW+iHZlwFmCnpX5vb/344
hdSK/2xR0HmquWozsAo+re7rIdaVrXTPsckRY615wtRj4xHguRiznMlA2fMo9DZg
bykGhbftRNPiLG3dCdOsrEhOgDMPn9ix4Ap51OyqyKveDtNvg77LNPu740LrL3Ur
SB1cjBGnjm1vJ+nvmkni4wsIFCP++fIBy+IcfM8PLr7evug1C5FOLtafaTQTCKtr
u+Gwnaj+sGAGHx5CIFbr+f2L1ZSpLrFtBF00gCv7nrzKfsEa8A0gC+H2jI1W5pxo
UPTXwQD7MK8ArzuZ+ubmfCvGK0xdmc4J1PvCsMK+ohMb+It59Gy5cwlf8GeNgpsz
hdkXy/1Mf+X6VC0jyx8R4HCSax4AyrPcxyPmAACX6q/JPCfb49fOa6VPzOn0+AAl
eo03KmqmVc8/korbVZ2gTprduFQblnFHWGFo6mGY6GK6bDy7ikHxSAwPYKKOZ8tF
fFClH7KjD2J0vtmG+w2LeSVyKv4GH6YLzjvNDppkqG3aUMTGyMU/KWSVqHd2oze6
Cvkul9Tgi7jljoraCIzEorVvAd+9r7fCn9mZ0/9EQsy6iFH4E5ZjweIDjjVjWKyH
eEE9yDUbj49VdWFN9vxWQYPrMey8AtHThgmbFzm4iIEmIfeqjdAKdie0X6CEnKQJ
hde/yridYfTbNHPtv9YD4mQx6w59A90XinFjhkLHZhsrO2VYbu95MuT0yeJgJxUW
Alld7evbXWeIYHVETXQinjvgiUvP2dUa/PKfAdI1hrpEjN5epG6WIgAl3LrwSLI+
UuLE49LBEFgtumxxCUx1PTvAnWL86jtTr/Hdjq9PtC5yR7u7E1KYVCMCYa0w00a+
zWgkaoRiSR6vZ6y+Km06bGLMuzCjmrQumfERbCKViySUl6f7XS3YyQpaoXVgnd8l
yREMOe715sz/jYG67/crIF4Ezsx/PhByjRBg2RE/VEHTv2CHfK9MOMzVWke2jWW3
TC7bE7U27GcQkZYT9jBmqgPbr3MydNbPhj2KCRobWgKxzS112IKBq0Gf6S9QYbIa
AZch+P9h0woV0iIZZ/ug7osmybhtAjU5WYYOfVhqXCsVa+2BcRHz7Ly/OWbBpm3W
N4BPGsmHse41P3IE/uBwwzD/SBdmpZTYGcu6LuZjR4avsON73dagvQj42WrK54vg
CJsbwpymcmCTgLIlK7S1DmcvcXhMWbVKdvqgCWaw1IoWVmZ6xIS+M74LbuqGTmWY
eclcPL58JljKkr4en6us4TnvZGW52gA489nuIYvhXjVWHj2p86JD6HN4zJ/2y0t6
UZNMN1dO+QtKh6bk1TZuzf+iS91PwMMtoqyg4Y1t7M+gUxcP3T5dsgz5X1XxYOvx
raJGG34dyoVk3rKRdUshdS677vf9HR4TXoGxMa9sqpRYhHa233tAVtRLXIr8ADY/
IMqOqJTJmpABQcVfVetUzZXlNWF/ps6O2570fRIOmnTs6MABMDQnWjh7bDvF4iH2
1FwehemuiZ0OhQDfQHD27BCxH9mAgCgj7dqWCBYR/DzWTvWp5PwpZ9wtFG/6IUV2
iKUPzpk5+FWhr/Wv1i82MTKmT6Iz964ZWk4GDm/sjP2NcZGHi9Ga0lBY2pbuTJfv
IE927An+ExAy3yT4p7dZQzijoVUnNqMJLAKoP0gNRVXeIOiMYTOZx0MCTbXdYFOr
dxypGuxK/iMKf7nezwcGv0QUGTXNhrHBiVVy4YNCWP4tPHpOmINVCvPGd9d3VlCM
/7pOui9Yj3BQ23Ga1Bj0hjJQuNn76oYjzcoMY3xYmylymg/LikATTCAStrXWWBzR
+1/qMVjYyuaCZsflD9j/N+wRYN70AFjqh65hhsMYerrKxOwv/3VOCliVMs0sAz51
i5crURkSyWwa9Ovy45MS6ZAIf2/qBrx+1/66ehA/sG+EXsxylwKRlyyIWDb8N0Sf
YB/Q5QktNEhFC5XUm4r/uOcZBQ/OmeNg+uohZe5iEJP4vRZsVUZp7o9gwFqyIBYL
F5apFE63o0AuTEwMuk6JDLnLcfELshQuH/FTaF74Xh3BuSfblRDQCg59kv3C8Z5+
sFZR5ZDXaO8xm2emSQi6smu67F5jNn+zu2+bqDPbn600JWWkQ5uREEO8vUpK4vTf
Zdabx70p/O68EN5b42MQ1dZgMimqqM2fOfuyo2VXWZtad2o9a1BSzYuPe1xMD9Cc
l5z2udGrlgcjZIuI+uI0EqOwDYlC7dqNkq1yH+PXo5Lt6tyLGxHLzw3tidllUGf7
cCAsn129tOePyIWQBuFdPLh+2+90cWcd99otM41G4Jo2hjpVTm3cdZQEGSSDaU5N
gz0i29mNWDCb7KLoW6JbYFtU1ksY3rsLXWH2MRbGSdGAtied+/AfG9LlgiLJYnZl
bVsdKbWj++FX6XYhoXiitUeBFt6CQpR5A1QkhDN6W/FFx3nK7mAcFn15oFsgkWKs
Tv1A1J83YcOpHidFJMkuJHCvx2O/62TfOp+eZmNsxxSQTikuaKHbWQFU38WpGqsJ
vMhD0ejPwsd9pb1ftp4na4E0zQuPxYgRnD5IDwRzddTWCMnX82cnmf8gFFTyo7bc
ErtbSaIybf3ghoaEh89K1Okke5E5+E9gQzUf5f1k84UAhzqXi5h+M6UMNLAYzo72
acg4GrIchuLq1KWM0OaKoXcunn8l0Kkfq4PModcBJ8AGs/ePnPjdKrMLmXaOHxWG
mn53WYEs6Nu76DJs9MhLV6Zb22AngZOCbQe4YlhqZkTmwm0s7dmXpI/zLOiZYnyc
2hNfzHM/SjRLjRjHDBoJIkK9s0QYFZoq6UwyJPjiEb85ayJKO3rVlO+O62xyxaeF
B+xofHqfIABSRu9aQxp8JF4fohMj+6Vp2pj6xtVlWawySveM5BN2SRNNj3ZZPEVL
0FszFiEOx8eUcbwptpdIQyy/0WhHENLd1QUFi+f186t5wkj0vn1sAUll9gpo+t7j
CR4SYLnS9ICDLk5CjCa4ntnRkMhJXOrhIqamd2G4cV3AosePcakzpQHMopi69Lj9
wcTrrL+pGoSV/nXr68P5tT+5otbn2azxW9G6fHrIegDfJsAlfeCp3W0Sl6MWoPcj
Xi6GExsmxOpn6B8v69k+KjV0ST/tYIfIEbBcdfPJ4pfJjySUkd5HVBL0ZHMPz6sf
OpgMpniVKRxISYx+d2uHFzvqOKCVZb4nRMbJdSRriq4H63te4H5YDgx/pz351sI0
wNlhw/lxYwEbYA7BKXz5EsRYWMY3z4EBIVlkUYgA0qUUqqosk8CTZqRZLGnWzQs8
cTdNt77yBrNW+blyZ3KOhPRs+J++UENfIHLk3dpCrcC1aMbGHqw/xPsiyufOK7TS
6WZLufRyWGBPytv/qYD2qck9onpYjNaTei/MSWoVj1Eh4haDI+hy8H5nCIoBj1M8
SRueWnVbrT1A2l3u29AE4fnBAcL4wJmfPP4119geSEWHyOxN0P2V17Bk/MUfWK13
REyYo22dtxFe0UiEp4a1+0Vx9sQXuxM0RGYHWTleU0CQo3bWXk3jBYdcbHv+WeCY
b3YM7fh36u6WPQmZ4soay3O4S7GF8nr1eV1zKl+1nhYpDeggz87fVZbitPljm9tr
lnNdmyHvzqz9U+0dgnojt1fZc+bFFLYnMcTIgxlYXiu1OafukxecGQ6+5byHr7ec
czCWCeGk071K948+df1SkiKNdiJrBuovTYcJqEtviKpiC/iI102KSYbI83Y5hqjg
sFnsRJ0iSQ5/oJyEXu3UcemQjXG3vxEPrqVziQ4D8IpicJIez7f6rSNra+KU104m
X/ZYhkEpVDpIoLdfjHco/fcz3s+4vKHjwFSZQCk+LEMgELa5rPLVTPdOU9/ZP1Q9
yd2qGkV+eVP1PHzaEFFFFDSDpE4Pe58bmthogRXD4DPRW0TEQj7z4pehSVWEnxCN
IWAaQ0YLAl8qUACK9Na+mjQjmvLP8aykjyuBDDRymhJdIIAnz4gb7zdK7IJJmUCp
QnVUTgHBaRBKX4ErO9aoHBGCwCZ5qTcZyAQaz5uRs538e+7w3j4h6PFdcKJxDPWu
Su++HVDq/p8tBZX8czmmfqdSmugEn992vDWKwrEickhtULcvg3l7ZTG394SgYnHz
1716tM63mhbWXkKLRxgQ3vYNTUpCP74ZrP8m1DRlCOt2WtrZQCiThAOfazrRG+M8
qdry3OPybeLGx3D5oQgjpsHvMS1pzDus+XFLkPEbJv9AhIExjuLm1sdbgb6A5h3h
B7HQayrmfC3AkMFuPzw1sEegs7JZiYEsXfBlyqqk5l8HCkjlzTBNcvV+fGg+3rcR
0fZbWT/F/ex2oDl43wxEabHd0+FZbpJ2GYBlhsfepB3S8J5sJtVppdpP5A/bu1MV
0a8rD96wz1HvVTK49dBNXMGM/IjQ3RgafLYNeCS9GS1s4jOEfq3XLx0JgMBMM+co
3yhPmCMPgR8Q1Ijn1cVvK+1FP0E78o7OCq/L7UMO1Gsd4WdWbIQ6pFhC80X+hDI9
cb3cYHvVCWIGG273FqsHFrAkASaaosgA4ugD2d/UlsmPx/n2QrboIfn0oLNJm4Cv
KQpFlAdEQ5NcRWVwrCLQjMIuSBi35fWw0eAXtRO+4f7FIXmdQ3Q8AAz9k7WO/+An
m6tz+NVAvq71K1O6xJI8CzLB45gNg9+vHWGmFmQLxWwVK7fxdnjHYUY7GwbCa/5/
ZEkEmSkQ9HgwqAFmSuy2a3xHciESLQLr+34bPKlGeXR8wGHn/JorGoQurERVJ7t/
/yHlTC/LzrZKe08n/tWLs2bBq9XZTFsRE0P3ubWHSbHEI6hgiYl55HpHH20l7Poj
2NCcyR1meMXEa16KFRIKnbmvEOEQP7rO9IwmHJbFy7HLweCV/1MMl6PWcH+27wdo
T9SzcEvquKcm9mh+QVCGqX2PzMEBi/QBkV8Z9EbCTXdAF37s1GWw9wvy8xbHyLBP
rAbUxEK53pmcyhdxBlsDerQ/6hDn9uqtuzaV5D7eewIdkyCSkEXB+Yp0LYKcXhxu
KmwnrN5SdaPsn+uqJO2SKSoA2Jy+xWDfxWpzLmdtW3e7ZvWuB1zCCpFqCX7g7BSA
axZWMLzZ/c96yBsz+RF5mmbvzNVOzE3eUfs+ZOdG+dsbWtHwNKQKEhmJVElLoQeP
lk7vbYOunRATUPdTjlcvhjynPiQChV7zvjyd+41c4wj+5gfcl6ZNUAtzyxdeQYEI
IgD36reZCJ9hhNF9KCKw3urLxx6gID6HcJVQc8awFNEtlOpTtQdZDeAooe5yUKG3
tF/6vBvgvZxaiyBHcPdNtSI6h8WD+yDpY0PTw9cWC8xiPQmvs7MhscJpY+l3b7Yo
2NMiYFyXWaK+a6SK5d7c6dYZqgP4+Ybr8GqmClinox9WySs/OOcjJ7UE5qhHG1ec
q7bZ/22TyrIRt6ING5NEaqF8iGxiBDkaw0T/ZbqnJTs7I1hp6djLWBA21zENib23
ox3gyvqeKi6A0thZVSctEUkqKQxngbxxBWTlM8Fb4/5oWOMG6QACsJui2wSmpVPo
NL5+o/4KRcbnurZnjdU+26a06YyzK6RmahLD1z7MF+5LmZFR4LfPz8OC7m+ctw4l
Ug0FaBFWAsFS8vaEDltPGROY5VefUpL3vtaTx4+ZRk92/2G0Ymyp5nONT+KsGHoN
m+PEnOo4HBpNPH6BVBfptt7G8+45hxT5uFa5amHXC+Y411hLRF0TJlA1T6WcW3ZT
nn7cn4ME6ymOVvsa7t4+k1dcMGTjH+IxhAw4BXnD8Cop8wWhQm1Ai3Xvvn3MadzT
6sCnkBSwDkr63m+QrsLGe41gdPKrbi++nFgg+pXXwfYAY8acXduR3v//xmrgDCTS
3wIsi4VhGSE5FZprupVdNujV0toSrKlLAdOIOdMeAvQYRxdLd/EiJsonsHcXL56T
FRk/+2jiZX/9xDrv0ydqsCGi3JRYEuSyYG360vHyH6l1IYg7meVw6Nwuj5m5hWVV
IS6vFhQs85AH7NANC3doZfWL1QesPKMDGduiu4LXI9caSJu/jDZqFW3os3QIbKOn
ffCBwJmQSC+U6rgb2vG76xhKJkS6eYK+rX4awhXFawlDBsuIIk7psdJq6AlgwlI9
zQYeiZBj/796HY3svZxAGIJovsCnRGSE6XQIihoUIRJco6s3L9UPVrQv7l82QWT6
z39Qy+Ob0DXDAmKGXWF01kbrMrBl3kqCl8tro2c7mlR0tlgXXdZ6tYJgzl4Lp5pu
0HSBhU8mLOGLrAGYDFgM01gcrSD17xbEa1s+1hB0t87uRZALg79FpopIgoC3lBRe
YVnsDSW+oqk2E0bks79Y+pw1EqRB6wlicVtLC+nMvsBpm1RxrUUk/6SQVA3cvbDp
aXHF0oKkvbjPcYg8SUqFmlkZR+01UUn+ATBiDY0Tc2qxKjnYUxLsbcXVRR/zr96C
VGUck+L0hpZLAeAM+8GrxrA2H5EIZewcjMr8BB7HOhNDb1LsTR6GNQ88aoiC5FAO
8DByxN0bBiJQxwYetouzZu5OOTVLmaz4I4mQGSycil8iM0Z+w8FIL6g66yhPEFbD
C0hqjdgt2pmMVIVHx46/okNfTccijr1wHCdLNa4Th+oP2/F1jKgEyXomHW0kewsZ
P6KuhtgoesdlIIiBKKWg9clGiqYeaz4xzNqWo8uBN4Dwgcg5pCNSS25J+tIjqh5f
Swvmslcjuhlb1E4YX1+aCyy6NNa8WwbNZi75quxCMVCCFO2u8ZPNNM6VYXntUCPQ
Y6E1Szgs1igw9k6QxJADYln9F5W/7qVr1MFw5yZao6V4/H6M1CgGv7+l0Vhybe71
sLp59Etl6l6GD+Z0iwH6Z+e8J1+IOG3iHX+znd+eGYhFnmAqSBcEGfi8MQakf2aU
jH9/SKVpfCHVGPGsoZcMymjpC+qZWZw0API9yCzDHR9Rr4ukuksDtQ2hAvRfbXnT
8Qk5xlLw8bM3lojS97hhs0KIcnseTpSrXGWhSQTebGKKJA0om5kyqvTzf1Pp1r7q
jkSWpKHrwNtnrbGbohykPuDNbigv35L+kbnpKXA+vKNHc8wVrdAq45XkU4mKG8IG
zSA2r+VB189JUKlWFh/2Py/8s+Qk+CttPr9uoZlUYJGrTLkR25+mbBcBkrq5Jvta
xFIXwefSjJSZdae0wmxEfbnWkRxoNKMMDIozYJQ+GU8n92JHR842oLB99rxrOyti
L412HhDdkrUB6Zg8FmgxgIirp/6nynL1GdH9H7qHYHV2KTcs/8O+AQ259G/VGsod
fXoJDPlDDkM/vwERlypc3nZTBexBJlxvBbfC5dtP4H1BjKC1bdQ027PSqTu5lgsc
CTZY+LZbTDsw9wUJlrw0TtfWfv2E2Z7/K/AgJhQvMoiajLt122V6NKFmV4vjqM+6
NCAJA2USvhPc+L+GqY4/3Y1dX7Bw708F9AanbEdU/xKVkH7RSow8KZ37vpGTobYx
s7eMjzCRlIgQKtTvs3tpunSVwB5Km2EhWnZbxdy9yoiehGQJvAKWDBB6j5Fw117T
JMaGgdqdvp1OAdWbZGjn5TKTek7D+hoB+M3tjY1tv7QAZopk3gp8UGlrU0SdCLJ6
JuyR4Eo5J5oavmHpSmM2KwCW9kuREdm3FVKW1LIFwUOt0pozM8BOwtYW5JGZhrfG
rOP+yVuv8wDZlQbX1V8m2Kn2f4ySqtbXKUPWkGGEAoi6tqtWIN6GoUmbWWlZcvb/
jvmWTScMGQ6b9b7Q+bCH5sONbo/Wo8htYas0KacCrj9ZmXSPaJ2RlhM7rOg0sJPu
4ohJ+rW6THf8IkR9ZIhGjprcRUimSgKnBJeSuELJYnXVpkKARnXN8umK77m/tar9
L6BxcofvgA0KYkWUMR8R16Js6N+ksjUY9JHMIaAxjanZUrR67BCjsT9DG+UmZOPB
giKRNBKl5GywzurE+7pcDT9aNhTMaUJpOYiUS4aVxLGpBHdV3IURLiJiNdOms1sf
IJm9Ew46QR2v7K8bfGQGWOTzwHTJ5wUlxfizEmA0V/abmDMwk1sqmihtw934OYWL
1rjEplvSfk3QxSNIT6b068pDK5orKY3l6K38/tZ/2QWWhO9n7pYMxELqt1LcEXK9
sPGnvcqUrV3dTiKQ1pTC+0xNDKWtntCcUAc9CtHcRilvXlEQsSxKVj23t6Hcodft
wYUbfwTgaxb9OBVVPufoUUOx3aw08p5oxSd2/TwKy5ARZAgQMseAHIYnHqHl0otk
z713+dJ0cKJjP1Vn2n+hPshkbmngWoqByvMModdfM8zaSwASSwr8WZ1538zBwUhi
xEY6/nXD4pqJmhka0FYbIGgfVeIH5JU6Q3hAhsLJA2wJpE8OARERcZ5aGx3CSECB
Kz4KxlRWSlemigSq9GI1qA5eTU2u8Gbrb7/4VKb/ej9umUDtr8Gno6BhnrTHwe3n
mpZAkCV4ILt7HDde0jOLhBJzDmkH1ipVD/Eh4vWv8JlAbNsmV63lqaPRxykMqT5K
msp+bcxlJoGqdq/n3IE/ewsZEBPZg82PcibltRqLt9rTzY3jNXGgzmZz1E/XLm4H
tyx/hT+MQ9izbAnxGzDh2jebxLAzzEwRRjuagCbnY7oBs+ix3RNwzC40FJ+2JzbP
zPdHkbg8EjtO/Wom3d+RCertq+O1r222R0QcnkDhT+3TuJDj4U2KAvaCzyODoEX+
xa4jV6X6kyySkS5TclSItTEFjLRfruFYspGV9SIUTQAx9Yu93jmlJ0LQVopUY/Wu
zi9TpUCGxfgae+bEeUa7Na7U6xSlri3LWd+ikw/Cx+dCvYMBP/MwmRPOrRUczHrv
g99j1TOp5MROT/CThGmhWJeay++tW9fdqpew2nGB2c5WrJaSfPsHJOuvxEF3zJQl
OqsU9aMNNPCTmboTDdczlfszCXlYry2n+D4qzwCiAqL4JWF4clSFgZ/p7hpFm+lX
pzF/JfG620NuJI6PrFWwmeZcHGDhfIhFbsFeHiBCLFrjB695nLKpSoy07n3aO7w/
LYP4JyP0W8Ke72C0uoG1gebeK14vJkHTqODtZPIY4Mde8dIvBZMXvUFf+FpWF3Ur
5Mpp05mlz9jGX2zCEMNSrDenQ6YOufrnkFd5vvbbMgiwEfcW2qcF3Fdtd0JOTp5l
EcpXsqo/7fCCClIt37FqUoT5LxRhKOa9jhuTHhP3AYvlZ0bNt68sH6FVJ3kNHqHt
m0luNbhOnhmUh48i/PEJYWi7rwDmmfeFQLZdNqz973XN04mJhakyOoOs6IKsINwJ
EzRTu3qDIsez6PD8PMdX52oQmV6AHJptjSF/w30WHPwJjrSzNL/AFFoLoN9OsuEH
GCT+ADl0Znrid2cyjrwE7HcQ+e+SNMSbQ0QGsg/yjKRbmr60Vc1m1H+5qdgg2TMc
S1m88pit/zZnTRp7BP19iw3jmRR/7xMo/+gtVYVx6dTqSMuGV35SftWZF89cmVm/
4ng7Ctw0uJ7VjBoYI0pb6e7NYSEGbBmGlwo3SBUIfU0HdJVhc38wQOfJGetV1K30
u+DQ25730gmTd3Yd2d2qNFiFUzWwc60x0jOFkHsYFOQJ+zLPl1Ly/tW2vajkyWPe
4vcIDw8Wl+J6Q7+gDnRVc0Xd6DYQyjMbBecliJjd4BMwDWwobBYbVY6Q+nLn7dlM
gweFl0ycTxQcA9m+gVB1/rs7MEFz4ZgIdCY9aIU2YCWX1f3Z15drGQarnxx/LeFc
mxGXs1Irl7vGyj9z+5ioxnr9hKAXGQYXg1iduQrdu8+szyiINlW8oRBTLhP9IqFj
AoZepDs17fL8C6Mk+Zy4LOUN53yBII3AhoG/4vJwvkqE2yutzOYKvDWLC0Miw6G7
i+5zzGYDrgaUBD5go1K2urWrAOj9TLsp5p69DLAuU/iJ8Mf4ATQ9FRXOB1JINTE8
kjzsEGU4r4s7VHotvv+WnoldUjLG5OSXIn0RQvnsKf+cSDF5SRWhljD+CKUybLkT
NQXTW7ORsR0zul/GN1R8myNcGqMBriS+ySB6Op8s/U66tt7FZphbz0xkVl1Fsg+n
BNxy33MLuSyKyYigMnmbsE+OKDUeHwJE6dtzGRDa/eAzT28UoPGSAxyqcycJhRvX
gaBoz4odzqegZr5cgoYpnqjvaDVUxfx3sXFMBfyg32lVLZQc/9BBJF8S2nSnoGwi
LxBMqKxra+xMNq8IY/qf1urZDW26gSH6etYcbwiG8GX80z2BYa3gW2KxLKS11RSo
YR1UsonvsG8D2WqWEVSomJ3CUPMWzHp8IUeBR2QJc4GQwvW0VrPlehKezWTU1FRz
M/45a5wUVuiNEkqidBLevOTlQukBYUtH6xiS48jf+h/aWCAFiK+tEu2PKxBx8AVw
lXEXmCRzrGXnHjlKavTUpEvMZVsWIEJEBPgzlzP6+3yZDwj0QSAaMAEh+6QNPUn2
L4GlLCbmsU/hZLs5lXkFFOqVn3Lp/czCcyjhHkPfr9F77nkEolb4FuufN8p2VLPd
2mxZnjVDQfQAz2Ify5/TbXDLrv7OVdAiGpnn52kuGgx0LwwoyTrSjngGSfQna9Y3
n+jC75G1LqiQkcoBOx9KA8wPGRmxTI5jXTrJpcuH8bfdg/VVOPBk/TdGpXj2RlEb
s4+SjeXzToLTA/CFLM24tevf7rbDHTpRAno/g0GEc4N4RDzXbPHnPsw9G5r18ZU/
jpC8ondKle8dhczo/kGsyT0IizgAWwAv17DOG6/79q9R1ChL1yHr+9y4jaogNwM2
GAZSfipsBwpLGusDHDrVS/6XFASxAMwbeqjPqCXt/48IrxeSzy+JomT5KgmzSt4L
SOQ+ea25rHJo1/KWlkyDeV8UXkpyTf3DE0lgvJePBUYw/A19V0meVlajokldPn2z
75OzUtClvfstckAp7g/AJamMC5LUUV3Q+UqZnqfPHnyAwM5ZlOpXH9QAelnMhW0G
fr43njCoxpgctF0VpkBoxXT/BzyPis9Pwuuc/bzpFaKDiicryTybQXoFAUxNbX/L
Rrkmtvun9wD+TBmT/5pymwcPFaWbOOCjohQsR1dlCl5uHT9p8+Us7R1yq3U0fYbm
FeZ2hshaIzC/PGVp5b3qst8TCFaQOxOqb03KSnfQQ+HWS10mLEfmCyVvtwoW03gV
nQT1fMC/GyCaCu/E9mVPFi3tXbSLtrwhjYbHTmVynOVfeX8L1mwg/X0xr8tIsoQ7
6GPgqf/dNjvfmSiUn7I5ja22dvOByQaYFlI0FKCXxJkDDuJwb2KFzjHEXX83CLLQ
xDJtoo5vikRxVqCfqTcrx0MsL3Lg2KoDtISgXkYkFM0OkKVfsY1FEHc0WGGsQgOA
DP4Eou9aTrIctmEWlT4+w6JjRnm3uL4f2yxqZKXGtN8mQGQIA35giMtn36f1A2ZA
oPtaGi5i7J5wtKfI927rtrJxd8GXGXKEIPCXc0Q2IsTTHwyR2xz7dxaehGTbD0Xk
gMpJ4cMa3S1EgSGZtzJOdxMoCeeVU33tfz8yxRtWGiNX6PuU+PC31aON3BdK+DFy
yNhhjEgxMD0XVR8TYoH7NQQpMVs/vYiJordWp8Zx2aevZlIU1SHuobW/fJR+Gkvl
nyf2JkImzUioFWKQuD7/4pBYIih38J4mlD8VhFaRIFO6648ylNaOs7lX6jeGXBZH
9Z6j/u3Q8+KHe1MaXrzYXrTMFhvAkJnjaEGMD6ZFVapr/sDr4Wn5KDjl1Ybdkw8U
HWQ07fPiihi587sEKvgKP92fEoaZqyg3T7bQv0euy3Bz6xskmYIHfTqbJBJn2EMA
oOX6pGCCUCGdlubaQIRWHriC4xRQrgkzDCr9sgZ1KoQUSM+sxx0ZlpXlsevw3k5N
D3D0EGsfZfDOOlJNRvHplc5jPgiDPJgNqN/S9lAw+7oXi+Yr26mOJmGVqW895y7c
yQbLFiidkteiwrs3EjWugfm1yk1YBYbi7W/c80o3l3WJW2XWx912nKJom7AswRWU
ObwTfTk7ChNgrMclFsrw/KVm6w/4sA0zSQB2RvmdWgT5Fk+1uD2PWnYboewVTx1k
j4OZGoUg97LcCEAFFXKeA/njaopCyshYqjmPMRpKme6k6iPD1MfHQeDvPo1uzX70
Zs90W9iH6GkisaEZCk2hgNgjflpvG6KMPvmIOGp2hJGe5Qhj8WWecsRilkz1FrM5
3n4ysZRqve7Kyyd75+XiblJbXnLFcObMpzMd4EB22QS/ruwy0lmatyCrMgCN7ziI
+ja/8DVhWGzdNCHGgkFqN65GUvyiChEPhU+PBEfV+QxblyZc748jQVwKyAaYH2kx
KsgA9YmAcYlOBhmzftFWOHVkcCeZuD2Oqu3hrzgWzkeaZ4Br1F+2v38WTnSBWR40
//NMwotlDEdL458bOc/uNCyIUN+T1ich8ulrg1QUEzL0LSYgAP8gnXJ+aLcdWCA5
puDFi03ujUpZE/0JTtbqOG1sJHUg+IIkTtZ+hKPD5J14/tp65UI9A0k3fn6JWRkQ
ZUayeLJJpD1OEPkXXI2qA1G2nnSm+KrXKJXCNgcJaOhr8w0XP1l/Q8BQsqzmLCkA
jf2VoYD5MTfrghFlee2TF6AiyoB/J7ytPMKCOJpWpSLs6jH1A+xFMFurJEgB+S6U
U04qp5qqt+WmG/vo/4AFAM92vhIMhEukGPpccMZB+tb2Sv9m328DKK5UcjOc9BH0
coSbJHN33tgc7DUm+LINm9uKuedVsjglc/Wwjy5CbTRtx6r8dn2uGV/qCk7MEdsf
x9J0GKprAMz4Qf3FgoApu3/WDQhZejmwdsGTS8Pz8naTlAoGrkqA0d0f6QxdWWGU
81evrarjgIq/3OWZQ+pge+HPQxXzWVa2mpQAaMcf2PQkyj0SmxpU0JGCryySszWG
cStiRceCMYD8rVsboGnvp9Greg0l10793uQMnsBT81Udtrgv7/EtGhAaX3g3DyR+
cVvAEic+mh68NT+/mFVpqA8NXn3idLUIoZGnsQBAr9U7y/hUHTBf2vKKnUj3oIkV
Pj6gBkHgb0+LnRcWhUKW16TC4kERFeVZlUn+LXlqdQ9rKahwX9tw79BIz7XxPP7G
ZzJxr1kF9nXmoU4S+m9vZav7l67pe8aAOE4jiBWXZqGcN6Se253fuzfWL+4Wd8Ni
WIo4HLZ2BDL9jIcXTcGKIZSRIzVK3LgQtdwStFeERJvUCzTJsJ78JOgR69UGYrD3
TB5kXq8QQQfAbM65zBju281msIviMND8xuZigEN9hAAMtLs9XqfTMw2YDeky0eEX
J+se5Kyh8/SECAPxrSOINmSoKItys08ZUwOuj6nzyR8d+6dCZBJTNNXoNsDlarMt
4BBSPhKk708e+Q8mBgf0wpjqFSck+OB1XJguG68VRJ5l3/aqizmy61rJ/MUzxTni
F2q5nVQjKpdgCuJQveaJQR80t2R+P/41r16d0t13FkQ0N7V4FkfhvNEwPsbvzGHT
kat0A2LAFJ9BTzCvNrmtM4BukframDqqjIebl6oWeqqc7OdXvkk7TPDLNRtARiiH
JsCLBAQzS78o2neucQXfytQ2wT71FL5DJvSLU3xzqnUBCjN9vXZhLc01N9K/nxc3
id6CJS2oBsh4tQZWc3m9QRA6LGstvT6XJ0ppB951zmYQQ4l2XNM+ow87APUp7o90
qV8jzw6y1/Ymp8DxSmlJ31zI+T8c23+4Hos5y066p5JjJSJD/DVP7xnGjhjg0UX+
uhu3Ku+8+BkdYZBhFiCRVI4dFjXKmqcNYtTpFxgp+S8OZp5y4H+u2wh6IsXrnE84
0KUjEgvnwMIO2svCDB3CZvSctbd+n+aVHRL/P4f7XaEASKKLn9xSbGfAEwEvUuyK
Qa/YR1XZEpoPmu5+SOPbYi2dcqpQsU4j0SfBq7pr/zUsra7DqXjD08xR+2zmBY0s
/pP8DgViU6Cmb9XJ7tMSIzH4yBasN18UEJgi0pVOXu4K7W4rYSIh+GjGfPaE3UI6
L5b8IX0XIEeIQkIBsPyv6L00z/aVK2s+Rm/loU6YaxJJVWJ6NcdMdBBvvkNsvfj1
AJ4vosRJGvo1urpwTWs+1rLLWzqG/9l3ex+UDzSi/dBvTmv/icyAsFGkoXdXTdnX
nu+QiJ4DyKkQe3TvAi1bpTV7LC3oMC4YHhKTlGT4es0XFry+Xxd3fnfte03iSdmB
NifQfIEEGeJTLgfDFbISeNa9kep0C4um22HA2CP2k0NNU+8uQkUdM+sMdEqDUJb9
0J2Z6yBWQK6xNZq9Zcboa1bDot/o4OMrCMZbJ+rrHDS/ZeZlzOwJNdNamBC5ngv2
P9mnaW4Bjezu2XGEF6/kEZo2GMhxT5ptXwFdWWv6F12YifZZIp/2QFZlne/OICRb
VopJKAd3j2n2GkcBpP/Nr9pDe3HulwSzOzAY/InDAtvVdq5RlHrFXTfnHUj0O8TG
JuD6Bbx70RCygbf6t1L8o9Cq1kCUffMfGr41cXCD3pAUp0BzzQVNwDjVKk8PS43Q
sONgXDLLowMWOySSuZTVkarpHD8d+QV7/qvszBYUELVMNFxVKca6e2JQFX+EBdp2
hSVTUeC47841NzTB46ujeBx3kMfFss3Hg+FXGxzT47uufJ+IH8yF6GoAYXwnSVo/
OPI+xejEjpkB/663VDe0/d8M9fkLuW0op9kBOGsqdvUfPYXdUCLNjbJK8aBFC/x5
D231IvFZ98uX+QKsVAovzD4uZ53yR31PS5X8yI2M9TswBIstEBa+Za9XbGVVY+jW
4aGj3Lpm1t3EDGMYeGDzOpRBcZEdyOntjrym1FnIandi45ZLMu6hGVfrGlI6H1E3
F2Vi6cxb5Kfop+sgS3o9I0HcLTfhSAoSUzTGV2x4CiAa4b9Ha6ElSLr+MY15slJJ
xTiDnRed6/V3uqG377IZmR4iGOMmt/DcqbZ53VE2549O3i8efXnt4CIVGdZH3Ur2
MXkA2wLv+Y2iWjw2SfRW2mOZuY/U1yqRtRh9EijX4SzAqPdrTJMjye20sxwtxOlP
Y3+WHUg7wtFs1zda6zIPHIXuVE12WzG7U3W/ZnMhkbRhQBURl87Mg93If3nd/7RO
bMQI3CdJissoDNVYmR39mFmI5SiELXSiBntfNczVuZEDf4RlBRC1KNuU62sNXkaV
DYl9iQx/TxpRSx/qUtfT3yNZ5zU8iUo7ReSJLH4F6dx3rxvV0JHzeXO/yZk6Gr6+
OMlO3liCeSqwVHpgIdH3IRiJ0E0bpRtGdVIAPJcXySqNjpXm8xExVzat7sEcI68v
A32DlUaAkHY83Xr+MimwqH10S29bATLTxPniHbR48FNyqYvOzItVoWiY5bfakKd5
Mep/IVl1H5eqFsoyYo6r3TEIW2FcuaxI2ow4pMVMXsn3GNXP0KdoxDDOvXB6ub2m
kkwF7HAnYJqkAhtg1WK+2/hkeLbKXMsWn9QELO/hnI/tpyQDNUymL72XnS2c/lOh
IqAFPQN9yhmlsselupfvFdthgDSIbNYqinAEXk5Raqd+/8YcXk6zQdttZGidHtIU
jslWo79v6yyiyYS45uYjQe0oJcuAXulNbdMICoh/9ZQYRWj/KVOlZJHrD4M4fsns
CKBhLgZ3e67VLKj0F1fjpf/Yx0pgicWrgFd7I76gJ1II4jiInLNmv/wTFuaWbhyG
e2y+gr0MdHJot92f4LY3fZ3dDjCLNFRhxtFLUDArHqMpZ0JtCguQzOZDBE3mw1m4
Q7nUwdpavW3Tp/yvdp0TKgO1E1xavR78bbPIZLa6x6P6fQydUf+ujgrf9VFn8C11
iNdaLo4QGBmG7Abm1vp+Lba+Cq5gC2t3aT5Bxd1cmnL21MBomoHunNC+cvlRpYA+
7zYB258gfRD5R10BM+tjZIkbQWFsQahNLH5U0D42TaroynKtG6P2lXACoPNAi0qj
XJlZ2VYnlyKl6NTeUUMzAtYUMNOaNOplZRVMYsaTi2PnSV9Koblkgaa2fo9VuM2p
AolIkr1Mv6XijH+PK9R+6ATdJmaJ8mw/heOXgHwjh4T7SkMesNmcQjhqEuvOZKAB
5kvSwou+zIkcVCaiSvcZcbxC4yCmNgda8u0a+RHrg8xiNMAYC6FQqvfVFy4J2fG8
+08U3I4TR8gbMzGPPBXsm5woS40+WRDd9oIXRu6dIstjtsOhZ/yqNTMgPoDZRqUP
9aj0UdrIrOHGra7YiT4bOxtlkAFbXSBvlsN5tVir3pnLkzZ5qfwORwfO95k1R7Q9
zS/Oc6/iCAx6tJNl3si7ilx+4V0jf+SR+pKyVHxAwXfa+B1tXMuLVNTGoq9sa7zJ
ZSM+AJSWjIbDsewcTJGKb7A4EHpda9vTqv1w6EKRP46BL1jNNU8u4R6v/N7LHvJh
9UV3wHa4uNoAYtK8BJDQDa7O/se7Ms3KAieBwAV4uD/UWDi7C1TEFO4PqUSmoZYU
u4qbfMZ0OfH67p3VnGx1sejJXIgb5HACylxpE/A/mBO4w+zUhJASiViRz6K1nip0
+e8TkCVw6NamqJhE9mNPPB1H01p09wUZ/mVY9UqkstkMRg2IvHgqnGqZFKbYN3rl
6kU/AkwKrvOGJCiMSrQCfqoQ1fRmY0hjTA/2pHLNVWnmc8mbeOkfJk10ZWX0IjML
SPXpS6A6CSxZvs6eaNToncc2tkdsvZXtUEpc+D4o4LzCHvzRW+FtvHYnpTx4wBQD
f5Q770o1JFQRU8mi3SRY6ks5jirGwzbdPh4JPem6utcIOGahq5ATll2whd2nxyN7
6Q0LeYs5EQNY18aSICayHKGqdPK29lD3YHLGX1/gu4FpekZ+m0m7Xtpinu9akW/5
391HztlJzP0wjg2QeXNjIUieC/XOn6PTrzJh2XvmohonOcng4StLhjkf4an/Z2qM
gXXy0+qykZUmxV235NQe5E2fNWMSCPPWiiuLS55unBQ6a47Rgvm9qn5jYNIn3vV4
/nCjmJ81Kqv6J8gTXKn2rzNUHhuKisCvi6qU3W8Gtv5he1zHBC6Y2a4LlHef40T8
qCTI2aLuPbLeB++kiqjdX0DKXFbS8uXGEdiMVbRNPoR8sW9rtzfImO2Ro31yY8Ru
DdLSvCayGZhqS6+4sV0UyuKcNp/ckRAeRiqCXiKs/WLnDB/zU6IoH6KFtPbe0uKn
+2ZqPrTRL7y8v/4P7rHdbfhFJ80552sXAuV9x0O6cjTU2t69YefP0vI0FWBU2fM2
xaEcBnf2QbaB0ziChJtS7nFP+4nwNnKPL+1Xo7suHHQG6sbVQKKDuYnUnQDGzQsM
+VHVm5yk14KAJ299bSdGOzZc4R3y5Q8ROg8sg15vqbQAas+jvrk/YDeYzp72MVC5
ehJVqQJGW5jty7ItX520frbFvJ3zFv+r2rzzobnGgP6NlZmwdTnXz/T92IPtGr7X
xbWHpfAC6X9Nwb4N9FhZfT4+OK+AigubOWCXRpIjAO2LzkvavRY0cO+nLliKTN2H
RuMw+UMW58aBU4YqlSbH0qNEfPZJQNeIQl3L/wBJO7lUFPoqYDJiQ+XSKC4c5hXE
dAhOEj4kJneqgflNjriQqId3b5jRCJVDBh5GPIuMv7wnD7oOw9wFcaH4WpvDuSGH
SrmvHOZJ/ndxvGXx2NJSasVjUJTDx0oi73JYzFJLDgWd5iMW7ZlOYJGqd6aG4cLw
5sJs5BYic7xJJJaNgNXnpbshQAe3c9056d+zrS07B7TJXUpUJ47i66ezLlITtJFN
/SA8uWQO3sDhtTjCy+3ZCEB8cay1ftj0lgIeyYVM9WpTa/EspIJpC6g7BpTXZxfv
GX7+RoAsGSEKAtcKr115PESSJVjpk6ZevDWdSyjFgWum2CtXYr2YxyDsbWgPW+2A
UeF+uKvd4MWPskrdhfaFgLwzqm0B/4wz855gaWkNFM6CkIK+4M75d4TgMtyQdhs3
K7j1G++tROXe3h5kMHbgec0FyAWvg7L3he37OmkfZ9IZnlZC5uDr9gpzVmMtOiWt
atoJUsbWSYGYa0UYpumOkjtcK2QPGfAuVhIArvO4ZyABLCFfZ7zCia3kA6rnRl7B
n3OYpTTJ38JhHLNmXPRGhRLa5RlO3zyKX5oYDeo7oRXKA9mwr02iQnGlLH+Oa+1n
tIZO+nqKWG9ErWCn5u37Qjms/mNWKhHvWcuWTYHvB1N7zlL/gAtjNNZeyEbbIy+j
m0u7K8CV6fgcAhTGhp/s6TEFKeZyj5GG1JT+i+p31CYks+nNacvTfxHDitFu+u5s
3L8J8DMl0Z5yTi5F7kvmoRqZUxlK4zVSQHAyQTWhRGgpjyfCEAUnGn3fkXfG8O4H
hKNEjeRRRw8zOHxQBlho4DFTj4K8vCDZUWTTn3VmvZCAyuFvRO7upAsBytogJFF5
V+B2kTvhcRiMlKA0HWSUBnanRXBrzihjaTR/rrzTE1FO6p3qCnWLTJkh5q1sIDcf
WM+W8gfvGIa+ZwbYiWyxMVn/mU1VCvpu2M/2KKMHsYpKqxrBFUR2VoimAzj4kUsM
UsGbzb1zN60sHI3d308h+YxyJZ5anrj/2NNBYE1HXPS9oLHEtcYYRhngIGaJ6oje
kmm9xZ4tEy+y8OMlfadXirV6M/LY0M4vkr1NLojVgX/UhhXLoTpukSq7VIH8JBEP
U7WGiIReiL5XLgEh0IwaecAZcob2R2AoYwN4KPpKaaO/GJbPk62EUGuSnY/yxBkX
XdgqId7IO+4zN/1m3usmeoLDPQThiYcEslPoDexv1Sreisxyp+kWgrsL59paR+DI
26R5kF058X1Maxx10t4cLwiAp9v3GE/nyHBmeezpjR6GUcTQudr2pmNPQ9y0MTIY
bnupRtFMIaFDumcylS6/uiEQw0UJQqX2yNbSuxsP3XBw2s7p3eaBJs56S/zOE3N9
0ibAn8Ikr92hXyVS2VtOtqpuZv7rc8lPqhV+x87dIcwMJ/7LnXOxmxLh08O0BjnF
zpRd0/9hLHQZb9sXY4GbpU2SVq11eWB6a/npRV3g5OnuNvWf79ODeuauWqNk+7AN
hjp/INvw9L9NE7u4W/EWioKd5vAekQpI1UOY00ZXv8H62gtGoWMEImYSWXP0OUH3
ei81r4YZzZbEGS1Uhs+6++vf/IyM5klhwNttD1BxAPMWgNORy1ha3PZHHgK6ov7a
UqG2o/T9mlmocN+l4DcsFeH/lwXlFJCNsSXFsoaUycjGUb76ULM/S+ArdRWp5Rp3
b/UnLwbhty2tI3wAcMQyowHtJs2eba95Chxxz4PKyEsAjO9XUq/3WvGoLbING/9j
MBIpH3ABX7VvPgQ/4g6JkYAQm5sgD/JbJy2OU7RQjHfXYMFbG+72jCGvS8JAXIOR
D0m1XgPC0HbaJ0BYLez8MtfZK+uftSlrpzlRhUuaynIManyxmuSOi1E2tvWbtNOR
dQzjaAIJUHeusLnrXxCyVM7L+U7r99t9jnlVJwl9OjhogqmXNkci+C2tJ51WBpvZ
rpNTxr8NMGxLeHtMf6SQCk08UnFzpfcjbN9tkYSbcNlSWXRZQ+nD2o71z7D0xokD
qDhrByZN+9Q7HQ8CEkZtsqrnrtNyJOmiW7ZqA4c47unwo8nA4SyPyN+6nuhW5AiL
nHWURNg+P9ZGMdsPv1i7jAFynXW5lsgBOmp3CjayZUWyHzg5GF4UX9V5DlN8gfO/
WJuBlIM91CJVx924cFuimc4ql8k+jE2gCRvLX7Bwll40Zszw90VdVTgY1IiUQa8J
lUdNPawvVW1SaV5IIXli+wGjEvaB4TuGXLd6BPVIAgGET1lb0CFAXPKMYVW/F5KW
c/d3HJ9atCB9SxloNd16Gh0PyROD7CPACk4za4Sl3z/qs/TNcytcroCrPrvKctnX
xj+StO+FDh0pl2h52jckXjbXHVZiWnfanDe/VZEc0hLyEIvIQPjWz0qF5qTNPQnU
75tBnSEvtiyTAopV9jPHl9Eo6f1H5WjZQlebr5ZIpwkOMyJXH4GUAU6dESL+4ZhX
aUqf9TU1glYAQye3G1unNskxNxKbNRuIGRzIn/ha1M5lMurC4AUVAkGFGg8Ztxcr
3XeCow1dtcD7KDRoHgJdUKMVDobsMBVEG9B5+TMEO3dt/2p96ZgPAKklD79O3OXa
xGHYnGvq8qrvvUrYdrwhHL1UYrw7Dez05EZAUqhIHAr5ytrEkMM0X7JJkq8kEzuB
UMCxPVBR86VxYjbSOhO2om3hDbf6DZ687dc33IZEyKAI+vO8tfPSZJv671sMazQe
VgTdlIF95+RmgJ30ATGLYJhZVEikxJGZor9nZW8x5N9/pABEC92GDCg5g7utOJF4
B09Xl+lzLnqiYxndwbB3ZFk/LDuRs1wacZ1PVWo+9kEm0QEtEb0NrKmjJzVA0D8H
W5+n1DS5YU92EhfHWCijGRBsJnKvsqaI2FxcXRa+J+tlBRiFkDeIYznw1zN4okkF
uwqPNA5qNCcD3TR3nv3WkM9Y/KdUgZBD3t6adNB/FaBh3lCtrgURf5YYtNqOCkcE
QeZcyZsau1Kiy+XXfOMNB3/1iv2L/qKEFdCs5rwBbz+Gf45xLdmAYOwqT/TEohgA
5NRchFO2/WF618S3FK1NMwhuWgdBYQrRNpi07HP4g9O/kqzvo7Id/IZ9GMUM94bB
VT/chQK4zv1CbKZa/8ZG5WroPByGZBICiSHwAYTD/eBTVTJaeKDiFOxrw4Kq/tON
cCG+2RJDC0U6ra5brz3V/y6oHjFQQ7wdbPVQtRI35mkWeUdNrZLdcJa7NsWfW1ER
cgZWU8TIL2f3hCybuuW7Vt2Lo9bdLl0dS2uzkxoQ5+u/ohzKkrfBQh8KMbhFeVAY
kGtnzS2N7LGNDotKNoBAGgWEZPukNL0iEPHrt2h+20wv3cUbl3GqxXYlVLyxGSTa
m14UY9cVmAuhhKgm3GXRATqH7iXu9Em88FTf9tA0AfaCU7ivNqBDvv4wU4rBa0Eo
yMhtqRdsGeYMpy6uIFyimn9bZ86Y9vchMxL3seNmEHE+tISprgrWmz9pL+rUPIuN
JYCAc1r2FmpUypKcmhEAOl4grBEv+iuUw0S3QyrJH4Dckn79FaOs7gC9bwPkWYEv
OjpMu65GiEzYd/aVII7OJWRE/axjwzEqaG5lAXDMZyEcIr5PuDDprTaztNeGnO7A
/+KYXOOMUoxMLSyHcf8PhK+5Oy7aiewqhAU7CU95wMMoH4WV7sj6VK3jYge86+Ji
mKSmxMhrewgrALGUisOD0jKYnZSmFiO6DunIf0UagnaZUsnvmVH+gbWJlR8ocdfe
hQKHObV4zTQE3/qiAW+VFsefLLN3bXdqqheVzbhEwjSKuyo0ayCHisfbBhsCy5wa
caHGUUXnhm0opWrm0uaBfcmAzF+QQ/ahhwRSpbbquEboHTccRodXvJ8UdEsjcZX/
W1aI+Gcv7IyKgv8qEQKz4xHpka7nqLYyWWrcZ9+ASpic3lLm3gRKrEEcTkvV48sb
37IN10rZ7IaDcV+Ls2gcLO6bqFD5fe9Rh7pi5ggHCJcoO0lCSdlKK9/u/Mt+0QnC
Ahn/xzv8a8Jo1iKVhhdjK/xWmIlmFubnYPBlJD/No2gvv707vVUULMiUYRV/Cs1L
IjFvSBsEEdeyRtoTtjxu4+RP1Njdw1nuT2wqpFcNE+HCxAlYeFX8g8xj69jwYPes
rP7wubdpIeaEfFfpbzGYgWsdlqkjpkfBb89PQjvW28pX+IeLxFEuYWSmSVI5NlII
xawSGr7R2IHi3Le+NMcXCy0snSwY27dCi3g3HXGii2tD8r3YHfLwn1124kzYqr7+
2/HZScbrGLrc4MLMPwucinQ8NnRs+lMGhnxPk+sB1CfMYa6HYUshzepqDvPC8QRT
y+ar9SwSNXVkV1Q9rUXB6yo13bpgJXTnMxEkJZf0F5tzeM28i+ztuJUrdAv7UYmD
FJOfy1hdvLWDAJBa178JZhdXvgztGuh4VtHFZ+SQUvHp7niR+SN1Nzyg3WQ0HaXL
kRFHsUrTyP4jeeT3xoQiUWko4HJDthJkglQdcqrasoD+kgjGpMCgt9/F5+AqeAh3
FCo+TJrqGIazHBcvVJxOzZiVTaOpn1lQz+cgwJgfOiH3Zjgt4j3Ib05PrWaa4UCO
0llzP/Q+nZFaqN/x0DTWozh9L3UgCz4jr0ZAYVY4RQDF17jfs4vmf+FKnq92AJi/
EeEcbKdKo+TNFGp5QQuxcNy+9bxSN/+QTWcy/qdHuaeHX3nMoOT84OqQ5CzDbsXe
s+CMn9pc1RyDLIoKXzheL5/uULlSx8p5OlEjcvuw/RIHPp1K5v+9HTPKk387JrZ6
eTzlugrxRlo07IunEvpD1QGYj25eLL92QLJ+92K9WBgf9Fj7DuRx0gupQNqaZP8M
usPqIKTlHezU4ueeT6wIWFGVGaBK/Mg3bwgniW2uO6ar5GKac+zyNnJrGavW4CAM
Nf5zHLkzJHAcu8798gbN243eSrferfQxRzFxNYsEMUvR/7gSdCvXhf7Si5n9YWg9
ToWeMS1L/y2nJE9x5qhAa81Ew3I+x2ScNZIeM4knTJKfB03MUX5zok8SPx+5Dqu5
icD1jX49+rVmGLp+jtNGvDLWkNZwt1qMmhOO2dSGlz5MfrcJONvbe77qQbZu1/dT
VwfsvwzjkxTPIhp4Hk0yjHbiKNOBahUQrttP32O8e1oqPVi5Lix3UipQcX8OO4jO
blhQkczOtpPSTHXi3rLcd7iwkqkrmk2tvh4OqvY3WwkEwvGljITiAciATse7Oe1m
ajx3HFl3UbXXKl9KTXd42oqFf3YVEXT7y4ZfiPDRt+cWlp+/xpzyO283xLkJR+Eb
nFGMxDYLHpeyKoXFJKwO8p0tn+HoLDxuGs92U3tTx/GDyAHSdsKVpibQji9P9Fay
wdWOdDsuEWqpqq4pkrfC30l/FXUrIKXbjagQIpuovdrv8NxOjGDxNkHHrUMFnfVv
rqCRhZryjS6KoeBTh1nHgoqzKCcJawkyKboAKuMxzQq3cpZoP46as70h/dCYiE8l
TDHbEidptpdsZlB3aOwu1wcyih758S60XfvCZqKBw5ipWOm2qoiVSIyNc2DTpy4t
TQ70PJ76AmdjvE2h1pmnxumYRZYALQpk4tZl+N4bvEODsAQpcvtd7qZg6UZydZHe
eTxwPSJ1UAtLiy5HcIoSvaJJwigqLNXoq+jeYLWPGHr8cjDUaXuZZOYfF7bOYBMZ
/kguxZ/5scuySvgRGIQSSEhNJaG8z7RCDsp906mg7Liurpdqc0FSozaFD2k+0ehL
fD4GTxaFVwj874dM704D0sNGxSKeqh1B7X6VKMBJG6nWJblmN6+MWLo+dvbThWXG
ZE6NJUHZjuf9PhPdLnq8DG25k27ARatYDNuBtDtBYT8Cp/GyGDc7X+m9i6WYDTpH
IjhtPWSPQbMkcmMHVUteV1YhsY9L8vC+IissQ/STLCjDpot6FO+eRKFet1zw9E6y
yutZn1kp27WWCZKiDFRFGC+KQ0aYzKPua4o7PRZbXt4J85/hG2cOgFoL0aERxbKA
j7RFpMkoSkJwcSLQRP4EyvTFOCzund2fjKtD3Q/VbkUkKog4toXNJQduA8Z+F94f
Xj8GvcScPXUJfygt4FzZ732GXUEKjV7ofmn0l/3sOdX2un2LBgq/pIlFaoITUJAT
qJ8XvoaBHQz4EBBfwM9lt0WRhEdrL3OjglOhOFPoRTbh2vaw2wPpQQBfr311B96k
0yzU5fsR7txCNyn3JWKGf7iqwF2HKY+vGRbgExEld47bliaVovByTV3P470G0FO+
HFaicHWdGqdKIut+H/XPhqZ0S+hFxLI9dXI6SCp02WEGTkbWxf/MlIsx9xxNDY87
iC3Lp49lGyBzZS7viteyf7MgeBCrDh2WT0rT4dlF3vsrUxorYkRjIBy0ZThxwkRY
IWJPM3grLIXKlfcdyVMEV7GeyE8eJWYhKSWB0smtM1PZly+K9Ofq38nrEfcTYxGn
uiLF4FjerZsBOwOD58WXpzJaC842acADCJU5T8WMVLJskDnu6/9vFyhdzdTqwFpR
r5iqeoqQkx9HOjij8r3IiVjE4Gyh3UpAegJKFfCnFU7Oi0A7/4C/f0+4aU2AYkJ9
l+66xudnydpj6juG3fV2eeBbJMIVoyquPjx50U2WB23gYB3mlop5u/IV5nwoaOrN
nTewbksE4XajvXnuqcl3eSUka0ehTzq7yiXryTYuL2JkyasRJ3slF6+zlYk81So6
iqoW3a1jO6Ij4yBLCRLB/IhQ3Bk8MZSar5HnqqjKSJG6YUbUPtww7KJjt/DapYR6
zMIi9HIf5qaqUEGKxq+ocHC3Md2Q414WWVx0MKDMuHYtDN60c9rs4eGVOD6p8Zu2
6KqkZDf1NVm2sY+TYsYQ1ht4m+TURgA9B74vHieAMWjXofvukbZtbJI6pT+v7iJe
UlXbXq7ZKmUmk0MPdvjWPoXeU8oKebZd8uMFX85xnOs93cpLxRSXcOVNRPJtKorR
gkG0a6EcKcjEu7oVpjayg+65j1h0Hd8zzH/rNSKNjZKzSfKFI7QhEHL9Igvl51lV
M/doBzxkDx2QqgzhkWFE/WRZFM9QaxbrDgKtw0hMoKRN/l/y1g5NXkM7N70BYgVi
8bwFhKZJnSEpKqs6bXaDufhHVy0wJpTllwjfgQP2JkxsG2YqKDfatfML7iQA/aXl
SAvPzfBAt4pBT213EJnUiSfV0KSTo/3+S2+jDlgW7hGlfg/cDnizQ28QBQalo2tb
A3OtJrHIfIJtlrtSvpNiPkG2lgHB1A9v8+hdEAPRZKF66QWoDbnH89cz+XZH530l
vkGK+EU3QU98cTTMy+RHGg==
`protect END_PROTECTED
