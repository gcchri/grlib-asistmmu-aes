`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xIGOEy6Ugbss0+6Cx5y3//rfLHd3SXPTchrWCGXbP6hYi6/6OU+Pn7AlrLaBYVa
Graqg8o1kVFKUSF2IrWD0G5/amyBwqYjURUwcCQHXhxZRFhmQO4x3tTMWCtQrrAr
XptOg0Xz5sp/eFdIvu16p8HQvp1OACFMkDE6KdtqexqnsxVENmQ6w7WmwBU1UF/T
Pek2RJF/EE7vk8Yfqfm7O3qQ7vRxGk4Xxf45jOU9C49CtcAJuf1NpGkoiXlLY+BP
IOkcwZQxoXzcJAWDV+TLiSXLzmDy63azJpbOjVIViZXfkh8mHJGfXh4kmL51kw9Z
8ko6Y+U8vpOiC8E3X3v4R+El8tkK5GR3Entff7CmqZaBjNVtyK4Zhekx7k1BjSxN
nV6yW+OVnZQe+kgpOphPv6p8tmXVORJ+YCSh8TxL49wx7j3d+uAuDElwH6KoHFCJ
MarQ2I5E4xEjF4dcozMxYEw+unIy36nCKBbAst5637jtzxGbjwsgQGfTWUaY/j5E
x0gg8jG3jAxxO2Qdw3HAd7R9kw+6oy901KXslcRkQzJl0lD4iNZcwlGQWd0pcoK+
nNLAdKaoraI8shiPCei6buX/AsHxpEMoK54CKH2DfGRh7zqkI9iT4VYAoLv8Xb53
0Vwnwa7SxkfKJ9Ib1k8G3LUShyTxi4WCNBkVxlMSrrsqaMqSVV1DLFVGO2NgY5n7
E+iY7OPUVuQ8BiM6Nd2mfdNfmV+6jT+aRRaGK3jszETes79a4HTCDHezId1ryS0Z
zOhDCdNcO2BP0YEXpoRH+3sXQ4t1vOg7rbxcReoJ7de4gnhU8YOxkI0KsMuNYxaP
His+uqV4UILcUsms3/LdrImPxbrTXXznei7HPKiFCrdEGLHs55HzGqU3dz0MvzPI
BjtEmLg2wzmy+ZMSI2bfUzZSyifrS/7qDsw/vYXXjpGv5ePsAmLGMk8TJPa6ReeB
`protect END_PROTECTED
