`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1DbFgqAftzXvlmIYN0K0wCt2fhRFtItATWcmUaEeYftVcUCuj+ONTQc5SOD9TDe
eUb8nIiEOfqTMT//s0tZvfi6Z6Ra6g4C6fOl8hXHAZr9eAyT1o+6ogCfweG8BXjk
G3eJNCPpLxBXD2C14X8Ld8D7XxSZCbJz2r76MsaPRVSb1jX6T9UUpEwXJUnAgkBS
+RR76zM1c3FxSVlQi7reIrPLknHYpwwjgR4YCnpDgt1hqUFsvz2/MoepFsDbNWKb
tsd5Nvo1RdIz0p63C77kl+A16TS/nfpqC+d1OnBlaT1q/56jqo0GdaC5tvgPY9q9
CqUIdj9SEVK+Gx0TfNDAMH4yQMD2U0mJDIsiPb1myKZOm8s0rJ/LI6bIP9GIL0KV
TlK/7uhRxNEJnAXmwVez0Vq8AwcMQQbl2VHstYL7znX3ct+gokgsmcAruj7xgCCg
XQxKrBj/jAtn47b5+3Zw1IqbtP8bXDgLEmM1njYrz4fj0PVOODKS2WykHJh6blbY
KoYHWQrDJK0EYfJA9D5ovp8ST842LmEAe+8qwP8pU5F/mXigr2zRjp8H182010L9
L5+ohcftmUKJvP7mvKGAsovR83Kv+XpdUhJaNjnbqD9cw6HUpgUKL7HwGyijPaX5
kgYt6J19Cr+LHm4l8W7VtQ==
`protect END_PROTECTED
