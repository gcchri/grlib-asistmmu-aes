`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69HHrKpTnEUYPIThdyacvZIqWw5+ygkRe8f2nhTRWsmBdBWVfKRM3H3cOTAZNzHT
MuOYaINKtenGZVkQPvMS6L0H+QzcuXdDJtGZB1JXcdh7gGv+g/9DBFfWlQzmguj/
kmmf021dhBZYMOgThuBcCI0xv3bNBbEnM9weoqb4zub1C93A6udRKMKPKbF1Y1MZ
2faUHEFxidwfTIKwX6lsQZoCYxQyHHeUXaN0boWSA0KIGZA1RyGKx9tY3YR1IyN2
3idPAPvZLdkoL25Bx8UJp6emgz6HVhxuXc4aZ2wQuqSg2GunY2xp57oPiOL1vm1Q
5hjrf+fpkwYCuDs0HCsYyyJ8fsXL+3Q5P5bBSCiL4HnSHkULV17RqSUunqbvn/wS
3DaCqmGTIKpro5UqmMaRfMja8Mk16U93PFpbOSuS/g65N/Ay3T58JuUiBenNxRKK
lLuiIaavBpNnKn5hNtZZK7VXDxsz4aEn8JuwYPOsg3o1Id+iHKaYWNRQ2mBZ/f5/
B58LXf9sbqekaW4RaHUR4lNJSZFdWES9CWrgOF9ASeHCafjiD9lX13GJLiEjJ9aN
XacbKEo4KVEFNlVyWqNaiC0LQsfKsqlmo6G4yUSJbfOJyMEBF9jy+/t/dXNgPE59
tog7oFS8YYInpE64OIMTW3BR52qlD12B49JPKh0ewfMpiFGenGgb6elzMnfoIZdR
eGrTiZBgwRq+wx2h39Ak5NSwxZZAHphrA2Hks8kmDzqHYHElUIfpREj0ul9ZWO/O
OlUy5CJk8fs2ATOPhTGkm1QjJEzbe3BKQBtgbyelD3lgsHwDOyRzoxCiUKc5W0mI
SxQxPzgPqhjct7ObdAQ4CJeBa72LTif8IFaLaPzly/uwMHb1XdOxIFas/geRLbEM
/Cz7ukN7z64jJlYAnA/4Rw8iDYjEhzNO4X3O2j+MdFDM+tMyPLFHhdMHJzWH0SJ7
eVd3TwqSrIUfnNjQFOdxT+XAhxYC/9cgDDVSOzGx8oIRCReEmyegqkbrCMK9qzIh
Wt6YRYRufVLY/UD9DqmiMqH+ljshh03d/NzKrK7vLRFOZagVg3mQVdg6X8c9qiUo
W+0V5oT/eCW+zD0nlKIB4sSm7r3ZNy0jDikFpIh46wxLjeqZ6tF42sOzck8Z9DK7
ggOtYaDNFcEmmRiMlG5PBIXJJpOZOXwySYDBIDn2Hgz7yFIujJk0ctGDpqN8kFxG
bhMk4M19f341GUfmLGWSHh9Yg78Kd216rtlyN5lN56UAI3sHbFgIaGLu2cdY89YO
Q1e8JBuAE8Ad7JD5RHLtT6LZYdRKoBwbpIoLhFdvQecMG3D/3VO3a3USsr72J6W8
cuVnAKpH+tGFxo83yiXxSGemyawc+RQfInWI+QpSwjVGQrrN/vs+YoXgQSFJr1ov
/jInMD0AwEaUJ1wEHLRCPTpI6q5UEazt6KW4178u795G8LOW240e8X7bI3OaKjeH
KLPO6RLrRzVJo2AixxrRXln4SWRcBvE5Mo/YRqY6hlPfexMvcjksBdjNRRvtdlD4
CfMdzrEuTQNIho4sca/BEIbMAlypKfrnI9pVsUUc7OLX51PtT4wogTZIfsM13x/j
eux6+OCWSI45383juEjT21ieKi9TAEcn5+pw48KsGnJZi0WYUNfgXv/UV8c+mRe9
fBQZ8ZB8i02Q4OJxg0T+Wc9Z95fKSbQ1MgTpEC+iXqFieJcMrc2OTBofLH5zewEA
gk3epbcpVJJB6zrIaQnO697v57vVvbisEAigpK4CPEFkllbQRNaxqMDdEuE2jsyb
h0N/BSZrMcPYFKugxEkt4Pk0tudcXfk/6aqmyQp+gizt0ZDI9qXpkvaIK+eoMAW6
QFg2n0DExmSfbfbC828PmhFFmT2wG32V7ITKPf9apPnLzRHhZgZ5gGRELHmR/jGN
OGMsoI+LOB6XNGs0w4WwvFBDSfaRQ+4yTOqSpqvryo/Exx64MNPwIApxhGBepkaV
ERiNOC2C7qgBNl0tKG8ibjN7BhDbkNz1NPeCSyLf1J3nB9HCnZ+xlBB3ueF4TOxe
F9ih1xlqaJGPywMT/M3/r9YpPS+NIsqdtL6b0nqbljJl8xBmKQ2nuRzUQTpcpn8R
NinAnSyXv5soAHXDWzfJgUwwDuQu0+/eir5e5dpRqzLeig/Dp1FkC5mOcRukrE4B
Y2lDFZUMX/OFWsNQbHUvdG9hh3TyERpeQAfpS0s67ulDilCikx3OWOwiLWkhYwxR
YHr5Hlu1FwOqLsv5I+w7QyKNmAk5QuM3Kn8fscu1rk5W38A92TPrj0hG/U0HNXJD
KqIp19U3QqODcYab/ix7mEbs+EZYPfyHHQRCUSLFZIMwcKoOFdD78ORqZE7PP9Yw
V6loQjWWoVvjRnA2rFIVP6dzjMVsA5q7sw5K5ceW4PXDQn6NF7jn6NHRjIx2hpMq
pVCo4+ScIFiDhZAzpgkq1ByVEdKagW2ULdTt4UsN1O/U9/AnCnuW/mAV0gyLnQoH
tvg77zv8cwzS00aZv1tkzeQ4+Y6FpjUgTP/OzP2HjIQOONgkoyoG2Fu90kU+Osax
tMMkN+AuQtNBJymqklx60Xd/D6yOBv+feBm6WOudW+lY5Pv8NuLR1fYgjUmec46b
PHN8HYKk3ol40w9BSO+vu2SypsMJiqnTHtOOnImmMp2SP6JLo8F5kUbkAKb6koVC
l7BCliQbd7RwEtunJ9FHYOLzP/sPuGgl9dVdi3Kj+mrUYvL70gUn2Gvuw//j+TyU
N37QEwfbjMNN5V7D0+1mjmO5zlrX8O9wQErPo4H6rCdDRnvwmYU8XTaprLzNBkTM
AcQN/vlZhxxQ06IoI39KydV6kBBSlhalafDTk1UoXJ4YWfu8pMsDgor28M6qT3r3
iUwLKdQRAJoo1LPc8WyN7thYzYoy5bKK7RPj2Mk1ZGJHQ+9hcLk+Sy61CUMsm7VY
isG8xxBgqZRrUrYGicXjacyQKUg5c47Q1bHeRrddG/XS5HdmUSdoxj8ewOhjzSeL
R2rgAPAy5k3NZngHCN6f5h1vWHgZ6UtQxig/LYIP56VtoXMWbPjo9g985p1XP0cg
ny9WcS0386hHyoEgxJf2sadgqyAm6KgOhWuXEDXCELoUw84d2J/A0kYAv4Fx1bo5
EC9kkPu2+o1dey4FJ8tl0GxrxJbbyGMRwypBygqEVHSvuCO4qvrFSRKjYdWZuwgV
tIKDcswmKKO3uI0jezbsDST0XSJzQ07jf375AGY6Dt4iEK+kcWb8g2zR16a2iLZY
Rn1INDkH1K1F0TqJWUtrwP1go4Xd0cn8NoXF8K9LV5JDL3gGRtEswagXOgRIUhMi
Cy9466PKDq76VKJG0ZE++IMmp5wIyx1VBLC1xQuvQ5zKHT3ZzQ8YzOiYxFzR+Xlc
z1WmP1psH49+aJ30xLCH/68W7eYmqOpGREsL0YfOD7VRH64JYGKH0wP6SBA+HIWE
uHN7eGRAYmAHO2x1lQ6u/HiReqxgcOaReIv6KHx5VUTdFCXRr8TFJb+yb4Y0eXnr
e6CAJziVNOUZV2B2cFjfXGL3LcbJlenIn4xTHdTkJdIotKCl+vUnrQHRfENFqeON
ZMmz4AyJW1gSiihKi8bEvXBHeWYd8Iya0QI8Cw/gz4jsYYdgDTySP3go6cPkh2nH
POQQjXNPwiUR3hirEfbkiXHPl5ca56wgK89KA5xMTcbgw4jZUejMsdmdB2nLtxLE
oLJAlh+LNe9bi3jri5GXdmok1AH5p+eGhIlh4KdaNVUJzg0usiQ8uVsSf0XghtkF
ckQgOpJlbY7+MTxi9dVsVRXVfX7aH9hzP6Bm2IUPNAsyl4kwj4AKFppQbV/T2HW9
8lL8YbU0ILEfNG8TFJdv/vsk/qmq13s93yJbbF/cu3qT0a+8/2X8BrCLciUzqaDb
MlTgh7gCOiWkiXEE6feU8Mofe9T74j6GIB1Tlgd2bYBZr3fYc+Upa+e5ncjRshYy
eII/11E0iLJPP91k8aa41VPIYCpJ8b2xOxJSZWki+om3x6yILbAzYrNFjq94FfJF
63MeJRU+q6e1bZUG4Df5x2nE17KkJ09ntpgaG/IklrTbHQ9pIQLv7wMSK48cZF5X
BGE8gq0tWokApb3vBLescVuHYmaKiroPday8xGO9tcQ9zXgoV8YP6yKYop2xFF0C
GKzet3+178pwwBGJgBpeQZNf+SWan6EUhyN0veJjf1vpAXYZqpOOHyW13lh8Y/Uh
KAdxMht201fR8ZGwGJoKTkjASg6iFLd6fshrZ3y5fQSMDahLu0UyvIDkRmgttdzM
cYtXvIUklmJP2dSpWgLRyUFNuPfBuJfJJ7XI2PsLw+A4xaW+c3kskXW8M4b5KNiY
bBjfgCGfVDgsqFyLlyPAFm21osx3pMWSicRI0sJKG4qiCxU5I6huzRv+3rB70vfB
whg9jjmC6jLuo/SipbyVGTf2HR97fHglinuXVDoopvvM67S0ZGd81L0zVZJKk8Yj
OH5PHJ12jHbPRxxKaTpYl/GyIG/TY4L3r89uS2TOjj1E+lQj8lxN+tS/LG85Hu4j
9rb1hMc0u1YNFRMB8Vu6BeyLjC6yQHt8Af2w2H6jROiBATQLyZJqFkzV7LYdDKRd
zrNGR/0XCCeqetvqAQ/5jJusU5ZXWqBG1m3Yx2LLhv/49vw/4ZpOUg0UV8UB/RQP
xmGdB6mJzMElz43AlUzrJBRTLCZOKsPBJDt3bAjuFoc4fpKGWRvO1MGn0wLFNB/Q
Ipfdsxfa9LExKgPM0CAv96CqWiwqMJyF6+uPh7HdvFzk/ymL6sUyB4x7PbsXq1zT
1tt1vNWxAEQ9dLdwAaMErl4u+prLYIEO1n0DvIg4Yq+GzQc6fewtLdannm8m53KO
Hd1BQj/68MzEn273oiJtvFg04EfLZDpXNSfNKibvuLnH984WF/tnoQscSqf27nf6
tjTqTXId8ykToMzPKHAhs9eyWmIW2UlMHPvjxZAJV48ex9zUTCwfHie7cpYnL7uC
aYNTe100wNjE2QrqsnUzEfuFN/HlmKvKa1IqbnBZm1bFTBWR3Ac0w9FJLrz+4ADV
cVsRxWltPc8jnrKlmHY5CuAegjXeTzhf/lZoyXCgmGajbhsaTEwenhqvOZTaoVBh
+i3LQX3cWb4kwrCizR0dUJNNBUVLDU5u22Glx1Io0qvidAYRbGuzkaqhDy7LxlY5
B7Yc/Ipuvp0ZxI5/51l0e5Q6GBKZpP/sWwTsgpfTXqi+RuvjXN5gpi1kwqYFLPRD
XFrKP2238QcffEqjUPwxd8G0KuemCsqcG/aBBDqLBBPs9LA7ovtOSIOWbBoTUI9m
dJjD6XZyl5CJ+hogKx66AwdIdYpI8H79QteLSCDlVZcD0IojnIwLzspc6RphxGxZ
7K6jloRmFl5hGS3TxGbnSxX9bO/+ovZKxCbnKayxa86tBIqxDcyqIaDG6PrESLuh
ZvcjZU00rJkXznW48/a3fST4SgPJdsnbgEfqYXjEGw52mjLP+adj7B88VzXLGEdw
p9tKu3mXxCT4rtYf8MIeYE6h41MD3R880L71dkZiaiUz1VRIeScMgYSdZiYfbWn3
FiBUduDOn9CB2b+Wz20b01TlZCeBEcZnRGM+AvfMygUcbXFYhI1IZHyIYhwVwQ/I
TAf6PhdT/OdH3P9tdu62wkgqMhoAm2di6jTAyeuGat4HvBd2JJ8UvcoUMwA1EGdT
BrfJMUoq5LobtnYdOgHbrIGhszT+nWD6dRU3FSq7ybYn+bZsI/AXtpjjAsXgZsL1
SLmtDkoVkZSMFDy/EbItBfCzUBGyzE9LPlUl47gH7WVqZ33CfEJNNAWFmK6Ssunh
Djzo29rmyBgnyYD+guIkxIiOLIB/niomX3ME7/tk19TRNHLHhMF73XcHfpJCoNHZ
FQlgt5d58rWEpAuEi5z9UwsN9fme4ldzER3kNktbjX61T5FWgbloUbf7SVhrIpvy
YEdXqN46+NgCvGEfpQZ25Eoz2r7kIpBU5qERl3Y6pelAw4v67ASCoCQEAHBoBQjr
jSlJ12u2aSudQlfaCEGGKAch5FsH3uEIRAe8cRQrxNuOeM7IaPE9L3zTgF802Lu3
yCuGaMYqMfyyuJXULf1QkwDyehEXTTTkg+M4iYWivjCQcQNeujbME+CIv19vVwb6
BU/quVQ9Bte7Gyq66rybWXRfwmpzrckTgoI2UqbdVGypeRVc6IIzZLLuVpta0JBM
YIY+kEMouNC9oaKHnWaxfjVYb0LE8jQzan/qsNKXxPn1mUk8ei14GLh4h2unFt1q
eHI7sVfH4hLhKrDcNVf3NXgL8raeXR0dzhJxPuXfYfXneAFfmmHJCf5IA98bXPTP
BZZdV4C156chbdLBkLTcGEHo4vWi7TIeUvi7W/i6ofEljKyWk+xcUVpBScm9E02A
ucZOWFi03KpqmjdsPKVYgVBhLci2OTdq/yKug4DmeIHXHLsCoPaZ22sbd8KdY2Vs
zLA1X6T+ZiJcf2FTqYtLDA0djCO6IZGiSYXcFX150TcdF0EpaneWmSKTvofTwnRX
4OQFlGr5NmmD5jeEb3JkU42cO47A3WqyLotFldA/trs5RqUgrNjyEAc6yo3p8EqW
QoyYpr0/4cdMcHWzhn6Bfdu63DAT8Tl5MkYToNev7ZnRDKyQlXq8+Tn92BsG9gKI
CaHUZ7syGc8aFPu2iaMqWNumTEJntGlHXl7z1o6v5LCm/CQnKEAkLIwleNnHUNqF
hWjkwmwXz7ZMs93pFHNEPwve73opDamOxBTTAi1zN6Ak5d+yQP/KZZq6Oc8IJ8KT
vZrTnBlQL0Ji0bfEJrewl5obsh6W9mYef8mGsB3ncqbhh1aF6nhG9yt/nA9VI4Zm
QRnJxk3L7viiOVkz0fJcxMwi5Iq7SgN9rHAOdbV6XPvpDdLBwq8pgCILAVA1Tihp
qG8IftFqVA28KY7pZ4P0WrvfeiotWk7ytmZrUaQXFTTLw1SmYie5QX9d3V+c3HVE
CSBlfQ6TYiVuBP1OkUn21pFciEcTuYV12AZEWH/qCOc2BXQTWr4Tli12vN+szOON
8mpuDeepXa7CgaEaT9BM2qpcNbDpyKUU/GhjSNdq5wrYwx679r7mdH53lUnOLAPa
2aqY5wEx2EzZqzFDc+8q/LZ9OgvrUC7LSDCMN61a9PyuE/IKXgUUAXAxHd/XcG7R
sInBYPX4Hf/ck5bhQpE6gNR6Y3uyEWbuDcz20kxsHO7du8a+sXap7tR4eQ8QU8AF
rma3dmdQAIVO41lQ65EWYi1JraYAK7VpHszEBvb4MsA6ZWYpFCY/h6kXuH2iSyp9
cfI38PdDvJjgIm9Ucj+AqNenqxgriBh4E4bQaTzW6u1LobhwRlHVK0gPEVc/EIZU
rLN9xDssdnkmDewBI5V5Zg==
`protect END_PROTECTED
