`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Pay+Sb+ZYNYrLXrNL+hjgWObdeIp8SOqLPC84BoQRNOwRyU/O9RKggH5oBR2nro
WamX2ttq720PoYHfJblgvvW2UHFxLW5/uc1+2K2SZs2TdSV/SYDc/26UijXzdjoE
AB8agraCTBtj5edVfHS7Q7mne3rLf6C+C/bW5ecVHQ0dA293EoFPx798aty1d1uh
qHCzYPlkINgA/FBjSnq2OgxJcV6g7Np+lU+yR58m+/Du7DFJnGR5qx0H4huPX2P0
gi/Eq2n1WnMUxB1G3R3su4uCvok8PH1gMtTgdb2W4Y/eNHWFST1pYnzUjCezBCZ1
jELecbpYMs+z+SOSwWvL0aCTWgTwIYLX112vsTMqtCSZjyvWqptxaeKLHiOTwD9x
5PQMTzSoU1CAbm6HsDWjI3uADwwozbbuEZLbqQpl3XrTx2MuPqHnAkrm+lRnB4Et
87ELrV29+7FLkKa5xYM8eXrSZFjgpe8UqGEe/Q1Jwss+mB8XbcNpEgzks5niK140
yeL7Xu4Ju9iwglF8u49oVdz/zh2qZSoOcttZ9LozFk+ga/so0NhTa2h5vghTA2c1
CVJw7OFfKpTihVyeXX4MMOP6xo2vmoCh//01wtNDo/G5AxD/Ce6WmOf6G43Tstdg
f5LKyFTN2f/q+vLtgxCxxPSrwshD1gaAWScRg0E37AHbysu0p7TSBdk7npk/hsQM
NY8sjI+5dtg5SAUqLX0q8U5fgnhx9j9MjANkcvOIOG5Wen+9g5SA/zCgrblxlacS
WhB/8460K6/kYW+AjschbNeOMUwC71Y0VM/gI1bthAeD/UPisUPxEURvZduGmnea
vZisgAh3HQa6Rjfrif8azYhsAmVVquV0b4IbhQlT08EJusvq1j0Mfsibv6kvG3TS
dBnw6gu5GMkmVVQngPVpVNBRAz3P8Si4NZ6SzuAye8qosbl/oljSes56K6U5BoHv
GJoLPuma94gw7Yrec+dStXTvUwagyjL4bT+UHu8jp/13We9L+nRRr/AtTaXumTW8
h4+oaa1/0nHU392NTKhW14fZJipbTgIpfTroNkkmRxJ5D/NsHZtBhoUAPhvi4IvT
zoFCvUW+WE5JNj6w1At1slDJNUtWxJqxAjdpZYy1ctVkbSTM9kg92cc9WsQ8tI4a
pa5jiYDWKS+RIiyuhEL6hDXC4zO0KMu75S/SjYZtkJT6g0mtf/Vjjn6kIRSY2Lmp
/IHWsnvwpieAITHopN1aDn7BLG66vt26In6Rh1eNfLTIBqmo+evnmu2gZ6QiFd46
dY6m3KYrzfrKWNdvdnxTinlpExclm5z13RQJGRNVHNulBlYHAAKQ39m7tphioGjH
zP4PHRoVPNv0PTi5d+v/ads+CypLiGjuxDs5syLsxmPOv4dDk7TiTw9Tk7u/RJAp
tIyLhuLOLO1bnX8JX9xBL3XiMDal6G2TJVBN3u9VWhRBqlxlzuLYmhvZZOHsf4TF
uno5zoPIHHHt1h0iaX3OOGkhKpeDF5mRfgrkYYCAwwl1klDr3bzs8AxExsZBtzRf
Ox2cqbQiGXMZKYY6yj73N8v3F5ITAPou2nBrOpJsyczfdWCcKh31jt5wtDpw4qTQ
pZqCcEBBD6n61WJ9a8C38J17qpMdMAZZcGtrcfy70GjZDjGf6mrpqfTC7+jBR7F/
mG3s2ZlBQgRL02lGIizHRw8sBc6mKeOih07dZXwT/EomxrZI+wsJR5ktcvD+W9ud
m/+GHWr7Szr0LUW53Ffefl2W3Lkm9BpUc63LfeQrWp2DNzPTrlBDKwwVrwCWnQ0L
d09Efur2NnoXwanulPr+g036whnKVTQ23leXXxC9PhZiFmD6zeS+SQrxyEF2RdFz
b6RDdIwjkmlEQHPx/zEgTUuTBVu/BvSNvz5LX/f2F+xa/wPQkRvbPzy6km9mU9Fd
539a078oRIIh+i23fhFPH3Wf5VTX33gwev00yyfGNzzijcFszbB37nTiu2If6bl1
vDAVYyF4E8ZAI3UTYGup/RXCe/mlU/dS1Luh8zpCfLlctpHDSSH15oTz3qvrTlvU
KtpMtFHn0Ao+TOGD/si7GtZbtiSOt+car5JIrb5sQJHctJo8zekYhhpZnSBtBUnD
P40jebMEvX0wovBHdRVKck+HmU4Z6tayvoloc5ITPt5bf2dmCAaGgjJ3G+xIp4gc
tbhHwchNVuqjM9DkjuZ4NlWBPRLe2/pTsE6/mOqcHHLHBUwwB7DHpdawrZNmP0af
/0HQngWdBp+dydWUncFhWumEouzETCv6WFyEIdw45rPvTOQOyE9tjnXPaF8Dy3eF
brYNFUjOZKiUUAj8oh/zlyoYdJKk8ww2fNKUtip7UlYuL45lCAZoC+oM7JX3K9aT
e/CX6KQiGoEIU46phYRJ+WOcs2tHm0DRYehqLupgff6dpMLytaNUiK1cfDJsZrqh
RZxtay4+hrPwEJzmj9DAZYLOUg66vHGTtnTUlqMz1zdoTZ9lHqONldBoNfGD4dnC
I7I5SKXkWDI+K84/NhRli/3OKrzeqOSixJ+1Vz6SoO6KGve/X10ObELSXRkVxOL7
BFXqJX6gxLPP3/eSDTlW0Hp/fNBAPjrPBnKOXZ8i0MudPaLOtBW2SfbnIeihf8IV
A/Ge0/CLLr0iIbTdvkuVeOID5VzudG2Dvj2WZ9fI46h8ZZdtFbUkVcScEWA7mqiq
HKdv2PG0ADdY5Vw+fM/DDGkeWwZ+jWYsk3/vTpPnFGye4XFv2soXW2wA0m/yExLe
K9+dSUU60O+PwNFpGMi7yrENv89m8GHakuVy9S3NLQHmXU0Jznn8l6Lzj18p+b5p
asKSrZYCjL/814yRuWXTJMz5jFh+f4PzuoICEk78UYggGXNTxe0tPZPFZQgIAMDm
psgZgIc2juATdbUZtEUuytdVzZhyLwWA9PpD8zd1gmlTc4V2FvtejVnzas3TEtAF
CYocPrmdSXUmZwf7NbMem72YnemqC/mCbTJxQEK4gUx1laob8T4YH5L6lDzYca2k
DkN6GXxTU6rIwrw1X9i3bpmiN0opgybdkv7kiRyZar+SzEjzTWHAriQ1N8F0XTO+
hVpdiYcbgDQhAaJJECqYiMRGE1xUL1UgcVXCJmQfUWVkUGzA7TxcFKCzB9UfrFTt
PSzUPRYjo+6GCqXBQxy9pyrpVPBw4oQleNnSzjGauf3908KqcU+YO0tUNizErY9m
D8AeyiPSwxBSP86bLlpkbbqOeDaREjpDmS40JiXg9XdXRNb1n5eOuA2FfRfNzfc/
W4rkLQtYQrbRRBK0RuH+hALQFrSYRbJZk7Uh+DjO2jLI0Z3ckDfv3X0yb7myuw9q
sANGSV65cBFgZ2C/olgQPJlKu2SQSzKhYLd9Q1tmPTDCUPo/Pu6GBoyOLap7chmu
XLZdPAMNiMngBcbGRosej0v7lNDQ8Hmd3R2XsuTW+ZiEibsE4IHqfWYs/JSntd4U
C9Z+zEWkToh9dTabEncmP7XOt9CKUmj0Uz5e3UrxCIL4UPMTM1Ffx0aE//796Fym
eA2wwYEk1tgDJNh0++Fb531zFqLw+YSZAtY7vrKPiBM826c89p5QpcWoTX6cJp4P
W325T065RFar4F5hquPK1nFEhBDE1Ow+8AFbshj2Jiaw50P1AWa9uq8CFKUZDYvD
`protect END_PROTECTED
