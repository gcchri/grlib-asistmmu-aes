`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLj7NDYsxNOknGLyWRK6oIRhOYMrRGgJs2NJhSDhHhoHE6IAvmnSGtypGxE34EW6
ohRX+LykKZiuiSao1KkHx53rMN9rim1nH+cacwM1jSs+2oSoFH/nzpkyAqLGx45r
09crO+FmySa0q5O2um94D3Ur9AeLK1qKjtxB/Vv70se1Tjpaz/iBIZIX1ByJpb0d
T+SkSOsNoxMzfwdguYsN6jgHSyjEgxyfhfyEZvBpHVH8h/t3KNFE/TkyQwResgxt
iM/M0quoaFZoHSU1zgzhoKklPgwtGHrh9Iu7sZ8UW0+tD9m5K8jOJHBJ0ktFTajy
xyS9eAcrq/mDkhCLo+u93kBHAZn5WOxZOOe105BDhOxyz5h79GMQw4M9ACDWbCb7
EwgFVwxDjefZZHZ0l07tymp2wLoCg4ZK+zcpnlpAFp2G2hfrMFZcqko9HDT18Hac
ZP8CtkbOhr5sI/EvoSz+Gb5QeUsLbbp/uAatwJG2x4cpSLbxafgWFvRb3b/xHGpq
`protect END_PROTECTED
