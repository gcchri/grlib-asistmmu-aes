`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VH0zjeN+kgv8ry98iCu/xeQBmdxRKMt2lIppTUffAUDXtCRscWJlKvtxnBSnvfg
XqFmmM2rHK+TD1+vuOwK7/wDd2g/XryDZ+XkxX4SunJL1mRJaM8Q6iawO/+LUvAo
zRHBAp8yMZui01G6NDutTw+BwXW2pMQdKN1IS6o3eHzfDgWWX06HmvJRk4Ke6K3i
ZqCLa/JWmgNoDnhVIB0IxPruhFhilX12Q7CdVkJK8PuTWzFoMC5poLkcDiLLvVsA
lszgBvqfv4IRrx7hciaKWC49xJ5cIb0+rxyLe5iaWKNRsa75lkeVqj/oNwcP+gJE
d6xT2EvALFE6KvTGAQTtd6heDMH6Yd59wmYC3GmSSDaJ1u1oM/TIO+Rr83u/feJh
5Yh5enzSVKlUegyud4ZY9DF1r0At3jtTsv47vA4JVMs=
`protect END_PROTECTED
