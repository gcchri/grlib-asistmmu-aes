`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyDPAJQ3c1L+AjWhPo2HadcTAe6DZqLrF5NUU+wsHe0tkcUkfyJxntivMnx42sb0
cj6/TU+DrRjrHlUxC2IkmPlq+MgNziooGI2Hx6jHd5Sv2JwZ4BLdaJ61P/mh8fdT
bfoS6qDxacTgU6nlZoZo3TjP+VPTuRwK1HUPxfUIS6V/gt6PFKMYJsZj5WAQEcVr
S5NXDvLEXDtanKytcg4oFij0AP86TRpD49qPsWrekMGAr17/2NamxcCUGalRUVxJ
4RoUS6oMETmcKrDRkH9CqcZObApwhm09kJFDl27TCkIWZPUepJneCwR4zEemcg4z
ld9R+yFTI3o1PgStOMkJUmwrLgdTjYlR08QlFY/GA8P2Liw7y7pUqBTcli+c4I6O
vy9taeBbvgL3RD0tYvQVyzH64q4lerFeAV2zhMoQb4wYDQv64dr3u+sMs3cpKpvN
BI/5m7bHdCVsjPQr45sNoWen1jNDUhr5gvaDtr2YuF+6h/HKLcZREEKHMD/ptroM
XNP2824rq0DhnK2jvwYrHeZwHz306NXuxeGPeg2bGDYd6yTeNPTRk3piQKM2vNZC
DV0ZFcC5Zv6fqdLEdwkDYGutSEva1t7OqqVtZ8q8zteKFWzAJtr5+7Tig5QBOh6n
Nc56yG85FIFohmhvLfKuMxX3IzMGjOR0+eOKPM+ItA604EiKJQ/Uv6Teeib9E6WD
9Z9uvOEqXHXRP5Ar+CJ/FUvotWTrs6ewxLlMQ6pquDWUBJupGUXNWL+OQLTHfaDR
F+emwws0Tr+jACxhFKsQcrwdMq6YW84qtQRYkHap4r83OVmEBX2rvnn+vL22p9F5
7ZUgF4/v9PbVxtd1cS5SzSmfqEBogt715JfTTfgni/MlG4cBBDCCTytEZJehWWfF
KOKbZWuLRMyp/woxDzumod8s53QPskhDizs7tuFh1nzOa2JeBVPpZgH2JaR+kJ2z
oAyZDnr12j5e8NFP6FmWG0X9p4aHPHRWl370LMifTBW03AuPeZH9zhD2+QsQsJmp
g54DPr5EGlnexlcVYknc3JP3TcyXCf5h20eYK79QfdsDgcCZGWANF1DVHCNvYRih
mA9Rws8M/J/thGnlWaiEat4y2snxSizjZbssmv6Eo+PrITnL+gDt5PuZcTm4y/MP
URpNgmcw6WNjXDjRQAFuINzrAP5T6Cm8NQizHP2KyUP2ONoDzUGNPis6Xl6JTFob
BpjGa21aGbq+OEi51pN7b6rsOePYpILfB1dhiGn20IGPVayCsSSQFkmBnpaF2a6F
g2nE5wIMWFpZ8IWwwu0m64O+O1+WzXXLQdLluu64p1Rj9BzOgCPj5YzXoOwmx2lG
8gLlpSix3HWEg7ni2RQ9e+IgSo9OyzW37UcIY6YKAnejs7fOx4CtgQzNQ4bPLZqs
GlwU4mSjNA6TZxNyrBE05GK9CLvJ34gpxCrAQCvXOtYBDn49zoc5YQz2A9NhTat5
H8td/yphOpRScMWLC7wprU24HSN2vEERH/c3sij4A2EvqGAfpQmtqXb/VVrPRpwF
DXtIMGsgtCwhNP/wUV9PT3yG0vp885S+2GmCgj/o6hPwJ3sVOXsT4Asf7MOykRzy
G0v5AKztZ/uNyAsanxoo3jWkdsToqhn6GDCDvsw/WXJpy5dkOMOAj8pCLhbUki1m
CbKrzl0qb2yiKh2MniWHqum0tvc3uHHWy+LA3/jAVJIAgA1tScL3f9hwsyN2EXGn
Tip14ZKTAf2vqvgrgDs2M7ber0CfteeiJs2pzVWAJAxqdiRtoHmmvgOfFgV4b0IK
krBj3ezIlsIGIyRuh/JOMauqfI6ne6IYoOZjc6h+RxwI3J04uCvyd32iFSnAK3kV
8jMC2k9VH5lx+f2wg//4UWnrqa32HIwNUgF9Y69m3UbfqBz2JiFjtIhaoT9Uc7nx
APKetP7UK5tvGUXZ585cuKFu6bMhn+BP6lKN5hzrmwvf9zdf6Bb+IgeQqC3Ezyb7
3zMK0UUpzM1vkbNjSMQZE0vSu/QnjWTjtc0is0lno4tGpK9ZXZUroOdJtf8vCy4r
snfC0OcV09T3P2Qhm0z4YOgoNKhkkpyTjKlZMVmO2hWKdK1HkcRf8lVps1VUPqf4
2ts5qwotAYcyFJyutBt9t1/UAoXOu/++JlyY2FAHB3JUNkrJkpr/1di//MDKfYVo
9o2IR2cFCP7ty3+LwWc8x5ABxIgG2Wj2IX8OFlfNy1Zd5EpkqLzLlMS3ilFZHJZv
tADG6ICBACf6gQX0ipbslJ5SshpOP8RGcumwKEe2JosVbi/I/9ouwtt7/LEtAhTr
FeUBz8HSdJ2VKLA/OEsWLWk5qhmUENTMYpZS4wn+Egp7LTTDCnGeNdfOGR8aZNwh
JkR0weGhPvlIZCGoY2qqIGWdQ2F5y33zyzrC+ARgKqjpA90dazdZ0+j99U41l1ol
dBx5BzCm03h59B4LZAYQRI0LasjaEXbqswpT5pbRKWIXGgBWwD3kl3pKj827NKNJ
IYy5XEMKiddDr9nVe5f4XtbrYghIQJUPbV4FWWwCWgfN2XCi34E2d6d2pJPYbGhc
d5r3fPfSreuPefEjJCH9ltVuVeJ/1NSsCCFgjA3/ztwdo34gzCi2nuFlq29iV/Ld
LkcxfmOHhQFqvGB7jzkwNm3NqI2iIRTv+sQW7z2AHegx3zz/kNpWzaKZaPPdJKO2
bRytAaFfs/Unj/spP08dAxrLbKRp+IjlxcXGhusbzMX+zvnl+Ixz9O/Ug6JmKjvG
GC8s2trtDmsrg9q053mlLs+tz8jG0Fj17vSM8HqERrhAZ9Td7YEwcKhUshPumj7f
o0R3HUdm1LhWAWAO4ZMVrzx5bkZw+CzN1ar8FB/UQQwDBzbvR5ygk6ucW3ICH+TD
vGdYOvarH3u8f+LI48BEWLRyHHZQUlfmjxY+95m8qV3o2J2moQvMjt9rREJynmts
tEPOHtv9M+sfqOh1QQihNs481eNmw565S79fQDEWxeJxlxzslMRPSNp7UkTwYR7w
ojFW/tkqOl2p220JEB7Ucxq+k/jkV4tAELkwi4g/wteNoN45AqXbBDaVGvhkAURq
VWbj+BC6niNdK8slzx2a4pvXlo7JGo2a+/TpSgFXu6xosxE+SdjnGvlY6Cj8Frc9
/5oJaU+5xcRA4/BorgAYn3iKPi7hXdO5W6M9yTe8HBcUPW2us/Urn9CchyOXCyxx
VQDusBssn9ZURImkgHu3IcGWE4qYaE8GjG3tGCUdG3kI2316lySsKLfR4aSek9se
nn8Kj0o/mxTN06SnEgAmz8+c3rtCZKJXc++zCk03sdHm016Fz0Z5x/NzY2bGpkwV
5ajNzYNWHAXb3EWmQGH7HNRrgU2ZQHL/erMO3z++nHIWRHmYupB3EpEhgSJQs8/1
Gz5EaohBjAGjMIRT/sa46saJ2rG0WWAtnPWfla5yz8giIgNxjLbMeKuV/Y/A70ku
+I/2qId41YVc6rxrpMDX+saVGyfZyA+nk42vvL6W64koRv6fKV8VvfGooiNXancl
1jaObALacRjGeyQrSQN3xLID6sDKibZkpuYLtC8aoBf7HfG9w6+dcNG2tyUXhkm2
TA99mju2VOvr9/QmB1jmC7ez2dMF/G0Fkl3QY1/X2rHlYl+v11Pzvs5GdVeqOeEB
koN/ZxQZOwvwQiM+jRbYhCuLWO8Hhbd3am/pdwwS0tDq4H+xsfXnUma8mq2GarEu
nOoYVopyjpqL/mPbqN+/g+vL2LhQXaObgdCkL+nA14JIgmyICQ4WFyww9fV8E6/b
9+B4wp2/s6ldyrtXdNzhOqqarpBJgQ6sQXNaHs3QfQ7Vgqjsm/TBezhr7bsl/nYd
qPGKaXo0IZ+ogCNiB3R/5H4tutt2Kc3HXYlZfEu0V3xlJ9atsvkrNKLj4k0mB654
kWR+3pRwnvpdyT4C7V3EjstLt3LB/lzddcuTjhYkTXqX/9hCuy1ghm4O7qRKURvw
YtpotSzS8PMVZIS+bBXqMjmKsxD/Qn0y9xPnWo2hR1K2lrd8fSJ0bIDgy2GiIkSZ
JChdtKT8Kai/dFYrT/H6OA1MM0ZUelIkXcLqlPDsb2nKUzQ/AIVnIfkft68hs+j3
pqGt5ACkCtjX1BMWol/F/iv75sJAXcRKWV5QZZHZztl2q5lpE6KZ+IT9b0H/tQ4J
pf8hanBiy6GsrTGI27GC1eq8PqMq3apQ9xQVGzL94zbJPOrF3B2LLVIGFoOgEDaW
L9qesHSVFaXAvpK4owBLUsc+JKlz3GH3hrL/WvyQ8YdK6F4sKttyJsAe8zmk6TIe
USD9yv2dSTfh1gPOK/wzosLwOUM+vgGsAt3ltFAuTyCAq933l338zUKxkPnMFOm7
weKtx/gFk0xGmwV45Vobji3edZ2QEqunSTRegg5qBlG+/1MAYv96X+/zxx1jRyMc
atrdsxlQ3Cjh7eWnS+1VXTmcRrFU0KlRZziMkcbd4cylXcfbtuH93hDugzSIIIM8
5abZbd7vgu6rKYx9EKHFZZtO/G3bFUdXvz7L3mnGJFMVg/QEYFINQU3yXMk7RT9R
nry3HDloyGmJ3RHwKzxzn/r5SQhvN+osNuBodp3YIqWeOWO4s725Hz60FbBfcfXw
0ZLv+Z4wQNgCRA60LL0YEgnCwJctWLyb5+6A30zvd58zKtN8RDj/uDWzRUWMpyr0
V7zpq4paJb6ZDFZ+23QECVT+vAue1wDGrxxe6ihV3V11wVdtyHG9z65v7LRFMKVJ
swQI4An4aB0GaRkwkj4+QNDmyv8aIFAAev4qYtRICAdJMTLvsr0FGm8rJEtgqWxN
be1aacGVrWw2aYRIIq5ZbCxEsffqe/yAvJDtHCZ26mFJl+/+xADSopbaAqreXaqP
2rAiAK6eOPJ3rnFyMSrDsYUl3vy+A2IRvvBLqbQC/wPgVG+S3Dwae5+BLBZYhvCg
OrbgXe46Wn+23uxGHpjskM6RX8EpBTY6D//5RI3qGBoV3wExxt4avBQd5BKqIAju
4iwbjhJDpLVwBfGUiPtjr7+cQ4M5cTEqWbODZ+EuECpY1jIKTYtXVwXJNrIp643a
9tKtpBKHdUzknJswz23Yoja6rmcYqmmblP62R/6f3PgivXpi8gYKzCCrg/8tM6mL
5pAfMyrWVVNcqgB0buVp3OpfCE3Lzh4J0kwVIt6lKPDxdfL3aBRWVXYOhkfuNdwc
42o4Na3YWjqiNZKnckezt20KBthUN5BtWfcMDuPMFvo3+KgyFUirEnJhEztZlf8H
xWcdFMLKQK55oFOLN48A6wfEO9FXAenU+zq0V5WfLivg6rxyGwpVa77s0crsN3N5
Pq054/dCt+/ezSyF6JUAPlES68MNU4VUlS+O02utLwur9o0Axeegw8DfA5E4RK9s
e0EZrXg8Mc+Ws61L+v5hCUt1lHPKM+vjNX5563d8pefPymQpn/7KeeFJpS9Fg7tf
mwf5os+ABx9v4B5mVOfdj6kb+MMLQKBciYzizczp1BsTruT8WLfrUOsBGHi9zxGB
hjP6byyC3YVbpzhv3bA1IjoTlwGkjd2wKT6a+4HSQxmTieQnNy7vi3f4S8UG+9W7
agHJST2366hoQK3bB6EZK+/emTEQjRn3y5vFc9Y38BBHCBiciA5jbwa9Tau8pyLw
T35Ke6uVCMbj/Vx5EYl7cRfCK4vOZ4rEksOyrRdybr5KMz3xDGWoPt9DA8isPKvL
i+X4ua/n77stgmgK+Rb3nROGy/VIPz35qHOoB4zdVOWEmijzSSXanFG7fX8tT9iY
RWlgbjjUg4Y4QK4byjENl/RyEDuOsppHLRu4769rXKFEwFerfFqvCVp/SDw5UePo
3C1422r/ny5rEHppLtSxfTQMkb2gL4kviVIQBM2GKWYAp5ZiumAdsSgxWrVMLzrm
6UNaG7XHlEv9DvzSqN6N+SFzdNIqVG2qiGmudZHiO1iNQZp7ueb6pzOUE4vrhMXd
2iSlGBdqHKTlzRjEysBTHEpb1BZB0+E9YkfbTIdqQedMMzOoynZ7ICjk2ctCalH7
8iTycDPi0mF1zeiUa5q7J4n9gc/J3KLdsF6wZgXL1s7dCH89OIthoje/1Z5fIOc3
8ahlWoOcEMxNbKvvAM20u50s4uREaHfOCs20g2Pg3mBZX5ANyRTnq8KLXvJYyFe2
Cu7RZusEyOx/wttYt/NfiyVKbvgspRx+JuGx0lt6YHmKFubrgMuI+rfRxTjerFk2
t86j2dBsyjQCc8/ckIlEc5lvYx3qI6wu9/xl4bq+3sOERYTGhFbOuTE4GZKP4lIH
oR0wXBgXFj7kh0E4sFEuAu9Wt3PZb84Uxq8h2QIYt3Z0fzcJONPpgFYz73Rb11mk
ZI51PA6ZJR1EGbhvyGq3fFEeU/wjIeKxqLG4TU+ByNX1MEkL1N45fcWfmR7mzHkD
2u2+LDDSXaFW0tQtYGoi6ba4+3r4CqOX9J58ehUTjj18TsPixKWCnymiufsnfiV2
APDqSK4gDd4VFAga/8I6IAjPA5XFH80waCIlGvFtejBLpN4pRutbWprACDU2t6Fz
eJXzrCB24hDADvLJHJPGAet9eKGLxBmtEmkkgXMmMYeL54+A9W9THRgjOXb1BlBR
K0p1KcHL4XPz2DhP+kHdovRibFiGsx9biFZSbuIPakhxh7m3iKwSHPi4Wp+Eaz9i
F7JPCjbb7z3vFQeb4AJSH9HdxKW62tNoGWnmycrMMXBdsMWqJkZXDzdvgw/LHMiB
TkBihIVvvovkxMtDm3csWFGzJlaEM018t9PJIAgWNd2yjvLM/Q+E9M6xkHzMG8+1
XxF5nPWAEcdNCRACUzr8kTOyi3VxZrPfh2Xf4y2v6mzSC1rjiWf3gUc2Il8zWDDz
Eeqk5/U0iKYjpn9q4lNhyVrX8KcY6PQTPARECPDUJCP8Qboutuz/rY6xK8cymMod
z+EHW64tBGpTFTOMIeKOpfyN/uWGHZFXebCayNV243C8jM2eFgx88c2Ut1+CZQlV
DTU3nP7Xrvua4pR1s5sj3R+0W/+2PIxhi+DZuct4b/DLi+WW7Oqz0FMflQ5dzPqM
4Hmrd7DG4znPu24yxsq9NxZegiAAKPbBtuJ6C7lrccDCS1nUEgqpEsGXFDNVTu5W
otVEAa7M0HH45eJvYNuab/3uf0r7Sh8InIkaXDJyuIWEsG/sqYdzzgFRlp8B0jT+
hIKWrnHmFDMxps5vPtU/8I4TonzufmXhopACgOE/H3K++sMGXEMMBg1aDCBvv2yw
0/h3T5OxtTULOHeiDhiazpU6bTnSL20e97r357iamwRLKNkEyBgbw114sxCqqgqU
t4tpa3rGBkkTu6Laom+M592rAb3Rapgo9Rb5rDXbM/S7kSaAUX/TorSC3rR5a1u9
zWMCPIvua7bYaU+xtdKKc7+F3vmkLg9365G1kgq+G5WP9SOQJZ7rUG9uxcGfkOK8
7h6a6flilwX5QDfL6wBlHhnIEYTyDn4jT+wFEoLCPviCA+JUXC8EA3Q3BUp9deF8
I1hYasdyBQ7wOrMVZyp7RKrG/8tPAdKNmV15UMaa0AseAR2dfBW8fRZLR4Ed+kEO
1miQciRH3+A0eKmkJ1nNukKgcLpGSbtgbZU3hr+a6YHZZEYXwZZ+zBMS6NGmgycD
EYWiSnyJKQTOvgNgt5b1YA+CxkcwbtZ0zFt2hGdnoZUAX/yzyCbUNtxc+YOXsRAW
RmIPyvf659kRC7sVqqPvKO8uPJ82sq5ZaG8wlX4JwLQA6NKvbmceLCtlT5eEV4fl
WM32ixJM+pMUrjodkXhz1gsWa/Jn3uFbGP07CxAvIJYlcZLJz12YII1Rr225kK/S
Byi/QIxROizYo4znYdrfOnjL+iPdi/u9mOXgdcXnF8C4qSpBNJg/9GIvf5xJiKpF
mg3pXOIUN/efMsrfjWNTRR1isfuVb6oRWGlaM3T59pd77WLEqGzDo6eJ2tYhfijQ
5/f3LBQUssG+lKYZmGJYNdYPa+JwB6/uUtE+FbB1WNODh3Q1DlaPeRrbTWF9FXpu
1Wdv2pO78qPh/9/ac2mAhyP/2+O/8wV9km75t+36xJOa70ON4fZ2/TCG2G8hIMG7
0RTqgGGz3jstiNFHOo/HKNJvrH+6WvN2/vDDwoATYRUsFdodcqaYX0EjliLx8pBa
MBVDOeBR8t3gCnxRhBwDia8a1bbQCp2Qa5xjAV8p6nRYLIUQQUSjKjODA7lGH9Rs
Vgx5w2QrCnIX+CqJEZUwzQvdvAkObS6Xtp6e8QUoojcndRNsNrHXJjvSYVuXUsc8
7dCM2Gijmb4jarEFwh+AdhHrVRMoucIFxCYSLYPurG8sZM4UQxNpHqLqE/LMY9K+
mgPEFqd8XmngBR4Ooh8Bx3FhB/0MeB88pfnNt0WuY2+nRA0SxYONGE0DXxfVPlJa
Vrv/JjfZ994Qfyrzglt+N0jQVIvQ4BAoHO7MaNhN765Fa4PhvyCFL854hjkmBHKN
R7GZSCVolMsN+UnkLXgAlVapWTxTHbI2sjc7CQLdooC5gNQV9FKtAXA54vcIXi9y
Tre5kui7Nf5T/xWRLc90KRqA8tJ7EzVkDFagypBPVHFU7pr8JyS/Z7GjyzOD6F/y
46ZYoNc0rV7ZJ3TJOdpIlIFPRnYViCS1erW0l1zsypgbuZCmQGIi+w2PrNlQMw8H
2Ie9KLf9JOT1xpXOdQiTXF7mupeDKlVlnhNC6X+luWu9MZQJZj7+AWeoOtd64awU
aUp7RodoQ5OYKj6mSGmJu93EluWc5EH3YLKU/gCo7ZPDidH4+9x3hRyzArkjYmIS
iWAERzxIfU3CfMeJntdLSepLU8hwKZuNuUxu2l6I9P3OHyEmLzVKDJoD1mkMEOKC
1Y2u2764ItaTSRwn0LEFSRMEMZvWpdaThlG9YyFAVhjcy45y4+YW1Wo4AeY5gspK
daAx3/YUuktUzhiKc6ROucwmommhs99IsBH+VUckdf5O0ZBrSF1kPCfo5i0679+c
lMrQtwdtsZ42dGVIraWfqqookgBgkQFwTOVRg9Tg75AZcIr4h3g1DOL14wlhnQxc
mP71YGmhzTJnjPk+WZvQSngFVNk461AKHNCcyHU1Ei90VNZRxZhwBoAZfHAupIr6
JtVSWQgCEHeDE2787DW39gVGmcGk7TkW4w/V6Sb1FHSKX5JyWMbVAdvLXsrNHVsW
6A8EFNc2wnP+W0JxpbpI2j8GN4/tDHEo0YTLpODUzifw7EeNOlFQpIgNqVaPxY4x
lNkGTIsgd1t4107jhsPgNFicIh1Sr0ksf+KsZZeRxpkAMh19ht8T4UQ/GykiEQYs
PmLVgODK3q9A1rjidCGT3UjnDkOGEshKEs1BIea8dhMYYnjnX65b9/KDud9wuXG2
r0EY6RnQcIU96+x9nZ0ctR1Q88p+A3iE/SY/IKOEoNEwxTpe6OTyvMqUwpp6D0XC
bUHn8qXFd6icnmEuMBKvaATLTPcCOKuJaolWfk2THiRoKB/AxryaU+FD1B0c4z30
BW/kNxoHXeNvt4cqfott0T4IyzJO5S/WxuW7vyd/JjzDUIiUlN2HF5byw/qGRys9
jucDMP/FyAvEw6nL0WL4wj0xa8faTjo0SsiIF13kp6qIXOAYF7DcgtlFAm1aP7EC
jo8Y0TctMrPgC4gKmRovHa+gCErvMFGF/AGnNjk+4qXPP/7/9alWAfDnUjfCE1mW
QqWH0c7xP1YcbevhOgiX4inKV+i3bkwm42tnFTvKRa0v28wGVj5mwGlUU4pgPlQh
cQyE/PLWD40B0/2JuK0rqRIhPE7iNBXxgWVtOzae6iKVCFFbd6SlcMa1yAGkRHYt
S0MxxuDq8ma/5gcSGMnBPKHACd1ZPU8y7S2ZwuBYsTXAspBkTpuZpqAPu8WfsAjE
XD5ZCCqPdJBO8oBM1HLDxxnod0bkGrBA+0E9V/9cwBBMBK2ckik+/uMyJZ+B1afk
NJAYAuLZXnXJZprX1x5ATrB3rJXFTLzXRjV0T8ThvyX8i5tiOsektc5LwnnJ4OuQ
anFHjdkDQB+46INt6kLRfHSdKZuyt26oV67EZZKNs3qlfLRgqQz7X7fqC7d3kE0B
HjNpHnGM3Rd8sCrRJaqcd/H6ztqslBs13kynT527FJL3nhrasFXSLaKtI9YfwaSH
pXlLQgPKO9b0aSCJuOh7/XouuF5Xqm+yucIxUdqG5n2zWO40oxPvF4imeKPvNtJ7
QiS9D4I4sZZMgRMaIyGYPDL1SH1LiQphp+76cvnyQz2L1S73C2eYOKHTBd/Ap4I5
2EIoeToI+QbRqyu4HLIZ89AsLhKrls/jmWwHbEEbi2Lmhg479XEoJDCi8fn/rnwx
xItlODgVAQvax8y1TPB4o4IsX/TwX50/Jn/skMp9nZM6OpDPZFYOVk5cBrqcHc3r
qI5B+Qs9DFBb+yNgNnmxi8hJwx/xgZ7snW7rxLEuFJKa0fPSXHCVpCrU4fhsfImY
htubt6mw/tDi44hmhabH62Gtr4MHuPM/T4xyZ+qLZv+Y3dOEe0bzsb9qZTM5z2Kn
wTcHs3t7i/YNtPcxsJ5aSIk44hE9Tun8e0/i1aPmXVTWk8TXqP0lwxKdmPg+Z366
3BlDjHqkTQuXOntPixhXrcGW1JLwFuTFNvDkQyY5IA7IYlTh1HgIE5OBgQuO57JA
ri2bmllwcOaR1WNEoodUiI2WgmkgrklGM96adfQUDlsqWhUiuKRGIrxwkmnP8sEW
dsH14EnNqClLQa5+sAnaSxgFh7ihupylheq1fIYBSSUmTXZ4yIBb23868qqUUtiJ
3yC1pKZx7lJhumKc6zENc8u43W0X9mO5ESRoYcthiq2O2neBHAj4suc5Qx49wHs/
q8+KPXWlki+1jIz/m3zCRxvAB2+u081zW88WNu8pDaoltEdgJl5rCGT69rBf+nWe
zft126lFRaraQAZcjaSXcK8UwWseJYpAbc6Kdf+SEwLNEmxb6YrZZyLx3ie3o7Ee
N4o41nc8jSQDfHSHWa2pRuu62s237boI2GokCLbCNDom6M5c4KJj8cxcsfg7VaW2
QOTtgWwq8/y1LhFCpe++0CUiS6Pv4SwmUW4xM1ZynYCnbCT+TNAqE12P8w5qqQvS
0uYOqh3ZQJ12YncR63WOdNqACZAdxVun0ehYVnHNhXu7Newbtae1dVYJWvjZNVgJ
vnJzJfirqwkp9JsQvbgaGM3ogTu1NxYRTyawD/VBOUf0betFYIpSjRyaX41dyQu1
qq9W0Og2NxBh55gND1V4jCwXcuCOtiV7q+uBzllz0+j+neqIs/mE/wHOvtfNShEZ
4FHUDRH9zrkZj/kSatM+hO4A0Xbgui69KafHxuoKjopY4J3bhS1oe0JW9rUOWjZH
1AxrbHBU10Q/e5LBKyfnyQd2a3AegeLbRseRVZDUbdtgLPsUNGuOos2+rjdObHkz
j1r+nmyzABj+KG8N6z+159fxRrybZSSDQmiMthZBVHcXwWSMUw+Nqk5b6JP/Z7SH
Ejso2U2Eozr59ykAZDOHz6ItXBdTD1D3EzWvfVqySPGU7L5k8U18Cej70O3ifDEn
9yZJIjaDFv2GcZ0STfxbMEbleToBwYITfbZDebfRasYcVnzEcjCVlwMu7vLuzzG0
RmetDTvkwAqSBePxS8X/OcNn5qRtT14zboLJlAvYYuKlX35XZNxEfeDNsWL9uono
/DJKGMzs+YCDy+ChabnWlVLrtreCnyC8VkfVqgzxd7Et4yxo1APNJSiwI76qWDAS
rSNZt4j06nDuhgGsUnSjgBimTKTl+JnnddRJ7CDcQIpjQb/Xxz1Y1Y3tYTZjm7MR
X0WZNCULuCxCVuOdx0ZDC1mQt1HWUTPyTJlAU99UqSkYPusRXnlIgOEt1vAQIt7l
38ePgGyiVRe+kChQJFlUOZnbT/YWec57/gqxo4D8OFxn9O3mQU36pQJhRfFWQlAW
YNx0No5lWLEtBApOu2h/S7JS4KQk95fDxTQB10i6pVNK4JOlGPjD3a0KQ59OlNWf
GRFwzC8spkLWLTaLpb679tnRL/iMqAaI+4ExlPMGGM90joKbc8v6InDmk6Svdftc
A1NHnOEs81WYQGEc0CPaK0vTTdrFMm3UiMw5GEB4lQL+S6RmGKQ6QgzcjBvoDqlA
Y1MBSk28KO8HJbUcfsPyKmwl27j/rLM1cEGkmifwDUwbCmUn7nTsWA+3MMa3spzI
6evVhcVJrS5791kvhleie+ce37paNaXEHfHDpgp72Jqep2HRhiJU6sZUz/pugX/s
ZOB7DKiPQZcM826k/AuBRfJTI9Z5Ho0dgXlna8DBUX39/7/jh4pHlLLOHnUjE42R
VV4F54Ok0SfnT/G3bj4+brkOWgd78zaWpN9qYMcNRpXgVfgErmK3nAfQZdBZ72Os
SdBJeM2Mw+lnj5d/Iyb54ZjxebExrCHoJ32/Kij78YS2Pr8x6MRl5yOeecQe+4RN
vN8IM3oguCSbjJ8RgKL4xuvAR+cUfKjak+3hqipYRLunI6VB9N+6hOcAP60YC5dD
cT6S3OiVJz3a6P/WXln64szlIyF7uDAK97lf6eHqLsrTWPsot7pWknJLW0MiNAfg
QzEIuRSEHEWieF6K6HGtrwFjY9Jjm3wrBHmbUbmTMCSNQZ5Fu0yDY+dGInQ1fI+J
gxrAXUC0SM+g18Lf8K6u6Dooh2Eh/slg6HdkC0J7JJSBjbIxHWJPQzwM4fa4ecxY
BgJTUbmcOxT15Bp1+hiuLL+Tc8utyhyWYLg0/7YfcFQi7faBj13LwOiY8vdxYnpt
oq6nBJv2t3VMAJqtMSbq2jwsn2nQ2RDTQRh8n8u+Y2yKCqCtmsTAz/7uBxGlBXvw
efBAvkRQq88N5BvQVAGV6wQCMSv5wddFuBrDNM5bNnkFASpOoSBVeO32z8Er0w5S
Q9dqqSlyqdk/27dIY3x/6Dr05gQZIz6sIGAPPguYvUGhhX5Blap/1nWp+3WAmaOo
dYs2fG6dOmzoh09s6EECIZeBRUYwgHRCxI22tosg+9qnDK83qKEtDXYDVMN8X8Ws
xpJdaYW2TeLAzwdo1E4lju7H/R68WgBU8mYTF1JfoACaM/gwjDCU8jtUr7NRGSGm
/RSnlxeaV6zuOXXZ7AZoHbR4QO2j3KEEfaAvpI626A5gMyHfetoHqxpL6XpTZEFc
r5Ctg/gXJIphC3KCOhWHsHkPFuf6mRZVgYU6/KaCsE3TzXwFqPhofdhF60HVdaSp
njjN8xR3DDHxlapixjw6FQKq2ql11m/uhn2FRjIDBE+5daFJFXycMTp4tbyAANS7
gNqDOy2FKeUWCZ+XsssPIs4MOB9Q6mLa0GjDnwI7cP83YBFokneHvDpDVzcTOr5G
kRP8g5A3MslZF5IJavQ2kT6Twz7dxvdKoYu5yhhBeJfCrrnpg+vyerInEoo9NsW8
zjkX7fIjKDCA1XNEeUT8Yz7A/kFhRHgnOzfGgQEiivgNw7MommezgMD+ZrcMnUHR
k1KsJcyYy6gvkQveXao6Kc9HW5J8J2lpe7hKCrbt2yYhg7bQqDKOeikSmNrU10gL
tleUQrxKr0qv9qvPZNwkYz8d8OgNNUZQvKP9/5cXDCrWfRKrlVBbBwQLUQS4lCx9
+wA3egmxzhAT9IHHH7GCZMfyV9AU5TRdUxr3+b7mTPeCH7NaHg/NspvfltAth3wa
qx/a6FRPZij3X0O6I5G76CuQi7G9xvuXVykLKXHm9Al83xNULW+3zx35oPhRKZaG
V8SVFjEUR3t3yz2Urx8S/GmCfgVPtN3XODVvogTGFdpqWFWjs3mmSv31rl3Jl0c9
jy1mcic1J5ljalm7GO3hf8wfuU+uZbnFtaLcuSNodaNSF4/QiZDhWN8PXiOSHbxI
5yV7zBaG35yJIfLi7K10mIT1VBv6GVhO/IRhiCUhA25tlTkoVKbY3Nml3M7iKvBd
gTHKwpp4mgK6CDJI92+X2cyYi2AftK+wcm8CpgjkfEkRmbTncLv0/NgOhay3vPBR
8ThIkRU+ghni7DZqvIhnugwRhDyCLivqmhoGlOQHU5Y9ktEDmIYFnYEwNuNvEVyg
JHJ9xHucojyA+Y3roPishbVdqwgh8HhiwtD2egbYTk91kqLXK6sn7ntfUsE30Arp
eNoe4akt79wsBRSnk3SvaOKUjenVI6/p/o4AP9p0Yb6OgJmdr6yi/vzQ+U5EoOJs
mkPlhf4L4p6lbKnt6eyQRcSaM6l9ohzc2KiupdR36biC+5vvkfxdVwY+Hj4v6hKq
8ExTZw0L78gnoAYqYHS9qzGN7qF0102H3NTLRO0SKG7u4UVkuWMpIE6nvHU4UU3T
fnybZTQMV/9U5UcclG3P5UG+46oQ1lI0LlN+wO+9KadM39v7KRtLYqe1NZyBpIZd
9GrhW8krU18RjoFL7JQrzCH9DAAKwGPC0rpUMG4MxvP2zgaH9LrH8y2mS1P1xCO8
WJFrMXNT2B0ArkDQgk8iUmBeZVNA4lpqApyR/UJ4Pa5lxNavn8JLdsZxNPOD6Fuw
2vHEDeD8A3zE9jfi5SrDuoOdT9Hyy4oBqGXmogKM/RjRx+5eMad9pyXijhgc69K5
BkuwRpg0e5DSvkr0QretRRW2cbdE1vUf9Ye9SMu2mnUimT7iZ32fWo6QGxo6TIdm
hP20OAAkzTxSVrrjATxZz42ds69kxdSOnAN3Jh3tD/DLa8BG6PGWo48RdCh6cqnl
cF8jue5Dv/ygUoBSJvjJW4xioyk1Pp6f49+4RLfi4PH9DDJ2ypDJ5iD5LSpw1cYW
++ieM0J3ZfgovhtCxB/PUZ2RRbsTjYaVDihkEH1stkzAg5YuOrHp3U3bQK8Mcexn
gFpTBU9WGhLd33wZ7iKp9/zDMwQDCiywphWsQ8kZP+on8mBqBWQXTAUvxkN4MgLC
BGX95LBARRdc9JzKMXPagIDOo5+QEluaVoKqvVIAeGMxIdeaB8ciMkGAkOGQMKbq
gpXo4mI28pweVhRai9msv1YIbufR9nvnmDxiNRpMIW4baKQjvD4iU03hfcxoBXxD
R3SigXtoiDhnKWE1YSKJoF67D7LA3J2oLcVgT5zWbaEMbXhM+wVGIBVdCxsPRx8D
KTpc36GOsaEixmZsl+yAnweCMpGQ6/iBitPGxWwD13oq1d7sqMuuNzhjNYT7BPGM
amUeqGBCQ1JdOW6PWGNTLxCGLpnFC4pEY0W4t0VdReF6ZxI2NHFG4u358acAs06a
VC8cB8GVXraiLk7T3I6jX3OcA5VG63cw08ZANyHHk56uXaG3rPMy4IDAzVgCWSi4
9e3RZMZ/kR59mb5/6RPgrNf1w+ILWflCnGLKnerdZTDLABcFJHKZdaaKwDo+KIdd
qlF4riV3fkxZ2psn52r99xUuNwAA40dHAhUtEc2nkLYNp0X2KPXeVGsHbiP7maIB
ZmQw2yeJk9MI1h2N3GhsmeuGkCPb6CE+NJKWnUZr7LMZIIepgTThNuM94MbzPZdD
lQa1xPBfheDiq/UalcIIvFM/hoicryGfrqQj2Gqc+VQGE0MxoQp73j9dxWunFZ5l
AdrMX3Chgb1zNMt7T2w+cKpa93JBbqzPTA5NgD7DsbKV0GlijhsGLTxSU8lZMM67
FNOanyoA5uFbf5oE6eG+tkY8HhWSaLC9jtODxEYNYBUW8R9KB1Hgx4PWEBjmNlKA
IrYDdyer0JvPRkBrFBBonhmZ4Gzu+zVjJTpv/RoynRTwacJQx2uP0m2oXgIk0tBV
wQzPpOVZTy1zoZyVmJjAbCLtAcFSZfnkiYiKKBRI5f1foVKW3dIIeI77/qMS3nUg
su4lTBGygTc2umCEce2eFE0NFrvG9Q4ySz6MkqbdXkyOdIv5G+cuqZlsYzhbJgUs
0Lp9Xj6uD/ILNWo5itSVvCrrleHbh/aWKPHbJo7fpMgNfgmMoZf/fyQ4+55EUwUW
XoWC4uCmcfJPf9iemVFk4T1IYs+ywBR3iOmKPHkmqS2R3GvVawWR8DIdKfSu9Ji0
DO8YdjGNh7eNbn5AprJ6BpzBWFF8hzzjqgzJDcBEO9tISFiDXG8NKNvpK+tjQbN0
lw+Gt4v5w/LIe0PbHTp7NT3pn0oxZnohMlnSSTxW1eMeAMhSBvqG00u6tn4iNq3V
VDMQD8krTUiZYTw8pnAEX+JwCdoEfdnNJ8Jee3XPjMPy6RPwxwRMSguE6Rv0NF/B
4SrYcoxiwvJvpYfXpYpREVP43HSmodiQIo/1mrS8X5dBnL29q61CZuU9/XxSoV/I
Pc32/ir7ak3xG6dyT1VXCPrDPsMi4FlfttGehqH1xZxf60Tzu9jbiAGlV1i2QBJu
vVAb96zIjhXrgIWDv/7mRFaBHDO5QpQbnCe3PU/EIbgaqtt6guoljgGQfwX2qHCh
zwmAfmz6SdlwAPAUXNMCxluND4kIbT4BLcfTSAZy5DywGxuuSfT7eONLA5eK6Siv
ER8DbRoTzMgAyG7ewmgRa2MVcEf/WIRlErr0vf7ibUKiyliSiSjcsB3J1XM4x6Wq
7SJw9Dx6w0ous7nVb/0J//R9bYoAO1RYHNPCbx6Woi/iM+xXLCfztrsXCPZtkptP
AhCWdA/ey+qakP2QxstWbjedOw2+jlakjQkM18v5Auqa6BDqH3rQGzqRdKU3sp8/
7fuCoO/zvtM17zxetjRtMAytScXYs0nPHPJqso3d8HO/YF2gPHimJvumXzj968Si
Z8RoxqWH0j/rnhduR3nFI4x02Od9qO/jl2HYWh6OtARaAVp9Qg5D2HHfdcxFR2SV
LA4AbuqSfkzH3+HYAyP+X3x9btgCEbl4CIUU2f7kNoKPWJ4Q1Nupbceu7OHkq6ru
CXC7o09ets8+tfrgQE+O+gA+CXVK3aPH2vVj1kGLq87clp4oTE4ErXD4cttxNJGt
EZhCvbRYUCvglzRsAWc/Iq7XQqvglvdYztEQA5QnDu13+8IUzYPRb5Cv4Ppip7DK
OPnJPtWJTLY6bgkqBOEa7cTRcmtQ2H1Bf9Bi8vU6n4pJwpauzibGZG3EHkeA5OwF
oYMOiQamTxWRV1HXXrjYEu44zZALaVge1FSJotKO5cgyvDFX/bbm8jfltRfQWFXm
ybTiWiZsXEJm77eE8zh0RCscuyH0nVIwvPZsK9SeaxP61SSWHu9lQZs/m74YYRET
pS8n/A6gVHxqhYaPH5vEN2hb6QuquwNOvjqVkJ3hAmCJsTfvYmbU3QAEemzDykM7
A7hOZZKn0SzG9HNpG1Tfx+6rwv9yB4veDobaVLy8CglYa8GP9gQqeGTgL64RwPzz
Oe3nNyNG1bGKvxnH44BUvSGZop1ibT//RAYdX8VD/thy146SP0MHutTAoPA2R+R4
N6VDLvJYp6E++ibuLiA4IAIFgHmHFn59F3NJkjo9ScjtCJOAYULQ6KwHb2fXka20
RTUI0cEGpQuUsnP8IEAkTZWOlThYF1bHStQNJZl+PQ1/qcXeViN7AYLnEr5U5drd
qmXEi6gvJaxSzcB8aLkmUy1XyYNYH49J+ltabImWn99j7PMPRIBpN/zyDQM+EKz+
6N+ZTThr9X8YPytKbBoJ1WR1uaILO7NgaI2KLSSR6U3AKz2L1rFYjBVEZv98B2Dl
WYYGf4oqW8fVKsuGFtBrr1FLbj2AJMkM6lMjUSEKKWS3WsULw8Q50mwC1DDfi3/z
HUAbxUgktzgwMSww50clCguFMTptyWIEsVM644ROH+WIbAkoiPYC8xWCuq3dhE2F
PBTddMLIG7THDKpC0pYFvalFjkFDB4HF94pE/lWX+LwddzST7XC2XiyYBWFicfr4
u7yfDn9AmtdjOU197lRBM5s52GC3pjMfKuVszSi1Jg9GmvC0x/BTbuNu2vfivs3J
BGra1dmQ1HgTjrjYWwxauT+uo1rQdViNjDejUfQuXGHSErSGGDcboBUhO3ynh5Bo
0ehKI2uZQ2tjbYmvVJUHahs2GD3X+oFAkxWM1nbIYgY2yor3mFOSkoXByCtEQxeI
HhReCQkpjSBne8U3uyD9EPdPw2kesleDsj6tCkzfgASo7FY3ofZZdFNYzje+h9mL
1dKBJqpQfwQE+FjwNYEIUQywxvHtWb8Rg2QDg0kw7la88e1KI6MHt8D2xQlO99VK
SrPKEh2dYThq89+xS2reSpLFKkEC7c/vIFnWzdUH6NI7NyDUa/mFKB3oQWf+No6u
uuKWjP2WIAOZTVUKxvS60jvf+r5zX6kRK+ge6Lix4mNouzSvq0cVA/P0UEAFhq28
OTex6d2lGHrd7aRgrSvH1YJlisdBmgE0Orr0nxuXSmv3I8ww4C37GU3EGzFWkZ10
6NHCr+MwQ4n1Lxmm37zTt0fBZdRIuNWgF4KmLM7JRDLn5QjMX9SfJUpoC/wJglpK
9VTus1uuFuIX+08qfnoFd7e4oBqnLXM/AbVk2dIePdsmLvl6/m40P5gxzI9wsSKZ
fw/04NA8KTH0c4GSzEiyH0JUO42ffbivDmJdiklM6fH7sfsJtpnksyX3rYP7actU
+4cDutn5U1Y0gBa9ydVQW9S3mosbNfgTDE56CkPgt4pPhM7950RKlupwIgXv3sVh
rhS18TiIIhFWU31q17xzQ+sW6+0ephuUGmkqy9RI1lzTFqtRse6dnubqfbRtYqbj
ooqb+OlXOwU2twVemuqBrMCUAmgHv31Jn5kGAuXiaWaPmVI8wL7sQJac6NlQ3F5t
c6zDBn/jT+t4tcSahNdO0LdLaayWPUG8LVTwdIdQ97VMq+6CwoVJQIDvTvyiM2mz
RKAbRFSsOV/bVPVrz9iUtM/Qpc96FPnBKlLDDfG0wGC9MQPqawiqkKtzkH5GPILx
6FI5RlZOE6vhw0EaNWYDLon7xkDWfubsq8dTu8DBkCu2vwYk8Co1AJyb3NBZ/W+R
1NGu7+FQPAJbBwERYBiYBL40XA8XA3cBD5kHrdDe4P/rx1QT7rzRVxTfAnSe/O1i
z/wincfIkIRHHi6jp5TFpYtTN2kLDJYMcqxtRnIUHrZ9bcl62fxL+CfTHPd5Ue/2
kaxXdDFnj9hvfJuLg4/2ZdnCoMPA0X6kLGTFjtB5Lg+1Cukc4nW/deDahbpc8AmN
57W3RNZuIt3OkNdOvGJgjyVHK/yiOgN4j/IdYaCLT4uOOY3OYtNOeonaMxeG03sA
aSxQolJQ8gv3WJ7CZx68HLX7c/HepwfiQbh/a0wezH4JttUG+IU4MKa/8TXd2RMK
PzTBgNqZvfgWZHgglp+OieCoVOOvOMZ9qhinpcxQbLvh8XWIIuxVAqpaKxoNrY4X
rDqX7gqPnMsDvWQ0ICCrx9vOrFMI5TOs6oFAgjgPD/PRoYFs0rsfMPQC2sFIXQ9G
XCxQ+tdKpilKcTgrJlvWJvS3MxvPmuVn0yW7EDg0Ct69ONXJK6FdsQpUrUE3f/kP
RFof9GycsH9abRDTblUqmj4mmndCrs8jnw55uaiYRVfpnpdI5Y7hQa7M1zG1vtrY
MfeclyJaD7G5LB+kJNFb/1eh9ppFoljo6jWNF0agES4fFx87UMEFx390Gqwh8BKP
qWABZJuFsresqFJBTZcUQxiCD+bpYOZEDG1ii7gy//dlD5OrWrt8nF2TVNE0VrjC
WUa60c/F7kJZZqJPiPCdRZGKTQlW7rJjq9HufpZGa9L4lJNzDaFdcNnUSf6SPtTM
68Ton4NmoqMt2eQcY0Ujo87TkhGR/J36XwJ+FrEtoRngZ19ckXryEWAhBNthfDrv
LYHt9anpT+QC2pXfX4v3adgK8b46sMZg6HM6CRq8MF85BYIOgN4Vefoh66/VHkya
rfDTv06qqAPbnD8T6JEzfcGO5jBiOpUJRQXsHZIC/7LtIBn7vywZN4sJ439eWO3a
0FXGUmQWASfl6SHWtVTfSrVYpBqy6aqL20Ljq0peKubvwwiZZEbyiMFIZkSCZb8r
wA3gnO8eAL4STIXriFeWmQZahvk3MHardXIZ6243rTlBYItBGPAYg0/zO6qfdbkb
5NmD0seayiBMvNLm9WqHhWjdxwpWlF/q1YUzv5luvm5gmi6LHezKu4PYEWdr51l7
TI0e4IP7xKbLYxMRU2vzbw9xXYahkplEz1tOmLaE5jxGf5xu2kuO06NoHalqzayX
9zb3uDdDeEw4GDx0nizEgmMjGm4jbmHVKhs7VE7Oc9gciX1uu3oQtlRMRQhmjGpy
lrvXXdD1knS+UMU+N+o5bvgVHCGWojRsS5/Ue8Jk1sj35U/oOLgApLxe8VBFguBv
/LRtHaUoZHTjTR1l/y7FA5gg2LH4HTH1q80QcT+BobZQzCbDspHPKs5Ka8yUxbcx
CtLLKTVm+U5cboXvv3HcJh/De3wUdTJMj3tc6xuxpscfZYLgqRol6g/YEnDLOymS
R4KQX727QUlcMY3rveoSLtwhSpBHhsHz/upC+Qd8fpj14a9qx70qjQYf+ureMgDB
w0mYUrCGl5L+MfNo7FEXUK6YRN6BgN8bKizwBwPMInZg5tNkd2m5q0fiobZXbAzM
UYTRovW5u3fAFJ7mpoXfn33YJ7SF1SWMdkvOpOaFH6ts/qZc6CTyAjP1O+ZwWbBZ
tF7oLupAndB3E0tg+f5nw8JFVXAu2HDzQ6y6lkkhnfKj0qUl+x/5+AXh2XWeRA4z
r3qGjfXnfwH0iwm3NiQYPA==
`protect END_PROTECTED
