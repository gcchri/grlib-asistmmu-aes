`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQaantDkNFJHruK7DFjbaDpLf45YcwZsJ+Wn+O2g31z5kforTcrUYyaMpsgP4TcE
v+7jax/NkQAq+iIlVedATpGNPeYrBfx8btk618aJ4/KxSM/rNXTSobubWwh0vPqf
PdXPVNsMy3n/SKXZIbN4GSP9zy7TY8J1eKoyqzPfyQqjgGD3s06gjvfjIOAUpXil
2tgjf5AvFNkR/Vk78R7c0vnmQZaR8cIrSC0B5BztOSanAQPU6JsRg30bBz8zKSOX
AMIEAPZDEY02m0Mx4UBInw5cHdWegoU/weiupWusTJqR2WhwKg/faFlX9EjbTV5w
kkkM/lkC0Ao3/yV4w6O5n60k3a7TwjMgG8mh9kz6jjnwaTopOJLDJQhjv7/V6sNR
bizxPr1FgaJ9n6+B1AJubLtrmYAlqkzuum67j63P0Hc=
`protect END_PROTECTED
