`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMBvaG8Y0Nt0xaBkv2nz3chF/ndE9djm/gzj9oN/AZbqJgwI2/MI8HrPK2N2b/UU
FM3IscL6Wgm/nnxuQP+SUTIHSc64pDJmoZYhd7UibIAJ8DRy2FpLZ0UJpDQnck+5
AJZMUsMftQbGPMry63kPsNUqGzKtSLoB/d4vlagbcy/Z9RcHe3kinWVXYazJhQAu
O9trhJhEPjlx/fG+Ye5ICjTAK3DbfX27Kg72FQec5KJHa2ejYqvXnMk5q+tfUq4n
JyBsQ1MxuCoeI/XDK6yuxpXn24rhwdJAjfYeOg6LjOMdIh5NDqNngoSBQkx9JJhy
M8iqWUyQlDz+9FwZrU5QMcdQ6eZDCTjQxT64YWrhcOYpQFCrHE80n7mKLsMV9J3o
iJjRC/3vXEgdRldoldoEe4Awdih5BD1Loor7iTLyUDWQsgjuUSGz+fJ0oyqdBbL4
ujIsR3cgGHe81Pi9piMk+l/upWbPdfkQAyxVyIe4RCugrchXUYIFM0TJVnK9278K
dTD7PmNHtIEDZOYp5G1zoyKfHl4x+uMgR8MKpGTftj5/sW5jG/S/DVe+dRVRj8h4
GPHKBBVZQ1GrpioCTSAoDtyprdkqYJ0HaG/ec+IXZiahGod9qZADH4VABZT7F/wQ
pOIf4Y2EmlmoA2CaUtTeG/gsfOLgDbht7cOFIYNNO1627F4QMhFw5m/+38UzgT8M
cshp/cQFY7T6K3Pnd8jblsR9r3CbBBJkT0ig4Abhrpk=
`protect END_PROTECTED
