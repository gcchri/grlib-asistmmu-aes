`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8IWi5gUje5DWqtAC+ndYpVVb5pyeH88EhyOpqp/jiS1Crr8nJV5Ctv72b4PJz3zg
avLoXesA4Dbpg6QJ/+YdxhKtVKZfSHAhsWC5shLvL4eeE9HucvUCt2Blt/snQh5r
K6YMTP0x3MDDunfBcxF1vjIsfwe4Lr4QIaE1lCJsem3xQbLwkZmHuFu3zUIEDF/N
+ZW76nk5kwsBGxq8jxnh6lHiqYy2H/hqkW3i4pzxIlJuwQq8dcvpmhumB/iwNdNh
OUiE1FTzw2TUpw/Pj2Oli3Nw+ZBskTXfMTBno8/Gj9zhNiBS+wfZTQA9TxAJZTwp
V8lhqemT1yRJEoMEKHQYXaYqt/KdqROIQVEP/6mAu8MT2h+w4eBbxKIYlWD1cdFe
gKs1sq4QvuEGtUTD/lL2aXagVNvv6oebmv+0qMmbSX2Ht/H4GpULQB/pW9ZVP15e
ZDCjgxfA/4PTDiaQIFQqBrQclk0cthAoXSrzoxOATLc=
`protect END_PROTECTED
