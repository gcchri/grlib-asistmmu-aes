`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ftdUY06Zmvn7pp/OuyOXP0wzwgIlq8Y/UVMs+DrJKBtl3TFmR6K0r9GPgg7SydX
dEmwh5p4U+Pl6KYvJoCvW0ZKRK1ynSo+Onw/JWv4FFZW4OspkwGBwJ39O4LY/6jf
5LimGvNh84GJrtVfu4BWQqeQT2K0wM/RVHDyty04OJ1lviBXFmvvCqO01BtcF+Hl
7YS0Vr+G41xA84FpDhnQMtGKHO6gqRl6OUKTwYjrcoEjBqUJw4UETHBsyoZWSgxE
Kth1aPHqubkLfcSSy3MPnE9RM04VsgPhnDLCH7220HA2BhSy6HlF4YotEyxcq4NL
kUsn035BmSxJWQCSqInU8YRmeoUZuByhn5xwcRSlGD46voJIN0AvIO/zhwkTQWeN
2+6eAS+liy0LnKwtJJ40D/OBYSYDH7yWUV7lu3rlR+6kDQjMBMgEx6ZacKCzqlV6
F6YpS4gAWtCIVI2zzNdHUiDJRbHtDhZ4zC5Sj5jjMY0YJg6NkL7OWoVN27k85iLo
GDjPj99D9u+ynKsRHrUpNKBSElizu5VNp7IPOfNsG4pPHkjHPwBDc7TTWxJzjjy8
tjojXHYKvp2x4ZtXA0rDvqJfau0peRiIYVoLb70/hiG6dm1szX9gUYmQfq337rNl
6AzK3Cf9UyC1Mqgq6auYn0L1YFK5Imd5684kGK2rHAWtourm7lXau5CwnKnvT4h+
oLDc0ZJEE07OT6gMkrYgRsefHgAFL5xJ1XlLcqhsmJyAnDTuUxJlLEy7arQMxhKC
x4VOq5zj9Gmgrf4MW6lFAA/8t5yaWaSf1qWnTdNz3zlfQpG0lcljMSt+5jSGpqp5
yTsXyNHLLcaGFz51GnFeJcU0vGgkADwMDrg1/qyZeDVhe34/znWrwb3jrk9LfvrK
ICkAvHTrhVHRr/1MMhj1+bXA0Sl7sEOiuClSpqfCAZmcd6kj29tnAnOtf4qjASBZ
m5dBJX07npPC+qMhgmkhKv+fpeV4Bxr/bb2mjHfIvVCZZKL6Fy+lNM8QQ8I4c3ZS
`protect END_PROTECTED
