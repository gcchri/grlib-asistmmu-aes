`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zA3eaNtIWvHqR4sRnTp2/EavrtBIkDobuEpxiJNHISZaOW3C64vkpmDNeFBb2ra4
OfgrWM6ehmxCFwjtJrjfna3y0teT4ruOVNF7QO+VhT3u4p86KKthrvN+yQhJh09O
pU6G+p6ToUPY0TH+jfmlEH0VQlGpJ67RNvnW4MCiyw+U2bZk3R/X4JZiST7eIQQV
LH0falVaK1iURSl9S19y12MapA01x/6FlEgNAftGpWGm6lKcFdzZKtl9/T7dfuhF
PDDQwwfmDGuvFVkCF0z1iLX9V1eNFWzioJ6PImVBAhZ0JyqVaYy+CiBPZs9PabPv
fEA3hRVYHHsDHU6PfPwiyB6oGge2rvLMAOidhNxcxp2nsiBW0U1q19MAJJLZmWsZ
LR+ddvK3Mju7zM8ybU5guQ==
`protect END_PROTECTED
