`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Dz10J+OBviTENWK+81Tp6sYCV+K1enbmsKp/kbuH+KZarx51Jd46CeCmUrYPVwD
Vwx11PeMKnZyYn0hXqcFaK5V9YvGhN+rXj2GETexwXKnmcHDUWbEhgYGlEPJRCBG
Lws6emIy9TKMVxkwx6ltx7FZDFtTxayNFsmYtvbBzM8gFmHQ3swoSgi7tXBfc4E6
TO7a1uQLTLQudPjR41JvS9AJHOMVPpn2dGw9dUqyf9vt9xfMSK9fJJ+FtY98/B7G
VHYjjXltQB8enw83s2Iv2pcwRAmX9S4Cfz/yV+DBU1j1PY7ZF+HITvx4T8j6sORB
4KZ12oTktjpt0G0AHttb+W3sWba8zIHjr3N+OdBtS9bJHKInjf6+gMM/R8HgANT9
5dK6nzHynJNLdz0Vd2mdHkHuZuL8kJ3ekf4OHP91kwwbB+1gKXvrcTKXkr5N+Cgz
uDe0bqWnaLvzLSJZA8SYm5U1w+LW43zGMP8oh6wP0EReXTXS0T2YNZAkusUgBWid
aIp/1Cd+aeGZwzAwVy4aFhDtZhRpaBtzg9UgPaXIeg+RrEumGmX1jLRWDxzdve+9
dolkq4FZuSklemgTAIgdiiwkPLyqVR6rFpjc7TZieyxMhYHDAuXxpI95e48UeV8q
F9MUTrOnVbODkYrqYnAEi2/Lmw1PSHUSgyKDA9BygYQRE00fLlgYzFkcKBrX+yjX
cE3uF1ZBBiO1AP/JAJlwpmuHVhe2ofhmVx+f8AsGnu4GPajResPaSlld9TA6yeNe
scEKSApmmdyAdsW1UOP7j2v5ZPWnGIT8Eu5hJwuxhe2Op02uAU/I34Xcp6j7v48d
rOo2Yi9KOgQQL2sqTu1iZB/GCslWxbeVhPQ3FChoig2tJpN/P1NeaYTrqqnCS4AH
8NemBTmN1GzgUWxMSPgVsR6QmrbDqVUIdDyCNUhhkwnhESSwkuiyQm+OARcnwzfX
B4fXEKnASFx7JcxOlFfJa8v4NiZjiKtHrpyzp51NoMBhDeKA8GPASJB9+cqddSlf
4KGKFXdb9EhVji6ZQpPZaku/jyM4FCSCE6+OsMOmrdwuniZqImEIQygf3OlIrTZo
`protect END_PROTECTED
