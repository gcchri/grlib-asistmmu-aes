`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1pHfvRnq0/XXW3o7QNVK9Zj984DdWRxi5fuxroD1i3VOO6CEO7HRIYkixm0+cP+E
ehOW48UrmuaK/nf5GEsnOiByf5AQ05jmX22zs/7bmrG0sqM85wQOMPuviUedWQhK
IBENEoEcOp1r/9RkMkjfLkwulHg8Ngcc5BEbq0VTpS1BcQUR/3hoXGXjtKFsWCC+
HiAD30v/Yg1QLXPrcKQ16eyMeZnhYh4hBNEKPxrtB/3zy5BbvKVVAOzjsCiub1nD
ONvB5vpjpreogkWJszS1Zqy4UlPdbylKKEKT3db/zQ0zDKo28Z/MrvdewUkEH5Qb
QN4li0MmKCK/nM4tOdkwLclB+PupBueyqlHrU4D+oZVg2HqvP8feOQXOcFEmkO2b
KFkWjdRKTOjMgzzN8sACDbGQ1lXmvxf/QYghItZXaJftEgTI780Yx9/ck/s/YFiy
PKGlL9ioVmtVO1ZcwLB3vK9ytBeJyExU+EfPxt3Lr90rFvCpDcv8KwcW83v9BoNN
dt3INljn8KfwBHwxtjug9Cd5P4ia8JGZ0YxmLEOlu6qUKDJmuPCgYvLPQZql2gms
oyYVle8rAS7m51ukgJmREQbDWpmVOallmuMDQLojGXhhjZ3isOlpCqsYVER/62Xn
K4suPGUwwNn4D8PxxnE+5TE/BJfn+U7JFffa3mN0Bf68HDc2Xew9MIQzadbmT1dX
hYwrRwjn/x5ECOxPXXzgD/anbzX6GQtUGfZfHanj+Eis3ZIVjIhxU2bC57ru6D4A
Vak1z293NeNzPAD5csVKUg8p2Nmdz7JzJxnRL0hpUx57MZlDesTbTbwpQlkUmaOn
seiycdTMJF0KNhnneSe0Y0WlfbGkh10L1EdYuYiDKOTfgMwkwzvwLJmPNL/mN+3F
z2a68/RS4Zk93Bq4QHktSEtTUzKkSduSWs4nXTjxiOC9FQgs/HLkcITQRi7L8/yh
OLANK6LTYbb4YSCb8AqlqGjvCmfv6IU+9CbuOZcA+c+iX/UXfiJhnSSV9t7hcOnk
eicWPnhFdkuI3auHfv9zY4IDcX2w3LEvnbFJmMmveKxq49/s7odiffqBKHbkHIVG
3pvMH4ro19C8IWHueVxPSM98+bHi54CnaJCjXiKqMAGKFq4unYuEGcYvFa5RXOws
4+TsGvxgEobc6SJPbeLlcptnoiriIhQnYjSk+3CJZZWlkpeJSnOOXq9x/h65xXJL
2ELQYysvUVdl6DMKwykzP1O9WzZt4IIj1iZylQ2tuh2rp080GqeJrF8x0J9BfBK1
Xc+Ku2vVZd4feu/aZgDqNlcpM3A6sLRAcvpLamAmUgrWaAQSB3x/MLGM1U0144an
cnzNb3N/bacS48RTBh5iefkjFM15vrSpI9mI11xFs2pteDMPgVYmJzAwEz8R7NQl
D1D0Hr99a/4QtmnSeGRPu80MqhixcFf0wrtygHI4Mk1m+xrr+78Vxbgf1+LQvtxg
bjekBUnQKNwOnxjOIopRjbK9PK2meNgCqA7zSJr9Es4gfrtIf0rPkVvdPifP5bWM
otMOudNB65QW15N0yfIJVOThHcNu6G0YAJ2MRM/CwNWQuBLAsRmlrXXxnL67UUKN
H/PahvYHsxv2vgkkswqEUJ5n0CKAKKTAhtt6zsMD/sherJPGGKTZHEiUheQhfYB3
gZlHaOQizcA6LZl3SpRvp0b81ko9mGQV2Wxx+APuLb5BSGRqJsmTq8kTvldtfJtc
TrzHwigiPuaxBMaSzfpL6DOtey4uh63TOLLCLDwVUYOexvEBhem/yk7K1h0CQFo0
c9AkfO3t2okIDMcdpqgaiK0MlAeBiSqDRD+1AVUGzAYP9IwIr23H1rCUgSEjMJbd
XAOV4i+9z577wf4jIF2yyq7sR92/BAL5N6mx4gjDyYu2Nt5QPhrzLSHXdJl9Mc+9
U1MQgXcv3DxaUnnpsk6WHVVbLRDfytQP5Jc4n8xD5vgjENXf9a/q5mMJjHptnGDt
yNNd/mEJJ+xUjBvXBO9nP1XuLmSuh+wE3YxHLiICX21nd2EXNCnjdwTq641VClQU
Y+aj8fp0yE2vrWSc5w435qumSq2dc0fuGjQSvpamtP+kjKW9+RuC6LydzmTwy5Rj
NeThlTaxDDeJRzumo5J6BpYliwgtxIgzTbsKZHwwH3gZo3FGhopwuUs4DgmyrhfW
3QTidSBf70ndEjLE//2RRpFfwlwkeuvkcn3aK9XfQgPBJbViK7FVLj7NUVP1DK8h
U2PuUL4lQG4utZmWG+lPfZGTk410oE0o2YmrTjriyd4ebv/tgvqGTHpwuQPpDVwF
3exBXYb7t2KGRweal6r/WFkgxju6oXBpSpxw7M4JNYGrrxtd7GyzMRrRqiTEps7X
/ZuPKQK0r+V7Zskt6UpfC0WZmFoWVNHjYVLnzspxirPwvqDCueCZBiIn0HOW8yvo
Uy41RYD5JcT1FXrAZI8OHdhSca16BoZHjyfFvIa4OYdktXnF03so9U+8V6HOtOKr
vylCRur59aWdnuX1uQy0ayj9H4zz0ZPJEeLr11XBW6oDRdX21rF87asAbGAkGz78
Rngwllw4Z3EXz/5r38hz3Vwlx3EdULwKDokWm77QSbeTh2k9WD7YecqVUJEcvQW6
5zSQWha1g+26stAeFkPZ+AmE9cR4GdDdJ8xXZ9D9ayWuEFBnCwNp+2GpsGqHsG51
11PLJb7L21mQQaRXf5GVMSJXurm/t15ixOpnaXJbUGiCp/MYLQ8jdiJtNvYlkbPZ
wSIIxULfDK0lY3Cl3nR7eBAMMPz4cY1H4BTpyB9PTaEYQwdhwAI8hQxbPJ26wfR+
80rTVsmhSG0kzs1ihi911swmKhNze2d5EDq/CVy2X4Y+GTBmoM9Nm6NvpPSA1Iul
L6vSvF6wddJelomcZ4u2bc9Lqv/IeI6bzTf4Q09sZSSgksWsI35fQTiN9KIVsJwI
LRlm/2ma3dGRPdke+aO4Qq05RTJmLzP8f8WbB3kuzrFqRgYldvxzNovics4H/Kcf
V20jIqdWLCdCLKk2ypeZ+5ogKazKPZ2jPxDaglWrJUIyx2AJBT2tRMV9KDA65OdJ
0ouXwIXJoyCIvc4Vz/KNfqdyBDuoFCL/KooUpgiGoys7RtA9erd7oxuyUYGZmZ6j
yHQlu4EEpqK+A1XixQ7Mo75sSIPn2djR2De1c0O4asEvY3Gq1YaAJAz9A4tPi9k7
gGeCdtJKOU1tUDwDbFuB75FclZ9sbn+rZ9gA4l/SVJHKxRHHQk6chEBgt1JVa1ep
acZ74zqFo4rQmPgJX4vieShfYSouqXyM3wQx38WPJvfRnXLzeeHqfx7VDGjEzGUg
ZraP4FbrKhfA2GmJE4FZiAOj72UOAEZvMHX5uqkPVG18p7WT8Y/NfRkaXnfzUNsW
Jv1YkT9pyzGkAhHf3fMvISjjcV3chFe45Cm52zZbegb/iyEyQ5BeOzdblG12CmwL
tJBl4BQxteUUmEXfA522tq/XklHCWpKUJCUEjFN9tVunyjlThccifiRbXN0fCMSJ
eB4fZTrnJ17psn2esZvLNvydMHnUjiE64Fpqt5kPwaF/YmlmiEVmGlL3fz/ymIiT
yV+P9wIiLfd+9KOT4Qy/vx7T4Pt8N8cIvC707gY1/xJIoM8u+IY2PYI54GJw1H7a
6yie0OGiGdevi1BLgEYWrGLEcEiev4bqDqLZNclGeS+8YDs7Cf8zswfmVAbtHaHG
z9XrqUrxFkUIBhSeXn3fp6jwLmWIV3Jod7ULeVvWvOvC6lMH6BKcTMXzLs5Sc9/k
CE3dGI9VMyA2YdG7lpM2osoKPzJhxbBzDVQ1yS4n0C1QASn9rWPm1+q2GJ7zjwoc
rBRSogHyO2EfsoNKNAiIMPY0j2Pv+6wXEIpIx/AgCvRyntHiuUoIQz9NahIYM+TC
mUtHX+snMUogilKDWqtiVcG2vviRPT4Tge0HdVMQffWKkrEPE/oGCXstRkOXLQod
pf4h3bbsTB8egzHeLoiTtnh2NoriM0nxf7o0UJB0rLg0wvl8O935cNSiHMDqtU0Q
UUBaW3EmmwUuYhYFwWxI/2wnfYy96Thdl6oNaULfFOvEwJ/QxAv3a8tS2fhEk3m2
UFYJKAoHMvF21gHofxptHchUXGE7zF03GYpA4lkLrRkD1941b4qj3x9kO7plv2qU
iuaPiSxTKLZBG/ef8eC056OiAacdslbuhdr2P7PU3Xa69DD2toZRvjP2BQDnQXK3
fO186EP/rC+QWroV/7P40PAhACs9wL/aVPV4Can6qOjnBE2X1x11KF2Xl/L+TlpU
ou4ysFzmlNeMtyb2vue1iRswG+tXX8/Oh7RUxb/egkYlMDzBAzHjpdnA4MWzRfsN
5wYM+bCHGh/fjPrYQS1uAIhsdt8hYifBfherHM/abC9ZNC/pZnkBXWcH3CYYL/9y
9pwm3ePv1O1VpBkJCNzyt4GNSvrm+KPj22ZpNb2vbcZBSz4kKAda5Rmq1XvdYKrB
bxHysOy8op14eQITneifsI4G4OfS/pCHSQrmdHZ4UndIZp9/b8UGyxvoZYHo/uGD
1RdG2gUtswH63bGGlxMBcLlCdbesYrFwfrMI6BqsIfJNg7z3pOc1CtWIf+R9M1r6
cffdigTvMWQoidq3q6LaoQ==
`protect END_PROTECTED
