`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpeQBHNufp0wfAfNHsGZmFzYkcsm99SiNGUl9WfQkKpXsFM0ahbmCi1+CVk7mHl9
224Oy4lt7Jdoo6/nyPugost2FWybUYKXJMiAs1xCWz+nvskTFT4S/t0pE5BduYys
l9Ym11kwQ0GtnuFFLYp5+5Nn56fbLNHrijqTHTdkdTqVtaT/aXtLRgPr4b+uFAba
lYihyrpIlLpLAnFJhmFCcwzp1gq8c0Axh6mM6qG8lWwD8Fp7fz6L/hWmqEtu2fKb
nsSoBW1GEfUR7fUse1eAB5j4DsDH5FNEC+0WjLOfYAK130/BrcD5ilJ/jBb3uIYA
Ok2gpHdoll1wdmdGBjTt/Ejoks/npdDt3Pr3CAsReScAGfp2+lxxO9/tLXzbVq37
ytiq6lwseBcn5hI7Z9syBTG6ItGmM6TaZ1ocHocs5dR6XUP6DWvDcHLXMSqHMlLi
jddbCfxR6WViSaGnxHB+zsYJ9XFX8xA20SgD4jZi//tnXFS0oKPH4XYiRszTVtxh
PiYQ1/UXbjL+uTx4z9ZYpPnzTV2ogbT8LwqJsRpl/CAxNTBZgHACMMpMoB8oQ8/F
kpq/jNdnRycimixhWndw/5H+mb7z3m91k4F2SiChbou5R3G9liGP7p6UoZn+DLRT
vk8O3Cf9qD/DSm7s69BN8o+//OyJOOuDq3LIbQzwe2Dxy9NjTq1YgbZMlR5uYEla
IXWFjZba8qkuzGyym20/C3VXUnNWoU5P2mirVENb3SQ=
`protect END_PROTECTED
