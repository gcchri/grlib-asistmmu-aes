`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVpw8dYqZTdhkI0oyPoKw0xfNLilWCGA1BNg7PqzIuXfHPba3ohw8A6AlJ3lyk6d
Wai0x6pLkam2yNhb0Nzc/CUZeiFGh/dbhr7FJtfGqsmVkJKFlXidP01j1NeIQipX
rofGGIhZaYvtsxWGFD1kqKpAUpBLAGAU23CBZspscffRDDVlYVcKei6TkOh+UdYk
8BRq+6IQu1X/7spNLDPLS/c1YU5w279ubTqojJMOBlUX/SVLokRlVvevX7UWc4Id
fsU5+J9pwyK8AtW3ElZybaxXQ4cqSLZayO3HdH44sVbxkAs0RMoe41SXlecU0s7Q
iHj/bbBBsGA3P134m28DXk2GVVQ3utte5lWGgNwZA7DeMAOYCXb/ZLIME5SiJBTb
66v2U+MrcDfX5IXQPmdDWdTpa88Dg5gGvwe4qTiKi4Y4A9KGIACgmhZDKomHEqSB
y3Og8GtxsRFlxD4BukPOrwlhM4xA0UVABOO2qS59lEEzu40Nd4XhxfbK3EWUYECb
51ApYJR4wJLHLlg+Wsr8qmq7CsUAk8GUHUAxUFVaLPCmI1Z5dBSMjNxYx/trAc21
`protect END_PROTECTED
