`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tCusmP+B2Sy2ZmjVirPcj/jSVkYKeOM1xnwZV9Dalv9jfQCcT/fO+yEIBKholaA7
XN4TiCQZ3GEJd18grQiApB5uXw1IVpCgtgug/DbsNqh7wlJdEBsphrL/SZHf0uXF
ZtS6KAXVXqhtX/pJyfIfm6kSmLxifn8djHesMQwGLsNHkhlIb1FcKW5SD3Q4XPgx
3BgFHUhVF9h0hCE+wHaMM03tHo3M3j8yekdQ6dbMjQy0fMZ+YWS1CjOJrT25Nw6K
gtlWFWfEItTmUXShCoKiWEp+HntlVi3f5gYZlSV+UTqo8x3ilMtY1JmAftM/0USP
YhlBCeeUrGf18JfJPFRPMUiYU4FKQsSnOC+Z6UEUPVxi2YY3lrkkDuvh0uTabKR9
JbHBsz3+OQnSHQ1rW+1/3H3h/m0ilkPoSAVmDrjEj0vUyUKlP7pl3fuYq/uxWVAJ
DAYsnhEfI3aXRtH9V2b6eugZl06WI769QADcYcaIh4nHfyZTgIVKvRyU90SfEWcn
OReykRZ0t5LeA1ErDix+FfTXY2cdG7ntOkIzwD+PkVq+jpulq7qakW/Yyl1TXk6f
2bjf6eyCTJqYte3deQY4NMQaAuEjG4/8LByu9Eh6Qpebl9muR0qpeIA64HrdNZH1
p7n6ctz61VZ21BmcZmSmnz/beO8hEVmBzzmcoZuikxQtr/OjETAbgJpAOwaU39WB
ZQ/rSBdG46tgxvbfgH1LZij3ameGnKFkpujtwkw/Ilaksfdm/XfhTviZc+tJ9t39
+nwcNB0611ZP4SDt+zKFgjG2VwM7B1AaXqzmUpgGvuTx3P1WbLtYkfcz6anhsIJH
GJnndtAN22qz/PlS8/IkPj5COcpPPlC5cpZnpTUDY/l7ZN4opDhGlFTmoNi0C96B
YpaX50Tnnn2Bu4CHv5FjcpUxGEWW8TnsKyK42IANCK71ioEvmGFHr7llfnqq8Ziv
ZFO4izHM+7qHoO+6LiCm+iAVh4FsxZ/QyJKyBMWmI1c8+epFqOAQBsf3rg7YAFwk
1usEZKNl+ipDWV8ALw2+H5trMhITJyHBzfFzH6PvKEuF6yE7f9xseZc1TC2vNYbk
C+2Xe6NOzx24BUe0qu89QAFkTaM4ZHtPk5zjCB8OOwZ8JKenxpNsuGBDmdFIypAD
FYaNTTkWUJBPrt/3w9I2tBxiKReMku6AUlPTz/nwFdo5+cfwZ19FXZXIy2yAzzD3
3xfQzogL8d/gm0VFC2C2IVaGCJ8DAmo7cpvQcjYla0PVMHVY1FDZQed7Ux2QFKp1
3Iu1pHfzjO0DUgGxL2ItFR+jqoMVG073yI9EtaeuGUzLfIlScmB0uoex0HStlhEQ
vU65PGV/FrG321SswV/+Jru8CX698LqXz6JyeLBqhk1qWwO1bPlUOso18jSMiuoN
5bCQO9uKhNJjqDb62I99pdDm3ZrAYETziDCX6bX8A25jVhcBwrAIwQW+vD/IA9DJ
zU5tXIGGDAGIJ+A3mlAXAclCswL0jCopuvpNQNTpVOL6t02T7xlEspGYbhLBYa2C
YuvfG+swh1ZHgkSQHaxq8B+3AstZJYv/BuH1x6SfE4BP77M4Il2hzpXt8s+vwLgf
AVKZED366BOi5OJaKCYOUpCjCsC5btfZF1VxyIYLGzNs8pAynFkkw+Sg/fMvEenP
O83m93uBsWu4Y3uvCzHexTroa/v8WPeVdlWMDRN9PLH5B5QOWhvrmZQSIYo9LsAV
Fxv/DL1DWOkSdXRQF/xP5UE4GPAuQ8NUPlYzvTBWYFyHoIroy5sRt1d4aOR5eX/k
O7OC5596GFONqF8gjNkrD4cadA9vykOjomnSXNb5CK8Klxswayd2Uwob/FMMSczf
qAd0Vg6vzt4FtkLlkJ8N0E/j5WjFG0kUnBKZUEo6AcBN3620iooMyGNmp78/1N6U
GURUMSrrCJiEFBGV5S1ovDtg2G798WOgNkqDlAVByaGnb7aY2DBkeqG47SoaUMCL
V+sd3Bt0fmNVlXutf4TNIumB1u0IS8a/+HpQzbbrkghASnyb300aHQeqn2wtJpQz
8003pzxVKLtCUOV5C3feN2RV30SUVT0Vo1cXA4gyttq3TWCT9v61g4taVVGOygwf
jaCeYPf9gQ9u8RqSO4EjOGvd/MuHk0ZOW3+mZCLEoHPCwUIbZrcJGLHQ1KCdalA1
ekBhI3IyYNAR8Ct/429Ij6ZtlzrE5ru5zzqS7eiNYAxcnsdRcf9c8hJeo3IhXSuK
16OkcN7guptILj6J0P93GtjF3Q4TQSWFED/V19TT80z4ncpT5M1RmYaM6t59kUEy
p4c8IXu+5WFp9y0ZXyTuLU23H3QLJvKtevBxBczNmCGRfjbSz81vf+c7lEXK+NRZ
lsWcC/SccOliMmkrsLRffa4LbvFTWbmVw/OzizNGoReSqZM+4nwQIzR1yqbeAOcB
G3gugc65k7f7wwwRWmsrKPquuo5cu0SpvQ29o8R4/q7Pnq93d6BCypR/PWc6SQhb
ASGss3tCkW6oLPdr2vd84d2ZmuZf/qvNMxJve14p6GnZD9asd6ikVRU6iQO9QJuu
xaZysI/ShKdUuRLflGsFNbS5g8cPhKOD9m/h9eZw82R3dwxixBqsj6Dshv5Fz1Lb
VdLh07q/BAC4dq/WBUpoiVaG27VOnsgK3qkwbG/dqteMk1jL9ky7foX+BYEY5UTC
aL15xwLHVdezZVxeUXNfwx6UWcUt/AbbPeLKGQJk7BCIfB6FuwO174VW7Z+T0G+X
jwmsbcwvGchkv46tPu+mt9svgq/JhsJVU2NDBxl+2gzu/gmyZVi+LjoGAxY+E40u
b4ybRDjcDh1gjo0UOwuyCi5viQXUGYgqUWiNwOrOy1L14yPwr+Y10cl/Uqu+5Yrx
dPETDvoIonQq7oVqha3B+HRmOQjP1DhpHn1C+PazJp+aDVeqvz80QMAtRcULq/xV
b++jY5nODnsIF7csawBnvU7yp94gnckn/uETCYppuLDO4eSBImYYols+cP8HXA4d
AISXYyFlvqCCfr6baMcwQd57Tr/TgSnewB6S3Gjd2E/nRVyQUhMZdQ3QJ45NmOcC
k1sLYVn9gIU0Km+JkmplrrkEL4CIg7LoMx4NhpwlTzyb9sa66NC22U6j49DrGFTb
SR4b898mav/8pOAZBRPnouqDvMgNHvqJQkcyKZaAn0zNLY64qxY2See3a3t1e1/l
CCWzCBOjIE+jVwidVtVNfBsBZkK9shu00b8jTA1Y5TmnL49Qe19PLtXuwlKaqnq0
NsT03nHMAPaGL1ud2bWQ3y+v+OyEJZMkIYADSDbVO3ez8HLOgfEB1e5E3/2kNOOp
EThA99P/hPyR6ikkrQB14BJvcvAuF+6FVIZR+flqzXKJk95M+ETZJSIkTKbHg2FQ
SBpiV7qlSNooAyU259QvvePYd0Ua0dAJj6G3Kpvq2SyZ2tEO54AX9QhkR9ntyDaZ
vDBPjJb5P90q77lbv/gg/nqgDrI0CLtVhUow3hY3xa+hPiPeKRkl1cXidhl8oQmN
6Uqi5qoS9U6wi5/WOCtm/Vy1SHXaPMGYfWCgsBlTeZFmKh0EsP/C3rIj7sFliwQL
wtFa+Q3yvo9eDPKLRuMPdMrDKkYaWqyaYH/J6THuDOxrMkJeQz1n1fC+zD15aRS+
29GSJq3jSZS9BNNTOLucngDo55b4ATgGmxgo+6+zihB4QgONXfSsbvaKqzP5UeOA
Sa8QnlUho9WRIHaibbXKQ4lZuX8G+nV3T3bIfnyHDpYZo8u9Ujvq0BbAUZkYooCR
p+dQVkTplozwfAIPd9zerYHTtbniH2A6qvK4rapoF+Mt1txEfvPsj2v1ZTP31Sgw
ms7wgzrkgx4P0qXupNLYLzilkTesSJNpFJsRi/2sBUbT2OdPh3qN3FW+Lw+iIISm
W8mLK1UdgwWVYjKjTn2G6g9fK3KAjOYmYK/hs6iH39ZwZWFB58ggjSTAimXes3sS
ETkpzOMmgxBab+CJgCvXIpRsDZIGQ3BifaFhP1+N39VFkefbKOjmFyUNrOQNk6mB
rbE49lODaYQMV/CO6qw1mN9CzCqEcLtu6zEWNFlsjW/dyNAY5QbeLlKgTOvuKJNS
F5rBnytM7G72Jpa/grZcqwdawxHLxGA5dYdyu6cEdoCT7WbIcuGRIyEVYa4iO0ya
kFFxM632mVe7Hu3HCziCKsZSzZoGGryxzl0kvsOutxnjzj35IcSm48/RCK4sSdl1
rtLBxCS+VCLwR7srSdl/PDzUFS44WbHhLCxzsNIw0002lqjcNnYtJU0Kv64h5iiz
dV9HegwBJVmTlm8AiVZ2wEXI8teTzdJtzQK110mDwrrrQUovbVxBwBUAKTZNnNrW
QGN2zBMqyWbuBcuQeDg06E4D6HshF5o+7vKCl71SufHqA/VJRz/ZxFh6iqpp0hs0
8UIbLLVd9cFuz8IAnsSBZsRJF/s9hdgqwosUgfUgI0QGXCLbmmjo3JyJuXP0kNwo
xwRk11Q299n37mP+SpIJYlHPwXY8sHSdl1iVziNISyidSFg62R7hfX2Fd2e0iATQ
g8Yz7rFOXLGWfMZtdhB3TsztWk5Adqo+vn0zzNiVHCxuvcOp/I3honn3SzKk2iNA
cImuvmcpSz8bNkSt2GnXTXRwluuMyKesZZ9UBHjVtaDGSbgkYGfPu0oHoMmi/BBA
P9DVEfLrpEaApvqWhphe3Ufh0lG6NME9+BMNVGQ+rDm2EsY1rUlQ0m4ximGbcEhw
WFDVlLNxgArKsxnymx3+I8IJnXC2QUdRfzLMPYFVugIRIMtNGMBE7wsh576AKCqt
K0cIZySBXHnL9Kiidmt47aTbRFdY18ZplchT9j8pv+lthMM6CFTxWYmbiMEYdMC2
mGIVtQQpSK3z6JPO1lKbU5n55rfqXx4n28zfJ5WHpRQTx3BDyoOhG4CuVIkSaW6j
DqxZ6MWJMq5pwfN7hIDguOyBUZIpbNa8vKPrYrXr3927VWIiIqYzLltW4Ime5MTk
YLFHwWGr6e2RMLhUNv5f2GQT+T/F2Iodv59sL98Ypjz8HnqoWm3Cztg0CSCRhLiC
kTlkk2ABzUc64cOxvNZVo9vu7wMF3Jck3JHaQJ4Gy1yF6xduUPzPc5yBZCwBe0m7
Jj9iQJh/CNaJqgModmEZLjb8n8b2aCZi+MabVjmT5+YjuiTz5EpRA8QbmreLEsgm
nQSwNTwUvP8OtZLObN6A9QlygTC4UNZQM3oPS2BrBcDpQyZFmVx4rQuqpNLG8k0s
ivKCVW1Zpd27BkMveBEyxqzWi5QHKfm7ljW1gfqNEt3lGg4y0jx9gDDz1Wt0UAE5
KMPKgvQumMgj1fo9H3SkdgnHLeU4+adcl5srPRbbz2E7J22yGPM4ODNJfcQaH1ZN
C6bBLajYaPO3oxmY6R/+HzcH/pJiNm9dSRJB/Vc4ZmcrSTbjWMNT4FQyNI8XSPei
yFkR3+Glw4khDvNHti6mSEVn3Tu+9d/OESVUpIQNa2anzC6fXdcC+Z0GsoqjIoy6
WKajcmKtq3Y966Hw6MeJOmI1/mZ8ViKJxKzUkhM0EsesZk69AVo5Uf8Hm36hs7Ym
eIuknHL6FxYawXA7IqnTv/I45Sp2oJip2xTP4Alt0jgrnsTo64ptfJ6q22PdHbF9
EyVb1G1negCiumw2qyo7j0DiRwXxLfwb4V+FTlnDlWYgMyBowtG9kF3PsY1RHEBv
lFI4kHnpMGr/+QdupLUNCXui30Ih2NxlczSgYg2hRlOHCiRQ8xd77e6N+a5Q8ok3
MMd4zXgt/4cVql8Z51SVDyOgagseVTGiTKKTDbp2rPBqfVxJBmtPLTV/jDzsHAR/
4KUHwpomFDmIZiR2E0WxEywyXZf9P5yk5kuzP20/EedDKinLeg6Dwgimp1dZjxz3
C+elEJlB24q1zBeZur7UHVDNzV16SU6W1bGRYRqNPeNf5gu3aEDQaHVQt4u8jEJH
gCLsI2BFqeYmFzjqTVUdYutPeMLav7R1vVS4ZGPXcaZkdt/JMBOVaG+hYJftdKwN
3e9XuAFEa4Sxol7WZKeKXrxjlyk0y1v9mYBjULaydzfVt24IDL4TUZUBogEL0Yld
1b68bYl5UJc8JznfovyFXIk7dB+rMf0Z/hCMesK4z/BNsFS3wMF+BHENML8preDJ
1wT8C2XOYDqeRgh/R85MzsS/2XXqGcscLHAFgrdH+NMQWFc9/Y2s1XAqpmcpMQdD
FGUyaRU3nxuEPOxWf0Fh1F+L0Kiok5Jenc27IKCZGsq+9smh6geLhEue30ECUmD1
VnBFq3bPPPdLQ0FwspSF0dvjUaRCK1mHgMnsDxqW2NChNtN2+BucgqDeglVMtble
sY2TjdNlmQWabs8CRZ8dg9FOBp7IUXgSK7lG70XDz7wBv7T0eqEtAqdJUFsX+3wE
LBn302vTWmNmVKj4GI6aT9ISleuL/eEjtKjAwjhgEIYFuTtGgeZG9BEwiPAa95Wy
fXDFCTsYvZr0RyziLUYXwSo7Hk3GcRXI5+WOEa13VEJNkCxbrLpvpYerGox6UF79
eFecQoiJSIoX3CY/PWfw7cXLj+EKUnxwqqpfCAEXay96oVf9l4GVG6YxLb+y3vT+
Defzr03flb8xeP4HxC2pZlKhE7AyGzuOGYkkNaxvhRJGYqUudExzckFBVtPRx8YG
kR7/1i8cXQNqyjY1dMaJosMAnTQ4ZvPNGJLWtYFT2wlbESd5eTdmXFnc3s6AaRQy
gbXNASnuQvniKKLscY1YqQlPwe+fJndSqrl4j77cwnMfJItsZaOum/4Uh8SirPwV
hc6PV5bkf4iVQ/o01PTbEHoARvfYafa4Ito/rJPkxEh0eiAJ9bba97dABj5uZXdG
a9DSLqQzVJiAQGKA+Ht7KctLGIeLnuYLYrH8k9Ibb0p6Z04EmVN90GMOLyinKYCk
Cd3Q3K/eJ/B0gZ225bAxb3ughxXn4DNGNS6BZ8C1juoRPlq/sF0Tp2qyOcEttmSm
woT0R5rWjjslEh6LILSevjZ/YysC0TkPEFKgy6i4CqusulvGQMDeUDPfrp6/JUMN
ceXvBLsnN6q/oGROaawLDD2Eh8XmHdj5mJh508e6hCFrzA4h7jcMoqSuTtCBQUbw
t5gWQrtXi6KCVZ7Vl7jHETIMpHM11F3wmKA/y8nXg1D35yQ9oIOH2o0jeEVWKjwk
REf2l5c2AGENaBaZ8bYttqf6RQGA8IYO0E2dClt7K9X1+fDBYsc2Y/fQvMhlaNRl
bFsSAj7RZICinwoag4Stgf5W4lX5mQiDVh7sDLS6BBlxyvaGoPmwtxTqtrHfIP0t
wIHpk2iMawrGgKuzoPG5nxesR4G/ghFcUXY7cn+pOVTQW7a1dDJoP8WZbpL4es9v
mcU/cWJ0SCzgnubwRG3dinY6Qv4vW74h3GcblGt3MHDCi2N3E6DpaTjzecpomHjK
b4zTivjYa0ubLKyPhFhJBMiK1maq3eXkHgrcNJZaeb7fQHozic0ukWuFF70Pr4l+
8fRgkVJcC2Khv3iwamAaMnncgM9IWG2a0Sy41mw1PXd4Ry6dqYFzBWG0S4ZzsQ7t
k0btnKorkw4DM1xDlwfu4C++jZlMoUsC7hcmYhhuDMxDpP0r10ovOkRmRU7ozoIv
+RF2rzUxCxcN1Gi71TFl36YTtpcHIrwHaujf5F2PYzFkxt+wvg+LWLBpAIreCpVC
5jd9ZnBQ+1s84Crn+Hx2MY0uWhR9w3Qe0JlT0kEPZ0DRpdTgQF67NnC/557yvyz5
blO3s7/5XDd9XQrjqYn0j1bY2+xdjg2IycDv+fHqAn0k8wyk8ouZoAqKImfFUhXk
25mhFRgmHAQOioGUwNE8l1Km0rfl8drAD9/WHMfCyLZnkN9XM1eS3GfF7/sB6ufk
vJ/f8CrBhrDjLfdB5rBCey7CL9CVQBiIRDJY6uWPrAyuDiA1UC1zfp99cojZETTc
75Kv8fpyHDPR5aHuA4jasslfCs/FfWVD+Y/DrJ5bEoMpRoQLPyXxEhSRh+ghXIF2
RlVmAR5oKE1fLzShvBaS5AANqqg/+6EdD8z9WtgXfnQfzhskja+vDotY39zEg2rY
+m/vOATQlic7+8Qx8pUrZkx4Og6lwVQW862Vi6D2g1X5oJ4TseTcZC+5QZ7NY4mq
8Izq9/UDw6ord6oCPfH9GcYFMmT3W5xQAUE8nBnvesZbmXNiQ4mppfWF2fS3/yhJ
TfU3FDCF+M10JYn1JyhJ2Ri9ZV5CMY0jqXP3sM269jBF7Tg3aQUfSzp32voKyCNE
hEhpiHbETqAisRQrZh8/PGUOH2bFB9jJ+W5LDNTV+JoiQHrcOXiXURvvF1ANVp9A
7JBQt+AzRixnXhkSZF1GxQ6VsSWYFuN5eqQsN96+GQEInwefVpON2LhApXxVx/tN
H+JoF/231T89vXxCtS/198hAKXJPVcml4SH1CxrMyu8FMnDcoOq4G4pF04oqfYt5
6nzS0QDzt7JdSD2vsC24XQdHpHoD5KD3+I0cQb/0FIgpclMQ8C8Ab7AGhmvZRlMU
rrBSmf5ClViGcxbPuXpbKl/GQyLTkOiQffbQANsP1d1xUzfATCsgXH43h0WUBjIM
kmKdU/vrDB6jn/QA4xwXSV0tjw8b+sd9Up7PgFkFcmptT9ocQZwGJ3j2eGY4p0o1
6wlOScfybdMsKmxZCUy2wbuo2bYPI6sgNmbb2Z0ag8o6hGt5Vo5QVn38+YHpr4TS
ZuRolJ0u0ZKbv3qIc+wG/cwncRjIjjKUxnoxJf1ZbNpRHQWhBXSzeDIAQPTOQyXJ
ibvuZCgohOkoHCG2jPimQqLbB2rsmfzC6ZxkTRGI8k2/+67ziJRLokvhiXmwZtpL
91reAv21vW9BDkdfIS5JER/mU5LNPrcPqxp57fUK6I3r0UA5BhTlA+iir3uZ6NzX
DEJG9ABWEjoASCegK1ILgIZsy+orMcAQJ1uJq4C4x+r24VgFUFWxR3/EijoU5VOO
4HcTOndmjpTK6GG/Z1zM5YCL8dc9B37OiuE2THI7/Y6Z1fjks7qr5V5PPwFqqEnm
I56rVUSPHCIqrWYIl2J+OFjGuE3L0x0PNVnBzoK2MwW2UdQq4hsQzRpH7Gk6+p/T
Vw7/os6VYCFZYmfaE7LWPNWjtGBcnmshqpOMTzPpw68dIZrBwc2VS9+JVl2HiSq2
npBjoVv3i57/oAQKKkIlVqd+G1S0ZJdxap3bcBzLXEwXgD74DudPoyeHgWVjIt3o
a5NH6S1v8OXXCXZvnl7LTAt+celt6fPFdI3gNVMtE+O0kE2eb4pPk1MJ9gwm8A0+
r+IXSGK/r4HbtY304Lwgkab3iPXwHKBT+cMD5o3HSS6/tCmV7q5MaSJDdXbL80ee
O+EPkvPCZJ6wrxdNYR6x1NSXJarm/hdJ3KnfkkMWx0Y5uN6qr65nNGqbjTOHXhzm
R6nTRoMGoFn4WNLWwYDWUvgcqPSU6PwgcPHqo+OINtOSY66fCtgUsVImBaNt0kNo
jDm75A5DqwSCwYAaueHcPSD8UgCSFZzMH2IGqf6aFyk4HCiuJB7gILczZn1RSgSI
87uRV/0JXJpQqdVCVk19PWOaH8kVnZiCx5x950LH4Ftahb+S6TmEYzsNOljVnJl5
okAVH3XSUzXwlhsKXM9xx3yKYA/gZr4dCVMrdOQeCcjkEJNecXs2d53iKDw0Lkh4
VGCRZuhh7cPvjnAK07OB1FDZNZPtulyDvfLCfkw1/QJQQrEDrHXDJ7xPlBiDrt4N
zuq88jkiPKdQ4zOOxWXc7Cj56O44+Ci/RKnNtouaY1Yh9HrBAUtAzDf2a1hyX8Sq
gg6SiLnNY99FoH36AoGl8Vp5XwqMv1vD9P2/LPYIH5faqwRnxm95PBDMlMEdggUN
FKZ9DVL9iwvlhmAH75cG1neEgvaDdCv/GHAjeOxssKW0NcMAGWzvk/Zso8uTFrYJ
zgfvZXbgcRLSZ3Y6DYnhAd9wQs0cgjpeEC6mS3u3unECxj8udV0juBWmbr7b0Mm1
7EThstnyxCB2fqkQLYx7oZvDCZVtx9H73W9K40sA6IV41Su6hnt8xg8jJ8/9Iffs
cA0HY2zVKsxbWsYncG9owzISF1ZWbRT3OBi9p7lzel/4Hi7nhxqP0SC7Dxqd9l2A
qcWshUiFLpRnIZ44nBNshE5pFtJymO1Ei6veJeaV3+Mm9pnOL/5vlB9bR303qtTt
aOKjUek4WHGnD6YI/9tKk9GahwYUhQDzxb9g0ndZ1kHi9jD87D+yBySVFI+pGKIa
j1FO8OmDOpMqlj7sz/4hl4hr98ZbHPvSEa0sX8Sy4t9Nxhr5xW1vwkr4GNtAdoYg
QpdPVU9tQSMGp0aVUk1KYJwuNWJWPW3j8rSipmwfdpxZ70oHhl00Ps3RctmaKPrD
T3zg7c4DEvAmMMzNO17yy0FqrV1M/ijM5qlDyHyxzJ0eOhRZQMYK7xvlBz3dCDcX
gAi9iABmNGpzZDoFshWbZHvDJTsqKUPqUN/ZGtzjr3qQH3fuH4l6TgYhwNDeabvB
RWOOO6dspDFlFAbp3cSBOqsnTlLXIitw7jkVKSJpjVe7VtY9JIovjcO+7ykRdg2O
Q9twuIU7K2uhIxpx8SsMloLiaGyOgY/xviS/mcPYbA9lNLdnXhI2xTShtmmYh1Du
sEcZkCgNk7ZBPFrnQZLLwNoXqCmlEKGLloxsLi0JOcKztwyzkItvGxQDLh5qcfl/
ko+rf3W8QzJ22Tx93jo8SL1bezg08bhF05R8wjvQdTtwGEqxTTwBXmdpUKYoQE9P
K/ds/P+tVIvXAgxe1AKVW3hVmSCYxQHh/WHMjzZC8cZ/ID1YVoJTxZnSD7mJINPs
9GgdDMls9X4ET2gcOevo6o/pt/lImj4IYjCXeMAz4I5FTiAU1IX6N8/0MADaIRPY
pNzhWuBLFfzbUqi+OoxdNaIFQ4BW/e6+U6XHh5vuNZtNbSK2A+zo69BBshXvH4xF
1Da+YK0YT8cHO0sSH+KNLRAyFr49yy9qhM8xT0s/wVAveWDN34n0vfa8/8bpLGf7
g8vN76/VdmJQmaG5hQ9G2utFoZWlEx4tfeEsXQdAn1cRsUi1zEnSpnNnh+5rxX8h
8a1q1VJ9iDxt8oxtGUMVCWnWykCODpWcYyqfFgMlTQIh/4NecOZ1OUftxhtdyCZx
QYE9rifVANysj6GAou2C8jcomVu8SWFAYR2CUJ96LEIcyBLt9Oh8KDYEvnF9BSQM
bKiyJjhqKzeEqHkUKhzEYoKKd4sxCk/bRJsi+U8TqsyWsssLsZ6LxkI6khvttDt+
tNQrEwy/9XLRHW+HL9t5Z15DjyN9ovX4ahXhO9emd5NmpGnx2VmjT+z+73hIdT9T
bAm47wYLgYkrenDsqgC8pC3T/1A2lm1q8yl4qtQxytidrx5Tj9AgJo3c0wlGpchD
Ep3FOOw6NLwDN7Tk5SNB0oL0ub4bchTI5aUG/4QUJlF7cTT3dD+Jp+dslVtQanvZ
iuc4mfGC/nmUXiOZW7BIQx0IoEcc/sEZ+R7XYnhndUX2SWFKeuX5+xqZzy9XaqDR
HoxRCXU5RDdxqTVDmLcFA0mGykjUQjdqNBhFWUw+e1fmhsnI+ImOQ5vlZDvXOOUr
7co5KY4xvTSDmQbO7TfxJo8LXeVkEnRdGJvGPpSLmYgEeAoBrbgGclj9xACyBTXa
HW2FhkPrIKR76RGBHlwy97BWmRIaK2yECHfELjtD0YChVY254glhhXAJbNpbZhZG
x7nETu76rsVR9GBVuFJx9ySfu6KaiIE1r0cey8K07XJ7pfCoQgg46QrDXOO9b5lL
JWqTnuBVe/MGLDO8xogM3E1msBlZ1g0DmltsVHJXcmwnkDbjAWtbw8aucz/mZbPL
sDQH1DnzWZqb4PxgA1DeY5avnJuT+hIf0tAW9sv1D/vUuVAB3fYQzRT08rI+H6p6
XE3aP6FPEeZC9ihPofIOJFgYuA0Y+EE9LUnGcXORuZEWEk48RyBu/SYGBlNWYmqW
luBIauwW96x2XLJHJvBtNnoNw83HDmFxalB1ZE7OCp2wbDGBKjsHRgYXBmPvZ0uI
toox1JTJB6ufiCr5sApfegjdS0nccqJuTX8m208jtLkGM22YRZAyYasgoGWGsUmc
o8tVKI3Dos5oBFOO7C8ZnMM+nKUGcFu22DhkQcVbtERnn7CJCFHn7jRqvfU09yRQ
nLYRa8rxm8yo5hslA59bIk8palv1gUMhUdsmwCP/cexx8dYXo63CM2CTa7LLKw+T
Luvn0mmA83r/c7kdeJdMH7tDlMWTVW2gLIN8XH7vk8n1kzIw5q5LqAgaEKAd6WEL
DEklIzFoPeZorL0FVN+IttQnfIHOJjA4H1t6rIdJHiszuvtmm+J0mTp4ic5eJ+6F
7v1038rlzpgZ2+1tqbAx7fVKCX/qAp4iX1CF5/SYLGDwXW6maIRLb8sp854SgIxV
FDOh8gr1kkn5XzaqoMXGQvxUSxAP3xk2znQmcOCyIRtJYp+ZO+HvbmjmOjaPvg6x
tX0Yi8GYy3AIKf99xIbY9OjAZ5T7K/ROddEZT153W2yobZrm+aGIgESEus2MU7v8
u9XnKryuXejXclzUWDF35Qa77cWLDQBMjKv5fB7sCgYXjUeuH1wnzrktbuV6LCxt
PxScFXv09V4rwNqASm7nq6Ug2nMV71a/kJaZCxZtyKNa4VkuZVNUiGQ4XVQT5dYz
G+1ZHFu4aZFdZoBj/6Y0pEzAiQ/yMFQ9+B5GBJO73Rzv9Pqk9jzuGJWs2vA7L4DP
dpdAHtPC2YN6TEomxUODqXH5FiNqGgYnoi/d/Kj460l0jOcgLgXoJE3+aWfFmhGi
H7ihUEeGVwvx/196AKsfzaSyhmpDrddCMaDyJ6z+cpyD/gSr4v2J5E6bToh9PvpN
HvsGNpPgsmRosMD18p90+v+Ut+8CJgs6d81JBk4MCixQHTp+yCTGpeb9hMXPmfI8
9IGV4+qv5H5dzEUt5bI0UIR+22/lgOzq9L/Ki33qhCe3d4+E/OfaWTmXNy5yvPcw
/dsVNNEXEXsf6CUBK3bAZvjuEEcbKHH/ki93jYDMPXG0kgGJLJNLr1/oVg1BE1MB
NhVIpWV44meTgHUP4pjaU9UWJUeQK5xdCdwpXIxSfKpiG0tgqdQy7HgSXw1oUHua
uGfg517rldPAUwDznriT7C1djYXK0GdvtdngR6ygD4oKQL2X1gRSZvpMhy0vQq3H
t/xMYpnLG60k33hdC4ucmU0mwvxzEpfTJxP8ar+pVUXDMHDBLmolKU9cmFT0RDSc
plEDEFG0HWaraYxOZENv67TifJVo7tSKZhojWjVK7J2opjFC2MGKJsHoaTpnpD9j
FMYNCdfVCcU2zGZGkgvu1b6icV5T4BE4HbtPqSF/ZVcEo+5Gh86AG7szIchnHBzw
fa2gOb3a6F6bkuVkH32JfjvFUvusMtFXSxJClNoXS3vnQPYW+lY1i1YZIlFCmZhJ
LeRBZ+Z5nfF6MUKhXfczJRK52R1uAPNAuy1+QXw6OmZvZ1dq6JLjv50xITPKrXL2
E2VfdC3aJ4Nz+OcGJ3n93lyJhiNL5fwEQcB5CNmHketjB7RaxgtXZ2viGKGIg66b
Eq3orYZocDwjGTWpAvbZI/GgKFQQbbFxdZ8ilZBYee6Caaa2+wx5g7lPOL1CfdOo
TMwmcWe/fpQuINxw3IOmm91TpBZw/xtD4D4S4o82EXpGKn0GwVR1nS5ohaMljsrn
D2CAT6hxuFF1KdxMRPIx8kv1zndMH//4fv19kAuZLLLXjaiE6oGcyVrjAeuJJ7gP
fhC40qOlI8yxwyAy+kT9YDwIhtmifC1nH6F1QWLjcba6txb15yTAuj/WsA6PEqDj
lGb1RpGCk5mdv055vLY4+lMHZyuCbBXK3cxpkjXtjkrOg1KWKLtYYvgzQSEcxzQE
zzOl6dNJKsl0YXhPmB4w8RE1Y/C04CRUB++wrXfaNEnmtwBuHiositedi+eFN0GR
27P32yEtat1iWh6FBQjK37frVSuN7bMO2TEzO6cby+7Akc6h4JiMOXVMOxLGzEsB
Ph/zIkWdZutTZ/QBLBkA92z+d70rJ/kSPPABM9fpNMS4LiKXibdSdV3dMmjNmz5H
nIf9TYvMWA7WBt1vX08iMjlhLi0CDBVmWNhH/U/Hg5cQJRetQ9z4ci+lKYnmd2ni
8preCX5xAj869p7HQ2C9HrLRe3VAW+KeWnI9BAr8+CsiDx0BFwWSDNIkvWU3eTYC
gj/RpxjsHE5GhSpYQbvMyjnlvbenLVeVX9kUqAPPProcFK+fEGW+FiPz/vIsmRCW
Ii+FKLReSa+TxTStTu3QKELu23AiZ9qo+g1n78KCGbfqdRPrn/kmJI7XBKJgWF41
HUqup0wKMCz3+8oBiwkJzXrGxdm6/iZAp3W19v9T3Xp2MqWow4nRk8HZkBCTPoA9
z2XG0ey5zsVmGKB/r5mUaBR8Eyjcohp3Cc57jsTWPdbx0Kb5F/4YCu8UTJ6iXCZo
sgVxvL7A3I9PhJF4JCvEg1seGI5xt0iSdpOSJuvbBxTpUS+aGCW4Bs3aZtRQFKUd
rdh5sIhgwfaX1ccqM3oHRqpzLKDZD0gzLVR1+26SK7I8i55YXiRH8FatWJHJlVck
7Oxy2QD9teRtzhUw76BNY1mv9ulKNL8KzfwWX9nT1gA9nCzzMFXFMh+ADLegrgFo
ySa9uYKyPb+1E2Huuq9iis3fEZPEni8btX9BA4a/bgUhU57v3sFnMtOdqIxt87Nb
ejqCYKZfbgyBqgrWVtrgkOQT167hvtCHgZ0fwi1e4/fDuzJd2mcrtfCCMgjCD4r3
mGsQJMMk7BdQRpfhXpdIAQHAWh4N9knwocPRfMApgKSD2Orv94SZ1nhsNucb14Ki
kQjzJA3ZQ3cQxDM0KqEtRwAH/eKebhODOTI+gQ1AK70AL/YjoXILke1s6EkOG0h2
0Cz2a288ZMAr95FuQDN4MMHXO/hVIK55gwuvB7GmvUXSD3I+4cXqCNP8dCh2YfRX
+hjVZ4NrbTNRU8zmA7tlALIl8gGL1HCi5gsZ3jBdTyJolz5GRjr3Ngx4KFvCPN1u
XLlpP8JwTNRxzynKJK09dsFf1gaThSNHQINQL9kcrd3xtGoYrcNTrpVHniADso8R
H5uz7cwpaY4GhIl12TGxBHsjQhgrHo7pMC96+pHtzSiCyuxIJV7LPZabnZZH7waK
Zc2Xrumj0ni29X2anb7HO26LEZfq5UgDIBsMy1lgOy0wlW1H+NkFybsaRkonmV/V
0kI8XDrYKHgufzxSZY/rW6LXcRmPU8f4pYyXR8nF9q//4VnsIENzT7UKGMzkaYNS
ErphZu+VaYf6fAWslRQ33MbQNa/qSOVNQ5INtJhUWU2PLv4tojCajpKvtpvVr0Go
7p2w8hF8ofHtjn4u9YG1daePSSGopHcgzqctJNHdVBzIwsTSWYHjT21geUiQS/uU
PNeHX2Tsc4dI9MZfntTZcAalNLRx+zEi5D4hvGeRyYpcLlDj58Lpz8zVrNGFeDBP
C6U1F30M36wlFIFVvhf9Pn1ZwjbwJk2q0lrlyxE1Q7WURdSBnbwZuowsE9gKrBBg
wBuqRfphIMY0qM/LDiS5xqD72EqDN6emOlM4edssAM91oC19XkIyZw/lTzpB1Cvi
`protect END_PROTECTED
