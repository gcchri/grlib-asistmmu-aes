`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C7cp0J6SVzwvtjCu0vJb3ayspORUe3cwdyDdyMtBkx3cBMkR+hllofddZmEjd+k2
sBVCmpqBexr6UE3oZXaoeegPVLVfa1aKK4crVes4IWmNn/mWWeWWE26RCRR1GOny
RDKGpFsF1IGBq0RF0YiKjwYwhcUSJuIGadmK6ECSwo9hCFXSApeE7XrVgG/+BYTp
KGhq1yowI9X4/IGe7ragy0775WyFXZoU1/wGG4GIj76n5QWU+RWARyih5froXTEN
uei+qbKmj4TPJiblO9HPZeII0K83h6BSRuoVqrdINiOnAIxiw15ymy2pOgcGSb0w
CPbLrSD4/ntUFJoDW0W/0P5iFm5X+zi+lEG3ZsBc32XBHcmFHW+iLjZnlvAFc/LG
ckBCAyxvmr3FbNpVae2wINhuLDskJPrFaJPk1Seyj15221WhTiv7qZq5qe9y2e9D
VUatnJoZ5cthtx7K6oqHHOm5kqBOjqv1Zms5QEeTIxP1FaZlzDGOvl6PBoDQRjlt
1RZO5OxO0uIRPYe5pHHTbVKsKCtnlLIkWi7UeuJCK4AcqiCiVB8ZZIRu3TKP3/dL
7o9qt4UfoUadgkTOGTKCXw==
`protect END_PROTECTED
