`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
goFTbYi9SEp+IMdgRUEOW2AxVI8ANLJxjm3CLKlbwe3c0ZnFvkUYOQ6ulWLs6XGZ
YfJ6b4/1RE3ihAKu+SH8/0hJDGTn238hrsfSRKJjee002GAV9mxbPZ159EaAbiW3
H2B5zXNLIgKut0hkKy/jYCl8inowk+eVhjPHqtby66p4Sd3s3YAmIyOZ2lNaBxUd
KTZ9uGBi152gljBdcSOLgZtFz+PsNIruzVsezYhuKwtGZDBXwIKsdnZec2bKuYzQ
ZcZ/zJcOzLXn3I0Ea1C8YXwvwRmaPhbhQIdclpoTx+uJ2QD3JGFGMQf39zokt2a1
rbK8axJkb+UKme8AMY0yFA==
`protect END_PROTECTED
