`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5JwymO6+Toh8rhBKPtDWukWZ+/W/bDwyn1ol112ndzrurMn/4a4i+1eeAA16MLb
yXgyiEweuyWNSrhUqL0nKH22AlZoAQFPnRW/DVpcY34BLOd5DksvtnfhpAvpOFv/
JAkiZ8PBNeCWa8PaD/HoToQDRXgweWFN63PvF3/q0RxmS5VRgszCiDsF1nL9mutt
oH7dSO2l40H3sUTaK5mYfbRd0Blm6cIQf0vpgxqNFyvhPcA8BRlP/bJuc23zmKYz
k1xDbSJyCFo9tOLxP3/Iz7f3/xInVK+zPyCOayHMfFFZI2M/hvxlFFkHBk3sr9Cz
WlLGU3/XoXm+8uVRi1IClAHRIKLLzJS+52V+DTmXbznJfuXoD8fIEfZzRo0/CbmM
ZSII6bxIniDM1WOBU2VaiypjfBDr4bcpCejXRvrEVOkc58eyqiJvJqV2GwWatjwo
+9reMjO029YU+qt7zebahI+K2ez75PJcsdzZIpZe5a/cGahlk809naBp/vkFv6EV
jLmiTuHnOxqOvTOCjvhH2EjrGvkO9pVebXCP/2XgwcRNgIUluT7fq2TbdRYWSosT
skyHJdEwOb50GjMNLFNrejw4cmUvZHK2R4iG5g+kl/PsXsUjlH5mPc1Ae0K63GaI
i9ZzT7qw1lEpFJ608H9hT2pEmanUks+4FdUA0v0xoIe8hXnlFyJeyYheAnMnUDKw
`protect END_PROTECTED
