`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iVWi6mJn5UZ+f8kZBOEnofe0GHe3CjTpby9t7tepB6P9YO8c3r9XZhrPfYyZ7qwm
bDBAJttGtCPwvPkTDJ9fbzEjpyM4ZQ7QylBiITQzHFEa2+U3LotYtH1J4Pn/+zdp
tpbU6sjnsZmCWmGfuSLyVJzqZtOvt2JDHdDdWoMs8dMTMK9bfiA2Q7/tYt7VZu/+
lXy0hOtJCfYDmcUxlWcYVxAWlengwOvtq8zrbo3Cp0rE10XCF54pewlv8dB8XDab
CGCpih0/het8aXI2CFfuCaSESBCaGgoTJvg4rcl3l3Ih74zhmx9cbc/hCNboK2EH
tJPXBVw7wRFrUPIdkNJo/LcQxWG9xEreDqS4Iq5Doozbw/B+aYS+GjAvp71cKZ8Q
m8xAcwHizSi2kNEY3UNCgO0i2pZHGbhwNrKtijHNZaDgzXjMSQKhCDtnXCwX2Quo
`protect END_PROTECTED
