`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DChOeChBesnPXHRthKC/8CklLc7w1zPmwrMnol2B6rIv3mLNm1cE5/0AZow9K2cE
C7DNHH7ob6J2dLn5xOLM/sc67ZBSj3O846ggu0TR1fXewY4EI4FyjsvmNaycJlEx
aAapc32tYenP1vAdr9MrOBh/zm5NmJOJzRYgSKs+CvicW/hNaVdFR50Y0pSTegdV
feQbJibJoV13i1p11OCVMty1ndNbjlzz93rjzw2Yi4sD8Vqx6oY4+0y7E2sajchR
/U+vyGNun7dhCpYBco6XZhkKTP/D1CyK/pEYGjpa/kvYV9r0odVfup83HqQ/X8Ea
`protect END_PROTECTED
