`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uPHSdZNX6K6i01uKR5YmxUz1c3ZyYct4V+mPvekIEsdzpoz6/a2UWrInYg7ySmdI
79ZEw+CSKe+Z70q/xDwDzCZAvvfCa7s/mTS5L8wQJe+zJoEyY4EGN//ixNQhm7YC
yzRFhqosK2Ks6NycEgXrPYIDlldkAYh/0D8Xtqw8qwf1fqS5VHDtczF6mMahiRta
Co37EZLgQ1tO/K0UBWWZhvRM6rr3j9Ec2RGI8BlGtGIMpidVQvcKpszpToYdDmUu
yqLMajbDUxYBU7Lq01//ZEvSSUlGfMbBTjNBW2Jyx2t0XxlAyNfDSGH2pMqF/VyD
`protect END_PROTECTED
