`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3B2Ucu6kxCaQRgjKf1W/5E1HN6yovhcyfRTAJ3rV9QeaYPAe1SotzauN3otXH58
CHNMlPND8w4gnXHOIl+7UDlFNS985hVExjzJfemIeBGuX40DRn51VJSFCkLqGsVY
gu8BlCCZsbZsisC9rH+CbTaz/3Z8Y70N/W2o7YOpU3cpskMUU4JSxIcoCgjKEg3y
iv6WdWB4v0FCWEiahFX5d/ORSYua2vojcIfAO9ALPXhqAfoOMq+yuVRje8nbu+Ar
LXQ2gWOuLj7tlfOGYF8IW1+7K6q0tN1ajyescGQzZvM1uhuUZMBCJs8FeSGuPy8n
c1xH1xxPpwinvO1YAhQlGzQLS40/qgdivfcR6uJxCdI8t+8ID+bFbXyNmjvQeTEZ
QCuIf7+pHsz5PcdPTMz9VlYdE9PjWNMTIdTTPsfNfQEcApPFfFK7gdrV1Au+wEM0
sr8i0/YALyBxBds3UXWrDrHiMoe6TJRm9s4HmkxVxmof4gE/wLFsp9A/7MtQBJwW
3/HoKgIwHL1kHoyGoo3uz/zaj7GJTumqfOuwKOv0TKk5fBAu52x9LyNvTOBZeX8Q
kkdj0v8Dm9ITHcyDFykmUA==
`protect END_PROTECTED
