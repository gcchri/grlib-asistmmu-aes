`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCXet/KcgWeo5VX7YR3wVrfU2Wx8T8GUmqJJS4Jzwrs0Vkg5STMfhjrFvDGzoK3d
Fqm3879RpMa/Uvbj0i8m5X3oB0MZjK6LqU5eQELlAfx4Rjme2rb1dnnQIcdYWYYS
amWPxdwcuo1JSD3EfZZuydC3a7l/khOK2DZABSHA6cmO6kBXSsyfRBkqpozLmsbv
2CtjpMLqqBND1wDJmToW6ArKzKq9H+PGElW1p3FZAcD+s0CngqY5cL23xNJX8sFQ
pcW5QcqvJmRRA5FKtbWk3qO5/CsnXtAkrAF3j1/h+T1RUeqa22KDKWrdlqENcF2i
x9PLhIt5BQmIVzp22Kq/nFsD1iPjdBo3Po27lrOx6jEUS3sFUJuLDIJsN2FUq10z
nKR1oyMuQyItfGAyyDKk/lwWsyJjgGl5BFgpxq8qBO8NGXutHsaTGIfp1maaLnP7
jP8M2wLIopxOS9FcL0w9dJmO2P+JC2rOBQXRbMBLlo3ppshe+7qAui8t+omB7Pp3
4f+o1dI2suDL0GPLM2reKqThU6XHHNSMyTbvH7dmMjTfQLAoh7OxyRJkpR/6aJBJ
tDNjwIbVKME2ho173xkpR2O6v/c+ooABM0GzYrzDIQAvDRThjIsoysJysogbSVAl
qdCaGWJtuccjoFsQQfFK2aAAI8IhG8v2GZF+LJGxRREy3An7zwmCp74/y0e2NYn2
HIj8dDs+uQtF3WsaShUxgl9Q0lmtN/pjnkUkq5iBtExlIKJZOWZk7OXopYR1i3Hn
kntQZeAm13FXnIh9U2lJWqmzt9tO2z7kErTdbonfe+38O05akYyM4a0wRg0dGzNV
`protect END_PROTECTED
