`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeHw5mv3bZPEx02fuVEUu3zOXEUqR8jyUjhScp7oxxS9q/Rip7Gn/S+eOMnHl1g3
c1LRn1p9QWjWWLPRe33LzEfN8Bzdu0s5m4mmqkD/9/cPuyCXStmYXMQw5JdVjODZ
braryNRk34S56sYS2u13Qdz3tHHs03MFabzntmwNLa8OevAmnyDz4Eq3ZQfAcLuN
SDZduFzgMXYVRk/BcHCkHpV2l0a/NY7hkZXY62Xx09uX3nhuwArVfn1XLwDdQXDZ
3BApIpMhspcLOYVj7K1hX66bi76b8/2uAP5w8Bq5hfZccz/G9KxVhuRNO2lK8etg
/6bay4ndW/vuJyTnWN6zrtpGd97RATT6blSekP2PhWR8NVCVFKhEmLQR9VMgn8Gp
lPJFpJvUGrNIXwKWj1RHeuuyiNotJ4sM5lu5HiAW23+8RYxeJVdxWAB7ZIBi6EGv
DitN1R7SIgb3YLMTa3/pPgGGlS+M+Kn7FqYK29mWwF+KOt/BFZb8CnSPIfnBDMhg
7O3Fm56c6rw3n8x3Zme8Tqv1DImc4BVrYChf/wZGdaXiCTKzmmA27jilkbhP3Zh8
dx8ylv4iSIu8gdVvoeStdjfhzPO6WU11Sfz7U5Nh7+Bw3ib2+CxQh0JbNOzz8LcZ
/87tvaQDXdzDMiCITCKalNb/MpKXEeKW5GZg0u6tJd62tRjVEfLZwj+jlW0at4E9
n4q7Ln0bjKtM9jy+MHMdxqsAciezbXXoYtsTHGPVVzdzoArVcOvZ/kMsKI5ZXNTR
bkjo3LskKx30NUFw7aUYtTfa8lwM0fM+r8P4VumvKlQ65FZlO6nZPS5d7CZmDGyH
z1fvX8mdPZ+dWTayi5yUJyaGWzas2/UIHqoZEi+tbZMezK7OvhuXok8KJbgch4Jr
s5qAXwg1L+c/E7vMa83gxXFbGybA6xJb6MZpz+xSPAyp343kX2IWAxNo2ENtdPvW
`protect END_PROTECTED
