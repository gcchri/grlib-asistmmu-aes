`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BKdFG3m7DoqcDPmlDYMI8O6TbzjiC/O1gRBw42prZAU1JsSU20e2MuRGZZRCIAQm
9eutQ0RZkAQ7z9JNUouP3sjgDYMXMjdaOU9hbsr9UChWFzOYMqCwUpOTUnj2BsRl
FJNTsKVHdTU6tRR31nLW6msZbzzmqDkerHwVwRJ7FsOpHa/T1rWNt/kPW59rJUKd
EBS4Cj7lZPkoPLLyJFWBG2TeBxyyQoj9SmxtC1H+sznY97IifcxyJE92AFugEwxH
ghGVHsMQLagr0D1+aEuc6GIXJNZeq60AhZNPN2lLJqjmholLC/V66dGIJEQLaewx
qswN89WfjeBzeChQYEwzhGL65XftaR8DGg0INWjSbYUjFI7AzD0ZISODTgnqoSL/
DH9HURK6TDA51vlmyBxOsKXJgPiLCzLpHDCGZpPiWV5T/vS87avEqrWaKlbUBqOc
eY2g5+dib8M8mWGZuqy9+PymCbjY0vMTPoHNwZUiUWC1z7hzI8acj4l/di8NXyNI
TF4P6UbrvXt+JapQvuTFKEe8eb0eFr/40sRyjeuunKYeZfpGxdlLKCL3IPNTveuL
BGFE7P7Kmfn+dABLLbV2k7afLXimRkBFmP95naFFZocrw9TYlmtZyKQ5dww+pXrA
B+wJZV+B9wbh3U5BVQVTd59GOkDJy1W1OF8VGLZU/7o=
`protect END_PROTECTED
