`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jeAoi6JJNhjB5r96ON2UZRj+ZlRIMEq0AmzJumUQzfBRYHmHTqFNW2XolJueeuBI
zKF+9BstWesPmYGLjL1NawQO+hzbqRtq9HCD73cEFuNYRzjY8ZoDtYs+Fdfo39DW
7jy70ZPBfXNRA0ap7UN7QYwde04nJE7g0DJ3EO/duh3V++RUpTIgwoYWMTJ5T9Co
HRDTWAlkr4Nb/fxPccaF4gt7+g4Omyeh/W3gI8EhHnuOJaSs3Wbczny5QnNVVuIs
xjXqNcPZ157BZFe3pacl8NcZqa6Yk5M8WbST4s0vQSL2rW/k4zY1Nfp3cNuXi7nT
tKLoLgUyi/YR1pxMimvuYOIPkalM8Lz8nE4mKFJ+9KdUQn3UW3+hE20fPK5uSkm5
a1V9mu/MI04vFMb9kcxCNzQgsdnet0D7gdjyOnm8HSfjhOqBv7+ADOsvtV3Fp1Wq
e2H6NdrN2UESfRjZh1LL4vymYwpqo9PcO5P90/OlPkm3nzqmJNRSztcQrQMgQtYW
8xKOFiEiplZxGXFAmYMFqsTVs0+TFGeVv1lKIuQfKtxQFEKq26OXQGwRon7ieWSH
CpxGzv8IKBSAowIv3cJFMsJCJk1D0+h/k4e3da467KmrVALlMaIUJTgJ7Skme7Jp
3XtKxPAcaCTbii9wkam8Go63YyXHi5ZJYVfXcxXmjkGQ6hQRBiGxFKolomJc0z50
`protect END_PROTECTED
