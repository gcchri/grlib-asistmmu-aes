`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LL6H1s2PFBXXmL5oDiS3pzq/NIZ4lYWl5cx0JhIDVnA+kvzmFYaYeaqEpsmDx5ie
vl8uMVXM7Xn8oFMss7sX+a3/8F4NF9wn8+qGFec+g2l+JysQ8FrVLmBg/HEbDv+B
UJyypt6dZUrEjHFCpNhQgQoc/TJ0EqUyNvkOZETcrD9gQtdvJK3qsnFXKfg5SZwh
v9auJkP96n8dmKD+d09CmL6oRYCLfQeWRYipMzZq/XT0v3DTXZeUVF1Q+Yt8oaiq
6tXLGin7nYByEVS/S5G7f0G9Qp57V8imQQN2DnC2ICXBTjbUOsRCPKdjbwaPLypE
6Jw4ijpOygNtLEo8W5lb0ribRGx58Zo3jgA37CpS57PycagFDPgs+9IunTTsU1Dp
c87F17e7bjggrsKuMGJbrQ1IsF38C8/MwyXLHxkK2SM=
`protect END_PROTECTED
