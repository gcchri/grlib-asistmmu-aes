`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZgeWogFhmH736V3A4kqLWaNZKqhw7r1EO4JIUgA6JM/Kur3x0Ti0DdARx8a3u/SJ
4Klrz7ZiqaxLPUA10GJz+G3hbl1n5jxsAUb53IWTeA/toEIe3XNtD+ODC1HJLtmQ
NjigyPv8rhTd4LzVOLB5L/SSe1E3WdQefD7aMe3+lyGCyRpK0V8WizU/JIOSuCDE
evqupnn8AOGEblzKZ6HSQjQ5ZlRxCcFJ/O9FrPzzYur4qGz3UloTQ0rFfaWmwfGh
qCyxJygZ28i7ZJ23O+LS62BWVhqLYOBMvKLzN2WP6t1W1KHQECz1tXWeOJ0xxpaP
C/n/R4CoyhkJF5wRvpjl6I2E2FYtPnHLMDOOgUS2TpYjukw6FrsyHI+4OpZVxDMa
ZbcxAwVpj5wf0zu5yPZhK3KC7FyEMAsPBhf7GhLkjXAlaw9RY7mC7ZPYTAHhcNIb
pl/VhvuOiQZ6+j7QF7L25UzMN1L8tRdDa/dR8ylJaIQZOrhdilusJ4xYWuphGV1F
1WepzX9PpCnoNLWCrBTN0rwT6Fn9L3buVFrkhwelp7TeQU6UdiXfN/mxNELLtlUA
EVJLpr+HqDGjGo7A5oSlN+0f1HkcToN8LtAmybL+55ufk+R6B+wyLKVlQSTs2XKo
6OeCfzu2XRR4cYy2KUxzDTElk1dEznF4NoITh5+FOfeFAyV4CImQfeesMvTcg5cg
bsXN5NAAsegB0se6FudHCLihvU1va1/GyMoHZevjrhvRV+vOfVrBsfxKunZuHqyE
PjvoiXwkfjT9B1asJlfATtTX+FWaMz9l/9/zn6cH79GQNMQGMbkq701kAWcS0kJe
kgq9isu3gO2Njhf3YVP7r9tcaXW2+0rPNJrJCRbdlxn/iC4x8R07RocbKjrZ8zjd
ym7zOlA1BAMo1ChqMZ1ipUk2zy8cA0obyyvIh5c8BJCMEWVVu+++6e5cZeSS0slR
3qfPx872mPeJvGe+kkRZbg==
`protect END_PROTECTED
