`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KDcpXFCECVRTfIsAMPNrsajpMmEmnu8L99tPh7L9w7NKIFBkqdbx94en3nxJqAKQ
eqdQy7jzwlJfdl1Ty7CMTYOq6Gp7CbpNdTFAArf50DR1XeyLxyZxrLq4gi7Uw+IS
BaURUmB+JydmsHP4XnFBWmFFNOIOneoQxGR9kWJJvEquKgW+3/PaE1558UjuuqQQ
KEUfPhlqlt5WsLYI2cne/aYEItgQvJPTm2ZtYqAtQFGy7ZNpzrGaAAQY5FMJTw5R
t3ofp1YGvr5ADEsOFRE2PxECKD7vxBgGOSm7u6GPL16N4lhPff8kMHmyrKebET1q
dSes1TOz1/2ijvssz1CBx821J+l7MPg+irc03u7uF5vP+uOteZftNBEfmsrEFlSX
DBBC/tfLBXHvNXO8XnoTSvgDFglQQ29179V2wcQSRlOzyRx1RltsCbeYEFsqj9ws
w6mJ1ShzT/28vzKbCFoG8pxH7oV/ygNf1mZ3outkudBPDFMP9GpFWafTKv7f5fzj
`protect END_PROTECTED
