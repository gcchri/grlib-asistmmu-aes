`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRP//zAz4oMpCuS4IwXKsTzmfqOxIPhmKGPzahKVBq5zfsJWpm7JztSpqNit3/ms
oW+xEn3pR7Efry3Vpfy936Geh/zIvIEiaVRQY44fE9TY9e343qkD2QOdsSsExmqd
ufgcrX+qY1J7VgdTz/IKAl44mQJ3iOOtHJFB9711R9T0pFevxr9eq7az59bPWC3U
5sB8V2PWhi8wcTCF/DpgKnm2QY4XFmM1pVni/KRa0fHT4ay2f5KBoD+nsquaxzjf
dv6aA9x4dZ8p1ahNXII+frLhwo8atfIv7D+8hFuPdCBO1fDPGBN/tqHJ2zq3/co7
lDN3JB9IQLJDrbcxJdRwgtbffcYjwDHtOB/oPZE6YKeNBAdovxmGNlnNAEowNpRz
Ug87TcwW0vLthSW57nBD2S+GD8WzFb6wHvs4Unbnas5geYnjbaWwttPLhZE+oQEr
uJnVeaWh8mgJVqpjtf9+syDEpI/Me65Y93aPT6C7NpPyNmHuS39hbLSoq9CGIfFP
E7gIeGiL+IPbZ4E2QdWYrnctNGh1WewrP21DFY//sXjVOnJg5mHHqBRovr7e0+Jx
NWa/9tqFi+MQb12BnJM3XHWSekiReXGUDL9qve7KeVXMyVEvM3IKS7a6zN8BJPw7
HFoKAKws3sJ30z6zRqe5+XcjY1h/Ulr9DC8XBQVru9iXgtRpECkcwcG3PzkUzvEJ
FfIH0fN4NLD3D+aHCWGmYcrr2GO+WtMd2jsi0xn2R7+mlXFyeax6zSVFkTJUbXpi
Pq3ldqDh6OpGMdWgIUXHyuL4WR5ovvPjQSTcxNGhhIzahz6ba8pthff00tvdFVHA
8qT8JldA2jdbmJ3nqeWolgNK7M5jR1FO5uG9H4QFsk+Rh6MMKtEOCeEBQU62K10C
n420S3QEI1zEutGp/t5aaOPrVZF9ZJhkaArH4CLeGNOQ1wm65hBhNk1wKjSLLVKS
wCRZOeAcGV5krIqA6mtYfTA1fmzaXuP8Z8LjLMV3mRZ27uRRzTzbqMKf6Ia1nb/8
SmDxLTuPHzl+oh6ZBvvk7pS3nnzttxkpZMGoAPiSzdx9UW0kVFRIFxYrVISJiqYU
0r6h0HkGm6guHE3w7HU60C8KUMR7JDEnnKOm/tMfM8uErB4G4LLgvQdUHiL6DnGo
bcDD78lRa0TH8MlbOPihKsTH9QORm9atRN5dmvK2g7xao75Cq3Z0kGg6q8Z6CFCw
DmvhB8qTexp1Osjl04Pb8vQOhhReXjqEHwzg+PcKr3v6P50btfcsThJXePDkVv4K
`protect END_PROTECTED
