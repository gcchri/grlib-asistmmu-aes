`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UVJmNID6C+9/WcvsXNNOX3hUfHAeIuZauhWHrcNGNM9OdkKVjZGhXuq7T1HiEJUb
hVxfQ7800ezLqJ5AoykKt0K2SJFpTSWRWL5Q1NZR8FtHl2ByaS8o2MQPQsTVsiC+
3mfYDa0FTU5CBaiEAESq+Pv435Y5clIke206myTCYtRePY94YF7UkvCL5Ba5r52u
6IkfrlonkXxabidAOnQjfYNOqfVgMq1nOth6B+8hpPrHm8FIXq2LQ982sdaS1wzJ
i5unk4BpkRMDwFZLokA3WnaBHwayciJ8OJdJhr3Ycl6ztMaPkP6K4jpk3rsMO30T
C/2loiw4FVMlJ/N0qgXQGF8MKEJL5U4dwhby02ifu5kUldt1cfM1gAFPmEcYX/Rm
/09wDolSDaPB6AddpSNAn65h5A7Nqsr45sevg1H7BM65EZJx5msuzQ8x2BfjH4vk
vkX+9/BXsbkkLdh8xNYxhZCYzNR2EbVW2LuWX2/0jmzJ+eDv84PUKcB72mM1W3KG
kdJpUsEuYHUz1+3qB3QpXrymNgcNVHb78wQCTqZoLnI1dUPwNI7U7VZwHACRMpSp
orviiEVvnwu8ObFTK04JFFUK/Azygud9HaIkTajWA0uYFqm22F3XD3kwNU5UBi8K
6crB3NQ3OoIda4JljP7xgSkX9eRpEKmmM6vNl5Cy9f0YYVVaKCvOREfSrP0ltjq7
`protect END_PROTECTED
