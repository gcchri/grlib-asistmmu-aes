`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqAOngONXqzZCqqcH+xi/tKlym5Omv6zdJYSn2dGassnmOzOXg3CSd2VWFvr2ywc
Er3moLvAbhz0Hm42XxZXLXaWwaEcFBVk9QZ6AlPTlKvIt18zeS/2lWxn3cvUmm/p
sZyv/qVoC9FkUa6D1Kw9McG4CWIAhlNaZrvDQzTOnpGg93oKpCdyR1awzdLkptC+
CBy0MfsDqAUIErpDpeLucK9bi4sAr7CYI8oNrDqL6hHpdzUE7Ke6xLwwoMy3Myma
UKIPHnF3O/G0K5al/i0NI+WvCXueDTlswxRkbz3r4TW2qZqblh2Kkfs09ckAj/an
SsvnS/aRLxxi4GAOLrW+MIzA1F3mZo5qfGEzrwy5Zwmq5Je43I8234kKe4QVXIBy
GYz7B1uSWi4O2OmgxOKCuyLpaCYP0Ajm2o7rTgSyjycJEgSYzDrkYNWQM5J0wObJ
kTuULH+Oz2L7gYdvuWqvRNchXogBDjnJFfOLUzVtGfNInKl4hK11VqZ5Gng8ycEe
Dgk6T+rVJFI7oKk4/zsKlCJAW/xsVNXmJY9RKBkrX2dbDAeEg+ITEmI1huI9qcwX
2PHcPD5a5GmGZYrfQrifPS0pFyZqqQCUn/Qhn93vZmihFIf1+IE0wijP6QNOvb/8
`protect END_PROTECTED
