`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BtJLI7CIgL9XGKjGzb4jW13rpT8T0pmayxKJuL6E6F2Y9Cd50L5qfbMCamrSzxV6
zWI0GeBeltUKjf8JIqv/LNaQD6wYdgp2fOHrPX9+M0tsvbLDxcXO3XKcQYQlctQd
L/Q6olAh/jM78pPtlIZMm1H3cdnYEouSiFIMHXyWgVcESxdEoJ7jOlLpZasODZwB
TdtuD8kc2trtMeQ/ofDQXI181e+s7yNwkY5eyPAunUSC20wy44VDMk786W9nbnpf
B5RB5fCTq/28GFRpj2BwYFLMHFJrTRV4QdPj589LtHQZ8w2Uos6b/x2qce9Svsi9
hHsuOBDBBvmcLUP3/0C/6PFKoIsvXE3ky4NHa7GcsVXScGU4pIzt5Y94FZ2TseeK
GLqgb52n9ESFgiFoDp7XnlZ6Z2xD63jpORyvw1eWZd5kwYKIep1ZnamlJ1i4Xmqd
KLSLkohn4DytK6j38HNSXtXiDqxsl6BkIqf7eXnir36dye9yitnYes663DYhG9mB
jlBlHHp1h5bWzwAxBFbP3mrO9R34oBgZvGFkImCJSpig+0J0wVKEeNwVyKfMytVH
KWF4mJczKZ7LYUHwQJq+mDKzstaMRbV1iJVFbLiEVesLQyLqdqB5xTDU5vJjGcm4
/U7RcCuSFnLPfUwePiHk5Z6GcjqTaPmy0i0c05Dd17w=
`protect END_PROTECTED
