`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3TYmjQABNCybMfI3sbzBCmDSL8pXSHpwHMuDb/BkIYCBXjrMwfHLuXkc34sHZjGT
miF01oucabvqyXIZsogHsL5GYBi4J8cdD2j9fTWZoDhF2yfkDv0ff5KH9veQkhuk
kzHGD51LMSrbsfNwMgj8ficvfFdMYuBQTrsO8PmeprF/6ByKWiyMgDAmJX3BMz8u
F2TeEMMoUkKPCkqtSxVklSRsJmvpYfl3vz9x29VNGF9wXfdX+oTpqFWJ4gyjkual
zV1gzwmARhMzkMvslYJknm51kTkU2TLM4VcpYAB2s0xVwZIPfKE5ZDYCwejYIu7j
0lvExeAdhBTWxYkb4GTbJopIYIbl3rYnJLmAn6A7jqjIURjTqW7kOYDFnNLvAFoF
QmYgkPQEhilYVVoD7LGQn0tT9se565V8e9CyvJaDEoMLbrgSi7KfCv+S65XMFl+Y
QPhvGxIMpqV1DAY3Z9hmHPKz2HYQMcBORwd39cBQ/KqOWnoDJflTD1waOwE5nmhH
LR3fe7WxJEa9sahpyvrDbz3imtcuXKY0bEktKsYeQHPPsyBQuZQoh0B1m3hbIQVg
i9VGRLh4LV06FN5UhVHoeyacKg8ul+P09TBaORmG3KekR914u/16R1AP6N6mA27v
hbxcxUs/GDuJi+0/BPSxxbo72YF1NDKGi9vJRMFGKCLzzw5UEZR4PY1DbexfIPfM
J/h6P0leHcm5a26+K1Y/+qsKnkW/orgerg1Wcs91OJH/gp216Ua1Uu03sjDpWMYM
xGN5Xr8sP2ZHfMs3oi3YlgJAFAHe8s37o0zzcrhB1ZPvlTFDXCy0KDFy1cr2zUxC
aTycOib+HPo1hx7PouX4kzju8We+k06mpKkcmJl+7leL9guL4XRkTxk7BV8doMsb
cVy9wGKjtDBUCd9cKiy/DH1EhSZteXOijDIJy1u0rwRe9dk6H7XNfcFgIij3+1vt
YDSXtYlgkF8LCalUOFwYUA==
`protect END_PROTECTED
