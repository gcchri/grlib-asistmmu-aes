`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFFwlPzFjx0dEwmoiEkyBrKHwQlJusUN91Y0lB7a03BO5GjYUzbdq7t7P1pGoI/F
4GJ/pviJKV4pBHgcDNe+5vZVT+1Tdh0Spni+baf6+o//56KXEFxf47YhxuNR/7j5
XUaa0QzKhvoTQ3a6sAIjmJSHgw7nbPC8uU+gisMvI+ZlfdqeAqyNECXt+YzzDpjz
T1xODf9SFhvpOcMtpEd58cCt3j6iBlan30UNn3yK/TV1CiYHvuGORfjd84WI4P4Q
OnZRs3ryqhNxs/0OtKCCJpl/eXDWr4znYmoPH237LkP9MagCHTJJ9+KorZzD/QdX
H33q9hdC/nUxsnGoVkxnZDCWKK38JMGRgy+W3ExonBGZbA+xtmR3/IjeURq9Nd5D
s3mGtEf43DewKBngwtb6yC5YABVVau0WUG5TO0+LuUKQUHtV3/lADIPgodaKaAJU
KlNykLrpg7XbV7F/SDtLydom0gDuXTzfQNpFu2e8Y32DYIjLXBYdwryaU7DEF66y
9qWh6MpCKHbPiQ1bjtcT/w/t+ssXXzou+C+DUCKpwubEgI0ElThyQlaHqcmh06h+
rQdR+qxfZTsDMFJ2XpO/hpQkLAV6upFw0fxNSkKbbKBT42G1/PmbNLoHnvGCOkt0
orjZiJPEjnRIpI2gfhGyb4VzgjinQGZOs6Ro4suQ73zv9MNffqjYp2eAU2hMXLzk
`protect END_PROTECTED
