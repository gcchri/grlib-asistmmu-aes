`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MDAvZUemWd4sXAzB2blFk7z6tXYo6bod9OyyAZf5mev6WU8OiVuEDrekbf/stir0
QdlZNJ0nA2p2BG8Yf5cOx+U6dIRpI3qi8x0WzKR8rsolxZHKbgHZ52Wcu9SGmjoC
AXDV6MHpIrEr65ubaZ6A49oyjcoV2uum7KsGjAWFcuWMJZeKQr9h+JPrXMuYNQnq
IaAgCiQjUTAZvmhvN4HOQiWu8Gy9d0FezG/LgE8ja7HB+MWACqlTOXsCIJB/4ys9
lvHIQfUw2YS5GFWUAIr+1kcpJSjbWfatEySs0CCJlCN81D6IcFE2O1u4MCldhD0n
JgMXar0iqX5Q3KN4mDAeCAiOJpdZ1i5nQqHfwbAoLeiTU9EZdUD7ex9WZPGTTYX1
`protect END_PROTECTED
