`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NOjLlc4rnBMp394kg497Pig+RJBVC/iysok+V66KJloTlGyiVeqYeI1fVfUOlIFU
hAvW5OtRpR1mHNTJuwH8Z4UVNuyGIhHZomv1gqhUGmRtr3oFh2cf/ZP4TuV1J5Yk
fWbdXuOeQjCL5H84aBDmfuY3o+XN93AgCMe/i1oV9bOpyscmPhMZJxZZZK0pn4z/
mYlTvPp8XoOIcL5SKgyApmJxo6J6A6VoE0eqEdHUpcF1o4lflQQh0uEN6ZOadjR0
IIOthe6Hx1Ws20PaPTNrNaBJlix23UoTKGu/9ZNeluGTA4n3TRoErMuQp0mRCq/S
Q7Zca79JRfZZpgngURIcZgfp2dpWRQiTaT8ShUrRodrtsnmMJA3tK0jy5slQuf8p
KW/YF2KIyJtMQVWFYUPUIzllEtVIzIx9jFFp0EANVt6ubFL6+lgyeuxRZNOYXNEy
uRp6eSI9FWmRqvp3J/GK0w==
`protect END_PROTECTED
