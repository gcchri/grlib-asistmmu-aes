`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmI7zDRhqHREOVIxgMfP+sd6UoT8l/o/fH7bMFmDYQZLXA4FeTuFWWtBGffGogSL
0RgUDBiwIRmG1K4nzk8i0u0HPdbCcV+gdnKPABb57H1K4bWk5KnEmSwAYLiqZYQx
VC3bULA6tOQkmBxQopS5H6NdgO3ZujnAvwmacHHHtcEOZ439+gu3RUe2+8Lif9bn
rKlJBL4BLAEXP9ah20/Kfq13CX0CRpCcvmub5jheMaidBM4q4xEAWzXcF1+3aktm
9WDWVxv06LW7xvuH3XfNNLxGC696kqcEhgDTLB7PgIYq6Jo+wCSYj6nDtwlshBdM
tcOurU8x9gDbDjHY6i1vAZo406nh+1Vo0LS9gi2mLgeimFgBM42tH6VK74SFvAM/
/c2upzNzoyI4h6w7YAxo08uMp89gEvyh0qjeIz1Nd01IBjI5X9i81p5nK9hKIMh+
bKdm64dvUNrI6xX2/MQ7sGeak8d5yGsNx8BjqZq5797fPfHpZa6PGfzf+XFTGK9I
H/+q4cqi4u868P+RDaK6mqMWV71o9hczBGcrhZ1FsqP7fKyBtNAkuYefXkeczUIr
4DB0oESoz+OEdJkMMMwPOLo18xQ7HPfdry45QexiqFdXueMjfbLqiidoEhlpOTFJ
uTPq5VUbfJ0Oa5B1M1NJs5UTW/9tjBwgwYvA/BOS5zFgkTxQPjcfhhq7Ak2zRvVS
xexaJ4IXaKGu2XC+VEbtgg==
`protect END_PROTECTED
