`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9NM/YYeEn2UkzndEcDiBhsmGQE8nU329j4dfblV2PnmBaoXs0WmrwHt/zmyzQSsu
3LLyZws6SHIK+0sNn5NT6u0XYlVVFV1MbFvjGDcB2qI7fZnFMyQqsxSmj58fElHJ
MN+iZaF1yN6DYP2ShOxOL8W5O7m8bg1I+ZAfvJKxJ5f2EJNX9PXociWrimbXCAWA
YJ/M/iRQccxX3BKiDOPbBSAkPk1v0aZv8Hr9v+brkuP2/YF2YcCwOFWzEXS3KfuL
zbHXMFr8p1XpjG0NEEExygXTbypUV0xWTUQovoP3vZSQlefxnIIHDZypjMOQCZ4w
iiu+A2nOu2w32bXb7VgDG0sehgmc1qrDuqFsNYmT8vLIjt/TtQLEeFDmjx0gbdPk
p52nn9WURfrGUzqktDfw2MLGItSZiQbMzB/hWr/CKOYKxIC9vkhokjCpKTu+sXUV
nb4z0Jpt++DNNoGA4jdQREJW2AfiNVGZewUXHrqJFi89q0c+Yp8nmLatLdud4tK7
RRpnqEZE7PsaYvFLbxMuU73maMJaYJUOUF6HiggICmg=
`protect END_PROTECTED
