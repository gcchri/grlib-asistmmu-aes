`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DH+Ps6f0BGY45HATEbApPIlncdFiLchFAAXtkwJ7NIegpGEXW8e0grNHRHPgpwbq
5l6B/BIRzuJZ3QB2so1KWktZVD1bYWqmrO5ILKqgc4siDbB3D0iJMXN7IshoRSRn
LkwXKCVxko8Qcu7PJCfqdhYDM5D9VT90VM+pZufM5+lD2/YB9tIfoF8vkjHQRiaq
6UkxiEfNbe42cLhKUvUnZCtje4XLFlxFo5RJa2ag2ytmI1dLT4B3n+NoCusqnJ0X
DEuiW6VHanc30pRJRikaISic5b8A2SNcZTJlwbcQMCYyalGn0uRqy0fHj0r8Kspg
DrmR05yXq1jO7kwDV4s5OE1ZapnBiu7m/OB3qWhjpfjDXdSwR5qsYljbAGzRlV8s
8iP8tjc7FTXb/agVS54wbMQdz0C+SMZgVzy3sgm7RXPCqBh9EPe4eKpoAInzv72x
TYi0WUiA2FiNCwa1rQ2Raf9ijA4nKMQj9cctDMM+FE4Zo713y3h8+QRt733SSvUL
mFdFTK3DEjLegckKw17nIoBfL4j6tpO6rzUafQSaIKeraERMcnd5WZ0ZQe5uzt17
dqb/dOqSM9bznFDwJkGs2uLrL7JGMXqSdY51uauUatZ8sm1AmSEW69o23+2MJQuu
QbQ47eVLFGUl5fseo7mopPqbyCcnFYIv+PomYe+3WhbN7XoUfpyc/Fv1S5INUiHy
TRZ34QYhg2q0yPBVeXn43KpoKFzqs4eJ9+YDf6GV451oGPo0fjnfpXsxcf66srnO
ccNyZOZENy4xv9nwQoHddQ==
`protect END_PROTECTED
