`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DD12nilQAbTGyTHow7WHBl9ztN64Wvyc2Cn9L1nqJt0CK0/zEYI/lO4i+fs3MS/0
Sz0mxi81c0fZqptLIpvVW+nLam1BbF3UmafJBU4jRk3XBbDdmsK4mTR+M/Q/2Rac
R+WYA21iLFCPe8GfW3Pk+snMZq2hwPgmFtm8SSPohkobGt2gPMtLaVBiMtIq9wue
Yt1fLqleqElcS3UbOXySOnl9w3pyXGL9GQOhGxpgtbDOg8KeNHQiHkTyK/HsUITU
hfDnVLu3JWBB6pSZ2nZ8Lk3Ky9ra9Iwh93BXLY2NXFayndBMLP5QQU1/HLiMg7Js
mBMNsL1oJYGdiNnfriRKejQ8RTAFke6drYl3FDLLdMyTu8zK3EbHX0ZNHOwQ/4jv
/XaG7VM0wDNFC859wmnb1MryJTnO4dO4/ySCPEIO6+YSo2813PGZ7uFmkx86gYYB
z7Gy2smhrEoD4lTRQL7s/3IiAfK59kfrYC4iv/vArQrfVOqVbUYEtfYecSaFI8Nr
3fCH1ZimlLaIkxRdaJz5hK26opNKUX1yz3R/xPg0VIHiNs0v6pIut65tSCtdkFNS
zNc0hwcoYpnm7ZyQyUKgD/5UeLDbwzqTHpdpZ6dwq7pYOpngbx0Z52SdaWt+Nzhe
0NnRo3nWA0ffYtha7YBfVz3FbYnEnBl4T6a6yy17jqjRA9SnejZCHvokconRWKVU
FV6EpjO0AiTvM2wIfpeqxLS7Rkuxm5DqgZFjsL1E2L3BadPVZiBXDr5xbjiiYib+
66kMOZG4KuPc7BvraP0X2od511vhJ+mGQd1W9A2s/ARpboXZ3cv205o5Cvs+zM3u
+VgLg5T1WEw217XvIHR9w4IKPFOyD4ioPgc12vPoNOpWubkhZIesnBpNTOsl8o6I
FKWQ5yV67M396akSA4r5jKNnpxOhiHGH4WtTkclX7Fa35X9qTztVS3pVrvIi4is/
9SXO0TWf4S348ZfRS7ewtimJWi7ga0YuWHegyc7/VzUGskAbW3OJqyMi/mka1T22
56DUR6ozVFHR246nRBCOYQC5EbqL5whp322xVTdvascQQKlp07YFVn8dmVVRTTit
F50RBD80097vg0MfBE0W7GYr9L35pV/vpfbiaGH4b7ee+q4TUuHl8MVEj2O3mNGi
/ZTc/Xaxy0xSKSj8X8UxhUtjL5yXU2IM2ELdfYLZeUNbBpQ/KEwVZotsdeAWAAdd
OhFKmF1E9HcZ232NHLXLFxmpTD9klicIU0XSVivYS4iUKnaBiW4lBjwZ7nKVQgkl
RJOTW5Pe7u3XaP1q44ayvcV4KdbekJYvzoIllewslAYpmOx+HbMp5uyoVi9EkDV9
PZPvqAwPI4NkqadXdx32sfbkRfWLOYa35vkcT4D9s6Gg3LOZBKYxsz27Tk5YBcLa
hX9MxbKL8aHL2pw+mk6heNiOJHqJ4xi76jJPqkM9pukILSTQh811ctGEoSTmSWaW
8XugkGj3WidtFWdGznLttcHtmdeW3h/yKTGjL/PkdEhexFLfANAewjjhICoki60w
eOwQghoiRAbhQtrFgK7b1xTCXrZ3AW4lO8NOLlZeh5bB+YocSZVhEZVzCM6WnRa/
ZiYGh0i/tuwBtjx4oFoHEBkAKzyCwvRn/1zgpjVQBzqFPWJ+kcANIUXzCSDksLTU
C3OjqoM/cqQmhdGqIeP6wH2n7d5J3MCEq7nHdGRS+yKwEL8Cc3r2PRoXN4wq9i7v
uWzOgGMfLDDU0kX94tTQZcgO6iwear9lj7WO7udvRZOxIMKzTfyNHOSzkWncHzG6
aRDU60ufGeMjm3zmDIwyK2t1coEq0mUBNu9Fn4Sfx0E1gFUXXtRN1Pbbb/IWY4oM
c3pxxQFT3x88jjJwmxje9erCfwJ1r7shZqdT9s2p19nCMnQUJf+uA31fgSnf1GxI
fnPeQNIRwLgQynp/9VHdsA3veMj2FOIOiEAyaVqcdPv4IqBbI/uxOdwsFolJi74W
FQGNxObUqcIz7bVwqckbbZgX6by77SmU2feb2FHtuCEIHrMGxetkQ3uR8uAx9l85
iZOGMJyiQfNkZQqupc3zp1tYLZQZm+svapiUV3vMkZ67W9SM9ivMnKmRZlI3cw/Y
UF6XW9jiYchuXjZMcc5IJoWD+VaF2GXedrQptWSbJbuh3BiYNi05y9mWmZ7KHJ8Z
od+EIZ6h/WnX+pcHPp9jAiEBaZnHlvKOHo3SXTSzw652de7jpJK8i3Hdaj1doGvb
svvtCwoSD7VoWzMCau4ptldhtQXpI0UVLWqIFKHr4q1c7XdTx2tjLN0hPrV/Q6zS
fGA+f/kYo7MTwTelyEO+8Wr3lk/qfntUk51OMblNsCsJ1COu2UA1Muyuaum9eZGd
A+c/QKNvYH5bHtBd1cn6mX2v7GLa6uWr8JBK3dPlWGFIRy1l1cGufwoShaWph5AO
dG4T5/ERW+y2GVPHjyQD/8a5zS3I5vIt1poVviJMXI8HuvEOk5u7SCAKqun78eqM
/dxvv/LC7kyfZADg1/g57FyaBGrQf010qGz7Pg3dfLJDNiCdliq6es35IGY41lp1
nYk6rDF4T9/XjHc3zduYs5QQsl7/+URexTcVTu9sJd9wqF0NSD5cW777ldpG7oV3
L06+uK+5Lc0Zh6c7g4zW56yvY4AyH+3Prc+hFZi/qirUr5hDaNW6XdEocV8IskUf
N0PLbuGiREF+LFDV2ZwrhaA+X+fj6IBl/pk3i67Elso5XSIc9A4U+yfFTolBNOYm
ECH/fxoAgQoKGilK1TKMbyc4TZMqwaUqevXj1FsuTfvSxtMMKnfclbvUI18gAiZr
RWK7bC6cWNDmGB8n2BsBQ+EPkc37HybTtj9vZZwjFpui5x9dVpcKludgjf9rl+Xg
W2RInE2XXPyNVmzQkIt6OjkHrfMRdupf+a3x6Zc9DuGeCnwT64m6LGQVNMk/nBox
ccOLQHvMr7BANfikIfvYZ/pn9fxNoRuoLdoO5KZWjGZlGAZbArAAagRTpLjPZtzT
lFt6mEEVUOvLncs6oFurqIuWFPui2yCwmRJuHz8aKq9utMmWCKSwwx6v4LG3iWbL
sqI6iqL22KnCgDEDrUzP46FtPo8rOpYueyI6Zn9ZgWwjm63GAo5in7QMIhw/lYa/
iFueP1IZl0BH8sS47Y1u/s+/t0gZ6vGjrn6+RPw8nmNyziCOBLNY0fR4U3eVapo1
0vHTiH54DPvTyJaGATmD8+FAusKDp++ay2bxGC3OmoaDBV7q/g6BhDbPLpt4OSbN
K/MjOZHT2/de3RPL3t/mTD8jeYZKoK0yHC3l7wdhC4KJ3Cw+ZpPEwke+jqxIAcQ8
p4MeRvF7opECrn51VdSrcEdG6Mr6Ar8oPxC+j9bEd8Dp+PkbCzPjnYIj8EaD3yGX
6vnP0+WzMQhdwXQw/bTUsAhvqGMPwuJ7+Vjo79cSAIwNkhjhlSeqYOHL5tJ+fMXW
RZqArG6swQapLOrRUb63/doTqmL348eQQyxXQ1fcG/A63Iig0RWa6v8E9dXxGl5P
8QsD+YXtd9WPiPLAQJCWHpz4On3sbvcuGIuTbZrujzjD8UHrqdmSpFB6pmDgRa8i
vnwODcgs7nIUWVSmCcrkoiadDVhKNdf2kzLbh2RQ9lOGD47WVPuJE+745wcyjpAw
umMUz0WhYFvFxKaZihQi0dCjrso56trMHLDPKCvAowD4y8bmOkUi1z0ikL8IoaDs
Md5xS0PdRzNhdN487LMNBbOY4fypAkOx/S0BypSFM+4Oab9pu1dCnsFEUqpDaEMs
2hqtuUMRgGH+R6rE5Fwyc4DEMido24bpxygxCG+Mxua22tIX/J8HcvWWq70kM4//
FBEp+b1nneo1dM+Y9CHggRxPgwwtF246nqs0MWUEdk6yZ8gnbKm8OCdSLlKggHxc
xJ9iNkYteD8VHo3a7xjJ0JiCgBjueTqE96EETO46QPTyZEruXRsXBTUmpscwnFqp
vrSomqIL7eAQjCul322ZYlo7f+oyI7EmUJkYCNcE7lFt4RKVBHuq/0gBdj2bidXl
DtH2T9J7rJp5oBpnwdVMCWdaFHOsxPlnjBphwW7GNcaLHIMCQ9Od+0aBtZxXJjeL
bLm+yUmvG5pcG1kawQpnDgMaFmdyC8CUyrzE2TfRzFdkvxLWLlL3euUX7dNI+ai6
zZTZw/L/3LJBGB2V5yF5ea0Lv2gwnmdqM6ZmjJnWG8YBlrG2VctoFrp5N7OiOXfi
brMP5wRqURZxmBBBhrMFz/uROM2Px30hpepofE+hTzG8iqVnCR886tfp1D09yTR8
vCCFEBE/7djFzhIJcQAWmk8MOMu3EoffQlJt91PEFOiStJ08h0b7mZpLdsd1f/Yx
0OI6jfTC29lVYMz5k1p0+QAr/cAyyqo4M+CRlWr3cyL0NsbPH+Qq5i4z53Q+8RKZ
vVyaexWe2fXdW8xwbMyPQcl3sPKUNzjeZStxZ7tKCISY3qeIZryimoijFadQ/vWm
faZRNPXb65N56uavSHTvXzQocwSj4xzFm62v9KWM55rjLx9K6BMIJaHRC4KRTAcx
BxuVmswwsVzqnoQtrrJ2f+boy6iT+uGaZ3H/w5OcGdgbXfq/zF7bqbhVREyZuFUg
2mzJ3sNqfhFWIY/85o15omAKTWmnPZRujJ1Go1Z6O+LyqMdq92sWeixQ3rMF1GC/
vBaA3Xzn6NxIHulDVKuaOswrcEPksxBRqlIuSCGmZJtuQ4nviNNxinAc4y6Y+Nqq
5yNCfleIQjsNUqz4yICY3eLDzNchn30P1twigzNeIxzWyj4Aepqnw4mHZJnvST62
/ughZucou9pMBb31bqZdt5iJ7xlxrHfDAhYzv18rn+01kW98Obc/UofFBhj2rMfK
uvsaoi0/eq7W2CYfbNGqAP8Bz57ppLGf5/B9oK+B8rvHvao1pQJ+9XTMCsd+QkEM
JWV4cQ4WVQg/8zz/qY/ASDcEQmnf9paC0efB9y1NjogJZ2mFh3Aa1O3VS8tq7RmR
gyw2YysX25bd/8BqGskndSltz1EDH/lMabGThxVe+A7EgaMlw4Tklk3Z56jHKOCJ
728uQ+scspl6GroHv/ykemPisdlUubBolknANXiscMyT43s8ib2Oo48RYbQHZShD
KpWUAdW8amy7r+qCHldfXBEBEbqIhKHqP7Py53LO4fzIce/AJw41+Y12Z3SyR91K
vezdhtAeybJVqq10dIuXJ4G5MpBBrFwmDc+rC8RiSRcv4s6pjGVqTO2qjUiyWps2
e3XshsVhh7tYJ0LNfXY27EhJeV0hmnq0vtOdqQPRkey2HsqHOebKP8NV+N738SxA
5MUrTVr6RqkzJOrzT9WBJWyvRuEe7xHb0+lT5rubMm84nug8V0Dk531iGSrr/gfL
NWssLlxDttgnXxx1QcTDmZ0VimVYpm9Sc/GyBwQhEC0eQJZ88typ2HWY5dUKU9Mt
fQpradiVxYy4y2w95rDYgXQgxOm8FZcjn808Ob3r9BDOgf/elfAkhKeXgF5QsMiu
E3IsnVHBUVFjhWqMpAwYqfGQ2ZZXYZYghWjHEr9WYy0pbf+Clmagk/M62b+oUlE6
8LPdTO//mZaogmayWv2JB47DE7f2rA04KBbEZbI9hphZnfQM/xIuKtvLmFE865Iw
WFJe+Ji2X1XG31Exebf7kLDL6alCmbVW8idOkrxxBmJlWiwwz8L4fqexdZXcHVoT
uoMaM9ZcDvKWEVAI8dOJBXA85ztqG7UCUzID7xnYyDwoyGgE1UpcDpz+O9Uk02OX
PldfrdnIGc6rqJPck5Yi4e3tBCPITmRevrlGBtWXnD24+mJjE4MP4Y1AryLQeu99
QZ4f9yCMHe+fn/D/QIy75zkgxJTSFoGmGK+WlvbVWywLrvptM9nMKWubI2Oas9ri
Hp/P0eeyg1Y+OnwDcN3ZaBcVeva+AyHy+DjxfzWY5IzCxFPG58pntPoc7sOVPlUP
1Vq1DJ0HElc0ZWJNRNzVlsBsN7n+foofizdwsmFH3H5Yt63Iu3FjiXrUNPGu7mZY
fPxILv0ymnVuD8QtDAhMPGeaGa2K4ApmUqxApxKGAAQ0XNdcH0xERbNnYhknQqxp
5f/NrjpqyJO+EDCItzQJ7uT3di1xzqj+h60Ypdy9GbtYYn9NeADX54VbhZ/VwWXb
xg7qAxr7hY51Bz2tBaCB3FNmEZojpzLqS8Jz902wQanVBvWjOjleqDbuw3OY2qfP
XwyE8ePWGGki5H8EzrFIUBS2eSp4p/PFiBNbBPe6zU1OwU/IsHmysrtfEx7wQhYy
jAaC4mGMHiL00SOLKn+u8QnWZWl/T48wectpoEB5gNVT6tMR8fyqcc313nw2pzmm
CHAIrd6GUEGa4hpflVO/BgOgndy89riSrwVG/fjtMP5VWLc2vhciBxPCYyKi2vY0
AZ12MPsLYWCjwOlsY8J5eIN8C1++Y7WeQh55vON5emIh234xiRK6GVsnIeq4kDHz
h3QqR3SiZb1aXo2l4D+Zyl7VbrZE3vNFJPk0Q5HtXj5vVxQw6R41p1wqgn7PVxUx
CsxFpOdzGxJX9MStYnHIWFdLAyyt2ItivszCLKLiczA+hNqGcHyE9YLWQqIcTPH9
Jwm7JsRREIVL/OdOZTbFclJ1FZUDwoQfB2AJqIF31HIzN7Edt6hBVLVFqb+X1WrC
Bc5p/d/TOdc2rsdoV96g31NS3b5v505hKPwqIGMyEAjlya/e9Y5PIJWEVvPpIhni
dP6J2xzXoBnA9cz0zK/HlSshHV7Fj478VlxJT39v+ao4kcEFTPT5gXSXrdfUjrab
iCBgTv8P6syAqA0QS69hRqA0JnVuph6fNiaHoE7oePVV/p2Qq0pE6IzsOc53Jrfl
RQYqpy40uHyDJHAJQ4TAkAMVb3kZoRtk2e00lXkrmrd1ILBNbE26P8eOQkApi6YR
vxuP3gLu1u5sMa+3IgV9ZVQpzs1MBoK8TCEsF/WG5AEUNcytFrKUS26ErIq6wHto
MOSOlsqKJvzIpiBJ94GcOFFDEecIZb/IbLqMShZQP9FR5zbpytH+QyKpbYc84WJE
HED5BrVyvU1F3hsOvyqgJcMymK+YtSjxHe9rBT9mK0lCRCcUWXWlHpBhNr33cSoo
ySLE0AOYW8FuububrnCcx4rxMmhvCmQtxCaXkBJlefmPXpEAF/Xo4KnO2sU6wHcE
bqESEk3XL9Mb/1EVaKaFtOXKQXGkL7TLSKgGKxRc9niUTrLJd5jRA5ISuq0YhiS7
qft38g6q/mtLjCnNiKu7ic0ZH8MYmadzOmx8XB27gCTw4cbNTPS9209EHpfoCEHH
AXEfqeH7PvhBq5xAT1Qv6vqew6Y6LvbEBJ2k6weYGpywb+9DkKpn0rNZLsEeF8M3
PI4sC/23qsHtdaK+VaNV1yoCp0dbzCubaapB41SqZwIBzkwItUD2jtrFw4L6c+N5
DZuhqJCJpDmRV704+mSjok4ZH/UJDy1Cz0R+3MClU8njiYB+FfXOGKyrWYafWTRQ
FHt98S9BqmkFayO8ugsIye5AvRma1vy1GmiNYItanRsqcUA5EKbNmvGF3+2M5hQo
`protect END_PROTECTED
