`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/hirfOV6kBVQuR1soxSh60TVUNYgVXCgt35HBUQFGNnEJuZrEPDxA3MEGTeL674X
ykv0Zs6/npOiofRwUg2aopFuoojj7tpUd5VnS67YDNJ6euYd++tvX9yDBcoQhTB4
LQDRk0xsZR+xjVjiUPoRKPnUzelCqXxvdzFHPNPt0kbeoKMteKNv0m7IOj9XiuZp
oWhancTp1o7HzbUMA/hnGDQEI/106Jh7Rxm/QClm1EYavlFryeBDDugRjOE+WZV0
3q65rwMU59bt8pZWWKTPTKsBS33XhSbxZohVf5msirxvMAofbaWvfFpbxGcOr770
UUIGrWTCLIWVtnPODqK+8r5GZ1SrTnTn2nhla9WBZzLvnTo0C2wyVsXumseVBXoP
SVdJZXwHHvRX6fh08eh8cWC+ZUm5UtQqpU7vfLdatK3gTy9TsqEUtvxX1mAYcfDI
lEnM3/5+9lwkAYkTOAeGYpBywaj2i5O4QEBAa5FxrqfuOQxxlN/awpktw82hKmWU
ZjiM+3u4PHqwVPnbDyk+ANkmbINcfg8UAgL9WwynOOYbNuQcqTiPmPLsxzo1XF5x
B7zKN82hXSe/hSpvHI690AXN4UvdiiTxGjkp9CEHIJ0qw8VBVEWMS34HzqAo+Kl1
inq84lNDdMpEipvNhX9Nf7YVdVVgS4Nj9WECdQZ6m0abYF8LU6qcU1HrIOxUOEFC
tmX8BsnWW0TZ0hR5G9DBcBbWOHMotk9AjtBWilK2kBAp6aG8DFieAs/fEZ3QuD/P
sD8CeOg6Kdw9Ng7U1VvKRxO4xkcEvnQao1f5Mig/qgf4YTtBzeubW4puFe3bQ/yf
4MQJKPNZhDU5GE6iApQcGY5mo2fzY89BI3jNaJ/IcR+V2yYL7m7NCycA+Onxxis7
4gZK2Vguy2FxJOnIp36NOeAIVb6Xi7XT+MPfPVyvDiELq8ZsSANc38mjM79n6mPT
pBiEIoalXOp+g2xDaN2SvyUZwyq8+XxHu/V77lYlLCij0qQQoH9vRNSSibgtpbIK
QaO+nGFTNriC+e4abf/68qOGcUhEj5/7k1fPb8NVzIBGDYxZ85IxZrjsJspQnPHf
PcC/Hpi4P0z5KbOPK8kWgNJGjHoKUR7Wy6vJZB73hXEVi421IoHMlyr/jc4zDtF+
IlzXDG2pQLQ2Hc6LJ0PsUCQplGSayzU0nyibyDCtq5BrhJV0493UKoENlKHTSWFx
LjmfTAWgwUPczivL3jj0aDaKvB6gGBqOYm9v3kDmHYJ62oIiXP1Rn2L0uUCqo4ho
3DBsFVKHunbHrn+9P8J+iXYeWgsVvOSN/BBBWBtSjNDoyfPhD1fP6VkB+d9VeUg2
MAjbBpa3KgkVAFvMNtSa05oNbDVuSpfthQenqRd1F3TxPjtcbcXoHxZdRSLdc9z+
5E145sQwiuX4+eQapsUxJXdGfMiRi8ZIk7AA/WKeadh867WXe7cChUNMR/Hd2cnS
SzfG73++sZNo78rvFUzLOyCwdQdhhC0dkNiy9gWHLDlQS10wG8S8Z8Hxloz1wMDI
qJnfv38jpai4SBEHxqv3StxfAH1waqcobMBsvi5fAHv/HPag6q9JQdAotFnec65o
KqUBpZJHQRib6PqfkzV1mjJIYdUiwoUNoHaSyxIBGssxQYlZcLESdiR/BbO9+Meg
dX1qcXNT1DpzvSlx6p7ffTk8yw87sREOLp3L5jgxwMnsIKGYQPpRy3s/5DYdZLxx
sJiId6VNlmJoAgg+21Di1lrElzebehWMVOXJkDjQFg0nzMQiSr0NhnHYuHM0K0B9
cZWoiMikmw2WHXftpm6fQhiR9agYsrPE97hxN2Xr2vuYN16CSAaslkNJGmDT2oe9
F/U7mDWkLIDzfKYUyqYwBPpPo/m/r96+ydneZAhJqvWCZVLP/ehzg8fjKWypimGf
VaR2pmNDi5/8TuPVnxFaYvA+tjByq1RSUn3JpCANkfNPRAWgLezj8PH+pb66t+Kr
+Krwj/Ms1lxOhukPDJ0gt8LY1P2X9NglplvrMncYK+slBH2AsfO/ywrGWbuZr1EG
7w5c8lNTi79KIIHhvvUQJr8k5zm34kPOZ/v0KC8MChyzKoY6p00i/ihFIxd7foRR
1kBmGrdT38ZZlalKBClGF0JMDcJY58kH5uVt3xirV54=
`protect END_PROTECTED
