`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yMR1lyi7iOMUqtmmxNjXn+vUQYgWteVyXdepKwi7bh6Eh4DUZwt8vfKeevtYDJd3
dT3JjKp4Q5cEikMa767nsMk579A+fhsth6wfSET1wmL4QiDU4lUn8FPoQCqgSB+l
9YK1DYaq1wV0NeXel4EueIogVPsratW0005sHj7gy457OyrbHZiiWNGMqnGOtz0t
wADhEJ0dDG8c2/thrtV9YKH69BOfrf5tDbGYCpCFoMlBb7GQ3ReXyvJlhLqT+sLJ
nAbVNZ+nEevhp0UYLWj/JXlU5Kp5M9+QX8UD2AWr2Q34nMFmx6evMULpOw5Li5xu
0Qy34ykoZgiMtvR30acPBAJlqW5ufdFUslossVmfBeP6dIuHEU/XNE7J9jjpauwk
D9u93fTDfrdJAM38g416ASQQyRIWYq0+XAy6avNjsPBuIlV9YEbgZNIa8AfWtpzS
slL4Fd7z23aVFytcX++LJkc18OsnOW29TbNHoFSvjSn1kPOQbE/KrIJ6C+iua1ep
lNr5NjazwiLsf6fmuFCIi1CLBXmiJe8QTHzqIfFiyd+TRWonm4o5mYHJIHlY6OPh
lYY0Ydrw2eZwvOUmALh9rOk2rHZz/UvLmXKC6BRDiYg=
`protect END_PROTECTED
