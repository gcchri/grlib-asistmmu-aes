`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ciqnEnXkp3DbJr1vekwgYXc88vZZnTgTFbQkNyxUi2ikYGkLET12B79rEp2cXQWW
4uknoBeMZj2BtPfKguLAhmEjxWI0fK9jlbtE0bajxCAk2TM3kFtdU6EN3ZRwsMrp
t1zKpihGRxAzKDT3ztX7G+5KJO6wU7WwqLEsENxl4LktDACjxe90D/vwrZ+DGFrl
rALF1bV+rX5jBGErwv6oaD2D6U0KLxthsn9rIwVdyL4BQKp5c+6zr9LK+JwuDUYe
a7a54bxmPwmAOEsQ8kHywcK4Yg9rCm7lgXPt9LHXEQiMXUYrZKxon43MVbxr5mvQ
U8uYYN/b71ch9KOOn5EJ/szcYZtRES8daBzbxd0BfMkLFtiBP7G9AbudExcD2pJP
6in6JEI4jJ7Teyl9UKDR3rs9/KWhAS8WHfk2+6SyLBlF/ATCKgEKD4eex4hL4+Q1
a4Mz9bH2RinPgWB5TJCl35IraVBU4myeMIYDqreidDuzpqN5egv5E7EWpZGSiMe8
qRCnwFeeZiw0s4N/lgk007hLE7ECn+ajs/OBhuwOtfT9MKgz2+L7dactT9fsNoEz
SaxIR4HLWXpdBggIWU5cYeqckVoSWB6EYCT+G92stKrs9QgHgiYTf/noIV07ujZY
+XWnQ6teMURlNQHwPP9mgFU/sN7v0QPu8GrxmUl9I4/ergiiJ+8CHM+Fgv/x8/R4
ypvIHnlJZuNMbE5qeuho3HZ0jIHYmhIjGkjUldScNPVFyVjcsLZPCQaVXH4Mctze
WgEgqLPHDlCZvkblGgaWKAJGt3UJA7NpXdKFmksNowKoVSlibCraHUi1B/sdiQBM
DQSF92b9txboYijvFxu5iU4khXTU7x6GaUpWZRSeE6F/a+noS2RpLYkntKwlcpu3
p2MayBehnzGncljrNtdWyVGIC2UIMrni1keE5gF1i3ukxszIb0wnFKR5pCR2G+WX
+8X0pmuIu1oU8GhcIczvUGr8Uo+VGVqPbT/bwKVvID8cscACPVGie5bgoC+x0cqB
WUG228bcecuvje/BMlaNNwiCmEF+4mThHkECnIKLtmRP1adEz5moWdwO/v1U3FVa
NEwZe5NQ5J9ugtrnx2QtwMMnhgHyodPiLx3wY++9l+2PKcebnRMKT35Nqrj7IGaA
4LABxfkR6dcvkeJAxCEf2bjRKIiaYpEYAy6gUTataI3738ygMaHQitjy/cK8uJiQ
ozU8bLCQ+/4FTsehN8Cj/4WpKKI1M55CoA11mUHipo6eGB9HvTGUv9XiKM8Sx9U1
/7zuJUwekXmihQsja/Ho7UWlD6FdiYXcN5pkEcdWjnQNsdOGfPMk0cLTRejNXPi4
N2vDInKiOs9BYe2gF2MjLdkHlsHyJ9pM2g2a1Qyx/SNRnZCdT+dclYWmW8s+kG4T
deMDey0VZ7PxuHpPQLyCtw==
`protect END_PROTECTED
