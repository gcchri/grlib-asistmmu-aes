`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5HSSizDBuqPZdsavsF2/hSrI/5rzRVUeYyHsF+cjmsutLwDHQWpw5eOSt7rFVxfp
GdrPX2i7/NjBjPl4CEC5pBdLj80c4h7RKV0FWQWEzY4cSiHCAyIR/S8bWan8E7wJ
PFvF2KEbbYfxPgV+lpI9KAhx88iVCRZv/83iGT/MTvBSo54soHeBzFDsaOu4KJQ1
i2UlVm4McWAGLKwCWcJtk9HGQDpgUHO7CiQUc67bOizmRjM46LfwKPT5KziseKa/
nUQx3b4SMC4IbShby3CPlcoNliMPjPRJnVINgxfICiF1a5y7Fxfp7w59RI3nf8X7
txBXufWM9g28gGSdPxbqSYd4BQkeNZzsuSdGvd4uQ3fQfS49/cCEBufcaF55JyuI
y8SqtvXwtoJv56BmUqGUcMFn3SNXFNkR96OwUjEULkDxWNAQI9jMiZIk9MR2J4B2
rAM5LKDDwq0sdO2snS05lg30e4r47phedjlFJsaOwjA=
`protect END_PROTECTED
