`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iU+ift4hyuyCUZtDoNe4AfFAk/JF078pWZ7uBegURnsdv8pmL7Ryv/QcyCd/pdPG
TpRRmS4ZmAR6Dll0DtCXroLl/yOirWjh5PyX2RHYOvOsiq/5i6fPrXp8kJxDOmCt
URnpq5LsxAuSyGZPfrCAx2MkLwlqR4GlHfXtohDEQVDzK9VWND/VZpPewGoHDIOL
0D/ebzIh8421v5LqVERTKR6Ij3ESz+gtw2H9jplS6ntch6XqhGNF9KBaa1VBR5sJ
lt1DSHvDf0njRT31nsLXyrBhbAuocomrGK52vZwH9nT4U+G4kyoDK5JUCz4bDv19
5A+f1Xw48unLQ6UBJ9QJCBMc1/2bmBYUuP/1on+HO6c9NR7HM1r/WzWd3vDosdt9
Rby1U6jIikjucfqwOA3vGrGk2HjDyhOKgsZAe/APY1bk5Yw2iDQt7rNSTRxMR5ki
AAmA+l60zlO+vfx4H9dUBBohQkFHgr8LQ0n2wUDMirXFzvu2tiv+ifGD+gHbikt1
08i8Zc6H+FYP0gD3b9k/bwsUVJo0oCbd6gwsy9QIY/LESRroy6Cxniq+HqrJevSl
QkLkrFrl5qPQ0EBDKIbCCVibVvCjBvX2dCY0eVqbnoy0wAI30RXo7XiTeLDUZkVi
nWeKBT5jBzs0l1X7mpfKbjdXnxAtyCrPi5fnO4Y0BKxJ+lfiHDUpXq7DpyIW6vZL
nsQoHQnV6s9B3EYG+mjpGfV9m7ZtuROLMiELXRPZPxrRN4QuSmcz6YrMeac5knhA
Rkl+Y6JT0QV5dIKdT6YchhWrQeaB5ikNaeHlqOtVCQILHv2RYW2qaihuQOU9DZRL
zeM0Agp7uPh7Mg0mHN5z7fzdzqhBYPGuMZNyzwqQKwtl5314G7i5afZCcw/L2ghG
2U+4QtioXrGsJ0rnw+cztBwkyX8hrsX0l4sMZ6Cl8JdcWGYT1hpC4WsPitefmMxf
f+M9s5blFQ+rX7U/JIH/WA8ADuKHTPOYPfPP+DlCgO/q5yHMnmkXuyKluFRW3ETZ
Me3V9P3xzaE7iep8PxdzXQ==
`protect END_PROTECTED
