`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+mk8mgDMKGcCF2NsxO1lQEBsmsRJ4ylA7OHoDuJspUZCe0PgXRR852uyzzWBs10
BmggSQ4pabcvvVMKxbkH68srtjN9a0zOOUhAqIBznwP9/jkOhBLptQ1L3zLgVAIA
TnfA4wEnSz4s/RrlCcBYVKjZLBAwyWGWL+GVEzdAMQnoj8EsLPDY4wpKVmN9XcYD
WqgvEgxmwX9WY3Y+Qntl6QrFHobG6Ty3Cs8vWWWgnmKx5BQCyH+K/13CN2KQZeB1
FxEl86sEn9Pj6Hw3nQb9xO3B1pX0hIbkpp1L7wjpO+DI30iry4CfUGBDRtp3UhTb
MuMFTQvWxVKZlJp2m3N4QdL1lXMkjey/qWRvL81puQ5OtV/9dbobPx3gazox+8hs
Ua5CF0lY8vpwmbuolI/C6aQg3I0194gSv0jU5K8h7ojuiOMxdoUIEipLrWLgYzjV
eVebwx5e4W2w9apZaENnKHy608wsA92MIIOz2omLakVX9bdQoU7gXwM3wjv20kys
qIppgqgVad8cB+pkCZik80OInQ2m6qmI9fcggDb7RvXMKILLm2SfDehAohkcnEbR
MKFDui5ET5ORhER8ktDWMBeP9iUx1JCiiNq9E0ETEbZTWQPYSJGV+tJa9/WPibMl
K7G43+eCJa33z7GnhYflrdO+QzlhD+lO0QMoHb4m3TeK8ocRaomNlsZhIeNgguHB
qDzm4+WLDLsdCLq1yyfo7Mw2N8aYlhAK61kYRkQx9Gj3FTfNaNLIVXp/yJOebnzJ
cRyDnKbIGRiUfG9AQLUU1OVSNkWcaCpfQTez368jLop1sgj++sDMX76P06Bvgshl
ecHPU3g1CYe4CPgbJuYb6pSoIjzTP8e3suoE57rXdU0=
`protect END_PROTECTED
