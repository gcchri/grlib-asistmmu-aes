`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mF0FDK65IfyGSwDzjn9J3P7qz+zCXO/sYqkchNUTb7SFl6diCNtF5MWD2NWwSm9W
+myKg65r6fzKgGhTN46gd9NsL/Lx6Qfre6Zj7q+HJyd9vsOMtazsLQarLByvaNuq
h1ym8FwwUBF+ywAwni9V7PU5rVKySy98Lr91Mh0AELjStcGg3Hi57xTz7OCFAOzL
xkF6xlj7M/PeYQhWJT5JXaLXj8UyE7my0RIqnNPeTe0Nc1DYEuu9KQQ2kLzJ3efv
8bcbK/kPi+ZpwPX0gPZxMKGwlTKcJfvbAGhElBDV2pMLweUznpGnLRqRLhKVIMJl
y77AUZYgLJbBc8v9XEsvvO+lGoZqasa9t8uMIApwme3QS0yMBpsMpLC0Kar0sX5e
d9wsV2ZzgYLwYyTTc56pInpEQigznukZNFjQf55JbX5jML8xn3VYVl3LU0127vhA
eAoW7jYSh0UqijmNvQiU9hWadwzYXZzaC0oRXq6fVBil/mbf9QyP9DO8TyRWsAhu
mec20L+KBpBLQdUEuV1EH+9J6idc+ePtYU3ZWCBPtGZ9MblY3qX/GxyXYeKV4UR0
Q5rf4/wBMwEiHLOL0coDgMv2in9dB5y6xD9mzOHHf6i1aD9uxkroy7IiRyK/acg0
1ZFX9lA2ol+Q+otk7Jc1uopHz/Chr4ohhFFCtyjJi5Q=
`protect END_PROTECTED
