`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
myxyk59HJ/Yn1NmHDqisvHJ3M8ymXQS6eLAIGwIR8I7kwHcTDvWWMERAmA2PTXuV
0HRepnL24RYjZ+XwfCo3TijceFas2tzkWJ1lqYWKdT32oTngPlneDU28/ikk4Gdf
VqglwVi+Bu+W6MINZSHHFJPZAY84YFaW24twy8GLf2tY+paQHxpr3amPoKq+fkY7
jvEOT9n5e8IVy8zLp+5TPh4fKkTOt+EaI37rsmvPsO8BGYM6DF4Q8EuQ1Nr47u3F
II40Gz559h1913KUr9M4HpbJRh+orri8KV9oAntFLP9gKEbLSPH5ktRvb1XqXkKQ
+YXIS/LcF4UoGvxmEt7Yc+vpgVsmYaU0D6W5sdH8LcX2Ka8aM3Fiv0qxOAsm17z3
WVB5ECLMgh3OBJpSQ3n6d4csBSIBjWRwvxp8soEefFbOAn49Q4ELB2a/Kt3ch5Hd
K1eR9bwB3XQBStvgEllxdKK/15E3QGiysA39++zaP0iQ9yVdFgYZJm+PkbZX+k7A
G8NwFP3oR14Xl8oGGdmXC/KVJPenl6jCnONI99ppgNAc4b81j+CNTfRiyk3qZxa9
br15DlAcH5kDe7LEiBholv0c2sMHdP7mHeZs/eGXYpU5+z7iYmcHJvd7KiKdLs1A
c3/g3wDMYtma7v5vR3tM+FBk41botlRXx5e341hQbpfrypwpQ+l0EHjHID2GXzAR
m8ek2vSsneSkSWDrjcgOFA==
`protect END_PROTECTED
