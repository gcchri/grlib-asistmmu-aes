`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOgVy4OnlZltN3sHlBksqjV4F2xVF6NUIpCqenuqIwJ8pjSm3meG53avwgiWPa7U
QvQLk6cxLMEB4qDQCAYiEJW/rixxaG7d1Ay2pjx6utbyQfj0KgihcE6K37j5Qfu8
9Km7igb7TB3zV2INWc+XIeKzKnCH1S5CWhWCTqn3zRfnTVt3VdzaFNIdgoolLvQ3
50dn2oQ/QJpvUj+8toFMuxdGPCljuDrdS3JZUmgNuYDx/AMLl+csGRRZp69kogCY
s7HB8Us1bYiEY9PgThLZ20tSQwINi/nK87FG2pWiyewLvCwsl/NJ81YZjcUgv67s
aIb9iwAm6LwHUuBCRSwRFkcZM/91j1OATKm7+3M3+cRhsbEE9xvMGGmqdwmTygxQ
Dux/ouBOzd25UAbdAumqFIU/EHmUXLSbriroYRGWqpePKO4F/FemreDXT+fD1KW1
Wj0P6ZafeBiCaAFEgL5C27rveT9TT7zdhQAdi8kjR9WIBxSXwixvzNm2/1KBIOh4
h9UqQu34FBne40PO9Q624E/H8CglM9XvingNuduGICNIlTHKqFr3GQWj3mOxtCQu
r68XdZCCftOEkB5Np2sxM39si9cyY2XbL2GOz4aOMWlkLb5+qY9uySchyi2LzZXf
Vh9LFfCRLplSl4CJrCHox0v+qc8IjyR8HCU7lJ6rC4zXBIHwdU7qvsYUOvn4JZwY
q7ALUJ4y8jKW4LvN584eWiT4CIeuz/Rnma0lxkcKGbA=
`protect END_PROTECTED
