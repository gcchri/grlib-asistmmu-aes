`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kSX7/i3EwC8fviwcV4AE9QO9tDiBCq1CTn6OsCN+qVPwrfoWz/SsheFckb7SZsiG
9T0uWtJlaOhL2JUbSdria+07K7NgNTJ+7A+igLVF+UtskbmsVt5LaIbFD5v7mxRK
uE3DcChqhFv0fW1X5EnZz7cqiifwRCKMKmOWUQzxSlJrCqPg7eyp/UBMtQZ1/UMM
K7NBvWKuu+g4PeUtrpke+h5w6a1F4rZlam/n/H3wI5zBnSt5ybnEHcHEfVG3joSD
rb9XONeRFj51epFt96o7H9ACD+0HeAyViLBOIHhhRvPOxFuVXpAy1rEQSWNIjDn6
suYIFnPbSEd1I31tTcK+PtIN7j02AANnf27o0xFXWzUqGHHzyhxeIvoRWr4JC/o0
XBXDuvmeGmVmN0FsywAarntr3nYaZ+2bzT2NmKqGP/KJH2j8A8SZekZhDoJgpwTK
0DYbzhJcSrLR8hYhJM/QysYGWi+geuXonIqrmBGKVopAHShYQza5lcGzg9nN+A0g
MdoFJbcSh5DuJog2OCSRQLXepmgjUrTYGlWhQyBv6xFylrhtyTBm55RdffxxAAI0
dAubNL1GNmnMSOdT9tTM++Io213ttMl21uS83jINw1blOSXtERITxpHBfhiG99d8
1zECTRNn6hB78MLJADjSeriRh7YyeBSYfmli6yeWXkChfzKZ1g+EYL1PsPoZy06t
tcXkaQc+newPwaxNWriVVq0oADCnLC/6+T1+cKdY7UVSsOgFpMk9tj16eOSgnAQx
umqYHYcHM40hKtulm+4cmF+scZYfxp1xUeobZmt//H8FugiwAXf7c2CFrMuY9MY3
32OdI68f+JjaBPh/sa/sbNT+W1MVDIk93ghbjsRsgM6JlDd7XHzkdt0EnKEULPcT
a39gCpyI9exGE5NsYJc2JLkWAU4l8OtW/RfKlQ/ySOaPsvrU9tGBCstHazL5h+JS
hroSqRN86npvjmqQQm4e8oCs1k0UbpW5elbt59fXa34=
`protect END_PROTECTED
