`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p7nnKuPspUZyHNWZZ6RD9QYvn1y1lxJNXCCbAMjv+bkQdcxqdIKIHSsq/f3dLQxm
8kCht3OTqa1f0Q2JtumDEgXZmBG0vCrNZAtkCHSLVGzu+DBJ/x5dArS5QIySoGQQ
tYe7m0d1c4bo+O/9MEy0E0pfMLTksdSFCLKXe9KHqt2Hs0lPfuDpNAK4BwqarFJq
S4U+YQxf5PIf77Rae+y5Y66TTc4NzqxRjgKXaTV1xz0SstNBl+wWwJBSLMsLN/Rq
uk0nRi1BYIxImYeKKkx788yGhDu8zC+ZdJ59iz/MrlQBJTRPDlzkNrfoIFGShlGO
ISFELuhUxkCT71teK+yF/AdvuZFilqx51Hb0SkPULooAmU0nrtPFlMw+QOD6CVYx
GDhUoQARcAgkFBlVarUovXhNjufpzFNYBPco5sB3Nkdn96nRDdF+aT55sOVB1Eb9
IKstBVyTogR1q1a0i07XGHOcdHu3fb/+7O7mq7xWhdNyOg+nV4KoFA6XTNSlK9pb
vPzw90zUjtzysHKKihADvQnUeUnONP9YgOL0TZZLb2oJ+swnrCOkop/ZePLxZ2BS
uNG+7l7PrqaJcXN9mvU+/IQij/IKRhBbpGcgr7jMddxcMwVhzvi2bkWMklAf4LAe
kaRe7D/BJQ/ZqZEMsKdW4NYAPFNTlp7+JBrtdaQ5Z8o=
`protect END_PROTECTED
