`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmRnESu4JOWYNrtv9KqRHUfYUmucrGpP+FW+j/S04n6lEcW7ZslZn557oePIrE2j
7U74HZvOh4Frt/1xDjcGDt8EJLaOA0piuP600mzvPtimcAwlm6UcIPmxmgRDhPGO
OXqCuLzKSE74elhrj1P1kF24D50z18AhLQd9/Bp+McPHbaFf7NKPL+KH+rO/sZtk
8ycBbgoypCZbaf9/rgFTmgYpg9BDMP6CaZR9/PxiN0t1uZ4JuIypqt0O0ZWoFc8S
y625ju5cHI/VQAAjVvRndthkuB/p+Cge5j/ZLyXbMY21Gdr+UA05H6UK8NhK8Rr5
Iv1fp4tw4W+SxAeIKLruOavfqhStbDUJERRIFhvt4539pk1dG7E5vwzYzFGJpksN
`protect END_PROTECTED
