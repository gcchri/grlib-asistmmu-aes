`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vt9FIfgy+XiC523QtqnrHJTVNpFZAQtl9Bt6vNHyhZYQdNwT5kXf7vTFdhBaqDLc
IRCpSVeIZbs0pBYWzu6F0XqHoL5RzS79rN/mJUXt9kszlbEfCIXRD3jzpk9b9QSa
bbnbeEVCD+4ALNU9xmP8NSdHhsO/yUkVkTD35Pe/wIWYjcliMRwFwM+z8Aipbrl3
ZXihL6FHKHnCbhynEuCLq2qZ9Q7INIJLvyXFVmm/ZtS0Z/lGNVWAJJg4bZdJU4bE
ZK6UPU3ZRj6iyPsLiqvvLtqb8SWOAIbIxeC0Akln/UZo8jNKNfatnGtri5AwNzUH
vVNvDLVlxQPPhPVE/VyRa0p4xEVLigD5XcE2DJUEuyxGSKl/j3L7HsAXKXdfxEgp
6lsy6rlySVrj1Jgml1OkZexUM7nM+SUrO5XKzeRtdhJ1H5LAG9x2Lbcvm0KwUnRV
TGy/pEzkwkThzBRAcPZ2AHfA7zWc4c0cHBhtGMBokamjMxuFcEfX3SblfAs31yX3
Ak1RrRDnDwR9qr7LRz1i1fLJqo/uNVX1B0bPu2vto0A77EUzzrcSgXls30FNOfIX
5hVnRyHw4LY1fDwnihj5zUEH2TC1nxvDAO9nA5H8T7z6J6IZvT2PJQOWuCRFflja
duksyw0sDuUsSYtS7goNPh2qbCvT86Ln7K4iUHc+n6d18JCW4kJxmZgcR6XuY/ki
Rom5tXDTII0xdSyzmoM4LwSozRKmYDPL3eIhgfd2FWks7R/Ng2psVzeUg7wuRw5Y
Bykuyk5USh73eWac1pkIp52TYDA2KXID61W8u0PKux7Jdk6QwvwZ7b2X+izl7cph
5nwfdtJdS09IVeUzT1HKP+30AHUFwKVB9x4qUZso2E0FaDOyo/zllgwGSEw/Npfx
SGrRcLdCO6ZFs1tY9mLDx0YGnFdycbKG2j9X2Hx6Ww032XGZuLdYdNuV5O+O1EyZ
4V4fOeGI+4ULM0WSOTUwn0GfoWpctWBz8g/ofLhokEaR/CwSotB0JpZbpX+EV7OO
KKbfc4d8JiTKHQiuNuy70YXuDv+esFA3Nj7ugi0pFTH3ygfQ3oISOJBAX0lGk7GC
TV47RwItzIUuYbQ79PMsTadxkOZDB6Gkr+adGouMNx5lsvzaqBDBZNbEdk5nz89o
0sOFxkxcXSOZSbZkI7Clj+1dD9zCVEsVJwWcBBCkE3c4OEhjdMmJV7sDGbTclykL
Vl9SbDgiXux+TuzYt+1M8h6CWcFISDdgKdDWb/TMOegnk1RG1msKHAUkvTm7v+eD
YrolVZvnIe87MEOk28RfIM6Glvu8J0m5lZeVMISQvDBH6jq429bKINvt+8HNEbe4
LTGmtTRKH4kFGh5/9ynx24fh8qBfr3X/lHTMBN1aL75tDVkBgqZryrsDO7hXa36O
Snb6z1znUMHImOG/E2JUF4PFmDLvbnyCJegyu5JY4G43O9/BijCoW6ts+V3T1bv1
DQbwT25RhPhh9JiynSm+E1OyrXbG4Nl5Q+rfRsw9Gja8MOSgmsWE7AEdgsUVDPvJ
E1VEjblaAovgq4M/m/xbJD3DWn1Ydygl/q2rdTAqI05/K3kXlmbUaPupzehExE2b
bmyFS+blnCcIaev2Pl5IZLhvnIcZ6MEv4pXXxuZEotwscW6OLnUKdba4XIOrrIN6
nY17x4RLi8tg38mPSnLo066w6rhCT5NnW+N3na/29VnYym6GS7rQHaD4Wvn0ufzz
qTgfeTNdb4eRJTxO9YLQ505l6hXK3u1Bo+Whw6jObSWor534Bn5L9YSv2r28FzAb
hHe5GxNkh/jF78pucmT+eSsjH+epnp7H4tWv9yr91EXxrM2fJPuaLoNz/BJ5euec
cvafkV1/kDPJEpOqa6/aFPIucX6Shr4cg+ydmMK405HGbnxTrYeC2ckVDrVC1P80
RVj3yepKFWKkE5g8LbO8URsvmQN7XgQK3b33FXXruE+K9kEZWZbALDmsauQqXC5B
hGJD/C+yQSBjWpcM87gk6wAZyg5yKIi/esJrPM/7iJmM/eTD3FWRzQAD9lUrKmKq
9egWplWVEIyjRbI6sDmUWlgWqxy2mzlnS7svpXqnJFhGRS2b/2OaFgwtYCQQ6HlW
WZmxtPxP7nL4D8jN5kTIKxQKbN0sZbRfzfjNhlKM9as9YrfsNvrAfXWpLmUZ8eov
10wFV2IoQsdxOJukxEhGS6v6raGyaKGtaW6u18VA/yHPHMJJgIW/Drh5EhNMv7hc
wkAs6iYSW3/TdA2Gm4ff+SHGQ58zxpJPO+diOogryczB7PD7uqfLQn1WMPt3qc5+
mPQXJNT4SlOYrjyAtbwzut1s5ugDut9x473BRX8PbC2gD48aLq11thJETe6jj3Jt
U9IUYDxKFzu22YCsA96eTIEpalhxyG2qX3Es7VmlE4RRKjNgjBWvho/u26cyCrrl
/nY17wYi3DBHLB1YFet/CQ+vVvRBrRlyTCOL0v9+HaDkLRn9FoPr7EBHAamigDg4
wMrMXkUtndQgsSsVo0KYLw==
`protect END_PROTECTED
