`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2QYPCxcAkmueHlNUInciTAsH7/GZQZXInBo08EHMaDsw8onlhoDWYlFUphHQoJMG
TtlorRCb6dqvVw1mgYd3ShHL6AvmRNDphDhHw8Fjhy63spX79bVppFUKdzoPC7Rp
qEw/y6zNchB46h/orQIy2Q7yezNBeHyahYchJ3zq8WtCSwwbkMBhOPsR9x6pn1EO
GwvQuowcx0bWrQgrc1PPiXhBguzRrPmuZHYkWp+gaVcacPT+L06yvLxKAfd9Cg/d
8m9WMWF66rNU9TB4vy8esGh7A5R21EKeSsYMDk2Jb1CdKJY/B879Di6PcohXGy2C
NkyIbajVd5/36wrmM+iMxcAdag5Hj+Mry2yWvjC9TumCXpkuJO6EZ5wfBvN/47e2
i3JyWH++rVVZtuET2Rw9tcg48fcn13XjAgCkXTVIEl+6SIl7tnYoyqe9oocKHCeL
/26AYp1o0LTmKUlMQch8xmzJzFETGhxti6TqrY70mMYMClCJJkWTJ9u+vj4AzhBJ
XHxYKElPeQNxEhllMXGXmmySxh3cE4LBPB/SgLLkrKyhxbfXBsrelmH3poWjpNkm
24/O60gBM3Xxq6bEYlm5SEcXqcIribBzFgciWyxWlWKqiE28M7hL9dd6Oe247mww
72bFnRmIQprFHzgtiDh03CHF6hFde2zd+UCXG0ivpASw6kWAMEFnpJtFNCOaVNbo
KLHCxKLzEewJe5QtQOWd4Ni4zlImZOq8yYjP4DillnWsPFowRw7fphvL/NDUDNe4
RjWBJ4yhSuOeoCy5O87B3dycLJIvYFxE1i3Nd7Jqq+qPhSkwwfmbpYBSUkk5b8OF
LoWzzUY4RX2prA+hpER8nZ38vq54El2zQKwgaIFL3TnduAxVKwdut6HykpuGUUX4
GvTV8pXeKNJPoh1dp81yW/JHQQZv3KJ0E2dC29dtUwZeCMDgHv2AHW2tXDjPlhd7
VNG2CpAkGqDDOCoSqqQtwgmsZMI0JqTjz549nfDv3tlr7DheODC6XNbhTyuLG3rk
8YJto4bX6JGBtNVKk2Znbq/v8B9QynRme/zD4N0wXjjNELVJOCKn+KELASeY9wDz
scdoezugidYFC43zRzTV3HUzvXZZV5sMXi9BmxnpaaYXa1rc8nyiEwtN7Jv5fkys
a9T0lnc1QFcy8cpwBim8HMCsZBxUMlPKZA2oqQ/0jAk9CFDWFhht+NDqoyZnNsG/
N7NxjkZgYKW+kb1jRq6xGrSY2iGqMYI0lVvN1UrHBaNdOELAArikVdJ9jwtomouf
BSU9QwxUYEHw/bJ4So33ZqzamtJBfaw3typQXVtUWt7UasmPTipvVZGpsYUsk71G
xSOQBfrFushFQd5kXUVcKOTIdEg8QIgTtrfOCd+OJcJxQRzUGRipBHisLCVyyR3H
wAhxaTJ4xTy+YuCj5QXLIdbA8QP4/E1SiCswcFziDdjFp+WL8VQxZd+xFUhxcatr
pEH/+FUQYc/q2i9MTg1zt6XfNE1KURIjopTwpLI5ZeB49nkfs0Hj9UYPoI5Jo/IW
jvVFSCVPY4s3xrJQjlguGR+0X9eLweaabqTsdAzlP8/7LgAZi6cqtkbCnyDTwLXW
yPd81Lv7Trb8uGWNUMp+pfe95qxxviYnto5/fp/xyNToWSzmXei/yNKASPodp1T+
+dv+hWTMRcn5u4B9a36TZm6fX9GJAPrFNnYL7zGfkWw7tF/6VT6Zr8FqnH72ibCE
t3tvcfXnp8Xz8cIu4tf+rI2zYBvlaE65+2ObI0DZfCyMZphK5UPxP6aVXUABN85b
URPDnzUZDMtrmD4eoxx+CqhncEkGIsX9Z/rT4maZ+XU/7FqQ8Pzl6Woa4OM8vzzg
GYSJuc1BjIrpGddnrnBzPwBGaPvIRB+t4SU3rM6YJU2vtfbG9g6izAAsP1hiDKot
M/OQkcOmeM/hJ2OcAR2tKxgPT3Bdh3lZR+3Mf4dMXisY23H740l5uzPgvUuaLsKn
k0pmqDso/Eu52VFNmYLqlyd29NUmVKspQDrl8RTQdjpCTHtrZP3wBg0yqGAO8nAM
3e/N6X7c7ZqdazrOIQmZm8LYvVV4Q/b8kjjDxdhz/NLw8OOgH0raVjLyFi4eDmd2
tQq3tWsUuTl36Glg/5urWTh1AByARc6u73CDMQ3MBXWktRHv9QoFLcObbOe4v0xt
tMpXfLC61q4MkGtotWESSn6UUSdfXsIDF8joVPyB4Q0cButlm+/xSG6hIo7lfpXK
7UFIgXW7VlfI/nSaQ7TMpZ46cq9vDjyYjtqdYL5FKOfXfWXPENFX1RYxHYRr56YK
enNTtJYbafhTa2SYYzTojpQ1c0saF6hEV60K4CPzAud7XwdbQY7TKjuJ+NW364Zr
RU4cVI56jgJmxbFkejSdksT5i7PQTa5d+LUmBIqsEEtuEcDXpSx5cEDisk9qx3Qa
IIMMix4vlatQwi/+VtoruPF9sHRNNi9hHad2E6Q/99ZTDsrQUSQUczpb+3wCaol8
a7NJehbsEvH6+Tlj70CePvs8a7+FWFh2+z+JxheSTXEMj59bzU+lUA8dTiJOhAtg
eiLK7QTndZu1nTnXEvUvwXS3S9M+P4dDu4qSNsqpkATg20XGMLFpjG2oI9pg4vFc
y/Ih5ti2dW+Ll6hC0kmlO5gQuFg8G4twYnawnU+Ic7qptd4bhxfQJfe1Dnbifi4D
UVvaSgqEG40dcian5dcYIPxYX9vj23XGr+vT1Als51yScg+gPVTxyc+kXPWf43Zv
j50sU1Jsouf/tFQ81xW8y7RRvVDMI77/xQiRS5pIfz0UR4Vx0kIeCnDqmLqEcpD5
vv0og4IL0Q1DwRs9sBE3B7XiiQnVEbDaDuhsXHBbdBnItL1eO94GqqwRNoDD41x/
F6KeQHecviKQXITxqxVR0QKLorMZ2QVGcJ9KAc+T+xIr1jIrtgHSVPFy0Rls5cSV
i7/RqpURXYOoBCNv1IMv3jmGrxzmdHsfM2ixgDs5mv16FKoRnOLNIHSGfqMT4zql
2aFtHqsfpbslI00sAIw8NyFmAyh86tAFGxbWrr+ieXUvAAUfkopZSWyBqhixMiiJ
CbU3oh78nkRkATfEZ4Uj25c98+fIYMiP1zJQAESznMBgHzEZN7BJnblRshUBh7bw
51E3B4DxLW6ZCXSuokeOwfWd6aeqhJgWHDohagJpToPaM3zFWJhR/2Lq4zKOuULx
7vnins1HlhGJ5J+Q7Mi+cyQ7FLYND8+JA3CicVREdU3b4aLlTP0eXUwJ1Q3HmFUX
YLv4irmXrnsiaqvrC/WpkBxQ8cS9oBpAh3WIt7GnuvBs7uBySNJqQ9T2PZdjQaIR
BrDrRUu80QM1DKMRiCUgNvMAxthFRXol4tOS9e/xzMYgp0x8ZkrxD6XIgL1SGDhy
7W543vgRg5Xmq5c67Sm2Jw==
`protect END_PROTECTED
