`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LbxAuPJlnRhX8Q2bX4NqzpOTKduiIY+L2n9FkzS2nIMZkB2Tz1Dp7rCnK9WUr3E7
8QTIjeV5S8HmWykM5miLHxBoViaFCydpvpcm2n1IQ4Fy/s7oie30m2RSvM+ZskBH
1BNE3SAkQQz8lsKmWK6awACBPjHekvpwpLSMBbxpwlNMBp5Ypio90Y8f35Z3X/Yt
jEvHv/46sxNd5MuWzkEuh5UPTSNW11A10CLciTE1sKLZhm7ySMhAYN52d0nzcjbh
HHp+qoAwC8Lr/v4xyaNZGTULyXMZJpskqVzqAqMVlYr4Zp1YDAUWQqIdE4YxHn4V
qgUKRHcdln/qWpa4tJ6uLn2mHdT75nmC+qYzSHsi0bBPyu4DAS92UWfuFD61jU++
8IwGEQg4pX+MESXjjGxkTg==
`protect END_PROTECTED
