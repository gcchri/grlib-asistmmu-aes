`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BB6hDFdN1j41CmTBOmh50os3Agdf3kYAP/xibsSEsTAIE1ZypMTbL3w/wc0Pmnaw
ynsexzzTOJuG5V1Mi3KkAUeBMf4vpnLVP7XHRXulUgZr+Ag+lzzGytbedJk82zbw
BFyYQfXY70UrEG8B+DKv418yIrM6L8x5dE7yNgzSguNkbrMtLG6H5upIbxRv4sOI
iezssIMsKtysxgGnByvT05p/nwYd1mZfv0Lpxl5oAqXtyA3MgG27EWNAt/ShW//g
K8vYRKWXDGY1sMc4+zmFlY6yYh0nF0ewpI2DNZNTIybg1nTTFCVeiMpIXm9fSiTb
Al6LauqOTfaZcCw23KMK33npJxD5yuwWvmlhtnXWrv62fD7kmFC62elbGblgOHL7
oNsLYHeQ1IdzKYeHQwozL77BjBulidqObtAWUTs2NUT/KnaXJ9rxVJUvmTJBljqx
nFXJStrEzQVvIiFgu7Ij8jdHl9eERWJvKtPl7szpkqmOgYMd6eyAuC+q9xSSaiCj
fOoQ6kyS4A82sAKQAH0bOobdPA12my2n9DyAv44xeQPcgvclogksMpkIcjpdAcBR
7IfX/u+yLpgSwY+m8tvlRcMHpNBBJ/WcnGnIX8ha0GLbWD3s+zn5i93XPHrxHeQv
ogUUhH0GZR7bEU0OegPzrTQ1aSg2I0M+Wol0wOOinK9GdeYr0rNbUG3Od7qvOpCT
P7Rbz5MWIWZY0Mp9Iien0g==
`protect END_PROTECTED
