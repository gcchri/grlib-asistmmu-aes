`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypwp36p9ICIuO8D0wzDA5ZCrpxK3jRmSN5VRvLZlUq49DBtCN6jRkK/5DmMlSXMq
4Gt6dv0KHFAZ6nOwzyKnoLruUqJuIK1DoiHbBd3TwDEuw5fcdbhqrJlSrxw5MVPJ
9yxo28cuCwRHIczsl8m9anAZO7YpaMyL0C1ex2KBXeu9h/nN+Jy1k0Yy/EJ2UxRZ
5ocRPDmXZ2PwIcOtMVkzpMv8D2c2a90IBMjMxwQquZZVwgs5Utvb3Wn3VGMKUT2w
AtHTQjgWaX/3d1s/Rz3e+5vKWgKwn9Vqkrro/1DjHca2QOv8hDy9NIpcvBb7wbfg
xXF9fHvNPSiocIQjcZ3TBWMrfFLADWtRH41u78kNfjK5oFkYhDN0A21+g7rie4sz
bYRwK/buSMiDjtzccdKvT++UTMpKMzN9uanuKq4wjj6YGeCCisa5rwn+VPW9HgVP
nu7Fu7/iQIIgnz9Ax7GdGuxlNmvg9f5OsC7HR2kqla5ogA+Nxu0iYF7vrNAAlqH/
vJeqQhmGqBhBRZ36ENv2NLU7BwfIchiSzzJFlvtWORenaKNwxyx6DzaKfrbWEsXb
n0g23rEre81CvyZNhjocdUjj1hLckWXvuMTffYOvSjYqz0U8QNFE2oTRXbgcUU1Y
f31NAS+7TZQG6tuyXb42jqh13FAh9EazLj6+saT8va3cw8X4IzQD9M6pIbXki6n7
rKa7Ff/8MGdRBlIgqYalu6jlJEON7n5M/a1JlyqDAPRJUxqfCuEpsupCRBaX0+aQ
ks3wV2+1IzfqUis06b2ECnnU2gGj3Y/sJUQI2RWbRsjq+xbu9gulRgSVM+7mZdMY
0kWWUGSpOvn4gcwB3xcNfxvlwr4FugIVtnRnIKgVh4eVvw8ZQG6rnhgO6qqX6eHs
VqZ8Bywwja4Cd5G2RvkWRAencNpCUbQajxkIddArhVm8UnOQ9YhczR6eqSley/LG
pcYfh4URVFGlw3I9T4sA7aFdCmgxt1Uf3TeqIYePzZ8RxXdUF2uAF8WsYhhBIQen
vyUHX/Dd4V7DS2Ucye5QVRGTXKrCv4c1ldQFOcXP+lACoOJo1mu6JxeLB37mn2gD
LpS9UHyaYV9N3no7Ep+vugiOK0ClHSy6s22Tu4VtJt2D4yqEd2pmsF+SaMP6mqkb
mUMq0nAJL/l9TsMgbV6LHmw1kr8MORqVqeSmij5eUXg0X7BuHOl6hOBI7hhlLn3g
wVNY3q6p+FHGCY8tWE6Wo4lYY4b1DhLZpZrcjIwTrNj5m0m/Tcp85/EGAKPF1oqk
avJTwp0EyJAHTAPzZS19Sg+cVYjKvnnQeByEjavm8p+bIM3TLkZlgrr/bX8+P/Ok
yV0+7VYeE01Ahn9J2ID8UYlg1v62+o1IQCpmn5J5Tk9qcMOi1GCdraey9YA6XyAr
DH8gJs/QhvA8fgkgqKu4uTdnwUE8zG99mb45ObNl9WIOf12ak+a8RtFHdo+1e4u5
LlKvcp8Zfv73+WVXsz6KMankq2POIaggRKhZyog3jsJ9FjljNprk4/aNFSVRoTTb
6B0PSwh2oObrbnhI0E1rX1CvZ1PPLeTYn2Z1g0AvV8bSu1utahkCPzqnM7+dMFq9
u3hJFJXLZmjwFWGflo9jgvCI5aEENaGCs+7EkiEAauGTSUfWqjDKeJPDX5N02UQH
5EiJtIJ0vWAoJHUBLY1TUJMBHmsGdwf4UU5067aRkbzk+uu3STW9/dZMq7qu5H2g
PSOXCyyVXEieVNx+4fbMyMoDVVsmauoXZeCQV99fpalI0nP1d4Yu4teyDQdPaTaO
gym+MvXGAI0+hrqk8v24we+Ix8reYkb8YRAWzKTdLo7jxdgWSktCYHG0YQZLZRhx
2YxU5nbayIEYyWfrCp1cP2MW+z1SZbrfLXhPrxj+sp8B3CiFfzQPNBAagrapnk4T
dUYNHENc9Nk67orqUt9tGXPEYq43y0A5nBg3goPYMMyVwIKsz1uZBUU3jOFpV9C8
6bMhvdyzq5XdZtFVll09Yji48ND3xwYRcfoakEmC3l2hz3LpMtmRv1GTNIqss0Jq
MKHjvoMOZR1NLGWkYuGUXFcI5+k7J9Xdht7S8RiPLo+T7xAOm23WkyR+rzJwzNuf
6HY6JKR3P/+W87DW5D7hz22O6WJD+kXOBjACkUMiZLeJgcjG9YWpaUF6MXZ2zlj4
EvqKJo8foS/OeWUJKQgcVQZ8J125R+d4Q9SmrqJy0iami1aB2itNmd4PXgWDMbIp
kERgGmCFcs73DLj85Jy53CqPjgxhmLFW0vFDLsk6TXk5EgZs+mLDGpP21lMv8ReY
WwVdXErjs1e5Wb3l3ejmkQfz+YLfUzM7DPlH+At7oFvkGQD+4gEGcFluPWtmuF+S
wvJUKC93h2KnVfMI3uv5kQoha8Alg8eYFVlJu96LLIR0B66ZMSMvGEhq9ykQPHj2
F/IPejW/P/kYxznd4GG3Ia3Pe4XEFb4JXKYzvHcTvvjEnMXMBSQEin/esvR2P4C5
++BwnOmTTUt5BesnhYOamKmO5ITG5O0jTlYhxbwUSPWSyxBOkm2144wS8I8BAOQ8
7Przrgi+iDC8DuW2Uw2h1GTtA0OXdsRzA7G6VEIXgM2VP1c5JsRjKJVGTQOe1gYp
D74h53LkrDTyZNxFLca9cAtjB9WVQYYJWzeytNhcaAmMQ6H+vss5h46zL1fj51om
o9CSCeQK0JwYbjO/5DNQXi9AbDxOVe/2gN6zCULOjg0qYYa9Or8/V2HapEjlCq91
vJPgiELQBr9yoYWdptbez0cLxdg6+jC4+mmTfl+hUnx9EOiq36/YTjcGHQYFrYPh
UiwTtWaFIN8FpmQXQX+rw9xTXjQa4LBnUn0gaIWbd3p0RlEm+8hChg8OsG6HQy1l
taHuXUDhixp2FHHlXDriPkGeRVhNpyVy4vlwD7ecTHAlqlS0L9i6qIcd/BLJfzBd
ze10qRAY0XTsasrQ7teAiH8cAKXvvjYMjJYWLr3/caJEFEzBTEGgfl5CglxQ1+dU
YGfPeab9oNhUWubhIGQCJDcMZQpNRXIDCFnESUbDRG1+T+Pc0Kv9wS8Gs07On1fy
Wigdy11RRsOo/Ec90VD6dhIlfzDXHaeIWxmAQiRUfTNe+yMfb1eXgmCWjQEPX7dm
3hv4Cq/ESoTLezPDKuyYyrh6d+Xb44XGSc9scu88WEiWdhYGqyFPGEUFx6aul0a9
TBIVBHqYLeiA0MUUR1eytP+dTtVUs/WbaO9MA6qf2WrPHJ7dZRCqSvxvj4fmzAPp
PjpB4PYMzmLXSaCGlkElkt2JKGQMpRFf1OM8oEOZFke7VuTt+bdrtIUyPuzf8OHs
RlT8NetEY/R4t+3Asgg7vrgKUHlmqsAEke0dEMODIOnsnmRpjfBXA3KQeGXYa561
WzGw9uKxM4XDxWCjpVFdevubAtelGbnXNSBDhQOEF9FrGpHdc9QiiXN+t6XhzwGW
Je35o8xsgEV3II24TP5rB3MwO7Oo9RNuLbN/Y21kkTjEhRZrstX4Ut2yMNLSqdCx
71vBAx2dCPLu5gIRmU/6/EwoEC1mSbKyHGwvFkdST1WFo/RqbCWdYPijSRJTogO5
tRQf9HLru5m+gsjXyUIdYjJgieAwP2I80HtCYNDaoPuWdUVkhZCm6LiDLTazOD/f
Aw8w5iPSDBP7sYrmq2od/PmuYoPY4vYzmL9PUW/KTdKuyCMLxaRf6heMP1TmbVlf
mpPwk79qJ2BTbA2/ICXNGQ7nnN32y51pOdG5ZixplQv4xS2HzCS3krKH5rB4YAsk
jIuWGbZb/xpbxuT/fMaTSk/+cGZRgMRBrEZXpVTsJmB9ahrucpgZMwIyKDxiJ1Jz
bhXdNfPLSJih6JFunZzJ30y1RElIfYtIXq2Y3jCtdiubSZBuQIF2w/f/31pkrmC5
elQ7F9xDvUUgzkAEcdKv4K9nUZVA6XN04SQzFsvca9OAS2KID+nBP1IRnxFkURFQ
m+/paqfe9aqDx4mntCCzRqfjbCFrpM+VZ4LZ1QhdneS92POPcsWkthrSp0ryigrU
P2z3gbPaRjNUYk3jmwMkbyhkcvbvbByJJ7XvuX8ruK/br5oW2uZ/0QyhujCP0aZM
1/DGf01N72V4m9vj3tWzKOqEWom3b3yYjsXwiZK6FNbzpzvCHgQ1dsTuvfy79LL5
wyqTB1j1F8L7/9RMWinj1MKTezQ6S1F/BoXhj9SjHSloXCQmlJP6DZvwcben+Za7
mWT3u0Noo7p+sIjgeV8Ru5AVMc4+NWiYR6xoDfmweTZmhXA00caGroh+mYyubhBW
p7/Q8T9XUp2zQU/Ii39JC/TQ4rfycqwlfLnizTEapEmYJjHH9b7BRw2scLZyfsS4
YxlxJ6U0Jo0SA6BZEfRlOYif1BWMZEofaZPvgNm+wKRzW/JuI+9vrNxNacg6JKWr
zkToAxIwFpT+aEFmJDyOkaTyk8Z43KwUyyIhHfc8+wbqHIcFy1g1ef/vE+Q2p+s8
5yvQl32gO/EBRyfOs280htkgel4ApcuYL3vrB5/U0KL84zHmAoO4HZ3oTLLjKyhW
Q6xnh0N/UIqILYbp4y7TMHg/xKYe//zueCrYXs5Oj2CsPut4u++cKaWH2Ksj180Y
/aqZMLmHN331hCyYUsw7dtykiDvwH2ayM6Y5lDhbxYWgsvgIfkiwZghujJU++a/c
8GkvHuTp21cvp4c9xNq1Ghg7TAoY/h+RsM156GMMBhdoU20CBTinYrM2BWQ+2SRu
yt/8oI2Fl958HbnWT3Bok+UmDaG+6bQivGH8h2saRASEydGyYLFknrmkGfHygg2Z
6LvHEVa5PohXKwmbX6Aqf9HXQ3ppo93qfpQM19ZuCRrof0B0vy1FFsgFI85Wd+r9
AzyX3ydzQowkYMdQGW72NTmc54OilOiOhBjSZM7tY9kvar69ivQ9LJ+5uPMWnziA
emxsdzPejdJvXJNqgD8Abx2EE+LlcjK+A6oJbkMNV+KCB1ioQxBEvbMeXApaGnqv
CZnFGScogCW2UTA191ThkixPORRtLnrQhm1I4yoT8lM=
`protect END_PROTECTED
