`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DlePwZ1PsPkCTCaEhWsYx411DVmzuM4Bfbo1YWsWuYOqJhdwtK1nVX6rEOSjh+pk
vkAVQPoTPAmLkjQApzu0HATdNBQ7D31ErsLwpAiRVo4APbmko/JA4H00GnhmvACu
123JMNRG3oBHNC8m1PPrIDD7ef4X8XCr3Ka5p7JnGi2xiJ582x1XuIIHvP+0r9Cu
zuhfQUzk5SgIQQSeYlbqliHzAEbBYuNmJx745bKAekKiu/m5i8toatqdjSWz4hIp
4Ns83LNntibRVHHmgZ0l+rbKbj7Awn5P8kBtjrdjBZRaIU5sr4+KwvppR4i2wo31
8j7uLlx1KnmTG6YD1sEYdhvAXYeJKCpaoZxB7xyFKmRxIyA80/XwbD8V57/NrlvW
hsSw+Ojm8rdSugW95ricbQP0+w6G1f8Qd4c679Hru4KevkTBkq6TBXtDWIVwwF/d
1twDn9wJNou4IWa4L85BYK62GHQGzH8cUOOT5Ukre0m2USFA9Y3yijOT6mjcz8D+
3X3oXmpRk3HqaiOe28RYEJM5Qu67/iQTUGwuSTN3EQeYwn/kBRoKU5EteJogz2jN
C9P/i1Uiw3c2xuRcxvuK7Ev/fM6gMCPWJbubr8awMb82oOFDiNNzaDN0KoaBx7TG
Tt3RKD5HXe9MpqOlBUNk57mvqARMAnChKDWhwB6dIeljM3GJaFj8H0A7Qgfsauz3
Td0ycC9fq1IHVGo6f/vYgoQnTqG/RwdfB8HY4CLyOtLz/SaTBnPDP9CkT8loPWa3
yDI5JwoatjvFTZy6MZlGynvRct5tU4Un4dSZiBWvmdj4KoLVS6L5XRfxiM15S3Yi
ot5S7rW0IBpLH8TlFD50QoAQtdvmtfNCY83T0m+GRb2rw364XHsiLa5B+MeUYDv6
LjWcSrdujIU8DMh2WiM5IMSDtCvSt9v4pO7eM6QwJ9U6eL8GmQBuHBogJ8U/GrIq
GgbHPrp16ORgDTn575PYYLlnWUilc8BnpjCqNl7bJwNWH957N2DD+iSrMhlOy3kO
dflbl0qqJeQaPYV+uWYbRGf6pxyQAggXNbA0GsY2qw7M+xNZy84wfusxEE2/efq3
82IW7gWOt3ewBiOnCu8B+ZTJGHL1J8TXSNG/mQxCb8Fkiiy4WvQlffTe+t1Ja5WZ
yHRK5RTbJlIli14zBitGo/iaL42bBqVP5HeCLdmqGBjzfomcUyEdSjxjc8ULKgRS
U4aBLHNYrHILzeOnegTMXDppJAebHtIung2MxV0WKysYlMrN35KryYuzvUykmPlg
NhPaIAm2W2GD9ZZ+03amHdiFnruCXkU1Bq4hKJd3EimqJF1aRH2o5BxjGACQStFY
UqdePPXJAcWLSmvQRjkou7532xGtzBJcuxEjl7LupFqlMDOl1vwm17BBoiUCkhFU
8LB1smP3+ispCK4scNJlGA==
`protect END_PROTECTED
