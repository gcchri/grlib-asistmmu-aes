`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oyv8pKUB21ZuefWq81HcMauQHQEzaIKqTdNX3cz+6zKJmYMC4GYGTQa0rMKbL2Qx
5ExjliMjHjYDRkNFd3ZxU+q+Qv/468upguMiMUoZIKT1y5YDNTMRUPNHRWIMcGK0
0lPNBe+3r9WtA5Srgq+7Cpzi/ELzDFQjUc1/O3dzmq7gpLJtYwwlk4Nz+WQOA3ou
W1ksjt18Z0Ovz9ue44RXqrUuCRLVkGfjyk+yZtRBzrtjEQadwAYtdulx0Zl7PRJm
Uvl5zI8qBgQ+wu10Xhq++X3RmtttqqMvgZIWl5FfEG2nngpiW0SwC5q7ASIhVC2B
A6470AAcj2FzTzW81v2QT++JHZIMfVkhV2Zo3hlWhXNBJckkDnvSdi9P9IW6DASk
48FvON3/DM9nahmM3AQikw8PGCHCXw16bCdurxnOI9YixsUzxsueUguE9MjRPDj6
3pa/6G7pKni5XsY1AuHU70X4WKYfpqvF/GqDEICo+UalMF6hKQ45XN/dBZMcTnMR
l9j+50zauX9PbRcaqYRmcecyZe/coDNehkJV2XYp5J+tqDQbmvy3NAKbiBY/3MQJ
RpoWARx6faMz/Kkm8YRaREZQ8UYfS2B8mqLaWWcCxxKRJVn9m5jKVkvtfmY/A4A5
dbs9nynIcIX81fLTlBEzvOSkZLf0zO9MPaS+r3OLLXxD3vcNT/YLCwtJinHhjGRp
pv3Mj9DITZebMvHRoSNNK9G5mXmc189Fg/G5W4e8BL1rWqxNNcDnauuSqY0f+Tdj
0sJcG41KJCnSZm5ufCmrA/Yrv6viIy+qgPYwFeARvWwBWPiMaRZFvCG5gIOlzjHy
W+01GTCvX/x9z1bZ+hWEeJKpk2o4Vqs1x3iFHhmyW6xoKOzhswQTVQG+vDH2f9/s
vKTiZsj9whm7IrzZRCLlgIyyAlqi9Ip1HGrkO5vqGg+zOKJ1yj0hFrYSMEn4vtf6
P2qwguMeTtOas6QoBgwaaNoZ2YmL2TXc9LvjC1VCnu2NshWtPQc/xn7QjtRzhRHC
WtxAvosWUSL+UPCEGzACNFRdzbuiKcaYd8bRa+8+hHNQI1AagrOdlB9GvLZOaMut
WN1d7bg0b53Sg6aDu3fWv6d/sx1nHDUZBqpaKPqRZR1fS984Fm4czOL+RK690opv
izvIBP2cwvC94ZtdcAO/dI1/tkY9dJQ3jADANCgCgu0qRRIarnP8+QiNYs8zZoUp
78ktXmAS+8NlwqHuFViwv97rnT35mTYshN7punPSqtW65BNoJIWHppJO6GXU2UNO
V2gJjAsS43wvjiVFA3pxFASwc641DuWHEgwvVFexbIaH0+AkTYbVZoVKQfjg9rPu
l/21LEI30tA10xEBUJ1YqV4SyCs+iYtQ27hpj0LyzEOjRPEkcp6hUOUY6UzZrlws
7Fnfmfm6zeAb/eI9Gh9KzE8QYcyKbyaLcXENEGKXhX6dYcA2tW3bwUFwkGaEhdh+
GRTYGr5lYAFM9xGj/JRS6vHgWGEzBc1fAlqnWzdoQBreHxOsUyeHscaA0nbmEC0V
8kGiSt9w/Y+53QZvbn2UNO/9ZP6OHESZntRpzwuU3xJRcp1/fg9atfZAWdDC9q/s
kLauDPYs3oHGjzPqv39exiVIRb90K8hPYmhkpEmytmUVCNCLnz0Oasmlgm8l+MX3
k1UizRDrMq7BlgrdUoE+TQhGEgPuE+coEPCQwIS0B/VxohIvAel57QG4J0C+ZMcx
OU7a5gshkhckRbc9CdNZ8wPEXDT5KtlLm4zCSYDzAya7OTD4NNRg9Mtj+GUG984w
oPM46iiG6YWhzBfdZZk/AkduM8h65B+XbfGJ9qPYKzoO4GEoQD5FV6ECCYPeqhwP
AqIdVkyuOokGxWz8SIIgMlDyojdjGdCnRIr6oqcmI81LoGq1zqPck1M4phD9LJur
L8EmSAxeJsfeNTQ/wB0SdQ1wd/zmrfPFqObUTRSVtXZFJdvhT07QwWj2bG818HFV
3pmYZxvvfjGNsoKBg+3WcKDKYFgo0FP3YlaCd647i+G0ktpDGIq/8IzBSW/ZoiZb
r0MeCry/iZsBPgYHls2M1gkvqIDa0B6NX85oFGgScwNwAfWwf9dwmaJluKtvaBIa
VvyiXgNehVpFXHno4WFy8dVPe6SXLOdN1T6IjrMqemyG+6kmC1CdUNvj8OsEAcWb
528+Ov/STJe1ubRtrXdFD/JXRarIVB9A2Ct7c3l2qUoqa1CEdTmHY9RkzJlGn+gX
+4JpAzAkT9jioRRWAoZU/uK5/b+NCOA2JTCoiK6o3a2HLY+vfbsp9n7HfUpynqWs
jh8KCX8hM0Wwk0kWuJD9bvJFLGyHWcfOWAOi3mp571YVei0R++UySj7gHb+m8TJ6
w4TBGnFIKRLxbkJtLb78PcnXeczqcJpnUzqWkjU1qdRs6meAxYm4bacQPIMCQL0m
tKXX1jClulOnMbVPd88WWhaYm7vxzWtHEZWm+ocUQdJ6Ac5wKRNG8kIka+WJvc2K
vx53+svd2lbQ8sfnAYhPzJMaAWcjvklQWNu4raFheqhSbh6JbI21VXPmQL/iQJ/Y
2mJG4/Y2RqZ/GFMJsOPb0AkHqtm7nMZaHYQaqysxWs80TLu53JWeGfA6MnOwwyKW
+V06MgdZ/F80S8L2/ES2OFTypgvZySqCctTf/AVYF2m6OqH7+ZCoopyXtn059OMX
HW2woTkldvmoxqM6FYfDv3aQDzoKaOyO1pHhVUmKzBFBg7WOCSX2Cg5b4sODnw3J
ZTiiEUZxV6tcLaWew3ZKniBPky2ulniyiSHMFh8qv6Cv/CgOcwPZj7LINwxjSXpr
Ojlfx5+NWUEQB1OGYO+hwCl75pRjGsO2ZcsIUzkp7sqxMcgDSx+lvxpwRAFAhE3T
EsVV002Aqs9FdNI2axSVqHjhWi9wbIaat8ugyjjRvv+UiOe0628znNScwilTQUxa
qeB+AVQFcIJIRYB5qUjcL2L6UG95w2XJO9UcoFZghZ1liUHoYVjKm/PR/aHdZTbE
pnuUBnihH5P11leWGVjaWRQXdDIHCITjG1FZ4K2jypybYdyNgM8Pa67rXJdBVH4B
j0GBXfo7bGEvKOGfBalbJJlEFPHxgMY6eXPTDTqv0bfQN/8UlSXUYl9TlPc5fwzr
ub0IhEudlQmcyA/YDJM1y+pRGf/aa6smeCGAY7udRKT5zijV1t8H51u5pHP4pZnf
6GSufzf20ocBukSN28bIZdBB8B8hsO6E6LKudzAE5cOFIVXQO2c17OqNaivlqbV+
Upkr8q/966grFh47nVK/2zfWeRYMkJ1q5pJPkZbJtjoqg55mQManZ9crtpDhh24q
ItpWR0ts4oLfWmVBj5oJmrNJ0p68aOx3N41iDbs9u1pPdsNbaJWFZ+uKCxK+O5ye
Qk/63O4A3TEgNhEzcg8WaZha1HBQkYNNCMfNuOAp95msic2OULrMnwZenAAxDiZq
qf32RGAa+mcEsKXogwkATWHp1BYfbquPadK7/A8BLbqpuUDKrAK+Hp7M19I+JJZK
jwXmCbf3crRP8SV8C02srcvphBl36wGQtpGnyJbl9c6QaQS1CuE75F/VgOsdzX5u
2VxRvMjeiugYRNGDBTnr2Q+sh8h2EwlsUKmlOywYMp1Vzj54lRkk2FTBjZEznwjg
q+WYBC9A0EIH+d2NTaEIeet2hZuaItPqCNkArXgIHWkx0z623sSCRMAKsrIZ/3jn
vaiND5WiSShxW2xnHAoIqfUFomjPxascoHjj5NUlnQSOq5EWvZDsFZfyrBqDoETv
5xmkLKylHWz2BnuEOFvtoxYknarT7E5x7rsPvh03Baogts5YrR8L4yKdBwxYcrkm
OZbVRHMc8n6UF+RLCkGvY5fJAptHKoYiY9BJ5PMzKxHvdBuu0oAayea4FVxbb23+
9XRj5Kb4jQXyBKHCzJsTUCDaY2DclJ1awYLIQk3DsdzRu6RkOSTw2/kvSY/QsYam
Qelv5+KBv9OzV92miNcNnX656JxPmm3n3fIfgrjesZsj8hA4W5wB9jqYAJaX3M0U
gE/QhJARdm8JG87P7HWqv+ppMMCQt2y6mrgJ4Y/rwukJrfw0+jeRjQ6FBkSdJUjP
W0vlXroIeX4FoLvMpES5zhBQOGnRxs1yU28TxrwmWVGIltC72XEL+KuJONdnObOx
Itq6yG6C3umYSeNPHh3ZOPRqlXY2p7sLGG6NdOc/vziECwt0rHITeL5tBnZnj2Cf
E4ZNT2zK/2Xiwe3hHpkQBGkrp1HJob6j9i4I4A3Q2ThGR8hjpZUTsMSbKltZ5csJ
25XgNxnu4Q7WxHkmf9PKYMTEax0lnTwTKpmqp9WudTL4iS0Fi1Ld2RwKuSwK2JG8
dRlEBVTtqwAxnw+CoPb0KSdbYvboxf7yi66SWjxYplZbeULB8O1w4nIjIxs7U91O
zRv/pTGrTcow+Hi4FF4laZ9xOrEqqxtSPrgZ3KzoEsh0MHnqvCgyn60+yM+2g71H
anYYmrxXXICVzvbQ17yo8f6JKogpeMbTM3QakcgoH3ATm7XM/L3Oy0lX9m6fmof1
qqgEAjGoAmc9KUsWpyEIlY7UcQqUbaJnnkUWG2AtNspaxWcTD6rkvNlYshO4wRrY
6bB88QFyZ6Y+5cvjzD+neOVlIdyLwHO9V+4gs+AJMXjpfqyOZWeMoYp7HOmk8OCA
`protect END_PROTECTED
