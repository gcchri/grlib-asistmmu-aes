`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nonJyeguGMKnokF60IleqKUeA5ZmKdclCc/ePWtuS7Sv4vBAN/2xfNYU9b1zksDB
t3Hwo445UHk8RmDQUUgpzoWoq8saN75neY5pNZU72+Y6VJ4KnJbWJZSSgBNvXxaL
mvkKusNAfPF/uZ0/TW9XwrpZ44bp66P9Klpahqig5c3gIJgwPEMnmvfiJ66sp04T
luTm7cVKBA6/5zhgg+cb9kZZaCtCKBx2dokI55W9LdBXeeEGeHys73rpULhxHFF6
XQvLI/Mt6sxssUvFrpa7GWs8jFEWoTsCRbcG1YrKauyyPy5jafMdio0koip8AYc8
gdthOTTLMOVfVkyPvW2lvNzrMH3X245dJv2N99MD/zUcmmgl5YyUbZ9oqQJlEdRy
aO4avCVWuAbZTmJDewWbSw/oBGj61XG8URFPu0I+RSueyk0YtYMTOGm4LzXH5DE/
nTnojZbb1ohpQa4SvNfYRMPOmoxQ+GA8BhgEDgOSmoAmiD1HTWQv2h+ugPCw/P9j
bP4QZRFHVGyJ1oDvSu8Au0i9iuO3Bq5KdVXW/tbQ/H1+ed5GBrTSVieJbdkaTWlt
VJnUzX8A+mo71fk9ykN75XpXMh1Keu/2gepC848JQDXr27mckuB/f5o691GR3z8T
ZXSMNW3E62XlEkTYN8OrkbHp2i3wToYCgYFZj5Z0MiM=
`protect END_PROTECTED
