`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ww8m3iUiwNUaScP+oAruWUoss56Fc9hN5mt0cn73Zeo522JqmHKTYZiVTsY72LJs
F+aBZOh2LhgwHBvwS825IYekuyuenk2cE6zop8joybUrH3Bkomv5J7br2IUx394H
XsKQ7TlzHbX78JFvPlNfbtLXCEKZSKyWDfJy7mceTB88wQbHfQqyy6GSkdDzUGlI
MAVJPtwyxUAZ8uPmGmdhKRyn+BjrGeMJpINVXc74u00hV/BTBbX9icI0obkRtwR9
ndviOFT81G9onC0/uW5M4sD3QWWMcML7jG+4VLiJVEfhsOi7uxxXQwAzVFGLKa8f
psZLYpO9SP+lwXUcDA4RjkuMxLoBJVY4xi2ZhcjoJDSwJ6RZFIBNd6ZISolaVTYG
COrQKKGYbNw8asLZWBCKY3tWRjehYoCXR5uRc2Gq+1s=
`protect END_PROTECTED
