`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KX/KHAXkM6w3MPhomlqpXZgnP7JO6ONFTSyev+g/3xY9zSCMA/9xsReLc0NclaA5
cEhmIIHp3+ikWg9oCVe4Y6iJDPjVbfPRbbL/LDttSEyysjZVwDQkiHf8NIlt7bl5
cwOAHTmBDCZ0tTrAI06ruBvQcH1UWCiTdHbnsO9lLIgWC7GpTwhu7X7EOPglCfgj
q0NCKfmBlsRk9R9er9jpy00vFP3frtCVLZy+rOU+CpyAvgNMZJ9sdP5BCGkKh4va
W45gW4u/waowJHObGm9l6Hu4uZxcEOrgjqoTjZ/f7qDkDmCLLs2pM1q4V+78gq75
OuUJ30xyZ1YKr8arf2FtAuSfdE0u14Yk4HTR6zgWkDc=
`protect END_PROTECTED
