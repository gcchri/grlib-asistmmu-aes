`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWmzwq/NjSp6rikDxAQeYItUMpC3x2vQvR2lCt1hHXDmt/SSLTRLi1kGIOxeIE+3
jfTvLo+pWp2XIpUddCcOuEohbGU64pCQZvH4kPfMQxArThhNyveJFFZL9aRzErL0
MefCGTDDUvqXOgXTDA1JWuCYZBG0A9XifdpZcbm3Ub9pETDnuwJ7BpfFwc2RPdIh
zu0yu4LA6N6B0MnjMPanxqMkF/hhx3lBbVdfcm9d9y8WTjCxEjCHbqp+Us/TKWnp
yCFIy3zEcD/yjJMpkXlBp1ApIjyUp9+Nx0yMYgwiND9ID/8d3w7c18WQ2ZEfHPWy
wDm6QmFuObHYT7zs2M1HNLUyAJRO4GFlfU5MvTXGIZ2lat4aMd/IQbb0T8zQNLlK
Qxg/d2jYL45ijEUjUl9bGSCt+00X21pEf/PVgU1HqnOAfBHjYOe1m7d3oN2QZBqi
HEJTzhmV+pvmvrn1VTWtm03yRIEM22eIN6dpmg7xkD+xaI5WCHOduMEOU+JtBrmJ
4duu3xq4Fo2GnzCiUPPjyLpWsRRmtpSUMdoMk9/fRMZNDrS6ZwWrVykCzHpUOMPS
fovLcK37dC4pdhy/7eEYeQWDAHPabrCUK7ACNmDjCzPLtPDLEeI8i7IwnuIgovF2
iq31nwR7nnnt9DZGM89GC8k8j9BdLAkO1to6/wie60ZPVb2Qoy7a2f7ImS7dpTEG
c73dMh2hxHdLa5AYXQm1E5qldJBgZ+6Lo4NhATciLso1SdBEZIyHezCUoENHo/bE
80i8kWqGsFfaTppwhpE9TGVBak2wLtPhJ15XX69oZ4Zvm1JGdThpmu34fCGofYDe
pSYz9+4JP6aTRnv4O3XFwwb3FL++NKgcZmRWf70+q6GuZ8JtkQOCc79si+78qe92
RrysQV/8phK/gNOt4wO2kZdQXSoZLd7BIksiLg5a7wXi3PkifO2+6c79a3yjE6S0
`protect END_PROTECTED
