`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
avJtxF1dD4jE9zue4cgkQu6/SRq9DkDbd4/A62HIXgFCbig07TZ51Qr07wUpfTLn
K4uPorCheqKlvmIxCyrPvxDDmMYxj4tlDhxXCJZl9FGhCIBYNZQBi5rrsNciQCIx
Coo++SSsESQfiJjgJ5LfBr96gGtNHntu6o4opQUr3o4PSP1WNuQoxCKRuccw5fv/
16uyv/dsAACJaJGsrNb6LsY8CojKjnWQepadd/reZBx1V9f+kWB+xLWdZ2ZZyY/D
p/wPMbeAUb+WFP4HyF9ytutiJkg3AAfynvlpTYeR/Nx+bALQ3M0hhZBUz9RnsspP
vLnPWfuLJImwTmgdBhfdXsEcUCP7RO3PRHrt/kRaK4zWdixyPaEfrWe3aIpMcmw7
r9lxEf7wau7rZ/DaEjh0t4HzIsMkFVk109zwdxeHAVcFwqBgvw8u0tJTGRnHWtPG
9+ONHHOuP0CJsg5TLaWX9Who8RVB8tiMyNz2Wt2fzL01D5UwHKt2mQ8VMMd6CGQC
h+SbcpubqSw6ghI8higDx3U94aiRqa61azdcozrYaCiz+8kcgJIdF3LOFmBfo4gF
`protect END_PROTECTED
