`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJgyhJU+YkgoIRv+jLAFobDeKz0YtKhCQiHfKZGQBQ4iIFPvgKFmhe5vFuYJaKvw
N9VPYpeimnC6rGixDdkA4U/N0hRvLzsNd5a6aSUca542LnNXbIVtk+VY/B8vYPUe
zulMh0n+M8GNdhu1EkYruA0f44axsutxGLyYEpcMyqvS3UYjoyKWhd34aq4nLPJC
65gWZJyMCnTPjukIA7EPjNaWC2DgPT5QaC1uAqPWVRlefB449QUGSvEcIHxH2x0y
Hp3MV4oQ3pXBFB/c+3Gz0Co0aYcI5CHhlQ2mRnFu7dcxlN0DzBZ3tFtNrR8xS8Uf
FilFbI5VvPrEpQ37IakvGg==
`protect END_PROTECTED
