`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+k5cCyQkIdtELQh/meY/ngek571GlAxek0cTUHbw/EE6kwcmedk9i0oiaMxU5VZE
BVvJnAKgjo/4p431PUHMRy660kNEC9Lq1gK5jYyOSfZHrMB/3s1pNeUBkxRM3of0
JhW2N7NzvfmBm/2jvcdUr9dwv0S7DRIkvrYRqeXSA3qmcrjRqA00UAD6LeMC+frw
357Cq+pD95zJJwHkGM3F0CCzCB/zMb4U0RrtOjoCg7jPE2ppfVFCqm9LiQo5xGPw
tUQj9Jug5CDn181nXyblPSQDdH1/y2vCToaNfMsS6I8v7o9iYKCB3lMlqV7cdTLp
uy6EkJXQWbTonwz3IJj9tYP433XKrkJGumk9V1urWwqGnm4C1Ib5qUHnDGgdecKJ
PkzFBTcnF+9rpq/3i6baQw==
`protect END_PROTECTED
