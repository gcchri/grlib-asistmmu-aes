`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/8OrWi3vAV21emtSJfJRVH8xJbj1p/t7o3DxA72M/wfFXUlPDzchmvGrPNtLZs0h
E7ADVJLd8rWKz4QV+Txaa4hlcJVPcMJGkQIROQp0IwjfujSrnHpXlRK3XegAlkzo
2cb2n4rVPb5ZD2qyfphXz4nGHsyi13tSVaU4slM9xvh6XOU4X2SvmGQfhK89R/rV
Bc/S4oClNnJxokXBdA8esbJerQLdvJDtbjjzLilzsv8bMr5TGjxSHg4k5LddYUoH
I+tNQ0aJrfVNwAmIzP/eHds5Y1EUWcBba17vmQ/JxdVPBMX0driZ+AAfor8xmRCZ
DjlKM1kv08Au6mud8Ilr9KwD9h/MHPpF5yNyNPZVtm3jRJjxbRs8vLKkEqBNcIDE
wefEo6iTZEeyxq9bvVPIvKRBKxs69s1MT9vuTobbDcLoHShT43u95LVAeOa3kXSH
e5Jls4PjAnfeqlp/GcxjK0PQ7J37OwhEBqi836Sv5AnaVeghgS2oYDKa+x6MFiH1
u3zXpEwXdPOWD16qz5GI4doYvQ1mZ+KoFvp1EE41vp2GqHXnObQR2G8HIyKrXXyo
jENJL7PcCPAlblihuaqU/tH9O87AsF66+JhOqEtea3xPeuGJFFaxNm8GeqJhG1fM
`protect END_PROTECTED
