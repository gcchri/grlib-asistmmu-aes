`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oNtJiDit1eOJP+t0qxubzOZMGZ8mJsSMDarLROZP5ayFbejUxH3bbYbrOdwZDEtw
SZqEVbhJF2RmtaPHXCs8wMqOa9oqcoVkUfXXR/9LxvrVpdJlBdclH3QiJajNiPTm
AMWpb9A14WUGRte2kijuwtVRvXo3eB84+r7kiLteOhssE832CtwxDcUMXAtgi6aN
mpoS7MR14sZ6KwmWyDUT1Qrcf+i1DPCqL85T5fW2hE6LTwmtpGapItORcSrnV/ic
vcETjPeIF9N1czS5RBkLUvIP7fU87UHPf+GbPJmAYxUEV7So7/gJ2nuM/wO1rwKY
yUkG27390nUdPbFJiFwHIoSdPGRf8A0iZz8clGtkeRPLnT3cQ1FWIinOI8gvNgEB
YVnHRedEDLRdWhEzsUnTaDAEQ8pmHLGahV8jkmeO+S/ox7a8hZxOhpzNxtIx287A
W6T5Lcn6U5DV55+pmtnQz8E3XvxTUqCsiHRUF69kuqqlzwJAijy2nfOl1YYKOoyn
qZGibKM+BkHcZPSW0KU9Lz8T6xxqU/rh8rWJrJAUtribgswRS6+qsr/dEKNQ7Kbg
+TTtxp2Le9OLvzWxBJjLnT0pc1wD2R2FyKt59IIcxuO4KtjXq/VGr+wcFIpSOpda
eEv2UPVeujcZMJANqwlghEOpXCD6QSxQVHoziCq6SKfiOGJd9gxVMoSU7xkboCov
CvDikhoKHz9NUC9P8Bhw41PZ/Y+Rd/oGSOl1CuuXofkh5zIDh0WEK3NcWpw+jrna
MPKVlFdO1tO1eSo4qt4t6G9wRV0cXOperdVQVOmNJl/enu4PkBrJTc4UvXx9o+af
TXeXnPYF72aEpWoaBXTWixbxBt6mNH06s1C4PFtV8PgE7Ub6hZOtF15DPkdV4ZG3
M/LNSQYO9WAc5UfQs1/BVnvywZn7UDjQRfCTg/CwrvJsbbl5j25T+m1iBeutEwUZ
X7ytAuzgKPXk3SmX1k+a+ara84Gpd80Rvj287Lk1jMk+7PVDgKUCCWlZgFUjoL5/
KWbfiXVbvygCQLU5CPimdfMAzTJY/9fIH1bHx0UFQ8F07J/JvGEBZDNAJDGlAIgV
kPQMtJIc09eDxNPjGezhDYDLiVVQpKkdRWnQ55X9MDKN1HElQuMLflmzTgHkclxA
`protect END_PROTECTED
