`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QxzuouiJyzndIZC1grHlFudQ8wdz3aZkRfI6PWD2xDeMnS2GflQ70xBNyQeSAWDO
Wx3crnKtiuT+mWonyeQ02s5HXkdUlEgW2FWfJLOAvp6TE2mVvCoD1FmoH50R/4Y0
B0B1X41xFMkF+RkFfO0wkkGREGnnUmUXoswGCpGq4j57ZK+ZTuSAu7cy0bWSZm6T
NrJ14/VC4e4LdLNVOjWTBouSj84ytqA2CGWzRyG4jNkq9ua+IkGxksSvfA26tnR7
DneEZpR7WdJFcJVUDhPH3rKvkqSakm6T+WykKVg0A/YOn3QNB8Q1X1kMH+WVgtOg
rnEfMb9zQ/9uUAEKOwiTX5bdJ00OcmAuaY8xu2/UycZ0g9L7+2Rdt49lDbmfzh3o
ytmj4AhFz4ekD1Ln1rrvkdUTTX+RKP2QOBf71P3qfZIbF2SdngF79Ez9OPwzB1aS
yRf5//pleQneHTdvgkmb9TtfoRC9ySgC8jAGJd9oC/x6xzKZZKkTOd9SSas5K/xf
HLrEUAAPbHX9NJZS10+wZrQQc1dSXGQlKufARICLyZICKybM2cR7xcIp5wE3C98A
6Tz7wrqOP0IG3l3ZUvFBBeNGJVZGOngMg+D7QaNuvXxvaHcaKeVPhanjldRl7FlX
xkc95tziMxgvYmFBHEaQ04wPJ0VfYC9wHnXwWQ6M2XYMStgqOBqKZQyMrmI3PmS7
gP0yLb2yicEGodkby84b84k3NSgl/WIGCipN/HUTCfk=
`protect END_PROTECTED
