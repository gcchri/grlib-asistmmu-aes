`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ItXoCcGPjcSJZ2fpj7Ssqei7ZAi43bJRo9g8jqpJ8wQtyBlxbpkvqyIk57H3T9sP
mhdccdJ0IFVSIbbTYXemonjkgJawm2jldVfLMfmSXx9rJtTbbHew8Ua81+mNOeKa
6upw1JQyoO/QqGlsbTYZdnXWOHcM5VsVhnRzu0Ur0KnAG2lP4NvXoXKL4LkazUUk
Uuu4Mo4J4AT5L+oICCbv9JMKXz5IbL+ODlkgKe/3jcwEcqBXFq5bK/MP8FBwATkR
xFD6RFZOKDTErjidcSMkZw8rFIq6UVHzb8Hd+2cpg6M=
`protect END_PROTECTED
