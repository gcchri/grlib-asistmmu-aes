`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ealzAtuFchw33Jq9XAMyAzeFkD4yhpBG+HxIvaKnRHOUGlKIIxyrNvh8+nTe/PbL
RMLXzqgZqW/G9K4vsecPt+IxEGDrMhuQ+jbbCV6RovyADjChN/8mVSaB2G9Zr0Q5
sIPQzdpuhTHznOF/qDeeszXdy4GBoEK0bcwT/vKeMu/t8FXsT3OG6VDW/l5psVqp
eVOxKi6JJXCk5gIL7uKF6nfJV8wQgBVYhBgtldjoW9n7v0MIb2gVtiTDWKh8X06v
osA+44SuRdLkCKfdlLWiJDzaEH1ekdRRUtf5mg1z2L+yt0OnTwVqb9nO0Kmch7w/
vzEYpbb0QeiPAjkXH1pnt6xWFF9nJBGe6WRlzNPGHpkPkdqmpXZMOLZk1hR94haS
tlaK8tPyf04CDdtTfIKgUb0qelpVw1I9RBowkywY1PGsxVAysw1qzFDrhAuDT/Ao
B1cdjtNvOwW8g87Vjh2OS6X1tSAqna7yASCT3i8RC3xsLxz4B0VemuKKT/g4FF3b
5bSLGGgwVBOsI9EjW12Uk5ghcB8a9p64NhKcjckKnRhyZ3cDLkO7Xg+BNUzpbBEq
OHs6eLk04UJg3MsBfRMoxEkPKJVHM4fuYARcKR88jYk0VscPCJoq9Sz0XLi1ryU0
RXtLcDOe3RFVFBMdud+jLu7Jw5tINtHQyOqj+Ornn00v03ZXljMP+T1Ocmerpyt3
dzshoKwVVvwHHmKGnRNy9bStCTfemcPExwwkodhacNwcny1/3fUCSa1cvU5enPtv
CSWN42XUJrzb0t1u86hn272OYoncRAJ7MnvUhjdyyqF6Je7q2cNt3FBCWbgTaZ1F
uttd9YMbGUKVvjmnNfCOcFn5h3jQRD9ot3xd6qLl3oObvKEIkRO0gMkwIYBdNvD9
bsQBw9WMqSXQqpAtbVa0qEB9vO1yEcRsMDcFWPvxgu4z3IvyDUB3qtb+cV05lCVu
`protect END_PROTECTED
