`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yjs3Ct6sf1aOIU4ndo4y+NdDdLQWNT0+rkhzEOxhkZVT7bfE4YJG7M+QFYR1FC/5
GxQSRmAUkiLsi4pmp5f4OwzsmjElXOP3LPYj9tsZrRRO/I3NSaL3soCVvmiK8/hh
192TFgWqvRRmOs5nm8R+Sy3R6PSj05F5QDvinbDC1xyJ280hTNp30bPnj1oAMKZs
pdvLrY4at5h5AN4bcvXxwrfSKhLfk0q3J11OYoC6b8i6/uVEoGA/EODmtF9151yK
J+TMZFQ5T3/tYStEsz7VY2DoRm2YuLO47sZWpjw971PwMSWSP7A6tk3MMzL5iuVT
UGun+n+e9iZNDqTtZZjmdQjuE7aSMuWFeDOaGk0FtcC9Q647+sdn/Dh4I8UhIYmY
FjRrkQ/orFdHQLPuj0kEFwtVGzLDg76rBnKwZG/WTfIpNEo4YrO6f+f1r7HBPQlF
`protect END_PROTECTED
