`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ln3eJY/+rd0b0DJ2LKiQEO0fOYSw7nggw+HFSiwhx2Fu5+SG4faViKovC+H1Hyfx
aCVON2ceEYYo/LOkyjsHLyfCE3iFeHQjAf62JAR+XBtxd+pymoI/fAwexs8P+FOB
U/lhJE22qu/UEhUiO3jKd0itci/zfrr06hFWJEgVbOPkKMKxOJD+4j6DKDFu+lPL
rHo91yRaj67Lm3nSalcrUYjTd9jDT17uK0Vo15nkfoGrZMOujR5ebFE6qmZhkcFD
fIiWLZXOXwIA4/UATJB0jvyw6ksjreN+cLlHetap0rJ8+QUj6qqJksn1T9v4VkE9
DWjtAmRTAgZ1lIj+VKidXCtw/4URqn7EcLSQ2n2LPC0=
`protect END_PROTECTED
