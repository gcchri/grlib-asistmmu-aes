`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
02M6hivEZTN6ztWIwba6MW9MV2cA5He/44/M2o62ZUnipOUv5/AT5p6vSmVta0zJ
oJXZ8O0xszA5ZsGvOzMW7NN+J599c2vvTlIsQNYwVuQA9GZ1xIn0EneaE9PS8fE3
xUQSuWoJ/8sP/Nkiw/mk+PgHjTtfxOsbx8gaJksJiJHKRV9o5horxAP4HxVhleRY
b9nPE+RuprCHxT8hZYQBxAnnMB+U2liWsMrE7gb/DBKGgeGxi6BvqIP9MrN2Hr0R
Z5fp0rSOa8YuaysgPYEH6wxm58S2vWuX7R+6XpIZnY81YN52Zdajnvwifjd4exUj
G7161CEMTzBke00+qwJuwR1Qmqx0CEkxdkylj3V+4R4fHEhGJIYipp3AyjSHCygY
kG20yBZL78eCOIKXs2vxh8iLMx1wYHeiPN8rh1hH8Cg=
`protect END_PROTECTED
