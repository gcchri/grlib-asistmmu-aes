`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ElJRVUi9bxHcIEr7brCmNfrALkReWcpO+sRC/uSXWAQ3sXGMlCTCpiTyG9y7AEY5
QBaEQpZahNhDuY6Vuu6PSfa9ugt3nMb0+yT767ZaGNVVqOaL9Fao9G2dWyxUauPs
TQ7GCuV0v+vbd6N7okFcRvZsZ+gKvkr+UaqCsSXyaHwGUaAMTh/2wDBsZPFTYNea
D3SaTzESCSyEimIJEYCBdm637sYtvCcm083fXNWx30SWOg83CuJckrZB3E3UgEiC
HZVN6CrmMNlkSRnKxaDdFsSNsi2ZgHMkOw1+sv3l5eavYToy+1UMz8XAwWf73cR5
R2g7emIKaz36Pbw236+OE618kRzyQDMMqbOSOstZL6Q+Zvw5XzTOOx05FT2aFSQw
FZFUFTyiQYGrsTlbrL3/hyCIMmE0s0FoDjdrmfJ8fi3Pn3+XJv8/9xekHmXZNpky
q+EMaoDn7pHWrg/nH8LaaMEKqYN7lLMcMpk8IaOtm3Bu7YMIR5E6779cA2Q2fyz9
6c0p1S1KJJVHtlyBQERc5jO81/siJ1SSckjNECjKbcs32tEvZOGYh9CI8Ly4t5lK
hvLsJHl/5gB6xUHFI+mtodtiSb3i0nc6kQ6vEf0A1Vly9gT3whCCjtI8JLRGGKpR
r+InEuhMvLYZE9h63eWZQtb9A5eiWxfi53cwfZ2iDoukrb8wC0g98vSpTIzA5ZJs
MCrG0ZP/TCOWAnV24M9Vv0DqGU6lzJ6P6ZUbAH8MYDckta0BQXAYR6u5rZvaWM4Q
Pn0lM2Z+2N/Ni52A64uhOws6Y0V612oOU5LfR5moBc7Ks95NLGWg6xEOWx6Y9//v
J9IV+qYVuTBIQfIXdgOt91aNUNBMvizWH15uySVCFrx8Z1LpNKVv38ZfhxbF55Z4
Gfm3xsQaG02zMavkiYhE2nhSpckNEHbJOWSQNVFhdwNqGjsoPPipOWEFsWosU2JK
EfsCkU6h74Rw39trbOkxTUTSUGGFjcjkHRWkcwU/5w8UQTubHN3Zo6jU7QwdQrV6
jBg0nwES3YEJEQc5O9Qjk4g1FeR3cSotv36c7JhIomxbJMwJ0TguMfx40r5guMoK
A2aXfdWO+lo1NIH6fiGhZJvjB1RsDj8KNgWOvSQpTk2JII70mmA/YQCbNbPHZ4x9
5LY6BKPJ3G7kQFYYqjkVQymqc2ZvmGLMmcMwZu4I+OqihANuBKRYwsFs3GfJz+DM
6cr3IF1CGrUHIbVqfyklKU5XYfXi00hc8bjeGU4pLaznjOmqXAvsD9qkp/MJww1v
ZAtaeG6+HNJXMyXBn8Br0yfrvQtjeroOSk9AL1F7phlIbLrrB4F/gCSnDiPcL9me
anqquBuX2Jn9VcpMx58vjUW18Q00fb7GraMhR9CW3MXN1Ev7dTYulNn+67k92lGc
G5GMoG8qQpM5ZTUOjFc2R9UI5V+w2P6lVudfzNEzVW8jNC8l1tU/ZCavOcCXnd5H
IgJ1+1wi0mzjBxy2KrnsF6QbPAvp2ypVdHXGEnn7PSnuL7wQgwl2/XguiuRNj+oj
pKyfbJrCGeJGhYaXZXJQkjSatEtq8PS1yNc9hzDl4XoSMlbG8xJ4/xg2Kp8IikXN
XQ16Gtf0CHAPUWqtbaXmUBlEBCVjW/YUD/m+D1wIP6G5psFc5YzO0XG/hVxp3LO0
VnFrxqdLyl41cxpOOTZLeqgu85J3kX6e9CB5GfIhaZRU3dl1V1MV3vAvp7QqgZvl
Bxka0M7CIMAcMtuY7XEtv5kf/E6Q/FUTKi0Kptya3HzUfMA1IvyopDLtnV5ll6hW
g960FB/y/T+Icxr9nv7tStyeSz1ytD/pvLrEHK+gBmqGA4weBiE8SMPrFn2j1/Op
PQwcu0PCbhvUpavJYtUSlFJHZa9e0XqEvIdBS5hvrvekJZ+PRrSkbj0aXsj0Efiu
zDPnP1FFjtJi4MNrR05kS3YvpFgD0j3PDTeX2TbT9dddpDSW9QbLrIez4EaJ5lA0
+ydX9U1B6VQvQNox0Kp7BAewWmZxbiX7wYGKvtLvPK48jiUEQ8shiJRqKCQs8wMc
QpRZQt3vEwPMe739SUdTAAysm2wpIWBJgkPg2qlMFNKgoHGkTzr35sDaefb9Or89
GM8h3/edwInIYpXHFmXbUipUO57O5vr2OdQl+qAU2bHsFh8iXIBWJa6zQLgknUQ/
ddzJqsemnlHS8DJSwVWKM5AtYURX1qMnGGXicxHSbYXb/VQHMF8mn4oexWlo87H5
LWzoBfsG6RZraWpOfjs5yFGvtIaLPCTCyE+9o3OZ6BHJ1oft4a/cXDV+bJOq5CgP
V6epmvYMURs5fvtDfby+ox6NeJDAOljb7CslC3Lfc2lAWMQkw8QEEKsdnoCqRbOT
YR0o57x6ezv1VnpYkRrh9h0d8YpK5rHSQWsEKlMDPOUcjPK42gDLXxEFHqqjlyEi
OEhlvrWQt8689udA+COJwbmUq7mpOHAKzMXAUDs2Oz7VKP4NpXGehYLI8DSTxF1G
sc8ZHDk2Qi70StJWqr0bbHeVanmi1nSS6Kn50m/1yhAIsz31IabmO3hmqw8+KgCc
bPXZ9RsnT9P3i7f0kGXDJkGYOcxYDFgKpXsOJp+MJaZnWNzR38ztGYVoESuRW7j9
LgCerzm5MAf1CM7RED///t9Uz4WwJ3y8CeYGk3V5sxWN4DwEdznPesEUOLbFesJf
IhuO4SvZ3ksklGuUogCfv+7d9AIfBhWKU3Rz29+wiibISFArdv1bRbapkIXaD98+
4ljfrXYIvReD5qNALTuKqMmZF63F0MrNyHoejm+oQQfn1gKdqrj2Nav1YZ+MMl+V
stryM75VWTKyVtbsJfqMC67Oj3O9P5LDhMDDYdCzO5ODyIxD43rATUdMozXLT6DX
4/0WHQ3alKuwno+PGllSFLP7kanA4gEQfftO5KwbOwlDhBruJiq5HoIELUJBZvgf
rhP3kXP9v5nx7koKzG1j6tLXybMKBv2fCJpaDoHH7GjelpTHlV4vzrsFj1PlIo3Q
TJ71sfVQTiCqZRMy/Etk1KzYWl19tZPD0viu+27SJ0M+hQEGsH4sA3lwH3klyO2T
mWLlLSfU2L071smsTNr2Rfe0A3J6GSwx8Y8uVbZ+hGWydGCqMgZ3MPFckA8MLF3Z
bs3vrzfl5sigRZFV7nF+ZwDKH28F/zmSBRsiMSlTE09s6YzT4MjxF3mlGUKB+thX
1v34KfmXufw3uOm0Z8/JWRwxpW3QrZqzU+/YsW1F3/z9avDUvHYlpQH7qK5juNr6
igCRlPMEvqXtrxkqsCy/O/GDxTuOqYd7vEL04zTJoEuuf7VGg3sV57oyPmdLI7nP
s6WFC9Dfkp5AA0G4nHfvLroBNu1qZCK7vCk+FF07jkf0bKK2RpiOm8RsiaNzC1ja
GQs3PEnKKIv+NS0+dmdbzf2x/rRQEtD2imQ4/399E6Ciwsv5IXxOqhQM5VGNr4yw
6/Brl+Uu2abQfojuDQhVWZbyz+978BWqYJnnhzlY3HZP9tB7OeJp88bmTTbT1RHB
tiOt3/4FkEitze8D/03l12Yy2YIqKhb12uK4GSzLwyd9k9NzdUVpkICL/hs1D1+7
5GwmjJbn5r2Y+n36HQFRRkv0mkh/SNDPlhSXCC52PTsT31Rl/Lms4v4+wiuHz41m
uVbaWXVRieD+0zOdr5sne+zPv8OuodUGa6ngeuOgm7f1BAtvs7cN9uPCvbjIf4wl
ctBfml8jUnJr5/MdeLNNJ24QQ7JjyF6YirYY4nnKbrl0V9xWcX2kdmTC5WLx08K0
lXcWRyWLV6EMIf1qiMjikl1ziI03HZ+rDkSmEKkFX+3ZauaaDcYhLqtwPNvEEJdP
Mn6WVSl2fhmXiXgHAPY3If1YwNrOLvzP37KwS9NiWUj0sHQRmLFvLnd6RJxr7TSG
+oRE91QCBPRyUzCfi2rmU2jrS4efdZs6oubB6NxoZxw8Wss8hAA0v0vL4/o/Uk/X
RcWIgUFG6a/ITyOEYJxDRIcQuEc+idwYylHeyMtRof2etwGzVOBvwD67IGTB/wd8
sfShcEk2DqYv6xqYKOrv3OzfVhd7eoOTyZe8mzX0zR+a4CZxL1+NhluWlL90RCq8
84ouK2ShOsN79T4LORdXWl4V3vjitrt2HZfUC5FRbHTX+gbkZe3G0V3UO84OqpVj
92x+qouSFuF6AtofKmgXfSNAasj/OXiN+2QnrbkA+ttUkXR8+SfwdX89r/WVHgXo
BDQd8cwL5jDjPTbsY/PGWn71wtmR7HA9Bvik1oAU/Pqt52oVXH8633lnqV0HtiDL
I9QJ+P9jFC9R8amKi7FsLJ47Xorior7pnZ69Vlvmuerz8NUjQIRVJDpQ1oU6lZfY
Wj9Il2kzcLBr+UyOyMzuGP+gC40sivLWb3pVJYDY2ZpnZvJXB850OnOGl9Z0apBr
KNhQE61210W08ZsgvTWyy4hIl5svnZMY/Wn8D7jR95I=
`protect END_PROTECTED
