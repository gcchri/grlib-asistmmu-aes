`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfWcudHXF0tL9rcNZPtiAD3OiEWVPFyWwFHRPLXHPyUyVFHiDHao4NRwVSHRRH47
+PGpWiv2qazdD41UwPGAboWQ37MRGkTVnukLhY3O8/pvmj6Bt1cfVdSgvC1mv7Mn
HiZUbZ2N7UDQZUUnjOhapZLeRYsOoCNe1lxpKJlRj3p5qW4u6moviArmzGoqDgsg
SiAXGNOfJDJcrRPv8hVAUrAwGfCDKSTAOyDE/gF6Fy/IbbpkplW0Aan9iK+fCD4X
tieW9s7N7L6bYgEc7JwxKZXF0QcHZoTy65wX6frF+H+fpXPXCWgwNCrEr/mG1eC5
moHkk5TuJ5WtQEtag9Af6Av/CLEZdLNEYRrnXVLqODWZQytjHPFXCeVonJOYuHtK
o41dpsWVu4DTBLxYWPpVGA==
`protect END_PROTECTED
