`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixYrxgsp+Jo3ntMny5nVT9DynKHztnd0TwUCbFoRp51fqf72yFhurNla/EMV4njg
kPcVjmG9ZeATK8c9MvVNTZTTnolXTErf7ramOXQDNs7GosGxYZNxL1B5f9R9rELb
CCoGLY1b4xrlPlugORIB1MlNffaSg6v/DUTyjggz44DtAZPjSPVQ0YyIAYyM+Dxc
klYLloXAdGMHb9gH7mS3GaW3GMDcck2haO1YDUOzTaLPhnFphLw2wLDF8bpKVL5Q
`protect END_PROTECTED
