`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ib6aiaQG6kdk1IeDewCjcwNoy40Js3SxSvSnWGPVO0u6/+bKlcb7uMX5tcx8xxu
Q5HUqzqHjUw8ITUtYnje0/QD5xV2X/ZBAszB8l4RiLqj/NDGflWSdTmcheJsKyv0
nk9BmOCfU/YLEwoO7tby8bJZ9vDi0QQ1HHOcV6UhMAFZWvykFTXqXT1AYL/QmpxF
AIYrk6DITPCIw0bMbGtUAhN9SD6Vz6mJGtFQMLy+zVQJt3B7Chwq7+MQVWzDlNNb
rkmGVudMH1Grdx4CQrorDMJbGe7g7qaDrafAUq9xdXo0LXXL8IaciinO4HmgVGwe
rYfnqpUoAsACiwU9tqs0AiDt64ar29YSoImaLP6jTsIhzyYRBAebP1eRtXJr7K24
ZVsVII65fxDnorTYcP/H7CAnrAoRVDytO5CjIHrQM7MDUp+ToLZ90mQ/xglGi8t4
AoyEuCfI79WN4wKGEKVmGWdjqm+tpzv/UM8suVSJyNU=
`protect END_PROTECTED
