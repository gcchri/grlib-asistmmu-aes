`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NSOgntO8JGEEoXPSJpICxja3R7BxREL2yj8cA3q03RsvrkTBIV0d42CoRtj6kvrp
tYxaoPd/YUyeaw+zsdVnkNZOlkly/EyqQCjc1YVS01mIDyXcldHvCnUEdnOr6Ma3
B1M+IR+aaWHv+Sg0aml18pVogaNw6J+1kGFFGt5st2bYPNovfyONby3h9RX+UdD9
7SQ6lLnUyOqpIt/QWSelLhGJgj4/TPYUgu36vL5Do0/f8vZKXRyIWel4KUzSwish
/7x9xyMahOCZf2/hBSBrHHuKVmfFoO3eio3RmsPWGeUluFnDuoW6pmrNMrqtGGGR
4DjGYSZSrNwWpKnrL0bCP3nTYn4oYO5mL9oawSX7jvCJ8X5emZIhKc72L/AnUGUJ
IeG6AUM0p/rdbYCUxNMqFEVyKQuePbj+TnBt4bbAiQe6XfQonR/c+PpSyBRZK1jO
Wfl+iRgCzT7+rckh+YQvoNlDODrJPi0aH2nrfU86J66BY169IxULGVn7H4jEANFw
tMQI3VRAfzHwSlf4d58p/HfUX8XKAsLOzNXT21s+IHxB6wh1y4btngpIVaVo+0bG
ZTz5JOmseZGKsZyvAVlcTF062Ao8xG3qP5Yv4DFctP66wfOKZ5TCM0Pf50bkfBjO
CDS3QoxQdaYOxOcDI6BGMQqKubcjJIvmFxMi9E2MZabdH1KNOqddaCJ/ofwRssbb
Q4AvKzmlQ6qWrjQtFJKDrvBvSOld8DPd6hq5hmwfx4UcJLOGiT+pjNGzcVtHzrp9
GG41so3CsAJ+5fz7k14DDRIRkE4GU4iXk3I8utjdvzQkMH//zH0ME030HmS6/EAU
WprRuMYJrDf1F/WyoXrFt0orKB2LKbAR4ItRUgmYkgWAituByMEuFIWsZQUDUSFe
88vdZXPl9kvIFm+l0DIKBATfjJRuNzmmDUEmwXLqgtB37Fqgy6jKngWhZ64VGkR/
dcDRHVOm3C6FtA+r2yf1Dg5QiroJtnDG4UfO5+sI6aYN/EcmDneITx1/qLjZ1Hgl
925gEbE0q/zj5xrj5pC8CrkDfEzTYyVA/ov/4GdN1OchOouvm4hb5OFUGy52Fz9Q
qi8CAhtlmR/tDklKIMYv+LhAxZsiu4Winq1qj/gIDj8SdhtLk9kgWdr04Dq85NvQ
8kc/P+6mD2hJbpuloa44mqOk1suqrUcGOM5upovOU85Eel1wH8HEd/9QQO8x0/0C
MUsIM785v7ASHPmvoF4xQcNmq3P73/AA71kW/dMd8Xk6FR1iswxSHkQWEv4O0i0h
CmzPaldU7LR9CQMeZoPg/VPLrA0gYnfgbv8DaHaV1gx/1ys9thel/Z6LLcuao7OL
pe7pMvzNG7ifMY3kzdLX6PLiDXcHYTrWmAtda+cElk4Gri3Ii4Kwl6ThkVfAEU68
qGmrWDTxKM9o0noiP8HdTAleIbeVRUyHGygaIv2iDBJxUW1uQw5gs62ysfR3r1ws
XO4asUNKzT7SGxz6pgQUPkzO8fKlyQ886z7K+KhGQtszPlI/hvwnY17DqG96+KqV
mRYKhmqZe23fj6YqTn1OcOfxbs+tvwK6U83jBtDONnsyMPe2oyXvy+9ejKIPvluc
hOc2rxK1x46ti6xQEnknQ1IgmWoGlxwP41xY2F6ox2j1RBVV7tsjO67pQI5Cu8W6
KI14AMcZDGUehn/ra6W7AIv68PVVqTWIHEC/AB/S2qpgzN2I2BK4padNSwQZFpIy
xRB2bMadApsN7G9e0zqsgqY3WD0qBWJ7OL3xFZPgEuR6FFr4tnJj48kSegp+hxXl
+/P62idgJXaeVznZKqvT8t7pjBTdU5JO2tOGUnRCqfThLtR8t2anh7e/8EEGJQYi
lXE57fThbvz4zbptuDaDeKpoFeFV4K1M80o0UOOX+ThKJBCd7QvjXKvWrvMfftx7
H54IZPbJ2FSgY6iRqOtiXFkXQ7LOaRzDxDGkRF52dB/P0K2O/Goig6JJubT0WYhd
VjfXPwF7U8u/zySRmp1GVR6H2mrkFgAmZBRpxXyiS7CLV9YW/hEpru/jRa1fgKhu
N8sSJntwiinUpBi8WlTp7FuZaoIyJrWgETMmdhUWi44=
`protect END_PROTECTED
