`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UF1FBOC4KJyL13mcEnmm53JncnOBBKPSOK6UiyBk/GgVBNO8oCXV1SXiwLh+y6IT
lsha4XSv5aEvKAVhIhATU7SK5sQ69AIXf8dfPhs1juTOrsJdM0P1ejXEbA/y1lVV
Y/DsYcERl5NYCAf/1j8yv5Yo0s83oFKLBlqPvfj72e3MS2Bo+IOVdAJkwkQ2PK8o
d49SCualhE+yBLgnRJdKUFOMYvsnWDpzzom8M5DdS/uu0oR+IdCgrfJBL18zS1qX
2mb2YVGzv20a5b1ppEtqCIQc1fZ3r0ZQATHw0+hcYmJKCBB6VgRsXEkqid1tY4fP
E1jHN9CuBBagZXE/tebV0H3VlC3QcOnS2N16rD9lvMtMBkUZfv1/7V74Yth6Ve1O
ttbcm17pBplEFEgtZLUISG127ibaSPEe2wJHvvj5ob0=
`protect END_PROTECTED
