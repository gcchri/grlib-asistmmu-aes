`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gp07vwXH141UZoJN6SueVvUXbQ2Tfwkl8plEKnxkNOaGnOH7FQKphuFy6V+6K1iE
NksiUjeur25qsvnDigy6JMb064jYzT3/xp37W/zUEC83l3cDtsVXrpPfRvNRh+/H
/gQ6x93Vh27+8nmeUJoywnPA+Zj7b629zsnNs1qWfknQeP4/u97C2oCJ+0rzt7Nt
GcetImJFKmAWdJ/7x1WA3j0irsWx/HAflgAsNF7qXo4RRu88dgcRRS0lR+YtF3P1
0iw98fLXGfd8ZB8Q6MdkY3TIGDf4CDUpi1XKDU7LVtU=
`protect END_PROTECTED
