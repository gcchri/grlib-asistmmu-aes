`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zKsQV8Cp6uM52sWfIQdlyXWIlRiMoEt3Y1iIDisaY4ilMPJMsa62a3S7Hkf9LLWN
MU0HgzEMIVjyd8hwFm99tNs8/77bO934GSJ8mAh8g7G95J7NTQP6m9qhssOhlrca
4TTHLmgCf5GnrNXsr0NNkJIrx+aHmzsKPF/NrQ99tdray8fUdjusavx7gHYjm38P
AQjzFBX8wLnHAFXJ0S3rrH7gEcLEI964K174V/Xg/BJi5BOaZ1BmK6WDMgwos4N3
fyef17vvnlijZaj3xFK/qCkyE9pnxGexa+r2XNB8YDqWRZaZpZQwbGY2DlKwzXh6
TzPF1Krhs9XGjTn4JTABH9PyIjFpBnyxt/1APyNYz01QXiIxL/4GKbPdN63oSLh9
QmmfhFcu6IgAS6jsA5vBi4M/FzCQIeqelFvxr3L5HXqTnzEuu7uYqvUE4eyB9JYV
s8A211968/m3GNrlq1gPmQ==
`protect END_PROTECTED
