`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nppGKOOoFnucj2hS2VWUVAQokLNcCbDppAunM9c+LllEL4tDU02z8KV3HMd4VXL
jZh2QgsMA4HitTihdz3d4COJNlMVAaVGR9dtGRc+h66C2cdDvNRwwYr0Pmn35BL0
AkIk1VarAvF4ULBAj0bZPa8whr4bKH5fLNegljCQKIbnjpxOoPZlSzMJ874Q870d
VQMFT2EU4FXh7jLpj02/etjJkSZLVcNsnEK7/xctS37DB4yjiYH2bDuVMPEKy/Md
TrHc2qNl1bSWSn085wi3U+NIiHjBmpf8+5mDFxnHDMuLmjqQeJE+y/qJyXx0J7r+
udCaigMAHuuS5EvW3QZC4aJzdBevUZEhek87asxI2KWpTxwUzsi8eIV4pArmAG/C
OABSEEzbgEKzASn1OFOuzw==
`protect END_PROTECTED
