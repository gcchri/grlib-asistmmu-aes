`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iN5wlOrPxXymFOdF/MzPJ1E2GlsumgDt7w6PQk26oSIFcd19TtYt4EZ7qJYYj7k6
eD48ponXPkKL7wJq4tK8+b69gP3jPLFDnA7XYZcX2578sqx2LcEjc1hvmHqPkot8
NQVEk+eYoHoOgeQWbs6gdkSJKvzX+ryv5kyYj6ncWvea7En1hiyc2H56PbW4WsP9
JUX1ktNzLXl03/MOjQmws8gq/c0SjNtXNNQjNPWhTa5WyiJx8hf+y9g81xXTPbL5
BjUt8N8msLs/t3PQOBwZD0MfXojM8VQOzT4nsYxvW55eJ3zbJER6bqvlZ63wsBZr
JMHrwg7s/k/Afzz1+suDcDImSREgttOvbFO10KMV99y9eD/hcy8wFGKeKFwpMxDc
4tbDnupyF9rHRFU+vT8wqlCDHtjLgSbJuPjs5AKsfNbGer08Fwm3CqwqtwBq05iG
2X8sEF3BNAnoSqqFdhhEOquoupckFEwOpNuMjNc23rXqDbUsVUVWwme1WJpa39nW
hPDO6cZ17o6lvaXCOFWz2Q==
`protect END_PROTECTED
