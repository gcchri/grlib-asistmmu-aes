`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bBCWzcWYldHzpfsLzCtCFbDigY4Ano6N7SqYZxGiS9q11zlHeyN79S60aYPmxkzj
ch/zzuRlJoS7yCXFvgMdaCWotfDgav0nz0XzA9mBbGizKu1rmdDPO4lOpNE9yiag
Sq5ks5UhG1WSRIwCsLnx5T9SgAoiZqwXmuHqW+UKFjFg77M67d9OKREr2OE75YhW
1V83R7f4Lx06YL3DcRoQuMQu7QrTuvT7sK0naYWSSDKfFD2CW024xTAz12d7Qfme
ktYwo8z2uBN0igUUsah0d/W4iBAro6LELY65s7KoJrwBaUEyOSpQVnjg5YJMMbtu
Lx5qeRW4eP+FAhzS6XevzZxr6Af5RKumgZ7qZVCQAOIQtSuXBawTEqZ4Cy6/VCbn
1hSax54zu5Rgs36ZmHjOj4iPYgIOaZjEk8s8gjnypko0+QU+L6EfdKZlqDmBKElC
dQ1jTIeDVzLW/yv30GTiZlQtOWtFqs7rSZvjScJ7T/Z+Ty2yN5xfernJxsK/eCcg
ZsWR3bWTsxEW3jL3lzxvKxIthT3NqoqISoNo7wUrck637inKcgk11aJP1WBngg2i
+CfANAJj0Zql+y+VKZiX5lxVmpBGPzVn1XxVasrpnOK8oKrnJG3RN7XQSCTANRbA
0htNUVqtLPFPHX8k3rXleF86jxi/EQgYmuhSVeUhhCQcPrfl+s5jkTLjd0atZSOP
DShSi+wIsUGMfsMuL1nO4WXnIK0AYCp4OZFPIqrwfTy28BPHjGRfMROp8xds3i+n
VRcGMR76UvHrfiXZ//oyc0SA2glxos0e7MCCY9nj2DX/dk9zXDodgNyH1uLv2n0T
a6+KRWo3DVM+TMyHQFxsZSX6sBLArEygQnHnKEXk6QO21MjYSqQriObPIXqpbhBf
xepJ2SsPZOCeN7Z7eWSzSc8jRC74GcUWkdpzFlpNh5K9ZAWQb/RmIu/Y9pYTwoP/
bHM2G2zzt7yaKNvi8nW5tPHmNJUdPUIPKBzm8m35955jOgKRFSA533G5uscu9KfB
GhJB0Hj8u0GtIpR7RZalMpCRvNIWh2RLKhgJuJwLjqKERocOPMobhijIgwtpLkKO
8wsiM5rR7eH2K4zTJ6h/7a3SEb/Vx/wLPN4ZsKHyBzgH1aQLjar6XFzCJKfePB7I
kAQrKyiRwRqKyFSThLy0MdNO34lhHVO31Xt1+LWqiKyTZPdK1rF0Kgk4B5Xg1quA
qe8PjQ0UDR6oJZXR9cV6tmXY+OBAwbs+fgjIGE+eNiGpNhxzK6F/3shAfBY4IyOW
NH86qGfBy8nDVA4n4ezGh+g3AGafDHxUY4dLzwgx1prznfpzUKlyRsZtpdPX0QI+
UaFrsFygCVO/0trO23Hgx87ETTPPGtP9vIf07xe9i4ZQp/82fMXQft8pGZf3HNcV
vVDMFr4eQ9cGsoC8fqjH0kp/E5acmR9aJtROOxZrU42bfSX1mhQ004O5gZk8on1r
U9dydB3zjbbA74sDyZMT1uXlcu6AnBqI+sq23nsLi7KDR9iXCpeTu/sOTE67vHHB
va0BFNVMH/uowcF22PP5gYd+fJKhRAquFuKSN1O+5y0LgMWATewX/ADCydg0xb9W
1lTkIfvkFi1912mdZFChNryjtuITXy3R9LMR5WCj2XQoL9Yio422CV6E4x33X06F
+xu9FzW9oLrvbO5gSo2oUFkw7a2AEk+kI3K+guJB37Xa110zSiVAqgEDLOwQV95+
dQXnEhJ5muoA6/hLaOPFgdqlhjKFoBAbdKsghD3cegS9jMaqmgiX1ql+gUFK0suq
7SLMr6hDyaEyx8s3aU5J7HsQCVulVZ5PeumYmH2T3P5Cw9Vc1gkvxaatiNQCyqTX
JkGnLUG7B718W4OXZT42P+0A2mWf50sP+sg3hB5WR+RTrbc5jdtZzxDQcToJ79DT
WgL7HdPOwrY+bDEjqSAL9oOncGWmltHROex39864mWAVfNhV83BuW3K01NNXBc4L
a8OGk+aojO42aLFAAEWFU6DSKE76+Otm/Z4cYNLZGmLVrROhSoeT8Q89hNx655Ti
o0ETSPq/+ecxuBPXM1xol9tNbVrIOixrQD7CkH4we2o3LJL1N82lfOhQuaB2gYtd
zz5mlhar4SCyNrq/ojzi6qOUizoopRnB5yvjE9MhISlCVzDFbF4sf8p4M+409lcj
e1uI9KW1CyXofu/3Pw3noIYZrDGMKuTzkxpHtUbyCIRtHgZxedReBPBW5yUGewlB
fBUapvWWkMaAwdY2GrZsORveaI0f30FnYvvWcG/T4JlQGyJxr9XdiKZ7BJfWH3Ja
NowYSlTkM300KoxkbmPctEyyhvXwdmk30uxJwfETG6g8qEv4kOmaE314qQVaD30Z
PpAUHxsgdsXNW1QVUjG92pgCxP9D8DIOPqJu+IZIFoRLmHrBWmdFs1mnxXrt3T71
cdZabFp8WJ7IF5MDSGkoYn+41pL4r7KadUrSyM7NvtZsyBl3aV6iZLB7Ejgj7eb3
uXZ82ktyoZMRskEzld8vlgh9e/FSBwZWqvOKwSjixARYPRBJzR/auvhXl0wM1bwo
jx/0MAJr1aMpMkz6hxaqZcVvhAEVq3JXf0LRkRE7ZNGYAIfvq07g/k0Tbe5Xl8ls
UxayxNKqh3v9i6YFzH87Oal2mk58FTMvrGg8ELLgY7VT9kgZp9irw88jgdTfnWU+
CZgL/qTRbRVg2RyfKhM252upLqApGZL70uAiUHjso4moifgMbjjr/e0FnkIQNIr/
3NHQjPnjmRxV6D58ACGxSm6LLSBY9D6yuVAcn7p9gBkUhYfvFqAM9FRhEYtOUxro
mVxcwHGHhn3RH8DQS6hrk9fxfTWoUgaxMD1wB2VitBLsWG3OF0J9ME/YURbv0tdJ
W7q+WxA0SpNNwf/tUg3gJaudeQU1Y79dn/axB1R7Z1Wiwikkrgj+EOGHpIdus9c2
RONEuoaSThKSstjg6PXiMdYSEfYiiyRhmPQFmVgAnUAoEPoyTt4r1gVaYrdiEb6G
SHWoVu+veHQQlCdj7CT7JlQK+plCBNEuDqa5nnrU/nbn9spkaDS/l9yk86Ozw1jK
c/Z28XLhHhqWX1HyeU23KwYthANV4ObGsawggicJm2/Ufcs5VZlekKL62efGKB6l
OYS621E0ovsESVHg/xtuw1q6VrfC9hMxa0vpN2RjIKcc66lwlmx5Ll5Uy/diUdBS
wvLwPqo8t8+bod3QOzvXyhcZrx4cjISMER3LIcTuWF/qIJZkYdeDyTmdlVfuaEw9
8yJQrv1kBxf8Fx9tMaOsst0K9e2heXISKoT9m9djrFd6zpMWGB0JtMaq8MjKHJnt
YeS1wG8Lh232ld7lMWj5OQ89tr9Kp5EKbGDPy0AvHGNhAWmTeGuKN2gWeRNp/06V
ZDBikOFF44rlRYg/D4kO3ky64dtcfF3wsOZdAGeEfchm+6TNIeAGZ/1Cs0N07xJF
32WE7harrsdq83JLT17VwZLWY3ZhCJHkks5uU1i5biQOVugSf9nFbcvFaQJuOSmS
HxbpLiYMgtI+Bsm5fB14tX4DaLhe9AkI3hDJDCr/liPBr+xjFUHNqW4Ug8l+XqfF
8CDf/xu6bo7t8WIlVSGKgmu9eA+s1Sqf7kQs3Q3RdzOODX811G/N7loNjAc/y4Tt
CPU0yeyqnpZfFQWUdOOW2lZ6TsemYFI30FJveqMHcuRHSV7B1xwDZKurQp3WZ1c8
DTmRMb5VQxF3oSodIB8GvMulWbEmnnBxrT84xA1nkwFtxSZ0rRIbF6z+FGkJZiNH
vGtKEaihaP4exRG/kZ4MO6vJxLW65Yv/Cnf4EXtYdcd1pejxIClz2fvkxxq+lLfS
IE4VEmoH2hHauwfahMuyJg5CB8Hr0ljYjRaZz0WN63T3PGCWwIIeC7SZmyBLG/Va
DAgjVuiu/KGlfh5IeLJBvgVtALQl8BgEG14r5QqLLE4DEsOscSwr4au+1FahAjxo
7lVGDzgtEcm058wIzlMCAVZZzYU/MGZHwKvsHC6OQq+WCVha+6L+/XoD9avofzLL
WlMTgDEvCHD56qIQ2GBsVi93UteVszZSXdeVUQ4csuJPVpY7pjLQLB1px8K8ACkl
XFmd5m5fEQF6S50TKu67e+v+JPo+Ud0MchlgHUWFjHppNRsPm4C3Zdy0IKaxmn0N
x5I1X3YBcvUYaXP2KZE+wA2CUVSNI2o0zEPL2DlWGmOD8gUBsWn5JF6v6+bV3D97
kli9uPsLqlhNSAd7gEJY6xFSh9FcKiq5OyrY45i0mnauoMN/7WJ4xDYmgPgZg91A
Vb2Y0mje/7BA8fhO3d9gDQm5A/5t7JEeGZfz0dwVVaKitY+cvQCGhCDP+7w1PtcJ
Ic/NzBR2eAMMjW7wxN6tKdfTOxJeCNdedmTFlufy61MmhcCv+wJ/RLMopQXihgCf
thueKqAjpbQJjSue4t3sb+u091Pj/s093hi0SX9mbCTWh+bM9bf5gBRCV/PCWIBX
P1wmOgPUI9uuD4veWhzyuy53znQ513BEgwt8c5K7u9SiIKVghx8n1CNyou0xGqWC
cmc11e/rsidP0yBpthXDtFtJKTW8Ct4P7xFUjU3/KCMCl7PhNsLo40VPXyHnjoi7
+9XHdE7q09M9bRS+GBI5OMLepqkopqXRdNpI/Vai7DGieyjo6KaUO+3aD9XTG9zu
ZZIRmuiqwLvZ7CLPpBxz+zwt6xolwTqQsTwGQKkyWoDfqlbxoIrsbjOIlO2kCsKd
8nm6napxb3btupMgwjGXsMxlbV8uhMyx3ZWRzCEselgq+MvxsWdkJFAV157meZRM
jd77YYBJ2mHD1v46PW060S/wRY8ftYZFX30eX8G00vhj9mhWfWKzwEy/EK02uaN3
ERz0gZmp9QhO5PR3EO448IMVYuhEuvsNUltjjSwS+p94mqYp7FLYcmXOsnmgQ9vA
ays29U8vAzpg57BrtrHoMgQlHuDLZlDHjSejdcBTMDfyJdFfyk0dQBCVScv/jBhy
PT7SLp1WIpIfeDfPk8frGhF7puLvmUrsC54KnihBPzSmCkwNiEsyEUyEouUdd4zC
u3NWQTGQiEy29WqwPMfEyNBXxZsc1fDMnhQQr54KGJ0ypacvhsl9RReXIU/XHZ5/
0HdQCnwIDs0LHsSOC+VpKsXk5De5vCd9BOwwyDHZL3XGyD53j9x/nVJ4nHCSK/Ji
4W0FyD7QY4lN993Icu0zKXtlRUyILB8esSeEgzGo/t5oMn0EIbqnypeiLOHkmgZQ
uD5vk87CAF1sZE7stPWusaa9mFmAXz6V6NtvYTFnVz2xXaeg2gj+U8k4n3PHZkaN
dsm1ggpvKHLB+9Ki4dexXjXIUHFsDtt+GhcnsNoo0xp6fMoM2KM0BBghujG0gncP
bLjnNvgrsR4HS768agvUfcTd2vcTjgPxdunNfg4LR2cLd97AqReLiPFsvaX1KwB8
fij0YsAUGA3MRqLsE1m302GpBiCqbsQYwJ4M41OVSrudaNh1osiprsVdVQGsnuHl
9Otb/XVl7pkrKmmlZzBnPgpIxcraHhR1Ay6J8lqY9OoWkC00IMMrlf7pJo0lQY09
klebU9ToSswQmAUdX+y50tZSew9r8eRk91VseV6q5OhUzsVQR4avsO72/Ha04G4I
rFahjogOJ1EGdwn2zVVfpyqXVW7zUA7wJFACxft8uEiiesL0RN1yhchm7iATq4DN
/Azc1Yp/RrfaDoY0lD1q16QSbKHv5KYtTFbiMacUoepS2nZsO4yDF0tJOzOun5Zh
mODa+di9YpukML6ZaXTkc7iDN+MjgdH79U5vr33k8PBYdSG2V99N5qCjxqKYcPaA
jZJxMdfyghB/YDiZMrGZzGkj2/Tigk1jvNDxauB9Us7cqBI2UsnomAO5vknj7NtR
FLYtnYec76DT9t93IFXzsWoAXxXFmUeiiOcz9eDEydtWeQCfQgjVVoAAcX8yMOGo
TtZAYpZfbzksECamdgZpSLym8T7AtIqRhjZAi3FhxFW4fts2iOEb5cXGOCPWHuQI
kSFoz/B0Zie621MgvGSV6bfQdg4s3p9Kp5n8KiqXV9fQWDVdUab3OIaAiYk2bGQh
knJBQ93MowNIt116aErCjYeHNLrrS2TnpEaZEB4Ib+CVB6pVgJfTuAZbppxGZDXi
8q1UmdhdaOFfHuj8cJSGsFyKgEI+zdHl0hQD81EIVC3o9jQdKVIcbWtRDBDVQ82q
G/hNyA1tuBuuWDYr9BK1gfsElKoZoctILx2bdZXGjXZoaMx0UAQ+fS4WYgqegx2e
qbxCWm/Aiaz+YyGUx0PQkzB8BvH8M3zpgd64RzBrIcRQJe3JJGjcMBSq85N2gV9s
6OAN1W++WUHSbwtuUzWjItS0sVjl0SM5dFUdTW4iXhc67uD1P+sCItrbLKadAj5S
R6np3lMfNfSOHcueZX20X+4CndkyIAqsypL5Kf8JwGblE7gLii8IjlWGIwm8KaWr
taSH274V4ghp8omfE1ISRxE5nF4Psx863QqPQ3BZvXNj9S7bwuEMnqgmg9eh4eu9
wqBr3s65PVwHsayBhPiiQrXR0tQshgfwexbfpnEGfqSB7bfKC/iTeJJ1H7ueLx0u
mPmeMCsWtW7gmPw/d43SdVpVRc1srxI2c6IwfRoEgwNfBHwJAKEh7p5A1WbsQuzz
OysCGWjRKwntvVw6c2YcR6Kb6RKpiU59b66iZ+OJt1QjYJ80+F0PtPZaKP31uHuK
QZ3dD4b7oHJ8xsvYJcCqs9K0cAs4RpLgip4wI5+oiltbrScpn5bninbKK3XGw7jp
sb1tWNTuHAEwevkeK0uRKp9rQ0ajPR/mzrNxnbkXpQdHzNfYf69lsvJCeJaLZwwy
qROYW2DmWZ0bKxiXeUo4hCcSkFgGMhUhQKUte5VLrnkUR4oRkwCIu1wHyUjsVRQL
VCfpzvDlfZiPhguWYmPyv24kbzSg5cNCWuRaqrPK0Mugr4jLzHdwprC3F9ZHk7DC
VqUQ2FgnbyXYPrzmhsrciypncqCwwvU2djtjzIunZ2Wya/mYiL8aZdMmGl4ToW5g
k3L/5UCJuuDBNuJg2rb1jUNg/F2fxbPP4o71G43YXAJuHTe/AiQBojyY75JaBBAZ
FoyaO8IYure0EZj3MwFm41V0BKXtkIWzC/0KmqdZ61yJGWxvI0t+4ru5A+lvF+Am
4/nnMfSRjrTdNmR7jxLyScyH6Lxbd9L0CDtGds+viVd+jJMTDnjzrDyEps2V3ptk
IXwsl0lp+L4A0Sfooq3X/M+GMIm8jUV6qXP54JNKp67JFaEclidGZUjBUaaRto/r
AKnAUgQKWS3dfIVnFSa2Bc4xaGfEvbXZ+z9aWPIbDknrg5uFE5apsiBhTHmN8vx6
bSokVFm64YUxYafgZ/lsw/E3I++LVso6HQvCSYRRwccoQK4Sy2d451/ZDDo+YobC
y7wWXeMCyEqLWTDA/tsHMqnySy0KPPailXktjutTUDdw/8hqihUrZooOeNNh8EIV
v/4Fm4VmNWs3fzVu7sjvSwaBQSlSLOl7EjTsy5YNsEoel8LUp7ZSTGMctZlxKOpE
W7VAB1bf2z1vewEcxa69dCJcCnaM1cTSrr+blw/ay2KsVlB/+FgodEfripTo0fH0
wD3s6SyasIWVcEUUDsbQCIagNNIYfuPY+CIES9BRz5AssmMK0x91Sy+r0s+lzed7
BmC9kIYjw2mlkxtYF031Jb/FMSP8mKNJprMr0RCYM/a4tyQaOjN7BgpcmAhMSAfc
CxVUoUAVGYDzxBDFlgoBR4PQu/EFbhRUKO2I8mY2mfsjWJnHz5rwKRh5bmAU8bXn
Pb3yDjD22RB6ArutO9tU0ehsGXFITx6akLTkxFk9LAQ6rPquT/feGrTI+oa0VefJ
BXuyt6/lg3Nv6LOINSh18EZd3Uj2zosu3oR7T7Dz1LAEn2VfP1OzugldFD88koiB
dgXbn/ZdmoVVfYb56LuLPI6gN/MyO4JvBVFIhNLZ86aPYZIn9uR0AkOjDvBL8hlw
WpbaFaZcSngIw3YL/lmKaIjLR9GLkjn+pdrz/Ezr5G507qgig1oVFfXH/orB8cgx
kvkzm5s153Lk0Z/X+t91FnAix41pOcDkRpKjy6wvR2VztKdWN9x2GTGpdqc4ZxHw
pmvp45RW56uIAHZtxppORSyGF+m4DR+PGuPDndeE2fm2gJHufbzyD6UNxl6sBrot
Xx0hTnLy8C3f89EhdnJ+jj1qZQlUZS/ZBEWbfwGTpt9pYwIsGHVnrX66BFmQ/wyP
MkzAF7tjhIIs+CSzEh3F2/Vjqt531Cpn2UJ+8Ew1g4mQyK4F5dbEBVPfqvMXJswM
Qb32UUhCWJdCYS5dw2IYG+Z8Yd6HWHyL6Vw/gxqcQorcdJFkptHmI6yEUwpSwguh
pFfGCL8NEbHnfFQfFcl2fr2xoCTYOfRmzvoXFz5d2ErcDEF9HsgaM2l2Yx8Hh6in
/fLSkoJU0euD5meXyLriwpsiGyme19QmeKb+iU7FdT8ycxYsqhJhHLtab+KM1OcV
U5DIieOhpqh/tdScihDhqlqPIz0qBlK9+iOsLiAMyCC38XVmqaKcyPEaUuyejdDH
Ga4FsscNCB9K1SgrOoZwGBjgANyGVzIqxMXS/WLTuOhE8344fbyvZxUl/BVaHqrE
qXF8UQqsmP78sPw6vkp9k1PV7HCDSlZ1nOIPn7jVNhgxEZQlgZzx2cFRt7i4QPdY
0hUijHaWifHcYqBqh8Mqt0xMi+Ox+3cnQXjQaRsaGuZP0ap+hYlKaf9z1Fo/HpTn
XoRzqjZWghKSA3JCHTrkLp8fD2ZgEYMB9LJE/OmH9MDQQ0DaYHKVH4Ms0l9geXn6
wbRigGhj1IFciY4YIgZz3jEaflqgqEw/LJl4o5TZ3/1wngwCsdIULVnF4DgIf/X1
WImdtNFMkLgqK24eqILD0WgjIkaAuhpf8sFnqPSeAQTbGaxXVOZiIeYxKdXYO/4b
J/GXPIapbXIablHib2KOds+jE2ZZ1S2ZbVJHgEzmbaMk3SO/2YZ+GETDmwN8WmQh
pFeY6GSv7aQeGu8RFOtG5GFqPYbv9ZoHSgFwXuY7h4M1BQFbNUu6pvsaV2YTXUzm
0QyO3pSWN8mUM8Qg2JsBvuN7Wuo8erQ8GOwjNRtV3T/BPK4Ozojlrp/rzrDACyBd
xrJehHt62RkT6Imveqy19hBSBCnHGZ092GOjbSID3GcpfxvYlYtqEbFZEnGiYRRx
FzbeJ4vzTbVkv1tkXNDxGww98j4Bj78y2CbGUACkX+RpL9iivJxR8l+AK0zSFJsa
ekVNq5KAq6SmGwE7zBHyuixN+TnRtLiyulTJureOc2ifCTDrM6t+wfu5T/eSuaT3
WQhfl/mYgK+MZ9rtMUBeXVvP1+KF8BVPFGCw704EZMsnM5WNih6TIbU0FSfYniVK
fKsQT1gdyyxfyUlH3M5cPGjWy/M4Ci8i4WRffpYj1EIF8NcIwFvRNLh5Hrr4UMNu
n/mWIMvRTrmrfQz6/VG9uK90oCeijpoydgDZ7vdh+r1SHS2l+A5WkVuiLSkyfBaV
+oGn8mr/2Izs2RqOpouBXG1h6nMDs3x6DgoZERJhT4YTCPObMr4zvUlL7bSMV6K/
3OTKRcSEpmllAPsUgHq1HdQhx1g+gaok0Wur3yEhuUlTjOmBDVjkj7enwsFFDWTf
h8LjmymiMt6xiM+Pq8rtF0pvtu7TvrkRnne3Y5zbWmRyBR63YGq/QhUpxOHH+Z21
V3qOIqq6NMB//bODFumYFC2W6XBBJNOF/cYSzdTTCyzr8w00tr0oLwLrPdUszQSk
QQV+5aH+N18jd6XCdi6NBvVepIlb7JSsfVM7GkWo6yNwaFoC9VUKk5SSqHFT0hIh
EYIcLrCkeMy2Na/crEqQ1yYZ0Y5MwHPp3S4vgnvhpR2MYf7mlSHgt+2sFfvpAKeF
O3VWrHMbIEPi/+Fj3b3k9OvO1OiXpQSGN3R0ACLdis8PBqLtgaP2M0EmsXsPgp3v
3OQQ1Dospd/CTvdtztdLdZcMIH+NKyT2qEg3HMGEnJq+ve7A7HZd8sXl14+RaAPz
fajE7FKSloa9UIm8aDMCOfL8xGTEce6Ih11Ymq9HjgRGEEw+lp0l9TI02NnC+4eQ
Y/wjarKWJeW0OGvbQW0MG8h8Ak+QlPdaR2rqF7ZOClv7vtFwtb9KRmxDeFcY5muK
piCVrWu8a15mFB1+z3KP4Ym/zEdgyrKPY8lx6qpsWC0EgWf4b7gflXLOQwM34ebO
xkjH25HJKTDLUaiHIOFK9pyqFyK0jkA/Q3RUgtHaVw3905C82waay4nh7YxB9M04
F4oVQuteumznbLGh8JL2l3S072k5w1MmhUn/NDjEgMmNJyr+QZDf1PxtybghW054
WkSwTP5wW1a8ZWXGPnTNwPRU/GleSzKCytINRoEWVfSp8Yz86Zeib9FPn3ffvq5Q
BKhHwO8QDne0wsNtY9ABYKn6/AsoDTOi7zqKOBIXqpT+8cVP/EPsKhbDh6KeK9LB
jPuTVs/V5dEAlgy4RBJfLvbXdvhE4LA7o76FwGmEDt74MFMbvkhdwDFjhHBY8ei0
9c6Wkbo40EN7wjQXordUkJj16oDd5fvjz5b4obpTVpIXVvNMRLIc0+lDls3be2W6
oYsexN/nJg8Oo+B433++FpbWyEi3DtlbXHC/R+5Pw7zG0TTuASfaOToyeb6vhG11
HSDtXHk9k0Np/KNpBgPDMz94KPijB2kmC5ceNux8lzOx5/yBJ4fmn2x9j+K9W2Q7
QaN8KXpfLLDskm8apz68cjCPjg8u3KgHjpD7NLnRD2P+uydsdvWPLt1VpVh9Qb0y
aWhjxyGY32kw3yZIJYPgt/03Y704acHvs8w8/QVBck2sHuCK2opya2UOJOCJzMv4
ig3pfalv+/peZnwwC4VTm5XUirkpwyL4rs27Kq2lC3V7YiiknTkTsNofrX2J43PH
`protect END_PROTECTED
