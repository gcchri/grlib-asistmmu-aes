`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JT2Vo6pC885xOQUMkIL7YwaZ1E/nLlJ/JczI8nwazm2FNUCjJSwUGj4gE6dbENxA
cPG1iNHzlGc9qCf5ackiRaIc/8VQRGDreW5qs/IVae4ABcvvhkD7MKHpD7lu58x9
8ARIjYVMBvYAYTFT/AYDzaNaAsTyhMgNdYUHigf69qL37hZbgeAFxRG7KMsk1wWS
+9Yo83jhDVpFCRQJPreCbWyd6faGI0qtXCZeOXOCq2iOR5qxh+i6p7/3w0D9iWsT
YXsqCrwJcsiWK1Bua2dbRYJgIsgFAo71z/souqeauzVdc+FyJAyvOOb6d/qVjPMq
pKonBZpt5tpXNj4S9fYdU+viv7dvJT0tNT6MhvODV2jKpOl5krWFlegY/DBCFjxJ
dfqXP2kgaRsWc4wppPlLmzTBez9OLsLSXZpQQJaiZ3/MasOFzNLTYJfmpuFA+H38
K3sZVdUY5xmvY2ma+YfGAEMGahcwt4feIqvLxC7bdYE4/62E7YDMMoJ7flj/7tc6
HboIEcc0StdE+R2t5H1XzsDPXuYDkWAzAwcVqNxY28mZjbM6xEQPYxkMgxTxJqIY
xjhmCP2Yf1KZOlL8FNpUsUqBPaY1VM1EpLNw5ZUq9T9TaWrF5CwkwE/EYuZI14ce
e75qI+MOAyFZU1RKhbRH7luQcc9bu+cRmRpsTprOqqHu8S5AWYEVP3RBmlY5vCWM
yQZprtdwPriuodO/c3ZGZ+QZAKCxYhqN9ovlx9ZclbJhIaWbh4Vo/+OrD2pUC3zi
uG/+ck0VWWzWNvDkbIdMUBUrt/PWPMhq0Y7NynPt0ZAtGBIejHQXUfdQLdExOMw/
B21BCohv9QV4RATw2+3ZNe+s/b1FTfVlnI7zX8BCPEH8N8ubV/paK6Rm2t19eTRR
/0pH4mtxrA5TniZcR0s/zkgz4oD1q1qExIFnTVcqFWzGsGZ1jv7rxkBD/U5/vyRK
2GFICAH3TcVUnUl0bNwA50RO98OIanY0XtTxyqzMbZJi9W2j3mEGU+7U0qvnpVGt
CDWEQR+g/XWCJGUivtT9tIjqRy0znh0haZOsniV5Mj0iUAgNPnYKF8rmcGNDY+fa
oOHbrMLQ/xOBJkAXRnMREkSy3bdIhxSNUn3FSToEe6Hv3V2ncIc5jzDCZ5ZywJhX
znWiLAVVl4d8aPU3UIhUDm0k/a5kUXTlVr6o71YFe+XRw4NMT1qFCQD+J35kh6Ir
l0Ha5o4OJSLVZznppNGitrKnMs+uCgpZLpIbiTnYSmVExr6aOZDFN8KjbuaLt9yo
hya+0D4rd1SZuze8gu1s7cwDWtFghojlcb9mkRQkcT3P5pJ1hWNkcWFdGuvuazM8
A7V7nyURTCm0FVH64YHbTTfWH4wtHFLlzIVKvJG4O8xyHCgsfmJPuH1dn3xIbNkk
CuCxeuK5EBlhagiSCt6SqiisHUESVw+mglVciqDkzARYguD6u4EmjdGmwocm9Z2c
mdAqxDFzxwZsStL5by8LMXBygzdAUZ2fzPvG4StQlBQxiu0GBmDtz16sutdz6yZr
ALTKqI8FNJvH51aCqEhNAvh4lb2AtFSxrhQKBEXtnbqjA0O51PTj2uBOF2u+xlaV
tSQCr697CUCu8n/DBD6Wl/9KGCFyzgb3CrL5l9vR5Xje9gYmgydXqR0B6vg47M6o
5clMNSu2nGwDGEkJmVvMO1AmYCZATfh3hdExL6VxNgNM6jTpnZLNdfnyLmWdl9Yl
De8haTx88YblodzrsR5knTQrUBVgTxC/BJG9O7F6k/QjT10ZXsTKrYLFwRYEBEYf
i4x2lDNrYGocYWJ18Chk1kayh676v4TW/5qQtzaird/Rzu/Y3DOdEbDuI52f0E1H
AQxuHkrI1mdwUXmwXGtelWgakscMFFq8W0J7RyN6RTOA8iuWeZXKXpg3L6IbX48T
YloKnJwd1Mbw2mUTpSuABQ==
`protect END_PROTECTED
