`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gsQ0xnoRoNtCau431wzSZyO8K608+BsC9GmtrF9LxQXGOvOq+JXKhZXh2IrA46vw
Sedpnj0bkrgBgHy8xFFzKF+8v3BQx3qgEMSn1qUpa3FjBrwLuFdVQJtyGsZf99jX
a/xIrblVbhStWuwPNqFfxcjNFPWmmrZQqvVw3i9BQo7KLVwQXaB6wpZdsr5oVBGw
gEQrZcY6+vtX5PsYncymuxMfvOaEodnt61xlbiCGjWELd9fv26BGXLxD8yDvDIj+
nK5pmmQ6xBlzHkSypUKhDrjRICLkb7EoaYAcSoNPztQAruBHOLtlM5sXDtP/k0UF
7PycTSWy++j3ox2wIOqF136GjLr2ZxrnmvRTQkkYZXr41Cp3FsBmklyX/XiebcOj
84T5oX8o8XB2CkGsUclcPgQ9P8MElatC8XH8ZEd100iwgqIdEnlbbyGMEj8gGk2W
1LIUVJMPiljpr/PDw0tr602g/pJZUNHbhR1AVvWDjUIyCvthcG1dpNS3j5Ysq/cU
U6xftZ/B+EOg3XylGv50oQKX8MpyqfmT6enaZG7xgxgNxokv7P4PF3+gwUZQ8mZ2
rEwb6jJs1I287n+1huvKNIwir3bwBSJNIey33yZ3/Uj5sMQUwIhuxcvn4cQp1IMP
HCrGG29mKvJ2lLgNQ9Yz756JeeGVh4YFXTxh9gxoVOTxnh3NEULb7dR7B5KP74xk
1hC+OiCNdFMOJtPiH0grzh2br011cbI/SSV/nmQ1kb9icZyF2Q12MFiltv9xrrco
h09rONK7Sm3eT0aTuSSbr6mj3lKqVtkUqXt5EOgJp/NtkkWRX5ABYCNFwoOUygl6
9O5WPLN2wvlRbUUnjRKPcTTvNIPdCp1IZ9HEnD/Dh9rK4E5Un4HefF/J2boyM2/X
+2stDjNCw1mhWIdhNbTgINq07CLjisCfg8jZE8q963a3Yk/p6wm5h/rAYlzIKxzQ
lR/TdYDRQG50Z0422J1GUMxmO/JF/cqLmu3zv0shLbaowrf6sXcbVcDqB4l3ith+
sHHr4KcEeuIVGiylkRWbUFIG36gKQmctuRIV1bYg2R45TGeh5sPEbv2iRNfjqTW6
HGGAahKRAJsS2NhX/684xRVC3cpCkiT0szWEyJZ67LSLl3cfc8AHXE2FZ64yiPI8
6liDGP7KmO6yYR0zRCCE6n+6vFGnzU72nfOM/HhrpwRHfAsau8cd2vt30EwFz1dU
5zIzKxyz5IYtUBhYzOUDJmwxg8/90GG2MSgp6GtFlELDZfReSV+xL1y4xeJjWChZ
GGsLnTKVx/zepj64puuF8cbybpq5e3QaKDnnKMQRnvHfAu7o2SiSSaTNOw5Ung46
XQQmLICxaCcsCgfb/mz74fJtzdVIGX43AKj9IMArPDmSu3NrwnHIDe8bqS4sSlr6
5oX/eWK9NgSSDd7WwNVwPiZko+OJP6d9auK/M+MFni06k1aA0vqbQsJQu6ZQzc7V
SlWsa+9Wsa4SfLDDvD/tMrPPCtbsbrmq0bFE8khAAd4+Qc3D954DlN9tLwWOrNtd
t+KR5GnNBB8pCRdECisk9xuSNHE3DnVGSYXpgcZ1ivjnpgyuaZ1n9X09zyXbTR8H
GtjzOzfy+7S//95G5+uMA8hScWceFxlY2DZDE7fdkg5eNELV+bs4K4VO0smvVWG8
HwqDDHijpIWCo2CzHDe0EbjjFDElzMZHMLGPiTNqIBSKEGX1AKMbV2fzm5pTBb/1
wv0P0WUXlrxSXc0jaZX7VVuQE2HvoJVXiEUseXVQZxeFjeYvly6KRanlvZBfPWAH
AX+gn1U7xoOuf7UAJ47WcmYIRTzTISV8tG5ydPuT2pY/M+CzRVQ9k32NmSp6kdKP
pAzqqKU4+Yvln/VTTbJp2ziKFbYABPN4lmlx7RCsiZwQgp18FSabLAiCQs7RnnEV
C0Lo9szZ43uX1hj5OndAEKsUdaFpcz2gVqwGQPjnplmUmXKVfH0f8/c/FgmFk/Dg
+/fMnn7FKf5F6u2lB4LthLzWBQH3S7rWQvyc+9PJ/N9E6+YiA80zptybbDYU38dj
Iy/wEhu5Hn4JotbktlhRC1BVJm8d8B0OoqabUc5DWnYVCbZZdNdbHSfnLQgXCDTy
gMfYUjORXtbUq4s7cGY6cReuCYnYXCZw9yN2N8WINE5VhyHq7wcIGt1k+1OOENWU
4azqb/0VIoA56IaMTHWRC42iQt2A+thWZGZUZ0DSyqXRXz1CsORrdsGPUeUNBZPK
gzCTb+3ValegcR0YlRJCQTWi/4XZ99JvanSU2Tnf/rmccAP3JxfdCg2MKahyYSaA
Cn710KfDc8MuLEdCb7DXOTreYfj6RP0IAKruAInSuD1T4NYLNdK5iBWFBmmUoxhZ
ae+wZHyG3WLUaKTfSVBWevGJaZRNkw5hvJCu/WdGTqOSzxUEtRHkKQEXM4484GYY
ui3WHMrPLBIEtzsqHhHOTYXKVnkaFUngtVURNVLrj1DOCQyMz14dXsLp/e7zq+yF
Hne3jz28WXQhG9+lDilhd4NuhD44RlCvIoYv0scMDaGKZu+2og3ZDk4ljoMY7IlN
IFOqjNgh/ZUGuWHnbSMP47kzM3kObhJYtcGLPgvLYejML34dcYIC+VGKdJypTi5b
qwY/Dcv+/hzVPKmcCZQhkPYfwkTmlVX0Z56ai6BS4XH2fjn8Nuesx8MS6vlJ/nHL
hpuKGCzBPv+FM2qS69f8g8O4iCzvq7EnmU6xXW7dZbO/93ODDeGx0RMYrmJFlHfy
8STKhwPuNgEq7H/GhZ/spH5hOFYOQgzgcVeRwcgA2FB1wrA2pZiCpXATpcGSwsp7
pNRNPkdtjCcNp5SNwdrJKUObF94PeoBRPBKa5Q9c0wkGvBNBJizHCabYumjbXjG1
3VXwCfQA8FXV9TZmqepmZPneY9h81u1XwwV/s0Bb+AYVdLVdbzbSpIXKYR2Ffcv8
rgzU+eM5RtFCVfwBjAswuMgoqdw3DcNNL3xwhSWKPYuE+pCJXD+YG1kUm2p0cvdu
sHyCTbOTTW2XuhS1Ba/k9CSaEaSYYftqgFUUWvfGGQZZTJ3qsAePCbjQnSOsVkCJ
yYX2AEvK9k+zhMlKKgQafCwz2JzczSoTvjia/WoQmK88ptklxDb+c5Kh7zIiumsu
KEUFrnM8Mk0RhXnN6rPRlvhLbb6o9zqLxzNLS/jG7NFo17KLAgb4VBh5ikLnxXtK
0B99GqLUkWPIYYMBJorPOvzG++JRzPtYQdbj1mt+u3dZk7mOPjRCfOc3b8O7GTDt
G4nGTDWKsiVrBskyY6HHAzMinZsYhbKVDNNm6hwiMk+jbaTH5IuGtUarehj5/riW
J5Ti1B6g9QzK/277Pthd55iE/Wp2LWw4n/ov06P8jh3XCbzNpp1f04E4tWx+yFiK
uieUq8wQ644yP5Gnb3gKKuzkp5GvtKEwkuHlaYpRqXB7/t1/Plzf6U0rDtUG9lQ4
xYdIZgzUVOd5p1u4poI/un+hWXrpA7xZDBuw87deBTSj7YlVJEk4EvudTC3Egiy2
AGKBaNKiyObJxGdNxcPsOap549tmvt6yBNQYShHyz2Ps9n0IWK+BLIvMX8aMmX6j
1MqRYus0trkEupUMtMbM534XMY2EKVQi/AgV93dcl9b9a1Q+r0SsO98ccTTZRh6w
8PIHmaNPNUtgnPV+eQ8BaTQ2bkg+688AItOlQyrzC9oaQEAdI4usblHioChTNVrp
AXQfvvB/eOUOJGAtKXBfOBp3DfsTJzMyGGYIsPTVDymnR1JyTPW4UcqbRN1iPOPh
gUop6jkuod6QH37u28lqbofrSDXZsCiR8qhDCaWGFvxfhSI01lZXAAXkzc7DFAQJ
i0i3IkA9Sv9Omr7L9Moamu69eHXlXqUp84oXiN+UVkdBiAf6P40D0c4/WmZgh2MX
qcwBGspKRSLfDUUpZ5pNubtD+jNdDrOAkS0NOmgaCeXLlI0HotKOZNjtMDNGtmpL
AsMnnue72UeFMTTeGzPYd5oE/OxrExOaPLp1ZC9yPjoy1qTEda7s6SHpGsNIOdMG
HeU8yYLV15Y8RF0Fso/WpR5hQnHeO7uoh1d3eAbUmtH44J/ijYsCmBFa32UvOnXq
rFKZCfMy4H2m7F/s4gmfAtiSsgypMvnsw9pQpB0H9CBBdtr2mI+OiYffh1N+2LNo
xIjcMnYXmUh+s5IfSKd0WSf1Z6Tze6Ecz7MEgGk+jwsgQNdhNpbo37WW5UPx/MFw
hz6ZSXwH0CzZaLJe1uJOVhVhBBuSZ7X7rqD8lkeh4q+fUy8DN0QYGM4NQGsza2MJ
XgS/q7ozmXGLBjnpEK8H8j3MIfdM02NUsvfg8tpyMAIy6nh/75Pn0a6nhBoO2rWz
5rsgtgOr91myaCeqVuya30yq5VgbUsK8YXaadARerMBugnxqlfqCPh6ARJ04OnUB
4Z+VEd7UVrv1QqYE0UHqS6vpzQxv/mMAZmTBhpgTGL47Cc3dnYDdgF0t1efzIQF5
00t7uMagY1fPRdeTgcdA5DG6gDQnHyKEabk8Nvq7peZ5naDC7cSExL2ciAapLOho
Bkb66F3hV2Eyd4Oyf0Pntyo6aEW3ULJ3sprUMpUKwwp+qP5tQ/2njNL1P+LFWyaq
EEYcozrDZhKXn6fBRkpDheA6ZR4ZekWKHehBT4qiT9VS42acs5Jo2FyEmbs+AO9b
7ycnMzgNGfevk5g4GFwh6bX/7zIYcL/cLhX971dy3J6iyVAsgpUNMTLDv+gN9a+s
sV91ENPEuXaHM317WLdmMgxTP+GhOCCmCqIYn1hHMse7xzG5wmBXsrChSYQyKsif
wGeLv1f1gHY1t+oQZSmP9gmiNszyPWuy9lOQfsbp2JW/bN2ktpXjn3y9MpXhHNAw
DVh1pcV8YS6Cc4FxYYgczxMfT13pZnCxbru7tUIZJDWEl6Vzjy5ExtWw0U7T03cc
c4UfFFBM6ggi9S4/V5J7nC8UuHwjccUO1ySfxRnP6bRDFa3dPtqQ6NJUz5LgaJ3+
Cm/JRAf1RpUBZFHT5pGLt3IdvHw5vajSSnhwSkgn2WDtD9hzIzo2SjfNlRqXN3Rk
FiQ8Y1bDA23zangj3QIgrXTC643XKxC8ewUDQYdJOrfxQuOpvptVR9l7ySmlSKt0
Vxp6dFfNb2uvxezfna7OAO/FKzckWkpm+rug5gyqQQvZAPr1q80gyfn7XogMRhBM
VnDDn7283roIx3Fns7D9K9sI6BwB84K5WmvkWkNDrGr5sIoPzHjCWdX513VmNwJe
7Bks1vXWBkHvEV/E1xBfhh5+9qUMRrRRil01UK+59X3F4ExlI0w2kD5K2gsyQQph
h9cjz6rQDgH3Ampghbs5jcayYOlsUFy7CrdrORQ6FfxP1Xu0WYibYVbV5JCVYg8n
8KnxoNYZ4ukJuUltGEuoUPc+Ma0YoP7Mp4xsb9i5UTstAcOYJMQ7Ex5Nh6BkvoO5
+0QMDcQfmRLx8iaFJN/xA0USmAMdIfAZfwQpC7YSC5HLcaVplHtmWTMC1yKqGiWa
sfBgdLumG/l3hTLaz2vwGCXGXpYX25Tgzy9/G5zVRzoBrG4el6y5fYL29sAoIkh2
a3qeYB9SVCfHsPttsK//PURJqaduvlFNJYhZVb4Z7LCzQxJAbo7+xOv9Fzdf6Le9
/nUTvpWABCMRnCqZ6Vi8wYz5WsqpmvHg7iadGR8Ah0ogJFTD8wZBc7H6cL5OKA46
K/no6vfHC5Mdzl5j6IOplw9PE+HRaNSQmHqg8RbZEgDHmjsX6FXXAh+DEMIYuPKG
HyVkwRjz9RWy0Xn9xqU173fC6+/Cd7vrhwwGPbQ3r8FkCg9pRm0xswF/Zy/cnsg5
IPv3J+fIn7dOktBcUENyArM0BZX7JIV2exgl2FaeDWaQ9yWgjD7UMkzXFZj3Kcee
qZ6Kqq55R6k8AcbTya6IqWJt1Y5XnemGY87mmcU3zIoqhjViHaAxIfXxRj9daGvm
9T+lHxbpG9Y3XIuwI9ImugpsEc0HPCdQjAdJXpUlyN5ifmIZh2LpQsBbalJVWSZ4
sbCvNPsA13Qx1twBq89c92n1NEALUSBaJKm4tXzwFVE+LdsPzJoimxMT4oRZTQSG
g2+dRCTSyv8mk8NNo1wA2nxgi2m3PWWn7OYOrccAAltPqovCJSpeELTC6oONqIZY
gycAzKwenefgE1YAvXJGAFGRh/45HCNUD8ws6Z/QFa2FINZhgnGGzLXM7UsAuN81
OvbcGxGVtm9nS95U6HMenpWb69X/cmzIX8uLqXarDFF5SLURb1eZCm79Da5vi+nM
99C4pSU2kJNZjLtLJLFvH0qXzi7zkKMJriFby6dJGOXl5Gt4EiZ5ko5fBebX14QH
AinkfEp3tgW1ttrkFBN92qCQ8wBR17x7QI4/NwDnAnZfXvRFL6ovvk3l1gdg6MBK
Winza7QUYdzKvCPKkexgMsGW81wlaEhfdxWj34aHfVoN4zdWTfl2+ORXhPmXJeeS
pXNGD8uLmvVMg+Hy0Sp5EjRjjtyxPNgba/Zj+L8j4xyL4t2vZeRAfF2HvJXAVhII
l7e8EnAttQX0mQYcORPDu/jyjZK1MJu1tI0xFaSLYf1mSd3HSYeYrQua4/0DpJEp
DdjKohs6kx7a4QBfE/NL+jMSLJPthKrs5pz0qwtV5ZV/SvBYKdkA+XSq6Z2VQWal
DJ7W8Ue3el9dLd3IahGATjIrYhA8s5HPCmZWKxptpUs6dD8E0BC4z9SFIQghjosS
idgOitOVTp3TJi+yKEjeAgD1uNDZGcLHHJDoCTPiyyWDlhMg3/90rL902q7jPC3X
oxRWjUHy0jMad3kwQ93Sob32Zg1aajAPIgxsB4OzkT9T+aB3Nvy+uenADtu5CjvS
MuoNnB1lxVrrFrY5BTb9NLngSOO/YfVzYKYjoxFi3KxtCuAXOnfCwC4HVl6Fg7b3
KyVOaYYvGLSphIndVRZId93i6aUQZhaRTaQ2bNLlrnkT8VQoBlNmpyLf8UUMMoQH
HgZw6+KMDPHIpotYTi9jYiuu0r3FP5g5BFXni7GGfW0JctKnXv1/LRvpiXikyhJ3
DrtsmFYg2/Ifdgb9P9Tz1AQVV5eXJ4wJJoIuZankzegts77frcf3Ts25prB4C+n1
r+m61d6A6sC9hyxQRFJRN4sY76mJM6SowRIg3fdPBCUw9EW36ZqY2iuScRkSRl/F
kMpg+aayIzlIAJRf7jYymG/Xbpd0qp9NYRQS4mzRusNy1Z+xAtVouxMiJNmuq6UZ
W1e2UNc4iqeim1h6MQx1XmjtD93MI30hADbYNuENN6CsWxF7Mnnjc3gQi/Ekayxq
dQ7+EZ6aNZi5f8J4Ta/CVoiDNIX6gz1vp55MnjQLk7HFBFgkNnFebXkX3kaTbwjK
V4BiSwe5R2JajKH9C+v99HXBvxgxPxQBJN8s8rb9rUZsQ9lQ4pZuFekyTC9Nwplj
TPUiJ37XvxrXZI2wdgOI6S1AKKE6KFRwBDAUl4JYtgPVtz5hqms95hRFQ+nugdnC
iptjaxDH/kavWFYhP7s9v8YAIecFTZkPcPyja/Zrc5E1Nd8pT+UsZmQ2TQLRi0rm
Xb27IGvAbVHt0CMZs+5MdxcnsA4vvZUouhOhpHHUrxv9E4rb9Vgpr46z15zOA3Oy
rtEhMgBiyb4jopio6kC6E3ocrLY+h+POBPO11NJwBRe10fYgyYNEwkODDAFZoy1o
F9NjjhxGBfU9Go1Oi7l5KFAftvZIWE1pkJwocaYTBgJunJVG0L4knSIwSU/k5Up2
nGAp4mM3Upefb1PjhreQysfluv9K0IPINgtTyNg12t5X/wnHMvz78WIMzG8Gjsm1
oiNFJfGqLXJ4ofYKVSPTIbjORgGImVdySEdUE+3woXKxmCcyTbpm6eaz37pFsQQp
vrXccefMJQ2UHcOdBtLBU3BLpEXt6zoVBOOTC92RoVxeajQIxnKCPY1kTWDlzHag
cp5GT4cNRxEFqjMK99BBdMWCKHf5HRW1JOB5s6wlWNpV5LsR5h1jJL104KYIyBGx
eKpDk7bm9EzxS9f+Hh5N7fjC6CZbttpHrmL9hyZBEL3b96y/zNGBGL0ojeZQy4SU
gtwomCE11mXBeElZT9ogvwXID/oG8oeDTNrkDsAy3RApf6fC6VEKseTURjJwgewX
2GGPXjXr0mNgPOXznW4IPCF/QpxmeLGczbZ7g2ZwalLx9uH1zkmk6RBuaHpwntGR
O8Oeyhael4TzBM6FwLH94XFu0wXmSH10a1wgxZP2MKkyDSlxnCDeWqok+0uKuiKE
8TupEwEI3dgB9yPtW5bo4D0rwtSZBOrXG/nVxtKK2s3NYJnX+oCMeZ/ZTHY7bmTd
cO1pK9+zSphAP9NpneqmQguRZilB18AaTP4O9AULyDJr5KF4fGtqi/z7sYBrNTnI
jnvog/9cLVP0ddNlL8LXVgZRVnld+BBswJhOkuATpTZ3mv6FABdAG2Sdb9Wysx2v
wsjUAJQUY2hJc166oaGud997bP7l6lWOYYPTNufBMMSKPUeTWaoFlCrLwcJgWrmY
YHKnPS/R1u01fT/7W9VYR81oe95F54kXAY5miy4+fSKL63d9mC/VoVhabbr3i9s9
FJma2LU8uBFbaBJ97FpC9CLdZ2RKAn7JZ4fRIOsnpvSkLxQ2rQD/RykzX7ZYagoL
eO2axxncp3cCE7RZHpfoWFpgOpTaL2vu1Zl85on7yRNLx3xw1DcGdU1/NPr086PF
LaVzdbNdpZ53ThTaJwryEpmmvIQWRgQNhEcyn/GDtBl/4cOKiNbH5l6UY8BjcbMF
uWTsyevJCti4mEwkHQXJwTro+LK0KmkgQFUwq0hupVSBK2AiEGSb8rspn1W6LI1h
bSIrV066asUq+x6TQ66LQlxtyYuY7gEAHvqxUXirdvoqZHlSE61cVEAzRtrp62/E
DduaT9/dINE9fbfaqzhnIP5a5G+ntKFKyWpFMRQSXupvlOJRFuQ4fPGy7IDUQuqN
jvBtXu4NZk/Q1XYE+1ugbbP6zsdN9a8hmBWsJnATIg/dSKGVWj4/+RfM1gP9gzuP
QxTCDV6lwD4eUxJT5kR+alY/UchLLdRVQF383piyaT5zaya1TwudgOcG6Bm1JkyX
mhFEHH36UZUVz1jGxO+zva+UR62YEb4rN/AtLdVnc7sfVtORlaoSvghbSf0MxAE1
k0mOSAKzBOcjV3vTTIxfi0Nn0kH29Z64+E0fLYL+vKp9yLHlbX2DHapvUEeNxGGv
T+DugKUIxF8YQfXidX+PgWc0LQsVW494MAvA61m02aW2JEsvanr3M6l9BE1dgN3/
EbM/xg5AzXkkYMjMJhQKlgDTNtU76+DNwjOptaeHC+ibc0OSEAg/YV8nSludwSfK
zIbdRAceOZokbwuV4cFlve4yM1XAcEXsI4cqJ7OpcmAKq3e6r2eCtlyxO+kfDTXt
vT92La6ikLbYuvQY5hfkvK2vQcDXYNsTcKSjTiBvqC2M5sNKoODizlCdNiynh1la
+ZrhnCUiT2eG5NnKcvx3JTXwVjoEjpxo0MSyMIDAyx4ZZ7sHNEk677ih3bVneyHL
Me76UtLl1vLbjVMOSdguzQYGFXycmi77pE9PFppnxsqOxVZrwcjBMEENQsdAQQgd
2SxpGUkYXk1AGFQjAVmJEKuhCMxj8l+5+cHZyMX5mCjbtIAREJS2fGAf2KrpoiCw
b7ZxOmmBORmqt0J3bsQjzp85b192cRMAJAfP0MM+joP5ZYQA3RPs0DdW7W8cb/x5
DpBSimLUqOeR0bVul6foYVz3ERfgxPFaX1BvOP0WR8Fa7m5rKfGJyiIFLf9sAPqj
Ardkm7kB/AFyXKhUveqhbL7v2Es3RBYS3eTBr2Yl0p0HLDQUl57HAC8Xs9oUApUf
LlkxA91qy1YZw4b1Rki20t14a/GjddN+ZKrVAALa0WHZg1QmE9dgVLjwX41OfcwY
UOwz+e4vEON7p4z/lscTND/FJqscZXWNh6NVhruotAdCGlPoA0DiGl4Mm39jNgGV
m1iRusfyFeYwG54ikXerkkld2pBIuvsPJSKwAp/qTAHdgq7P6oCAS8yNd+AhwbM0
OBfgGc4UeWcdULs2Lz4HI6QN/MxL/zRSwvkA/yWk+UHuqulrAE9LCLO31f0oqi+B
mGFUkLxMx0TdZTbbrb5IPlGm+vZPsa6Mr0y1prUtxZXFRlCvyPvhYzuypsrEHw0x
bsdCb+1vnTQLt9r0VHnv0TDqIGLMJrhFQW4qXDr2aFE1wq9G6shqI6x4U65XD/Qg
KFTwDD89mXdMmwy3Rr1K//Xsh8Q3LVxAgmncZUgGr9pHpoOmZBrBPqHYgPNoW0Q5
Vi2ZHtTYFtJFS9Qo/UWRJh4QrPm1NjR+H4u0j4qPy8JYbGx35SEEmZ3+ea8nGlqI
FtRqhoJYO8E3HiWd++d78oGnbPHpRU2P6lwHujUPuitcgUwXqPa9AXNiualqUxHR
JQ2pl2L9YbBIGH7d0EqKdty3A0aMoX6lMlohDMdhU+PiR30DdmgO4A10DufykcmJ
DIvbd8p5qpSg/S0S9IGufA9DP/Cp3VHw1cXu8XjZXGPRhuE2sKsFNhqUDGgSU6nO
hTdyzRgTtK/cdyFXSv/A1BdvlSQYkyf+TIDM5uKvQQpTg0lNM0VnfPuuL02jvYEX
LiMjB5dAaLo+rRSNLo2qNpz3Zdp8uiOEnLLbvbkJraNENSluopVkw8z5X9WSgkGN
P/KBe0I1zQ4FBeLZgqh6yVxgwNECKEIIXsUVpcqrF8bvucE4Exi/qzyFU5gGL3sX
q05F9cDZn/inXGhUWsc1p8DuKxkKNIoSlF4Bxmm0WwFhL0m+SL8XiYVW+UHgMgwi
OVtgy5O9PI7Vp3K2ac5Nr02aJxNcmE1KN6uWeoSQpxRacstQFv5bqPmzqYQYfF2H
I//k0YsXmQBaBZeoR2W+9sznN6WcGEHq0P4VwM0rwob6SNdyxtOpStLkzkWi+2+I
KGqlVga2sEDAiZRAzdVvRQQ9x3UkoOrXP4DhEAAou8p/7dfSJoa+m73tSl7Mauny
9SVgFt5CmwQeoVRwKVgY5askDyJHXuE88d4NRhQ18W862g203tBtJbozwYWzJYMb
06ckcPpGo61Uj3LI4eRYpq7wnb6ow+cdfazIMgdDNvvfGaVwuczbwFKMLt3wx0DE
yiTWztptlvzDeqelxkIoEcLcEcoj2yowaJQY55sVKFAVFj+nAxV6DU8kVKSFeO6R
Iuz1orAbfBDWPaUyHebTmhykd41vfgm3UEHvblUYPN+xjWYZb+NttGJeYZUXJbst
h2o0pXGYrHPiStwcDLz2x9WvFN3JsAtcFVNK2O3CltQet1hCljJZOZO6k251CqAj
6GoF3CC9sCE/SvQpeoLedBr8Nq3+R5MqzMtygYgujAQuA4LE1w/nuuJtHy5aE38l
XCV8RFIKhKG8JmeviGlNOcOM+mRNGE2BwqSNoHpX4Nud+Ohosvscq8L1W/JjVJAY
I6Jw2+Uaw0kU6B8FuS0TFS46+d6pZUr6Ml3yvI1bikNCxC6vdSHYtbJwVeTo5xi3
p5CQxmf+3zxIbAcYuFtlCIhaIrSmWQn84UheX7SpUm9rPEAAckI9t4t1gO22xG9m
uzTpBCOkE4Ark0U5iCRaSmFvuDWFhxbl3KoLKvhk02wDNMoOmkMQ76z86YR1Mrt5
P35JZ5GbM/Dt7xuHDwHne8AJNrnl4hbeD/EZfxZrc5B+/b0N3aXqPQjYJkc5LniK
SSekk4dqpxlwLXiyzT2sfBfOw7ySpElZ9Adlj+E/MTbW9aZAC1RdJO+HmMolAx8U
09meOPFV/dSdKMRGvNYbWsOdun5OTa4SNb4hnk9UBjQUKAbtJ9QcGI+Sp+G2I4w0
7ktByfUNTgpa50wCWx61FVGhxA+PrgbX979p7Qnpx6HHqOrtgN7p4x+5c4xKn1ao
qgTC7bY0P31JxHFU5kA/qLhW359woI1poCevyFRdU2RJLg1yE0gL92qX2GcUP+Bf
SXVSt6a3lGfOiLQoGO62GXpaUOCcuUULzeYpbNLVU8qLAEYKy9G/aTzDCG288dLO
o4xD6Jgz3Cjma2oQ6qp8rirF5YhzrDY3jqkCo+tczNFuQyE5SzG2VGE7t7H8H5Xe
bcoJrF1KdyMF1gAtKccGk24g2EWH/xlS9IDd1yN9ADuq8qs85KBFIir258tnPQ9F
Myq7Jk89eSm3sguWIcp5Gjm26d9kbcAdzO1cbRybCmhA5wCbq6KMZRrEx4/6Knn8
TA+WPubejXnumtNenys4OinXs5iNG7411ABtPiNeRKUX4N7NM5C/304CMAJNnxZ7
mhHxbuBjsl7wV96soBriAoFmIMFuc7yf1WvmAFPeWAzFY+Ral0mHK9rylTNm2RZ2
qoXTyeoUtuNFPbNYNPLhWUflw+/fP9bmi9QFYCSjAM6b9OdDQvG6+/eIftnkz8p+
nKFQx/ojsRWsHqmoH96HJcMAM0iXedE6+z6OQClRTB7oUjP5MrNUs51dvhi7SsaT
Jqimu/mHTq4r8fpTqiaBwJtcjNvxO5IyYRElW0hZuUtUVf0amzrt2eiW3vLCsVbs
P8zX8DFAGc73pktCXPhLdtE+0SzKHwQBeiwAvpZ9zprgVJ3WbV4g76xbQSSvwGSm
wkzgTtVQBVyx3Ql3F3fC0fxHwRHd4hwsBO/a+zjYdpbEjRibQ1ZtBZGXfg+fOVaU
eoCoUboAINLtU+OHn8PoAXR902+ro1RZaZ80SuYL8KzeYGfda+yrT4ke15SycFNZ
qoWES5UBKD/9SNTfl0yDYphPP2HaPV5uMmLPrcTSmg7X5XW6B2vVloGXSxCCnBDM
jNofu0H9pTpiJn9fHUBMJZrELOTvFRUw7GHhYoOZdRXA7kuWuBAmBte0++MV9CJe
1zo3/92UiSUjLWRYVQu4A4lMbFBZnLqEe3Aerg4pRhMDEfhoj1a/nazEsMNedarf
+X0UFw50zXjb9JLwhK4XUOokqAEsvY/wfETQNm4iNVd2slyeiZsoRVKZWCmdBzNb
zYrLy5G8a9IVaO4Jj+88gEkJzN8F0fSCYc8I8bt/we0bDIRSLRakJijb8JK8DIEe
3wPJWQgRb1FcrvzxbvBZ75yELZz79y9Oq7yZt1AImViPqzMZscl7EOIOY3E9FIzX
Zm0lz5Hp+OySqV/Lb3ZirTytBEmWn7apMorckPLrL0tRZalxjczlPj4cBvLHwwQw
rGQCSW9XsCEPvQTb+Q0sXyTgHJExlHuzWir2prWfwpxlyYm/qCWwv+6ySmbpF6qG
GI64uCxm7c1Itx9QVApSjhu1xXTcd2YCt9oypQScTOTB2sVxh/nheMEgp64s6HqE
XuaLKCAlB3cVPv4OJV6yVZnRa+uA0Cs+O3LIRKrR5/MrV+sqx9h+RkUHx7dnT/II
Wsvidc1ZTbuqS+tcxVNrW7A9GmY9O3dmx1d7cx0F8zHh80tMMsxS8kja6jbl7WyF
89lard1nZuD8JRi6xEfwB/jb5abiyuszqLU9e1vwdqTDWCNA6JiptxvXr5Xb9InI
QqbcPd7MGPlN+v2UKx1eh4dg6TfLPmp4PrWB1Bzj6InY83x/5KdK03hF6gln7jAD
O6Xs44I1Wo4lBBQEz6x5STnYC7LS2eQ6uYGf7jWZlvMJuAuss/y+omDR1xuSRdOB
3VU2hgisrs8z/35HMcivNIsCcVsEHIVbReKUyBw4GjTOzx8EHmm/zjaxUxUdfFM1
S5vxavBZZAVc1Dy6rsv0ebhui5b1wtPqO1j2639+4UHBvKRzCt5ZME2oJlNZX76b
ctFA1t8r8NaliwwxG2C0d7n/XfpW3iUiF5fPaE+TceDhKrCytMICnABdJrVn90yP
dUdQhn0fhLlrM/KcR+U9Izj2hr0MoOYgG9EcAFQhyNTaC0sdZSzgPcGrp+EwCjAD
Bh+dz2rR170FqfQtjR5E7Fnlsp/0we5aBrl6IHFYZtGr04ZdeSINA9KOSMNYVoFe
2oD7HRsqMwgWIwSo+BVBhwE2yoXGaIprbeKStoUsMU9mv5yIWzyt8hUr6rn3UqDs
kgxItpSTlWWuch6rxOg8bKIF8uIE2E/QWkbmFKADPjc2VnyWNpEWqqUK/ev15KrG
Gx9PZA9dHX+dQJ7gh8/zr4TlFDDg8L8KOdg32qz1ICXWRGTr2u5PS4UDx/pndF58
JvFG8FA3PkQUKzYZVrshEnJb9UGMRMTAa3GbPc/xbLAOZi3C7BRhFGcsfP9aRXyK
TD0SIaLF6sh48OP5muXAKFTXPBrd60vEqPXUVpbTGGkyozH2WCq/EoSqLg4LS5mS
0lNRbrohVl+3zsyyIyJ/oQ8xNSoiH7zc/ZE9vDWTpeSVlagHfg3FpOyglzZw4LaJ
iMaplUK5K0oDOBjceclDv0Dbm+hottQT2gSSleMD2dPQa+7LB9jKEOqcXowRW5oo
jNlSHuiBypw7XZnkwoMkgov0gGh1PpFRB/jVpBQCIELGTVIu4d7g4APu1jTFPw6u
CBFMhljHLB7DV2qAo6zhRqGclSGcnrEAVVTHz6IgeQ8TTnUeXQsK+usbX7RlUq78
ELzcbb1jVX+78mAlCrhgDRg1cdRmGreGiASqPBpL4bc+xRLBxrUPMlgclofBGBnc
sPKrs67DUyqL1DBoyzATd7Rto2ZLx4/sFNIOUdb/okIZyBg2VXFFzIZ/bumJKilw
00HUpLmoAZD/KopkL4cRCmuxcg2UsRQGwHrrpbobgn5YWKe7V9FpX7mh2m0FQA3b
Ar4T1+66mU545WnW10rTO7cJA4c1csxttCAC2sCUiZwjZ1Ug5i2GLlELZMPzSz4Q
e9PNd26E06epg0X6F83NM4wwM5kkIK/3fNHGvo/QOei+G7nx3mwSETLScqu3f+Zh
/1Tbycn/8Baj3P6ZcF/EFyaYgkmxNOtHizZqW+wJHjBFuaKPEWdNbjlfAZSHLsLG
zN+f7AhOfQykcLmKdVrDn5JdfE5RxwwCt2/73XI1rQhOFYO6+dP/aJuvg5K5kaj3
rB8Nj16EEOyxABfIbHXhadX1l/sGcCVuaxiFkPaAn4WABXzcSU7dkrvudmi0kEwB
Dh2YrWl9q1c7ULP87erbFsU9NPfSVv/7zZT15p2+GXNrEYkTVs82YzRqIyjNjyUP
h4Xlr6JvoPVVwMF50vZpCb895U0B2UevuJ1t3mQupj+fwWYsOTZfu/6xwHEMb0HD
IiY5UBtpusXFddZ0tVeC+fBBVwZUmeSjLK8tJRMKGwRAnX94cDSR/J1UNdp+5u/E
Nak50rbQGsq5Kt7A9iBKnPSymgL5mJud41oBygVkypoJ9iQ5sbqL8UWvUwHgbsQO
UuUILFNwQAm6obxzHiCGLqSlLnbVmw1rBaL4HAN9Poq3c7l+IgXJEuuFanZrt+4C
X3UHf9EqSWrFPeoeLa6KZt/UM5xOSCVwAKf1glhIKdI71cF9Hbepp4iYOIxcnPZN
iNazeUJldNCr8bEdgvifG8/H1QigYZojDf+vZ03XpFs8UJq7X59WRcG3wbJApIot
tT/N+k3rEwGLMRJLyOadleic+8ByZu1gIp8sCvn8PJbQ7QYBgRSR5pzehx60RTC7
6R/L6wFh2BPye8EosoGsICEglZjQbAiqjGFLgqAAdb9tyEQbWqkcELgCnQ939iHE
GdXs/hY8gUnvCSAV0EyMnmqUtj8Cs2ajxgo+mYqZnKz78PVMDddcSBDyjH8eP6MS
t69rwaVOEJx0LNPXJGAVefYnJ1FGaxR9cF4ROImgjSO1Kn4ILNMh/OqVUJREB6rd
e/nAth8dX8vTcZ/tAk77hn9oW9Qft5Ufd6ffK0ROQU9thixhWgSbOCpq51Decx24
7FAkhVOirhiJoGPRV2L9qT7xap81WHFJkP4RY3o339KFuMu4rHIE6e0oN8iLm1k1
HwqyrZBfTjDeR6D2i7L0RZsIfX/1ECogAdVJlpD5MwsGkyoN5b28l7Kk4xApEIYs
FZStmY0Nh7gSIHA00JyVbzXshB3PfyfolxwaL/Iksb9zQ/k01VFzW8+H8/kKS5zO
xhXX5scQp7Un4EYYJr4X4V9Xg60YI14oCT++nS2wbZeQjvFvxn690SBAsGCE4ojE
oky6slW7DFnj592EYlggXtXSdLPBGJ1Usc9ry5hGQ5awr7T1qKsOE8fHVfVj2O6n
xds2wOJNhxGomRZNjsjh4v/mp71HwhHikWJOVMyrG+QE+VU0Hk2LXFYVugbEDkT/
ecNLfQvEeX++b4jYxk6gXl+EhDeYdcWH23bu7nyIAWmzNzNcagva7zGj6TfI8pzU
ujBXt6GJsOMAcmoouW4ml8Ivn4UftANIPV6YDRwJcV5qdSqxlVbns9Ia5husABFS
e/+W1lRbu6ABAjsaBsKMBsLle69pDBm9psFggv6Dt0+vTPgLuJc5qQaQ7qGS0xx9
JwcD9Io7rJt/3y6GsNFflH0C2P1Ve+cqMC96TT6m2GH5WFzJxjwiAcDb8ELSkd7Z
ZtdBavWt1st/n9O3qKh+Fp5XJ/LC9PI2s+WUvL3E2Srq9ahhefQdChpOlRcAXFuV
tQqAXB43GPgJhzT3oDY4btSVijKdyDWUtnEuvuA7Npns9Ux2V/6JB8b30KRfoVPw
EZSEH8S5qQg4AoaV/wGsGK737QJ3jGu12m0Wb5RmZufTty5jW/k5HIR6hwUWGpNb
r1lbIspKDDk3y4cAP+WsCBIH7zNlbGkFlX/h4WIQ7r2d/N/26X0rfmv8/EZCeVvY
iLIgOe1idkEMq64Viyb5GQb0Wh5Gw8NTUpHV7eS7c584NFR82MlvdTSIZ/0yvE4Q
wARNKQmyg2Q0VrZ46aTtSadH1fvtSJTXqGzDqNyaiJIZZcwqvxSALRu7f3L/8DmL
2Uo9PPGnJbT7HguMPQJaWplrwNE3Ns+ci4iPlM8F0Regf6gCe7jb8Bq6ymurhRW7
eCvHqyHsawxmAm5WO2EV8i229nylM/0iE1i/pIIMTWihAURvZJ0trDCRvIgrxQKF
cp3gL+Siyc+MJChAzYpCKOQb/hlVExptipq9mdq5/cc5Qjadm0d009cLez+pj5Ht
X8x7GulzCAeSLgFJcswRnJTC6aOZLATvUP8NZmBSOSvQyj/+vx20TI0zxelzSHFl
p+5wCAHLgPu7B259QKiYcipVNhzoRzxL/KUDQVPbFCs=
`protect END_PROTECTED
