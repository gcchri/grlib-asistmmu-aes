`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DOyIgHh3BArmz+WwJ2JG3s/7jlbVvRY6yJD1zK+e2FCC8hvbUl6LD4Vcv23K7ULX
f3dgYpShJkmA07rD/HVUZLVOyUMxRU+aQSxVDRF7Qf7+ClfddOjzJJ8aRtXrZEFi
zw5rPJeGE9cy1WFFOUUMPaLaiz/ebi4Pn0ra4pQEv5dF4wWZYHtava1BW98EHMCM
/Cp4YcRryTHisb8K9w4ZpakOrDHidL1s5y2jAIqV4qhJZ0uUWEc8Gnz94DpTQPkT
2K8lT3InmPKCLxhEA8SRYtW4Ph9eDHY/cdVHHRRRFyaBJZgfaa2ilrF2Y0mC036h
dKrI/j2p1UBxhmb2ICPTTvMG8TH1Bf9ZjI6rq7UIPHwYijxHiYAiCibTajHBF5gq
Bebsi2XOqHYXJsGjF9xfM36Xr95c/RJ1NgolfEmXZ3DlP4It/7F5VGiXphY7UIn9
TqgyT+h31bqFnffDbuJ2smM4Lc9HE4wk6P44MHwvl4Gr1w5/08rjf5TQe5IVMOgt
L50QeqccArxT7y7S6BlDdpLjG6z92/neyP5O120jkYF+SkpTgg2DCS3WrSniCKYK
/cKw0HGaCJukgjMUJPg1g1EgOkWmdZkFQMHvGVw8T+lwOiEbt3KzkmnthK1mqmDu
ZPLxGI2Zvb3jfjbaZaZXcLFaP2rZ4cakM8qImvfCmw+b5+C/31NfHULyOGnCkATK
rA/j6FxPvYAVjM5IyI8i6wk25lwKGgEaCiD5rfNi3oH3fg89GIdP0GX4X3rGl1N9
mnq1zdtNEJHmKHfMdyNRpX2q8UQogdbsAN6hayUacQ1GeHwji8O6RNh9lj9NIsW7
EZo63dzA+W7lZROSWITfIuzKsTxO4y5U9rG/7mXt3wpD35vVLISI/vYij/zwPd6j
AXlN6htWNPe1jpJoPM4drtD/UZkpX1qiqx/eEHJe0sEqkdjdA9ci40MsbBf36aBs
eoTKu2KpSlzvn0mJzdZ+2vS2QKeM+lwv4MhyCxlCXJ89vcAlACd9w/1brIB+j+Ph
Xj0S6pATfKhJYrzGv/MfZtudY6Y3bWYbfk6yKEoNmNNpMEl4p2QIXeY/5F1aiyJY
ckF9QkvFhGphOtG0Y8+hymxe/FGA0rsfNGSE0Yu3Y1Zw8ynnRY2pfkXDRu7EDdVJ
YeM3wB80KGe/5ur52mngUcCUgtR/t9okZjcHECUAfIT+FhHsjp4uZPUS/Be8suqC
tBtForJ1DUWYhBZubsl9zFLAdao5DszQoBK60k33c7YYh6ZAp6G7tIhlPTtkEXd9
kyLibeP0kQjRqDgUg+G/PPZruCyJLkpOfkWHIw70oz8YRumTqs56USX7Hop8Nywc
UPCslaT4cP2PkSCS7KkTSKo2MHz8ZmdxlqoBqlybMN2zOhmlX45ZnJQSdbrZo9Ih
IlTXi2BuxSzneJBZorzpF6WoBpInuVtHFVdaV1A5TwBZVPEMTmRWoOXN/aNu8z3U
BGwQOsWzsDeQteVfVimZ7v2JUCbEHB+zyrctuh/hL4u6jQhhWxsKYGWX3npnjO45
J4nrhE1Vfcgd734/BX9gizuFjNToMXFK8tWJg23pvNbDA9ko7l/gg8Dvs0Dx/h/U
PkkCWndQIqNLG1MqWh7yUauELNwo7zOa4g0NAEFsSeaqkKcjeYmUj76hn7399o/o
trqHwcK8494+srLgPBIIcYvyWG3dMGohGNC6qNxru/vdYKOYKIc7kwiTi91XFBYq
OQd4vBFpJ+Tv4+97JiTq39iz4/mObGeVTsGgSQiv/Uh5Em3eZS/gAjxcZd/yizYl
Jgg93T6RXNg7RyWvEUE+P9qI3rA/0IwNdx7i8zeBMx5hWe19djyBJj9hPlLdV6au
vqF1aVVBmdzKb+iZGw4S2ego8vxWSMmuqKJhSYO6tdYZrvWmMBhgxVgleiIOwni2
ItaVKIsLtJdsu0nDTaPkLRjfFNXRQQULRkKjtYxUoX83aWKSWEAAtVGSLJr8vc7r
dB7BBGbmkEq0GQH8YiFgwmXg6/tIH0DJyMEUyUXVSYBuJ4bYMZnNQJ5I9XKLU1K4
X1Zu10qe64SnJzTaVpTUlegBnWSNwYgLOJYNgsZLNgB5UqRTBh4zpue2ZA5Ns+30
0idsxolSE55HrO8bD/QBVxIGXDiP2itFzOon4RCdQ8jKtYb1v3ecX1WgkLEv/aFj
9phpobB/kmDC7d53uv6p/UuFzmLU/25PmjB2AIZOOAeNMkvbg3le8BxctbDmG0ce
+G3RJVTWfWRt3GQpOJf37fKKHzIaYmW7z/oKi37+WGRoNroCpENST8AVGxTe2oRK
BIWU7TU8dac802cbaZLKYWhbwFQvwMCKUyneHEkLBZHLQ/u1UehLzrqsPkC9EG3i
7yGEHBwId7bovxtqPX2yVHkiA57/GmAasUiiT6XL1Rm112KQgJYBGz3qLHhIg37S
mQrxCRajos+R8GFHJ645gD/sNwzaTS5QuO8Wbyl6kZAnfeUjupqQsfbRRPi0cydf
zVoRX0Hwixl/PVJrKLCr9/QGcJ13fpHc6QtwY725XVOX3rfja8kPdtlgKHz8C4/P
59MvKzCeeqENkELEo2ktc+JTe5evV0BAdQD2UZz6vej2CkXQ+17qfnruzRYXZYZx
QvVAB3FhyA72wmCnCFXR/uq5z3CrqQ2aQHOF5pbx8uynxmz/O1exn0QlSY+LYjOq
CV6HD2Jwhs3zXwuwAyHD8ktVfSGfzgtCiPnAUjTTbZUHwP6yC++pAZ9cJ5POwyr7
ORF5pXpUefbSGT7XhL4yWq1D1xTEE7X6IqahXoQbxdeIv8rWVispIDM5HI01WRaW
6TyqqPbS4BlFUmlAqmOkfa/Pz8WSDqpCETI14GN0n7sNB8LV0xaudlp8Txl7iOVa
9Mk+E4pEEXZ51wnEAdIz57kWA+VoVmfQlAA92PMV1tR/r2RNeoPpVPcC1APLgEEi
KzqDJIJcqEds8ZABEd08Y/Q5SPRJbu+RejuK2+bYZc++h/0PSGEdAjjKZZfmZPNm
lqx69h+hDzWIYz5dYAs2RxjOo3W0yXdJDDLsnpOJ8rrnG8mXtFQiz3H+If7OWJKI
KMT+BM6zzCamomFMx9EELUPx5kENZv13/GmaQ7ZRxCwIRv0PeOdwIYUUL7EvChj0
tDHyDYtWRnKCbwoYa9IjdezSrBLUH3ThAw6+s/gb1Pnpa5LvCRa3L5iIdYlAyna0
9cdBZlCjutmBkuXZ+9exCXTfDupFzUIaaQdaxXBbLWXmMqYtXpE1e5FQUFx9vPKW
XkHtOp9bHWCXLdsBmOacM2ytZFk/TTcAQ3ugQJy+MxHzACk6aYOA5VkKTHJgOXM4
wAwXxzafMMK7BCI85yvLSkHssW3KE5m4lH1H7gI6oVqttzclfYeccM5H50+v6w/3
9aCP6sXGZOnPJ6yTWhBPKP3vtZ4HeuVxGWw9fefHj99HD/ng5IjRv9vPyx0WFQcH
UbsV2tAcQ93ns4FJNDy8vmyW21DH8ocyCJk0G2evxmxrLpqcXsoquRz4af0HKx8l
oYwWcxHS0tFXHk/EeOLqEosoJL2B+LrozCaxG+TqViJ7S+C5OELq96uqHD7oESmx
jCCVMjju6BNHdp8nL4TlmLCh5ylCH14LYQcfnX5FsrK+Wn1yAnMfsXn2buNI0K6l
`protect END_PROTECTED
