`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QaNR9TYrHDYjUEVoiRnLtVUnuhdPD3oabYlWn7S+iSPX+QRIXTnQBmwVNFZJPJ2u
6+9tklaLDlxFOxd0extcIbNHy0ZeKuO4cpxJXxdLnnz9mRynlf+ydB3uBc03GbZ8
BELwdiebhlYVqrj5MYfscpfohWfB70mQIaWOoU+c1wt62c7Ni4wsL+uUxUxq/7iD
sSILRoNwT2Fq7D69lS+s6A==
`protect END_PROTECTED
