`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZWC4V9iGGLUE8VxyHROljFdBqXyvyCkCJ5jfaNtESCv4rhBjgls+5r2NlY3ffOY
747Bzu5rDW2eMDAgtVxY8LNqk1PZaKr3FWur/lv5oeOkTgNSurWRqm5SB7dms0pK
ZVDCeRVpcFndbX8vlI79BZjmnhVrMuGhkL5ss6SaPjt9p/VWEp2dOWO6FZjVK9wN
7NnPC+5/jKxibDEGttg6rkK40ODZt7ebS5F0zGmyK4TF4BpVRv5yWOO2zaQr0TfE
DaF9yzi5XyWPNQOhR9aWxliqBwrkA1rC32gW/GSL1+WiCnap9W9cikkgzvjCgvGa
ePxf0FJBb7H95vBKbE5Ep+POIM0IHyhgPRyQTQT3JOLfnqNwzamTV1rxl5g1JoP2
01UuooQelcGcWhfPK6CKMxxMbG4Oh0dRTDGZ6NIBxu5Djm5s+Ma1byRwcaRosrT1
sHMADFC4ckhJ46Xr3jHZ0cDFFcW/lgqSDyQbn6GkyBU+mOTjXf2Vdjv8Md5hb7BP
jg5e4+zoqkHqzhLxl17qewzJe+/vqK7vZTvTY9zGuzLnpzXRF2DbzQSnu15BdkMJ
b/cAlgaq+5H8UXgo+pUxnoee3SK9maSz1KAD+ayObPd3wHgHgFMXUNqM4g2qi4Sx
`protect END_PROTECTED
