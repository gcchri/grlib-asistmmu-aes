`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YDhGIy5u9+4OFSRNXDxy4ty1uwU9AXCde9IneRZ29o3IKt60ie2qzWy4xQI8p1i
LC32wdibGtJ4iADRfehd45EtuU1xVYEJnGtLi82axRecPQGLgYcKgacsZjaOqo1q
BXSPGH8/ukvYkXv86TpcpG9aXlRWyG9KvNJJx3CoclAy1LBEpN0beW6DK80sfqdE
c9IqPW+/18HFPuiGr3yWamnDP/kt5U/4NsV+tuNX5a6ebHjGo8GGj38Si41+m3uo
3GdYmOICySXdVVQWhs/FNcPxj3jDfLXMeTREUFINxlLjjzGqkUz7zYTu7TNSipKt
`protect END_PROTECTED
