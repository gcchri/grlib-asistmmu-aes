`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
20k/7ZeQD8WTQvuVgNxn1HFXS0fNP8t4V6CzZ2X80qvKFdaBR39+D446MN6NUFEw
aFftEfIn1aoX1xK8uB1+0W4qP2lEMIw/xrKuUAl6ntLuGMVJMgu04dvAgIcRy1em
/JUZK4VRxNi0rr9TzU+Lo3Vswyy6O0tebEtC/wS+9GyjMohpDR7tF23waw+geOc4
28KQ8eQye1dj8qzvrnB2Tvh3wsniRYdOk3i+ElqtLmx2oIe0jPDoq3d/EuNUipof
knUfjfKCg5uZ9GtFcFHuskr/qkr6Ii6hSPH0ZzuKmgLCyG5c2sVWbxADlWkl/Nw+
7if7j/Kz12c9DBCYgf01S6g/2qFW71z8SGaAMhmwr8/GQWa30BbndHkv3TYSJfSl
sjbE9+5iSLhPv6a3qeXL2EySkEofEaLcYs2EzC0SQfZunhz1nUWJsibxETWbxaCP
/L9zDJp0nMG0ZeTK4fWxJmnKdTGlCFWKBV2bHrrVCWM=
`protect END_PROTECTED
