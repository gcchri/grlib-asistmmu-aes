`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5ATIgXk6+vbhlRfh204HQImMNI+G+1kJ9+hffPA/SGzB6l0WCSRvNVTRnS6ofah
tqE3cPJ15iCykAfC0CndRqH/y5C5ozWCYbvObqOB8zgSopqzmPltmkk7NrWnRrcf
bnQN5eD2Ena2xMAa6Gj4brFYRc3cyjhQ1hCp+ZvfZamVG4rmSWtseDTMD5rRkvTC
5asT5MRXZUpImfrkUlDjnRv/ioFJuj1V9vh7im2tTdA65I1QRwDmSpVbgs/ExBX5
qBS90VjvNO+DC9ab7HBjHuHJMDrKUrjV6P+JJZ7BfwFDudvwyttsr8UPo6jVRMma
HxVwDctJlSNUmWU9ZFfu2A==
`protect END_PROTECTED
