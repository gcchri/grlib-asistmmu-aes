`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7uHwxs+aj3wTX+Rh23H0+5lzFRws9hNQBstChO0gxNTQloEa70UHtpKKFks5uNR
7+Pgpxwr+9E/lfE/V21KboEA26bA36DYumftWu0a/21/AUz8aEmq3SyEg4SB4Dsb
sqlWcjQmdF+FQZzNykzLi4xjE07wqGpbC9qBW+8pJJQiQkdTr3hvHEpOKwz5XkMf
cvOpqq6n8OABt/h/A6mUI+blECmgNaVOpgUwSrBbuoULJRP2YyLWjWqtw8kZp/kJ
vCfZGjifpHEPf7EryWkgZ9dByU6E0sLaiPlB6JB7gsIvcFCfvFvfcDVF/So/NESB
g/L4ZGlJfp56vEaWOGAptD9TGI6O1+qGFH4e6KxcoK0vam2CPCQx803RaWuhKOvj
VPJiKDiFxsS7FJr8C4E8vWsYwlB32FAG13sgB4p0FW9z38UZMEnglLTd8Ceb7NCQ
1LdnntaGFhSKYzgDl6Dj4WKrQMZ5sBc0nSx1/mIYkfrJKyG2Ndl0o1oxMqhxsFRO
eLMkxbRJ0tOcK59ybgv1XlM0uWMoeOwg4G4GowIfo2yHkmr8KKqqMOTPzwmVrmLp
WHx5I2vczz0UNZr1hwvoRJxUDk0V/oHleJkPwaIntFZqbkyB6kcsocjs+rTWqofY
I96NynLpilXoJ/YGGj1nGuTjnukPku1PQM6IiaRR2NEfBs6GMbuE0UwVsJNa+HsT
SAvywusk22Qsq4lO/xajCRMWRNpl/qlYWxycZHIrNaL/cq2kaTNn9Yo03uMMN6DF
siDv+EfM0RnhvDhsl1nNEEPMD1sKIjEiP/lMzDZ87aNKqsPJhgZFwkMIE6d/xwMF
tm4eK5Kbf9mu8gCa4mkz6VgpLjlyL4cNlmSUhVrS+Dsgja4hgwDKA6iUZ2C/QG4a
1Q5eEg/HoCIXZCR3+M8dg7aYuFpjWA4f1WnAgU+j39g9mmHM+jkBzZmb8B9gbj+F
UeAySbNWehfm52C+0xvQLUx64KdoR+GRjm4y4z4Yu5otvofDg3tYelHWFg6QbWGz
dKgQKRpoHiDIUdBBuuPxjV6p6WVsD7gTn9GJ/5LJdNRDZlDvnR0SigpOnG9BFMwi
lBYbfAd4I/PT1X5xn3fWV0vkDEJAF5AOEUmQDbmsgpf44q+PLl5taOewywv73zTm
7zDhEin04ravqqCifGyvEYjBuzu6UHHS5sQwOWrZcSd/3hhMYRBptZsqNb4ElE99
uByYi7vtIf5J5flleoTKV8HtUjC1emtl+Pp0NQ6gsDLIXjN24Wqz33iC6FR7xLNy
xDHY80EeIi3Nm8yWFX8mPaz6/9SSGXz0fxYPI24sXsd7Ig8OJCko+xMmlZZysCO0
Dj3spEbQJTZd/N6WctljVS6nwpNYQX8DuCnvFuFMJQViQevCU6ovlMbxKTeovZqu
BnuqWHkRRYX7ny7+9FubmG+oHvmnB0J2c3Y7HU36RDoRpvESY3bYB2MhjyzzHldU
aEUMDnXcMNFSzjXNJr8qw1nSBr20hb8Q7y/IALiPUYr30PVM/7FXdrNCsFS/40VO
eNFWTZ4rXIpkpVefh3vNAKebcT6/3GOuARp5/e10/vRkzoewq88Zzl9+WXiqiFv/
3tVJefit/t+wjbY+TUnEf5XFTiOHLacRXMeRe1leqX88zhHOWdtaKukjdKJ6646T
Uh9INdXDkI18ya2zMElB8ZyK8LrcG5MIsDOaRyiFVVAva6EN8Nrl+zON5Algn3h0
2erVgkRd692tCUDC2GmY7u6KOf+VxYRIr5ErUTbaEvQXiTvv8UqRZANCG2DNNeTE
SqQMMPMzbUn3tgRpOwQVbyLDAiI5yQghszxYAKhyP+DAMqqzcpE+05MOxpf1xf1O
vhhA4y2uqFbVYszq/F/Keu6Wn+gR/GZ8HSjLG1eBKiSxdEaP1PHSbmms3hT88tOF
+r/oplInizMWKSGwZjZtjnwi7Kl+9iItrqNfImXe/D3YkpDc//fRfjtY7YF61tb/
siba/Wol1d9wVxuE6RJFnUaM7AmN9LO8Yh1LeFEhXo9z5daAZaDH69UpPDxviEnK
/O8bVe6DOjfhHJefsY5AW4Cxwj6t82pYfRC7jOfdk5mKIvvqlWGt/Yh5AgOz/y+/
AMD9sS7GHm7Ap4hZ5adrEIT7Av/jPTcZG1d4RxxrmM/z75EzZUTUyYAU6xpr9ONE
YmHguFDbFeVrzv78sSRzyQJ/xWZCTLCfR+Jji7G8zcGgk/MxWz2U3+hYEXpEfBsW
4ZGsJpNX+FFgX3LDJ1sH1IY0CDKSpJ3yel1kpSSGx2cMXo+QUzIGlnjzYqZMO8zY
0pul4bh05qkg3Yo89DUVFqUuHJ+RaXbzvFv7EwfGOzAI3DA8C8o55j0uXV6extSM
j0zNrqdK74H/0qurzus1CqUfm/2ZO3dZTnikMbkf7ScNuJPCbApm2TYX52+pjJ+i
oCGLMFXvJjZNryFsxBSJrKMf6H6xyzeQXsLnZbfFXA8Fns2X2uYOVdSggXJF+fuV
Q578vao817E4yRxaxQK69XFOXWciQJh/3U9fJzqQxizH9TPsBBBspYJeSh4g0H6K
CJFVGdZe57KsBDA2q6tW/Z4SJOyzjBiAYnMeavaudZWMILF4pabLS8iBDPVW/s5H
uk8611fuFyDJzVzErWp45J3WWKR25aJ2Yliowug1qv6+oqjIRHrHvuNliFeSMbp7
33MdHgrmB9kRy/jS514UyZb97YlmNeijkGHawNmhKhdkgTJ3Ko+P0uAXtDH6UTyt
NNkzXf7YhLdGLN6h5AvNZIl//tWFHRvcWBinhuzD8S95ARN8jQVJXgO/dKiXkXXR
//FHYy9aPmfmIN422a2csqSsVxzLu0Wg+/CQAR2/93yQLpKrzp5m7V5CaN9BrbXv
V/8FEf7O2Ta2Lr6T1BZk+Av4Vek+wE5lHIH4G0Kfcxgi+zFY8erfxU9o7ONaQFRE
zEXGrnHVaO2y3y4WAcS9gEgPhsauTeBnJqFIIFiyvmd7ZQKOPMilo0OcIvwYqh6I
bH54onPWz1EO/hfTyM+571PldXjDGvb0dW08buYfPdkGbl6POXIezw8VWRi3kaDp
/Q0DQ4wZ/COYKKkLdXd2rW5f1frAsyP7JwtUKmbPp6hUzBJjPlbxuAsRHS+HBsCR
5oXdv+GRRG5jE+DhzL1lrddBVfNmljcAqYka0oHeUPXCsuGv57/LVxYWg7UNaqs8
DFUMK40Hiplcs/4id2XsNwHGI7FW4kbxxi+6mYj9kB9KLQuC4C+HWx9YRTmDY8qs
momZdyKosdN7X/z5PIL6uw==
`protect END_PROTECTED
