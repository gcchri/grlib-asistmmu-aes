`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QYnxtc4cy6hDDe9hzV9l3k8MPzzKZ1gk1SxrJRzJZc+hrUkFY97gKZYrCsSxLHys
7xURnjjgC+94YII+O4W5J5T0vCLmqwU2zutUCA/ypiJZ0J34rMM/ftbue2qn4VvF
Y7GD+M85bYqxG9nt5vz0SlEwqVQNS4uJN5BLyaVU8pOvvlyOJe3bKH7wFcbNKKs1
bl5hJTd2pUVaYC+dYwsdYhM3nJsj52Mz++xNS5MOvWb74wEpxo9cjy2UqbrOB+xJ
7cfClHky+/0Gxh7rmowrwYb2oJj0oXfbNjFo85LUgDcTPb7pFted0rX5+ubf+5Ff
SGzUn/w/pEftTFx2PYqq8S/pzCs6jSjV/tgGR27I5rX81w9WnvLLOG4cVY9HhSiX
YBvFzEGt35iw06JSYt2hReuc+Z/6Y0srTX8icz6QA7h+7Ex7ajyc6IS1c8/N4IIt
sdO00oafprCgRyaaY0QmvZKTh/PG+meZ25b3pkMZZiIlK6QkdffJ7k3C9kngcpzB
C2J4ulCuQAsDZN6Zo5mRtbt/OxfZ5XUYopWX4gf6/oij9nFcAbc44i7uenlMsVeU
Cm3M4jCzpmgS1INjghDRNg==
`protect END_PROTECTED
