`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSBEe+CsZcXn0cwscQeG5TEv3zCzEfiIBramoIDA+7aNGxLqbppmE/+0IU/IVudd
xdDVQ0DmAXCb6u7+vEYuxN3D0hDXN2RyjXbxPWziCy+d+jC5WeIWiVqKKbJCS6ed
fuiCj8vUiJa060wekx5lgbh2J3/+vvkBZTssabtgHTkSN3tALoAHvkNE3SDfMSAB
EwVQpiKhD8pndTYMMyfEPTl90u3+0/NUHNERCQZp8Guq1KLiW3Zklckam2Sr2EvY
ilwMzIXRtqUE99nHTLZqKz/EqUN6kiiY3eV4kLdtI9wxbJ13671Sl3sXc+P0tqY6
X7HD6aFKu8Me1fpAk2WAIIwJnUkgWi9EZoQnUXH7dzIPOroCejVIDEePr1D/rLkE
2opSWj8mdMwx2JiwSwqnigD8s20vI3HHq/MV03hfRZ6yLcTjsCgFepFBapZEt09V
cOUcrPHFZKuNEi7c3qYrdGHf9eNvx0Szs42lam1XdBZh1rSt68fu1dp1uKZcqAAa
u5qIjgIgo/hY3VlurVb+2Txbcbw1/9lET5nWIVP/pQNVfkbmlKPrVowQgDQW2AkV
Wl5VAQo9lqZ5ZEEYZbc9qyk3Aawn1gblbFBK0deM7Fm4DI8QC5p3Z+9sbphXuMQD
2yVClrvAK/eUI03V80X8T35QEfg5VTO57ql5AYBOeD2TBRNflpF1fjqp32FdM0FN
glVLKOF96fW0RrfKtD+HAz1uwjirRWoFrhO2rc/+VCdIbTbDAaLYyMCBkqgeImSa
XLude0C5HzglQLb0tR89Iwzl+iA3MFVyvm95xW9Udln5R+KdflSaZ4ylWtgI6BSD
8/P7i8uhLnNrKMS07lzbjfOHef7tFngZB3/sNNbnuPiVJoEc2u18P6Xe0ztpBx0I
amsThB2ibuq4sMlrMgavKAgumiNW/0XYKuj5qzE4sjhNdNgh2f4ne7r9rLEt5f88
rKPXTI73XjPNWd0akV9A+qSg/4+J9W5LZn8/LnWekCrIUYcqXPy6Hn2cijpcNLs+
eApSAqBWkw5HAFl9vClVVMAcPMNFVz2oqSQXOb8dSpOKAVjCLp1i+QihkkCdkkL3
g7Tx8YSlG7/oaLvf8IPaIckLAmywLbjZ6aL9wHZWU0hF3eSIqIP0qglQVaoPxo3H
av+VfEWCAUSB+yepmCiZdhOnkUjRz72jhXutfRFJqSJ0Ig9VU7muRx42INwMEx60
hrXjJmsYzmmZ2URS9ofduKev/QTUqobeZHVcdGot62OVaNP3cKqMQSXYx6qLvsmp
YLrm487H7XlSVs1GfA36wVVxYb8VsQFPi4kQSyh+t2rYPuSTs8q+R1Km1CcVYR20
k4a1rQhIZU6PPmlxjGcPlKvLPC9OnL8rC6PT/pDJtHeYmQkX9LImbDnX5PgSRl6M
HxmW1+4bBrYCZlo2VPkTVIxrD8pi8OvauzeUbf+JK/Jh2klpiDjj63qKOO/5cg7M
Td2DmOpEvFxFeUwtPmb5buG1o45EMrTWjTyjAw8IFr5N9hO2DFbnFfaGBNGnLzow
bhcRFZaUerPb3lggqtlLjBiB5dI8wLisq7VJBbU3ejeOC4aWnWG6qF0ebjWv8ykx
PBje/yKMSYGVUpRg5e/bFj3pg3K/7UDi/LKN7/aY/vVG0SC/1kTq/6oD2A31w5sV
fj13GBXUCSvuIsGSnoY3n8NjmljMdkyg7qPbAWZD/oelmDcIk8VCojfhvNJGP1e8
0Y0AVJGeHgAlo9oRoO8kJacU0sZdrZXkXqhzoj6kkgroHhSbc2w/N4nB8GX8u6EP
OcWuzKzC7kOXuu2ZXG0lzxGveWYW4PtuF5cHPA4QeFpkFsLWIcFzk2ZPMKwg+sZV
QRQBhO7Tuf0JdKYkIVtUa+yQY3AhRID6gcN16+V7DDBjuLYr8rAonPmiVStXRjhF
5gGMi83Bm3Q35REhDdOZfUx2imsINCl7vN8rHxVS/myFal3YfRnEVbQp7Ico7JbU
gdUwZqkT0A1Uo2uSekDsdZcrlLTuJG9bTRBNcfpQ/lc/ptzrRXoztWbhMafB2Djh
vpJm+ZLRY49uIOVDE//nQhLwEMkKLpFb+wepOCuB2wZm2e+l25ytS2S+uHU7xg1U
UKhmzutQmRRk01AqxuUuC3dulQmWuemwBrIWK/809feqBb/rgyJjc8XDV28MKOtD
l+fqAbQ0iMA9G8zhoriNMet9oRXHWhED8F5UY/WR1mHLILmob7lxPj9HQSBgrmp0
TrUSjRn7G5zPnHXRqRBUrtJUx5TBoZRSHCoMb+4aB1b31UiaczdScLbZILWFhAAp
/sbdqpixZXIvcWG/kqbVFmJ8kFqcgfGO4gUcJGNxcRquk1aUWA919xwbr7FzZ/6J
cEbE1LNaAqRvoJdv4QZPYSNvHe8GujVCX5wvpJJgV7A8x+S3bhG3Iq1DL1sQy8+8
jGZGoeVPEoJarMUXTd+3cBoqKkBzdhEbBnkxSOsuFUZpojazEqpKY2tvW0xwCvX+
v+ou7tQaCojFa/ErW61v+RJTuEFcw7yEjaIUpjgzFK1g0yQU+y8PdY29Ofrg7g9b
pJn78ywI+vCrR2fbf3CXacoItT38uIZjocvtIGPetE7HrROMlAMZqewpu74aDcqy
os6YhYbbPDKyuF7C2F8pqTSQs0zbkHMLgrcXt00KAfx+dpdIxvmJuF61tHuXp+zo
vfXqzgyCFjl7ZYhhKSCMGlquaYL4d4SnZeLpuivXH6b/V5kLiaiKIAlVLvx/0QJP
7eZu+CQoJWnGnnYwrWBa6YFLwh8PrtE9trL0nErlH11/09gm/UfoN/p1nmaBHL6u
I8WOsc+r8SAJ24T+nIghQ8isbw/V09r9n2jVUmizjEISzFewSKTnN3qEJrerS2J9
LeS55iLlUkV3pq6iNwgbjWwO9FWHRI35lr2XkNEbj4f+dZW6vzfkhNo74ifSx+xA
GXfq98wTtNukmiH5Jx2tHSw9JDcrjhYZYRNTo53wOR5ER1WwtPoD9yk8Usu+QpE0
EAiEjbxg6IDxRXam92/Gpcv/9BTwjbb3khxuwAOmELpIpKwUtkqUTpu5i0bojVwS
Ab8SSU6LnYP7h6SvOmJdpB+dCwSu3Wjq3gykSwdGukuCn5IMmjUBXkqss6iuQ0Cd
CTkPqZ9Dt9cew+p26akup7SXy+oWdS3lWZmE/mbwwlDP7XdNXXw3c5A5Gcadq3U0
t6BQFANiQWvVYfuy3i9di2epJHXGIRKGCI7w4CGcCaQa00uhaY1ZC9Lz9gL7o+Iu
joRMpbMdYBGn6EaIy72SKEj0jxQrEMTilQ1AiZ48SzrKl9/SYG6OPKcbt9agreBR
ZsxeirfuC5jT3/Pk+iQbAETJRcD0OdPR28N6WlWKzCFQmnrP0IhKZvo/Z5xDtXVZ
9RHzU2r+DVqVB5rpbDdtWxnlH9pM0loh6G0hxYmZlNsyWpyZrUnrO0cTCE+JjNK7
b1dTLIWizsrs2V6pVjTcPoH9J3oCEkJhfKgUagAOkHY=
`protect END_PROTECTED
