`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t0nrSBCQDFG67JjTak2mfoC2rtQBR+dbKwmn7sEDbElsLXH5x96Xy4y/12bgY031
DHAaWc7HfgVhnQDeGqfLsKr0pxM4gH8GHjoNlI/hkz4YTQm0daNLG6xXsFH5TJdN
MRQJR2rFdczZ/gqj81AaLFWrGTYSL4RPWGrybmCHxmyqmRZFWztscwyhkWzzYuK4
/wdHjmdODYi+hNTadvMbscZSJVm+2+H+zBu81b34/66nrIyNRyB/Xrx0NA2R3BIy
nMJ54WjpXQfqE+T7YbylZU/oyoqeo4mxc9uS3ybfHg0=
`protect END_PROTECTED
