`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7IglovgWqluMrAgzOuzhLmR30lcVkzcyRCGbjzY5EJCFhclgqWFP3NBn9z32s8Z2
LKvJCwlyUMe3L8oW/+VnX/YxYQ4zyzLtPp68OBPCdBpMDV8a57ZlNM+7ds8zdzYb
Srn8+jL7RuCLZwZ9bO3eFyun/X4ZhQOCBJ85BjTKF+mdeL8/h/zPJz0kYxXT5yMO
9tBT3pFrIdGR+x6NuwQRMw5vdF4jisgAkMmXPUB7RvffPNRGu4Qq7jY35MnJTB40
iHL+qlzsellTcGHbbCgJ697MYJ4WmSw2QmAl7lyZcml2oIW9rJSG9dXpMh/OgBLD
irHoqHVO4+Zh0OD4lKnN84jxMDHg+1t/MujKjYJyuQeaG4p9O/QLumWItgRZTJMw
7aPYI7zMeZzoa4MOVbQV7l2gTzDjdtAXGZMfACbYJ/7a4RzS+qdMfsJLRO4SPIW/
pc6fav6eLs+FGydME81WwcdtyyN5QtoFgKum+/FALLMSiBXDtgFVtFvtNKCCfXcD
Fx1bd496hGdZE7NWyVpk65KPR2Ga40m/MFO3WuCd4iQtlDAtCBZfyM0sOdir//Uc
fnGqP/WsUaLAVCGagQseDJIAxN7zHtxv/owfXTkoahjEnPHF4QWhp79YsGgswGTm
1NDk93LtoBqFUhBB80XFN5R2/2QQdpz7y2HMI6D3KVFFqE1VDMsIcToBHZqEYAb2
2hBzEKUYkk04lbsaQhs7sUEquUl95y+pAGkeqn0C54AEgwPzSTsGhsLq2w4nYOqP
trJJ3riJmY0qnkkzGqFfIVPaMqa4dA2reYyaNbooaxmKQ3ztagTdebp8MK3/vcEk
0YfJZscz02NGgLvO8ot+ZQ8B225b/T4PeoCPYnkZNbHJyK8O8VExyho3dhaCIxwq
6Dmkm4CsKvZSgO9asotg64WhEhF3t+SlI9XYqUgS2tIy0pNlHHQI9RsCaxB/JVeq
vjgFjeD7Ja79t54SqHE/VRKCmPDw1uSsKjBUc94hYAk2GM6rTOl5+GnDVcWn8MxQ
wxvxsm2xEAsBgX09+WVcTvxDXASd2VipQJqL7fvMwfy7llMWOY+l4JF69D6Ceai6
4jFXIo8+q316N48X14McYGzxNxaRt+BdrElogdojTHkiYcPU159rvpZWTMCKQkSg
`protect END_PROTECTED
