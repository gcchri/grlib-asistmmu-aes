`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1e43Le31yJWr0UNhql2o3U8mb88vUsKPjeD4C0ce6eCVvNLTHBxKR5MkIoVfAAx
E/fEhrzZC2VihtV8TSWb/Udg3ChRnCST5hV1w5qCVz5oH3xUSG+yRh9XMetfZis1
KOi4PyuYNeSMpqR9LtMvgySR1vEGP40tyG+xmt7T95zBWpI6Sow4f272WZyd8yDk
R/eM/DOf0m+0elAZQUWK/pFe750QBapgoXvJ1xl4E6LJ6GgxexNQKE4SnLPwIjQN
IURI00uNgmXxMWlzbpBSi+aghP6aKaeG2B8KONZOzHW3asvTaGBmfuaG0nvmdwD4
vCCjZDvkKkpAaegfGHBSuWPCXjjJ1/LFd42RuqnmU63uyUaoipUaJJ1egXFMZlUl
OHVsmel1GBxqc8ixL8/tDVphrXS0p+WVPKR76wQv3MVJhIExP55Ftpfuo0WU2/+e
sngWQeZZDK3Y6dXUxLWhB0bp3BW9+I5HZ3qQnCxxxRU34C3e1HPZtIsx4Z6M0rLo
`protect END_PROTECTED
