`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+Idr+VMKjf7w2BiehsqtKio1KlAHicqBMbMhX5dfJwy8LoXlawKCb9I3P2trpS1
DmJ9+grjsCcg6tEJq2gUkU3NwS0bt/1R3RyRjJXMLYkogvDsRoOtEQLfBSumOE2I
WdrLIQFn2BLgkGpLp8tttOXt8oKDI3OBU51fGFOTpnh9fmL3xBhfUI6afOZNuM99
A5pxNnu9K+0f/UYOjQqTUptlk8nLDBsRWV9ZZx8rR2x9bzeScjc0hUPibLsShJGp
7pNVKSiyT1dtSfOEUFzBPos5zj+0/8lM5B6uOPWJzJU91c+lY0AbMO/yio7qF8z/
Y4rnhyGICr88r6CXvB+3Jp691lihbRrWHtbI8mdHuHc8b7/AsG+rY54dh+Rc7j9O
OqJJOG1Z55wgh5In4tK53tU7I2fhUnn31Xpo8qBZwifyuuJnvfaR0aWC6T7LImpS
IY+PeEi4NUKh61TtkaD0bSoErvPtKPoCrIfNa3Ss+TUlkKYAYcRFG581DS/HF7V0
XmErndQoKHSGcDfkTJadRD9c/qqLCpcyrL6+eZ/FOiR0126ewK48oKsNeUF38RJQ
GooOKc4xjxtKuIlNP7xGdcMtv6eWNkjshOLAObzBvXaq8Lf3TKwKUrkAWP9hfOl/
yE6KkIXX2+0fHxjLiL32XfMTFlk1YR4RWrITijvHDfmHGsleF2Qv2q7tmhIOtzMd
pxuzv+FX1U0cv0+6IvBPi4lLlvZbbJSEepfS9G1znTt4W3QUGUp9LrNJfZ/PODz2
Br2YCa1Inn8gpOoIy3JclO6nXGK/vsGeUnNQB7OJs0Ws9/i5i0r1fLBs7pNIZCo0
E0U6UeaRNwq5MQql8OkNepp3Jpa0XTna8195ODacPSRJlfX51w7Fn1uZWStV3zm4
51mimumYGQdZb+depJ3gbmmHACKnkiVINBJfvUUsSSnqKbo6gDbPhX1j8kKpbh3R
xYEdwoJeIwF71pFPci8pVHx/qua+2K488KdwPyx2C3eiJ/DF0VlD9mbccjsw8ge+
6XkwcaudkNc2Tn2EcI6Mpj4YYb8lH0x6mNE9ZRha1OjlS0SpgWVZoufbjRP/WSFB
ra4aj9phWd6iHj8H9NaC1hkf/zhxq4ycNp2hCBRvY4jwd2HcHdSYQfeldM0M83sz
`protect END_PROTECTED
