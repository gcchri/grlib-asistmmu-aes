`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/A/C3LIFdO2/rmrixo4kSORX7+MMh3gnyugo2K7YJ9u7j4W5mDGSB4uQ5WoD9ew
1k95zfxopJV3faWW6xZoy3KHgqsxf2RXShMGaayA9hXI4sM4f02QNXqTKRSnQnJX
+Omp1731b4v4A+THFnDCr0NER4FxTSfiyHZd+Inu9RoTxFL8abSY1YqiqWsJ5+L1
alzHVVF29j+kgWk9XPwF2A6O+69NZOfarmUpS4MYEhcXXT4bxpil/ViBf/hx3txs
5s9LaM+yknnB5NoraQjMH0IS7CmoPS8IMbiW8oFenju+USSViB8H/S5zq7NyUzyh
NRjh22F0ER3cuO9VJDqhCERQo3j+YwYHxMQmPiwBZRR+qJBHGbtP6rNUyah39o2z
KOFQbNbroaovXvHWnTa+i12y7vpOSk46G+/24nnJdfyLWvLSseQzURuy7hKNtdBW
m5tyapBwzdKANyO9ojTmTgTwFezL6TmSvH0CoRNHqZHE1bEIgKDBp5kA6didLtur
75eUrll6PTFEQSjV2H/hRPH69HWAaN/sDAEQTMeLg5fmJH2VkU3O9EzBPvKMYmKe
`protect END_PROTECTED
