`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocmkZZvcKUY3RBqYCB+ghXoJ0UX1Ke7buibq01CA8bdIvo2pGUxoO02lvClT/fyg
kmLR3G0ZHPvyh+lCEAP/y8gXTuPGlU2t8WXMEzLUw+lyfrXrfVJFSd+vmWdzG4P7
sQq5+LtpPnK34SDaQSvCBGZoIhT2W1AZsxFOW+Eq5K4atrJiag4vb/oao5GW+3ki
nkifPiABnxoEOAk0SQwmXtB8N7k/FKf9KDm1xfC+ycb8KcXkEMC0ymWqU+RlCWmj
uuXWLf0DiuA6cph+/1TELat6eFIceqXX5UoamsKfdK+FXbh6tdtmGp8Kx06aaCjE
/kUwoRqdTFtHHI3J80HwxJJ8BzFtt/kqDtamRiPfhX5tGCHKTobEOp9GYS/lGCDc
yMw3JyOW26SvWmY4sVdKlz+dbN6linccvJgYdjFM1t08UObXYP7ANUr1LGkPH5bl
g22OXOJPIZ8k08QT2A0uJ7EHLlHYkaoVihKkSdxkhI4eW9Y0oAUB3NXXJ/3h3Y1e
I8wUQahJPAOIAdyZlMQvktJz6qgUSBpRfErpUZwWdmo6dOop6FrNwTGXYH2PThI2
gEQpBlWifpUc4OutJaH011POM1+gSVbT4gxx1msgJrMST6gN6AkEdWHXJ+CARWQ3
Z5DBDLIQ7K72gDW3ys1mJfRSILuh7i0ZYMJaZo/+prTYeSp3aM2yimOr3Bj3KKzY
NfhaQIxoC5KMJHyQat0wnH1fMIUrtc7IUTvKavkHmdmO+QGiH+58dCY95S9Nf3Fn
O5UERrnUsrk1qpjP2C8XxlHM8Eh8uJerKIdkvpSt8RkewW9zrC7xwXshj4hlxAek
+pm7GQTiNlU1WcZrJCC2chxpg6Pqk1vQB5Yx5Vs4T8OZ4kkvKIAgPtnn7kowX4zP
ensCl6yHtl1mlXWsStqf9drsb+4hPjV0cViW8Kjureche0NE12yh4a+4QIWwy+aQ
vX658I3PAa9rGGaEhngYg2ot9F9O4/Voeu6rnC5GMhA8oFf7IKKIIWgInJWGKwtD
Vh8CH0z5xXiCRvVGTAVP4uKHTUP1x1NBR8qppTDNoYzL8IQEgW4Dbp1gwhYH2X3g
8/M49rydKYDBwDFHSxTuTAbHFm2wLUXZtkC/PxrSdYbU1HXLE1tfb+npLrqeMUj8
ZU3tjGnAq+EjZqhYfKaNmSJLxhqLOUtURj6ugNVPgKFNiGIJVjIpz0OOShgCS9kB
i3vLVl0bOrSU6ig5AmwnS3xgQnoy76iJacBZJicg2wAV3fJBZ1lRBsfKcrDZo0Z6
RJUA89mewd71r9yMf5cHqUQHf/bnsGeQM9KQjv3QG4tuQXeVjQ3dsgYoGAQadJgG
lgM3V/ed3Smvvv8G1HwJFQ==
`protect END_PROTECTED
