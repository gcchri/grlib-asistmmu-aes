`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+6sXvH/+28eumb8yY0iCiTHjxJ0XPxDpZXCwjIj8h2YjJf6CAYpp3/Js0BelWhM8
/qAU2uGt6FQMf7aWk3dXZzJtUbBSSeqlhvYOYVZIwEtcu6XnWwAg6ssI1OO2CJj6
B6O9c6BT+OKbrMqKyqbS/iHh3zQtM/HdKx2AT8MGmoyCbCfuB4jmcbMomUNpqUrJ
rrvQZM0yknkM+yJiw6v3TBHM/Wq9hhtanjers9q7zdmmRLfnRwKzKXQ+o5y+aYPZ
tKl2OzGkva0H4XQoi4ehAJC1jZzbWJT7N2FVNfsDupn7Evz5lvCwGgWtXDIcZoRR
epe+tdXuZPB7XHSNClreFauv2QgR8Uv43FRrjxW/kEJ37myXlpykDt0t4zRDIFcs
Putqh1seGTjcM1mfKaLvQKEles7GOKfb55JXQgFDCK6/DumR8THZfeeuoCWNH3yf
V/3+f6atHR4FEXVD9FUHx0LfueVVXV20j9CERHsQRmM2iHPIbq12j2foAJO+LTs2
DtL8S5Jjf6MvpnmCQczr8zLQExf/Jz47mlsPhf9/5RIeYTtxTBnWGk9CDlnXp6mB
0N5Ga/1GXCEddpxVpi7TnBJ8h0955Yp6UTmOq9AusFB4OKLqKCLMKtNj2tjviFTV
/ib54av+gKdlxU+Eq+4yLF17At9jxDdWf3Lb0Cf8/fsgZwHnSKMHisdkrhJvgzwH
k20DL5TNxp8UmzIDazp7q8RplpONskH0CxDTh/+aqTjySDCgIEowyFqLomeoBlTR
F2JE+ytH30jwI0ldhrux1VUPwCT2chK7+VB42ouIdJlscIxxSkgO4J9bNYiEWcmh
vm6gKBMgKO6bE++Y6Q2tXlv0t6OyZcRr6b/c6dodLgpxh+R+KXUVS+AHHeBJFf3M
jDlAh3O1kHBNl4O+CpzxIA0rAzdY5K8B38gA+kvIOBQr6Wqbvnam9Gazy3LimOuQ
lxGdiBBWGgCt2ke4er4wISh3MRxBNTS4lrWVFqmodplD1PrWAT4ZyTO9a+0Q7qmD
9RC24mcX97VrNwMJR5JJjaNx7YvACb+wLvQbiEx5gFjDaadQ2Mq2KZFAsWP1tKS2
BG5GVxuLthq/EVtklL0P0uVH2N78NVMcar3J4twdtzAOUuhVJF3i+5MpbdeUofhe
8Q7CWHa3fCNOoAYS+KS81Xaw5RCjruwF3qtY6lY4MOIVRdTbNnDKRqTjFXUMCMHa
Yf/cytHOaAyhpQAJo4XMJVA/hPdIUyihKqcBJTcOrcT4Ie8JDjrJ5vu4lwgbq+cJ
N/b0C17MSZlw20ceTJH8aGdlVRf0qxJWfwPdjOLE/W0gPOO70H5IdQQoqHpkk7eM
4qPGccnxcGa9MDNQgOUpOL+HxiCtA/GOu0ufkVgkPmRQl9vMQJUtZEUX/aqkBrKO
Nk3sboGk8FlrD2fEi2CrD15oSv/bTSqyKHlgQHcCPLS3Tkk1BaWTcHP0NGw2aD8H
B2E5us1T8fqD0xpeyx+lUY2XYqtvpAKG/4DTSFLAliANYEuavQkZN7LnGeh3Uac4
ASBJZYCp0RIgWhsiI6L9pkzGNn+LDmtClOG/1CESi5ojeOwSgbJ1ILOU7mM8PcNL
DQtR2bJEi2JrBDtMjpZZIwjtEX/xP96QVgHTWkOXWjYvuRTpSrFGp2UP/rdg+dE3
oBHmORrKZEEhmSbdXRJfkua2KnM1Ub8Exta7geRO6WpL7HSsc3jKbZDVxQEyfpkW
iXoLsC0UGxs7OKC0kCJXhypVh03csXUkTVVAPtOGCLklmjOh4xHvt3Pl3tWoYCMC
JO/7BFFYPtJSHVku0DKKgu0Yi1uZsAEQGyhqZNJnxv+eHPWSkJu3AOYxwmOFSgsd
`protect END_PROTECTED
