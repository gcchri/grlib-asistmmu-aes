`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehIQutNl38Xa+bTlfgDeI3F4LL8e7WgaK7TUv9ynV9xjUM91BK9DsibBJS6jP2RQ
QqxOx1AAlmhuJdhrll8UaShXvBuT7x9Tnql6xpr0h6K3PQR4hKpOdlUF8HraFNur
xQ+dP6o367bVAwdHhBaoSigJWKOMggjUjI3GdTYR9kLrAnFm7GEJHQv0WQKgjb+V
v5FfaFfe1LMwzyxSmTNH/MfClI+Qjfyiml0QiMZk5BIe8r7F3Bgx82im9mce1MCt
pdsg9cDtKPGtVYdlwlq56w==
`protect END_PROTECTED
