`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zuTenyeQiIVsRmEYdlfnGbuVbxZov95wKBGCTVb61zG5rfOIEPLMgpjeREMhkptb
IKsjqj4AONM5LotMFgEh9FeE9+uuvIMZMNhyGWXL6wg1uWvGBSId1hYFL1ZOWJIf
cYTEuW5J7UwJX9sopsSWlXKRzYqtOIHITzEJownmt3b6rOMNLJ1SHVJBY80955SM
4x+2VhICWlaGEKpm1GSggzt+GbIOD6dNxnFF5OzzWGZodZatH4vY1hZCXwpP++M5
CzMi0vmG3XudEbTJf41nuGfvNry0BaTZlBFXJHA+C9WZk+vsLFbEAqaGp0WDCfbn
2E+yx+JE+JlR7/iLByJYAXsqwA+RNvacO0YJQk4/dk7+6QAopn6XPZdJzGzX+APc
tDD3Y86qkJ+FqXDJlLlaU0aKDlpzN5WBfF2qRKIrs/MmarsvVC/KAiSSORTgtvvz
TCHLS3U2U9Ab1b49gL2ZpYjggbcQ0VsPLEtYy2BPeecA0IKEZANiglioqaIHyr20
NGFPOf80we8luSeq3NuZUJttqEI5sssQ0PpcOu3aqKnDO8S626PmGL2uEmbqdWrU
wfxI6KF2gcxzvnb08Tjm2cNsPZ8Wb9uvf7IalTSdfN2xefhwe6ZRGpVwFvdqyoCy
qUoJDJK6wwf0wmkvlh4gEVnShJ8ngRZyWrXGnTtQu+gy0fGZxk+mptQ4ANQEEJkp
3j173rP5Uva23ZFJN9ckmN3bok9B/J5mZieb4Sc2ClW2oJSjzRt+Nxh1LgDt12kN
9joiXTnvgL+7qIpstIZ6jg==
`protect END_PROTECTED
