`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Citk1YsCDg6KuQkyKKoMcEdtDt8lLnIbMCt9hundADJtwKdxs7bB+BRFf97X4jP2
RhjYiVYF+7bSge7JMIwhhSGfBF/44PdlHuhPVLKLAzHdiMxld4805K67bHOgRt3r
U8pR7WIdheThKRsHlGJ2CMnXOZS9AI86Hc/AawTnQz2V0RNH9Oquzx8QefIbEcCQ
9L743PnBaPhpNJ3vefaWe+3qwyDdAR7fXX0etwuyuFTQM83zsMMoJ3RopVxucQ1o
HYtSP8+beetKoslIvU6JmftLgJqdhgE5UkpJGE4MvaHqjpIVIryNWIEp5tfZoygJ
GH6TPgboYFFsz2ySBiqzLlH+dr+GCFaXu6mTe97eKu3U+LjLG+2nBr6+dPlVDgtl
Unt6o9je92QPezPkouQ21XCH5YTyWBHoY+psjVhVpGEgYtI6wtFy7j5pMC/bhLHf
jVGOV06JNpk0r2DgK1/Qh7AyETQmLfUESWNgZxC468tHaXJcxxzuOg39nGleRzGC
pTx0E44oibfkso/stsLbLl5cJ9KJ8wlyudbfRDRSlzt++CgaCo9gSexMm1UY1Gur
MyhPF1MS6L3HRBTHapL39J6iC+xXFb0t8JDHHpMhqOyRSsgUiRNbFo/2w9jqDpfN
+ZaWs9pp54T0y53oqoh/JJyfUk1V1VLAtuXw9qNCdtECVhDihqnD8JwVK1ZhPRkx
K+MF2PdfsPKHdTo9yhlqxq4zxpRUuNP3wmzQGV+YbgwWX2SvFJtIhJwdSpFxAW8J
5hMTXJJ77zmrXD/6WmGLPDALMbno7dIPKSPBzXNyA40uBv6WiPZm7Dg5GTN6WiFO
RV8E9UYvth6lE48EDl3br//STTDt214hr/UvN1zHHIoOSj+xrie9j4kRah8mlo4w
tZIJeqfTfBbssTeLlnCmZloxRD3GAFTiEZc6VJLXlo93xO1jBMbzTNwoOWmI/Own
fmpAYUWdy/AiUp1pJW65myPw40bLW/E+LeSC5QKOTZsp2TiDoWo8lS62uzEV5qty
A1h3Y0CZVWOgGRBoXlDSCCoEPOYyOgYA2AbMrl2ak297s3CcIlUdculZ97F8WOAJ
5+ZZ0tGFaKrsbjMsoGoXm9SegecMeg4mIIe3HsxGvtFybrndOYj5Qobvh9LAvB7a
SngkFicxyUZKI4Znz0yqhQh4vyaHJw+bvWUSN9EonOVEKJQnPI7va8hp1kRPdF++
5nNh6lYJxbm76vRiD+rgoia7Q0j9NUXRvJBTvfX/syJsstF8tn4QwfwYEeK0IyHK
/WZmNXfC5iOj3b477VEsHkq9j4UDjqBhNvLFHiCTu2EHfnMmckWfDhWDqHC5SK2H
N2BZJ05y7PkNNCsc9qjgIJXzILYrrlN3TEpJ/oBnUfE4SawOclqfUpkOTIYZ7bjF
nsPyCta745svlQQbVwrZwxdkVSaLivGcmIYBrCwQ/A6RXNrizT+jiPvP3p62wm2o
TVoZRJ+9US2kptq+k74rexisSDt9JBv70s7COfvZ2bxzSuTiUPcThvPGT+A8d0Gm
3vbSJettvj7NHlRPz909FIzXLgMxRJBqlwvMJBod/FYzLpsePT2Bl/3acicfZb7z
bT+S8pzxTtHWyRNPS/luvxPYWhdR94WBecCnLyBAGtwSiagHAr/6hOy0ZVX1/h+Y
dlwMALe4ng4z+LrHHNaXDHztg4W5uCbApRPtleRQ0Z4Jwm5UW1M1FCv4cUMnM/zI
43mHmlNJ1InJkw9qALs/mzK52/rS+09ElWYMvyTep3r7AvTuSVcdicKCIpZ/f6rl
zBpFinSVGJAnb5+cgAFFqsEiX6tGPk8Y6QmjxksPJuDmoHTbgIv2wIMi3qMHy+t5
DVbhzLDl+HyMhrod5ljpnRWpk6f+136q282Fje74/ADrsPIn6kAmK2TNDdvaw6n6
zBViBGktWBAoc56quLvJWBY/60d5XIkZPZgdsfRhrrV3UAfaXcpZ3uiP9VY0JqHa
sixuVamu+sOSshTfgz6WmNC8r7FmSECYlpGwl6Ga8NtPEniOpRfD6zOqxpIyNaWv
M8o06HPmrYxTnLJ95i9dGlSftCMOr9NVE2WmzbR/cPeFnroAnb2l3yQwHvU1F9BQ
khUeD5DKmZdJ3NxikUZ5efQ2EdekVl8ZuzrLPETR6NAK6ZYBU4raNF191YKrsAxx
wgxEkiFmmnAiCtmlZoiI4w==
`protect END_PROTECTED
