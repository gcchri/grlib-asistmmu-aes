`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSbfvN6DZYu2naKF0+OFszqTdNXlQMbCFV57ClvfUKiEAj9iZg+spMJ3dHrpMxID
yMBsz8tI9nGGQ7PKivBC+7ORTnA1l3pI7RvoOrQfdU9GGhB2lAaNOw+gHTJGUjiG
R+K+mcSG580zojgTDZl86gU3vC7xaOoqG56++STeyny4vnrJP5OnzJyDoHhOMcqM
iDjnr/PwElLql3TWqxzH0JNRBvIC52+2y08iw6bRvS1ink9A1cqUP6hZmHC4euj/
nPwJIjDdw2yDpFb9fUjSQ2+ysnZat0KTtTTyp50IRCN9ml4funRjmqRD7UaEamYp
KMNfSh5RLpNx1x4GQIIrFyuwUh7JcJHVCUTnkbjF9t4cxzVFV4yKyN+xxyWDrcpL
IwkUv53ghdJ4rmNvEeMt7DG9XUVqKL/Wyu6a4m7+zA8=
`protect END_PROTECTED
