`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkV4vunrvj/ZR6mXhgHPpurBu9cZU7k5rnzCxchdTrktDPDbR8yhKWqvsVGAnADI
06jtn5WZMTRSn4P2lI3avLAEsIgBGbARqhAvnEHgG7iEeb++Yw39iml5UaUTw9CM
hPwrUiXCbb2/luqVRn0aGxrVy0Q7S8/PUWBDjJfCtNgGbRs/0Is9gOOpXN7XryQd
NiwgVW0R3BdqRMWwuBLNNpILVzvKmpSBfmdyhCy3Z/rzS5HghTJOhi30jXeqKj4d
b/SRNdbNI0rhfelEYve9yHKRxTozOY8hkzNQk3O/Pomg6b02YGhrzs+p0DAzPnp/
Qx2iRhSPsXLpJ433xyATiWUj8Q1NY+WTjW1tmK6+yRRfBNbPdVMEjmxUrKvoFLNG
`protect END_PROTECTED
