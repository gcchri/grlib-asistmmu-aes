`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yT11+p9O+5Hx8a6pYJe3wfo8FgUa7HQbiixWfR0VAkr9cNLCsx0AqIaTgQqjshhQ
f3hguH9MGM71cthyNzXlA441naIsEfPFAX9BIspTBm8lx1I4o8EC8w0wK+I2Nqmf
yuDzvHKtPCHKbozTQdeGyG7DWUi6FeneGZ9xz6yFJIzQIW2DY18BX7GEapj9pYGQ
6UWGgDkHcux9ZXW0MzYpODok2bnFA8OaazWgufhmRRWLvu1Oy7/T99HEsE4xB0Rh
x10UNb1tjv6j4/jdk1GY73sgpnQPCrizig6ukaYraa9rHFZCbyacd+5HpHk8wc03
bYYuEAPyYqVST01Hm9ANjwZsPkg2pIRrDnE0+XcKv1tgszc+e33EZMeGnrxe2PS0
/lxnQeCEGH/oQ5ONG3zPsa/uB0z1Vi8ULJuUryYX3DUBJ6RmBuqnqU2vzXMVdvIc
yYzMOZPwYGCkJz2CsBV6Y4LYrbF3GJa8czroQp0uLaanXMkfVuYe/5kDRXM2zvF3
2IsaWxNXfn2CVbcJ+J1wYsAipTcQk4wQAKBPu1b4VT1nlzMx4oJkWHZHW5OB57DJ
aSoFgQUsWG2F0/jJkJ7nlOe9BsBa7KE1hMVd3Vl78noaBbRsbs3ZLFdPY3UYCcSj
G2l5gC68VvUatMXzuz7cRWeaSJIohMKucJlPKSAiFnLPrcosW1N4JAS2aTJR1bQz
4u+K1+6aT/dhPanggVf8h/RbTsRCakyA8fPYtqYcIN5x/m2o/0IN88lv1Cjti3Mn
xg6II0jUSWMfQVzQZ1DmNtXcZVtPZ8SnD+AEEcHK2cIHfyRWAh52Pczz/6XuUqVh
mAptEGyAEv6sj4WtpWWmatrxJlGF+806m2FrwYlcCmwo5Oy5WLdO0ar55FjRtVSd
XJpDOgpeYLl1k34Kj9Zlu4hXDF0bbI2sNX9ioItkraiJFV2O3TJqshSfN8GkXN1M
Gl6WSzdbhuuMx35CSjzE3j2Ao8plUVoZTD5JA/SCYYrT6cD76f48QJRiZtTHHAYh
FtWBxbqCj1TJjI9QAEqyx1SUSeroobquJrjZP+RWOvvczzQ4E6Nar5bMAFlNzyAl
ozrOe0H+pe5Vwh8Dz057d1XrITdJuY3Cep1XxVkk5TudLYsYMqJK8d4otvNQqqOY
Cpfh9pu+7TLgE0s27ECQyFoD5SO/e2CRrO4s+ywpmiIvI/nY3zJ8jRB3kCyB698P
VQCGjQi0NBYedjFQv3mwjAJ+1rujp9qZPFoJChtaqi9+vR38fyThGeItZvT+9Iry
HHwPrX1TbSLFx+aq1/v9jBJEPrC9Xex/1sl6Knmjtb+pk6jZihmacm9DPhrYMjGh
BIsgCekyfEB620EHhjgSkWWN10GwV3tL3b/XXxSraNOvlLcfPcLuqpueSG2lQ6Wo
GHwmaN+Hnz1bMeNJZab+ohKNpbfhve2RjsbvfNd3ZRP3s8gqAvprQZxrCjur1d8T
xgcuE5sN6fELuojkk5Nu5AlJ5BfogFRcomh8T72xEzAleDUGXT1yzEigwoUaT6nS
yKUs3/aUXq1iR6n4d8ezl0QlqoY63e0+E2vnup5WlR1v5ifahZBw7WjDXPMkSTni
UNtLIQowijUV49b/RXv14vh6DpcIM0Uhm7XuF27mXoasDwbmOpiqEzLazc+SFsag
yARoXZKlpugkaGEWLdNUMG4G8gEdmQVjkOEfFWs6KSMOWRC5mQohjX02hLxevUS+
HnhlmCip3lJ/bVJIBZ0fdqD7PaluZ3YdfZQUGc08QP5u/uelFKFq4KHh5GHuxxwU
gHzFafgrBhMIeNgEFOO8JXyf/j1W25ptr3zIFvDXxzy1EToy7SJmffu6sm4gRdnv
B0FwC2IwySgOOqid2Y/TJ1DjFAKM+5FMSXlVwL3nMRFNnw6xAdBZnCd47DVCb8uv
SviHsVSIlPW9wia3A9rLX70IUj6B9mr2e7G90PascwRcvTgkqKMzZxgAhxuPvGmE
iV6H+WSBvi52d3HYNonXMSoVwVWfmpzC6vpMcdKMAv8x6pL/0ueoOFBg9cxGyB1q
jgOfT+EpaToxJY8q973B2syjfzcatmhcOCwQVQrxBQpnUTieXDLqSmsY6qtSczfO
mKshEfgAqQtEzLdQBslPrlWzRtMLdRxa6vXFMaaqg4eVCmHRZPZF4F8ueGJM+JHc
rgU+B0y62w29nlh1+OTGt+Jz7pLzmNtmVxluGXWGs9RKejwI1iEN/Zsy7kjEnBrr
v7zkhT4Q7NqVX15mmCUF9lhs7ZhoAl4K3oQ5PucLgaYGVWH+PAPQpJqqK6vw9g2e
+U2H6tT+DwDkURTFWdxMAF0Dk0dZeYSfJFAgx7EY2rUk0cB7XvmvZ1WCTQyQb0WY
r4ulm709CFF49AwM8pk3kKur3GCJsTeexiYELo1cF4LFZMhG9It71fmU1Q192azV
4tGSYyHCt7sPxILUIOHGn16s+9TfSFoR/aH3h6w45d0GJqOv7pGOXr+KWQFR9ZyA
ik5v7zaZry7gPFItpIB1oz4yNoxk+lW7ZJarRVVSvoisjlAVxMndLEzJpyQO52SI
FaqYQlqJkab4j3ce5rzffeblBo0eD/HBfnH2oxkazn8kHy4DBi7/x0f0jkqSnRyU
3MIHmKF99QkL7zxhIg3W57aPECpwFy/oRyB9XOdLDP4ZaDVOJZm/U4dC6Tx54gNd
932ckdgDXaWg+lPy3UmS1mJEMzErYR/k4r0g2GAxXWA0i+5Csb0/EE0PrNJT1qDy
TX7Zey6sONNDQcCQgZ7aw3TL8m4vKtNec8GgCn9+pA3srtMJfTRR1vbrt6i6SxKM
nT9K9ws0NFNC4FuOIWjI0Ie4NDmLoJ0g08xAxWQwCSJIDofqML/qmpI7FmKjkyXJ
WOXPUsyUgxuslRKVElYK23JuAMpdNIOTmKXGWW5Md8CpFSiXqeDu0KZs6i3FFb57
aijmKSgjXjyFVy2ZpuzyOAkFRGpQpUwpyFH6jTOrXPjV2YSJsToNj6M9C3Wtv9nM
F/X3rhcGr9ljHpCVRade4vzUik/YibP8W29rssUc/G8lTcBsY0SnegKF5DL5WUpF
8J+Dfow7+GPesOWfCBAhuRrnZskfvw43rDLX7ynTbnxVqqtQm5DK2x3elDmlFpU/
r+fKa9nkiSoyoVS0F6SyDYGpq2KoCV05LHGeDGafT+DutLpEDKXdG+dbLK5bqLSZ
nyqdZPjAeXo2tKfYoibRYpoWojRe0u3j3paq57DspdcMLQbjGIGVgrlIsgW7jWnd
XsEer1/uQeolHlK/BN4GaDTYbaNZTBzAKV4CXeTCIddXAGscMF8Yn0AgewiCDNoi
EEnZ6D7Yb79ZNX/VgdW+DKqolHN8vOHpIEzrvE/ULJmcVcZGTADmsf4w5CBWvoY5
1OwWBsjgdggeG2ps+ULNL2b6D4IVbE+FrqCHBCdr8Y26hACKuQGW19VBY+Oiu4oa
1VKv2nc01muAx8owBKJnNEH4VaofdcKx3woAKrXjCqA41ojRFN15D9Uzs9gi/2yn
TbS+Um2SpG4mEoK9ecfMxQQ+wqZ8Pw6q3oIFtC7Q7RLe4ruSxnL1/+uSC4WtCZV5
aY0lWoVSNDmSS0KEHV61lUgp96yuc5CNItrMeHXWTO+JKKKSHo45TEMOZYGx5tXu
ODbR+D9KdTiCED1fCUnnZZ/fqP1Kviy6dE6X7hbR4d7ABvyhHCzbiPP4+B96mE7z
rmr5OtI92sd/k/TG6dp/7PYa6V72dXuflLP4C3b1ThEotoG57A+12ooBfJKAVSc2
0Gx8XfxAi1KKLw/Kt6+Ee+9mSpMUViPCUq2OJMl6koR8tvutR3pG39bb6ZJjvxZN
vg2rEYcTB6jrV9D9NnY7kVFe79owJYAEbEpIosT04nAMFHz0+Phj0SSp7jQERu5E
DSPTo5rLLCuKmeqTvwGjJTZZ2UHPP4+aYjxOD8N2+xEhtGppqMvFd7rscD/Ki4mP
Y69zkjILCb44Xdj7HbZddGL8xY2oiVLz/Fm6pXlIrS1/l/fTRvFHFUTXYttWwq8v
lY9MSlVDdbk5UXRDqqexhxDRscK/77MMUtvWZzKQyf8YhzxLBtUCuDt1qBohbbkM
4L8qjwn2zIYvQPfd+1YfMMOursofVXAEl5uZtU1L0Oakxb0feNr6Mzcvi6hjd3BW
PWgbRBn3e8gmQ4qQ/M8Fq40MoS2MBHCo4tMRvfHP5wGsvdVq4QMHtLyICSUoCyvW
bPyOTI4P18cTEwY3Q4f2gzTNzRx9lK+YlkIh48L1YVqXJUFJ79lUhkn46OwYFufQ
cKE2EN4Cj43vRYkcjtPgl9I7CRsz99GGefXzZwARY9SJ0H1KB4xgbF5F5UoR/dES
s1wb0rFZWR08fOehuSU7SEcJq+XuoGUciLi3fGjicZVMlhGDODZMdRbHtWekAFR/
gEjBqWfannsWr9RZfJID/sfmpQQBqY+gmubnKy8CCyemI3T6otMhHmM9Dnh4EaGa
rGwpuDwF08xJ3tTEQeS/MbQ75ObraczkqvfXRhxEdDcK9zNplZxR1+xbWoHkvmIb
PJLMbDJGcErY0dIeUdi1KYjBqZY3v0Br7jWa4uLP/fWO7nk2ZBn30sjr9BmvXHfY
P0Eii7mx4jGmLsNjF2RJHyPgyCiqpmw7I0hqvld3bhg93ETe5LCzk82Lp4FYCd1r
nlLrAedZ+VlvoNkJyUVuiRCY2Yb4gS2p88zEENprCvGPiezhMPdHm+ZFHKctrNfb
qIukknoS7JTqFyJxA60oi007RHS3wvdvk35Toy0XVsi4/p0iWIH6LhE22zLFhr6x
uAbyK9l5ulWsvKgX7vQcdpeLwfJcrFzNAgX+L2Y5ZOmlr7xq/UaOzNsSmdVxfxqf
dyraK93vLHpM5LUvrGyHBe7h+oZEHjCegwphBnkSR6/2Nm4CKHKt/2rOhTVV7Sv+
gAxy/u2pgoaoGERduUxR2W4ZiIHNM/EAPKOqetlhH96HEswen7/dpgAfaialLtpv
oRhxGHREy3X8WmGVuPkO3EjHgYXgKbQt/THNYWSmgHydvOKLBX95QKipP5DbUb5F
obRYt6x5iKglpKrq+QwEdA==
`protect END_PROTECTED
