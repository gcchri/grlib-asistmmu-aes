`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qEvQIDFFbmLNJi6I/ydJ6fXfFf15neF8BU34F82aG4eo7tX7oromrscUIzkvQIVL
uqc2Q3TG/e54BeBvnCHoSs1q5OqnEpDxVajQeka8rLhybBn29iSNJ2MJ/VFuF7aZ
xIc/g+nc0nbBGlCvSrCiUD12F9W/T90E7tQQiExpoKvLzITOFSkmLByP7LH/f4EO
aFl9yVZwRO25VON9Qhr0OPkc4Z/RoitFwRaNbYpr9bZ6HCkrTC6z7bv/ur6mg3qO
0FyJFrIXjj7L3nd26LJQhA==
`protect END_PROTECTED
