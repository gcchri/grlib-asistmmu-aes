`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGpSOqpR1I24KTKA3z6iKkyXAJf6aMKterEucP/UHFr6vqK/dAyBMBh0G+CM/ABT
O6wZN/zyVIQfyug2ysur50WNFt+FACz4zta5Cx5zFCRR25WP/7MNneDzv15gFPf9
Hw757fSIOqurcj/PSRwzwaS7FIOpwpoq4JQS/93KNl+d5DvFsWiMNmD/gYGkZ3x/
e/DeD3A8T8EWzzAphjbB8p78tDARuEbAPDep2yAVp7Fx530JcqrZZVubRmPBLoVf
oYEEniSk7pzzETb4T5p6Jf2X3i/IqjdyVBoeSQc8E7RErtaViVUsX83+uMsqjTLc
6CG3FuXNdw7B/vuvNig9nxEEfKCsR83MHOBcMktFCWyjMqXwyO8dLBBCh68gVTED
W//zKwOjyZNmsG+MvvbAZw==
`protect END_PROTECTED
