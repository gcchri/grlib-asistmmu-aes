`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HG73JO5V7xxjG2lk8695bL9EMZK2GVJiqJQOq3QeNGx+PRgEoNmoj4OmTjC+076x
ixrtvyRIktn+baG9iy5W+lruw/9uUGqBcVzoIZor42O/Dp3/0PhYR4Mna1Mj9DF9
vc+1vDWraSwC3spKTVerDCwFPHTHqb3yq8ghHa1C9ACeNuu9F+snKa2oQyh8vZ8Q
yDLJAU/emG76FMCKFs6ghnA3iYjWoJ7/RWs/GiXPFJPHeUO5JCPY/2YnIxqr2haC
sGtHh0q+RZRq/A7+paQvIQOsTECGYBezOOWo65n5nytIeGl8yZRIrlmIQDnKmEid
6soLcOMhpLnim9XkCF3tUqQ2d/sYLTRwWPNgm2OGgNab8MBnngJ51vUmoNC3fm2q
ltvCYvRuC8aJIyyWylhXTwZE1lXz+EMkM7MB/D3c8j5JmX7k4JpxQ3Dkd3Pdl3ck
gSiK2dg5vurnc+M+tOGRTcONr/gGvNDilqA8ECbgjbujICJ+Ry8bv8f3UhCNd/VF
`protect END_PROTECTED
