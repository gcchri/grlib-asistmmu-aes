`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8pybwuMepiqwshVPhTa93OH97psaIlnZPUIZ6g3VYGmruxtrFZewORzmqc0Pay3J
jTKUMXjCV0tSPdIQ+0OZHvdI/IAFIuY0XYis/s7+/te23cEcpzVmwgE5rEb/me9V
zFtHlALKIoLUdusMNU78ZgIuB3VgLTfvaMyKqH2c0iTLE46uVVVavom4klXvFIwI
qoZh+V3uDiiS9Gh4QLpguwTWxL0OK4Jk2In5dH7nwFny4OkrSK0kWmEdhWrDpmrL
zVJQG2gU0q1heuS8z7DKk6tQxiKzNIa6wyCVtUFDr9T8Om3y1PVlQKh4owumG7AW
anGWqwEbeelvXBc25thw5KODLZe6hv9TtWL58vlr0G4x+uwBOjZoBzDdDYESsPJb
HF7KIKUOBs2t21lr4Q7S+pW/VTzQaat5S6aDaD+tmO+zaPO55V0OzHk1pfpNWolB
Djz0L2EXilHdKd4q+H5toSAL6kYZzNb6d869O83JE9VVbkloIX3c4u7CtOflKXJm
+iVEluDT+DuQHC6zdrMBhpQCxmH0V8pZC26lEHVNPL2UBxJGdoLO0Y40sL3EFZZn
GHNbye9H8fLhzhTakhQRLEQGgVjsY6L9cdIlH4ozuuKXnJvi6cwN9eLfOfdsyQTj
FaG8mbLtNtLm/DhgzjD//XMwYQDW+Dq/f624erVm4TLQa/F86ICjulY249st4C4P
/zVyDiViQhbhbfPwCYvV/2j0f6MByRTKIl5g7DViJI8fjr/U5bMetU6GTt74652t
0szsOE0eOsp0b9PqOnDSSg8EF9lNjkjmZB94I7CG/ucyYSuZZnTRTzCj91Goy31W
t7gv2LYHPonfCl+6iHZtEAePBpKEmK+xpAe/MV9aTBF4NOxtGYmPGj2ZgWoRp1Lk
BafmqVlxZB7wRjO5stoddhhdnQXcayFdoDvFcobOnveRMKX/n2awJ8RRAvXoohVv
0VknnMcxX0+mXL2PrncabpOGKLfUr6/20TwTa0lPkDb6AM0wDFHlYKa2lZWXPrAO
BU3m/9skVUp3FfuG7h2BATdk5EjQNtMPhTxHBFIPeM4ermvqPC6qCvui3CycFugH
/0yw6AwwcfVi1L+12MSb2HZUyh7TPJUR7KDVytfur6iOpkk4TNtx3lVu29CODa8D
SsLPtkpkNvkOBRcj5KHMt3xkhXArF8KuAP+blAERFeo5AP3niV4e7V7v9DTiUHRZ
6v+LXtg0gDQ0n/4vV8pkzI9mFo2wjp5lXK08mQHZmo2SJJeWgehuFmOa1GR6lBr0
bqHCHGztji1c/X6561MJa8FYh/JPsVLmCwpdRpb24LdAPbrVnapsZNfZkOYy7HCN
SSK4tTUE32gc2vQTUv0twnEHD1u++16fNCVXaj6ZGrnlfelRwRO5+qpQqH26YvyK
a3io6Mx3KU5dawy2LxopjOZu/F1O7KQ81W3Fb8hWw9XJkPuh4pjyEQ9SOxw+vPh6
`protect END_PROTECTED
