`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nav8UX75cNCLdGEG7wFlZbljTND3x6rUrQry8ySi7ILRw59a0wchwwUW7P5oPeaq
AhRuVCxdZYCC6jwrpE5RgpEHlye2F+p1GrPgHzerrmIqaES8BfxJany6opf0tsgX
Nhz77jSwYus3Zn8FkitmmnkBx2YVVLyUmBWofVqphBogXrP9uIfQOhnP1FLO62En
k77iL3pKMSTDCMbZpEIGMSoR77sqXoVxOXRSA1Q9I7E58NMuZtiq/Lz37MzHjtkG
Ej+8FDVw/2N6YoDMKp9W9vWBwR2H5mFVBBwkdtrN4kMKhZk7Pw1RyBaTul8+l1Dn
cNNSXWxgPDhh9EURYeEQao6x2oiEg136uwDFB2RarG8aK0NeBMPNemdZwc0RWwxZ
+8PcBifu9CmZ4D7Ky1dhQE7IxKNxFcwGaD7o8GQTPvP5bwIPPVcs2naYAilotjJA
x6KfPSTiH7sh0eK+seqUHpCW/iYrS/OT1yqhngjL4hBPShDO7gI+K/u5QSeLgpmj
ZXnZ7BwsOIysMAdztcQ8lsO+2syRC8BvyDEKazGogcJpmIri4WDkSXe1vTbNwnmp
XOcL92eUBKSLB3X09i0VjcBo9UULvd0pzUgEfd3R/8CeUQ4HjVYaa7QKjFbOO2z6
NvalUx5YPa1GODGROzjFLAORUYY8VYhYKfuQIJTMFtpJiMn2Y4Y9q/ujejSSJfP4
N47UE9LMLQzwh5W1d1b1TtCxrDQcOhxKol5RnUWsfLIo/Se/MwOA6ccUhzJaQgPr
PegED7DW8ujhBYedCIWEYg==
`protect END_PROTECTED
