`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+A/sU5jgViHNzWQTMF5AbZDbP87CkIgu4qfAV4/6QiksJr3atI9hoKFbZ6oCnJKN
Rt73C9d+LYEnGEIVixTmP7qkRCtoD/Uk8TP83TcQvirRdhqbl/nwvZdwtjq6KpfO
GOWhaWkFkWlFzzGmoRkCfjCeUDuF9x/XTS/kR9WGIYBkijAHs3W0wDbFHYWB+8BZ
bxpLBNiItQa1vW6YgH6wNOgg5zcTOrFB/4QmBH3rxcn8xbUOIW7kzYcxo2jMDdFE
pervCgS7xC7H02OO2fbX7PS58TNofDEKL3BnbaKHewpQrsN10XRUbRAqc5x3Wxbo
SDB5z+wkWF16wV0869WA6qmDWN5ZALWWmI7XRUkUy612BQ4/Su06nWZ7QStTjJ6y
qIgiKIt0zhNGGPMjSIz8QCNlMyCYusHkBQfu6YaDvBpGfvSGdndqf5JTXdJHKmHf
VkiosyZlmZt02EZddS+NidZ1V9tcuDwfSy8z4ZRaZ832/8XizZT4H0priEK3TB9S
+e42grIZt6FsVv1BeraXS8FfhOXn2X9usQ53BcnF8cuqL2AhM202CazWakRiBM+U
Cymzyl77ziurD1+OwOzvffTJV9itVIqW1YwiXEqTmVWDcLS7Nk8zCOWxjh7Sn7qa
Sz1Ubzi00PWQIkm3ZTychSXqz60D99szdH5CfIlmIjvXDhq0fTv/Im36/xnuDv+4
jeMJtcsGzuLHzrsoUne6z5cMB3RkYEpMBaGj3TIVja+owgYiPyANBQbue0NjqPTg
4uBdzIe0VjdX2KfyUNLU2Tm8koC472+S+88dtuXB7fziqrZts24ymYfH9N+2pIol
QAPx+XC3A0xA7G5p5AqZ+ykl+/jfzmKuIbI9Msh/bNatLcuROmCCZkgRQ3xJRBor
9LNn8gK85DvxKmmo3dl4HG3/ESKIGt9TqsGwRr4jE+WVjJdpP6nEBNcDRPJz64pk
6MvcstVMevDMEI7KDguldB/iWxkK09jfNR6XOiLBIVvyr3vKK4MscH9M1lraMpW7
miGj6X+9K0F2bSbQKpwLQPaDfrqryC+A6i5vJc4FJHtseSTWB+QOTbCBu60zlINr
cFxkeVxxq3nSbvS8+1lOajJZb9hiYZar6TsykN1EoLJxiZBvk8iTSxBq90xHgemL
`protect END_PROTECTED
