`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BekQRGuHrw7nBT3TqunTKOlTqF3fXNIuNLR39hwF8nlZf7B4kukvyHxhDXBnwfOi
xD2fnI7ZHrQqxUJ0qEeZcdinvkP7Uh8yBSnEyeW+6hdRLH/AzJdZofKTjLS6qlD9
ccX8H+bP+JmXvDy28AQRLKNOweL762tT9WQ6aktqC+4k9PpUK5JA5HhBxr6SALFd
wJDaj+SQchDL02fuVIEZDlBBvI0RO2BtZwwq+9yGoXfh333FZjBqOSUpPHRNkYS7
EJATRaLOQbboAhNitZJtfX+NG681t14H8LOSckgMsR+wz860EHtroGXhKgAn+lHa
ZUcZ0O/l7QtOl3pWDd1V5QmOboP2nDvXL2afhIDFMyy7x/xLiEJYSqGFU0ijriVe
s+29tW6CIJVPPjN+zryZvf9XSF1zicRYkTxl5w3V59W2xXCIxhoibyaF7Urne9Od
eIULOj4+7d2uQVwGhjSoMCyjPhODJDUIC+Bq63oOjlpA1JUvXlH++f2cKRWaumx9
FUuutz67jRfsfFnod+/3+tQbfZj1Tau0AMuqJnquUb9gjlPvxT9zG4WxsCd1b435
BtgjS/trx+gf82YAkvZ73ff3US28x34LYEEPgyHdamKXl4qflDNXopkH8aghyEtr
y4S0v88/hrK4vSBOKZDXzcaNxtDULRZ7hViV1tyCV3IXVoDw1NgDkupvBKk8fKA/
fxse+YitAE81kIbdeZu0Dg==
`protect END_PROTECTED
