`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+S6rEieuksF3317wM/HBReJqXFhRIVjWoRKcYTgqenumD4kYf07yjKadvaeB47Lu
rHMSta8KqT8Bec6xHA11gag4Wjbg12Cu9822v+9RMz3AGlRu+GXsAoNSzbjUgN0p
xU6Db5F/gcyHneXP07mqC4uTNof6hb2+ilOCAEOPlzCwu1k2GyBb7uRvwiwqAK9q
VvLMyFv6knJRLJCg1sEWvk3PUgIV94TJyYUY/hIpNmItiiiILoPmsRlVsUOD7Dx4
iUNJo3233FVqoEAjPHj6JhYsoEMTKch0z9HjGLMnnxC2004fMMhX7D3nfenuQFCA
esqoUJlDnU6DjgV9DpRlL8+4s5C6Hr+n//NBPMBbBA3wYdZ8P2e8qX0A7UOOolIk
3yGhSk2SxAeySNvRXbev0ZOlsH7pLi6/pglH5em1iUaAcfOHkg78j3MbfbHvYZM+
`protect END_PROTECTED
