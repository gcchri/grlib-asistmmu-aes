`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DmYpaNRhERUHQhik+rzEgSwTRhUDb06yBi6IWxUktcoXJ7nGtdLDq+UlW4eOaln
bL8sPpmPyVvQ2mR/zAUwS0fn2z6z7qoqJq58R/7Lj3SYrAKbqQgSqkRiEKUy5dsM
awKjXBoQsj4fa3WV7gemLPUhBoXAEbLSCLpufvOT581hfS775zvUKSDMGujVAAZE
0Brb1jFrPdCEPQ5SPOQ9W2U3ax2Z/Xs7EWQ9luz8okFF/zAELJx3o9arGPTh/F8F
bpuayt+zdbRIz2nt74hhUfhwu2VSQjiaQ9L5Gf/gtnNrmCvbdL2rol0swopF6kRA
efQa8Du8T6ECaeWY6n7VzwX1F8N3HtBFU8muOMZLnH9CSxUzlpSBbpkBkdx6wbT7
eSOmbKYnvyEAA43X+mYaN6gXJNYdgUdyWgp7BJcQZyxwPm9eEPcwvYzwvwhBa6Yf
liFDWDi0lFzEOg53M+/F7wgsLB7D84I0BflexaSUUjzEbksHCmHK4Upt+qcWKc0t
Lpm5zOXhg/kEhxtH5HjkLWyCoZXBMJfaizXSauwbSPtaDVWa0/KB+k/v6FX/fk6w
dNPaJQR0yaRfrkI/zkS1eT189s1PHS+usIcEv7vEj3ACsEnE9E19bQRA2VkTkOCZ
PS41DCRASxsNDFN2LS2gTdXdQaUQP0HPq2QLK49kjFWAzb6qMKZ3Ru1MZC6QdRgH
ZBWvkngm+IUvKTwdyvbgnra3z57srQqLR9SDUnVpFTwcXNqMd1oA2AKrOdDKJqRP
yntt8yBKRs5IrvekkPs81Q==
`protect END_PROTECTED
