`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NuyUGU/Zrx3FU+D1GS35IkClXgLQumFI6lSwoFVpkcHxLMWGIi3snZvhgYHoi1V5
8XJ1nj+M1Wj9nGQ9NtHEmOrx6x4RG+fHj+Ud8c65bcXDjCaBbWcuaXN5XbDknVVS
UYKCCmP3/w/5iq5ZTdpzcNqYZmKA3jhhtxanH712WFl18aDOPINRPtPROCYtIGDW
UEdt0CoCD6iAmP9Cm8y1YyQ/z1qauX9TSwNY51Q/KYy5S493DK43DkS1oWBi+qFj
0k/J/XW+L7ipsbP65BuyRlGs72gG5dqNhonUk6rdWquWf42A+AALim1IkHAJnuTR
9dQtXjgJAnqJ6qf8YIgMDeoqITfTQy4iEH5DTv//hjI60Je3JAv7wfpk463Q14YU
LiqTWPSs3hdHLOJdZzVzpHnTenqErvv9s4zuWe2GGBKiXF7i6Z+L8QRn0gh7hdky
HtHEohozU/YrESVJBkiAfPgJURSkJ+4r4SutkPyBW0vk/4XKaLYQrP6vZsoGAGsN
`protect END_PROTECTED
