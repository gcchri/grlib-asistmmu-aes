`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z+V6obOAgQfNF/afkcfD4RzOudLjofCdUvBNZuN8Sy2cO9v/yEV4rcSIjH6O3PA/
EIjHfS1HByJJbeB0gMPX9iIWGoT56rsHV3tmkK5qJ3qlci/YZC8hia4LCO98xopg
66sNvOE2poK5Txj4UD2mZX+prrpuVJfi4gxdoxDCm/Fb5YaOLcn6/tqsnMKOpuiw
DIHjK1MIiESRJilbr6Z0x+gNC+rr5vT300SxWQDRJlJzg56iTBLGNaZe88+UvaDu
l49Rd/Vlck+fBCkcncvKkQ==
`protect END_PROTECTED
