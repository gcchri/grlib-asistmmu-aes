`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHR48RC/e78GgxBm6HCSxwPWRGjd7kHGB112u5pWqKWnNme4sx1abiIU17TMIPIn
w7fYRoiFQpgDNerS53+SI/yZvGwHodQyBra0VcSRxTJ2/e1IFMcxdxWdyjCskjMC
dBW0FYb8wfKDpFOmw87XhNnsGQl9zFalopNLdZZsC10erbn60ntj9ajnuG1q7pwR
sxVl4F8h4U+GWtbJ56ltVZabj7dvXuZKKvS1/4w5Djiy6gQcv6cPkInd1yjOrfzR
AZ5lOkmzm0s8SCNWg474z3VuyJmsEJK24uZq0mTNSfBCHL+6vghOMTcDsaFjevPq
41DAWeLow+V1zqmSjy/szA==
`protect END_PROTECTED
