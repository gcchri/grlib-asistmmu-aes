`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z4LTOTkgsqaTIrQl67sIENCb2HepPgnBsdv4cEgrWXgKRVdcPxmLznp4FUOzsDq5
NKkn9uIz6x5ysfASBy5cYAUAPDm2ZD+0wLFNNSlUThaxFfQoR6ea/cj5WODfIt69
PXhhxP2DLvi8VBgwlkN1wejvlQsBWAsMdgfTGyxJqeZglkhRbEDpSWZiw8KDg7Xp
CR442KO3NAnWFCdzQ3Qs4mex3lsu1dc1Xsapkki1c2pt5PMIJauzQOiqrmED9NCR
/0Yp2XFX+FaaAySiF5y3TPiKyQ2iSHDaRZBYekuZHXXZPLhB6cPrEd/7UiL1KJKB
2GGm6A1eVQWMFP+0UJuFJm9iaJ6lwbfcJnnXUJqIIVjzdP+Dr/GRqChk3FKM+DS0
dMNEVCii5lmbY0BqXHRkhwpT6eit7hJqYCjSFLhFJ4RDm4VzzgXAeVrNpCNe3n27
`protect END_PROTECTED
