`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1c7a8jo51iTt6NWH//S0/STsN4tzZD7loWoJ4u5tfxCfgTftusjAiVtDQUynM+km
YFOI0MBWHFAsHN4By24nDTrOknKr5mLKY6GE6O5Le1z/p0YQ5gaGLfwo+SHFxTRA
8ASFFO654OfBm3mJ0fOCPFbPV+cM7Egx3C+1njFjBMdBfwfCs1p/HAyLkSKdRTTO
6nruJEpYj6AZX3qjRv0bV7OjqOdDZi8S0jPCkuUUOf2T1Fsb+HDrXw4IRyE1HhR0
ovgMt4v4UXidflPQ7a5DoWP+vG38hTh1hjgoutSPiC/jJN1f18mSHvVlcRj19DWc
3S7BarR72dAVe7GOb47vWEwUypTRzbCJkzH3EhRwuBI/xSVgG7HY1afov6ClYb8J
9I9SwYA6JyRafJhkMsTJJYm0zx/Bd05nphNAbJ1bmH8V1/xcxeFnWiSQOT2A6cTA
fSu4QWHRtqcsiQqSA72EKU0oXPCCLTxsG3gVjU5w+8G30UgEJ1HVdzrazB7srIfQ
pt1ZcA1Z6cAXUlw7YAbiuO/Rpg/F2WgOT7RUjR5RLgtL0pARQTWvqhQ2YmJRy4lf
A6o4PEeuD63K1vpaLOoljeUF+LMsBAi0Ry37zAnVp4Jalv5yJrP3EpTboMqgqHzp
qmuZntG0uMUgrCKWceFKwiK/+VisYNVlst94MwqFr3k=
`protect END_PROTECTED
