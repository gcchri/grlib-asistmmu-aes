`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DhOW2RbpTSiwiRzvPCbKCFTFp0TAQod3HhURS6dakpp5sCEyxXckkalHSVrmCMW1
QYyRLtEGBwQu0gGHfMmZaV4ziKbFFCG2KUTs86UdyzcUpFT0v0+GyCq4+jyaHjwY
/GAR4vqkRtum0yGlozvSNX377k63rZPYaw9AWsC6UJP/ti2U1JS6MtR5ZCBKBxDm
woT8hxZCmvx8Ivf/rJ9llFvKqlf0DHMXe1KBTRydY2OSrbcZI18sku4rQkGxBAtN
BWzMMn6O4aWsOPEwOt5jtjW82Amfx+YlYdl0E7mwVPm1YTgGUbs15Zs4/FT2WL49
aYvf47OaOnhz1Z4iCd3nDuQ8XPcWE5zsxIQLU000TTtojLHj7s/tms5uq+0X0utD
XEhH3UKvQvhe/C8GdAWQ+K28rS+QTlTc6Ztq9XnbdTWeUGSYRNqirbJFE2MKJc+w
SrgNWa4E9wymRwmsvSwLojIMJAfPNK9aDmXw6DxWzEm5gt9p0tCr0m/8eMJ0Hs8n
wP3Lhce1gmuhMEbiVWbXC4gPkH5y5hda/EgolDGjC8E0az44OeYb7kEP8rxGAKtF
z0FDEJa5o91P7D/2KAeexDRckgckVbommxvcnN9nE7N/IRBFfWWMIlFQg40zuiwY
amXOK0+lDtpNVpE2KKnjAy6628OSlLRRt/cnAeXn32vM9DxZYfyJGO8S6i38ISwI
JhRi4WkSPzGo70+BvTiG71u3SaFpXqxjKvZHrCnJBsDyIiMus3JdbX6mguFpJn86
D4SzlyGWqFUSQ4TIgn0MRw==
`protect END_PROTECTED
