`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IjD5YzpNF2mRx2tXKEsg9iJLAB1H2GlsCzlY9oFRsKtE4vgOBO8OH6J8kBZ4nrKj
yuneDKtsv2waCnyBea6peDPIDYCVE0PKhQE5QWC4uM7M8o+UlwXsTEwq9ffAQswu
4hx0vyYRAMe0nfXyqizaumSjuqepsbfzu1/2fZbifv1KoV9rQIpYdhK6zFjZXBJT
Cm/Dav73nqIAM7zTV4E34VAe+s9FOpJUUCA+WREG6MtE8ABg/w2IGdGzcOa49JLG
Pn6AUOpyIDUNtNkZJeavm4I7i6c5hWFKgMCyQD7rMHLZH/YtJqpPkwkhlH/NfagE
JEEIn+opQK30UAJSzBhmJRKZhNDhsK0ji4qzn+HCYI9C8mv5CSRue9yWEzh/jv0Z
Rp0pNRf1vKOn+rSV948M/tAj809s3dMN/FCc0/3IOm184hwo7ywqQdaUn74OR4U7
m85z1C3PYnPi0CAVclDX/F48m7kjAJzyXX7cXe4lPvyCfgRrhzRDIT5+t7O8ZA4d
`protect END_PROTECTED
