`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVpYUc+hOnjMheT4JlNX9Qo2qxuBi9GGcI79hE4/dHBNL92JxTWa2e91vf+g0zz5
oOIasBEljl0aw9Au0mifc52FOnvq5k7pLrI5TyUwtWh69AsmUnZBbwXb5CFBSJt3
5BBH2XL6m4T0eflAklqOP01PE/lbg98vprcHSgpBewo4N0A3KpDECpzCThlWOlSw
f7FqOoYSa93exVa5EWFOirDGlMR5fd4lqa+X0fXvU6sWkqFdiHkh4sZTjrnHei5g
`protect END_PROTECTED
