`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNcgCXyPzusTYCyB2G7hESJkQkbvE6cMmjdONZpj00adUgBFhkad2Mxz+n11dIn3
qFSMznuGpfgIQX+dehMWu1Zs1sPkyfpaSdMeMDw76/w5W04ibRtRSKYzUInS8sqA
0eJUWbe6veNjZ9WKXLoUoMM2WW8bG612xjZnGfgRUkcNCh/WuNBrMIP91TFzeY78
nqfdXHUHybTpKopVjoqc7RAJ4TvUDoVJPCmTMUvCsp3OjarCiov8EKBtCXw/9NPE
/hR2SqUodljSLev5AKMG1V5ZD1kuZBPfuXkIMmvsYpU=
`protect END_PROTECTED
