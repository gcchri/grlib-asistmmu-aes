`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GvMxCIF3DliPLlx0zqOrTeS8LwY2mRMS+EuW5SUEej8kQd0/vYy1ttHSigH6EDHk
gFlo/tSDcCSGJRToeqB3MD2jDzdh7amIGEs5uxP26UlEUGFGZ11leO6Hk61ScMsq
wKGYdt20chQp/TIYaiU5d4TDBVBZepg69vikPJXbvKLsMKfxdfiMNdwLNvU5jc2m
v8xdDLHFsDYJvs2wl4oLcUacp+ZZFCJyWKlspOZQcW5RzRYxxylwXeE9hyO3I3Vh
PSnUAVvLHy26a4p87CUFNzt7Yf8Qbp+yJDFkYvPhotoR9r+S3en03nVUOXpaopKR
6B7CO0zUPveQoXrUii5eZOm7Z9XuhilVlqeU9oF0T72CRfu5diWr+LtdS7/1hpDy
/I8FPLziiVrPtLPKErsoevQiehI5eF7AY0FfoZ+G0nqvuEMdiaAQfuQFWmV6qSa9
`protect END_PROTECTED
