`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1BlbZ3rBRbYGrPrlFiAXx3QetP7X3lnihLT9+a1Ybd+wTApjERgyJj7L0Uk2Med
KfrUIf8FB28bM7+Lsdjt7EBPFqERcMDuTttRwnQNqgkd9ByeFoZGYxC4INpS9ByZ
fTFbWbyq6NtKYAbRqJGIWnks0xGfHI4wLxVtoPlQQci0hlKGJs4Bw7i2+iMD2H1l
3Rl2BETyycrQOOOeLjEozOxH3ejhCmiwos5scoh+pke23mvRJkhFRfY1R4pJL5eU
N14dEcpstjoE6smMVJzp+7THSTOi2PTlVV15Zbwu7912CPmZPxu97BhbgwMmmTod
VQtKqU/VAfEJ81tckO5dCM8vR1574d/UyKDceN6lwuFxGlLTffqIQV7H9s3neKmA
3dSmRhoGmAJB+2eaFvTh4Q8Yklgzx6cGjX6xFCw30PklC3ffxFfx99QgczmaH1zV
XxDQemqRVBveA+yJrljYpqnpDpaGQ7f4c2nET08NMrvy4M3tcF4zf6TtMyIGbOSj
FSAAfP3xsebglnVkWFhdLCt6YwBZOzPmGjG4mldIM6HUpRDAsgcXPZVxyTIlnH7r
zszqng3dnkiZySl/uciKJSPZ/xaYmePYNg1WO7O5DfxZCzlNpEpk/MZDTpEplgrC
+F7U+6SbZBZ9PLAGZhS9UMhLIInzs0CV/73xR7MMGKbvcLAc2cPDVibplGF8pnHC
3DEEJRHW/l3MzVhA36VHjRRiTYRkedDtBWsPib+Chv3ecigCGhNvGQA9oh2Qglfj
BadfrP4L/dOvWfZe2vgDnbQrc/UFXkR4gu8OmR9nCqk88lpaRkEpwrWrEIFOT/zx
IfKgSLsG6M7Px2Kji3ZPZ/Pd0hVdAFH/5rrdZmV3Q74VdStZ8Em0PJ6t9qylQud9
DbAAJ1dm/v4/eQ4TbDDjkjCyObJrTzXkH0MT6ylHn5bK7tfuQTkb+I9TG7GCdYk6
2NC3CSxiQsZuWvinbvmFt9dsTuZLZmJi6YZUbsa9BcI=
`protect END_PROTECTED
