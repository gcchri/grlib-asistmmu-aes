`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+JkwQNw69aL2vmMFJb5n4KYkhyGiQjiR8qoiIpCr+R02cXF75OGWwLmkTDUk98M4
JmIV04X1EumKCmP3Nnf6h/B3WYJop9U876oytZbQjo8SjHFfOAKb++9DO+z+gtcI
RarvxCW6kpN4lcuQeXipb9FrBzwur+/pZXz2E2ci1Rbvosvr45ZIqq7KhcyHIQU2
mr8dOTOIeM+bkt86kwG94UP/XmwyGnATg+/4uu+dv+38hZnUEAP+T0AJ3ICMRk57
NZoTFwM1OwnK7Y9A4/+sh4487VzJwW9pw6fSuRpwZQ3eUNef8gTiIOM1WC96iKpc
b5ZS5ehA8QIlhSnWjUp3OVD1s5go/QAnlLoZ1vXuO3qP3bu60TOz/fqe4Z91LELy
Phm/z66LkCE0TJJBdnw3fBUf2x+eloyOpHz7JqVUTy2C2N/f5N++tyRyutbV6r1h
fr2CV3yy8UHNBywiEWv7FVamPn7GNNdUD8b/uRElyGcpRYhWS/N2NS+7p4vb4fgU
+BC93HsNbVbfl0lDkojW8oJiRcehIGhoEOOgz8rqOM4=
`protect END_PROTECTED
