`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqXtaSL4jmYjquui/AqJadk9kO1IEbv7vVBmZtQXUP4bn9Z++kj9/HpN3F5DHwrS
Bl7ChLarzT/2ni9Kj5U3B5mG490cB7t04/z7+DrcEeg59zqLt4W80XspW7z8f51Q
vLhPXerbSJ3GyPTBmd5v7/swzKk8roL/MqorKjoIkvsHvak++h7JJ4t0K1iwVU6X
2PvTLjfCx/BaNd8PQ2g6fKFGg1PQDl6+M32jg+PPby1eISyajCVfZHe9S3TiGSPh
nDNvBY//Ck6OAipfuywNhoLL+bODJTQhiTBIWNaAHKQx0NNASoWBWUGC+19h6JTh
gqY8Dkbcy2OtQw3k9fJjMjgQgHdNDl+iR8nu21CbEgmlwzTlU7QEg5zoanASLkTM
Q5UbOYLo1YGAcfVP+oCWs8ym3sVFq35ST3HlvoXW6iOui68aMuSp+g+/trcoypr1
nVd7Ic/e31MliZyEMUuBzLyP/+tRcPGIbHVyH2p3VoIqTpRVLLoKR7MRui4vUxdm
pzQZ6GJQlrp487vFI1TQPw==
`protect END_PROTECTED
