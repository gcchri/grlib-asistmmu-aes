`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3Ai27T/9bdcJlKIKBkp1z/+LcJR5j8Xicch6Ji5MCz5Iu2lWdaThin9b66ZEQzh
2g+OFXifxTEfl5FRgqi//CdotmjroNj4JTVr628+yPuPjQ85JpEoiz/NExhEmUjI
+0LKD6exT3E9klJXKI77Fxe4IY7YU7W7cY/wCpZ3KJWvTXTSdcX3LPCyb7WPWdkp
ZF2lw8utfFDaAPjvvVH4edjVH4pum52ij0K6oy8REMz6nmjpuzezB6JFbK8fKYqH
5HzQs8qwWAL4UoAMUX0/+SUd3dQ8OrQLdAh29Blt7VDaZg+w2foRFJIIpUytSOCN
tZc3DPzO38LGuwRvkcJMEQwp3s7QMWP8MKowHeRtzce0W4lAJWYUtChbWejyUG7w
b7V7OO6dhFkylv8ZUOWSxniJqFqkupF50q9AA7ibCSYUzPE/VegpynvXYXVB+buQ
lZ7ueAzHZ+x21MZyTZha4WE7X/fTtyrT51mPch+emKYejkRTG0phdVDw1QgDE8tR
tTUUu+lWHizuef9be2lZ2/WXikOvFnhWX6PF1sFR90tqBeUOLtTYrFATrRBd3qo8
WVzigZFGxfhErUdlquKpL9PMd75zu4BX1qNu9rbYJOfmcBls8qahgN29HFzx1WFA
VsSWBO6l20vrBLrN2ysh6/MAKhvSz5dp+es3JZOEcsVaWi9sR031HSQZCzF/L7Yh
ZdoOv9MvLXYWULdsMO828WtGmOaQ9vzCAsb83zRZNQ0H3Z0q6SzTqgGo9XxJwyc5
TTVn7ZsTvZkbYFLuXiNKblvwKEiWZ8w0NQhG92D7hXYqdXKp9KR4tTOjeR0mrMkz
Ui+mIo5whE78zOSMrGuDXG024nYFRQP/rU8NFuFjCjFIGUuoX7MKo7emIocf5qp0
nBvTkn6K1dLrR+HEPZcxzusW4fGhfd56YHLRZaMUlBM4+UkE4q77C1F9PhYCTeLA
hos0RWmVkAjvClZ03XFijLnxYShRxPoGhc+ljltmjBqcGXFDhO6PyIcyzaw1K5fS
8FnbuVgc9giHkL0rV0W+oFr1oerbvfeBcUjp8WmdujVDKeDBNjrV1CSQTig5rwOk
5B2aKqK/If9Qb0UeXZF7cWH0pbUBuM3xsI5YQC6C8cQGD/nuWE1rIor9sfpbkQiW
efDy2TS5NgX0Wq32qkVybgDvzjD1H2bXFBxl+gkcPKau8e1XgiM/rpO+JCEhhWKC
GEQNorS2fwEvrfOuafARUND7BBPp12tTp8/Pn1zUkfmz2UlQ9UzG2UobzC3P2WFF
tWNT/TrWk3YkXLsBFax4uI8GOTokv08GqF4IIOBbED93TOSrFPf/nlVjH+BIQNI9
JOijrS6T4+HUStrXFMo9Yu7Dnw7r9PRBc2LgLS2Ij6tKkh68VuPbt/EQ+04eHutO
+08r+SdmljwYSYHe89SgfoIQOYm438KBNXb84nSzIX2V9I4lOT38O6tE0Sp6M5S6
DW0C4i2FzH6UMISGqTxMqalX5XuIRgkTSqMSIP9zCFU3ChK7ZCT0aOADD6OrNgZ8
IHmojdsY6ndvoVrugiyn8bF+5BDJO9ydczh5GJFTp0KO7oKQxCtMYzMPe7o9Ijhy
QQ2wT8MtlV1DIfHsr1sNTD4qypYubs5diLC1hjN6StxOgIbi3KT0enn2J0bcWUVT
3opJxjz+1fjVBH0yxhNGXg2IaF9dKK6EVijnmiD/LO3ZQKNct3y0H8wB5Qq2tdwR
2Hh5CSY3eSJWPf5BNLkhpE1sB9pSRpB1TI5x6z3v9Sxm8lv2rMZSOTcRXiwT1IoK
CPuydrfobUvjmtK8yqvk7YZvZPd5Gc5b/1j+u688rrgFFbX+qwk2Vn2q5/EHo3iO
IMRIJHSFaphEIRXcsn3/lTenLDlkg2YL4t1IfWpa8SKqmLVB0/zFLzHZSPeyUR5E
z1ZypWBXw7IDf/WdHwnt3C+F9rPcbyRUgoRIDw0QrCkbQvx9nPNlfUFeaiosLM+U
3QFHJCRZW2Y4n7jiNWWobgkujegRL5uOF7a4A1AROLYCQcrlcdWgFhqzTzxCUwzS
e39+4wcd0FKHYSkusWbNn5Fvz5lxCfpeHrSgHMa3icccGUK6oPkcLtGydCAVTIPO
/ITnIA81fDIjKjkHyRSMe8dlagfGTfT8GwKZ6KJcqg41PditbQIY0uYv+L34lysy
GlvvLTzjiblkAFQ5f/AyuBDaR7kZRcSpWvl+8PG4Qbr71klGN84YW7IBFDUib5EM
qG3rmXdyOGQAH0Iv/U52kogi/YKjaHUIfpTfDPLHj0noPf7yjlCUF19BRxJONTir
VRNow4qMfpfc7DfyY2bETZHXPZdTM7ij10SFwm9I/dsggngfI3xAy5sNFs6ss0aV
4fr1IbHsvoC2MxBI0iz7uMjttJAZ29l0I+x10g3+7H3JTL4Ojk0vBdnUS946gwxg
6rypkW5FUefHB5VxYAP+J0sgkC2YS3MAAypTdn0YRQG8cLTxLxvYt3RHnpz075JC
zTx8r0Y0raRaInyCRi1k77eDViAxWuCqFm7UIGWAYe3C+GV3m/H3Hn+cJpovQsSH
Xk7tTHf9vaVxRB4PQpllYnMj9gIt9VKTY6q5dGGq0jfl+WdAhS8aE5iIVMJQYvHz
tkPnbePqWNqiq5pRjxIMCA==
`protect END_PROTECTED
