`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qJnt2vMLBXWdHyaIdVIQPZDnc8+KMzpWX4TT67183S0hKix2IeFcXfU8Cdr2mgy5
0Blh0tOd87M5rE2rCEsNleVpZMh3JciQksZX0UXS/KR04Ot+JjDxeAuiFdsid2xu
edjqIaCgEQSOgLp1OCnZYeYRWZsPv6XnyT4KiT2lakpNFScFKzowW0cdQodkh/GI
oOPc+OQAHJdQCQaLjstIP1IIsPD00TD0Z7DqU+AfAlyWaBrKRmrDkwzA6jaMbVcW
j8tcFE2/Mvh2zj2347J6ItNV7zxHmvBflrfFaV8207RGeTumKWyUwVNQDKlQO9eR
XRRmrwaxqbKFpf27+fy+oTEY46N5us/bvueSTNLsD40wtsCwCloIa4ZjWmHICclC
EdDOm2lTsTJEFZy3jVOP7k2XUXRzHy45IGQUPNeroPI=
`protect END_PROTECTED
