`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Kclk5dSD183Rpxj1ZPADJJLdEd+jbXxkLIkLD3eVN7W5wfmJToEtIjc07mRz3sW
OBfqsjiNVOjayykKQYUj2skO7MA7NmAB6e7JyTkpzoxkkl7GlxWy69psOMMwQZsS
a1HYoQV78PMlfJm26fg1LGmHD0nINJzC2m+uqqBa0m2GrfCC80iiCNvdZvNpPOQZ
hkEj31fsJxsQivCVNXBK/oeii/naXWNp49hKaG5PeQl4dEPv+451yJQmNgGQ2iOw
ZoanNKi/xg6njcYvRTBOLhot/7YGrlK3ku/dOr2sPeL1H9bFqoBJNGB4++RHvbKX
rkrtrZnX+imc4Y8h6WJxgjhG9G2T2M+XHJkGp0sY1AGqg3IGK09dfiXt8ILFUxHL
D5HsZ7ZfcNNNv0SPi3x08pD2t0e/VBu6B+I2tb5cYVEnJHs7/XN4MoT+LtZ3MxXI
SNkfKfNsrbgJ//EwiEeusGYGZQ2V1seVi6AhAQyr1p9yNeXz6vim4BD8DBWp+MFA
DqQvWsbf8TyymCq9AqWhQvNxwDSsfA/hIFhdH+W8vwUEKBfS/NlEzyrrSeL52SSu
WtxEy6RDxrT9oLh9M7tR5aMKxZ31COH0AHdGo+3woclPajT9eF1WTa4YlGPIMurg
VjbKQUFTytDOdqI/VH8mpZ/MqIsIUzfmd5mL12jBwlL9Q6Rd2bXpF6vDWS3HBqaJ
zrQKe+0iT9ObfRE3ksd8CAphygh9CwU0Mdzetyd4J1iHu9WpL2oGU7J59mSprIEy
9j2hYG39g6VWnG9ySnUyiqtdzD+OlgxX+3mhqTwNLjYD/iQy5HS91wAXpqURjz/G
wmaZjQpisnsO8Ilh992/EMx817AS4XN1xCMtjBheTntjrRlj3cU9ItZrkH/UsVF5
/imycFeccLchAIPoIDZXekHbOI9JeuXoQrOvp5dfupLrCU6W4LMtpSf84vizDHAp
KjKkSzVfbeA+Obe30t/+odo62VtHT/vb7YBD2sCc+VpP89a8xIB7POyogVHQv8zG
b6gEOu8pZNY2n3LUoZCDWaOoqKIyX3voV0whctkKNqCLsDaWQo6bpS8p3fG1v9aX
YVGctM0GCQ9bF6axsjCJVzC+z/9Vc8EmW6qpNKOCOlhDHow3leqwovPzZGOxyo5D
WBcemyaEpxiviRbOKaCP2kzDAjI9YxVyo33KAxkC2eWd+76bnz0mzdHyFm9jS+qs
HuIde2aU4yMFo+fyAMOTytgfWuGiA9q///hJ3kAGcyCl4AuO0VGD9lVqMbEepwiE
4OtofypxIR1ob/mRG5ZiZN14GTWNSOLDgboOgWw1EM6gg0dZss1F2Vj3GnJaMo0b
SDZjTq0UvcxRlHpbOXlq38a73xK+4eHOk2maSfxhiF61HOpnXD7Mz/WBT2DUOtYN
OWBBCxlnXNgqYgArKPHHdoEwSsGoIzi9A4Z0yw37+T+ZNxLU+xP8dZ94gmPD+vL0
5Xw+/zqVfwL0MlA27RwjdbOSXVeygDyYUnckPgJVWEv7cehS0yInh5TdCgEKH0YB
2YRFn5zxvxNCtvPiVMD44bR7cpA5O75OlTbEmirwKfCPaXQ8Rd09Aj9QproQiAic
9gPj3AeFLC3iUZoLmVFhmGM8HyuYcqukQYtRzITEKShv3UlAWFEuw1aoJfFRbx3O
C6+CA4o6PftJHq15TWJPhGeozPhZk7KU/huAvevRZgseWrDQdYvB5e4wRUNwhT1r
XSCcHK2JVlMD/ooQwtwXPWsQlMmFwMnbmxu/Ju32J1lZ4c6NyJAvgTDZ6YdkW08X
/0WTic1N7v1Tkcle5/klCxTg75Xa0pRv3WcacA9v0vDI51T67HTBT6LoLWDHbBvS
w7FYoAz8o+zbT2r//eA4i9yIoBZCPq+8CHS8adp4zRdQ4c0okFL4sXEWkOSFPl63
j0i7c10+ZQBMh2eYsp57vDho062y88h41TFU2knoxTGua3/EzDQm4DijTOQhyBGP
d7NbwNhY9wuVWoHypdMjA5H2FmcR7TnmB2S5XB7yLdCTjDYKiQGkbE33K+QDeQ6c
HfwlYwzJ8SPHKGIMPdcj3ez97Eb1IpG3uFYx528lApEZB+sqB+FhVc1vJpK3e/kM
4iMUc/eZRvUB+BA++YmBOKoFzgu7bwd7XUCazzLMU3hBx/IK/0hmZl7zd2XdiYV1
vjPPlEThvkNMwihriXBZz/tsfrR5x1nTQzQ+RbYLyKBIXGVAcK+/VMaECKARLKIx
UfkmKRaJ4/mlyeVQ5UaK0aIXkFZvpR+kTeLWfSjgfmE+y/BGulCsDgoARTPVb3/D
7VdWiwdRpLk2TtzE/pO6FbGVavZyT/Nk+u+3KRw4qKoukvi9uxxfYqP/NmajlZob
vfX0IE0A3gQQjslz58z1PrWmJ+/ysK70Wupo7R/DH5OYYeVoEfSxSSfxeDqn/GjJ
LRCWkl7D41Uin7vkyik6YTfUpeDOb82TYZEAoMbesfDY7g3+Yp7BVTHstfe+vGzX
me9KrucKCFS53yJ+7elC+g9820aiw/XTVRR5GCK3Z3YIBmJC9whyhVeoomwuSLW6
Fp3cfOtP3JJiU63N8PAh6oKXOR3t8M23tq0WL8xHdDgKIBhwqobSWS4s486RPE20
qr4Eu5YE6992YFNs/IzGnTqqgMlKVd3ggxOpc7jaU6ZpFTVpJgSyG8cCc7M0JKfK
bYSTVQEt4C6n7cQOZiOw2P4qL4M+hZcIUfC6+ImcnO0wgYUMb71PjStKvzWYGcsg
cBRgilkWWXdODfuU0yRD/WMBnn1M0XSeswW8FraRvvJkweNNwnBNVxIP0ZOqxGBU
hoGr7OhHYxNy+ICSgQ2w+lOME0XD8vpUktg9JB+Osjh6/962d6mR0595vm5D1Z9U
nHfYZHFwdoJOjkX0fW3+jqPakZciEss4lhl4qF/g1JooPqD0AjZy6kGE40eEvMJv
M9XKtFkDkcZKOiEZvFtkDS7h9/ZbE2s18N3VeoX1fIzYaIPdbcZO8eSRSKJaetDz
p46gjBONSz0Dqaa8rNQxTjDgCk8aA1q3lDqP8WUQSJH3kfBxjyQ9dkgBx+Ixvn/B
s+kZzURJnQTlJ6WYLGXgkALc6c4jSGgstHpWeD5KbWs4X/g4scIbDaK1xT3qUZs+
A1tTyIEcTSgpnTEn5pYr8KeTEqOGEuiunkrz85bXuWiZXXBF9eoQ+Tym8svffsLl
EMLUxAiDn6kNM2rJaZJR4XKquR9HR9S7n56eHLG44VxhVCjXHPtMx4BUNh4zB3se
W+j5vEZjr9bHCNgIlnuUCAKj1TYHZ4eUcomnkax0rha0WMjlIst9gge4O69tVFSt
QQ0tqi9geutUGZHloZsHbzOpB/tY6cEhhgpHshJ7it2951ONH6Qg9ztkNBIcvWhx
4TZ6VV7VNhk/VNpNgDX+5ob7ElmS1aHgz9rqIGkwhRMYP4fsZCLcP4Iwu8ahTLOt
F3KWffYtvPP7PVauMkq5eNKVLYjGDw1Yb9K7siXPbu7MJ45g7i3T1E+2Ee6h3lAs
h4u+viuYzTenfWzlUIW08kIl8YuZZFyETdZvplSHu1/gtr8AFtzDPApUPwlFA5Od
ahfX62q0qnMC3VrQv+sq4WlUwL+hHLip4igGbp3fdUbn7lrx3AFPsq/szUyQzkMc
Bj8wOYbR1LfjvRjr9v9AdFGEQdsW+gEInhzdN/1BNWCPUPUAWBu+P/XeQXhHq0X1
qjrnyQFjU6gFN47tJeIoyVh9q+xhQ865o5y9Wyr5IRfs1UUI5L93bfYbaGdgqn/s
bBicS1pXW3mWYWtZiwjpVZzAhQg0SL+6XJ0XmY1/jSLBHstC9oQGn8mCPgYDgRJh
Mc3bRvTB4yxYscC72y8YUekOYmQ0yXRTzdUaGwH/5fIPArWdrNE1+ro79T4nWk5e
qpZaDFBthC75xzIDWZk//S/3PXPRvFNhZtVwLq8/LJ1c22+LrIOpkCEyNeAf/70S
6AJ/5kaFlgXSmfGm4YAyBYugrpiH8QuQm3VxKJp7ev3VfKHDcJl+4KYABmDpwCY7
3l74aJnzt8M9FGsfQAnKo0GyD+8UjrdFSFxqSyxbLWKvwk9bHCXgUGlmw9oOSyMt
6RxCkR/T8GSL065XTOWVx2dvbf7ksjr49ZNIVdKGEUF8lv9SwFIrnm74rISnNXax
DsGtd0BdDMS5PWAvkhvq56J3wJ7AjD6OGnOhr97rqFBkJ1BAJpw2Z/Uqezf2dwuu
RBhJHy2Y01LJrCZ0H6TkK9Es5I7y9nwQn5qsg815HgtSXymhRUMY8vzDz3ZPJBJi
8IDUXjJgLF3x6H1OAawZPcXjMGk/7EKbrRNBU2EXk1dSvpEAn68febyRKrmBV9Wb
SF8+rOuRkcrr6csdG/b5EzxB5RYZ4whUJ7aK+o8/8BRNpLQR694v0XWJ5TTjcnbw
CK2Xak5N3QLwC7V1He97EwmFzt11Gr2tScRHXMJhVRq5+haW0xAA50Ox9l+ZC7j1
7XGj0lo96AP5NRwDMNlOfLayyfnKA9Pyj0tas9H6mK0C0rFOCnkbDhwk0nuHyP24
ICc01uQOfgEfZMPh4ciPkSr/fXPqnVDEUFrqg/ZBxQK7d4CVDekUs6s6EZIiVgqT
YynTa/MfwRyiBWugMM6Fgpts8Eh9gGOIIvpp0nE0N97escS4w+z2Pf5RmgCX7MVx
Ki4KdsubeXQPMxQMSvafHWYA0HapYjoBFTti35puerDxHf0ZSpoaRoPpDYC1R9ox
UyZbn1MlNWzzaQYe/n5ek/mFzQwsKLqX7ebQd7hag2PswdpVqR8ULhUVq3rq58l9
9gVZ3EOrYvUv790GfazUGQtsrl4n7qoprLuR+2//tJzQQ7GGMBJGnQSLLvnWG5y3
fWdiryx7/XIG1Y9sNGcZv5pu0h/OHVFQ1TiScfZ7sU1RrawanzP8y7jOOlUJh83k
0t+vMxgkMIjWwR9HvKfu9VUDZxNibuludLHnRu+50MUt1INl5tDY359GzPk580lM
drToWKhLaJbl5pfgRwg4mUjf80HIvllqGd2UlnSbDkvFVtgmskry8eZyPzg+3uZw
egbzauYkO4MxGctqzybmJchOFdN9+34uiT6co1/U1Xtkh8PPE2ZANSTSM3LPTUHV
ELcV2gwcxZnF7a/oXVLxJzyvOoXJtWvb5QwQ1ZqsGVOhJSlcte654Qf52HKBXPgN
dUSv0QH1THdqxAeixZRvNmn0L7w8lAkWDy6zG+kJqACjZb6H5EXMKV+Q438bfjit
IwysMxcR2iVUl3TZRE/RFM+kWPyA9n2FfliPbOkX1z8DoBNR4O4gy82VfALLiAGo
PJKEGzWratebYMBFR7KmyQug8HhmqPUI1C55RoUl19YKqlEDBB1pt8Yn3HCbwUT4
7Zkur6TzmmKtX0E0LI4ZYURKS9/bRZFttDWk7++LnNXqA2ZKV3bRS0a9V3HUu0K5
hHsaUx/6g4DbNDJWaYzm3Q+eiW3tOYOUwvmp3+VYTr0KpjFDMb3vIHWGMyN/V2/Y
t7TStZtEjaGWsWTc+frqJVVUYuJ23w49hEPdEim6rPR2Y54qD9ZejSM7b3IerzXE
HjrzHA2SrqRvWl7nygO6tNu1Dr3cFt055x8rnYZ3G/+QdCGTeJThRVk/E6/6APCw
ZKdJclZ/AaX5J4JhXLFpRadTmV6DzH1o3k7WWHbkA4hfLOotwfwGIGINWM36kYrU
9ba/e2M0JhEMRTxPBRP8tYviIbkNr5yokCO+FaWxUbo09DYvfgsXkOEERgpLqy0X
RbrknKlOp5inuJIOVlrAWw2550tWduXE5SKMKBZaj6mTsCGrnpIIG4WrsQJRddvB
v/3hIOa+8g24BzmhwughAyvFAojWoLvN4sMgRMi81S7qvExqMNiWmXG/ZBc4r4JC
hsqTBF62SdcHWxqA8wos4OrHdu9PK971im4X1+h9v3RvpF97PO3LvqfkXmpSsnwN
WXIOk+3u1JEOrprvVLVD/4uuqp728rmf0jWU713gLPZTNv4EusIWCkxzV/2fzN33
8oxcIgdJ4iBWAcKov5ApzL0tYhwwfFLodb90eW1qP7cXccq+QNhbfosVqggCKKHI
/8WFSP+e8E2lwHmXAaoT4VwZOjKJ1NukVs9g+fQNtJxBhWGgWcXtot+lDD8Rj9Vq
ZcQD4VlhBA7mTCb31CzwdMDhYpHisQ3FKMExds/syb7P5jXHomK6qtOnNnqv85/h
saTKatLLNVlvbpUrFbmFowHynAw5MQI5KbiJ+5knFquRzgdBjcUM9R28cpk541BI
MhJHHp9bwP2ex6VRmjbwMm+EAofrPyfJ38KJ9lPZcnyy37nYgUE6MHpxwVp2fYft
inVvuSNsyHmHYg/i8m7z309VnzM72AitKyoIVIapD0TXTrdyBYnW7H5eWIs/4wfY
cjCJMYelxkqYfwYqeRvWp3KLCmndMmF3ZCpBi7YQdXZNQzf0EvnODLL9ZQ1G77gH
C31nyHZWLEVTFEPuJl5ziZU/GpwAvcJkzKKWaQj0bi8hmckj+UdVdvUXZjzalN81
aCUwDlkGZAWhRh9c9HpIlihww7WYDi52NScjrjDu3dhnAKfedfpuNNigJpiL9p3z
oGOCe3vzuHslQ0ot2+Dc9Kea6Gna0ru1dYhmH1WBu1N7UvJTkDhEFOO7tOgvTcYZ
xel8z8EWPoE2XyvJHRHhQ9tgOMbmRHXjGr2LB222ZbhWAq6CORryMh0TSJjP+Nyv
ZrJNRTKyn97xqPZcnIZt7aQQzflyC6FgD2mRa3hQgI+r4QpVJxKmrSsRsUl7B9rX
tIDF+GaPJ/TB44AqAHld0I185+n9viXA/cbyNB24QaBOo3Ax2BaYzbZ3lcRmuSwc
w5JxR9To7zPk5nIZtAneuu238rysJ2Rhyeds9RkF8RNAlRAmbq7GIIu/+YcmttSX
OJp1UnfxF1UutRHcgrm9wvUx9/QWr08uzKIh/73LW8m3CIj8pnXyioyuwPuVN5Dk
oLziTRF5fb4kDh/SH4n3s0gHLCm3IEl5AHROdD8B92zo989MuK6CSsYR3gCaO/Qc
JBJtyXru2KXwR7QjPq+196w3xMvP6k2L589Wk6G5jvzlDR9SD2FWH2vL1bWCYzXh
YKQAu9UBqNSr1CKTBN/Zq3A4Bk6Era4fYnxg5fpBBGm272qqDZIyjs6hl7h9Cxpv
1e9Z0hx/wqNy8Wje+0jD6VC1M5VLLpv9lRB7Oczgn03wO9V2jff7aZI6J7Zb/bvI
FzLoOl49+lcjSSA+iGMN9Zreq8FUcP7/PlE2XGyySxUdlpQCZCkHCYl/2/m53Ir/
Tw5Hy1fas4I9bRQS/Y1rdHJcdGSmv/3m790cvXp+FXxeF02pv4/UYluPUzqfcoiM
+3xfx5D5vTOi5BxWQzsqMc7u98a2s42mG8d6m5ppbg3K8ZpidIZN2rVyARJhfmHg
3fGu7q4LAQ3awgPGfjiJ9OovNPWipjH+RTgus1pQeXt5Ad8LkFVyylEH8m7YKboz
rVevWAsWOqGfsas8J6QrvbWmzqinOflHQJT1seGdVqWBWBdjJ+JXJPmtDuIeUM6/
gNHrseZw28ZemXPKfxt06sG9fWX/cMpnnpiNC+7N5s7SY3vrS2oKHnLMeRGQJnuR
oGs3qmzcauYxSyHkfMqDRtlaizMSkIDaNsQcLqt9N/j7tNpKC0U7nsB5I0SkvNTx
f6gu0P6uZ+kF9zMb0uPE4wEBJoTbmZoVopKaEhlINrfjqVLVxl/cGQoO8GityGHi
HVS0bA/iHrkV3NDZp8h1pL+DIffWaayyUZDfgPNMqgFfH7fUVyRLcqAVKjr9HVDU
pm8/NJwlsswnT7iLC7cnCBm3zj/QA4W2pAoZEiPKvkqGZP4OU50+K7mFYB4PXx9F
zLPxFdJmPzdF/4zzVzXl9dhaUUxKhwmKf25wwGCY4KGP+k7CcU0A3j2gBHz/nP5U
y0/EqOoseS7IbwHQ8kEf6RBtlD1lOOcdKYYnn21Ly6wAvKq92Vxr3fXONa2gcyp+
fvHD9+77kq8WE8F41QCiqhqtsuf8NryuZuS1fgZr1yy0lkJO873zEMi4B+VmB0qe
q9ksGNHvEFuBH1yPEcsFyoTl0sd01ava8u1OjpQQIgWNcDL/14zmr+cM7qJSomqK
WxSIBx0tbjCRH5DiUsfpoRZBUX6+hlvSeZyB8Uw0BT8SfWLD5MP0ruu3brgNM85R
fiV+kKjblXe6a3mteUmzJaWeoHkfh4eVeGmQsh3nSmzW9jRY86WBh9sA5MK2PTkE
TmYUqpcLMF9KI48RkY36w7RHZ2xKGPwpYOcTL4wVoVEonhDIxsJqxnpimmtibTNG
9zDBo2uoGwqcUfUMInJVDWwL2mz29LgArTxmXtsZoDhWBaB1kV6UvywROVXTjc9E
mFLJAanCK7ByQzSwVJhMrh3VFL2OCrL2kdI1dljd68sedt5kUDUpMQL91h81RQig
DXYiToNwV0AtR4oEW/ql4ZtGfUE8lbdbrqq9tZaegKlxawPzewr6S3jdaTI7vrkh
maYLZ8iNBunTgJrcdrbi1bCNDOxbSdeh6uPUm8ffImAg1oHfAThZCE/zVF8FrEYP
eZUqh0Lxk2nC15jKuRc1PMYEHaG8oltG56q+uFxfFPvXM/Ag88rxqPmCdhG87rvO
NERkZEHLhgJJw6sBr1Aj/zpeT1sXlsTxGcL18WYpGTk/UXO/qsDA+u+AAq6v1+5s
PtEnZ9SPM9L/hSruvKw8xvzg7ikBESWTrs/O+Il1YIFgUsSVDM5tOetak4gmEr/g
gJr3id2F4JF3UWkaBW8XPK2FmHCp06CfkanLZlBH/JSDkjHHBeYlq2jDCq5+lnJn
/srO4EWaQOFnberVD+LdJP8rvpYWTXVJKJnAhnqCc3fmuUnzPa85DcIP7HAjNgFx
CuWSFac51imIrhaqrRaG8HS0EhWb4ptj5z4vwJIat2e9sCUX90Yox/xHbkGufNWR
0jV0CqUIqFQDrtilBlk002VytchH7uldsfctWwjuqhTg7HTSuKQiHEfKe50kYzWj
JcdrvTTYALqeUvOZiD6rRdcL0m5xW6VZg6p/O0fKX3w0cRx432LIGXtTFnRfDTuL
O7t1eDBNGiry27wUwGnpI9BGymoQIzCmbI4/tg46N6VgqmDivgd6BRZ3b7aIf6G8
HDjaKFQONVLT0a0iwojhOMmpYznnLdi9LApL7gmGiJdJFCeovraPAZJmO3GhBuTx
5HASFbvbuRRHdw92+3Eq1vjVWfm0XBYvwx/Q4IMPjl6TW4RcsdNqcdO4TSd4c2dk
cFMg+BmDBUpfNtO/+3ff9a/YB+9lWk0qADGfbc0f8x9ZdCpNmanYPYm1YAfX1yov
mwHZlqUaaigwUBL6pUGIQWEIbyY6hlzx7VffYMwpwYZOaZi/Lt6mzdw7H4mK3/sR
2UQoCA6wk6GhOjbzA2wwLJxveQH6xjWG6NuHMQGGsBwyOk/hG3Fl9Ru1RZBvRe5O
EbC1L6fwEFq0kOx+s0vsMVLXWTZuFvxxnQTm6H0fkeD9FFV+uklYWi3IIX+WMIyI
WACbyY0twc/BfKywzqh5nMGTdK58DY9L7vFgXvQQTqfFNJneKcCE71T69qJdKxva
FxeY6AwqAzGIN1MPeU15iT4FG40p4lJU0+38F3Isc5QcPXhWFRs5s8vUH1PfNut2
rYiIlnQhhtnZ7Z34VJiViC3Y8TjSm5tDliiMjM/+f1T18Ee/Mo/4+ArMGYuZi0vQ
N3B1ONxIo4bDxnmbHvzP2hGMZetrgLvKP/dc60pt6s6oLyg85S5dmqVkj2eKFSLt
CQPzs5XvJZ4J7bzKaeYl6J3wvJRExg/ARqgcZiY5gKa7hHa/YqKqqlPa2R1ktwup
2phy5bwcqqXc5EGxtigELaOeLo2kqiYNpHKt5WQqgrV59VhASfYzzMbLYkN8YOEs
9T+fu8YlJBv8cG3I5pHshd8tZlcUuQaOYkNhF2uVJoIXEJqZnKWt3VYCnK/JGLCQ
VLsEtrzlFWk01A2rUlZGdTreDokn8go3qAFboEoMaDxXOKZCIsdBALaG3SKIKstw
T/Uo+Qees1XbRKFzjXHefWlMDAfiLhxzgxwmOPDjmYdYmuKY6MbWyJEGVnrDj0oU
WnRvJYV07w5Gzt6o8/IU5K5Q/hw9OTYcvHDZ41i8xAcgCov33xtH6o2JkqNGia2l
KrnYbKXWUwkyvNBqAvRoaLdgsFx395oZ/8mtt6TbTSNJ65QRUIBsFAnseEgQZl9n
pstIF7g6VhENXeKoKxDBEifM7Z2sMOPp6v1161ALaWZhgDk53AeqY3Vr4BVMKSYV
7HIL+H5BzSAHKcjHs3aypHkbmfe0ODRr4NeNDfVHA6RyEmyHPeQBJhddS8dqArzg
kz375TfLvfWbTKTJIuNeKuFRmj9q0G0noVFkYOBZVyOmo3A9V1RgH+v5318nS1FD
x4vcq+11dnriProes/xlu1n5icFgx5gzf1CuV8HEtx5NkW5CNxzMZmpX5vd+A6pZ
PCU7T+Q4XYVL3YiAnVUcyLvnwk+RpV3SmJHKWBvfiQQFI1W3DVqAnaneamD//xsm
t0VFJ871BwOlXRjHx6IK4XC82Fd7HbJ2aValirx8FZsTdJt+j6UaxpL8Voa8BuG8
Qmis9nkcR/zkWAa5OGTqih7DYIzAvhRC6v1ZYDtSFMfJOdrveDsV4eBiGbY3m8q0
f9/e3nbiSWsqx+sR+3K5f0FCxFV8sdsGhAO/YVDVQB0ghqVWc0cj+Ie7X0PjrV4I
SCUQl2J9/6mMABkMqb6tWhQ4PDmFHxV/DxI1v29t45Vhb26hIyPyw9IanjvUY/g6
ypnNoncZy5dQQIrEM2+gl9U6P16V7uXctreeOo//raaceCBcGz5/fKbky+t96Rhs
9RUuqFqIq+y+uDIXgwRNG01EbnjfqVJwdUZiY6/WkOnvwe2hWlkAFBb07wiemhDg
uEe10W5s7vanp0HL78H3VyOC2PHSQJ76pVR2ipFnWbipSj+j5hvjQIVs/BA1VcYG
HFg6QV8Gy/nR6WEq4pkiQlytHB4REMak7BZlw2wzWYjLLJnmE5EbnCP7eBeG13FS
U6c7SD8babFbYKO5VEH1jdIuOoE13HGwFHj9v6iJ5awY0+KszlBLqTt5NstuEWPd
X2UAFpnm2xCqViNYbMxGEA==
`protect END_PROTECTED
