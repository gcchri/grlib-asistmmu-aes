`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdh23xJh5uDPh76yZ4FFQ2rFORGlFV4vFLGV5SP3xHhyr1xgyBw2KC6m5NjIG+ob
iG68xIqhR+oQJzoTms7BEe00YYEy+gnFxpGKkn5I0+bVw1gTSDcHRbOPvK/NzyCI
iqkpuMZV9Ps7DPczkJoPdJR9S5/EaHju+rqj3woIUk+0ASP83BJnTBtUgVncgumX
OL45HyTTpl9Pui0jozMOldcSWBvJkAiUZdLYzgG5/z9iRMRQ9a6qf5FGnWUuIfKL
yKnKsHCIxOgFyznyrmHiP7sPYQzTe1/I0LgYrZLZEM75VZtsg11fZ6OwG1CGH+lY
QePtQJHVllW1NLuoRtELZ3yhGZyOXlDWSWCoyODgjcNuNH4cg3QV4WQ77QWfdLCU
eh5498CTXo/0UEmG8ivlovdFlcRG4IG/TJjUUuopYfvJyiG1ADdUdDmfdo5JdM0M
tlv5JtY8OV8ycpuJTwvcC9b7Ze9HcB4iRgwKSQpKD9SB7evEiMyATMmAATKB0DTA
HAQDMHlifCGekEbWFdEE3mS0dP1QUt67Ji/dSqYhfuGaO6DZFtV7ZDbdBUU7AeQS
+pHYlW61HJnAyD7xwnQlTUp/9InY5+DTO0fb3bBZ2JD7Fs8YTTdF/HPfEYFfPKxN
mojFJFIvkQt+wDQ9lgWFtCtMxOyS1/y5pWnLB0z8D2y4D33HV0uUVjSISC7iMJVS
AiuKURUYjBWDzyHJT2pz0eiwuoUH/eqkYQuaO8K/JVJ9Iu6NJNwufINx7Q9UkBAx
5ynsbQtMjw02tWx7bvH2OSyKxpiPefm66KynnhIKL2DfM5N6p78VcuE5S0kpdAxO
o5RuII3BML6gHsIaILxHJHkBIVVpdY8cBoTrLSKYReohd/K+rmCicpkKhQmf4nph
+Pt9o/xQ1GOxx/87clzqwEyKy+gSGynlNuiyes22wAcG52/vykWov9eSQN3lB0IE
edso68AVQHfmwKEBtEoI+y+uqgJM0ZyCLUF2W1OkV2fsXZYJkqHf3Ib6GoG1hgZd
IzJ71/WQoL2Cgigzof5v8T9Ai1XtVpfWlbwH/bNbqiVWF4RFTCCtbsJWr/q/YfsF
1Yb0KpgUyfrmJvOz2GHDSAXn9fHuZeW9QLRcuZcg7C3YD0PeDzhaAm8Rw7j+H4MY
zAYCBSKzrYyfKPlGgmWcvzc+oR84tkDip03RAouQWe6To1ZKc4NcJS3VyyEzuID0
S86UtUocb5yDsRjmwn5sOFiiIjjD33uTmTMM9Xmn6R2lBdMZMlLbWh7L4pvu0o1o
y1M0MRPXG9Tfkq2alW+G811oRVpuqY2KAX6RGflW9MIlx+p5ZKqgUZuymJmgoZxp
7xWwg9kkH6lL2L84WA6u28SY94+AETF2PByVWnvpwbxeK8AaHzszzhVzrk7GCwa6
nvNivaOg1+oUiRzu6E661pb5zcj+nyUrik55hH3dNwM/Hga6HhWVs2VydWVYYzbc
qvQAD/m0hR4fclOa6ff3F2zr0TiQzONY5XBXnuZD1Zl0A8E56Sct8WF9Kfr0zLiQ
uzZbmHsYMG8LMEnrWH1yGmaCsYYxqB9HwoU+laceC1VBdhcm3XGzwIq6p3JlauOu
h9Yj8GOgJYFnphfKs6dQ/x4vMA3ecdiWp2NEUNMEgcX8In8mAu6wM67dZFdj4yj8
7Q3S60ywTknx6eW0xIOlGlzvl0r8WtpueEPbIUnZH1OXZf7l5yx5w9xDudis5JK/
5oxWwGpEp+0Y6OTr18IenM84Xl+M5St9MG/8W64JQDGuEkQh8+yoEsPIbmDVlyNQ
stN2k4InKWoXjmAXrdeqSrrPHqD6Zem5Pndw3+TmEH4p6aN0TksbftTfyrZu7rFV
IFlNY4jkMwP3CTNXoNM3jEdVs9AHQfCcr76Tp/QtpKtU4L9nxMt1KXGCak99DOcv
Bb09srQyoRo9xfDR/nurtZy8JA9cMB/7kXpP3DwL019wJzKaNXSnm+AhZzWtEHLi
E17liWwHW9j5MlvlKb9qUnTSEnr7WhB4K6x/wuJaWCrB/ebxSC9hFptCaY54IFLA
P7QJ26tIqLGc/aZ9+bG9GzSTFDrzVckexqdpcGFb5VHvtiHl/jaMJMP133L2VkuL
5pYLW5vyUkfFXelMTTuX78c/W8H1b3cz0X4IM8t9LRZVzC7DQ29wQS5J2eWN1vm0
3Ks8/SE+JrLSnix5OdE2cKzTJ6Uq72tVxKSmLQTLy54wseDFBFVT/IiEp3SmslPA
XrSvKb8aeecqoSLLSUXLmMBChc1fd1hce9DDGX6BPc11bHaAF9yqihKHDbtBCRdN
Nha/KH1/BMoCKjomS0mMiRZ0W42rmxpYJHJHvX2B2XiTUv5bPVbTMcby9Q+TfuKg
eE6yseJCrEZcm/NZAhXw5L2N2edag/HBLtRony/wd+pMiXWMt+vpV+b+W2ilMoRX
FNY25f1t5C4gnkgTs8zY9B6nwbwGCROMbbyNnyLELQcp7is7BdFk7e+eDBCjMxzo
LrQtoOb+upiUPVRP/lYwO3Ofo2SKnuxx3RpJFh7RrpIarLFn6pnDPqS88i8RzoGc
q95EfSvZi2yrYDMC41eoTaDOVMc25kuvC5m9bI+w/c9dj9YiUEm5VB/mqA969qPe
fGc6gPTa05b/XCr836vWn3MywgVo2HKwuGJLJd8goF9h68KT2VDu0VZoAWz/airX
MAxFR0D3SnCcAfjtrJWjeu6OCupQ8Z/YxXNqwaPQuRlEKPw8e4QFtUPg/53ao+Wq
FUdm+ldHGZP5WZIXELpZ8ny2TODV7Xus5tWnR9rEl08Hjlx0nEaZMtC+MfbMPCOl
tqCFmJK8o6C8AONKydYxhFo725WYFrrWiC8r6pGRRGi6/5Z7CXl39e+uqQ0i3kiA
9KCQD7J/kMB6C95GliotHyu4zEK5EU8csJYQKb15CxFO253NPSXnacepLo9e2Yla
pRNdjGaY/MqK3oAkjxUUBu2C4LeyQPghpLznTNPy+tHMpCnEcavdNbx6nZ0pOqSz
QoEZpkN/dRUi2ImTWRT3sXkCjb60ngWnRCOMLcOrAZ4dPWMm3WV60zJhUqzU6b+U
hYRbI3jODmeS7b9en+kpLZJ3I2kC648ze5+niBmutKAmbGr0ZfpqBJAHZELHO3xh
kWV2UFLfGOy2ZZ/9EtQ9OVxAvhF65sJjxv7iNXk4fPdLzlOfph/JllsQIpsFKf8n
wGWOMpQxY95z3CfoGEnCveXk+nJcNvS+Wv/+iUh/0vczjbUPvm+Pfos0IXmUl3wp
AuI+q9fgg1sbKzk1nGRw3v9BNYL6Q8OoOK3a8z5K5UxThkuD8AfuqZwxg4yw8YBJ
HBEHgp4t5WVJ1O7cnm+FvDDwjtAfhzaGMquTfxoi7NZxhfHJwCAh7yKO/ZyWMMxS
LeWniCRxa5qbateOpeLTnP7kyy7Gy81oERhy+Cg0/S5fyn5JybLaYII5wUXVa/cn
0+RyeeD+RzohRyXxb8DLra6VsMopLV5/ohfZvZFjea7IL2lbJsI0JZ8csHUfeOWj
CPbHrNo2pX2AgVPYplUMfd8/e2tIwTcr5rAqAaKM3852rGcD+3UV8qhodf19xsvW
7HugKT4NHBNZ0U8zl1/IY8hpCe+Vzr9u2Z0xjya6+5ZBbIR6/q7juU3UvnIJmA0Z
KrZbDbvAIl9Q8E2JF4jQCN2a5GgC6oCry+YllD2kY2jgAGB+437Pjb3BvES5kVC+
xzeTniQKQRckS5C2zsfWFxLUu7gvSj3P1Ety1ossKYtxunlinasjZLbHbQqZKPPs
nk8KnRanVV0IWHv9JlCNLX9PMX44SFZka9ox7XxSEGnjOgyBgFNLlyz0AX+wDQ8Z
VHeg+TgyMxPOUB4Ned8WJ6AKpg2hN7gyLC78gDRT4AnQdcZHWhk4UrTYp4P329a1
pdUVFnviHzy51dY6C14K1QD6m4/KSb56kUCF2WVDhyxQbwZQRuLJC2jAYfcqmkmE
kps8sdb+9CF5pd3yYy+hfZPtOd3e3oPoxz5ljz5iOnQJew0TUiPvOrvr7KoJdRZo
lm3Y+OF9jUEZGsxiGhjevwY8etzwv8i/34D+u4DRzr2Lc259k2BxirUhHw0WAkH1
1ynM/f1q++tNHToiqh4RjfiBxhxIzwaS25IDNfwz25MQpsUZG6yIO/3c7V0S4uUD
jIzHzAMXm+DeauWjHjacD8aq66qauxRHTczPpClTMZDvFrzG52YntJv5Ph1eLzjI
dxDyRG30wSjC6HhohebFwXzwa05y89FgnS11amSfB6qm1bJMQhzd7yzBTrKlSuEm
QWEMabhznX2U6ItSvgQepoNaUU+I4/A0NT4a70+b/djtbRaGfwaRBMY2b+mkZ4C3
a31V2ckL7de50LeAeItQBe4I1kZEPKlSZ627UG08DFaW+Jm9yssrJyy+Muq0PvG2
TkXUP8RKMq9qgDCClcbknFgA00DBLfhqFLTcIH+ijPzbWTD//EOST1kJRhZZetFe
glC2PDTfe6CARBBQiWD7JHP+eC2ohVgZfAqb9DYEi/8ISNQXn0O4Jh57YiVZnUSw
jdFv5htS8zymjKZVt1cW8lTije5WrRmdQe0BW9gpkx4fKB2v75d9CkcIuL/EMe5s
zU6bfW3/Zw/K4hEnkKm5+wkpyHJxwgRdgkKiq1hOv8KGaEEcHEWcrZKYWgtO8P79
CVjfwpG22/sGagjTL6UopGtwFKhb3O98aIpp0uSk5gJUpSCl/VE16zDFHCDEbBXD
7CK5qa2o2ljhq3aGbZkPhMcw8bpJfrTTqvFfKrKls8aihOuqw+xxbatPN31RNvRN
AUbKFrCSX4HvAWUXt0j+yFDm3MzaG32ATRP4U/Bgn1lo9ypZYUEXwMqgVRibbqvK
g8/AKPy9pp2YcTbI8Mnqbe3Mt2GLtzXuHAMFTc24dUJuGia1yvcsONEr919KHRHY
NiMFlVTJxpRkyCaYfYK1nspEBP6jmQ5L60k/oRMhmcYMmRp3gZ5rGWQ7HaTqbsBX
v61U01hh4fFCS5bap3WVWNsDF5xtoX/KIvKWDnivF5bYvP6lTRzfBjTz2/9pj2M8
oan8NDA9Dkj+k77zI0KMS00kmqCrRNDU9LuIonJ6KaDZtXJFsLis+oNiJfqSOpdS
4gZ6Ch0OuwZsK+fmOGYOa0BiWTvt6yET1yFWU5YM6O7KcN7c61LbdduX7627T3TF
ajWsL9w/1gFLz2KjL9ToGZ9teSGxs7XX2yRTejudcyyHBu/Sn+TOcadUuPpt1rid
oXomOgA5QQ9DwRUwB3l5GXKG0lvExgpkiwFxtoBnrSZ0dxRF99jRD0FDMn39JGRO
RC7c5EnufQgJKOrxzqpVvckdtjDtzoDgzIen1ICwNFHwnXeUN2grcaMSXcnlFYVo
c85RGBgo6VjToZXCCP3PicmPixP/d6MtplJ2tOcqeq7MAQl5wHXphH4xiZMB3WTD
Qpw4+2Gf+8oaRCwhiUituYWzB4tPjnzM+VMeUgfMKW+wq06tk3zALhd6MG/Pp222
sMa0pLyhs/+bWlp3f12+ZhjKFKqzOShd7S0nqcbJwLlacTi2mBPmRt4ATFdNFlu3
5nrhDs7EerGidy3OOP8oWlKUZgQRMgvUY9qxlQJnbFU14Nb5ipk9jxYNV6pWppNn
2oUasj8T/4tmTvs58lt20ab+vjCCyYVVV2QOMfMFDEqOJr1cbIOHrDJh55+N1rIs
okMB49sFnAt2/S2CPP7xWfRkn22z9rxibs8jOqkRbInPUHFW4K3DO+7iye9ilY0z
SxjiNrZDqX6Sz3e4yoNhPOdFVzz0+by78KxioOPmkI8LkVTOg/2JK7DXXTIkjyC5
msBXAEz3XYAlSD2HWEzSn4azZtWZ7rJQ3gv4weIlNvI3bgSS1bjExCTzc7049Ki1
FKc33bYbnYr50n04lYtspdmLSuH130AsbC787oKMRoDr2UDpVCl7nC6W/coLCUg5
8zbPSxv/XJSZJXQAUGV93RL7m+itwgO13CvLhdBUMfJfsSJNOw+XVZiu5UCBECFq
qJVOjCeSfmgBxh+TAXJi7jl5S+ZmKbpI79TUq98r4tsotFDftdu1FLv7eaWJ6MHh
R7mhOEkeQWgCa2QSvwAuW2Hg5PbkHH6gwa8QzkUtSpM+1s5cJo7zDGU5bHl8gHb5
RyniNNYC0hgaDSxZ/JwIwcxfS0EUzK14eTI6MyGCLaVGL08l33cbZ/Je86qqwPc2
Kl0TBGwi0aWEwmtGBpmMhUhhGdJAsoUM7ryDlZhnxtO5HLFepZ3CyqbU9DI40NDv
iT2vIBmQencwdDObr8aLfFrW+KtxYe2eqaLPIrBRw1S6V/5JL2MQN2rHldMGXs3c
`protect END_PROTECTED
