`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3eFUHSriSSQIWw7M2MpCHmRzKNoEF6WGgH2YFL8ogdGOatxKdCislzgB4m5iKN0
GRw4ZV7B2CtsKGVplVjWOiIeKKlZgMWAOKtdQPKSGw/ye33vPr2nSkfHmMBcZsa0
HWuxIHf8xAgWRBgSkGN0IwM/O7JHEZzdigsnuN/ktj32qeo8CjMNXRS77v/exQER
1S5lXqsU9ewSAY/reKiPg7psXXIhblRveB/fW2bGJqYRU88fQ/D3X8qEdNhpRor3
biFGSr2+5mPfaXXpTZjnDsfwrsLsnihqlmvxsrQ9RuYPAPjY05/HfUhDOJ2XL1F6
7Ww2XuLCPxePJ+O7sjzh8nrpvL3fwoYRpqmqYECrY4hJ7hxaCbyUUY4FQna7OiPr
xW9RP6sKjjWsLwa1Vm2rphiVf+BjPaEJ6nI0JRV/gBqbOe4J6HsKN482nZn15/Fu
2QeJFGW3sZ4Kt6q5LjqlnkFjZAyB1VZcUvREvA+dFaiXV5HinASSuffMlAl8IMho
`protect END_PROTECTED
