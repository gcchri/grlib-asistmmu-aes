`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bjuR2TmF3O5IF/VFBWC5xZRCx0KabwWX1dlaT6xrdBTNlIRYPBcCFSY8bZdxtiG/
kVEAvinczdyFWdrfR9VpJjmxOfVBPsC118rCuDDsf4CGkbwVFidqjeFPujRlOe3L
QgUM5hxiZ4IkYyshARxu62oV3RF4ojuyjukiRMKhxKSvsTE1lLqmMVXsa4/oeIjS
BxtVBh6DW5qcpdFlHZHSJr/RRxw3CQUT5u+qwS+GqpjgIdgXL3TDS4alyhJ0yU62
Qu3Y1OxC+P1ZC8Se6MC++AiUyyWeQ5ttvlsrRPp4zwuMPTiKNKNXmFbvyb+cov38
gzPiz+9hH46wsdjBMWERC6AxHkpQwI2JDjuFDN4baDGqRCancjN+GRaiOUQccqG7
mo9CLuKpt9yXbdK578IFIFRNDicrEjGxV4mWa98FCf6cznJGq4t0RJULLvz5ovFs
6fU2W1E82NjhmYGR+i1GwSo+Sy7qAUAtHy81cYWigaZ3W/xOhz79PjJlXdiQd7Mm
0nRGdWAmt7OnCD+DnDj5jstN6jvswuVQQ4gLGd4i7jbokiRVWTegN9y3hSqIPHKG
SWK7DFgDI+js0W8qDlnwl3/bnF/GUipbk8Wi5PWWFJHJ+3vMxLuPFi8RC/W3EPqn
edjc89poUw/AIsG8LI1Jw9PENGnjzGTZtd45RXWSA4s0Ml6EL71dPq31q3TwokHj
FHxA2imi4kpRdnmvfbCa7CcaESpYo9iOL9x3UqXApZpR2+r/5E4jVlXQApTUTlXu
hFENHGqRPmjBH5Ulcx9u6Mttdx1EF27MXTNBBATC+HtIUA72nNy41Y6v43bItyL1
`protect END_PROTECTED
