`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ThXPxq770Phni0ZX96Hv6hXOZceiQWpSy3KuOhWKZfM2wWbpYVA8id8PU6b3F62y
tZ0LHnk9dul07KQBd7lIeYl/OBZpQ3vPL20z6kCugWtJjyOxtdDg/01BB3harGQY
kvBgxoaz+cMb4Wh+sCHCKqtLKBPc6COZh0O/52xd+z/GXMmAEj8ED8PkAw3iuvmh
l3sc7Jf+iaLVD3bqyznx4Bi1bhLEGNwZMZFJzxAwQ74blEmHDlBwrMNj9pThRYiV
dHWn+wQiwOoh+8DEOvurcFYivaDucATeixaAGO1C0BFvd509d3YvRB58M8fvH+JZ
W2e1sgYkk8WjPh6aNzcVqwiucji+3wA4ymEtG98S/Ulwd8RulR1wll4SJcVR4GV0
Z/dxbOqR0SJUX5jW9UHsIJ+0tHxd/iyKAdjhHuEYAUJBKpFPzGpzDLOnCNb/aiLu
vS6U31Xmx6kbub7TfOLyAsiEZSgIcYHhezuGCKx8jhkUVJ8P37QO1oQtm/eR1vNo
W8PifkvtipKo2NAhGkMx53z8fL8TDkTY1XgXOxuFQYqJxWV6TI6sIXO7ysbYXkma
W2O32DBQmNeeriCPGTaAx3TWsDT9Y7P35Ibo88Dqcme/OnwmJgVfdupyYZfHLSm4
WLIbubtHLBCDM53idyZk2A==
`protect END_PROTECTED
