`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jq4M39X+nNmd8vFG5sEZik9ifmiN8FsFCi2s62M8fwUvxvu8xo0P3JASuEakSiPA
nokRv32xraUoansv9JKkEF6rSSsCHVCjONKJUbg7lmNJ5wJM8mkLqLWio5QmS9m4
N+D3uLOkWPlAqEZmYxTZEDOATc5druGZpueaEPqqh25oyNKYIR7oWfGpu/o6blDj
wAfWbo2GMa7Q7vRrgeBiOXVLlK145sW7NbHdMJLe5VYU6Evm//vaKvY/tF17MNCU
2xZ/Q/daehghSjMle17O4vdX5UiE32v+Az34RZh0B/eboFqg+CymFXm0jvHpUfw/
hcDGs8S77vjk07CoKt9HcNJSrV4CVBdtsIcXclKcIwjp7EQq3aw71adkaDvhnqTP
VPpQMm0irWfEpYESpwo1OzKPpy68G0XMFme6FQvwmhg=
`protect END_PROTECTED
