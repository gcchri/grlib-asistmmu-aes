`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wkP5jWKWYMVj1LeOv1uFvBRp82Rkr4GKr6KGMa+LF54nVGjJgpxvpoCzaQaj0FwO
LIUEqKJcthvZ7FHwuxXHlxktLBYmRyqWy17+0kHvRsBTb72JC7gZhYhpGAIeC3Rv
nLMFXhGsZl8UNW1BvaofNdhTj91Zo6uj3N4Nz/V38N4BVfqNA6ThXaLUuxnPIck4
1OiqGJp9d64zvAA6hpheFQxSfnplbEsiMZmjoX0zFNWePJjGtdKFccAJ64VPe7+x
qkV4SxzEu7fZopGXCfnN/p2DLRMYEiah3jjQ75PGG4+sYk29wmVwR4Zzmw1wcYIG
Bl6R8nYJc1vFkABHbpu1xQnCKr5NNsWNsZNbiO26W7E0Q/5AAkjqE+M3STDONzpI
lQleutDce73FZ6GjMDqOAEvoUNXGMwJx5owWlA0eKMd7S5R7UqjIQDRfSbcjgX2p
`protect END_PROTECTED
