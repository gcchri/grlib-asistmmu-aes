`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d5ZbgfPtm6pTaWOWmoWtCscUiY2kb0ZvV5g+92s2wQDOtWGbYZJfL7glQEKfCpE4
132TcxMol6zObKnHaI/mV1LPbIZcgLVKxjOUaXnvQjeIwJB6qVz2FjTtbxEivEpX
Rh+n7RgCK5Rff1M8207MwqRNKwSk/T+SkTdmYeU9+w9SUbEA1yZFvV1Oa7Y7P6t/
y4H4SEIngz4FF++vPZW8kmckIk0TWK/VlsHjoQhmhLmqluXU+64o1M2mM2zIVayN
PWKfZbwAg9OHN5M1y+3DXpAkj0mpwLw1qt6YqAdMD0k2GK8OHbwcqgX2WPCKlLVc
SZ8WhIj5494gb4NKdCJaoxH70LddowRvUbPg+IIyIhljxyJeaQ2YnaC103HCDzM2
xXe7T1UAhVUGJuRe5o8gstaMbNeszOeHcLcPuTgDp+7UDZ6HAu+z5qFW8KyY9enw
RF+iJFIzk+2tj+CmyNqh/RR8s5V1qzXToBAnJU5LVAm6X2Gj6NZUM7xStyUQ6j5J
xdnqrkFzvtWsFFiojs38g5yUsTdTqnymvlBDu5aKk+UVlnaEBgK9TimQPnojQVG9
OJd2VBMRHhPWrr8EpiQqF760mQpl9ygr7q6KP1eAJ7jZb0rXqoEfHU/VfO9tm/QE
uEwzx8/CuSZDvPtKRolfSQ==
`protect END_PROTECTED
