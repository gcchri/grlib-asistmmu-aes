`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b9DYoMdhG1fJpRfjJpwpVVVmm3/vL8gUA/OvPI4qtvRxsyHM2Jc3AhV5SpcvOn76
XNFt6xGv58tU6JF6cVfYPSBQvnMvifGW345354Xq85+LSGXw92n5GgrjkV8n2sdV
TuLZCwvgq8faoqBsEXYeQnOVfCbsh9CU/nQgIQzI3QlCVkS92UT1Z/3/ACD0Q8YE
4gxr1WHFgLIoMht/F/5L+jIGElIOzHuhbbZu/v5RIoW6DjBVGzm9UCnf7Pf2AWa4
fLRQJr+bDBT6wK1ryElocjqop4TONWBjBtboRlvnCEHWXQQMvCrHO0b88aJ4opf7
zBGW5qFH6aJHo+CBrAny4rBKYG+LFCQOJlysguZXm1ke8UMwgmLQSV1wZYtx3uJF
8CE2jYWl2RX0iDYargQkNsbwk9Tru7fEt2BJIMcxJc5EBnp6vn7AY1aEeoEXYXoV
90+MDVB3MsKb+u5loT59DXhYCHBuzB+/homuErjAMnB51hhDD8MYb4IYscsKTyN6
lQeYEBW9g+wwSmzVAgESzY+TUZ1RIPsz+rNL7qEwiDfCjTjIMR49MqtNLwQgDHMM
VEbZoWtRjzVu+mMyUwok9pH7CpuaejnpATyX5FVLFSNFzwpZst8DNNbPvX6Zz+7f
kZPhQRGLl8W13oZA4OkN4d8o8stSYRAeUKXTf2+5YRh+D3IyGs975nHBr1PsqFgX
i3GYimxews4ehVPOMQU8Yav+8k7bb/iR0LrJLRmtVHscdogfy5kmEMHD+Yi8XEMp
EZz82VDsv0t1CZE5wLf4R3v7A3rioMBmCK/smGAjDaTIebuZKvoTw//BBAYJ2nx1
jih0Lrwb2umN/U+NJeIIKvm/65PeUaxGpNs/pvvSX2En5HiBZCZmGZTEjc5y0ZPL
qSnPlwf+k0T+rME+DC2LL4PH64kOjmDy9fzkKsMtp8894xQF8V8+oVomHUxD+hag
9L/qTg8r0MQjld6NxKnre0SERPocW54I4M7aD4LIfoSKzeTsvtsBzf/hFCmC/M5T
sxdVtLofN471Xb/IabM8rSkfQcSolLkudN5ONN5BbQ9edItLRHbpPiH1Zzxy2N8x
0jkhPCJs/wTsjmIhBUAtc7BekV2MX5pP/vZsOMyy+WOTBBP3aTpfHu+qpeRd2dM0
bxjsM9W+4+zhaU6xMEkGI7xIdwjsiozhSKXut6Q2Qhdq1ttl87GId/MXB9EP5f1S
ucrKDVe0nkTzSIQVOtHjqP0qctBm8c/915Ozb0v/DJ+IrUG/vYfBRyH+DfYJ1Yni
mWZC6LXi5uaaog0YWy8/gQ7W13IUQ/wDyur28C+Y37ZykjszNyrWLH6ycxhCc/4f
8dwKOSm7zoJxS4afJWXYqaPDmIWVr0+9x+InBZxJS5b+Rr89MMpUDl2Zl9iiI6wv
r2u4hs8xH9smmc4t4MWq+DQKpId7mxEZ6m26/vvjYSrwToHkDRpL0x2b0FT80zE0
xl4cV+ZVEL89DbMRKX9CwKv+TQPkgV4FF7YtoMc9KVa194K/Zf++EnPaqu73qbPN
D936eFM+E2hpFXs4fq1q0meD1jfnG7Ubfjobg5UHEeydZYysG16q+j1V3Ihm0qv6
1QJVVOdgiPkbqTQg4JEDfTDnjKWlEEytIv6O+YV2dzm1eQqbwD01P4pdn+Ejw3A1
S3pnWIlrdFt2E34NEDQ8A6jzUMj2skUezohDvXQPlq8MBeSI+R84+LKrKtIubyL9
U2iaO28bQWtjMrGqReIMUZxNLsaM+dr8rcDop6+/yFzGPHEpZSJm8687dFN9c8d5
94l0irvqS/u3bjqFMyviOjD+PEONlrq3QhaBHXtIy4NpxK4At9sJyM8gFCmMrn/N
9LkdzC1wP2pGIikBAkbt6b/HIza1PcoLlaX5U30YZnT1EQygtfy/8iqah9TfYkUh
caghC03oNs4H/u1MJpshw955SXZtWHiNoTpG6rguoit0OHUUiLQbcAqsOBGl5Nl5
xBokjUGyxjUZl4Zveh3rInpjugTXhO0Sxix8LuIRNp/3YEEjeFtKtEascH5VCbyh
PwMIgcJ/5p6SH+wHVZSnzUi5lQW27ymaJFvPFErG0eFLdW7j7ODVxs2p1NOpb5q7
Y4b6wK7h4ncWehktHtEj0Koothl6HSnvH7IRAwS8w9O5x0QxVJ1cGBsA7YQuyno/
+f427ZZAfFMofngwKbKpPnzpTdgS8zvo+EZxRwwAIefxaJNDzzU8FmX1ECmosgK3
gg58P+MiM0qxgb6v9amtoL146kI9W5tYDAfM1illsY+c2Wc7DRIi7phl70nDGd1h
8hoLr5FxU7QDmu5rAyiS6eaiicQhgLqnVjW7OqZ1G6Qcz/gOw1HM4wbQrLepe88F
IHvdI7oZYbR7g8QD49QfJG4XUnUeYjHlSiPyeUHSn0MDICE7YQV+rTMoO58kjKWH
VsRJYtmgBnRhcWdLFQnU08DgvZ2unUj0vtEnL4UutWZqrEj6eGc9j/RtPj86O77G
/l9tfE7CgKZrNbD17XZCl459kzPaFMfSAuabtS4pLrrTOwC+hnAqu9FpBdxQr1Uo
D38g/CgYozjp7xHxjeqhKUSG5Vswq6/wxWw38OCXcnj8/6Af8REN37mj5B99mZT9
S4vidbEizIdPN/nF2Z9Dv3zFWDCfZ/ArEUNn0jozdE5x+HLhoTdgRt9XQE27UjZM
QNDkpY+IqpocpvqqMS48R2Kj1D9KCm28kTGpRFGp3QIld26wac7LtOUzEeqW5ncM
6HQ4U6JNHY0Cy1JXBH2u2WpiqHYOorFtWPKqx2ltZTXSS1IRsyWg/wtJLrdHxU4r
D1ugJyvT7xDS+F/I0eWdsThQIhLixpyB/S1nnmbxlxsUZ8nZ/IZMGuVoDoKH3i4M
23ABOSkJ2DK0pw49QfOWcVTPLa+9GYN+nuYhmwj9GZOtYxMdoK//VVPEPpY9YRl3
FlJUN8Gce8P9lxmh3BW9Q1a/KSLWvM/1ulqpT71sS6Pb2wONx6QC8SjKlFuOuwFQ
2uhuObUf6jXpHFCmxq8YgscZKmwSfxrHvJHmTPu0BOqdqjLqYqLQkCcnjwltKJJx
JsALIDmpSIv78U4YEM6tLMjFr51vReS85SEbOPKdKjphyvqyW8a9uXqTPcxsTEFm
qtWGC+6iE3GGJosXX4OThAhqcxVSeK45YPNtVgE51GiKNFbchcn7ymyy0lTMXDKN
t3M11dEAPEmLtcJVvPppf69GwKVA9j88BhnsxDsmmCzdpvNb5MskjjNKbChcFlKt
OOQVtOKMTifQTda+NOw82//10NhBONjjN8N4KVV2IwC//aJyeMPbfPgQrgwB0src
HLACDDjByvaiH4I3lrWWpeIxDRmxBxMiTRavNamL/OlzLmaguvCMfDPdfOQsaMKi
qcDtRkqmU6qiv9hRgUckEaF/Lluk9tnyqFxqikXU8IJzEX9O7f/kMUh9XhSV2jQz
P4aPiRYV5OZgzTzdJgpGHDRTZpobVCJOitbX07b2qBKVzsSN/nuwnlX+TpBgnF50
2GDtR2thKd3mVwJKfXelgmFGJpsC5YGfNo/YfgD67F14YRsw/o1t121cRCQ5arAg
4/qVW7Vrzucp9epOxRBLc1JI1OwYGzPKuvYOFExLIk7TAOly9tFtWf0MP/0JV6wg
`protect END_PROTECTED
