`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5maCsDlx9zxMfrjU7I1yn1ngHOFzXiT+1MpAewCKyce+W4+Fl0gG359g490d9Cxw
gK6dFZg9vaTgM1e7TF+Pf1VqQVB5Po1VPw3En9PS8fj4bTRn1aQIKMMMXnjJihui
GM24841KlpzDOdTxl37zk3fmMxu/+N1xKarOQg4wXS7KY3wrw1RkrbL4yPrh5c00
y32tCq3ksDoR0jSr7+CDj7bAme2ajBWQK8+TA20wnhyaZM+KWsU8L1llX/KkM2yJ
5EYsw1UrL1z7MB+Rtrv9P9ezih1QYJJNJZvGVTg7nU0mX19bMpLolk6Xdaer4e/f
bnJbFo4LoZuYY/eP+3J8LOf4rWKIR1jdCGX87tgYYiXpTE7harVEdHJu4uchCxxX
qzeYfDNrZEZNcjZlsdwgasiBjilwgewzkvPZN0D+lsfXZ2Y0EceIrJtyoTkr1py0
HSSpiQg9438WC5/AvVbzrbo4Ra0lNoS2m0tPe9gdRvNB5vt1g2j5z/AzG0jmp9pl
0TE4QyTlbxNydfRvY1i/smKXuYJ46WMxN6RDIQJCVyaVCj5XnJPLBp/zUGxo0UKd
ruadaJt1QkD3fj2w+DIdILDLw2NMiMmRPENZsjpB2EIn5OZEeu7gFZKKDgOqaxIX
/IU4Mexzz3pChg97V5ZRM/2+WjhWQWZj4LTJmKPN8s7FMYextVQnu+d0hZ0wDQqC
RU2TbP6Rmc3/DKBZimix1XlQZUBt3TLQBRnTwyMeeEPclL0LJQqRKKZVtmF5t97K
esRXw4SqOuDTKNCP7WB0ZWzhDEoRfojWNtPR4Bxo/ak6lb7sMU2jGcJmDMl1YMuL
nrESoMapkohaU3HRPpTqYFHmnO6Yb2Pg0vj8FOV2mrZ58KPygFptVUQC7TQDAhz0
Gu5GiFz+SyCa4uUf1iGNW/HgGh4o5owrStj2jvyIvGC9pJlPKv7QZjqac7Pcu+J+
QOp8n0dgLoHqM7WP3ho9D78wTda0Z+T7VecF4WCn8yrKGaWjuZMi3qbl4AEdXcD3
`protect END_PROTECTED
