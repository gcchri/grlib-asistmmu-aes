`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZqiXK+j0Ns+q6D/9x7Sjer6JRgHxqeFD1nmQlSrXZsNRt6dXKpcOClrVBoLydhU
7WwT/kXbo8j+D8IvR4oc4jDQjRW0mAonkAQCUwApw+9Xp5ndr8rdV04YccMdDkRo
5wDpDgQTl3o0pKkC8OVmJGEKnuapI2WRKczei8G8XiAUSA3tRU3cyY+7e1RoeuA2
Qvy9OkwbYP3bBEqaZ+wkU/SuNGjDYp5CdrVYwkM7qgQmEyBZAxGNvv8/OOvT7fm3
U2gDOI0RPHye/POsaJWko0ZFCcRvtdxbzNMFr8OhIQj2aEa7waGo/r/uq5z9A+Rh
p4yCj+kiy3kh1167LoSMKW6mElj6p+e2nqRykiDLuY7giZvVrBAIv5NByhI7HU9E
9d9Qt3Nf4nXTE5aNeywmmQG3hLfjOpQeBGnoAz2FRbCg3CO46HSrnodx4ElwtZzp
HrM/ok+bYUgXdQEbH2vNn+2yQ8AUEbviAXrOsYr5AhB16hFtnzZ8PP3l+6J0pgHB
oR4cHgUkEJzj58h9bt/BVgfpBypcq6Yxirc/9jUWMA5c1+nm6z985yWXRehuj3uj
L1jsq4QpkknacawPv/H2dFDQ+zijWJWR4H45Uf/xduToxTN8LYAb+kjd6AzYCTGf
rW1rdSoz8l1aCFasJCIv970pNRIjaMprUJfT22tSm+L19bPLL5wDDbKKWXJqslX8
N5lT4gkO9V1dTcsozhYnw9IEdaTKeZ9iuFE7wutUDSJh3ZjZlwy/m4wuvy8JIhr4
LqKLTQ0kzNUeJcMj/ouxVxrdXpPzFwP2zuyzT3/IFQlJg4qKK3qAAkiRTl9Vs+ud
mrpX0HbFtrdHiWhX97TRVp82ZOMd9VOKD7SvlzVbUhs=
`protect END_PROTECTED
