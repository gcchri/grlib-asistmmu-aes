`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vot+m+0DFPG/uIPC3g2ACEe90J6g58IEyIhKamGgGB9u+aU+RvnKXgMzyPiQq+8s
9bg5J6+ok50iaCwS7TjTXHzEJGHWgoowo0uyOr4jS1p6dqEjWEMBGrBZg/baCm5t
J6CKfWSGUFENxUtGkBwGMHdU4MNTfiHMYAwiZ3ja1xltVKrJ0BDyqpWPih8FdV9G
sKrx+tTTIAiwVtx4XvHEpx7PM5GO/8G3XCMYkJl5pMSIB3DmsDx4iGHury/FZ3SS
G5LxscbpR7R0B+S63p3oww/RYS1esh2YddOG3VtdBQ8dIa6s5qQ+WfZtHa3g198e
fdPTlhkruCovpHBIWYjRV31B9U4ct6O0Y5P+NdvUF2HD0NxAJYsBwpDyR+EaYKUa
R9QnOl5IDgP6Cmqcn+iZcJNhMUGfiLVgJ6Nzb/x90K4UN5dZb/ORzXN4BJz4f9dz
Ir2QLUhyVWcIUgJWJyRXzU7r/WV7o0a+Vfujj7A4ZS7d/DzYNS1QbDmdppRBsHuG
CeUmXNdi+ptDDHogbuk69aRCksB6iEPGogbkdTiNuYokrq3frFiysmV2XyGMa/oj
qd5sBLpHPGbHlaf4zaC4ZCmtYDZeOLf5DTz0nFS20K66pwCAkQnLMTeHTx0/fJ0q
lplWcXuNnFiSFFkAQ4XqT16wUR8IxEukF4FK6ugxZ6MGFa888ZKINs9n0H2pFpBP
rG3rN4FcG0G07l5oI+wFM8NDjOZcy+HIae2siNl5h/MTVgMmcltsj40HdPrQH123
4diVTZl4L+zJpogswSJX8poJ3BpqrkAs5kRNjIB7iQfNR6M400pT7I4i8ToMWs5z
q/Yc+uaXld/V00XIJNSAlrMZg7vtM9n5rZU+8MiXzb0tyJtMVhgXaU2KfJvCsCDM
ycyTrd1iaaR6KZdvhtstReC/6gp3VDbXpBst6cWd8oCnXHstj3QDWzh7wx8f13sk
`protect END_PROTECTED
