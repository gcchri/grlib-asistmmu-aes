`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LS2mp+w7wRVUe9/2M/fPuPXPbdyFWx3BxLtYHzRyhBnbP9OHjbBnGBCDNhbaEFNP
T+59GOg/H4TZa6nykFxQ2M/7ZzXmEb+RNJTwpK6boQmtCILXZfjJVsEEhP/k0bCV
PZITYrAJ5zrKqkbjnCEiwDmgnDlsFCHwCmddYVhbqCXW/J98bSsmHCE8Lw1Lo/P7
cKvY4ljMorqGD8SwFxFzLd2Fm1v15vi/noWAYU6amzCZHnPpZELi93XFaUd9NhwJ
F440Ap5MHnUKZtjSiXwFcbbtPNowskpiTrrBNsP+8LqzBjrxxksHbpVbdbkjg2ov
SUon4jgQSpTtiixgkH0V3d578SlJPcmwhAXD90r2twdOBHH8QJH3VEEf5e7Rk+Ol
gGZEJfvu6Mr1wshxIQ69YC728U4FQuf6hNmsm1Z46wkcSZjF6dRE+5tgEYylNp9v
b3/rYt4J/zru5rdjuuamAwdydc2KuNqalscvvEZadqmbntePWh8yo0wKtSwQddwm
5dQH//ERpYhN9x8TVLEucG68hiHKkb59mp59+MVHOQ+L7t/4KyE6AGtOX1us/BQi
8jym9aE1BOyH6I3IwRDN/13LSFAXl11+z+oPYalltGuPNnG02JLI9drXUPvuPkDx
Qf9yWMLvPOveITSLgNfB1lAcU2y7HTPWf8e0RhnHHfTQLwHxFF8O2jz7dz+EgDpR
CreUK7lxkB6Kyxi5QMpNL21rG3BPU/9tXErZmE2ijF95q67wdKyRJFi9DPT1kSqM
nq6QSeqcco/KjwESBI4bxIXGPYeYc8cfWVZcG8IjMd8R9M+qZWUBHnRwWXNzCrtQ
4xTcO1xHbdLFS5BQhi2lSd9cfktmVyhq01BjWtwOZzvLBg2F48bmNboj2Bf9945O
sXiVD4sBV66tcLxtft/z0zoi5OEpQl17UkhH2c46IS12IiBoDgI3klcVCJqOeNYv
P3mr3w6lhxHV7QigPVAmm+qmMQB0vvXj9QPX9Av6W+4updfM6WKLs1CFQmIaIe73
hhR04mZP9y15nsvpYaACWeRnb4FmEp9UV8R/kidK7qhN9QHKX5J74t6POZr5FW8w
nTvkbN3Iu1H5zdn9dSNTgMQUa9j7dVQrQg7MlrJK80XODSYuOIXzVn0G5ZAIlTuB
fHGMzgw8Fk8NjrrQ+6NOjZHyxhXgm9LLzTKbJ7b5JQv2mmWxuh7lHCvC38tTG45i
t63qIuD6hQZsikgAJPxChiBqXT/kCGuGjOsjVG0XijeLNph2t3yvlDvJiDxgdIhX
FGQdBj6ngqVAuFqHiOjVRt8LYIe+8fh3GSmtjb74tE0v+TT92QZMZj2U65mimHa3
1a4zwvjUNS/c2cAI6Pf1iUOlh7MLa4Fy1nPyS8hhOfiicA8tg6MShDdMCZWTeSKd
UUXn2UeAjMt91CblShUC8OY5o5r0yFIV3L1JvC6ByIppjk7zi08dk9capx8oqL2P
MuwJndUeefU1ESDsYNde3P4MOgHFeo1RihgmXc6JSNWOM1ofx+rMPXUQdSaTWiYz
nzDIKm8CoPvPbV0GuS9tFSlWachnJ0quigEHHvhQVtsPvqJPYpflnUY8PKYfngfZ
Vexk8XJW/P0GUY5aAINRSqXdfvEd0KXTy6THLVlVXE8W+QM865i3Xil2SlV8kaIp
PuMAuKTWJYyZ5EjB6LaNaHsePAh/xM9miw9vZO2c6S4q6I9EeN5lW4SnScfu7mPE
q/58zoNNCS+mVxuknTMmYsDxPxDhXf5kS+S/JZlL9bRfaCGSx9VHy7J2qLaSi8Un
EzbjkAZb3HVMs1oA9/Hz2xNOKdlXy7BbWVdiUsEFZYycMO/XfU0Urhw+Hj+cQDJD
VTbulZ1RoUf0GFdwk0jI4ODrRv6C6W44pDjilPl61IBUYStn1rcDAlypP3xuZbTf
81pIKWQrYUk3PukDPAa1urGVxaPHWGGOoKXr3FqjXgdd9G2ZPYUHImci4YuZVepT
9JA2N6P2A1xZrhMForFezGx8ttM+XDsWbqvDG53T/LgAuVsuCwk3yavC5Yp9p4sT
7gqPz99TTS0ja36daQd3/XSgg0D/yThyfqr447OssdWa7OPdvhGMGZj1tmII21Tq
SW6K8cRHAbvtrWhB8z1cktXScmMianziZ34of5MB9e1qve4FLndshII8VaQc4ZGB
x29obi2tTsrdUzhCWYexGusMXlQ6PcMTCcLnyQCkm4FmykEHfXHChWMXqdu2Kky4
Kz9bPDXpRwqOWZSCvUbFEXq/7TYVhw7F/9zswTGvQkY5o7W32eieDJkCHjTJBSYS
DKnRhYZnM8LsqZoeaIOgS+OD+krOotu9KIW7gYHmVgYfH0W52KIzUb6/aX34I7BE
w5Gkpp2dOArETOdwkCGP+eoLCR+0sDdQ9+jouF0NfdU=
`protect END_PROTECTED
