`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qr7esiFTdb1uofi6/JJ2VNrVPq6FEnauKiiv57U+V1Sxs43sqog67JoabXayYWeB
9sPMu3YO55ByWzAw3XmnKimsb1Tf6+h5RIEGDDG5layJyJmBGi0HoZiIIVjrYO5E
zYOffasJ3VGf301Br7/aEI3m7LS+HoJNXhK4/XpWmpdSTpta2bVu2i78bC0TVIFl
OV1Rq7I6qUt/mWjtsf+JVumSRD0w14N86yiRVMArbhlmQj8mPi1JGoJzhZM1kAGU
BVruWu/cSD2CfzTfBbWHDgHaem5yNKt9BRsBa2GIV98/bJHeO+Ei4rnUZ/A9Blic
0XTOoXvVOEg+I3QFM/h62uj/vYEzzKjWpFFOpBnGE8z0R3yNkB+W/1E+4IaXRDI7
0o6T7B/5xP8t25ZaZesW4BUEI488uO5tKBD4rYoh201FAkc/m27styXJn/Iw6/lg
MzVJV7zBSvhTmKNUjfaQjkAPQ/xj5F3xO75H2Ia75fUKBaXFNA531BNsC7QkrB1F
KTQdadw3tPTtT9m1fiRe7r1nH/rLdUZ+bH5X7UxKJ8ZORJFdU10+IUbE73Gl1YiN
GgnEb2mL86KfZMYoeZBgKtXoNLlrkKJmybzDSh0pd842qHP9DxS9K9P5YXc+UEx+
LcgR5+q2GHxglMVMI3Dy3JNp5WoxNSyWtnvDfO4FG5Z1DGjJBuT3Y1BShWwJvVEc
0ycVawqWMJr2AFYGM26mp1+BkQ7FCjMWkgWO7pHl/qk58Kq9WB5IN/upUxYgCM+Y
F+klWhgC3K+49V1de2nY6w==
`protect END_PROTECTED
