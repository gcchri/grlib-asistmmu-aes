`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0kQOetfOb24QuNlfitCOUyqhlJnWT5ZpS/FsE/f2PF9vu9OgL/H4xvJW9roncFUz
q4MJXzhP6loxermgs7GGubWGLWA8gVOrEEYeDCgpbxKDfDBwPI0tOVqZc985vvpf
Oj1NkAjkGZiY+09EOwg1LT6SgO2+WYMqOeBleS3W/A3P1k5smUL6ZOkPIkOZPAJ7
HsBNlawZwHT0blaXW1N51FFjatpOjnsJQW4aZzC0SzaygvnRShhjIzJqrqO0F39u
A5eUcF5MoQZ1imI+knK9saq4BQVKRfSqjZZG8k3aRKJZcROxTgRy8JaZUfcVntpe
3SZcxObS91CtzcnKoJtIGhBWjmX4eToWy04ojUUZUFfC+2N2asoUFy3021BBnFQz
VBjvcfXs7tZZCZjCX2eDpA==
`protect END_PROTECTED
