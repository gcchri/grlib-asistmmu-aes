`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dec0vymqtNO91vpmC5K6veVpZgC/lEBc1PUmpo/APIrC9udkg16dQDuImdSt0mCU
Spw0zinoPh2ED4/ItASeKp+3+EMT3X6kvBpM1hGaRn+iMAD4h7PKhkK2mPed5+mz
fMLRsS3y7yTkq4guIkpS0wtP8RoFx4SHuZAUnzQAUFe+S12F6MZPhm+5E1hItSm7
90M8IviHHivLe1HsJBF0kFx1hm61K7iDJuL1l5GoCjSM/oNM535dI1MVIxMYPMi+
61U0IDFG2z7D7+7dh71aNw==
`protect END_PROTECTED
