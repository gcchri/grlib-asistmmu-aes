`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s2deDyvuHF1dy2qhO2AlEjzqzEMrZxl7xMY92SbIG3krGTuOnHeLAaYJfFIKxyDE
wmomD3pM3rZ0rATkQwiZnIJ77SZJmye+VEjoVAYnD31zbJ7e28rTB73av25W2Bvw
Zn/jTUWpFQB3QFfAPvaIZEdKQwyJe+BObEbuJ815FgPrsOil889aWT4dpnAROPjR
qEsfai/iAfspfQNEzuOSJlAKACpvv/DStGaDzkcjLouzupgxpuDkcEhP35gnFVj4
qYkhzLICVLlm49Lsy6Px/ZQBFWpAJ4zRZnWbb9jp2QqSdSHOoO9dy9avJmQOUx8U
AXXEpyCCdlH2lDHzDIqmNTl6gNLAhyxTewRhF/WQIyJXKhN7KMryXZTpoX4B4bvY
M8zwZwY+mpLrsux3A3VDY0MQIgzmNLT39S41LdQoGeIY96XnwGwmOfzgtjXiFWm7
SRXwc9x+b3RF9m5jP8BX28gasWQSyq0c4NPUVFquYiWKsWVDLRFhyhNKfgBG5TXO
ytphf3+3y8cklzGTCGCHR6enMUeLdgBJm+NUH6jupG6z5783hA4MR8AR+VV5pMSz
`protect END_PROTECTED
