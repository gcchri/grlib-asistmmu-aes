`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RGmRq+Y5QDVgSI4mpeiYr59TQCNE660e4KFBMrCja0sX/ayFRswGEwlgNZDnH1Pj
4dpTqyjT3SrQ4i3pldSmtleDkrgJdMcU6VQMNo5jgKU81cU5zKK4G1DYgFVS8Z8t
6uXKM5rdZPwq1Wqf9oOrjqHMDs9aJIiiUznuVRDGsp2rQbq3YSKubC3Y531L1IU5
qqNHbSEcV9pI4rlAwANVyCl9oagzANJVpgaQJx1tX/yru8wysH65QiLKUz0rePmh
juZkOkxtHIQjgE5b4kp+OpFL4YAcROt98dSvbPQtmHObd5uN7YUSTLO1dTD8+lWv
jkwnFdAYaNGlbo0hzBmHUwYHK/8HRjcJJzj4rm4Cmei04HZNzvcWH9+Bt6RasL3M
HEdGiV5yemD95rVp4D80BfjFHDueCmbhAIQve4+Jew5Up0RgAM6qScnD0kENq5Cr
SwndFN5gF7O4T0PU2Fk469ZCm08NJfIqF08YswKeujSpiGkf9MVCLoXZCWg4GyA3
2X3q+5WtvjUVrAcyFuumwd4VUakSbZMfhW7nvA8S4OaLpohx3nOP+w/YMpRHlJ65
NjkgyFbhtEAUoWyL0dAx9tlY8NG4zfg2z958nAMt5B+Jwdonut4/5MdS31+3YlZU
14UzLrA4dMzyGaFdyD4yRmAOC7FOE6IUU3clZ4voC0RFDl/9KpRHn78SqVcVdR2i
wZTmBaVQZihOwpf0G6oF4j8CO+2AunxLePCjz19bMWKxBSy7LkaYr6y4UKrhKIGv
H492hSpSRNVBQsCnKhG5H1mcgp+s8iIgxs+9YM/SuWOffwOarZ1OvbgGcSdlu9/f
b3J0MTwvAViRAjTrLRd4weY9M+5qWnCfKATIvjplp0JQ34yvqmMCoZ44eayQ5Zeq
Jg/QksBo9cmYkLj7eu9x+i92N8dTCOySzbqa5ETktdXisVIfPzrmcqs6tQPPOOkX
1J+0mWeP36PcsOfXjvjuemZh14a2qHkBp0zfaWSRYac35E++jFeymlCbNylxLEaU
BYvTXd5u48yahqp4lHFaakKmeT2vrxXoXYeX4ZASiaXGhJeYqRfcQJghgqhb6wRB
b5mkbKmk8H9g7wUxN/NdNA==
`protect END_PROTECTED
