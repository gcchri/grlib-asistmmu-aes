`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6D345nKSFstj8Lz3hTqd5cnBFsS/pzmRP1fVtnzIsoxzjVNuC1AETaDP+LbfgTxY
T+K1q29Z9o0sGgWFmkOUvrKo9exBN2m8txl0aQVKSATQoSkmbUh+VcVUHijGCvBK
/L4jTNmJba2V4pZqPX4+DCCWGtNU6hdL5GFW+Sp3UXKtihcnUqxAn2FS6NqOs7pK
o0zh0RLQ2JCBNydvBNu0tVa61mUCWx5s7roapsn64NtbPnYWtSpewZEcT4s1iHOk
mxHznBpKLJzw/D/ibqxQOW3kbNu0KGrj+wlaof5/mENNw1SdAXeX7X8gm7ZHoAuT
`protect END_PROTECTED
