`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t6jZ88NELTB5kEbud5S5K096usPEHWirCupfbhd/DKmS+BqG+aSx9/nImyHfTsuO
caIS65xeJ4ZLg+aAhWd5ObFG05FWYO7EIGepNW/36Cd1KXPe4rt9hxpyzVlOvgRl
IJsNwbAkSUN+yMMNDJ/D9x+zVITbMkLO5rZI1vC4AWB7mftGBt4t4waNQNHq5XOF
6FBDZS0h5SCGX/Q06eu9/u4EoVJ7m5TpBd8Ujbbv0Vwe1gU7JQ+WcQeJSb9IsJfZ
+E7RZSnYR3pUTwPi3qqsQdFog9rhB0ouqZ9GEe71NETqDsdvuttM/0CFh9b36ZuK
DORaqttGFa0mbqqnybzbqQ==
`protect END_PROTECTED
