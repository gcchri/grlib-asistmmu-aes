`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6KMz6wd6ntZgz8W7cl5YG9lMaL0SbVPLFex0Exg+ZakaElJ3wNkzJzYr1QmrolG
SnWLgFZ3CMK/7Umr0IoJIRE/6dakqy5bvSgfhq8+e1yy0dbtRmPHyIQA+0MBcwRQ
PMIDem2rsrVXliF65g6HJgc3k6uoJ1ggde5N/3VpcmagrEk5tiaSPXbgHldf11QG
G8AKitsoSXRMhYEGbXCpv5d6f7xLE/m7wHBuZEc1o2983nMENiItQ9Q2P/YA1kxS
QJEyzG/PepTCds1uV6VxiqkRXEaHqj/ajmbPVWzHEVIt+hDsquoEHHG3cbksnIiO
Gx54GQgOyzQhWcXM2itEj4Cp7rxfl2SwaBG+7/wR41fOeNTpFZMoLbNm/I/5BI3L
qN8uQtMDvNVafVjVJUZug1yzuxnpKWmRRoFmlnUO2lCKJrV0PAyBhK7Jh99QC3e8
Qk0osp4T1ohA/F/zUZHPSHOt7GQD8H++XM8duXdara2N5t5KSwnN4zmD0/PGEpEP
MU5eeEiDzRCzFdp/BYwvxyBhxW0BohNjEqdvZ4yusnEpyxKzskYeRtICEfJaYIPG
13SPQwNfA7Y0J+tDBJH3RHlsgua8VAuGJHllBv9S0rRZcHMHF5NhfPOArtwsJLSm
m6wZblVljOFCH1ydZC54UKRlyyzlrmbp6C2TXGF8ZPdNa7oE0UFUpx+uU6vYPQiP
Ueba6J87w1uQf0HweXBxw+byR2X1NfGSmBLOOa7c0Z+qW4AI6CXOJT8Rb7Aj5quV
eDo2G8Cl6VB/MGL4NYftyQYi34WdWlSQHz+uhox/KTUYNzyGZsTuGXvETH4nTA+x
EESJEuU5MYH1MXLnpjsQkFJPvYZ0lq3NA+9PpWqvG/hx/MYOpAjW01N+NXrYWKIl
GQzcdfhPQ0WikeWEq7KHZP4F6vTqnytpEUc4scnGgdGJT71PmaF1SaccEuLRm3N/
Q9QWr1pvqY29JuGjnGizQkcFIseVLZQrQutKqCsBZ6qm4ZLratha5tcO7mqtORxS
B8sRMlIl3+xWns+xPnAy+Jz+tuxpReXqjSQFFJWYGlHreC9qC5/incIU+qSPcDJS
8AMvc4SC3KXlQjvq2K4dqPjObSN6xtRyl1OyytyRussq3rbBcD+ecEgRhEhBpC7n
`protect END_PROTECTED
