`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3CrKTzpzfR1sd+cdzZ4fHPcyK6OBC3U73w5hN4z+13PvlYlP4Mzkp3eSdznHQEd4
gBAKzapeypSZKUtwAeWEXPXeJ3S2OQG4SdzXPlthtX4t6MUWsHzB4Re4L+A389rk
UYkSqADItw+7reyXp7XLsolXUAmhfFdjSugweMqdmmlwAXD/+mZ95Lt5bZCT7J0V
xWGSvuZy59CZbxh0sajWgV0CGJK4rMMX6m7Z9kQQhTtGy2NheuH1px/hDQbTrjNK
Y+obZB/IzlkdjPCmBtOsxkiS5qgZ8WFgPuK8ks3AWxBlhcIAdcOO4V6um83/Efnl
ruJ9qVO4m3oUbyHTtjs2xCLIpeXPIcrLXKOVAI/DgnSH6+fTiNJZNqePoOQwHvPm
h791ijcHn+1iiaQeMnD64HJl8fgcGrGzg7A4olSqu0M0VSN5JZ8dtVKSBSBLzVHW
LSSVxoNVaot/JUSAWJGEaXQnVXvmyY9DcTwPBD0lYZPKb7a9mQ9bFvpyjnMsOJ+O
OZES6NNT64QeBt4BNUdKo7LChuaFlAQxIxTyY09GgYuoDdqtSGO910m92I4zjKrU
1eCZKG0i9tUJeez7FgMCl6JudPdIMmup3j+XtbQa64wRQcW6yA9OqmBANwCN3YDZ
TjhQGY9yw1Gve17wwJSZGYRo6Ui4AJF3mBsDh7IGKYp3U5bUQj09msqZR98l0XrU
cXOuk600v8sQFDfj8SjFh7nFIcQ+/u19OaMkif0xbIA=
`protect END_PROTECTED
