`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u1FlcplcG9HSWrKwTLGHU9MdpvcMlZcVwbdwhPVtZ+v+TWU7IbX/jv2lC3gza/Yh
/s5FT/S/dHU7lly+YVVLqsVpPHZNJ36Bik+7yzzQnAWxCryzj36bT715mkjE7XbG
FfFOMh8UzMTBSQORnzjF1jKcxQQd+ACpuJbDDO7TEoYth8VupBAAxltxA5M+ONRz
Yhk9vK6sNPCuQQGrTLGWi6TbWFfGg6lVPX0TK/eapWi/lOzOhEJt05BCEa7UHGV9
zJyZFWFq1gZ5i1pvvfq2KSH0874TveG4cyM3a44DbW7TDGEX9R+4O9S7BD9NcTnp
24yOiPNGuErQzfpiHrU68RjX/NVXoRtIl11BypCcQOI7arpc7J6Gc9RkncoBbzPT
`protect END_PROTECTED
