`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S5X9jYDTrRs4J9P4gscTpNfJGE8r+FTlx+sfKXjg2DH1oQ7u8zTuWpbRAKl8GySU
C/ZBcjQUCNvYVyFJ8smSw6K3RlOED4RifOSHj24yj2iNL4ghQcANShAzKi74DB/r
/SEVZYQZvZzPtAzQIekBIkbxnk7zNVSe21pw8T2sep+1bbwEIpja60+8x12CVUK+
ASmfM9mmiyQwoaY5z4E3vAcmACwRQ7Dv3AaH5VC+8mvSr4LwVB0h2fXINSDMCasi
WlOmc5D5ZkQkd4jawVPUr+jkwOwY5UbsELOU5kBPYNGY5OcwukJi7MSB0x6CyiYZ
`protect END_PROTECTED
