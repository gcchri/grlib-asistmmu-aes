`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ddIlsGP5rUJKc1PGjmbNqnGt9H6qUS6CwAOiG54VKHbsKG9gq50NMXMcqsHBfEND
mqQvk8mjOxeT7kSjLTnlf4kEWagtuzqwwix7RPe9m+Mt/tFMOMYte/0Fc9slxonl
N7JzzqmlLw06zdGeJmrivX99ZU2jTji/jl/VDEj4Fbsv3F/1zSGOkVEW6IG+kgnz
SlwFGEfAK5Jnyd04RTkbShhkkJhh6ySeEPs/nOvll/M5YhF/pYwiUYk3BduT6IeZ
5Td9x8D9UqUbyzAGYf3W+p/VIKYIjXuNEBxAWHrbadRZ8RBjJenCh391uW9T9xKN
iSMMU7AlqpqdLFpdoWVy01GYYUTSP0kGiAlNfRzktUqdq7g8ZODtcexZfNCaoGdq
LHBMGX32J+DBvXRvDGNk33NiwUiC/vbpQT/xz9ZiBeEfXz4Q7VJy6qSuLQc5SwRF
E4jkBahKEWYr9xdsBZwojZupuxQhwT+IiHr1gvx+JoJyiBBPnwHkZyoWyi2biQ4j
bvSi8ywuqQwcIBWnUR3rfBrdrLZe2rT28CdJdGPhwYgyrkEsSKwnnNg0otgLvXkL
jSToo5baLBtEtpMrEChrIT+C/v5VPB4E/bY+amnhl2TbsydKZjQtFPxaTO08FIHw
U43zpbyqNSP1cjOOojwCbnkwMx4pqHm64K4R7/hJ3mvCKKsb34zQZw25i24OyQ1J
jQ+C4Ywd2X5T8mwa9H7NUMXowUUK92H2e9l9k6ZzY2m11UW9N1ITLtiLX+0qEAdQ
q9OvgbvxKpGLaHvx5Rl/WH2Ct9gse7qKNS1s0yIsMnA=
`protect END_PROTECTED
