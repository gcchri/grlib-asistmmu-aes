`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNUJHhqU1Ib6csHkiTFSa1fy3tOUSwAcarylYcwbhFNKFRqloIUwjGoRV8EO35JU
7IpJiZRctXAMo54Zg1JgTCiHNr/wEVVk0939ilA9gdkdJbs3hYtxSpayZFpt1y1f
CWOYHsXDqI1YI/7F5wyedV+oYfOdr2bgG4TrmVXhlyCOegQUCgADxEjg4WBlohYg
IOESbox2pKG5ZCoARxGTu3xoyGUG2Fe7Am4uqwfLyFhX6JaBtCC9utbsuFWPrTXY
hej1ItOVvvYWzURlqZ1Bfkw55XIIQO9C19vDnGuPQkXPFWsLkF40mepBbbJMjjmU
51vf8GVlJkmMIhnFOMJIqjr6rK9d0L+VuR8thhHqweY/1j/M768sxQKa4RLB6n9E
ZfwpMOZy0sn0qM3tBqLsN/M8kZqpcPOspROUvdGGjqz2EZfgLTi10IHgS+TzT0rl
MfSu6atfrTkI03uRqjqwmlWU7B7XgASwBepy5t4QC1GeAvexhWYcS5pCrk0o+gUZ
5bhzoF7EkNG9h0hjnY5uN+q7dFLCmgR4URLC/nTXcCw2BupJ4rfVCuHlP36VM9K4
Xkf3DO/EnPxF7z0aEaHrj1lggJYetPcx8i3VzHRQOym2fu+DV9ivMtYsWKEzKMBK
jOcPGc/ygSPMMTHY3C/MWZoNammiqmeyncy5h9rh1DQ=
`protect END_PROTECTED
