`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCHm9uX1W1wyROwswk2T2H26cYrnyM2MMh5DNWwZh2INO7S5nB9RuilxZ69xZIcL
G9bIYwOHx2+Wy2xq3yJr7XagyUJpyTZpTX26Ap4DlDI0g7fZzlQ/xCDv+frQTwRm
0WjoQVvv0u/LRW1OqVQ6Ir7ykfLkpu+3+Ya+3kdwkqknWgWwkU0ZVnTSd6m1AygZ
Xim8Sg8JrRqDRhQt7nNnz1XDICPwolJHsV7DV+uKM9rfB1ROzwBzCbObbL8L0Cxd
ZHcHE6NH4SWB6lgcLBPrzoUIYRKABLKxXZENcj/UsApa3q78FgLXE6peetD9S2sU
CNP15txeH4pUoU4nRS2t0tmEogGISYXKD0/35O3jFujdtg9ox6ppWqGfBanNo9bu
oyyzcLru2AsZ5IHDEFwwOajy7lE4/KBiDeNhDByqt1k6WL/6/WkI8nM2ZQVJAo9a
rrh+IsOhio7B6ygMy3kowCC6Oz0VU1ATzr5b4yxUlP9mvdreDAQLC/5FOStPk7b0
74/7VnE1IIrmxGJzYKg/tKPk2HThWArDPyvZWGKIzH/H33qkj1+5grlo57gFdAzg
SH4JMrtLkb5Bqt+2gBdKOp0kNU2I3ECvQDoBRx6Q+XIkdtKRSs8GeXsX3XAmBUDd
ps+HwMC2gwRtHqSUdz/kp96UEHxVnIYZrbrzc28Q4u4gfT+tT8SR/uDX33+AzXXQ
crwRnnQE9rflsnc+oHYSlGElovwwMpc/K+c48W0dhu9QBdij3lgV8OAUPdJFMEf6
IEBes6C4cMZp7dmDKBXI0JfHpD8ih+qwtz4y706gAAKcI79Ugs5Hs5nGZpjMld9s
LLP5K/NIvij/3yGFC4VyKZ8xB68iWH2sT6f8u73BZN/TkmwK0SQJH6TaaG2/WQXO
q6loNcR15YmXFX7UsW9oTVqt7k4MHTIU+tgi1LFch+zK3UwMSx0dxG4kDgRJSPaN
`protect END_PROTECTED
