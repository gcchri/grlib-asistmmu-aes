`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/t6qSQR43QZ1PDfqGQiXDHm/LSK6wAf/Mto5vLyh5Yn3cYucI+oFfm4bhwkM9E1M
FsDD4+/IkDv6z0rd/MgZZ8rkHy18NawlycSn7QlxNOXtoAO/4XcCflc6upKs8BPX
ILYVmjV+ia7UIwHNs+6Tf4MxnCP9JQszmxiu0lDdC8Os+zJ7LRsW/9Qnrl9oNZO5
uMunbXrRvQWecePOJLbkcvhnfw9JfDnCSCh+GI7jIucCa7HEIFh347ILS9apEhuk
OzDyjbF3gZEeVLNJBT0Kq2ZKf+NptRB9MDhddfdGWyQ24gQV0Dx2VMFO+G3lPudV
8TBiino9fBiFgtSF1Zn2eCUC9bc0ytG8h+hysXlKfjWLTyao1+2ADzEdX2uASE3o
Co8U1LDuLHnETxlrAyZ8PQ==
`protect END_PROTECTED
