`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRdn/uZeLuMaJI/t6aXcfLAtfnHRLifA7MeYFX4iSZe1cFW/3GpUCbSiEFbKqlxw
hFy/Wa0w+sWIvSLRWHdma+wZwlz2FV8ACftyGwm4LQseADl4rvGr2OWBY0+2ia0d
WnbkAQx9gC2HsP77CyGzZtsbJ6UQP/vRcenHaEtsDmdVGJKD8rFtibFUzlRpcy3c
Yq/iKgLcMc8j5nAYk0+5dZnZ1Tja8hA3enccBa3FfKxH9wv+NEGPzmflXaawORM0
oGrXFGJ/MCMjSTONvTfiG+EP8VCnEkVQCKDVzx3jhAeV+aK5kM8Tj7HkxmuRxijv
WSHNVz54cLKk9KxbcbzXG5aeRMDMkt6V5pMZAYRiS4AHgQS7EyypGacoG1jAa/Hv
ryzNMHHUs+nG7XfbYQ5oBiUm3VHI86DzyMihFAULjk2KuPHDsD6rRwLBscpMBxdG
Pl1sMfZyPie9GaRPfU7EVk/VB1C3owx3PD54f+mK8hVEffY7qCH1Yt3Gi5G2RFo9
`protect END_PROTECTED
