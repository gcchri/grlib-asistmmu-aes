`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aXfxSHTN4amlvuYy+wdWc8qer5BG8Agqe+tpy5FD4OJ4QcRJMSX5yo6rUKh4O9KK
bBrgyTH2WQU+dlwvl/oI93E0Dv+2XCISYXQzOipzzVooYNeZQ+kdZBzRkOoVJ5Pw
OYbuxirh8El5yXRuoDCFxy5LWhzNWOGg0/skfN4MXvdw+QhR88aGcE+lP5YzfCyw
HwvhmSThrV+ZIxvntVhYVUCkdmEdg3+FWSx6hPyRAsnvV10AC47/oG9BfMbNh/g2
cDrk4NUXAy7XQYSzMlOyMq0eGUMqAOuwhBCYvWCMnRWXpJ3+lNbie+zkmvdHDDpj
TomM8b3Gld1EQ6aif80iAmvJIRQQoqPwAxc2ucCKlf0ydVHvW3YZT3zuRte0Aagh
gMXBk0lipDbgwH85xozvAj7wGhRHLewPPHEe65E16bxUmEPNl+YGPF2opcc2WtOK
`protect END_PROTECTED
