`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8qE0GKGQZJJnA/+psuyuyEI0KOg4LTzvax+Lzp1RNXdE0wZwirlactZkytmAus4
8Y7pL3uVMY/kyeTknQ64S+erY/Tttz0ldbc0LK1navaGY/t6pjOnXUuaqPPhhgZJ
xxGj67tzLeGFjKZ4wvwVBCBWbIOXtKiWzBjaAXEplTrMXKNrxj4ijX2ZGOlGULBM
PyRRRWW+hLValrGGtV5Rc+nSltK6QW6m1QpAwfernrfVTuq5Bhl9IWScRq3TzS9w
gwLyvn7NS9gUb4/nsr6FfCZt56jY1Jkdofpi324zEKsBtqif7V12NOMiV0kaFt2k
hkTvHJjHMMWEXLlkgdm46S27NmOWevGbw5TSY+96zvLOznNNFP0NeP71TmGPlxaf
B5Ay/hv0kH4Csw9Pd4tbilp9YLxjM8LwRnU9CEBs0OvFuP5+okAEMY+n2+6UhFvc
vbJEIpE28LxbnBOHMAP5zdxFgqhVSUFI+Kpe0fCftW9KANCqkyFkc0DjKiLTb4SO
AhSXdtxvmaF+zKVw5qOI9//QTDte0r9NmNAJ3GTe1nRNXBjx0GNIlSTMpajxM0r5
hnPsnfzVUpeF6eCBGIAPxQbPZJIAooyEU0AFGf89TCdAsUgTqWoJubVhiGMTLRpE
hR6ZlQJibPyLi5mirhjubWhh+iWzqQDophaSdrkc3P968MnLMZHvmf+XMEAOMYIm
wnXqmqL+7erYCyQ6UolSk5ZKpoO0p0OAI81iZAszvB7TtsrA3KCN2JjLpI/6HS8J
vcS6UsOr5h9D3aqxRyKHQGs6T7DhrLrQg/f5bwJl1/6NzU76yo+53BQYXDUryp1R
6Qbl1pdPaExy3g/ro9Xm8KeczwN/a5F3fs1Jl/BWmP9A18YqA+scMyAPA8mtpnKq
vv4kILiFBLfqflq8JWApHMo9qr0ld6wk+BQfZYbbuz7LVDIn6b7ewvuoKbfj5kiY
gYmsJ0vyHlpC88iVozn6vpybBndW86yNHmpFjsUuDAGMguLejnrb6EMxEWynuOTa
M18o9Pxnnhapu/+C9cl4OBNFQQUshtL4nDkiOrvnJjOh/Th+Qyfz6V2JRTxPtred
PYsiLGH3UkHWnocDInUZoo8D3S2lFkju81LvY+VficE0kRtr+vw7+N62mXapKFxG
uVc/pSRivaiwuQ05Q09JfvCAqnpUu3ANI0f9w+3B0xQeQlsW/sXIO+eNSgbRPJJh
BBnt5Ax83FlSMX0e3YYT8C9Cpx+ZIw9AEhYYTsVcudG3ES7BCi2xLE/fwrMZm1Vm
brTdFKeIIJzrsY+ZHlHZtiRxsOnVqABRoF8HVtsm5lA=
`protect END_PROTECTED
