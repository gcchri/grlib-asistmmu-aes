`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xWvxbMZzm5DDQVZKK5+aHTGA/Q4a+HIpoQUm+LVOmOIFDk07rwuB3libvfPOnwzl
xXthE4BFSLnve8O26FXxWhmx8qhzB9M8VDgEl7L5agt1qcvbWCvBFm45IH0sG8gZ
eWjOdcb+FcxPQwMm1eh47tdEb530Z+QEkU636I0P6p/mzfJ/plL0DvVkaEGKgYBw
4eJ2+6eFKlIhtgme3o2jTPWpwmtoqYRWm71Z2/RYf5zYT8ksxaFkD3VfZTGu5nVT
5gjfLpg9S+FSmBjg4VPkno8hpT8s/LYbTzSWSOxK2Vim1jXCUCSymL28caeORQDE
iNM6y/bAD5aMNT5OvtlM/HVg9o+QpvbCbM4RFlocJnjo9oDkb5H2Ej5XV4cvztIW
Z8+/FaQhLH93v0yemb/dQPyNbk5WxMN5h+LavoQQzlwmI+abpqESlGPEZu+Q1Tr/
LjYgC2N2vbfGitsWhoCro19+qMZKWP7wFPFgS0p6PWEhKKBw2Wt/oWnN1gXSyAvL
VxedcasKVXBr1MJZnrFxoSmISAXRxb940pT9IjGJXaFD+aVgz/+TskB/u4gsyv/+
rmywPj2NvHHDcM14mweMWrQ2a0WRWGNfx1j5IbJCafxHTg0nwhlAeP8Wyg3wZ3/C
p4vcuAg6WHa7PUSQ013dXb+A03uIYl7eR8ywjhTXSsQ3+rNc2EX+fh6A2sgipVph
07Wngp2+KpqcIHISIA8AnZnBn1spEbN4IPu9vKR9Mpkg+gHC1LWRkIAUJqeqsl9c
rKRsWua9+3jiPWrFWU+KycBUwxzUvWl9xwoZAAlyVbx5rg1T5ZdMft6YnbLJ+oMs
u98WA39boYqSW6DTeurBRTlEcXuc23c2/nmvotGO3tzBHQOYt/dAUMIwxPvHO9Ee
`protect END_PROTECTED
