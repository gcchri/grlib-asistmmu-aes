`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Flku6LqP6MjuNZnn/oMCZGOgYtGV3XZd6xOpJhZHYmeqi2ZqKdUo8KvOVlNnK3vX
f4cUcIg8UYYweFMqy/AsZTjuEEp6uLjBNgOQlzhOnHRlu7Pbq8x/WoyZ3SI3UHUe
A7K9m4P2OJJvhAo/WlOsWOqoSWcdocxcPg12MQAEWVrbWJ0x0KpbYDgrxwNkubGw
Ww2CMx8RVEVZTefI5k/DAB2fzWLXIKu/axtL9ZFCk0au291+y3nf8pBm1ZcuaPFM
0tweeGaBgg6LtCIuOT2oOlOrNeQ6p7CdACB0fwbxTyWAIYOJPhq+qmR3Z4P8ea6t
Ov6hzZHunK/BrMl5s886iSJ9bcm/4KOPaJlqcxBJ0mXRRt2kH2DnBFxMzfIN2yB5
PmDG/qSCe8tN5l9pn/umr18Nbqs9a3AkCVackZLzvFxG2HzZepZs0l1oVXIRzaL3
SO2Car9SSo2MSocZSlE7vocKFP2IlQuvWwcTL2rLQRHwykD6lf7JmJ0nhcImDmZT
`protect END_PROTECTED
