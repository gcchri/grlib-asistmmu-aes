`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+kSXj/tNYlFbS2RJOSHmHjcvg5mwUdLgDEKsfUSOnvkCz2Fw3YwbyAKmXGg0eqBy
nawl6+jwG95XBR3kRUvEGCH1nN9PqiRgqlHiVrxBcxBzlT+d4XzOSbBxMHQcCGPe
eJOx14hehxmIVURzP2SCTnfPMeXw3jGuX5F3WzQJPmhT+Oy33znSZ9/USP9U7OB/
vDkwTRtdcXvDd9Bv0qFOWaLNhSTBX3CW/Rdxw0tiHTof2PZCB9Ca+39JW2mWi7Yz
dHXnXqTCJwSA8UY5oMBqdkSnTsFWpSjK3wtngaSWbzRDJGgXkERGpU6B6eWVK4qQ
HwLe+rghUyIpcHrbVn2Lyf1xrORL4mBa55L0ghqr85rekgrQVhni1hYHl1ym500d
U6LYe++koLfgp3m1VVMncA==
`protect END_PROTECTED
