`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AODb8tWc4Et1ue0o4H6miaxN3UjOdYncoomU4mT5Xr1p3YcnQ0CVCsQ63gYwMQxy
borlcV+HUe/2+VhhvGnOEEp5F42sLBOb8WYa0arCkbbgBAQxy7DDfl3PO7dybni0
3gyaoMiSbb5QULQ02u4QDpeQTZIowgUmk6md2cEVSgUl4FuwqRweRoPzk1EFcQfF
E8CWN2YdZYNxgfaewPvoF0KzanHDjfE5rlHO3B+cnKLaZrMAFgF9GZdNIX6Y2ir0
KVTK/vjY6sMQFjJiYaIj0okEunBoozRrGmWr6Pkz8kGZYWs+ZSiC2+oRpVrm0bpY
s+d9d6f2NCMFU0aYAj2iwwDEuCBL8b22gfSpjeYSo5oAXqTvXd/MqB9xJI+A6Y+v
Pd/TgHXUfSVIxq77n17o1/+lWyCHdX8sQXF8BIdlIjHxEhqaQA3KaoxzDE8bYGgx
bEYdio4ZnVzoJXMVF1RfNFYw1MSp01uxrkSsCoKCdvhy4rmH6lZvMVapzOhZeYEM
h3Jh8PtyDuidjANHvIFTgq5bZcKtGW2b2NkrkDz1+r1qPcuLLccWKlARKgfgY6e5
zTmMgtbzkM6xcgaI/6a7eR9JIXsAiRvl5ShmB7n+QO3EWkJiGaDm9pW3z5OeCXSu
FSM5MmTojXpO3UDT/zTi9xpGr116k6txVlEXCya9DK2Spjgu6IcCNJfI6wTuOwC5
iQv5SFZJeOvF+ghD/4EEVMNGxG2lkW2CgKC39wutbOAWguAWgeSDvku0dpreSZJ0
X0idxkR+qIAlvLyrrVjoWBSnDHWRN5ZewFLSC0lId3Dvk+eyvGJ0M2PV1umCdfDN
eRUCVXEEpq46JtU3NmKrpuxQo/x7B+ffbQSqWbntMWF2rDhGZV17hjKAD3Q5IamG
DxS6HHCTZQp8dTMKDlBlovihdOBjCalfyc33XPX9lc55uwKLZn5FKaFf/uNj4FaY
2Q4jYmN/NtZSYFeAAOekchci53ea0MmZFJNqS4GfElEsuDVW2vEFJbBQPEUni+jE
8aGS/sTNwweWjfu97y/iSbr1NUq6vFCB00EQ9A6zzLda8ugCDNdnQzh6hheA1Df0
NMm3/FkK2/hnm8wbzABbMRGjqo/lqsSzbpsGHECWj5hSTWN13+ZMTMXeiXFJhTaX
XIqdr9BZ+Q4mNgxRUeCzjmXATyRHNDocze74naajKPPVoTmx2eclf/tu/IfTsv5f
nQ1S8xzfgFEmStOF+8IAUsFrnAil8yD3iMVfr4EWx5OMd49fh/vsRaTJQcmJli1A
AzLpiEesq200Zu7Kttjw5+g/9icjLb5WT0cfCCVN8KFnLjhbpaiyiee5YuZtqxr8
D24y2c4MlTwpFL4UiGamEAP8UlN1YVeaqjwDEupsQbVHNJPNiQtYYA+/IACkE/NU
dAkNo972TtwfJF6yaP429tBnG3xu3mqR20Lk/GqiSs2F16nECeaUpbMtM30N2/57
nGJsQxKl9PBLxjH+iY8THt+dj7jcndwypKVWCfYBnZyTD9SMZchVu85bE9tsAIrZ
PqG9sPudLlINhMvCc6b6vfl6xzGvfXeENY/aM3nq0mj+ZE9bqadxArYg7XQOHsL4
iWl7G2AixAx5yjpTE3MBu7uvVIfW3wsSzFRnVwRzcGO0kbwYGOkhrazQHWNHtvOm
5yKNhV8ERR1cQslDGkRrwwM7o0LKJG+ABon0qfdCE9vlYHk2n6GbDf90mOMwE8Za
xJQwxLLTpE1pMIbNc9Nm+SXk/zhkZqdeeZ882oJ4mBBmhV2gFcyX9G9CHv4XT06Y
e045NYqQbrQxIRXjXkiHlAYR7ZjZ59R3VrHGgcBIi9dlOmONSVmNNvhapHsdJkQT
s+v45VNA2Uyy6OqSEWdpZehMSnBJPol1w+9LymrsxWmwYHJw2YQrQgT1v7BsqpCs
jkuScgiLtOEkxkjrybxeKapIMN/TUJGTGCDPkZWSJJ8JJGc7Vxkz6AmkiA5lGXAv
t91Xt7SsxUS2ls23UwN2LGyK0+xNMaUJE1MtcOeCpkg3wCCljIBQ3eGObH6wW8/n
92qkeMEzs9l1x5Q9r3mF5RBHNlWBR6KBCS0mrRHYoMginhI1Wu1imcZf2PMoOMah
z2U4MZl+liL+JKE4GzyDdTZVWH2i45wkfbsW48cKKgGVl8tcjQzaByGjhUwxFMx+
+o0kt6yaRzDVScExnTRzenmQurfodt8MH5vIryEroskEdFXlAyC7aH7X2s8VBG4S
Rj/EHgKOufftPGLdtIE5sq6/X0D43jOf6CzVNbwwvGy6LNI/Wul/T0X9lJeTogCl
kK+N6p+xOwmpa2i3t02wBoflL5DAb0EICX09tTkx55EofRq6CVm3axj1QK7XvHay
B95elgxThdSciy5tYH8TzOAPXKn5kZvPlB2dPZeNo+75TkTZsD5cTQ947vYUBxz5
6b4h8XhvkZFCqbq1WO1YdhgWU6UAEyENaDzPjwfE5nK2TEk6Or4NdOQvepVEtMe2
U1GdQ6vswU0aPte3l0HL3O0ZxaRxdeGMLWYSOiMoo2Bx0mJkyCOe0CGfsOmDCyoR
6Byq8Wo9izP8oIA8xH0YXIouKBmtk4djSzxiHYxRTpnmhj8oeS2hTzrZN9is3KPS
ZTyefNmsFeJ1BbJ9hIaNnUAzZ1kP0k8jz0vR5viTMZzkMb6LDPtPZegEz0auv4zm
hncrSuo3JnAXvfKdKHzU04PttTBXBBjO4f6zascamJ/gAtC3OrezHp9kczxwUEP0
uep3BoOWeS5iBwOdMtzRVqhJEQrRUMisuiZdr5iXqDjZZbftMfUrZmwey1QmgQL4
6+0vH5CIxfSXgIfHfuhC129ZhcJkrmxw7wdkNlRe9x3hIDN+8mwf3crhWJKTo+V3
ryh5Zuyo3qV0LyaKlZM+kM0n6TFjM4sTGwVj2ArQLrLBY/yAwLTScYj8L+lTpAS2
lW5BeUNaSzfvqWvWRD+FLLxyTPqB634PxYV1xNuk2pCxEW6XlD1yVgIFaAjXK4AW
6/VrrEuwjLbrMB0hWGQUMyeMdHXob62E+IbSE3yl2GlVpzIw/+Kv7zBYZCS0/y5A
O/NTDvsL8OSTpJKnMmeXf0bIGuF3lHnh9OX3DKH81ptw2rGp1vjUSWu8mllS5FwQ
da7XS3kzq33dwvaDmNYf/ieyMDwN4xmh7U+Xpg8Xg54mzszCpSspjz/D1jYOSI6X
OsVnPjTwC2jFl52aai0Zso8akwnpQZSr8392oRdS0TK4Y5ZWk4qJ4xkQqlP7YJZ7
Jrzg8HmdNU4awUlUWA6fFm4rB5vwSlT2ha9LZj/qDODUKCyiNTc0RQpeoaKPvHmK
BvIygTdvuszrM8Qqv++UujRv6dY7VaPIz8bAgUvASRq5BiAyyzjpvwnyF9r0kd6t
0ewYIQArg3w1MidN3rrmWB3x8Uc1J06h+fjc8yxe84Zkc1aqDSeTAeRMYwuIrIX/
eZHgeh24zz9N7jjtqBcrG6hUZGmzUYLhs+aJo8GuSqMmZlev/70DytdIcpa6xNcA
+UZ/g85IWwystPdWy2TaFW2iGzuBrq7D2P9dXRzNPCbxF3RalmY59v8XBbUe/7X1
TFPsKuGMii08VCn/BYJ1rKweqi0PPSFfoZ9yhtrUTD/ac6ojoJifOw2Iam048U2U
LxHpw8j9pnxxo0Yz+ECE4z8cJWe0T4NNUYoWxh90VX9jbVZgakAexEi/EY9+w5NO
l307fzyfJLoDdt/jKnpKUv9IfmKFgUH0vG32VH4njhEs2BjQFNNeUEU3713IXlSi
UsaTDO9w7+pwXy2Nt99RvI7VqxfIHgHUecITR6gRvOeuri2OdBhMc1dHIp+lX5RT
prfvU+wRmr9NpaBDU6Rg/w6FCC+SuRxbQLiGyvJzO+9vgxo3jFIUD29jJdOrtRXn
Gltpl3ns6Ib9BewD/+jXU4UjpKfyxbcwxIo9kEFYArxpm7OAYk8CT2VIaI785gEf
BQ6caWMuM3O6RytPgIqSCMIO2fc54S34NDU3EggevexZG0CDeSHSoNu0rxOwnQEU
0W86ZC6gkIt6vgRMPF8Xu/hgblqBEdjfm4/jlIrsF/HKOfuqQTCTbFKb0QV7SxzV
vOk4myhIoZrap1kBbopXg02xlY41sn0zjh9/t+/b4fbs/vSh7qVwfHYnoeNcSEX4
vHJJYksFHTWBWxun9p/QfwRzqMwMohYgsqjEmgKWb9F9VOAigchKjvxjVF1XS6mD
lNgP9cAdykdG4JTUEYVmvva3bBW9Tsdc39WHCGnHs244zxnUVgX35vE9aizyspsH
/HWVzHfBYQE10IGsYcbVblqCVhp8AmLaqaJmvbxB+uWsHUDlBWuZ9OUyqNsndQ0Q
mu8QOGA58hN25QZW4hk925wVcBguJR3ZR2ikOmMhmKM3am7uuA/uz+a4Br0QvtoY
AvM3GCzgWPB5wGXlEemSMhgScA8X0Eu2iB2tkkBrn0hHPzf92gVus4O/u+okcC5l
UlTvVGMFplHs0X7C5at3ZNdetTo+iB8nux8hNmQmBeiqrlk84+4YAV4icmY3yFQp
Dn8TeMS/mJJXIfm4CNfit9ph/4wHvcs4DTMvUABPV/zqFb3GwZYAJvbCgzFyh3wb
aJdSgsKsCDDVFUdUS5Td29K71hIywTt5cKQJgtkYcI8GboL+CxmLhxTfzfI6Ge6G
Ljtne9fyDBr25U/NK3muy4niiB0Cel13pwduBZPSiZqLsl/k6udpY2Ow9MDGVTZx
LZ9TiLgCT5nSnqedOnHmTqKDnjRj1MNeGyjSWi9JVYP6e0Mty5GFYRW8Ynw47kgN
urcSF9KpfAys0M6kUn/3t7Hst72J6OfArguastJD7uUMEOTSKg0BvxIMa3c0HzKj
rVIGvsY60qWiSJl/oQoOJuKDChinm20oim05YGFi78rxDVc3gceTLSEpYp6qzbCY
NUvkXwv+2LXk0Xl1TV2KDKhM2TEfzn5lNbOpDmsWl561iAKL4PWelc/yTEhoGxDV
Tuzh091VLZNTQjAT6OOj1F6cbNEEj/qZxVuUD7mYcT5WDudf29kwwxWxu44rQfaY
0Xl+bPz5ILnkfF/erE7nzFfCnf//tl/WOHD+kJgHdN/jyNyu3oXxeiVjzo2sX1xd
3gdkZNMeMuukMj4BiqdaoFydrgRZM7pTQfOgp7xg1ykfaZIvQ6gS0kTg6UbB2BKv
FHMDMEidKlve5bXZMjJQ/4JtPuO6GuOWD9Q3Zxz1xKJfMqtvPfOjM/GLMNwE1QW7
JocgyOHOpsvNa5b5pyaNOI1nr+Fwkr6dHjl54DTJFTR+xZvbTpWkO9tLP50i6ssR
eZSfgcja0ncGpaGOy19fDMM7IIrUON2E9MB6lJg1JuMhJTA+zKBa7ZuPa5pa+BwG
MKTXSL0oxWprbHJAEzb7MJC70KeF8t/5ZCeXOvBJNO7Zyboab4lt3p7JpES/wCHk
QvRld/Z7NzhdYaX++w7E2g==
`protect END_PROTECTED
