`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBjZ4tMp5bCdFuJfWcM10hlqTjW2YY5df3uapGkJpTtJ4vs3QrsOwxvB1IQUeKay
Lygy3Qu5VV+NMFiJzXuMAfM+Ge3gNHeIyAOhLMjHcdmrzS2Zo451+4s7eV7JrCmV
mOMy+N0RMPLG5DHqZuGoadHTxlNjHOLTYcB1MHHbMqxCaltozRMqoeC7i7wQu6oj
FTIg8PElXhFLMmWJi/cjcBngg6KmCOLShlvIezhm9i/BbBYgcayV+v1yNMlFkjhy
EiDoTIdkEC/4SO9Q/uEwiEtljAdgGMIgdgDr5MmZO/MHrl10evUi/tw42c2Yweg/
0JC5tDR8VOB+I8HIRow4fNSQIb6+cWa6f891JFXPdB3Atdl+6FT33UnZZNhBhCHa
gNDCJaSe1+zHie7/ZmB1jlkgUcdsgLz1uQJjb/GXN1uKDdZJQI+WJMAmtsChyAYa
j29RJQh6+6ytw1g2j64t0chkH6lawz2qgAfs6VWFxkla8UZ5qsJaQY2tQinBsko4
Rc79JX1a+j3izqci7vTY5Tmb9GzQRhRQ124X1tIFHUJHUXodxVAx0VcKjucKDzZt
RzDL0obvLh9vgjgryB9w6CAxVXOyBKoLJOcaXS4g08LQsJG9aPMjhbB+Wci6AFpm
nVWpkYU1YGR2+3QbHrqwGw==
`protect END_PROTECTED
