`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cmxm7fEvbtIo+ygl9BaWvIayP/cf5i1Lhqz+nyMGTRFNSH7jBdQEHgh9SLT65L7g
vRswdkh9Vn0j3H1wKe+Jreom6Cnp8GxP6KhprX65v4xJ0J83EPlN9+IWa7kaDLMo
Mv6cKNMnFGlauFfj5Ypsj2QQDZ0U/XWFx+u6ms7Y1q7GlySq2eoVKx2pwyufT0oi
lEoePtxufKXcmPs/hueGh+Q7N3U1ui45uLarO3yIkVSCq1Q7L3JWH12hzasDpukh
4+lP209n+hoW687ARIQhG1Js40n3XHScLyD/PCSojkegq9kWfQGvialnCFiny82V
6TJT1XEn+NBy0QM+K77kvwQ1BVS8zzAHuFgATrDVT0w2Ily9PvOQbVh5edD5yfL1
m6wYyezaiqthBhwkTUDwIPA6HVNwU6vE60KJWm8IZFLcSSz95mg3T97x6Agnq8je
6U8Qo7Z21eXos9GjnUGVextuGEtEjJYVk7j2AKfXIobVB01wPOAhXsw7INHmP40N
5KMCdtj7Zy8DJLAeFDKBE6NW3l2skg23WWxWASjtGrQLok64GbvKEksrPDA5sfF9
W1/hezmD6PmM8fMaGUbfhgJzCpk7HNxPbloe9M8QSzj+Pp3HnZodII21892HAkge
zu/4a87bnNLm23TRSO9cAtDwbjBJk4BpgTz1DTcp2A/geBmu4R3s5D7GcFWStBK1
GESY+d2w9E+i6AfuGFX5SNxmmmVsF5MJaXyb+wBIMp5sRqdDIfK1gP74/pdfxot4
Kvawa53JyRzUAkllX5aMgfg2wA//9ARpN96dDjIER3AQRWS5NWoxJ6bFchMjF/hu
YmbsWGRAh38dN/6x767HghKEWEP5qamM8MlzkgMpU79lU0hLXfHdzYgC2NISDxcD
HrLEhJgP8v4+ZrRfFLj58WFnJPM/Tp7lBAw5H5jNWpJwJqTvF+YcNV/vWsMPmzDS
`protect END_PROTECTED
