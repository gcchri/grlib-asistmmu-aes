`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FjEbPCNSFSVuGDyeeyV1WF6jtM/zDgeJSttgVEjqPFdieaLtIEushskhk6b967C9
+mgXcdfiFmu3lyTCG8CMsJfUiJD7KaYPJn7n2W/4fwwIMpG9YqL295q4jNXi7EUu
XmEQhoPrdEMGt1ll9tHt39GyPTDRQ2wCvwGPDGkF9GFOuWtZYVzNncdjgMxRzYo0
F/41O6ZdbxvhobePnu63AWOwgffdpKbJF9IJPWv71LtZ7uhWrjZkFeAqybWK6FEs
Fy2j4nv9vtljdCsi/5vOazoebPG//rI8u5rurHZeo9OKYrpPWRHfxdeef2I+cdk9
RJTfE5RV/njCanuFCWxZgEfd0QbeC0H1U6xQw3n5AaYFxvTjeJudQwD7rsNIkAjY
jQi3Bllaur1tGvpDup4UhkFx7f4MEPq0wmoRogxYh0OQYvVYQZ1wWoSCZER6gXX4
qMkAMwyhffbi2AZSmfR427eCK9umZJ9pBqGAQlTFKLU/XBHE2jwuuXcsfNzo+g54
d5cXjHytf+GMJf9eQepjAyKLw8qc0jduiyf5Cb/oMTjVte9QGDtSKC2s9xAVhSFj
fOfaw8tkM9jtR7f21Yvx9GP/Q+RvsCXs9ay7Ek1Xn0+TgxeQdXuK+m/s5ptAwopv
wqG0AB0f4udK2vMCT0Xn6GCoo7aCQ2OrmGSS/kHVsKMBvJXiNq9+fzlMLBHf0IHP
UyoE39kfWZ4KjH6CboR+Sl7CAG4Sa4QhH+TCio9gYXuBc6C0oJVBXWRPEy3QcHnt
ewPwTFn+ZrqJmqbbMBMLf4Xrrhl/M/RKb4F8Uf0aL5B3NcERd4c0An3vgjZxbTD0
8idn23rHdduzwULT2orPRkyvJmEogdaU5UwJr6c7/0d/NyT15tO2VylQbpBvrnMt
Ltee3/dal7aMgwKJt1UtaZqKQyJb/kNne/AlxbxoE/2JwU83G/ZbZqFlzC+pl+IX
L/mjBauj73jUYzgMuf8EMPX2+GssbVsI+js7su4W3qDr9S0SZphCcWVTo4ticgLw
vxYGbg2SMPjVFKZGR9RbySrSvUI/yRyz68RacMCFNW6mG9vcm9qo5+1j2NBDpd0G
raHLEwWPfZ8kEjQlnOOEW5cJGgCjzBi6Bh73qIaV4bVwS6QLrX+84ygiVAyWwnCj
sXnARr/FJpYVLpfrA8EPpsjq2dw6Tx5zAACJQdkzIleslTT5N0FPpPKsq7/ZCna8
XT94sSyRILA6ZeshFevnaHjLJZSr4XSXbzZUWx5DeWjFGRrZkcdlDb3yf4GK65jI
YqMaytJYslxvQQpACjXsgCU+5+tvHPB1Rgn2Linjc54SBYe7V7JDmxR6shEgagXf
/ikzk6eaxZWKbEHY9VZLoKL9CtM/B2/Bo0ZXQ0u1AbOIIlMfTE2DnCVuZ34Tg1cU
OVwrNf+FcUJiRwvaKTcmzdvTp9mup/AcxTWEQt7OCRoipec9HPzt/AV9PvlNQWxV
`protect END_PROTECTED
