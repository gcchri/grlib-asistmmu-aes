`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bY1yzgXpCc+QBD9Ckh7yDUGN60AmgHRxJ3eIoUdA2BH1fGPTYWgLy5q3ZkZpjRrl
XnDvYMT7ej/Altx1S4UF8aSuLwiuNza6qNKvSu8MRllokD36VvTPCnp+JGufk6LK
+jRYJjUXni3nk3YG45C97oCtiJ/sLghjHbNhvgpwNajtzuBPmeMx7zHR/y5xyZZm
MD+6OvfioPCi4B+txQENStcLgGQ9cpeUhuSEvebFo23404TBgKZICr1Pz6dpvtPR
I4Uo6vRYeFBRArIHJPba2WyhZ7guWAN25ux1UELwB0CFewi9XU1KQHsbpB7dV4xI
KSvThDBZNkBVOqmHCGnAC5DHD8+PJ6NnbLizERTxdcACKemESTtvlGRzV17agGvl
FxVpuQHfvKDxR2EXWu2NLtTHDJzcknqlM2gOl7MVdlijOFJqqx3LJQvtBRJAMbbT
`protect END_PROTECTED
