`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+MXHvdHarjSMz/SN3sNS2CPzMhGIM9cLdLvTdzUhg8Fay0jjYB9SFEx7CxxCPjE7
eiNWsdRXH5y49FZIQMSPNIKC02dJP5WWGCyFHXVU+3mwXbHmGFFoDwyzqFV+1vKJ
2OToRoZsxFWf4Nc8fYoQPZ0XOqUVJWZQWfhVLj8votsMUF0zIw8ss/c5aDQ4UWmD
g3ojQbj1qHVqcHdKOFS+5x/UfuAiDVbVhHUdG4jgMP7D5aqUUhNnTpVPtKBP5iOm
7CfeWjmA0zv7c7PpjyP+lcxFIxnaOW89MnRiWkytMYL8aIBVCJfKPXIr6Kga61mY
LJXLub9APbHyMfoJy9vy2ny19HW6o/KPoEAvQ9JVOTi//W8xUViQrgNvEjXaXkJ1
46s84PdtufvxwD53LjfAOvuzUo27UIst9FAqh3g8U15LENb65ifWwoeEw5amqxd4
iPvjp4Q3F7l9GALKWV+/4eaEpSSL02G3kj+ukUcZkoAQhJdp4nn4v6GpoOc6VMy7
f58g3MZkrP502mxLwCma3+hSUU3VYQc/HGQWevIzp9fp4Hlqi7PJEomcDsIumT3h
zAD/pmsuwb21o0G30nUle281fUhaHTAvxfwDJU2uiW2YE1pHFfyBZp9MM+kNxKey
Hwp+sEokJmJ57fREKtgIxb54vWB0MeeiOXWrgY7kAbrj4z/AlE5ym9ap/ixAikmu
WI0NPBEdWknKsEln+kwBi6SsLPfGJDjFZ5CisKAsKRkB2/hU8R/GweI1CT8vWHhm
V4TfSDIcKbMLUJVk3Y91Av85ncMNPAU5hH8wd8ft3O7JKYHTey76Y6FxOYic0XMn
Ut2cl/+5RPutjNHeF9H3Uzjx7jWbT0vKZGLXJHeZ6RFHHP1/y6P3d0tKOz9MR1Q4
Pbjqc/16OZgxnOzw5Fq43+938VffL+7x5fmtjKJ9jX1ext6OZfTslYJB/mpuPnfu
cILu9VC1zyCIN1yYKNj7Uoo8HnUkJ6OZyMs8YQ+TIsD002uARQs1siauDDgPjR4N
F/iWk9D0SOci6U+Bos4T6ADaUfP5/hNAOjziJvnc5OOLkKBH2QawuKFKb8cbgAST
kuAcs66a4bCdrTvkrJ6bT1xVg1sIJwefu9JUQUF+5AdwCueSLeE1rNE9UU0ptQuJ
aEJGpHgXCGZ9ZLByVVu+CiAY3ysUOyUJyoyq29uNobpMKKt4DaPti2yMEE+vDQ6R
SbzN4fUJ/l2zxL7tLIaWQvZ6ZnAxtEwitVxrCsu21vfHJFpkNVUpfj8nF6xEGeZ0
jSXZvBFwIE+SuXmwydupE9m/f4QqbUiGoxeloFBuS9iXvow+/eb5Mk4JC64dng0b
IhYumMXqX41egc6dxMM8hUePxgEVaeuDvtV0cBExun8a4IcBNTnVS+SXZk4nMrdm
LxhxYvoJ75M1XMA1YtYsJs2j0/i3YiyFB2T1dw12/eYrBSfQC8Ax7MKhLnfDHk1G
vIdtIJWbCxArYaIusO59kFwBttMx0GGyzKiMoVm0Du4ybQMtYPKvVrdBIzGwJiQF
GDJYCsoh0vECHDdIdYcVogEJAoR5Ju20ccPqLEujgm39vOzitKFZFCh8Yr9N/Bph
1a3mzytnOd4Jl/QelU1lIBzDQ6ABi+hdDTPXvXzQ2YRKP/wRKK9Ffx0BeIunSw9v
zL4FQSb02anxps4OI7s25QIPT3qeSln4nv+G74NN6yrIxYfTq2CEIpIxWAs6HQf6
5QgnF4YyqlwaQKjxF5wIRkIB4seDvH4vBIGRKFXgv7+Vl3fBkuvVf35quShSwdXn
CMFjyQyZKRjuRe4JCHKsoU7xy7Ksu8ECUnFLff7DFfbayXgxBT9QN/85x9dRk82y
KN9CInly53x6MITM07MneiBv/aXzTwFVPazpJzqBbbgqmlvzpDKhgo8dDEGLa2LV
jEXmqIVzvuq0Z9dItEH8cQnz01oJeaGOF/zaG3f2YZ30TDxynPT5rYCQWq3Wpmgs
hkxg5UaxiXYM0OXHWWEGUf7LA8ZhqxUVDNMP6DUDLaerQEHkbGEO9Ugz8Jo8Rl5W
9lHhi79gJn/MJKZWCqqkoQOn0ZxQ1651uZlYynY/Eplc7Wq+GJDFOT6uL9hgvk2g
Bzne4kIVHN6edLCFx56wqtptkMR0LHbL1CN14TPvql9eNsBw2nM7zRyFkx8Fl9/J
Gi6DjHrcxr76bQxZ0gALeO77RMx7afdZe0eayOVWTHkbybP44XG2UDQD835fP96h
yQGJzNoFndZ4fGjjPBJ7UyijB/1pxLZ+k5s9NY5rdU3MCHIYaGy6TAz++Z6RdBye
yK+DA+oKI9p6UrTxNuUC+XAD6Y55UEtj+UYIPP1lqtMLb7uMdCWziHMPpfcxoULi
3mvuUVXQKpBLJEfFieiKH2+xr5wVQEEc7X9rmtXYd26bAv6N+o2cFafRrZjN2qe+
coXdTrN175JFKI5VrPgX03EOktzzJHrhdmNn46N3ctel1A6nHeSrIdZA7ph4VMI2
6gO+E3FeunjSzXs869rCQhLqO0gHyfReZe8d4oVJ54n0lX/doh0rcPQXSwGrrgse
71Lwu32bPpUdk21dy0eUQM8iAc+wEMWGbY69gXK+Jc2uqHL8NjCOlg5g5nqvoV4i
CHzn7xIndEcf+D4a/0jWpR5i4TB/I1qHK/2JIwgsUJwiCLKcjKELpGxtpEEYw1s2
7+jJxKHhgZ6V0Zl9cMt4/dTU8oijK4O1N1Rx/UvfvUti1sHZ52jVhAWUFINSihh9
JO9PM86G42BPzCkUSikOtCjKecOmjYUmetEWVC4Wso9dnLgbMsw2C0Urkcvrp5k3
UXQUG86tFW+d1xIrGHSdMiIUmrgE+wDy2tLy0OfuVXzi9CZHj1VD+cwCsZAagcXr
F3CHsgTNqXqiCQBwkp8mj1Ge6zrLJ+lnNDiwJZMEGqI3MCBfaWe77ngEVk16dyfR
3TPhs3Je6eyfishkaMMvY+1vNkJNmuNt17YXWcmLVtskJW79ASIW+hsk48qVGF+k
OB8n6Go6loqvtJw1XUy8UI/WLbGfQ2x0aDa8QE4/OkOJBZrpk0iaEZbFF1TdMi+c
gs6sW49SF/tVE4r7m8URnKZWxmPFTuqi7nenjo3YUfLKlqHEat2+ZrLV7teLeYp2
8T80lauGQ/uJ0Y4QG+T7cfL/8ni4UeqN2sVf9Z8In4yZQyYlmlaEpx4rvDqPwHpZ
Uy5mv9JwlDj3lUXB9LUzrAih+wd+3WPky6yEWEKNfIM6u/JxcB5ijrPoEAQbMIO6
hrdq4UNt7NN3y4gPnn10/9isdZCcxNlAUK3IIF+evJgpTEuyKTSqU2VBOmvkkMOd
llczTWoMGymEhS9uDt5Tcy3buumvRk2gGT4S73wEhrGKrGYGuqE5UqNxR4pmvP81
hGUf/2RXyBRXBfU8NpVbdp0QTfupg7vKhsT9cXA0PMOdKCCXbFp5d+DbTRMMqr3y
i3OAM7BXQolQ+Vtq3wyuacdiAgKzZRMyVVx9tNoSbKjWxOgRcpGs/OeN4qL80pfi
m00xXziSv1zsiMuSmaBvUQGmo405B8b4Bu6cBhhKTcWM245XB5rXK/UO0X27N9Af
CtCM0SVZdPC2mG8rUqtfiyBSUuWfr4AQ3bDc0tHmS9YDxB2nhVUpBcKxYBMHVJSz
hHSKrGw41j5u9TpNPn7wr1K4gdaHNOvtw6cJ65dtxQyUnNzfFxDyI+t3LJPpB5Bp
1V1nnqRNYe1tfvnOflCrT7sQu7rsylOtIE0isHfmlJEchHKTa9gZbhZiacY5HrYP
YPKF0wpvT2shmHzf4hSlLOn0KJWOp1wmKfFSx/V5Qz01tauuSWZ5Hth0Jo8rlCy9
F1nHM5/nPu2D7xWhjB7sA6d6LgGsRWUcuZsO4bGnKlOZDRCcomlPllRyoWN6cjjh
IZKmnufwC5XaXh41WtCBhLbZozOjieeizuETKbVB2s3R71NBp3sE0BW2DxsXcAne
2R8Ze4mrHkYgM+EEWHhI9t6PfN43+1cLPlVEge/y7zfpdtOQgNJERamz3vWbOGo/
4pkdhkpwN3QAAwjKQ1UDV9moqP9WzV2U5jKmH0S6b58Be/bL1LEUMfyTVTEVGBPF
CsFA6HAHFo3pk1C0FqPrtl/2bXI3mQuRqoo7uC8FgtORROqy5Moz3NItrxSyspXu
V1m3Ev0JW76SV0cAhiBO3DWZtUl9k+nKEDVwT918Tl301an2LvLY67ml+Sw/DKOZ
C0lQN4/6eGNmKkN0jeDtDM2wq3bPLevPz7KMGEG+l0W81VHHgp7jTEM5YGw3FN7Q
vEpTdhRzP7+ZQ2SppjY+cN1w7vVKzidG/MeZVCrm29URDCdkn83ay9mxXSuXoH0w
0OYwfLOeeDJS3L4lrph8BcYPzphaTl8AoDMiOyNCoE8FHzo9dJmaOHNW84DMZdYs
LxGJF+8kEk+rxYV9tA8mHI+lYgCTxCCUKQAnePm8vMgVJTW7atL8qPtHDvYRmfNS
ZV/E0d1SSLmlInuNeMUzDSpYUy4pCphILYfzssommXhKs8n6RNMHAiPjJOZiEa8N
x8tr9CJtrRLcF3/67o32TBI9b6mKvncIVsz5dyaV/olLE2b3EFXue1l16n8rDbuT
A7G6aI4O72fuxkveZllRX+nK7cM/BjQw6gXMZ/xq85svEC5vdq/pq2sgnO0q96/u
PG8mXFH9rlAv/rn7ZkauGG8T61YUIQb6ORo4ADqfJeyNaTM4iML6CskiZAdZ4aD1
UrzOcQM3nbYi6MsWQ3KAskf9LYhBwrzGA6sr7MticFeFontJdhXkUQDb1qSexNYP
gvVge5sWv5smmDAXagO1hcBKzl+AJRxZnqIa875R15MsSi9VEFkRmXVhC/NI3JZT
A1s5MH680lpjWexBfFuQe32naIN2JkGPzaeP2wqcTwIw25H8SLhdjSnrjGMxCfMZ
0sdvXyLtIT8Liie0uUzK4W+Pkm+P62ZyjEtzf5cPt7eyerJfxUTBPbHD+PqIWyeA
9nilbGnNPewfe1zpsNbClyokGEfxZkkcsbj67w0WScih6gzdWftkiodW5hbmIHKl
10F7vOwaww9jox5LM1zeQQqo5d9RUgBgSkpPQa7lIXjfldg/A4gE93aRf7evWLc1
gdL/2BngPTAx4KIc4q31F+I0NaMXpJp8keXLGJBy6NUMfghIpCqoDIQ5u/gHcGQ9
3BdOMdOrJdFh8QnsaTBrpz43Nf8LzY4zct/ikZWVNHDmW5NsBebK8HHJYNDpt6y/
qEc0RU2eXebWKplPeD1krLRHyQGd1iR3Fgmm4pHtKhDWL/Q6TBmi7/Uz95LhzOtn
MA5lT+RfKFRAUfq+z1GVeqoxpzGFN/o2CrCsWKTN2vZWD+5cgQHLIXmVMRZjopJN
cCpxJrM4Z6RNO5VKln0+RBizRVpfyUKkOUX8wjkeDJ0NrascUMKN9BCeNucYneYf
23itshWM3qiBJv11dwwMVFmU6dK93RiKZuf9diFq7/w4yVHmxwbT/uwWyvElEYLN
H6ZS0v8yzWD4/WZQjeJdd0jwcJacxJz9ogbxMrVxI9zTaHl/gMuswXb3a1NrUkwN
roAUZ8PaQMFwr665FZ7tMmjT7DXM0x2j3pkqifhFDoYCgp/joKCGONoLxkF2/g7L
O6NrCTpdZHxnVSC9Gf80okwX0W8rtDYjyCgChrDbk1C1DUJ+ypYM/U5HOE+vZ6E8
djH7WAnXCwXNa/MCHXWyBTuyTpUpN7dCfVM7aoOYMzXHc3VlUjT5eubsG4CqJcT2
wKu4yoSrGNv7d52rih3t8NrpU3DdCi6hzvadQ/kM+EZuWBiJsahr5Ag3XEW1DiRN
e5+CV3l8r3QThoss5vcVDHQkm32ROTuxc/UEvhDbdgOJ2voRR9+1mR3SinLvOB3S
IdhGkz107QOGdqlDi5ZzPC4FhGCeQBxo7n2KXbLmvi9N8E9TiBgNvp0AInPPnWjv
zarn1lGiv6BNez/gsTUJE3htmK6GLoVX8vSsG6xx4tHBsCcrCMIRjNxrEXD+9j2H
S50yw09IIpyGWlatmUfZT4Q61OeG7n/AREsTBMLaim4jkVfpLovhFIFo4mRTCep5
HHDsb2EoWH6mUKWk6Ca+8Udmmr9kMzOv+Y1Yj+OE44y0UF+8mat7UBCZDX8ZeieF
ydLwJhx9MW2G/GAtmkm/tjRZpvEp9RtYvMMYWNAH6sgn01yqR/HO9bgEV6Tuwa6S
CozlByVutHno4wkvgLjWwjHAO/VvRFkzsy0brON/Tm5YIWta/kpgUamYwzxTmlXn
M6l2NzSHR+QZOJXwBi11QQNopl8j8Gx5sNCTpQKu7B9Ga7eL7CmLU/e52LvAFbyF
9hT63a9/QdBIW7riIlLl0bzaAuoadkRhpu1T+0OJ8BPkb3IckvnlGXRy/Hr4Q8Ab
N5dvZIERuXftREQLSVReN2yACc3/cLdXTIQFhQgJgSa3ZBTIwK677sHMwBovG9e2
SKv6PsgaLNegzqKdYJuJ5xRdX0UluO3fk9FlMwn/SUhuMNWX20LcZfAo5FO2hliK
pU4nxnD0Dg5Cp5R6trKKhyg3XAdFbvkMdL9G+XcJRPe5bx0JyrhPBEVCctLlosjD
YBvgny0QQNKumVDU5VxtZR6bX10o4BWffrBsnj+RVoyONTiKP5PZw8umXzSui5za
tkEHigQcpULM/YtQS7duM2Uk4tSLtv9ebcEYRmESScXTz15Hsvj7cPIaPpjF+26R
jjT2WMu4T2DGAqNshihPH0+94LggvaMscORyWgL6CCXWnDot7XLEEG7jqEbRyRq7
YLqOWFEyxHN3xuLI5/jnMaVSqzQ1BnCUYsT9d09tABn7NOgexehUnZkP4YKGpYCv
C22qJ+vnt8tbXUPc4vFM8fhSuCE7EXtaIABsEnWVsjOp6mqmY9057olI8ovmQ3ew
YZsiCnqYyjrkk7Fc7kFPmgqAqJyzGf6UpVjLbX8uQClJFZ05E8iYXyf3FBzhma60
HbUtSRZYd4mT+EGhXQB4Rt1xrxeWCCJ95VNuiY9h59PQ07HEY2ZRZj49hgBA0frh
wULX8RGJDxBcBwz1VoB6UkKaxlwqfatBSPJggaQkxiPI+pHRJrsaZt/MgmaL7xBe
3FpMpaHHc6eocMJLCkFUtcEgcUwt7Y6YKtfTBAg7nHIwNGKUX1yHQEE9w0xLV0yE
vgeCcfocJsRmpsc6NUygKgUOD/zKYcDEe0Zt9SNDpF19cQs1XwZN8Krz2thvRVwY
nrytcXpBL/RAUxemgJCdWYZddPrtMwgGpM0tXV8myAL2YqDS0ffvJ0eFmlSEMmWF
F+GJMlZiQwpk+leDkoZZLj+tGDS3VJzhdGfmzbAbvm7uvlUtsGe1AeFpuDW/VoQR
4TQeSLx/IsN6je/uOnU2T8UXD0K2k0x7oyDsPAosTlUrC0mDtpTFSBkklpK2iseZ
PIw+aNCdZ10B+AECqLRX4O2vglwlYRkJZrITxnGoz60hL/q3ttFpf4z5okZPYoAc
uHdgKlHAF7OSEq1B3sM3+7jQCOuVOg/26XsaaKKoOfd7EIz6Q5nwTf8ZLBMKMalu
wMTwaDGm+6RQhoFj1MoAksQRscz4YiODtWL5AwZPMWIlNYMUJZdfmCIt1JnbFI0s
XltZrF9sAKlOQgVdlSIYl7DXd55V0a6mYib6V89rRRbV3V0qAd0WFmYghkf0OCD1
duVZhFmIyxDdSP7kraRZbfm/Qv8Ras+Ax9pc+/gTBssMrt1aLh0gtmQTflzIh9cB
8NX23oafUeZdg1nyNMCzxV4YWpOw0w7HYeCl83EoLMAYsCcHVHNosDxerpooQr62
Unvp7iFGadTUfDw2wV9abrclbFZLh0PcOU2C5E8Ta0FcOWbaG44j+iWa2g1KjKbN
Q6wb/6K6//aQVnrkuu9NNZkjWIveyi+JwVO3D1rIoQ2muffgMqMYVp0dZJHTFDwB
UMbdI3eaq8Kg1+Yq/hJtv68eHAnOsy19w+4VrL+IlvmVC9V8lnRaPtbgfhqTmblp
DjjWQCdpxna9KsmwCPDAoCLR0pke+IoBWOgcOyk+rnLpvDcld2nejfzgZZ3/yJm7
2Dwtgwaa8Yl3FUXvpjZee2ofMMKwo5+nYdSa9EnN9ceWP3a4Zl+yeOtwJ1qwIhka
HdqS+ziKGealMWChaqrDx1b2vDX+4u2DmDjK/We4ZiHP+jc1XOG9lviThXyeS6LW
NcewTGrELojLJVI/K9JdAOvEBD/pRBfTVKI1mufvJ1rZZQwmCHpH3NGEEkaB9ogo
GRO3bEUgMlxPY/ke7mdxkhO+xpNk9EdILmfBvXGvQMX4ftLP5cREi1qqeJJqH1Sk
W/CbKGtij02P5lVw4zvkfgamlGpq0XBlplXsbFlDPPHEMlCCFaZvE35SwBIIJWv+
lYc+PQqZ3oFM/b0JK1Bkg+hr05tLfeyBLUe9ECfrUxgEKiAKe2tQlpw3AkATrAN2
PAX8pwT9pRLlNkGj0vLKgNsS1LRXBrahAJec3muorONuVMMrtfD7g+oMFxgQoa65
A9VlTjZJuXnAY3XQIn32RjlzUlM7zQgQ9X1bIfkUY2lWPyLdhwyVMPb424lLbHKl
PplGeldFmSa5LONzAj+O00VDRcTgqfSmr+yXk69eJ5IlO/JYlScSOgca4a8qSdjR
l2jgwf+zVzxPnN/DDbcuCHpYGrmQi13E0CdB48rj433lh1eMOGr4EbbN4oL5fcNt
w84vMS3TXxMgM73P+nxF0x5BCtVkuoZiGIlsozGI9I6m0hB1IhqvYsbf0eR5BB8C
DR/AqKL4+NewDJCdKD2eZALUvOW2TkK7gtkO+O6VbI/z1cP+rAw8JhsjrzJUwOsY
MShgSSlwGv7agdxDxPQR0/r+tQnM2ucszPPphEC7AvfXjt/5iTFlxQBpC5mma1+k
MmCq5qK7saljO2nPspu3/9jLo+1zv6OoN+Zi+zsUzdg3tdcD6KMOzj6KwdK/qeJT
F3H2lFlDuCg+BsyomkG2s6HmIEyNfTFvFSIGxwYtg8AoHAe308TO6NLWIkdV4RgW
4lA6G1qsOa4Sv4WrEOSUsj7xYa634IRjgXfsLMqCbE0GR6/6gzRtUHkxuQT44+2W
eP8/c+LvgDdh+S6IzQtPwbiHtSx2THqgSCgtd4PQpHRK/RbGjb9OZtF37gcl+6ES
A99/yZl1or+7NrOidE8b/2r41I+dcjGjxaAFMM0dxBIaCFj+XjyHB8cYQTeSRwJC
qpXLera9mW8wav+tfQ72OHNHUEQzNBhHPgUys0CUOlSv0Qifzbk2mj+W0xkDHVM7
n2Z6+sx503YcFSXDI9PbtUdNfcQVprF/JolbVTmMJX4CGsWCh8mrNvkzr1Hig+ss
FqXsg32WAHJlVKQjf7yYOzlqdzUlkulBVLpa59xpQHKRODl6xXQfVWgArQAHDCSl
9Uo9FDk3i/soskY1wZFSSr7fMGVq6+gTADMviLygw9d9yxDmbU5vmthNYSv6s2NS
ZsKDn8tZl8SPGBIVas48H4LjH7XuvoS1YvvIVcho9WJQng9rpnnY1PnIWiOvkDdE
Za3pqPFq0UBqbVpMWLXbBKG7Cjin9IDSaTIsP51cfK8s+GW1LYglj9B3fPcU/SQt
reIZtNX+/NFOKPCHp++kyVRlarP+jYM/nmxoiv2m/Fn/zdLlWAGlogkX6qBSDX/Z
eyliReTKGgqpbAXV878VmZBqgmDgdd1F2wTfcuUiPzY5SQfRzQ7hczawbuag06Ez
CvbM8npModS3v3ustLO1g1ZcuS359dCPzKkEu8wqISKjtr6bLD1TQYg5me2m+DO8
0R9XJhgjsuPgxXuRPyzbclfjsyE3DkdTyiIt0ichs4dy9cMgko4kMo8YfeqlZVYQ
C5fPYdTq/p7anZ/0ncSc2tckXyHvr3sAlL///1AVRC0IjhbHItIjLh2qT6gfuCGQ
Gr6JNkkENeq7f19Tg3M93FXM94YUQklapuu+r9Z+5b8zqp3VsCv2HB2XD2djZxYt
iGfp12MViTTdPjpxZj63RthpreFPrifEl6o0yWZymtL23UWp8MQAmlmjleG4iR2c
SDxXXPM1Cxlg+igO5vYRhgSN0+sxVvpcAjF0GnfY/bquvy3xjNnlK4pbnezRI7Z1
1a0PCLE/Vg2z2bYS5yytCHJvFB2x1if/2qIEsFVEjerY0exaOUG0wACMr33PLQzv
3d5gOcj832bkUrY1ZPV/QDzJZAWzhfN80eI1qUSceo1MmtXr3t5lHSwuCgxiqKOR
snDMavOqmfwzatcorzWRFz7g0goR2/ScNySGB55aJRmT0O6HffOrFWXndJW3YKDe
LHmn36/CelQr9SDCtGVOYHTSmSPUiL4muLI7Zq8xjx59EpNOlFZ2j30Dn6D6XZlP
IBLwhSiZl97Ba/97setPCJBo1ehZtspC2GmnhbN/7c9b+XfYNaY+DVQYX1wbebE9
7eauTwKqf06QS97y1YDKd+8IKgcSPgmmgCgh8+K4QD3ItbPuYwG9JiVUGFxuXCPV
JPqjQ7vNtL8jdQ7TCR/5J4Bhzx4yItvY6q+Rk1YlGv2yWVk7HJL5+MXsxF/2KbBp
5H89T+DeP3J5NJZOqF5QEa0e94DPLy5rF8oxxWthTrzoErPIkWVbiqOyUe1+qZ92
p6lLWk2EDoQsQqZfWLDNuBTUTjBlC5c7SvzaMDFVlLy7ZzKIiOPDBEz6FpRII760
i3eBpNagSXcKY3XDKToFUlLItg8njNf8xqmorx50NhTwdDAahGsXvhLM5LUg91U+
CsnNxC5ZxrN9L7JAYX6pJaTU1Vt5Yzh8+zyqJuc3u8usmbcMFTwK7XOGssumyF22
SpP/y2tU3z9kMz7wYYMEdRt0IFtW3JD0yoElhDf9+l/30h1Qx9c+w+dOm15V3nAP
BjSKaBM/g5ulghbMhVI2OaU9dRTlvF11OJWw4BRa60J+nzc7mKJMaNi5kmMG9PKu
zLgG4fZPkuGL8WJsTq2dkffN2DDJq6w33AZqgV1p6EEf1IuTuXjuArmP+u3ufGrm
j8FOpMViAHz6DH8QFCWMRYGJO0VkYyK/LKRqUi9XQYAVGbanQ6vAvlKKGBuNUgKI
WEZRcHGk9kwqF3s6Q5RddN3H3JCt3ikfJRP85WpkJvBn+y3SSifOyecOBIML3w/e
624myx8ReZnjaR+cmaWWmvMGC0qZxdrAu8NoCdC9XskX7c0yS4kkcZjFDeySeYdX
MxnKa343PAkZ9y5MQpIXSrdmcm+bqHjsw2oKu49o8rq4q1jNOKHAtwSiDXdeoxQu
OnwlG5zRdCDWf8vuBhaPKnIPtjBvRddPAkSxbKd5ya/tRHpczY/SRvzQgtJjxRYU
F4N9+h1yrE7qv1n0aapueJfqdaKegGx/Gd7b3UNMVfNSAjLIs6bMEHYLK3wuZzXG
gJv+sMMbhz9KFMtSYk9GwfnkS0/FcS86ajVynSlNYgn+1VBxllZ3SbD9Uaxodc+F
xHJEfp859MlnkIqPo/VwDMrdLhhE78tmUx0aEL6riPz9Sv13UgrcWVu7n1BCMz9I
nObKd0WKb4Lwb+uM9WTm68PVhZgMKR2OZP01dECq6LvHMskWzpp/PhBa8yxqUau9
efERluB6SFEB6N2EDMEIWDx6UlN+7fes6x/9o3lVql1U4o0CQb8/LrN/mywkpYL2
q6vbx+dQffMUmwqXBSrk7UM4+lK2/HToGyvBLMt3EPv4AEbImpLXPhBKD20OuKRg
RH5nt/98DPi2c94W7q+zZ03xQtGpqWMH3TPU+/ce8Nuyn7c1wTgiie+zh5YsqbU4
HbMEFC8Yem0aw6IDYFIC+sPzI6V62EzRTl0rxQ7hnDMzk5djCr76oqyYYvf/glnL
2//kY9vn2shcEm6YE/k3Wh8AS1XYRLXxXAeKaDRSKrhRCS43sRxK8dmfKxF5p53w
sDNhmjduC7L4RFp4rDUFRLbbtxhs/v9L5tz+cFQvffx/aumV67+hMmQ8dU3oYcSC
26/h1zavuTts48eOzX2+mB3ePb6J9hA2aaogLR9NFRSUlPdKB/qUBhj7sIDAQ51F
LoFK1KarbFzZVPlfvMCyR8VeNBgCbpAF0Fu0gDIbZ+BucF2AVPOIVRBc4oJI8d5K
dNWpHqvC657iJVoI0hAxhCvWuQXCqM8zdCA5HmphxJCgVud28Xt5rkhNVCnHygR/
CIIteDZqhP+vP3AS72h0RjY/4Sqeef3ertB/pPrzexG5qzl8EYAYzHnkahZ9Vj8B
tYfNRK4Dx61szuL0bmM5PM+R/IfqwrbSQ4oSSX/tq15x9FRY0ohTD0O1FG6oaa41
39Wsf55PF5TF2VWLxuh/6ajpkER/o2tSbOYGJH0tmUb7TQ86SX3QZHArU7sCnx6V
gWGud7jvDvT+wjQUF8lNLudw7W7jB6ZEC0TTO0aOrHx9JNXjik9n7+Op78fiwPQZ
ESvDzxv98uC8BQ5yZuW8uxxmfT+pJN11VAPZlLrsjCiOK0ZFmYo3IBM4xHjoacNU
hqsPZR80utMFiuAT4Kzpmp+5bbo7MCvLY/V+GRWRfpi0fO6f0PAsUcqqAH8jjKBo
S4ccsXgOVwnqv5V7xpj1qQnf/MkjaahOL9omP7+az6sJBnSl4sxEcL6wqdpdMy00
1O4FgGDU3+HAUZayM20zyk1mAm4ChXgtTnmTKv1YjyfV9jjnvMvdGJ8wwsYwg00s
YfN9ie5xWdL48w0KGvY716Iv/+ZIjkjavNQaxigp9o8AdNxN0qb7YsPZGQiGpdOL
cmuXi/ZiTPXald57E/Lv49sa+nMmEwWRSLi1jOwdG0gD5e1yiLEXNyR84f7wxYo/
DpXuBdNAuPu46DDL5/pax4X8wPRWIcfaSv3PCICEWDZEyOMGDIAdleuOltGbkVCX
OW3Sngq5ujDLGcF6ZcZkR3/+Uzp2HOLADgaiZhiZRJR0NzuNs4ZVPAIc32nFJS79
pos/MT2/BbwGkenXJPUMXlCY+92J8WZY+4xwVGqj+zxAsIOb82VQCKcTrgU33u1S
sd8rdiSIq7EtUhDZuR9pRPSvmTvKxaEVOY3bOmGcO2N/26xAGGw+JYjbT5sswUd7
FjvNAf2/k2gTbPFChhHbv2s+GN66KxiKlmbOy145ofeb5jnGIX/SjpIuBmKmctZV
ag89NJVCK5rocMndD+ynt6c+4EebtHQIY8Xz+9rqkXAVzz274un9woT31woJPiXo
C1W/e6GfR8L2zBUN42ntMwLOlyxoGUsy3dLEOWJ1Vww6VZE7iHq1mfA/fdtcx2m6
HACNXKGQVYcseZ0BJaoqd7PsFPxEmsfjxkOzELhZYKzKKIsWBpbE8dhDnlC/nv4g
ZAXRE8h4iQD92RGix5tHbVO+fgncDA0AR7SI61uScY4/an+RUr9Fr3P/jlwGVBzq
DXVqUzpg5FLIFxorOQYlEpkQt1wLbnSfWDHW2mzIjZSvd2VLfeAb6WN6IWY/TYTc
Mia/Yiy8F42dJuxSqtENjEHXsUWLcD6WnvaIjT/AcpmRbnldQ6OPb1YwnjgEfBPa
kMbeOV3fAFQKXjPeTvOzvqPIGkwTR8ScjUJb1xb3zw4olpLE0K2xoj80o9+vR8Gn
SmPZ3dly5ofMR8pqEeys9c17tzbqy92ThREwH2rQv96OTB320m3ZXb26ZvSt4iHl
5U84OFESg7MmpTFuTXFw+6Aake7/4P0p6A4meqGmGMwa4Tcl+mJ2qyKRFQ6gWFzs
57B+LL5TydQuPSsm0mLMdZbNyOeodwyosCUrNn8hCPWxQ0mFuhIJjRpfx0h7x9cj
+qS7zXjcpViw6nQ92B/ZNIBwpHKA8HNDmj9K6hpSbOlE8kuUj2bN1BP6UdyykX9K
Dxb5hF1V+fASJ0KwZsGw98tS3qE2ghJpW3VRedzxYYI6abJMet/+M6Uw0iCf6MSH
I2tlu7+HQjdNWbLjlqlgCEy6dNmp0nXEZ25t+3X2s4b8rTpNisH9Ql9Sa0XSt/qr
OOQ4nj6zSXopgy4vx2eyMRWPAtmPL924XnEC7wgoPPAqJR+08wOnS4hwpCWfb3UJ
3QDXvDQ9E9rmrXnzC90X9QmT7JtVJvkR3DpYam1HgDYA+6dRgjc52fvlBaHakSDy
15/nsJNykvWujv0KKefySx4bZAGlrUkUFE9QJlDG5DUNi5FMfenAbaN9zh/lT7NP
cbmLbgnCngiKnI8eQles8L6iGP+Hn4rK+lFsdCTQgEvoh/FQqUuLr7hwj2YjwV05
GavNi+GWT5bF4r+kHE+tdPDO1MLSQD5mkQY7DqnAKIBaPdFdiByj2lXZX/kvzMBr
sufhSaOl3M1L4uJTl1C/Gn4U1IszSXXpFrlM6Fujoyh6o/n0lpYw7TWEV6fZM7IP
Pt2ur6REgX0aOlYAWcI3NCYcJyLivAU5EZCMeh29PuUy+zekbX296+wtdCPeD0/s
8DJuV6pePu06ksBwjprTE5k9UvDYNKwUSZVAqKIuNI/I/8APi2qmjCJnsa4SYgoO
aSfBInnJ154ge/hA3VtiUiLF3ht//hIAUV5PgVer4RmwFW/PcfmwsZOukVbQX/5E
XHQEpxgHX4Ko5ry86QOLyNkh+3K0M0rOtjacO3OHfTQD8m6QVAkVV5hunMwtfp9l
3WbQJqldaG2eU+fIEtdPVjsQ/giDzTUQPyQmZpOPKuYP0iTBdJ2SY0GpfpjXMYj5
/r5NRgWLNt8ebxXUorj7jvW04kgA2mKWNRADhmhxPKFygjORGBiuBhgyVnt6CFVW
MmtSGNFX6fmqSAcfSEjbvrhn+jsc0Hr6lWqasGfyTusbSktqXtPD/+fSUgZyrRYL
EN+Fv3V50XBn3URDOUCQtod991+7CKn8G7lC7wZl8tVGNZCPipWyBFTTml5ZSyz/
/UETFVnCbZTq56eMXTcBBZfgIQs4l6zra4sTwJfNjGfNPzo6BuNrXBkRDv+HnO+U
MwFkgejXGEc4wkhXCL1Gxh5gX5MtY+Jei6UNGY4WfE5VpmwG/2B0Ov9jXwUtxYqw
KryUZSVXQI1NmHFRFggSDosayC/gFp4GQ/sYwBkCpWh3OMtscbD4qJLkpIXIfdmI
CMUoyzlygRpZQ6opznu9G3oqtALlckGrdmbCWpACLtTipzPe7zr5Hj/hChtGhLmy
GqL915wX2bFrd/kiUacrtOtOjbRhlxNdvBulNghg3FApSw2EwET091i4/wcxijpH
eh4lTrEQUg5jZSektJSDyvtNBBUZaXTMHeaQvnoRcLK3fbKnvT4VKMVXIIPWltVF
bW6KEP1sAHnNNN0vKBO3EntDkZ0NbPO8ky51s0PnzPtrNnJ+eAGouswOhoF4K7tW
GoVPdC9yWghtKA7NiPqr3R91vOcmgF94H9MDzg8yS+40/flg1iAQNQQ6K4E6o1rH
WKYdLQFgvdLOOJuOcmDh05j6/oDeCCBHpnhEZWZkKLuhm4+7CiV/ouZ+yE1IaHMR
IkHLvozGMdgy2NyUksWvLMbiNd1cYtznFDX1TR48PExHFPYDFcBRdMZ+vcwRl2KV
CGI8w6zRMFKweVeDUwYZ0BbkHg3k0UdOlfUAbhNx25nTzG51iXutQKROVBnjsnK4
A/mKU21JTGjHdYf7XlrlfyihNFUn/m4FclewiYe1kEN1Ppy3f3qQHnZIJRNrTEwd
B90ZqfotrBWUktFmod9rF1x1iAVlUoy3aFSOi3ErmjzCDRESjKF68Gpfxd0S5Ziw
cU8xO83sLNdxFcXObxen1yqUx3kY/eONhD6uZnLq2KrXgA+BEC1E6/kWqRVTB4Bf
ixLXRZcJRIgkEhLQTlJL7CZhbd7KdHV28md3I1EoQeSGBZQ0O1yRCQ03P+R8ODNd
W9zQkdqA7DsnLOcz1aTJz6AqNl3DYJnXqOKdOAgqdbNQ3kFPZq7lXXfbJJama4tr
vaDqPoT6ZF8FPpWUsDCSwcu13iajk4V3OieSveaj54RWZmcEhpv0BygLPsg9ZMd2
srAikKCZls1mzXMnlX8ATIX42su3fAT7CEMWhP2jNvKM8sCPB235e6ksuOhs3ubS
g4ZME9Mi6SZhxvmbaez5sq61FPPKY+G2JdWfR1IJL9ZrSKMaeVAg8h8i/eM5Dnwq
OGbY4nDrrSVwZmRFc7NvrvlcHoIz+JOXIpDB0iUAVRDRfkBCaaY2ZLfX1UC+OuKH
zTEiQSpMKCY2d6qvkNDJUgjMFwMVNNbYiV+Dvw/zeYbEGCNAi30mFnAFu9ZYvc9f
/kuOwyhCjTgVPn5BDkjptvL4QAANBJylu55u1EDR7i5DXfc+jqG4SWaZfv1UasA9
aD4F4UYg2PFVIA9o8YxgmbGmDEBj+0h+dnYCVvBdLg6n+nyC6T3F0WTCJ5W8lCsb
RcP6Hnu7yQfDUOlsvYdBdKkl4OJUrL/E+0nsnjXBx+zVt4776YYbxChCFnFMCa6b
9WjOVBhEr88uwdYwGCfRE+tGA9i9TBiTw1giE4tmSu2Bkcr5hCYcr2+kN0mrPRDG
imbPf3W68vwG/D2ydMnMzjnc2w5godjtVIzulv6Lp7RV7trt9cd9OwP8xfE6iM8e
CpfMDUY2hFcYDBpMROnnkGsFMZnAf5xq60Am0W/KS9KAklElsfqJt5sB6E3ZOewz
8X3cy7QlfbLe360kBd7GBDEFK2NF+I6KF6bfjQJJOAo96PPPocbkRimgIlu0ZVld
wTDMO9R4nOGy0ofXzJTzEDyzRnhTqx9exGqoBmmLBZGjESxNbU68xQuiY3f3N4+Y
CWR7k75Siof9j1BqYWNKXx7et58wU7Jz+N/46ri8sYnsDpzzYFeAbrofZdIr0d3R
/X7ZCKNx95CtvHrnVwSRNRvtcV0UM1wrLqLAgnkHCsaIJyCkv4+xWwGuGzrJvXPu
huVcnKr2IzUaXy0hcU7FAp3s99Zlf/5craoFoYTBedUGP/fU16ybBqeL/U3VoIUy
2kMDnWoxSOdajP8TU96UzPRibERi9xXL6gS9BwsDaa4+yItAg43Po2qwu2XtJJEA
XAXBqN02AsXXtpCVmvlMuws/eSYgyUFuhmMynWwFDU9dqncf23UOY6SEesrnyFtj
nqH/CBy5Wcw6zJ1cvvvKxCzuC3MA9meoMB9gfvL4KVfoKctNs2TytxajGT8BlIuB
V30uDKyWRDAwkJgSwGVSVcyS64CZisiHnlR+vMIQRMVjoVR9WlCnbkRuMpcBY929
O5FZ/VLEPxLuxHeJrDjMR5qUX/dWb/7Yvq5snrw+qLjO4WRTK3uiXq8kJ1TpNmTl
UQjSBqSh9ZK2lbq9H7wK0hm3BdeNv7HWjvX2vbRfQ8nQ0Obf1wi1al5juHhM+8+w
RYlPYYrejHqJ9iUkb+IM6MkNCYHgdYs9h8TKszeK0MK9lZJ8VYyWBmDrDCzrCh8G
Rq1uVIZbX+NalDZO/XMxaYED5xTP8gbBBrvCw4ywDKtnPWZ/8+wXHX//DMvQowM6
/fjwG1ibU9dY3pqFPETUAAUrA/ryx/sW203wgtbZLhMW4uVrcRKOmkV/cT+JRwWL
5Nx/ibygpOTnumULZS0/AnE/nEPLtUN5D57P0zIodWYRv1YE9rfnTtj80cuLyzi4
uaps8ZgXJ1aDeSYB/arPUSg2AB8rOK94uCr12YE9TOKs4L+lZv3gL7TPPAtK3EJk
Moq7mjE9Edel2x1tDUFH/++QBpOCJSk++0WSxvR+l9Al1B8/BGu9XjNKJnqfRU1Z
DaxMWqdfO4kcDZAKxd1OnByLut2GmvBEk3Qa6BSRQNKTBhymT6a52QlkV+jpBcfh
4mThDeW9ghSk1Aw5ZxLJXLgG57Z9IOcJtr1vWFklnSA7yEWjvFo6vPZL92LKV5dE
nAzEbuCHB/rrM2fiIYm0vyUgpflU7EF12/JNmX2/H6Fp+Op6EuvHXS9iPVPq0YlQ
cSZZ40+VXWMeiJsI3ScHFUS8gr5/50RCd50jCUO/QTUlIkMPpQrCbu7OKaggpiEo
Tz2wTeYh88PYr9vWI+gpJw6jH2898H2b0iJ2fragNdgQzcupWUAt9kfcp2mmI8ni
X3UA9lZsT3bGlvgR2VcbFMkEQgTDuCtuS1xUgZYcE/lJzS1IMnDXoGH6aQ7fVAXO
i9sWZXZPHqi8AmpASixfpMKk6cLiNR7EBFEdFM7yhLZQDsQ7gTrptT2dCjAK5zbh
nn9SCMN87fWkHYemwbZsVc9wHOSTCOwlfCPUvE8W8swNzXjSyht4trnv72uneevl
bK/OmU2B4GoEA7dCg9bxIWBeHKXB27FPbJF0N++ZG6CH79jWJQZd4Kt0c2s1FeF8
kVcXbZqqpj+pT8s5FAbDfCDbGd1fnovZD9RgxXOl9hlTL+weGDTMyXhyQM4KaLpi
8aUBp5kuIEM7+AAh+sHpCkKwnfBLJti3kOFU3Cf3ETnKiz82Wc+/PP0Mo/IPZR/4
MQxIs24MG2W2wf6UheCWZs0mVX51rnA7ZueIBYN+y2FSNW68y38tIYusZ0ukjXmN
pq6v85EHc+EaYAR78fQ+F+NIj0ItkwutP0HlIXGuRqnRNqJxzPcvrY6sl5eb9jxd
IBNMK9pq0IXFW7F/c/TaJmYrnUOir5YXMjj9bn6fk6UQ2nL0IfqMmdw5qwxLkh9j
p1f/HFIG1EAE3q9lJo0/nno/X4j85UOTp3LRjTa2BWk711VXycatA/LiOZ+XpzqC
YHoE8Umtj+m/L5KG2fWlH+w/EyRdrrIVggKspgP95nn+9jp1amxY4M/B15LTWt85
f7NQWzIpKFBPz8+rAnP/GCSm/BX/dlvALnovYAQ2L3N6hfS67LHDd5g3hbVER+r8
Am0MsIStpM+i9nVMUE6xrvrovCgvn9VjEEYkQNjHpMivYQlL0rNB+nfC7j0eSU3P
FZTjOBv3JbijzjAKrjZPGu6bWU5T9DdKg/h91rJlfsEzwYfOGqsaem8nJohNpdp8
FJEXLsSTT+5X3J62bRqcML4oe4WvWiQ6ZPdBHELkmt8xqb5knEU53w+VP4QIKnxs
qHnHJnCx+4I/MVPBjJ90l+dnYuBiJeokopTZHgdPpR8VgGb9EyejajW1TMM7DDXP
LyqUbDqUoUXCaMd1MqwdoeY8oh36mq9tVI0lsBZjJwX8bRe/DcBD1tVZIcEwZmwO
LNxES6aX44SAEYzNNyoYBbYHZnmPEN08RggPfIUmzR0woVVOCEY37rJNdyruVUdR
BAAQ+PRcx9gDvbU0BycmO/gjkKSC9OdHtP8u+8AqDONmvU1WAJed3xQhz+LdJV1R
kAZgnbwMgSnJ3+SbEDEtF2Xymmj79WHF/XGSBvS6cyS9yVCeuZpcXFBWHqQBaTEr
BhfjAPTkQkEEen/jTV2++NDPpW5obWfbrCEoZtYw1pNppDOy4hEJfqBTUg/41wpF
vialLkXy4HMwPCyQA8ZWk/GiGpM4q4wDwTBWRRxtdQkvuy3Xu31E5GMlp6l3Vgvq
b4FOxVcEf2jSJM6pwyxOIl7UR2sxwvD+HgPxntsIvzNurqmbZu4l+YNEv5NGtUyS
7aU0tUAUDUsxlsKG1lH62shxsIjRql92QccJwtmx0i7nz/1tFeul8Kw3Wr1dl90R
vxeORcy4f5f5YW01OdGVB/VUDrKdlxKvCKPtxhoV4WpNIYP3i+vZtMlXehqFwt3/
yHLVGljzfKnBf36ffHtDPKTw1pfHsBpx4CMeX7M39OJKqdOKmhQWNZaemUWYQnZZ
DI6dGrIKssDj7xCnE5AXBh4q9Kzj+dcMsIWr0rLNSJIwkiZpCuFpHcKGI7uEff0S
tHQPDtno1thmvsrB8pJI6g67v3f040iICwbef6LYHcv+5RmOcuxHzdCxR9+GZ02N
bxyy2bA7TvkF7Bjs4l21/0mEsRFLWcSFFQt3oPxRinjSj0vzt7gr8mJve9dO9yS0
xnerCg7tGS4PEBBUWL58jxiMP++0EDt3YZMT1Nn3ftSfeRTvy/0oNYHj+koLMS2Y
YO239Ritf27/6Z/AXEBuhu7MzYULsdsWZR6AzS52kJ14uBCmC4UJvdvP6+bsVfd/
Ju64lWjuQUcBaY9Ggi+he8J5+9FOeVdRziwpMKy8+6Lfc+u26xXAnN3JQvFKL6lQ
Q2ezOY59h79hMtEfyLpKjStPkRwLYoRYtDPT12FBFfVCmRzGkVGjawPfF2Bkmssr
9xAwaCnTuJcg7rH6gCVkL63rIwbu8sHiDZZmSqF6HMYJTvm+7GUcBhHOTOsRtSG7
uJIWkyhXhNpV8nbb4jgDb6zcySO7urkhWgcar+NWb8c15aPgcE3f986Xjlk8DSH9
ZpVz2RoQ9aSO0s/4RTlk2j9HX0Ibxb+YW8EYGNP9cJ2AFQLDF7ZWwwwrxnwtcFBR
nWfdjt7AhPo+y6GXmtBRkL7R1JjSk1EnrUOilWQB7Y8nymRXfx2s2Xr0zmFxqwv4
/5kFsxNWU3+TIsSbiW8IJOsDtfHTnmKm3EkL34tWoa5fzpqVFDYzzqn1mgN3QdJG
bu+51DblLrUo44QN/On6RZLzk0h4Bg77Glc3Sex4piyXNz+jzV+6VcMRLmYf/4EO
EJ7wWnxd9LwRy51YIRmS0udlt2Z/TGg1Sx6oA+sso1xkf0kLy6xC154Kh5rb5P4V
ga6hOTtxw1eLcx2T7H6iREKlwe3xaJZXCBUGNDv1HcCeDeF9e0aQQ61D6N+UEBhy
mafUN154Jvr6ezqbehIgAnzLdr2fjMlQROLslKMcQeqpGv4BYlqMqCIph/aLLDuN
mYrEnGrMVuQyTFJNwOu5v/CNSw+d/WSZT2KNOlc2+UIkPlP6oUzNu1/J+goHi4r9
6X5StgQbhVu4ASFLEmTynOKiu9Z6sWqkLuqR7gilXKMompYKKaWC4tMOiw5Viff8
kfKskMCng9gz1HT5arEYuL7+R+nj1t/bqB2yEsYtT203lbSX3W5t2Y7cTAYwab3Z
U3n0ZoNNAUkQicCl2EYXGQpsRy2omZu80BdqABNd389NLOKW3VeGd5kxFx8VpffO
5TgrzhivITpCCRmjBdwOs1UJOoa9p82miae+GxfxkCAJ9gFUf+v6bWIr+W//kKUd
/XTmgvBR8xOs5ofox/uMUW4DPDJu0ke2m2SIWLDRY2hpkNomtGZ/qsgr85hPorGt
ZMmjJO/Fb/L+0iphK7NTgqPq3cvpVYUSXjUZCppSa71wJ8KfnCHfEWtk9txrTMVA
S4lAPOp87z2DsI3g/aiKW6xJcNR6SGaJkxFtPECT0USvJq3JTPIO770WCu/Z/lI7
h7PQcHoFHD9Udrjq74IOf5e3ha7mZvZ3mw6Hf8YmHbQm1q/V2kiLIFioeLn4Sotd
LKK5QyWuWCFw8sFe8qrYqr4qayGfj2/ZVVlalx/PFVnHkm6PXxJdx2Vy3MJfo90r
NQ6x13tTyhGdlK3ULbloSADrqxKR2TbmoAOtc33nfp+WBKHTRgocdwAVyFXSJp5r
CTI9Yim11uk2TYhouNTs99+zgnA6O+u+f9tebWnepS0zByxe/xvFzUFqhOMZBaz5
7IXwmQu0/upAFGCmfnfTz7iDKtrG1b0Jv1vykrxwblXsBl6EVtN8PFIBzRw6tJQT
HjkiJZEqvqtub3oU6jESN441ZN9Y/2eOtscp5sWwbwe9jJ96tz2lNJrfCGIscnnd
OWiUqAdfMdGcajzFK10vLcsvk/sqNGnkHiIiUsWMMGBMbgR/wXdczT+rCqbXk2c+
frUwZDqKKCzZoqnDxMIH2MBJWHEB977UaDVvBHq2sb1CiQmYebrffQq5QVHxnSuY
iXebi3awss3xg5on2VzqmtEZ2u0UOdEmBca35Shz5XQaR/lqYaP4UkSCmuus0jYX
5FbFbkjv3JB+57acr5Tpr/Zeyat0P3YUc5hn+bVrc1vQlQvLz5LV0lQI39LrfNBB
UmdVNl/saBy9wdnSXNVmy3RpBD+mWPzO0jacmr8CnMAi2LC+78eOAE1UzafXnQxn
Urci1FXe6PI7/ND0j6FzggsQcj3oCr2eiEcmWi8KnK0pRHYweudPFRiDgOxNwcld
UuCFQmS7BZJVsoK5wqem85wwetxYGp8hveh8zcjkdMl0/CpbsGKATostlrdS58Kf
+P9lNAg6UtCrmjNuThALqsE/84KM8TBSzajdROzQXGhMEKZ9bo6x1LK5U19tzT88
xnRLvW939munfqiHCp0Ofekqik86LGhACx2+pK4O08N57o2ZO7pdpXc0f1X8rnGH
peuaaK/SVcg3FkaV41Hn4TFs5TPmOFdkkBO0SMSJcZdafWqgGZ48uyLXaXjFTrz6
GFxd0JvQFrAAj2nQmjHwmtJRSE8J5/rdpa+d45R/Ro9BkxiR38Qga01aKPOjYoKU
RAUu6szPw3Nqu9ktW3eLx8lf3X1ilIKxQKsWz7/CZTa+oljdQY7dyGeR0Z2D108Y
zcUbUcjLD6SyfwUyXMILxtcGkqTjYxPkn2XguZIMZOYAbz5aUqXAlxMEZ4v+JD9L
j/g+4BedJCjOjkyboKPTFaXWcgzkmWk5kxhXC5SmbUVm1LKHbtBwYkG5Hl5xG7ew
uwfwDD9lCVPltjwtw+t4yWvQ0gmwc+FJGk7vo5lDrs5d0rxJSM2+ROSrQ8EpVipY
yICrOsMR1Dq/HydMcEM+ZRDO7/VvyYBNhpoUDVGv6YFHTrlvg+yR9UL7oATBx0Ne
elesZFWuHWUPi6aCT1xn+YWrNDjmI6X/FYincBJ7OLSqOF8ix60SwnPSlXfV36my
ba2jm3t05lm39X5HA7AVdxVTGBWGwYD5tKrur/1yVE9JcGmAZ7NzpORi/KkRfLzA
Ei99BApR9R/WNDnQ2PevCwG0enkvLGg6/PN9HSRxEJJS9szJtAakE5HMj088cmM8
EbIvdfixnK9TPlF6dbYMgmIrgorwDKQFb4muFEIaCb8w2//HUypFwOyCyjoAI54x
ZHRtt7FSXFAm4lL/iM4EARwZzBNz4lNNcWuGR1y5UgLfT/kVnax1zbABamjv1hRL
La7cxs8Eq0UrzzlkXsRpU4N/BbqPLYMnFzEU/3zCnUkm83H3ycSLeyHJ3xF9B8RH
pGd+CG9Tx6fsHMPKSUYLuPtRjG+89Ah1ktAjhCQ0/iQpgdVUq2ye6T95Vkvz+fen
R+XIZk/buSNOZSlkkZDYA/685gqp7qLqkuSQcrnTv5gKqLY7HD7pU/0zvV9Fosvm
oNLVpGYsJVe+reRkCbSH3Rukk++7AFu7QNhZpLpaTqz99+fCtLcelssRyZHadbnY
jp3TSg4AERwTiwB4N5bN1KDVxoDYtzofaO6bYjxSDbymtUvHmvED4evE9JP2Cac9
WiBv6wHNeqJXyv8h5TZRRwsESd+ZNgBDeGUcU8B3ZkHDB7o1a9hf89CLLP9bimu2
Y9jGSHQ2emSuqT8QlzLKyzbUPO8Xpe/TMtE/XMGUu9fvoi6/95gTcU2itM4cfbk7
0RpzXRzy6n82qVHAZHwCB28zfyHyROEeYJPYn/lj/XMj62wTAC1KVxAJQepeogMI
qVSqm0ThdRMKahblY5eaRValBIZVycaqTp3HuDB/KkFzDfcRxaWvwNcejd2gJXhW
ukYz2Q6SiGbewSayNmm/1qZRZx5OONkIoaZnF57an62wkHRUsMqz4DbsRGS/Vlzz
jh9RpjUG/0ueNCIeAdT8/l+OIFbpznEXsJAbdQRLphEV+D0DNW5j370ZBEGvVT2t
W2db+CqfXwLrBsrIurphf4435St3qZJ19as7IrUeuqqk69OGyY5NwEQ2MA1C2NMV
Vi3l4Nh9IFzGN5gSfzi2dacWkV44UB4eePLuMmpHvOs2RzMOhKV4mt476nL+1ikf
AfBwmnNzgNNvqzjw6Lkau0VMTxiQVI40kYk6bK+ms84ZdmRj6i/kcR0+TRE0LiCD
8eSXaxnr8RUOJ4BUN8g7SlBIWYd+nc8YNsPHivHfXb6m4n2ZmbsI4bVMcXd5IqzB
IDv5QCd2V4Caa6RGdLAu3pdnCAis3tWZXK92LF6ptSLHbYtSe/LKqaEniuG/7x9C
/l4mydWLD3XacPwaBbZJNLF1HkycWD3WR1viU+z13vw6DFPmuBIz6ZH7lHRKGt1j
5UE9YH81C1ZlAYAbmpqtpVPLGrvVCBeZVvcUztEwo9v2j34EMjo4LDceMLCQPm6i
O8Eg+AQOe6Iyevl+pFTH8aDD7kSfob/QNslY+2cViqrLsnSJRun4/PvdZm/Yp9xW
H76O14R7HkvAWd0eYsk0rb08IM+7wVDXqSBNrbFrpWxYoope1bA7xZMlrOTqCOYo
RHbLU6jsm8px0etcI36iGXyfk2qq5cPZUC0zrVWt20L1KK2R9/jxGiqbZa6R5dLE
oh8aRbZIUWgSFW6CcXTBDfFaLvHsilWmRkcUPWo9U+jkyX0CahVdW2p+SB05cvaA
TEy6fomVkm0leZym6HTPUKtSgVXSKHs1hJHj6ktMgtg4uWrBCo/DtUGRy4RvsiwZ
OY2eQ/D7bra9dCFV+EbW6qgFkTt8oEZpJH1v5zug9WCDOXiEJpqu6kDdAZH8dglC
AhBAC/kei8NsKptioOH1TEXhg+4UUNJXxxvDf6EMAIyW05rrfQu9LypWSAYpfEcW
xAc2EpPl9iatnTnBe33fLHX1h0Dh6RR4XPAovdIzsXpoG4OwfPfMFOMwQ+pB4Ntd
yPHen2paWzGXKdh3VlV5TStUugp5SzpEYEnaBDmRILy2zVZ2tRH94s/psBjfGpkK
qmItq/9U3mbDu2FNgEjWtF5UaqCXY3azLKDaFVTcF1GseRTOuH2y8KxhnHb2R3mG
on2KG0wv5ILZjln3acoSfV5uik3X2Wi/HvunB2H4SrabeV7UH+hP3em1lE2F7bxA
P2y+xKZ67FDcy9yKAz7snKQEex2IOSEPpAolFhqBUzz9GBwj3OgY9dMBbbQW4ji8
OMoMeLH0rTZe3elz0T779ZY9xR/eAWyRyJaJLDY7j68fNRPaEE+l2kXIvg34mtK+
WFFI7XaGAco/x9fvPXoDUBHxZlMJ+d3Qu3PRkVLJ8W/QYQ8suid0SyHGBV0zwE8R
lne08mKtj/5s+6AKPgPdNX0+goouBdkFWnpg85JqpSRsrV5zNc3CSaALsfVQSSTa
vaUmigtbgWrbFpLlQYRshGzSFEeLNOOZyTOtVcGcXOHf9VrkPOBEarvE7fLD/3FN
5KdfJ4WyXLEQunGy8B9xtk03TeQAX03syGXCzFQYPtS3XQ1SCiI+t3tTxoWA8qGM
zTSvC5aIpBRHPeV06cY+Eg8hK+XEFNny+iMQc6DyEFnOCEl8TkV01THcylAkbI4L
dSjRuYx3eeW/eWK0xbxQXV4W27toY4ZPvpGNipD+XdPfs5yXEH9tTzfVrck1o7AO
KmVIQDrvyayJ/d67b5xEsIPNYqUfKCxfzEe+9oyQG+3ndPcOLIHCFKvG/lKxm3wM
y1sFehmqZjN65ovO6wVNAE6E039p7ZbDGSTijItzAdLjKaKJsDxfjK/LL9MAtUf6
UtHLDs6BAB/n5+L4C2bGC2HTQpIBthrYGwr8z62TsqeW4GLcU0Ql8jUTHnqUuUaZ
e7X3WfjSMMoH1l9s39+FS8a5XGBj486tyclno2cNFBuK2HzmyhPWSR+d3TGBolBa
LdRLLktn0s4N0EsGVATQ+7vVfWvn+n8zKeMWkyGH0IzR2R2BSQjnAfb09AYTEcis
UXc2snfgPf9jbwCl9DxC6maGoPJ2V9HeSagX/ERbgsVOK9bJkzGGTgsfl4jHGLsN
s3objq1jHk+Mxo+gP8ilLkvSU0KJsqB2Ow6O7zzU/oVeak9lUijGY6JEKnbL6gXE
iXpVRheFTJ6WYyGz0KhM27vH8SKD5iuchjOYfxDrl47TMWFNzk2kzIZQbEOcgzCO
2MxqSXDP4Dbw1R1+2gUeXDOjAM/2lbnPjOMlHsE7XLe+os37QCpf8310KxCX+W9e
UPApomR20mwPBC81GxSa0rREHUEJvOwZIx5bibwG4c5KK0HuxEjmIv+NLbmAn5we
ZGAm34lhz347KcF4+sSEhLOAAx6GsYvf8PjBVf6v8BF6tLOzTwsVuYm2ioGl7qw8
DMTdcLTAqUGX/sECgjq4LWICyyooL2+ctC1CTXmnMY9q9JvNgSrgnxaK0/u0S5cT
IXC3LZZMeFBTKlelSrJeRVY0fDDXeE6cuP+hVV9FYbJDmukCOCwiPyaalAs/PbwF
/fgSaQ1pTxaMVYv/jesD+GNvV2yNeiO8TrUcxg7BUEHJnZMzoVf/1dIaIx0zg6lE
zruPEJ3t2ICeoMupGylVtx/ycn6g8xZffTT5JwkOdDuV4v2EBF7NSmRnBUKqai8v
+6b2xp+JkpDdLfaZUDbZF8CUBhaE7wqRzyW9UBnvupVVtuBCOozoJVlYu1NueA1e
jqS8lwbz1shGMNmIv0+7g/4tZ25IRPvm/4gb4BzdoCyRqP5q79sLWu1Ab0EekiID
/grtm/RlCoOmt9AJf5JB31imLuXffb+EjlpOsMi8bTaq+CyNw+FhlraBloFLSRxA
pLlJQipBHKVP6nfi5upYDPfGQNtUMtfK3GxarF/qOc1/1k+2jjIig60h9y4lfKuW
t4yh3zNwAWpIyHy2/Ls8ORKSlqQHeGKY+/cwzqfAeSbUWP5aDJbxjric+EC5QNXj
4oxnDrOpJr9GqKEVohSIRdZUJEQmDZC2SqIE3Bd+W9FIZ0FSEyevsXjQGqKTGIuf
l4QuK4lgDE5xT6E1883btbv5n8jtxbB2lLN0XxUY4Vfyj4wbMjic/qRzWGbR7Q5w
oyiqXKoZGoFuXeRsMvxk/aaXguvUPcKvMeBM3KuoLBuGICLSJ6/cXGLC5I+eBYuU
OTnN3DnQdtF1tTpxu+BDIDnUJdUev0cr712fiNX12s2/o7xA/hlkIIWfLkygg2KO
KelGkI82tQdJ5bY0p2GebquDN4jWD6zGu5foqdgriUif1Ruzks1UkKFr7LpVJoYm
TNA69WacYwVCqHS8+dHDh1jNpokHk0aFAOShqZVdi6g49wncKgNH2GR03jgr9fz/
MH+4UeluyVwCxU0QNRk1KYV79cY3o9k+7Kx7/t8DW5uI5Id0iZzSY3ZSKaxZXUVp
5irt6rL49AhkWI68EBBvRhyWMiT3HGgHv6of02EoyA+Xgvg8USQ+p4p+AHL8TdjB
p5od7jP8Nxp6Kj8myC+raUIQwxX/rIrXe9Pn3DU8AXNpkgCeyh6Fwr+ub97I0vVO
MjBo2oCBLU/2dqeEMTcioesCfmFk2IwHBHVYrAL7QMMXnqfwDRkf86K2qiYppeLf
w+UZmFTU5VzCOWr9GsGG+knI+YKyeCiUKqfe8LhPShUdGwYl+GNnnGzKcZWMht5d
5TNtz2tGGim/lTSL2BKCUboTG051E4Q8rZJQlOiyWchmQ9yd3fLS2VBCtrQkISdW
FpUA4GHq6Q5pT7rQx5QQ3UtvZ/VvP/25ST/Kexo+SgSirLiMEYx/ZNtFTbb7/AHY
RrFyeJJAAAh/zTRG4N+cJMwAbCe8qYQeMxM69ELHAL5DE7JSro5x/mzlZntAtbZX
QLucVpUUqU8UX3x2zD9xhmOxWUrA7Pqc5Qb2rG5He7j9UoWLBTIsRAQtqRrcLcYf
1Wp8qBt2nESvWHld3Lh8JUgF7N95kHJC7Cy+YS2DdyZ5EUJ7x/dtDA9js5a8tTRO
BTgj0wRyGD0CrZBsNSUYY8FpEQLDFI4deQV5EUb8bIn1tZtGB4LrcXrKOKQ3pAKn
XoBEdMWvxc+dAVDK4mCoblNVCgjm83hxCHvjHKRzo9k2oXEa6XhMQRxkLK7R8Yxl
XLCpCl7VzbHz0AgmxmeY6MUVQ49U602B9OjBkT5S94WA50dzSeKIfdJVSzbbJu00
LiIslg546XVW8K4f9mMKRB4+/sjNkMzm4aTWNdIbUsT1mx4Gb09eGZ9kd6Hozydq
CjhWZLdYeBQwdzO6JqiXh6x8AhaE1c2k0z4dzz6vbJdK7+hUjOMHHDJ5jWtFs2j/
o/PBZGPNgppjoqM187HtlKm4mYEf7OE8XHGMPKUYuGFgeistGJdwzn+Nffg10/B7
2DtZoCZC3R+YQGhmKpwqtzisKb+pTemDhZUkptMETsCSjwQ71VWLIh1Jk9TmJo6P
HIIR45t4iTGYleprYWjD39kFubEZv1q4gafPUXNLF49ygir1y/PSIMPuAL2Zb0E5
ZGhUpAzxZgJ87oFSk/FbHjIBAz8PmpsL3mZINJ2aidApnNgjjCG44b4N2xlyXUWA
0SrIQsv60/HUBlM5IzXR1uz1Bz4GToQiJmO6hqN0QWuPsCaakJKTfUbnXTZzXfSs
1VUXonxYqyPQmIEMV89ubEiOnmwaiY+KsvbyPtCH64S3NpEveGG9msvXZp3Aiyxi
X82MXl4MsqM9OPpG1mEfLmIfdQdwsLodNkCtFx5YHd7YproXLk3wEGC1ncwl9uNx
B4jujA0Op5XJl7bUuSrazKX3MOCcNE+rAzcWxE73wUT3zi1NVHIHx5y2CPy5c3/y
OXruXBkEV9A+gfoYdjgDSIYFh/4nE8YcF3VzuJKuINTJFyQmOCF+xtqNHYvFuSIQ
u1QL85BszIhCndIOuWbhwao4YkG4S0vhEmafg29z7+dGh4XIoftAOGPjsga5ApgJ
P26irkNn933iT8NujbwVavqP6/3z5lIc8Wv0fwgxjZdDZw5hcyXj2ZVhyXW5R1R0
tXa/bLxgm5fVN494aW50/F4YLR+sCIyyM8HMfrSZifHhX+uJin3y3MP15cNtLz/X
Mw2Zua+LMu+Ss/zUcRyxVdwiqyS7TjsybB/h9P4JQX0KjhF0XHVNiXHYXBX9X64W
ZAMtYqw08M3BrNUHkk8qL0XvvoK/UAspIbl/PlmvZQoYggT75MznP2WOe+rQBYNI
J0A5Lx3u1t8ey+YTTcX8ilm9R0ScrgKKEqLDysruxw0ACnJw2T4qvwUgU/3RRk2I
dQ96rWMeMdMUEBNjQ+tE4Vdq0dWOdSJENy+PXC8TBr70q8qVaP5Rg/LxCc//e3s0
jE1+XUzMFS5FxgEffpy36y5zNS5tPmudHiF5KPhGysz7k2sKFenJnO3nFoW2arYc
JBrk8dgHEQguTJDXNA398+2yYjmwt7Xvshm1d7E1bzNMS07OGUNjjhJyJF5CPb4w
II3XkVkrqJSSUCbenjmaNMX7KuwHN1sir8XLfYu3cQCYLTXfHZgYpzdpw7ZzsxDg
gnjhsmibdx3tYmYXWoqXOdHedYc7LjUBSD+rmD3Wu7GAoyIxACnRmZXylJzgHE9Q
zJ7CRbeVXR/j1Dslq4eFpNi7L+zvRYgWa6KzZKVSUuDV6aNZBIruVPIIlNxL0/LC
X/Jcu1JOzfNt0yYUoWl5MWQMLOLA36j+BXqp2A7woF8sGBx/21bMNjGujXKcOV1k
Fqt1hmjCuaBxrD7mX4Kuxy98vWtcttF2BGAi3QXXneS5A3YDT/SWj4O+EP0VoG2C
2m1SyXeNhSb+VTe0wVe56SYeH4LsBO34nYkmiGxM8/rNSHeZP27clDOL5Cmskr9v
vIgQk/OETVX/T9s407geP+/5SQO23k97f5YYWOOE5lCnckf9u8ZtuiYqhSZPP3N+
NgP7N2BCuuACAXM0HdtZi4Uv4KYmRuN8zlZuktVO+UeLrx4q+9R97fDbC5rVXmRk
aLFLH4rCUanQHImIKCQwH70wiFl9SvpWm76YYcz4wMGqFVDx93B01n2ZzJ/MQKpY
apm2uL0ZwI0hJxp/9gcsayH3ZOhXbxQAxc1KCcOgZK8N63RBQ3cBQs+4hISLzUew
tfLad+Wn7Rq92l1BG5pzmXR8mfwC5ef8oblgBqj5O2eSI3a8dCFs7SEyYM4M1WaM
KK/CJmV5u9DfysWTGb9NzbB0iMXi2sMSsmlpCBxAFWapwUa4RVrNri/drkSWGYgX
/19C54OtDQnnMCUG+yHeC1RnHZY59IZuEqU5a8ZxxiIpH8L+S1JfBPc/keLAytdj
69WJK/hML//YY3/9rnWQNHRVNVasAOQUIqyu829K38gOtC/CrsX57Dq7cXFaDPn+
EdOZWShqZctw0x2MK49scEA3lPzytd35xkL3SSwnB4oOJpDPvS4kErkvY2lNDUhN
/7gaHA7JIUe8jqEQfFDA86CrOHASRsCRPFfSlm0RWixtDsMinVwRRmhaglXtshTp
LuhhlwkzYSJtZmytqAfbfKm5goFrg+3uZmq1MSWSACtnXuMjvLUlfqtWKgh7DaRg
7uYe6ji4HEQbdg/rVNEj2RPzWOuIj8M7AROj4mxMh0fXQpXVlyOI82L1BJke0+NP
LsvuGGcs1eBSNcbBqMDcWsBgc4sQYymoRp35qMQS8rQyE0hR+dKKRJNfHa8z4XwJ
Z0qLLMnCISajbRV7tjxluo0+y3v27s+LoJZEOQKHHYH5qCVHoCmp2lMuci4Xi/Om
StXunjdRrNglxaxpG3Z43/EFFoczN4fW8+RNXJP8TnBj1pptVIJXTrdedD+nZXv2
s3s0LoDpa7GrT99WyGrCy03JcG4khuZxYZydEHHpPqTrnS4oSjcl/lV/gOp6pXew
FnxplSr55FAfMtiyffqFCfWTF5q3klhkpPNkw0+A3+qHXvvPlA3s820Mh3F8HncZ
FaMXx8U1b956yYDYDpM2uHRqPKJWafbIDbv0D/TbtMlBjlhf/PcxRo3rEGUGyNjc
JkY/1tr6DNwX93JP5Cg3gmgVwwvgBLNR74R2VbxY+Yeq3AoXu0FJlSZsxLC9e3Lx
bU9a60WjRUy3X+JyihBaSLdMxz0b5lQ3UnRW4/AyTEs5wNSHsRSD8zCALB17dYbF
dVJEmDfDNiS7HNW2hcEvTJ4kptn9KSQcm1blXWufdGdzZsrFo+7dBnWq5BPukSZp
x3MfeTOJE4ez3G2NeQIl/R37nY0fCZepbgA+lTOAivsBC32hY25TNVE51UJ+Zd4d
E+/XeFDlI+USgR0LDgBX3NmtCoglH0nuoQMrCoB7DmAAA1VpV2YJ8VkDFRXPKYbg
AQV57F7ZLOZH/mc3WRQ18cZXy6vFpvcHCxYyVSuHhM7Wy5IO45h2i62eN0UVxHt1
o7RADlxWP9a2/Ox1ozg4sNXIzb9kRHjQ24cGk42kes9mf0xwQtOfEYlSoRCF7V3Z
PBw1gV7/f2T0SEDwGIuXLNqBH5Ufr8++KXDYBI5EOTFM2YBXzt9B23WK91XBZ19B
UbskJ3INlvac1PyTAWExGYKQUaNrriWkwhT7RRzAcuCLXqC0UocbJKdok6lJX/sq
x/XpoVk3hZeC4GijATW4sJ8DVCpxuo3s2jYMT3/AytOz6QvPE359aj2Ry2X0HNQl
95Qyv2fgJfCAdk5FzeJMWOS+R2APf55iIG0hS6tfLaIE+z2p9FsxFOh5XruHx/bX
eQxoeN9w5obTRUu6RNZSDjPxf/nycw+qmxryX5Ga+K0EvsAgi5vLh6woHyYUUisl
21JHMoeeGvlfJ4pBYqnrEMNZDTgmWd228dV47lS32CH/M0JFhS1dutYYQ4UA+Ueb
3dufrxTuGhHJOHcWiycjc0rubHeX6l+vXTWVAWxh8F7J5ZilmU24VFLhNbed4Smy
pQmYbGQ6uMiddyEF6Nr156IoU4vfzYBc0VOV/4gEJXPJhY41ofrhvu5rtj16jQrK
JJQudGioIA6L3BGz4JOsx+HAgRoluCr4M9hBW3RMB0vB+QVucdTCT5Z9ibbiv3We
NXscwaMSRBb6MsEgtcnpzyTyvDyeTUn9KEux6PwTGjYdmhoZVkGw6Ngow7r6PMZU
oFtMy4hIcbN0dT97689XF08IRnAcpCFqSubXge610J3cHyAkE5SYQ4pcsurvRMgp
0u2m9xU29utlFr7jvubCL5FQ4sA9V8N22j4VTd1c3a2Io1SiQwkz6pgaWzkKx0w+
WXsudhFa9+YixDdoU/n0v8JT+zGbvhzoNy7k1TQUCkFju7GW8/HxOCh5uqt7rnZo
yHFZPjhn2jLOf/Od/vT9PiOsXLrtcaJHv8sog0xIMGohUQlf5LdRQLQqDdKbIyIv
IZzUgSX0N/9poQrjE5JGXuG5BeNoHw/CwkY/zHXgrwp7nTaODsU8N7iyq+QZJxjz
mjelmdsxunTG9XoQAJ/ol9LdqEB0EJ9I1S+uFt2GGSN2O8rvDqcJAxWVze26PShi
Js9va5gld3k/akuF/QNp8r3bM1KKSoQhVSCuBh8OvkbdTgsl4uT6OAbCN9gmnaRN
dHcpMVPwGtoRYLRzt7Fh+E/8dE2fSgjacDKqK8DTojalaQHVLhL9pGiK9qy/rnJu
BGAxyA138fW9vzuDhZi4A4NTuH9gUCZy7jiwc9Vo6fFxeOjuF8mD1vqbGpjG76pm
Qi7x/hzo6qEfHIV3SGYoOSKmzgpN2wqogL9DySYOy+lLhgm95cVXEqcP/JfLHCuH
0gtb3j/XQZbkQalPLTUPNEicnO+DdQy7vicnhZiOJIJfuOfED2irrNkj7jZVAYBr
MJB0FnWjtXTuJ6nvVS8ouFE7DBHm1B2PzzBW0m1oDUIC9hKsCy7MqSRu/XnaXxAy
onizKYCgga/YHNAjHfwhxpnqI3q9MuTHgmaz5iQMyU8n3d7MvGsH63G5dzU614Wj
3HxN8yIZdV1HLGtAW6Wk7y/S34FqjkDBhtxlJRRa2fk0Xmt5Tckdy30O4VlkfzGu
P83WY1fQ/UmrE9koFLSdMNqBFDZx/If1dc13JuzzftIzKfKxF86cINiVGf2W3Gap
DJaVSvx42sckPltS6JIuhO6j/BzqrnxDTdFDIBep+u4hMwuwG0wDuSA/3WzPv0jQ
17Fa3UlaxjdGQHtFdC94m7ymREFRFoC5gFxKj5G37a+mrxXWQ8pYzkxQJbTzdj4m
bwgIwwBMGS3mqPD1p32hnWbQt3mGWNVAXEtQdMGUMpBi6QXxBxPtyDlFlhbUeGUf
/Q1bYm5to+2b2VETLWgKYsAXANOG3ZsEPRBfUYxuUqKhzP50zw/vEJVmNGIbrOgK
9KmbTft527ev7SmH6w9wrnz4yckYp1ZCNanx3r9CM1GtRqpAb3wv/9mVes5PZ/3T
TMtthqxoll1gET6ehGMox0H9uumQJy6hBfnbc7JzW8VBqtDPnt3dCHzMxSo1zc6j
G/yCtt7wb1di/7UC1NKQBc+B6fu5se/MQLBhuZzQAxxEaxaAnlcVud5/s3jHkenk
3lhddJJwhLKvHONkcYlkO0pLCAfT8OFHc9TiOjty+fx1CqYfIHbogZUv8cw80a7f
LEWowMoRp/OaPdFMxf1yFaf2+s8mul6CJ0iqSH6h2/Z4fRM3x8tNpQgmEIazHE0E
87iWa83WIaxD8l8ZIN3070/fvJiZ5IbBtoGHHxSNxLAoyA/GN86tVxsM+yaszZWU
vUsru39dJoTuAAro58VOQAyhIcrT3Eqb6S+/kX1kOsDz7pTtAG1fX+AtfzoZozYc
GY10BbeZoE7LJplmtPiamdhcUZHbqxr6uBquCaVa826qAGEc09+F4FOmJL6YLFIl
NdqXy1GJ+lfYmmvz/wejRJ/Rr7hnkYNyw4M5YMbrNpKkwekabBvhirvEwCYKrXq+
xq6bJcKCkTWW7YI/4n1cr5z86qKG2qP+9sqj9Gq/WjwXZSOwiYRW2h6VbSyqEFCu
oJqLZ6HBU6TqaCxWEwvLu0bdaeAouEGfNQy1V8vvPBacJAAiXYMKYxsw3taPEEBC
tfSKC1KTKdB78eukx3Np6kxUQMTlDF8vzNq4xIWJG9ZN0xI4U0eaUsLs1O1SczXt
HVXnklKyHFXiiNi8kYR0MgNcnKmi2llFuj2knfikd+kYOHQOTvfaAa/6pQr3Oor0
8Fxdju8HYSVXkpbq/BbILEDlX2dcNL/2y5Z6fxSzrHmmnXKMiRQ8Ujo8t4MK1++W
dgwEEz1vEbk346Y+Nrk1IH7OEdH76QsnTeiu7QQAvm3awLsz//4C5YogCu2z82Ma
Ig97LBq+jXlZjDgjfzAkCFV4JWCDvBxBt2lkeWOTxoj0GIoYHIgCK/m8XClwC4WH
kpUfFPBgwDNyjVTxg5HsmJsQCBtWTi27cwmyPmfeVGrvQJf+cZH5d/9s+hxzH6Va
DLx/p6HCtRngxPPBOuwgpd37nifoB1lc9GYfLFNVHgHp4aI69heXmccUvz3zgUQf
xqaDR4ku1jaN42Hs4bXDFr5ic0/e7iohyndQgH236YlbvshiWAdwDUvsoqGGYWYd
IjVRbOVsc2lTYpPZihJwYJlWmQz27wSZ1hW/k+f6W5Z95um1EVrtUmZXZBMylWfN
h+iXIH1TBp0WhonqCCRUQfNB2aY4U4n+AS6iXwJoYLF/ijZJWBhpLm1OQ9iF6kuG
h2fqigH5FzqJE5mXe+EwDV1thsNWl0uBG6nbEYbaW+2yUNE2SJPbCv0FYFdrStH7
W7bzFY36T4pfHISCqdGcpTBYR0Pl2o08YzwHlqd5gLhqQRVczhbYAt8WXM64WLT4
72CKQcfxB9x5b9/VduatpEfnBDOm1KUSaNGu7o+NlIHupSw/8afJqLp1qGbtBJkM
pbdGEbXXQRvgVVp+QsDwulQ6bjoqI4WksmdI0afGgUEUG1rRix8txJgMVJgUeHO5
d9KyBfod4DZzy1/2WqPYpbZ2h1buj0HjQEbZ2A/uHjTfR763HbfUExhNzL25mUk0
JxUassFYzdSKZDE4wizZCJsIUN+MoJfnfXXeB3Vu7gH70Pon80Xf5A64x+e3vSJr
RWV8gYTqYA/pwbUSPcWnObY6Th47AMWLEPxL1SrlmvjUaYApEqqRlCsnX0J+2eFB
201tfG67vLX9kirc/AuwuWiKJtxhkMvVYIenDWxZWFPqbTi+a/qW2xSSPKxLZbTM
bZUB8ALG6DzzbCY1L/MW2fgz1BldVO79DJvXA5dlarA3bxiIq8rmy4/o7+aAH9+B
EOlNjp+nXby6M7Jx4yCTu3fLOroCkDix9+Mq5f3MsqtE2c2UOBS9CNh4a7Nj5dPZ
It7xwvq2nnzyPMClg7Xnx+XCT8I/OTT3SDVxZb8o8Qs7B1nh28GEhdnMGrOYIKOI
8keaDeKmqIqAmyaidWUmIrc2GLCCFssbmzp5dHPSUbKT/Og7bJqOShaKxk0ECCMk
buaq92MBT39kNzAwB3+IELNvbeIojaYKXi4Vt16Wq8GUR0SG1WZzbdMVrrrmBkLW
twoti7puTYmdb9YQ2doFpALnSVJ4cK+t4aWOocfetCuO1GbxyMGslWDlOsdFpYgw
M46XQGzby/GIYFbLSYOEeG+YkAYts5+Fvambsi4c0QYRtuOOufdgmUXYcWF3VM04
TQfJAirIxyBK+aqwG7t3GjcRh6B8g52iBxzO7DD2nzLT+cyaLHpWDPW75GdjAeDb
zx+4qYEIbdy55360dYNapsLBXsnK59b94oYOCVw8n4Cbcb1K33wIC9zDoOE4+q6W
DJAZKzUkZDTbwpl1RdJVlajZkbnIjqUruC6kyX2l0mLMuS6aPdr5ZfYYKI9z47Et
J6HVUbVf8NXRjRrPS8+/eE6YFO4vqZgbpm2Bgh1otrGUC8kPasdiiHUI6f+T24Ps
ts54T0YZroW0cVuJXqewosV0fzbd2JKmfJBf2O3TwHSYgNbc5Te5vx8LiREH+otN
BX04EEBLnAXVXVvfBsz6xEDZvr/it5x/Bw6qQfThDT3neWpa/GUkESsu3DtRndip
Tz+GkrLOq7WxFdby0khjX+rcyQ5BO2WzFE/TPKgqleLvpQjG5kZP3knSiYPgZVwJ
eRZ1bji6L0j3mD8Q7VCEjFnJ/0Z1V4mOE3gqwtbl1OqBHXGU65/8hCuEJaRIguW3
lUXSt0J5a02+GvoKg9O6nbGhl8x7soIXQgAzhcqneEOtNl5ebj3r0W9T2lJ0UvgE
HTA49aejq7K1YAaKP4/5srXaqXd9zCxVPudOZ82T9hDt5nTBnoL2/3EPTfDAYVr5
HxwBWnAWjI2czOnUWSz1LQz05yOLqeHNf3kj/ypDzjdgpNevfoA40MOstfdDYaNe
mhC+GKXIo0j57fsFEkRbZJmuOlvzyzaTu70IoYXXUiWt5LqQJhvtBP2NBKtVde3y
Mfl6bLsD8hUZIkpmn+3hGBnfZFcGnmoW+qDIEQi3TgEDEN/9f5ETCZPfjVT89ImA
wrhIJXHryYFUrPif52uKjFwdNAgacmxiD2ZIv27p/LgTCECrXycQphkVqveuHypB
LHImp4F7xKxkJfTPvjsBofjxAbRrQXK5MMrxYaQRWadIXEvq6lyI4nJeHo0JaCzh
F5TWeJw2CerYvu4z6cgnvijzXbWTy1OMbPpRB8SVFydOFl3UNUaAsA1WtFX8SEoK
ACyoFYyQXen8xrIkA8LsRoYhEGT9RN8wwvw6WoqGgudY1d1/chy+eY2lUdDnsc25
3lk3kWiQw+UZPUi6ST1xnruxLouSvSjE+brMa0+vYC4s13wsy2LZbsxnsBtCb6dC
K0mQheDrpEYLiULV5Yn2/ur03AFw7sjq3T1g6gO5UIcFet39fSEWeLnG59h9tVCO
1nQvYkcBDqDireuRcVomI9KJnoJSRbZ2zrR5MtJ/JwR0NVu46ov/k+eD8PmukVIT
dWruhN92mLexfm2QkTcaxIcwFdxdgQaPySYZfffnuJglRoU7gQ5auCkWJl9fLT/D
7whdqbQJTvS89l+ArbjFehaoG2zOEaw/XHOXE5Qbn7/7/cCainDbLHYdEicB20z8
RashXRasN/RTAF+vbqfDN4e/SaAP8v8NQcIRmq/yNRzu3TP5XPHnxIgZV6uBVTgX
K0L2kMBQdix7Ln8T1uMahbzHc8TarJ5QZtSg92RlgbgZmYpPB8XnX6r00NxiHJKo
atGgKSGnluzc2/n864y8fskz5sB0QhY8v5hWbe5NV0V05/Z/fCKMRjDP/KQSarvy
SQGkDi+D7dDSTtvEsrLRRCsc5yaH6AfvwOrGHXboTOpP/n/sPHD4FQG3naiKSDUN
BF0Um0CBQr3g/gnIKjfdBzVvZ1hZE8xcreopUR/mfr8uJT5v6TkaDq/dklqvM6sb
9gQnBTjZXw9uKhCjXvgTsGecxfvSsEjVdCqWgIO3AbPvemGn+OKBeGferW7c83Ea
PZMZfrORYIGN4La5kc/7vUxnGvP9Vq70WMmF6ulS1/b+4ctK0QKl+sRW54sGgzeA
jl4nh2zpTyz/yW7AQNbsKYSGBK4ktuRymigg/T4TLrc/KLD3J+RSi53U3TNRCAlF
0VntAdsUY3Gbn6lsYHyzTXL84NJeZtAoAZIRPiSAQqg+OHAkldyipz/HIqnnR8ca
YsTVRYbYgzH0o0iL8TChd6+slz5NjChwOJab0DcvfamE/mVqtueTnZKYHf0aa5Mn
JWhs+mh0LnTEESp1Qv93DSQzXySfAPmHSNm7ln4jDF6S0lZewKa2FHU8cmLDk1OR
dWlzWWu4+AaA7UOOpINulLLcTvBBRvfoMVEdCrCYEMctbd45JPEibf7EEAhL8OXZ
YFfk2/7+F5S7yRo4jrUfpeNeAvrnWGR38t//vqcGTdyaCkMMcRjnr14MhvvARueH
OtJsCoirAbxc4bcPsoBl6HcprXH7LU64IglB3f/jXlDOtzpMpldyoFx4QK0smBL6
ipXJ3b+S+o8yYjjtm9d4YZBgKUhfXsMcbTGfCxc1TFCCwjcM7NqNHRh5DagjtUuX
m5RSU2YXG4iKKHEUp5qStFDMRhG2Dm64LWxTYOiQGv+V5d/RBOTYuGciiB3Pb8bC
cA1I/A0N/hUJCMJ0Svl9XKBgf+KvzV7TmSJZwWrP/rrp8KFvlnMMVYD4HofUChQ0
e+CPyQUbQvcErHTe6mn0eCFk8tvo2nowLramD47S1HncaTbP+H/r0gtpZVmwv/j8
wNrQgESoCXNBeQL2sD90hRl4nB9LSBC15tY7Xoltc8adXdM30z7AnqJzdFnhc3Vo
qndjWUnJszfshRHq/TtAJnW4v66mR95xO3+Wuln+AW97N+XKY044qbVZfLc1QEgj
hyR6tcaemZIst75t9rLxhfZxaQ6jV/P/3VwYvpvnKMchycgZgRAZRc/gou3BJCDs
pqFXSMGeXEa3MQ+MJHW0Jc1hUt+2cxVTGbIOvCwZcS3snspSixDxddgAAZWxnwmc
AugowM8htKfoO92yFQSoq375TherxK6wR7if3c7jp/69/KiGgwQVSsUT6dHE3MH6
upZEXXSAah4T9H9AEp82TbH1shwPJP5H27ce0Q0r09xNOp5M0K6v/j+Z2LgZ4HZY
5CpcrJRSw+SFYzvq2toaUpnPWs/5IRPYgVltNfz3HrTXqJqTCjnM1LeoiEBmybIu
J8wmU2O8f+iu/boNxzCAedlrYkbmUKu4gPYrkGCJAz0xAEdavolmPmrUyN6IDfxE
XKdg2fvjrZiwj0h2wlbYqJe0WLqUrLZ5SqJWvLmx061ol2RVg1N4TXbdF6/XjLGV
km7xyua7Ad86c7QpRKk9aWxv3hNUouNdJgzqt8hRxn7tcjqMeuZKIUIHIzJgmPNo
EBhTo/um841CrOk9PzVLFaACpj9BFN0m7GiX2jv/ecf7WcRGYe1waxRYZLDgIwY0
AoGHl7RZfFMm8JJ1J4Pwyvhmzw76T1d0PrSGZntpmXzYlj2oQRNz5/HDBoQOokIQ
QThGDjfOylK1R2L1gyD7xpBTUySW/lmeA62FoXUK5m1ch+SettQ0fYsyjNDHDk2Q
643N+27dN61SZrFL6H0kILD+aSBw9NXTX6x67HEk9CFwkTxdnvjk+F6vO15Ox6B8
I+GxBWlYYcWUpaTmC26X//J74+6BvQL0zoqNfbphoR4fSNIKOlwzVlolwyMd1jmu
kRC262YOCjM2BTIdt4zu4LVQvbRwvQlASJmBx1cBdGq5/D6fuH61fcDvndTu56kf
c6ssY6TDYThpqAQ2RzR7sZ2D+EaqTZ7MaWRaJKsL40iTi6zV4JBnXi4ysHiYi2pe
EtHh4TDDHr2CW13HERKcO6C+qijFnVOZiK9Zq7It7U3lMS0eSCoeJyj3BkjbRyOp
AyBIcpqkVAj9E0BJkO2TGBCT5qlOtttcgxKSK5ev/FoR9i67FDWMnavTiVpkdvOc
O4N7kB9at7n+SxWTnFJTP7+gKCB5h3PKt0Hv2KZ0hdjSTp6yU6BYFCue8TQxY7Cj
bxSoFbubr3s3C0kZsRubHz1ZavaGajgUeizlIxr1wRcTWSox54IMt6oqzvf76lUv
/HrjICLCro6X4sRnW/e3ipquWZ4kJPx1VkMvbkCJiqdg8qszNhjQgrfpOzBVs+Hc
I7oZmUvT04B7VeV2t5ZT2Tf0ZfoTOB/+GxJysVC7uSaZyEkdAXQwlaOECJ1m65j1
XKAXCOiSSuuLdDv39gLCa9xHPY9oCl6SIz0Y7f4/CxarpfPq7OhEhw+6VoVGZpHd
0jIZyFOLAMd7t9Wih2OMz1N44mklNfQL5i3xTN8j9soWDfj8bFuaQG1GyL7YZS0q
WeaucfhN1wPI3cmsqTSKB06birmp/lyedKvvjthAqHD8oP0yFA5y6VJP9wXbO0D0
p+WOMiUoxgGE8EumccyKTGBwbyYtT4K52g52ZLnYGT2R3Oo5a3knmr9QWi387kt9
AN3FA2o2wlWC9Ex299pNxAKRRKxdVCJTa1RAgGW7pcXOg6dEJO1BwhPmRayiwn+o
F9lP5FnvBGj+6Z6/HPMNY3Ws+0FKGbV4dA2waWwbCrc4sbdDdPP8P/RwGbWmuq/F
fa2CWPjykNAsl8e0tsZc58BJjzwIwyo6kUc6A+K3RuF/oz7JhAIcILCAfOTsuqgK
3xWseialOacF4O6gXCc5ezCjKAe+6aV2uT5zh2ixNM24o6iM3D3Nx3RtTO4OW4Gz
ypiF0C/632S0Tmpo4RRpD2q5OUxY0Hk9w9AeSDNqiFa3EhknCWafvvjUadNnEr+Y
M1/cWUb6y+VtJYxlxE9BpFr9wPOnVrvIFh0mnKs/FaATB9vWA7IpEmZUyEHOFzba
bGwn9f7Wkp//cHVNmg/aLk3+W+7f1nR8gF8p3UB01FySHOir+/QuQZyV/36BHKY8
JJUKOvNgY6ikne94HY+iNr5vM0ukNk+01Yed2AjCAZw1sxzjCmYJYxySqn7po+VP
07AeP86ToXteMvgIPoV99a2+CpRMTJOChS9cdkxJCRx51vKr+fDFK+Zfszd8/F0c
xfEIq6s7mcoh8nD8UeixOIvG145ecu0cEFBBGyKUtWXXtQ4R/KfCEv5R7ekGkg14
VO9jGF9PY1LblNY5BfAprkfIPk/lygkl8lAxaK5K66t0YtYbDQE+WMg2TmKbZUGu
zTnqVDnP5CX1mmqrv3un7VEzBMy5jz85CxYrGZ3livYuFkgouRTHSVURuWlTg0j/
a59e9OaNR4EdmFHFxOdA5ncsqXY0BBZRCkLtD0ybN03h31aBNLAWqesjct9CPxCO
hYAfCfYzFvQIBY2susSRtxgPbSGFr068O98wX80ccifz+iKU0//VfAHlVPzvT42S
jj4KYNWbRzwIDAqlJwtHoY6xqpFTgFh0Q4FJa0kw6mKxPxGKLc5SbEGl6XfuZNtt
T2hvDIO2vi3KJyzaEJ5Nn+UeESuHETF2syxIu4y9ny1nMw32InE3loqJiBoGLuUy
aXtZ29260LPmLLTXH6Hy94xlQvj0cMd3xwwrQav7kIfMEO9+8tEoQ14SxW11J0E4
rYIpl6sfUkpEgC8GMDqOXUZ1kATrX2xdG51CTerh6+jbF2UmwzkkeRLM2xiIYrZB
w0FvtxJe5rs9BdHboyUrxGCig6cTqF0mt99OXt5ESfzLlGWRdBlRm5oQDK0N9XIr
r1yKPcHBDuuxtKU2zYGbMLeQc4vfLNCQSVLfItFUkstyXOM4rCs+gQhTpbYjyrPU
gsQmImMvr6zQFDHBREAaqz+glJY0Y2YaPUOb95xzNcSaCK29Py6jtexIr+IH5AFV
gIyG8LmMm3pPdjLfpdp0NJ1LZ16Yjw1e235YOWwCPmpu6jccucnwcZOwpvN9zekK
2fZsNKU2ff8YPxQL6p/pWcMkwdTQTL6koQeBEl2+p2MyneP6GiMN858ibID+hUNl
0TY9cWBcLG25WtwlgnLaMwpm6aSa+GKY136kTmJEuE7Mv3M5//SmrdTB+1wXPTe2
uQ5GPQ/mXQdQbIB4vkY3svLu6wjrawe+GG2sbTA5KNdBIwaZIXVUyQpSNJDdwmcO
T122P8YhZrC3JW0+xyIOBIVxzaZwp6DGawOGjw43ybwHbUaQuNlwYMg+2J0ZPukz
JU2MD7qWtUisyqhzRb3IA/zRwgFnlufl40Fj7iK4TwPy3eyUxWBygfAVeeyJLXb8
O1dKZkDVDJ24zvBz3kwJcxgDbXqglOU79KdzB9EvLgU2TFWhpvRu9mYIR2+ypiOh
5L2UWErocabyYqvPj2ZO3y6sHFjB47QhVRp5iWUqdQqYtSMAC1Ylgca3EQRFYWAA
D/IuPm0i+r0JDwCiJp8sVqPaoFPrbWxXHXiY04riE8MnVCt3kZPhD/W56iVaJ7Kw
VqIdt5meDm8p9in8QDzUwcOK8QGNIyaLpY9yv3SACsrC0UtyaMODd9h/OcHpd37L
XJ/77U4qQQ+nwBydXsHlN17oOB95ZnXZfZsW+82gWFzCo0qOUkSaXT88GixmUkF1
yxec5x04WJFJEFEmQ56z0lsimnlBZCjDJvt7D8GNzKsHCnVfp2TmxkRvtLP01tEz
XsRARSgnlS2WdOf/lQin3RlI3/cJ4pJ92ExjHkIn9wbFH6TFkAoOw9r95w7A6Sg6
OlOyT337jfIGY0VsPNvlFo+ZKG2GJFHysw7PDNmlSmWCnYU/9hCIaAhvmQD3n144
hW6BkL0bDFvmiAnwGfftOuq0X3cdfifLTR8tDtdake9SxAHtM5WxWfU92wvBYMtC
k04TelnmKNNcocgTPEXbAUtMUE//d3VE98KRgnukVZzORaRIaZkD62WuZGZMmqRK
UvRPQU67NNEXYAAtXJCN2bC5VSyL9Cs2K9mX1AFXzB7MfB7qLdfMVsdo390TtVV5
h/F0DytaGK6H1OgN6pOb+ct+QZXfZVe1F1K8kdCnNNttoKfkvjXWfxaTgkRizGKa
Kc2x2yuZIe3hE8lXeeBzi21ZpB6lAajQO1oc9Knm4+/RxiI2fdWFz5NeIn3ZxWnV
HMWQai975/VNirswdalTb/AZpsCWL4kzlla/kaAdh3iK0GHCr2AnEDDRlRPd00WN
1uPWw8cWtG/kYNiLWCdpybLdLl8G2h6ztCyM809/wStBykykefSCTy9VlmXDs3i8
hbaprOZMKml6hons8hW2NNAKuilHaSGpc+hcx/+T4HcTQ0WzUDVBHq+JKi7OeHWd
4V1yAwo/ApO0rfCffb3g4RcVL9TJRqITNZQeHEnm9P0NpCuJGhTU5e2nCvj+qiHa
s/oq2cgDgzZyBz5y99clJnhNgaeIq5PnvfVC6TYu5BN0DuWJGGYZQXfCHxNO1Bzv
fg582KU4/+LJFvoy9OiKSw/CFabS9nfWwHUOZ8o+qqgWxlzL0MZt/yAw99s/cTkT
MJEwKqabYW62poK6pPp4ity949RAtmUyfl609kS7Ipo5xehtZTyq2jRFX4t9F8Pl
xb6BFlB5Zwrxlf3WjoU8LgVE3lihL0MdXCZSY69jm6hX8MiGTADFqh+lNFrb/6aS
zK/8poLz2moytt7odVtOPpeo0Cn6rNceJBKMWQ1iWqL8kM2VHT4tx/1+cZSBM2MC
Z67GpOG7u3o3/F1BF1NBMFCYgvoiNDgNeAwY3MuO8EVjLf8u7CUmhYNQ/WdIQcR5
L1c2auGl8B68ZWKbcOdYwijttA9VtOERPHKkdj5NWqQLXOlJ5KC3I+U6SWLxkAhS
5iOUueZYAzzIGsdbiRXRVZot4uR/UqUu4MTvXe7HStByxrIUGR1W2IfyjwpDViuI
MLYu8baitiZQ0L5XNwZUuhNgCG2oB2ulpiyI14K/qGDs+GiSZXxuOVTuGT4wkATR
zvzXjb/PVPVJBY/ovHTKznFVvO2uh2QJREfzDAaYRrm+zvc5QmtKzPQRUis0x7Fx
nCEuKJTxjaYw2RWvBiUxGHADik9x3JEuqGszHmowYTrG2ac3uYDV3IkjRWrqZSaf
FBtFZdWB4q3fTuvLCAom5wfbJdnFq0jy+5U4Agtl+mc/I3F4lKT/8nl5y8WfiXmh
HrDWyFLW06AiDB9gDE3W6pDHor8A2sjKA81peKR1EKbWg2bfbMym7Dw8p2fyyN3Z
panrvcfn2wDvtZpuTDpkH+hddk2gTsAo6gvCYnkFHsFOaXfNHCWLsAgrSbKUsP/m
3g5ylq7jZcarLBsVN6x1lHmcwCONxt5sZCY1rdF9JhLhseTTJWQKebNjgUb/autd
Vaql2tC7T8tHZ4p9sxfx1uAE3dnu6EXDrOTvMqi5ALclsdLOaQBSVo8SvoAHJAvf
UfOojk4v9yNVBkDnsCu/GRKYKFkJPpQnevn543L6E0cnIhWPhFdj0Kd+JaVeq0oy
Ew16D2MBaazpdEhZfZuq7+EmiPJWuW8Nzh8ImsJ+kxaNK3Mgr6iGtY0Cplp9Ep7M
euUMzgYvEq6eqz8dwooQXDRqVAL67tiWKLh7XnUEx2VCHqIsVzmZ5rm33/Z5EYD/
e8UvAAkgO6pypnWL5ttR3x+dgLouzzSj73lCGuk7/FKZvyYjwWcXX+u+zskVUOgC
12xASZGSe0uJ/8diLUXTb1pYqz4q+fSs8RIlxZjz4W9TgEXxzxKSVNaz3vEOAi/o
0zi6RCd46AJPm3mF+lGIGey8c6MaJwYH3ImTi5T5JqgCub0or2C0d4ram28xtzbi
II7qrU4yYGpYfP7kWHbgasKV3qZ7MWbmv+Ir5Sc2J+owSWF8cW4rKBuFIO/JW89z
RWb1hu3vKxiHiKTVmeDoDbi+vDON+LqJD5jXfWqUazKAVYkX72hCBj1w8C7M83dz
RM5TfCgI8HplD8cVhTcijinWMD5EzWHS45Oqyox9vXu6XiBY4E59wrGZPQczHyGH
tPueVj8CKH88jUoa9FS7t/tojUbDPjRIZo33/ijISsdS+84zwTyYVrheImeSGJIA
sj21yeA9tUNHsln/YCvh9PrvZydq1VzxLfM9f3UZ0vcxh477qZdhidXVBWa/jy8J
kxGgvz3A5byGEsuFILShY/uqgzrGpilHbPagOCq7p+ZWS3rDodvtWCy5Rsz66+ha
qyKQrHtEbDTmIwwqTwAZgkcN16Bbd3nfM1C/YbuAf0+VZjNGxMrN9Yk2xNoIgi5g
IUjp+X4eYndo21/EglrEytyQ4AKrR6YICT6jbTtyjCmfqUits0wsnt9GBHu3jY0q
xQkVN4qApRFSq9+NgISnslGnTpYtgMtuGXxr1njZexiP+KXsYj12wGBcu2yESfgV
AigmSy0G4hjtUHT7KngHrxqNx7MBmweDfMVIdJd17O311qhIFb9yLhEBCyZykqP7
OVLMeEvARRtm6WflB0O6dir/ZfacM4vfdL+g1m1lI6elXCSYVggGbh42ql+XkpSt
gtIPmgJKJ7F1MQkpZKP0e5W7L/pZ4HWyTiQmZ08FMUHNdBJVba3SrTXz1w2AxVZ9
Q8+SEYFT4uOQjIxC9U08lSz4CvJ17ObyMEf+AaRrJseCrp80QWepWllrm+Mf4hid
6ICTDds0W/Qhd3sIo6yoacvsbyrZXHNrvPc3a41tMJNxyT9K+CwTbTzLL4XlpiPc
fB7HrR9d8UKR8yUHP2aA37PpzdANrmb60EvgRrwQ6WgPP2tvuIC6rFABBp1KQ0+P
sfdxmZ0ybsXfUx+ecBl3GI1zdoGyy4Z6bleGeMAPdJW5Bq2JveezeGvgZfLFwJhW
gjMSmQwKpaAIChQYQg+Rx/JTBPaFUD8a+vD9mPe3My+CxRn6tDDP5MGn5buq7TA2
HtVb0oBtPQOk+weBTIry7CRPyqZrC0DNOjyhsUjPFETmb7X56jmubtIXtZJsN88o
//yj0U72URzVNnBEqoS3wB3ld/hZdU7C6SSXUOCrxg6GFfAwig7YOskBw1dWP3gQ
ZwlV25+6ynn8FF4FIOpAtN9WTJVmAXx4DRZWivfI5+Qj08c3x8QWlF/xzTlpoPHq
HzLN1050/kWsjNXOuqJ70KnapIECUpZD45iSzdP+2OL+F1JWXGCrZ4k9/+zLDjmu
nMUfZWVZWj8khLygmOTaRrZJdBZTzli/f4/atLhOjmcBGFh/koB3LNhyIkFacs1I
o0AgLKf7pwk/llGtw4eUMMbLgPuTvb/p9k2DTIdVdBKP+aOjY3+MWK/gSY0PwgIG
x0ibvjdTPwVjAvVidPt3UR4ZfcztodyM1Pdm/hWhwiQ9dqOSi9BCMZkGPDN5zt6D
FEAn3Lcl3KKDKIRLxFXfDF/qViZDPpdUKOQ1V+Eb9Ym2lkI0cPBmAQTAw9ncbfi6
8ohcwsLm6XI7qk/SvNrYZCm+g36WTYTt2T2ULLahOGGx0bjkBIVHFGHFfHjEg20P
ZZlWXvT443AgCWPms9K6XIwUz7JxikeladlxvVtNxa4zt0DjdXSjrf//5qAT1iv0
BHQ6eJpH5NisQCUi08v2tdrOQpe0PRU3ooqnUFUhjcLwato8ryaKO72Pa2upNCmu
ZQ0I3RXScnT73vS8Pn5E+TLyr+itqJeujUzPHSc64DjmFlQiX8TnK6amlvt1i+k7
Y+VQXhFC1J4ZZXxS3TwCAHhmTiCEN32BFBlVDKi8xAtWnMeqSAkUgzi86wccHi/i
oH6Gfr42lpkr9iIJzCWJwDmVz0Y9jxWKkmZhiLzlU0qfmShqUoYs7iVVBUgEG39+
IMhLBsuftezrgFi6rRcDsD2fDH3eg+K/s3debBadsG2tbhBxozGnHfqtnt+Kycvc
IW0LKYdQuD6mIxWeIOaQS2paImY8TCssunTSU0BY9gc8NnTrhwjQsTSd/uX0yUK9
/5JY4W1dqYgjiCcDxs5ZrLRN67guZGs5SCrWolPIS46MqJVpzXhkpplxJAdc0WoH
NjCH/T8KToBN3wH/5CMPRXfDcnQ5UM3GbZHGvJfHGk03nwyP7RlBGK84L1Mk9mr+
82O7V48OaF9ezSXyotEIENaIKyF0SWMf35dZEiAQPfsQd29zEcP65OqeSfSybhP2
7rhGS69mHNvaaUpU5jdUMwX6GBjz5tVxEB/SxoH599xie8qnZ61jRmQ7SWod+rt/
CIyFoXZ18KmDnVYwki00W3Q7QBkJUij6UEWMGlYq8qMQw31NMITSBQwDfblOCsWi
UjyH6s9az8BvgMHKQzW/FFIjnKg6wum9V3ibUVDln6hV9z8aXgBM0W3yDFr6/fWl
3XgiTr+KZujC3K4nrO5KdFnbbkbtW/K8Mq6jWT+Vg4itNF/uYPshR/EHmJahxmQf
ai9ZeTmFcW/vJ+hi2dMiBfXMVbvLPLgjHAv5F8lsYypCk1ofyAabPOVzhEJQ53Od
gwbQXr7bNAplkThA6VU0ADl3G2GKl133EFF2WkLliqTrMm9GNozxiXCokaM9pQji
FGaQ7H4mRBNlnUMyZyVS4vIqwnYskL1SzlhA5BBITtnwWYfo+Tib9KvwmsLj9O/B
ikUEB/4hO4ZMTuoRLDV/+TXrmIqsFAwsFof0Daj5zg92OnTzgdI+1XSrN8xdn400
JwdASAEILdLO92zSsVXNs8OrJuQwkF9MnJAMjaI3Bg/ObnvjgiNbSbrO8KPUusoL
5RTgbXwBYXcSmBpzR5bc2J7av6UpCm2dt4CIKNDMwOwdAMINJqaPlb13YkS9EtZA
LAZj8htErHJ+XDd8Lg8kYuJxqLR/a5VERUggb+Ctp3VGqZ6KWVu5E3gAzHvkGzIA
O1PifPHsVhsUHE8VDim+XXd4M7Zx3DC4/1lDiTuSRjkEm7Xtmac/txD9/Hv/7pLz
fGj8XAwV0eFOT9yd5MJrn4HYJr4KBgABJY9Xb56gtPIxY67W8xA3Cf1ZVfcnm+tX
DTqRUsVUEOj/7iwDsdqAnyGkDnOKQskIaUxe1p2jo4l/aCkN6uJr/SKhqWPavD2Z
g5f6t9kq56x3KYFV5/9dXwTC4mT8HS+UoMFq3jCx/vxyduTmS4r3Agmal5pn+mv1
UKj/yUJrlVuKjaacfjAbScALJd24bJWUFhtFtgkdxYKj+ph9TeCZNEwvuC/gBkvR
tu9UXxPsiN+gkaZDwRoyYsfT0eGq8rMFRkPFKL98O3R7gLiqQjoUYzn8MaN2ATwv
T8tmjQmjH7Dk/C5cCCFzoFwVYc0TjillXMzbgpr7gBJUROA5xcVDeHm6XY3S6HJe
F2SuaKNyg+s+3C/wSUGwOprt1XtTjNbwkqQ67QmcHbu1hDO8fMjTvP/XZ2jJhlMQ
KShvR/dAwN+1FcJOooBumGiYg8Ylv1DPhCtjCVB5k2tgkP3CzwGkXGMu3thiuXRd
RRGfdMPFnGN9r7k+8YSTxc2+AP420qYou/I5EYAnHNBTFkx6OszocIpt/RKWxXbz
nCKirmhJ+x+71qGsuoxDxtz8X7RkPcH7I/S4X9CdAcG6ikENarL+6gGvMKTX7O3B
Wjvq0JltKybHM0eI2jzacrAhmsHBQNXhiMFFoMBTonToOCuRYmmnVOWLNaBqX9Lx
Pdy+Jrw0/Hd7IqBRLGm7y6L9TGX4ucmQW8aut55kDXt+PQnItM2QeWDbBoB/wWv1
Q5J0Qao5U9r4GeLgqzZIUnYiwkQZw8oicjLSFU81ODz9eeY+DHYgkieupUJmf1xA
QfDhbzZvKi4I2MTYnlgEYNtiGkHieHe1Ictl80EBntWFjrJHE1p/CYBfaPCWAuxC
xDzCnTiVZxdGzeLE2wq+AVv2g7h8OL2CfzyrG/EofXKZZrNXBxwchiDtU+kaP0nN
Vl/6mmmy0qkef50+gLxTkjczscphIRw74vN+hXgQWoLZMvq6Iq7eMbW7sgDtIJbr
EqvSw9EK1GDj6U0PKkoOs28BVjQoDLm+Cafzr+9p2vh/zww/xkA+bEXDTs56let3
QLBpNwuOC1zkC1BoiG8ZkE/ifxwaSV6aP6XqDAlMVEEzpAFnYNu+8J4XUfwunejJ
vnSCtQWWdbU1pKqd3S6gQJlgBhtGrgTaMPt/ZTWGuymDraW7dW4nYZfJ6omlNJDb
DRWQ9QCUIz8loBEbugDRWe/Lb63j6yQUMU8wCSzO330VooReTf4pVOjrXVETqMef
r5DFc38HyDUUad5U24lks9xj3BRqUxrZsW/ZIrg75f7oPHybD6UCyhbX+e/Ac0oM
a4F6i4lws6SDfQSQeG08ywMUrXLdsJ+GckvAAoIm9LkUEwUUKMo7LVZdhQe3459M
x4JLP+W2YiG2Th3py/hfFUdye324OiJ4KsMnc84WXtHoHYWMmgiYtNu8xiwVpAwN
H0jA0KcbiGR4F+eAxi14eWu5cQoD6qtLi3HWcIC0RnwJuKQDhpkBOAGAUvm/eZp7
iFZ5fkQiuviL86BrqBoCEtg6bI+0fzI4z8iTR6/tA+zzVojGUv2dxIbFWwLdQUkn
JM1vgXoywkT8vlJP5y/9WLhqOsrQ99lah2BO25tJWeRurNCsXjRZhHBxJHxS9Oj+
jQlelReKtvxKMmtOttFBvW3nfqw9GR4TCWeX3sSuiae3tsHU1SiaV4VZi2KMrsMF
OMHsgaLyaegxrxh0zpGriynq44AkTxohxTTAt3ggjyyIK4ptjS+srPwp1FyePceZ
g/Cy5JGO7OO9UqWrWMCjeIywdjWawl9NwubU3OGWJX2IYY7VrcvfXuQNJapqM0HB
lFBeqofSatFa6FCJu/UPk2Hq5TwD6u0uKzoc11v3sd8ZXrGwAF1rfXBRdLFJNH5d
M2Rn5ZRCCbcNFrMJ4DdFqVJ74Puo3GJDNBgW08Fvo/fQR5J67kDFRgoWMC5OZbdt
D7D+3dIS4UZprdpivXB5OLzwo7DEh71yB5jtfcRCmGMOKHGlBFd82AK7uuaIunty
JSyXa5JTcuGypzGK9bnsgenDLkyWMzp1dQaanco5yOEa74Hi3JvssOHnGLFBBtKS
`protect END_PROTECTED
