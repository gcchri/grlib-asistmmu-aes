`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i90c8pFssHVyQM5jGwnWYcyExvdE7ex0Q7XqmqjR8eJSKx3e+ipmq/Ai8w4Mw4C2
hQbF9e0ENAJ4HLin5frwqbSknaEE1izXyI3+Mbzbok5NpvsOSfcOjkha1t+CHntb
00V3Xs7IYW2W2a8C3GsIkzFBwia1TzfB506Oy2MNoi57N0JAlZH7yZlM4deSEe6U
5fo6CZ0ksrSBRvgWlBhM/FDAZRDB1AqVZXddfMJV9Sc2T0CGHmoV7j6LN7ix4yMe
/2krT3ixygn4sZ+PNrwmewjO856lBQFtRs8kohHYIpGQ9ArOklPgVAnXLhei86dv
XFXMstrjbmJ/PCCkeGj5xWrIy2owmDxgaebJwtFaENVXaUdqBo9+FIWgDV55Wvv4
6oOj+dsJwEy5WJCOcOt0hLCFBfMQtW7QeZ3OlKdZnHDpr2iDXzVzYpJS7yUwhrYl
/cnujtFr5sadI4ANU4/dugXX34K5zxfJCFf41XwIEbWGdQruE+KMBpbwTL1A9dVF
FqORgR/+DOZIwBtomb8drkBNvJ+j3yEiJtFXCmlpdsUkuk96v7A6pLai9af1b9FO
WkcxAqz7OkK4WjrGbK1DAwz8fl208FH9AryN5wcPORI11VCYwv++tiJq6z1Vlehz
3TpwPzckH+o9NCnn1A7nDT26ASbPGdbBjf0xv0GNi5MrAo1iAfpmD4WZD8R8bsnd
IPb/EgFDJs8V8rO1wERYoOJ/lSR+84W1c131tPyKkXzxX3Y09d6hWpfqo6cldBGF
XDf1DqKpMq+vFHjrdxj1EyzMzt7AMrrpSQnarN3HgeA+yqWWsk0axMyrGhRhxaDE
rS2CHx1oTiBv1YOdad04zWDp8NNaenFePhspKlmBQjBdXm6loNB+xhU9PiJOSuzz
`protect END_PROTECTED
