`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdtesbe0LzGPTA39IkCN9TWQ9TRHzYN9PMvx8RHrBPoPCxUAoDXG0YkPK/xuwv6Y
nXHA3WFuCdh+nqh2JqPILiPX8lZd2oAF5+fCq5qcTgsssueY2M6UT7JEPZej7Pnq
bK6nNTIKmUY64vhB/Y3wkl6Qkypx8gSw9V7QxTvIedLq3XPXDLAFY1NPS1atanZ2
PCg5R7May3x5XArMWVhdkDB1wjmAYkNc9zo5hRgiOGusr79mStDX0QIC/G+Vn08B
FhoaadVJs5ZnwGJUMlp4PVbJhCEhTiLvfRuHd3s59JANFxrQ8PGgZ/0pV2HvPc8Q
DWypg/0VrsnddGThVH1wsPfZqd4qqvP1NuqSOH398VHDY//+8uhsXKgO3nkTE4nl
XT7lde8KpEer25gSLnF+nhXyU1tc3rxuyEzPnGBy8sqSbI8QOg+w3XRlzSSAwFgX
mwinwCh/g7E/GSy6XYlawBDLqOy/zyNn+QdxZf8RyGDA+0BfGuR/VxeHxkio2xqY
SIYl9ER0t1MTBefAzDjp6c4rdtoNxhJHhonnYNZFfzxMsWrB/bARgB7kRTZtL20X
Z2D2GruCiGNp+NUEqhyxvSXSiogvcUEzoq1shj7YqRczUysWrMVvO3qLW+6OW37w
tLgZ2VxuJxjvEN46W9Lj6e+sLlsXWeQk1N9bFWme/K5xENSjqXODEbVIbQDTYPcl
7PsdFJ5E20bMa8UUHC6wXF4mnCpn3p3jM6mE/1waMgqk41BvfFIssGG/n+5uPLnv
n1+eDqLlx6/QqmKrNPFWHT8G60rb8IxntCMsfNjoccGGgr/KnbISBrWrzoDpM4Eb
2gi/AuHGELo4VqpS6shPTR4Ge7AId7+qpeJB8t3f0Y8=
`protect END_PROTECTED
