`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ScH2UmhXFyhQrJI1zbE4eS1q89CqGDECfmGLi+EGHwIoqqZgAeNGWk/tpwpLmTQB
JqJ6T/vNeDtzwjioNfp/2Uv41edfLqo8oHrEc5i9rCzIb2PIzWN3MAtNxXkmt+XK
sRBVXyYCyADrTDZ80hR71+wdTqGLTBZej29z7qd5btE6o6qvKl1jnGMtVG6FZpXv
1JMum7kCISJzxatOiBj6rz5qeicQeGWkPJdL5jYBH6BiI/vExEe82tjQYEmd/6uE
Beuvnr6nU/REu81KlfPAVYdBVUX4YQ7ZPP5pfDoXh+3fH8XXIbz+qxAm50B8WfvR
JBre378R3aVUo+42A5XIihvi4+T+DzZxiRx0xcbkDL2tpIml119MzfV09os+aUie
yajeLkBOsxqxY/OnDt8JBlxgtVDz1B3U9Nw4i7mzKqT0OWNOIw32pk1w5DVgdaDB
t9ZaJtbJOHCYacoP4Zo4bwXMFKipV17u5pb6PspyuwXUFLuaf9Z3czRjC6JwLQ4Y
fGr24bLD0IjjEhorDf3N0/VbPDIsm+HyvILFHZXoN1glOBBDjyxwL3QX+qFTBNz8
4Ib8BMrXq+m3vlikx1oRcYCMNpCgnvdihlK/WIG9oUGttb3SRc7dS6eyZOb8HQ4m
c+lNYZBwLdRV63G5EM5L1BrQvGQ+khrF9eWCG2n7R4p/eaUiDAYuWNSBCLIYW8uc
v0KuG8lwIs6LB04hy+kWL07AHEyditRwQPhPR9UuCcxnuBrH1Tboxa5uvPltYDR7
5O7KtndgPvsDb4X+9TneBhv8SKcOPvaecSTrZqh1sf8KBixlWGtNI2lPWZ6HREhX
sN75a/uL5XmMZAgzwwqYL57KCZ7qDImMsmAE0kIJTMu1CFM6mRV68e/tIcU1+v9c
sSxwHhJLiD7jIrwhaGuuMRy4EaZ/1d8/xaedz5y6Mm7S9CEpjBuBINhng80io806
eycsIKkziYUi7LdIVeAh3uMNpvM2VzFwKs6yGC3uuKVb+0/mbtjD4sNiRxJzb2iJ
k6UgOwGrjRX4JqhiYovz6m5EeH9HVO01EejJjd86A5ityY2ZaFjUwFLjhFnfsMlp
F6X/CKe5IK0am20x2xOIyBS9XQJR6+Jp3nTII612DlP2+TO74vJCBbeAqie2Cbha
dsGo7hPf2dASTRBTYUJ04/E5i2q5KC/sTeFvuU9cRGY14BqK8t9VAp6LNCrAhN0Z
6v2f+NkFTPThK4rSGexzElCrbzQCgy/LT9TfYD6umJE0++q2VGB7f3N4kp0zUJoO
e50TS3zH7EZKUqc0H9LLk99JGX/SSYvHpxPsC56Gy21vDykM+7R5h8/jDvJFb9UE
ZrB4zxRmC0AJBJ5SEFs3LwD7zFmqfX42rHHRyAVaol98jANV/i9F4H6LxCMJdrqO
eBxB2fcl4jKLnjWtmJBLDh51r6cOtpZpbGWfCwziqNmCP+XfzyKKEVhdU7qOTrFo
A0OnfmSrZqpNH8mdpkf5cSfNbNo6WZ+B20rEd6mf5TVfl5vZmuwKhi56JCaiCUpw
3JzabXOR4wU9pBvr6uzMWV5vsRxxDt1kv5Pj26LR7D0R86wvWKjLVAtspTR5/wxx
gNwDxeddrL57WWMHQY2wpWm4hBDgB7XSHSaxq8z6l17o2Y2I+NXusNEq7gbsfsm/
FK59my7tph9S9WQkhuP6GyG6d03kRwyEDZm2n9c4146WE696JrvSGb5lPQLYOgPe
R8wYVmgVTTT7vqQ2w5qf2LDJ1o4tha812YmT3O1O7pCFr67DbD/3UI9VAVe3xECS
AdaLNMIYYj0oatK6+lkzr+KPrROAjzbbN1NDWGNXZDo=
`protect END_PROTECTED
