`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3wck8IF8ET3JEpO32DqS3mnfj5a6aH8Em8nYIhZI8Am/iIOom5RfZfLdG05iUO6j
JXw4kOTdDNUtROMjNGEnLhZkUkDp/ouFK51+vBn8VrJXvIV2q2Xf+0dW1KzH6rBP
EPw8BdakwKR74ldLXmNHvdEfpv3Zh4gEryB50bh5hVafJOzR/nRHD0fEobWEmCr/
PCrw3aByJlHJsvxT516Bs67GoySO0QnFN1sRs7GGTC0gwmt0Kl9VgbNOUDY8Q9Rz
ePN12W9tFLYFt+yo7snlXBDnmTsXbOiGHTLBEo03HFU0KiqMeXoEG9kilWdXn6hX
gUSfu5g20EnT+Th8vtJN+OnDrDaU5ODGgf5/yekKzIqbF6PKxXEQ+GuqYhhbms+3
m+C6YrMud/ACK9pXhJTMVeYannYDMzlpg+8m79VdA2hdM0wV38wAnyRk+YYLs61r
jpjCnX4RFp33It9XOUa5og==
`protect END_PROTECTED
