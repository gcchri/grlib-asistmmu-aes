`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwlaR+w0khUTSjut+PSVuperfDvR2X2qYX1ojnTzbqlW1mAEbdRRScBWW8bI4hLY
uMQQHrUZZQZ/9m3xCUmAsOV+JdYb/iGrzUDHl+OL7ndswIP3PHb94MCBNpfSZs33
Kulg3bKBjo6SzJm/VeGMNMmTDkPLipeIVuq4pk89in3rfH8HB3j7k7Mgc57hNLtf
iIsnJfoC46iZnFxPB1i3sL3RuTTNDBJyQeRo/X0ilCTzYvZqJPkxQG8AmX7X6hgC
xN0z3Es/YU28fV2lL2R+ekjyXDOk26lfef7srON6y9yqfU3HCDhzk+xuzeUOSSwb
dCFCaUbYRBEbUOcGDHT/DTx9eylmSsm8tQ1XJtjKB8qNiom/OG0GnEybX+GIWhFV
kiMqh4iwhWO3Wtxm/8+N5Dq4yNEst5kDaXeXLuq/b4pL+m+A29CTdc/A8Mj2u8pE
bJMbxtvpThUSM9FbJL5gu9Nes4ThmPe9KjA5Wobf1AKIMU3RHxoLI979t8mJaDuo
`protect END_PROTECTED
