`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4B6E3fSKGR1tK0wEuCmdDqrfVZbAFZEgYMDo5fbnTG8JHELEzoDjA8BZ/HmChhg1
U/56UgTfaSCDP5MK6pkuwuuEmn0M1x6GSQQbcOEz93Xxy5Ghj8CBQkFuPSUfGXdR
lujTpqzDdHIqe9ED+3Oh1hxnhhdmB+x3ILr+E/G87697VKOaXofbiZh5go+tEB2u
HGfu4loCwWyseJQD4SD01i5zhNNEie3Jg4xoIK8gIljIPzYNIeN6i13OUIVN3e/W
X/HNnTU6S8vH3xjD6nQpHJ+t4Qjo5sOUXn/GcuZXx5oEyXoTluUZ3fp9wTPiUnCL
uFjlxyK544cBtpoQSvsZiynTeN694q/PurJQKMurA7E33Cz5qnzXoj2q3MVsrA2c
H+QfHD0VJNxxUStL6boEBlpbHoVa2MQu7UUFws7EzVN35DLo+EoRxOHsctJriYL4
Y9fzMsS6Da5etc/OiMHgXts+p5wGGe0XjEo8kVaEZtWO0P0RGWxbXTpmAvEh36Ni
3m0VY84SYIcSyhN9SrHCe0Qs/yD196pzcB8KIObKJMRsI27iYRqFXl+1Q8XVikeO
SZHSZrUR6i8fahKDgi36GqacnHq/jgmB7F9HEXXn3+bvYTNKTsgDY6GvWbOua6qz
6JG+Lfuia8awhu9BCHZztdJVnyIXlUNg0FQ4v9Fi4/qhGje8TQovftJjbxoTUgEe
DwBaHYtg15N7MgejbVGisbbSZk+KedbQrVdbtNy4Coun6u5GIE7V6QaSPpabJCNU
4WoyM71ZQkVSrtuCmRyH6r3nsYPD/jN5QVrbNxhlUyogUTF483BB86pIMgjFEyvU
7SH56hCH8dUhnK0u5PDCALQnBwA6Vsy5IZuBvv3dbW0XhQZ7Z6tiScN0riydeJC/
ozDadZSQV32YIluVFVTq15TxB1/2wdUfptSNJ1Jv4nsW9N9gF+3Nr2fXpmUfi9zN
RDDywu/5RYz6a4pEUI27ArSutN2Xui6gd243gicjMss8xQW3zJveoiKR4W/Wnh35
Y3vAPtIb9BOQQqYAvrgoqC2H0gRfRXL3P8oyp+yyIjntC4dOvdq540FXJZEibrsj
amn72Irsj7Kyz5mrbvrI91oKBK+APlL/972w/41XnHGAImIU9qfzKGGC9+cw+snV
Aiy6pZavLJaMxtTxb5547Mfkt6GIrIa+1REDvYBHje17tnHeo8F00UOUc/TOF62h
PLp7VwcBq371HaZYzsP1RHiC9BQ7gBbNIZ8vBamjxIeVsWtUpqJhdXJ6+59+mRd0
KAkBvreRvz/x11b3ZuXIBltvVbRt4gWtSA/CgvfXwjOP+4jLPZxgq07JsF8etikS
y3nKYrV5VRFEN5SYjecYL4IIQz6F4yIlnWESFPLf8CishA+MVv16ht1Fpn4Q/Dmp
s/BI5+oysCMr8bPSxPh0lxuMLQxWYd9/qu5pkIoaJdbF1Jx5s+74Xxb909nndXL2
6HLuD2VHXiYQEnMMfFTUSiaq2sgs4AzsgKmRXB69keeZFXUgpJeOuH0BDlI1g3N5
9DyqgUwv0BXQMAhcG34HcgS8HBe1q7Ei3yWXuJZozKQu6lVU5ZjKXdMIJPzKGj6B
w13FTBm9l8NU9/OBrEgFFEMr+lBUhNQV5KKE3b2CwTneecIyQlblhYNQIeM96qsP
jK8gM6RZXG1yLMVZ+j4a1PXR29Ez85Z8H9bGSp2M1PBn7IKO3dV/P6nnH2ejvdUt
MkPfowFFHmqsWcwfzFe9D99cHJ8oL6kqXi6mlfGvsIeFTmXsxSSFEWGmdQ+G88zv
Kr+BqUJuOWPOpu98GrT6Ijgy5/oc6hqUOsxaXujrDnaAWDEx2fmUNwB4NjHaeD2n
MlQYN8KoxV5wCZdmS6u2lZ1rbVzZv+Og+jnybCkprVo25bHtsGoPd214nk9zdmsn
Pm/69CF6mn+9kYyJ3fzHggelKZQ35hna/gTuPdF2JaPCvbytG+xZ9EfZ1tRb8Y3B
szsP7ls2/ZSh5TOj7MINvGEQEghcqfe4VEYCefLgXkx2I6ccFt7OLzk+wXvH4qGD
j2lJ37RZ+rzPtjPP0oFuieXh74W3yV6sU8se/VUvQpynqv1KFlGhadzTVnsIU7sN
FiS9U0R0259lZ3qGMeq1K1VgOJMpKPPQbDwJLgh4E/Tk3irg4QtWMXZv2Qx0l94w
taXHlf4DSEv+8J0Wo1vKWXNJqrzHl+eo0GZOWQmoAXQJ/AMzr9Kz92m9AvWzA20u
s/w4gnPdIWg9ELMwJJTJNlzLuA84XGcXUgYRU+istzap9FWorUBp1Ahvitx9uadf
LEVL5jP86lnlglzrtebQUehW2guA/EDeVelvZKHM/xckJ77RjSujhIj/jvbfj92N
Xu1FF2+mE0R6LZjP/4CagMcOXp1Ijt1wa+YnGMSdCtyf92vLLfofX1l6/ifmJiaZ
PuT4mPqU4UAjtcjH7q2dDOeALkuNLhoiKVEKSoCJr0fcEItHYduLb2M++P8d1Joy
LPfx/sEc+mDaj6HDUO9I7GmyJx+hfkJ9prl6zNZO/Fp4PMHfY7R5zWQN9p06m8H9
2RFRvNMgz5nqzNe4YrQyGxBv5d4xt+faB2BkhH4yi5nfRwf44RoPZpTrjxhFB+Hf
poOwhy9cTbdICW+o+B8k4PPxwFp4G9muZ6deqkVc+Ll2Dy7FiHDY2rm8Oo6RD/tZ
+agaChntxBb/Znr0H+KoaZ6/mpllW7IbkNr5erlntcoJLKXlMofv49UL/csrRK0E
Ra4RlYF1gPx1PJBWU6tnp3aZEGckBT+fkfTRyfz0PS/x7Gmf9Mat6a4LU9iD59nd
2EdSeR2lhAvb3IU/twhmHsIJKynFDcJuxmiZrfEq9m0njEMkOqRlrWviHKiccmSK
yfLzO3fyHW/d+yeYq1eO+yvOldH41+maXqtH4I5Vw3prrPv1+DTIveddamtj52In
y+WUNNMUUzt9Vpqd3sC2RHAAq0extjDoPyEWGIKw9oSWVAf/yBqmPZkPJpGbg/If
0Topm5wIod50cyqgCA0iIpOmQRQ1KZoYpNHdnjb3d5G/X2bJMjE++ZrmYjH5ap5s
01kLRFoHCnlEDcwD3tiaA6sRrFtIzdyywC9tDKFQPK/KdgdC8XJlAVHcxIlarxTR
L/+4q0p+MzDcb1U3XDDXROvTk3nI7zhnjNT/9jiB22gnJP/DjUpRfjTI117+qAXs
tTnglc1mFpL3iaAFCh/ljUeCPkjZnfWbnvlHIRb73xADrJGxQYEXqYbAhhe/UFH4
SYz+TYp1d90yl/Q7Vr3I9nm9wh5k/pD9ICP+O7q7tMNTUdXpjGAYOPerGHt4wIJf
mygPwfnf0sicu8TxcRHKqyOnqKI1WahduvUJJvc2fqEPauuJq5vGVHDF5eSzIrnH
cvACE6T81xTMlIEaubDKfhPf7cVq8cMTSmyyT/4znZsPn0AgsFXfm8BK8OOO4Goj
52VyBGcecHQQxmBnVmVxyywH5nBsEjL+3anT3USNrUJuDURxj3e/mbUOfx+2+V0t
y+R5XL/CDIRWV7J3R5vfqfNOmdeupVSbndosi4AbqYyBpp6OfQsAvjnTythqfIx5
NKGF9nlwv35dpAY9nnWVOTGf4utZsajbsW3EBnsc5q2NHGBjZpdrr4rpXg8s8iDT
ikhGqKLgvlbixks9KPiw0lO/g0TL/8WAzCVF/KGkTaq8VvKwHAmSKqmIaUYruasJ
e2I4bcoV6Sk8AgDIKEXCTN8peeCQ8n3AMTn6ywmclHAJ0QgAO1G1aHsCLD9QkN5Q
tM47vHsPO+HFzx71lE9W6/A/KJEDykN6B0NIeHg03Web8QJVX/5T18pGbjq89wj0
zKT7I54kLyeEVnWtSJn5j4+Cr4CUAqdtbS2DNYCdHdZkrsJYwJ0SjFOQHbtvZllp
vMV8UFhupjo7GfpZ+E+RLOuXFeFZCtSxtfXbQg27vVxSax3mIAYdbH2woODs8MKw
fAJttgWSiW2Y/C7ADdALsB2DnsvR0VihwJsjEaOJ3n8Qh5fManb2OXDvB5anajz9
SwPCBI0plNYzB9s5DyY6vsnwWz1I10sFCLQf+cl+K9Q2LSu1Y8se6x30EgtpP5lZ
I2AVm5j1f8mCIHBPkrGLLaeg2vrP7124Z7znHM87qKJ8m1Czui9IDip3NPz2mysA
wdMrm70eFcXV1HH/JHTjZcdDRhFbuuz3lpRfrIdw+jHc/t4b8Z+z5zAtLabl+mBN
nUtmLMx9QhKooEYkrHhfsPN1InFbVgBePowlEV26NLNpFq02Nm0/aLogWNHr5r1R
nEEY1TIryeEvkMB342UaaOgievUI+eGOsVHmv/Y17Jv18spnRDLiFisZSb7Pqzjg
TKXamCEdhYFUEvExOnaYAfRALJhOrCMQSOiveK498I9fXg7w+zcNuTUD1flryY3b
Lkp0+vdFsghGfYeA3QftrBz8fnu5OngDcmT/mAiAHWAGrLBGnppRvICHW2wKyCzZ
BbEPljpA7dNgDHpqskXDquRVIsgDvGgbtsv1YfJc7VKXdemg0kkszFPm0wJ6vp59
IK0PvKpJORQxFIIfgex4ZMRk2L2poXR+ly2DT98wOAn06ERiby1SAvRDEsLLf6Uo
9X2uPUqLxNBeIzEDQP8JLPmgtKUSSIP53CCmU82MlejSQVEsyE2pv+OK/CGjwR1f
8t0EBEuKZMt6xaP0oHEEpqnu7ew3TOj+FH1H5xs3EfloXS+RaBoTwOLsluDo+Llg
kDMrNMRnQdDKIgvZ+3hEC20MAJSJhmqVDd0uMPzmZH8fyqWLAxAw2A6e0aeF/ug8
5VXERCGB76OGYrPOjZ/S/zQwE7BTkZTiR/VcL+WwZyMIPJzCJf0Cdv9af0nRDrE+
0mPAq60ryZPa6zBwnpjF44prgX9/FTGzUW2yjfnEKc7BBZtEGNvqkJr3i5MeFziD
RTvBE3nH808pebM9sMNLnQTU21ma8yIXgehyt4yinXAZb6y3QXFFOCSBa4Da33z/
NBK1Gz2Nf9pD2AcVkLPQGYURCgU4xYzkxspADdzZqG72zFfmPp3MLXbX35PMrHTq
yhenPCkEiONfushitdnWX8H/Jgeh3Am0OoxYoOhoo2JN/ptXOa6Bi4e75lo6LrL5
9J427BAKbRrxVq/6dUwps2BpjXX/DX/HOWiNDxzPOmzeTf+2jbWZCWADHBkdk/Wv
PFKq3R02UDtgQVLuC+By3w==
`protect END_PROTECTED
