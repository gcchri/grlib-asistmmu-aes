`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
himvloSs7kok+Ds34HvYWGKd8MbkUOupXtsBWWYQzMO11j7lNpXyk7HgH8LcZqWz
D/gLBRijdFdYoEVL6pudjio+GBN67NtWCHcWkaWdar96V/ZakvcVUrFm/XKZabJx
e7nyIxt5d7cSQpcNsffMdr0fOpP1R5u7MuozsXVlIQceNCrwXH1yGzq9V3fjyPs/
vwvqMI2W5RVYHuZthO2RT2x48wxMSDABT99cENkS3KyTmQxVSOyVwhO8iwUKUITm
`protect END_PROTECTED
