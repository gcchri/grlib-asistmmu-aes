`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PReHPWDxBjS8RYIgGCvy3Q86Nvnmu4zPeiunHC9AU5LNj3eGy/zFtgF04b1u5MPH
XPbUu6v8iO+nMLEU8HbUfR1YA115JxpxqFtQtwD6doaVg/3Q1CSv3Z9KHndAiiRv
y9DAwSqlOjQ2RCrXTh9nit6cOtsCURZR6LNORyUivrew681wcKQyV8QDQVIb2vUt
4IuUxIg8IZTskbRJGoJL30iQXzGzqyHBMP6BGLfd5yc5forR11JMuBimls77tF+x
2xxXl/8zqoOtbjge+O/KNOjviPf86dM8DzIvHt/n/00qeCkpP6r9LMQBUfTfSSPU
mm0zvW8iz4bhDdxEtU/QsqFXmGUhW9swx/Hw8ZPEJmMPlzc/0j/F0piWyWb1m9sR
Pz9xhf6CTPuKA6S2dBlCrMIRk0Gnz86qHi+QowxhLOcImQZBtt2EvusUGT+AJdkr
yTzudUWLqfEVALShYfUwHfdUEtGJYcH58dfhvRu3dDBXT9sylMlJ+tc+q238RF9e
wZU+2QG1cyqtB3oe4DhXC00S+QvLBmWpqzQrKutahcv8v1z4YnbhSeXjEWSB4FxK
SzP//zRvTILADJTDudOlTx9JgH11TxyvCogNTDAkfUGWJqrT0dz4FizJTw/QfIIE
A+ppR/MySqCY/tt5gR7WWYkNU5AORtfEVY7btcfmVC21ovAXIutH2Mr1Khx9NRl6
zxkimK58sJBPHBKmjYOR94MP/4nTa3NkssOZQFRVP5RX5Roo/mNQoYPzcnr2zIAr
1W7/1u27a2NDuKGyOBnS+m1oc4+lC7hdl3OdwEGT9d5mS2rfuwBCo0w3D9CzcvFd
dSM6DLeu3bnKqMZco3cODw6r6Sg6qncqT67sqC21feq+Kd6CAEA0u9iuaiE3/22D
oqDRZQ0b1/sL07hYjDzDXa4n1oUx21/U/KTjVj2frYK698/ym1VPSyEKNvjkaH+1
0v5tNCf+4vVXex3JnPyMsKO8aIAs9dBpCaIm4dphuSQNtVggRvuUGg7trVbt2cYe
AlHoam6iIzGemrMUq3Bfy6g9LxMQSIZ8ICs00JDr7/XXo9WYcIvJg7FYMTRi/PMK
uywM+eTLw8uareEFObGCY5PNmmDJTpt+lg4oTSCVDaBkaNXBAT4ZG/HeT9SIl03U
b0CWO5dbJdT5+YjSwZJIsPVIq6gLx7V6gmW1LW6tZ1ljrNrUQHx6iE45PrIFNc80
1zRgkij44VFDd+dXA9UAv/U1xbsHG9DxJx/O0xAyECjvyBn3ULwu7o42tSuhJirB
Ex3z7fjLNheBxwF5qa/XNBfVT0Efb6CuqIowVvb1GhCfJ6UvycvYOKRE+UVKXDV1
/90UOgb6+V/o4mS4/Ae4dDYUOjo3nyOq1sxRz85dU0QVZC7LwIsPw5PBzgoQMZnx
yfl7vX2cpuTDQuFCVkDhnCRCU0kTvoPf3Js796QeocWQSqmDXlgAVZfSOpFAySTm
x5xJle2wNPooDqGvYQLsuwZRqxyUL1Sgsnmf0nXrRiVhh/Vrpl+u4WrlrDk8qfM/
m6tVhUR/RQnU3e048Lxkww2x1X5TJLT9dDCny2V/RCzmPq7yyZrSJgIx6JV/B3fh
km07ww8Uz9s7uuhKTqIahUrU/EmVty5Hg19y/IqfXHEmHTp3iEqY5+9WJgH0DAxY
JZmeeRvdNEHwnnkUMWbMMm8huuDXbjN8XenNZ8d6XNpEolTeKJGvjh8vfWuHpTB6
/SRVioq+vgo6q+01OXsIHPW3ZSokb9Qg+GQUdGq76Z6Hv19zZBt/qhlLUm4M79B7
nSP3Ssc/a4n27AIHaJKYh+igmVIUYKRiabvUWP4HVvZR8/CYE40pvkx5S6Qf7MXA
RAQcN/TZ1CMdJpUE8870INwYLjCZt0eBuE2W78bmAoZ9/APilbnTEBMP/3lBjQdc
DszU1QAokONO7ImwbWoN6PUi/ih0fCF+YyMDw52FkvQ68ah4h/Lk4zDZlSGx7s+Z
Wz6Fi1oI+Pinq+CjaBe5UQkiLjNWudCnOeOtESyIfhydzI8geutxVWLZihDHzjMl
8miS9+RJB31AfcRkHmmadT0mgn3oUix2rlgEr6DGArBHdWcejXCn75gp9RFYH4f2
jD+YQynwTylX1COayHN/a+gWCOEEgYDjl9TDLuf3Sct/Q0EJd5U724Ru66wai7UW
JQLOWBjTBTfvfgcDA0oGFEP5tXmNqVicjBOjVJk1udFfKWFzE3udIAzxdy1YdeBN
p1vknV+gIqJJpc3R3KO09HEhhLPx9nlIBWppzX15FPcwZf5x25UbINh8qKHV1XLw
hMe7N2Czzofc6eMU3XrlS9sPoA8/Q8Klr3xz/pWci9fx3pnmyg/yjy6WWH0gsk1A
xxzmnjGmvG+1Jh+QYy4TA7+VnoTodpIGL/nnxvHx4y+87xadbMDVj961pRfHOrnV
0++eXezX/2h/HHwTFrYRFEcrvwGlmlreCm/NSzaLkCoOG2ayWCUCeUSxdPokmfFF
e54KLrmbls0tT9LLEVg3ED0ZQE6YJIPHw+CYdKD/VrdEgKV584TqMxB+17T17AB9
CIySUUK8thxUNcwIHXHvAEHm+ZnUlgLWbrL/JGhvzwcTwbT7Qxmy53mFKR+lqzsj
SHsYzB57ZMIgFUDkmIqANbwcfzcnYXVmFHNwhFXTowx2K/T7e/YDFl7nVKJd8nf7
304itdCTBIBEIthMDU3j+yfkBLZkZ2XdgGQi+Byz+Dq0doN8bpHnRcMNSMPgkmSf
LJARlt/WJVH59O9EBe0y4O/SSqy/+0ZhFJhpreRwuJ2gKHGpvFMEAlDBYhaP7FAD
Y7RSUMxfvgoR0QVbg6K5HHH/8ArsvXYjO+y7CYTIZtWP7GMAbbobXMUpapCyCRnx
gYzXmjHO4grCKfLBfkCTQm+EmnsJfssNUMCvRgm9ZHqmCwLAuXh26nxFItjQhE3c
Nc7CqTuwncsu0834LGHZ4JW2oYpUJam/7YF6JkU5Jd13Kwhd2dk+3Uw09egi3izb
AHy55u/W5uPOd5TwcU+4rbcQ5Mg32qMD5LWTkTxHNrOHNtOh37Hn13E3oXCEQGCj
viVXFVlSYgGn8+Lci/S3qptUTNkeaOE/32zSwu3V8u45GqC37VDd/DzJd28B99VC
CppPArDfzoqMuQjIZK0Tbj1IEiCPT2X5MQA6ap1DCRrd+fF8YKP+FtStjRIXe/XP
U6yJwotJQT+nA1GgHY3IIDcruAFP0LsYuMZLyeMvlj4ROMWghwYt+KhnzBuoNwAx
58yFEjdNXodHtk2DbXlXpPJo8kTSPKXcr72x6Z5SN//hTQPxrEni6+65KxToZc/J
BQVvT+dg/4cxuFR5067/dJE7OYAeDUbSgrVCbt3J2SIDlLzK2+mXW4pDqlBshVhs
pvhxAN41ShvGgS9+76pWN6TrCmvBqHrj031FGz6QU3dDsuKuaQ8+jmHnqKHoIvxH
6gh4sXKPgMp2xPg5lUhOcCDUxZrw2JaRxUTh/fhzCFtobFKdU2t9cBimXGoAVhLh
bKS3z7oMOYuetx/w/Bgl7UG04A/rGLlLVnIadoFdHOaiJOcGuLDXU3p0P589rH7G
0w72eS4S95eETDyn5/AE3CVp1AMutMNPF+cwwzZhStz/nzMdXH8CQ9Vk6qbCumtN
mKizVf1jTIfv/pT4+G7+yyzm8lVpEXltl92IYteAGzMIKasG9EmlZS/CeiNAlT2G
Uwv2hjlTtBAwD1fO4Pu6Radfz1mvEQ8iY0rhlRDyzl9d/60iIToLwaa2McOzpddv
84u414vMNISqqWYB+4io7sMn6zHp/9EVSeCaINlutPVnueXr7WM6EQ4OOToRL0uv
Aeqn9m/g3U1VBkPTEbND/r5F6tUkDqwgRqKdyKhBYRZBK6yIqfq/r33tGNGA7zMd
vPgTxJadl3BeKR37Qc0b9HnsIjJIECmP8TjGp01fqo1L6h+d/H2620R8B/LFzPfO
6/+2nmNTXBHZRig8dMProX+EfjbVQY7nmUO9XN6ukcEVFpwvevJR+gk1M4kTvNdg
eXfZBQ3WSVIVAYKeySWurdIdHD3bzOxQUU0JvE42nfaVfez6Ke2galYMkMZtpQNK
rOvrrmUPk1VqtH3F0E7yGLImIGoBBzABlhazh+coUUPPB4v5JMGko6ZP7aX8tcPO
Z2w59c5jtwWVO4EJQxIJP3gjeXPt6OCX4xL+gj+d/ybVwFWxhrXFkZRWDXrm0B67
cIUSe2rZQecmORAsNxJ+0rUEnJbOx2EcRwWYPMx1rkmZbC7oQALhHclvHWazoZaZ
Y+knrMjO5CBxHsx+43ZGYkgjWm/6+UJ8xnnPJe48cVmylG0vLSqH55/Y60jcwpW/
M2KvTllHY28Fnu4ePyIrpDBiOBmEhQHfqA8lWlFzJtKm4XhiLdxzsJtbzkv+ucAn
Ax56rnbEheS1Rm4+nGinVx080/tMtWTKOXgEYF4I//3FWSHpyajTQv6kqfJFcWe8
GWk40n8TT1KAyyFI0pT98NHkHALhQ36FzLzm7z3KoVpEu5OR4r60Y3iyTbpk8zVD
cbXvLls6g9gZgBN25Ixtdthy+opMG06/ELGiH63QIJNuH0mxoVpxKtnUHjytBYHx
L1VPtO/U0mafH77kPDOSYkeeN+uqEU/wE1FG2IW0TdD1jyRo7LG3bEl/KsgpZ/z3
OXo+1vagn7SIPwAlDr8ph2fOBlsqu0Ht9ir2Wddef950AJJ571FxuNFPxr16NrHo
7b8GzpCrfB+olAlMHdI5mIXy2lzk2h4JzZbsvvkdipwaQlPvlzrq4hdNWQ8dl4Ci
gaoGlRVODV0r9JVNq+3/1TZLqxF1FRE0wd4DQ/juamrmzvzSdnirp9Lr+I9wHVy3
eKzNlsbQD4THjRYSJp8hpdHJDrWcxk/F/vGV28Uks6ysV4g97sx4UTEyu1UU85No
FnRD87DNm8FsWZCUdDEZLJ6F1yMClQ70UkojmjptyHWBrGunmpiLyRjgQqBUK4Cl
AsedSi3DbIz8K2xAQm2ru5J/2a8SNohds68GU3mHqgpb3krImAYv9SQukUcIQT6p
6NKlx9enHFUObDjgz2t5cX9SeHNfBP68rupi1O5kvLNNSC5PYx+66I0zFLdAB61I
QujDEH/hp8i/pzUawnDqa1YO2ruSR7+qqve05PY/U5lA1WmZ9s95jWo5Nvkv8/lr
aMWTEs6+AvRQCf95sFfFJwW3zpJ3P0jOLccuq8HlSsBLefHlPFr8equXjUDBslSm
M61DuJAKPskKWOBKUZ5MToEEbaTFm2NE2ITDRXLRSUH5H9H58/fuZRrch/tb8uZO
7ojZVDRnIm3vvnRl74TZ5uZhhFPgSr5XB08md9rktcM1FqGfO+MHi5+rWIzjUgVN
zTiPw3EATgCuXAXAt86iQaFupOy+9rO057AyZ+iv2qv9MbLTtjqulzOb+laA0lG6
mhqEvyredGTjwGhuvuetOCLniZrad1lL/w6AUPvidP2r6mb1yhaHn+E9hv3W9vR4
kdmCYeg6Ed1fhPCRMrHHPU14uj37k8L9dUCJBW4oghim+8BuEkD5YIKJ+/vHOdLN
ErcFVztP/ZYvb3j5k/pyeEni8b6ctCGhG6ZxOEWFkTFpeSbK0wWMAAKKMg7WWXro
g0vvcKmYY+xSohKTv9l1SED6oFuLL21HbU+S7i9C+YDztw8uRNa4GByD3h+iRth4
MJb7oIhCwpxBATTrth5PW4ALYCN/3n8Jjf8hGUkYbRbyxaZQzqqAEzkAyzkJSCjI
Si/PwGRix0xGyN3P6VJ8I4aTc2epYZiOzGZ6BfZ1dQa+PlMEPmaTLTu54Id9fHTO
x9C4rW2k5E6ZPfNaVTcX5sUNGQHYOq62lrqXDp/9fbEoRdR5/qT63TROrhwXY3Qb
vEO/gJwbLr9M6PQqAPtbxsMKwaLjx4x43TAWlK2JU/wOoFjyScTuIgLfXbgop//S
Rc9SZ6US8qCmLRkf5Ztz0NRMihVlv5JfUibavaMVTQ5PlJZIHBKAtxruEub949kV
Gn+CITqjjs+b3arom7ZfRtqKR3Bob9cwVMYXZrEbm+lzXs7p5Tet8ylWiak0Btqr
8lgCWKWQQAmxFdPAYUkrDhjPW4SBZhtkrXJg/Pi1cBrXwJT0wRgN127IxMDev4on
DMmuZYuEwXQQshNyCrZvcumYM2qYWV5WDhYVEvcoDdmtrLDCwJyUVvYBL2hslOna
nGfgUSuNd3FENxhqQ2UzQ4uDTNxI6/4zBFQ1J8lXyO/fflh2EXJQCsIt/H2cXsjw
m1sap8V95nc3PG7P4U+zuQRVgmP7JkTK+gQ9d6d4b9tN3ybUwcJBKYjSJM5djHOe
8WS598zgX4ILFA+8Z/cA5Vpl3ijsAPCjnqJUuVglIH5vCynm/H2VbKlNtaohQ5X1
L6VOcLZd5/xpSFnBMMzMUDaLxRHL0y3Pr2AyhNjzxchTPEm/v+n6eXAd8xfoNvpt
ck1JfRudf/SE15BeWQN6zVaUsh/4O4fj7yWWEJ5OFwcEZWhTSbasuZTO8kkweOdK
gzf0lC73m8Myq4BxY9v4xFm+SQjGSb9gmvOHhIhssuNUZNMTYWX8Z9bQviFiQE2g
QDcwvwedNWgN5ypulBLPd/FoiZz1SPyGihtwM3W2uODxOI71njx6nDU6wegqa2Ly
6tXbG8fqGlCXMs13HmpsNBrwvEbcHxPw2ped+eb8RnnjcqVDPgz++RUYUnIop5Cz
cI6AXZBQy4JYFp1/s34ohbGtnm474anoGP41C06mhLxJGsz4Pe+fPOXojMgi2jsS
RLT5726GyapDNAy6oJ6QiAtA8cbojS9WACBfemI1aQpSzwGySjGI9MV6h7PWhOZP
9KNnq16m5/mIZIJ4z9f3M65qw5W2zjLO9k3Xj4KLvHLT+f6PRxMDDZPyWk2MG+JI
SIaFuB0wiZO8+LBvjL200ojP6QXvkK1lCUVghmvL3xG1XBnoDucLwXjAMiZ4ylxc
9PJrX6j5PjQncw747+EJYWMDZXRyZYIY1YCyfgK5l3WsNeO5DhQ+HvjN2n+mSkhn
EOD1bj4+NZDeLqoV4A0cj/bc/Y0/D8Io89sIn8OctBhqqrAdtGrMRXL+OgK8b3nK
QflC/T1In/UUDa76mEZxymWGv+KhLDmHk4NF9oAlfL3S4UGmKjelCxKG9krrBD4f
Ku3grjwP57LwhIOMo6P6Mz+IBL+eW2FQbqZOLP2ar1Y1Tg2mS/pKbjmrPvfsFur/
BVbObHZgLtrjcOFlLKLvbuIVxbhzshkz9I4IefKsj5D+Hdk1PwjzwPGPqULkYBSC
YS3aWHoyvYFOR35py6Mxf4U5TISpv/UgRuZoquh3tslsF2Y+AJ7CnucuS7akF7tV
igFHx9QfQEnVEOEDW8fIUnd0Z5HBfukFDRkQKHxw/n13GdpeyfNVlFyUE7eW6ZF+
u10i7r4JpYaA0sRFkNgk5FXX7DmMcK4ksDoXF362cwv5ZoD+XN9P6P04SWlU/Exf
tvNYH976lik8L6AfenVsSM/Df208ytajqVwkqLNQJCUUvEISsq/hNlqu/MDTPYmH
ZVmNE1bg58mOO2tSYp1Pg9kqmYocNie+lc1x19iV7ozD4cG43MJkSfpEUnxiXkHa
CT08waKenjjoQrcextf8/ickqHwRkDK/JBy2PV2fo88LoKHu/VNRtu4Yl3QGUnrU
pVS3xzOEAdDUpcBz5T+VcHkmm/reasygkJ1ibqYyrvxsaajEp2GPf55sA/KUQnoI
PB8FmEbIbOX5/4mD0pT8NQ4xvPC5pIKMLzEJCFkr1IxBMw+BVRJikQRTuL18rs3x
ZiD5B832qSradmed3fv9l+0Ltxf/ASOadxoztMImz5TfDl2vY449vsqFfWiazbWI
2//Z0bIhGnSkkUVC5TpwJS+HEJKTg/3k5lctp56/KAieRksuLELp1uwqMXwgraiK
Ehw2xZvKMPhH+6RJhFB/4lTCxQjJhzYog2fpw/LCPCwgbl1Zu2yW6F92uqvblSiI
KdGT+yG4klYkfRA3AHmmrlWCmncYBQzogSYPWvy2FO2oaKldZN8af/Za8ALLLvuZ
EQtCK/OuGSSDTH1D1PZ5M3QN3D+oSAO/S2Lsaqrwyf73aB7zSofYgI0JlLIhrcrX
SvrMR9GvZSEfC9aYLfS+WUjFkJF0g2ykGs9v1HHXhQOOg9XB3sD2L6Ez1FPug+Lw
UZOcSfBnHI+P5iUBvLgfLi3QPhpE9qrfGH2oMJo80AUo5Hja92dyAKnSsCt6TgYs
7nKtkIYYQ3gT0m76zBoy78+W4aUmoppLdfSbKQHarSGDxZ5kI9Z1ViBrmVsRuDML
r30KmZr+oyil42lOZghy8CCxtpoHNlM5UOnA4n6tO1glySu2T45gz2siAEqkhEjC
6nFdYc6CPVmGTL1gp42T5D2JbJJ+nQDeVFny0JjgNLRMLxWZE3Y0kQA0WdNTCyun
XTh0lyuklgvUuwoqje7GNCstrb4mn7PtPKzzjSYN6xHBUscbOjfAqtGaj+WK+Ii9
63iXc57+Boc+5pmXDB6t5BesoRKrHX8Q1xUmyuNvU01ugfXKl5/l2XZM5ysLLYp8
teRX0uZGcDy3Obub8/Yx1UHyjgkVFSrvujCmhBwQ6cWHVJ4YR5VuNGXngXmxt3l+
TXtb3U8G9FlrcYNLFGeqASwTaNoqF6EX9bbk/zEKwFSHss8PxRtSDEItImtLzi32
PtXvNpv+qoY4GRoDs9NoiAdXZI3wk17R7a6LoIccnJOC9BkEqxkUkBjQF1hqx25/
jW3UMt6HrGk6b4/FNMxHZGeWYMnGKXBnpH+XFVz1wT8U2mONQtqgVLRFQVWn1VUl
097pek6HeTJGL0C9BL0HnbGDovWEtvedxDwCU+5cKV8enAREX3xW0Uhcg+u8JVn9
eqSolFy8+qWFYVpNxxEujckEscCa6KVUPyG1nFSzoz2+oaxv4d/74CaeNRjFHCFv
3+rbLUCw+XUhv9ZA1eKK4asquKN76OCOFwY2eR0xHrmZSZO9uQRDLBGqEeDz7Fc2
9STVpXctTGbT4mcD2wQuSDycqlmtAz5cxhpTXmyBBK5LZRnucZiwPYyXI813+SdL
2gzGsmdWuFmQOYNhc3Mqr6u/dHsVMKpX7+zEEGHU/Fxozf7LJH7kWTAoZu+mQBVt
Brngn/2W/XO5k3QNLkQppNu8+czY0eSneprs9viuZGqs70LUxbvqaXBpylh2lbvd
wpwMImejhaMZ+IL8Z/B+pNJxSrDd0Lj+zPCcVX6UowyTjJbZQCiTpAad1Rc4eBLE
sjQBZsi/kEqd2gQgbmtUdVailxiPZklQqrLNnrUpDpq4B7k78/F7ESlhObXKLv1T
3q971E5jNYR8ilsGDjwPLaOGv8AToHFQ+5Ib3RQkyNAA0NAx1YKwj/5EHGCCAovW
n7Sf4X5zCOD2/nMt23blsU4mT0HGGhFVYUM0Nu2ZKjunml6oZwqRej+RBp1FKMj3
NRYtm3DvtF3w5XuH3UY4RDuzAhlgha9Y9j47PA3xj80W7G5XhBTwifEw6G1fMkhS
SxOu1EqBZdeNsN/M+w9TbO5bPpczq7DwnDiSEg3TjRIPqvCIFAxX1EpsRz+dlVX+
7ES7qt61jk0KaCJ+lUONou3H3zjn65i0jLopWoWTWMgYjuZU3RfqMMe++7Y4qX09
L+mnMG4j6Z43y93ECdcvFfraF0XajAqCd8t1r6akuNPJWM7MfeQiRA37gmzLQdks
hw6CEduMNiNeNbfim0jkTeQEi9/x0U/mB/GLLrWhY0WDEluNPzMbCkCXcnBGZTzz
cnsREV2wxRYbPn4u1O5PIfTt+H0hmCDWBcBXvtWPxIy9LfW7TZDvx3yF0QM2yPsY
mZOOBkg8GwcVHOFadKx7D6jC4oZuCQ6El6Y1XnuJXitLO2jMMzg4NP4W8QArLY/K
X+BXA5PkAfTKURn1VO/2/BsrmFTN9FnuuCfmigKpYdYiks30qnZQVYYzk8u7TJiw
RjcWZs4PdFU3UBHBeVBI1eOmlHVxfygwD4QkHKZdp8e63Zli+cB7vV/+4gunuT67
VgElwr7vsMjOXt2teeCMdhlDEmK2A47HkdPsfficZe83ktOtHlSWmpfio5PtVhSl
C3bzY1lPo1aiiXkDg1QWgwYfqLRGZKdoKlEX9SVMHOJU2SFOTXboYgJLPcuNotww
SeIa95XaGrU6LjGM5HSsiAVSZFYzTTbMDGC8nM97/LPaE7f8TSzdI77kSCQ5IS+s
l0uN9rNmYkeqTb1qzUubMPYOpkDxLRDFz54UH+yEINBoHKqAqyYQMsl4w45638pO
hddyfLezOkia2ZG5NgDquiomUOqwz0ph2FurcKysNvLoj0SAkmCz5aaJwlj+kNrx
mvSf7kYQRkHKkejTSq+uksCaefD7bsp/ngWF5rORfpB0hXsD6F6vtwAOih6VtpXV
ojvDNNslN3c+QNnD/K1IyXGmsHgWErdhekyrpOobP4LbQHFA0wPA7zc3NnQkzfN9
PH8G01s71XPxbzuxezWfqIpSlLaS6NeSewsq2MUm0DqAFaUR6RFSx1551Dz/07DD
C1ZZAoHsKYI9ofSEWcDZ4rWtZPhTHNDAOp0ZqdTA+ez3ds5AOah4zl9aMz303CXa
so3sQoluNkQwRfePlP0SqREKs9r0bhJL23pwjEu+fIXu+JcKxfslPaOVd3EM+ZeO
En36Quc4Da8QlLNpK4kan2ATi6bgeLVrQcwPQXbT+ohNtGMZueJ27avIzITIi2PJ
kKOSZ+36GHNw4Qv9bEwyYZBmdPa35MzF8CWJyStBzrzK/lUYocbBaGUwHcd72Jkz
2hCp3/GJIa7zyXdrt1V4/AChAs8BQ8//Y/uGphSAOlF8BI4sL1nv4MbR2/F2glJA
UqQE12bMXXirvu8f3AU6G4GL35W2MixvXGYN+jyihzA5IUxuSLyIilEtG0O4GZ2N
LouMCXZK86COzCQsYDJonyZ3hv2pZHldHb3QUuhKqAG3eM2QopSh3hjLgrzqJ1BP
+5OifSSftRTR7avBAG0go0V8Mi9V+eFRruA/tb4RAbHPykTemZAeNC+//HEGMkMY
3BYVI7lF56wFahfg7LuPbgC3fLvromrA/vmpkvDoSPY7lT8I5/wSle7vdjU46+Nb
RE4BF8lGtbLnrUG4uuxJY6u3zD6XtEl3v2u39rCSo/eAdXGEF+xxMw2nllAV0AxL
rfyguTTOEMM7T8kWTm3czuk1HvuMyOCeoUtBqIh+vr7Hb4N+FZu3mpNt6spCBaPB
rwdPcj1n40dP3guoKd/PbwQ6cokGF64ARfKKgSKoC5VA6SOlIK0vqFaHr/nYdidX
9NEVlfRrTedDAyRkuEFjeN43ZIhSHXXYOq/5sS/eOWr/YuQ8xjWqUq77a8SMRD1m
jXGRO5xBvK0EtM2MupAMGpXgOM1PnsVueG5C3+wiW2Ns8s0Ok1KtBdgiM0SbOOIj
mKbDK9q+GxTrZS/L3YivFZMiaSSRRWNh7dPsxBRSavNA4wCGLgR/nVlWRxi+4r7c
meXgs5E8hlNL5XNNXFZTq7Bfc2h8nRcyHg7dPid039uCHtZqYXuYHkJAgQ6G8mLe
/YYkvvms6fI0mUbkKXh9ZuSz7uQbQaKQSovL2TM/1B5iemnEFW5WXIxzBIq5RhRA
fi9vutUYYzPBw5pEtkMfR+MhkU8EPUtF5Wp+2N9enxbCzcAmbiT4pfn9h1ltN/dY
MiWsZu63axfERERs/AehhCOYE1tgC8PKM4veIDqVuLlYgj/TIJTcJExOF3fMGv8l
iZnUZTHxwzTBI+wnfEBQO9Yde4S91omjzobkU1sNw41JNhXuT+WZi4Q/weKpXH1g
TMTsHZ+ZZdLVN+xg0p5QCG4KVNGm5ICo6peczK9/Ujr13N3izOQ/XI3kDvvnEozZ
UjyorGqzd9y6XQa6oq89yUgK6o/lJSryJsX3odjsJ69Yti5czchowntODKnsMwYJ
GFsFMBWBgZtAZgbvnNcfkEZieVLwKZx1E1xZ/Rz9bSHvwHyzK3SOklZIlFtRBjE9
QJWxCi8vpp6QWkt77BrlGEAE2hezwTD3FPqUpCx3w+lWtK3SiKX6wjoZYFLZx9pn
UyhCXBJn7Hv8p9QbOYa7MvIA92+108XtMCswBi9iNBwIJpizuVtrQqei1KViFUER
V5zJtTEvQglUHsrKsnjuXMupuXl7Tv3fsBKeWYViYi9s1c43WgS9nSIsg6fEYyiE
n85c7gf07PldBlTUMWTencmQzucODqR7aqIRvP3bD4FdY9/Adro2QFwpYn84Gt2X
gzTtAvqDaMZGV1hc/lG1C1lvtEyS7X6nB/We1kPf3ME/UURjpKU6GF2AW9jk5e9g
5M0WMDW0JWG0VOTufrDda34vupPI+fm1EriGhcdkNOSMPLhRyahP4vXGeG6XdFxb
a0AFFK7Tdf3TkzfsRc4k/D31uOuYBML0+VuJ8LIE9TeroQAz26+OYnQwOWLRixft
ho8IrtZs/TbtgHUcaas7UF+r11F1QABoiw72OnGYStLQNdM3kBtSXEMhDdDvRYkf
lYk/4znZPLjrWKL5ADbh7l+U8gBWOMiNCDvVHh74OnbAYbGngj8ZOJ1L+UZGgufN
hJvrJI08vjv11XIRoToi43yydpajb8WKypZMtoBFvmAfCZItFL/r+IN1XMCovlf8
YAEjIjzEc+MYCjtuxn47Hrik1QWhEvJMs9Cd3aMlcEqhxV8x3ZXt8KJsZcBGsl4o
lXk1yejQlx1tiA4i1WI9GzYZWtSL6CsEcTbEYY7YNttK/ERkGhfye5Hr9EIdCEoU
g8tajexeedSE0jkBPHqcJwEuZD5uZYx02DsRfUau4ccNJpJqC2yhrES3T0/RL8SI
+6CeRjmH2GjYDZQ2S5bvGwu14o+Lk0qqG7yzOS0/JmwugDamNyg6thAqxCHp6Def
OPbwD2az2QUE0ODoOnKCScgtqDeOMAY9TkZACMjCOtRxzxFgnfairzSS73OqlngX
wU1hHZCNleXB0omxMJnJouQLgxUNdtezKAWa14GqtOs6MLFUWuUF74859tyc/kcO
Tov88fwUZonLAZOoZ6LDAEfK38MWtQaeb3cJMhgUMJsIp6JbSt9ylJ8+BFgoVSLu
mNFkKERH73fGCzuZoTLy5u3FPLGm1p/8UHv9OIVCCG8mAM0XWV5oIVeMiBFMgXFr
27VmHrjW1p7LVaiZPnmpGasOrtY9U29TVQ0OOKWvh8CHUgPJ6Yz3El/RK0bAlvhB
cEw196BrBd7wQmTvNXdSQBYhotSy6828VGIPhIsA82c3XQoRoKa5NYbJTHNsinp6
w7gCgoKcfKP8nTh1gzRhfNsQsfMtq9FMuFvFnaBNCOipc0nMrQL6KeG4bbcWjdg/
6rNnWt0jjktiOy5zMZFHCWzgM/AYWRXncvTdJcWw0v5geqnbbn0yFK3EVyAAUzKW
GuetQEWPsXceAxpBboYpxzMB4meSGS1gN+KjO5uhj4PVAM/3lPzmHLVrpiN+KHEy
Ck3KkuDfjpyZHrnzgbqLtNQQtQOiWMXt6yM5Ww6zwvZqPay4JHlxlpju8imsiUSm
0iW/eeVf2nKICfIwH00uReEiY3r0FzlJtIdrPx6ZLOKfEVvo9DUOJiRk6RY4Nbms
gvToIVUqas50kbsdvo40gV8PczgOBRxT9+at/rlVjHF1V1xBCa5T76iJ2V/l4dbh
vlRDRnBOrt24RggKvAcY0znIzU3uGm04GiGa0rjth9PQXjPwiL1nvp7Hy/M1q+2/
iqK5/AllfzG+WkQvZVHp/IfHQL65oDw6o59T90SfeyNLREeUFPqbOSVp/HiIbYuN
B2qOtT+mjHPoQnckqlNe+BTPY6GZZ/rABk5cA3lrYVgpVQmiqFkXEXFpRfyvEXqO
TJCTT1thN8mj5K/gEAkJc5HhkLRZoMcqEBk8baJ0g14alYy3tlHAgEFxzsJmRM8G
/8GStRLi1wFxdAsykILPtjrNM4rvswkGiYi30LYOwZCX7E+MxujrQ0Jm3GV5IBT6
33CEwLrnHqsKKXcOoRCCqWclMx9/tyH2MxmzdjwzWs9oSxH2v4VPn/SSBPPwcIII
oPQVKLWcCjjeKvLg5orjkoIOTuDX5p7+2eH8tWe/07Kh7SdYvUDvUWbVh/OMxlyr
K5jawxZIhU/4WqdhiSF0eP9GtGV2+C9c6+TsaXfF3HsJZavaFIz3Unt/ZVRzt8i+
Wv4bdeUa7lpwJS5zcUcXefQ+F3anI06809Wvf9XG1raJYfeJJwiQtRfkYMN3Q9RU
a6pDCBwF09dUjfUVI+V2/klPc02aUszGb8zAhYa0taZeCVGHkAhf9/YOh/R9+glm
kn5glkXrtrOIObKoPGWdQXJ8nBnCur9r1fUlyj3JA6Bn6lWBh8hluXNqSWOc6ML2
5JHZLUmDO19rkVGy/FeVeXuB1guoxDDHERLrPaOBwF3msm8eBq9TGYo9Pl6B1Hld
a44CLF8WY9L25yZpUIrcni2gGg/RDiZtlGlPiiwY+i0ClgYt7AecO3b0y0W5XIsv
h8ucUIIhKt6oREXzYjEmbprfxzXAdTGeZzR5HtAi56eSvQm1KpsUcDHx3YOKlztI
u4mNRzqsWnJxIMcToV5IaOi0Amp9TRU8fQP8EEn0BIC37ZfHSaOC7QEly6NcXjk0
sGxeORP20hfOWZfFm9UkEzatR1eJu0WTWT2VncmWvNkNIXu7ce7GMCOBL7WYeh5G
VeJM1bjFAtozGVeO6DGLoRu5Hja2W4jbSaxhT2IsAZcdA9ONE9CFLpVaJo1+8koz
KWuKzOn3aUr9ooyCohuzzeNnBCzu12cfubKCGMQ2uJrjMs5OhdIx9IPEx113iYHj
jO4rgV1x/E/1TQ18dw2rjJsAI/VfzWrqJcpyTBCUwKpelYC1gWw+8HswnTnNHc//
I/8UJhg078Dd6wAAUPEy1A4FjuKSDi59+inO6V0h7fcxL7Q394+RxqOZJ35qHs9z
SQvfHv0JyojrCu/o6BLEW9rEDDXwH+p3oT51W4TMItbQmRYcTYCWYjVviUbKDJ6s
PhMmZuIqdrRiLHf9jbNOnvJ2tHY1W8gTgMmloAQutp0/4YEg8ldm0pw9Hw6hQ8//
q0vWyw45AhtbjYPjXgm862bzUoL7aJusCIaKhmBHjy3hVxOYjIwFgcO9gbXD/3Bg
NU5rN+54YeGFjnq4R2l2f8aydHz580L40XnmVYfJlRc4RLJq5LskcsUfkzRUazWF
LsOMJ3dcIZqSjlMxMUKkb4UBJW3CYGwaaSmAgfwIr7K40hKGNAepw4NGqZZxO2v7
jPNSMFaZqwyjMa2b0XqfmbR26End1+I+mqi3cq/9FYpKDg/d9B2keGFufDWY6t7T
OkbOI851gGxchfeNqb9XZ9PmKd+SSXoJu81O0kaR6BsNKSs5NQe11KP8Ow3G2dY+
hWIl6roi4hpJBgLkpb/rZbjneZo7axR7lMWyuDb68NqXGChON6sj5Dw/H0ceurTo
7MdeDCqAMQracjX1muzGmF55f4J/Z+VuyiWDwE5l43txnNCV7x69IydqmeBCgnPk
LYRErFfLcitvuVqAOuTVVyR+h9++cQfPWxwrNeen7h717MRuS/iR4D9kAEyDI1hR
OMXZJuaVvBNbGVSv7tfWSIEzQKijEGNM/Q86CM+t6SBVJqSK7Z+bmxm+uNyYle52
qeJMEuHrPw/z/1wFZFbucYj0yCuDM0gUIbMAVS820mHlgSY0rfdSBDbjisWOa9ly
ivMf8mDCc6PmEZG3RdGmuXfXmUhLV3Tu1RHv52zAqPSyRV6YwEcG1jJYcSYHNh1m
4Dy1r6byNZbalwc+tD59S9DSTRjpnWy0Am0kdwlT98rakenturaDAzpuqilNeP5a
kICD47RfZTA4StseDeMQtO52kIuD0GTT6Iy75k7MowoOFlTz0eb04kB0IDz4MAfC
2sTb8tUM1IoOHYgWemcJCl3weSaXYQrOZJXbHRyNXcL103Ag6wfEGUMlPFFSDjO3
PJRb/37c8U4ZYrrqrOiRrLimeM4ma0Y8jUr9yz4qKNRqM94TcDL3+xERxtZUNZ4e
unoBMerfzQpgmA8apqrsumYCh7bU2DWLgUKYwcF8Bppi5C4DGO45e/LglnX7U/yQ
Jsi+fk9JhZTSiC/ReLsmdzO4f5j7ipb3AeFf66qyCPII7MB5g43HQrrlCzMZsxQu
b1k2mRuhrn4HjdPr7jcnmqm4qEYMLLS9fDLr7meizn32WT1sBxeBwiPSDCLvc0tK
nCdzdx85BJkA6DHpnQDqmGjcDCNRxtYKvIgQMvGVek7nmhU4n3U+oohao3F6S0uw
faDLZd+KNqS1ETo5LtJuQDaziU606rOt05EK6qkc4AV7O2zD6rfj/6K0TUOSeQ4v
rNC8HjjtRlPQCpTkAddCq4XXn+trRYRh/QYBPhg1s/aG2Qj6qxPBJ775gNdILw/m
cD47f104T8uOqgZ3w3b3JWOFCrCLSgGp79g+qAafL1H2Jiuggcq2UCMhbFTdUxgW
3vF0efFl+T7M1gIRzloG6GuoIG0O6rfF7VK6czIoyGw/1CADQO/l/o6FwV/lXPA3
vmnnlnEXSTsI/KvW6TcTOvVCTRVwgurW0ElKt3nv1nUC1dG8uqIy8hpJRchs71+L
rK23qtdfmyQYkpGmbn7WDI/VE5qwv9vInl2CqJAdE/1EbzZuK0CObcTBxnCQPEDS
bf91wR7vY+1IhJCO1Ha0tcVBeP2WzCAGvFmbFuaTymDapQ9Ygtf0OVRdWemnOaYk
guvQZShh2HJf00TJ4Xb44ObS2s+OSvRUCjXYH7uysn9ikK6e6hS65tpBeP1sLOfI
txyB925C8LJ4kSINCOHjdu+nJyCLTFXAyTK2EqT0Psenb0uGrqCjxvGRMHKEYEou
vimKW2jASdCuQ65dJWvZcbVULNlxKOpxaEPGjp2n/+QVi0vJ2yz5caNlTSCMFD3P
1t4mYDabfcjN8fG8WOJYHMo2pWnlPzweWx6b6OZ1qsjBu+XgocR0TePKkoa6R/9B
cdx1xxPm+hSg4go+BDJ3DT5KE6ZEBifPnrK1PqoL6FaZGXKtpfj7v6Jmz3No7Ekl
xhWl7V18EAOe8mrS3dSYbtwxDZELkPTDyNBKromcZzhbvzupV/pzWOhjYJ1ZZAlX
eLIYGA1DkSETDjnV06QtZZcB5dv3rHWDYxrK0uKUxbiNwxxDfS8QEm6ZQT7F47Fy
iCppeIsU+G2i10bfH8URQUP5j/0d/ZouoWy4YMKP70aMGv/3Ud2CX9EPhs9sTCTj
+Q1cbMudxwgaw9zUXvnxfZ2f98dBWuscaH2oZwJVzFFPY4NCGBAvLc8w/y0ZUrTp
SscmRWwtFJs692f1uj0Ko56bpb/9YRXYO/8+RUc2ajg9Q/izv/O9HQno/vntw8Sg
barxbQ/MWy2VDSHfwSQYW2CaAmw0jn8JED80ve7wpfP26ZoUxXdPZzSIsBLk7zlh
Z9zWbFf4qnQaDYlWJ5k4/Z3rvISNODA3bbb4hy6CXayXwhaW2rqmehWiS44h8jLI
SSW0hiVPxWQKTmx+MZya679pYKDHNtudLBh79vnoPkU4YYRrQWAZVNWSxHygjEf7
OsiJOhIvZP674L+7/qjNaD85N9byqrMgpRqdnKFHa3kTDfm4gx3YydvcmAz0P9im
uRLSh7Udjy8/pe5FqyBBGIY/jvn9ROjGp0QelyzmHQetYy4b2O8G6MqCKuxkWE45
7t0sr8O/4ndMrj/OCsQEJHPi4tpdsJMgPfGmS9ccJoVtMlfuLwRITL47QpkXT1/i
DZ7ud8TjuuHaw1Yhid0bdd5OgnLOOyHh9wwbREBxB+GSLETltDzKmCOjw82qRh2W
cykQGpvcnvtzExe5mM/dJETDe4qWEM+dkm8FzRwTP5Ir2P+eL9cMKbNcbhyQeMBE
pbV3+GzgsvAOB14T8/3OMNlms0jcP3tzWMn3e4B5YPnVSviddOyfqJiTPL6ILUPz
lfDTISC8jkZTwZnrqLOf30HpU8SArnzRwjxlN4j7iRN+RB6l1UE+ybnpzpYmew1p
guWRQVwg4Wbnsf7D+NV7LlkfpH1AqigUKpLLCzVG3utrGYefwyxH9GJb5h8/ADtr
Dv5MHhV52aggTwJux2rqJ21jSxYT4GRp9nMKjTApWLbbgvlfqXTvtuPGqcD5LA3Q
J2fm5BHOD8mnQuVPiKbajpbukP8O0Y6dN+1xS3udyq7MIqXiqoSZZadz0z9pcYOj
ctjLICx13F8ip5sGZEJUYq12sxbHIC9MLWxh5shcTnEbPT27ZdKKLWBvlGtCIK7L
1YgXrKZ2OG2pkBVCtSttRXs7Jg6lH3ChBvjRs5iUueWBkmcnFpWid095ZRxQzFsw
yPhPZJxei+8LV25kPXuE++1cQNTNiedkRJEMKOgvq3k39ksVr2/7ViQCZ7F++CnH
xRo4dh5cCP70NMozJS5Q53NS5kK36otDPPSRirKIYqg90F4zyP9ncHeF8W7uHui4
GM4/0PsWW50w9EiNrCJLk+alL0jH8v2z9hZDpxmZ/uN4OKeOj6hTWdxE6Sdbba23
xzTbZBQ+Eq+du47kB1xtM+BOZi16Om14t+105JPs+hVJJsPTfGnaQnkr1HfFnEOE
BlvObEOzarcRfHW/tPEJEH1J+yrLv8s/mcIcfqQgxwIntRN9QVKV6ukQgp3/jPlk
mJR+qlwKAeyoXF5YsvgyjzMBd7QN1boThC7Fil8i5qHJkwrQzA/zCGHdFPYpeTlK
liX7lhZnKM0PqH1eZ4LTnk6T2ozGyujkiu0Surd7+ce928dz4WvHOAJ2+F28gCfb
BjCoFpF9hl8OblxeuNuTG1Kmr8zLCsgtRepWcof6QxSFgQaOhz7TRCTk2tvUEP71
CRUvoEfN6aXTGRtbuLDd4hvJw319g3F4/kLAU5at89cwC383HoE45T6MdjHK4pof
RNjHqMTtusV6YMaeT63VOCBn57Bncr6V0IqbwWG+EXr5q7ojP64X1jp8Zw2kQf2N
hdUCLOjNx25xdIctDgobClg26A3NgaKgijgCaKoLIROTAOE1pW3nnWMw0VuacCUS
ZTn+Gbk2Eq2EtRllNUeRhDwQXLd0jHvRxIrdStGvON7XmRhcx0A/Ul7kQbTBGwUS
XYeRM2sf+X38oJV1PS7xp+iEdAe2htBTXV2aBr6+KZhRrK0w3bRlWi5LzfksH78K
diiojwHxlwMdbl9qcb3ztFQx4cKreAzBS5IGPiWs2x27r6WjUhs9lnjq90xpfY6A
AfD5sP03jv8olnByRwJBwaZRbyAdjsCst32Iyajw4xaUUTWcoYeqwYN6E9yfsAxP
D7ZhriKks4pKxM95rReShG6Wb6ooghspENn/zaUtfPFfVoyYD0QBl4Md65EgiWkA
pVRIuSPoaXirVcWAcv6+Nds5+z6nIeXEn/lruBFFDElNgRFTSggoTYTOz3GKxTyE
yYzBpYW9ltezDf/+w4Yh/QGKsS+g5TpMhPWvYaFUJAJXhUFTgZ3z8Pb5H7NnLBK0
PiFzD55AmFj3TQNRFxyPCsraooiybLX0DTSowoCb3+YjKv3rLECwMJ81ecNWse59
bTtEk9SSLWidkQyf4zZ0ZlFJ9ipwLzhAGZsF2vUu9wbQg71QxokWVVTmTj9f8QyT
BQlM16wQcPISBWPhN1Si3IKIzkTW4Y9r6QPT2FkYllGBwUHBIpkZnsnx+n/IKtBX
DQpAAPkUWHc32e+f1BTVP5DIYsofaGFth70OatEt/AI5yx6zyglzM0jxEMfw2ShF
Tal2EnJjWX+3wa+m+uScJ0/jNCWN8od5/osEynP1cO1j9SUqC+AKslnqhFA+blO1
7xhJpFBaSitkHp8+aaKciUZr09q5cJHmz+Tw5Vgjq/ZA+Nch7Sug8ju53/dQL649
Erk//fFjMWX7zp/W98zheYjJWvjCeSyDJ+GQWuX6QeDsLOnqdoelkFrNH26pB2eU
0rQ4iwc63RHKY60/8DlwYYX21oop2SnIaYbiA6VI2FPYPmK+FlfF+aJZ0D3dfp29
H1pEmf7FNSj1wusb/QAUPS2jMwidMClwUT4wZdKrT8mnC4766Kqu0oO5Y3Kv0EkP
kg5ZsxuRFVV5V4jWmYVyrMk7CPMswaxPqL+cry3o78j1Gub5VTyB+6eEQd+C1jMf
RE6F3uSjzWNymStREfHZxF/e81xr2puJkkpAmkyGX8sbEYMTa4UABTE2xO/d9UEs
HeKRLMJh+jhHOacpyeIm0vf4n8E2WJt6xN09HxkE6XVraL7THpOJNHOyK3aH40YF
m85Yzxiarb/muSQ56Yz6pcrfg0cJw5s9oAt4PdOsv2r/ARFghvIeM1IThn6cDCB6
+y8da7W99h0ICB4jlVG6b1E9sOFDBsX743Z1fTMXx8m5h9IJHwS/WfLQwgYz2olu
VcrJZyxv0L8Be4Iorng/GScRDPdSiFalzGt9I07vkQGKXOpXJQ9zbXSHHq6qhOfB
35xYxYOdK/nUIPmOhwHdj5/dSFzwHe4kbI9OuWGR3CO9v5lFsGt30sdSsm3cDZhz
/S/Y1N8UF33dWbWMr9SXQ4ZVUdNlvJnLIq7bfakQbopfcH8P2oln0YV/5IeAT7At
5qJwvb6dHWOekN7vz8TSCYd7S1/N50DA+mqxRtQNxLVkUfWZDVoZsLwWhHxW4n/w
ST/THkiaALwxnH7bqYQvKrBr3TuOWtS73Hpk0ZBXBZBYohEPDLf63Vq6nxpNvek4
VWiad8yeTX+7nHV7wA5rt0F0M1yiNgfF2KtcMI+PeIHqhT7sU9O8R/5mUWe+oZ+J
OsQceOhnqt5GWf6K9sVJWAo8J8IFV1LtFgdM+xYB6lOSIyN0IQHbt4O5Fqw7A90e
SsP+iWrWF1VmRjb9Mk9ljMH1jbqU/HYi33+KLsSAgL8RDyp320lPH79XJHQt+0ll
NEpd98GTKq52HkkvzQhqyVXgU5xXNgYQw4VPT4N9e09VdYSIquRUbZVUjYUPdeGy
flNwQWo+OfsseCp8CSOOK6jchlI57oCa6/XwY1tm5bH90MxREEqn3FxAaByvZhSk
MmjYertFSgNfU0QH3c3aVrH6fhUGYi1gdpFBlCyxal02y8LQN77axG6dM+hMNyWr
knZqI3Nuy/5w/H2WAhcAoRBP0kCi+kbOmTxau79A7qdG8F2p9Kwa6ppSDvRIgLBx
yxR0O7G350S/ed1RTf9o/uMj7W+RpNQnbvEHD9u3J1XpGwzr6+1AzyC80FXu/TEd
/D/jS4EypaAS73fEWimGXGc5hQvk1DDFCfCblYMDy7bH65rJIWgsFcZL6JOqT5F0
0kXpVbBPC9xcIJfB+8CsubYlKiekOtEF7U57h7O4C5OO9hXCJx9v95or9SpG37kz
tFw+k5IvdIMBqOk7/ZsHAgT+v73jagBt6FEhcussSyNA7Xf0wZ86lPPXrZcNAYSk
73YH+YXcUEhvtkLYoHT+Y3bNJQoHs4wNDNMrg9tmFxufFMVq/RkMebk8ms9o5UAy
Kim49U44Z0xkGSu4zMqlqt4mFT0nbx0WoTbn7GZdJMjAm8n5ECdvy/IaUDV37Ml+
9yc4Maumiqriy864wPSBTZ3wliNA6HRzxrUEmTxmX4u9aGuy++1ZbynOylxB8uBH
4VsKTeX5B3rTpQZ4xoUGkiiL7FSf5dCqQ4+BfXGIaidLDJ+xQV4ytQRyPvkh6FZ0
n/Humvbao7d/KBk2iZ47B2EyXGMpg3o9Y5Te5ffwtg+89mSkk6FGUS6MNV7JdTr1
nmtKOMj3Hd/mbGM41kWmm9Jx/CFNsVd6rLoOWDNS35basX3Xhw9aR7BFLrPVfMTO
ls6G8hL8482iPnM1JxfZWbAp8sWnNC1mxs+upaflu4O6NrPreDRsNnEOlxPpNwTi
pZ2NytiRamqu01UsuOryrTdOf0IugKMYi9NC50kIDuMXLckwyoG/yPOKdLSSlM52
VrYV5iwHzicwLw0sDq6n+SZac80L+WEnM7msupmssdLpgwxaiNP8TMHegg/YUv0S
VJ4euAcWdl6kdeyeT1hf14HfQTX6/wpVhVqwE70B7Py41rhFzCh1ax+uQ1mXFRBJ
5xarCQwchU3CBGsCE+9Lz8rYunLBoDtaaRd2Cee1UG4kr09+Fvn8pEAjsFwYXg+u
+hvygXnghISDzcqJDh0XJQfk5n/nPmMZmpFMZXmhkVJZG3KgmF5MSSg4/Ambe8rK
Jd7ltkyKArC9xqaRzFuH4bdG9SlXZDyN/WR0X2qWOPgU23KDu6BmZ7bkSim2R/sk
90UQVYBQ3eSrFwqvCYIBkj301jZHl5Syii6gNYj4UrIQ1CQZFQP1pCBop1tNSsmb
s/KZcrvVONWZyOIkmAGKW404mDLqfK43y7yvCNsWSS9AsH7YxwQ114MK/Nt62+E4
Kk2BTkDqxkUO3nMWFo46jK8VIfBrnwjOwmf9Z+RJ0hWAF5mhvs0H0suFJA70n8i3
udBDa9+W6KaWil8bwDBSkvX+NoYDvq8bYs6t7WbQlLjIdNentbaxUtWF+EeF0V2s
pqaTIzz+NdtnJxLzJmONxuKv8dnIwsC0LSlEihujm6w/T6TdpOR8PphN5OZR395A
LRcD3tqk2f2yE5DhUSHovd80YTlvEra6fKZoMain0rXvwMoq+tclqmkGDBxmRtOr
MDCgMv+i/EEGbzJhrilrJmx4iVrnnyRpXu3qFYypCrP8JrxYKit62q3uut+DdBRm
Q/EkeFCiW9K1fjikWV/+q1S6mX6iw/8tTaDes2Wv4CKEv7NsP/GH2jlzo+uFmsbe
NQmBrhQ/QHPZvi3Bpyl988pd7NsQdzbrV9LMgUpOsbOQhN3rFSE80DVgHMrmS+wT
/kFFxqJFJkTVSf9YAVcB/Ce9yX5lutrU3rQBriPOKl2TmKND7BJQRyRtkZrGPzt8
mUXbKioRL1WJN+XeIkCGiPfpy+lN1RkuItgm6cxm6Ejz94rnahpRkaNx/Q5ale0q
vDNPeBXOpHRCTLCOwRpkwfTUUnjTt+c9M+jovsjdO2qRPsiZl7zZ2OJ7eYfgAdre
bpCapNGW89LsgT0KUVOxlt2W3hoBMtKjSkMULTvXe7w1xJaWlhXcNU6ZOQ/T0G1l
Kpcue1beDlGgX37uvbzIW7PfzA6RzdOdp9f+ssfgpIvE1Uh93ew3lj/JV0pyOGL5
XUb4tuDfRE+gxuWYOz8OtH8CJq52QGOF02FjQoqaoOiZFUcbPxKKh3MfIBlRweqO
EqAiKO+OZCYCyg8J+f+EmNabnD9mMZsyy1WkditbyiFPjln9kJ+xFXuHB2vimN8T
fHzQqLdREdZetlVe0kDHLbKRk+e9m+hHLepvaBW7AMrWXfCCPeAWd7U1gjwuXtmh
tt9Q6H6xMOb8Bx9i0dKLIQRzuD1+Jn5/qyXfx5YfF5w4783ENdulpSpbgIl4SQP2
ice7+OZJPw5g71MjGP0FRtsmyG7CXcgOFoD5G7+JF5VYjgap7zeACuGoBOcVvPz5
7WF0BssvRi40wo+/5v51poKCPMinJwTiceOhqHarQV2cxPPZu3dZis+Vncgg9X4u
BKJLDpmkhLegRCIHSQyOUD6iQzxxXx3jfmNX2Xr3cLegyUUay9PwNQNU57231YNm
LPa9+UMpQ5eRTDbtw88ubyyVKE6oko2haO8gAG+gOk9iFMkQqZ6i7C9+q+08jACs
1M4mx10Ji63WQiWMoGYJ8PZ206vDiyP7oZPgFS7jV3tSoBEdYgBK+HXGEvP6BPIi
yigHAaHy91Rtw6OPE3zvEKWlieVTbd6HWTqwiCq+aWGd5/bac3p6jkpC87pl7lyR
oVB9yzn/EhGipv0xGGcjultBKEOKR/0wM/+ZheqJUSUNWB9IhDluzPr6PIDgQ0au
PeUNdoUE8Vj3Sy517TDZSulcvtLmxEgxFwY9qUHxDIDKF0f8ytyBV1ZEX8ulFGyg
5y+jg/dsHEjgSU6/loFhoyxvcp8yBT946C7u40G2lAGMZIbZt/rIHsf/e+4pBeQz
UyIOk7VHIW3pNUX/Vfc8haOHiatFr0ue/pODEXggx+tJxCU9S086SQItLNP4EADa
yKarM16Bm02HF2/O6fbEr2mwhYl5xR75ZvQqmu1VXqqtGtBaTrQsSZk1EB0uqmkT
Kceu3UAwRifkkjlHBNlXe5oRhXhX+xCn7l3oPqx8XLJhugcYAfdDBSqYMBgnYM+E
KTnKji5WaeEOuxBjF/Wjo3ZD8fLVRjDhpK6GBKhOUeT+E7APwkBojbJI/ikJ4VPb
j1KiAEt3a5YaHCiDS0whmchsonKxqQ1ItHIn+inElkWBlYuNYd3GFlLs7aa0rQjz
dPiWiZwVUhLaf8KtUQmm0Bl//RR5ClL+L/AedVGJKeREKV7lipDO1zF0Ppvfi3rj
j25n5ywbrKepUc2l5BRX9B1yfLe9hMUXA01aHxqxQKzlCvZPXCGP22k/JHRze1DT
53pwRs+NuvsW2IupD7bPglfiHbxbRbuYFZk0rFYEw9FkZngd5At+HBYerRPs8I72
WK8owpUAuyVpTa5aJeoteYqv/VeG153KI+sZ82qm4pl0oWQ5A7QLjeWvP95+5Gcl
kowVtZ+SxgMDF0s5spClXgaiF6b3IqE3lCwotdsRd+vUrsX97eGwMnoqdaqIbyAo
iLNQzO0GxGb0sgC56u+/kk1JA6NbD/M82hhlewI4jMx3kfDPl7W+h6hNYYTAn/Jy
7+Sr8TEnfzqqIBhkiKOQx6ZEwrqzSslM3iOZLXnohSOIqCjtNrQi98qksZpyWyVM
O1itcMR0KB7wjFWu/qQrWM24avAkgUgyVNduICLGnN8E2Ydm4Ztg6KCinuJWJ95h
d5BLScjRp9E5kO0axtFUd4Wyg/jzNxPfWdE+VptW28bookdqHmgfXGWULUyGjKIB
YRkWnQOwXAuCgk+LNIih5MEav8KDKwD6cDNlpysifn16oL77CLG1mefcgyKTh13H
Zf66ccBCZQYhJ5oMIbX7rUezWlhpOKSCDljPbBphg1bCdSV4b6l2ndvUJ51pFNaO
ngQSZM0+s/67Rx7MoQfjItwpLIB+9GuDrPY0kiygHpkFDZmYV4MNd0C2JLFCiHW4
4sBjAq/ImjgPk4Was8yWa5gGyf2fpRd7exLwyn9n6Yoip2d4xeK/AqGkHu8Zfg/K
0Lxbt3DU7pSD9Wx1DfWmbNhF69Sqk+Qw97ObUL+hIetPp4Zb/mmf2FCHM+RlQgRB
a9VELRuGWu6IShFQSBND4XWEO6V8NqRRtO/UiQWUFpAEo704BYvFOPTSz5oEVckr
Ri0mdJvr4T21vPN9bGsNs3xXKSiDtZI72UiiwTPt9TiAKqzUxPPqG0fuogLN7flF
MNHnpW/DbELGjkag09Wc6zjUBAmC7YNq3KIuKExV9Hg11cW9tFZn8HXqC503hooG
S1AMOtChFgVdgcp6biR/Ky6KPGNCJk/UaaG6HHNaam8S8TnuxuQY967JUmShvK42
H0BkSei2Y/YSaZLCmvLOxYBa3xKSqhqE55CDaVEv73XY8bPm28SA0C5/ic7VMNgE
udk+ccAb4BkEj1I+aPb4CGjst8CDzx6JbOigJnEur8pIb5v6+kc1v4Zfj4eBQo/K
eX5GFIGk5ty9x7x3u3MJw+lyd93LZeAMvK7Fx6OS8wErX4nF+4MfzIy/1HmWzZ0/
4tVWN5/mZvJsblb2NEJFHBssHodsP51b+dXkbRhYv2ZCUcoskPC38mDNfGt66ap8
NHlsBVVRoGUe/4A7ExzOUJZpj+MYw/WqCOR8zJRuKJtQLe13OXv6Ha8a4jhpGlVW
nh+UwAQNigFNvOuIUD6fpynQumEkLyXL5mZ5riPa8e+4duwQhDHbNHqIECffYGfP
O6yxuR1pkG2VdEHQkaRIE6fDB9fLjqnFN6pvm7HQxaJWo5C+yhs1wjrqK9rFYnG7
mW6pMrTOdC1LWqjweY1bXsttl6Zw0TbEjiFyhA2cVAepL88rZmeTbUccLtocI6wA
jO52U/Kslt8vQWQ/1gckyr1z1O89On7lPIp3q3bU88ggoWcRO8pfEFPzf3stY3nO
bZkLlyDYhcCHaSPmt7I8mnaThzs4i/vrrh9kaeeZyyxIwSaSoN0QPS5Ih/GfsCBL
JTV3EIylWQj/4I2KBwJNGOmqvyvRPLGoGY7Eh8DAuulOsFu6s760aFl6cnEWBc4g
HOEjtHE6eqXSVeEmNt5jVvJmkioPwX72O8igo/rd6pbZrihshAqL/qX7JeJHj/GH
50fT5LbV2Sik9WpH2CPXlOijRM0YQg7O6G++76qP2/0CcRdJx8DTbjS9Qik6ghj3
lzRMp8Oe82jUV4cFbqiSsNskm7Obz7LByLnM7ygCL0ZQ5tz9Bnl5L0adjwVomBnp
tzzf8Z0/kDGiGEpNG5M35sT5hN8Kn3D6tIdumBJxnBnwbGLxcgKf1ZqFEwGgYkO+
JFckONDsfdTJVGgEa5bCneD6VeWnqVHeD9/TwHfVSNiQoyTBrYU1G+7IHEFzoO1u
rZMz6+6Hbgf8iNT4a676+Tuv5CDjwQkiB+b5EYEZxSPP+Uzvt2rncCvWEvViZ3XV
r2YZokC5SMX0pdvtGBzoMWvRJOkomubpuCGhq5ZezLmyoH0Qa59EnP316kK0XBXS
SgNsW3qnAF6TnaikWEexzK7sMOp25fjLYspdYuQoSD4s5BAhqF2ud82MGdTjNmO7
3I15B+ggGcjL/vkgsq12k4H22tnJaShUmwpZFciaV9wKk8y4RyP2x1WCzAk5EAZv
0vqwJ8DZYH5/TkfW6MejINn1aoX/rDcSv82UpzTNiuMbVmax2jVG/3S806r1P8mo
tVwIqrDE7fsPkhl+WHNPQ5Y1CqahAG66BOUlxFUIIMNLNLAhEaAhykAtIkseHllp
RF6KnI8app376cJbnVh+kLww+fR1z1dB1UBCA6WT1FMCk5dGMdEJkNafNSIm21YZ
ja3OvIL6f9/PW8/X9XaC4vqAK+pwEHEilpuNrlZlCqN4fsm6OAoZ004boHwqF6e3
7OR80pO2xollEpsAqHa3uSn5gqCVK3kYO4iCGZQPFvRWVbQ4ujyvgLmmt4fcrNyk
+iJ+ID/6jcDhZ/wyg/Y+/t58Fy0pONnlgRdyj3H6HEaHOByyUuLv0fQbBFQEzNjx
KqtaG61GGqmQC839iBFbTBISP2mx9CPOF6dAQP2gfGrJf9UJmUmkl2/thYcb4ax9
9hKs+/m6gUjkuya4+nc81PBu6xw6zmE8D5cCkSePTUqt4ZOrvD2yRpr8wLo8G/kW
pHKvItBaQimSN5Ussxk+45LNkSjUSvd3FVOUf+xw8p8PUqkdSmQzco4qPVqbxRj5
Rehl48RT46JMKDOHLoDkV8r8msep47WWLIjv2zbmUJKdrSIvFeqc3zEswFrwhiWO
RrX3KUq8QKQI6DhvYnm4rFmqYpHDGT4jJCZ9K/ZWDrpNiI+Vy1H1ZwE1noO63Lt/
isrlawR4UaPY230VMW0j08XS988wSPMfW0VaPOird1YUUFo4IoAvsW1Tjp8N/38M
cCnRnjz2eABFy2iycv6VkaCYyOjQ+15aWXZUqwsmpLDaHdGREFnU4i77kbgDEHqZ
4QpLhzxhibr747ef8rl4l3m8YNhKdOmivK90ZPy2mq2vfGX8hl39t9S2AAz8gmHc
dFKgqLgfm+6xWO3YDj+WUe599hYBt8xjqpd4pnCgWgc1aJeu0/BToYaOLotDAO+f
M6gcJpuOKbQxN/TokowuYMlJHVZ3Gk6pWrHPBmPGzh+M68qrOcPTy9Gwpuok86rE
Jjn+BMhaHO/5WXfbNaV37a0dJTFPy22m6oatT353A+LknmaQP4o7t8r3530gUbxV
g0ML97+cZw2aPOkVFbM/+1V2CfzUwAym8QKiIkswtvd/eFK1hYOsG81bJB0mOPV0
uvd5LHE2tAXqC/PSvwnlMslVEjXJZ6K07OihA8eDi2lf0Tbnh5opWnQf3olro8r7
iWPP5zpCUiSjPvJjV6Dktc8tRTJJZ9+FTHlQSjGMXx7Fqw1E5mNnipQhOZaIw8MO
/dxMkgq1ht135Zu6pPnhZT7F5HwMJmSNTxAGGw35vUQsec/+VgX/iIjPNlQR8+C1
q2hjwWli8tKdi9Qv484jWV5L/Lxrhx0QaH1jfW+UjsrOAqk8rLCJlWGloOPIvkJL
XLUY9Kv50BLrGRP42TuGDYCevy+3niPdLRd2UEfE6zIEZjVUDu2nVntcYx6sv1Mm
8tKA3Rw5dnrA0Jse4e9tlAerDHtG8LoecDKa4JHli1NfdojAXmnYoTqI1QwNxDhd
BsTCm4hOREYZLkOOAouN3cK0+95f9o/C0AA+NwwiMcNT+mrrIWoq5OJmjQAHoMCE
2v4/LVwP4kyO3Khtk8gIioMUGJRH0AKL+/p9vz4IX2zxxAMIiv/UsW+3TOJ1nlh4
xHKdgq996ppUl4uyI1E3GGkRxFg2INxpYcHTPup/Wwpw7/Im6qI4cDX8v0v3+bZG
fcmWDNkyXUV0Z8VJ0GpzMzRin5rL53ONwqzIuFLofjyRzyXRooiK87tg3leg5G4Z
ZXU3kiHB/yD3fwMOesrPP7ZPk/lvss76thIzoTGHDAks/bdYlzbB7d/2HQuyE16d
WM+Hari3k+xx7xwFnl17rWJrZKIzRItODjg/AkvAmWq+IKNY4sfICrZDdkvmQaHh
XV790EJvq1YVcUz7hLuMKLsf0UqECGKxKX2aCmPvkOkFDX0kt9N3/VkFKMXrUxJ2
zcEEPx9yOWT+etBSkYDGNG+flFj3w5RPPyVkh8d58vIl9HHXPZxqmS03aMgdnRQa
K//tXviYIDKpRecCUh1UA42r7g6Dl2WUeiX9pkj6yldhPEnWoIP1YTiD4wTtzx0Q
zLHKD54iebO3CbQJU9wB9vtemXBWybHu/AYo3murzzIU0qHtt9hW9wc6uMYEwRVH
aXxM0sAO5/L32gM0GrQ3XbBPyssdnECkvFDjSpP1uwyGmSWm6hs0etfwPwKku6mR
yAzXYUnVePL7SAQ9Kp2Pk9CSVpk55XqTOOfLUBU3kXxZxJyQEwGvmatABqm+IJZK
Rg2eCq2F3Ed9P5I7bPIL4RVyDgEpHtORWIJklE3ucRitDt0+sonsHVcIIl1CO+im
zei8pmIUWhWCKEGQNJKvoqdF+Jw8naWu9gDFN7Pkm3dP/YwuCor7Akk3dTmNlbO6
ltiMzNNuqtlGtLaY+z3TEoOr+icxaGDxuBwLNoJzBEIUGVulhs6EexGHBsSW4+5K
GlWbISiaqS06++hrUhX+jvwfG1UpqlCc8Sl9UXMdbsP9wMUhf1EnemqwN8LvjM40
zvgeoja0pdnHxSiLGK8wqm03cgsbkgWJu7KYZfHByhXJLSQMNBVOkG82Njb3Yzgq
9DKLxqIiV2B4Nlhy7qEMgC/tWMtmltsnTay7NNDoVTXfEr2KXSL3UaLk0AquCYPZ
T1FmvaUCPeRdJGX6mIAOU5/si8bWi5qNzWCcCSrOQqkOiAHUkF/J5KSmX0WVPLT5
lAa0AXTdg8VC2suOCeBuYq+CDVT+tcUoxg3iGbA+QNDbSII8X9j7COr8b3zGLqRH
d/Oaoiar3o48nCJIxMKdJ6CP8BqX1XVV1WyjDw4zrhrEOAvFdH55UsHXEGZkQ0zX
yAMlqn6YU9F2JC1S9xLkDDbobNn7jmhLDiR+m+tjsfQSkjV1pq66X3bedgtxKoyr
5P6RWPkTjUOU3OYF2G0eBSHcO4P7Y/8Bi8dD5N1Uwvjkbadcs8r/OTmWsgU+ilCl
TVdzsGdhle7cDkHZM/tm8xMB4nnQp9zOWExxIfdDR5odKntFIxNQBNReA98RSK24
F379XmQGby0GwU7NbD0ZX72Za0CZTxP0G5g0xjDc3UBQfHxR70/sZvfRY3MYmn1Y
5KjzZ0Z8DYw/i+bbrMYOn/2uNPBk9PlsCA82cPGpX59tMMz94XZbh5m1NGF/hoFv
CwxBtwUAlS0/HaBJBfd07S70l1p98Sb44aPLu39LjyCkdLCDa5AqHtz9D2DyEJEn
sM9tQeOWk0tihv5aENmE+N4EL5B7bpcvXaugngwgMkMyOuumJPUwFkEpiKtsSIUw
1P2Bbwru/0ZIrzLVEH1LraA3pWunJpYOsW4KzdqkVpWveVkPqWrDvWk5+xzrFTIo
TPQRcFmn/V8fJTYDb2iafXH5P5A4dyY73OvtZz8uMqQHvhOWhMG9WkUkmYCBZX5T
W2J2GUm5tn3LaW+7WkRGLrh3upZauH6cstfPcmezJwm6LtI+6UYHDOHd54ZBQbrO
o0wz6sR5QiWbkSPf2o5RIIv3R/brGPq8y0LE/KCmALHlCs9L0qIE6XSTXzXJcBJE
UqsXYsM307Pd3K6uD4tVopAHZo6B9movZG/W/P1axfaNoe9N0TeaaaSVZaWo02wS
oyC6yScY10sjxg8g4sRm/ZnKuzF9/MsEKATbf9Xz1PzkoE2k/9avAGyaV+uSbD4s
8Jb8jD8gf0hAjKxnsE2V3BmonH5UGpkDNM7HhjldDdSYjax74v3P0g0tGilxUa5n
H27tIPmJsg1ilfptCSq+qEJmMrNuxDk7J936nyq95NDgDspeB31A+JKbBklUwkrQ
/9g4SGXyRSl+W/frKwK+maiJmUb2CAh9Oaw0DIOQkWQyk8RcMOydT9GITb5Tb9rD
yHgSBo/W38BE8cG8h5pt/u9bkH5Ej1CtrF73aPV320u5HZC9DeS9FuBAcdIBMBbw
sILEH8dHC4JS5Y9cOKOy72v+z2JG21xOvJKQBlUhxdUxcd+uH7zCCCeKEZyd+LTv
o9HC6IoBc90bwK4rEFA3wel8/MJbseEkYOjaNaQVVppZZzmtZPfI8Zw0wMpUf2D6
PChgCQkqyOnWnk/Du5Txupn0rV1uf/7a9kVrEreoaSEzNMDpxaKwYDt5KHnVhcrz
uj6iE6yRXTSLlVGacayU/MoYi7n39x8nuWk2OB2D5pnQEC8M6mVPUEV5aSGYz0hb
9bXmUik9C87v5Qsj4hLDluFxUySaHSuwTqIu4SQQOBu26hR0uPvbvEUN7wL4hBuW
FiL7QG5bfggEFRcI7CdLCICI50TpHctWN4g2/TT2NGolH+fILUx92Oi2GvxH+2EB
T077OINRsnvQK/kTQmN5nufADUxKzNjT2KMQQah9b+woCjc234DrjIIGoQ8O1XI3
pGYdCmezY77KG+vCBZ5PUc+YdrPBem+qOgU6grJRaIo2BQtmGZz7nxV4lzLK35Pf
ordJCDVPBZkBdhgfKsvQmR039XLyye78hDlML3uLhhA67N/Z9Kb99AfFa0n6Jm42
Eergq0HVc5xMLr8dH2VizFaC3X5HU3N9zukEjDYcSeFcKrLJvxa6+zge265fEbvm
l0dIX9UjapQV7BMKNJdghvrT9ugx/9uSqnLSnFogHMQVhx/THJpAnghFPvuyX2QH
+UqffgcoxDYNLRsGqQ9uy4vWXKBIFMZmxeGX5KXKkeL2oMQ3nkxjcvehcDNUKdTY
BUZiCdOi3jeqY5HaASjkH4EXbJxYHWn2HZK3Ale+7P4r5jjMtszXYge9nddPmN8C
Ianl+c7IlAysmyUbULxdvMa7s705Ny5ola2bdMrz+oUN0yM3+W1OnsacdDHK5bS8
34EiQbGxueqv1BnwbONDy3wi7Fs3aVdLrszvaC4/XUjh1tfC44BgptZdksp2i9d0
7PopPTGJiBhYKH7jLF5G8wuD+gWl8E/vvUPdKNM1CRUwzwNIOoJHxIvtbKdbSjaV
xYExMeH1JUfx4KaXOGhskkUICHLMCIv0s+lY0eEJrnSMsbuyFK9maWCxg2b7OTqT
p47Ir96nZplWACR/Krc6ieEUoiqIwdgjQe7cvye57YYu7BBjOTeexpTKJLjOLfJz
EuC9Fz2KJOXURKscvn1hzanRnTmBpfofWMTD573w2f29BbcFpEWJsmhHZNoPa+oO
bnsl+4zakhioysN4B0FqVLXu6uRTYArPT5S1a0JipDxm6c0nmGw6HWTJaPtchnvF
3Q3SQniJOIDvYZh3jQTzmYEvzgVYcl+5ZnGt+YWp9RavonWSwqB2+2UiWtx1b/Ai
QLr7YKYa2KZgekh0vomySTU2gXcI3WQsIuuGVH7buiqhCAroU8m/cay4KHvEv/VL
Rs1z0ETd/BZ5s8R1OLvwi817YliPDNN0p6cY8xwDCWpcykjP8Mna7wOCG8vhSh57
gJMf7aLZEC8sTQ+uTF1hJdAUnj9CwqqVjBfNBocCYp3mMzv274D1qTdDNn/mLLLP
76wTH2s8qaeIi631TrbJYKzKbTTezEA4pjLsJVO5Uu/SfgGAoCBmSJMunERLB1Vj
sRCUCQDk0F6ETdTHjsCD7xfTEw/QDCPuEbWO7TnSV7Fx0E3gORqks9tLR2nPdmgW
I4orClxmmVHWNNzHareJ/YXL9c13y+42dbtlin38LEfVwlxaR1/oFDJCynL/6eTx
Ml7gCQek3EyHndrF6oGxbsH6eJqGQ2FaxfcNaJ36WLhDdEwvXbZmZCpo+kppEkcD
6uy7bkrNAEFnjPUkUDz+sYA9ARdHTDmxkL/sTl8V1uGGEk01qR2oIlxkfxH2QlQk
qYY7AgBBNz2gRTH/s9Dhx98rDXonjRJhc3SXcZF5x8jJUXVWlvFPYI3lTSlszuo2
vvjYWuCTPXsDFI7XZPbTRLAWgzsQox2Wi93ZPDtyLCzkfxZgLX5mLwu+eRcFQeWd
8vikTsGiBQJg53ypscq1mdZHpEaTCyqUu0lq2BCz9ungQft3pVDyDZ5Z5s25+cuy
oqACk/4DAFHXeMZOjtm9QwCMr/Z7xMdTyB9ixFiat9ykYdCzzs6gy1Zo1ct081Zr
R+GaQ3PlxpFt9wnr9Lr5kF925i5PrbPNN4ymAnaGsGe9BOL4y+91QXAhR8Z8YzFV
TmGH8hPm+aPZ01ypYz3yPRWc0CQge9BhTBgeWIDQEG66k86UtyyFZDI8WYgTnXpz
i1u8UiOuFmIQ9lP2Wsvk+e7ZQXP31+TFirXyCw+vllINgsAmkpshWRgcSpmyPbcM
KygoXHFU4baOP1L5V7+MwCR9UEIvV3Hz4KBLsf4d4GDL3zYYXfU7vt7o9KoJeDDm
+8n6RAHwGOazlg6eVWoDIvrDWx55e5Rle/D2x8HP+Pe3XP2kGg8ltVupquagJTUx
i1Q6zLgHltfo9HULuK2NVHO0W1BifthLlPpyZnKUMjeqQFdgPJdbHeNAY+bCqo4J
pTNCCTzfV/fs3fr8XoJKmOv7fbmRyph+MpfbL3K37kcsaqhi3/+a7Q/qOm6WuSS2
HOfSFMHQxh/g1SjbwKnObFk7ptuuONeQiWg2grynxBAAi/7z3Z6Z1B37xWyrr9Uo
PBxyXBekcMbOca/v/J9CYiKSIG6yMFcbm09kfqAzRrEQ0ob4QV6MFPE7joTBVwTr
tXdSNXLFTSKBWIopYUdn6vqR0SU83vVwBMDqfSxdNtnIBMVqZysw742Y1dGEwwT3
49j+Lli2JXK6qj4zD9MTqIKnq4jt72lYy1P4j8hn3ohHsdD7hRWP6OUFL/ypEQDP
ord5eNXpBs6mZYaFX1Ug6ce3t0NVxLKcQyYfsPyctlKxuJY3w0QarAadPGjlzU+U
DAFnCI9Kg5dPcwfpV3Y4WzuOOkws9nEfvHYmbFNmuGrC38VZ3FKANpB241QKybuY
kUU92o9bquyk3aWCXGav/nn0hqCRTriUUdXCmZP/FPThoQEkRH8vaPJAkbVspG9n
3T9oYlGBi9PxIuvWLPPYE1uxl4whOpIQmBCO/4U3zPkIWzgIDzkWCiPUMsrsJj+9
wtQpzudUvYsY1xrVK1hr+GXONza7g+4isB8g3vNzDCHpv7NmmVxqNVJuiAeBv4LR
MjrNQJAB8zqi8a93coSnZnXcwUgbXmc7EiXw0Wo+xxSKOrpapIEDXKgavo1S1X7j
9yW+CJ73dfcrgDsHnxj11nEUCgcw0We2822IJjq6urnyKsphgS/Nlj/rOxuQ+S5x
oP3R5WRMFZ7BX+s3DbWr+WeOrG2LngZr7suhjck1IHvy6SatDHo47F2euLISRRsr
hmr2KxVIDn+3aJWHERUeAOS7b4xnxQusjHI5liyF6v8sSYU0QA5gv00yG4tY6iu3
6sXx0w6+hpkeRaqzzyWITJEvCFXjcupfawh9k25MLK8CV+CnjFCVWxrikQpsXti6
iULHH+cpGUhPde76xfS3oz5wUp2YZ2EC8gkoHB23rx/OSxOBmHlpf9NOZeZnmGHn
+3E4x6yE94hqbVWYgzF6xhhpqBpANSo0Laku9UJKY/MN5HwYVdbSo+7zebSemQxC
bCAdMa1UcVgyTlJIzRCAO1hdepSJ8bEMVHF7KZJYnJIqeq/MBYE53GtveyXALoTV
2GtfmAWYU8px6yj9YQQfEj5o5x10kBnRJnmxkRNjl49YRqgdZFUtpXYpEtb0IU53
25VitXczheAwaAutHd09DmP1hzVw58Wb8trUeUntS/g+qy1Ds93PvqxFU+LvS4gX
/daw3z6V9t3TpPtuVKhZLWdwP4XXq9mVig18V0UNyvEVTtd3tDeUFLFh8RF/gRAz
SI93d9Lf6Uxx+6o1e8mE5NL6sF21ZQ9CypemJrwl4kolCcOzgSednAmvM5udp3QN
fCOi3B+9qybAQ1lbxzxeJ/bcps/ywmIdodh2CkiQToznbhVm9OI7UTMRIqG7HGlL
PoLyJOPURhJtW2MkColoy1XtqeFkbSC5hshhcJIk00rfHw7VfesdQVTlQH/QLiwN
dIKFHxVF2SsoyDiniyY1+F53dxRs6R/rs2rW9NxnIunWcNcubU04u4vO5wVvu2Qf
RmClXWHe7hb8X9QvFzGZO9Oj2h5H5KEaZzSFGsPwh5VKVxxKA2nk9Nbib2tPj6Ri
zOdZ5Orj7CHbNJobn+/saDzgdy5zlpyOvEN3UOVQkxF/GXqy92dDbJWmaF49bqXd
GGx3kSj3236GHiFbqNyYotpijlDzgz0IfSKbJcYKddXLGrB7b75VNawIdE0RGaJA
o2bSm7DXXwC2Za38k/LSc4xtMfTTW3vIShGstewfuYqqXWUxrWFMphnOVkcSSGwo
AuWu/4ijVO9oVXQDcSmx5JdvQ53PsBQcRljFZIQoZYDEOmtiNMdPM7MHWdyL4LkL
TrrceUlQTLfuSURcSQcS4YHHRBd2K5ze9oAxpvFnKdV7d8cj70y/PaYB8nkW0pRC
1FSNbf0WL5JKa0mFcAbJz9thtYTqsLKNRYCZOQzrx12xnJkq+MSqd5WGLA0U+fd0
YqI7/zJBhX7Nx2y0RDubUcriGB1s+aCSOHMNnwppz1C0MhTX9/3LSPp15DghcLG0
2jfiqBbbGOo/tt5Q514/VHnj6gZPHPhByoQXTSRqyC5hYPkOvQTI30paH25oNgDH
xyp26ibhRurV5/9xbCWgRIUTJhTaj0F+VglqOO01f0elPsMrY5u3kSwuMABy4bQM
40EqPpweFhEU8TBu+7cjKz3A0oJaJYztVUsax1L7IwskzOX7W4Us0R18MGNBAPTs
ucuL6mIfxBpkM0QOyTRuCIDRtXcWq6fz3dw2FagpB1SIL6bK7SSjKvRGmK8FQlNy
5L7XseE7qG13qVWZq6RPFe1pa521R3U7DF89h3zQ6Gsl856fR+Gh/kEDvkP1JbNH
EnH5lHrR299Bt+OuUmrLI3onTmiebwk77Kat5TTimVQH5diNqEW8Pe3qonLg01Sk
Btb3E1Lwb8O3c6yIpTns7z2sqBQP76G0LuN1VsEyMMYT1cjE+O6A2CmtTojxYDF/
g86N5IRd14zwShZRS7OIyICk5g3JNxFqVEihKEVbXX8k9VVRJ81VfTUE3EyyIUlH
E4tmd24E3dDXj3hGD3nWxF5tg3H/8pMmzkRB3fkzArB2VJQynq4A0ESLOaTP3gXT
c9I9VK0wOjDPoXmsqbBU8mXe4wuX+VUwdNZK7Q1NpinOQQemBaJyq+dOTnt52R3F
cIr3LvLfKCznW9HZFvurhRTPcJVsOT8OHtyQinHyuNGxtVWv2hCe6sMgMGdSPb7p
L0IZ+sfVqT1FEN1pqEupR3OzK+0qYxwaaVMKNCoj4uILGqw64QbQFPQ6jHaOYcI9
Xrilc/Df5CQFCvep6cm2cJq6oW7cQ0fpmyNh71kDEHLtCH1aYawVvTYImWuI7DPT
u/AN2mtE+X59efFrwhUwMYpijqHl7Z3EVN4MDX7fqPAX3Uh3pwhNgXHh1cAyF04G
VMny6Sek2aSA9kZl22DpxjCoRg5JJbmrQ4iuV6Crseq4FZbJ0h/oPGx1rEd+N9+w
0i/G1LbP7INhohUIJM2DEnrfdjV+D0sw4kQyNkXMwSGeGwh5twE+g3/9oG7cC49R
UI16JJ/oeW9PD7N6N3k2EoqG5b2vBUDVY4f0gJiFD+tXcoN1ifwf5ep1G/r+Z71A
txHR1RrLVaxtn8TjmhbScopBHtNcNRzMeg+FU9WpnutEAR+FRFWIfAeJ3asKPY7h
PzM/WfekGNmMUG7k67wKiZJJ71TIoqreOpCaEPKaPIUO14VlxSJZNpJmaLBSfxTH
a388rQuJRA8Cilweiv8ez5G514wy+4y6h1s2VD/mVNiV1jSXZedIQTH673MM1U1O
6EB8f8N6Js99bSFTcyKfa6mzwfmBIdoyHftcn4LjUKwcM3Qj+u7y/1kvzfWeJgGq
9OsxVBtdmJmtR8yBM3o6W52jbHD6C4Q7J4vShed6BwCdiYhMujkif2VLnPgDmT2o
nYW5ebpon4I8sW874WNFn9Fk+s9h/2xwS/3l3XvF4mhQBUqkyNXpP1TDu+htpKLb
XuSJXfwq+klE0OVwZlvtRx8j0cZ2ezDB1ziH+VXDlGY4NCW2s0wrTLGdq1nnDwHW
Ns1zO3XHp7Ri6t5aQGX0NCfEF/68DMNaRAqq5o3r4Q48m8Sbh5ztzO4NiYeNM9zt
xbhYBKS4Pbrph8vqoj5W/aHfm3oFkdkgCGxWVkYKojlTK4bHEh0NY0iRgzm5jHnN
JoheJuf8fwHJLMFexc5Lxx2gl0wunWEmAExPVWQ3NgiIv9xrjD4OaHHPSRcY3zqh
dVuTzwfXUgPzFHiQ/A+drxqcC0dsLhXWOFyx8xeJQgUeyFs3XmgdAjjl4GCS+8br
dlNql0ydFAIAID5FJ4oh+nZknKKmxY9MFyzfRZCz2mHeFFaCGmJAZYVafJChTlhM
OQyYMS10YJ/fU+6IlqlRbu29QitsHgsUSUZhgBMD4dNz1PxbHU/XkEaTS6w3ypge
/bdBpipLSxx7eXXyO5Nj2e/Q1q18fwML5pAOm/LA3f3yS2v/T8L2+Fu7xbsqIjut
Qpr+CsRADW9xUVoZ/CU8pECRa3hZu2IfUuOF7etpcjJHoYVj+tonCB899Wj17WrV
qaM9cqKzq+xxyqI7vnBGqtAR7G9LrZ1+WHi/No35WPctvOtmReXqdDH1juOUS6bB
ufHkest+hmRQaLWEyZrgdV52D4Bg+7V+EkKSXmpycitFVBFc8/gsk+iL3YM3XKxv
Vac2x5obZIbVN8rNKA3TejGEiOMVFt98aAk7kqw2kinClpCzYIBWa4Q76Eo0WQb2
5NqCXAP9JXymnvqNcXOoL5f+iyw+SMn9yvj/82IKYkKrg/qXPehx8Aoj+CWdizal
mKiaY53bt6F8wEnP1iAk84YZFuQ2yvNE9hx98PCl7PCUJSWQsm3+0mFwHnaE1iPn
kQPpTCeJez608sJ0pK6nSV2mxVyt2i95cCb3im+OWr5CzDLkLsiMCSP8l4cW4p6F
ADUTLhogCVe+wXAQWXokc+aOAXFfYlytozunh2esz3dvMRs3hOlk1CfrBUQEboMo
yrF+w2xGCkva+e97Wtn5KvddFKb6DGi/xI8EjD9Sn4EAJ2WIhreHKHrvgrrd8n2K
bPiaZ1zoaqzEwFLZLUpEhGWf0of/s8CxAntnMmbDb6yN09X2fNqOm9IY8KHxLJSZ
Jc2/CYvGX5AqmU7dijwIuCrl2dnofqQWCMJeqRqob9wyGXy6mwli0vXZ8T3rpM0V
sn+Pg/KrhmaD0x5TmaGcKBOFJzacSrd5aXBmYi5jN8GRc1wzpTKAL4wMeHNaort8
o9selQglexPrzbLg5cWEeYuThY1xGQyuJ47KXcaoo6QTA7mjWoL1f4d/93eDl/Kb
1BZhdkaCrcPyLDD8OCD0APbp7xJYjbh3zaJnAYe3V4Hf+i7Zf6ZnD+YRvtC0Oxp0
1lAY1Wb7RkGpdQYiyTxKf4jQaXKIONAAKaKjuh9zVQ/VGkQBcQNS95rcEMAJ4gAN
8zVmIVd/o5KTdEEKCiCLjN/lIO+OKAznPPP6xUAElaBxLuno+PMuxVQaOofpj1T6
CfmWh1+FAVd0owxY3O80CfDfIP9T3kBcCRk5KOGqDRA7penXyL+yJlJBcnKjXcKI
W5pxOVKylpz/nDpO1dPvVk2vKN2At119H3WqojjtuntXFYS64tPqWO2pP0PDjxBB
vGnG3qzlQ2hGVck9NXmdi74ZW2E0lKY6tu6m0asgjvaKYBiNaLUQ45jj92KL3KgB
m8JCCMyDkQqKsIbOj50VwNVj4+S/Xj7WId359lOzlp7im0fFNCpkHUqXALDKGRnx
pyB7J5AVa9xJZ5LzL8qr5hOwn3Ck6Mbab/3hzn3U/OIXZFjbK81bH3ZWgdRZ0pH5
VkUOjAKyXe/IyTya2RW0WLPojHAoLCkJU6v7CubVk0m17C83fcFNvJaSS9Z2XUam
BrnOLmgDRtsMll3goe0JaGIRt/QVPhc11JxRP44gu6bnhxRHiIEFUIc3nQy93xAh
+RrDA1VHa7yQ7UnlH60IpXCIiQpGF5foJ0wa6jIM6ogKeoMSsZ6mh/T2ehVJugaU
56qeRLdxQoHUqa0CDIiEaWrwabswT8caZlNCPuz6AXWGTB5NbauzxdPKh8xdqGK4
FDTFlyF/yw3bjOvjqyMOvt8E+QM49q5RUr004wFKAIBdMffy9s44FMp1UVsxV71p
SQfUu5w3vObm5pw6x8EkDTeSsTGEQsTjH0IJoH6fckwxBSOv8K5/azm0LqGj1cR1
6owWVTaYR2+PvXCfrW3vsH3s+dm4HXK7rGrOspjyrQ3QPcQw7dy/G5qWGjyN4yd8
VuSdTNpUNGusJpI1SM869z6UY5izXABPFrvBn9ed4f5TUap3aXWANefJsR/oZFTs
kbF4dKJ0/OVmKwB1UwdmoWxllNxEC+CbwK4tbIqzkTxH0kDLZ347cGu9DbHBezWH
J+IRGv2jnuWFmIIS1S/nMRSynaehBTpT2PWVro7EDGgjOXUKJ4q8XN3P6f51tY9L
eUwItoo+XSEjlVif3uy99gjO25UfH+3aI0IdT6HZo3gq0yyACKLR+WzB+uNNgE1z
Lgpor3iWJbCR7UVCPmburIP4mqrk63wv4UjYH3Ogn5fT2BnpzTsyAPN0IS8Xc1SH
F4E2bdVrA8kQ0Dt1maMFuAx5/M7NpFUUV+GHUgJ+unE2fpEfO3SRnSaI/TVVApSZ
btxGd2tsUEdK8VUcvch6KNiLlmrUoYgLWbA+eJBsAUfp2fmmWdsUJGVxGXkHPQKO
+sPUppo6YazBmhke0GGzopg49y46SCdjXdUyy0kF3GQy1IsjqIOrDVKoZODFcDEg
hNGYGAohVc3ILZKh/fYhMuhGEvLIUAgD7VFesZbUE04r+eaSojSjGLx0ZBawlu8f
bQs47OSfNWasH/dUXMYuqH3nA0AR4yPLCwd8Pzic4Y6L6h1tQOLz5EWVC6CiRjhU
hnfMRzc2SASmjr0CqGJHxFBkru302CLb+AzpMMZIXUXlFkuFpEiZkXlzIHDUsxPN
bLbsOlx51DI9/8jR3bJDXOumBsRaPiFiBiCcktP5O0DANCUwUIpEq9nJCIAi2g5D
YFfz542OF59z066UzfQdbxvxwVktJIDc/Dm7zlOceJ+e7XUzr3HbEyrWE2Tsw4dB
mBGrRSWN6gT8I4Lqz1SWY1qsNMZW/7YC/ill6Add3mxGfl+Uv4sqeJpvr6R8CBBI
cPotefWJVrrmBN2LYOVQTJGSiOkjE3KgpPOj/WQE2Gwvm01m7Z0aU0KzC5rFwqql
17UTnVXKG6BSXYiCD83GmoKQhJMKelHpg0h+4jvqsAmekFRpnWuw9Vs3YYgr5TFL
Hl/7SK2K4ge5goG4+nECrYxVDtO8m5mw5U2eR21b/2GeOtvNSeQFYnHreFFoB6n1
AKUGkiROMLg+TmymS7678NfJnEzql1y1QlNSS15KlK9+u7FuZP6qbyon04pJsIrx
4dOedtDI02Bd5nUj4re3fdIrnFU5xsf5k2C8xJo6Kfif7I1vNQ5wI15LGhexWcx6
eRJ197YydceDEvQWSdYIX5NUSPaV6r8eG+UKOAzLrGHJ2hy145xw5IP4/nxdbLt/
aQdLY8ePF0NR7lBjfQ8uzL0q134wxJtYN7IWpZGVionmdtImTBOwxmyT2pLNnJl4
OPDHUiu/VBdsyuXSN84qd10n3w1OwLURbajQvRJgpKhkIk+B/dP/nZ3DMviPzMrc
j6DwMkRPziFu/z171fupAQPg464gv42RGRQnG8sL015FL6+PC8O7yzzHBPznO00h
RXgrgh9n6h3XcTzhUSkX520qUMRJda1zpFbC5kdgCVlCO0hMLYE5fgZxtzykoYHo
FNJQ7aD+AqzucdfAKB+7HRBFu/7iDKvvcZG5Ai+HmdVigzHiUTfd8DIFEpAwZn/U
M0XVS+TpCpiZXYwxS9SqSOEvvPe3U2rV/wxNx9YYPcrY6ilMHNHFvbxwDtwgVH2U
817Y5tiIgY3bUaUZhafa960LGE0Hu7W+tsTz/8O5LwxoTcVSdAxlzwyARaH052gr
vGHVBLLmbmV7nvTQCfyDHEpHhY/HkG8g+AXlWPfexICRvFiCwjNIg1HC9Res4Wa5
z2ODdVQaBHZy949C6ShAxddOKKsIyesnLEsNR9QrRSGK2ZzhccAoSU5HejJvuUFo
Cv8gFf7EKinTOcpIKRyRNPeu+l8npK5ezgPDxMi4/jRQozAxy7mftSeIgZkceMO+
djz19WpY85ifd55M9dzZEEr4UmhaAN9o+lKNZHYQ0q9t/Bww3PDBoXE51srb3IjW
AnBTqCSfd7hzTMB5QMPa74xQ7fuEY4RWt++tVMGsV+ZXZL7TyRvFKg761WXOaboC
qmzEwQ3t+bygBXwvdcJ38lK/B8NvC0P4f9H7koLH2q9UINwkFyaxF6kseWWbISgc
L26gsGF6XdNmYUW1t6+mJStPbMM2ekxtgZrdfKba0nVzy8VxAWilw6NwbV4km5xk
7MS0N8DxDCh1Nfp9nIGmjR59lBjS/jxtFwMj1Pnu/BDHvp7tNWgFAVLoByCdnMhk
60vFU8hassnR+w+YzSofMKfyQgYVAO7uz7dFaF/ntRJsh3VfyUh+Xj3Xd3d/bv9k
ENphgFVhvVh0dthrWRTvf8+monnX2YqWhzJTO3cqyaKbMO4j/U8R2tMAVubMQ5wO
jH72VhYHjyM5aEZbtSW9iAtNsM6OuPncfU+c+ojZ31Mi1NF8wwb9CpT9ul5TIQs+
1q5fOUO/Q5uIVZPtDOsXHE73h+kVoe1mA6OBqRYn4GSLqF0RqypHLRRaJT9QnGJO
DBXZ+iv6Ciza00fgz64jnQOUayifZ3s/8cPOwmDWo3TN/lNhY9z25ZfHz9p2eiZs
GCI5bz8ShiUrk0t6pVO+M3a+XnHg2/AS9zlI20rti9sGcPgqQhvHs08oNqzdRnEH
OBKTySAg8IMDTVgiPyobM8eK/fhGAybjLplYr3YQUquFNy8Fv2iyecoEQEix90wI
+xkMwWm0KpOJYuhDH0ofZ1ipBQvPgllCbKNS56uET/hyrmegWQnhEcxb9xsWOoBK
l94lRTwqyEKSosIMtpsNOB/8YrnNSSqzAS2jY8asVoULMNz9Mxv73HwYNzwZBNeg
qOeSTo7xZiMMneLdvolz19lXZBZr7V0jlfrGoQp6vQBT/wbea1k4iKVnhDYKWztc
BRuSpGksw62r3gNPg3/2hUqFFM7iDc+JEoBx/BB+UzZkPllDbGv3y93u062tTLRU
2q7loKG+5S/0Oxzf8oQkY0zP8sHot78ag+NC4v22PRuieYjbVQTJFGhxoCbrt+J5
s6k92Z6vZHWd+uVbXTtcQpTebWUutkPL9bJ6JdWxHJ4Ff0yY/7Pzi8VZiZNFYQsB
1uqA3TBeFsPvI/9s4JVqW7mmtrICgRotnvmQlqRAOPdlkcHxBKNTPe5mm9qvcKUI
yD8/OQ62AihoR5MNusXHlYJEZcmh7vLU7mTZVsfTwpjJpcwTVNSWxOPQdS9Asvsn
NnElsQ9d3LrV/dkEhz1uPPjt0IlW++yfps69yCKqDVaNXPdpKpAshBp/KIGdVm3q
Lux7uVb4v2wsjOO8LpymZ5OJNUt5wV9qVT3au/mhYVJXJ++Th1rlRyExHhsKSjHz
rD6XcSqEiXlf1lbb/YPkZmRPoKBT++S6iSn6xbUAb2JUCqtYytRgRFbs7h9k/6/a
NYFFgg8QNzjtEdLVgfiK//Mp7POvMQ7p5XYvNUTxl4arWpAUeLS+eXc+hnhdMx3n
45HKQywkjyEUunKPZYBRQeGBoNt3i3viMuhzNLkARP2aI0Hb543CWKAhRvbsQSXz
wkfO1yxUyOA9xpIpzIkPPgxFR/eb9A78fnHLfCnfPpL/tYEOAMYwUhXJvqSynr/q
ibS/loKF6DbAGQbmLuYyIf7X2i6zKe2hMpD8nBMTs+YOUzWTlKodEM3aReVTHRJz
YmcayVulMMQD32FiyY2XMfCOGz+NXb5ij6hsRNgI5OABWMdhvprYdwcGdzSt8GtT
z56CW5J50Zjrnx6PcCJBu/xqn+IRzPP+IPMkNTAj2rzDpUs5wbuSaqb6X4UO/mj/
ueUGjqs171tl2ukFZ3hUfEU/uHVnW7JPOLy3LTuDbn9dFRR0xI3NWOVRMIRQqM8K
1jyJFqnJaHHF86cBY458Borsb3UAA7S0FLFMstKt4FbLhOEbqv+yNcBi1z37zqwI
RCpJhYNHVVs7GTgboXQQMUiNcZ7O1or8XTnzirSyRJKH0Y0Egi+2XVyIT3gkHjZJ
YZhCp0XWGvWYTyaAOopU/BqcZCDhTqNAnbDysw0X2n4qX/bhu0Q6zfkXRlrMp8tV
2MC+gYTtnNB3rocJ0diqNFZftXJIlE1uAyGe4SEbDd29SYsltlEpPuMi57OjT7+S
tMCRmK9QkF2plsqUwVg3wx1l11Gbv65abFIF2WehlK4K07xFWFLNGO9lEBRPnUCi
N3mWZkSKOsbh3rwfCxUBPD58t6Z3GlhMynf0sCb0+xPeNOKSLGQsDZooBtK29r3x
vAG3ZIuPw4XZ3hIjW9qHi7XXPyEMQ7SBuMuT4+AtAMPPDiDcj1HhaXln0K0LymMx
m2rU3s/E0b/xRaDDyRaS8+lMv9z6Iz1zMuP32EazJ+nADcZDCWvSO3d99ATZTcXV
t65gjvm11GEIn/qYEGFAVzvYnfR3lwkdaO0fCWEE//hScHd4EIhkXvY135S3Gj3D
KAKN3B505hNHmCuAOtqghmWGZG9uPjIH5LXPZmUG5jcQZWAWc+TnawD8oPKjsa49
GfBLwr6QpSkDWxIGsigO8OeHAL3dYou8LUANSOWyhZHHEpWq7BT3Vr1U67K9alUf
SRsuDHMYSPQ/Gak6s/XskNVDx+bGSJTfcz08zi9dEjCw1VPcnFrXHtV5SBJfJsRr
06lij3322PQE9A56YeKnf1E7ZueccwqLhPV9+bQZ+FUO/AJ6pIRIT5FlR32Tss6Q
oHJy/UJd80k3LOGTO8CIB9f4KtXoFQ7o3giY/bgiQGKUz22T4+KsAa/g9ik39cfs
+XB1sOixTGmJDml1UEi5GVo1Nwr1paRvFswSfI1XQBix4ffyPve9SDCG8lDOFxxB
nZ8tK/vaJ6JU8rU10OibGxlDj4EAAXi3QDqiOJMFJ6rit7/xiglLa43ViEAkdBH/
GnS4isIPSnTAF1Sd6KdSAqYa/0o44zb4eD0HM7EuZ3Y2fSEtrxOTzIBsa1WxeBhQ
wHLbD02aclNV8/fRjH8yd6EFRRsPmPAtHpTOeZlgK12Q/KtnS4Lb6yIMl9S3CeZW
EkOAlx1tPe/PLbUNZf4wX1vg5VBtlwNiDVgGga3jn4wLEJd8mbPFTiAinrhULsZD
dBltmnI3bycR6SsF7kenFzt0948aUivuPJzWgWWLk9qiiahOzzOVUoSFaNV/nfw8
92cwC6T5coqlpEHeBvSWAD3h8UH9AWIOIlEGcMHehyTxUoNal+Fkoa9jjGUinE80
eF41/MdeFRwQpQKQ7RIgEZxAUF+cfNg2v39U3vGDLsrUpnKzC4EjpYQ6PCm7hXPd
SneldzfRt3VGFTZMwHMNIfILx7rc8f/UQzXnu0m+FlQrWxBXF/io/Cl6BPeQWt3B
SLpBmDOfGk/VtJprqfk3R/kungLPUwavLuiTNlOnYBRLETn4J/QE4ffej91QFjvZ
iPGvcbM/lfx0XCoQ0GkNQ6BUx4syl8VGVuA9R6pz/2Ig791hpJNSfmPEdwzkIepS
5QWXitgDjokIdoLWOBRrRUJXbxAFIfvwSNFy04T+U0BqkvyqDBig1I+o1vcsIJ66
htAwFYkiMUBDGSfb5yPzo0GY1Zdgr1FeIU43VIuuHcIQWXiVFge7y2jP5yVGYYxS
L460KvNXdGaXjhpFA2J5SSJPHjUPrn5gXtAHh27+PBSCgIQrJXK3SpXnmhGSgySz
ZDm98K3ogIAKVg9pUoCnoPEn45NeknRJgbyDnCjh4HIkaKOFk2E7jDw57jDaAEAW
0bmvaPJVG57ueN3CVJyh91iIrmk9uzHBT1egotldd6cB8xKICVnDThHbaYtky/NT
ZZXvFV5J6lvrCTdjdsx7rZ4fAj/7jsrZlLS/8F+AZM8hvHLHmq069C/WmvACW4EV
G5NHBFuq7OJRvXnv89BLGM0LGx/zJyrAVB+oyroUqFyWJrJvQmLEgOA9RLAKamhI
SDmXZfG1nztsJ7n5nfWGMMr9ojES3o73SuSaoCfkTescbceFKNpDeNvr2DpNX7e8
TQiK2ubhx3oNRPFVi19ssFy1oMZ4Ox3GO6OMWLscG0JJITNItJicXYgolzc2qY/T
FK/mn1o3Xc390utoFzdvwd/3KlbfPuivcwLLy/0UX5xy7hQyPoPljsun6jLg6/Fu
3rhMpPhGG9XaeOMGHyPsz/4KBjLlHBFal5sBzlLqp+7uSpUyQOUV81n4+hieBW0X
4urmAAG40yyhZoNbMqZOcPltRBm2C7T9t6aBxZMF+6bybPcJTRFTgNeCCcXZvhP1
l757ikb1C4TFs5cLurUAAyXwG6EsTol+RuPSldxYWtJe3o5cDBFk6lxkKoWdIAC6
ieh1mugtcd5dP7qgUljw9B6jvIIVW5tysrHxDjMmsPfBifGnIPVQyC4FVLvOy0Ha
IS7646YHzfKusg7FtRfuujoFFkIIUgBEvrMNguPTWeG/ZvN9C+r7xsWnd8YJKuOv
jLP7MSrszynw63PLoU7779rq08WfdtwPTdT3jYM9zuJQ1DP+6Yt0C+1wjZEF4TWT
5u4vJ7eCCzWCB1Dh92UHnN5LMIVPQt1N5XXRyFXh+ceZQfK1VQxylI2QA8aLLKNK
MHZ5x/6H2Hy6o0wDjY4HwNlzeKOMYpf6YxxCMG8oazmhEmNyCokscSFENaUc6bW9
h8hEpctuf65BEvzEPLlWjutjf43Yptsl4jvvaVlysN1dv0e1AUDsBa19NKoj2j9H
5zroWzd2CH/f5kkc0GMznaCTtJNFan35e5B1wnHfDqctHzHa8w+wbFVB31sw5qwd
q8xDhV6l1/iS8iXVzVwOyI7jfefmZYXjgAPi2X5zfJGOKDOEdhafjNyXGeMBOVa+
nERpRVmVI1M42HWVU2fAq8hJcy5+9J58xVfzB8iAZKJWX8beyiiQoagAQFA8K1Go
sxrn6zKULluvJnbN58xwSEsRBN7o2LCFrOY7niYaMBlndZI9p3/epuR9McAsfSrt
IzB8X2rdYsJ96/lQ+uXjni6oxp8iRtYGOIYsSnUA1U8rJv3oxOkp12gV42g7piDw
ee9Ic46fLV49rH2OKNDdtGIeLwn51IeXGTaB9acnf5nblzsTHeurQOtf4UF/x2ym
I+Z84Vdbu5cadt+PSf7VeP3Vdgbhc2vNbOsHDkD2GAPsjnpHcM/Nnfr/3AaB3I6o
076JV6DQIf0z/bO7JaZefjJKYlkjP17x3I5pet2cPIQEJl8ky49IGSzkUcpVve+t
zsVjZs3HaDsfpyc/vp8jDsoBJD3S6h/qiGI55hfiFNz7lsjMe7RiYDutn8koqAbQ
EKdT/EHbofCZxwkzzcQ1ghZRcVwUQc/PdtyJIyKTyV2zCzQbwZh5iGLUW8xoXjbh
mBw5ZJjue8ZzkQEI7kJ/m6FOoHsmTLtZYd7o/+sgDnALQ/6OrlBxjiWCTptzYMfc
hVMd0F9PVYRKzEyWTkHOIVKEOlkKLnxyRKwBfX7vm35J4ipxDPSRBlcbbwskLWJE
EpRoa04SBNMytF334helBZYdJ6VZhhXtuGzzagGuf5w3XpJDA6DTm3oDugiit5Gt
w40XH9LQxd+AwG4WsuCLE0RxwlYjILpLuBxcTpgeGHbfKIG45dWAfo51sMcjgZp/
ImLGtXjcfUdMPciskojmOGCuJcTJx9d8u39fMoI4UzkoGvnqSK4ErnsXflZbyIk+
/CtpULFOAtnTTYNRUSDoRqkzN+C/Oxbl4u/RlErnLs/oT182yA78b4iHd43oK60X
ECrI62Zvpt1TJeCl7KwFF5gVuT2foHpO8JXmV/Ss2hupgrr85MQxPgd5QLX9xT3b
+OFzwRKeW2z4nRmcWLANxJhHa+G338NyNfNvsPGjZpRP0LWqwjUn2DHjv3e8HomA
EexgAQIO+RYLToXcOYl6/MOF0YC0GZnT80PCEBSqqhGICOfp43lwDrxHoXmIFPQD
tgDl3rBHzXFDXKEdm3ZNzZ6s4iiYiYQklxyIiaUWAUrDuIPi+83LsrvudJ9/Kxib
R+qj/pfFgxDLRhylLyEWOES3aS3SOexKISgnrAKgzx9zVOCa4MDKlvpu2vgdRe1y
l+daTwtQc+0h1YhdFmWu+cLwQgjufHD0t4Dkkl2A9BGyHFcTZsWGIHhbgcjOGL0N
ccquSKTSl9CAs2n7qqCbHREEW68tEDdP5BHXzFOjzpk9h6ILL9YWqwp8dAjKemU8
oZs/b4cZw5ssiRcmImnhU8/Oc5XOYZSHYD1jhh3aiWKfH8D2t0fGazpr6+mPuVlz
OD42YXXGJcAmrFW4UxKwyKW/7Ld4xCUGk+r3u5Va4V77EOJPr3LKXuGRTxUPBV9l
b7zZ27V4znN02G3DMmhWB6RD8ttCzWUTqx+AcWQPqQI8oztU3C9/lsi9MjUAaJG6
r5JSjYcdZA1XGeXntmTtlZIjX1dn+pDn7R1IYZWP3zDOm3CRrgMcyNCm7n2Xze2y
txf9cQw6EzzWs9FqK0NVnPHvkQe0o7h9HgL0eFQNeM/YolE7YWXS81vnKnIP7RUE
EyA1vo1E3rG8ueonjaBBflOeUJGXd3wjUiv9vHug/Ty8lGVMJVw+9z+QnybZ74Ie
1yd3+GYQesU46Rgdg2yFdMHr/gT//mjM2KpjvKfC16uCEkveofgDmSU8YeB4BtmD
BSbA21+XNyahkaynVdldEZaGu5vWANyYkNpG4BIwPlzClcma7f4lmTrppy+5qfgW
coc5eBvBuQiNVfzbG/TpZwNUOXOP/MgF0ynLX4zvh/pDgKCNZRlQ9835AVUmU5yi
hdHgRJyh3xhIact6hcd+GtfRCm5qIaySmyEyH1idIR0Uaw2OHDHOQpkhHvtwoQmx
DA3/FPatmoWJpEDzIjpnaIYK3EUKb5zD+tlbeZ9V3slzfEvl0RZWs2ey6GNSJ60C
37yLm2H3qhpmfyRFSh/NUbQzI1h2r3Blav9QWQ7chdaShgU23sCyIJTh5L8/9OqX
BQAMyhWyz2vyLHsGk+XVbe5NIocamVEE3kkDCs6xCzAEaFN2YtMq5o07PQ5lCGvh
qdmL+W0n/hP/cW3zMf7EcjweX0VJjQAFd43GNn9B1zTk4ewJtc9k4glIvuW3mC6x
cXdhCtALpw8aE7EM0NrfHA4uchSzGNjoAHH3Ds7MSP6Gf+4FJsEyQRyfUvKp8N61
qL+jQ3prtFN58aYqUcnSEqRVYjYDks6e/wyeRLSIWNQh8gyKNEiHxKGAmIl32Uz+
mLAwHeMUmP2+TmA/xlmvvRCH5T4odYH3tDWxaK95W3ijRNsYlAczM7cPHjMzp7kl
eLO8DMwsKPR/GJaQY7HgaT4mVXofd4HIrEIHb62M3ecJcUlQrb2lapWJfXjie0Fw
sR1QJ1mEIQdk8KRDSTHzBux3X5k8rrMtQYwUUpsNdCKGNcUSMC9ahOXJYw1Au4uP
dKgsFd+ONKDgEO4dbN+8DhjcR3nOt3wreHe73HSsh3CwzQa2qt75R+fCj5UghQAm
i/Q+j3YgKyRZW1fRChKvF701SxRzJqkevoojiPyE5MHV5Br8SOSPSxxHRUwXkMRw
hMQiQP7LHQ2Xo+KbjV3bsmoM1v0fyreZWDS0HK3f07j9zEXMnpPc0pweBaVUcW+9
F6gpyYxhFLeAt+QwVLDC86nN19Fi9VscrA2jKPoBUulq45H3+ZssZxGHeLWpFPxJ
9gZ9+OPvhmpNY58mok+2948vWiE4e/NpHo19ZREKGXbZqjHy2Xe1lF4qEdC25U+v
jPfuxhEl3Ojfgvxl2cnTF5cdZ1ETfYC/5SX/h3NiYGpKX4+tm0+88+zUF7WU0FcA
nj3b/bXGOIp+PAz7Dd9z1bijK3B3RSlvTc6XbAXiwZ+te1P28g+EG2kQESelIMoX
gaKZIvg3XJIno7zjiXpBJ7xo/84XomyWfF9ZsPYqQYY7IHPlWlarDivNCcKdnH+D
gJpgGDhHnxZhaKGxH7246dsmSqk0Ny6Ana2WgmsgB6mEe/yNey+1cgR4Df6SonRE
Xs3W7yrVYVd7i8v9SrF8zNeldGOEukFGq9sPnyYiEQrTtfubjejqZLDOA+BW8jTf
WT95NifBnLorjW+u+kImpE7JOjn4VssXh7Ms08uinhLvTdNYeayE0rGuvJgKUam/
sx+vIOxiIcZhWUfZ/HEsjNz171I/WwYc1P4wLU5+K0V3xV1UHfMRFtEQupmamGAJ
w8sR06hXj4Tg+A4PnEh7mPQvWZ++HAecH1nN01UuHBIb4IKplVTbE80oYOnf769w
cu0N5i7DbPu+mXkR6hcQAfXOmZy0R3lMSpNEQSPgJknBYAPSkgTH/5oUG07yyCZ8
6O2Ayx6Fcz6OIdWm+As/UP0PG6vftmCvkWBl00+8o/xhZc0uGTMw4YWbrFqdiQnD
KxjcZ6MvqjsPDSbtbq/vyuQBbYm22RiTqxcISsQZ9A5A5/oRYpnwnuL/EzCv2HYq
LqX3Ry8AWkO3t0HMuk85QNfu/0kqnfHfuKzK/abg+O2z/EUm1x3vJ/rkuBBpy3ET
czEzpGrlm+B3hFUFMVppMnDyUkrgKjO2ZFAGR0UNp1iNc7PmiwqSEMTXW9Cde8Ny
K24w1WYCYuvNfa+VgUAesYSA60XvniTUitb1i7eniBSdup1MKkVlB5eADlqlI8Ic
NXt3cItj3qhC0GT6bke/71ZM/UHcXoyD+cJ9IDuZI8S/w1NAbP99bLnlPGzRW5Md
MqMp1RZkbr+mnWxPGXXyi2CkbvEl4JVmADBQMA8qMUhjIx2ah5Im1UkRKf8GxcvW
gsY/UCYnC33XVTbZLQ9f9FuCImCyWm4I2pXteu0lyAXI/ttlkHYuravVELfKLMEC
045khbh30/XTM6JNt4/kKy8sIxuNsvfssYg+U3bLI9+kmFb8O//7xi/3TvOiNrFE
ZV2IPE0w9MXhbrFIFN/fwNoqJ0QlMLAXqWEO7GawTnSQhopxIm90PlUvPCDdMJ22
qxdAMMWL/hPgAGpa4HAWhlYvzyLIgeegPf/YWrfRc7RUOZfk3PU3Vbux/SqKMhRw
XKGt/QTwIbAWlvPROCJzNyHTcAJXcnmDcTcstUik0cVfC/uOkqW0FQ4cpJnzcgYp
KRxJIyIjWCI/5W5kcRudjl8PbA5FsJv2ufMYQp1OHVgfjOWiLAG4NhWValixzWG5
Qjc1XSJ9/CoObKTMyBDMYt1YdXlAtYxX7OqaxcDOp2+SrnfU1rQNK3Gwyk64rtAt
Pwc2X4zvftjqqZHdr2WWvpNSfteLlKRYfRLaYUkDg+xrG9ocIWIMYYxpXiJP8mIM
6s4rBkL99USodbXaeBC2KBc9EHQ1Pt2WuYNOhCwDi0Roj5rc6Tlrzx8ssRuQmUcf
YZG7U9KjThmC4+lL6GzJRjATR3HjyufML8lFSUKsju743fCOj3E4fAlOVM7r4Ohj
ABwzlmaL3jGaW1HZBwbBck2tIlRRYhzaQ1/ZpXgRTOaSC3ZeDalV/hPYZ6vca65t
gY89HpahZvpdN4RW7RzCCopkNGBXW3zA5IlGuTUnbD11bIBPky9xqKv+jGSuOWCF
87jymdx1Wg0UgXxWQzXktGSgYJsjRMC7Jnc16oiFWekZ01emyXjzj6zMnb9cCtpB
b70M2QKxsaF2QGrnFV4sOLeV/SUgdjXgMchhZ0e5HjSQgkWPCA46fbOdPekesA/3
nrZB0PlpJwwRVCoNRd7Fs0exkqLZPLJEdSUaygvAYxiwyts4w1LLcp/5ecwiH5Lm
nV21GNqQNAKIpzkH/nT0eWaYCIfPM79Vk+1xs7/7Eq03m1xVmvubNjzfwFGxtmlJ
OpZJl28SvcwVHcrpC3wmJ5gWgITwqN8BP/jScKEQu8agCyBbEH9npEduCNpSXFGp
SM8HFYYvdTsCm48xB1r5+2a0MQtUnFbkroyNrCjZ5Frzy3kw/gzCUA20oL845/S4
WGfiaFfg1XzdSR/8J7q4ZC2GmQz40d/VIllGUAtz0LmD7EcCopfxE/9mq5vRt6HI
VAQxPNXGvdADzR6+Uq/lVgmkkUdJLkmqftB9/O6pQYisCE/qZzG7jxCfNduALL37
3bxxxruNDoZ2fGf7woWym8Y4ubvLwhMeK/nMIsSPSJfSpmCsMkUCuwU/SjTpJKNm
m5azMdYa0eWC0sExYjfqNSrCbwlRmer9zptONdyD+Pbx3QfcfK1zuZljNHR5JZAM
5AYdYBJMK/oWxc/u3nINaSvPqxHRpo0sBjl6dUa1wzLkMisWKpnOxwK8GsYGOSDr
XC4wF0xrWTV/yXnUI4dZsryWeaLNLPBRTeCqBvZxHkllibacEuYWH/Zkj+KGZTC7
CVyl68TAe7deN7vD9uCsXh3FaUARNwm0pvteca6yR9Sx8SSP908k9nFlCV7BnGtx
FMQ0EhYE5PSEKfnT7zh9i/zx+Ra3be0+HC/6zLrhyzp0AGDRLFE7XdFq983ghTlz
a5RKdyZtWjv5pxrKnQXLHVMP0wkuv7Gj4i8T40jHfyn7+OgavaMCa9D/vmZVDFNE
fxNwa7VZlfF5zJumTC9rCtMncD33kIUxjCkH/uunbXxyt5UlrDhhKtrZ1vsygT3U
i/BqA/3S8O+KX5dvWJLTseJw9729q5tyrUt8JUFNaLBhJce0mb/6Ez/4AYFR3Vap
gaFrs530hiVtoSttIoSXB9cRxxUlZf6F7JzM6x2dWr/MqbRoEbm/Jp+xDYVhVc1x
hfh76yVAl+yegh4ASJDkXeZze6X8TMkrp/E8+HkKd4V9w16dBmIrIz/9LeOhvATv
kDS9dGBNDc30V8SfV8nWZXhBJtfY9B8EaLYQVJle9g01jDwJphnpBAYzISJC9Jfv
wqlw6f57kLMjum65ulFV2M/8597XGZxofzMl6fJYPstJ/bFVTjqD4uI8ZM66kTZK
4zJZhBO0x5mKjaG+sT4/ErjkCOjOMQCGTdP2muI2m/WlDwRHbYtsxbRFppSrLFEL
pwDOals3jRxzdF3U1CyNGDzNoL9735H2wt3krvJquR3nJQYXbBbDlqhk+6SB/4Vg
7pYGh4jKHgaYfaIdOH9bTpelTFP3CScHfdrpznGbaAR/3w3g74MTJn0ybrWVcr9s
cZVXEfkT5KQvWJ8HmMsIm2L3KAjCk/hV4mwsS+AdRmtgRAStF4KSLuZ5elcsrQFg
gSVobHwLLWAHP3m2RzOpN5Y6uNKoV96n6pnIuNxXQP1sHSKlBjVBInhHalzM680l
b5VdhM9d7m8g+n1LWdcHSlRVuOc4ewne3gtifyQ8e8dSIrzir5UxANoFFx3fRP7X
Zady94Bkng9r3UtcDQQud3AU/xM5A3OAVDJCsJcfTvtfbUrqfKA9AsUc1iY/crJO
/+tFZonxq+riCOfmaO3IKmlvZMz+Y6gIE6rp0peZ3xq/nnjYmKVrLjp+lzEnmaSC
8wONcj/sHt6EwR2zo7x0oYBIggL3rTsXthj5CkVJexgtvEBU41SRMgnJ43+i7cGn
cu9dEsuNKqWk6Fdtaxa770h2sZdnG01PBwCRtpTQelB7WmTe9/Bn+LLWqzCueD4W
6MDJ6UsL0k5upwxn9CT6luFFE4GRYbR5GIZa2wx7M2Yvw3SlYf79jwCMZnNKKqlP
VD/kyQv32hFyQ4HXZZvTKJLvNsYfFpMDhC63f2N5oL/5kFC5iE+aNngL1PcFuSUp
TNyj/cWOGqWlHzS17uLMQHD5KvK6M8A+QdjI1y1VRxhidZKRXKlJ5v+KBdTUb5a6
i+WOmA154nBV76oPMcUskpZ3dqqIERIL52xuqMcbYoZbv9q/EnVPfny4jvfdPUJ4
pU7ensNET/b9DhaTX9PPgWvTfyJrl3VSXS5wwXoDPr0V49yg1oHlznqR3Q9a8nk0
3TKefu4LYmSNzzd8GRbJ4JQIc/pa+uGXljbmMkXknXU8/7drmxhAgXIyrjrGQk7i
e6IuWAcvWCRXqakWttN7ydGM69Km1pNqPpKqQm8p8Q0wTFmhrEo/O189XYzc4rmm
awbKuqrZgfvUADmOmYkoCT+Y+WnNqnQeFFjQfOwCe5SNLboeI4hsULH3mcyW0/VW
3j2CFw4tDXE92mOcF1cwV4Uh8DEz7pwlU61m+gFI6+A/RN1zfCFlkoBaMvKUIecZ
PwjQLr9N+MeQAIDv8nAx66Q5/aJB94q3Ly9j6T06mJ3y2xrQwOHAqQ9DojOZsMmQ
n9pJbWf/8xr3tFKnc8u1UjfIP9TqdTdhGMEUVq6sJxZNp6pAwLbcY6qEOUwAOp1C
YgK3ikxI22d/7y3UAV9jJPxU9qzGf0SgWNOdcPfo4GjMdljFZNEC4WtUs8BAmp/H
TbTafGWVVsCNTV85Hp8jVpyLQPKOgeOvKPlCYRgHytVbURR9W5vFkGNChMoKwkUR
1HCH4fOHaWb7S8qWq6xjFravlqLAJGz5Mm7ojT9Jd2VJ8LADAedUF7JLhZLROLxa
E80Y9QwoGIZ0/Rr3FAVZ7IwXgaOHO8ZmIyevYogBhZ0A0E8d+E3M7KpARXFnOJCD
TX02DHcddRS5T/CPHdrxq35SRPO93NYDR6oa4ZW0Sa8oCiRJ2f6v2HtE4O3QI5Yz
26yL1knjZ396ZaRSeVDuABk7PcakbbbEtqwirkI5hBeBLv0dwfTTowse/OG9r3xr
3tMHYhGpEDvYQppC+Olb8mN6nmQVTTKEeRJdI/4ar8JBd1ygPn6UM9bNd6uD/gjK
xrBEMiQIblT7k1uVPcmRCFkbGMisUKJQaecj6DpuoHLa+PIoN4kv2WBf7vLO8to0
DtAagvrNbXeVqigKwSqGTcHfaX72CrO39BYTtZFyUAKtw1wodIJ33Uczt60/mEnM
/o39yAAOr2ctXjPrehd3SECoela0Z2WuRKyqwtDUg49qEP7t+sv6iDLKquXr4UJy
bDkAdBIGkoQNpcZrttydsrZQ4nfDGyi22OAn4te3kGR+3eft/bb+XBX8qdGbMmeU
T7BvQphglYI/uOsGcNFUHAU95PYMtzrnAts5BRvMiJTaQjf8v+J1vYWcA1OVFzwx
jeK48saZYf5Kpg8MID8fDd6pyhIt1QBwNkFSFyMuXboONjV/RJW6FMkrw+cDSYFp
sAhqGpimKen+RauNEZstGkkwK/2Mh64UKeTqDUuOTkoKQbblX0ruQ9aUdDT1QDcT
DRecfDWFif9mli7g95k7PYVOXqzfKuzxojuqYHn0MXWDAvVe4xi1a+K7Z1RznPtn
HCT1RTbqJrQ7mh/ZybxzYNv39pVN7QldX4F6ODw8a3SpW9GzMhlLEX7ORLEHbp98
TFytt2X/Yg8ikrf98+t2q2upz3Yg1zIjLjz3CyF44QHcLkCIymibsRJq7LfUZ1Y1
3ZfgZhBjhnabMEW0KWuWPibYbkjIgqxOdzPX8OtG8tY8pT3gzdJ4lbytynQxNbmb
qqpIx/4drq18IkQHRmYQWxoI9G0+ok8npZ/DQ3oDFdqE1vUB2gsOmD8UAAoaJ7vj
GG9Y9xa7QzVTEvJxsyuPRyd8IeMoXTGOgu1fh/4ugtQ7ZgcktjdiM+a6PdDqFDJk
0cu7K+kuwevAbJLd4O52D7Mw3ZAPZgqU8hcMQH3wD+9TQlu+i1dxSYbFjFq+yHOE
Tr+uFNTf0+R+B0AKUTOmVw183oK65HOp9zaX+/piesJo+LbBW0MRnLCdTLvSNj9w
Ms3oNMcvpeax2rNn2/n9FSDJvNAfGi+TnA3m7G4HfY+dtKpgiJ6Q1baNE/b1RxKi
mlVatY1iQS4ADRsqF4r7ajmxKnodr5sur3tHYZfqqAgFLwtDbISBTnNBh0l43C8k
YkIhymtECGrj7rQgYlpGEfZC/KB51vLyGF34NwgakNX7GRah+aX3+Mciomq5jhaT
wa2EgCjB+i2mB0evfLdeib3mKsfOK1wB1S6M5zQLIY6yYwk6gEvwnW92R5sMxLzE
LcAmg1f514Fp2W68a6angfBZK9vxjH7Lagk1dZ4QEy8iN5YfFJ7DvmW2tL2J6XzZ
MY6hZnWz/67tNMmxOnEf48ge1ug9MdmJ9oAn9+iwZyioiFk1q2YNzNx4RCUqWp78
x1tBusuTsJZ5/o4htxW9YfiSn2nmjICz4Y2PaQ3cXsPAaf7sDQM5qFOYEYtc0mhq
ks2XD8bDEzn0cY6D9e3WIermaB9jnnmx/UStp4bfYHS550U2pHvAqrRiFvOvJ/XS
49WY+0BXz2GfM+Ov5geikDnJsWeKKme6/pc7tau0FP2TYKqwCx4NH44CRsGAPKEi
gphs7WyzIktiectxZC5H0McP5msdxKhNsY1THybiSz9AWRqq8A8VATcA+VRu2szw
WXcM7BhhBFrQ0aXTrhf0asyabiyTJK0s9yCMqGAV6fLOvd0J/pyYR9prYAqE9kRM
oqg9H61E1Ga6H1+Rv2YDpIxO2GAaqDMYuVnR/f7FwsVUZS72eAE/ZrZZKPgq+m7b
10rHr/w/bA0LCVMRN8j3ya7j34VZEc397P33G2y2Gc/n7MGXP0cEU33g4fzWPu0N
CXS260QOeBzdEiJcWYQViCNtI97PCWSKvpZU7CZK9xkdKAcrS3CELYpcwZakHN6y
1yR75/Zh5E8doKfjmkrhBzj/fZ3ykujoLfs7WGMpLtsk/UCzJts7rLlybWexYKMO
XFohbNmVKTugtdxH0ymjDcv1l0jJKpLtfsOSI1BB5lWqC/k3hoQ9KPUTBv0ur5GM
l41PPPVtVJoafhDDY8X4HjW5WZSJOI7RVPwmgsw/W2UGZuX4UW8HCOlvcT0Wer/g
3XAIP/vf3KgrPkN2BG0Tee7lXdC2SSeiQGzOMe27WVA111p8ZFe53904OFPoDOPq
ZYsi3USwBsPmI6coYDj20vVDSLTOg3+zBLQJc5p7uTiLFTxRR3frTBCBNFHa8+03
Xa6RlrQD9vU8sIkx6oDrNjD62ZFX/fuE/01b+rR6pRqgYGWLGsxvx2TYDoci50/a
Zx0CmNeAWyEndr8nsKm8v0gk0zm64pcgGR9JjATbhD7k8j179WPPLRx/zaq6vmdv
kG+5DRqwdQ/nccUm52uti/EOgP5naevulHYkuqOf9MevAM0d9Z0Iird0CUAeBV7e
3EF8eoTdKN+0jXzCZb/MLZ3owqrMs4iEAE20TLbnFNxlCwfO8M0I0PDOrQNNXzgL
TCtArgVcTJipSSv4yNotWB7Tlyf3Psi6W3BYLj2ZKMdSAwUwucVarOCIm0z3DJ2F
7tji5BdcaJSvGXfHk+V41lWqIJG1yvsLfjthXVza4VOf/gdMJ+WwIUrwogL1dirN
kT9nIb8YoVd4yZDe7JaRp46kaJLEL9N5nutbQVDr5yPVlxty2fTaWELjNcVLzlmD
FrVcL+5gcWXBZTep6YH7M9fSmEKf85Atnx3kI1XJngCa2T2uTprkF8TnYGgmozk3
L5si+VRB2M4l6SIYdxpVqv/q/cFRuYy+awAnpfAeVMRqyWf5rtJgO71JcST5nVBc
hz5s3L6RdfFi8lQzcOLndr547i1z8X6rekjyvjhz5fDmS+bXYszC3wSSeuhGLnKj
Cf9E0foDfYZ7eDeJ4C6dnwlRajvcvnwb8IFyIcM/pV+Q+5bBmdzpXOMQC4FkSSU6
IWOIvXpGSWdWOHOKEqfS2PVMCO9FmPq/Y4z05qTlDjOhb2hVBqVTM2AnW7rARb++
u0byGVDrlGcJovAaIOlTsu9NLUfQ/vZAPsk0nnC+/ArnFSqZjpwwls3VOCjzkbwA
wnpg8Z7++WM0vVlIZSsm9v+jLYk9SYfuLwrMCbXB7TGkz0sJ2zPg6/Wb01Jh0mTz
hkNKJl7ppzs3EY5i9FVPSXQkwivuEcK+8GWmhU9EDn6twZvIke2JFzYikgWQqwtJ
AgUY1snq3/I0gL7lyRXpPBCAWPk+//U55CAdh7gfQ/EPrQIw0Ay/YLxPjPDsERcJ
7HQUsYjapI5hiQ4NhL8M5lxBnHA/M1gsrbegAqhnlAVM8NjXCQJG+IlHTDnlfizn
OxRjENLYns+BKQLTKxbr/rXghqrDHQj3yodJvmVXH6D06EkQnOy+WKSvbOMSG3m/
LgUq2X7CFKQe5aGm1z9Wx52aGblrquYzdY3UUDYLPTDJ7oZEFJomkaQSWC2Pdep/
/W0UAc/+VUhr8b6XQ1s/Ur8lTLTh06oEiy3KLz1PrpLsc+vb6PS1GBPV+9ElPtSM
GUCovTYU4WI/RHDybcF0KjEwVugL0kcfVFpot0eSMJSWuZ1Kd/z9vqrasoi4xqZN
EsnbZTwA5SHdiIwQg9HhYzGsr8Ig0tLtDeHvJwkvsHu+g1VxntBevfz5kO6iBjvT
U7n7I9Ix3eooUeBwPEW0Vv6+hGMXAvS5/MXUSWbHHf2tNMeMU9XZceJ8yvAmJdXc
Bc/UbFpM1v7j62z+Qj7He4w507S0M8lGd9LAm1l7anac40dh16igJCysjh5Yyg3f
d5H08w/W6znptUgohw6AmrXQIS95z4/efckOt57pOgRHY0VqOqsjyT7ETFyyuCxJ
plNyG1oa7dXztGRnsLdlqzQuHz9NzEOOrrsnVWrd1pn9baaJX1WYpZnep8/+EMLR
nZq6Vl3lD7hVEk0jtJG/VyHPwzqZwRtHmXK9yIlsVHlbON1ICfK32Kn+6KUTr1II
RSElgrU7Lw+Bf1CZXl/IIKLiZ2T26Wd/snIICBfe5t9cupbK6DrzoCxpZbT9uG0T
F52ZvT/R8VPa4pXprBfKWfHiwwEyO4rviqY6oZvCMd8HyPlVHRlYxP7bOIPEHYVU
9hn2L4z92UH9Qb2KQP9B0RKZIkBVhTSZZcei6iqoorSA4bLhabuVa4B1O/f177vV
o/zE4uuQ9o0yt3/Jmoyn8XA4NBPR5aq9X9Cv5LqKVGtXuEej3sUHjqeFyoe56W0q
H7DSPavTNF0SqRh0GKGP5w4IfqrKfZflcYHsMwfAhAxcV5cN+pC99YplzQViShh/
ABWfG7SSwzAf5we864UVwcrWOOOPhmFROiE2YRi3gS73Pru9QXiwSPSA3NDzzqBl
q8KTNBSutlDWjjTiHtmYPlzv1NmjbNmTW48doGnwK6aFejBMLJKXXAZrxE2SQUPN
qzTWhHktbPskqAM3uAyykXRheb2fR/tOUAjqr2HfolU44csgSbjVBFFpDVJq6Wes
1VzXc2D87eiFv154S4Ofl709kEVX6GpvJXWc6T4rBAuoro3yEfsT12zt2a3DdaPi
P8iw/puouhIvOe/zmXqCh3EYSpQGNyMiNjknvTXVQQm1vseMOI7EcEKvgkaXdX2y
2oGNEjIIJYl/Q8xzgensKSNmN9x2ciMlOMF12GLX1b3jrKxyolMZLJVSmJCA5Fn8
JJkQq1PnA86mWRITpbvQUhAPJHHMgVVZcfj+ISmvejQXibLgyw8BiB/qOE+BsoGx
LZ1Z2p0r7S60Hv05nIABnHLqw6X51AJmrHyhHJ+jGakCw91C926OV5nujl/dQHcM
GHjwqBNUQv6aifRiGlTUnqcaRkBPMG83UBjE5OL7xRDSTH/RER61lguqvt25pAPX
sSyvLgiaZRCsV2zvYDVrguO25h0fVatWThBcbt1IP2MnkzTkvT8AioMNS/VTzA+f
zwh4tTRiNxx+K7uc/6L4gVEsBuObFhVIHpQ2Gt/sKpoT8ttf30FCJ3GI/1B7c380
RiBxwBlXMmoIA3GpXGa5zMG8zm/+QfpR670fN7fu0hPtIx7sfM+Ut0N69vK2mL12
oyPJpG/dUcOQi3Pqf9+9tr4BaTjOnobEDxDezyZIcDnPP+OC66bkoMZAVm3vl+bm
wZ8qiN3kxc2SfYJtSyvGggEFJGf1xG1BSJNAIRAg79z/LbM1C9f4YkSiIcLRL758
MTET2DCmHzD9AZ7QpCJ+lhCsGFIQDlesfOElfmG4ggytpihCm779b9tr1icID5Aq
IEv0Jsnf7ifJ/iu2tIk/JvkR5rGxxMzKbfX24QTXUPpXY8De8QO5mCmkiePXqt5y
To/i1C/jSgwm7dXrSJnezrL+ICK/L/+KSA9VQqCYlF0Ttj9GGNrqhQdpkB5bsaza
tnqjhu4SD5rOZhPPLAmepQ2JvYd8SPFhZYCYMSEgHJHR25u/hTs1vQFPyjDgF1SD
qeQN99MFtvBT2emkU6RVjoMjclr9CCnkUq6dWwTUSOI9dlfnb7BRMYbWziHtMtMY
SCV6nx7U/sIZ8yG4eNsFi9IVVlaXWTgd/erkVZRGw12ldqiuDD7GOhL+yLKqoDpN
v7ZevN2KcQmOW0N8MqkzbHCI65n5qh6Ri7lZ8vRbx5OsNQkE8G+D9UzKp0tRs8Nn
KgoABi2k628zID5LDxFZ8S9hOPW4JeuXDhn4aIkolQiY39pdG9a7zv0sqQftZvsv
iUH8/eP6Kz7whhspPjmyKRoNm7eW+jOTOi94qt8Csjk0Ql9YBgCKC+wAnotHMEjL
Rmvojj3sCxVjyhliwdErUdFJBNJn/9VQ2GcRnAqQbP/No0x/2tpcX8jersVpaFO/
2japp4eyqd3TWq2rMPTSVYVTnM9qAL2MNtJ+CmxbpmRcLIlOg9GC2dCVqF3esWRI
8wGbr0ZnQO21RRg/IUU2dPLVsFXzNiu9Uapg9Ya2to2wcrzXRn8LqGVqCfVJp1xP
1WaePZb2UXz6RFMkqwwT/7NoIvyUVjpXKVVUnDvYvGUV4y3X1umtqI2BKPzHbQCB
OsJcsB6/DQmntNjfssT43HRMwJzeAhna2qED6QbNVe3U00FrzXLUowALxK+sA/bc
YYgg3N/G/zOS7Ncl9qFbTLCVmfqT48AJw2c8PJYgUnMFsOg90U9kMoCQlbMyGku6
t0BacbL3c607M8TjDDVCmjphIt0yLDUf6A0pj1BoyovgiBXrievfL+6Y5cy36d+m
RUIsVwIFD3yLhyLdbPeSHVWX9L7Ssi7eDcouRNePleTkp8diRmxdygJ0U/8Gi0d0
XPhn4tm7iZpyX8zGc44mBVytsNVmpNEd+aQRfhzbsk7HPtg/QjgNEZ/9zmedG0Mw
I4P/NPu/KNT13YGaT6IYWbR+AHPFGRIucx4pshTH3n2eMOjKQOcHbb3JAdnh0y6q
E+B8zUbJ6BleU1bRR6CGR/uIjY7ITzTcNClPROrcFGC3Wum/UIwap7yvUXpWAaRV
P3cx8N36jWtuPBJ3zFwK7w3kO9LbqyV5/7CBkGExLx1XfQ7JYd8PT9a86QSsOMd1
DInNLHCylyskNsvsabe2KRT81MGsBaWMBZF+3Cc6UEV7QpeBCeLxpRcvZbUKLIf6
UMqzQ4dcNQ7H1BrXrg8Qcj9hQ4jDUEZF5wiofwHHpSA6cqF5n/erZ72Db15ee5EL
uqKJTzgGTQLM7hiIv84MRkjHEMjt6p3xmJEvHRIKpP+mdkBobcPOlP1JWeANG68x
0L+Xh+ImkWZ0FzZgvqlblBNlHiaAhSs6AoRbXmmlnCvff+q0NqPXMAIOxq+oPUF6
W1GCrambjkwVGnH1j6CTDzlndYQyXyQx0Y1KW18SMgNCCtpALYmEy/kSKYGSP+OC
tVYp9x3XZpJw4G+g7QYxuzBaVOkPEQ5pp4Bj+A5aPQo3Rhw8K02liC+vwmCqdqpp
nnpd867eg+TH2QUuAJY4DhW1qnn759VCf1QQfRd37AwL/kmMFXDlUIsLjQy6A4hZ
JEGL26K4Cka3IzUbtQ24wKiPLtavI5poVey+lVN8tG9AMI8YENc7fhglOlHRJohB
zvnDmBz91mUqIA0/S8xZqlyJqfovy7EBuvLmjsP48IZzkbJgaVLwSG3+5egWcRH0
KTgAzm+MZP9PB2r7PGwN1rXbKnzVY+YOu2LA/XnNT2bkdgiyl4BknCxyJq6gaypP
t5WXmm3MLxtnwls/Kgog6Neya8CRj5BowD0cI7H74GsXjRCb6w7p+JmuHEsbivYN
K5hYa/9vPRSwnsQOFyG7DxVuqMCKUyFeOkL8e7WxB4kvKf5XyBzcNgdHAZHDgMzt
4jiLgooLQl0dxx07jXLmUxwRP4YExEEEfEcVmmnTYVTgYGyqVtYR2ey/S/3Lf16F
uDiPSPjtliSH60GhNeCcbe0QYc9jEx1Xqe8LijaqnVLGLvz93JxxbcbeT/AmQCNw
TyBn4cSAwTHa5IDbjNY3jevkDPXUu+rLP4rdxmzo7vHezFOj8AYfLm/xovY0ZNln
lJOMJI21V/llTRFI+7Q3umV0kgIcNAvMOLfkOpqjoLxssFRFgGgdjvdgSurgJT6N
rjMyyFFuVDaJyc4UofqO78bDIXsZ6V8jlR30aKr8O7jWoJkvB4vtLEsLnhgQYJQj
0WCUI+V/jJ5y0HVUmy9somXIE3jMVNtnqyNN6wkXlD/GJHavfY5cXayFrr5I4i8a
Zrk86IpmYHU3sLvL450G9p72b1nI/LBenvh451KsYq/51w5xTrMUfdqiKx3Ks0hh
jtcH4+DDrBrsI9hI2L+vFCNUGDEUx3ZTDVBuQzJYNj+JtdaxwWrK3xJkAY8stxZV
1sR2dQ1KPasWKouLrrJiGHNUDnCFpd28Qk3WR+EcG7A8NoZJ34XO7owxXcpGudMI
RbUNbQIO9qFdgzTePKZC0D9iN3KuDirgoVnZY2jQQAvcdioWhnG/CRg/X/9X9rBl
qPmBAf2FUfNemz+23bfHA1iHwh837ALJp7OXSfCK99xTGwLLXWkX+MBHmpScIuM3
2vrYKGUf9MyBnrkgffDJ4ln12DsU0LHk2QoY2ilds6nj5sRXyCVVHX4/x+a6PlfJ
IYVmkYnKPNRogYyuF8vshQQhXDhSZBLIFQzSW8+eHtacZzEDoJpWClSaOuBrp+Qh
4+Gy64ovlnUmmJcuG+uYoyc2R2tVhK3nUyhtaPPGjbAHIoY1EdxHcMrkxUasSRR/
M3CNg9CrWR86cnc1LGJVeTyn5O3K5xPL2xm/2cMiAi+gDzkiPz+wrz+pBLSf15mS
2LDUY0zNMhS/8Ct/IKCM1LaaIAgiDP21CoN4xDlWHrQzqgt2iuu6pVzGXfpYGOth
VQ2ODhSO2BpNJ/BXgmlaOsirD7VQ5uhb2MVjDHOgA94LmbpS642Ek8b94qTxPCvj
aUgtb5apHk5eGIgDxhhONZjke7klreO8caCTHHueU4jD8DGQpJPMqBwG3QAxN56N
C41gsCoJz7CTcPuWsKWIpKEHTjpHGe1yPQIQqaMyk/mmNu4e9amBvG4SkGZbJZ2J
NCXWBkEJwhUBP8BGnD7C2k6s0IHlFd0cRHuf+/Ni9X6m7apDWn6pwDqy8MT3KhNX
tRRHQ/u3mEep9KdvbtN7ZtDrSRVLUGKG81l3MUWd0lMxfj+UIyauG4dyk6QOBQN3
JSLtXU7nsVOMCLshCLyQ57+9YGlMxgLOt2Mnwkk5h1Tu0bfnXOhjiVAyJ+VcnMvG
5wtgeYSY46hU70KVFBg+yPjncV59LNnC39d94oPbSAa7+/IEVK3W/akIvgWiuu+R
dQ7fyZr0c2astcXYF9gDSxTmLBLvbgtL0QBKrYc+QNusJATPzSpIQ7UrUoQk9WZk
qlfLfhFIB9OUeCyGQY5dcnk7QGmDCgJwd5d5XJWzzeARlLHGesL+HqL0CaRtML6s
xyFnfZaSfDVd0BnNCbq4nDNWK7DYG64jDQXoE2LYu0q/fUJqACEi0juIHgRJ/Qer
6nqw71RWy3Ex3KsAHFd/TZvCaOgeTagXu2RC6K+Se6oY3wBiRkx5pOR1J4WakHZb
lfZgVSev1qHHY/31G3r8HqGR791D8/PWaC2QGP5xG7J+FUzRYeCuO84H3EioCCd/
8UwT2p9Dr7JkuCCAqo1DDdcluyfG5nGuLiMXLFEgmao+ajt4KYoCaQZkTRWWc7lM
+91/cS6CMz16w7U/VatOeCDWW0ujKNXOfvJyLDceg+euYQd3LIfxe6mF3Q+UEy5/
DFQH5Eq5yQPoB85vM5qm6GkQTvjCYRf15ClZiDhiqQWgh2UZEUgYFayI2m50nGTO
nLnoEb7Ij5t2YSgIHcXl1v/yWDBR6sHKh4LV4YXu1lcHUG+p2QPH41t+7HXybfyR
oLtfbj6uk0bIQ1EiJ8xeuDwD1WY7Ol+R6avIy9zDPgBGeKZ6WBpLBLGi5VAgiNPF
gd0rQw4Ajl8oMi2QH8NVHIbvs0x6cHQNUD9VeKNqYhBqGhpq5xbK0HEv1U2z5qVh
bxffPhgFAjyqmarLjo2iLKB5wS6H8U3EVv4XwEQGfilSsWxmt+nNkH5CTDpH1IGp
os73Sm8Z2ctbKRaW4qYBPafmVb5uW2FsT+u17j4XDYlHZ6R/DqKgH8K71WXsVlEH
pNaZxDQ+1wW73pYWmG9hm8JigHveVknx2Ee6Pm8+iYLc+bmwKIHJRLMA6WcVwU3t
MKL6k4oJbYSXS1L11Y5JIPiRE4sFmT979XoC8SkIvNDIYcIj4tv+qmviNSSNTS58
KQd6kp6L1U18qnjsael2TWCqGwvTr1UVNO3ulGR9Uz3y/UFRM9g3dsJwX58IAddA
er2FiTokuTSn1KptDX36MQFeBrRf3ARemuFUNReG5n1etgfgs4I0TiK9IlT3HKpO
eSPZaK1NoOx5rNCoz5j45MokbeX+pLu1DsGjA5lafkfOgKW6yL6WDP9cdEAARphQ
d0eyr6pne33zvObXsUP0OBaRa5nkPwA9vZG4FkIHSGaszqvyWjp/Wz3nYOcleuka
0fwHeZ4+u89gobRzgXruvgr+iTRnkYVALji7Tr9xut9f+ezxFG7srz6u8c7eWHZs
3HVtu37N1hEuq1lBUQzDyqfFuxw/1xAf3hct7U72JshJi5o8mPUL4b6Fow/Fu2p6
g4sCQtR7BjHm46HhPi+DNFGzDC1azO1ACVaXrSd/3DXQGEhSljAjrsjD96n+wZjg
ppZ/Tp6FOtaiciH940FutXwbQxoGmGusa0Iej9AdvCOOZyNywD4ITg964SUgF8im
QKjTDc2JeVEX5C511ETK1yffYevl57s5I+0LvvoJjy4qbzCHROybHC3Xaafl8mG9
eEiKb20ymWfS+NBWKJSqNiOYniHgA/wNbGWoEFDDAB0mm5KTaqU3ZN7dwVKb3Fzz
VcJ3IkGoZg3Md7F1+a2Lar6GCx/vmU2r3a5w24qIB7a99ZYPJ6c+yx9tY1Qx8jpe
ASNNDyYQ7iq+N9spaHJcMsM2iF+5JqvMxlk8zvoLsKfCO7aWk0fWvRe83RBCFVsT
skZJ5Sfpp9U/8Oi7M2Luu/oLWT/nTyvclu+CUO9gKfTV1O21NJDhLSQxJPTPZGej
BefVfQ6MKavCuB/uKi28gESvATQDRYs3kHGPPxGqMIoAXQP49ZrnaOvBiX231xv1
j1UbsXqJo5+AM+ejqVj57UfzErgyQ8b577LD5eR5bpzvjITZjjCAB8IJm7wNTbSO
zzAj2zNJ7OP0YEsU/0/omrI0AjM7yKMykhfgVmzJ7ghs/tHFWe0mNd7mmb3Frr6I
GRFqV1YsgUu94sg/GkV9tPovzlVqxATSXzE3gUt7xXnq027b4wNPgH12ZZ6aGoZA
miSL7zu4aM6Idjb51tySfrH2M908oi86s/u7IGuXrnuzslQbgphSXYhR5WyF28KG
8g7bG6ni+muQLhN96r4YQyAv3gw8JgItrnbW5ymEwDl7oZKDOAIZuKDk8w1Lxr3w
FuGnQS+RwZsxj5KqByBY1LiwdHBiqAHLqiofsCFwh5cs+RQ5J0BDFnm+2CYPq6Zv
s1ju1aYfdPO5IWI2tfjW4JVsUy/VSpw6g+f27fu69DCAYqNNvKPzzyfTYVTyVNAY
aDBhP3x0c3xqZuxJxUWIiNcIJ1ehbvMcPCFHpQ75/a7foVId8QkIwJQY4qhb/X/M
orxWS2PKLm2760XibyTg+4Dm7ePlepSRbLWaAY123v4wjY5nwp8ntGTvQNr8I8CG
+LtPfdPB4/TdUyckUNMBiQhQ0NfeizeGU9uqvO0h60q29uGJX2Phg3oE83B/X3L6
oFU3n6j0D4kNTViS+S+z+BS8mJoYJo3FpefrlaiWrUpR5DTypd89ZEkXhsqO7DHX
UAVAPQTa6XP+wHEwall1tZYHhUzRa6E0SRbSAMYokSsc9O5q0BjllavEXlOgYt6c
1LoDiKTleZE39ZA7EcPu6/sADlzSrJVtmX7lTIdrun8Gvhy5Ely+4HMC6x0H2KXH
isJpLU4bJWh0RI+mmwA4hdkHO93NcKRZgGUWNAMG4O2XZ2Q/aB+pNlQEXj4Id04V
az7Nfn41hFMXZ2BeNfB1lvTvrD8pieH3C6Yto4dNxzStz1NydKV9+rDVRHlZ+TdO
0p3XXn/hOmeXJaghTmND00RkWuIn9ytaiZ9TzYVSmK2PMJUOQvoJsRlaZ7O2cdvl
q0upLb8Pvl8CACnTbNmlGaAwDiUM29grzskWdtbzrhOGw1r2XMRSejkIDA+rj8br
YG49OVxONtBGuiiCLdjIEvFG9EsmeKD5DDMzut2Az1JmlVTtMtXBFWJbqUrcCXq1
uM1TwV07O6yTn3i3GpZKMoznDzl5/BNfxXd354p0U0921L88J+KdifJ8Sak5Xl2O
9LKe8Wxy8vDIHWtOL1o9YRy+5WLvgbPWkobVSWBt7NBZ+AN4VGF9gkPZxm6e5hLT
8Hki5yLbpHJ92F3N1y95zm2FG++fcmiuPPCV2D3xmzkFQNxY8PjlP0ZXfxZdDP6T
9YyomFPdmb6SQryfOFw48cbGr/vSsbOTJqwxRIByYscsaGyfdS2CuAE35lJSFg90
aJFyEsCNEMqx14tNVz1nGXXqMjLzSSt/G4bgRpxERmUctOS7wuHz0nT6WyQxdNkj
9ySE3ULGc8pWuQK9rg3JBntG0zsTKZBAjh+SBVVwDMuJqfUDFzOvm6jACkRBrXbG
SP+b86JXpNfZcABKAwvBkAcL6UpxzeMVR35458/RQbh+MT1bVuy/LSThi82ZEL44
RklSxm5NN2THGuq8Tw7g/K377c14VfALjDUFHUI+UppmaIz4VocYXsveX6UQVgO7
bR0Nzpii64XisoAjI1NRwOqpMmyGuiHmsyyoV4u2X8VaU/r5ysLQ0UJjxqpxDZTV
8FSeWaubP69nXwdt2K4I5kTRAgf8jFhAaOK3GvnlO7HwVwnMn7ZU0/iBY9tV9RE7
FhFe10wccM6/WIWNypgmVHPYHkztF90c18bPt1+QflSI1Y51cM7mKOTYG6lSTSeG
LQN0iGGexnCL9HTjR1+F3VgbKI/toLgVn2/rGgBNNE3SLEbp6yAbVoEc96ozBbyc
rynkrCBAM3RgIOHfDEhYiybzJotqt/BKuRhAtWrdNak0AeWhNoMCCW6PwMVVX9tS
tUYVSnSKgUs6igJN9eWIGigQqMWNgSzPNNxJnmTByGU7a2hbxUrB0tlqro4s/Oof
BIELEGCA5kPagozbQFX+nUIz2SADToG+9349H2bbYDkmcDPsL7scqHkgRZZn8QKo
2xVXdSVMmh01IBOVqAd8EtL4TanO76s4UGArlbw3NMtuHXDF+xWlnSDYsN0gXEZ2
AVAdTMRrwaQZdRnGpnnvNFI9OG9xMScO/CecK2cp9fR6QNZSQ2h9/ts+mi9FLNiq
reXrlmGDG0ZVKt/p0LD2ZF96Zr8atUeATi0gM0Tx4BetlTqigCe5JNKY0NZmbQDZ
Ps5oP2SfLSLNry3SQlN2LM0e8oePSbqttJp+oI6yIAUqZJn6gnLbMI/9HsG2Ceqm
9aYVi/B+oTa5rjtHEXvGwcYdjDB1X7QOm/5bOv5NUGBIAw2K/ak/QBBRHr6ZODSN
NYlnAOKf8q8/fMsL0Sk+oG9Pnius6NM0ps7TIHUDxGKKtQXuWegDhFyYe7L3pu2c
oMEvorI6goL2RNbjaKpPFIkPeA15zRFta0qgdQV4jDgjGV1BdHVK+DKZfv2FaV3A
URySuakGmwKPqEz2HNricbqTFJwERbVyG7HLiwQl0Mh408eVa2iWhdH+f8ksBLzz
PFqZ2MxAWZG8ppV0qPRS63e7jqZGwaIMWEzFjRRRlyRr5swJ2rBJlR3Z1Qdjea5k
XDFiT5Pp7eGTcNsbU/KAcUq58tYNUjV3T6ch78fbFvIonxLlQbKJehYW37Rd2OUr
i97EP149pRx4H8ji6C/mKo7TJJQmLxChMmm9xc0EqG3dDfEwX8X+/ydKts057kaF
XV4UeQgINfhhVBsH7vvnCKSq8KN7bZ5+tNvLx2vedIxoHorhjq2fFRQfCSmvg1r/
F2FmqL/qgI3YOj+LzreGGn27y7RT8VwDqSdfMNLu2OkSUO+6/ypFfeM9/m4+7b0I
KGps946UxcDy5Qd1ka5vQeKPCJtffBfnU7EchRr/qGKF2ty6xFkM03+H4SwrjJK4
ClfybpgCrXd1e+fFUN0+KnBAqjvR+4OSjQf8wUgYOFQLC9IGf0xxRZPdvFT0LRA7
UrPS4EXeNJulnhbPmjR0PDK8A5DRcS0S06P35vAvM6k34eA5r3TYO7bhc6iXhp0X
S4Rk+xAKG345ajua193ApoekjFFLTfGfO5qHwpdCEGCyRX6torxMDKifmCDBYnTf
S/ZjECIMgl/IbO2DvKeiaBy0xbeQsIo47KIYF+XvNOEPGGC/DhJpS+MOQrErFx89
p0oc4woOmHXvE782H/0pWWsxCBTadNU15q9msvc7J3d6IEeHgeLYp+ZQugo/e/Zv
3Tkxxkk8YfznhsJ5+CgjkoAHtahQsmOobx1TSssXpsavHEaIeKurNeiW6KvH/eou
okKEFCGFw0zF7xET6sTS48r1j+fZvfFzwQKRMpjjJaMT8LFOcyWHtI8agsDjVUMO
O291masAMSkBibHTTOMv0Mxfd6CAaXg3s03f+SHwq/RfF5uzP0Wk4h+xO8OET/II
hcOqwzgTWtxcs67DEIk3hzeN2i27Vm8jiB8IjYtH/wXPC3DdSOzJNBJ46wTIU0eD
bBfr+fUlGjR8F6fUrvczx73D5+F8y9CvOSG8haTpu3OMYWL9xKzhZ83op6gKcEeZ
2eVojKYxJqsD3DxdFtyw0PzEUUIIIXf5mARswRLJRvGJgIHQZfKJXUkc3p6LtnU5
773TdkZGPWcxEWKmBc6dFFf5W6P9RYhM5/gETEjWZvaA1Pt59Gzm7pY9zQ0l6l93
DMwtl2cP6P2nAIkbuOeU8fDSCU0z2zbB+VXOM31oGekMpnYzcXDtQ8g7LCyquxG1
XRNnq+TcSoJ8UGMP4GBox6sXuVWSnW7/iCr1Hll4/Mv+r1QU65COCkDvjwjhCQYU
EyUhpvtTJcKvunYKrymypY3w3XXZxQArxmDMtLTMqnWcKh9OxzZKZlXBb4He8qVh
j14HMlv8kLCVE3pU7CwAd+v7BfuAtnMmD3KLCOfsiaIi8PVvlKOpV0kqCQVTpCqv
9Sbx84I0ht6SqbfN9+G3JNvYLZ1u0GMiA3woseWFc/w0xlCZl2J8YSQwjA1xSy19
L1tiU8jDuPeOblOEp9xMih8hdiz/KqsPz/3HoX6e/wrqmI7QGzTjf40ZzlntNnUc
b0ALBf0N7ZqME6aVu0eqKkxUsEjLp80yA9PoMy4kuFKRyuVW3r8KqwmCArf2fip3
R2n0WBnyS/ZUuRpnVIJ9fCkcDCdsrgLW5ZQOj9pOVcBRU91czbwgpygl4rbh5TXA
nH/kexVKdJvfQ+zdCr/X9aQOSqXsrZRkewgfYg+nbY2/Wp4ekOoydDM2M2+rGU7R
WatC9nVcbeaJvMSALS0bIxnsFwi79bLtedt1Rv31HziI6wQ0iso48x0b6U8JEO+O
ukvZlGRp8XzSKj/NnH6qu+gW9y7gJP59tKzER7Tl9N2kyq0dHlgK255MIYPnyu1m
k2B5oHKtcvRUzZeAP+7fzCIYc2AyOmUus921gjguddYASEEiwlZ5xjdKjz7faE5Z
OYjVYVam+hYZF9AW0tkyWqicKdyyMATO7i7aEUvB1oxuxKhLFqdoRaQZ1gclUxjm
dTVrUXCkxpoAaZIAhn+zL6VRqdSesszrIDUl9nlwNlK9q+Xtg1uUReEI1in3NSqv
qIa93E9pCwKzZtQZ2gU0YR0gUx1CDw2wajqRzjq5zfZVvClwQja1jpT89PGa5IJ8
A76CMNLi4YMiJUV+K4VtDBQz+jlurtsIRODUxkA/1KaP5ItxfSp0aD1FUqABdINA
1HydmWjZWrsJnAGgrwxKTkt0oEyema6pLHoPvMCJ7XFBHkulIS6cvk3FaztEt2+r
L62o0EBaCPjC0Zc10w+262fzfio0/L/e7sEPFOzM7AhHhF1wGXSYoozi9a20KyYr
Omt1N+pWC9bl3ytg4Wv506bQ2WSE0MLqzgGl8/xmo+OTNR9qf+kkscXCFhytfvcx
55o1tlUnoW9ujTfCCZYtRC2qdxwTEWr2vDUHZ1GX0DYMU+JuAfAeZ9IALQzfsimD
Z7qKLIJB2jKANmf629eC4FCox/5uDmZVjREOfKB05kPFLZxD7BPJR6RgkvfyMmmp
lzTdVfTcMUGHxV+9SKJqXw3H3ZyGd6CEOzSZ85a9bZXenEthc+tge/J2UK7CLASR
7r5HbXUpOwU5LyBtij/Qso+tDmxV5gk5odyYndxxAxAGSJFFd7p8jsWbopWNFjiG
4MHhfspQqvstliDKQ3fE5ev6wMsOqsqc08jKq9frCL5stv3XQ9xk/ANmrHePbHEv
8e9KG4qRTb6My8emS47skoNm+EhLEM0De/hx2gbUaEabj9bg3WGct0dx3DqZtTSf
w6H3BVj9E6hm5DsjThUxhcDsUAkfiDUsTuYRNeqSNeNzztJh70C5IbG1LEbL3gAl
QMdAikHf69nmc5lDslkJh4XcyNwthQvAvXQibzBk9YzFoVXu0x6hHJY3dK5Xkp0y
lRq3QelDiUUqOKXUPUAJ+C+DSxHEjBXshI5eLQpDrMYV66fOXSkP9XKaPLKwj7gl
P05HLtHMb2NWBgKGvhj/CMDXxC1g/F3jQmrn5pwyt/86+86t/wcSeZwkhQA0psX6
+5ltG51JSvDgsGWBH4FADZyVJSmTryo9VYUxuJkMgMi6fLBdpS7o5XsY2odRYJ3S
QpMBYfNsAX+mu3/i4EKr9H+8CeAnbDbzas4NlqswGRIHdKFfH/oX9aFIYCLkMZ5j
gMIC4VYSOWfGTSPOLgXYx+ogyAaIqW0Uct677QNm4JNz9tIvuVAQu0Y8OpZFzcQa
hcxwMZN9RRw/wxaqf58UWFMXeMp0aqUNkhKfGbRLEfiBLLjlVVBlrRpscL4x14cu
47PVB19/AVCWruv2Ta6AriOPeWUyB+5inTsvGNK6QQrc8y4T2MB1LiYUH9MGoClw
jPxveJEUHmQBGIXIzLRUVmrtWAj/tnnan45uWZgGUpodYk9+fgSiLvrx7sL24S5Q
IDAOtljoo/nvnOdJO4eFkFla90lYo2wsCIxdpv5hgTYDrss4y7PvXAkCrI+OuVBN
oZIfnQkOQFyjBpWBSG5uGUUqCeur5u2Nb0wRSAIcHROe12tg5v6tw/NBCAf7iIod
lAY5wbHD7wQ1dRPAYCb0CVpBg7w/mnm8WJg0y0O3rNMxOgrA8+ymSYtXQgHxu9cq
xHalWZxvEIWi7hABBk6pEVD6g5tIfIe6qfHy3ZAJMCHK1d3jj7mQDZ0JDOK9FcaZ
kdy8Sb/WwsmlemXuJDZzZVxYGHs122axSUahIsszqiWsRCWG/z3lCyUtRR2KXGGD
sHwcmYq3+XHFoYthTHX5/cPnfTL7p/W54sAoabld8kFJKfEca7DJ1kdhSyEegXUk
dXHBZ77gQYygf6HLtJATFjAIKhnO57DCmVugrpoMZcGRQQ2NmMWer5EVYG7Kvn7O
Y/p562S13B4y+N1Zpsku9PsNcJtES+/bMxvmkVTd+L5uBtHS2sLba5GtUhPMCZCO
kUOAQ/Nrp2ZqE8Ww4Vi9sN0SvCsiwz6WGPRHoGTlyc/oXe+FyZ68kE7cTnirIM+g
IHH9IthzVGoDssnrd9hPz0qpGjjC2Qvq9PKYdSFpvzNQQ9WUVALLRrM+8SuG92H4
2ms53+/rL+UQo7LmIH0jYmZQq20rPWL/6fVzPjXgcIPdyZNe2FgsQoXHanE2xoKJ
k8/Y+r34Kf4KwxLytuhqpS/p7Eb6+kMft8OM6bmvh9T97ynB5YyEkk8x1PTnPeYE
BxUTtzE7ktWYkj8okG2Ds7Xku+QtDtFUHexKSbMcYobOKyPqpPxyhMCOhoJJAfwv
IhG09+AJlkhGA8T3ETIwAX8goL1bdOjSBr0kNikCqPj5hw30DEXlG8i+pXhXFoMA
YzBoFnHQscs581bMKmf3iwzGfeuIyMuyuqUUXtMtQ1j0+fxU3BPpLlOPC1Pi11h8
Bs0C1hSZsnYnDF+WicC9wS+z1h4JROK8VnFGHlC3gqcyJ0ZBDBfdfBraebDe8t3b
+/AgLxiliKszP65nJa0oQi7IGe5xCLtmhkNaMMR2OzJ96BVEzqURf8gOLouKmmGN
yTKxEFC/t/7G0UhrYgUDC8aMx95k8mQ4bF5DVROxhw8XVvZ/Xc0qGjEqZZSVs6Vr
r+lhWl79uJOCYt9LOaCpK+fQUbKB3ATdubHXVL04ReySHmwA9lVavFKdqNyqVROI
h9ctmLTvyspapj6IKAypnqQYNE6O2kwjX5gX3bxW9HU0kveEzF84JUpsJz3SXDtl
ZqY3pG1mzayzsbo9uStxfsANjJBRKOYy2/KlgzrNhYAK4Ep3LQ+D/lJH9mDX5awG
PfLKfqK5v1q6yPChEJxDySFjckFln1/lro4lYV2TKARI5v9UorUySBf5cyeYFN1O
xc2rGUqO/F6PVO9/iFTl6EJ5dFSefuKo2DKoI4bfgR1Re9gE2kMuvrygROr9tIfM
RJ0qB/ClPHVRo96sMUW4KmxRwgmhI7S1E8a5rf+1AGAhdm8ptVnQrVckmL8/o3hP
oU2RuIVfT9SxLek9FKp9Mss+injYhPBmzPWjaTOb9IcgMqPZOVfTv806oU+X6tA8
oas2ufVSvWZ037OBeZn6km3aARZaS7MQ1NC27vrzDaKFd6RAyJaweuCrh5FdTv/H
LHhUkolO7U8dVxwRYhNhI4v3MbGtq5i30eF5NqxoouPUeBJ5KGG8Hs6d+8QbZi9H
MsSFYfwXHCIYd8+QuKAtQIsV23gO6Iwfg4pGCewdT79La0O2bjJfcKKnZoS9/kbW
+fO4Iguj/+jJ1A1q3dRofW8gdEy2K+XCVZRWOusLFExzdSm3l16rzJ3HJ9724EKS
L8lQR3W9P2VoHJm3uTiNxJiKRfh45YRXtM4JBjHPiQe+Xz76LaUdksgCr+2O6Sgb
7jJIiWi5Y8pZ+hLacLelmNEOx30bc9a3qpWBpgOUqWcd+AImBpVJWEoWP1xeUa9r
EeqDxkA0Anqn1usWfeJDTcXVy1nv9WKG2AzErNw7icPlQnPziwOuXrruO+m4WZz3
rncadq6UuOmBa2WCIUaM/fWKueQTfT5xdktWRjX5OwdH1rXFzpJvCAP0WbPnXYiB
e8AA8yEcr0BH36n4B+VNXvAvDP7Mnz2g/11LkRi5TstYK5kxYleRUgS4+7/pC8NK
BvkrceOZX74xryqwUkXqPCTwTx09kQgestqvAP95ZU9PldRHM483omHICJybpIUJ
zWH40027+iBGWCr/LxwbxxuClscNlTwVMM1BJOXFPZIamuZC+32/9G+qWcoY8fF5
mIqYrz/VbsCatWxi45pdpHASNT2wh4wQkFA4/PaBleHhvRoBBlA5YvRfSyewmnvV
6B7ofvmwJfcmytuAYQxEk2yDlD7Zw2WJRv/u1G2LD+LBzlTaZlbAxtYkx2wA/uWu
ToU/eSAuZX7GyVi1jV7IQGI8sYZDLkDSmJ1vYPBroeoo35MuqhMGYVm/fzmzrPub
HX8J2CcC7BfC2L0xWrclpiJHQrZR8pLV+8LV93oWsSfBOT9YZnC+mW/zUHA7tYwL
VMvJW0IPwnJLshcLY/cF4lilPaihyPfv72IEYJYb7J+fof0Q4LlbV31z3izCbHm2
CeuyA3KXUjanVI+ErivzH7EK8NPfkiwJXmnUz8A0ji9++Bph72lUYUAM7+egx0Vp
nmZuIRdvF/aePwIG1ZfTAYv1n03J6gj/b4KHfUb5anQvQUEUDCCM9zsSSjxJFU+C
JRsa/irXneJOf2LP3C1aqtuWemcXqLGrU/6MauQh9+RWjWE5xhH1PYZpyLNjwJKE
jtlNyPHHIVXaDGRP3L2tTQg8MPyoCSSw196B+pp+VNJ8FMsLJ/xFTBD623ibvPpk
HTsI08o/beeTXbi4S1NaIOBDOmzBqLsR1C1Ex8XXN++SsG3DP8ZPFrzMIi7rkKvR
bV5Lcy5IVZYXACEU0PaKeJU23hkINMEfwvsr4WVJem+kKlJb2FNmc98jEtWXjbEg
W0w85K6HGJxSvbOpK50noIhcgRF4fDyFuzZkApTwMdq22ImA7uGZuUTKbe0giy45
uAMK8tdtSg+ZXSHk4lsqY3A10sNNR52q9DyoOlWb8e5OjIxoTgUVScpZHMVttnfz
TAQzvJoi5rAzM+3cwSg9GMQw4WtGtaZ41aRtoF9RkdHmIKD4LyNZcBwiHpY2IPzY
mv63pxamzgyzFIdDRuGnlrlRL/PAXRIqP+/m9ateL+IyZ6MVpt9ywJIRdQpn5rI4
bRdeC7UnIR7LAY+GVypHlQNbutavKDkaavoD4vah8nvs9qaYTcEfAdHAFAPZedXV
XyNm3VPkHZ2Iz1yGAIjVquHp1StFHz+0EC4mqmU/kS7Q6H4nH7+c2TLeZpRiV5mw
so9g77f5jKUEEjdz5XLTNp/DREQba95Rh78aJ2Skqin/QLoA6jHrevtm+YfbeLTh
dSK/KPWRBG9+2S4WdMj8OFSXEktnJeydggRtMJStWk7JD3ObQAVqTBDO2S78QizK
VbJcmptKuN8NCvMi/jY5h9thqcgDXBr1Fd5TxDFowx2CaEXJvzrcC9lSqnS3r0jx
v7ZyWhEQzwBZw6DRv2Nn1gKmCDVR7vpsLZtycDttdjY1/TMb9UqLUEhANZ8OPrEg
HYzhmo6U/jln9G7k++2K7pC4HiCNkRVAIJL568QovQi4QTJgX6BL4Qy2ZaYkHTmc
N57Dgdy0drtsQRzzsFpzNPoP8G9KZKy6VYfzwizzimdqDQFYPb5IGO5Tc/Pq6aHZ
jSH28xIew+l8gihF06IaiJZatKrlt8mKQaQ1FUYQ7F7EsW1RwS85OYsFUUmfa0yo
0tQ8zSkzX0wHDQ79IOjNEBmO+fvO8RDt8GtubNkny9zcWlOl/lBC4N3cqkABT7Ve
/iZngezLeqFXYAqafEiQsBJ4/5vWtPMsEGXq+h+aTEjvs5yXYe8Ce4xUIm6zQQhx
T0wxf1zvdo/fbiAnV+7NvX+sLL7NYyKH2KXBcFfS2RFuFbBAUxmV9XTQF8R3sPje
2gp1YWNMz/UMlOotvwJlwnK2KJjr02A0QusnFRvlXC4vrrRprGT1QVffYiK1Hs8T
V45o+HqjxCf3R4vAQluPOgRJQN+H8hYLy/4J74pVlQK3BB9u+fjQpRjrUcDkpaQb
gDJy48rlstaen6ZdJ2mS4+PlgCV5ZMiJXaE0ydkkFmx1iwfZTGOZoGsmd51OpesT
w1DS1qK5XYSsufM5t8jIeZkHGud9paxGsKpZUZ28Pld71UiOLM6gJ9vekychf3lr
YDSIvimvFr4/h63F6DBpU06YHd5aX7OrsQn9DgBBG+6r9IpS7NeblFjNvkLct779
woHMMu+USOiRmX67RGam5IFuhBLGvOAGW8Jq2Xw8F8n3uHWlB9wnf+Jg7QaGCorg
/j5Hzuj2aM6+EyAIl9XQF1zK+vf4KZdxrnegGYHu6ETpnxhzfBi1B9AHC2cvNOcr
tMQouE7A4LBaVLmE2hw4XxN9/UPuw3T7InO0Jz/exyVzDskB82F+e/Mzsy1uFLGh
o0ZIruGXcedxuBb4WRQ5GZdAT9MpRu1Qi7g+kjutye50j3Qdwlga3EjmkZHOJWBI
nx9xsLciFf/SBGiLdZHDW55nuk109HZNT++b6X8Q4F0u++B7pY/894uL/xUlJV5p
YscSSGRBM+6D2ijrnnskoO6YtNdntJ6C+n0+mJzF5Jue4PagTdS1Ub+qME8CdLfy
V5vFktxUHswNL3CKADM+lGO0OWJvGoDCc4ScYLzofgIZ8JVw51+NCkKC45DhYmuU
mj7OKgzb2vLTAPm8aqD+JjtByaVrSSG6JH4c4ycdGZkMuXZbcegbKFi9TCO6Fu8C
dismoQirWq2fyt9bQIazE3XJznc4zsdlXzOLxnTgCzPiFHXbqrPrDpkEeWq57l9R
MpnwrxoKTAGadvdiyn0nBvv7GeJEOaxNuqoTGMySPgxhgR55R3EeG4aTxq4wQUMi
iDQ358TPJiJyhhzQrvIQg05qbsLFVQGg+vaseTvVh+zafEm1YBVLxZPtXIEs7rYL
NM8mje664F+bUBKT2bFRQcy2hmbN+Va1P6o8UipaYowahZT8RtraaX3Sz+NcSDmW
O8SvO8MeMAAHsz6uRHFI223GxqZ85BRhUPKX7kkS43qBIAl+xvicmWQExCSdn0n8
xxqONm0wgFWpxbgON4G+To/DUSEvN4CmSODLPS9aCeCtNU8YhX4iylZnbk8QUxY2
WUj8lh0agjikdrZ73lza5m2e31KI1//qMWk+1v46snYCPPcMYtKmZr889qBZd5xo
JT2i6O+J/+TSRn1/AxifpmouOjd5ZXgtf2bTbs8CTZyUAGkw/DuKmG0LjZtBeCJc
sUaItd28rdjLwbsEs5vAnVFMmsEHdW7dnezkIdjhME9keUwc3zoYanv60LwzyQpm
W2YJQpZaeoSstVZt8fjNmGm38n2SLWth+1E2to2oBSVJKoPbuRZPf6JgfBXqE6Oo
1YwVHc0tWEefwUZPm+EE9zhilX6O/pfg2KM4LFOADaZRSJowkF0HUW3wjIPz0q+E
+hUef6idk/5uhb2/IN0iiHu7f8abEWR6ofOrfj2hz7mcut1mOnmHAaG61HdctVkE
GfmQIQ0ldh5BWIMhy3iuTlDaCVy8GpE1ApxhWQcjT17wzjs707yEp4cJRzyrywfT
XTOvLNZINnbsPIaAzoD4ENERoRGQ8PzDjEV0S4HG6doNw0/sA/AqykasKEjXURcH
78mP7Hmq1/p+m4wxlgqoeVu6LVEhr0Ftc3+Miya1Q/PfTXkHF8BW3sJ7ztQ3+pJU
G1b2RXpvMb58S0YeFpPCU5Ga1WK8c90KEWjp1FPSFGGa5g7vcU9R0LJakYcj+qhZ
z6EA+kfQf0XCY5FnuOInV8i9uT7io3kD1cpdsG9/j1TVYLPq5I2fcgN7ds4Ghr9g
P/XDch6ugzJwUqfHWkPUmLkFwflkxy27xOud8BQ/cQ1ztxCmYyAmgkTWoNuOGGLz
d8MeTrAPkkYJozsRpUlbt8npr/4rh1Pfny0574qM14788a4vwelCMExs2e93X8ii
FfKla3s/Yf3xMpdA4ewT3kVU6UNMLYeQyoX26KdKm+2PApB7ydO7MRSa1+jzLMfW
Qsce15JtoNatamBX6ff2ohK3Lw4hMmOXvi4hRp76EE0GLq+uMkjCwmTNVu7rteFR
05bTNh2jX+tTQyLnlkoNG7511eewf4vPel/k6yGuYcIl/DOXItiWPdh+Kobvyd3I
SDSd1tJT9zBr/niQjsR/9aoAr+6P7G9pqjsfZTUnAqye/rKxwb96Ql+Wbn8SpRnk
K7pbs/qO6NrtyqSeYDciH5G353ceXwspAuyYIO0cs2L4WWXRXw2+GnyH0RTwDl2K
0rDT+lKSrPgLc1Ltl9OddwgoSfwpIcv71SoOIG03HXRmEWTLx1IUs3N4AO+/bfJ3
Z0vrvqBbOuwX8uGHDOfD+TSBAutLhczB1NnDOEtk2aS02gUUJmaRvgbfjrrVY6D7
CQA0AGA40sptRy8h/4tQLcVFQzpuG2TrUyR6sgcbeFZTihNGzE9uCXoQamHEFYWd
+5PEBw53ebvg9v8HFK5x9fNDdA76uRoRxrwr0aepipFLHVvmn2K1U6ivwq2/h2y3
85/ZE0EfF+vWrZ1YQbM0Cci4Ca+2Vi4OY+mcvOLchiTB+LBF0QJFSrnDZvkWSVet
ZyFCX5/OsaLkGn+HTADlTNwlhpsDQ0tnpIwRKid6LSAHpHBfZdHqKat/rBXkw91s
fnWfio8YS1J21a5iqRVCBMMzBVXiB8VVVPXvYI741ZZdOc4ZJfyOzFfQx0mXC1+Z
in66frUWDPQ3CRsdCq2mRj4y4/RXqy9TEKaL+a6vuuNYbjptHZjgvR8QFGbMJ44v
VeErZwLv8P6+T/Z0JgWWmcWJot6Sl1XX/V3g70hH975YsuEzmI606ah+WGJXyvG2
dHK92e3MO+e+IEkn8isCkKsgCZi0TJAhMSjCGYr7uREAHO11GI7zjlIgYZNMaPm6
gZOkeAiKxIr4cfYuZJAbmGU6zwUbkp/Ga6qV4YgGaBBbEMq4Repx6myrGp+NYyeg
HciZR4viEUMFRnBWjmFvni6seiDgPM/RF0l4/faTlo/R43DN7Z/UjIATGBk85YhG
LQa816F2V2URA+PmBTsfW/SlkdKYKn7JRKg22PMXBC6ILWICNFVieR8+cvh9VRus
xnq0xoCzle4jIndnwQdBkKF7JoB453uK7ic3elS6tlFimeyCMjQ/i3RUKkWqxBB1
KuUUZj/J3L6WOjr/sbaAsiKBT3DRJf7fk1/cGeAv6rc76AAJFFoM/kS5WrUYWZaj
z05GvE5XneaFy7CEbyPuZVu1jkl2lZHIby7AeeOhtn3uxw1G8l4HDEt1mWJxbkUU
ZwrclTxmRY3vsWtrWRYGPWd/Yqop3nP6nNt/YYKxz1oLKF1Rwe4EmSSX0Dwp+8Bm
T70mf8cgmQD5pfBp4p/0g4gaN9SsuzhFLgTw98bJohgcoH9rWV60jJQCAflgZ7X2
9hW9SMCqSuW7sSXRWZl0zLAaCGszb2ddR3QV+GzdCPXEMIoPr27D6BjeRads1X66
HWGBTEGPrbE5oSqnfZDf/jQdG1ta1JX+p/SsSPbXpoN429MsQ9KrunJyKQ/xGsMJ
m7SbDhCfLpRee4b4vWETX6W7Yr/XU9EwENzvhJfSHOjDSHYc5i7PuA64k4N78iEP
0TCPEButzo0C3ZuEbXonj/Wjh5IzSNQ6mwg66/NK0oliqvWSj5dESQpPVGi+rKk5
6zPstivj2vc//UqaIDUU0eLFc6UZ9iPoNHRzDccP39LrUD4pMzCjuzttglRPH+0M
cp6YKEk/FgKkaZUGora3JDV1ivgoSjQIYVl4D1HY5QY+b8o74SL7Sa5SLjZANX9x
EUOpTx4CbjwVecDouf8Ts3axCyt2F1sgiNC7dM54y/PRwZ4fd+fOigu7uIvgLfG7
+FTGhXLeIsDkFQlKOSCZ/z6hJKKslwkNIuDCywR9LkVrFzr/23Z6GiCoU8iPn4XB
ND0inIlOP3myX4u5W5Kkp+sEXnCqjZsWQ9H626bTS8pI7DpzhIwasFAiFep7C3YZ
JokvyuqhhpwYryCu8YMUS3fDYPuAfieW+RE1FV06ybBG/NGBg0SARtIzm8bW54NP
CqZ/s8OO2ZkJpLnw7a8jdgZFoPvZFpfqQqXOg/X1udR4UVOsFaGJeM1vagbNzFI1
Et8dzum9fn2etQ7QQF24R8dMQIxJE1XPpoX0EZHurrmxJt3bomE6th/vcvL0yqzH
1N3tAUUgg39OhDBOw0wMeTmciElhpau1UcgjPAR2j0/xeVgKC+kb1+QebsnHKIEY
M4bI79DyadncDCxsGk6aaSnoNQ3pNKUsVj6GkY+4MwDwdqCvv/w7ancT9ZLiKoLZ
WqpG7qDhhUmPPQ9ruUPPhGb7zMOwyU/OoGn1P2gAwhNx4PvCny0pcmhVmoSN9jic
pDrLNNVkIDTH49m32UNLa4dybLXP02Xw3fu4F5IcpZCZR7gEfxtqIb92oqNo8SEY
LwvQS02vqvBWC2Zx3RBePqz60DfT4/aehlZ/gH3c9MnNDab3uj2B7ugFIIqyOpEo
cYTvHiVxbPpb8O5Gn55XW9F9J4puQwxYNz2AmcyGvknyDkuIHbsKSYIAjdJJnTSP
3yv0j/Z5H+LXzUc2zUIf48bBA8AwVQw1tGdf/U0ahvZzGNU6vpS84vQ1NCIo94P4
ru2BgJ8kH+LBcl1a7Hpy4dLjX7vcAI8D5q0nRn7YKncJWVJBoOQWWGR2sS8LlUTd
P2BjxS9xofUDNZ7oXBoG9AF+YbhGPqxXBU+jgVIjban4iEtxHQ1JbDV4xu1IMSwZ
nFvf8P4aVfd8xN4UNl6fI3rnoywAtrBW6HAbGEZcLKldnnToZNpDf97I67tIte2Z
ZF8rwvWQXpVaNCFChAbXgqOkfkx/Smfevnu5sXGGNRFo9OW3jaDURTUlpJE1WTIv
hVCc574EvknwMlID1KOu8mI90d94c2JuPFshAy+c0r5HzQgXmhfj8ANWR/NE+hLU
j1H5FpU38yUqJI6MHKlv37ooj5zJ1cSVoaA7F4WiKTyaudNbmDdQmH0z5V56lhwi
LFB7rmwmcSkwgW449r+ZOVlvhmgoj7+n7Fyzm47eksUX2gRBYR5Zq2loI5OMdQoK
eWCt1jtM1aTick2Ql7Yadd4YtohGzyV66D6fqNZr3yXvkZk24zlyl6mfpTDy8x14
gAnHrczQUAHhqE72/LPi2sA5PWqN8jmcrqOcMgb5aJRmkL+DglNpg/XjTlWJmlAF
owde5whFlOMP/PCQ0/eIvZJpOCrVAeoXKSdI3BgRPPTELq6cdyTdzEMs1pCd5BLb
g/VtQqhefOSUUqapMkToArTNnfacZTv158g+eN1U55xsV5kVHz0WStqfKhW+wDEn
iF/wivwWqr/Er8I4M+04tOBFx00UTgxgBUjc/PJlTo/st6DX0WtDy1SGFjpR0keO
o0DiRyPWxDYcgaLiFLyZXgfi++ekgsPjjWvog+n3J64rZ/jU8e6RNW4HR3F/nfU7
cvwivyUGjarVOlCk8rZ4FA0vwoUzxPkRbuOCsbx9r2Zfj5JtHRgouS2vEUG5MfE5
hcnJN+dXDLEWeTGNNfd+tppQ8zNjRlYF2dk3OB5agjjUvSJh4eUuAUPafltHHITV
usKWk88o/yamBAbUWcdShzTtKyvpsnIpj0goY1ga6U6YSHcR+pCR6SglLX8fwJqV
2wdGocvQguDpY7NYBcVLZc+dtTH8aPuUVAQ7wt3GbjCq4ULuCkqhifN9KJ/3nAus
krKQ9DhlNp/jf72C3PiESaZDc1bPqMELVur8fZNGELMrI9N+xm0GXDLYuiGE+qbq
wBimvJeVXNzmirLR3z8Fn+h9hSS0UV+v+cXRrqthBLZA6NRMIeAmJdwVad8d8zAh
lIqAX+bP7gVmJeOOW2IRyC13+Ub9iDeIm5UgQ32ZJgCHo6k3agAFz2/JVT3R7tor
o6UP+aTCDi9fiIpr0SDcKsm+KMEjacjsSgkyqBkMjcdoDSqh3jKmYczx5EvsndRV
pFdZ7shFXxkmbTnwuxu2V8C7Kx35ttHiLKg8qPEGQXiDOUoAFdhgGRSukM5vzS1N
+svOD19vHwj9JCkjaPuVA68SaYnssa/caBgi6C4YM7pV9swDu75wYeTccxbjVbiF
bVOFiu/nM7idIv+z2ux/lb1p1102NK3e3yBNDTGLtCoCkeFeTGPKaXkXCKXYAgS/
+D/iknRO56642G7BfhRaakR6K39sRJhOV4yYzGbVX/MBfRfzs+9MAXczrIrhqPxN
MHJjalF7Lr7V5/pmwDcZ/MxZzoZ//BGnv5R6aUi9PRre/0if09MOlKOsfB5J+2zE
eo2vm+LOYk4t5568RIIAEBnPihQRMHb4KkxThEH70gJQW/+TlzQVF+YqSkJmMOsr
f14XXRfB9Z11ICLF4P0xrfTqZ2+xygaH99D7MkEUG1/G93T+SbvfNRoJz73S27QC
DTP0jPPEC6+nSsJeWgSS4WYCtwaU4VBfSpaZ7fxqxJjtp8J4aoNx3Cn3O0sokQna
MSmUlFDDoytEXgQGROfXXJxKL1NH5R7w9Tmyb/h6qSJQEwa/bLCYqGVIvbmY7vRB
OCk58ZUu2+3mEEvSo4BUp+1EFpDpD6/BEWy7ewXlRw2z/pzjQUUFKoLUKfMe5vJc
j2JJKG3UXezy43yrHqzfhntYeG2p/tyXCF5ABu69tHyQlkfiHHfWB5KsJQIn5cNr
NdEr1Mq1+/c66sPy6X3JGcitHTXJI9C1gF17R7e28ZZ5WNrc02EEtebMZhCl0Y5t
YbqqSRr5yqBpLYROQC/HAofUaMIyww9v+KWTiL3HBLIGJM6fns2zemlKAMVHdd7+
O/uo4L81md66eXJoeUl8WJ+b1rK5iY/Sp3qTKbdAMPi0Rtuf1EkJSx+aTPYR2cHu
j4Yb6kGpFcOXu8PQGcm+2DNtjjfY06jV6MvDqTLNbHXf5nthd/2RsxiEp4hlIlmn
HFW0n9Q8746CI74ncgcu7HvKdlGedMpDR48zxaZEywYAkCfm23M4qpsCqv0bU3mV
EDLKd72u0PoInZwMViua7facCkFzP/qoQ/uGz5v47OJEGR6BegHXOQxPgpWWHdDG
x4hQup1FXvfGBu6QZZNCMmKU7MahlPLnkWmtKU2nUJM1iIKxp0eTRzD0w9n0Mw1r
gNVVGb2XUVsHUo9FB2+l6WO3TxeasoBX9HYlk5LgnLjljnWbgBdsjG6rZEkKcacx
84negKszt2Nn0sZ5JymJEYOV1CvXDhnLsiXtu8q4XryUmFn0sE352h6HZhSlMNol
yH9+xvE3N8j2M7VKIiAIprQ4cjDiQKFnlvTiXgOYdTY6jZ1S7ygChxg+miefkOx6
tEXo3KruzSSMgrmdjKLPD4jJZCX+XIvW/MGGaM1KQFW9qC+yTP8PGcr8vlAJESR6
JzM8It0ChoVSyIzQUbMPBOUKrUp7jdPZqPNfk3ucnMuCf+AaOGEiFUJdVaf2DAyA
eqZzltf/ws2UkKyp5ohNQtO0lXFDGcZGW5UGyZdoczKevjsNJOZZvCQ5tfFPIru2
XxY3OBBVQ3e/DRiRhYrNUgKNyLBfV3c2ccDETXspd2mzC5sg95TA3wNHdJ3Jg6Jf
jfe2o5S1TIXYGlmMvssIciTbrF8lLAIwFubSN/fm2eIVXH9q0O2oAogs224hWAXF
tzq4SCFgQT7Cm8AGfpIg0S0jfgTdNT31tvldwPKkxg8o2V9ZwcGp0w6oD0umDjpV
mO+JSdKhcVeuj1URxCXNXjQQAP/OeFyg6KcZSUf22FeA8StsF4vWfCDzwbaTyeh9
QDdmsSDKNB+o/gcnVFum6atpbFg0TqEMIg804bt/vLCTGzhI7qyH68uBwX8ovVZ+
BlICb6qnqchnqodM5MIhgfBcDdIHRyyidP1gNwZ6Gxf0x4kFfeMSDBa00qY3cTMo
2PUJsivmM+jWd+p4ZK/rGkEya/o5SZVFZLmzXowMF9KR35Z/aaXd4u/F5h117fP8
O26ks9jqY5ZQdGObpIONRn2sEJBN+0GKQLgvRkTfqbEfYjOTNgY/L41qqYOI5tAl
G4InVeptGjotwha/d1DT/Z/i9FRDxMZa+6IslApuhF7lWmb1fdVCGM7PfBwJ38sz
zg6jwzH4EKcrNENeDZVafE0ANDpNs+CgaiswOm/RAlNjTkmjA2dohqv7zUBVpz+v
h/BMBdqYXAmvmsVeRG9NL7M8U/g5Rf5qn5akSWKQ6SmkudVN6PgfeetvYhhObvEQ
OnGDbkKGVbJWTrccvcFT3Vt8HpHQTbQvGCRKDES3ob0JLMy6TBMi8hmMe1xuOkll
3oUfsnY1XNfGmB3DwZtAUw3OQO4VOmJHTXe/tGzyNBnm300dsbYwdRgg8AY2/53X
9QmArIPM0qDmjKJjBEgc/wuVwd95pwJmaCQPGHeghZnThSgFwUCUQn3rTqKSvUD8
uu3tugO3rQErgzOtgkEwbgU1iroztmRt90bg10urf4yoPKNVgFlXfd+WULR02cCT
w6SF/JCKS02K2midZnsxwEccN9NL5N/xyLda33eX3IEhzWJWYd0h3GvSUvssTBem
kQQ8AldTtZaAXbcmWkmZGeKk4fZsrieK5vsFvHwIaYe6bRvHi53PV5wx6nASP8KR
Keyrr7mIehbCymP1kgDhLnzXP9wyXJ0YgI5LX2DKd7cPceAxKFfzRmSSAfz/X/vx
JuIWK0CbSm68Ny3Xufr5lFs/LM+UETdtN0wMpnYKpPqJQisVm2QpkkJM2S2cgKfp
qaz6KTnZ4OYbHOnVt6vth5GH5o37RQ0zzBpqSe2dCalGlyg2ynm/YOPt41DGmDhl
BN1JXmQs9djZx2728XYakP5l0+VjonwvUCrMa909qs5321LF+lHF0r6Wn0HJpZhX
AQ1nRlz86M6RJ7XTjSk1hdifMIIuLNvitjHhUegDOotc7z46RHT3uZQ+qkw6guhH
rqv4DCH4eXmOujQzynk5jqaGbKMMVgECQrSeG6v4GahTXPs+/GNDkoepOZrnD3i7
cZl3LtGtR20gJVTMuLZ4BOy4GHnBb9V5mygGNS6T94keJuNrzAoUBB8HVAS/56vO
v3h0ElWax++hSQVXCnCAMDjwfUjYPo9wjR+fKxZUVXjQNfB2+JUYdDKqoHYqtpDJ
TeP+6BsPfHJ7P8WN8zo700kzDOFVBOJWlaGmEtVvRvVVfrZWHqvPrK6zjidmNMTl
CYkNtmIHtfVcKmVZoM8rDRvyBtaCVxg/b+GbF++xbqvNehMt/BwWIyx7HyiK2QRG
o0Ydz37E5Z1uD5i4PuH7SaMGjZq8GVMBr0+6r992+JmBer9SNrLSK+rM00pVj4p1
KuD2H+pUIgYgdISKkjE6IfGRgiXfPN2X78hA+jkcWay8dad6vMH4OycvquznA62H
yD63p3gNRHc7xLsukhAsMzBTh5nWRgrJrhgrnkrvoUOsinlFDIJyi0MXjILmIq+b
jpGUjrlXBas2/TaGkNcnEOq/yoJkVAUyMMFjAP3QEshErqu40c/S5NcsvnBNSuyl
Lay1rikjGb4nk9VnvgPa+402louB4euxbTP0P/VLConLw6JGdSVhdGZLwl3CYWZa
YRGAyNpvk5VRZ4Jo9ILhFbJyUOzP8RYVxaDqwShVDAmBjohHp09lWzap1jJZutip
L+xB8n/e0AmiZz5o/bUp87kqi8xDDWkVN48AvRvaFViwr1blkhjloooLQRuoRb1c
ld/ZXxEI89Ph2cZ/cqIBvchxjtn7iAYt1kKsL+1zfYqh9BLuHmm1V5+rNzcYTpWP
wxupep5DZ1YfKL+MayAjeLxCT6PYKsLZexgg5lF/w4BeT27/Vqr9UFaks6DrkC2k
zHaG67j6JcuAW9vRGgZtfvTTk7bb+I8uEbs9LNGC3NR+vw9443kK2R3TUHdKSJ3S
fXpseiytdwmzNsLt4fENh/g4cozxU8zIXZJxXPHhwcmSn/sTAYtd8n5ZXiyatFo1
KGi28MVjAeAw4aSbW8es8jWa7NCdKQ2GXY1j9C0cucsL6hU5iUxxOKIaL6LYpLoz
RLBN6YXOofqBIuIMaERCIq54Xa4vMJROW6rY4dR3e2XQDJQ1dDll63hD6JACmYZW
c0VQAJsavpFW9jw8M25RDZjKlaTUQeYHyzy0PT9suCJr5sNx+q8n6wtEN5DNna9K
bBZFu69VF4NSre89vSHGgHtuHUMUmfA/xearPT3BN0dsx5cRhbI2BjP4d2zlB175
6uHP1+GdaSnzQzoUdKBzfuAX+RzZmwT8l75Iobc2CL1JMHD80SrJSB6J6CMTWEkx
tc00l72EoapgFFr5/NBVWu6UaeFYjExVpBQ5xuO2ZtZS5Kz+Ags3ElakWBaK1kWv
U/JcEQQwEpYsmKu9LHbfFsGPui1krNXSzPne3VTEKgWZJd+kFJyvPRP+CbLVmxwD
UQaX//KDVM9B1610uXFMzPDvPUuhEM2R8YKnqrzoIa7UaKUSrZB3hyRYMJ6KR2Cs
Fwa+iIKwIwRiGbfgSMwoy7WmuAoC1l1Jg04YVrhSlxUWIHfkChtH1l7d+wjTO9hF
Yxi69mug+tyQJga16tmRVvKDNXFdvkF/cEg+syH7lIfkJILknH3J59841zfoaFD4
RnhASOBaZxyivpqSa54Ue+XBkT/pMO3Sd1OiQSxv2YFfFCZ7yLqrJN9JXB0yKOaV
sqxBezA+2IS9xSLsK/OhYmKETAz+XoxdM9Q0dsmdUZLfnWQSP29yNs6/yyhpFGzR
D7XG2pTUCO639tRH42iM5AeM+by93pIC8UUT5Kac8hOsF3Sb+GaBMgxZyKpff960
GT11pa7wN2TSNIK9c7o0n003qB2LiAqf/HO9Wk+HX7XI8j7+RJYwMGZgScRMlnEf
2cZK41qRSiPpSGEnq8zAkaWghw0QD8W0eo/UwPWV0VKzkjbW+A5QpFxga1+Z68wF
5S/IA46nv7yXmU6vLR3NqALmPw1FFb7dn4ks+gKDMFRznYK4Feyi0e4/7vNz+Y1B
sKCEvZGAUgsj7V2NTtUQX7inpPzyQas7h5+pw9M+uUw2cK//5P09hK+wIuanqR9K
DUL2HCH6vsEuxInOl5g89fNjfP3xg/GhkplpixeVbTWoef32qRTQGghMPg883F4y
IY5gdEQas3vqV3mWqDeWI3WFeUmXTnZdKzMsB+JbD27qDdwsVLousgwcG5PRqHWC
3m+EGyPCNsqAuxSjMY4P0803kbWli099/GFPc3UvXYNwdi7MKyeBdVsNCfnqoYfk
8zfxkXWXodMxYlpdq27XeMmqBtRYufpmSnbbp48/D7knukyTezs9zY3jCjGwvGvu
fAbhILDog1jGWe3Bab96QKX03TKWWLQeU0iosAbfXBROHXWiic8UQsJ7zLvDv+yt
e9p3ZEEUrn3osOKu43xa6OcHK9FhPvqp7WH1Sx3IfO93pzR35dXurqHmd8nCxIkQ
JbYN1v8zvGNxMIzgOPsPk4DRpqj2hTCuiJcEoqMiDMNEg9P4I1b2sVKjVY+I+LDN
UX7y9qjgWersQEmlq7/mhF1FdqQhvzlINEDoG5048Le8LhYrZGU0iyeA6/sWqWUI
j2bPjrcYEpjviY1T++xaDFk39nHbbEz4CO7DpDXIu31ag7b9+kkC5dB7XGjLRQZh
4XfHqweg0X3KzWBb2AgKupDSAnB/09kIRf+gIwedaIEDPhCc5oXB+slsFp6g7WXd
y3hhfYlnM8KCTeQtYK/4dYDlCuMLCBfAcf2FdBjVjInrJ4MLpy24HX9L0BVSC5p0
46vqHteh0XYgoNpSM2v+W9EX+4w/nnSRqK+ZjagaKjDL4dY3OgngQ5VNIWkasHgJ
bSlH/VHqN17ee4Eb4xw4m/d7eKebIPB1veYpUDaokiDahiVlaXUZigRTX4KxG81t
WgWg+BBbUUyFfboXMPZKaCxcuWI/O7/0bNFxc334oCHGAVjUwloicCldrX17TvuN
arMuGsIi8z1I/Lvmqc7lEMR8FF+Q2k/cdeaAE6WCYP+OqhUK4Oqgf1BEwetrv5xc
jzciReD3HlsJJKIsK5PnBvoCrLaRY8vGkd7MVs1N1yz7sopDRC7a/JBXDQMF2WCi
IfWOIHs4O4tYnLKx2TWg+Yc5vH7wOhB2w+h4fdSuXmyp5YceQQJHHIokbyaymRoU
zPFq5+3dMjFFuaMHUxPCmYeGY3jJCN5vmXhjF4qHqxy6p+xxdNPBxFdcU3dwMJ6G
2BJa1hUXQyxmGUaKk/7lJw+lVeH2IDzlK1Nxc+7vzUIUfURGFa66PybVI639S5O6
ZCEzmn2h4A4DwNdznVaTnsJmOp9O4/wuA/Cge0QaSN7oKgar1sBN2znhO8ddvln3
r9ICPcIcNGeF3YPyJCEl9d2eTxJxw8fFAKuqRJL7umC/hgc573FVvkT3zOBvTGgj
616i8F0EA0DO6xGTPXCYhhYUt86DqzNmR/LxmtClfmHcslq7yMIAkfcurUFAg65S
+rcdTio21YCfo9K1GLhbiuTBQFOkOEdrB/z/WUhCD9Q8+soDXU7Ey9w3dDuSjhRu
c2c/SbeaiVarUxjcwo8l96unF0nNr+yRA222RPvaOSpRKqtQYvbC6EyMxuNhk1tK
S7jP0HYH9nmiPxsblCE6fX4Bu/zxP0NUDDMqUowh6IlECwwkgBTHQH02hdXWxqP+
p9hjzAPWi4IZITjGkVqetkjGxCEWr+xNNUSkjZA6iOlSkDuOYMKfCBUN6GQmkKZo
fEUnHi+bnrLth0UzutGpTH9X1LmBxkSqDwoh6GsLIrIM8Uv1JV+ov7KMyDthL5ir
TYzvobJOT3t1X9JQuF1pVplRLj7wc7Yjtu4FkRsWE1seacbkxyDr1gDVFv22BJVz
fCHsNnPzM820Vy6LfvvgjnVAKEajWSI8ZpF1/0EopTOIB2NDzx8A7acp3tKB/bgd
2A5n2qO94GcyT0R7E3+lTjZYkUad4YXaWRDkOLwps/o4yo6Pne4Gi3Oz2ec3q/9o
M1OyjT8TrAUIYKwQBHOiIegXt44ZmJohsrAk2932JGss02hqLadO5EKGJt8XAYhp
B5jkadRkezwCU0Cg05W5qF0OYJwDGjwFsfyakg1Ct0bD9sRDv/4bCiJJWqnGbESp
f1XEm4Qlde4oYOjREzAOTzFgPG9WCidaoWxUtQcJkrKj/r5aH6O/gW/pAe56yUIM
wEA42MRJgzeOQlDpNwyY02djajJDpaFjtBhKItWuCX+NpByJ3PTIEMYhH+mHGWQS
SELrxMNmBnja75pAKiIFk6MntuBU8uKNwnIXHQz4XFmRxKDv8ZN3RQlv/gNfg5if
lkZfA9TfTXLzwlobVn1Tl2/PM6ovKENK7ppeJMV8DntcihpSmzd6F+/+rIEKk0DS
tvGIwqU+Pki0sCdclEgFzMmrjmLkUEW85Ti+po1FlibkdGKbMzD0ZuZB5m48ZiZb
5l09HxNkJPIZ2aRWjj1e9K1fBI1ZtdBlWpgtdp2qgydSsUp1ScYdLHLSInLdek/1
mBkhZ033HYJn1cPTLW+IP+SoIfHfeN2CyOsgUivDvIei6Um5kGEDTaR5aj8Mweb0
hnKysSLixXf2TVKql51kYp9vzM5b1IgUQ5QczykfWuVzo1Bm5D6MQbB+wHI5VOO6
A9O25n3dK0r5hbRXc+z7wJC6tSnvSl478ZiUhT571beKPN4eb1/Ba0xAnLSF8gPx
8ZpRdu/NPk8btJJGgJWSyFa1USC7Ej+ybyjfeKxRE8jrGugYalcxZJuKYSwj9cPv
MQOLcXF/svBjaEtaoX63/TF0Dxm2397yiyNWUcLCggWVW9bhweYWLH4ecsn0xSNd
EMcIsCvV7NfMq2TYrHnYtgVwjYqtrytm+X9hk4rWF3T8L17XXpHLcLlGvI9bal/B
rI6Qm95vQmMf3EG88vEEDFKyzYQcjkXF2OJHqu+DP+KwtZcSJhDeuBdyNfrlzaNS
oLjD8bDhl1EmxQKfLONN/3d1Zzh9zImE3n8j+b/2rxnMJeGNHmG8ZU0aYToUCk3O
Px8kCECzBvKGKnJyY2DCRxo+S+LZ8AQRrIoiSg16Swy5vRc8Ade56xzHORFXXe32
htWCbJGDdyX2CQAaIgX1xKNVOifWTcLhd6jIdGXM46oiICq3tX/qa5RTIw41rNw+
i6ZSnXw5DGCP0FjwwGlH8cQAe0kGcCGXQMFJ4vWTdyXEPrzlI+sU9toud7q6JrJv
zPKf3L99KpkoQ/FOdaXPkKhmiSkWQ3rms5cC10MuX8lgmizNwMMkxKASX4VBZD0V
YkXJk8114EsKv+EBzymMXBP/gTQiCmeYKl6JF6W571jfBtAHehVLvyhRpZlVFkHg
DJLEGvTgUbIyy3cRYHkJCdTCIVh/ipyZf8G6bopcUnbThIJI2py4PI3QtNaMb/We
nwc/LxcBpLddI86fw9KH41s194G+psyVQsL/nRE6BKJ1w1Z/q8S7gJ7KNdGyUMfd
PfCUDTc4PNb2LnJfc7NWViocJFGQcLfssslSkR10r1BrJTX569vRKW0bndNZiUeS
O90UJ2FfyxW0hm1yITikYeNnfIGBR6ugqg98Cavr8Ezva6stn5PyLg7QEk5e4gNJ
ZfJcA6swpm3fb0aCQ2Q52uz7q5IWIWlnRMw5/vS4pAq+33AYaoak12p/Hosiuk0B
YxKp2QdVRlcApoLzJreSu/PQyqP87vHSR7VTgg6SkC2IbgdMr3Qw5rZPhUrUJGwe
yoFydQpR585HbNRiauFttQBFssp9I7GZ9vF5nPZmFLvu5JpbfQbE7SEoK5uCCEsR
6u5QDb66WV+zy+wJJdzsJvCOzjAWmnRrEHG6OQzuNtmqCPH0/EX3a8Bi4tZDHB2F
8OIjDxL3me3F7xECMpfpkdKjT71OSuoez+0vWfFVYI6zOB39xop8R0m7eM56g7Y7
SfUCPJsOPLizYQPARZhWj1D/IWAFv8/KbvX6v0BpFl/J6eGAUA2F3nZccX/P1zHz
bbWSX6O42wKAdzRGSTWej6iquBlcRBNy5KrBXng66MAFkjZMAPf7pu+/q3ZuQV3c
eEovflBJ6P/C0SvqNVNfeHEyQbUUUEkGcu5Y21DZeTMBPJgnvVHGKtbH0yK39BzO
A7i6WczSclZ3BEW2h/hMfpH+3atyE3hv7VEJvEXC4117zhaJFxgeLfR8yTpXIaC1
O2oiUaPuybzPNR7mG7+cUXo28jwcYLjIHJ/JD6t3HKuIQLZbWclinU7I+YeNT8ed
N8m/+DN9ccLbTGy6Xms8NwSHDIxmEg+BJDXdqwvMREMxtZxQ1Qg/HMMFL8I/3GbH
xNv9g3Y42ltB1IkNCDsCEndADTUzVRi/9xI9pdf9VaDP+9u40ufAo5hEb944SrhA
iFZKyiGU7p3PFkK9nc6vyFDTAVDLxvLJ8a9yIkwjgoAYiwkdfEl4jnOSspOExBeB
RFeQp8BYEF0898CuygajcuDD0H0rW5sGOz6CvW6IHBEnFd7SLgU0HeKWZVDCHCHd
uY2aAIUSsItS03ZO999Ud9UTEWUYb7ESVSyDmcEGTRNTZ3nUrE31tnWO9AdlQv+/
aAdoPuCVCyV++Ye1uDHrDdSYg5EBdzoVA5Fu2PRLyrAAPfICS1nhQjJPNNotERDU
fj0oHgz/cnARTGby8725drhBUojqwkfWiOM6rD+C1HUArUucajk3G0gQ0dfJkfPP
0s46zxNGOjsTl+Lkiafd/kWlkgzSt01s+sy0uBMA0kXhW27JMgH6iDsfgcfbkAs1
TlevTOVbGvlLCTctdXQsaTPFpGNLre3/wuDgckJxCwnMGCDQvlf09RXzWWhkVnRV
eQdxvkkLj4vp85pyfmXerjocrBwJYLtzSQjYgAh+4WyU1j4qJflXlfF1OV7eD9j2
tnfE/r69qSO2L5IUX9OG8LzWgVraxFaDqvqPIFgmDY0XoVuoMsAAVO1v9zU5W7+/
gFMrzT0Xklzj+hWXCAYVRJ8SUBlifVOpIRIfycb8pugmJzLWRJKCB51vZ0LUBRKv
ymzOM+JWgBD11luCJJhiH2yLqFGGTkJg0xIzG4/U+5XXzLlZiZIYd3bFC6rYjpND
Esmw9VN2WRsFGIKYXZjso9zv7RWAqLYu5VZHYcUaeA9uIMVXAPtBuPt2h7Ed813O
dgDuGTRgM0C3yQfpARAZ2T8ErMJi0qZ83waPQxpK6CJ2UQ4rk9hfLD61aHp7gR36
OzXrJOpwKTIsZaE1Tnj2CQx/2C5M/KlK7p32b4drlCyMBFvIETc2KXHLc/2noMFW
lyDnSyxcyJH1sfJdwosC8+KZe87QxHpRIff2G2VhqKeYV+S4uzry/re0SFf3sM6q
JXULp+2lva3cJjTc8exTA9JgP7XwDWreHbf0QvHnmrYQaTTVL7cXWBr7uUUlnzje
q3+TN5T2+zThL2yucLy468/489wLxpURlHXiOwFvxkJb/iqTZF6FKaQHcGWXAG23
n+1yRRw/ebjgBV1A6f0GpO4gY+V6x6poLwZ4t6Xne9VrKD+VtLaNeL/ADc2bCe3e
fEVi0QbGyjt3krTMoptamqYVHSD9vaaJDcbMasTWaOkYoZYZSIe6T433yjM43d64
P1gQy9OoN2xx2mHAgoZHwONys9UCtBBFKLd7QRroEEIYmmCq/nIDJv4/dsJMQcm+
vP/Xf9OebtRUuSIe8ZS9JS7KCOx8l7vEeHwfGZbGbjdsBloX1XmSMAzuhYPce+SS
iMwcAnCl348OS77nrLGGRmPQHF2irhwm75khscew1cT9+lCOCgcB/YDTIrZqK49i
pGuKqsXG7RfckkWZmi+YOIyH2HF0RFcB5cQfs0HUF2V79k1Kgui/cMz99XC9C3Eu
WyLmU7I+Pg0r0wsHwA3WRTk7sBEpU6bL2Rzt6eHjZ8amtbEaAioclGdn4iVa5aD6
5kZxLbzPs/bg2rPxVKmtBrYjjpYueEhlPVB2XiONwqE6nzaganEM4Mkk2FGTKbWn
qyoYyv+OXvAkechShi8f2rCHvKtab0CC+Jsy06MubhFlE5vx++wnqnWnmUukmRKp
ZYdJHSFfbhV2dnucORjK0Sbr3izpyZvWOhfgF1I1JiRDVOAEBOhDLsbGaaFnqpRL
brpCrhXcXe938VpMrD+o5sUbuxBYF1Q58jugEr01scrJltSpoBjI8EP+oay9fLtG
ipwFfAVlDQtCwEw1JOnAPjEHvwtS+fjM+mR4CVJCsBf292txVqvu/3n65gCpH/EK
a7yDNDU4QqwHc+JC86DxLOGj9taNlTcENrOa9UUJcas+LI4A7JlKf7bBa28LwCYr
oo/+zR9/0mJCqVjnfLoxBUrrLJMfPuHRSvILbXL+5ISrHG5f9XJFDe5zXcKZLDal
YmcPfp5sFVk/WNJ7nsqyGNWi6paagXty7xt6dwtZyccCOcnwe1hO1lYGfuy10ZS7
97wT02gTqsn3ivHyr4BYc5xdIlfJeS1uqf99P9iXG8Kx/yO831/FqBdXuYvO9tAD
Y44UP3lRBWkRCSlMCAZ9LHEj+WcfADnqPuc8A411G4/gjshkRWRktHM0dY70g3x/
NwDv4CTpJJLhXv4YeNCmvNpWkJKE8ZCkvLbD2Qkt0tRRuZJ1Q9rdvcAmtt+epYUC
o0BtUZIkm5Ega1VzQhotrUDXT40H/BuMuBv4+jBiV9FnIbKMl2qiuymMtixp4l+J
z+kz8hBJ24soKSkQI1fqQAuK48qSoiR1yxy8LwV2EYEiMg+q3Cx23XbC1uF321nJ
HCWXBF8M97I0vO7gfTfEM0Pr2R5LAcGZQJY8Ev6mkEItT2SdAjkjwtdIgh06J70p
PXKLyO7aMipsLsmZ92+bEsPtBv4E2xhX+e2PiMHBXo7YI3nwurRk/rsczpmsTkdS
qFO2Zllnd7dGjuWcPJQiXTIQ61B5/a16CWrgqCtNvp5ovg60g3oKELsR7nNqoEx2
phknVRor5R+A8VBl4506vA8o7RN8Bw6f4mH5uz65I2ShmJesNIdJl/MBYvcpVaw1
TN6XOlLCge9/gfdrWg/imBFM+cluTDkODGIGLR/AhHEIktsL4S0WZ9umwpEVDVU0
rq/5AH5aafOOhSXm3on6e290kbVoqXEDXcvZIsxCmPfXLJjQbmUen9Zd2oRWnbgB
eQjsnQpmIsjUcnscxLToorvGvJLIoYTiSM+vu6/YwGp8Zxd3GBpdP7I9fmr//tk7
N8N+wPSOyT0iW5zXo+Bfdb+09AVyogO8nGyagI/lmaYBE/xXgW/smYzUchb2Z1Rl
sFFNt8eLwO9djVBRSVp8CdGJmnx5kOU8kkMWroZrbhE1wDHD78NmxnnEWJ31nDLE
os9hf20oq48F+o50d9I4aP6YfqUOIYhAqTckSTuZVKkGhdzH9oJpYl9+QgopJ1NE
hqd3uJCp0vojlaBafjlReVMDHfV9npAodkhqF9XMK35mYsAXZTu1XUxrjuzEWqsT
nstpUQrs/w97CqFywax6oh37/0g2yaZ/3zoMUYIJGMAG2GhCwsmuqAoB2pC4nH3S
hs9iTP7L+/GNgIgLGCrkxqpmb2X8ueOubLUkswmHwytEhNe4YGp78e9CGpcUT4QL
E2Hy+c0En/7T8MtnDnR7hjm8EJFsGgU/mLL2t9CdJVVah4rIhxh9hlYsSFwEAN5F
sgoGpOC9EH+Ym6hbj9bcsKlVy46Uou87vZ4PDD/VKK9xKE8z1V4StSJwJMIL+fxA
Ng9AFsPJYk8A90d1Yq23Awj4eL/Fp92jmKYj1ytAT/hGUFi73cyR/cu+Y2jEzuip
D3ZfPBI6JscHcnVMH5EWTTd/bY2k+eo2AmcHgXd3dRS/LYKz3Ge4w9EjFCLeGUhA
vqXGvxeatS2yRMgn/c7Y7Ix1x0AR7bTtgXcpu+uVJwjS0t4pxK2FVZQNJhx1ZGfe
uMdZS6VXvLzGjm/IV62dx4Pd4+XTQyjT4XvC/L1Z90pbX8ZV2PaN5M3t9omWjA2v
YRu1yOTIXY7c7ukK3lIWKEXDYUj5+Eb+52X5It3QToTvlR3CaIseUO/L6o/7GHFs
L8RQFNYmvipgIzIK+0JSRVSfj5jzIxJoVZGqByq5gynKbHZX2DMYutkfa9Bg5ymu
85ZRfX8x1s85LXaeOkla48CoKmKEDp/plqRk9Xkb9rXcmyjtEKBlt5OybQUK2Z53
GeeVF261qG/9fk7Z29wIS+w+4nuDNqwcoBZqw0mGzdCryb1oXQXPdAiIGuITHe27
RD7DCiEYjy2pbriIQITswe6AXGG7oykBJOycee2/Mli5msP0fXCrXFF+cXPyaHL1
jNI9pX4tp+lxQ5r9JF6JGS3DctYqXMgRhivZdZtVLN0cCEKlBVrKTwm4LJih5+DU
X0V4+hi+1eYvwpOkJ6ZWOMsmE3yJpRX4qxfYg29vOC7HHuVypIQKj8l3hgVmu9Yh
Ksymclv8i1bkB2TlOfPkWs4JVvBs4OPoO0NzKyTL0V0xrFPVAzJUEYJP1aej1LPd
J1R5IG6NSslEQGAXuM9OgcubwJDHzCgmBE3vSO4cxmkOA/xJ7w7a88lbfqjMqXA6
DSHS5C3fBL7WfnkHVZszVfu/mCdbEFLTrqriTuaW9/GACyUEFmwQmIGcOM+wOd2U
4J57u/2i7rvQIX+rWWelT2qWdrWrwF8/6kprxdlUA087wprzUVv1K/P+ZjpVE4Q1
4IZBW2RjaN/IliONMPPOsXqMS/hYhjEEJLLlkvnVRES51JjNzkABNZqruEI/6PPK
ZDmtCHRhGzme++uLThB1EB87GoOR57ewn2KVDCdtn6RyyK5Q+AybEBpWosWO0670
/7ruukndwFDuTKOmR54xUC3Oe/ypOiEaUiKNV/SVnj2KvtizDP1oaZ4pSpIw0ydg
n0BDLy9gOYRHolHfvt4YJgVbZiVngRQDRhwuZ+DT0+Cocc/YckiF/Li+MBaanx06
9aGcoxipwGcZ+wZWMYZTT8Trnsni6HHmthe4JOWGOoyIQRZoE6btJlGLa0yd8EAB
n3ZtQBAJh900xqrzh/DXJ9rzdUK5Iv5E06ZQSe4J3PrB1MRyhQpGu8vUj+vS2Per
/pkuLqGn1e3L5c+BNRn/8bRihL+gRGVBGQlU2SJQXSU+hlJBnyEuzV55aDvGPVEO
LTPkHFYa9BcW133VzUQkxnGar17XweFi35ZVCYHaKR3gfmMzKa2U53nJdZTAgnWi
VzDNCVE2pEGgnhXSip4VtFpmrL/xNiFJh4hiXYexvKr0NlrlXAmtdcA//s2n7FuY
Qmmv5IK7SidqMMQEBsoHyIz7qLWGdC0kmu2WO0gJDpsQ8JQgfxcO3SupN8k32knV
DtOk0l8bDL0ytxBHOx0wEAubKT6oiuj/6c3oUC1IDVsDeaS1O/hz/UFQfrDIA2Xm
RTaFD7Z2TDrl7QH8HieFeeL8JwSLt+coNYtx60+zP5/j3VA9daqBBcbVcYkdOF4P
VyDqZZvhDKWA69/jHZ8nsgHWjKXIy6CzTD9hZtvOf+1Cb+Ho7jz8R3p4c/UEOsgi
c4U1HzwMMttkwpovvEtmbdnVWYAK9oNAN+QUSudvE6Ujyc6jQHVnCaceJIi/eXWY
KQwm3KMQOC7VRJohAvMhPYQlfcB1YbovK6jf41E3LJsSmJTGQQLFj/pcNkntqTVN
Bnd+RM0h5jIThvOIq2qTkrKdYR0WjeE1L/MTlEPCKGIsgg3PDwYwDgVdVt6pr31+
wNaEZgckhcufjf7GVzBwB2eMeufvAEKM8H4BnPEBlHAT74XQ2OoXjo90TjL6cQzP
kd6kqKbgF7SnNsmQ3TNrkTpSeqgI/ztDrnnj3vvdRWZrcFcqenNESxhj2zYAf2p4
mQ+u6UDb907aRa0AS+nZrBo9LX8poT8HgpQNU4SncOiR/9wXVPjTowhNQVuhWfmg
uMr5odLkD64JM5EdtLpPTz+7zPchPWqsJTyHn1AN8hZrp0Gi280BG6GEW3cKnEDj
eZcFe7NU1/iTOfOOU8C/yHNKSWzndMqKwpi91NwiYdgkbvLqio87kQwRj6J0mmGd
ntiK4Pjw75dCn5i7XoOipTaZDIhNcFsNBs64Lu4AyStJZt8ySo3hLrgyC/TuDLf3
OYmXqmy3peyW2u1DIfFsMmax65KE+HkzElEO0qAOnRFU2W2pi6yTepfmShjk5oL3
6Ej+hqstpglK1uQt6NW4VA3p+k1dDgLfV4sKltSv3OT/nX7+pNVdWlEORuL/b9mb
D/veIWw+JIR0TZ3eVGzyoXeRL5MymtHxjlSKQOP29wI4KqGHnn3NJLKMqxFNFobT
r8rjiJDngDMBeP4Qn1JNEb5/SYlsKlTqXYFtEOnY4cyr8tciz7TKWbNIhXPdf2Pe
lgJ9obXgytAVA8h0EvRnuvl64wY5EaMUrPCslSKoC/XGLidsMY+hdD6v9VU+dRoK
PWjZa4OqPJS+CiLHYnGP+yZ127ENbm+Yp/IMMfH17QtNuEcJkf3UrLtatL5145Uj
x/N6Wqdeu2jjHyZ4K0NvgVLJzQzQum+qQr0bgXJH6aN2y2RNu9ulmOlqnvpK1+BZ
mZU+xX5aLlZYp4RCBhylaufrF2RBG2Rs6fLP/OEnay1smfSpuGPldPwPe3wdVC1K
YiZPnDEuBOcSat++QhXl5z33VFAeJAFCtqHNbYYZkqbYJ3vzmi4jymTctX4/dPSN
4x9Kv7T7ufjiD1X87EJ0LNw0Vq2DGvcXsmdVE1lvyBdob1MfO++YsPv1ryf1OmEw
QeTlE/PK/74lMEaRBLZAqgmeEhy+9cWTqgPd0iRCtFCsSxnvG11IoUMd89qyMu0g
zMb+Vc0b2ah1HtSe0nkPIcQuVx3rlgiE81OSAjpfBPSzCORRqavBfd0Tp8qMTryu
FiueFX78itgu2wblqdIZWnag+MWQVD80U/YdGNkvQl00ZjfHeOs7vl1OByKPPQh/
VE8c735SpTlaG+rtLu9eQZzQhse5gWbHAAbwrDUNhRbmk1NzOndG92/x+ci+tJE2
Hf3JfQWcfvGhyJw0/ubgJ6T8E79fl1LIfSJ9eNmAF7yjEpnI5IjgVrFX7/qBh9n1
QKjdC7vVwT5+hADCQWrNQVgAr6u/Bfuhumr65YReVBH6p0yYOdGXZWbjenoRLaj6
HeiFJPQli63CfjlJ+IM0R9zuruyfiaIKwJnJm9eaMaTtHZcSYXfku9Xz+jZQNsSQ
HBBdfyqh7vqmfMjRPz/Vd22ezKHpQUQmZHg6Wy0zwQFJCoRNYeNZrXRT/ct3Dl8N
98H7zy7fFMfrl26OIivsWRVrI/SYBLklzMuH8+NLobRFD42Z4AXZR/WbqrJOuHFg
w7wlhXEHpmX7w3M/PkAQj8FquXU3VF3h8bhcRkpBQXPf+UZ/MJ1gI7d9t5SQdHiy
IIFeLQu7MJ3Droq+F9J40O7D3Q9Pk9wn71mzpfmHLooZFR2NSAUs4NAL7BuGzhF4
oVhk1RW1+/8TkC2F1aFi0RV5YZydf/7hkNmcgX2InsGiww33JgujFPEDA3sBdXZY
hSYZF/tpo449d5Mxj4k8aVz58oblSxQmqXj5Fvod0TBQTRay0Jeid8781YErEpxt
gMKDe4XEdX9wwx0mpJytxHIcbJSM2FQl6t93GAHYSqDPkr/XlQ4E5ugSbKFK76li
Df3tdw1Qc8PRJBFTIYMMka0aUVPn4EOWqu6moULQGqKKDGiyxtjg6dwA0peRJHKo
Q5cD60O/xIZi0nIb2e7SVpjhOx16APP+KPy+jAkvKzXS/Rz5eNujWJTp3MkFCBmT
Mr5sB4iEXNf/KM2QUKqVevz6ctHNZyFZRwR3uubT62D5jw8Cund8xG0AVtZrdA8z
CC6uXVsvZ2gEjfrlmtpVUf42Ons3B8JG1i+OChPyMhQ6iiVehtgK5K5pphZ0U++o
rrlzVZ2ikSSWIIs0aQnq+86ro4kIAxJo8O/xGFBdPmeaMQiQQaB5S9UUcs+iXrDk
tOrhAu3b5D4/AwiYGvxVpk+uIiOvc1ybLZa7EX+Cm8P82iDArSy5cJ+OECXax/js
UeohFbppRiYnfsxk1qlHHhJh6Ceki4x8mBvXqBsJCM074jNI19bD57TO9DV387pm
lIfUbplxfugimR4XdUgGl8EOj/LS0eccc+IeCzKPdkzjc2VChWO8s3ceYXunm6YA
zi5M6TIa7J64bVs27ZaA1R8uCOQbbkXMgDA7G7jY145tI5IELQ9OCLFNz4LXgNm9
CFt7PQdrGqFpLd3A7JhzqV4cOWIghaSNeKyDi7LYd/2ik1G1GhnBxu77NqvX2dWQ
XOpe4fb2e9cZvKmr7JTkfdlmGNWuWcIwsCyaFmVSdnomcGz2VnB2reVfndREDS9o
AcdRVtdzprpszqJfoA0gxn9+8ucqRTzGlUsNNosztjo8HgDHYvm2NeYNSEpt1bvd
EX7fMqR/kqhC6zMek2ReOMeGzq1xsCz8TSEYYXJUDZ2uGqmR54h80x8cKokqtO84
G3Jw/LSGZQHM23PT7xk+MAajecZ5YhLfSO76dEGuPrHlK09yJYdvcarxUeexqcta
q3mIovZiVP0yiZyEjtg1uxBH6+UAZG2DPm1NW8Qz0gJL31RgG7d/sHZ7I2oE1ZX0
GBBTMOnUUrw5fW+EZWe4nLL9qXli9LCyiWVhsB7/c+s4pUmmkPAnoEhE4GOJKsAh
hB6ZxeuPfnBsVGzzoWy3PQ==
`protect END_PROTECTED
