`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94VI2IkrU0ROBlaT/dFpvKnC+OS0wR3aPgPJR9RdNXPmgIJ1FHzo1ioKphQPiwya
8+xDyYcGhGmgVohYuMeLIwBgLUynENxgsUaRSpiz0YYNjwQ8JDG2VwrwroTCa+8N
c4eKnS9W++CCWRXt4y80GYQQFkut26P1meuNTA7B5M3ZswxymtYdWO7F4FOh2ikF
RQwd3aTGXWR4mIQLSWp6MszPAr2vsmp6dL8OtMYI7vgS2HzaIcjObpoiEuTYFpOM
SmHzDt06pTr+q+kS5CvNqg==
`protect END_PROTECTED
