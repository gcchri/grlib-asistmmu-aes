`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OARtFl+G4q/rXWC7Yoo0pLwqPAJ6sTbrLuaxDdIZppo3FnfRQmNs8lOOlyP26HNE
UZxdrX6Q9noRAX9F/XNyPS55xgXvJfrTe7YFhyJKc+NIA16l1jPT3GWBicH/aPPJ
S33YS6XajNuX0pG3dvp/bTySBQFclxEfNI5lsvtPyhu5NbbqeKweBOiL7BzJPEYU
JtBEUl2CztVsW2Gx809f0ETiH+mTl/HxT+8FEbkqdsmvWIjNCdRlVxRKQMRtdKyK
UZt5ZRtV23ptM9qj6iWTbHbPiJm3swFjZMcUkJePIq1Oz0c1fbKbtJeC2SfZYgaa
48OSShXCSd50uOG+KSju4Q==
`protect END_PROTECTED
