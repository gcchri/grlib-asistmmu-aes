`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUH4uV39Fj/v3W+zautiTk0Q/WmLznsPFNuYn+9t46/JwUrq+Xt2XfDrTKWTQDTf
gcvxPLQLNebVos6txf3WQjsteqHT2xK4ruK7j4JJh7f5UN7VxB95fKww7II7FC5O
r9kCrf517fN/RzHGQqVj+ztpT+9+rWynJ8Cxmoeio3bWMuj9F9UZewNXFF8o7W51
jCvMF9jBS3Mw/9II/EWk/A==
`protect END_PROTECTED
