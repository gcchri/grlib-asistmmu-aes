`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MiSEDg7H2VhTngRaKX0QLMYq5dXMI70ELwWCC2MB9C7fn2kFYjzfanTJm/Vko/hA
qr3dW+iXb5GhKxrJfsA0L9Q2k+PGY+epFsUDOz3UEoMc8gqZdJupp2dqbPy/xm35
SnkHsfnbNUAVPD/syeebVPjMalaJkGujNu0XOFHnU8jPs42ypkpRSQ5XDAuz9X6+
jGy7LTrNGJ/MLMtNZ+bBDKLW6vSN/ttgmWFpCeSPBn7qjMcwQj3OKnZ8WgmM46P4
6+CMxhC2pRHpXv5GzAeXBiFcUKQmazza3dBJWO0o1CbKlaxUMiJ85VfLYX4y1ZMq
wmIETcDy/ZRcF5Q08SwSGaaXarmUm/6Amx9TC4/dYHfGofsyQ+oFRVbtAsgKJOdJ
Mwok+LNJuI6Jjar94rlXSWjH144k3PpnHhOFvo+BpQg=
`protect END_PROTECTED
