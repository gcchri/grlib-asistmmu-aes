`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBwC+Uq0vWrjMCGFVBeKlx7qyPmpWOOkSPa78U4X9M6YwCPM+Tf1yNX2O5e3Niwf
6iVjSDVcV/pcPehtMgmAMhhQx88RiLVAyk3LjhemsMO8k2111i+2LcblirVBrJ7n
X0Btap+O2e1cXD1VICSd/rsHd8tp0bpgtcdsVlk9jBFaVAsJqSxUgWZEfT3YxkUe
1DWDFlQY7ubdtmzGZjfuCic84bsF6yZB5GUlQRlGzK6NGOmDTJSg00z6zXO9GuKl
omuA8hKJdWH5SBLTITJ5cVFAp/+Mpu7/dqRbC80mYaQ7gNXOBfD649fm38DI7zml
WuoeH2EgHiDRTOr42rQitZ7KGEKazfkSn/PF44xNVNDyf2i3uSwcNP+HmR9Y6PMV
jYLi7en1D64om58l1sM9kbCTXssMZElsuJtnAD6bJ9nLaIP48UO0p4rfKVTqmncw
j94fyORUDNLlx8DwnWUkFRslPX/qkrsTjg4aeNUrBHH6/ckeV3CANQCP7g0D06zg
rGxH9vcVi9RnUspxuakCOEK7ySGROzVXfbG66vZ/3dm/N0GcpBW1lhR+M6ihm6Jc
cKXVIKExiPrdV0ZjmLBzOTTj3Zq65cf63anwutm02Rc=
`protect END_PROTECTED
