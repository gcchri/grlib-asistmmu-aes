`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
epl7VEKNCxt9m5Gk+Beww6TQ0J3N1VA8vJmDXOEmjlsquWPUbbRMNBeC7e9vscRS
+l+T0rd30Pe9cUdxQHE3mo3GIaqHTWpRNspy1OMZ16aD6vU5c3QmDqKkrbKz+wOs
zQTzWR3dGfTReYwTU0ZqZovUNZMTpxzlfg6RSyJ1lhiqq2j0v+y5AA9I8bU2/JUr
EcC7yA1b66zSW+n+ijG7dBCG4m6t6Y9G6p2n6g01e4IZRa8BktEsOBqSit8pA4eb
+CV/NgK09hnKyHrAzFR6n4Rk7haBK4DsQAJNVeJWAYp4dzmFRZXFJoQlIkGA22pL
9ZImKd9VuXMlYwfSbiSeHuroBP9Kex0/QQC5yNF3kTj7KUcUC4BS73JLnPHt0Y8G
9QpmqAwRKq7tdwfpfKKUnEdI5GG1+8YBKdYqwfZzyLdf4iuaEpQcGCl0HyOVoXAI
BAf3Y/I0LSSgj3hEDxY6G4Fj4/NOhIC1HTY4T45aK6raz+wVts/z1sHkoJCr6tbN
+my0j90p8VwrBzwcFU1vz/u/kjotC9MapLEvvX7KVnNux0WYVFKj8pzx/XJKSjoo
7q4hBb4tScNu4GFbgv2Cv6XRSgqq8DvNxNgwKzxa205n2CpgrrRwcCycaSqHU4Cw
wwGLECcnya4zKJZQTTnuQT61ejCM9ObiqttQeC8k8nIRfZgfmBhDha0uRQzB2bDw
2656a0Q5RyqIsLBa2aPIGXjv3DmR5PlNP+3Rj/RUhHe2iMoBYNIkQoW9RvyknFrX
aSGeOVzCx0xkD9+rKq1ZMPbcrpz/BQj0h8JYWjfMTC4CLsY5jaLI2xpav6t2X1hc
Zn2AKkXKtkW3c5UZgOQcBNS61kD07MfUSMOLumjh+5eNlWEY2Mpn1jQWUYNL/JsR
RvXpzetxQOztj3DyfI032HD2Em+BiL0CrVua6lU9bXORdELuztbH78MVzeKu1lsc
MyyIsrryGcedaBVT7/Vhf9SVyU9R69plTjZtvKBiHSBPJO8tPwv39t7SgEymgpkW
hb6mhFvB3GcY5tv8jGDWnK3t9V5DR3WxK6oAm720nNin7xtcrnmLA2EFKoB5aQ8n
FrCoIJBjBfAJ2kua6CmPGPz8OEw57zvS9y4lmvM7WVe9u694Wjnx1NI+Fa3L+ldU
3l+ZmoXLKmHOS1xS3175OElOCCLkQktpogvgUFT3y+LyBXL6+pmc8BHqtk4ALKeg
Iot2iRULOWwOxrW/yqYdhQ2WcqSoA1F3kmtpME0cMnqizcT4gv1f7qJUPSwuoKLf
tWdkUClR0YH99so7oxTGmK+nNzUXK7VCcLBYsX06uCgF3OQwHLA62j70jBKe29W5
j09RW/25okgVZhzNjRK++dPp8jDG8i2z4exhR2eL+XLJG7KKcfjwlLEx2Wm0A+Ed
gjl0QRZRaex75ZgAE8JROgeQsZc5Ks6CC7eK9FS81etIKT0CubAAUv+Mn96fk62p
RTvpLOKDP6MTOxK3tpEQtS8hHl7Glh8NXn4JUg6pzVas+15PUYPMOj14w77N6R9B
82aDuVkAsss2SrE5Usj+ce38eMwJGNF4cM3klMrYrzaTDE94lH7gLNySJNuNxBqI
ionE0L9Jfi4EX9CiLYlrA1K8MJu/C7JnbbNJTXr6elR1icwSW6w9YAMO3zitOySt
G3IEformBNJiwAq2/5QbdCxZG+ZCcV7PyFWgF/y9bc4HSpuCREwXNSH3V48mJ27O
aVb9gLIbn4lFTVZ+gxuNhNZ8UPnEmRQfGuex7T/begwM3rHTQuhm3J0fn+hbqoHP
UVaVAc6MfbBacXfrNC3cw8wCEiHEPOScZ4BvxwSe7tySipcGUB0oMDTZ9quB6enc
brPbCjiT1Z4mDXoKPH7lqwxXjNjC3FwyAyZQs1VTHMJ2118mYrSaTB6Qfx87k8n9
CoZLPBERma8oOlkNwze9qrDA5XialBgS94zaBnWKBXh2wh0cgOjnvc6n9KC7NVPb
+1dbquvq4wU7H0DgbJDABzqi6p167wrgSzV8O0vurfe6G+mKtojmnc+//U2W4g0N
qY3+Uy/dZhp67CilveJwV+7cLfh+5GLIbadGtS9IG2thpKst8eDd9yvgyoBMPJ7u
FYEckX6r3plXvfG7+Itna7dR3nKX+519aHEZnez4l/RSJg2oudAZyi0CCpjhFutJ
2Ch6gae13cLyeUlKTJhxSlLuLuJSlmRpHaQJ3rq0iqPq45HQB4LJp3No7VE6Xpd7
VS0PquamXf3wNOUR9+vAvGjM1KU3KSO5Zk75o4jfCR4stc1tRusMOYRLcoji6Dbc
8YqW8x5pinddUTnBmqApDFXYQShsHrcOGRDHzsSzRzDWgucnoxgyXVSndsfXjJIn
91L81iOOqeM5w6J9GmUCdiiMcrdI9yBUqvFQvM39cHmDx05QxZgbAE+pGeFwb3KF
mVW74cqIkSAIVZXdlqKiyvPPp4CGY/FiUIgQI5uJlK3C649vmrLanX8vJTBY2M4Q
xhJwxhFi2SC83cQIZ+8mAs0DWPve811NjaOUcGnVFBuCEc+drFeRCn72QBqQLPtz
HCmy2Y7y2yB/l9L0C6ocYcZt+rt4agCqem8OS3RL+l0M9ZPozWdSrcT9byebwY8z
EM66FUe01Pw8lCUs64aZw1DY6KLb+3w2LIObtHK8Z2IDY2u+NtmwiFFR2/YdCj60
5rK3/BHiYVobRmgyvJxDWPch5d823FIGrXi66JNbS68qCZuui0TakDr243BKwb8/
E0Ibmw7OJkWAhllvmCukep8M8GJwh+c3ch8styOghAECmaMgOS+XwAiX9eB/YBXR
f+gFa8rOr0zhX9/E2PVIR2mSuyeIJABSupUezMosM8exxUvruP2k+i71u0eyuJ0C
TbPZPOEd9F1Hfl217RHIyLuAWtzjACLM/yRnKzOYidjGBaA3eYRT7TPezG5NpyVw
/3Y/cBwUP1IhqIwUVeCxQF3Ii52qZRS9mLJDI/KGedonm315heMnghCiXZoe/4t9
GRLBFrPJ/qcgWNqDsxep9t1jwWEMcHad80bqDs3ERnKl9fhJSiHiuNlZdPQWusaG
bmIypPdY6rCpDehJqNm/HaambVguRAN/IL0KT6A3gbzgGV1OGSw4MANuergMTKYm
wkiLdbfZ3hhRnPYcoahcWT7pK5En5EdVxYSytSOjS4gSbXMrCj3RgPsjn3UVj0u4
qIqk8iMnfslvWTaArJwaq4/NgZZlkLhqjNTZRby1XANSyDr4vnPSaSSoJhul8Svn
oDq7gcDG/JZexq5RNcWg085ZvPoDgQMV5XfFKFKuygRL08gQ/fN49CHLO1ycoUIN
t0cqZq3HKHoUGIXRAVII3H7ye8rqGxxaSUzqGl12CxDeNoHUyOblx5jG9/6lIDud
NSqItPBLIguju1k+NDWi4/L0eBRw+eFXMiW9c9oRSuadqbuy6+3ZajiL77Gho+aX
Ht5qguEZRUyRlDXxl38iHyQPNYWAgE4w/i9FMkFomFlT98edQd06skT51oSv/xTU
rhi7LQWRpj2t1Zjw87fvvH4ExS7yCabNXXhAM9fKccJlmrMmoEG7IUHHQ+z1ZHHK
0n0epHJYmp4gGWPIbwagZbC05unjQWnmkooi3HokIXVN7EzfqNrh+OtJY1a1Ce67
eyv0NCPg7b3pjJQmfdKvilR6PKvexBXA8qXOLSEtWnXcw+eIyMBWbTbUBJQ4kzrv
7phjumoaxdq6UPNfa5zdrVthbuzyc4RG4ryGqsB8T/quuwZsYBeOed61u/HpgrDG
Ts6xayJFNdZQ566S4fogxKwWuw+/QbG32n0ojHsfahEvjiB9bZrSC2J0V1n7FOyy
8PmUmIrrtpyJKay7xGQhtZIH1f14ACPsHIndOv8gsmhIrJpsfL1odCkpyy9g4MzG
9d8EWcbuAyCNZGtuB+B90iAknaw5O60DT/MKc7eswLYGA8/RBvTtyx0OlqpI7qtx
ErmcAoyuc2S2s3kPoknM9H43/olbP++5B4grESu0P8VGiMFcuf6TWpHvrmaBH0Kx
4h9mNk37wAjxRhNFkYMcIg5f2T8wn+Ky9WOvds14HUyCcPIfV1u55vajEJWxTkhU
mRRASRA1Bo1/gTYtLZ9txb3hcO771TcSrgeBhHpQmu+lEkgJ4DlNZuhNF7UUD+pj
CWWgtAejNQSzERmB7GkuJ121D+ixplHMfq81p0O1AhKCGl+vnjRxVC2kgUAA/J33
ooX8D/Dai9FToMXZUxVO2nobX4091L43TYdupcquYor3Gn6DJ/gmCWnz49vfzhPs
6Vhf7LGIpI4AHfoOLSEFov9BsvmC1ChSU0MNaU77HVZ4o6skSE927wNij5zKJvfp
05ob5BFSkNCBdRTFZz+eC7dNKIHlyJYEFR3AbvhWLZwUaCpNJYkXiF89YbsS0LQJ
poeAhszwV0y6RpwAjaoJVcfuOmJn09oTRSnkaDlY63+JhmeoSwUw0dlJ2SlN860M
H1sEQHsL5klGB/URGAXkLC62RJIHyqTrSMAtM5x+o7ErAhfI6zXf5uNEAOncLpz7
XNiTheC+iHTXZ+3QEN8L7SrYD9XIU3kzHWjAcIC0+kAxFvyf/AmHe8opTuPAgtTa
zL8JfSZ/31m+o2Amc2+momRVo5yMeWCXKGAoy7CoUxEFyhNPjY6Bise1ccgENAqm
ZqVq6m3an+E7D7+QUSZjrMNzfPj6pi/qdkw67mJvHjd4z8TNg3pakw+dRjqNS0L/
HFins/aZekGLddPPFO6lKhPcevi+Be1jom/mq/Fk3NQGxrt8JFD3eHqLnCHQNh1x
QH2Smjpq4I+BGi5wNYAdDGurMOnhXwGWgLjBpdhEYd8u6bIY47nDz9iVsNzfYBRR
GW7mQ2RgluQhzvTcLSYmxmVElmKw8B7BTnCqUAU+ky2xJglCCot20jCTewyz0Ue3
M/Thv80XYoJm56qHVzZ/q3C3UUFPOc7H+2cnZYOlVnXxfVmaMya3GD2zSN8RhT93
w4uQt0R6ZdJBS1AwZgg8/bLI/BlQeP7aZVZosZ/5DWZ2rYfedday2ZZpkxRc/QLZ
mYL/ISgaluzrCs4eicu6zNaVAdruQNwuVeP/8SfyHOJBAmZuAnmh03LniCH/rhWl
irhSsPbsnfQ9M2hxrTz4/iYEHKbJ6Vi7V08fbIY4bRtIgmWhB4QYdkNWYI2iYCOK
qCYXml/piZr68p+TxF+mepXuwammJarHUV4LRPxvQoanqmWnPo9VC2ELSF1Up8L3
MeWqmWgHJllPtLc5asRI4qdEqnIETGCQMiLL6ODHQDyHIDRQprCUxi4rTmTG/1ks
XPcBGRXGgfmT9a3cEs0RRT09nEXJj/L2Sg4+AeUTQE4UxTFObicKqq7w4bM6aYUq
Cb8IB4fNruYgo5YcC9Jd19OFLFyjZNSZsNIoHO+667fc7AVpaN9a/R7zipdsbGLK
0mSeVoWNH+BnFa6wbeiBUI0sgjxdq9pLYmycgrFMh+mNlRgL9T6gRnnugaVaX4Eu
dD7u+7ZB5alyuOI/0cKjyTUG2N/gDzkrVlxeXIpO1BVVAHhgfYZZjta9VVTAHN+M
Tfmw50n9ha2mR4PvhFHfi+oE44IWUnQ+Pgw9TYGHnBmEBZdRtwNmNUI3hHCxZv3d
sWNfELlDw2cCvO9PGWzaZls2RXWf8P1tGhuizKqkCMaI6U27qflKuvbwhUVtW5dl
VdxLku+czF5+tR67PtaMGNKZpb4XeJNY6+LyQPHC2TzYkHczVh6/0K//UJLHYASB
XwaRRFMIiWFdrYQNDMh+O3qouQB+lRGXYIYIUEwxNIOLnDaEybuudfJzU3MwS50t
pHfQuN+yfOxtvoLf++CLuUpzuJkKS5w5Y+PBZP0rOvnUTaCN4Zera659mdqX2ocN
iUBH4gkudKdvzHyVD0eTOyTt1ceJLjP5q8vEFAkQELmtOTkyfdOxAIyQDoojKUj1
bpNMw8IQDt3zijUoXfXbh6dgRfNEzCvyeoAIqteahuQcAp2jua4BERB71BKYrfn4
wE4sTLegKzGRvMPirM1a7o75Rt5OwD+b+6RoA4gsbTr54prPV6XCbtisSL3bqIaR
0VWu7ljCSxiMe/lXPx/EqlGoroqaZLOSQB1/ul0WeavU7v9nC73mlOwQZ5CNo7BP
GZsSMedGl+hNcwS/FnKXMhMBCv9ss7+SIwOVIQDjrTgUcQz3RRdTXimDf6a3Ypht
k1Tnd+gm8XhQyQ85GuIddnvI36rRRa1+rLx/IVYp+TUqTJmbVnM83L4HFT1pnge/
x+DD1KvDRBe5JSAYqUOo8HI+Yz1EIy4lnixFVJI4sJbkuMtwdMe/swaMYSpmKVVF
KGDJp4WnTZHj/hA55X/5+c5N+cQb6MvNk5Dh12u8UszkxRxTmR/0IevSGB842s8o
bWkyAE0Iz9LYJFRYOhK+lMn/wpsj54aTafKB3LiyL8GjLq6NN2BDIBLFoknQmNZP
HvkKhQ26zCncp5037juDQHqjTAzc1uUMvP4kZQ/1WpYRz28FiIRiSmfaU4fIFOOr
7g+XA0fDZJuyV+RynkBu+CO2tf1NZfRQttN53nZdFOojKLOUfHiT9xbwyzVZ+Kfj
cnPvS4a1HyTPf1LxCGbICrrPFukc6oKytSaOUtR4oi78o8iIgvieN0hmynxgAq/E
8Et5ybd2ho0+H+5YYSIkUKrcjpgzGMcNNZtXn6VZ17BIHksYcD58/bJdrd8ipwPv
0+KeqQhh1mOvVSEpk7lrWxVPaHlWjM6nGSzkpaTo1kdmIMR3h8Xtp2I3Z7dxa3Eg
i8sTc4eO7i432bxzV1LPJgEwYoNshmg2PdtjM+FofSwxqN7imn3tc1Vf1VgtPJmJ
e66f40MVuGsoSrLT327DYkdK31nzQzYWEaDe+ycM9D161UtcuxNoXQbNNoyAt/+1
1KQzkvXXhU8f02SDHQ/1Brma8RUFpEVsgQANyaFiBZICgDA2Ph0uFM2b41L9uXhD
LVGbHhIOCGIgAjgGQFKdE+pFFOtLnaLy1PaDPFR3LGTuOPnERaZHNu4pxlPxsFFo
m2PZUNr9O0lEh8/fxdCYhBwM26TjHoEHPBuhtpj2caaAq4firf43Lu8rH+lP4UX7
AJf7x5EacZgGlFdLtHIiP0sLIrC9A1tGcSRy+de629y0w7jyaQ+awFrIkalXNoMA
iBrfyYalDqdkL099clM7hn36OUof1jIBX7MENHvDzwV0HdQL2kf/+IslKHkaTWFk
Vr4sGvSPB/VXjTLmEGA5v8cSBP4FM/KHwl3hk6dWUFWvkpyg+PhB5XZSqpgePP0r
qAhgi98rv31W3hHmycFPBTi9qKc5fAItZtw2vhbEnJmzOOlOx9qyGzcn6UNJGMkY
9vIlL1SoQGt2So+w8s0l5hL/eoj3dfEZ6ZiAO4D2wYJJ20F5RSVvlXZKCsNu89Sw
oTguNgWdJ4rP1C/ZH9pmOTFZc+lzjLR5IMunXp3T7rgGjhXecXqKqh11bJWaXGB9
9b283Bgxbgfh2PxSjTfaPBBkVVasrJ6XGjBps+WXxWnBpt4bwTQu/Ub/PvMLGAEC
yNawjqdUTqlfeJj+98ZV/2P+YRXTRZeAfy2gsptfa0gbhOM20fCFkXdH46L5C+Ar
K0Cdum3o1W4+DCCFAGpf4+5UznkMftS2T7UwJz2aifs+ZwCcWLBBht3CrlaXsxHh
bChqGotKDZMcZm5UMBRmgdycpbiMWnln8UgRSoLFTe2sOXZ3aYmz8ah1Q20xxydC
DjeUjtKT7nsv+5KopPtpY1y11t2rd/O24/c162QrkchDt/g6v3K0JISY+fwmw/Bq
w5eKRliqVKiMTwFOhxz7dGU1ufK6g5ma9Hk9OaLID/vWuaPIubRGbH57zjG46hIr
56VHA3+GD3FhIm60hjYuJ4pPt0mZ4oIIcUKiARbgnPk5c5XRB9urHihicDkQVhy/
kd1lmS/nvAfJL+Wsgr0x+89G1Pm+iaGJIKregAMVCkKrRfRUuRZ6VVrrpaPD4TeR
qmn9U6eT0wWWAamOaMzfoCV8gdITEAUg2THAXqUSKzxOXHSCoIQvSByoKZcJWG3Y
NfnA6w5JVV/9cBWMUTTGOIzzhGpW22KNZVtDtqFgLJcLut2j5PEXQjhjwFLzVopt
EHWJbHWMDEx6OsMFlxXyGtiYgAS9TlboyYjd0w6wFyE90eSraA2KcwOCQVJbEWq2
gUloP7C8gbPbl5n/dmLcwk2XqCqWZJ5caT5gsbtqeU4lmmTBQrQ5cQa+VGmEbvc7
CA0DylKS+2FpQCo/y9YmBV0WnNnsiazFNEZW19Z0bZbE+QdW5SryCES0/lCTz054
5SGYcts+8CstEVZYzfv39qLkMt38IZ+ZR6p06E+zKNBCfA8wS7uUC+R6IczWzMQb
CJ/j9ZJBPwtoBJyuAtqG67u/NQujVaEmBqbb+m5PJH3P4y7xUFWTkHkacDFrCTYl
cnbcT54T9MsQPEuuPXb16/C7bS5eYZxmVKtKQPu9bszSvJzewcnS4v9PYVfEEDrf
Zd5HHZcJ3YXbnRZQpeIgBsKDRHsM9Rf3ff+TQ4TCLjfSjJGyVSpRxpk7ThD4e5+f
sUWuFwUpursNA5mGxJiTyWsM5Y+TpTP7KmcjYqhk04EbN0dqOiKtj4Z0RJjM3koo
c2V9iumJLCK45G204pYVRr0ejc07CjH313cdLGNvOWtPipNGdMPhJi1qx6x55mwO
XqK6YczYZhAqSIi/SfAEYtp7X3IdjaFpnFr+0CjUOxz6LDzD4j5Vgn+UwD48ZWVW
q9xlAW9gk4FeEOiYSPHvtnjT2LWkCLxNvMp8eVCLV1EoBODiJTu4i/kEzcvPzUan
+sS7CRij1S2+YVHi2G59/uQpWHujBeaeag9PDk4q6ai42eQH7Wvc8srZt4Miioku
XdS7u3xPb+KRQNMAgJzem0B3nLj2VXqFnMSwwCif3SEdwR4zuhNuO3w73krsOofz
7gdF6J/KhGaIBEpoIGSv1Aw5d2t2P1FHRYfAR1GpGEt9xzV+DGxtVzcYOomMHQpa
U9OqQ8T+EyVZUVrtJZ3davVQDR0G0O4pYzK0EoITcF4c5bm+TPT5++Cr7EIZyUKy
TU/OjXPqF30dYUnLHTBBeMv+eEOhd4O0X4dWJjnMDhUbCAQC+zZp/QL8PiDH24CL
iKcxUhLyAzRWIVLnQnQ3+bF0Ht0ECWo4I5KwVogINrzswSM2a1hpNU5ZcMPSCgvk
TYnkDp1j6U8h0+GTcPlT/6TvqTT+C9kWhOF7DkrGtDzBD1SEGAktInatitI83Pzx
oQGwrGO5T1kVgLmda1YPB6kQNl3xTIyCRt1r7DA/QPmnPThV8b81OSRWjg4O5zVX
d0WfhOAfTj41DZYJ4A2xOZPm1SrhbDuJsdq0JM/gfB2YkOabXC8PQ1/DLikABVPN
/28NFv8PKkQqe6fz7ngYLH8rd1XD93+Ic7Rnx8bs8ULWnC5RnEaYv54kxC/mYTGC
VLJjNy1psrACckHtMGDbIlfjlmB6GGHLnJO1yo4bQrZDPnblftiPP1zKtbTPBjs/
LKlh6lWi6hJD7xDsdLFtLmHFy0HNcmapKoml12g428QqPFmu0UrC0+upvWMtOfl8
eN08yShQj/q+WSeXApdAXG9FGPZHSCrPpWGRn0dPzszKx+09FQBlzi4xBRcJyEbo
ptw0/zD5AcF/nv5j/cICNbG2h0P9dF89xkPJFzuby/cDxoLWfA5YgPeAgqHirumq
fW9vOQbNq52Gm3SmbBetBc/8n9VBZ+5xPkIqaI2ErMOXIMwfsHkNsPx2amNdLQE3
joAEXkoZbHeiajtIcPFpzK0j26eESXdsdhaS1Rkh5RUI78qon5o2R22HuI9miq7B
6WJClDo/b3JNdHjdqrCAKP6ZbbC419G99HTwhoaahrSaqHtkkScg7gCY20NKxA0m
1tmw3mfhy8SrP/rtrMggZoG0jRgJod06F1PffJKECCE7oJz2/oJApyxcFQmTyxoZ
nhvZx94MAjDYAHm7Cs/Mmwfw/eIpj8JEJb49K/J21gztjCZGN63I8qh41U4qsYyx
OvF7yYkyvaGqVLJqU/uPPMaHf/LCwDV8llB+MeTKZQvxCeZDRTyx0rLzjTrQRfu9
EtY8w5sFjhzKiAYlJgbMCFQulgfxxGVsEuWw3kQ+a7xPTWbV/PYVOYdJUqlhIDBN
WPwqpz/thihmcE6ilj2qsEsbqmqq6MYvcfAskwuK2Cjg0bVUbRWkQA27rM+4cXl2
gIX/BGue3AdcOj/8Zk6fDIMschdFHioif9b7BMVpCykfJOn9HuGE3IlBhh2teDoH
mzmKfkuynqusu4uPF4oDKsQEjEVhPEmVIDlYCVnnmqMAJqlOcYr+ec/lYQWqs2ZW
4oqJqigvLb/NuLWsPHVBk0a55RYG6MteazF83yK2cpHGqyinGw9NAP/I+PHbp13t
H64RrskQMyyc1Cnx9YDSeNqL2/xIMA7gToWnztaKLj6t7ktsTvOakISevf4z2+V+
g4+G1+/zzbiYlWzINg/0KSTfPu/MSQgtQTuVEeAdkXaXWnhGCcGQRDgGarijFnUd
npuX9+m+3Oj/m3Dr4nAQ3uStnjxvdIXojH22dGzLkUkVdPhxyaSs3Ff5Rb/PdARM
5VGbUzp+sRgNpGq6KtT3fNtOfWps7cAJHE6zRlNINu385mlREB791WAc63MmL3fY
ftU4XQ8l9PVfRruQcKB1a8HMKL+Y8rco1/V6iilEacTjmLQInFoVN0LewKcM6TQ+
I9TyIr38edomYJa17UPzea7RplBAYm4dk83QZx8F6I+p2zwr7HsPn7IO9qiXD6DV
EcCO7uZhICMKffasLF9b84yG04QzeC7J3woEY7nkXpoe4GiXiz83ujeJW4Cz45Si
W4qdh0x/3Ngj+hSAGISrOoRasA9lTMcWyKC3aGo9vYo0kfFatsZQkFnyfCBQJ6bC
f2a8e0iEi0fle0fpNfOPY8HKuKRX6f8rDTQW/CvGCwpEXiEX+VI5w2ePnLuO53Ir
cIyh4h9XEUIi53QocZG//xKEa3XvY6HRCJr/g4oBKbaASaVWB0qjPzIxWTpYCJRB
ZIdFxHUcOadIwm3T9H3H64qAKRCA2dqZ7koeJkb93QQGYXhhyqU3BuLMTmOpazXd
9xeUKcFqDRljXuAEbVOflIzZkLpC7saj3av1LS7IPffiL+ngCJAp4SFwGDDoaNcu
X4D7iN3TjfL204y2SENTnapLBz6Od5Vk9bWxKIjlv/3Z1GoqqFoDsXD0g0GkARFH
CjHAc4ThjNBY0yxbTvSIOQ+6olApEyn6i52vIfiKNA+ZNfczOY2Kqe7RGpwxDgqz
v5dFMJABmyHjfSV5o2S8nmjJ55U0gMW5Z+NDJK7Gnudc7wnvR372yRxZpYXKwD/5
bTxJxmj4joKmrR2lJMwFRLnbHw9jAMdOgqEi0H5i/EwiLTu/Xq5pJXyR4j7aO5yZ
70Wwx9XjzFb0b0FfsFcHiB+ad+WcOQW8qPClWLrW6AJhx49NBWXM/RnX6nOuyd3U
PRSvJmLsa+Kb442MZVULfAOUvL+jBWcp/e+dxsEeCh0YkHE+IGW54Lp+2s55iPM8
BongpenExlSqL2N37r3EwNH6U0H63vzcpovQOZhMgIlECw4XZUlv012BKyUutdnb
OkIpdut/1dhrzKljMoOp0qhoVGHlBE4z3igYutsl07nh2BENa+lcx60ffOffii3R
KSd8OUgQjFCw4I+i1Rp3kO/zESf9yqiwUMNBOyQ6hPTSu3TFH94myZMWHygWkQP+
Lq7QqwDDieOFskgr3fCHkCSFBYL1MHf67zyfswKDeiDiIqW3x7vuebaTExjUcWjo
/NG+tZsph38lAIXCt1jL/CJZOVGhGke9onaDjKqWDLFuDbZFzm3mbB36KYJQt1IW
RpBCzL1R6lS1uMX1ylk3rMlo55BkdDQHpiEoWBTdnoeU9iFM+SphmAF6iJiZtUy1
kk6R23LX4w3KkyN2zzHhVMUhAxxOV0KnWXuaZdw2sVSSEmkN1oeAHRRIUPLJPWz2
Yhhcb+CcwMsi0jdJYUSotsVfPg74+KDJnkYv57sB55oRZxpjfUAiuygIOxgc6+PQ
cFjLx9OVR4IYM8ESpuSjwz+V36lQHq7ymXZKyB2bWvZZ1aKhRgn9isUL+gxIWPPI
xhTTmgWLbQ8A3zoclfVZgECSQOhVIAV7QvdN647hbtO7SIWR3GVQ2tTdwcmaQJL0
rhqDX+yehS7NByQfE58GgsbrMhXH8KWDxHYdaVM3rCVLNO2/Br7LD8EZNo7hWl+H
p9nZOuqP4RfHCYtJzUWLDInz4tUFQEGpSxKyV9EXugChS373pq8R3tyqDapWwczM
MpXtwp89+TDiVObsje6Ok8jcS6kLzsjA00XI4JadxHGPL303p5VUx/m/abw3RbeJ
lrp5XYY1+ufRk6PAV10/ugmTXePEFFFLK7GXppMH4kAEJKjlR0ZPjItkVNcBg5P0
AYCxGZgk/LVrXlajhY0JKccZe6laETNlFpgbiN/5+uRw0sSIRvAgUr94Gwdr7Xb+
lyeA0AEOXkiTTnx2LuVAJQqKxM2ymc+oAMrByAlqytdtqaSrBl7DYHWxrrq9l6fj
0V8TqJWtwEGfIqGlqgT142QH/irB8l9R98K5Jf+XScZzPhMawYjQFGQONM5ncQLL
VUdqhYfPc905piDZKldi8GSandLlUnra2DKMayu6uipeBBSwdqmBv8zCqxlkKgiX
cYh9p498Iyf1IzzaT+XIsa41qlyFdViovg9pM6WLXqgNEu5g0QWZOk8TwZ5wFG+S
wtZaYzTlrGxsAbvBFbvdv61VUzhTjNZ6puyAuh9g9F2ppD7EOEB4dp3XSRaJmyhW
cAZeizcEr1pnr6sqIRsQ204jraHMzKcdM0sFBtZD6rNKYOxC+1WV8xzW7dYMgKuc
oJfu1v+Pr6RLV75EwlwK2yYStGyZRWuOZFPbzY27sc+gz/FQjerljnSVgf5b2iYL
iWfk92mTDiWPAKh0UVAHZJEcgTqo6Xy23uL6KVeeJhthyPwBAnkOTkVOvD497NpK
iPPTgdIC6LMKnRb0BQ8/XX4JTFxMVAb/ZKCA/t404zRY3jmabV7v+nAqLnUnbMni
RzANijoVlbAzS9sZLydjjJQhVzVy4pQ8oXe/pjRZFr130lDA4st1CcnBBxPeXGQE
28jhZ3PYgDL2Nhhy1WzuUin4TM3IKe+10AcJT2f7KA+wux8s1pTZACPgR4/e0Xbi
jcSeEnjYAsiuNypTttJSC8RvLGWRR05NZprW2K/6vwEd/rngfv3tFspDyqw3IBgi
bbcRw3OVqNX9QPzOLn11FR0Sei2xHe9b7zmfYDszuLydh9ZCT0QGSr5k2hN/JcTe
h9RGsCw4YWDjyh/rVM3B+6PFsK7QYRkJkGZtqrVa5nALe2KaKjJCTSNfwZ/z+GCc
i9PMzOoYW2+/JMHSYoKFnr37AIdGtFmQWJmgiUG4/vlPGgiI5OUYAI6VzE1FeVeh
c1lMkFn5kj9JdL4tfuet9CIxQCogJnhX/QshA9mCm3MQUK34ciyy8WcaxmISGCmg
y0d8XYsuP49ne32znOmuwnu9+flBd8EbXIpfdMwlke/uleajJZUwmuAzRzCcAK7W
fWlAepGcdlu6LNMmcducbwMdXAOhEi2iCSzindwMcKeDbdCvNYr1P1UVYEaT1fZk
ePwBdISbPYg0ribDMUHiALmukZDnxlVrkuSl/BqamJo1zfuotU11mcz4PTThV51m
5jNotiZiLOUmOoidTwhOEjQR/n0XilUKHV07VECo/vdaNV9FWoXlIOLokZAgKSur
A+oxA6O/EnTSgRuDlXjnKgGoGywyGzFkUbs6EbB6xhZgF7VIBXdBvOqBIVaztGXP
OA+yL4VGFalrREksDacYIOSxj93eqLVlIYpgB94I7w+59hDJ1DSJ2sGWraXUdS7D
Ykj+qnkNVplcF1GQJdCLMKfMVhRy/EtOzwWmyYro68xVR9p+kXLc456f7j4eFbzA
wi99PHIrSzyhQZzbTCsZp0et4s5iCLzCp9iudjZTxpYy7jGDXqZW94xy+zyRy42p
7h5jSAiQqi0btCgnLHQDAJkySsL3DCGfDIaS5LEZdDY5Sgbm6CeEVDDXu2vi5Bld
98rifc2gYetFGZEyLj2XUIImlHNS3myffGlCYiTM/dPo+v/KylXwbKRVz3dRPxD3
fT2Q5ByyND4EdRvnoBPTgVljwTy/1Z+O+PHgTpUztu5ibthXeizOGg/EZn24Ymyh
a1jRUm9WcSCVpCLv5BYyVqWucbhzq3O40wjomuCr2JwKeeR3J6Kv5/GHlTNgG/eb
fJu/XbUZvFGmnOR51XuVoKhb+OW9O0MdQH+tnhPS6SOLtaS+pfdfqPg0bT5Q97lI
x4sFTO8iNRlL+hfmDgDU18FYFVfO46OSQLKKArkZ2o7vYdFQCcL1FOWMMQBX3Oj7
Vj7jZuTfQXM31wslLUKSb/1wAd1paL/LrDuHGYIroKqx8Ix/YgPzOdyO6lquRckA
fFUTXuc+XYWhGWVu71U9mqT35ijxAs/35cQ4YqQVcXs9hWmaS0XYDuoNOipsEAeE
8EW5N2dSIlH2FuEzeTl+d8/UAbflmS2kJsljXR/RMYeYVxGA98oMrOI2Q/3dTFSz
Jv4cRr/2TjekzF/zYrSzgTonO//FIf00QE4ZMe5tPtHi0hwBfAZI8h8g+060FEl8
7J5FUqAeL7UORL5pVxmXt8G8Am7o8eswz2j7HFkYZ1suJYLRAhqetKj7yV3zAhsz
WkSO6GNjIq5nRmC3cW0ZpKrEs1qaYZZ7TLg2Q9oJ/DL4puR0qGzkoAow3jUJNhfr
cQXdyDu9EvQ0ZvMjCc988O+t2xlLY7rBfdqw3Hr6hNACv1CSHtcTpuHpy/5q/va9
PFfbXqhUIAJjOhJZugv2i3QzZhu964yexU95edivw2VZa2iydLMa5rVpmXg5+MzF
uVcSDAHou5IoKKdqM/AA7ovZTI6/jSyAJhyuahhlfOcx7Hf52MhMyOPqNLQJtT2W
UKNjxGlnJiJiV+zG3VGEv6JjTaMpqSa7SeExM3mL041d9gsxbJJglsUDGQkEYWAX
z1knpRQzVdZDgmWw3+ELW+gpl/E2TQS/DQlDXrn/eNF+CTEznsn0HzaMuGxKoh4Z
n0kGkUrzXE+X344KwQxObOpfQ1FuYXZ8/YynTCS9M74t0mEiMfD3/NdEudLVoSi5
U+EbiA0IPWDxZWb8dyl7DSQrCt67xwNow/aQknm3gYqNzKGXBkEtgTOwC7CIWjzO
HM68JICErPOlRqLzXaunRbWak8rt+uPwOiLUEsIkom/TJ7/0xv6kwAupIes+whfz
4MThfj7f6rNTOa0lSZaYFyAAFyZnKMoHOaOzOpur6kPAGNYS+MIWrj1A2cpd87Ue
+2viVppKIeS7BMxD6u5/+ho/QRx24jQ3od1USAouvPOz2pSrgsdviWP8yv/00Nfy
g2nj83b+ho7LKCJUT1JfQlLij8Ft++4LnfI6Yf2x4hi1XKjTLSoV0VK7OqMHJfra
ikCNQ0W59qyZS/Zgvyz+veUTCJYgSBpsGUs2p4oPSpPPAtVNQuQMX35t3xSzCrc8
Eiv4siVpdiOX1MKX9wQ6DN/zXHBwyo2VQyUSWw+vGtynB8S7DPBUFv4eJGzhYlLw
telxavICr1Hccvcywi9ztLPFbh33A8bOc0jWZvOpM0CckWBuKccmRu1cpjflhoS4
072VWMsJUW4Akuo/7AiQdWhdV316RLNFUwK0ev/Zi/9LDq6h7Ll6ZE3i1s23iOuv
klyFwP5rL8pGZlOEF5nRY1/Fn+lUTNymwdcpCHuoeJfocakEa3r830ZrohFEO/Fk
r1Xbmrx53o6Ue7yXIhqUQ3haFugSPA266S0E0JthIKwlIZFBjDjsHoJEG3sjBwdp
Y01P90/oPnKqCYWujA1oikB6RIF97RcysIOL3aCz3KN4/6G/PdB/RsCS7B8EgZYv
WwX+Yc1LXEs0K/qDomR9DJaQdGFgNsjeGA4MyTIJaUl8F8LvYt1mDZylUSdmC8rn
1MPpD4rJlcatsMcmRw3RpO6YmM7jTW/idzF/cOfJiCT71h0iJt+LMd5NliAHfOQd
FNNBWhNAMgTG8jYNl+KXyfFHwbSAnvlfw2lQjcNQE7BeliKmaonVIyedR53IW175
nTsR8b9PpkJ6/E6r2Gz0nV2Xtp2FxFJOyAd9WUj2HEV131JvNeRkZW1A6dLQJv2R
/L5j2+DYNE3XtrNgUecJvNdKTY8uPNzbiLOAJohofiupf45wz3WCQ6jPXgNGuKV2
x2QddzNRKEuMH2gzveyWZ8TzWVBEcaJVe8myt+Pua4IfCL4a/Os/H6fzuLRdM+7Y
oJzS33vpiVni7umUyzQ/CKYHDoGTPFccrQCLkpmx5Co3IIo6AlSnTj3tPT4pam4Z
Av/BI/6QUy75X1bLrPk5MM3866PaudJmqdTM0r4naVIN4mXeSkR2YmZZ9UfbqWsI
SiHl5ruMfsg87/GpT1ICj/EYVOS0Wh6GROx9D0WA6I2NDbHJ7hBXx2K6qylfXtad
NF0pNQFhsyhe5sRfumyVe3XCJ3PLi/ixoIyGEpL88jKdP7efAC/JbywWZBNIzDqG
EQ/lha7Lm63Td1kpe1RLov/VlNuuRazzZKAsDbN3vczQL3XOMcFjG9j5Op6m00wb
IX8R99hu8Ap410ogteMp2MSvQqFLRyd1+s01ZXeEtsuFTWOqFM0IMoLo099qT/Gr
iVVnj0psc8Dr3t2LaNhZ4+o6dLGckZdhLSMiqe7QX1ut1df0wmKWJFBM7LZkQi9e
JGIG3OHu3bNxL1dPRwx+xf4KF5r0nncMKF72RuxHXNp1Eeus0WDNxpOE9xXEv+gF
9Mg6+wWmvfypZBrVig9+Df4a9LKvhsBPRZU76WC5UThRmDjIGglZVwkKpttMN6yT
E5KfcCmKwIIyizre4+fIboNtW86VWLS99OE7iEWtjahFiAyXsiHsEPIWVCSd98rG
t0Tt3AdCKgZCPlJfErTeTwxAMroi/BmCfysf6cz15pHXp2l5Vc49PlJafv4SCkLF
bUptEVL/1X/7IwXhMEbmqVczboXqqqVnbAJn2T3kI0hV09hV97VH7wmhZGqcBo2d
9NaGD0tmcxDpEXAwY3x2Kydi7s+7MisR6Xa81WLVMgunEV9Uk6CMMlt9YzmzWxrv
uHYqpsM0ZYbfHaqNuNEGh+njaTm5k9P5v2qDGrL6Sd2zS7qC6UJoXJaxGOn+0c8/
CjgKvoHI0YKGMEGoPyfgOqbaC55D57V0CjujIf3/JcJZpq6DFpVfgOOn4oA02bkT
4l2M6/UhO3abQBJRbGQe09zDAmBSb/X7XQKt0IW8gqWcXLOcdtRRme2TQYEx+y24
H1b4zLWJorFdoRoZ+RBpSCYnlL6ljw4ORr51SAVzaZByyAIqPBLQzdHBtYror9ch
gRF3yrrL7YqpFBrCKIcGF/0qeXxKpSp7coxBr5ssZBwxlqwGho/33W8d5q/HEA3y
xcfP1d1/tWNGPKDieOZyihjctR8i3q0M+RcZ/Py1qYwpxPcc1I9t5/nxcwgtBPe+
A0hAnHOa7fkNwHLe6xYdF4zAuEfmSbJAt87l4MP9CTFEVCQcZip4+80nizNyX85O
PVftO5uF0JdmLEC3vdz2wSFBi2tP4fQBS8Q5fP2rmaSu9jHy6/Vzw1iOLgVbTSCd
lCjYdYLYBcniRkczWHUOj4N4yl1d1WZY7Cjzq3jAWKk=
`protect END_PROTECTED
