`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kiBRC9z9POjMO6fWPm5eDzD5Tb+A7hr4FPno5AuTnU6/kXQW9JUlFWmqpQ6zZPQ+
jRDyFiYAoOt8hj6huKhRMxb0Kwr4yxXyLr7qbDF4P4ZB7NO9xBHXdNmjI1LwiOGv
19XKPM8zU+UCwwqopFKF3a9QevvQEaumbrw7eZm8Yw+b2n0iEOLKofb9R+ANEen1
6qnry1/CWoeRK4+AP9ovdH/QRGsZi7xZ+7QtU1AJop2rZbbkGSN6D0RaYrI4GjHe
HcCAdus/pBUCZ52bvuKJXRMzsJ9Sqk/9NvwIbsAxoVs=
`protect END_PROTECTED
