`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AbgXSWaDKyeAZiNz7hHLWJMIopRAU7HlCniXgGpj0i+RHNjnTq96O95BazCCnpe5
C+gCYd5SaLY+moPpYZyojsweDvahgrFMsNqqtxJ1XTsUx1BR8syXyeKyvjIuE8gn
Y2OkDrZ6Xu0hZ5I0ZTXsXNLsWBhM0Qvzmse+hDz8KlCF7Yc+8EGH3D7PKPSgN6Ge
C2l+JgHKEbw85oC9PIQHlaEedXaTFeZ/dUhmH883Klq2qmap0aMeAqMbBJ2PQzmy
MPVJ3zPGMKXA2VxjJCMBFpP96IWx+jUChWv1xc0qEVmUoiu9GYMEmZ8cu6zzNR6M
jkFi8XbvS1VFcB1ZDjnytuphlMX98DAmm6JxFXT63ADzQWUQD3qwBtKwiydm2dDi
R8OqhZIsgnsWTvohdOnErqXIQS0j9t9C1pwIV2U66JqUctFqGvaQjpJqWqMvZ4sK
SbL5glEKUKtO+yufpwA/ZTpMyy4LE/wzIKzxf59fYqsuKW2O8xEV3uBs/DuOs3eL
GGUCHqp0L1HgKlNj2ZlmEOYsAQnw8lkkk2KHuhnjhPYEL+mz2QORfg6y1rSXjgS2
6xaetFbnN2q314iTG1uffWD/y7aQ/vluL0ThTddD5kRRtKCsqH0mKWF2O/i92DMm
afPfyRTwwDY3dybOBDodB5r+qH6GiAZmkY3MLQ3vl9cT24iXrOcMjDrBKhnx48Yd
DFVlmSPWpawE7dC0h2sndZngFb0/gMQFh6dU1hYxuda+meRYrKdzuIQGYa95VkDj
bt3KxpQZ34cUr/5PwccUQ1W1fRGEEufsleG2jPUl0M3qx4iQqdELXLfYDq5HrnvG
YepzSfPdx+ecTEl2UTWzlct2y/+USg1h5+gDLc158puNrDuad8DutZGPbAx1lfls
B1u4Pdz+EWVjd04YumlhEdjQZo/PTHP6nSKRQ6tPjeScFhkW4Y0zp2clAWIzFjDr
lFaQfvkwG3leUnquPTxUIs3LIqdpVEueXOx37xvcz/Y36gVYWPjac2gH6ajBQBjx
WNIO6Ddwg8AdAlSfgfowZDd1J5NtdKUd+G5IGqDSwBsmoKmr/m3JeiQfDbY347PK
FIiFuH85ANx39UH1heAHnj7HXjz7D5hGmS8+BYFzNpAjsnj63/fNBdx6uPjkvjJC
M5KRBcbaT0Y7myV8nl1v8AJgyQRZ3kAj9JoWThtjq19hKy+3xhy0VFDu8sSBG4Py
1Zj98YESrayWOEpP+JnMz2Xlznk82/Tl1F8DMXU7VHbKI+sfyEKct+Hbxg6jCM4K
jxWdsXhFrhThroGK7KXZ1unrY9gEylpUt+pyEu3aUgwFPSUwfPhGUwFmUXBVz7SD
nieLT/S95PVz0F03vvokUImqrwy4D8B2Yk6AFkYKrR9PM84qFrpcXWhafS0qM+bg
mWCxgczvyo1xTSg3vbcLcfReuv0RkQ9KclVhlnEw4YFEsFbq4u3QlKNR//DH4OcS
aZFDNaT0jBCl24IVLuHKn3S/fft2xRYZaMTE8d4AF4cmSkAECbNyOFgDeVzAUDG1
JvQFq+wTv8JKcsr8wy6Wap6e+dgJbLxbYDFJeUj5lNOWfBfB/q7ksrpNxqPNMUer
4Ni4spMpWHC1nvMcmwhTK6TUf1/frTigNChCKgdO0wLTDx/bfXBjNJqJNpz++HNO
l/Ms+mKehEjnwW2htXiwGHR7zzlqgpBy0WqyP9+YIqVStNpFFDJF4arlpAvJPgeg
CYq4aX/oH/NdO9g5dl4x3yP5bVX5t5UVX56BzNdJbCiYqZNzVE/GQcaSv/SXGYmF
Wl+sLtoDqJ74yivdulxGUKxHzCSLhUk8OFCjyo5uCwPRhPbDMIyXIx08oBTWiALq
mmZ6nGdotoKCtgEXw2G42+849YBA0DfE1btZYIbRNGgv43MdxtqbHjJIIU/uCVoW
pN5+iv2kWSiWBoW6wdCeIg2za5FyyhytuJB2cz8RJoILKSHCH7s9RjdFHbwgbgGR
nxs3vqMy87SxQIXTYXNTpN0qHzJfTEvbwnGrPz87URn6SF2VW1rq1JTgfrkIya1C
Gu2gqYhTK+MGSKLY0uBpewhkiEzZ1iD5LmqMlyjKXWQPH9x3/tAt/b+IGea8IEFx
HNJORZwsIUPicLzlQjtQGqB+onW+SxBPSpvFlKsYNNkt0HnThXum8KwhSa8ucKkF
R0KrUM4hbwnopIVR0fIjwb9P+BOdFCgBEPlT0pzjBTR8OWN1pAOpwaRsNaq8I1TY
V1LjNBmeIT2Zz10uTSpfkQhlItT5cKs//ttR5+tuL2Gx4xnETXWYs1iwElv320nq
jiSzqc9NdmjxYtloN6aZB/yemH1aPytLgQ4qkRdldP0SeT0nvANCKbvPbgA8pMiz
8n4H3LIMKNRAXb3UxznIpEcVQC/3qZladROJSEmWeYUdo4t13lZTQz9DrnbyAk+K
oIlSb8NJrN/bBAnUIaR/7wmDVyaOIyab6/goqpyYb5nJ4Bj9p6bkTsUlAMSOVH8M
ZzwVhcCC5iWdxKONtRF47+gHBq51Al6Ci7KIEA3gKW2RDt3Ij0FNFxCjcPJsz0fK
Ab+t9PaGN50Hi5iuGei8G3sh7GY3cN6x1XTpGfVdnGNwcAIctQrVzvEZ9CYNjedM
jUYKSanh+wsAbxlwuPyYpwfkDBvECjLB3xuSLjg4buT2i852eaamF6RQqj+Oq4/j
ShWATdsb6wXIhPhz5XqywQcy1Cpk8YE/LcZHLhU9kgdJoPxABs+YehOwcbJutgJD
GeaHw1QN/W+AkLaUpbXIfcxGoj5BwGAeRTtpHIKz4dOsdViEp2V/yDd70Ld3lZYn
r51Ra2jKXYrN1URddt8JNQ2ptoZM4ORL0dPUEnPPJ/7DKSJzzoOKy/AX352qTnMF
HjP9S7cVorUXxQMcwkrbgqJyieEOqZ9p3/p06clRlm5DQk7jvKu6lNb4K20wI1fd
6Hebzec01YuhX+PcV0LeJYMXtUdJ8nCI5NWPKWH6bKnX87tJbjMsTsMnbgK9YZ9o
LHUZ31LcnF7cvo0TFBMyolftVTYHC0kulScYy/w9ShY8jn7wncCOTRQJf2wq68v9
ZpS4WgYZTbbwQ/dufCZM+QUaK22Ti4EVJ4Vj0b22CB4N2WPLWKB8abzKNHNEMJ1q
uK0Bsmmb+fwMRs3NWLj5m7tVHHSghn0SUznG0kEittHff/b4HiBeyFVmrsM44jfc
8ZZeXjTfLn+i5JPG6zQHs0ZCEbxYPMZYGsxvlXq5xHDAmm+y/r+dCWUHIMUZAZCM
oKg7X4xBYAZh5LyaB5bcJfJUdt5pSqNY9d/CR02kO2fkJ9LB9SSrSWQPqCy1J7yQ
DvvgGxkPhsXzrV/vfIA1wmH1A5Xc2nKSmlSOR45nD/IigZyzQA8ywW0FpzZrbbEK
9J36gnSzXa0CixeFahBSUALTEjnKbvaK6VblUU/TUadcuNTZN9zE4p5TjnylwhIL
mp4vyWsR4aOJx2fbEqzMSadLtbqulyfTJ5WvsrgWjxDTYgpkHSTl8m+ElE21Idzj
GJu91Yj5+CYp7LmeOdnH/JXOPi6QTr45DTOatyGEVdLx3xz1Otafn9vhFuu49xAw
BmIpO+vwK+LqHJuiO3pDsZGfQ6xB+JolG5ysb2RN9bKXtIKI+XqW1+tGd8ridFI6
Wn1VNvEoHCnxFwbZX9WvHDqsd7Jzk+x54L94Jd7zmLNylVIZSH9MeyS8rZbKvIFf
A+TI1KVgxJK6UrlIFEO/4E8VzfVFZvgObxMKDY+ouunTOoXohnWRcec7UQl007EJ
H0hReVlQCkHetQL3YRWnmnmktIGrJG/UKO8Hbg5cLsjfVM4MWTl404/JMDPsoLpW
+ci/BsLXr19rYfkKoh2echYRh08CWxxXXXU/TkMphxiDnlgut1UAFkDFItXm8KkK
YL/en8z3nv0YAfOWo3rDdKrFYsUgWx3ptaXjh+bKVrPKyWXnNn9QCIhcj/9LQAVl
bBtXxKj9AGIurVvT4gpxAiyPqc2vQbr7s3gtpx1AB9ocKQllkLYUx1uxtKAAvTv9
kbpvHAK9j2yMJ7Dnchnr93pU3OWq+K+1hqxbqQjj8u8HIWHAzzOnt8uD37JloAtc
i0dqfec9ki99HqhodG5qHcQ0DAT1BAWzZ9N89sgasuzQFEYjP/nVnKiKzNRWC9Ay
rWNYl+Wwhrs0ySSK4JKIL2Giln04opS28X3lZ/ZXXEwLvRkL+ZGbS2p7CH0rnr5r
1CQXrGLDsX1+J4RTIffijLuQvjdqUDGzQUKJqmCj57usYshUJ3DDmIeRZwIhnNj1
JwVC7ygOg9OVYLxc9R0ffllhiG8zRexndn/f7wO8HvTseZu42T4u8L0JLYS2mm5W
GG7WyAJShdAs2iiOAjFbNn1hcmi7r/CWJcgzj6NgzUaRYI92F7fwag9ojTPJO8lW
wU+xRA2p0kwREzmGzcfA3p+RtqRqZVR0rc0ExBDusDUxRHqt3mHTWNt7cHTFRJa7
qtpixhOhW6jM1ys4u3BfQ/vVlmJVrHiBVjhmBnHwYDW6Vsj5/Wjv9J48rOVB0nwd
XCgSc1tJYIJVchNRimBvVuLEhkPjHO/pSDYZAPFlm/ayrklSreYJ40nsKXj4kiRa
ViwGLqRFHTbwydrBkiPYk/cPD695aonmfOgOHD0/ApVesLVOT/sAWW+BT7GlVyE0
L9zBQDPSdKiAIGEWtQ/koiLI1qDy62t4FBOIm6or9yBZgj+eWalLFPu5Cnkt6pLI
I+Oxbg1v4U1PJoNrp2bhBz++1ssdaDLqBOZPN/lK8r9KUjQmAhQp8lBGTlqTF5NT
x+19GwOZc3CjZpwtoMe+COQWAOGjXweKRhlkvZ2ZB8tM/vZ5W2JvmvDGFpaXNJmb
J6nv9mRHYP9bXybaWIWQtWiXBeNB6wKT1nIqAVVCIOk/XUvpDbeO9VzSqC1LEFe4
sNnvljpgq6knFtjZXHypGhjuFwO3fvxn/STKU0BzBDr2YQh/7mnEkrHkTI4PlsbH
s2rJFTPuNx8I2NqZ/2EBCvquxpKgOetYxCUlUzgoGUTpl3tyheagP0zOS7VliWSy
aFwVtpXIHap2Sv1Ty0ws42+143KV2O/vuY4e7/qZTXNXCTxu0G9tY3DKmuCRb+Hb
WW2Zuug2aHyvbNitIn/yT0JzCamqwk1Z4A5dGL5Gc7uezY+48C51g3QZBw7Fer7o
6D81XHWk8kYfhSj/0asscf/wx5vDt5ZaVMBgxzoITI3IOiXoBprjsSVy03zKP0OO
o7Egkl/0DwGe7RDISo2Lo49HypgM8m5mbtzdmauZxXsGOPJZ4gDiLGOlP7WWKfbU
zgdGVOOJp9R66nY/qhIRbJ2DAVcXFCKKXzNG8iFSKhKvIjAnLg/FzRf1ug17q+t+
HmNIsg0sji1hAnw+2/tSpoBfz1Kfp4wPMjGwFTapqHhUCPL4LPuz7Xg0F4u1/eOE
fh8Dv3ZOJba8rnlh+kN5jFyfdqrOm0ZbYR0ACbuvG9m2S00XPcJzGaiLbilyzOrY
bl3R0qBZZjKUIeH1p6TYTZhWE++kBG8wDBJHWNGPKJaJ4m6ibX5rTycRXhHiqR5z
umS8fXTpc/db4zYECP1RdU6tm55k3CkrS4SaI66gs4v9B2pV3X0+y8jH265KGvjG
1u2kqCviFFmlsB86i1S/djKi9szlGbJgPHSgxl9ogFSMDAkG7rs5IsJuTgh6m3gB
/7/ZjYEYrPfRqhan20NyedCjdGqu5fOLhkzvs7L6PHMzmAvq2r8uR7mHcBSHROdK
8ChvN7aoVJFIvRmj1SNzYaemKt2Ik4faBy57qQba7QrJjuNcb5vhGPz55H/2I9xj
t0mu8rCZEocBgImMPiLo5UfU8YdeCoddREL2X7XkhRyXn6aRN9QibsIs91EKpGEo
JpDchdpo8g4L98j+23SiEFzrUPyPXF00g/Sj2NGy8FbGTJpBw+mmsgCbWIKRdoGT
kuzODUDGyysHF1MoR8twR9CA9NUqcDuOwZzc4RZD3UEO1a933GXGJUkqLj1AtR60
rDxk7kgWxgMeeb5+LB/jph8zylQXA/SKqojQI+15zmk4tqRVVJam6X/XWJKybI3T
RcZkAt/2mRv9tl0D0ZpwWwsqmzhfkk4dDk3RveN4e9w4Biz095kx9mbAMCIj1XhA
50DpDljH8fxiAxiqitGGxEcQuyU4+moplewdkTN8d+F24BvPhpyILktLQRVe5Rnl
NpJ+Jj4jI11vYW73TUbQxRPiF9abbPYI3dnMscnTcALnCJ2b6cW0q+ItTs82SZni
DZ2k3SoqPj5e7txtw/5NZZ32eRmoGvoRoIrQOON8HCpKe55TVCFztTKK8Hr5a3pf
0NRjcOBEEyYHAokROv2Zy0ekcW1Jk68lW1mrqSjxSMdT4dt9wA3g7WIdOH2aUm1v
qNWexC8zhNDZHxhoi4SXEAYiU7v6A7pcqFcJwrnortnW1NY5vcsWFH8YxgeoCNJI
NYTpUlQzL8t8M1avB1B59QKllbbh0RybrsW6rzRsSSsB0xMujbtj8wAW/TZyET6e
78KaBbLZV8gWIF1crqDW6yEai1/s3REh/gH86DMbAxEYM/eu8QBxgDL70stgtXWw
GANLVec9wPJDrlgPJi93fB6N1P+EOy6Jt7zlmH4DC+Jx4D80SMJMDZLGCg6iQELi
xZiltBhsPDp/gYpUOOYtJKxyjnws7qlwD2T/7mSivcHpRRqpQfadS4HBmlRA9LUB
85Ip4tWkQWN1nfBQCFGplzTkjKJVQQLS/8vc0wnSW2VhAJ/0cvkZL9tVDl1ZKdUy
Uy1Ofpde6YmGHfX2ywqsJ+Yt0itZ6YDPQ77EIksbHXzMyi0GP95DlMjsri3dgpSr
2luD4Xg6qMXRX3lLYBLiG6yga1/AnDuQYkOx3qT0DmAt/NqmPu9PQoUlZ7Rq+vQ/
eWz0rZxsjbKMPs/gD8/AJrWlAl0VLvYdEcQGt6SSocxlLEuSxpIA1dpIw7umfCvr
1YOb75ePFQxpNZxE91tTOVmSWf+vrpXPt9U6AKLl3qD8NLUQDsIy/T/FIZO2h2mc
5IsD8DSYX5OLGKJfnIp/hfjvV9epWdnr1IqUVrXIhtKYhTqd7XCKk0jqDhdQjdgv
DXHU98slzAEvVWRG4QWXDZRNOl8NyQUOPCXKkStve0+sJMQmx/qPLWq7Y6MAvcVx
3wVF86oaiqfzQwBjDM/FsJyQkNHSXL2xDaFPO93xECoZmW49SenqIgOG081eMvxU
tQbf2cBKUjCUifep25iqKft9gEMIOX2KxQQmudkS9O4VL93LH0nUEgllX8Q9q6YV
Ojvglad4gA4HZmX/OTHi/bqr4hqDxR2Vb6dMUxtm73vSnCKt7BydoV6VRjLJvFV7
c7cmMaDjLM0I/Hci6J2eYGbOvU9RDgYyjEtRQX65t1fk/ouRLpspBLRYXCrRWMgA
j5MDARKL1gWu3ZB7pj0i+ot6ECu5ypZg3NlbE2N3lYxxqsZr3dbpqJFHLkPkq3gJ
7xNlL/FNi/xAeOwtAZvTU5BPWOyqVIcikXOhAaIVshT91xrtQ4e5q3bn6ye+5mpv
eqCNOsAwjpHvCxa+8gEtAIihx/VXSDMmGfxKI7oyJjR265C4iQASuELI7BVFQ5Bx
63hO688T1D+D43tbmiKo8kT2WTLkW2L5qDRv6y0c+VUSThYC7SsyU/CMnlKaVc66
NdacoquFG5BVmw3n3AqDXWwm/ZIPArkcijdjqbyXsollc7lngky+2mQnOu8u5xYU
RqM044KjTHYRRqezldNtDaxLGlNyV36yq7gLBdamvv1aqJ1IS4vviqtBhZX+KBrF
jvS9qihT8jjVYc+cl2kyUGjQjSy21u7k3AjM2wKX0JS/gomrYOZxnSwsT9GNMCxD
5vx+mxzb/2Nzg7f0Z2SW5Q5dDx5JvllqGukc/khDPUH+ObvJj8gZ8tAgj4gx41RZ
/cpdEE6nqvOkJNfXie3kTYsGWzaBijIv9rGoJDqY0rU6UQ/rpsS44lPGdFK3XnuD
Xo8Nrp/JxOVw66hqeipT/83GrWVUgTrpGwG1cGNMhFKk4MJeF8H3KvzWfe5xqotj
Z5gl8kTyKwM6jAcXgLjz45ApToIW7CNbPG0wuqdyZZS/inM6CYU1uC5ONZjn0Cx3
mb/G5A+HJRp0vRbPDBhRYBIKKyOwV2o5VQ9u034qtJFAX9XdPZ0vFxi03KkJE2lg
XVhzexf24JyBCEkqxfUjVpb5KLaHTJi8UdAJHHRakMRQ4cNJY6odnbdtML5Hotue
mfBAdD8b6NLCa01gRh7VHLyY7LUVRXz7q28Y7wP3H16tbP5Qov1bAii/iXrm/POw
pCgF/AM2z2zRPqbzc0Frt/fMufcgNzHGGhu2Htfma5VRAtlEPjdhJyvJ1BGTW5Pv
MwPwseh3tiyo+vRNVCv3Pf16j+t/8bgDvMCUZmIpbEyESVkwQK1Lh07NMdhrbT2T
V0OXyimkuIkM2DJmurWqiZB1wKO8XdLsVE/EUksoOAiVQOMSEK5xSuhRABWgaIGg
aktFiD+P8oQi9RCffLlpvvbuPYYk9r1qrvdSYAZmLLhVLW1Cabo2K2oVe5ewyBR7
Pqi1tkZPB1hNmgNhLsBdCyXECEBN06w/TLo7K9sr4rRBqTbJxim6fqcNasbc6sjm
JMZBXduoyEuVcZTRVtOWD+xjg+KDFOnuiuPYPkXsaRgEnah+hhqUFFkVQBIuYMv8
vqhV55teYiJ5QHrApYrS/0hYUIjyqOIY/v0pDuyFyjYicBEyX+JG/uXk2sl//oYA
GcAL49L3aypLQLEtnkH+f4F2SLaLKc8dMtcpXNUqVzl9lT724+lGlsnRTY2sgpll
26T183UxkYXG7YY8Wz2IBtZaQFVH5F81QlvEZLvJzS0GVVOiSMIA1hEa+9uJJvOd
urCQ+y07ANYvD09RzyCcoy3oTCFlNEolf5rl+17jnjLYzjle55Mt0RyyqGOi168w
hNq0xarppwvteeN/ldW5FxKmCD4ktCsLpvNFps27Ypq/yToEXU4g7DPEIGfmkC/+
gs9NK9loRnWu2riivi06ZdpxpnvhEmT00oQ3Zsc9ofiw21SBBQfjXaxBQm0+caT0
odELujG/Q3f4nYlTcgtluWkIXpg1EqquDZ/jthxvhuudJYIfH6EqQ/XGb1vxZFzw
KgurDOYGYI/0nIppm/zYWzzoyC7F+9NSocYfW9yAsBM5bF/Je99s4l+acPYPBGjw
QMJf+0SnaNtX+1YlG+GT7p4HUeDd45l0WGICRHE0IIN9eUeWskNvmA2nogd4MLKW
etM22AM2O6O65KXc7Kf5sLBuJ9TaUiWGrH50woQTtmPEhfUGQjf1wCVZ+Q3inAZV
b2Jl5Wzh502BCnYNAxCRSWLQvOOK1aXyf8wlOhDBlMPoLwboRbw4Kq8r/aZ9cJC0
3BwAHjTdUlj+SUKImIbbvYdT0I1lXB0OnGiwEF9Z9SZP2OcU0q2HAjsgQ9eupmDu
B3+t0pxZQARuhOFqCFIalSIaUNRUivjeLLeDX8Ym7t99PxtwAqz54zvk5N8QajwU
f/AYzUDEs6a2MXalFDvg//oHFdbHP4P0dPeAQTxT9xE4f77+9tpMeq2+l6jEMqOf
daRPV0zlB/RwXJrUZ8E3OyYGaPQl0o20yiAGfAB46ifBHWnuJkUu+wTCkgo5lxKb
A+Z0gmiqtWemy8DRtfBpt9Ur+Wd6hywYxvsh1Y+9DiiGAPO5pYdVxO/sxwuHtZWn
48JAOBq/lYQ5wGPT0sJqKVTcNjcQi/ehXldAKmd2NWqvLVNOxpg6vOjFthmdYoaw
pf3AKUjMOhQn8RWYfp5fcyh+Bjka0h0LHcOTKwNvF0S2ug9qh2AfnjcAUkj82WSx
sKMTaT/9sD4NAAz0bFJOpuSz1lQGLzlokPKzQvoo+ZgrQgGNUutw3wG8LVAX/cGG
Ik2BxmIqnqRbKB0mh+6ddYlqcEVE5yyx1aQqqpZh/NooiGmfFDu0VWAuMLApfTlK
JY3W29fXzDR2zdFoEFlhjbSuJOOeEGGKwETb+mdQlVQq9yMprGC3B5foos//Jk2T
iBaC43RgYr3PKHb+pVI57ACSipwBH5E5TBEY0FkWVINSU8Ktt6lq3omfLq2ttIrz
wqG7R/boy2dGbdouWNv33iVQ3qXeT08RiF1RL+R/AbwZPBw53wKK3RkMHB5r8w3p
9sWigxSFjAN7FV7HXuuw5T7Us2fqJI6vJfZSgiSDtBOEBxgrztzS5qpox6m78LfU
tn34o9DquDgslxJcxGRAuT604ZnMutIdX3uZ+DuCke3PVj9ISWwBE57/ma6y69SN
5aoq7YtCtWydZxZM1gPmO3MHVtBVjCC0Nq1EwDguzeV0e1hdhjPntyW8w0fYbw8e
62LeNA9dI7fgfuWb01nasybgn1DPtGJiyYbDa2y5PjebGC+dsPfl9nxuQaR54zKp
ChroMYlsAuR0F5ktLHZWHT0XU6VEq7Nk/SUFuVKY9Eg0NT75TO9ewoGB9rONRDrz
1dU2Ts4NxqoCOt4nMizS9+xNTQebqNEAA+9PwvyiWCpWqB8TSRHVXPQYdioM1BlC
3xluaiDJ/X6dC9PysSNNRyIQVVAXsuHTInYtNdK+2JA0KA8XNjt1V2WyXQpgWVPe
Ataf7uA+U+hrV0ABAgan95BoLYuQCI9X1aQNk4X7GR6pLg+v42cRg3NrYU5pwICo
RHQxnp8w5RDt6Fh2M+Nmp7OSUul82xv6LE9CrLcSmDvtDB/E5wudGzt5BxjJzRWj
CDwY3CyiExfWdJieZydlm4UwTPAaK2MWaaX540rGmzYszAtWC0j92g6ImE7eSBxE
xqm/fYeRJb5HssLzdefWY5i0QQPn3uaoD+2tvTYL7/U4vAdCJ8EcZ0ZVXo3ofweO
l0qQm1EpOl4Dh49NMT+5Ka08WfvXEjlab7+/OaKjqV3AfzzEXfLEVpAFyMBlav0r
HC/rlwzL3TJgTOtWMhvnNsxzlBLY5vKYLaIHqCL6Ttj8TYyjzwggR4oNCpfjIEFJ
h+KnItmh5yjpr/ZHD/aOgA==
`protect END_PROTECTED
