`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V5cx5EwMpSjgMNeophWkcLR/G0VcimgNr2fW3RlkgiprUbLHkuFapioREuRjW67s
xDvZmXeT/KDIUZCvP+rpgPwXRMD6ccyKgvwZBliTkyely3zPvszFN/3Epm7AirxL
N9IKMfJXLRmwtJHgjzekuJKK25ogr4pYjZ7he+q0VwB1Pt+xdRKe7OGfbYNSpemu
jDuFu0nQc7RlapT3nJuoPD/4/cRJpcBm2Jq7O/t9r6aQhQd7qidEUo5QsrO3lazH
evFZFqPNB04XdsSGS0+Wv2ICIEfasfouzUF71ecywR7RIa8rnKtcgoT+jolnL5VC
tZ7fVLJ9eLI243kMNgaT3qWDryZT4VnLrselBHH64Qs5JCOtTwVsJG1Ko9jhm7oe
sQXY5rtd0FSqWIasGJUCEPVR8Sr0O2QAvF2Mdo+WwF8UrgfgnfaBsJzg2Sn7Ttq4
QrKyCiZlYpV/bZXHZjd5SunprjtNYEKZhNHJe84lwRZLJuR9r73KwauYFRH++KWy
79QK4NVsz/M4MYAcDmlepoIDiXjYOh0qGr5CZHOcS739zMAUjQqInFe32GaKM3bk
Zs2hNHynFWam90um8oVJekNxf5WOMeWKaOOCmKsWUlJJhD4C6Bz9LIFjMUsBTJGS
bg94s9CpkBFxqCjcWRCmov9dbVCdF36QY1ay+Ch3ZaxwBfB4EffPCzjT5pJi6N9A
2wjGRVmP+QjRSMezCK8rqS7tZzuaJewlx4DAxxW61JLllWcZFsDwK7OtUgLPLogg
R76IRmgif6GawLubc801lMxvvvHk4eCoDV/5g5+ZOqAtHsuEc5Et9XWK+RyQX9T0
`protect END_PROTECTED
