`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pC6tuFq3ufs6E0nupFHQVInzB4uoNtcY3dwtu1mauNTEnOIfHxonR6uwMPB63OS4
jkup4M+mi56AySZpoY034AnLWCdHo7ieqtl0B/ah25P/oJzv7qKla4P5htsg7C1X
uC6BGnsI/9sYBZIuXqmR4+hzmXNFz1RuA1l/ZghH2+gOvN0qlqtvj85my6092NmZ
kIkzLwRmprwb/5TK/Elp9WiV97sOkx3RXVKWaw5l1oCBAD7MQX6qhEdZevSO6Isb
CO2IHV+1zdPWhTJzcZ0im6S9ujMOscePBwcaMoEGu4IsBLyk0hnSBrvnQcy5pMKK
3T8qCHrJUD0tkDdx5tpMAL/RM/tpkG06GJJzQjJNxdrQt1PxqKWyM8GoWOO0C5N7
WZLtxldsGT4rctZ5vMi+nGE+FAwsQ4hk7g+bdEB1m+AkuYIVtxhv8F6Sxqye5amw
3naAn7hKKabt+r0ytezKXlsLoSoRSo0RcATIbkmCqIfi2PAqsXlI48x+FwxhB3OT
KQFLtM1Hy7ke8BKTz37HY911SfoU1/IuUg6MtEVk77jPruqI3a7cqhX0jZAUidah
otlp1VzmfZBlFgGrsfuFPkk04gEYuj3EuJS34pqyQOhiPMl7HpykJvzaoG+N1dDp
`protect END_PROTECTED
