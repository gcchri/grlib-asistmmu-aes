`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZB5idJhdKW8eOZM/3atm0EV7tIsi3BydzEOr6PPBRDxkcx9B0MWp1k6iv2aMJFQu
/c0Jzl3LrF33s2ur+WBfMqUbnqS+bUAVlIoDV4TJt8yQ19Lm977N8phFxhfems0J
5jsiukPQHoxsb78e1XxpZOmfa3bXMHoRxhy2CDEG/nQxbgDBIpJhNEBytkxcDPJp
E5JRb5fN3q32P9PfpzKd6Xt+Z5ioD/XDlRSxBeRI0qOMOUmpvRFKqZgXNT/SYR0V
j8rlfM5ji3upS+Uc3LSb1Aa0kHepd4dfTEnuaMT1N1fiZ+3dpQ5PvcXcpqLv4cbF
1jRC+k+FZU3oKdJWh0lxfI9Ub2g/TRm1FYpm1eefsviTD9SGKL+eVvvK9ZtEla9g
N+QFaQ+oxEmriGLvNqw6RRxizuLgAydjG5xDZoijdSa5Iy1B0Kz64F5hVRDX/yL8
EzZULA9xl/AMaEjbryJaWkqo51feOYMaGsTuBN8GL9VOzI4QLV2vlaYJ1j0WdYIM
nEmcaV77J57L0iaGH/1n/BiDM3Eu7k2VzRsOpyeJ/IrEqFHwEMzy6+dShYYutAsq
PSuTrqipehVMCgBujg7mRaQcZJr6amZrYgHmGRwlrePCmN5KkvwwazTVznQcVBHW
P+vNSklumbd3Pn+g+5mwg9+jOyTWKBqFapb8a8iDxuFVi/d72qomM4ucdMbW9jmm
QMk2h+sLGD46GXvw6YoC4Mk1Lg0VN+OTS2kQZrr0GxPGVRzO5Kxzy9fVek6D6rYo
XKVWXUs/M1g4d6pckreNnh0Qy7OZpPidEcbviTJcCy+NgQ38Nzt8YHrtboqKDc8Z
adc76oApbOhPKLsGuB5Qg+S0dzirAn6D8tQJ9orueIgEYB30axs/Kc3Lcwn5n5Xr
eU6utijr52ZWujdeFcGXxY8YRA0O3Li4DzdsMfZkU8Tsne3/A9/Ilok8o3pxKhvT
ssNRkheawRXurJty4uItWlCiYzeae55f7wE8GMRcIdm5OLFZ011Pm0Sx6OC+ogiF
`protect END_PROTECTED
