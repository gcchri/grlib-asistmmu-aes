`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rze9EdqB6W2TVI+dbstntamnHZGy8OIwCnxORGENxfvjXnjFoULPgXgMjp2WmHvm
cokapNvnLHGeBmoKpG5xnFvwUWsaR5EQQhiKH7y2yaxdJG+QRrFiox7Yr4l8VwkX
yA8k6qYwMBZbVUGXZbIR9m35tMbFdfG4QSmrABtZBw9OCEUPbXbl7L0ityxyVwJi
bCHsTxJweVEQrah7eVF1LjhK382FiEKOlBhO4gwJBj0Tf9L5YWSXQ0xrLwyhEyPa
3Ddslo60K6TKQrmCXZP+KhGSssCs7ukEUTUfc1h/1HG0w3NknEDQR+IqeSMgWMNO
Mp+iDRtdm3qT7ezdVPDcOadAqpHhZ58NW4VABhnJQARdpwNOsNoBp49963JutWLJ
expaqDe+aNvekhDVzaXrsngbzYvwkS8EtUD6dSLpdN6cTRTckiQSVj/oMi1VRlVx
gE5nsXUDZwlqTW6/6W67cISOLssLoJ6fSjdWOotRbO2tk3/hdCn2sb+HbLV7dDCd
Kp0aGrbE2YDeQU2653frMMWYuNbVlJaawXCYg06+FSh+NHoKSHlTn5CVUjMBZFrp
w/MtWMpC8nQjB8CJk0VyBZmk0ZxoLjAxqYcivjPgr4IJQT4RxRzYCUnWGBwNy/uB
+FxDFDjqKUd1wyb8vBNdIBVc6NrslLRD5P0bvH+oCspIYuvLelinyPMFfTPA+THV
Jwkxe2jOymp+w5iA2q16ud9DoOoAo9CbmgdC7U+BjSg1DLc0cLiW58y6qNvXIlOB
O/FNITUVAj+FVMYHQbr9PJPXigCYgI7rDRoF8LdJZTpI07zmCHk9xFp7OJzNgv2L
jG4GvyW6zP7kHPBjKNnqxquniG/WFvSGpFOmLQZJccjKa6Wg+mKRQkSwQXX73Sgy
SIg9LVGvNpXQfNslseoAdFkNoTlsX4wyyZk7X3qFeMctiBw1rtptVdyfp9/LyaVG
BFpRVL+Mss6l9lpHC55IYkZa2CxAt3vbO8LkuQoDfY6FGkc47hbmqLboyQO+m1c+
5b8PemYfKTaLCt76QsOLYrUrRYiI0GApz41S8Iur52L+26acoLftcIWioxCazMlP
pC4jAOiW0J2F2lr+Cdm4qfxQRSp8l0/KNNSozH+8uOslVXbASxPUy7NdZIZUo6t2
NZlVFdte1reR1exBrMrFbFPYnTGtPC5igrbGKV1m6UL/W2Rp0s6lrfE9oW4NB03C
lA/CwQOhkWBkXGkIkhkwGV8GkS42B8a0UUIMjrFNze337y7/DKPddIym3lnNqKrx
uwTu+QSCLJRMxUJihFbeGWJpMyDffTYtfr8LEfee4bxWgpUco/BPS8OMRKwihwel
9MTRYOCXH8IvLhWsj0oF5W5Gnz4IcQTcgbIKl8tKX1AVGzGVGhc93RzkyzpcVePE
mpeoEhY+C/Kp88yqwufSASjf9c5sO/PVtqEpqcNOO2TDrMFQggEjGogxSUdDN+eb
/Cqo5REmcqOwhsgCUxUve1ztn3kwDBtT72OdaGmWznJq3y0/CvSC/SpVqSPjmmsM
Nq603lU/iF6thMG0Roe9Tc9oDogb92GPQKRDuCb9FOwsy4mxRnNdyKnl5tyx4D4P
VrNy8nlbb3kO7MOAXb6/J6sxFKlsG3xQMl+zyCyUi2I/W75XvFeCCU49ia7wWdGH
sToI5jFqv2aW00cw3LqQZDEZWAZ+cCsyU8jcLeSAZOCmglzeCUJXHZ6wnLSgTjAY
yvDvGWA3IfdjcqPNlnasSpKOKysA2NwQWeppk9gkCjk6XVClYAzpYG+COLjETdY5
ZFm+KBwG5C0JO7tQ7Kn3a+RzIQiTpX63voc+1cuUSCP4skQKTuvLQ6rMjyTpN7rX
F3pmT63d/rAziPEyLQY7Meu5nVRVj9y4foe9ZyZ4WDDF3tZgqzLFMtAaUbGImUdf
O+kGrgYFAX4HA81yeZy7gwhccFAbKdkddYbFL81rY2Qjof5zy/hKe7/kx4DKgPSY
PZ7zWljOBJLOdN1ZhIqbiNLnEnxq0f6Mb7ZTHswT1yPnxGFNCjfAC9eQVmr3auro
/J4qD1O/YByvP7RKyFPvZm6WgmsCkE8RWtzU+6p7f584oGzQhnmYLOmTVhyRTYb6
V0N+BWo+yJo6as0CZeBqLQY1znNYpkvzvcIt/wjRv1LhDnpTPlI9X7dagqgm6hwf
HL34mD5vfK7f1H/j8NynTdLXzzkITOsB/HBc6u9tQQNopqgNAMWIr0D1JS1AN80g
ho8ORxl5oRYfLlhKJeMmkzdxyb8PEDZyxeLEtoKmovRaRXYYmvfa2qcGGjswty/D
EWIPe1BcdiaCeqYzNpEmlitMFOwuSIHE99eHLcv6b494oARcwxHcGV3P80nrHBoz
j2h4Mxizc/+Y6nw7k5uXFhhK1KNXXlQkY7ZJD0MbEro5jmsrjhQLHqYugo7w7IZr
0jsfcZprCVcrzw4/0qKIzSiFsPLT959UdguGPIV07qjxUiRijozX1WnjUIOW4fpz
ntmkL6hJ/LPazQV+WXkddTQmN2V1J/h1L2ZrEPeLpCjspNIDMI+XSbsAzlipkKa/
78VPPnCMroJkV+NyEHJPXFrds1uIzG56m5mDQVWBGVzUnzZsf0sRwLJ3ASfFvnEB
DRaAf5eOT6ycnewG4Z0MxoDpXi3zjfkR7a+cbdmYNXu8pyJGo6z384nziOs2mcB/
9q7IoPRKAXrDbZfKxWBWb8Uy3Ml71WhE2CNp35GsiArcPNNMFMPau33PgL96RQIQ
pY2oZhxtw2xuVQY7HVk47PF2FS7r09W6Z8eev7l9TbQYkWL5A2kPwilUL6Wn1oo1
/19Hc6JlvU6KJJZd/24gRCVRku6WYCk+Zfq1/EGqqWJ4dUIzQe3KY5dK5adOsyMS
QQ6J3mT7ojFhDUS6nWCapj+Wwa0fyDF3JkQkP4NpOuY+w20wirYy065G3ASJ3PYA
6n3Za9ZdCioipXddIXs/79YoV1/V2UuFITPQ6LkR444t2TaFSkxA4osSzoWke8Ar
9LLX4ZEw46an3B3t+1aoJuEdXcoHv2gJaPrz23km8SgIj7YRp7aoZKwzlIiwdKp6
lzplPkFz3DbE7e4VXw4s560JUaoWW/YEdOv5HF8kETex0b/+ExRD5JYYd6ZjqzHU
eXX8wnjG+VPC3ft3c8t7zPX4bjh01fAK5GK5zkjqMaQ875ANJthGAPvQM2bQy7mb
XfQ7yjV1ulLjferWRGHRSjLO0JhljZhJVgUqsNZU7lNMlNavIA75uU6vBucpbmQV
sS7BsLAvdY8womK/JFWY4p1ZxO9nUh7et8PT0LtMRnHRRBPProM77T51bcbh8b23
ZCMLd45X4fhzi/DoaaC1vGBW4wLoOav0vH7g9KtZOH234mBDMuuLQJlfkmTOpO3x
EC97aibFrGbVXxDKs8Obp//kBelLDJVBZMOmSkDyzZ8Vr6d3KebghjVKmmmXJIuW
RqCtFW0kpfj5UBe417+sCDz/cmb0gg5dFlTbePLLtQqwxPh9J4eF0VaXiTw0aJEQ
7IeCvApyq6Jr6w/Fi/6MkNKJASwe/pwa03bKqebhpgnsQp5MtLkQPSSrt7cZPETN
cguYJWRYOQA4dPKMbjubfYlqb6s7zHvbQdIuk5keJxDPO//HwE6vv+mJfuMNwM7c
pjzV6VVxsw5naeyQkFCs2dRkn1ZEzpXeIMU6B7o6/9xu/XTF6ZxRiSbaCrph5590
LRTuA02jNAmWKVXx9Dd4vape9iMSCI62whiHAZ/cA8IjnZWE/MEDdPuWIYleRzNB
y+xaosY08Ml/r18Jy3GQuxxZTosk8+VyDmL817yTqk/FzL1meRI1SaST/4JPkpGR
WsBErMp7/QtbLASNCehjomPir2lwwgZ3/Rh2S2OL0SIpK0FSDVRtDVrLkAaSusXR
WGHZKbREY65sTIgJ3tP7e7vIaPevlbsUhyJIyfu+OI/bkOQQD/tIsXXzZKOSPOtT
xJQnE67056AUBit1IKDh6RSJGsiLP6LXcTUlbiGG4ftiG7razvQzZTGkc5a0Wp7C
kiUWZeN4OgOGx7kruHIczopJ4NV7CaDDcs1goph3Umb6/pSftqWXfwT3hyE+oU3J
YAQks9S3AqkAK6lUsBqlUUkpWca3khjn4tLKde9Qud8c+pctUWioAlRkdYNVsOfS
SUHhS7u74Z7/UQpVXdWpw1LXt3eQF/PJzyE+8hjVlMuTT8coa+PQ9vMWI17WfaxD
RXyLLzzSq98JnlWb/JWi9cog6kw/kQnqh3ygwnHS3OqIQhQOrur1fsvKLDJe9RjR
dVw0kOvknravqPN/Dk61UG+HpjwOE43MxkBpNo74V2dtGsQn6A7c0blvPVCAy6VE
AhYkadyvbuR/z7LvGovHTiApg9ZpJaGOFahcdhIeTuXxwrepROagG2ZkCo/NdZit
rYsMB6Nib6hhgM0BEALg/3WTLxNjwiD86cmXoZDJvpR8e5HuaBgL38BxwmheG4qP
Yh3nhc1MSs+VmPso2NGTlJly1N+cKr2rVx+F9u8ut4fIBlGgstYRLZlP12gBf0YN
Nw7/UO3dff5+2g1izsx3r41WL3nqusex/RB9NbJvBb7kWOqYpTB7lYq/bLYwzwhW
cux7aTdHFIEpluYt31My5luN1w7JuJNGA4ulDmnojT8RVL5MR+MpRWvrFkSIaKyN
mBc3HjGG96u6z7ODIC6EKeOEUUBIrG6QbIxap3p89Ui9EjaGyxJLS+4/0vb5asEY
Eb4+TSiY+Gt55jDPrBBVgsE4hrb2OrYbNiYzKznZfQt1KoWYIItQ8S2AOyoX6SAi
OIbsyWXt6V1Ww3rjZlSwPgZHCM2VYsLKI7z+J8hoc0V2URnXbj27UmaB5GHREprD
qOH4FMor5YsQE7L7LA+NBkIBAaGq92e1xiUzYZzAHu8=
`protect END_PROTECTED
