`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x2mLaf5PsUxu/13xl3YyL/BiuSb15Z+MeJATK2VKVaEOFlCITTMcXb+ilaTeGXI+
DVs6MCphbibHUhmi/7TQahsjUSpxEE+hlTUwwAFM8jVpDm+3ZadfagjkOUtgQOfB
FU4oB8qjm13t3QvULXNzvGjODsZd2jRAC3t/pKvYD2iNA6FjsM6n9NF8MU7BDiac
LJjTyXMZMiw7g4pG3v7u6d4isQ6DxPBJ6h6F4jmKfX2t+xTk20wMnJXBa+sZmyWm
oX5Za1SrWB+VM13166Jr/qboKCTLUrEfDvlLG+qyrgiqRV35+8tbiz6qjyWwYhAJ
ZdDByqwmmqQQjmpdkEKkrck/mi23iyLJ+Ia22CQ5I0+StoGbeOTD1dnt4RH6xdYf
eQX663wl9IDIG7il56UeCHzUXXevYx8yYAzhUiJk4EeuPqTDizqefjKWyYwb8924
NmUi8hKYxTzYNZW1SUbjRqtljfx3vkTGI9ekb+J3Bus=
`protect END_PROTECTED
