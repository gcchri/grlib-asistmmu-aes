`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMq0iK2sxaValt/wiwKXCvRbj1GM9j9kSWgxDclKr8YFGmXrBVYt9aiXMa1j5mX4
8rjHV7KvE0jc0zEYzZhNKwniwiq2ZGlwGvLMG6Ex2z5cjO84zcrIHXv5/u+2Hlq1
bN+t+KgFUzkDNcksHnS4IoELwypK28gstwRG5uefzM8qQwnJKmbiUz6X2urFbTYP
EUDy5DHM/nEK+Z7FnxonaNDeRRvzlKodOYVCoyMgFLIGZE1XhIMC/AE8xpLcCoaE
WGG/fn2riho/+HXTTGJM6f17SsEYuspwqCG/o0TpS0nGtnYONFlMYGS22kPiYfng
80W/SfhCAJKZ0Br304Z4AA/CKvkARON2Jm74T/o0bPvijymL6leCfT1ksPhU58V5
J0SLvvcV0Q4nQ4fI+0P/kidZqKl57Tg/gno/eAlx6K/ifL51Xhe7YSjVPtQz3HdL
CZBEYenWSmq8MGzrC4bZkW2dbrkIBQLDVxcK4nhAzWqnk/R41Ch6OLHnKsNU46pQ
lNVhCid1n9T+2G6Uu+HSfbfOJUxHedU0acUYBjE9qzklA7KIGZ1jKEfxPdhIdg5p
TtNAC5ySlii3Jg5wusNe99mkx05W9P/kzqDwqljduCY/21cLhqrFwFTnweSrC1Gs
PY5GRmGnOMt9MnMZpaUsgSCnKM8MWskgLk/zVhyvSFioshzvL4B/F73fXaBdjoJx
Mt0Ud/Z+UHkTrj0pwEV2hUW/cf7pmg8I0PBV0oLD77X1ealRSWBV5GmEsDK9kW9h
ZOAyexEyuT50vL9cLphG2mkRY/52F+0P6kLE1zQ+Y4vTx2fhBpXWKvOppH6X6kaC
s0VSefPLM2fPn3jQNfPwmoG9dRBf8OuaVU/kB4CFJubb0P0wcBEhlMh4ICWB55cF
jYTJM6mF2myOaI7kojktPni65seWZccQ9JHvKzvFX9eQckutzQjT1HtTG7C4XJov
FbJM+b9xSo/5H+jG0/Eo2DoFbI51WQThf0Jm1kZg40GsGg+P778VGDxonjFTceZP
I9UOqQ7jW+sgIi5E85eYj9u88m4jbswbt1KPn9xlL8X5OrRPql96P57xbyGg8OAt
FEljp+KgCth+S3muFkdz+meU+1+He+aTHHXNMy812eFkXo3vokqxxDdZ9GysjH0R
sSbjfcU5ZvTsJZxojWng3AK/zraoLK2GMtVNuOKTB+sG6FRF+wGZPQRRJS6xymwa
itU/FQUSO+fwkehLsft8CTEksE5ploxH6u1bFi2Ka9uXC0cOU9JOOw9o7IUCAC8P
X+cgDlPQ0/1boozwbox8Et9WDjMWIsZhsVFbVtbEwFjYkUSS52JQ68dF+yE5dSih
9BElfOcgG4RBH9FemlWXbvLfps2PrQ4Q1dmnu5gZjm24CxJVSVkbI7UsgVHLI0LE
skwrmx1M918Y7S4LD7g2+OdJsMh//ZSLf4iAWxxsXFz/LxjcfbbSirxS5VV3q3D+
zN8rK8NsTv+8ccUIa1qG+uY8p8kadX+gAntg4zeBE6pvPQMkZfpJ/y9vdlOinoUN
be9CJsGc4X+t8E7KEu79vAaUst8qg1+fwn+N91eWBkUO0AAGMBJQgowKVPYZt7iV
fV7JuYIlyGo3ZUVgM9qPJKGirzB1yZ26fr9aCQ4ryeklU/gR3hUOpdfPdbnePj9V
vXBMBxSubSbzQ7ADMGLOlRQXtAD+ruCQMZ+xDDUNY3Hza9aTbRzuEJp/GnibAvf0
uFaogDKjLB+VZNb6mRPQp+pMDrAQCP0b0op4roLCX4SoDCL0yQ2z7WLudRlxYJl7
L/gNqr3XVdngDFJsMJLoqhlzKW7tVdUzoueUNbsxty0lefwSQK7KGAB7yjrZhiGQ
Nl15PBqxqmdzOTQVzhQmh0qf32IiDQ8cf6li6Bw+k8M=
`protect END_PROTECTED
