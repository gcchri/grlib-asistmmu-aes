`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t5XF1kXjE/uxdAPQbftUq0rGjXDQ7XVR4sNxB2ySyBRye2dAqgxB650X/bNLJLuG
+b1JpryLlZEEhIe7uZ6ULiQiJHxY/UKb25rt6fM0xV3sxXBEInRVzxRNicCvBnQh
Jc4T7mlvoa0KYtzki9gTCaw6fTbiBZ2mjvnJo5i5rGdhPbgR5y811aY9ivuoCXNq
+eimx32LnQmVYXrfRkXMqi1aXdF7lnawKD6JGYhDBIyxzmxjXc7tJd044nqE8AYx
qJNikFrFUl5qGGWMrFT64BXkn73o61Kl92KhObfULtHN0+qwG3fVImbDaBXJjusK
b1lteGfVvHPA1M/yRZawfrrcBGNtc6TOlQZRE/QnEXBMQt0TCqdrdC+D2+3g0fut
N66Q+wQJzX6QznVAod1VnzE2aA1anAlcEb2osb6IfVzF9zfsSwlRZV1f6T02Ezni
hvRLhQMNG/uP0x6fFFV6XLegi4Eg8+CbntWhdNN5U3riggMa3bneaq/7A5YuBapQ
40Cau74jiirOAKQjsdJwbOnyrD2JP9AXAfbyIDdOs/AJh4EGcm+PUcrk1e3JJsX4
H9CFA9uT3bt2kYkepZJjQuI5nrvx8nBpg3aqb+hlrOV6tCynwkbSnCgTgSmS/eMT
q5NG6TEEBpNmMeNPNg5S2zwxYXlz1bL7SZnCBIdm2di25PsrtWdodAi2bBYGlwob
8+lvfueHLmT1LYmWUyqjmFd5dOg50+3f4eOQrBKLxdGb5St8XdCCdhz8izYMLkAH
B7bOFzFw699srNVnfkM/nwnYTLqarFKWETbxOOAogBmnZ1ZdSbWSazoP0fMkxzL5
igNTlRBVavH0Gtwy/PPnGztmIz8P33FQ08FAWqJuBl43WPAk6w/C1eLrvbzKCOVk
fg6bA2i61sC2//uyb56DlbrFoPnKQOlzw3vRA9nbeWSACT+jHk4wWmXymKq0DEU9
rV3iq4xWjgO7Tnta8aBNuN+KXEBzmUEd9RGyrEAJJGY3LmBPJkm1A/Fk7tvxhQ7Q
t/oafMEkKFmT+1foiJrGH+VUEqaN/L22809HgzJ3GbvkFJbyibLl3Ge335CzvHmX
F+mLn9su2iCOUTHHC20IaxAKnYb4ZOsLxRPGPsZmqSSlkNbrxfPhLjZ+aS2+b+4e
0kb8Bh0AoUcKZfuYV3D5rRPrEU1+vsWtnuHgZ2LoUC/9EbiFDQkzDPRqPEjwjIoM
LSp0y6VjQqt6Sc6GQ7qG5LqdXI7wx5NKY4UYntxwRT8ou/WWepVC3CXRECPcnTDO
cPyj2DQ+/t6+v4lfPsfTC/Ye7W0fhzGRvbH2Hgh+S/XUHFwnJjlhxOslY5t+EpRd
HJe/Nfoa7jDnTaGPK0WoLKXs9vcmmrp6wqL9Jx6KNJ5Pd0vGyt3VGjQVCTj4Ysly
vfLDrPTlOpVyruu21bro2bEKD9O4mHRzY4/sGZR2umWYulU23I9DXLV/p+lQz8M7
f+jltH+U75wkRxdM3fW03VvlZLWWn51zuZbnaGYYRIJ+WWrBxa74smCjtiuoIn7r
qkyFpg+1NjbS3MIq9EBofQvjqr7ITex8FJ/iZFzzzlKM/sKNOq+kU12XM7hW1BZi
j0BMQUueSoE/O7vJPyrC8CGMZXOfm70vIinfGVSmuIhJTfyv4NTzdEE1bmzuJPPV
wEwElfb1gJuyOdMM+iuDCQan24Av4vcvnOEQ26f2IwH9BpTSCSFRPffqDghMeO2w
bPnZM68443lF2hs4sV+m2ExiW9OmsDt8MtNA8hc7MBk9QYUafxjW+jzPhdHsmEWH
GHEu4YspY0l1It/v5FkvrCe3mkYUInw8susOmlx2lslpTUEJ2pFSfxZiDZhWWqrM
yi6R8bjl6TSVA96dSXUNttmyWR7ay7EaBKA+jujvfZb+2c0baGbg9HXUkp5TaZyI
V/3GZljabj2hj/L6jGUmypBxcga4dDvXv3xM2phIo8izv27L4GZ+hzAiGD3Paxti
VkKzRNGMf+fW53lHxUEpnRXNO3qovx4UpF7+qOfHqIHIUzbfjjOtG+jU0H6SEgD9
tWIQtDsC8FOkmN6Hft+tIhgjDH09lvCSgm4nAL75KLDSGmBH0H+0qw8jWtQePY9A
sNADYGgeadxt8hcL2QcFy8SyqqLFvukhVa7MgrM7J8O8SoaqSLn8kBY1KLjN9Wok
h/8O/6LrHxHIrRY+SnOk3hG4souBQyujleH99clyEwX6ngnKFuKTlkSCprKY6MVd
VtX8PMdiex2oqAiS12mdmryUxE7T2qZzTt5zm07wEZ5W7EjE2RQxBy2CeISXmQvk
mLYYGLThleh1bIM1vZfwS9AIym5/uQ8SWxpgS8Y0tGIl7mpi7ck0xckqrXv9sg4e
HmCfZZHnQoVCPzwWNVk5it13Bc11ZVr3Ny+x3TL3aI7kafG53JGVXVNuI42PdOZi
Fsw9pga6noEoPjmKHs6B6SR2TzxmrkljkTAmIW2XKDEj1QlflGV+AfJMhfEtTW3H
dZrVElB4UX1FNSpIlr7q3iNiV8OFhrs8BZTJFwPdkLnXC+DSpLXUfnE5S8Ogzaj8
LRREJCeiOtegPQgT2DuJnl7tB08JvaXtmdwHm0vTBYXOQo8q1Jajgd2VBwjardsw
Ftt1uil9xDlD0S5cRs8V7zL2YUVWr0vt4rpfS2ckM2ZDGqtbHR6MZ2yayzygFvow
Gw0lg28H9lAQX30yaCkoS3b50Q8jlMQGb6NO7qRCKjtuvV4l/oRUDz7jtT9/uJQX
b/9Znaxw5AZs29PqPa/gWLdz8iF93mrj9ETYA0c2i0vefnTEAcx1kmP5yAqiEdhR
vSA/BhvlD6y4Ee0+uc5XxxvT3YQUbhNLTEdAB+EjGkVN4hmRyy6KL+SnHKE2b4vI
rof/ToG3DMCiTkl5piaiAsUaAYOiOlvutDCQJIilGjzmGijKoBUUVh2yxixyvM93
Wdl2r5jTxYjvmHOwugLzv2OlvIVQsyEbALnDKHDQfbvswUTrUJ9EKVV7yFx2HeAO
hIyfGvKbYt7WqptWN/pQiirfDA07umDXRuQCrKGKbtpeU10JsfwYEofBubxGKt/A
0ziojutaf09cU9xZ2HzNgHQoMyzH4H/wU5BaH4cAG4UQgxycvA8m+2sFZCZpcvn6
L03kuiZ66IciqcoJsiAtEvadx84Oyit0tHUC+HQ/K0vAIVF82hEv19qd0mIePmin
AbYPnvt7gWhMe0fTxC1BaZqxh24CzToOzfvMNzYVxhoeFHYb7VH+7C1N839pNR4G
2wd0gEinRd3VtOpl4w/z41opVLfXCzBMzNXkROex8WCS8G4Sxme0sM9KGmZ3EzJN
l/UWd0FpoFKTwFRcaDUdu81w2E+PV9R7ZJC4Y4jhbgcxvh67Jdcq4PJJHu1NgtJx
65TJWi+94PWfSIFDGhl6Un/moMm1uzFmAS/SDnyZDTd+X/EyRMDzxndps5lDmEL1
Rqx5eYK+xXGeKLXbrYYWJe930+3+Aqc21937MqcorJWDZWG1gNglENGR/u5q168D
z8VQKiOQm23eGFHkswzup5Shp30ZT2EKeMVwKP8da5MOI93IvIY2ZbkxEPfmFGs3
HyQ1NUkra3s1rHuPWN5CyGTEF1oqXJCEk9i2iQCbrwgzek99dW5FRLJquK85x9va
OngSJf982mguCSSHmlWc+nQt0I79OS0d1xWHA15HS68rH0bVoCZeJk/KhQkjSDUK
AFvZK0gJWSPNaQaSQchrxdDaebVxUPNHykY1Fi1s0CLX5ALKWU+2F1+/l7PejcHJ
ZVLm/dUCv+VVM/MrHgG6d2enkzYgE3J7NVldaGyN7ooCfj/uVL4dP5yFwy4+MhZf
/756d2mPGHIehBq0/uEhsYYL7Sj5dx135csnrY+aWXXyDGZiVvaZCd++jsbUUxQI
H3pKk/n4RqcVHspJmW3WysUzJu+rHYSWxH3mxD1GGDp1NZ/gDJ/qycSVVpYE2KRK
3z4+Ff+GMog9aZP3oeHv0bjI/pZtnGEWv1ROhhqeleUsXiFM/fylV/OV8bZteKyh
hwnmpwFAkOvhIOonoQ13dxGORi2vAuGe2spmLkR6decZiF/a7TAILOo0j5kkC40G
/ckCs98lUP6OroA4sHB2A3xQJADXmSK69le6wY1sj7S/1uJkFIiZQj5NaJT3I5fU
cQB7R2AZMhVAwIYwyvVhuDXmPQEMt4qa3RaswrhlIHQKgRWUYuQ4TMag/3pWK30P
ZKaxf+nTshybhJqaK3dF7XPJK2VT30KSpkmTs7FBaMCn9uWscEoOTM3gJ2DIrXv1
BaHJoNiKfehFcADsQV3qMGs6GYxjci261IBi4SgO3j9ug5uNi11oH6TRYZ/SX7dc
+RqHLfUwr+/x5cAAe8B2tPlhP9jSHrmDTK12yNMFJz/r3hpmki8l129IRfbSj3Us
9R23cDlbSaolE9ceG/hgqd6iM7wmrJJe9PDdG2RMbr2Yv8rUJKmzhSCVz7LX3L+R
bsBP+i99zueF5DOLzENhXoIiyJJ/bUXvvvf9jEEsR+A=
`protect END_PROTECTED
