`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RdMPgrPD3/lDtVp9ECc67L5bw8GHCh2T+eFja362EvrnJL5L5hMaNHAXWdZSGVU
D5Q0NA8vZE8kzBxMZxNY4u1T5CcmdeaSo+gIe1qrTXh7uISyPkM/9fmuamvRnpdu
yTxFMAWSsIYCS5yQYTD334M6Hvafva2YNK4sgxsBqknYLJlBqil7Zdk1ST0bJP8g
i6w9IP7CJ1Ez7mqO6paK9P0UWYLdi9UJGN0MfYBnxKtCdtOZbh4U9H80Z/+Mp5JT
HgVYeVVVaNgh3lsO1O3jtvwjiLb+O77EpZpf/23A6pUJwhR2cjhGgpyRapC77gfQ
Dqll7CGvJmzh1qu71RbOpRzTfC7SsgzUDirkbkxaldzQdEcYS3Jfjq10MAFdISuh
xtWtt1y6Dcd3fkwruQfNg/QHp1YkmjT40LeHPu85L8OXgUrFCF1X8KLsGH30M+2S
0qPEIEXBvMI1mVf6X1/KG4CBUnkHomiMbOcDZFq6jynOIeXCA+voQ/C2lIaySHu2
gvXP23CGykgh8JUc60m4E4Fe7frSMN4WUZ0IIkjHYkQfxzcSPm/CIPsj5u3vW3C8
5wX5TNXGDDXcFxTvFsX7DVjQK5vdvxFkIOtF6NcE0VWLYfATF6smZRCA8SJ7j1/j
xrLFRneFIQKDloDWEfTN4ayXXm6bKvv5Iac4ydSi9Qk=
`protect END_PROTECTED
