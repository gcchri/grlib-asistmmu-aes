`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2df7KPKP/+Bxt8Bh8tKyB10vXv7tJOlELBJX03nkijWvrW+1OG9it/Z/vBvHdKp+
jv6QSiwxsixwTZqraef3is5aphs3NDQLVUjbKobwvdivsIaUWuPc5K9hS5TLpqHs
Y+0hXEZVgbq4Ws9AhcqfJy6zk4PdEz6tdB7eNKnRSrP4uLnhTGOZT2zLsqR2rTqU
ky5sU862wXWWVgiy9soE8FSQ6KCgxM6YDJE15n2RtJwa0J1R5CZX2xsVS2rLCePH
rOkiMtVnq1mxga/OSccW4PdteeuY4TvYMP3XDKBbZTani0DVGy64SIit+5ihXLbu
vjbaXf9oLe/rY1gWPODb3s4AEzDFBDrIKEQ86B8w07YTur2nksONjxmXiGP1sK6k
WsE78Rkxp8TE52aSrbUrOcfIyeqs6dJGt/7EaPT6MM2QVm3Zv4G7SLpVyK5Mo8GQ
2ISXmOhpEw/GuXArALG/KZDE0esww/j6VghMV+yFVS4ZwTmaDfkYN5lTLPn7xzmr
sUKO+bpcshRTcTn2Xksi40VxNQX7ZYoRj4/MYsR2syS83lvW3Gow+i+0xi00dYD9
BoqtmViqecGGM6Y7ius/3qPeusxeT91t8BOUjQ4RvrIsdPIwjY+A2RqNfMP3ofUy
cnpS7By4edQ/iEWF8Ice//HaXY0RMGRN+T2RjeUjIK+U6H6fWJGm3yuKuFNarsxl
D5NnIRuE8WdBscYaR0sJZTvsdA4B5QIDo7PxCglYuUanLHDG/P87rMoPitYud1VI
+R5NzQ8U4zuVspMydAioyVGPj/xYXWqkp3g6oTqYsr/4ZiTAT02JzW0f6wZMHxKA
mfLtt+JyNkkbMoXCkvi598hKHO8kACLV69ATJRzfqkrWcG79DoyUAk5V2blOW3CE
99Bj4rKzfI6CwOBvacBwGFHr7WxMrTLBqaKGBbE25WjKp6O8mWfya/bovW76xDYb
GAeRp6T8yFvFXRrBax5mrXTpSgEYz7qGkXE1YNZ4gcxiidS/CQnuSX91mkndAzbi
Y/vtcMA76A4IYEG+11R+oiM7/5ljZSn6trpd6O6gPbwZ4ZBg37kJ1O6rsJxBBJn3
JiFOJiIEBlBfeQc+8CnjH61ftH2oLSaxuuuPC1XH4oxod4YFbELSG5PW6L2n1eco
naS6xLV5otO8CwD2iuBxdF80Qjf749o6RsIXUYY0Ye/QsuyaNccCtlYtoczVetBk
bD1iog6YminPHdPBjAqJObNzeOfv4445BbP6xONAQFh6vJA7hsaRWHCZnu4ObP48
44Ryr+vbLhvDjHKKwvfHV5KubLd6lTJN8BQoQ1YCfIo2PNtqXkstP228LQ/7XNcK
RSQztuQ4HdnopEGpsu8Qk09Qo3hNB5PDuGuomXj95myCgbK3KyhjNYwF0ezgnaS0
zXdbqK+c4BTEUC7zO2MnF0ehfWFLe1JfYdeL4bJcTQJh+sdLCX6GHRhC8pHn8MTK
IzAOqrv+6/KkJNpvNhWP/VXsMUfwUFnMZfG5JV8ehJvjLXFLIkAYEJ/dY4bblrbB
aJRKCYyI/RHUMmbTZtzB8ZlGAU+tILcG9eXyu+Yth1S6timTNB8SIqmhr0XVN+0X
1DZDVVKPeUlj9Yd0Z8rrk2SNP4XDwnn8FRrWCKsaGCIIQP07rSxvSsB9S12anYKj
YCdXXXhAKIkk+p5i+bxVQdCQaKAZ1yCSiZ9DLHim3UtAbrrtDaQLbKxhKp9d3EmU
tf6ZdcALbWFTBfqp1w6CTvpVfAcWaX7UUoodrcXxa7vOhST2gZXSf+ylmAJRNKaU
T+bKSrdOFWbd3BmV9asXXOYXe+CYcvcAZY9S4W3zb5sa6NYz8uzBwwzSEDUTMygU
BWWYczLDPLF3d/7XECCYkgUHkgaLiIpzsM8a1dpj05sK6HBBNVLER5t9vxARLrCh
gkyJWX35q5Sgj0Cpzd5eYxOFsJcaYnfv0V1RFtsKOHI=
`protect END_PROTECTED
