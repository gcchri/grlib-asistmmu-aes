`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVUHIkl2jczOgSAPcTzcNEYkIJxpR7BN12FooIGbluCFQ1cpI2embyZHdyyv6ywt
i1KhsLM2YuwfyxDBtaWfJ/fzkLZqXZ2Pocf0R0NlIbx77UKD4HXpr4WTwTZoD5On
Oc/rq/JLXis+DOop6/W/vAuEyU+ptVu3nwHYJz4lKC3v2sHLPNvEqHSuL3qIVD/B
xSWL1fMXnwVXaDg54rFJStBsz9mXldt8d5lTzlajAzZnZ/u8wCcmswg8mz3C69yI
SnTVvKrCddoJeX+3axAsxS+gVgHbIHFbm8VfJdT5bbuO+IWmImtiVzoIXjcaUB7x
vw7ywdVC2K7ucVTbWOnU2qjDZOmzXiJaFVsRR4oKKSlf2ZzrDLr5gc7Yh7ZYorhV
Jt76Gnez/1PPRq7Sn95hx6klcDOkjrqA6uFzEssMj7zOCqJ48T9n8kU+M8X/rk62
ok6PJICBORLUTDivN0TC0b9dIppBwNjmuEqdywBPfaDC34LPuHj5mBaVgCkJZ2uR
D4cDTX2ePEHL8baGrSoLhOb9w9kGIzaZW+ufJJagO8BdZJUOZ+Nsp6B4nZ+9gS5A
K/fuUQx5isga9qXjJO/LJ4X/dHv0D4WuKqTD719APBRjjY8GOZXvYst/66gWZ+/A
IAeKBpXHIC3kdavFCxLdLzFIrGvnBxZxuUUpAt5fpSCUjGc2w1RTq43rL2pj3lpA
PMJ59b5XnhB5TDqr3MCc7cWzbLrhUTB5SM840AQqLWVQ84vLHanH58NZhzzyGn94
oSBkGxqODmo4Q6if0iVz4Zj/AoL+Qke/tHEHoIjmHU4vAfo1MU3Ckfdl1Te85pX6
nn25YQuiAeB3D1p5sAiObGg6SA+LkoU0Oc8SHVra7/t8ZbRDQjYrnvRwsAcXd2od
/aMRXFeo4eCM0qZzeQHOYGLRRng28j3FUu50508ZysuUAtq6rEADHGbKQUJrljM8
N3ztFaS1uZvzdX42U8SRYVh9iTyNzHmD7zWadDs8BIRJ3NKF4ZeHWNxPq7FemI7S
kUKpvWlMacrtvKkANOQtg9DOYocOZTaNpbZ/rVt3rHr/gqORNwRK1ljxLWiXPy72
HQKhq0M9sXg40YwwulLzWInyTdUqs6619Oj5Fu/tWRh5H9XJ0FPehy+YslmQt44v
APWDSKdOnbzc9ZvFR8i/6zL3PaU4dtYfRHSYbtgf6flI4622qoGaag+/RjUwhIE7
TqSLeFLdOKIaKECCecuDHfO7Z+/PBh5rRJtVdIj/3RqbVxItWYC9Ge/qy/ltgVSq
`protect END_PROTECTED
