`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SDhrqkpVVyT2eRfYhncWiRPOzMex/n/uJXCVwqIpany7ct7bVVaR/Z9eWmEsbwFw
DaN+WZW4si6fIFmaoN8rr7yvUpBTtgZdDrBD2mDR/EhjXH+jW7dLqOrR//iBnW6I
6vu2ZzlYzm/N9/ak3rtAido/LNG+ExfEn4CutrOIhndkLF8YnI4RlXgaGWTlHZ/9
0WZboYPI6DEG8XI7hbnzB5Jy14oLKFyraf+NTOjqxkuDqBs87lWfYR1wFypGJOK0
xTcBU1Zi3hoVfIXTJDrvh+v7usE3ZF1dziewR/MMQLZGanRdk+pvNvGcjAXLFS2k
Pf/fPKUg1SzJ+UZWAlnndcMpun7/kG+751vcsfZhS3IOGn0TM5SlrzYEvTVZd1tL
+KNjCckm6NcG/9up7wVo7zZL0Xv3czG+GiQw8WiTiQf8igeq2gw4BhiHUjQ3zIEC
`protect END_PROTECTED
