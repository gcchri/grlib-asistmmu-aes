`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+yR0Bwy2xmsrwFsIsafkOLCx+tpWx9hKL3GcFtF88S0UfVmDXh+FX1sXSE86OqH
Nrqe5i7o8aLzoWNfi7OYqIOwwGaGr8POeY96Nyp9d19yr5ZVmCV2iIBNFNd/k9VO
RAFMQtc2gQkCg7pQK6qPdwmGGlScPnznMe8ocVWcdGN7YC7ImwASIscBu8jSaA9s
PW7miFxnkwUG8PhkvDgSGz49Bj0nkAbzgU7ajvoN8j0eSsWsE0ifhGkSwkDi8oOI
xYl2OWLwAVMI9XMS8ysANH8KqqUgfIxvrQBo4MYqTI2XPj1mE8Aqhll0ajKcEWzC
`protect END_PROTECTED
