`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oWmojzj4D0KPgvRHZq6iI1B24u0lz1wCYj+29MT/u3PX1KqXWfzCroaIGMPFkoV7
djLB19cjsm3pVVddktyRjwzweEix/JLX1luCItvepQNwWZTZfnNokZCwkNUayNh4
/Eq2Qc1EAQNXESfGtqL2TMtYz1Djy/DY/7cO6RPTovHq+/pO0NaOuvRVExty2VDv
Xp2wxgIaE4Q09GFPbHhO45xF0HaYuApeHyMoPIKMsFkdtAcAxSrzDUEQgYwCSTRb
tAXEt7Y3JGcLhaOJpI9ch89ifA3CB0JPel5a7l52UuKMGgLYVzLBAg2dvv3P+MCB
H0TnTDZ1WYCjhbe/5G4ZPjOcD/ke/Edb4V9PZ76/+JLfy0UEioEATR+kU5B+3hHh
ezb6X2MqUafu46zA500/MzoK3Iv3JpKb11nc110T6rCP6NO4usJ8wi96eR3TD7tj
9DaWNbtFnX/3/55cxB7QL+RzlU8FGNDpkIsC4W99nChnrcjmyE6smY6lVjtz4RZy
uzuYfonoOq7k7H2A4qIjcjqol5sK4uwwyNp8U07cgKAg4EQ6gk1neFEgB5EXnvFj
aNhTgEu1dlnA8AhQQXU7WlLaG5kYkT2AsHP5ljV+AzVoXQ4O96yHSv/V92wZNC+q
Bpop7J8IAv1ZFNvKSEeB7i2WLEWXaVD7WxR6atWLMlLh9KUig/aXtDErzuBTSXCu
GUnbu9UHAOyso5bvdDb+f+IwBRqc4yV2AX5fvDQ7pK6cnAFoPrZreB1bke8iW8YE
H58s6t6ezpbK1t/15r1a7w==
`protect END_PROTECTED
