`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0atn6pIIaizUr/VJLD/l2s3k9XszOFZmi/mDjmAxLsefQW//3HxXizJCzjawI9P
NPJkXGphnAxnSWlMAttdHABmiUqxhlMhBLyIMLSfJmUJD8kackrRxzs2DGa39260
0xfzV6GmP2qEezz2ZjjEXA+oIsaFszQIJxgghAMVj1gOlvLytuVySYzVPKxfnT8/
QPbM5auR9gSFoTYHNY6VNtGhWXFqtAIBJCRBqBd6q4OY91SftsJToZgsmFAmvmAF
WobFnJpPmfW3jR8N9YB/L9euwUhHwJnrhK73JIFCAYL8DqlapPY6qp2UMfdd98fU
ai6qrB0TF3XS8QXYPtOnEGi3rxwCeYp/7iorftISeWEBXgD7+43gYeHbml4Zf8g4
6NdO0p4VqNVBMn5gh3RTOWX32+JGmM2XbVYDWDSVR+w=
`protect END_PROTECTED
