`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
crjjXsf1urUE6BFIx93iX3Rlr7h2qbe/OXxPVx0a9PWurlAk1VnqDPtgyh6LrMXs
cUmOHgldm20E4AyMZroHoXN2yw27nxJCxuobZtmC8wSS8lukJdFJbM4uUrMkYNfZ
8vLHcd/Qi9k9PkOpeN0xIhoAAx3y9CTc/lVS7MouIyVgOpN6Aqfloh3aix5ntRbU
oQly1QwPgCivnH0P0QloaohhoNHm2lrkQaNLBYQnyzEagPg9o4VN6yJRU0bRsJ/h
7r4YmkHCFz1ex1y0EGJHejD9IYIscg75/lNsFtpcJ+caU32OhZ1Eeu8gdj9AkK7l
/VNTrvd5auhsRqv3dCrdlL6tASTJoV9tCqiAwv42FLw8TENBnrFH1N0NIHuQWrpm
bR6kXlfwvui9IChpLltuNLhqhbj0DzvfYdaA9QfP6zI=
`protect END_PROTECTED
