`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6cDAmvpJbL8Y1XTpZ6x5Ik3Z5NoUL+AWF3BdqUkPl4zTsa/roWvHYc2DgrZEcVdM
xkF7ACQ90wjQSahIEm+dn850GdM100KBpPwiFQKSOCBAcb9XZp3ksvHsebxxIyBp
MIgPspPnvNrOK5c3ztag8W6q2LN/KYqQ6tn+nKf/04v0TrUt7O18vXwpclZ97ROH
x9z8NS6bRsYUFi7DfIHbMy0u7wBwToXhr9tVFLiwgGd4xghBG3XtB80/gXcqN9Ds
CXcnz1g4PVxZtusm20LtT44W7iUHaQG5UCWpjTFUpuk3gCN7oKXlve4uhuyFM4AJ
N5J425TqQV1eATMBKsUC+CLnlEW4UARe8/4Rz8XSxRtVDrQnE/rBkgPwPoT8YT64
nCZPICMytscV0XofFQOZfX2CaQVX4IFSqRUxrxbMC6jR0gjJIUaUDnpTDZS1W3yW
a1YZK+Jmk2NH59CTTSPhzeTuJuTQ0Di2FQ2kpYTfxwDAMq6o6X17O4t9R3+Yy/7f
gTveW17eSU5jDZEeTIagESKjv6fH5UrtCFGQd5aBc9tk0nscfc7N5ySA+hK8ZPFK
zUMi2+j3J6fIDsqU/1QhCZWJ5BEJSoAPjtXHT9VQdoDl3Be9lPUEaBsPXncMwO2z
egijhpYFqFyUI/yo/2n93HbIdaq0POiShaHpQdSZOId/rZNCapZLgYwnPIgRbFz6
5M1p4NtImdb1X7SBRy0xRUJIt/57ATrGLkKkBGUoZ495WIa+8PObY1wbXgQ6Xxzp
jLQVg4yEejTLQ4tq2G6j1MDBNcCPfp/Je5GgNl8XEVvkEYZzU8IE73XtQLl1eAop
wwQrypW8up/Q9atT4WMBsiOQ1bhOMgkI3GciDeXhI908qnGCSaXCqwTB83sjoi2x
x5iwxz47o+rQh/sKhtvoQTevIj9H+npmv4O+XPkoOviGZ5sINDdegz5PZaDSQ3lD
CEcFWtnItmu85wUYxZxm6AuPdbsvZXUXmrZaJSwkOecNE97Oz2tT1k69Yi99lVM9
KijS7kQtl5MY9W+BPd89rw==
`protect END_PROTECTED
