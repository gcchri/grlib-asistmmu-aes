`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i7zAOCAq4qAIvtXy9jCW0Bssw/OPJI39nFobRkzZvh2Dcm9GWI0FeRCAI5paPBdn
9Q9DwM6tW+sdzCtwNtqkIDdV8PWqAE295gf6AMtgf0FNA/LnNCfdJI8+f6X8GO0m
P8RKWHo7DYxFrypg3G3F5ftLQte2CSyftmALPa/So8uQJyKZtWSkoLkS2rX4XEg6
in0wZVj9Twh9hDpSm7eQ5JG4zXWWdmln/NlqYznJf1nhA1CF8zOgODKKX3JMgVHI
FkKSPYaC+8oMLv8CkIVFtWxEaQQieeV5t81DFqYrX7zjbGK7W4zE3mVSNksy8y4Z
YErMi2CP6bQliYXdgEhvZYOBTC5BGtMXqkp9BedNTOomqwftHVuCs15KrjLAS8PW
lPK70JbdXclR5sAd7z01pWdUdrRtfaJXFwA11EwGajgDZz++ZWzrGJ3hFsJDc5X2
VBkxw8tapANPz0okxQEQKcemykiHXJYbXkMuqEtCJh5wg4uh0BoVBs5kcyA75bN/
2VNCLZQMnaolvcjhtH8nNynoktRhErI5TjxBL6unRvSUymCTA2nimWEpn+964rWR
XqkvCSC67BJ9VDQZdgIMHIt5lZk3BddPbwxyCcJF4xffd0/yTmGrSqIWEb0AlD4e
SwOSLGYhpgBGT9leq29TN21G3b4E6EwMwp7VKLMtN1hawu0PcRBc/tnZ+S6Zc43m
/tcQktdXendyQmUXfGogBLkvFMg2pa11ZmZ+xMVstrcIg2WJk94nsA5epywXSyA+
DBTKq+mzUzJMnMiPacHPWdq0fXvdT4xS8UWmVlf4bt85crdqC7Zq6q2UKe/CwTRr
GV4SFUsugmXjucSBZJfAk4g019TM+09IU4y49LF1h6f3rS7QVT0vKqD82n4Q9/JV
`protect END_PROTECTED
