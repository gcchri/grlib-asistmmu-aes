`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBfbJKrYuWxS0XjbfLiwiRcvxQPnaERT2pBl/NbozJ0uacvbpnmGhsPgCnGjnKv+
DGiD1xvLpQpeBSXv3kowNRY/hTNrn+kh4G10QOQ6nhs8/NoXbgpXtloBjzFGEbsY
LOIPydLVrVYjwyd9Kfa2hZDEF7JPHRsX6SyDvGnd3fJrIC9njxRMNynBde9RillK
G4+xaOjZ1IZeZAWv8Ruet0kRitUvY+rWpHrBfP74DmE3gcKd0Z8muVbNXxWf+YFk
Lyf6NTfg8VbJn1rJMJNPYisLehI+5zNHivxfIN+Lqr0yDSvSjgnDtHbzPlSVjvuN
ZImQH3KHN7JpLO/w1ikSo3vpOhaJZ5fvSCCqAlJmCTb735gcWtpnjHESBVskchyJ
`protect END_PROTECTED
