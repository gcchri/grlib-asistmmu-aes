`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
msoTL5XF3BzgEWLdpveXO1gk4WtZex5Lc8wymFRUXVRuWJWbAZ4yg5xrZPdOsXC8
YIz2ItaunR5Q20+2duQ+jeyJyYdoHxVAw71eu9f1e1yJ3T1EHmZJumC4msL1HHy7
i3XxPkDLBz0j46ajcSMP6ZZ+3hxWd0pImm/VoN8an6nAkBsdLejytlsbrqEirPx8
yVVlVdMA8GxrnpvpxlDkAYsZeeW8pUte3J9UtLNN/nrfMCwr6hv2seO98j1ODSSB
EL/RFccwnyEeOYv6NiWOaRB1qvLqcPdQLp6XyphuNnb3MNRBEOtHJml2a1ie5fW8
`protect END_PROTECTED
