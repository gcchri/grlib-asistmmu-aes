`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ttJTRpTU4tvxNDXI68xGrrVI5NNyfikaGb5gls/0S7sD0U6rN+l/HRRzSvkOvcUd
Bm3gWx2XdnCKt76+KZggaI85SCQG8AIlUluUaARCA6Fz109YtN6n5tMUpuE+vCbR
mpzW78y3YDSFkPjclWK1eolo7zlO5T4gDx2oHA9igBegUmvrhpds40TYwV6q/sWG
Eu4Ds/Tz8jKAb5hHKUP/wdSDz+CfFSpCqErL9WTlcM0VTSgYU9t2hNvH8qgwKYe2
Xg96FAhJhCq6+iYLVX3h7roSYj0v60P6un6GAZLFtojSsekSuP9GKih+pBIc+gCB
`protect END_PROTECTED
