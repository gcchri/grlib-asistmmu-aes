`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7EtBxjCkrJlKOlvktfqSwYYiUTBhlpuh07SqCAoQE3IEJZGdJxdoA0wnKWwZ+TC0
8pui00bMvcVdM0HS9Uu1a7EB/OUS+9kuub1T2oMSf/09f3zf/AfPlJdTwVl7gVWu
7XuHqxMtrN2BGzj7kAJvctPYE7bYOfmtzye48ujJpuMzJfMhnsNIrrmOmizJX6In
j6dhndNHM9ueX25kBGmAXaRRE1+XCAokyPdYXqt7phmgrJfSGUJfSmO2olPRElQo
+76k7yw/hLclQ4f07RB7KKMy6Q2uM6dLnlxSW3D9RQxt4BBvfNBej3TMoDJpy5U/
kM2/C8ShNn8JtybcxRIoMjcsCg6nezMPXJUYm4BCFe+rzrUOxXOj04r/WcLv9Jsb
Z8V4IhFd1r3qCxexO7eBzTDxIGK6xDcyqsR+Njgs7W380ZkYL25a7/qMEr9tsIQ6
b8QClANGZWaxcIo+2XnSwh+TKp6jnWQj7dzOpXPQ8iuTDRKsGR7bzqxkktoDRu52
8Z3nlZ3zAM8QHYutOZsd9izWkvnevZ9lEVXPqvWqebwddUvWARSyNGFtA3wF2jIy
TWGQXUoX1QHada4Ep7lG82kV9LscgUgPx39sfOzFQfV2nn3baa+W2/AhO6Ut1WPA
z0BqxmgbxAcipJQJwCOmCd+wONxy0rkBq9hGLvzGk3oG8CyTgWaksqut8/zfrOkF
nVwSt3Y93kZC9sBi1LoazFNqNBm/5jWV6MxYGVtmwS3sV0RekVQ6leye0S3phUxk
n5+4PLLGlJhaou8K8pg6xuSu6q8uCmqjQX9Er2vVmx0tY8npdgL0ESp5bv4pb3fI
o2jndqDZHl/Sgg/ZXASCYrkjTJvVoZtddugujq3crHunmL+2VBo2r/SxALwoK1Cd
D2BWh5g9t1cQ5xrp5QhPtnxcpCEiDaJww5PH04OzomLcQrNi9YgpT/mfn2614WVf
lNOj73oBNxiMd5aPTXUwRpgdX8Y/nIqIXQzIDU5mDpkfTdDZXCsq8mkDsTkfebP6
7l1HSygYzjYBCJXlZ3E0kBUtbp+guxESwNryoHXb2hhJ9f9C94rA76cJjfu89otl
AXjuNxIuCAV3tSbq578bQda+nOKEmI6R8ncrTSgfDkyCfrFk63gKbhZEtA4xEyoV
FFo27nQTUVoCw+xhIYVrWsVxFuGjNsQxWH8Z0nUDtUqYYjmUNtaBl/Yb4s+LpvWO
mIxU3QIAR+f+GTdk7gvwWoanJrvFBSNfFmqpn/9d3bH+vIwchKaSIt4RXyIa/Dw+
HiIbUYiCW1FZL8Qmn71Lk/giHhUhseDSg4YcxSrnh3z3njyFI3DG37jt86j3EW0T
jnMfAl+IpYJjr68Da3mc8SGMOfv+O994XSLY7/vYIRBwU6SgmhRH05WO3/k3IiF5
aNvnyJ7mToY9dO2IPXn4zlLdFx/u4CtRUW4kDr0+w3JnKUi9fbQKKAI7DG3IrLC+
2pEO9YeyoRYSvAAu7FFJeCKzxKnIMUO4XfxWYOb4RrOyGi0ChkzS8Psdt+Y/bQbm
`protect END_PROTECTED
