`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BoQLgvAWlhLR7zKNBEd22IazD9ka4kAuocvMGCKlYpdL13DMbMPNNSF0Ib+N03jy
8pHBleuQUUHLFH6jP0me0JtS3SxO6Ersi6WLVemrgN39NNH3f9ycamPbmGjk00cQ
x3JUnP5o27ihHJ6ZyOaWyMAO+S//0FSuQntuo/c6r7wy15HBjOcbta9+fY+ZOWEB
0YqqTVhE62dBuKZMPCm5gvIw9sjgHPO3RAtYrRCB8AEwp3SeyyQSB2KM3xHPOOyD
FvjsCKPToFlGavjFK3R1R6MSkMzyae4lJPQpU2YpDZAlPtQrjDLE/3Qn7xwIlEzj
IGPJq7/S/J7qFITUP9ew7bKitFau3lQz7eBQehJDPS8hLrl5bgtJqiQ6uNzuxBrs
jUZ/HOrKc0nseDp+Ou9EB/ub3Wkz8AuQGFgxVzCf/70U10q1dDjOa8QtEVY7h/h/
kbiH/BMDl/DpOOVlmg+PSSzlXHCImtWmc0E93uVZQBD3ew0o2cJuBzD7P2TdlPsX
ucuy0b+f36Uu/p8m+THpwyE6CN7CxjNBPfVM1BIYaFS647EtMv60LUhoZgdjYPFp
e3EJ663Cto1pzeYOKDmXAYbCFShOltWlD5pjXpfAeO4uAoUHmOgPS5x2nkJnEoup
60nBbUYFE8f+zbl3iSfCulXshwuyXBn+ncADXOBnpqFtd/Xgn5pEN4fFaS2F5u7e
uAjSeMS8sxk1ELavwBjDxCkC3sFbzW4M/VW2SIe6WtPaHJLTZhtBJD04CFpMAW3M
/V4bF8rCTLY6gqbA0lXPO6yzKom3q2ZRMYAO6ESHQ7zY7FauCq/gSfpNCJYNbru9
CVUYCzGD7ARqb7KHTolOdHwR1E8RgSPXqLRXCto6beVtSYB90U4PeDQ+c2QpLVsH
s+yZTk1h1npVwjrNxyCdsrp4GZq81DKkZRpwlv6jeU+tksYD/5QpSp1Qu0YXw12f
C5hWsDrGRHoF99HTU8BycL3jpbfMQfgtpe+R8aMN4m0EXJuKZ2hMAZFKNiGv/dNQ
WYj3i4+1LwfEngUiEsDbWKLosNwRtaSrqTqwk5/5YopFi+KzbKqaGCcrkT7DNABY
K2Etw6+EBTy2bI7iCgl81MOIgdoyH8VGQ0u+YpZ/qBbEc5sImiThzIQ3GrsvlrTw
fqMfODAGKzei5ciV+ImMc4TvqkJ4q+FrsibspDefJK0/NUsUuD29mI7IE4UfTHk4
N3hpyEDQbv8uJl0C6UK8/uCBBo6eYHev7C4/uCz+ewRLAV5+jeU4GejtepDg8QpW
57glHrX5zRO8URKvfJYTjPW3yB7oh0UrQLn7P1tP4oUA966hG9wgy77PjyDof2dp
Glm/ASOyo4NvUDOFLz9Tth6BkHNlyjYwHuqkWIZFtgENKYXeCWr4DGPx2Y9Pf72P
GsMuraFIonZDQDQCZfI7S4JDHJhL3U59k4LtHJREHXEmn0TH/jYUkxEHaXW8LhcV
CJG+7WKlG/8AeMk981iZ+xtCZTXTTOE8PL+KI8m4qxU02m1d/2WHeb5EFhBnrUf4
t9W3H189I1GiQz8+1FVrR5fTwrqbg1zArbpfTA6Nsbx3ZwoC86hxhDjOp1SU39Te
NdCh55LuuyO8Iz3pSqwzEQouN8+L2h+YFTygVd96O1XEQP64K4OjXp8ANhEZORdT
jjMAU90u1bBQyIm4Qj1utZQoGKoN1I0XnuzJNiPhP2ueM5deVKytAfDVLWQpgYCC
c/KVGrPi1eSanvjhCuqs5ljaFwSTh3jq1DleOOy1WeRNQQCLWBv2toIaoDcox3Up
MEoU/LHNctHzkuwqKBtcIo3AZEmZBBonLwcN/iW6Rq/z3HFeEbvdCPGWw+O859nH
ndsvADbILpTxgHe1QQz6OElmFJYfpVZleEyAQsD0ZpVxcdebt3EfThT0ElWngVbP
eTy85C552ekzy/g/oSDpYtTVqXNYj3NW21tyjHLcO9zRe4S0ISh2RQGLIB+OXR59
IJ3YQU8WaN+7VXIKReUurt3PWbZd6jdSurBAk8v+794pHGd3bQzUhxC+L8VowQzD
4vEioH3WIrfbTLhs1ZSgU59Mxzfsd86DJRPszu9E+NL7Mnqs+JJxOOAniHRPk4ic
WY4eKehWAZTD7goBvAIB+/z5wU2fJe4VxStIMUCr8eH0gUv8wMI+czf+rwNzyiHh
ltyWV/dPHpJ5mJw6hmQnm0GzExWx2Jjc8fuWIX90afy+ey0AlIQNri/D7BjaQlPb
tRfNXEY8HhGuHQDFe1SRcz+if2Ih8wkhNuVy7072Lq3NuAX5R48RJai6dE6xLYtx
oEvXPY5qabeXxj2HDeR0wVh+ZSraEv0yQF8VbjvJGA86Z2ReU/w93Y6NhpuDnS2c
7hNqBhdpvJJPWY+ilBFpSOJAeiwJUVx/Xvmp1+dWZ26PR+G06lgdgOrN1kCtdUec
ruvNvK9EdD8kR4eoFYgnO2OOrT6Nlebyibzt2ZnnMdOfa0KjupnRMsDLUBdQxxbe
7pqs4NrSDWoYv63n6V9SvnZImyDqbxF5xMhqoKyDlcG5u/gbAqcCHJm9rEzxy9Ef
Y5u39WBs7sHzh/i24KPCX88s5rHdIk3DXu/+LviNDwh/6d8Sqo/p3XIw8B0/zc8E
FezYq4eiQhe7ziVXakM4nfryL61LLsK6h9st7wfMlpTtYyOUC6TSfigN/xehKiOx
2TbLcmjzy8yUCoYnzVUAnfQqaW6G4H6Rj6X0h0pO+veQwFbgoMmD6tc+8Y5U+WJz
+wKigAqSKsHDB/0gWUWWcmzrdYHW+09JDz/WQd6+02xQLllKtg03MXhefluPengU
fNSpn6vu1ThK3cHcruwwYmqFyUbnK41/fKemINZE4pb/AZTKDPa3sHKZO9CqIFQj
qf+2au5srod6U6cDgqff8jaCrTouKAU1t+ZQx/s52upizcL7DS8dNjjxadPl0Efr
mhB6AlMzRhZCum9Dl3iC1gIJs6f9i+yEJez4YnG+zPg=
`protect END_PROTECTED
