`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ASF/PVrwpN+d3QtnECnBNRnnKyOqASn+z2QcOSObp9aogY14pZTepGqkAXYWwwt9
JEvrKBMkUy+C+lXywVbKeEVY9+8V96sSxqJZSYMnkwDls2NJB1pAkuHliSTnh96x
rEUndCDokxLKZA9sq7wUWu4e+4fQa84VPqi35XIokxZAp685dhD50X0UEy42w0UA
Z9LdPc08B2qzhl1aItR64DXF12Jxu5z4vczw8zQkvWA4YvMm0ASWuZvCsX24rQHf
1V6De5bJ0z3Q5mmx/aBvrimaCzBFqYPPN9y8+n0cZFwgAFnzG84N1DLNl5nEuJSy
Axq3vn5wDU5u17yOBDtvcg==
`protect END_PROTECTED
