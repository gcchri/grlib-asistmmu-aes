`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1AJZRCoiiH9Ce8290F0kroOGKj9Q/Zk2wjQfqEh7p75fu9M3pOtzrNmknpIEVqVz
IGVkfwaHsqSFvKzr1GZBhs9ytwGrTBOWQNUgHjwOcNZVbUoSfy5xN0r+Q+OOsOhc
qSqbZ3ho88B7Ql3oGDifAmikiK3g8eZJMvQFri8ClkCAZ+/B5RvcebeFZQRO4lI2
+gEBiHD2UNCXtYlv3sD0TRUgRE2U+1snFcEgV5msgCuU3g2StyrTWyxsk+10NY0j
PJyWSd6F4MINMeYwfxeaI7oWBO01KR66wBuhHqMD/4nrxsFg4YJTFzgwsBILemEQ
P7Y/IKgYlQRAX78q1/6UnQjTSBkvKGxICTaUvwl4GXT/OvT58xQbgRvH4fFEadvU
e4yG+sXoPCN74x0ohfElfRcsDHtlrYNtKbbvN5KiX9fD2a2fFV4IThGogGEbM7gG
LZXHqGh+7NoDOugj/aqkTcEHvI8CkN4mDt/yG1hoCY6+YBvzfjPNB76eI+B/MycF
jBFUvJsHF5eGm/l2b9wOBuBktpFaYPENLMW28sYNbtM1hUsQkOjuI+wdMC11CIUX
Mq2250i1kLrDXjpr7skVdfMFNyBvf51wwSh0HKsW5iTgGtDYlawNjRZN6oC8HPFo
o0PDzPHYJQDiXtxCJGPYeem1lIZrZ+8n9/ik1BI+pkK15JhEPNvsePSGU4APLxWv
nqUoyT0/oWHG1YfBUVuICkl+kjT0oQwLexjzj4BYVZ2kxCnhBj9V/Ga/03LpxvvF
SCn1Eo3q9BXvN3ocbLygFHHZN4IYHHaynS+QV0DrQyGlrDHEKHIS/ECBQTUzxOxa
BxyhDBpsWLqLC6+9//zrHRnHP26mSKPPTWgMG96toBSEYQLjDLOr8nvy1qVVhjCA
X7zCMKduPPQf9eXkkyqBDnnKq1pa4IU7aJvzObaa+FT/RblQMmiTjXbGgoAa4Ipj
FV/NOlV4g7KUB0LY5bLRXkrcxlPXv25D2ZKhDZUZoG3yx1sBa+S9uRirkOpGuT2I
C3vevFN53RmB4Cx26/r5EmPuTbtcoiCFHx0xfwyfVR1ka6IdYFCwuXf1Ll40oFIY
+r/DDbfQgkr2AbXrBAH+3xpwSYW2I2urhFo2qCPCHh+vQBlbJez7IZAIlbfWH+UT
wg4M6/sBisFaIRa/4NXBQtI3c4ZMQ2J6k5/dhuZ1tbvmyjPZkm8wl8WtZHm2yt5J
EHRlISvBC3C9SVU8oJ3r4sPAL0sjSx7y7T9VU3pd+T2mq9yQecw+SOG1qZvg2lh0
E1MBAT9bdODpKO/Xd7yUU1FuyRW70ha1BlzWXvfuzCCNEucHFxbq46iOCFAGUNPj
EhLA1NvPrJK3x3t4XZR7/bcFLG/iZKoaT0tG+uibZhYopSU2wImh3AiWXeGavqJ2
`protect END_PROTECTED
