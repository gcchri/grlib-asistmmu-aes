`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6f7lg3UQweZ7lJpEt6urzIC1YrIpX6IirsXqu0bsPXIj6zwFsARTbRAwYnIppqc
9UOAwk/3+axrGTBlZlPqFwEIWRkQWFWQeaH8AxkaUSo3pxysxj82unU6eGrF7rtD
aZNV6R9r7SkHCkE2FTIlJZ7mpthWFT4NX/KAXG+fZsoUs/G/P2mfyXXKGWEs/CCQ
v9IIskH/n6TwJqLc98DogNKWsxFuBqEUcolmn/BSg0VNqoC90og92lCoFrWOr5vl
wtF0EFEalPINzlHp91mCasfL4+4qfy/BmBmQaqnENf07bBccy1LUuYF0BtG+JEcR
vFrGBvjOf+xzPChpqHwOgrtetKWh21vguOFKF6rjNW1s7lMHwhoZdi4pYNnW2s5r
`protect END_PROTECTED
