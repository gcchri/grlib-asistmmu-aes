`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rq1KoD9JPGIAuTmSZZDpzBjELPIvMTW6hKkI0qRy/h1qgx6T9GT7rLfSHA4hqp19
ykI5fiLgFtLbGlo3MWmyhqLUCh7tLngnH5e5qp8gp3eL45fuQdzf02HjSIqbDTSC
ZrJchNB29+J7bm9piZm617WzO4YXWH6mFzs67hnQpI0BHjLo8cTOAXVp2EGlTNgb
Xj0sqOExs+9ia64NdF1Zq9WempyW+8wg+MFLJojWh2zw1U0wpcEBh3uhhmaKsYZz
5FB/uFuyM9z1irb+cnEqp1g74CnpnAo9GxLyQ32y7ANfW0+tzLwXicqO3lM6q5Y5
hyJEeovWC4dt9RRbomW6bx9Y5UGpehee58jEK4p9Fhb7P+3KVN1GCpll7sD38mT8
z9qc2w0M+WTxcDj/IPyYuH2B9lQxH+M4KPYvO6DQv80//VhHWZo5bvy1dFwO0/8O
DleBUCjrMIrzIvB/LFuVEdp5PYh+P89pBE5NLQrNi6im+oQvKkwXVWqHf9Rw6u+p
15ZeOGgTODK5r1i5DG9/C5KCb2xwPWaOJHfxybEiTtUY97MlG9z8/zIN29/mveeO
NjVVOat0ZVE2xYmBT1bAYUVxZtIkrkdcVZgG5gAmht+zV0Ck39ZKKSJz5li9xPRH
e8L8fS7R/jA9LcIaT6DlzbnPFomlb8L8JMDDhAAu3wkCHtolEzQICdMIdtib7dCJ
4kQyFnYT/2Zi/b35qikhK1PaYlWyKiI5zibR7bdhP5I=
`protect END_PROTECTED
