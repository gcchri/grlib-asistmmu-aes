`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vE497X2D4xuvBC2xdHsQSzHpLNPxEtk5spDeYZVxY4Ylgm6YS5eXOLOQDz5fY+z2
2VXQrZR6eJAEwFLkMmnWybCQ0UOuPW7d1iC5wm5i361yev/dWho4zYRKsRk4cgIY
hcQ4kbRnFJ0D3EDbLkYdN8qXzeOfcm7l3olB+VCnYUil4NBg6LhnN7bWy0atyMvn
YwGb0Pf1cSX64ucABJ1yO+pPbfhfE56R1ZY6SQEe+CjUy8ZqtAH8wnZy9vNuL14o
0qfVLZCs+60INeGpa1ntW9o/98DGCNJbF0Ci9lCmMr21QkVnZggIltOGsYzaMuiw
bJ/di8TKl74eWSmr20mnpoBC1EM2TIMDPV/FFWhty83ja6fUqvsrNHXchxDiQSVE
LZi8sfoTaJDoBNujBUXOO4THVTOYQXIH4e7ipR8uoFo=
`protect END_PROTECTED
