`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qx9MR7iegik92aT2vNE34EYxwquYdfG0dSZL55Vh5DSUukIioCvRZ+RONNaC3qq3
sLlWIvcJGQGaYoZCR6AFBLvzN1+xJki4VUxbm6owF7Y4h53O/tInZQwI4wHnguWQ
Mb3mHF82PQOaALp/B7mBkuyYkhEh43MQSVcH2k3h6OqlY99sK98goYN/Ve/k4XnT
qc97BwpzPnYPKhhTdym7TnTlj+293M7ozf7RJih8ZHRg3kMRky5z8UZdvfYaapfA
ZNvU0zB3SiOEAKeLxGLqZfHnp3fDfTuLOa9mdbxXfGUkwdYe8uU0p8/30aEjhAxL
/vz+6NT/bCTMMUvqPwJCEx3Eo+AK1WflUO8ArwOFn8upIMsmhLrYxhl2Nr5ZVixn
YoArbIoUI8T4775oP4+sF/8pVtjx0N8+08NU/V7V6Cg=
`protect END_PROTECTED
