`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aiGoP8n7Iv+avgzUUFmy++0X2PR+3tleT8MbTUZn110nj2pioR5/sKvsqtSkI2lb
PUp5dhl+3IsUzIbjAKs7VBnoZ4Wjrd7L0YhBy4cQA+n4Xdr1DBF8ATnZlDrpk08r
/9tIOesSWgnEj7do5uk6qK5SqJo2/xKcktYBrpEHej6gOlH5BGOy0MedhdGgos/7
E9cLlS4jZQMQD8clnvPc14FCFt1oIBd1oQUCTK+PV1prwOACvmHWOHRkOEyLIKhc
zs6MNvZng28eU8WdwFOUdzpQYJg6jGNmud1NT4Y5ZSVc+tsCPOGwrtxENI0Io+Fq
8XDE3XsUZRmS5L4iWMMGkbDYs9PqeazJZ+bUuBFPIkFTUQ+s+RdJ+WW6d8rn0HWD
mv5kRMT7Et0nhoClmkC/JsPylRZdGhHVyT9wlh6VZDHrXkx/aEb955rHMOPLHVJc
pQizVt5jLtSuPhs7A0x0Kw==
`protect END_PROTECTED
