`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUa19YKhhu1aspRkaCHLc1Nm8XgtKpnZK/9GYLDiUJt+3/KO+6ayv0OjGZWHvfVL
Wo7GDYd2xFd3vfTAe1x5G+UpUouFc9+AWLdpJOg5Hv8hQzOjoTVvkVqZQJTKKZUc
/uzc9P+uNhrltBokxpybl9wCXsXECD+MIWf7mDUvwiiZLmoJPSNND6Om3coHHuYA
7mXLYPVeWn/SCeoi/SCoI+yV58WeF8NT/7zMpSKdGVgg/3wDQ6aUkecTABVHTkDM
R4K7E8EQVGIZKEv9gBAtrulyZxMp9+/40HH7uxGYUsW4+inN6muZksGgpnxNLRRS
Aw7kxUSIeSOGV0iH6ZyCK7kTwjLXkEaeV2dCIZ6cHBSm2AtHEQFw02R06v0nR7GB
a9uwH478WoXOxIYfcL7qxRsvirCw2PMKrHdRQskQwGhPjj0NM+F4N2AxgTl5i4FV
TQdeZ0PgJetPfi5zAf9iJbn1wWSPRXW56gIzjNsB3iy2xGTxDZwBEoX4SHYt0/Sg
cbXSMUf2V+T1FFEGLygwSRLcMwAe6jrOfqA6ztI6nwMN3s9z7ixHI1tJHKKm56CF
gl8IEbkOIG09GhFR7LmddEW6uDe89gcP9zA4favnCOk4SiWEBqssAiYHlJovfaB8
4gmpIntKOBxxZNJbAj8QOts2mBXoTq3PrH6LYnJD63GWKsy0DFrP7lgbtfleI+Be
CDt4/5PfBTHTPKq6dIQEqSj/MzQSbM9IlrfeRTtpR3v6kd0QNYJjyXggZ0bQwPmn
boWxNt6BEP6ic2ylFH4Oyk7FJ4OH4dwHP7RD6f9CpCJvJsm4P4KHcyjNlRta04HY
nWk99G7dT3Re7wvlpCZBlDAcIvaut6EKNOOj3CeSAHHZ6yamOu1r8yjIWrpMVaWl
DGkoXxA22ppQI5uCcLNB27UA8tI2v1pBl+oJYj3ZA9QOS0bZqa2yWtmeAd/1kkGk
njOwBRSDqvOLwWYhcGm8l+L2tEj8GvU1TFAN6TXeNsi9NcaDTGpvKyToYhZPseg7
UFolUFYz1222AIa6gyRmDXwjmWEzjO0OhbYrO8XN9Dd29ectBUivYMAoUnCqyG9A
7k5u7pTolOWYVp5o6Fq9JChtwvp5f8uKxNAh2/NSkOO+o4XteM0oQthQZArNPCw7
p10FndzLEqMTKPbOBE38Zg==
`protect END_PROTECTED
