`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xewrnYn2RRdEQOoE5mVQEvJFpFJePyDDQ/erjFppkPjtGW4MN0I7jZPLFt0ONWGA
l6iYYFRGsAvoBc1OT5TwwBKxcR06Fwo8jkugIXWEXrbwQTHPfk7gZv06Yt23UHpS
X4+FlKez62udkiddUrmBpb/OJ2X3OG5OA/gKECil/gRUcsOcfJvcfFAWkgCgw99Y
Rdw2TJUs2CHCMsgCPrV4irp0cIRY3J3ZZGXiEpFghKmlTmNQRTYy6oSc9cB++ugu
kywKeLnpS7QF7CiSDuxUOEb6zKNfb0IOAI7S3/cHJEOAQGLH/MFheIciIcsIWWf4
eLsOkjcckmz2k5cQkQi92ouI6uPTUk8/hbnvAZw00BdTq3x9bJJUKRpOUOL6YkOD
LiqaSsmegrAMLqvwIe+aCciZ3yORtDUmuHait5z2Abw=
`protect END_PROTECTED
