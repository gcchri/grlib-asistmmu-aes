`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsNifhyVi3T08NnPInybbG3EBiakeuU2esKKG6gVuy6r4+TpoWyTG6RqeijPWwuk
+bVuiYu7crVEirQrsf+MXg7jggykQgH0CZvPlpO3IOHkDLN8cQME8tCk9bXviQgU
JJV82Oh1FrLK2phMkHPxQXKCUAPcDXysA2vAFPVZnrtJvMuqYYB6kepKRHijkA69
yJWjf0hO/QNv1LdmOvqNhwqwhXZtpvIC2kzhMmczOJDrOJcH7rf7+M9p4sjE5Xjv
gIXZoRMrwaOTTea+LDwaP1nHUtdY5p4OXC5yd7bbQJ+CPDyI2wFXPmzTwW0lZPmP
ftpawtRAZ3y2Ki/XRIbhMqn6HyZC2skKsGmiVCvCvtEWaV6KH5Kpfg9/5F+39ot9
E9K/E3NmGYkt/D09jC0+rYZsbazYX6ndSDD8zTmsofpo1m7l7NkR9wx6Rw3w8z+k
4KzkpP1Sn0Ox4hWgLv+TBj0JfEleSiQ/DvvpMGEHLB1/3b21uZEG42ixLjGFrkY5
t5IEPVd6WPhGbrJyfyDCSl/VqD29aBaSLKAekSFkvHa60NOq+OyVgxDpWL6n7nty
SLe++61T1QTQCD+wA7mEIk2ibK8329UO3RETI/5aiW+V/7Do7Vtqz7abxyRklUfK
ar/4rpu/HJpbDSmuphxerQ==
`protect END_PROTECTED
