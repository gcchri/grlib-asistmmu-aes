`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HWmcg/u/KVJXM+a+S2j1HmVhkAso9O1N8JGVLzikOXbaSJFp4BQ6h/kACEfBusBa
pEBqreQ1jC7mWcmcthON/tV4jR9EHh2jXJQER6IW/KEV1Lpk6vBvNwDbd8Jq/vJ3
DkVoUWZVyJx/75x83NigaK/kv5nz7VSN5UmVHD+0U1IiKngTkiknrq3/192RHDGv
qhJbwRWuCZ0YImOjPWfEPqQciZ9wHSQrJBkhmeoYRCQJEpQg6nd7icsZEyPuXaoI
oCiqASzTbERpMta8ltleefrZAL6DwxSxaCbxuu32FXjFxUx2nZvHpvgBNL7BEcCd
neslSZyz9U6tGAvCe9v2iO33ie1pLFZ7K2UKo/zpVOyE8rCQ2GwynTybCGBDkw+r
RCISVD4mB5BqPZdInQjydBGsm2QZ15rbXlUHMwqtBZ2J/ykSdNWOHV3f6RHeL7uT
xsQ43u63Xrng9gwgh78mRsWctY2Hj6t88MRD0z9TmgooIn2F4Rrw3b1Opar/tVWO
3CGIRiWV9/DahuQRLOlyhk5sB6wSKU2H8ZaMn6uF/VmsT1ZtlAdfA0i++FfkcUML
avaEnZMocYQ47hFQcL8fD8BOnxDkxhqFYbx3HCJRm3+rBjF6xtMkHieB4rmFa9zp
U7mXXVLaNqzOlwj4yOwebvqVJkDfSMRiMMthW882chazoZzp3pdN9o7CADF0bch2
8SXCejJJSzgGhF0BZu49srnJNNnvmbqA7KOfDRG3eLHFMtDFX7pca4swpuYqKG7x
tFRN2j735XJZXilsCoOJjIxCUEklrWCOG+u0himE6r0BM32jixJWg/hEssaREDc3
lpkYXe5faaFsedDoE2sQaBQfxNZU88q4KH4Q12Q3xS1ctqOV0Ac3dhkVKFL76lXu
vtgDh1Oi/zEHguNvxGTHf6k9YuH03Oikgw8CWQEiOR8MivwoyrJW6M/h6Jjcbvwl
OsUBf3CIGUu53cwd0qiv4holrPuRe6ohOb82V2f0SJuApw/jLuCRrfQuvnILgd9O
wT8YLltBNe27tRC0l3KhGieDws8oT7vStBeGNhy0ehMkiVNeBO8MCV8qXq8/BbK0
qMNti6YxK7UUDxtsIaxTTvLEZS1M/nxaRA52hZhZG2EExrtnkoyNlpLfsKze6abo
lOv6I7HH5RmMvspSbio9u5Ge3D/2RsQIVOFlZe6tmh3jShi5lZdqvZ0iAnp/xMsa
gazLesx1sKMzORqjnTtv3YexDc2VzX8TKSgZphNCNs+b/Akmlx7dgWEgPSjlT8U6
ow0y8SfxzAmY525KHYG3NAK+Bot8psaa8QeleFK3ijfgoYU93OmW2Z24R3w7dqLt
H2T94i4KoGEpjFwcZRGxX0qGqFF3S04Umv6FnzUJSJTW9fO6WQeS1tq1kAsuHfb7
XpSRWYZXXAejvyf0C1P/DbRuKmgZ7SL8hDheLaPYUaFHfe/SnvpnPgkXF7R2vdtG
+ItqNponsHQws8UsKGfrdM/B9mB2PTeBjudbIE1jqj8TTKj8DNyE/U4iTIVRGcJl
16JTli/MTkVzHRG1uEWgbKlsIb+7LmMNyUlJLnetadFdURLyHBjodKF0D80HSo7M
d7pDZvNxiRhJ+n+pxv+w/fNgbEVY2noqozUc4bWJI2t4HH6fz5Cp7zEsOO5sek+g
b1FL7pLU6Ms3kIidkK+9zbdP5pZ1ewFxVg8A0sMVm/pi63EN+MR5afzxmVF0I0E9
wcIeL/qgBIt8VRgx6sBgA1YXrWQqwblWEaeQExk7VfD2gVQ2ohCDhe8awPUaVLNE
aL956dbo9fyF48K7vNc6tOrn4B2ZFxpul4RkYkEAL5vPdZ2E4lw1O34vuVxpp9r6
ppu3PtjXoj9kRYmWA75F9BzH6rZfqEdez5hmzm9AdfTy6/fyzXR/byDvqiXZJ9ck
Ez9gpZURuGLRR9TXzRLAhdyE5Tc2kPYqUbh/uj379rZKOP+kJJsJLIlS2RH/i8cU
moB6BYtLVGBzYZcaLTrstzUyfYu10pR3Fq+5a+oh/5/QWBpi8QYnIal6k/mNzL6t
KchsmSv4A5/TNFV4Y0sYZvG8KddxTdVgwV8Fc7PZzfDqgjNZfWkxIz82cN4n2H1z
87/XTJiwHik9N+DJxylw0C5sSt+O7YBibrg8tC5zokbQTpEkdfxdzpGhYFzCq0Vy
yR/1dzMdcDdepz8368e+AsmEZ0C1GJ3BHnLWX/WOujPWK6/+IyWd+UN5m3lJPPUP
zrV6Z+lpd9sWH50OWVcyiob929Lmn5oXuw/UHLVm20B/zXYhswuyxtAp57MwlEHZ
lZND0iUGM7xzcuK+y8xc5cJRKy+V2aDHPa7f/ZJizXY/LcjKaa5yUeUM8OzIwFZ8
jefow8zY5IOxVvloZPLje1O12pHqOb8zXQp5pJ6QPEoqhjLkshyaOksHxlWuMx+L
mIPO78zUxSaExlbmWarKK9L1iA3DGM22fe6Pal0yGw4qGNDaf0EAbnxIQQZ0QSZU
sGKtjkGlLeiYqf/jfIWCnrqe21SCtlffxbSFWaXqy4+6IP3JnsoQHuRVjg4HEOcM
O4PY7VusEDgXakVOmRejWsahiMTl9VBAS8XLwVj1WY8ByEFO5VwOj8FE7hj5X7ik
PiiKnSYSFBXrwxiEbpRbHCCqBmdAdJ2+2+UZFLNtVsO+co4qEmmt+WQrDLzbdMcp
p9em3UdZpEYxNxnyDtjh+TRF7uvlpJCP06sCkNBm8es2YieFA9p/S9/xETIbKTLw
aGhQx7tw45dSuQJTocGrKK7b7h2GKoZ4m5E5PBWoeZAE47QI/vOpxM5OlGZ7NXNI
lqYaC6IeTcPYvTf6wFbp6di3+0aqSq54mucfN0QCfsNaMD56MGHYa2oc6MVIEmDM
WoU6aWJtPlLirFkvpxEgf5QJkqVgikuhmX4EWkD4I84xA+hQ1fPVMI2UyYxO/LNp
XnWe8dX4dSrOJTr6rGpW7g+Wa7cvqgZc4YSCBS7jWt2NGfuQRtZYNZaSa+ODBrSz
NABaWVOz/tR4Yljt3f1NAz/SS8Mf3QA5o5ur6t9m0bGYkbw9xrvMFidz78kxyje4
lNQYgm/pLnCDkyZ2hOEluCaCA/IQrtgnltRZ11/oSbj4VJKmaOyAckDJnI1BQPYJ
CwaqKQ7fyGHvzmF1cxbJU5/p8h4oaZa74MGtLgbCpW3d73P727p8U3iOuLzUnpvA
vRp7gIqB5zCZVlEljmMsY/B+R1IWEFsyMeiKu/oTcj1A2Cd0rAydyCv6EELSS44u
1Q9Bw9asaLbPBn6B7qKRw5pgjCY/Hne7mKFm2WhXFGOQ8xfi3aOKGOyIy1JzF2rT
+m1link68ohbAZQ8Y+tew427dQLjeN1dQ618Zu9nGsc0m9GSHz5usIYU41jXE1Ud
xBh3msQOAyYKE8opaI5eMzUzkuIMFO2I4ms5X//9vEwfVer4CLzu6l3K8ciW52eP
TpHmHIArMQ2B159Zn09gx0WzG5tm7lDThfVB/vNMxhxYACRh/8U983ms+9dtgfdZ
TSVV3/N8id4uRQbA7rs8zzrXFrKH4osJ2LfuZoLveoGcypjnWkRWXeNl3FwM04p9
8Oj2Eb0S1GcfZZ/Q732qJloJKIrCICq5dAntnk1V8K0mymnz/+b2Bd2l7kpi7Jm2
hQXrl1xAmC+X0yZQY1avN4oHyTFQKQWySexR8BQJHN07KN8mZ2xw85ox8xndC3dZ
NXHLyRTRL/jKOSFOJuqxe2dKw6gn+Pt58gcMCR1nrlMko2XeoiKf0ulkRq5hB/G7
LdLl92L+0BTDRhzoTRgpx4lbInzc0Jlq+ANhYzcKzWLSJatYDC6kAmlmg/zvQSPf
2+gaSM39Kj8XkJ1Dkh/yTo2yyFbBJw1cnRMTvohkD/vdRdrguhFxu433ZF6ATkCf
/by+Y1A10yYHnx/fVx91Hw+mzQxU2IMv7OIkWQyvTEd0NAQL/TEQUGaQEqwZv9sd
p5vM4Kh3hb/A81RXnev91PTU6xnZXGS/zczT5vqUCPrf6ptwxFu4875T9BYv3aVc
8VbCVUj2aIzeYD0WzYi6roebmdfiEo5jjHQeLFIlHqmkYLcI/fzHJBVYsD5nxAj0
rMp9UBS3FwVVwdCGGMo5KTwF3KR1B37A53a2TcXeKqh6tHUwC5BHQfJd5bjhaJGp
a7vjFMSPe+V4ozPBQKKTcreknPB4dnyiuI4D1a6rLhd7rLMUfQs9AY9wRZ4IBtS5
VVjjm9QRKH0yWcHxSAtE4nU2PUoKB4Pcc7oLso/ZEnJIOGCfovxndDQEr/aYNhMs
rr1jcJYmsDGK4h3QYUjzzYd6vhSxf89Mlc0m8twcw4qxWmkC0qy3tjC64zltZORS
jXZ/hljgZI2MTPmGMvxVmU0g5LonaZhTUWBr9ZDyGaq4CZLUfLtsTlgQH5hdjTYt
VMAOUb0m1oFHTkVKN6hbT1li24mPSAIWju8YZ9Pu5vYlxUUYw4RpnVZ6QH0dqzIF
5RDY1+DKnOYyEN/edPVdi3ivvTXjNghii0PyydvdFaNoH4xZ3grOHcsTSHzGeK35
AQF6tG+7KqTw9DIWHAqsygG1fRZDpS1EdNsItvvTsnVXSeftIuicXmjms4kHVjIP
SHGFi1SlMRLkRZfSmR2Dsr9binjUAO/ebPvybHapBCOy0AJ7cKoygSfWvEP22WK5
CWyk5Kooa5arH0vvV6vFS+H0wzW7D58r8K4CLlG/BG5QRXgUA8SSVzC2LNDgqhyt
c+tBhkekmqlr9qoTRSOTF9U+btiFVnJdHPJN3RY9bTEkyDD2r//4rXHJ6996tocs
ziIyEvOUaTaVG9k99YK7pSV31XKk1B/cS35Hi6H53BfoQGGPG6QxKS0icEqnDPWf
a39LBqB5v+JlW68uFEVp6rUCjLA8RV8q2tMwrOxagePGGN91jRKnPGKzlz0erGQ6
YD5PjsUrPDjgwagyK5ac+8jsiSSRPebTFXll6Cvjfj5FPC1gOtWOdwbY2GA1vfFq
06naq2PoGRM8JCHMq3bkQFJeG8qiLU4/gWau+bfJAEe2N1opK1RS+0wS2vR196+0
sv4bnMHTF6gRhVJ6OP7sES1FVbYAKlUdPcJJOoaWNlnvpnCf5vNto+VX4LSEI72y
QPIndkXEl+AP+ZKUV9WBWtC22hT9zJbnOCu9ywgvtuy9qvVQyFP+6nu02VCpr+H5
ZuhJ1TusU+bEK1IcC3gSicFPZD2Oq9fewwsOi9RP1Bqu8/QgwC8Aize3aRFm7hY+
w5tWUnke0wv5Em3gNt4FQUsgNY8ntH35X5ztliWOThO0G8P2jP71zBCD52Sqpwqf
jrVriqY7qC1BEPrG6TRYJxNYfzg6ELqk1/cKwyuSWE6+Xx29GPM7/bMaUmuzNhZ6
WCTJFK8HF/voUA9TQ8R7qB76dgfsFtZHIF0x2BsvMngVSvsqzs8VKdvly5ZwqWMg
2ktA3/Od9cRfuX7xL1EcnuUOW4TLV+KXMlvxNZeKKv4euPTXFPLvi5JQ3/IsRKb4
YjnYx/rwD101RiC4cdcqGE/1dKqWIus41EfBkQU7MrfYhJcdHdi+v41W8fOi2Z9Q
Lsy+x1ZTUkTQpo8v3FmdazqnXsFG79z0l9N8fUKWHuWMaEEM3CY6XFahTFkTXXUG
EL6YDMixdscMPEnkRf2sHarRopFRcCVnxNSEfIULm0vGwmnkP4H94amhmqiZo1hL
p8hVNgRzewOH20074WcpmIAWpyypTShj/Bi8JELKxLW7YgWoAuByAOKF9I/zubbI
X/+7zlUTAFe9auk9wD6fY7QFWxvP92gg0YhqlUCkfY4Slahm9T2w7kJJCpK2Yx5K
cJdbPXAvC5BURk6vKR6fi9dezdXvus+Z+IeBY9IqGyxo9tyPLN26A5595OpNPsZW
lpevQWxANImbu8yJYdBCasxZLHoV3Mg+yOyj7aFEVup0MgTw8Fr1nSb2gO1llqG0
YbqfVptfAsuXTYLJe00APlrttG1kpVWkqdSsMXJ+GbUFuy9bd3pEeTf+tAnoSTtu
WYMen7U1BptVj3YtmTNv48ylevyD+HWupdWEL67vPyl2kIlFKdkFTkiCjroAlv7h
WPmDB1J1w8JPTBfubDzU2eRIgR25d8/dnmSc1BAYQS2ijgMUbseIbNCqd+v2RJLh
BGbLnS+rsjzUa0X7jvIoSrl8/z9E1dUyWdJMY7Z5xXHmKyjxeEu+shPR6mWLwBsX
oZpDNhfvio2x2GiZMm7lIRqkBbN8qTm3S/xhZjClahwCXzL/Syihc+8ffl/UfwBb
cQxvUCZ7IdJsJUIfNQK7evm5RNSwyQ/NDEseM3VGL7HSLp1NBlzVPrgQbdfB8HEL
0giRtQqSpF2mCwkLMNzLNB2zLKefCHOMj5R7j/ldHA9zRhp74jvNTSC6/JEzHgb7
FJXDNtMZKy5zwr0qO/lclGZIF8n5doXhpN0c1H2fLhQxf1tNqp7Gh63cWDQHJiV1
GLLkmy1oDW+jgWU4/vIWQZzjufrP6eLpEcqrV0lwkaOzbDtiG60a55AWlqFsfEc8
+lVrSqHQyMFhLp7n8WxEgmpjPByyv/7a6ISDuE+Z3J9/hz36UBLhvPDHoUi1ijQl
F05CxuKp+AFHw+5R7E8XhMhRxrK1bJzkUqUBhD3kEBF8U+WZNumwYbvvs7GysNcm
ss83724sN5vt+5m3DQB1bq9IQU36gvQUdhDuwAJGMA92yVE0zqaEWYsLpqH4WIvN
Xu63HlOPryUOyKJ81UFuj6gbuFMhQCMAnGFCYCEUVyMH2z5KKYSLiwCtqI9qNCa7
aBjRIziREkQaWwbNqRA58HZd4+Xbn7XZVestR7umr5s6v6DaD5HL2XbXXJTRKQeR
y1S0ugjwPQNac9L2eDYzmaRSpxWD/z+bM1LfW4ZyB8PqoCy9iFdXAYJbyiK0pQET
EX5zdjJggLUbnerEGlWfA5YRmq+F8DaQsGVOnSIt5W2BjRM4WdM/RdECiDQ3QHyP
Egc7gxqyqJBjHC/hz91heTx2y5xix34RxEfbg/naiQK2eQd5/V6lxNfVueJ9Ckxm
Snqr42UWEb16sUKoU6e6d/u7V62pCiQFtp/FFAGDgNhiwAf2CnSsYcpWQrBFSXeR
614A/roCHdULlRxN7GO7qZT85lAkY/gHOHWSROK/HEzZWbRbbowCR1BYYi4m5rTd
7HYjPZakVz61f5B5IAecMPWGGLevIZTPG9APSwg8ktC7o3WNC9Jt8XYpgIgeu4TU
euoyaPc5mffKHrCdEFaulZTjT6h6l97H5ZLGofKnDWzQ9bIRwKWUvEICaMn3enp9
az12dwqMvUHrNtC08NYSvkZT/dSc8y72ogtZVDq3pmLeHKkI7nySk1gL0Jf2PtkD
akEEaT3z71qK3jc+w5vgTiB9qDmGlC5cY83wwuMCzjhgMWU6CqWFUSN1KC7nl2n3
o8wvR/NCLoE7P9CBCAXXYktF3wSySZ3Y2pvGW4cCcs+oqmzLZ/OsBeLjxIHddoOv
kmNMkFG9WflMTgJ1u96oXodP9g7AsigU/SHQOr3PwhD1OFvDkbg9WHcLT7vNnyHJ
+YIZ42b5GfUI7D8eyFf4M4Mm1+7b3oMbzqUz9wgYIdAv31fkmHLRE0USOfd1Bqfy
fUxnT1xjWX58Ab2gLOWR3EvSvw5RVGgie+r0FeEJlyjwzWR3hf7KnWY6v+cAXwhK
2ub23THB+Cr7E2879dSO+u+r0DZu9MecE+FPebXiiromliIxR9WUg5h3CE7JfKbH
KvdQcJxwzYCIB+sxb3CSYCHtKVKG1hBR3t5ey9hFlCZ/TsYB3AzbFuhVn0Ucobe5
9I0Pw+WFeZWSJdMckJ9GKXpt0b49/VKnjCLW9nKeYIPW98rvx3l3A0xCNRsaDEoL
MmmP/8KFPVrRqdTwWx2Gq+wyJS7c44QDycVmpvNKc5yHeh/5Y/8j4t+k088HWI4N
wWvdyDkJwcYvigQi6Q7nR9x7LECfX5jaxtLsA4f/Gf6PWUXn4HtESMeqOgZkGcQF
jgzAKiKlY9wDR1Uq218FqffKrihkSdAhhhFsO5UlJdLx+FsT7XAStmv9D8OgDJ3t
3mUq/Tc549l4bVTceOWxlIQepdLmq7/HIcrJi1fqrHkELmedOpBb3QVOKpdEpLno
eHdVgX0cBxJn+XLuQ7dK/kSfljjYtEJqgNz3WasrEGhPK/amXo0nKZFQJmMXyOh1
V03MHXYbXE0nYIF3sQPHLDwf6xGeMN8yqU0wR8rdqT+tXz6lXO6MnHY3K0wDDRJf
K6dapmyGfy5z/t0H27h/hjL5J/cHfrdL+zXD3/80jofT9v4lk/zh5DGxoycvVnSm
ew2zSfMx0F9rACd0qt8cpsqKBVBy1JSyhyKYgBx9j8Z6c7kiB/gWCW09HaY7xysJ
j5Y8JloqdAFQCRjtI1XSwxVS9T4tBNyeYGLAux79amN3RjcU0Lx8vLf8RXRCE+zl
kLkVnS3HQCMbOOb7T1y6R4Fe9ekNCNORHFUnnet6N/Y+uUcj0t/IDCFJiVjoi+Ts
GP9B6RXK22uD3kH/yNRU1rDVoGObN+4k9S7BevbC5V9lnXYlarYWwj+06JWlL54O
duhiJunw1uYcx9LF2eeKrRylIDsI5AIKuiDNMNIFuUfw213B0AOWKdh0RSiPJO27
I1qiAkOayLQ3s8kCzbE4Dj3DtWK1dM+E/O8XCPX6NqwmR4b6oi9xGPxOBtDTs3LX
QCjTNas9wbb+UfQS0GbLwgGuBh1zs0ea7wQV3cTPloebXWUqhqHDNeu0Ro3ZY3tw
b+DKYIca1iS0i6eIlVM3BXtAQ/s2aqa658nDsxZiABhsOpcNoGRH5KR3iNbHs60T
ndbNXEvB0lmXjMbaiuXPfujJ36FEm+SAnxZS0mvtZTAm6UoY8sXZ7R2ivWfVqPKH
aeUXEst88Lyc5aGEzf/50ptjQyYt9XL0iM58jgxAWYc5CqG55927L2ST4pxqtxlR
d4yn35YZvMR9VHwOF3cZpqVHe2IfAFYIx9m1M5542rLA9yg+dzW/GVMsiP3bydKz
4M86U6igt2pPY3B0x9xe7DvK+or+heZBuzsxRp++8c5AawgN70o4VhbYu77tjTqH
xE62t51hqDuapNAbUjulU6/XeHNeKK9XtGm6SQ/viW+l1SkomOmCrojN53kqap46
E4eAyAWi3V9Jw54UY2Juvm7TIJEooTSFSprNcAlsBEguEJB9aUL30WYGEFXhU072
ZKij4ND8tBFaXjo9NZ0dpMdAOzW8c3EMosRqM2hzl6yW9WgNaGhEdJaXXSOuunyt
HOVteCwvxEb6Sc/lflxwaCZk5DbP87EZWyTh2x8E2qWYK4OQjOZfvZBDIwj6xwct
8WAoM9zQXJLmevMSMak01aLzEttLCxNOAFkxuWlAbZt6JdnD5LVDfl5/S1e0rAfm
BF3IMgMXnntOSr36hMoXFkISHCt3G99vjNVdT/G4GD2xnHI5P50QKGBZJ52kSZHQ
HAS54Xmc4jj6jOUeW62+aHWCrGCfv1Ft3476DFpF7bavV6xp6HjV2XTXmVxITiAt
Ss6/3ATS2ADEfn48A1u/EiM9ZGZxyeNEVso7QFP4mIgoyABegj0uFS7ez+TM3Wnj
zm+lF25o4t1ZrFpclca9nYoE5HL8n/LzPxCiyomtLr9Yb4BybK3hpYYkEX4DUCeY
fm+St/WEB20nzjdKLjqJlGq7Mwg+9tWf9b7Y6s+/vhlhtbBn9cfNj9/a+pbJNitm
wMGHbrljrIbiycM0Ecj6ULxWGzRzBTcqHyUSM3s4x39XzboV+2L8AYpK22H7NwHO
WyPZ0RG5hs9Wry/KMdUkBqP9HH5A7mbCq3vNZhnWYxP5Ftn/KvBTL1U9gaD4i7Dr
Qu/2gtDSUmBN7hqeBx7GjRjk3M/jOGK1QJL4c4AA9wpBOlx1TTN+TgaEybKOFgZ4
G4ov1yG3L+xU+9rHiE40n5tjequ3buPkk3fCfxqLq3P8Zsxr2s2WKRcJWyxAMLxA
1zYja9PRAUdNBZ/+/3yXJnBUnJsLtVgxI2IjyjdPlTzl/QQG8bcj3weDedUrHi4L
/dF6w6ilc8KrfV+3sl+qcQlRHkEyEVPBU1tTihVEhdQPWyZr9t9BKajmbHHN2YRE
zu3VG8ocZ//evW2D1STlBwz647ekULoO+R6NHEqce2qbxho5hZEt8BIRCKNhSLmP
YII++NU61OUmkdfrNG5o608MtvVCetclxlpGh4a2yB6MA3rhL35BniiXzt7htk+9
NPl7RhUBwAvwr7ffKlVj6l4KB57TL+ZPnND8eXDDbBDwWgl4TgTvQtf0c3dYCwlw
mguM3iGeNBUnqwpSWwJpeqbYLr+TSjI4Mnk9V0pnbY70Ekz8SCQaVXrNvDBdbKdz
xM9MERAj4vYZ6J+EhXH+G91yflTGQhWer2CTxNeCJO3E2gPJ86sKyhw8qYMGd8wJ
G+/9gkIrKWsUqwbc2XalSPlHd3H0odH1Z99QsyTfwnB+6r6HQ2DsUX5xxyFjzx9H
XVpm9L/m+5u/fZ3DM8N8N6iLB22UwE1FFNgYZ39M/9/tH4MIImYu4ZhzKLq+IWvu
pChT8WQ2jqvJeq210WxAglDXIT+67Ij+tmADzuGhDMUZ34UzkDZNnTcg3jNfs+8h
zS2yvsPbd8NSCVB2XeNygw+SiRdXdmYnoimqE4nlHKXFoQjz3s9/dltZHKQcn5Gw
o5hwzcntO7ce9l97R9FimtuEenY/hjCzX/kO0+HFnUyhSiVGCi5e0XR49Fi7OSaw
IWK+gI6nRLtUkuzDS3ShsZTEq6Y3tXj27EZwcnFfMfBsDKQSqV8lJGBSh2Rb4p6U
5FivFUxwY0FB61B6VYOwy7Q6fhcOcLyGpDnTFhlE2Q5POI5t+LnNlKuZf04vuGkM
lKWyE5IzSs7NKOLCiWEaayb8wXL27/BHbNhRMnOqZl64t2Phaol9kO0dSj+Y5xvx
4Lapbuw8g5MrwTdFD2y4JGXDWB8PyAF4S4/Phe5GNLk8EvaLvN9gAP83BoLtUVG8
QsLs9Faiog5H1TRMlSLg3gBIXGwGyTn31hnJU43v6XHfQ+2E87pWsHf9WvsEX7JW
EddMH6QLm3oedt43eCnZ6EaPoqAD8JMdhBz3dY3xXI2erbu8/bjrNCGumBaLA0vL
wdh/92UeRyqVV3I3buHNiu+SC2Zx3klzwEJZjM0ogQNppRIHo0rv1RGgfbZlIMuJ
hxpHxavnr43OeLh4f/aQn+vIkXq/czejyCQCdXup1ViQPEVtcao7g9REt87x1z7k
+HlIDbTKnV2XjA6Q1UMX/aXsRCqoVcpRjLu0PVQw35gqSB3V5/0Z9GHh1HO3LqgK
M5LHyQ9KMEOkOkBF7Xlb8cuIE8GMG7HDwwrT7W/w42tSn+BBJzRnSK3pK+jUwchq
hubGPS999UVFcB9tQom9kpJPyGbJ6sjCUpBzm8SHWUoKf5iabyR0DZJQ6teHx3XO
0ibXcwxo+TdvbtpYw2mTUUx4PQxNCdrrtCjNSd3Fe8mw4+iRRlVrZntZFwOFk+EV
D7hCMvQoKMCoq2LZ0+g51CDnZceYS8T1l/MvwJ2yfZTTp5f/rImRhFFYSlfMFTwr
4AxrJZkUVv2OxzaXLM7I92xmX1U0YEPUDqk6pKiBfxPVs5FwruZBWw4l9NtpqU//
KhAVkearmSubzqM3mfU3yvtEmGh3NvDSX8Kqc668VSe8L3n51foyzJdwdh9mFtCO
Y5Edc52Ybu7vbo8iUFyN2Fo44yfkM95LeRtQ0l5r8ba6vGoNUZj9Se/313iYRHJK
w8IZ83PqE73uhRvDkP3V+EKALeQMpIXPzcNv8/J/UXZ2ppytT0XiTRBH+KooOtYY
6KKrVq+EN1WDCGmN3LKEq7LpgHjFIO3Dh9n1l4kl4orF0EYP4GCpXb49QjPMjhdf
U7No2R9AKLfIJhUBe01tRx9BUgtog3hb87khK0EH4ZaNcbvucuCiaQ9fSM4YfATm
lZH4jBGOfPmMyI3DJ5LuphQ1vYG+oRt4ZyYoC922NjWUKsllV51U8Ph2Dc7mcene
sF6CrdDvyO2N6afBqw7s06ERBsbhIx0gJZoVzA4xhl7HjppXGtsCGd1R1KmMT1XQ
+Boh82FMvByFoXUgWGrbBxaoNnzgeEeIKGIB1fPRofIXyScycJURNHdffeIAPUjF
QUIJSgKWdyotgNsoKMqHSU7oHTmBKCq5LdEo9drM75r6fkYXUBdEcwKUB0uJcw9R
pFW9Rl/uqCCD/nPxhx3oOXOwq4bUqayqAjF7EJ8G5lIMiXMsWWZifDvog79P4jQu
PrXxtMS/uT7Vj1trw17hPMdj2hgnQke8pc26GF3V7BJpVygQYkkG62Ch/zEWceUW
R7j2Gr1yYBvbLBHn8yZTRqeumGsuWvsMytHgf7NBCBf2d4bH6XeX6IGO0afdVE//
aGSLsXfOQcEPkK5H6nU4FJgXq6XtWqU6QM4pKMTdx4tMK40rojJhpumwLDbka2MT
v+zEg/xwoJUXrVNWo4TWrODaW8v+NwFaMmoqDMrtJQ3uml8PEB2jKlHT25y7Apnz
5b39QAKaE5B2StVipvnu2M82WfndmKECYZQ4m3/CsrEGOs8npHgtHlP37kmIbPNA
D2/dfcWaXmd6d0QTrE6IkqFhRcKDtbvrbpfYUG7ebgk6I41FVFtsxPZZyVZPXsz6
ZLg+7+G+4b6dPqt1i6L1gQ+2XHDZPO2MKMhJorYC1M4OZIDMsD6y6srK2gy2lY1I
fAdyUVnvx4qtIOnSkc6sGMXr7kKnvXGcsVruRnlrGVUW2gDPIr2rsF1akoW2hQO2
RNxDMp26QnTCg+UaXW+iVrKNy349JWd7/UgX8BBElngPsw1zcbzSE9PGGhtvpyFu
SFGUJaCBVq5U3tNc9HPIAts0VBnXAPu0YR+1JyoXc//ZUKHLjsqPFqGXPyYveArz
RsqtX1/2ZHJG+bOpX7s2B0RNlE9qtkeGydebELoYPDRfaiX/kY1GNWeUv5eCEEA5
GFOc0THNjIUlTtkiPBZ/I9bkrZ9QRc4PtpBq2dTHCwPJabxjraO/0PdBz0sDeqOe
NQrQEVLZwodsX3UG4QDgY+56RSuPcpbMS+EOIEH6hf4R8DCiDJZDuyzoq36du0Pc
jG1ajhBsaxpVs1CG8Dar5Us8hy0HqRD5AfshkW/C1cDektMCB+Abgrnw0a24Y74h
fQb/AJpBryJ2fdXbxybLN32yUSpKawTAf9OeNGbKASC4AlbeTnw2QQ4PSgvLAkI5
nsAWdzXpFTuRAAxAyQKb2fMQNiENDopdieQ+qOYqYKMZDZDNyD7NJuXY3XlLRPTn
2M8+8ox9LdycEKDAhby2tPq3/ASy2/UAAofKxYOV9sYxK3zbURfsuPvws2uD4bLa
heQYExq7ZgEvtwpZeaOBwTOCbeQQnBTIwfqDH03VrUvZi9dqiAEVKEJCBPnVk3QL
Tc1J8FuKRgg7qKwM2Xl74CJh2irIJhRK2sbkK/41i4NoDgLO6lAXGno3xFeqpyJt
P8qlQhypZrcKsvtJVZ95ccp9LRv9U+Z4BSObNOGZk1XaPq/3mGVX2tumlPmqFxN6
v/0OhMb5zne983G0b/9mQ0uS6xlLYhRUx2VftYao3KGMEAnTD8ePsYRpP+MT6eDl
uafjPs3lgmfgr316bIVPaIDTUmyICHaBdBLYVs2sswAb/quSGJ3LzLzvLCdJlzqB
Bxb8USMYVrm+GIXSTYJwunWOEgKhcMif4bGUyyKE4jgHCT9ojBct0lDdA8veybfe
Grk8MvfdMfT3V4s+tHX7bubUP5iWnroLZeN9maflzWMu3i86Y44Gi7Mg2zQvxO24
tNlyoQ6xPdEd78T7j6k8Sd8epUjIgKCPeHP5u9hXZ0nMBXUD66U1m4g6yS2LeKjd
zr+5WusQQ+kFwmiOTDU6J1cep3MpRQMcB1WpPuQ2ePnaYpwSppJdAfyk9k5EDTGp
guFiNIStLWT/C9BzSGYV0yLnllBIIhzYFc041LyNNMHBVnLO9hcGW0mFGF6MMfR0
zuUwlb1ZNVut9zlvE1HxVKzpv5h6LUr2GuSFeqQD7Nb4PlNnZbA4qx9gNyOgw4R7
oKE6VGqIMJNejXDpwtVeKS5Atn/MsyuxvisKbLZxBA19v4MIKTugQr2AdTmYUp+n
gkJubBd/TqFp00UqBP/HqQ5tBvLfb+0HoyEQ93FL0SaZYqOLIcr2lAey5mox1O4N
MNldTupo2SVfG+zSRkbPbuXXhYSvUU0YMYmipIZMET4N2sgXOUwKmHMa04vGSZpz
ENaK+tiZJwFPmt7Z6xKHqAWByI0UfG3u4dD0WDiBKWRbeVjiZDg9zK9Okv6dNJBT
0xAa7o6FLihyqte/MGKTiD7ndLVs0sppV69rtU8wO4OJH7Hjkeu3CdVnPLzcZFgf
FJUbcRDFjfo5Ckdf6OMB/6WL7afkCGi1yA4Yew6p/rb2toaOZBj3KtwPtlob+daR
LHcUJ0xsifC7stszXg/VnC8CxhoggqyFNz0WNcsjvu+O2a20WleuhIvxX/cfPITE
f0vQdCLzVFl2p/qLhr2dCJtjvp8jAE7yTJAwnUwHb33LVb5lTzdsQSBBtz35O/Ne
mt1FofribcdcKOX6H/UU79ifZBRZ9ZhJCDJcXXrqH4LZci1yMQBf2zHjrKs/qYMd
7w3Mw/Z4Bh1h1BZKGLpYnD9WG94pAuat7eGr5qpxryicS7/uu8eB17aDYuzMptFj
ZbFzASqJ1nbpWeqtiS01Nh3RFy0vbebf0HCRGdSThSUKIhEqfJ/MT5PfItwO6Off
Ggz8auo1T7K9xnEnVzBTHj7qUjQmfeFoLp6nrT78f2ump6MAqYsCxO+Y63lB+1re
Y4Ne2hr7Vg0PT2joJw4cxPqAgpYpL1E0rukc4rJJYQ6UbPb8TIsAOFzQUW20ajpc
AGBMwfX+8ak1BlyVbwWpDxzDB9AC7ow1ABYF3Sxi6KLw4PMrliRPjAQAeeSOvzE9
Niwc8z7AqAHS8XccwsLAj2n2IDE830e+YMQ+zohKiokJJct1BW+LDkvnXh/nU57l
dCtisSLeZAC6JRVPRSoiaLCcXR4KlMg8+N4xSq4qO3PTpZc4SmMXZ0G0ZZ1LG3aF
yxeZIardcYqdvANQYX+MOicWKJiWQewfL6TcHWJe+Nlbc8wJGcGdclchTS1P9VtO
UzPIie7t9vyjkpwOOA1aVDDw20jmlZY086ShyZ7tRJxgiO+ovLmZzRPfkshSUOaN
Mr3xjbY2mR2t9EyOxxgmcnrUH/Z3fODyB1PBRPMvfuK9HAOMF3KrgfwDXfgYUDJc
Wu7JF5H2EDAygqgWDDf6C4B1ndmTh0JiqQdr1d+nbIURjv28llp1rawfpUqyaVFT
kjsfrSTQEt8PymXoez+Vtkd9kJR3/YqOcYxzRj+LBk2w7JJJAq1NaQDaNcU8Q3tr
ztlShFl0CoH4VpgDBdpfssSnxH6enosd5GMmSUCV9ZInZ8BF1y0eA08hXsydZGh1
xDbjy8mctfA1we678PMx27iTgoEFUqx28+ebV4OqGbLbkxoHe95ywDSmiHLBoL2P
mRuN78fnHua3smhOykyWNzBM/Xz38RtO5DInKqmiwTen2gjZIHGcoz9bTcYHPlQF
R6nysuFEnh2mbt2C8k6iP0u7Aa/QgdcizUpybSzLFwMKugO+hNrAbIXhrt7vJc+z
8oZ00KzzhBJModZaGW0f/qkn1+3UGSODoAxpgISk6ejhEiFH6leZcZwX1o1ppl7t
1KPmLX3xLuJ2cfFzYjFVKI/nnXLfMdsGL+63qGEwjrimygyi1kEqYgSo80QlTULP
SzcXRmnotL7/4WUHiSPupvTGXO1ih6tD9GlBB1Nk/pKsae9dE0l1Q11PbcVPmLXR
4HzACszPC2BH0QIMlMVWdTRFJzy65YzbZX9ARCUqs9PIwSnkDpL7Exp6pwT7UxZQ
ZDuuN66zkN5yR1XnvEZFE56upnxn5uWLyS0cInt4zAinSR+jEuHWFhfxiHo+bp1M
x+B4cVM8ZPSmB1Cp3oDUtk1Dk1iwd+GPs2cuh4y9skPWNnuejtMK9Ftl2n4djcN6
Q4YoxngYf0/i7K5f1xl7mghlSF5gObXQnnX0dxKnck1+LX+KnFfREjOIKr2Fxmi0
sWbuwPmkV94crHf4YmR1eYzyY1oNRT8ZEnD3OBgbMcj4gop8efo6BaoZblyTM/c2
XfYgG0zkw3+h7NXdSZPnOXXK3xn/u+wAGVGTIxE2rsgxqplrlxFCsbBtNd3/f6dh
rawea1mtwH9WqGYNWwjEzWaGKTZgkBzuwtqm77axrHFkVsVbjdwja9OnfsBVQD3J
FuCyBa+85W8T0r1sfyjQpfap+VJOsGnVUYgnNe1UFMZs5eGszw9YUwW4FWmmswlk
9VeMP0E9tjcZ2BG3fpq6wQwUjMOtnFsN+10kNVlg6vwHhZXdQXdEQ9zf0nF3mTmo
PqrXML5LwM+EJSqNbLoOmbmWK8CheWFAqP9HPCofLSLOyXZ04OglCPK4CQRFaNBn
WN6rzX0d33+x57qeqMLA5oBqMgtUtrZ52Ud5PLCyFMSy/BN5jEHPN9do2c5k0ZP7
6MWLMKZb39RwE+d4i/J3lEjuNZrVgDBp7gAkOc9UZe9VoR8q+z38JHA2BZNdTV6U
dtCZ1a9QupfA1YG6Cfsx0LhhyBP0GtAVx8/27RiKf6jvWJ3MQzZ2b8C40wpxFHfX
Cp27zwWWud8rruFZaLZE17sjOU8Jrk6uGIflD/98T+IL25KkSws27XAxDPhX81nR
TDLs1J6CLL/okiU7SG1QU0DtBZS0dAynIHBoZ/Vy1SXwFau9Nhep0EE/NXTMUvOL
Re65k2R8f963gvtA12PjIpOFQPGZLNTeX8MAPuvssbgrNRf+1fn4vDZjR1jLPAqZ
VQupc8XaHApFUB6NQBgcSRfQssBIPrFwv99JvuZJ5DVpALriWWAq9y1Sg96LGoOg
0189yxVnFZT94frQOD8rP+DPAddcOGsvE8vpzRqi0NOcdwmSTmYnRwKpbJiqv8qb
HCaH9/EgU4oR43zDEmBXCGT+Cfg2/siiy3fj52bJwDXDzAfxxhXg4n88OkUu4Oct
IMoMV7YIVvoMoWXKhBjWp+SFXOyU6XA+4C1/7c781EXcXPytR9M5EaYIlgEUFYl7
tPeI6NDZybBb5mnGcelrTpYLfSL5J/ozX0DoeVZyYpl6uW25M0kQbMl/HYwtST/5
toLoo9XUn8D7VFWHkQyriv79tq8Qhb4CxUdmz2MjKjbmb8exvcQzb3oToLpiKnjn
oKoYtU5jYcdUvV4ky8c87qRfTYpyHQQRp3Ul4AEdMy49GAtA/Nkwq49MKbOE3fis
cNaQVVMZTH1hgHH6jLnNtgfxZJECFNsWs7KEVAfEJpwWX7utydaY/HPiS0o83Euh
nVYPpCJiV2lNJ/VuiqEDd/ij1GmGLPbVTpE/6rhTpdXKZAysUqw1LpLs//JAH16d
R0fpnx1myKiNOpbN8+WMPWtHtqlwiVJ2I0WQ68Z3Ox8bzNGB32U19VlrDb7bqbP0
Uwlpe9m2gmG6lJsV6BbdJRVSJs5ccmC4nGLDlgKXkeEoGb6IK0n+fsqFmQxE0SPC
Lf0cILJFXmjizw3zXLxVQLVwFIcoURPXxUt7C0nnAb7BUpfMr/wgTsI+AmefWjHL
/warkYV/WGg6FGfhl8jXsO0HVRiOInVQuIS302UZNRfx49jWuDyAY08K0rhF5ApA
X9cG/KJD80uTWCKRrTyGytB323jTrVlbtPgSSu4CzjYj8YDSLN5Xbq/7QFPtaTkj
1M+ZRjtgNJ01lWHB/UllPuhA0MhmFadDWBlOt0ouEchCL6r7nhNdk3h+EP17LGX9
NYYsmyciTGFiwOgaWb51maBPTY8RsWMMzmXJrrx1aiPiYmPBouZCozrNufnpKMw9
6zATz/G2q57HYZUA9Y+wsANo5HTrYwcEoIOEjP2HoW3jJz+4/hFgZdKH7GGg0Uz+
t84PaG9X51hDpn7nWD5ZLwPnR0rOFmiahUZNIln9ehDkIyWxn+oIHBrZO4wfJZCQ
mbRLPv7ex/3Koma+jOe4t+jn1vvaJZC/5XygaAUhf14SsAyum3bIjFh38nn5dKrC
achpTGFgOA1mRoxFLPENfzfsauC2Z8fWSC+9iUxopE2aFZDhQ4kdfl/0NJ8eXZmJ
fakQeogP1E0J5R5MOMYhDVX2mvWPpy96RfzeNwdx8xiguStGMrrvAu7MlD/4eGyR
ejEwqnOl3YUphCXIiXZ5RWHA+jdihdv7HkUs9dJeI8Wa6OrJ+t+eXopLzqjzplBn
IYBm4xBlKTZsutJ1ie2fWalrxLxtH5fKItalAfH26ns1WeYuYLLdz1A8QNHs9Atx
0Hoq59Zy7Cr4RmnXEbm/ow9QPnFRG9WboSH8bqjlUU0l9UYijdBYqfaD9Y4cPi6j
lZ7vfmAIo9isVKRfJ2bnFMxC0odnluOZGBc+ZfW573coQuXF2Z00qUH3DAbnMF0Q
lTyMSTLvvtuw7Q32J9p822ea3LSOsKJxd+nb4QCxLpJ0jWReP9c60J/1U9hF3Zz4
Yo2kDN+4eKYgla0aScWa6+mEQpBz9kVuEKJCnLbFya1L1UkBqIbr0xYld853f90K
T3OnhQ3rS/pdrhfTYJXXgem9h1wJeEk2OMZh3Uv4pv7zuijyjFWjF1wB/yrJv/nt
70/r1upAdv07u+M6HMPYt7EKeTPyp2F+RxlgnSjGXwhurf6BGKwRZ/cIkfdxsDvG
Y65/rG6wCscDlmMXn84z1NEuH/47nTVvZCNlAC1jD6fnqD1+ov1CfOfVFCFnnihB
Yt+QaF+XiOQKCZ+JaOoLkEazAaYedMHmXzqRC3PH7BqHQUj4HiTNlctzt0T4CZsM
dTgLaa9Z+qd1peU7GyG6yt7Qrc49150ANmCdOVCtSa2Hqw9srbIGDH8HeyB3frNt
4Z+nfBQL1MUxnidr2OB0qxysfsHzxxg8wNa0ASrzADZEHmPzQwWuBJgAnBy1qNsj
jLeOrbB3oNm6jo+BttMwMdJuLHA288pOM51dOP3M+k/rDMiFwqi6/a5cNVuVV98x
iPWY3xpriNfUhDjwUq4zfprrEyCdROaBokdtxJPVaV199F5KIW9V3Lnv2c2g4Ilm
2ZHMjf2Z/9oA+aV67d9xomxsSzJ75kXWVWBxN4Gp69ueZTOLAqiEgARhQCTHd8Pj
pCkRqcoMyF9ig9aNqgWnH2Wy4cI1wI1JjWHhH+S8y3tYDBleC2SXqzrdFKqffjqT
5lhJH0PkkarSEqix0OD8+ND9jB6FXrRKJ3m/svnpcKRp1mHRJC5UKnpWfxrqxiqa
evhx01WEFNXbvlbB6WH+azzJXuThE1usRNKEegQMYzZ9PGc/0dfbhJg+S2CP4QG2
bvV/64xUq9lNC/5qIBEn0d2R1yAq12F8wPATanOTlGGF4oqqEwlry2WMer/OpBJU
9eH+NrQ6pea/YfWFU6LiqjvEbUpR7kqV/6gw8HgpINl+sK5zJQtTavspJte3COG4
nhLTYUUq4Aqfa5IQV0FuEjTmaPcdSOQ5+3xLjVGxsoMlgZG5/z2mRDTzA97ThnaG
5VG069aXix/4Ju8OrGp+L3YBj/lW2N0gUvpGtB/iDSr0XntaLglzT3f4MIl1UC+t
XP5Y/JFJAjj5FH0Dl4mN+N1ZOsN+IDwpEOG7Jdzf/3aFno4LdYfTXnUEMdzkuKO1
9YcddnaFAHCwmA3bKBPF6NGkhUCDWvcc9nCdMZ2xLivVMkhmeIcdcA939hCmWz2N
STj236BbAbyAUCz00OJBB9sKrQa7k+X66PcWaB+M3zCE+mKXSKqI0J0ZoPeliW7c
brFX7MfVCVQExjKnOqaGJqn3Xdo3+8YY/I4tL81zJ3wGSADruqYDqIxBnMwkODBE
V8UOkUD5RLQVSsYWZMFpsrLq3PpG5czbqmSBTiLD9/hI6fIEI2NfonSFO3vrx0tb
22kRNP14pIyGaoGO4rWIErRGlZ8PGjUg5sOyG0wws75oVm41b0hOzxAc2nJDS02Y
CA+8u26ce/dTfP8G7QmN0WJ8x24CGH+0HlP/r7QNB98Et7xS/sWH47/Sz5rjPiN5
M7sZYpzXnACnMTsKP/OleNkSzr+wbOI6mcRYr2+CGjH1f0M97q8RL06O60FHS78N
dUnyFZR2mPU4Xur804rXoWKh2IYYeGYQ//55D+23qyEQPJnCKYga/A+MtaFEd7eN
cjcy0+2ToOAqElpKsuiduD6joNWkU1psfFrhM9SzEobyRDFlhbqEsNMtdEOdCbAX
YrkFcFnaHg5OHhfW6exnFVr2IdeDsazvkLYkvOAghdplviL1gCvwbdQNtCvMca/h
U5ZfEvbJhjemCs6wva65EWrIzQ7uupHaFePNMr9u8pNALgGlBtvZdENd7Y0qDE61
YdEwuSUa9WonHtCb/UemSAIAwiwFitq3RGsOX7aKWe06DyG30CqnlfxyhcThkQ+x
eWVA68DfljXxq/LWi25uWJFjpxYuKmP/uXxXeFQlcopceEm1TsVY98GTlnxBuCZk
F6jApA7UtIJacFVnORosskNdDR6XMPOfa9AKbfglnDA87eKEgplLoHG5luQY5BJG
jbu51BtG5yc/VhHUtBpKl75BQ8BmlP88jSaDOVYwpmRxn038zFq9tW6JuE9TmA9B
aVQ6EopBo3hF11nIuA1cthRpZapgU4zvwIL5TkNILcC3JYBPqp9peHlEafKte3E/
8856KI5LgqFgi+31N3iWgjDgBG5axR6Nxv1CFzS2ruDRucVnNL2Aq4+xPS4+KR28
pmQcy7E6fLErbz4W4mK6dHV7+p73GO9eaj/X1JBSO2bSkhkiLrO69Qkdvt8KtEHf
av8NkEKeEYUdcN9A/+dbLmpLcI0Vmm/HYi6vQOhBG9gZNljI2lGqjY2HGjXV5jHo
aLDopB+vvNjod61n2bF+i3RTAF9VV5ZJFoS5ig5uIFs1VXgSQ9EsQo+RUB+a7urN
G7DQWZ7TiMCk2CvwZRBEunJt7M6UHvRz4segajRuyzOpJBzvVX5WMooxaImgt8Ng
ftvrcelyXOuaofFH446ooC+IxJ5pRD9hk/VBBL+F+9stf2YvGEpRW0F7R2AqWWVW
485MGY0se5qlAPJy43n2ToPbbjtMm/sVSgHgM5t8rxlu3OGE1W5JoJzldeCDyfcD
2i/j2/IHg3LML9nLOlkYbofWtwQq88dTOVfxR5MfqbbNieckpWVqZZ7O6Kj8A+pF
Wdo91oT8LKEGKHtEPrlpXfRuNXuDUYqbQqyuA55MWMCp4xd86YZNiHp5DsHKrdFN
n9pw2z7YnQ04r2zapv3RMWnVUzgRjExAtqwzAGdNIQDrcioxzBwCA01kKi/zGuvL
laV4mq69eLgQGRo49nxNByx+WclGxQbJHfEODLEICqlfSbpa5Zp3MLQBMnuuPESE
5NCRUNMvcF/Sj8uBsFTdwbQ8dPWWB3PpqIQUN73uYgXiRx1tZU14EMsm9YT1O7qm
VHiGSlAgQEDgrJnfYQMi4USVCzziqXcEIkmfvjtPeOcPWAtQSAJzt250Rcmcw4Tv
oBArhZiVDSPaUMSTeok7l/B9K23PeIV64TwAtxkh5Gr2ySJM+Ckqe7iB/cYJsWF9
RIf2sF/+fWkNsUKlpLwhOpFT8fyxXT8z5iYSoULODSXV3oOvjXAgMX1QFgbyEEcP
0x5QfAxoJXSv4X+sK31bZnfZdKj63MYav0SstgkaM3M+P83JhtpE3w9VLA55Swjq
u4Kp/MML4to2THBlPOUmF+0N+I+N+onjYlNNib7D1lrSU3gN7VDAhND8pLP5l8L2
tD/0iN/6/kfluPzKNWXp65Ji5zgsg4MFPGJWs9qbBG6C1E+JH0Y8PvALfCVedba+
rNFwOp0gVo2xpx7Cb1J1AWiDMNuBXMe5veVxBeFKgQnkLAxllZAhU9HHehBBlBc9
zX8OHR9NRJJ+wl0n2xPLcm9m2e11rB/UaHRZXuqU5laV9JXQFgXa7vTKMPMKgIJd
vFdwW8nA4qar9Hh6nFR6B3WhZ2hAYeoaMzzMth31OlFBKj1mRKshoojMfoqJ+bCr
6OCVibjfMIMq1FVd5m4uhZbQnhf90mqk+mJVj7+84e4hJ2AXkfmONvo7KXDsKshq
GO3nzYkGQzgn1KxLo5wHFi0mBRv4Ium5FHnVENA+Gonk2aiZUoX16eDp4ILWWtH9
gvnV5fqExLrl1E73c4jHQwNkAgDrQK3OE1fcTkaD9ewYiJ1X6yPjt0Kl38rhin4u
r79hIqQaHZJPDIxOKsKPZIlhcLjk1SrOAJa9IGw19kQ5EW4801summlaUcwixoLf
P+y1a8X1PQWcwG/46snkveZHN0z+q3C/pbOmEP2nDMBQfLT47KJHIUmXls+x2RbO
+NhYHuXaTP5fDyPYthMk+Liyf772sEGIQ8D4tZMJ/VFs+u/QlSK6+kY06qTl2mps
HW/mgAQo8Xeablq8e9AFY/4KCr6FIOTaqtsqyQ7NMxIzv7Xzbj7KUKi8KSdBlXpy
sMQgedx6eyYc4mt7HwR6xmOqzIk7+YJjBd8ekCE1Xpq18ejpA2XzKK8qGyPjS1j5
QmyiRqB8fZbncuMKWYTXorXcYQwEjpoF8Lb30FkjEsY4+Ip14AnYzOZgs1kzaSS3
y8Lz9X3OuSuaJU4qX13qtLVNbMA6RoVwgJt+vsUcbMGIaA4BepT6qYeT7LDMDCms
Sk4G9JeoquhQbXCRPalNVNLiPKurwy+6dFaBEiZEngjPN5OO0xrleAwFiNRwIFGh
W7Jx4DTnH4LjocKWxd/tdAKUf1Xy4OoZ+d6eX9HPsV6zthn+LKItgskG8IV4RnOE
crtnWuyGlSessJV2SaEB+xvmLRX1ysdFS1BdiZh9WXW0iKmHa651S1woDEccilb/
WSWuF54aqq+GU8klYJ0splZoy9nMefv1AHiT5t5nN18MqUM8RTSUPgwgnO/AxsGv
KmH8Gy2efsmuhhizKYpoZrO6Tp0FLDy4w7Tl2VbLQrRPzevA+cxtwYrkB+ap64XH
KcX3QpqjIlnXoiWrb8Q7ZTwhr3/4oTNURR4a+1y+Wn1vt0vOApNy5MJPqtYBP512
jQ20SZqLYq3lVoCzqOKeC5OfwGIUy3o2JmgXUoTuyMUlfl7hApKicuXSekxBl7SH
o6YZ6e4kpSrrf6uY/mgoXBH7ZtzqBYMJjAlcqGVSk5Gp+gWIw0Oielqka87hXW4i
i3TIkQML+HoZhn1PVpdrbWG5TTWST4fgNwvYDtnwm9/90/OotllDJS8UEfTR/GvQ
QpCPHzUNtDGAi13iB+bJRMVjGhZvuxGLRFxSOKeERI6DmAU2SIbC+W3zpjXdLwpB
yDtJvmnWjCHXdg9DaDqq5wLUjO8/zKSbXTVhcTHE0XU9IYwI8FT4KNFdFfaXreU6
mWlGde0v3s48WZz7Ub2YssSldixpfHN/IbehyClKrW5OediBVFAQGTMhoM34e12+
XSad4OfVz+6WHzFX9adoeH2YKEL7VVRA26ZQXgGJOjI6Tjicshp/3F0bwAkiPmOT
6imRYUw3jOC7jCQ/iwz8aGD9koi8UkVfFKR6mUniuTkrztOrzeKvKw2erSuaTIrU
i0dN9CJV8gW+5CrSha0VFIhGZvql1WStugLasHYcRF3kmnbseJXR02p2oKu8MO1F
xQrOFD9F7qeCWQ2zUrxIRjMmyeIUjnvUvzWyllR5ASQRv1HKcqzde21hILygOZco
xXsyEgG2MNXXvYgTUxVh/3pEsigAltzaWDGAkyulpRKl0mhB3wP8f2iMLQOfkBOC
EITFvUbX8iA+agwnqClYQnl97oS41S5+oh+HFUHqk8PdpC3Sb0BGSLwCXPTuooW7
at8wDeW6CQLI7bPsy78scos1dDNlESmieaZw8pfmaphi8zJ3L4dXmCC3t1Fo5b4N
0F9smVHmyQDLUrLFWSAPDBT2d+kriO6yp0GYOudJlLKyPxTyGxVDyIFcBDZO+v28
z06OoVN04zJLO3OMJvAyORk0tmny/mO8OGNr50Uqyf0etiBoAUj95T3YYnBlw/uJ
iLY8iBtAj6cqIAxwQ+MZrKQHfuvGLx2NHFoZDgGmON1c41IEpJmgTWAEMqchg7uc
v7IwErLo3zUBpDxBiAcoXIzaKsvYn8ZvT1dbVnynfDns/7EQ0EnQgogRkyafdLwN
2ajzLtWqdgUnuGJh6Z4hVje58Ca8ZYzRNC0n2R7DNSE45jNBDhDgC+qXId0jc7Qo
Gfp86W4n1y8u3Kw/j1g73yrfAQDc++4zaypsCd1enBhWUpeo9MsJB+nDlgy6el1l
Q2lF5kNug0jwZE9sV6r+KUKjqkrUw2WD7SNL0MMXGTcDa6rB72NVzDrJk8/4WynZ
tRVyxalqOF1G9dJciemqWyZvrGekwq/6qVcdUESEqEFl0IUosRjkwQQjSr2GImtv
njpcHulwwNLyTifNPIfB2m15wDbB3xnvj85CdjWBiQweaZKDVIfF95sDujZimLoW
D3g4kx9NcQ7nMEYGbs0OvQ/82gSOkUEqYi2q/RJDjIMmQGV0QEW1NnZ9Z/GUZdfW
KMnJlZ2M0XU5I29JgK8q4aaEJaf02IX/kvom+B1SdMuO1XZwiTZeK8Bo5FIaDnIg
mTToZOT1m/Rp2gifkwEg8XspDLVRo8U2k3YVxOLFkiXQyf0jiMZxm6If+vI38Nsj
tGLlOuGYQur2kS0rW88LKiCypgiB7MhT6kQGbexpuVkvpN3JNwP9aY5OhxjVpvxx
FUB1B3svhuWOxIiMtX2fnhncEwYfXVw9KOEHzszQZEwA1w9nCmR6dKEyp0XBq6CK
nlRmuf9IyjYymT6LBvxqpZQruA/upO9mAh9c08rnfV9kKEX3rTA01zea1JWjMKm1
kbMyTGL2fCllJoyev5kKj6PqYnFWUEBU1iVMnfWxJS9SLxh1To0yGZcJamvh0Vyo
62hOJ2U1s2a0b6SL5JpvMMunbqgLSHFzyb1lUHEbsLayhYNBrU6N0ezKcmqJ2aVk
avYlVDyu11RtHhHIJx5be3tm/Aw3n3/lDwp7J21GUh7vwZ79+RbgimtL74Va/Bk8
GmIB5UD9LIHsCqsflufgwq76Nj7NEwysgByhJcYBlgKBBBPdQJoh6XUyCdpqb8IZ
Z1nUbUknCHWaOA5vgIjqm0vh8rcm3QrowimmsvxB7pFrwVIrqR2KUOio+35vyzxn
5XAxlGubuU8YXd7Ub3ThmKlTkaQa914QH7O9dwp0rps+hamvh0nLo23EJzIunScQ
17/0f50ipGSDZDuukO+6g8iPMGcFri5T85iPSJ6iRv4r3vXoWAfOJrF0pSVIMSGm
8MI4raqwSdgZ9S0y4RT8kTTTSaoZzwY2ram51ynyozcj6Gi3VkVPKv7GLqmele6n
MjfKpGo2jWNw/GTn01rIZYf7Q7lOOmJDbivoZJxO7f5pCXKq69BaIg4ickwKnSx1
1DVjQ2zCOezXOCAno/9a2W8O/ejZD8pP1u/ETMFNJWO6PWbDr1TepW+9J/4W4ckr
iUju0WGpfYodG+ARZb61ai4nWOftiXnn6i20R2YjpQmbd5VR7WULqkkFtvYVYRrb
Q8kGX5WwQF1qzH3eLbH6LvwlZXKnayCPBCoSA+cQ0CKqWWvMOOsy22eXhMPj+m2X
m6/x4I5Ekp29JHDy7TLpAYXbgIbOfPlqsHK6+Z4cnh8EHWGd+NXISB0VkJ3G7Zo3
JxFoO9S1owTz7JO+yLOPRz9eL95q/BLVAAYNEbQYofWefpwW9rbyLPN4Cijdqzcw
a43E874LJJPQXQNaCEjw5f15adC9CejmCuwkK6gIpcVmXx1cxVUFbiyZ6eJb9gmE
XIxbr03834hFS8A2/T52cAn3lcHT1UphJlJNSOOyxNNfPGowEHIS2FSXlsOsj+Hg
x0GD1V3Xo0AUSxYmQBftCZcIWBGRab5e7j/1lhkgZUBTacIMwT4dtMV3Y1jonUtk
op2cz/s2azR46VUjPM2JHbOzqMWiuIzBvWJYfeEibpA6iKbOJuVM4QD5nzN5AohL
XZSm0Th4J7289NG4xJGHEDYiGg7ZMIs+KVQqH4IrIaR+oxzP/rkVlMsyK+eaT9rK
H7rsViabgkD1b/X9o2dMOG2Pctz5QJQaIE3i2/DsumBL/lK+B70TVcPuMox3CCpl
Feb7A25muGchPHiGnSDJ/QsjPZofWIh2HEVwqTCLv6sFv93CLps7zAkdIvKWs9MH
DcHkr6QgoyZQguWeG+ru1tnihcy0zCGmjsDwfkFdgv2o5qozHRgpb+SN9+ePu9va
VsRNfMrTSRurEEoYwIMaUd+IHb/+jtom4disy4zfGYK1kzt8Oz1/Jtg/axjrgbSP
B/S/reFWT0WaH40O3BVVhHGX9Ik9V5Gibk/YOGfLqt4+9Lm+Te4UgH86x5fenNrh
1S4OfYznk5SbvAsJCcX65A37DjEMb2StDXWn8dDQY9f8iTZumDaKMMGJRb1U0HvK
s09tODfs0zz6cyB/DSl6NvH6VtSn2Kw/mKGCyC3ewb8PD/Z8y/qqTNOpmwUyoimU
gxsblxzt8VIBXSAqSMsor7SJPBt8Cz1RnILbYVFMb47IwGjF35SNkdE8iL39grSE
WKxPc0qo3uFGv+SE2iu+A2xT+M/Qew1TKf0VKaiCiQjvDMu0U8GvvbIFMhDyG2xi
/OrgZ1qL+g8kIXgis5pBm63WH/fIjgAisB3RhxalU8T0udCSHwBGD/D5Hj08RM+x
tJbhk5lVskcDCh3TTvXQ8HfCeXiJHT3gVeRh2VMV6PRI3Y2wIvNsgpJE3DHIYybU
QqVYx6Kd/pL5r1BRQR1TlgbFdHFQ6QuwoobBFydJe3gnLwGgrav/76OCIQfFEh3q
h8nQuZobT2CE2j1h9L55CKoyKZOAP/bQJzzeeWYSYMro5qab3g90K4PjX2v90+di
iZhsZVMrcJGF3h+iq/X/2syG8dvxF0L7QH24rb6EMRvTONy6dt5LHse8eX8qdU2d
+jJrABq+tfcYdI31xpMvCjFRfrTCwfbN2bfwqarJCJBCG5sFWjsOvgGVUGQcbq6U
qLQf2K48sHO5SouOfWRBCUMx8sxAQbYbB7j/S05f4ICcrm+0fRK5xxZWTtAtJ8hv
3HsgbAfEw1eSYQd/0/HS9DcCVQSX2YS2HxrOdvV1WrbYgznGR4UAfSBU5D5qAaFZ
K4qt0kne/60md3cGEEcxHcKSpKb9wvKaAQAeeRciGlqkkP8i9o9y3mI7/pZjtHJK
W14PatzjQCa1qA40EAS0zXUhGxXRnkGLfW4Tqq5T0rT/PrO3YNlbwGB7VOCzywGY
EDIuYx9lw5JPlVoQCAywwhBuihQGt2PSQsaqwXkXq7TMMkdJ9b32szsKv+ZX9aeJ
GstoTj1WS39awl0VgC61DMbObmmCVsGxKcMt5RBLgxqdcACJvAtPeiR+Nd5SUQHR
AIPYKmIS9XyYYJOy0KA76GacvTLvb6PkHuZh7gEpakzNKKA1MyKYgmA6Bt8qLOqX
D8Ae3PYWcJ7SIsgR5B6t3TgF1d4NUoXqSmIjUsT6MpZUiyn6R8b6wNTPikvq51HH
QtrjJllGZXsA+cJ9tfRI2JGARu7eYBzn9VRoqXM+FE8VG5pf4oJmTUvf+0UHpWzT
C5Zx+cYtGiu88jncMAn784qXUM/XsgMOg42CbuGOjCvEAQuMmYmStzPnB04/p+ar
iGS/7f79rdUorZBq/o6eGvu/e8mnrssajIQWI5t26zadDey8oxatNW9snQWRo5bh
RtNXCj1SqeT49FU/AY7uCkJD2+jYZ6cxHEsa2tA3tE8ISl/x6kM80Oe1hqR+Dy8p
RLrbGK2kzGQ0XraVfaH0IQh3HHf7ko7sTVx1ksd1x+SBrTz6q4NEVoBBLc+cWKT/
zMwzKO7+FXkGtU5DyDHgXOzLIyQ+0f2iWxItIe97n27p+7LmOtoqk0iYdjINo8R/
WMmCCX3eWdbXslpB1uNA7AiPXQZWfd0Q5VFpIqSxD08Pm2GMeWXJ4Z2gNdHWVCwp
pCwPRA4uF1ekYAa7JYlmDe9YsvOcpMnDAFA3tZCD0rC/oAo64ThXexRgxRa9jvOi
UezNc8qOD309w6y9p/EY9CI0IogWCj1wZBRXrvqTYb1FwoNMqv8QoYwz3Yn541vl
52P/PUO9B9z9LA06q8E8jueT4GSdBGBIcgW8cuuiaAh+H6i2A/WQSH2fR68k9fhh
vtd/gxmp09NT/kEPhrfbEKer/pqe+D6gnmE+YOrp1AJSjawHWj2kRrfbslpx4kQi
yNBncfwWRfvVmn90TVpAgifFLUUX6ByTre2jputoHLZJrXjW/bMXlOeinU/aHUQp
duEOgv79FIJQ/m40vKW3dJ8lDHK4oKbQD5CuosooYY62GHFfuMbarN7vrIs7r8jW
Gz0J8rthW18RI+72bPLdTBiNPwIXAFv/u8o3ZEpD9aXJ1iCP23ISaZcqNOJ3KfDz
ZOFsANnlFHDKDed9lVHsJG0HiZMEmo4YVP4+v3nZLsZ6eUqDuK5OufyyO0J8EsJ2
6fKzaRUUUVZrd9g1whjxaHXR4vg2B5tOn4l2ESX1Z/KkRLbjRyrDkO+tvYw3+X2y
4YiA0WU+XI6zis4Lw9f44bXSfWPTLAFS/Fk2fmCXfslpWA9DeZpKiKQm3njeZi4p
QNiqQIN6dfPDc6qVMblvHEVrRgOFh5eCQ7KAvzHkxt83mMdEVwZ0U4Q/752Vf+2N
eKWIyAN++j8drq4CGZ2rTSR8Lyh5Naqj5hjzmiVY81wKyU8lo3DkvDWpBBZInq0Q
zCTpTY3PdCee6zcWCws0q4FUUGHwaGJt2SEi5SiUcCKNbal3jYjqqw0qaVEfNOit
Y6rON1fEQL93YEg5IXKQwsObGI/fefVSopJP48wuYO9r9uaKsGBpuOpZH7rn/cbQ
fDfFnKiLuCUPRqmoxtgajFnDS5T4EtyaN9zfS4voHQMB16bHeYSeqJGemjbLRZoP
VM7L7Pb2g+/JGjmfQ6af7DPHOHH0YPlNOGaPI8OMOwnqIweDhTlM0a8X65CreZFH
HVAPS4Y8oW0S+FTUHEXDTDTfOY5ThgkESSoLqa6nWeeObpkYSGj0hk+xUhMK1fzY
eLOXTno0maS3GvBtFNrSaydu1gMhjgrY55aDeihsUIBXF9BWtIYJuYK+nilCEwDj
j9v0UOr1phLZO8oXbBpSGAAo0vFnQeIPA78m8eff0XJFk86Go7QAR5DxKKMX1BuA
jC39MDTV7g/QMeIJSksmOP3LS6NeSSGKbrpofs+HjbecMo1QCyD9FuhrUI/tIcC/
uVRf/Vgl1YZeTn8JSp44YLe6AKtqZkAQdSNU/hSMf4TZJ69MeeQRvrL5b/xL8tMn
TazqWsmTCMELPboyMpkCpwD1dA1SurHSCHTfpecutvhY6Drw5MCuEBLK5GjluTqO
4dZMXHPnTSCcjuEwc8HWhuhckY5oCa0YJmwTjBB5y/fQ2eCL3iNHlrOORD/jZa9T
U0JE2fqAeInVps16ViGxRHhKrjVlOZE5XDBGodTI+kBJItvD7ACvpNLtqHx7urK2
3qKBgG6BxmXecrOEwgEovSIkfRCKgSb6JFz1HfJcXEmhjQ6CEpbwrkH5dMNbLU41
OYJ53bLLigUIbv4K6+4dINHn6ZxBmkwHfWYBYSp4DV8e1G3de+JmZPr3RymN3Ipy
/eUsV2HLIUyw9WigFbH0JtmS+JF+0Ga2gcNa05yddQc7H2S6msVViWyyX2NN15oe
i6otmG38aopdDADgGjITnbkq6UaccX5Ojc9hWnDF23TuV+x5uW3Ii5wsYDMTSXQM
9IqK39dttcwLHuRWLN2XPOUXgGuqb052VVnVGjikDAGgP/AE8BrX8Hj45sDG4QFK
5uaMtFvjbjWTYwL/AAVkbWnEfyHpoGny4YNH+sfkKINtzeS3PerQ3BdkUt6oXM39
J0AjdDFHoPlj0jEeH+Hzorrxa2LQ6Duh803xvQn0RFo6n2vZsXrHO6MFz3wqQ2ry
3qHgVpxG+dPEDMMVI7vfyJXCdnRJYFSjnsPmvTl9N6PHncwDQtpQo6V2Ron8E8d1
feCPM0wEWzVi/Wl3lQ47QG3IKyT0iMchdzEu7evKZhvmPEFOhCFYfkPYndHtS7PL
YdP0Yha4QXtOtAVskWkqcFDPKZmmKvx7B31Uou+ty1jpem1HZvKx82KxIBtt5Nzk
ZRpDOhlqPCCf4W0pCXEs5Qj7x3DG5V11u8js5Am12uvloqmFdI3qYCb8d3+Vnww/
L5gM1GOtqkXLZ00zGirM4KnTrYR3lykZesjmAgW4tU8obgy3XZlM07JCFLtWXTRB
ulH3sTmgT9MzP3XQPpBchubNAItgwahCaA8KBBHwTQ9fIxNKpSRc71tpiXA7HDAC
xUxNSVu33Zv9lvSZ5+Z8KA5A9TFks3ccom9a+aJidWO+Owo7aXWx32aEaPv3LhlH
9GS2blNU5R2i90ZKfTrQ1VqBOQD67iu01VJI9503lNZ7AlvO/0Apj80C70ocrt4n
pQSIh9iLaLbn6+frTR+i/QsTgFjvS2Sjn74LFQNnbZtAXdM/Xxkt/CaVt1TgKldg
Ji/sQZesaEtS3WWhz8GO9g+lR3sqPgLtAHIbPybDtIQQwT8NKt0E7RGD52PyKjMU
Ofn8G/v1YVRsh4vjPDdiHwyeVlUEzSQQp9XzffA76KQwSjuvaRnrKmZnkIk90qkM
RJD1TWZ5TuSBfi4bEtdyg1vEMyqp2whwbR2jzctgqecsjyD/k0V6vOy8de9sdbya
EWCoHW9uHPooN6mvyqlDsZHQ4J5xolCXh5wV4TwBbxs3gftopoTY7hmJ0eCwLeCl
nlk4rAbeU/FuKSUpSdc9KO2LI7KoO2llwNZ1GZkLDPNLCk4YPX6R3Yh0rBcQqZ+b
46GMeMF+WM+JBG2uj6As3NLj1OIinKoNWFAIybrEhrwBvIGKTfXh/ZhSLD24yplK
aUeKNZJWVu7XXLKsnnArVJOsJuhjRMCb6YaZ1j0FkQAvsq7rnIr5R35MAfKY4+aw
PEEj2PiQsc6BtG7AB7VVSbumNiwAIU9vjJyuyF01I481CkMZjkbxx0tfTD0cnhL3
iLV4iK3ZFHqWpurBIsi4NK9V5Jb3Kkv51ni7E9b4q6OtxWMiqBiTzmiF1kcxSF3b
Aixrgl/ejkqlioTVf3OYa3XuIL1b0PPDOTYOlTVvOeTkgolfqU7/XmeHpjLIAhzm
CPxzgwbUizLsKQYHZF9V6FwOuGJvd18jHkkCqjerfuG3VAfKDxsAzidwHxEpZ9eg
E4k+HfeM2gLOxp4DZBBr5md6pFv6oLIjzXOfRgBaCVAzXaU2i9DnP0I1pIYPjizY
jXB7kvTGGTZXxNpQnvdyeT3GMCzQxi3P6AJWP8ydWttdASzf8/sYpcvHo9OnGdBS
B/aNZrG78/fe0Kpwmjq1vUauvZg+8vyt8L3bry9c/I1o//OTNFU5BPRlxXbrxUH4
5EWT4lYYfDurCG+S2vHMP1nzvcDzM6rzBqcKl6kS00ALiFT2dsx2gN+grXT3srPO
TKjte3udY/lSHwNtKEw9LHSLkGzhn2RWer4BYYR4zKd9E5drDyf2MvtFmVmIeuQO
cqSlyCJ0zoA5zGT+w8k+yO9+g0pTdeXJlpDksczWMTW3JW+JPfLtONkEsTPM3xyJ
mTPwqREyAfrGJ2JcCYhWbCpNhRmVIWV2sKDBdbHYOmnSMAOSmTgWpAgZtX9QIZqM
Zf4k+A2KNvtulqJC2oRqhYs6mLlz4kfAjrm8aCn3bfIg4Rd3lUmCINSU6/y2r9U1
8sHg3GuotYLF+9B0zVIHzQwg7k/X+/rVbk9f1zDKhRHJT/d4fSyV7A0EbW3JFEJi
/xZ8nskdBOkKNtxvFtLqe2uAEFH9OonT5G1eMkNS5IsFtq22s//UrF9HmWB3avKL
Hd36EZMlKMB/8XKbyOXPkZPyCXhZgrJDJYp07BjnFc9k9H/6FmEfIOv1Wn/8s7uz
jXU9WF9cHBQIY7S7x/0W3s7YHiluccvE3fna6fPjgkL5Ajfk73OLkSawX9cY07of
SLrBd6GQ4BI+YKgdCt7oQfqOWwxKNw+StPglvHGx7sh/ZNbQW6ZytGj2gwW8WTNZ
JYs1Kh8hEzBN0xmkjgburn3HwkJaXjDdiW1X5oLEMORckXpglHRMyAc8yhrsVzpk
cnOQXmQ2zsxw8ksFQt6ziC+q+K2Mm0He+Yi8W1DiW81fKsFvPam+Mqx8uCMdgrhm
Y4XZAIlQDHbvpOhzPBInfhE4hH7BXkRvvUylTijL3QlE13FL7f4T61/pRfoeTe6M
ctrw0LtbVNv89WZZ3kz4YKEHTWHfcDhr2Ook6ml0XEBZeGr0UDdc7K967HwDPGyj
8G9/2xWMYpiT0/xvqFvx93NrzEhm3+OSNLLKZdO9kIzeABN1qrcvjfDpkE2HFQJR
UzyZl0koThzKAlXUkhJXKis3YGUdrOZ/fslNz7L3vTX00Ua/3Wz+6YpwmLY1ggSa
oQ9IF+Krb2yFt1N+QFnlC4asUARe0VatSPkPYM40NGnFfpaySmIfjNbiZTayQK7y
fWqp8AZ+iGxDEpWhssMO8irEea49Y12XyhFY4I/uCv9NRFXwa8B452ATIwR+2rcJ
wLywqx4tpTxQw71elmP6e0JcRmjC+m/kZA6vgvhQYMD6v3LvRzzXf2c+8xD5KXEg
4+Wlc0Vf7Cibi8HyfUko6IVyjInXQ4Wd4Vs5AVSNTFyKM5SaoUy4VUOl9aYLLw0j
Su3idyrDonSoPrET6oFAHoQaAPbioOjLDmpfKyse+OnJzKovDH5t86yvJrhQk4xx
CIStZZU+0pkZmLhWEVUSh6JmAEeeNl0AmFr6Sa51yRJg32DUQBkYv8SZIlJucxlI
xj+H6EM0Ky3VJVc2fdeUoVo2neG0lelcRZDnNpQwRqR5UGAvdHH6NQzze6GTazp9
c90OjY0f3KxxoODFYDLBSc3bgQTAym+q92ROIfjnakPIMx6ojM1nenTxI/YF/BWY
daqdXnuvzqNwkrENlJ3dr6++5v5eflZ7INFyDxdCbr7Czpb971gVdQ6lgiXOAVK9
M1ACPTJjYwzSXuY3jgzDN/LX3hdarc+ThxDtEOt5nx7WIh9P9Uye77N6PTWDN7eU
LUgmPNeqAKGCgvn23Sl1Lp6pTOBIkoPCIR8PKEh41LzyQE9sXiYFBck67M/OK2lw
KkY8IVnWXHBljMrEFvShRbDSRrkTo0GwcHLoJf3u+542tQ9DxH8vD2KarfjkXJjT
hIRlAQv6kpae+6emCIS97YrN9PrPwZjmCi5nmWlYIMLwtrFD2xbS6tPKJJM3FtHi
LZduuQuqHZkTF7/J2ZXXTepeCmB+VaEaWj4bG2kNjUUjlxluChauMiCEF0huwvjn
IggrpP+d72oKIMPX1JT5FB+syNmWkW4d6RVZqcW+v+7LB2AHU1ALyaeg9bLPJ8rh
tM7v+CVFAZMM/IU+GrPLU17wWDdKXu3iLIz4e/S8xbQJkC9BqQursspN++G6GqUM
FcB4BsI65vdVktllco+bruWTm6jYkiSbocZLhRt6uR2KlGZlbyCki1/boaFIfIwl
kYJtX7FvDrbz1kXT2VNV+BHTHw07bXMYQ5gdwcC0uPE54v5O5OZ4QV9bPY/kK95Q
9ziT5gSRBblGsXaCdrRQA+9AWyT8F4dcFcg0xKgJOsPmI5NXSalbJcrbnQ6uFhyM
Zsr0LiTW2wlHMxwFX5ljLYUN9YFmx2IIO6tFte0N2V3C1pD3EETRmfBsmOMPTttY
YMNHK8WfChuky2BuQWZZtgduueUWfv8U8lxIV977KOFC02yeoxczYK5u1JGygAtj
b4RSVbA49czlQtyFVViZIxC70wxqWptuYQFNfS1rAG+o449cbG4eaBmrpWCgeeOg
gQd+f5vqZZdvqrWog6LsYoEl5k+oo0o2VLtsJfBasWV5ySsbZlPA7dFrdK8qMUbB
PUIRtNWOS/TZmw3CuCW3Oh9he2QUxj3KBTqTfibW5WAO+1GzREzjMO6LA2/J/A8g
7b4aqNEd5epM0IsLpynPKrhW06fGohus7xtp96tZgVDbpRJUS2bEFy/np2SUvLzY
p8v+DtMJiuTruQHjdnkoMZAkIRf12dW9ueY8CdanYYYIWdI0DCLiiOxX3xAHhBx5
zKl4de/qfmeeWOX80j0IHZR6Mpowj8/BSRacxk4W1Qx/aVgEvMp6aDhJNJuqjdfq
48i6kpLYbVljp0mnyHn9OnuZFSQsS1P1z7ly1IkNo8ip8utPpbu1YgCKkAXybdZ/
jNeL9ilQEKvH2DePSTWVOLp8YTD96tap8kNmOZytUSsZmIDp1Ax+dG84XDiHt2NS
6Q5uT1fmeEI3tSL7B+ZTMkh3c4BuPTcAeHP+fuHzL1Q5BZWSj5zWPUS3Hbi/0lgI
47rlGccn0ddi5aHgHswH5APbc9+b7nlUIQC3/ZSNE6j13NrPsu2pllc+ohUwDTft
oJ6slFLPaz3x3P/IRpDM5p0i6PfNB8R8uhnd3hhOzcGEwDK9E8N+YGsCcKdQ5OjL
TaQ5ZwL3XmR6l1TGUGOKrf5FSFzuLmjuoSHDC/cj3xMkyW5BsMRYHqoZ1RqSCh3/
alMpFNRqbYAyPny2k14XpTJwLsk+I2cF7zdb9rGT+TstHCpELCK+ZVSeYQ2udMT7
sjQWsmcG13uP6hp9r4+7YXWDl+lQnn69EBtzHSPHHYaSCYNBUeSVjUejs57vn0sZ
YUIyNSNzH1VCHLT84ZXR2am9TUru6O23/Jm2gKtNQDUoThXv65r9SRxIO/MRmH3r
4VA5R5XosWzaOCp8oaitq3mCumtFqe1ArfaVU73x/fkQlzi+xf0zxhRVS+YuCH8i
Vhn83LWyH7oMSOAsHfaJJa0N5OHMbZDPxDHxy5KRP70JvgI5X1Uq0hjFfKB3q124
0UWab+g5XJTnDQMuEg3OIJWXJqZ4MteJypeJuns82+1erwlZAYB91Iia0kF1A2FO
BRvhHc8f8q4qYq5dGvP6INznzYDBgVaJwRLHd7D9/FMlZ61rZpjGcpOqVnAAxhbL
6p7OX+tCSbd6Cejs2o/LjppJx+xH8xY2PrwbOW8Q2+SYU0Ut3meqQVPn7QtwNu7T
GIrKuoTxB29A/jH0e8606wq9V7SfHaMHKjrHy77ykUHIxTNvtp4hyOruO34gLQTd
DU9QxkrNkAQNsW8n8EQLcgAbR6b8aRfx2/bijm17cDrJzS7IQHbo0wIr34Fdhb7Y
8LBD3YFglzi+TBcIvbUzoafnCMylTDFLWBXz9ck3bWUmdVwzVlO8yp0Ra9pEHxRe
DBmV7E6L1fmOW1f1T78JqO10PEFKrv6BmQ4eYG5IqFquMMiHxgPhFc2Jcwl40n0t
KDvsQCzowZtd+gPceTbOehkjDYAhJ5skAkbBNX0iUredtEGMmdiH9b9tjUfdY2hE
Mc+eqotDa6xZ76TydYFcKmSHGBP9h6TpR66gIn12G2vLy6b5YLkc1WHxtahVFK9J
sB4d8Ip/8zlwCuLHYvgT7MAgCUUXSL7r04Vn+dZ1RJH5rDFgZMrEt3c4Um8p1ll+
QO2w5SrE8xw5XmJB1bU8HvWpinN+cGCvyq5sFJBscOsu2TVdWTPL4/6bpmxE9ToQ
PwDvO/RFcg36naiaE2s6AGAvn6O8kiIQsDLcaMz3+Monhc+c+ze59QMsKNbzUbSp
W1GZjYVWUTO1jlfwx1cY+TAURLgO7YY8s4WHwtbHjHgTDPbWuDmILPpLx/I8Y+ct
SnzYmHXLzRLW1FG2OpYMqjzaRC/uoyESz+NGJSNitUK7do6PcX0Zyx/OR4VEWURn
nDDCR3VUBmTCtMwrBpg9Z9e4+BklqKmNk/9QHe9YKlEkloUbcYPdp2Nzb30g2aGw
2ZFUSZdIQkjKpw1I6+T2K3K45g6cPD0G191+aNnpqRAt34wtKqXAQOmJ5h+L9sZ7
GaIhoRaVcagxLlRwc+FTRDK4oG/kLIPOplVfjWJ7bf/bCmRIaqUyBMrwWMviTQuk
hnDwqekbqyFF6cAkE3aFe21VQoVSccdTavrHn/qlqKlEEZNAgCKd74vutQrbjytQ
C4rgCbDJ4iNYaL3r3pdTYa6GtrfIT8vfvSv84iqXzmdzd0HlzORFtdEp1wdQB14Q
oC7GB2pVNLM+6984iOalHJf9/sM5haq6oF7yw6oxhiWlO2b60tC0DtcHaeolV8aX
zrjILnaqTG+qGJ05LXEjchC1ORHDyJYw/zR5PQkKRs1nzI9z7cd20WCQxTwq8LEH
jooe3rDmLZxWE6W80T/lYmMlHGHV6oBHtH76XKxAR7GdG2eFScWwVL/YhGqN9u4m
UayMIy6rnwTIXD1IyhCQkWH10mhu/wsdiWMP5N/y56Bxv3ZC+Co8BmwijOqFXwD8
shUpyUkG8uaoK2PF5obUMqVxmQlDt4MLxxDD0hK0+0VmjXSQR4P3W2eSpO/u0ray
OP1ruDqfL++3lBN+Z9DZy28ilx5RDs56AuMa4qabdI1wYamap54CVPrHIu5krsaU
g0NstWJ7T+Na3RZFohLmK5W9bBe+uwhdirnMD7fkrpM6TgAeVdGCGTj4wExy/UCF
ZJD6JeB81WaM04BWe6aPDptNJb6eKYocU7OvdbUTvUqJIcPkKvcydlMit8tSxxyh
ik++832HGRkQzXywOUwXFv3HRDDPgjJvvZ0r8eE48zCoFRHTusI6uBEuw9mMGH7o
LPTJdauVdM7C28Xp+7ov9mkh4a30q++OOQ0rrz8AAXpwv7l4mCwXFm700AXiHZh+
4xLx+uuJD5yCxnLZhHyiF2EfnvwU769dLONGhWwzI0xkB6QDvaZzcaJaXWrvUWCz
0ctfUSHTCotK3jIkxIf31yJZT99OeFyB0Sq8B0LN/hHR2aVGRihGfTXqrb2N2F5I
RofFq98iRYV09kGiX2pppycsRwvUuTxidxj52uSqNIDYip8BGaUtFcHUYcUENVAx
m09gWgOEVbXyLhKBbe1wy6OYvG+gZgtu7KZ1veJzvKPY8y08UVnWiwJIDdMDtSqG
nkZd7EurpE5L7JrtJmwT8cNNDK4PVYHnzgX0IY+APXCQJPiou7UuKPmXAe9iCInd
kNN6cU/UpevymeAXct9KyL2koKdzd6QiEEANXGvfl/f8NkZDqn598FMR9NRUrPqB
XSZhx1mJcpsmNDNSPDOKDzyXJPArSMvuUtItOrvk8RP006FTyy1cb24DPbdYA1my
3CaHxZ+Swk6oyBDW8AJha9OPBwTYuslhx3FRn+2LfEw7FF9yBhoCiM6ls02Ka6Hl
bnyn/XKexv+uVO2RUHGlblobhuJBOYo4kdP1X9Q0k/+9++1RO+PgC5wMeIWG5rZt
k9w2fsdTIGx2ZsV3Mg/+tULQPPnAOnyU2ElAlTJ4UaIk1H07/teySj1KJWRN5nMt
EGh+rvR8HIGAIt0rXQpUD8fbSwuI7e8EWa6QtbQ97rVSXiYgjQ6h1KvYI7Zu1URy
4CvLUImnou1iP8DMqPDDcje7IVhFdX6ONQ4wof29pnQmVcaWKGaJZfWXfjynVplj
E7NhBebCcknBxPckwK1MTJYpTWczl0XzQoykFTvHotc+MWUcX0HOyw+Ipz+kRkvE
ldU//t401hUe81U7u9HPw7ea3CVXXFfNct5bMXqwTOBzDGu9ujYLejvMiyJlb5ZV
XzeqBzE0OrZRDq6JDH0YnWwt5Qj5w3ZzIWtUjYDtWfp2EW9nom44HX5ra+leTExb
PYvwGP5MChohKAeV30ng9dByKygVaSvV/M5/d5j2N9ND1+dDIxQRVAi+0SMnbudy
HAbcLaLdYzVM4HgpLI7Mx4CyiO0uPfU2hGyiSU9Ake9ISaTDODKhs3PKjDD3LUuK
1WVoudarYeOQN9kxe9Ma6jFkwXNC1oT1d/rzTEE2VFmR73o9Oj/7LpKk/kTbYEkK
E7hXZIDzlNkFKkF1x92oRK1Ak7iC07hu9vzUfWwNHfQ2ibXB8xkZUOicbgG5F/i+
2cNBcNGdWoDFezB8iyMgLRhFK7MDR975ayR2+3HhM7x0rIyMMUwo8eJnLpdShNpc
GF8leZdgl6+T9znUEGV8ajh5iVw2xoRcemHZd8LLTyRKJ3GwPhnUEShR/Z2RJ9NO
VlYUsQ3pi6+VplVzqyLdaFp83PtdqX3uQxm/Z1yKhNSarW79+50wW3uSls9G6PNq
0bswvI/zt3O8W5JWAKWScEHETWp88J5PZslozi6RlcZJD+3jV84f2scCLQiK6sjU
cpbsyy/FxRniYgmPs3A5rMeORc6M5v67GQoBbTJEjqEGhuhwns3nV/mYJNu0GvN7
UfX0zwS6Nn7zef9AaVEFWiDt2QHNMUh/w1g33VoP8dTJzjqLxAt4nmCy77Yps8lR
a7i6dacFNT/zx+0EyGbS+EZLf9RTWr+DBOmQOGDN1c1lHGkmf2h3oKzuhCrvxHWx
5v0eJsgBiZmmY84oj8q7yXjkDNzutbbve3uOODvFqkWtDb1GoCVu1jHB5z8YJKu0
tBQG7tY6VuKaLROEgf1SBk27ExGztY/1IDQ+KSEuaaFxZOfmU4lTtqs1PdEagCH8
+wJqJHClcRP1D67QIbUgff9YuxX0Y8geq0QLsWXHvxqfr7zKRWHtF9bJXE1JmBIy
LuGLoNJRU8QuRekEXLsM7TdWtXjtK01Izi1fQecmGCmN9LokzOJ6KQqxQwcR6raM
fPFg5mZ5vod/at8ZjVXFG3/6cpIB0MbgcVN4f7/EgC6hPe51xRFqYa0nRZndmiPt
o8jcA1j2M/nDMCaW4U3hB6W55b+doCgNj1KqQJDy2pdFc+eRWV/frJE/MEk0h3e6
8hdVPJxdvJooE8Kc+uziDOQjMq7uj4u8tJPsi+pyeRD5qYbbagtp2S4CJ5tOVdy3
TUxAzf/OpY3Y1g5j8a0EZ4N5qIcAaVD0kdq2+oW3bUT7Ibz0bcESUALZMwrlf99s
8pYeuCiluCpJ+EJhCc94jCy1hp4+2E4cJV0HZqfVBUXXeAG4RSvlTwikm/vmNuc8
KWwsTfTwKZ4eeQC+4GcKpNAJ9Za7WunKfr78Qr/UuSXosZ0xjymrvX4X2VT3vDF0
1nvz2cMkmFHhI7gPHuw14roEBIvbvNx99yYs01r1uzrWvbKIqW9QcoWpwxLldHWE
IZxiACMD2vR4Imm0/e2ATjm7gPYr1cTSS6bl8KFR6enwYs/U/4ZNn+s1H5Wnc14D
V9YaKSIdjKFueznn5QUr47H/Fob45gY3vSBryYMY/mY3OJAtJwY7O8vfMCLC+DP1
JvotAsw7MF5/jmF9cTOpkrK/Z2hZacyI5JgxECtw9tq/17QDNjWcPz8uCAS1aCtr
56vWkBq/tmY5W0mY8AHJI/L6LEkrbqbsla5kxJ5QHeTBjr22fPjaMXIV9773W8zI
4seUESv5CpFckASNYfGA1jFIuDBt+Vbs++gFrShwNHc9nQUwaV+ltUJLWWGBaFwG
GZ8akmudpPlcs/gdactsxkWmZp0tnkkfy5y3nopz36SzeV0cs7525yu6lYwsBdkw
GO+U6HdjHyXUV/8MT6kd1BC1wxfZKWqOwAbncozspSzyEFh/CtgPDW1hJytOcFIj
4C2sGUJqQha5Zrb+p2evEfYmPDA2ADprQDUtjwA+e5mIENgPm/KHyvRw2Zubwbls
ItW/7UA9J6nmV37vYfuSMdBTdxan5cR1ddsnXBBjGO0xoFebm6mWNrLXssXaUl0A
inVFVeYYXmoEGckLIk7fxQRU/JPGwLapVL4e/IeSASj6mTQrv+huft7lhsqNH8hJ
l1RE+e5FiuhSzb7Llq5u2IIoOzvAC8s17Nq+FIgoI7ET1rt5neTPwGad8UCmqdtK
hWhMt6xOdw8BjasY/LMt/bogVVS15VIa/9lf7sOp2o4L97yUVtdAKlTTa4QCF0mI
og7F5hiVq0tVf243yrOB2OcXk2L59J3utZstGk4FrSTNuq6Ym7dmV/xIJchKvPTu
eAD6YWIdL8WisfMVG9b/X1nOvQwqQDbnP/DCjhCAsKMUun/bFBdaULYvw0wyty4C
qB9tzw4FsRVg6zSs/3SCIoAjISI9gkNh7PETsgnI7BoKyhd8jt/kNvddeXgIyb0b
/ucvGYPR274fSiHchiyTHLCndzWMyXnbS9isCOCkh3WjeSz9UrtfTq1v1kL82h+4
Qt+yBf79qT150x9rHfw9thcgkX1jjm/NzKTwJpWThabcLH6qYvL53kmlKpsju8Yt
natIIGQ4Ovi0kaNPAFx1aRCattxLrzNcX+ZuFezi9FFQ2IMZ5Vbyn9tqR2ICE2sr
foqhVOjhuRDa1nVIQcLh87fZq0vLuDd2gTTdwJfrMjSbCYlZjyrwKFCHDsHquJWX
SPbJmibn7qURnsQct/0JFpbygId1QqnJSpEI/fC3mw1V9mpxgxUD+JiJEBeZKtXO
T37zIJTxAUXCl8ERFJ7Ky/xaBLN7zV/eaz34UnEo43rwtN2CxsoH7Ajp/E/XwpVu
21zhSDM8f7BYJc5mkUSbLXAOz3MMvXSrKtd6y1mHgLXR/56W+v4IrGqwpFUvJ1FL
1C+Mt9Q9Q2eZ846WsuzhM1aqrEnxzlJTFelbahBGB/k7/C8sKWUa6HWumGMd4yZK
7zWuZxnuBQAVNIG6NCqcmgLomSlxDFXEN9+yAJ0V96tT3Z9WzO22mT2vF1e78DcA
d5YHRCy9mIwHZrmCXLRIGXIvX/vzNnEBVzZgyZCUx6cLjMK/6WAUKTo7rIDSbU9B
kkNRD4YrMWi/qRZAm1QYW5ZplCwS4q0znhiDRFYskLvMDA8YH5AoHUncUZYKMGmk
LkiU9es4xixmQWL63rWiZorovHj2BsIhnLAX3w6om7u8s99wfg2T+5gzdx8B/QtV
RKr5vdwpPIl+jd6omEQMRNe+NToSYna4ZPr0ghAVOS7UO1a5IogOYVSgddcluJs/
yHp5sbm1Zaw8lpd1MT0QzuCRCDWieR66ARvJywMjSXJES2HN8Ca9AP3mBjzAIKhB
ekX+SadWYYuZQJ7FuTD8KQR41yOLKEnBXbFpUNRdY0hRWemTSBQDWcV6E8C8VT6P
qtKlvKpzir+G+pD4Xpv4nuvHr46LCUHE46UuYcEpTeHsmJ3IyDp+PYhWsW1jtbS9
tzdYzdb5efJ5Y9z3E24FmA4buH8GyRaiGM7T9IBxS2npO35LiTPTgcKCy7PAhCj5
Kx+HVFFkdzedQ9hqxzFXgJLyQ2Veb4S+EFAX4IeK4gFMUPjS47RMizxBPUzlGkPj
09YQT4723ktvZsTXhkxmquxVIpu5kvQkA5kNxk2rzHyoCPiPF25V7O5PkedPk2gR
bEUxnwhLmAzyt5J7JTbR+ToC45zmjlFHJrCYzBZyxALlqfKY2I1yLHyp0C4COqYt
xW6oHzdxN6Eb3dI+Jqwi+nOxFW+tI0ApX4AtySIQoQpmWPncqtOq1C+vSCKFjWw1
bimh61E6xQVQ18zzd4HuNfYdRgaunCXVGBmw+AusQdL7mSya/vTmFHB3+fMTfEZR
crkogOmzL93ybhB0+TyvkcOEHRJAiEXvmmsbNy39k3U9N7Fkm/eqHhVAL7RqAPMF
06MxtnQi+oJTRZmkjJEtFNAgUWyZlHLnZGpkZrI6BNEANpu/dIBPHzElHTD8mGlT
nq6rwnvr7BvfVxQBhG5Q8S9+nZ4s+BqnfDYUAmqfnDB98Hm/PKEIYsyZg8sAxaMo
7MGZmrGpxO/SrUhvS0KNcFz7NuzNwtlAGQpBKAAVcwB8UVHtw1Z3I5pAvSUtxoLV
mbB8zNDLeXagVumqK32RHSJbugBEwJgl1B7gupXMc0MOnUshw67dJewAtfcXd5cX
+IQDHwLQHCgGY2CkYDSyPcGhy9CR7afTV/gUO9+2KKx/ZriUINtQ9Vw1czTLS4Lu
iTfulGSjxBogIjRgZndKBgx+XwAsazn4ysZOH5lmNlzTurlbQkm5Xoy3bvrkpoaR
H47sM8AUt862aF/kcUllV5usHZAe37+FGgN16SzRqDrp5xv1ZCSkLv0qeTWOpYFR
XaOIz2ZdKg3bchq+rqqyS5Tu8i8YX0e/ApWx2yZ0eVL0IZLAvFIC2M3tQT4Bx4LZ
c57cQqArECMVeGaVWqmSNjqu5RLKXkXz3W0X23RT530E7YnVayMgpWjC7KfZ/xlD
k8m+Ke6LZTqT0OvzpVnjhTgc/p+wXuZrssgIoqmPnXJzULGuN0mpRmwc0XNoCqvT
ClQyVyKMO7rUGpdpYWRQ1AbmE4Oo/QACUlkUtc0lS04FFrEp2CfN6ArcmswlF0QI
HMdzR3sJNApE639cXE0BXaDdxcQBb8jFtmrveMvmApR75DQtMQReo5TCMkEAaKGD
OaZOXeL1BZW08qC6T0OAJ3pxJbz8hGDaSmVBgayGNrK33B7MlmRHJCAJZI8qJoDS
3JLT2cNk2qqkWcgtjPaLuAhLBWu3ehSfLkJoafDQpQ4cYmC+nlo+IuZz7bsaF0xR
9lAuY22OiuA2YW3eEukIxyvLUIdIM1AWE4yMm3Rjwqq1C/zzl5fUR15T0HKmSst3
qVsPocTkfRXsm+XWQF636w4bTKFydmW7m2EUE1JpQ+jUCdhhqTw1LCR5JXNhi0YX
ekqfXXuAMnzAcwbYftruR7jE1QiurVCD/PFp5ea8JtXlm2yFaF2Ul6D1qjHCYPNh
d/zZn2dFBJQhGxrfLAGiI1VMjeBHeSikPi4Lsxt+6BBJQsf4TLS9658Pa44RVCIS
t7WuCzif2fdkY5Sjn2wq1jBdID5KdryktNAKBcyrvdTp9ESjL6shuKpcln82zNbf
sl0k1qQPjnGQgx9IxbqwT4Uu0fifgUtHRDh7wfAMZz9RvnrSQ+ml+tBsj4JRxZVH
FnM9OWWpjvU26SWPk5LNxTdG0Om435UfTW6atUMLeyuEkANkKNuMZhx5dQr3Na3a
3PSjfP/u1X0XMq21SkIN25pZOcqE9nVLarLYlpcCNYk8VZt7PoytJx++OMZdYU5M
DuAur63x6xoQZJl+sdi10H7h1wCWdQpTP/QHfLv4S9wPknQF0/FIbsbm2SdYnRYK
/a8URbS8YSESNEpM6aiJardb74dQdauVyjc3B9Slp3b0s2ZD1XcjhZGoQNwWyp+/
QqKhw6QOTzazmGfWRNXeQxiXNAdOkIslARsB5E6B4iaCKDS/Ba7WH5ldimX3tH5n
N30cOs7H82UzPnjZgwNV79LmtJjk+X+FP+14eFp+1lWpllvp7bY3C2Cbwg1YYW0w
fZAFt/4PHSd6p1GX/S5u5OsPPBop2WeG4Y7ZRCE9a8u2be0NQ9lzWA2DG2u+oN0Z
jhlW0TTLpFK2V3xlsKfduR1KNtrx7Gy5K4jsPKyb6En0GaEUnaPCq+il2xaehEaf
9c/uC1vacUL+U5bUb659qZvp6EafuIZf6Uvm9/rhOYGNOTutsMVVQmif5urFrDY8
OqH9vlVD7wSVwYylht5ZaWXBd3PCSyuVA1lx4Xk3W9fbbrmqgrVY5y9C5ZVToSZz
D9wjtePIoNFJdWaJ3NyB3v9Wcy6bAl28QiwCZ/jjOpwWq3YVkrXctIifRvxCMSKB
X/95y1Qd+wOs1jTece+MsufTOUCQYmtllce+09L7M89OeiMRrUHsUDwqvaihzGvS
cpuFvOG+UPRgzl9eQHkHvMrHk2mw5EimBDsypW4m23e/ocSJSJAsPVbni6d1P/1C
LpD642Zx9oIP3xyzYogWCgOA3+k5BnuLVQf9thrGNbh/l6DqkPMtNszygjrmeO17
QBTIvlPqVUW54THe5MR0G3jVqwU+xCwlo1L8wb4aY6PIOCJk3th8Yxa4dVc+OSEW
MwOMWwy9hFbNWna24sa3nTPBWLblu6hwr74u60UB/Q/AhlCFCalT5B+NUP+eTZkr
YVNA2f0ataDAjt8gAAuOQQXIW0mEy2+vx7aNfj86vb14jmiCe/M+9b8axqKwaXm7
tOvqEqvowWb4IoHpWumFOfDxECpfVL6kllMXAQB0zvkEBz7GloqOhJjQAE84lISa
GxB04/hs5YTYh3+XdovuBDOcFJBo6pIdasgVx3tV3N9KVmoqu5NAxsF1zgrgBjp8
VxNehJc+B1/K/P5qOCpUvA/wlwrjRxVVYvF79HFUp3+fGa+UdW1bqY0ED3wtqhCO
eiqAq4PG38CJffvNLEmcQgfoMBIeRricvbVdAciM44BY7oLqaURjGteTEMGI5Ibs
VmkNhGd4E2amWsMTWT6MVLe740AtHE86HI06w7cstAPtO1z3aO+Pm6iVciKBN7q0
8HI7vp+it8XRJma74bai81FV4M12haJ5ylkxgkqVVI+YbyrAFsGddiWzBxt6mjFY
+mzezJxGVu9v6z7k4b7hOdxTI/yGxEQlxqqOqcDfWmdT+cB119II8Amof0zHUy1L
jF2S/K1Y7Z1yI4X7EAZpWpInbbOdpf1/f9uWGi6yDu1xz9n5XYjbadrptwqsIa48
UZyJaxoBpKq4vD2EVnd8BBRj1aNckAIGEYQKx0hBmgIJRoPxCLvxZCUme+dVUW10
H03AJJ7ek+Lq6nhA/Oge2OWzPXs9rCL0HsNPE49/uKBjukvmzyXigVvO4TULWteZ
ro2fHworVOxZW6tGCqahFWoLRuw31Ge/t0772se/ZDvBJb2OKKBGsRyysJ6RWzAz
X2wq2Vi3Ej0xKBQ4CBx59Enk63ODUoo5zdc03dKosdJSxdyAvhTe2/eOU2Pt4pMh
XDLUwIivDVPaLfrDiaKlKrYehF1iGhlTtqcQC6gG1N0/ZHAf0OeFIi60hw49hNpX
alEU21ZaptoNlR/nFnRqqbHAnGGt2oUiJXYhjhHAi56DwGAqLYpHJmKuE9/PRAMO
RI2R9eumnnX0dt4nHZGXM+qxcGV/R5OGGjdKFneJhCKekb37icr2QxlMqUO4DO2h
cv/vVvTEAKR0yv/qudd3chns0g5QWma3lfU1PzKzhVyD94wyZlVUsusrdli/GOS0
KhK7Bpez+/FKctQPbc7AJS2wxb8jin2CVE5sXIMQRM3ouw72+qz/oNAUbxFUs/VP
x6FDDRK6ZJybMPfJBfcKq1BQhIeOZ5ufWAXJV5LUUNLQNU5/Kp5MLLgFSifMin4u
CkOn+qqj1i3X1y3beCQuGR05lm0YuFbk2ZuGiRCGX4fLiXrT7mF5C8or/GRdNQRB
L2vD+U9F7C8ZBlDpdSNph8STzp3oMU+IqMeQ79X3POsITcxe+FLwo6+Wxd54Q7at
WPLCYWjowOnxJVgAJd1K+oXSFeFWC2eD3K6SXHZ3J/YEd9msfMmW3Jq9JEpPwbwW
pRgRmwPZyApe1h/quWyEbDLQkmtsDb34Y/T9+M0YEagxrzrdtvHtwhZMZHocw0Ew
fBJfGFQ3lJzpdkq/VMLhgH5GLrk1ZmIRWJmZLX+tsPl/yqWsjKjfrLzrcnavkReW
Vusmh/LHoR5bGLa6P5jXQiZ+l1cl4GbGQeJW4KVPI4qCQY21SOTAIMnplzqqm95z
3k30KnFk6R7Z9KizKYqy7ATE0nBzb8ONadWTiBkU04oxk6YjVgAyK64tp5sqaHcC
r/nkGywovr8eocJ2ULTLt4NMraK07B2U2kSMio75JfZ3i9mgfv30ktJlXIfSFN1s
o4X5zrw266yPTeAMtuEP3RqOjZvG4mbFf07YndyCcHLvTw3Wmub1tkOQY+Qikap9
3RZF0BMX6pG86OdcG7cZYixvzFcIh5gygHqF4JYrb9bbWpcs2FfxT4VWKfzpwolN
QIJZm8xOVOtGv+laUnetBn5KDstgWGqKvbaQEXsFCtqoRcTdcqqbKptM+JLZFSe+
frHK0swjwp9IXDmqv1S+dUYHXWs9P07JtSE2v7CUjETrSyrgbQ7JcY4hT79cuO9N
EcsLwvOue3gce62fXYed9LpjZ34/ha20jH2FNDdgrg3Ezzo1vA/LjPWr20CzF8sT
0BLgpm8oQr5M+dZx3FHF0TPXu7r2EWxVAoYhVScZfwKC2gichq49JA7748Gp0xg4
2KgZ5mOYO+m0ClZ1cUo7Hqj+Z0I8ZB3uGX5sDxv6rXvgkC0FrjikiLdfqgzebDc2
lGmM3wW2bVbRe8DgVJmuaR5RJtjp2VxRbuMEliFaPXpa7Zh6J5nnkgcOV9Dhsrde
xS+E8j2Ys0NefXlx8UZAMLJvhgJMRv2fDp3cM9pqXSX5QUHligTnLI0PDwxLI13W
UAzCqjSZIzBlT35LPJXw8eWwKqhrvJ3oJJdeQOdJFyffiCD4WVto2dVM9q/BbgPZ
UU3G//yjhujeCVi8k9MrBfxQBpNMJLJLGCMS8x/+WdUGN4erQ4j2mxmC16D2+nvG
MRhR/j9X2etzcIX7yv6v2WSZx/984dgKd/uQxg+xr/4PcQ//pzLb/H3u1MFwdDaQ
jTQpPqxgh+1BNI8dpj0m7qpwbC+2WBMRInXjjMXz/EPz5CzagCqe98e+OJY6FJRG
lnzbxsN768NJnkpMT+k2Z8BKzTJ9OYADHl3fxnWuy4v+IX4fRMcPRRF+y4zL6+zF
WX6Xw4iUszqGSR6pE7iBCbLt9WHrOpTqFl/Tc9sJpFV19t6+y7qt6yBkqbGYxMYC
cBUIphcuVc0G2BscD89DljtNVSkGAYUqBQNZiSl5iBKGULByDmECNmSUjBqef3/q
YZ1XvOm3a0Lk+6/FzgoKfo8PdlRfS4M1nHWU+n26DFu/bp6I8P0o0qjeSx2JVyrI
K4+03/FaBuDXX8Qb9h/Bu+PQmnwryUnINvb4I+DGUt2CFDldbHI0gCEu16yVCksn
Y0CYI1te8QbMKfue0sBa8WsROambP6Cx4hI++NoZLM7oFAkfJQDGTFDvHIQYsgdC
40l68xvgdlVhG32Y1yOxqU//fYovWWuiKcodrbLhZiVJ3OIQ90TRrRvLp6e0lK8Z
NlB/HqFV3UJ0PpEApIpBuJEQDqMNS4Rg3O0lAE76m3CHMk/3LTo/ntHOunKh+rAs
/Zw3VQFHV9pMJGePPuqJPXCxQMNJlJR01CiWg5OHbOC6wWpbuoIDyv4xMGzPYXHA
tzwJvxkxUIjVabSkxHzvbiQkK0QqnU2br6Rqt+3xj9WpAtfSHR3vL0FBvSyAFfoz
Z5ERFMXT6MiYEEwQkkNXRWQ5p+nFp7niV9eLr/OB/gZKocU/9oeFtMpp56GclG7I
4KN/bCB8fogdOYUe6Hqj69eJjb3BrmOyFnt+PIZd9QiKjXkit9Xhxf1Eia7S19Pv
LeZ2TnXqYFoztV8FU0NDLp2/povIpsaBW/u9siSMs2jDU6suRvoVxfzLOXrR0G35
dQowtbYVXRiCJwC0D0LE7n8YDgFgsjcmYDfA86hZM38RkFOQHEBsb1OIdGuPNHNI
SDMwXGYs2NZDR2tv5f4J9ucW8vTIiJJoD+PvbuN3oDqbm1xyebvGBlb69DRBwJDP
TujYoEXdxYEp24TnNJuzjhDR5EqvBMJjmYbzA3Qa8+ohvMD1z/frTACQbWkzHNWV
KBKc+2/+r1PpM2yZn2oFeauvqIQK2BPVizJqJY+vpQz/dmo7zIBK0OF7dqss6Aw3
8Fua0JeEJ7Xv5EVBQ2z6ti+LOV81bXf9LaDf6tuhj7lfy/M52SjEveuhPVcAyttC
JdY/pK7+xKF4wqypL7lFIREtzJUKQnSLqT0CcEl1lnmsz8MgGSeBAA2/qFLFJb7I
ILPv+3gDWBFG/sal4m9y5T1pka/bzCih0pR+J8aS3o+jxax7jQTva3eMFrYLmVZY
0FfG1YkovuBmT36l9aPd+Rq9QIqTJPjaSmaUNfrsdAlJaEJBK3YDqdJF4DUEbNTC
oCJZ/SVZ1kmXOuLsbbM1hMd+Xz76A3LhLZhqnuNvFO5PuzYJp68GkkU0lw4lMfpr
VpgmLoHEA7JUaaaZVX3RIbckfwWbBrlLBNTP1HVhVcIyrdlDya00ljW4wlQ4f5PU
40GXu9B4SiXkt+gykDfJVeCCKrmPf4jjSXEtEMDjfZS5Td7K1r7GCeLwtsK4SWmJ
EpMCJcqn11JMJodPjVlj7Iy/0cpYGqfN2iBKG4wT/OyjUN/eqwUi7Xgr14kcZfH6
ORWazCyWRTwuxpqEWf5PQuEo8qU5Gek9fJcCbEVKPqr/F/BQweUQo3Ud7m38Ia09
mpZXuDMk5kQX6A/Q9PD8MMGXBpUMoABg7aS8qM3TUd2k1iUL921xi/JTfQWY/gSk
MuuQDNgkDRqUtTFgyCXLUcMAhV40ELIuH5AXbs/d19EcBwyvs/5T70oDtDRhs4Nh
+CXBvFAYQc+A8fkLN/M/lPG0ZDxSRKiSSNAuFOhgkfy9x8e035NxVt0WhD+0E0e3
Y24v/3eIPjUTIeod80q846ROACyD3DOaregrzxqTeD1CZsB0Vl/AC1t02x96MJyw
4XlxCliZuMDatEqwZMorVT6WBONZE4d6GWWl+YHziiKMEMYnkgEKf6JqE7hvMbcE
vc6sCyyzFUR+vXKuc4jqJ6eQWcVk2cVk082u4WFxd40ExgcalUQ13d+Q/hgagLpO
GxFYjBkbbp/+E5zcKZw0GwWDbeKS2S9nAJ3GhelUzzq3LEB1A8xcp1QmeeSWDIub
k3/PLYnXM0aFRPy9eYcK4uVMSjrY2mm46RwS2HLezsLJziC/hCvUUMl9t12ynIXJ
wqG6dTED6xeSLMClKulRkZ2FchpyHqIV3hXHrIIAg6asNk+vnAVc9TTXTf+SkPlH
R1FWKRRxJEePtHM/BQmZKd5mMCXMxo3HssUF0+yMER33EwWRkz7AJlM0R0ImCeVX
qzlWDj/vuvZBxUJs89I7Ie2+3dLd1qWH5Uf59TbJg8nBWMfQ+EbKkE2+r2Avcx72
LtKh4E6hu6Pp0Sk44YCxqVoPJzXwdDQmVlLoDT5T+2HTIbsrp+pT0k5VYKdk/F9e
DYrzgMHroaUnZB4e92Rk1VdQ8KfTtaXZoGnB0iy8dWIsOAWNzminE1WXSVg26RaZ
Rt6f2CjnCnsuikm46erm8HKtOd6wZHKWrkrrCP1MLhgrVPw1RK7IqNit0eJ8T4ZF
5cAK3apKnsG43CKlaY2U7JT7c/mG4ZAh2LGupEpaR1VEctC0G9ILhuyQrFpTUQPR
V/bOUx3RUKovJX3xIiiiRwUJISXHD+4jQywJfBWuo5SS6QGFq+N2SLZ5gmFpUL/p
3flowTyeuKEEquSa0B6zKzW9cLn8JJDsBdKV1061ftDNOfT+m2NyMqI1qdWs44xf
CpGutVd0NO71OzfHK03bpLrf3/MDTZr2eQ9vdjUaDHKZfmZD5aYB6IR94WOlgQMs
E6pwszwwuoJqwyb56qPH0vP7riYp6Mxc3uGrVi7MlLl1Cq3ZDLTeNZFdi2KuVIPH
6JqX51XSCfiQ//5GgW3hj1b2Q2tC9XyZ1F03YmBzYkMMHX0C/aaRxnbGxsJ3s9Ma
XPN4gEULFuZdbxC0niR2tOlxzQMleU84UOe+LKdxWtSs/ZVofClUQwN+T6rLDWKU
UXcXZgC911eyhOv5iDZFuU4weweDtLrx4Rz/XWzGA1IQvHg0qwx6a+t2WraUFKas
YNgomAH19QXPDny/vWr5k4NUg7KiNDd50SnUZSx8Zw0WktB5ZWJ2x5E/FbMpgZH3
Ktby4pBPxqYgOSFJZwJBhjHPhI+8ctbyco0N7ALjlzLMuM4XJ+/lpg5UbO8KVTRf
ULQ2nmfVo8Rvzc0lqkfTlDyRaeS9fu+Xq2nbGKWYSxPwYkzx4wD7Qy4rvuHsor38
rVKtcI2QJ6yPjbtaIHHRg1Pw3F7vjMNW6GEM+mYjCX9tfAf09g16PRTS3pwpyiF9
pfdpF7PmfyNKcNJifhwgSOgqmJ1DslEohutLvJWyMjLVbV3X2Xu8RX3F8aZKjHJM
e+gZ5blE62xCIOLKoX3MG2ADP8HnN5UGlQzC3nWVPIscky7I2Pp01LAQZ06xFWf/
eOY4Kwj64KuZ774yf8PvP/WOY3CVhKuSYzLizgVw0XzDIDjWcwoDvh8nmDYhR4k4
QyQOH08WI8sWQBFS3IsO4P4Q6nu1g8r+S1kL8uPmAHNIFdhx34Xmm0TRFKL/SVD0
nHQ3d1GNGt+A9ld0IUyVrCwJW5wdc2lT1baWfTRMmxl14mCq1/uSvIxsAm4z8cmU
qfWIGo+1acU0l5VKuwBwqRK2EL60o1ZocabAjWvmg/Zg6HiAxYT9dgBih6Qw1x0S
IkXFck5bJZ8M/i9riW8wna2LtQKBaa22KnSHUwy5VpcWU31bFWmEKo5ClZo1dUvO
tD9LVsr9FSOaA1VZ9ZvPL+NrMaJvpQSXjtY07OQ57dq/kMNbtOhR8e8Q9LTIa+qI
mceh3+Hfqvx2BYEXgJviHFEMR7Mv2Kb201FSeO7wCwuGq++GtAfQ0WGpQYcwaoYK
Sc08SEUC4oCjazEJtjKPebeeXArzc+aLfhm3V4XWCkalBXTVKeJRHO9bz4TvqGQU
oewfl7991op3HLz38odmBeY0o3wJyqQz1ZI4xlqD63p5jHgdeKUPHGceIC+C3p6l
gjGpq9paD74kT6OUlab/6xHIHjU91mZ/8lBTrVMOOrxqHnMIj2lTEo5KkTixQ7Ys
ducSNL6B/GC0WceBTk4CcdeZ4TRVCBX3BRap89br6mI0u0jgHYPiqUnjyBlihA1V
Efp67qkSDdoJJjCadGjtcdOqgyyKIFm/kGF9w2r6KrZKJuz0+W+lrnPBfL3HyZaJ
wd6+yQyuSbr4K0voNgYcfP2pNbDnHu99zlf739ncVjDhP85GXEfNdE+BdBYQSrZl
x0xZloWPYjv1WbXpKZ6UP23yUXiZXWOrp3gTlvCVVjiqW2xOGI/CdAgvHSbhLBT+
Y5kYiiMep99siSeEvmRf0Gd6JZK9l5BVSqrhviCGvsN3L0e4VrOgukFFP4iRTAYo
foK7+/bWtG6kmmXHAdLEcdqpBYM6cmE1xuJSrrTLslyxdxq1wRt76+ANCNVIH3Cr
h1Yke5W9hJ9YRdyGENUveek1vNl0YKc3xf1Q6hz4PWMBBjw2UpQ+HGGlGVjHUO8j
D3Zazd2nn29if4CGw9QFezdjl7I/S3opQAN3X6YCINIJe7jLo8g/+/iu8kKfAGHV
41nvCd9ZIzS+J6Eo7moPTP8x0kW65b95DZdpOsIfD8Z/Oa97XHJSFZKJ8mkvHlOs
4Sl+l7q3HnOFJ/pSQY6DsYsNdHDsxfovOjJBftBW3ivJohVq7ZhJS59ojJT3H9Bq
rrdzH2z7gBWz/XoDwrU90ooHrbtCxan3Kfn8d8BRZCIkGDi9Zq88dyTOFfxzK/Hz
TkJARv0GKyPipTFwMJBRlU7pJneMONUv0rvEhUS99VFYdXxDvINQ04kkmojRtRgf
pPowtj2WaOKDaAAhiHs7ATTnQSe5F8bcjF+n6pYntnUYh8e7VzXOvMllZdIZFP2Z
MN7ZigMC3cuZOiGFrFqprpgnYIKv3Qew4Nym0sE6LPDUAHH5qERmKCK8xr6LRyc0
pmHXJmwgW2gcQQY/qmJCe2E4MB8kiphoPnQ+lq7DfHKf7c6E3YHSV41B7RFKDuvb
3NpnUUNmcDdMPhuQKJve6FocNHGB3tyJLYlAP4dk3oF79tFGiPa9QhCSwI2LssAs
eTX0Q+PPcNMZkdcrLCViurWRV+nPXMF7PSd6ynMDd2CSxI+pMqDF1dgFZuYEEobs
ZQKgCEvYU8Haz3lnGqstG12H5VwQXIAuqP4BFLl0mf2Lo6Uq2jabxOWrogZYN/KB
mTSOtbbrs3r8jEkb8Nun97d2T5LClwuGcYbGnJXYC5kJP9z8GhcT9eIgegZ56VBz
6I4cuCw0qrBK/vECwwldA6+W1D6+V0luUQ7b5H6k7YOJXkOQnGhC2kmMvy2XVJYg
l6hwkKPQQ12dg8qMha0ASPiXeMT4j9qYDajZb5YCb17wOJsVn1ODEPUTh8K5/Swz
RkLeyyNd/HzS0FmvNP4+v3eZztu/HXUUvfzvedK92MUuHbv3LzRotM6761x4Lzua
g6Y9y49kvszqxXmE+QbhQPxbKPJDj49S78qPE8tphlJS0RZGzUW/poSn5WMDQ3zi
LJcccq2Kzk2tA0kPxN28a4B0TQ91efLT+cSLp0i1DUSV80uBfNvxo2bN1G/8nOqu
SuiOi+As2L7ziLgjr9+N42MctymUQoKMGIk6yCDS7f0pitABoS4iVi99QVpPJ+PT
RVRzgkZk8UyDVTVMpx3d8/1oVHtD7XajAHoKGq7yo1sI0gIcFNz6hot4Y4oHS1Iw
LrQrlntBhFRn1E/5FGe+HvA2LooNpZGHxtPTJl96+iWSM4JaEQhKJ5UHocraPwyx
PVbMDQioIicyJM5j/acnB9iqwJBAp3Yr3X9mTbAIBgx8X6dm1EqxrnOOayVJEdgo
rLIpB9JU0F9Ua+8HGijuzzSayIeMa/FUaznRVblrQxIH1Vm1rBjwhODazmrg/ulr
CiSmV6uPD+LVJpE7NEjtyaF5w7toNs1rB7XDRCcV5TY7R1m2bt6x6WpFE3kkcrrr
EA58EJewtaqtI//BvrFfuPVFs1nz6mmHQuWvTAkgaK9gdE/XtriwHGG8ZU+JfSF7
ALoDpUCSr4/8ntdnLuRViP/TgAdTePqTmu0LdF66fdm6WfcUem2Vi+sBDmqOsf+D
rZqNgqjbmu82/2Z8HtIhFANZtsX0co1g1YemUPwFkC4Rm4PAhpDDR6L7WzOUhavl
9bNYd3lGB4j+e4ZXpoHzB1OTQ2AB+9umMntRmNsemoQ/Qc0d0NIlT4/DIPMq5KH1
3+jlMJ+PMWph2j83B6CiXGme4rN2sa7L5/7TlKKpsEhCaQfnMAXJXQ6lCJBA7LRh
0JlRUuEAdjLHowkHGlSPm+Dy/q70kLBW4HV+FgUmfhkNuqXnKp9e83nVh3RWfDjR
aKFT4SdAi70BwYsb3cyVVtLRIm0gplt8wbcsvpB9G09XQBtWrCv3mMJBr7AXmIt7
D3kAmGdQM01NqcPi+8qWxrrv39GHMB1lNtOD++Z40+d3IO2k29Adt8n6ETG/9x9E
boeY/w4xNdL/14vwQqoExQH+iBwxsI1Hk6PRcwxwqs4hDu6oMTRdRFeL7Hh2nQ58
o4kwT+9jrPyiggCecdviTAJ/HKAPmKh2rHh/rwATEOFDi7PLktxkIlzteGIWgY0f
pubCJ/gHo5ssJ5IxebA/udnT+0oenALeAFD/eWqxsI30qOmUh67lUzZn0lK93nQB
Lplpt0a8RKP7yM3SkaZswzqe3lt4gtd/u6MV1xY6xWOIwLOb2Kf9WNOJgk7N5Pts
bwnoUnLPPOcA4xI6KTACds1JUg5LmX1n8GmLsxOhEzTadxDHtU56UsleN15oS/tx
MjgYVoEy9JH8rO2+LKaNRN7vt4c+08dnpBZJoHXtMIUGRaqNH+Ri5/zA0Qp2Ik8S
6HZHiC3TuAAFiaukmxzVg8O1usWKPb9iJxfLgx83xg5C0YAVamkQYmD4VJo+Zu60
DPoYvXsZ5txp3JTAfvw0pxc1lBnteghtsD6HqcItOwpXDBHKtdJC+Etj4ScAWiig
E6087zF/FUyhSBr9X1nWu+sSWojXzq2oCGb4NRFLd88D3r+mHBViYeRSetnI+TM1
PFaPGj4JEuJ9zmkn8k18F/Bm25j31E6dcQvDvrPKatpswQF1oZQLaDNdybzXIzV9
G6CWySJ2zIe9MI/8aTPLpEZoBLkOuBkga4+65/FuGBurVh6z83ODDnyU1B9VZvqV
4sT3X/b612mcrS62GVwUkutnGs3YP3RcatxNPVPifuPcXouAxjgW/CJ+sehssU1o
FNH393XJiUyegr/BXJ2YS3J7ZsLJV2gHMMDfFpAYWADALmJC82RaWggpS8n/Huvd
W8+3uCi0AXeusXQRLa5UEI1n7wCxZnwzjRosRmTASxM4NojEFHDmjvhOn6mESMLT
oIhrIVwgE1AWiKlapm5bCBqeMwvs3cnxdmnxHQp/iXOAsnnb+bc1PDOPUBt2q8sX
nwl8bgNXiVPOwST4E0NaTz1+LcWu+0vmWDUibKuWsXFTkItuRZwUr22ms8Wh/lHF
bMWlGe+CAYYs7AKN1an3DAXjfbZcZ61576iBA0TwhXtjt7+Gi7DwGdfIBIcQv+Yf
jKRqZqaOHo0vDQ/VHl0hDbCtK3EPvM/X2YXbOKixfNATwmztECOM0fOIVGIdfq+u
vwxmHqaB/vZYMiGvYw4sGo4uQZ6mGfkIIfaoWg6aCCm4K8mpEsorirkCQqleTt7i
TZfwqYyK+IuSHzTE4I8NbkjNuA9vJ86lprvK40DfWH6Doc6XsOG0ZNIB9U30wlvZ
QlkiaLqHtJHpFeg4M/QLccmWZum3SDSVP3erHXu/NrQRr5U0p4YZn+txxF2GRfVO
gKMpnMEpLOpjIUH5NH/4c1mswzfgj0UNRHoKC56PW4aIcUKZVnacih6qmLBlmDul
WCNb7eStLmuml6FywdXZcAaGeXAZFm4xx263NzvaEPPt9paYbAV0/J+DKbT/V7Wr
NQ9/fvWiQ9N6Qebi5cy67436EH7y7f3hfFwz39ILk2aXX/SDuRoI7vFBqA2i2o42
SE+3316rw68o6ltHnFvCp0dGbkIJXPw03SxjIUi6fWpAmGkyPZdyDracqV1hlLPM
D/vHcNuI28EMHJM2+PsasBzzaeUrrqYrMsZ/zrsvJ0+PjNCcdDu48Q4ladZ+QGln
pPinP+N50xvhRHeAL9ahHYkivLam7qeoeN+tP48dgA04kjACJc6QC7JAPY8XfDMH
e0pSgjL6jZyr2OrJISMr2R00ujOAfRB5cSeonR4X7eTT2Ijlvbw8HdTi9GTZPKIR
X6AmP3wpwYMayp20INDWmEkSqoorlVlepqNWljnw2LzFPLP3DkZr2FTldMm9nXp1
lcIug/ktCkyj5MqSf7CE8tMDsTGuIJEQ4TOqEFtoQ7KwUpfVbOhETg8ZhYuDAtfL
fYqKgSjcbopX/vxoqqT8ZiEwhBcyZzLDqrYyAuOOmteViS/yLS3QRSXzw8U2A9tR
mTnTLoptz0l62Gs6LgvPdG8Lr/OKWyzqy2KquIq1CuPoH8F0I+gq9gmOaQ5NFMR+
5yQU6NMH9LgZP/39LqSSJuHTziTBxgDEXDksym1K0KnvNSQECqQh9wM0wHI3GcXM
VtB8ufhMMptFrxEgB5yKpJ7DKK+NvnSJMCKZ+L7IYnpAyRwSs8R/zP37Jsd0H/eL
oKu4sgLhG6mGf8HXz8AmNZKhGgyjKQJ/v3OjAl5KkCdXB27EPshGwraEVxVMi6Bm
OBnxrq2XsBrpoGa61CYs3GtiQqZkiJ3QIDwS4WsXgEa7s9TnFT3efrMt72Rn+b9W
K6QS7K8zh+vXwb738fc6Qj67Vls6zogM3vkqSVhiwKbodAm5gdiG2WVxYEvEMmhE
AuSl8a/fg99Dw1mFxFrFN7EqnHbObwBhC//5fLF3GOYtCK/mhKUphNfBKfLu3EAN
4ZRmILRiJDZsBxY5yPVvp+fYJtj8CpBn9YltnH26sK0gUH+wN9KrE+suqX8sh0CJ
WlUW1tYqmfjunU5WDQLV29Z+43xdfABx3VeTEMWBgX07jhnL3wbijbmTV0h2nKMd
IKK6jlCVGA5du1KXIx1KY7Se0pOjvS+mEAi+jlIkZXgIuRr3VcqUnbnNX4zaWI8W
S7+yhxMJXDwHiT8E/Czcf2krT3jYYF67YFiI+2wGw//HqpgnHpdvpmIAr2nxg1fM
lwG+3Q+8PgwMCYsD0I+nmq84+UVPD7RBcgnepRT8LQW67saAh5Qd1Ur0Atl/FOCA
ITkZPLvmo/zUzVE2R1c1kS8tMCtE4ZtwXW7M0yAeQg90CIDRSgHG4zX2KwuYFGru
fRh+vYMY7hTIUYYxreX63ZAgkL5V9e2tcLaXk2u1GE3GsHSUNQN/P/TZeG1GpPAm
g8BJn9usJM64gmLfsF3KTTSJRqzvRjAfV0pDXKmONigVoOM/NH/1aOiNYqMwp1ox
yMLG1Ff/AA+sttRc97BX5fs3NQ2m1ODqa9qxuqwjrG0Bfp+k//tVea7aqr5IZojB
kDNjbWnQLw3NLwOI0wTzhB1l1l9Tt2kjrK4ois22OVN/ygPCUkhDBLdvG4x0xiLG
DxDMkx8KR7CGZhgVqhyI4inwbobeEzs3OFs2L6QiOhax1llQtmv0tHj8AkpeaHLC
CNk43IZNt95KJRf3tyvXI4wFxEqyzwQDdQkQt6pxnXZnPXUepNkn5EkSSbGAGyxr
Fxh2xGe02q8hG/PZDrnDe1TfvKKpzjsXY/DyjGB0xAbhRVuTosucDmsTkCfNv0Wb
eAtufRDePPF+Ya6NiqgPdbCtUmuvPEUqvvbilNZXo8XdlYmZmhQPHf4TnMxmsHlN
oqvVXX3dmWcY/oGD8L1Yjq81Qy7ub/AqgLjhLJU2uSyAvlOErf8bQ3fvrJs2fwBR
IkcYRLdVmV86cu5N6CHw1X6zlbqJG+d76lZhFfxwo659QXj9awM84sdWzOk/by7g
8XKND68rwhma9lBuORKtBKhNG92OEnuER5Qdh5QzurmLYlzP/2oep9R94W23EcOL
7XWovR88K52edOPSbvwfvOjFNvxKhbiidccSH2dKKP2E1nW+x/xMytF3IniPEbzI
7MVQKrFEeV70Bh40uzGxV+8UGk+3HiXXZAikT4Tl0ZZR1n2L5JwJ55uDd4tY2eGA
08b07Pqvca2LKr/DxiuIQtCdP7hRaTfNjIz3sK7e5TJjTRErODOtABuYG73vrBEg
lLoHhcRmjzBv5wz1lCsvO+iSr89guAz7l44OehTwLw3YYdHQ81Ez8WA2t6cz61MN
g5tzHCFMxiWnLjuSQRirGUWQqXikBErVwaPOh/Owf/JOW/bRo8EYuolUW9lWUVro
pBfS+fmFEE7UQW6MKNAy/ySd1AyByJBJLmD9B4/e1DbM+8zi7D8xg1AGalQqgZVt
y+VRL5cvdhn2heFt61AyyXh13QMnpcExIiMU+kTQS+UuoxWsfQ+pjVj90NtlAcTi
uC/ZObIJ3MJDsQHv2loq+hF5zo/YmGJm8Aw0ETRYuIqnDu0tKCd4bs/WASf9Yb8b
xAb9y162VrBwi7E0Rh4jy3AHE98G75R9ICLjDBslZOUQ4xdArpSB/eXcN3yYwldt
QgdLx0SCyLg6CtZbIoHQKVGenU/yvckAvjUn3sqan7sQW5joO4GriAreH3Onl2fD
2NGMgI2XBG84YuGIsaCqvJ68+hS2dnGIZmayRBDjGNJ146yqaW1lUCiA7yR13pCr
X2dmcNaBdHnmOZ3liIx0v7EBgE+XD7XdbsHijLutn9bQvzokkOGkpexZkfXuw7tL
J9dj0qR9GQ3+3F35n5puJyTcjCDN7V4DtzpyrgS7nJO2JcV0crvBy2f9w6KI8q+h
p6eV63da1wcdSdGTHQcQ3QkcapSGoDC2eCa6XGFrXdX0R2xQzH1RTvdFK+52L1SR
RlFHx34rBigh40DrIn5QGW/54yWTEMlxuwBu4wqTEKCMIVAJEncQXLZn0QWaWM4T
vwHUJpxzl1WobFbhKZd00J+btpZ1JrDI6Nmn0OGpK4mGBJQ/cus9J/f+JNsQI/1M
k1lsHbyu2NUejFHitzjQIgP/2N0RUvlnV3YzCMR/7TaqAumJPW3NbbrkObxfw0sP
1dtjOMe/nFLJMpbGHf1BHnW+4S50hSuAvZ4utOIYtK9/25x34o+h5kRS9rdcTBWz
IVdCMrHDH7KVPe2OFnE6dt1tIaG31WCFYifeFaVKjtjKr9XypGnWK5mXLpUhStyM
TNHcdIy4/MEz3ZqqAvvGQKoOXcwFt+zDZPQSFjww6d/BATrLv+P66F16yKac75Cx
i9dnztSWDUrFdjJEHBpaWxFl+4CDxEZRYS+OLlMrIjyDgQUgawSSNnx7OOJmz2t8
ibJr2YiwVDl4SBcJJBaHre75IDvLM/FIi18thDgSY15nnkKiJ8oofRhDBIjRLJPi
3C1JOw1d+lFyujYDAmerPyIoOwPHan5IvlSY8Oamb2945IUzLwkLDVj+8eMBYw+g
qDnEWc465oMfbAeS2scw5emEGERws/xkedRHrUcINgPfJWEEX2jRTD2QbdJQdk/a
4AuTMUSXbSBlmyTn4f0v+ed3vNPuQHb6BZZTa2iWj5spAydxl3gQ+g6KKQzNK5rY
dw4Vd6umb2RReZLU1blkzO3Zrh1cZHljwzIWIxk//bGvPwfMKIWi2EYEAPOqwr0Z
uXDWSyYk2VcRhe8Tp6I9bIz5A6DTOA6mNaORw5NLQ5BbyogdN2Gnmt39XsAu3fts
J6cQRwPS+HfVP0YJ2TLF0jCjf/ixGq3n8WKJxvw9DPFNL2nqzTpusmDl3W6fyC7n
UYpqVCpkdTblAsP36BcWFCCGrpVWcm5FMhSrm/8zaty8lvw3I9ULU+gEGTAtAX4G
raZWfwLerzHu2EXoanzSnRh396ezZzj46ctyd3VIs/WHXSMgvjq7Qi5PT3veeNtA
XVe5Ou80jpEl3z3SzqoypRyGPoPyurjIpqWtKihiodFA42ebVU6/mYbVjjLcnje/
ZGLQIVEAtPJaYp2wg/HvazQvSKt0s9rFBQ+Cfgpyu+uGfBD08eK63SUMuCU4aitr
IJ8Pbv6SCElJUgdj7gNDuUu7nSx4v99piJOg4Zw7DdJDibEutkgb3gxBcy9xx02R
nI/FSY/Fc7WZAkGWMsEQOYHACzTLMY0B4sDPgX4164pSc5AmUasbl36exhKbq7+S
vMbPgGMxJ8Jm4IKKw3zyvDkcKVwRW+d0452XNnybsQ+v8p3Zy0hwMhHrcC5q/dET
Kz7ZFLjCQJAJYLhjUjYf/nITq9hoX0MVEp7pA5R8M+JXHO8YoU1YZ++kfNaPUXKO
EaeK/IirHaSl5L/Jsapib5DH7jqWMEx/YUyTmqERDayuT20P7TX2LcPuu7smVrbz
y7be9lE4lkP2FyQMIE+6lWhwEEyQ9+T9HFGAYcZnwDWEC8CW2gqvxIpBiBKmXg27
lFy95NZRgQS3C9ria9UAAl7CgL8jOEZYN6RF2YPtnL5rEwDKNPgIwvTwoXG7HcZx
sBsJ3/68B7QQKdV7amd9R5YQgSvzG3sisU8nK4P2L3oErMCPu+1O0oLCTuKSeMEx
4/2625C5MwviTpeBxEbdQIDPgRuuQfpWPcNB0xZMvse9dPilL+3DkwqWiM1NgcBb
EBDUs4k4OybzDRIiOatlfLi2qLOdsFG+mb4R5ymsxm9LyKuKZ7sekO9d8hZBmKkR
tRNAbBLtTL/wZWz8sgldbXhIRk1O9AUyculWV+1MvGuboy2DAHrUEBHtG/E5VDwq
K5aSH7XfYxY9RPjFtYNiLYO0IOd/8/hsqNCwY1OrEgNzmSqrqXH+4V7618566RK5
9QiEY0uYN1M/b3b7Tah4Z9PI/miKsHt4hCLcMSPsIPk0h6RPTirw+LQ/+6tzRgOA
j3+4ibno5MmCJM9qcQwVvzV+JEZCyrZ+1AD98Vrp/n/CR8AuuJAhwHnnJCmZoSbp
I668BU13pjeFTREL8sqU6o+S6i3W395FYozyl8kPp0z1GzIvkMUCUQWl98dqMFZo
H87IyyRGo6HEqg5kqknNbzh4rjLWptoj2ZiX6q/sa50e/aJD4UIzlC/7kGlgzrxV
JdLYDk4O/OTW22J0mL+th/szBj0gyWUIaV4VcVUiReUm1tGj2RP5e1fOXBTv8n/d
oiEeVJUrRe9gcmn3vYb8KSQcdhXv2gkzjno+9cpqB+G/KAGdF2YX3fipR6uWrZe0
V1unp5wy+mnbCUCHa08n6BCoVJVHCwJaHxZ0rDFYw+aKNf1c0O8OxO94TaHdMn/m
Q+jW0cArSpuRLoXQyMeMa61EVUZVtWhCDMz35XP6rzocEX4p/sIgmr5tbOG9hV4h
yhJS2WI5s/NswebP0tJ1tsuzJd7Y0+Q8pOqv2kmApLfX/zctPCyXwoldaahKMQhX
YbMF7fvIU/kjxkqWDI5FZST7oe/Q8IAFGuyKXG+8iKmaLy6CQ1n0BlPlXW8i7QHI
QjAm8wIELF1+2YorVTQuVmHp84wf8YwvQgcdNifSSm81qMk3BuMvpSbffbHW1jEl
QFIdwtHQPp54Dqj6nIo9Mnkfoy5eKd+WX+Z+K6xZjkvnMV/jwqJo32DYEiF4pXa2
RJl4UPg/slfnfersQm562F84R7FshsjfGJ0ZEFZB4eFZrVyC0NieIP6Uc3AmWqn7
JQu/ydqkjbGDseg2p7zCwwYN2vXIq4bb/SZNVjhKJoazY+A1RAzRAscgaHrzKsUA
MYHL/3yC49DhKQQ3P6AjSZ2HL/yN0x5q8qJt3tA6MnLTqdQViUyI4MS/z/e9ENjz
xuXjUi1x+jnGzSvGJNHus1sH8LKKGgY8ITRXG6o/7zbVLOqvuXzWoYRb3+US/KqN
qoWGMZ5JLmZMkFdI5w9WDCS4Spzy3rS4brbNdaaOj7VXZ1xmSa93D7XqyXOVm8QY
GcKmr49p3Hd/47Ym6ysNDKCL1UdpxD/joAk9oLxtfC0FbpC5qMTuuGFvh+bGZ70V
geORkwnJ+dxnVWvyuoiyUWQ4/hFVvtRhuM+7JuHjV4uQ/4uktQTcUhHs3PglzSx8
ITS6cdpSIA+VFvLD9ml1GGyUW+XN7HZeuwBjhLMvvEbgXWNLufB/RtGyT5HtVxWb
AKoKfdBKM2vP7Xpa7T3CFoYRS+fIKW6r4INHxA+Yz/eXsGkQMGpmKHHWZuLolcxT
sgkwzglGorZTIk2WWO3yl0qO9FHS7RhtfI2G+l9X+gOGR+lll++4IE/zW78+fU++
bthw++GPYXWSYOhyIwnjZ1NWjNZUw5szRxy3n3xkpbZZkHJxGTFk1x0JzTN2Wv+E
7XM7fSgHWs7pNYqjeox97TmXfKV51Hkw6ap1CgEFf0AS+TeU5WD/pdhWMBXTXR6O
Nmv//Na9ilWE0ywML4VlFf7gnIr7S7mRDDR/MSlUWy7unjgPNJ0x/Jmk/3Bihm4h
NBx1PMVWQJoA1OyOoobj3Myeo2N6QlR9wSIAn6ONwoC0k8TRjTIIqdSSMtVveHC4
98WADCuOJvjhzzeSKrl/S2zRPFNje/IuHfg7ejOTlDHBW/Qdjk/LkaQuLrp0y7hy
TKE1f++t/oX2OlSKmKgc/Kc3mor/CVJP6xtNFZGLoB44mhq5hvl8Br0KD2U7TDct
ulCHY1+mn6wlMrEIFMAQ6dG5Bo4AsdwxaFB5q0rIVfMualCuAsrqPJ24RVyraTZN
KN8K+ImU/EffkGRmSp8CljuiwNi8myW/wKvGlR55lMOt54IsvwlsqtwhKjyKNkGu
IIiUMQgL2s0W6YL2rSIZS8L5Fb8YhoJNOhIt+8iI/fYpqnsqysPitfwoJJXLD0nS
De0dsHK2W4J84COg+X3rmLOPJHByKcwb4jc8WHL5lo1EjQvqMxTpNt9+dJC9exZw
MrZwgxiQJvaCRxclRnTdkrmm3vHbWo7g3SEU01idx/P2KfcUxWat1X0QoN4VIqN3
DPTXbgzANV4CUsNKq38xsvAopPqO0/NzpaXY+F1R8gnSK0eWRetRAji6KBChyHEE
qBaNfkGcSjUD34uCytYex71tnerqgBhHXP83WSm/WRwFTrK1Hji0xKmPdplv5o0z
7Z0BGylbCHbfsllA2MogL0QIjFnEfwzBjl1Ap5jxjaXuauuYyJVR+8hLuYlsIVfi
6A/8c8XnuJEEYjY04cmsw/EENRwrcrBqHMB8ntYwfBqlhTFZ3lKCcGH2uUbBcdAb
7NiItlTbwTT0kAaDSX5PV7gzLL45R8Mv4bslcPTkBDJqvMrerhwOlU3wlqpX1/Xr
+rapOfaCZOwRn2b+Y6+mG3pG8fyiBW3t5brIB016M2X6HyqezZoDiKYcGsLqH6B7
990KFm22WaFcAqRJbboQxDW94soAxI1rbD04zEsNjv21Q+KaQHO9VX1KZlkaEOWa
dFjalMeD6fnPHZtFTeYRYiLwlvBNlCjcknSziOXfLM0baGmzJe3H1nmPF3yP+uwG
tVa13ojbahsN852Hvx5uK5jjkxskQTsDJd5Ccg/bn/IaCgb0rTyPqVFSu+Cuz9X6
o1KVZsDCAr0Vi8x1Kqcf+ivutOJwWPlrZiLBhyS5+8KXZfl5mLVH4RTOv1m2zY7O
Ite4MZ/8lrG+UuDtxgiwGB+HvrrKvtpKkc9bW5m8yLdi39GPCBH4vXUEZQIAeBt2
Zff3MtdZURxHGyaSn+q7rge7Rtqbj/kZHRw3Poxr46Vr8Nofnr9e8hw5MTOIEAhO
8F3txdn7sSEnBrrBHVAG0v54KFcgG6iOrED11ehhsV+NAzam5Hmnm4rbg9JrPFMM
PEzcF3CkrlTJYo5y87j/9vZ67bDrJmihFSnUsKW8qqVl8sXyL1runT4V4TtOHe4m
ZKVMxZx8okOLbqRi+Co3u2ol2HzB6clMCUvfQioS+lGUh2dXJrvpCqIo23X7oiRf
a9FiA1RFvlDJQEIoBwF6Vv5+UB5YryI8GX4EiG1DkaLgkxFyWwoapNyA1IjktPaj
S+ea47Go8cOBHf6ek18LA9SsHSMmiJxbVL0QhbUIHBgu/xlu13RAuESlSoivw86K
pAAao2a3PNnWI0ZJ2qWDVenG0//Svzs/lybJGxjuSSnFhTUunmXlFK5zKfnuMyV5
ilXY2EQcM5PMYBBqOL5vm1R9fMOJGb4303TlfAZqOZEF9i7WdLzJZeqX+xmvEHwP
Oqn4DNzj7AcUPmyIYQ3XSe5uD8v5Ch9zj17m/a3Gux7Mj2KWVM+LhfmVckE8gF8N
4XdMGXal9U025u4Bf/ixBsytJjrOJZ6vj+KyqLdRpuc5YZHVtSHOPnzbnCaNiTCA
pTnXRucE55N0NhN0FbJ5jNawTwv5hQSFJJJfeu9p7RAgWzJUUXHC1yzdyfuDdsJ0
Sx6cTVI2wcfsOxgcn7BtX97asKRUFfp5HQwQgzen6IXc8SuF6QiVyJ6Fj0HmLuS9
J4bEzbOQxONCfD0ZLiy0pxPIFmzOWE+k7+IWuWqzM7qUFuEbkujybkETpNG5mdll
dzsl191k7UTHScU5YKkXeCNkZIJdylqskVha4h1DcqlcdEGX8h5tlUE6wabtwwX8
nX604yB9NSseGhEy7z4bdevNJXcKfW85ChH5IKPPVTeTXCegatqSvdFWhWX3GyIi
KSUKF6tGXF/SbEJiC17E4TVQ5vd/MUUhiDw3WXKG1s1u1In+zal3XaRbZOrWPR5D
X75OX5F02ABIwEg+2ZiDYwimysjaj+Ka6LaR/0DJxNFiRrpN3gAOK4oPdn93Nip5
douur21yQtkFV2rDGDO2bx3YAHeXeRwOmVGbkZTvmpoTSGZvf5qXdRtoyqwc2aJJ
Y1jQXH9RfDlFpZ2dXmejECgeeTgogMuQvmJhpUegJJRC+P7k/awMbzzphaJ1a5yz
IKTkxFiZhAD0qd47vX2BuNspD/rvLtzyyL6MSrZFVJJ/qL8KZscxVGBc6+FepwD/
fRHA/i1ywEhHiq8tY+rt7yh52O2k+0iy4ukwjHktNKUr2KJFq001iR1C3Id7mw8t
xqUXIfdatX4jmcH6gtjcCIvaUxdwXJ9qmxNOBdLD3sTeOvIuvAshxahgSvrb+iD/
BP/U2B2nwPBzqMPbRx8cSpOlFKaQJLuH2bRySqc6lfPqpJJ51E7AuQf9k6+Qb/d7
t9z4PV4nEUzVFqN376SeHQ41cX9l972xKR76s+c648NIq+/Y+/bl40tLTatMULaU
7E/gZDo5ZIbJZAwcQpRLe0T+GYLBvnxgjBKNXyHe82ySgJBg18RViq3SWWXXJfWh
hzlkvkY8WtPDugCQ7qk5OtyOziOBaX0gVGVty3b9GASzNri1WsGfARzt6h8/u3S2
VMwINPzIfiTWaKsiLH4KEyJDkhii0s3VDys4XQOTyCqOSuzHPyubq8HXR6e7mQ93
fLvdDXcRp5kamNjsO8gi+C4yjyPXB9hQr3QPvrtPY+kVnAWTq+4dDSTxT14UgF2+
C4TNyE4wWOtQIBrMPcmlF1DvOayWS8kLvjd7oSCdzWK7t9NKTUUeO81Lwum8t711
gdphK0M+j0uoHuIAWQwl6J5WV5XPnzc0F1gVKB8wOKy61WVReOIWT+3t2VrphTME
jdQlw1fhWcDEV5deO9xJNmPg14rT/PxB3rhz5EGqCwkRCaUrx9vKZiUQ3O/MBvWe
m3UzNVS0rn/l51Ye0VQPYfhbNlHOuhJ/+uBYLxgkzk0fcGKR4TPD+ex6Bfz/JSgD
WnjlCHfD4XWzkYNvrZp8uC0Ig1q/goJWMrftTRyHb8rIGRLaRlZ/1ECKL/m3llDW
P7imnpkF1grYYayCJ48GNe63ym7N6tWNSjpUvpgPAU8U8P40eKR277G7C2sLg1vM
gb7BW8o8xsgsJlNwchv0Wd7edyDIXvJSyA0R3NmCuFxzObAM6D2nmdhsG6qJeuTe
yBb05U4seshH0eOYuhq529hKuJVkhlHf5C+wipB/jtYgSyZik84PBZALvFk528Kf
54iCF74hSrl8lv7w+gPyDBjonCcQiVdn6vse+phxOXweY0stpY4Uat4A2sjbWGRS
sMK/oZDlsRt9nBPx5/803FOYH6333bZw31L70WwrbBnDbySdTi+u1HFUfTJZWSaU
OUJIZSIzjj83gqgX9zGzKRjDt4RPnes5D8+62bdXIzRX2fz6cUP7P+tTx4oQL+oo
O8WMfiIckL471WCr+BGUWXl0Ko/DJp1C9uU4xWADtxTAHhRJhXiJMIHshScYi6q8
2Yt8qoqZNY4XfGQfg1da4p4wEibZ0wu4ZUoLOEnY3QE1paJXJnld9QodL3FT8bOR
XSpgVz08Gw/+PItmqXhdB2IW6R+pbvQYvSf0J3SrukFAPxGP1jtS6z5sDmQMT6xf
voCnKtsBpYXFcLp0MmbfaINSBUjFDpFlbobLYCCLiVPYFS/HJv705iRjwdJd+O7l
u/gJKXJG3chP5JoF2DjFvPNF0Qh6ujFDANbq/AJBqWUxwQsMzUWwc8LuUech+acD
owN7y/QM8mwxePcpTWy/kaFpSGsmPeOf8On364m7UeXRiSx/KkXrH8T+ceq6ATk3
AzcfTqarHUBlvZMPurxWwHrvQA1pBTTCMRqeWlxsxhRB66VtjPZCGObIptSlNBBO
W1CSVg5vjQzVY/CgZD9VI+Lu+n8xaXaRS4QsxI2K0KHSzT1ATbOGcXz5+8SIJUEL
F/tEH/3P3ZKiPAZrH9FsJPE4azjdmmdkQ/AtklbGFZDt7ocHegjlNIrQq/lp9Dza
LqKKt3t24KNortMYn1/uJCFp5+3Z9OXb3NjHm9IO4bieokPAONwVFUqBNqZ43HCv
j/+lW6P4bVciDBTny+EUphBTx2kX1GGkLFfI/SvmjxMOhmsvtTBVHPDQ7yVh72kC
+oi3BlbaGEl+P6Qx+lfHKvz0owOodFhFcMP+mc2ioY0gxUMTm5Qj3PrnTbgR/BhM
6y61rAwT2cSZOSqEx5m+NYJXr1r0Cf+Y8N6QTLqoYMaeRM4a0wS9CG6YaKcH3Pk6
sh8uyRjf1GqhCzQ/Jp1pn6pPv9CYq4v8IkBDblNRWlMvimsiWqhowfulQjlMcxfZ
ct/7EVXNXi18S05ID3FkMIKWzm+RYGVwDJDG4mnpHZrvr/kW0aQMqgyMhruqxE9Q
qAAoukp8DNIHfVxcONknMyzRw0vDqAQMIPsijRuymuDXNiN+95p0sdOi48ONx9eu
L3ECNlO9TwLbOWlxZo2gyQjVMjv17kOSGqwtfWROttRHCzwhM3PpSQ1Cjz3eLZAa
loSACq1+zqEg2Pv4QJ2iuDR9vmQ3Of+IN6Xz8XxBPvYNiTp2OmHQHZbr4s8YPooH
HhoApqNwH2s8wcq42BD85IYkQuQ83Xs2bAFhgr8VYPEIenMcBd5FbA1bfCEzVbQL
+0b8fMw36hULTsMESbuV5CJtzKaIC07CQKpt71tU6i5zI+xDOljMG/CINqxL4G5P
+Nrlz+Eo+1ERmbbng8Y6qUjVfuyH0+Tt70/GeGvuMes7Q+J+qCLpDg3HTTV0CNYk
JYrbZERRtIT9GqibLh8wLn7tWezD70l9sClQ370A8IfmaqOuVKIZpotIILHmobFz
sMeypirutALESfkpY78Ey0ydL9EziAo3YKYCVfTBresX+GVpp82QZ8kfnBf/SKSY
z0sCW8fw5N3BVwJo+F3QFDP8I4hWvHSPszbKsNyF/DCIfDNDQqD3ZyQF7KsO6tbB
/LORtHdafQ5VIehtHDR7iiW32M21LK1WkPK8cr8LASjke8BNZDjfZas0uUf18Iix
QI5Yzmt3G55oFq+Sj1HV/ZVcoyVttRmmRsKVlnxomFbYEnzH6WvKXSM2DOpWq170
seW3J9JTPAJ9Z4OBvSVPdQ9CA06k+wuxIb2E7HZOuFrLImR0UAyTvD0v5ctCszQj
hnk9PpB78y5kYPMc6V8/mHyfnBA+dimUXsfYOUtklGVAOKleWCK+Lde9ASv+AJrF
q/Tkf23MLgdmsrHFzsA58dXrtiatzrdAEhxsvlJoWOHfEofFEQF0hffntm7FydTI
eSIVv2VegJqrwlfHKG4K1o46+ZidrmbB4yf5sooaPoY51meVOqRheNimz41uLRaZ
qsJGEiI+ftRyibWvuQToEBASD/rLSrb8/Hy9EWXwunb9q0Q9lmUf9wuZ51H/cblt
xvOKQtsMJQZApjFB01KlDvTtvSTuqx/kdm0Q6YVjsq1IF2nF5EoDbHMfkKEcvvOS
Uwg1xYfc9cIcCbMMSaXb7kI5fpTiyp4SoOlJK00p3lIczk8GUv+dQaZY4pZDF0RV
SAcW3vhN1Kb3K2q1v+QshhwVd5ovvcSTXj491BOc1Taa0ihneo9fys4t3OcEGuj0
+nSG1BtWGeYAKxRCuFvKy2BMszpYOhm46hLr74OiDZVuGaKIRWakzMGSK30vcNhx
SkC7aGTcIC3/yfJMoSIjyH+udUDUE32K25IEzrKWQAUszuGF1wPKfRxDd2wj2Mci
2ECR07/SLhpXqaENFF8ZO/mFzi4btGwz0YIJW6/vhZQEe7nstZy1yK4fB1RNqMba
l1sgrg7sxUlbF0Pz49AAYnVcX/qvtI0fQFi594rG+p93P/tnBdAZOheR7/FwfN5s
6z0zmKsb5IhkfWAnjc5YXmWSxXtRtbAa7Um0Bm5reTeCn1q21Boh6Ik0Zq3XML48
vZBduvJP4lbSZ4nhUPgfHE2o1cXfN2i6O8bBNRzwgndbOMVFDWqFVuVjsIQrC3wu
Bmrac/zdvBwDfDvIxJKU9ldnfAeOO94fzpdOzLGi6+ZWNCayQB23tWBYTsDFL213
Slng84sGNjrIDqbbSkJA/DkwpwBEEw2BG3FewygUa5Niry+ui/vGQGDvewF1ZEGD
/NlhGSW8jYfBd843uIGoJCa1U0FksJn1ddBJevceRDNtwldbNYQnBMfQ3yZpa84R
GOBCiXVXMwSN21gXvUNGF54cc+oDEcR73ruTPJM7l095rqq7R1a56Mg28gn61JgQ
BRV9E+VwIxrD8ZCEujfkC5eZWx8AXRyS4nZDckuzfi+jMOG5rtdk5n2Jb48S90sF
IMZc2JDTC1semTX/GpUdSVg5YaOLFAZwMQ+9typM1u/sgjXxdm0/Azync2n7Uhro
QEZBopEIhlX8pVhrnnZgvCCFv2P82Qbk7aztBFq4Lqk0PsviL0sbaY3OUrg8TZ/Y
ixFUoKIG32/0djBzMWgPMuPkqYiY2cyAW43h4wlpx+z8zWFuxmcfq4CMKO412FFK
VhEQDGLO0qagStPnldQ2TdT071pg2dGrGeKOC6W4cBxF5qKQPYEyNUyLzSqSEQUv
oG76ekC83Hh6flnULO7Va5V61w5gYJlGG6YjY5Pkma6dct6qPwEhqfb23LkGKx7+
s41wwVQcgAEEShjdiBQyKk5XB91G7RWT1sqRF0pzMQvQHIPjLGe2PK5Bn9ox+/DA
+reo5EDp/CUEMrrOdJWM4qA8ewsWxHvTwqkOlK3TO9misSrTXehC15iWYlmwNZYe
hiPHmsgEzXRkWhZEaLJrQ6VoHVOMMCrnba+edTypV7Sz5ILho5GxTsXH6Jkxs4M4
6WC9Orj/+7dCyOuePC6lRZf8X/DqAYa8IHrD+5Jlu83YnO3j2Zh/7Sfol6aH5QBJ
JU8dCUnOWCEF0DRWahIq5uG6clcOa3pXNIp2MSmDV+/UZsN8Cta+0FJlw8s/B2AS
7+P0ybypIfimqc+BUkbEp1PtQZySMB96kkZjX5UMvgHfWPVa/Y/R04f2juMR4HJt
B5fD6fUKalekNX8BF9Rd2b4pGryKdPkHExFPmn/y73YVmE8/GrFfmfI8TMr8FodU
ABeu4Sli5qBi90ESSERbypBNOUL++EmqqPHKBBiv4WVscRpbi/Qvz0Fl6qc/hSNa
XAG4ARx8Qvcb8hDTzXt0EDjVk350VSnJjXgO9yHAB/r7mvj3fp4J7eQz47wZPIB1
I/iajOAaCZejYY0t/r9xXyhTDF2hZkbn1zpONbC3ZMKXpoAoGbwTIQrW2H9EScAW
AGiNL7BV/cVHb/dhg1A0Bd+9PVE+tZYsV+MxVSZEfK+wXonRXNl12iz/ZN9mug82
BEYKH5b/xQwObF6d/rrVpSy5Q29dsLqzyq+LdoznqaRgzI3vDQ6k2RkN8SDl9TaH
Qy6xV9V2zYFgc74Vlkbjx/rV2T/DiEXKBfDldH1N4DGuPl75ANmlsa6jHY9h7Ko+
WWC/LuDRcGlX1pORng6a6I0DpHtU0zd2DpVIaE1whZLDNWTIhMsuYv9hTJnK4lF1
M+fyITjMSCp9mTdUVPq4Rs8gM8Of6PAgn8MP82k5QHopn2y+WWwlzLgLqvtchO4d
q/KPzVwZPlRbtw8ZHWk8QGgOEjHLzTrWoifCKPky7r+D0TKraY57SlGJLtP6dfmx
cC9WLolY0wWo4IUXjpB8fdGwXfd+z7uxsTniKh2SrCm1xFSsMEqVrgt6/PffHM1K
W9XPNsCOn+5v/cIsLv5yLZTYxY3ggonTUItSlckQk6JmMDTYlYL0xtcJCcxgNImM
SyvzRrKm22KgTZE1da0wvyPP2gU5nN0gpff2fssm7B+kGrm5CpNyHxOW9SXsuxDV
OPYj7rKYPpipPQP1o1013h+H0VdFk6EC1q5dCZS2S+ZR7wIZ/ODrvscavbw4Z4kn
mZbvHMEHf4tg1RNm4l7fPvVLABsY0DUPfNbVUOmm8PyunZN4z8a4AxxLBOwrk2q4
i62p2Vp1FcO02w21/T6lEPshYrDduPd7FYQBB+AyqRe/faFQak8WtyJ8mPlhiY/o
63bt4TrhT+7tW7EYDIHGt3z9NdkpqRHdu0f3/m7o0YskbU6kQ03WwrEQxUN9FCT4
iqVONEx5MlVqKUi3vqiQpZNS2yky9OKq66ofaBxay8DwVO8+T7rThSp33n9cWpgJ
u9+cvxXo8Ulldqh7dhPtbDRCD//3SWO30lSN6svuMLdGIF1brwrYCNkDI09xn7M1
a6He7jZ3G9jY+dvWNCA6Hn97oCIA1PjTHPWdHf9JLP1Gxpc15U4QfPKgL+bL+2yh
9kDmq7D4mxRhI4q9Lze1KP6s9Q2PLM+jPGgquWBXWhclgp6vQXfqNo1GV4hqLNMQ
4wqx1mHozOcTIk4Tu0va1csXgoW1TiVTZu9Y2roi/HjcIz3VRhxpSNNpNVCvLrWC
oYOJNGy2MTaTSzG9+SxxyWxccZJZIZ28AQG53gOr7MICCEleCTzTgiKW8WxW9Rkm
vvfQA+1xuNG43VoyQjIZoEWVW5miHwfd2r+0FGwJB3fP37sny5JD8KBC0uDSqel+
qM4WVixjkJUGhpDLBtJ+dWXtfgyNOOm6L3dnT3ELwPJLusBxGxN7qiZjwXn0H8lm
CT4IpoA2c6voyf98FV1KlQPNmuLpd2diK2vDm87w3tjvXjVyPcxhrElp963S4MbB
rTiBRPuBnQERAfS/08CwWkpWd/+o/u7Ggcz/hHzimG4Jmuh9uteHVyp/TWY52hWk
+5vs26gM8a7qCm7i7WXTADaX2uNeIHTLrBf3MykG31KBHa/oZt/xHWm1yc52HLhP
nAWtDGZw6RUkZazLA3ZSi7yWAqRQv/Cmd2K69F4dwpzA8xOKRCp+KAVcgPhWt2t5
1bG3+/5Ubuc6YDHU9dDlH94h3h1RZt0V+CRT+0tnxtzvNr3QgWevINjwCfNjuUqY
Mnml2vm2dRfWgaOPU+yc6WeuOkUOK7Qk3YuU67CWdwfe6mwAmNYtq1oXcVXC7tIf
IVkt3w/rCqZbn++CH1DQ8/SueB/ppfYIzSrzaknpWfvna7GzLosKzOkU9sw2Rldp
X6m5rJNZs3zPZyRnhIV8wz8Q9L2F7ZF0Ghqa7KoloEtYVWGNkoznMZMHwXuGSnXp
VC3mCZjwrK8JxNKarOhCG6Ok3I0QAcCQEVkUS2UoHYeLcQ30Jgeuqw5HDtToUfyz
NOvdG5tWBjgLFukcepC+J/Gike1I+4tXGwSHvA4Qn8bMSbkvidWiXujH0BC7L+hr
jRf7dhYHy4pyyMAodOyx4cqRGeqZeHn1xO2BvePbp6DRCfkLGC2SPbcNNwmquvYn
e8kmRh2UIn9XlyEKnsVjALBUsa3vsmQS/Z6L5DZ/8k6gzGMEAnkF23pu+uA54lQK
KBn0rKElmLOz2tCyo25JCHkz5N70ShHeYOHKQuQV2kB978wk3Mkl6D14+vn7IPt1
5A3VzWA81fqEfuTNByHG0+uqaNHvsZzhiwxXDQHdptiB3Z32YWZQkF43IBWWdEvt
FCNdWYtaNzmlNmzZy0IjNK8wtDO2Ku1wVmNtwO+dRLFpH8AbkpSgUDikpISquu+9
VvxpZSKklPf918YblTQTPhKkFgMqBkbphAd56wJFYnAQ+xp/zGKSdAJ3uWqSCc85
qNjuwfVJEPyqVhSJ7FjURnJ1O//zVWRCnUdWxHdNE+UWLY+Q04wd0pi7vTCSS/e5
PTHxZpCln1QrP20oASty0BQKXvQMc2RudOZZDBovz4fazE2w4mZgOJMzkp2Zok34
ZzwIrtn/IkLXk4pdxo2XXyI6h5TqlrIqkhiY62AyW9N6FRfqaV4n6gGg+tUEsVkD
qhmUQm7iyhO8/nJn1sjirwZJi4pswMxjKh+duW+oj23A+Chg1QgFSW2RlRn4YTUo
KXNAZMNcN4we3SXvl3+xt+BVJYiD6tYJE5rwPvakCH4mEm3Chae969nme8Qsibbv
0JUouSMPxyN07vC+DmrwuaGOgKt/czFRitwSB0NiC7U9aSUUfXt2h2dth7p5/x/w
yx6GF44Ceo203fVd6rKXcrvZS49f9EKG1sQsOyzh6TbYsGZFiKUvK4+tTZWVmn3f
SoczDRyg/8SMWYI6WsA9GejRIAO/2ICeTmFYtYoHPNcN/eQzBzMlzJhc1Qizve0S
0+WkoNNplAVABXGZoNGrN3AsTYxaRtfVTSfhk2szxIs2RkWbiph5vd/UHjxgv3mZ
g2qV9f5FKItRGgMURS6VyXGPCgmDeJmwBECf/6UcycDAXmQ4nfSXzlibitf2iR4N
I4v1DRKzMrukPsfddNVjH8z0ll53wXlISbxqYkIbDT8i84XJxXMg1eJcso7hF87R
SQXgbN8+Xab6OrFjC4ZOKyxnRtCowEV4pGjTjNv8v9V3Dkux+stJNy06c8AwCpUP
zrWWQr3+lviZqS4uCHQZXXL4zcY9QUEBFRP/3Wl2IXiE4fQPXc6C6NDkmd+2cwqr
Lnr5poy9/WoGND2ojuBPiiuQEdf/KxQII/oIfvfj0vqFWdxF0xlGf3H7eWVcQcXf
6rq8NI+dEk0C80TQN9ejijDsCAEJp/riN+4yUsJ1TTQyB0rxybGhz2S3DJJbXZGc
d6p9P67v+rL5AvmisFHh1tQVrE+oGBZCKpv95YK2Ne0SS1rY+M3fdm2fNUJrr8dK
u5U6dMLh1TUJy4fz5DEi4r+642pyEbXHq4dfSbJdKcR5m4KcDLw+5X1krQGqIC3z
G5UaX36KoP1sd472dh4YRsj8ocWfRDYYA9OBtIG8cn9hemcuwIuKqNA9oMDKzRMB
o8RoHZJEk1YNAVntVXZoXkhcM4selQs3aIE94E3UY/ODawVTT5kA25xQ7wOHP3hE
OiQ2P3kPWB5v8ITIc3vxnzvwDplv2iSYYsvUT8Z+FfpN+e1+wl+QC5B5NJ5i7yCd
azDa3oANNAdfkda7btbIzkcxxDBSqNsNqQ/ZfUmkBYYbsvIlFdvNihMJalRcaB2G
xoGAxIwHRp/YtIqsuWauv3ySgXfuelSxE1vIXfGgQGILLTiGvOmAi/G6ctF4kFMt
FpgBbL+87HxPcC1lEKtHk+00pImdMyt/y2lcQW82vdrw/MICxmvVxSNEnlYeXKZO
w1TWuLOgOZHPEYU3lPup0KkVCAUNm1ExeGS7J9kxCrC/SyQZTOXpY2f1jCjyFTLm
dk3+lbIeIE+ylKnDPduh0XvQBPvRueN+TtfE/uoa3hPvlsHQY1pO9zlupkJBTeKI
RV+865OVUppC6J2yYCeoJbBOTr20BLFgobYBMNeHwEbj4jmwg1N5aE3v7uSi3jz5
x/QhR7lVupshH+1Yc29fSqUfFf3BmNNO0k6kdBuKWYTlzky6XbVL6PR7fLHS4Hsk
Gc1EuxwR3UvQT7c7rYIURsOjKFslgBPtyZWIhA9NiYBHuPVPGrT1CWQEvmUoTtv2
zjxL8dPjfhsQbB/VSBCSo4ou6rsAzPKh8Ev5NHiIQgFA8p1478DoKZlHGyxrDiJw
nQz2dI0xc8i0G339Ylp3qwBPkkOVloWX5wR4OBVTU33+mda5CmbIWC16I+IRMoCF
dCz5MHf6MOmf5/yM7ILGtrn6niMmzYToTb+NIikwvQHO2wgUhvhDd5iEmT4mQWqx
KHe7VuauEOenMrSvfSrPQ9tqOCwjxjPVasHSSI5ryKRYdEEEk5BZOFbvhphAIfQ+
CzbWX5LuN2ZsuLi4v8w1s7w5swAjQUHKdL6F5/yFOfd2ewSXs/T+UqZsyr43TbnL
H0FRMyGoRHhz4WUSYvvs/eOBrr7DU3rvo0gDW/KKZxbZfL3X2KOfBIiphoFNF8Vg
+pOJyoEU63wnqWcWbPx2fZ31k1hdjOfldP+BHXBKv2O6dwCRCdo1CBHJl06FSgTn
MntdeM+x3e/r7y8g8HN9xP5hwzfU5NzSFkS4MAhWhLZ6CfeZCFg2skpt/3EuuUqU
f+0O40JKdEgKkfEWAO6yD8HLRW1z+DFhNyFniunbRaF69//L+T+4+8SGiaHysN49
lsoTbzD9L019H4XmN/vD2KsxyH/hP4qXYM8WFm7qtwcRCqkyAE4hnTUdhnCfuQl9
zWRc0Fq7/kTMlNyH7zDqV9zrYN/ccd1djzeDcrvQ2EyMNWM0ShTPi4Kzhw3oc5eb
JWO1HkWGi0uWCMoBT5f1KqfZRvYjQrAbsagyiJBHgkEWFjg6QxmlrNoMduEX+utk
lvdPzHBSjOI41nu+pVP4trK4hAfi2Vlp0PtCOCrTMJyrcnKl6RyM4yPgXjNxGC8y
ApqbbZmhXN1IIRw7jkXYiyBKmpq2d7ee4MgyUBIAHrbj7g55hHRvyS/34voZKlb6
b0pg+4CcTRX9tWKV7F/5tGVSVE7lSTm863JdHH/NBmWHX67Rgbz+9GZacuyTkhJR
MmwJTHkJnjBl1oCMkEo/ljxtIxiZMn3lBtqrm4fZNmkAKjt44AQX7cXIYW+gqsYU
I0Rj/QYLTJaswAqmH7Lw6bRT1R3Xkb26ad6tBLMMZnht2djZtuggzkpoLoIUBban
0zkGe2WoaJEqPhwo2u299PidbNALA2+gPORDpojOWuWYZxWDXfSrZ4qWoEdlC4mZ
rdH6v9IIVUTBmZeq0i7wgTIGjDIf627LCuJcsCWfxM/3cpx/wDcvCzmk/OZF2vn/
3kckWsG3VUGLi2fSkS/3SZKH+o2ZaHE3Up991hfJ1wotlrmeVo48Wnv35wTEe/pz
NXzikR2bGIzjoKpIXPBk/wqPi7Murj9FCGAiJ1RWiHfd8muTERQuta9GbKRMERo9
wsts6iRVhpZoy+Q4SMUMfI2SFymLqP0mVJpGHd4RIpdqNv/JStrxFn4Zt8dI9o+L
nASBy/dsTW7XFHm6grdqSVfG7tw3hLgVu4f36osGogsuSRPsXNP+ecsvhDeFk5Lj
GM+9XFd4zgayL8+Tnlztalmr1iVuWf27qyYV1ky6AxM+2w0exbvn2fy+wBYidZ13
NneJf+y2yDes3B1WlJ9mzBiTzMo/IeixGUC2dYZdqNxu31FT+yuChm6O8OHV3XI6
m1jeTdS2RBWty6fnlCTYcLnnzmVOmZWxvMI4pHeb/Dn+Hb+vETjtKwgYkcypIUli
Dz8CiWMRxesYj7BNJqcvLdFkLdD2kbSR0hRqduyYynhlv95QK2TDnjS0JuY1MTyN
k4nuQpztF4GwAEb1Re/XZSiNvIHDCgsxwZdqMLCizaN/E3LrOF03PAKsTNNEA4rc
FA9UQyQEE1AetcaZ5IIvvKnQAAQkCdMrFS7l2hw3FF64GYlWjiw0TRtzrUwcksBF
zEENo2jwe7vwAm0/dKYWGtt8BScGvDTVoJrYYMnfA9m/eYYtIr+NkDUBxR4Wx5To
mFknkskLXC0yUIesVzdhq7kYmwyW5woQbjIUbk81nQ+BP7O2Tf+uONCr9FGCtCyb
1cGHzuxN+OXfSDaGcSffCEcSO+SAZPF7ptQHVO8W4MtSMu1LIx21exApS3mM1mSz
fs1sGXbWSljwMMjaDrC9WY75s3LZ4Nxsscdat6NPtIpLfA0zVfWL5IivAgHb828k
ofyuEK/0n2kFTXfz6H75eHiIApjjvwXdhtuHAZPoV5vKaDCOUuzi7Tt/1OgklGXL
RtpdbH4R0GSs4xAeL8Xy8fVxdO8JvVrnRuJVwVYKRMzhJJmweLIjfuvbZjqN7EPG
fpUiXKOwCdVAKI5j8ybkaHJ5JYvS3D984BTptUWNT3sitpTMbDxjeZC6k8kLVgbV
57xTV3ONxBKQw/+osAnY2jVZu9s6tZOCSbKbfhtzEReA7M1c0FITK0N9oQluQhY6
j+DwNt/wjXOABvGicpc/sQwQ6B8Jv4pzwZCO4VynWPbpWaNjeHhCiNOJ9X1lbxB+
xBEbOHxz7C9moxQmZm1oklqoACEmhlQMaCOYfgWnyNohR2LTuJWr5B8M4nyEYlmY
kJXzqibJcu1t9ra5a5zmcY+b0z4re7bli3zJ1stkih0hqNznPg8uXmALOqSjd+He
NbHpYhxwPJ0tp/UaABCsslZXuEREs5ZEazlyc+dh5G+bKTYH0MXJasN+kvDdvbSp
fiVKmX/izrz31hGztxIeJ8jnNYYevHC1J5WqvNgv5nBPuZBZrXYkfYi/WN3DeexO
R4AknBAUr/Rx6sAfrfSIiUfqVXMQXomKlnb0xB86zeE46i1JpsyzVuHkgFpMYk2o
gj78qIAxcAv+/LzXVMXWUsnuwuKhMbgELdVp7GCLxRXdxJsA5pa/IH0Euk41/t4A
xmtCHmwpSpJXV9UGGX54vmPX66hPHOQXc74rUeP2AbtA/4mhRdKlp42pN7Y3uD7r
mEOYF1OhmEuEeSy3MPogRe17PsG2PEo2qcj9qA5khFd3AKuwQ0XDcevZmD3QeR+W
qxoVi3kXVPpqxDunSmmqfzIViQ4enZN1EuCdaKP74ylGYEcgO5e2VzGXQgEH8MYr
zPXphmKscBeigy8d9MYC2fxkudBxxvoKjY7BG8d4b7wZHN2Y+25w+uetbpwif9wQ
foQEEB/TnWkx5CLZQxPtm2qZzkdi8H0LwxxAsQ/OxZwmbRwBcJb7hljADNAPZ5w9
QNsJhqi3/66Rajhitq4AJmqcJa3468eO61LWBO0525APK1/8aJ5Q7R7MrSbQuI+C
BqJpQevOSnUdik7AmtWxxIvIgx2yfusWrGTNtzO/oPL4riESBjpYScV7FYjdL/6N
UJlrT5ioZKQqCwkZ5gv3wlP1eIRENkJSaS3WIyeqJRXz4cZr10QhFLqXHKhqFv0G
9oePSXciaKfGzftxP7zH2G4bGl+PQ9uWNL2nRv5RidCdVCbr9dtNoh2pWT/ydGpp
YVY4Bg57NFt1rMLmSZ1jsf8xn8nFbR9k/NOjtUfAAn9WkbCuBaTcpnKOiPmNK9gD
isnS8CdB4nLXrIMMB2wGyQqHZsdAzKZLdvV8wJi9tqSxfmB0DZoO1BfksgMJzvAl
J2M7zaRob3vTwRfqAebsy5GMa4zbRsyseUUc+1SQBZhnlqGnmIF5qz2Nj3mV8A4M
SQGMK540uVLmjAOal58/RNnZ+0lno/9pcQiBfvnqiZx80/OTAFzjGxTXGrEwiW3+
gwUkOnwF4yXpAbr5nZd/eBhw1GYvEHoovtdu+XVeWJgmETj5OjFbQ17Zd0AAJkPH
pYMfx4az0cz8gLs4C9NBtSXnJBiAknlPLWJOveMW85s3jg5scCU31TXhPjnxjpSZ
n9RV1pNXxmussaLqtwJD4ycliOhoqSuHQ7zzcnmbEikMsARDwCYjDInPERyAlKT7
hCEHv0SPUprs8FIg98fEwwL2xY6XsA7I0btx3aYXyFHkgKZYXADPC5Nn27171czs
9jI9M7m6tVaLnEEnCLN79zy7FRlAaJjc1TOzK27ubP2I6vZZ3FM6ZMp+/ihNtwD1
tUeaQjfaZyRNoThqKg4MkO7ioiFZhIRMkDEYfq4llc6LmIfVdwVi0IdSrdQ7ikpl
YoDE8k9XINIpNYiHE/pgG7PlAkm28+kibYnMx7hmhKTH3jSjaM8SNpSB7zqADysf
tFifjSKFodvKSikc3AiGgW8V52kpTd4KtdWkEnQvs8aYJPkml2BEW7hB87VGL9vT
zImLEuXFrX3Zokdn/APiaE3gpW83WRNDvyCTbvXw9bFFGLnwaXwhYI+fShnB1+pM
N+425pHE5unVshWJLryPqu3DxYKNGUSEQyG4zIwemMcOOZtSe8IxactsmmoOhwa0
8es24LW5UBcoxU8qKng2wu50V7AO6opNtLg1dYycMrLuJIKvWhMXlsm0yxdNgZp/
tTYEfmPxw/Y9f88NSCn7Q9t/zY1HaY33bTgnw5SpecNWM5IM1PJZMo134A1jc1ci
dZRxeZ893USAf/vToNMyLsuo2dWBSzEqzjWjwsQdgyF+IbnA0drGKMpL0Z6c/KD/
mq/rFWYtNEMFFHTL8DydHcy/yiI38LlqEXPj9/oB9BokS2iG+jJJpntbmWMUoUSS
656okgjZb+yzIfdWy8uRzAwoqpYBvREMDmV+hZsVKKF44ue5wf6J4Di8LYqODc3H
b2gVyGIECMhkoXM/tli+bvQJZWSRG4foT9/e1A8eLQbfwy46MOKtMKwPx6qIJ1B/
Pmjie+kP6CU8EeoloJHspLRyVzJ4dJtqRAtmwAqW60+VdQV10eHWruis3lr5L23e
Pb0TWywJyKiqe35uq8XNhYNhDY2mafTOJna2ULs4xU+Vav2LvRBYyDfa/RLCk8uw
rGVJi6clBujRMp6UTGM9OrtApu+ZAAsKOJW3K66cj4yF3xeFa2I9aaxfPVcbPjZX
ylI8Dt/RaI/8AqkV6g6DkeFgEqEzqJ7ejVWjvv6ZiTPvHCjBy1IDn4AYgnSEPBg8
F7RYHf8o0tD9cXQV2HpHAVXtqrZRvwgTuRecnITBTVBl8uSfDayocrs8tUfr3N5E
Vf0Y5Bccj991E0dotcbgU34qFiw8rzF00mEwJW3E4FnzALdRJp5ISZ4NIkL5tEq7
jI4qjUdwYM8fPMrA9SVIAc+YG3P5GPIsdf18Ueb+ZJhnFx3UM3eKjS+aV/WyK//0
Nz2VOU5WX/CbOf9iFS6yRTs5J4bOzZ8IIJrHquoPHitPnay6a7Ab4+5SKdWwK2eK
GkNwdN+5KSLyLIQbPVcVjYyrN1nrakeun6DsXwb1I6bEASoPhl4MK3JObST/ImIM
wAmQ3Z0+es6XgS90b0t9oiKXrdgc6a8WUBNTxiu4OhFkSTuqlmbLWpNeeg7LLFIY
LGN1qA7aaMqDQTvKSplLK0bMUTdG4XX7GQ446Zln5JORCP9R4xqtAxfCIRnLjYLP
bVg2G35LewkbON+3oZmWYTXcd6/fFS5mt5IYtkivkm90kmCV00Q73S2focNDp29C
ZmUaIt/bJxzCZ1GUJxRz10D2TZ8oX+fIQaqwpz/SgF36Ew+8DnToZj8RygdqTARh
DzQoo3kxtscnviRSn6uxESUbmivJfV4NWnhKmqrhEiWgDvoSRq6vrdL0YY5nRwoV
mA3LklH4CtQ1G01GdSbyhB80PABxjR+IN8ur/Cf+0MBhG31Wrxiq96FXwbz5wQrE
Qhdw+ThJfszQ4Xr4JdnPW0xHKFzw4cX6xZ8HNuY8qty5Hma/gl0iKwzf8DGhGtIZ
kEdS8U3KRPMMh4Ynaagp3C6fESHF2iezoFuC1/UZZQiqtC44U2aGzUy9Zzu5aUSo
EfaMo36NauDP4Vk8xT6yUnkgDwnV50ne/ouo686yo00g4Wz3yDcuEM5EXjvgCxqj
hAcl0nQOXkHAhE6rnmIUBHbCofSzx/51RIy85rzKWhHDQF1IuujipiHA/cCoU0sq
zxNNhTdlgaNd5dvWaSwDkfOOfKIp+PFbGrfmi1WeD2IO9enAGPvOSzI7Iz4hV+6j
MYtOKSBIkRpjoTeAxSVbLTBoYZ9VnIfx8Q5EDy6OgTcKsePN/2TRVbF5DYzt1Eh/
hL5i1SffYBQOw0N1AU1beR7xVb/eRWBJh4dfc2rVoYsvjIjwF8M1vuZo+UrWl0xN
BeiPrY2RABbh2mhNJbhyEqIqgt+6dAZ9yYms43SWf+QOXHMxubYwALvE/dfLjUMa
Rvigq9kYSg3AmC+nzPOBeZlE79pG8nDbQmIhA5HP+Lm7zUeqRgXQ9aFXsP4SRZRc
p7wFbce48uv3c8eXSfiDUmQsaGf/eFZjNfgU3JOKZETKJZ90/E0G9p2NSAopDjcl
w+bceIYl4gVPcQrJe9rJdFw9tONNDiqG+EDWP5FH10IDE4xqxWRSLrx8eNDdyipU
rXknSyXKuggt26DRgMsRaHubvAf/A88NF9PVYL/HNqlSSCt7nTm4rw9/AxgYjpY7
Gy/LWKy2A/BShdgD3EnYrLHesryIjffqFjEGKKNdDGNeksgzP3GC3uK+bkFDn4Ax
x5oi6R5JBO7VhpPjwkUKITlu1C9K17wWnSf3Ixhuv/o3Nkk6ItYjo2kCG8Q/kHhp
bjwTR3jQcrhlJbROTtRVWOQM29YrJQlxrQTuF65o3vhiOhE78jnTBBZ63RNjVs4J
jcncoZ+uXpkWfj5E6UG7Dv6uvStTzQQ4dVsf1fM7z6aXlRMf1zCR9pcrCVM+0Yoi
ZiRTv+3DTohmy6TiSCgxppv/0R563r7mM+IVIbewE98EfTJ3O50bmByQ1ALIOzz0
VBDMbCpN3duipMeX+CSAD7XwU1/ZYhbzouX/d7R56XyOoXsygKZGznLvs40y7soI
vHmuAsXREaMmPNQvGgaCEMMdXhdm0iFbm9vksSAgcRR+TejjEnfSHUfeToAPzsij
rQi6jx0tC3Xye0q3oJL30dO2EvYCZJ85h7nxdXh/uWKPNSja2zNvHwZmVqyCJ0QL
Js4OU/X/40eOrSemjpcC8rnSpzJRt7K9e5/RupnTUtcD4/LczbAkBh1jMLHkuaL+
diXciuxwl7iVWsYlyChcyrNycm9VRVd0lumLW2EKaB0wf2B2UH2Ug8/N07GDp92B
85SHLtE7Tk93BtqrxX+cH5R0+ql1bvWNUP5jbSN2vGZpAAo+O6F+o6AOzmOXxGQ6
uekxriHllAv1vUFhhftDHvbyRF7fneLaQ3t1qygu6qmHyAbNNokBhcGzlRZK+tfF
l2joQkqBS59CB253d+6dpYSEWhUMyftSdMg4dgPBiSk6E/IK3OlicFTXqqaqUZx/
0GbMlFV1dfeT0Q7HWcg68SMEXWEstlBtLmj4z+7weDlOSC739cI3BVYku2nucFnd
hq6nD9BC2DCx7B3/vd6K74q321cF1iPHJB99/NpQ6a7FhG2IsL/ZjqAJqB7K1P9R
x3vbnRZjn7/zLty+Mkcuead3hs7pE08wGUl8143eaNxkJyAG66uKbS2tcsiESMiK
BgOHWeoWPakuIwDNbQivmqsI+JU8485bi8S5ycMgcDA0g3qRJPw7wse6JO2eSRyg
R+RcHhVCmFAF5HNauYXxqyXC4uGqz7opyyra0Itk7kN0Vn9FC00ZzM/3HujPiO8A
dMto7KUH+vrpPyWTIw6kpPu0lOyovCJ23JEyDkYm7lMS8m8GQef/PvLJXF4nVFMx
+cOVW6XCCvNYr3aKoY0uPSFR2t19bfbalyybr42Bgm/dH9YZTEIYgEw8A6qSteF8
hY+7b+8VhtWoJ8nBLMZtLFhR+P7nviC3Ut8g7dCtspKEGRndRPwy1kcj2ox2roKN
hnV8lIZJ/IBdiWkz+/4+5024dAwnKYcGlZYBIFBHCNQGCaQLaAtyS4X2gZWYqKSf
gX4/6ZSuetPdz2zc2mSSZSjMVjb28xUzqPl1/CQyaA0uK5YxroGh+AXtLdzbI+a8
f00VcZq2oFUSQ4V6KI3uGj2+v3eleBOWxn+CUuuwDhgVhTANkNpO3WVCegCijlN/
C4SeqkOVIj45XxY8DQdlNU4NSqAfRmGp/EUUz7mXSXX4FwwpTiAtF2dWpFIEww/l
MSZknBIu699H64AvUggIozZk6TBT4J/TETJGx6/eV7FjL5PBmNnrczJkLcB/Ib1B
X7mgPyRZ5D7Z1yey4ijYii13vcoOz2eOfOMfQEMSacWq56IBgooK0rROYtylyywn
Tb+Fw5A1/c4xSLcb6wR09q9Zm2flHvLubnZwNpLOJivrEeiyWXF3qB24Sk0gl06B
XL7FN5xI0bDNBMP+NbV3r1iGo88ii/Af6tAeAWwlE0iSJiXi8vchqmEvuZXtly/X
bO1X9FsyaifbIpRwFq75vke27FcIPKMQxav6fb2fQO0GYurdcQisY8bQSm7pmar+
keBUMEQ4eZUZ1yW4QlIeiHu68kpBT+iq9Ogxtgy4WkF+0zPiNllLZ9yMKp3n+3BK
4VBEZ4Rjqrv3OHX8E5l8OxHYZDxbebkEh/s8v1AQedySi0XJVSINI/Yy/y+eoW5G
nxL4fblkAq36EfCoRttKsTr3pVIRahhs01x7MKCMQK6ewVCLn0zcgi4a1u6b1a/e
lk4mInIr3tgHtkgdd7USEj6aC1nnW4wuyMflBS2/BV5rhNgwZKtDAxp6EFNje6WT
ukHJopyyIL8GFThOvFy1JVF9dP2ueRRVehZCmb0vjKixQxMtt5SUOGntA1vaIL7I
UhQFaZBV/GPOgl676iXP40AGJHywHs9Fl/giKobXBKPVJ69SBp855uviJxOiNkOp
yY+zhpncviyrlBGW3dHNINlJtdm11QsOQfqeXjHjZCnQA67HVPKG9wwm1+U38yCT
BgglvuXY1x5P2jG1feG9FBxw/ByRF3GfhAi5oLnrBRgSIcqrL23uWF1UDJ0jNoSS
vxhxYRclfYvEIKPS/JB57iJafsca/UNiDb60F4YP2j5UfVF3J/nZqPnl43gS/Lza
bWtLR6ng5KDCsWTUTi7uj1Ixs1o3NueKXyKflCA1xcH/zpq8nxu6bEcjWHPR2kmm
fe+JqjYSL2aQH+EwTILmM32h+Czv8tUHNSuhYVW/3qDA0qyiLZ82VKYwD2RFOR5w
D0l3P49hT92kbtCspMR0Hcr8XQ9Oy+K67keQFxAizu5/JPm7R9WcQqxUub0+gARu
2Ll1IFLJw7ztXsvvsa5D5jlAQH44KdHsVtsByZvWFJz7KutXc4MnhYxCAvce8i90
z/5/aHLWK+OYWI2U2b9PW2/z2FogfFVXdK4SuTHpPL/1J4EEyrO8qVbD0xz5Qbcq
/7CFePCKRySKKFfQmxy6wLb1mNvur+uV0kK70arPaoP8SlpyD184s7phPwMSts0o
zVipH1gSxOZ0UMnGLpbLdWF+xkGwlgC0ctB0Vlr0wS32wG0WqK9mkkiEjgWb7TjG
LQyA+vwrDXQKK//3NgxM/i4lNR3HXJx4A2vQXHSvBfAOO3WDhJatzMMSPsmmU4p+
Mg5gyxVPFMV9TEHBIBMORzDczTtaQX8WNl83f4pO6E5nFZ/qc8DxaMg1upHB+lCd
OrrHOgckqE4ZayCngtSSJcejSNuPve63ZW0ClUnstnu+YWG+GCuMXptLdPJDSDen
TR0bvQfEehC3S4APn70IQXhvrxZ6aZp0nF6aizt939TfwHbVtQxqzBaZ3vZvtLKi
azmCeLKADeTHRyuZkLNlGQOgFEOtAG7ml5FSjHMyHlr8spOLpvxarjp0CvXkERJY
QKdmOU1lVdQasYGD2QcUZ4PoFGpL4yqCCaAwIKikQuqj93CRXbMgdWFNfyzHBMal
QsaAJynzc4jGiKFcWgRKBlGaRzfDKF/XdVisgHg+pcTu6FscZ00nTIdFJx3m+IFw
tXvcMt1S6oA85jvGYWYcYD4dEyS2qPIPagipxiwfYh8Ij8lJy/M+gZGLlBWulLxt
FeRZzWO+utiBjlp8zeN5lU7G7jllPGlXmF5AEL4Sq6c+U4ynxrnhYPA99PKO7SiA
k/8FU/iqYDqUrHJN26Qin8d64UgXMmwPnpMbCERcoesp9U6jxMUNWRhamBbL3Roj
f8kq22Na3OC26Sqo32ZJZmqCkzA8yn5xfgi6UYzK1Yoh2xUslpT0GsKnWXh6+6OG
6/rjDM1tLNPF1zMkMm2TdMj5I3rI2mWl27FmH4SsX0hVxUgDVCWZwRKTYj3mJmbP
5ritLlLty3V5jisEU+69Z3cvopnLOv1k1RUyPlQeSD8pltGPgPIISSm5xivsQWXq
6b8/85TdpGwsUId3xB9TP8+Cr1GKzahfO9EXYL+ZOrb8arR5hU3r9KIXZpXFNkZ3
YDZfo7fvHLTYI9AaGWfTMp5IenVJ5vswPht16iTGwfChJ+bmOVY+zHo9oio1/m8p
r5WDhPFnpoECl4WWQ9dRuQf6abePHNqgYxK2kDkNBzJ/ehYSd+0goVu0WMFx/b7n
qnITeWQjgNOXnqG9zXaenj+E52eSu/Ndcqp4lfQRsjObXvRRwmqGt8qsaGTrT0A0
YZcJR/gmdPkFOGYa3GwdQefZgwv+K1nNZEK5WvqH7Ena+NKADeQRRGZMaN4nR8cZ
Mj0woO7FbDio53DUT0HzFuWU34XjZTFqb4UdCxTeqF5Z4dRmGn9wGc0l/XfG/t6k
wikHLdOCdYdnZzqQZFl6sbxwc9eUp6aHDWp+U0Y+I8UpmD/Xd4SaTgr8zp2k2W3P
bZAnussEnEdknKkwxNU5eUYDznKQu1oBYfSBYSr/7w/gPfLKIX77nwHUYeolB1mw
HCE/UWG+ahJr8dgPefsY+SgOPetRUBoR6D3HuWTri73vzdcB56Sery3nWweH69wt
M7POFLZFse4ze2msd4wcSPMCrCdrdF9f60ron4qSxiWrzoXPQE0CFgy07mClVtuT
WsULuMr4xXsQiS1QUED3kfMUSdF9DQHGBYDpy9T3Yk7tXk99hLXchnyHoYJLOyni
mnzyKxrCqhawIgBDyJczma7p9PMxbDK4Pa+glV4EX708usgd7wxm5QJwqEkO3/An
vsSyIDUvduPyTjAVq2Sn5BBiHLOwRBu5eTaIjmvnCLuwhLKoJn8B1yzFghTJbo6G
RFp+EW7vkg6skDtwCLUzotQEo2VGl4ZlOGMnQ7OwUyGU5xgOqXpmhQGS2N/lEEAs
QxKmxlIlQ/wsJQ3aZ98BKZ9+glt4bWC7pLbsHCyHqxo5xD/7eE0gCBPfp89dfie6
pqvQLgS5KdaIneLLDgGSnJSQHrzQC+nLFyNxdcLdGlEuxhj8tpGSfzEl8CTHqKVK
vMRkww4FmyNOtXnrhaMMX71ztFKPxaCgmqjwtodV+o/yYemXVowPSh4SyHaSo3/M
5RSBd/GM1SuzTpUbN/HSeHc9QeK2KE3kbWeK+I5r5bQpJtD3ZQaGdj0spnAqnwuI
ZbtQuQ9DxCZmwJGLLS+rd0dqTSAujIENsf52nXgOpeoeI43ref13YJSwAzzF9ZyE
tsNYJK0EWnbtOnhzAWrbnGxiHad24RQFTYexikBkaS6nqBT9ZMtxkKfkfWL1pZ6m
v774ckfZqJntOHEWeNVxnT+BAzWwFn1w9TkzBx6ONvuA2tshrIvwXz/6DK7NoUuf
f7n4JUNpK8C4TKUpn2sjnxEPJHr7EZtM8gNeNYOzwXw/rVYh87oDg8Rk6oCjL4Ji
UsnzbPfM66KJaFKCzGwZ17za1ssqWYKG/j0ordxEW2Um46S7Kn0iMLlAT+0BgtKp
Lcc/U2J3Nv9Wgw53tOWY99v/1luMJmA9BrXmBVIXqkKb13Tox2VZztAQpTKqTk/u
b766Xo7DvJoQ4tNOJF9D/MtFF2hYhyj5P4gm3rYhYUsFtpmoaQ/gDgoXKf6cefN4
xi5roXq9VKWBV5IsqbcbchSPjVCWRoHjMKDE9888A4/z38Q48kdtlvQjaQ5c7O2p
6yGwNqxfprsgg10LJNCbU2QJ4XizWPUySd8PG2Sdt5AvH4U6rqnsaNxSkZUxlEAg
4AyjjFmAQR/Lmzd7wQ3c61F8nE8S2THduVsRwvbdmJy3dfe38hFrx+gWXreeqc22
+iWh1i5qBH1pl6tjnsjtR1wiB/bKqkvwvo083Ki1QRunOXLshW6IwPvM/tg7I2qU
hmr+/3CwUimCmVtiC3Qt3p+O0FLdkXHR03nk9XzfvztW8lNV1qgXIR89BY2snFAH
hhCUVH2QoMM3r766fVjUn8e/iFoEnyikh8tY8DIa7Qu4Rwgi9LIO1oANSwPYuRjp
inGht4somIztJgc5DpGuncvUeAhc0yo89Nb94lN9r61cc5KRJiI/6o6RuWAoZtlF
bsuDgUyInKc/StDbPMZ0VZ9mjcuSJnzBS6cPjAmYrAzTdJPI2sKnioweXS5dbwMh
3UjHenuHTKvfNQXJc3ef292RKg/b0FqetXhuE30/uYFzcflpEgu8eUk/9PJgPdgQ
/nNuwT7gb6srdvLc13GNI7yIV+XjzE4FmiOkbJosYJI/22LxAesWH8lSUIZZjozn
LwTaQHWw8ceH/HcqBBg6ugemUHI9ECA3bhNLyWdx5r0bHf7OZSTA5S05gHkomwdv
ciXBjy8Bips2MK1nntx+rKk8/yBod28vHRoY39pQpbysX3vahJgDnS9QZZW/AGUz
i9FhGpDLsOTZA5kxGrZyVztOZSNH5Mm4827nutXtJmnrIMGOoPcaSIPx+dqUT4SM
584CSeuPdjMBtLU3VuwpffhKlVmZiIESPNmlXQRsOEeDJpsgiIFPVZJWzgE/s7Kv
XnxB2EDN9gkSIrm0GfwgUZLNrDXzy/BCE9teYMjLgieGyT6iS54PXistA3czvoFS
/9HMeaiEZP/8V+tTXco2kZNOLJ3Oc5gSDT54DbEql2BUjUUQUMIru5smJA754isD
Iwl3MsXfdnvTDo5DT9Ri8RcQEuBWgUaaC20eccGNTLJr07qsUdEqu9L3aMyCgjza
YAQkgD9K2mDEBVza9nNE6gLbfN20IYZHVd3+d168cx8ghq6NB0ZamL5JurncOpc8
UMXW+8j97yC8ibpIMSB8HNdsZzfCMeb7CunB3i4N2o1Xo13CoKNwduCqTOZtvS+O
Zs6Lqa8gyNn/2zossIhm1+Mxkix0oRqMXhxirLQJ1OBSeu3VO3pQ4HSPRofLW8Xm
7xg9V4eOZ/Wpz9U+7HSqcbA5IfI/eV+ekaMuMv4RMVdMvCgfBm36St15EY3kkjD8
cB9EefqGM+kYwzP6G5ackzU1Qr8Q960cXN8ojV5FbkjM/UkSlNpB+ronIbJENQXk
X5naHMTxqiGeyHKTlSJDmN0NcmHA7w/KeVB4wgmPmQJKECjIsojMOGVKRayyH+ry
rl/rhybW9Gt5YpkHM8kKeHHrHCSJemuabUXbs4ulFaTIca1ohQXO3Gd2HVz5uwQS
d3FE2dPqbj/cIN+bO/hy6gTbtmE38Uixvqz4d8BfHgvcgGzATobNKMnV19UI/FeN
37z/GbQbz4QlolIPfdFU+bNYa7PcHYS5oDjfpHwmy2YtoLFLJWUKClnVV3N0eZqC
4x0v2u+1k1ROM0Q+Vzb/QkbakKw14tM4r84ya2dRNuDdPXy2SQTH4huoXaLD0SpR
2+H9cTmsPpjTS3FPg0An8OR4k4kKPl6K6N52WIa1h8jxrsQ1MhyvDZmtk3/vfR9S
T6ga18kpYy18ATq6Gsiv06q+ZAlr6g7U/NQj5WCe1hyZf83SfbrC50ZopFtoL6qX
hz5rjgNNG7jZdkyqZA210qWCc2HF6qG2CXqjltuprmciWf6y2f4P36gVngk6t1MY
swLZr2vgkKimLQuyIygpa3Hp2N8QrIlMDprCla/Hn8qasO0b1+9wbDWJnFkyygM+
TyiKu/ZP7j0pddNHjEJIIdxruOC9lKwB2YGRd/zNgMui99hpbN81nX3e1sfH6aHN
GmBcx32+nOXDVEGU5ezOUYU2sAGe+f45o+OfjUQrtWXQXpuKRXgAyytYiOKqIrYA
MGyf51pS5jIV6tzdoLstixvLVYVDWjoi9ndX6pHWaLiqJj/Dwvs3muyJpkwNx3ix
YOHDbq9IqMUQLumN3eU7VVt8zweGlSZani9hcjXkjTFjEsCxiLtbjj2b2GJE0NRv
4Uh0SOckv2CjdKr5n1nNs5K5x7ql67wDUolcmW/UYYDWw/3nJ3P9Olbm7un1AH+v
wB1Rl2ZidoXWt3+FeiFRLq7sv5UpGGkuqljtzm/KRtgkezJBq1MQt4cswRiWq8KU
OViuifx4st2ZgiS0h/Wyx91XQnrysOX03jtCrnUXuRskGGyqkmZKfxBwtFP3+Nlm
tC9NqVtORjTkN1Md5kZ12FurViY1QJfFtPqvwRj5v/mGzMtaaj05/W3N2HuFOBP4
d3OXZXxNuBGptqCsx19Qcm1MwVZQj2qLNHS9oKO+M+lTIBveb81S11O51mVmWg4V
DtYcBPT/siJRrSDzipzoPBIATf+FC+D0FkpG5jML8cBm3n2K0NohL3yYBmRoSMqo
it2ILrCzRtqUffN2WslW8DVct+D3yfhjnse6Olag42L1TjsjdLawrtPEETSqwtUN
UYT/o3jT8OUQA9AwWltPFecpZn+FsvUn0AZoe86oeMpxLSdgFL6b5YpgyT6Gf9Sn
jC+2mtE0vG5QxVCXGl7epSPFDm0WEWcJr5lI3dwWA/KPGz0B3BjvkBhY2/ktvaHG
gxmPWNDpWRrcId/LEGRj86Pu77N1YUiABCLA90Zm5xwuLPjv7JOxjeL411/iX6+b
WxkHybX6MncCo/OSYpqIkCWVE3iBRdlacbQ+Q1Tx+qyOLHIZ5+zRCB0Osik37xHK
r4HmoM8FF0SJ+KGg6ZXJL4QCinMSIEk5cymeRkF26MhmogVKn6rV6gsyNRtD27Vt
nKeyTMHR3657oXch5TVUHtKJ0QjoJkdZv0lscW1NKGas+hBIjgbbGCXZmXgyo9WT
qjwsIoerYf0eKJtcamCXgjki1rP09Q/hkI1zSbTacxB7vYs1n0QJfZdDx1dfLkOf
TlMIaWt8xgDLUYg0DDelfrHu3lGUUHG+6hI9ADtTaXQAdes+zmugoNRIQOTZs3dd
Yco+vIh1OjW/595/bVZ+wKwaf6ldUW9gnfJLH5QjO2L+0xabrWTRHySxSUODyJIg
nGAlmzgW6bCXUsKPNmgA5khPlQolZQs7mwEUAo6zGOHuNFmMVgOnS5lfGqvcFFyG
BWmQ4y17RmQScpzSbYB04cfOuB2IpDhLti1B4TQoXTJEOoK3mYgDSEnnsnDNAPFF
TCt1CFqhDCr97E7oo4RtnpM9DRpHCWVAPcGsbfk2iyu3N1iQf1J5M/ZODvHE6jBO
X3Qtb7piERH/hrYOGHyPM+bL2xadUHTLsCLVfAedjP48pQkLizeSlSLFm61oISrY
G35dxjuWLRLElONbNBkJWx0HXYAH4n/3lHHWJPMahzVzfk7cw/kWv/YoGiHE1qz/
bh6qUWLD0v+FGzVJT0Rm2tnyfPRwXV87TbbL6pMTslhff+7OANCVOisM8+IyLjgG
WMxxfc9R9NOnLvX9cPV7pXYFMPFBVuAbdCANWwZNFHKwrVxL+8EULzCTg0kggdLg
R+Idegws2kvufBYOFgt6qtO5WmZFwL2UhiP0gWHIzKJhjhEh7quh2LekeUs1jYJt
YjbmXdMYPw2Ff42cQtYDFoXGIN9IOJwBXcbR8D1LB2gsTVdb6BCa8yjMyQMQFXCU
JJU82KWNLxoYdSgc5/9IYthdhvzpd+DDDKKB3UukyJ80Q5RtHoMDmI8yIvMlLpxK
0C0XHi0xQsXNQXBu0sMMA2ielSocdza3lw54iJ90AO6vlnxhyCDXgOn/kY1p5xnI
007msOObE+pMUuzWsQZFjE3m3cUbSOIje8bkw6ODy9RDg11iTQCggx3PQMJvI7i4
DuNqLqr/H6lWenTh78apqmVfW1hpUIwKP7FPx1Xt/KQu/X/EP+2RXSu/MDJkAYvx
cs5dL0J2Q6kxUjhnr6ZMjT/f/p98y8UU+hZzX3mH8uP6sYOVz2FxPpqchBOCgzgS
D5ENeR4O0dCUHai8LP0se7Rk+0gNmLo3vkL96t4qvjkYMw4SWwAEjL06gpbXw1Dp
u8SqBo2YPdF9vBmNPJMAb3UhyTYwRDPdpKOm+rth3Ts36akchYpnh3iSbUxGRhxf
T3MgTGxz0PSWXubNCvNF8egbRet589AKZmh7zlyBhCEdeFWJwhE7U8Xa9VA7FwS5
xey6dZB7J1wEVhmyIMDhzGopOn6eCXtUP+H18WCMW2yPSp2UBtVDwRRl1uUQXDiR
tr18bY/gMtJZT1EAhetZle+V1DxeLjfWOQoHCLqeOB86EJLgZt3Lkxuf8AXMUXng
qYvhYZ/8tNighCJDbfSmWnWcwDODRp6l7BpBqHFGvmcjkdRdFrBd1STYvzzcuobc
HUVhXfGF8z/LcKfGwdyeubKVfHfNPdPVWVNYrkLgoGP+KZN6wkc5jEOdUpENpKlA
I5teWYtGhpNj90aGJhf02PRMH2dEXaexSZPA6uroHHt8O6bA4fwfGAH9j3v628Ax
rjYp6RE5JjJakRBjIc29Q5mTvSYh3a3/ATcCITBTWn13LcMgAN94rrF2VzT/pGz8
sZGDwmAKMgRM74BgLJ1VX6IL3KAgoV+YBGA70xY+5skzp6I4VahRL8Pi5K7aMpH/
fiW0nuOO8ITIzjnv/lb/xvkiPxMRJNqY2DiuRQyIydWnzX+d1fgcfRl2piEXm4yl
3cmz1SDvz75bxepSM08xwADKDkVjXsdwJFSMw3apHN+7rtA8wGFKXJcPfzzwDUP8
UKMWEmoFVbpPLl13tjC1FuFPOc2oB1Gv0fcdTwC2w5BNs4ntC+iPZU78kljZAJLb
sCPUl9o6JTWiGd9N9wBqyExH+yS1oR5F/VvDeR14PcNWCnqYIO6D6tDK8I+TxUfJ
6lNMxJhYJ5GJQkAeuLncl/PXxjIKQfa8TAVeTNBda+SbR6KQphFayB9aCMZmVbA0
qUR0PBdm/L8rYnnFAUSR+EN99DrmdtvhkqsIGl8pJNgwV48Dtl11uvW+7WspeyvE
bMI4vZZJ+WCjqUSqUy21ud+FmPbuO+Bw174hA4MOYD8UTP4wYRXKQhWye7nnXthS
0D7KiFVTTzMnXBjCsta3/rZHmtdUZUXd65rdxD09azGINwGOVVVXcU0VnDB6d6wZ
plePdYBNU1VZtNL3TfNF70hizuJJxW3mox9+wCTJIIQnzs3sgx4Kxx1/rj6Oi5UK
HrUbu0XdRrkqxv3gYDbxMytuqo7kZYjuykBqdqMfVf/uilav8ffRr5u0TsUTfY+J
JrQV8uu3cDROZfnZvLYDib+/3kn3ZB0RiEep3QkcOfZCa1mObwNAwlzSmVon5HAy
oYSyIbX6vj677hHEND+0TPb6GHE2xMolBQK8opCciUvX1gFYNyhK4RdC9ok4TJ8B
cqYithMNLGgWwWSocmrzHqb/j+bGL4T5hlQN4beLTmuyrAEFr4FOAnuVs2MgbjjL
NZLX5vFyx+IWkrWRDEtObAlMXOURcPgNHWDuxWodrdBVG8AE5Ln+qZT5LPH/CSn/
47FVS4mL+wYIdKjdGZ4fZomB2a1ONVh/IPQuOV4mnaqrYbe0WsIBKs0UeUagHcxs
dR//nqQkF/d4sxHYUXaJQ7Ea9ZOryFlZlIl2OHjLzodczZeDdyspX0FzArBr01XW
3y3qwEYRHRVQWCpEnJ39M5ocEx2RGhRFRbswypwbRiteD650wfqBTkiot/dy5AvX
WOrILNarGDJSq6t1kx/th++wE4WIUUF262S/bqFk3jRstbSq1QZHRaGeRcjbjRnI
OpqGGSff/qY7SAgCG2IAIX6/MZAiG46/kgeZY5U13BpYolDI5HvF60FGxduY3CqG
PcePfjdO1pr5Vplx86D+DJABCbQlqVvQ91AyJ2eEzzLq50y+JEuY890Xx7T6dZPB
JN8tDzOt3yx6HRnn9JoqSUFqjtCP4LaQBVNIH3f7nif80GMdhviFfUm19jLAQ7d1
waxFgYijCXXrt/z0SonS2qhDwLFfHJsZ5JuRwTOhl7jToG0+clbUVhW6shYbC8aW
9EwrQu+eExE7MTffOyOnMlXQNuecmw7DaCIv1ASyOF/ORRMNuGoTugzWXEUYlipP
14oM+/Bq/NyBvHmaM5BEJkoKmaM9+pGgxM3p6Xz/H1h6o6gKknrsn8I/MQBwMdWx
tlrFmTS0QdRKQa8vCsR4ZzgdJ1Io78mY0kks9Moqe4FCmhew3ZuVupb1iNTWMK4O
/yqcRQNqYJ0kjGM2ZtzOKHHFyQGeJ5VhuzDNEVhcHv7X/AVeRj7g+b7c8RXrUD1n
2/T2OTvZEs7Ig0qIxndD+AX3zgcKlAw1IMv4B3DGjdeYcsrntMRXRu/qyXq354yt
FwxwCn9ZtpXZKRqvuMB1eh19Pzh8HnQ3BwzS8pmAJFoU/2QMPrEroGzWTkATql/t
WVAoH4P49DXiZ7f+chdGktVflRtcAPPjwXa4HqjXy6LVhv0fxVZGy66CslgEa9Ff
a4K0fucO5L/LlSGCsaLaN9HsGfcY6Uvdw+9mOwk5/M9IIoTJXo6x551aQWfpS367
aOHFAk3blndnrNSPXkfUpQpIf9O9dKbLsVu1Wm+3fGLVrLSM0P+TOwKGeaWdI38a
rCDiSQe5UAw3AxqQxQf7pt2990SaWEju2I1G3cGP+mwLvlFWrJkAMy1a52EkUv35
6dMRXXgtPSCMwK6r2d/bDejea1JKD8g6UyUMonQhb2T7FYpzTFpVUPs8zxuEhdMx
DUGZlTB/OeYmBK8z9Y7DJzPbR34ODhEBcEI9tNG69FYlRK8rOc84G5+7puTR8SLD
xsqLiBRqgfxI8yXgLgRpmdWgvxk2p4F/l322sZf6CbCCZNKf55/d1e/23wDNyfv+
bJY5abbrqlhSvbObzrBBHw5/wJesK84TRiqXN2pFOhIxFZXr3x+WRxIt05BUVXOx
yEI6/247zQkllIZk6vjIEm7bAQV54zbPYwb5nBcjasQISYm99sXwfAfs4o6mNavi
hdQl++FxenlAYWtIPkVlmt+IlM7LZu5Uh3r2xWSSlT9Gx6tv/CkELtNO8hDQKuQh
9WISmiLMhTsn9mOHQr2a1TDm35KW+AbA4jDiS1oKZHnbpbKZmZuwcfsnfUhahj1m
fMXnMofVwcKluDtsG93prHV1i93lV91jSVp9QAYwJDoOwRp2j/m/xRfd+8/YmCzO
barz1bEh9oT1LZNLBTTNDFctWJ115AUgG6jiZK20npaxAk4aJCMedPL24g/iZwAz
YtYfvyFOyPWbzraMQDdyc4gRMvCakKFQbdy2LLjpTqT36R8tzFZbgRkaB0ZgIkqD
LNaA/2QCB+3HCLBj3rsPYdu4bzbw0knP/0yr6cpMbKsAb+fsdkId8sIxJYMhM6jE
2/oYm31LplJSDugTS748cnLK4ANZF29ya7OjDJc7x27J/ew0Heab94J2vqHQDO2D
K0FcB5+vT/mb9HWAV+Xi2C1W6JjvYr9qoFvhCJE2HPqmpxygS9zL1lxvTq8P4BUZ
wCp2cdDBqVw/OLUzbLSZMcOM2kwNOgVcw67VPwB96bfAft2R46d9ba4lRYvs3rGU
gEKGh8gIJxxWtESPdJ0GbpY7Qi0YkwfB+aZHemxuedSXKJa+z0wf3NOACLLf+rJ4
u82yyRMezX64wJhY9CRUgNkjJl6iWglkJH5D+H57ln70VQlYPOYFzh1HxEI9Q1qt
5bl0fsgvv2RzoT+CbtL8LsQExC7FIS7+jXtFH2soxf1frfN2p5jmgRQLZ747AJ+c
a2p5EJSZLOiwd0aH4aEDsjPcmpHwb/qiGOi25g7hP8NrLSgemAyXLsvfgqhGP92Q
701n3IzGwsooAPmxeEGkIbDkq4OAaFxQNuE+kNGzLXsOSCuLapytjsStAmrVYK0k
vh4ic+4A/eKHEEFHzhZeUC8+DJBUBpoc+gPIQVLfv78tT8rwc/wf+D8HB4XBTIN1
yK8f9lwySrZlVLGGGUU447KfgnvDlIUFp2remQkz1TFAnQQA5GzorOTQ+4ILFPXj
Y6OCw5/DqIgTZqpb3ULVDwaWeDxTobitBNv6YbADxKQdNqS0fG13O8OnHO8sOGiU
4djsovL/EXvi8mK3bB2sm8jZUy44pAS4zWlBelUutdBHV8qBNvNh/yRL4oJXN0uE
U/++emFlwKKRAdAIV+tts0CLcbiqWPx9SG5TngHVfVAqsvrKTB/jxVMhBhlSti+y
f/34zBiF8fXPTis+uVZBYDqpgxBpirTdjIRbAAkwPXSwsPG5AF9X3GKJziCznjCK
ouX20TjE28agKhrlwAJfo5MTjUlAdZtU6nrv0XUhgiOSxUAO2ImgxVY3PzLJ2GRD
w/GzzZz4hxEI56BuOvfL6pFMaVpQBsX1JHbcRcYynMy/Q0XR97jbss9JHueri34k
SUM7zet0a1ma+BxkiUGkxkMgFTKNI3CVBm6zcPCgQ6GJgc3ypXvbgoZe1SbRuI6w
OLB5a6rNRlojBPwWyk27+E45CXaAWhMM8kFCjvO8zXzkK5ax+YQreOSEhZbkG9x3
AHB2eFGMyXzch2uME1lm584fSWcQ3ccpEjZ5YTZk7vncG23Yg8s7szxS/Er6qNHQ
FExn+EencMlMDD4wm6pP3KFtv41YJYk1tVEXnsnm3wvSpuXEVUx6ypnDdvRd8Gku
7L0mkMt42XmtdUYZxfXKHIRCuZwQUfZLzpTcNlVrg0LBxauyrPFFX75YeR0tkz5H
SStrXK3xgVHcK6qGe53z+3ENQPtoz7o+cIZS3lkcyS7FoGJHBotlirEInTyt2M2d
BJlIfnck4OfzwrD71bkh5j94ApIdt4dNrPrCmzLBcQ0gNTZjcGICBL4yKL6r5aEn
pzL7RntP4VOu9JK5/75P6uG0zik+YpDO/RexcgGrJkEKJWkkqmZQGMEPk3CbVBu3
nOpDA1pghRi9TQx1O9uv8ag0PIBa1oeOU+p4NcRl1vW0dTteXh6UGlHsB3/seh0o
bcbIJyPDUVDPhS1u83HGPCLXe2Vl7v66bgmYlbFSEVDJ/VxV7ZF/PWcJEFxVVNCF
7MOtDDzIkZZuhbAYVXVBGjFVRgL/+L71bM6KVa033caNROleNPoBAoo+XiDHqJSr
vJOfMfhy1KCQTf+3NrFAUoD701+mTqw/mT7tmcEH2rMELzEwxES1ZGCGt2dDSHCa
AsBeBhS4STSn+1BTJDK4SeMdMQWLgsVKttfXcry/WXgjfCTvm1Oi7KymUmFUXH9k
DrHiwL8WIFat7aSFmxRA05WzbwADjXzoW4HP/zzUckKDkXwiajpOgTbvi0I1b0vb
qBezPU1JlHAE+aQfPYRerbEAMh2ySDuaZl2h1mQTtu+o1pMpABQMlsXFZJKo61US
xiQJMAnbnGmoKCjY1n1yKPetTnJ9rhTUqjihts0FIUndXN/qYGJ4oR31Cw8TLaVe
6dQZV3yURLajg45l6eJPGhm79KE/NZgj+NZCZvPTk0xHlfYtis6m8Uq2pxa6h5X2
RiS9ktHWkhkruDnYz941Pwc0b6tkU+Nty9x2c61weIxFRbwQ35zQsBDfO1UANwPb
OE2zJEYHbSUYJT/Kkc7HKC4PQi2lRKbtdEL5cpJtzrwKTuXmoVj+rRmw13hjJjhT
+WPH1+8SuJbiEMUGDzyD+CkwJiKzgjgAdVDDReMLjpNmPpFyn8BBQCKNv2q+1/ra
GglNuG91I4iTcFi3CbV8vptXb7MosBnqWsf0+3zWjHmEG8nN05AuYc7KEDo5KpZI
dDowEdD3lul6pgk4b0DebWK/Bv42mbdKJy9dYGqXfWJ1062Txm+s2hE+1DrF5Wse
WfujmYAAXtHx8+tQB2Qq/ky5KwFHhz9JAKRma6kivf/t7RatzFqEsHv/d15XcOXd
TvbU6FCcTeQZWkapu+nk7++aKAkyNP3GhQ1Xp72AN9OC+nTXAHjWmyqW4Q3ld19c
pLkwjlomLFcd3muHIURYn9tKjGQh+BzEoTYW6Lps7iUzaWr+wQ18P1Koh49PeAjs
rizwvlO5pEsKQwK+C1baSCl6NMk38lKKfZwiRhhGAAEXcd+tO1JgArEgVK4Te5CQ
l5OSKyUFS8f6ZD47GK05UOx+xj7cTZbdtHS+0VwuizAXQzdYE1Mnq6vvUvWwxNKr
yeWskwMZzTa86bvmXUlHAEWgCHgGnNaPMY5ivLYXKbmhI+rTDZsaNJLuFgEW4mNp
Z6CkiQV3dzh+EO6CQfB4b9WSVKHhJWPyYMK8zEG6hiRMjdlu2OnvH+bP6J+iDsrn
0YWoEFNSzBNsVHAfZYukvXc8RNghLVYQw3fDTLgSfHBKzBOPbpM9zZvEVGvemejt
1oZ1qswli7b3rllVN6kQ/BI+XY+0y/XnzfcQADEEDVQ0b2yUdKF7fkRoK5K47k6S
zv3pDeRAmwjCoqiQhrL6/jBm1QWSbPFFzh5xxdr2ww5DDNKj98IvrCBc0s7yYd99
uTH+i/k6HJen5AWPToNiFOfTftXctYppRqjLIa6N58+6OS2AKQX1o4I1LBtQhdgb
9fQ/wJefJG0lVledVUWdrF7NJ0HlqJrxxHdlrp0T6LG6TGQJ8rBDrmdS2hiiST2g
+IobgKsWHGDcbugbrpj2RsBMRiZJdr7OWxO+6LFCBoCm8HjVAbt+AV4YX5d0nfTJ
gh6QE5rOMh/cF5aTj9KKPLNS2ZpF/I2DL66F/+juGiL72Jp/vFmze4cFW5CaEqlj
UWeRHbxhUuxPU7jnWsGR2nmd2Cc5c2ylGi6vVS5w9B65om5aytLo8KBdjaAUEBli
1ZNtnNv9V99fi7wpU+Zdj75cqEk5tRJMUQxY1p7BXkt0G7xuEywqFfjva3KM2TOg
1OEJoLQ6o6OmZDGZvATrW14NhV9McxCgQIGRQDHpRKOKk1j97lodhuVuJrLo3+o3
fN6exO7tmhxUpQ7r99o2HvvucsV5JXW7Oo2fPh1siz0mMTtaaQKlv3dbNRRvwB9h
EG/0L924sVhSNTWd6kkdfvfUXtEWUik/gksgsFy6Fx+YwKHZyMy90YrlEZ/lV3ja
OmQA6HsBgBtlahRt+TCBqr/o8zfoBqY/df0NxNAOVR6O/q/UAJ6zg2WeVYfwWpdJ
bkadsfClKKmUuYIlA77hn/TgqguSLzjuXo3uxjnLccrUgJ36ixD1fw/6yn5WNN/9
bfXD5nqdQfFkQtffCRWBhfbtXGvAWekZYXthvp+YF1PVNxa9BpEqe8GRonqdNTtX
HLFp4x9G0vjx5TcTqr0aru1N9Hr/s18pk1eOUDapO71PoSh5tt7w55tHU+BdjNy0
e8rPW9SsgbenkazajES+2RXnnj7K4BgvrEfCZ6eQJ5D4BRFh3aCFiSjmFVWFjp6C
SXhiCXBDymoD3HGv3/bR1SwWihXeVrGmDO0LCFSHNj1F40kAZvhkbT5lpqlwOyL4
wBCqa/IX9zPV+FfWisp2Y0WXjpMOIuqKC52lclm3GmR3ju//nyDJxNc1O0GvgJiO
0j1pmhQ1N8hW+5G+epswvfiY9UMg7SZJMczfiinpm2gP4Dr7C/fh1nGPqlP4oUIu
9Zd56PU4xR8wPDcAVD9AcgIhhGDx7VYig0jWb9qx6xh+NmNr0p1pm7kHDdX4+34m
F/ShwSS346SroNgZq86d0B1+Q89kcQqeXXumjEdUMyrRUA18ga3DfglUg9iYhU0f
bU3md24RwHxtTTsKnuZwYuhZNdtHb1CurY8go1k8h8fJBbtyBgn3MCyQ2GWRu1qt
PN2fx0KEp8rfZEofzZMOb0B4UMCtxs78vxCRj0GIuJq8pueZWSYqstqvwn4Epm7H
3uZJ9gu5AUsDdSJ2fs0FbaaI7Rk0Dxz22KHWu2Sg8R+51OGhLyk/JvBuj7wS+0Rk
JEdd/NeAGfqAVxl8YurprSw2fl636aqeqyhwJpZeEKFvBioifrYIZChLvjZTxpLc
kDKfi0g3bWC60Lt2ghs0FajyTplJcYKzMaj38NFscZzKnC9PaF3esRIq2Q0LwWsX
4f4DV42oXqOy12IUdknSGPqXoMICVxrbKWk6WJA9wQ92Lzvj/ybTqw4wxQ5qoKmE
BG1eocp0iJmbCDF18igMliL5jZ1kSsgk/GGu4PsNErDr4siCf+qhcGkJ3DCtQysz
DLjXma8qdHhQSxtepnLJ6h8s74kxEMfBN++00X/RYhGQxI/xSbiPAlK6tqUyIU9X
R8hP6bKROAmhVuO9GV3gKIIG1FSbyf8fZj2cJQdNlk165O1oTv4uyuP7FCqzQRaz
L9chHq8+RMjirJ3WAEFENbkJ4k+z98twCehJn2Lq5Dyh46/xGLjDZTIgjieRoB8h
cJ1r7aMaJD0RbNSeh1owXNSCqUkEgfcFYIzFA4b6NSpRk6SPxx1YrSKkswcpqVHe
RvVUKBtDEsinfayQ+AdgBSksqdmD2rtF70qQGmusQedd+d08SZSFRjO0zVHKh7T9
AxyQtcrpGp7zvDMiPcLJOL0iETPaIXV8BgdBuFOo02IxGPhcIJvD1j3oh6EI1yRZ
J4Nsgt3pkjlTKtmVq9pdLm1OuSQREW3+inoiCzXahzRYPC5sxOdUK4Zx9W5LTCQg
cqqD8lL4oVfUqGsVDVrFjCrkgY3cfh6kfiObEigfgoK1EWSVFejH9z+uxRRwmWKj
EmMSUXexM4M21RHM8rr+P5kMgaIoKzgd8YaIj/wJfixOIQMVZ8tAeIgExXE2b1SV
VhHIRHSD/90bC25Gw+QiHkYxyC+CH3Bs53ltr309LGAgFf6kJ2NOc2bDjwI8DdbM
lwjANQqmgzYh9wFXW7mML4O95Ql1mHHcBgHPXT6P8A8Qpjz/T55egNxtfAH0bj+o
YT1IG/WbsYwvuxUkpTwGiLQQXWwir5/iJ7KAYYq4RFEKKBgPmenYAM7YyXky7Xx6
dkMJw7L7Thw43Wm28pxjPv2skW3UgGncpV7hYR4WyIRPc2vF0PPlcNnmfuKnbV9Y
12hUAEdEJeuB8EIYmOFpbOmTcejQgsPEpC2IA8ZhyYnIIEcmbjLgOLv5zgHMR4ud
EiJaXrRVlRaAhJegbH276hXBY8ubE3bXfDy4nH5VGWzoJVDG9kIlP3dZ+DpOCeHI
JtuduxW9VErOSbzqvHN5FSQYb1fshmT2L5J0UrjQJbu/g4TU/DqbD0CKfPVGwJPR
1WWMb+ex2/LdDuEYdWmhpKOd5b7sKqF4kI/coZwHNw8SsOLawGl9N1BYKmngi7m0
ZUzy86rgjrFIxe1bBLcPNT7Vr8X/kizFPgecmrpuqs1sdyk9KYnTyfcOPjuE7lEz
R13TEOrfKEd8BrYuVb60GBFM5FGUVdJLP70SbajzUazzMsrt9MdwjwuYZ/e23rL4
McZik4YMCO8M5Sz4SsUUlwk/ivYXemJDW/Caqn+wTa64OsY8LKh2VWLF2bliwODD
wiJJy8VwalwrTCQQwD4gKodRhKDW2MMEsJmd8/S5PTjR8Yl1m13p9ba8IhJ9Zok3
GV9w88/ovBLh01bq9x2IjJiLxvDjiuLCnq/bb9jtZtljhJXI1RAvrw034xBCFcbS
j9xy9F8r1FJcvztGYdvAHxEqQf7SDC6PvO/BX2LOZpqYn3ZkXW5V9mqC6qaaoVr0
qJvYVTEhDv6cAadQWDqCZVswU34j0OA7dxnhViqx8LX0rRXB7y7DRulxC575/9iH
zjiDCdvEmNJpSxbYYhkV0Bv6hj0DroKrkUfnKwovrqsp5HtuIKgAGmNYtVmdCJeG
9T8ji1EcL8WNYkEoKCrtFDdVImI4hxTkpx3rnpr7xuqpcTRJ2fblEtSti2kgaMbs
24qNnmoaQCO5ujVu78UfERZRfq6ofHzn886cW8b8rnAJUHG+oQ1jSbmcdMivJ6jX
upt9XPto2g8oQBveVujyuT6sO3ujX4xZM9Th25kM4fbsdj9Pvm3ruaxGa+9kWDI4
QMwZP3EA+3qHw9cto4Rh5oO+bJ0dSkFfE9tfdsny7bcR15U5QH8jTyqeO8/rZD9k
Vcci6saxp/bn4M+7k9xJgEwBZZJSgrDKhnD28L4MuApCXyOAJgGkKECUwNmBKjZT
2f/bI6YNcwWJv0+3JwDiNiA+bHaqofHBynkgnO4RDrDPm8OTccELSZxs6O8AhMkZ
AOFgkMIFOlE5/1/mo1P2iojM2tJkhRycGPfcJinq2+wr5inW81tcD2NuBqwo7Nlf
B9TO1NYZr1R7pAIaAiCmn+dv+MKMriYgXnDX6irdnJmMUbuINHiNNOPlvDok0LgQ
qar7O5BMNNI5/G8clHsQMP3pKVnRepg5zCWAgreTo+R+BiupxnTghql22T/4/eJB
hwMhbyx6Az1dfQCFlFCYuTs+IdjblKi7YKF/m4mDyN9xNU0NDb0DhpOEb+NkASZL
lje3s2pP2QhtqG/vojScoNVPyXeFAbE3DKeBQxaSo664h9GNupijNqmbMaImSw4n
UW7TzOX8/E1OPVo2sHix7IYnWihn2PFrlgngLa6GqfCVoe8YQjgUiPV0eB2OeE6x
jA3q2Ljb/rsNG4vgDmAVb/i386p/8aSd704o7LAiYUnjWngFOe4JZWQ+wSRDKKeh
f/yNTjNk4Fmf9HyhG4+5VIvOg8JnxoFms5S+zVQkx4OOm4/YVd/qP9JAhE5RRwbg
49EKTUB571Wj8vXiKj2BDWF8BHN4ZuWu1++N7Z7f6iFJ34nVKUTMVqYbEDka0BRY
BMHW+Q4iliMbBrtqSheJZ3cVIlhiNtIctOpFY8Sebin6Ep7uPSOL9KZm38/FT7Mh
KsDBV/sdTtAjRYeGtZlfWGOKLnaWzl1KjN6JHVCfwo29gv6EoIXYAn9OYHcJc3iN
5F4e4Z3l2NxiFDo1qNNFT2T0CExD3tWmAQncfD3QkC4hv9paarrd2c79HKsQOTuc
OrnNsYlmQUut2AS99dn91KuRY7hyLp3vcYWiVsaiptbnXM5XiwcsE90NaZzEWmeE
2te1Y+fjEAIA3IeQERGgTG5v39+m7bwM+dUlR0002gHZrODBDIHiEORdVh0+iBPw
6KcrDdU/zCM3DS06IJkKH+SgUB//qgKJHMt0GEviw3glTKmJPpYdi/TikFKm5S5f
JdrS6Pll7jshsdFXNXt5bou0tBKmrGhjgQRrX6JHrHyFQMwKpaBGvvyulc135URP
SGi7Gxe6C7iZrk3PTqSJMits0OPabPoWqMjYrfBsfw/s6h3XLaFhW19aIL2YEnVW
ARc0hmcqapic3x+1Au/OyqdD806voipkg6oCtBkFeocRLic2R1h1YnFvptUTOvHz
WJD2t+BHabnExxWl0hwbE8SIQN+Uc0HCuy6ZZqbDWE0NQsMvCEmeMzFe0hlJP3rw
VQw67CSUolgvfRSjKUWyu3stQAW95QvqPNuPoj5lL+KCh+7I3k+b4NvBm5IHwAfa
7xp/9pPoy6WWS2pbqwmZAggtM8Q61jySADVRC+xFRAKsni/yn0fU9WfFzTeVtKcr
BUN8IQWZoW7LHBN0BKHR1JTrp5t8iEj5UscoQuLfXS+kpvSDKobpykv4x7Bg5d7u
0VO8UL+XvZE3RouxSPmT3Uk8xDkWfICgikLtvjqcSY7AZNkb68xFn5YrTRfrdhMC
c7l4v8p3NHPASKe7HeGMEVSKWOBU3V2i9fzCsJvDOd0JnhJJBJeTae3+rYa6ZYLC
PmpwCxIIa9VfBRhw0mqiA9FjvbiO6aY90GAww4WJBZ0IZgvbXs9yS2tlLc/lY6Rd
Oc+bNHkwQwutfH4mVDH/N0JWn56EqA/pK+hoqPaxXcwMWNVs0MNlBH/b674M1r6Y
FEjnsOSu67nl67sc127BwagMY1NG9N+zu6OeC18HNFREwcy3IYtOEeTzOtT45iks
zgy9eAHa/PNgxACeSM32CiafM/h4XoXQobyTnEXCG+zldCPvicfXCY7oiyxLNFd3
LaStB6dWdTLzWFmVvkHc6k42SewnCj6Qeqx3Oz9ijEJYPkzRkl1LoDgnnd4WbbS8
1xbexAnUyKy7wcD0mXy5QP4v1q9/REwosv/MYxNBBd+9dX1WLgL5qqWrlzCk+EAs
ZmQQuAiClB4H1jkmDyBxtXC9k4gdo+CIoi6TnGEEGMhA4bl1wyO8KIyowLnALk8E
qq2qkktSCmaJPsTDZJqxL+6iRGyOLK3BvxtncnxA7b1G6+pq5d3L8b2vLmXWRxh+
tVrP+xc0ihGQZBaloZwOkjFZ1Swz6+7uIO9gRhYhT79tNSf6cLeQnsu+Z5Dyutge
gY2LxDToXGjRPCBfwNlevr38PAJD3TubpPRVYqQ7j4kdk7gqZ0LeIVN8xhBtxSxJ
H7YY2826OUDBkr7OEnzfed3kK7F6WiLhgUHVndo15hxwN/fnaXeopDt+VUNp+5+v
9NQuHRy66/pVTtJw7bKO1we2nfW5UmfIzfzzVPILjeW6GrU1wFQpi28VglNOwlTn
onI623SuE34zGiF02UCrr2IDqmHAk/Fh6R6naxud9utqvOAxSYV02HUTU3QEiuw4
nWicVWvtkZxoX4HnT/9kidbki6RngoV/ZhDZ/BTEVkT8aeZp7FCyucejOnqwEZQG
kAZCkwK9w+xp55isMMTcgYGD6Iwq9aYy3ZiwCGVhCasvU9wtT+eH3rrDcaZdCb7S
RCIFa+VcirIBxt22vLgYegVTyfulAjwhX87gIE06Pv/Wpgfuso75Jf5Z24CrGSO1
UaaKq1xwQcZ1AV6aopJ4Of1NpYG4gDxGN8gx99XhkfGNsQbSNGMCJVie/BBqLvxW
cciOUZv96Oja0AyWksB2iQ7INCcyewlQH+3dDycy6l1kbjbb7uTaMKfJKa1pc/kj
JxEuDyBjK/v0rfDVYyXRLBGtTZGh5nQHBHTu72PTdwBjDfwS9Hwh762TgtNl0eZH
Lw/j2/Sl7vliZxld5heDnHcKwtgYgQ5A+CS/gXjJ/G/Z3SFojTHgUrvA3sgCgjGN
hE4m7xhowBnugD/lFTy9BKIyU7/7O/5kyf5FlssEUkKr+Byx/81xJkUD48bmr99j
k8/tnJwdicGySOCTDMDWb+AoFBpu0VoOl6ELoomdrnyEjehZ5k+//FNhPCOuqB3F
2Z89Muhhu7ir2Fv1ZLdZGjPMCG9llQS4wdNr7sEtdl3veMj02BjQndmc6NtrD21f
jldgdrMtoqXl2E3Rxk/ajwcNu7dnJziGdMscug7dMjNnZrErJco/kiHUxlYC5UlT
P8Xs4fDqA5+4b4JvwE+lsdLUVxsVArD96gG7t2a4w9cRlYOAg69CDI+ExK+jMipS
peo5LwTacz2+H79RnwDBx3rFtdArq8fR3Of6xeNAMYjB3veXpCpD9quq00qUXzo4
Rb2eijun00HWpOYodycvxMHZEmVVNq3SdbGpECTi+4tfrkAfl3jKivSccZLKNFpt
BeGkTAk+YetoCApJnE8vm8dlDxOA5jtpxSv+0YIlmJKZg/3paL+z27JJYobZyiui
UnTUPPov4XfBvG8IvlG3r1Le5HLvH81QWOAm1PWfrGbc8UAl8M2zPDLclRfuZ/i0
QBu2OHE5Ju7YYC2QTN8rcE1d8SSJCjtDSgV5Atr1PudFyLt2+Bo+cjmsMckibotT
UMvubd74QTckRTKry1Op7eSlFOlQ7628IryKDSKjw0LTbhCG5opMNsxOgh/z/Hn2
nO71EQ+XIzvqq2gQ5ObWDB98NxwuEqtj4rSbGnfy1Spe/SWeBT33GKN0VmPq1s5p
sLpTxOY3P/Oq9UB2nT1nS3lIUCJCJPvMQPubN1WgCkE7QWmvuktnq9bycxjWQJ/H
zpd4WOknvPNJWa2iJ5wz/F6M42EBY6GdVPAto5CDETg65D1sXXuiSzNK9hN/xoeq
EJ3tNm9APyGMyfo5pi4SodQxfP5YgJNFKJkuqoguhPQQHnNCTvIt7l3gSZrBp2fx
fyEHtvnTD62wgcXSqvm3C8t4k5kydyCIfRBBlpAoHMrYO35TQ90T4bn9E/4pt6Nu
HXYQAGNwLMZXLM69HqM7gsH1ZxijexZEzkRFWnGRUXGdPnpWVKm4UrOKQI9s/O6a
XmUg/1aHN4cXarpV0YUPeaJrwgccO58fxdamjBS4qX09wy1568qZG7LWKztqpAOF
QSEbtBws4wROdoa/39CJRQ1p7Vt6cRpBGJCw4X+aL8VHYf2ufMu8wW5wHYEbPuiD
x5rxLIIws9cqRHFHRH3RKnbjSbHSDy5chShFauCb7J3vIqfhNszYHCuV4wSP82qe
X2685DvYKL7M4c0DmItyz+y1e4yq1ShL1U9vZ1W/+OXZy8nsiDXSTM0wIX3tPlU3
ddEZH2A6RxdGWZ9oc0b1pYS5XTr4x25tyFMaTLHDZbOmPUOoVtaJeteRziXz1rLT
D/225uWvo2+xLfXp+jphY4cZv2qHe49FrOP+NUN4yJzVF1++8GFptUg0cB8iwk0r
y7yGXFcuUCFc38SXRawdSqFYUYWtlH8xDxtlVltuaHghjAcHmsWlxyGnj9Pvu+n7
j6KUkqmK4xaw7cEm4XG7bK2WJWRgYozlqSF2/VudAXx23tH7jgOvbEte/6hhtIXm
Ai4Nf/ICjqOYf87mOAn4j4cHwbQxH7yLyLy2E8N8eBAy88azMvdsXm5dWNAylq8J
MUAem0yEiQ4T/bnwe0NDvXUBi8NOArxpAVM54x1FIjN/INCljSf6VKTZrp14/sp2
DzLmMHfkvZgft9Zr6P4b9RIZuOOy9LmdTHMzZRjdyzO+Yw848hNdM2N11mzWCO46
DT65ajatIFjCrMq+Byjt/5ohThbLKQ/Tu5PHQXYXGAycPtK/CgdAV5pXBQp0BBaY
nj0KvVD0ZXc3B9r9korX79/T0z6TqVBS5efN5wo7tjDwAJKpXWVMtR+OOWCQZnxw
8h0DVRKinMIxOL71aZxftTpIp9k0zsj31Dw2SZGeqGhs039quP/R3vgxly2Te6P0
I5J7UIvO5KIwpmDCgH2gJfZdVrkxq4s7+iqI7follDuREXuudiJ5uiOn7Vp8NEYf
kakDyDoYBQBqOl9+FoUWOL7q6hdVkOn6j1yOJgj49QSGBXj4hSddrgSd0THDHKh1
XdgdAFheyxTVWF+5OYxgT6Z0WraoXw02AiBW2kcEHYFZU9xMHYUbzBM8XrFlOG8v
NPzagIbEly6PX+qleX9ezwq3f4B6SQjERiSIoCPE4fZcnYRq2y7s8tKiMsf1UQTS
Ai17npVkdReedvWvW1d2uz1KAJK61Ocfjj/MaMaIxzLzelibUhqRYuYxNakCyNMr
z8Gc9QsMcdsFDkcYvDLldeE+oiDu0MLRI1B/Vi12Qecy/x3tBqhf9FSfXHZQrL2X
lU9ZskiDT+MrZvU1eqBaOxC2R1sfKFongMpe7LEbve4gtOT6VK9Mkgjo3+poKb0X
xPEZJNw6todZSGkkFwEe1eWgvgv+hIc6XFcEik+B+xuWgv9He9DyZ0XqmuPItesu
slESmL7saDb9+Z9D0f+La1BrHJRTKDOrEOlSMFMfkJOid8Dukf72g732L//sQ7ZR
2vTrTYuAd0Q7WRA1ypoy3ybMXjae1gFQn02jJ8Ny5yhc/UR0FWtmg4ugsCnEFmE9
2kzqBWJZI55IqpEOWW08SblDauqTbjN4fF4oqOO3xqM0hNjLxpOASUM49ej8zAgM
JBNOKQGfGiaBGiPMQ6J8mLsyKFGSE29eA2ucoH+jpxfzWu7JHBSupzwAaRuuqFlN
lIW7H641ALcO3OtQR0nd4Lp3tcfZaMpR0Gf77fJiLT2XfCrsmjNBRzbrTXEWFQb1
hBiZ0v+yS65CLPSyHOyT0ak7sqrSqe8oOlscuwfbKBRDYXinTxT+mM2wfXMD0vUC
uRPVsbSKqieUtz9I6pqh/LvO/v+6VQAEv3bCRIAXfhdlD3/fXP8v+rX/tY44hDru
cd2xhngm/vPb0f9DAZhNLg4oBfL7srYBKNjQ4uvvmbkSgHyOp/d2C+S13qRAaQ7v
1rnUSKm/BMFsJgoX6QxkefpTHSB7zlAgXaIx/oCyk5ClsYpL5IVPCEAzYcsDh8XH
yKV7AGFoRY63qANGF274vnM1oKal7fAf6JrpPYjS366QQms1q5o8LkRjjBZ6ytvJ
3R20DIbrBXqHqfYlup/lvZ7EW5/uUZ2NnjJXHdG3zlkwjT2f555j9Eh6mqwPiHEI
Qs6B60E473hCIQopX4LlQKSaKqS2OCibXKgGoj6Fs/OgFZoUOVpFAg/pJyootOt6
2SpwxuKUmbtCr5twcXrdc9RJLGYWA6q7QHuCac2ZMI1mnB1+H486e8kjgGRuIXS0
8pyoZtRX1axpamqmwxagyhP2z2F4fAa9Z24PZdrvVeVAi3R9jJsCEN29UzhB65Tm
Ji/SieEkCtwe5VXTRds9hzBUjsbz99mtJ6f5ovetdTyywZjk5i5WinAc35GBgTdW
sdBJAsXuU0cit066rrD3lrSYYt87OG9Np/zpsF7M92VJbMsoi2k5RVcdLQ2KkRJs
Y/mkg/Zaz7hQ7XpEBOcgleWwhgaWWitVsyUm2741ixH4R2FQlIbOj2DO+UvnK3Gw
fQzXZMxQQAIQfmM9Nur/mqa0c4pRDMWasqhVPrWuTq/zyU8V3Lx4apRBeQKD7ixQ
NYr/HQxC01/RkyXxC/PA1clqkiRD8sxzbcbeoWyoiSG5vhOs3vfnkgzw2Ch3ApP2
by+kWDWSOAzO9s4uVXad/82kuIJWXIFzliTe2L7VQbGgdspfknjcU7xA+oXJtR3l
gYCT4uDQNYNnvA+fDATipV7S5ky0DH/vh/GR59g4lPkuLfHrzaxHXYM2y/y2GxWX
LPWlHq7jNS4CYKuKWPGn/kQsLxhiCoEx+NVEFeqlducDuZ43LKfIpD1UyfYq/QyG
zdV5m2VImRP33te0sYDCTLDUuhEtb90x7rpEfLwmHDE7rWuiiCGtNfnkXUFQwjTU
c7jU+uTkgSIVvkRMstQUAZg9+ADTtkDPz145eh3Sxuey9OnpxePPV9tVg+FQyxxE
JgyiCxeIJh1JgVMWY/noiq1SoSD4s3UKUiUinfaE/cxZdFvIUiL95GgvVDMx1Bv8
OV5vjLs4vtL4s3R/7PkcxlAKcsJsOTpuTsoS4IHGxt5T6LQfEAx4ZtGh4YjBTgkl
1R8Ul9WWbAHQ5R42M5Ynzcq/k/3MunHozevook9hRkI9oaC5W6Jbe6Z5iLLpOE3k
lu3IHn1XUVwBBh+9BSMUsSlLNyqs0Gwpfbphs3OULE7+mG3dCcoTF1eiOKvTZP37
dnEQfmBUbXKUu5NZYErpQtoBi6OVR9BsIcBbXuq1DSnW0VvwJ1c33nHD0JHMHQ3r
cSW9c4Kveo7wuBtamIfEHt2jpyJ9z6p9YVqAhV7mbvpRKoKSK/q7pD4uOa9Rm6G0
TzbUgkiGaHUD8mDVBBgkvj5K0q2sEE5HasvitFmhC1FW55ICB43cYJL0iW9pbvQ1
gfoTmHt9KiaYEXcI5hBUirVOUFw3Vanjb7+uY5SCHZd8V5ar0OsIKR0Jurk+UMCy
sWClrgaOPXtMKqnL9vgvvRhIsNmcXqtJaboFz1wpDD+tmiPylQyKiJx318/YPwTN
k+jdMk/lNAW76TztMyKexE4LqAIO4QNVtWWXABoSsXrIheNxBvYzu9lVVmb6HynP
xXwL/eVMHgq/XHeDzm+0fzGMNMxhW1yDpL8VZg1xM3ThI/KKeZgEFz3RYvwuHwAM
gJ+ArABkNmmQKCn3rphh/7OOcD8c/aeLPjZuBV4QNifiIcr8Pnubh3Yct0PgrDHc
5js8TkKm6acYNne8BX1OAZThbyGaHIQHphzvmKahyKtucN/ubdKfKPDX4BdMSahu
irfoXnQUPu+TrA7eT/ckHDPrMc3fXkA1AHZjcFhrzHTN+vC/KYNAdc/6tH+uaoS0
kSHNqQ51/YfMUy+OE3Vp0gVnr84aItzJiIPXfuABFkhJNroCRMWiugNKJ4RIXqE1
wulEL6WCky9UN20elBydPV0At6aoDtaXb2Pv3YKHx47YhAe7oXUgPedNDfOqC+Bc
40wj//KObEtWyzwgF2BQxcoGGn+jGcR1ci9YGJZ7AGc4H5tOfmbc9SGBp7un6O0X
iwF0eUbTT0Dn9j7uVhdDmrS3F87m2KD8438HMMrjHEC6Uig/DUWZ2GEINGswIK6P
fpchN0aGdOLqYgyFGprdrpYHXvdX5Z/+ndGm8TGnHtdAVJ3j9ufMriXFvr0wvmj/
xjdksCzlU/ngWem6Jhbycpz3exTQoS0tmAXkUAqh4Lp83eWYpqw1dBharA+URUmF
ypkJAUhfbEvdsWqAvz7jxlaOEDudoIomBRUzPVpUINUjXxvdz/8y7XZHbyiK7cb/
tKfUYwSK57dzeFsztpE2jclJVheI9aL9WaHuxX7/ygQsQWzMDl9+8UZham/QZBBG
HC8l0it1fSMWvmV5amPKh+T6OAt1QGg1KxXbJkHUA5vzn4mx3F6UhRbxUoxN2N4B
zGmeGG3LPxaWGWUc+BiFHVbW9emu1NoL00Us8J4PcjhUtBYHX1xrtLCSpVQFz06S
EU8yCdtJug6tiX81ixpBxb5R0GhODVfgVTV+iEZkvDJ6yHtgQ/O74YFnYtS3EdNe
vLNCT3nuNZWwiFdBlQxuptuLR5dwChEbGe4XgKfkD2co52xPlXabbZqCmZfLdKoV
LmoO/QhG/ev7B8P6/OBy9FU0M7s+49NfvqPCoZNI6Y7L8se8c34XjwxJMIkgebkX
oN1wUy6G9zYTIxlddCf1vzi1X7raw43armvSGQgJHFjjpW3aczKglQ3vvHdmLXbE
d9+KIVY5joLLLP3B+2xw/byYMfc+KRb80YFJzHIlIW78lW9LlROppoqXT0kHe/VR
iaJBorEI5dnUHSsrsEYflf2K+uKKVnXyXhcw/8NWuivJn6MOYcUGo1eIMEZDnhM7
IiuAgYwwitEuyMRcDSKf7C6UQgR7Qxqph7x6eCaDmpw7iNy1VSFGXYsxaZEY0zPf
Ex5UM+SN8fzpkfHzlmOkpzyCzBxKhxGBe6DKDvnYnEOpx064t5Z0zUZYZtsPL1R0
hxm3XWs3gHb8mF/CmmSw4bwzaWAYF6z8pCxxbrB8S7ZThMosyaDwp6LRTQMtJXya
EdXXNAf33cj8X+4iJW4nIM0IJP9j0OZwjkFaADYnZVxfQr/qMmR3pmlaU6Tdjgyq
ETLOyKWshZUj3tcIHgGcTDmzUb4EIGuRlw77/td91kLERYZJRyHJSd79o2T4999P
01U515F+CFlbZXQmJWI9EHmG1Ai15skC3m9312NYfIRcNOiKwAfIseNktBCIec6S
KPtNJ4su24J0gKuAYAoRxrb4uLnAAdL/5B5aV566vWSbz2gt/IJdnvlHPp+g+I69
u59uifx+iYs/h4rg6HQl+kzfNX7PIQrzxhGNx+++ogcOqLuXxoMCIWQXMjzg6VGp
0I9/IhAG9Dh4IJK20AAKlVQHWCWwjh6Zo/vBZGUYIyfGvhIGgYWm2+iqQsp0I53i
aaXDN+RsuAPNuhyU+2ZbQ6gV/4ce4Uh0umQCmgLMyc60lPtW6gKiK2xmnr9xMTeq
eikWJfUvfaN/NGx0cJ2r4pa9T7TJcSYR/VXSJ+bKTE83ZyZ6m1PQAfvbuavKWyxp
ysp/NQ7dBEZW9tdLzS3TSN/UNabg/+pw5JlBvbpQ8DGNDe0gmx38OLWQRlUO6FuC
TUXOo7VjB8hMHynKc+/eU4JObO1DinuzygYyfk31mg/uhFmp9RVKONUEfO36GyaQ
fAas+4+ebJITPk/ygv4odzrTHYnGZNZW9QY8RHITlbcUc1Z9/k/e3ZScUouAu+Ji
kEqbKik0xZQA7WxZ1NNK0anNueSp4PupQ0MawuSZaswRrtp7csmK87M99k9R/G2T
9r5GL80YiE37pSTzF7G4XEUJggiwFVpgsle8TmIbs33hQlsjP+Cwt5OAM7hFBIjO
hRRKaAOjtg6cUNYGvGIhsHDNSuNV2NszvDbZ9sfGK+2V8zU6Ls9zdPfNznqK5/TG
zl/+EyCaZLKzWlibn5T55GrV8gP73mSOyKxN5PQmDPvSbCrdic4fTP+DdBvw+myr
oQ9xXNksffVlE2t4Fx4LjiqeQi+FQI2TmfZt+AlG0UXlCQcPzd0Yb5y87y4PYNeC
drQrmiv62AjwHIIfra6RQViNa1WYbKbf8aT4syKJUsNaQLBuvc9+0x8cYZf6Vrfs
hFAAMMOyZm8tF6siKfPixx5GAg5NkYkF1pl0eNtaOiweS8zMhvcmaz0xCQ9notUa
uOz20pT5V+3nTNzs6MZjh0+arTk6sW2Zodg44PFoqC2qQHKB4EJgumymrKxJKwKj
hLbpohVKcIguaMN1P8ZgsInqbMatB0m6LUKwMgdZgoVxcTWAMS9KR+xtrftJNwCa
Z223QDgBgwK/iGANEN4w2nWc8trK9gJE0V+L5KpBf7IwTfIqEin9u1uZwh4G8XnZ
QoQk6qZUgj9QS4LbKs2lGKXSIafKhQIr3M0+qXQZxl4oaKensKMmQ676UvMh3SCI
WE1vM46YhrsxQ3ymIlRsbErr8JQfTs5ws9TpDSMaNM3t6Hyq9dPUgHv9DyqEV6xw
u3UUWnZfajrCRaAtAK7qB0b3XsxIdmUnqk2uvIom7xIpn0WG8hmgUmtwZ4B5/5Bp
1yUGdB1Zs2dMoaDwUave+O5415zbkbsrN5CxLuBEVUcxT1ZLEwpmn/hvWgltmiq5
BbMB1yu3aeXcuMh9FDyWjBG2S3RVmtf9GeZOtO1JdM0EEnap6xClyK/7fI7pzYPt
+dTSoEoZES1NSxJeNT0Uyn4p333Cs+Mp4Cg85DjHKFzuSy/S4CGQGGeTcKBF487S
K3Ktqd7SgbPWB9xHJqe0OyTRNOoANHOcrlBGYDOeoA6aOTnoXt3zGb5Q/gynVJUo
ypNPCkK6ZTmTF+1Wlc9c1Zl8OeyJGsm3/AVj7ZbIlCfziN3VlG3CbYGsJsFnwchd
sXFD//lfss+rKNL1+GvN2e9l+q4IJutItEnSRCMFyKF92AqMZwGWC1PbhCbozOcB
rXSKbmae7qqUfsFEKqPx6MyxFqcSOln+BrW2yzLAOo4EXOT2y3SA98yYpc29JgBT
xdpucogPhi+EW9OUOH/SenP2+1tQyUV1und7VdGMv0k7hsU7h871AtVhV0kqyn9p
FGZrOg7Y/GPH1KR38RiDhho/vSms+YWATjXwO/bSe+AxfXZMiRHh3mHPpPdAUE46
SB6tw36UQsZ53eLnGQDzESY8bPxpa3CR9XcE6JfkzxbGSPI+wmw98HUfhQvFJ6Ja
QLm/P3cMkrmTlBz/GFnY9Yp/XDPchHmd/OWXUKwTgvVeEY/wENhps/osyTQ+KqBT
m1WmZxY7bOnXxPfUvkEMd/Esrd1WGzHIh0q5UKySBZlI+H32V6FaoCa69dXzZjbR
OJAN4ABszAqTG2asNO7KhVwLRdgIqSog8DZBPdwxrPesx3LDfSyEa5yZ6A/m38Vq
1J0M9WitsLEQPl4H2Rzp1kAHBimb8u0FsermqIrif8TXvEWkSyTFYECNs0q/IWWg
25OhSadRSmLPDEI0gKDaqiMwhR5WJOueicKhwG4ah9VAY9CGo99PaKJN3GAG+Xxk
kMPOj6g8tChyqdS5yUwaZ15cAaICkXcGu2ea7MTP0W/w7DXsX3wkf314UjsxYq+x
vWdQ2XYev4t41cWGZTGhc/YwSiXliBxjZ7O6todQvNxKiZKKp3gSdSYxvCSkF0dv
2O8/fwdVyy85yUTtZP5skAM4aExNZai3HuUVVYbMxlWQEQzN6FFL+AoncY8gAlOj
dokMa5Ous0L/5poQqKcQxNhTWY4969f7qRq9EGsZagCmgc96+LyFhpyVaTkZtUPv
/PakZINAIic3xSTCGqmN16gsyEm+tTYKrCaSbNaeDg2Wc5reEHtaVXXG0Rzgrswt
CTYtTKS8JOr/Ppdojo5FmhvEm2I2tDTyIS0vv2gmzSYlKW2jYniX4JyIN86Ruff4
peOZTYEcJ8UW5j3F8F1ZmLj/mC7+C1FPf/ebjfwUUo/ZXZXp1KoaqLATwQrSH6wB
3t0en1/yt5ZYHPfShRvHyQPo9wMaAssUqGjI18wm/hB9jGNWLWPMjx2dsn5I8w+7
DVleb2dFPH/62ACY6TgAkeuA2XQJMn3QxPAIruM5A3dRAnF2mZ+UOvtazFN/5U18
XLnFI3DMKmw5fHibbjV911coN6ODPHpxOzlxlDFYUI0IrqC8fj9JxVv9+iCXOtCh
Bz8V4Jsb9nMWeB3Bxl+ulSdueWMfLwzGKsaIPmrQTi0/pOLO5w6G3pZWEcxWC6P4
605BCQI/kf0TkQgLXS57s0OwjA4HF/VHh076ZnS/lkRg/tnQu/lFCnUiaUgTWzff
HRFaj5L9yIO3l6iEkgCtADuoRY5nNdCqY3ZUeaVyNwtt3OTDy+0bDcq4TClfZZxW
PZsfMBitKPJzFtaF0kBmfjxlOfqLSIVgAsmz8UtzHqyxLMZT6pP5cCRPq/VNEGx0
kIk9SYW3EXWrhHqVkIBZgC+MM2Bd1Gc+WzRjfxBtG0UvOl+KYlS6JMCduwg9ZD4e
RfjRlH3LYvmvjJA1BnZ54GnXkNEcro3ap8vKafHaSixqBERlN5y7Rrpebejtq3uP
/OazKO2hasRmlPWUKBOxEOjRzbPANXaZTTB9BwMzvVMj0vL2RaazxoLBkX1tat36
7R9Nqf6jE1pgVBiWfoEAgtmh+YjTpTCBxssHo0DYpA/kw+KyI5rRcB+l0GZk5VZ3
wEOSGXE1Oh0Krrfa5OLmVrXgJC9MdhV1gJZyjVd2srxwfAX6Q903AKhC9RfJeWpR
yckqAfMbGwb0bBoJqNnqREkUYalYoJQCg+hDcqfCZyhM3w624T47RqNEdDXUxMlp
p2FaCPqrsH2i1E1geDylH87+cpOsLPnI0+3tXct1aDCW4vaMOU4I84i2ou/RWlle
cxkI/vO/BhiPjTskFJTRtelwjFBjtGEq9MYQShEXlfVeIzE4InYBTc0UW2fGLxb8
Ku0jsU44pRzJHZ2SztxHYYBO1mvdcRYCPTclZQ5DEzvHEnyHZPs07TGhPPHdWrQO
DAvEUraXb5QBo7La3Z264Q75KN1RHDUxoIrL3mZCec8hKSKX4PRfExr0UngT30CF
LDBRlERuY+kd3uIWxcCmzEk28t1rdbHNMbMhiFMwpaKA4f2uGFc/aqyEVMJ8bfN4
HxNrtLUQXmQuj2bzQe/waiAFG0QNK9kIhp7Os4NxhuX/CfP0/O3ZDhk/Kx5cXlLT
8guz5ItJKMEJyCTuPqYWZyzehVdp3wDvZgnXxWwXhBj20W4MPPIuHQ+DyA4fDMHZ
4XdT4UqQC+Vjh7rXq7FWZmMSq3W/wpt9ULncZFX21fcpkp56cqlYsIpRlkAeSFMb
I3+gfhoq162i9c/jNVFH1igI/om2U+lO3IDRTB2c12vwniH2PtEj+wmLxOgXUBr4
vy5t3oBFuIreRYc+aRqzJ2ZUbFNy8m6VMRMfam9OcgLHdLJM0Cwh3ucCu0Di51x6
85FWk63gIaIPAtCH0LjwUoRYe54dcTWUd9eLSSwKivFi/fwJmJgYjF3wgWEQ9zAC
4BbqocEn7ICMyocuXTY0d+IXhtEnxjhME86oNYlBkKKzZKz+n0ppRn4wFELD4QiK
PteMt88LB+nkERv0TMHGGO+CERUSD++23XEm4oKPY2v/uYaMTqzJVdrUAqrTsHlM
aTATdPgCN9yI93WLsN3jVIetLmy+lNmnm4DOIByp/pmboXsQPHwHYTgXBPHjtJsN
kihD7yvfiIEv/bZjIS8yuJlkyewmhbXImKmnwkcm4zfaaM9eqco7OEP3iSfrrFuI
Gj1MWhonExKcNIxVc7dXdVua0IBJfJ9rx/+UAa3BnHm/FikLN4fu7pUFDMmyoflz
GgPM3dEMUmo/wNgMAKEFKUPS6AvmBKnBNp+F9rcKDHKD526pg2STzzu9HfjXl4Zj
jhWwnn47lB0SXl+3a0Ii6ZO9yWZt7g7SA7w6xk3O8xVOxp8FrkKsZqPVJWeUNe3K
PFLY65srzk8Y22hROvXL/PsoRtljn9JXbCix78QPc6HlvM6Wb8PRz0xCmem+B61U
tw4F3ezcz3g6+qU92yYlzsTYU5r+eSfexwFiC43aD51FOnEwM8i/W63+L+LhSOsE
QQLHrZgTIjWDkZ8QSVGUhG5tkac3Dg9G+t49Avtm5taqsXu9N/hNfTRh26za+B/1
eoV5TWiVjQLgoF/ZysCT8psXdtRHXq7e34koLJ0ZbzgPcIkyeqzizYONWvuY3KQ2
c+EDPMD4f7n0POcmwNZOhOHKXixFnp4EnPCLmlYcUWG78gDpZCqSOWT/1ZRbdVzo
P7B/i7jWr5Au7QtctQXuwtwT4k12aMzgtWT3ljxeFYXmZIKIHD8JYjnjSZ3QSFmJ
MRWrX9dPIOGWRE08RxJv7aCCahq29wdZaFjxsSz6PL+5nvjKKKl989R8BWxblLhr
Fy/dJpANyBf1R+3FW+sZJxiqNW65xHoUstE22BY/y8yslOBAKP8YcCLrggU+iH7M
8kGuaxSvOWKdX4kz/lyxUR0KRDDpRgQeQ53zDznfuAh7dFrimYuRxllyZZJeuzMa
hca3kMuoDXfsLJ7fIsGeNpCUgOFI81kgH5KYA1cmhPqbBoCxQ9qK6rjy2WUoS9rJ
DYiJq6Go4LQRChf546fyUt4EdJjbVsATeAtrOTh07IOsI6mI9NzhjofKKNwQiG6X
tLtl//cXUHcZ+Y2gTvv2eE9CyZO03W+PINtcIQ9DVD2nkOF7/7NDoGT/nL23ieWg
/WPkWQXqSMTAJ2vUioUtwI4fDK/wOXCPxV1qSN2acKtHxZ5V/cVka6mB+P3Uvl1t
bGUxl/4jhZcMnVb5ePUUltcxfGMrJSUlrqLRx5fI87yXoRB59WOzfrijVzAaoY12
Gn/gDNoqjeGUpUJDeKbGxWCJ2KYRtiS6RnGjvYqrjgOUoSodLYp7Mc/3Z6DWAe/r
pZB2DV/3IB+m3ehhX4o6inRqyGxNN2znsg6sCOX5YulurLO2Mui8Xq0M7bHqFVQm
AvECcfSekFkRd1O5qovsWnj9MW2KzyE1bu3VA3bKsph4CGXRAtBAJIZRgi4WpPqz
S2GFHYi/uPDwhu32Yf5tWDc/5uX9LdYxS7O2HkK4++cT86tbc+mdXNtISf6qviG1
RE09gtRssA+3VvpM+mq7rn/ddDjeaSQSzzZLWPRUegfcuPWODLFI52DXu9NkB5F8
oNarQ6oaDYoetU3Vwo0/QNmLAWjltEN8R9nLB0jGNcrEFLu603wlBgPEJC2uTJVe
5QEvPpPd9sU7jxAEOGl5qPqdpX62iMhMj4sQlObKbtRwgD9PKPvE9of9/kcNtFrD
j5VmjONa3kkrukhSa7aMToJFC2Tqzw7Xx/yR2QcHqFExjCaoO0TVM+vhLzohDX0G
asdBiKR3GFnBWUIefNHADLTBAyL9BzDfsgGRiL8zly4oe6c4da3LS1Tlw3Kg01zT
kIHFVC0U+3+zSVCy83rlbDjDsK3tOne7r4tpN49NoA44YFM4aoH9lbGtnCM7DS5N
eTfb25BAMfAcVBLk20DdGKq8W8ruBBhEfbAU9B9HQkHzKkjIHrUuhsezlKdSFVEI
lzBbE/QTB1tGjjtwqagFj77ohfS8gyLWT33Bjr6BTcCjT5mIUga2SXSsCnx9VgAt
ayKqVb37e4nm870zZoqKjiG8/pXghafJt0cbfzfQ/ou3jHC0lqdUE+79C60bo7v2
1U3Yls6isv9jh+Jm9Bfgt50NSg4hhXZc4S0zs8jjoZq4Or/sB86e8zd1XK5ii7/r
5bvj4GCFLOJFciwULPirNhLZzi/O8FpsfmAQ3ymDojZMC6JUrj+V+1P9lb4DbJHo
uABfnKFdmM7VJx3CxhyZH4VeczQRRjskadCa15JdX841Zaztri/y0sAQifgHnWG9
WrFxvFRCUfPkTAqoluTc9koC0SWk7bBKPzzQS1jSaBZxVgERlInLQ9uCNLVGkMVP
IH/OeBKe6jKaLwxUlqdz/lSuM1Ly6tgmdBqJPcRJL0Xhvm9eLu1c0qJ/K38hcoLG
52oi0ZSA9qmy45aTtYxatwt6hpTPAYUaMrPixRno9qttRb6OloXkBEufwVcjPq4K
wj8DwE8PeF6GxJkqBpkDo7keqPwAufN5X7weCe+KFVx025gH4E/egfcussvjgttZ
KmtO7aKy9n+3XEG/PsSCkeo3aOwecW4Wuc/lAKm8JMsTQFqkcs38BVPIm6eDw36v
CbdYJw4fVpumOEmXg5rWkUBI1qAqDkazarXXrZuVkBGF2S5qFlgn0wwNb/bsSfeH
xRDp0dg/mrIFhEO6r52Usjr7zWlDTtH998DzQLQHBiKJTBxqAW1htXdt8Xece61T
iq//NC5nyHht9oW577qwDkINO5RTAFe4UVJE0Im6nbtYPewiXapSz1TqTvwSCsiP
Gup6mpq+00ftsz8ob8ElrIwcc0DA1y6/eK02CdphPJ7cK53/bR90yZcksY0UhVMt
X6HZf4dB1BAKhDtZ88cub+NRqHk8vEsrbgizcl3Aj8BUp+5uMBGLGG/IWK6wkYq2
TyRI/VPwrbdl5C5Pt/XYjv0UrH6kcP4Luzi8qkErDuwniIOvONhubQMXxp38ox9O
YZ2KPhzhI60GNnQzidEQSyIZR0aduzG2b5H+KYtw7aQrPhngV6RRg2H5Hbjffk1P
ChEWAvSjOvxv/01psW/nG5sYToM5QCA46xq6vP6F1x/pa1WHAga9NhUxUkQs7Wib
UoQc+zM7Mt0ktap7tp3hqOn3KSDrm6F4cG9+1dvP4xk40BaLTAQ9GOozz8QQlpwp
HxdvFnEHV+SMrWhn2q+q8m+Zwr1lecVZPJdgi+GA0GOv8o/i+TN7KBU6PFvgN3gv
Or5envuXJo8lxsfwEPyQM5G3gsmYtCBSTA0ipxhf3ZT7iOHWn0LwhGcL9qDxCWuc
8oVUawtyGGhyPDlil3AVaQC4V40WLsyVauc3rw7ip5NMgolXbQeQkmWS6sbhp/O5
5uFvW4dzIWQ+tn3myMIY0yGAl10/Bl/UNAUSxKu3EGqCkhuRJZ/LvlzpUvekUapr
9NPIwLLvgjgj7xmBdsAqddViFKq7sz6uHKI8RVygejjnVxnU9sPHKrxDv/kfmdrU
91Nhxk1NCEw+4ga6LDYOi4FVzvjbOeck8ZLrDBm+0q6zdcW7qHKv17JuZGS+Eocb
A6PzyE5wC25bisnLne4/MzaB5Iu/I80EDhWVU93W4yedqs+JMzkotZ2bi6X/lLdu
cHwwSnkZfQHEgTsJJhgdPPvYwVWZlSM7HVA0+XrcZbNMY+Mkp52P4KGouXOb1Eq+
MQXchgGynwfOlJ1PlFNbKwO4siTvhH43tDG/SkgEwg1ikdaNJOZ8O1Zi6YwtBHG/
8gC4YoSbe7O6T3PzyLH96AnYo/6cdXx0Z47K3IVSJXpG9w3D3LMN8ZD4afyN6V0L
FtUiEoQEE/++0VcvvquO/h40KBW+UjmUglhNNkVWYGda4ILr8KWTU+aY1mbzNIVc
IH3pex50D8QX+eC3S/g+UB4iSsHtSDTEvMw07B/Ku+4kBnGDik/apjBy3RnQGXyy
KaTLUVTpVHbwiMcYYW8LxrSd/EDQh0jrH4Lfhe77w/2dJnQwFzg9CBi1Dvc16w7Y
LQ5wocqAfjRXiNzqx3Crve0JZAEnD7YLhd9T/6UrevyeLxzRL1fQZozTaoZ+mGhl
X0YxWjmI3ZFGI7DGScd94qJ0zOdI5GLRg6p3pMwX2sieKLfTMqgQa/lt/WcknIp4
PWtmeoVrX9A4ADYwQxIn9OM1jAzyA5D3neNTc+PM5DKD5QxjOk5y2wbb9HwD6d0W
OCHn9qA1W/ekBVN2Ka+U2SxLl+zzuqRPXmUhVK7eHYVUu2lPcstzpstaTzaoJlm6
nZh+UOHX70uxVB4GowjBbMmiadP6L5XSmpW8u4Y95vNjVKtbKXv2uF1ekDUANbAz
1tO9SxZwa3W0W3zSwrn9DFwPlXLevTTw8VrFvnUBiywxfNMekwiE1N3LFNnif74k
atSfm17VjddZef3e2AHXnWRCALfuf43NyTMBK+kUHF9Egn5Q/z9FfMssrtxaNjnQ
M3np+VZIVevADRyJKf+6o0xLKKbEfhfFKA6eBdkiGQmcSF/H1/6TQrTXE1K3ygu7
XISuGiuYpidKtHg9sqb0d+yWuMd6JwxBXbyiYb/GsJUYnRuOOwVjomj9EpTrDONV
BtVtzygcAGdnATuvc7mOK0sO3kIfJ/viLoy7j7zXt1+KwneBacB7VHJmR0XyICTv
qddIyevj424+Stusm7owkiHLJGk4usun4MkNK+tTBhL0qq8pdHqHl0xrXVofH5OJ
SNBubhHktIBUytYW0+VlVRq9dbzLGlR5S7NxT5j0jQ1LhJejw/R5NxWbYbiSutjk
R3QUjaZa9VSR6TJ4ojOlBRKE79Vu8qppLxwlAYEUDHCxXy2FVhqJ/D/WiJp1pTyV
He1A/O7Hto1lZLv/qc9fXg1yT1Z7VpuWIj2C6+HeAEuTukitqEYjQpbKDsV/64am
UIr7nl9hr57EU1a1WhX8Nd+6vfz9BE4RKQI+C9q/2IEsSMUlIfIpsqp2zh1Wlyi/
XAd0Esy4WSACa3CSjD2kR0JATlj9jcEcIsHDB18nv23iz09uWaeI+f5NvAUrIQZK
T5/0uc/kIYyG9ukPNa3gD1/xPiXL+CsQpnfB6CxeaW/uNE4pQzU4fd1YinF01do/
Yv/yZEDT7Q2V1dv3e01CxZCqnwM52+1HTegDTLF7PKneL4sXpEqS02ZpX8r4t6fV
DScgGluAkgav7Oj03pJSKw4tCv5UMjlT+WpCEdgeAGfi2aYLNEEew3u6WcnWWgdp
GefOH0GP9q38AHLqcHSy8JYeIzCUVd+inlYfTw/0eQCSBDouRr/ytlG2jSbuPyFX
ILbU0+okPTwFAE0mONZtDGwPGnt/MFPGApGLYcXD+NhIQ4Q01chNFo1sWNSQPbhy
cw9uOlyTODJoQTU+mRWpt9JZ72k2TNVO7hJ+W6tMIxNBSqtxWsUkk3D3fCmI1ND9
pKt3gcAEU/TE+1aIxTos0poNafseN9AsPBBGGNvva1C6WhwL8JvsHBsHVi6lbY/i
AiBre+h1GjzLH8ZIdzIbYbxfYqdpqlIc3/+KLzhsCLG4r3G9buN2mdf3KeaynP8o
Du4fTL65ruClHu9cfXpmWMpCB1CqHUuDLGYSNVCIBa07+pUjydniynIiCQmVLlSd
aWPCXD4+eZQty7iPjJWPzpHh20DefochR3rhLfmqBZjzuZmDw4qwJi6QKqJ3Rbto
Kc+OI/JZr/JXYzxLBvaoVrtsgENmkif1KTIANB93TSt4fqXeDMn0QSq5wUGvdYE6
+eb+QJlVrchbP7kbZ3Xe34gyeCEYdbOhlsIdQKI8O4B6HtlYkxGMCNnJX0J+6qO0
c9Kz8afjcUbn2r21NJxb4e0QQ9urxB9ctmtjBq4wlhnZnMR221LwvW10nL9OXuw6
TpFGP7x/VKiZj6Tgt5Ni8I9m+LW5dU+vz+QDLKz3bMfu6iwDkEWMmuqdhvmenns7
1JpxrbQ+LJ0gYuMV7n/1xpEoDT/9vBriA1kkpuCzDAs1Apn5u7rfnIdYMWsA8Dv2
+BKyUVF3qt6L9/Oy2+howImjwEOeFGnpAaTyvtBxQItzm5FjALwH29MDq2m7Tfv/
5yJwtKyzJW7i6H9fA8uZjh9wCrkAxoug/g225hrtNkj7rJjlwx/Ghrj90RkHCiBJ
TI+UYk4XT/TourAhnqhXhalqK67vem8K/c4DoUE98GMVx0TXsGRQY2/H6RnDl/LS
L6BQivRfvvd0iRDpK/IMFKcyZm1pWruqfghsata3hevJZ8ZWvp29arWk1XQMWkXt
8tkCWXDxvXBODxoHHCEV/DD9ZUy0SbydG2pf75XflKB0SEn0biGF4jH52XIf6eV8
zp0Q1Nfe/wQmGV794GFmol/f1q0cWOhHJnRAW1+VaVC1mq01PZBVVg3yZObauiWp
hniCei2be2qHxeY0PB4WDB8YYiQbZCqDbHB9FRgt6Wni/Po9y7VsNQRiuB2tYUYb
VSYXBwYF/R0mg48r+NGGVmxR49n5Fobfb+EirWhH/JXx+rJ76bR/ntPpmb1XY8Ps
RbKMiQdpeFC044jacEFQgFVwEYIDvtzMn439mLdPqm0ZhqtbZ8dpm2xgB7r8fDZq
L6IOQG/3UKxMTH8mXyR9GGFJdxZ70XHLw19HiimpekSFgxQz1gK4Gkwer0z7otzR
n1U4ZAUWwTR8D8MbrLkCGE0LF3L6zcoi+95+eGKnCXwmgd3ngvTBL0RIdNFJ1V9b
snyKzBWVaifoaDJS48jTEJgD06MyZJ/O6idMYwp4Iy7YH9jrafEm10rZSGYsyjpD
dWEearW0NzFkMxHWKiu3XwF+HfDcrVglVX2zssI43/lkJoPoDdkUyKhVJ//YRFaw
Hj0G56QbKBoGVlv21jIlxKnt0jcJemm/dJ+W3svxMWHJQHy9ajLQ0OPeKZpI4zKo
dTBX3e3Bdz9XavjGeYhA8xvlm0Trf2f6mMFQTegmhR07CnSbRhzLeZTJBAMcpHz3
AZ0VzW4AZ1NtzwZLx4Zh2/GCxq+siD2RQkl8YvRyy+rcNRqElPaRVdo7edfmgwPk
q11QMIoaAxqjO8+oUKxxg+yXbwx/pEGuyBpJQ0kScNbJcpRcpwKqJcC8IGU7rBQ2
eandPzVSzV0x2/YcFMYr6vT+0V6wMisCKzV7TJZ4100YrUh4MBoeK+LLaBBnjwKZ
5MUCOffgwUjZ3fO40yMIjN6vgDdBMHFG9BG8S0sjLuXwnicNQTtGh/H7je8zIVru
l2b1b9oc440aCq60eaip8vmgfCzi2neGhvUwYEM2gxbjQvGqkgMKWsNk4ZrLUCEg
q1P5OfwtDElWGPPhAKEXtd57b7azS0VdH20GG/XKlJdekloIvvUhL/kmHaP0maQF
QEUvcbv7AAlbgJfdSRhJeO6JpAQ433FPTkOkGJPL1LSQzXhLNtyo2xyZMNu/NI+u
eXzt3b0Gk8Das6X3DXD2yiSGMOdwVHpxVWxN/luEDbIwSCyyEbkguy2jZtwXUfki
9w1Yo5XjYBvsW7JcyeHhrWWElgjiUw52tJv6CtscN22qb0PAyvChSz2kJ6EtpA1b
Qep8qYJzx0eIZbfkqSvvL3zndAuX7b3XtZ8FDT1XofyXGPgExvlDICZwLgPFhDdC
peuALRFjEP1g8PfjRDAugPxqR0GxFqxo7unhz/8n0s2p8rOfo5XOUKY5b/TMlFZj
mRQYM7EELxY4fV9vkVmJpLdzUvIEf1LsQpivtVXorIg4rax2gtQlAmb54bRjhKYB
8zrE75HyqpKLDZ2YG9gzmA7doZSroD+F/6D5rfdUso1CnKVXXlxp6iuVEJHjerXB
J4JmnhN5nTxWzHcVXge90TVhipwFPWKleNoPek16/jNZroVS407M2Bt5U4tlo7XE
oQaCCT1dPkd7zyTIBwTluolzXRSYuCAEUplwQb/DV9f/MtbtCz6auhSWPScg4BX7
LGLoQcQOYazRp/DCcqeWFXIZQ8+LARb4Le0Ra46XZq2GIyb7M9KGADDtEWq/3Agg
cNKWVJGRtw/sNLQvz+9tXlfZQa8Qr1TdulSb4ETAZ244eulbLNFBxk2P+4prXs8g
sOJFzoPuEl9BX32XgQLH2pbOifFUbkb1sKP2jqTf9VQNyi6LtaW+qZk5oTdzQdi8
r+5ynAzCef9RAiZHtyBtb4xfHluM11Sqo/hQM9C1XC7wDOT5A0Cd+g0fp/7HZIbe
lyCvpgDk7japd14FdS8tXDFt68TmwanINwMWwztw3Q45081zsWqiwAWGKwYVXRGe
xpE1L6UNIiZcj7WwaiOGW25wd+23l8OW9i7T5ABFze4EzqlWa7OBBthJ9zY/EE99
NZc8mjC0IsNu+qPE2FgKVDtFEGm3wise1JpXeOp1B0uG5k6vGQCUAUH96A11NE12
m5XMO3jUwsuG0eFPxzSnbK/7vtXDtdwzLH8aod/c9heAnLpyl9ydky8ukTbs8cCk
B2ps8B/iuGMg9JeivuYp3LLg2GVMc6JYUotQaSBzEHMsRvLhfREXI33WyB+eKl8Q
6QEx952B2xr0K8/ifqcUK41rFkSJepiRJHbvMjHRSJRqRC+pz7z/JwMdMakO7KuC
ZbuVmQYDCrpV6LkQBhvFtHGDww3tLv2s5l7duskOKPTDs0CczY1xhsidklpQfQ0b
reX6ZU9gFyrvQHQ+Irpyb9ABdLC1s/okdxWHU/XMhfkJ3nfhqa5K8xo27BCSxMMX
zwub056LQzvS+GMYbpF3YcbY1v3KECFTanuaKWFhEBHlLRgfnORbLFic4OjpUkUC
mY1Wqt1+dP8cqcuwdezuBQHCoe+xN6ar98WSH0W7Y33Vljfpo1AqNog2RPhcaK3N
IY51nSc+8WmCoJmrlbobSqZs/jL1Bpjgor9CaC7Zfs6jq8AJHM9BRJZPpDiGOsQ/
igddoRrSMmLez/+kv0I9CcBHTvzcUvHONjzt85iFDGzeBLfWPWzSdp9hYQF7VzlW
XtnB8mEvOnHqH51+Le9byuwkq7KvpSn0ClLtLpL2YakuD0IxL04QsJtUvrhERw5R
qN1VE2M02NV4f+L6pPj3imqOJjVsXO9PnrEvIMl2AGMU4D2De57eGu5PV/FQXOmj
j8JfSrQRDTr73dIt5B+AriMcALj5gd9i9agoVRPxFHhcd6indMhwI1H4troMrF1w
ZkYJ4YBGgtnlS86OYWI/wwHzmDJj8s5dTxux5xbuCw7KRuXB//uKTV0OgFp/XPiZ
JlSVBTUEtWWVOO9XAMauNA3VtE6GljofyohBMw3aAkuTCLXd3BfwHpJPYzBDpOT7
8LBroxm6YDeBvVAL0PYiFw97e2mivo1+l7WXqH5SE/J6A/dWGf7iX2xa0/OxoIT8
UDKq/XmSWg+XVkVr4LrEd5ncju7AzkkW0m1UARHf61lRQwi3dtABpCdE0AHOLQET
ZKHXLxEGlE15EUOtvu3DPHwGXF9tjn2WI+qq+knYDrMgO4N8xD0hXBWE1mdofh2k
cSsQTM4ZFDfZaBUQBrywdGnbHmHRYFVXRk+uay21yHCi8TyHUHYjnbuwuiftcF00
l/smkIyiZArzufPusiiBUBxwvBlLQGTDm8GCqg2khE/ISXEfem5g/D/j1uSvOPju
iQ4FdPXHE/bLHwrTplObyiHKqsRPCA9jwBFLz5vtfYsffsU5CxEFnZ5z2YH591Is
VDPcn9iNmlAdG6/OmwHenO2ux/MSCcR+ytvPVVKb1DqERfcGUqYUnH0jbUlYxJnm
Lwq7cSRrZIaRTUzYKkppOkWwaRc3wYdOEDPSayhuka76F1A5OHIURmlvAzluVKNb
hom2S8rGq0+HBq91Goh9LpF3gEAuL3/tBwBFN++6DO9OQD6zKpawWq3etAXSbXED
+9WoXTVr+foYslUlXp8hgJD4aMTnVWyvXJgyiG91g+y6Tz4T+0uPKR7tL17gS3Jv
c9xpiUcJD92CW2ay+XTvy9xlaOEcGQ/9OSzQgya+gy7s1QLbpkF2n4s8FepcAyex
ccpMc8WTCsblMD08gWOoyRqZxYBhPxVeKeYNQNVsKCqrDEaLaFq970X6QfLIHo4S
ji5eigCo0OJbfBjP5gN13UGR5qyVsY32BQjAr/UIqrg5XrCqyIovtU+8IQjTl7h1
jiz+Xr+wAw6zwIG4KRqBjnhuDiyIP+w8hzvJCMa//n3RVL0hVxrf86VujwwT74Uz
9imeudMXpfEtEahbEQrz8DXJy+CdNuGMd/jxsl9OL0RZuyd3lzkbZaHr1D47nfQ/
FV81GqdhRbWVO1uuwV3r1zS1VL4xCEBLo44Ha8oyD+Vg2vC0KVMbK2ahWOwArsex
hO0RdJRvmkKy404VnmLN45+uiUj/8FMLfXYKJjne8KlhwWhhWwh7rlnFYE9Ojqz2
4Q6RpN37MWaK4gMtBJKIHMknHVY/kIKlgsvzV98Qw1nXrpx0hks0PH7PyCAzd+A1
Q+Mc4VkowSf/IDZcBnHEbZEfKAyfS7xYzxrQnP4u2mO8Y/DbFCKuVTkuACO+8yWq
DivZT71u8LFoQqkPSCc97OK1UMf/FYPoNCcTkiazIqy2JSqodLNfVmlB8Z+GV/Rs
Nlf9Nia8tXqFY4LphdoyYVrUxIb0zOIh3RvNKAFwUgbnAiJEObrWX+fmxvAFfvsz
Ft1VVyGxAOTFc5gBdpKo88Gdfvk2AmajQGyvRXmLsKHwqz9RsF+51qsu039k2pwF
9brvW39uGjVNg8I5lQ/QYY+JM6fYpgZa0tCKSaxpYHfJeg9naLZqw1q8gl3Oryxx
TwgA5t3L2ytQboc6ZWaA3VJ7mKtMnZc/HMeiUOBS+/t+yusjV5juDarR9v7wqpCG
0fjoOa3n5V8qXEOjO7odTduB2biQESCzg7PGRLyArV48U837HxainHsV/xIaPM6e
8V1KaKYdiiTo2OHHpmOh5knQmIaWo33A3iB2VjCdrP62Il8bqwwp71KDp9xso65G
zVYYSyEhdmxfogQsbYOc9m8abrESxNA/J46Ejwc/Kozr8zt+4x8XZ/FxogCTcZAZ
F9JYENTsCBaG1+SXROC+Ocx/g8ZQnuWp3jfVhxE07PCD+iNrQXve7URTPb9dqXHm
a4nM4cwwOEahsVNBzZJkP7ouxoynz4p0rv6XPjPmHa0L4nWdhUREY7w/1RwxxK21
w4DJhgtAwsP92uIaCH3JokS/96ADj+CumXIaFNH0KW0ICS3lBteXmYtadQjTyNni
ORfPGuFVGM8kEMaqzacOKy952/mDrw8wWxEL9/yxGfGAlzHXLM+Q2J/eKt0FFIj/
OP+jjtu2M4RJCo21TWRxod3AWQN6QIm9RW5BeicQGBafEDFZ8z1ZMNb/KU9PQ6pg
LR+ZtllX17rhwxLROboS3LNbQpWhMXopYEtC1yoydJvQ/1H0r4vfb84QsfxfsKSh
qpy4ScgEXLpRbnnfFbLiBdRNroebOGl1jpbyJwuGyQXKm6Sadek0uJkEsdTxJOgg
024ZMWrzKP8LdMOQBLT+79yrPZSH18zB9Jzl5q5yQsZ4fCAEzWL3WMC9leC/ad+O
mllM4UfDmsZkEK4f8rI7LTukYZFqio8m6EuUEyWx8IJ4L4VZeXmqCCrPhUZ6uqAR
W62uiVVS25IFlU6Au6xX1ruZjNhClGPVZmHvHmEG0YrO4faA+o1wHXLDrS8uNV7B
ICDY4C6Cqu+r4C34jrDh7WuFn4QOMxCuRHwLoeLCDlebVtC83MyOey/OWm44xay6
HDE/Rwtm4xtPFhWCq1Utd4uJ6z2lyysZ8YIC5UNJ1ykmvuyZh3VlpLMxJ4Y8XgBP
0gjZH/UW0JxT7pU6tGYCeGX5NOPbpk1dvmseStky8HmkhAXpU+v2gr/anBcrKmy/
oeMisT27FG+uW8+aqrJVYiUOszKeOcR7oqh/9qZ9T8RBag3nknCw+vzaZB2kRAFS
eTRO154fA7/B/diNuT9QK+AWR3A8oiBTabJ9JjOUMDDtBF4411BKBasPkI5hYuyw
uKkQO/qmA+95ClQDetjsKad1DWXstfHhFtb9Rva2I6LuAm0N6D4Ayx1yxrMPb5aq
NP/7iSo79ojV2PX9PbzT+Enn2vE18AlGHpqoL2krl/+PGz6zrwZEEdSD7yrtuXXn
Nu1ac7APrK/oBIqzrHA9ALzrnsj9SIPXmcga8/DatE2Sedapabjf+9MnRsMECrlj
by1pb2Uoj4O5zAkznGdI+/3pxhe9n7o60p2pKPmpAT1jHbM40dW1zr7BnO0xtv9H
AkfwAL+f8msnLS9fm+QZSWMgC42DW0g+1zMFPX4f8iJ/But486xLQ8P0nc6tPt1R
2QiR4IFl8T34quS7btEtaAiTgJOQWeGV/0LeoK8q2py68fYM4m+xBITI/8UgRF+A
GaA1Rlhk0Nvy0C2xFYmNkwDow3+527U2F6jql5IDUW6sIaUsyu7oo8IyvjkLUCOp
ADkZr7yC8rHRvxXA5ESIPu5d0mocjsLooEi9laUQBOuxDAzXPeBFT6aebpAT/bo1
U83WXz4kMcXV8S5obAx04az+z+s+J4dUMYoIDM5A1N2Zjkej8rXhmKqDHpah7Klc
scaLLHnFclpwbhsm5fHx0HX09e8j0wOEU5hrLDfTuHvRYcOdk9kr9Y6jc5qqj3TQ
Ta++FsqgkDC4MG/cgWZG4hj9ub34TIdaRxsOdUN5YQxl4VozwBsSPuUq+LNROJys
doNQZLaZMXCHP+IjWD8jWE3OuNuMnigODp5pE2CJ53ULz0PiHhN9tNkIa+MY3HEo
XLQo//qCrGZ4/o1eQXDn12WoZ9iOVXBId757wbtjRZ9fwgOMdVNUIYNb7n2phQjA
QW6O0iMZdousAVvIbQUdKAgVqtZB4hBxoAURRr/SA0yky2pVuucfCgYyof5Uu55E
zOb8JhPlH2V5xXsZJtknzr+KtsLamSC8wkbJixUXKnK+naCQbUcRxLw8/gRBvc4j
4QfVQQEcZl2kJO/NlD6Mpgn1TAF95LLrDrJt6GAfpFoLc6/NH6JVHiD4mESbcdaj
owWBCrbbXCdymhr98GkAMe1j6LToIuhsrneIXUa/GwTgB72tncKSOHFdTTefwsde
iP1WJTCIIB0Sb7VkiKHTsF3dUPUEwMhjmmsSknVmyHOtJjLo+35OB2u6VewWKjNs
dDsBgiwjs+NlO5QOyZbllR5J5OTDla8Ml5C6jQJ3t1/Jkh+S4vVNARqXMhmWUxqD
zBeWr3qkyYbNtlv3GJdPHo/5z/fkyByhTwmLAq46Egsmt1sM7OKIkG21cd6E3R5+
I/EA2rCQn2C968QoICTLXrnJrC9tsU20lb5ortVc4i78tz/97+WJgm07KQmkT5C6
RXjP8CIeIvGO3EmkwWHAdG4zf7N53TVOvQU5aAZ+7ZITHo4Z7G7KZyBF5fQr4O+s
IvftgnA8V5DgIUcndCujZzl+51uR0KoQGhv8FNCURrqxfaKisMrZaNriT2pe88DA
0NiWfychvNkNAqk3XpxwjOa0nTg/Dk5sm1sETTn+AQ+HCToaPG0ieIsfoJhamatB
0hKYw2g7Zwlt1cp79cd6rkssuSTfSBIazL5eO9n/33YyaebE5YFZ+dA2h06k23Zh
Atwffj7AP3U1lty0N4OkYkMezUEVTUQ2J8ZVRhyILrwBi7S9ArP0Xso+V0T2J9Sq
fXS3h3iWhgsCAZHh4d8mGmHhsIoNsp92miukWJb/7/YJDBgAy6QbYgGIF3oFYyBl
ZCNSe0a1fV93qw5fg1mttcBe7h+dGCWl/HyNO3xKTf9Pcqa5EpRAFsHIKq3FpdMk
KM8ChliMUFkkDulv6zaslJyevaekp7CWnJLDnxE803C7yx+4UjaFockNd+78Ilth
r+lX9OkuiClAG1IwtXspO4Qw376IJ8DyfkVBCPw7daKB3HvLPDWbm/HnQANGi87/
wO4/QMnrwWTsz6Q9DXmyZB0+MxGS8abzeAK0bZlSC4le4QmwGG3ATMQaaIL7KLyQ
GCu3VZy+5282P7Lnhkwg2k3rFsx7KfC2YVAJ/rqmtaf/kNc+riRPSTtuTPB9qTan
bpZZ8E9fxaLRlKiT49/Uu/2jSRukpgDz6jXH1MqccWkeAxFUZ8FPstS0N5qQEuG/
CGO5iJC41FgfQ3cjpuNxLarTwKNGaqf/Btk2UVPrSR6pjYwWlIWuH3Ca66erjlyu
VleHRRB5BZo1jPHGguF+W3hSf1pAXzZ4S1JVR46N8A1l6mhWjpv2fiRoW0aeVwHr
St0orJ6wD/jtrm4kUmGa8LRnpVLyz1w27Oku1TG/GcA84aZkuyPaKPeh5qw0SgQS
BZbd2ADtNqSUCE97It6bdLOTrPlZmjHux9eSBOSDKuuqf+/b7+msXfT3LpMxaHHM
k/SPMFHdBcu7wpbg00wSG36d3FYp7mXo3Mbo6Tc4Jq0aMgyUMUGf/jowPHTU+rcS
tIIt3YeygCs2dPuou/z7zdYLwdAI3GC+/YBorPW5584smJF3CPXuVTwjPg7wTsBN
4tG+0ecez3DzCNZTqaIH/BNsaLINa4yMd84sTGtb2Erv0aM4AS3S2uIPCUlFH6+j
gSY03GzrIdrxtYjjvkh7o6cY8JY+G0B84echreFSkb9e5GUzt+KDRqPy+HPO9Qae
cpRfBZ/7s1ckiKoEVE3tLFL4I3agc8BBABpAxbWhBFo1WizGhOhTX2jd1g4j1G7T
bXEjgdK7wkxCOON4HiSsi65LL/r9Z4jLD5cLxJkfl3Uw02sEGiZTIks73dcd78NU
rPg6F3tbA4KWqg3aDVs9EWkAsPjyiVBtRVb7DBko+/2PsdYGLIGr2tbfo13inHEm
bt1dHyxKKQFfUd7x8ORf/wqfkJMdqTcV62feH+uS5qrOBz37CatdrlHUHLyg5QeN
MNWqHlrVDIZzph1r0w8uH8diDawgVB0ClfWUb9YwWInOddsW+LOX06TjmwmeFHCe
d7jbnfPKz5jCJUrnueyT2VDU0IMSGId129mPoDOWl+Dm5WqaweFo7XHc4rpLogAM
Z6cUZMeMP7dpByarpemlk35cHy8+wU3jjFxhULu0twI4u/STZCff4EZQ8zejgBqX
CTzs4FzYNBDSgY/0jJEf6TVKWkzJdOG5JlaS5h0neauSgUHyZhp+nPi8mgF81RiF
ei/31GuURvjciPOFs2ipFdNmEEvpsGA02GZnIuCHzlZpWonGdtmCVZUMrGevvT/S
o020PdARzmblGO9DoCn0phdzo7HjQriMfESK+gWsDIE3O+oUgH5L77/s8ljzY6Oq
wkRsCEJGRylkrhEJUwcIY3C0P9yrLpzrOu01Mnd7zuIpPSdiZTNVpIIgueqP2/MH
CjTNG59TCEpLXL/g50BfIK37Lt7lSd6GyMvERCNtlmI36/WFxq1gOj9pCVEsC9gA
o4xdp9mBhnMScQx0M5lX4nJeZaYG14gZ0Wh1v2F1WPOJOPV6taOOg4NVEnXZj2zd
8EYYomHBeAsAKJ/JrIIp4zspcdx71AX0Xk4onlJEEnXWOI9hDicvEc7WOhNSaKbw
IqaU/PTPjTKiFDZX7HbnsR2miCI0rp5AHbAoRy9m3XuC8QkQoR44rEfJQ/qwFOuS
g/GcNhGSrNUVGlYmtipI0WrDC2k7PAW8HT6BQ2+2CgoI3QLG/3yRIzv9UbZPrvln
UL5E+fakEsi12rdjfYdQzXCPRDfYweR6KJmwTC7ud2GGmM8Aj4/RIv/1fdbdZl2O
3uVNwKA4UJEjKQTPiTj/Rsz7kPBagrxwxVcuOPi9p3Rppjkho96tZ1lT3ryKcumH
gQk9OgZUdzI3OI5uD6GeoLtPE12pckaq3UmxM8IXVith7BotJdwgnYsnkAYip7zA
cjyUd8RtoYV6IzqDWHKf58FG+fTh9F5rAczbwaYDCgQKqTKpSI788MFPmWPjNJlh
Sly8Pt9QvK15sS4mgI63AZIq4oMLmQffPeYlVUvd5tjmAVL/B6cDnQpAL0aFmMVN
xMzbUsQig5TUIJuPgNXF50yeSO+/S3zF+lzfNUKBmezXiONclydN0MBU8hTwAcSg
sElMk+1sPgD+eYjhGjgTmljjvRxltlSFqjJ/oYM/kryw1lvf3Ahfcir6lFK2S545
bfnfL2ScujKW/WLaJFAy7ST7ZNdlu8Kz1h942xZy96HkoXU4t2s6AFAffPIfF3IY
hmbWMrH4TGk0D8KETVspOIl458FCDmD75QxI6xjPcd+O2nHz079hvyQxKimzmSuq
+KsGjYjrTuGT+H/wZpHUZlBSlXi+ENK6xtkv/O0ilwoUzJMpWRrLRtwyM/A1v8TB
4toECqyz5L92bJZwvzkpPz6D2SQFw/TqnUR8lD+761/ark4VDt4/9WED6Vqb4hmB
XC7yDN0lwZhw7MYskII9eF+bKdb2sICOiwhuhCVytjyQdPCPwJvhzE6iSxbYp3PP
/eQXu57sw3mZPj28+XaXBXt3bZudUWhL5H9xvDmU6chPH1v5yPwCm3l3y3xkfQH3
2ey3PVDQYoEXUZwLHp1q5A9WKWRyXnaveVX5FZv91MSWLa6bX3+cbb8GoAMnKkCo
hxBSTaBNThOSLoV6ojIZhW8tWUwMvBDXfqHNq++eaNJBFMBUbjOJeLYEo7JfhEO/
2DUmanfvTPc+r+fP2eZFUqTZMdA908tn4RztxU7AeTtzcy+3xX9HaOCxMypnJpm+
uKPEU8mwVAQ4E7CsEKSTE2og53c9l/EZPoPv1i3y9S5Lf6EvfEEYhAdp2q5rzlus
MEYs/eVWBi1Oo1ijPZhdD4n5RIx5rPnD1gz/P2y5YkZ6+Kl6JB5TNCIZBGJUE3kF
cbbFyzyGR1APyCkOsBQHM4RRc+RpSvBXYEjZXxJzIxjrs2kz9mofts6MjXhemx6n
cl81oZvsfS2LvStrZ8sa+D3CCsPs+GCqqG/8nYWiqJx5kQmPt7tzrCTSmjqVu5QV
wErs4y52EXmCn9vWe6r7hKzSXVeddh/zOiPQVIzuRJuddVKJJIF7icoXxdgmMo2b
dt33e+z3li+IpD/cz2ARlU88SGAFffJ2PoxdIRf3Rf3NzrHIhPE5gqt0WTmzBGqL
SdI66kmDgfF+AEYnnO4Q7GNR6T1D14DLrJluNMztmgo0L/FcXnoWn4RnAtoNU68p
b442ljBneMCcCGj10wN8mgJCVGZUvMI8AEiXmf7nrCfyMUwo3aXr20l45ONfddQ3
qPpaXNloFC27mORg2L/chxSLvluJCf3w0DgHd/QH1QtQ8tVSf2avZAgvgJqCngs2
wDzSqdsXWxfj375XXOFD7GuZ3XmYrFX20wrNhVJus5wzFYR7LB9qiS3/osvLKFJ3
nMLCwvy5dlf4ZL6HAVjItQmSIlOYfuGaNynAoqQQ9g03yeJoFqAlp0tHy9wNItQK
yWrSCvl5jxV/xBjTTXWa37Hco08kW9H6wZ+X0Onc0JXio8NMGbL1n0HO70W9TGqn
Ud2DDTqM506lqwzQcX4dY0JKoEpFgChzXRFOzZt8bV5cEXF2b+DId0lfIi7FXvEB
BZbBNEUcRZI2Fl7Ldv7ZDoeago2qtrm8oeA4dIiFK6OyozKJgseAKSKic7RcOvFw
m5lARisop/jlOHB5envxxPvv6wLG2ytcC2j5x3BanP00PY+DDJUTpCCTPuzOyJ7T
vm5s7GifgiWSYIN4sxXaWs/K+85VkHIT3WErX3izYPSKvyd1tbmxGqeYHceWUKFo
9PQMBU/hQ6FFQ7cnTb11YrNVJRs5Pxsxbf/Qj1l+FFgsOHZ+7fbJkKRZC/blo82V
dWg2DE3MEms5qatj5l0dBjvFVptncOld0MewtKASoyBL0gOuH4jMWfvYUeej+2AK
LhYA2fBEzmJ7b4RN7IHVsDcecwlcdpq3VNk6XgiZ46lw86AKaSZqRpL3tDORiMn6
+lCvNjH2ds/I6zToAf5rV9j07l+xr6vtIAC3rps2SjFBn6rFnyCKcvr1Tp1JvQ81
kj2TgkUTrtTuSHbvKu1o6X3moCO0REVkCJWC9QLirpxEfZ4WEOi1djUN9lKrcvmh
jKEhYf0/ODfpHJ+P783IAqFhe1uW3TSiYYCnDwhEkWNyFzDEtw03qMYD0JbIWp+d
XI38G6KqxZxPT4vXOwZZR9x3qU9rx/tnZqDJtALqfDN6YHVjVyxoTEK3Rd8wJrlN
cNTMNX5pZlnaz1EHlht/9nl6r+r/inuDUVHIz3lixMDQNC0NGXBVg9LU5wve0kpG
oR6A/T3hUy04PpKOkjGSRRo0H7XeCS7Ylpo3VfUPTOAexpZx+VCBS8nleSfGo92t
HjaO//ZQOBV7agcMDc1sm+abP2qhLsN2/5XO485o4yXtqmGhB9v1vgq+FZ0x2yyx
a8nTFbnHPmNygSJd5P6wNUiZsoWGXXnzebCTXU4loM6kRZAa1x7GzNUwF0qfzSso
RiCTbZVw+cpvvIy04bAebi7HTDz2dThOkiT5yqElEVu17b6E6aCUGwLkBLFZL1V6
qeWxQfCN1b3VRoy14sMqfWad1EpbI+HsKNf0NwrUTKPd+nbh7CVAGNUtBfsAntZM
nrwIXeXKg2U6E4tfGFPI01JofMwCP8tFEWSp6rGp9QrniqLL1D4mqFWUMFcFoy3A
qza9hqN4XDPLTzntFQOAP7spDRkbHOe6DjFsFLaqlvg5XxiN8dVFSKGdFzAXKch9
5r2XJUqh3DrHU+9xZ7vZkrpgubM9Zqg+CuTJziEHvgpE7pOQiSPOYpbNtXViARYI
JiomgZRqm802bi0oKm0BZQfIC9xwar8czmasEM+J8vBS8xWC8NA1Qrw+mxzrjbqP
uegfT6v3sRZzF7JDnCorf6RfMXsHu5z8PCUDy5EkfrPO5O8TnQt+7ODcovKhgfr/
XfQDfwvXYBT25C3sEnZiXZXm82pGIWHBfJ/tfeRGwcUu0BUyUaHxL25eLnvjQMg1
uENF4jZsczrHQroTJBIDYgnndC5SGY+Hz5kX1oLHWEWkXGeqTQX8jG4Z8IB3JvFp
0RY3uxMMzA22OBgv8MyV+dMIoN3mbd61remxwsOmBduSFCiqkkngvCuW4jWf688l
yweQyEnxhJWlgmISOcrIv3jLJSJ6x1CFxaxR1P1iXVnQBnRQ9AXad+J4orryoiFE
SuN6hmEa4rdyHB+kbdv8fQGotq4IZeTAIb9waNSWBjV8ciLoy54JUbQvKcURuZBL
biRncY7TPnvkPlIYZ6lEXGuwkGz/jpubvJwUGQ02G7cPtiJ5gvka5JJCrbcnFjLb
TNwIA64/JT33rEiLE8mDt0ZBWZIrv9y7R7HQn5/auYHi2mxFSw1XwjULzEs+AMTN
/+NfeSQ0rZURV3PC5W+xGuySRrCii/h/AyOVZJ7X8fWAwtSlkXy0jKPLE874LD++
41JDxXU0r+hQiWvQGZkrxlVhzMpR8qmJ1T7KSFT58gxIxipEbi4p2HQvz5dvHOXl
9SmRXeIPjpUwfxq9Ab/TZD65wwBE4jTUmVpZez7j2BtISxDoil09hKAGQg5dRk9k
zoGXiDOb6L3AlMEmfpz3OUty2KfZ7arI5tPBpIFTz9U/HsxLgs0nAPdlY9qZeN2C
wRHs1pzZaDuxSWMm8HYyhvdbxNz2+/i1d18rVbyp+aITPyLP76zW52gALBkoQcWs
F+UPySIqviGvoFisLzbImGrP/SAY23rVk94Hiap9/bzb+pcD8mhP9syYRFkDJNvi
aKdhj5W609y+y84EFlwqPmJZruUguLf8QhDqvSdnJTASzH6r48lEVJbSfAnaubYD
VVugGEjG/+lvAhThVO7Vjrsf+tv5LS5Dou6YIUDvVKE5+ngemhkE+KNoWkEibsT7
qppe0AkcoFYpQ1O4/Idofdqn4cj228lTlCLkTrqS5z1zhyKqxdYfA+WuKG1uRQxu
rEgzd4pg+pwobKNBSCAyh9HwnS9UWc8zqD16Tjq5jUv+gGqRa+eRKoK2iF9saAFD
rD8624yJ5csMB95eCvAkefbeBxcO9M2Iij53BrpPM8wmrWbm4hP8GC3vFU33KI3W
UFrw/5F/IoW7h7vhAXwbtqBT6tHoiYbFRBOUR0v71CPR1sF0yoxPNQ9Xp+FHmSlI
T8KrerV4JZyQajViY0eflcEULwSH5DBukjiPvO7ocFtu0+GHbuK+5b4msTcRyaqv
hMt4ftaQtKIcKhvZwO3mkuOIvCVTwCeCzm5lL04SC1HVLNZqH/0IQiZiPFUBeaTZ
SyQbCKiuxSmJLF0CRFZwZkShOnXoDjEsjRydPVZNE/N67MngwGhVCXx+iO0B/J6u
nnfUQzK4FSTr3FzXpuuNIYuqdb3/Nr34ZjQEz5XYfsc6wbeZOCTPdnoUVkTyhC/H
tZ0rCzolgOpDxBclZYBaZgA4O0TQb5Cm+82hVtgRAuqlaiR5cnZKmJc9FNSIgyYG
HBIVBrubjUBPPgc0t34qoKHPFb+wbM4pK53oMtY+R7NKYt2IPKVHZcGQHNhnCkfX
73k7mT4mRahd2M7D6o4MlexvZ4rFzB6pja3GFIbRdkSoVfS+xZGfDdUD3suKSvRZ
CMa9JN6cWeVTZppUM5Es1Zp8jja8o52hLF2CycWCJIUGbpcFbf8RNp8dHuOi53xw
pnxZ76FI2I+pmyno+XKIQxDwc9S8JTT0N5V1QVv3FqcgAU60PfuEpim6v5Fs8iyO
q2jZf6mtqw/X4zwYdVqYArGfru+GEmjhCm9YJ6JXXhq9bs9sbhz931TlrHDnCp/H
soEbqH/GGHAPQY3chQAXi59lhUhYEJ4e5ePXNq3C7R5SQ8R12h5d3nRQIj2vda/4
79FkfxBhYikSv2zOqcbB2jw7rOwxe6Tlt6IdpRcy6xNBrjvopSnMEEzrFKu1SGcW
vo2SyOdas5LJ1XskWg4lgN98Z3BtBgGdV6qChFjNuahkt5CvkKdTrFyAu8QT92Rv
iKjgTT4oG+EGeY7BHe/ZiYHjj74Blh0J05tKYDilFX8FbZSiSLKwYxMQC/Las8jB
9L9BjXUDUgiMj552SY8Tc2I1yA9HRKZueLSrdQFYuQLtzoDoglNTyHWOXzVSC+o8
RG2hvxhpIUw8nBrJKPKILb+53BoJ/rmDXGxKJm8Vx9JNw8mupksgToUbW9vlcFT7
gtrpwqDB4l1qX7XE4O37Uqh6w71rP4rvYyUsOEMV4bVCQxoSkFNG8dJvWFMgI4z3
j1EL2ad7N8ENlV0BTMluvGmQFvuDzcW4/ZPGoMpOQ54vyKoFCUsK4zIZAd0Igof5
/MZc2ms2glS2yuA1R3wMj5hNPk33rphM6WWU08uJmBr3ZPBio6q2DyuFoK4E9+VE
67elWCZyIXTHt5QVljHeVdqUc6t4a9r5VX2Wi7Pybc5mdR1OIllkOMeJTm/oMBCA
7Rjj+g1mp0B3I39FBkC8wVpC60aqrgqQMAk58QwI42CjVv1pqW4bHw45U4PIBkTM
iNUdCDiOghuZGbY8l1WbwtUd1tzfZHfm/LQ6IyU4kGq/jGVrjN4FOColXt+YRPKR
FG7bDIxO7sv/N9lfeTy6d/XTD7hUHFELg0FgpE0IRmjQZ5OFNRW9Yah7r3RjcBE5
/PE9l8Cp3izeixpd0I/RP0zQKcg1ZpiqOgN+Blciw7uIyvGJl/UrbVIrX8qNTaeM
rmnLB+zomdAP2kzIUDEgPG4nN+T04dh8q2ZEtGv9aAawW9QjAWcZtQEi1vKnzkOs
bfCWeIzJ3FB9m2DD5h0s864cfQZMP3Kvzb8xXGuWfc1zYhWoeOqdp9M8PE0kXSl4
V2nRJbM9kkrQ73V2bQzfW8z5hX3fpkZERQ4Uz0/pH5RkQTb5/cKyH3lOsJau515l
7MyyIolkeZpzhMQ59alXDJ8BMVzZH85H59zfM6zKu8gp4T2KR2uI/AXXIUhcsFl/
3FJbDiMi2I+RoO4O6Tf6ZfsCap5AL5YlmIEXSfueuI3Fp6+q+jTjHf4J/PJ/rkk7
3NqZ6VNeUgnZ1xmXIyJA6HoPysJdoXJe40W/ZOdRsTCGnB6BQJsIeJSevwj2rkk1
3Q9Le9J4fNvxeeLNXklse8HD/yZ50dadcsc6n64JrVU0HedrEEjmDSwggJmjI8bw
G9TP125FhQo4E6LoWofO1NNzdk2rVqXxEjiB6KI6rmDWkirHKKoJuklzleybpFjx
ckwmS7EeCU751hokMJ2Kzz7WDukMxszSKL8OZTAjZvR+WrUrOjTA6IDPIyTBABMJ
zxnHa7mROmC9sK2koa6sZ04xgPEZFCMqRGFo17TpMdNdlhaVVEjCcSuv8AyTGMtf
/hy5bsqmFOn9+q3URGASrL9M4771bs6pdjN2VI3JzjfSQzQ3PNtuA7OHOFMO9Cya
xRrELFSfRKG37k/W6PDKx6fJOyvwj3IVTQn5wc2mxjUvTyHMpytullF/kSDKBNL/
EsIdyeTJh1aSiS1v4yIAkdEvfDmAeV6Oj9qGNnn+p2JDVsvznd7RKvM5DkgsAZfR
zEg/3ApbdkGcP670x4zkx8ECcdVzqIuNiEJtGCEwDaxjDrlICUyD5ry9elPPhsoU
+rM+sgl7W/U0u4JixK6oLsfEgXiSaIREm9BO3nFpEk5WBPak2EgqDVUtijznQvmr
b03WV3l+HWT2mO0gzh2eZ7tDREexkKYHdmwFcTq2Sm3fCo02pktvUfzxSEozPDQi
uJl9B7E+K1ZMONqgBxdZNeSQgyuaNfCFmBd4p9GBX4Nva+D2UUyJB0Kahy4ycoWw
rWU/AXywgo2cYs55ZzTwb6ZaxSJy339cLbZ6kf4qOcy1m7EAmhLubyTMo0QX4XRi
GjkUhWwwgdr7Ot7+XqZ0IhJwuihkWIOQfVOCpLwZyNuz2yQxqXQ7ooCWiWbTVmcD
VXnw/8QvPK9rirKgJlIsml+MiXNxkSKKLcRMAyT4Pu4g9EhPQFAc83fA8U6F1ncW
Od9Ffq+7sTtYdpAqDM5ytKuvPh7TMIvvUi9znsapF6wccBzQUWbQXNAC6uH3LXyf
1w/9m3wvZwhgPeP2oej8Nw4icCKNaod4lExZnozKuXQ6QUdf83acB9IcR8mPUVa5
jrftuL0zuYT7XKexxH+ejXmtoKL64afWoYSpb3FVPad2/3YUB6Lf7AeYt6wAWfEt
Udj/1VqzMcgGJlBqf7Z1GA2MU5kD+NFHxeh1c+zwPNjdYykXlzlOVS2llPPS2Xpc
Gt4KS9bizMj5X9ww7zBUvZGwV8bGrtJKO6hLTw7TH7bDlRjEata53v1AwSxtovQQ
6vQ7WC0MM66zeBBbVZ9acbobpgrmVKrJkLR2+sHT25Jq2z74LZWRejvcL6N6HGA0
+d5TuuWVTDvDRZ2K6mvJIXIqklSWNqO/nT9da1xsC2qfFcbUsKNHfsFQrSrYhsh4
FbP9Uzrr6nvB0CA0qUFk6xjNvtB7vATBgmbfMhMiJmazPJDwIupZuC1r0gqJEe64
9lk0awdsnwlCdqWvw6tbI5M1C5VSbFQrr3EERYw5R0W5WxH4CRcxol+IZXDYtwVQ
31yQT1Eshet6xJE5ApSOXLo/3s95T983dAQux1Bc90sJIma4ZVbixTVpkMS8tfaU
PqqPRi92ZtOzmvc7u9G9A1NgC9mM9K2kjc3bwB5P11oH+6Zs+javJLZ9B6qSX2w/
Vjxxk9XB+YNMqbu4W9naBOhFaVuC5AXgpzMQY6svInjlrfoEMDOBJ8GILI/IolH/
Z58AiBF8gWuydt3shcon84EWDPwu1AKpnoBJCzRplhibga9N7Hoh43ELuDioWJpe
OiB2p/ApwcOckuxP71XBrVachhKHApIpy8kF1qaQwPliHV4rkmLAl1lIIhU/X58Q
Nr4kEd3YBLVwlZ7HYmc8ft+2BsJ6Jily/T/VuCHpwZQyj3wpBMHqRUnH8EJEKsf5
HfOSOo6jJh79TAlbFz2JrQF6jXYa6PaC0cLKIpS82Cj9fkfsmQD0iOVfUPxDDKKR
u88ouq4e8CMVnz6w2N/vfYx6a2f+Z2cUtjMAPaqgLVM44lzL5V0du7pCTMb7HOSc
Bm3gOKCMmqdwGmaV+IKNMCm2sG98a7H5p7tH25HPmBpUckscKCFdeVPTMrKlzTTX
bHlMv5Dk/Udf6m5iIfnpdA8KS3oPxOTNVyVEwy6CZNADei0alVW+jKtOVV8lzzgP
e0IObeGpZpqqBcsYgyIIhank/LBJewXnARVLrc5Hqa7C6uyn03DpyRPv6vMqp+dl
sJ4clss1BI6/X/uyQTxJOcAwGgzk51+lhKqfd/4GsM2UOJWclPk7j7hwinvEZss2
LW9fQey2f7Ly0/JzNDkFDsg6eRwRFPhVtTG8b13bDteBsyLesRUnweDbDRgnNlpq
gR3G6I4s3YhJ6dskZ2OQ11o9pM21teVrxmBqVGCpjLj1AhD29k0IXk0NKONvgPja
zX1m8EPKHkPj2gUxlfhETg2xwNJjWjjEg1aB3zpMhp+Dij7WlqKyFQVOL9dvOcqm
YnvRUYJyHF37uCo6OfGtMS+nKcM+SWeEbuOeIrnHZkTX+AEDKEpHT0ESAuRQebh7
pZt0Tc8SYRVjzP/zMQK27K1+gKiZ2Fi0ty1UH2GzixWhU/n2Xq6UJ+om3suRlWa2
2Vja27KaKq+xHRy+U9jVeiV/bBRJpSFiHzrRn9oXiWaU0T5iRZuiQ8DjIJJEhwlC
3DKxzLPF9WYNgAccAi/Bsb1YsnSHuno93v+d5WDs5V//NT/9dX7EuS1+sM5yAyCb
q4UTKc2WiUcxU/tyBRmGezQp3Cqa1hW6rlofAfGejgpsauTNDp6qtUs6zi5DQaKd
XjHEWs7slm9Y5fa8vuR40Tf4I1bxS0Vqjqt5OR8gUrwAI2lY4DC5ES3zzPMqqZxz
KR7qrV44r6fyIpOdZWmBbmYemqok0XxNu4407HITgWExhcfUI6Z6zHHfVkLwrp4A
jtcAjAcd/2bkCpnvkKNKrymapGEYxRsBcKYNc5Unzr+8+Z06fmNzEhVB3+HGmVUZ
M3wqEVmd3VH1H5fVFKRQY4ArnIh/WJJJWkb+/oxSLtKEkEZZbiWVMihKwV2PjkhH
mL6U5+PA4t4yE9+UCNsBzRjuMTTTtUX6jtkclj9D/j2wm1VoEZr5VkfKh7TdXmpA
XcjVsegARGw0pboS0Ei/WR2bvafSLWPpAqR5XoUFfVTUVnm1nOx4J794raqrXJKQ
AMOowWvxb+L3f5eD2hwFc6DA0uzZSdM6t8cUiE2OG2e5ngfRp3uVBQgfH22myMyx
CHneEDsNvon+wc5dcGLtZR/nLvzbpf77dd1kmugyiMxzP9wSo8wATO068WiXbApD
FBVeVVBaAqCscmdy/b+5twhy3ccJFe1W0Q2vq3Yf0ltblEm3dPJFjcJgB3Axy/LZ
TNC8iLHEHm4Ke+UMNZ5vSKKdIXKxlTVyFuqvxrbkqJAaJtrucpMwl7gAEL3Br2+A
6d1X4p3X62DEcjYaBTfsYkaGGxjUctj3YtOPMF0FzT7Iv3myu2QDYQOj/PDfCijg
4bCQymw4WnB8qF0079mH+9K2zm4TqIUivh/us7JO/BEIhzjfDwvUwELaPRb5T4xS
KTIAsRyWqzJvt+ZolQ+ltZWoZl/bUI1UM2mvLD7VG86XbrHzEmIa6x7oz10MaYl/
byfQTvOVJn+zD6D0xLRIdWjD2my9tRygdfEkG1pAKk493GIUdRgO4+A76x6JwIEN
6GTLD8czKc2TYlJiM/dEyVTJN866omiHiT3fEF5VuwPIoQ5ITDYYwbrz5PojbG9m
264L7Pq3MJ8o29Ac1cF3M+9BGsk2v6InsKrk1sofAqjszExm5aWrgVuJdvqS+nvT
fybx5vl9Ii+cKThNmlga2CMp36VAxk1KurqyuU4WDT/lWJw4dNg5oPlOHtuCZEAX
y/Gua6B+NMU0e241XeY8RIbm8joKGcqw2MiT1iRMMvoRLgYj1goZdhTUbvnSYwRi
YAM7r34dM/cGY+5p62WqjOdilWkG0fQCDc6UTjPSzw1OoHMy/BDJaHB4078tATK/
DEKtLbpMFgP05Sf0ybdn7qks2ocwL15/jWpUZdNR9p/mFcHeg9KPL3+8+aCt0jq5
uz6aF9iHGBdlvw1BH5YUa1st9055O07ByWiGJ6zLQDnsWefb2i+OMTn2cLTrpOgB
6ozZDFN0AZYLeWXBHBzkjtF68hTCUjr1ekdbgny0hESUAdwqTVfd8/X3CC35RqGd
azwa1WdNXyXy2LmRHsMIr9bJoY6HmfG+V0BR8NR7CYMxiIymSZjuwx/SdXgMNOGF
tZLr2vs7YhHyVyFZGgSjBa57TPCPZubSx/gc5QbIcfPU9VC3dRd+M+omNGiTmMqH
GaH8xppE6MzC4FUPgZM+Jz94LWg1dk3Fhl135siGfma6yeB9RuCJAPju+tjatNU3
i0YBvhdrAUqQZsjXyEVNeDNnaYlao3I/d1+sCBBYhYjy6aAXrVo0hPVtgT+O4Ykw
RIyKIIFQTo4W2SxwlZzHy/G60oEUVFINJMiK4L21FkkQqhGWgC59rYWU1KEGiSca
0YsYZelHEihNz93siqfbu5jllxwvmC22cs8sxJFPJ/mBtB8eRjdwZYFcGcLLsbGI
1AFgWI61ElaUMWkAua5ZX1IjylBYm0XG4Db20AXL3aDehgqdWmnljWMyW8qU2azA
BnRAroFo1EU0mDeMDOindpdAZJFSL395UXq9X7YswM69cMumx6tYAdqhJ1uSklU1
0EUvnG14SJ1fmPxtJH1dgSPupK6MO0A4MmZbnOIwWSu0f4gIbS9i2XqlMq2w8k+r
gSG/35ZsMJ8OsAN8RF18uiOYt8ZeYBmYaUsma/HNlWHbWNQk2ktsnzOub0ymLcyd
2JEM3tZ/asDD/QxfQxsYX7U6+WZa13LHVjsyKRhmyi0NgfNTBqhmjEOU7xrW68yy
MpssZV+HCpUTFZ2GBJJMrQdtYGz41PIeWy2rklwbGo/2tDkHtME+7bzKW2kREdUz
tyr8X8f6jmy9CAaoFxGKn7D3neSZBF8xG9PQXm7uqEpt+b+p+WSzti5LZS8Y8azA
hlydQJ8Td8ssY0uPqxpJo6UVQbxuky2WTAOxS6hPIhI9lHGbTTvq7m/LzsMp1S2T
AD6j1YyaqCZj81yWwOcxKxbeodfd1t8GzQQN+eXnP77Z+I0U4WbaJYrbT+y3tEEQ
eoZzgiDRUb9Sqmu6gUS/VcQacaYjARu979CdTJhsbQWrnDSYGklIjSSlmQv7MiXd
2+YPSG0DLdevAj+KUAqRwmReVhy1gJju+HFpMhCIqLVQZ3+5M6IJzrfmVkZ1Ip9b
m5rwboCAnh0fa+e0IGT5ico5kXcRAsYKgZCGL9ay2ZrL9j75WyReA5ejRrDpBr1v
ljJRomrZcTgFlgMoViMryr0nt4LQxiNGIM6KIq3AYLgzRNK39RQzvSMcEeiM2d0Z
KrsLb1v7+kSkw0zdzX6chdsujyBJ3I6V/ZGYt6mFTn6wkO2vcaIlEE5J7JcSLP+n
s9vj9URmCemKSje2oFGcV1BMkGrq4GNod+ruQfK2ieoWq8oXuyf3IFCvm3nKw8UB
cuI06cejODCx5hcH1LP942WapAlMqc27U0iqYF3Codq69r82vEl8UytFymkWYfgi
cPssHc5jmoe9Bw/ujHmsOKgaTSjK6UWLbt+GK9YxoYU7dYdxSD7i3cFjWORRGDg7
0gB+A2PZ+1jxKUvhtUfkL4QCzLqvNkuo0qIW6+3LoTpSWWmcStv8i2MVaZ5YqlQH
nB7NlRasMFnno9BHrH4NGhlNtlv1j+TuYSjGcRI75BOpBO5LjG2yYd4POaGOUKOZ
TgrDU4eIcWhOtUG6eH3MzV2yMcfu8S/HQQMwqZD0SuS4RrCK013zT6NE42/N8V8/
5TAJjnB/2KVIzSZq5Nvr6Om6364/HmIGD2vLqmE9ZZHxt7wLAgIjMmfJqAaX1Zpn
lnEVmB3gYq5Jh+QgHamfKBjqnfKhpN4jm4mYqn4mGi2ZanQ8DGg5WhVES9IPCgnx
Lc1A+a5hUHNhFQXipAUfBxxegXCk4PRoG7Xt7oLSteoXWfeJ75ohAhJarY407ca+
1DvV9c0CCkJZXTMmffnP27oyZE4TXqpiopNHMfJ//5CGG9A8Y/x2343NsvHLUNig
ds2ecpJqcdEIirOxz5+8pUCOj6/SEJ/Bu57fZkwzK+mRQ2oI8bfzX4vrfPAfDTk8
IlGJCp6Xh9NiqJctWmT/i9UFF1/TGko34D7O/WVSeCyZKq8O1gwlCevv9S5h2woo
9tduekhiO+6bQC5IALMY54XPRpBzKvjreXQmWgBAxWAvuqLxdq7nWqwQ/FqvcEpC
/5pMuB45F0e0VyCBv5ctbTiw9z5oh7cNcahs98+JL1SIdgw1cLIThfOZToSFj8zE
49TVNSWD1GY4M0cxjs+35uFcyMn2NLHDWYhldbTo0Ug79U2rvvG4E2Tx01bYPdXM
oFXARPOfn7//FarM9YAzTfYKtVPhZLAgDUN7MJHa8vSMYu3Hjuh3ns4EY/30hUqo
9UR1qktcN7YfIAuddg8lUz5NYtcD8ptKffDB+I4jlAxy+9oWkbvBxqdVAhcnRcca
JbMNyZmXnnxNq/9hvaEvM+otRcyc0JsUm2Kv3wto9BkA7SGuldB9NYQwlfG06yun
/v6HGC7uZM+yQ+53tuIIoZth2oKEtY7ekxMMXfQ0tcpNyLcsKtYRYlrHE8ZIU6QG
wnI+A5PvsvCH7LvGTNi1Yzak+ChLnsOMTxhX85ibMJW35Jnn8EXDNNqc5Dg9vdrm
ohJV4J3gRaYIgg5Sc4uB47xKsEgc0ycukwWswu/JfC+7Tu/g5Txrhoqj+7bbPGWw
Z8kZmsHzsxAA5vozVfwun4ANhz0sDmZktWVGXgrWfeWV794r7lB0MBf4/o2Rc6Ea
4v/XmZTKTKsjkHq04SZSnTW2fHp/vO7TRnsNIz1Y60JdC7N+Jc7e4op+wV4ciUY8
x4/71G3fxoCVHEirQJs97PzBZz0eIELjFltNQvpP+F61pi4OTrVKOpiv/9AGI/lN
xABiCgGaB8JHksHt9L1duMZ0HNOf47PUtWa5KAYDtnA85HMbP7MgGZLR0vnKF3e1
LJzLk8JcbYGwHjqME2WkVwDBPlxnMLYoAieRsI4qyuSGczE0QPeVs7skkv1ZCgDf
smzACILHUYx1nXEjEv4OqFoDxMVUBnN08ky4vEbhevPHqKawe7O6SKn2qWgyUay3
V3/wuQhPOjAxqHI3p+EwcK5EFzRWc2hqy6ox0K4IKASnKaRYYpcivDkcfvtLO8j7
vgn48F0ayRU+fRyJd+4tgSXDMsVjAM30GtifLIYZj2BJ+jRPHvE2uPdrYcqES4Gf
C2LbLnNlhn7WBEDzOy5LDwDolLiBGC+VveEGmbg3IoVhvrzr8WzzPORor3YgOeYy
AUmyjYvKO3sR3p9Fd8gDqpDR4IOxzvlXuzuLetFF3jNdXytlODagpzWeWrcwmLOa
k9kZGY87fH/F0c+0p0mxFZeuVVUQ9igDqnDlxTLdIL2YHHtttyklSWKfWw8PPxg7
kYnFhz0CnmFSz59nq/C6g5VYttJxdaus+I+43FVo9lxUXcAjkHQJ6+YIoIB1bV0W
73T7vLXzmL/ZZ24Jcqm+uJ/8m3rPejhSvU8tD5lI6j7+CD2DPKiuvkDe9jwaL7gQ
WyGiFVBlgPqurtBS1lj/rWFBphOOTQhKvsf06idqKBPIBxea66SO5J7TUJcdKFLb
1jqPpjRwmHISdoFeinB3MYwhJJRHf7ORk+u+iLM4d9lZxPHhM1DvLynfmBsq0Pbu
U4blEa3gqpxZLfer+9oma5/MhiNMe/bHqsn8L00GjEOy+H4K8ZaGXujjXIU6yYju
T0UavwEg7cSgrJL72+2QjS92PXYcAz5bQbG4yryZp+CxJpcudti92uHNpZrkhEW6
AfAUG5JoBBILKcy/KnlN2RPvU9JkZLbHgnbYrsJfe7D1U248Bj/FpWCnmvP5u/Lb
U3dFKO4CkLUNSE8HG/PhtlXK9s57Rh9gu7PEs2jJcXqxhqh8TXzyD3rbmFRnnsd3
gUv9SnOoYYoeiux4tOhMpPs1PLJdUxGNypitPtC1yZiPoAzuILXMKAm0jbPbsF21
aGNsVlVopGG6ktIlw9BZ6EuBu63lrJLvTswGheaJdmH3eM6S+4t9nWsgN33a+tF5
JAB7yAPNdHAZu2GJjvmSNs41TkBLocTWr98w9AtBfMmgh4g/363cCshDE6NdwDvJ
7ovPB6+3UtV6nhgjSw9zVu3EgI+mCOomCeI+zTxXhjUagQCAiW9M0JLuE4611Ktk
lpfGY/C9biJA5skxKpKvyrHew+OV03UUaH1FJ5lCYveqoHbOU7dqqBvIhYQivOWD
jMjcPk0Q4GhDaKQW7j0pK78tSroEAPJ34MMfTa66qJrERvbbG6xMOEYFQqo5udsU
+9VT34inanfVvAB4DKI456NZrIqaU6raO475n170aalSSSFOajGfl83CNla9gvh7
goI2HNUsCu0QUCervX8wlc6Mp1yWn9Zw9LUjaQ2ugrA8wvmxBkwWJJVWOpiY9kGg
sl6ypDjPv8EeKu1uDpCmHKcKKS/4YXWtQJudU6SfcYjar2+XginZgbOpwnwhoTTQ
cXKfES/ukV1Yjtx279mPwaA8wsO/w91IU+hYTyHCr3S8rzS/cOqnnYwh/HF/wn5h
xnfmAyfdeWExhLcl48rqwpdzDaWfNWXEdKnBJxDGffgT+2TVDikbGVULcN18Mvwr
JwXPfrRj1RieqrsCR/zupjlpjw5CKYWzr25HmQlgebm4UD2mr0M/DOjgT2/9Pe6o
+/71GxPr0RwUMvnw6RTduoqYbK1nj3w70zxAmyDGoeHAddmC75oh/Hg/GCW9PXKt
GETTRqv+x+DNgcmnixVY9cTdKya5Y+ws/O3IVsYepSICBm0lGpvZOyWdPsrBPkm5
01WWyo1akJ6PsFl7DwCUlr6EXrx1M2MxMF+/+ciJnztOWKADwTP7HNlOxGte0vr3
uwCpfAHOUurmb2PPzYQWs1STXTXz6rTzut8ps5/Qt8f8uSvHUQVRG5ZjHaZXertZ
W/jB4RRpnMXWRof/6Mc30+8hJ6VRSJmgk4nVKla3GcGW8CnrbA8cfS4Paj8+knsu
6Tvdpqw1dGQRZ831xwuAscnPKSsvaNujftZbd4imuxVE85t1/cnggK+IKVhEc1M9
leJ6jlD/Wg3Tr5RCNZvgm6NYdlbI4nDn+c6Z275kcnbjnvBYDH0+FCAWCTDERfha
7IzdX75ppjAWfVUisEXzUBo2BXXWaK7fiCt+QSySj5SKcHnsTXPYeDg1yZd8zPYz
EQvWCZhNgwQAh97gVLTIxnGtmgmNQq7kOwmAdjREn6o5ZOKwqWjSRqzd0LYxWG0A
RR2DBSuQ3qpnIU2/BWBAyyamnPVnDT8uRp/nrnldCgIe+RV69/3sqeVZ1biFVR9m
e6axk24AIjw9vcQoTAaCk8lTPl32dciCm5ElZuebd2u5MXrfCCDZD6PU3uBi/2IC
bbRiw9LoMdRgGGkd1QQYodkVz/V9z327f7bJLF1EjnNdB9QjGAicZ7JrgGDXWuOY
RW3TZCxrtD8P2E8zZih9D+kXRG8FwGsaOPKHrf2V9m6gjX9d1yqhW+POQfRIbckm
dtWa3YTbkbhKYlguMV77aEtn0ye7MtaUBLRRtcYv9nVUdUM0NUK5XHlB704dSVzD
atvuxXm4ieM0dVE8VW0L/z6R7R4dEC+kwSnNMOxgYTGNeO+hEvZBfUWQKIwtts1L
XXbu1g2xkduqziAjIZ7gkSBnQZ4zi6kamWujD4vkeRrt6unrZtgXYwAO1A8SnLB1
vaI0HPXmM/xRMVG/SWyHMrwDoViHomOBCkO1qE0h2h54X9Oh2SVYI7ERjXUAn8zA
aobb3WnYZqtvGoA5vI8i01e1P3baMZfSA92xYh/q911tUIRL4UPKYn852bgchXP4
GADm1WgHcjkyz/tPjvCnjmbCJpHEWPQKObXEGTxOWPjmjZnYaAs5RY31eJr8PBaO
q9O2y92dV63QdyYT14T+v1XBSAnTO0Op3u26hBhRXkdWBUponpyuCnFImMb3EGNq
Ep9acLlgkzmDlQ2cgJEZIT2El3lTfMqUN+l1XIKd2RBky5+djegRyafUmA8r+K2O
KjcI8NUbnIWZ8LgBet0d+OQLqyWhxaBVuwv9w/PPvGm2cGm+uopSDoKU32LnapC2
Wt8P/3RQGUTkvf0GrJze3VZ13zsrVfeggkxN9WgRB/eISEcCI/jfvy7njnDW+3WF
t93EerXS9Ubv99ZeS6wpcgPrfGeYeBriYKB4L7JGEYwcblaVRTr9KCe+50QY8EMW
XjiLFz94SkF+/cyrMs6bj4E5UaMqNZU7CbjMNbBPwKBig4pYF792+yK/rsZFAt0e
5OBtAX+LQNqOfvGO95ljjCuzahKaWYKGJ1dUVkGhLK1ZDmR1nmNyDNETIC7yF7fz
pNb71nvYJEYZCKgE3wvTcW8zoNUZtnXrw22F7D5+BLcjkxwgT/W2s6iHa2O27o/U
Nfzw/yZtMWRpvG62BvtEK6Manbirohgx9f/HElSDdh+zR/klSGjH74NsSpiUhot/
dCQ16Ez0RIwN+kV9at6zFvFlRWUCykl6NV8kC/GEy0fX+im+CWMONYO8q2n27MKV
IwlDUz1/+bKtvChk1Bg+/vxuNIsUCMsXPGny+qeAr7ReWC3Gnl2uGzOrc5dRNl/C
+IpyMxQPgd0UbWKZPBV+wb5NRrFBKM5RzUE+6+9+irI/U98i33q14MMKctjonKFO
IjeTKW+kFMgYMgc81BEtcs4cO7Ro/dp11qP/XgiYfxMvjuGuAnj8C1ZH43TdDscq
lVgF8Gc1HaPYxXJX1o+3Xigvq0uKD2cnjTOLy2/aj9wJHMJ1kOhXYw/j56VPwQ5M
ds2Maa6vYAtCbEVdaGtyc0g0NUuyQyJcEOVXfHpB2LDOxoMzcN4ec/WmJIBry4sH
nZBICq6ml8TMv5JeaUQWwkOzI4wBIMLZbLTROiO9fur9rMEKWzzRsskPiTYXvCkS
EU1L0uTlss0asAma5A4SswTzktRLVTcapE8FfmIW9ZDV4HfsoEV1xvJEC86TeckJ
VNqg5JKkmV0jetSASEqzPFJHLVfpdc4qdXD07EpbOCkd/RjCBnMX69GlihGpI6r+
HOHKVFA7+Mf+MRTX9+aZKbm2A7ddtsG0CAFFBuwII/2+p6tB/F6ja+Dal5eLn3tb
dl8EjBrKumFQzEISUCtXHgLDgVgVHsAmPJlmiogBb9o+qZVOJW6I0VlyOxjiA4V9
PG60Nowefjg+voTpNCc0YlN3vvF59xxxNRg48LAwifk4tOdOCBKKTsgCGHt3/sju
3JnOzzhonECI+yQiRdtBvzyodajyNEOkEJfa1CYqv0K6dx71RtumTJAMNcd5Bx+q
3ppUFI/Z7gX57lRiuYlS4B6qddd4YkCz+9EgjgAHp4s57bEFpi88EnvDuOUrdFY1
Px9txLjIIzd1isvqRRYzCYQ1DWsIGU+0YuuRNu2OUEAVw9go6nLne6wayzueuTOg
hdXnctbxKIbvODz80578wEO9AjH+5MYbuf8pqSNV+y5W09AAp0cHzrnveOosaSJZ
zvnL2JC1NLXH02uw+ZIDH68MspnYVD6sS45wNwh3canmtCZ0QXX/ZZWEHlCv7pEr
xq7fOB95alcQN0TPySZecTS0r0YQrXALamrWjxNWZDrQCInQUK2ucM+nmgEv/cN0
9RO4vsz7jZPuhfLTukDWaynXLzwtuRktfm9SUz/EswD0D2yCmYquZglfjvtd2c9w
IBoue0bMQit6QDwEbfriBLS79ZDuVWkVLx33wEZA0jUx1W/W7ZY/kLBI/xXDRmS1
V86vxgVE25ak6wARZp2RanDZpD1obkRt/Ps7IqGd/amsk9Ij0U3NOBOyiZ7fPw4g
gkE+N01Z4SHLpKu5FG10kHzlgc84KsDBMJshDi7RFi0erg+Vw1wCCQNTnuu+EexV
lQHWVtximTuFPNT2gIrriwceKxdlpM8Bbycj0guvCXNg/ereuEuE9GsV2SDPPPz8
yzer4rHGdTcq2G1vtQ6JPu/TgCIX69/l5P0fLQ84v5Xzb9p0am5ldUbeiKH7ld3U
s+R0q65YOykt2R/YILcQezo77gWB58BETJ6m3Xypjn8dgYRyLG1ccHlHRqTOcByF
cdyR/Ya3SHkZKoMcFzI/vFZd3s+7PALAm27iAORSp59msiDC1xL0a3qjHLT7uJQp
DKEzXTbKWHTj9G35inZIURGOg5f1Vur/1zZMiLGpKuPwNzE63HKgP1zxpKZtJiaJ
+smaUl5s90wF8LD96bMEVkXODTXUNKpHmrMuKql0tP07rw3i6GgerOkEdTR3NU4Y
wxWNjlvlwUITzkhEj1n7CoKXrN5Z47nsv5LQ/C00Ie6vEC+QgzbXg99mq+XTU8PR
1A1ZWkLbdubhMr+P2910JLFrn6VHEEFVoxd1fGtDQ/evw3YfSeHoFBSmN+A4+qQ9
bqS67BWNZ5IxSXUSnoahUqwv8WdNMkux4dQ4nkwhxloNmJlCTNh+yrfeiBSkcy26
s1LlMxb/umQkwn+kyHrSI2b/JMA25r9KTvjvR1GpnVF+Fpieh8Ex7M0a9NoWZRFT
N2a7Jv8LTrY/lE3hj8RuKgCX4XMmyfh6VbLi7o87rK/SOr92OgJ6FEF55v9fMC4r
QVIBQfRtuuc1gndWw8yv63cXnTys/lbbR/nNB+xOVD2gTyQc1Ya//4CDlSsD7F9w
VmCkzzVqRnLBkASCdWJu1iYWmJ0Zq+FVpLLnEjFFBZYaMDcZmOe/uCdcL4wq6h3U
t2D8KIDG9HDxpQG/Uv8wlf5CtK/9C61WnATU2jg/Vt2BXLLG0wfMCH1CwmfaAr/j
a/YnYJapmwHwqQNtuVM8f9EIj+MiRL8/xBFvYZiafKmy/00xQS0Cc9Zf63VDmdr0
WSknpShNdy8UkYemeHL2Xp1cWJEE131koyvM4qDcWJ3e+IRTdpLFWMpUOZ1i9JVa
5MqY4LjHpwZnlM1WIc/SUo/2Xgah8e6IKU2Bn8I8oJDSE2fzKJHzv6oFgiQ/yQoK
OHqNRLS46lwqvAoiaBvTmv1TiyGnUdqukvzEZ6lswPu1BsVQTrf5uoG1dGwIid4L
Ml4KSmMS78v3wEGHwoRoH7E0j1WvLo7sgHOO+1Ibgysdl1o7pn22yqVoO//EGxGM
fTzmLQWcJXSV8UnN7oWMGytazp5vDU8/YequcK+kTJqLrr8N6XDMk5iIDCx5XI4t
XgT7iNniSN2CKRhDHCGnl8JpIDa1M5NBoS5cFi3hptZzTiRUEFTR1kGihurmUdAT
9ZLobrcTI/ZZbWIp4rY2rDeapAX5KIOOLkVOHuCMInHKQZI8nNieoV/ezEoVATPN
vKic1oPql3SCMSSe6cq2J/CwDv+iHhKyrhZnPfJUGuSf91yOdQf+mo7Iy84C9gBy
sgNHlK8DG1PZVE774ngJC0Ve0lmvUH8vweTXxXBD51YzXsgtsUc8TjPze4W5yap5
8DUCDw59Fz4NI8BI/1gLmNtRWfEcw472SPaK4dTPO+8yVpLXkpzFBlbRl6Yu7Zrx
G2WfrCGIpyPmzvI+QntNknHmx18AVXSqNqOSrQoam2y2FsJs6Ncxxx7Q9VPOyIZb
x6p72NHH+LYMEUWRrfmC7jG6l3s52Kb0jjK0+Ogr7H2cQY1RrUadvhz4fkXUbRJA
wrQOa53Bt/RH1E7GEokxDWuqXP9wxSmiBpWSpoZWgCLo/EkRwjFgeP4JgqIP7R56
d3zxolcHpOPRU87PA15wyyITjsjjOKDDbPwc0bYle62N7d6m/9KoUcYTNe9RveW7
DMi4ySrdZCcaqE9jtK4Okp0WGvadvR/YAg0x+pZYgQ2yAUtJm7WdDahohYtl0rNL
jrSAloA7YZtE35g04Q0POTVNqzLkGg9unvFL7a4FRBc0j8bui03oSUtgN9s+Mt5h
C8TmJ32ngKwbT7Le4iLaIYXMkpyDNGx/PZ4D/1RtfUK7yKg2+xIOGOPGqXKUbeZb
lf+uryIchtKMYX+mFLfkBYDWl1wDSigBGg1PnzZIRwqpXp2+RDxRQcYYv8VuRke1
qjQsSJKYIOB6XGbF83A8hGH6URsLHRuuPQjXJlvRcqdFRUrKq3mbn6Wl/cgqb2gL
6oKrAKrfevEUgPLxS3QmqfAvKGr3QbaVyN4CCPQzQtao0Cs8Y/tL+sNZ2gaJmeAp
V7kBJFofg0zGwGklA4/QoXxzgzg+xJQEO2keMPJ5f7Z8k0aZtdzSb83XTFSRbclv
TxecYmCuMepJYHqDU9v9wUOS6+/I+afXQsHEgXzr7OeRfCMTS+R9plBreR41M31H
I5eQ1AKFp1YCgS8/mh5+1rB2bldQ2wH5lejDShqxpzpF9/XJow7qomn8j/sQ94ZG
el8u87b8F5f+z3E+5hoDyeEJPxwg2mX407LHNmJwCy5twa8ZVHLc9/NeuVV7Xurn
bABiuAStO/NOrEovR0nq6HMJIemwEz37VW6NdiMfKxjIXByJcpS3DODCAcefoeSz
qXSPfPHHnZO12ZAUBw1kqJLyYT1u+Yg5N6bL0eAQovS4EEfrAk+RNl9gyClAnsUf
jmZ/yyxqou17A3izVr+RKCMI94DUXeyYSPMDKHgfG28xQaNIZ/j4VtX0dFH9SqG9
OxOsdR9Q3eFlSFRAtEMryCB2nVR342WyHkTH+9RukG49gzOpljFkjMr0X32YDNmV
Sf4KeOnXwqPC18N+dE/4/ziQL3gvJGFBCrfRsYOT7yBOGdvTPw7Cej6RUzOBZ8cn
NXeukgHaCw5Ai0bO/NXTWWZMxsRiupTzBYG+XMZkJQgcR195mHXaVFwEcxY4F3RE
zDC4F1h5ryZANhi06D4wEz3UCT62dh4nDvKqvGQ9CFWIUPwmrrPWRaDbrR23Z6Q5
9UUyIcFjcULTUMEz/VDcUgplv98vp4xpW67YWrPOpbxqIknkIDgyaiEx7gPhETbE
XyB+B6ORL9IxnajpQrTSTNbWoCANaWTdIeqcifZQsgon+v6OTg71SMdZUCGl9NLA
hUy7p67LP0pDSDq85GBXpyeRTX9EvlY3WNYLkKmV816EdVtnrzS1zmBySVmp9vO4
Ca8j/WWAdK+XV2Gm71Tnh/byBfxOaYjehKV3ugQ6xroTjz4TGyVJ1Ant5z649TcZ
/Cya9NaXAdnFd27VqPIRlkim+TWffKrya6+iZ58Av7hvrnZ248W3uyFPWmvSDnLW
RZO2WKZSAqEvuapu+gEsrx1X+zJeK3cR5d20wYD52pMWFWFcW9vs1EQaK3IuYaZJ
83+Mkk5/4dX3Yh0Y1CX+1hyviwG9HT8iGqYLh5DGiu+A148iTyjCO8kcTQrAKtoF
NMbIUYVGhA8wdF4VAhg0ZECfTyFok0bFOQ5j88TkjKamOQIcHupD6+SqvrScC1nJ
6SahdoiQS3h5ocDYevLkcm+giOe2ui2DNMcKcfZnktm710xjabKoSkqjXzm1K78b
ld6pUVPklo3TqfFdOnuMRm8lj8wXQmd06XdpULhJ2urwT/yKJPCgGCjDZeGFVr1b
84fMNaHFcz4AWI3iky42aGZRlFCyqsG/UaDxs2Zx+kBael3SWC4g16/pVtFyJuGr
f9sdM8XbF93DPI0ypiMQzgzRRlbWGCHFXn5mWygRW4AZfZ6fKEkOiRO8ZKkZyPZV
i6Uu0cWHiiVVAAJJHEFVK7ToS4DHxjm94u7Bmb+T8CcYoNYwtu8rhGCoDdI57KFK
sd1T5pyHfGvjg00etVStqHe4gnzYTaVp+EVI+soZtVUOgEq/c0WCvtTjSE/h/+zF
NiCJH4LhCdCxRtaf3vUhxXPiXL1Aqaar6HaJwFONxZrhycIffqTZWvT4NEMQzSKg
Ns6NBrHyrx3RIH9lI70jub4KieBDhfQ5uODtGAuQt6zTHtJFx5qfrC30fDHfznUE
kaxNTr6llHJiU++a+YMrrsa2xtCXrKRAlta1alKoQ4yuy8jlVuFs7QMcbzioO57p
yyBjb6gQ32uY1W8lZCbrmfUEQIuFruLxPFMfHie8oaVi7muh8uH5ZRZlUvgeP7H0
g6OHYElEseDFqH/yr21z7ZfCDWI2y9SPT8bAObBiYHfzwHVh9QFzFwIg31/DLAhA
s/tuhXtjxyTMtBCCbIpNGNCpn8rv6s4SG8zkpZeafIcK2zUGZXxoM77QQbuQjnCm
D4Tr/DqoMOJVtI66ym0SFstkO8vesHDmY4UOsdt9oR1rhsaNipYl6VfZv+8ThWyI
CmCDC5HQaxBEqJ+87qgGr0oooUV7gRP17xnGTifpyaWn+ND7yPB6qEeob5li43HC
DcjiKWdLMyWmXmJdt5jpvrFKlkiPBE55IXBZTDY3TgM71J9bGO5QzXEXPSFM//SK
CPDEunMxMKXbMe2zj7d/EFK6LDbyh+6tQM3ssCRAzR4KVos36/PsEJ00uTazYzkx
d5BB9VtRod/Nwg8Znk0qGPGup0gNS3DG6++Cs+ofM6LMDB2rN/RQdKobVLY0E+P6
Hhfnl9gVMHD5hakvm2HyjVj5sxV2jwpjQb6W9Uc+l9CutseBO+U8uUF27yK3vkZP
K6mdsasvK096/8Kf1u3/QioYazfIWNfPlQSOAWHKkfCkqrDcSWFFKqXB2brOXkWM
R9znFsVAuO1mkytdw5Eo2ImxTENUIXhj+w9+VUv2bxWSPpHlZnDyyHBDTB3j8cB8
FujERJvSwlgdi/esBA15xfreHfn7PX5Ziod22jmrsGazPGSjwQHiKkpV1x7uVGqf
pf+nFYPUoCxq5bKrx9uJPPFiogXcRjZLBypD/Vpz8L91gko7IuewyeEFm6H7LB0K
5f5OBQMowKUG6KSWXQXvi/ODYdltWAFd2CxVrKLdV/eBJqJEIk1YhoohTvbROMUI
sQn2dy9oC79msRBpmEFbQgRUf4MKJIR28n26xIKaQxOGKxWWeBYkQzTzI53WxQZo
eeBHVtwwr8iGU2yIERYMr0Io/K8fTdWLmrqLVYWMmPiCIaBcM883GHdRMtM0zHDh
LUkf1V8wroigiq6klZLQAHVssp5sliwlvrPA+7oN63NPyx1gJS37MLoMobt5nPje
MrhlVcpRp4CM2WQWwGfn8iqBgbv529lJTfgwWdTR4AYNr4O2NbGe33eY3v7UkBF8
0Ueoyz57yrhhD0V6s0M7Lu6DBO0Wsnbw9RLFwVVonJiFdbtmPot0mBLkNXfnLFPa
pfPb4uZss4suFfoT8Zy1hI4Ljj7o1o2RcDlHPxRJwvbX6viVgphG+68BN2SSGw5i
yL3JxzrpUiAWk9BODq7lgXvUqvwadfmQjxJU0fieu8HpWFNKL61Yjo2J3/PAzYLD
H1+fKsrRf6AzcdFZBQ+A8x7bLMdiqYMdlFXdIgTB6P7qfyNo6WlHT51Pk0k+ZGQP
dIs8NVd9CUwZPhwo6tav7wC93K2WOl5kZKSXgjI5MoiSV02zfxVS8zzZJqkB0zUq
OtQnT6iSU4r1Nwvu2XeSVC7Ugbq5LH6tV5nQ9n94bd6wEms77FTbx6RdxoFNWgLd
jC3BR9LCUSKKwyWV8zlh7QIGV9BZcN7myOaD56zHQ0oe4ctacDvgkg0Rbr2iYlmt
edV1dwX19WH4fk+olXlOC1V/qUYmCkIQcDK9e++AofF/zi7nNchu414Ryg2IeQYE
Yw2/irCLEKmQvdGCe64nn1bDEqp9FH/J+CgEhE3qofo/Ndd8JrAEGPsMulXI2NPO
GLj7D/hfGvjtOndfxC2RRra0wWsxs8RGle+SjRjqljSpDIlsjIspJO9KT8lxapyT
wIA7BKAt1kztTdBjHAp5RxxyF0gHlHFRPAZKpah4bl8W5j8Ehyg+X/EJkDsJyDHc
NH5deNXAUlapyYpZ3rHlmmjtD1z0C8ixJ78mMxnnSMRGVUqQ+0+zNf8y+AhjmsON
LvrP5qpC/iF+EL3N4VhvpspeRY/o5E55s8sbaI5E0eKoeViKFZfWxSg6JMVk6xei
PQx+2x30+/8T/A8dzqBBmbj1Jp4m5UoB1IRIq9deVwzZ14IQr+OLlvi/8pZKoBkZ
l2ZIdzvHl6cp1ehvOr7LqqV2REe5AVKEiIdbWb47Pl/0MK5SChLBkvO4k83nlCjW
GRT80dXOUnzysSs30t9IpC/UgohOrVWAoDSWX5vFUfIOpPvE9U9pZofQZan+aX1y
uf3wA1hu/uVUeq9VLJb1cAqNlqjMHSA82S2IsbqJut9GLxiYeItZIK8rsruVjG7l
YBmPwXIwiVU1PXyD943y55YDIaA/8ugjR5CPwY/O6xwEoAbTbWkz4Nk9STsQfKih
PASuaJUsSEhVnmHVpTXM4+dNev7VxabOqJmVumNipRa87O+w/68gjdreUVIlY7f2
dcELt+cbFJrYLMtt7PuBleJ1rXomFCuA0CyXz4xRKVZeA2Fjtkke3mgnAJj+acfT
WaQayXAsUkRBs2myakX/AFbdTWfP1URkzLV+WOxDypTtKrZBneOAsmW7NWOl1sQd
JNb+8KKTptRP9KSdIV/G7elrn5Icb6BLXeu8VG/PKlZJ3eS2LQvrsy06Rk/iKXR0
tCwUKd5gomhdtDyGqIWQoF5GvKIZHarZUzZKzSR3D/OefvjAs2ifTw5JRHqJPBxr
d1mdV8FqsUIUzYN4AMMAHibNuOKgtLfFStEuytj23CbBrxSFuYgkoiyuFSeergQC
NMsXdI6aiAwmtGhhHVWPE6spthdWByhtFS/SLN9MmU/aoWtlpE61N/TWFBuJ6dOP
zINjgWv1dI8b6Jh+VAxS0fONTm8APqwYC5wBPKV462owg0geSofbJUHySVDEA501
sYylFaLtUJ//xugmj0FxavW2RYF244olTTwTXsnuNDG6yUuLFhFHTHYagNfjDjgL
UOA26e8iwWRKe8bR40laSVRZc8qafFiQjUdoL+XPPpD+tSkLJJt+nxFxLQ92Z7o4
+HJmMPL+l5VLSEzx3UIjd3UBs+VtJnMUu6iXvoVNz/E2G9F2o6t+tnOd7ZCHMahE
cpNHLlDaAVgeRPGnvnXH/RF//s2mASwTvXifI7UnHpOpQZ3rG7dbcSUNFBd8d7xj
r+pvY2zSD5U1FaDbTeoxnSYLZGfTaRECjvjRAm69BPFDDCaOQiRpGK4JywL+GfbX
YOGjWwZfH1xJpJ1EOKLDQkWazplkVshVskXLi7Qu32STFSBGUSiNHBsqbtXSs+n+
mHu+kLruPTVO1xQQrT4gsfjld7SOg9icXcfMEoApiQzu5crQ0zeNpMPrI4H7IEUy
1dqtfNr+qtAbCgC+zWr7MBPkYZ1U2Q/JvICycgTClI1QB1Os0KkfdgfSYInOnP6J
GNxVJFrNokXhyCBWHM4wmg0PGLxWQvcsux5YPcRrHsRLXecrmBp53zuU8ISHEBiY
kKLMIbaX2PFvUAa/aWHRDDm8u64AC4GaNQYzbhl0RxWxybwMH0Cnt7/+PnEuV49I
mMgr7RCh4bs+f6BzDIFLv4E+msEv+LpcP1GjWO0E4215ROR0mW1aHATK4L3bT5wD
9IPPvK1rN7y4cLK9/fh/botcAO30uGuBK0h279vBI0ApTc227dIK3BwM3rtyGpyR
yxZ0Di3WwICWHZm7tzF5PNcXnbp/1mk1174bZTUCsy4ElvrP9aMXeWiu0SRD1JnO
Hx0Sbi7vmAKDXLo6sYJFI8EelGdM6PSlzYxmAVsbFeUr6re2pfIsduc9tYVOZW3g
Afn5qiNZ8i6P/b9w+V+jqgxU6sN8TeU5cJRWH8rV8/eO520198Bl5tzlQBU9rSZT
0eE6rVz88i5uxT2TGRLWtaYUSZtVurzSd3su2/z6Dc57YY/nMAQZidHeIgG9CXNs
ulKsVZFRy/9b9esYfyCX+Acr+h/WERAk5+YjzHcpOSx2M2O84g7YezpERZc5SLhL
Geg/9MI5x7YySveJGTD4t3lIsVVr59pr65cVIAeRaWYQLzLGYuosEibLiP9JlCfl
0H3lulJxdXE29bx3i16mxaDDPmBgl3+5qccuP2y0CnwUbxf2Kk2KalhCmHeeJ0nk
6fvhmJ+Y86Yd9xcxYPCz6yBT/2UmtDim2opBcTbec5iZnd7q+ISlo8U6Z7GQ31MM
QwfycxTzSQc96Zhr2Tqe7zSfApf4D09o5QhywKtQk86iVdKH6pdmB4RMpa2yciOz
UR+LlHqdS6q0nNnHYKmCgBPNgSqCFMECYXcE5DFKBA/JieShySTAmN8ZhLyd+buS
MxmBF2QInc75N6W8ulyBGapB2aONbKErF5+jfVJIS51u14klRF2eOOfY4iR/2PJJ
J7pMApD4Dg1EaSI3EaEZct6UJLWpBBoMGkHUgQSSephlhn3Qkk3r4DEduOHWGhcy
iB+RNoAJ9IyVSTeQWhRzMLwAoTRQzwn4y1I3ac+dC0ZNq55/5lSBewMJRWYlgmAD
9pn9zHHOhIHTF7F1KCdtdWC2tHUBPKjdKGALRljO5N35+ZLfx+y66YyuqbKB4Apo
YaxdMOF+gKF0CGfhMCNkj9LBmGZgvvXJGKb+RRHzzfMiP6r59vhBz9LDYqfN9v3A
x9Sf3uv+6CDHhHmp7z1x1wLTdlPRjqopdpvw10L4wPt/+FEe1Hs1ZCbpxiEMUM2X
KY6CuJlZYAnnR8wltHc5PJE7q1VXbLXcXkUxOL6KOmKXA8PnhWbGSHYqZ3JZF1yU
zwtds1MFkluo6nvxRcgoNXPwV29+wIoLNvE6wL7G+fcvjNVC95KSY+VbE9qWi5kb
ofT6PtlreCV0ng1UUotyDYO+x75DSQwhCe4VwUgRan+UaFRANugt6g2whC/2Iura
GI8nU4ioYEqSUOzYc1y3TOQg+S2MSAGhcaqlmEgXcdy3Kmv36bwsWvdahBoMTBae
q0jlsKrdnNWsDa3PRoWzMqgxM4eyCMIywPAV7sFdqA+0phuKjwrR7NAkPdIWhdKx
O9x7HJncaloj005+o8QK1/SlgA9073Cf9qG7bI5Ws3iVfYup9mTNz8hlp/JRjJHA
mRzRnIBAz5u2XZ18nEAdT7/2uwkLuxiu8dmLa18ixJZhidEE88cjSEip4lYu5ELC
xWXE76gjd3lTLDDS/MerwpLzglUQRtecjaWY1YQJkUiDYZzrRMZ6keAlgOznDCs2
K8+BZGhcTJ2rDO8SphP7BC4a6DYUTpSmqjt4AZAluOLUmJWc/2bg+vhxykgRA/g7
YZVTPDKVEWk6S/V/mEDmvJrNTBNcpdVLbt+442SLjZj6AiV8UO2rvhbEkHlORTb/
4+89+60iY7fJRzgomz9g2bVDZQ79rl0J92B0NLCxfKAgxpGYRKpR3DKzsDdJSgXY
hKPd1JeqjltjFPY48eIZ0p88lZrcAtiHikalhgl0GZgMnCi6Rab49Eay51YAti7r
Nbz9OTCaL39e9bIsh9xZFRx46lvPdhsW0KNOhL7TvBgNrt3c9wxjw4AP8Vs4+1ju
IkZ8bll3EPldOyVoYUwQKaDBorVnAi7BtdG80bvAXWUmwS3U51HtGluaaRcw/VJ7
I89t/DIdCyAZjmqBROoqIum1SHghBs5Dg43RACZk5UNIanEXx2uOINbM693ixBpo
1HVNswxK2KxNj/SEaS/mrCl70o7AATpVGdGxjvWpwFWxULuk7jTvoz3SIT3JHMyM
txd/T7kskDPt2WrhI3eE5FAeeV76TIwSDsI3WutOYmdyJGnkbNfZgSEtdTVcTuZn
AqKbraBVnm9Hw6E25eMNaqRGt+/zZMvu8IaPv6DDdAqRhyyc+j0yySCzFj6utvOt
ive7+c6pSXeUjnwm6yvJcALL2Z56w7CX6wdisCwZy1k5GjwksT39frV/zAEkwHl5
ghuhszZlZ4g6df/WDs1WpCsfkzmBxZTv5G7PitJCkdnpYvMlHkA+OzjDTh9wJVcq
9xR38GJXcbIYCknUHNIukkSVyCuzrwUh4HTJZQ2NU/NvGU0z7lp1Wh5sz+ntCRpL
w39Pfdei2SHkxZQS09/QTvr5VMvLNimTmNYU0BrhWNfKXQjTZqh/crbSjxT5Lx3G
zi5S9918IJ1slIVcVYBZAG63/iOn+o47uf5M2kW8Mpao6z8uH6bjvsbmQSM5FIhn
qgIK8wXM4l1cK859GNGtVSlKfrjd23mBmJsUbWTugyAzr3a+6qJzUdj3STrWT/nv
OtrFoHuryvFqgSzjtcKgCgJYPMu3u4uVHvsr/5KiABanYltZtBfyFa+JrTs7UON2
FW3MdznDds+XKu6akqfC3eJMS/Sft8O6HsIiwqXFBK1EjsvOVQvJkU7cJ7Fr0Kx7
0HwDM0TJlNuSGMVLZ0hzHt0VCxcT2vxVBwknX5blmbkiCsdCP84MI8HPuYhjmzEZ
w4alY82LlyMqsnz8NcwNbz7GgBYql0+mdoRDG6mw3e0j6p88/7iwYoyp5X+UuDH2
0s4+Qe7oO0KUBABPqHOmjnT6RS3VdHMhWyyEMderMKAJk4aB/zbdDwlHho+kxqyQ
u+hF3W1IlFXgpJE6e3AHGu5cAVueEAHjh75B1dP3UhDcY/cG72e2Q2T8X4f6XqNx
/OQTTJlg+46RyH4zqg1SgOgTQA1D5mGZC5csjJiTd216/NQ/mUx3YW8XbF6tPoNk
MR1G/ZJIRGvQpA4XMfE/nvoVrczghmZi+KkRQhSIy6DpLmM138ytD8yyCHAaYXgU
X7n+b+S/hiNbwkDDWd1xj2fEaSn0TIwParVH8QTjdx30hMS0+Gb0Waj54PlhffZg
Mk43RMGnAkfbK9gOu9ubEetqlUTRz88Ob5hfW/XAanvkvzyXoiyMkSYxtZV7GDEQ
BSgtBsSYpQ7YZp32ITA7eykcrUE1L8azG3R40wztA2QoHtRK8fSJLeEPckqhaS29
5ekXxREv2KJaQweXDYNIaSswtwlV4Yhx9wlM5nLeVq7qjEMVhbIjeLoWvMNbwos5
5QR9ouIhBEVV0TBaDlYDJnDCEmJ92BY4twzMw5Tem+3LfpBgpEJxUwmG/o2XcW0t
33NQM+ibGJEB2VM0YSMvfSSulJTw9E5SlpDceLPssabdStVnRLzlPErVARJtNHl0
s1Za105GiUodAaUNrEqd97WVWmRAS2GBqH6j45e9f5CmQOtI0vc44cXg1GKKsX2L
d7qlTzhJESD5ZPdFOXArhsJ3Rdd4pgqnDzi7+F7zz6vReUPXgGZ6oQa0tixmZ5tv
JZ7l9mLx0/nL+5eVyhmvNH72xnNCi5eK4Rt1HrF4zL8RsvNVnADmazJQelhx6QPt
k9aXkRv9QuZ9WRyrDePoXlX47wmJ6CIR+mCXrHyYvLYDNogYk8XtK2U8z6mohqvU
tZ3y5h2flrqXfPotZuVKkxr8QWgyJZfTHOXk57nVWlRydzpY+uvGm1G3z1EIec+M
QONmv6Pj5uwcl6OnaCj5IkTWeXPSBh3/JKv9oRg9m6lCXYWzfAupR9n6VR565CRY
YZjp8KCQT5hj3o5qjXXZUV/XkCTKI620qjLBjoksrET7SCC2Ov65Vj2WI/0EZZOU
QGsGiYbhiSyclR2fWPY+gfD2qzET1GgM+paFsDr9cBZ2SkC9q4WAksXYF7cmbWJm
Zy/77LF9veJUWsoPiTzRntOHc5t0O4z/Q4tMZvRnc/GZB7MxFmcDfUYekbnNldll
lDE7oxiB/cQZb2egg2eCfS7fsKn0AH6unAd5MOAYPPGuOZUEdyCh3RAGQID/cH1w
8OFrefEFzdJZdBjqHWHMSjGkrU6VJJMB0HKzs3FSLtKq5TlHss+xNgPWE9LkrzZx
M0XA4IDqFjMZu7C3VmfoU2DNC/Cr4ru1EB6x5LgkG6+6mPw6+tkAv8MbhnjZnsXg
WiOTtTICY+gqpz6oMLWd2ZutxnOW8ngmX4yvuqvlQPDGEN+10O8ekkgCL3zkaoGf
jkpi64Q1E9IBgE8opWeGK280E0kwpmz7MZR6CUqOVSgzgRU1pTJFZHoSFiklsggJ
tCjT5WBTa+5Lxfg1r0kmi9yClDXOwRMCspoZzNoSq3mF/Zli2qNDa7b/CusPyc6Z
AFtPumSap5kvxmU3kZPm6Obk3PxeUA6o72WlHoKPyIEhojf5XKR/KBg/n43zyqok
ARdZJOb8Ldx8io+9A2xdarpUKZqTQRjuirJIWENXmm+j9dcorNimx9AC8Drba2Di
j66aoVsEB+Q19gmTirL01lKeqk5nZHQ5LiHbNFfE/XgT5rXqynGhKr8TfBbZDMWb
MEK50ya4j1iBdJATsceWT/TvNqyCwygGXS1myWPkHA0OGk0EzgGF9kAUmwji1HMV
Kb9cPABB9bFLte01PGEH8jiSurYCWquF7QQZTvBZztW4mEYeRfgRWacoI0rQm/Hx
suPddmOi+9QCpMw69ueW7c6YcPNkH/QZoz0g3jzGDbRILx0gdOuRMQD377SwSwVh
dajRMOSh0X2BNXhUvdmLqorqUrhUsYz8XNxF3TEO3vmEUPcCPSSZreiWxQmMbCDc
onRaUQ3JIz5cv71+L+LbKbAoakSJa8+0ngxX0M3iKkzN3Kk5CJUHt7ZbBqaof3Bf
O4WB2qD9UPt43AhZmDmEYSj1NQoySAwnlyZsVjiOucPIGTpvVIkhMllWbmA8QBqx
7nD950R1nZGqrxdaI9kMDVjtKxgdAndkNoD5M9JvHqXfWxyvHDwbNrHL9C4Nv6eg
m4QU8OS/pY578gsD+Y1fmqqrtejR9IeN9dHNCKnSI3R3rTqzZyIvbtuOmogRpnfr
WOJlmT1gdQMR6vcLit8/RjtpWI0Sinc3LvwXIHdt00Xdh0iQCpctvq1pX3ZMcVT+
wZY1ksBhOdr46Ekvuy0tG1EfDUK/npGDMX/d796bxQt6zgjJA7mVfIWJ+o2KTcOe
A3GzRUSbsQ6cBAj8C0dXDsHtf/WR9KefcZX3ByvAvyaoZAsNF4K/Jcc9VvEE2mdu
UjIJpu4kOxd6tT/n36C4RY7O6uM1Yx4KHso63dgwuSXMH6SUUa4iqBEE/ooktrWY
zip9A9TAJhsG6SlOw1hGawR/nKR1kxMfVUSEc9ZG6M7ITKx5fMhM+CzSHp1IvD8R
WIFWPNE8oH1vFPHMjEPWWo1ahYBB7j4uorme/a47RXxVQ+sqy3G5wMvT78ovi5hj
WpyMc7DBZVKOIH06XLIjSgg5a8lYWEk6J9oJXaRdXOThD7CfJKj3DgQEFL1yx+7c
2mCTbLnzTT0S/7ySCYndKPuH2t+YimpmxHJZDxR0aRR1pYb9d9OHWRLdHRnPX+AM
k5GDbk+6H4h8Zw+uybqgV28/8FYpC5QfsydKcl0IHpR7hW0+zXbSrHdFnASOR9NX
hJSKVrlvNXMzy9cq9EZ2VpGi8pXlRK8bAGD1OYLvqOlrdlXn/aQs5xp4EXiyRFZE
ryo/ZaKGdtODLYqmf73KVmykUDpQYwvAv0uXkqevrivxBTsw/etfX20ml1tib+QP
EehcCxRPHPqnnVfn5t9xeCoL/1sBg/aVnHLgGcCasSaYZ8pRpISyKH2dib1JBIcS
ZKL3K6afzDN6/wR8vtmiYjQaO0MAyzqB19BJfeiUysMtPozkG6E1mBYjXBNIzKfU
rJREH5sY8mWmMciRKlDuAJfyW3/rtZxFy2daXTFQSS0tKCZ45+rRveh6/FxDdiyR
3NcqAdzWYKrogGMvIUOr7RqIS7P0/iiA12dO9Wsn93A4nP2ud/4/+bBhpbijFNOd
r1piv1HzcSXpKxhwHtvhEq+iUXl/vwpcTHfRznzAa8/warJeHpUXLSoDOJ6lax6W
WdOiGb7qRx0Jck2mMTIS3BWkAAQYG2evDkWfZrfWOIl4gJqa2NiS12Wpy3+7ecyC
/73DGfBG4v2YqdeYEBUX82iktwJYOlLVbQwB5qBxm6hjgbAmopCVDDwkm0ZRmJ2S
nOHGfT+0jAxcAy1Gps/0MuehIDyK9PAiN1H/b2EKauZiFnygVvGEHESPz2oduDQK
wsAitgkJ1wtSUUHMdL3AzLVfmKrTeUiux+BsyrGCVovFrYfaepWpMRMVFKq1DeJG
ASscctOuYNdhwUlTrExXyRP8meMrPux6ZOIs3569gMQt/oVO/Jw5biuF1Qept2ps
qFqNN8UZDYtcO9LXMKZpnSMqqSfByWMO95aTcDu1bP4xGokrTF6+0sqLaMV+GEeI
ri4CTf/LGb85TAe6PKm/un7uU6oeuqIrZP967dro4dcKqCkNlvNQooPrx3jmUNp8
bII3f0utk2WsiKOwin1MWr21lzKCc9EcdDYKKD03BjbYcUtzbpPrLplq/Wafi4Rz
kzJ3yVp4a103r+MICOD0wUNnmZI1PeSzc36TMOeF8V4+qIxqoNeL6U20THmkTJ0K
z26EBsdrJuo5GgsIXIhkU4Jj2uZOQRBVVcZSmgzsUko8m3htDkKdkwtUjB9HncbC
cpazR1ZmgTsz4mXc49SToCyl7jZCkJZPgW+facUu/JIpMQJEyyAbZJxy0Dw1HMyb
kCRzfvfp0TBjMCjDBbgL/6/UCxuHx0O9C9WuaVfq+5eI2tItQgHHm/nZyY83HvK7
yL657dzJEnxYdzCzi9ugFHroNvKvss1tZzJbQPcw6fz6H0B2dcreZvdUu3FpWLjy
x3P+8l1wTzkHvkCrpMdOs2nIqOGkS8vzUnJcrwS//D6IrXsXvWFkuPRv54PK1zXl
dsn7NqIgebclWUqSHCXCKcJGiwRn80+htWJXxVq/T9pJSJ8AGfbCRVWRNkIcyM6N
IC0/Z9Rulf4I+1PF8fC4uSEaCMCGIo5CFeuQyvU7u0jKYD1y0Cs5xo3UpTKlEZxq
s016uH58XSxoSP04Z6AHy/sYHaihV7vK7xA8hO1zoCsuJLP0ttbczXRxpoKYtOs/
/aHpgPiecf9bFGL9mT3NsMj7bd66tioJZeObwN2ZMrXWHC3tYLbtUwdwPbxJdt9W
fn09ZVoBoku6HkAvQaMKizh8Xw5du/Km/SSHYccYLWFikr/fwIeT3uNbFKdige9m
6bPsz11oqksJvMo3aAPDpkf//cN0y3Pb3iVysjs2y8dxZVz9+BeZkcKHI6nHy7OT
2sABAZM2rWKpI5xtK1awOmDinP3U7fU7sc7PBse+98R7mAGK4d8Ed9V3zJWxvHKg
OQB1Zfmcq7GqEb3JMFJ2ZEfV/NdfxYCbXmxg50NRoGYZEckklQ+5dXK3XVQ3Sh/m
QPIkpULrU7KWySFk3pYSNZl2ac3ckPSo4KUCsTi3WlyJM/I9HEhMO8lSU38KAvNk
UeJ0/4ayHQrs/zGtB11xHcEoul/0K5xvIGahc0Wu1+ARaDm7/IM+FlE3UTT9tRE+
lpt5J41cF15wvu3swIDxpRL+7BrJh3pZVjZ6Ww1wgKdgJ+CdmV+/55FdWBqWzeek
Rn6KfhuW/Y093VVIWW9VRkwpCyNZEfy6tjYe2wDi96gbYhFN2fvq8dlM6tELXNHR
qhsZfT1zWsIQCCs4YHT6VQGXSzFs4wZYPNx8ujig8iZN4rTauQ65FHCop381RTdb
HiiMcws21gUqT5QDgx9anbADwWR5A7M8g9u660ldEaP9jbEiBTKPrUzd1egbycQ/
9hbzH9oRCXEqbURKgbhj16HLoRTU6bbeVHFtcNipGnIGYeQuHK32980hwCso6PJ1
u4qm5obbf2xpufZ16jDHalFLWwRrrbDrm2HXbkAcMlruzx/v2HPgWg2j7F+Ci+Ol
Ac39EaNv84WzAdIf2/Z4aw4n8NM1/czBLFppUyRIG2Q3WLdOPMhsBvmsAmLZ25/d
YpxL/fTLuiPzleoDpv+LfNMIc4Kt0DQwvsEBCT7ELjhXNDSPzx/EGcYxW1AvCYpW
bjK9F5rvwtiPqn9ZeZ8sPoCp/A/qmmmUNRvNmLHdq6gkHjetvsjJrKjpz64wKvxY
1oDtW/YtNFXRoiWgWyn4x4J8ToyLBlZz7s4N2+uy62nwJdlVjPtPo5sKHHLnDVb/
f3ZOF9ld8qntyXt0aZe7vPj4vZEUaXrOTxndJ/g26xjMN7sT/KjkXR/jSLaGrVmB
NXW3VIFFOdcJx0F2Pr/5tKbHx3z0gut/70boBDvWJb56kZ4af07dbCaKHOfT5TtW
huYobbq+6jIHTDLvvLw25QVqJBdk8NASrMoRES9kwwcevGUVa4rO+0e6mUDh3vJb
ewfUYHBt9urBf6qhSoFKaDSQrkExRcqArqgtXA0vM6tQufCXGajYCPnEFtFkF4AU
BAng5cV70LZ4M1Zn2+r1Z+NDDioJmVeB5DJghcVxGCHnhjh5hDHtn11DYMxDrxzX
A/qL4G185fWdfyugHeLNGz7Dzb9L/QowbSQqAVk/1qZkzshV/1hw5wyJYua29Siz
i5gmFRnB4p6h6eTKihPOzvEgm5UWqFKqgfd5pigZszQWXBczC1dPrMcHx3DoAY3h
m7/SJx+GsoFYS6b/Q7Bc2hqehFcnvRQ4bMW1nFlEgpLoP9RRFoDyjeDObNPbrcVI
hn9EPial8xFmD49t6R0enH7qoCYb0fW3gCzPSfhWcE1CStP5+xG/wG9ZqpOaT7O3
UtcMwYPoQ19Yv+MgucBSQtvTmoOZZFL1Vqm1fpnNZUI0u8slfsSiP+Fx5MIyzHH5
SoH4AP9F7R9W/OTzU37xWCpy8IBifYfAkula5uCubbAkqaEmwgc11FxMPOPH0F2L
LI9fSoWEV0bhDqOS1DlRdpsz3Uf5AYeAmu+ncS1h3bc38zTKXaEOBRHbkXPfeWIP
K/ZiZZD2sFzZNya1F1JvLFWZ2l5J+V3VwSvFuVzW20acWhcfjISjRngENOyV9eUV
2ujh5vrzykHUi8uahLhtfepgDo6cHga3j+TCpolGyNPWo9z4FGHDy2nYw0bar+Tv
4sL6RDBDX/MNHJL4O04Pw07S3i1MHt6qDM6OOvVHNlBMaCUQJXu85yOwE91o+8Nb
wCBAHQeUR5nitsCHrFuJCRUY1QMfuBazQCvp1ZMBZxJdUNOIlhJgPPt3mBlryKZz
xQxYzRxXitFUS8YLhJc1vz4oLtl6lXY2Rn7mBDLg7a88FxCSfo7OpoBzU0/+dhps
DgrvWeJMfK2lt2+xK3DaIDH/hDjDrzfRzn1T3h/CPxZcdzu7eHr5q/23H7vBgtFQ
uCL/AjsafiS0FtCn94IEkuTGnItV9Ji0qtSGZxeOlYY5K/UHWrK/vKF96FwY5gSO
1VBBKlDZSOgSace4rX4FzityT6stUDPnrTzSrCFguwNchApVaqQyL2xezuzRRi3r
AjdkjnbibiwVwZukWt/VOGtOdwFSFVQbJwrGiMQnhZdEbNrnm41eV+L+tQXnORw5
ny6knp8FZvyI9qraH6ypFsJ9sLsbQZhXxeBeZXIK361TWrwrBgcLG/5QtTpkqMGM
/CD1Y2xDUC1R1QipDRA86lU3SpYpk2OABlbAJyABwMFoQ6GQTFof2gT7n3pEdkix
Sr/LQTCC7+qywpD5PpZtp5PQwEQvd0ZJ1Vq4PDGgqvmTD7WGQ1NV55mboKRDHPg8
iRkmb8mTrAomdR9hbfoCH1KCyRn947RFffQt48H2QgLEaFUVhDNGOLp3mCGLo37c
P7TRJ+bKC7AQSX9oHhEDz/stnTP3Ou5tBmm76ATd/7K+aU1pXzlvNeNENOj5jNo+
wBxshIyK0jwNdwrOzwrBD/ANivIZVe5wZ25YrX/v2d5diRAyr9z3l5S41MgdpRqh
V/jPODzZJli2essDRz0SkML5HA50ao0bkI9q5wAQFpMijfYLweelcs4xyE/pC7J2
MxORTMXfI7bxe/px3JLReOsB40UjaKTj6/SX2gtj/SNZd92ew1BKADFhoj6s0RwR
Fgz7oh6JZ20hjcOSRybL6iCeDTMTcrpTofSfNWcywHAaTKkosVwthvWN5Pm90ReX
W9fhGHR4U6EhtGMJWqIt+/oMQlMtLXXqYPP7rZfqO8xmEzMTmmVASLNd8SLvjUKV
WMxmXMaY9LulDLdLj48EUzU8KzQwUu8ZssjwqzOIojWQxP3JKMEX/6qUq83Ou6k6
qaqGiC/VyCwZgyTeh/q0k0+by8afuxXnOnArJ/S28bJpZVFaKmws0oqR3I153N51
zrrzgBUbju1O9l+d/XDdm7+jejBBY1sJLL3QOMLBsx0Mi0XbzAzwj20CangoM6BY
BKe3DvlCNeoEJvCM+0EOji7NLd2Z9iDiSR9OCIsqj+IFQlXJNQMGsiLk7APJYPqt
9S/CKmU+MYJAJ0tyC7GugI8ojUST9glfIZB/cKX5mLgP5G7PNqF+W+iMOxKy7eJ1
wuw5KK4zZuUD9l2ng35OG80TqebjoPnfgVnvN3qghtOmx6DaQdeho7xZdVvNgjnq
DXj9CLS5n2JkHYbpXprv3VLah9xlOl+Uh3hz/Dgk2QOUVR6eMC0ZEdBK2vNVrxzF
l8mpnkLvL1jmHjDHD0PEHMDUagUC7z1VJA0HsC7Xq6ZQAYJY10KGplKOPdBSRdi7
B+4zzdbVwywZQZ7v1SO+VXIVKTWLd7Ux+UthBWetI1aW87BH3jkEPbicCkxkTTSI
hnoKhBTKqXXup1NjdNZ9AAeECaC0euuhRfSseO5U74BYcNpc1/GbjIZmyev4ISdC
0KzH+9CPAe0SvWNN+4as4xjnRSjoohs6giqwnNUR2J9VOhsaEVgc/L45WAYKNQEc
JKtjCwJyhMddQSuqX490Gi7lPeeMllIhzfHsUNHw1l498S/APQihM2vvHzFIjNMU
xBeUJEUIt5ffMBiaopu97G5Bdh/D9PSZRt44zzcxK+waB8HmumUuKLcGZPufmeiG
3h5rvSeaOLSlaDW31xczccRtFZMJ6hQobxjicHGiFVVfwvEAzRHbz5jzLV5v5+JT
ILRwuAkvcVfa4J5edAsUok8r97nknV1qyHmaQe4tbvUki3/MjoSKmlM0P0wpfMRJ
vqk4kkuG7mVGjwuEyBdvKG1C7nIgtshQbk02u13uwkjNY8l1fMBc4b4Di5AmQPY/
VPfvh1QP8+mSCPUDuanxYnwqWriXC3csD8yVd7AYPhwq+IPBMvt4ObfZTJs6lpmU
rmbGgEbAukEDtAZ5bddcrmJAuUR9JvKTrzuhC1fSGw/7rHOyrqoylr2PeKe2ESfH
yaq/1Jkcwf5D78G3PUimZeIsVcs8vaWX622tQ2AehWeaCg1aZUCuPEgUrkOIVMSv
E0ilG4MEzLfaEt/DIV/bjJ5iuHrp43qAEznrBG9Gcb6ZjC3QpH7fVX4El0pstWKC
Be4gTLW4YFjsP2atqep6u7DMMh6+8VoIubYzLvAoL4P7LEV6z+9DRnvE7E3NhYkZ
aqo/Zj6jOjng3CWEdf44Jc03D6MsxSXsuawwUvkiT2iz81ojCwuy9RMGpVnFp08d
J9I3ytQPG01Rn6VkrqrfAjoIziStnZlMsG4p0t51UV7PwrjoReWN1PGOE3UkkT5I
oq+OLYLSOtg6/lvnSRlB4kN3sfbUwM/EeWd1vRDL7XzU2Zn0457Lx1DbI7xT5BGS
YwEUJDWU5R7o7VYuBR2E5X4qRTewG/WxBHtD0Yn0QHDpSrSSvxfQeFEFYVg9TxIG
v6OQwP4x0mo6CdwVle8/eBx0BQBX4IsdxMebr6PST19LCXMDiXc4PW3QLCEZYIF9
JcNnkk/78QTeU1Hwvj9ch7DEgOHZvUmLC97ceA24yHwrtbEZ4Jw2G/lgefQs6aFs
r8KmTdgiFpdcRbSccUoRh1pge/VQiD58VIihzEiAUHgnqMjX/mRrvRhpN/Q4X0nn
6gmAwJOAb4T94PTw1IcZacCWlgg7Y82sP6tMITnc+6lehXwqIzUVr0vv8LoMipNI
2q2vHK2Wf2yFrLhAht4eISZIVVkXrGUrpKVBmuGa7Kn1sN4PLOh1BdNMS9VvYSpj
UluGlMBAO6hOoHQ10PsShLHzCzlEGu2I1BKkdQUENmmROM4Isb342irNbwQn8Uit
NY6n02duNsSrnr5LVP/9a96XS+jdcn0NCSi0UGxQtmYUuEERxvRqTuXzXFe//WO1
6F4jirtG/bPUM03LSkp/WxwS33ky8+K+12a86VniXosiY1AY3WIUQPVeFBIzAJZQ
A2Dnac8BHYAH/dJhDRkfNm8IWJwQHEcZT0yQ9ZYlTHVwUvJEYWNfcl/rAkXxTis2
NM6EBIlsrJCNWyNp0T/eCytEnRDdjlC4SExpo1y5wZ4xGjalGjEJW0b0ymq0RqeP
c/d3fnukbHgcCsHK9cLSXCADGTeiRoVFdrskdV/sGa707wUbF+V23/QGXMtHSZDt
q/reJY0/a04G/u57njp0Z4tdmMgWwIvG5dRTj+CsTf4p/aQF0hbohhgmV5qMG+Nc
hGPpPRDaXI3QaWV/P9msWOq5YFII5aBkkkqCNZOWMR/xq/3Zfiq2hHXZ+dmJRS9y
UTIAXEvIbvWhyTmpy8cnTVZl6GKwKj9Omc6U5I8DaQh1IbElbSJKGPhqQGUFrM3o
CiSRaZSYKuCQnuQrIuE1sGL75cTKwIG6O/zx7yudfudkWYYm657vJQyH3XVCDi5k
nl2hIBji7hkS2xv6LtEwAdwSL0zYPg2duW12cB3TwBJu6LPPE9bL6PQdkOk9KBWI
zRRo1LMnFo9T3M9i48kw/+qXaUO1rMh9LRIc679stZK3uCbnY6BbIm7kSdDVsJ8v
qm/FR7x2TW3NSU/S2DdSIDUH/1TNtLp7SPdo2aPgj+mAg5a8n0X8LpjJrL+GHrel
vWZVcLV4hAYmHHa24LfUQSG5TuKxUOWuVAX8ueDF09J+SCR/myJ8Yt2JdCUHl0sj
WvIAkU91l/whLzvl8j4JGCZscn6mu194xKpOLsRpfz0+hoJcrq4Fq7QAUI4XBF7a
53gy1QURzKxA1xieXyx1Im5BRXZ2Ni5y8KXUCJm9aMvChUa33lP7jUK8M4xsbYBc
y+g/zNxC2JJJYxaAKN9pZHBEqqV5YArDDr7U4T4YHxF7fetJmaN5qNcnePHG+AN+
SV9vlAQy+xpwV/0JV8oNvel7x/L80et97GYByXKL7AtWXucAfsie/5F4pJz9tueK
/ezAzuGcnFiQamyuci53peXhMX8x33WyolnMAMQIbX7duwIBAVbDK6e+diWH16L9
EXyAL7VEwhDGhyIXZE71qmq+y/BwObtsBQ+JuN3QdUhUDrRwiT8Z0o2lHi18OLlK
jJ+F5sV8x5TUn7dPBNuOkl1NMghfOVfN5NNuFVbOIFG5biM+BiydACAQ/8DShbXN
1lAj5pTCnrhuwldtN5EPf0TIvypPtMMd012yZ7FVHt0XkKG17BGCzSUEj+VjWVOo
o3Q1EZr8BbGtT0EOdk5Wvw7XWjOogqw4JYiMPvgvXhQtTYeeP98tK5ONGn3zKxpK
q+QMCDBilOVKgr/b7Ibh2061AAREd9VYlBwJiHAeiWQtRXLjaRo09Se/CIjyf+8X
+aucBfcGgp3o4IKaFEUbM2JCU5sBzoc62j5ed63gYyVY+NvvljHsH8+hFR+GV2Qb
+Udzj/alvHczrKvKmmCDXZCLUfuqiTU9CJMK0Pj9kW6pKyQkn7tcABIFDPpbXxdB
3Y+Bs9d3itASKhuwGvuTOpEXQWZQy9LDlD3tzSuANp2DWwLUme269VZ0Z89xN186
tZNzdZDh2S0f9XxPoxY1yTdMUuJVG8Sh3GEc2fLga0Ml4Pe4c7f5o32v3byaJ0qA
N+0+FJWDXCAyEaEeWfzPbCtSwIxm7Dom8tvX3dBAO09ALsi0kkOeMLnMIUKwa8Gp
LYI8UH+r3ejv4ueOQohhCFGxlHO+wxllnqDXpOAprGt4+PResK7vwi18j525CtNe
3gbDyTBvFauy/7BnuK1C2zoxKhRu6d4h/orXpYGbF2kQKrGBUMyzQDoGWRX1cY+D
htQNgnkAJnUcBjP2B7Yfxi945fLVSL0YCHlBeyBD7r8XWQr7vlS+c79l6Cyo6sb2
nle63i25NK4CASq2oOwHOTsI6E+uW4wUYDWGmRO/ykyBKzzlQ49SaifcwH9zKcYZ
e1//5RgCy5YB44d5COGddhaOOMQZZuCyXWcON4qgrcdrTmIA34O2m0n/t9e2/CaV
UGqAAEkde1JhhesQLgYgaFl7nlgW49fLTRu7895OFLOQd+KjQBDc9KgpI8I8UNab
P9/po2yCf+61HnfWdoL2EhuX06R4gd7Stea/aHeuftpRC2pNj9dZfL2s22NDpdQx
uv+kXK2KPHab6vs86d6MIjg7ehB9seW4L2kEURbkku0G7xAJswVH4l2yqSagHBd3
WcHSFGrCg120F3kl9rHCuyVHDnhr8f5yrlkm6a/cZpL1EWa01oabyA4acOjUG0K2
wElICaN/OwzDOBZjOt2CI+VNqrDqpyBr0p3+uztWTnjbpeC9rhsADS+GIinL7F8+
WtXeWHLzv3vYWg7ZGjaGuhV28R4sjrJufsOtteqk4VH3ZYwwLyJ8aO3FfcRrD1Xc
dKbji3BPdH8YmPVX+DKPLr5pjYz197ibUDVfKx6g7gx5dwR4/sCD4MciKjYXnw5N
d7s92xjH6miwC4gBO04Zp0Pc8SM1ycfwAiPdjjay4d46G0oaW1C88Fvvd0/pz3m0
NzsUgv7XkkT5Gs1uEp5lem4kSBwwqowDO1kybZHk+SZ68RcOVB3ZUs0i31vWV8Po
FtLwQClRZEk7ciME1WQdXx+c7hgfa9b7DO3dagk0TwjdTBqdiPhgeJ0k5VXTEw9b
dyys73Z15u546ZUYF7TDwOkeA1xffEow833xnt8uSV0wbSzx95YDgAA0/5lh9mEf
FlouOlhhwJBvKfF231+6aVLNzaBCEhOPOBF959pQkEgs1xEbMh0c0x5+Ch+0kIGG
Cosv3FqBwwtFpjUsp4P7xk/IsKgfogX7MsHjgRX6u4LzB80+gnQ5zABARbTHldcO
5lQqbnpbBv7PiYlmwXoB9D/YOL2qMM7eDYD4cN7FZWE4UUVNNRJSWPjYdC3mzPzK
ZmBB/YWNmsmgygMvlsoOqwSP96K/y8DvaRGSAs2iRCoEi1LjUDesQJ2z05hOhTFf
xPCl8oL9EIJ6wZr7P5nVk4/yZqH14qbKPr+MR/ihCjdgLmGA6PjoHWG/b1bGO4fv
9AYPdAELlFDQnh+qLcNAy5i7VQ2oCz7jeNDCNmOnokejvTn8AqZiDGhhja6vTwtr
+dnOiFwEOxTWHuaDsixzLlIitymWZFtiVaOgqOnLxFQPUba6vVB0cKGMAjPeqFkg
vPPhwuOYsWIGrMT+PYl9LVMzgB7N1IhivOjiRCi0n+B+Ued+1SuXcUSF6q8qvobF
1aHPmF24E7Wm+tYW/Fx3Kl3br/tz5gWnp0i11MVuSobFiskgmKU+l2hduh090CVw
h+rHPmHRkOa0m9yAkTgOo9Wmnq1mUWcd+WO+NlKzGu4h35VijAklvT4cKAA390uB
LXujGFv7SYNQJeYM5lv9A/9AMRA/5jmbU0ZXi0L36oJ+woGRUNY2WXnNXoBGKLKM
2T3OGnhkDRK0u7w9Sv4BljaVIb0z97tovYz3b7LPQ0J1U0sG4t81aR+GExBj3WRr
KqzwaGP4twynp7IUSOGN7P67rMfuAuB9nOtrKzqeYeylBDmc0Xcs3dcuTZvzdwqa
mlkcV3dO0CHhQQaj8Twp/U+yoNAjvW8BKq+ekn1A/ZdH3d8NEyGJ0Vl9nCiyJ/Q0
CEGw1L8SUFgppZ+1e4IX9hIVuqleuEo4CflefTfXMF9eQ/Zcx+nvwbuNSAZIDRX7
uRYoEY+aOMDdEigkU5fuKI9VrfsjgLm9nO9cgJIoPWnv6YFHk5CYll7iBXJy1Wvv
l3xDsn0o4Ncm0P+cHnHX1PZ8ffI7XOUcD+l8QLKbMiOvbovAVc0lq8G1W5rUn3/w
0GgE9pCMJ3CC6lznxUmVcU+EwVUy+zF487fJnkTqAr77KJa+bld/uNSH5U47iwkF
WsGaYFhV4u2igCJ/wffs860m772n+BHe67uEnE8dTemSSCxtrXsSJ9IKk9v4rPxY
S97P8f5FdnjkovxJ8qjIVpL2V8XDBSTrhBXx5H7E5xnpmXsAK0KWh7reT8c4j0nZ
zwg5l6OT/qupTP9YM4zo8sp6xLc2uGiPNjnVbaD6iLLhcMMPTjk7Lcfp0D1vI2CY
n2+1Y6Ffo+2P9/yQwO2lwJd6Yx0QIlBiLHpE4pnoDi6iPz4OX51ytiXuolZkvOAk
NjS0GsHlWn4Nq1kZ0BxqmFDv+qDakDZUHkbIklIvKGG2pem5fy9XQwuNyh7syyOD
xR38w0LopYEcgTyGnCxSFr7Dg01aJ3qUdOsNS94jT0iBXRExg961rwhh8Iv8sbho
KT2/EETNGqiQg0HlJB9lukLi+6aju9CyTAfWlQIxfLw31kLUWH0m8K9Ioya1YB/p
RuNsjFnZlQjpatZv6YOramrotcrDOcir8elfInXWIQFIOCp/rhlC4UGDM0clsB0g
rxPGRLC5B5+6sICV1Rk8PlG7iawVWQn4EXQbFVJcVXvCWFWBLpiUuVKL/EL68FvM
OPKtOXSy2NLEpotKKnUj27FVdzjWd0O4bE/TEO7ekq+XH+YUA2D4I4hPU96Ziwy0
BDFiR+VYRr1S5OPfRLqjiLUvnuUpRye3NK9wMgWi9f7RrD4iBJmb/6r+7Tx2YP/P
p0NRI2YBdpGFYMsseSBLmtOkflCFYgdk40qg+6dj/9NVhZSEfTBkXQAquWVopKy7
TQC+FWEOBRqYDHEzIXzbmhi0YqubCm3qKIM4uFkkedirPRii4wn5hGP9+rCaXR/U
jcPZoi9FV2Qw6/i1TmX7pga4GadW2PMRj8YzqDvyp20/bCDuZbmLVvFxYR4Qp405
ODsIZlH8UTlVo4XdMdv2WGlBXGFrjou9YutAdYDv0zjEiBoBgY18FWVP7PvnXnRK
VSgZKQnVoaMynBrOoPj3m5Gm5zZlxJKZxzA91/2jZvQbcOYhMLPSK7+HvPjD4VN6
8+9vFAgoXC3K79bSqPMshCo6+dPVVQPUTWoPRV4Z7I8DJ/FvZ9EeDwIaPdCjVlwV
taej+h+c5Ccy9cs+MTQQZ/tFzmR8ZsyaONhX1AcAXcHcETF/nv73MvpijwgLFozJ
lH/2po+vqRcUyJrKM/yM0VgvnUBlVgnWKE0Y/T/3r5j6Y4eVvHuY7AqnI0U43JZS
aiz/JdcSgZxbN3PeOFbO4s3xD8FcEo2coHqfTDhMssBLVHiJvdUhVHhb2eg30qUm
AWvwCtoqzhbVJESMK5CGswq/sLZIj8A3tQkhPay8zceBB5Adc9nQSYn5Mlsiz+Jg
OfBXfE8rFtjZfN5c7DAQATmBvRLXjfFfNC77DYAfbKgB8RJhTM4xWSdGbv68B0fk
+Yrj+Ojpf/BSLo86hN/RTE7AYk4oNmIRJUkO+ulQfgWwcfofKJAxeYAvRuzfJM/U
8zSBE3mOL4KeK1YXbkX3DWaJ9iEQN/WQB2M0IN/D8fhVIJBZGlwL/olKDOyjF47p
FFjV2DbXrOzyvMc6JH8b3Xmc8izhLqfky0QKop/3nVhxbNOmJC470lzDF15zxGLf
TCmmYnnPvJB1uHE67fPOOXFiBdyhoq4uHj9gL3g68G64wrOlqBaxMWa8jxe/9zR/
0cm/g12miJhMFVkQXC50zTFQCXdTpdpcvDm6I7YUIxQ+wPXnfuMqGHOdki9xRVw3
wZZneABhQOGP+3yA9OQV1hquSvshiFtTUGt1636lbLJUXVsdAAinfCrpMm+wBIrh
OXlSAFLYpciSQCwMH6wzgAEsBuuk9uzfXNQhGcs1mT9B0jTVCRZrEJCbtH5pOa2y
f5JFq+IRFtWZ/g/XEyNAFg+m6+z4u0zmzFhcf7R/IXBPVKnO1Y4KiDkrYsfCMUV1
HhhegcNSTCt9lHaBnjFGDRW1H6JaWfR05uZD+iSAE0FySSTaNt/xVYSOFIApG4qi
A990mqOdOR/zd0H5q3SgX/TBPWMFk/vUEC/kqrSoG/yctpYPCDoVCEZrqFeh+BNf
RRXkFtC+NUehDHhM24E2KGeVscRUYlO05tAeYR7LD8Fv4ZKKAtfA7wK4BlNgq7ff
e5JNRsfjXMqoiiGqUQnrfb34P1hsAcu0YdcEvu9jZdcrDzI68srjNa2QFA6unSRB
TGS+mSvusexVLXfnAS9Nmc/CSvP3tmHo96pDeBbE8GpdoHP2l5bE3vB6ZokmDxtM
D9gceiQRXx2B5VRRtKN2fOkg216AHEhHspneF7qC1FO9897JFoK0O7Pta3v8yl2B
lXJQkK0RkHGVRj0K4GW5+JEkQjjHAubYSU8Pnq1VjES36WD7/Bmdrs8nixLfJG5L
l1DyyZfUB34EOWqshZ7fNJ5AqOEgTD+DL35J4xUWM9jbW5wMU/jdIiX8nNvxahYF
5rOdLzs1knl9ddDxlIbIoNeuUFRH1ijmgLc+4I7jBUaC23ZZHh8oMrBlSJmf1VPd
0AxByHBAakzZRGyRp1u920jKhaUJ28FF8JyAs5LrBR6yvLW9XMzGYlmRQwWGSVBw
7x4V3TogWu2uFrjyN/c1KYsagcAu5SnXpW1Az0QrLlt0exHd6YziJDKz7zF+EiEz
5cJe7nWCQCpm64CSKWK+blgq+MYdVaQlLgAGxsa6sCHaLTn6cuJJpzoRdf9O5jKZ
fv4QmAQxR06/oSqrSsTHxuOX1sjNXNHQigJHtQBlCVgcNykd+6d5FCOsMdinE0kI
AR2HBRJ9dzFjwFGjKPIqxIKhu/YU79W61nTK1sgu0omnPZrSLVQI0KgNhkKKmNbY
oiNkDbYnprr6P4Gxo8EeBXeauvK38AcrsBw9pSfr1EPsZbaIbSkH//m7kArbMhEm
x/pXuGNm1wSWbdf9Qskgck2NTdioeLSL2Jug+Bf1Lrkl+gCA4GCq4NhhMn+KbeZh
Jd/rlU5xOITYpi+QDvpQquivPCqHSSz10/6oKASQcwM+XmMrlEowJzoINV5ovllF
VjbzUHg4GvqtDl4F/pYkFf4HKWFzvmfdNZMPARx5z04q+j1fHmYJojZ9GFlXZlEh
i21ZNeVur+Bwd3Lj7boSwa3kUoQWLZC2PE1m+WuJ0U/02/Xa6JoP/IYm3WOwOLJ4
Tii5U96LZQ7u9wUB6+rF+M4Mm4KDjOt6yXDpZcqKujnx7WqTuGXpQez/fOA5m7z5
XhIS0gOORsmMI8EavoSl4uYVgtcbbqdabXr5fb2lfi+80gI/tvSFAPIZD9Siuzlp
zR0vvr8vIBGT10jBZQeDZ5QAxgbV4PUGdZMUXBGKC9B64b8iQ2vN6R+le+d8MNtV
XdSuUCxIA9zByPoq4SHU/4TrEE0t+fYjk8Si2UxCkzJMGt6AdZZ1wSwe/W+j3E5D
sarQXVXK8KzeVJwtKaVMnyReXvarRvHT9rR96o7mmBK4slaWo5r2rDENkAkPklRe
ukLDpBPwoOluv1xz/A5UXCvjtj7jdvJt9gdPdyCvRNQYlzrTGkPkzcWsx3A4/ZAm
kHh0reJNxmye2Iq3DVyk4iFBA56UtpS6D+Sem0xFda7DnIaPYzfGW4bdGaPcFAMp
qm/d9Tcuxww1QwYthuU6LiNKCDrcE5/fKp/enQF+JUy0xf4EMpvlsW4t16lmh4AA
Dzca+hhN6a3kiBHHDBa5euDc8NfrJ8VLsyunY+8j0enGkxnoSa7bGwS4IrFxNIRZ
HiAXIn/YMDEhSVbCagKO7cmsBCPyAH9BNxKiazw+eWc+5N0rlyuEZld2b1ke+/MP
EZMVo7Xit3FVTkpii61FDLQKvSbt15SasiwvjiUIWvyVo5A9yvPMpxEIp21nnAZ1
3p4r/kauRXwbZx8DmkgJjvtGJjrkwr0LuypCi9Pc757xUYP4Jhg/5eXnJYw2M2/6
f7QGV4KdKK7BowLOU/opsAmOANaV+rKMeZN9AwpclQ/ZZpfec9D4s8CKEKew04lt
tFmLwP5uQhXI0NvDu6A5yeFNzrsDeXuJw3Vsf2xjoAZ8niRORkYGRJE+gb4prIWl
DILvhqcqOIVfOY55qI2FJbXxxjhMlsnysZhlMl+YOXY0Ykqx9Pirk3HJD7z18zXc
ABk8stHxJuZpFZqdvwFgemAR8hbTYoQU6U5r3+SN3NazFjIbpt6YuYE1hP35yHVK
SDjoPcCJl8zI2bzVROL6Mjgw6yvtJ5hCNHpRfHviJgjrQFcvQjX3qxR+NVbn3wV/
0YTnBW58Vsl9xIPfAM61dFjFZRDHN7pzpdtcAkXXZYQByGmZJKrqvjAqeCgTY1r3
nt6moyOAg03mS9xjBK4RnvsoukL12OwGyBd35dcfGYbnJZaJnBdydIGvB6DKO5KI
bJhT7gCkLwNak1Lf9wTYPB9nZLKwhZ+jqoU11paflaLTYAR9kgp68qhpi3vHPQAl
+s480x44K35fjyqPzCfBpBUCq/O4rRPtC7y8pfxUYJ/ISBUZadBet9n4b9PTA/KS
xwV7TOnWpZMCmtcUFsxCNpocBhpTTEgX808f8dAkPwEjhWTbxFikxh2m9xo67/Xb
Il5W+h5+hKXx8jMIrjJUateQNIGdn1Z8x0X5FSlImx1wxYo+I+78x+2sw6ss8l7b
xhwi3pclo2tCYdaDPKKumkbgp6nnyJ7n22jdTRysWyoXqKjx3VHTEcpLaMBILN76
jZ5jJlo2Spc6pnNUbMmBhuRTvI3n6cvsy2GzfVKk6YePltxBdxO/+s7j/AwakVPO
ylhyRMoY4SrSZUkoFqnrSrJIUKCcZN89hTrlWuIF806ymvXJLVBdTORsZL3z5zS6
VcFSggIl6/+dylch95/gz0VrYlIpYSL4VtBoDu9njH/g+2KFALrcqJRLvyAfEIYd
Gy2LzpC7aluolbGT0MqPx4jGqFXK4qQMJW81xfUmQlTb2bbeECOgpPO+D1rzDWLm
1acMrssmk/A1Yen6dMWW8kwckXZ5qPHlP26FF7j6jw4aQvUseFkttrXVtCrg0l+X
MKLjHnuPPMe5Kf17YjVNxnzAbWYcQ6e91bF0HKIc7Lx6kShhV35ZYBtOdU98ZSLi
YDi3ipuZT5IQ11c9qJy9Y/PFoIAEl7MRMNq/poLSoqSPHzu3dumVZ3oTI+MEVPBT
M/CNduhgPPgWPrfQ5ZQfVCNKTsKQBtPDYzne3M3qVrspASNFe82jkKsqayzQC+D7
QE/Dbn2EuvAEXicw0pVrYp/w5ywnEjXTeA1y19TPLQGjxRCFjHAESvPLi4a99VGG
7OFi2z91S3IyuM2GLfOJKKvy9Y0mqO8oioXn8TrRNcNB1DJQ1IOhAZNQwhBbsJug
6gcFE9rrs8nos2+ffViencIolhnO9+gwLuy729lN2fVTGLb6FJQ0VAuuc1qXiLua
LyM/dg9OOBcWYSL+s5gojOd9K0PlqW787xorMZhzmwK8dy3mEByEN8kVMHDa3jF1
fkjktRKoKGQ4dF3MsuWpFUHcvav/zpVKB5mVN/8rOeMa6MjJHkhenMoCSbB2t/Ug
r1ilBFcH+R65+L0+n/aa/ZdwFgOZ+n0YSPWJXwKdfw+eDatTAerRF94t0MpxPAwJ
zBMAhHe7noW6h1ECQFehfQ/Lrolbk6JPxwbHmdXyGdiTklYaJgfMlHCW0xvmJkVo
RPYQZP3hgJecE9+tk57eFYxejK1mO1qlkXbPvwOBJrfyEfjeuzRZjKstblkiWZRr
jDn3tRw2aUc16ORWcI9kltpW+CW0jw9p1L4sx2pRblVfpfhD+StYSAR/8mfEiGt0
n5Z+biJO0XZt4EGL2HcnFmBE+s8J4yeggW2Fwv3mat0eQNRRoorCLqdsZQ5P375x
GEKLuobqfvQ3fIlZBGg31ObZQQhQxTO1K1gvVKlTXJbyMxI5eYNf1wWnstTCjcB4
KdjIj3yeZzv61xkyPKVRFuBo2yktmEBR1XZd0HibHCm9dsPGOO/L8E7dR7sjK5o1
NCqjCHlKObeEQ430BrJTD27eIilyECUvyR8Gy2t5xX1+Rv7MILPr7eWhUrwsLAHV
5tic6pHmPZM/SEHmu/p/Nsv0YepYm5YwzK1b3WLE+nLl3nrxm3Qd/G32aYo12OHv
Fwqd1MS4yuOrkwX03qqZOl/DhhfwvooRUTw34yaPmpMHkOnyBWw6q7O+cPLIK5dM
6E+jGvdsrN+Ch97LQQu8+CrCHaKAhthE2ejaUi+e9djPAU/Qf3Zv7zRUEyV1g+1M
FKv7ypDFUiXsjMof1BLzpH6NUtBWFTm+gFqej/NlmGZDLFTydgP80rkcViRYZwuK
V/Wt7h/q1IuFSrZuFVuBTTYmTBOmDbi8olj6RuH7qJV6oTIubtd0j+gk2J2e6kWL
xVwTbxU1HO1GeVuzVeke1BGDV2Dqzpd5TvbFpmfuT61HGPlKRkWQ4FbsgkF/xV4s
3jynUuxgk7JuZPW14UqgHCDSUwk1kjdgYOiKOCKLN8qboF40dLMu8PA/vQb9p9Fk
yDJB98L6H4Q5mkZRdEm42I7DbTly0ci3YhCM93Aju/F64ohgLWZDsWsU2cFOyDSV
pqG1J6wjN9bNEWLrba8OF+WL0V0JUf+cyr05fUT6fTrIkI7jeqdWzlb8HH7fEVUl
zAMBN++EhIRpBwPBUhg2yHGtGJRuV/Wm2C1HDh/RhAj0s99iRH4XRAquee2SOZXV
eFQPdzUAaEycUy+A5K/I7rtOlmgcjfKvZE5WPnF3FNiXv277ph/FK+bbcISEcyYB
n8yiqH21/eFEecMzd4Ms0g4egm4Whqw5G9K3jTytry5eh9KSVOws+bpi0YmyX8OJ
8karcY21glyTEUqjGw9WMvAHgg5n+/5dObfrGgFTRcFQTVT+iYmt42THBVxrIkXx
pOdMs12MM/Ha0wk9oqJ65GSZb02wMUpvnZ/hOYJOyhBxuUbiXoKmqWC2vnznQp1p
CQBHQm3r4bZqhz2kQHECMK9JB1P4zOD5kSucYlpMnSLHqguDmAnnke2PZoizv8jt
YFg3txNMwjWRu/2iY6miDuXTHIfgs7cmaIc1f8TydcF6ghMlsFzbr2Ic+KuZiUYB
Vn/R0GPkfELvuK8eVi65bsSKZRIzGMxANbK/IDoE38cLIX6aXvd0aRkolyvWAKzR
MVhIuwM/ma72I4xhPrdKhJxc/YkePY9AW5M/lxTqaiQiNoECiRm3drM6r8S5EIOm
PI+lfqq7PZD7Wq1B8E21ReIE8onvlF7utTIZnU3aSs/7GV0SPohzV/WGik79uqNJ
NYdMgn7AaGhWLwcNhLXZ25gRNlZZhxLSjQJ9XjgzfWu6HEplqWbv2rWWscr9p7ZI
AqNUrERGZMN5bT5WVqnFQyF+CvuxU8JelI1fNrrOykfEeUe5eetH9Bn5Z1bBgzKi
ttpTxWYm/3TQk1tpjm2N99rvpCnl5T8TLcQPy6Ek7U93aZfKHwS6/QsUSwi+Bj/N
Ha9BXXZY34uix1P0j9UbYBJgKL1wQa95uOEDVkTA/7RBLFtD26lZg5c15VlTYR7X
cxOBE6cUNVwffDIt26ZdEQdcQiaGpV/P6G7gDJWHeulmUDTg/Tn6hLH/3+6Zokth
iSwW6yKAVXM4X1NdA4muW5Fg5l6MljAgrCIEUKH/WCHMByTNIoW7UsRhYNHuqjDQ
mj3O0fIfGweAWQyKXYdepAgZ0p93BfTHHKi5U8DV1+/e0pZU2UshX/fwff39TPT7
9QO1jCBWEPaXumldOD2FPj8wAMo44yKTWqj/KKlSGCl70YgtXFzR4pzXxTtA2ROt
hSrL7dLjLlVmNQR1XF1fDq2Vo3IPBbPxfB5hnmsb9r7jpW4CxOuG4Wdg5HYg+InK
on/1GnWB2TXH01r5mNqcnu6kM9qcsNSEc22r1iPOuoxrgm8UR1xCAP9kWzE3uiDJ
D6C18P+7doFmDAmdhH9UjTqcGKsOPtZF2qEvwXFZ0HVc9uoZltX9JwoYohfOxRCG
4P5Z1rsM7IFlFbBBXN5o5tp56//U46NMahi2/069dW6jYRdkcCSO1xj0/BqDp4fJ
1sOyt8xSQ3sW5qgghL5XG5/M5P4IhFrB7mJbjhdrbW7xAfdFKYGJ4NhiJ2R5Jo0w
njy+Eftt2UosKKDLSWlHkfVZNzjPvbE9gSaq0vhxxpGPfrymbpq8vOfugsq9Hw1D
H9I8y6mkQh7erCxi3Z+P6lRS9xiIkrLm2oWDWKEHn91iLn9rNy7AOw+7E7CtoSVB
suaQz/851w1VOiUddQmaVxFyHI3CGavLtcJB03XGhatZ13f2YyvH1K6rbG86PyKP
wiU/8Bn9uVNJPN/P6k27xxMjYJaYt6M6hn7dh4EzqsLuMnv/l7+D5eyD2ik0XL2p
ySUeB7xXmM4+DVkRVljqGYRx8cM8aWJV/7JHxywFc1gDSIDnieXG/BmYDfk3H/Sn
618V9cvMm/YBIpvWmovYMM+LfEmd9jHDJV3yxjfFBj6luqw88T1hwm9IaOPOhfH8
HhdcwAW8omEqrnL2jT+2j4rgOVJtcKuyq7nHAJNsdAlZGIIK35u4pi72uPLH0XFq
qjgbQ5g/46kn8+lNn8ZdBhjYZxR4XCUpN3FoCl+DVvVJlP5O0nTp2gWvd7TcouWN
7ZHGKOxBZrcnYsxQKs3Sf3uoGbVnTVTlZ0cdCE9X6bWflu0FdAVs94H2ToUVGSGN
DZN6KHZCpx+T/mwZfIBG8cHfecSYjqllXIRnAQMnCn+pM5nyenzudvkzoyaD8Jou
4PWM/W6zzwDGY58kIj1mDJxnvyG0TOkQR+Apb2rEOMQ6VMLVV1fIjVxNwetZaaoN
zbqHZIjOwTn+rNDGxq4ex6OInwRp4XYT9sfw90v1FD9netwurTd/UqNpJSy8CNiQ
8HtWbN/XAFOXsvZaKi7kIV4LX6146VEH6KdgI9RWFlzvbSHh4LO/nDE65R6/Jxcv
NZZi5UkWc1K/pTW4xmEZVvIQkNjazWSRM7QMpzk/Oslr3IMysyo1Y5f7YGbePkaF
R7P5Jbmue5eWV3L0dOsUsZxdsdWEsUtFX4cbJZi9e+mtpZjKeLoYxow7lgolqcIj
YYwNl+4PHBwvCFVGOb03fmkbjQnLUPssfQc41T53QpbTnJzrn/gDpBEwp1t4IqlH
QMqNU/C9btlm69H5DJxSAgvJjQeZbrYNik2nOrigx3hiXAml8RF3vLgaOvg6J1KZ
tkzZy2rPUUcdy7X4/eRHHlPueEWQ2TwKKatSrcIZTGC0gGrfyk9rD16K5iu+nk6a
6/1qAscbFArC7f3jA8J0faVgPiOV29KiOW5IAdY5uoolCxQMKATCyp5nf/QusJ5n
qyh/U14/nrDuJttUfz5ayy5PR2pgppF77l1AtlVVeh9Ytb+w0E6l5HWDPnwSWi54
LDXb2hG1fyn/uzVEiefrR2WF+B71GKQOvqwI0Mq84h9LXZS3Dy9ycRElX3yv0EGZ
g/JPlg9tSHHEtbbC4XSCAOW1CuhHxM/GTGiGXz3E6rHbQRZdwx0LPGaTvvHAVdqw
jVXHoMWfzb5rBsbLR5GrXTL0GOrqGgrFvz/NPTNikAiUMugD27pVt+JMmShE03Ii
lNVxgA2z3on+YaF8JlJl1Ls1SA+mpDfpZFtPTxeYimLeKnq2QT43fk11n6+bF0mv
1FsQ+pav/j9eJwIR7xAyXyObO3gMSUFzstxsjTT1EqJf2dCsIfo10dabNpElHoPt
gMHcBB17IEA2YybQyE3TENYMpoTUsu88Py2gvI9C1bhZiaTcpAIn5XBBDW3Jb1Mg
9CHiTIf+Efjw4ROeJd5EvvzDjAkydo6CSW6nrcKGYWqC1vUALUVDEsqK0fCuH9St
2qW9PyP4UnhGHOL3X5sHK0g20qBOWKPJJqB9f5CZuYQ5pQIJ3QuTkCoL5PsUhAiu
RX4JvBOe2nmtPMM2orZgJRu1fgPMP24eQk2W0K4P1xPi0Q6VKpQZ8NoCsy0VWVTQ
NrrBtydr3jOP02K4NPWjxio3/rlb3kdZToS2KDUaBjEguM7rdAOLziNrvZ0iK0er
6CQFxoDJkKwQGdkv+XttKWPeKM91oJUCyZhvryS1fr8s3o+7fJxnEJHOexH2htPf
esIl65XxmakFppUpCvL93qYjsy7WQPIjaY2uHHsaA9HRnkVFFkA+aloei2NvFQgC
K8wWjcE2Ydl5iFWHDgUd9nedw+YURNmntQQ5WVyJ8q/8ph5pgZBFL5Er9tzT0VRS
tSILl2E8hvcP/4lLzuLDcAOwQBgiJ5GrYLKLpTkzS/wCHvYvS6QaszuNeof9Tlcm
U7PIa9+65dktKofohRMazSffDtwnn4oWv4d1dLqQZp46qAvvamcwdV0UX2aw/Zx+
BVScleeS1tA/pa30/VbTsCVH5oVoONYKWIjZU+Qqd41AWJUWxeAaSHhqXf3WlZF9
vZFeRKqCWX0kiXnVeuw1+ev3AkNKFlvnjwuN86jBWwoIC5nIOmZHGxIL+KT/bA+G
yNPuJhAnjxQhBE4N1WUVF1WfF/D2f08FTEOPlY9I0uNXzRMkDcAdFsZlDj/1i0at
0re6Cq2qSU/qQZ9GivNUY5PWUZ7i2Pgxmxvl9BdBESaWsYNE6xLEFqLbyYt6StCE
cxtw+jSDLxUh2/AQ3uXny5zEi6VFvLVWe4VblI7q7d+xtQtg/tPkrQHE9evHpf0t
EYqRwMv6lQZnuZJ8zXjCOqimWOKcolT5cwGhGY1X2d3OM/Xmp5lmWy4zj8jFySdu
XAYqg0/jXgTg86qoe0NagkfcSy/yeOaxPRSsuP8tK5+Iw2WNetyRX5CRiUu1nQSe
njF4xSrxOW20h9UPLvKVv1OM00OMJU6y6r/sJazsDirfRIWxW0LNexVNremXY2n1
q3cShWEEBOL96vVWmB81698DhUB4IJR5mfpJyB+JCZanVgMxqlIu3UAr40VQbCt5
4rgGIZTLN8/G46peFIHFQqmDGlNPRJ/AwxqWhDnLV02/WRyEaz2qJ1/wg1gwGJ2Y
fTHNWRIBazvOieDVLc2svw8iTjZOZh3rf9t/HPvxkb9ZC1d1RFd/i1Pu9FsLUM7w
6wMgd/f2KM9Lgut6WwpsR/B/OEBvV68ZlACCxxdDPRNZmqnMJobC2KN/ACGSEkvl
FcsXONIo81yS1tKa891aemxHpfqkjFFcC+4CJFuzdOZWU1SkhKop6QNrskJX6RGr
4Oa7mZ8xgj/QJHIEkwX+SjzPwy/bg1WZIfkYkQXCR+QTdZdawzgiIGWr6X4L5P6k
BSjWPKJAl1eaIGTT7m+SFhx4m9qyfw5GxyVeTklvedgmXyB4I3gq+5IJh5uJCkS3
izkMCLhtk0miVOMwajdpO1Ao3N6p3PRi5dqsfSQsadZ9A+6+8tW6vvzshfjkU7yF
dA/nmAi3ZVEscHmXwcTkbXrmWFcU99yW3mWi1AccH0xWmBJx6okMwOwgWbZHxWwv
BeHZMLUy885+Em6/QGH+3kczbikUj0k4wjVPkegJV7gqOjWixHDNMDA3GzsjMR1V
2F0WunOtrJ7J6gO4XrQHJ9Z6/jppNIG3chM/g9m/3yBZOO4f0EwmvY+EtfvYUDfM
Xr9+ori7SZXzruHJELuQU+IEDXuFpsFJ2XYClPQ7oRMyI1oUbzTashcRuUT6tUa0
wA24Ss8foCHGHpLrWQKqMLxVzyxYl7vDLL2zGh9jU8QMINF4eYwON/3GKoj4OONt
/NAjxKgufyb8BaoBwSyI8V7oGBcEOtCR6qsZxwVukziLtGfO5O/spVGEIytTysXG
Dpx8/K1BAtGwghhrO2Q8/tcx4XLMYaDUDvmRtt1K0XnBfGCiucvs4XWfvsWxoLoq
vPHKxqdt0aWE2iu9O5T6Csd8wBniAg/bkCXBXy/3qgyHRc1rh7FEtd1Vf0BFDLWk
sdQy2ItbrV/s5MKz19UfdbbYiwtcI2Dh5h0qdwaGv7wZDFy5YF5pDMY5FyKHPkG8
X+3CntPsQa3nnx6Zlj7s2czG4BSQVn7S5FCsv+se1GL54ibZatDRMaDmTGS0Samn
wTcVXJeKizi9k9XUnQpH8f0wm77SErNSx0dXbYzxJ4pvPXiCKJZ7eEcv6nvZarDn
BEU/nI1jplt5BwLjrtFIThPll/muqMx30Wv/sQt7Hyq+KxK5vmfUAJXVRtuYzZYb
+5QpcGQiPIHVy8FwGz80aABUcCZEb/p4nlqVLiWUAWOVUNAf3eN7rBeosM7RxTvL
0zDM2vWyaM57d/LlhsHXUVfmWFFR6vr2uIiyIjODy0fC5jsU0NQwxoEjfrHMLkiy
w8HarMQfI2uQyFYXo6lFQM687LaXZKYTaUA4wuBVN9S6497+VID8IEVtsnmdWKnt
bR1741936uUOWoqTR7Y+1hHZUzCjYH5tyxdC0sKkpklj36k4HTtKFiuCKFNr4db4
YrRrl2CnCiGJYEzoucP5U1Oygt48vI7fnoCp8ZXq78jMpc7+iadLEMISC58BmurF
W6Ksodmc5ZAxtw6XF0/LMJ90dt4dehKmJrrkPwe57hN5w7pDcTJEfCZYVgmzac3v
N9YBxDuX4BzcH3y37p7a77gg4mc+IgGLM/ibUbv37q5OstdQK7KGkocuaIAA85J2
pymwwL4XwpMgRj5QQgd4lJmQDEcGnTnO5a/2iwKtSdT7RNPXpXngKZ5epxpq6FgH
GDZCJGz537Ppyrknkt6OJISdO2jobfO6t7gTeffst7b7K7Qm/8onaHbtrPTVxKC1
URzkmZL6B63ZY3TVH6xcdC9qdrYntfGPbRgHe9VmffwunKgsJvaVC4njewfzGicB
cUaEqbCROFSEESoBZIXeQPEo8THRwzMR19nhnOcMMI7VpjWaMCRcIpv5BzRt5VUp
FS0goRKJHLlR7pLkrrHWzBj1ffWkYtzS/bMYL16BsjgIjxiFCcfT6FJlxFIgrBbv
MuuxatrmquSH59c9eexYYcUdDc08NqntZhYKJaGOfUcYHtoXt5lFIwqIpZPHX6hU
0g4co9CKO+8MYIoRbR3ft39XO8bZjsu+i+fx27fNsPh4Eiqht0k17ck945LO/awi
EHuphuWBDWdpXDjMjKFQIt/NyMnF6//nIuQM3yc0y5WZTTgdEiMNRQ3DNG4267v9
gP3SpnHMCtK9yyUCJTg5kUtWWgi/FfZd7yocHVdyX9JdCyk5fTGZYoarqGad3npH
vuJiC3u/z6fnxcRMe5IMy4loX0dAGvr3V4RYLw+4JsBL6l8HlyZE1XeJK3PMSRIz
V47ys/17qTzCo7kmv7GjfHB8RYBS214zGaS8bAMhqfm9sQzWsc/FpQvN0ZR/Ad/H
lktyOtpTgjL3B2M5xw6pzaXO6a5IPeomlhXhNA9e9/f34RBtxJQzAVYrIb8bbTnB
vYRKOkcnPmkuvw8y6kpm67Xt+FEWKBeMc+ph0h5322tC4AhLbfNibCTH5vzEuzLV
ODIZsqv1HD2/jS2c1EGTbXqFCEu8uVJbXOx5h9Fpe/7wA9wmDENj8RcOaUc7R+uJ
gMwyYe/25T8bo7WJEqEkbK9WslC3QlRdenVDgwVTKMCw/wEY84fVYCqgN/b5VKeN
s//YUFRMo54JY/Aocd/k5l2rrqDBwxHyYk9UP+hdQ55RTsMQuxlXm95yCZzsemwy
KQJlA3hOBmrhuUvfJmBXPSfzKnuDybcDkZtYHyBFRHFxldadG2UFMzjsLBp2fc6Z
He8sHSFXmKB4roSomc9xpULtxnMSKfgPhs4aR28RFwq1xujywuJ3L7M4mMb16X3E
xfgJcpUNTEwm/Qg9s9ZuxXKzbnYhntFyRJ9VkC4OAh8wRmyNuvMe6ADcLf9QSvSS
b97Iumw/jb/QqIAbgxEUrvfXk8i7lqVjh2QLfsUyEROinbflBGb1ixkmU/bFXsdL
y4rkeZ6+2fQyW4kfecapuAAie5J0/yGx6S81Rn5R5/bYVW7AxmLxBEap6TlrSWuo
WJarMfYonvbMTDE3tZlV98WySmuZv06+BIdsDJ2bT1dQK5rH/MxnZDrcd1X+J8Pg
HXzMlaQFqs4WQHlI4kvWukdsCL/zi0pHZxV3pkQaBIcBgTOJi4B+JyF/OOetGlvB
RhMMa58Xc/ivUwgjfW2SKuZopps1DVktQTP5racaMDo2vGNDM6e830PozUtBOM+r
K3jB4CZNBjypvjnMRSluCiDkYyrNML6X2ZalDLUuY9+S7rNj/UVl9MrbkbNi7nXY
4C/9PP6F2LrH2v5pFYNb6GyuBr0Der76Og9/p51xS3GHyoRibZa9h8YUB7a1aQ6M
BSgzRJRDoPwtP8Ivni4c0phyGGJUXhNSKCD1j1P1AbwL18o5N7muLB1G/NBpSNu/
cZbL7x8iAj59110L8jAz7fJWcor19fAkZK3m81SrfYjZHud/v0BxEBJBqxVsZC13
tc4oyhphlHVZOBvTdTl+4lIFP++84X5lYPSytAX+YM/G2R1cofLHvEv+ZTpyXU/N
D766vSE8QV7YKBz/WzLySK3ZNkA/PLk8cWBufTf8rxCId6M3cY+cBpz/0J88iBam
r4D/2hSiUbWkkW/uF1HmdhSwvg7+2NLyUa0q+sxIzwVOlkLf0t5xpcMQO/Cuydlz
ee6RraVd+7fEHsN5PIpeVnub8tgY8i6TE3dnClN/0IHbNWIHSsAkPnReumA7D1BR
FyFxoFQLtirNSlM8JPB8R5SXgKeAst4DHnPK9R5Vg7xwnjudzC3yYRilsvCVh7pc
57h5d+zXDfWfpLjQiKkgITbweBVZ3AY77AUpkF0WRg8oQI0EstE/tZ5bfo3wayVx
KbwKJamGheL7Y3xAu+Ia9uOmklXds0kAtTrNi3jklN8ipPKjIvxS6e3EfWRspQVz
8kOO/P7ZBDgq0a4zLroKi8z73xKPK11QLLSzHolAVbbpFV/Z7+y5aOBZuTnMF4rj
kXkg2IAeR7KCwl2t7B3yjO+SonXpJbT/EDqDA2wXogiPA4j7/tqjxH0AgOJYgQjE
+VSTW7AMEtyiZd6bqrVghf9fn7FfcKIIXv+LkIDk1lIy8l9xCaLqVnrEBXtxxErg
xkcCx3DvsAlFiVP+BYI2QN8UT64i65vAi69V/D2CANFagEh+Iuk+OxbUDPeR42kx
SIt3MR2SCvadggR1BqGCv5/Bj0mUQeaywqcAonigcy1Bs4Flv50ns+17b0OOJaPh
55PY3O+dMT9QYTad7rwRSCeO9jZjqO1/udKDST6Y9e8nTbv3PA5+AMUtCAbOzxzs
PZ/GvDs6boRITfdKqLavZsykeF4JXqXsCfTejFg5nJyNxtG0ElrvnOLe6NiQH6V1
Ug9rLOgpI5V5yvuUPVtipsXkdHqHQrjPw/Kq9+uNWU4dEBwQmV650OwW1p6ZCkpn
fJvUQ+8WZe6IAHGGGe0c/V0+7SQgTCtD63FADOFIW0EqVofA49tekBFzp3eQWVhP
CdhnoriBYs3/vUQSlAN3bl/9xKcGOhFxqAWefUj/dnaiQtchH6Vh++mYZxSUNDY4
gb1Z1H7xAIMNZrdCgDzih+3jiPWVhOvqIs+OAzhYa++T71F2jjorF7jldZzK/kaQ
5M0VSajplxKhQ1qyPX3W0A+gAI/oYuXerRyocgDazSchHipV1Fijo3R5+7qf/+AF
Z+WZbucig5FepJ5d4DRBZSt60ILpTeecRmtPfqHJEpvOq/1fp9HdLLavv1H001ZY
MRS5fNtk5WAYbUe/IYhJpSpxOKBXxGg/kiiI9lXgqiYCRC8mjNSexO+DVf99rlCU
1eaLcLMLRs5DxwQRsjtBeGzku/SJFBiWy5DXa0Du++rJSFaGLRz60MwhYdvshbAn
i2ezZRTqNao4Z/OKkzWA1jN4vVVttEsAu7A70Almfc2xMjs28e6IVGc8ofWrteZc
w3p+z4pLpjw7MyAE0VBXt5B3D64hBd2PttXr+9a6NJ2WCt05nr56KCLqL3krpkdI
EeBmXK/C4FH6/Y8kl20xUNSAZJoMMdIr1eiaKLaYjgG5pSXBx21n5QB0Vn6QhPDU
zhmdCy5eqny9++Fc1KYG5/hP5RcT2H29Va4FSEWw3mKlVPVYumdSsf9xnGFiNjJ+
vCmzP7ngKhHBaFJl50qconiGg4on2TwY5fhepGoVh4H4uJqW5NP4yNqF09bIyArS
DHkB6NPsy2DI8v9Ozw0WaLrPGythTHKR5dCekCqgrA2rEiGittTpmVZZydPwfsx3
ONfijnpElu3zZi9UjlaTmVzeTjIuU74yhuC6GTURmG/VRB/InEDRWh9YtWysuO7r
vn6+3dcB4hy8gdoz3wkbpC4fzUvtutehuqNQsJwBMFztwAeZVId+8W7koxXklwhC
xEUm+9FIFB0P/nd0PRB8F1jR6JDLhFJuGrxLi5jFtoMVcxsAO32Mr/Yps0US9Of8
o9lEZTw34tHh4F+9OGC2pE81hL6k6U9EcSE/wEcUNHs+mvBrjkAZXXEfIAzdTB1v
b4m9BmqjrgBrq0Txs7KXNK+h3ozN0vnE2fiY82a/k4IYB8ST8+/kzs+W7EHcX/Dx
CMR024CtQmJ607lRbtR93dhd5eRZFR0xcbnHjK3DRRsOP8LhKj4GYWPbZpiR53qf
lTHNPUItaHZpu75DH1Ztv4nKA05y4W3iRUEFQthBWwon2IpW3Nh27q8VaWl9IXk2
bBsay/TiuFRSVYpByaqpNT0bF9xUaaFqUXdIRmcVo4GNf1kXAWZtb3xMQU0Jf0ax
0sASF33KgUOFfSZkHJoAH/MHnJikGRQQoDn7FgvY1WAetDnY3PfDypScIq14iQh+
yOmsi/L5Grdz/GyxQ4L0o+WtYDw51cbS1e/EtD94Yk1ldUX+HRX+8NpZELCy7H5s
yuJiOOSKzCujEL4HadIysUcjFpMtzsD7MbDI3IwhXbFqr2gYxZbzaWobMDEtzGnT
m9x1cWcojkc0mKyZaTsIWwAbOJ8938+8eIqnoD2ByzebwdZTs/8aDh/oNwAxaXr1
SLKSf0ezEyLIp+sjN4v9J30YTFiFb3faINdNid4xcNuSTKjMBB03bSM7b7aisIl7
nB+cU6cwm4KvS+RE0ts16+khLvk6k7H9r8Wm/TU8rNZGamHTz8tK50s7zKr235cp
mYQeB6xu9INbE556a6vk01yBXJMKJGuru97Atgl1e1IZOpeRTydedU1ova6QO1YF
sICxpXsCUSxxlp41jm+p4IWL5Dq8XzC3W+iNYpGJIXVYAO5S3hdoLdvD/kJNvyEb
FrbzpcB/fdfoBP1/fGNya/tmh/9ubOD433laxsbuQ5Nddsp38Hj+Zk29OBhbDbVw
/YLZlpTLMReKP8ge94O0YLy+Gr7gTl2fMv+XszFvPiWciFQjLAoZM+P8/CdcgD5/
uP64SOk2c/1/JS0oMFFCyr6hzHValGmRMCc8HkCAnl42y1yt9q2XwDIyPO/t8wYD
u0ytrifB4IO+OFZ8OxPM0QIAJoFImPmHeOVA3tZPDrdCwJLjE60/atYBIhtEf9xA
D2RvDoRekHarP4e97rT/zvx2LWPLhSQK819hX165gxPFcYa7yS9mmX34NniaPwlL
yEsSsYMHA2GmqqPpvuCUClmrKNKiHGLdrVg9v8eHNndFp+Oy00cxnnOKtYnFaUXl
IT8sM/rL9PWd7jhjXVaDpzlmOC03nzjFs0Qus3smauEag6NzWayHGJMVh75yPnGZ
H2OPZ35S2DKaCxuTkjWgO7RKjt7krLWHgYocnXu7q1cXMS3ZBLnV7Om/V9Y35BRb
D0W+3XoIu64bI3uqsSzJdRCjKJJ7/DeC1HSVba0n4IAQY0/Nn7zFYY7oxMEioBTf
+JBpXvtc6kGd9pZKZ0Ze89cl2oQUvMSG3fbH2gJegnIe/xMgsoS6loJgRQhqWR50
6sLaPgVsn+UH4W9GfrjABmIGVzgL98IoBXgWqKzMZbFC1K7+drlRfipFc+lFFkVw
jVgeqKLmwPfCBbBE6bsN0TLlepPetWzA/WwP6+o8KcekSTcw71hZcLbLMdagJXPk
NnHfr1j4Dgn2FNd+H1IOb9t2AFZtt2K1JgITs8BiZjNbN/pcWNlVjVaUmwjnIrrI
nmJBW2iRPk4fe3IJw19pib0n0lFm00qsNqvdkABMCByAGLDfNTZeT74GKToN0NBh
oJ/X6lPx4ZCzuR3tjRPwLc0bgovxD7guVkYUWh89xh739iEsBMR0tb0FRuGDh1U0
GJGB1epgSshvyYHifmEHTzdL361CyJMWPUN7O8MXtFMVnv5Fn1Vig3W8d3HLPLyj
ypNUGib9V1ITQPcSJ4nAcwMdMZJ0rOB9dw8VgLMtZVt6XR3gyMZ2vfGl8UvAgcgj
i3VUZ8tbDZOPWN6JHS3+5HBOIMGWWlItwv1edaCiPxJDajY8nFGdmGQCrpvcfxpW
xMxQc1GgnUi1IwqOhrU3zEy46ar5OYnvSpb9zKMNYo64sybSM6rjgG7Df6CdAWrC
Vwum175adXysrQsUC4bjdCr5LjfGDHqXZ1/DOZUQyYM2VBuz+/rm2UMt5HSxtdpG
er+3VYBqbkjkP0MVm23ppvJVYhL4wPmBbBmeQ5Ijta4+XFIVmjW2SkOWln03mDjg
VUYvzK0w+F/lcBJAAwl1kE35RxMWwaJDXaJ2+hcUPONcXqjD3wjBxBzFWFaSxoTJ
KQT/S2tR3Y7oZGE9IumU1eB1vZ7bhW1KSaKciQPKYGvsw4Ws85VXCFs34vuLJkTB
Hwt57etFwgSuNRsgB6XfTEcJYRs83q+kPNLF/OpWWFivPo91q+W6qAxAAKcAi9p+
W3cyAimGYZE/AzZRKXf19Qmdj8vV/BYSEp+mkd1kHsHl2hbOeTTetjY91AOTPXfO
pP9BwZ0hiwuOz5K2MTPPZX90S38dC+QY28M2r7HthqNm1CD35GZCGerNslyJUj9h
a6IqtdHI0d56DYogfWmG8l53LiUqAk7WT6b3Ms5DtEj8v6kislKy46IWqlD2ohYt
fl0xg2xaYFUjLauUWhk2D66oquHKzca6qHYjnMamd7+uPS7t/rtu3sjbudu+3tSI
chtmr0eqfZ9n75EV+4zic+CrQEAVy07PfDIF2dZtkcIaMbLridPcd3Nsi8C+jytC
CBGTNNfnAJv+cQd+Twpyc9oQvl787eqsXM0avbQCVBt3p+iAxgPRt1GakqtLksPe
gbYjuCqnIf5wkx2wizMeci/YrKQkFcw9QbKVF5gZUNfZXNrJwNHReYKuCH6OvDO2
7JuxQx9/EmQ7l5f2u50PA6yPbSHgp2b7W51YdXRovXzZpEPjfmfUjkTkfXc2BeGB
5/I94qYRiz3C2HAYtQVrnwf17/4Ic/NseU8FFUElcnVzqbK9tCyr60hH2gda65WW
JfVTjFZL+i0siOSH7maYfjsENzSP9Q/AS+eTNhPiKahg6+WlZcikb5DyNyULrMjt
6fFdmMRCUePqU1UCCrpJ4SGmQOiY1YBWcWRLGfmVbVdUbXJuIyf2WIwLbX2iczct
WvEN6n3v9nexnjeKXX9jqidQ4vl29rhzDxKKi/cw9kJqW5FIfYoltHN+kQgoNd07
BYMJCfhCjWAQQD1oBrlZH9Z4TTPd6qj1M1eHgz+zR9qdN/67DW65utlozLYhBbZh
24+4hkQzN7x8mYTvWjTkR8vsySEKtGiUu1GyUBDTVhYitKsOEDhSP1ACP3zYJ9RK
K+32hm7oAtNW5mAr9Uf3AXL0m6TY1h8axQQLx4EPIMVlKCOCrFE1BRhg71vg8egP
YqNQ8BKIyGkhp4MrEWEGh1iu//RDm/elP8HFmYB2gzO0rG5wIGn4EjuRZrf6npeH
kbUWUIas3EQIiQpfj6ye5L4JcK2AqN7B5dIxjdjXJOW471pYIc8rWoJqlg3j4cvm
ijWTSKmR4IIYpFT0rFMfyF7JhIybVaHVYhk9D1cl/aqO7VhNQOubYOtdsSoxMQRw
IPHJl8MYFrm+knXNYa5hVgd2tzCJ9d/QW6w1wm5XDLB56C15rq6hHpPPV8qhXim7
Jc9Yp2+sYU7EiIwNIsYBZS16Vtwq5EUGOExbEjB6xWqFZ1iW0KwHCnYoREUXp27r
p6/Zdcedny9UbIdfjJUOUJOZKRn0KXeOupf2iNSpejW8jBoO7iw6kVvKUbt+Cf2M
Hgua1BFXJzoPyReznZdx68jlvqD/R1HAFwwWJz5HvVE7cYkk/pol662/WWkoWqmO
Mp70es0ENzMYk/64mxso7i2q1hY6Q8sJ9hyHUxSWm78HFDW8nzD1AdTQBngy3q8q
9/zTYzWO0mnKCgayt63R1Q7p+XYWPphLNhTkyFpy7mumeOtsYvesiERka423pgC3
UE+6kXG8YZSJGeUUgMy8KnWWvYRBKyNFFPHWHY2UNdljMyxaenrUF3J+iLQAtnIG
1iRg9Huw5C2J5zYsUimoYtm7Z7deHF81lejhx7GcvXFNVKz1QPU2Jiu8Ef3D6kqb
cJyDKaPO2SJTlsNUDG6uqR66LluiPGvY+gBAXWLZisYnR2tqU3LjiItgmyXDhQ08
5cy2ObEDvrmc8ZD9HyIxHqRxqZbG1x2vUt38C9PEqmnP/jBAOhU7HunTntPNrBCC
iFNVsBu0+f5Qu08SArYSOajeCIxiK8Ecsx8w3f7Fwf2B1Wljn6TDLLwlghbknsZW
VdgupnTwYZHSFjNA74EpSNeObDHpJ/i11yyFeCKJXqk6EHhSZQh8QwHnvBxkUfZY
xyxX/czeg05NLquSMEBUIKPE7ZzIYVOwPzuXadvPW0NLnqqC5drhQ6EJNkNXvCRi
vOCwipdEWrwpSphc6u50OA34FJgvte6m20SC/1ZsoHsRrrhhzBaQ+9DLgyfTSklC
CAxiytooRn79nVYsH2yRhYw6nVy3jhly/dX9FqloB6lPs+zX2DVpEKvIHx6IhAg7
XQjIAo6LHUay7LZbDv+P1mvYinJdLVdzy82BLWAIaVAlPm6ZWHqcIAqGDU6WwMPt
O7GR3VwNEQoldWFVbePvc1MXs9ZWRv4OQAcQbhY49k5MsD3lgwG4JBYgnIm7xx8j
eTAn91xdht7Keq9Iel379H7D3gG3WnsXk8xUKT5moyvZt/yL4uhWtyeLiWQ8WBHO
cY22hyZglSSeMj3H+BnGUz2QciAO5PhHFwJXZVE5SxOeQ1AES0fxXeAH5AMrWbw/
WhE+U9a3PxpNoJUavR1Jutg9Ks/U4XQYB5QapJQNnjxPW+N6VTC9OJaT5+W0DNB7
Y8hRUOhZz1Rl9mxMXt0/LCkZDgVOgQB3hvveQROOu5Jyt9RIWBCO9NUD2BRgRfkm
vpmnCPr0viOf+eYmZKOlc/1C56eVNfFIMMTreCC8NTjt+um6vIxvxd77uZXaJeUY
mWneccpLCQSABWG6YJiFFpJKY62HQLwlaF0fkHL4aE1e880K+vqTQoTsXsc2FNb+
YiXtzK1G9/sXnwlXnac4IbMjBBtGwb9NAhRh2X/F8iYIgfyl8KlzqDfTDnakPcDZ
TNP5ZbvlvNc9Y3Kk2XYzxgec7CVbPavyiXDwluyZMzBoV8xwLWBJn9ZA9ltUppqd
Z3sAjhBNDMsmRiLCIKwrsz8M1v45HoTc+wQBlozHpm2Yf/lp7vxIBr/YkZO+SkSC
vU0zqc38t2qbbec1mFN/9Dg7gDdERCgUFGkbM4Mj56xkWVFiI3uf8PXTfNtmf7EF
d0p5RVUb7OeJOBtNy5hiiRRCijgCj5WTSkdTbqbZ0xYwcCjOylZyIJ1m2iPGaLsn
r+g8/IWeAYowdXFhnVtpJO8ybwif1KgttfeWA+sk5f8VRBUL4FexSldnQcVVFl/r
kXGMLw/O//cLPM7sCXYkVx+11ELan7LNEs5PSEcUkm2O6W3W+IqmNLHlsiLFXS/j
irFNjVgmVwYQVafu11fV2jMMBX+wyqcrk/iV/9iIt8KCVwfFYmSlwCUrUKSkpQ+i
t2KVnGVulyi/YRHiGmSZ3mmyVC7ckxbsN18DGvVHkt3dVJ65CPQYAn3m59zhIFBI
WS0FKHtbKIvdHisF9iHfLH7iVogrJLWXJnb99wXr1XO5Z+uDacvRtZgEUPFvJFoL
u91HmHInhSmAif140Wsw/RKq7LmZU2zfdSKyPZUOZoQi2uc3WMBklET1yS/LmnAu
gy+cTGVtcS1BuSQnjZp1KDb4ErIuWGLPjRFrgVf/tVUYQoZJJCCBrSHzHnhJpVSN
mDvSnAY/ivLKPRr1YbfRfHMHQlTSteziJHzcVI48o/GyaK0bhHZraZf6outZ9F9L
KVcozKVqmp8eVedjVPkQxP95m+YP9b+K4wO1R2REFgCbsCm3pUvdYiKOfcJ1nRyU
eG2iDF75nnVFqAxK4JW8oFKnklwj4MlJBx0CczfpgX8UqxD2BsZsFxaHUCeIjyIF
udA1LY5s9kE7pZLf7JeIpGWY85ljivlyUuc2d8sdjqGFZGNawfe1WRvHP2l2+yfn
UWKFjj6wU4Ufmn1VnFEZqjtDss2jvjh1sbESxIxjwGKK4qjf+93kU8jcgf6IBqj5
6QVQQmzTNRcJfNvQTMkdF1ql35SrIQuWs+KgH/7LpW5plD00KhRXGC21lGKy3ElT
QL5QsxBRo/QCRCV6C7Hm3RqYyRPbjdGYE+wfR0PekTluplBOkIeXAF1QEFB14md6
Vz45G0kjvBg6JZFzynS/jBR+WIJUOWXxu99a0ibooOcTFlYi6l6WexTbhazibf9b
0fsthHWuxAu8fIlyw0ZGVGxK3sK0JfrP/A1c2PzxYoXQO3gPWRoEijl/xUSTDMJu
fJTtINJhonTbLFakkKUwrySTib3Ez4RAE8R4VDfzDmHQMsBrLVUb9tLPnxG1uRGH
BqezcZvDmGwu27UVk+nCBxqdx6EG72gjEilv+YmhuQiPJKYxKoH3MtHd3ygPx5TR
8jwNRLRgbmOTz/rfviYqdGI3v/Ok4Nf9d9H/vW9ST6CsOLOSc0PDFTejto/qkF4K
hgDXXhgDL+I4QHcIEmQxF26VwrdE3KSgh5qXG/OpeF0FMDOvdAVhCGsb6E7njHOm
r79Pn308gCo5NW/j9C0jK3eMy/zEQOGIYspxtet/4I5bY+gb55f4BE7vN2oEp1bd
tPsUUE9iwabzcyFFLA06D3wNwapzsU+8zM+2obFAH/DCET7B4yUt0wtKbsTqOk1O
4cEMdYWSHVA5YBGhnpMSc18FTgmZrROfqdTRVSFzedBDz7JB8poO1KwSYwoTb2PJ
RnGJpgqi5D6Nj1ryGno7GNvwQSOdJf6aRXTL7WfQKIzgY5CkawHw9LH6HH1E30T/
JrgQWKzuxVqc5s34b2/1Y96AGQX/dCaFdTRPtVy40zow2OFF2sJfgZ4m8P0xGrYW
7Ah/hDeirIaW37GT3kGpYt+bR2jV95lLTIXWDK4CZV1C8If/MziYU4P67CDf7ZgK
ADvS1SQ78Ltyz5/fvX5un/WN8yElmCCtv3zbgMVVBNonlaHzDkJWZKln3afXoObk
lepw5ZluYu74L7G/Im7VvtuhITTG+HJ3c70Zi8umTyeH40Nt/cBD9RIQNjcYcGSQ
a5QT4y0LYR5Ll2OaxndM11rDIgrAg/BV+G0BnxU2yg7Vi0WS5Du9K1Jp7oKPRntV
Eb9r/abvCXfr3kcuTaMXY2MaJ3Mx/87N0uQ6AOX6ARCF5hQGrv0rwUYDM10iq995
ZKtDwL3HNrWzV4upkCmu+8wmnUkllP4OpfyXSpoW5sZ14uIlv1DIpFzsO94pO1QB
K8ZRASSx4OxintaIs3zh9XtpJFoAA90n95T0+khx9iTmlvyXHBKnT7YMphhoEz+S
CVDhI8AbXEDG+/L/RSjhrESHrqh8VmymgYTk5zV1bxXchETuW+WuSXuql5eNW6qE
kawOyiFlTroRicEpegwMU7acGqf0z9kKiePUrKHOZ3zt6jemg/pinz+CVQPOhmB7
ig2x5vSeBzI7HawzL3PQQeqJgz3JorhKkKm7W/EUDUdNpRilNQ8a6BYzwgEQtHrD
1BVXKxML+5qpxckC1ch8znca41fCrJqS3k8h9+Kuxs+0GQMqwHDHIowzPgYNiayM
7IfTveu8pb8ES6js32RcXK4nAC3frR3v7u9aBuaWsmBgiMmTJLW2bIRjAkcW9mVf
ptHqZrozBdV34eojhvNKxbft66lPKTdXnyzDlncYyzm1t66YFw457+d/twvn/Q7Q
Ee77bOZI7Q2row+xkRsVwJAPv/CP/5fYejl7Vl2jon5DQEdy/kHX2z6WHU8GfTTT
qjXZcRjusJs1NTvx9NfK8qBP0RzvG5+B3v1FIcKABNqHYf6sA30zMGa57adFa2EJ
6C3V5MtwCchkPN1Z46nvp0gur+dRjsbsuTCXLvHDm/vyidT3M+xTgKOHjhh1HD2S
Vt9WdRI/CJ1bv07MebHQbsKccxMOCH3uCrKqoxbm2VG39PoKkHNwBvApzZzE1lLG
gK0/yE+6qq5Y34KZJSz3QPGlEKotVlW2pjT7POwvXd+YM6CAO4NtEdc/p52eufAV
zCgjcAUw8Abz+5286J8SBpXQ8cjvTrtQvZeAJZIPlop8q9rtDMG+blhHzMWzc8BL
V+K8IEKd52JOXKuDeae7YTwOsF0xzY4lR7pLa0nEZpHrAmTX2NxqZp4KHgsgXCcH
N4yWDRyWs6tjA1iTlJEUKcj7AZf1IAFK6DEjl420Ct6HHoH04/W/nEva90u6R/ov
uiaDKwGiX0aw7oKjb6dN2hnaEk5WHT5GgvQ56H7hMPwIwA/KA12QScDI8PvpAADj
xkTdrQOWt5Nbwc4N6JQZpFscTDPxHv/ybt4iKTfohDPtnC2aHrubiz5BxhGGxpLl
/SCH+MbLnRgGmnbJQ3A9RLzFwhNTp9wmpdkZJqGm1oQI4/N4t83Or9hi3dEIyHjx
5OtjvpeWPlFJ0pMdlTJupuztdQN7VWGID5DzSfa/6hr0jmRtd20pq2k+P5KVhSXY
vXP2Omu6OYsb76rLcZv/4NXp6APpuWkccgKCs4eCH6cWxUzWQ80680nKZhEu4jJf
TJ+O2FVgBnmG5KdjTaWZGO2sopTWfPwvErMzsfEJ0GjVZJwcjhHG2bHFrwe6vNle
QpWB1LCnwlBWfDQ4j0UbMq/S8xgVe6WgXad4yGtPSdrmdWJzPFLMycKxy2cCbBy3
DYWVQJ5LgVoCNH+htZYAxk3dkmmhWGvoF1W7kr4LgIJg21FJXLTZSWY3V/l2vfHQ
yHeahM7yyb4WG2apMNmJ2zXDvBJdPWIAMOZKjGyAWd1JadoZ92JR7rP4dKoe90Ds
1FfDMNU5NdyymeAlwlgtA7Fc5X0ElImEAO3bI/JcRgz5btBRjNwQoLqzt0xTVgyb
/0EOnGxeBKFraZHAljTx+4e1nVj9iGLfCSNL0R5J+4KGK3DHCL4acKBAO89m+C0A
BCTFMfQnNXNOyisClcBJIWQrk8tFf+OMfnnV+rXw3DTGWlmRb18/+E+QnUhp/Z/5
DcA39JxYQShy0d3Ya/wabiDNh1onnTUQQpwIzSiqw0uP+AXWC7zbYeFnmsdfjI8s
eg/7hCGvY3PY6SCf8uotqFzKGFJLxK6JtBbPfGCxKHWwjHuEn/5EYJUBOUCqFHQd
yWHoig5pVbnPFvCp/G8WNTjApN55vLtuMVUlGVXUUe6qrkBdpOKAuFdSMAYKG9sQ
eyR/Mf0yHRGm/xZ75+pVBbcgChKQuffiiW5zlm9NoC/2Cn0/JHoHcGuYrrnyUkYE
ckYhe6cLHReHNmsqBbMuwFx8f5RKfKwYkzx6fdwv/FjjboiqBxaGKL44QIelnkr1
DKewf/GnzG6D7b+XdznWBUl1PR5iCw9/alPJ7PWCYfvFiqx76ZLyEA/Y8ycIKe4k
SzK6CvgbapVWgIeK/She5uoix0GYQrI9X7I75/rZuZKXw6ZrHI/bFS+rWx8zgKLG
UrU2/pVxaPDwziL5Ey7RnVivQpuiO8l93wCn/PmCcX3WcJbhNWnDlVFU8VWcdxMR
CP1yT9IEs2iddbySI4Xy0iqGyWeEIYrzy4TappV3ixlfEyzCWjNuhZZxGmBvP3In
4uf9JxsId/pKlhxMkPPDOQm/+SDrfrZlovlBZJf/aqX7gz+Gz8aIbBjThRjwbDGR
+5UmA2Ex3k65X3RPvWn1koZfLly+x4syXYLlN713I68bdVhr3SQ0F798Unqv/9Sk
u/rDZiiDkdtuLHeEhNSYhWMhZIi5Hyq+7b2BgiapAkEVj0hE8qYGtJhqCuLDUjR8
szwl0O7F9oQdIyytrbJZzWTJYzmt/fS1r1pcusSpdsBCTLL4gFsHHwoSc2x6aZhT
qEnjshczx7KT7Avuyw/VBVz6oNBzbr32vQjxFZFd+4foA1VYrGrKf1ks8yloIfuO
jWkfBD29H/R/xPhb9tucAaVSTah8xQ08m/2Nk99WDP1S1PIynMF9NxI3Z5XFyPpA
DyLtwZJiC6SgavxvRsXf3ZOZpAqW/dYoHqgotUmMI5n+GX702EsvrquzMmKbts5a
XfuwTn3fS5Yg+O3XKgvs9SaHyeI0bvcoMmxLdddA7FWqJitL75n8x18zcJGqPh2Y
GlBji1U2Fpu3dqYo3QZ0SB7EROebYs6lnPTVwguo/OXWcvskssAVfaG9b/J3zaeg
9i1nQ5dioB6ZhkWu65EcnBkT2wWvOJQcvQk2RrOqOsm1r0852J3mdyZtKXH33We2
RMovnvF4AQM8sx4NwH8zki8q4osp283nXrfyAmynKgDDMgojzLvEh6wdm0TZ6Bvh
hNG8saVwEuGNnmy+FEzYxMSewyzNuQlPQGnQJ8pbDKCyMuBdGfXRgfFbIWWbb0zL
pAMajzfqPZ7XXEA7spmER76pBxGMQtBv+5SWDymvHnCXsG5lCdRnZq6ir/C7HuWK
R5jI4iSV6JCrWkooFcA+G6k38EajdrRKnfZOCwE4N6yL1rzZGHtJJ8USlMMEZMbG
ijoRgfwZUWzBz+4ynOs2LUS+fNwPJ/XKqeEtjr343xckXeVx4Z4yBFIqm8uKocqB
rtZ46Zu9UZYyzcDofzkkiV1wlwoAcZYlPdZ5I/cWLiTrD3ADerY9XUe5DaFqizOB
zdDbF7+MEYw1Ad4VPo1XgfK3ypQeMH+GeMWBMwrkxBtVIeIakcBfBWp4hmVOvahB
zLbHFXZj+i9Q0QHiz0Giouif5eqSmbj2Msn8/EOajyIw/CbBOr1ziAbs/fxkzkoW
YIcb4OITZAbJGPcvMSRibHnE7zaGv7pOqMOPVoxGIx463gzuqQPOLMbViXS6/gCz
fUgPdF4H1zjdTPEhHuTAsxkK+3cHmYoPEanzDK7XCP+FPNPGPgPlY0P7OGzuprOz
wCyn+R1bnD2ZbNNzHLlstLTC9kBgF0DjkpVwgOCiXVLaWzeTmHZdqtiY5kjIP9jF
+yAFdcZkV+kC3JKEOSsQ5FQeF0yeS12x34YW5I0yI+Yfsf2DHogzxXDijqngNWEU
rSibp1qvYCCquqpUL4HmJVik9NYZg0W7uCVRWFx+9zx5fUmJqbwSi0s6NC1+bX4s
ncZ5MaDKXBEmWpTf4K+xAFvSLhBBK6GSwF2tzr2jdJjo0v1LMolauSiqHIL3aMWy
kLCL800XhlUs0biMxYyE+14enX5Ex2UQQ6qQjrMR4fc6sVIXjk5i2tgMh43iOhaT
/vt4Z311hG3d7t45sCeSj5PFUxrp3oyq0ScXXvYWxZAjd77YvsUo1mffyl4CwlAn
c3FtZ5UWhI2s2sy8DFWK7ynwRjSJpaTxJRYpmKAHajkTCFNTr3+5j6eOuDddN+FK
3qFBxBQ/bwg2QANODSAAXeF/5HgmLMjADnIANseSOsIUptY1mjRuL/F9JkA8B0Cm
zcLPE+pzR6WQut7x0SpiEMursAQnd3RIXAIMegG1wNEqWpOxsZDw40COzuvrJzMx
w/VjTW2znK6z+nBC4SVHCtrfv8ypqyJrQpOErH5tdru2xJ43NFUkO0QimtzHRIep
4l6MI1FnRW3ZZez3iD3wdet6YCpAL2GmbFMTy1Ls0cQkCOSNxMVZnyMqaU2Am64q
0TGx/oo5+22CsfRl19JBxkIP53oaJ3FVE/Yqr3iseo39tRDpsBywE9i2G8wnso5K
NEjDM8NZmyWDfopMFwMHJPn5rHt31mYjq7jlBF+FZZgQD3atLj+vCJ13M3fwTN/a
70z2T2pHIexqrgZfpoW+/9FKXT8ikP4WEl7uLC7FfL0C9FCxmEU8Wnu5Q0frZ0sv
DcEx3pWuTgfyqqd8PXG1YLcprCy4zvJMbamMs7WWtXDW2yMvL1L2Z3Z8kXvOrkbV
w78Yfem1GNTXuEklB2JAufChS595zt824N97au9XJ/PJ9OPcHrFQgBAieoIXJX4S
RcGabqWT0lFBkYmvP3IziWzq1dyvQOFmP2siVpJd6DXg0jqf948b2ZV4xH0m0LXF
oZc58i2PmxcdenEimgAXc8G2kkhju1No03aqMbVNIMR6kCzAsZnaaUbhr+B8RPfm
Ee6bi1/1C09XEV/HkclQRJUrPc3igxmyb4S9Up3+eTyc+s/y6s4DEOlTinuDTHP1
9Ya/Fjg6mHI5CBnvlf/n2LWbpEvRWCdfcJJXC5JGZ4dnWELrBY1Ov3YFg83aZoT0
yfVr5EAh2k8taONcBl40SBAxbnfw7O725e4h8Ax9DZbxdZqB04M0uVrqDyV123dD
7jW//QtIpVJ7JoidtIrXm/NVs+iYuE0cj4uvYUDWi6sqKXYFbA81oTfwLbyS10/c
bQcl3tWLC44XSoLCSVRpF73yP4zsXsA3XXsb5iOsTEqodfcr4qr/xhQcvrzh5Scx
n3gB7gAzSZy69HgyfvxN0ICjvzCqzOhnb1woio/7nljHedcMRSzCxTV1RT+9Vg8K
K8S/mvTZpb4ClxmgzJGQbJD+LDPqR5hm93kP7YkcfxJ6BAmQEyYdJmusEudIrCt8
1IIoddnEh9p6BCLgB1ew4WrVPm55jwn3Ljl7zdDgxmd6YScraqOOQhmlk+xkrOaa
PuqNckjpG+WnKxEB+IlneQmF/t1NKK/7T5LKJmgXNqkZLBTZTqusOaTJvcd7Hur4
zloMVSb4D0RDet1Tr2RRVTuE+uWWDJXY9rDs08iFyRVD/a/7psj/ZBqm9ZQJGc22
jCN90J5NBFn5JS666e3eqJIdgcKqtJBHuCqezVvl7hBxHd1gsGT3sbbiy7lI93Nb
iud6S17Vz/KZ/S5FcifWBvKH0umKjYEb93/eDVtn8SJnyenNOgsb4Zi9nWZaHHD4
XDGs81ZVzlTGmO5voiRVnvZcig/FEwPaJ08STS+pFADCYKI5JZXdPYLoBDcj8zXv
0uyBIlqvNWOp3ZZhReJDIv/bJaiyZin7ckLkybSiDEbofdfKxMCySRZLMzLF+eFg
VXDddRomvuiM3V3yWxdDSXDCciLJQmrgGuxESJNnT49kApR2CGXwCtV+pZsPaj4G
IUSq3DOnb2LlHAtlNvQEALBYZFN39v54gkDUWcPmccbvMKR+E0CN1176sHWMdPCp
nVpfUk3iuwY9M559HCZqzlNIKN+CdA6/aXUo4qOliGKXmT5nxMzukoMjMJd2CWzU
+R5lXZTeqdUHxuHw7JTX1Vc6O3O57qzrztUhaETVEVWlawz9x/CiF3J1N7aSgLO6
abm9QR3KRJZgdn5v1p0pOClbq+ChXDqnKKtcurtf9TQlDfKCeS0Qss8tyqswXqcW
R96BDJqFby5VOOzdxcPnvch6MKMeMHLqsO+Ozr516gu0Qq0DAxCmMb4YVa1qSSM9
KJjwaTisYBFkbP2iXtWX0Mz5RdO//vCOanMTmz4T5NikWf7gGTk6SP7uaMygjc72
heZh+qktSL54xJusQon/QvNu2fKAXVZflEtT92yuvANzzTu2G3lmx+mogLM7BBZr
noW07HUYCoxjA/Xu9KHK4uFy5wFaD9/plRIGyZqNoXLkLacUxfaq5cIeHjjbLf04
oW/uvxJyeSGCJ4Clhr2aqF1G5vk5MJHJTafVcP6beEiKpl1POEqGmxA1UyTK1ovV
w9ccTm0nDPkfkp7bsg5Lav461P2taqATqiZAMw42GYwEW7Zh+uAdyX6rwRFnd2w7
iZYITRQf0SC10m3dZmOdaVfaw5ounfPKat1ZdkehwAshRZM5d+G/Pa0WBNT3vT+v
sujAcygAKUPPNe4+EdsNAIK/rKx9LrziwPLwd5NsfJoJFFmaetzMPz5pwAAmt1Rm
b+5IUf5uTlISGP6sQvcBJDbwqiMI6susO98QoDtgL6YjMtxH5P8puKOk8dWBO9Ke
OTec00f+fgiKeTSkNrjUz5PCvWSvHrjFDpFbDbGtRur4mYvyAcUZHBLwA4LnOBgW
osB1BuihFHFiyCeyknBwRY8zWWpPeiYZqqDDo0jrvpKrDIK2qf1ez3OdPjNhtgyj
C4FxD5vwlTcf5cbkURvn+H4I1kODwLFWS5cxax1jDE53LoBCpZM3cjdYieOIheaK
B30tutasBq1Gx7uffhXabOTm42QToIzY34btiNvFQavQBJLxg+inRawxDvbBLL6l
N4BhzsOks7dAsnXHNHU1dqsfnKiAbzdnF3qwFP5zd2TVwStwRCRYv1WO/IqfAyW2
2KlmZHjyGCo9i3Vc0iOvj+ar3/TMmPGFQPZj0KyJT76XdDNUveMIO81KIKUAWewr
vSnGiTRkMePe9FfDxsv5bvgpenUlL/MNn5CNThwACglNbW/qpGBpFN35aVBhj5xZ
ffsFFN4cugIYc6Oh5CsefayeToPX8Z+/mq/bSxHCmvQa1YaoLD8CLevP/q9KbnS2
xcFd7Z9+YjbiO9hUtFekV6eSKP6+Dt9SMsaGKrmBCpdrWqoBUClBtNsLt2qIl3GH
/tEMq1eLhMGvvlU80b8LyLjc4uCHhJ9f8KbNrfudF2offtL000Bw5SG77feG00/l
SrdzypDrrrUOxi7XwM6hwM6Z1xjP3347rhBtjYEQg7SBaY/wcJOJ6KTgrv9O9B/2
ZM3pDc9jd6ySl7B/3yuIXEnzxkwjiwZaxAfq/BgV5AaJ6gTkaJnLiPQD2f/Rh1o6
RdAikulumA/SNALmqV35r2ES93mGePoSMyN83CXq2EDGfdzaOxOla6v9pySEfjzz
8xYKbToTzGflLEDKr1QEBn7PqpRiTm9bpMZMqyj8p0ic5AJeRSQLwY4wyUkdQOb/
Tsp/X5fnQSCVY9Uf1dk14SbVBMAF9sFUWoFMQwxrDT0a90g67GifsLEy9s3bUKBo
TZXYi05H6IvyhEwquRAStAFr96J2hyJXWlqzdIJcLlmKBvWx4hQ6j/wGzwwV1nga
oji+4+2vaMTvWfURwmV+kq4S04it8pWRKuSZfMUJaNzEid8EMzMzJXji8sH85Xwg
rnW+htseRX1rUXooENvXlyMo4LD8HLyUxQSmKUYrdTm5kezUI6aDCpWpJZYL7ltQ
zyxaGD9e9pRJlg/w8wA2gj3yWM4Kg7nxQYlQKnWZtqVeGrPpZV0szkcPaKk79Svt
vEkaolKLq5f/IbimtYOYMvW03Q9+t7P0bU5VTfueUR/07HKp//SKBfgHKnB2gAcz
hQ5pbUagSlWM6qPml6hWUTDumL53yWuczHulbixTv8YaRyDGPI1aldhR08B384ff
QZE7KTI+CadkZqW41txoO1PB40jxXpgKk6Y+wiIu/Uk5pSakavioqp/LvZdmVfcN
aXLngFJLnAii2rqf65crdHgUqfygFNZ2eDshvW3RPYYPIf6vDKH1YMHnTn9dmcNm
qzrvYTZwDXdsrHDsiS8ciGJBydPuiqpl8Urvey+Wk4QJM7QUldrenh4mKhbL6NYZ
RtgN1h2imVtkmmTyWb+9cBvwlaMgCNy0S8hlBhecvfTqJTVqArc0BCtvsy9TgiAz
MGCr6ANlDkgOsJOVJGwvvf5l2H0qmCagSYxVxnozVTBpPD4U5/HWephIjGMPritr
Rhi6tLIXim93nvZ0VxD2X4BaD+hcwnNRX67mgeFlI40g7dEOtKwyZI9LR3Xlm3cx
j40e/4NxWIGLJcQ2me73mI3mCC5A2MlhNvTrpyw47l4Jz03SS+/JuGf1rWRQ1x8x
EeQQVhHAqm+mSaDsy8LVFXgMr4oAEQ3c89dJS/PUfgtB1293vtL82s2rurUaM87f
P0vZ72psmnGK15AGa+kypYpoKLEiVmOpLb5RknsSAKDTkdv22NOkVUEgAOFzC1YS
L2b1tz3d5Of5OcA7DBn+B/2TJBEaiW87VW6jSqrywlIn9KK/6zWaMOkWyiFFmjJ6
45Iy4zKRriUc4h4aq7nmCyXJkWbbUiwCB+cpUdveBeg+HupwAy8loPzIzdcVkcWE
ADAjmW4DOw1Rlg7Nm5sQfNVDZQWHCREkufnX3LA+Rbvieq9OAr/82MUurd2I1Vmd
tcL+0LYEiiNuULSgPmvGXBRVNY/sHExH6kaXF9p4cbMl+Dkr6fH1n49YlMwqZzd2
AouVZ2NlM0iEwb/YVUSsRHO/AYL+JL5VUaIey6j85S60Zd/PMNT0nKcpnQyoEvXv
4KvxKIQgFSENluJzhg1n4yU6NxNEbhQRpiGY7mCJSqPOdQVnxcIgMel0jAQ3Bb/2
CNUqFL++heCti7sADdAKVf40b/RxHxhVzwjH0eLvUPk+uw6/QZxKaWHY4kwxflqV
AVlo75cXZQMbkpbRaXTTgXn/NOzW7pC8YBGPGsqUuofGA2ipZZZRRB8/nbChwcef
l9g452IO7/nv4eTEVAo8zR/Ro0Q6IilAYNZo4zsX9Kcg1y5pdbLbEtWApsoup698
dyBm6YTgSzmhZ0F2gii2d6drm3v0kYXLRhty7nRe5pnmZLKtd+qpoT9TCgLwZRb8
1SVcEXiY3JlRJqWvswMwj4B5B/7WBnFbZmnOVpHV21taEr1uK5mkUQp0T1Wl+y5H
dc321sd7b9X3686kl2Gkhk2QGiA+RDwx44r9wBh6oVQDeTYq+0mljEdW2yY0rXuN
SXl2DY/q9aLWmAHw9PFHM6e2rwZ0q/xs8XacSq70UaWjVaqUiX/t7Up4rS02Z41k
kzHjO+iBar9SzCtG4AYs2Z+XFkZdg7na94lwPGO8m6G9FnTWmvgPUJUmohCvt8PN
EqSFAP6nk6RBAGBE4PjONurz3/wySXbMNwjgAGrBAjNbeD5ZaEHG2UlglbIlhqqG
qZKvtqwhtOuqr+uaxBMWkaOWZJGWMyUGiSMFbpxoUHwIl/6JLy7UUCFZjf+tb/MO
Df5PILrn95murrNbWqPJBO/Wm6flGjEaYkABGDHBEw70k/IQtdA13Wdf+M8P6wgd
4llxjnaAfEgfmnEm/s7UtZJ3iApHio5YwqVx6NxjYYWuaS4OVNYHJ1GYxEPNyqpS
Q3W0KUsQ3OBUhpDYxZmIPOlY8lkLoh3jk4xTIC40V+wvGjZexBOsvdwv1mkov05g
/RUrRS3yeHE4ugCh8+6v74STEIxkGFEwsLz+a9RVxkpuIEFCWTgs5F/7/AlT4Tim
LSV4DeFRLEVaiquhlXBhq1l0F45c1bAkYw54Y7mc2Xlj9HVYw1Sq5YqDbFXsTk4Z
gzpS/0RKa3XqqB3rJjCaQkkr1yUyq7unkiUZbEkqNdLX7nuNrdUC3H9vJqkcxq9C
ZCkfX9sOz5vW5SQkuI5A/LG/bHX0sSuze9WTDVjbLxgp8ED1gNlHFaW1RoDyG7bs
kikNVQXy+pgXXCo3guqKD3bszt2kci4UXEQEfLZ34GRKMViUO66TTG5p6IG2acXp
bv/ya02K1R9k1NYwbJ7MY6O/Cp41VMbrGDIYIGLzlx2b3AY8rvnrbWOSsIKMnYXF
pNQQR/AGlyQu7ZhjsMzSNfz08tPUrbI8xJtUwoqrv7Y5ibT9da8ISavZGJbdo3Un
irdWlPa62EpFOIRl2ec5YRZsbrx2rrrVQOB55zmcHfeUDIW7CvaC85oPAnRX9ySt
Yzw7spDtQDVVjWAZ7o3NPyBT22CuZUCTIm6mOXzgnruY8Tr2XpItppbWerZPWB2K
3brYX/j8NW3IjevB+1G5bS4w5xnZOSQbQRiR1FSayhVRdEz1p8NWyXaCUkZgBEEK
xpDSbe3uJ7Fnf+NQuvl4kxui46RJ9YidYvU0OKhw4uIwxwVY4My1FGG/S1OgwHq2
XWu7ant+vWRwOQ6bk+viY2p+O24IV3mR9xIdiWkUcHJsv2yd3Rd+bbcM2wiIfIVX
7x3vpGt+OH3cbXmAiJmFHJLIZqfVT3PcK7TH4HKyTqzxYSuK+cgw20zK2+gZydnf
v+B3/qnTkW1uIditGQ29xy9Zo+DELmmIegPT8Wgb4QJPVCnHivcW87CPtY/yggLJ
vTAWXUtTk+0alIMFzkq92dvfDRICaiDDj8RpfVBq36dqCa23Sed7abtOO401PM5Z
zqAB9vgvISBYX375bWQ9XZTDLwUE3hKuNPKXlCmox4DHBGcPqoKHVpqMY3G4d4x4
j52jN9ShSL5AKJondf5A0X4TKwMpRQMjZ07ejr+yJiajMPeAVGn6S3+26v96uPn5
ZEnv9JQbNxb1GXOlhvYXljWMskBTbi2N+fu5AqFfxmt35pPLYY2jXE+r03ATimd8
WKPFe5cdW5Px3kZFZEu3Yghv4JxY89mgY3Jhd4670iE5NLkdQKx2jH7M6NT9e82f
bpRa9vxcbvMvzbCV3htnLac5zbridRzxRjA/DTBFptGnvqDPJlf1SMODv4XefoRA
wFZ6W96EBxKdPxJt6E5Gy+u6DCm3z9NJbXxoorl/fJGj4L0SUj3HXCPdYXuZtthR
Da279d0/2JeIfq4kkB4eam+hYoIoLXqlsipGDxilAQh/YSOffNnwROAIPuZJxXXw
izG6XIYBe9fBLWDn8/KyS9oDE9rL+k8ok41vjbY3XRc4oPCC+8p0idx4RIBPIjET
PXNFmbhVhvWFO6/3mCOH8/Gs+3qlvVBLZpoQilGRBgBGRYc0Ws/b5tftvNbjtmkY
7yVvu8MtjxYwButIGCKPbLOz910nIb14EJ2fUxFogECdfirg8UAAvLeRX701DlxP
dsKRdN9HBTPYNYy8jZwrONYPDALPJoKJxRREPHai9H2mlJkNYEbDDGp5SVMVmqza
ktmxIeh7xO1j8x2zHzL7SP6mfidHTpjFqXF3dzd1cRXOc7IDcArL+QXtQy9Nrrbt
DKurtyE2JBDxZPMhIZovhjZD4N6xZE7czj/tZgvgoBqOJU7neE/ZLa3a6d/jf8/F
sRZMSTUcuy1nUxoFmYFWkajz8dTF9JWEUBRIygn0qLw5XySJ2WJcytOFhtYPMxtC
WRPOV2R2AAJZdM3YLM2Vscyn7xONvXH4i/FvCKRxsuRDdW7lv6Dsbbm1vP8cdv7k
tqrdMFhVj7eRMetaacd+rBEwTIM34k51L/ZwwrfVGlE/Xtss5FSAas/YBOvlelIO
PXIWS6OfmOiRGJZkzW08vh/eSgAVLB8YGKCEZi7W9bFtmvADrRzFkfZR3ti48lAY
PvwfyvRPcWxWpooToNFBGtuSeXIOoIBe6P08e2sQaKwh6NVBW3PjRXosn/6XiJr4
CPzYoi8XJ0idx3sYfF3QXteRtlYNAfB9Z851ye3oOcBYJEjMPnSxDMaMDGtoq1qR
XBO1ifkXrbInxSzeMgdZM1Bi+4qa7RVo9z5YvCoOYff5oAUFBg8UR/uU6yRoc5l8
LB8hpphyLnYKdIOYhcLzGuoYltlxFaerC/Gs8mg9+mM4xqATXwVpQnj7iqKrhzCJ
8JCNu9Nj+LLBXBWKg0BB/uBYRFu5/ejNEq+E1MuSuEZpb+pya7pqImf2tremQHjE
tcpn/EqLdFaq9gD7060Q9bqBgmFqqD/ZcEaH5UWl3MiMKQbX6O+bJm0xnL3Xc9AP
OBUlcEYZ0KKn3AGYdBCAxuvuMbV+rlTk/++jy0Brp0ATVZzRwJ9PVCXPds5Wl+WF
qwUiDP8P3eXv5+voUf01SUfXhBxCsItsPTvq/cwcJWCgae2RAAx21vxVWoFeYbb2
V/GJHlIvkEV4ALYy0tonkH8wm65bFuxWkSgckgN8SYlOVpMZ+gemrH0+3jwWEag+
NaVqnJlRa/I+ubUl3Mms+Y8w8sMZBnO292VVIzqd3RXQ4jrWeTmQXwnq4rg98O0o
pSk/a+K+n1AgJ1pNrfnSnJgtf3HXp/t4qxZHkx3IAkFvDkTPByq3ALiF9cZE5qtO
ryGSNNOpdggdXH22Tyrffqnc9hqBdf2SA/pce97ouLCfOagVGtvuAjXHHbSwh/ei
wX7t99Wk+u6uAK9pPe+T+iTVRCipCBrYW8tRzqToEFX8Y2/JRseUXwH2BuIekrvG
B/vK9GZA2lw2Sood5WsLQxR5UBBVnna//hbVtv3VfvDhTKnHzht2Vgcd9t4ySk8m
+RbYWZdAfmCczFwRJ5lO/uzuvNv8RL38/2SgKtdPRFZP9P3CV527xq+s2n180cVz
FbXQM6BEfT8ftAm2tSHIMtZPbCb7gmVc/No+XjSFF4T8RotlVlh+kFKLphcQzEU3
w7Lz0QpCb8/qD4MkDimuY4WjxRWcNk4kWaZ58K9openh0M3Q3tbB/Di70Hc5lt3X
F5qhtehct22dj/nAW6oDT4QRmLLU89u1rEE8hZSW6Zy04/WxQJTF5H/g644jR7R3
YRmo2oKiPwWJ6WfR4DxtezPvEVkasfgf62RpnMbLbvwu9Zkqzd0iv6UEzI66Z7Ab
P/sruNP7XRDG1X8uCSuQ2dGNdjt5zgUFj9mfFv8dsl0VFxY2o2LssBD8QGFqJJ8H
XThIM8RH6PnoCzcxqAWiGZya+3M/tug21c/rRdzVvMAzLLTMaX84AhEFfN8WKKkP
IM9pNMi0pgDOzH5r75sNVBil6Ej4Ff8qprWsrRhD6GFn9+JLB6e7CxWYxu0PT98r
fbbJlu5SEj+dD2tZUiwV1kEtRN/fgTYEXHNvkf5TgjKlJVMZ2HPSLrXC9cJeGCXE
DRxAVHerK9Y4GoyHX4kMZiY7CVwiIeY5cV29/xscy+9Ucyc1aWt+BCVA8EvXR0qB
D2Jx1nP8eS91+k7LiyKePCOiaAc7ZUHbS36QlnSFnGoKeisGfZ1Gp8pd5tZJRlE+
zp0rThEFqtQpMPnxT97wz1BgHX/aRMXHSW5DJiq+Y55dgukDx0rMzMldcqtyuFFe
BToa13+Uxfnszfyvl8PZC8l1KO3cbY5sE3BDfg4tdb4bWoa0YPEq9xceaKzcyXk7
A0iJht24HBXLOKny7w/tflVMtGbAuLVpnNDp5Oz852hnpPoWDIboxFY48VubV+rJ
uxOeAhfdqvGo3qivUwTlMosNoqDfIXw1fuc77lv0XiYLrcyzchqAP8+SY/xi1wBv
GybRIqj2S62M4r7feJsbu1rWWrt366hbZChaXayneQPrbCceDcWKbuF5lxMrxt3B
vACupJuKbXWJrFj68+AO3eBKFZEQ4/jD6D5snHolmFc1He+DeoHkzzhfOFH42YB7
5dw0ElT7zbr2912rsthjIMDsdrCUKYc1QM2TainZ0Yhz4VZDZzvhzWXbVNLA8I9t
I7W3Cx3/XE7xZwsvNbJnTkFQ8HFQSkOGq+JMR7aq4NsXC9eGPw7u+YttACcjgHPB
qeNs+0t4Yn6hEsvM64tqxumhr8gLn51HpvqzE2N+LSRj9o9T/lOpXuuKMCONmdVJ
JkkwRuzwTVYIr49rRzLdJ81gf5Z4cPtEvKgu3dqNVIgjDocr7q+hPw07Jec5Uq32
bxvHl4b0AJkOEqYvB8n7OUN0pVoPUHmrjr4KX2d4Xxz7l0IyNHYt2umUeudp9SqH
eqqwRSLwbjcDYEGEdk2Tnpwu/jJfWCIH+ghZhSq+bvQBRdcXYtDc+WfSfpkiBLYd
5Rp5VhtU/zsUcoz6ckQXTOu6GskQvud2Ud03KvPREckvpGJAe9dE7bD5sLjbt/Q5
pcnEyTVvBaUv2aIBAUrbaXbmwY8bM0JK67MPwxCX0h1F3XJ7ZBDR6u9vWAfi3NrV
FLtfEtHkooLt2O2ECEAMJn/RgUFeecrbRYwg1kr7C1VwGQmB5eCrbkhRqtOPepJA
lS/Z0seULefTfDV6587kt3/zT9oUWUmjXZinScjgVv4iFCljEuq0YgQ2V3zDLGKa
htz0SWoc5FElOqSDALiASUOIZbjWAenFlcwfGQlpjF8oh4c6vPikUhIJk5iPz7YD
NdB2gPTGUHhZP3P50fqAWd7cBWV0SmIQNm6v8toy88CwM/SceN44etpbTJyC1Dt5
d9ZS858VWWmLL38iqPnt6q4N9PT8otCgGVY2gw9egmBrC8LDAbUdcbqH8n2v+ui/
JS2lM3JJu8B8ZYdAtuepy1JhZu0Py9xXPvIHc4AYrtpvfx1CzL0MMqD9VfmMTI/u
AYlSgNwK/e5V/CYtlvNPMrm3+ZawhDaRpQ0vOOODQCR3+MMZdTBIBR2Bir3Uurr5
PyZSB7al03ytpEXWJ7q+r+9Dxar+iC50rasmGmqlEEvOd2V9MdJV6tgdqT3tZgJU
2DOFSf+f2/0pKGS2Apsdq5RgRR0NTksPUq+yIcmnNMkKjzYMrBza7W+AjaQCkZtD
W+6n5S6imDYqNBhyAtRdozK9Vv7btnAsnJacWckEM2NBhmd0XmNlvJKoaw6P/qAb
len8D46ulNRGSGN33d3Yl/E8+rOoXGhwvgdL6xULGXfDj7A59UESS3gyN4o6dF7L
xETsAGSXr91U8dUF6z+hamb1YZAqdGqzHef4FHP0zmwFppfcdBkp/8ywc6Xz+7BL
gpwPLBhM0UsMvEsmrexyzkLr4NTg7yCi9ersWzkNlHCq9XYTn2rXIwE8rR1KGOU4
pFFlpG6wVvTiS+Hjg7ZfIsBU9RloNbOQ0jL03bAFr4aBNxHTUoq7D8Nqxm+/ycbl
7r9HtQ3jd15MGazEksU6Mzi0XAl2cgHpDesehRES5XcUXxPRWdH+oaoF/to51yXq
JdiOKFAr/KxOSurCXQjkJF7L2NjbBdhx1e1veUoIoF7WBqG683EEcclkM1EmmwHM
/aZf0FzpXrz6HBsiN6ER8DhHONnccKgT0l0xQUklzaSDD9eyhnGxcxtHC9isgU6Q
3AO0/RZ0oyZtO8kxYkz8qyXicCmpVoGBZnhW93siRSwrRJU3Z+Qt1OM3UUUulhJX
SO9NNT9cC16HSx8f/Yhy3kIlHKJbL8KFmQux6Aga2cSm0fJELKFKBGu3B5wP/Bp/
5vXb7PvNgC3uYC1IkQEpoh5qqRnwORK+CTkgeTCdhgeTK2R+5jxg7TXr49ysMR6i
CM5VpL4fNqfjdRpf9Z8yVUC1tx4bWTtob3oy7QDW7oS9VsTS3ctajgXjY4cJZ56g
b0I+ZUhZ+26EmGgs5TamlH3oyTZDC65RoFsptCuPpwAvz3a3tup1tqHte9jsUwtv
AS54lXvAo9ZMiMmUA3xJE2Of6LmBIg3Ijne8L+tv0Ay3WEKDVeFPlexlYx6Av1iV
U6ejCF5ZEWTID7i7WKGS/C2GDA7g+Oyk2fdaLRoEWK4s7mEdFGl4jEIVW2HV74j4
p1tJ+3sVT7mAO+MoEysZz9aRBv9Bk3eQgRuyxeOM6bvmzCpZVvYhlSbnicHmYb0+
Fj6naF9znGful3U80tF1f3rBa6+GNClYGkxNy+OofTg/eogC0dtlmx801w64Eb1M
1Ps2xaTGAAIYVJ5XKxGAODs8JNLvgC+Ha1b8tdzxsNNBE+RNCfMFjxNQshZ1zZko
MNhp9ny6Bzhp1P9+9o4AEMT2K24hQw/coDWbOVUs/aRmef4ItQj9UsljjJNZHRMu
yvaLJW74KVyv0SEA6J7LlhU3pm9oGrgM2Rm2bkIhzzw/WKvLKAkYnjm96PIm8d6j
GP8EPp8k+QBTmkn+pgFDT267YZnMSyZ/hR0j6AeLWAi6cS1gY8GnEzKxP3atXXgw
CdwZyoeQzCRojWjksVg27MrFpkhOBUIjoK+CfekVIK98RT6cBeKu3Npq3X7sjk2L
PkQa2npZW0yRQDH9/xb9R6MRcQOKdopJkwmFrKT4fcp1zFgaHn9FqeA3iOK8nhEY
2DCOsxUug8gFggxv5uhm7p0XP7sg/WXtnbVn2RHAdLG6fsURTfCmI1ZKY4P8S0go
QnR2Eggo67UYG/i6oN6mfY4eY0JdoKOtPkVwaYEX0Iy5BGNZB2Km/ff2uw1xqreY
jon2I1VTCPzpRI1xzK3atLWMvSPsEQwoWOZZByxLmPwqdK+h86+1HLo4RKBBTJpP
L+/vk0UqaAnLhMNrBwGZfhp5enLDFP9LYSab8phyauyoYnSF/FFHl+i5upEbPjjv
hYLcygJc7M64fwZHjZroNGka/wL6xqWMwZkb3kYTyDFlqpx+vUIl0GywkuWnAjb7
+lM/UQIX/gT7WPEmn/zrhrjRUQqiuTMPqeT1zwXK4PquBmdoQPTxdD5M3/29/HDn
3SUAjLJiO/RR+WPWZQA8i5bqLXH8ztQlFziaH0CACK3LMwi2NQe+ncjL1CajA4mE
j3EWv1MeqDSedWpFmohkYdveWlcBpgqsRWr+2npTISZT8M2x094Y7ZiwoTH+Cuuf
zzzpqIRy3nd71UCXhJoSCGvwf4diuEdMqIoonlHW87MeG2oOk/j1Ao8W4L8Jv1tl
zf/mn8RAk6mbzUweZKegSayrulUdkYnoxFx8zFO/ka+ilS9VFCZTPOP9y98rls6h
by7kNd1TY5r4mTaYpj6ySiD8gVonEBpYNBA3QRo6FszBJT4sm/4rrzzI8n3Efpdt
jpe/HlIbsFk7EDMZCLQZrHdza6M6UoRXhQJmY7i9Jj7WSj3+Dq89m/gIfG05Hw22
2bFlaLDl80Q1S/aktKRVTyvKWj1DPR6xD3Jh/KbbVIjfXNqDqPfztDkJZfMVD5Ot
cVvyzSTi5/qoxzyUM6qWUTYfpHSWJRmV6wqYtDwPgVfDdHQcCE7W9kuq0CAYmqiL
GV03J7OylH1px16i7foEUxLl+lPF5vhaoV8c+pGj+fNkh+k5jd9zdWC7WqXoWDfR
G0b5/hGcNkf7Hr9Rw89mGTWOSln8PixyyCnT3ig1bsG+IHKDl1DaBaSBR7465ybL
+GpZCYGTBJA3XH35tLjwFqchy79ojiVU4HmQOIJ7GMzspnzvfsK+WHmEOZTcpX5u
A+of0XEft1+NdppQHGTtqQjDYcW2BS+cbOrSBPcUpt7hf8dVezVO89367JF0E5km
QuPaTdPauc6cqgx/Mu+0gEzI84z0/8oRTuy0Rnqz74xnwPSzZlidMHDpGCjxAlK3
5hngqpkDGNKNXZeBbq01oSm2nQ5cyLEkWesDAXPFvsxZ4Gq2SbF0nvE77uz9m57t
Aeo9a3gLBHYpi5Lk4S/SwcRyXoirKlYkyIYSvkNB2PIO/o2DNUDlf24zObkghUA2
pCKra8cxTalzUqAsePdJD2xAlFuIMJHW/FnXM2HD8/bqDsZngCQtqEwNReAgvtP3
iiAWLlhC72bOaTcz8QgAnt6fYIxn5oXYOKKANn5fYmTxRNp8OB44ZU7CZfgledAT
TyqWjyU60aL4qOjB9aegWaP5SnzGqg1TvpTtQwv6A8GoG7oc8XHQZjfAdZX8zjgp
Rlr24ljnxxNEYC0GCaIbifBB1nNLWTT7q3NKl+ATBk+/LxUWkIP64TBzrbEm5DEQ
ottiIKDhgS0Lgb3/tRLjLjrU8sZ1zH+591vFExW4dpASqwFn3RAKKOTYMocbigna
aKAxj+zSdzrpn4zYvM5cM6ShD1ludAfMjZI9ELTmsjHFRzbxdvbXHhKiS0U3yCM6
WDtKfXFwPrX3orTuGv92LHu77w9DonvxwjCLEb0HbE2ClwKT4mMu1nwlga2reKZw
ood69s30/BL1GeTMEol6JvzQt8bwxB46YvRbf0/ELYfD66hTfcNycwgi4Ge6bAV6
ykndxTlZSrQeIkq1hhGDTcTERXF6XE1yDrmLtX912vqLtiDD10+jQGJrYG6GXCl1
u0gePp+GtEOvwfb8aGA7LOw3e3f2W7hMdoWtCjebN7CkBgut3lzi/b4xRWyyt/sp
zBhPBAU8mFAfeJC9LGkphoCldgbkfsnX2tdJJILOoKHpTC1CEvfTbAMuc7Rc6O5y
Zv94s277whP7Gm3grJ3Gw2JN3CKVqGTQwG5jEtSrbAreKNHvWWumRkBig9Ixy2G+
WWeeCO2PbBSp/dl3rMo+sj8gns7k8pofQ7tfULF3Xj8PRRFDs1qecRrfwxfvE9We
NMbhRHizzMQO9UHpb6aGdnbCFgmImIVPae0JS7vcZLQF9Gb7kv0EZQZm+eL2PA+m
VZMJVI63Xx6yELH1nG0cDKMoIj1Cl5lKUna468FSuSf6WZPloZVJbqXwD8Xc4dNZ
Q/3qiHRRIxEziuaCxkYHYbTfBgr1nFGVUp46BWJExK9oUbX62jDXuZQzWfvuRf5p
U115oC9h8qwKEVkKKNdS7dYkhS+wQT9C0o6xHbs7qq5XEfdXwUF/ZwK1pospZtp3
/pz7/y52rfn89flfjslFqP7Uu7cco1afkPiNsQpHu2dy+77l0de6dsiDe549HdXk
KlGAiRDFQ3pZNtyhTwPhaNtK3F1fkxSvZZiQAobjfxDYTQBy1aFSGTQldqqEhKpx
yOY3z/xkZ8BjK0boIqL5vqyol/VXI+flZ+2wjupIWJ5jwkf7BUZptVYVwdf0KCjZ
qMWAQ/zy9L895tBwNItDI9o1JJCZxV5UwTMMoMVFMDMx90lRt1FzUkmNT2q+SK43
yyyNd97p/89Q/aLWcsQq4OHwipe+7khCcZOArABlbqJrZgy2751hOhdoDGskihfH
yEgPTUY3Xmf3sW3tR0mOADsL3fpGbKtqdm/bNeP7YLhFIPlwpQuWPt723Gx6AzH2
2lYVidrbW14M3wLB+1HW3ZYULQgEDJd3f2qxhTgdMKuUphHiG4iCV8kAm46oNy6C
oiEuJYnZtqUmCz/PLyiJW2zfT15m8FTZZs0mUowt7gbH4D4yC12QlAbwbYkP6aNM
BcuBbYEJONR50Jh3J8n6cyzGGk++9lsBkCDIU7PLTya9SRaTgo4SU1UuzXsuhy6c
gL1fiXqxUwAIlmKH1BIBYbDNV2hLXVPkh40ydnV3n8tEV2QL2Cq+H0q0twZ/y3X/
phcIS7NZlRFxpmKrWy2kzukw4sCec//TzkX/2r63sIVrWRCc8P/92+Q/S0EAgAKs
C9hC39deLAJiCGM8hZZSnfVRvAaS/dzZx5ONvCRq/lAJEIP5EmV+BYlGteCI/3IB
ShxENU4KWLpMctBBi1t08GXn0cjbiG9Ra/CLKBkdwns1ZiBXeFr0yh9JDOHRD27V
kWrlX9DwZ6NXErTzy3A2ylV1V8YfGcvP3BIkUtklv3yWsGjvHIqPqbVgrowsWhdg
fz9gzv/gfCsvLo7WH9YrryO+CpO0AA5gZT4hSZcHUWlWfNH61lgF5TXdHAEpN8iN
WbKiFJ0E8XRTaspViIgcWRUi6mW+kDyMz4PN6UbcjO6+G3vQQBgrFFgLURy0rpL5
bDCEofLizITJB87+5y6/bwZ3ppLcwWvCEKilZEAJZ6lWe8aPncfiC1W+pYof91mJ
/hgNzTVbCitT93nziiKHM5U44+EfPVPhaWrr3VidDJ99I2Uk0IDYGrm4eR16RxYi
lWqMjnfQpKIWAmUnD/KZ0uAniiGtXMME/WDzjEszNv9lSFDo+tmoMd8oii6oA1Ly
n7XxRuXAGP6r7FRh/z3UNadcTw9e9GcIPIUmvYRBC8+bqWT220SEP2eWRQksl9F9
ES7rekk4M0+twXdhcBZpU6Q/i4ejo91dRH8a8bmlBZ+FiOR/nqktJrb7QALjefOj
JSjskUmz+vkzEvP7fsFGEwUMqicTXAwne2y6ICFwH4XHk1EsC1hUKVD09t+X++o1
WZGZ+buetMEJWaYvyaWLKMryuyherLA8pmQPseZolC3NcfUGBBD3BxXOTrMjvuMQ
zfiKImWslrSnwhB6iwr7BuNr0CDLcCkE5E0V5HA0e8qOuAyUpW3pgxwCL0GgIRfZ
4w/4kjuEHD+LqCofKrbb8ptGIDWvlWtT6IS2VLWa9gRaoZmezwox/6giHFJ4j57C
oGld8+7Deartr0ljm1WVwN+JkT5UdLq6gZB9D+bEp0wm5MSlAL/2bE7seY3XADoJ
8mZ9UJItmDU9zkb2GiDLgT1i2M0IUKD76ADxNCr7UdYK8gQAXpMF9bJFrWpKW5JM
Zvwr8c1PLXV4N0Dj7YOG9hXuYyT5P4vjLlHC+KMhw5TtTXnZEx8RtKnzk6ReZxFb
tXX0i291O3TqhMHWCn1eNXO0xVvydxlIDYalH+4QHGcchkzCuvul9WzQTfZIWB5B
cd8YZoIW0are9LfqqxDKeqeV575Xi3MYTFoCulWz2f7dxdW2OTXuHqAlK/qRC9OT
Sb74MqMlwKBuR5hMYkqJQMtkpQ2lXsvjWG1zqdHxIl3uJes1WlsUKgbY7WY6zFGV
58MEx4w7MQx9CpToewdiXQK/DyRjAgKiNp1kOvFoV17405nvxzOrYDjpiP5ei0Ow
u4JT++KUdQdMhjn+zWG9v25kD/4rH3wgqozupCG3ielyOrU+8KgzO/7IbayzwTJM
nkM6b0plfiutl6ju/y14haOw2QmWna8dP0pJUHx5QH2T22D5Tdfm/bpEqp+HlKgv
L6NrVBNAcoTKGOmruw1Erabqm9Vvyb3ZwjS4UYWEcntzzMwXTaB6WAcO4nWQuVc1
QO9u9g4VUf7uzKtl7QAhtPQihnI01/4sHuLyS8mtHuiqNEnOClgHulod7Fy2wbJM
kIffnCLUV0lJy7G6wLjIJGqMo9i4R5S85v8EbBC/x9gHurOTKG6CgBRkOlobB9J5
5pabfRR/WQrdjrOXKdNH+H485r/niVN0WblB306PMprulBQ2VhhckcrAoX1r/0ND
y4OGmgOGCfdNyppB0xNCpSX0E25z1rJWXiQCXXSAFN4XQajlyzrCuHpMf1zOjc9e
UHh8Z3RQB+yZGxQrOyXn86/zIzP+UiDENDEeh+IaKsEbEFLM5cYBNbu2Lqx6FkBC
k2pnotO4aLdpWB9BsV1waAbBAi6pX4f4jAi3Nh+xSyKf3Andz/QWKdqfPlUtkpIb
+pA9QJwSzWRIxn9fAxlSxcAkWT0k2l+Sqrxrri66B6bA97xidsrzv35Q7C7wbQUk
rWg8AR6nL7qbGTA1980yHVcmhUWh5P9kVtXHthX71Swn4ZkxI7aKbeIXgQK+0ro5
HPuwUr2hEA2YeeeIkdLrqrhbcbPC0l9YO42wj0cZIuuo29b8PRebXZyJ5iJ9itcm
WZ1NpOE9+D6JtlSRY4khdSqImTERgrmkbhlssWuO65pzRhMKb5HKSdytSVEjmuPK
fBG9dADdrMPtoID0+SztpeRhcRqdjwja9JE1uDJYIEmxHwREoVI5hohjSGnnoxQ2
Ccn9etcu24ngNgcML3HY9ystRifqR9zhLSWsKKnGhErddgd3j3ehIqDxcV2QT0r5
uGpAktTIAApiHcqVRyF4vCiEPknrwGYch6m5DSdcoetY9Eh6rm6pKyF9kY8pgUvT
BhqIsjqrENJNHlljD85HL/DD+3aHOMP6lFchlrWEGlIKTILBwljA88E6wYlBqv9j
xVF+baSkJH9FyHRfYG49nNuZX7r0217yz1iMh6gzzRsjgsPY0kARssuGOlT9QhOZ
kWr97ZvD8OGua6EVWEBtGmQmqfj7L40Cj4uTzlITXWQk3ZIq/9ez+h+hpZJ0fY2s
xjkeTkatlmi6uiKco8Wckmy2Gx1rB1brGRqunG7MuggoIvV861E3IKE+JkG8pQ/l
1FW3qCTPoxsDDXWyEH+S8+6uwmdwOpk8KJm7Hyl4aVRFHc5WYbCO608D3U6Y+snB
HIapSIFmpEp3CugiPG2TE2mMbyhQA9WaG22Hwa9/7O14v6SswNM87FqKkfRbA1Ly
A0bAVipQBoL3XGCV9v72IUgqk/l/0u+jDA7VxyjDwnLGPPw7EGx8hHDYHW6SR+6n
WbKUVQkDrtmpmGtODk6TOSeNAj26vepFseEH6K/hapQ+imdWH2xCTMiutAh1B17I
MkiDQqW95n8i2V+YJfutd31SkU26QyzVQaEDLN0+xer4SMzHu+ILTO9+LplcRn7Z
J1pRA2pwU9c8yFVTq2GTLD//6USUIFhASaWmpe+05RozCDP9ll18wYg1rPTRN/aH
CdZ2ZcWJiSrT+V7GiOKYrPUzQOdWiUVS2Psow33EY5TBtlOt0ayV34F2yY8vd7hC
w2oUNwR5Ukvuwt41BlJO4AbreivZRoRoQD1Tlw5RISf5Qso2CM3UZNT9yRiHdkGT
w48eVm/RaQOz3c9DbbQkEQokHaUOFNN2Ogx/D5F/Smoq8i87CntZqfqDgYhSv3AN
1MQ55q8SCUWJ9b141Hh+kajtNP4kT6yDamJSjGa7Ce9/B5aneEBBlH8CJNesPvCn
K+0o6enetJfpUxXNw2QojmPGTc8Aa7HKH2ux1enpafAnSu0av4RZUA7cgyJoMt+C
uqCQKFznoG6lqTHsk2WL5gXB+WaUO/aQNUd+IEcogg9Xr8PXj+pYwJKIcfV3jg1C
5oh2ym8lRQPuMAhp6D8EU/uaEG+lBNCa9RYg2jCarZZdAyeQP7OMuL5MRr/k6vt4
SNRljNPCRw2EPGbcQItkVqljalPL5x9+EESMB3V9WMciVBkT8T3OkwKTawiXuOYQ
xuuFUgk7BdCaAhep7huapSl35R91DMcKw+KosiLpz3MI0o6p3673S+T9H3UrrmTv
Dkiwc0mkuWpC7ajF40u0NKJypdBpI6bQjaZUz5HdLiZE+J07Az6Z2+f61GmYo9mO
Rmiq1X3ueeGFsJPIU0sGvqegTImjdvv5UCfn1iEhj93oDhOhsMVK2AwbPsQpJZJg
eHPKjRrgsBghitRhUXLo7FtaCPOG9iUfWdHVYzyDm58rFUettcwEJ0zsEI/9Yn0s
tuhk8q7Es2dqNA0tO4TX/DslmH/YioeukVMpY0xn+/5jfnp+nsC+1pklfGIb2BaU
uLIlaxNSSanJOi8IW6MrEucKYv6BMoBGpU+lAReLYnCJIRK/ja0YVlRX7GwjaTYB
H4OpBwnPZwOLyHDvwWpe4gmjGy2BNhTo9EsX6z/E4zas7dUdoRIQJMjmpJ6/Tqfk
VB2TYjAlmszdXzhldjTIzvZeHwgHhLJYpP7pc2HOZhPJyS8ywVIUQHJkI3UlUSxL
GRGa9yxBXxpwkNsHxhref7wNEQy35qnzPbH+ffeiC2eMRgyEVOfXj9N8btcsQnBV
MUnLEoZvt1B/u/6HjjirCEkcn3sNMDj04LQwVHmKuVQFZtUpETxcL06gDMDI08vM
6oRCePEZVu0HQAXSNlrmL7JyO04EDoYMXzE5JTPd38KIBnyVbJ4ArmmOzSiGo0WW
QUNS05/NlPsTHXNBABQx9JrkQ7OYu9NnDHnDEM3sMsTPYMVPy8i916bfh6Oa/Q0l
Da+Fto34Dm6+gjInqf/40CR5yk3j/7mRwUhM34Qz8GG6Pl7IYtC0EPYLsakt4GC4
38yUuWN3ZCkt2PjjMF/KwKQw1JEVOt9Ju93QYGelfZU/UKQGLSOVJ2Tvy/WD2IE7
mw7oEUXwSpo+Bv1ARb90QtbVAp2P6XBR6+GIGacViII4XuAeJbKnApyWD3xh3BmJ
ZJzjjge4ZdjqWbhI8DgJnB3S+tlOz0YdT+R1ptZiTh8v+239v6PO3Lq1YRi7XO2a
mR81ftoUW0+UPzTM+9MHV6ClhcB7FMWnlI1edGHs5EYSQLZDh3cijCU1LrPZRhNI
5+7oXhs40EDkg7sMpzP43GNP8yJ0gHZWFFr58NzDqQRC1LaRAFAnJR75OeysipoJ
FyI7k6SiPl76NeBq5B7z63eU2x++D6KLBo5y37xSld1oQeHDOAKL0FHZgmfuFm2q
T80lVBw5M/tdQynpD85iMWkUpp98ojnXB6yL4Lf78nCjM2rRHtjVbMZQMj/dMnzJ
W5YL8/GkLpCXByVrTraOuWlNyDksGv6yIuKH26W+mlQ1H9OyzTqnSuYERj0p91s5
ehQhHQGUAQT9SP7mF/M9dA48+wIUV4w4FsievJAqzFPPDuYGIgaXD5f7bd+MmfSh
1IfIMxBdT7YHz8Kl/12k4IEnL/8DXnBeFQe00HlW8mlUW10L7uszCTFdfHGbEi8N
Q4DsoI/6RBg0sxIs4GU6aZp4IVwyZN75pIQm5Qoq8psUQL7lRRblxYR7bfuFClzq
3frK4o0J13EYQ1suHxxCcwQF/+gZJr1pdD0GctCIO5UEpjFWygJTMquOi1ETrhJ9
A4O6heeEYXtMK0lZcxu92snw2BueVP33/6dVSGGsp7BmLk9RCT+pAfKyfhJHahNY
oeX8YZAs8iGkBSfOr7d6xE/hTsXchYWIoMH+NQTBQrT6zE4lqGjeyrZQI3lrzShD
LpC+Ni/S35Swfob1dPF4pYbQQmJ1vX6fctHufBFkGNEAXXP5vTuLv/WTEV0ErYKd
gc7ab3PlA0dVc5XDpuqxbBQQAols41EdwL7wptOZk4mLTRAAovDmNsJvBi1yFCte
ddxkAU79l875xC/IhEHaXcQHNyWv0DX9dd9Yu26VDk7MFhvtLn0tvQHATYcMZeXH
OYHIryRR0K0Fm7vzdii7rm05yJsemFe1tRsjdrQ6Iq/Q3P8JY3MzCZTXWwPXVY8v
e7T9/P0FhSFDrDI3jjJT2cmyvgVZbuoMqqkmkyJENFRnkiYQDJWBB26aQ0yQvMug
kfrCh4dK6oZswdZ+vpC4ztrOHoGKZ3DJ1pEmn3sHvxqjGAd2BG6LMXRLkv29cvVP
U8lyoggekoGLrquoUT0ORVdhKIA0CPUXRAahlMCYvrCmAqICRVBm4sfRfhGpYo/x
dv/LSeAwZv0Nx0JQtWkFj0wFEEZw0rDyEM7YlS46hpbdM3UDWIyV0VsMMctnSyiZ
BaohqJUBabePKJ41pmhlB7MSr8QdnpypG4fkHVHM79S7i52sH8AIJ49vDFjC9U/Q
tLoolm7YF/v1wrAWebYTCq/MaSvqd22DSbi4vk4NwNvfHUHA1ipaRoKnKL/N7H7G
G3vuw7c16fB/oDeY5QKl2xMbuMr7OCowSUpTEHlO4mxCP/kSy13WzWYSZlxWJXIR
aJ7cQfun+/Y/MTbl+l/ilAn1IMzR2puPwvLAqSr/m5OezupeDHdzZOPcnP0cc9rv
HUMdZMwl8oXXNoIcewfDu1Ir3weC/zn6pba/b1ep2w3eWrIj0m/b+/xKqe7/2u5T
YnLT55yYDUYa5pmIag3sVe3DoBPuVjEdCS5cLguvVBNOhtd9EuwWUJJZe5mvJPCf
/f2bVDy/cWe+m/LZL/rhP7zsTHPIdSolxn6AzYXifZrr/tRJ9DIQ+eaY8kAUoqZF
KvSc7U258E6CNP9DMUW4wzpT1WK3CsCfIzvIBWZgpAZoY+gaA2maGNOaX+pbStWL
NeLeMsdcrZBzWDIl9Wl86pFzaP01MPWaoLIxzdRiKm8yJId2sJGO3nDQeYCR/cq7
njoY1iJq1bwznU+7UFWeQ2VcSkv36BhMmcTjn9S/GAMUzj3SUD7I1tcYD/dmRZXs
Gx7rkWRQUI77ZN+d/OsITMSG0njUdYH0RWFHlDSFztzrRPWZL9/Wl96ERBjqHzLT
MnVz2/Z3435yNcaiWMtGpMNaUbt+p/Jvs9fpJtxK8Gjsx+HKGz5EaY/S1ecBMmqD
mHRN2mMFVIlY0nqsKqyBnUka8RRwVrPmEYf/LROiON9DMk2BPlohTw8+WZOh4G6s
mSykmUnRbMpvtjMXkPS/N9WTmTJMz3KJQ9wYJ7fFYA4ALlr9pqm/zPnK5eAd6dQF
DpoFtgxzDOtrIJh1K5PddOHeNEZHZfV6wSmoskaOSUoMMlietmzENez/qG9DEO2D
AyHS89Wk0tqU1NQxacRkPmRiXZw7EGD/cH+Kud4Qen8yj2rYVFSJKBBFnJFxV5kq
URmp5s6JPfviMKPMlSO4czu0OqFJqG8Cn/uUIV0J9LJGNxxn+VbLasDHrheBDk71
Jg/oh6YGgODet36kVveT2n94XC72wcbO673jsBkqo5tb3QlNLcLFXWT+UFHssKNL
MwhNUWYrcX4bFe882nYHpFgkI1n9yBN6FYYQ3xvyYvbMNBT7FfkXLoLPcihvh+86
3SsBEyIO3dydo2X4HBDt6eJKaQz2+t9RdUZo/RunKy/jcnfAuKUDM+ZzRXiU5UXH
Eu8znn5hLOYRNwvG/O2ot4uTyh+J2R7cuvj1zbGNlTQIKAXQpnldolI7tv4VF3QA
RAc37W4G3mMMFu+gVAGu2O4XJphQB3BEBuN2W7AJxQyH3cWAsC7pBirdessmZNcZ
j7Sp4cd8GagF3ZQtbTylaDfiupZWzPUSg3PO8f6VPzWwYr9B2b3kXfJ8ZRS28jrW
RNm+aC0yi6uJG/hns/jPxyPkVxyW2+4Qfrldt/DqDIfc5Fx0wvvNrbl3Er6GeKyx
nWMid+iZFfeQaKYjqsbXp3HwQIP0SZIXXP+o27zcA6c5KDdhXMRj0uWtOEDV79AN
QCF8IU5MNFhooWWRgoEpm/HRNCX/2A6zXp4LTEE7T4URg2mAUtyXBveujkZi1q39
lWAjDebskrDienKyaWnVfoA7N9OgqhcxTICetR4T1AeDMaRjUSRuO+OGkGcpCx/L
8Ql8WsUfrpr/MundzY0JXobgwAhY+yiWz8tvg8eBJUDZzDFMCd2dnifXhq0uqikx
RYfC0hsJj7sXbrL29D1/ToWULS03GhkLZVh3KHqTzJIb+VhJEF6DeJtGQbYn18ZO
p/wX5nNljkYdagvt8DavdOuttkbPOOhjrqwwwOGKNHvjP2rPpChR+Ebef275nkMW
2KLfZrBpqQkkrkhR48zUQ13HUaWz8W4oCefKja16aZFmbCDnskD4ElRdpmZu86/j
aCe++rlPMnLYDM8zS4yw6K6EqmnQFZgGBilzrgTznxkkCDz4Nbw7XgF92bcj76pp
m19V4tgZyHFGdDFI5IxhwT7zRK+ISkvqCZumgTuZY3qJ5PA/EKEs3R7ICL5oVxGX
O1vuo4Xyw4C5yFdmvMgl7eh1kbc0sivyMmq2YWnX+8smpN/D6vuxTJg89ZagDaL1
a3OHtEmj4Ozik7bpjPzE9kMUwqFfRaxAL0W90+UG3E2uKLZ6+wG7Q3Nri9DRnE4N
uMkBsAtPjabsRFHNsKn5XKd1/+j9EOuUjZzhddyRzS3wNp3AOEd2LOHd1kCwIChO
Wurt2+nndLV0xuTjXRZ6oAVlozZQWJldO+qGgquhp4b8sz0ZpQaoUZajLwmXLEKB
q7PLMatQhLk5B+1OhmX/SGLrLR4ec9NA9m0Ag9Nve3jOeTiA+sA2O6CfJtbmLeDK
iFyagqGcXlhk0jAQdceVR4B9m3/b6c6Yr0ExFlPxnWjigkLceY40fp87eEcbnzWs
J9Ka255bfa0uKddbYXsx2y7keXX8sBzD+WKSg1YcYL2J9+u60Pxur4d1QXBaYIPR
yyJ2lv19bu+p/0v/7jGyYrYgeerLK8H27dvNLb6HcR4tKAjMSDjN5+J+s2p44uUN
KqG0wjtRJyQS9g4Gg1wgLzKLOUhzbNTYSrvddb/ovNtMrXq/9bcYvzZ2Sk1YJsJ/
csGT+RRWkyTGGG4gUtjbbIAHhJQZhNGCjfcgvplpFN/yIOdxx9JBFCJgbM0gDVYt
YNy/YS3SZlw/YMdnSDDuHTEs8s8vToBUDits/3BnojR2aF7QYDJIa7F9F7BLbNRt
+LJb45CL6Ez5PcxUPq/1k9MiAz/+J9HUbvQ4ElcX7drKAo0puijNQkjMFEoc6LZg
XTmG1SEK6ZC64XWLLQHQQCIByiCpT30A6qS2HMS8W2IuBdmYXHO9LFke/fBs5hsE
zftaMZbCu11m4exGat5fDJWLnqn/zjFbofJsNCD8THGrJpQekC7qbvhGS0FBnw5s
sr7qn7v0GlJmVKrRIyP9dJzLvIWOkDe0w0UOlOvbFXURpvRX/Gb5mX7Jth1z4W/E
xwbiThzYUmSVvGTSvVTaXGxFYj3g0ONyFAkbop3CUPv9bQVomEwy4xrru7z3ZYUK
f9Vrpolcdlz6ywyZmlxUwk+YhTKtFyob82cJFqQUUOLSnGPGH1Qby9kClYUsyR2x
thfp5SzZ8tKIWetiiWuKpbRMtYuIN/iSfQs/2BCPxV6HlgkTP0lEZUQnnURwf+Ry
41QfFp5ACmxNIhU8me29y0mas3XOaKuMvwl2yYSajrIasIQoCWdBG/6UHd2zDZc1
MrUnACl4cajxFD4U7ZJ9JfHNHBkp9K8rimvpB/xkoRZarFIqfi8vnaDsoAwIklq2
wa2os5C76KNe8hymtbxXFXXw2lb3QRG5Pa/JmM2tyAj1NW9UO1UVR7lo3VKU3G6V
m4rj0aq/pYU25ryOivwrFfIHG4Ur7TDpOhGB7lUIVQ91Wb0OSc6vYj+OEoQjooWd
Irp2tk0y/fplzsdHsJi82xpaCN9FGlt42dnipxsqkoO93CWw6hwiXG0Jx8tnDK8J
WYA5OLz5f7E6JIxE5OxoUdAJ842CMSdzGL/hOKi42S7A5o9wW8kpux8sV1/+S7G3
CqIjU1nFrhXa7YGyGAO4GAxRdjnalTSlbHh8vUDySABH1EqqWfSQX6NtWQYwWLnb
nkwIOE2r3irc9d24nTx+xrMCBBmUJ+roogdw+lqDLxvf5+/A3yyn6yMRPXNJH511
X41LAAF1ukq1s9Kph+zTU0BAHP3BMEDRnihu3Z7LRe0TGLvDw9ec1twD2ec8Sb31
T4hKIbuG7ATSBdICrI6dZppXPeRDr+RMpMTkdWsgdKJLsYO9tnyVAOF5yEEJAaVK
tHQuxwmdjojCq2Hruw8ECYlUq/ssg/7bywD1NjgA5UegJey4a7magxF/Wjx8Dzlm
1+deqFw1eOti58uG+odf0llt3HFHr31w3GsnTVNnUqBDbQf2ULfIhV20Gi3uEBDL
UfrBBBUk0/WsP1ddHX0lYpFNebo7/OPAIe8wTnRDZpwi2nw+4kxsIFBPxybePKvA
661pBsGDsNYy7IqCfuDH3Do004HQpb3mG5wQJ76cxBLjW1b7myOd7MJ5YhrmgL3c
gKfKoVSUS6Hd0V0jKlP2HvMGffKwtFyhyw5GKALo/ZlFI+cki96pII8VXHP5WUfT
5FSIL6z+4F1t1Wiin8AtA6r3M1ev04hglOs+TDFcXgCdZv+sk/t/P0p5C9sbpML5
9lCfV3vS0BsZDbw4wm85XlYG9m3h7O/8DunAwofcnc1G5ONELoSy0NUFGVIMqnVy
550yKZX23kQ9/8B7XZ7OXeQO/2UM2rh4kefOy07QmxlZoSHrS6Cy5X5UDJRAplME
tLm3aW+/hQdzM/UmUBbpumxljplNvV8K9ZFhgOFVQ9zkCUPOVRP5MowFF8FvA9ni
g1DLHhe/ZNg9+wQLYw15MaNc52H7GiuVE1X8VgDUeFNDGhNRfVGC8l/7VH8i7Mem
002ZOxGRUhvkcpPZuq3ND4lvjpt12ua4+KilZSjyA2OScNU4MaqJbl7tgEUMyxQz
MUacA1LXSobHpHO2NNIEvwQfcwkW4RIwX33fHduf9r+SZGzj7JLMqzYpw2w4Lmle
uiHnmkNuh7jeP7xczaV23AW0W0gdJAZ+4QHY11SUCVSf6tJMnpC6Kqlzcqcf4dZe
Iypvmpl2ReD8T1Q3bJIwBfkuzcqMoDWdLUWdKG7OsZp83uC+oWL4z4H8x91yJE6u
4ChRnSnwwLj2Y5MI+y+bgHyCA9MdFGzUlPeFqO/i3EeMwHHx0cX1sB/Y06GvcToK
EegejkDS8LBwjSjnsOmMNRuDANuHhZtQnST5EGour3nrJTlZHXIqKdknKcPZ6Wgt
QU9j6LcY2xh9qSPhm+fsNXMObx/8JUOQhXQB1BChgE6h/onfrn3OBLVOYQ/5zglH
6xQbueW2/dRd8/duPiVhDt+uZSgTc80TSzER0JiHyvBXTh/DuwAInSD+zTcG4v+z
WfRaVsON//b4RFq+lXhaVwf0gBrGub/WM0kIGWRbSZ83aqDkaVSELo8AZxmIIMW0
jbZzu4O49NbX4RCzGnCbWSjGMrWaFk48IPuZduYq3qCDRY1vK0qSpyxm2cP/qKv+
CL2Hpu+kk3v9PPjP7zA4Xexo3iwJoa2r5HyIwgACZ7TlU9PfCyalBsnpfVhuYj6C
kGgivE92etOKx8KaPbmLvdmPwF9LXUIAXI0WMFgT75l6LGyQK0CK7sKAWSw+pIF+
1MgNEh+Qm160h7dtmfEcS03/HL03KghWQSMaGhgEjUfm1uMT7+6JQHiFpy3wIxCU
LA14/tHAgSKXhKk4yZ2ajl4xqRfxJ4TCeT6Xa5Un19NaDyS115YrHl61TOoixnq9
l9xrtd0a5UG+5NBQYzpEt9MF/asIAhEKM0fdJoIplLb1towgTuECSRcHDtUpOR3y
TIAoLD1UGD0Fbg7b/MZEbOE121VZPdbpwo9u3jfKEuMTAMiRDGDcQldDm2L9GKJC
bzAxHjqgQ/5cvNTDHBy3Mj+VQ+F1hXtToCZpXw6QkHx/yxVcGoWegNRTDIMqNAtl
cyuaEnBPiiun54bVjGJIap/c5XK5fUhfunH5bdGF7i3YKNbKGKShPtU37oxlaIjM
RrDgcSej9CbtSWGGxnVod0V6OCISm1mujvHhgmMuyI3VYbKKI17igrq8wnmxaz6R
smkyM+2mlHgy71WJ0tufyvfzBJe7yUq6GHAb6Fv0QnzNUifqgFRWcUGyHCtCjVkW
DYK/eSs71Wd4FaDLk79lOjSZ7lJwi3M0msBDkOh/gj7lRVxNUuWfEeWXjpwLyWW6
X/TacFAs0vV4tD/Ex9v9eYFqzdoqoLJM54R7GjPTTEvZy5J9cgcDdRFq/1hkBDDF
+uCrck+wAJSkzOFICjndISs+jtmnHSM2+r7MYGv4TEi2rCDhP3H79xg7Ca5Xt8r6
MIBVj51r9E0aC49Rrxo+ZPU1QkBWJNQ+Vfdgu562k9T1zbYPvGy736+q5r4DHMLO
+NBLOHJhpUsXt/3LBJQFEKNRweTyI+V+ZcoAazaPkR5tlb/BnTAzZiXD8qoj4ca/
7m5f0CbcIym4RVzWAm9py3+k5TxFKgZL5eXgm8WzJ5xDnKWLDVLsk39OC5uSqpRV
MjClqkw1XRWwRK3MW7US022RVFALBPre+FNHq+oMGSWgmsAu31Nav3IoTPcDUBT1
Gy+ZdwaVG+en6g6efJkjlv7q8piOqHC/98zj73+tPHTrvNhuXhbPTjbJuRdUQfPd
znD/O560gPXxHRdUjS2/UqN5XAzJ03KRV5kGydyef8dUpQg7hT4UTK9SN4irNxvQ
3MEYuHZ6k40v8rfWKc6VQvAa3zrNElsq6VFC1Gc/kx1dbHaMtOOjelKeKmMVMhZA
Vubaoj/KLdsxrIjSGPtqjNM7CPefAzfXfr/mClI8crzLs8RGQK82iaKBXgWjDild
9J9rWmGn4WvZOkjqttDzzYu2D+jHeX0cFC19TD8MlqgmnjNqSq0vU8gPA2EhsBW2
LpbbPp2Bm9axvl28kLrt7XBf5BF/E8wvjCPW+Brc7Ib5K6loNIDxyW+0vQJze1b5
+uE38yqCllWtyiQxf7LN3OSjGGiBG+DhcT0+Qh4t+24+LW3wM1tNrePeExCHeDCR
HHvPv4H2OXyPqmS1lEOfyDLoEtggTpamEgEE9iKgQ9LdcMP/9yTb1c5tnQLIM7Tt
dFSnkbXN2srmZjFjN07ZWb6O9hNrBY0IP3VZv5SarlUeOocY0q965clfuAUh4aiz
eTXOvtCakqoK6VN+9vZtwzYJxqbZKeRS/E9ayPCL0ZUqOem4BSDxsM6/aNeEPtJu
qcMLXAHx6+Xgti6rE6gDTKRx7TtiDjHrj9Pza5Y7dVpiuysyybN4ugVdffUapcPj
PJtPH2pQKy+ru5JzxdQYufL1iCMyXq5RQjsZRnCtJfckEYCuvJeQYmvJQnvFJXgN
4sfffPHnaBPzOv4TlK1rKBR9LTW5yVd8YC7YNSbkkg7HhYWbM5Rwq8eB0G8nxuc5
6z/+UgRwfIl626frODXLbDwMfp8wNhSs6h+ew1S47KIPZ+3hQst3gfLY8qBuKFEC
tklbfwxDo7gv3kVDSmQ9VsykmMEvoJAcFzufAcUJ8wNVzKlCl2J+LujSro3HOCh7
CUmXr3i8zTUU2qOAWb6WVP8XuTkGvWDhG/r23uv/fzMxOnrJT1b2cXLmBXz62Dsy
4wotsBEcwGgkj7Lk+xLvj25SX572SHcBcElz3s2fuU4vG449185jN5Mk5uJ1W3dK
PAjfLUbrTeqvDQv0XIoy8QPrWhEWIjwTnz3wTitar2vE3zCql4sqcLuLF95Kl+nH
TfPtxIrHyrIrbadiWn/NweobGz7LPUvkt2U52pokSUQGhvzQQzHrPg6JvWNmFji8
nBDFeI6mdfxZmnoXYDWyCyXL19oMK3f1ga75nVgxshpd+Q4bT8IjZM4otlHqZ9y8
rxJjGVSe6YRmuV4Qi3QiiANbQq6xD99HSiRDsCqzNdi7knJMbe3Z5rb9h1ByJWbm
p1XJsmHhbtLAHiDOu2ijcGRYuFNKdNRv21ZdScOu+YxTQemwuDsmSHsQcmFoVkB+
sVo4AajeQpOIpSNNzdrKRpFxTOaYqGRjXqMB3pz3a1G/WverdYbXfc8KfhxdFPdL
9h4cuNEe76CrrQW6uxmH9RHvw6bwhUmPJCym1nbpoIWTNAJCY/H3B07DRDXjYH3D
TU9KjehYJe8zuwtGZKVEHv6akZuUGI12AHYcg1BzRuFtuGgcpLiE4kR5aLcC8fy+
lveTzCnB9PVUVaQX+SuwEzeU4/Ek4NzkuU0180gYoqebqPnEGGFjFHXkzVAOuHJo
MWgNv1+9zD1tAuGVBhK+Uh2+NwqF5fWnGWLM7FgmDm+ERXTZRhA3V9QnpY/geW+j
3K9OeAWEwJq91BTHqaXAieX1tOazRVo6tRQXVPtNo25kWVtSXU5743PkY1vchVkB
Z27hyI0qJrLzRKx0Al6wNZoUheK13pk4AIEOueUPKueyxSJ8W9DE90cgzKV6yTWx
Bd7ZHrPrrasJdOkyRbOFJaY0JB+3KOrCbCYK8LmCg3gFdQvj6Qi8VqQc3hoFBJfH
+tnCu7Nz95gz+cHFPc+g7qFHBhINWlpI+reNwRHqOLLYBaznDmsN1iJIkC0yvRXj
V29CYWOqLMIGkg7Ig9ABRVMmg8S8UYtJ+f6K0RgDN4MTYZC7QphtCV9C17tSgegl
5QjRsh1H+/Uz6HKwllvjCDfsUjXHLTErM36Visfa+aQeuksCgrei/MRiLlm2IZkk
xljh6cW9mQRIXLtTNG6rEb71KkWQhRPnXPhL9jDFihr6NfyhF7wJ5WQmu30gkWp9
S+uFAVV2SKK2Kfbr6Gve+LTyl3XNtEJy0DaWHkXh11c9b2PocFvcq04PDv2Wh9jy
aGUScjoOBr3Sr+cjqN011qQZIVhwlqVF4hoVsQpso32MNpfbPNe98uoN3rH3vKNN
WYf3/bYCklGnkJdw9N4N8G2oGiSd9/goA4UM7TFj9DL9OzXEuQk/KmtiCZGVijM4
1yVRkoeWxgoV05rmlYjIAHE6JT7tZ59vQirArwxyvwhhm5XI4OVnu8YCWY+Dlvdq
tyuCZlsHaPN4VbxPHwyDPqpM7xv73a7LfVpUg+af+438n0vW0JRgort3lv02v2Yz
vcBsOlos8JRQWdl79FtUZQiBjx3Z34AkxzYsc5Z2l3JrE2pZ4NQpRYAQDZTvhZ7F
OZAfChLZ0zIFZfvH7GOZgHPZENMitNo/+epOOaPrgDKkMuQFmgtN9jDCCet2yn/N
ZXzWnAmlMI2ndCDDmG4QGSSwWXnbInlEkQ2uByNj+te6wG9sonDR0iK8wdg3ROqM
TJ86sLw6/8JJKM67+hfNkAro6r7F5nPFSd0qKJdCeJmOngP5qc84o5mvVRlruvP4
Tc8HlClhoib0cb2QMoE2aM1QABZOUDTySivevUKje/SV5V9Pt9/9ycOx/wtxbPEI
B2GbB8D52YqRp5B/6dT7Ul5X/BAnUerij+YjYZmftQah07gDMtrCB/1O/bpapoJO
KhwVRNHZLqrsyUQqMt2nmGSFzx/C2h9ynyyraAvbB+obYjYyib4GaCIEbrBLev76
N52rA9Uk1DQ3wP/x3vjkwnqSA7LkCb6h7f3cW7T6GTOng9k8n5U4KA6gNuoIEw1b
LujJOQWCUHGVTE+b8sHmTIHGv/kwQiaTRdbq9e9QCQoJ74xpVCCYIR7ay8ytudoQ
4ldTYM9cqwXPOAZMzctSxmvQXW91V/Jr6TKicpnkFSiw7d7roVW/4qTeYvu+f8zm
clacBgzfIVi4o/vipDX3ctARBMMS38M1l9O4Z+pW6G6olpiabQM6Z2CaRMEn4ZKd
W3LIaMqW5j+cgHnYbaqxmeHKJmjYuNWVRHlIz2yEoFEQitAGrw/N1Od1mGhsmcxc
gMyi58DIHPKbsVKJUUFsEKFnGTn+uwWuLZuJVTViCLM105OsK838ZT0WM2N06IKz
sL+9O7lgvyTRi5GWob17gPb4kIGuxBhGxP2/1GG7jXFJkBWf47pPwrf/aoRr67XB
srnidvftlw1z+IKq+9pNMdJ+joLLDW28hfgd60XBGcX7SC+erkL215f/J7BmAlIo
r30Cbg21NYxpkO3uLPDWVKY6GNMUXdqmsecn2lCfr5i0dhtEfz/d5qTk9QIuMFNb
DWQnrptIfsPY2yqB4zfyv/0mnX1aTHCug4xIKP+tGj9xJoevS+zmJuKuFWuNxOee
YeDR3RoEivFdBC6Kl1HWpZNyYH52fJUb6zVwsxprTimYr+TO+leRWZ00Ez1UaUJA
1BPxJ1bH6tS6b20SmDkKU3Z2ZAdOKyOmmoRXmLkJIIon7wlZN0OgrxcTkAh4uJK2
MJxEuTltK9SOxRvvDx9YrBSmZZYm4Ztn4W/Kr96SH7301VdXEAZ+Og6dW7BOXWpi
ErV4bFR4/INngh0z26AB98vLFldIgIh7DExarTo5s1r3TVTCJabt1MZ/IZALq27M
VBu5Yyt2upiBI2Xv2wH5ZNmxTXpVWAF0HUfR1U9MA035QmWhmhLKqegp6hfg1kbL
46QvgYIwQ2LR42aX5zwrgiOnvF5cGYiEy3rPDm7w3PLvUeGgkoEVWiX6pT7vkBlB
sxEnSWVpLyshmzziDfk6scSV47IBMb79RZrJCUL+FfhBzwMa82midsWr7Dp0X+R+
BVWBYn7GT+Ef/ZUgvXJ3werFCd6JrzSH/htF7kp0HeeoGSXrzBw120VobW8Mog4Q
1JosY9Lj7A5wN9i6V9IgNkqcxJjhncAVI5NNvhc1MD3V7WFjW6goxId7nnnRcwrt
2XTFfdnZhnIxi0RvHGkTrl+ToSTqnmCIXZ9i83P9LhAigcsfI0g7q3N4DEmXGWv6
0uu+AeVeCL9bPIfR7yBM7kWziyUtlHWG2VFiyiUwKdfLu87B0SGxoFmYGIPbvei7
aH6Up7nlgI06DOLhibW6GBAOVIVlpMiW/KFmh+bz+UIsN9Xt0HIq+4uf465KrP2A
Ovf900EsNgHp9dtA3BCm8oC0MCRsWe4kdpsGFoYsrXcTskym5n9cgOSVBtazvGNi
3AtdImGDFu4NqcrN4GCVnQqwN2vNpYHOudLKl4ujxBqJbff3tAo1rlFMKBHNmO7U
2Tn9emQaeRWJ2XXuxJLtWf999k8CydmxqYxMX8Ob4scC6rrv5kWB1P3xz+TZJ6fI
lyBSOhy0dPa11fe1baWouDjMX0AnOFVuaDR8s1fzLa7FRO879qjxE3ZjKZoN3F/X
rMWI1LQZOWlwwZOSwhOV9mbXSyZbCUAsaOZENyfp+kbPoDmHv9zLPxtusDx+y10w
CkvuSA/soGS6sRAUc5UeeJYbWB2ENO0DdIxfezKS4t61gofgB45gyRNEiaaqZyPg
v8THtD41ixmaZPEIvw1bJPCkohFXUsKNIyTHILx3XQp3cVCSas8bLMggLXBORvRX
08E+Or9zqaZE6nq6YRwCrLxNdd5xNfmaN8USMZZGx8DMsVPdbcg42gUIw9Y8TJU0
W7Yabx5gMNNRZrzueWXDieJlU2hUFD8l4nOuXuqYoPDf6PYtpfV7GoXP1ycxrouA
OCkUM5G+AHVS23x+qhZo0BMhe8ignYiCDTL95e28Y00S4GuKmLfMxyK64hVjSaTI
u4/tDx+KuoQIj4Hb4l6M+VwyTtQ6+U/eGYNS1BaW7v00kVnvXWU1Qz5PceKhz191
Els44KlM/m9jlm3cT6mUdu61Xm4hAe385z4GwqN5pY2vPiNoj4BXSUjBV6QiacsW
nHQL+LW1DD8Fvz6RPJoerygw4HlSCk8/ozjN++atPVgiBVx1aDlsSmvqtE2jYHdL
GD0UI0MDRqN2FEwr3yDVow8APr2brDQQHGqPoSEDkPu5iUdsoQZLZfLvRPByyBoF
YkA64QTak9JL4pMHK1s6qgyENxphSDxLfeHlYhddJsRBYZD3Ge8YX0qXhE2LlFlt
Pu7eqSiJNCsaOQTlDv2TeGdDH4UVS8p6lJ+CFmk8bZk1L+llcanc8rucv/EVKGv9
pk6Ii66Rz6/LpJMe102uWPUc310WDIANX2c5uLBAGgTBWlYCs3Y+lsLqnTuXj0Il
SQUxIlB/RkiFrsUWzhZo51S5vFUa3A8CVEtpLRLR8ib6H45uEY1RRJJSOwUkRBq6
fAxydaAHc266mMroHNLmv2YkQu/6lhNXNu/NXpFCbqbRaVrTr0/+SDKT/R9ROMV/
XoklPyVQzk1rb8gXN9YS8woSPt/X1RKW9s6iasYBgBf9OdNdu6a+FosnHHoTj3Au
UrT0Lqh2XvVTMpLM7BlTuSRfpJ7TKqlF7eM6bYM6BpDzmyeSCK4ouyIupls8x7sS
DsDluAbLh65enr8DxiA+gIFef+rnj6SQWX2DdPIhgFVMW2vwtyZzyd9MtdVi13DF
HES8us8CdpG50nMxmeDGrWjekKCH2aMJFn8uErbd85JMKaQbcprVaMg7E0j1sdue
cNr4c567c+HgLyQsyJzNkL+ZHv1dRHvi1ZdSAivHPF7QAKUQ0A/6BVshMNac8gEm
1bBfHuFm/JFBMn90HaGj1lAklSfuVqunWa0RZMiY+U0jsPOZGdbSi2M/sKQ9qxYr
m0umcUtemo1lXVRiMR3x1n7OpX0LqXnJz2EvA4sz2b8fpZhYI8tQdlekr5v7rYGM
9tT5MXl0BCvA0ISyj7Y/UIVlvetQmRxBx2G5rxl+IT3qOX/4bmu6SsJ9WiX+9Ol0
jrd9zGtNuunF7UttvjpnLJ6XnZjqaPdiU1q4DHIkGzQ0jZvXbXXkRjbu8mrhl+0c
GYFEv31bU2+iWoTUuGEwelFrnkI2pOZqMTwud2xOkxf5N2ztKVMrowioBlFZ2c/k
ZG2pOR1Xttbq25zXRIoQHz5gcCG1qe9AN0QvbxFZE/0b4Q4cuj9WlEz2IrynrWjz
z+wEaj9sinn42Vd795n7kfl9yASA1Y+wLEHQCx6Yz3LmdSI37O+tDFpS1zQNp3nt
+sgTireILs8Uhwa2Czq4sKaPWvf+faH7RLsPFnRqHOwkBOC6DTB06EfZykOfbIm0
lx0JTXDgZCe4G2oVkY+vBCdfghrD/ukorw0ob11ojTDrgXXtBHSRM9J8oD6Xfc5Q
qBQkANuvFLEr7HHtRzffS568P2xHixNYvskwURsiYTaLLwG/GprHNAo0s54bO5ky
Z1ku/ewKcQfU/yE0Jj7EiBx2BxaFxXJtzlbPKtzNP9URyfxNLfX7cDlO44m1oclK
luLHKzJmGjltReLzThEWXpwazIyuCkOJBmcgsKm1h8pe7oeyR7e6+hG3irWRT7xm
dzC4NmuSagDPq+Q5K4tTNr1TCRYzdEXyL1IF0wlBfB7C9L0hMP1rybzzs3b+9sq3
RYcpSmZEDJ0zM+bZztKFMhvF89ZiIdNKdZM3Y+UDey71d2bjA87NqR6/lrVRdswx
A+PRv/39YsHsCBAhilaYuTQ8T1bm4e3YP+tT0fYq61DtfDxCpzeT1Ye0D5dIrplJ
nXnHhe90cih9CTOgzmyk+xWE1O/BYu3o2BBE/R1iAmCVxF06SEdxMWWTVqIND/B+
Zu5AHvUnQH24T5ExQSoUgL0r9VORn8CRxF+uHmcT8g6l+iMM6KgF0b0my18YcInR
3WcUjqBehC9EoXmdlwwPoqYhl7H1AUKY08Hj5a+kzidhH3WuFU0Zu9cGBFbBcGRy
d9oWljoo9ZoM5I98VyYNk2xdxb8CZO0yFO1oI6NgIWU8/euszUqO7Kvzh8QlhUbn
HUcJYcQCoiWz85xLgrBXky/absHXhv9G1s9qTOyWU9aGDlZzlxemciNTH+js+SVJ
mmLOEum14BnTDHBunt0zoGoWg0twB5r6s/3bK0g1YMqyCvZUm50/KFrGm3ajJEkx
4a6Fbri10E+tU3rjHSNa27gi1gS4Wfc0UVGY6mV8jkbaEyp+bpSFRvSp+bfB62jp
8zphXO894lkdVXA2c1W0muqlJ/eRe0jnExCH7MHM+sRkgmshfXSZ5uE6n1EiD4+a
DAXRFgiHf3FalEPzTKJ3CCb2foJTtJme/1X6KcSQwjAyMsjuYJ/wt+Ov+UtDuSnx
Wv/cPrmXHU1ac1EJRlMwDpm2FngIFYa0QOicCDAJul6X1pwJIc4j1Pd9s/TGXMwa
b0hiLC/gOwG1bD5u0aMLkhB0mE6wlW2bf/cSoNTFAnXKGcEF/2vgUO1e7NdQs0fF
39Pa5iCZ0GkTRdWLfqcPAxEL1B96tu0fiVr1WQbqxOwmrC3RdYou9rtyeAoxU2Nc
iJBnbPi3xBwihz+iThrjNqw1qd+m0YLRfbYX2uD8uDhMqKyC0K5QKpQnpzGkwH05
j/XVjesA26JTHXXjZBeadWrBQ9BZZBqt3Scye/nRxwA+NM/68V3Q2FAIIIynDiLf
AqzvWJ5PJVaJK2VGtql9To6M6L/A9BmvQV67rHH6RnNAOXLD0lD0DQY8O+mWwe3T
vCFy3NFuY41gOc4a/+usdOpg09olkzwNMxzXjR579D1NRHdM/3u/P9t3Y3+MXIY8
scEtkLG3UR0IKZYcaig3jE0d9szrUtjjtfhMTOqtvf+FtfPw9LkUyoc6/IkM1BR2
5szq53ZQwXHH0C41HBRRxiAaY8R2YKaTcSeJjALIwyAOiJKBQkcIp5/z7mASpS73
QZKvaCBmyxUc8/DPtZUux/6r9BZT4MfdlDKUGvkcHErWy0Z3eR0CXZg61BIKQm1R
YsCf9jaF0QvOR0/bYZhzJhi63s1O+8iMR7js5FTHfqc2w9brfp4/qo0ouIP8C+Gz
DKNBXyxMrRvvwOxeWr79dsrxop6zMsqX6yiXzmgN/WlT8DnmXgbApN3Fhv9b03Qb
XfYqQGWfCi5BFREfa4dqYLrUX2E5aGxA+FehyTGrMjdvX81AS/n4gflIXg2VZkEo
czSAsxdXBa+V8vQW8h7kjlPokvLVACJ3ccbSdIB0siZ9tgeJFC2VMdCF8abnWzY0
KU4vR4uJL1JGgwtRfYSzs3VqmBuSlcKzvD+QxFyRtPOMSOWWThVYRaVoo5YtZD/X
aaxHU3yE9qhDwvNogfFU/bQTANbmvM8zft3U+Yh8NVqmCOCB5udGiWR0xG4JLFTp
6krlxXLIE/d2M+3pun4++WqYqD/gAY7Tc9rAlC3j9lek1VCZLggUW6V7VyaPm13l
FHSxPRTfSiV8mJymwQeGvOW0H5L7v7mi716Az2kTUROJsbGkwNmi9Yru5i+1co9h
wg1s70v9eJymBs+oqUkV22FXl13DsfWARtRe6fuETlzUpmB9dzwkzBWyTSLOi0mo
EA2cq9fC7HUJUBF9+vgxcJPTcfLvnIKLr8fhaHJl0Krj7GBX+PGz/16P2+sa1pxM
Iw90MObtty0bdPsSaIGb9A8wGG0o8t+1dWkscFrdSH4jLLuXIYdvPkeYJ0Moefu+
D6XtJTxcsIYFdSpgaMH/ujT6fgETcuB2NNGma1AYZWDqVffaU9JTuIskZ1pwyr77
+64la5F1B50UZB/+3H6x9TGBn0E17wpr+pDFi6OKRVfnxrrO1TUP6yYNP853Fx5i
cZG0LY/Z7zMeFi63mF/eT2z3NhDyIFKeMS/jzQWUhNrOfQudkDlqdIx4lujPXviV
TBSzhAeBLO512Hlx/HcV6VWqQAk/7MvUve7WL32Qw9Ptdmb5T9AmZIQaXPwK6aT8
/PJwk6/Ty5NZBWNc4JK72ScbeLRH92Mh787CIqHBrLz+ki6Ccf1CrzYpN13kMHiS
QPqZ58UF4y7Jm/rOTGlRyw4uFdHtWYrbwX26bmgIR2CRLuHajcucvQ40aAvHVcvC
MHn3jhwIG3DQAeGrYGwLs/ihP5ZXoFU3c4c3cPEVERzzMETDo7IC3WiBSQYD8w4v
P1bx/KdB4ANsA0a5KzxGfRsq5bPISjLAlJbPAhkV1BS/JIjirvjCYmkgu4rZ+M+U
0J2kWclHYQMFId7j7TMB06PP885Y47ExRBa770fFqv1915bGxAFj8ZgDy0vGHn+G
ezSm2Z/SCJwjbkDVJZ45o8suoIavtEAl2JxPSdM1SwcmQ2QX/4higtpHwEbLGYs4
zC1+OBjGgyF4prw2f8Y7fvwyKYFLTv6rHTOZYSvLSVlouIfAFUf1ivnrs6ldftrp
G5jHro9Smzg/jSpakrXu4/vo5Gc+KNFGS+J2oe4PRgCp3sN0VVOzazmla/qhTEm+
RX7hNbPxAIyvNp+jxs/Yvsy+MxpwRuBZHf8xU7VpNwJyiqln/mgkqsX4RpqgF+kO
PIvdqoXeb7hjwGjz4WnjEsWaYqO+2Tz1RGwCqqkVpkejZNyGuomf7IIQsSmrKLaN
l/JvRrRWnwviBEDfDLxW6JmK4/H4LV+DwaUFxMgCfPYywUiBnDZYl8naWHXmHjTR
BaMBHONeghe7j/xLeSvNfm2scsmWVOzRJDlsSUhA6E/IQJVwTW3NjoCdmjnCmtMl
SSsp5yadHrcRSRIN5tMZIYSPoVVfyE6mekBP4p0KIWiWo6a8JZ+Ztb4qJWMadB/D
hdWw3P8US1arTNk24+PJOhWu5+wJEqrBIojnd+JQXERp1xQYT9psC6QZwNYxwQKF
+GPucNHHhkdEY5q9A35jmgAIj02iX/l17wOvUx4n/+nSFbhOmxAyEOCJ5xubd2pJ
TxaDIUKtiHWrfh/cRgsney6cyiXBEb7Xc+dcImdVDJafBbxgbu5qj/ZP70tcuUR+
vAM3M/oTutJRrDhorfl8rADJAcd6FBkMQjzpjdqUmUxfHh6yK8xhsd11GIF3jza9
fC4UYKdu5xmhHpS9bRBG1CCcZvAitb02JByr/qZ52j7aaReXBQNkxzjCjeOBENoQ
OMTTFOcc8ZOx7qJ7DMwZVFqdH2/xKrC62lBbCILGugBLHsyz05zy1IAJVQeh2nIR
La5H3Cgohskce9lN/ZIkOPA6CH/ufa7aPbBsGcnLYFG4x3QO5HUr8PLs14y1HvvP
zdlppcVfo77xY5tl5edEJyEUUuNDmfiHQq/pGpPDJof2pqouuspUh0a8qtA8+4C0
a3YGjPazfO4XYyZ9WYkTl5WvDTo8rlNgqywHGryDW9J0MaUSVhcEz1Gic1u+dTm7
W/bTmgmFsaxUy1cRniBSH3Ug5xDszBr9/iglewi9e3Gp0KPFmE1LhmKh9ft8vIFQ
rs2xD1m6A2Q0W87b3inSIoY+B9G8Z9V5Eh38bQ4AWb3KiripOkSiheVdsZcTXzeM
t+St3esjQzmOfn9tOJmlijGhvw3rWISERgQAqTzDPZBER7JrxbFtHqoGov7UWdVj
N9rRinn+LPZuTa/Dxjiw2tinR4UNoALm5g0sj4qnI0GjC5l/I/II3Lt0VjkRxO6q
TPURkon+WzvaNCNJtx6h9qTcyvhxz95EcW9GMO8Ul+EVGc8wTcJ7GbgfSf1kIew0
maMr0RbbCL9ZN9prANKzPNYiLZ75fBX6zY3o1RV9l99CMNc6UjnGaLCBuZM2rR0d
ngr2pgU/idwp/+iXgk38oxe2R5eZLaiC48eU2cKxIYH07fG3lbnx1foN4u4Gv8QF
aAhJ7G49mfjkpoYt8bCrHevOed7bs1IMXHTvR6NYxTRrZu70ou++JYQDMRUJtyNs
B7C7FDKsOc3hoW9rw3YxO4jqOaqQm/cVcZUvQbzvjQdao3Ee4g+ea7PXVAOI7fnd
wc6mSRILy/RpjZ7vR0R945W1Q81w3Bm//vYIRKYEi25BmdBOgKarUMjgKR7rj/Bn
JA5iPQKjmcbiYJC8qYdpQh/DG0Wo1eTs1CFrIRTDzGi1Bm9NAEyKz1pTjRI5hYAt
LzlC87LVPoj2bpCLcg4KHIoR5niiCrU9fkWN4KP4mRyw8Ders315Frr3QFsgj0fn
Sj5tbkCIBMbozLekGHpyP18ZpPRsbRCgm96wT0Gu7r00d//ty2Wk9BTL2bdzJZxL
CU9rPgyxLFpf8H5q63w6c6LluQ7aBOJ177smE5sPTHiO61ncBs/syooc9tPYyAUU
cG6ZNGaFHgWKRt0vIerBB/txtwb3UJXWU0fvj65ZVaGra/rTFuY2zTPjBwMyXouD
oDZuZoEh+STSm8znWQpf8C1DLM/+lg5kBTQhzXx2uxsJVfrdxcX/iksZWCFoV6Ho
d9bRgHxJp93ydNkKFltljRt8QjhD7T1aYwm2BcntN/ElSgftHqWdMLfN69N8JDTK
h3KpeIL5LTgN4j5A3lvZr9W83l15q7tAV8QfHPB+c2SCufwSznnN1tVPhrdJSQIK
7bZsSjJl7jTxLfB94GV4Gfdv4ubn75APRwrs1l5bREXQYzIxjUFlglVbdw1FL1ff
AiPS4SLQvCGSCA7dkgZZ5WgUZlg+Vs4rI+acvolwQRRQN7zw/Z8ETfPQRxPJJ27e
EIJEDUgBFtU6pUUVRW/5w2odAM4brmco9IrM1YY7lj65CFMly4hcpvfA+xjqfnC1
lDba4WNi6CPvjvvpTSuAAiP/jQStBwIgf/4XSsKBy/dFIhwZ7v4rOLyaOGSZ4HrB
rEmBAiIh9tXQtaiiqJJeEOwvNT8Q3s436gj1IncZjcCUfCof2U+m4blDYzVr4Ikd
l3UiV3F+G7WG1qMyBCMY7MwnA7oZNav/1O3SpnCtmuKeukBkU4xg903QumpspnYG
bkp+KVDHBQQBY/zeHjRT1kL3EDhWsKYvMwEl3iR2E1VdiMZFcaiOnK4ZAgtcKkP8
RNcLhPF5YauzkhDSnF2C5Sk1Mx0VHAgZ0jSupnYt0PVkIFNqKrfWpAeR+BoEXLAQ
yFOHLgjDAXg3YMPa5hQxtApzpJovisXjMSb2Kinpgdi1piOSNz4oEqUnaCyavRgF
oQ2D6VM84DETZC7MvlrhM+KiFFyRXQ8rFlPYhZq3xiGYRXdyYE5BYUvlUvohv6mB
iDFcuy4fi5iBDLzOmBU7G/azwOQqpz9UFS+9HSRbE8ehMkWUp20qaYzJ2JQ4bFZN
S6SeNafUge356rOdI7SslmHXEcUHGBgkSVLZwQrrqXhRj6qqK2WH3RS1Qy79C4Hd
A0Lbv0D+X1JXYqXZ+C1+a3T0Gr/aLGKn6XhflaPvPSHY+rXTJ/JTgYVQmxLhEBXg
tqS3EtKLm7UemOK3nU9fXSYyDjWNi5GRDo60EpRqEZCy4RsTlgGLwoSF+CkgqFQx
lolakD1j1oqjkduzN3MAFx9nY1r/gZ0HA73iwDKUVMVbxlEY0ADbfSRm3crxans4
11CocQazeNZddH44+eKFPL/9itbzc/ZuO1xtssB8Sx9PphMgRaRub/Tw+oToo6nG
wYjMSz7opZAilPh2viAgYcmn6uuPlM8HpaB5fTu6JB1WG2Osjn5Qbezj9hwzsR0F
WR7Y4wgZVJPNJWdBPertdyIeTYoZpOcRb/Dh64Bk9uOlk/mTcjJvW9r+xY7QAv3g
Z7ROqZi5wZ63nKVUl62qFVUOvJIyJ9OJ+Ew+8scbqmW/8EXtwyGFsxAeL3lHlhRw
VM6MJSxOTw6ssRQEUGxilWzQUxIYoD7UWJ6ZexeJl7y4aLZrulIARgJNZdW+iMsM
B3I65ly0QU1Ewiy3whlDOy0kd8z7uCLMDneEKA0wH+S4uv7Da6kG+fcImOdOawDv
n0cQxOmyq+BZUVPjtox4uP5/Z3Syto4noKRXxXde8RTuawjLN8TBrPEc9/fN23gF
TDz3XeXZkDByuiR7hjI6ReSErcLnNZsK6Ql7fJxU8wXcSm4qF1RIBmp+h9dlnVSq
M/BqVtVbDX8Y7ZkSS644TqSI4NeZuM1rsJaPQWtI1snryhPRyJ6/fy4iDBSmvk/J
IFEW79sQnapXdUnDlGbnLqNRKdl6PncY2l6oKIExbshU3O2w4L06q+Bf2ZxD2O0z
k5QzkKiGOnAWawlmBdnpcYix5dE/DGFEAcorITuWBfQVaoUz8ejUdjdTSv/QltxS
/HczQIEz74F4cmM1/ZyoJE03Z3Eo0ALS5VthjHvWCNaC0MvX92m5aWJVQtHF/MR3
jvpZ5VkQCCssHZ/Pry7HCu15LXo9/KiNV6zR7y6c8BvQWQsnqjM4ZLaTWjuBG+vo
MVBGHy6BadxM4Sm1WZ3UTANvGWZYdJ8P816MCJ48JJwUun/9kbALCrludEaf8gk3
su8FoizJRI8FVMBzYC59LhoJgpUNzPjEtY9BHc2KaVZ4BR/MKIoXzmCP4//ZaoT7
oigBqntQiAKvP85AfUEifpqL8+c0E8R5KRe15ON1pyPnQau/EZrAsF4wSC3FcCc6
nCDtjRsxOSqmJjfCEAfj65D6fY9jDPD8zeJKqjoRzFEpNYecbGlg248iqmeIh5Q/
g4h8fCJlwz5qUFafBww+hm/RN2o5UanLRoMRm4CzccrXsTTOekeGfuTO8QHeHTmH
j2lKgNdR5SYwK7oGRA87Lr69qnPQovHGfTO/EDzNSltFSm7NiIGrzJMD+kDi2CXI
lAtRawJbP1ebF38sDMUP3G3gOIDcPxFHnKdMhr0Yimz7jTpxVdeKeVtVv5Vt+6Xo
slnbWZk7WT5ISGGQmaf76cUmZj+wMUWJKVpYvxv+bTWzwG2MntbHyZm5oVz15LaA
XVAQ2WjcMUx3kQMN2eW2aVEi8OAjQwHSeY2dduS7rx6aDjX/JCTxZvg71hK4g12i
ssirnPoLSCxWBUWspXigtM5w87s9YX6+G9S1OLetSnQKVKD5I7l7p1WuxP3oCDe4
Hq0js6xhAQJGgr7Fr/nD1t0qpHND7WuKdE0mXpvAOwTgKBpeqA5uHsH9B+C/xD6G
fIVPmAZjpX0KNw81GWoHQGWBEZGQEjVnbi5iowuPuIJ0siE/9qoO8PQLTVOVgv72
LHrjPjP7vfGa7rvx04IyLIpMbRvs+CV9T3hEfZS3Bf5GNofChJ0X6AHkYYqTEq/U
CPmouqKC5OPWZok2zKtdQMxZCyLmjqemXVSyp91V8D/HUDp+SXKnTh500ucQJqt7
gvBGIyzl9+9UJF4x5N7rOyMBhCieGLIliCEb6XpBrc8nCwUcInUzRYQvYuE+smlJ
BxwFrTdiiWAlhSigMnrGQcSY8gDSUqtfB9CMgtw5aQbKeVM0oA/cCi+p8BJraPHb
q7vHpgWwNorAgCxlmbHGk/wcHfBnQRJpPclhnmSVtG6TWs29w8OecSNBWvYMoLcH
et7OqUucLcndzcZvg1/K6s08ux+69qDcmiazijvVKNq3B3RiP68kjlahoXIZkO2F
30HltDNCSHdfyn8A/BmRJ6K4st6mKBvpxkbfDevV2cew2lv2gI2aec4svg8ch1y7
R8FdymrMcGoU2FwEPmQnPm9F+ZlSAz8C1+uCB6/KqMpeo0W9dOqfc5sjEGceD9aj
4LOEuFfwXkhcuaxz7sx1HHpXJU9sfmmUuNVjx/+sr/WwQ5p8861MMOcA8CqkIUJ5
28WPnvWO5/tl1yiUZPa9V6cgRfQL9Oq3FfHQ0kRrWweOQbWGW5dmHxGV9EsB3EAX
7V/ZJjDm1YaJQhoNccHX07rqhp9bcpTE1AFXv2U9d9qxwsEhhBil1FZmwUhUSrRd
NcFTQbRyswn4BkC46latgL+P6C2lcSFno08vOmO9/MOaRqM3pBElvWkwB+P+cX2P
u6Lekw8JCOAWc3kowQNgg/mPYepquAQrqEyE2Ydy0nx1q4qv4raVcEprvHNNfanq
zkZbXk8HnmwW+ML6XLgqEF5ZoerYkkdPzAHTlzblphqt1Hl+NnaHTY4xN+PYuavO
RZTdzTZjj94cJjBAlLL6l9+el8ikx/U53HMcn3lSLxXaVh9kSrXtYzmozYOimxSQ
xafOrWaTHUhOtwNF3ppOzyFSVB61BTv9ArvB5nvuEwOaPviLVbT7q2tQ1kJGeawV
3bwFAazq1/+CPFoYqob1HB6PTOADKGMuc8/Z07iMji1QMwvsmk7jAhnCRJE7l20E
t31LPVHjzSDSrpkcGplAANZhU50WCsNHMdMMJ8SVj2XBkN0udNgX2Kno3n/cfSWb
He0PtfqIFRbkqlkvK6pVFXojefJ0Q5NWbr7h5wM1uKPItfxj8e0KyI7N+qm8my6O
cOgtePd8yy+Ozu1cMAakyy5yCauX4H2XNhgZXzYsZoCuap7z8nZUStMtE1xr1wpf
I8zK8Df5v+ffscfy4HJyWYiD565J5G283W0nOUTqg6nIpv3gI5AlPBTTsQaKhy5S
lXcAbMOUEvNztGeYvsub98oSIs3h90quXNW0sELSkkkNp677dPSifWMZVgU+RhJC
+lhL8kXYVYtkK8+uaPnqwUGoxcWz9V5CQBD/VeX0eGOI+7vfs74xKIoat3FPIUa0
Np/LDWtkVcfPvpeCmQhJWsLbdAZEY9Ey6j/s4l0O5hZuM9EJRj6lH4LQ389p15qs
H1ESCY8mp1cOO8Ek7fT/9id+uTlUYyxi/x7fQZjoGMtLbIYw6I7f2SaGz+p3BGNY
DQtr81BRGQJqez14UYQb3ycTlNBDminE4vTrpfH2sXaFxEp92PmkDh6TVMjhG4cJ
zdlGok1J2m5Gt/Tnh1eY4z8Wpzmq9SGJIaXLWUguqwDrNhIKDZjHLGtcB1kRlV4a
tVNEDHmEF3yh2JasXeBraeerXm2Xdg3puRINEDy80UyLcr5rNdwvpBHmhRjNYuCt
9++dW5+LqCSQ09IStjiLdFlv0ib88b5nMCeKtcwM7Xv+KjBJP7LRgSM3KHV5tMfc
LeJ1T/DNHmRIq+Ee+tMsQKysJi+YQUCaqH/CAMARV1dQI36gqN0sMY97GTdXOOnr
VEf6Ng8jRAYxna+ofz/FUd+YgiQjj1KeTQ38hCmNS76KmjpivtO3fp1FgZbN1ei/
h7ngcDajlTaAMHn3qGj6S7as9+mxcqrsz0eqbePAA9ducDhbfa3Vt35dYkdjGPog
lxyvSu4DY8U7AKQmcCMJPlpV89hs2QRFEMYAJtxk2JMofp9/RpaDze5YownmmwKV
Hc1J78j4/IXv4UBUXaUcp0Jr7RwTjVdQdTIkLtQ8rJ23OVp5PQdVI0iUF1GB1DQC
B5s3NWY2bih09e6iUl66sCyRys2imMcJy1IgVzMSU0/ShJbsvStuuWipd+sYIwLb
sNLkms6y+oO3+GHeuxIBJPzNaS5grM4qL0j8RjFzStc0XMpjjNRrwRBstqKFpO4C
ycxbGAtUyGu7pZmqgam9eDWC+jC9FmFWxmalFXE0CaOJyCsHzes0ZVl/a9qAHVa9
5EoXicWqHcm+0sTOSH1mKWHhmuA8x3CxTxeuburgWsxYrZOpWHbPNxpz8pAVewKA
5gIX/qHjhBF9lDt8m68kyfaI8EWVnMrZiXnVtozoMFS42REnoqCkicZ5E+bpv8w1
8D6svdPbbNHyKe/gAwwCLZx2FU94H2/2jo0wwnvpz/kUWiTuwfTaXe1m2d4fbVYI
NWQp80s2/YyBnTBd9affXjrF5GopDe4KXy9mEEt1tFlG+OVstL9RHfWZ9gbKROKR
1S/82+M1tq62Ru8/kIYpqIS7gy0XbQZ4VerqI0ie5H+TRlaTh6Np5f6x5f2KXAk0
wxjBzv8hBCqaQc/vlVouTKtcSTPiLB1ltzZmVTyqdtUT3NOl7vLSMKjoKe21mAEr
Zf73GpmEQB3+c7muCa2KO1KXFVUmKthZLzdC8mHHUl9OCrQQZN9nPmlApBLzF8Rs
mo4Io/yiX3Qqkc4pALmBeyq8b3wiusIFBEZzR5YjFfGqBHgjNpNi3gT/doI8nIyp
TS071jToO+5uZJqmGdMZ+4IvlapJwmy2fqiSazGCRB0QhkAf+tzQhDPeG/Ycdh/m
GFQ/uorDmF6pJIrroU2N4a5G1FipAbnn0jZ7I+UzfkeC5LRkSOiZADD+PHcBUDFb
41wdyWMLGL5JLktDlz2cF00En7d34boOU7tmcFhZnmGzDPnKo90v1pf6lzyhFu5G
LGNQNmWtiWEctt5ScKlfU9LXLHPY+/UKSDoCqekBKxBvWIwLrhSIySHj8CbsGy3j
lw9Pl9I0pUpwx9+Yu8NG+mKuKl0OE7LWCprsNmPbyJqfyGw7OUe7DAT1wXtdHh0o
PMmjWtxjK0ltEOd5cPTv2bQkbCn7pyigBZd2xia7BaXfF597kFdqKfbqaJIqzGnU
85XKOupfK92Qs1LiMDB87QDmrMuuiUDm/mnrdQT/6PZ/wr1iJwSr8R4py5P6hViG
/kEGshj4utuOv60F9MT+VwYd+a78K4YxpeupGG8yKC9FTpADlM6pSAJ/kqGA0ILO
NW2vPtT2QUaNBWKzF6O0L5ujQZdszWNlZLMlM1Nnmh9dfCcvjrYUGsMRaLAjMpb4
sX9HubcIOdu0NgOeQMdvG+KUDxskysxB1Y6Gtu5CctG75ICDg0vCwMVl9BgjNRww
iy6pXk8EpRUE8J6c7B9RcYxEKDduWmYCdU1KYshSlR4QTMiOd86e+p2X+iSt3GQY
t76dfncOZIFE7jsOWLoCSm3ga8U/7JTemDaDtC02Zo/KzXo22kLGipUmjkWfGusj
nX001C8euKXgHRhGw8hfvT+z+UEGMsbc+zIbtGyh6yeEdSkKxQiyrQESfdjodwnz
uGkKxyMwj2XNCVZPcJ0DSblPgclwSX/ENOcwiKlzoTrUSs9Ifw2NwuenHRkZPZzS
9s1EYUsnL4AQ1hstGVgwMaTEULu5fYV9MDuGwW1PSy4n0yDEGb/f5yAR0d9Ra3Mp
pW8pEWzBrMtfOpi6Otzsh6K7TlaxjXCqsB2/SMfa7YL2lumUhvGtSlepFq1hXYyH
L10WMJZ1/C9HvTPvg+VM9oNfJllIg9NnoZsWALC2p4KlkrJ+x8zwzCcg/qdYbvbX
ZlhYQiWJd2RRRkeARISJRA0RQJvvMrANxOfdS1W0clHmMNb3PzYxUzh2znYc6En0
5Evl/YltyUdMfg6cOHAkxQ6Zh5jdkxm8EqLJIEpGuKA/AwfmZ0tl+L1VEGEsvrWU
kwE09AMFpTeZUyRDnX/1bIPPBz3oC978oIas/1sMwOp1aA+K6mhFgs0T8H8A6Inp
wYQA0cFpDxyWgsjdzUH/ZjWGeUYPb5Cw/QiUmZHSMPeiDQdNagutr1cgDAQuqmpW
GwGYaLVFhPGDdtjRiu9DM8oCKIIM20Yocz4TodxXr96NXqu1IQgv260NQsMB6+Mv
AjNuNK6oGiecL8KsFfhTeuqmjB86NLaGkLQwKFi0z51pTeHddTTzbT6yRLO+/+bX
p2JreIxSmOSgihyaB2kkWRrt8C6Ohbykc85AdDegv6QQajH4M10CoGUwZNG3TKKA
40XAijSJnKdEkkvoulzjjWxH6BmHykNjiosFuHdeyMCOUGM6jpK9BHlbCq+AqZTw
yIfMg6LFi+UPCoEU8g5EhC2Zgk45A8XfkeZPfa+KrMrTJRZ5IzvIbAyaDPIhkFn2
BuROeq25Z7hBDi+RndXdG3/hezpZ0ucyu+s5B9BOc1MMPvKxOMA8q+SKIp7BAnlm
2KuHGos5CXHvKgUcxpNgUYBT5+jwEjBk+cv2dr8nB4xRN6+0/CqRhhdtCDDfDgsA
O3s/DIE5b5vkj/vYoXo8+rs5g2EZ9xSWD8YCgVhw2HqQ4RiQFyslOBK9SeEe6Tlz
OpDaFR57sPYLHCOzZ6KYfK+4PSB/bnkmJG/kER1eWrEqW5LdGcj7+mf0fzGolPo2
Kmh+U543MWdy4spzwkdukRSNhy12MtnGyVfo0ilocOizAVppphayeKofd9T1okGx
hbT69VOs2tUWxA8sEAu5XfWA949Ei3xopFlTxy1p+59J5GK+uTV5NJoWlaQOq2Ip
UDDG6L9Kw5xKlRswS7qTwOVHo7ON1QafgAqVo6i186BHDHeYCfZlgz2JQutUP4lY
v59jUcvgW3aqUCH3Ibj+bLSn1jxO/QH+ijlDeuLG3J67Sc5f5lKH1O+sMYgNTrT3
bZ9k+9U850XmFmBiLCotRd1S4xI4if0jwHsQHdemmPoSQZjcphCFFsJQx3Im4URG
XsLKWnK2c8oaKzc1EouRF/2CV+Oielib84Wl92uYqooqxzodm4lXmdHpfWby+m5g
rlpEvBhb+J1eZonbxeEUprCQdCK++yGRXpoC6tV/O8z7uDoeC/ghilE24ZfjmSzg
jVilbFmt5ej9CYvDo+gCQIBDcyuA3uvbLt8ixaYLMQiAQzqNajZSuI/RjukHHJqb
U6PUUK32aGuancgyKZXpxdOp5OZN90BW56nJE29Dt0RtaUyxU427KDtAgHdZHc7O
6Moqmv1HhhxJb4Al0ZjCdamFzpgRfv1GZpnZ6ZpYA9TbvAWmQ3EoXI2mShts8Agj
0CQe1S25PikUm/m0DMYqNGBbswb6paIKA14oGrVira17J2doJ98Byo+qX5Z9PY9T
O2mo7DYcaBh1EESm2Zs2WbxVhXD0oG569dV/GxqZZPdDjqboEWqn3iNqpEjk+3/M
1aeTeM1s64aQxYbWprzYrHDxG/wJgncMgb0JPFNNjMLU93iulTfOlLyOx6tkBLlp
N+BopWkI9uQ1w8zPNPd3v+chIdgth2n4ccciDhWeNBY3bjFzFCSZxd9QSg4oTxjz
8ZFiH0mW0Da3H2xa6afyO+9sXLgO2lGmHfFkYEOe43lsIQYY5xywFHKl+sIxfDtL
zKmbhuIJeTGwBy31JwpvQq+BqBpB30Rt8mvGGlXK462O5bbZW+KiyBoW+kj22MaF
wQgJtEbZDFJjUec6lC2CGX+oDT7K2nmkL9Y9+/NvxcpktA3oymgMM78NvUW7gG06
mzeYNm7rNi02GEtFbdAeiSAfuquTzOqofOHHeYpK0uh1Zbr6YtDE5nS04qnQ9G16
iprBwtowMZBuIYzz8IH9q4aXW39NqH71ZoQk4TFsVmnhdhwR3OUWtgENCUzI9+4c
V63/MmN4QZqeDiC/ZmxyeeEc7RhXn50N/rQy3feTCjvc6XKV5gzuyujIcK+zMazv
0cagnP/TwgAfmxhb7eVFoKm2LWOik4wQ+sX+0s3dixvm1bQROxNiq/+kbmyNQih7
75Cc+Frv6q2TBJ1Qbwpzfp8gG+PFZd5UaA8ZnFYP/GYqpvSrpSbnQ64zSYEB1If5
Fleao+RZMVLUKU/kpc3XnaROAFYHPpzCC1MK/xoG8deG1QiQQB/H8J6gngxk4v42
MbCnH6nsV/MIzm/qSZqaVFLdXoAbIFnK6Ht+bn6xER93eab3dJLTpofC1pFR29c+
hrzx0nncbLrKFFjFHamBa7MkIEqlhj1BAO5coqagiCrrvcDCS5MyVnGPNb3QF3vD
DUfvG5LqIjns94n4d1H/aRmwNW9AOFfZCIncPbeOEV6bVqRot6PSwM5g5jM8HgG9
Bdy+7bDr22WnTuwj2OQyqEPktQfaqrlmdb6zezBWL4/kZlXqGKqKX9lvkVcSC8oM
g3CLqKgBrghqYv6kZIVR50K8/GhgWBz9s+/oEJeXLU7Zgzg8JM5RUGmVEZJBIfED
AImtZqMEuvizd2zIG5Empt5CrkRuKgdNQjt5BtGmOkpp2mSCSa/4U099L12D0wxb
mWmvW+V1z0RcoHBDexps6Cq0OuVMkta3UJosbehm+eCOmXgdvzMHp8q2/pyEmfuf
OhZAQpAgbpdpjhz8uH070bPjofjRmQaoBpmQixCRbZQzF2QlLh01GMCWCfU9MN2+
yN+W8H+DY+5sHJisznqbEFtlkclIE1r7MsMHkxZDOvgzgfzLfPPE6FVcXuYr37iA
GlmBeyakxL3zGl+MqPt6cCBtpl1C+xWObJPM50AgNrx9TkmeehVG25pOV17LHK4w
ZqT5x5bDMtIDZlNuDtpOhyA01/cmyLq7cwvSOELq9C0lNArbYF3Q6iXIobh/Rtgo
wCawyZqJeC8GCaW96OEVLhpa5wHk+UevxfrqQS2wr3Y5KM1AKlz0IF8BLnNlKa40
5TLeBtNH1aZwfrsyqmnFr1ranOot/IDjcQA8FqKdQd4EwukKbnMK2Ae7tcuypzm/
gzpn4Yeqiz9nlbQjKCQE0+ESOTr3YOk51p/eMDKfqfDY9cn12EmvMgY0FhlGAk9f
GbEG74HheN7lVY51fqt4FOJDjjxPxLZx0cZDeRlP5Es6WBe3L5HFhNftBSS9pHQO
sIlFInhvVnMbo6gAtnYYQbEQxMeUXEY3b5SEqU8J3EPppTie1LHE8W3Bmnst/vI/
b5WUNQW5+gEbJGjsBOYLgNocQwGr0kRnnKRwcbe6Lq7nUr0Bm9Xqny/MqE6KNngI
yr60te2MCMPo6lSGAblIY3DOXN1AYa7IRk0eJ4P4z4HgolvtXIYSHoVLv5XAhKSN
oFnzLHGH1RGDlB4Mb63Eo5MCOUOmEiYJNzb4zpfcWYtsGyD5QFRfEuKqJIWFdKFJ
oFGI33lzKcnpjfkZ0w96wvLQOT0zrGz3YPW0Bz1rr+HPlvnQjk7zW3zYQcltA0nJ
Tn+PRFDQopk3lsXysx4sKshdexVGx1Xzt1sLkh/9OH8NXAQtiacI6L4FUcj5JLBq
T860bdcE4QhBiyvfk4ClRgWdL96uxGo9DikYUDgeJEmnL1eIsMlHNaKoalDCEPnb
k/AmxOu7WGQzMTYvPRMliwA0ba5RJZADJzz/Bkazud/v9iVNQjRat2TIzOu2kldh
4M94ItD7jYvV9ju6Rt+yMNGqd7rE6OjV/lFwSK0yiI8FKslJuK+095jk1TYUwED1
tZPEfup5/OHaxexXATEDIuXYP1H91Dxn7HBleoYC9EqwZ5mykiAjUIaFwHmLdyyS
C/DTOVk0uRU1UDQSn0kvAbSamCdWw+hmoMi1lxlw5vU3qtYS1V27JQ62RhLmMIMS
/a10s56DhFEcdKwnMbLIRJTNZgjLd2O6pRqkAfFCiAZM0EVOIwxhQY+Hj1g7v7tB
662Jzik7/mgSE8sIO3zG/uG2z9XiHUszM6iRMRw+j0PtahUlQTIZBYnxzqFnbNv1
tVYBblNtD0FC7jPiy+3ftm5RoHapVlahx6N/4OOt7YfpKD03Tjy516sVbmbWUXO+
nGUxmbC9LgwelNnVSYE08pIsyjTO+MlCvwTV86raTF+4odDUzf0DKQswKHXXQHz1
WTkW1LIUvRvjOQ5q1eLuLXP+9YoP8q68B6T35WnavsYfwA9Qcz9TSkZdmznImaYY
MIr9jGmnILYUAXSopKjrokx/BlNlNF2+oFUO+8AcOp0Xy4bdX/As3zQ7F8YZNOa4
w5SnXGGvyLvlYA9QthaIeJlLUJSSG5Acon9/pyFGsKsXBtoDN+IecEDFcCoRx395
NhkKSKxxs5XBNlTGusqcnZh54nU+HSOHu1PKLgfFNi8YIlqLv+N2ypDW+645wqZ8
IQZySIQx8EV2BSw0JR4ofo12kKhR2MvsPwV6qixH7g43e3xnQ7nOGL5/6XnZiDfL
tktCcB+sNGC9kUL+zN+fk3LsYiJemoXzDEP4sYZec87e/GNOlfOF9Rl3yNoUHb+B
MIsoJboqm+OzA7SGEH0chcuegRwrthTYslpIg8+4C3q2OGfGf6C8y7c0d1oOFNsM
houw7pfN0YkNNkL8KnY3YPoCb6VN+Xl6t4avWiy1ZUY0DeEwmNuABhJQ/FOyJq/t
qOdoXkO6GiZ9FRmC/ldZ51PHWwUKeJZvgU+3pw0f3MmgwZCK7eXgSLI1rZIoRMEH
4LiLn84FhsRlV8ThwxljOcjBq2Ti5vIvdLzhTBZrD4gJNnj+uDwGCB7NySkYMFPo
mr2zaGl2zUSwqZlbSAmhvv842Ccc8t4Qul6r34ss2OhRMbpcKODN882F+4Pc3F1k
jLMDCFcF8VdTZZm80Ud4Bus5MEChP/1IigfmyuCCfSQh3NdVI0xCd4m6FE4eRTli
8O7G/cDcEop8nwjbBKZd5LiIoDylUxJxlJWABxobXb7MtvNcmLbKiDaSreokqFfR
KgdtAjrouwZ3a5Ti3zfR+KxcpO3bXysMZKANlw5xzfHxBDa6TR24x9MJHsgVM2Zd
TtsTM+CeCkTwWiNKk/hLEsG792Chh4dbf5glDGuJA/b5CntLJFU58ifrEQtPB0V+
P5Ol0vDFVJ8q5I5yZcTmCdRJ3wwjiWAYAS58EsU75karHYV1VSpSwlQoaUoBT9AJ
bCQsuoNIH4r2ScNkmc4Y+t6Vpk77KdU9qfs2m5Ss8MR6+Bptlk3OasnLvgjcwhAZ
LpmJaPu1hHUmpmyt4eiQYDlkZ5e34XaZMOnJTY0rqGl+ARXgGrDpXnLov88Hx4hp
gkYD6GTmva3f8j4Pfgnc1rZ9E/Bw77/gVsvJqlOAbslR7L7g9qrjvYeALfIl3fr4
B1i5EyL4KdIqsi1dEj0MiknpO1CTmqMMJVRKABT4pQXGfVKZXaw35iGTGGplwgIL
hrxWFSzQFs+DqaeY/Aroo/JczFwh9SohnckCT2FrqZwFnPZIHcNMZ7ec33bmidHn
dLgLnCTniI+gLSj16GuKhS2WPc956lzqPAnjH8uCMLBlV0JAD4vxB4tfCp4NwTG0
bm7B3xzwYwcjdoJDOTbpAljW6hfwMuuCCsE/VVyZoBITCrLvx/wCO0lqaMt7M+36
7HVO5vlxeJNxC9FpmfJvx2CJgJXBo2VPPt+GpS4ZGzEg0A2SX/+kUMO7K7R6kBk2
gATuCrpRTMUqFORIKNAkXX3ug+ihnkpaLkg6Fk60vlOUg+XIjNDf/J8ghWu10YtU
KtV6DQT3ur6lxTRVySyCkCZ0smxpR5HMgRNhwNrPXc/TEsIzf4hLxwJbKeMBZDvF
6pmR/RKTIrDEf2rdzvYP90uS6eeDpnwcRZ6jTjqKpR5rfCdLi7bPN0Pi4hPM9b7I
Uyp2zwa+geJVoG/j0/rXHApLM5WmDnfL7b9fndijQFU6cZ6YuyXiITouAClKzLPR
e3TE//Wy7JHsZ0k/XcqKFPzGW1JVc5AxBt0rjJdeop8J4Db0yN+0x5q1fGOtJAdT
yCBHIKW4lLsGiEJeUYeUS8vjp3FVZW/0+I1vwcuUjC8N9ugaYrORxkAbBep2B2G0
E/ifGOz36sWhjcaRMpa2i/4UWs31cAxhX9erpBcs33bD7AYO32cgH5zk6mXiAELf
0NU4dDg6EZ408LxKaFkjzcpXmK23wtX9y3n1fAgEQk2fjK1DRJbTAqj1NvhSmp+i
gSqGsMvcWvGvO8qNSvS2gZCNQaPlT/qq6JNFVAXqQ4et9NywE7ksWLnsosjL4x24
Kf1hjVDom+lKPmBRel3fR36UzExEL06DO3ho7SiuHrXSCxqBaATBTAfT3YfkRo9e
zxHEnjCWkrZhcPvQTvglVybnkcQAqzDDlXW2ydLlp+9XrSPRDP82PA74nNFJZtTl
lpq+FTVLyHtsM1xJiOXoyLoe0TCxxwaItLD7t8QYJcPHql5hl1HHh3Te/3oSpYrV
zdDoxo/bNuEOjSbECYxkOJYXL9G5NmFXn7zpTdT5is29UDkB4ZyyYEk2JRMtxf9a
LgdZwfVvcTuy23dqHpM1d+GfD8YjNhXrVcPk0vYeYvZVwH5RHywMavNzHgfX/g0x
EwD1f7iZ2vf/fgSmXoHXXsZQdEeP4vrYxnwSZUAalfMryOrEt2KFWHH+p84Y0WGU
hk7TVb0h12sDrt5PiCMk2ztOJzBhG7AG2YOu/mSEzjjYBfDJ3EqzNxitCFfAZszl
8hh4y0peGWV1k40/Pl9ZtxICc+dBFLMgWICTapvEBO/XDIYODqvLyHB1wLaSxTST
4gCSMkOilGPMjvLvKatGlgyB01wfxGWSUt/NDVskKjzspSLZSHHslcUMRf9MRtoi
9rauxr0GwqZy73b+OIvLX36BIE0KJw821W3Y/3t/WKmOMBEg8SBN33gARu0XFi0N
g1LpKn15TX8YXkODF6jEI/Xj6un/AJCOyekih6IU7igVkav9Yuk1MLQeXjbl6PWF
xW0zoWmigK2xB+aGfLpb1g5cunvyED+TaV/zgsaSoiBMXmwEepWMX1DvIujA1RWq
i/xbGn1HsGphpViPSv6ejGnj3mrcGSSNKyHzQUpkG6B9427iWwwlfkSlTRjdbqC8
EYbXJD6px4K5CgoGgLLp80+4laiDDIBHSQnsBuv9s0lnr9S/qNBxBLqYOGHxQ0VJ
kg+hDlX40bGudDvVcbUnC8ayXkWcDpjqm2ALV+cynNAOcPQGXP539hzSXd8qLwDw
Ar5niYNX+34jnkGyfyhrE96o+suaH9lXb8Bo795pvloErzZHqTsBuaZG9m16JrJw
o1Kan4PloGEqpY+FnCoUKDO7j+dMmiRpcynZmlZQr3VDK9KU4kN0TzqAMzNfwOUW
6Ak0gPbuU39M7Wxv6FnSoXoiUhAkW5qNGacRO6I01gP8NV+5lnyGnFy57CoFmKGQ
y0JOkW8d//DrHXyKZSM5jVdKAl/f5MKqhX7RN5ZtQZADlvz9Xr7GHAxn47x5C8rd
5BbZbBH5UsGJtqcJnt0GjoLtOramUA81I88LGyGbNH2dPQ4Er8sHojQvqJHZJ2mi
VDa3oalpYHOnApSJTwyeb+lngTZ3vfltH52vgDPRXeH4dVnU3Fn9jlE+h9FgWOSs
EraunX3fxgx92dWy/rHYJHjm+tXxxv10xwA8sQ3nGSnm9h3Htsi+Hk/KL0vPfFA8
Y1TeMQl0iakYkViKsEAjIEBFrtepJTsJVzan+zk2WGQmOPIGIAplTJol2BZT3dcm
CthWBc1AVupQvIhx2prfyEdpY5WjIwIWoVtMF+ZhHSnf7TJrEVviCtbfpm9bcMqy
fsTh1jtiUa8poUo/DxFmtqwFf/SVlAErykuHGhAJDiLLHCJ9JP8H5vnhsgK51iLS
k7uPtdGwcX7YryphAPtJgOM+IdTb4GCyQxv1XjSJtb1CfGNPUoWzZLOgXBOYv4xa
al3bDdlbYJcfMVcR9vNJLmQ3n4uakP53XpOJe1gwctVx95P81Fv8Ed1EZPJNHwgc
3HAMRiF7rN3jgafGfrNTmHQOXbj5k4mpLAqEc7C7puWWhYA+9KYG09Agm+B1Ewjv
K1P6BksHxnhbkCrVpmblEpQevvwlgOV9zUJKMRM8tdCOIwWhFS2yrnh0J4Pz9da3
kuhr/QRScOxIirLGSjjCWgIhRp5nsAsuKELEKdqWGYIAQ534GjzKr8pks3r07J5F
lcA1GeD0JyWjPeKv9T2Stv9G8i8ClRr39Tobnfl1KXoFX68ToRawykepSdY1DF/P
bthuBJHcK593MiOJM570gZHvIwknul8p1PAPu7MOJnd2W8PGSGy+RARY73pH4Q3V
yQgW9nn+X3d3U/GT0Je4sIlmxrVMceP0Q2oFcIIv4n0kGnOXrRiHhBykffQM7Es3
Bio6oKnvelfeAoWk+/Usuc5Atqpw36jGO7BL0vgRMn0XwhEXqFpmO22xY08W+hqj
5YxInXldV4/ku3eoHNdeegrauAJRd3Nrf10WOtSDx3XTe86ACHpIxSuQJjEQtDh8
gwn7NGeRhzAWdqDatAtcMtgfDO77T+QZ+gJOv43Pb4ccvwSeqgwpcY7q84NNmqnx
GDHRBfRtj2wPCLsRdioTgOAEO+FM29xqhtNaTcGGZKkbLhqS2YPYc1YBzxcfXL1Q
k1dAmOjcQ+InwCirI62r8KmSRSOFCYRK/mjJ9c0wtnvAWnBSTTLYQoD8xMkUc7DT
1D0VzqGIMg2UupCHjgcU4hs2fEPiIzTJjF0N8HlEeFvPO/ktEcz4cjeLdthDqyuh
LJK8gs1gL9MPogxCnV73knH+uLYo7o52MRzKRlYSOQnnrKEbcOHrLl2kF9FLnu26
h2hKRaVVJvsrKvm0beMuA2vTXspdlYcy6zdsZbrFpenwb/5LYfCa1+eQfXpcVAsO
AFkHwqvHZFmqzqw9XjBY4vGo25WN4tYAGhQssIqjHSykQtpNvUeoalRwOW96H/Lv
kozjVS+3ABhAMJYQfsaYG47DnMa15ulOG3uG+GW0h/zqRPm2Bn909FkhJH+qSG+P
zuxLCz4EG60U5JvYhIyhuFN+1XzKexivZJSWGrYvjyI4YdckOSGyBGh6PR1zRClN
jgNs6Gmn9pL8NW3/cepJHKHU9nhLKI5pbm/A6UWGUMb4KiJcsMOL60gqeb/W5F5Z
nRe22hTUOtxJbstxpugVgV0ueOP51NOQ3lU9z8e+/eQu0UTYOdHXk+CJ3IGW+zfK
eMhpZWfLe3Pcn0DOGKsU5V9RnYXT7lHM9+A/yJ6J8eo8N2Z30v1FRnZS7JEiSCfv
76i1Lm/HlG5eRagTxSPoCqtWgHpWe+54ecEwmdHkKc3mMoFngufGG+wJIu4PljwM
fU3vMBaYT8BNwKgYWfABdwn/8GCrrXBsd/hiLy173GYsna+b+EvumXY7B8704j3K
8hpfGtxxSfNvXcomn+rArNTfJagXYsOXGkpm3mxt1xe2hQKYkG+tXTE7m1R0C6fs
7VbZyssNCBQrnFY++JTKrtWq/fruK4GOw9UB49cptnWzjNHJ4VK9MUeqFwNCt4kE
EMgZyQIGUBcN1nBvfubQbwrul6V2KNJ9T3oOcrMwwhzm73ssaLKck1m7VtgXoIrE
WjaqKHpJcR3W+K8CtxPyJ8IyCXNiU1+NH57BaoaEmuXRUgvKweAcMiETUGaPTHNj
bSpKcikEwtPqbNOUmjSrj8azaHWFojpJS4JkHeWOE8JylwdJQKGBibHaPOsYMyiQ
WQCZot8uN6/moCV4OQ/FPabVFNbYjUt1GnMCO9C33T9TNtufZFS1AdmreliU0zGL
VNwjGVPGMrzpR+gg4bMheC7GuFJ6JAqxFvcnq6Q9kOZivBaUiozEKI/QhhR75War
jmVUYM7CIPGHwMhNinadNNMTXBqcnpPAuRrBFfCOI88DJugsf9cdUdD20cEZ9qXh
jmdDxS/f93gDRas5KyhwAMZaJzLbSeiAMuC+2CaWpHGoV7iIbSrJR5CtbqpHnuwO
jfITwvvGB5xAWraBD+eUK4jeSha3kZZyd5kIP7rRXSuUDRRFVbrKMrliP8upUh0k
O1erw1NPuAF0fF32YL6HlL8vSAduI3N07watnJcJHnQFbx34RuEhMmQsCidDwMyC
u0mluBOPP6peKlz7i3Gg33K8prF2tTBPCxlQQ4hB8vScyKXXcLsCqvzM9piOcfab
/QTkDCyRYlkqp0HOUUac8LC/y6nSRuU2TN9RVSwAujht9BFmVaXvRSvDLdUlMQmg
NZF3SKDNx3CAYsZ6yEuzH+ClpxsDgu9hAioh4ZmWcpXYTcw9VLaXTQC24pNwpiGz
9Q5v+rQPlNQX4FvaPcRct8c/UTzrphtJ+QlWYPIgOzn50zJliHUcxl1OeKmtMwZW
LUPiDs6BSAaMjXJwg3zaZFhXu+w2QUJEpLnoJVB3u1sYdtnczstVU63vNjRao9P/
fx9jagEYEEnyumK4AIcoYZmTKdaPEJj58RwW4+jDQ3/qfDRkeYgk/S9sU74ukJCX
2FCGLgciILWT3dWMbN3urtbpnULp8eHATOgbgYAf4b/H/C6qPu34kVdmv1kJ03Cj
QkuZnnGuyayiy2AMsMjZbop5E9j5pLLIkNOfonB5OUSVAbitkUCuYlx/I4Ux+CCo
rV73+HOfQ/00K4Eugtdo2crSDgPA0uyUyebavi+0R0a/4Ja9SJeA7IqBf/WAx5iP
3of2/zdSLMlC6ZTq6+yh7AVjCo55MPfsk1u0S0LxB9b34Mx6XsZ9gBQL+Gg8Cwjq
AqvXa4Wx/AqKw1LwJZaN+Ud2ovcrLVv7BdC2zc+khywEI+Uk1D/5xC2JX2zdJHcP
P1MN+kqDuM7Dodjz6aMP4EL+/wvKevFOkWsMYlfA6XIVqiNYmEtW/RA3k0zuEuJv
+smmVn/giRYWc9/MULsT6zsDrGhSelK6M4WqV7v/miL7ZBTzJYQ7FZpDZSvJz2cj
nuVRLueMptLqFwdmOJLhgb7EFqQjXHNX4FWTot2wGGMVaRxGpwRSXngGPnNkVdfs
LnJpuYzRexwmUmkeSaEA7H0CYZYPVwraD8tJkwG3yI43cMVG2BYeY3E1e9zXKxvn
pyQ05E9evNNYMZIHO/Exl7iuOyCSFIsu7i4U3TnZth/nGfvOXAKE+MSivxF1Udk2
ne0qAxrwyldnop97pmRsIc+y5kMWzZa0prezMaBOkHVH3Bt8nNwttJnQIZ3SK2Th
H0VSGnzje8YOE+JGZGRk1Hhn0WoxbZyHzehmLNmAByI26jpw8hA3t53Q6D6cgCu3
paISbj7/YVIJ7hEkI8qT9QSBLgD2hvTcBSVCGRHrsmsCxqavQKH7/XdSNhwTORSZ
Ru1Zfhc87dQpTGb3cIIg9Jf9ObCunwfQdUl27hpkEbVVxvQZH4bLdUuMbR4Vzte0
R7aUvk4el2VMv9muxZ2jVY/LGrzMZa9643hTBCmafYbWkoPPMfm5RSnTXVWgdfoe
zD+wlC5b1wkUpHiYTNsV13PMrLeB84udToOh9IVuodvv2vumbwOFHVLO3ybsgpyA
mLeUwnVM2GyZuPxlFYhoXO01LjxwHrjG3GTd/Im3kU9/4f3VUtN0ylD2lJqLXFP5
nq28bBOJutlUFFXWILrjM5Znohcw/HAVt0YkWs49yqveUTZ3SDB3nUz35A7NasI5
HtiWtTabik8hmfYtcmgAE0vn4PHSObXO4IHJwZak9qB3djjg0/FqhIU01Ia/352T
TPRJo5nKbokg56UCN4V8jB6ClUFxLBrwU4vHhj35ecx0pGZQbKz72gO9VoDRvlxx
QL2fpKjF9d+n6Edp1c958IXZpIMJ/BHZbdmbMqQECqFDXiwQDNw6WWAD7uefS8nM
y9ee5+rQN51PtYQj5HxBUXnfIdLF6bSE4M2fD8pEJhR3Jr80mYNymNbkN4TsA+GE
6r3wCfm+arPP9hZGzK3z86ai2DfM059PQQ/juO4w7thuM1QaOWkI6QH95tsuHhwW
+Xr7XvX142cH3woavKxN1NUGSoQP+favdkuo7Vgb+IvahAIWWvECaVn5nNQ3WsZh
4aL6p449fWowoSH0zk2CemnTDcD1K1ne2V1ULvHYn1EgrKmgyuWOyBCRMbEe7NcA
I9s+oOK7Ghot1s9MB/SxHQHIuW2KL0pYlzaDTMZ+eqIxoZBiuKvzJC6hvxUGDFFK
OXt+1bQowjQxisxAZlrAeE7qRxbFJHLSr0kmyw8da6MCkvZOCUXcsPffiuLgsWEg
5iAqzoUXEaY0gBfFe5VL0Q3OxW5Evvyl1UgMFAbhyP0tCVfu8JG9lMmh3SEwhOjA
4syBN5wLTLlTKTgCjh9mWEQcCtbAWdjiSXtb/f4TgLnWDNzxbc1fltXx86DPEoEe
PVpLTrvgULLmBbYkzzu7MD5K+BExsfBtbu7hTpYnhz4nw52pdYFJAQa1JSQ1OJam
sgPaKS/7ZaXnjtN34Uasnc9llZLCEfvLZ47DhpLYH45rehOqQ3z6qIew8wevd/Wa
QdnpLfDfObI3TYdOl7DFesujUzVKxMLFxFAI7lz77+nuKO58uDK8czDN+5ev96zb
AT9KrVlmnGbjrUO71Lrl7x3sv3hufXx8qVTRBznC4FCRFIau5iNfgB0vcOtzBw+1
NsO8haYfGBqPvtxcFIDlISO00+WdAOd4QtVXuhXOupKkc0/+UwedPhUXQJeEOXfV
AdZjdAJpTFOd0iwDOVysuhyHF+SPfFnXLrqLZIZJ7oJYJvpiKvpzVChNObVzxobP
iL7tFxTTMAZ30brC4SpTGRuV2Il/+Fe15r2y8ar3ioBAgQQMjGL8ALmtWF8t+Fc1
DZOtdDCdXOHU/E6LIVz0kO4TPWl1DvbGQi6SuEypDN19mhL21QfGRdjrOi7xz+Iq
cWCGUAUy6BoONfCg0X6RoirmcPbIt6HzWcOSjjC9fND6iV8dpoC5lPcdR2onuIyA
6gUvkZozQ+HlCjuad9JpI8YHQ9E3aUr5o52Vzjnradw4i4JFnUEdtu6I72z2aJW9
ycTuZsAfuJiIvpQBVsYpSGn08P16h62/hcHxV56FCHJ5EcMD4VOX9vvSPgYq3PkT
XbQfcWqyxnUeSY8xggaIYy0cmVgd6hsqhwiGAlvpRj+zjYAY7720n/xEA5fhDIcF
hkA8AXG0b/PmeUT7kWHf1WOjGN7IXx32dUmdngJuSIj1yedjufn7oaDp2LGbg8H5
OhTpXIxUWVXPaDWUFD6yWeJhJwqXYgEdaKpdhb1LVTmczxkGSZoPJEWct1vd3dUj
ZJloctW7ZFW50u+g9Hjqf0g/WvMcks+uhXP0caTe0l2UUBgnWX74khP62VcR3osu
B9/1vU11YKC2u/rh9mQ0PvGEfF57qqy17wjLmWHfKBhujvcMk2dp4ZKYOglSmjoN
8pWPtJc1LO9xi9Cd09jQNSOJ5nL2y/sr9Ih3dkOUqYwE8wNMkSP/+RtZQFDgknrB
F4T8fy+qhYJOFrfLnRZxGJUQ8lzy06ptPuMhZ4ukCdj4bh67udnvvUVz8jxKlwyb
LAM77AxOQtzyMqzhJN4bIu4y+lCCH0B/7VqvAQqKw7DlhC9PImfLDPlSSl89E+q1
Qa33Xlu9jHcDdSucPQk1ud78+MANBQIpt/PXN6h7CfVRKgB8DCb/6JT5kFAWRnfa
cV3RWgntznWTkR4DRF3tVz34iAf/FFqbamrGLYrMxGcfIe38KnTH9/ySE84laxq2
zNpu235en0xvNaFwFUiCR9tYyGAQTURPRD9CLxhRpLpsx6uzCXrVdpM3HZ6sFN3Y
dinu46FUPL5kx1pSPve7uj+mFJDOUyFy1sPA/m8SPpPh6c2ORABL7UKl1NDrkBs1
T9MVpJvQGRE7K1Hk6unaF3OaUHSUoJAnxmL+h+ILiAkrJAJAhNJAuPJ+LLKGxWmu
CSAg+RzRP0t+625nhmh6BHikY7fdNl9V7pv8n0Go+YGAXd69uC2HdKiPbIEVJX9g
d37z2/zxsfYPnP/xRZ+w+IhORzIGbPySKX9dHNmi4ILxszloA5MVPM+pYJP1ND86
Epzf623dSGiga1NPh66QRH537BkxikVBaVE0fomg0f7+tYQS2iHSIAvVn7zfDGJd
qjy2Z5utCT1IRZg0oYfSYtaOGoG/QVSLfoxLJ1760GGMFENSLzk6Q83Z6m0suZwL
OC1yC7LJ7f9hfkc6ShVvoQKAIQB+Of5b68Rp6qTtoByQJgCpFbUPNCELqWoZULCC
0hk76k3xWJEIDECxCEVzyt5uQwv48/lbbDvhzIDgJgWczL1ECn6HYvDNsaajejsn
/WHSwy9rzySqY7TpZnpDYvLsUBQ0rguoJDynhbGGwWtGqqJfBFvkJjFALNNBbrzU
SdJSy1oI1TFLBgquJphY/QnmOuU9wTQZghfmRQJQx6d01D8YT2IjkBQ9vn4ZQ31z
lnFadqsTBaAIFpWl7NRJm8+wk9Cp2bnwFYP7Er3sSVo9nZubfXUihRlEu6JwBdBJ
OTmG9AQThx3tTYaBe3dSuGkhXGc09CFkpbr/wLxqGJ/TW2dntHyHmaGOshfPnrnE
OresBxGp0ixkp5N2YAvVlBCHiblV0vhWMDnZiUlJNyjjViNvV0TDdqUCJuoustC1
GijEElLlq5sbPPPTOyUDMbO41qFhtJdPw4JwST6Bp6KRQePHD72J3yqNLJ/z3wcu
Dt68QFKzWfKLsanHKrk9Lm0FYai/qVC45F6gsCv48giFhdbn+WpuG3Qi/rAsgZ9P
1MMCAM7tGO1UIU/Tn6t8V1NxbdFDVbM7fPswZiQsK2dUaT158vvtku0D1q3JD0fy
L7x43Da/PitognSpJ/UXqFON0GFx1dB/l5WKadcDUkdjdpAU6kDjQxGoLNlyuVhh
UPUszlftHxJT9tfnBDt82JYn0rCjClpV9TSioLpHTUWbyAtp6VG1wvWXbtJcERPB
6xjQHiXulZpuLECSn193OgntfhJSi+3gqED1vOn5a1BSGOXMXpEMHJJ5MpYVllrT
yntJMPF7oakhE7xXh4+ar28YwarJia1ckY3ncAVn0rBoXPms9YTm/e83+6PMMv4h
gBgRmwpg3g9N87SL0YrELD0Y5ot7OHAXL5xxvwtLgLJBtWkvn8Y1l+qr77gHNvgu
pL5RNdn+vVwNWP7DlLA+jfmeyzS+v1fwkpWYZ4ySz1AhsqPo9eLJPSGnehrcHuMb
l7Y22TprBn/Td2RxhCOAG/Xm9gSj9t+IkF1uB/6OdRZQiknyVju0xTHg1SqFJ6r7
n6nNuRtj5186V0NPuYN1B6eJMJQVg/QeWsp1XVOWKL6/tj9stnbHwQnTbfJXk8We
aGKyyAmokk27u0HymBPtw52gVfsPL7iVmQbB+7317ln30LPDqnRneo8PUM7pB7nM
l517Pu4A0iKklRmfyYoIPsrmBUk80m+Pp6rHYsLKFgOQtq6MAxxftBDLv4C4BIQh
9DFZnyLthoFigWagO/w6NN/MG3poPZu1/G7jWCkL7O/yaAeLoGWOt9vTyPRrFLs2
nWUGXLsL6mfBOdQwDCVqtwtAAN2j/I82GLVRm0LNj791BhSR1hqqbbIasRJZwIiU
H6jMwXP01Mpi2A85FtIFbMk/oGa7VHZIA5oUTbqyc6j/1QsydcF0woFqWAk5WCkS
8iSf/02JFMW2F0gyMr7Lbfuq4LBQYWf4Bo1RJ6c39REJ+EglwwzLyW2x+wCi/rMF
ZjbRHzQ+ncvmjEeun3wMOpDsDHesa7ip/UNPvKI0AOZ9ka+XDyBEokAFAItuQpAU
i7nF9e3bJNgddyCjFQPhpSIP4pfSq6Z+S8a3BtQJOoMJBwr4xKCxQuHDlJTIjbLV
UbiSzzux/OopNEhS80YkxA8VBlc7d5P/YLc4YsnCtz9SC4uRfLb1JC6297sh0Lvo
f9oT4zfZrM0CGgws5dk5w3897Lo+V6BfaD7ITYP/VHzLbwKz0TM3L+x3hlSEjkXc
fO1/2tDr7IEqfGbCAldB9k02CxgG7EjxQAHADcfDDJHtz9DstG5XDXiY5GFWuBly
F1oNjiC5wlmenYsUx6ezJVC2EiV+6XBiQG1uviwik0CyFRkfAKQSyA1v9mSxOHCs
wyIdn4d6wcFqAvnFwMwauFK+eVHQNQmaMF4sXLEwldhYEw5gXspD+BcgTLN3Ui6F
i6oZdeLOZurw/8u7ZNpvlwDjLhYceJMivC1ufUBs0RtTqqP7iLDmgBEVbYWbpE5L
Qy16+vX+AQvyiMD/T0eUXje6T7FsVROBurjZxmUsRrJzYQmp7TVY9ezzeY6kMFMN
8HrZWA4yqGoroFYhcQqA0m/9wVn0kJ/I5CcG1nm+1f5aYHXHXcwytxR9+zGl/JZR
Q20iENLUD3ryuxsnvKX2EKXAbeknCfIhMdvWV4qDY/1LIhype4BrTZY902cyxlbG
jf8Ht9vn7HSpdEg818clu56IQy2f1PpBgjfVuCnm1TZ1bf0OG+2a2d9uaEPZ/xVR
DKxQNkoclhFYAg/33SFQt52zgWBrMY6V9nusu19OM1o8dy0fwuotAq+5hTXebucN
mQ42+xhs+qbzQwk9SEAlvu3jYg/FGiGL1YiCpe7nqwE364Vrp9tOMdi2v9HSKIgA
pFZT5aO0bLECWi2rT3co6shbFbdc8murdW7sistMdsUNw5KKKev/HefN6CiskRVY
DeEzSEsn6oOFD8VRfhM7bMvXGrL43ElZ4z+6cMcjtJS+QGpqskO/Ssa/yw3qHDxX
fBz8TSTox8DhlahgFoV0NQM3QRuVv8kTSmD//nNOkYOoFL/e/BafCG44DSj/QGzp
1733DGIvY6l0ymIg/ylqYvqtYVGQT2eevMJSvzvvZ2UOikrNCtzrv0EDD8zF9VoP
aywaY/dDXPXCVPXQTSgTF5Z7Kv7Z26BLpfJZ8chHel46SkramaJ0Tm+njDLk0B+/
LaBM1f39vFJi1MTde7sKATPrTLcevdsuRx9wPxSM15UNLVQTggZ/g8FaaVddlGyZ
DPbz1b+ZsljIj5vVNa4k5n0ed/50x5vzgcGqgabqMS8yF7FgTeQBj4ZJjPQfBOs2
4Eb5LzHhZ8OfD8E3xZuFrzJtQthBm+t4gBrvOV4MMUXkzWnGhsVYvOAumoToOaj/
jkd6RTfDRzVkpXPjgjqALPI6hFuwqD3v7mH5oeS9SXgIA9gJq9WmTf7L9I1LMDAU
eSPrPRzk4oH1OlguLDWYiYq2nyZPBIWCqWfhbycc2YGJ+scmQMqfK3mguKh8C2vz
qsjpzoJKZVFylJwtiWuhwlng6lLENaCuqpqAbbv+sEq6PChPEHVsKHzgMPlixr04
YLuy+rB2yd+R/luXwMtHHXq8IOpa/uMOSzaLih6ShHplZzjqsKlzP+lQsd50GBJp
XOjdPXgB6sFwIN+6iCI0SZb/YG41jLYlo6kdAxBZ6s4doAucwGctrEdPv/vDHx6R
nwpsSiV6Zz7jHhe4wxc6JAwAYvvoa/MmLcPrwPtRYajQ3XtM1R7Kh3CcC2S0mFfL
P5c02wPIAfZbQZyrTRgdo1lvGuY0CEVdgozobS119ymP3Bei82NxWAt0b2DNuuzR
eD1IAHZkFajMFnGtWQbU5JfKQImzPGyn4UtFrhf99BLVl6g5jCMK4VyhwZZIQqG4
v+Z6uFk6gCtDgsl/d9a3IEHG78OkuFTHd6J3wZi07yaWtrbJKoyiDXoPgZUbCZl4
I7L/N8etfa5nU31kGESeCz67YgVQEVc5Wbm41SpXX2PQ582mc+13OrH1bve30jjD
5v23ErJ7W+mXROXuTmlXoOkegfsZ4UT1hImpHCAvsIzWqR9YANKjPhf8LxRDq4Ur
r3JHKJOWYoZoY+HYFJmKG0cIN1jJjXGQhVZUEjB4vewxtztI58WGQ/KAfwy3nnzI
xr/AjR/b8cTuYc2J2h3dDx5GNzH5jftYesaIIBLEEQ+aI9r+FyaVmR+Ta7v6+bjh
HXKtaiCpyoFRcbHFkE7JCvFu43TdKP1U9vQCIbf7qKf/IuLd3YCzI42YWARGTPwt
Iyyo2PIT8YHg6gYkQ4UV9rTMYEtsqMhHQnMskdsTfYyXv7cLvZWHb8E50apxlRKR
rBxAAlWZZfnxSLZEmFEcnO9P1Ga9Hys4R2eiDIASd4MAJZvC7TMsCYxiulPJmJc3
n1NcEEj6Vf9EoYv0FEN+m3cPtSXYnxQjSetj+Zz403gyxZ+2zH18/IL5xSEQiwpH
n9/dnsN+RbydLhLL7WpJlmOac7Mnm+DgmFCSjKfglpEpIUe9lN3Nw/2If+vTQhr2
F2wIdM2Ss6wipt/Qq9jo6zSVebYV+kMmBjYyQxQcbxV+jGmDFEgGpaREpBi38+Nw
m9/YCRudTyWpbS8bXM9NZA8oShoyfZGhD8J9NLsgwM178kkmURbNV3TNedbJKHw1
aW/gkDRQc+9rwfcyHNzhHhTyOhUwp+vCLoQUVjprXpry1D51BVzUwK9qc/B8bSPl
oQKrKkujP/p2T6dx0h/MlUN1jpWwTuTdJKfx1kRF9vfqnJmdBzVbuh3P8rdANmsH
4sjts1fAQ5jKi8tOftcMoxcWxUfJCsu/6jSt2ETGyPs1r2941WZFxNT96I5HSaHK
6GMci0Vt1JcxpPOsmhDeqg9ehRG4rmTP3qLevFEaUkbE31rVUzWxhPHexU5GsAqr
Q6yEGU+IR4l7+UxjT6MLA6DNojHXbYTqOFfMLINXfbLUyEfG90JzuGxXm2OtGMdC
7K4Mm6K/nD4kzwcGSt1ikHgGZe90e1590r8TCcQyLOct8hGZ7s24PINtmWSmHOJA
op1OtjGnAhBYa8HFmZwNkkIIQ3tSaobmSvhAPkAt47UB6R7z9BqkBIvTE6ZWRqdN
l9ypoAv6A5LkCqqEjSdaqyk8hSG9shNdPf//gMd/FsAvcl2Eno/lglcgY8RpGV5s
FgKc+shHinIajmG+jsW3vekRYWa4JSmKHvIos8b8p6L8AQmgOkW7gxKPQsgzTI8N
K6/fTISGM8r+fz3+hxP3VLR8zPyAmeNyryc4UPSOjmFcu6v+8g966jZsdiyjBRNW
gr0055dgumeDfeQ2fDWIfzYJ4FFJD/iBsBKsLErVqwvYMaPywWTSxB1T32xjrtFr
P/kw4VLmeCe2xexC6tsJQMcblizvfHwoRcAYObA2Z4up/k+vO97qtLled2/CG1jr
As4lYq2fK9b1ZDwDm8xiSnN+XpZiHH/lbj5euH9wbLWUP10ewgz40+HD3cippDRs
8zY2ht4SxQM8X3JStQ34seWK/QczfDXblyWl448Pp1XJ1wYLWAsMWZBZIFQhRj66
jaNZHmAa6ZFLcYFAoW1sP8+UCXiBe0rxmoKhAPIawHHUkH+GKusKEL051k2MxnL8
l6/cevs1jnjDarqXxayrNw0M8szJeaAhjrtY6xkBp8YSCtLLwpkWQy2t5hVJFp5K
Qc509bL2MH8fuegXXUk3qa1E3IdSy3z1DlESjpN38mUsi13wLQ9Sv9L2bxx6hgd8
dhnzw/urJetSYj0fCZ8mqNO/ut8gceRiMsngYui0hXJoqCU1GSxlZX9u9KrkV9D6
vmZFt2Q4S5Pwp1GdHOSE8gbfbzM6OBUBUDwXXdaX3Bzo6Uezj5H9GcdKJgLh6RkP
2mczpiC+dxdWADQg7S21YFVIpHPFk3mT74C1IrgxzB1qiCXz4868J70fzXSFMjqd
5h0aSmA8B8ygPuN0rdnZa8qKokJwk7xj0zRRLVKmIdKBbcXxIAi5k9YPRAvNKA1F
2tpK1nOSUqboXOxSZLYn2S8UpGpsuR4Z7u1Z4cRv8i+DoH2sJA79JX0Mm+ddcJ//
hEKY2akjGU/a2PESTp8OJlVxJahrEumbEGNjPcIdIYKJN+x/OVtNOwO4XYGdrq0z
tsA+g0zUaRo/dZdBydBE4sdEieRMaaKMl1tjyIpS6l6aCJWrLZC2cP4mnMO+IrxW
heIMC4nPyg7Oq19b8Zg67F67i7rhJSiwvcPhS8Tmou+B/ukGbhitEI7tRGtCx9oe
sfZTsOLrjlWz9TYbn1NeLWUrjqsKEgQtPDgebhuueC6gmergVnWEeFCYoVmKLQFg
TPVZwQ0FtBb78vaTuoH/NBQqqAuIubtjvutFQ44Id2BYIZNxAbrIZnZ7GG24G+sZ
LtwbDplh+P1KZfX8oCFsr6qyxj8Teopl59F0kNj+lYAzfwmcglFx3ma+sU7bxTfk
4/XaxNYxs58RZyEWPcX9fDIJx7uM0L7MQs0GMehFhqGPAmdamxxrR/qe7+ibHhNi
ktN+9N7psauktqrg15IUC49OY7zzEB2r7g/ChHcsVo5+8dsXzrqollPoGogIRMNv
7fcVne6yc7MkxaXNT4ET6lgV6Kf1hbxxSudllhI59v2TBizFR2LQkHmXs2LXPtHX
ONVVrHaMrraEZqRNaZ8Kc2OeyVyU6XmqjxBi4pamO86fL4+F7WPe9EFZAhv11uv5
0BTgpGXagPORUJO93PKNnpyJG1Yx0wXEN/zKs3gbC0amO8sPPu+6wsZ411JBkzIA
jWOwG8CKgwXNdbMC3b6XLLNhPweUzmpYygNyJZ7sREIcsaVYlRoSJLtsfwDBW4i1
URgkUHGcNJ0n0j3GvYAdixbs/8H6zdnDtpJqnt9KaR4ljlQO41xe4wwBBZvO9b0C
rQOkmvotLPYue1lj0ar5eZDfIOmPZoGyd4yIzXbc/HsKx8C4zh4XYz34gOkTXOGt
/3929UUJ8Len0KCQHlNY2X6W1ic0qrRPdBpU2H+/wv7cg1ZiZYFBv8mpyXHZ/2mf
tl/IG7Jrt019FT13h0eqQMzaJtBP8yfzV9hOfq3k0hCvacWhHDdlqrTTn/qIIM46
auXvKwwiXR1upj+7MzW5Q+Taw1LJWBxHdTVAf9YX+3yjJATRgg0hJM0WppXDo5Xv
AhwoZbaPKyOPAEkDlOw6cfMLHRKM2jVvJXFKzPP5yNX+CrR1ik8IF9XQEp1Nv65A
Z/9QWehUAf2Ftwl63P9vQ47NrBJFfudXb3rEoOqPxXJaGDeebMeBWNZSEc8wqc9+
EBjmKFI+QcN3iilMtNS4LcCCpDjnEr/IXxU815TFHcsmS33mumQ26JPHoOWNtj7P
49nl1jRpe5SukXhIBk/s9iVX8tzu+AKrGssCsXvbSgBtdmaUYawC6dYYyXO3fFvd
QRl69GiIiEhJGjya17/sw9opcOEo/CiAadV3I/99dgxWRGPDAIp5/0wxfs5olTir
PLkKAPaYF+NAWucUUaG6CFmWSrXm32pIC/S5YYp/rDfVae/N6iZpsAaQpQljWKBt
TvnZBqNsqw2P9beQgeNE5SB9aoWrZfzH379pkpOV8/PiSS/936WQ/nS3+Jt0MkhW
KMmoxW4CV/fyfs7k13H0sgiQNsgOseb1K9SYne48oLpT1uuqBvLYxtfD671IH4Na
Xs7zJvYaT3IctIFRBooXtz+WsWOukt6BPo9o+OcSsipmMDe4L8E/Z559RAyLdefd
XaXuasdKXKpWwYIOYmjzDxC76p8kqkk/0Mae+yIacK7PznGAKsDpSmV0VXlJwToD
MgcB9B7V7ZuUCrTkOryZ9+tq7QjobjJVqSMXhK1pIuNexzgA6gp0jVxrhlRNH++i
Xh4vQQZX88OgpgijlQnc5EkJqkYe8rVN1OjkkzJxZdwU+v540w/T0g84Fn9MDaiZ
0/ACxXXyjZIHyPAA5oiwpmSVX8D1APXAak8gn4n5wXuXPdNS4WPIzlN2eYH+8RpX
121QYOg5CjxItw4q89mtSRFKNqMXboUO8RE9BmpUxaxpVBdNlpdGuae8hiviwFxC
lhGWPxZUkxOmgFLXzdnK14V6A38AcJCd1vpyRvSy1uoQi9EBEIMSGOdMuxmxq7yL
2Z/Yg1RLp0s5/FQRCTgGStfunKXsmSMiDyaLPhIZD7C0P4id+u2AHJWXkULV/5VB
Lm35HG7P9RWatihnJstEGAcLxgHhQVHbV59NYZJcivRpIISIVzuBvozb1T9aakF3
UnC/jVWy3ZCACYd4yR8LFqVZBxu3RQX0m3tGTz0s/RpZU/2uWpNEg+IThSbyxx/Y
ZRqWlnCR10HUppZtdGyRrwzPoS+E2/ldFDCglnhBZ2p1UGd5OZQuhZ1RIgFE7KJT
83cLvIH64woCTbVrxeN3tZY+TRKsBCxoItMw2N/t0wHP7WKQMZTzEPOY5jvyREGw
WcPGyksHhe5NWPz6znvXUgsfxNNL3ZVUk2jZUOTCi/PW+EiiOtmwOeGdbkv6FsFh
lS0UJmjgm7ypxr3Jv6jueuzyP41FfI89EjCegFYUUSEu8m7UcBTvJRNQVJMRRIlw
9aZ95Jc6MmLRnB8SBRN0yIw1HunBAz8EqhceGzGgM0ErzITRvO3RCSQuFNO1QdDb
FN/wJicqP3dd51LAlTR7VEZOXJ2dhBfzxo7RBgHkym77J8zbge9rbxSlYdt+C1BG
pbA/BW7HwEL6SRkjR1j0X83hHSZ2r2qLbSxmBlHtdVblhf0YjLTmA0JIwdlnctap
GyHFBZ9pBQqzhZQ+uW5mIEhvKF8TUr6tw5uua29jzbCrR+xIIzRxSZtxouTVgZzR
YviVsGqIx9gDp1mAqWmc0G2Rzg1Lcs/MENLX9vGJlea/oOiD+kTT+g+lLGnrMLW3
nysr1vd2sXFOP4RzKIM+/jQyDJcioFZqxtIBhQPJ7xBGWVSOuGMAvA0Hnzk5UWMw
C8+l56O8mGXKY7LT5RUSWaJNRODX50kfQllbxsVfr71lw53F4AM0fOyL86vAiaqd
xvG9CBz4c42CADMl1kuVOQJI0QSGMTT1FL5cwf1C9OpnaFqoZFU83pVZeEslNwiZ
78NYM/lgOz5JhqMPzj8jbYKlpBwTwZb8nTlepFGB9IZhp2n30qq/T7c/IRgALJoj
bkVo545eENC3u+vyM1IDWlg9ubW+xsMPyUHikvmTeKwDTT2uX2SWqEtSpTwqWdQB
BhN/mcuiyGNCGm0fWSFpn1GVO+0wgl6WZ7OyGSPGV7AxwsCiYVRgo612kVcfu0HT
BK5dKvfHLyHPdwq2ZR4s74ZYBdkCaSeYsxzsdGhCuWUA49RBdzXK1lpcPKujTkNh
ss5fi17wdalrtpYPRcS+ti7ZH4YYK3b6Z8YoW4Bou9q4xCacwmV0v844QU+3es0f
uUqvQFdZd5y11nw9HVJzEjop8LZVPhXwiNw9UgKQ/S8jrds3ppDJPC8CHC+MnPMW
hpuy9EgxzX2aG0E0P98GonaXk+zjYruGzf/kxntCYr9imZrCerdJCg4VmrOqfzdr
xybG4sAmyQJLnWwYeyfhP36aMlIEXxmFoZ/Qm5LIrUV9TWyr3q7e3Izas9gC8Kr6
9Aje4Ydo6QxsswdL8sAceHPZCL4oJQkECfQ9RDOd0AsE53Tiu/lyBFZd6qLMU7gD
GJvDjNBQwmOJmiYsUWY5asp0ChxsRBnAJnRr6cPrxZvqIGTypDRsfyDitAQCtDWw
N87S3haQCjz8PYDUYWz5ac2XKGti8s4CIqeYZufEVTquWX5AMbuZuNZpk4W5biC1
PgaQ+8YZyBBIvaQvnW8Ujqj/ZjSzNXV5MWYvI73SCv4E3RYN5gS14scnkIfNjxfH
2plt0j9x2gaLexMkHS4r4Ahnd9qR4M3uoaOCH9ZbXTJloUfN7HwgY7ixYdvCnd/5
NZ2iEg/FzWmdcIqQCSQRr66Nd0WX1kDif4C58+7TMMr73G/BgNS6UMIXCPOE2ieO
7U+t5CD69fB6wnpLPV/sOwObVtwrzSZ/JbOK2oV93/DSEZTFTJQXjrz8ranE/ow+
OQqqUbYWGo+DjQo/B3KieOMTuhnL47/Qur9tpRukr/2vACq9UHBUwYGNrEx7n+ie
yU76fEUshii27bS+19qoBgKqmX/G2scoRuSTq6eeGgljvtkN4DdT3nnbgWf/imnf
Z7ZRl3l3ABF56Pltsmy5crFMq1devfI1u7ZTP8a/7QO/WDwPRK4+nR0iKs1cykEZ
vJ7QfnpMdGms7ktE3U0mZVeSm65DVLd1dcle6tcelF8OMHwIR6lH4v88LbvpMWdw
ZsNnqS0cSIYrbbyzuP7hbRp/2UtxNxVdFeREFzxLW6P8WD87leeHv6u1UOpiSb/O
xeAO2CXFZyTzorbyh/D8Hyv/8FHuS9zYuksrpo4Hs9DwG36vFhPjkoU9WEyqkSWn
7xBsP1CIW8FzldfvRFG13Oqi19U1noTtvaKydkcF83XloFu7ahwKaXFMA6sRU37t
4moEWotBYESmEkiavCUC5MgOyQ0UJv3SkIS3kJYqAf9X1iyPuc9negafaQsLkJ3A
HpW2rMa9hHm0hO9DyXS0zbdnqOUrJVwiTIhhsPldqTyMwwNwYh3CPyan0zF4o1IW
zfKDqWNZaQTOojL0pbXc2IbobDKAxGq7iBRV0IwwcY80vJFid7FGRg7xZ/MnKEkj
T5UEMv//WJjYh3aPBtck2LKKWuwQc6RE9VJEnKMJGs1vt5nJFUZRsJTVx3ApH8CJ
l0TbfjcjbNCywr0wkMwnWy0D33OCbTdKNGU12XOCSKleaXQwhxP2l18I6Tj2FqpK
Y5XRtpiOMcdB7FpdcciuzE3O2Xa+H34iOSn7VTxzF+fnzWDFI4XcT2bTsFjSzEQF
KhbiTTRw8+EUpVVjdB/Xu7ZmWqKn/xDfluM/ONUXsZ6P+31L5DsGjP0P6oseAxo6
wl88KmCw5kqlzVUBPRdC667bcSBxeApoGrR4mViey0EPtLNv2slphR5QBeQzpoeI
VSQAEuTkQU3V+JVPaD9WYsXn8nzTO/KMpbZakfD6DT0DcUCj3qwYkkZoXtyj1b/o
H9HkCZEpUZJOPg+PAvGf53ye/Sridc+n0OSLBLY4n8u+jMW8EAgdhvCkBdFOu6xz
uEUEtuu6fhzzijoKA6tkw2aeLNBSdRtIiL5QX8jCVH9M2/4IcC1C5TA0aqOUekeT
Y39WFw0MsIISj/0unyGHCX8fiHOHbhopEgTEIn3Y2Til12+UUqrZgbCz4HdRK0Qq
Eja5NyaniwXE07AGeUqcMyW1iPL4hjiO7T0J/zJXz/FwGP/JtvD8kGMJjEXS5/Ge
N9Z/uCO+f7pfoSwX3DpN42OUd88bNu6srKA7Am7UO4PgnvB9YqphpTAB2MkOMHgN
YTrR23p02DQrIhgfu18Pd9XkHlYeYKFnxCB1R3JOjkvGUjGDTnDhlmZvnWhOCnNN
iAU7O1rghMLiH8cHqBb/sEyfmFLgTpvNOdPQvjw6C01X3W/nY7RzleazzVc3SDpk
8Y9Z9AtCMzNKJaKw8ywa5h5a82fVlLzBM2QufoHz4NO7200eif9gQNVkXM3eqPNT
yK4bjRdqBnJBFsrZPth2jKuGYxInNv7migG5GABBUsTX3B5nzy8S9yRovW4eZCaz
fT5MSSD43+u7Bdx1qOGzSnjvaP8UB6625Km1A7Fw5nZCeSoQ6TsO/7zKE+BDTIr/
XlC0TWuU9T1oj84iW5iy4ni1+Ymrb7FpJb3YTVj5wzZBMqqZsfDub0ibqEEz7qmo
ik5L3UEpvXapo4mQvY9ui1t5fvXrJalN4gkDxy/QVEozYkLFWGi+kFEXo4Cjrr4V
v7cnTWKOzkX24L/SKZAyxzfWZMe9D+/FCZL8hRB/fah1Bb3WgbNs6YBcPWbQjkLH
qpmO//XeFU9szl6FsOzN8Vt8k9Uy+u831gWIIVceh1bGE8ts8LMyM9dmocPvHnNd
XuSIhhpAcCg8LR0cNLfQeMovFwOZ9DCJjuxstKuaMVVYB8NkxkOcpnEHeZ70P8Qv
M2OKDDG33lxWqHajDP/iNMPYb2atrTSVUCj/VyRIrvFWIo9XF/W4PzCjYRi8cAyj
TSGkTJ9tYC4FDJ+3HnJLKUzU2KSOZVcP1+ursbUkduYBixFJi/6OUbyccVm2QPZc
jzTjF7qw/NMMMjW4y/6ATG4aIA9eLeQ4orCYw7WXe7/Uopsl1dw9Jir4//MFCPDj
fH76EpDFVqOeRHPZ+c6SF4n1bOdm3L62+RkLNvAFPNCR+/HM7kHFDpkk/TBpLDmT
q/2IbRVVnHxaDPYx7Mpgl3LOybgScxRImyMVSEg8hYmD9pxZBYKWrNboMZ1IXn7F
7D5+RVAeh4Zl6GGCGn0kSeQBKolWcglzlHII3LfditN67rFQX/B9cHpOAI5CkILU
vNdtm6wls3OADEAefjbNmeqr5o26psyZNCdFVCzgxRDRvVTXjWFh4DtRw/+VhO+/
a3wmqWlxt7L8jHweaj7gWCuZ9utdpYoZGKC1MQGr3MQKmSn7+1yYC4+TqCERLEZ5
ucF4dGnoiEcaBJ7Rm9u9/5OV2+kpX3LJ5eFHSNT1ZkQN9qd+RlyVlkacGyc9RfeX
9YO14D/EmQTnTzTx6yIu7woA4A3qBRYJzLtZYNadh06SLlu5k+G7n8jXwUiK/Yg9
lFZZxh2S4aNGKjieygt1yiN07RxwGOv1abvETX1/A6FElPT1iiInNgh+aOb8Ppb+
8BBJEi17Pyi0pS+nfR94c7vaaOdSkgGskCfwGyT/1jimLi9oNXDFqZ26JsFj+Ykx
92JNboQ03mQjGuPwH9Xhxc1rmglHZutMaFSubTPcAzkQ98q9Wqg3ew+zuhqmwiNP
3Y1I+ap0LFIx8n+gyndxBeAIkOf8A3ey2kcB9lVjZ1rnpVN4bAF13JOOmk7FhjX7
EiOY0p00zTwaWLscifbvwmdv7beE7J788Lci18cgh95e6AqsI60gIhPt74nkpGhf
pShAs3e22gNEAIzgvdQ4naL8tOHdqqRcfYTcZRDKs9ab4YsRsBvq1t66oNU8R/pT
8rFFef4xi0B8bd+Dx7C+dWO+6zDVEx/pWV1QdjIf5GG+MuCQmHFy9OOMLU9nkvKR
9th+ACTHzPgF+tWyFQTu0zp8+d+mjRd05jsQGXCKzHGk1kl5W28nLDtgoyH66QpP
ZWbp8/eQFoTMX5BSJA7I3z7YRf77plh2E71i9KZBVm7rTFnslv8GsZttfv8gnv10
XJZSImHIQySREyrVSh56avWNm5Q3G94jHcVztCuDqiMSe/8Emb3m+I+to3H1AANd
1eoJrHY1qQO0XXG6X1O96picZZ6RJSS89k01mY9pklcWbhwTQGR8vhVYfDhHM14L
LIdIFCi0B+pSKX1w2WyPBD+3GIaqaNV5OaWt9gDqw0NtA+JlE9cgFqiBCgFBUojL
Cbc1Ul9oaipDlv09TCz54zPKFrpsMgqMNYbd3CD+vLQ3QkjHFeElEtwPJd141FcK
xjiudG+qX8z6s8E7PisYFpNRWBIuskbTN3Uorc+VD6WPfntmFcnhyLGul8GdCqvl
Rd1RQsTzStR1D0J8n15Sf3XYgufS4NGa8saMKcY7G2Vk9cbdjrJ0HP6oWFy6855w
x8ui2DE3Dd35t++628nUNfoQbQInlKpSwKZt9MMNiU+aYaVWJapJk+imYIEHCZF0
w84165MVIrvuWbuVnKkvfFXb8KnNfZ/8R1A033/4NsfcOluz4tTty2gERiLvIvwu
IpFEeaZJoknig1nYahNx5g8D7zJxM5VeuVYBXdIK5mBS9ItQ6OhfKV/pCScXm88n
vpWeA9yo0Oxox75qjrTjx5WHG0tR2W5EXWMrhdjgLeUDplvbrhLjqZKfQfo8lrsC
UWeZlIN/J6fSIF2cRIyTlOKz99M+ubqMxiipYaS3tEbNGzaIEuleT0D23dcXK5nB
VzQ91DBtCghVjKqpgpl4vjpUvtnI7ADtmohLTRLoRrqU6wXyHenYRfngABenkwUZ
jTdw+cmUOBUPNHEOWTNN+WxklURkhCyQtdT87YTUfagCbpqXy3u8QigSEMYK5by+
1DjtixHjrsWHmy+SU7K5Go2eFbPt/uxfcVLdAMNMExVRz1VATuhrLf4MBd6voGRP
x60ZtL9k0Iv6tQVVuCTztvrhe1/PndqBH2AOkNEzZLMArMVYeSGnvAdjJmG3DQ54
aWgxART74BF19eFil64qMY3z+RlZmEj/BKr9itNHnIKHa22Mgx3UXcYvBEyFvZJB
I76bpXXN1yy3cqi/w/hXp8QFJrrlrDLg6PE54lNG3wDcMqRfS59Hv4GM4unt1XY+
AJ3mvEBbiPAWEOB+k7nFuWKUXB/uiCaM5GdUDzQmqAecoUkG5kktmOauVOvDQZXM
mCvABW3fjgei9KS/156+W3HIo5z1pdIcwL3oQdLzptUscaQhE2ZCW89H/N+WfvTH
oT8nzjPdWK52DB+fB1N/rqzY5bKbFoUa45R/6uvWQnP421IVvq8oF+PB5eF6w8tT
u8272msEGM1FmGAaV4yVnpGCyo9Do0itd8wY1lGuySj4xC5NCdrYZvLuOLAGU92c
4U8N1OaBhaO0U0yuWbj/gshgO2i5GZdfgnb0/a3/L6pUZyyuv/Cw5bmXwtcf8D76
8BN+lGGziV2CfhhOC3BR1/4epEQTQK33jydKFGOrUEAkqPyLEGII2zRariY4yoIO
vkjR9IM2I92hK2xDZj7pC1sPtnoKUkU5BAftZ1iNeEUV319bVWJT1u+32J4ZF4zL
cm3kAStdi1niz8GzXfMVyo2QHhX2EIbWCs8KBbck2CKUsD6BXyMJxoh6mIANnIGA
M6G7fza+x9rSzk/dycGoFZT5OStKIcsHbeb9dTagJPXX7x+nUP7RnWw89vzLZl14
63Yho/Pf5fDLvDJyiecFgFTgxGd/U7RMOSKbQ52bFf2evChESeIVld1DSHk8yWeV
h2RpBLtWPSLOJ9mZ1dWd/hUJs+CD5tDUOS6Q1SxXtNHXfV3mxt4be4GFgsM7uDjB
Aeau/rIZa21On46l/Cc/PwbRN8p0Dv/Dqu7RGowrZ6dLaoh1Nhpt67EVWvlefR9w
mc5VxGFH4cxuomHl3kv0hfm9uv0N9Az6HIe0ggnIUr8LW+lk3IiWib+tldfGGZ3B
tDpGuOUv9W9z62iEEglu1vpY3TiG2s+oEBRaXjNqOXepdwTtOZXmwuQ4c/ATa8oe
jZSnBMMlbn220CmGnfJwEjedzpxYsJaD9DQmxfaeUT/ZKpG2mCVrh1u5eunNtIkA
UR9ds2aRu/xzZm1LEYgtiqhY1lMWnUYr3WUblFHZomW52LSJyIsfNXGjm8WYvzcb
dTz07JTtNq7tOc944du7YoWzidD1knMS1O4SoxkL3eVmR0WFfD0G1lIf0NAHIugC
68hU6u6NtbhL/Y3f51SQg9T47HrRIUSwHBQaXxbqdZMABjNwCwh1CHNb/NMacMTa
vUnVQ4tf1amEky6sw0Kq0dfHsNM3p1C9lGEEGmwdF6c4F7GnVfDo6/8EoZVmzg6j
kXP+fiQSJ5opPIYme/CGLkdpouOZLamm+KcZ2/18hxLiY/Wim5b28NS1AT4yGRBS
PR1TSiX5PF8Xgl5mEmlkZ5gtftke4kQ5ojoht/zUqgdZrsqos0F6Ofy5sFXq/8yK
5WNqHLeejl3+o4uAz47ChtmFCXT0HXPmy/NOSLK0x9mlzXJdGQL13LKbFt3OMWzx
lBF+qRb14aTDY9pH/R2xt+nVL0QS+B2Pif/DF2dA7axsXRYf3jgj0ADKI9OeSQhx
RLghCFI2Gs9ZREnqRZvAKIicfRay6dlCuvBJmdNZzxefzRkMNqn+gDH9c/ENxb54
3sUipwCM+JBDPfnwkuviB3ADfGZ126xS5CmU7f7K4fAF1UtV2h2JdVcT5sVcPyeK
tpt/Aptx3oVDUs0oMZtEdpLdOlYixawgAYd2sAubDWQGIuohM61HeKY5XiZauln9
jnbEdDkMWeiihQIur4zHmdYvyOhTX/3NUB2qpX7/mcj3ha+M6er3Z8XIURyYG3QB
5owSm+ChQyM+8v79LP5oQICOzb1FoljJi95GfqGc4k5uufU7U9VtOTGUFkNykGHr
qvTy4a/2BDXQchsXfEx3s13GcXbTNmfZUbzDISHFRBhObVVYA2tNl7CXZcXybspT
MuS9KdcxYy6c+bXr8EYBVpeOOBIn6mcPyDnjNv499EgHvRaetvh2n/VwyPV9FpHx
36+IaHbazgDZB8yHT76ri3BcAfktgxRh2OJAw0KszlO2Sg31uuoJp6hP1vGPuSGU
ctvQt0vDMUXS/TCiIbdwpNLNNldPXyTbl+N5ZxTw3o+Tx9rHBMq5pBtWt+e/f5zM
TNKLobsewR850y8B0ACMxAjqjo9FKlI7Wsrz52rU7kmTEuCTOUFVMmsChcdpD3YG
ctk4KT1ixax3xiHDnwLE7xklKQjWbMmJMgrSi6U5fT1f4s7oGhc97n19aeCOO8CU
tpUaeNLDg7kdefx0N6yvdUg8vbliR0/0hzhxfDvTAmmwn9tPMx/ygT9jru1n3sNm
xCmmnNW92dtVk1qpMPOjmf/cSMAJxO2c1j2ozMsJf3UFBrNY92e9wK6XrSMKIoEF
2NWQH0boQWxYjMX2HGr+lfqCIFRZM/tNEwsQr7h6+/VRJdR2BdhOTuJLZo3g8BXf
onqwIqKrMn9FmMVTnvncNkGgRikC5fH8TQ7YLinjT8CiQS+pwpUqyvKU0FpkTIXN
e1TmV7Kx+de6rDtntdb0CaffUZylRH/6mzBL2SGbBAsIYSybZOM+rlR58mRBMJuk
4ISznkkzXeRT2xNLmkIOVWAcn/caZ9dcJMropFRPDdW8u+AFinb8v0CxjVwbYOBF
CqoyS0viNHggRmEqVnNdBm8t33yMoSaSwH8AqNSFlvprkd2gtewyja60DDu5djJt
4DPoSlq2W71BL2fw2GHNvnO+6OH7H4JX+qqTO3x/kqxsd+WsE3cewKaIvNJK5TXI
eBVo2tajW0p1Umhrfcq0iy/6u9VSUCWJYV59k7GRaiVj4ly6VZU6wCYn70PwDa0f
CW96YpsIbphH+2vYFEVjFy1wcVcAme4pdwgPfqWyszfnuxlyOY1SAhBfxfdfUGST
7P/iEqKht+LtUKsX4iIgbjoh7IbdkR1PZRkhNee09DiLP537zY08tSR9vDRqbriq
DdqJYWMIfntk+FdKaH5qCasubadcFa3dq5JBPO+SFzLQWjHNdoVRmB66dLROC/Aq
rZw8R2s8SYGrAsWdzuPAjjLUA8GwYOzW69d8mAUTVXo+KWRhhbv+QYYbQEDs0LI/
ra45I0UqnbX2WVaiJbehcOFiYFBGTc5Qk4pFc+qTDVHDZQhvDdI8fFh2cy3wJm68
aOmVEou0WYglEghRYOrU5+sfW5ax6wusCfT0O0QpjRsWWomZX20SBFXhPeYvrZWZ
6u41jiuw0sajevqsb7zQkQiqRLJV8GHGGkchXAaS3gzF71DIzH8HGc0lUo1pQ0qD
fEYwIwGESfRfik23JNwZL6jod6lUx2IqrvrhlVNmS0nFY7jxNRPqt3WbA552wqge
p35tsTgN6yBeP8YaiSW09o/HstttXHwiQhVciegXC2NJyRfmJdxQ6wNJI3F03lIL
ADyoRij97DY5bbROWTEjwuJshkLqjJEjA+VMmaRxL9Y/RkzvyqZ7Nx4iDa61JZSH
90gFQHiKsdzyKixR6d47MjT+u099h3AI4V8gqG6zIkJh/JWGlcVhaNsri6KC8GAN
Qq8Madk4NQHCcQ+Q8E/1X3ACxX6fIussapRivtMPpn/ncWdWZA56nKgY88v2qXgD
2+JbkbESCmxZ835evukGns6Gg7w1wUmRRt+u+LbxrDJEHYR1lrp1wPgrdYCBYq0+
c937eZbrbF7C14e1C/J6IKlxIgsLzrmgVwLn5JGZO+WkwSKsgxlQ37srZ10b97TX
lubuXM1TIsxZXgGGWYL0ExTSaYCTOS/8UA2lmGOOIfgJjERjuHQxX0XglgwdkeF7
49w6UBneUCzn36k5ehMG0r6LECpLaPgqqHhONDRDfz2lO8jN+4rR4TUMMgnD2jcg
SyPHUiMVM6aoWhuN+GUCQbuo7DmQeu2esjooJJ1zIkPaU1eVlvnF7EQBEYPyzICU
pPV92KGK5cdp9jRkGLrxlJjL0p5oV254E7k7CBj8L24LHZ7IliwQCYVKmT8QW/q0
8QOgwvTPH1K+iAJp8bx/tsj0+zBqrRSZdj9aIfO6W26N7F2ZGUwABPV4XU2/+QS9
DeQV/YRRGmeZ5YQNP1lgyGyBB2st6nEWf77M7bbZWMrmNhL6BhbDOE1TvvNMVOEg
CddPKQUO8doMaonN+jtvypihJrJfiyyzbfQbdHMeV5Gf8o163hoDdzWJdDqXDTBH
PhpaVbGAL+p9Lq/jn+kGbytvk6S1KJEyINiZFEfQ48JhipS+wglz0eSFs65zANwf
HfNEuEMoOlkuUa6Q9Kj6k2lKAQZLf5yw0JgsLL9FC0amf8EuosxfhUtuMuPpV+HP
WB90j5Vm7NBN/OPe3W1rk4Ti60rOEkDAzuAg7Bj4uqjKe76LzXgi0B/W8U0ctaWY
I6PGuIYEO2mMDHODsdRDGRkuwt99PhtSB6z2dxuvJN1C+mBFQbpefS6prajhMIo8
qiTILGCkwcdA8qNn1yPY9ZBYVaF08qOWXhjCJhQ0behf3WrzdWdJXApTx1PzYdZa
0IFwLFAzaIRBE2jdE6/SvrQMA3FfCaSmdyTje0vHj6Tsp5lBbQomsnWtpTyWEOy7
ko0MuyZJE2+hQ16RSFM/FzYaarbH/UGfJ/yj0GrKK9+s3vvN0hj+CXvm3Fq+05n1
ZktJmdwPUahb4qn7v7drjxqCSmI9WFlNru7EeFnv7+CS+EBe4QSIbfbwDBn2cuOa
7LykHIMDXY5InWYmR2eIdAF4Tuy1XsC0tCNJy6EigPAksHxIG6HE7xH7DUB36xvk
fyJWjVmVaEQdxttR6CSriglLmLNgtqaZu2k6M5UX9lJkz0ocO9jZ2FYE+fY8Vb0o
VuCsv1rsdvgSssqr86mgyUHLwirH6P+KxVhu7dWoorcluEOx1XcphVpTYeTZEq72
prhsPg6xEg7q6ddqmjNbHnLclFsYzCJo49xXVGqEcM1XT/efUGVSouc7DfJeX+8G
DikP5gr3q1KueXAXuRLYMMYu9YpzqCeeRyGPBIjaQlpMfZ1/v4jdBCMQKEp/VloQ
ufeiDNZ7Qn7TImvwrtL+qP+k7Tv1DlurrEd68LvzoGR6K+udc9hKmmJmiEAZBZW5
rpJhWK2f6xYC++cUM5o7Ycg3wRTur5OcW1vrpOfnI8KPj3mIMwlLVBWzcUTHhfcJ
91Y1sbIssb4Fh0v4yvChQQKpdJkbDffp8tKXJyNq4ddyPCCBabbV7kDNN7YUeO4t
pALdPjWdwQSVu2pQ2DgFFn6rzC4q9f3wxE+Byr8XjmjQUU+QLkHwv1MU2BF0vQty
uXPFLqpHX6Re2xp26QRrHY8CDC0YcJObl3GAdUi/29G8TtJQkYevxCDfXyeBH7sV
jKa0C6F0xe4l0mu/H2G3PyzJmeEIqzo3y2oivelxB14tqAIfehiCfEw+7wpxB+yH
yUwf6H9yhe32mMaqGzb0e287b5rdNb9C3kIsbYCEYHPuzAUt4ir1I+gV8MN33hEd
oYq8aW5kkCXYUtqB1Ivjf/DanMSSk0V+MjhpjXfVHTvg+jKcNAIgn21Tj7AxyNAn
ocrLPdg8+k7y7FruOpjkvz2CHeDwEj3uBkqzP5NLuaCMst0UODdE9X2Ui1YuGIK6
TgQdto3/tiDUlkRZPRILH9LjHaquQVCG0DcqoUGYPybeK1GYFN78RNJyj9OIEfEs
CL25QK564/Wmo6UEFr5lrvHUMXaYz9Mbx2oK+rSnxOAwsvI6KcpiCLclwh+bq9mZ
3RlTv6kgdPrcabvfOIn4PaK9+I4DQOYWlodiALF/2DuDJRe+slpu2xpNBPaKu/cT
4jGUkCRLHcVMImiqTeXsDijAQNXvw5ipCzUM9eH2V4GkjqyDRB2DZue6GBJNRfQt
4IUVRtwD3QfBnzT9r8uMiZSbQr5Yyy2i9btZlxVFsS5Yrtv96ieImbxmOA2B9EQk
2HPM8kDwRwxmAATSsJ3k8OP+D4S6fEk2q42hf3uUvDP9Xprsu42BZWDJgy2JKgXW
I3qMZi5mES0t2BoXXEVnwyTehwJR0w3TbpXodgN+hvYcLNpkeZPzyXjZLF7DFa+r
GB/qWajo9BpbAalLJ1LQGxBycSI7aQyZ02M/U8gZD+EJAMODB2rFV5JW6hnN+sbQ
oMVoAou1NBVaO7hkP//FOveIj+xyavmcjFq3UBzsdmcPEv1Jmn3rCNfnnaL6cyn4
xREvVIjmNbLQmtKz5MNMpTJyzOsj96SWbIM21MCtMVITgAWRgvHizIxeMRytCrvi
jPrnUiGx97Cl03fhauG8v/X/bQNd5a9VRW4VpVYgBSKPEQBTpGLJatfzLCMxZAkM
98RQweHWtUvYXaJlHZ2INC+21AaEH3aL6c6+Rf6HUMlFBOO1xE2MGdcFz4u0Q0/J
Vz//+OuaLo2hFmCyHMRzeRJdl3Ar+UiXyRE5X34mg9JgdIGP5hWg7wwD24AJOX4G
jt9EWnRyqpCyMtHpLmoX82IrH6ecA56I9IT3F2eSzgkgsGxEBx//9osaziB7Dg8U
XKeg0bBlLA4M77Bu6fojexo6QaA/1AfCMVVCJPbgBdMKFS8MtjV8uAUZ4m1zfQa/
W3IUAt92hUyzQCrcxuZDm42wxXzHN+XZ1rpGUiAf0Q/BT1QDjEmc99wOTvHToBAF
GRs4pe/yPNlOPWLAVhXXK9piAo+1KrTosb8zGP345olJBo+vOurp57PgCaOf76tk
2Uc/A+ubjDONq6bhpD0MQo+CoTRAdQMOATKVFOifnSRwOzmbRv5xTU2PSTdQnn//
x4UeLcThx18yrg1bzDsB8R4ZFdWcNDNKf516hBC22CsdOjHirxSDXwI61XEipio6
bYbIHsTxaclHNrfifpZHCTFW6ZafDpJbD1yG4QAHDM7E8eV108QTukMPKWII8xfv
qI64T9ABp05clrJvYtdLVbuuUcJxA0eMFg/k1RqAtcV90XBjaJf1dHyAiYBUQ3VO
WMldz0BKIJnEMSBbBaOc8fSTefFdjsvtYo9LKwF8RkESmT0aLsmYq5qopZ3hibHh
gx/qmsyj/onPDPyxKNmi5BIM4bsXY/+s5YvCm5xDKCA4gFVq4+6x20rEsQltmWld
eI14dYsWb5VaVZOiCTarm4DGLsys2cq4wlt47XNPDWnYB2Z0xojriTEtbCPEz4Ui
/FI6JU4+ydwYbcGE5C2RjtwdjxnHsX2KhiEpEx/+loVHVJZNFVlz2cyfEGSOPuCV
gGpGUu2kaIOatT7Savnm5xBSOrgAzEEpqFB4YsnOJQPXfmBtcQxNhMp0dOacj7S7
S6wcBkbGrM0e+jGlIzX9Q6WD7RPTwcq8AxqlJnH7l7aZS6jAAcHFeLgyOPy28v0h
N1It1aBFDJRnZB6OfKKz7n3obnU25rLU8+L7NQcu2fLtoQTrMNTZsvcOEqFkyeeh
GuFHJD3AHmribLygeEoH7EMAL+QpRCTGpFlz8qAoQD8Txt710jmF5SOoSqiY0PGI
tp9yEteTyCovAug12UtTqwxd/J/2O2pJ9KoHcP2Krr05U6iiC6OELRqCoZom45l/
+dRbX8GVijrqSkDQwOztZ9wPSbgYRJ1Vtre95mruC84IHdAyoTrboOJQJWCYpaKE
quPxyA9jSZZEQs8v3rzg6vF+7QEvx0rAaigO+RMj5HFcY257FsWAdbqojhkOLMEe
/JD4ypk9fneJQK0/N1gvW4mBjcG58xsdvpGVIbLfX3OohPYf996H2i7yYIUG1RD3
oE3/6dbq2Qg80z3umHI2D3ReG75QZZqolX0c36X3zDC5NugNuacf4h/45ZESRsbK
UETWJB34nnHXRSz3QaxOoSznizw5x/wDk/L+APdv0LdjGK+mcF/q/v2h+EBLo0jY
WHQ7UqfpTTMOkxWDR9FflDarLrcmP0M+uC/nkTi03blRDxDcJU9qeFOZencTfrs5
Olz0VmV+UIJJPWg5/+ZWyzBy2VuvRsK63GbQ59NQpZfalonBeK/3XdjNZscP2iWJ
u6V15S3xVdty4Mx4QzyV/ksetbUr4thaBYrA3bVBigaTTvpdVlF39+H4IvAaljn5
zWYpuyyHF9i940c/VbRd1AqRDWAlv6KI8hflTM0WGyPROmsYXRYExAEf099229Tf
vb78kV99cxrVrhIIVXoSSFPROxlnaM5Ibvo+NZ7weaX/RNp01iSAboD2VtuM33Du
CDJmoqKQJ3pjICfgIziil/nWgwt9NUWb07/P61Ms1ax2VpXzC5XP/bRCpDCHU+bU
WsSdFJPboQU5ahY4qfqTO0KyjFXy+oxkSMfXiwRv7yXfzI7horfyvG/JPZXowM8d
XwW3lSBGuh8D2GZkePRUtN46GioO0lcibXq2h//P5oSGDQSstXZ9LuQ6kXYL5jD8
b+bWAdn1cpo87kdGc/nVB5tUMmrU+LibqpNY3Hn2rmW/W9BuracfGrXevXHvLQU3
GC7EcgzL2ocYcHcuY6P1RHyqam0ZrGHtgXJTG8R8TuTStedUrnziFpCgFT72e7Bb
vbA3WkFBWrrvTzioOVT2bn5BntqgwVlFAMcYKA2MSZPiirgCfP6v2pJpadaB+If1
XyQRVDIITwvcyqKTCgvGKHC2a7qjt7Z4y9087RZ31VC9XgrVXetS3hDWITHIBelH
IeWqG3GnBn/aWoqiZLSjDBnMhIFX2S5iUCSik37dP88c00y294yNz+7aKvjaxfNT
xXfzihjWny68smlMoB6Vy+9iMrZ2aav09QAv7o4FqKCD31yE5pH3ZygyWoJDg2y+
9AIfpSilNLprtVn+O47NxjqsuaF4PX8us303BmIkGboxji8o7Z2QECdhP7M4hb9Y
yvL9uHBqg9TMBIjTgdnnJBjUIzl8qFODSZJDktenWpJGMWWpYTG7OswrJCSsZIzz
pkQhhHS6/atnlTNzFE/9bZVkvPqaHdu50fGAiPHG+FdvF/ZaWlYPZnwZwQR9mDwZ
eJxaSC2OEtOvPN4MbVryC8oCnZcKmrFt1KX5/WHR27OfFcALWFtcEiKFj3ZYwNtT
Mhj49CUsCwfXvLaAYKqh/wSPJQ13emN+ijykG6RMkR9OmXE7YDVQiOqPQ93tJKmc
/NujFyMfhxA20NM8tenhamkD9ubMhSX9iugW+9/M2OQJR8eN76sQRVB1ioE9R1RH
bfHAxNPX9rXMr11d55B2WTatpKewNPvZn0zDHlWhbcQ3DAB0w4r68DblE8ucjnhV
v5W8QG3xF9t4A1kBXHWlaPJ8fRoTh9FPEnRrf0QgTCAdpFqXSg1ywISkiwRvtpCf
cxysRmV9ST91h5wzNRcb2ItguDtvhy9tGfBlFd12PTitqIGd4e/huXzB/4LV70Jo
oYHAI+bzko/fXdemioyYTHAMIO9HkobwSER/yQwzfpDgxJUpO6PpA+6BzoLBkI4t
6GN83V5vUtOOTuqOIkq8DI2F4kDShgnw/LIszjB0BdOjbTJg9vf0RGgQ6Vd23Fu5
Yn7p9ES8n7gmu1IOzBzN+knNhbIABnCVq6J4en2sdu6xUbtqQxyacgdqMOxVaxHR
vlSiQd5L32a4BY8qop4Yilr8YBRr6sg3QmSFhVOJLVF6TiJdPoxmaPRcLpynNcdA
KQTxzxcj6x21nRHTXSeu8C+RKC9MnT6nfFetneDSh651xdyadZ49rpQiga0spKOC
/e3uAYh5Xbcg2QVUYWwrQ4yjyQ/yUEQBuLkk/svnlSyJc+puZyzTj1eKAdoYh6XK
2+/vqwDqbRVu/A0AY255ABbZ2HxfkwM8yJfJm5JAc3AfHRuu5mfcteNN+s1EngV4
/Ec6EyFYYD9JwysgdEdHVfaG4xf956jlzoJ+R93x7csx2/jY/mTwctRd7RevySYZ
SQqvDi7zLjew3yxAex0PwX6lPdnoCDLjU2BcoXZ2N/Cq/HSYuCarVJ3My7XtGrzl
m2q6LGmChmtp4Cb5FMqlf2lU6QqV407tBJlkQQmrPccPLbWE7IkqVxRqI5Uek7el
HqIQrJqRrM2WXJkpRByVN3X3mWtTnnO/6pTch3pKSSnbB7OmRAc/MaV8+S7DR8V5
ePC74EL0oSZ064VB9WcKbWRJkOqLtYX0+DfzP4OlkbymDobfAff6w0MfbEvfHxDg
nelhuSyLMe//obh1jm7YyP6xwqoFuM7jc3qNpWJHHgDoY4GG1YA5e9e3b+pFm25Z
99xHwv8k/1kvGDWzphMTcQX3Gpsx8r91+UAojK1qVDVnw71mJmWDkuVLBjVO16ky
Nj7mXkhXeh6RHU2iBnOYKj9cENEjp42xAV+NYz5ucHGmLbqa/6AXxZi3YiHkVPpB
jLZDfo7WE5ug84LgCB9njPsRzgYHEw7pMZHR8ZPSu7Q9YzmXfM0k+ZvLXms7xNaL
b9a2+gv2v0VWwUyEU7FZPSCBWe2WDu0IJ+15MbrDvPiyeOYm1fJiLCJsvIZw9Bmu
nD696zZIHAsLjCt4qisAcDy8sKnmT3cFmWZ9y+xsLm7HNuKW6PSJyN5On4teAOSp
zw0l/+q/IVH7TLERgCSUdUt4hDCc8zMPYg44FtaGD4PYG7SXfnS10Gn7HYP1VSij
g4JvNMRWpUhcPExA7NYkZX4z0gTuSwh2R/S1FGAQEXFQAiHqG4QxWiXmbUVOII8g
Ec1GzKIhNhwQfQcIy2abm7xKw3nd//SPqdL1j7UvtVtCH3qYD25lovcxoO9CiH3B
qdDNgsE3TI261BFljdekoKYJ3znqwBboQ7KIpZqFjXix6VzZ2/5TR4Bml+C0eM5c
2Ss//FS39wyrwCw3D8+GKnAuqkF/ElOpPzaXIV456v9DRFLceRQIM+hiA0jyAC/I
VF5P1KKyADLe1Y9Dlazu8kOf5hOfkeaSU0/zJfJH8RISuAW0j77ovBYMuClutj/P
2uVOTzwV5dRBI9tju1q/clliszhwOS2Yzo1tUxTNzHFtAdKN5WnbJH1AorjWt5n0
jEhj2e/YvFTPK1OxFQWTP0e6olaO5QAXzPKjd1EhFc+y0marZBQS6S+zVkgFZv87
SDUGwb8yua5jJRqlw2fhZBBUPj/fq1oNthxjve8tAbV80AYVlCyk5Uz7iASMcla8
f6lLuL4Qn7+lfi3aYK+7jC4ciSbnFpNP67JQ2CMkfMK7ujJiJE1wbSONPG5N4CAi
O0t6Naoae1BLY7n9wquWEZ+VM6Ra/LTLmySokZ2K43kS9X/1mSO1n6jZVR5oBk6J
HOq4fSq0RyY57GxPRWmp65dZlf678vaB5IM7JuPeW5Dah7QbShk6NgoKiTxP7eT5
UeYfjBdt1hpf5/aM5yBopNzoJ10JoUCnv2fWOQoS+/kMm1/cl03V8VXgbpe0JQPm
upGiemXJMq/W90XwPXrj/Ofy8LMcleiNKLJ0NkgzwqfvNCIeQYnh3FEcd+g2poaj
sD5+IozOLP9UQ0aNA9FZMi3tDtIfJh4BSxtvQ8/TAUj9Ssj9H8NLBiV0owRkfmyr
b/o6Vz/tkc8EMKNHv5o3ny5cnKBPi1iDdLbk9IBendCZ3btCMb/2Kl256K5Z1I7P
FucwFJGBXXGNUDf+pszTzDGnr9RqdExtm5fVnWREobKuu49ORcPi5RaH0toMzSYP
f6uP6mtEJlqjIGYfNeVj7+qxrK9mzEdpfqtAO9X93VbL797nMj5GB19CJRGuoy+c
DAbxdSKQOXdt1+jPNGNVahYcEki2BzuEudxF339PlgGospOWCLygxX0n+3OPKhpW
msRni+4I9yLqzfhyJJjFziL5zapVwFQR6sYXY/jprzehULISdDbUQF/33w4kTd71
EZc0iCPcHh19v5fVabfDyvFk0K5YDYMtWsX3RHLl3j/FoxZh9tqSFa32suUvmEqR
gCv07w+0cg+oYyzH9s1+RYluRFM6em+sKhe9h8ArLrNGVFcyAvZat+okwxRxMjMO
ickapN1Fy0cmHTTkNS5HOoTxg7uWQNAhyAMTJKCLAwqN/CZ1fCy8BckcAadVAfPa
ogD0nsu8Li9vdyB4rBNMmWcfdRU2Ixu851UbkxNJr22ntyCjX+vjXCypJ8xT3dTP
NBbYq7Bqp7q2MkcD4gzEn9Agv7CSxQT+iSQGfu8Z3mSUu5w6/tRWRfB7eA5Vf3z4
FY9aX0bQlXKAu9fufG+iRuCn5sKONB5qVff2N7i84CH08fjAiLiQIeZT3h00IATy
zl/8BDTX9ncon3sgUxnaQUdeyWoR72c433G21nTEeZjXJNDFL7i5jklGeklg6Xbv
8sc0GzjPRsskCmT8GgbDTrV3G4s6cjUUQYtcv2+T/jBlkDw4u/CiJeQFnhrbu+x3
VeMrtsk17lP+Rc2C5r5BwroFIZMFqlW1SntaDgyNsWQfyVAxMnY4ssVE53ZdvCyr
1zpYiK8mTwYKPd+iql65mSORTWg1MH3iJXAw8MmNTltjV8UIRIzVdJP4p4eteZJP
Lu9n+/CpY5EP3CV7LyXcvAMWSjDV+eCMVooF4/Lc1KjR3ADWXiAj2vK2kgF769Fn
Di5ZSBbIeLQm2fQI1y3kH7IealMuA8if34CEqydogg3Eh3oDaguIt45Vak7ZKR0X
nuJx8YYYprQUx+U2B1fOn26ogb2z7A4sr+WbCqFOoXLNB4kbwyKtCmxiSouCDcVW
5jixZ16STs5nUKmuJhnN6Dy5n+IVTkIfX6DSpmuhgouFZM4ne9UD4hvaZy1762Fw
zK4AXalENoFZkEtBaE9C2uQxB+pNqj7sIuit0o0JV7vUy5sH3U6MriAI9zYi59vx
O60Plt9bm4b4jrUxykaiieQ0DAu1cxPvS1lU/6qz/YCq2X4x1oBLqeR1lpIPK0hp
OtaJ0GWSeTQJA771It4JuULFPEmgbHF5b/8KWqHiapCwrE+4mfZE3TucxS/aQI9V
lIeISseg+4gX7GAPVBIprZENDFUXsp6+3k7v8f9MZ12grr4AYkuVjeIdCKoCoDfp
wuSrG+oEcmsw66ScPCH17HruTmOccz0OGo49wq6YHChoT0/PUi6D8TNNKJ39Q95p
yuULc7/8HTMhOc+6uZZt2KZ5myGcVjd2qvAkkV1ozOmFnymqxLPQ0cAzHaZqgXDJ
2X3oFP2fAYmQVog7ig1Wx/kgssHQjB27gf4Xrz7cQMMdUBc0HAcSK5e1/HlzCJCj
FyXkZFmZTUMu6j81zu0bVQF1+UKwnUg/eodc4UZgU78dyo5LnBRFFLbkANfcxxDV
Xyvoi+piYW3VQfOs7w/KV+urQAJ56MYwUi+YXyeRXvpE0qVhUUWPDfWDiPkGqkin
Zy5+/raSCwf0HH4sAzKfWGxmrOdbllEJk35PkEqg3Jzi41f2r+K7EQ4sfYPt27/f
ItWHjhLcQME9kSkkCfku7ql016uyl1rpyBulUZkBZfni0K3rZ8mcAgkDW+E8QKc1
cb7NhHhUPoMccBUOxcv8r8txTjgpY4jSwFVmCjJ9Y389OA3wUt2po/JRwIjBQujg
cCSAdwGR0jCteejmWF+5mKOAo8I70EBad2a4p2bmDQDScnB/nHD/minAxfDNST1T
dTiTJPMMdn8O8SkTZpvhSuhwwiVmoyqTnhrVxszE0V+xfXvjMSEU+nOTM6vzIa6J
pSRWF49VTCDDP0FPmKNMTH44y5ikuKlvjBvcHgdt0z7wEEHA4jKi1kQuG+Uk5Dmv
RcqYQbVGLXowpBKGNgBG0vlfswfeMhBoPkNIrWxwu9Hb+r+ewjeGBG9/fSbpjrcn
OMUcUranqa/J4ZrVxqgxvRpC51131ZU3pPrpMsuP3ZePHkJjz87P2GFIqPVjiR7D
EJZHSgn2fcU0OAE/LKjWzpP0n/DevhTvgCkJY8aoco+o5cU4ib+kcKTCUwkgEPa6
79/AsZnc+OpadXcyauQ+CsEkHD6fWw1VCFUNjssjSvASvWz8hh+PmitL4LK5LOyX
9UpjCjfvOoOC9qBrGldciY0fxmEj3EfeuYvaJCInVc8UMOQEkuy+M5+cCGoh30RM
pTTfWxM3bF6QIhoAvjkNGiA64uIwMlVhgVzxX0fjHmwnLnsLFT1Bv9YGO1DBGoqb
a9jyqMw5yaYmcYSeRXO5A9DmMlL8KvkSmqYaIAmgmqWVsggkusjnIlz9ad8rgmrz
fCQwqKYa1asmLs8ziGArf3+dgD1HBM6MSE//cmziXxX28YuW2Lmu0Nit/yKkDqtN
Xs/wr3rhNnAyD2M05WWMwCj64/tUD3zlJyx4NWvoA8D3rk6nJ3LLWU9lVy0M73e0
+iwMlSUNBD15gC8JpL+PdyCgJMIRDZkn6k29L9JJ+w4YBkw8TDjhUyo44GLlOk06
uDijtTovFsj0Hh8nxmiUgT4mFZAx2C5FIx7UmwJJ1sXgPBZ4hjHocm/Iav3DQKOV
MT/PaLg0MNR1ooNA7oXJvw0T3OZWxBg6FktcvHF6+Gax71orDMojRkeBTnUzXtJ6
WEi8FgAxDu04QWPkQsqZwN3s5yXa3VjaL7naFoNnENUN3Hc+t5g5ylm+Xj46OTem
TJEopWDV2ehQNiqsJYFUKrdd4qRrM1NIe3aPhaxBcKwrJpTGLlU8LwtPhoTLkhpx
GaUYtAmJ3G4HpOcf0aK3k6WJRqAgSuo/LxcxSwSKe9MtwpltXXE1nQDGQkg0XX9S
eOF29S5dmQpGLJfKVwDIQ6k0IdWtF+P6Nc22FvaLjx8emROTX3F1EFkPmWSh2pNw
gqkvqYLeXVVDr8+nOkn0vmGIUv60nZoEhiv0QNS8fDA8zd6ol6l7CKHQmc8QJlRd
WEjcCxtZTE19UY7gb4cXL6WZyUbAUanoMDMnuWmG9lOMPJi1BIC5Pybft6uM+vCW
6cPOu7YMletrHtkCbslK0O9hUaNUzQqUDq3jfO1oMhwwOes7oU6DIjOweqwKbYsR
GVTLLq1JhpOM3wDq5vF2F9GO7nGC6FcLZAoxuZ1NIg4AtdprvHyfhomuEYQUaauZ
RoNS4c/c5tZqNOK1ZU9Uc+H3GzvFasyWzcY7ow4BXSyWrMMfAbxzY5n3ylcIXrqQ
aouhKD2Ig7WsP5cJXjuhUUH67EVaGi5LR8Aplm/qZ4VHymCezI/gJUk+FgVVyjTn
89N9zYSwKxAMlr8Ws9SjLtUmKrYr3sbb8cWgw+cHtjyx8FDGafq81CYfQG0LQiR8
+gnaQtpCh76C28zwcQRCZ2PC+08LQ5kQVrrVw91OhHsHXvtx0gMhcBzlzejB9e70
mGNW/G/1XwL0r4Loqrjp+8UYSlfRzj0Z3y/RRA0WeWq0QBbNeDwzCFh9IbcfvFi4
RN+zcGt99bRGiGaJHZt9neTOaNEPjmhwQ3LO8OzjB/f5bb5fAYY2x/kasluA2Ikd
N19Zr4VgWjnwxejug3NeyU1vO++AUtBZhQ9H8tdJKFk67gpUcGz//BvjYAQJrI4F
MY8vsdBEtotr99BlZdecS0wiazzODmDJhT3AXwV7+hjJA5FTuY9UTyrwb2pjZC19
kUp8SmeoR/dYL5FLwgBGj11+qphUcPKD6biiYxl/80SyK14afhnujM+589/Ja+5E
0M1rQu1z6H3CmWabZUkiF3fAjjo6bFwF5QiZjRhOKArx2lzzLM6Y0hy5Tr2zCC72
dPyB6qYrai4n1oPHxTX6z/4+rWfQzT4NsCAj47EFWvSC0JqbZz3+LTSqJozKvkQw
h26rE4NoHgTYTUS9xESfGBDDTFeDrR0TmMNe/WGo/9BeUyGJrrPwNQGAwm5rto8n
8u5oSE5VfHTiiOIu9tkPQ14IdV5JLOAdMAsJihGUnClPdz9p5hkPnoHTQpuvpjP+
MR4viQv6ME+sqzWR8bjjhiA5n43mwf5QzRvmuff8K8zTRUmZxHYCoDQRShQDZwaM
eAg6igDQHi5ZxRLTNkvMZxlyKfriT37CPyE7ELxy3k8RshH9/BGEBJopNk1B8VQb
uAVvS4Oceha1f+FmGa1ZFBnc2/pe5AdlW+ITvA1ZY0PMo5dvRYJZi4VoT0M42TS3
Tffr5RbLHKBf0MaxeGgAO9vrMHX8OWBjbuqsr41txblGR3BvH5QjxXecMg58fhYi
LxSTLwcOJc0t0ZkuQ7xx5WSofVhcP5YRH0KmJUopYTEEleE98EgrclOZssmxXLVC
95ZISZPku9NZTaaliYb68utrRFGXHmwwJ/jfPBM/lrGjZBxnTRhdG2lKHlvprYO8
uiG692LUk3p/Zebx8O2wCBvHrUaYPQTGry8YgllNXwVpnnqvMPLxvlXtW3jBzCCD
X/kdg+bfQ+UENGPsVzasG4SjgQtSJqpimEyoS/OzHKbJIlJ7cQWleekUo7EiOZRP
UkOsThjUHPqWA5LJFGP+HA093CbYyETRzSnvLpFAbLsP/Z6uRPeF+3IyAuqhglEV
Vu1gO7i/aqKWMG+ul7fo3RAWy6yvJ428HOzFEmoZZbLzo0lSTTgNVU0+yItypYf0
XUZmc/jxccnh0DaVslkfX8PHnIKyZ0W39w9kuajFghQVgV3afqmv3VU4BmwPnpqY
3FqF98WU8hkCPMiV6wLa5zlUuvs7lAq1RIu7LJNdkHyAHGlpzw59rE1SX+tUPcFW
1e6tvJn9oPl6nCMvcOxxJRfFo2pTosToukmQLCTbn4wKiTR/ODeTshUvOBxgX9sE
81mOmoc7D11T7diCzD3zvUgmAFnbfUUALBhygTSGUX7uT0q7L9GTgyj0TCUwNBN+
CT4jl8TmG1SCRSy0WdJ+g7sz5n2rl53VAvoKXpbMs3FF+N0L5l4QeoN45c7b0ZJk
m0wJ+T3ti92IddatP1OxgcsNjBj/XNRXUekIRkhNl7qbX69MOOxVANLDWsO3V3j+
zRlAm5qb4ZHde6dVbSU9pm7aM9Wof6l4O7BuFp1Fu9FDU7GyO8py2Ft/oXf69LWX
eeMxbgLVZ86McNeiJ8kLqLkjqv5fO01inMzCf85lF2Fm5eK2I7f/izuW+n0MzTmG
uW7lRaOLXiB9Pddw3El9pWDYLlx0tf8Vz7N0cfAweDhndgeC1zY8pNZa6MP+3gm4
n/E8uE4rlKfTCgRvvka4JwKHwp7EX8IDAb15inV8TkzOkAKM7AT0XXeKodVZmfGd
r20VraOqQiyCLrb+bnnsVZbWL0pHXlQMu9ejAxebG3rPwdWygNUjK/WEzOzL/zzl
j2eUPwOpjG0MjNRem2tfFkFJN8514R7v/WtSFGk2DmFQHlpj04SwJu8Pr8O9YkLe
a/MgJ/ZhCCcIWXkHcFIw4AQk/vJEkz7quCdNyr9bu7zTsvqYwOWBvEI1bk/tG0RN
fGKANVIjZxlR62rFwGvjDHLUVSqX+Hz4jQz/Jv9AocBmmlzBvDIiSTksDOANAWp+
5qutNpBiLOlC183uaLkohgT7hGmcYozFZpgOphk+4VNGUK1cKw3PMWc6Ml7CAOLq
+yGtIzV0kipmgQO6ynpxGdKI35RP899YSoKQa81Y19Hr5p1bauXpu1U7aYbsFdJy
ek52AAtfzvk069r24BNnE4OqJKOjAKoxm/lEQ9iQs9Ax3f3ll/Ov8TtqMzmkO21e
Zkb5e4H1uPtL7sTs7OLp/6cgDkMaswBj9JkogH8qNnKduL+i2O9pkukBK1tYK8pO
eMTbksuHS85rnPffhncsHp7FEfEZomMEnpr7HVDknqao/FMshe+sTvurH/HVPhJp
2UQl3SCRgznpFoxH7a+L6AGzaPfB1LuR6r/rJF4j0mYsf5mpzpVeeBwWIJXy/TfQ
AlcGsWW2Z3Ju1tY6VS4cDADTgRfr5NKrtaABv8HNwjY7CGI2zDzCfyXN91DpeITu
TMJOfd/bzlczKyYQx69GeO9os1ng6THg8H4/p8bWKA5sf2BTUNkjJCLb+Zhh08y2
0/s47pL3rMAYhGB5BTfBrBHg5McPswTESO6ftwamWIvuD7M5mPN9MF9qFdcDwL31
5EPVs1fQGMzxScBwQyuQAoIaIQNo/9oW60359xDJvFms5V5muP1bXEcFLHgneopW
4cOIa77vrhaH/DQr2UHj8iQtdORCyBu4oYegrjBtjpDMrB9sDz5s6YP/FdpDQgy0
8q8acK0sVhekTVT8Bd/96K8ryub4f2D1EnF4lQB3UpTY0QFGIIpY5KOpAG99gM5N
B1HPF/SHsBWGHHNzqgXKBX1sORMeriajI/y94ubfA6jkJSIrLUv+sLCqPA3MpVXi
SOkvEt0U3VgV33/tcGM3eSgexqangsudlJmPUGT9q/75aXOa88hiSvfsMJkLJGdQ
5PjYol/+2q5CuZSf52R/mrPsvxJJ08QeT3m4MEqKKbEHjKuVSrwOp6AvAeKzCQoN
pQJdI+ga+CGDarcgtI9hSXpjeX+gwXha9u/JIioycp/1gSK3pItTkNDQJ45/svPR
O7Q383s/k4RUKKQg41y6vbvWk6LkwRlcDAWIrvyHAJlx7YhW6WrFdIWXVKshDT/+
i6Yacge6q6DQ196/ZAQJOXa408n6/6Zz+lEAP7GOtoKZODat1TG4D+EaNFau5F9t
WxK4ZcfYKp2QtQDcwzUBqR7u+umNTiDpUiqR60pP0sce8svR0DfgPMPY6hxtRsO1
7o3Bi1Q2S/bEgpHjMB8O/7jq874uRejU3GnDwsDxBXi7nX3gJtMGEulnOW4TO2u5
2iQwGJv2IECyfwDyGSb50ymN+tbCvgCC+dBXbeQIiqA/4BAwBU2x9EbKE60xs8hb
47WJTyuXSiskvAYI1CrM6NZPAOQXHbhFWiw5iu0jQys8ZXIwocRg1CblqpbBxTfw
NMrlM7xuKqnlgjexi3lr8Q4OHkxvDn+Oe7mbTFLQyMmL6hg34bUi+sFZtICniwWQ
iG/dd3EKFHpbPc379qUcdOlEMl5u03Z7jFIw5ECm7qTdBxdzkB8YbrE0zzn5LN8r
mmlCRsKL/USMoYszHa8ArwufTJVl0QJMIK4+H+38DoKBDjxhEIgDhPweqK1FrhY8
Afp42hZxFIKLo4Azfc0UPvqWvsr96EIm+/j3/uKtyOw5hnIU2H/wFUnJ+6/IMSOG
XA98bfiRuMeLHTorfF4rLgyVqdW3l96kaZsg8ZrM0qUVKiFwOJIeRY70LwiMx8qV
WaJc11E4lCNHd3zh/oIgJ3G7Xl6nd64p1e9b1nGrwHK7W19gTk8DwXHI6HnoHETV
JuRlabba58BXRMIHqLhJ7iwI9aPFzuOJsC7Xt0Nl7atwnjAaU3lT/Nn0VjAJePAt
O8zm4tns3OLoggsZXST0ICKg7Uyew0cz0+b14JxUDzNDw22v7laP+NzhMIrrpSkQ
GEAb2cS8QM9lQK+vAdph1Th0bQ04RzF0gmvUfZ5GC27/1i+vAMrnGATlPd+MOrur
4Vb9PReupAQ2exhbWB50Rx9JDXj7GxEZTV+rlHXyXd9vX/o+Euum/C0zYi0egFcV
Ct3UqSGrmz8CsTNJ943qyyStyXJSJgPxQ2ENY/vnbv4PcyeIswv0YafZQisjpbeV
0RZb6RjN4O6IeHvNTM55EPAIEFuQk8TlZwmoUxFwZZkMQqQBCGhaH1ozSvUr2f7h
qyvH2C9HN2M7gQWQjJTQOFMfUvZ3NB/7wgiMs3XGQruO9/okG3Wrx6/KMIsAi7Y6
GvTmFop4YvKoDqNupJXoqFzf0OKUqp8WpkDQ0KJsWtGohBRaNJHCbr0aOW8WHUn1
sNwsziGIpfAA5Av5ugNIgPiM/2HvtGPVXsJCnMyWhHz0C32LPKaRHEWx00j/WK9S
wcf2VUU+7T5PrFt1zXSYhMkFKt8z0LvAoY8gjhKckyO/YhWUzkqsj/larZEq6xa9
EIvhahkFFSxKl6dEGMlcnLSg/B+9dN1T6Y1XfhG6pWNdnc+ZRnVnetJVzLTmSJcz
fU2g5WyfyDcGCQ+NE0NXYGJL1MnY+etaESftVNGruGZnDrLbdRFnyQcDCZFrw+GC
k3Qn3E5C8AG73WQAXQz3IrsXa+5CmZHusee5H0de98hae41PsT7r3f0errLWPk6L
0+VO6/2tQruUvSM6mIiRRTAr+fKPL7CPfoYSUEdVVQzVXv4V4bwPdkIIdNBb3Vqt
yXdkVpbZGvMPELvTxt0h7qyPpZ3ELPOSN4s5+w6tjLus85eAT0XM2yOvrjYg1fNu
XTS5VdRdvsj9U/RsK1hrnhNKcyrdgzeRHHniQcW0t9V9MgP78uJFDqesqOGXBWdK
i5JwD/z+Rz6jJN924DibFj/Fjx42a3hI47ksXUNS/nwurvTnWJikgAnFg45MCIgr
kZh73iHLjHCNGyoaEmOXQK8DQFG6U9GiJo5UvbhNmO8WKExG6prE6JyoQLT8R+xM
xnJFezeVLuRB22iqzYvIed+XJnvMHOiJWKgkygf7+QRvQJBNK3FJwa34la8PSwIn
4VuAXm45rhHTqsr0xnBKwtX246vPciX7CWo0ju4Clb63fLYBNg1tCVCoqZGw5dOh
EwMfMhPNxCZ8gmEyBrdC7COPRDTd2oUccMJ7xW3UA8Tnt0OZPF19mqCCh0JhbK6Q
cGj1K/UTCeTwUEwjqiUSw3xOwIAgHH57tFZvXkAhgIInO3ikeo4fa1mm7Mf24clX
F+d8K2pnKtZhJaEfSK2Q52KvHYXmh3xABnHs0rofa8QOhaf+mTdVlFmt+JOxCyVg
vXzqz4aez8Qr+gop4hkcX/u45U5kAlmGQvTdDRqrAX4kTvJ3Ha07uFcJQ7orqH18
lfECzB31t8VKVFyrDwxbcJMnvnG2S+Sj9ZzYUSI4E5L//Bk6Mx8QFtOAlB/pmopw
zltiPvnnoByDncdLYAf5Hkwzi85RqjHhkiS2kJ2CFZbUEHCuFlhbeJEF0umIo+1f
d64aS9zOTDe1Eq2ubIQNbBxNdYqHrU2ov38PFfwZGtAoi1S3N5V+d7wf+wJdBZKC
h1kyVj/wUqP57TTriT0Cm7qRR5TtQ30rhjKdtGlwF6yEOP/PoaN6GcZ9L7OAfPok
PBnHNkFHp4/wvNoIXzohFIotoWyDkmhpdPiVX7CkQW6iHQ4jnE0qMT+cu3SBx5T6
9sTf6lc2SS6fz7TVjzLzMA64/yIradrqHtYbCpnnUDfUF8HtP8V9fle9AIjMWIXC
a2XXXyy7fqj58yLijOzkl+ZyNHgqdV7pytFM9nkyuRmtz2Z4Jx+zYXFeR7U63wkS
p1KJEQbSs/fJDY+pAEu/vjHcq7Glmm13dsa7aXgZ1Hm0KAiFqEVUeykdH4VyaYvr
gCdweOdc3KRpSTEXeXSq1MLO3l1HU/PIS9tBulLpBgncEK9VH4qNaXzegiBVarcz
z6pzefhOa8vbROsI6VbNT+FMaSctRy9QGVmEkpV9O6zJ3Z03bxqkrygg1iP7g9HG
SlogsTMtRH/ND1NDnBAX1hsLXH52Rv/pBvFeK5fpzX0vD2EsP9V4Ccw/xrnW3xJR
pz4RMT+cTJD7TkE59DsED7e9TGCmfTuH/GLbOuTj2Yl05s+RE435SzkA2fUxDPbk
TyD6+qyeyQoPRweqwBI/THlm/fMtIbehqEGxOHaw/YD6n8Pix1gKtqExxN7uihnV
DoYZoQH5B0aWTpB4KxpJ4hQMfP2zQF2mO1C8SF3oIoiZlvU4EdjozB3QWkFQb1xb
S74uZklO6FpU07lh/2r0yR1VuXB6wdgQIcmL0H+30Gz0AvIGjA5G9G+DuY9Rx48S
ZdG/xfEpASmUqGYCb1JnQMEkHRBF13toybkS6V3oO8D8QEk9t2Mu+L3EFI9l1lHL
xT6/YjjpnRgKmlS29Czl0RJRO0ZALxMa4MuOhMuob4PfP6ZhNfriH44PxmEeRxSr
NuOPRpTDv6IqVK7oWgCDH7LQlLTbXg26dLilo3EumnYr9l1/rx/KcPDOkiEe00U8
yR3vipTAbgDN9+6O/7xix3MSXGsOJ8xcl9sSSQd30vQveMXTciE5BiO7MxkeeBMf
awIOQZg+RrFM3ncVDok3H8woD6w7prEDbztUAS52ZjKE9apI9x+njl+FVN8r97rk
d6lRxySQ1F38GBOSI3vLt/tFnyf/p1kAZrcNEMdaFgPeBIZnhZ8eZ9ZWkxaF/itr
4qDupssqxi6ykhwKk7lbAb4Ur9omY37ESgOVSBKAPaYdn+nlZtrlC1earE++bZYU
w5p+Ay91az8YcEKa0a44hZbPU7nqWZqZFjNIeReOWaQH69jCYqCfL/MX1x4Kv7LE
qwNIRwD/tzOJ/htNIUUV8lrqL4s+qzCiQUy398fCuRJg1r7Ah1OWj2Mz1gGV2mMK
y3sH6UICjg8HK3L0SYHOOdVd2UqhwQm9SIfaKSXih59OBnKuId0yVeZ2od7psGwu
Cnk6OztIXBSKHowhvfR57vN1g6M1vEIEf3d3Wp1D1oQwC0d4x/gVMBD/HLnqbE1+
xvP6763TY6rsnAXhZqEiZgpyNb+LZ3CeHeAZL9gWBAxLeOYJuIR4dMiiGbBXqt7P
2LSWFqHbPlpw76WAGw2RUJfpjNPkRLqPsHSuWvfz1YrDiK+wq71Sg28ksqAceyN5
QJ8SQi4djtXczdREBAt/+7BfFkp7VKRCKcnpCQHOKik0Dpl4SDcJBALbqLz+aZVz
L87yGdiGX71TlYsRXy//s6edXmjmVsCSJ/+TWQtTGnftM/qd9nAjxWfVu9YDy3I8
ThlGrHi8Ndf3L9aI+1HLUtQgvdXrsFlxdyEN3u61OEqtvHjiDGt34At7gad6Es6y
4IsELcd+RUmgfjO4+ajGW2+UbOUq6GJ+HXKdine+dXk15TreBjdKbvKyBx/Zw6Rb
WgTqKu8KhhWMWDqpenn6zL9wzMazYeiunkQ5BY47l7fcmqPGjg9N7di3TXdI8PHT
bMLVOKS8Cg948hb+mq2f32T2cpT9tv3p8VUQHvVqfKLi4EVkKvvIPgHrvTIbz2eP
aCI08/iQnWHlWS1bHXF6IRNWzV79JTnfhWunpNTWYRmAUNiJSeJJtTacRjU+1bcW
xz6SSPSNtIE9UGQXgbJgXpuBsrXIHJy/xx2plBx72PZJM+ueaxnQvhJ7iUVAnStC
kiCGbEAGS0XmM3l4kJ7n2BhfwjC1KqHE+h+P8z4TSuUOKq98gsKIU8gLaSNI2aEG
oaNlMjuqBQngtr4Zf2C5HkIkYnpacSrdxKhkh+M37QrC8vsUBroPE5JkcH6HWSdV
V+FM/GWmrbMO8KhdL4+/u56YcFA1C2mnEdjH9ZbHx7QzsIOeO39hmkk1aMDD/w9d
TSJ2eYcmc5V8KhsVU19Dpb4fZY2DZARfXMhRuVO2rA72fiNFLaAHebflmMAHjeSw
pEhmGLwVnJC/eL3qjxDvZVBhKNbt8Tme/T0OWdx0c1IMJoSKvU1uRFfYS3gY3sJ1
jHe19IqW+HR26RRfdYgqfeoAR0sD1lGaVKVbAFzxkGIaw0op0xRJr2bMJMcSWLed
m3vW7rGT86sHDlX5llZsoscp+2meGxZTWgsr+2e2vX5AJjNv+wdPEcYS4Pe8U4MR
BS4fKciH21OxuXfCy8XXamRx0p9YYfyrHZIdKdj2Umt9dTcAw9AVoirYodHbtvEj
yCl8Dhn2/2tNUSmAhSThOBQbmaiGRrIh7OKIvAkrS0Tyw+w1g4jxMx1tWKNnr8c0
BtK/wY1dzjnPP6Qmp3HAg59jR5QpahTlB6f+h8opw+gBVd4DJI62ljQhTUd4qW8e
ghGevkyCT2JFEz2D2kJ+dF20l4XF6wGE/pVE95aWEI9ddEQCvjtb2x1FBV4TyOqN
SOj98Cz7qJaINwml7eWxB7dGuD1/+0qAniDa6z2BySR8Ux6z1oPsziQ3Iep8LlEh
JWDJvEXN74m4qFL0ybND2Uye2MukGhBsRZ6POGqj9iXf77LPZWti8rLXv/Gf7Bpz
mBnhh9ip3SRsDKADs5valIVOzAbTSc6ghfrEc+v7gVJeSoJ3FuTfezpO66dN+A9m
5bk79KNRbaT27D3DtVWd/8q5WSCFCDDwZ345OXYBvbuWar70G/ugVjSi4BdqVFj2
vGKRSkqqhS0IP251mkrxzJEsHKsvQeJ7Xk1HE0/PtICvpmeKBerBcS5W2BEk9E9/
rf4lRSMmLRWA55CuesFW2oJJNAuN658BotfkDslThvO2wlHFbHcj/mFNFvmFhA8P
Goq7EDnEOjvxqKIYeTEayWz2TUmQmp+GdrsF+3QsO6lLMJ61DRB7NjKO9F13+RIn
npYhc3nYnOHZa7hyBqsgS+wSIlmvgV/GAx4SERa+f53JWT/tvUlSJygoCvAidBWl
M/mPk+uPVvMG04LcWPqeDDH80ssUllzGcZTwAdySzIKkm3qL4hp7s1FRejHMd/Oy
0q11tdNVjqFLeRlLWTCX187eQGPNMspAEv7+dPO7W7eVh6A14ZA+psW6fOZb/edI
U5XjqfOiWPLs7fhNIIAEwqKSDBCwZ2aGaedVhDm4Njd8oEtjqU3YZH4bJq7S75rW
N8c90jJFnGxB6zK2WratV2c+bNlcnNr2rXtxr0xGtyCLpjXMs5Hd0yuzKXrNZbV0
Fhf85k06g+v/8RJ6RIQHi/kKT+FNof2nJGKsNcrIMlsNZNLSi3OFGuzysC/nxrRW
74dpU1CyyUKrArBb4840NjNlCz1WSr7wuvyDmXLskeRWLkQQNEOOiiAaQb0cMgfM
ZyNEHnByQ7+QeVrNAE9my9/ln4CBI9xEdQ8Hasbvr3HMlHcg5HsCnzNwkAwVOGWq
dOiCKGhX31I+RwwgDBGKdHdGYFmRiuMN70M/c3/mSwHabJsHGvknISrrVf+bkmsf
7EsX+dXH05AMl+zybRvTLkp7QK+UF+GUKu85ORnOHf2rx333fhvlWkqxtQDUzCOZ
aZNeF0AWbx5XOlqVU40s9PfoY2BknqD4doTRpIJ6iNtJRfqNYYnKV5gvg15Wz2Nt
gPcdnnG8Rz6mFxPT8NdZMnlAA6MJzbBlC/5lVy8KJEPityfXuDuknLi8j+6OsGYc
VWSO+n+s40VnilmkHi89by+/3kpGm3YdJLA0zZ681CrufnutSJ87H8EUp31tJoO0
9CxqCDdg+HONrwD2fLQdU7GzCZH5EV1QGMOSmnOWyKt4Lt/QbxRQ8aFR+4PaEho8
lXEFZ4EksT1peSAIieANtuEPxLyA5ZEwOgHT8vLsZS5bUicUD1Hje/LA6/AfVlCu
tfCWO6almperJasN2iXjsbPANACULKUSUiU6CekYiavLLCc/y8E0zJjZPXXYcylA
VjNMG9GRU9lTnnnGDE6p32pwum8Xy4zNNUXOnOB5qC5GD7akdgHA/558ntrPnCp7
E56XPBksD618eqq/BXtGASMBTVM5wZk9qyJGW5h5jXkDQjRa0QDXMGc6eXw6UX6a
214aohvfxfbz2JLaGjrGrTqPPP4kQuNt5baWO/xgarIabR+Kto6eprc9qWHvceQ0
0esjRRFYy5mamTWRuuA+bXsgrhvMhcArcGzZ8esjGZzPOw3p2gk2xBqs+MZzrkh6
no9tg/TrAR1cZT6OqXWGJEfBqx61vEXHJQyf5N5Edrlgn0cE4D4bVRso2Fd492nu
a0zpUv8GrkVn5RK2NHeuh2R5ZdnoEwzWw9dLp6xhaunJCXBgYAQN10LfxuT+w0+G
iqPNqFvpMIP553Cvj7I88quBkB0ykNq4w1vhMXwAqHPR5KOpp3jlyd9JCTc3vUgi
O3SK1tcLUBZqNn9QqA8s+ekoJPgrZ6SuJb3nqJJfzswXRbzFE94GSa8usxvtTcp4
ijodzFUBpvjrh/I59eyI62K+l8tm7Z27DG5wIcZE6zUXP44ZsNJekXOLTo3peUcA
/3SFqf5LnA0GqAWY09CbEOYNyGR4A6flBIS2iqTp9JLveaCHvrJsxTR1icW72iq9
5wLkrge8tz4qVCnJdpOT7HYlNZxM73oQUop89QAYqTVfA9T1rq8jutTyE5CY01tz
e/Dsul1rPzgrwl8lkZ1NE9+cRzTqw6QRJyAHXuw8Zn9DclLtaoNCKqdzC3fnMFtw
pX59BRAg4x+e1S5rsxqBLV6VZJw5KLOycQ44zX9S2o2YXe/k3zG07PNhXLDWnAnI
gCp+syKrAIYo4/gbJROTP9QC0hPsbsLG4YQ1W88S/LQUCMkRvn/vFdXU9+oX7Zp6
E0+sO9odd4NG+piIMm8F0YklQ5CHgRk0cfzRTvSBOLBqijtHYOw/4LX7MNRVkq5k
zDFc5LzePkfz2PvBUfIBnaVJjkacTdYAS6B5qqPGzEPgJ7mDkqOlqMmtY79WnJRy
6Adg7idW4ijrzX/MYuHl4SaB6PGSym0KFS346WZXBPRBLYSOcYUB1zz41x2T+Sao
JF/k8xrnqZQdiBbGTwFU7DWAnxkKp0cyQosXpPgFHqT1JtMhl7RZma9Q3SEK3mSd
JxlsP8XMnPcdFOrdOI3ruTz000msmwoic6ubd/DgnaRqqn9nsp8VqnpaULL7J19P
/59lSc2bcWv8iWlwGwTkZ1FCsUrZ4TzuQ333DU7y3MOfH8qk5rFyQ7SdbiiLLlFx
QBCqA3WK2BE28gHBRw+jtkuGbhiGaCPmU9aTYVvhdq1AUScg7EYDu7IS//gGAVQw
sdP9xLSpPwqF6C3bg2d6oRYs5kTcro7bjgt2akAwWHXF9YF3P3eSy6XUbudxqNhP
+VnbvyHCopdJxi7JBK5IWKg9wLEZCewcSMSY7b9/dUfdE4lSlWWltmK2B4JEUAsp
1sE70+Csw+90sW52ZjQNNDLoXp06DYhuuhjcERJSi64/6E9GfeDaHzgwpN6d0pKd
NKS7Mf75yOihnnBfTGp5T/A6vkgKw/gKp1EM9YfFnU3ae1i3zdDyO9os8lDpP0AL
WM97HDTPnWo+BeuTK73frjXuOx41hHZbBfdwQUwbhtuBjpZcI6rgfUMFW8TIyY56
x/+8bZv3eWL4x4egBNiMJ8iC8LCMvRdHRn2NDtgwLVZ8AMyBkHKgnrRXylzrEE+n
eHYPAGx3vowqyatl5y/VsXI9kgSNg935xVwXiYsjxogkXmciJ/rKqyPHjhwK6gkA
Xtd4vO9nXTaw5Sr6sm+CH57jJ3j5prFd1JFJagyZb0QJ9sHxYaJN1UjJMBxMpjwI
7WE+zUIgQCjQFal+ewpkfB1q1htrgrnr0k9BPY/cE+10g/PF+EIA5fLVKIbgoXyb
VYFqMe/GBBTkCLffzvBKMG+BmpncuwKNqM/NqVqwYKC72UH6CgPIp6z5z0+sN+Zq
VRzl4ZE8al3x+UgIrMOnwzLWj7Lr1CxNpzLzF+0u4/5GwL4oIfZLrUsy6wvLDgbF
pC6CR+ml6ZWlXusQbfTMQQiq1cEXCDHoVqyMoO9QDX9pn+vz9/+Kr4XMU43MIurB
JExwv4mv3tzl4ZOLWWQ+YatWy1UL3jx1N6Mw7l5oHmVOJSwSVcMYZIgSnSfIZTU4
GzYLpL1GTotlA6Xvb//9+WUoxB++r2YubDRN+bWlBEMu1/S3Io0PC4FeoyChFrhm
w/J7oA6voq5Q410oDILOuK7rHWafAG6IOsJ5HXZcDDwuqH0EaS0tjmRwwHVChxZo
Mof3bz8lY6eHl6L6d4znZz5P7jb/I6tGHNbcfAmQSFCux8d4w9/bPUSscCbZeSOZ
jDvM2JkMa9DqZK4Wh241KiRTIqg3AbV27HmCmyfn4OXRORn/n59rYE3gFO1t5e9F
NcAFfhR8BCbTv8Bnt8gwYYHSzgJhk/H35A42fSGC3MeEUS8HbwUiEY4B3kCaMh4g
4oTm2O4dDFY12toP27YR83XQ7CI3ITPbPO5nvEYmMKaIKZ/dfCbZx4n0j10Mc4jv
8dfcqeFikCvDwR31SP4qzho/3/+va9+gbFtXWAZ87jH9x3lDUoYLcWYh9S3Xv5w6
glRXJ61tJ0tLLQ6rYM6E5flEwOSxwSYTsl0OFM+lfhwxb/STzaC2d/o07KnMKE/0
f0Wr5oVKYCyNIa/cFIWA7YSg6zUxBeaRH6mB4LKXO3xq5/RO6KsWSBV0pSRUSxwq
Vv6C+69h7LUcvOVmSFqvnoa9Mi0tjRdc0F5bX2phibGDZlGev7mX28jXBw6GKzT9
GfJ0E6RL/2jbJtlmVRQkdV8y+rBRfoxFOTwawvTFO8xyeaAKVxOprR9m28g45HV0
TaG7gnBjGfsXJShd0/bRa8qM9d2MppSyuI5h/jcPMKCS42Ved3/L2LwW89L6XR5l
Lmd+eGGHTZuwFmeVqFCk1CNTqJoxyZElg6kJBIdaDNQqdvGz2psS6oEkR4p3s+Gi
czs9MRYT0yE5VJbR7H43kXREy7jPdMXyigNAwCG6SqfuG/ANaTjB07Imou8qd9/G
dKaEIGWYmPhb7Of7OzRCyHM3fIvPD3Il9/KQvMgFdXprP4GIXtHA2eS6mB1Gg1P7
ER4WUe2HhffZuIX7bJn5/gdWVVhS7+wT497DVa3Oa9YQbkgIsq7u5G9HPmQlQSYE
0LVdLySo/Hf3wbOHlfZYaR2GslQxNg/A1R2C5PDVuB7MODmi8wZNkgzYfWCq9smc
9qLL23sSkWmB3/tjzAKAgre2UNEpR0yaU5YBi7Etr5mxt+I49fqTNdfOoEfahkJb
KfbInuzkAksVBG7K9y+Jap3NsyJ+I+z8+T2MfA+ctxxdIr9856p8fPP2VANxt8kd
cu5BZpKV7vpnukXp5UoLX+3DbjWHT08VFXNZxEsTu+nTLSLvnpGYtMtPoXRlBBqi
v48mTBa2luKvumbYTP7LLj5CCyHcf9biqFSWU0IE1BqwHGC68Yi8Vc6MNBHyfxc9
y9tw7iC/XbDGCNjW+tM5vPiW1CeG7UEqgQAM6xai0a1hPGgwyYmRK06a6HYxPm3/
rkpa8uZKZorTMu3BFTRWCec2KNudYyRjiiTwCvbLU6SMiw/n5D2olPCWwL6IvDal
mjCCH3TQGZGpGAJoqIySPSckPDq5vsY6OHiYCY24NvJ6HyAE5LV4Z6EaXcglAoKQ
FVXnk46QsQ+QdYMRpNdU/Jhnkv722/0I66+3Ejc915cKm4YXuRkLs5oKYDVRGRLv
PGHMWf5VNYIykQDh9YJfX3/HwWfqEL8nHPbBueIh2ngOhmiy7M+Bt/i5y8ddxT3F
k3rfGIQM689mC80GwwpfcHdczvPtlDNXu4SjTnuRVR4cJVyPXEMleeV7tiRkJSkr
n+q57crTKCDBXlxpxApGvw+68DXA54V1wsIM4OKybWpFhqM9k8zLCeNH0abv0D08
DycRB4nZX3AnhUJVeGajyB105sBuo+5FsKW9Cqt/xfm8QpgwSqptCbp+yYkLOLVu
vHDGgER1ILo/BiiQek34G9Kvz+RAOZi0UiIIqXwpHMrNDTEwL1XHnnzDzaMb7Spu
eTjm47rqTgdZ8NFCn/YRb6wZyet55a+zclayu+eE+UKDt91JMkiE3ykm2JerfN4w
nziLJdvvZwVsagZe3p778pt3UCArjKlhQWaKxYfSXOLBNfsQICMIWSQriP8KUR1m
nsypSOYnQeKJa8PNEVu4TKmZuD7+S34KXvugOeZG6TWlvVRDs/Jbmya+t6y/BZ8f
4qBVB8zGBlTtfJR9TozEYelgtgUGy1FZt6+uk+HMSXUwi1l4YbFk1jeStzKKaT2r
0H9L+hSfKWT2IXmK/3KuE5/Fjm1Q39+vhQbk1J2WtZK75btAj2f2eyhH0EP3OPTM
B3SfPBZs6k3ogVHVKALOwWF0kPILVx8VeXr01aJrgV46dXXTZnocqe4DOKqZHEyJ
ohSwx4ZQy7+zDTSiqPXowZJhVwPD/DgS2JpGN5GvkdT+s/K0bwGac8qPt0ecJbjw
sESY8WpX+gtXd2vrDucmpbf0o3ugCX3nVW7Wo9i+y2YJqS/po3jgTyxAFG76QWbK
ALkwND5XPNCpVjaY+LfKEY8DLuDMzZxMiBorMA1YPn4crHP5RFJOnjWWIG5YhcVi
HthqlgIGWI5q963/CH+5ekDwXaibfm7NrVlyAnrErPGvHeF6PwahZwc9XNlt9K/F
1EOEgHOEHvPQonEhN6rCMMO5SjERXe623KAyVliuGdAMBtppiYlB2ow/GRvYnC8b
kJFbgQy7S31w6IVh7UqI55//zTKTXzY6xICk3mVQENfocfYutV1vFtXfZO6/gsrU
1JpuWskguW0MBdPhUz75RJ7rxW+b+oXDFAFPSsEKGKb0xwIWyAeqzgcQ5l7RAFAB
9aBNDJLfIsEiw+4M7GBrkjoojelPFq+GO7dqKAcuTb+b88Gkvmreog5zAErVBH9Q
iDXHzX5sUklCCwISYUBXKhBT94Q5a2TWT5jX8q7QkSai3jN2AuUUnjCjy70nF8PU
t+k/rcn6MBsHxKnI1aMb+y+hgaJ184sl8JpGe8WmsEnsV1hJcHPg4qTZSOBeKPuS
x5KjDavSRm/0fHB3Wu0iv9eVyaJbXFj7nzMmu1QG/bi/aQq0EUsAjf5S7vhDlUau
vtNgZOWv5XtpP2f4HzvLY5dfBvC9HM0za8ot9Wr4N5m2kG9DoNGmaH5EL81Bj15/
K7uZrUGSpITJiwzJeUX30Nidk7y8+0eHblHeiSNN2atwygb6qShFfCj0xiwfynr5
5PdyVv39j2N8Q92bpO0EcRFh6c0eZ/o5xW7JRhwGSZtM2azpjig8k5WuhIH+XW9i
rZCipo3gLkJN7gDqpCGt7wIIFxCnd/3FNtZJeE1ruPMomhbmRlG1Svwrz9beXRZP
9bxNDaG5ziwG+ajm01bMV0lwsNahldWHiTmix6Mcxuaazi2Tyt6nBHHPiaKnZLRu
SQtl9lfDGGF4yoAp3TsWf5gWDiUeavvGoCsVMO5DzR1Lgzt8j+s++DYH4fUlqljh
Aa0DRd5bVciHkW1Tr2HUp8dhxni/erxKsxqxv6zcDiWSzZK9qjdWLOSt04hHk9n6
xe3jGq18YbKmXAWfNUybIV0SzwWNsRXKiWfbiCGBj7X7tAizDiaHnEOxU1k6gbWK
uspgyvEI6GFzrS/fncQUTuuf4TIeyp2E2dzMccwQK+ndssC/LDQCS6w7HbpIqGkZ
ueuha5Af+dlXGgPUg+w67rPr1XYPvG7DpnCBidrufj95tdfkzLohvJkz7Z/wbJ60
mw7il1QJZIYX1rc8z1F/mRhGqARtxU/b9IlR7osmnCRIZ6kQibkzj4/XGYgkiX7q
9bc4Wtlz+npTR6Rr073oRSq8cJdSYrXWOu3VfnRzpjOCqy56e5Eb4x+FepGgg4uf
0NdTbr5EP3JqzKguKY31lu9v2GAFELEKmAjK3it2n/oL+sKUvc0sdQZYWU15f032
KDPLatpKZsoWYpj/tVk4peAJ6NevOw1Wbl1Z74BV0/LmDYoeTZar69aSomqKBQXZ
RvytWJLjwrWiHB6XNn6ThWR7USZPHEa0hdy6pI1SpbcDYeET11/OT+zlBs53VPS7
rFR4fPst0sdlSIjtv2p0XBcRldE7tKkt+gldo9PQzS6ARBHwQWsCjyXYbGhAqfYs
P8eoEhkrV25e1xj/GFckoHqlVFwyJ8ue17tM+CKKxIhUtZv0UIWFr9rE+ruRg3zv
I/esxyhLTU98453/behCqVuoFPmzOQRpI1dH+NpQLRAaRnPny8tB61vux5CcvRh2
XvxX5INbV9G9zQ+7T8diQ2/UJCnZc7KECdYyp6yT9G3nTJFtinjSvy4sQR77ZW7A
5pFVxFk37O0rPvOBMeRbkS7SZwPyhye+NUNd2FcOtfFRcW/D9cNpqLKN5TxenQOp
WhtWy2zzHb8A0qkeBVMwMrfgBHeXuMII8PC0X1rTy/OOKzilVRTt4Iz80VqGYCvA
Hq03gN06wFS59pkiDetzvgRW2le636oaxskB0+bgHKlwFxoR1+2hSxglhFUgFYvB
BQGIbayMd03ZbVgk68u0SbYkriFOnTIDCMq2s/a+Wcy4DBSfwa4aiQLjQY1DCXmf
CDHoq7I2E6iRsg+PN1o6CLlMDkTqkIt36y0jduKpMX6fnIm/acgH7kiN4LrH/5DV
3GFG4SCURCRm2wXa2UOkOFNTzyJQzQCnN7BzVkRozkg2yOOyaH2RXIKrRkTn/QEj
qcvfXmx9CsTUYj56X7GCvbwXngI+DvSNHhlIxpeJj5GXxO/C93KsmKiDBdAZXUHx
b021WN4j/2ZYnuuAVyvVStX70Kf9MkpPd47l2KAY7GNst72FGsZxrIJqe6Ax/94G
NdXQRBFbGmwEIbsioVrJxc2kd3dq8auPSYS5qPGWUPBZnsDfXyemtEO8tt3Mft0A
x5M3oP4ybH43+OJ3LYDmPJqmR/GAbE8a3SM7kpiokRFil78omQGo+wiCavtk8IEC
248cTjjBSdswOQZgpNqR6XAyH01S4lzasTO+uHb0CQu/oIUp6JkVmOwv9ErJyPlp
`protect END_PROTECTED
