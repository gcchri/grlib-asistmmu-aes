`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twY/9TiwVr07jYt7QvmHY2Gm8lVk3130c1kz+U8NOkI4OZx2a2hPo16amVWrmg0+
LiKB1f3LetVW5tGeWMAwKTq3yZojX2fPjBxCc/fy50Py5h8CChIlwcbrqutPmxGV
v5wiYTkjno0OlOEP/MzVDCi0b5XSkJ9SlWZhpDw9QgWImDtiqa3SWvkdfczmu+wS
AuPyDp/+j4shrv3kCTnE3zZlkSaLGA/AWSkk2L5n7/4vMjT3c52Dqi0bO0kRf0yu
F0ZC1dPrxvm7490DCN08BoI4GsvC4z+Sz4NR907DrDjfpc+iB4C5QiZwMRilxroI
4wQ9Q1t5ErWlSD3NLqV7aXFz7Ej+8JP2BuxIBIy4MKandlAIt6NQP0VhO19hKSR/
55EWsulJFgaOPDTIT0VpkIU+AsP+myAKI8xmVIUUOYGB1qZvsvOC/vQDrnO/uhjF
cJh90JSqb4G90O0jXXv1YOcrlCZV3nFFANyQPWsL2YBgL7pN5uLAjuPUI/cVQvkV
Vos7eW86Bq/2/+kS3Pe+COObsfAvOy3qOjVpVznBNkir3jfSAjwWrysbbvY6C2qw
B/jfgUa3CxMtvth4AZn23dfiFmNqgl+WUvDYua8j9GgUlO3yDQ10pS0+j2g1Y/WW
GVXvq0BvXIuaTwZ8IyApYmt3SImO4PJQe7r6snhcock=
`protect END_PROTECTED
