`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bl7SDJJbEOiuicv9IBSvIQODIGts70bnF42+CKDdrqV80JFOgZ8zQoISTdG2MwM6
1h2fnw37Z/R7hkY/JP/sNYxD0HplyOdEAlTp2SrI55JefK4OjOhv1dF+Kll7qYve
ZOe/ZSKajlDVUCJE0Z+JLxKpUZqY1HcR5EHwPtdicaH52Sof2wsD9BkjswVDLhFi
smh+vaxUe2pAMXasE7v/q0Mf3yej/JSP7MlwUXbR5uZ3LdmER4MEkwXRUaOgu7xY
R+GKDW/b0oIJvcaXbvF62+KAFrTlvuuIHPB9iIPQ853rMcf/yviLHrU7rASvCjTu
4UNzEy+XfF3aOu9w92zk7YTwXs3sJPAm8cxyDbDwrMeN5ah5Gb4NFreU8r3B8RY6
iOBXtDN2Lzb0xAd3CmdNUPjTaDXFBVB/foKxEflDj2fiWwz1dYHRjU8xLKtMgYhG
nPQkbM+0tvm38NQQhcqzwB1QIqqX07Igvt4j7bdR0v1992u3zDCZ621pwqmk4ygU
VbsUsXv1bqqOwm+gZKC+IHVlIEptwl1YpEvnzcb4ROFsbX+EyUTqzz7pQqvKntBK
KBqGIPx3uSKUzhrToQrHB5ISrJGNkviQ8StCJ+Fg8kxOe2Nc+613056i1ynpe3I/
1gYgXdROUnuTKGlZXrXES2EsAf8dWAX6itWeivjKxZg=
`protect END_PROTECTED
