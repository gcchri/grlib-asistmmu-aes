`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GxeXxrvZFEtHXmp7/zZLynrDZEoOTFDg3hZlt25Syezu3mYI5lRyNX1vZlvI+pdR
jkU6DLUbqT1W34x3pDDrkQGRGAzzhw8nlyQS4DIXHJCkbxELETFK+zhPhUsM0Je+
fXZbte5DteiJk0+XksOvj+0LdHuCfDXdHlnnXnJupJ5st6dY3Hzwsg9KGEJSXZUH
9edSt3kdd9wy12p1GRx4zAMi4gUgutp1tzVu6MnEf0539+809T3ctJWayVMpOtKg
8fz+Y3lZ90BfaBP0d+wx1tM7PIJgqG619G7e7x/VPJVFlKisICMiQxsO/RgTlabL
Q3TtRCIKelyfqtG9jhfkZWT4EDruHD6M9owV2VI5q+nnzREayu6yillCYng/SFzr
69biXajrrn5iP9DemI1c/U90W8waxLcUCSManvGwk5VMXZZ+TSWIDAzNH7kuP/A/
PnBg+SAQLFSJynpem1C6ESXnAKgm91pGo2ROlXcHMBEzh8+huP2I8ouSdOeGvf5g
cfm0bUNXBKGLNTkYa+zo9rrgw2uFLzOx2hRCxCqCDvEqnZYgK2LSq2S10HLeciFf
0MGIPwMFTD2UHM+0utf5ygVMNZpNGf45+avzT5k51OjV+E3ktGTAaBnE50AKp6zV
YreXEQZftmlDV/EIK+YbqyPXjXD1SsMIX65idDnBm/OeIoULLeTsvVAAyAIYnbXQ
L8QHIWGHxJnQXONf0fbGWQ==
`protect END_PROTECTED
