`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N5fZfX7/Thl9J4fBtARYVhwbPWSREAtQjklPwCWTx+QTsvu4kZJ3bEan3R5BKCI6
VZvxD0Fq3I2+oGNvuxDFExS/IsgT0put2I67GIAQriNQmfta1hGOQCjma4LshkEE
EWXVPrhhptmYaNaG49Rl1AJjWXsbuBa3pJYIfJ3QhBVt/kjM/FuY3oGlQuGfoEvQ
GdGpP695LsiSrNzyj7RfhI6v+qwkNnEr3G2fdzMoRpIv/K7OUWz+wxbVDUh5PuU6
wmeEJPHVH3apwTv0RDcZ+mU53vbyWbMvbzmzk7jwC6zxNrnRsi4ozi/BCTkEto+C
Z0DYWBBnRp9ug11VxuCZWDOPvlOv1YBu4gDy4F/uSC4UkxA0D+QZ8LhlBHwqvlVY
55phKbiXAr6ygpNzLcPAM/jC7QKzpyY6d3bT9dMSDzu0o9KpayBlfUkcteN+TZ7e
TC+wPG9UhJbe56Dtbw1XONe3Tt+kf3+pfg6ftC1uMmsyOLoPtzObGAXbZv4ZnOtJ
4fgWmhjLQtZngE6junw15OLE7XuEI7D1xFEMDCkFnoUkpCLTW9YYSOqaKFAF2B87
17XpLgohVkdP/FeySNA9QggQjCL/yQ0Vc+mVqCqzKgs4mTQKkpLrqQ5Dl7rS8wua
`protect END_PROTECTED
