`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6aIsw6nSmAbsq6Z1L3J8yozr0q5c7tkeN9Z0OcCfSIRrfreb4eZu2yaNOBna78o9
pw8xrHXA6UPiklUSYXg2PQwru8a64fLm0UJ0hiG/s+niysBI1YKARKsJ1JxEadBr
NqilctpreO7xntyxQFSMROXCPFdgwaSRZmLfUZZZZPrOWMvXvCmrvWh7zu6O8/tt
cx9ls+OsPBtDTw02XA2d8NzW6FobUg4ZpvDLW/qDWTTvbdXZN66iAjmXsy6Z46eE
OzRiV2Zp+GOI2In7cpIuz/HWdnEbygY1oZt3vDDujXL5LFslBKC4//2p9HZ304I1
Ea7X5zlLUkCOJXIuk6QW1qHrRyW+Q2T0E//7/Njaa9Q2JBfWHxRa90zMvscqkzTr
Cw6L4ejWiA1yVUiL4KPsTD55k6ceFgjlXTzt1a2ZCbTIiYbGgLaEZd53tODL+HDY
dmybQpwvFjIoN9+IN0KABnuwesN2qcZOA5MaMjjnNhJ3z5urZwLcE+0d+k2R+65+
`protect END_PROTECTED
