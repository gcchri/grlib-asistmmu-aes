`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hivcW8D+DMq+W31MPaUjzj61dcLNmTqptWEHLmG8h72TxuuudTPI7mLPllcPShrY
EHa5lvIScqeMXTXPLN/31AOgkXZRsDLPiMHNgtaS6jqUMTTdvc7pEq3Dhu/7ANRS
xGE6Mu74RRCQgOE769dfeEDnCnQRQC9W/HFV6iS/l9exymWNDtaT9tyUhnhYDs3Q
VsnB1B2wgl6Tjc9JHPugOgzZa6zoC8n4qHiOgXrapHnelJTv3L6M1lOT7AL/4qEL
WGV3kara0/qBpTNk6teD9uaf6eaikqptcarBbQFqfHw=
`protect END_PROTECTED
