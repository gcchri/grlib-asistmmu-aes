`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vWIztHBtIL+aAmGWkRfrgHCWhu/36CLIHsPkgdJeNsNqoe5ewPShjGWUgccE5gYS
nFX8EA5gctgD8MVJ+FuEQOcWqBDCNV97O0iRZVJZwSgmZUfQeojAf3Tx8aqMRh37
tqWJKqiwSGn/M+9pq9HCOkPAZTXSx+M0Qj4obnKZlq1fCF9nriAmAscVOsQapup5
8GzX07PDXnmLpvW7liWf7dW1JRm5ZpTp1fl1V8WMTBllWjhD8B7CRNDpSbGeE3kW
EtxS9PIDXgsOmUrfjYjwHb+P249eJfqhMZ+H15MUFpKJndkBeS7MEo1HnfhbhtDO
eL3ZQ31ldtif0pp7pToW06wu3lYysMLrBo6EqDsgZ030g7yY5tvwCwFyDea0/tPN
roYx53glDf8oz8JiuaTaL5bc5oBVPjOVZ+2uwxXrP21VS6TURMEka73XlfnPBN5Q
asu0etVjwUdTMKnMlky7rBtb01Zt88pcvFCLjbH7vSsbkQhlANpzxgspTDGV986h
yJdHBLglUMYhZ2FAX4e+M0uwpZMQpevLvAmTPxUlooddhGSXZm47SwX1v/YGvzbm
wL7YDQ3FcUbGU3GZLGfaxw==
`protect END_PROTECTED
