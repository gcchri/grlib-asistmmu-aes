`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwREkORgpSSZju2JH00Pl9AZ4DSyIBVuTcXCspe1yexDiI1EWTGeQwSiRGz+UL+B
dF6kwL1/rXHr6fShS/SrshhJvFwZ7VjXqJYm68nWc9IZwdLqKPZc0dwBojPCWWxP
ILNZzQgNqEUwkBp6LYuZew4sPlD1ryU+G0EETugBtAX7ty0rikxNTkqg6S4+xEiR
VRt4iUOw61It0ASFGU+qrnw2FBqZP1STGPTSsGEJxyT8RGAygnjaP8A3K+UykhWK
/QdN9IQKZFtBLngncqbpL5kQGjLy0RV62DgpjRJ/2ODyikrDPeYcbiphC6P0PSDr
HhJoo0oxqrTCL8coC2PGkizQrIGpQK+CQwp6MxSvwJYKVOVxppQLhP0Ax3gHCZkY
pAef8FcBs/VcVgMgy767cs96doRtN4H/EZP/3V4rU+1zwaKqEkLAkTEXho4g86sy
S/mb1lGL96kqjvJVQFwoU3K9q0wu0gCzc69JRVykMOAV4Ikc8ixcMUT1m7GmUVMR
CZ7fmfgLb15jWK2YF/kYK0q+lHPmacldEjrYoemcgdnSJuNbp3aTtWaylnypojKd
wclj8vNqYNIT7CTZdTAW3MrpGwtKC51QEGM/+X3o0TiyLgVlfjB4oavWiNnqvEvQ
KvCNiEtb0WSgX6DMXz/rSo6rPrbOOu07wvvaVLLoOH4Qe+/PFE+rl0bRNadTs8fC
WhsGyaN3U8dKiOhob2FHIC5JOteQPGaa3sBmj16JG5G74foUynWOAvMQ0C8hjA8t
boyXHLZ9u9qYaJpRb7hpAMtcv9EWo2eu8jk2F1d5A0FXmZpVX2207z2sOxUa+tvj
VyZfDuAynb2mOJzHYdd2fANZw3LukQPsLm/y0ThIGUIaochbyBzz83wiNYNActfK
uNtWXdYD/FkLg9HIw9zyYPECwwUQNBc2fOxBFjZnZ/s4bP7JopMa78TUQg9dQ2nt
Le+j+xcd7JH0FQhqEG0NHoBSysjkm5SsE2U3hat1yRNFQjiD8/BGbOYZTi3cAOrR
hwlO8TxHjpZfB+sF+cB8jiJChjazRoU1GjfQgeTAxNFgkxDXj6b30xh7uVUE4oy3
MCQdBD8LeUr9BlRvk/BOiKI6euQBXFsDV0sxDSUuLfeMsWjjLPngJh31nFYIvwnQ
WantNAUlp10tqjJkKnHKtL/6kq0JJcXHFSp2eL/Z/sT9YWHLVm1Z4GmnY61bjeoZ
XzF+f2Yivmpzm8jw1PhsiaRq6E9p7FMMQYpO020LO+1VDr2T2WpPMML0SjtGv9Z1
nwuWF7/r9wZezUMkIo3v0vomvOSXd9eq4IIlJvlfD2K2gDtVXX7PL1TE9UuhFGWB
AytqA7XFdojzeGoZoUl8pl1N02hYA0b/1UItes3Hj/gZIGymUoU4HDfyN9d1PwVT
Up7Tv1fUf+yr6bmgvmLMENTgK5udZX0xpiHb0bsVH28y8/Q0L227sqI3IqL59caK
lbkv/qG0H4IsfuyNC5QLuyO988KWDCrnJuEA9qQoDHecfWidWd+sjOhsd5SmK4Hs
pwYA4WoeYUfiHPjb1dVAvMUiM1z89Ou7nBgzCBhrW3BroWZ8ql8lP7mU+A7jXTwB
21ojiUHGxVYAw0XeTGxKTRp78C8V8NI85YD3IT8NFJIoyWNR/MPljTGUZSFCnh2y
YdW6wXYPEhvfq38muU3QS0bIDEsYYatupE3eaFmZ1R2nkF8dPWgLmtGvKMa5r12F
zbB4Qt4FmLzxlAzTXfzHSDrDqKPfAI7DcC5ZpMLjANzrW2/6FtnnPIKUnIQSldD9
uilMHErLCN8WbJ7lEoiZgvNROEy9gs1opYZU5AGlqAz6IhwcWUsE2jXvYqfrpdQk
QyjvsqNNOJjH74Re+EEEl3ASKoCZUpWOqCsBKbDAazvoEvVdfVr4jJpeQdqwtI5P
cGdondtt1S6O8t6Vem8lySSco/Mwdi1Chnnola6dv366q8gwxhD8IOP9IkR5sGRV
o6h4t25ZvIs7+RtXcqqJAlWBNzK5cCSyl40yK3ueyWQ6OrtwHcbXkjcSOMDsHxMF
8ESPVC30BTWONhZx5K62M/r1QbrW//UwXnaLUAsm5kvg0QlUS9tmev4FJvXDrvwm
GMApDhY9EddF+IqyywvUYvKfJj1nKjtvKTOKfnuPsVSuzne685vOo6ODyhUX5I2d
BO6nmvbJCYzEXGMrrkik8kuYE60+fSYvB5Slud0OS17gEaKi8ja7uRv+lfM0mQEW
DIa7ywJv247V/O9g59zuBwUzTlMvoqCdN0JN36HmdSid2/tamYiPqg+cATMmaWFE
8CpZ8Y0i0moFZNX7d/rwj7lZeon8W+WHyZW+JBccg7bY4G0ME9KnJNqj8BQHwDBs
fqIq+b2ivsuIAMN6lh0TDvipFGlTmxdCJ/l41JFEkSeUTpQW1R6f0+nrMPZaZKEk
tQzHC08zBecGczRUuv8Iyxg/78rkLO8r/UTMFQAISfR9RzOmNaCfsWP/QLZqj8oU
g474azbuWYEmzjOGpftDSxbQ8va1I5BKPbccXMhn+37qhHV05bWzCZ/F5Lla14Oz
qwykMNNxEniktUjCOFb/sfVxPPa0jsQCbEUKWkGjxOIbcok1b/W6Ggvdzp5kbA1P
PIPV77kZMQ725X1lqTsxdz7jmxl78Qdh6ZTgVDlb5lhmnctLyjKkxZICLNdoq6Sc
zKO9DgyVg1PEGLqYnZS2NT+PN7QDM6m8qC6NbsOyPBJGpaa5G4A6Zmcudzalm1/+
az1Diy6gNZuZO5mpcY4Um9LUzdjh6FDf+95klrJR2T2g1w2xbSf6mropRA2AAbMO
XYJchscT/BS98+nUqhQereCIIWXZqnzJ1M7BZQNGa657/evAYBB0oS9o9tq7s0y7
h6pllfjvGW4ow1nlp7mRc6xsRu602uRdBNddxvvuy70AHyK0bxtK5DGl9IHpL6fq
WqGZaAMPCnwzzmsdt3phsdIuv2oo/UAn9M38KecKYg8KRuoL58dP/iV71tXwRrUT
LWLKNCnhkgaAMfabr4fO61MRIjXAHKic7IcrwNBYfz3Hv+xe9Q4e30uMwJc9pA8T
Ym15MPk3rpE+WrRY1sFsMLG/JByEsoWmqLJE1xZ8MDhHTnzCK3TZ1I7FDNBQZyPQ
r0uUMOQCny+BIEcdIyUvvxhrSmggCMJVPfVaT8YnJ6rMyqMiPvIw41198YyyA+BK
DVBjzChT6ZrhEfsQ8BYh8V9wtbBoxPX3Sv7bH/GDugZ0E49sqvXoDSZ4d5Cco2Wd
gZZvIcgHJWmJVGmAUPLnHTFbC7NkOSrUV21xEywyQe7DBGwH1S9VY7viXVD+WxLu
UVPWTdSJJCdA1CkDSTyZl2CF6jGqB6iB1RnVB6qJa9WqL69Z2xqBk0PstUINs5n0
rkiU1+Z/O+Acshyu5eotiAZazOmSWKrCfpkHXMCIl+yk1ekz3/OGFYka8Qw6lG7i
QNu/1xZ0ABXlH5WNXkeWcczH3nHH/9VY8GMUdALNHZPeTAqpzrr/pHjwtBnXFYsc
XFj0KVelVQ/qguqKiP+JDCbt4+1cVmgNwD6fguE4tZuYAysdXy9ihgWYXK7cqmYL
cKjTQxAtNQjAnhHeJN7ehTWrCqoZXmqHhin00ozCR9kQ4qyielLtawynqaOBF4ZM
23nZnLOcS+o0rAGKb6QgndA8VNCyC/qK/RrGP5HQ9ly4y1eDZWpDu1XMU7x8+wg7
5trO9ogd1Hp6XhdLLTW0WBqO8mMyW32Dt4R27EcWdhHqzxJLyGFw2lwUu80a7+zC
nlRGFwp/WpNAY80CJetA1jz5kK4TWVfT8s27K32U0XO212jw9VvD2z1XAlhtITXT
wrf+4GzXO9kXlBXlaYa9vvT0rNt70NDw5b/o4VdnnfUJYyLLxwGzUEi/shZirDnt
m7yFGn+io5M+bj5hRjcoSfe7mMMRf78of2gYuPvldzIEdEZ2cACOTB40ey3je6Sw
wYFuHgjrVsX+sdXXwEhgN0eT+jIrL9u3J2xR+JeDhrPqhJqp9GeX5hbEVptOBtPZ
TrAtqSoAaVXU9t2XJ4gLp5K7SjJKfjJHJPG/XeNg+BdwRmycBUGyOiNTbWyiSD/Z
M1qKEdjMkDDzlL9qvs3Zh0rod2zS8Os1uYZWs/x7HXqiagJuUZiqp5DmInLozIvn
H6FTeFNR3eSAaG2DBNM0RZSsj3b4u/TasNHv380UZd499z2A/MU+lTEvWKjk2Vjs
bKuu2v/QFWf8I4KdITw3tUORO4/n0o7I1oGSkribjyKAEFQidlvHYFvnm9xyegK4
dKpgewdMwsKSgmEp+6HsKZLX57VwAVbXK4r5jCwsKslaIQYh1WwfCDv2rzcbRyEO
aytyQAJvQv2muNkmFn3sr1z+U0Bc+bCykC0lmSzO3A1UPVhBB66kEHPJQOtg8uHk
7GW11R24EWtdClGkmjsi2KOg21358oc2/VNo+c2byTQIgWgTYDjnXG885sQs8GV2
+XOiFuNs3rLPpSLa/O0e0NC6kIE/ha/e3M4eIvOK3SUpN7IDSKPEjPnoEOF47VXj
XnMciAKWTkquXxmFHRsyFLlm0SyPjJqMeSEB+TNpcn3eV51DSDwYtJxv12hko/9P
3sVVMOnyN4Ne/P29y89UPsN/ppIYnJgTToA1ZGOtaQkhNRcg/BKaeOP6cTbPCNwk
xxixmMxgkiv0ydwdKW4ko+YozAIANBaMTFIyvxIVorJtlU7mQS0mmTlJQ8nGwzeN
ID0bR3m99RAT0aRL6fSHV6FThGSB0+y2sGbkPBUNO1qcKp7BD2RxgvtcIKbzafoT
7m7p36VwRduZVZr3fvATizPKpAHBUl9vKoH6FcEvLwuDDFgfFg9uwcQ3DaEjr+Ov
qYb9ISCbPGzPk/5vJJqG3ICw7+x/hB/JKTiocq/pB64Olg6uyxa09oWnXwEZUDav
ptKHh1E1A0JNQTeAybLSNtp0A4HgWpPua3z0zFhO4aLbblZEE4YjqCAMfMcyNzFg
//lD1hJE1KHEWg+d6vJ5HtWbz4FSWg5JepihTRA2NtNSiQ7L5ZNQ3oterZ0SYcMw
Kusp5zYyBa3zmARIW5/Mua6hjUIh63VB6+bZbq/yVQlPqXVqlve7H7oJqW2w9u5S
xGPtahXOaSlIm/LqwbVka6ws3vknZ4TMSwt+/YJLQ9c6sVVxVBda7MptJRMeMP7O
9xLrwhJZuQeL17ydGJxieSG6OBfsFmWLvOF3FMCl8c43aaKtCDkQ8DzNC6ijaZMD
e1Bttzig6t2ZH9NT+wdPTdxWNmaCgOwR6OVipbXeLs03Bi0WbZLhKEOAcX6qme8+
tnsuAkv0O3L48tFfLc2Lx2uD0hF4Ir/o0cwCddaUcdMWmDxzFf/KgZO9SmSIiImQ
NCAku8byInKND+Lmf3WdRry1wpWPdQIUH1DDAbPq/NaO9vT4LhA7f1FOuLrnHWjk
LaEHTxRm7FapCacSv8yixdeA9Pqe9N1fJvGgZpZaVwKh5OxYvL/rSUfhxe5eYcck
rHLMgUs2QFIk8fXRzySP7qRp3mq1KCRuNaHlzvSG5WmXxOeUw6GGdnuSN6HqOxPK
ItaWZG0ygcyx0BnfYEpgsdUXLufTpVP2tyvpIWlywYIEBbLdFNpZpoOraGJrAFwi
aiKNtT0DI/bWSNKiEZTZsZKhvhxOSOprEXcRqSD6wjIFwM5q/wGYOEorHarfwm02
pbTuXssQ02vZ8XMtnSUwCal5W020M+74C502Q5PGyAs7X1m+GL5Mym+geMs1Zu1+
W288HYd3z8zNgyduW87JM4HX4FzxDSlnXFkRpqpULgr/BacHlF9OtVL980PNhM6T
AZ5254BPmODShoeSNFSwepzWyfdD+Ew4Pzyy4HGYUbgT3d+hge+8dukQfmJtPYOs
vSjmvme3VGY/vTI6AisRdKy4Qwd60dz1BRZoE+1eAD85tCPNIPW8JgL44Gmx1Gi5
IgiLdIp5/nDHGVMA/kYqoUgWtmjTDP7BXhjHiw7AL8LBJ5seh0pXrY+lAJ74Co/p
EwHUuy6+wetA6MQBQAXsEU7ThxKxEnAX+fzVRsVKpD/2hBB6ML3TRiAOL3mEiGM5
sPTgIjHJ4hFzt+mn6Vow8TScsZAEwloeYRQkUkgcxtDdZTzKwIhkHnNAMkIzun/a
FFI345c8ewVvVVjcB8F/GBN8/5efbIaLntAylz3EVALmd1XLHRE+aQXvd32Lnj+4
TJkXEKxA89yUsJL94IGwQhrScxOCsnTKoziOl8B76SmjzE9dNXMFPI5/Sy1Trb2u
kzSqq3D0q1I1C0/Y4soQ67al2egQsLXYNtSlLT3ouuKBPYQVnYLv8gt98K0W90bP
nDYcG08CS19bA3OOKnP1YW4a2dWHzFzayKDH4DnORvJGyYGUwBWQEky+cU4L8Y/8
ECsV/mtkDkZrsT5ia+SxQyXJqLzFOIrEz0GdPS1lZnZpXoAWYm6/Qx0L8UKWn9sz
y0ZJFTcqbd8n0AvumfwjOzDNgfW52p4v3bN6xWK5Li8c3QafK8dJFrwzxa495mxT
2/sUS/hQyM8AM+1IR5dc2Z/cMtB/bPsbMnpJ1y4IO6aS6Q0pgSXOIEnCx+NVlWas
T7xISdSa8d4HdV0aB+XdaHMz54JmhIGH2NqH/CPyYuPGS0To5GC6rwRTjz1Ar0N4
XJCEPMl6lKJgyLypSkSBWNKak6K+9BClkUQoMj3pHuzhhHQhZSlYx3mUUQiwED8s
3+540Lq5uF339jQET4ZHaGEmfMivoWDkDrtN21Tcx+/hhCmDSzslyFvmZGrH4syu
rreYtLgcAmOTL2V9wY1w0wqiIK4at7ZlBAGs6BTEXVnIflOMklWN1IOH3gr5T42Y
ub4DBeJ71tDsV3K3m5rIdyV/3jrUO8TCUOrjDaSb/H0iSYRwi+r0T8rVwJmQdF+8
E+BjY0nVBtSR0TNT9JKD01DV+AyAHWQXutB0tlr7yZKVwAHJs4i3ZmrUUcgJWjUO
3fQBrqIVUiDSPnv9w/6eCAFdL9J+EfuVUwhYfwlnwMctgmyfSHUYXDxg06EeZOfL
JXIhPF2pL+3EDpsprNDgs/2bCev3vcdHPmSTuToIKBkdqJUyuF1flAhzdHKL89Wx
RL6ohRAX41IKeLNnXKvbLjETFZo/h229Iv5ZxCDXOuq2zD2GiABN+ltl+K4a2GDM
ZShMRkS2guqhU5rZgKr0PNAfRN9msfXUI6BJlUbWCa5azw/UTk1fFbFpoqQw2bhK
nhiWDQqL0EpbQfUSHfh+opa2m50II2U6WhJvxgsg6/b7eklJ9vwwSinxU8xxCYpw
83vIH5fl4qsOCMduhogrNm1l3/wlLa1ZiKpMiTt/Kgeov82JcvihhPW0fbgeqJXU
bm1pQqDitkz9YZLLFWqKegWNee2RvkRGbQ9AjtaZ9M8wFYe9JtJkIGnaBFDXLQR3
yoBxtlGFHbFB7o45A0FeU26FfX2jlJlBjTULUYEkh2AyEe2Mo1QG1GPnOfDQ1Rqo
FgYh2HW59DxNtpXydw2GybYlaE2KO0UE2jGEsJXdYGJAEoWeAR4q2h51Tq8w4Viy
BBlZymGLvCyAPuRLYokEMLA3YU20WR9mNBGEvd5ovRS4GVgCRaahGRXnX7wUukbo
UhH0AQrrmFrNY1HYkP00V9GQPXDMLlUnfjH/8Mu+xxNyXdyl+Gzm/sciPGNiPUzi
BdXkXEuugSZ053hiNI1Hsu4rWwNo5XUNTaf/Q6L1wp81ZFQ9l0eWFPOPsi1qfKpJ
tjs6bwkC9yK3sDAS/LxWxFWE/6Zr4JJssJj6+aYoiRIXQOm9+T+pGFiYCA8+Z+zC
QJSDsndZgZTHXa5c/5abnQrRWJM+WYDJ3kCrLFttK0RCQilWhUjGAn30tmJNwjOf
bpPgRYF6PvSihZN7a65KBeuArS0ypBCZINhZPkC9dBX52rKdcQiCogHbTioyfBJW
qgJcoOsvU0JjQ+szToE8qc7gEZOhUSwlsKu9aZrLzNhR8ZBMyBxJFDpbHk8Q6YC8
sBLXHfd290VX1zIsWF/gGa+HL0WK1DmhgY8FBJAJRO7v5hj2/UZ5L2TN235ksnGw
R0E8qUZzG77GegVNUnWtVAllzUbxNTzu7nBJkakt3ivrhb+c6Wti++vmzUUmz1Qk
wZOfLfHqgtWJYHUXJbNPyAqy2sH1c7YztWW3kzEjE8r9p1EwfZ+n2mG1jbsjFeni
znGrJdlx8ru28AnXby7fh/zv4AwSNAgXRIhQEoT8biesquHYg4lhhgFKdrniCnZh
w/EKkipfAq0gs94P65Tv7UiUfk/s6B2Hhi9GXAU/iJvFjAIpHQP7A6nSSXYGCzcm
kDbn3mAaGlRO8MSEsplEakoVDQjauDCyCLIRfGhQ7TjUoPLr6mXreCr0+sSxj4eL
KIHr8dTqmJ4SedAbddbulIXyOgXwfzd3ssgJiQYfaVjm/TH/y1MOfGJbar3oUnBv
cH1nPlQpfg0Gis/85kO768TGLyzR48ZsQhutimUK2l3MrRkwU9bSzeNX3IJJbaoH
P9IS3q+kq37QCLtbifIsF71SaFgnYFD19rGOYSEDxEXfJT/hp1wxGyKEbpYjDMZA
kDYM7rlAbUXGmwT1xTL4UxSAKsg5gdm1EGkknxSbZOliyuz0+SgdEPaXU/CkRGxd
onfv+Le8JiH9TY9t4GOOJGZz7b+RviH+OCxil1I26w+9H5NFn/DQdzRlAZVptQ54
QEGozuJEf9waAEO9ruSbCnGI13JbP9fnWkH7g3mNz/B6+/9V1FC4nzhEzABuBONo
FNEOR15nZy88PJPBlOh/EflUy2gSW8ZlQCXDFh/0jWYPH/L8rzdYHBj9otdQsUxu
WdNCmhqUoDAo8NR/YLvX/76wuL7bm7uS3cxHOL0bRUCH8/j9acJGAsw6zvK9VFNQ
P1qCoYFYxpGw31TWCUVjYGtOtTAWPDWjWxnaEC3Ozde489nbJj0Q+OtI+RwMaSwD
rmKUxQL63gq6LZ1xn5MHcZmFZJQLbbqrfBYzkF5/XvB0e7hPO1Frtn80RdgsXpeh
mu5gUsGROoPh5W4fAq4pX82zwd4EvIULIk0cX9ChEvQFrJpn35F/opBP7fZKUf1u
X3Z7UavjV15G7TS/F/86l0HaXc4Oq5wrkGAs41Ew9iZW1H2Emix2z75rCDY3QLhx
WaVkO3gqbowTCWUfQRPxucf2Gb0GgoofIpqJHI/kOvWQ+/2d2qkNxXlebwila1QD
38/fr4Ia1NMM+luzINJ5ox6V+gCvgrsSTRK7O2f4+AmJvXVtP+Ki0TTj8bfL+PcD
zLVCkif1lrdl1wKC+JvUlOpVcxDOT+MYmLq9nML5hSMwLD7hDOO/BTApg7ieyqg9
IOBLml2gp2mB41xxSe3ATtgq1l2lR3u41akhyeh9IUJEVBKxFoO3SfzBrEZf2LMb
sY9nUXT/5BrKyjgxCqO0GRHlyRbwlV16C4OvzQtU/69X6758oNRm9QCrzX9WIr7Z
PauP/slx2y9mhrpfQbklkSmnkkr/MPwRtEegQMkHnBAfcOFDsAubrXmR7Mu1jrja
s8T6p2ek43hc2wMhZ7XQG7eCw8xfpsb9fDEkTcfq+ZF/oMJ2jL16p2UclvluO2pG
9Gkoz6iCx/f+x13KOxA2B//cNSymK3f7K3dwWbttqZeCwtTre8JP8Ysz8BWWJ91F
SEItWE7n69z8FQ9QswV6pUU9h568IiXkK1Ei277u6YrxtBOxRsI+VkOykyNC6Fc7
Vde55CEiv6Y7mjG5scLkKhwqoXDZqSooJORMFLyLW+xvLOejlnZyIs95J/IZMGJv
cF+vxFNR2WPjmwUWGuCQ18y4bu6uJombCrG+s/qx5IUj95fiuZkJo4b1D3RdvG6P
aabEYFRr7z18D2/Dx/YWLH0k/Gq2GLMJLr8vxIlZwXWBme60UNIKimNNv3ykNkBk
LHomUJSEhZRlh9ivD/N2lYKV7Beebp6ySKVTRdBYzEdxigXia9FE/aeKZsMhMqFv
s8PNxlDd02sENalIHEnFq4cM9+lT5C2biRlTax0PIYXchl7+Npg6Q5vtff4T79/g
OeRf/+Mulb4ZSP9FNm522sh933KChIYQrHjnEqVGd41TR7cixQhcsmrI12Z/b6U0
rVyUV2lFAVbnK7MhWaXhFzmFHRHTRIIvTkDbvVAaPMOAd7piPzGdj8o2ilfq6rvK
B+Xx77oXc1DIOvYVaYTLy3TMbuxu1G/PdKQ5rFyV6iBVPx5v+TPvEiMfL8qa6Hi0
LR31Q3GXZSxXRS+b4NMDENxoC4zqdeFr5bkIlATw+R0NOrqTXNLODKMI8UBjwoPk
ZxfpbAeUVoVO3vENGgyDW9Yz1sB/2/lZS3lu3XKvY5q/7yYi9dQ1XpZlZbNuKdPC
i06XUQ2m3yO1kXNt91RJ73E7iFyNPxEtgHYGYRK6Xfxi00M2b4tPik99SDzMKnGc
ucuxdJjznPOa6NEsc452kkT3Xh20/x438pqACmUOQTDcLXFXMi9ry7HrYgHZOE+/
7dyAX+r/hNauj8CjMDkrH4iX/iSxKeFsj8qrkOjGfznIWL7zzMs+QgpIGDINIkSS
Xcl9EKTvUhgWVDBhUAB+HIFqD0lOYYQHBTV8U8r2bUlGdy+KU319dwDsr5bMtLCU
skuadvexsx7xBuGi3Jhg6tj80EUAqXc+R+NnOHYCJ9rzqP6v4ein8fDScKR/fn53
3sgzC0b0XA9h6YOKnPVGRZpOH1M8PvicIpSlQ2mIxGCa+pqkkrEC4dTwMCACR1MV
p2sPgypbSmmiFnf0ADZPQaKoNJzYGzEanSPAb6Madp9JaAHI207QaNJ0cjZyjJKD
SyHJmVxDmM4anfXG5YZOPxGA+RfHg5i9IXNK1rFwe45TPhgbMc6h7I/Qd6sZMuUB
jYma4bbpMPiixqYAJRHuyuKT95cdpba/kfLznGhi5j4/mwLjLQJyHCZJniQ8Mj1U
TymeHoI+3yHpPECRfNt9x4mSPL2ijdrgGPi33hu/3SV9B3xx4yzaW+j8cQqGfDrP
CcWAVLARwF6e2wJXCpTg38/Z0SWOd9oltqZs7Wgq/sD9hwGJ32KD+UPONwwNFhMe
3nGA4X2XSiG/5KCEbgDs2eFOH3BzxRTQCp7Is7Q3C0DLy17xJenVicx9xKVl7zPN
S/6jtGN4keAE0N2A383ldVIB3jNKcC2wDkkTjyCREJzdWcgnHXy4kfFy/Zl8IA26
5JKHaRaCk0og9a5PF0HQJ3f6rIEvpgn01FUwiNQ6gQYJ0af8xHtze8nYEtooEtvS
abIeamCxZ8oFt5+q0qFjAQiERYVUjHzb4M4QWa8fT9/TwmYe0mE9SiMQiTsGR3if
d/bgBeE4aqJl8RnFZelKvBkQChWJreZvbg1SbFBDkO0F61q+vOMIXFkCZaknhW/3
TnBI/mAKLojb+EFj/iIzInAl8BdbBL+t4oZ7Z+KXGUgYpTK2LWma1suqgxBNDlFG
Zf1gQjgX+Cjxv+5NjBju5MgAsqTVRw8XVl3Rr4swjRk10mDirz+xMPKLx+aTz7Hl
vhEEpJ5GZyJs4JBvPrUTUWoqAfp3S2fk+XmzX3abNXPeFewy+Tf3+t6U0/qfYBci
xWcIMxAevT9HTx+lrOD7C2Ynitx5gX6G22kTZ6NuYk24GbGzqNybvmO1iYIpR/D4
5esWqUxT1WWbMpeLC7h8k4NjqKCruWNudo7ThCHm3t1kcXbUTm7HZdLFONhPI3kC
iw2n7I7pLiFoaDmqx7wW6LewSFaqS3a807WOADglKDEBIPuCHRHvEZGTg306skTb
b8mlLfokU16BTGgbp5uJ/bwKAsYQwwgzltg/wF+uvZt3uKue9XG+zkKBo8dJqN41
kRIDDBycrYJAO4rHWnYbSuMT2dQXtdJplfc3ufdoEvW4I6fH5iwvWw3mR0me+MmH
o8ED13YN3o3cOfc1Q/vUU/mZzCQhCbagUcAAbZTs6QETVejxiS+sH1FV/1maQO07
2S1XbLH1IwOCOdFzMN4OCM001kdzQ9feCvTCkN5FstGZh8mjGrkrBlXEonSZIfNL
gdVjpL74+NQxW5tuoLdgJfvokeUgKHhBWMusef+daAoITeF0w15wULvEzyR9/1xq
spHzKst9Poez6X0nDKvehnC+PmxmhVecsjpdMxu7qLiF/wdrv9NMTt6Hz5ow2oT3
Ii1H085Ik/BXSDzMFPQ95eStbCBAVLNSeoJNnpcozqitL/th3zaeCv42VF0WQ5Ne
mPWzoAFrnwfCWPqJIPUnYwHZ6BeHvZeNBkr1e48mykZQC97Jw1Tby7hOP07fiMLK
zmWcim6Tn/UE0KS0ytI5NRNhVkdnLLxKgav9kjxIywE3hMD8x+4n1g3qEII/4Mg1
EAIp1br9Warw89wYC2UPOZW3wMJiVY576RfM0vsmpPLudzcBcrvfwPF9+7al4uOd
s4jzbx0GILVEU/FXF8qEzd2A2ZUwsc8Jx19wViPMvrH68yn2JRgU1b4GOPmhqHpN
f36iGem8Tqo+8JHkdBrSnic0Lw/yh8WCGns6kRX0+XS+qvYPutHU9ZBmjxwJ4K6d
e7a4IGxAtuzCVuhQcEcPDTRXkLHv85jl6n0JR/6bdvvV667KjrhOzRDO7kjyfUMZ
zubPCJyKoTOLq3vVD+XsNUXlLirX7Elc4No8u/F4kHB02KJ5eyHF7GQV/sehwvsl
Zsz6ITUwjbwpZlW8uR2ETaBH++T3IWVE8vjR6ovOcp38cZJNBuk3DkM2AhDGqlyB
vXB7sfb4HvkfEtSYo9gk6J5KaCLKuMyKi+DdfAiqSPMrdB8Z+argamsVaxMd+Gnq
z+rwxhbVGYxsWGHDuBukH1ObKXuQ0brZq5MFybCJXnPiDYSCAuTsOVFDVQkNOqbA
fhdkljjH+A6Yu8GboYT8QVkbX73XF5I/fdwgsRgJZ+mi+aMmFcaN0cZulKJqeVdX
mYyBDRaDYIBHPJO89aI0F2kfGgNnkLDLCMQPRbUFUnANVgEvOuPc9YXCFjTHpRlI
lx/lwpS6y7CMzLIqehhyeK5gfFO7jes4URhCoDTP0e5Kg3SKgbRFy3gLQUKy3jZu
GfnrWNWRdg+4jeyncxUyua30HosvDZhRUPoX0Zl7q3gNEx9Opcq0bG8RgkIf3mjM
KlTA59WD65uRTnRgcadUjsLaTS9Bqs+plLJuMaD5nVnGEcOKhQBS1toaZx7ZqzqS
AjXtNSdHHjIE+gG4ZSrillxJdMXvSMVkhOcihlR6XBABPcHm7B4TpMpB3sv6G1R5
PFFNUHp/OhLpA9Zl7vZWZ/Qi5UgGoOR8OJGg0tzYg1tBqQlKDrOvRIMkLtx1cgqX
lkiDHKxGNwjmGBLs0ZiRmAPpsYPZgPLLejpB6+lhBn7o/Z+4K1hXcYJ3hI518i26
UOrnFFVnOzGmy1yxJP0WELFJ4UxFRELS9EOJy1fVnlV13/V23GWKCs4bEzuaKqYz
6M4lDFPba+wAB7UFGI28Q1pEbfmCU++fku4w2MMIZBYeNDSB93I5hD1LF4B3Sl6t
Q7JmFkLqbrdfa0vE7D+kVNf5pMghXwRnd/veEt+KyPhL0cBTOMERIwIayt5nbm0a
RUtfwlOnYxSl29wymJ0xix41GxlTf4rD+QjOPpcLvxUu7dXm9/Skxu0E3iZ7shm7
+YmLmHR228zzzofdAcQNBBv/TUlxbcTxvj7wMSXpfrSRU8ENY1TdKFD/tIvlgz0u
LnGiOgshoXGe/JTuKDDsA3VagUOOQGcaIVbYyWiDLBz8Q0IALPwd5jqmJoYA7xI+
pO4PHCAOAQFEsFv1UlQ0Oa7UFadQOQoome+CFW0UwI6JB5Kr/8+K30vOkMiVK+fm
2FRmWQpSUaV7uh/jftA8iuIl5VuQh8Lu3SRb6VshhxHZ4ezfViYh/DgdVszs6ihy
SMbz0Nyzo4RjmEGo/PYoJxV2y3N3NVaiVwXCszi2eujMhkJ8VDplE8u3+IxiDRY/
qx6gO/9wdRoLQBzMv5IiNqvKu+zv0jWOHSVi+JkQCvgPqMZL6wqnZ/3HB2+WDDXB
Zn5XtRjX6ucaop/kXcbRQ9k8xwqeDJ7eVkHgkRkaC22J144iu5n4QCB5UuvGDK7t
BY7QKwf/RlRMzpnU8f26yGhfPDnhP1ziDksL0VFJMhKcwnlPl2zYlvgxyxeVQ5of
Z1OHFVHDQ+9zv7XlNrw4UZsUDsGWseCmgi4jiAbykExiZuDEavd3VH+sXaPWJXe3
hh4f10TB48awhkULD+/NbyU+7NyUSpyQPV0xUUVb0FV0D8gF8SU5UJEEjoAu83Yo
MxrTXiwF6QtgjAPVpOZxmjObLzfDvB10+LUH52n+sjxMY3k2cNJVkSRSjtbmiuCL
LoJgBXuxi3okJJZkXF1IaPD8Zr004ze05Go8ImJF5N83LV7SlHsR3Gv3VaeX1q6/
8LpS77ftlQGTE0nprswPeRZg+Z36Cj9Ruga6uiBEBsyIsISOMWCoSeyvwBFXs68l
DsqQScswh1z2Ir9TIOBkaFP838H4ADaD6rn9pGLjhdjsvs0XcckMoFoBZ1zjErsp
K7nOytPSLUD6kOWuOxrzAHqs/BzUwZ//DQoBnyyOjZDWzGvUSZW/MbR7KDSWYlsz
75rWMpMkqTz4iLeInXUwh04irzV5UA/T1ZQFBWK48Qie1hZGw03K2btBwbz7B4xb
Ya0g6lvdPeXv9BPfBE5n2QlGlLh0H7pGaQTJceLl540UE2It1MUjvDULyfEP4e75
8mbNNI/4FYRoWB/ffKyBslbySerw1mn55e/joyNJ/J6mibIyspWIp21wvDjZO3Tq
mqNzVvY0i5q//snD2lMJytuvY+I0sUva6tmWAfsi5tclSP9poHi+TjGuqjV6J80Z
IEgpP/dmIGqnYRPDv6bGMvzDA3kzp0pyJM2maU16cSTfTRWW0uR3mRB+3HoX/1Z6
/KTaVKK+XS/h+5/oXfS4FJ/gWAQ8LCWL4OcYG+MvML7s7uqgIBDTf5X0Okskj2c6
DYzHqHPxMZlAmBN6Cr2KbHZolYCIQBjj5pqquaCgkLWmCuMtpAUXlw3FXKFwvR/W
Pipnztep4QJFn894hlpSCQHqV0ApnKICmBNWACwTCTcJqJfNE3tf7sa9he/ZIEGy
WbRpjUG56ZCErQCJXpHUUGBtEhGZT8MZoA44oOceFS9/MLlw/ihFMyY2oDM66P6o
hPq3ejul2Himix88dVqC/xlxm46pOEPvKUpFNqwy2un+U9Sqkxz22VCpa2CEZ0B7
CzFdf40RQLSEq9yghPmRVIPwUtJHPTPVzvWKhdFGWPdK98FGgmi19kJ270lKEe4w
1R1wu4kNxXkyy2JB+0oC2qyKAKLMrq90jvCNLODbFxqEw8Fm8Fla5YTCvHMhwZ7A
C+qeJYFEbC6hB8jgtJSSYe2XP/emh74lSK3KLypSTCK2PXzHHkkqwJ/oJYr20hpB
G/BAvdT4dgB8wnujR/uzm8luKKC3bs+lJc7oK8qFdvF0PuuScWZ4HyxJIZjJ4/71
6pZ2o3dCup3obaQSp0b2GhfawFfwkx5V+T6JY5opYNATbEfzc6PdGjpJ0Bfbxi7v
LPjZEU++5t74la6T0kZSB+HT6PlEUWXvFP/49DGQexUoSoGx7oLVmC49pLgMwObk
jJDewqblqzT5Za2cnXLNa5/DT5vKO5aY6Ol61maX46AlEmL3g4u8CgrSzxtOWupS
DHkHybgvxrsiNfgInfxTB1L5+49vNG0X5EgtX95MRrciNg26cNmUMHyZsaHcN/T6
p71gAL/U7EZ/BswxS/ydA/EnwDIEtDSPlDx2KhmuhgLB6w7mrb2xUkDnfxEy2z0n
eRbOC4dnOZGlWZwSkk1RqH0aNByMxnCmfXqnwzIRQ9wDKiNyzzBN/juqMlkrN+DA
pS5BF/VjjPbtsHOBBdCvr7c3JZNVpeqr1deO8U9K1qnsfVRAS9K3KJqDtw3h9R/z
bDieGFg9ueKPXwZcNtIF0fhjRlM4cyUsLigba5Ts6FMgZTGpOe+HMhb14qhZHUyf
DlkPoztPXjQj03aDUQL0AZAFOJxswGpSIU+6lJWij+63GfiR+a8u/jqnqrhZcI8B
SW6rL73rHo7TeLLA+6pi5WitgGBG6bCjTCYmgHUZxpZSRo87BOyeHy4jAbW6Pqxb
ONs50dtl8FnQNxlmg5HHpgIOeWziVq00aNYWQ/lx2BjhO42K/Fu4Len1ZQ+p8oHz
Tf7Nxz7HcZsEh7DsOMTvwOZ/fMReWGRS2ksgFLlukCtpgC6IxdcH1pHXw13B4fJd
mPgAvS4wWxKQYH9pWuAfFwhI67H4XdkH9Cs1At6hQZtijS0x9ptH/eaHfmuLgd5+
fvXd9ezbBEK0nTY+Wb8zIGWh3NrA+6sSkPdlgRqBvXLVfCR0ECF3M1Qq8Cm3lF85
JivLzYTTVlwqVzTj/QBOsZKNp20LQh9Jx+6Zx7eHCJAYAtqF5fmmRKYHT46nYp8E
RMFZQV8KmgThZQ9PomY7PrPb5V8GcUQAZLAitYLM2TROulQ/LrnUfsosv60a8pOO
bunP8lhby0jOvQzY4SrIoIXHSuqQiH8v/6v8uTiejtNeluJaiikeTv7r4zt9514D
NK8iLJJt6/SLHoPHfRC5jHxswOVg/ldeMU7jlAtgJwT6WKfwhrCqE+1q1pBs61bO
lsiOfD9v/2UHTQnGUsn7B55r0SrrxRiI0me7Qz0Hai7RGXYS8IYybN6fVPrZAw0L
BjmFmdCPG0JMhO0CNJAP1JbY8+XmM/RaqNKc1J4YRlg3NYa1oq8LxiwxTxqvob19
6uYheK2P5653s+jyfU2ygi9XYyRMkKX0Wt9lcfpGy2t1LXAhHi+CBzP5cCQtB9fN
4YPT+IzZaxMqJfYp44cWHLxOa2Q6HRZHRX1cMS4ld2wsm8oNtnYln56Sb7SW3zOr
oIFcsJYfTpLwQCXASHbWB73W8uqWSIX1EvBkFSHE1lN1yXw8d6rt++gbdUseJNTo
7qgBOUOI9I16mZbmof51EdqCOROOMHcacywxpYiFWnomD7G1hrmHzf07BpyYE9PK
g1x/UJLTDgwqnXROmxdvOOBKu/GpG4jR0WDwxGwRArcQCq6yIJDTcPceOhW3ZouD
rMXo1gbcVRtg8SjQGrVxZCNi+uuZimYfEB4+h8OZDtLRKffOZOyIkfTW6dqFy/wC
HddB7JnSQRgsLtySr+IittyHGrFYo+LkA7mryeanlpVPhy4rfHAtWHS5IEp33JBd
8EjSWJByU/hoelyjhXe0Wtyp7Y19TnwB9upmbFhDxpiFOTBTClEi6Fq5+rrcRAqB
yF31+fEgCShnalG+JuMLpdbCx3pTs8aHXhGxnY3ri4Bi3j8IdyxWIuzJUp12b2MH
saWV3E7RuB3juRkdmI9KTMzLqKWmWboGqaij7Muk111LqnXS4hzmJ5hDl1S28y2c
BLfpmCM/lwmAGAYPV1KFHf+QBDFWtLFGfGynwcIXgf6HpX4W52LanUxkWkNslTJC
igqL7EtuOSq3qhcdZ7BRA1pddTdsYSF7RNlxkswQK4ocZrttfv5YxLMRqupuksou
apgiN7UhoELOKzLyl4nAOBjs/0zN5WcVOlYP8S36fESD37K6Yzjg6alVNPuEyz7v
ZsBDgdw2DdNkKrXnfv/taAjGefNB9mJZin0O/bJjkQJIybmtGTrrn1JxpBPKEpLt
xRpIfOI18d25g4GwLPXOOL+9/pBZ0ZXgy/Efh083zeQQ5ELqR84BhkDw10f2Jk4g
+AIVLpMTv4w0A/XyKvlJMRPt8dbE3TM4WsEmfppEG3cg5C6msiOaKZ5IqH9R3KZe
cjgOsI84bVV89IOG6uTiM35WggRj/D8pRo/Bep2u8FKCSY3WdZUs1RamqOZFCpWu
ZN8n1A4OD1WgkApCqSbNeXCLR5pNSTDETuQFEDwL3y4JJ4ZYr3Az5K9xP3ppBGvg
RiYq7ZzHh3VGtfD+zBPIPVMMHgxFtqqRUDcsha9zbWm0p37EhOPwRgxML0IV0U6E
0zIYPGvN3GosOQcb9+DiHwrZGvdnsTqu/2rWW+3o8+/whdlhAJiCPKd9bxdmWW0l
+nie6DdXQP9B7QOPYigH3GiuDLbxee0f0IcD03wTxSAlcNrqUy7458x7rHzNv4NV
VNwTH2iE2sh9ekPghDlqp3FIFjnyk8g2+CQ5XTwvksuaRDIz+A16ckDvMAUniINn
GakVq1/byQhfUI1kRZncolTLaaaYU+W+xOHIZuUE0xggHm0+TLSYLpQqeOOV/2Fo
8kE6jsXfyPQwIc/YLObbebwppi5p2bsEQJT2XmKAo8tMsy9ui4HsFkLKS20ZwI6g
UKJQ84g2hg/AkND95e37cV3vjoEoByp85cz45CCjzKK6yDTZd9BdGm5abtOzq0LA
HyJCTiC8dHFwLmQiHiuL3V83lTso7RCaSHbexfiw6z9JXF5Hsf7SJhoYfWhBv+Mw
uQS3yqEuuSUbiv5iK92YPhIdyfDXSGJGzSYsDWC4SxLA/FE8SMJNxO4mfp5OOblX
+Cqyev5nx9oexi2a4WGDaHjUILqY/eF21bndmFrhYBE0VyyasgCms8qOMGgrMezx
mXPxj4EK1eVnzHNHkBKJTBtxwl2FJYfKYXljZaho1L2/c7WjHZ4ITij9aUhorfqX
4H0bLB2RVzP7hUDgYe6HOBwDP4KqzQoR/5onedyOjrkQYlQJWkpj+LHVhdIA5ydm
dhf/mZ4DVtGoXwKWzIfu3WpqBkH7CmWORI785xT0JEgf9mSb9kV634Ft2aCtVFor
82rWdc1Z+YzWcL79rYjuia9MefWW156L2oAX1XQQPDTR4audZnCcp3mEH8fQ5rkK
hlLhXGmf4BGWqSWMZoUIYSLweNbQn206Zsx8xx443iUZmU2Uu5Y+0W/ega3hQTXK
HBp/TYGWQReW72Z+pdr9AICl6T9qjXJGli92lsLWV9OZklntao7jUAdDniO4iWq9
3lgnyJfXwAiwQW9HUJRRo6Bo3+vYTE2KPKaXvFck7HnCBJsMFLOARJYwUX7WFqOx
s8vG6I8TKF3gJvcKcj421cjOeHpl5afYluIV8eL1nigcFgCoAlx+3ZytdffaiyiI
BYoyKO1E+DemTtryTuSDdFuSAFJAimE7r0QOuGxBYW5jgTwRcUB3yHF/76j4Ky/B
fkXE0XTQxu3guB/rkide9a6foeAi5ifm464iSM2MubykxfXlq6+FEuI/C0Tvu2mv
/k4Jl8gluHdlb/FfJ+14kWavzLr0YrNlYKshUytNtgBKuMWk/Aluyn14pTdIzJKl
9yr+4cXDZ+WT022aih9zWOtUEP2YXoUuNOjkP+PXSWLlNNu4cGBQ/rkDgzHWg7Dg
Y5GRi9Nwbk6qqB77Kd3/hNOpYWIUp5zWwrDZBahtQ8ShKr8MMX/Zb5e5t7sFBlEM
p8/tw0SXOmoNqAunfwPRYmOQkGYMxm6TGj/gfZwIn6ZC3ybJz67XFIYjAL1qjYD6
A0GCoSakruOTEceh1wOLrxqgFzQQJhCPXF9TfCMCkbxxWA0NseCl9TcQbveqHvcz
v4JRLjVmpDtYM3re+y2uUXN3T+xZ7CCDHgTgI0NA0r7cmJRIm3sllXzC6IMvMfO+
0/hw0dtsE+cYen577froL52BjoFU9gbWU5Rqzl6Jovnnh4A4ur8kcGkgMoCGvjJs
pPmWsusDJ6kxrkTn2qrai5jTls4G0cJH4859xKoMGgB9QUbcX1VDiRgjdWrGxLj/
F1RYOmbx+PmgQB+5rfA4fMq02OHQyxM3at+bdkNhld//68Vv8AMAMfpq0UqYY7lJ
acTNdRX4LYcBr3cyfz2kBIffwnh81qYmh7bH8uJ3qRsDrKXWvqG5fAbtahmmUVdB
N0OcDvhDjzMkle/1dg2F/bZ/dtQMM3uOxDdsK/fsvxWPv7q4KmsRziJF+E25EuxK
+O/b0cFddbM9VAqelvG0mE4U2yq3inapnQnvwdAjrpfLJKWBbdr55K7KEVL8mW/g
7kCUiadYaW52Q8d9COBzW+9UzmKvNdrwm7r9qWOnsRTsJUGThR+TunVQs4xPAnn2
TNzbzopLGn9eiF2NHxCcTQ6OHlq4zd0gF4LqVBxLIM+XV3cpxyUYIiHMTC+Jd38v
bCwuePbujHwLtHh6683iGgB8OCbvb+DMGc/hqaUaHyqc+AqQdcXsL2jrMJ01nrbK
UZHYR4ZBWCwAFpsOUc01L8c74G2B5ujISQH/vdtusOlsUyI3E3bXPe3xg3pq6Ra0
RsP48drgkZdfjKVo6UVwPvAD7W977FyAt2GSzUp6GQu/PDOhJpDiu9gJvujl5N6k
lRGDloexaDHK/dlZ8np3IJFfLk1dNZqsAqrxsYmyO8kKdqiPYwPC72Iz9b/Cs3hU
ehmEExFLFvr5u+RYqb54XXI6WzoDVg9Uem8hry5jSFXCWwE2X/8WS5/BbKSzfE1l
Ax4fEqegJY+6byfmwVIqhyAA/qNYPnaX8enX4Hyr6bocXMmu8yQ12eOFOWFxE7Zf
DDFyItGo4o0yI4bEHqQF6UJ6OAtxT59R/TNAntJpRVWySEY/SHguGNLRE35JKYX6
CBZ67GXg+Mdzw67tzbRWPQshgHu8OPXs2V8wsaAoy5Pngba/EOpWu2UAYWGd6A49
DooytRxXmW0y3NFPJwZ5lTEKRSQ/5/dvCsj+6Ht4aNwlKDV6bTMfzi0dJWEBpiD/
TYgRnbPC+DdjqITQ7ShQtweA8Y8TLXk/fzVNaeLxHDXfpCmtuSZpq/iDqDQe7PmF
hQ3H2asQlO/SjRoDBSwSyiPVDT+elW51atLyDsMsBrOr3/2kgfH1ijE0ha8JSnHr
XJ5GJ8F4Vpg/77uG4+hS785NsrhlgU6QDmu+KbVBxpBEiKRrXinYoSRL6K2D8vi5
2vp6jFm+OBlxWForCU5+rZEKLR/AtbyIjYsH3RJeGTpYecGNrNKysI/1ylu9Abz4
6VN1pHN9CnvRbWfrHz5Lx+COwtUogHz71YrW47VqJS4zok6isM6kmQCQnivm5upp
AzzPoB2ZvCq7wMyjv8p4iXrDnuJ05uhut6xp91z8ucQZ9f+ZKCDqt+eEvkRDJbix
kJUSwHLixw1F1D9Hd2daUZOHaPH6xd2dDArqATiv9+6GB1Q4MaClskPs4gA5Xwp/
tryk+SWGHaGEDEucA/+C7l7GInjF6zLnPtb7Yk9Z96Oj+Tq/tGb8qZXldqTnOzv2
G4Uv3oMZGcCi21iad84tSTCOW0eJB5AnDrDOlbQtqHJxDffmNAlZy77nsgfFt4q7
KARE9jUvP8+AobNt8zrIJ7WSipIpEFkCinnLWAct7RBB7ysSJWSfobYEDxWQpYhJ
1ilZQMcI2UsELXHNFMNOXsmFD9/QVXXAVs9EMRImjuWj4qupGtJYiIYE8g1LH18b
pM+/7fjCfVQ8K6vBHKWqVAQ3SNsGkT85H3skKyOTbz58eqQMEbqTDg0v9ZFu8hVE
izCMcAn2Q8Ht8rCbt+Um9x1ElghjKKbBzKbdEB8evYLLRRJOSin3IALgD6fvKM5d
aJfw8Efp1L5ceACdEAbamzh+dTojnBD+mWxuQrR9p+YaOQCWtTOIcgeFDtNY/dpt
f6YC2Z02jGBKrlh1QR8TUsjfTkOnM85GOT/9AZQfphSiInERJJ0u9nng5Ls1+aHB
bHazO7jA9qEHXNHG+lBODOS5xXX9AYjwanuCI2OKNwZREYf9qfVrNM0l7F84n0t2
OKKA8N3KN0hzSAYCPMEHTtMwjptXJKRKqBf0EEYPX7wATac5VUfmBRav1UFNhA5b
hoaoQQ3mEtMwHDl5N4nET2u6Jtzd0rh3NMl/gdEirQVfoLsaG0plm88b/ioHzbkP
SXhI0oeH6PGHQDtNtNAe3v3BAV5BIsdwI5t60UyjiaQdyi6KaQNZXsl28Xp/EiRT
tJW9TC8dsgYEb1kxE+XYWTYSc+nVG5J4B3k+dddzNLFIZj9IY5tmGot5EzFmW9Lm
sUycb+hQwQMGSya4dkaetVB4O1nNHBM9aXHKsCalKwWAe7MJKu7Y6r4FKdb9cWzI
kD4kJuXUxObZT6nI3uTTF4uPxOQ/7bAucrAxVCEEVL5vbXCecABuEUtm5etQRdI+
3IYvCP3W9p/Qt8aCjhuCaoncE9UhiVxrNHszPBi5F5MaVv0MANAS11vVL/awYCX2
PJkkGd9vEtbx3qHTctW5aHvVd4BrvyNfg3xPiZyTk1gJJVUz4b/ML3OMnm0IWElp
Huhoz93DSvwFw7Phx7CzFBQiKcfks64PIi3DZTrhDRh46Iv4GiyJWoWFmGwXvzAJ
Ql8Yv6gzzv3e5uFM6xWeE2LyiUbWrD6VE7O4Z1LRyQnU/DFnVrZ7QGJoHe+Mj3BP
aaCyI1XwuKKd7HJxPhg6gOdFy69zpw+RWbFbksQwVX0bQRPIb+vkMCTATDbJqvLU
a0r5CKo6MaoO4oitwJobEkYDGaoe1WEFXElS0WeaGDwOgkWlnb+andgvEwfqnaXl
gUCSGa7qzDBazZEnWI2BU27bmXgIpNYyziD3oXxSWgDgi9rKGTb2U2i+oDPxi+s7
uk8ujWO20WLc/OWi0ec5vLSEpHejSzk/YyTfgl7LeXuMgkUfankAWIWmAS3FjEFf
h2rgiWjSmOeYj29RJ8iypjd5aqrN8kOsOgZ9P0/Rh3+3CqH2BeUZ88gET83fNYJQ
V1jTv7aPiTpL8iTDdGCZAiaJ+yR2B+4aVu4eYHWfA3jYImj9s5YJc5H+8VFsmnE1
aA1eHEaNyh9wypoFCjUp5q0VgSfC8G5HbnZTufaTMjsn76vQwC9fZFxe1kCgSmJf
YyhJnoeBZG7YTDOP0ANVwg8X6P6eMK+cdOLOV7SQCS4z6tzdWxeOkVYPR2cULiaC
nXnse94VqJZi+HPjfpz9oVuanB209/dMOSfvHcLi0gE4EnbUB7oBO6qTp6fSyzgv
Bsw+5k/hZncm6puun93cIoDPLlc6vSEJhqoUZSZubtL/5aZFwSZLcezKbJWSkL3b
q7DtSESYMc9hfNtUeNr4eqUotieoFsinhL/6jSpkPWZRZTbHGyYCpB+/I3biNONk
LFW+ScguwyAJVhupAk/w4gsRquuc46qdeKxxYjazLPok7ZY8dytqGYK1/UXH7GwK
KWEcvtPdpm1EBXcWIH00ENh29uZ8fZdJsSa01mMEGTFsEn7pfw671mDJKh0pgwHM
6kfweirWisq+AeDHWqSmTCOEk6TgXYlcLz2GmL/cWRaBQliCqi4uMkiD/WUMSpDm
1Hk7Kbs75XDS+V5ZCPJSL2dtE5DU4yw7JP9HPWmq+hhI2CVfB5LE0E6upLtS9YT0
9MtGz3a5V6E/t+pENdr9DbMkyx54cSsGCfnANEdGlYDpOJA2QUOSfpmwPdutlrpQ
LvRTgdWegftIvRZYlWO8j2cUlzjkqtLfHh9PyxBV20HOEBathEjqxFzbrbWqrTys
tuAaP98vbgZc3aM9CbG8W8H+IvWMkDXTU1rCsGz/XlMFQLyeLqZJSTzcjk2kXsaP
QeT0bJrvsvrpWbCE7XEkrSUCUCA8hs5oGdXeOdh6Sf67ydVT4jt+Jm7TXu4GmuGa
m8v9XF3AX2jT/vIECtYPTVuLjijsYsstMAGADpj/ll145w0GsumSKAPMHocZiDja
+Ccx3mhQS3KK0E8J398yrbj5tpRooDzEUMUlOAFmjQy5pb3ggvAdyq+CNTGyOYmY
ekrmSoVBveyi3uUBpRBQQ2MlZ6MgvDZjMbswnttUbWhReAjpVjbRFyJwIpF+CjP7
UHGyAqUAhE7MS9l+2e4s+WOhoA7Q1/fLzqF+m7DD1ZepTD8R2bn6LPyx4GkFlQyG
4Ozq5IulXbaODtyEerUQl7BlaZtHT1QbuuyxK9S9xFnCsnlMeMyfyS1kb5+FZIcy
JsiqdppjEYAF+UnstTgkb0GF+5RiA92iJoAY5HcMGITraxjAyzwVpMmWXnScLCe9
m02QZyc8lnBEzHk3KZQGQoM0ORf519269pbOntkVJovEgHUO/WkDnRtAJALx29rc
0YD/Au7hIJkqdfhWPcFbHgLoy6SOrA0JvESSwa3EEUN4IjJehOJiL4A4w78W0TDG
TGqJcT29eJLlqN6bspLADY3higv9l1I0hNr2EqUOGpKwRlqb9OsoT90eoBAznujD
kqjRxYaTAkk4prC9qbfFyEch8DvH4v0LYa4FXIptlMVFaBQXH1QR3PuaF6JnWyRe
nIXR8jbufAL/NvQVUeeN8UfTd1VSgP0VxBAHN38zEE9U9eWnNZ+88rNiYxJk2pnP
vm9tWr1PiqPwe5d/cFPfJKgsLjvySWlzUR6C21bozdvlOmGl3Yd6Xnkpb3XAK8Ql
lYSpzMRLw0mR441My0ynppnAIHUl8U5SeQ9DiqsY0aPXw1gA12YEftP1XmbNEWz6
8fLvjQri9wINIYhni7NQ0My+O2mpqY/QSkM3OwcGLKJqx3XJzOOv6wAcjVZrzPj7
Ai1WwR/xUQGjCc+lHpBtkiPp7y1EYW1yd9G8MqInGIq2W+85bek+0YHf4l3tcinq
YvdtFmvgy+2Wkiwqa4buk60qcWJ6BpoD0w8Q0f6wz4bBIP0i/GZXWmZPFr1EeNUU
7lQBacwy0DpEOb9hYpXM0++Fr8b6ke8zdADQzTx66iheMBSwUBvRj3792TR+TS9y
3Oe8LkDfcThmamJ4a6N7K6wQPO0O8MH4SOpMqvV/ab+DADb4cCHm2AMo0andHX8L
LOTlq3j5vf/1Zx+VXWllt6d6GSgTE85oPeKob7oQnDv98EuE651LBRV//9vuqTaI
Xqb1HQxgKAXGnvAURBDKDI30KwJUugHYX1EmZiahz1Y0Xm3YM43zaO5aJr6JU1pa
vfgHOnuBHT88w9SpL9KU1705HADw7k3yCMAYRAGrIZZdEP+6xuClKfo8VNYRrw4p
SBx2eWfu9BDr1wJztOLVsHxWTNCQQJyhfFwUVz/hZdiY6427eHe8U+qXd241P1gV
D5PzQtZ1aGSQlP49lBvpiE8qWXPB4nf00X14Ejxcc50jV6JGu/M7bfZcRQptCKAq
cR6QExoBmUe7qc5KlAUYA8xn3wXdfBT6/PSzFb2dVfx0SupSNMSf7crblZUJWQVC
U0R+3o95vhtOl8tqpAqwkTX5Ugaw/9iTElAUazlFSru5MLWnSf+OnLPA1BNihn42
qEUmGLLZEyC7k7Z+y36+61SBz0SnIJNz55DLPD6tcsBTopC7SMrCBhsyGqc31w6c
A/7aIxEnSXiZJeLYOzfGH94G8gayT8fyF8GINz85G6rc00ONcqkcTiJUoaEC6m+2
3oSlyT7i/1e2F6Cj3+/HpFJF1XEyCovNlIwvE0L2sDRSFpID2W+2ugr1VUvOxH4E
TJ4saxvHo3xVASy3HW05HHJMrWO/xbbiZTYNb/qDW9OLOjUmHb/74MRZ7x/YKsVp
MTpLXmFIYis4wvntQ017/5aY0HHo8XLyNsEbLizHo5ZU5/ue5A4EOQn8h0CGa/Ci
5N0k2dPgSpeqo+cB/hhB3ovVeYVisXOqfkG7T1oEJn7yqtGBUt03bSknOrdDdzb2
ZiAsPzDlIIhnuY58tprZg9q1xhFrmadN6yxO1L+EhvUNVfrtn/WVbyTKP2rFmIUA
U4eTwj/Sj5wXzcsJUTm8BK5R1RlSZPSwMY+j6QgBz5zssAUZRsPc7BXQJGSJ2uGw
GgkjP2RJC6vjMpAc3PX/gu4NLevFt7B04HnTpAdvHMZUtE4LQ3FWKX9n3rS/9gYI
QloVj7a8cInKmeyoLayg28MLq9Seho/0WSdiRwLmPPPx+EFQIgQEDMNIjRngkDSD
MBQb0/DK6xrr4+4g0bq88uaTGuBC3nxsRHBrR2SXpZsp9Ibl4KD4FEuVIe52GaqH
hkwsPEDV8606UfTTZYBKbRPJJS50OxlOcak2SPOYEWZM9gTGIp96fSXNTPVoENqS
H0ejHvuld2NU7tqCxkMxK3kv7CvftPowX7HdjibK0bEHz/rS+jSscKaBeUeVhvHS
ftpT/804ugYsBOlbJpHtAzMr+gLkoWdxdRqFVwckzUqtcz30xJJhKK0MVMCsChtG
LKgF1rSDTOWnlbmVOSO8/q10tZ50S09W1a6LGjVt+IzdZyO4JTOzc/qdlx6dsbJp
wAmZbWxAVRHXjZ+ONLYzoT1c9eYo8Cy58whsVfaz5uwejj7A967JiEti/fucRL/U
ilbYiZtvjRnbsj3mJqoinHjUFqI8Od/zdsZuR4+oNaDVLLPPqLla11kiQN0a8lRc
CPXRSVc5aIPBTOkeV5gjtEbALQwcb01MUuj3vqjFBF1kZQSa6/yAI1wxdkNNeCzF
QeWWag799hBQhmnUO/y7W4YxnHTIOoOXqUpAufUvfpJNICNouJVPBRwU6bf/twTF
kpEYSV0v5lrsVUeCrYAwrPG2koibOsQ1Eec/2UBVgA9qF/MXv+s9fhuvj8Dl6jsH
yQi0CgS4rg9eZzm9XvEcbi0TYA0tSDA5ozuOKnhywsLDAzYvMvZdncFcyD7dyRNJ
T+OHX3rHM3A1ZIC9CWmY3UMc7mAGXeCA5EiW/Mg1hsW/tXAbj45GzMDkUExGdUTJ
H6RD5QGNb37ZYksPwxbI/2xoZXeMb93uCFr4dkh/43FhihSFmqJli6mTOFniwMrq
5aR1ZD8+w6jcozbHfTcueBO6TlWYRwrG8AffblD5YhfMmn+SaFKk+97bPK+6qjIT
EvYdT0nYPX3u7Qdy9LxScW1XjjkgQvlY2XF/HTiiK3nhva56jzLw4/0Vi1krO9C/
7UpoF1MQXES7zfTXvtI8iIHh2mYX6EZOvwJXo6jo0FSUOfl8ZIiYJ6tUE8LcoQDn
W2f8VgeXIfQLTQ/KheQXm1KD5v7y3sOLOL3v43gTMjIFnDOBAFa9TBYXxeEnb7mg
jhKz1fb3gLabbvpK8YuMduuaxHrDYiLNEtvH94Wm//xc7QOmaJQAl2JR18G44j20
1N89SRfegERXvMJKPlVZ4XAAi4QMcsX+k5UAINwxbigpm2O8m19edbMSZVCNDeF1
2MIb4yU1rXizBoDzIvY67FyaSDQSovZF6NqqTtHHl+sJ3ooX2eWWJPcp5ptSRgo0
q/wQlqUs2kRN7M32CB8cU7jNPc+PvkTJxqBUa4NvX4w387+u9FEhPPVa+orITekZ
6BVArBg8u8k6A5WH4xHi/aTdMpIx/F1rxEw/VQNM778HjVoa8tzyC55UaZfeTnfN
rA5ohuuHv38eH1HrRIecSdnJ3wZWYaHzetbSntPBkge2Xjc3oocQZifgl/78x6DC
yLvauqnVm8zymViUodlQcdNw2PGDpm9bk5p52Kq1jdgc3m/B5XQRQv5KLEXrlhCr
6cT8W2sdkD1Re1w4wfB9TyVKHZQ8saSig7PzTn4AyM5TRMTdRMnZvWU1oMrY/94M
SO88YDh4ysiFdeg+Ov17GD5ofwRpr2zVU1GtBcbaFAdhcmExHvlA5E/ovDAu4Ony
D0KSOWpJK2urnHalJCnAjTNaBbNm+8lCPOn72jWT2TGvpq6h8pXy5WUEwTqgjVFP
w1lm9m7htzIBxxC9NLutdMYaTWlkgWkYSYQClMHKPfRHADP5bD1gycsp04fxRHPX
rvQALv+j+Jq9oeR6B7j0FzG9E//hIa/dsPHTEydMJXkTGcmRtU717xi9Fcl7sF+r
3YI7G8hOSzntlqcoXpVrM+ZUdOC1HLqLNHuEHFyUVtFsFx0eQ4WkpkQshFz6hMOP
MYfUECaoqAsShkSf9ENpCrwH/i3xE6efwChf92DLwcTM+OUqqMfBXOKphZofvBPK
J6IA7hbGUqOv5G6hiEiWK7WjJ7lQPVdMEIh/yXCfb5ZbaNn3hPI1FVdnpj9W7ihH
2rjzAaHdHF76p/4pRK37hC7/xFfZz7APYHcy1LmwHII/NOC6TQj8sDCoCWdSxcIR
cQZO4eP5kH1TysroWHeCZk4ncubOyrzEKwFgC7c5hrK/LHuSVmxfLVDQizxuajiD
0CeRbGUXhpoWtpgT8qkkp+doD7CNiWOa+vY42VhuRqbSldlz5srJglQ3CK8WVxu2
B1yKe+m7r1PLJ4w4cBZ7ZofnURl6Pnm/dbrBuueOq8YxOy7/hCoTfs5hWoc7MG++
N3EfjDDzar1qVzDdLRrDcuhqwqQSbL9bFmSFrs6T+8VDr1x4YUN5gO6pu4Lko+ry
cvXCsF0ToqryHFslWM4u4nZijeyfdpYzrrPCaYwkogxlAzhNljevzMQuX7Gyjo0w
oGfwAsGqq3dndwqTDFVExtr0D+k1+etDPCy32koNtwitsw1ZwQlRY2cD7DRriMyt
xy8KjaDEOLIo+iSCkkoNxoOPhgArAxd/rf9tlLhqDKeIAqDxd8MlT9ddB/ozKuiJ
T+z4S4hFfofDCD67ptWlkxwecvfLBT9r7ukWvR1pbDb1EokUnpnkBCkcv0l7foq0
mNOEwTfe2EasyvI7A0I3hydhcMRRx+hCc/6wLHVznP+EAJf+uyDf3qWgefjvUMoJ
RhcjlARsu7KiT4m/FryPHtRVei1vprIGIHD8MkXC03BD4/Yn5sb8jbPxfodSvC6H
j2l8y7us/V6y9fH0RM+IR8IFnvVhjluFzdRaf86Jh00jXdb6FeJhdJTVGpPiw8QL
RdLRGQIhGsITsvTHLezB8os7qTQCrZtPa8KZcVZuWFoOdo0iU4W7oqBqh/SyWpC8
EEVLUi1qprfuT/3PUj1WO9aROcd8mGuH9fUDGOdWekF/UJySWedWepcEFtFUj0GM
AwDtZX3ofcuoFWlUOHta6ws5cnNxrk3Llz4JzqpsJq/0AbC5b8snRClk5yJr+z1s
xK5VJtepwUcl8+XI4z1Ox2b+oQ7gXej9+arySQwxMucgtNJs6lkvWD6Pbzs9hdJk
LSlzaJugICRUQyN5inZ5ooKjdhzvo4SwIGNwdQze2wGHtRGcdjOExPK64y5H63rI
UVeqXXuYoKDVP818Qqk01jJWf6yHYVs5+VloDOihoJXflht2sMLRTOlP1TKtq350
0zxySs0JzFP6b59CbjuDSE6JZn8aCxluWjwx2/0FGSAhfPl331LTSL1Bb0XRMLNL
RI/teasZ8xulG4IrPDrbBy6DCT8K6wQ6Q5yeA+WB2XaPrVQtDGfTiuBB9BJT/o69
iYkNeSttG7UMgYZfheoH+s3xcW3ETiegUatb4wkwmulq7l5NbxtfeClZ6QkHVUxA
r4YuJwLbS/EUepnB6bEpBQmEwj+T3v/EYkZDcLhWn2qCuJd66TuaGwRx0gFNWPXY
xuqlwJcDvN0RnpXOA4PJ9sMZwhj+CYAMeO5YPLVJFl6o3MEkHbkJgG0IRvfn1LgF
r6Q74zDkgs3M3yElo/iVgBYEj3vE8a20hvhLU8VUWtl8D6VQYhnOQ8cglqAjpgP3
JRBLc+PIGY17cF1wu2+bSTRosGKQ/A+cgyTmp+AfyoMPOhmmwngkGv/e6lIwpD+G
5LLUcTNVSCZTUPz5oNF/W8Hz+3uRE/fz2c4NvGbW8f+AVAXpyCBxNTQMtTOzm4EF
MdlJVB9d17XYTW+Q8/xAL39afe8XVY/EXcPFKhbGsn8X+cWU0drm1DQ1CDATX5lV
SpAfWZPYOoOec3mqRIHHwWiY6/5VYblFD5lj41kIatwPekXWglKrZmme72HUhrZQ
w+HgoBOPZJj+5ev7l2EH2oMVo98n5tHAbEuF3iYvpYd2qJ7ukvFXhTq8vqvhcHXH
RROVrRhbWYvbRc2hNZLzCEFLvE4T8eXudiUIkdrSGZ2gZwJLHpJiD46HT1LT1/AF
2HjQ4kgkoXlKySfYURAycooopcKXu+My+2gr5umAs4s4TZvmmzSWL419N6fRh5h+
O7WtkP1Bb4mwsqH6vvzRlec/dzyd5m0EvuePm2qqhP3uk06M6hWHn/UWLetRdf1K
0dD0LPY4ArJLpx3I4L5AKs2yVH8Vag4gsdEJxgzk0Y8ynNVMkBMcW2pQ6dUEq5EG
CBC3lsFuv4dI4aPQvasqh29ILZH8shIfvy8UKPXHuTV4MXDooeQqM3Y5y9Dv20F9
oasf5hMO/VpbN4aKeOoMOwDzBg/jATKtuXJYdtx+qfN889ElgNpO14+MWeQ3/ruy
f54HlNpD32u83TsJ5kFD0VpuOdnvEjv2k2mdlhjeUSVKN5RYlWqiQS8XVezZZ7Y1
c3RqnkOmKcQymwFhD+5WdodiMCFU7ZwjVcejbBM3F6IlzVhz4SnKgbA0H3Sz/vVL
NUayB/tosx+1GUzMk/2/nxMviVYrttpgL9SFyxwYyzhaGTmShIfRqffYcioewhx1
qpXDJs/kmcOw1xsrFPTTsVMMA5MZwJtV525WqPHFXTBKLq1PHLBm4EW2brzt8pRg
Uh6E7kl7gNQBEghvqL3k/BI7XiWmNdteOtj0diTf/xlHS4y5AR59tcjdx1UDz5Ad
WWqpaCObm+Kl5G0vtnQBcD3UAalRW5IKcuf1DO2rmdRZ4pRFqnUuhAPOArikSmkb
I9g1zQTpp2ubMvgcoM1FaioTh72ODm+yGFkUOVbO9oQrLrsQaLF6uD+Qq4c4fs1L
c4c7wIY1pVzZpxONRmunFf2CmzJRUwNx+qtsoqWIgu/3L77rIVRRHSMXfm06mDCW
X+E6VhMBhdZwUqZlbcvPg2T+v/B7enrs+8tfng4Jqj0YLAhuAE+4bvCTMzkJy4iK
EMVzYUA7rBTQ0IUVFSrLYPsYkgZzDc9BtEvRRMMnn16fsoszNhJZ/p8rdzfxUNWN
FrDdgNVB4MpKyOhgfSIzVpnuacVMr/brZoqe6eTM3SnBWtWKSraXd2sXup2nwj3d
KZNNKg7Ju4IJ6kfE4aGCfnEgnWZ65ZQAAWCdzuBwIEDmEpnKa5pfwcRuSxc7ny/L
OsnOxaYkiAHcl4dlFst6l3MSkdPsXCtpU7mOUITqHhDt/3Sx9BVu9bu9KVEWzFAX
2c4GTzn2CSBmLqzkM/aQPqopFwfoJ5YCqmaSwFBkkU8RuLqhrxc+ADXpw0d6UuNw
JR7wFPx20tMPGNPih7Ix+ns9zRYTJDEYm3fgHFtD4z2SD5nNarZMcv/poXTJcqaY
jhFeNa0Tbi6qBydcGbKcanoJVrgorobDd5CKvxbr3rKPo1zbBTADdzzH0WcnguHf
Giv4yW360wGlJLYeULyrCTBTfKqkxG5mzEKfg5Y/K1VohDyiAbFpSSRO4WRvhwNz
2l2NIFWQ2GibSGTxuoDXL6uB9U1sPGXyqadz4iuVpWG/Va0KpG+JyNLtTFJKMkJI
HXGPb3oTBUgdIF2MBSVdbg5YUR1wvW2mZMvyad5lRxZYAoWPCU5hkB1+eo38n8uj
solU6OAcujFHfW6Vo/+TlJq90wEoXoafdmc7I5xpHbb3fLqcsuV8+vMf4lZ6Odbm
QWzIJvnYfURxsBRKaFhni/2xwFTcPKW43uc1t/BOCEl2RuUkekkK3Empqm6+2/qg
Eg2F6Joq3ADJdPBkC3cbP68um0gcidnWqBkdWRICdkJstUKE+lp5pd8wnCgzc0Oe
KtWpDXkUPT9idEK4wyqMyqoxflv1Yyzl8UsIWNU3eZrAIH+uWWByUkIYWkINOFwY
Byg0JqcTsUf77do5hWU4xEJMoeLBLwvzd9wpGa0UklV3PU2oeBnHQzHDoBx6DUpl
DIHCvr02ICikQ6Ou0mS/e8Hzzc5zns04moV23VYMgCSHGhwd7QlIEtojLUyjIa5a
zDUboaloXwDyIilgw2wqX9K82vA6B/oYncHhAvNZas8DG8DkX0Wca5DDL+sto6cu
Uy1zR5O3foGOEe/POKphiu6TDsepvCl3ibtY7VY6cBMHfvbyqzSG/jrPBjMq6Fsu
S8ke0pNwitKs9PZ5DBktLv4YAjkNa0kCKNlztPWzhGw/ROIDFPLO3mY8qxcFCN4V
w2bfmEuNi0IHlhZ31K2KgF5VOv6MRSQMJeFqXqX0hUSNBNK0IzXBYCAx7xWByawZ
ChuOhy3xGbSsjKTMQrw2qn87o01GkS5YgYFFjC+pSoIAIN1XrgDYkOE0LnGPv+z4
w7/ayyvQPVBQ9K/n8z4GznE2mOcecsy1l8unIiQQb7hQ+5aokqvA9XbyGlMtLDg3
ujPQdntPf4yCKJAPQlc6yViBZAmlIUhGVnhidGw/7ox2oIc5aASYXFyCGWwrd6DX
Z7P4gnF6L1sC0lHC3mSxQ7sKizHtt1sBpzyrSnQe6TEm/+jAIMFoaCdOopW1BCY+
rbolBS5THJWD83kU1g1yvl6dzNoPviHc0mLvICdBflxe226MvUhAtHXpr8zc7xmw
spjWTksDxRR8vvIuRb1f7wUF3AutCBrtf8Hs79dw4uPuXh8Nktpj4WcS9lQ9ryQc
63k7YjVxwWUXZHJPinYWBz3NipWTQ6WlYcCV2IKTvxSIMVYA/POoJasyYXdlNqgt
Z/03BrWd2x7UgfOngsEi6Hal3Ht7RtOGfjv4dGb18j8dosJkW6SlDgj67FFL23Cf
vHaxfBj50fwZiBtAUcgmaDh8qgJOtTc7yFGrNJu7ahqRGPEFatqbqxTSsaqu8euI
Thdi6pXstFrLbic1cxY3wFPJw5mUyI6Q8FxArYM5p2rMr3rVMG1rN/+5x2lgVXIM
J82FFED5ZeUALtoBaOIOg6fQcdjhrtEXZwQI+ShuYPNjQS1E4B+s8id5MW0hiB4o
iWQnM1bPhfZFlAlOm3dnAQ36J9EStpxvBH5H/34SrbmjDnGa5fgu6Rud+M31kWb/
s6jc6ayM0IigZvPrfL2HR3BibwG6nxUAxzgZ6aH7xojvEleBt9YltGXj7XQEWgRA
5gLlWdZ/XDOwF55JjZH06LO5qit3T5f18yaikfk8gwBgvUzQAKjclf9r0mXCydgo
g9SSlwt0XBycRbTdaTYMWwi5JcEp9Ftzymmocqh60yFVVh2ykMRbx0KVBtUj99UG
oKEiLCeWhE2B0TrWu2MgDNEgpQ0TRFUmhz+VQ6z5UFHpAjDzoCBVF3TDfAEGioYz
pQrfVi0YPFjweekwSodMRXS0HHoSjQizstoMiKwcYEsLIeR9Sg00Dr+rJoMMkV93
TWe3oU1vBj3crRnvTEZwuukIane8MbcLhfsCA7RiUzF0RwzHqd4/QW+47mJ0D388
7/Tiouoq+azk6Xgz+uLaAKyTD4uV6kxNQzFUAPcE/xOcQ71Vk04rNXb8LhzLuguE
8CDOY3y16mLIZi6UI4AMlytVMVABt9SxMonBqdpf+jSDa2y9YZQncQY/X0hXSncO
ht59O2nyKklRCPBkAVHoTUtnjsq+5LJ0u/gAGLbxvcBMSRj+8gPX/pBLabM9Twj2
1RAM5KTJo6h5+CpW5BfRRun+Fk3Qz8kUEH45jBPtJNp3gh4vnL9A7K0QVCboqCFD
HVJtdfilBdGww8QQU/UsbeNN2i6TrWxfUdgt7bRI5JaoeZmsSi5Fcsi4WMGZO8Rn
dZRLLLWZWCd+gijIFIr0WDNJ4HLIdfOWjpVOY/T+xswX0TCqdcCCx/5nps4+9vQt
49rXqE2ROoaMqkgE4HsCjY5J4noFSQnkG2Z3IAFNn3jeMeu3d0RHyfz2ESX+EqqG
w4crJUPKns89blRIyxgMxu6zrLD5WMY4wAtmOh9/lPH2ATAjGkDafK0AI4daNTj3
5zR355xOWhJrUdEx6wn+/cwbBiIojaH2dCMvMn2i5PN8OxcRSGH10pJuFAqFd+e5
kIO0LkElIrj8kyAD1BFk2XcTJYKa0ZSUngIrgr90FZcjUtAshcQGw2igygZM+AWS
LNxrd4XISGJEQgSrfQUdlUv/9s1UGXQg/zMRSx91ffF/13kk760vSD8ztvL27GNq
xW4EN2nQVm2wwFv6yxt5bXhiPIuJBsyCVDpkxnK86mRKA1VCHBM4F6mTw/7oio/w
ymjdTlD8pSPdRis875nEwczdN0DU1qMBvv1iW++22jUI69LrpAWtGlPtov2xB9P4
6AEYpwD9orRkpUJyx015gA6UFEaXaD0yaCfXsDEVWCJC60F58dlHIWS8RBWfSeWR
3OUzC0HyqFBzhc4JMrmzua/JrXe47FZSE+WKeWR+ToTBqgNoJx4nVJF3TnVAC/n1
1wLUDwc2hvlIty3yBxvhx0DL3IoGVUpkFj/yHwUY8VqR/CuqFb5YnIXHkz/Wfa8W
Lsmg36JZvR/NcwVQR018ksey0z30wNE4SkZTmxh7HC0QKRYIjo92jcMOsPs67Ggg
cqpdGHTdsHj38Mwbsj35+cw8Kor4s/AIJueP2i6tVU1nBXo9FVMDY3LYv1L2sLNF
SxglxCNdXBuoBiL4Oq8cauTNLZgpjwRF+D9c2UZzWzo8aUOQGi6J9HVbZMOhQ5xM
b7elCcmlLkzHnWBQeRyxrfCeKNVzBbBE0UxyXmXMDl4ufCa+WewiWK2KWcEaneMk
UhqeWrp8HuoUlL4sZMbvvXF2yrqg4KksWygRpA0vV3HUGAtymEzC35mR0fY4YToH
Kpial27zfoojrIwhP/KtIjpGRuO3Rg/lqNRbls/jumwg4QHWRx24aCsOx5ta9lWo
Y+/qjurqOcVz+ne06Ac27DreC4hI9dFO32JxnfBAvhWJcaudvYAOlBLwSHrY3amM
UKHh+Xg8GRBNN1IW2ndYEJ+0mOSuANEvcW8RyI4g4t5D8dDzmwaTdQYfQa0LpMyx
hmyDtsnTFQyEuamkCpThmYBsXBHjSmpIkNeeafGY7xDQdPceJd7btgoAWfIGXXis
GKkgV0uAN/kbsMn6YGRXkb2YPRifFPcg2xd4DQFUZZ+eH5rvNG73Bz+Rd/fay7P/
yhWbT857sGR/19VfgFEr0hsdGtAHwncJuYbuaxIT2eE0oDr8vPTq1HbDaME0BD2H
86XzmknHoK+6BZKfMsp20wO/oZ34Fn9BGkQ5QY78UCrDQUFdjN9SU44E15HYIdvG
ExjYKpUnMMFRiRjfoY+N4U8nWWZcRMKMlQp/wNoA7pITAJHAgrNqMXigEMKbR7FR
mV/kXCwEOw6SAtuC9SO0UwPTqn2VBbiP2ME63FXSByOuwM5pVnCN+w0EMkSmtuCB
yG0LlWWFVTAC6QUHpYl/5l+nyXR+DhqHqfOrIBUmALFpisbNJo50w+IyXQbVoyLt
xYkbXtWqQWaopKuIp0UaYXwCBOptha8FufQWjdrM3J5vEu4lJzasA1VtnFEOZCwg
+ozKINEW6wf/ZC+4AN+gklbhT0+j/ucLsP7QOwUmOJvdzrqeJicqQ+yN29xw6s4L
J/qHa0nqE/POnNXFm7gZaewpfYmYX9A+jHT97flt016oujrj1ddZUBi2BPGDNkuM
3k+n8YTHifDTuAMemiCpNpSecm8x11PpSNxCbLCXxmtU9hZMV6Xp9yA2zSdYzCEe
ccIX7sUtWSZkklcG90gfzLNBXEbaGBz6zT76t16VzY/cPA68ti575I6xGjZth/LD
A51HR8uMPjXd7yfL2MiWg90hWmRi/2y3keg3yOZjuiKGtyKs2EX6rZqpPjVEReSm
w2oJ/Zz9kp0Yat8z6eR9ugOHkeNsrH+1nDo0qUGITL+Hxhs6LVwV+i3Iz3LWdERF
yd9wiRUzevWLqT4nzd9L29Pyla+IdTItjB/Um1OwWDTaICxGrHItRdbJsLPYgRqY
TsvGOia4oT9JNzrhJ3ptaDlwfcU5gEKfqiCrApkmFJK12tHWTQbv6dcjYWe6HiDc
LZNowBv1zHJ9BEt7KlAWXD6GZvV6+7gjQEknhXqM1Fqz0KxK26fBWotSpVGfT9s/
NkEf8NJ2c8UwY4y758LECNHRf2cQ9jE0KMbp81yo3NHJFpzdCnN9i3G+Bd5HMQ5K
XRe+anM8WFJxTDBn34SAWLaq7fmnCwZWV9hDYwjVGyCrzQT5c0lTqMZEX02/eFb9
3EPlmOq9shzU5XF1vxp86H1Ysxy8C0iqOjcx6dJTra9fbNXN9M/P6B6/UYmnE+ti
pPvAkg9Nt1+DK7dDkiiF5ArGG0JxsCwKGZ7eMCwkBgl8xwJmMeeSop/1Hq6QHqWt
Rd3ingZ9n+Vr+vwMe1J8h3phEMtUV/0gWPoA1s1ecToKd2C8Rz7i/vwopY5mjnxr
jLiMxQsSOweSfj52ymTuxwD0ecxjaaqr4OsBohdDSQ/vHHvKhaJ3a4VJr0jElmqJ
Z73bnmLkbiXizWYhHB6jHXJvNZkWD9IPpm7QVoGsXeXeQEBTmSfWSt+bSA1Pybfs
uBhithcD3aUnzcvqBqldyx/kkhYo/PZDVudJvTCZborxcht1naO9KZL77WlxpUU2
1GFQKpO4rFl+EigniKQ3pkyZE2sQeLHKHIQCCfqhnZcR5kz7R7ngH6w8WX088697
6FE7cQiML88bu3sPULi47LCinAnz9/33G9I3+AvdbHBKnPmPR0WmZShjtIL4da6T
+PQ4fl+CEmhWhnpJqv0d40d4BIbRPO1chwkDrb3QcO+l1rb2SEw6ZTrN+rkeB/Dr
gtzbLUN3RJVRDD5gljwu9ejefnSehQIDu8SXkR6gaEDEBnddc07n4qHYrhRMuuIT
hMrziRCGEUmH7ICMAVv58mATFTyBeS0XxQZgdoWHweiYYb2cxbp5EyTVLu5lzfgz
+Vsi+xd4giEZIjFARxJqMDCjkyfi87ReD+4Dxbiere3KmgicxRN/r/c/dPdgFSrC
GW6387ySP686ss6k+Qmqo+b9BkEQTQPMbskW3i/ssz+86TGZRExjk4K0k+ziYLDa
nXWxR7VG+1JXVc0CtSFGgQhPd/u23weXQeEvzRrqEbI9Peq7ytxLz2yJYlOD5DI/
i+cBSvwhbn2luz9G8jbw0sWiY+TuLr//K3oLd0I6KNWaNaXaSC41gVq9dbyzj9T8
3/BHI4q+sieDEKY6mapinnUNKQcg1DplkGgiuP7lyMeVg7TovYzQuDQf3MgEKTQF
fA9F4AZpVsPB6vusaQ7FmLehsHHiAZFkTiV9nkx/iIB7ykH7ltrf5zfbYHGZ8QPN
Re0OBaFwG4m2XmZdXRcFe4SxQmtU0jfJUrmQk2zJm6LivO6vDYGGMb4usDPfHLMe
wpcN9NM0zgLE201FXXDN4e0me3m0qMDI2yZGTVENFhuRFYqkc7QSCXDYAIeITexR
uY/CdvjjNFm5gHp6I4qW3YoeaTO7rpO0KOahIptAPTR5rr302wDOoY1AocgEj5pQ
EcFT/XxRNoCGqMpvvPhcFj026gHfLvP34zs9gpbHpUVIWT3H1BS0pgGQtVNQ0r7I
3wmFxtxfNSnT+Oz8V6suiePgDVwVYDHEGl3GIqbSAUJXTvM1OilpFkrEGjkqdk4K
US041HF0Z91C4yG0EiemLh+FL+MLDPQ/UtKV39sVDxfhLuinI/JXymqt5QTCmsJK
+CrrTB+5aWJ0bPVJaPl9bALh9e1AZ0IWvs9UFKz4XAIRKt4rMAOxLPBlZALWcIkQ
9/BguDqhmgHVCWXz3IDN5C0lHzlKujKhihKUJWBnRDJYQXUcUgkRQOcHNgPOPLE9
NC/AsCWOviPSYIGai9aL6ZzZh4S8Gm6RChLnpKRBJ+FNlrPbncq/N7kiItuGNgYM
eljOevxZDtPgh+deY4wco9rY0v3BcAVzhJquTGDIBWEKKaGK6ScAGzOFjc5zB6f2
cvi9uUB4v9f2t+XPAFGsxsJAtF5JXfnc3Cq/QO1QhLIQiQN/qpg15N6AfqZjWrDh
bHfcozUUR39VJicLUYYOAGJktw78XS0p1COYLJsGmxstp+px8zMdrEYtT0p6VtL1
eH+NnZIrCOCcmN4hbHEDI5K2MzVwuXa75j5GsxDItqjWXzdDxaxtU4J8Rc6Zo7AW
DtGHDJTT8lvyINC82lS14NbZkH1iLKbjAs5vpbZx/0ZaJ27vQT5+1uuhpSJieOmP
ar64Y8sA9NYL7qL+5pud7bAabrg/pp/BgDntEpSnvu61gcUZLVbuQbRwaP9VqUqX
TCfLUdwpz8i6XSuVg4u/Wml70m8YhhTriOXWYoqh4lDUAWzDBYcnIdL14skAsRjp
5IobAfT2OuBZZM6B/9ieimBLUdCtsVuxvMyx3bXwx5Bsa9t8cN7cMzzcXLgIB1fm
0HK37FFZ9CyTbwrsQZAPFEB0f1+CnNkJX0GE3+HFyZ1RPYcC+p9jvBwJkWnbIuZf
fv8xQbTurV4esTimnudZ+DGsgu1+jtVKx//MBENrv7lOUAQ7AlaUgk7fV8nR7v62
42gayrc7+e+PYDXzQ6TfYEeNYdCjovKDBRSlzgOsgjV1CEMI6Ts/3+SU0h3YBkTu
6jiXdr12ULWNKskPzLElWt7pIsvU1m/QTQut5DKuJAJtp8zDfFqzj43Sm3gTMOai
uTpqG3F/IKLKxv/fUt7Pvxr3OjC/OMrXSOnF17ZDRqv/m4W06MbiFRHvrn3+Db3W
M3W/ZtUAFc9OkIJE7PAYc1XmQ4Ey4FyoCF1wZkgsZAOobrAO+CnhwYwr9RDMtKzp
XAqQP/jwL0PSSaITIoUOP6sp3/eiWzDq9cYRj3IrZzRp8n4pHxIOlUtRIeEBxYl2
ruaSvg4UyOKklIhhSXYTbCAdPHbUh8W9Kh63x2kL1SJLbwp8nq283EAsRpHuWNoI
tzM82m5CMJu6R8HpRk1BAVwUOfD1r7U3xIquecqJ9MThnnCyVLuP7mCxrz9foDZW
Ut1jMSlVjI1KVAXUjFOUtr4XEYxyxRkpnVGbCx2VM/rIsKdLudq3eBcgjsLktqWk
GOdNHrpTul0zvEcJ/lwicECd4XRgCTv2MsfOkQ+WOv1Q47T9R042rdiV7WFpV7vu
5E0d4xoNw+Ii/t/nWPuRyGTSCIpB/jN7yFzhnES1dYwwNMoTA5lchQ0QXqTQRsuN
Hcmf6jTi0Sz+7LEeTpfJg4/viqmzue8fp+1y/KLB0wXjTE3AnMItxiXwwHo8ogiY
HLQXt5AM0jfpHczkn6qKqayZCQkiMp4Q+roqRih3C3ZqMy2xqXchremIlSuE4pyy
B5lWlj4Z2oumzoVqH7FPZlI51de0vS36vqjG3Z+F0CMdOswczNgfUrcmmH1eXyDE
U9WHOf0RYsIqI98zCLsGyHXCymIz6UKgd1vxeiq00PBvRh6GK/Y2Xwk6jZ5a1QDH
4Ithc3yDgZKbLfzu2BV964Q1VRCoXMculBF4pdGiMBMf8zkRthFky5tjgWWoJGet
7kzQWXeyj9Zp9lKXd84l4lNVm1TqNpmA61I8ImfbQoqDnfrSVpgvb6zaKBzX4aPu
g2czSQpw7XLVNhNXwx0IGQrdvfT4J3fQkXExfYIiJuvvcMdGGRCCoWO+5rxFXtwO
P8oYYWAV6ViDtdy+/sip3wHSxafH1NsJnFB4Sz2KGYRuNZmqDSB7/OtyIcA4kuMk
UNS2y1sc761s5VMPjxCB9bomda2h2L5ofIdSXMyWUZZSACagoUj9baYael7ItsfZ
rHc2y48n2CcEpNkVsOJSnhT0jsrVmczHaCaAW6PI33brAvnohwxYIpZxcT0dXCo8
Yq3YeIUmd5+RVSDVkmw/4jOvduA8AqlB7yHtnk6YA6OtHeElz8pbymDRfAyxmFsO
/R2zc5t0vR8wBJUFnx0VsfIubq/l9wqmQhoRmnoXWRrE/zdTNUtNi97diy/iMwmr
j+DpoIoXKOgaXStIF6L9dIw30stE0rrduI5MLe+q63XnsU/llukJ4d4xMojOZzge
T9rUFhCmTyxmx52rwlCv9dzqazsjqz3WbIhTb+zYgfj8vr9j5DJJKUDeTBu2J4pw
xO496pCJc0VTrgwsbpzOz3Zbqh7rbgXx7U/tdqB98ck5L+/6N4XlpgD07xpVsgXy
haUlezzzi7xdUAFG0gRrNEezfzf0l26n4f3ugikd5jiEzsgvpECnAg7ccfU18KDh
A7hm7lW/dZyPE/Hc3Rp5DuDlVAuQmmVa1dOvdYVnxwZkaUOc3vcYTgRRGgAbj646
eOTvf55lf8aMy1/X7hKKFb3fooyyrrFOXANKWsC3z52E5hFA0iRVqj0wXU4Yuhc4
39Pt4dIRHTBzSDj788fifJLDN/X2mJAhp6QssmTPXXPXUR2NCltuntdqWyYrPNy+
oTT2YT6aedjZh1ZB9a3MEImadjfdjZS2dXnlQYGPZfBQJH4Wtjts5fHCifqbzgiB
/dlZFaKQqYug4RLXfU1u5ZQyjFS2UrA6xEIfMcIyuVr6l4l+PKQA7PbvnBDkUotn
wswY+hkG3C/nVCpgqUmcyYhljvkvgFJT7JpxJmx/SyBjBtTDfLgi9t1T/NyQdQtr
DASulydzlWCz7rho7wRBVX8LP1B5D7Gj76R8SmmPJA6qHN9xqjoPaS6z2TQe0aHh
QFbh3MmKX53EG6JIK/J4p5FLBBAB8vwDJHtOOJQK0DkBIAZqLOgpKf/d9yrpo3Ib
c8Z7yVJVCqK7USMcAgfAntfIWU1E0q6xqdoM3ykxKOgptW8Dkv5VOc/jGlurBfFh
Wo0IPRg4Lh8EZ+1nKefXuqOqNOxw8FO/qQg9ZmHkmGMVxQdKQNnNhntl1Ngn1Sgh
F9n6dMWF0MqkifIbGBF2kn2Biwzk5Oe3kjpFotZL+HdCwNFdSoFO2tBH9fXeF5Pu
PYeZGEhG+PcsgxDROLpTQjnvytzUHR8WW6dmTCwJNndM5vsTxGAk7eXblZqZuGH9
y4eYKqdVPv4sVyJ89xKm5tFmVUVI1ka5u2V44kuEqpwwtfLEzQlVjmv2JNGglQzZ
cbkeyuQlFAdVcGUTf/ckV12xpLa+LItEsuXZTkIsnUwuCBMxhSgf6j55zaVsMB65
Zc9av1J+osd8fMC8Hdzv4Qg8R3AijcFzUBkVaJboUAFwgEgq5Mp9h3zdw0Qxg5yl
znWi3yqhnApDYzD5HYJnTKLQ6+4+7HL97Xu8Bxpmec1D0NylVp04i5+8wUSXU2nC
bHfqofLRQDeXqQJ4H0oPa+Tj0OncfUhzXexaD4eC0iHYuVpcrpHJItMnx/deGwUV
K4cxlqpxPsG5DiLXU1OCM6MX+JQbxqpk+KCMF07KDpKtNlFJqNvPLTAtsTFOJsKg
UglAOo6+vudPP+vbT8srDh7yp859AQljO6LPT9m5kKw1Yyj/6BLqpuZJGfVMFBsm
ZIUZXqYYhrLqFxjcvrNLd1sFYYHlkTx7ZRLKDXHjZFbq/HZ+k650/xIA/t4/E0OM
RBjuTCrxzcKGPAVCsJ2iR2dxpo+l5SeXktECE5Po9Xqw5uosifChNfzbKSKej5JV
uc0dp+SjEsiSNa0daDlSpWJ37E0TGuvMAHRIV0v7HZ9u5sUWrSr8lBqfWV8fxnyr
sVxqHDPZfPp+aQys2mRpUoWCptN42DiXk9hF85opKwp5Dr6IU19XZvv/uvQwoT2w
DkdQJLPAloBLIn9ILPFlui5OBel8QX7ViVziHGIi9Ak1IPUDiILttlsmPHkohgd0
CRB47US1fC6tI/Og2vo/7IRb4QIL9L8qr/o2pZGXEdlbLvwBdTzdnE3d7zEqlu9c
wOciZh2oi8XSspXLbkndQbChhH7HzAaG8in9ykFu/zIYbfi5P0+fC3rV7XJd0yy6
ZAOXwsKslCOVX+uqirAeUwwQnCQtYxW2/cyTH9YzHWjpshciPqLW8jrtg7WrxqEP
FA2VJ7pwBA8kMvfmVXlnIHhfr8dHhXmJ9XT00MRCoUwMgkI+fCfb/Sj/PRiENjoq
OPDGttw/s1yCeYvRmP01E32yVRwAFmuLhgEwnktk8G4UlZY6fxo4sOh+84D0WOs7
Bp0y5y7voWZyjScaClt6CyZdsNnZElS4mBeNTaOK8tprvlfFpN9TETaA+FUZz+Rs
wejKJIeezuNOW8y937+WtFeWww5UNTnVZyNhE7juQ3tSBWyAg+zUh5MUKP4WVUEx
tpu6nA2ui5vczyQU5yLjf4ONbESn0rzg0mZM4RXrc5AScEczKD3Z7198Plo+/3xA
A/nTOcTier76fILaRrRBvTVbUJY+Mqp+CUIDXfn8ykgXJLxbNiLV3ZIVPiaaYJuH
2uCanpCU+3Gfn859Za4JkB76iuYCKeBmmqLTCpo1+rikhhz7Wkus4AJWP5NN4R5R
OjZCiKB7bYSx6tVb4KSEoWO9SUXPzYjtk+ScwnRwNC9OYq0480QxLNZP347+j734
Sr6jG2sIPFONBH+jpi3eJFPyQwb74qW/DJkUrYrgNi5Ki+1zKm7lzKhSavwjaWk1
gfQaXL2mGMx3hIemhiQDWVEpDU4INlqnV4M9nrUu35mx3qGbWWkLUxjpkDg5vWEQ
KffglGAk0edhmsIRHNwwfJU2L7aBEDPqhUvEb2TuE1S7rMe1Ka4YxW3dW+enc5A9
hs9iU3YK04HJwbjER3g+lJ1uj9qs1cTBBaD2pOKQNPzw3MifSl7yNxy4lzzjyVrp
pai50LxM3+KARaryuewC8mxD2S8fPe7DBi2zrCfv4O7IJSexrGuEeCUz9/sBydm7
8YJHgg5C9Rs9NUdBNZFFrm7UgGobWG+wYyoHZCexEFKfrWU6PszOLdDvWFczxAGp
H6iNin+9slwNYcYCskydNAm+gbeqd8fd5CElH5aQ4mdKb5cNBtBzmt1ExltysXap
X82aDd1lhjUNjQTTDUgQ2+8VOtwbjIDQYbZU+s+5WmSoBJlHnj72D1EIz9SCyZE9
J+rQU3wqs5oWOtC/uI+wKg4MuH2e7MVjDkCuAqURP0b5YLU5HrGkiKAVafn1Uod2
9oD3QjDwJtbIdcSFVOwRt9GtdX4RtyhaR5gAZDENnF5yYs90Cc480bBkPdb1RVIx
NJT3CG3YBk+IKA73nAmAW7T60cfg+tQCVmNPp4voRHHdIPTZ8UJm3cxZQthtFC6C
KCGeA8KB/iiVpSl0AH1QQE7EE+VbgfR3mtLG0OC9mQNPiY47oD2p/PjB4l3ewNqq
HD4/A+RjqpyLb+0kjzRRI30oM/7D4eYs71fqHYVZpLwP1FA4u2hRuNdbKLgKAAS+
yjaZkvMueazSgtzf9oS9xEgyBI/iUNUyM6CT/6fW+2U=
`protect END_PROTECTED
