`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlnM9txam0rH+yMXstEM1s7BYjDVlKlfg34VnEY/NXjCdfVTa10BvSKwIzX/7mFj
jdH3NpfzQB/uqV9r9kTZ5xKBKhF5hx7+/PmHOn05Bs8rg61x2OFnFVX5pRrRD2xe
fqm36BS1936mmTkLg/jUBsnLGduc3Zv76YzPbi9H78qwaZ01Btx5d2oqDKZ1vUK2
pDQ3oE5dv6oV+TkG1zYUZiw5HTOzTc1vEAAjim8zcRjAuHc7XOSiozsv8oRO5XSo
XP8xKCkaj+20qLwFaloovJwk/gDjpfwqVH0lQnqLu7JOG97fS5l2yjCnnmxN9qww
9xhdTgNJx2KAHKm6wH9VqqFdgSWxYGQARkbb8T2/+gp3sGwfhEQi+7fdhvb0ZWBU
ZLZrb7rf2m46InxvcYZi9cwjh1C+WBjK4v/LHBjgtayxcvGSvE5lUsFqov8cuZsx
A+C3D9c98YrjLLh5wkYzeZqzVtZ4bhDpEhqiMmk2idgBtN1MK0GDC2Izqzu7McdD
IRmiDN5kcmR/pqvI20Kt1Vpe7E/iUH6ubGB3N/epkVD9BOBFUSHG0Mw9L5Q5j3q0
aBiNzWGEtq7N2Eqf4AcKQg==
`protect END_PROTECTED
