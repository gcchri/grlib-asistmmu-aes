`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m17XqEP45hDSAqaDudXNotEaGgIiVtplo71UYsjvWBXLCg/99QEdzZPkjSCcucoM
uXbAZvxbCMzVLaJdx70IC0p/te4BtvPw6iNlO5MBXuBMLrnlK0f3UwoV+Lth/bU2
S0+M1WwECWu/cK0/NmlCHMwjHe2uDrIQxJ3bItYrqaIJfqaOVtsgCsdPaju+NSz0
iH+y8B62kBwL4XooYmKwWxr70d6qntlVUjho+ulNU/cGy5WEn0cy4Z/qADj+GmJ8
sE6ORnLk2XzPvgdCmpogJUBku/juo5HYoWf0RcEGgXMb+pXkpSUqAhPR32Xju0mu
X8P0xbjhiAXAGfmQnM5kl+R/heGMuUR0NbuQ1jr32s5RUSILrHb31OC6HC70Orp9
pEQAo9kDlbvdV4s8QqDs0xyPICWuMnXyskhx5ohc9Uc=
`protect END_PROTECTED
