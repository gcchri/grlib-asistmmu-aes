`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kK6WqdOonvBuxaNGKtjkk9QvRBfjEOvdDI1Qa5AmJWtxfrZ51o9J29hgFYEYOUZ7
ShJTkeBSBodhqKR3Mlsigs+LpuG+iiAkcn+QZMsFY4cOVKsPe/+oxN8P8AGHcOYo
80NgLiQUcDt5wUgmktCj6UJqTw9Vp7/mJ/yErEqyAZnVu+J2qCpM7rnFOZ2fnfxY
P1FIyekJdOgPYCyPcW25SSxNXwZlq/PWQeYg6l0mSoQ+r3WnQetkjmK8b6+4SQ2M
KmaApzHKuEX5zUVucVJHKqXXkObVHHqhAK9BRRMm/eLgmYEEWKudG0edewHe41zM
Sc8gwKdQQpUf5ImgsRFHAbEkHn1YGPY7a2L1a1i5QAtfpJBLP0696hD64lRViTCq
IeJOt7hSzkrlEaZVjZUKFEP+5X06SDrHUJKcYx3L1CaJd2a3GMj6ykdbKr66uiwZ
cM8xjIj7QwbHI5OkOIF8fCFiv2+Ix/GQh58uX+mXlUQW8PGOXPFRZIz6FGam+0ah
kwcA+u9eJTybCTza0tg/5QseRCv5EQlKyM7XqZVy6H+/FoQr6jLUph6MR+TogSrW
TIyPtD8lv2O8LW0m1597ajQtY/oNcVJDQ/MF/+pDdfPC/mz1RKLutyqOTYQIi0Pu
OOjvDSwM3gLEU4zngh+CpuwQqx4xc/O2/i9mwnKDcCKyTXwSW33nuRJUgSF2eewH
`protect END_PROTECTED
