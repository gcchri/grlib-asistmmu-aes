`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fo8Bch+7i2RwW5Jn8VWMmoXU6VQtgLsQifNhr8chPoSQTdkksN/i7lQI5wnPPJcm
/hZOY3CuTMcgifJziOL+uI41VL6fMxVfxm11X7WQFzC+uDvAip4+h4SegUSt+TCp
bmDPhEyFfCTSjP/SMKoYeqsDrUQQPbtugmZC47uooU48EQBlS3yJGDj9CAjiS8Gw
EuE55vnQZzOWMXGVX1Qc95WHhQaioILLAnp06qSNP5Vb7CNjU3UQFmDejzvtAYN/
lEQILJWQQy6bAkB5Ejavo5MvSLWocf71+Q02io47qPauqruEZGq+fiV2i9VNzyZr
x7cUxigLSZ8u7iALcMR8spPRw75RG7FvSFpgPozGD8PzZYM7Lc3hku70nrnpuBqI
zqiacUX6i75MmwcXjZI6Ji3pw9uUEPqqCewre2Q48S/EfVhhNRTXt4Li3s/11Wyd
`protect END_PROTECTED
