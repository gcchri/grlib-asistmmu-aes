`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/NXwJWOwSR0P//TNJq0MnzKQKpYl1vu6fCu/eMNOUvcK4BRCelVN7+iV4KycwIOC
s4ZUhEFX+nVrq5zGQ2h5hMobgP/xJ/oI60Kzl3chsqBk+ycSEBq2+E06FEWyiNEK
hnySrMl9CKKFvHyEv2phSDdYybbmGBrE1WZFxJdH+BGIMK6bQYnTkl3Fzo8vREur
jq1Q2eSoxXwcQK1FsL9O4bg5WXJHmWPJxKnXoFLOCGyEeJrkY5/kBigGhCc1gpP8
ZHDsVrgURDNiaf7a75Xi7mqvUnv4rXN1+PV3zj2G/AkA+UAj2nusNPy4i+9Rp6Pa
`protect END_PROTECTED
