`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2KWzSZpgNzfb1gnvxJYbUFGD4WCSOtHEo81Vm0qQ628uSDU4gv+I//dsOerude7L
BWckbSEEJSHJ6b52MR3HT9g8XegYLLiuvSLfqC8HVTvojuWrrcv9+c6sPXiknYCY
dr2aoft7FaESJq21otf1dNwj704JGV+V5mZvJX/kwitqDuaw7joyBO+Fq5noj8kD
U0xfMvJzYSRT4b1EaDJ8KnI4F7H0gISvFInexJ66hwqV+6KEDXoBGyoeSVDBh1Iq
dUzLCSp/PCQLBmuqs5N2XIgQh9w11vsvXKACl0rYXZExT5uHqpwgm8TtszDTA06X
U1wu6g8Z9ZLDjYvOUHHX1yjBo1KvQhBzTY66LSVcW0MW8Ex4u/EVDe6RaBNRcXwS
y31WQVSsS4T4z0owaEfLvfMfWeh3kLltuxZ8gSfp+NhEXWfV//ejymhSOA0st90n
ftPCT40dylWbxkxA2Y97G3YhU090jDHBNFgarplMOcd+u18fjS8+bYAzrQOmA866
zvLv8Z5+rdzODB5p/ml12TtitWu0prJ0CZ1dBnZ8PF+ucyUNWnyHLabF5moNj/cT
HDytd+Ic3EylJdPpIq9EUcf4eoA5rdqPlXNnmHpOj+4M3pEDRJOFnfkMy4G5kxx9
LtU5NbAFwvqlnulfjhrfENznNHW8xHzkMflHrvV91JXnlzXzAuWEtAD5lfVVU6S+
cXBasrG4Lm87oK1SiwvjnMSop1qIRNvMQ8chZXAxgt6AdPt8itLT4VPh/PxdabbL
vboi92tX5bB31ftXJiRy7VTIuupTUce4GAQTMZi3aizSvJ5Fh147wXZvufEDBZjx
FpVyWhcYDVJ3Cx2DfSKUzZgct2HbcHMKg4/7C1obEQmSb4j1xk4HqzxnnGf6CjMI
F7MCBfp6H6wDX6ogHxptzhvp+yHtNDRSNy+PJ3j6MbDn6TjmaJ7tcSMH/IgoxsvJ
woPzKEKoAGD0i9kDfk1ydH4KMT8AcICejE/4u73dy0l7JayveE3/TSQSLHVs+Vp8
AySTMX3xPyTr2lszkzqlcG5tKm+E6XDPla0Ev0FuHD9/+NX94Tax9hKBV8PZVuMv
6gYAQchzFN6pYZ4g3Krshsz6z4Ks2nI1pI09KKhQ62BZtDIDjm/oaOq5R0VAIHWJ
0rI9OSP3yrZxJrRrRgmVdrYC1IaHJC/pmroBPT2CkIcH06DOX7uSlBsM8Hrp/Vlw
ehDLLzfRyYZHnGBRIZ/RugS7ktEbWSz7jBwpWkEHKluSu33H7oxh2sVn/3DRw941
xV/l6Wz4YZ9YydVixp7EDQSzQZoUzrvCyb8IDSD00+5EoFpgwqHT+26QdYkX9v7H
9aCNHXgan1fTRUUfW5i6tDukgQADafNV8E7GL3+iQZBFjo5YUq8mJ1EAKh+7hNsx
k270dFmvq3KenSZmK0/1pMaNhjPhhx1gQZ1fk4msOZIdahUZGYsYW1vtViwl4fnx
uGIBL9TUJVDD68Bq1SqnCyGu90z8vMkR4uC+EuY1Hqe8AhsqS4r1uQJIY2RW7JkA
E7L/4Fg2S6hgO+imIcpEi6K0V/pbbGxdAonGC8W1MQ9Od80yMsoRrBzov/OmIjFk
sazHhERcmMp53e4TKIr2Qq5KTD55wLC2MGS28QdqRr5Yl1cY+sC7nhYF8zV7p0iP
XGLjWKDpCIuwncMnZxQFJPyM/62w0J+XKnbu8BQWfPq5Ez7rrBpwB9+8NUb06ZsN
9vEq5h1Ima9EGN5AEOMXuXwwgbdlHMMR7vTEpzrLwlrKRBs/KmgH9CXNtHswHXxy
D2iWT9L+YUmXU57/NvxxFClv5EmicA8rxPMgHcTU8LNwxcNqsT8sStykO3KCbhIM
fFwtHxBusbF8AbyfV5H+g1HaNa/pP/HJp29dk85ZNZ5tiv3hczrCk5XTvxOXIhnE
puMAxBMRk8AzghaI8ouIpNHHoGodiSXWl+oSLwG/9S86cDbrx+Ca2BG6JlPNb+IE
0B4wbW47fnyehf5CAq4PSiiJcbSEZPr1j/78J7tIxOIL5CauCJn7DAatRPTSSVug
WlflURYgEpsMwLJNqdoBsODrArVd6Uz1nXgZhNW1rWTPE9akonCzwrZaAHO331V6
I86nLi2vUez2fNG3T+xyAQYjwvxIkWewhWKycUGQYh8YF8DsWFMB9t76EoiMKH+N
XY5S/WCE/dl3s3txcgfkt0aXx3w5c+Xqc+Ctn3Q0J3etGi1Cbcj26pgmo3kd91Ko
eL9u0NP8fXPmHVPm1XjT1tyIKkMdxzzdNuzAGPdilMFZhlUDhr9+VO1tkedr2saj
g9X0LFzF7M5tysrp/FaRwnDYAWxn2KhOSvidaLLi4DI=
`protect END_PROTECTED
