`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Of0wjXKWjNH0BlfIoy7QN77FSgu1qcYfQNCdUw4VR1VLKhNHeThbDxLHhjmUHhU9
3igEC7Od5n/lXN+GqJYvogw6d3vA7JkMzIJhowsZRG53dZf3lQ2T6G6Yk1Er2xaX
9ZSeL5socjIY8myCHH7pYRdlpDb3HgnEaYtIUnn/2s0Lqxur6zX6tYo3oWwuE3Am
e6TAHtgl/cXu477sOz4q5s5fjhpO6x/9064eSr755Fmx7wYO+wbKjKbLcQLuJVCH
6PGFVcEWjl1Z38hjUb5IphItsdLMpMpDYvMNv7dCwD34gIbk73KumCtm1XaCh8M2
/n3gl8WdAkXgQEnjujyzwEPt/ppc/YZXWbz3R/EveufbFD/M7de1gCvPigB6iZ6b
CphDxzbb/0EHnf7AzBysLg==
`protect END_PROTECTED
