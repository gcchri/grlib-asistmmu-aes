`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pVhfnnoguzlYdWFCDm60Mifruq+i+eMakrAxajNo/kQ+26WILME0pIzc1M8jDaHb
e/bgi37YMvPBaXXvCpkwRB6Ty+1ATfXLlDagkHkgMG0tFrKTiqEhyWVsYtcwXKDB
Lcj0tOlr0k8L7NL2NN4JoWBnE8IcQH76KSYQIZssBebOSoPoanx1mqkjU2vrvItJ
cTEawUX9/Lf2IdFPRvXFJRlGzCGRyWRdmR5PO55F8uVpGRCUKLpu6KW9Q+WU9Zcj
m3DNr+JeY9Ptd9zdywVF7q6x82Z6OLI9eACz+5hxPBeuJs+S1J5mWlkmNYw1F4pG
3xBzmbiUKcFDsXEJsgYrtZmimN3Kd5EgxfXn4LmxIQRSPNLmFcIAyMm8qq5Gee/U
KA4zNEiCh0DMBU4ILqLYDLG7Znvc0rXZSw8U156Pz/5/5srcN0fbOqRSjrBWPQD7
bbsUQ+tUUGUypAmRH3s9IUy6NhKw+cvRm1g4x0MbYQZzs0CorUaJpUiwcjEYAahh
+eOHFo9we2MTkV/HthP3StXpe1x3p19aXFyfBO04LJFqXzhtwW8BF9NRSnsBg06R
kIIhhcFbS/ifK08ej98hSPTZrypom6b/kPEppfQpNUHeuDdlOrE36IXKmAWHlYe/
tOK6If1vscz78BnzmvE/3LVCnP2pfNZ7Nme5GEY8vLc=
`protect END_PROTECTED
