`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4bXxpSWVDqFS9webQkNI2e1lsVCbSA1MQU4ITLTqT7v3Ax2y74LWf7Sd1oL1oIry
ebkmw/mcMVRcPvVicbWKOlQ0ZMZi8Z/7wKFt9GTDd0Rg37g+chuj+lyBmmXHTfVK
RoS7DlGA8KRCQkFTjR39S2Rsgb5iVqH/kkLVm70V+FfgQ/9yuaFnUtxwBLZr9Hof
OXH76io6OjA2GlA+ARf8u2MZcgGoWTGXTfQzjzcBMh5vZjqLBxtFdrK1uvhTwGl9
RofnGjnGq2O03sk+ZRYgOir8392L7HgoOpofSte409tCtsgjgLJ5lmK4Y6FvkEdm
if5/tWi3jS3WlFpoouu4NJXYkAqBUp9ipm2VDLl6t9iS4u68YGC6s5EIZ5awkkyK
GZj/vFQc3g/uPTj1HRxcViOSfxMlhgnzkbJGz2WAR+AmibG5t+9uWOd7hAbixPr5
ea+TFW2t0TJ/Fu8cU+D9UCW+6Z+UDoi6M6eEGiACievI8vZYe41jWUjt+4pxYv2Q
YkTff/x2KvPt4ojswQ1HSQMoRBQgFJbyf4sjBra8lhZ881vfOxjTg4dYApbeNrHm
QSYm/4W3x/HT6SnRd7o2YFYCrDWi+eFA0H9UHELsR5L0bvqfU9eB1ncaBto2QKhZ
QzhoybVTjvALKVT/D8RD44ElP6GcI0yC1pmbW3PXKZQTdhqNsGhT/i3XR1u9ZMlM
/KqIdC+WVLTv/wsRvwhs0fTKG6clyBUg1glxVrdYlNZmbQiLNROozAdF2GE1Q1jJ
zQpzigJlNmyFp8oQ5QXEcYWLAQnVdwm7qQDjElB0XCg=
`protect END_PROTECTED
