`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7xzUnhAJtm3oO3vhFI4X+QDGf9g3jMnjFXT21CvzuM1DoGuf4Mkfn0lm0O7PF09
WH2gGiV7FfbSF4zmbZRBnhFzsHgrbsaNNlP8jDjG6+mi0CWFNRU5vGw8cnAeO2C3
mqw7lFLf7duqJXZu+QBEol6PQDkuWoYyGT/Tbmva57O3JP8t0VSfHQjimqXl+QDz
QA5WV/COol6yTTvt0A9yimwnZhoc6TatvghcKZwQWoG/96wEM8mSm0AZmXZJXD08
g0WtlDGjzUJl4oy/GUCntg2PLzu0kAcLK+qhZK/DoYHXnFF2e+Y7FLGmaKiEoa08
Ob28OOAGTkdKIzU3ThnfpozNKHtfu2yKKBFQ1dLE0edVnCqLmr1nmeSEMOkP0FDV
CLa7XlHl2PJH5xNVOCJQ2G+omZpGNw8AcFGe9AhFWEAof46ulK1dfIopIv0j/aA7
sNdWoidyX6YZC8SqLb1qrXGvv4tDHsyx7pNOkCm8s1A=
`protect END_PROTECTED
