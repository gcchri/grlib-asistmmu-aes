`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fV7PWxCkbWOIwyfCWVm0bH0Su7mwGicG7Mvz75b0+a0+6s9Nwd/TTGsbaoeoz0SX
mhflyBwE64Zrq0kygLZEzCpFgrGCAYQXTZ2fsANg9qCX6M1hwHaUuxwNEi9IN8do
I/nPehrlqKoCriZ/7G6fIuXEhWAK7ws0gBD5UN4OG5HqgJuf19o+HUKX/102Lia3
Ki3UW+vbAAUxr5Z8TwsUWSC8tt9VGKbVJeh6ySlPkjxuk6vfQI4AaZLHwbJLa6p7
lHVJImrc9121XNSuvYUIYMhoT/1tinqEay+3pUB6VBauMCpL1GGCCGFUH8o/TuKh
B2Reza4bP/aO6fRneQlWAvdVfHk/lkeqLuqgtgDmZqgiaUJWFwayt/ysGBzsK3i+
6FezhskHwxS99WhVMQ10EHFIasEKMaahUuZ9kCyEVobgNV1Qc+L/xBSWjPsXOgpW
glB+Nt6aBGBPqcb3SoUW8uRFoFK7WEDaO23VHr/1lAtzrTahc+o34mW4ka2Okn2a
kOowC5exZ3fZxvGCQrmE+zXW2NkWaFEUCd9EJsJMnqOA3zgpgdd5Tu46Mo+TVr7n
HTwIAgubdAK+EypwZzzn9QVMWv1sk4yhEjruG70bP78+T1kmicxCVlkvbDXZcPz6
6Lm0d8oiLzUI3HBpVS/Pm2bQvg31jcvglI0/WQctuVIbcVjU4CkcC1ru4o/I5HJJ
9FK6n1jIjDpwil58AY6lO8LbOKuDeoOb90OZhVlkDdW4tTuuhkuqDy+LjxjriUgi
OEJBGFedkIt8kfABq+u2SDt6CgdAAqlM7ZimJK9eMAXSQiHzFndNWA+LVn0Wqam9
fmuVWUe35bc1emNi6vSdLvc5J3U25dTaMuiCPMQsrkxTd5NwgM+29jVaFk2Ml2qR
uwXwTyum8CotzTSgI6E9gg1kFPYJuf7F2tFoMdlb9lSAKdIVB4RWuXo6BOCcCNEL
`protect END_PROTECTED
