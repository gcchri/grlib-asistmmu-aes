`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UvkdOMTDcjJODvxPiBSnIBcYsgdySCRteLzKsyTDCFXcJOyl2Y4TUomxFXcEOokj
de1XCUnk9JoZyv/DMnbQvIxQ8iqb8MhEpkVUMSCF6c8EKtc1kmq224Q1LCdIEhpu
inZt3Ayn2TI5yAdm1yBGTlp7eoSFb9ZitER8hs8UqDEaS8Gu3HLqQN+ZCAc9KN5C
Hznrx1qpwsQHUkVsLmHIz5Txozhxas/qdHK7XCB0oo7ydv3OHR/J+9FwT63HdyyP
82pAXW3O6Ukf+BjN0moCXaroyiTdb+X0Q8hvmXb+vtjNP/Lf2zKGGBTOZOig6vcM
MU+iWTzeVkTpSQeBQdipq+D34/SCynSBA5dS2QUTcW4TzW2cjxIH7RzLJWixcC3N
lEJNlzUYEKzanUsq4tnvEChYOhW8Fb5vPrfqtm3npMc=
`protect END_PROTECTED
