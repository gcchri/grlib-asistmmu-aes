`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4rV7EyLnDT96pghl+iwXYCmXjtYxUBmOUMUiz5vA459j3G2/v1un4Bp56qEXsq8w
S9cAo856CcAURp74kNvca5CxDuoynMUIrXqtgu+LEPROk4kJuuWXGIF7KksKkgxA
wnCx4IUypDpfQs1632fCYuBFhIg+wJ0AOrtXEb7W5L6hzyLlkOqOHuMpq1ZL426M
qMyX7aXwJnH9y/w+mYYF1m4DsEApaF7CYhKQF+g1FM8TRz/HzDtKMnJKN0Z/23IZ
DxaOyG9Qp1uL8cR410jVUg==
`protect END_PROTECTED
