`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9U1f5YZ4c+H82qCspaDLXnvM9CwXBp4NxXk8kzcFbro1E3luDYLFnuNtjiaA8F/7
d7cNHIxt2kEV5qEkX1uGWGDi+1rVnd8XnPZf3bYGGyb3kfewHWF3n1WRJjJ5QCwU
mhK34jLmwKiYQF4kmXsg7fO6nNlSKQa4GUCfxkpNax10xLTSvLFPuy+WO1YD7yY8
ifus2CHtAJZYKTvpg/Cz0nxXSyFMhE1Zj5tsJsYBrJEoFsubMpfCZ5o6Kel1UH09
/qQSUYn80j4taL56p6GjBnTogQiKVAMmGpDOlLx44n6aD6HQIe+0VU6fbq5M+bTY
wvlNSOiWzQfe+Jd39Hi0zjCI6jiHafvFE0g0RnbLwjaIINy5Y/Hu2uEM3GFhbRYS
3Og/a029aqqdf3OEswqA+psZ4tO0XeVOCnfVVH5/W+aS0QZ4X4Vr47B9swD4FZEB
3yXUdtaHWi7lX/ZPqNrdQgFDOwM3EYHYaveJdNjVUvo0QC/pDvrWe/3Eq9/DnvTH
B3Dq+6tQhxlQjoVywseeNPW5Nbo0tlfMiBFafHiUEFeBxV8+Dcel7dM65aSLqK0r
R/1pAqQyAwh/tebeyc0i6c7QhL2IhW/WnclbmmdOV75GiHV+npZY/55uknJBuch0
OKNAXTMc7xG87CDdfHqOZbsT0FmjFxRB8A5AlQ9kyrk4KIV/4ECi0B7r49MQBxrn
nRYrowCZtpKZldaccpUyWe73kPM/XtI07LhhWzXYc1KdlSYddw2lnz7rV3xu1RpU
gDpz+68T0Cjwz+stE0AOghm30rn1BSI/fAFHQMxgMjXL7plQgkfNTuUtSnxGv8Y1
VRUzXXFbX2RPbHCPR73TYssJZUmsUb0SHhI7HfsBS6iqzVc6sx+XYU4spGizFE/F
PDjIX8vBcKTatGh3/ZpRAuoIXwICnmmZoK1k0Cx8hHfxiLS0ujsLb/LlDSPYZ2J9
35/mb8I/LE71qN6+V0lS+vX8BpttRWy/gI4YIieBCB83TocWLq8Mn6h5pDhTc8pK
8EwMWHqYvVdrozdkBt+gq9UxhM1fYq6wdIDobS+6v5uRcJjdZbOYQBGOGN4MXURo
`protect END_PROTECTED
