`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZzbPkpdBk2nXgNWTBVvDJVFihLMurzNY2NFhjnzHgZhevNIOdQEATQT/64f3HzN0
snbEJQsWQl1vMHA/GiiItdL1ZZSUm8f7GHtR37LoH3wP7OLvIEfQkXYJeo99yYNq
q11ruyEWGfQl4d6TqUnYv1zBI3YtCe3v+Qegt7GLhcON+QI7KIpoEiK+gd+Fa4Pw
Oe5l8eRWjzeCmhFGoL+xKdDf99BlU/fhOfslmY7XHtb6cprwF1+3P3yrxIHX6kl4
FG7N0RtXTVWoP6vWMF4PsVCCTzg4BvLWCiv4eKSDfQ+15JSpBR6ESQOa7ifwJXBA
aZnIsSZUqGGzwrSJ9s5SQbMBVoZuo5H6A7T+y+ZRP5XpW9hncroKfX6EmvfxSbeE
`protect END_PROTECTED
