`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hQUy3+uLZ4CXbfJG0Q8UA4vdq289N5cGUXiLzRPN0u6I7k4kftoln2QPKl/FmJ6k
9xgS64Ckkk7n2P6WEc6CKbS60I6UUVJCtoMk76vJgkBlUeebinc7iA9gJWKmIELf
2lAzC6JbCntWKOcRBh9LJM93EiJJKSPD8nl1vA545Wj11gEdlFfk6VJVzs4xCRSv
fNGA0xhlLYRwZ8jZrs3sYMfLzGh0/i3OmZJUU4xII93M0N5Cr/Ez2uItO9ZpmkTf
10ob69W8FkRfDJ+uV+nqE9GToEsMVLYP09GrHKOXGx/dcQZRLWD3ct+rtBBbmfr3
bSC75/BkFPt9CHrNMm4NSoNd4rkYFkJ4kOAyS5V2OxOgLWeE1jb2qD4xdMamQp96
dPBC5bsEEsGwGX7NDxwSdapLPu+leJoz/5E1JRTkwT8WOuTKsFLKS7Ruy9HVH+V9
6e1NwkvsIYkFrh0VLrHFcmCAMZNera6qLK+MbD+CyQs77OPmitY+3mUAJPkQxaiC
+yA7jHNBt8qrw2M0Vt8oIBGj132QkyUdQf6osVeuKXt4+UfaPKkfr8pz7Q8r6h3b
`protect END_PROTECTED
