`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gw0WT5KfoMndp0lD69pnNbOhcOyLl5t3Rm887A8Scq2DiDTLs2cRVw+euwRv6hC
uWQj0sYJ+ydErjxccFVkNDmrDXCgbfutoTRCaJj6YcOahpaCtvA7P1Ux4F0BIj6X
rDCFCPPTJ/fnKqcakgMSxRhex1HBBXPNpjcpgyfJGYclSRm70j9pHFXXcMgGA4CE
KqcxY2B/Y3vkaETZYhcuhyeLXb2kZstZ9dKWzTPWD9pIpjRgVBwBGmRMkBMlt5zR
D7v+jd/bJwqTxYD1WwqSqLe3AcH+1W7bxpD/jFcqNaHCZ0AqU28LZfSWCUyAvCUt
NucyWzB+mjunYXpgA9qlzo9YmjcoMRpMDAUuqu4uYUZjmkpFlqRgrowjQCxVdC7j
233uBgtKdlRA2PD29mASoCxQnagaLtqdjjor363Df6S9Irq/sIo5jAFxPYKGB4VR
q2Kje2OVn2wsYBmoujjBhsdEvUBpNLQbabg0EWnIwvjvimns3nIvFaQwFBWVNld1
52L77irVhb6RjiJfwBsKSeLHy1Cspw1g6VaLTjH+55T+mqR1yDE/tCyewTDO2ABy
01vgw4iUny5D3Qeu7C9wdxiPM5BwcwV4eppuuQigCXZkQUtoZpPZnITYTnJdA710
aM57p/1BTYFw27bCT1yLw5FJkT2f1uoA2XhBnmMyeE9Ah6KTMcp8zchPVMmiyPb1
Q+TS+Ki2WeyVZBUYmG1XfeFbDM7oyPX4VRiF2J9691vHDbQPvXehC37n+G55YBSk
sTOFW+8z4caoFPuglL6+qqj21+OJAbvc39Byg8FP/ZkazmCqM6Zl9FOPy1IShmg5
zuvZUbU/iSJKhu5te/zvKtrRrhUiaTIyBq/zqadl1avlExBsDBGmsVMNOTomWD4M
AIk7S0m8F8cdlPsxnzaXhzbmqPkFN5a6K5fczn5tac30Q8zPO0wWtyWmGrxjupBx
wjLt6YoVkXh2DICycF9Gj0OYx81CH2M6msD2R1LfibJqOENldYmSVBQ9/0ENRLpO
tlCSxr+6SaUq71VMVRRbFWo/+s7sBmdgw1v1HudlljfUMxymoRjYQZFLTqt0yGtg
D92AQMExecU5d0o5iRazsLTe6Zw5VHOrwWwwliXQy37J6z5OY0L23qrx4Mtk7FQi
fCTKZot6noREeVE0gZj0lsCm6V2rA44E1gbG/2Ep752xLWyBpNdHuJR9gF+LvYCF
FUgGSlL8OohXd6p46k5rwILVWMStq+fvxGRR+2i39ei8gz8s80P4ZSX/6Vk28SNO
HjqUnXHvH1ovXW83iM45KdACRMt3Hl0U5h7wCFjNfmKMM9nyJrloSzbaQoPCnOyu
Blv474ifNnd+7cCiI1Lf+UZN0RjFjU2fdosY37t3FWCYt3pxXJzo/VbgDcMVio9N
6tbEsnOrbPSBvS6DTS9hyI/Lrw+YAMey4i0WZqjj5pkyGA3A4RPKgvEPFeVciWj2
R0GHFpSjD9DE/97OTODSQ+YeaPMdsw45DodsN+GQHlOVrzbYw3a6l0tYGqFX7OBV
y/wesnRs1LSDpph6BO309iOX8irFW44HEOvKxnUCdwnP2lizUt4JMY9OXUZEdG18
hnA1rW1dD9liju19yVnWUYEpUnttpkQGMu0Sbs5udquyrw3L2ydCkUbQWzA3p1Z7
Ywf7erbBV1ggZjc/jEZNEMK9exlt4eKWU5R1WB1k/gwlQ+h9nXe93zis2Kwsgfq9
4xAqI0tlctO5QUl2BLnMFiq6Mchkihdnyf8Lm1YxgqLnrsMTttLGuzxI+ESKDeA1
s3LZ1VZ0vNVRhWwh3AlqJWMskj8suyA8YI5Qj1OBNQ0sBr+RQBC9tpwz1QwCp5/X
kzpAFcQb4/+ruy87Kl7lCD2auwEIo8mVu69LYcq64MxL/+tuB6yeq46YKkMUXpiU
Bzb9T4BAYCHSctqhpH0TJUufjWxytEAsKpIYmQUM3q5rCBjLptP+FyqhP1e9H+NA
O447Cb2RJQDqsoTbOe8Z+9KinWaI5Ftr1Ewk3le582UZzu6pOVMXwPah1HMOQLvd
aQYKwtoPlVlayfd+P18+34ScdokeRZnH8Ca7yS7DaQUfI6gdeeGYjflQi5QQ83bG
6KoBOcsD3mLO0P1jsX3Mu2cbR/j8bwp5VDyzqDynrREPSArySpPQta4ibEBgGdPe
qTJ4IodRpKb6W+kQYBnKwu+KKr35Bpy+59Z7VFERE7oURHhgukdxhJSQ963LGFyy
nIOvzWhNwHGAL2buWrHFK4fboFeGXvLl4/S9bKiXC/RCoRpXmrhZPXvxgs7UUtDS
/4/2fqj4LW6hcEeQ2udj3UIzRz0nxcHCV2RSk8QLnwbwVJM4ttilZZ4ml3J//dGe
exAFQC4fO+PHjU9VlEvxTwOfrF9WR+ThDMiX3YEl/g20VCGRpnpIL60KFBaYIEI+
+pO2NKellscZDQ7gjSNnamgnqTL90FJrRbew/kSNCFXKMd/LIMo6AO4iPSesH+Bc
+5JTZIQ5BD3bVV5Qf1tHvhc3Qb+SmeF4qbsENpuAtMx6tFXWXaM9TqY1ho/WsK/k
uQKtFMDwQjOqFaHMqXC5qeQExrR2Yw7efbi5fUM7CXiQAdhUDj4vYQU2ocNzJJqX
miAuEE25o2XdywmvvIPxjrsKD6qdaEsVtzg9+8ywPlCLYQ0pFTs2xC8sNVo3r3QC
E8bVdQWbRzG/PdNfdaC3tJ4PRXzrPyb5iBT6QXD3lKTajmdkIUC72BBQXBc+6oyP
JM8pEVn4yYxCXrSOxRM1YvKjpFqF1Q2mqV8usoaa07Sy02nwdHE9I+CM8GXGUhQ+
jjy7S71O6rp+0kQKyI/69rjRW5VHU0VHZT3+AqWpXq7nQY9y82vLtp61ciXMGxlW
OKaCHzRGP6idVr+xdosiioqxHWkiwZaovCv/5Dd3Nz9zKmIG/M9LuGKkWkPcUTU9
ihEbgSQWBIp1EKe0KORDODhK+N9jtcZa/tt/+HDEYtzHwFkEQDXB8MybsBA3wXvG
twfblSa6TYndJ+YeTm6VUZsZBSJPiqgt13rNfIQ42CJEW6ue4BJj0INy5nv8Rl3l
qQpK5bFgVRNO+iTgReI+wLIkfxAOFi//GeGEmb6wr2aopsj3flPwO73KEreT8eGq
0PDq8zSkI2AYU7HAdsqZqz27fVE1D8mZiaWHK01Ma59QvkZivas7eSqDBK/7H0QS
FIaFQmE1SxOWnhJnqwHfAq9Chvex607a87orIEn3Av2tt1/D02EncDrGlLZhmomq
eqD72y/URLa4qz7fcgP+s3jNz0I1HDZMKrmejrkS76eIrsaLVSbD0TFPdvLE6VcE
xeC3dADaoI+kpi+UrYKx2ZYPQmEfatQvQwTgypZKPpsujpvawf+cX5pKIMFhP5SQ
4O8xPx2MYXjlVuPiljeLVdO+ilr/ciwnS+B1ym7Do1jkYnbdv5r+lLEYuaYHzxZ6
E3l+q7sBOjaArPthAjILAyy2mzezv945Lt3VRw5Q6C+FdZlDJnoy5/qrqtLu+BpQ
RSkIa1Em47+2uYL7yW4cPZMUjZBnzREdYKwj5s8vqWM=
`protect END_PROTECTED
