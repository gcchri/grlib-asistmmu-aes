`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abE5mfhizK1ePsOGPxS7CSbLwrV5oBTI3XGINGd0GTw7QdzhrbLrn6zmkuWXsnqM
+j7C3LN54fx1VuzBLJLgpTXQxpk6fQfhJwRvVSHJSKJ7dQ997cjxOnoW80myezJM
oXr5Tu2lK7F4oM2ObMLvp6g7ohYMuF+4BNCHhMOhE2r2CrTUnQUEcOR7K902ry9B
2JRW7vi4XtV+fBQrAgbHxB/Mw4OEVJptjf8bYF5y0YtOFyxtSGI8BZ0ECVwhvJ+q
SSvZ2pNGGaAJD3lcZQWDnNY/LkPzDnr3cLB2tHp+J5kpIcZfpRYZXIEClmQjMXD2
z3hW61TAnvXxxrvRlpiPz69l1V9LWdUTm+0cnPX6yoljL6USlz9+srSNyImdsYk9
BaY4dPGsjEcgCBpg6vL9/iAkj4+UDaHIwsXgTT0sAvrj0mmkEKogKpFR8wVDVKm0
of7Pv2CCZOS+x8QWSKXeZA==
`protect END_PROTECTED
