`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ak8j8ligNjN57tuaiw5J7eHIauRVhBG3h+mpalvtXo+pYpYGJMlaYvszzLupJTlJ
N2S0PH3NpzAA2Te5R28OjR1R/3JYwoTwuCyC9/tDMgKiA4CcrcVadlzdM2c7J2gc
U1/2ijY+/qD/kdWCsMJrGjE+mueqNF9Ou0jqvZfAWtYNmiRkLShQ4cqCfwriWI8s
gJPcZvHPdtWCTpZZ7M/BHqGTbyDOEq7eOX1GW53+PlRrl+H9in3clZQO0whYVxFl
ub4l3aC89At/8SyjGG+XCT+NJLgetRCQksPMjM+Hwf4K+LR7Koksg3HrD9QQdKxz
eVpjt/KcRrk6T6zt1NDdisQfujGFSBOS0Xl7AcPRJhSlxNoXaP7m5yTzNYA3yJY1
GRUtPJqCNHxSmkFvNNPJ4A3W0STx2JGEZXYhMY75OVGZ07X99DFI6ChdoCNtLhaw
bB525PSvRKWkoBTDRuwmLpHX6eDlj5NYAgwU5BnESksfowLF7SEb8mybvOra07t8
9VkS6Jc8dTteP1dqCkKn6/G39VHU7Yb80t0xsoj0kFXPe2hD+4ItgQXD8o+L1lWa
ppfjdS8Kttz1r5SletFm8R0cmeFk914XD1Is6VtmwomsQqA26/z8qcqgr+neg3cH
XR21ED1OjHVWFC1SAmY5apKEAirRxhszEYXWr24hz/92xy0XhiD99DQExR/MDDZ8
sTDZ5ys0FIfIQWFxn3SwexyTkHjTNLfrEtNHldj3MJmjxalH0oV9A5KdSbpoYidn
`protect END_PROTECTED
