`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XjmWx0s7QDCOxgNV9F2qhPbPlzzlkHF38jUdaIzNnoeIYrh8CmcNibc6RlSGO0a2
pv0JWXXGJHRQ97YK604jA3PT1znAQ1mrOucb84YZLZ0gtrz+sywFqu3rbHGQMPkI
vVbLMc/GjyCpLddFgKpd9DgMpD1k60amh8QBhMe8xTdGex8IQSr02TrNsARSBmsk
xRFojvTJIlBMzBlC1mV+1JRbZczWv3AR9XTPDGjNx0Akq9gOIKLOeehTJJ/FpQ6l
oQ8DzzqVjcsC8/JGtAdIKgw+6ehvWk8EMxS7l1f9xeMD0XoTzjObUQA6poIM38Rk
SGQxqL8KD6nExyZrlzLcGSxc1w5R8bVIM9Lnf7Gox30qXMSG37YYMPLYOMzXhGjY
M/pWizBfLIDPhCdRoEQN6QhqrTM651UWUIKpufoJdns19AaBVgiJ9qLzcpGyXLse
bj4q8jbq1nT39sq6e4HZhFVKpGrOvfn+aqTCuwJVraIV+lKVB9Yooobfebpuyl3O
s5xzhEUJK9LeQrw800eNhIpXh0DqJnN7F5pXh7k9b5sqMdqCPLdCqzVPzvImenu/
UmRlWkIA/P+wW2GOzCuAtbi2nx2BO5sSfd/pbuJZK1rMlyzOi4dQri76oISRRKp4
CJVV8qWuCjHjbG+8AVRPLu2ty/sKTAS7rjDlsjtcAt/UNSHqmhhb+icY0ZTjbuK2
HWvyKXadWaimedJWBzLAiTQyIsskpm9KKsXH11yCZfHUaDJzTgnkQyVd37wH29pC
xBbiROqPBBEHKv6j922lQOIhUBbbk7dg/imNtWgTOaSOdzKcOTQCtF7EAw6jJBDy
rEZC1w4y/fdIN55GmKNRjEAOhSJQagwlJh3hjGiit25n/8roR2tk5jmZyG1PFS+e
w1yBuT2bfzf0HG0zhNikp6EtlhFZM643aq8PWVtmX5bLzvd5TbF6nteEErUVrfxC
jE+TR+hWKmP770UGPSXCMq8u4d0PveDZKbyhrKO+U2AJMdHelxQArx3Y3j429Pd+
WSie9IRpyIamq7ACjs2Api4FE9Lh4C8rKp6gBTF0tm+Wnt4GoaUFsQJkmwT4SHTe
+pp/1Wgw+/IOI2sXeGR75dop5q90F9lF+QW3jMnxF/Rx894uR7FVeoXUNh3vC6SY
u9iN7D16tuA7I1m9xyCqBggCRiVAl35IfuVd+zE8iexbRaeneJ4zYz7CAhdZdSnj
0mPG5DMiT346cA93ClvWhFkum9An16kIlZd3uJKeUmBBkWbJ2Lf8+Kc09qTw8ggd
H6Qouz7hkR0iNmmj3hnE+uaynzZyWWfFKo97sTScXH9uJp0Wmvg1z9v9+dcBr7Zi
x1mKl7qu0Jdcu8/xE5Iquy97U26uUY1Vc3/w7jDc8kgDjgRYiJl6JVzAre7ugWYb
VHEZz3LnWwbp2493xYNP7fZoNUjD0XvzO4JvT3NgRFo=
`protect END_PROTECTED
