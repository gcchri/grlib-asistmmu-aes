`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cnhZ6YgolEQ+fAFErKutHHXceBnVGblhXJBSyb5aHUW9JrzR5Bf0jwFpVXDIFhtU
D1cju7k2+lfkUC7ri2WTfheIzflwfKPawQgs3gFbsmPkm4x3AcgPSJzzzXK07hKt
56LDphLm4fkP6CgTGHwN+aJyjlDG+UJlcXCK5KAxNLV1PgSLXjvGCmYoT1XvqChA
vTY7JGAqaH1Xqs5GGl4XFe8jnj42hZ9og6q2iuwC3hPyYK4DDA2ecJXqleX5LOLZ
woEa9lXL9qqEjjA/A/B0UeIlTlF7GTQpttT2u+rtqiVw0pheFPK9p6aDVuHQw3vJ
uaH0bc3PFNj5GepPT1gvK76oJjFpBEr8Tkgc/dGaSh86HmHJnFAhCgOss6FvaqO1
QCw8LeYBynB0J8H3NzNdEXoz4pi/MuShlLOKjPTLHpuAMd+l0M9CaE1pSTKaknam
QX2ypHTBk+gebgdz7vtI8JFlSksYzqT5xgZYZ4hJP8xQtDvnuDKWRbs38O3gwC3m
YtPKfN0qucqxOLpDanZw9w==
`protect END_PROTECTED
