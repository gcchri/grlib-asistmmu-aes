`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jx9qsR6CW4Vx/LYIRJUGmaAN6UPvs7jwATuoHvCuFsPgnVgEKT+h1oH8FLO809CN
GRADSfLlXrktnbqJc9CKmYIorQZSwdavGRUVYPhj4jhD7vWjVY/IToZteXjetx79
8gSqXnGZxgFhz65Kg2pXN3BXuIlHUuYUwuDRWYppu2VHdHliCthB/O58qK4vCjdD
3lPJGjrh5MbXcuBYX2ZEttbolqJWMcOR09jrmKyU2+L53yqiLRTYF0GxpmvJkhzE
i2t0Dg4p1Y1xulOEP4U0r74MLSm7Lf2XU3/qz40Sl7V9+RY5w4W/U2D8jaAx5wx9
xr8hfTPodZfB0SvSFlSDtT0uoQ0YBIl53T537IrLX9krtcRHM+PEWrqOBjLT4wDT
jVo5EBYPZKkNOFtSIheO+qHYUXnaoWVtzFT7LfhcjW1Mu4IAHtP9vHv3N+dcqNgZ
hB86rUPxcH0yEc5vusi7GncdKJPW30mD+0jkDsOIOZU3IYRCzSSsRnhdbN/l7r1E
Jjw7XitOH2m6T9ZDMMn8++sKeAtZWDH5V9MLXFAo9PYSSKf3mI4KsSNA8bJx/Ys0
VbOKUsiCqeMYD/tANL9U/bJl07ubF8yu0jMNQwPsw1+1z4tMn+FBBRvWsgG6Qmju
CAarVwgAoS//R7x8S3AV+6fHIQGJorqA4ygkWlWlXgnQh3w/dPwg+Af92aLLlFCS
LGq3MplKPEoLFzTJoJiiUuU4dxYw1nz4azWvDx23vsQp6DhPZ/wv96+cqbhpjjM8
IInnSgUtNd5KGG9MGoH/q5n69cEnHa+NJUA1Z9ukRi5EWH4LNSGuqNMqRJL8F5wk
EEReuUKQz29eLzn8doJ3leUwe0xz8P4zowrZ+3eyDXUcIWMFD3f65NQ5BREYxDTh
duW/jiRDKtA25YtJmPI1LUgQpAbpZyoFRz0W9bTG92+YxC7pVUQcC4Lfz58bDtFV
zeB2TK3phShWMo6zTVknDffyFQ8+sJeo+JXy9a0A+PloD2t0h+sBzvJo5U4dgAuX
bPf+OrkN0GCfur0rxV3dRqlgA7YLrxysz77DwKhieM01Ssu9/CTUIGNvLOKrFOoG
34h2pR2kVBPdmhKbMe0SRQgraSVXbjt4xsY8ur4DauZQierPrytKQE4LLLcavMvc
YsLE9gCVvEg73iYi1Tk87hTONiwCCv08/4BPDGjkFhdsfIX+uCbrW8XfXYyIbOTP
OoCqRFCYBnDevFeJSaBfk+nVZPY+v56k09v5aizmHb9aKWZYGG+MPGPZMPRWD23P
ZWHl4CZ5taWlIinAikFCq+OwikKKqXvU2yp0W+oav6f1L9ws+S9obIkpiCcF3wg/
Ocfyz6A2zkI0iLdfUD75qK1b5CDJeWZbymucWVNhCWG5xOjGVfsERtgRbACnd1BC
bGfP2OLib3vv3wP8+jHfiVQ609XiCBejiroMz1VxGz7KqIfdnvPxtGtKASSao17Q
8R4QWnmNcb44s77P1MyaiaFMt4EufRIa4tOKL/qPDUk=
`protect END_PROTECTED
