`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9XulBFJYljITc5AJtFS02tjjKUZacZZoSkSTgKXklZ52yvgtojc9HVeeUq6aHtXY
pqmwuSu7g1ZiiLyBn3Ga5xJf5Rg+hqEFlt6gLtfHOmSsUxIYdcOYcAs09oVcgUKr
TLedKOlHdNFYQtl657DkfG5q4j/ndHMRBEu1IWyGvUgsaHvC5PyhlREArNEwevlg
26cPcnXTUaYYQ65zZ/++mhlcrodynA0bmtU3GWIaNXi0WhAXKd7zjeUlZbb3jj4a
D5Q2WG0jl9BzVR8UTmfHCb30JOXwI84z6pfgzm7Q97CqR+c75rhVh8CrrsxxSwff
8FpyxW/4e1l2PftrSK7eUBGubvUQtML3heWVLMrDJpCyVTGeIWCowp/iAQgZ3QJd
p6ETVHzEeIweqDLQxPBjDl7RGSjaHWXS9mVdQzJfPxx7Gyv7aRPj1l5gl1L6euJK
OauSkdoRR/NpBgME12ONNuyVtbVo+NpM7AT8oWuX9A+79owFGdTGYGVgqaZu3TxH
eedVNAa6aAWe61GZyCI1uADZqgvjVfZOMOnS1d80QqWAoHziPcgLsyPZBysjRl3K
1aMorkKOkIME0kwfZBD4CGUD8+MHSHfbSvr0dU1SxM1b5uW38wNuB8JXmLivBoBT
7aB2HhSoHePNpWkfywXAm2PNPycL838QFHrcsyFe9v5Nf7QOsO3NDyBjJh5WFxsg
7wmqjySv+IBnFrM7RLaeOQyvVSHkGCp7tW59nb1p1Sd+Z5ng2noSnH+q3ebEaQmi
EgpV5ibLI4QMBnKbnEzRmIRHN+y/9dskv2llfKT4q/mkjxEZEF4ur9i82DTJI8I2
IAcxTmi9cpWvgnCxzuH1VpKay19mrrAYGk/VWsCJXHKbYg2MDgtcKaQDwjUAAddU
K1S7izcZ9TD5545Mdrk5AdC/LGI0e4410dExz7d6I+ExMcoGao97HweapAxJZrZ8
v0TZRQe7w3iRCuaEZiA2mYsVR130oyMzke9/kLsRhBZwtNzS3aDuGaVFvoYKciYB
nLxurGq+aAZFLfbvtnogLoH6zi76UhP4VjQU2xG7bCrmz4rDgLJPG7LOI67JksDN
Fcf8lyWFGaUJiKXLRe+kGe9ijKLBgszvcafCR4c4gmmDk7n4JQ1jcdEpxP2iXSUh
WHnwIP3PHpgMRXTuLeQkw4H0gFdHYxUedql99kb/vUvW7LGUdR/lUd86SmTjVrEX
iS7DenknEBVISjhQTiG4nQ==
`protect END_PROTECTED
