`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zue89fX/PaS/3COC2RMIiJPzDb/J2vqK4egjWYHy2s926XKJKx5TJ7QjRVU5aMAB
JXycZSirAPbXGTXemg9z5+nk9h02iVRnv0qxSWuVQJGaPwS69NDeJ+ODV7QYKgmr
Fzb6gKaZXKTRVuDvP15eEcV8lEDjkr/ax3msBKrB0Zs4EHPShJxPHl8IgILa8RGz
apzNQJTkyFYtJV0w/2uXCzlx/Mv9e7zheHqTTYiK3ZbjgAojulrCXqsvbi8EUD8E
zBIFdesphxLL2iCqjmEaDrypjg8vln2TiPlkwERv601Z5zJ26wfnE3SDx8N4wVv+
dDLSUHqtuKd0MPPdJ/7b2ea/GopVdkr2knjHI0BtbER4Q9uayQh3l1KhM7vyvDVq
2HVgzHsmbSkUFl8alJmOSnzAyCJV1Cmd2GkZvhxCOrET99+jM/yhkQ2DFYzR92eT
RKVonvyttvaDuKGJEcW23KxejfuMSG9IcuQeNc47KcS4WJYwmfjAy2Una4UvaCqf
r8CsYI+NZWnZKlNrePqm+RzBTPaTPuqTPmse1c3C/sBUpCvRh3VtZf7bIG2WK+02
jlztVZ5k2HtITxRb7z8NBZ6p/idpTyN1OWXu8qSV+RjRPuAHD1O6C/DKHK+UbB6N
YJA0oIvV6C4BQXYqMyN72azF9AmtCbmaAM1t8ycdgXjYyEUDHRwx5iFZwrfv7W/k
V+FqiqSEU3aYtFy/+Xa0Rr3zvu7fc7ee200y6DgzIJlss2NKG/xRrV82Ut2ooASu
veGVqnm1lvg4SvonCfkuwQ==
`protect END_PROTECTED
