`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djYj22QdQ9TAd/OKOJhoM3NgTbPctLQ+ej+pvelB4j1tBREVuiEVnSIrBJPQQmCE
k7e2BUkseGeQxO28nUqW7gPXLnBmjmf1X+Ee6cqef6eRCoeEI7kT0VLRie6kjZ0Y
GbIQf0bbUNY16m1ccVWD39WDRqaPMTXBob9QaOkeTC/ZmBg3Tx7Q8wiEfqWGPb7y
lsVsifDkhI1FPfdEFsHoaM8qcwkiEOpTxQlSERpJ3oNUVkB54iqum9rdg55rMETn
Ru0qLEZDvxb0tvI5P4aEjcHQBb9Gvp4WqpxBoDYRMwY7t/2dgWFfIm085dkIj4Pk
4ZX8/PS5vIZN+9MlYA4YrigQbUNkSDX961+bQW47XQoPTS5a+MmO0j7WCwL52LRS
pr+6IC7ut0TwRlZoq/PdxzfrC1cosnq+M83s5kXn81mnkd4LZhxonfprx+H8O42W
bO+yyDbCg5H61DRl/WohH/eoHPoW18L4CRsbMz6wpzhqmi6Xa7UrMcDwTRYgJhMT
bndefmNVElX2wRo3Ifl6qwjmEPG99o0xkjNqJtt5+uJ6ykjUKzJzKCJicmsFPj2Y
GLlMMHpp8YMQ3wUoN1CEEed7oRYgIedqSd5rVDYIY5ZgeQkXYsLe+8AbhAEBheQo
O91FbAI4b2gq74WV31YLTvlG/RLMJ77NOBrVAxaMH+pVrT0jJ/Dh/RvWjjm8HJrk
1goghh+2VFojg938mjZqjeRMfx8KDkW1WDIhWlqSnsc=
`protect END_PROTECTED
