`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
johX9JoxVaE5zHBvzzGilNZHdqa/lD0ZqMG1jg8/iHvqVtiMsDTOla/P/kvrt0uM
qaI/y5kg2pCVaG35MlphxpoIua7jnIi9gKJHM8F6WDLyGWxX83NOwHVhR4y4Nrai
cHlQMrCmpBF0O5HTrQpq/fCVTFLytF+qReO9WdJEs1yP5v05+2aeLR1PY14iHzOz
TqYTUw6pzv1AmoTsMs6Q4yzdT+nfP5Rp1/ezc4TPq0v0te01Mu+8Ip37WswF0rEh
TAv7iI7xzfY+5SN3bcIC1Jbf+vFmABKEp3d5M177yyO22bU4r+1/Ov1vvB1wW40N
3LJLPPW0cwUO8+9RNxNnrLO6aSW+Ffoz3Z2OK084cGYktyo52f2ZEm4pO8GF0IBK
Qp4TH6/VZ3HyikrYkZ1PB9rgSvXxWDG/WqBGoctn3rNhMSt0/ZDtD0z1UZJshCQd
AVYf7axXO1EC4IpZm+2CVCJ5mCwx6IFySCBVGr0IydhesLB4jWjBTuzeScubsyyQ
`protect END_PROTECTED
