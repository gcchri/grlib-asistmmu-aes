`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJ0sYC9lj2GAaxvLfSHBnD7QeQUJ2IWkWjm5Rrer8pOvUoI9omOoQNoxayIDSU+1
TvbNt8UrNJGwcsr8pZ8AzMkafNgqjpb5EXkx3gZebCg0O/JZodZVwJvPMi6/06NM
KKU6arYk0pQJqD/m6FzcpXlHPdBp29Up9hREmHqaoEeM2MEeXPklGACFM/t6K4I1
Y5xpULCtjpvf4Y9320Y69pALzrrl5XrwcWubNsWp0B/uLnN2c7wDAjb9c6oBcSx6
9p6HIjXWy3cSAffuTIxgtJvELdqY+o+FALx3WSugoiH7mkCLUDsTHrp5PhhY+a0G
hVxwsjqbWrnE1WlUR6ZR1hNENWiu8/w9W4rtVqK8xXrp/Eey1FJPDrTAU2cXdXIE
O+lkk4ZEX2K59utUvl8UtPU1UpQIKk+5w5eltCjiR3dH8LTLzMW5K2oXamBNUCEI
Ao4Wwgix7MEzt9lmBYyw0ReYXLjEZhmNt2VsC8j7tFgZaSdHXDn4/75o0UMZ3Ecl
yQNuNNGhaQomPN2rZdBPORaIaQmoab9pF8+wm8WSTmCcQ5CMCbB22fwzWWb3iGE0
EwZRwiFwAhr6sIy/2mIgpd89qmB9AWPVdWDLhOL4UmecfSMYOgPdZbkH+bXwaalX
GmnJIAFIEKqlYEloX3IpDRu5B5H85GPRdADWdTC+d0ntqHadMjY33WBWVj3VU0U5
rvnIMHOwbjaROezEwN9wcf9++fAuhH2XQSV5ueEU7mrIlJOZbrpgr4TeTpRfB/Mw
MMVk1cpHvufaViQVN8Og0YhauHRHgTDDjuTTjbbxCV5Vw/pSMbkY0U+vZzrld9pk
ehctv7b6x3WVdRdt3P2cZ9jMoRHyz+oySWgdK+ZJ8GlqNZ/Avy4YP5B2siDf3tAr
mkwznMpImW2aLzoKBjryq6XU9fFtVD8g+uIdnoFQeSLzNMm3AbM7EDmRG3RRfZ3o
gXvGWabEFJgOjcC8V8s5dwWOa48rF140IxKnC3LNOVT9SR/SWwrzBHCffBdDeN0I
2YESv0uz+dSVUKfNJKjZWjAkM7G7pwu8Eajmhtv1SpEdpbGH22PYbMV16ZLrGRRu
5LYamM/uFNCt9knr8UjFT/dq0B2UC8jU+cT3+PhXCaR5I/SokViPuMoUbk9h9aXQ
+2IKaWf5IL3oyVeLf32EZQJPULEorMt7uPtcAUaZ3Jp7JKDPPuseEanoFd/RzOKv
RqoOW+W4O1kliFD5VX45jAB3ksKabH8sSdMitJG+XfM+FchLfkuDFntqlhZs1pRW
SJJZ6uaJZy8Jv4/g4Ha+hxvSrqxVudaTC2YdRZ+JPyLkzzNTzYBbwZDIveYxpM9H
LxnYVqMZWb93mi0J6kUVgwt4aCkTPT7Wz05KeCWZnAs6ztipglSXLWEOOeec086M
uck3ZfNjjEnpd80VJ+vevO+znXDmNp5H2/5Mk+7U1jJq0rHRMgriQ6kBdg9WLfQk
PF2qofbFUB241tB7bD1AUbSmz3qkK8AVMqFpnQG+TmMbkXEHkQq+Ef5ClxnL39n+
cv3zZzVUCe2oJTdUYSr0vAoeFS/SXsqIw+9VODEKzrGDwIN8LFv7CX/YZXiszE2e
7os2eig3JpCDnLFabXpgC76Fi/j0jBGm3vq+ylSA+acfkRPfoOh9171W9E4bEIwp
GPxCdtUMn6t2tQJaT/762210keQPqflcnaaDU3Pekyc7RHmTRWGVvPzqRQ3OK6S8
gsej8l7NRBOZVUlWWDhswVgpQLN4ge3Iwq/9I2gHVQ7ugdTkKwqsZJv5WspwCV4x
ss+e1reTQObeFSrZ9ArcrsNMUPeVH2DAhII9O5Ketjr/CP41U1uOgJjDvMq4HHKr
4YjpRji6/zXUBQGMugaKlErxUkHa/kRMDVpVlKoG6iZwtO4shjmHk9Idw7cy8em5
6WJloNlkXMa8YjVV7pa+k85/1bWJIFCc3l5xWsiMgqsHS5tCdunkIazHqk8+IyNi
vzZtkEzyzzblwpFzufHcRvrosKRh+y4wm6ZDsXyQLSr/UQlDybfYc6egQDvUPv4F
gGnIJiCuWOl/z37ROQsNrBETFMPy+dLhpP7XB9qrZtJwx/X/1Ec8cgHcKYQ1yCGb
o84KHQUu0VYQHnjokqigJ9Fvt/3vylQ17i7p9MV9HavEK/4djsvIVEjTbDRNAd7g
oS8xyapcFypnLCv7BQBE7lY873CqgVHlpU0j7TFDVh3zTXOF+4Xloezifunkwhgh
DWQyg84jwKLtFbUBndKewg==
`protect END_PROTECTED
