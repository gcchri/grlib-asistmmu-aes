`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cAKdkJ5I5g8JAmYhg29IXuOHhmmMJ0iAXfEf4fnxPKa9FjtJyvxQ09QT8gN0E9g/
YC1rH/ZyoGWYtq1eZmjAfubr5AIxvcGR/nYUHtnQqi6++ZXjWa06M1qqd4KLWm6W
aaD8Hp6mhvNqaDQmQ+Z1eoLPVNLWeyBH5DSq1B5QxsQlQ8Chi1P3yoPxSC3gd+6M
eGjv8rHClIUx9OrcHBBz9UuGb5Rd+7bA6WNsYetT6Q7GNgU0UtGKUduwkfojtDpx
5JSKwM/fq1iUiboB47Gnq6aiXCbtCxrcZTfu1lYzt3+50WemVusf+F1hqhQBuwEi
2yEazIpiWQS2JlPrGJMwqv78jb6yV0FT1dpuxL405pKBFTpSZB/sSIw0xH6PEAIx
lGdLJlqDZ+fhADg1haZrBg==
`protect END_PROTECTED
