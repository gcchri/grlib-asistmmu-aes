`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m09grZMp23rEt63ag9r5JNw1KF1pXQq7OohlgaXtpFRt1GDOXqF1ru96Xv7SlXSs
DT0EolsU4CJz7osBZlMerfsopWi+gt1ok4HD2UrYh3eAcygooRYm3NsrtiuW8oO0
J9TEXXl91IvFIaqjXOSdkym+lTAwtaZCe2MtB4rj1FtCXKsRw8erNF2nGoPoPj1y
vunUUxpznjsBH/ekH4JQU5Htw5ua2tYmI7OUQW3e0rxzEmZJlO9sR2hchJgeqHdC
d3BylQdFHW+lqXTGBKKVovYtgxEcb9UwZ2faJW19BdsgoJjjGYBp7+GPmI63MNyU
XSY8JcbzevCXei4aETcj2ptPzq95IqY9ppqR+SSSHy+Iv7V7lkFLqoi88w4ZnT30
Hv/Q2GQIoyEOthOJ8BqTh3ROOmMo6MDfxrpF3yQDwcv+fQSxDwaaLwAdVZMG6Rrq
4VRK4qV3texlbzvtOa8tJGOeC2md5ZJ5MRG1JnU5MJs=
`protect END_PROTECTED
