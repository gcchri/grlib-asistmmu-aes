`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fsrUawhqNco28ij244I+w0FZHGw+h7j8M7rM5fLtO6l3UbzMTXi8RSbP6ogRmDSw
vSrEEegakhJoc8Upg3YaEId9F/+qsH+tsQK+U6HTuT5uacocOT+85h5sIBbHwoXp
D7S+W8ArShd2dgP5ej1GV23nX6cgS1qz3L/V4JiIjWTe6hDA7lnPF9r/uPv+FxIV
JdrJGwikiEIEsWCnjJw2b20wM47zC2BepHHYs7uUIppVzfkqrCTN8bNikSEVcL2A
IhTBAW2DKYemooCAE5eI2ZYdj9ZZHKdvekmDnVP21d0XG4A+x13dYyyPewgtwbSf
RJ6pvzpGvTO2mVcOF7cwRwEEAPUlGnm8eV8wp+E6V9kn+haCZmaZkfKwsAKeI43M
3MK+r7zu9rubub7rZnrGVzVLninRhEh5SrTOdQ1mz2o=
`protect END_PROTECTED
