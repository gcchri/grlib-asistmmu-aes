`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jom8A4+QabxUy9ejIMhh0qyvMIejEYiTpkobW+R1PDnqW2imIR7OMnO+HXOuqeW
Y8sWUHWVx1ln7ujRVxrtzK7h8CjW+8h9CVQp6oarb2m7l2CUGexeDRX0Bf1Z6QAd
OvYsiMUcaK9ko+KD4+pe7+5IE0Bt3bqAfv47TYohG34MEcasZrmcpALJlIZjX1lw
ylXEkW0jHdo7RKLEECFi99lkKxRgIvz6eA5M7sKejwwy2cHC9L72zasXdC8ljYQY
`protect END_PROTECTED
