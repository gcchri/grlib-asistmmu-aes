`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Wo0PTsKt3KxTWjY2TQDzKqI0yetQzGOKnrwkmXHYMdPnbIWIOAKzT1bg2XC9c6T
awOB24znwNYEAHkJpHfoECGLSBZGJQ0Or8MVpaZ+9IrxP4+21spZLWFZk+kXN2rS
mOyGNKInQge9Jf4Vf9cUcpuXBEOc+NPxnIPjT2uZRaegzEWFBAvw75+xOpevmbab
oPSRL5SL+xOh9qAzSy5tBdh1u/zfjvCRKVOEDxoFdw4XN/LHahnSbw6SdoxMe1Pc
fP6ZEwyqlo6JauSrAHb2eqXBVLxfMh/0MtuQgF2c4KiY3qMHrZnZ4jV/DB+51fcb
KX62I5s1u/9/Q2MjbZC8PLWaX0+ss/K6NWbZwEMlOq3CwjFPGMwPjFTqmIA690+T
SpswDAIawOJLynrOgcYlaJLapAGpQlwqWl8Ddu4Ap5Vkoy4Q67PgWvrs/vhrzFTU
I0l/7/NzqNWRNoj0RCRpYYldL7qzm5vUPLR4pm+y9PRyhFIqdxLXLRGrerDJBu55
`protect END_PROTECTED
