`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
usfkmWlVdVofO0RJnbnl6gJUkywe+mgjcOm/tFiBLDSWyJRGeUN8OVB9jGqIPY5l
Xiwo6Szxo9J2hiy93wb6rEl+Myj2yEvzSb6FS+2OpA2ITfhYvaZ86R4CenBmlXnE
SgWfeXeFTtexIIfFSeMtsDawhRzfq9X6nopyTP+cnX7dbfg2+z0NBLjRdnVdYLuU
9XfzUdszk3UOwZ8b5e1GPu6VU9J562iWCGr3vOaZEtYOzDlX+drrg4KhuWvTlVke
QCt5kUEQiku4JzLTQ86XCM9IWZ8N8MwYCFoMZbey0ZdqVdBFxtFlGJsHq5As/fY8
cvqewryMqop1A2h3EhakLtnwfu8dPua3lQtoY38xg7vOkw9hhtYjXeNBu8xRXL0r
tdfO+wuP9LWuKGciBSoP8Q==
`protect END_PROTECTED
