`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMlzQJDuThTC2SY5uQYDTYEMVTfacEhQTzEdmJG25tibeELauGARKU6o5LN8egfN
9XNb/dMDIgIvpRu9h3l3crMYKijn04inRyr/awlAFEPf2TSR0EXbJt3l6+3uHW8Y
RMI18gExS6IYwzHrKE62DXj96tglf6duPsHwGdodaK3VY/1Aup+0vFzK8X6h3IKg
OlTgtnFESgT8ABOVrwkn2EhLMz+RAhjOcmtgYd6A4QeEcw2FSHzxESAk+Fpe301p
J+4PBPIj+skO1ioKFocmubr/i+qZQR4/ubrGuAqF6+HJnX9txacMO94WMabqqWp6
o8oYcaAKk/Ig2RAG2wyOWrh9NyLcUkRRKieyP0DByJDWWy29V5vHNDWYEPJpbMUc
`protect END_PROTECTED
