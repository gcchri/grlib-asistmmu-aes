`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qm9eUWjEU8AyKc05r/HYTYXuulAX7eOh/wvmfsaTVRbzs4SyItrtmLOn0gqw7iIO
cf0F3KG8E4oBIPkFEaCUkcKzp24AkynbLIE8sFFF8PpQorlMhlh7zC/OdzC3D/7G
RJAqVRGNXX2Ygc3ohCBjbk2/hgzQTH65V9DOk0YAG4Jb7HtGNm3KUCzd9arrC4Wu
GgqwrFlIt2w/+KhZSlnQ3QNT0EzTqrMmGxfYFBBwzLWP23lJFG/RntxPj+BQwUcX
mG/ufodzvng3Ebto/GaWV5pnIQZvbrId/AfL8fOAbxteOfjmd+8CJeqMYNkd6P3I
5vyn9zQDcqlfIijvMZNitXCUZQ340rK++C4QepCC/KObwYHRgM90Y3H4wwDBOcXk
OOA0ausr1xC1ATJIQlck+QpF579MtlB3jXJ8FvwmrEs6rmZexub1bw582buXnt1e
pjK9/uWIpBQIZyWt5y9FM/DlBzcDa2MD20aFenwhPEQ=
`protect END_PROTECTED
