`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Vhi2i8IbIdDbgsPP/f7BWjxVBynVe6MLsdU0oUKN6PpVsDeIZfV634KOcECZca4
U7d4BpozS8Zl0RfLKg2I4JVCB7a7vXCoWbXj7ef7477LJLExT+iqQEYTgLYXr1Ac
D86FswwFSYhJ5HBDq6I433voC11dI+iwd8yRDu3vz/tXyBpBY141QSPHlg0dSOO4
pOg+Y04gagC224xEa3Dv0QkysIjuyu4EY2fbAN+ZXrchHLh8PwsUJ6FtbH+7wSJP
N1M2R1vIW/gBEDq+JcPyeEYVW4s9ajwBfyLmYNDtbjhecnUpEbZmjcuSXveYShVZ
ZIJgknMkFsME59HmFEOPeKvJiRjMo86VTvsU0CbxVSkGjmUV1BT7LD4Fl57s3Z9T
vmaiOadjElXskMFRZb2yhCh23etQE22HdSJtmpKYuwQ=
`protect END_PROTECTED
