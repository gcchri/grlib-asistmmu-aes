`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oFTz7v7NtOf52OF8DIOK9cjKn6X4e8K6j6z9s07tp1WGw4fcqe731mZZPoV4Z0dr
ATgaQYEuGTlKhrH1tkQegFt9ZTWqn00yG9pnEZDVnlU4keREjehXH/hIJspa+wec
Um/bWX+s8VLl+jyeUJXxZB0WdLfZsroVndGqOJ7X2Js+HRuHUngWjjiMTxWX1RDm
x1EUORBnjzpyJ0rMJbwxCsIM2/k0uM2lCLs9APPVfA0jxUSssKR9VTf00FmwVBuw
vabS5u3HX2mEa6FO5qkXJiNhBrm1suITfAZMfsCcAWx5ndJy62NVvWslFU63o7p7
VjsWyRGwJBB4XY3HPHzPbw==
`protect END_PROTECTED
