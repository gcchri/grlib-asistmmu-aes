`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LAnC62r5b3oote1rMvH4UMrpAoBwb5kYhLDquypIlPLLKYs/5Reo+09xLYKzB7Q0
OCU4cL5JPs4Khw3sy0pI3WDqinvoSLQ85KuSHOfC/8AOs0ws1SJ/3y9zT32mGgx1
zoM1hBgkfVSn/7Gtcz1Ld/PVwPzBKjMR7Mn7ygvR9Ofy+YU7gsFd77yUSitwRlPs
HGvwBlyYqaSfeQppgJseHT1MHblDV8aqwkyqJ17xWgtC7tuiO+W/TJdsAVZOAgYR
1Z0PTaPX43Xg+7FivZEXywoWhrN3Bl/tRdGxDyajl/4tbOGm4KnpVTXlV3vTYP6m
NALJoqtBuQaRjpQrGsYD3nF4hpZH18i5cEaL7xP36b+jP4f+Px58Vi4Zc1nAEpmy
9YpeAuCJSw1J/CZle1fKm0fPNGmpKT6VYB0jq+rqKQg=
`protect END_PROTECTED
