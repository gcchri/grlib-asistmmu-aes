`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HYMZ64gUKc2bh3/sUJl/luN2uVwavZw4dQZuDb1ww0w7ruu7YTyIriVL1jrnp4Wn
Y4+MxMEwSHPoYsYbiWoFNE1CuVEjb9WaQbJiA0cxYIavgvVzY8OFYhuDFBH3TBj9
y7Zp1NPPKKc5UBCMUfWtTI1U3h+KKJdRwk1JCxYOEi8s2s/yc6QjepiKvaexO8XS
tKNqVr2AwF6MhsbkDhW7TKdUFs/Y5V0x5CTtFIF7f4JyT5EOvwsJMvTI+CJ3OPz9
xc11mMb49pGOXG8vnEWTHhxJ/qIdAWpM5MBQ3IwWGEhfHACAus92+DPNNF1v3VG1
Ahc7zUDkNUZ2XEx7Ta2BhHOR8MyotPX3CcP+FjvkVPJLCA7zuxM8C8bEPvBsX8Oq
rclirBTH/ohCsSjxDAsmu0SE0XntwzvJBp5zp43UDUKiNXg3Ii56jLGi84U/DDVy
z0o44qA4V4quwOrosYvOQ9RoqN8wUlPNkZOVHae7JdoTetNZI7474rpViP5dekrC
f4ZaR55ylTTXnUxRWIywOJMZ23e7tdY9Sfd2jBcMoNPk4RgJ7fNaF6NAFbLU1Jt9
yxCyXbw88htzyamDkemncx5D0sxuuGiMccOUsyELbFMqYB2eiKBlV05SikiRq8lC
7cBulXwsAdu0qfP+//gTU+CcMbc8LsnTIfY5GjybzDK8vwlN90MnASgX52gS/Dl0
wSCwV0+SDZImqNYXSwwQIM5oHlZkLTKgq87uiS3jRxc2e2T50+dGL8+Ey3XQaAd6
n62/C2HC4FNYh6puoNShbe5eNaPtic5gcBe/1f8Z5vHkjOgax89WZW0WyZOSO+Lm
tS1btwP7tb1Glnfwe2ajGXSpEMAQ3gzldmcDdwTfIT5LEjlEL54T4Z7UYwwRilKc
UrUKoKUMknWWVkRYFxzJ4qjEqhkVWBl5KSD/8CG2N0FE8SVTake1H/MbF/f8RJ5H
5mQzAj0rjQsPG5E+Q74I/dSFWXeml/n1zoT95d+kiJsvJOn3hyfNzCpU0wZydd7O
hr6qQGP4G38iCJLo4JpIzOvRKnc0T6/ec7yzG8BWB33S9ZYkT1dKxHsFoLQSXEov
EAPLdjGQ6GebFcNlVpx5q6zlUAZ7f5p9/V0bCbXYDivhX+1pBBkFkIA9BA5lMPco
rPmlC7YVY2Y2bv2zn/u2KIVxBzvzX6RTSgWS96O74hbQOH5E6+tGpTQpbUaxlkEa
N0vnRfM/6dVdwDeKmgn4tcfSd9bkDDNH5Ac+w80vbP8mezxP9v6Vjv1GzgfEcXnT
vso7zNIXhGcnUmZrWa1+BBClIVprpUcqFkcW0b9cDNDYUydIUUYUP38CubMQq+0I
YZCYpnpgUiKPrhtVi+4QzFAn2U0Rl+0fVHdDt5oLpukjUxJzsA0oxNEhIBjB+PkJ
8SJJCAMjF1WzdSJeV10LIxEfw31q7aHlc2oiW7IXFt58omlyovrg1ufFSYTEM0fR
6rDXy5FUn2ovlhkelw9YYQ9txKkFVE5X/cXuo48VS1Lqm8gsTeD78Z5vPcPU1XAj
YCJX9XxzoG6CYaOq0r2OuE7Q+gc3Vx/sPbOf6TTq6kuflfgvP/KopwdEcStRKHJU
Rxh57NhZWCdQjowH0inceZiNeEWzE37HIVY2I/ksbtVwnC+Wbaa/bhe15ol3DlgM
TQT3AoKWo85WtsFzfy8SsTTCXBYk7Nrq55W/cWBnKxTK1znlGmpaYKvOnjSMmJNF
MJCihfTg6q0djDPq7StqVbZbt/uwSKYY6yia5S0X7oPqC4v5Ds40FAHzJjM10Lp3
dxFTZ8aex/JmEzh6NQOEnnQmeV4sD16CClQzouewfATfML4nA7PIi6qM9Ik2baoP
cxpf3yK9/bLXS4B5DyUPGiDJ1r5yV60P0MDic/i31/7VS2y7r9VGwpmn7pAQJdqT
elXuySmhWVQSSvpDBnzPm3ONa5jbOzqzf+uHS8/lE7qCZVQXDb+Mv8jBO/AS5zvu
324nnkan9YpPNSTgvtW6HQ==
`protect END_PROTECTED
