`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ssfw4CXWdEh48UyzHQ5LJ8DiRhKoKrBfsmB0OdE2Afaa3VmjzR8CSffzpNIk6ToG
qSF3xy+giQl/Le+60+SYm0gRfp6c9aceD2x0www1by83b8hmmINujZJlSh03Q+Zd
n2LkFMhMQpHcfPXSADP2UejXbq4AmgDOg51ofgfxKkjd77mQQtLDdre5mSA6SK5D
6N5IgU0c+mehVtL6qMZRH/k4n2XZNmzWCQ4l1zyd+Cw5eji+FEUwdphWgUv3IuS8
MzyvlHSAaGITy5VNmM3v/1dR3iyDmTgqc34oQ0Rak/aMXvAXIq0rCuesAtZylrSA
pa3u9kRBZ70zcJRiS7Cd5lpILUKz/sIYqRW1pb504Ajz6qCpr3Vb3ZBXp26WQtbW
mln/DtdP6rX+FdePvV4kT+nP9WB9Gb75JiRYKHPgfdWBYCKHcjVX5twQZjGhU4Um
G3roXyY4Mvn2RtEYzG3/7SzNSQ5bB/xezrM4HHMO7TkY7SXxCv/7p2m1jbJTb3qZ
lGbyLmyGu9is27em6jqyzrgj56sLZacSFK1tYPD2oTO6x+VT32U6Cc/CynWChzim
NCzHjne+F79iXqbTLSunqqJ2tlleHmxyoPmI2fqIUMm+TnIxegfk7Gq21vo7N9np
I7i/apSiy8Vo7pxS2b9y1Q41+Rkl3CG1YienbHVAySQWidfqCQD/KVf4/OP3jNHh
5D3+xfQZ8fCiaxBnzHvg7JCBgvYWZvuKPBTUAEJFjO8=
`protect END_PROTECTED
