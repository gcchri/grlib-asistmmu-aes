`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICgivQ5F2Nv/RTIqHnEv8+RtJCoeGxWwVd6hU0VgxObLNh9mm4GxdzrdcREdErMV
E7UUzfIYhuu+8++pgUapcU3hGi09+KoHfOtWbsDj9JApAOQHAuWaa0xzXDmIV84G
1sE9OlkvcT5Vtpc2Hk9qsfhribyZT+PgnLFOxSMnEtvk4/N/Bra4Q0wwEGhPVdCa
ojy+FHSAk/EJseHOL4Yc0Ir1IuPOg4GF1DS3N6yk4holF+3mqPUlIjjO1y3X1R5v
bTRtVZ4SW1jQA15mSJlCLIt0El05LJ+YnJYt+NtrFzcmNghjuxANS6C4blR5RqKj
Ntbe1sPuyWewcQDKvW/hKw==
`protect END_PROTECTED
