`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N7jlRduYu5cF714FdsuPU2v/nYOlrhxVIh4CzL7yBD3QQeTH3LDaYjjWsJQxqRHS
vkrD5K3EV4vKBgVV9Mfo6MmTngvk7rkJDiRWlxZUBBzLyVTbeTfu7qdmoBFckOSg
6vvwDLfrM06xBxT8ksTchBMBlIUZOTwPc1NuXx2ri/Lbu9crcPfX53IzIkFiG5R8
DIzJiosPdTrDyxfnw0jk0ElukP5ZeXhVu9d6QofQLNL7Dv/FPTD1Ltikf9U+c6H9
JZ7C200vio067o0U10XgV24B0uyXPkuuHkt6wgwzZTA/vNmfg6KDU+j7EM76APeR
`protect END_PROTECTED
