`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uKZYH8UZ7gIvOpVMoYwrRBHLqInTkedRskDUVKVrRnHwrt0+kuKcXc84wX65PS7m
jV6P4EA48TlRIFDu7l4+8BWKNk3BnmI7C6s8/Y1FYQ6Vo/RfzYIFmuc9QeXeU+ee
LD1R9UdLXngINhUZTJS+SWnA0B3vD7NhNvN0KnnF2IK7zryeEv8atmevYwMrGKcw
Q16X6g9KLkQG1PqZTCM49Y6ySheR86yWkxIQJLxD8YE/fhZ6eQmrCy+X/SZvtA06
vpJlnnWJ/NSt87kH8YzfcoeCoADNyA8vTueXcwaODf4ibhoYwZ+/TlgnxQ+Q8FAM
glRN1zaO+3bXDMmvySQ+6gZA26guhNxgnUBzHnw9hJNrr30VffEQHy+tKmSumIs4
k/BCaDzpf2p4JdjRHktT1XdiDGlM07/o72t1WDXV6Eoh7e+y8tc0J42Qz8qQIigL
5pDsCmN/z7l2yvaWZfQslHEV4fEjiqWXIPhZvsgjhCn2Xt5zO6JbPgIkZcKTyOVf
NeZf1WK/Y01+eFVtDCXyOOiyQZk0xwHaDlnwxSggOZI/qR+kZVtIU9HMecK/bdwy
rCvErsiVLQDPE+Sp9Ej8OXDqt6qIqKtfcPwg+Qg0TGPMWIA1MSXk8qbQF6X2MZQN
mc5/VX2r2vRrFu47il++FheyyE2XABLc4OWr7mp6j/g9bBkL5U7f03sfeAss8JgC
YDyA7EESjMzkez4r9Fm352/NPoGgT80Ao4Z0FBLQCzGThZ7AgRBKpO7iYD+JAlsY
wvwq4kQB84dKJS2ZWOzKXQE+e2UwDpRiUUf4RWaDVP6MXHc31ytutOnNOmVXXDiW
V4687peLCNlNItLJaA3uZ5XTEYWG2U0aCsmLz7o+cjjezc9JDbbt/syf9aQeLWG7
XvkOr1Fj+b+vJ6H6U6yifrgBk4fjQ8PUMEVFL/CWyjU0vz73RKZhzA8qAtiQhtXA
El+yvAMFPaks2XXWhkaq6aLG/RIInaiiSvio155Xab1bOwCfmecvP+3TcWDTGhym
22icWyo6AgJJhQC0g8WbMqIkTJu9NXxSmKwQCD7M6NXvafmETkk6FK9tmsyr1UAf
7ybnLgNDCKj4zO7kLTyGgIhp6H2DHFH1qO40wWnwLyUVv5X2Ck9WBQWMuO+06ReC
OU87acNLeCSjEHZFlrnT5brupuKBmTOT+FMtOZDyU8lHNZsMdGYiEDYB5UcjArI3
6vPiQsXztQOHBu9x9urTwQjriI110MRJhcVOD/puxeMIR+DlPFb0EWn9eIptuUw+
RzgNUEum1zGxKw1wD1RXAIujfVV6kRHS+326h3fLHhET2qVzP2wAjdoHmF3GRx8T
AbtKPJ356WHuvM+s96DlJhvLPtMKQ8hpKoQ1gQxA1detjzRVe6K9Qe7v3ttaH3AL
a+QrY1FyWt5DlrWZenjYh8DkMplIc2mcP6fnM71EBdfgRp5H50lqTpgFeOnnn8sV
O/0acfN96tU89CPL5qNTVpflsyqxa7CCaW8ksU++9FRv/mNLX8j7ipBHzKvV8tGD
3ritLg1Tj88uIzcNh5PH5mbw6JAvfYF9hYTDNgbS4lRQ7xeXQ36niWEp/LSnmqm3
wTTs5R3YwUvZromu0XvFhuunx53ya3Yffb35pL9WAKJDhgma0Ah0SqTs4WLH8Ef6
46VyinlTTrvQHawhuY+EK9X0YVzb8pr+TScEK4svr9guVCu1HZiCUc7kYCZ4pv5m
RJcllEdFjCuTHhQx08hvIZJt7MqBOEd2uNO2Nk5y/R60sYOO7eXh7ysN8GjERfR/
53E0NRYIgnsqJJrHpbp5FNQBvycpshEgs4nZC2e4EQg6vzLI/+Mr4wIUl1I3Gh7i
MJK/OofmSQDtbcnw6jRCjXgU0Pbx70QmMUMmqffGMR6Ke5ELFTPjZIOxs5ejOteP
YVNp4hR8t4hgNE+pvyKh3ToSz1iSXZ//MUE2+zVHfGxHZIYWdE/IMKnteZUr2OaK
E6vPqd9/bpmzR7BxtFVzev+D/GFESasADKopdqCEgn565H2v5YSONhRRnsoKkSCk
UBny6S1aa1r8akARCThRJKocP8pTDoWzYt/P+JFXfrQR6m90eZb6MnVLDDCF1Iow
T+GzoUO5r2c00L9oatypmYFZg/hDBJI6jZvx7ASuGHmQxPRk9gVMzOd2jxWr2TYg
g9L/7F91rrVT6u7tVd47XAzfbUx5DBKwelvgDPYdOLFp4RVHhivscPAKaE+2ZDl6
v/YtIN4CpvY6dmoXI6GC1WEWAJlvuk77DkW/h7Lyy7C2H+kI4vL1j3rGEvDu1j/6
MmtwndbBRXnw7tEkv8tcKpBPa5qdJtzGFEfXkZSrtyuOel5t2i6cQuoP/+/SpOTE
KHvriTNA92PmE3u2QoH3SLoWoL75GE9HJzB0l1r72FXkk2aJf7+yzNkv/Q18+GWk
pawB/pEKkspfHn1E5fW2Ko6DbJM44HKI3w87go10rXXq9Ny7uqQywonYFNviyKIv
BnkLraSX59JZOclwrEO9BQ==
`protect END_PROTECTED
