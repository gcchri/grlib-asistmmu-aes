`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BII7p1VFrhdIXpjnh6WdySHz+L+NNFzsmFV/44t1J1vs63ml16RkmMB/zJWQ/Dlb
P+tI/FqMz2UhS3UfJgspCgmH8IbTtDhfUbwmVf0SjX5PhsIq85KUOnTDfdYHjgIN
/KtLM1Nf0yIqIfMMHKQN0Q9mnlFHdKsZxre/D/yzgi4/TPbCYhHxwljb39JcRExJ
2ZRL83pP9Q8B/hCZo/3B4O4El6C6I+i728yrphOSeRpF9JPqvHanH1ROoIFu3TZ8
3+isXFFVrVfSgvjKlA5fb2epgCncxH1wXG9jEnSFNbRuoBnT5P+VRuXPxZ/ZmWpp
GRHxEvDF6UcwXqwzVHEZmJTR/klSatlrGb4JHi25Kafd4VEtNp62bzlGbEK/R4gM
bYsT3PPi5XZ1hqvDrCtBCmgSZgWbbzEVlt0s5BS+OF6kmmUUfPzow13s7FGOgAIz
K8Zj1WGTsgXYHWMaVe2nq9fwrl4M86Hw9Il6+vUOw2fXTgqkiJAsxpjmsZndgzLf
cqejc7qRszQGAmhXi0VT9SNp2dEMc6BIlVNzWKPWhWAgvPVTHXl2S1bh/y8aeSk9
Ah/UpgbbveZrB5whDcWmc1q+G6iY9p8+gNFnsS642IDQpVQzAbeKjz74thd90c0m
QsTBt2f+ODZ1VLzSkwYUjSSuz6EhDc2ObvRVv9AZNkw1fORjW+XsOhxRCa06ebXN
HKOWTIw7ZqQVciiV4PDiAv31Qspye698Ppcy9tct38PsA4SaANdqsWkZoFkvU0j3
s1XhrdDmtCbC2o1uGngdoQ==
`protect END_PROTECTED
