`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yFY0OhXz0R6rNoTMN8RAc/Qr+wKN2Sl3eybu+Sfgmgja3vCB5Yi3P8at/323ROIN
+Wj8wRfDfsLDdKG6L0KKaxYoXGjspYEgOf5uoZHscvDPXXQYFvTqhz7sdKbqHQBA
/VLDza9kHNqlK/W23i+H28riG6iTeEJFmM0DguZCMYzzlInzEE7KwTwWICwGNfUV
2+b9VXd63xYF3Dw2+NGiDnBsCZzDC4tUUkSVj1nvi/REkaMxPeVic2JC+FbNWsAV
eTZxWVJwcPu7eyjt6a47vccr2vSmobS2okGNPm580ph37E/3TciQLAQlXxOvFaat
eJ3D+tX39LVzeqbhECNXlATjPZKwP1NoUiC24KJmgDvj80Ikm/N4BmBac2q6WCmn
Iz07uOo0Y3j2OI0hXM0q/OGBaJhdVHIlpeL8WcVXv/o=
`protect END_PROTECTED
