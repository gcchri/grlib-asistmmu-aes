`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/VAm2R8jO+LPmd7m0sVYrqQkHEy3VdGpkoxu5ut+RnWeGI32uH0jnsfc8baJxlX8
0sGny6WrJgB7HBZ1iABAWPvDGSLT2tSG9G12Xebrcky33SEJU6xp7CniHpxBdbLX
39FJQ5w73ZvvAZrhxhQzJJcgTs81awG05TSza/0+1ZUbRKRFydW2VheLyIkKZYs+
jIxRgxfuKKQwDSUccswzOlSqiFDDrtQnEpzXwImme7Vf4HwstEtBpZIvs+uItU7o
6lPcFdLuWT1XR7cUoJXtDCQU3bnIZ60gvy+zvak9HyVrEBhWalkxh8L8d4IrlgJz
uCSNFNf6hh5anCx+UMGcRYsBvuE7Ho9hyfsEE0rsa8mqZrcntB8AMPjPvN7XiOMo
GDzlEz5wawB2q9+Njc6cKBHzUXYQH+L10xTw9Cc/hNXGN3ZyMwodITmbjGm4yrZ7
+heLFbfSOQit3cTsx9YxC/y5jnFBrOHoGz63At6egjbx+iFkF6hSV3OriLKSRt3T
VKAE0OmkAEPa25DBQPADkCg9aZAcXqeoiyqZTzedyZOq9zqDC8nkFrhCDwqFQQhp
FZViuedIg3LRQNctrFsi/JmhcHZ/YlbGbf2TqiRHg2kLRDfZGUB90j0Oi4MuK351
VqFzH44py08jT3S5/9OoGp4PiwP0GRX8TerQ9UwxbO+jk68mu0TjiXQa3WcfkTz4
9vGHQGCVcbTmvdhPPzwvB/FmooI2RLH5G7Sxw7xOWtKYm9eAwzMsoGkMxjAw9Wjm
32p/EpEgIEd5vGbR0MrQLc7aEN34t2uzsrJ8xs/0CwYPrgDR7UYs8C5UnrfIzx3p
bIipttGmzH+oaVOxnN138jXErvAk6Ls4wHTTtjllQ50jcu96JVNpTrHh7zTYCTOU
E17wYtUu9+q1e+7VPSIAuA==
`protect END_PROTECTED
