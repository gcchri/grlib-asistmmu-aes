`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hf8M5AuJB4L7wkA16zOZj/EYamBhnRd+r81dswMKKVWXFD04kkZksUcHFzbqugKh
VwIXLD3lPMLBd8dY8LLauvCyr6/u7crs61f9wM1r85/2SS+UfZHngFRodJJt8pIP
xPDmYbGPGO7rI+M6OMNLE2a8MvsuwXrtJnVVtXmUHp3ahrtLU4juN22oAxHWZqg3
+nmixQQf5fiHgWFaDd7L8QpUvprq2lvtmOiYTXSAAnhkMKQhy283KPu02okMOv+D
tAnI0QsxnDMLBXAm3+DFR2R3iezuTLMKQE/RYd/mDtpM7WnP1NpV0v+Tkjn/Kjvb
i8wtWtUdChF4SGAAh42+EY+68TQ12PQSSenwY68YcUI=
`protect END_PROTECTED
