`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vOXwI4mERQzK0sFxA4sCjUJyWdEgt0M45MUvg2CWhK7Y9h6uZmz7nzvBwi2aIrl4
CJG/SSh8SUiCw9CXr1LzBWsoeJ5hMeKcjp80Wo2WeWosYScLv2LygGbAUEjmJeFN
EP9Dc9yqKcTt/RfLC3TgGxenSvUFlohrOTO3HTfD3/hGxr0Imc6ru12vLDNkt1if
9fK6BwJ9/gKoJZBVSL+V1zt6Gn/PCcjbljD9dhzXqAXzziGrQf259k6xYQlXwCLB
qsBpSen0ZX6f5N0xLPIaFI6uKhq7rqcccJEigRQEUlQqw84LhSjkCSWBpRpgvtZD
aEOQQuA+EhsloCc8ZPKOhQOY3JL9jLZ9Ay/q48LjVWSn6FMWf6K/LadycG0V7Is3
KJvtqwaSYu7B16a1o8BHDqh/meL6UvWLCCOJsL2wIsMeG1jsPT0SniUDwO+bRgv9
5FidSxUMcFBrr/g2+QMnHXxWUeJbO/uWYlHQAIemtKS9hfvA7e57DcR1mfgDpsCt
6gwKqyljniVNHvtby4EP7HTyn5lAIJxPFN14uKfSCI6XH2a2gxhdWZlbSlVEJ2QH
MPwsu+vLq9DqZJIie56lbh8t0WxdBdZwcypQ2+8TH35aJu3UXAsCZJ3h5epLdbL1
8HwmDW/7EcwCFRBBCtzNjfzsKgAxdzYHKHUfSGPSrxX/UBM5BhcLAWTaHj26b3z4
YF9618I1L+Hdz2t+wAEJ2aAJ8AoOQFkswJutZAG0frMLZtLYvTS2s+Bjg3WfDrF3
x2HLQF1W59L6xWi8/4K0LuBSLabZYMd6iYjTrRZ6lVryOENk8FfyNb7fd2rYpb5/
zaagua05lheUx4WGkyfgM0zcqKkQ84HtoprNwLN0ciH1etDduidF9oPqRmkA0yj6
X1JpFlNdvzTDeER39sXspi8ZU6Foh7d5MBnyPtwklsx9MK5p49q0OaHHm6WvczXE
OvV4nCFHk+8YV8/Aa5iLrVZjc1O6OKxgFcvz5JY0NrOBQYQdoCMbop+MjJQmE2tV
oKX9zpAcSxR/9YSAqyp3FHNGyGgEWUuu1t+uyBRTHLZcCpvY9ERzQ2Oa0z65RbJS
dWAZACxejRCclw2CWq5X8FaDQZH26Jwc1dx39pOGilJJzAatsII+fX9qoVwtfPyh
tH9nmMoVVWepGtUubFL//PPIzGc22jZkpb5WmhRT/9+xcl0jRaueLhcSjlUoSZJw
5LcdoNx7XvSz2ImszE5sDNCHZDu5rHEyeuCbQFLbxxnxOzkE3l3g8CcSxn+UbjF2
8Aa1odLOs7pHnGcHqZAkmfR2nlbGVr/vh7ZN1t6+Rvv3rGIRrdTYu82TCPVbAXyj
6SXHBOfTA8miUlODV0ni7W+DAK83StoHE/V7HHR7bbBpsbiRavLmAezpI+kG9kYM
u0BuFxasaQ2p7FEuuH2lG8HcDcdiywceor979dOV3n6IdhsNvVjRRhxCPZ+K8LSW
WdLTGVyfOboQRe2/0r7hTE/ZNgROTzxgvPZ3VUkgCfXWJntYoSCbYLFbhbGlxHmf
`protect END_PROTECTED
