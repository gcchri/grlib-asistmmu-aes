`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gYle2wjMRhpRxCmVk74gXhzWk505Nf3LlIJ/41UX4ecSYNuda90Nl6aInJOphoUM
feifJ3HsmwEEadJlIL0AQUZUVMUOrNHRxTH3p4oqMMZUxhtD3YSmni8ZTRT0KPX5
iJ+9e0BXMzD/e+f5G04lVZoTd0jX5EaNNNZrg5Ey1Awggn4QkNGlfvKAOvfafIwW
Im0Kgd0VZU1Py8DrlCAdl1uMrhwRDwXUXtonoZ3syZTaXK1yihW0yWxaJDa/CxcS
2E6hnj5EAKM7W8aQba0VH0eBMXgm85g4ATbHPL46UiYJ8hJkSUaXyJEomYElmDVy
jbQChP4meWVvACjFRytlgVosRDDbPKyvv4Et3IgTpUUcDWOGj28CmIjI2IF1v03E
e7Xt8B63JlZ0Hs/0uDmZX1k8pbY2YR0FSZNH6LaCFbRSedBWJLW6y5QRIEtptQgi
a/JS78tTPxw7GA6fIKzYQ3IfG5k4mMRw+ONV9s22Yd9xMnMX2Vi8wHXgd5JdxyvO
O6J3zmzqUHinzKWzS1ZeVcvTv6rvyu9DEOfd1/aD6x2F4uFBNepYxfgcKZ5hEZ1A
Z570i/SYNnrVBIrKvQYcHmuZtAFK7ZLdk/xKatcuHtM=
`protect END_PROTECTED
