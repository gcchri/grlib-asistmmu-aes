`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
En7veCD0kAd1Tu0nJqfwo4U1EGGd0zMc7+Su1IUFzIrqlhrh1neA4/gUe1qZIhqe
GMS9avG0M1lugGHkhHYV7FTaBdWqjQg5O16jj8EKlvaLMiRwktnnea7zBlMupmjW
xDtLzQgF7bTJDCeHqK8P1YkBQ24WmNMRLPOqk6ltUoiybR3P7B3EE/04OtLc90gl
WrWuQ0wfH9Ql9FlE8dpdVwXoLG5W1Lmh5beBgyaavApKDLCSkwaKQ9WeynAbUPtv
59X9ltDn3/lBWDvf8XV8G659JG5lOYGt7JcQQWOz2ioebnq0P71Ui6uXWDmPqVP1
mBPxcXJXJNN8Gw3oMN9IN9m3HmJkykR7g19mQRu1TOKEduAgOff2jOVVrz8iBEFM
lgF+3UTcjBsHPwMW1ikY5BpytFJx5OIp0oFBXADBQeUxMeJm5Qb4Zp95FFDFWOzC
`protect END_PROTECTED
