`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8USlXog5xjOcAZKuy89lCSzd0+rH9KWOGSCFBXsTT2MU7eJnfSf6PRsN/mujZL+
/ULR16xliVt0bW1jDRYuVSHhY22TPApEDW3Xtb9d3XBJkcDYGtosLgW/RSmDHf/L
3LnoGoFhs9fQnJuZAAwzhA7ms2gbb0D4IW2jjr8R5ea1T2b3LlU/RzLBlpNVBBAx
kZdKJSJtHnKCnKjZLlHpbkr1VZjOPAcU5rhi+1sLWhxOBNb9Kb5GK3+TwyEXK5+y
5qIvamOgCX52196mtkLS3lp6ZC7kaZlEQCGofZLjH6WJ4xq1f7SnMMGG0T5iiT5d
/OyYSbMImc5HabYzMxVh4Cckdd/HxU12itx6gna8n5XP7HHWJRcPJSUWHfhW8NBJ
0C4N5dPJayeASfEYKadhUf7YymTXvAlz6vIpD/6A6SoKvycvpHn6n5qgZLwN05l6
zek197gS2Bpo6XRIpsTNagotLqVWEUbV6Z4Pt0S5RF9lFjwk1DbL/VHi/M2xR6zN
k68ig2Ug8+7K5zDwwh4Hb0DMBTcNd1uca+0Jsl1oRQ/Mueh4dszOfZ8Wo9pYVLMj
k6pbwZ9ABQbslibR8lZOyw==
`protect END_PROTECTED
