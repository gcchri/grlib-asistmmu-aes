`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A+cWwfPnwAut22zP35pvgE7/KEFkOsH+UTMbzLnQTuOq+lrArnOIaWQ08bSVjVfG
2cepZEhw9KrWW6Ior5Vj7DCcFEN1xIyxTbvZ2whrKYSU5I8zhiJeDs9dTwjF/xDO
FO62TZ/pPJ/2s/zMICC1zc++nHtb874w+RlsCSUxgsoHkSZtMRy95f+JanA6lxxL
OlRxUsMZotyvmoY+hxjobHStA1cvzF6C2/vBt24SGzitDFBJwZ8PIWgQfq5cGwQ4
2ArwBxrv+h2CNrvgoLkzoqgZtRk62w4p5DEqp6nxB+do6Rw181SOPxHY1rwz/HTp
Yjlrp4ZxR+KETeIphLjeWSlDytoW1t+gniJSQ7Eox7TPRYZFBFOsPeZyqZ6sDiQg
JIjKC7ah8NdmiVXxIjHwHQ==
`protect END_PROTECTED
