`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rlUYYCKq860bcaCueU25yeUzcBWl5mkkkDVKEjCloL8MBvy78JhG6A/9xQw7DJOw
EZYJNn7BiH0EuJJ3LINdxSf7wKyu7GEinxjVf9UY63TB3nlZUTp+0QNLJVr6P3pS
0G7x80MNbRSYba9VXC3DoK0GWGOtXejDW+NAMmtP4Yjd0HYy1skpkV3Yrv1B3gqu
i//TX3hg2hgC/Je6tZW2bezKRsvECos2oQYA55Q3ilOlsFqy1H9rF0PWKx8vWszg
t/FlOoampmSTMSu7uztKo8n4X0Xux8FrYZNTq4uMo26lP4ob59zI6kCuAeTxYSFd
d6hl9B3GpuXtx6wHAnepEbJ8nzT5wrLZ4E7ne8yWNG+MV7XqGR8dYsskl8PLTwFj
`protect END_PROTECTED
