`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hzfdPXW0r4GD44Yq0texRODj2CcSioYLiK50+8P/5vHzRFSyM89/aaoCUMGjXnYb
CaMMT48X70w7Or/pTQWaT6fKa8ASEt6JLG1rLBdpbzY3BlCDK+mdFXy1tiJJy/gZ
Z0q4Jqd1IDXn8YlFxwT4lg0pFDXmAt+yoWuURrZkip14qsJkOiC96PDEnkdoWE+Z
bYSagHToB5y2OVKlvZtVYSS/dNT1DmuSNfxR0Vwbzx5JQYZiOTbvWvW7J06zGZlS
YFePPPdO8scGvpNiyWtTjsIynTxrfn87clAnQ7Z/n700uy6ocIm2uepbHfFb2doy
blDqxId/JWUf5/luqap1EghukYIuRrnwJW/5f6s1/6uyu/g4HG1xu+MAuxinaNNV
nAeE2HAmmmdm6iPz8mJ3Au71q9dYxw+l24NncvQFORP7f+Ybq4pHhd9LOxhupwfx
qErTcHw3k9+hn59yvDvisYaQYKCdKeCgFeUOG1Z77ZfuFjHSYNA7ztQc0YW9g04D
dBUiKMp7xl9l92pmZmcF2dcBAf6j7OJzlCqa4o9JOeQ=
`protect END_PROTECTED
