`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+p3BOldDzy6WIn9xBBq5G0MWsY0ZdhjXCm/DM6ps6vnoxdZed7KaLJFlntGzx/Oi
x90FKDuF+Lb8X4Oec0okBt8EKopNBdxc7KjOqD2CksEA6jigmOByiM54IWqAQC4e
8ROz3Zjrwx7Ox7LxfsgsVRignSKE2pgM0TRemxqDRJP8H9WlzJ6Zqeza7SbilEOf
XozY1gegic1KW9JgBGoQQx+ieKWp9WkoFS7JZEG8bTAagMZkvT+rQ/r9p+05Rzoo
cVRiBwDnX1MTkvmnoLdNJyRYVDof0mzJ41QltF9VfEHDHYmfWEvRIo2l4LQW+K7h
4mdn0lIpRFU4MmEmXrzs6E5y06fj+nWhp3rP5ivoqs62Imhmhv5+Po+BnbslA6Kp
CoyZg8voG5SuS79LebmM3fYXXK7fJAGeolk5rTX0e+E6jPjVir3KBGMFytUAs0oG
HG1aLylNPEgcK0a5rrrNE6tW1my8zu6ROVdqRns7QgnHWiduqW7azBcNPGEuMo0O
s51Ei7jR20+A8UpUPruNPm5urLl/XjAwqlYV683XQkyNL8CpiPlD0W+PDPzxtB+X
+vhJ8lCPPfosrnWRnMqaUxri/lm/mr3dyZ1b/Qd/4h6OyzgjD3tcqZHWyOOYFsxi
`protect END_PROTECTED
