`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zS0ll+Fa59tG6gtde9CzHyJB4yfv7d18VRzRbhSD+pp3NFxhWjyJQ1+E/WBcI0GW
cYyGEYA/6zzKjW7PytDB/Qm4JlpQ1F9jNowFe9vjqS7LPpZYadljG2GSvwHm06Ep
i9I4WkwM935oBruCCBWoSTHW1OFdT8QtxGb/iKhD7HxNyRVrt+yKeY6oHpVnVl7K
0KDnw2F532LuWO932bMJq7x6dEPxiHrkG2f7r68L3b55D693rOtVy0xYIHp9SrZv
AGEBIHd8KfRN6pUHfuU4786VKus5o5cpWQuWJUu/+J09oK1Fbe6XspU6STgpizb6
4RwjYPWyS7Dj9KPfXL5L7eWKo8y5oIk3gEWMzAngSR7nShpB3241QUpGIumPy1z8
+wuk4saUaI9Lyai0kurVHj6gPqR4P1uPVDMn7x8z0V1yrSPXRjJPYgS15vPKE3Wu
DacDSGBLsJgsdWD4Y0TlC0608bmu3Tn5HLwb3UpBQ2ZJRHL0dHxA/58aZmvnNRbZ
0Lx9HptEQs0VQi24AouWe1el7+vks4LcxK7umfpzIbhW6xyIbQ9KnRl4cnnERqZx
74+XUhP0lehR7vd4I8UKz3aDZaslhJy/+mMWK2Uocaq3ofc3Pifd/qSLMKX9jyjA
RaFVrwjMxBHNRN4TCTb2s5cORrFfmiwL58j4l4K0BGe71zq/2yl76ZI8fftxj4zj
T0Cgsr8PDtzNctOlNmX7Pbsa008fyn7r80QiEzgLwTvYzldsLpEjGoUbVGYTVlRh
`protect END_PROTECTED
