`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTCnf1rW107UG5v7+JlR20XTSiEPkDC/JwpKKraY5PpoDsegWPjTzZFgA/CJio23
e3OgP+Q9k32uoZkcs5Mn+ZSl+7RvFH7B5q5mCSA09wdZL8X8Wj2Dwg7yfDPnjglH
pKsLHjBPXPNrtHZ9CxxOHqtahUcTf4uYxwOmRbmIo0Ztl2x/736HEGMQdYVg/NSk
mSWDkqiJVwWMZp6d17hN1Pp50iCH/VhrUvo1oJFWphpsna5XYq2HLlIH6Y/glDKM
YtD6CHADgcBz4x9kS8dAQrEb7g8vV/v/D0uzE92i+2AaEVSTNehdTU4mHYhFMX/R
j78W5b5F/Iz+/Jnm4wi9xuwxLHt/0tp59griyC5CTwJ71VU67uygLp1A/4tSnPr2
ejW2aeAoqUrwel7fh9oiwYBC5893UV5yM4XbHREutYZIhdjoOJpkVYHi1xJ/SLAG
K8W3PbGeibeLvnPZ94wjeByuq1/UsHLqW872N2SxhlniKDGfRm7+zlKMVIzAL2+i
YXC0DyOF5z26+vGwh+pC2NyJl443KcBZhSQ2WEWRdVEpmmwpovy2Zg/8TgXni16m
vI3bY+hJ1P0TzFJwnHPbQVogW6EVAOiSuAc/djVbl5es07YcMu6qPEzpo8zA2PIF
8k7msCfpNHXXST3ruiis4gJqV1nGA+U+ObMqzGMQu41FFanK7b4cqHHy17QKplen
lCvxahUMhxrbOYb0oAOHZCrRt3vpfSR4rrFr8ILIGtcZFVB8sy5vpZJvSjQzJrgW
gut0rTWWha8ZNJw7m+VtJvdGKW2XPsHDkXVK21Hnp9SCkaDwt8UlPpKxwXyKLaSc
+oPHB41X2jNGByowNsdcgYm4Oy7hyv0CVYgtTW2z6w5H5BFmQqaN5zPwRRw6chZL
qG19a8DYvRxLMYZCDoVVBW89rgamcjNDShvRFkTn7x25I3sgpE12zSVhRStLqjwe
YdN9M7lmBvmiUW7VEJOwKF8iKnxz07FYL1oID00wxg8ECm+rQR+T+HxdkbLYGg1+
ib3+kG6zJ5jyzlpNUn8lEiSotjz9gexo+lsWnd5mbJBSQzMRD1w7Kun3DcuQEFQQ
4f5MzarITCbnQiVpO8xLxxEbTvRSSV3fbDs1jO55RONLgR5UnT4fGSmsm088hoKr
SLJLxq8MXDHpbGoGWkBAkTFgBEr2SYIrD+Xm2gfVxsagpHoIWqO13XDuSGlEC21u
zowbxW4InXV82xSIFxnXDVaGNBv/eZ1qjS0svuAuWl8Cqyd42sjbnGCgnxvMyUzC
51+XIkKqfd2ZUrAft7KaE1R/IOMVnQ+MsPdtAE1qBit+F36yfZ1o2D01VC5omrwB
ehiyTeYsa0SGgj97ZgzP1Ao7S0Ile0055yTMQ93Pw0bbsU6mSJhEQX06/YuCQa2q
v1ha8tzlv0k/R3y5Q0kBYok/n4C7CxfQy0PEnlsMzmKMy6dA7MQCd1C/MmCIpFt/
rVpQuoECoS33HH9tm+HIMEj1FCIWvKEFCsH7TEv6OFbNrLtffDRql4P2Qd6SzLBw
jew7RtcEgwg+wLsBOHTczOjFSaC/u8/Qbx2BITQOhChWitqmB6J6mCj1SK1wYbdc
`protect END_PROTECTED
