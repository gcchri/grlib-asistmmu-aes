`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QF2d8SKEspbHCaVUAyqp9XqiVJVwQR2vqu/s+dvFR09U6EEE/X/7/QugC93qLDGx
zZn6trtjOoAyFCXv1UURcSx48rSa0S7Y9xlgqteHIec/VZifivj4aZIgFD6OcboJ
+PktDZTPDkYey23YpPibaRoUfRCpuiskjvyn4JWZMKkFdnWxQzxuJh13Ayk+YJT7
MvMAGG+Fjw0YPQJbp/WyvLkfhfD9IHOXN7fg3n0QmKg2L4vHgRdfByFTVzwi5J/B
EQMd+RqsHsrRmZKVwTIC8y7ZI72BFofgZs50qiRsrVnbjv9/NmIlA1NWrzYWlKzf
yQYw8NwG1Q2Q/2W+WZGAwZkAMhsVSFIYH0MRmKEv8jpHa6+b6JVdNL22R+jIJswB
dsb4fe6wiGS3i4gbo/4u2QDLmbwbhTn22q0oh/wh5FDeOwwN7JjrK73UttRnjHta
t6GmfFHN5xgR6ttx1aRl76zW+uhheWvNMRKYFlzucuyMN7gXkdm4UmL3TCkmn0Ve
UHszG1ZToheiJCaAs87awOBvSarakjNyE7g75OKB5rgDwtFVhz9S7t44QZ/HCDNB
tBzVDasHQztGlwiwN7dKoOQmrpNmaGh2EIlmfWvrtmETs32qQ3uOjoGhnr/gjVNt
fkCNRF9t69+TuWBZVbSrJ0SBZKHdOV5oCcWErkiiCP4JVcI1ZYXv+2VkXVTNTAxh
bG3d/yi5U9UG9jcq2hs5u21rUxx9F7tmDKP8iGAzpZ3UvPjPx2DB77qp9v4b6b/r
dcJGkw/8kDwIaiaxgTQes+1w1SQbzSlTfg66Nse3IQtZ97/3RI+pvu7BKPmaF/AJ
QfIVG3jkErS4/LAwYbqDpZBJHORfJcu42oUyCdi0jmgYfLlhdLvYMd2Le7OTulVv
RjaQQHI67bRF3caI+kaSfURCC+80KO1Y8LNShzX/kzFZPuCC5h9W1nPhFKFjPEwp
NYgqcJdwl/+0B9raVVHe411DJBA3K0f4jzJV+XZtJ+zo8WqokEj3WhN4hjZ2KtdF
7mPwNtiTx2siO8fjG/z7aWcXFuSlAhnQOKXL2AN1n6T+k7Rh7ftfkRy93AbJfwer
v79bZ96xf4eD6CAjh8IswdG6qh/zKRFW5NJd++xlsCsc6aSWcc/eFYA1Vt6/oSaw
IMLg90WPf3IehRXpsGqVWdPmNdzZCIjstPaOzfKRy4h5M9GoojdH++BNQxKcRx/p
HtFzEczYyvNfRYYcMx/G5g==
`protect END_PROTECTED
