`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZlVXwI4HAy7mYw0UWqQZyNc6JME9ovMrPDH2aqZaa8sCXszhkYRhod6RnWCDbRs
FS+0FNHLh89RvmxN/Hv1Bq9uD2lD+r+iBXmLUDP6OSrcdiZEao1LwbnYxomtzVDp
kMFeI0k79LVIOHLU9QcT7sI/74XxZO1t/J5NWaLxrbz9R5lb8JVdaGAGXRi72RIJ
NIeQ5HMBksXj6HZ7rDDzPFAubl8Ktv+9F48uqY7V49Ipp75Wj5wPHJqN/J9peAzF
sp9aT2mkNcREO/AgYbD+3JBynt/rP6CMZYNdQ+Pw1B0Y03lsClOQFPORVs5NrGOE
9ByajBAV5reHtcml7+75ZajrJuP5ZkC7wYIV5JEpaGSbUaiXVxXAS0XaMnf1ElFm
PPTjH+DYqEjBgzkemXfQgvrksvHmls29cpT0sb9iPcFM2djB1q/5efEUG9Ns97j2
pbHPnevLUSqy3zlxzIMDapJ9SJpNq+difdT9RCtrE0RD+5Q5RFpwwZ4YtGbGtmev
hsr+Nacz4pXdourwniwyzmu1s3BfpeuHOsTVzv+W7A0x4bGf9VJxPlRalXcHtBma
+fwKaMeXDJK0db05iu+uFhm3XQKLktouAlA/NRYUgLMGMZ+oHOJfyr37dNh1eomd
wHWlleb6k1WFkGOV1SCrUQY+3tXW8iDCb2ycEzmi+zKsAOrlEmhOGjnAsZ+iE8YI
g7gYMkD58zEhkoU9K/8jn5Ejn+vG2lpW4+lj8GARSMWTvdFVoHDgqtQH/2fTPpL1
44DkCmaAKEZVn+GV3uJ2zyRlu/Q4T0fm3Ku+LoFJBq4sdTaRKyCkwCO1/GZTIJC1
V1MASthl2bn+4vrcyVcqq/+4JdGRGwjmLvn9ehyYKCUMzoMqaUmVpOPbC6mqEMK3
a8TboLiWYGvaC3IPlmb/3DN17ROCMK/OYWN/X9H2MDmHZHp6TQdgCQAgrzRIAO2m
bMXxudfTmSmpar6biKqrUmYti0mQhFBTeiIzwg8IdAggXi5P1xmEYZh7S6tcvmvp
/vCi91Wu+hb6negzxMuRwKnpP09x9qdTkzAEeXYG658mWQlUve8sDFoD2XazTnaS
ANzWQDXH6EFSDdZ8rvjhlDfDnVeUJ+yG0McmKu+IgpnXMM/NIOKA16f7mFuaWOPr
tg10vjcDf0k6ajhb1DZmyI9d/8oiJDrJJFLcN8heNFO2a3pSrrxV2cz5Hjl+8tgI
9o6M8JcVVA/F34HzquzsVS+srz3kg8PySkZFDG5Db2NRYZ3ELIlA0yDiVGi81msh
X1CN9cK8RkQdItppaZ6rlSfxL5rxv3FaNxU2pO7RwEt0SrgVDO9Fe/+Temu/YTvO
papZSSkZzy1t2ZDqBVeCuZQg/HiSuwBaLaFgwDtINk7OHatGZ9oDK/752q3nOH4E
rE8CuvbhzsN1S9Pt+uSKBmuzqXvZLIfcbgjfjkTyz4pDNaq1EwdheaTg1J1rFoIy
shAze4aiSkJ2qZZ0Y+gDaZ0b8PLg05GDdJb7OAP6xXtnAsyEdFvmCtSExSTl/hE1
SV0M/LfFGIc3LwEBm+qj7UrjackmH/YymYHiSkCNUFbxKoG9zEHjTG1qLbff45LW
PXWkJI10VaXRI6IdfyJcj0o49GYafeBaprJUFgd2/S94hxdGQeFtVWK7D/BLYSRg
TfyQiDOH9O74z7CKo/qzHu9mbbJcQ68/w2/93AdolNJHbKDn7P67wAJf+uva/mov
ULAT3OQdtdOl+LezpmWBbomXjBRWar9R7YbiXXdgXoQQrYnpgKEaKHLdJqgT1ave
Asi0zhwVG3+MoL7fHeeBd8iYy7sf4ImihCRCO0G7u3EOhmp68KeGgZacssSafOEk
8tWOhHydqHtPIQLc30S7UTiCBXcWLYFr7c0b/o8vTP8=
`protect END_PROTECTED
