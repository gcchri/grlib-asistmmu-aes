`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Fbu7AEYOqtLzWa9WQYpuDAsskdas48jQFCdHG2uem4igK4yoJcakkN29llXPza1
vv2DJM/3U/A2qILy9yCCtCZqYZy+qQJqgbvcePzhYyh75kCINdl2N8+ioTEH/v6x
dwy3+FptpC7ro0ApmkRbJIXmPauXqdDsikN8ce0v0bWi3m+4B6PzaQTUjCDiJkQX
27qN+kzo1LW+H4NnF1L+K4vOp0rshnPj61H95NjVw151VazFw2UnqcVsogx15lEI
e5Fp1Ag47STbbysGVIl9GY5Tcli9nWd+GmVqV9hhILiRPred569daFvo7rQaz46o
RVHGr0JRDSxPYdF1FLKeEPAU8/MK+Yl/Z8xIdT9oao+ihNg16Qpa//KiU09vzf6r
`protect END_PROTECTED
