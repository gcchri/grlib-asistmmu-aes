`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JWg9fRKGXUmwb9jbFQOjYmh54CAsRSKI47L7Adtolo+4KRCp3zGofsySKA7i0I3B
4qslbgRgrVCGkEe9xobp6abRkrllXrTNcdOSeVUi+J7a0J434L9KxLwq+QRRbGJ4
IWGhBeE5JJL2tS9f7LigqfQV/tMwj3zw5PgB/T0J0YpcRmEEUX7+8r1ninERRuR4
zQgFwtYcFjyt9qhlWzAIdiWGDxn+Z/Kml7c6FU34ItZm1iMLIfKinu4Cs6ad/yTM
17i9MCSQ+eSjwCS2yGnkcw9E8wviwiLyodGdRfB6dQWDJ/cWLXdcD2sdww1P8eDE
z+D8Octlz4nD5mtpeHLOuCN0qMEkXLJenH8Sw7jc84S7FQ7a0uVjA+FioQP8gn11
P+M9Rv+7DM1gc9tzw04WauL8k2x/cbcn9wRh/mfkH8YglI/E7E0iDSufjDjrmuaB
ugphpXOVKZnnxzpliCzLivqhn7GTluN0cJkQm7DZultQGJNdrV6tc40nAhc8nzvP
/4J+mzYg5urGHO+d5FF1A5fkk12r/pMPBLii569tSkeyIjg551IfFZNNG9/DdZ3h
jhVTiQ994CsgmoTdEdBNPcdlJ8GhAskF9Nh5HlDn5+SSsjGoULJE1mT4s+XGS4P5
SZJEqzqfAvp4mMVKmsSmnub8Nb6ewqzmmAXUqnm7Wse+9kINWQo/4TDL/gSNp989
4OYeyEoAoQU0RviJhBD/8QVqIHez+HnoqZrNgikwCxHpkFbwEpYpZ0W7FA+FKDY4
dvjrZm4BxKQ21KiI8PDWWSxWve64JnrSTYQSZQcJWy+mUyiMVvjqJkTt5k6Rihil
SNZ6r1Plyew17Lgu8Ove7gc9d/k8PZtZchPbQ25nTayg/nLeR3jDwcKLoqhZ9Ugh
MhJEX2fivYq0QkmmuC+J0WiYI0pFY31DDXKzNrjXAeOI9w5W/iXxH9yTAB7UHEHu
PI8JChJIyKEv4xbkKYuLPEmaOBGe35UKFLLy/BIPHXGgpGAdbW4D3X5Byw//K+ym
O4eEFNJKRO9tm9ICItjpM/KA16ZcXc7/wHTdas/blfGjeImbIA09Fp53IR+JUUkM
BOiCmC6REp93OsJVMEVeHbz08XWpvi5uLa9CxWJwhRuE1dBUpuCZ+AwGqO6h3Frx
cO/zWArIEW/kmCPicHVGP8UiB7MMYXClE+M6Ipbog3+kOn6O9EKyxc+Q+90V0wmm
hbRFtJhW3404JOqxnEgs3tFwqpf+d/dHCI1YORbNZyeJsV5E0+OxD1WHiF47E7Go
jAgHP8Wb1bh9rB0cCNL+4gV2DYhXcYfCKRJirsFcpIf6hY/DFr+lKpIXNHYrLlrq
J8D9NVUcziLiydyGI85ejOvLDrmkq7WgQPu/efoLiE/zQ/+131tSzozc0gK8yySx
uDqGZDXZ8NgtxCEPp8UrFaWsvNvUbcTvD21noGq1clZN+0FKPG4VIB+dMUWXVWos
1JiGPo2UvWn5RWmOYtPbza0FpTke3GQdgWxWaz50vnAZfyfbuKwi2dBdGDve/SP/
6Hn2VQrcY7iiVvsGsPjnxMc4mrqSqLr0KZShCa1i2qYHvnG1tSs3zMxE0mWbMRuy
ajWN38atfh1J0nuspktXYiCadXyo/QLOBC9G+LDSFL2zA6OzRoiRQrVGOEUUQSol
Zy+xqc+uDVGGSDlj2upov5m6OEyOjcJEXbTs1Jw9/Tq9YBxt818Lc/4yZcJRopNU
4WzHUSdD9NYzmYnSRFUAb7E3EriSQwhyDE2ETDQ2l8/ov2sUH5qFwLlhObRVNmdr
`protect END_PROTECTED
