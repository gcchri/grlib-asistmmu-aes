`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iKEkeBguMjiY0Zx2JrQ9M3bjodR6ZCJ2QoU7PVMF+/MAGApGN2b54cR541+NOnHD
aOr3XYb60zFSHJx4ek6ozQPSOXBISFjkms0IBRSTj9gdebW94DTMRK8zf+R5gMAW
Nf9LJzhLlmJsmrcESqi/1lwHGDcvuFKjl0eBiLUxRfOes2xcZF69zXJgcIjtYkJ0
BhcEArDfGgvwI+ia5HX9M2d08xeu9gU4UOVHK0IPcn6/nJkMkRZ8Jt53q303FRu3
E3dik03/LaWv4xO/1HbBq6xgNA8s4CQPjc58c7Qcvyaw+XRZ+L8OSWuZ6uVHlV+t
Wq7O0bVujIYjRCo68H6i1GOoJWe6RGasDfdwNrFNhXsKGcS3MoqwniDvqwXdDjdM
CaiZBMwHV5NNxw7uwpB8TxRv9gR4XoklUIXYVaFGgDpy8ws/OtWHXb0bj+VJUCi3
pdH9W+OellE5MGKcwOdabbq315KAAQaiqYxc9CmGVkY+d7KE7mcGf4c9KjjYZCys
+Sq9LgeXE5BlwR3BMUWIOeEPA5ek7L/eSFxk2DlyoNpSnnTaf3ETxUNn8buCbtk5
l/ZG1B+1ytcRbqC3oQDnEBoqmx2sEsxVtB12/VvP6QW/H+uB4G51yOIFRK8bfzzR
XYNvnyKpxDK7270/leVRSA==
`protect END_PROTECTED
