`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9GgrH02F81di81XoBzpsYseJ8V2YSsKDGdHBLroH6IQhdPGzW67y3TgCXEU88Gbu
21Pe9c5tk0EdOtzr24aEc3Rl7V7yMJjzEi5+X7jHzVFlduZQa+KWNBo3VKKQBqm2
d+5yRH+jRhDC/IZlZe0eqzXZa/RU13Tl93hMWRBNoUcfcZwGGr+AX5Llf3qE5v3A
829tZkZ9BhsWLDvgFqDKanUfpszHGCbeYoxdaX9zsuYVFL24IXuT4BFFvDPUY3W/
ivUtEHe3aR09jK9H2Os66IvU3dicSXWTuRtAJtpR7yWnAuypK8q5fQZMFY7cJYRp
UzjngIbhxKpWcs82x+appNxgZARsxCBYs9nB1ucutMjmapVTdKTA5TrJpfQcMea4
vHYPKiGGMKnN2BCBviHQHosSv639YEBEq39lvx4Ngra9inqBveh4nXe16aBofy1w
bBA8ayjzWhphHoZ/uxRadSvnP8oI8v4zDM4hKWpD6Qbg+WeYF8lAbEbz1WFrXedT
mPC4gz9lLv1Ov7UmxLTqVQu/giBeRtdmdGsRlQ6W1kTZioN1Fn/Gas81MuzBWkS+
FVxESEXXgdpv2ID+fs/ooqfg2kwZCAmvd7fSs/LaFSVVCMKbXMa2HJE045FbOtDo
7u2UbdV2A4jocynSLbWP03mMgxEbu8hGEaaam/ogDmdO183MtxWbQ6cqwANw0TSa
TzX45LpdiZVlXqmIj1gsc70NNBH7lVfoZFGa5e+O+343AVnRy62nCf7/rhKJ8vOr
Ec2eiPklC2gt62MimYoc9ovxu4zGM7XCsOHqbkQx9Xg+78JAKfD7f3dlL5Y/9BCO
F4G637GXj8gMnZLhI6AjmuPBExnvtq1KM4SUxRwyADlPCYZfmPzWf4n/gH+8C3KL
NqLontVHgvyhg/wwI8yNbgjWsYwJ/CN7XYP4KT+MBT2IpAsbKMPVBFZkeyAWvFfR
6mhIh83Yo0Dv36xWgtKp/2Whao17SreFZK14prE6eRJbeCqnXlnOGo3IrLyQIMvk
2Oeldx4jVXm5BFlHQAjtx9ZHBFDMP6PT+6kr5klWHiR/kz1JIKRW/zU+xLCecqsO
KVgHt4q120q9aDc0JAr0t/Sm47z3jQeF3qPIpxefbGwsCD8zzPOwEFktW0HU8Fi9
kIPNmQlLFXVxDgbMsCpbNGv+FE3O5RLjr8MmBxQSJMDCbi71uPrtK67vFaKlU7Lc
EUGM3ynO1w3WHjroyynQYim9WlEosfVGzqTiMjKHXtRZS4DXZHV+yw3tNU3B2l0x
ZJhSyEXQC27O5UmSe7TiypZ5bJVEgBZjjSATUokyQ3kRWg1O/Zpq/Nz05nar+B3M
exWuJY/MxAMPZHy5rmire507HaY1EtrWbvaQzdejR0WWajPn9uvcpr2hlJ/tWYdy
k949nH+Ca/JI/HJB5j1uBNYbSrJm+RKl8B2SdcSzds5iTkQqE2u0EYisbg4UBUcR
KhAM933lVn3C9F/wEda1J3hi7o7clqAnfqFnPgeimLRJJKvHquwIGjLsc10v4Q3/
0d9SooRcoYvToc3KKDmFC9WVP9fBFz0AY/LEa8+VqdxeKCsSnk93uvpKSrCRMm3R
FK5LHpyvHJeHk2sI3rB4gZxjZ9ytVyxXBCAOKKKweg1NtTwy38RCQctflyw56of2
cVN1FS5VR8kvF05tnPyl/fEnHSY7VOZX2MegL2PMNE6snbjciD1vK+rjyAPltKWf
tche2XPVsfBd/iYICfuRoRpzYEEjWBBkV+5s5AtwSE5I5KkR4SSh+wh3WmCWmLCj
pFRmy6jGrHaFfiGWN3kimZgFhljiR9zNfJRQaetin7F4C26XkEuPvkoDFGSEx/E6
WSI0HY3AJnPtDGUtpLACpePJmvbYs3bhk3/afPLEugvYRyNkqcWMYVMdGJPEc3gz
QIBQAmckQICvmm6fQaUc2J/aZh4H0MTPNr8y6uk4bMa+bAe+o1JAz4sSPe6TlXmo
JL9war8HyVOc3xHxwgSmifDL8nZcJ69thTq1NQGoKJA=
`protect END_PROTECTED
