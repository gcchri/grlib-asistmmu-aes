`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B8OrdAFULIctHqOJCpmiD6Ep4kPozJwn8YMV45VsV+r87AG2v3aZ4u7DAk2UpZF8
I+gN6AQZiH1F2NeCCqudyDIVoXtMwwrX56SKJUGvzDnrg9C4YRMIXCJH16JSWMC/
VsSiMpBvWBHMzsDICaW43X8KucadAnsjCB5WJl7pluG7xuB32I3IuRE7HTVhnqp4
d0vlAR1ZhbbeiPYBljcbcYnZAuVXYM9ZONnbKfNrXtwuLMe1ihHUD6MDs6vk2XQH
hMi4QF5nDmx48DmVhY2xdxK52lfgkJ4dyfdaiA788Vy+GPECZqQEBE9m8XXgDFUT
XDHAef5gTB6cJzcZT3fTIwCjdEfTXHK1q4PkCvP5ARI/auJCetSJUI+ZwEc8aLoh
RLohpnJjEqCecpj080cUL3Mn5s06CZCBSL9gYzGlANvZkrirDIhweCixP+cGYrwy
hDp6lSrhxE6QdsYk2u4GWBWavoIA0PHI05pjkz8TblvP4Kt0uNtqnr9oc1X3ued2
pYNZv+XraJLod6Wf/Sfc5I9cEXF34I7/cVYulp10uScWggnF0HcaGxXjoWlmoQyT
`protect END_PROTECTED
