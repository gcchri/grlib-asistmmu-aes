`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
so8mD22pCfo+XEdfvYp92Iznj7TVX2x7dJbQJTrhZTC2Sa+W53XybOxhLKuZu3Ag
YUr28B3UoMMN4HSgWUWOdQxSG1Ub6rvvifySSbAfkhXwDgsFC3t35TNTRi26lbry
NS6PpNxGoqwQOXwLVwodA3Fq/cb3/rsioufpPLaWAtzupZKB2foOq1BE+JUwQjlB
cqCqUokvsHZ9/1CIreNUKZLX1q0z3j9AhAiPA5axTXNr42Gsc5JDBWqtXRfiJ99I
rDqGrvpEYpzfvnJPc6qnGQ==
`protect END_PROTECTED
