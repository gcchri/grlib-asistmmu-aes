`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GasH7hrGAd/gmSKkjx4dPaEr/7p2NWrXXo97zZ5bDKrpSvazjoCTlYTHBYdFvobx
j3oX0RsGvH/K1Au6JpQEvxdf7k+S1if3S7BwzEFMZiqiBjMBsT0IkOe/7EkQZPoh
zAVoUURTGE0aBqRvQ5XGDa4S/ElUWsOk4XxXdBedrO2c3IGzX78muTkh2jtXId0j
yQeBaElNwEp/Jjo7SxaXJsy3E7eq+qiMzZs3FwhsxLmqCVGZc/OithlDNm6/u5In
TMsWx+SM4Vp3sO0RBguZ2cpN53pZ5oenbHOFm4IigYCUvace65x+zx1smUXC53bX
/O4TKgeWrB1xd2TkjUCtp/UyryoeeC4GgsLuR1rPDTQX4qOMdUK7EJ3lUnwaeM1d
21/YnTJb+CiFolT7HG3C2B6sflb0/kWY2tWuqaY+mPH8t8pdm5hco6RAf0xKzMbD
17i9ZihhSg0FhIXfKAE5LqLtbZkIBm2nJWG0YT7GkfWIlulZjb05uF/fAqg8QgIU
ivYvfbQe3XmiUKKT8+5RPnfJ2M8sI9EjHByNWoQmYVPuLEQZHR80vglWme7HhH2z
AcvdzucfMKFTLePPvcNYGLFMSFN0oA36X5BYI2BQbxIWxd7U/1jT1r+pYcuuEBUI
jsiha2IXg7g1DOJq67t4iSMk2sQrEgX8VDVXa4Zr1xd1xDhTm3LO+N4GDoEDcPc4
wbMWF8RMRh6P/E1TMYtS7VBS0P1QQh0m8Yl3OROvZ1AAtnoecx3+EH/M1DXtWrVj
jMVlyzA00K5zx0uVQ5SsRVD4GeW0hpxMXkfyDfaF3RZ3p4gu9T8n9irMs2tZupQt
cuMDEPjM1wyvPy9XgUAj0qs0PbpagGmbQZF6n6D7Kq2TpNGRAV2Kvcmb1rpVquh2
Vtub5PYKOxosDnC/jpsjbnfajouO2IUHcjXWpTojzjHDFcozBFAMQnAp7Vq2v4m2
4rK/MPHYMD5hMOtPeRCO+Dwfs7IMZ8tjQef+NdTKk6XXiuU06YXe3dtEZa05DWhJ
/OY7OqQOnqUuFc1Hgx9MJr5uvJ+ws9PiRxL4Y5co1pltTwiVv/8GfRfiiCtg2GRW
S2gjWavO0LLPD7mIjIJ++Zfockg4vgs4m9IlhPkaSPc4s+EqL8LFGvwcYicT+2ja
iB8C57rL1W/dzLrEh2L+bB+rRQONSSsPWiJ2ZZEPk0Mb86VlOLtmIFyXp87aQ8Et
po6isFdyXVtFvqXk/U/ObVE7DVG8RvSX1ghzKEZ7szU5QmqVZkTZztzuEDn8gkfv
HwI+zZn0nvg+ROdAiJhMKX7bKOiCYMGbYsMHamjhXTeqvyh2T3LNsqSifPmBCpc9
8AX4BqchVgUEHvnqSi0FH81awKyH/SGwKRZlWn7OkOWc4aFGXxz9ba+8hV2CfoRR
RUkyxmQWrp9iz26EahGDo/NYyRAj7GurGq2sCVyDkFe3Kgvp67oRswBP01W5ZuKD
emh6wUOLJjFKtOe+qWsYYqJtmUw3wZCb8/TePCb9VBmMmHjH9bXLLekXRuiHk3nq
8HNj7Ok39N7TzILhyddriSYGCajY8LR7y3xZPh9GrPU6DlDrcBRrHR1AcXxMQzCj
hDgERyvPRrOkOUialWtFeNhiEsrruVNRmhchSAKrlynG2OYmGLBvkvf1c5ATnJ5U
W6YXmQE+hNduryfiHnrVfTERq4Gp7T9IMaM2bh8l61rLr6qJh8kti0Z711F5hZnu
vjJ8OmhAEkT1zW4X/4yx6N43/JcwoFHmoNLkno/hkuXydtCIm6zn9LY0lfWtqrmU
ANvq4oDv1+49NnILs/CNGixvi5i5sW/N4uYiVTyR1zj2kkknly28vJmeeccY2376
wtW98ZP8OWIMM6JLkaXhe6nrKpVLxf3I0XHPCQ3aO0/aE2bchF7eb5RB1+F+9RRO
6NbAuEF6Ez4jNO46qKAIE0nhdQ6UIhuw0Jon+CEYW3iroE6XwfUdLLabamp+JOdz
zKh6NhLD9b41AQQrzmXsO9U5qi7kJ6lMBVRn+dupyj16cA8SW/FL+cp9yjByAgRX
uuSdIr0eE6g5d8R5FS654TZ1lOqzOSFdzxwZ02xi/ZvimyZvs5PhgZVWUotT4+Ll
eRNfeVHF9RzWV/QxtruttTDU/YvpYKWHUShUoI0ewfdBC5i05GxWGFawgJmlweYe
ltS2X17L3oHsCVGGrKMhn7PnibIBv0PCNLJjEV28qQMvt9GJJsA/BxMvEYhi1M7J
nKvDdYdL3iQEiSrN+8ErZN3/OfH6TK8MQHzvIa/Xt5YuDYVhhE+jziMdrdBmIsTA
quDPLVr463zKkM3TDl0NWNRp3WrIXrkXk49Gpd/dfM957/Su2fdl4gGaC64VHCfs
vPiKnq3f04yhfo5oU00w/a0xHyWM2vV6CND2Z7XOJ+IiHNDD48xlrtg/mFjIe9GA
G8t2BP3OedgpxiaPCQl7h9ytaMR4FW27wYsX8Um/tOJ9SMqjTSySXgf8ni4Gp2mm
boHdBX2xsUAtcdJyHlQsfaclGvCVS87XxowY9ndxwUi4S9YVQNnx3MhEluLAjGtV
QzjYPZXorVEOjAtocpzJj1AzHOmz5f6tVcy4UJx6PK3nfM9U7fVshHqU+f9muTCF
RVLlWYfh1fdMlWjKMUmYRO0NMvkZcupQCTRHVSDpGzkUnJzvLveaXwwYwXDZUyWI
U3CJ7TLKYa8GvNCQJ8a+NftWOmtG2XhhbteUH255BRCe4fBtBM+9swzMcjqyPYhS
e+kZ0Bx0n/ausg3L1R9IvPVLWod640knK3lySVLXQKFdZws2HlmSjZelr1KtZfZk
0DD8E1FTDOPs29UiloG4IrEnRF55ubsnBPRI/VBkA1eAGpurcYEy1vw9S8l+bag8
LX5iTfM/MikSoukLZ6kPIcoXnLalYN4rY5LFeL3p3kzU69t5Or2E8sPcBUQhxMsZ
6g3S1PGUR8vkXEbzLMcGQoG96QogQLn5c24FppwTegAcnAd2u784qlrklrtOySBE
3t6QK0K+i7vIKk7cQIuQnDlEecLqDr697BfRLMvTJw11c/SqRCvPI9WoQntlezei
UJ02m7bxwjLePFGzsMtOE4M6QAxeFLeixadrE79L57wJ2wtj18zwwJClDtIjNMOq
6o4ahpIyTJU7N/F1pT/KMy49Vt7HsmzyhMsoFLQOWcGvDXGp2bbuyfEXBRZ1iMQm
mJ01b5UArhN7mVfDZyIrL24PYiVqMsm/mtTvLEho5a/wICi5EvYJoY74Se2N880l
7kX1+ly+4P2UdxLsL2oLXOnTP3DwJJLykcAsrXRuFd3SSkugAZCZG5zJaRUDpC5F
BzA2MljZpar9aXnTumhNyKH3WGbPP1wIAv+Ju7CJ5/aalcRCetf1uyQSoLSluAQi
9DtOAXTILc/DYgrK7iwewq8iUGY6SfeBbNCBMI+dl/zz4O3Vc0PLPJWoZdEAQ+el
8Z375CTiDsbfEH5pcHRtT2/zJVw+PfvADMGfhz8j1oOZjswPFsp2DeagReOgggvc
FMDW6HLj93ev4VvK6g9ueJgF6WrNoMAIHZ7I9VfgjNMGLmvWRQTD1WQIEHs6zsDv
YqCPRCBvCT9+jpaqMkCkLx+hLUJKeFqkB5+l/kiV7K00j54xfoiNw3h8yFKA+V9B
4zXK1j7CTCyO6IgVcvwxn9yQnCjBsEYrJ5pPQgeWZGntfwRF0cYQTHBT0x8WtC/T
lZdTA7CHGxKb3NKrBFBxRBvJNTkDZt8DxuPmEtGnO8mVPzkrVl7mDIePH1BbtuoR
ZAvlRt1gg85DILZcQ1+PfA9L+osPkJRjRNF1c5/1O5j8P1fZh3KB3tKAnWI0vXaZ
xGO9x0XK0HSx9fwI5GceYCKf/jmXeleM/aMbFpscnrnqWYu+qYLYTDDVeCPOMHqg
nnuONlT2EFPO6mS479Kw4Rtc8I5pleHMu2KRUa/QBOpSQlvAbIj4n/uxHG8r8NN5
CnluuPvAeMydHyyyflx33qYU57jggPXcfGiNyJlL3Cv3urDFlvlFjk3jYJnsoiOY
iSwIE6T4DtmqcJAq8MhnfLqYwzZ8p2y59n3SrjhNsPwRfIHd9c1SKdsgfujDbYqB
s7vQVRsaQSkCyZuoBaPkPSr2aHqPFTAsm4iXWmuAe/Uymzqpq2UdxvJ9gcLM5U2H
8JfucCSGremBHympD3z83EfpGWqpGxZ04P2flv7Mcr6KlXVX2HD/weY8skXgSCcE
FKFldtzsjoq/II0hCtJnZhhmeEAKmquE9z7Sb4yzS5zmnX/pTxXzTiqzcNTOKp+Q
JqsOcLrw+GWxrhx8Uzj/R+6u0xyUIqhCAFfZWQWnN9dIXRSFYHlVpBvR6lnf3Z29
50JZ2AyjNIPuz9hcB/pJCf17WHb20Lvg2QUo5INX6Of0MsH55TFayN0VE6wUJPx4
/8YjmJ8359tf/NKOF4UIGNAHYWIfM1Rl54bwGHMrMqG0k0ZQJjcOdoL/mA8qx4EC
agIGlTj1c2+0plPq7YCGSW7tCvE5hkeUI7XGU25bTK3F2xDpANfR0/55zz1vkt6I
GZVqd+ESW687bpvWX7N3ITtdf5epLSxEzvB6wje1zdUClf055uycrTBW6WyO8KNU
wVsRMNUf3DFg7xivZrYutfGh6rHOTUinjym019ZnOyMhSU0GrflljqDG/6YM7TrB
KnRcBMLAolfmziP3B4AxiosWrK00hy1tmluYVqoKl74sXPSln9Jlyhl4qloiFFGT
2OkhFL9kfNbXcsNVyRZGXsh2+rgPZg34R3UXSh48VhqSnOWKDiOqA0VViFg6uG3H
iM5lraottK0W/fe/JRlS7Ea4vgMCmF5QRdT3pcfcUk8DmaHcQVpRzCOGzi92pWuC
unHmDWnNkuFK3EwmpIpy5xB5gnYwjBXnScKgk+FaCek0EFDMZSvj3NNOyR+WXvW+
g+xok/xy53wEOlibL19ZjzhyssISUGl1SPHmJS1faOMyvbSNx6eXMnyeryXHMOBF
1zP9ulWlMjlThx64Tq+7sHpbBQ90S+GMLiYFcPuUN9okK/v1zTrX1UJfNspjb8/Q
cgRp0+vuGUB8QmAW9Pc9Y7IKgMuClMIXRRc74RqlDlvSxgok302/H7iL1OFA/F59
IU4jdduOu45z02hZzmae7hKbbOGbSEFSr6xW6MzVHy5xgXFvje9uNUuZygn95DN3
/f2BMoUsBP5NHb1HePlBlWD6McIsSnLLB8rSfnvRakt6TfPsmrZoHt9oPUxW9YPF
3XtUe8ArN5RoURYWLZ0Vde/Y3AxxIezz8hRXusBlcZnC8la6Hwq+6KB8N2LVxW9c
d58TEofBUihCGkKRyt33ZP3kqEYTo2yhUHGfjJRG2NsQkC+iTiE++ueGTNPAtKZD
eK2izOZyja6K+B3CHulnW6eJ8otNCICZV3Sdi4LJL4UWtEaZmSgO6kAzCR4N7a9J
/kP33AXvjWJAL7o4gMxpAl59rYIxsQyVJcfo+LkZbKjzJOQwdM82MFJDxRjqQdNf
BCdCCS4GVp1QPkwYKpXSXkF67vjZrNtaUCL6N+r82f/M24WNqyhAmONHpfyv63B5
YYyDXrEk6lDev+KKv8BHQyugQnxXBSrNWmGLzGSEmUW6JVJOk572W12dkS4rBPIV
ClqHAZoROjsFiu7VA/g6kINkGZWH+BJZsW6B7s2kkZYsZgkTyJRV95vnTw3qOB5G
SvG3pVUPttrIlkmy1j20bdajvyWTfaSnILwZUln0I6+BO7K6GiZo4voQxzpVZvza
9Noo9urPDwSf0okc+mwpVsF0kpFJuqbzz6+RvEMzWtw6Htgn4x5Ydqx9K1TLiV7P
JAL2xw/tIJPGmJV4xFbkzoaxtFuQxOPgMYgin91EdwXB30RX4wmg/k6QbEzihLz4
kapf3m28JC/Xbd81zqULazOsuZBp3ae8yoi0McIgw0lcaGlJCh0g5k9aFIKUF5qX
jPluzRgveVGTcyd3Ce6fA6o+cITgOYOmuV8t6iikZ1fj1wrQo5SnG4PnXeHpF3mP
5C28/3zPj9//NRX1mlfY5sdPKY2r/Q5ccyQnCP6cLTmdO7isar8FjSW5GCSsJz/p
VZY/0O9h7ErJ9wbrCrMwDc1abGtB8wPMSUJmQe8yaZRG60AWXQCwD2LQsDXw5Mlp
fOZ7F1atK0EkLCKAilp2vLmhJE95DdPPLskJrsfhVVwlOBZ0TSZkQWEYuaH8Fvml
XHZo3vralyXbGLqYl7ociJ2NuKyhbBzMYe+LibXqMxmBCBwl3/aHwFCCB5kVOKYY
SFFLQ1RGmhn7sOyGGiS1clfUn3IeK5zWYexiQlTBjYKXxV1pI43nZLoFaCNOUYt+
XH4Wn5PbC3SBRG+hYGHs/he0w63wFGmDfpAshVgc36LVDMGKbwL9ivmPGT5z3y03
FgcwtsmULjCx8+kLG8sGHpLYW2UnT/ApatDfPbBVcQndVfI+AdKUsbUAeKnsXwGs
3q8F8lDJy2g3br3JACDsJDICUbPRlk0lgZw0i2IoMRECutH+hsZVx1oWqWqKTkHt
CdpRMnwQqm+vctWa8aSzD9zV9ebgLukzFLiZ+DnHSz1EHd9Rs3jPCf7zjshQMRmj
MuqafoowHk7LJCnIy0x2A/hEDSP/yshtuQu5lIwa1WAAG2C3g4OUyDE3pw6Ax3JO
izkw8t7Lo+6y7otdWGRBwtHKVKHvIg1nGoViiTIrLAckSd52DOXL2ov9BGDSkEfU
OKA8MlaBUZ0LbjOXhtGBl+4Xb5BpLYKvFngXNKr4YbULnd5o5Z91aX1eQYJhGn07
4YBkmifYfkHDDP0tQXk7Xl1FzScyhjS5dRyL/wWNWAhp0Br3BMpsXpe5R2fsoVCG
1Iytlkbr+cDUVv1TQv4Z1zqwLzQsIXJU8bkyW7E4ComyeF+nUIjmNR45iG/hxD2m
pSp8XRxEyL+6uNYf2nRF2+h2mX54jH+1/AAiYzewftrXJNClSolyQclePqNHg87u
+y7xLZ8u9wnZdyjC1UO9/MmwoGy9SkyVC/StHUMtgs3RsMpYMgh5+fdd9CIKygZ8
21TALhJ4uYdRoQ6vx7zAWAs5VATPqkWNhWaXYftAFzgcRrKx+qgiBmyZ/eTCOVnF
0Nx3CV8QxEansXXKOnnG1qZ/OavwYBnI9CrTWlwt0fha1S0bRY+d2VCUEeMlktIn
t+5+dUKzwQ1Z7PQYBZPLilQ+AIWj6hOZMGmYmHItYtn+8pJI8ZtVYdd/c0xSlxPn
TgiCmR1bEcy0kHuaFWheRx/FTkC/QkWf3zUvYD6EvA/JxNg+M5iBkzRPluI8pbuO
UG7jy7pgJ3nYyzmRG7bO8NnIxioJaqdPq90Q7v9LCBFmJrSuEsljn5NG2LJnnDb7
AN+hl0Er++vUoyqAKIDB51zS9DE/1dIbcRQ2d6JvexTLMu2Atp/GVvN3yXj4wPLg
+oP/FvxEzuLoyUff+FxY01AK/Md/U015/3Zpbn18IXMTc36E4ZJq5NQTR50esPzs
x3mHYWjCBuwSoRcisQruclBImec645K3hey3GDmvFbs4q4xbCyZAUPyKLtGAKqVS
LasMqVp+4J4AfEH0kVJU6rQSwN8Bj6GmkfeD0CS5aQRhhB7RpqRW1t5/w2Ic68++
ij2PJS9QN9SrqanNY/3fqCjoXQznmA67HYnpqlKUzPzeadRUKeR2MTVp5oiPbCWc
2pPGqyVIeHOrIxycb0EsM/qUTwz3TogdiZHbHiDO711QUvkjWflj2qmm9ngAIYj/
fLMTxFDxTk0RDHIc+QS5gDAtnmdtT4z7T7g5VIWAB2ycvnTOYQN0MTpBSUQtvz41
s8bb4rcjNTfQotveuCBOpE2RddyqchkMgW2me2hXBxUjT8vP/BOt7xmKDbC3/TCE
0CunAnkn+uA3TdX5+wa1E6KoYamxymFmn8eDa3obzicilltpHBbYqBjI+Jghi/1u
NzrAtgLcPgERQEvS9t/HRyuTQYgiGnZ4zzvuEpIPNW7L3Ooosf1b18u956/KKn3z
hYtCQkwYZoZl0yoDLIrg/Du3dv+gc6oJqkovBeKVsG9rlJYHwjQCwIFzCt0eaBwV
WNGPQO6idGZQWtYPXhTD1iJyP1tvGSmXZXWG4dIyD4ZHFhlCp/xXsxKgLohQnu7Y
HbgRCJmCT1/R4uSuh6ukMoOfcU23JMvg8Pt9zYBqBAvT00ANDt5J+v4d1vVRNaNa
mJxuq+0FUKgZwktZBLPE8ucj95zgvf6hfrbaUr4MGKFNv6hVpJgVUz0c49vKC+y9
1D/NHJitIUXJwaNARw2HVKM9gJ2vAeopNnmoV+fFNfDYqEHp9D9/EhniJq96PZes
OWGTDu7q7V8JpQOLqitKa6D8ztht82mlph3ZuKDS1NYhCIm0sPdwilVsx9TC276i
xhaxcYdTEkECikDmRYh5hyKeUuwdNhOnKNy4BbG9hVB7rCrXl3mtQlqGmObtBU9S
kzAxRUC1M1DnJtxocPY3ztQPgpJs3Uv5ZoAKojsPytnQOnT049e3ljtufnDE689E
lbEpSKHUDgcIsmYwQmZhgtQUbNkpnkB6vQ6AQLemiXo23XJ21O7O7oRir/yJirJn
Viv+RtLEM+y+dEgIZEyk54tE4R0kbbv6iwNocQnkUZXD3d6AxsjXuoA3pXdnCri0
eZaJYF0fWP+pmHSijbkhywAO3SEzkcfKk6UoHPZ7w33Mq+K8LEszJmnRI/pu2WW+
dee9GbtxShXfolgmE/BWuHyDnKuKEVXU0HI990YvCafTrmCl1BdfvGGws+8KAMba
nHWMfQRrPCLlBr3Ov57L3d/1NLoQyZo/jdZnYJbp838iuDdRzhyPnrtl65Px6wko
ImQaaF7+J/LUr/5pV+qzN0a6coY+p7iXiqUagwzQeeIznhnEqvpipgTY8BufOIoW
znUy7BWtWFkI87RtQVz3QxbJD+bVSrBuGRZsEPiBVB0EH8tf30FzeiQG6K5U+Qut
vQNen7Hfomj5uQ/A0noKdfxoVn7YrazUOTVjprBlV/Xzt+VC0Hmthy2/NfgP6qVJ
0JDcYQ1aJHaDotoFzeoLK2J7s4NgNxvgvmKLzOCwu0xryCVwASAfDCjSil432Og4
fQ3rUpNtg6GuaabhBJI3PXsPACCitTg2E4H1ScHwzDwuPkR+Vq4eYqQQZYXh/xJu
rdHU0EGN1YXdRJ1ypvtYOVm1M27kbwKPeJJxFpoohIWHnhKQIEGx6QAZu93lbO/A
WeVFrUDT5FrhYl404tJmgDuQvBlTVSOqlJ3kG58qyD8FBz3WLXjiDsjTbW5zOJw2
zVtDBwjjudLXxsGYIS1BohSNhfTJ82ho08ecerKEQOGG7mMJBQ1gIP+UDOi86zaK
0vRTpta4DG8OIweu1EszRA+cYEymXNv0U6iXz1jXGSHwx4l4rE7i7EnaLf1lSXgD
VZ2GU8JcyrUw9xOX9EHMczEpu99mo95W/Cz3CyQIa47XIOInEMSlFrmkcJQ0THRY
1Y+92Dl/lJoVY00FmLVbuDa4gaJwpQAz29DnWbRiLepRiadhuabOVT0O8INIbbwj
eYXVFUKFKFDDGZ/BC2HQ3eJxLnMAk8Gq+MWTfnEJaC0qumAKTatqmH3BTAm9a0Kn
8eLTKpqGaiSaupyH7pk1T5LT3bbki9SPpy13u45Nj0wQrqIpdbdzbkIkNQGA8UUe
z3XrvEgKMuKvk6daDu/N0Nh6t8n57CVBAshZb0Ha+YtMOBWnJtdGJNAAPpYa2TV8
GEOynqudfJ86voiZiUuSXg0/uIMNmXuSlEYofg6JBDrsoTQWRfujmJrR+tNfuaXQ
0s2E8Yc1MdNeX1LM8+bqmINzKV1EY8/8PBSK84w4eDbc6cHQqOCOhB0zMBwZeJzw
lLkdENs818UnoCAefXZpZWvIizhOrFqlZtO6+oJ+VYpPAu+6WR15WKFlC4hMy/rS
dYO+CrwgfgQaKf26BrW1vWaDVMZ7UkaX2/op2AOd+TkcouLVlYgAKKfapmaCJMF8
41yACyZc4wuLZ27YewT2tWxMqPbkLkv1TUuOafuju0m3FqvN6k8mX3xFTER8QlEr
dr6Kz0nbZ5XirZDxlYeDvxeuKhw+FpukkbRbNEs6CxiY2iFypg3v4vULZWryQYiW
p02WFT+0MgvPin9e8bYM/vM52ZbbrEJOoqkhfkz6hpVxixJt4LfEm8sU1T2g/lZp
XG/V1qCAnEYjtw9TylRUXof12nHUv6XSrq3SehgkQMWa/wx1gco1YqqWueyMxH94
HmnLlq0XrVkIWmmWHEwk6k0+8yotRH41AFBKrdy1AxjlE8j9OjzEevw0KaXk8YNc
0WTJbFPFxUR6yE3yw8upKw+Hsoy1E+KVcS6mjlx2+NXdpgqEXfzIeIeZdqG3DPAo
wSo/CqIxy2PySupwKSKQMO0wFXGfnlc4j4sp4L6s0pom/3nyBewCzxy2vHJTrHKU
Q/3GpI8bJx0weRAJqO3xNxXxbc94sWFTwn8RDSrzh221YW0jXpZSBOBVg1lA6pXB
k78A2opRqmeNE3rNMOkchsXPHcCI7rxqptK18smwxuh/C5zZE/r1h1y52VO5Zbja
D8pJ5KT6RbL/TCBNE4v+bT0SNm9b6uQ+LqH6/nu6XAStiRl0zQGhr252pxS3F4r2
RTa+h2kOJN7X0oXh4ixpcDJRXSOjX/d6hvI4XpBkFDt9pFbRMCWXcn6bYEb107Gp
tCCYE/HtNt51rHAkDxKL172oSzjyXHTwEYQcLAH9vxyRWIitjekMy+LHx14Zy4mi
NlbtQ+Ed3uuSqqzfO0KCS4QS4sMvVCh38f7ydoUw+fQZ9l/KG/z1XLpENx4Mgihe
fX68v38iLqtCv7hvHZir7HkXnNb29DYJi5Hh7XBZ3KkVIGVg36KXfRyIZ5hCfJOt
k4sAxhd+XTmhcNpOZLqqymMsjoW2XN7GaAPKsf714yV4FbTbqRq31+qtNSMXnlhY
bAVl89CJoUF9Zz4Hx88ZYZ7VBiBg+h6EQkPS+m2nmlzu2/vTCcv6pQ4CBXW+lhum
GymKtl3D3JKWJpT/mOoXmFoqrkeKOODG+BEBSmS7UsCW20I/+Bmr2Z7rNzzunpJn
QCqwi/Ku5iTZcaV063URU59ScT17ODY4DjXvVIByHBOatl1o6JBZPn8Hj6k8VBPu
EFRBUFMEXVeYlRLyfFqw3Mum0ILYzICIDBoIHxPUczUnEgOnOqZYqeWMOuU0Pa/O
qfex7wiuPagEFlGUNbvujM6wLCSGzIP6qjNhhWdTUpObJ8LcNUhLtHVhWDacGEba
yx0F8Ker0XZJYTi6mkiN8D57MwUW0HqsxvD8hn9PzCA8e84xjk5GWqPvaYbHpVTJ
4IJ7aKf0jFpPqiOopzzNBfomuvTWeNqqts6xku8PihbPeS7+No1ezWlwqTO0Ze4s
jBu8lY7eMdFMI+L1gqfRrkf/fTw9fjJx1i1LqiEoGM0WYHl9Ntu+rqPSefwDlkVh
Df+t2muSAMNpIzwlIrhBxqHPSwASadTktyWSKW4qSjgGHLPJaU9CDzgMuXVnXZGz
65Oj7lCaGgj9zbGWd4P57GKj1JktlheeboEEVgA3p6xJjv0x2SVSE2/YuBDJSTMo
I3wQjpcwtpLl0ndrCPJdzCL0UvWoRX5uYk3nCTTAYVo1qSLKQsefXI7RgAtu7gLU
kP3N4TA5RG1yFfvxM087vd4lstDlFtFgvMPO3xixESXpOx4sfxjRoQuoyVBQbqza
zxudwOwu+M5bwdZZQMFfjCjQ5F41Q5qaK9lBbKHhBdE90HAxn1AgiIOME6OXrd8T
NbHlJ1u9M/dtwbufQEQB8ZRKWjkoD0hl58+k7wxpmcZctCQ86H/7G0+7nrGGTeY7
UuScjROsaR98xwrCMUQveW49eYXsKH90taZV519yxDooXPs0jIor+G/Aw+zVtQXO
H0ZLLMPgLj9x/u1nb+8mD8XdAbSxoHFDJksqLi+eqUBS0mRnhvwjV07yIWTSZJC3
d8YyFj2JkQ2kgB7C66DGr6jtCSsuRAcjnqo+wv3qEmmXQSd2eCsHqWqXiGKauF9B
Fs+RHjy0vlbX027moaSak+8cjczQRwRP1wv/YZo/FszJf1kuOHdI1xq5dWk7HJhA
jEzFy4vBIX8KWbX/xUkhuN/J6A2NMlK3RX+3cpk1pfr7aLq+WSm6fOTIXUMigu5M
U/JOrgUajSE2KIHhLyj2iq/DKxJotZgXj5Fho8jMErBvAtORAJjKfi1/t9+mPsFK
qYyv/uw+GHUgOSofjqSFc9W/4h6aMOS/51y4AZGQ2s2VSzW3q/u05WCRRETgaZuR
RU8bscp7VdC17aojxlCTedF1gkiYsTx4rOEMsjYbTHGcDP5B1zuOoAaCZpwn2mEZ
ulRUy/Aqu9DaD9LJkEXJerF9lraykmaNSGx4sxOwzo/VLf5CB2Y8TvwlN7axmE+H
csq63ykKvnok+h/5AHZvRJ1CKUUsjSc1CdKRjSmtu+RogZW2QedtMt8PoFJ/f/R+
cLbdJbQXilGBL3n+1eXtJnxIHFW7P7ykNzeW3hPNbwzPDWFMRK2+ltMYqKhiPVje
A212HR84EhZ0ixvO5BRZjLAaw5QDQNCkFEV0oWRzmrSBjvFy/LPteZ4J58FouwUw
GJk/Oj1Ck8AB1VU2ILg8uCbSY5BKuhegyix2Rml+p6Ca6yINRMKvG1cub+C9CT7O
GLiDZEK1yoU3XKk6V5KGdZz3bZgkhr4GeC/km8zWcrv0qRPmEPPmlLIsvGBav77a
ZP9IPlgue2nNkJFlYF2wT0fn1NZgcVetWulv6E40q06SYI6gRhkjSYfi+9FYOKCl
0MYxpvGsT7vVpq7euyUNU1n02q/dygWb/Bo93a+M35mIdNEJ5uaY1RKiTdTn8nj9
AZn7jmYuOdC4ASdkxYqfTOGcbMMVrbaVxrRIkeN9WkOZU6i6bI6xqT3G0w1dyFPI
tqqbklG72K7n8nuHi64dqTdcxMc89wjG9PmOMbaWJL1UM08shi64+F84Uepj6Bsf
cN4l+p8JuhfSrRC2EQSD9PS/vwVOnOF38ZwVFvtWL23sCl3/wOoc7y5UnZwojjFO
gIBV7tbd9UtiDWFM1BMhTNcnuFpcfw2mIL2m1sH6nBGalNyHmn3Q5NrbDeWWi+bs
pWu8A2OstNJ6JMBFTbEk5Qz+nSNBa1klFpu1ckTFE0i6McR2L1CzrutoF/40FAAV
bQg9RBqgeCZ9Tlfh2tkwpetZ3d4q4ACm4eyJSB39Xj8+UEwODVS4dNl+BmwFzsnr
On/QDamFZUvYXLD36s8EKWUziy2PcGVJchQnDAgW+4AcoUjmGA7dnRyu3S1isFw5
3VUQ4GSSO9AC+ILENusuK517OalO4f7kyq30ieHMnCORTl8Uut1SbozAAiWHBpkk
UYO8z//JekRy//IwJ0tdAnu9E8BtG8+SqFghMoIeKVD5/Kde0h8uqQMrttI5sPlb
7FJcOnCPBEhdwY9lfMlaBFwZLmaKBYK5hE8ZoImy2XPscHDKcERTrSoSLcHIhkpE
0lLUSGgoRY7kBa3i+krFIeGUAhjEuX99N2chNNUoLbVUWo/9fpfwOYeY3cnh/ER4
QBYbYnnc7IWVJzu7GpsgOB3aKHqH2nD0Ry6/FWexE6PggRpSzG+uPz8hk//7xiTO
MMAjEAmD10AUIcLauGXy0Twl4H/LfDPWVe8MjYboRHXKJ5D7xT6vW1VqJTnMsUip
mixMRkKrxG7Z3l20Jm2cmp/6/bhVJtdn9tRQidpYUnc/5aUpZukWmsiBtyQysbxH
SU6go6B2OoeMZ8+kemz00H9ynBTHiBm0qlJYnE1blJupJvL7S3VbF9Qz8k/lGl5Y
RXyClTXjcyaYTmqgVrvQ9tKcV5O3GoH4ybxsdK/GxWj2Si0v0PVc4J9iu3NNs0IG
D1HF+PI0tPkjwolJ1CXyTYccoCGV+ByVuPeBvM4c4oN9knWt+29aCuR5QISS+5fN
alBSM5eZiJ67ise2RQG7Ors7VVkECtL5ZmPlt/dnL2fLX1+UFtBHDs14D1mEaDYW
PuQIsbm4ashNWIUYsMq8jxu8h9++NpozE3PLrtWYx4oznjgQKA3jnaGErtbY8Ti7
zw9M8S2XmZpkbGe2wjudoO5Qo3vY8uBtLh1Gu6B+IQet8stK0J4JVd6GGbOGjlPB
4NeYEtHOowVOMSCKPDtCwRsCtIfpRbNNslxfjGtkcBfFE8OKfV9dZLhYidn8vZfp
e0PZP/GDS8PGJNTIMGSY9fAKmZo9u1RNoccMPNXjkJd2ew+Dx4LudK4Os1YBy/G+
el1wDMdEgXw0VCuBdvxwrB1pRGFxr5iF1G5H8E9H7ScOaDqsoqCgh2dAHMMB3rHl
e1Jc/JrkQL/Sty5OveOtg1cpUixiaEqcANVw8YOgNz/YtAUEgb2xKXIcM8bfqJ4r
FfcWsRYauAbUNKhs80VJJIrUNuYkK6dx8SL5bVU/Ci5kmWyLC4tOVpNACVRM0mi1
rzjD+UjgFsSyQpYipE9THajZZbzoGcR3bCoMsrMkdfB5iFDJ9d71yr0CWVIXx9fD
xb38xcAGCNgUdgTApQSxF+mO8jqpp3LjBcbmiL5Fplprxn/0tFCf3RGguOJPBY8O
R2awP6iYa94hKbxrtsafDbJeUHkBO8bdizpHluOTvsafjlyiL+TcmsmZk/mVguf/
dGBGosP5mRBHJP5EXS6b1isxDLiPaYjog+PlshZh0vGR10q4sCNvLDr2lFDq7kSp
wCDQfhwi9IX6ufsW06RphRA6TMh4x3wWDZXRSLtquFjX42HtGuedWUi6KbOgavtY
QMypMMYep8CJ675gsbRy8wH+FlUttCFtORvTr/CChdfCMI0yfqrHs9eLevhmniew
xqNgt0/iFzJ3FAGLqu9UZFL26X1NYq6pH6zK0qiNLEF5YkELGDG3LFYYxAgyhBCe
fiibEIMZLiTMetYbIhLJK0UKGGVYvyh7AYBJKmuR4kW3i12AxmMN2tXUcCrIVppM
FZrzFD/ThH4VwIPLSt7sraTQdXyeJHojWEzdE5Mkkr+/05xtbEPL+fe7a1jGwhhg
EU1iepVLR/u9BlBVe1VhyC1gGK6y0BRBBtd5fh6bUfbPP+FmjP3nv1Agbl6B5Aqx
iIGadXtkfDHcLwkFA+Fc+8RQi7VNZdvLEYp7MV/2KmFRqCTQTl70RgV16CAPcXj1
8F4nStsQf8l1uB/FNdrTParWGno/+8YCH8dlMTZANgA75mOxz82yA/dvSVR3Je7j
iKG7tk0tGw44g0bAPQwooauRtSnygg52rm8NI31FAqERN23OFPyjo1Dss9QI39Ma
QMCTTXmBUxoGc3JDR7+EyRTprGS/M6+T45CSjJqZPbcDSryXX3tLn9ZpfDqpJQ8X
QLIBZ8RHWZQQDC5bbabSkglROLM13r1uJ14J+zFsTmOWotk/F7RgrMH3hwjlet6F
l3mPe9R6wV4l4iaQmuPZIF64ZMYFO+7nrm/9Yw8m6hl1YLtBZGCSEPGJZx6cfp/Z
2UltqxSaEErQH8HauGW2/Pascvb/xfHUJezrTczaUhZZ6d42wR2Q7kiCAFbLjWZR
YAq5wtnGVCsocqJbqp6mwq5kt7fznghTs/aKbWKDb6rgtzBoWJSqCZFvQVF6oMRO
/Sxko4muzX1b9z0QX8xfvV6WUh9nmokPow6UoRCOq3aVnjRCkjQpPE1pkuuWBIhm
eO2etnGvifrbBXsjOxYnMXWsPPgpDHVSRhQvNmqRok6Y/cu4PsbLOLEcS1wuRkxT
ENRuUgA4Lv4+5sTQsISBhTseVfPtUxnXsN7aCFHDvSm3uKzQqXraGuK0BNc4pX9F
bAlXgOOzErIgJrP4hPm8R8u5SXRMJGMPd4i43cUuxA2X4LpfK979jfqfGiYaPiKa
yuXVYLL6CpBFyVNKwcjBjz/dPJwxOIXzp2mmTFt4qQnAIsx8BYQY++WEIPux03ln
mfXd1UVV0XNHP9fbqar59TEmbKulJnqWXJO4khQhmq/oPEQkhFHtiTdM4d608nWc
DL+Vr5XS6ZSGtDjrBBAITEKlWHytS+viZNs4aU57bg/a1c468SPKRwxfP3oz9QYN
hs7n82K2ViJ29KHCa6ASGAqtfmleFaLXGg4WslW8UQvN8RApbOC8R5IBtEf37Kuh
xWNaKwrMMumD+a74yGRc1DAOBTMN7K+eD/wIlNw6x/9cwiv75dyZFD2Clr7MBym+
xOE3MxVrZ7KsOdd/ePaDpuRx68TfMt7MdVnkDOFK5dNl0i4upy1DBDFdlQOIe0jJ
J0pGQYFLqJaDU9YoLDkrhNt40N/bfZgwU+/2+jiUlC/BkfjUG6S1f+e3a2ID33ic
6t5X0i5tFEjaJSenCV5bt5xGqOVJuah40HdMyth/0TmcGw/0r0t7EHVU5aaC4+hr
HQ8W/5Uri1/m3tSLjHIrjSyMogyeYVGzAiY4U9wVHkoe7CcCo0iAVQY0J6+Fu/pN
9BlFZpvZ2M99mEIKvWgd2pmsIIexlKhY1rOrQl63uJ+S84zswRGPDK3VmJi9jwC4
HCoNRQaJScljBs7kv5a5NGChqop8fhYaco54QdqgqiYDgHqX73yjHVtKsZKsA7fJ
L+YYwmftSMTbrdDaiFR3OMQGkCjlKUXOZyOLfqVXvXiaEBsmANnA6lyG9lAJTWHH
NyE6J1DTmp8fq5ftOvP5h60axukS57I7uV1jafrrGJaD98UXtcdT2z8GLxtF8o7W
RyBHv/E1w5f9AJpre6rxhEBGyBO2HXF4mfoRRRGHrSiznqmGuChFo4U2cIqD9zfs
sDZEgHhtIhkUl+L9E8sPPcpUlKlxDgSLeLboY2LVOGf8USSUDPppDp7Eq7G/gWfq
z/cFjtuXY/8RHuHlXQHGUeYS31QRQ1DV/O1gMCqI6az2a71HH6khxMfAjsHKPC3K
1ZOVjPy1FOEhsUCJR4Rtao2qI/1KhXXAekjHTXIjy8/CNMXYmudUNBEHTglER2EI
N1i5NkqeSpPToxJe2qJ8+eHbRJJS07R68RL3cpl3XapdLp1HQ9gAzfWGqWeGiLxB
EDscNZcvNme7hXenx9BeTLHdvqdqAFiwe6Fe4quw8byVJL7PqNPFnn4Hro3ZgSAr
vcKevw7F0HAaMkv8iiHKWuQmCDIDzwIlO47saZrsul+kYZpMka6ICBRPVilkYFUs
hEM4Nnt4pamCDYyuH7wLKk5zRcjRM46P1mdbsHh0iyFRXPyZDFdrmxk9Lrp/xE7S
H1UYVRAcLIdto0kcM4yU3w0yAq37II1aNPOWxtyHxjKNAe+QSiMYx+5Xw0m7WFmj
K5pddWHDIromu7q/kd93IELTnMeykq3ylgRcOdXMH6+Ose1XPK0J1QHlFuFXlY+R
2+fXKXPH4P66GH+/yJkqseIabxm/rAMZxGjRdRjA5Z/1HlGsfJoTx5HX8lzFgHIk
ntV2qN+I2SjbNhlGh8sqSaWOCzNCbWopzslh+Bwr9WXLfb80yXbhgcY9LBC6dYmM
VGOfJwUDH4M5uT5whv8JZF6X7p7G3/yhkw1JAoiYpNRX6CD1R/TRoRqcbOOHlRHr
uqxy2cTEXKj9J/Q7zSgEJFsQVHE/3xHjgXs+5zaiM3Govqb0+zanXzVXHjpZc9+L
GwIqqH13rjZJaDN1oZD1B6v4yH8f1Uq5uh7KR7H78tvNWcXR7u6v4F2yqa547C9T
lQUDjObSpTQUwzsqsppvTW3f485YztawSPC8pjz2Sv1MkkTL4LCnHIBYCaq/4N+f
enhPO5geBmPnIQOX7X+HwWAIBVO6AJWnQhsb0TnwSkB1mqDLfMuGyVcUcNiWO+8S
dOVzmwvMCr9YqvQ2qmQGS8wn0ee7IdlpvZPk8/HK5HpNrjQ25c0ay3PND2lCNNkz
/wWkWYoKbfuhRyx6eNEDRSqLGyS9DgddGmRbuFhT76hFGyXRH2SoGRNct9lCQo/e
tMBB908u7RpphP0arhFimdOLMrWhzUn0Pj00wl1cipNYfaU5vtgq1p+e5AhjwXh6
vZVD4bD1FpZ4tgv9GsG/uibAc8RZB+3WsuNgiLdK/24EyjTZhcWnAcImosuMLza/
KYsvT3lRqnwCgVo5UCUPT7sUsV1P9Mq+L6tdxtSayU52Ji58rEBfeI34e0aCrJbu
wQ1rT2lAYKAZmoo14LoESiaFkJ4AJErBBzC6yGA5Y1jnO3+WBvuRo7QGyjGUpqmd
jxAByldls+N+0M33H6cmSPZrJYFsni+dl/yyrQmLiClE89xMxxPUwBM1bHnCSsq1
TjXMWT1eHnzCtUqSoREO+fW6zNrdgqP/+6UIKdIQf4IUE6VWiwxjz9mHw0ZsDzZQ
vqJuNPrSnLH7+TcAdJB/a29LoTY4ptJd3b4xdWgI2LG4eCHTrP5R59sS6rfVOkcU
Oj3ELMTY1gs741u6flFBIr1likz5YtLbhMaOTRWK6cdC2yoH/thgT/8qsnPp+k1u
OQWd2bF1PAb4ldl0rWXaz6Fm6kMZozQyt9zCs4dooMeInzU5KOsyxE4wxt4WD0zM
Jm7ZgvGBXNmYGfFj1rQEkR6CfrxTOfjgHPv4ExwnFC9xOAfGnCI1pYQxFgnT7xxa
VsHpDe0um1Pzl9hHhOeA3AeoDKday4BiYeGaW5kAtQHU1L8bINNYF3BGPF3L4cyR
g/XqX9b0C0KaksmMQzyyZ6EYbZ6vuMYSDxcLjOPkx7ZAPZzsRGhr0GxP6kwO3pnW
UfnAuQRCwgJNe6gc74LB0F5g+EfZtmxSg5ThJCtT0ZTuWIL7m3VzNALIyvBmLzw4
c9X44+r7PX3T6BIndP/LsZZbu0jtxuCG/blHMrxyNg63jtJ8M2h9iWt9CWMAB36Z
cSQVcCAY56Xq5dK93lu8BPb7bsLtVTd0KXziCoAmZEeCK1yYSjtQFvKe5S1b1Bjh
ZBSFOa+Ud8bIzdFRK1U8joFp86i7IKJA9cITZ2ewu4GuhzJK5NtWYJVmUtA6TQpa
EZwsI5HwXmVT5Elleakk2JiIh8CYo77kAfDy2S87w6mmepKHr+RcQfB49B/dUPt6
T5xUhPqiz4DB2TpS5Dn3oo/OE0gHPUy+HuQIeRyRkvmGb1d8DxSON5s+6Ul2spXh
dd0csr6y10DUQEcvQIeNlQs98Scg7VD6oB5nZDmiAoa/0rVN4Vi9yjScldJCyjAs
uJHkJItrCu5yQqCfUJD7j9Q8sC4DFR9Mj4oOF2cUGtWEnX2ztu1aaSXDZ5R6oYhE
jeAI3RBmoeU+jgfbipV83CLuaXxFpWNSHVYb/8SJAVwG3tYqHDR1KigtQpn+xzp3
kgELtZM9fUoy0/bNX43PCrfp4CU9Hw0fBkaEGEliX2WZTeNxOxRVxhQtu0QpwK77
oiCn0g1WrA60Dj2JByfQbCK9jG+xUQrJkitYVeMN1Txvk9SLlSPVNRPEPg2voQzK
srYa5k/C7KrOFlo1JCqh1Sz5w/jS0C8faz+IzpqQfc1YlrzkGCOmEcfP651k9euK
fp72ew7IxJJk/tY7tkZSs03ARLS+eR3ncC5vFM6VoQxQLvUBfrSQp3VpYp1/5BMo
D3er7jXtarOGC8xLKPksymQ8YAs2v8qiMvNrE7zsuJSqJ/yoOojsssu4hWS75ym2
218t/bwthz8B99AhhsGguSAByRYq5wszkfwMbw3ORMJzP+5nlp6jni4dX0mnJNj2
Et483N+ebh91K72GyDyWaQePMgainQ26d//rj4OhIuHOfy6gGdjnDpyPJEM5QfHi
pChXD64lX0R2QCm3egbE/R1XRgqHkKsuk+vJPsehiB8JfKNM5VBkyLelx+6I9H8d
7cNE9hQu9cIvvImR9tKPZrUkxRS+wcD5UY3TqHXP5fPDqWism9Bd9jk+dTnWrFdN
zTUZUub23BQeAvT0aj+VU4sSJz95QrNClWfYr8fZZ/REaJlx+k7fCQ0/vW7u0i+T
qbEFUpMJGJOz2Tz/o9HwzcpC5yU84u8Z/TA7UG0wmga5B6jvtFmGqKHFAY8PpUOH
Iz1ghFekz0S2p/TfhAhAjmAxqQThNnMg9W4yDJeElzOg+7yehKEkW22TruOsatuE
XHb1ObQoxk8K4Uvbc2IY5C2PYuwRhGMGogVCbnJJJOpGybtu427lYJvEh7YtguCj
YDcwOqrqU+4tFriKtRCRDpjAoFvdCD52yJv7fwgxd/5c8cJi/5YVJ+10NVjWrWMS
ojczWfwiQAonuFB5CaLImJt0m4YbqErHggjVyjOSU8/RS0Cq1qofq9PIzuHcfg1x
6B2yPw7VjnSiWwtjbxGLJw+ROYQNXYv5ZYqkSNCa5bUUvojNlGmXIbGtmVqdl6jv
UB05f3TkyPi7Ct2ALbW5T4IKS+VoUkfDKIIOcUGmnrYBCA58VR2zYReizusgFbwE
XWgJfH7e5H413U2tA5MShnB6d9fYu8GU4YvZaXOkjGY6aH9YiMPJLNbEIp/dJr15
+5j+Jxu/pN1tnn7hPofH119gYaIsM6jV1QvmOhslzjlK5gsp+dFboAxQnethQd00
IUwOliKXezjx62OpeheRQSP01ZFTHThfLo9GC3FKfzOFlu0HBNCWtW88zYpqfllT
DCCSwtK3oXnOXdJiCeWYGAKahGNGxKrer5YijDf73bJPlccwQOotHBqBe3kMrUd3
7hfWI++NY/lV3Z6L6PGwC02PUzUO3NfI/KI/kzxaekaexMtPLIidm7xKK9/QZP5o
/N08a3qrdhzCpqxtG+eAr4FZ26Tgs3YpGTEYXDVhHDb1UI2W90l0gys9/oI2yx13
gxmwabDIZGSjN3aXxLGowH4rpvY4xlL/ljCfvjYEmfGWmlQt9zFmfeduyEyxM2IT
myfMVWsxpLmOv7DgpOa+Ttb7dlTwYfphjng7Nfv8+D5GvOpWGHSsPyjhIidnuPpA
NVfkI0aCMF6bIXfc7OwbsAIkA1AhfSSjc2jA30TKFx0vCERGWsdogRTqIdTh3o20
rmFn213QWFK6d8yQ2m85FSrlBx/rj0A8sCHveANiZI51RluVm42uGEUnOQ4+K+Vt
oEOSHHVa9rGlWVT6Qfjz+bWAnp6epYdGGrGrIEaIlKSutMpYGz2a3K7ZFnbw/z5I
bAenb3PYCtibzI0KHhQSDNa7RWN+DoFxjd9Ya8Gw9H79DATaEPCMP80kfAgE2vJg
SBSRSbpIzvBNRTpDP5P4Ldvm5rd9XmrR95sDuvjc58+jIDvDNSSz0bHGCdPXLquw
rQbfV4NpU8ubh5Ve1LD5OURAeZMtjT+mDZLiH2U+8fuRGg7GneqxAUFjHsgbApzM
o4gaZJVbL4SwUqIXQn0/bzk1+1Cz8mOHKxy+kXbeqkgYNOg3M+q2JWwccplXpa5U
kt2+TC4TQYM1Nb2insWcZkGrLzO8GEpToD5HIKhLf+z+poE1dvRMkl6WndcrYUSn
vFMk67oC6nJfvZeQAFEW1tGRUUTRCB5YgJKdiPs+RlIhasKjGgtXFAqc6Xulg34/
otR3hStUK4S4aAkw962djwdmspWolmQe+ylZvsI62eePtMx8dfE+J++2a16iH7tV
9lenz0SIyFt2zD2qvIuh4HLVSCzCbRaLjecSPdIlfNMewfSa0e5zdtb9Dw6e6rY3
mCMdMDr/eQrepTWcTOGqKFw7bnf+hjNtObE1CyJsCG4LLSON89TyBCG8pdEM4ETX
V0qtTBEl1hAsvXzzaed9lmWtEUddz+blF3sQLinG2Dcbwe9mas6izEdmNVuQaK5D
fjZM3qyyFKs2OTH7OmGrTP3oVlWenROlakC9l5laVTQ1pwegF8AuKead+75Rz9t5
seeleZQjzPmvsAYPz34Ou1dKZwPwaJ545xgB11tkKzBSnRVFwL2re9WUwUhurbfC
P6VkX3mGMp/KdaxDWIpbmC131doRkIV7R0AUCiEfPm4tFtMplloLRHnGg2AJD3Kh
JjjfwyBS8qR+cWvQNAQL9SkqxmcWF8RwHJOMg4mQ/UvMjWBl7yiFxwd2HqJDX+/o
f9iP29we2Rn27PlpSoUQdMwH3zqpOxSrgREhDIJPknzqbq/3CaQrSxERKCDe0/ub
IHoNpzFXh+P0cyRclcVd8xKosGxMbUbXwzSb4gVlkshdmXbsbSn9cTMpjnD514Yq
66+HaVWkVNMcIzbdPRak5n20w8/HiRF2IuVRduKLdSa0ryh01nfk6u8xzEkVyyO5
BSVIu7nTWT4WbGzPr2vOQ/OWO0V+t+9mHkld8Yu8lavDN/0w0Rq1xOfp//PEqRI4
xdABw5+GTd61aOGG2aqC5kTemgZKSqWtYLQwmcUnhBFri/FtTGsftU/ggysKsFFo
CqSA4FiRd87aqxQBA8EZjBObtNe8RkYv/1V96ebf0A8npLnKrU8DAk3f/KyZ77wa
cpMmdIkgFIIPdUNVJwPoFbtnZGsH3dCkWrDLpVhcJAZ1tuFeK+P37Nxs9XT2Wv4C
MvTRnvZ4Jj30t7W0BulIY7ooc0mHc41vkQrIu6Q96YXlSVPrkHW/4cttKA+VSitT
xtP2D4r50zaFQaFHK9rde8hYYx+dwVNLndov6ORlQIzu0WImpmZpylRYgfT1pCu3
WvyLhTfDNGbvGIEyxN8HrKGaU/U8OOok5m6wlzA12iNyoya1KFWQ322X9u/Ee/op
Pe2rS4MFsiYVMtzL0oBlkK2tqp4KBizDfQ9xXGtWVm73lBl+I2vIJ3mb4+JmPSUI
C/dDa2ZFNEG2DSrqo3bg/j6gd3eBKAMarttM7b3M38U8wDutyLMUgTUxNWdI67r1
QtKFs2LyZE7Izg7wlbnmxr7dvemx7K1DqFmuxbbK9SujZXjT/uStkuGIWLEEPaFA
ytBiBv3qe0fd7OxyY58lU+tyvtqaFx5PSG0pFe8luYoa6mu9bJccrp1ZbwpKBked
jLiNOUkGYty4ECkvpzEtDqKzH1lrYqJf6u2TSlWmcwzuU+XCbuw3CXT/0B3jislp
JIv5ss+Tbz4WLAPmxlNgyGvIOflEG3VYv6z3+tZGDtZOCVa+NWHnXMO9WAOPcT/l
OFcjyf5N49ppa3xpSwYEsV50DXWxsVqFLYVMOOzi4s0upheuSfkRvmw3398Z7uHS
nB/hEOKsY4lTZtWzZKv2RTok23IygNXr/D0tjRiiuJFf4VuruB2AOF9UMLpTZCev
tCfKsZ49Q62rR7PQ3syV3odGXJmX6ZZRc9GZpQOOq0JBGdHT2eOp5NrDNbqavFSd
mYhJy4JSq/qlFHuzhmbphtIwapbapt7tkSY0/C15yzszGPmLvslUiUbG0fwb7N84
gyhkv0Dl/VL9Y5ekn/b6d7F8tc0VkbEobX1daMNmWY3+fnM0NfYS9bxUXfanDGGW
gEWf4q3ujg1AakpJzmFhEezATf8Mvr9ca0zNB+GeXbIMu5ozvRaaWIsStVE8mLKc
8PPFktAoJnbb6DCdkK/aQDvFMpcNgoelvatJxY18a1SHcuNMtUowBKXQrP+pc1WI
dcHsPjlajMekm7dGgaW9tBG1H/vBl56bXP3rF5dF8lCBGCZRLtGK4mm/cI1KEjwG
KK7sfkFRtsxcogb7WVxOa/hUAr0Nsl6jHpugrRlFN26lwNK8PtYouF0cAr8qGBzB
+NUUjFQJjtPJB/eLUrcQJLBg0gy/L7RljqvEFmft46234kXdiDI+Vc8mFnd32YU0
ISUSlFYOyBEjf+dGtgJ8Qn7EUjFf2WZU1F/KljYKDlbV6EVcXM08g+LiLaXfqLPO
Rq8LJVyBOEoB6Q9pAz8YFbxZdmDLFkfVm8WtxsJm/d+C5e0gwo+sVCzgqFML1WUO
tpEs3XiVsErNKlmM5X55lp9ffVI701qzsS8JPLearUNwjn/N7iHYKLGTSSqkXp1B
4ha7UD4vVeWjzFOTgGBmDWDbgDz0rxZD/OTciS8JpE+CcUeE1lEGU1wfc6hky1/k
FDQvWOmXdACZpcW34alG/OxwxfjPFXrpfnulJliEu58jpVsFTXFvQcK4LfUei8h3
fiIAcAkutYRnC8Qx2Rv8SOFbGPyVPnDlAgtpdpxxvwINLiLEtUy1FpyKMkYIdLth
7dpIScMGytfNLIuRLarRcoGSHv9hA9p0WQ/odDMoJti9I2gRIEi93n3GxTjPWx/h
3yRqnBnJRxOPTd0TX/7u6LseigtLjqXRyxOOB8bWLMA0rTPZfKI/4ZknRvmeIEZo
OoSubsbjrZxIesV9qzu2V4QinfInLHFirjG5+K7dNnNoSzF1ATgDcbCUUNn7pHMB
PBwNVyaAmYz+0E/5f+G9N5egnkfXyWvPAgsvebfxEVu/rXWshSHgSeZYQKzWeWbj
7YHNu3BP15Dr38Rx17+fb2IawWFv0ua5amXEjiQM8EuixyY4HZkIxX4WV0Iwptrh
2Um+7YgHpFfyJx0wyXRc9CMsTv6S2/T8JSgJvqR+v+bjAyxaekpPl+NuftxgMjwx
P3z4U0eqM8MgIhkv3FafyX6cAkBV0Haom6sNVTb8EBbeOQokkU5cpp66XpiPiK9z
ZblbXkmI5AAEFwy125R4OMsRaH5PcUwz5oE1EceFo1m4BsR7NmOIpMkZ/0Bb5F0r
HXd4ylNjowLi0dmvcOP9AV64au70+fkdzyhu2xPdhInTl+kvQPuQc8H91rM2SpKe
zlUGoJA85o0L8vBNduxH2Gd3v5E7iSBDiR6wHFaPuEfF8v6j8ck+Ql2JrcKfREaw
lXwp0UV2P/RWDMAk98k7RKlD9iJMnWEDAG6zBiGohmbUDehepsta0FfedUxq642X
EkdN1o8GQ4wpr4GBPsXP/Z0/kbr44enamGADCcdVrQjgXtK5cLS8+mad3YqT4dEY
m6HoCFk5Zsouv7JzmwIi4x1houa+Lg74ibwW5jo/HwoOgy0IVyVrvgZaGWkhV6UC
R+jKhf7h+kRATidfC+59Wgp3x3hz1kKeljrzcqDt17vzx+09LpyIYItZK5LojBRQ
vw6WptRhAoNG4+fYe39qgfKXAq30njJ17ou/qNRkXN2sO9LVoGdI0ZwEq75MPU2I
yzpnj/VazQRpaQW9Se8npT2Rnog8UkhBcU/byweDJwiZGBTYE4nKJcCcVYEiB9Pu
0bGhypnUVDqrfnFtiM7a4UnN4surmWQ2GwI6iEkfa+8llhYdqcOlgzMI4AxLnK4j
qM0OMQD+JURdGXCkmqPZnIzNsPWnrEa1ZM/8OKWzEaZ0KG00bPeSnEkBN2PIWKot
/WMG0jbGCo6G2+ZpYDdNhk0q8FW0Y34yTzqY9Vt88gX7E5A1JnafM3NJ3oJAmsFh
sEIvRvyoJJKgFpKRJZnuUVFHo6YLRSZ1FOCWNvsmrlKJYXi7ZHXLnmSujOB9oWBT
rmmOt34QdKHpmEh8vl/dyFRDN5nPmu94IYmdgDf7HQwUaLjLnEap25AY+trlmsRs
emSnyMuGQgMSIWfg85MiQ7i1mE5ObaJAvTMaumKMXewcKEvpuFc3Qdvi25D1wLGB
GSsZmyjdoDH2dzaIeWYkBvIYS7+09B0JgmArjW3VYK4N+ABTAC+nGGWU1chbgdT7
+LZmqzLNYShH2SN1PK7xQ4z+dt8HY6Hn9mOCWM0N0XIR2mPkWhZsoM8cmmGLn0jh
LrYVWH1HchOzou3An2/D4a60h8B3i2XjElYpHu6XfGoILz8FCNXWaQIsHgScA0zQ
1r0xPL0+ipwr5cOfQyu4r6jnYSCIj+HLcz1na8tYSWEQKEdeHl8SXYvgJYS+gtEb
fYnANjZcKyPZXCOiO7yVIQeGqtxKV42Ao6VC1QRHc86JG+UnFIUl9owsHaZ0hCUn
TWVrlRB/eeY2rqW/yss0Nz9cgaHlCX9T4082M0EsmiSDPMK6UYXCwpx3bvaNuQBT
F4oF7MFdgD+cvz4eewZOWW8v3rPAq5iZB/Kz+sbqWt+uYUJkFZmciKC6N2j3RdvQ
XGeHnSACnguAoYyFlRdD8+6ZMbZy4BtDczzCECI1wkEqGWjQBrSOZH8lfempiKzh
JOGx+2XtmjLcY8xVWCiYHKlvKB5UNBfaif3ciLS9ACnl12TGXT30PWeD1lZuAfig
58YW6mTspQl/Fjp7gDN1SbztFllFLQc9SpnDDAkZmABJF32VcdXIa1fHAs9j4rkE
+cYwgbveOUDP7dvwh372rg05VLtRPl8zxTucVwn+CPkbAAn35pUfi4+/i3rEDJ5I
8jOKGksIL4k4bqgXHnWc/cw+kosbFiNBnbfVdDco7YnW1R1EmHiEF3Rg/ZUTfbgG
HWbQU3vlIWduG1M8haZCjwifiBdS4nsM2s6My2Sk0b4p1bOvu5JGrE7MYDRorGzM
dsEb3/BQhzzS1ZTiHNPwaPTUhsO+WtYYfW710La8vL08asAa/UBUKsM0bOzxcsse
mtdvnv9M8V9aql1F33YwqzGU4RYoBJ0CLEuh6k+vuc7xJqVeXgV1mEnMtEi8XPTn
J4tJpH1eRzF4fSJK1IkoB1s44pO4bsiV8Ilk6p0G+EhFYp043j/kU4vR8ijhwZCD
2jFMu5numuMS3yBzzTkikMELd8RZz/MKE5ZDyRqHytwSByegRkAIyELELj3hYFTg
8AvwTSjgWfAg/1fkCwMnX349ltkzCpxbKxPqEA5WmaaPS3Yq+iNGze4u2fQhIRCs
YSPBoadXH8Pt37WeMD5agDgrqDitqn8er4EeACkWGwmUkENaxrcjksw/ZYHzqpVn
soUjhMfZa4VfF0rfW3e4JTIAkakJz6X3bFbeh3MS9FmOsF+RfWiq0R9lEgOWUZGR
rYKgXVxdb0W/7LPQ33wMTbX1hpkCN17D7YpK9K2XjGM/8nzqVKOCo3f0cwPtF02z
ZSseekdZph6+PDxhbRbiCmdT7u3ZlezDkzqKAspaVbHDfYmy6rzG0k1Q9YVGhBIC
2CMxxYic6vCu9x0YODwaIsrsq9wWettwNY7QMFraeuu7SrwC+RIi8KA1vz47uVr/
pImYkw5GwBI5YyFqgUgE3RQryU1chAJcWCjRa4sdNPfvJ2aIAnsvfE9Gb11sCyv3
y/z++eMI7vOGT9V9fo5eUGPjMiwwV4dAnsSmUQ2PSySVgd7TZyXBPVORjsKm8Nej
3ehDuxu86L1/KGKbEBy+8oquKzIpzrjCitp79IwIMN2+OhQ+/wjH9Wm76qo5tll4
Q2rpto8Ay96iMwYAv29Zu4HwqM+rvkGwlkM6gfIo3LfacFk7Ef6uXADl41e7WLIv
ak3YtPSgGUAryKlwFbLHnXfD6vVvGj6nveo5Lozd50aO3BgudioZhbGXS8NESa7I
EGV06ToEenwtDu3xXMFqfGTapyteW84kkOup5tHS4VIfZgg+3aFCU4Xl1Q5/Xlfe
0F3dTOjqLSM1xh79HcJavC+qhWjE1nPTph0N6e1vEZxyaDQQw6PNquuECLJIGK6Y
GJKujMkVLT3K5VTiAHuVbpUx5+quASaT2G5MrokaCkBED83MrVGigsT8S+UP3fvn
yrMJApyrasIdvtdGOUiGYsge0NiZquIMrfarxfXSjWIuI+CSmEvMNF6J77Snu+DB
f2E0glxFJtHwD/dJhWzCWAdAV7hkj4Pc68R+tjtIKW+cvencGMgZNQliszmXdyAC
ROV5krVxfeunpslsgswijSejiutXM5B60OX2h5Pg0pijY0CvP/AnlKviUXY+/TAX
PtJWd3LuO51aossEctuLd9agAe+Pr5Xi9t18N2bg2aFk32nc6hba3hqt8Gn3iwXG
DK1m5qK8YTrWaopXzDYrUYo8Ot5oD9MxRz7l77p3eQ3xutod56E0DiTzp1/uGAIV
HtrMZPncNh00PpvzGuMf6AwVPtMablts+IOasqVxph857XqB7RlSOzqJ4detJck1
bs0DSl7PQgYJV4C5jJled8zU6svlawcmsqdw14jzTc+Os7n2eDCKpCcUNkAm7vbW
3jwVkUXEEFwa+cyPidNvmT80WmbjuNhXrChOzgZS5GW77YH/vuhYwEgbxhPlaMR+
+fxk84NSKt9PMsTglTNcMi26/I2zH88Qrc2DGQyOhW9f9hEs2tChCPxSHi3zNFVP
lCGkz56NqctrlY34GCW2cM4ialuZobe5/8huZdF2RYRdK8y5y5GsPmlDKJ4qg+xS
WWgTSG2vYa8DvTA4nzuGY9CyTBEM4LPnV89h0e8/p1cFHxcKlAzd+we5Q5DPKmQv
W7JTIDyL+Yqz5yZmboBj+GhHZQQx8Rm012kd/rmL10hDRpGD+ka/uELfwkrQWIFt
dOJViRIGF3WfREXWsbM0+6KJPXewA9tC+PLS4dvmMEudtnOfQjYXd9eSZUAI4KcS
kr9DlCfcl0hR47crItpfOSE2gdq7kqqu5mRgJl9kCSiJSx+kYMGpq6qGDfoyM/TC
l8bzBSbYJS2VQ1IM7dZHwTWlxkphcVQhUhOidLri94wCakeV5KguVNS+ewxCNR4h
PoSBa4/C1Ht6B2yESqDewzCpfOEJ7/O7yCVUZmKDvB+R6yXyeJss4FzN9kGsjaRa
TpVZtM0XDlFTqzGdXpqCx+qn2OoQqdEAXiog3WyD6Cet4IrhZlfOC3e2tWZE3piO
bxT8Ud5wPF8yEnjAQQsxFVWaUobXbWaFim7U+/eZuc7jzNMGIQ5ib5IegDRbHCS4
z+2bCZT9itz4NzBmllVURiybCCiRz5KIVMwlXYaLoFmqaiXMiTujENrY6F+vV7sD
9+X+eguzRdIe2howLxM7f2TKOiyxeLo1Ng/YGBkAXtyadb13YfDiyvzZUOCnRZLw
hB+z3ZDEqqB4l0z5vp+l7iDnbVQyR6rA3fMqGWppfejEfD7KUof81Xcv1eOZhPKV
eQX34krsy/jIz1C4g5EN9csEqSbIkA3ObV3BnBUWZV8JaCJ3ZJF3CcNy2BElwT+S
IyqAl+JVEqplHgX4qJvgHVc6vErNZjnM7CxzIqM81i0NkrfsVIrC67t9w+gybAqg
oqrmALnAX9XGS2y3UTLfKdJCxlHMAzh5YVc90YbGQBqsUlZLCEQAVSfq0juqXr2h
VDj9p9pH1L8MtIadRDyn0WrcGBKid24uIv64t7/ahhFjoHakMXfDsXmRYOyCPQGu
0PhwhoFLpgi6Jq1kl5utBax8FPXr5frOpIGSPdCcXDNmdiiVX5O35JnwGZ/ec/+o
8r+I5yuBkFCG+mstdcpzd34xTLjcau48+rfBnNwNQGAk1Z6vYk9/WJCrGsurDn/1
31RA3HtzQbQjLkUBo32fQ/kZRXpRfMQJSKxlc34qyTP7V/2mkXvSNfgYOH6w/Xw/
JEUOyUjVOmSkCk+NTowNvFEUwNovQHAmjMxeeYq/24JQ6diFBUbUnVHkb9ZQfGdq
gx9IXUfFdAqbDwPxTGb7UecdFw6Q9a9SFD/6ZY8F+YgF1uA4aU0XgmSmVvAq5IDj
b2hEdpj6D51/u/7k2M2Es/UtRcXES1tz7Ey7DbyEI+arGtUfuola87nB7eO7/Bbb
/Jr0c5NxUqM6u2YSRp1zZOjJGUarDU4qA24HbWZIoE63TxQsjYLp09kOaZE0smgG
YiWWxyO4NmqPGKx8PEcDUDX3/wNtRPrMwbygsOievUOPpOpicUj5/hsHogXqwZ52
T8/fG+SP3mfRMMDjxFGiTg==
`protect END_PROTECTED
