`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGGRKOkeFgxzPkfp82mCj6mBO8UYgLewtAXAdw76/S7sFom1Y61wsoNR+1RhBmWz
vTWQaU9FcTxnv/EujKrQI5sBqRqBLCm5FO5n2A9gqDLUEhBO23i5HVtpbP12QaoG
Phd2JkP1uFCf6FbSkBrEAd/cMazmwbfmG1XWWphf4bVmAX/6LXNxtTkIZh4Z45QR
t5QeDWl6ahZZFz5Nx2A9XGgotuuuPNOgndYRbGDnmcG0VaHSXnhijS0SAhz9x1OZ
FFEgc2E+NJoB9vAFq6SL07x2+ZKUzidxmWxpa7m9WFgaCfIQhOSd8Zj6HYIdj+D9
VAne9TKuTEUibToVQ7K2rvNPjPkedC9z2W7KynRb5/hSbqMvrU7z8kZWsCdJZrW/
r/6++a3+LlyPYuRMo6TKnenQTdYLtMIo2uPURWFMbhoOstarjpFkQQaMWhUo1eyU
5ZN/D80GmYflKkU8lkGt91v2R6oy/vg5knBj6/5qtP+DYyWZL+VFm28//Xgnb2ys
kUBrplDf/rw3dpi+ghKEA9wLSmaU44aOaXS4jlK0kcpk5L0zefq3df/nDsFr5rtH
tDZzaPTlEKFM4y+ioyztxCGiRRzSJedV5LEqwMWssY4Q2Tc4DCl+0v0tFYezFD24
Kkt5M/hIfrPeJXJtjrHYNg==
`protect END_PROTECTED
