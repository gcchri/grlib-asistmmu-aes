library verilog;
use verilog.vl_types.all;
entity GTXE1_WRAP is
    generic(
        AC_CAP_DIS      : string  := "TRUE";
        ALIGN_COMMA_WORD: integer := 1;
        BGTEST_CFG      : string  := "00";
        BIAS_CFG        : string  := "00000";
        CDR_PH_ADJ_TIME : string  := "10100";
        CHAN_BOND_1_MAX_SKEW: integer := 7;
        CHAN_BOND_2_MAX_SKEW: integer := 1;
        CHAN_BOND_KEEP_ALIGN: string  := "FALSE";
        CHAN_BOND_SEQ_1_1: string  := "0101111100";
        CHAN_BOND_SEQ_1_2: string  := "0001001010";
        CHAN_BOND_SEQ_1_3: string  := "0001001010";
        CHAN_BOND_SEQ_1_4: string  := "0110111100";
        CHAN_BOND_SEQ_1_ENABLE: string  := "1111";
        CHAN_BOND_SEQ_2_1: string  := "0100111100";
        CHAN_BOND_SEQ_2_2: string  := "0100111100";
        CHAN_BOND_SEQ_2_3: string  := "0110111100";
        CHAN_BOND_SEQ_2_4: string  := "0100111100";
        CHAN_BOND_SEQ_2_CFG: string  := "00000";
        CHAN_BOND_SEQ_2_ENABLE: string  := "1111";
        CHAN_BOND_SEQ_2_USE: string  := "FALSE";
        CHAN_BOND_SEQ_LEN: integer := 1;
        CLK_CORRECT_USE : string  := "TRUE";
        CLK_COR_ADJ_LEN : integer := 1;
        CLK_COR_DET_LEN : integer := 1;
        CLK_COR_INSERT_IDLE_FLAG: string  := "FALSE";
        CLK_COR_KEEP_IDLE: string  := "FALSE";
        CLK_COR_MAX_LAT : integer := 20;
        CLK_COR_MIN_LAT : integer := 18;
        CLK_COR_PRECEDENCE: string  := "TRUE";
        CLK_COR_REPEAT_WAIT: integer := 0;
        CLK_COR_SEQ_1_1 : string  := "0100011100";
        CLK_COR_SEQ_1_2 : string  := "0000000000";
        CLK_COR_SEQ_1_3 : string  := "0000000000";
        CLK_COR_SEQ_1_4 : string  := "0000000000";
        CLK_COR_SEQ_1_ENABLE: string  := "1111";
        CLK_COR_SEQ_2_1 : string  := "0000000000";
        CLK_COR_SEQ_2_2 : string  := "0000000000";
        CLK_COR_SEQ_2_3 : string  := "0000000000";
        CLK_COR_SEQ_2_4 : string  := "0000000000";
        CLK_COR_SEQ_2_ENABLE: string  := "1111";
        CLK_COR_SEQ_2_USE: string  := "FALSE";
        CM_TRIM         : string  := "01";
        COMMA_10B_ENABLE: string  := "1111111111";
        COMMA_DOUBLE    : string  := "FALSE";
        COM_BURST_VAL   : string  := "1111";
        DEC_MCOMMA_DETECT: string  := "TRUE";
        DEC_PCOMMA_DETECT: string  := "TRUE";
        DEC_VALID_COMMA_ONLY: string  := "TRUE";
        DFE_CAL_TIME    : string  := "01100";
        DFE_CFG         : string  := "00011011";
        GEARBOX_ENDEC   : string  := "000";
        GEN_RXUSRCLK    : string  := "TRUE";
        GEN_TXUSRCLK    : string  := "TRUE";
        GTX_CFG_PWRUP   : string  := "TRUE";
        MCOMMA_10B_VALUE: string  := "1010000011";
        MCOMMA_DETECT   : string  := "TRUE";
        OOBDETECT_THRESHOLD: string  := "011";
        PCI_EXPRESS_MODE: string  := "FALSE";
        PCOMMA_10B_VALUE: string  := "0101111100";
        PCOMMA_DETECT   : string  := "TRUE";
        PMA_CAS_CLK_EN  : string  := "FALSE";
        PMA_CDR_SCAN    : string  := "640404C";
        PMA_CFG         : string  := "0040000040000000003";
        PMA_RXSYNC_CFG  : string  := "00";
        PMA_RX_CFG      : string  := "05CE048";
        PMA_TX_CFG      : string  := "00082";
        POWER_SAVE      : string  := "0000110100";
        RCV_TERM_GND    : string  := "FALSE";
        RCV_TERM_VTTRX  : string  := "TRUE";
        RXGEARBOX_USE   : string  := "FALSE";
        RXPLL_COM_CFG   : string  := "21680A";
        RXPLL_CP_CFG    : string  := "00";
        RXPLL_DIVSEL45_FB: integer := 5;
        RXPLL_DIVSEL_FB : integer := 2;
        RXPLL_DIVSEL_OUT: integer := 1;
        RXPLL_DIVSEL_REF: integer := 1;
        RXPLL_LKDET_CFG : string  := "111";
        RXPRBSERR_LOOPBACK: string  := "0";
        RXRECCLK_CTRL   : string  := "RXRECCLKPCS";
        RXRECCLK_DLY    : string  := "0000000000";
        RXUSRCLK_DLY    : string  := "0000";
        RX_BUFFER_USE   : string  := "TRUE";
        RX_CLK25_DIVIDER: integer := 6;
        RX_DATA_WIDTH   : integer := 20;
        RX_DECODE_SEQ_MATCH: string  := "TRUE";
        RX_DLYALIGN_CTRINC: string  := "0100";
        RX_DLYALIGN_EDGESET: string  := "00110";
        RX_DLYALIGN_LPFINC: string  := "0111";
        RX_DLYALIGN_MONSEL: string  := "000";
        RX_DLYALIGN_OVRDSETTING: string  := "00000000";
        RX_EN_IDLE_HOLD_CDR: string  := "FALSE";
        RX_EN_IDLE_HOLD_DFE: string  := "TRUE";
        RX_EN_IDLE_RESET_BUF: string  := "TRUE";
        RX_EN_IDLE_RESET_FR: string  := "TRUE";
        RX_EN_IDLE_RESET_PH: string  := "TRUE";
        RX_EN_MODE_RESET_BUF: string  := "TRUE";
        RX_EN_RATE_RESET_BUF: string  := "TRUE";
        RX_EN_REALIGN_RESET_BUF: string  := "FALSE";
        RX_EN_REALIGN_RESET_BUF2: string  := "FALSE";
        RX_EYE_OFFSET   : string  := "4C";
        RX_EYE_SCANMODE : string  := "00";
        RX_FIFO_ADDR_MODE: string  := "FULL";
        RX_IDLE_HI_CNT  : string  := "1000";
        RX_IDLE_LO_CNT  : string  := "0000";
        RX_LOSS_OF_SYNC_FSM: string  := "FALSE";
        RX_LOS_INVALID_INCR: integer := 1;
        RX_LOS_THRESHOLD: integer := 4;
        RX_OVERSAMPLE_MODE: string  := "FALSE";
        RX_SLIDE_AUTO_WAIT: integer := 5;
        RX_SLIDE_MODE   : string  := "OFF";
        RX_XCLK_SEL     : string  := "RXREC";
        SAS_MAX_COMSAS  : integer := 52;
        SAS_MIN_COMSAS  : integer := 40;
        SATA_BURST_VAL  : string  := "100";
        SATA_IDLE_VAL   : string  := "100";
        SATA_MAX_BURST  : integer := 7;
        SATA_MAX_INIT   : integer := 22;
        SATA_MAX_WAKE   : integer := 7;
        SATA_MIN_BURST  : integer := 4;
        SATA_MIN_INIT   : integer := 12;
        SATA_MIN_WAKE   : integer := 4;
        SHOW_REALIGN_COMMA: string  := "TRUE";
        SIM_GTXRESET_SPEEDUP: integer := 1;
        SIM_RECEIVER_DETECT_PASS: string  := "TRUE";
        SIM_RXREFCLK_SOURCE: string  := "000";
        SIM_TXREFCLK_SOURCE: string  := "000";
        SIM_TX_ELEC_IDLE_LEVEL: string  := "X";
        SIM_VERSION     : string  := "2.0";
        TERMINATION_CTRL: string  := "10100";
        TERMINATION_OVRD: string  := "FALSE";
        TRANS_TIME_FROM_P2: string  := "03C";
        TRANS_TIME_NON_P2: string  := "19";
        TRANS_TIME_RATE : string  := "0E";
        TRANS_TIME_TO_P2: string  := "064";
        TST_ATTR        : string  := "00000000";
        TXDRIVE_LOOPBACK_HIZ: string  := "FALSE";
        TXDRIVE_LOOPBACK_PD: string  := "FALSE";
        TXGEARBOX_USE   : string  := "FALSE";
        TXOUTCLK_CTRL   : string  := "TXOUTCLKPCS";
        TXOUTCLK_DLY    : string  := "0000000000";
        TXPLL_COM_CFG   : string  := "21680A";
        TXPLL_CP_CFG    : string  := "00";
        TXPLL_DIVSEL45_FB: integer := 5;
        TXPLL_DIVSEL_FB : integer := 2;
        TXPLL_DIVSEL_OUT: integer := 1;
        TXPLL_DIVSEL_REF: integer := 1;
        TXPLL_LKDET_CFG : string  := "111";
        TXPLL_SATA      : string  := "00";
        TX_BUFFER_USE   : string  := "TRUE";
        TX_BYTECLK_CFG  : string  := "00";
        TX_CLK25_DIVIDER: integer := 6;
        TX_CLK_SOURCE   : string  := "RXPLL";
        TX_DATA_WIDTH   : integer := 20;
        TX_DEEMPH_0     : string  := "11010";
        TX_DEEMPH_1     : string  := "10000";
        TX_DETECT_RX_CFG: string  := "1832";
        TX_DLYALIGN_CTRINC: string  := "0100";
        TX_DLYALIGN_LPFINC: string  := "0110";
        TX_DLYALIGN_MONSEL: string  := "000";
        TX_DLYALIGN_OVRDSETTING: string  := "10000000";
        TX_DRIVE_MODE   : string  := "DIRECT";
        TX_EN_RATE_RESET_BUF: string  := "TRUE";
        TX_IDLE_ASSERT_DELAY: string  := "100";
        TX_IDLE_DEASSERT_DELAY: string  := "010";
        TX_MARGIN_FULL_0: string  := "1001110";
        TX_MARGIN_FULL_1: string  := "1001001";
        TX_MARGIN_FULL_2: string  := "1000101";
        TX_MARGIN_FULL_3: string  := "1000010";
        TX_MARGIN_FULL_4: string  := "1000000";
        TX_MARGIN_LOW_0 : string  := "1000110";
        TX_MARGIN_LOW_1 : string  := "1000100";
        TX_MARGIN_LOW_2 : string  := "1000010";
        TX_MARGIN_LOW_3 : string  := "1000000";
        TX_MARGIN_LOW_4 : string  := "1000000";
        TX_OVERSAMPLE_MODE: string  := "FALSE";
        TX_PMADATA_OPT  : string  := "0";
        TX_TDCC_CFG     : string  := "11";
        TX_USRCLK_CFG   : string  := "00";
        TX_XCLK_SEL     : string  := "TXUSR"
    );
    port(
        COMFINISH       : out    vl_logic;
        COMINITDET      : out    vl_logic;
        COMSASDET       : out    vl_logic;
        COMWAKEDET      : out    vl_logic;
        DFECLKDLYADJMON : out    vl_logic_vector(5 downto 0);
        DFEEYEDACMON    : out    vl_logic_vector(4 downto 0);
        DFESENSCAL      : out    vl_logic_vector(2 downto 0);
        DFETAP1MONITOR  : out    vl_logic_vector(4 downto 0);
        DFETAP2MONITOR  : out    vl_logic_vector(4 downto 0);
        DFETAP3MONITOR  : out    vl_logic_vector(3 downto 0);
        DFETAP4MONITOR  : out    vl_logic_vector(3 downto 0);
        DRDY            : out    vl_logic;
        DRPDO           : out    vl_logic_vector(15 downto 0);
        MGTREFCLKFAB    : out    vl_logic_vector(1 downto 0);
        PHYSTATUS       : out    vl_logic;
        RXBUFSTATUS     : out    vl_logic_vector(2 downto 0);
        RXBYTEISALIGNED : out    vl_logic;
        RXBYTEREALIGN   : out    vl_logic;
        RXCHANBONDSEQ   : out    vl_logic;
        RXCHANISALIGNED : out    vl_logic;
        RXCHANREALIGN   : out    vl_logic;
        RXCHARISCOMMA   : out    vl_logic_vector(3 downto 0);
        RXCHARISK       : out    vl_logic_vector(3 downto 0);
        RXCHBONDO       : out    vl_logic_vector(3 downto 0);
        RXCLKCORCNT     : out    vl_logic_vector(2 downto 0);
        RXCOMMADET      : out    vl_logic;
        RXDATA          : out    vl_logic_vector(31 downto 0);
        RXDATAVALID     : out    vl_logic;
        RXDISPERR       : out    vl_logic_vector(3 downto 0);
        RXDLYALIGNMONITOR: out    vl_logic_vector(7 downto 0);
        RXELECIDLE      : out    vl_logic;
        RXHEADER        : out    vl_logic_vector(2 downto 0);
        RXHEADERVALID   : out    vl_logic;
        RXLOSSOFSYNC    : out    vl_logic_vector(1 downto 0);
        RXNOTINTABLE    : out    vl_logic_vector(3 downto 0);
        RXOVERSAMPLEERR : out    vl_logic;
        RXPLLLKDET      : out    vl_logic;
        RXPRBSERR       : out    vl_logic;
        RXRATEDONE      : out    vl_logic;
        RXRECCLK        : out    vl_logic;
        RXRECCLKPCS     : out    vl_logic;
        RXRESETDONE     : out    vl_logic;
        RXRUNDISP       : out    vl_logic_vector(3 downto 0);
        RXSTARTOFSEQ    : out    vl_logic;
        RXSTATUS        : out    vl_logic_vector(2 downto 0);
        RXVALID         : out    vl_logic;
        TSTOUT          : out    vl_logic_vector(9 downto 0);
        TXBUFSTATUS     : out    vl_logic_vector(1 downto 0);
        TXDLYALIGNMONITOR: out    vl_logic_vector(7 downto 0);
        TXGEARBOXREADY  : out    vl_logic;
        TXKERR          : out    vl_logic_vector(3 downto 0);
        TXN             : out    vl_logic;
        TXOUTCLK        : out    vl_logic;
        TXOUTCLKPCS     : out    vl_logic;
        TXP             : out    vl_logic;
        TXPLLLKDET      : out    vl_logic;
        TXRATEDONE      : out    vl_logic;
        TXRESETDONE     : out    vl_logic;
        TXRUNDISP       : out    vl_logic_vector(3 downto 0);
        DADDR           : in     vl_logic_vector(7 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DFECLKDLYADJ    : in     vl_logic_vector(5 downto 0);
        DFEDLYOVRD      : in     vl_logic;
        DFETAPOVRD      : in     vl_logic;
        DFETAP1         : in     vl_logic_vector(4 downto 0);
        DFETAP2         : in     vl_logic_vector(4 downto 0);
        DFETAP3         : in     vl_logic_vector(3 downto 0);
        DFETAP4         : in     vl_logic_vector(3 downto 0);
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        GATERXELECIDLE  : in     vl_logic;
        GREFCLKRX       : in     vl_logic;
        GREFCLKTX       : in     vl_logic;
        GTXRXRESET      : in     vl_logic;
        GTXTEST         : in     vl_logic_vector(12 downto 0);
        GTXTXRESET      : in     vl_logic;
        IGNORESIGDET    : in     vl_logic;
        LOOPBACK        : in     vl_logic_vector(2 downto 0);
        MGTREFCLKRX     : in     vl_logic_vector(1 downto 0);
        MGTREFCLKTX     : in     vl_logic_vector(1 downto 0);
        NORTHREFCLKRX   : in     vl_logic_vector(1 downto 0);
        NORTHREFCLKTX   : in     vl_logic_vector(1 downto 0);
        PERFCLKRX       : in     vl_logic;
        PERFCLKTX       : in     vl_logic;
        PLLRXRESET      : in     vl_logic;
        PLLTXRESET      : in     vl_logic;
        PRBSCNTRESET    : in     vl_logic;
        RXBUFRESET      : in     vl_logic;
        RXCDRRESET      : in     vl_logic;
        RXCHBONDI       : in     vl_logic_vector(3 downto 0);
        RXCHBONDLEVEL   : in     vl_logic_vector(2 downto 0);
        RXCHBONDMASTER  : in     vl_logic;
        RXCHBONDSLAVE   : in     vl_logic;
        RXCOMMADETUSE   : in     vl_logic;
        RXDEC8B10BUSE   : in     vl_logic;
        RXDLYALIGNDISABLE: in     vl_logic;
        RXDLYALIGNMONENB: in     vl_logic;
        RXDLYALIGNOVERRIDE: in     vl_logic;
        RXDLYALIGNRESET : in     vl_logic;
        RXDLYALIGNSWPPRECURB: in     vl_logic;
        RXDLYALIGNUPDSW : in     vl_logic;
        RXENCHANSYNC    : in     vl_logic;
        RXENMCOMMAALIGN : in     vl_logic;
        RXENPCOMMAALIGN : in     vl_logic;
        RXENPMAPHASEALIGN: in     vl_logic;
        RXENPRBSTST     : in     vl_logic_vector(2 downto 0);
        RXENSAMPLEALIGN : in     vl_logic;
        RXEQMIX         : in     vl_logic_vector(9 downto 0);
        RXGEARBOXSLIP   : in     vl_logic;
        RXN             : in     vl_logic;
        RXP             : in     vl_logic;
        RXPLLLKDETEN    : in     vl_logic;
        RXPLLPOWERDOWN  : in     vl_logic;
        RXPLLREFSELDY   : in     vl_logic_vector(2 downto 0);
        RXPMASETPHASE   : in     vl_logic;
        RXPOLARITY      : in     vl_logic;
        RXPOWERDOWN     : in     vl_logic_vector(1 downto 0);
        RXRATE          : in     vl_logic_vector(1 downto 0);
        RXRESET         : in     vl_logic;
        RXSLIDE         : in     vl_logic;
        RXUSRCLK        : in     vl_logic;
        RXUSRCLK2       : in     vl_logic;
        SOUTHREFCLKRX   : in     vl_logic_vector(1 downto 0);
        SOUTHREFCLKTX   : in     vl_logic_vector(1 downto 0);
        TSTCLK0         : in     vl_logic;
        TSTCLK1         : in     vl_logic;
        TSTIN           : in     vl_logic_vector(19 downto 0);
        TXBUFDIFFCTRL   : in     vl_logic_vector(2 downto 0);
        TXBYPASS8B10B   : in     vl_logic_vector(3 downto 0);
        TXCHARDISPMODE  : in     vl_logic_vector(3 downto 0);
        TXCHARDISPVAL   : in     vl_logic_vector(3 downto 0);
        TXCHARISK       : in     vl_logic_vector(3 downto 0);
        TXCOMINIT       : in     vl_logic;
        TXCOMSAS        : in     vl_logic;
        TXCOMWAKE       : in     vl_logic;
        TXDATA          : in     vl_logic_vector(31 downto 0);
        TXDEEMPH        : in     vl_logic;
        TXDETECTRX      : in     vl_logic;
        TXDIFFCTRL      : in     vl_logic_vector(3 downto 0);
        TXDLYALIGNDISABLE: in     vl_logic;
        TXDLYALIGNMONENB: in     vl_logic;
        TXDLYALIGNOVERRIDE: in     vl_logic;
        TXDLYALIGNRESET : in     vl_logic;
        TXDLYALIGNUPDSW : in     vl_logic;
        TXELECIDLE      : in     vl_logic;
        TXENC8B10BUSE   : in     vl_logic;
        TXENPMAPHASEALIGN: in     vl_logic;
        TXENPRBSTST     : in     vl_logic_vector(2 downto 0);
        TXHEADER        : in     vl_logic_vector(2 downto 0);
        TXINHIBIT       : in     vl_logic;
        TXMARGIN        : in     vl_logic_vector(2 downto 0);
        TXPDOWNASYNCH   : in     vl_logic;
        TXPLLLKDETEN    : in     vl_logic;
        TXPLLPOWERDOWN  : in     vl_logic;
        TXPLLREFSELDY   : in     vl_logic_vector(2 downto 0);
        TXPMASETPHASE   : in     vl_logic;
        TXPOLARITY      : in     vl_logic;
        TXPOSTEMPHASIS  : in     vl_logic_vector(4 downto 0);
        TXPOWERDOWN     : in     vl_logic_vector(1 downto 0);
        TXPRBSFORCEERR  : in     vl_logic;
        TXPREEMPHASIS   : in     vl_logic_vector(3 downto 0);
        TXRATE          : in     vl_logic_vector(1 downto 0);
        TXRESET         : in     vl_logic;
        TXSEQUENCE      : in     vl_logic_vector(6 downto 0);
        TXSTARTSEQ      : in     vl_logic;
        TXSWING         : in     vl_logic;
        TXUSRCLK        : in     vl_logic;
        TXUSRCLK2       : in     vl_logic;
        USRCODEERR      : in     vl_logic;
        GSR             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AC_CAP_DIS : constant is 1;
    attribute mti_svvh_generic_type of ALIGN_COMMA_WORD : constant is 2;
    attribute mti_svvh_generic_type of BGTEST_CFG : constant is 1;
    attribute mti_svvh_generic_type of BIAS_CFG : constant is 1;
    attribute mti_svvh_generic_type of CDR_PH_ADJ_TIME : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_1_MAX_SKEW : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_2_MAX_SKEW : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_KEEP_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_1 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_2 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_3 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_4 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_1 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_2 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_3 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_4 : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_CFG : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_USE : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_LEN : constant is 2;
    attribute mti_svvh_generic_type of CLK_CORRECT_USE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_ADJ_LEN : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_DET_LEN : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_INSERT_IDLE_FLAG : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_KEEP_IDLE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_MAX_LAT : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_MIN_LAT : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_PRECEDENCE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_REPEAT_WAIT : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_1 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_2 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_3 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_4 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_1 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_2 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_3 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_4 : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_USE : constant is 1;
    attribute mti_svvh_generic_type of CM_TRIM : constant is 1;
    attribute mti_svvh_generic_type of COMMA_10B_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of COMMA_DOUBLE : constant is 1;
    attribute mti_svvh_generic_type of COM_BURST_VAL : constant is 1;
    attribute mti_svvh_generic_type of DEC_MCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of DEC_PCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of DEC_VALID_COMMA_ONLY : constant is 1;
    attribute mti_svvh_generic_type of DFE_CAL_TIME : constant is 1;
    attribute mti_svvh_generic_type of DFE_CFG : constant is 1;
    attribute mti_svvh_generic_type of GEARBOX_ENDEC : constant is 1;
    attribute mti_svvh_generic_type of GEN_RXUSRCLK : constant is 1;
    attribute mti_svvh_generic_type of GEN_TXUSRCLK : constant is 1;
    attribute mti_svvh_generic_type of GTX_CFG_PWRUP : constant is 1;
    attribute mti_svvh_generic_type of MCOMMA_10B_VALUE : constant is 1;
    attribute mti_svvh_generic_type of MCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of OOBDETECT_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of PCI_EXPRESS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCOMMA_10B_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CAS_CLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CDR_SCAN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG : constant is 1;
    attribute mti_svvh_generic_type of PMA_RXSYNC_CFG : constant is 1;
    attribute mti_svvh_generic_type of PMA_RX_CFG : constant is 1;
    attribute mti_svvh_generic_type of PMA_TX_CFG : constant is 1;
    attribute mti_svvh_generic_type of POWER_SAVE : constant is 1;
    attribute mti_svvh_generic_type of RCV_TERM_GND : constant is 1;
    attribute mti_svvh_generic_type of RCV_TERM_VTTRX : constant is 1;
    attribute mti_svvh_generic_type of RXGEARBOX_USE : constant is 1;
    attribute mti_svvh_generic_type of RXPLL_COM_CFG : constant is 1;
    attribute mti_svvh_generic_type of RXPLL_CP_CFG : constant is 1;
    attribute mti_svvh_generic_type of RXPLL_DIVSEL45_FB : constant is 2;
    attribute mti_svvh_generic_type of RXPLL_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of RXPLL_DIVSEL_OUT : constant is 2;
    attribute mti_svvh_generic_type of RXPLL_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of RXPLL_LKDET_CFG : constant is 1;
    attribute mti_svvh_generic_type of RXPRBSERR_LOOPBACK : constant is 1;
    attribute mti_svvh_generic_type of RXRECCLK_CTRL : constant is 1;
    attribute mti_svvh_generic_type of RXRECCLK_DLY : constant is 1;
    attribute mti_svvh_generic_type of RXUSRCLK_DLY : constant is 1;
    attribute mti_svvh_generic_type of RX_BUFFER_USE : constant is 1;
    attribute mti_svvh_generic_type of RX_CLK25_DIVIDER : constant is 2;
    attribute mti_svvh_generic_type of RX_DATA_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of RX_DECODE_SEQ_MATCH : constant is 1;
    attribute mti_svvh_generic_type of RX_DLYALIGN_CTRINC : constant is 1;
    attribute mti_svvh_generic_type of RX_DLYALIGN_EDGESET : constant is 1;
    attribute mti_svvh_generic_type of RX_DLYALIGN_LPFINC : constant is 1;
    attribute mti_svvh_generic_type of RX_DLYALIGN_MONSEL : constant is 1;
    attribute mti_svvh_generic_type of RX_DLYALIGN_OVRDSETTING : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_IDLE_HOLD_CDR : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_IDLE_HOLD_DFE : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_IDLE_RESET_BUF : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_IDLE_RESET_FR : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_IDLE_RESET_PH : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_MODE_RESET_BUF : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_RATE_RESET_BUF : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_REALIGN_RESET_BUF : constant is 1;
    attribute mti_svvh_generic_type of RX_EN_REALIGN_RESET_BUF2 : constant is 1;
    attribute mti_svvh_generic_type of RX_EYE_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of RX_EYE_SCANMODE : constant is 1;
    attribute mti_svvh_generic_type of RX_FIFO_ADDR_MODE : constant is 1;
    attribute mti_svvh_generic_type of RX_IDLE_HI_CNT : constant is 1;
    attribute mti_svvh_generic_type of RX_IDLE_LO_CNT : constant is 1;
    attribute mti_svvh_generic_type of RX_LOSS_OF_SYNC_FSM : constant is 1;
    attribute mti_svvh_generic_type of RX_LOS_INVALID_INCR : constant is 2;
    attribute mti_svvh_generic_type of RX_LOS_THRESHOLD : constant is 2;
    attribute mti_svvh_generic_type of RX_OVERSAMPLE_MODE : constant is 1;
    attribute mti_svvh_generic_type of RX_SLIDE_AUTO_WAIT : constant is 2;
    attribute mti_svvh_generic_type of RX_SLIDE_MODE : constant is 1;
    attribute mti_svvh_generic_type of RX_XCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of SAS_MAX_COMSAS : constant is 2;
    attribute mti_svvh_generic_type of SAS_MIN_COMSAS : constant is 2;
    attribute mti_svvh_generic_type of SATA_BURST_VAL : constant is 1;
    attribute mti_svvh_generic_type of SATA_IDLE_VAL : constant is 1;
    attribute mti_svvh_generic_type of SATA_MAX_BURST : constant is 2;
    attribute mti_svvh_generic_type of SATA_MAX_INIT : constant is 2;
    attribute mti_svvh_generic_type of SATA_MAX_WAKE : constant is 2;
    attribute mti_svvh_generic_type of SATA_MIN_BURST : constant is 2;
    attribute mti_svvh_generic_type of SATA_MIN_INIT : constant is 2;
    attribute mti_svvh_generic_type of SATA_MIN_WAKE : constant is 2;
    attribute mti_svvh_generic_type of SHOW_REALIGN_COMMA : constant is 1;
    attribute mti_svvh_generic_type of SIM_GTXRESET_SPEEDUP : constant is 2;
    attribute mti_svvh_generic_type of SIM_RECEIVER_DETECT_PASS : constant is 1;
    attribute mti_svvh_generic_type of SIM_RXREFCLK_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of SIM_TXREFCLK_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of SIM_TX_ELEC_IDLE_LEVEL : constant is 1;
    attribute mti_svvh_generic_type of SIM_VERSION : constant is 1;
    attribute mti_svvh_generic_type of TERMINATION_CTRL : constant is 1;
    attribute mti_svvh_generic_type of TERMINATION_OVRD : constant is 1;
    attribute mti_svvh_generic_type of TRANS_TIME_FROM_P2 : constant is 1;
    attribute mti_svvh_generic_type of TRANS_TIME_NON_P2 : constant is 1;
    attribute mti_svvh_generic_type of TRANS_TIME_RATE : constant is 1;
    attribute mti_svvh_generic_type of TRANS_TIME_TO_P2 : constant is 1;
    attribute mti_svvh_generic_type of TST_ATTR : constant is 1;
    attribute mti_svvh_generic_type of TXDRIVE_LOOPBACK_HIZ : constant is 1;
    attribute mti_svvh_generic_type of TXDRIVE_LOOPBACK_PD : constant is 1;
    attribute mti_svvh_generic_type of TXGEARBOX_USE : constant is 1;
    attribute mti_svvh_generic_type of TXOUTCLK_CTRL : constant is 1;
    attribute mti_svvh_generic_type of TXOUTCLK_DLY : constant is 1;
    attribute mti_svvh_generic_type of TXPLL_COM_CFG : constant is 1;
    attribute mti_svvh_generic_type of TXPLL_CP_CFG : constant is 1;
    attribute mti_svvh_generic_type of TXPLL_DIVSEL45_FB : constant is 2;
    attribute mti_svvh_generic_type of TXPLL_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of TXPLL_DIVSEL_OUT : constant is 2;
    attribute mti_svvh_generic_type of TXPLL_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of TXPLL_LKDET_CFG : constant is 1;
    attribute mti_svvh_generic_type of TXPLL_SATA : constant is 1;
    attribute mti_svvh_generic_type of TX_BUFFER_USE : constant is 1;
    attribute mti_svvh_generic_type of TX_BYTECLK_CFG : constant is 1;
    attribute mti_svvh_generic_type of TX_CLK25_DIVIDER : constant is 2;
    attribute mti_svvh_generic_type of TX_CLK_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of TX_DATA_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of TX_DEEMPH_0 : constant is 1;
    attribute mti_svvh_generic_type of TX_DEEMPH_1 : constant is 1;
    attribute mti_svvh_generic_type of TX_DETECT_RX_CFG : constant is 1;
    attribute mti_svvh_generic_type of TX_DLYALIGN_CTRINC : constant is 1;
    attribute mti_svvh_generic_type of TX_DLYALIGN_LPFINC : constant is 1;
    attribute mti_svvh_generic_type of TX_DLYALIGN_MONSEL : constant is 1;
    attribute mti_svvh_generic_type of TX_DLYALIGN_OVRDSETTING : constant is 1;
    attribute mti_svvh_generic_type of TX_DRIVE_MODE : constant is 1;
    attribute mti_svvh_generic_type of TX_EN_RATE_RESET_BUF : constant is 1;
    attribute mti_svvh_generic_type of TX_IDLE_ASSERT_DELAY : constant is 1;
    attribute mti_svvh_generic_type of TX_IDLE_DEASSERT_DELAY : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_0 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_1 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_2 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_3 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_4 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_0 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_1 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_2 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_3 : constant is 1;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_4 : constant is 1;
    attribute mti_svvh_generic_type of TX_OVERSAMPLE_MODE : constant is 1;
    attribute mti_svvh_generic_type of TX_PMADATA_OPT : constant is 1;
    attribute mti_svvh_generic_type of TX_TDCC_CFG : constant is 1;
    attribute mti_svvh_generic_type of TX_USRCLK_CFG : constant is 1;
    attribute mti_svvh_generic_type of TX_XCLK_SEL : constant is 1;
end GTXE1_WRAP;
