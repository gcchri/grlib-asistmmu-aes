`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FXgVDxnHcpMEgqxo4NfZE34VEUSF3NacknDVdygBenMmR+vyBN/ZVJtymWuBXKgG
WK2tnACIIburttKTjcLwLtj+ZINLqukMo3ZQmf8cu5jie9uXes2Kf6FRIUO3d47t
fcL7rdhw5WEzpwdCM4po2WTnnV+hR56aVhHFq2vQ9yNF1eADyN6/j6Hyw53eQGyU
dUB4u0JkRz6/A/GOlgBpySUbZilhiNy+BNwpmx3lgPjbr27b9aVI1sSNgSDNvTm0
4ZR8Z01svwYigrSeAfpHtd9x4LN5dmYYRxbStPzwmnZjOVtNb+yuJ8H9F5AmGP8y
wUpGIThrXpFTUhDCAk47UEFELiHCo7Brffwe7CqI6+ECKkL68LTyLLPRHSmeRDXH
bA2Yk+0mUkN8b1zAIvaKDhhP4jEnTIbK51VDm3IkJpzhYH5Is4ILygncZWNrkYAq
wHjeY2OiWczT8t6a5FbCk9VqvumNHGGNIuzA++1tmn6g+OiSBQ28w43rlyd1qMzF
A4GZG+np7ZkrOdG+DJAncVeW2JdooqqWdOblmBH4NYTZknjAehfWeqQJMS4Z7RfN
DltPYp5kRSg+Fe1n0eoeEZL9N4wlWzQU2CtZo6FQV0hAKw6eRV92PqMDH9I1qxbt
+KDcb/PNhG4GIeEqWUJic6zElohAu4nuEW6cDvlQ2hf/3yrdODWFRJe+AsZ4cnLl
/NvXiP87OJx9kWEwCtk5CccJpxyQ49YXDSkpsQUS6HlSnwCGClTvW5WdxcYwDuMo
tU+6wg+cTaxs3O/+Lcy3RfnKlA5wJZ5mihMAgRuoDUVzQJaupRP4hdkM53/+CY75
5OeP8HiEpAO9lFFlFfD8S8fWr6zCiPaeDaFoygDjlis7YLuRIDpa1sZPVlt6k3+h
Hdn0H3rrVcBhiur2wUU0FKG2t/hSsrWkubkwfnbMdrgvCTElyZKAm6xmAJcp6JXD
QLFixnGKnupM8ij3j4urkw==
`protect END_PROTECTED
