`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5XuDY1o0nSIZkP5u5oMlbNn91ACYzj5hO6TZlJDqk4cldyghZDgzc/JWN0GG0aRf
dzZ7I9oNZNR8oP44IIua8l3iOHlA5oToAtO6AQUMQvA8w9RF+RJxJ3o+3Nd5/2Qu
n7oHITQmjgozrhr5Au01i1C2soct7YAjgGDcbGJNslN+B0ViIKXBNN7B5DFABs5q
UsL4ZbSA7SkdO5JDneonULEVuMEFX9UDaq8lo3NgqJ0VIQCXYPJMVGQb73Ps548m
eGnUidRrUK0V4YQ9nc4DX1WfeCMC2J854z2HhOswkxyXUUCCu2KGqUPKG1E/X9F6
+5nKVDvNJ3THGQQFGT0HiDqLTAhM7P3DjqDvnNcfrjNxWR3KKgB4CfYfbR21XFf7
PFXIxQyvZ/BnW+ww2DBM+ZC727avRwAv/Waq2gnLutbaTUtEXPOnd3gjv5iSGtcD
hTzrOJITyGCYIR7EhAMdru3WZhO03KfqJMyZHNnPTSdN+1kSx5wdXNEbsRnkPJ7b
mUCcHah7Xza/A7IauDzzNxlFAZEktYQN5IO6QCq7CsLdjktCfgb3litp5OPlo2xp
W2k1vhtEJ3s34TstQMj13YZm/tFyobrn25wZAlHJwKLQz3aG7dlDOGCHIQW7dPAT
wkvrURlvKu8YmMfv+STNyiEgBAQ4S7N7qeZf9G/I0TCpovIrKqp+I42HNyLNOMc/
UTruI5aAbvIPSD0PGIcdJw==
`protect END_PROTECTED
