`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wo255VBRPnTynPOjUOdskUDmY2jBO0AyQ7gd8h0H4weduE8WCvYffgZXdq58sljT
FNQHbuq55MA22NavMj4DvNb3/eowwC4XXyAZ1fxpw0EL0b3k9eY4j10DEVLWFAvU
++1MH0WD1rf6LnEBia+Dx63GjAcP8EhUlv7uOxSLVRTGk00oC7gIu3aHCEPSyZXk
OTS5VCtS4BZ8zp79ejToUs8RkCcbEXcNyZ2DctJnxwKuskrg5qJX6gSHMLm6j0sG
I36FdhTnGbAWfgScRvDPlIvNzzHCt7XgLc5DIQHqUxR4dp34z+Ohs0N8Gihb1sj3
rqPWUSOql+qEM4IJbjbPM2IUw0HRhjDW4VoRIht30eDGPi0di2km4U8loCu/mny6
PfALNBD/JjqAFGPZhCip/g==
`protect END_PROTECTED
