`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZOF57E5pvOUlawo/7uus70FjHFzJqlha1CWPHhc/vrHzmeoReZ4SKAN0tull6Msm
oJ5NfpDWUac36BPsFBINf4+xcs7G6xuHZ4QxOpRriPMqoIU19Gd9v5A7QWxwhtqQ
iJ8s47JZhLC0BWn+VO6V9fZKYKYQwH79n+AQu7z1r9p7xcfNYFG3HKG9zA2P1dtl
itIBO+yWvMEoJEcmnO8W7wBAL6Aj2MDy+LT+YggcPjBO2X0NJbQiRcJTx9nhdOyX
24jmULqOs3E5B7Ne3nJTrvxwN/ckF0116ZQMC6yZ96Q=
`protect END_PROTECTED
