`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kL/ylNTtbbtwO4JNZFauaubiV90Sl/o+/06GoFgUfgZwvOXg9RsevP03ssuMzSh
gqZLi10Vas1xaJRVqzUd31Q5AcoCm01fsvL8e5V5UxjjUPi7heAzlnnWrKha5gC7
TN1ubGDgjB7lmBrXFZUmsn2Rk474EOu2Qz63VtwY7lx7xQBdFRgNustqEru7pcTF
34guCoFsLsRTMcSU1H4R7Q/tbHC/rSLunsKssN6qpNmMigtnxQhBbBlRK7E9E1W/
FvzCnWYmDNY9avoyDFIs7NYTF9mqUpjPbbq3xXuQvyR9o2Ug78+Cn24Qgr2ZgkyX
sPM+6EWVqE4u2Umt/nhNO0DQi/z12jDRShn7D8tPWZ8YToFjX433SJyBGIyMiqqI
DnJ7LyA25zSgmeRknBKYTUMICSCw2RYo2pMam5oxBeQ35TI1+Hbr93U9cNgcZKCs
QY4TUIngm/Nne8XsKfpUA1aAvhFjnrw/Fs7PrgRAro9TT7wMSEag30bDy2NeX2wp
TyFDww+hIaTrVX8skzPzPTKrskuZ6mDkuZ56osGLDBksrqdHzvtHGlw8uuqkKGi3
pqpDUea3Du9DV09xq1tL1zjKt9GIz5Xy3we8KjuYu2aWEHT64MCK4+ghCLXBZqSF
1WrfjM2wLOdpHrMQctm8HaZmjSZLQI3UED+lOVqhwfZe7cPfL73eo310nSDKy2dy
Ng2afJA8Ie0gccCEl4jACIBEFL/BgDnSd5NxrdH3svocvaTGVDJEtdY/X4LulWGJ
vhFZxWWGGG1Aausg226bOQrbx6HjIUdR50KaszYlgoiVapbZ22pigjPM1iK8ZF8H
06wFB721ABCFCBjukFu7rY/lkkubX74NsaEJ0pnyNZuKtMwOUmbVzCv1emaFo5M6
cqjwppVONAzJ3Vdjgu8RA4ZbGjRB74AbZcae/w4LcGJBDV44dboIhqcqxP2oDD6j
w7r0bXV9XYC9l1WpMftpoiLgvrkgu/eaA4+MBSYYMEnn2xKMQds/GEcL2DAj88AH
bllLiIKfyhEn+YEoYGZ1YA==
`protect END_PROTECTED
