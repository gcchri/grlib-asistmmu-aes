`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Op+14ghyTNHd9Fs+4zF6rrb9AJ2B4/s0rZohpaPgIOLHW6eBbuapZQ2u2gpK6q3i
QkoNpsRrdypB79DAtNvk2zY3W7+dJkV9g0gf8B/kJedY7ZyEFawYD7xncqMHLXXC
hokj7nZ/aNpMQSuylq7CHEr89ZU2IqZI2DlpneXE/90hGLXYj4jX0keeqH//JbPa
ibzGo74B2icKqZwpTLh59IQ3Q3zUCvB7YRWqwb+cID+4NMZ1rQa+djaF04ppRxQJ
7ZT+xhJHzy4VEb1HxYf81aWc1jpY+FSTu1WPK25OIQmNWIdyosfqM5zCIuKRaRYf
5XjSBERwzQvx0ZnYchG+WDyo6DIyBkjZb+zt22b7M75ksniuriWolVho8DUnK2Ro
FLCJX+wo8t/oiTc9s/+bDhd2sSpLTKWGBg8gxuaNAps=
`protect END_PROTECTED
