`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XRFhfWtqfd8ZQf9aa9AbqKBz5KJT7/om4a7kascAEloiesW2yN0Ka620KExUJGtr
CLQKg3KsxLI2uY9UkdTydgdB4ZrF12X7CLp5zmsAI3L0faa60VHCxK301P/MKGIg
cPUQOA27AM/Te1JPkf4TADtI77GzcddNuz8RIsvw+RqK0ZnLNTXKbhZhLk+VhfzO
pIJOthNsj7TBxvMeUI1buB6DEwozMXAGToug6PPDcjjgIpyTNAWYb5E3e9Tpc5eT
0b9OpnIdj1GOpjGliNRSjTpiR+khk7KKpu9izuh2MHylaTfEUDe/qqaRpAfiJ+LX
bz/zPz5XaSNiLMkEiKI6+TlDbSGlR7BbHKhUUgB2pa3S33vKxglUShFCeHa5LdE+
HfOJLVqXmKk2q62Q5KlzIKmjRhoVPt8TU+YR3kqC9qOeeLaAkAfjm7cAdGsFCYL3
W/K5vbxXct1R23GWQ9fcUujyKkCuBaiU0KuhnGiXTz8=
`protect END_PROTECTED
