`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7gK/0G5LOJZUf7xwq/2Le1RLT5KRc1Rgl6+S8edDP3O9hNNVOklTeExaATpqx6so
GsuetwpLfe/Avcuk11H3fPN2kOyzMc8hN2VY74urcmcXAYVdFJImSxOpnRRFt6RX
ztEXNQvan92fujcGin4W33S/rBVDygmtrJKlvrHEDTtS1TQ0NCE6liW/dKTeho4+
Wgd87L31RiV0Mk5Kax4miYT0adSliRI2XFLRxGIdjc4eKnpnTjxpkrbfd9EcHsDE
Gv+KKETXdnBB7QGa5dQaROm8ajoDuHwo+LzKE6YBIdTN59soe3AajHq8rYQhUurN
jrxG/fw4PdwYNoGtPulrnluv+KMwyEEqvzTG+biuXyKGcZDOZNPBA60zfF/vcvFa
ZTA53UOPdOe4YtlCax1+0VWO3pwk4eVgPVYpxKORmxUbo77YKsVd7m7B2FcgGqea
joLKHSuZZphc+ff9FZHWzuT2wrgpH0nUKiB6TKJO7rd3+vrTExEOmjMBHNCmdoWK
sO7JSJS8M/RdNZ2P2ksZP1yngghAWuldEgYyRa0UV1e5f+XwX/k2F/0l0K5QTIwb
LEHQXFme2OHkOGLNonBfK+arsIn2kxG1JPuZ16IMU4YlZTnqDny8HiRUZCUlcSgd
VUxJLNFiU852VF0/s9FVkQ==
`protect END_PROTECTED
