`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAJFnWvFQ1PAc9kb7m364jSeUKgEJaHd2awCyBvXHCedFXRK1YWjrE7S+kFpxUBG
OrrklGABxVX4C9rsZu44u/F0716HTKVEqLO+55AwRMj7MQ+9Zcp3gpsNuNrk7l25
H5BgK9yQRzRJgVKNnUDbl93cHfzL0EeqKrc+tkd8aDp6UmIWLMdO5jeq7bHYxvQK
THFeGbhmCGl4s9h1e9OPrlCxUWGaYEmMIDCFymfjMbsH6brBEB+5VWxrcb6hDuCm
Xp4NOs8rh4wOUlrg6kg4TpAc+UvSSBKXKc2xNRgYdX/6vmNwgvZk8CUfhrh/NHic
UKb4WshShpvyvfnXjRgPw5veSoDx4CzSo535jzdcy9S+RPH9f9fW052NX6pTNHKW
9C23gsL9/CfukDDpidOAX3ZwmK5uChX+oVrilYwsphiQYiTNzIreKTWTvRZyohPv
kJrnQqHGiNtb65/OFJfxHHlE6Avt6aHuX8B9LXn9g21Zuo3pdMqMx0al7A10Dm6G
XFJh8oaTmTYnrWR+o7PP809CKu0UU1b/yIIDl2zaYBqsIGkiA7quIyC9xl1RUFA8
+XL09pU3sHpuahqvlnTNzse4+i6jaVBGUQ4kso3R4uPLiNTNQZLCD+6bZ/QQY6Ry
goemVgLaSOCO8YbwzCR1VJrct7qMTHd5xeiIXrYgUavOXJ9wHyWt/gldnj4Wns5j
1AHNFmghSLtR0O3dlmvBojyknJj0boiBaYMFF3EAxZXn1O+T63yg/rXw/9alXfmL
lwod6DjF7jWhU+zsm7M756tp+6DH/J2wI9e2UTbhEJahZWr8g8ejU4946E0evglK
Rx/bfVyh/UlXnp7SS2/xYkFiW5fMSf1Gv6AMmiGIxTwtkq0qdCjR1+Yw76L9y1Le
v6Ebsk4UnWZSkxFaHMjizwDyQ+B/9neGX96yBxZMYsZ3GbKg1kqZH8haE76RqGbz
TNT6w/9R4yv4npXE6qkp6t6EB4ILvEEVXs3AXSzKnk2gYFLVNpy6i3fdbHs+kntT
5xg/9pqQ7S29BOUtcoaipbdKtZO6jH07upOZCwcManJhoOTA7gRQZ1z4vnlxPBLv
ADLYgIuKa4yb0LAlrZLTGr959ORDBQcO3rvH1ohTkJu2/LTw88sZJkYTaupzEIiO
/SiQSvgtk6zqUOOSOKDhtrRxKQyx/iob42wuyWMNdqoI1rBskduRueucSrmC//7y
elsgwsIuWDxbE+Y+W166BSBPwRvcUTCAJkPbZxJLLxT5PVwvwE1mRlqph3i3tduA
zTrUlAlttaJp1IDAAqhZ1NGKa1YmQ+sCjgRKTTGuGiBe4P/mIER1Mzh05YWLAi2F
sFq9yZSsRZJtP380Ndeuk96gEXOIMSkMBo8xFF1aDwLC6a3Pfb8/NhnIw2Gi2m7r
DMIB94o34iwBxejInPGFrvAfhcMg/FpZ2fFFwMU4aliJAP23vchkdcNPmdjWR85V
FIuEbWgCCMfF7oi0VqlyTXHv6vJeeftBIfcKrERDpbD7pI/zEWArfR4TQ7WEONyJ
VJn7nJpHJdsYAJPn/4nZfIGJAjiWVSTqldpdd3szdZ9oUPsQsRaYl3eW2GWhHBy6
YX6DMQUAl/hRGwQqLbdyZ6U3HKr6RjmUbyMzOpldfDgP6DvE/HtghrKAgDnXWG4/
Jivuq46PBLZGN7Edq8SomgxbaVnNFl+O91hdsw9NZ6CAEFf2NQTZNqLwkMHRLZKJ
oAA6BUvaepnhYo6dX0YpcLGk32dRHMpbSz6vT5lDcl7RAkTtV5kSAAHRMRD0lcb+
kGB1vnXq/wpobz0bGlTztwF7dGdXmmFulL6oQlgxri5zjc/QKiYhhFNzi/RFdtGI
hGWDM/MaF7pU0fvDOWbnf6w/3oKyf5KS8T1jaWptxULkHLUg2fH4XVgILVjq1yaG
F+qxk0pZ0445qj+ssEpA91UvbsDJn/Lftdb6cO9zeb/4yGsCYBVkiBCdllP5DN2K
6gUmc4bf3oO2bIWLrx9xm8RGbqor2iBs+cp7b2OhUg8RqQp72iESQA6qhcrp1nsp
u/saU2D1VpQga1QIlSLSv+hqmGIp/I47nveHvnZym/WHS56z5VHzB2whRS/xq//8
XWoYP3aDKMgten5amgdxxOTLgJcNLYlC1WYcghUeu6eekre2Pw1aYJRr2i7vWT/J
0t2VtpQSeOItwn3ikcLpNg3HrWIEuM/v84hWq1hehsrfQaJSdXWPkRnWZn1EpA1W
GrVgwfNigWXaQGcKdUm5/TQYe0qnNeAxk4I0fc3wfBTKeGm/Ffi5JBJYkQ01ytnt
QBM2ILCFdteSwwMc/B7j/rlWcQgM8WQrcBXYCe1JjRdT5Ou+Pv5M7sI8DJ0IpMsY
s8RBQj42HZq/DZrC2w5PTQjiD+M5dLIXp4euBo3NuSruHwO7V1coUpLGFKPLISuJ
UEWOcJzDeRRpQ0H6T/8zViuYRdzxi2JzZfLB4cDwVw9hXzqZ2oR9jL2Umk7OC3MT
e+YBrv1WZdK1pMgL6P4JgHK5w6cIA2uylm3onx0yp46FiUTMUGl0Ocfe/FYI2CTJ
NpFIFlK6QG76qAHLnb5UZaDmbtHP9cks63+3sTGH8Cy/PSNCa3m9a1V036bMZQUU
2mpU1s922m6hIzRfqm13SMIeL7XGQdWRuG79w5cYU+5QCmSPPTYFfWFKTwyaqhG6
cJBTL3VbAl9jUsshZEIMCaM2W+03QoFNyF1M7epsfGuPCdzHxKkn7nEO1TWTO+jk
MtKXj0x32Js60D5WwPoeVSZdHQaVX1lFYZ3aBoHTYFikTmQNW5VB86J1lw9aFC7s
qNHTnbGSGb+xBPxgKBISR8uO6FZsuotNaunoThW1gYepVvQgEsOMed+Hy3liHuTW
8imenn75Yt9p1SSWeJ4bUUOzyIddDqwOnRyTdHZ2+Jb2fwl6lJC1hXjcZ4ks83D4
3Xw0RDV4muKHeJHObmR8Bv4XtzwJe68pLrv90ZWlGtLnlMjbrDnv8WvQkgLzeWP0
skShjsQc3bSzFaBZRF0ZtFzvc0qRsWfHz6+p1p3MxGaevbjC1IfPBpIOGa9xxzLe
00Fuo6mFYB4TRH+mkCgTKn0sWVsuM4skQerrzLIyQnJTioZGMhCxz3mddDRiU+R6
97Fg+oZlAuH/u7z1u4zIet51vCEOj0gDmzdk7j6WWoJQutZac7Mw1G0DTFRVZECC
t9Dm9Vi899kKos1kZB0Z+uc9b8MKqwmwSsrGteHRP8f6525TIij5X3IVOF9AL+z7
1vfhRp/XHcPvZvES3Y2bgjxTgKt/6d3LH7vSxsOhGcrjUuzvYTjJXEvtwtKkOpKW
tNw1RWOti2e6fkx2xhZVAEPl7drH3MX+nA7XvZNHupmvP1y7b6nd+gL/SW7XDTs5
IfhSn/HE7tJge1cdFCi0D5UoKdc35Iffjr8qXdULfrFZDU8l9JAAFkvw2B81bPxR
JO1F6raBy+wEYupdKogr5VwNABjt7JEJ+ESTMIDVV9GAEJOJHSR46GW/HAVLeAri
/QGRVQ5DcEsruD2iIdzwmm0+WM0XjEjDqfbZxjEXySfZ3pI6PYrFzEUsgcPwKYLq
ddh8dXWyogudJtyphrXrZ0LBjx9yD6HRH5KpTMgkspg1qXeADvfUye4QMPjhgij7
2YRi9GiJaZGZf9QdS+VfEP6kj+eYWFml50HLAKHAk9xapxkH0iFFMg/kWKESADK4
RDrP7RcokPuj8Wef/DBRtunqHaJbwQSnN2FHOXTzRcrii5aADNJwg665uCZRJONj
gW0IX/+dn4PUzx1wrd5h8RsGGR40hEwP29MkqOZHHqgbTaMJjpCqaUWxOUct10OH
RC1eRda46tEEHegEcyFmZVsicR4neArGwca2dnMFQmVfhpVLSGFvoQKHLrJDt5vO
RtdCD0qN2ElTv8B3c/lNqLo2u6E+thZyjexJQ7LO9xa22S2Mp8ne9ZMnsbmZjBuW
TeixRh+92Od9ck7Kn1dJ37BeSMhC04Mf0FwM0gUAJcEUFtffckUb9+8sk/weRCMX
lQ4aj8m3r8JOU6w8m8ztBoh/aatY/U7CX6gqT/pDfqcPiKbRP1fxHpmkF/3WnuH3
KzUTyXyZcVaYL02jMLoM7JtMCIMxkb2qL32cOcqBG+W3TzktASsl2LMRnMoBXVh9
u1Ph6JCWtT4RTl975BGfaVYeSrjrEF5GvZqtVMOCT2jZzrtb28CY/qnFvw5Ugby0
fZi/76gj1lDlGuQvHE9NjFZQG8PutiAkn9/wJ3X2Nv9Sa+EPyemmMg9qUZe6p1ZN
Zrjy7nsno0jNhUzyVabB3m/YaWg81Vpcqiv8MqHw0JEfrvqLKlYU8FtjBnnyWyxZ
n2b0nGM2Xb+4fL4mtFQr1owcQNEhrja4I/ull4Fup5OIbfeHZ7oItn7AVdVKUGaX
5miZMEWoGYPuDlgakmR3yXiLtizftlBYkNcWuj1st492FHB1H1shEzaM9GYqZmPr
A9oDZEUmqt8GF273ee6o57Sv4SQcas44FYpKtA7biH1BxPxMcwFnodViYeI4R+yT
6LAK9xXWCyWrjjoT+YpZ2FYDZ7UzhPwbEvNhJ9p6X63r3RQELlfrJhlLSyVr+CHM
bjo4ts8uukaLvXilz6F5WDzZBqfankS4RibkQGAKlqJdGHvudHMmDoiJdfKVXs3O
FEt+JtcSAPJqtHVb3yu4A0sOHgwVr7SQOz5zE3eliMHeKfyXSkNwoUM3ppA/Sd2u
GFrX7zYPCfQOy/wTgAnx0g==
`protect END_PROTECTED
