`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BkbGuhOydeLV2kxulllgc7RTShA7A+wOFQaYVsH7uqFJ+jVoRFrob6eVu+kMZetD
qZV+Kuwz0r4uv2tk7qLVjxKSWAe3u1DrscfjwzH929vFWZSkLecqoYXmf7qahXYV
RAnNTHPRADAvyA3toyG+oITrAKTaf4eP5X3rdw+QPo6mx7aLluQsaYLdBCpA5r5c
NSKPp62HHUi87rpkCZB1Zfqlm+Z6mvXO/DBECRRlNrVHRDb/HrYcAh8z8axm7SK5
ux7JroGjhJZI/Vv+FsiSrptJmud7XQ07bAIK/82hZGXxDuXc/XDfo0HTisTPIJWH
3zJThY3E/B/oUbBIDEZ6oOifXQH8ycMVFCKYDfjdvFNe9SiDH8iG/V6y/Q8ZLagN
HNtiZ4B3VUekfsm5jGswGWTMn/aR0xV5g1cD1MVpTn6LZaz6qfnralR+uoK4A2uc
e3wa/fgn+Yd7PIrPlV8wRfhFsCx56qfENYuvxTelEVQZRep8CYBvol0K/N3sxavC
KaTb6Z+Fi5RWnueaXAYZ9C8qIMNpHI0xf6KBRzBSqja6Xi99+VDeb7TzlrQFylDR
CR3aHJzqyWb6GEo9o6V2U+jA8AIDmU4VsNUA0DV7opYdrj0x9DipLYiJxYaCugvl
3lfelnD9pXcaYX49OAIG6qs/dCZkXslfnbwfa8lDrnptgzD9DGahe+RxcCwHMUz1
cO9jcdiGw18s6Hi3dG+RXC83y5v6TAqRgJqOkDEb5HU=
`protect END_PROTECTED
