`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2llNNYlgHPofSrIkA22rMHTeyXoU4Sg9j0vUGcLu2LCQVkgnNH7Ej3PLaaVWwqgE
TeRgUx5IIUCYmGANH+ap7259FiG2+UJhIdVkYU0L8ESxy9kRTanIyZp+/SKBmKuN
HP4tc8T0usD+RlYzJBh6y8DtKcZUJ6J3K2T5qs+9PK1Ypbc65FXr0iO9T8FlWiQb
WQY+zyw9GIZ7mXg1lILGuIdX5fdFYe+9xvaCWRfEbG2afU946MvRIREZnsX8IyIm
ui3XSmzOaggb5rV6uSvZICTysg8I2H2No5XtFjmi1okRi2pC2W6BQ+T6CKlhJk5G
nOioKOSVzfCD+vD05imIQQqto5o3lgd/8TMqkIcMcE9JRFS/4iiyuCmhtyDRkzZ/
cLV9VtvICdiYtGqO7vwNkVXAItaoT4q1L1guOFGhiKymuqVW+fcQUjDs9UnLF8Od
5RK2/oTktmWBwCWWS6vs4g1csI9QP2zH2eckug8jsAlSzic69pIeZX5nBSwTnHjX
Xf0lrLpXWoKVGENpG+mRiJA+TulxU9GUHfaMdJPf+d/+zdVQsECCCTQlWQx/xkuV
kFGGY5GzdSePqvUSgT9y4zYTybi7PZ3UY5v9CbYg/Qc=
`protect END_PROTECTED
