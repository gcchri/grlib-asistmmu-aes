`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJpfdKLoiWUa9fJRroEMHCvUf6MM7ebn1sy+m9CcOYF2nGaWTBM0CC5p8Mu1ykqV
15yVAS5RlK98Aj6f7QmWxnQ0BYUN6ySqeK1Db46plKb/n2CdVLdy7aCgDwmK0ZB2
udPMtpKFulbYDilRQL39rJjaMkjA0UUP9mK6z/882ge87LKYCMzby7p8vCYCzlsP
65ozds11IW/yCp65Fwtk979Cyv0n6CDQA3oP0iHFBq6AzdTry1b9uYSdx/N8KR22
1VAKADPtRh7Z7dGcXJabbuIhfy+PrCaSDu8WaKIMPg8V9fTxCuWfcm6jBXTnbYzx
c56GHd/heXiuFNMjjdwXAVHOhSto8Jay5O9/FT1iE4rYBHCTTlgjb8ZRYcE8R3Mp
YuL7jYdIWSTtlZzfFLZmpkr6pIeG48Xa4k6QxGEM7yJ2WnSv28bE0zE5NmA09d+l
bqvnmtV0KBVrIQ7uXoXyL9Axe6HaVVeuIfLJ0O6RQfGB7P1AVzFPe6f+VLoWcl4g
`protect END_PROTECTED
