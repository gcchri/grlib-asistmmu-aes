`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkubsm0oBo6Kl4oHt5xHi5i5Q6OKyrhwgsaZ3Zs15mCJYMgWYe199bUIk2P6/sDX
NaKjHkbYjEJgV5UKCoQj4fURes9qPrSVFzv5aENf0+oMrmyE8LRr5+1Nj6E1g0ZT
auhnU2hBGM4xUOMvqQYNjnuwQplzDuoagTmLnZJAREDvjvJaAyXdA5nkNxifENwk
fdivMJikUZ4gBwHjUEvAPDXWH4xqRDdviaSfk/jUx8Pj9aWdqoyAfBAruni2MSx9
VlqFVIpEG1bVbM+7WJ+uZOHo07IT3UqTlWJXonLs0Q3alSQzgVuske6rDps6t6R7
rZafFgQrMLqeNo6CbNn5Todn9gmIXs/gtPycMfySYaUDQ+oLqztAZL+H06DF0gir
RbPOnVV5cwd6FyVxAk3qEvFmJeDm+btBDjX9PWbVm1ag6D9423FqjdX2rS7OiVLg
ND99sYJHc3cR/KShfuH9NXRHz3jFCjXPwEO7E5YPtzrBpE8eAqJhGLEUboFgG79D
8ieRyL6KKVHxmfTH70yBjQ1Cb37iNvci9lM0EUj4aCKtgXDdFr2dC57JLKQKwmn5
f6W8cZGxkx9er73XsUMUF1ZDbM0EBJKiclcCQuQ1eEoojV2A6t7t3sYOyAQgg/1f
5s2MUgBZzneogssIxBGURiS1m2+lSvxJ3IVbA1ogk/auUz9/KKFphCPyW78kSJb7
U+oQiESpfYRx2SAa11+psobb1GFETXviqDhkS0MsM+EP5VbAjH2Xi4XC4k3pbcgv
01HzBiBWLwPMo2knxH94AHeeFxT12lKdO51ha3XNZNb0OxktXQXGpoT98HirXzX0
wvQ5RFXy3P/UEClya4/5r6bV5omt19VfbeROMbr7yvnWEt5pbAJ3awLjMFhhTkas
oNSfKI3FJkNkAuT7x7KC7ncJDZ1Wax1em87Qb7UKWO89Vl8zlod/9T7Ib/qKGO91
aQrUD5E8eXUZZ7vaZElXow==
`protect END_PROTECTED
