`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Y+7j+F/88ZSUhKDpppH/XmuwCaASAdt2cw/ObjAaIcNcJxdZYDBKHmmiLPDh5vq
EzyQe4pPO1mEIFqXdrFKWG3uLgVn88FwTJN+/E8ftaXcBqYj2HjCu8ywEEOkY/f2
RGfiSRp+xMR4FtuV6hgvBe0IUPH79/PsgnaHys2c28Phx8MgwqY+HpCo78zgShee
H3MHrxAtM1EA1WbOsUhlbBSV+pUBXEOFe7QFLTFm6REjYm4dc4p1oavn1bBt8RHs
vSjJ21V8SnYrM7W93MpN5AWE78/2yl+orLQgA93eKARyX+GE8sgAipupqZJJ7R/l
qsLBiBZhlH9CykwOV0H4raYbGj9LLHHSUhPa84HkFagOcOs45IHrnBujiyjeDbKm
ejDAtN5KTpDdng9AVlVGNAoqugIX5W8xdukHDrFuQhDxotkJWXduKMWF7HrLJm5e
E3NrbAByM8PrsvyAS1dXiTjIrhLglW1l6bVeiV83dJYY6IUzgwhxTLAkqyWiLkjE
Vgo3TcPYdzvtqr5UxrZ3gIIZ+6rtWdu4gBYm5UK0qgau48MpQWHIfAECMzKP7s4O
`protect END_PROTECTED
