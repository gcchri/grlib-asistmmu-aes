`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DtmrystzR+Mz7VBncTmO9m/dUf8fMy15pkdOFNjqnfxAbhTmOf4wRYnlcNuHAhwO
GQBvmKOe9I95Hchv6yqOS4S3LZDpqjLa/AGZZPeTT2QRyh+9y5jxCYjwZDSRBPi/
RxJW/0H6s2crSu4jz4mCvigKk5fH62zSEU4cJEIAndkvwUvFxUoYJSGeE1E9kvLB
MaNHxQO1pA2Z/hTXioTeRKHcqlyKvY6q1aDqWsrerMyPCGTKjzNJYMPuO5vrAFAX
x5N3CmxACoxaVOSp6Xhpoce/eBmOCWW8mQi79O6rM3lQp+lQXpeznezkvuw4ls3Q
QR2IBFQt7SARXpnNjUISlsIr1ZwVdiwBVK9mjWzTiZJ1cIPhDe1CgvQciwqG8Vbh
jElu3k7GMJHrAfISWvs4Ig==
`protect END_PROTECTED
