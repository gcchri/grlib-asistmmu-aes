`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kT4U2Jw5fI0HSx+3V0c1d6y1s5nwXXGhYpmzy5PsRWd57pbFjuCh4276h+R3nVSU
jDDsuaxHD7cqmW3IasTc0Y0fMvxfRNG478eWxdZNuoN4Kdq6VoXcW9MEU+oU7qv2
J/9gVowQhujF9q2Ifb6nNs5DxPKboqW/rd0auR0TBrIkGb+5l/0HuhW3pqUuVgyD
z8dcM0GtlRJOfd7MTDgrUtrwESEQLG+NeHrdTbefViEFGKzfr1pN53Ly34VN8k8e
HZRc8zRvTS9fjG990E5JwX8asnga7DCYEzmSuQIDBAml748ZM3DTLRBQ72f0TadH
N4SLDDXN7pDIJCmsgKM4O+n5ay33msLKAtbAd+ZTRdf/25qOJWqWZUGhilw+qDNe
niZ4Bnw0G6QvyoRkgYNqiEO6IRTdOZxahplurgEbuZO5gOrBKNnd18PIgRv7D45o
W9+Ht6H0HGks9r8onyuvehNmH6VX+3a2tQiiNc6Zep/EYRO6nTla4BQLaFdj9YWM
17t9hYCW9fkwRyq+0uXy6XgcFLhdQ/SLTCESRJVTPfYaSJjaupDbCyqiLu0KHl8x
tPAPDUawMNF0NRfYxsVSqA7rmMiN10CqNFqKggmJCU89wT+O8cXECzJeKuwnLKRj
HEYm1rJKZedWO+vDS7ZQxH/Fu5yZlkqqLQduNOqKD2yEpWkcS2XlOJ5G0BGQhAYG
aDj87GkSgcpWsHic48rGg5EAgSIBRL8gYjgaQu/lK5lTdqPT7QgYJ/O6eu8h09+e
JTXMTs2utU4xAWkaBqwARCxH2MZ8n+Lol2idlSBMc2qWtWsIaF19uPeh9kXxUf/I
7ssbVy5HeIeL1lt7oxjghbZDAupsLHNUzSNGq6K8Y8N0WSLoGVN+oma4V3qAufHJ
NjKThn/rsklk/B+cl2yiMpFohd9YUz58VLoCoogjVzdWPhpKXUyXOVnAOfsOB10U
K50PpdxcbPhDfqlEFiBYYVHgP6TY664QUSaq6hftGzubUcyiHpdK5X0O+E8LCnEz
Q3ExvJYhwZxgSHsWNfzCyotnyFAjqxuhPDDkdMLeT8GeXmCxQM4MfVZdQIp+sBAX
d7IgVKTa3YBndM5/Z+e+z6mLTV0HkkOfEHJgYaFTO93bOHxijlhxOeOl0/qlT4SQ
XmaJjXknBGfJe4gdHFGlZRXa9onD5IjpFEruzXLML25S3eODHMq6C4PQhVWpmwHv
Xz28f2/SMd0RLaWxVHMDQvr378V5mhlJVyqfrn57mBoZ8OhsW3mEzVLWB5E/eBpu
RC7WOegugY5rqN8D5oA/LhWkOPmYZCG1JCoJcuwj9z6lVz1HPC5jevNw/IBXgkZt
Wu6cs9SEXqD84S6UqiY5jrBfyz/KItRi6Iv9n9hlR2smU3IMuqL5yq4K9FTP/Vk+
Pgj01xF/xgVfJo8/bcVuugxrWhQKl4dSO0HLFIoNvRlujqwj/rc/VTE5yml6s9Za
o2LxIuTr6TLwITWZlBFBJL4GAICaUq+5KyawvN56cBURYJ+8Sp2OAaUa18ubfuHv
XXfTAX1wXFMYzwq9V/OY95YKwxkTarpZdOfUJckz0AR/y1TwPod3ziBRN2RMPkmP
tAMC7BIUL3c2f0hny8n5ANFC2y9pH69HktgCJqLteFPssE0Jshtt5NiYwTyOFoi4
PfesGi2pFUfFuNm+nwWES5n+luhtTYkaKc+uaJp6eVQ2Tn1FptIvXwzE0cKXA+Q/
0wARSUJ2ruK01LT/1XJ1dTOGbf70bzKVcSFo0zNNC1tyj03IekiLh3UQHW/5LGMw
3zMBkvsc9gXLA+wO4HIbe5Lpa4pR6n9c/HaMswoKljRMPW2Yf2hraSXD6O6io1r5
WgOPGqndOGtLoFI3FufBqSIbXsxO4eq2lb2mlidySXlErZLia9IxdG9vOUmnutVm
vFWexoGg1B1KSxhurr4EeEwVgawW1xRs/rIm922BI/sCbz8dJZL+87i3rU4FEuHj
aM2CnAHrIKZbmi0PiKC66EDc5nT8M+O1j3i9gFKDTXoBHT9bSmF2iD+4yt/ggABp
HWevRKWkoFOONjS+dlB47nNWFnkmLdDMA0AfdmDELH2pw1hHNPTkcgQXIsgGeG+s
O51rvqeI8ZhsKP4N/zG+G4/zICWpOnXpP5JpJcoluh77quZcHbQ60D3oE2+YX/Ry
9ZWBacdDAAUOinkOY7F3MC/yq3+6xT/wx+FpTkC4bKPf7N/W8L9HfTeBtdrHd2KA
bbgJFSQeuGL14UJF/tmtOmH6nsMuEoUN2/wmrA0SjCdhnwMKTs8XUommUpeoCLNj
vZnwWNjGxhtxNi0vRZ+Ptl4CQU436/OTnhtwkfeY33Mp0FaSnqls19AaOv8Nte6t
7++p87OovchF0hkeNB0FFUBigPP4XFVE3EuguhgjiukfBSxj2Vksw5txjq9r7UuN
KHAcexid0oKM5pKXbPHuGREqbNyAkik49SseKedvhwilNNCSZ4cD6ErpzQYC146l
AO7cL+SEMVz73zgZzf48Jp5uwrT2RHxquTAtzfQwOchn27JNpp1z0vG8wiZ1ALbQ
ufjuyRNd/yJTRX04jN1Eluqrd7zREkulPG+FDnB3FKIOkdpWv/ERhdVcwUhb3t8T
jey0zpCt2xqiEZBl7HBDmlmkDiBqHxaabXfC3uzZxcRdzbb1etQdD1Teww74aafN
DWEBDZ1JolfPT8U4Uy7ApRtQOlgGwSJJ+0Ps3au41L97QaAnk7z/2vwwNPHyf2Ld
0R2aANMuOjDvD/wZUmphSOJktXitQc2hi3R8PfkA80rrVtoH8MsdcjT8kAqcBaBv
bKDAMdxXnCgi8EX7WWc7esr+IwKd9Xxz+ToDA88z2P5WeunWF2iods2mXViCbZ2I
o1fVS/bwyV0MxbSXYcYuXZjMzhcaKsW/vXu+4rG97OyzZxpe0ed/Bqy8Keb+QW3A
2pTY5ykUrT23gajcs59DocMcPRTXq91SmGUFKJCsOpqB5Utoc3U9WqrbGznIzgXE
iVV1EEP2xdirnMyXsQ3wJyqf2OKuoEQLZze4/I9LwQhgTeqdpTRVt2CwC91K0q/W
02ULKGupknZyJV0eOB+GEBrZxdNhneXF0amUJiE8yxZ6X04mM9I+WKYVbZblaTea
Kr1EHla2vYK9PFztLiU4hpVsFGKRwCDVxmal4jAXcVSASYEpJi2hWhHl7LLXjNGZ
MFJWV1NLO60zOSOZjALZK4eRIZ+8crkLnftj/Fa/br1qwr8BURwR/MSZZudNQdJZ
C9KP+Rv+8zCICnuGONJVrcBYVy9UuEXf2iSZ8rAEvblL/4S87srp9VoAgWQvP5xk
ZP8KpmdYlWK2K/xD4cacEvZwLjGuWpVPh2tv2Vr9DbhLmMaBZZCGyJTQVENUIfGE
Vr5JHNx8Cb0rV9OcBGPAtHZmf0wc4IrV4g1gjGTZQEC/deZN70LMpBP6H0H4O2lM
T6f/C8ap2EwmNPYhmVcjHcI5JQj1UUPG5xQzAoTnTJC/hvbqAmYZW1er8+pBrFdk
SWYONb9dpGU3V7QLxZCcmb6UbffKXgjgWBP2eDH5OtQ5c9G3gylfQfgNlay5c63l
SeLWrBzVkYBzxitRYwjYQOyEYpY4mV1Lvu1rL27PqH63QWlT9zjGPaz+GjZI3VUY
E7e+LvQetYdeHys2w8cyiIajHYwRt9BrKbciNgVupjSD2Bn6iqcwnbZKgcCW9kNF
DGwOFzOHIgEg7rXu2OXvAD9mNyjMWd3aI11/6E3X9mVEfgs5JzhE5cir1s+biBMN
792LVCDlV4zivrdtDamrvxyvUQ+Huzg4R2sZ1CuYh1OsKLKD53xZh4omhLEgRdfP
2aDKVkRW/W7ENzjmrurHNeQFOMOB/XvP+76b3mONGw07Ir0pJ87XGp8onl9xARKs
V1Ae7sqlY15BS23t6zjqdtuu//XW1NPv0bq/wpL2Gb0pCLV3UW1uzk0aTvWzqelC
yV5ce5z2ZUWj6DLqbCGGgt6R57yYefo7CjMytRP7/cAsjCUn9gvqY2DLxOQ22W1S
sFENRnJ46j2opvjcy3/jqbdpk8mszhS3ivlhX4CwauSv3Kc/PlXpFti3bKHyb4hE
eX+UtVHS7WR8lAQDnADeMhA7qqaw6aglq+2CxuvcYBRnrSNCjSHRBYdUv/DoS2vF
ZW5aYdU++wbH+vZUXLZLVGATcpqiwscZ2lDpMK3lSNtX4tzbk34FRgt0k3UXTz0k
8j1Ux9Us6fHWbsSjYYIi9zpZAsfK5c4jtKGt+9o9WOvrexTMOW4B7+sj8ZEihlTl
yWyMRX3/uwQTJbww2Ip/+X/UydGA6VMuuad7FeCm/qqYaJGmIopgqrn9fQT3vJDU
c4a0NzAvI41mVrJTO7h5XetKcY3K7I+5DlMG4xJQXCE/35c85NaYgo4sfXklq+io
yoEEftHhRuHTyI4WGvQa984cYli6mVs8EL7KXRl8/1PuAvSz5FJxQZb747KFe1Iu
lwUqD8FWw3pugnF5mUD8ObJ/w9AWGqHucNBCdak3IYUm6d/o9KEkcKBn3Nn57HbB
P5knI+4d3HHmV5YCSyBCp9DrALPTwuNmsMKk5sxi+xYjbDqK0JGlHGp7rG3gK+zM
+YC3ZBUpno7vZFjGY/hBg4LEuKqhb8eqjpsi+WwqFodtv6eD3vMkqt+rK/wo2lqP
3+GXzhrl7ycsYPamOPm926b1vjL8fXt/FMHAWQAQg3Rk8Ek38q5Fca8FLoAee1Rq
8hTJZsVLcPetb4VBClHO7XtsL4t9qjZiMD5pbNn81jVEL70isM3vrEfNsyQ1PhSm
EZkOL285d3HGgc6SZV+NKqtfflxT8VeFDszIGSQ25WKC75T+1a2i/wI6PPn1DVo0
CjwHnICG6mKsiNF1sq3CrBHE+lES8OfSh70b+lB2AbUkl0Bl0UdMBTXMomgA53+O
BVs1kFNgW/R9kq9xhc9W7bRjyFas9twuZiictUaCUhz/lWuZUEJnZCeRvRjh+y8J
/JLPYqQS+2T3BY7lgU/TwZDaIBnFJBImAIDi5AJNx+O72Q/1xQybyevuTGEmi5wj
LjsU9rmYJ98j48jOMK4oHWk44HXH+ykwa90d0luGLSDybb9L4AnqywX03Xtehn+x
aa3ZdAXUdiG1zOlKNdUpUkDxZLmyRF7ccjmvDmBi9BzQjLoRuHqs+LSao6iGAzH4
IcuVwXdX5e6sFhKJnr//gzpAwMdBPOTwp2XF8Uh1v3A9Mbjf1tITdqabN+54wZ67
YU/fKtoRSjGVjujuvOMnoMRMGiL8+GAVugCoW7l1D96CatYeRDgdBDZt/eyJ7JTt
sChf4sd1qyOJ9aeajFyVPx7rQ0YpoCSItwvgpMnVYFHB7p54PyTQ3GcOt5edTK6a
baY4WZ0MR0xyziREmKlB/zEt3CFqJ3ME0EPZuPOqOxcdSGl+3VcTB78ejwWUuVtK
31RTszGI3bi4LytCcvCFQ/VDqIfUkvWHfoZotQvYm3/PtyVPjLV/fYLU1/POxJpp
Tm2j6iY8n1x9XT7904/3z7WIvSrqJaIr/yN2DyLO9zi9twLAiXkRMDbqLWyOO4Ry
PJnsU18zadXPTaQ9NPyMuZ7nXcogxsMBwaUBogY2OemOJVqZFO1PRjmAxaF0quWU
SO5k1Gr9UrvIwgTgyptSUJC09b6iu+6k0HiEv44QbLmusGgvcicH4Pav/f+YZPF7
Kogfz2UUUz/jK+vNXrBxUCxSeRi5T/pJsScHH6ki1SiVRhUONDgmQvYj0iuNCICx
nYD7gitVKeF6R0T8F1KdMojX5kA3y8yPsSJsLpNuxJKgzAmFQHo3Au7Sj4ofvCMp
28RapAw48jumchOHYoqgsg2uLey7CxwGmt1a0/Vc0ZSi+BeQcZotwe9bEnKSHEnt
386EiUh7ftoxGECeZmQYyUNb2iQ3ZCUmX5GrVkF9kd5B+v3RADOWMycbvp8JCGl0
eYqic0Zc+EFhR2mxcXTPPdRJMkna0qq25zFEY6ej9O1oa77Ahhzj92VP5IaHsqUr
URaAlYh1BzLQHDk7pQaxSD+fK9jqNMi9FWFFhY9k2Z5N10CkGeN0VXBUSmVzmwEK
uL+oVJ3FTU9hH//TdELX0Mi9rHM9tOXaeolpSQJ0qRrP0soeRLReno+kB4zlKeEp
BPgp8dpoCFG611v9JLNmzhwSCNGCz5aXq9nBoRivjaEB7m7rOzPPL72vAtGqJUDi
zDJeK/Qc4CrtrUFzeu59q70hoje09aXB3zDpSXa8JTM1b7E3EA7Y5fXlWt+vEX4B
t1Ik6X7fpjGMlWYCh3xYEVSPd75UTHqN2Wmq0CbRfq+xyPeImhEMMEu2b7ujhQSS
6IvKm7tyZvuB8wXE8W2pSUSTyel3VfHLGi9S7xrpiVYKKGzhx/lQ0xQHsH/960FK
AkFL+6inBNv93QdeyDaf6Z3UTbP/KUGLFuQvVt0/x2NnKDEX6CMpLbfVJO2AmulT
cJBpEWe8j67eDs8SRbZJOjc3VQ3cr/ms0Qb0ymbd3JdsgMd4FDcA/GXAVgsWrWJO
QNPqZ/NqLYy4D4YWYOxNhnY6oOdGDzATg8EaGBSNm7r6VYZFR35mWaCSJmp7Jovu
DItGN/w7CYQZu36z3bMb0PJPNmg1OhlSkI+PLIXL/oH7W3TKt24GSXXLHGcFSshO
QGzgLPMrNsnqjy9fq6f3jp0DC7KNrlCRlXnloNtVKkvs8pPrhKRvSPKQRWDfvSBi
Vbl9LkONlzL9Oyy/ml9cLJ6uag5WftGMEXdRQHOkfpE0oeRPSeSSKtaPbhe+gWGi
M8dAOJamYaSD1j1HGMXw0MLUMklBrnbvkt5bmoW0N9ynKMM87QGZTzBlonhGa9TZ
CAUwO6+u4hFdN5qaI7VZMTM2oKWUDeXd4yhxa9+MyuKE4UCMp6NmKLkeGTnFA53Y
IIg4tLjpYue9sS0KXmb/8auW7BYWWSn5yZPTPyrCR7mW+5325cLlDFrJ/nwFJAEY
hhBcjd7IsAOlVAgoqtueBRdZAIZGwFd/JnNNq9omj8YispZX5oy3AW6ZdhP7Vc6C
9JoeyLfJRhMslQR5YUFQ8MQkpFTC1s2bVFzh8NwHI1KhXcSrSA8XeGXnpE6LNWgi
wE2C7N4B9AN8KYltNMMciYfjoeCbhgagEPXEQlsMChG1KUex5oJ9Yl21wL5+YmoL
NEbNyhjZwHJvOyfl8n62+w9BnR3SNXkO2RvEiJpYMZFQ1PcuS3LP1pyM2N6zG993
W79W/kX/4nbIKafHOP3aQPnOLMI7Ax7BXhcKhfCFfxhB2o4n92h5LUfrnFYp8Sw+
bdt1HCsPqasQLcKG+lNBIQ0GpgOr/BllZuKRto4wgHn1VvifUoa3jJuB7TQ93KH5
1aTjDrkTAIwwflvS15uObyCjV7yOoSI7l+Ko9I502ihFUEtppXL706S2xREveoTn
i+fEIb6ve3cKI4k1nmoF/KIoHw9IUMFIILLl0v2AtYBq7fiElwtK/9YcSwf/9RSV
zdsiv1HWVgK+WZptFUfEeF55PGiDWQnNER/JNCvUS4uULHujPW9DbWRPic3WXjtA
vYiwNAy7s5mGOyJ6A1eM8rgGR0H5O0VtvZkGwE3I+nPS+LxsTBUuTmNec5IiFxu9
2+Noqmfmb5s5CjKVrmYvUNYUnxTZjQ1cJJ6qYwTGUlD654Xu4Nk7figFCFRxvVQH
RtUTGGdXTG4a/tgMi92jyBdN81dlRLelkp0jjQol5FA35p0P46uABPuAflDenraB
duEUA9FKXaztr6Il54aoq5dV/zU89B4sFB5c7vYxFsMa5kIiRuSLJr3+tUe4MfoQ
hWxYo76rwB3v9Gh9PAdeL11fx2X1wmWYxfAcK4lZfRNXsJQkq5Xi0BD3XvL/hD4Y
ksEcFeSgvILNRCfEocmIdIpHppZk3c6RaO0bRpXDxrs+cG5Uv9tvE3R1gs2/4Azf
zRiuNRPcYTQxAV32akb6ws7MY9CmNHp92ggK+1GRx0txqL4lfEN4zwgakowuUuYN
qWoa+WtM/yo0lWV5tVzbOo6gBQnOl9bbxtbJ30eNLNHzkzgX9Z+5bnz3rvARX0wK
7YO1dM+CxxdcMvL6rJFDpfmxOXHUZrVrB+XzzCs+aFT3cC/6+4iiE5r35+48b/di
5XYZtKs5Je3NPaVhwpGox1XsmO5BnGj+XtUzgXpDrWFg0MX3aHA3xp80Wi++sWZ7
G8ZhLnS3jNCns22dOiAcf8V1nU69cUGLX5cBqBAXrRNCAKmpHpHi6Gl8Gdi9k9O+
rQZx6TX9nYpLM7d7+i+VE1Gi9mebJ9KjdXsG6Q2L6HM0ZAYDH/d9BEOYgotLi508
zWRzX1r7Yu/0No23AC4TpCQp/99MN8WTfv/0XJTwJtKGva3ZXalFgYbBh18kOqqF
s3Fl+27kslOH3XRVrQhDY08HoLInoBhETqD1j+V9lswngeWbWBcFHvLLsdJ6uquY
KTIHFqp78iRBDyyfe47/ilS2GcpMWU5+Zte6243iOeAd2mP9VfQZyWLVn89dyPo/
MN34UdN/HfUIj/ehgqXgfKX4tqK8qEjJ5mJrFQZKJOPH0DDmLOTpXUlWVHIan1oW
3kEBrx96PR4usgUTEzCWr7A1Dv3u7AmlNPqTyZrhHTSZqUHSHey6nibqNE08YdBq
Dl5buIqAd36NbZx0+axvk5ojcifnYRMffkSAP+thwgrZKpRMJ6Ht58lFpCFCh6Oe
ri14cHl/cDRGiA+R/jYM3IziDRyP+lusOT5bnKautk4caTS2b08IoWteuI5E5Zya
Bb+SmysE4sJ3wFDbjXQVr9AzVQnZ7q82Pgjpcb7sVRzyf/zJ72agV8R9UeR5dDvE
7f2Xd4qdc0CLJjThiCSoU6BR+1h1RKBFcmwWbG7eFipKCOK1fnZgoykpzQTxYKrZ
NJRZ5MxlmcKKXBcIuUF1Hjxcmt/hHweoYzai9RIY5CKZLRJnHK983VZtwDRWzc+I
DWM45yUtRVtYiGshVUELW3U7wknLfs3xb9sVfyuEwxRNB3quz9Oyd8+zTXwVjs7k
NiiJGO+HCqFY47PPLK0FOaeFi3V8mPA05kyg7kjThGjXIjUwqhAqLsC3bB7wZst6
azBpKsTlFdm+qh2lt6RP4NaecKCHbsEap/vPnyrhWROYPGX8/+vRzsQQvGgzfqBO
JWyxDICv6atcYu5F5mxidAl8sZ7dBAiOvKJrIJvdvMwjx4x4mhVZm1yniJLhjtLG
izUsl8MXy4soXfwGgYqjEdiHr2BvgSYE6A/IaBkf2bcLgj+Q5aZZ+V279a1VgORC
Zl1I3QApg6P/pP1OSNC3WsCgrjUMAAb5GeJCdhim/EfOFbw7Nq9+tNHh0LCSwFsC
uoXZFERtl1eUwws6cOShPtMyxSyeWni2PamZpPtrqqa/kqR3qtQ+Q0R0ad2KHNS2
yaemttQRqjJymdG+903v4OjFzAlGjWTX1sznJXvBCAgROLd38iwS3tD58Xx/ge3O
Nocdra0L3oHc4kSuEtHX8nrdq2ukyUgsgAYGfyTrJJGnT0BpeVlP0b5BQ7OUcYtW
KcMZ3qVe+aXIxOZLxZ0HApV/TsTf+7EFFoYjJn0KIwvK73dvbIj+jw4YVTQBNMJl
aJ3pWwUQyA+91mjSUmGleMuwjxC3GQIPOQ1dlDPt4UFChjf7xLVT8G5yng67VUWN
HaTCFGEuTO44RgIwOtkxk5SIyfHCAtHadcTP/VKvPw5Bc4RXnP7dbezmmpEibIyO
NNV0S2y0iR0b7xcMMAPDwtov6GzXZIcMBtooxC6AWpyLw3ILKPExtmcIQ0jbd01q
xrKHzSqgQFbQswVfwzq2b3FT1x/j1K4pbT4vH99k0evQFkcqQDhAk922FMcc1pVF
hRrkmut+9C8LlX9uUf/46raUMVYumxaf96jQ+FuMowwJ82NKCERq5nzRn8rHQB2+
YfT8pkYAdKM9Wwv5ZSbpr5OY7exvt9RZrknQv2kXModK5i9ZdrTSxF37i33uzy3L
jTRyBC60bGw+02KdwbY7pIDZsHPEvTwJ0e8ua9wrMC3JLZijI2ytIvieaUbJGzNB
qnirrnAZKPGbnnq6U6fPiXh/AUWXulmdFdlz2rO5r/iK5/Zdckue3pkqx1JPpLFO
JllkWoiNpt+44roEF2SNsSJXQHlevL3Xww05R8ApNsdvGgvo/sZKanMUgALWvg9G
UtBh3lZTKm7BakyT6wSdjevtby84Tnuc5qfbx/tCcjB6Yu0d4dR207R/S+RfWVgX
9dJCnMg8w8UPuLRwo1NTuEx/0yY0FQmwJclNoYHh48sugjEWjyvSoHwoGqhQyN+G
6L0zrO6tfsAFsdz3Y7Nfuk+71eAtFBvR0o0Gb+XfcJFGI0fvjzyhFrFKxalP+P/K
FDHf5qY+a5vO5CKm+muFgpzi2dwCDUn9+C8VqQnL2XnBLXvpnUbgJkjdw1eRbozX
5SAqTzDnYidIrJgy48cTS4OjCLnS9NFn8awyNWwdQJS1oT7Y0D2ZAHKK83UAy6fP
1//1+7AkSUvBykhyGp7exh5y0dIFI3IwilzSAHj5Pmy7oD/4iWOvzB6U221wsAck
5PoCBHXyIPGT/buQ66AzW6pMXx/WDT55lXppAYIqyBqqUsRgdcJHf7E8rXSh/W+w
z8nB7tEvGqp7lZ8chXnccrRD/5UgaocS5pRHt99p9SBpk6AkiK5T3XR96Wgjd5BE
Zutu7DDA5vDcviLXBbG8yMfJ0pLY3fY4SUlAqzcSdVtX8YAtwTFkKeRE+rU0Ii6y
trpRa1XsliwuiQhT/0iUHK2x6NbIbWPSgI12fU0SuNZ0zRM+nNWtykOD4MfDNNwb
EqPO+MayTJ5sCsRF+BuL89xyzbehxr++TLPfXQif0r3pQZVhglu1uBSHmxDD5DZy
Ow/rB9J8v+Yq7nIycrOvraZQGHqxsIh1vTGB8WPjvS9eXE6KJhRHqJDA9G7gqxc/
mxP1RWy2O0l52/uRMXHWUTjjk+5Yo/eWP07Vi8iA6jgM/5eOBAJ9YeYsVZZTv9uQ
zkGGFUpicM+bryKmq8XJ/0Ki+vTi1t5U5J3GkjXE70nqKniYNBBeG7AySyCCfBFq
5WukwMinxW7dCOlq1jOXQ3NoEnmIUI778zuECt+rfchNhBIbPY0m1IqTXDtUi5Hv
IjkvRxy8+Wl2pWMCYCOEA2qap8A3iEL2ZO+eg2UXZ7Nk84VyJPl9mCUS2H7UOtpS
1uhNnnKCi0PZf8lwEJIHl31WHtxce6D+np1ATgnnMBkYTB2ZijdwHcGerYPw2FAr
3qMssDvY8uauu1sF+y3z8nAQwO96PoVagr1gs2sbD0ki3eC+2jL4bYRYyaMRQZjU
0SbfPSNjTFtABOd8vQ8BosDr+THmJoD07na1tUdag6j3XKxLsJkHaxXbhbY9yQdj
bX5fMav0QNd5+1UKTw4vZwbhjUNB46VMmXw73ivu7RKjTwlcOMvR3vBV1WFiIOD+
GpXmBfzJI5zunPg+raWxCRmJH5yggi5vRaqljrHGNQoN81uKqVf90pJtME3vVNNv
mK1yCY33thqPIGJ26kGgNP3pZVm0hhgUswFf02JVw4adH/2XIOaUKa/SgvZS9JiQ
Rory9bX1B8rNjGju3j2PRbk/1qoI6SZRvLBbzU3kmGS6VSLkvVtpZcPjO9LtjN+5
yumebxd1bM3kOjPzTHGbvCaUoL7eOBU685ZYYHkSFLRHlDWO9AX0Y1l+phVtctxD
YJBXwyzjnz9G8hHzYKWZ6MOJZCIU2bK5JSlf4zC2myzOCRZLHDpuEeH4I/H34781
/Fv9aryhqreg/2xoxqjkr7zDoDc/fvwv7/OQLG7t8M8/K/E8Z/zLf0JDTCdGytsR
bks6EBsZhJ8zzaJzBIusvyarKi+N2b3dT8R4p+FKnQY=
`protect END_PROTECTED
