`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4AOZIGLu+NCN4e4s4r/hgpy/tmR1exjGaR9f5xnpDOBUUHqSXUkKKdvxofq4sam
CWx81fCqULYw+7mDD/1GApj1cBjz+hMpLa7+vfBpdS4leQy8+BLmn7ZH8w9CaDIB
CkMP6nnabM+U1aVvz1Ah2l69PgF1kkTmwRa9tVqXWUXDuY4dRddRudCZmvQ9Qpps
SrwozCFe0jBfaHhfOsVBmBiJ5Hr+HCCMzJ4QGm9MVWiAk2kUZK7IGBamsgk5D18s
IMOwEOSvM1/o/aKamGvAz5UcoWd6zHHl5epQ4lGFbMxIcUde5m46v/2EHynqpp39
meQWQ8534Yj7ftMML+KmcQ==
`protect END_PROTECTED
