`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzT1mKix+XnsXtMLFFDhn/osqGqm6p28PlGawudZJr3BTYGV4Q5R0z1FOPE/Hl6U
dwIqQpyIAfRJVsQeySZRt1w636sTQiktaLweUhojkueguc8ljQg2wUenb96Mbyad
QriTCvPkBn80xRmfq69jc3HAotUsWycBfvQA39711QW9fdz/howpGzVlF6NO/VAu
AUiYNAjnndJ3t0VJJkDbyPGX33WdIQ4pgIZPtsW3xo0WzD0gutdHu83IuXTN3rd2
eott8uBrsVY3bMTYzuxOuiZvyQllBDQcrbtafdBrE6/M9hSYDv0V5/DvitYiCXzU
m0JSAUo/gkcYLekStj0TxzWoH1jOJYvbRIX5Rgxs1myumE8yinyRdh+xtZz1siIX
K+16WBvpuFqs2cLoeulQipniRAY+3UbRb28P9H0vsjTZm9Xci9gv+QpaTwYj+npQ
w+6OsoYTolQqDLGpRDT9Sbqgo+Ks1A/mTiXKmRkFCklqHtebUAso9eMPTo613PFV
`protect END_PROTECTED
