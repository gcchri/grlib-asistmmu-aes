`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mfy2f4bfe3TA1B3IFZ7/+CwZuIeLBZ5NM/9hXa/mv5wydpX94GEIkJt+1HEVo9Pq
Uusc0+XRIYdImyuImpq2gDRXlFKpvqbjmcEVrIuinPeOea6W+Pg1LHAxXmYPxp7Y
LJX5RrDk8cdsZ6Yc+g1Yf7YkYh6bic/gZxzxqlSOQ8TgMIoqqcDPlmZeXUaucjh5
+loQXYZrZZvthRzTr44nV5nIdMkbHAu8S8fZOQJCiQiJqf0+PGZ31eKpYQPE6mP2
cXWdl2GaPTiXuCDJOzVOAQPm3inldLoiVefVnhY4QzE8+EkBqtKuaNhMK/A6lgsm
oKLRgU1xZ2IoTeZ7++1Abg==
`protect END_PROTECTED
