`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBNX00RXepcUVh0RpMuy9N6BfBqdvtOtU25Lmnk+3YYDLIzYvBm6M3loEcYieoVV
nZJnBiYIIra34rd65lRUipYCNTkM7PlQLieWsKUFuSf0gRB1NfuRh+DluOIZjjzN
8TPL8sDd7V+F/Ay9ic3VDmUrw/RbADXS1wfsmuoxiQ/tEdwMM+OfBM2g0CTvSxqn
tXUqld91AUC93WZrkDlHNz/PRSdi13vo2Jwz/JhdMCHVuKEPBn7UfZiu/hh285L3
/ij83uXDd/vh0P2lJ7qdc2lap4DP/7t7x99qdqD0xdTljlNpWGtnzLj9eMqwVcZV
tHCUV7PI/g+TowB1dN2G81fu8AyrmEk/Jv8yVQPZ0srqa07EWcANh7n68pcg+PKX
TwQ6hW2uaiHn3KL7Pg3Vvw==
`protect END_PROTECTED
