`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3vc9SZtwRbcF0InGb+QxrPGG3LPYgY3lVjv2XXi77atyKXOBtSSUwiWVFtHMeET
zIvaF4YoOa3p9PjF0U55rlGiiax6oK3Gzq8VZ0oYk96W6JWvDWeXMRyWN8YcjXxc
ectgymrNBu9Z+PDoYI66PjnVZhmFS722mr5B+W5ONbscRNt2ZnxePE0ECcU2jEVm
6qpJzsBYvDHcOwYx9r5iFDq7Y9Q8kc4c2vmd4SAZKSdJEvh9PaXTcyN4CiSZ2r2l
nX4lZWc3p6agwgbh7VJ/ETvq4Zw/o13tM/07qa/h7HuOcQtMuQ+FFI4tXv222dt3
FGCi0CsMfR6W2Xhg1mTGV64Sl7R3rYM7aIaoowAqWDEO/MwK8VpEzNsFzJxDKSlj
2W2RWnkSrIC+x8XYVkQIlA99hptTys73NYiJLm3MNg2a2D6GMimKj6DgehYeb3S6
fzqx6O5qYisVpn4JalTGogeotCLcQYBfjxklRnuf60pWLZ0YVsd7zj7CTnH1cOuB
`protect END_PROTECTED
