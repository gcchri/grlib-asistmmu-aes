`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2XKKs79NxhcmgeiUEdRT/fhDKLRjPXktHMGYqDNN+QiB45rQWXvSmfUExAyuI14
siYR9vg2w3zB4xrM3XWCCH2PVO5EuxPkSQCf2qWRsr3R12Dt2YLKDGnCRxMLQtc8
kYa9L96cb8eLuIVOQExePSuGyBI8P+KE9NSaUQi908i4tVpedfsrM/NOwpibXhYu
+n/t4NIYvnR81n4sbTXFCI7PyHf3G7GXp+n6HfJN1ZpEVgY1ZF5/A+PtDc2QCgki
chS/pgrHEwrG9RxxBb8Myfil7hsq5COK1+F48F/MVtUBg7o/BeA2kwuZD9EdWeCC
TW9ebNH3flqI301zdJwwC4Mmp5qSCY5yVpevEAAxgBETOxarNhf6jUhy73jKBW+3
`protect END_PROTECTED
