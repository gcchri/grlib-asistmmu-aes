`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hplGa/KxrDvOWat13I54m+JFoO75Re++NtWLsKYsh/c1ubnnSfJtDceyzyMZLdaF
n+zYthNZeVk/2Ht39YiI2n241FsDy4LmtMQEtA5JWZJKttROEa+ggUkC7yAjeZTj
59yp7cCNggDw6AhhlSif9GZ+oKTYYl7MZsr0vxAM4GAJwnV/N4BwoZPOUWhv+B1q
ntubaLxDf8htNoBrZ4GZm/bWaLPswpMjmscWGNZ5IyFkUl6eMQqKzZtpWYKyzmK/
5gEXhL2NjQC73TL51i6ncdmtZcXXAMc97LI+qbRsI22PeiQfqCC26XwHsgr3Owf0
TwLmFRUKRr+vCNUy1N/rXJDgAAwQ1Q+t66Fxl1OcT3zWc5yi2VMSLugvq87puKZT
55F4/PfntFkiXleSHvModAtObr/6j/erR/+kRyncQ41pl0ilk6xcbk6WQYLG8wi7
uYlif6GBeTuyMxWzMxN+BY3Xd6MTY3GLzRLdx3Ghh2afuxQ9FGhNpHzui0+ambH3
L6nD8qS9KegfOMN+zyC1UKZxrXtAqQQuY/IMquFMnq0WUorgXRPYK5VfC0tUM1tm
vl5ujNBjxMd7+oBjRgCMZMRVs3u+r/2YeWG2LX2n9og=
`protect END_PROTECTED
