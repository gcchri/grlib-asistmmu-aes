`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNVIGFQVD4K/rzy/eRVxgNJP214qJi/QZo60sk5lVRS3Y+gOMgighTZsZNpuCEjh
SJstNPL+OdRHc1ljUWBcNWpqEEhxhfnyOV/pNjTr7w+7YbaNdciQber8tPqCoHdl
hXfgUs/h9wJZYOCinM8FuyDrgkI82DIZwhsWEjkyHDwvl4vCg2s54Z21GbfC/cib
Tfcfkt7iTqwNL8DUKau9+8Zl39ghM6leqXV2ZXpKx2W+F/E51UTC10GWehj42IBg
Y5dj5Cm6HDnO6W5gUF3E0g8ctt48iPrJ1hwrUbJ9e8LGMblUXMUGbzDr+BxVR5LT
159UZyQ3WhobCwt7puzRshxNXAqdA3XA9ELfT2le/fNfrtu8sr5uW/MEHChJjHz2
UMqPtLGj/bCzrbPuWI3v8P3uR2pkyoWic9M+pkOmykcjsN1suLHabsnSjmQ6RkzL
Ajf3wM4m1KFniA3t4lDskbxQFDmsQCpVa8c7fT7nWQYfCJpINhYm4b0SHrniYREw
P7sU9yk3XRYvuo3qUbrRXV3SXGgRV0y0iXo5RdaJIQ0ldJpAl33ctXoRqnxXRgoh
`protect END_PROTECTED
