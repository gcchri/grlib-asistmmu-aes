`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UT3D1TGXbByypDyIuWgiqApZGBka2LR5DGzTwN3KkszAAXse2DjqoFeNc/SZxWJT
ZobQwqenrxv2TksdH6ZEZUI4nZ7rJeVlRiQJNqrLsoZeUViHaD6Lm3F3LhdvR36X
4RYH4eGpALYb+FXgbJQ95ZGjFl2+HzD35jGmDnblLBHv7h8PhnFHbO2OhqYC+H9F
ZFF5zWKduKoRjo8x1+qKHFrWAwoI+pBl2+MuYOpDHW1pwml+xHOLkPvq7xGMGMvs
dl3+wOi2jxLs/0mtnwWwKcxQd0nmeVwMhlS0j4HFl9Xwc/fDY6ytkgn1tttYlykf
lkCTaH9e3Dig8Us9xA8F9C6owFnNOYKdxNGPniLq5H8E5b239+tS0xCbj4ilZKKy
AC25DQvjkV3l+ke9eZzWuUMvZ1tZJ8QFDem3FJeahDGnL7PFYYhVo1WpHXn8NVh9
CszRrZp8RReKqQPYYqQNU3JpuHFkLEhWw3Q/2TwBNokfWG8uBf/9eE9iR3jWN3d0
cGxiMoS2yBKehLm1WmD8voX+iNEStSBzetTgSZnm7QVILl5MZyt1IV/DjzhMB8Bo
sZRo1ql5SbWTc4vWbMzadmd+9e/XfuCO22avpOKXAgPek5HWz7Pt7UGyqVKo6Jrx
L/wpvG9wy2jQUpEoNrb7d+m/t8LhtPSKThJ/jtziwaENE2v64h68VjVRvTF4hONO
tmMY8VQsfJGCFZ06KAE39vxyM7TosAG9PK/ya0JtHWdiGFdVyNKM5K0E+8sP4+BQ
y9L9p1Yzlo4RuqoIEifF73koJ/475CDnvMjnjse3GbdYksZKnHmRygMueTTSs4I4
2WI90O9KIuGkPYx8PfYJnZhPqsqFo6VfvWI+IMtoN66zXQ7vt/wYl5WQNLxhjaP0
mddIUhb4ORUbLkS58v5R75nZdkxun7MvyqcLY78P4KHgsNaU1zxzDEOFOGQChwZe
QxdigB7yCdTF4zMIQZhJBRvJAdWl3AA2SIYdqDPrvFMYcngsYNKgrrbPno9nIH+p
7jr1ZKXBHdnCMQuihPHAdFSDDP3OLvLlHe+oTCgIGDeQczqH/dG460ftg1byKAS+
8VlisAISv5Kf214jwZinwCvPEjyX0akiSNlziM1oVeARf63OiyH73uHeJju/fRjq
0PnSDQI0vT7uR1j1CxM/7e0oaFA59pAI2OBIYPGLrD3SmwihgZr6Uh7ffVZI+b0N
pIGrGEG0XB1tKP3VVSGhhOihApIoEECE1Dplk4+VdQYMu3AxNKTbOCvRXdaKNwUZ
hefCujHhXSwS+Z0oerPnW1ToRKuqIJKPHl/70ikY1Ghg6lG0IeiU2sZREWeH/bxy
/OUcL+3Ra/euatudNoOke86HoSTchMuF64d1rtaHGcVt8o5t1x57AZ71BRoCY/v6
qLxDYrNiVt7rWl6MMDvZoftJxNrFAEIcuy+QGChgQSMNmdbuuvBJZakLKV6VZPpX
XsV2BuoeNIpPkItcFu2MdcCOoVDlHKeHzj5h1/Cg8l4JaB7e3E+4V6cOtQGYrCGS
8v0KTgqg5zKENy5ScJ0L2MZbocN0NUpUsekGbaha6eF15I/lmWsyqO0sJDKfyozd
smztWz5agjLQ0D6msDcZvn6zgsA2dONni2q8cb4PenmUtU/i2hNWnGxSshkRK92J
Uy0blvB11j5NL3ThyfWP5g==
`protect END_PROTECTED
