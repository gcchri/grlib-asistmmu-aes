`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3eJq2rJpxI/XlQBgSX+mPk3HwlitBKqmNMi6Ey2NcLoYwku5S9oHcjP5wk9DtEL7
bKkhtd52HyOLo43iTKj8vVyt7invKlE2r3RKCzj+d/eIbXqXuRKGMjOwjbALllPS
MALgIdlWPk4KgKU5MqyxP5NNepO31xVeceC5At2ERHsaA7lCvXjHuQlDIOJLru8y
cBEh7L660y2/3bTLcaYWwaUI3d2tUBhsCSsNN9rcDbrkWozQveR22YX9EnGAlJP7
hNldpNEX/9JBAtOdvySCZMPOeBImVzLW3GYzKfonRQHSW0HskLYnNx7nF7bl6bLh
cPE4ZxviM5GDWwADd0M9PcJaviQAf0lSh+CsglnXgL4KQNjXGF9piejWN+5QjQqa
paotKHFy2x2VwOla0Vxhm7grv9e1ga6G+MVPj9AMNRqs1K2TivgfyjTYzPLh4l4V
vwYrMIfyMScxeQ07Q+2w/v0NUXUTMYzK3nl3AVk6hqHXmCps6QFGZI8aIf10vd33
`protect END_PROTECTED
