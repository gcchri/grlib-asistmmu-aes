`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBq9CVdqa9mypQ3COcihTWR33ME8umIKNd61gS8OClfok//0ttTxS/6d+AOHiYJt
FU54l1+zf8tPr8Nd7Q5AOaNFl67BV7/+yXHF+1kKdnoz1WUY/y72lLc+5Cqki9OD
5jnFIVhvrox7nJrB1cavgvIxmGOeqD+2PMQamBPq9UYvtfIf0EojWr27elU0/89W
ALHI2o/lU7f5G0J4PrKtsOB88ck5Y8GyODMTXM/QzuchvvDVesweHAdmwsA6Xjzp
8/WQIVMslhs7RhnqhWdnUQRfwmfYNXGzIS1KIVwXQtpJqI4T7NASYsRDEvaH6rqE
iywMuAwENNqWBBIRrh+9q1TEfbcE/n1Tfb17fuUKcgxuHl6pTNBOVetgHb1C02cF
1XUXhwW2giDeV5wYX/WByC3fq8gjYzKVNBqT+X1Hzcj79d1ae1CE4hRCXd+mKChH
`protect END_PROTECTED
