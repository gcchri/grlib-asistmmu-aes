`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mY7MVysvoVdxaTYL2QA4JCivrMH/7w7hc8UE3SJSpR99CEoseVRu31KQJ0+X+YIF
mRGt9mqvaE+VzzHDfseUL2fOt0X1RnAkbTZaixHlU9yhqspVC1+Kq7WvPa9aJyPA
XPaHDeT8dCu5i1uAeT4PWSrOBQk4o72ufZAMGNzChBHCo5HvXu9pTUK4ixrYuKGm
X6rcLNNG1fF6q6nD8nyLEZlb1p2j3hk89yjeSIYq0KNtqKSWDY3Ie/rlV4PLX7zc
JDHsLVavWFJaMOtEkjNaFhniBblV1LejAdM3OVcFE6XO9HUKqng4IraEL+ulKieX
eb6RWvxjPfQYbRIfcxtmi6+LD/MAadtmqacp/ZPcQ591Cd15mOC18ZXgIKS6fhrw
/vWu3r7DP0ouIbogDO5B3qY7SrW1RsAvf/mioQlAVnprHYqHNY1BsOZ/iTd27iRU
XPgNSnkVu7VrmX37m9GDm3ST3sl5gJz+qD6igokddYkb6y2x7gNyll7Spwl88F46
WzEj//8uaBU9pD3lDw6mMDVOocd+zM3TsHGomtUgwkLLpjO+N7MeEb+dhCuP9dhD
QeQZI8L7vVDNli/G2gkiI9PGoEkyFgZXLPIcSdZzl8vXHaNAgbElMWdiN/2APGV1
V9Qvcup3Hmj8t8FeVdmHH/k5AHvd/k4VqdBQp3HaU3JxTW1hwuCJQCisjMx+ugdB
XImzKjVjay5kVHm7COtsoQDH3QZGfCIw2IP1UlirXF36NvdpzOlsxr9RTjeWpiMt
c/f9FmeEaciIuRrV6NA8pxvEFKIvn2BAi03b2YWlZmY=
`protect END_PROTECTED
