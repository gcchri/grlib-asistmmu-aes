`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
75NfGDcr4fE7cW0qjVek6w35SW2I7PgaQF1BmpLKtnDcKxRcW8liCCG0C3wNmEhc
Ex48ZhzDAKAZlgxeZc/FFbfPegy8HMCNW68IyOWUfx2Ls1iiAVbD46KD+uU/0PNj
3DpaGmN6TbvuuKusIgK+axjjuthFV1daz2pb4AB8jff/5RMcmCqDPorfdAIOpJtL
qe0u99xUIGaxqmFcbfRnAzz06dL489LVuCbQAhA0U0I7VXSCaIDr+CNaJGeFLWTh
rpVixayY0IKky7K5nyS0yTljM6yYLDMWIUuz2XEjLUBGulsGV3Qy8JQbvBAnBRht
FiWZZQByWxTMntFLeOJ1rluVAzP3i5DdC+hgQzRjBYDb7OiTzN/V8POvpLgq8Ljo
RpU3UNTfKbItgvtNuSRot7tgkUdpx574nFcmnwmLL1RyVpYU87/LATFhI7mydnn5
YLFl5oU0BDYLcnxw1RgiKNhFAtm8itHa0YI3wPNnmX6xnyW50TBtSeDWZmrzbx8W
t2q80IttEFNoz2mpXIxQe6uG/IPFxO7QTkCrzU+ZfnqNGIkItz4AFlLPC4Vd9Vcu
fH074GT6MmLXhFIaGa+/XWnolN8rSSxlnVWDRtv6SMLSiXGuGu3kaDWNbXa9mpw8
2/x7DIsj2tQopZVNHGuDgfW7MDIM3mHLAI+Y9MnF2Brz28h4JilT+dtwvMxl0qHt
c/0OHBKxt+4Ltjl278+X4bv/iZK4GCq3Eh4KsNPr9SQ+kxPgdPfYGA5+EaaXRKMk
4g6tjQrxU+KxnvZpW3KWelmKB5R0QsFbO+1VHNtgFF0bTRJV4xfZapCnnMdLDKkU
r9LlQEHEm7HxVFscq+teXi6kMV2RUe6pdnmD6J3yv4h6FZBOs01zysoxoV4k0aqK
Ec5bf00RZ4mYBsCvXPXTj1WIao9eGSgpSrJKCbQrLnkxIsVACuZDqDH00TA/8yxw
7pmJrDQ5s0dLO93K12+X5w==
`protect END_PROTECTED
