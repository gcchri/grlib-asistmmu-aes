`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YeH5NGmZQlvBwM1frRLlY3o6n2TDJSyJYfOpJu1DlFNsD0JPCGNXrVoRXKL/iMaC
KP8OguZRpOWDnOo1gmGPfA328mDKPUmyMsKWAfGySEEoVpHeXmzjvc+BPwLsNKTR
MAG//2VVXBT4QR2uwfNxyRIY8DDgtMaDEaxfb7YntzRVXaLr6zl9jo8qUvSxs79E
QG7rYzQg5Rs7c5hC4edQqkWoxr5fW5eGoi5ie672/kKyg1oWkAlxg1dByusINgi7
z/kD2SwZHNqUhr1GIuL5fTPcYMHeWgCxNYKvSuGaw5quhboEv9l3fGj2Tjt/bN8M
yaibh/pB63icI7e8gU+dbMr3lSAX5YOfxFskvZROBGJDM9bpQVFQMUaEmFv1rSB2
bz4EOR+EVmotwvhxTJt/6aJ3tArjut9TWvYSrLo3X3XkCSkcKBCz5LAeV5XR/igQ
WlxlU5zc/+fEd7b8p2HyzNhL8ESli4qPpFY43iCzsuPZkCmeT+Os0leM9B+c2cP5
HlbVjiHONdBP8ZTRUOMivlIUn/x6cqNx2/rqJDtxAhUPdadJMD4UfLX8b4OmnX4S
xh8dCXzpXYhqk72huoRIPiO8FluvKbsZIdjf7btL8ytygtwAhFE3q9UdnEO+SL0k
Vf0BAssS/Rve9mcNsZopUYf7VjZoNopWk5NuqtOAqx1brFOVDVnxK3CYg3vz1mOP
j7sKgwEQr3DUsy8L17u5OQz9mJnVxRXfFrP4ZO+uk/O2Pgtq31JrQC1mOyrzXo+A
2084VkpeGQqu8Hrrtp+jwrTIPdUmaW39OYQ6B9CEqQar7/cnbfleWtFKv1E9yAdZ
4Wc6ZtZ3UyObdRzZKa+MY+SA8m+XH7u87dLakUzlR/sj9ChB4KxCegOvhw0q56sm
QPdCNJG1aQ2OvTWL5GxJVSN0+qh2N9CqaJb9Tq8jTvwGh7/pYv1FMQNJL13SCCI1
oYfKAjA8UOanNzQqxakfQHh8huLA6uf42e+9LJcH/a3bUC91a0LeQ2D0dHgd3mpD
UEndcpuSUVl4OhlUL+Ysa915DGvc09j3Wv3EqJFyJiWXKAaqm8i5YS3Cp02cCq10
AZdg6D7x7N4fJgC0PCeqrhlUed8T0E/UfWZwnQ5+l5eSifub3Ll8+focmCpzuagg
E9Z3g0MYm/sKrILnbIMQjq3loMDNqb0iwGDwTbrqiQrsi3oUKDC2LoXVlEFAZkbC
TL4bp8hS1F2QHXULYx+I9V/I0uCyV/wTySL3hwT6w6wVfeQKdRkoAEUTYjzdCYdJ
/Ge0HmrekHSoe4eFQ5TpO4pvd0yXsbWki3AXMgRNigUeZPF2o9DKhMV6icw9v4aW
czIuWNDhSrWwBeuuJwMB01nmLVSZVt3GWY/iWoicmDryn97UW9OGo5nsQS6uUDGT
dX4kvX37AwrZFaaAKhSlMpCnNGZZVaEGIi6Byhodu67OZ2/9Mf74/KL1JvdlhDfx
j4b9Ajkq8+P4oJPt1S8yffl2szzlMLZc+L1H4i2+ceVxvtf6BVAM5TELxXD1o86r
a2desUcJiX4AEHew2ZUa9jfteucy1N78N73JUMLcnlWXFGyt+hrHgRDoCO5VTaNV
GGSF7lc4Qz3jf6pbj753BRfNbaXpAhIeJTcZXvowKzzgTcd8DzauZRcar+G2dLGW
kDuwI0UikKoOL6ZvWQ8nwSE2jcuhBfQHJzt2KbFOlU4TPHwLwd35jmWRxNN02/fI
nrhADwwPe251guRryqGOn3P8c6W5k5L8pkH+OPI2OYnJBygCGdJrNAEO1/0sblF3
KJEBRBJGWaiHpY8+oqUuryhZrUF4Mki5+6+CLblPZftMv3nmNsyLgG2CBA6OLjrz
mxtVZKGzlOn4TC9pbKc6Vd1/8rz+urajUNQqXACHxPaweI3vJl259eggG6Fcfkcd
8JvJfLNxYDaWmaIRfbLX2XYj7//7PIrNT0MQDHguDO9xHkIkkJtPpr+/GrRjTjrQ
ZFV7csu+hwuh+I5F6gsvTswSI5+1zZyVuQy0w2O59zO7smipUrgcRZcTNXvaHZpX
cUnVHv5z0yCbHpqmD0aLg6yTkylkXJdaiSTpkNkSAeFq7LxZ1Y+29dKnRmicTI3f
7/s9Gk6w8wlwJPSgVD13EALMLpcUyZi6YfjEYIVUmQmk7Jc5lqlGX5EVIxTUyLPG
CQyADjvL7bE4f3/UJAiblBIqGiYS0uefe6anoyOloLOWse3UyTUFyXNNWwy4gp1t
PZ0RSyd1iTfx3kGbTzwmJcq0ly8x1xqMA2Y5foLH4xxk4zopyaAl9zsV2f7N0aaF
Z6Tcm3EcTStPzLHBVbRO8vSEdLIoUoklffTryOr6GMcNOa6iA4WshqcQXvU6alPD
4B71X1gd+RbLCFdkPt9DM6zor0I87+mm4cMoez6TZ51Wz/hTX6pbIYr0WYXVzYnz
Lb/vygmzuuoR72SGfA7tUsI+09nrLMvYB6yPuW6ZBARMWQ2/VfqvDfE3j7qHVGlw
ZzwNq9l++TiYdMtKKluHRdlmSIhFJ13ZCVA6UqRvcy0TPNcyhAQFYbN6nkWTiTfO
8A+UUQsVcoqdM7h9EabmIg13HYV7J613fk5tI00CVYo1pfH2a3DRwVGUmV+FhsI/
tH5aQn+bcWyqGRmTYP5eBIywaDRY2b4VypaWDkaF2hrHAcyooxoQH4TplDh8LTdI
AkTv0FV4rL777CQW8RV53Y2aHxBDaepoC93yA6Mls48doziu5Z6E7Wv1jw02PtX2
aZ6I6j40G21EJ78EmOPamyNyqzT+mJNsyO82XZOHNOu/ZnJRexvVqAwmsMFqn81G
RTxGSkBxXhvTNfABywpaE+2ldBM6DOMjLe9Wv50ZJpx1JRVFQldlFmvZ2Yka/RIn
rSMXO99H6AXNFEorY8weTzmIQvUy42dwYtMA3iBZz9/QImjoiYLI98mvjrD0/u4m
sSHLl+jPCJuYL/s9sWZ5KsMgVnOkRr2pAX8aUGJBB07CQUOojrymWQsTEg/ndS7G
3XoYZ41Y5CeI87CJXZbu2BeFy5dKSU+kgUCn4igjQJBrCfBF0ZWKZnQPrTR22TeF
4l5kPL4x3uiZLoOXPDpBNJYZE8Z05t7bAosuTGYh3hGLO7MsLWJMYSwGc5aPUVcn
BYu4n1SnPZ34B97klettaICtPugslyL7yPlxWxoQXBcqF193iIVKKdTccwqRbGgf
p1S56gypWfsY3NUy3C2e6Hn3A/d47OPfSE6crPtbOS0=
`protect END_PROTECTED
