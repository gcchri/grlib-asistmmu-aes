`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j1XS+GsLx+viKk26Z/tVn9xbrDIj4HlBSUsyhPZpUXPEfkfUakaRjAeiUNWYTvTh
yFHF3onrLhXmzrP6oKnGTS8YST2+pw+tfXJnTuYapCitYzWEJvlTgbkER6hAh0ta
VJsJVBWVhfi8NcPwOD/Tmhj5WjUMeqyYrNIV/Y0KgAklR5JqmcdzWwrRKxyjM6bL
Z5perNxlDJGJJjpRyc217BlHPAclCP/IW7zK6JE2FcWX/GTyLmKjqEVKOhVsDjPt
Wt7LLN4uTyfjXV8BKVd9sku4HCFssxNDxUAN8xOBnBI=
`protect END_PROTECTED
