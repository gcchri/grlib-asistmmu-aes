`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcgFQaZ4wB57QCJ+OhIKMp2f69VZEl4nF84lFm132JcRF95PvZ1UCjyZ8DNWvRmP
WRAFHe6SeQ1To0Oh5Q3cJx85WSJsWSw30SSVfWizmM96rGXF4uCI1x+5OaahXy5y
aj8SjFV/bHGeRStCwA1HWo+z9lRBmdyIEOIxoG0vHKOclqsFpkIflP2zs3bgk38U
LM+InNGpEr1K8e+KZh/w03aSs8oZAGmDwR+bJW/x6UHD2LWwl6eUMbaRV37QXYDG
zAlLF355Go6UV4IAjs8+WQ20MgOIoHeotTqUoGjTmGZFgHLfFDGj5ppJ4Bc1xmHR
gsko5gOlcfoNb5DbjU5wql5k3+nxqG5auWNbxIXPM9BWLZRxYuz4tq+Mm6PbJwMP
GWAxAXSgXPDKfBa7D9ZuwWW/aZdv8/cNohIzUL3vMZJoCieaw2LbbVOmnSbWt+yy
DUqYpSfQviG6LHto2UA0ePSQuN1Iu+Og7UX0nmoBd08gffRzmI3uccEj7foKIJLO
jRIPTofweNwPc/uyVnJSwf+vuS7AkQ8Kb9OMPZX6y896ob00s1GynvDtm2KnXB8G
+nb5E3vFCeSnlFKLLQT1KypMHsxkm6l2LcfPFejLVYtCd3AbKHvEoHsQcuQlFC2P
slErkDo9D2nM+2IwQCzX6EQ7UJdjut59iWwrc+VbhwxqhDvhB5qTKqe/FgQ2ki1Q
UTmbTfNZphvFkhOAASzzuTteWKdWJRhNIpWqztfuJpa+kLofPd84CLA9BocXp7sw
3Ikge6vjImNbPFITiNIQ7Q==
`protect END_PROTECTED
