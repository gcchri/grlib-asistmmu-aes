`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SXjVkEpPQzw9zWTa7ZTAup1PAOH59/W9QxpnYGY5XF8F/uyo/M3aBLgSLCqLApql
+zjCMQOEyhlNR3HgQznTuMYxpZeJjFBvQ0QbZ0c7B4PzAHd9P3gydijebb/ZbCPm
vToHfl9YZb+9//jLh/oBpccej3uPENRrP7mI1zs4Lo7rPOwm2qzJUsbQhv7KPumJ
hMPhpjM/9xHIPmzACAKLNyulxLBm4ZcKsmwI6/1nFqkjI8EpNEdiUYMV8ZsJ7BoI
PUspG0SeaGRAOeBNsJgDTQ==
`protect END_PROTECTED
