`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SlSpCeXm48W/C0LqMOFs5S8CzrVqKc4QnegQM2gcrHP3GYyrKge5zAb4ELYHYMKx
C8AVoy8nsOla8Y8of+mq1nlJY0F0FNx0579qprNbJvuai7amUnBZQ9avBeiWyKnh
wHQOwJ5uYFNvgTBJacf8n2yRd0941knzxKEIjB6nCLLsKRyYsTAOLw+wr+9B/iE3
wV3VeWWIolEepyzHBPP3WONO9ddHK0QI4q7YQXk8EFdQW/y9tJ/TtiAXm2rqSG8O
KcEHjffoM8VR8dn2Eo3VXvDnIO+SB7znX3gRLE2lVIcntnHXgriVRIhUEe8zLteV
YSXk+nC5ABsz5XizQcGCyM82pIgnUfF50yOuDH5LG/RtFqGB7mmZrid+PzRFiAIu
dg9kYWQD7X+OxJ+WCZN4vkQgL38E404En8ltIGl+b2rnCasqk3KA97xbZwU8zcgl
M8wB5SQhDX4dAorKb/KlRDUJdYvYW8Yq8vyj+mnGkOuZVz6JQzfZWq9nIQ02QDcz
X2YdrJ7rrFJAVpC6BxWeiJ7WcKdWNcqLbTowgfoy3b7C9SFP+kclmCczR45nYsFq
k0YjWxw+V3Iup8q1Cfjg2tdse9u0I1PhH1C9CPssm+92i7aTj6Ee+mFIQHDNPjCL
OQ/mHm9aLH6bwujUYxz+kIAA2ouslQirpRYj8B/RIYCYjs2jvob5vllU+TaQFgzE
f3xtLrd5IxXLk4FS4m86T6x1IdaYZULXhIms4nVy51T60t236uuKTOSysCcEX1xb
/jwH18d9j8UHvAk69PG6kpaoRtInVDE9pc+29G4vMRkIgq0/24DfBxHiMclqaJ5x
wc57eFJz/zj/im3AKaz9p1+nGxsXG1WuUpICDqI3OKXJ7jm5asjcGmNzAND791t4
wkJb0zZZfmjrgI//ALWz7l4/yYu2glh4i+dYH9K3XkxE+LE50VBbMZ6aUXLw51Zy
e/XbxD9Vw0wV2cl/q9Y19fF2iEhUK237gKFqJV5dB3+Wp8k27OnJCeH/4+YO3z//
GQfWkmSXjEAjSTdJPDTbaR54c92TdbesuBCK7YKiXZj3DHi3lBkL+RT93uZIsRyR
LDTPDNBTc+14vmSRGkkkTfFIVLlz9x7rG6hQKeGZQXI0cRyMJHwmQInOlOZ1Wabm
YftkA7v3sxUb9AL876idJA==
`protect END_PROTECTED
