`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hq7NEopb12qsnn3nGOqdnrLrzZfktQzQUbjqrv10cwO8zt8dfZ3CxZ3Z47KlQDoo
xXwd6M+Ci69Mppbp0QSq2hZgFFOLS4yCjq5eSnRioQr2zFWfifICXbVPVPMuaLwz
zNS6/ousIO7wDsI2pcWsmTPESDlmS0rst/UAK61279L3B08oedkFKYlk1PeUSb6L
KmsD/qDlackVSuA40+2c3nxEXCxoiO8+wekaaZYWnlEk2WGYARCqnwdNReFgLHsi
QHxUtZXPdu+vrn6utnKLMKp/ao2JqAJsv283q/uTTo471SgxGberQJswKP+7RiAF
UfI19frF+050WSstNtlrFqPZykqB/1rKe1+OEL1JPrDCwhdc3VAvooCXoV1DozgS
28cJ4jafqvr1yuuH2oKkPDTqXyhCM1guFsZWrBdXydLSq97Ky4n3yxqd4KXM1Crw
GVjikEgNMeWlx2lktTCkHU24sIUh47wv1Pg3igk+615FqSxRh4B/AqwrkxC76Sec
Y+ebwBva0FewSTHl1qzH4U+BUazrWpcQSHkhjuYcDDOA4+3vxqaecV4sBhYKX5DN
yjWWkCr7HvP3iCYK9QhI7VOMybSxO9vTcAWItcVb6DPbl9G6dsyAvmBXTaaV6pMv
RWqTfFDbuwJPdJl+QZY3inck6ixGKzgUWhXckHJcjfCTqKhB7QRxV8adgqVPjW3u
VezgCONoRB+fmxGicvWqDVw+xVZCb8Tcx5PCbuJD8D572EpgrnJmk+eV2KVOtweW
jNSlSOnC4x/hRxoD1Zf507+ZhCbq/uzM0swaxnAAWmYFBN4S6zTEgbDMEAIo2/0M
JOL9pBeqaM1fgLrZk7mplwE3WOFmBFogm7w7KbrWQPaaJk9IXASb+zr7vNDGFT9U
oe2o6mxgE6D71UHX2agL4jmV4Oxu4lmbW095T3yBzMu0GpTvfPzbSyzOtWQQ37Be
RPaMzcgLHPC4P7ZtE9ugES+TOx1zYfYztTOh/Wf1g9wuMEkGr1P/PLMyfAvfAevg
Ujc7JCBwvzoELsLklw9hT6evsDZyLZGwOwBSf6TnAiDH3Y1QHrDZDPnQ/K5MfiIU
zTBzgZQoMXUqzSGnQ/MIJD7knhfP+w5ZQB974QRKDH2Zl/FTRk6A5SUQciA3gQk+
7s1OefqBvaf8b88EfDTnX/n7QkDGN+a/BCkYaU6GLW6HdjfnQcxLWVgcsDxtaBX9
/OsBTZMm7xmhycQUbRx4Bk6yOgBe7KKqHrrl1p427mgSUON+OQiG6TPj7pV+gbwn
YSkpX6zllj9vWT10Tix8r6EzUK899MzuF7bG3FTD3u7KlEIvmfB7cJr5UO3KP7VN
XE33LSnP6JLGtn3wkUnui7zswRAMbaUwl0NMRS4b2mnaHrQXFTHaIt6l6VAMrVFU
vDc7w7XuPvlefi/LETwX3eM9ypYo0SejeOcQiqjsxG7R4+yRZ4rpesDtJBr8m82U
LCrPwE2V2gl6nf5IjOYU6Le8TRSDJ+sl7DUDYexaTOnwxB/2cMSu7eBHYBp1DkNA
HmpyJHd7lohTmO04yPsoLFDYt+Lj+7TpHh3e9xpypRoGzQzdHnctfdxI8Brswve8
iMS3d6+2Qkxs9IEn3/wiZnnMYrH/ZwIzooI+cZLZTHnGRlESUCPvFkgvYPkRB3e5
dwde5rEHa+pVUd3lzlcjuwSAeIaCrgmDWfWnkXSuTY9tTzKGfHxqGxBzTXb08/YB
3mp2rsL6x7cAFIbjMe0WB4TemFTQSyyc8i8JvLPKdEItDIs2YXBjDuJtOnzchPTp
wNUfO84Ga0P+Qk2JUqcdD06n64++3qVsM5Dpyw4oH0IdbfxD/TXnnnb16S3h1PTv
u8CmJvp+kQ1McKP62wW17/jWcHDfpNRdflIv4TR/pTD4PWzIw6srruuVmGfk1XQn
omlZ+o/tJ6wJYrLLZOSSWxsOKQkDrQ1kZy4oTYY+G70hiZe3PXq6sINwTk/5gAFy
WxyQ7pRt/8WEsROf9qRgSGfWBcBUDRZsLkz+TroRCdKk4GDnCUDU5nzRGpdxTuAn
eZOGVGEsC5Ptl4reEzJRZ+eoS5aa0BzHFOzM2OE7pPWAH3J/iappVlR5giVLv08S
LQg3ldmnGowmOtJVTdteS8kanYWN1Al7x06DPvPqETFVAt0APsaZVakQG7nhbcta
kHISrTaiV4tfDu18tL1BZaJCQlDz33dK4gWWaSbSGep8lXdQXahO9G39ahT+iTg7
T6dczIFlUhgB43IWVv4bfwOffKcAU7UzRETC3aA7ATl0XVKH4uZOZD+ay7Qm09UI
8RXaPQBMhNpxjPq/NjwXmxbW5L2DpQwBb6tQueKeNThVYo5X9Ct/5mOjmDii6v1G
ezPUlVR2D4LCz0ua61I9VkoyUWaPyt9cFMihbCuSUagOem1XvurxefWQWdab8WQJ
PfFbh++JoLlzktGum5ghHrqpUuNfUo3vYu2+bnwpdzTwNaErRVMwLvqu9gpT51BM
17dAjwADDoOG7NZYC7BtjeK8jnMyWoUyiyogJl0i9WnshV8+ZzfvMAkjwIOQbpGm
zMn1RwqoBqakXGn62+UbFFa+AzDSKn6nAR4Nm/yGKfvymzBmvkKSCZKBPCsZIsbk
fa70ll2sagT8WGQrRJMFTd8JNPssSTiYpxysL26eHMYs7KNIKrhmC4XfPbhFB+CV
6X6W3UUXHGvU/0lHkuR+mWFxwa0zuRp6VBzEJn2AJt0jc3bI5uudW7Ey3Sgf44Vy
vwC5KiGDZ+94Cc2Ij4VHSVW+pMgpafJhs/Qw38+FTRiLPXOv/Cq990zYH3a3uKKK
h6TkPXsQ/ln7yqjMEpbjws9QmocCTP5PDl6gForkzSb1qgYzVOkKojsPaxp/43jT
YmOgLn2OGGZFlJYe3lImqUImMVjU6s0N0XZYeeqYpp7A6ap/ZXRvu0dSxcpyU0dr
25U2hLJjW9XcsN8dmwgH3R43tipMstVW0iZ9bIDyst7uc+rtUu+a4IjX4D9T7EsS
jT2ip51EOwxPgBdRIE7uZnYXH6OVBbA55LhxMEAqUZhCblzMe9/ufeOjdW6NLL/B
7/HLeOoD8YFe/VC9wRBE8D6ab5dAAy444XJiLjGXa7XerdWPT2x0vuRLXaQ1b7Pn
i13gj+i7O72/1qU/SCZuA+rVny5cYQiU1wN/DfO1YpY4t96y237Zlb9ywOmWVJUj
/PSywiZ+yB3pX2QWtckFfxfOrZCz3rGgJhqL0+bLyo8/RLyKzEAI/LlqwpQa6AeR
C4jejIMhppm0dTQ3ajFX5VcyOxVWF8Bjzp++APPcDg6bV6/uF7WNrX55kiIuGqcB
XRO7yrXVmnTAyI+heRoJ0gU1/Bq7wH6ZgN7Q/o++i23xO3JwNQ451CocsICmEOFE
5ONdU55j9GVlWR90y77cqBq3wgmgtowWIziH4iYsX0dYCTpBD4AP+Ha0r03+4Am/
9y9ERD2eHv6/Ly3vyTW7SINCGsemSWTLsuAAiFZOdtZXEubfR6WI8Npi/fxoApVy
7zgD63edtmZjDnOWkiHtV5fUEsVm05HwOFbyROuCV9IywixWj93+tkxtnmGimmiY
LoIftMNRw78N42ooRroVJDk97HvJmkySLpadTXsLo6+H3tHurztyIhG0WEV1vIiH
GlmXyTI3qdYAINtuFcBzSQJlUZPrfj6gssYGOwkLrHZ5hl/1PkJC8xHjjLunbajw
C5QagWizdAQjMks/8UNiIfnWREJx+dmCpgxJfPKhL/xEjr5vERcIreNvx20jq3dz
wER6hp76fqareMCegBdMHtHIuVfuDZNTcGVt9wEtWMbL6HfInGhiRJoAO08WOkER
YuWR5qsQil7o/6Lv1mKJHgs7woRxenQ/GbybSGFf5q3IcGQYAngVttj9sjZ2rpv0
2NFGnzEhHAbuygT5Y1o+f+QZYen2Rcdv3HqrgpXr3YHnxgEqpF8VGoJt0Uhqau1+
bOBeaRQhsRNB9kS83UDMvEmUw9ex4kaLBhJlCHWISBCmPEkjYEkdjCroSFsGSK/F
siQDsDG0VOVhvhUnq6BYTyM85S8xi+SRsHSPSTpd8A5gM0D0U+ALSg7UpV8jFPqA
S4+exYlYbkCspw4yAB3iWMivmagCrGJfwrn4hZNFIzEqUho7uC7FKnvZ4GWZgqz7
Xhj56rscVSMDZe9inZj0UTY3gFgNQt2kXFs3+p5KfD1V9EGszVO6kVN9Kb0Kz5tG
K/EJr5m47ujvNTvVOjopUMSlf6VbRb/tOXTLDpa4XXERXBOe6dW9/U5B3GbJwIg1
84ttXa1FKUCazdsti+cQYprtjh3snZmCujgvWMLUa5V2f38Vwb9MlO4xa1E1O2MR
H42JYEaewRU4W4n5w5LSnCk5OAcDvZFQOmI8iEsDDC2f6FGvea2tG1UkJrtjgqbO
qMc7j0AED3kb3FhmUJxCbn2ksgRW2T0X+e8k5fz/M7X8lU9NTmeqT9S355IsyQCV
ZgGTQLhtdXLs9F1oF4CTkyWPltQ2qD8aiDHEM3Uz1s2FkjY12k3Szsm2gI/gtuKD
3WAc2Pc0vaYmBtjA5HKAar05WdBzeudzDIxkE/NN9YE0K/9tby3jSuR4rnYGfxzH
GFYwVPwyC8No0iNDc7rcQ8lt9t0dP9GInFj0ZREUk1EUjd3BNTcBj3hindUOZ/CR
fAR3g2ikLaan2dMX02Yx39jIL6U/1RAGGK0WGIt7wKdWgGRzuXKCQDycyp3AMGQ+
rKexvOziMJcJm4lBp0knOF+WHKMAdQK1zAz9PCj1q2RJ0VT47HfZlmR4wLs1hp2F
ttKK0AsbWjxsI5MlllDqdTIcbk2stF12cuPvh8tMg0hnLygmeF2DDWk7vl4bDRmb
49NK8RICCeJSlEhO1wY5cwXywYmUj9H1bbp0x7mnzAGR3ZsSIbWXzFM+Dsy6z13i
QPW0UiM4/pPHnXYGlESec2tOSEFXpqdf7/zB3rUJyQ6sFmFKI+zTiyP1CWPFg61Z
bn3U5yHYQFGD5mMviOOE7lFUvwnrn4PbFaw/DHQvR17plY/8378nciwPZaY8UOZn
0hEr0jga7eVMOYsPWzm+LlAzGkZwGp7nPWA5ucICYjyVzeUsV+yeXfis+L6JYkfD
WtoQbd/rbdoFMfxlamEz3vCFelWIsMJ9uMVftXCuujGWwdWTjJiSwl6pKNalWbb4
AMi/WmVr8v+7LpWam2VwvijTDX+F7pbO7I6Te7/7B5P0QsmlBDXV4RxxInJaWb7J
0T0hS/yEcTwfbDLTqe9jK+WIJDI9Kq+7fm1HrOjxCuXED9JAw4t1q+/QTDXJgwhl
lgQcrMN/dBw8jhyeIg0KjGxnxbEw8Oh2NOqYwgbUfAwypn9BruieB6AGnCc1wXzG
qDaX85NIfaO1AGmrUQhbQzOfShJqJxMjOjUD2lmJcxuEcX3TSyhU9ZBEpOB7s+S+
zGEuD/NCx43xU8Vq+5BoAK/KEoLDUNennFNGr0/Vwg6td96+o+njgBPwbJBKj3nK
hQLe5rQM5V8y6EIjnyVlv/JHsrVsTWaMze8zgSb6I7sUShWT+7DFyO9spPOMgQEE
vXERe66CoWj8gnk2HLuhyqO4G/iK978ACJaUuGMKl+5a3bmpSGXb9zlvBj0iw+gt
s5t2XlfRfJ6aIfqlk2WpE0tJoNm+WQjkVxfftbH863t+HcZvGwYButaVh5zgWtol
LH52wd3+7tRQ0akpDXGzRAiPSKdhJI3oKqfryLJEa0MdXk+PhYbASDZRuMYRZxdL
AKDslWimgTs7MXHEsjeEJS5Qyn04bNryy0p1yZdE+2NHAWQH2Ne1G5QMC2dIF4ua
JKlRe3s5QVZXCgVvr4XJ31zZBERc52DkaMf5Wqio+e3C+qhlX48CY0r3RwIgR7f5
njKhTT5FVxs82jTaX5ie31nEb3S09XMQZtFL2tREOWwtqpcpzPc/93ZWCfEQsifI
Uo/IZMus3sx5C6QCwoeV4fd8BKF1dkBPo65nsxOE0yW5oTxFNtxuOXdkqQ0Kub8m
gEVFdPe8Qgr2pIXfmw/iCsyhAxt7eijKIkZw2J65/naky7rFCAjzf8U18kEvLtr3
xmdeZR0L20wVU9WucWWmoZRJ0TWu63BhHZGmRsFz99Kl9U17FNgJ2Cz6QGttBTNn
U1lGikIlyBVw0ewZL4QJbDH5Dle5v7CRSuU6MEH0Q9RW7Ld3sGz2HZxlWV20ytAg
GxU5kQEfnmqv8W1K/1z7zQZpSq15EICoQr/PhwQ2IccgF/829EXAQeQu7qxVTU7A
WtUtQucVJwDhdBiWbO23oGXkpMdtL7c21nsLMq+J4gMScfxlmj3F3fli9txn/SC5
eRAJ5zGlfmKX7BuRZ25je43c0XbIJkyHnrNjYWD50aY+p5KWXiEWpfdHbxuFFzN4
yZ9UJb40z9/I5T7CgLSN2pwE+s7CNN78/BSP7w2uv3UWjRhzeTxAccU+3wqvVtic
KVaHiKQTwKIRWgLyUBdGbRTyRau9as4PtMYvLcID1Y5unW8paHXW0hqnbtakuopx
6n27a7WFXZvAZ//jNG3MhafyzjCSYk8SULy3Ia3kZ2p17cCiHxW+GR23LqzqWY+8
qj1IGpXLY2+jiigOE8g/G3TWVrhJRejT4A5oBavAYNFFqSSGAJg/tXqxQUfns1Nb
Le4NaWKAXDa23t7v/htOkf7QD43TXUgq+dkeVVsEsWRtcTNKspGdtnmiKiOigdnT
KAKLMZf7nG6wDLPpgu735mVDCBM1YZIf9fQQ+fIszF2PM0n2ZV9U1Q5zVoYFYczz
C6THbzQJQpBiZwxJyOYyfedud4qT2WOL5vhW/EafncZHrDf1rmL7bWL0HchG09Ee
C7Wx2ci10H8SMbwBCcd3Ee2rBQ9Jdv3TuEqRyIbf5eBlaAT4rNe/spWg3/r/GDmF
DR0KTDsaS80ly/xXUg+Zh2ZcVwn8X+qs+7GCeV40nBO7loNEt61v7+cCt55qCn7E
nr+F6V0kWLLxH6Mf/vG6bTMYoOiQY+QBTVKybQboaWyUoeOev5PAlqclLAix4iav
0xCI2Y6eSGhqHJ2Zl8AIM7yJSP8whEJNfzFU+Cf7MKhXb3rDq8uIi9HelsT/g+IH
nkIzcpBFDFzGmPOeTGK1ran+kgcb6CR+18qYcTnQkowOBLXGFN1vMkxs3FeZbXOZ
JLaxKdYsijLySvo2EOKtazIqqHiz/i48qJRtA45VcT0qS/S7sF3lpGNi8XYHQWKF
YEjvWo4XPVrtsvtnKPMj92Q1mrX5q0wtTDeSAxedPP/eTH8RCLyjuj9AQpr8MwXM
nxUaSa6Fw07vAHdpuxt1jURneAa53K02H5DH0u79Y4FM6eWnP3i+KnhvFiZKpcrc
m3Y+hGESNgx4Z8nAKUONwfsjVrMIT2ZyzhpGEmq1WPo4unRVb0MfD1l8Uj9LY0qF
WcKvL4VXSNAzXn1LkGlJGFgH2wGZRVobvnDtglq0NuFrPyhU9QplZYZ45tSfycO1
4kCL2oMaf/wAKcTLekTu14OEla9nigmp/MBlKawfNvTd8FqjwVPe7++IHgBYitoB
e+OlLqFdkMt+AMYw0vMo7dh01Q0CaG8Za2NwE8PMD2yG4yZQPQagtzHBbdsiZp3q
GCCGItYzeNg49rQQs1v8UquoUuN2ZtSm9RWLPzlo+OPq6PsUNXrkAx4rgNnr/yIK
LyauKT2xTCLDtzBmHolpQSaIHBttAcjmYkUrUDnTCdO1ITTf04YJeKrTCHIUhYxK
on+FUSqSagwwudp1CS5wV/4wR81vBg6Dk5SJOl04K4uiXt0PT6qAxNdbRUGUHbyn
+CFEkKCxJaqHfEyhDpvS+W8cxD/48MK8fay0V/RyFIL9y8ZIiVqnIKliFGb3y0Lb
nOTaSB5uTGMcQcRAjEEENLKgvPWqOOeV0aGOFa4a7JB4o0rbg4PDbBmdAk5XpMlw
cgGbfDQdj+wyhsCAGyRsHOEsdVUd/V4QomtbodziztM64FMTDLR7osddHkZn8xwX
MbSmuaFQU+LPyIbusKg0ZUkKBuDpkkV5yJ9YabqDXiqXr0lLCByJrR29haC4Jmv1
96mrAyeSsSoQcoPkHgB9Zxp7KShlE3CMrzxA7RGYiA/5VQGNtuUBxBo8sivUIG4e
ufItCeLlW3Dw+v1ZANTsL+lncaj5t1WQiEMuGd2dYNiplhLROXvweo97863ROJr3
ldKBTyXsxJJ/7C98mKQ4n6/fo9aryIU6LG7A93IKY5IgOOYNKsrTLPO/GRQkHoKd
E+K8JE6znGM92Zh0ySDqHrSAI72AOwZD3WfxLfS3BS1ITp3+3nwGt7ibGde6Rz+f
OyTOjdWC90683bja6G2K0wpiS23yX/phUJYYTzY8USP0oeHZtcPhCC8mvBItiSC0
SDbVx+rryvkiJpvdrWQ4UfGxOOVH0F3Q9bsUsUN/nv2t/pue/8nMGwHUp+LG8AY8
SuhiY0XEmHePHFPrC2lLyKxHb8fmrPfRME31ru2YcytAg3Od6Fo0HBBDaSkZ1Maf
b62aLmlKl5Qs2lUMshaVPNraFFOIZ99qOD1bN8mG8OzbPWPOaVXhR/Lif2QVips7
6J0d2BONPO0/wWMObbh/9Ho5Uve0YW3ZN8RVAwTBuQ7ruq+NP00LoWlkAUMSSMcv
2fUGUjgEEBAloa/E5R2wazcYwrKheu7AMnpXgtwwVSx/nUKBWJflYcjRcoUkVq4Z
FcuPBGU17kOvQ/BCirKTNZgCULya3ZgwoOP7SLJM3l1nBq+cXycz1sCUxxpDYFrm
YtDL3tu3Jn0sXq+SpPpjrrYoVr4kkDHI6n/LX4U6xuONLifdGuh2nxx/YaoBys1L
6itIdLD02TrGuKJZ4QK0IdPezUX1OM+lLfJ01Gnna70YSI4HV4Q3Yz6yjCOLshWt
5OJkA9j62tgcbfrozUUoZKLdrm2VyofrFh4FfY3BUwimjZrM3CXdAFMl5wvr7LYq
7bKhmP3Fh2W98A3APcE1d7d0xcSV30NofD2otOyZdJ/rvOZTR57I8eyuMmGz6Vle
RRyv0mvoMLJYUd7IdnuMcvVZ9v64uC+PTjs1rgA3ofskJGDnxGRij8l+RY8TUqSZ
FmLltdKhxNzR6adXAVs53WqOqN0gWPUyIxic5S6YrFNaSzR2GmEjtXXblgtQG9xS
GL/7j7FegU8C1XPeVwByZEieC56GvgOiUBoRAi0QDQOYuNzqhcKLcSyGwb1fbjED
7VB/HZf8p4iV9abG/Yax8ZhSSad+IGLoA/al6Ujdc+d90xi9WVTMJHwfIxiy7EpM
Lb437B5UAQG8Vf/K2KPv30Qb3d2W4urbuO/6FTCy3wbjZwmsgRyyuQnjIOBCjLXB
250LLWFp7kpqHEsq7/sf8WfBQECK2EHUa1fXC/IIBXH8rZrBEptCpqBKxh3TC3Og
O3v0OzcrjbJtkyP2BVZXGUoKtHP7fHb00n5T15UPawsPtji80ge9sqfU1NMa2QjR
x9cOC+oqGZK/EKohiCg+qQ1fgr0/fZw35mgHfpTH4pLOxsSHJ3fa69yLFWOARnmm
Q3enomeDdJ6uRh/FgDr1DClQJ12oCXQLdxPK5sqssDQ+8WmN9R8aWTjjMnsCpflp
vfhj2TB+7x6CvzmAv5/7anqwC5N4APAe9YFjOQgLHEBUg61JXKuR9DmzXefWxBFZ
07LwTOJwG+lD80nEa49wzIVdXJ6aC3UgQbV7LrcFlcEA4vQsPaV6X7mR6zYgFPEH
l15YnEW4XnFsSjCd0q2Sj1RjNuDbw7SV9HnFcL0DAgIN3S/gwsabrM5uSskieW+6
/opBo+Np9aYkbU/DTIJkqbbc0bZ1ri9U423MeHpF2j1HKGYJGtsXKqgO/MPSNmyy
4KkSCVJcBXlQt9lo1KLtIEUQPP2EcX35VZxKBefWY2Wtr5TGLZgb4wAli+H+vuCe
D9f8DiPrpBuACVsiFtG1OdECkm9FzKfmIBIkEdZAm8x4DZEetle027tCH4qDOrFM
HeXdppLn6s1g2YcRlZ/7P0rf4SXRdx6KyIeGjSlNP3hcOjR1mRvOukexEpuWNKGi
WD3XAfopKsSNB4OHid99anv6ptOEzWZVXZakh3bU0DlIsYprnuMbojH3Z/M9xVf0
qNdseCGgipjn2jRaeJrwRmsVCLKhm8UIwaxBTjdiuX+Fb8Gj6rKef6TQRA+1I92L
Z0ApmeZhgfKx/CHNGvVkG4+41jsuRBlTAifLfUVo3nhm12LVgNb1cm69eU3xmnlU
YGGUVbiZXR1kvQU38nSLzOGf0tCb678TEbFHxrKi5rQGpmB/p6XYpnCK03I7CR91
b94xJB9hqAYsvyUKzviVw9oH4iPxsNUNHA1HeOaxQoMfeeyDaf0gtR42O27ZYHjU
ZxCjLAjtzOqy1HXNdajAgqvWxFAnxe1meiMZbd2YGsHj4MTD1DGzRiTL6icfcdW3
1zrMfmiLLOYy/GqVuhzPQEWnsOwxQFcntEoRyEkemaxTfcrnlE1L87GC0HxwBZSe
GhS78/Jf06sJ/LZ4VhkbeTfQUEDCjumE4/jaBS01We8MRC0PsBAMJYH5dxQ16kEC
iq5hEY8/0vnbWHKZwovLPlgirI33H40lW4PXavXyzkgk1pKQD+CagNnZehhWO4D/
cFtvo6tlFoMFX4wEGKFWBcbUoWK6sTH/S9wy3VGl83OMt3nim4/1l75zY6IupChw
M7/1N4wO6Jz6wcwYy4VR1kOT0aAB21iNs+g5TUmapTD8pCwLi7FLjRiRr3VIWbbv
PqUqZR3N/dMH70HRmt0YpQvqUfR9MA3MEMKvrnUgF8KqOUBXe5GlHeyPJOgJc8aA
cy/f+l76+zwlWF5hrjJfaDAngsxfrNERJTuzTtRNf/tXlntXdOklRdTM2/yVDm0b
w8gmZDTVwnZyXPFikojeA1K3/8/v020zMCx4C8y/5hQCq3l9lnnfxSi1z9m/zETZ
HIEDnDw3fcf9ZIH1S3aN/bVBnzmu2fxpfWQHSicGxLf+qcVz6fXZj+BtNHKTlt6h
L+HznKVmvDH2MutOYZcKp9xBjaRuYZny/YsPKvRGtxUhAMSydzlxvCCRPARS2rFk
yPY/rSsi3XDWY39xCXQJuZGfjKS+RExCrDt92okIRBOVUnt32D+A93sEvNFrHsvG
2rAK3B1FBGGS5sJdJnHN0DM8743rgROWsXVm9he85qfFX3voGt/WIkrOQdVbD8F5
ZiqvLdaHcHQrW3JN27saZ8xsMal3I5YDejBKTJmH9kUmL7jsUoAZH4qpBA0Ll1+0
/yhyqBnGOY5GwLLhIwd4WRFH9mhK97lsSVU/j0VyDvnnRjEEmvb3cj1GdlCOjg07
veIAukOuWGAlcC1RbG8/SooVzisJJu/saO0O5ZuXFixkk8wpgzGYki9H52AQk86C
2nq63MpdPsh279Wax/MOXNP4blLGC39jDl2v4t14aNqXfcoRqMmfPz3X0QzV6HKy
baPfjHwLy8qMMBMTHUByxN9e8S4R8l7CgXeRePUQdeDE09lwQkqBvCoEuGpDqdGk
0ZzUNJ++BcA64GeRBOzxCOe6sMkAFXEmldH6IHMzUlb5QgxusX890bISCO/iKW4V
cM0IUocNKx+m7rxF8KHzad3GD1IgDBXNoGUNW6B4xTaevtrPs65tyo+pLROQhPxq
LYBQYMYlqdEzPGyWlepZWvqKCC7nzDesxgPtg/12fVuG26vZIEIB3qG/SLt9Bq78
dfAsuAfENzlAP1SRg+nTBC1DZQdtHGcfsxY1K+fogoNoDIFSVXOmG1mZNvOzkjJA
03ZhCpSbpPm4Y5G3iRD4LA646OpFuOQ3eWsfNKCuIQXmm3r0+LFZTKPOltr03xha
NUomdgCWJMvx2snj3gdfgTV/uscgO7v+pv5vCQ7G5OgbnO62SQLy+Zri1SvsuB0a
KIIxHxnN/NszAit3z4CaJmbAEqBDogRN0Ip/YyeP0p/CZo8SedBm3sanloJoL2ue
ZJNNEYYP5O356jOlDk4qsMy6QA7Te2LkRs4C++JaoVRH5iwW8AaLAs7+tuyhuHSN
yGyBneTDsdV0IBajL/qUFbfPt7x+1SCMwN+0ZuuE7PTQcau3zU4ULtEBlxeWblzh
A0rawLcqk4iVR3SFzxxacJnpg1OtZTB0aw4mrwtzDYK4+gsKXiYQKxm5FbgIU8WH
APBTNR62uiTrUMOqUrBvIm/qSnC/9Phn+vw+kfKiJUFU9xSDdRQE1qpyJUfWsGx7
KyE4cORn5gqGtnhQqVhTdHdWSzoJqiGv2HLtdxfg32ANtH0qTa9IU/xYJfZPJ+rc
0lcbpdkH+DisgMsWn/1ytljV2R2sMNMp775Ik+Kc1M1fbw95PVYjx+XZAxrjq8gJ
r9lXH2oSLSC612XRGkg7ZglnU3dJMK1Ax7n8+t4e1CznAAdjLnm4+CPaYZ0xgQF5
Tog+VyyOQG6SVwTQYfK1sw8x5F1XtxFrx26B5ZWJ7t0OG98WBNDsxXZn23mmEFs6
YArkE+KIusMscAVF2qC4Q817BJp6rz9k8VUm5AwkGyyuQSY2CVvG9iZJNZtlphN4
9841FULR7IgiFC5Wxp77+qiT7muLJv8gljx2uBNG7DeLyBqW355e+ILp3uD3px7+
fMhjZl2RY41FK2s9kvuWz/yqVcZCZWb6q+WOPHfUIItKvxkUjBoxu2uSNFriIJXy
StFehGhI13rJIeZp+ou3TeF5t9H4z222T7cvyv50vi7H18XHI+iQjPURadplmHIn
yIJBD/VwT5MQmiEgAhE5yZGoC+pqYXDqi/ZabAm2k+YusdU4z3xzv3ruEdPw9QOl
+/fGmN7tDfVpgvSUycvDg1qvaRwkxZJSxUQe2n/tgdlIUPEE3qmY7CZr3QAY8NQo
UhNelYmDTXf9OBw+5RU9E+SfhkrPbTO38i8BgVjafK9lR6SB3GXCvPCMY8YmLZYU
/D5PzplqpbTCn9SOXm254FpTyBMrwhT2dw8xklOHQE9V0XG4+sN/59RgETdcgdSI
+zx1CFqvvIxD1P4HKDogfQyPMmNW1PyhRWewGXVD5UwhayEyggFI+y3d1dfJO/xp
9TMCCQTmrI64+6qxNeBNDgkPU2ZrrzqfTj5iqgIr5i64rdwJx1WJtzwgXh7gXdrL
l6lftefxhxBG3GdX9ITp43jE3mtsItlrmpT+SSadPXEbYjcXnkagZokiBmhaBB9s
nI04X+y9cr4wRZSTOToOu0fVYsuuzVD8B1r546eOZPZJnNJWNO4PhybAHN9fnVix
YpYzzpdyRaaUZLTEZuMH1/dARQYeBI6qD7bGU54eYeROPmmLiwO1fGgveCN4IYQ8
M5kpxuMJyFrtUANzXxp9a91x/wXa6n0ESdLa7Z/KLJb913Sn4ByL0ixMRrSAr7d5
s2KfJcFe79BIkL5f0co5sMtWoIJEaUHAn1RsBNTnwuppDB0er2KJhol2nLe0a5p8
QbpCEicoSIjYNDsF3J2t4fcIGpV6siCHXVajoVYNql9RmZGpAjXRJDgEvd6hgq81
8VI2DCnpb7u0Zpn2lPLvCS2OAkpL+k1jHUHRony6MVudU5u/AnhObWV8ABt5NH87
5txOKovk1Eg8STEciP7/tSRR6vUToqsO2MN64igBMEWoi56/27D7RQqVqgB4FYT9
N7oE8IiEjOrNXAllU+vN1yKR98SYYLpTiyUpAuKIHRHDIffr+0BQXYsszzx8OpS+
8M87OLAJ+yH/O4DUST9h2n1l6d6OCDpyubYhYJP1oYoJUk7gdpoikd79+iq73sAB
BPxu2dJqr43Nn6N9PYUs/JJw/F/Kzs5u6oWMDZb1UR7LOEDPlYGUZw/oKjO70FK2
P7pnvQtmqokFKvAxJcBXXwt2/gVDm5171AUI7JTUz4I+QHfitnm+HrVfK+jx9+Cp
IKJn1KKorO3G6BYe8Bp2ZHKwYnLAicPmst0M8tNd2u927kGZkr1QoRWHUIZPnL9w
dVFEdrCjf/k7xtyu3XpVqvKP2mZXFoxxsZgx19tyS1M35GDlGVAKs9THW+SK4pJl
XArX8cn/ZUQEyujyWbQD4fq1Bf0w6Tn9MZFd0SCtwkIM2HzlMXix5546BODr/YR/
8VgbgqfkZH7sO01l4pG44O7Kd/cDRyOwFHTofrAlQ59KoSZ0PUZp4McM8+LG7fHC
9gRHGF5+/G2rREH7GitW3EADJuIWSXAqKzMbpe64zZfszTErKk+UGsAcndaEwURG
6Xi9MsYmT/8lMqToObpyjZ3MB6/MCmCFGlUSN18knT7Mwf/ZNRQH/AQ4f/APwW5y
0cUd5/mPYSGg7LF4G1CPArXgQDesJFYvKOy6PmfzGJd3aFXDoD6J054DHEBHkvcU
jHaDaDNC2YTLljOvGt0lFZdQ7fcZLRh8rfCFkbdWxGtPdDoFDGwSzpLygrw9dkF/
KFB826Z/XSk/gQ+aCuXJx+aaprbDxLwd6fk+9eHVTO1ouxv20z7bBT3dkCDotKCy
cH70haXCq2PV+FTmMe5Q/krzjYuZbzeY7HisyQ5Nj9KxboJf0xyxEZYev5M6TEiH
6YnL8+PFkaSQw78erhwDADkyR4+zOR+AIdziVwd/vIG2PW8iE1drId5q9cdJb0Ve
vd8ioo4v/cIPlbG/xKqjtwL8Q2drlysegHErh+rlqobQw9Fd+okCzf8UXIQusxWs
ZjIjcxnxsOI/y78D/fhxiiduuIz6Om5GqelMRHlse8hpTnvazTUrS/DEDIqWAEte
U3BCJuCfhZ494XDmR8L1N1C0Qx3doUEpqUhbIvcieqeRs3FHNxF4u+XWrl+wewqc
ROEyHbdqQS4EGoZfyGX5hSLnen+oVXgNWCWO2z+q2hvMwz0mrT8L1a2fV0qxWCVQ
BRCNK2t/fejFc7q/PHNgbip24LnRhDy12pwoLWWXTH/bDHW9k3IN24iht8gchVQR
dT/ppw7F7ap0gXxAP6uzSpL+zrB+6/eBbAdvYjWqJ7j3JM6N5DSYRiMMctgcaFqB
iIdzMQc2wrb0SS13xj/Xo//xK8u5gJI9onYvkxRpR+pwv0stQMlHHbok9vXf95pQ
E/VTk+MihVvAd+XRXqv4q/M7XeMDo0+iAoHP0cQyq560o/pEvmkrKorkZCNkSVSm
g5+Zb7P1+pbXsOc5uY2rcoDXI4fhl+iuPlHDx1pYQa3sqZZIvigjD0XnapUPvudh
Yw0NxQ2wSe7iMWVuBFQjtqfqT7ORy6BODqtPlr5QQ/CWEq8xKvnjOjJqfe50O1vC
JloQapsB/rjDTdV+KbYjmWOatlU6/cHX3puYupWFq5KPVWPzcfKhhMUBbC9dcQA2
1V2xiFJfoPAUzKAgSwbvxiNYbVEyE7XxpxDr6gxHHdIIEI2two3j2p87e2kMieTN
fEOY7ozQ1Ym89DJEOYMcLzUnJitJ/sWFMGlNVzopZ0iaNTZwWQLWb4qNZlFK6WpZ
sIbmu25ru/IriC7iTtG7fXyDuWSu5hLUqbwL/fXC7AtNVlx6NZ5Dd0ADR7fadwVG
A4c7gjXBTDxyhjWj9aZQrHvjotcaZPpqj4dwHURKl6IXm0stcvUptN06qWFrF+dP
WLGm46ILYfdRKjbfjjVZYTPIFpjEfpGT5XQvUKRcgNa+FB/R91StCG2IoXzv7et0
SLJ3EDnU6PMgbeSTbxHAwOn6V6i/frwCnKXwOzAiwOorPQlLDH7Ffmw+c9KbTZM8
tjzu5Nb6xmG9T5gVgaPw3FXS0/CuqU5ehGElpODloWKbgBRMcv7I71zmXghKWkEZ
SCMvfk7R0YQ1yWvfhDokyxfPzEU+k4+3MxyETNSEbVBi5wfM/S/WpZ3M9JuDfI7Z
DwzQPdvQTL6QwE0dkDFfzn1q4eb6o09c/cvNoTFcreIBeX2XC5TFtjVaUCRhqMGO
LKToea6eTldJiDo2p2Ar/b8fo3bMXvw8e3JfgmXEEA5uFzBbmy8S9pfCx3LxhLHk
DvP4h0Iu08RXjAMVGXg3B30HH6y5aUfNaoEFPS2RtVjT2PvOYU+O8llrjXgnk2qf
/mWvlUIpTVGQWmzadqR+Imc7kUMR3lvpKln/x3NsKfRkNbLvS9dowihJPO7JP+gz
NH7LOt9LOhdWR7ljUimUoBzJjnO35dIexZhKF3sEo2MWhhFb3Myr0tKLfPHtAWpw
rsJ1TLNplc1+n4VJPSf/ur2yYiVgoCpE8q7EnRgRAvbbvNQBfU2Pb59TxvGVOoMm
WQXgEmCucdUkNcf5kOQM6JvyDZJnfhrUok6YZAd5FgbVkwP6ORhinhyUyA0eRt0f
OV7OUP/n3xFbcmTptgm/HVK6kukKjOZcd3i5AJ5YjWmbhBF+e+X6xjIbLaWUNYKO
lgs1aS4TjyGzcEqlI5PbpGSZF/2OrSeT1Gdk+oxSQT+l5AXBZAwTKtKz2LiCFRYR
bRO3xDLeeg9xzqyQGo5qfudWZfyNrsQ/ocOKuRVkJYXdMXIbF4KBlGuTh60mpJnW
bDf8IoinWT7EGrm2T4CjdBltvCCUCjImshB7rcRQi0QXuS7dTk77+OUY14Hinvrs
3ohH6Idim/JEn4PP6QRb5mAs2JQmnaRCS7HJnhWQQoeMZefegQfmIqdWkRTdWytS
gLChx7hdnZ07OPMlpxOOLys1g7fZcSSjNdVZMIll8iXKWwGHwRzPbpYj1i5h/dqD
poNu83KPpTfZ6F3HjXe3Kn/Drlz0+OXSBa6RteALJ8XjbE40jCfHVHK9qDS//bTO
yJYYrW3+wZmBYf92gpLyyXVFyJKrfmGY6T3fPhiE8p+88QakVAdUW6qeKHkDOq79
glqgYE5Xvl6AmIhvrZVnxC0jpswc5Y7P2Gx/RHFfTfodufpjZydVl04Zr38cpU25
kwHaA0b3bGwH9MsTOtgOQ+gflW1ovJ9dHWn8FEkh5fi3PwodhWDvRkz5QCnMYcnx
J/jjkiUL071PuBH44ImaxNhQhetfakQtiqaLj6Xgf4bdB7/wI9RbGOaC/QlZH4eH
VFR9f7bTa3xm8pKGv0mWNqnMj+1godD1bJqGxo2fl2vHAEbucaBaxNaoXcpbxPVy
SFSqYld6xmsCMNnOweOwFZEMZgj62FzmC/J07hHRoX0RdOya0jduyLEvOasSQUR5
d1M7JVpB6ZHyB5deZl2Bxcse1tZhAWo6IztdCNchkfdSqC96h7KC9yutFBAv00F4
ngk5+QVLVCrq9CvpSeiiTPduYQEk9Zd9cwQTtb48j4CAjINA3oBBgD6eUndd8Dzs
ckLzXpOoFf2k+dyQhl9HQiXz4psgs94Ah2oImeZ6BbPOq3hQH35f2OFj+R7G5u6x
2eXUczInvcpPBPq8RANsWzUmA9WxUoF+XdVG9IswO7CnlOnO6naSHE5FNOHmDW7E
cQy/70CKY8nmIxRWsXIFzbsxPBiYL7DiLNwFgDjmS28LMawNgiwzxH880KNtIQ6R
/uxnZa3ovGoB+pm4+5p+xkEInVKRatg4lAFtTlcsHHnWlrLRJUt/t/zWrVycg/Uj
si+tRs8JHgvSaGTSCryhOahI1JLJQaQ7Z3vk3+h1bvnbrF95KUMOspMZ1C7oopEQ
E6V5FYlQ5MP5yVo5cpT48CmU8rTGh/PdbSW5SynC7kthKaVZjZ95qeuZVYKQrG2X
9QgqNixRwxgNOwH4J5zJmd30G+ruiePmAKGbP7Q1625sJjECOExo6JF46axVnDyD
OPJ8L0CUvMb2j3UT3ozyGE7lvkvDhYfP0qSYBJ0a94NbbuFxrAVD0bX6sdEEqe3R
x4eDRCXHQl+rG6z8sWoU3tFwUVdRUn8tcUHcYsNskvxc0GYzP5QJYPqF9fjS3E6G
nFm8TUty8WxGsKQtAcBikvwux23EBtiNYLUc8g34Prtmq+zFaEfJP5YAO/JVwpJB
CtHCT6Xz8yYtx9XQiVmF3kkbJ54Bon8t54K99MQ7RWPe62F6msKq/Wll7nxl7srb
G0Mc/3iAXCpf38TO2pQJQ4Py9B7xrjo8LWYFT3pg7YtwC9Cq9cDy4frHKnyLR/Qc
9sGlocYL/l+zJ3sG2qNZsP7AfA0udckCreTj0xX+zA3uArK1rjWOBk/EOXdLOr3E
cMG0eUPIwwFIdSD2z9+fBQUYN/dnhE0fLDEj1MiU8Z5I/67oJCDnj9yRqv1lor13
9WyK+lI8/ivv0M3Rr0FdEZ/GgILC9FCqXH6tpHLIifpAR7cuDTq/qRIKj9MOII8D
qhEiwDHsUbSjyk3Nalb76E1/SiBKc6axOFysW5Rcsk2a5KIhIwi8nDp8msrxX+Yh
NoyFowgLbO94LLGEF54L6lEqWrnN1X7RN3BiHW3r71c5QlJVsgBErBvb25gQF8wH
8QnESVMIrLvKa9j8rLURuGHseP0+jDBSSTa2ESmBsIt4XKdl5scIOK7LtRm//S5v
gnWISoIhJNPOSx+OYhfZtXpA70tc6MgiBIouoNJABJQITZg9RU1IoxOKRP3LwQxl
HdvrR1VA3HBjYk4MSy2YVoGVdVd/jEuaxj0gTmdSjDs7nD+cYEjgSpP48xqOXV/P
kjU7ho73x+cpN3W+41LYgJPpxnyQidu1ck7DnycjHKcVatDS2ehcCCjhjQypDBB3
ssQ02q8j3Q3yvOFiAALePUK5+pN7b70SCHDM+InJREk4qBKXPngRh+KHIGWV3DEY
GXhcgOEvLvmUeh/jRe1VzQSFY2Fa8PVDq4tJcWYw5/MuBiocJWNE982y2CAjj5Cn
B4m81a/JhoPwXZxTAfRDmerd76OfQqLpMHfIWMgfN/bbJg/XnIRoxj6DUNDr0i2p
rplEcp+ykTdGJgVMg22H83rYG9tJaOYV/UdV/k2asEEkoTmChUeXG61Y/yLdsgJ3
nlgvyRC03tXeKVKgpRR1+x68HwOh+nDbdSDH0ZuAoeSGF12ZwVdx/E4JOI+7ytkP
nmCgrycq0KFMdcXLEwwLGhI78HH1mjZ/s0gRNW/7fGuOWjF53qXbJsRmYs23vWGN
rV/nHSbyw+qS2cG+omIz8OK9sG3JJKgYcT97fkKkL66kiA38TNMG/FmL9A4e2GMg
enQN0zCwSAMWoNPhcyyuHIhyUGFNwoR1eScToMaKS6SzEfi+mDXM7/laN9un5AHY
3a/aE4IlpoLBoNcl3SRIwXyjBZWYanA9n7YmO6rLBOLJHTNi0Dp3fnW0TfO4Nsat
qkcAPZE/gN8oQqhcAOzTQul76zGuPw1rbMrHVPMwH9yUfxGkRtOE1WlAe1NMTpEu
EjBXy9aMDAlqLibg6AKabqH1cFy7Rw5nzXAiu3BOu5JQX7W57Z6ki0eP7IrI+U0T
1zUjsnMkLZHaajHfTzKgrxxXhjkzqs1w4M6bY4mGTzg4bhZbkxw9yA2TWJq7Ylq4
Rbt/IRSi9UVciHgVyv3KvktL64duCI6Nu23UDOrJ7pcfrOV9HJTy4CRKUw3hmcY+
Hmyo1tfZsjhW8WF0qna4KCKNtgyuAIWNWtwOYmWz9zh+LNhD6oG8Otksml/TUcEK
O1jQswMxFQ54C3CnVVXXWAMRcEvpZPjJ6JCSyxF5dYHwhtOo4M0PD30AuIX/f1kF
oFWNqZkWfX3LU0/aW1NFaAwKQhR9Q998OAYmWrhRhIhKZTi2WQK+E0Ko5y0jZGS7
47vD5bcmDV313bsj0E6lV+paG+uMmkj9qsv2TBxNaNaIZd60YNW4XUZe0AAAX5Ri
fMfO+99uZHmmvXo88ossmp0gBbGxee7we/BmNBeRdTicTWcCogFpaZGUbrTsE4Ul
+vahmfvAvXa/0IHCOZe8f8xSdyyQU7SOSfQ+SU3LAi2vWl4wlwEpvQ9ogp+jwzjE
cVQ4r+syevuvdKIO/m40sVaMhu49fgFlG3od6upyHssqYPSdE7EHNB9+ZY8Mnns2
kUfvDhuq2t2Yo4XccjrwnjfiVPUlYqfdoRj0u37+vNQ1dpTTZGVFIyjtDQKZwajr
JaOFetxEid6fs2UJVNxAsfp5pIvN045hGIOA3TN9Z/fO55kUUuaqe/JiOF07U0Qm
s5krKRlSU8wjDPekaJPC8hNzMm8ECkwN2nQzUfQKJ86Y/6AH6MrDAc8cA4Zd9q7h
4soG+oP9MqzykB3ju5eg+IcppU9ixi6+dMUV3/u3Kh4NssTcevb2ieRLEclHh/CD
+39kYzra4bzGtUiaTZazR1U0P9jlH1ussMKvVR0YfM+2bBPqvIXozLVlUEADGw5L
YPdawHIB42VkVgKahL9h7LTuz0ztq5nk6zI1KgDXe+jxLP1NlkwGRALO/8VdhFXk
u+1B7GtQzCjTehSiklJoi9E02/NRAE64SDMO++cP6MkWEcIVaqe9xZLlVRwpsz4q
NrYeuZoAymo8o3fm6hID8ZzG3Yim2fs3tSJeQ3u/MapQZ1OPcnmRrvZ4dkvBzUuL
MbmiFMPAn/7DAbOvF6lm/1HDgS+miXa95u6+ahe/hpvMyxuMmqVy7JVaUuSHXS0S
S71oi/19OUuq8LbmNdt9hAomTXiF7+td0UqavdV0IQxVwdH8/CHMEHf9bBfsrbxJ
y4/2NEN24hqLlvwjj0BIqWywPZDlQXE4HIQWLo/GXTS/hPN7Y0wDpPDnDQSapeWF
Ih7V53B71pt45vu55W+QRJ1ahAhcK+c6EevYaBViouyUErd2yq8E8+AaP6PbRBlO
QI1G50Jjf7cH3t4bFc0BeHOM6Iw3KbIRSix4IR25t6z8bF3Fz7eg+YLpLMjTLH0g
6bOMpwgaVnkHz47Ki9qLfVh1gbLF5IchfjNNVea9eo43eUgJZk8li9VpypaE/2NB
qwbQk6kqcxnH89Jnc9s43NTgDGtCc7pjs56iY1x8O5snPeh4al5WSop9R0yUUbdw
CTlsKygNTqk+y338OZ0EkIKnvaA8KcrRx0ZRlAMjiGrZTbmJNJMsXkzs4rZYGr7z
eCcPeyfgYdzSfipx/qtG37F6AUfsjXJ0zuWysS0jQtpQPKKam2HdMXJnGFhh4iK7
7fzcJ+3AL/91brjY/XBOE7B0W8Bdw54/sjm9RXzAjiOYQ6tH5FnzLMb1Sp6cxodZ
u7/OtYJj0zJfySOEmFJO/TpBrmoPrzO5DDF7wYfMfS26gzYsoIsFHyifvLMbNoR/
Qmq0HuE2uFza6nqsjsWNrgLxDV6CV4+6OIVh4tk2iHNxigL/AqetB1W4vGuSnH/+
3kdNwnXyL/p4FHU6OSNtlV16dtW/OC8ZO1ABdNCaAU3TVHGBm/KoQPYg7ZlRyDMB
ADrRy191jDCbHhTUqNhsMfjxOL+Cxqb5MNaT5RerUhIPMNQBoeEQaA7z5rx3MMtR
In+hDdF0YZETUEnwJQTj72GDt8eVii4IEQipRqtFocCIC03kqUtwqbuyiUWY+bbN
xY0LUylA/Ap3CcMBGWgQz1QQNu1/qmdMuOT9a1suHqoJxCY82w4ctKSaNqvp6PMu
vZGCpUNk9tRCIYWhORd7BhJL/wzCL6bLCUwvSefpxjio7+ajta6PEq8mq2w8JdPi
WR9MfGWXran4k43ENNfw6BKZNmfqgJpNsHGQY32nv1+d1ToYaGmab4CzWRzn4bYB
xfaLudswmqWGxoEUuwwpV0sn8xRdxDODLDkZc/+/hzrbymiKZCNoTDLcHNzXG330
mjsdDjlNXopwnit4zZ+zKOSZ7qtlq2PpAejvAloCtEkotUgJKqohnFtNn0uLadCT
QfpyH/Y2JJhdT4cQnRsFeZ3n11h3a/MeTH6OnzJweNpwWPZvMICUZimnEIHp+ylT
EWupd1r2Gd5ywS/SigifCCUn5BDS2a7NjkJ+9RxtwIjX3JOAReoLr6PIe7EaVfHC
FzmxaQB3ao1NEVGKuAY/ge/Y0E8SDjcQYquHE+DqV/2Mlp6yCR+ISOprInqty4B9
jZF7vZigEpTtOkzC7HmZKg5bvPeiGOkcKkhUrX5OJ0IOVPKWRnO0WVfKD2ZJ4E1Y
Qh7/o6OMAjgf5rIbCVW9KCfXKdNDK5YvC/H0xt2+C8gJCpsboIJyT0/hUcm1IiYc
NzjL7VTNH6N2+yYpNOh9UW8RIcks06amw9QeOyRQNfFbNwQaSdrE12nGh3S5NtB3
8oZKayybzs5jZKSt1WFKNYwfrvIWG2liRX5QQs9+t5W806LFpls0FcpCgsgRNm3R
37kZrIr2mouxtiYj6WQEqa8v+MhmOXFQzGkXHPXcGB9apNfv0ZTdRbbqv38ZC1f1
QZsfTfzoi9xga6NAKl4i39v8+zArval17U5GahZJ3LLAlMtsNGi+d8x6bTfvgukF
rdv7kU/r9PrTsk/1jGWyfvhKHanKFW9h/JEEtd2z3U6t0adN1SPsCq02wpcAh6xp
weoD8jZHXXkhKWsWxHWpihRV4P2ppdn6XPZ09wCVRvwwyoUoipLyemmrjT5MI2xO
oGn4w1GX74Of0gKmcU5XfzCF6OXdREkaYQtZ9WNyF41zLSzJGxjnEwulRri8wweM
JaC+vW9OaOAlsqR58na/IOmKnHyyegnikYpnl9UXZ1XSE/TjlvV9pLFJPdqJB516
Hs6qzQf2sOLNpCehiBmtwqSxLlTsVuQSYmE+Y29KT5QzOz59UMor4avJ5hdrqEjS
iW/9BJm2FLlhrSycxbovomHMAMXBlxgafZQrDXfvMTEIDH5haDFbRC9wFj5MUfTC
nclGxgoKqtV8US4jpktlC8ClgrNpxmecqMx0tp32vhv3wmayJekbZU9pDgEncJYI
zt05vf/uVDh5XNrRkrkDl70kK7zK0FMjXF6VHaNYhyB8XMDnJ84bHbSFPgxwTKSs
GGc3jWPlqpJ18aM6ih++Kv/hn629u1BvC+MH9Hjpv3ha37A029kd+WKk3B9rSTaC
vRclx7MGoaR92cs3E4yOrMxZxwYF/tPyeDKMHi/BT+l+LS12PzWrdQXkPz5wPN7u
AIP83NxJ/r7X61avg2ROxHhnq+tA9Xqj3B6Cnilitq3Aniqg8cRWqZOUwf6cYILs
UZx4CGBJitHe7Brh4iP+13BsSI7D4HUNgQdI8U1LjWHkH3oBZTszxJKXLkFYfvam
fUKlq02K7f6x2fh/2wgt8dmyhjCoNItN9VExHThGUv6nSryGI3W6RtE9T0DIjGDD
LoHiusUWrG7XqpGH90GIPAYN4C22yGAOzuVgQ0868qmmuh1yfWEYqO6Fy2My6GCT
VebtbBqkNmlp6nM0a+mkpuDJdMz6Xqp8jTwEnJsBv6ts4qjIdBvK5Pbwa+ZkH1V0
hXkAZJC5OKbCCt2lt9VOD7+U3SxfvCaec+sBUj2WuOrD4c9OjTRq/vwQuln+VHE4
zTk3jmzAZ+BghnIAQcBWxqRM+IMRq1GM0AEC0Qea5C1YJ5M5vB/0pDkc1N3CZSxW
b5evMTsMsG+8n3TPULNXJROOJSrYlgsAmmn3cQ1zR69JNHRbEH8IX7Rc5qZZCS0K
YeAQj2nBEeAkCxxO/0WNKJQiASwaA37fXduW4R9oRDcstofF6ittQ3tZ4AotMZsr
0lJFdKOjpI4Jwz83Ia/gp4ea6aCIvNQhiawcB6OllD7cSB4dFyzw+mVS0NRnWNG7
cJlNCRHuYxSDIS+FRltgfUzldwsXDGYgwD3EtjSDPNKwDAsAGuYXjMVSrEjrigsv
arW5zJyVLtZkqWIHqWn9p22k0/JIg1gDExdrllZYQ8S4iGadN8TR/KrdNHjZUU27
msjCTDC+0P+aIzawjKTQT+ioLynLOjUfu4DmahaGxtsKrx0q/PONHPXxPHbpUehS
5SPoP+Xle4ZMzSP20B15tIfoLvm3d7JPu20iJb69t+2XzY1Fz/puwT7CC3V5Xuf+
LJwrEJ8eipFt/dyfxfcJTJoA6/u1ZyckgFkwLf1uSYcOPNZm/uQkAKWvS9lSJPqB
JEID/F9l7DPeF25eMRK6AqH27W0vTAw80uHCsoOLmthDW8WRpiD4F6YqDF/5ak+1
8/YPxAyJFr0zaw/W/Hb/VqhSBfugYH1/vl0qBJnwf9Mfi072Y9E9I95HIECkNIpu
65i1/Eg/zVWurtxhrxHTh01amrf4lGK0WViAB8UHXgI+ZugyhpHWIP95UXEJVy3u
`protect END_PROTECTED
