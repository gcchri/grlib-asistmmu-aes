`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
by3u4OOscy58TS+uaLXsV9cRumIHc3OjHWahnLs7Drvoy7sX1ULWUNPHpr5jqtdR
+78HCHYynors1z1+vORhkZJnpKJxrc+n4X/NWdCrOz6ZtpGpUE9w4oVk9yojkaQk
XAdu/5YJZGH1x1b95epUo2fy1Wr/u+pF3Cc/qt7LgbqhoboTsFWOTW0A5+nuFv5v
/86cDs69DFWysC52s1WLqiXJpgOqPybs4iLbabKHCVzmeZtJkRNODHPjC/u1I66L
yIeGjr1Ks7DG29RrMrtLezjOo6M6tKCnzmEUPhc1JYk6eP8hnseV8Ev4fsTgAP/P
W6WoSfxvXi6be0jNpW0D2xz9bLYZ+AXu4axEEnh5mK2D27iTfL9xh7yo0wQTjQJA
HwUi/iqoM5+243fXEu1eTm21j8ujWw8kwbVaZfVV6YeuCTjl9x02NiTvB8/R2X7N
L/xUqCXKdjk0zvugP+6bOW848/uOgGX6XQ9XMxk6CsLEQD29qRcVehLJB4KOl1G0
LAb52TBFH4DWFLUZlWNcjWSgOlmQbamDK1ntEPZUl3U0HcTsEPGVSrnG5fEeG+yk
XqkRONaRFymy7MOLFPF4qyNvBrUYzcd35Fp5L+pyUb/5m8dwSOGc5if/pgA/ELqB
xbaUnH2fdlgoyDc/U80mEZgpA8VF3nhPqkgUdJGMhnvd71l4NetnEuVHUs9S6b3I
qrciIuZdlKVI4JaMsGu/r5KthtCIn9fxtWWGbqIOWYCBqSA1skfJ4KiWx9Smj0z9
wCXfACI4jFe7ANBNiVCVFw==
`protect END_PROTECTED
