`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EsexZROXFtg4kdtLEUjbnBdpLKuzPrccj9iC34b+2BuQR9NmQ8ECDUprL8kneXb/
QWwKGtFj810z+pOs9aiHFOWXm4/j9l9K+Qw6O1jFSE/T6monuCVTUL7yFCWJq5yl
b2qLB8Xdq4fNq0k2s/BOw71bW1X4U5QN4giSobQvXKZD2wHBu1VGvniRj8tJ4Z/x
vYUfS9C2LBi7FtC+ZlNDVzzAl5/+aFQvbYhCL2dw5kEMGlcusYryequqHuiqUGvy
/3UX2zBQcw0gYfBwp0q5mA==
`protect END_PROTECTED
