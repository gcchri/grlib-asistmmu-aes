`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lEMxWVpGh3XZVdandmW/vP5cZTvybHarLxUUonElioxW23SqwAg3kc5+1wsZesyj
up9KaNNN8z9UHYjLO5ddHSSO0f4LYMtzGj9OtVltUj7X9OQ8bSqNWGRsuhz8Rk5N
LZR7DIj51mZqf75+8uDzYYxtY5eMMqCjJ2LawLr8e9WFvHxb9FAttl+76iA+/jxi
fDlSl8ptouP0TcXvHFNVE8FVbyEMCis3AO5j5puxk2EbzLnOqtPCAJuTynNfD5QJ
fO0UVtZd4i2Ypc9q1jC1F9atmOJVYVd4uGvyQru/MHUk/Vj7gqz/kGNzR0jwvqZ3
nRHdkbIeI+zotbNzWsFlWmdTKDcLX7p+NMcEmg5eI9FH1nAfZ/xMHQ3JisY8frVb
9QbhKOJREIxonTvMfqK0adBj0UrmTm/m58go19hEPcSwoS13C232fSl44P08fzOR
3RIfEm7QfXcPxMbeey5TOCsja137snmdGY34Jyqohh/8RlL3vVao948RduIz4dxV
2AJ2VYRAvzoiTzzboC0YSPKoXx5GJ5Bnu3YvhYt80yw=
`protect END_PROTECTED
