`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GeiBtrQdtDkCcAJe7ohXDwFfOycH89H8cNkDqpWqBxr+OdEnUFREzITpsgrFybZ2
6BiTaEO3zROI3+QWQGaRwo6r+IiEs5W1rTby+psYeYw7NtRQRLxElIzE+8q61Vgf
60Qfe78WgHjY55cV3hLBZYc5JWUzZKds1Ngt6Q9TRyj0vUzlIi/mtaEkC2DBqVOz
EDJ9AukOglVMkwk1posB7PYcCFGmAvcoZU9Y/LPZy4qcwj/jilcblzp1hkH2St/A
nEhwBFRLHaaqhepHIuPaCbrueln9EYF9VNEvRwrbkzYniO2qcSc6nvmVC+G/8xyA
U1noE+L71gKlKNQ5NjKeJXlgCp7gMsC92UePEbvY+F3ekfkmXSGtGtkJB3ZEpqii
`protect END_PROTECTED
