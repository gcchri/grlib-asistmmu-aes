`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgIiQ3xHLoD3V3UMBV8HP2/kOPfl1ZSIhpz3FdkAkg0MDU6TEtJ0gZB3x1udgs65
/LNvBn/ZOGEJt4wDcb+PiDpTTSJMnKfD6WK/ekWGcQ+Ho1DFZz3tg8Mjhn7UAjQG
vYzHcUgWo4/5jC9UT400uZwbeJ2+Xpz+UoiZWxI9/6oJSZmWrZFl5xsSueRg3ljS
OTeUwygFzzidTGe9O6m4y9u6b+zKFwm+MQ6H5hZopSSsWqKIruxY03GY5Be5jfIB
+/wqi8sT8z16hAfN51L7i5k8A7r7Dl6u9QAFqfBDAajf9qQPE6AXuD/rEHY6Gbbf
D5y6InHXWBfiDZ4mUWXTEvCqy4G+OD8dsY1vnyTIBbARsWWLesebLmL9T0xAsBII
++rw9nBYM7zUsZPSSCvxW9FaUH0c/aooHURqh2MGO7aHmfqW63ZazrlZ7DUiUiNB
`protect END_PROTECTED
