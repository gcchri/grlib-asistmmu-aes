`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiODC4/KD1GUWSxPeEIHC1JG7alvnTxFjHXqHtm+A8TyEhoHWdWJK5Y72bL2F/SF
YYW1VtPtcTcostFg+9+VsGEPOeUJOmxB4q4dQETr/ivCQ8Bp/ncI4wOorUvdQmdu
bhCBD7bKkVXn9zhENOOuw9JnTqiQ5SEh4ULaFXHufikTWHAjUnedRWL3rTAiwoft
FLm7up2kvJhYZBsVTeQ/HBF6568TCRYGhIbo3vJ5AvIppoJzXCytZRHnFtviA5eh
ti2XCDZfgm4M3mDJEAapphrRFPZGWjuHFgFfXy2qQq4ntXdYLIo8wATYQ7Icex7Q
K8WkJAhfzRQFmqo1kETr+nl1x5qvn+T0D0OnN2CR22ZVRo0A0R+IroYNcfwuL0Qy
SEeuLuRHCqEFCnNfs3eYcQ659ZmU9DR8pDU8Ir90oeGnyMBTcDCBP10816LxysPh
gb3lQC/DM0myLJA6pln6pU54qfJcDSAODuflmfq2JkHuW4E3qGAmidVq7Uo8ZCm6
jOxOi3bDP9YEu8Ey6QyPI5XbIgAPFdP2LS1kXiTQvoCkhFpvgZj+fuumsrx9lZth
c69HxJ3iIEhgmkc0xW2eUjgFUlqwS52OzQZoaKvtikfpNfh6RbrULry71hxWUgoQ
ouiHQJX6nBIc51qBHSq3ELcpEA5NkC+ILMhIasJdIXcWXnoqiDVbTRnyixoe+a/a
f0mbhiemD0A4+bDjub7EMLKnHAHE/6h9K/puRXU+OyuRQXmShdp8NR5S74rc3u4t
0CR/keX8QTLgulbOwuXJpLPwRTvCnzhHxFw4pNdv/wU63pO/76KyIkIE64m1AIUk
Ju0In8XYiigHHPKHQ1octj7xd+4MPz+W6SCYn1igAJHqA0UIRxXpr7VCxNwTgX61
tDqSyCF0g0dRvbTSk5EF6SCvl4R/xatewIRuT5yDygMoNTBG2hJ0H8MwCtd6Xv5o
6AvWI7rjIQ/9fMEr0Lk27RKgL5MUSTWu2hoqaFIiqR2Ff5c12goC2rPj8GPJicOJ
IBHhXdjpVlaA1lZVLcEVillQQwnOVhRkNK7jpxuF0K7RgnGiJai6RUqK7Mu32AkF
Va8GUX19YT8UZP5Iumki/rI7mP3I95xVHJOTzxOyBd2Srk/Fl7FMP3tivBy3cRhz
7VlThMVuHMg4bRs+OLxIuKIVhjWeorEf4B9KTV/y6J+AozM32EfrgAtzXJRSAw9a
nAjd5rO6YveM1fOlpyJGJ5Oq03cJJSzENPiTv2MVgb5Gb7wlYCvOaDb+xqRosZ9Y
9j+zd3pyCicZpx7bLPA7mu+GTCGGyFm6K6ksDPPm14veM98a251UaQm8pAxgYt7j
P1LOpAHP4fSpbNI8Ldve6w==
`protect END_PROTECTED
