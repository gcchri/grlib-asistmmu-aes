`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3fIifyQ87GwB54xIwbAxj6P2/nagKzG3Z9ReCrGhwCfxms7RM1JeeZOyYQ5hUOC
dEu9t8Pm7WUt/+u05Qrj6uH0OY0IYwaaHyFKuWGuWicNeX6yU1nZuzNzyEqZaao+
zO41KYnTvJUMRA0t+cxXPAayQ5qJlOGB3L+jLUkKqrUKeCQb3c26SQiTKyW4cA2g
t65iV833rU9exNFemk/OJVjEo2qMn5Z0iu3uuoC2Qx9EAUgBjXbP83/tHMI0JVT6
c93x+8HdIE659Ynuqjk0nPsDalgVbBKst70rEuaxMqlFFmAhF6ERNNEEAJCo4yn8
QW5BUgqJcsFr5h40NXEXPqgC7nT0Rn15sOrG++n1O7FUl1hReNZ6HG/k1y39tGul
`protect END_PROTECTED
