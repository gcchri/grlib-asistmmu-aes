`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djuDmzJCN9dwX571mpD2uW4lFm0IlKo89TsrbbW68A3Pa0Jb50Tevv4cv2Jo7N8y
l0GHB2XYAo737b43kIpgTQoXLLeOljUrBaoL2Yr4YDmAupYbD19WD1wagthwZmSr
icJ7MGQuzv4JG4tiQJZAxr4608MELgPzIHdKJTnn4DA45Y2f5WONUDM/6bISaNVh
jbzzR/VJqH/FXRhKxzheWOT4nnLjae+tDMAG0HoMKZ4x+gmLcWAKG56/tEN3RJj4
E0W8DH2MUz147vf3LESsqqnN9c1o1z4mwFAoedxd0bQwYyga4KcEzMgO+DmA5t4n
Q8vqO4IJfF4l76asCzFkkwnxoMhqFlfvQwjjeeWVbnHWgD3PraruE6p0HqE735Q5
OBSegpuSyGwzcTDvyp4GT4WOtAKt4e0rtUoe5kOhbvRrAipsCf86Q4BKsI2rnOpJ
VB++0ITrHG8VK0vCwNU3kpKo69Pf5wlYhUz46QNHES584NWz2rkVDXEatJIqZ/4W
44ojBhaomvnVG3M/jsOyRFlByQ9deGJBqNYZvoOnRhacsmubowAZrLZlEjBqA+QG
P7S8wp5Uf2pHFUtxQwm/ksAMKDRAzrxLPOR4SjwHR62W6T8FreXp4AI8R8eLivK5
9jo2EYq2BIjD32yX9oBFjEdhLWGlVf626hZQM1kozJU+R2SGZR1cXsDAzTquB/FY
psWysNPKu7W7n2JCgLLxxxQ1Qjc47eTXoZtP01DOvpPllbliRP2qiFe7w22Gcefj
4tHLeFTidm6bkj96TJahn/Ecuz7zRbmZqi5RvHY3dwt0AE4sIUuLWEo/uf+1T6MW
VGRTBT7W0HaWl/i9wcnBebhkNFvnYIRUlE6UmMxKFPvQA43WEK8J6BImZKhljZrZ
ruaUrrl6Uwjs425qUmB+lO+vgpQBruKyjpPxr26ege4097JnFMB+uaJw/ARHe/cj
tWRqxBgkLgIESG489TbCswlneYWH7+OKKWhVf7pl+TMQujZRPsXdbK0V2lICO2r/
+W5ezHsH5+hoIBl5wmPFg9q0fV9sthxL7zS3x07RGPr6pwekWgPtvvx7MkpN3oC4
8MSON+dlKivBtkh6gFPubdQ08klFYNpfqZiTdmY/TcSDporyup5IoskE64UzJUjj
FWaJgK2yUCWNn8UJShxG1rEIX+kPmOth2/3kmELva20hbvNZ7U1DFVLfmYEe1fz9
7ZYiDnWbMnz8DiVQjec2A9ynHKwL9qj0n66AVThXumUhZJbrpdj3F/9Pj3royK5A
3ky9u5Bo25mHximbM3FInFqEmpYA8Dp/aYmLkBY7wPp5snSJxzhmqmkIxxv7RY01
LbXIlQXrW/2yLutj31mJhkPOXo0FWVRBzEnkOy81JjV+lkvQ4sVJ061gSMs1aObf
rQvipHh1CMg5k84Kd/auvTWjb+fzCh+qjBWHRClXoIu+g5usVepAYOPnRfEHtJM8
+YLcpK5ssncz8i5n95m9Rp5G+4ZHpIGMw81Ssg524QYMXBwBsIFhXSIO6hXFXXxN
GyioIzz0O/o6J8EYwJvle/lEd3sqGkEMcZdYaUmyVUBVFlaf8O7E9i++5ZChEhbS
WaviCtqP6kiBrLk0B+QjyhsBY9X5q2qFCSdHxjxA+XBIffFsBmNhAYJZC8OgdEnE
BPCGjFcL3i+BwiGi+8dJ1vsDkiybRZczzdxZVnZioyg1TkM9mLiwh4ufFIpj15Mm
nJrPzft/sGJCiwVK3dySke+/GaiRIfsNfroMreI8CFLTL/ZOWirq+IFCzcFCuchR
B3ZFP3gmxBQFFQyRP2IAcB5SunW9tfrplwiSyDOspP4/ZepMItkP/X4xe+IY5tOF
cwL2FvtAiXUpCQzNP9q98cVgdYRW7MMO5SaCqNw/WmxrsxCbeqHPmLRWkcc+EdzI
EgVFfK1OBSjDAWBcTfhbauzOWUu6ZGdEN4ljLku8K+Vx3/7zTBY6Qmwzyf3IK5Lz
9WK8iEjUPSPmFp8loamVPnLTH4yILlgf/QtpALEWAnkQPgfKuO/ASApsMdjPTnnd
4jR+FOIqZoB3m27Dn3V2zEfkx7qbmOcVGDsthwdAHtx2PiEad0MrhZZhzlFW1Hic
/uIwOioXemB+vqQZo2rDqCOrcfUCxaHZypiytqMnxRdPC8RWLFDMz911+BoQQc0d
TzsU9a9zt/Af4c/wN4cHj13ZuFfktAFywa1+dAKgrIicquyna3KNV3dA2Q9NzVbG
0/+AYaPsebNRVHkefGZmbPLlVUkEhmxQERgi3cgTp5hObAX44Yw251SB43NPgrEt
aPqAA+VGsfkLVd6F07Sh70e2X9ZvOB0wIA9D4RtNmwjH7vxf30+Tqf2gCeZJJMhH
YyBHYAyjtrv7RJbdbDs2h12NXUrd/NWQQ0/2aX7bJGhto/3MegY1a1rhdu/O6VaG
gz838fze6NXZ4lVHh/71YXBlua77nGf+9uwFjha34fSpCzopSeBx0U9lP8CjnjYm
FstetffEQYrzUbjg0csP4CYB6ss21/gIDvMysbxydDvy3awliTpeQtLCPG64S/ZZ
4sDZ7S0B6ZQo0/JTo86v9IeMPi4s+oQgtUS5ZaYpM+DYZ3HGOPTZjj/ebltR3w7i
i01HIJ2CDk0HGQ+L+tETLTLyO7wyny1ZEnQ+aCKN5TzGgqKu1bF6zEnjvyWXVz8V
y+e+JkcO2ZrtB3xNDBV273NgoKEYdoxCX6Xv1Btu3y7zEvJcFFjJGjziUkNpvtmk
t0pwjsUSPy/heF8LXpIR3czoIHUsQyc2mTHXQlbzDVAgScdSS/05x0Qv1pfWc5wf
ikXx9quQCai622RjUvWkEixBW3c4mTFJPG+OmXFHfmFxkp3mzpFu9jvCK3wp4wZ/
TcWIfMoyk1ZM09TwQ7ogwM4gptL7Tl8DWxkHievkt1va3pPtzosf0dGql1KddvXQ
gZCGUacGvyzcZ7FN+25gZuhXbnRwGn22+zcZKS1q5UMx5dUvxO56xYg2WueYoRtw
HA++jl9KwApfAEe2NIlMv+vkwUvIKy+72VrL9dUH6rGtNufodKnaFFGCiDwPjmF6
7AIB2Pm9YfLQ5sEsL53i4jx5F2vpNFc1ExFAVSzkn6kUQ60PSUE9/h7jgva2OREn
mA/YZQDJnryx2QfU3CCN+RKEj9Hf5nKKLPg/Mr7sh/cHZyiPSVklUXJFi1Z7OeuJ
t6lu0sjus/Hn/D2R9ATA/626GKsRG7FSV9wsHoSwpJdTFrSqW7o9J11Xu5sffYnM
m9fNfc4DqoIjeHiw0FpvhHg/fyaf3Eg5aseY/SA9fbA0W2mpa1KjxaQcqTIYs98t
6hCoSo/mA5SJvdOyCqh1FMWJtv25YBhp0+hgiSkh3iLpQRPvWAMOfbyUT41FjfpN
NlcQSMS0VxObp1N61aytRO7JLScCcyPXaCAxmjT28x6LbGJ/1ayj2v8qUl/dnvIM
1aDrtrOMEwREPVglePcSLmVz7HFP/dg1A2rCL97XBEJrsoIjgccp9AtR98NTjKkK
DyDWm3ULcaV/JKlmWnlddrUEvVVyg95xtI9cMTrAf7G1s/3Hzbu/Dr9A6IViSz83
kaSCJWs2sGluedXCzAuUJoBGTP1ecUphXdRy1AZF9qrm2B0lrniq/4VNzJyr5XHK
yfIhSY3iEAkNvZd0Kwn6rJ4PiK7f8ZsgmqLFl3Yqgke28ZSMZDjx5dNHjPIBZqL/
lLM7x2Y7h1C3fCjAnKwdUBCUV1JOrRF+9+Z2Dv9V4pmm7FlA4dI0vtfq4iXznd7b
XqYCHfXm8AaFHtDeHuztZNzP49uPkoi+hE7sD7HdNeVArfakOn08xUcbivMj+cNa
2qaluoPLH+kpT35A++73qmDeN9QG+k2kYItEb0WOY/ovn2OzGZjTvA9EHEZW8faj
oZxqKY/F+nQ+/mSQVoY1SDSoeXKMllnMlpnc8ZXMxe4ISadLq7mT3QkUqX66k17j
dA5XMtxm4r72xOdS7iHvzmXlD09d5Frb3qm1zpRjsQRJBBq3pa1kdH5FSuN97+Aa
sngo29YpgYteRJeGqfFEmS6uovcHmDmeve55403cIGNAZwONCJsCTAlQpTSv2ols
zLSLnT1pZSsM4CaQLUKAqrgb9llKNtBeW5DfUYxnv7THYCaI9ldFFLql6r8meBez
kIu0wvi8kQgeqLfo+WjZrQ836w52fDD0/7oxsrg8vZHTTTSeDthESSyHvf5YZE1S
BqCzQobSVCRXAS0rtHAOTa6x1f5LuO91dFKFDdfGKz5I0ni8pyj/qpZXg+muXLMr
OpF+pQsjGm/NuqNWRAnJPiH7Y4nHFwrC+8uffQB8d3YCvb3Y3cfSbDExQLNYadiK
kb1O3JIhB6HrjWOw07uBfoCFhAcORIRwD2kFyaGaIiZQp61+llStwjoEoyw/GnWp
M+nUHri2ECaFAoisVNI0PBQa5V8Tb4CPCbK2fFK2KlRNSwNO/bD8KC7Pqtl8j++0
TMaGzZ4xR2YiD0KdJMEZX0mKCRABZ1bTUQTJgEoNSM3Hz3FMPZF7/nlbD4MW2ot+
GbaV0naxeaNoVSLFcUpOZCMx2mY2CSh6GbeijaZzYAT/HrQNXz/iH5yxxJ8Xip5r
P1QAZgGH7fFFBvY8RL/rF6T9hmoH3l3Io1+GrIgnCdp1wVDcU5Wtgyt+9lGp2EQv
miYkoA4NUmnSp9ZIyGapUiX91djQtD9eCSAZN3IraOBtPAY8EweaW1K5YFuv6mfZ
D5bCLZozh4AVu0F1gECEuj2XFyZZM1H8tdd7RBb8koaa58gGklBRN3Cu4MkpED9b
3nEyUskzb6hZiJXHoqGIkqv7SGO48v4NhKj9tDyAeiZMySrO+Ws9nlyUWS+nU4en
gop3l/9/T0moB38Yhr/yjMVoD5TIcfK5JWkUJVPtNurRggw4u4l0dwD77IJjQl3d
6l1EVbGvobwn4OuvTB7tDhz5bNwezUuaF4PiSyCTut0BfEsakVqORDjDX7avL8qa
tSSZZP/Es/waS6hdXnovP8jn5a4AkcVAwsxZKTFaoU0=
`protect END_PROTECTED
