`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8f/nGd8bsJeZtnNUSEGy/bOz6fBuxzfsvL5p/t1Y8GZba7Yja153Jb0b4C2wzJ/B
qNpEJik2nQr4s1hyZtKpvGYsbJoiRGYbHxHa3kVpp7L1NmqK+gZoojTBE63SMGk6
oExXdraGCoLDbd2Odmu3jysgmk1Vb3Rj6HCc8J+PrDP6Eb467rPeAB8tGkVrqueV
mGd2SaXZLWZ66660vxfHfTnoZ0KSMjxu9WIJBsUTY03ztGWHmTz3ddxF8MSJkHZz
fOTkwjF8H/lf+hkCge1ZB4Hn4JRlFsbXhsTWzTuUHWJG+KmiFEoJMaG0rsPkvCvn
1XMKqVHVlLpiuBF/mznmRm+QEuWNCGL0d2wRDlkkjFMpsJgleIhsWvstM0rE9Dgm
WSkLlPkihNPKsi98Uvlc94LC3QvzqEKTTohINI5t3zrGyVdnD4mdKJFGFUAgmz8d
yLRNhsagTlD07MqF1CjdQRHqIqPU+3QFrpXV2Pj5ktxwEH73d5TZoRFys9nQOdSs
lLOamXjDfBMDbcmwu9aYBkbAhMPvT5YMBrL5JwKMREhYdro/v+KRL7t+OQEWUzXj
PjMwl+w4SMWZkjBjh5/6DbB4nUFqleiTMUHfAn4hRCkm5gRi6R8m2GKFoXg08FrC
rNL/r8wXQFyUs0Ac5JvsEHGzPjYOEvtARW7qd0JmTLwW3LETfN1uNSI1vUXwEen9
1QUdH0KlbrQG1siT9FxX+YvHV8mfRNKm+OQJAE12f8hbslAVsJ3S5T6Kpkaq3DhD
j//BYehsLlSiKtVRAS2sy6OA3ai7T+OpycxnpsvbOfHwrDF4n3dWnr0tZ6g/zz6j
2bmsdmvob4JqHcYnr5O36ACY8fXEWik1aexhfpKgOrnyy/M3NtZRBKAYK+1BHqc/
j2uq1D58kmmPB8wDT4wxCNBeZSTrG+HiexDG/AWxCFi/b6VUplaEVGX4AmX7vLCM
nyhQOySPDnHQrdqaXIFH2qUY8bCIxPLblyNTXO8506bRAolYl+b2415tYONOx7bl
GwfGftiDHLJSWPyYDbkiQDSduwkKOYUN6O9hGZIadx60ViSsVlZvXp/OpQxLqTuc
WScbGNQwiWyIeQKKlZH5c6zF5pUfMolEys7StA/xAsMRM1LA4ud61Xq1PmyWe50z
g5iiwcKM1T4TJfDFUZPaE/LnZpdySk40ZmVa8QUEwD8YnKM8bnYMdt8c1hlImTLS
v5s+YO88HqiL1AfTHq67zjHu4IvPx2zQCZM9p1pTQq62jZUegWPL/J3ehYVLVnEl
BKAUeGjCTg0zUmaSRGqLKQanoK9KslOqm3kzKEw/m3Ipyu/ugrsBCUYQWLRaL9An
mGRRsbx2xI9MOMDGB84UGUweUyp+sohJq3MdD9zXPRQEsO2TY8pradoElJlFQW38
u1YbWiCNlAhO6v87YKt9WnGj9mInZ3R0vERMlmCkTbTKlEcfZFnIMSy7vQel5IuF
pAEdYZ34xv5eM8LZXghgTxabNCwMq6s6PPstcO/gnueJiJA/9bXuvISYJZJ2zhMc
Kg9TKWpKiOAPLRCSYWbLrA4xtluU6D132RxyxBeAOxxEF0+cW1XYm0XdTgztdPld
56uh42QWKMpkF+fxGUoP2gKCJwB6Yvg/3vF82vkvmbcROkyqGGe9AYmQ4VuOFXoS
HMFciUgqACfnOXnhJyPECYVk2m5GywkuU5kNP7mJq6ew55QLSIX+PCejg1Iy2S+I
OsLYUsfxj+UUd3pthFR0yyKEfpNxdMSFOeXD7u+H525ZsSC2Gg8yIT+rD/EmbL8P
f+2RJcgVQ0YQCIfLOogWsH7A0+RTrX3kIXXf8g5r1pi1uccOhNGncIHa+/oAo4Vd
B5uK4YuBu+7QOXo6UaQ9jpXc1D3OVU4I6/pdkI/ftx8HACsdcKx98dN6G7U+94RE
WCCK1cjZWPvDq9xTj/rMGBoMr1WjBnjexAYDbM1T/Po7G5qMBTx1NNhYTfKaqamC
V/ONZ0wvleuTXYc9ywxCtvyBTIrASWpz9pQUeBjkCiE9gPz27lwxQAb/muyATgdt
vn/LsPxfd4kmGVafAOKCEzDZX5DU9ex0O3OQBrA/cdIpYp3RxD0f6VyQufQJ+9Ez
bC00OzRwliGfLB782cPRM/uQvKpPX/p6TryqwsFV9AbQntO8qZMbzBAyu/hxumFb
QAPv6RqcRjMPfnBQUihWrnzDmZJYClMU7KD7KILTU5MXUkRfxkffjC8Lt7Oha7Fk
FEqxlyDEwXKzRcBkK+0SwTRQsJgqy3SLAT9FCD7CuxVtKJqTit8BdNAPbs7qkjcf
R3037x+TIYP0TdEHdf0M5TzmUcoSiXlX5ESZx8FQqynylXGNTHm885yKyOtTEtkp
urtkym3bjGtJgehsPtajnsoifHodLc6ktDLPROaDRglBvdfOU/9pn7TH4d/bgAQw
NrRY3jJShgpJsQnSGWAthJMGtFUdwg+IhnEtDWbMC9KhNaXv9wVas8ZMdQrH9xo0
YqyUrF572wpS/aSbppOQcQe5ZaWkFuUxjZ2wTNQNower+peafD1/hhf57SAgOIGh
IXi0Vt4r47AjnlYKgdHxJoWAzML6UerKm54MgnV57zw9DszDEn+fq7sA7+ya0a++
WgC8uTo+UMwqD7Xc6RvMvfHdR6CPJ03Az7XXC8KHYKIfL06+NaaXBSrVoqCvv94B
rr8NQVv6Q5W21EvLITzBjT9yE9uIRlFb/sWbBEf3ezlnpwhB5jgDG3vQ6Jtmcy7l
IiYrB9RXJMtVqvjMogIDaQxFUjAaWSMLt1cAY944dXbW+LOIzEeLsczq9R35Pzcn
gROvX2GCSRM06NIuwrqiugNL3g4Ft+a01gEgEj+NTyxzwOZmpVBX8sV3wAMRclAG
IJ2QflgV7OZXHW6q8/3WWROsrsPc5mLKfOJYWOu0tNjkWq7hmCp/CKXEvrc+nL+m
Q0DU4qJQ+AeBrsUcboD91hagc09eJuLLhbN2Vx9V2rgE0GLt+gNV4BAz/foYO72a
ruVnhuAUWxPj0lg6LlbYsuPLx0Xod//7pFbZL6NHH2roYOI4Jim5ssJ3Yioa3iW+
kvlPA2tZgDgULOH4HaILvQSxeoQ6xEJSuLKoLQ5UK9w965fBkb4Kkn7glvcsRScc
xmT4kKWgwlBNtbXZ4T4buf7F7DY24lay0kEGEAYp6X8=
`protect END_PROTECTED
