library verilog;
use verilog.vl_types.all;
entity SIP_PHASER_IN is
    generic(
        REFCLK_PERIOD   : real    := 2.500000e+000
    );
    port(
        BURST_MODE      : in     vl_logic;
        CALIB_EDGE_IN_INV: in     vl_logic;
        CLKOUT_DIV      : in     vl_logic_vector(3 downto 0);
        CLKOUT_DIV_ST   : in     vl_logic_vector(3 downto 0);
        CTL_MODE        : in     vl_logic;
        DQS_AUTO_RECAL  : in     vl_logic;
        DQS_BIAS_MODE   : in     vl_logic;
        DQS_FIND_PATTERN: in     vl_logic_vector(2 downto 0);
        EN_ISERDES_RST  : in     vl_logic;
        EN_TEST_RING    : in     vl_logic;
        FINE_DELAY      : in     vl_logic_vector(5 downto 0);
        FREQ_REF_DIV    : in     vl_logic_vector(1 downto 0);
        GATE_SET_CLK_MUX: in     vl_logic;
        HALF_CYCLE_ADJ  : in     vl_logic;
        ICLK_TO_RCLK_BYPASS: in     vl_logic;
        OUTPUT_CLK_SRC  : in     vl_logic_vector(3 downto 0);
        PD_REVERSE      : in     vl_logic_vector(2 downto 0);
        PHASER_IN_EN    : in     vl_logic;
        RD_ADDR_INIT    : in     vl_logic_vector(1 downto 0);
        REG_OPT_1       : in     vl_logic;
        REG_OPT_2       : in     vl_logic;
        REG_OPT_4       : in     vl_logic;
        RST_SEL         : in     vl_logic;
        SEL_CLK_OFFSET  : in     vl_logic_vector(2 downto 0);
        SEL_OUT         : in     vl_logic;
        STG1_PD_UPDATE  : in     vl_logic_vector(2 downto 0);
        SYNC_IN_DIV_RST : in     vl_logic;
        TEST_BP         : in     vl_logic;
        UPDATE_NONACTIVE: in     vl_logic;
        WR_CYCLES       : in     vl_logic;
        CLKOUT_DIV_POS  : in     vl_logic_vector(3 downto 0);
        COUNTERREADVAL  : out    vl_logic_vector(5 downto 0);
        DQSFOUND        : out    vl_logic;
        DQSOUTOFRANGE   : out    vl_logic;
        FINEOVERFLOW    : out    vl_logic;
        ICLK            : out    vl_logic;
        ICLKDIV         : out    vl_logic;
        ISERDESRST      : out    vl_logic;
        PHASELOCKED     : out    vl_logic;
        RCLK            : out    vl_logic;
        SCANOUT         : out    vl_logic;
        STG1OVERFLOW    : out    vl_logic;
        STG1REGR        : out    vl_logic_vector(8 downto 0);
        TESTOUT         : out    vl_logic_vector(3 downto 0);
        WRENABLE        : out    vl_logic;
        BURSTPENDING    : in     vl_logic;
        BURSTPENDINGPHY : in     vl_logic;
        COUNTERLOADEN   : in     vl_logic;
        COUNTERLOADVAL  : in     vl_logic_vector(5 downto 0);
        COUNTERREADEN   : in     vl_logic;
        DIVIDERST       : in     vl_logic;
        EDGEADV         : in     vl_logic;
        ENCALIB         : in     vl_logic_vector(1 downto 0);
        ENCALIBPHY      : in     vl_logic_vector(1 downto 0);
        ENSTG1          : in     vl_logic;
        ENSTG1ADJUSTB   : in     vl_logic;
        FINEENABLE      : in     vl_logic;
        FINEINC         : in     vl_logic;
        FREQREFCLK      : in     vl_logic;
        MEMREFCLK       : in     vl_logic;
        PHASEREFCLK     : in     vl_logic;
        RANKSEL         : in     vl_logic_vector(1 downto 0);
        RANKSELPHY      : in     vl_logic_vector(1 downto 0);
        RST             : in     vl_logic;
        RSTDQSFIND      : in     vl_logic;
        SCANCLK         : in     vl_logic;
        SCANENB         : in     vl_logic;
        SCANIN          : in     vl_logic;
        SCANMODEB       : in     vl_logic;
        SELCALORSTG1    : in     vl_logic;
        STG1INCDEC      : in     vl_logic;
        STG1LOAD        : in     vl_logic;
        STG1READ        : in     vl_logic;
        STG1REGL        : in     vl_logic_vector(8 downto 0);
        SYNCIN          : in     vl_logic;
        SYSCLK          : in     vl_logic;
        TESTIN          : in     vl_logic_vector(13 downto 0);
        GSR             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of REFCLK_PERIOD : constant is 2;
end SIP_PHASER_IN;
