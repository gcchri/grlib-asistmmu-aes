`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iKJl8OWAhQvJ5OS9IAP6WMPqmqUoCrg1uawRRvFc6LOFagfvg+Sp4lV/+nY5h8u4
SxQ95sSmxjMlhF3iMYkysfeL0Ycghg0z09WM9Fzve9rrXkMxY2e3ywW13vDE6Lfy
HtgsZ5BFExQ1J53DUVPTOW+oc5uLUrd7ksCpM+avSIsCqJGxJGF5vIY44LZCTu3c
Ziglgy1fiAluu62vSvBby3QIuOVise7V5J25WCFW8LeBf6w/+DVS4SxlNqe6iS67
Y57ugBmrkzQRAma6ThCMtF7KH1eyvyYBzABQPYDHHhQ8J1AuCTEu114nYVZ4L1I+
sqeYIIC0w0Msp5dVIUxLJ/Sny1lcXTNSFeKJjTWtAO0Qe+7Z6peyPL47SB+Cn5ya
B0+CPRB0O8aITt1FW6q9EnaHShLO2zTPHYBhtaOyEkkUSFLbQX3oZGTALatVA9aj
g+DYxsOydX1XDaCw8J+ZEagvhqlyOHfpsyKyqw3qFxepVeR+PTMaRWtNSjgYOuLE
hprnD8CxqnhI2/uQKxe+TojjNLBWN5JvSm7Qg3mQOqGuqbA+bQmzk76vVo+w7aSo
VwSx++KXCzN6ox9aCIWtd87CfZYSDOl+20uu/V4K/usmyAmUJQnFR1hER8r/Wbqk
Ee/C5SnUTdXKDmIyci8Tdg==
`protect END_PROTECTED
