`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fbyfmYJ0aSiTaRIH2l8lLbggiy49djG6TxZyoA3sWVbA3fSilNOrfCgGmkqQQoHA
+TmafrUq7wedvYGakOpoYLn6avLxzqXSMRCe2sfhcNNA3MzC6xIhOTAsZSmrt4gy
GmihPGjCC1LcxAUqPTOWTP1MFgzOIyhXND1mlnWI3RzFXhe4aFoLM5I94ZO12kfQ
RgINHqEoHxAaA4HZF1RPonR7ydFnCxLyV3kJBQXPwQ/57SrPYgBsAwIlTnBeCrzW
gIeCalA0GQLteht5LIB7YQDn3xRTom/Li3AA7RQsQ7bvPdhDafbfVMnrUxJLLNpd
0SS6Z8XoInb/ntz87bjLem6TIuNY5P/eq8GVC/qMVTmMW6X/RRnltui/kO0KMDom
WDsUQf7QaHBsmM/sxirAiTt2p/RIPvOmZ2cn74salLccRkMuwu1xDcXyVDsvz703
SLSj03/emYFvthFw/JvT7vkB1ljLDM4tTRcW+M4/BANXKIzudZZrUjMGK1dKMPeq
l0YMitqhjhDa5w3ZB5FhckvKCACk+/kjbCFCtlOXA4U5gdVznpnzLZ23TynXQ1kk
wu84cKAnHfPTcIIOGI9O150ePhainx1Y0dyf217tFSN2gWrJEQiZV9pb1fNZSdsn
hF8vq95yhRg+VwhWJqwW2A==
`protect END_PROTECTED
