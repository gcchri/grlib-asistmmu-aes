`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5kRTNR8IG8pb8z5iz4PFBSxPXPXJ8UnhJwGuPoP1TTKh6RgI2/VZK/CF+4sx65fx
IYwVYgjrmfSgG47dygjz4nLYLJt+qkesZAlCgxBxCkaX3ljwsh2k6SQ91NSws+r9
azqag0cxaBRwv6Ys4JDHRkrrf5zBQ9abuuN6+pdSU3JXyp6cVkDZ0VIgWL2tvZQ+
nmotpjddr5GYgmGI8H3CZy3VneOIU6O83LF00ZTtpoahqWBz20ELCgbFKZqLa+ps
3UcCyIoZbQcSdTPfQchTO1MQrfi64gdFxL8se0mw/zoTLTFknnAXelnmceclCDsT
ylmnG4rAPCOFUa/ERLtThr4uo7++98rUA6ur0swuYjWN0szKLAU+UnHsQCSpeEOc
UHjQi8578mVCXElJujYgBPtJ4FQF2UizEJ2s4UuwhfmFNrf0mtU/STFXOtqDLkHj
v/VbfIhiftD5viEa8lLlmmOEpvlMmdeDGrqwwB+SXXEkdCRX9NlFhKbGcvmVTQGs
tW0+feovb3eeELGNQfb7V4Xq+g19Po7HsBAG45CTkavHvnY3N9oKIHoAkKEECiXn
+y1ryI33xWgBNSDp/3uOEH2/zTOHvACfBVHkkUYXZANEyldnw4f56W428sdTigXu
99nNErqRoHdMrE0yrzYgtQ13apH+9Rqu8jj9L3MBpR1V7DE4S0EHSpg/AB6KKr4b
XqfTYV3OJrgUq9LGRppukSo1WD/Rfek73XRhEwVGzGFCSacLqaeu8vgJhgcYBIjM
gHqXcQKcQl+aIAdnPfj2XzfNvprIQO5xQ8Yel0/JZeL7gvaGDAa4QJPkfs4O+I+N
zUUv/JYDuidz24+4aVLk4qXT0Noo5UKb8EjDcw4wYpvFUZTh8pdfIQl3mt2nsuw5
v+V8TzBWZPWoGEkyh2ujKBNQ1vpZ/Cn+PFaHOendhIdpWHtb9X7+7cssvGWVwqxA
fzbRiggdWglVqN40NtPSl/HgAa8k58oT1tw6x2gnsykfJwP7KU/0u6YkVEae0tqF
3ep5NyrBVudyNKJlm90ScP3uZAlgLqnK8mpNwSMmaMSEJP/g1gC0VZx2qtxo569Y
/kDM5PTeKO6zg+I6GStFHpgL152Ow/xSK5Pfd+I3CRN+awoqGmNxHsA+UiXRGrtl
pK4UAUeI7EqOeD+5C0cJzWb6nM9rVk7P7e1UYrJ9iHQ8ZaLgoVnmMQPv7kq5BkNa
JW3JtX/4bnxv0JFl0hwH9tcmnVkjYHYOn1jT1RexYBBYInM6bJUA/2TY15kiGZvt
aLXHbDw7i8oqhV7Jeyr6Vv3hyts3pe7XHKdsI/FSu5zGfwC/agj3kfV1F37AeOmm
SUSBt1N6WSuBRz3PJo1/Y6gTLTTTLONUp0v9HUXW2D8tDAUJ4z9gXCCQfJZLB/KN
LFeJV4u2LsaLXVxAQuvZOOZgzJzrO5KuuW73lXd3wuW30U5qTnhmpI6Trvb1mf1G
48Pll2sQoBzm8zHQf439wUSvv5cf9D8U9CV1uiKfkGuy/twaGLKNEEyWRFTz6M8I
VPQMf3mlRyA6nGeYPZJrJF149W9Mrspb2C5Q1uTat4zJxr3/D6djxFfe+195OogP
8Ggy5iIlEmqOZ7aMwEl1tVaAeKnrK/xu8seXsa9uTFc8CyjgRZywdxQbZRIpfEdZ
VHyg1ry/jxGzbFY/tGXzJM5z9eSbII+eFOvkT74HcFfnB72iKCXuwwZ41hiMj52B
LY07ksJ7Qm6JG0eRo0UAPZZOeM8Tbpl7eE/moaK5YCgav0A1m1cxHBZMh8d/7ske
pFqchSqso5KSqfR/Aifg43d04HCulxNzwSRSCxZqbeDLOyyKIAbTAvuwsgwTP3f8
cU6IANxO4vztjiMjZAmxx6PkE0TdNDuiNHYRMUI8QDNyfBE1HOcDGL0mkDoOhCli
nPCQmo/fBt6zHwE3/6sj1ZaZwyJQXUewl10KTupRt8BY1Y1h3J91ye1K80HU1bWK
IEjNcYSv/a6riURHgpYWEjTm/9R+kGRamWD8GT/2LpZP5JXzSRpSwdRfpb8o6apd
MbN0kBI18K+3HdDTdkA86bdDkWLDxhluXwx7vIlMw2q8TSEDp2pm6rspwlLS1AHq
U2SxZ/DSChnKJ3VvHBbqFl9QdZQVy5qpWXLy260UvSYEMCvSn4xi/ejuUV1YcwJf
GSD/S/xLabFFIJF9zeMBuD23XrZymYzqTSL6PXedONPuXFqonK3xbu1b4EU3cknL
tNJO3VoBiZMbkSthTlQ2uBwqIt1QcDg3ByOwvNBzCX759D5Kdd5Jpy8S69jAegst
Wmuli56ycli/gdG8EO7tlgwBLLUJqikXFMlo6wJrDoSMhehoEv7JU6jEQhZblPzm
AetlTTFB2jc6lrIkL1ECb21xd8FlujdsPoooBGOs9XKGPDlGiVDzsv4A3YtzJPTn
TNmPSPkB/W8B9gABLZEEOpFT6MICongaIyguQK3wxRRic8wndq8IOCG5NzobHc75
pYCowFv0mH0H2u4BET4URcxMJpEJLuRtBPbLOfWt+VTghzcblTCP7hl12Str/oSk
HLpHs6Qc5IaM97oWV6vcotrD7s8fvj9SEWRGEmhmdYfsFjGAMXrz4kNJSPSKAR4s
dMaBnHsZWMbc5EXQ/1/f0g2ApLyOUG2eAU2NWsefhSkcVDipliUw5SKtfH7YMXin
V+pH2rNsfIQj7xk9lnkfYOcoqTGDRGhGNreHmsxdQ2gQIT7tj+uuloDytKVYDPPr
myYdok+Uesg2gPPUQggxnttcvPBhmEaTlMbuS3+LbQmH8DDFJQzUZthetz4wkmwJ
u65pj9MaxRMp6D49VMYcauXRLu5WNfgrsYgiM/5OkB2Ho3tfNJRArtAGGdqV1Wt8
uOegQEhigYejDjmN6gINhE/0SQYng0Mg0J6SULoWqq45eh7tKIEnfs3kYmTlbKeq
puVvIgoWFowSLFkojr2lqkokC7JTvyGy6X8hf895k5fr/7XOBmxAMCq9crEJqWYr
TrlgegtOr2pfP4h20q7zcpvn7G+hd9nNMMFW7wVEPkAPemWC9of8W3dm3HS8v2zm
ebGueIeVeGIY391czDK9BqJHMGzLkz8rMqE25HXHaNR2ilWnzGuHxAHWx2MC7Vh1
1xpVlfv2awxFIdlYl/JRPKbMkKbdJw5aAesr037qMUAd3arD1Q/gGV9cXgtyj1OK
99XlTjLhFSH1d54x4YQa/FRkxrvyUaPf7eocFNdGeb6uMaw/haD++vzRdiih1eU1
wEqkxcRkVZLX2+fEVeD7pZK4VkSzOKEvH8rO59/qNnLexLQGPuMvz3bAMSeFtLqC
`protect END_PROTECTED
