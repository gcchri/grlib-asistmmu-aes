`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VYXJyaVzoxPr43X8vapDEZ4jHdWvVAESxV2MNaTlsls+nn6WBIrE3d5Wde0F9xVd
pAUPClGmidtoYmQSDzuPRdF3RVY+BMs3BO3gc544PBMmboU+eNOs5jUc+DKYwh0P
FyyQaY7qjOue/hmQ/MFg4uOHNQ5+VoQYAhHZtCwaWEsDLzmHlvCrPTdIHzLpddUH
UAzfyTulU8qRzTGf54rKXLFK32nMa3RC93/S18Sk9VTPLA6dGoC59EQaQnfke/oM
HImPnfPcIrA4ZSfBAR/W6BDqsuoSxM+XgjQzqPUYYN2H4Y18K1GO53tCVwb5NqOC
oqD3wCEChtK5FmnP2XIbq7lyl67tobqwBf6gUXujC8WA3LXwlUBz7Sh9awvrtwab
WAouyqLDK1a8jnf/90B6WA==
`protect END_PROTECTED
