`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOoW4lkTQub7Ej0Kav6jzrjSnbIHm12v+6A0tBrgame0yNlA1uuUdNziwNc/66EZ
QpL7eYBkQA6RpQG0ew+L3yTmEnKNESnz18r/mtjB5nDTuUs8Tu2AlnNxhp/nR6LI
gubAZWIhI15BabZsjGXvzGLq+5JHoou5uWQe/KIJFcCF1EzqD2Ob0znETr5Fq3aj
hEKjxfXKswOEHkdYjCr/aFqv8AGnFBmG1aqcKH3elLCoxDiDvL6pnC0XzXJRGgfm
fe0wuODY3NFYMBvXQB/NYcKilwfwT/5swfJEwa7pSFzneJ/fPZWDhILLCXORQqp5
tfR+ewroY+Sbr65JCVd4bqz8ZFc5YSjSzxfeREucs7qtH9UklQuv7BtphxNzzJZY
4slT0gNS4fcxcxV/T3DwojsHacanzqLviDz484NQzhxCWd+uFQnEVArBV9lNin2f
5ytACcimnHyRxAFiRv3AkpLce8DeEaZq3EyFnlpY1Fe11dbZfWkwI4txscbIdqgm
APFQUaGB3hF71LD8Plfl0C890/u2IRwc4e8DeeRlnmjHGEKLAAuSGZ+DAV9VfsH1
THnxnL0cs5+TQq8GDfFL79RNxPGzUXipilcvb8LczKalZhwIQyXSEYrtvqJ/LobA
1Fny7nhgd3AtVrTpf3FcAmX/KcdkCyFusb4n5Z2YVkDTWnnpV7V66mKwcOxAuo9+
DR9l8l7i401/5inkcf35smjeUWapiZj4qd5SkjOo/qFiGMfxPZ2fVVQlVtxe6bIa
scA+Umk3VG+ucBaGN7hIglNK1Ucg0RB+dN0DdaKtFilf8n0YEaYggnN8guwkQNDp
5cfoq/Ofvu9g9rNgozrsYv9i8lDmbDWvzHkVMyHwFw2ZAKsVOiARJ9+wO0QG9LJw
awKcdFYzfwTPdq1mFq76kOdCnFmb1+r91PX5VRB/qGw8A+F0YOAd+WGDu4p380j1
U1JanLlIZPk/aP4aq5OGYiOoD68r7z9eX1CjLBTIJ9Z3UxjC8DwG+9Eq2cGpGsPe
ecf2cVwALF0MbVMooFNPdiAunsJKOxqhk/uVvS0c2wJiV//4HBtpBdzuKeudbYjB
yW34+piwpv3xU+SvQanieqE3Ue0B5IM7UXS+DPqk/7JUzO6/6m60gi/BkmMpyA2E
IT3gK+JOuwoBZ0wEqOriGIDAwVwsFFFTj2BJ41bdIO5m9iWzW6lvcCfn/rMLWOzk
N9+m5yNLhs3lqUAiLTll9ub9VKHMgHHSLdjJZ7KhBtWssgCVt+tS/2Hgi87TxVU+
6Z8AX5ZAQI0X5Xq1T2dmb7/9AmyzXeDSciTBVXOXhnUxQnCEnuQ+tLf97yAjO2on
kKZpxrlZd6eISvCiov2hRgsluQqDldF1yrfmBn5WSTU9a3dFNa4JHKasLCocuTz2
s3jkbU7E2LtUmsASLE5M/kSpp+FV2u78RzRlUyNhzk44LkCS9HMbAQ3dHuSkzJtq
KCWBXZvUSBY1dSdSajycAUxE+KDhs8ejW09e89sVJOwPOs5ea9/n9VsNmcvzHVWL
ZzYHDL/vnumPjr0U0j4GR35ITFemY6HlPZuHarjyGUY72q2lffeZU6RDXmsCXz+h
Hs+oKC1J6KtRKN6JjEOZ/TBo3+S2s2BlTCPrEmF/IHZFbQ/Kuks83X2I0K+I2AnZ
s2ksC8y3SJrN9da7I83Iy6Vv3YQe9UzJQsjsL2YTlfrXsY3yzpMJvqyRomcbZQ1D
OXO1/UWxD9nWacUe/kybvYra74L/XnzgP/OdWT5V0eWynyKRR0jxF9PQdR8PztKK
/x3ZhHWREyqTn2XfWwzt6Ajgn/nrLmX5QVvXbjpKDtO70bth1c7ZUpnl+lnC8QnV
Y8F/9XZcjwCyaFRWVcPBmKL3nyxruT8ZobnJUGU9nxZFd3CE6mt2T9l/ARf9iHqd
F9zlsOCts/26VnUKAedpvyx7pQ20Wagr1KEY9nIObt+C/9zwqFEeHzOkXquZeGnc
WsJuqvUMwsFHUBzI6QZpebULHKeD31ZlNev5N2sPTXADRa1EdTWS2DCOMrm2xfk7
8/hoCYWUcloRMgW5cNnBJINyh5nOgF7fFqLrvDYN+kPx6rh533mnwBIYq6TIX8Zx
0H5/UBZGHsOJrVlPLO6WgA2NPgIpiMgmSW8wYH1UeFzqmU2s8Bfi2g2Pm+P/38sD
UJsiHSoATEqP6JVJIIvabwXglQ3gK1IJuiopOnR9rYPczaHK86ptoG5Thc8PIyd7
ZFeglDnVbYOZvuFGKbtjuCJrJiBOF0mkKNEg0jajMddP40gi2u0UYHispQrLt99N
HgWDZSgOMOqrDhkfyhMaPV6s7SvWOEtRwavCOd7qK1Dp9O81OYoHaT56e9X/Kk2Z
1O7P1+g2zyTKGx8QNIm7Dfgej7n2+F43vGcd2WIPytVxvdpX3YI5qHDzosqjMuJU
mW1MLtmVKtIHQzoC9Z/xMA/zOs30Bnkb2seFAmDFtZF5H8lsj/fFrttNfnhBfsll
oYQUJDhAI+/WzCqQFfTIKkQE/ZNqWNXW9a/0Kf23ZFWjhA+QOmSTQsj5iMLSQR30
xE/V7nqPBFFad5bUjPonU/IyK9EoyvGB12c7v3qnvZ1wz8wOU98c5uO1efHW11PA
AYkWfNzHGTk4aRFj+71vpE6B8dp5mDqOoiqZC/Jx7iYudx7/7fPn+6Lq7vfS6Djl
KQmFXW4da7NyHsUpMw92h8mg28hVitwXbZ65ssy/h0SR2fPQNUBLsyeITUcKit8C
c5VSGM+054JBBveSSj3OsTiFl/mu4m6TXPin2O7xRO/wII6wb1cEefPeRlQjOoE/
tKaaIP/MZgoiYnLu8ARUohCR/uKMqJMLzs5ADEEWeh27mlvV9aU8x1u16MECY6zq
LsmXUMTZrO7Ywmkn/tDo4XdNW5kr4L15XSB2C/Kl3JDsDAjoAcJnYhjNVwwKaYjG
uYYbGlIuyX77zeLfu+TsX0s9hyr0cjojQBns/3TH/RujMPbKLBlkQ4dXXnj4pMMI
Ziba7qLv9FYxJEUB5QHlBlNWR6V8FowymFJz3teRH/IDmwUUMYSqAhJ028UuYWak
tCHVZFVsM0f50C2oD/4YZpKsFPL12hEU/6aQroY2HTtBtFlBck8tXUC9Ci6VIyk0
8ukHIFU5SIcmjRKbUrJcT201J9XwSMg5I6wD8EYUiSxUYAXbibMiuE+P/In5DQWO
AbsfqLgY8le2GlheuUH71wxvE/Xvwj9ZLFv67q0hn1IM7xxFunmpVYycU2aABBGx
siG2kV5ZbL018UwQzPFHG7KGVCZg2gmKLlLcUU2tiosSovqCYGeX5liMI7+TDoiQ
p8pSveihK44YkWbhHlJsW43aw44A3ranjKLhSPe9h3nSPVCB+RHLVsFLkDhp5CA5
8SmbA/f0NhizRftA3TATeDg4g56sTx2NNuYINV6dJjjhT1JfVQgjmOU55Nr8aO6t
q3/I97st+9lfaa3lTkdToD4sJr7u41ipI30+tS09iqNkCOmPYPUrqcoPgyCma5w2
voD1pdirLplw+UskiZheFITPbMXvSVVOSFxMtt/PkqHBt2GiNWhztnf39Xfe0UW/
MZZ7TNTzT1xmNEeciXUBmxdnqd+FTdbdkfJT4UMPAJ5MLnKcXVPB33I5nSiVT0hX
ziyrRrNWnWuhX4N6GuyT6l3xQm5GeBgH2OF9ldIbwpHRFB3AejmhyeonBHOKrtKh
PgsrrCJqOQpvMR4O+gkh53kzNPegN+FkjNMeV+8j2LVyFEBpKrHjrTej/bOA3nX9
z2Plbm2zUDIduTCEN9yYDt3oB9p83b8pNrMYlooEZb7Th6w/8H5KjUfJLzWV8ASo
inmkbUqexY955HgMIDFwGwFUew+bLkEPMcMlOZ9o6hKokSEv+GXLJ1rt5RgltXln
MGRmPk6PjtUbXSNwhJPF6lKAaVrGr8rCQuqtVuY8AGmpOVhjxKGsb0tsf/6+Zbtn
GaiF7SaCAKnTfCSwIXBwR0Y4IXyvPaZ0Lxrd5wOHA5hWwkWI0G6vGydVhuD/VvTH
YXwggWqA+CSur6/DYnSLAHf8//pngW5bKPrJsqQUTuXEKToAH+RLlI3ft/MpkbV8
8KmLtr5SQ8TbIUKKBHTZOn5Th3avLGMgtIaJzadg6lYILFmQp1omVOGfBBXQQ+1A
RM1AZ2j2r4iHEp0wJK45u5NBN7kgrkWhAIdugJdDZntvEBzz4xpB9nyTNQ84SWt9
HCY3Tbw8xuMwsOpv+32l3uTSz7EabqX28e0w2OpMFe+5QSwVHeGhGQcC+C2/YMEb
XXaNuz/G2qIUy70otIU7aggIjda7d7Nal2BHnjYyK9syWDm6TAVFfeOh9j/pQN/4
Ug9e/yHGJqPcxXvo2T53UyNHAratvjO0dSYMhe3GThR+R1xQdaQukhzPMl8DRnA4
N3TsY0JiyCFt81sVXtplnh357mtf00NSnRxdJ1txdcn/8KgUiM0hrOBJmWbEkyKc
sG1UMgKdma3hBaWDb+nxSoDDmjonagTPK+GPp5B2o7jtrFP9yGbHDy9E192qQM70
F+A6FMwWJdJ5ezn6bL3NdZ0ltaqoKA2ysmxeNCP1B0gGglVl2eQwD17vGZkvRwWG
HQS1IKN83GBgDmbdPxDvLcrrrGcC4AFJAy0puw0pugXgq8i5DnhyoegkXVjImH32
kY+TdLggh/IlU0v4QIlgzvqGzSOnbUVNonzwr8i5zqrWPvg6ZBGEmfzFNW1eszlW
L5epWZd0Xr9MjKgTUah9DDweezpWzJUUObIXsfVdVmDgCZellg1RvnWGSnLR3sFF
wcvjow2VLdnFy3TySpfyDOXYHqZhRzI2nKgQ0To/Ig1E7qwgI3Ps26Kgj2lI3llV
FdYhIWGtZ/d+8M+WlFpWHc4C6aQX/lmAhsY1/4+18VSlb5yPyr+q7GZKtV7RLw8r
MK/sTB6dlrlOhFCYObqff2vH/fG5p9X2VezfP9ANVoIGvOjVyQ/4FoXuZ8MOCyle
l5ZO/GTGxR4R7m33r18IeIedmXJEQ1NEz3BjCX0+GIz2fKloA9T2v2n2ccA68Gwm
YO43TyjHvVtFWOoHia6UveqXm0JRl+mJvb8PrSxS55dxXuTAvnFoYJFnPLnSaz4c
llPzaxlauGr/d6NFvBBVSaFfWEjHyHsQr7TIQ6GcjvGNQzU7rWPdIUGr7FlzuDxw
SqUC8OomQdO17wdJdmwtx3CizleeWHwiTu0riNaAH0OFuV550X3UUWVh1aVW2vRK
Hysoh+REcgRZx7wuwL73SURnIokw/yMhcURawzoziD67xq2IqTKT3leeyat7jpDJ
6SsTreUMBlE7Yu9TRpMsW58Sy2ZPuGoZO/ENbkkoTSJRvJmZ+wLeEjKZcDBPTUc6
jSAok4y7UUqStwr0x162GJZh3DVzBPSAW2TKECn2DIODR8uO36zL6Ff0+zEX/tNC
gUmdkfDI6z+sH2qwBGxkzzKc5Dqk9aY5PWTV+LgowW7bEnzAPBbYzVBEMpf2MC07
UVksviGwt8ap0ZxmNZR12ZyCNagIREwKhsbFTf3doGlrkmA/Zk1cxFW7WXC2JQOs
4XSKkUD3JNVEhmjgxh0bL5hKBP9Cn37xKM9SwTmlT4HL9to3swPgWMLbXNxmiZvw
hP5Hl9vQytzx1e5VWxbIUFO68+ZfzlhJGgq49/YsqP1t2vv6IdD7yvdSetrIJOyj
q5BdZuj4ThmUz2G7LpsvwHCbXv3D/EcwwlRaTMyQt8bIRplCM/tvKw28iF5sfD+Y
b3Mj6rxg3AhatQurxxwJE8AYuJ9JR/slZvNQ+uGH2tIF5TqFrJbb1+Dcql3VCe75
a/GItADk8gDagXIFXfAzRH7UF6ZTJfedVPgVkuRaMv2pcMY3a3nJMSp5v9J34Jcw
omiLqRUJT3OJfNkxMdEJLMt9CU9BaCPJ12V5cGWVgXy81ByVaKPYCODJUuvCg/NS
ZDtJPJQvUuJp/AQUGlfoCClA/eqtAQO8HqksbzCY/rutK4kWRY3B0vvuvxnb4KKK
rObPCUUtBBU/LQR15eiFbtBsIk+4bjGSs8ldCvMXqHiknwbRvC7SxpzM5ltPdApc
XLxcddvhQ6jjNvpqV0O+Idka7+aWFk1FxLhFGfgO3KQohlUmT7URLf9uFEWmp8Wk
4p8P7SE0zLTL4roTzLpEZbvcbz2sOFSV/zQQUwuUDoCyQim5YVbIAdPvW4SAhUTI
02P11llSopVJDY1W5Bu2EvvWUN6pVo18TknWNzb8nzNImwUOWCQSNAw5eVx57Uyx
5lcUDBZoRmXp/ZCQqJrd8uj3ob87c8//8QWAbUClu4EXBLbMZAieI0VJRT/r4uNZ
esGtznk69l2/dHdOWn8fCwjlpA8YduB6IFwzvg3arjHITpRG5dCla9u8IExtdwm6
gLruV73bFvRyEB/ViemA9a0L4WlrRYbrALYXC6sB5oa18XDeqyGMpT58ywh2jzuX
Vacpb2N7W6oYUzF9YVfyqDkYgLtBNyfaiQb5HKV7SX5J1A2tqu/hZy9C62f2reP2
l1iaEZdzE2y1w9zhQ+CEGpMZJUA1nAiD1t9HHFZ408Q4PTbtPQ/3VZ05UC4mkcJF
41Ltd7UKmQvdEvTf4ALqnbb5gXMGItRSc4xWvLtqHwWtu12zLbSOn5W8PlnO0WCT
sjnjyJB+2Hx5/Q1pc5GaZnDH+E9LaY5xjcBd5I3gAUGW6o5RCuv3c3XoXmNV+gRE
ukgpJl39gL/8s66fFkrQfPpKuvLN7dEXKVMcNUkxP2s9jYmNYtJ1fDbcZJCZUj/0
e8m4AoescSrrjDO7MTJCjkQoYJfHFa5Ll4mGpF882NcU0H6nMo9A2iBifscP4kOV
94PLLjVJem06jV1EeIv7tFJDwZRNZ0Zp+YvL4Dd0mWXeC3UmnYoSxeHIRq2Mf7zB
674UBnqTJyMpWMjRHxQYYohEHAFdqLZS/BtD1lX/hfumSTzDS0M0rkD4ZA5Yw3ax
J/OeJJsb0fa+idB+wrzmCUZCZBbucNXorP+GTAnKQQK2/UNvxPy1xkPjkbCf59Kh
X7+z+oIds3g6hD/NjZADrBhlEWAAklE7k3iSXJA68TfbMV++xh3qxf3aR71QWI7Z
BYZEzGCUYre3IhnuwqT8m7zull9dMRBGtxYUS9vqgXPr5SyPD8ov59lhsB/EzcDw
D4cyWm2w1ZrcQQKbGv4qKkqEqD3PXnqYJnTSu3anC6HXvrh1Qc5L7t7bY6yWwn9f
KJlnjBplxTV9qcc4OmbheLmB8SuI+y42HFsWsnkbPxL+w1ovefDPlTC2tIQ8m+GZ
dhiHaGyzjesRMnQHt8ZMwRZj1sSLbxI3hHRh7565enxv3Xpxvuu0rn569gd0sij/
dwx/10FKBjdehxkmnrUMqmxWLONBwg3zkod4sg5pM2q6aa5ksH6EeTHA6uG0j2co
sM9FBaruZF4pbRBxTpQGA+7E1StKGOP6S5v2POsEuP+EVUwYL/PGyt0dI31V1gAH
mm7IQDnbkCVx5pu2fmrv95EmpPk4d+z5kwaOUKHq6PknRYEKjMIB67X7VwpQLcs7
X8Fh5IkslUsR+5iZ3S03CTyhhJga7YYO5qjSvECWuN4Cr5Nq+aVxIR9dZ1Rj7juo
bCL6VOdMVIWS55YPFSnkCIyUH5Etp0nsqH/dwCNw5MQszZw1S+wDPNTc6Zn2YLrE
HwQSif/eq8NRdS951Cge5LeLWH5dHQdgTWgTqcy1/L6ueY1Nxap5P3/WUnZW+0/k
lf2tJGCrjVvPtvdA10B7snFGvZu7hXD+Q3rOlhuPHwODkUTOva9o/dfVmnajHalf
ZtP3uwq8cO32mhyrhKAYY6UFNkVi3n5NkBH3KqdxUShpv310cha0XUdpovaGTuS5
vyOEyUt+21aUFv9LskJmViyAbXmQD9vX0sRdHP88CQkewF/85H8MzD2dlNsV1qcv
6uj2MfPgNwXrih/iju+HGTDpGMcooRKkPvQTp5qrDPA64Fvck1Vk36iBWIX137d3
8r/CPVTSRJF/BRF1tFFbvYKm00BiTHeTeIqTxyK3jBjYS+aUzWHL2L5jhOzGVE/p
puNVUTfWlneGQoRkb+XwVCWSVqVC3U4po6FJsLojobLM/JkPsc24yMkDjX7VJnzw
hv+sk4V7ftIJ5xbj8xVp2ymt3DmDZviet6Lg3YMZwWMwX0e3KI9cqolU95JpdP7n
bVSThMbggbgrd+fDWZtCEpyJVsdQNNuRldiWPo7rpcGQtf8Z0ZJ99yPGbOTiZAoz
1pIZCgeTbMKCT/0cDVF4f/dxpF7CuU9zUgzzYmfSfH5fTlQK251R3YfD2/eYSNk8
I0JoNDiPQB4VsJGbvQUIMXXvehR9gxQx4iBoh2+sGuydqMOSf03seJjvCfzbWLVu
z3tHjVLIKf2GXqfcurrMDJfRaRUCocFcPkkYEmS/Yibug28PE60e7lvtoo+uAe5o
rLONpwfQGGDpTrDzNQqovIC5IqucPObUQFSybxvs39iNPQ4fQOjN3RroN67nFJ5S
mYyGUy57E+dJErVrE4vT3OBHo+q6G2NgGrdogBGsvW14Fzko8sGpNLxfQTYlS1CH
M4GLqJ5ja1rZr8uCCHTHmWKsiaMsTFbYYpCQD+XXKH2t6tWeHL+DQBJqQrWQuvpo
PiuFqXvZox49uvimMBMCvEWXFsFdeYkBdVDm+wL1TFz3uGNHiNYUKePq49NZSVIo
5s7sROqhIMSHe0TTyxE9Lj65SKEKkuY3Jm975vS5KdNKzZu4pMl6gWyew47KftYK
vB8eBR+HG5Ds9z0hnyhQ3RYSW5CcUeGJLF9OrE5p3j4iZbH1wR5FeS/k8ZZ5ZgM3
`protect END_PROTECTED
