`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEqKq/cLyN+iRNPYIublxWH0v7AAJUnyEjuuMh4ZuAE5VgOszhoQyDUCwzlqMprJ
faT2FalKvApoZRzG84+qM8Tx5W8GwYBARJT43iyUQG8ULvPyxqPnjn2VdoShfi4J
rGSGsexH2pOBjHCJQWzRlg0QIgfO6qUrY/Na/GTUCYAjJ4SfPRnDSwDTJF3BXsi6
CDPPnbLC7GAJDjzIvXjy/F6DYu6zMpijlIeAGIveedcCucwcg81IamQWj8qw1bC/
ghgmUyE8LGWIa9epzKKzc1VDJNsrME8jDR32FexKGByRFpc++tzhJQjKjDEAP2Eu
Jyf6x3BD/634l9Gv1cF9Mq7fgVutXGku2pX06UCg9uyqZ2uZMyI6ggJb5usW39K2
PJC5MdUV8RR1d2aekCz83hk3r9C55OdJ/aPpv4I3XG4WXO8cfpBavBkO3b9yESsQ
796HSzYx1vplCyfbPu7jJFqzIo7++pB+6rNEvhbqUIgkKgK/6ooI5ePuW93TuKD/
B6jCjpRWgdiw3D9Ef2m70DkCEzo9SgM4/EYHuS0zb+f+2XTDjpNwxXvaAX+poMP4
P8n3bgnhUSUxyqIEMcWsIkuPb2QCyBerSKTfjb2GOQPbFn0Pecey7j1tWe8Esual
ySfdPvqW3IMEIurilWzCGsofmU+vT8iMei4dAy0WePAECXiWZP331YizyZLVf3PR
mQqp6u84nws7um6DXAnwCu2iXa6CvMoCGMpfvPm4AtX8R2FkgeeRrcHQWgd15mne
xXKL+aWyOYRjYO1TZWtyQv7gJMBC/jteZELJ5DwArXI=
`protect END_PROTECTED
