`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SLqs+ENq9KfaS5rUKIocV9WvR04aEWCEKoaUUWgb/vzBndx49X9ehBYfS/BTZBtJ
9sz0aAKEjkU11WBWKAY8JPSOLPhaVtVLVOp/trhr2It6/NdJTVjwtfYBqj/qLAM1
wJzzLsg2q6cUkBeOhJNIwIlIhPRsvDmBatk+DyRi7yeY1KwKTflmEy9YYZyTuJsw
ETzIP8LZvt+w602NtfCqpcF6R7bnpy5nt4tgVLbuYHDh4GAQPbTOuGNZBCKEHbPT
QK3O26VWcJZ0GixH6glRyW0XkCKtnglwVtaLpY7RzNZufTkUunhirBuHYeEN6Gq0
fa9yley6tKEz7lbZhB4hhzaa5jgO2pS+89oLicsePKTO3Pk7hESKU80C55lA4KEL
LiTlQySUrN7Awx1N/lms7KkPMlVapQBFJHS1KHOV0s2Pg1c1Nwd6KV1dSje1gbfo
I+gitilM5Ae5W6FfzirRtqy6602MJCJhU1LHxyupIGtLxFGEmfHEvhh/UJuofI0g
CPTwUPs3lgqYM97DYuCiiQ0+GmnUla0WftZmrgJlTB3setInI59naVJZQ8b/pAfb
E+AZTLZg3s6pwyQ+tf2+s7Sgce3ryBSOYEctMcZaDxOYERAOL6U8EqkCgw/1zI15
9cCvecbHk8/zklAraTndri75NQ/SDW9ALZQV+7BIHdU9UiN9MEA8FCRDhfwVR4Nk
2yz3kCzIz0ZV6/y3doqWTU8vkLMJgYESfLCN6v9tf0XRYfgFfP641XP3S0/ZZh0H
UpSwnSFH6JL0Xn/t0cBWLrjcnKE/DwxeVceRR51v7eMdedzjZARBxZbJmJJQZqUc
IIDkGrb6gFQQDLlHFp5+CLhQAavDU9EoMRpSr3M3a1YWom8Fig5r8CRhXNQuy4Hp
Re86yqWGDu8mYBuIdAsfDYz2dSgfQ31em/W9VvEWBINCbj1wU7sh5AkrJOU6fIZK
V5vWhTv9nlNsX+5UagB0/IJwhAmFQnjT9avMdPGuOHecZH/iWYpQh80cvWmH2l1N
YH/HN1Qd5ZnNONDsrhWVCJ1xL/LD6dxxvsiMsp2H60F7eD750/fd/BuZ54iys0/W
87xsqmRtMUe3uu62scNYQ3jVw6Y1Zi+WvJTJzyFFvFW3R+p44irVuibX+qk9E1gI
P9vUAIYFX1kX718hQy1K49s1SKNqiA8O3mIsQCIzlb9dSaQjodJtLVXXD1/2n4xf
yTc8vK8+9N19Ed/BO/zcjDn6crKjXfKRDc+AHcD8xcD1UV+bFtmtOzltVhT3qFJZ
psHh5nxHBbJFd2ToaeL/QA==
`protect END_PROTECTED
