`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GvJ+ky1NykAHlqaeQbE10ZFVE3y+r+lsAun0HTO9BjaCehhrEN4QQArn/sv5lS4K
NehN+xGqHKRdkTp6lolcANzPBt4xXdpI9W12ejSwKp6//39moT+iZAh2rtJEA6t+
I3jyQanOD+CmfWfQuxD4AaHabeWpE2iP34vWpzzvmpsHUZJfr+3JgR6hw2hWoVCB
6n1rfG4OW8IYjxyqFmAZ3CTl1/d3qZllp0FTxIgHUspuzYnxSZet0HXxj123LBM4
EEJ957uF9o5kSVnJLe65Mg==
`protect END_PROTECTED
