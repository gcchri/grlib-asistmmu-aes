`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+TzsKdll4JfIfTnviNV0kHg+VSj8pRrHjVqSENicJwDIMeAsuHTlBKSU8TaIDu8j
zEES8nMU267lbJ5oZ75aSngJO4JemGFAigTvVSmj5LvbB3R9rP98qQrs+aR+DV0k
AGyag2KHNbJ7UK7/SM+TzYWMP/cugQyfGlNtpV/Rh7hcaH+FyVSyz26Dq2xvTOI+
FrpJsQbGaK8YGgWoLsjn2OA+BeVI277L7zMe0yiYG1Li0T54GrP2s05+lefkTFnC
D4zy2JNE6Ts+HclLIWH5ZMuyQdKqpHcWA3Nm7P3w5lzoXv4Plznq2+fcdvknFDfZ
Cj5X5UtPr9Cg1Q0w+pSxFNdZ/14+QSwa/CC6RRMo6P/2bZdUdK1ecgR+2fGhG8u5
llpUxl6gwxsk219Sb2e9dg==
`protect END_PROTECTED
