`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JGgiVLsyu2JUNypUaW76aAqhkxgejfOe6rNf0ZczmtS8htQA/jIm92Zf1zc4jCFy
o+1upTr83pXiJmrneqFMYRWmdDwDIXhCSZEEuHXyKjoYulf0yc6/Y9M0XiFVthoo
MJL2Fkij/Pr5w1gi/pRY1eBc1LV/02gBoW/4Ed4LIjTM9RGW+FDbf03HACt5jum3
q8okPT7afnMgky57zrJZAhX726zk3v9J4PON7NI49nrKsforytIHs6rYTlcxb9hz
/v+XPjuvfRT3Y3vkZm/RZL4a2FaCPHckrOcnEwqU2TUVk2VV1ZjFfnt/VPCHXAUV
0HwdwFzRHmLVf9U0p9UHjhPB13/OJ2WyjcG11W4q7yxqR71SYtx7W2ZlD009XvWt
2kajkWXUvQcfXE147dD4ytchIMlba/i9XlGQSfzP/7tmrbZpJpUK8UhuhHXo7BpN
2nuPqZ9rIDUAT+xJfelhE5nh8BxoKhJdUbp6mHQAnbHY/lneEqhyG9Csl26A+q0L
QJquwsNgUccena2jZUI1h1R6oqQAtEo0EJJBWsCGJEC4NFzmTX9/lX8ej7aOrHtK
4xYlhP7zpuAEUo8dxAWV2xP6woQDSeTm5rRpQdSvssaoBdHSSs0iIyqgW1yCJXnK
IoQ0I7Hs22GobIZ24383v8qbSHHmASk9+UZ0iFEA3oIShUsiB7+eYwLtrXpYtGQa
u0ZqefjFe7DIl1AFLCqKuXlbNp8SqGAqUI6uWJqhoH/1JSF8ILtjqKdeIhrNidb9
L1IkvUmhYBIcQMaFVnd79rHsK84QZgMhRUc5aYXiO9id39E57OlPFpP5AdoHlRa4
1+LeZHXq3X0sk6Vc57invWPz8Wv9M4uc42JCCa6RQ3EYhryvrlZa2luZ/xMv+XR/
+rEcMbtg6DPGoFhD78WKkrrNJE1rHNbRn709nEH4gVH8tYUcD7xlU2X8hRYehWl2
ELPIUPtyZjSlMQohkqAtK9qohSunyjvvb91ViSivxG0XxVJdKpkM/Wc2daS1yrHB
`protect END_PROTECTED
