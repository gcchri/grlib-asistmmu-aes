`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
34yKoixl+pmdbc0qQ3Pp3gHXbEIw4axhZo+byPbiOHv2TRITsjtci28A81zdPi37
PKhUF7SpS8BAfiXkvNoPZG4WNB2UPOkDdrqCHt417/Vjd7zEh6oiEsMydFcSFpfm
Z6+zqCa4/4agFJrcRQZas+BU0b7WbAc/gXsukOvV3RSWeB45951r4+Q3eOAJnSyl
e9tLcy2jPBUekjixT51jMkwMLn5MDdpsgpGw5sajgKx2H9G+ZUAVKZyJ2XCqWB7v
zItDASRnT+GFgm+nyCGKpo/IUm0Z723rwLy54AkEVRmWvlitAVuC6iCKXRiY6ONH
0GjgLc2UrKiiHZz/ZoLiarkl7iKAuD9EfWallFEJDQqPmv5ZL5Qyn3uNf7rgveqk
RS89diduCwVvL0S5ukx3GqFiQHwtrQBQG+0NpE5ONkeAvPBdnHR+WYA5i6GK3DhL
ricq+FnXOp5bT86qSnUaSIVDi2KnWZ/zRkbGqnEE1MsGu9b72t9hAMIVVhjy9NKo
Re6bz9GjsmLrhJlhkV68ij1yPQULqcdXtcV9fPqzaLtbgmWZljbdTk1Cen0tLTUt
hqzAHjmJLqW2nSi4RdmXvR7uKfdxmk4M9CBrLKp9bz813HI2lGRhEFcN9oo10vvE
638RmywycfiRP+XjXO0YY/podArXTGBG8CmnfvVaS/g7xPEREeB/oguGLqWi7mWm
kYZOlPCgHahPzOPo3pvxyeVJETi/OrdLd4tu3ar29YlYiKzun+92IWDTaiN0c6hT
7hvu7AyzY/6LvJ5SAlSomhrThYs23InccPQmCJQZ4497AK4ZX22o5Wh/820QRtS6
vEd7rJMxWAO3ImjsCbX2pSfr40olXKRwzmpY3jEEUAtuKgf37wECMH16spvt5uRg
3EeUvwTqjG3AXB/aFy/YQCaNAk/9N7zS32U6NRwGyXuAsvoyorOPZAlcUxyRwVj5
vyCVjwPRW7PH1Go1vJBKZM9g4nNmjlfw3LA0JWQqYlnWQ2/YwZjU3EL4iCN56yZQ
8UEF5yrxsKzMMwKUiS0V+iN3Z2JF8mIDM3pY3Sy+0uuU9fqIPIaw9/6OUIf29CbW
6vIm+7rYnTY7VOcwy8RGs5bk6wd6pvLbEJ3M7KCs6lIrlVygNg0oufMGBK9exJ4w
0mglRRyY+639o1znspYszX43dfDdx2UtlUXN8rbkFOGVDMY02BZ8v1zGReqsdHQJ
Dbcz/YuAIVprv0gBD4D1Vho9Z8mQXCPz6avlrZ3w69zN49Tl32Bhguit6MmdrM+N
IXJAO9yG80XUBZ/lUytstPUIAt/OML9IzdvWQ1Pz3hyWW6pSF9aO1CA+0lNTkii9
oSeNjKn/02rmUUO2iljGv4PSAnDgD8LXzeZ1hqTki+tRJJhOd3sTtQl5jTQ0SmD8
5VASszBkjutsArlnObVK0509Q5pL4+BFB/FtU9AU311XkSUSjpuCGu7aDB9ax+EX
H4E1r15SwGfbf9nr/YOyVmq6SRrsbqQqbQI6RLgs2R4vpHeVlDSeNQYVgM6Vmi86
aBNqiR+zzD/g3Dtf+T66fgQbNZArjIJAXePm0Zi321JZsM1zI+DhjYG/Gc8yvSws
5qPuBMBMbz89sq7Pz3qeqGs4+yrBr1fUDT01QElN+8aRzrUe2OXQ3BdaA4K0RAFM
2Jr7ro71GmRmgfIix5csSx2GjHqYMvJWmvmXVwCkcZteJuA4JtghgcUFre2BNxY+
vygRF22Oq8BMz8dkvNqyJcj5Fk5JXjwOqw+zvB7tql8W1C9uXbA78r23Jwr9ZipS
1vaI7GihZ6KP/dFQ8ftYjsXAo8ZkCw4m14qi1e2n39oq7OYm5IvnOqQZZeuBI2Ts
TrbrFajsP8tCk0W16XLxTQ==
`protect END_PROTECTED
