`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjah3fpv2sU37ywFhgshSG5pU0rkvU066Dzf7ej5XyZKHheR0EuUpOVbklF7H4mv
o7AK9EFy8c10+QUDfisCtAXy1AfvXKbIYHSBcCeEDiWrpJTT9xGt7lPuen13ZKSZ
ryQr9jwlP4MX90Kk8ttITsuP4YYOhn6z+RKiDWBQoMXwKnLNKC2hCjRzI50BhAxn
+89s1I3nnerd5eyqyp3JvHUXwq0pXslemcn2rDOowD/MJqfgzMpZ1p626XjVW0It
Q3lTSRlALYI/A0QIQTn/SS4kn9XyTlSSK278z5oJM6SplmaIM+b+HDcJmmS8pA4f
T0AvgTIJCq2KU9qC3VdTuSsHhhEH7A60bieavuxZK1KDAgUAsOOsY41uM1U7IhKf
RyxG/VxqF3+JoOVKf3XMMht9C6atkK00HktEGI1m25CnmQT3wQBULupic9YyZA/m
jo4aypSKlBhC+oTGIYTvoivuTpyxA+5h3SnbQ+ko70mfSpEuAMIWtFHolqmugaNo
ekK43M2Iuzku/kPkmlhqucA+AtBeWBeUSgMCYtt0c1K2+3wwQV+DdJ0OosnQAX7i
IXE/q41hIv0qEM3eeHIvdYIbE/ilUbiE5tRpCEqsP08=
`protect END_PROTECTED
