`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b8CIpf4CfFODTGS9SCfkRz+Kpjx3XG+IN3EKZuScGAHSbRTi/37YAO5nvizZ9b5m
fcynLXIDoZiOqcFq9mveMjThvdLXHYU/5/E5k3mDDn+ik27C0zDmEkcoUIyLjX0V
IjW32aM/MCcAjuHG9bVdpBL9xLTI4sckZlUBlyycgZ1r7h4Lfu20LKm4dyYLRxEQ
ui3M7jE0ykHw79MuH9wsahUzA5mTsLTeax0AN0qgVwGSxtpEqaB6eTYNHcY4wM+0
KpHn1T8LTjJH+NQCHKUj60fKbIqU0qLdQYC6bACPw1froNkIycJ00DEBSVs16rR0
4zZbOsy4TqLzDvknyuV1/TxPQqR4fVgHxpMrBcZ98MT6vYWsAZ/2EW1/h87frgY3
q6xT5CFRZEffTD2/+pqvF8l8d+gklAVIzB+X5p5iKHAvD+jnE5C4eh6BaluohpSG
XDO8ESfyhvtJdAjpcML5c1Qpw2+uujy423ZOTVsVu3g+2wYWMfj/p8cnJOz8EUnT
c15j/mXLDwu3pwzu4qpHTxeGmwcnBJfs7QB9FN8RtuYn2a56JH1cm/K+iZqsnkIN
BDze2TFbMuk78udEUbalxILFwJtWR46X4LN0xsYBuBVvKA82r7jgYsrzhXV4VaF4
vnBQidi4Zr5Taq1tUnAbN3o+jM5OLrmBQXLSjmuV1ktprK+w0h0KHOMhhv0KaHbM
cR7+soR552b45hAnQJzzwYb6gxCWVWjxdzGfnpDQ8sY=
`protect END_PROTECTED
