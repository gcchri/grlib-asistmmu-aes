`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHGcLSE6XWR50MiMsUSr0fWvAr4M844NkxX1eeXWoUtCZJhQv/iDHQrv7sTraEV8
xzQ0cFAG+mlbXf/dLzCAdxhdXYQys4w76MYdcjzr+OK5qRv7UNZcOw4mg/eyOv8c
WWi1gr3T7+aLJyqcMVuAWZG7e813jEsEaNBrDNDyKpJjplx52SDTcCITwZyaztg2
W0JQ6plxEjBJQmsMFR6QuOuq+nbCKzXnpKofG46fLxz5QQBoFmiV7NL6Bj5qHV1C
5eiMeHO4SQa1dJ62W27qZEKukTBZpvmP94VBIQp/NJ4uO8UHyrr+mR0cFXDWKTpI
LNlRea/XPfwSRD+IqTZD5zJvA3CiTjcN16szBCkU95DMrQPo+5DAG02XSMEagu4R
QOc4JGPiLikZ/HakLIBgQ0H601Fi6wlKZc1sdUhw5uuA8L1rFO6Qeaaq4HfyKR13
+GADDjngaDbJpj2Ov6BNKA0Q96OgBEJJwWXZtWV+cp8=
`protect END_PROTECTED
