`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPE6b6Rkl5xJ6H9nV9RVDQX05YK5xHICF2X4LSUjqspV3tywyXruxT0zxZkMkcRH
DkkUAcKBz7cJfUzN2IAhG5KUhw3453EJfAqmqrENtmKjoWST7bpnjAa+/wAGh8t0
rN0H4H96TuD5DI30YyYlJq1TITCfgAuH5Rc9cbbnB5PVMRg6AYi9yFf/PNUc6Q46
Mx8LVxKNd6fQ57epIZI8z37/t1cbSqoekz85B7liWHoKs6/0/Bn3hDn0zFridYiq
ImRHI3nunkRlEmbIaL3u9g==
`protect END_PROTECTED
