`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpa47RkxiYQzh6DaeIHNCQ/fhGP9ro2ObKeCmxznEsDV+2n1Oa5ikC543YqpUGux
3osxXGN66WwYfPxAvGaybYxg9zGDl22ViM4uCpSGgcMWblJ5yCKws9SpYWHsm29D
tgrVMr8flafQwUZZgfLyfsS5eAznUSnIku2QtqJk9jDw27FsjFmqq8DDkAtSltWR
bBHSDMlUeqnPEggA43M1MGJCTEqigrHM756rWBtTzHRLmhW9XewplVjeedpSWPef
dK3xMxjazt0wKMMNX4GSrCnGxedcwhhVasEg+/+Vcv0TL6FM5jTDdkWh/8bRiA+J
AwquXqo4lHNqYT8SQOAlkpdcAHb8OilWh1xlL+9U/coi30Z+d/UW61qukwsQ50X9
AyzM4O040h3iKx+b6s7UNyxyjFPb8nkwORI7HWzqxOygkLs57VuLiLn2y+ZuSwZD
VKOF9PVt7GmH5J7ghOQq6eOQnSH1ViT/O8nIbz1mf2aicMaQ0Qfp8PdL/N79D7cj
PMIQNA6g3QiSIG7sjbpbJ80X8Wnz4kst9IAwDOXEA8JcBYPP1vTSdWvKzlH2AgR1
BEOQ9WUrGlL6bvcXQ6zttKg06wxJ1ID0V41wJuOYWIeiS/ZzTYbp3Af041HbnOxS
C6e4nWSyZo0CR3OaEMvM6yTkPziUoOjlPsvXu1rFxDB5sxkJvai9dOrmxghk2HlB
a0bbmiQP4SUuNFFu8hWhbTOs9M1EJeRLSmZQkWbX8Ku/GCELvyyyMopwS5QKNeAZ
bmhcJIZgR2IL7gWWhtTtn0jGbLrCiakL+H9WB3a7rgnPnTpN252Lqi2XNrX/tNZF
wNdyvREEzbv2cbjkdF6/p+Z/YmZe6w4yWKFMqYKrHo9LCw06DdI8kfkXIpCNUROH
53X/Hf94fvZPNQVqRCLncr5t3qSeBrw7Y4CcbS/oSihX3rylSOFGItE/+UoguAKK
bzQuYlHEbITNExpcEL45flCcfQl2GjK3Myo8lpXsW+YA8UYEEz0vXLg+NzIdA6ML
T+0NNzDSRs5mcKWlcFHJSUyUDQmGhQX/E/0HaBJYlCaN06aR3/TgjkMvTYvTCpIg
prjVt5GnN9L+HvX6l4bDWgcQWTDNaan5Gqg9WnwE78JtFdqABFuHetNi9h5ibVAE
oFkJ86NxNFDoqbwAouh2wpmMBFJrZ5woP6wfUv8YbS7CaDpH8Jdhb0UgdAAIwD7O
Zxc4lvP+0uqxfr396+wbOj6PToxu/pSUL4mMXVGjkWDO//p2iHPXqr5Zst7iYuVA
f0JYlIZ2dQt0JtLzIXq2DJoDbo5xGcb/6vrzJKog+FKbxh08HjIr/QhOg+S10I/4
tfrhKnvzPMiYj3CcXEkMMvMCkexpCVtS8bokVU4R3CGYQRx26H+PiukXIacl3w7a
8haCNpQaJRjqTtq6ys0tOOHEHh4zP0R2+cSz6iQesCvrU9j3xn6t0Q3HmJl05nhK
SLGEXbDhDpPlNU4MTbMwT7UhcbndqS9zbdX/i7EnKwGYd3XoAIenaX17PX7OS4XO
lTnM9PtMhhKRRYMYxC/t3kSDnt7wvEwyfyxzaHEmKMybVAfm4jV/NFCSbtwjN3U7
0ELJ0hx2PI56aXOvl8tq4x+TBR3w1XD60372UneuGpwaySKFShZOwnRYvdYc8IMj
px2VTos60M3Sezf6xwo740qCuBXsBqai5z0j+ZZHIgGkrigGd98gaZzyRlCYUIxx
/nvC8qDPCOFiHUvgqkdzFC0bo3eg4N1eEqdVAORjYor1GZ2K3A/6YfSS2rz5au0a
WMUrVGyD5TuS7CSO5gF+dj4P3NpgbMP0MJeO8pvJ6UX3jGU17Uhp+XIu7+ryPy2j
`protect END_PROTECTED
