`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TxbOaAu5Bz4+M081aXvvYuA20XbQZe6t78q+BU7y9BWEnUEFWt0AHR9DQMTLWRJw
p8F5d681VW0cTz/j6qnvuayzehueiGr+BdzT3WRV9RvHVb7zktFed25S7KmTxM0X
l1vcHa/FwZWlvJ/BiAMmhZmbAMiAPToyjBe298SDR2X2qfhvWty9906jZehIArDW
qCLWmcF9xnJxyvZJ3IeskcBRtGddyhCCBz7PugR1sCJMnz7U31iord15BoPDokhP
SlAhaPs9tW0sfyaX+ZM5gEAVOb2inttw8zeV6oI80k1xuJL+rRNwsDoujU6rqtwx
GBqVxABZmfZhEPi7D7vbclseZGPoTiaUcuFCMUktzO19ULM9rap7TOMzWld9ehYw
Q9vxvHNVpzgbk+KdtDZm2qHmEUNsMaYfZpULvrSFHJEgbhSOykkdv5kab9mZCbpG
DlwT1JieBLd497vdUE8yMEr2frGmSjCIPOJWQSGLijUcjlb5WIEUVJPfw+CYgmAS
1Lfe+S1qpVqPRTRJuLZu7gWiEKHrWORMGeteCCMXpBe9Fd5fm8OSc6Cy82U2nmpn
DGtP5a7PWMXdNAtVzUcxbnu4mpviEbEM3QPbELW+9F+/O1vplvKWA4Funm1jDZFL
9D2ofVHoiDqasB185fg5UI/Lta9J/XnYi5No+xUaUcGOxo3jiBqXI04UGDx1jWMq
SVuBvoc0ILHAM5DBM3zIfgbR71KtQA2Tck0pFk6BpBDYQ/hh19QA71/K/HcR+Tac
OhBtkPpksXnMB2N10SacP/HXS2eRAgdjMEd/jm+tAOr6YT0aJZb/P/jKbufazExS
2wRsK0C52K+sA4cNWT+a1ameKc/kSiaeXqu13FQud0KhxGibuVijcLcbvWhgFjUG
0csiqYeM50mgvBquOKRTD1gMg+3CX29yeoqeqJrRmdD33gFalFkj9I3mpNwjA5/k
JGuhFe5ZNaVyk3G/o8IQiKP68Mw33CZODAJUSiQ3Ec2X0wYouMHiPKL4LeY7/7rb
P3qQkBHF5RxOy7xAICLLJ6hFWx+bSOStXwjG/hM8gawMY2jN6SeQ3QVzDXcsx4wr
AGNeEryUI3ekEGs4O8yrNjGS8i5j7LwXiLLit6RbU8JzUcOuyrlOvQbLF18RZF35
BdSnyQ3vWGLzU9v+dwbgLTRzcqszNgmVto6oInEcjGcoKfeU/MQgv6YEq3o031KI
mq7P95XFpE0iPl0PJpNjE6Jey8phBFMv9fEDzgRexBwLEDmX892scGD2bq6r1o9w
vSF9YvruK1BpkWYC98p59Tg9FeLTtKMTJt/Z/pAlnzaefNE8BtRxbtWfpvQ54XYf
bbdh8zHBxIkPdnb5ZNEMVef/Pa6+jtsenONM0BitdmvqHfGZheCBz9jfIEjTEbKo
5LtJ3dRaCGUcCDc7+f6zE/cJykdqUJL7T2Ra8X1nBWtA91pfuMUE89k91ZJhS8a5
ZuOd5Vlao0BPPA934e3l+/c9VSozNGljmWqtJHI6bnSD17aFGJ/Ck/Qb8wbN3hRR
lbAemKZaqBU9f/XEZk7x08R58ZAxBK1cHixKCc/lREhIDl9d+GNpyJ8sL6hfY637
f3LLjNmhWo2/l4PsYrAi/SyKEE4vGFvDGV75Y5Aypa8JtZNSobNzjdEqGD5WGPrJ
OUNR2nySmdaz3ZdVAw10IuFlrbd4glUyXI6okmc1A0QaZwLQts9NsTMDC2jHlX5E
vOgQA/QjH/JuwZsNeXS+yOCB1cDWE38oDZ7YBflJn70HNtsHAuFOZW2leA4mJ//p
wmJX1YyNyZE+aXqAfZHT/iwIpPtLI3MZTXaHoQciQo0iccqowegKszOIa3/2odhY
wilklmgYpwlBRafgY91l6pJiF41P+uXZqKgR8yUdgtWktPPMyWM8OrgRBlMlG8EH
RgUqrH8itCvtBCVE53BvZ0bUKeVTx7QKogwREK5dx1fSiH7GnLsQwJKKLgRUptzG
MGb+xMftnu2n8CclP7uaXSic1E7Pff1+Q1aXRs3LPOehytYQf2NZiAj+uIj8yDYL
okMYsZZ1tbArsMe+PgYzM/4UiYhXGQ0FlpW6UlUF7B5kTHA5mjT1VC6GUfUd/2Hj
yf10SUe4+ecxf7IGugYgVsyI6uJGAMH92PAuZ8FgasYD6g4MYfCF+6COEop65THH
/ncv99pA4KLFzc/fIHnRdPEhIm1m57b/vUODZPsOf2Uy0Mn8uFjRAp9aOmTO4rKc
WNESdNnoy5ro629ufd1LPhAXYSyK/mCABR1YBz92KCUTMmklTtQFYHerJ8sHaPy5
TvHUaIMihqcZ5FfubMPTYdRQTtNl/V2E4etucxobXVaHOf8GKCnykLpyk7GzbtSc
CGyeYJIzM9qnaWxBTzRJ42nQxEat8nTyvMsxITMAQUVr35I/SVFO0Xem4rQfEYB4
xWCb3wh//ZVLt5qXOAbMGvrswnWepW7SrvAJbW5ssYbZgcKwGdZNdI6f0TU5LEor
H4qaJaLH2j9A2SIrrwJnnXu/cXe7lHTEbuUigb4o0muWAA6enQknQPT6nd046qdL
qwYD3LJEstadzfQ8gcdWjcXRhTZjKmiWjg+cxEB8J6WHmgtChNApCXJLox5sxO2s
sYbwQfr5hUMexMpPQCykUsKVl6dC/WuO5vBcuNG5U2DGLqVbmeGFX2FSfbwtGeqW
CA+shgGzY4ggkD5vcZEtDAN/6f8WqqnYb4AIflyGrZcEVJ111OwHRxIcQA5/MmZt
VnY8nPUYNEnKdZcUnj47Bold6AjCLfnVDh4xok3Ff9QElNZhQkWjOqzn162rZ1d7
hL3Xd8qLwcgICzeoytjyvH8b8AJJEquktyJ9EPF1UBwdq3SFQt/izQM1JvqGn6yR
KDBRsHJREPh42OYgaGQ4ijn9uLCfHx3+OBYswSveUP4yHIRu70ZcVK7NxmFBE6Lb
yQFCbLI6x32b8+tXWDh9MtY5QjakKHExTz4V54JVQFo5N6BjMd/pEIG6TRvbbWjo
nVsCB294si0PZItrI8Hr89APjRmfEqII39KTNFJ11eVzXZPJYDElL0ZRtX5F61mt
0FjwRG6f3A50ogZLuiydNvUUczGGwjYTloDq3YirLQDgGyHlp3MPNp6ymCocemvc
TPS/hLTumensG+9MvwzXwYGMPOmcAo913jhqcE9/+680C7hRntaPSWZuGycT5k8X
eyu1gZIlghHbqaQLP0WvuMaPcT3mxPddbJIssL0ld7UoLl3T/bxfPCvvfORH5Osy
nG6LKbp/PbZbK3d6BLp6zPoOlscbMHKBZQL3M/b4ylAMkH8HJK1tcaGcEfpiOTGe
8jZjpQnJQVVwBGVJC3C2bto4XjQahKyMAl0cfiD44lq0YT+A+jaXmlXg8xZlYsWR
4+Ac4E+M9ItdfFqIBFrLj9FDOIinRzfIQM6Lj9hTZ0cMke5ls8vekASaLyhWuwul
3Whrydn8nn6VcJc+PmU47fGnW3J/2V3S3eZTO2QxhqDDvfrGIdhEfeUUfdCMeqvY
b7O3938rzJ/k9nqjgoFwk17mUgMgOyuqfNXCBcPnlsyEU1uWlBBnI5WhjdqglmDt
GqKte9wus52EslCwVftD3zT0M09XBSWtyi/U5xxCrhgYiz1nIEL87/EJyn6X7AlI
Pw+kbgSINgtuZQ3IWG3VXxL0Jg/oEdRs3V4btfVatlH2JpymLlSWOMZbLkeOGhDr
lHb99+qk1t7aCuHnCv2sgmVuT5llS2kxZiH/+idIqxtY/s53w0Se+khOPlfxUC8k
tpgrzbQ8eZ7atGvA1wit6larzO4EcEPv5MTYkBpHK0LFqv6lk6HAIIec/u8JQv6l
nhppxJt7qQkSCEwLlJBNv+SEEAQwY3XX3zDl9GUS7NuOitDqKx8iYETzk6MSo1Kf
qBDoGkkQE1H15apWkAJBwSKRZJqTg8VVDi0E0LkUSqVsC7XrKQdrbol+ZWpdzg5e
gOHv48Hujn5iCIKvgIaqj0C8XGZCkAnbCzb4kXWk4fTwwjEHrapyBICERrXjDkpE
D7mmDF7D7iArEDdAwhxlDvGAKStYnLo4ocxuBWujrhaSiwED83QXNWd0k7Vcz8mC
Cg2qj1hO9qXT9EX1EbY/Skp4dNXtoVAjhKlmz3Nus8oTprfiZA2uLi11o5mzP77x
PLMppfRTpVjby4ld19oDOA==
`protect END_PROTECTED
