`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cm/iJjLon7KQB65w2H2+1CY6KjSybbUY4zOWL/3K9hCc6SDoqb768G+rjBrrq8Zn
DjKfXLhQPPAstIrdDc14FYWXMGqxGoU/W9HGPDAxHcWDo/nOBUcnk6zWPmXNfJVy
mhU+pPtT6okOCWh5VboyuqgYshqDiql5dQW7kJYICBqx7lIh17gGuTDWdj9ihOHG
8YzMpSLr4MVFgU7F2PIagVYMZtUvu8f7vRgOU0QUGhxpqmDDJpSnirHN2PTKsYrN
v80Jl4CqYnhwWuiVH7lzAlRh+aBtFi6nvAQMJKkoONA6XLCPwdCV4oWebp71C2ht
EaCZT/6mLisSRXkdwgt51uhtDsKN2ZPNo/4mzfB3gY1EZMjTWUStb/tCtdBkw7kj
/FBu2hB1r5UL51FdVqE3XZIyOCvRo0bM2QD1B/Og57eEi2nAd0P2iKP4v44Rqzgg
RVb0MaTRe8X99uVxjrD7sMmR6MmM6JlN/dIUCnXgrRBvzjTMo3+bSNGFFgs6wmk0
fDBC1r4FQz8jWQcG48hsND0ZsLoTJE4W/AuYGFPrsqUIoeRnQsuS4sJimrruMisi
eLv+Vct6QG8TFUkovs4fbA/rYXPQOmF334ccFpFDnugtWar/q7aEAkj/c2jKimRR
E1JULLPE80RDsSWjbzwN/2wPQrVHQNWxYKgsB2DvqA/gl0yG4WvA7NIZJtuCYGkO
Z0fjk+TV5IEQXv5IZ7u1QvY+BBmyJowOLoH3szed4f0EbAOIjEh1leQ7QgiqgNXL
TOj4c719SR3UK2pNsYjSN7RQXSddsbBOHty0vw0niyvW1U7PWMp9Al9rG++6LjEB
1ftEQiWZoSGH9yCkdfyxO1IZm4teX+9l0FNLVKJZ11UWCjk0QVSKA9rJtULsCCJb
41VrLakNlSbngwwVnx1x/Is1d5aQ2VOd9ef0jbppBob+R9fulre9O3hBpzKSyQ24
erkjd0VL8/cZq5CJADVbY6NMjRlzCrzbFyYt6O7W5Eu/3KGpvvJcGpt93IwGi0kq
Hsr+L/ek/ORddlOSheDAUkcc8RjUGIuUb/YaaXDsonN6HEqalbKUPmGfNV+dC/o+
kV3cAW8YaUl/AfHsSt4M4vQeoE7LO/dJH4VQ+2jiu0GuiVeuOTWZ4JxhsY70pM6U
VZQr8tEIgFM1Q2Lekc2Kbo8GAuy3Tooww6uxyH2EGadNgFE3i+eweJPOLaURBDyw
AflL8uvy1mTUQVVH+J/g8bN5npLuczhAEEcUG8LZrkUdIw5GjlgBx6CS0A7MJ6Ls
uq8c1QkGI4ajG1IvL12M6NR1HP7ynuXfc/ZHcbKZn6r6zGxwfa6ZhduTiZyRYmbI
KUeCYXGOoa98CKp5w2w8iLwTsy6LszuZ6nk7UyJPD6mENtU4OMybawEFZ+5SancT
iKobpMManktxs49Sct/3gqaKsodDKxtPFeClWGSMJnRAUKtSOVjUnVBIQG6Rm4Tl
KGF0aD7XrWralZx3FiW9JkNjG27eDYxnc2BCbySbMnZslDpTQN9kXxoHQ7ugz+w3
vLIP50x1SFWWRugQnyAGW7szo9brsIoq2QUeSGAJHMlPb151b/rhe5XGDx8a3CoQ
5bXyWfv+c+qS0gYYg1R97+z2b3xWd6XzVOIOO3LXkvLaGL3sqFz3g0hrRZLQ6h3/
5yTS5GuZQq3iGibwfM5WZr6cxMdMXGHmy9HGmlaovovzl4U07XoUgFutWKk02GLO
ftoIpbCqHilJfKcU1mjkyKBPscgF4SFLt182cW5dPClvMjHqPqihNO9y2Ozo3IOg
iegEFhyL2I4LprnUqJT4BSpEag3XE+/M/npelottKSEwprzepxgDNj43cT41v5CD
XDgINe8jBHA2u/TyhtzYyBxxGq1hJ4ru7PW6uQUW60wKqUUdHzwByk42ceo/W4zU
MnbeXIZzSzP3/R8nVTNbHZdfiubELk9dmXU7L5xrPG1mF31h24v6zoPEu5coTPAt
ZGdiohHCx3wGNTdPKvxmBfUaOigORV5AR5OLJHx2C9CRnYaPLK5C7mU0Wr0ZmYbK
zeN1o2CIYKNoVzhQCEtzi3U2ftMpRw8JD4FbphQnSLn+XT/beX+7Bgn2nCyDI0Xs
LQ+oo6vS6PUCkbVa189CWkEQ5AHxnQ/g5RzzMG90V2vYR8h7ppUhjdvFXpdGJ9sX
Ma6Drtf51SZ4uEt5axzSXpn5RyYQhd+YBvz4wKdv6GfmJLn7LewzBy0sbA1mak36
R+XAG3EzHEdRS6s6WXk3EO7dhPiDGOGNHRYbfU9YjVyr0fjCKBCqvjjBw3qKgBVl
KhYs8j5GvZG0ryo1C5BXJgoTzueXNoObiGptzhH7P+VJ9A6iBlC1Jdh+mrTndOWU
nG3ziYyUM9P519wZSa0IwGyvTDUfvXmSdz/UHl7Gn30yifExr1IoVxd+jVYEH4YF
eQb74WWX9r9/0ppffvkP1k7KhbhE+vMCHQQCp7EDky20BEoaYQ5fYPXSUL1tvD4U
vy0t1paTIZZIzJyXoTFEOesOsz9zLAaeYGIC+a4K2yxWrJDtgCcVOc8nKCJ2OiKF
RPu5sscXfgQQHWAJhCndkWFwLN1ZZpGoE60zfFu/kwHjSQwGakZaMS6VZu8pLZG1
ELCBZ8KLDj9QzYMvqYCHctzqMQi9qZ/ZLwRNYeycpdu6QOrRz6RuV9unp37A6rxR
grpCvFYim24qYeNxwRV5aZmiEPEwkVH3b3+KTzcXa5n55GRMD/B413sMSi1xUY+Q
xEeehVljWf9ygiKWvnmJwZ3b4HrACdiJhJosiftUyncI/hYYDhf163iHlM2U2mPT
yKiXFBh8lYapnc8GPuAJ6EH/jFHx0ZFxRQ35Hcf1S6dTXb8CGHUzYbyyahERhsSo
ysefLjsktAFsGgSYAFkisUxj9fQNoMZKc/HQexaVMfmAECWTXFvp80Smu933p3NV
J9fBMjiNBWfL2YGkiskhnEVT8MRBeC9oGLWRvhG7mgKehazyBqqU/XG9oPUK9eWR
NiQURj8yzBdrskWaNJaqfpMNTnol9Su3Y16Eq+AwzGzQIioTPO7jIZ182unlx4es
/06T/tsvimCjIZhdstm2ZE9+4fZJCH1fQiCZb0zm5R+xv9dE9U9cehAXkvOr57Kf
hdn2hX2FwLAkeqY7leg/xaN46ACPFH0L7aH2qpQFlp3jgzxuh1EJ3swjehI1ymxm
9CkioaMltKOrVnV4eQKle3VKvl4VTLPVdENTPhJiA3Wz8WiPTwwoQi9xXkj06JQf
9qjGFsCa7B+EUbLsugTTL0jx7ZftTsFocNN8578eTd0i5/lwUBowzaA0tntjh7SB
uaOn+UCzWiVYnWV+wD6BCg7QR7GYBeIz6N9g4WwCXELyyQsDHwUFw+Awcto8keQn
GvYcPGMfFYwAQC3UBYhsUl2KLHvowoGCPwREkJMU0fQ/mWx6THiIsZSTCg3kmD4v
txdJ1gYIY1xaMm+NCaZgkW6CypT3iTv+NQG6fYbZXQ89NcNpwOxbO8BSZHPtXOaO
skl1KrkTWZPq3D9Q+T4+ApacQb1Efa5KAXvMNCArOngNhRaOQ+qM4CI067cBM4/7
zN5iW6pCso1FbGBUoeENmy0EpFB3KiA2UeSA5TVusw75poTvA7LronKyWtKvmXpP
7g0k9hIZQVDbR1LKJiWdOPDCSSWqmyX34SrUQUr+yibtXTuUag7IaH5m7AwtMKax
V40yXlGB9YA1QcixH6PLlHE/PwmPYcd3FQRWR9Apjn8MA/RBsyK7ULSamIJklCde
6M5njoHDmbrzzQGsWjuATHOp5jvviU1oRZ2JcYF+YUDCHv7vsyAsj9GdshTQeROt
FpEV8hWIKqYTnrBww1ewvklQ5J1NTMYh8VdKfnlaHNHPXZLE720fD3iGJgMiAA7c
jFKDpmCLwuYheHdmNSTuvlXuYIjzqPK7Dvbe/FC+hNrGVbEEl4/U45v69bRqGjaP
UllRFznGY9wO8SZJAV2cnkgVvJKXYPw7svJJR2MWBv+IQ6xiTiS55LP43Bfjr5Uw
aaPkwVZFcwvT2WMGNjdxqYYPQoci4lgquzLz6WMvVjLW6Fs4ywFNZ2hdmZ8YGLqM
jfExV9lZWqnOqWoSAIsD3jhEKTGeA0hhuhNUD+BE01ZgkOTueA15gXD3BVQCMaWx
EeGaPL84We703gqT6oj2joUUvxyU7KbwP/V7nRr1fuT3Trq6r/z0FHpWOJzPlmLj
RvnLCepJSOadQN688oj3S/M2HPDHA2MRGJhISeb30diXiZs1Ye4WeQ5ewOawOor6
Dg3RVttQJKXGiUOqTpQS945LVHtgFxLmrV+xiTBiFkRSignu4AIWzp8Umg1Rb1aK
Ejhk1b9RULez5ElOjHeo81BQWv/ZbmQks6TsAPXT35rhFb6B2LsswpML3fnYAUMW
o1E5V90xA5MF33fn0NLCzLU67rMFTXn7Mb8zzPMUkUnlRuhPDzO4Ekky1dACivWG
b9eqbq8B9xPhg7SywRxtjRmoK+AxDOmnhwLb7RuuYYUbvbsFEEpQNawyhhUDxD1h
fx8XVB6wYv94t/0eYcWpbHXi3NKXCXuyG50gNHI0UzMvikr4OsZLIhqjEoBzlvnz
HTWsxAVjf+RGw4jPNmQj3TcRd2daWsbG+YFFGgrIkUk39tahhmRcuidhHmNzsqRm
85XtV1toe5Smc1SP21sIf4SitsQ/czIH7aHCiWfhjbRLjhl4nDqyc7zupFsjxNVL
ufOasJcW5m80as0tD1gwEnS7CKfpZVRfuV2FdYi+8OTdAW3zB9WkIKyKBPae2Pz/
CrvowCb3+X+HNf8KnU+j38B7Y3EIu6AshiYj+zcrAQMvQ+psKRiYqC210M1RM91C
L9fsTU+v6fNpx0KEcKxb+ih9+yofVq3aSpem4WtMdTHjn29hPbJavDERKJirUId+
O1R2fOhyYNv2/wyd9MT/iKQQt3Aig79MVRBRS7QaSY9nBFf0ta1XyMzwswP30y9K
OZnR9GN95k2UshcHZdHPhip1mRTu1lvfPQzZg85NHwk+NKol06C7+EmFaiZEhs6X
8Zg3rqnFsuwq1JAsV9soJq/V5wImn8Yb1L7VZU52hCj18cxKZ4XBGZxY9XwHGk60
O9JVV9gTQKvtiQNrVEgZXWOH8ZjvPm2kS/c8z+/P2Bj8AfFoe7CxLDyhSxg6VxFt
MXzebOPqy2csVMse4wF8IuSoO8C6CWjDqGK1KCjj7tHRiSR69gsnsMt9FqEEQjgD
RdK0C3mttcyF8fzuwD7h6U66xE+Qw19rsDA1GetkNTgbQdC62FiSDpbBEhcNahAc
9TwNb0OXN9vYHRNpnGxMw8kablflJQb9/hsgpwXq9uMEeucoP38rULraZ7naD1mR
GfgMCukYJrL4TfCDI5zXfhWUN/D88BeBvNkKG26Xc8iav62hTm7vfibYRrKZTQLX
+oZrxDP5nifSy3E7XHOlgWGncdBru/rtRNnt2KwipPzVMpwEtaQFufeOn1K4ZFps
doVZHRkowfZs/DAv5w5TvmXCFsOxP25d+ONdQQ4ok2af3sOwqLueyX1V1bAb/v9p
G2E483JI6QIHXOa7PJhDMTiKUv4EstsoK1w+o0CuW+ZaVPkK29V9UY61mcM2Nkvi
awwOHii08dcRojMR0qWYNuXtF3srfD+UiA+crv93pAisdMyu6qDqT4KtVBeU2H8A
ccc5yH9GkudkB93tWx6EWVjyS/PRsl69gjGRZwrd9ilQuYD4ClLgWDw/hsPUkZbI
KAvACrODUZ3/b28DArd0GwsuRY8QnUVdS69O7AtamH7REGnEwem7a8jE+GKuO6Zt
6hN83vma05y2YsgY0ATCKPFwGHmFB2Cfn6zjzw0hRvcxK9lC7VyzQA3MJUo0FEWH
DFkYrMA70xMIVo2rlMOrFmdhrrrrMCJ/vtSeETz+zI8V9muxCXpR/0E+C4E74i3k
eFN4meaqlMqifvlGqKIbu1ENbP4tXScIkuTQJskfG2ObKo5+2TgQN1FcSyl8dBPE
3+9QnX+Nr3EdzJHQ2TQ1KgkGJZg4eDrj9yBX07EArGhyXpUhNGLHaakOwgwNgCvq
0kB20xHt6R4V1H5dQKwwuEs7J++OIbOj7DBOtmhOcgxw/z0+fWKboTlRvLCLRLMM
krQZIlM+2iOTgEG4az6sM3+k5k12WxPqq5oz/MPnsHdVHMPLuxw+hIT+KjmzJt39
81BtM0uADQ9zZvfP3Dy/pCwmhVJOcvrvL1Bw176b/URa2vaGSydrqarGx633XXE3
hScg1i6i+wNspknYLfMQ5/C1FVclT2vgGZhCH7srB3K7xdjErFHB3mduQ1eJsdgV
/BQ53C/8pMItuG7ozWy2gal4RDNEH8x6KQPBhciINtO76Pg8CxsH2gyytD5Qo/O0
t5Qj89L5JjbYj2mlJUZoOwxs3I7eCdqHt4hdW7Nsr5TBuSSoC637ic8UEpMxVhsI
lsfRFhZX+dRCkwHjfNFD7bsT0V02CJcNPEM6xsHvqY0oeU6R/XDt8tItAlK9INfg
hv1sZg2s8Wl3GjRWOyuuRxRhWIt38PCTMzgelfC1yPv4HHZAp2JCV0WDwCWsdFEZ
eYcTKsBnhtl1IIYCSFkMf2YxZtt8tG4VIYZiTdS4xMhtZzwoq/u3YmjAWlspk0rR
2Nh5GUHf+CUofo57TZq3DpL504Cifh2726j9zrii1NbXPItOR05Rnf5JPMY7JfUU
POLi+2T80LIE1GbyxtxTqx3F7GoEtgkE3f6HB9YkOcPMNzyeaU30zxD83Ccsi7/5
NphjeXg3L9vuhMdmwsj+3GsTsjjglY38mZgLe9E0NsVJ7ZT6PQc/XJ8y9H4y2hU3
GAYrlfTPjcOTupS/xUzaZPYiowJ0BXciUK3bP8zl7g9sbKrCg4MR6abXaT9vThcC
MYmmlcL6xaK6ARN5xY3tKg8rd+gB7j+3KPKE2RztFm2+G4JDQxb4YW2XpMwIxKxg
eVpSpvtLX47MBK68JKgytMSTM/p1wJlwB1GBrpoHGXhqRU2XB7nQQ3U1Ht4mle8N
DtnIeusfftaslctCk7OtYHWay5ek3clbjhDHYhMyaKjWOJ7xHmI1jm171u0163hR
/EPnDXkeDsc+JtaPZ8aLOWWB0gnmsgruf3jx+yfaQjzt5JqW4+TP/jt5hyNhQVAy
WjMf16+nnX0PTVDBZ6CJpdNdyjVNrTN4Vn1IXXtW6welAu01WJ5axMBrEorOax7t
yZFakPlnt7TFD8kohZlnijmC+3PG80CIno757gKg1myr8kW5Od373/ZIESdt1wny
ghmfPEBIn80rpfFXot4P2D34bNMYhi4c4DQg/mxjZn6x5kv3PQfX2QYp97Ckysy7
EEVrOLuOn05dGVKciCkZTZu3kExkENPkCm7CuJwGrNZ+TCNsH6Fanp+Zt2SKG4jn
s5c3T5nWBOAqElKX2v+3S14ZkSH3sV4y+XGBz4bAKEK/jGiE5T7NtNB2ADoWjXUQ
0JiplmHmf+8GkT5LXYn305+Ug+Qd+Ls0RQ6FYdli3lqFMU0WdI/62Q4UcgJKe3ec
rYAi2lNlpm9cOxtiuVKTmmPbCAJU6TTfBVo+aRYiFoBw+2ld0NlEbIX1cscB+WIn
fGP/WiVisdl869v+jmsUhQ9Vr0va1HdbK5rRytNLvIK3/HIxnFU+6crCGjRQM+wr
f3xo244zJBoE2K/l5t5QdOix0clBVyCLZAC2TvHKA8WmIXb5CtmRaohzsIG/12MR
VZ9HYDPm12uMTh0cXBdk/OrJcXYx5IT8+LlQfMd51gdKtmd56jKGicio4oQo0Nbd
ke9mSoIShw121Q0K9WWo6MP0J6gMpOoW67a8IbFth59vIcq60+J5IauaClmKWd8C
ORbbRXdNWNISEBdP2C9cbSrDw+US9Boh6tdQZ+V5pGvWxwQjjYQGATTJKk29VpxQ
CkJtUX53SWPKI5HBIuXILzj8k+GyRojsj7bTk/tvC5hz+JYnh9+thI1xm2gxOYr4
hXAzKxxprRc8+RjRRRMpmK2W4EMOc4vXJIw+6HKlMlANJYjUrk6sjngX8hGE55oL
3APbwypfsCZIoMpti4yleU4tqhiuXtbjnDPjXN0W0quRJVrnvfdtgTK0J615llD5
zetPZnpGV3NDe9ZXUHJGW8ejuLPZ9JaVdo4b8esssiwPt2RZcMK3XVGqveGCGvCc
7hHejRXhESwriRqZTyjWnB6BJDMsmdEjsTb5nEDkBuTlKxxjfv/ZsCRjrDmlLDab
uxe2xgo9wX1sRPM5scopwG/0L+QiPdU+aqc1SKWbvqlGZ31UA2vYtDsTL9geKqde
Fl2+RoKVMZr95gHp5yx+yZvoK1l+E178AYXvLF8S60N1ERD8xY6aT5JLviCWlTpn
8ho4r9e12OT6lXWuX4izEjw3BwXI6NaAZ9p6i3M21osFSaUPsvXqGufSMo2Y0Cx9
iUm7PD+YhcWSvN6uJikmZL+RHc4gxoQfcCHNiuRifzk+XssmpNijbha9OaegJMZc
1zqlbdPc8KOUd1XwQNhaDV2gQfmrvbkPNCfU0pxUlO8MkBX0Ts9lk5KEHnUBcGtv
9lAH0nTHlAg1+W9SQIEdEGcndY3bp6psqw+UAc8N7LxorEz2ZjKjkAm8+cobzZxD
EpaQimZhFn4sU3xdiPHtIi6uSESJXfcj2Cv4EtOI94TP16E5Petls56k7dqB9v5W
OseVJ0AUuABbznTFUXTP0NztHhyO3tC/ZKZTkQtJNRqkXZm/IQutAhWO4v/ruWtL
bGfADzCUMS4KV/gNpTSbC20XUqoXM//MVYuzBIbf6GsHz++Ws3itwqJ+tp3k738W
Yt+ydO23gqeAE4buZw06ZECuxChni/FQINU9rwGQS4Dz6r/iqa5HGNBKObwj0t0E
1Eti4Kmv3EJECthr1xlYe1f0IIBHGgXppeunOJ00O1p8ddPwds+WmkO2301D6vs6
PyQgF+0NFscfhjNBOx1k9QZJGpLo+d8z4/nqcHFAbE3VN1Wp3HNaFR1LoxAZ/tEj
a/OP5NepsBq3M/z6O6GhuuipYEoTNkeIzwvleooxx5HIxws9lL5c7DGT4eTBZfXy
4ThIvuhCbkgWNhd99m7mo9ibntc9Sa12Vt7t9hwEFRHkonC5rWPh/4kW5jQjl8Vh
LpBakPXAVR9kWM37mtkONR7SkrhnXVhGuuSa7/0UiNqKkUQsOyuA/hH1bzzYJpfe
2nGo9DVjmtLgvxq0ySzDivhaln/sGemrPPchVhhZqpeDPDzL2eryMiDn/0slu6FC
OgaBBXDlYJ2nhCp1CdmQJDh1BV/yYwR8Z4afadnhR5kDgmDCkVbcKeT1AI09VoSO
PJ+z2g+wxxI/9cdEbYJM0DNbi4pNGoo0Jas58J3xbUP18iG2p1hctZzhvO2XR+F4
OMi+6kHhU1LOjYjDR36t7cyhg2tC7csVZR5bM7KvBU6nUf7A0jSum1HJAcidlev6
8T1+ldivb1csZ1unkvPUhFPXQQ0sa32C8Pfx9SkfDqXM0MUoB+qOUgDgKh0X8WTA
oDmb96jp0DfbhNPFdVulwPPW8jg7xUZVIcIuzXni4BPXkKwU+wG+x5GO82bqSRNW
Y93ELXS59hT2Gh1w0vqqZINQKJr/8mKnCFUwivmFpTaCrrKkfhTkzQTGSpQbDoUE
9ARh4mCFOtI3DMOctqCyhTbx2/wmPF3gEVvbXYz1tPZOGpaE4KdHKyAtIYw5g+cq
MZkfcm3twYHMDkEtPCH5H5M/P2Mp3Wk8V6H7aFq08i583cNuWwAjSeN43fGcaJcW
qDolxoPtuKP+EzP20AfVt4z1aEko0miKGtfNvGuHc7jB86AQ2UPtA5+Id0aqDVZt
WIQ92uRVrUFdNz9CM1h3rkbrhOVV6isgHTGf4Ce5wpRvAC0InbDGlvNWQJyWFr6J
Kt9BdKZdEhGR5kJFWi30lGXKuZcGysHEi6xZjNmMQ75mJruD+6dBJfD76sWxsdsy
1UbB5wgKvTZf9Az8N367WwPc+7TO7RPW3TDpyGJuMbgOJaJ4WL/HZNltbUD2DQgG
DVFp6U930v/Qe309NoTNW8urY2yqHo511gaIK7BUSSrUTdKEn0iToMlTYWCFssEh
rtc+WZsbTtMwGGl/JKJv2LtQfqHlevXV0L77VFYbqUE8B1qKYCfWeRX2esl3hszd
LJYH7Z9pIGzELqnScZgma6H4eK/ZIeQDs6iA7HJLg4aTeqyXAyBRvJZChacex1qJ
D0TVzfiaR0eFHMR7uATMNChFlkarVA58y+z8l5e1jAtxa3b+zPEdWz7seVKKIVKu
lhX7kU6l3xtzYtw/Ufyo6wD6KVObM/o0ZvYQvs2n9K43Lss9DzLrkAcRPi/tD1Ht
GzuBplPCCxZzJtzjBdEjEiGMnFMWtk3BidkXW3XLTZNmX7hGt7c3fwf013+jfCtT
IHVSSZzNl2NFvI/7j/RdnA+qrgp3PimWkhfDKW+xAkVtd7AD9RxgzVATGTTBRnWC
OdgsX71DMpNsDPHVAK8uYBBubLOBTykyiOD4Dwib1gHrF7LbSRXe6OyBmX+rgLUn
5UorAEnRKPiI089d1dOx/1PNAVOGmjH9e1D8Wlc5c4oOi236JIrud0ccQ0B+RILJ
LjsP74UetbgeYHjqa9ON4IBqkS1N0mj2c/2qyc3Kx1pzkIREympOlbINLK65bpwW
i21OX5f3HVfzApRZ5XKowRMrHI7WxPPHbAJzi2hOk21ymuzdZBSti9jKv/NnHl2B
My9K/Mo+kVF3/zvll8+Q4Nj4R8gpSUnmIQFduAuI9deI11yyLxtkiZPoZerNugYh
dfHq7zByCFyvl/LgtSMUZSB/xyv0eUHh9EBUkZcFQ/6pQd5e3lRG/UViLtA7MLh3
L79dgD52nu7dPHSD4Pttn6P3eh2X5tjCGgYuKa4IVoM2Tq9WzmqXFER+vI2Bh8i9
xWgyYhVS3kpDdEUFiJA91/eLaBN0249ldJcxD7mnqX0k6URNdv072VweC+7HGi13
vmq3oJGodmWl024Ju/o7kctJiPoiuecGta/hLpq7U1IZQeHMGPGUFGxxrD3uNBGN
g+UKYseoeWoKmCwMzb0SoPd6Y1q25NeDQYm/Q9kOkJvSnVRDzgM8pJqYheS0Lqii
JqKcHr4y3fRi4D72SE37fEdgwBKhTwYhIaieLIxY1Cat2R2YW6BtGFrj3WQfqNXT
eieqFavz4/m4g7oE6QulxSJt/+83qECtdB9jgGBxDCthDh9s8/oNC8uMjRfWv7eO
yFhmXMRvgisfH5V6Z3ESSlqfVZMdjSaK+EeF7O5i7NQXI1clwEmZP7NCu3kymyEk
jUHNqsaZdFHAcqX+ySfru2o6PL1BfCmt92YK58ww1Wjy5xYoMCNzY6kLj/Fg1bUQ
O3VlXAHp3lYKnRv85WJvbx7y4yY29FMqrYG6sSWAY3npEMCJ8GwyY13SNA//X0I5
Boe9wtpYY+DpwtToP9pZ+GDfzOv5z5QqdCv9zKeYLiK92cV/+22MCXvF0hDUYtGP
y1BfPtml/FFBqIah/ScUMq+F8zrlyQMWHfkKD0vspSjAjn8QheyrqHrpiu3l+52M
vRr3ptXee0z/xfnRh4lY7b/3g8mlwaCfVv+dOEhqEz5IzYeYmeUQnsjXjDlCNuko
Wg8uzEmfVBozQdimIrGAH20YjLgDKnij9klPCa2JKNPYcHp0o1R4KL73GyoVavxD
/n015CP50cz3tRZ7/RPt5o01qEgc2QcmbFRGMirv2ZMljAvzqgU+HRqN9eisepQx
fa2dnU1c7jIknWIQmGaGWrIqbR+NOKPjVjnr424aGI8uz0rimNWkDqjDyTKiq4Cr
36Qsnw6JnV88QT+NWsohozqVDo6Cthoe9TJmOvbFCA1AeOyVqVSsSu995chJwcfk
ETLJO0fOK9ycfaYGgfZyzZcpI/h4sCie9CWEMYg32/0AzLgd6I41JpNmZubCgwQU
DHawscq0LPyC7zvlN8vUpq50nO51Uqu6RPH4Yp6ioWsjoV73Zx8nboi6Ft76wRK1
rn+YUZ6huBSa2Z+VDbVvEf2VFteq9kyHVc4Ke+13lLHcKeZfBaCKeqAMJOebJTms
BTxF8uNOfQiilh2SnDXXDw5p2szLkAC7R7IpdomOAt/11iS2HuQn0Xg6TioC90DS
8CebA6FZSHujUZ6tqEJNksfDsqmOP1mZjAC3Yu1TZYTI1XCUYeFdkGHJC3EbXHJ3
iMxuw/LqavCyEAoDYB5qJH3SwsGu0sF5P/53puSd0AXKrYVVWyxQ+w6VFPZzLDSV
uuXOiqDVNOD4RYqz6y+CUIkNw1o8QEnKPuhoPF+Ssobzq3UFPuNynWmhnBYhI35D
0bEAR3WvJ/ceOy0L/gskJ5labckIkl5MPVKI1lF++m5yNj8Odxo7c1/noFrRKV24
gBteev8G6uEtB3Avn9TPfcaQ3EqL5S6xM/T4sFsc+dXlkkrmihyEsx2KmFJsGCVn
+TrmidjAsN2ioKt7FQoXvz7JIxcXsWEtqMwPT6raHUvWNOYRfuO7dI6tKRHzc5GX
98mvVVXI9yHIvTzP2JhjB5vUj0VfEuxoa6EbcvjS1aJBHnZk+clPw/Btidg569rS
rOURrAFzIcNtsAPT4+yJWtnFOXIDBoHsNcjATBuUTYxlLlVTrJ59nSVp2iJy90TU
el03uMwV589Cw0MY1j7eMktM+9uKXKr/MIQyugeSOf7QKOgolg0zMAcg8IzjfD9I
OOmQXLt9FhJBQAtOKGAkqmUUrutaPqBP47MNfz5i+A8azIJTlg7fuQgX3GMeBQ2S
ARs1USUJCFl5So1Cp/Xe2678oYYoT59b1VzDxk/9ESpUpA84zIV7MuBNpLniFVU9
eIIbpznKLDMHBktt8QHbkUwJ4c/x88d2jgM+lonJ6Z3gHI0brXwn9t0uixnE+06+
4C6IXC9nAhu4gp2AD8XOKODeweCSYd8UitQExk/ue6fARykpHe2oTg2/sUrA9xlW
3dCYj44k0JdNdG+vCwyFoJue4uBMF+AcK5Q7pGxQZm28FAR4D0hSDyD2Qgyqcpud
rLaAd29lxwl+qaoBB1frA5SQeBOyny+k9llF8NGBzYGaU1M+2qpFlZA3cvKyp3Tk
0xBsXJkxO+Gdoflq35WN7GsVJWT8Ok47eG03+8Iw29sNNIOX5SBS//z3dMusdeIw
YMJ5/+iQi+VxR8dwwoKkpZsj8qjo9lWt2PTRHDvUYp5xSwVylUl1fTFx80nnDAg/
ctOh9etjcdd/JEcaMktKVkeFKO3pkjxmoLwOqjAUJeGA2zZJihYk4liYsU+y5HSH
DMHw/kYtrAh2KEKWu0aYiX6K+t0YadZk9apm3vwcYEWGRZpQwN32FirajYkjDctc
1QX/HSboLlBb1A99y8N8i6Lpv7F1fa70S6khSgsDxbMW9CCrRknmH50OVQDxeqxA
fft+ropBLgdz+bWdsKR/Fdg9Vzi8X9RLFiHL2lbGfsXlJ0A278KUbtpk+aiQzUls
p/P1yEqyeUpDIpfWefxktYY7INRcV9vMy+gxYmnvcbt79qbdMJFXrH/OuKWbxwXS
rMGEaR/5S4Z0NesesNsaViQCwVdcdWIHfNO+sUxFw9twW+zYrG7Mp8JI4Y8w7vIR
Hi9n1tX3BN+cJENhEHLeeA==
`protect END_PROTECTED
