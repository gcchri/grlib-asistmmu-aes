`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78740c3UR0HqYq8hZR+4kJPAwRFxDQPQ818HDFjKyr+7krgXlIeCokaINcn1XVqY
4XQy/2RXMyJs1ABApLWg2TgFdqvwFtJ83DMOZIvn5LSz5j2GKYYkKZc0gUi4zkzC
bCroN+hohJbCjyflusDUMAd0Er1+ZK+8CZ3SLKeXDx9rhrN/l9QNrVPyq8YKsBMT
eQg2Om/IowJdSqMAT0e0jfhC+7fp6Ase78/82KqF6CPYlaFCeGluXeJwb+nQXMQ3
7Om6ZNCLpd01YUzqTCzlgr9HEiFOwqFFKDAPLqvhmNvoDmcv5vruQxv4/NzTpBx8
OLLGVazp4A5qy5UUXkV1f5njIPUAzrK+z5nFpuEra3OeonvIuRGWovvBrSHmcdO/
h0tT2urjZicVK4Fd8QQiGrMgFNziguulw/PuWNy8D9j2VXArmid4AXiLH9QbxIOf
SZ3GrdHV5MNOFGJq0z4kQGhD5MV+uRtusMeL83a7urzm1bvgA/DwyJLpjiFhiKWa
6eE5YaukLOrO3REd/o54HKQQidQd4Etj3Fjay44YGDAz+PptDqzrUy/aNRnrvxpQ
PHAWZUjxgfrOJKFqpncLllveGziFb0IqrFmn9G418fI=
`protect END_PROTECTED
