`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gHM289jaLWHVCr8w8ivDsF1EZE2lYQu77SOzWnAV0Sce2UunrPSN8Y3p4/yPWHLS
nKVCua7waONn0EggzpeKw+64JzkBjRjI9oK54oy58nM4uGBTvdwxSwak8lB6rKOy
gdCwJ4fEYkv/VnemOgmPqjfCLddstzd9dMKtOVTIBZ5OLZ9nWa+C0PUEc0LLxN1p
Gk4S40LT98oGXAdq549uicXV4sOBYbJ4+fiMjJnZeKxklDroJOYQtTNa1pdAmKWH
is5cEncarFgZObxDlSf9C7rGoAVV0TFVykvh2RCbmNGhN7hHItyif85pm6azumW4
DtGmBmYVKWSEyjoqDUwJFWE2eWV6ykGkYb4zh6scEL1VcXOih+DqnXY91/Ca1gzj
r7OYGu6osyUNJ7d43raqcTy3uFdXI2p+HD/lb9nvNecxLWXGKEJA+3GfCwzqYIn5
D2Po5HOXTXYiRXRuYVWF8eDzzR8EoTnUFxgQxFpfw3wWDm9+j9q7jmo+mKzPMipr
Zs2shaduq4miykTP8w2zGU6N9WlNuu0ixDcTNJM2t+HAOoxbXS36aA+RPbwwYT/6
5O/F61yHRZzY0fUa678LjDUtha+Qi9h0qxACRFeMGswi4tqwBfQsDsPqybG/MeH/
/R0/7U27P0H28yzW9PgJUVPRkRENdW7tgx7FujlVU75vkeZzvg2THRDv/0tn7wTk
`protect END_PROTECTED
