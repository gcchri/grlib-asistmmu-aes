`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xyvUsUob+TrrKDULNu1SEBAVU6C9E8PDBQE2sGgWgSKWvLCqKqmyzLnWePDUqJ0g
quTGMDdmhsGKGIoFJD2orNvYVysDaPh7uH80RmDLjGRhLWtdKA2LvV7r9+0/+5Mk
Xr2/wWVglh/+/JjySd06J5Qk5F+wPby8eHKUG+mAlreTETh8PDTJjDpeNDJ1QHKe
9mN4hHkzeVpg+SOO/1T3B0WsbLiU90fIRpe+WFDI5cEBPUfqv/9TQSJX38e0zs8W
+NB2Y4Ei6fWQj0dQjZaND4SKq1gaATX7Hkeofi4EYb3YBI/cA9hvmPAv2jic0wQc
maWh+1SwB80dt4OphSGIkhaHSJT7VKJS7ApATe5pB5rWPuW6WfbvBrCCTp1qR+7u
`protect END_PROTECTED
