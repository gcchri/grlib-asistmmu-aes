`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZEj5t0r0P/M9/FXi/1AsFDe9NtntgDkyY+WVl+gbdhfF324ionerecyujNto3xv8
gJLwEk66NYqMuVH4A5iNs2E7oHHzvckHkkZwj3zF9tWOLXZpraYlkF+TMU+MxZIo
sEoSih/6I/Wil3SmCut5hrIWurlK8bukIzHCky7XWGo2kVdyJsqb2vdIyRH2v6Cz
AYJTwAvAa5PBsYqPHEOa/GR2lx+KjsOS+zh0JozGAeU7fkcNB5r1/y3DeI9kbdB0
6pQ+HAlaZ9qi6Nsp+U2A7YnSEamfOFsT5RmUBKoz/0uV/apBlA8bZQipjdc8gz1y
yMc9R75iVWAYzItX7kijS8ubxzctfwO1EDfQsNdwqUUaDVfXr+lpfKpw8H5aGOWk
/hdu6nLNnxZ+7gkpblrek01YcGVqrlV8fLKOUDK12d5VWvfhgFgvmLvHZkLiP0IE
WiqrzEPtzULFGbDcaOt9yD/RLWsKZLb7G+L/ha4xF4+6U845Wh2KbxOZx8/lCfVM
6pfd5lHTmu03voOK8bRy6fvATVkFun1EfeJI5OE4+MtY6TCoPVRNwXyo8UYIePFK
HWLq54hs7Od5yRgE6LLpwJ0KTQQN7tySBQobU0c0gO8nGMvDbYNKtCht6rlbGGfJ
s/i88eMhTJfucVgmWtZ32iETlLPdBmfRS98Dc8G5ReeIT9ZKjmW+8yPiOM5YY1r8
+UaYerngOf+nWTgO4Y42SA==
`protect END_PROTECTED
