`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mltAcvo0hh0OXX8EhzisON3GfIK6NHd7OUXXsl817ghG4Zym68RTUmJ3kwqV8oha
qXnuQwavVFd1/TaYu+USbPZ16T37GJSM2syw6DmYLtQe9CpP+WtgCQ0iqvEWRftq
CNPogcwAp+wHr5Mr9zv9Kqu7af/gAO6ffi06NC6DeBTJ/VpvAvwvX6kHIRNch8Iv
6OgELrqhvYi4onxXvSin4k5yQcSP27SsmWLbxiY1i244Kki9M0CaaXaYmfTIJsZD
tz54Ul72tuDwxd9PtDwCt15o4jDOxDZA+iFZoykrgEOh+JHLK7zLWZrz1jXwJkgV
e1lR82p/JwOSagyd0TNpOsYVKOhExhjQgV96trduhl1fx0R+LfHAsdDS3nmJeli5
UKjfAP5UTedBEu5lHmV1UyLMNGjULvo3/pYhiMyQlFU=
`protect END_PROTECTED
