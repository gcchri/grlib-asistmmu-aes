`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rz5XGCmp4dXMNzgBAsr+6yQ9FKSTB6fTblTFiX1t2QBJjEe9RjuOTY8550V06kc3
xSP2hYPxf8wuSFFVeEGjFndTJrGnA5rRxhdKmPkdtSXgps5VhA6GkPcHl4FrTpTT
GWJ06RhDlFVqF7Ox5JJtGuynTAQAnyMAzRXFY9gd7IXazCvNdHHFvMzI0k1bRm3x
oO3u366PPxzEEletovodDkRWyZQIXY8mSH9i/TMxESJmstI/SJpuvPqYkbhJJ/hv
HmKVv1mwYADo9JIu3N5WzvjQkVSo5d0NZ4Yvdx8ta7K6O2ZlRKDyA5ZpvtLMfjXa
hLsoRzI85zGUTk1sY51QrITfudzN2iA+U3DuTx/l5x8AYIxLX2bkvcUP80qO1tLZ
LmW/HiARiRZybztSbVl/qvgOrb01wuUGFFrKqgoG5n+ZovlbiUt5z5yjH0j2twNe
9UxnTvo1Quoh7N7EFZc+VDJztARvdv3eVsTAh0z+yTZ7Ds9v5KAnF26+xkTZVpWW
CCfQNgPMxBTtiWW+eEH8u3PNZT5DjyjvxyAM8kJDFKnuwYlF55B0McSL+N9il21L
+fOBl98J5L2a3H9hyK1tIY65L0nZCMFBsGr7IPIEZ4H+CvlaS1ouvEVJzX7MSHFp
V+Iib1W46WattqXKbaXlS2flS0CGwLw2rk3QhJMcZMq1VGzHYfpyHnTwtXN5dgt0
Yb5sO6axJNrAVdJWHdjcZs6jedi983+hj+t5rPAp+8mv4aZfwaK6N3wyeituoc9C
`protect END_PROTECTED
