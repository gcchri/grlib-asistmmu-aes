`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Or1QXK+DFpgGZYMQUrv5LPK/wqE0HrM1bSnhMjwO1FF+UGC9fvYpGqSk7KkR0uuz
xknXcd04Puspuhhx5K5fggIJ/cfIcGhd+VNtAtie0/6fAH5i7BJQVJG+mkwMSd3T
tAXIQXvGcMvOkx2fyOxTeWdC5XCZ4d0CT9a3J49zUpck9Oj/gax0odpmZNuhyQPv
a2CH0XToJWcChw7g7DZ7wvDVo1O/tvXIV8wr95nSa23FSTBRBpKGSuciRgAbJHGd
3U/JI3YlWnmKJgS6in8TNjZoxaGBZ3jtfxWGlaqHLhVZwXY/7B8IIfY2nlke82hi
HYTydASeso5F7CA/Ya3m3laSqn6m4A226F6yL+nIrT6Z95es9FgnpDRfbBVvM9mt
glt7TEk0XchyPglEwvtkrQ==
`protect END_PROTECTED
