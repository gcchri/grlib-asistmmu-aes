`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVzPVw4GtFWnqdTHO/5NIGkviuy6cbnuD7WrYayzy3Ec5oWoz/Zd2ut5f6gRBWHP
Z09glci6nr3R5BsoU8Stf+6mK6ikK9GYB0iHIBetj7xHKPLPau/xWovVCPOvO4Aj
eYrMqhaLghUaC/Qgdr5rJqwjfLoG34evYdgMm+5301Opnlzrg68pEXEd1IGjxfFF
3Hs6kFvHl1n/pmKKJ/k9u1z+OBPpXk3b/8IGru35CjICIe9IY4PMiNjKqlyGnScV
rIkbauWkXPvHtCGeTNHqtoWvqwjCQ7kdy+SMf/zWwEEI3cBmKIlIAo9a+nxggHTm
gZ3UhRnA/WjRp2IlzptEaLcuvqYJn13H7V48bmFvV3i+aPrhVkkMDj8OAq2591XY
Nt0ZGZz8rftZpneBmwqGXpfnQHwh39y2cFyhwN3i0zKTocvdueEhHqFhNW5GtIYC
u68rsQF4f3YSNxUA//ZH9hrJwYqi7Tc6kkqyiUxyCEPTDbbZx+j+N17VL5sp3dgd
EPfBAe5ZoAgB9VRXhR3ox5juqKNrJYSGFp+NzmfcpB+MtYSsiZSy7UsaKU9bMSsf
Vlum65/yIq0DlP2549wiZuOv5NAUG+RZz61X0IWqhqEP9Q/rHP1znEWKoRNm+V/R
2RoRVBKntqz3HmwLX67TmGs1ACAp8fKw8DAunrtQSZL2ffAHUTGxnfTiHY7SvNlf
WcEtW5LA4JuxqWcmPaU2rY1mGwX1UG0Zq1/M9mAsqWtKeKqkcy9/dV3YF/HbrC8K
j03AU3k10YjNv+DuuG9htEwES+gFmspkFus0J8YO+BH9NG9dhPGfyDQbs0udO9Dp
oMxeQnZlH77bCKcQY5OFcwVABQyEW6x4H/2YCjL6snzVZ/5I8xbcRCZDEaRCtKWI
w3ZHcJVsh3lH+d1jKrBGuRG+eq4iBMC7ghUbGqVIFWqnZ1lRKlSZLmRu9HtXykJU
9HzBiM8oVUbUFUIlNnFNI8cviDC7M5hwk66b/ZrjK+JSvpFISpxe9hHjpehkprP5
`protect END_PROTECTED
