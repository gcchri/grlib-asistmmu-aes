`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzDr5H+GIV2S0AKQ4gokFwb6ZcOkqtI7vZrmr85zF+fJOOgemQwSv27JTpAusXS0
4tMuBtDft2+hOh+pPs5GlKEP9W0Y0XEy/Sd11fMNWdjJ8IGte9p78qoeF+xdvkaE
bJSdjsmXarhhVvCYRT0rCWBAzfWaibxcZWF6rgNeGo1ojwjGwcnAXNOSp3LlqmMd
Gkjnn0IAXb9AoDiD74OLlFuyYAIsWmj5LFLIHDIU8p55haa4Z/GZdjElO/Ip8VWt
Q9WYRshGSBPBPM0LS33YXNLXC0nCojFkV0FbQv+UCyjt3dlqubWoDt9mCgbktPYI
6dEMFC8Ke8PShn4hqWwbKt9vyLn7yYn6fs3snWKH+1dfbIcnlkQCN8AaCE4arkln
KZEZ5tG3kJbB+gaXtrVpS877Rnr2Ac7deZmUqaJYgoFhFY59/SdKlWKR4e83uy7N
paHbckeLi+jxIB0fMf2gM8fEeWsz06JamANR9uTF5ZVm7wNbZZdDsOfbg3esFj/l
1tvNiEJxLfOtasrO31fMdYbDnmcwhu4jrSVcvF+RjFrfzConkguW9bGAOj05rVyY
b4FCLw13fcOW8Q/Of9VKD3a3Tu79Igcftsb88ddbWOWxm+vFIaoLa2TtKlPw/yG/
HirMK/3rLDh575RNbV5C/wUk4X8qwDuuHhI+4iI2x6Bu/5QIuQ+bPT2td9qdrOIX
GHDwGDdsZBW7+L7sZLTOtEroUFrnRGyVWuwhbHUTxMiBlIozmrrGWPizV2xERN2v
t8oVkuIXdLZzyDHRv90DXXlx3SUPSOgOcPZ1cFn2TvkKly2PFSceW2hXKVLBCUiW
ULNGWc+/d8GmPLWY21dM7RR/gAGhHRHftbPZDEQ7NZ+5ml4PmZhaXJoUBwkNYFeB
IsxUOkjZZAXrAGxVC2a6/eQoBCHaJWmJeqdrrgu35VJTG8XB+Mw6SXmCvwAlmN4h
VP8GCd3ywt21wBQFxqsYBmOFHOy5QW5CntAkmEhZpRFGmw3SUb3OgPDEXm7sZVc6
gLDtjoYWRNVR+LzQOO/zkzPojpuM/7G7D09Un0cNMS01IZTse+RkkIVL8JoMfrIQ
W2BdRkXWPvoeDADQRsQ4kCmQyK0cQ/iw/q+FXVVTHc+94FErb+ombMsNQKHivDjh
l9rQYbFrh+EcoAm6oAqEKj9YbrECzuDkBHJpV5lZL2DZ5+6yE8upQAeBXpGDBOaH
J3W2l2yk9+aPIEWr30hJaXmKnSqhV4u3BFqvv5U8vCox9OkChlT8ri43nOLkjP6c
r+lReMWYNJRZqXgVVYTZLiUu9n6NaOJjDT8mWD1FyGkpQeB5vbjePx0jTFwLQrKL
UlVt6bGaRbe2Ou5j4/+TQSMMTgCDbY2pjTnSWuV4PWOsDWY/1NzSgXkDUonKkKzi
1Mo/wj4F/n4QbY3rgkqLOKNjNyL7Yrdj/EqSmBT0F71HCMPahwOzQHyazRXPXW2K
dprzhLyxuCLc4+EDwUDaRR5rPrjRFvR4uWhssjRLxHBWE+G4v78RIBKEmxrM4pYk
q/AOG5ArDOx/chWKUA6FUilCGCxBAuYaDbA/ZVtkYbdw9JmWFxymeIfFWfnKhLEa
MxqhkKp1jkzSFy3xS2fs7BaseeUDRxrpXhasudKBzB9yDVUEsItAhml8HXp3zyof
5GvHc0VuF/GDdYUWgXqt+MNDpy2PT4hoPoNIyEM8vGZHZgTyqPDK+jeWDQuKKTHU
kP2YLUwPwCYy8amuIJUcORCZiy/jz9thexhC0hvVF+1ndstgq/8NSatkYWR8XviU
vhpW2LoC95zXU0Mmd3VGZ/RC6LJ0BEfHP7wgqmyNUBlwgYYQ8QN2Z7mtH7ToKfdx
TMkmI0bv0V5CzzhrLTajGkq2owFIi1ioR85mgJo2PY4iG7IdUQIMcpVAT3bHNJV4
3eIH7difQyY7vsYGcU9peN92nuGF62ocrCpluQftqUZw1/v6wfvLje/dj/FAeMcy
9Zou6Wot36aIJJaOUqpdIp5HFUKn6A3DSGRlWue+3HMsybay/qzMDvua2GhyC+Pi
tvq0tgecysyoyAL7q8F1L3zmNEY+/lZjsQHVCbPzYrQfCQ5fUOxuHnJhBlPQAIGO
GSARH2mwj0p0yqF6EH/5JbAaEo1RQEERR6DalDz49yJW2gR8QHYa74GOJH/8XLy2
kxCpYn8y9yT4MDbCmG2kENIc0vSdQ0S5uKX1M3RYyq39gMz5zZZVhiHFPfacrRem
34hgvXnuHcFBtOXMgvJHW11/Xo9b0ErrkTFQ+lbRqYkiEUrod1IutvY1bdzdmg6e
MB844ZEPts6wWikOAeD7jttezHUuXvU1qetrg8ZM0OzJLlutaX29vbZZgJD5LBIP
z6+fWsCEae5fFZWbgV2pLmTVioZR7k4wlJYDIAQCxaUPdcPHHwr7qCp46LF5kn7g
HZBbCBYC2EL5xCgF5StJt7OJPUhpPNIMvv5VTBR2WjwlltaR5dnBhTvldJ+4gIGe
1nURTNfg5wxAk3uaF3f1Q+rcl6tAGMZvp1ZVPmkYCDQovckHUv+PegSOKBoy+fGA
/r9IvAbwzg5YGgF3DFkiTBRw0hwCZ3o7b9RiY7lItMk/H9UlYDabqgHP8pnPaMHv
OH24/sPnYFfkV4dVNTj56rSyXEaCCQkDPiQvX5DHn/UdNJQdAYVt/OgMeywSQ8PD
fXlwa23G46XtoISgO/X65WLSmg6tmswFEMR17JPj/TBn9kMwruiyLlAD7qJFvQWm
o/eSR536ElgvJVf5tsz7l9eyaU3tLvbZPDmzGO3tAMAy6v8rYflG382mo1UyFAma
rkzlKNNOv+Kf1/hzNRwslN10SZRm3sZ7wBCWqPVNGcjiTOSwrVrNYgyv923CRp8U
dJuZ4/XHMl0m7Q+527X2xG/5rEaZrqmG/ib6ThgqzzxjWM5VOwnWQZ1XQM+rY9GF
GIdKI8ZfD1cxHFudch8dT4kqm5j3bZnXLUyMd394MVF2Y4cdAA9NHtDEVTf42cQ+
MyiA+sslCE3dDB+/ETcz4d0E7mV1aFWuqMjLeBA/L33lrofsAf7K11XnpeJATaz5
eK3oZFn65KCEWHmTcRalmznHIo9u3oyf/kAEL+GXP6nEJXZTtBRTxeOySO1AAgSs
BDw9qCBuXSf91K/Ws/brf9JSgZLGaINm7ym5fsipiXV41IkKe26g7Zsqx9/ZjW2s
`protect END_PROTECTED
