`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4AknBNNYzmleclVRg1MHpcSTzI3pF1qQCI3aJzjWHMng/r5pQgZNgZg97qAPuQU
XLh78nzrzUUKl99Pp28jFuThb0ltg6V6bC0ZXrGHNVzbt8ywZazIQDv05o/LHV3l
Qx1sN27FaIsFaJ4noNsP/B0qH19rfek3AOATyUuj3OlOnaTJqtZ7Aya2OyjuhCna
Ro3ZyYh2ucjUc7jZ4ngEbRTflyg6+IHukv2zyJG0zMB6uLETeoKfW/5S0oTaLEXV
/W28V/zyAF6tjhnR/RAfrw==
`protect END_PROTECTED
