`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
St0+NmqEmVwsj+bPJkEpkQYBLtnmdGLZv7uglhGutIoY3Ag1EjzL9VehHfiIpa96
Y6G0cyyXhUDpEdowXHALNoggx8/hBPElanh5XtnAMjVv2iyFF6EQMNz0jgir7Z/d
nKf4raVdOa1u23zfVcia/QuJCJx6ADuCobxvdEi6C+2yjnnP6SBj12Kci/e354i0
3sueI6iNQEWoaZe0Rxg3jqqX03ibdTU121VgqSulA41SCzWIFLYJ8KqRKOTjw/lE
FhZsn0k2ZgRMW4ScaXBkI4FSkMhxU9XhASh/IiiU0C1P1p9YdJhm9V2KCN8LRSJW
J8wnY07uE6IEGzq1yU+P11uVN0GHIy479CYJcghiEWJHEWjcksfAOE4+gY44yYHO
QLfpobeRLcYvvQOn+g78fwlZTYST6HbOcQ5cbGc8Q1DGIA2AwcKM2nvOZ8FONolT
u1GM0P3meq1838HP4bATSjjSdFumYSFPp97v5yLePCo2I8islExZB6p7lBgsBqsz
9a310Ew+A+u47x0bD4AqrQ==
`protect END_PROTECTED
