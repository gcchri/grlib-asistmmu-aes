`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UoIDXnVL9CeYcDKCJfK/FOZ5Zs9lUYwF1gkOJXNiJpRPdgJHV0KE0/7j4B/HrtVi
zxB0ElrPZmSt5tRhYM3PN4+OKElzftBPwZSOThzCr6Yx0Nr3YaKH29gW4Fpr8c4n
6i+HlkDapaSmXoGIxnVotGPIgveBwHQtc6hU5X/Z0MpEF4Y0qM4XZjEiCQDZ+Pz5
EVkXmDxSr9YotoGHqJeuF1m35jzZFFIhtZtvfs5wd+tm3P9b4kw7jLoADyk+wTS2
48DxKpMZEYYsrGtOYRKDtmD4dZILvvPH/Uww7WIJBxQYq0jzJMJEW7BqrYB2Y7pc
VW+Z0mT86VqK5Avt5fYkglcwErht6yQlTxb7Mk8JJG5ht+pYSSVuoMXI/VLjZt/0
ggsoOnI8MzqkpdsmMll2eQ==
`protect END_PROTECTED
