`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ipHZrqwdTWdWv5biLbugogECuC3vyaRqWjamUe372cmlqp9N7KRm4YTNpNuIpHj2
UX//NNbhdMY1z02N4GG6VzeQ2kD6KJ9aBtyxII/pIqmcZH8YoOjZwnsOXHRPUj2z
u/LO4NshdtNs4Atu+4PIrbmtI9zUukLnFmxDnR27W1plAD3N+OrmXTwrMwyI1gSe
WSvpwrBsT94nA72MdZP3dOEQ/fc2nqxNhDTxk5u6SKHI4PhHEL84JjtxXdpFwMUl
6qU7YVQCv5AVMbBV3Cf64Et5llx3f1OR4xavw5WZDRhopg2X4Q2sGMzZuEYnRDWz
2uC6pVlBrCU2YUqCsTm+JMAZiWzpTa7ECzgZ2dcJBrhse8P3M2Yy5xJ2VDiDOT/+
rjqvRKSOEstL2jyohEQrZswPbebDDWT6ZE1mnBTFN8Di0cLY2XUd85Q9s4OGtWj0
C4TyszyxufJ8VfgDktMUbDhsaAcV9AfkIyHykx4xi7AAg+WCZas79NmnqYsTls9x
VOqvE0R8Q/HjtD8T4hrhFUJ3O4cXaWhKaoM2CZ19J0m+fGY9Ec38KaWiumDojw+t
`protect END_PROTECTED
