`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sci8vo7niLx7qWl+kQc3esaYo93HkTkQkDDmAbn1JmIowJagnRpa35KHdNgYhwQ2
1ZfXScVt+kmeyqyyYpnvmJ0CB4lz/IJxM0gotVutIasNt8ZqPnbW5wI8vbtDNQB6
FRxYayrRxKu9ZzL5MICWGCpzhp5ZjCmp8UYCSAxT3xfCdA6hD26NiSfLzQsinifQ
X0ChYCkVCaOf2s4WEr5N6sgrc+ysL0yyDQFhmH2Z15Kb4z5uP9aMvcWFeeiRlzCU
sN1v0sqauwySB0a7yW2T0a/3XjH+G6BDzrpvGNxT7s+YcDCa9KZXOSVwttCl3Rzs
updgFrqxkABkeICPZeleayuZZ05eTyFxMePQ34yrdDYj1akBDR0BTZH45dFx702M
mtKo+VqJCcer8kqCyJ/sYTWozL9HH79ZUUYIsh7sGEsalSwSfgvGWxzMl57nt1P/
ecm0xCF/xUlTBUJ1bFQ6GXtMuIQ9BDjBvs2u3mOchbD2eMO3gq8fMZYrYSuf/vGz
RBhnX1v5whCSRrUgEnDwHepRKfoRlZnTz8SAKcqki/UuocjPU/Wa+dTIgN+oQQjF
gldon29lGkfqknj5ApGSORu74f4M/+lpPbmaTf+3PNvUM1IrxrCq480bLHGUHrSm
b43Y/zRN+4qy6JCeyKxJC0ORMfhyiycUeV1d1I6H/SOg1yiRDt74/dfuJqw9IXtc
xQ5GEtNggFp0jERzThpaaLXvjb47ktFmPmwnP4Q1Ovxx4y/fOBw6NDXiOl+K3iFl
CmGnxqs1LXHmGr25HGvbm6fL17Qhoz2b2bFfQM6aPjdcsb9T+4o5GIWEm0Mds+H1
ih0jNWzd39vbP559ddvqxEDzSbJ2b3LmN4BAT2Dzy2HfRORSjniTiEXKwU422yZ3
gctyhc5kBmrXoG5XHuNmoA6NwCiOSRjKvywzKscO4YKN9VU4bwMWpyTO9EygXCTA
v5gcD96Mk6tohbnb+gReck/5ZCA1AoNpOnxRaAxeWp3LqNsKSVyDESC981ULc00/
Ig3EqrL35f69AZfGPPDTaKpYI+VwggRqYpAd5N97Cgh3FWaosfIYTjNN8VIj8yYQ
r09JYAhduV2cZa7vds/3Ct2Lu3TVpl/tiJZMEP0iNUdN5w52imfAM8M45St29TM9
r/stxbXvmZh41/6oEq3Oqg7WSHqmGsQcoGYEb2JdBCcgYH+F/OY9ooSZoA5hwn3Y
qzpeROa6e2kmfoUQtKEztlb89lZO/wV7W/58C1taF1R1K7Y1CO+78E/Okp5UIjq+
1HOqljjtkg1ZOlY8C99it0x4Y7V/FUZXks+8o4AFP00GPdLruBHWpmfsmaX9r9RC
hcjzu+aldxrbwlgiBfqMncxhpyHx3jUrZCAanvgVN5MAkthNdg1qkHJRMTy3zNdT
7pIj5wul0+USioYfaya5HPuM8DCmjrXjM2b3U0neJCXNWOznPhEALdvu+89SaPMV
WQkTz96pjFN+6tu3hDpynLBNew7huehM+oTmyMluc28=
`protect END_PROTECTED
