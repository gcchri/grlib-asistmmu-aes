`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6rJtYlPDRfE/5MBBVvU3xIN/ilQDI0XF+K08sQYUradKiOujIhmsPvv4eFKnFmr
qBR+LONiaVUAoM2OBSHGb4pKL6/pPo/8VoiTWrHyZusUPdaLcYt0A8iSbYHLvz3g
EhOTBgs2Nj9fMr8LiY33IAGK3imZ6R1y3OdBJHvt6j7nK1dizEGTLjrbAlxNENvE
iGLCa1tmq9IrOFV7RnuD5R8J+8Rd0KFfdvWKByQVqiZZGC7AEmOD4LAGU+Gcektx
5khLSMWk63r4oBPV7vVuDtZeKQGyczxwA1oxzGkU/c0HVr9T5Rn5Vm5ZiiO4mcBi
FgwHdptSQyPGDT8RnC2dMW3KAcQKg34tr3UbhdU6wJeTFjQRPRAAzBlRtR8XYKCd
h5pfA0gnNXdmreUCisJDn2kXR5Jq6+B/6vIE8lulpOjNRI7wieyTWGnAHzfY4cSn
Pt8VWStDSsD17RW0fG9QwW7WTPQkiM76lT82gZ9DkVgsUOxJ6YU8mUT+XJ4CM04J
3RIcNPKsAAFieDxX4VkcCRoMQ4vGZhCERwYi2QPTZ2b6yDYvC93vysGOmozq0lP4
ncUo36QTb8huwTtowtpxtYZrPeNID1uFmvcbR4DCtLcISHrXi0ZTs+B8wgatSX/u
AGRb365oKD9n0ZKeBY/gaE9RZhXSgW/3Vmab/1Bu9pWEAgV9kkhtm1uO4bcGQtYO
iehCxicOMK5fslnHKOnWouUMoc3Pcorf3ElEi59oFNoAanVRuqCHaUoy9HjHzLf7
fmNVRXqa5oabC6n462HgzG4N0hm2VVq2PeJqHKErhnC6LgUpMr9v1/15S9wyZzwE
imvM0SJ1f3Cc9g4Pz6BQT2FanQ9iokS6Qo4THKDsL1kCv3OyRCqx0haJVDb5Tg1Q
Um/37C8tOmpQHpUdD6gV+K1UBM27UYRVLs3fbq9lNLxhMSiFCgLMIopc6lQSNy+v
J73zYs+p8d3FgJf99aoozOUjX7n/B5rf9nYu6iBAcNa5nLOdspaQF68KJtLcJiFC
p8jfYa9RIswhL0omXDQ0p0h1c+BUON0CaRv2PqrUt2/QNMFUAC9UByRH9IIrpvpw
nIW9Nns42hVSBUZEH1IEz+XvwTXkJahJTLRqnja0FnzHMXQCTB2kmy6C+aC3jl8S
xnSMPB+vQqxEcuSlRxnd4Xs1Z9ibJWuFnmvYYrbWbHyZQ+OaoZo4PytlnjaXNX2c
HKEtTkarV4SoUlPRJJvtXtZAodCpzkHJn+7035zBizJcDAM0MX0tGnRe3uiCC7eU
QJ6iTav78D+KFhwVc43axQ==
`protect END_PROTECTED
