`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jV6LTDaetPVCrV6Q6fhj/KcABnyK9qEtOmAAnUZQYq5mKort4NQ8MIjZBTRlbC//
FG12vrnOgixH3NziDbRJYXHxJV7G1ILJPEEsFHOc/kjnZByKeINM9Jjp/Vdr6yt4
AdpREOvgFp1yJf6OqxrxETLW21wfTZwU7vucfWGMXfjzevbV4n0sTsJJECqxYybg
NcDHlwKDny4PzB9qz9wp0lZUNrJ17XvZPGnVqySRKR85NznzTwS3g5dgyRk3J6Zw
my3jRwTd8cOG6fR5VY3TlD834E68/GS5wd1vamodXTTM+XmV6N0zAIAWyLMyN64L
mm45xG2XwtMsBeXc1hgJDyIigBwv7B00n6KI+tHN6SNDEGjGtkY0Pm/0ARpJ1wKI
yh5dMc8X3syUzG0U6aiAkHLgWqJLQHIdmRrkOJri4cg+zAes84aPoHirB0JLlm8i
`protect END_PROTECTED
