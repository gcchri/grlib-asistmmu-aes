`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82E1GpPKRlkk8V3L8Q9QPwNQxbdAQoNjzxeo+fRTGr4tncyOqFM964h7xSGKiI6+
PrNC/VnO95mUFjgeL0z7J7I/4g7o6hCWzJnfqxXmUblHY0ZeqIV/PODmO9BRKTIZ
0Nc7c6lpXPv9tw8Lj/4ELABcgmQqhLeqje1tqdJ8llLpojTYu48ZeOm5vuAXEnJk
FP+r2hsAoqS+8chm38dnsym3IKFa+O5VJGommQDSIV1uGRglfJlDSqrL2TTwytLo
JvP8OizCznEQ6gdCENIVvrNsvXH9OQ8yqzRb+sfMh4r0hyCcyoUiKQltoEMnTrbi
rinwRL+/zZFjDdDdBYKiCGBOLOkyb3uWisuuFR7yoyCiOdycLnFzO8DgdoUXPEl/
aeqzfbVxq5CdD5gg/y4RzJ5ggsyZ7ahmm3tkQB8vEMA8dwFAIebMfx6rRNnmAKBO
qHy8D7E51vR/xZy7THlVYZRuUFl1MmpwgjemPmmj34fEFXw19Njr/gqLG8al/Qt9
4kleytstATIphq7h4Xg6sNP8wF5sZAV/N71vLvhNzwL8bInCEUM/UvE+k07ecVK+
dmibvF9SPJILh6kLFSWT9yirxYDcGLaJ+iNDoj5qcs5VEx6lBQzBIefbBVoenUgC
ZdGN0IzBQ1g79O4eKG/s0tdrNYNoQDvasHUfvyO/rKRSfzBhMEL49z+tGy1S6m6k
jwVK+7weSIZ6NjlupjPAlUZfwqBL1JzJSo4iWGROAQMHBfpTvQl6JpYhgTNItE6t
3ZQ8x5iK/FMqMJHCLwrZHeMbK0qXGRbGSkWPwzv8nYElyouCRNnHwfM2GVqPQcj4
7H4YvUfae6uFttkBPleOIXolALBcbGC/1VsNzjKa0O/8B+2giy3jfwocEDDHg7QW
LA7OrTwxy4o3CGb/eH7fUjz8Jalx2ZjWoXll3Vur9nBZSM+ky5VMG6G+46tyWdir
`protect END_PROTECTED
