`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BpynidJAqn2145IaPep364HzEKYGPwvg2FysdPsm2NwkpTb0vLKcm2sBy7Hazvs2
vhfHULELVQ2m5Lu+5i5tX3r2RGIEb+Tu5zIqom0yYCr0Tl8viFxJ28guMQ/HsAdt
kTI87NniIWuA3XW0UR1YzXQrOvhI/4r0xmLIxCCykawTunSBLo9jMVSl0hXqJrGK
kSv8zxSV+kwgziyHxnL6KREBnErxIggJQNTL/rOKL28z4bsxizBdJHUc2M/xYF/X
3ak4vvRKcVrQ+2py8kt9b0gG0gYMpqIxDmvcSTP02WdqT+7sk3VworUc1rQJu1QH
o/M6//I54B+bgvMK6ZRBh4zr2nnQYA0JKRzqugl5QdcZSBjX9XQHXnfCpjsz0Rrk
icoVM/z14/7mejXlqgpTQrhwkLI9WQidZzyStA0hi/7vYTIzoQcDaUk/ysSaomyd
2e++a5Gr2wvLZp1F0BDOJjxKwoJVD4YZeqWYK42SW689GtE9BS2+dqok98GxS2cW
ZO0uouSy29nmRE/JkTLSmIWcpVxu1rMWs294ZSWiEyfkIQ+EAEMyZdbG9F38TzhR
72haE4RDqLlaV2VcHceqZ8q8iIUsxX1iE9duJX5u6xsF6nVhAv/RrmLkdhaax3JP
ey5H0k3ZlrKU0YJFDjgzQxsYupEAyUuupapEknrIP3GcKC31PJxB3BgEQaw1mivv
`protect END_PROTECTED
