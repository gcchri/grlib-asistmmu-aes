`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vi/dZosv585ZWezodLE40ElMyjkGqlvc1t/GAy3m0627NRkQa/g4/JweIRA80n2K
Mp/KhSatsqmoaQkhwEqqgrlQcFala+S0OcQ+vn6Cld30sEOSjGIfhUJS7zjE/R9L
qptef9KM1FtOFxZHynevlb++p4C0A/bk8S5uUxyTP267MK3IC8dWRllp66x4PwnA
IoMXdNeZVTvkXkKtWUAv5kC5KKehQimnbjCrKUvG40/LNg3ZDLD/WbhsHJ/yTQgO
4v4o7S3yQPxuVnKlErKDfF3QECuKJnt896GO9NbfoHXZzEyc2pOQYVtA9cbwRsby
fgeCeMJpGPI+NTWDhz2U3nfzOc7DjVXX10/Z0Qg1FfU7yXLKhvJvrd8i0LHkwk5u
EaWv839C/Y1kTzbEQfItfQ==
`protect END_PROTECTED
