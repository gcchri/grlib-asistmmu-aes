`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A63bUX7OE9TCVP1izEFBbTmS3HdcPhpnBrpitDe2f99q28N/48cfZlZA/ZiZjVzn
0kdtWO0NxLLuAdXhnc3rNK2A4ne+qowGlD05NxWh0vzT/vHLejXHl3YsemvLKW/H
WolSaH6bFqviLwGF98tjKLRDEqbMSMcL5Kzgj47N0n4m2mRRLKc9cLNvtLKe081H
tWcAZ2pkSP4MwDWpRih3VcvD6U92TpGggIylXeJ7qeXF3/qH2CAwl08xjvl9DqYd
hQjZQR8W++raTuv0oqp8q96h/ZYVeYBLIZvoEdft/qNPsINb3Asm+cWdLp8THV/7
0tPoeIFlTQ+FCAut1/998vEfeRyTrd/fKMywYRmOtJHRNLm6e0mGt+ji1D4iqRAm
uEmYYXySBAq3lv6tb7TTT0MQlK0kFrg1XAPpayKPd5odDZDpprcaJZ5zyDpycnQP
R5Ra++eCov7fnKL4tndrHkJdhr2rohEt+8b6uS8tsl4k3YIAq0RK2jl9K2WSPWc5
OsuMKJ6Hinum4qN6vpl26SDeHlfBkjb8iky3Q3gUdl0VxKFOIiS8ms28kOIlB9WY
e9h/q2UkIfl16VHVeIXfeDX7DmEvhjDKh94vS6VS35r2Mv+YdA3HCpfVI/7FkGU+
Dz8/feHpCNqVkd1LUKRgEgQbagL/cOzn4OlE8Ykx3SYliNpRCV+K12BSPWUFUQNV
xz9FzHA4dY8/7b/0oMkKNb/Mi3d69ZyYrfFs0nmBGjyXlJO/4ST2QBT6w0l927rR
7h7K4gb2TgS1KilI/xynYRvq/d3KlAIkGDCjFH9sTygXwbBtlAUc6jAU2mgyfszx
mwDjHux9fD+fO4fKMXcPxa28ziSQifavERRywwSJFHFm948vyyy8iYFWoJBBxeM0
muN5tnIS/gv6d0tkX7s6QfuV2IyaYPaDVcN+jkZN7ZZr06HJ0hAXrv4DDIKeQgbG
jDrmnGnZkCZJFzJZ8ZqFbb48Jw/aK9aXnrV4n17OVBOlN4VqlrblssSfIFIpWtSm
ktCJVcIbHX3sIQWP+c1sLgpXP3Lf0U9IpRWUBzBCP4BHuqmonf+oohwSoLKeJwVT
Ep8atZU2edLu+wTkC6WUl/1dA5xAPdfwfdW1h9enCcI3V1F+fZN9QDAJu0KLpIM5
iiZezw3QA1wsaG9JZMHzSV2lQ0VNGU18zDcqxp0RZphZGET+936l2sA++NIj8ag2
acze4CWZ3pkqYJsEuU4oGlgZPHt3pPgEHGakV8jQIckhwQMBfQg9fChAF6lIEFXa
aWMc1Gfu50oo8CAywzsYz7NMDTJQN92nnbze79B0sIk93gavWO9hR3lnemA9R1du
XsmVEo4xQlFGDgfHDT/+bOGeKGDlbz9dy4bdY+RrZpNzRj8QSgYyPClWUUlQNMVE
knWBT7oTxUAntWqxFC7T3hf+tA0ubW4qvv0cRRFTrY1y7juY7x5+cHQTID9IkBpR
Dw7Ow8REuGHiWwBFQnzuYOiiY+iIvFYa0aJaHsI0rS0haGkdLRAf0kauR9nO0iSF
WyE+8jTwmON9xwWoGlecCFP2tqCPMD1zKu15tVes5b4GAlN7f1u4YV7vTCTyR0en
R72XaVWq+nSc73K8QqPgsP/GP1WXREajTl350lVp9bC31I3C6aPtTrJUIIO6ob1g
5C6W0WNnVaGYuba378/7qqzZtrmoDCSCSL5nPLodJSkVodbXpumTzT3LHMUrAZmD
/M7TS/LFmrUWF/5yIaknKaM1B0dxnDWPEoTQcYxP5yLdfIRMmPFLH4CCNmlscKfu
3AMofGmF6+1Jr1jAEoZfZqz7bJTyDrwCg2YZWGIues80EzjzygtbbTHw+nhMyxIx
BiqQEqBZXzjJpAFfs4slFWO/VRl1+CahDJ8PSCS7NA0=
`protect END_PROTECTED
