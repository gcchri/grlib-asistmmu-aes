`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKU/3MobuvmktRYtBVNpyPnqbkgMbT8F0NzW2anIKUokAahzdgqidGxtpqIuCVuH
H//LUyhN2GxB17bHOX5lkcnw2I5uOWQ+aulMGsJLcRwBCYebRBSot2CJEnAs+4EI
qpp2Vp0fqnImx0H3t5UHxXeMR35zp43pyaXA6KbMBN4Wta4etvYiuvpXfmaDippz
G5lAvumLt9niqVMTXp0rC+7TZKs2J2yLLa3eRIrZO6B4ISIUzDV0TcWax7buor/1
IFNAXxCkm+5Xgl2xLglQ1A==
`protect END_PROTECTED
