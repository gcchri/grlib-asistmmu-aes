`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Wj1zNEZPEcWB7ikGezg70xnlpTGFqBqW84hj5qTSIPAlFFp37ouoyc8Tt0TLuPu
tT1XwncznKO/dOYf6Y+ftXE2sW/3Yk55xuvComiFvuwaPwxiRorGQXGicn60HJaF
9X+ONrK8mKvx+c2VhlpJYrTFm0fCm8bgo4QAYcFKFuZlzTZJb7CcgXinvjXHQncc
cdxlp/QuYiqGX0liRPLWGuHp+nC4UC/VBbRo3g3HVLxKt9wkveAvvGk4dONeZD4i
//rt8bmi3ps8mBJVr8dV/yOH8U7R5kWAT0Ej7axTk7iIKItNdTa90p5N0RxkYOMD
BTTVyeOlAxyX0hD+fjHqjRpqaf2abQJrP+3eV3+yJcxXh8hlsMZ7OpBNghN+rPiF
DC+VnfFmEKp5PESfCDpFxQu3cJbnJR5XxlP0riP2RbQ=
`protect END_PROTECTED
