`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+viCSlCRXR8dNA2YmjRtirq3k2QKQdjLCfI++j2C20yRgtfMlQjxoxcQB1G/kzIA
ue6xU4/m375RhobPjiqTZ3SD+vaMEVFCqxKhgBbrPx9KjCgaNcdkQzPbR8pSOU5z
UtdZVnQg0k8HH3s96h+cyrEK/o6e/JDyPd8VOFPc1rtmmaUJtWpf7ngN23RW1CCx
WcA0KzS7XQIHlJaYwDhksD8ZKYmdixdeZzM5Rh150MsQDeymo3s0oSvtLx47Kqv3
oXmnZ3i/tst771FYv6rsFM3pqP19myOgkMDoNiOD1fu5Bj1tYMQ0Q7Q3ouoWx4bF
5rZcZqcCaM0IGLnfBHzXfD8HZZgMyghT7jDxMAYIJ9Vvp9ikVBixAHwWfVoyX3x+
OCvHei7VE4hpAK0JTQ4hsA==
`protect END_PROTECTED
