`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vlFaoki1jlNPTlcCmjfd5jzQLsiC21hNY16PmHLejdd4dvckJbXsCvK+syahkSW
K3l0/p+9K0pOXd2EFU0tDGx5bPElkCEOSWctqiPdv+mlvYQCrf0tri1xqTHM3zbc
K12J8cceBYJvPBFOpPYcd/D+5SVFY+RV8e5GMx350O1i2OLVFCJL4c72BKcnv2ea
rqgX11+jtlJmIzKaEioFOTFcO39L0AHMSYVCE2IlpJ9comq8AyLgVSrOMJSOcDY4
Yos9NdxbhmAWn0X5ajJsmMsc/dL50lCaHx/slrsX58inN4x2jPYL0sOd4UNMwruY
ap7OuWwH12nRp7Pd842Wsg==
`protect END_PROTECTED
