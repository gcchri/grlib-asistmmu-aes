`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rrUt1s6uf0nIQ/0yIP2FPE/7g5fSjdsg3COR0eFlfF0HFMDIiP8rTnDVwz7JNlHs
PuSrHi2RqHuSCVpfma6+zQ4k6oTo34jEl4c3FF8LvIgoCGUOC+b6WpFCiLIQuH8+
ZBFqZh4W+T2dc6uWg96UmPKU6KmEBuOYbqkqwGd3a3zqDZO+/vWlEDMbWSs4zt8w
viS+hW2nxUYIqrLuTjEWah7tE5jq76cwCsVOx55ZUcso65lGC3hxZ+LfiE2oXjuW
hALVoWc11LVQdK9X+AFC5NYcU2dds2WQCi7Cq4W5/Z25ULyfxFR0e7+CgY5IfHIh
qEs0T621UqyuUN5bU9kR/ZEJHblSOI23RSn+Aa9mMHeAJ6kPO5MO6l2KPPbtkPNC
B05V9ZWMu54L0jnSunFfoXhcb0UTpkh9oDxXgYb+QhWPR0kBafRz7qHpj8A25dMx
gjJ8u84ExrH3rJwCEAo526l8zoKLE+1sbKVhwFjOPbX3uCiVX9HH7M5J5WfCu+Ii
NATWowa5lALa4X7xfbekfYnxAtEzV4JZoWOU44zeLYE=
`protect END_PROTECTED
