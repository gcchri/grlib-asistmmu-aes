`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JRc+aNsN++LcYDw0vNn2UNLpYYVNtmAmXFGLEurKR8kCeJ7RPJnUJ60O3/h33OuS
0tP8yzB+xK3xhiqShPgkP77/Z9ZPzBVcgXXjEt5X9H6Orjmu/JD4F3xpAUWGqQLB
wkMwpR8XTH/WS9mmLzn51mEt0O9cyf/Vsj4FS50+9u/+vNlT8ZyBWdLnN4Qt9X50
Hm5X+TJwlzeNEsD9yUWJOVFoorY6/hdIaedQVyH3rZUy1IBKGIQIyqKBWqsrqrXx
zSKVpIMYbV9wSOl3idqJ5FVUhc8XrFlbL6+Vz4+wnpBdeb9sXcUeiIsIC9oOLgeb
R7qvT57bdqRyIGAA/Zd0XUBB9jFASEVw5LF7XaYzRHiJwwh6dGYZNKP23nvd6UJ/
BB67EDNTGTF1fmNt2EYoR8Ao3CqZbA02t0ZmBPGZIz8VY3qr91VXDDd7/+b1LEvW
+TpIKuDRzxJ+2ymHoqq6U0zqE93EoSg0oUc93dPEofTSMDLaxm3fzkOFX+/iu0+y
z4R1vfaVMhQRoZiqsMw8HQYgOHNi7VO2tGEix5ageaQdCeBSUkpM8hrlfQfGx0AA
Io9D3zoLDk+nHTmYby3VAVXSHhYzXNLwSNKteK6eE8TSaJIFDYot8TnY3R2NC7Tb
aMoHtRG5khBtae9tQWSKVKPVLUuFvUbCXWHSAmhXHiNZuBz3HOIcHZFUh+T8q137
mp/tU7atipvtdskzNJ/D71X+Abd5PGPMmtFABTBu0R5QgMs5zLvIW47C3sjfld25
zQOk39I6PehWWCk8q/VV6HTDSK+mnLexBc/ZC7Yi7dNQar8HqHp2cKlJjotSSyo3
`protect END_PROTECTED
