`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMH0aRQvvkK0ez/zT+2K3MdnPjBiZdg3U8ipTjscnkdbk1aS6Wiy8Eu5t5KOBXLF
lGW2mSdKKooRomnuZADWn/CSrXQM2s9I6+oybEVsDQwDkQjxf3RCbdTtFWDIYlvV
SYudJC4yz7APvo7E6a0bvTfc/YevPDyWmFt62wB3J4OURL3Gcr+BYlspJpHaYyfI
ZtsAiBDWLySx+Wj8cc/uMV0/CU6ZkLk53J88i9No7ItyRmdpn9YX4g2krAGO9EOx
L4utfkcUz9lf0Zy3Vpy2/4uuvtuSjDK9UP9Uv2CFOU9MIpI9IWAKlGNG5MJd9Wv1
YPLlysOr1d09fWYWgHywoVsvgtT4ncuPFBNtnzsM/xHaufRm4hcFnc8Ye8xQ02L/
JFtIIOo72ewyNH3VePIZrpgZahQzP26BPggXILuiwCX/YuKA8us+ma/h7uuWEZtu
VO7y1/c71r0TJm40/2C9SMmudh2VNkQyHB7HwutzSUivLJSOlDYA5yZcyNJ9aOza
S3W7ZXiiGtELqtyRGqcbx0OY15pmbqEhB029sPNGi/fM7h8+KPiLkYMFu/RjfzTX
lkxzG5JU6Czfki7TjfNmI3LiG8WIjfrhPy7mq5J28bPbDjkCkEuQsmxR2xk65z5J
/1pqiVJZok4J5YX64zoU6KPMaE/+mx6PNDi4HnBhC2T6Rtjrl0qt40aPaBulBYWW
alOhdglyQHRiPsOPEigagV/sjqMSKvloao4jTxjE/xkYK1uDyQoH9Ksp02lZcHMX
yaoo0Qw9OIytjoGmw1Retv7KTeY1bQ6JSl9OimlSPNDscwSQqKnkYRW62fTRX0BZ
3RUoG5h1Ten0DrYZYYt0TI+gT7g+yWFHMhG1+hDUAaaQbHGS5q/dO8+Sv0RgyP64
YWQo0MDJadPXQDC32xhq1MU2NvdtWuAOw1dNEMu8PbweAn153IBhb3968niOxk8A
do4VoGtJpIFAzusDkRHFA+aJqVsc7VBp2NzaiQlJWr3b3pRGnSpCY/KZaVVapC/X
KiyVeBXCX3oWnSI2wnZknW4PZu5PfPIJzOu3fycptYwUFrJxHtRcYeEI4d+ophtH
8+Xl31uljKUUV2C6W7ruXvC9EqcpHL1PwQa2kftOcpkUuNaQWWq6E4FaA8bBNGS1
uqh9eUhv5sbn6KkgUZ+WejSorH9tO0OJV5N4p+DIhQUH9DHBjr18oeZdinX2S5vf
d3j0QzFevxL2F/FaKIIhkAMj/77J9QA7aLI4/haoG/epq3BaTUfVWIirhitmMgxX
OK0KRBge2u197YaidXlKjvBaEv51GIxIln0q0gZVJw50C0N6wp76a9tyaksRlV3j
yQIM8FwrFedJqnSd1sIQ/ayC1smnPGn1Z/Ew++AT5xZto9UgFfIVqVED9ekOdHxC
XgjET+IGoP2m/iQVDZmszTr4EWgwZNGfOECHAhkYM+8XoRaW6c7NztGQiUZGJoLs
QS7P/dQ2GfEcv2cpWQpTslU3Vk5SE7jQg5ahLgaIlQqIFqcRAGXnZRgiWYlx+9gr
Q4Xtoz9jVXioPWXn5ywa3eoTb5iOsBGLjcxZQPhLF1AYJNu4oEO1n8a90UJHpWW3
frJ/4/56RZOhBl9I8ledKD9Pw2BxNWN3Pr2tBnh2LXtpd+T/cY+VbNdtTVjCz6yI
rPet2Tw0b4w0aqWgEkTL+HivWAhPui1tUDwgHZg4lJ796wHdkKJJumzWyYuTCR7v
l5utN0JuFrTaHSNPtrfKfQ/IFwfnzGoQQGmcyDvV25jUqGZKtmQsLzuwIOlqGc87
Kkonhgp6IQY0rqWgpAovz+qjVqA3f9OqHCFLyLhSuTILaQVT/GUOngmA0oxsCFqj
2zY3+eMdLLHMhR2gf0GcWhKFsg+u8wLP/KFLIG/I+PPqhneF8Xa3llWUroFXbUwt
7DdEj2enIrIz2IQZAWnSrektPkpXWLoT2v9J6BwA3yXNTfxyA+xecW0wXi6Y4iPq
xZHjk5GuWoz/Is4lA8viJ1Xf57umYSpmRKci0v0cJowyFxdO/AYZh8ScM1Jv5O14
2uvV4F1rnt9Nxg21ZAlvLrNJL1f3E68XeE0Hhn2z7BAL/nmabgfdh/nIO/1smAZB
BHQJYJVVfggtoHJmJn3H6SSMqEoi7wW0aRNJHtY1WulKiAGRhCZSbZ0gOL0iTnkk
S09xpAS9QxCvtvdnxhtR1J17QzPrgJxJLCuoQcOvH20IJOfIYeDEyMvyfouGIPpZ
R/KnvMU40OjiLIqhEgj5spAuHAjYLgTkgs/p2WDWMdhiDqswrB0jjpM+qOVOH1Wb
0CkuPMpPOsJUxBJKa4X/1ZoWLWM/jp0nmPX+PUp9FoGY4RzM8DOH/dGeXJOLccC2
4bniJzT8e6XERaY9x9e+VHR3jR9sZsTp9ue22FKexNqSuoGP8PRL55BVSm8h3D/t
JAKa2Cq7OFkEIJDiZU0kDZdTTv5JUQL1sjpYVSJLBNLGbAxu70Q0v5HUU8PSZAc0
DujnvzIRepqDgYXfo99/DICnhe1nnysb1IpmwFrLHyDDyiUVHtUhV2+OGa+MWedl
FrNnyr0TqlfbqdbLE6L18YPW7yI4tyksz4zf46H/f9I88/2QzZNw0u+EasyvAmmH
nTcWJyv8UilA493wdRO9Ojz7vK22Jt62ADzcpfONB3cf6hL6KVEiCMil6ywGtQ7g
uie5UwKk4a6szkczPOB1K9nGJFd8Qda9xaeDE4pZMfDDZZWbz1GULZT+Npn0HhdV
Bnn1LcWMY7YF1t2GknerOBUQbp8k3Rahe5Eab77lC44/j8zJzxzbUEfxvdx1iBkt
fur9wdEq5zW2IaI+P4VMUpvajf/GzF12FW0VJn+lZ//AXbFYfBkJnM80IkIL76gh
OCtomfdKCLiviK4sov2yYbOmK9DGYWhpkmnn323dXMvyr/dmwe2KKOP26fNhMpaN
lMUXOz5xDYaji8rz8kAtSFysTnog2FwAMcNr/bGUr5V5WcG6YtsW/ZmaQXtMplVv
NgHBRPxiwVF7TQiRlhZfZ+UTj51NMjTUNiUwX4fvdsmBXq1ttg6FwgdOd6GSdJ9v
A5saVVULu8xwygMiDMOhJ6+6DIrCzDylOoKWoWbD8cXC+lMXAOEzeZO7/2SsoC0d
tctuUL/i4oc6fJhj5K1QMu4vztEuJyVWZRhlbLFgHMpXI/oNeXTTK8xZeD9wtpnN
jTlccYFe5ha7HJF+senZxtpDA8wFZrGa4Pk0vPIw9PbJmcwCcDlrXOw+6OF7VXob
XNpdO+UmAhR11FwufCjdeGDgK+HzTzWdUAfCG+xUkaQ05aO6xYK9du96LHikyy6o
BUZHj8OBYGyOk9NhZRkQjLljCYZUccI1lyff5Q+Un0gh+Cg2HhnAG9HXbCgJUY1Q
9AU1UjkbWXCb9G0H+StBGtt5FFYfI4lvao7+54sr4Cmavu5QS1gi+YlIQfRTWzKI
SxWbPA7joY++BW/iOy99KxU1mG/l4Qo+loZPipkksL38Vl/HWb2rSBMwDdztxNsg
2qq88l24QNUdOCBMq2d7B3Aabxh5xNEvrfLS7b0zHcxXdEzhCCtrbmlpiqaxvrMT
Lt+rdbXrRW8myMVL5pfR8pJP2coaP/+1B2I9EvRY7FP+H/Y8myW/5Nzlmdq0CoQS
boLaX/gf0RA5faqq34ktfhFBKmgaVY5mg2YZ/pOuOQVEOWXggcD+Wc7SGga+0LFK
RMKMydutZ+eM+LJf3iGrs1UyUXKbMMEWAwjhK0OPUs8pKoNViaNDadRFsk7ajN4H
`protect END_PROTECTED
