`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0AJyxu0Krj3525kvsusWtfWJE6ArvKmjlP0hc05L8QQQpoFv5VjD1ThPw4c3C6NT
BrtkfDGsNZuCZ3w7k7HZLxc3V+wPCEQ06TkTuj34oD8EfaAVlMKXKQSYZlWVjPWi
d5COaXPqM85P/fuqBuhFZLXg2QnO/p+gy92jfJoANVx/EuzvrvTpApgNKHN/67s7
RGx3tf6FkQmDXIFNtq4ogZWiodkrjZo7cVsetwKOuVscSCadAsd8XKB13Zzs51UZ
9mQvZr0q7eoCNi3dfbpE0XI+MgoiNeKFJXnF8UFVEYPJBojwJ6e24elOP9XKzA8V
s1WzU5K7Jvo0Bo1Esx5ODINI4NwTjDTHOx4AltEofsXm1TROfHKq3Ail6tZI+EeC
LQqCgRt09mr4tW/cU0c7OlkL0FpT2mhJiCNundyucJRVPuilkc5dX8z3kRANW0sz
CYdA8LH+m0B4bgCpvCpAUA5zjDlBTSq3gKNwmpso9naY+iwZsLy2y8BpLmCYhIPq
`protect END_PROTECTED
