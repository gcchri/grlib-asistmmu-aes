`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
an2OlO9qrWsI0XA54so6hl3wmR8V4qGclv3Wh5ZtyZsNDvZh/V7y2D9ihsR15KZJ
cjcSjIKZ7IW3bk/dWCFxX4g1EPh9U2mV9e1dL1oy7RkZjaGI7ek932dg1RSX3ok0
tY4StRKm1/tnDv2HerfSKMbHnYrAj0VtlmIYkS5ItGt5EE1+mb09jr5K8gbcJ3zr
JzUKanoUGt2cr/HU0U3Ms54hqIgcqGBzVtW4ajTN4c/bp8MGOHVa0vmAoL5ROhpl
wfLHNNM6xbiOhQEbX7r1lwgmaiVaF4sw9wao4fnX4ovynVNgcpTKCAiATglG5C5C
mKBPwg3wo539Q4b1Ldb7ot/o4zT41BBycUAJPP+G3r7V1ZQEtHqsSETrvJCSs/za
PvpKwCXVxKv5oicwDkzxz3CpUEAdo3CMwFVsDzFDluz0YH73VYvgMpO/TRgdOnzZ
`protect END_PROTECTED
