`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y8SWeEzZQ6oOMI7uBNWT2AFXOKMUOIMHxHhx6cFW6Q+C8Uou8raoX/xW851kBXnC
PswT+vZofFLihhq6w0CmNfe1bpBVrGHu6WeYQldYxNU6bHWsRmhdrrEQoxU2ZEUs
9KKxCSoimSuzjrhpJncKTBLeaUGJgM1rkyMV+8hUxHUCfl4+Z/2JV7p/I5y6INZF
HvGADdNka0iZkt5OaqhVFDY5J3NIgj4aFhKe/ikFjJUjYctntROEPr0rp4Y8VX90
R78NESDyQe8EWU+YbfSAGA==
`protect END_PROTECTED
