`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TBGrRJYJj060KFuXxvTJLCOtEtW9vDkMskPNkKrYPDXI7xE4X+2ukyE4JXL7IpZ4
DJlvOI9Y3eCWv/ieUk0dant3eRTLLuMCjaTogd3b33lOdEHB44L6rWjsYQIxudeB
71ROMn78pjU5Uw0SeslQcaEaH6o5TEPwk0KfKyBdF+eaaQ9tw6a2OX8YYy4y0ebm
U83sJblmh2OmXIHjDsEL3BfVmSQQlAZ9AwhbxRaPeFLt/Q7RJ7u2IV776ChBWC26
NLbau4DV73kHYwOFvKY6unlSi/qsv0LDgd7jPocvSs7+McIO4Ou3wG4cNNNjhfCN
TCTvCab8KLaiivHOCGhN3GBvmnGh3vX4lbRwN+qJVUDmg6MkSoL7NDcUQ5T6WUwx
/pumCO4/dy/qqMaw8Fn7seIntrZ6Yv4suZjYeKOIU3LCnZqUtPfto+g3OQGd/Nod
ajUXbZkbgoQSAxWVAOONbqcNzr7XEMWO3+ZzpR+xICnRfI5uDOagx0Ork9DC/XjM
PsMGyGt0MRh3v0T4JtEH/L/gwv8RRpsQorFXeK4t+gDDpplklN9t6GlK1Xm4AEBm
Pfv5yuZIDQ12oixnQNJZ746WQgd1w1tGjazB1xtgLIATjNxsTKjiE46B9JNjO7q9
BptOY+HHMtRYoTsou45/8A==
`protect END_PROTECTED
