`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UXtDPGipkf+qg/6a+H425nf6YJhD+bJ2apAv6n+N04mj9WALV2YWH/nwTy/+jimo
4WrA6Kq3zwcIkXOzPytR/fmnZXy0uFXNa9Asb3F+HeRsvzDHQVQIKNXL1bNRK/dS
LUicWPBH9j6MR1EGMbdPuhi3icsGUb7+i/+wiWQ2MEjJLNvXjeFQiDU+jIMZZaOF
22ZIViMrv8w78Qn9NnIRpWfijIHHs5agL6MuBbqXzmcD/L8qDKQFWwdAshrYQBIl
FQSE1hkoZaGpLC97zjZfb18s9sAUnHZPDHJOPnwQMJt1fGHmeEnOue/qa4BKLRc9
gGs910a90zrLd1R+Hf5+XzLWWWYBpxxk+65xPAFCeHuMGwQaIaIkvF41gCXp2orU
WTX0/sYIcWvSadwe9UMyfwftMXhSyIq7u4BdBgOCVFKUSg0RYxQupgm6CbtrUPM2
+iQvy3SVHUi68PrGLZUNVt9qwoDPbJ6BiwK6PLta0hLrOeM2H8YZsfsmvTnehMsk
wKZS7N4YVmsbPbpiZNIA2bUWn1xdtpQ/2UaBCIQxwJ7KTtOFxBayxlFTCCJnhA15
ncVgjHQpRcgOAPBtU7JyrVv8T8DCVHKA4V0/NyoA1bh4zmpqaLoH8/EgURUfktvL
XE4G/KTPjWC5I9RSQKOXDetSozI+XxpvYdtnwftAJ45REnyej5qYat2yFr+jHaYJ
OAO1dQj19AAKxQRVhkdkkGgp/XQK/lAGvd0Ev6IvWpoRzTPgMqIJ/fpqelHzt0d3
fvLIUkuagiEKm26FLZyToxHvEV/8BcpIQhJZOQjh/Q4/oLyAAE+4GD9DK3V+W07I
L8BcnyEs1JhNx92TIn/6+N1MTesho0VVkJc2Vo4cksFF39QpQ5rls6QxsJaXcc7X
VbYmjzjUbqFoHrfeLOL6hG4GAGVe2UXsJqNbKIHkAbsNMmTHDB1533i3vOBCbWsI
KrmBapTdXOb3MMgJZcjhEntLyKN0fAV5VCx9oQsXgTuZihQJ1Rs3z4xpJCicu3Q8
JTd24OTvrLBAHnVZntjiOIUvrToJUnhQWV3RVfdRHnAp5mZ0pOxNNPgEncmtp/jz
WvG+gC1pwHI/+YvgtFW/QZMCMgrsbsNdijPrWPLdZcWAM5FEqSPEeichfW1T6JvD
iskjnAk7pkzG9oqyyOXrjcZ/C9zhaSWq8d3odl2hwf/i5exXJjvhl2pruxa/jtlA
SExj44qYQYKWZy704x/Ev6w2Gd+SXKas7TJikw1wgSrIxZSb/EFJCsod40iv9l3R
mnuxpEQcwT/m+71RXRMqEaiCz9MDOfTNw/ALasbJeX51VGLcGOQDXt1NKLseLic9
kdq15OtWAVDZttVS+UP0Lp5KVmfxdAyB6QdT2y0FD0UrsPlpAq3t1xwm15IUEtJn
umd0Zs2yDvQ+zMC1Wn0XoWMUsK2jFpKK2lyrCO2VHF1QoVvVdx8Iit6G9CcqpMWH
x3+YZsaKNKukPZGsLNByjqBKSn3OlEyYuDcbQAqXv+jeIAlDbP0w7ky2PLPgYe3i
3gvgKnVXc8a5mo28IZhGJhfyKgBl4PINkkCjm03dfm6Ol1UnxdyF+wypa5doFMdT
O+OInv7QMCrVyQNer+IrsvATDoXaQDKW1dm+5IDPdJ7z+Xi09ah9DuJL/DSWBa6h
kqUFrdIUJd4wWn3j7r0U00fk36gO/UxFDKNQlGMfRWU/zTPMv8cIPbmT1/XifOT+
m+bUl6LnAgYlYp+2aWwtpYeie3YY3akjYOZY79EtVTqJGrvuH0mlRosvXhLvSl8G
1LOCgBBgi+VkAZ4wj8vKznoHiUdCFodjUsU0wryS5FB35nudIiONbFEaR4O8O9XV
`protect END_PROTECTED
