`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiBCxkLRyDAswKKBpMD/dizDYMoMaape/ngthqH5S0l8XByU1AqPOBjdWCO49Mvd
YJlOlHatVeJGgSOnc4smGiVo+ANAckTZDiaVFJRyTue4P/egesgJlGUeroQCCr8x
LkG/8Ej/xLbLGYQ6VnEGEPt6T9j8uPhs3LDlGdYcYLMzo+EkvRxPu6Pl+jab7xMo
BDjX+tIUuZ/Nfm6/1kY8zRdGB9m/nCeAzqWBGN7pvs30H6njBt3Zvwwucovy1wX9
tPiCWyfaNXggR+8ntj9K7bdN6lvtLeaj7jr+nfep94ekuLgULJiTB+NfEVsWQp/q
ytE+bcsdovQYqkG/RfGPcNr9hoaFMcKs2vqh0hqrbmKpGAOgeKAdtRjo2AjKQeb+
IkmUEZCTfNGixlVb6Aiu7Q==
`protect END_PROTECTED
