`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XBn8Lliv59/gKSIQNRXA8y/gkJd+Wgcd/lKXl3CIplL6ds5eDXIj3SUlL0zVQTGf
nE0cX6lnHJ4c1xGqlpfuIG2ZGYtty8tXDJ80CxdV8Kvq+jc7eFX7oN8iXcWvhqpT
GQGYjt7C0ASxnCXDALXeuqmIiexHNBDnzf0V2pwmauoNr3pOhv43zXSpyFrmLNIb
ioiX4SY8Y3K8JXbB6QMXyeUF8WusvoK7dDu7tg17FZIoChQRnz88d86AjlxhbDU0
nHZHqF6C2X4LMikYDP261g==
`protect END_PROTECTED
