`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
be5BdpDzOMu7IqSmxbcrqa6/uVvfx2ig/W8QYyYxZHZJR67RNAXRt/Ttiwbmo64y
CedadsLa8+yGrOwdraTizN3Bt8HH3dBuIJoUHI5PCJv1o0v4waEXQr4iTGPUkmdT
kKzzQ+vhXT+8bhK9b5qb54diGL6QkY4mLg8aP5vKU4YYr+NBz+wgr6ioV8xOdfRj
zRvsfdzd2kcneqi2y5h/u+xjoBOMyXmaDWnFxGy/zQysSA9ZpLbKiV1twNP2m+qq
tnT4B5EUkr4e2CwpD1iDghUFfxR0kfakh79S5EgeebGN4VFj8izPKowt/b3dVs2/
zBeq8z/VRxcFWPzXtvek+yW5dOYco4o5XVjKK53rE+qBTe3DYJz30OMk+3uBz2oy
mvuksopIwMa9i8YaWrB1yG1535uTeLvcVcJAb0zu8hOD6oyWLz87I/YoTVjkFAR9
uEa2Iqj22xFOTOlJ6h78N/kIekI77kbNuWfuAeMtmEU58RQ4IYLSV/cUESq3X8UM
4EJWcIn+YFtXLhBq5KSDxEtFmbesAOG143akBeHrI0AxuE67SjnPmKMMtPpKdo+A
sHn1BzrQ346f799YTb0+7WsH/23d9Q+oMUCb6RocujMrVAlygDiqtd83uF14AgSY
LDfkH94uWtQorKLDlPDRH6z6xPesKunMl4plmRY7KslvArh5dK+NhCyJ5aGc9pAg
w+mKr/GaSzA/iMqsvzyjrZy3M+tKHsn6lb2UD5+2viffyZBQfLKzIgFVPFWUffQZ
1g2n5T+adM91RekUxnXtGXLIPGdk7tzRdo9QuVdZ00ziffwBFDFe4JDF25ZSY13o
96hDyJtAUkXfQrFpSc6lC2wplW1SWe8XpCZPPCgAl6gD/m67NEXOInNotx38q8Go
bQlODp2LcNzrldn7jQtGKQ1BqK3qRBHlMC61/3kA9OCMqqhdCc4gXwqPQPJRNmT/
`protect END_PROTECTED
