`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5My0yzop56A22wpMa13AQRVk/h5zvAIOUxzTeMp2TY5CqDU4eLGsktZW46bXYLjN
UOdsgahE4FvQ/PePfLOI4axm4Tu176OOn/OkLOaRpkP1lC424SPzGzDN8liJ8SvO
1VwM5kgsg3rq3ddR86aet9uyaONjBMkdXDkShlJyztcYSfhRugAzjygqlUrov+KP
qx6S4GXNGr4VMpG2PZ2ocxO8K+ozJu67FzgBSm/DrxcyqtbOkJ+U1SaRCyoWsIhW
uznK/WXlnxyfP7JKQQQfFvDYwC9zQvG8EXRZReLDBThU5E8VynRgjqnn1q5wB0cx
7J4fp1LmL9LWVrfKcwu+ZLrBDqvG1Wz2rd5FbtEuh3lZi3931RfbLQyOJCoNA8ZL
MVeTLhgiW8wJYFEKooOocw==
`protect END_PROTECTED
