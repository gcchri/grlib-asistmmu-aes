`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QxOLnnDB7CUZyCZvQYI0c3UCha3p+O052Y7HmgJvS/D9CJzI6J52oVqZEMGZxGof
dyUAShvSxuLnV8DNM6OpnybfGWZQTuntzEnJMPYhvacgLc/YJADCBdpp/HBe1I/g
3azuHo5F4vAFxzF6f79uJf74PCVOYIaHNdzMPHH7JtobIpIMycrLBVd7oksQXI9G
dXEEOZl+ZJcn9x5kT92lakwh3iVosHtTmlJwOTswuGCXgX/yddTF1X9Lk5gAOyzH
3R1GuEmOMfDGrge/or/A/IwvqZR46FZKo3HbXEZn4m8CZOdUgP+AKeWmPvpndGhR
283buV4h9VzF6g73yISfM/ARR/pq+NM1KFE3RHO2vhXMMZIgI6fTpOB8zE2T5wTT
6O9vvAmEpqF0crCWPAhVQeErLPp2iFkhrvfiiJbhj814pVIWRkshnWWOatWVDZSK
XsMBXe6RHq9Q5gU+rZr476+CaRxagNmpoEzNPVwnFgQ2YlfbTgthPHWZrUPBr1Rp
yVfcJf/kc4CV/UYbtwNdyJsGwwGvOJPO8Xgj+mqg1f6dQ6LJBDEfdvvMD1/tvzUH
HxD8YHJYaq8KGK6PADlR/Jer8JiUe0XhboJhl2N6eAv0GLOVaCvIzjtz+Jg8ksCZ
XCnmPVpsk/E2z4csLdgPxUHHYioteaChbO+GjrTdEsmUX7QRHIWx3uf+bhRSaBzB
blhlc4N+ewccJcctbH+rJpc9O0Nz3FQ9HGWWs4xXBk/95mgRBIYiNRZkzmY5Yf7S
oEu148gUpsthcQogUv+ytsLX52TomonqUAyG58eY3N5PllZLslhYvgjgmahco/tc
riiOvm+o/fQY61akZXMk5roUhIoKpchb2SENgMI/D4cncRhiQndmsE9UYqL3wuJt
U91k8TgAObwMhxOhrl52NkQEADGQGSxvqPOkwGlKWwHmF2v5Yrh4eCaR5XwqgEpi
qXEtL6pAhd5oAV+yka9REEYp/yndpHV6cvd8Y48yfttyeGH967tcqPSuTgIGN37g
OLR8MRC7T1JDm/jz6wOw8e2XJwaeDRaM1NcxG5yZlv+G53icadMk8nlexYVdbX/h
`protect END_PROTECTED
