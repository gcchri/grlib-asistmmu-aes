`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdi1NuvqAo9WVSKGAqituNzRvL+jLuLfA6vU59SWBv2DPNhv4TiZMMUlIQo6DFa/
bDcb5F9n2p+JsHEbTAjMxuXc1X7AZ/VCQfLJq2qc8NsExppcj0iEON6hVP+7EI9y
ZZYIRG5lC7KQ6mbQat5WseyitLbqlMfl4ALdauEelA1eP6O2ZhqImFBeSmAcVEEI
i3+hAglAS18DPM8+/18PK2WbAZBqLwKOAiT8vhbkkYd3/6ZrIPEMe//B8d9qBNjw
pHa3gAyVITGvSb/AEA7SdfuU/WKakvftl0wWvOvjMXfuqOGRlYeunaAHWqCA8wCJ
PrWkXrnJRPDBSml2/2EQmDsVuhZ/NOYAikyCAxtGCsrlSYC5DbWQdfepRX8FzC43
FJwJpnStIO5PNuEB4wynHA==
`protect END_PROTECTED
