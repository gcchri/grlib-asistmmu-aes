`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eGx13ahE3i6CqFDSCVXMI+lKpp+5bkr5S/R68UKm5NEN9RULCbk3RcPu0cKfxOi8
2Gb0MGHokrTlVcUxdGklnIpBr7qLe1Dm6qot0viyTOjNI+cpnRrEAcGRF7k5L9+w
TgOME/G5oP5i84CGLyU5EG7Stnz77CarnZoEbsxVpTKGiLdtK2FkJMS9PacSgcdV
mR4Lk++KFdjkzBL+dChBGx1JxZbR0S9D4L4IIxe6Pz+vZdf+3xOlaUNM/1jHRVYU
vwgESbyOuJGzMMqX6u5fHaGAERe5Q4ES8DFG/VDzs6xy64kJrqzd+c/uuCHQBWBr
lD6GeuVEu0tN3C2K+IjKeDqGDXIftXRsKMQdpxLiWLdf/Sj1F99gNG6EDG3Y48K/
pO0EHmfDQklGsGo1SdvRCMBpXXFjtrxbJv1dCxMX1b6WHC/nsVR0+avOC+wy5avZ
PmVhBILXxT5nK88WxjPOykpudn8HAAQU1tyH/w134KtKxzps11tOWmjUXN0YMTY+
`protect END_PROTECTED
