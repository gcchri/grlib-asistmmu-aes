`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1/OyL2LKd9Rq/uhJy81A3q2nVBEJSR48QBZB2KANW9DYs9+6jxNyBnXVCxuGy3F
wUuVoF7yBLX0/jtCI7SqXrwYcI3CPlbCXRO/URY2p1Uis0U++JLyXGEpOpTTpTqx
P0H+F51090SRRJGLG1E/JMtxPEQlfnkkk146ejwKyiod40ChxxL7SUv/YCsdTyMs
zEQStmBv+oogY1YqXKSZfE7hTS8NDcjKS7fzDbxVDV2upUcXrk8+yxkfifAi1PTz
P90SUQwly++ET50cRaFA9oJ4PEqWj+gVK7O95vGwBvoupIH5l6T7kaYaXwgoxeNi
YxLooLO/TrctFw1xR4ZVuO7MCnNam0wq9m3J0naLo6cDZEJrGyzrPlGRJ4iYL9U+
mOXkniQDgJybv1p+ywRFZ+a5lV7zFrFMRm6IwQ37dqbFfzWnhY4Z65Avthwf9KBL
nmJvlvCsJ//rfoxPsSIsjRFbTijsIUarPhj/Xms+M/+0C4PsrfHWCUnjwc5Vehi0
JJXvZ4SQA5hMQEFh55k/dlbCLufwLyD9fQs1/itLh9L8b8L/E8cDZm8lv887ZjVB
`protect END_PROTECTED
