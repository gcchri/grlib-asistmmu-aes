`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qBmFRraXKHpsotNfP5N02xAgb4bi1cbXQs0PdHkJz1jTQ58McJY/fsNmjh4AQEQm
7BegYcuXCoBTne+MoYWQ8iZD4HIyEfNpl7Hj9v2LigkC1xrw/mj0du4S2k1N2tjN
6qJekSBFajk/EFkUrcNH+zIAJ+yE9wHN0HoqZ2I3TntY6J/twQTod4hOdcoFNsuw
5gO9RbxaUCpLr9p2jBVMHWuqHg/PEygAX9otJ3czG61Oc1DrJq8UX3Mje5j5Hkei
3jcLv0keGtm0q3c3GpQ++pkau38lldOY/+6VW2Qqtkgf9uRGhRwJN3BiK7g8GMXA
tXGtm2uj6IqK5Ed3Vtum2dm4WYLZq+Rxx1Sw0x8LdmiMF00IFDcqWJudmy2glHMQ
TkQz+Ffbff4vwG2y6kTZMAgvHEy0NOmwevFdOyrXXVYCDbRlS23Hxnmwb2GfxioW
yjQ7rLOcpHbx1I5oG245HEY4Hfb577VGbkHN6OFUuzE5ye0qkpZue4LiGsZ8P6qW
cd2RKaZgyyomGAAy1WosaeSTBegYPB9nquogKqqzS3os1p8TrAk5eXO9fOC+0B03
BzxPk3l2Zan1yhlqYdroImUa0T+HrgnKrzOzSGSwZHOTliRxfXLcRNKkzeXbznwW
z5ACmBJclFpqp2eF6Yq52IXGckc5P+FTIasEMuuIRwuK6eXDYiLXPUMc3jiAsUm7
NTv+iIHNeBK72AFibUioBT1pnCb7t7qivEAWTKT1hQ17zuuEnqnqusGnqSkstYhl
ZYkVBzTMVmpJsbya9DYsR3gSQtYLqiH+XDnbondr0GB4JtYxfummYzSULDabYb6I
IF3jPnfRG7DNjI3bp6/DAw==
`protect END_PROTECTED
