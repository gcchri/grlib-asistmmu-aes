`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6s0uLAOdsV3sK7+Hyu2hQUj7Pt5BL4UcYURxz81nBqhj23Jc2z/GZ7e5aO6CIIzD
v9CCjN6HNPLnuaAuGwVGwyu2Hu+ibU3Aw5DEhDalCi+X7Vt9q7KrBWWPJRBy/sLK
qOU+zWcXzRJs/3QWkXP+APy/MTTgZimXDiuUbA0tdvTg4kZid0U9K50WJ1PdmxyX
NuZePav3Z590IypKTQI6zSd6Q+p+ZMPZ9irFupuH7ZcTkWqOP+wrf4f1Qbn+2FdG
JYU9RxaDZQjuvnOppZOqq7ULNzDn8xwDCv8Ya65RInnq/KZh/oDEVlCjcJ+AfiD4
EgCM4N3MqpWzjQmfg2LLpA==
`protect END_PROTECTED
