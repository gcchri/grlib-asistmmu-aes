`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yu4DdAUI2xTSwi4EZC++U5T8HkrA1JMSb/ioWAt9WqvQ60pvZYu+vHHFLpYvRJlS
o3Lc91fMYeyhritbjFwSZuz/bTh9wIvFUkSdGCd5gondoSDjy/oiYb8WvBxvVogU
g9hQDt4AFhJvKmi5bN5Udbyp1bH1JnNvMbaFk2eh20TbPnKLKHJXpYftJ1BAo52S
hcBIyAx1v/a9nALMcP0zg2VBQBgnpy8vzgU32mZ2i6+PVtW/zrHosh7KSbAhP8Ds
olqqoTn/dYQtR5sD8h7hA/2JMfyRc2c6bLaTZRneTdZxZb1uKYPFFDnQ2JvoOfoJ
PfZxPP9dvE3/iy1+ufsP4Vo/3oB0IudmXfGijK80+SstSk7okm1V7q36AakSPPCv
n9uATwEfV6eDiGnFaYOrTIN0RPcutNwEgqBtrtoZM+2CgTlo2A5zKMXt8MMXMjpI
ZULuQstzzTTSpYdDokbqEC8OTwxzmOb0VGQRZ8Ku8xmJ4NYnqkxuMl0b13zmZYbg
etDQSjFDtO5wWO5mCvepxhT825aonwf0h7NsYHGerSyYu9CcSzmUT4ZdPzXFmO/f
54LY6yGjidU9hvkryPu9QICRz9ce3PRFXWPQtSqBM0cg6Dv3skrgGc0IgUeVAzBE
7/gtSVY4eP2K9AHX9y/gVtFtXpuEFsYcX+Ga/R81KAY=
`protect END_PROTECTED
