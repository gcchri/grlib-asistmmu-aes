`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BePO9oIyql8nFqcCxcjZjhIVDVpEsrvgiURQxbzbRQLSjKkJa4VBE4+3gNq9wao3
kSpnR1MiZWJdQ2YtGF5v20dnbHBv8h3QZXmdZdcc1kAyxAnlffOMH9BldL7hxRu2
Dj6ftFjUJacqlhV4nNVnS/uI1qU2t1Bd1JWu2otR1maxJD5eiTxzK2+7E8BZwfk5
m0TMvhw8L9/5NVwfhaGshZAy5lHYbxydW6YcD7caK+2sBfMyiQ/Dx8Z0RsDmOV2J
/XkQDzeKu7uXojRcsRaBZ4xDA/aBRohezb00wQh2ON4LtpY7XGPV5jfHt+jgOaNF
a+SzDYnDJ8CZ478uXhaOVOpSfhpLwUwq+IZHesqtq9MelaGnmj9ccUBNRFOOgFHq
u1sBOY8Ud/tO1pFQMZot7MQ5tGZgh+yZPggwBV2G2hKVIElngJGkLNP1sY+UMNYC
nBaRpR6Eo4H/xEiAtwTF1JOYzk0W+B9cQiLjzEPfh3OWYeucaHNYX1WeLfGOisSp
Oy+7/qBl+sKK6XyVh/Oxv0iqScxVCbCV0Ogiqb+QjfDq+uqJij4qCLtqZtXYMJFL
a1fqrI7lvwrwcV2koQDazneijbexXHQTMj7qavHMrmuhUE/BX9+TJuDdUFhBFto4
cclaxizkytjpMb6A8ID+GtCObMv06665mQP8LFSNAlypHgAOCQMd0avQc7md4lZ6
yDMt4NOYVi0YCxoqg1FiT5yfL4MHLPVA7LHAgSpysog6b6oiKylm88cQaKraRUv4
+O6KaiJGQuN9NbMDaS0x24Lczr2W8obnNzWoYqNQnkAMMLMZsKnK+RqCx0CzZIJf
S9bl3TXrCYuUduIcIa3W2iaVOgjNumlvSaxKOiCHIvgDHRo+tKjLaABe8MTzF456
mts8xImPGyIT8KGFhabFSbJ21ulMnC95RL8ebfwhki4Fb34dfpmJFOyb2AM/bo+M
/FEs83n1YOueXw1Q7QzFpsOSCQnjNAceSaaLVAvJqkvs6zbo0ce78RzP+fMXySNi
`protect END_PROTECTED
