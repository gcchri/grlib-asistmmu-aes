`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnvaBg77DdfgluljP5lIt36AD34cH/WE8UsDmW1tFZ1+kxletN72O3x1q3Qt+kix
Pj1He6LmcLCaoFVA7BWnF6uLfe+wwYesAUgHayVS49LWfSSSvGI8Z/hCVaO3+qGY
yJDLg3iUMIJePUYqdraDL3SXL7gTv1802zo/x32TRJysaT6GpBrMu0bz4kUPDiwM
Roap6usqA6GgYeRWugRKIty0myI5NXtsD2xD611OqeqrARTrXMHm1+3lWlBmmb7f
FlkMn0QUZZtg1PNsuFH7d13G0XEKHCbkZm86Pp5UY+IGm6tfJ685Sy0Yyw9pgS0E
il7dWRqQmboABxogC6r9ZsFIW92t4B7w0oLU/twuAEmuDjsM2bIh8LVJFMTee0TM
uKWd2rwZCXKfbylVOd181OYhTr3Kff74Ljk2+jf9KRTVC6t/tS7s8IGyEXMBa53a
YjvCee9GRkFqxneLWMBmiTc8RD+dcwVTR4Z1gVg2in+8OS3/NP22lewWjzDhdSgD
yRU6lTch14yR/ISjotffS90+xq8o17qOfOPJAaEeaa/lQcHykZqbBy2cgG2jco0T
FQzMUCZGXqmBE8HRQO9/LPpOx6WxhDnDMwo2LKwxix/+H3edKUwBobQ4BMOGIESZ
WkBlJFXo11/aa8XSy552Ww==
`protect END_PROTECTED
