`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xlGEwpPKOsAyhLZdZLVnXE10X6u7Lf/KM1on6PNojzTbIrk4+ZDOp1hGHC8WAWEQ
LjfWbwcOtCqcDML3MghqvCSlbbMKbeZNpxOJGz4emjLhZwcNMnQnwXixiZAAUS9k
g6y0VF+PT86fsod/eW/XhQXMdDPYrAZySc3zO4CGBvhUl1JHjd10gYfF0M6tXBKf
Qk3sWkuxS5IyZbnwGHKURavREzszxW7Nm7IZ7kmDhXeHgCkn88wLwUe/agxUJHu8
A+kahPb860SifldVsrGW6+sm6HMBNR3MvV+KZt3x03EtmyF9QWa7R2lG4CtfTs2I
RAc0pQo08ykUrQ153fsJ6H9g26ggDhUlN/eD6V5UvAd9D1HbmJEX4tzB7wMW5NA8
PvEK24gGXZscHmfPFVMg6/h4YjfNk+hAbnd2GP6/xPlncyLUCbHLo+EzVxsrHsIW
2OqKJ0CnPODThK+DtVlUkV3SxP8pGnInshlxpuGUZtfq7VoWlGcL0OVIILczs7F/
W3J5Vx0sFP7Ymx4/TEgXAlsoq/aFU/suSS208PS8CUTkoJlDe5SUnZ7oXTAul9nR
Aw9OVqSzQlktlCuSOhA6aC4fAZGqd2vf9qi+6OXnQvF1ODlaZjDusq6PY9zT6+9p
bu+LDfNDRws4uVklLwmq5JKVl2e41YEcrKq9xm1Hg6sptDu7k4yTTTDe21fhaOuX
gPZD7RqI6s7n9/rZHqK3PqgqWWzisOoLl1laheB9Kx+vRwcN91ohBxJvD1I2WopB
Lme6P3/wjWenyNtG5WT0G5oLYYS3WfDZou7ZM3FEypsUZSlMthYSnZKShaBg3fRm
RNqLYcJslwd2CEsrmXVjZ3MuZDRAE6jPGMfEhBAACcnAMAqBfKL1VoWbDhZ86IW7
IRRLeV8cdPVWoFiCXAI6+jfGtKd98bu9YcqgHoYa6jc4uEKRLJhS9TpFAHlXjh2B
tB1IaNXwngEZZ2KTOi6ioCONGGjLavNMhSUhIMUkU5G8wTcxHwXfZJXXloNQIaB8
KttNMf5M3v288cwbeg2Tp1T++g7C1OmWJ3cT55sUBhZE2xLficamLEJIzixbV+NP
hInNvoQb0WaoHQj9wObVMHH0dxaovyHUa1i91HoeztsbVKWXx8rNiOgbbNTf1V00
F4hWNC+IeH+nTwrrOvnhkQThfCCsd7iXKVUl0I9DtxnnKTlwX24ZixjjLFeifrx5
Q0w4o0yoV8/SvQ4REj5/V8VlfYPS+Gm0HeQxHf4pF/pHTnzR+nAAxTEg7VGOh7iV
JcceWzUm0+/LdK3Ul6pDtD1BIOMGKp7tq2PpnaDmV1KK5XfrDw453vPCfS5iNirM
ppA2K5jkr12zU/eoiE09jv4p03njUnq3p8iSmENAVe6JcMn3jfBPE+rAbjWj/VuI
pC1/MpF0sIHBdt8UwVuJOdAgDOEKgraQTLf5om0W16mpBL7fD+u6mvtjp4l1rjke
6LgQh+EqCEM5FqD+Qb0HDPidAs+5YQDkdaK5UqoNLqw4httglEelkBCX4sStlm68
5tcRHzcA9r8+igsYGJ5R77L297BwzOjK85sG3UKN4VEqZi47TjZO4FZon5/+2J8z
BZIQwt5RkSDCsPHOkRsoA77+8tMB1Gb7+EqZuwXuwb2Z/jkBGTp6W5VdZrB1EzjD
H0oHUamMwC/bTTADvt7fvfTbbLNUWqy8E4fghycwH3pXSAAYsj3YyI/Ckbi2lW4T
XyiDOybK9OZlc3rKowG7YEHehRtXDXQlWQmv8Un+zh6J3iM/mLAkhedOh2iUH2j+
fEHajLPbvIh8KxYEdiKhJJC7Rqum2ufgPFuLUxKXJlEZ/92A6+FiPH0knCnfZpwd
4wF47/ZQxDVcx9TkyHg+xB42xIfXjwBXjPIsK2hsM/+A1gHxbHiZ3+X7dg0/la4w
yp+YtBywqunHrs2gDnzRp6LWawVi5PFnodcMKFsuGciDOQr61T3o6t0T6oU8FBBq
T51OXDnVFpA9jGB8i48P6UiHHncKXW54Z6MNTGIHPgHsInf5LDZfFEH1pEl+vgaP
G+gVGmzzPA8ZPg9KH3ALLQ==
`protect END_PROTECTED
