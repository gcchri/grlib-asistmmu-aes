`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tqE4rPF7V1RDzSV+uniYL2X7FLedgNX6uXMmxioysPa/PPx5j+VQ3yKpkQzmS2un
Mk1JEi1UrjAtLSFPIE7M7VLIvfsfhgVAmw/gjDig9Xg1tjclGCUPQIXRuBFzgDmr
zkY/fjbGP7PFrCtTCpSPGwpFyFiK8O9IjPLV6m3w/qc+sIymtZjmJ/1ia+kF3Mvb
oMkPRkkSezAR60hSJLxEkCLabF5IvnlTvPHQH+oJXNqfW9r7ct4WVU7M6bS8kT1E
+zn+VN7N7s8OI4pND7J7G6peIkxOT/5tOUOc4dDlypkocah8QKHeUjwEDbIKcNrI
n6hfu4fFHF/zru709agF/hHmAPNF1GP4svyr2d4u4KTH8GBqdlyCbdgKiUk1CBON
wsrIDtFtgnQdJJvtNWtZi7nVhmD2bGZ/2v7NOh8Rt1Dp9wHXe55L3oOolubRj25N
LceXQrE0TTn2dg7Pm5HqBAkL71xbziAxnCmaSJLZRgwCgXtlsQ+erq8+ZsrSJbrU
b7pPtS7tSQXTAuTxG0eihdYXx3DRhI/srMAvlSqU0crcBu8ZZNDKrR0xwJJhLaJo
uWJvlumB5v5TwZtUNyIO3hB/KEoBun+jOwTsjUTpN9NMdvTZ59hymJGNenORO4vC
BhDoSXvJs0toiL2v3t6qoVbQRSsrQfBoX4oJl3Z7B6ggYKkm6TpV/TZZ5FY9PLm+
M04hQFBelOoT/4BY+Nqj93LC0udVDLfr9pTqR0oZJtI=
`protect END_PROTECTED
