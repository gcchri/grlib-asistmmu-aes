`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4w51RUFxFbMAcIzbGRLOqdzxHJAwLjTRGIQcsYgrpc6ok201nxbxZTfXxdDAJ0Q
w2dON9w4iZT/goM4ykf6WfGSNTfJvGwXwvopYEtNQ9cdMKzVVBdU1Zl7pKXvyMZW
GlWAF5MR+sfW+SsteUG9YMkv77hZw19t6TlRo4ceJsfspEZXchK/xA6zCh5GsFPv
I/MA1rJ9IovZJOufQrWJTxlph7JIUKlyu/Px2S1g8qkT1368RUi0tPr4U7Qyznx4
fjzetc6yclVC6wdN/QDVt0wYvgk7S0t8BAQiBpyoEsIt7E5F8v78zLif+bYFuLRF
I4gdM5FRV4+iNkWMWtpI6fWN9rYEC7MKm8/AFU5fQ95wolYugvqMmygmREZO8WYX
/aPyNXqSSbNHrPsI02t4gnqm3c17I8wS2oRWZSM6xKs=
`protect END_PROTECTED
