`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZjS41BaoqYj5sjXqcLWAYrVYH4An6cV1Bjng0HHJkR+HeS/66BC2bW9kEq3RPT8q
CSica5lFacJT1Ykb+Gv/4/NtmnRJc+pSWec+wP2FkdzVy/w2eshsHdLoSj2XDdQF
WAd2cMIXe/yU+QiOQMxoEtEkhfa+Ww/ccUo+Y0vQvizcPFGL0MeY99wJJoQoQ6YH
imSzuYVFAoE1ENmXkMQD5WoQyKrW9L57nI5DP5R90lkJL6vUafmRces9W/GvbIND
VUgk0oK7DF7Px6Gw+q9lp159C8h+OFOLs8+B/Psr1hqaZahRLNtrEn5Cox3SHHgW
xNCxyghF8Yw56dR9I4g8pW76RTi3gts4v/FXyRjCerC6CjwMf6JPYc8VU6hbQ2o+
YljVIG/B/llJPAcTeeXLGKl94frA1uK9VZuONs6CGS4=
`protect END_PROTECTED
