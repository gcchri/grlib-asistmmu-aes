`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CM9ORH3VQIOFvnD98Hdre/fwODUJlNKc5Rx+7XiXqvvs9YKoOSjq8Th08+5MAjVk
1ImxFhQxw+fEXWXeFpkGNs7fI/x4GSaoLuUrJIWxOS+1JON+R5+h5d5wJEnY7jCb
5sEJ0wAf8nguO2DQj8zu50U/jIgVq2NPDKdg31GQ5du55Uu/Ojf5jBTwaj4Tg6E2
EouKjcP+gyHwz19PIN6pC1MbwBcXBLwe5unIMdqEozTbaPkEK9N8K7QN4b8oikqh
AzRFonqbIjD/kPypkUkgb7iHkJxrlQ5OL1hsI9qO0TnJrucm8cwnXlq0HOGPfYKQ
4QWjQKH73MiI+nsrUOjKLrKL5VQkADh/ssYsvIe9bGQl+2CH2IJmuDlmdM2nZvK6
eb1T6a3gauJhuEG8W2Fez88sgD6CHytEfgrckZ0UDYQ/Bf4miAEyV2bQP7GrHA2h
rTsFxvpMArjxEZDdlxEOHdigbFk2r+4HDDHBiD8CSiUg0o0pOrPhl3sWVJ27MciV
w6OYcWJBwz6tQTT2wayoSAFpbbsdbxKSy9r0KgC5YsIaynmVgKN9qpfI/ojrIWRj
nOJMaQqGLZ8ldy43vmxh8Msu3+Tvuohx3YkURFzwzV4N/gBgQc/iqPMXWrm8F5ng
ETtv+BLkUy6P1n/wdvwSiLxGmMxff/C8p4JFSf+3Jvlxxh4X+mA4EixxPXZaXMop
KGJqfnyrii9JFE1OL8qUNZgxO/joCmHfduBXGcsRAjsg55L8NPLnrPeT1Ibe+lKl
FXluJZKVBfOrSqoR/aQQs8BVMqYIECuUfujOgmCXW3I50hU9yNdBMmv4/fiZVkpr
W4bam1ydx49/Mmu2rJSM9r+MTpDePjDpiMRFUmeP2B6wM6sBXu4XFi5iX1ZvsPd7
ZG+YHNXZ14u5WCLLgIFEpCpQpBJqM4CFVMC2Dfsq4mwnSYfCfVXf1wRyZ2KcoZ9L
kdoPvPLmcx3lLrpTrmMTQEOy8QeW3WPeflG0Yy+tmpgRk30OPsiCbEvFS/ZAdM+C
HL83FU4VOj1ot+a0ZhwLkvPCremoA1KM5EoySMIMAKjk5w3jdWWE7WD6gxf80zau
rhS3Jont6DtMMalLMywz0UzsRmHp0uY2s+60ezzGFb4EUPxbRQUQ8dAZe9rS0fyq
u/jyfuMBrinp68gZttSFn6gggoFe3twvK/DcAWNKiaw6Madf9bps0aub224Qawpa
XOw2J80YUfc/cTd7xofttImA+nL7dIcP0IOKuegUZX1VhJ3bUTL7ckhkQPjUNteg
jvALFP2g0ONrrcxLi6CeshYpvj6KrhZvhgCon+ulmRB7uhLUWnKkli32KqppVueZ
hOZTJGJBYOZr1Sfg9WseBgKoz2M6MYgo3524AL6nvQ/0krfs4ymUdLxBBKLBxbUe
Bc+VBn4XgcSrNbLKocnIvaqE3pK2/ZT+5V1FSQNHKrQ9LiQP3K17f3x89npt4ibL
yynqs0S2OHjsbMFlOrcb2cLrSnAellbDY3sVr6r2ZvUlwpROvRLEeLofN9MKH5a5
h7vMPayTgTtx/y01WPiGwMA8u4Lycdvzts9TVwISB4yDeX6zjrO7XiBheUkcfLKC
RNhImqASwW2Tl18TavKAcX89LSwwMTZXqDKENXNIhTrarYA9RsM2djG67c5XkLdy
khoFpDR2J+YagsZJ3Qe+tkOHAhb6Meszw7gtLQE9EYwKA8ZI3EPymwvPknUTFrRS
VRA9IOL+/7XzSzveQ8fLZJsFjqcpm8dCGvFIhN7lQ9tyDDKd71TXYQopF/PmlEKL
kSSjm2lbr/t30uBy4gsa2alXUNC1x46R4/B0kL7p+phlEtydSSRTQulV6yID9YiT
d8OVrWgokWZxCMTlDZyE9w==
`protect END_PROTECTED
