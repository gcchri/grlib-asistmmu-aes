`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxdfcZkHB6e75szfeUNNI0D2EplCD7BqSW3qFTpNNmpaeWc1mWn+TRtM7m7a+d6Q
jOIe0aekNf6oehbk2lPfKaVBfYNrYHTTxyWJkBO+etgGZmdxnrhU+abhmXmsB1Zu
ckuZRYzROChnxKJtLMJoExqteBxwB3flk1NaCLyfZjVX+6YJfAjsay3jd5FT1IZN
93zMkpdMHg4RD16a13TDrEWy7CKlY+YDSUNkxG4AelhNnYiO5MjMwScTgIkcQzw5
QBV8wl0JwdyhB+tz1kl0c3iq24zFsLX8myvFYbnyKwY7xy5XWgtqUupdDj9ZaElW
T9wy2h5R2LJKeZvvsVncBFg5prv7hos/ZSKoKW1YrgrGP8SxghtfFkPZh/QvWLxm
kNY+dborb1dbdseaOK8np0QDqGnXIgfupeuF4RuG2nK06eiCPjRVmBTMUgMpUOAF
RM7RhwIYIKXvbclYU+on6dpTKKIBwCUkJla/5Tyuu6BUaSoax951guDsfHmecWxP
vmNqaGO1++Jj+W/Q+ZXixkZezgcFV8R/eBjJyrh4HrzG+M7z7sCoDB/ljNXBO6cw
dx8hmtPBQMKtG1E+VlFL7djFX+LPB10rPz/OKxs/RDrZHnLqcVslfMSpPt8/4wQW
K0m94e6GfUd76y3FKeISRkuvW9DKwm5iUy4EWKJsaw8NLr/+06yUFJzG0xOvgSVs
1yLODPsP1JcgIfTB4y1bNMXhtWrBTYg7UZazes22QSMag+nehvFsLgIS53I5NP23
ezsCPQQKPRsOEUbug8qWgQ9SRYbKoU1kwObWbUR0c9M7qJAVMJ1NUZA3CJ2AjTVZ
IsIvr38nompJJB/ofjCM6g5ElKcZBYI303kicZYNrhqp9h3toR5CRcOBzKEbOJcm
NQGdWKwetUzj+N3dSjtMfvuFIbyKXdov213DWBq5i22TF4s1kU8GEfrdcdpm7BmA
gr72YPKCpguhawoUxSave6PNGKEq+6/QX6HXSQ8f0x6UqtIkOm2lrMTFJTG0xRKT
C4bG3sV1lJWLfIJzLWKCYpMbonAwqIbeN7sjpdTSgLenBpQ61hZ1bf8LLpTIOtps
57YQ4BRG3FYDDULLMMn7yPtIZrlf3u6WHr0XatN9jZyWlAMMIUp5opvId0TndHy/
qSRNki7WkHPTC32s3whf6gBgCnbU0SoahKhquPhcNzfk0tx3hEeezWmpF+5sdRsz
mprF6tHx2ehexoiyYhAqFXbrhJ+fXho2iqX7BL1mcJJM7swY2A69yxnlLqBCAbqJ
XZANE7JBKQizOPTjrmWa+w==
`protect END_PROTECTED
