`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zvep6btqsp8Ke74XEuZdE8lUyKHyfu9jhfH+6vkistsELEcQ/23o7otjKmd8BTEx
GDlvYZOmz83vYP7GElTG3XjPwVXYTcizzqFkPAug9D0iKNxaXHDY6lJb8lsDUKKc
BJ2pnpZng7lBcrJ3sreRrbQVMeardRase4WYymY00SnzRkRAwNd0PFK1oqZqUgF8
GQDVkq1n/BZlE3jWgJBPs8OCBEl3ozf02m/KJlcL95Fdwwpv7ZhNtQiMCw9R5kbt
iIFQzb3TCUcAP1I90pZvSiWBbybpusXLUZIWJnNodiY/bpoVW/tT+DI0PhcuVK5v
Eq1Bn4Vf03FDJGw6tcGXvrzlVB+x/anFDp1UNwLRf6dYwhjWYamrosC5T9exV44D
Z4SjOV0tZMxnyC8M7KJEfPioHs/p0EBozxeqZH00aB0BoFuvK5rnRU0rpC6FiTS4
imiqNQybUKq2znfR+vo1dRKJjXIA8Ng0CEJt/Wl5kzvX/g0AqQweyrqYHV/wr0iM
Ob1xmznjvR+0lExKl+NWPCPxfwR/+gtmhUgft8oAA2YfvSfN/yAwjkcCFnEtblEl
VL4Djw9OFQBekmfeIT9oHzDdkNhyzcTkMxFssB0VDMuVYratk9iwaMBQXX3nuJNK
KmBJwJ5r1B4sqk4z1I2oCAq8ZwOQjMEtieQfQjAgigTmL0Kd7PCa0d9w7Jy4wCUy
/WlMmk6+VcR9pO5bJ1T+CSfbijWduPw0C2vkJ2pLAbeF4clc3fqAaRYgH8we25/e
OkXwAPsywvwSvEZKLFykzBLPhbafr28LNxz3zbNkDuQmmrkoKtlQXIu8q4W4lZMm
9nMYsK+2r+NX0wUtXpbQClTsTQ4twIxetFjzZ23/zYDe5FDJ2qdHmW2YD96T36D2
4F4c2DaSvhb7ljwKPVFDyg==
`protect END_PROTECTED
