`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CRO9ou2psEO89WmPu3R+3/QSpkBhFAJ2lW7sJkFlTjGna1J/FlCzWDT5URQB2JZ6
WMnkFlOCkVKi4zLxtyGd8bXxm0WojMEZFBaLpH5BJk/B+0v/2rAh05xUhLqPYCWd
rgIcShE5IJauxzMqU4nOlC6O43teSe/VBVHBdSBeLJMSGLVXDco+uzi8AuRiVyaI
1OUrISmj1QgO9XC8LwhSFhYJOeKtclt8jqI4Gi4ZSOzS9ms1y7kEBKyta/1YG6Od
YnE+e9wahGRGMOgsuOWWOCvIUzpZzQLNfKTddP08MpglHWB9m9xcH9h3U/0TkHkd
XOEDV0rLOUzSUvim3rz4VgpcMIAT+N1+BgzmnhKVWvxHEIR3E9pRLXSKEBkotWvw
o3dILpMth4Kia7/E4boMVMqcknhEtYZe34Jhpj4NBZEi38jQxe2ETiW8hBfhxvQx
`protect END_PROTECTED
