`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1G2xn9LwI/2QaqY5gtFCCMCh24c4IYv19ON9K+LF16ellgDhWRACMPvu4zazTkEu
tnRT6FVDfFZkPQxCDErZC29sJXg066iHKfIjPkdlSHjNzbejz15Z10set9XEfM4p
U2P38HB8jwErBG2rUXKOS29K9uk93U1J7cYEOORJN+HsiFrUZyjR/ARs/xxrQAWr
TIJGurc2664cDZ6EafOStFqtLWJFpGfDnBcibIhd1k3LS0PPuJdPTYPIV5RdUFDE
1v/BQJgjikL+ZCgRCXEGa9sGUE+2ChW8XP68ZTOCgRpaoP0mWwHY+IgBNEMRCXq/
ZVAIaeYjaU61KVeqI4RzyPvUvpol8lE/knUOZEOXVyXXVm1uX1hZXbcL5NHnwe1j
4flHCwES+96kupAntVThEnWVCRY2vojJPgVFzn2E15XtIMtbB/lDz9ENc1JiGgJj
XNsDQ2U5hqyZhPl/9muuBeYuN+eeO1AbVZ13lxy3BPMU+MsVgfY2O7YygYv0cziH
DpQZ8hDqbZdmia/wqfauxPHB+CGFXmWqG+9S8hA/ZhyAqH73gnHLvnoCqlbcGYpL
4VqxxCCEHFHk8o51rXtIWOEDkDK+E3zHL1616fCN9RpDYzGEGkjWDXD6UZdME+q9
PpPpDbx/N2xvDoCjSF1qD7lPSNNp75Yszu6MIYqHgA3wQZFj23jaatFtFXAGB/4S
1ovhRRG1h4uFbTyd3361k/qWR6hcwU98UgP0HcMBH3nKe0Xju//K4lNB2XXnCe5J
r4yhY0PGf63xdVBRo85fUIW+Q6FHhd9zvWiiXU0G2ZDsSDBhzZoPcL6UAR39GiFt
ODby/ISvLS1lCWrNCshhL2l+NM2jDHkv2i2BFhWAM+GYSd6/sbNZyb5EYuY3keby
5tyobUVBciXcb/bFmwD1XaLYdOwEtBt02qvAGcSi3ydULNJRTOPOr0XkWgRFlkG0
irUD82i9Gq5Q+NYINDIkeqr7izSZrJ4GXS+nx5iEd7QHVZkAOH/NrP86+sHx75kK
nmwv9iaLgy32DexveNbRxy5gO9l7LvHzvokMXbYLSB7A9BEaVCrRmpc7AGm4Bnch
DY5VL1zbea6gHcTToNVeTm/H7jFLTZ18Wiq6HroTVZERrk5oGbA8iAhqdmgazV8j
wddcWVdiPVpTBsXVK79MqO0aaVix9LBsoJBm6bnnUssFwwIBfEB4wbhfIbkuGOFG
drZ671s5+bUfLje8j9D4snv9avInkygujmuVyTqTK1A5tt4VoBUdHBTmPS8j8/PP
DRF6/E8Jj5AdfUpeD02B8WT2OniCGdAEta0Pc3/8HfeqsraKMeRF/cWGSG2w/gfC
8OnVWbf9yoVoQb6zrHserKm0hPVBartMMPVF4OqDHt3WuFxfPSBj9qBWlmKjYpUf
/RfQpM8jr5l882zvA+ierkybgPLiKd50OKhsKyfrHrsiZol3or1NnR8df07RXSym
Y/7fWlWODmTUuP5wLQYQtVd1xy3OSHdScYVigTtkOXY3eK2OW6UFEwIGS5tpOWCt
DxoDamAI3nJHNKfcqYdzIZMK/Sxn4g6mszNwO9RN31g3qaY8dREp7szq33/myM7i
/dwzXWxFYF+KjPr4B9udhMUUNIcxUEpgYGX/qaDb/D6znSVRPEboiJBQ7ls4eSW3
WtmXQ9j53MgUBV9b1Te2Qb5S+0XxT1Lpjf6s97mREzrW5BQ7s74i8NeMZTfn7CDL
G/vp1Z9lK/KdkFZTjmbLryfnjY6EF4wmHDVAWGjAslxKy3NlwNs2XqhAxxCeQFw2
vHlNdCwQAE5iPep/hjE9vbIiy9Iejo2izcgeu9SsNdSBV4DekikNx1yOdE3SmCGV
iRubEHnvh9/wqtVYaaYCDs28rjgqAhxgdVQCRLitk2+SuJ1rRZ9CvgZAv/8nmzbV
CV+Pba+78QT6+1DoXpWoB5Jjk6lvFKu1QlZ2qZwFfuUbkH3Yw+O4qBC9Q2F7yi5L
O3mnxjCSznpvFlP4H3fByZWtHeX7yoc3R/lKr4RZDw3xCqBQBFPW7xJtdmPy8A5g
K9EKJ/SB7h/2WeuJvUjEkxUdvyEqv5/XktF8JfDx0EM3gj1S+sUzdG2vyiT1QHsW
dUsG9Bnutie7WsKW1dIGVpr3KWg4NXdXywMef4OM4OUrrXDp0+kP01wBnBEe5kQw
/fGhWqndzxK8Js+T+a31KEXVFobCQOh2pz6ZK8g8EaWYv1+C8uD8y06WHUAgvD77
ARkOxHtvkTaGPl8JQaBL8hMOON6kO55k6dRSZ+LwM0z4m5+1lPg5DQzmvNE/dp5M
DgWF+yQwTzyeuhyP/KHL4ue5XjEypfjCFYiT9rPT0KJKc/aeh0Is2Ecan7EaBO0Z
YtHVFwuFE1A/FHePU5FHRQofTSg5/JGwPG/w5SSmgjzwMjYFnO9ZgYzfl2p1AK9S
VYWDoAeJhSUp9kjYs5sfKJ5oG3iEZ09jGlV1Rr+q39tZf6vCMonL92D9g/brn2WY
UR/e5YJfFcIcL+OeiuvNT3beGt2oalK0iaVUz6k34q36Y9ooFsBqzrosrreeaIgD
47IhZePtcuVoo/FxBV+akTnTGJEaAzDewO4GjWzT381C/syxAMxfCxyxacilwmA6
IYO6P+5B1VJmhSaKFjTenyuBjEKDd9SMhAnf8AI3ZKPMdmoA5cPIlD/Vz4F15QVo
`protect END_PROTECTED
