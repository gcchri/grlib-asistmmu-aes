`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1f4c4mJjIutymyTkw5KOk0yHH3jSRnv3Wt1tQsFXf1deyTKg5LumV4bl+ZWsGiAw
hoT10PMxlGyqiF2ucmVSDN/XEezKMY+dbJpWFPNZj/c5WQcQCloDYv1e6515uQkC
rAdRl/mnFR4sDNEm0yMHlVUQjjRzcrY702eEEH+lldOiDrGOXIHH4KveYVRCIKro
XMIbCMpXzdM2IpCwt0VW0Iu4XWcOR6iCGNBNIDMGtCbd42kU3m2BdRcdK5Ci5SRq
x+d4MRSZcCrlOyiabWXlhw==
`protect END_PROTECTED
