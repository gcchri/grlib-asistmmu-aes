`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/bRoYWUp789FWQ/G3nO92mLhn5kuNzkIR+y5CVmDurXK8Q42rsD9YZBE0cK+QHF
QhJJzC3kgJPN5IfIZ317c7wJCGsEJtHipboQJBdLCAWN6lECTkEOaPV0jS1zZDPP
mUTdayBWl8ecgFs3ynQguR+J1sAATkVh+HLNt1bj5rQsO7LvwU2m6bPKbE+1kqct
7oQUo3ARdfPf2XTvTpbTMns5A5uFt6z8zhj0T7xZ2ZMffSEbyXOekvKpbNqeCa/7
sN0yw2AAAaiVEFHgHX0WGmtpEWENZ9c/xhVK+nBReAAf0IXleoy4S/xbdNX3r6lD
5cDjxtAQTphopwDNXRMnHt7hRZk+IZo551LXgstjyswdVVdcx3vHPLR5ip7sEId/
`protect END_PROTECTED
