`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6mtj6vCx8/N/asXwyCPfM8VaI+K6heYPbWyEZJVf6mH79bhHPK+/DIsEiM2ZiEBd
a/fVG6EPl8CdE5wNzX53XwPgbPy+xJkbnoDzgQQd49mW9/Uwcr3KXfCgFM2AKiXr
/TElV+6XqK0J9hwZWvlOZLsbZVnIURhH8R8mdFPyyw3Ml74UgFmeyK7Il8s9TOJR
FXO2kAJ/RzkefSQd/+nWT9I3QOsTQYfhqymSK2JExPRff4gUi9Hme2ZlUu8vCvmW
MIskDekQsYZlpDZf1bRaxKZzdnInh9VErbqpLBDTQHYu0d+daDxJBtRp9Z3b/WDh
KPrLROfniJrkJ8GtsDla4/7ztL19h1BaZDg+XMwamM4h+ClReBiRxjmgdRw5sMF/
aB/7E5gIIKUTp3sw1/rZDICiv3EIlHnNSSNUvdJMPqw=
`protect END_PROTECTED
