`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KDSoQSrFVSs6PztsA8zzWsGTIf1ExvMrp2S/4zrkXdYXgWxyQLP5muz/tKvGcDEk
C2KNYYTjxyRaE+C759XGVnsCXFUdfn2wZw9AEzMeAFDWP/SXEL0tVOLQqVxSopGZ
24F/7MEGB34lmVw5TBWgfNDFtn13OfJk3S8W8VfG+Z+z5TcdHUQIgWc5qMb+u4m9
ojU24ywxXQ9meI8ZjHA1teNt1SnsYEfMmcBadM6PjEFdnLkz6fFvcIBWoQIa6rTh
RlyeiDSsKsbG6XfNEWlJgNO4PL72H8COKbXHzu6y5ceSURdHF+sy8zoZemm5Kr97
sW0xbOsF9n3SvDlSPPdiuovhQR3XCqwl8aWWRMuLZbQ/HwuEvbBLLrAiyldRUt0u
cKALkwSaBo9I0EPi/1wz0bkHFzUyEjEi24NaPSE1g7Q5oUjW3S/k8yJusaeTBuQP
yYVC7EuJRPO2XnJSkZbd8pHxWioJuse4LzAIeVU95FXmqC3+QIX4WaW2xX+PoJS8
lwjjYwjlUR/uJcMEe5Cy8ICjeSOKj5Deg98xrDgJIK0xxyLoe4sCFXM8GTjLgL8d
lTqyEbaYLVuKFJvHwqfFPGnaPWE/vbgbenlE8WApyfL7X/bvtToePKwv7+67t9Gl
4x6gZJ3l4l2ED0td0i5UlbvYDx1T6hDL+AukYIxogPyR1MVKJ/Z4JBGaNxdd2DC7
63OC/NOInN2Y6BL3VUaVxODCF5oXBcb8eeOvPedxgHamjDVU31zRPoikZwE+twjD
9JBlpbfHQKFgZ1m5Aa5NZmgziLobS+lDmQ3dHmd7N0dLEKsZj3SyJ4j4RM6vaamM
e80vvFuGLHC00P5+m+Kas8YWcPSzMz7g2Nl5A7iLzALDEPOBiudxS7JzNAPiLIYB
eJfIYjydQc6L2z2gsn2Uk03QRoRK8NBJjfFeuteyTbCEIv1TobJWXKuFiuD3GJRS
fjhhpfNX92oEBhSRhDj8+xoc/7SOgpBAJ6PPoWfV7Fj45iJYd7In5EEM0Ze8RKVJ
JU/jO7QUZFMe77Ves1vjpaGrg5LEP+CBLwxCeLXTCBcstaPiIo7bjXGZZTLVfZhw
dt1LgYuZlAuDBvqVWqsluUGOf2eOSShIuj1nThQMbUcmIDvqIrIHpqIAIhABBMbI
LqNnJ72fUj7kQcmjRoi5IZjj3VRu25a+F6//XR9E9zy55/7WP2oe/Af3F3nq+kAV
zlahH7HW1BIdhLhdgg2u6y1daV0Vf1EHDKaVLxCoPC1QhB/2cRgMh0zTpJ8z/5PJ
tW+X6vO49qTeTEYd6ck46MdUDR1dmJbnZw7OvxoyaVzqXCB3t9YH9x034BSvLdBJ
MbV9db34OsBPSbe4KFEHwEQjvfU6hEjxCPbmq8T80/nVKB8hdxf7+9CgikCuHU+z
KcRqi/PJhMj4K2MQVXtFCiXFunUw+hSS5/vgnFYirZqGKoXJ0ixGwR4Ele/52lI9
P5wuJ29OkOoxCecBXIfaxa3puPEa38W0isOreMwB/5uh+UwNalDkqFgzXfIHvBLK
ZrbUE67JmbRoxdYm5xmoffI3/uK1RDD9Zb+ALKXzQ9/7r9+heaPG8VJu5Y5GHbP5
9/NED7OOs4WBpPNCwQuQTbVjfF8WuSQxNoU5LMmjh86d5e3F5YQVbw0gRl76FuVl
JWEobjsQi851o9rGFYMlg6UPo4Mjg0tO1uuFurwypEKqvtY8IaLf46LrfTAeg3Cu
PKm6tuZRzQUo3CK0UzlqeIXdvzcw52PuAS5EfwdkK60VXDgZl1PP0LiDD8bwD65V
zdlmxo/4kOQa4UP33tRjduB9uq+bl/Uz11V3aw5wTPYSMYvsJpQ/Bw230piI2NIT
PxO48iXWpDpThoXvy2AqEGeNMo0uHxBgB+mlZsyO4skAqcP3Euwf6sG6CKo6q6ty
yY1/tkLj3ClufeU1vkjcj498i9X0GApxoX5QscihPnQj+PEXw188OyHWLEsEcAk5
Bk3Gz3xMN9/0FlIYyzqtX0Jb4Z3kyKZtCzNcVNtSoD5kgGcsSiZoYcZ0Ew9H8XWX
mdBa8Z2iVk+gAr77OhFM+phMqxqzjdseFhi4fVSe4r6v2aN6oh6ofVIx9B8146rZ
M4sGlCF33wqm4JkRCGWUJXpMPCMGPrv7bHn9UiCGVenB5r40lW/GxDEfLZX96jZP
L9oRfCMJfm4DikfLw0+pAvuZ4ougGSsz0YDS1WdXqPaS3Q4wMwXN6EkZZZR2Q2Pj
DDxCsLJuYExSK1EmYk6UkV+HqssF1YkWl1+QRsoZll4sWbxe4YdaQLAKI18YbDyd
Z5Z9A/kWp0XRVIp8eKy0CRqMwAF0yYFhpfFPdQ19W128rSZqCA00uXNFwUwilGw+
VEx7NjJOEsge6xoEzDWD1H//17Wn1juRdIi2cKkvy2F4KLUcNMjXIuBnkU8aZ3ef
vOe4yIzTa+jSKKMw6xMqNMfbbEneq96c9ezd3RL9XJ+YKfBdY8FUa8dlA1VFQr8A
CbUC0iQC5Fqec4mnyn4jr2Qw+2CKifgQhVCkUICKANEnoTl18bdNgCvlNlI3TJTS
vUi41dxaCGIDFx95UIFr8S99WBmJYdfdqnUu1ZykW4WlMk9NM5Ol6TbYDcqF79vH
YAPYihj4iUJs/ejjEpNJTOo1KScDoizn107gtel7OypVUM6nX6az0MV3BXgZajG2
kc8UlcpA1tvz/LtGce9B6IwCIeNVihV447jRCjIGpjdAvCj42lM9+MUQRjzjQtIw
mPa1mbVyCtRSPoYtuyxNp10OMloyMTl2tDTmkUkoxgb85QFrZ8adYDr8n+J15qVX
vPpCoe9G0eGgCus+iiVWkRqvGu1btgPfj9g7+PyLjcqEh14Rqk6MpVR9J3hXk8K8
iLDMNdCnNBlrVi4+24M9Z+bGd7DcB53O9EvZGcMe54unX/ZM2uonoe9Wkkp4RQwf
4kDMZ+mHlaUB8uoEvm6MuEOSUlOJj7sl5oOiNIrlZ0mPJX3MYI+e/jjDtr3SU7Ao
8WpF5JrRx31ncloA7GiQqpUdmRrpGVVsmy3XOoJ2csdf+aymATopbIoCVgj1k6Wp
NuwfAnhVE8m92FChtSr10h++jkQur7go1Yh38+isV/9SL6EB/g/mwIElFRL0R1YB
qEpCdchVq37NWRyjr0CPi+WSdjqMMfmrerdH97pgWuEw3OgVKLc5DJHwNMFj+P2Q
XZLzqOkjiabzEUpA2YiGjh5pgNdNSXpLnGQs1Xejt5/Xd9n8ETH7i0kNOuPAyriF
BTUc/tDeQz9TrHE7lDJ7ILDr4m91e0nmx1jp+QG4Hhnzf5ZbKs9gUBcVxwxNmtm0
zcjdR2gjv+KBus4+UznMj9TBqHBpByJURbHlbk3Q1iJMm3tLisZEfV/3nszmd/wd
XM5GzzmypOcoy2oKeyomNALF1XEfjxdyo7K1EM/U1X888iveQ1+b4REKSodBAIHZ
efec/9pOvJkR+aD6Wtul7YXq90b/SB7Qz9bFPwYjT6DYzA5nOe6Q+0hFtTOu3acq
dvPG88C9wobTD2HZaVS8T1xi78JAQPOnbtV612KGe5RLnuBBtw0CR/tyHaTtu/LF
cnLIiD7hgQYz/Zptghs394Z/iDXLl+kBJy7bCAepaiP+TMu/KvSRnvg3ZfHvo3mN
LACs6aJGP5bzC0j0/Hws5QUP+i9FlgWFVNCWTN5DFP7aOV9NvbzaF1DjewIYrWYY
C/dQvsBukMCtVLC4hl6DFp+yDyRLjYrYmj698a7C5B1MATQzfC3sUWT7LBU6pEuM
nf9lwGe2kSaXyKCtmjx9ktMaPGPL50A6Fm3ZjFnA3mLG9HGzS9+Glky2wd2y/MgC
dfrt1XQTeoH8b3lcGVCpBJJTS2eA9kUH6yvwK9hvDWSKcFi4inogvVUDaviTANN6
sEBnjxZdG+fkklMAZkO6g9DVqpnOTMfw1NcXcyR+P+XR1ZazwZ503Vq5ZUUI95Xw
JJt2mpH3yT/uXFSq9PGbMPAsDqrV948/RAjloUbpx7goJ4Z642J3xtat17pHbe0e
AOcqHzVHRcBczeF1ORhsM8PrkcwFZ0Uo2JiX62f6J1BAIfmLN7GgMk0ajhIZPtM3
A+7mtvfne+qmGlJoqirBy6dkDtMyQ6SSAyU9jgE3q7GQvYJE6GfJVvmG0SmLmjK6
fdcRq+CDc2nQXxH5q1y27n/5GB7GgrkBluNY8T3jAwTXgHaUXtyPOlcgCJGYbzoe
SJX8ixgRY0mJokt1NV5olGT8p8t8ioV6+CnGYUqlVzKzB/D87zVs4TmpgK3JKWnD
ohvKLBQ0lgn87NzUmKYaiL3JHaGDJVKeA55BIkiNz2T47OxS+t/nVcb9iQawVuXz
e8FZCTlew4Tg0rxw83Vs8z0wMDkgPKWRSy/RrVV6nDSgv8eJaphw367YqH9gmT9g
59CE2PwehgJ7zT77aYiLSKq9+2Y9jNl8vO48egnGlPungT/ABRN3WExTVqZR5ETy
bwSg1t7RvKexawNy3JkOTjOK0BK8suYd6Dpfvf5HtQL77wbp+BR10lWLUWSC3jeD
gus4iKVEXZogNHykNKdtm2GDhJY1vGE8/NEYDH9R0mXMDQbp6cKUeGPr1LMx8TNI
C/1WL4RkyJMslcfBzdsISBrrBtio46FIbboqkXaGVBspJg+F9gX9sYsLpn7BEnuu
J3m1say6tTJS4lOMiWiKgJRLmysnE+sxaVEMgJ8RfWnqytTdlgvtY8RIFej9FRjN
CaPHsuFe7pa1EIdaGIdJRo/xXZQAZt+8ghod8fjBop2MPnxW5PSlPrWPMBUUCjG3
Kjax8MhExXrm29eDabTRPeUCuqZHqf7AbMk5vbu0M0Qz4jVECoNQirOfDyY4AwpV
q6cDkmTRFfU0GRMWolqzK6JyD3pE3VSXrIY/j3Bza6CZQTH9Adw6pu9qMoT0AmwJ
DpToMbUEPxmTivKPDWRcDDKo8bK6p2k9w7RQjy14TmTB0Tiztqaxs/F/IrdHPD8i
DujkjwiSVOxudNpecdS5LZ9/eG359Qmi/kkOgL4fc9H9zbzFTsqvBBYrb6okGmLz
BK91qBHPgaZmL+dENtwIDhMNL6LN3lKzFkUIi5GNdliu8cnPg9yXLdpzRUOMf0ww
vP/a7TwFuqWNPfTlaXAFo2hbh/NA9o2foicVMrTZf1491jbA26jShQ9JRyJpa5c3
BuNVW4mRRre9erOVtoRgKzauGzSyB3KWBahjoAd8CfQHZf/iHdnBjNWUt7N4mlp2
Rn6ZhCmmWHgSideBzcduISOD7SGY77u1ec1984kR4CqEKc7C/wbvDPgeUe0yDCOh
/Weg5acTC7uiXr6y4qbevWjALC/R3/+pHjwFztNeMHKttzYOOBkAzJnYi8lTv5Vp
sUs42Zle9VBELppB0zY4b/R8SNM5NdRzWp/EZp8CQ9LWVfd9JHQb2ybgEknncp+n
umdvzJOVQaXM4Ge+p5WBRGV8d90EIjQ1vSZzYvRRRug9QmCs88h/1wFdZ88Z466c
7S+vRspSPkRBqAF8/q0xU2Qp0aFhKpvV9WZickfLusPJiYa3yYinoVC6ob18NhHt
Z5wnbRO881ge1lUclyNMKcloUaVcklGrgcibshl4loUZiQDwdbC2QZs8U2fxR/0M
IoFH4QsSKguu7kP0XVMAzb0+8n3YA9LF4nstZiTnwnMEL4aIfoWVaGv5epYyky4j
zqHHUJuW7uM+PEfrcwry0Rc8f1+wFewifWnaOWCAsUOII5bmDxNFSawp9o+VVR30
SBWFApI2A2QVM7JYHJLKjorBnr2jC4kvJjqvprSJohAcGJkfBzDWoS+pfqioDVli
V4va2leouEyO1g/RhdYcSl05mOHggRaxORJFRluxx9OZ7u9a3frfZQPelhNlix2S
+f2SE2pWPG57LoWaQdfp68L/GGZpfzffSHOhhPlqmr6a49UCOPB/AkcM6f1exGtH
U1116g0nqw3+WUHFGJMWeWIa3y4TNVhXSj4DdmS/eyB3cX5JOdRoBB+9sBO/8zXE
WqFHrHLWOOIJsExpw5aVmwfnE9Mz5Cmoh+kI15QvM9drK2rkur+9YV+1c/amaWQu
CyYiXeScXh2nhhQbwszDPczpKtoxBKAbe9f5HVN+755iRQFh+XykXsm3k7DI+Mag
+tquTUbYVuuGvU3RxX+BVXfsBDl3B/8iFFt3MQeM5GOyQiyhTQ0cLnU0qW7ctWuM
O5C1aGzD0dVZVYYeR7kV22IvGWxGfGrfNV2paZafUQym+8YyhKwe5R5gBOSoaG09
7/2eUvjnzoIJUEFZO1s+8h3FDxB4PUKsqo4bg+PtuDxYIEZ1eqvTugtFfF1AWLdt
GOPHyydu1IlLX3t333wWbtPBpf2j8wwwj3abxLxvz+qIcc4qIFcnDuHVjADAzKSP
nuatyeGEP8zSDWXUjOVvsnbnwUfEKMYrJ5Q8pXKF/8XePNanFHetPKVyV0biAs/e
4ysD71pXxjTvFcq549iTrbVaAbHpqi9Q5c2CQS+GwWGtcp+KUPCPQerAobzOEHtT
rW3N7d9Yad28iAZ7XlaCovbH36k2OKxwRy6RH0im29FD+oOpqEQz/zxBTl8NjHUt
YTD7SFk1rO68iwzYRAJUmqj+jS+YpYnRm3Bqr7qM6tR4RWoD5+GUiDnA7BTZ6kyg
RAmNA5o/EI6SWrv7rfI2THzc5ln4BdculQb1oWlLgMZUL9MOJYR66yL/Ja2+G09Y
z8Yj22VQXTmLKVJDcqMMUsT4//W6SHnM5wXmptcj77JV4iJoUav42lHAwxHuWGDx
b6nLvYrkimXO+aZbQiCYFvwNLgMPL6TMjDnGPYVY57KAnFokqgQuBlXF3gsWMzxc
9CDEz6/XdoivuJBAM3vVYadcf8utQUKuusLjFyRXzARwkB3UtwyK6ieWkH/AMNBe
j+QFkISqIG80CjUZa+QexK99XTFxd1DMl2KxV26YwC9ahtIEwV0vwkHhy4uh6mZ6
TERI5RVk7YNKqlHo5J04Z3jCOYSQ5VA5rY3krBDDShu4ZBshITnm/zigQEn23FUf
rkuNjejlVtEjJTVuBdiUzjolYl+xO8/lm5W0Jk65gee5Gw/KNRbdt1OqZBtDuShu
ujfEG4rVKCPRjJnwDfRVfBqNPufifA1F1snjBc1xhiFeFyFJvgK+LNr8sL01VLe4
DBqXbIjkIeBpuDVWqEJsFjacWV4oNHABz9t3KvTQ0HHQQGGBbJveDvRxRDRD0Yhw
6zwdsQ8ooa/zYMh7ExbM0vTqwqgUwtmSEohJI7EeJyC1+jFQ4NjC3SKEg00lRCCi
KQJxBlt6WWOMAgBp/MLsVBJ8QRJhkdgBGav1J0WhAAFBIbzYortufk/zBseRKlIb
o+AIqZyCYGU9vDMPEoyizzNAMw6+cA3UahYIqYSVcAdG3USpG3Z8C+0Dy+U36vaT
FhbN84RyZGkfly7ATIzxsmh1KIb9cEpvsdFETnPnr1ToIdfGg0MdXjrtQTO/j2yQ
rngRKDl15xF/fUwxaPyUL5wsq9X2WmUtreN0nuC3YPzNL41B0ciQqNQJpxbSwROm
HKUJ75fAVs+F3+EW4iFdz7vg4k0OxI503voFG/Tvx2v5OkTBAKK1k40GJftIry9w
rBRxZen1ahisa4sqVH7UW3VYzA/Sz8XC7XQ23TYhNTmJQaz3euMnrmBfYbYX6ZQo
2+NwOZM7d0DYse0t5ZfUTmbCq6e5hiaHi0R9fUsSEJXiAwQzTcCBQy+0y1r1jDiV
1XazOedljflm+ygROG4mJgJYUbFgFwsVX2Q5yW8vL0pp0+XWCrSBLAbzNXS70LDO
sdB8r5h9GC7UXWj/eEUIgyr00NvIeetLr/NfXhHlpm+cokuOAwQOoU6HnDvKrDv/
KoOqKrd+Af4f7JcTzEjyMxz9mPiaJ+1FU8F3fSViP0jg4OnOMWTD/+YOs/IeDLJO
TYKla1K4UMdvqChM73FQdTZlsVLQS1tR34V4pEZo/SfSnyiVlzyEeWeyiBzW8lmB
ZlMItTYA6ND4qj9jMQfG3DxsAXecoKw3qEZUfyxCRSABVKtDfjtK8EIXVCDp74tX
k4SZbVyDvW0wqDbQvHcYt8c36Q85N+cmuuWRa+dPZkWBTVHIFY3aJ8z0CwSqkwvy
ZXc3lU/594dVr6987YL3uE0FDFeOgvO55pXQdq3k+rPl+2d2Azmru9R3XCH/okwt
mXD5E3k/T/he4ett+wRpi7jNqnAlpLejEczd80H5V7QR/yhj5tvqtVLsFM/aPC4O
V2LSmfN+CJxUhhT/wobNeidomPesMBoOejRt1/pGoPZsY6KF04VRjy8LAlSPuXMm
I+sFOAfNsG0wnw1shco/mFUJ2AU2xGIg73F4q5fGEcFWzMIuhjxhacaQsPBVl7L7
JnRRkRdLTw+S4EeRWaxsG7pnCwVdziIQqUmXDkwA+EU9a9qQ85F7P0kpviBgSbzb
cAO40LrM7d+SSOfwh47DWZ7IXacdmjuwr/4jonk6fLP0qM6Z/bh02Hm7f0PzAiHJ
SA9IFcBnjVPZVmkOhUQEGF833UlOFiTuakfc1AQaTqNGDELlRY8Xbk3OWZnqNL7V
9nq2bopqpIPlkM9JYF/TZaQgqpUtn32DUit3cqTt5aGflasdNWBMRmaQ15+G1AzW
ZG44AeTz8XV7yI4kSkEOkRrsd4yIzNHfJbSPJI7DjrBVFwl1/DuTz1bB7BtKUuZL
cMsPmcU2z6eaAT7+H7zyZRJf+3RanhXrAvteF9yVK34y/WwNvt/4JOL8JlPSCMu8
Xn9Bl8vs1USiXX94bomVDCKHVz+bNPp7VSKWxahBsRQpspm2tpKTINFi6hPtid+8
VmpzfshfuykhpzJeIP1wyvdqdCxbNh9CPdt5fv0Ma30JCSSWVgowq6d8iOR6Wwfg
KUWiYiovb534AU7tmxj3wz3J0vkiA5QGySVsbgV7/12pq79r3z1lMgQ9Q1PUh6Ai
v6VS5CV44J7Koknq6XEENuMcjSTdiH5qxC+dhfel9OgsNPIVm73mLAktAl0DA2kl
MelNlIj6dSxUu568gAOzVfCRZgImoBENHXzcDItmNfjBbngoH+4hDO+og+wKJjh7
kmS+GAoe7gHZHq6N94s6nMj8x08Ryvfud1os4bgaxtqAyujJVoCon+mrzn1WPA0a
NjoCIIyH5HJh+DeZvMW6V66WDV5lVAaxGKJ3LjcfDGzvZsjjQWTQNPApGebmS+0B
dS5ju4U+59ZufqnZ45LQ6pJxUrbuq/AindYOUgAaHRRbr+MDNvxpVO5Evd7SkOMj
akZVfpgiSg2Ii5FXcupqp2RpZjwIYCuJGLw92Gj9uEMdhMLpALa7us1dFMlsBJKm
bhE455ThcUsqv09ZOE65B5Q/bzzG1XOrm2BRcDnzM6ZIq7B77iUGGb4ZVxQKexRl
C662wxLKYUXXb1hHFC/aSGYH6ghDfDTTnXCAv7T8PtvBP14MNsE4w9zcBvysJBcs
1X9VIJWxqxozAsPN/dUBx1jgy/1JwGygYfVAfePRP5nQPjMVge8ltIGncEn3E6rl
tHrTOiL/D8vAOYU0zyXHxkY+X/sd5NWe6HHmGsAGhlo8TWMCMS36J/CN4o30Jzbs
GEo0kfXb+vLSJ92ARItYhqR3h0nyPXkkFMfQdlP/NEDJ6p3V5tZxXXktAnnX/G2l
4A5cO874wsPhgo9Z8vgEjdbVQaNhWFh7XfGMzRoxCl+0+QKrzxUcyjBkXmAwD7xi
ykvQibg05qAp0sp5NoUAzvdOMydnbrZghg1oL/Ms4FZVILZO2MVVq92VKyvwzyZ7
/+q7dEtw1pbrgdjcgoiBX76Y7g0IDXEnmbwtUX6WLhiLg/3rY6g/n2TR1bMnY+v7
ukoXLQu9ywI8cE2eNQSmgVfMFFKoeNPKypth7gep+Io9sDY4L9YUowdF/K0Acwva
I5PXNxFzm0jPPQdaOIaAGBgzy152ZlJeUIeY9cHrHYXv/zbCkubzQXeQD/KUhf/T
BWYhx2Mf3Z3xjFlK4uUQkOGnfyrSzGT4gKcyPM1gXWmQKtZZCcula6spslwv6Wbv
j1wgMDy7uhm1jCjdzMvgqlq62JIaXX5daTeUqFnZnENAsDzRiEd2mO9g+5oarWEY
Z94mRWB+tLl2Dn2K8q2Qmtfcwede2bMtNk8JIjidI6Wx5xCEi+hOc/RPQil0gzlV
KC94ViH0yuiEYLxTHeBkeJr59Qhzoy620JDe+GMRUZ+93ZU/oujAgBbCToUPpkgB
+M+bx8lNIR/DqRlHVDM/wzqrFTyUqIQHouOnxaDiwlH4lUQYipY3AACHWPpPIGDq
f2DfzwI1qHmgt+59yIg20p7gldY7VIXXa0tnd4pa5MgMH2WZA+7biNeKAQ4HuG6y
yK4x2H2MqxaG86E1DyFC6/ha+4cqtBqmfNp9c7Z0ynPY/FHDNXx3DT2hRp4pFpyr
puzRZm/vNzPiAAuU40/g+jqtWJhIocxud39qOowu6p4RgKdX/08qosNSE+lUeuu8
6qt3J8oPIDJygrH9Fx/r/6TJll7YkYeJ1fsgq4asCZyFbY147gF1kl+bg6LjcHdR
szt0wJXwxdscYW9Ux9WhYT6ZfzyztgRWPqFfI9X3p6MEXt/YfzrVwXT9WkBmGzqv
SD+/ksP947nJW6ZRtNBZWBVAdn6FP/aSq/2ElfQQKZhmD/ibcLr1QmAuL0bgkZS7
oxxSEJoHbyBOnjUJfQXLtZsF6Wh5tN7lf1x7C/z/TKiLGeaGwS/iCanFbkbNCuTA
ROoHTS375HjCQPV1+X/WMoCWND7twZiRgc44d0NlGxWuMIPjg8eRImIKMETeGcH0
/tMdIh0dSKSxaJ4vg3veHpjqPWf/XEZA0SDqty8+9+z4LeatMXmOk6iKsvjUz0Wf
2wN3NZD1DdouJuJtVpZ104RHXDhnEv8BpIL2K2q+768CAS5dOokQvnuY+oBdfKUf
lQwYoFNlDSd3OlJon+xycu2+E0gAsvaxOVWwdYM1s8IAcHM2oB8efMKXa8OBxIlk
bUz03/dEoMbcU6SiACUS8iWVyPB5NDLaRfmBHYV5fd19qOtsJBvZ907gyd/x+CC4
QLvhPRMuh10GHLKdqNm4xxEarxtKij56xTzQekA2is9Ng+9/pgfhYLqk4yB+yiib
IuNivPfK+fuKEacINoP5UzFN6WPICS3+9kYwxBa47H44aH+7/NBmdXz9J8YXB/Ho
Da1R/8oajxRVCcBDfDtbi6p8VCZjEucrU7MlhxFv3WS8B18cI2NAufWW6LylYAQ9
sYiE/YVNPQvM6cMrflnkrdZLPc9TRNacnfw4Mm9WZJwiF/L3w6/ZoHzHffG8QFdx
/IrtzI60l183BKYGBbKasi+HJ94ZGZrJBqAuBxNU6WZTlQ1gOAa8y4aeGF/feHW+
dgvKZCv/Y7v9TVQC8lHwBkIGqyeRn8I6IkxBwe+zghFzqF046fJomQuNx2oS1YM0
J6pe+LIp0H09JxDtFjDrShv9EsO8HfBU1VKTgHgZD9RaPT5mRN1YSNncB9P5gHE6
cec9CFVz2QAHcDQ93A9EgZroTnEbUtz5SLjBHbK+gTCEbm4ztnOGmUD5QmA+FVab
RpONe7UV1T4EUBmcQ4wZTkPVJ87deHb8fsOkbqTM9WHFW43OzXgaEbpluitmQq4c
YsTIpK/ZB8wlxp5JoWiJ2aa7/OuD3V3bJOnXbVQHcHYTmNbaMfepkZ6gE46U2JN5
FulQ639PfJiPHJ4BD7pvgeY5BF42BPT8MPBlBDUGxoxG4nOaU6GPak7kf+UMrIto
MK03CXznxqK8GkGLBx6iSEGWEhCwSjEvzkHnXkXii7EsJ+x5LI4q6QOYk0pEYD6N
o8Bkxmrkdu9qKbsRGuOnNVlmPnwYy3WGTweYREv9qzFk0cLqaqxX+iLTEjWkAoaQ
apC4gZjE/G48n1T2L3Oca7tiWDpWr9rsBuE4QvSTCXLXbtQ+3SKEq1bZ9TxrlTB8
zFHPvfL+2o3ajSHB7TCTAyQ3PHrhzumr+szK4ub+xhW8ipUyO7gxLX5ht3HUHqiD
Dmg/w6rtN1ZIStX6uzvu/qe9DVKXxhkzGBo2e4E5Lco2uBoA3Fm43M+G2tYlJODj
Bi60xqz0CNEKI0lMob6xufJNhN99XRObKNJWyoJpIz7pVCWG8mGmiSgArrJgJCUU
/H+MMqtK4jcB1vsLnv7F4tY6XpAX8UTJXBcuscW2HbY8ixREIcnOYGK826a9JSAu
Hs4uPyXUEB15R/ELyqDUY4QyUgueCqkfboeSv3kWTAVNaUSpOTCU4l5fL59C8NV7
PYfWZu4S8a2bLZ300cjyUFCBl40qpdBqFb9X4MqXsHWHvwmRR8YRvFvG1Pwn1Xh0
ss2+fZwNz6SsS2Hvyj6IZHjTJdVs7SMsL41JrOArXMioncx2MO94jb/8yCnEtI5K
za98ZW4MGe64Y9IAuX0xO9cA0O5hE9xSzW2+muvyyh7YGhDvsbBYrww9s4RYXI9U
xz7hvkST70e0YUna+Pxe3fydUoa3cKUEtWFhHnOcDyGSDtTG/jFq8DMbn/k9Rpvu
V0zJAlcC/xFcs5CbBbweSj4wlJW8+VF6el8w8OXxL/TkIofNpSz4Og+xpKpd5y2D
B2uFgj//dIWhQuxHCK3f0Vqf2P+cI4ECN1L/dHypsx5yJxm1v66Pa230NjW6bPYc
xdzKrJuBls2zbcdX4lCjHH0pGA3W5HjXerJiFW5Q9f2G1j01EvqTRQuXyzAedhYX
lEExO2OiI1cyWTimb8MPsUTzSM7J2kiaftmboSA2wbbmvUjI5h3UPY4iKTT5B4Cp
ErCyNFvPbf/LobiwZpOAHmiXEHp522tZxzD8gmB1wS3M4rBm7Jg336Hm+sKlE4Wx
MLHjwMFaVTovi7AtCEuHZ3u2ihZd1mjo3STV9/vj+61xk1FdgEah3NCjt5VtGBt1
oigTdC54XRS2OVraYqlNK8TXtepciVVpnEW9LlJfrxzUZm6t0jwdlhMyzAqvEW0N
tnbIyhWz4cPqTkzeOEoMBLFOagtWBXIlmabOINwm/+1ImQ7Ihm5mvN3GM/ZOQ0is
KpkoqcJzLM+9+Rzmr7GMamSdDpa1tS/YDb2bgJJY9qrio4VYqgzaF6Gy9wnSqO9r
ffSc1lxSWJFvnxeLp0maGTJA4c221UJdg3pdnuCHYH9s+5GIW3wm3zdALQRdxTT3
Cbo9YLEiBc8lYWZiDLZkqRyWe3u2/dFOYYNf7DdwlGe2C68Q8YpWl32h2eq1XZb4
t7gjEut4ugPMbpfvFo3Lm/n+jAOIuaD2CKZorAz7cJcKAI7EKAhjwM2kqzO5EW85
Wxhy9jcuNBgxnYTSV12owAoXsscWF7zpUA1zR3UbfBCBwr6oNh6FzQngjuuUTblp
cv+4aOwtRjRZjKrzfO4Ltkslpa4k5XlJcBOlrB3Z5qQikggBpE6rABRMNdhdsCTf
XzJkUaNNB2mCK1sqNeIfvNUv2dn6fa1AESvIXmTys0KU7jjxUH1qp1+b0a4CMvPY
VwWquhmHyYGNz6qEQTSZfOrF9jpSiQF0dtqRfD7pfQaeVbfR1tMGEgPUlcvDb8wn
++/ZihfikaeWxFrwKVleBQCx3J55c/AzpoDC5YbsmPdrp0nTqaQMCi4TVavs6c8o
4GM6Er5aDxtL9ebf7DuAEKBj53C89vpWd6AYXnrVb9PMau4FTIxfrZ0cGNC1DnJE
914wKCJR4lpsc6zEOGfQLqeGRpOsapRmXio0BlkziRErgTIY9LW6Mz/vhigDiI0a
bakMIg+WbaoY50oR5nhElRcaRzulqbFGmnJ/Wm0pGbKkHoENSjgCi3fLPfQaffKU
qrvh5HKLDtAjm8LFeJ9O1cST3JeAqq3scd0wbbg3ry8t1/fp5idseNo1ll6JDapi
NE14dzyIj+tPaO9+F1CEbvP/GEbfyhnzTNmDbZPNiUBZtQBLSQHDN8P2mgZso3WQ
/BNRy/dvR0kwstfNFBEj+HAda4WGsrOrJySjob/AAFq2QhOjDhaz2mcdInOMT057
pQZiLBhxGSAcPDSByulpvTw/+ySWJVbqUglSqiIMrT8iQshjsiKPZ51Og+HTPGEp
qxqtGwiSnBcRomSnFdcfcTtbc9XMDt1dl8Gbqa+ZxjWe/acj9kAOXXcgvWc9sHsy
SBtHREHDRAcKGYD1X+c5MDZeFU1wiubOF65BAayDoIyHe5l4RD0I6bnioSH8Uk8W
i/HmYu3xvzi8IShU2kBKeFKRTtOVABI3bZNR/MxNMhkIhEdTaZbuX+MAueGziSPX
RyIdqQhQ7WZjmbDbBGsObUNvR2SCyapoahhidsAMvNIZ80Z7sekm6NCwlh99bHMi
wruJGtoHAQDHOaMcI6rZc9gQsdxRnTHFaP6k4bLzVKkSvoHvYnCdRu/NcDQ2sAMh
MyeFbMIeQe2EChvav4FPu/maUKxzwhZ/F5VGYUpKrTBLE5r5Kar0bkyOhHwL8HRa
KV/PVhhgQ9PYtXc0xIt3ggwbn0KBtTJlr/K3Zqt8hefPXM1YWy+NW/Q+m41s657B
yX8WxMdUZLCdYmtTtCJLqtUlGXcoK6EJ+fRYoblOMr5vFczGtELHmX5QxINi2jEL
AY1O/lhClkBZlWp/gCJQySpBQk7NuNSuG7EGnahN0uHqx9SQkHTrYtEu1Ajrdxg8
BpqNsu9TY6Ez16yE0YcT2C2S+Z/dtriP7Ej1WRNLHlkua0JGQP5sGFD9cYItnZE8
7peHByzxNOltkM17xf+0vfE1gdzomTaLlysE5pCgYFuGAEhN7Y4yKeJRQNUSIHBD
gAwBlGQXu0x1Imnb2UDktx4AoTQgiDenLbRHUaVy13RAMHrC8WhQml126bpzR7lT
HuzE3UmeQtSiZLHiChqjfAvaBAbM7LI0EzdxWmmdIsLj8Uiv4NbpaezBaqHREOU7
FgkxkT9eZuuIFYT+Ekfa6C2y2+YuwfV1t4sRUXfJbswwPbsI02boc0iy5rXDDxlg
mutzXuQoeN8PLIYBjVZXBpKSVW0sHOJzemeknrvVUeFmQQj0DIn+G20qdCvagHGP
zxCgVNwRs5tF5RTJ4IN4sVndwgz1Dk2bFWetCHa+1mzmB/rQoL5NwJC6hBTrjl8H
B74KwTeVTCOlEXxplgrN2yVkL6oquiYY21I4BMgZF6pA+yo1yeV5qmAsCjM0fggg
eGHeVlsIqvR2BqUr5faOdm8BAa9f0jhJ6YAGa1jDmIgPRyQ5vjCRvHtyma9fa3ZW
66H1YQCIhoiVtA1bMkMGP2x3lzMmHOLKgJPHpb/ALG7qIj4EXiHhYTtx+2IclSp6
n/yln9DC8lTFVX04zkhH92aMXkODrTjyM7eKsDd9EmSLSL0LDuyiLDH8f2I/eXQt
kZpThT1RE4/jRlXlatmHL79Vg820nqv1eT4jxtqIpyqJVvEmpePnsNcRKg9EBHvI
5zsGl2HWmQibQbZ0lJ4XM9rEVblxrDiON8Uw7AZbBDFFS2ziR5/uXMmOC9vyXaWx
3WwgjgSUpF5XZS+qprOYoYUB9XUo/QjdNL6qKYCNVfmiBhcFduFle/9t7L4Y3Q4w
FOywe+Wt0t6E5JbmnvDDbdtU7vU3norxfVpL6gIfJ9iMXprrZNktsLs3tpC8H6+Y
BTOuuFZtuFBqUMx4zcqjrtYTotAtCAyAMiDRhZUSlfJkGfajwMDPZSJDNRcoKIvG
XfiC56fUY1Rxp75RzXZ7cdbLxp5bEkFxZb29GSasW54RIuWWcAjSGtQtK8g9H3Bw
tKukhmA3JjOh7muSklwPDpfr9aM5SEBxHNWxgkw722TEv4DLA9XAJ2+ggMy5483R
JFPZQTFICqxRbKz11LhlwVho7IcCL7mpnfIMG4EYDVHC8W8n7lrzEwMzSU770AiN
lpELgD6rp5Ojy3xfRCxO6OU0cbu+ONZE8xHD0yJ45aTJtSfY85b5nv1akPZ0wfuo
zVh7AjGsoQ9DXjTjIz1PBUSk7ii0ESGQj5rqOQE20pyqGXIqetXopctZ24e94iYD
+HFO5AfTGAp+Ut2+wjnyRL0xPADzjtYP2DFrQLmdmOj3gU9DRJBURLUpPx2hy4ak
qCXjPOjFXeCSR5HNSmgNgW771FKZ4OS7rGUArK6FKZCJ+HP+h3G6lRHOlO9UWhdp
Qadic33hSvYefFPplk5/bG+uPg293ZElEiy4Et5EPGJl7CLcHMGVguX0W+cokXVA
gNJGGFeYkkn2/euFddFsB5dnctxy6MYiMkR/26EOszjddsTsDem1mDK2Y56v2La/
xGUIDThhLKE/nJJBX8BsOOl2dlMzNXsKMBA1M37gV8Y+GbX0NxqDKp2iq8zRmhKq
BdgQJ5N9sSNTn9RUKG8U6QiwZSBr0pLE3hrWD0eV++1YVnX0pDIUCTZYNuCjuQ/D
Xobo08qbdYar5AFZA13fkm9sHaAxpfXouppOMCSUAb1pFxD42npa6KN7Y0YeovP+
9ReIylqRG0sUaleo/ejrgupHXA7pvIyTEKdahqFbvO2Wgsudx9eS6oWAJlM7jMFc
OCk37LWDDyZIKlh82Pj9gIOZOHsux8s8AxOYX9AqQ3MjVvsQv3Y/SxkcwjGz54Gb
1vOUE0T4MAdz0XR2Qm2wkL9QKesOICjXfIBLz6uU5TtDce0HZUmB81CyFQRg62fZ
Vpbk+x8THqGgDt8JN55rdTsT/mzIX2Sa1oY9T95KVE1TlTbSwbxXrmT289iInOmA
pSFGY6cz8plY5tTtfYs+6z6PYRcXvsvTImF38WWY0Q/FCp7CPRO06giHnu4yt+9S
w7biaMgYlBfgyBJ5deRI+j6FZjf5m9UpvoDuFqxXdP2Vp7KuIDeQTedRHBZB8yLO
tGGtJMtqwaFMJSh+WZkCKKl07J1zuE9n1lyLjxessxmqbj6XCrWOXuaBA3q9ser+
GAtvdGRYSf8mnsQI3TyTIy3zLhY2YROc0DcN9Dy26e2EM9KPp8wxUmCx3574/R40
AMfFv0X+Hz8wZ5GB9sKRrhme/nOMAFxSb4iKq2xAeG0D8q17IvoifzUyHq10Fg0G
5T9brk+8kanwKFKRE1NiDXmA75FLd62gH3yjLTfa5uTTcry97dp2WWPbE9rXNBby
3shu85mOf9UCTtLSxR9yjLuUfeIdqHisamSOiinbT84mYWJUkISLwBWq8mjEzVJa
DYtPpZrwCvveNywwVRDtnxx4yd2p2t+LL3X/dEZaFmn9xGAI2VAfGab+dt281VB4
1g3OHzk2ReFt37WmjmHbDGlaaC9tbN3YSJ/UlAiXUAGS5iwurnK58m7/7xVOaBSH
BUYknpnDsbd5hwfZ98ThOHhOrLsrVY22151zYo0UIM1DKObQ8UjF/PfaH3QTGlBI
okL/NLvXxPtFYQU9zj6jDLfrnYtVaVVC1HOf4TXOKUvCXVhjRaBtaNUIaBGTfRAQ
3fls49LY2r77bGIdNcvXr+0s48OCse7C3hXQztgkcAU6ZADOqk2g5RhTkIn4P+Wd
o1+WkKJSVux2VqyLzTVvxG8pNRhx2FQkFqeFSw6KRHiqmrgghAE6moiiQzGuL0ba
+STss6bIjOZBaT/rjr1ICfSZZN3oUOyDzYlqRMfHfKgcgi91EQHezVNWiW3G4ftP
5XZkuD0UMae96nmmJ/CvO2Rr1ZwC7zasFFi7zj+O3tPNkwUVpuWOCn1g+3EPbpGU
qRUrORKmef+YWiIPvCOcpvdNrgSfg1QCeOuZdQbip3aE+8iLRDLjvgV9zxehJxlI
cX3HDziIk7PDjbnEeoEMa6dsi3G/gs+CUXM//Oe39h6pEJmg0c5YzRO0DS7WYPPY
JxbpuEqCa8BuyLvAyl9dLzt1wHLT/V049mPBckgOrRp6Je41Z8DN29l/kiSAnHy+
fFehV2IfwzfH/mVqPdaoxrUOqjtFEkXEXlUX5JPibyVRdH9Q8O/hdiy23i/tVJFA
6OI4ANj76er+aje1JmfLoKFVxPuHWeBhpBb4sC9QyatFag/Ch4sTf9ss6Hgfvyo7
DPz2erscx38c/uw4hTw6+hAHUK/AUce2D3ttwzEcOheAcLj2Szate5lufpYqGYXW
xtr5SfERWovJWlfZSaNI9BeWhv2TJwan5Ov4cq61Fa5+liDNL3dlW5gEOV6Rbzvq
rmX/6piBTD5piaiyyNkx/EgSR3hHqyMMbF1iKHK4BsOP/1PC9/oHoS/a5WZGApdc
t7QlnaG3iJtNUXM+g/vOsqm8VDQvu2ASaBoJk1nuKEO7nLa+x+whidy6L41774pP
xjkH69bopHr+8t5LFnBeg9IKeRtLuAfkeCn1f5bdsiAxbTILIPKTP8MWxCNH9ivI
biJjQJLnWdnaTpwYTo/0BLWIx10nCODmqWdX38wEnWyUcPs2GA9rLQMnebZaeUrD
RFlX+JaSH7fqBOyULun/PJR/5VeJJxBBKqSvxkiMku1AlcWAjlcGG6trEJknZq4i
tfUCJQepcZqucDQXSiow/7m4JZUZZktk74mEkk8hZ3EzFL67tlgoPcRhrgPWijwr
1p+aB+Ohnx4ZpKZ3HpeGSZu/icVDXFgp4Dqc86yLpdK2KbKVZAzleW2U5IBEEspD
O+TAGOSS1MzqhYKntrOp0VUUOmh2EyR8BQ51eBoeKAYt0Rq/wm7UiY40b5WVI78A
Eqtiy+wZbxJQEoQjku+m9K/KxSb0g/DQhbz1c0hj96ulGup5pFeYDU+O4WHzpoZ1
8Trur1SJK9A+jdHSDZ767yiHODmfVBuVZAMFsJzazd5CLRVJ/4/fqcwzLuLXpaGL
ZsgONPdJmCDE9NONnwjNIm3ybx++U2/E82ULDC4wSJ5VRsJN3ehwpP+QszEaKKZJ
/ZnWF5YKBcBZw3VZEwy1m7HpzJIovTNeVKl8Pw9UF1FZHBDGeD7+NMG1Li2Xu0b9
eKpUcddGaN1p2/g1ULXPGPrH7QfsTUUOtGkNT7+B8HL/fZWd+CS+bMdrIw5EhldI
Ex+wruZUdi4h/rqv0AhIDOGzIlkZht4eKRZ5cnXiugS7I3xy3s9HLxs8OQ+g1+mo
wxh7+UbHGEDIgTDQV8K9CddwK1Sg5UCq2Y9FhHn+hNyUYvHAYtdoCvLoJC3bmVGA
QE9/hlxrZ97tyLku/axXFBq3HfvfDUW8QpRIIvL1XCGTQeEfaSHS2bocD/ya/xM8
evhASRMWuA2NZFIGmlQujBgRNdC5xbRhMAtj4Z2Bu6fBkZ5+mqAxK36nhpmEf+wU
jwNQn2aYIyjM7zV5mPyh6xfS2QPrrhdz/MGDNHHcEiU+5sr0jUE60ihTU5JDLjyE
S+PS5NbV2Tf8WzYbp670f+mAyW0tfqoMl2VODH99kN54uZfCODkSjAtb4/qRtFJu
KujHX5K8v4kSyENqAO/ePUa2FZ1yuOkwGzOwQLN7VHxFGC2WKB0RGxBNbnfzqc8r
Fqcd0OBvMI+QFXYqsuIU6HHDU5RLTca+LntGfmie6IfjzCXgukLFCzq/1T6RA1D4
2URX2QGoLZoyLjV0zfFkuVifJ7UsiWFUY1FlLAwX2QzN1nyN5rkvuX5P1qjDPTud
StGcl7Rf5szCWN9mk6Bqtegg4XxAmUnCnwa4oRQo5MbLEULvdbwcOtoR2PGWxOD2
Toaf7POBve7wTY+Dj07irkGE7SI+b6v+yy3cytIN5IUt7xQdKAz2kdxtO2O8VES1
C6nJOOy19Q+g0j/jdvxgIW5K4Toz8AlKpXHqAMOxxYbY8+056kVvnqFynX19CvXE
6dZBW/5gssipko8bSJknBQrs85lSaL5P2vhI29xdFF9G7Lt7+blVXBBmfcWlwxYQ
X3KEm9LEEYNtDKUKQhmPzaZQvczIzUe/izSMR0XwFRqUlQBkaExDcIhENNI+VOmE
ac/+5v9wmZ0QyNOdX5wzX7vmykV+ZxkwljPIlO8p5tWgkHA2/tVTWWH8hCEfOAEB
AAsHxQe87nvP5UXBwMfBhmbzoqbPpe+PgJZ4AWQXAj8iXr53mfAbx40GrkUnezJp
ASnv+wEAhKqAXyJVzKg/8qNw5/oXNZB9rfiI2BXYWvPmg8fh+rA1T2F9/kPo3ZqC
6p6qsRjNMBUXzDWVg++bXmYsTy4YPE4FepdedgV/So52kfQI/nZD8ja+/q8q2g7B
w3TARTZmlCfezuD9JqQ1rafmYWIy19AzT5TUF9TRAsesDtiSgaGL4CHo3BtSgwtd
pBS4YY/CoB54sJl6wqJSD5Qu0ki0FxZWesCv//FUlxEOIY0Behg+2KdAy3ixxGJ8
T9hoidxE6/5NDAPRQ0vsu0rnpknVvXtkdAacpsVSl/XgumiMojpOHr9+umWn0oRb
LEGqkiidMYg83hbFUbiFio8SW4v7QRGzZIxB0SwIf7GDMmPdvtgvZ+g5u6uqqfL3
U+Exzsu2Qo7CivcbNdpIur2F9gA/SDYgw79m3BQ2xTxJ86B2BPmdHBbDomgk9lsI
JSaeydndbUuVQmT6DTUR1KWi7KJutNaBnWcyuSd5awg9HfgGRoBdXCSfPC5MUMBS
jXF+fqB5I1nYJYKrl7YYHm19ywNdHvsyoYyeEH5bb0xY7p9rMPSa70zX/i+StF1M
OSV7/hZsrge+D4s59xe5OmiOmAAmiQ6oftfZCQsH1+oTOXEb6GHXfV9EN6kNFbUm
5VCLOF/zCUGY2t/1HV1/deX+aDizFROBLvoFAItJjI+xClFyFBT3lFZ87k0+GMXy
MAV1ReBnKAufwsgm8KApAt76ljl3i5BVIbjVAgcyFAAqlRC5EpkLjXeB2Hs6BkxB
ksMNXIMWL/8BJOua68gtA1twB7/bPV9N5plvt399N/jWdPNmKU3cq3wvkdvubxs7
5bkSRX7MIt8nKer+kBPnF8v3pM6+Sm8/HEp7m4oDR9/4Or+U7Lvd0n5Yw/pzgpUC
04GlDMAmGd2xPo7oG5apb9cCSRtiAi6tRcoTdC+oEsNj7lRNcxb19rW1SRgn9IkA
PI9EOt42KSeldj7NQ0+UbP4FUHYxsQAVZKzDdxASmRV8LPiQ3cKQemgejHyeBuS7
JAV8PamBfXMvZeZ5bPeBI1XxHcbxQv41rh7+5lhAXw9DDNnxa47gU9HGzp4U4aYJ
nMkyHexq8FWAMH/63+LAeMVPrJ42ZdesEslQrLMrS1dSf0swhKn4UFS0A7osIQA+
4G1Em+VfhPtDjklUWrbBboZIcGdIEuCSg4ciWmRQ0Ds96AcvCbxFT5slgxNDKBau
vzcf0NFFOoOS/2D1TByTXFSRBC2Q+yvw5XDrRJm4wXOlGObY9fb0UkrLYd4BFrd4
RB0jUDMrw1oSM63M4DeDkBrySHTSm7dpWvly0wDnmLJyKpJ4H30QVTurxEDFRb1W
KHWoV1ySOQVDgWj1KQXmhoua4ITkcVDz+SgF225Wd46FXytn3tgJClVwMEmlngcK
lhfMHdYAuArFdRkanMVK5gNyeNWP2kzA0UZtNU3fS4zvA5GxXB5if1leWKSEBjJv
xal4UW8vrCR39JY5PIpPcvEKPCl4ckzBTLClaJbkbH1OhlXrxQlRLqAJEhgezM/R
5/Orvrh8oZB8Zgi6RCOkbe+9YEbsZWPNFeWtmp110IsH5hOECp0IkcWHH5/hQEwo
di5Upwt4qPWmUMgiTgF15dbWOf22kVUAV36VjyVu3ioAOew1k+cCt7Aj4CMnHaHe
OAAZu43a6cWe1Wh5TEKO8AYv/AAw5HAAZARBdPTlsxL3pSaFNQTrp429PiuXPP3/
NvCY72kf9+iuxRdibDJbx9LI2figMO0AOK+FX07j/ob3yIIrux1ay5Dc+24hRazQ
TaWB4fQ6vPfGx/s1KsPec+QzyUYwbwXZ5KbKqY11fw901v49s2uQ46J2rUaF5wW8
864Mut7zkkh7jUxE9V46KhTo9Ea+b+LiOp8wQYRSUDnAIjgQSv5wf2lGFwYwgLqT
cBKxyH+LShzTRd9ewUir+bZ3vv6lruqaD/rKsxGd+XUIK/uKgvBx5bY9uYxYB9rF
cdIaQc0usnWGkT+t1Vt8Z9zbfltHle/E+k60eScPHKD24cDpBiRUP8dB+i57+5VK
PCQngN3xKVeYkxQpYCNCciJ6sqbSAE78f058oENvMOcwYmmgZye3gYdz1bOKJu/j
gzB7ppINBSYwUoye3xNxLsKnIeQj/tJI3qJqaTLtAwFr2XiSHFyLA+ziGoh8xeiS
WuJukaQk8Tp0Nc2R+a0lZlnehgrJu1vl7WS5hriBJSsDA0P1k+j3zLOBsK9Puv64
VEcmsepsF6nyuyDn4ilheoJkk90WT/cRkm2R1aG5H7QULeSag725soG99PSBH4tf
J/8HeGGe2fVBskTWY5td/rZ+bNSNqw8douUPYVcEONwGJWhB8Y/lMtTk5r9iRWpz
G3EwkEjvLbLMjWwunTEGl3JAl7GJEMgBI9TdKhjDENwwo8BZe+LzyFEw2TOy5KO+
6eC2l3FH9N6bFTlC2Fslvs9LGchK61zX2gzOMR2lWdXz/0T/lcFjTSaBk8bbnalv
y7cfbMyLHgfeCUOyb5L6zDutZrGhDNKzxYWaHycc9Hdb7kSQcOj5mU4NOk3+KvJz
6gw/oiKloz7sZQpCWSqFyx5UTvYoUaN9ge08nOpe/K4a76mLdssObiSwCWD8VfrL
D6+DVukQWQTKrbv/qbj4vYi0GqRv60hcXbY0ekARwkVhirLIwNXjKxq7ozCatPCV
LyIIm55T1rbgtlODjjTOFZeUb7bW9sww59WMJ1GqSe0v3Benrfh6qCB3CvmdmbQT
GyBhop7usrWKqIHYpbTomCjEKoH2gcz8JhxpkJDgFbGBs+wkyW+SurKUmPjuaygv
Xrj0BQ4YzOeNYNY3KGJOoBc32JCyMg+xM9aDkzPb6yADva01sXutMVTemKZKCPrO
Dxm+kB+KVDXtQEVlpyD7V91p29A0EtgPcgNBMUdx388gwX5ymuNTp+so+lav5nZi
X1Ns/PHKupP72Emh//xAREcpXLZYYvPaQN9hRy0o7thkGEP7DenDlkQap9tQkPhA
BKspa2tAW9xivi1gtOxJeBkp0LQ6hhlvASJJbKpDK+6Lo3qgY3c5rbMHhz0XqMYV
8o70txXf7DlF/7ANPtKA2TM494tgsLJScGXUONnBWNmYAGApuDoZfMc5914paK8o
w8SuKIBaiXZGF9g8E0F/FCr/knlL5IrJB8dm+v6lLWPkdqbrGJIB10Jz9aQT/1RO
ZbmltzdM9Numed1oPQV4Hc9d+HvXARBUjMaSQSCobGdrszK9OxflVEHKN93KTT4z
ij0SdWQ7HxvZFI8ju9mHAp5RLZhXJeE8gf9e02q/fKOnPggWIhdCnleysQ2Tzw7+
0xFtvb6cyT5fVTJf/0TyWqnk/+l7nWDwq8s9W3Y+/K+/ejvw4oZmUi6MF0Sfr5ZL
uvco4HNfQtT98naLFpGIlQQH+unqem+gbrqu8UW09pwP8ONeegLrooVDXFcTguEV
e+5CUEszutwJW49MHWPQHX2qiL8/BBP/8oZL4/Mx/Sp5AaPjLHGWzAnfEkIxz30y
opR3KnwdNmcwkr/FgJhbchDKOL8kyuRW/jjVIHb5+8tg/t+rBkwomc/7018V4RXm
6q+jXb7QYErQOtcLQpocxDfgLVyl4th93V0MOH6+uRyMx+aCracvBclBXpPQ+u7Q
ZiMy14c07EKjYixE3yQcHdev+MsGgcIfjnfjmMqs9JPppZjnp1aUM/zZ9PdQpJtH
qKmHfKnVwq0eCq8i8je2xC/oQ2pgW26ZEuO9OOaf6wUXKw3ztMsLmUywpYRGKUUW
SrF3oAaJE2Y+OsBBGsmY2OFBX72hnuFYACqLZWbC/PtFCJC412ErZnZXmYfx7IWf
QKiPJ0qkYRxot3DW5ntcToaVn364WL5SvNzIUZGpo4Jx96kM0adYFLE0rymULrjG
za/HvmMSZ9x6DX8hqY+At04l2bDhgoatPkXzHjYvNIJC3eAYp3juygxBUC/Kp9uV
pRLW2zOVVGoF4KMdyT+8hC5d9OgqFEMN+HmYR8/xmfRadtu3ukWKlJeuaxFNwZBw
p8WwyjE+b44iuAE4FvA/nZRHBMdKmLdghp7CzbX8R7Nh1Rs6n8bOY2j37XMNcuQd
o9R0l5qF15LbgzHObdIrKNusJg7Fddd2AJqiO0SDjoOdwrGQzA2kz39bPY+tY9BV
xQRTUMSVKycVtWIitcperbbqCdOL6u71irZ+T3k7UqJTV5BVCyVs0BbKYiB3BwxM
p0G5hZvdfJ3JVGiYS+mbcvdlNdZOwQQ2KI0vluKXu4yzonUes/S3/4esDVjuqLL6
Zg9jkF2b94PP7eVRJymD2+pxXSq9HZ8v5yT1NUkOraiL5070MaJlMIMaa8cMwrzy
4mP9MRFki1pMQs+uNXEMjP0nCYkcxistzPSP7KF9jyC5d4fCaX4UrqzKnb3297f3
KyAGL7KhEGePzHELiHYop29P8bEoXlwJjfL+RwVoQv545nxTbbPnHVFf0uh2AyuX
68Y3553w4HgVLbfOlaNH60RiXJJi9H0dEgVl2mRxMyzZdrsaGrATAipe2cwOK52S
C1V78c1hg1V7tuFWXToERUB1gD+36CTlNTM83jHbPVWMbvrYl9ailKpcvLnpmwCl
vfrnlewNOPEE+uQhoh2QezydskUID/4nDeWHSbu0X2M5FsPViGzYwZfqTv9Cbetf
20y5lWEwx1FZAo8ALcDI1VumL2GW5+6ho1xfLL2pDW6l7xuUW06QJoOYXZM14oyd
zSgJGPEsZA3T9YJbhpZnrWl4tAAFc9CtbdAgzI8RQPNNpYtlvIGe4mYw0Yw63w0B
eFJx2/yFZKayMRVKFyx6EUOc3vbzBiK8HxxuSz2V8Yu2WuVpUltsw8U+A2UhbdV+
/cN1mLmST3pHypauRX4PutgONZRz6LptBhZL//VHcEB6Buar0dRQTb+0zkAe6063
PaHnqoAKy0Ka5rln2t/mGG0KHRJe3OVkmz+jqi2XLPFXZuvPBGJn7lx1rN5y2Gz2
dZ4MifeY0MrpqJRUJwLh6rL2ydrJni7uPA4rD0VWrZKC1IJMX8qNsHgA6NCZ/8kt
Ru0Oh45liriFChNdjl6uk/bq/Otp49SYXZ1vqHeJQXhS/qkURnBi5c5QXwbnalYx
w8GY5GW4MJ4VSJB0wS9UB0r/MooNwgm8oa4A6ImspdWlI4Q299OP563qx8EenSAx
6neKy78JxRapRScOcC+WLkdVe0n+KKlQz4D5OSPUutY6HquzAGd8eFNwx7m1NTc8
2qgh29rNEqYnX263e3M8YQXOuCkQD7pj3Z8sffVFgIgfqShaPdmC6/MOzc7sMtkl
8PlfK6MkaIUFWrDnur3Fm/LbHM1SJ+2YI5WUt47wV/1QVTxf2D9mIgXA6EqcTOdC
ZAdL7FHMewTqKCy9+yp+eyiOswkjEedYMzYn99gWb3TVpAAiTRerbrZi3xZznU64
afeG+MItBX8SfdR/CXoOd9Ce9mAkdY67f8zN8hPCl6FsYX8WW3wiQb8mt2mE3ltZ
l5q3z30aJs6OHUYS/jUVmubr5ONBkmcqVyZRPErRiVkyTI6Tf3bwcr9hLpDhmiqS
2Oi21o0xBsJwxPHjiKJHL3IvDG6xjYH8ay0NE93L4ojBBUX9Oamgin96wZNYmYRd
dSx9mt/g0mimaGl2nJzfVgaD0IQkuVuZhUZsiDyrl8wZRlEcC5xNA/b5zF3OD2Y5
bHiovF7qwShZnZapde1akoKg1OcQ3UxUhotMZT/ugvfBgf2QcF+SJwisoqol2Bum
xh7KZsplVqn1E/bDUDoE7NKA0IWClpp7jlmPRtacI0/QhplUUM9rjSNfiNKk4ua3
4/d86lnC1GAvLK4/Er4mvaMMSjROENYeXOaaWuvx7GpDtyxg+cKj8m6CfzhbVJLT
Um2QBO0xbz1sS+fXmFy8SE9/UtVMw/auaVqgusxUlcfeEYVaf75dgsu8Uc+Q+gaH
ASM5v00hoQ/E9Riq8lErkLOfJE0Gsge979DMTrnSTyCFwZD7zea7NHm8YULFvFxN
/8Om2bgyQuB5UAHhP8nG0tXm75/ZkqqGAo7WT1p5SImpmEzpVaUHlVHgNEyB9GWO
S+HjB0v20IjLG62+n5ltX97nk4qe5gu57q3m/EQVMyucTxTG/30Hq1X+qk2a9kyT
UrKC9/Z1MdE1G++BLBIaKoHBu09WaAsF5czbsH5GJckF95nNGR4DFb6Wdyu5XyrR
Y7EroBnf7lA27liY8En1bavsB1QeElnJFKJTEDOnGU+CFUPA2BWf2yIrwgGP9ep9
Ityc0WLBoBDJiX7hp4gFvadwlB2kp90jOTsPR6luHYYZyHPAQapLxcwljVp1Py5V
T6FWnA2+JZ571FN8jmz83xnwTU4/29cSsAMKslZDipbyWzAKJ2e9Zs2v9wvYWO5g
dLZ5TX9tn0RPid+iA5ChgGT9A9d9xrKOd1Wac36aTOCshRGbG5j2Tx9TSeBN9KgN
JKaQw/yolFJ7d7hjAEGEc2HT6u+IHLYF5uomQJLTAXUTF0nSZe/FrhP7+ErFrgEY
nV1JP+lW8MmevacfYMDjIJxrGTSEnSot2ULDPZLUYGB8pMWaeN6jgRrVDpVstex1
xc9zSkjFd8sL1sZlWnLfQXzEBjrcER8EfdgCgFhHZSYwczp8JWGDx6gL8KiLhXsh
L1w9Hw2nFEjV8m+GkfqgG9H9sMBj4c6O1av7i2s6ltGb3MMT2QX6T0zPUF7UCJ0L
QSlgDl7E0B5ZINlgdIJiARTnfkIHzZ7D/V9HPfnCOEhjkDkyD1fv4L0rbytLDsKm
7IgtjCFLOuCHPmtva1RnarUpySI+WImZwsDNagj3JA8o5Idf32JAmyUqai+idgXh
zMBUOd2Y5rBFs7BCL8sYwGM8fWHFC1O6f+EOe7mbJfCB3NIxUKngK6qULb3CBoKG
xdzyiiMY1IJ4G7aWfSDOIYV6qDab0IyqFpLGLjH1AtHccUCY8V84yjnkoI8N41mY
6As9q3EpJA9blg/Eilyo1aaYfFahBYvI1Dvamuf9voIgGZ7CZflHT1+1jPP5CaU6
/KBz49UrbQMMNxsxtMKpFFtMTYKe9ciubV43rPVOSsQD6msDGmxOT5T/2smtaaj8
u/BNNh5sfiY3/NM4CzJs0Xhebydgb3T6y6aZYGzrdVOg4fKRN1XCsSE9KraoXIGU
EgMJl4aGsnJ1vbNf997F14yeusuZm+HPHAHvywrMJEm6ov6TjtCy5FlUTkZectIB
DxX0l1isQqKJ6TAdSsy9FTyCi4wrHc5pMJwvGnsqCuSMyfbo7aaWFR7wNoXgm8Ip
qsY88rdvkndfQ3kui48l4KahU6XI0iJ+JsTEqiIQ+i/0KKPwKVzZz65JeoGlBVZb
pdXhnOrvAvfpctqOImTwGLztSp2f0Wour3mij2KcV/jLkuOdEwMCTa7iUQHN+NfK
5OEbeNtfZlQteC/e1GB3JjnNxzWr6n1kOu6V7dgSPhwysp/EZKGDrk06RP88arRS
BSqLkr3w1IRaPoKZnSdJhk/o0eJSdAyFHhgGSYeMBF35KsGhJT//i2NXpLNWlQeV
h5aof5VVFBIU3J/7A34JpPfbp5IKPwsH/K46C4adEQMVVIjd7C5UaEdVjP3Cl0QR
jhpAJbrq2GxsYk+xI3eskGcmqyv4wQMkjoVWeTOUd3evXoyAwVd5NirFkBcIFSpj
8lt8GMHck6DzL2rkFRQJGpiDhrCPmR/lv8+gjR8ZHNKf7J7x4q2L280N78prl4Hv
bClGgjXD1aSsAz7EhbZ3SUpxjmD4MM6WnB1KYIzEM/izxTjlRgPL0FVUzi+u1EnF
ft3uPtV/xKPmuLR6RXulq3ZHNz14pwQZa88lvG/Uvg1DAAysKwxm9UpwC7d71HtX
bUWbQC0OsPEJQomgWJ7u8Ied85G+Xxf2SnedascGGbW0jaKqoQn3TW1OzqAF58Gz
vxICGhljCrysiKa/0Xhw1xXHTWD9SkSzdxPPeETxi8HXMII1nJ/ul8ppq0LebRUH
C2NzllXTFd/pjhBDE2jan1w9XnaTNvQld2Qjfc366a71Kn71ZegQKpQr1ZT2HVel
uLxmxmxqNeWr+/EPoB/K0ZFWDg8xA+IOAd97jq+jhR3oHCRs0cb5HATHiA29DVqE
GSl31dVxd+F3AnmtjLP2wguLklv9stZCi10mQrEzPYWr5hgsz0R0OjS2Ut9rqiNr
Y6H1kfJ/GhrlFiqB1rQWJGJywGv1O7Zn2Z1ICpUvtroN2D6PmNlmisc5Oj4Oryci
f/tma5GPULz4sg3ir9S5KJsyUE1oV7jrXYANOnQRmwcyg6QW1bFHxH6YIYv3v74C
PaO5QQ3ApnhAVaX546bcNRg+tEkt+Qj8LrXrKno71pYpFEJCrdW62zTaI2GyDIvr
BRNJMZr3ejNqLOyCTWHN8KqnCoCVhRSA8gw567ywBMICEcBQE91PWkyj30PFap0r
jHPUfsXLR+5W7C1HR2g4hQfULRIwU5OMt/h3KFlf1wJILdYQLRWbgjzklRz14Z0L
yGNo3w8xkIFg0OWwcFa4wIfHU05jY34j3rEFMcGNy0aV8QdLT5skMMhx9cYDPvaI
oLcob/oAev3nMNIzLMq7ZP7SMddtkrun8FZcaI8ZXxFTR6BhGAOCTZi6yhp2vZOv
a+URgcxuA9HiOzqvVtC4t3gXff4aPiDNC7vQpAjkTQEXAaWd/EZp9YjMLYXtwGbI
45+xRNZClVulGkJpYvQt/CxqiZ73/lffgHZMtAS+Hg0Dxl8lGqgd8HWR2qn45NHT
F7shSCR3R2sYzJjtAJ10kImnVjj9sCuUCWN5oK5eBmkCDNX8yGbkX7IkSde+Q4+R
t6ooIDDg+TpiIauwm9xUSAOhXanBBJ/yqcOjB1I3U8iywjO6+rYwpF1UujnYo9KM
mfvm299qITDIya+NLhWajjliweA11BS3kslql2uip+ilBFi4+F9YOwhPQJEIQFs8
IynIoG4u5OpGcSHJu0F3FR7ZmuwvO9Jdf1NuOVNToHx8/b0vnJtKym/9Xn1IZ8PW
/qstV7O1YEBTXk7v7kBxqriNK1EwVQRSF88CJENCO01J0uomNijraOkBKtKHk99w
GkiwPSpoapS2yM98R+RTziaxtdA/m/Yx11UTQX5liyG9/6pGIwVQsyc01GRzKei6
QNmlsr4ozlfoPNzxuXln2I2tSU5owPkEBMATCiD2ChURDqZZHTi5Jd/RNQFnEojP
H/Rj8yAZwGY/j/6Drr6nFs9gOPF5YzxW9ANZL2K7eM9mHwS8QRk/E7TRTYtsOt6i
Gh2exX0Cy62VSA53DL1xVFaENlbJDDhi2/weUjTA+YA1g6LluPWD0mO4m4qs0dgw
dckBKw269ReQQbVVou0pBQjXoZLtF12WYwwI6N/Ne7HJf1LNFOL2s/DVJ26mQmUX
akxmIUmtGKrJgxqxIK0x2boPGUUGUFBzZA/W9V5CIP8XRBcgWS7OPDMNnq2J9FdT
iQMvURp046lnDvUUgBpR/9C+1KEQmnEw43Dq0NJyu46iuSXWY41No/zoBWwQcLmV
MA+fUkft+BZtdI0CzAeVlyQLRAQ28IqLD3hwj8zWksBetw+Az940rjWkYemt1Nvp
f32UQ9Kj8DtIGL3/Vr6BgDNWKyAuPAJJPd0D/iOAwmWtPnL2rgZbGrii2VUMJ3zh
VDXVgdY2PrcOJ7H137Rg5B5FopzhNqB+h91l1LAhcD/GtSPeHg9Cvla3fki8jpo9
+ZyauGRakGlyiXDViyQC+JHeNDClpOr6KfAczrLPzu6DfxEUlkWH4R3NKf6dC6qU
eQVHcT0vLCjxHjhCL7tXSjPnKnBawG26n1ddHPJXHSFPoDj2IN0S3imBorsg9K6y
DwVmIWDTnE2EsstbEar7XufJc1wS8Tp9HXDNT18ezCLZ6wPRbzcvh7OCc6naKXow
pYzOSubi5y4Ha2x6V4lcELAODuOLed0Vkaj5X1oIRO1NpeQ2vtaou/ljN9nj1bVw
Ics0smzwu0Ojm4qmaOinR8oHey+U/SYNpqpngLyn7CsvhCeA6LAsmIqRZN1PdYLS
5ZZMefu8Ibbdxs/ZQdxX6/rhJSRyUS6VXKTmmg+EqWUyMCBIRSUtkeufhotTlvwa
SWc4ZttCf1dtM1sjoQoRZsNh1KhnHNHiv7AEg5V1/CGiXjVKS83tGFB9z89Cd32n
HoRMXIwTqz3MydPqDOs/q1UOxHmWUI+WF25P+0cp2tRiIrnPF2N3CGaDttlNBMvW
KJlFwckpsYcBnpKxaMuZ17Jdvdt4uDdC/uapJ2HuWRgv8/2vOJ1ikYrXjGBQ/Obs
okSavO92oaSniLMqYvb1Rw==
`protect END_PROTECTED
