`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLA8CLLJ8Qg8wsf0/k5ZJE7jrYGrwpubMOkK5claeescox2RS1h72GnncINsrHj5
ZZTa9ugqCDTjQndvf7XgAq60unQqS2C2D7VHkidYLLPe8WrWxgiPPTT6I/thowg2
hggua3VrGy4XShnwx2F66IuqU6EDvIiQ4foMHYQyJi53gfEUqye2LKbFecg6pv4b
BalbLuxdO/CQW2+8jJACRo5mp6ixWbVA5Sij2HhcB3L75e7VtoMz6GdjMdW5tpXL
1MzAzNUa13qBHsYShiR7Kor93my/Clcw+Fh7ITuTyIEzv9fZk7rqpoyQeCm4izdq
3sAxqB+/61zwxmDdHgr5kLkySyAkjR697tG9YpZaFqiLYIju8x0/Hus416yYBxBm
d8ilxiLitS/9+STSr90pgT5SrBhlauL99/WyemovTTqSAtpJqPP7xkLj+TiU+B34
MvXZEPLVNhrjlVzYxhosAia1xAJiqcQMe8qOaxw1i1pSAun7VEB2j84B8Vnc5vaB
`protect END_PROTECTED
