`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A71qlrTvvBLT72d+9o4OEfg3onAmNHXCQvBQgmjybgp2V3/dlCTJ8b3QCKvP46nZ
exhgbRCQtswnL+ij11/5eGZfxvZxZobPj5sbExVl5IaC+PXEuLlAChSji0aV4YG1
MXdUdg0nds1Wq1SS/JOx1+Ov8DyxTgWdKoR24KxCCalrgVd16x2+bHjULaC28KJr
rGdgQEIxV/s0Y2rXBaKBHXVSzW3NZwi2OARwAt0vREdsomnBoMMIhslY5whXYh38
7RCks195teflFsZ/X45EWe5BvUX2DRNYJLsxhUWJkn4MQTKaU+gbabiR0mPRdzCM
gjEeU6sRhBgO4gJWqx9E09MjmcCptDQ1QuU5IMykBEsDIWEmAxwugMAaY5r5f3Wi
9Wdt4Y8gCHVgD1ldp31dLvUagLC/5gK2akv2EX4q+HzxfvrToLmqbuRT/zkNK8F9
`protect END_PROTECTED
