`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gSwbiAShkNUSQqDInhJssPGcwPdwaL1bXz7c5kW2dltIe77wE97CLruUkfMFbEQI
xD7E7TzBFFAbrT0dOwIb/glmnpuIKg3FzkV4EvqB9vDj/bZtNf+Q8t1QvjHlObsW
uG2bmR1O9uM/vGUVsMnwokiq8dM6+AmUJlSKdr0ENixzyJfpt55NigdFw6tOMXaR
qaS0eXgbOU91moZdsVKPw6ONPZ8Sdq+bHRiS7Locw9+HVc7to1HfOL7+ylSMfPrW
CCYqXzKXtZdpA3UHf7WW2VqxaPdCyrdQlC1zaWre9w9s6NU5UaulERTusl8iOdSf
TnAvr2ohjj1uFYNjCwmgFKQIXCcNu80nRZTOfSvLl4tloFJAeEKI8W+9dxHTfr8/
9QOjOnJ8UFlT41vvztLksUEX2CYzN4kcyFC7T7ssTsm92tCQhmndqC0TDdsl+xEJ
EEEgFmdG7YKwoGXubqpcZOWoKHw846gt2T+0P98Dr6mhKtWwiZqBZcYCqDClRlN8
R8wkLCDABNbdx2acdsa52nDw3Z0iJWl9EEdIah60vAKFzVeG3MXRJlHl3lJJEAZ9
IkoloR9GDrJUe9wtTzUVUhFv3JuKRdGBcO0OmyNPQHOW2BPzaA7WH/DM34MYkGz1
FI+pV/ItJzGBaZixaJ4+fxHusRPKGi/lsV6PzCPS9IiUDYNkgeRcZip3DFOMbvBr
BrzVHEW7+/b2NzqOeLsdvQ==
`protect END_PROTECTED
