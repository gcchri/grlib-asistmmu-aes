`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8FluiO49eLz9QjyJC2ZswbNIMrtq7tlaSSKSQEFgKeIeYo8KwNvsOqsNnxgxdd2
1ZvMsEcgI3sL6a2h/Dvs0MvQxk3X911N1XTKReOs4ziTHR8vW2/nJy+GBUUdNuEK
DbowJymsgHqC7YOq5dFYMNHd7vqKs0QNC9UBv7tHP2hylRoJPt7Pigi7FsXe10mn
EzQmUn6Y5qzIKnzs43HLpWtmPvGAp3lY43qhHCsbOtmmIXvDKmeEmOIKMe+QaqIc
nhcFL4c/k9ZBUi4HL9TgjfgC5ITsyCOXhvsHzG7dv8DM4YVEHN063OR0RTCCak2m
DehVaEsquyWc7ddk0UZkxaOpTt3C+56DSbM4VqrfRrb6JhhOhqpIkwOXPb01BKX1
`protect END_PROTECTED
