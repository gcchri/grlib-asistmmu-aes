`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AegnS9D5IPnZZo17kk43RIk2LIBuqU2IHsvF4RU1oevL1bJHi6VZ8/5tDRZC/Spd
ItXvG7AEvT382OJW2yUPKVYxhqY6qtpOSOGhyQeDmP4+DKgzNeJvxlG5xMOjKxzu
HHiQvvdNUq+CEmahHNTMBnojoxPyQtiAS3F3itlXVxZQZu4gOFfAFuxksAJkSkuO
N3kRRNAYf0x74sT89sd/84sN3Lh+sRzm4yBXKCH3yn2LnT3mN1n16hUGK8FMxI0e
yo79ksRovF9HHTeSyLWGRc3ml8AmBu7XwQY42MvsVs5j+EPvJxZ2YHFexuID5dpK
6UqVoT8ff9RD+Z4R7+I3Jb3AuUYT1bA12nfEikn+0xz+1jnqos32nz1fGe6KB5Gg
zOvAka2y8tTrwlcJM/WN3iOktTAR8ZOf7gbvQfJTA/jg6svqCYleXVknFf5Ex/oL
`protect END_PROTECTED
