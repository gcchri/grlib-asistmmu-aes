`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDDghTCstf0yriUD/M+BaEhaEcO/p0a+787T8QrafX6aZVNCx4xvUUPee5tOSN+Y
LK/zcVU9MlKv8Oix5AYWf5aZBo+VUhwsjNODD8cP8QIxYB6Hapsrscx+rhv6vuDi
FCM0GPPdpt+ItPDPtgnftBheYFFu7v41QMgJljNL/jaydap2UpnfHGUgg5NAx57b
jZ1ex+1xjJutwq4SsTrDRnbbUSeegBamWrZJT8RcQzrW0bS6kHTG1NX2X40KN2n+
hls+TmBRPuH2SoHmdzucOrVxzi+0g4bKc3mI53KfCe+JCIVkNuUQ7+lRnBY+XLTO
9rJNJJ+ZCBOGaZ4eXLg4iDDMglAvyS24g2QtkB1MPcXnMEiGt85VdBhiQ3WsuP6H
beHyjJmZ+2K3gKzjfZgO+1oCeMQsSzz2zfYbkvaB6pMMf0GbtMQdmTasMV+YpXzO
pAmYZYzGA9bPK3TpYhz9VHFeNZIDzOMT882mFfoEoe+Ak6/Ba+iN86m4DYgG72XI
tgKSkdeWXYnGR3VbV48KANmZfccy7YVyEoAQ6PwppX05ToQKjR9B+4rWdSTxa+3N
qz4yDXLwJmfVGFH5CAMSZesGZto4kHBskFKB9IWjpdvY6wF+XiT+Xu9Se1RhWCs5
pUMBTiec1Ng9wT0iti12Gx/izHMPabPBM5VwLQslVw1sG08dRaKm6hatx74p2854
ncahTx+qnTnZHL9WnbklyUEuGQ5XWuax167e8UPymQaSvIlmJjtwgVIP0Pv1gE1w
EPRYCNWWLOwvHU0omZb3hQ==
`protect END_PROTECTED
