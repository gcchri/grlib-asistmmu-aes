`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/cS7refdTQDesX0Kd9dxUOKXolrau0JecRL++slO5617B0VUEaMQ4XbZJ0JO+iVc
sgknjzshYMF1prCFB7g5s7SOWVgNk4Twky6sOyHGvTMD6duwxKLk1ba08ET7y5AP
fCrDoLYyvFyLsEKmS3BxEhhaevljHUd9VXILEP5VBjKtT75UoLtg9NEWVCBNy85b
KYv6gcn/v9f0vqCwZvq9hX9KaGVHE0XyIeV8G7erZt1ZLtFRgaMZjdspdM5bCPA9
yzngJCdP+ZhetnxwEJAtenEzlqKqwDO1O9zcMLeLwNNwXvxG8UhRU/u1c6mOMqAv
rU6ZrtlVgKLzqPBJ+yXL8L+qpfLhGhoDrahJPd2/nAXDwTcnBZWNBiuuS89ubmod
8fJi/gK633873mKCuoDJ3QTulNAzRP+3VU/eP5ll+Dt/2RAnB5BOuS6s01PtCefW
aDiGwX6qug8jZReBR30YrDm6pFyUTemBOL5MsOX8jqJOncSmipOW6uWqRYrX0XcM
U6Yh2p5RQv02CRcOcxPp3twTARgyVcwLtnjEDD54keo/Rh0a+iHv1uyZgpx2oMJR
TrFlPhGj9XMlMb8XQXYPfxrce4Makr7Ig9PIAYIHPUpv3ZFZZw3dldN3/I8GpNnx
whutue6Tx2xblDBKmgPdealFrakDmQAmlx5HatbKbo3slvmIA/HSoO3K5B5ptP5e
OM/rUzhedbZGY/kNKmyXgiPhHl1I2wGdpKIT0fkEqcowPp2CX5pPF0Zy21ZMlGBK
Wr4tJ4iFbsuJ4BPy6p6s4vEh2+2wo/BLa1GYVfPy1TuvNtSrwfB+mb7YNhQGmigy
7WEM+49jrl8X357w4XVQZ18mQqm8iW80R0EpiQN1oGP3bMYhBF7zlZWZgeptP1wn
9hdqljKLAqtTanZOJRnRUVJhiVcW+al8I7EKjwK7ao+ZlXohOoA9kpfECvIwXkRr
zttdqqeoMgm4dAG2GVw2ZLCIjdnz2Yj7iS3xUJ8y5EpL9Kn+H6x79BTlAtmb09oh
nJf883nDvgzxHMmwHkdAKXIz8+fnGdGgBV2Gk8F5srsP7T/1D7AxMnFuPkw0+LH7
yNVheccJo1mu1czpFrgFnlsvgemCsF5dbk6VBzlM4ameKwRwM0km6TPLrByCJkRK
r53VBGtsc0lfqry7RQLOq4pLtEWkEV+k81QvARzd0Rn43qemmyAyVJUSnq4KUzdd
NVAwgifqnr5UKORhGh4BAyqIurnVci8VrrD1BHTQhjxYSPzhZVBO3yQcrFNYlF92
RguWmHS+0jK2xEslfuBjXe/XuTCiYFL66ResFO1QNuHtnLYuLVDRiTmcxRrCE8bN
nyjItTUqDdzSmJ5UN+sJ2yTvHjaFQVxPFIxelRQrc2vhWEz8woQjdwc71OAkFf+B
TUH4n3DC9g7SMIsd1GOi3gKl4JWGJ2DtqXa3n+0RGaxSyo8gMRFu+Kd1yJjFhYdg
o0QZ33XRgC9XwORXzMrEDxMgP83qR6lJxqqUaHbAoMiFb/W6o3rWbqkDqzerlXND
jc9/mPDhxkO8W0eHToRpD63EpZ7P3apEa0jFx4g2SVwNdiKP9SCf4UtSxIIq0r1k
+KnUHYI61gcp8zGpI8K5HA==
`protect END_PROTECTED
