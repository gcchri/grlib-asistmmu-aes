`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0CaJ1aVs5p7s5Sl4J8YhDz1l9N4sEI1MulUob3i3oz7lC99mm8oxgp7phyVjN5XR
wva+Ao2E7blqo43FLQzgPMcxrMXsKgQu+pfJI+ajbN9ywcuToPV/IR1avH4TfT6x
Z3d0GgNQGaORU53+p2d9Hy0WhnJmLZJRywy5258KFSdN6L/+hfX5kpb7OfcaHAho
u4unGwlaN72wUhI9RGkzuSBh66p3CTY47XJVIJEyqOz3UvSqC9u6AGk94saR3xGd
9m/ZCW92nwahN53KrYTvATS1dHvysNg63Sg3oLZ8OfbTARC+mKLmWkHyG89ituf3
GNG13snFWlQEy6o8s1+gdRcDUiEoUyzKtmvvS93tw2VUSgN66Hzw59eqkQqBVGzr
bZueKw9/s65+tTX6OqzrcyG6cJg6vTivdMESMBhoFETdB3mJKD42Mw56c+PTTOCP
IR/Od36lgxcq74oYh4z91JAbTfM4KdyVVPW6YLsDuiyh5/ur07kt5uJP5RQ7FYbr
0L6yDtSIiZKtYDf4Skw1JoANFcjg4Ec3glqXmyV+Lo2BM49s+Qp45xuWqa97rQk+
ORDUHT7etUovnMDii3DL6R5crDMgte/dD5iljpEWIRkrLxYTfG88HAAwAz0ciHmz
c1FxqCQwBLNZS3JjO2mmebN/UXw2YoxPtRfS7c0dYtrY54f34+wWKR/cf2dQDQjp
PogrxTQP45rJIrfTZODI8o5kCl2Pe6ShtWbU0CkWT0+fwWoc3uzJX4bppIMogOgv
YkJOv1pxaHgMCC0B1UjKJcBwPX5aIBIlDCohKrMVvO7mtr+vCLsv+fvojR98XwZj
PnHr3AAgicFrkLPFpGDFq1kUNWS1tkEbBM9IJ39OsL+FyfmJyAy1jWtaqDmJ5Ayy
GjaChVZRz4KntkxOdwdPXC+MvpW2nxuSlpNcnR74asAXmfkse1YRj0MwlIxNEnaf
IWiEZlGnLpFw8YY787SVjXlxpdRHGcp/aun0lyhVbzsO/JN6IAqIAimC407fompl
AoXjUCVhfU4Ab7uhuNAlIeOe9up23+eSceQu6PxYehzFMdd/IJV33+Y4scAOIs8u
FxXoDK9ZBraqi9jntQkUpIIzgcwD2MKvCmxvwmB1RDiDcDXJkKU2iybCoAdvysIe
h9SeMpecZjWaaqXvfBr/do3camZJuP7f7n+7quYgbi6wMcAZKb+cZqu3tYXMsg0G
MRVDiLPY69HdL8KS9Q1/lSBLo5RSfR7Comnao89lSVxrBbb9Z0e+D8ilBPoxOk8p
`protect END_PROTECTED
