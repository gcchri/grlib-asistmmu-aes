`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y3gOVWiXhAK895HTyih/Hhkr6TBqluayzGnx60oedPVB42MIGg19ROt8pR5mRVLW
c622nJJEdbZC5Ttu/ppCHgHfX5X0M0SA9ui0LDnGm4/N6dU8OvDK3VSgXTJ1phdG
EM0GHZLlnzyEi4CMb3RLFb8SEeVGDaICyTD9S+06UHwFESPu1GmY2Sjz3U8lOQ+M
QWhESAgCBJhIIoLEh6yl0cHiz/MalEl23+RoM/z9tMc3+zK8ZzdKNnCjgIxBZ/TA
9nRqZKsdtkTMzlKq0IjOFcdSytWyBT3LhEps/5rOjBqMBagbnPIJV2RpH7MQKk9Q
ue8yhFpTg8+ZbcvSsdIAwt4WfVZocgsdYVTs7gjeNYGVCtVdsCvypvmAYYo2fe3J
olgSfvVRgL7jo8SbuiaYfUKlOeR5C+dgjxoCE7pwhGEVYGB/k5n5F1Cp78NoVWBE
yQ+VnY8Lm4h/3j/RM/RIekl0dr4jsOKeuHAak9DaVYORAIpMrmxLTU9Cbaeuy9YD
eo7ZOoarPlapZOKZTfjitTETEDYSfvpcEkfo+d+eHUufWip74iCVFjoJlHzPZF1j
oyeXMmkQMhv4nygGxCfRJIBuPDjvabMcicmn/ifSDMaih5eMc1c9hOMHT+Nz2g7K
kCj+idXC5r8YaS8Q1Emv61kUJlYnE6l5IfI3C34O+m21OHDYphJYEegwrNq4jLvs
iOdCr+lO1iSDRnRzXwBp2kMbfTWqdayA3WDcPU62q+qIMrgypSCT/vPYUVaQ2Y9n
/9/J+E1ix8RzXwGETSRVYX/YE/KQW8N8jT78qme6eow=
`protect END_PROTECTED
