`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jus3ZZuNEdEmhvSjnQX77hRxgLQyDaMSX6YIUvkQ++/bz2c+qy9oqZzvj6nbtzAH
WFHTbtu20oCc6ptgRcYLaHxxVyO/xhdaVVwZyXQ7VEyVJfHG+FPomV0KOlYSesmQ
ovx/l0ltUY/+164ntrm4F3Ufbx6ekTO34mMVig2IdcdIHc+h+XQ1kBOc0q5uMk10
Y6pBCvgu9hohEyYSClsYWArjbDq24jylLD6m4AsWF1HPbswS560BOOanZDt67yIj
acLaaoE8871VYyzYI30Orerq0X6GWE3VKtMLySeA6xxJRfqIGme65+EHjmBEQQ9B
kBJ1eotf7c+BK11kM6DToWoFB9mKjbee1sSYGeOjGhj6em9L77v0d3IoOjCpbC5+
OoSb861KCyMlfOwaVJTYAkgwrISG/s2rB3GNu+VYQtKDQoY6BexY4NVEdVsFW05r
EyrJATZ8inc7qC2tVREmXGVhrdrf0tYOssIHljve6Yxd5tpDoBsAccac6I5kGTFF
Ze4j7L04E86xRJLulFUA7Va447V/JECvjmeAjYovubQV7zaVBoo8+//ZZKE0+dCl
eZiklKvEcgIJ5A6ZqLOZ5GCZt9mqKL+vfiGASbPKXkh0Bht3snfqOI1qhltVXTGP
UE6brDMOdyjyxZ5r+oykoC/GURMxpJrzuRMawN1Dlsgb3MgZs3UuosbGlFxBtmFC
zDeM3pqLqSmJqnWD38xkAUERJ/vx4KPJcXPb/3k6NtErG83Xg7Z69NiAhNnDorR2
Ge29sqgG/ap9sEBVb/kS+hphbdORVW0bDdpPHQYHKx5/PF0FoWfUJ6vFaQD7MEst
K1nL4rshFsVCkvvKYy+WBvWTWW9lol82X1PgKejxMmuRMDPnI4gE4neWwP1X5Rps
iwol9wKrIMeDJJsaqyNbI+wZ+MZHHNEmaiPN0LTaMqMAGqtQRHB2GKWkye0Wh+6H
wgogg29v0srOQfyZ5K49yKBcSq1ipRM23lhP2/Od8NwvCGPDCrGiIKZS0nn3l/av
7YwEzp3M7aZvmLSG0+ahomWA2KVrg6Z3XDoKg3KE33wuNBKjhz8EcXnJfHZoNJS+
M0fneC0XD4PO88VsWwXijyqXjgLS/hpZAjxLK9xbcecIRdWZVjtwNDlTUYrziy5M
7lTSFxzNab5hhZo+9/NHESzexogmAiw/3kVoQHfS5kK53mZ2u4DMczdlCzLRSg9J
fp3phm1lGWkYZrazubPEWie8isftdjijZVwpaX3lwCwt0Cu4WCQkCVEmMrgckzOY
jcHmvC1WAwBQoBxOMQVzhI9far1Ry26SNSwTXPn+2E2nEX+HYbR3JtRtJZMAnb5V
pWsgjKqC0b4752N9r+Nl3/XtHW934eY/8b1grkHZA3+ac3jy9dRKRQ62zOaqnfRB
XmcsPnXu3EvxlFjhwFqByPceOR1aissA7zJ2n5x4q111/3aRXc3DuyMlQWe05qft
JohGknXyQoofaXrVBoeP/CTmlDWiaGQrq7D56Z3AR84NUqY2Y3yqq7OMN/HZTAqR
/DH2o5IjN/Y/CEcSBs9pr3nZmupaPUP3qVVRtrKxYpk27c86l2r15bWPGUte7GYc
9gP0ZfSlZfJ+OBs9WWP1MzTHRCw040hliLpRjZ7tTBFEbw/L+oJoW0fZUN2M6kIA
uV7mfs17WC0oUx+W3SFatXaODhiki1SqXzfWrGK0quUICtwErAyOYLlN5V4l4Rmy
/ZY8cRXN5PeaQW+pBjbraVixnOsstpDd/ljis2VF+vThn/vUFQNxhgJTAbjbF+qY
XKfObSmIoQMqWEplbJuIGjMs0T6FRx/QB8wwCT7UrRPCM0ZWY6SYEAzIapkFKs0x
DcVWpTMy/PP+732wnFcseq9F6sA9tIGD2ebLYHg38NVTTrBW+4lg5PoIoFeu+Tg6
iAru+TYj+I/tYqje2WCAyKXEC/PuQgjRDpqkf0oyGtrgB4h++YB5zuZtrRSenMA7
SRAZI4BT/g8zsaFNYNBHmd95J5A5LNmSIIqFZ+l5lg4yYz7xYLn4h0T9IoASoV9x
eXk8+1Ld4UhssI5YDZ4xa76CXutoBJhtCNU02z3VIcdcUH/dRt3Rz8Y+thwrRH5w
Ed2x3lWSt7Bykf5TdkZZKAVBeHrEoqlEqa7CSd1Z+FqPYt86l/nSh8AY+FupHejb
O/tJBh4sygZ2orGUE3AHLljeyJHjcxJh8PeOUJUDzDu3oVhhroLYE9QRJO/3lR12
NTxj2ZONYQAo3DQxN/MXdQhup+uzvHik3VPFDyX59IwsYJj1GN6Rxu5Fw3YbY33I
V/4njzRe2lQjdrFg91MWdcuEBUE1Whqo2ggrcT8/azezHuc7Z0/p+kDlsQhuPfWt
F5M8yjXT6lhaaPn1fNfpSng3JEgdT06RH+KLGyf5vN6yGL2GqKVCqo7bv/qWhoB2
E/R13zsnaof16AtASdzLFhejra3KOs78zWq7aFhiJNb8S6/TrZ8JyZOj4JLbul73
KHwVMR5QW+ISU/XEHmodoBOW6fstUaRtdNX5Gm/pvx/aod+tf0+ymarr/B7q6Rai
f6EAJHB+TbhloWLuEn6WAaYjODDyLTxCyaKSVuvt5/+Otff/G+6ay2K8aMDbdKkX
AumYdM++VeyD153npmQtSm1zkRGkOKB1nfq75InWsyg=
`protect END_PROTECTED
