`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8927x8kivier+0pCzcQCVuPYBUwW3Z4BA+71eQL8z7ZMCbnti0pnQ4LHZOw0Cf2
InDSw7MoP5EJgCmKaN+Ha9Yfa7M4wBimAt8GmjaSceZ1w1/0oOdcF0iIu2rK6fAk
g45FlJJ3sBgNWD91jwTjzI+cPL3Z2JAcJ+djbCfJMolFt5sbhQ2ngK4k4BcrUaMi
1Iu363BLEb876zYYtljHTqf7HyrtUaJ58oH7cZyoPKcAMFMsYyJwZmvmVggxZ7h/
bDWdiqKpgQGoIoCgb5zCb4Cz9sINX9Zs6SCexn/Vlg96THs+cGnEyeBCztihD9pl
8MarqFaIpDiyaWIRE+3WZ4u43vckpdYHkgK9NGnuB6uupzJZ865es+dL7Ywm4EzZ
mB6Xr2V8Qm0AsNkwDEoknuCaW7poZjFZ+YxGWGXy7ahfh8cLIc6lsKfCP1g9+sXF
n4ivl2v8D3fTw15Kjp/E4G7vdtFZ0fM7UvvD3vq5hdMNF5HzxO+ERX2zRqjo2cDK
kTAdjQr8+KXLMAP7QDK8bD480eAqfzZ1yGyU8pl2LLd+3wGry+u74Y/nKCEGNqCa
lNgMaxgYouZuiwuEoLdgnSCffT9ApiBQT2wDI0bFYS1Cvho1gX6W9URCZrMRXE86
CsfDemSRjLMBLrVhgEHhqCGFav+SskYD3UStKnh5c+uJj6cJxGHPn4ytkZLr554p
`protect END_PROTECTED
