`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lfsNsC34CqUzqZ+u2ZfdJvrit+HMf2t1rEp0VdOZPnyKrrf+cJ0fZaL+Wxp/tWGD
wDslU7boa3keDQZi16FDHHt1xKooo8IxuiHS6xh4jvWq5bJe750w6rtSDiccpM44
Q5iCi0SMDqWo8iFtqk70smE3ruHDOY5MA9lEEXgvmBHu65Eh2SY+7Tw3wa4y0cCn
8qDvMW2012Agx1tjuvD1fFEsDRRPNMtRjbAkiefSXOWOjal41HAiV7DHAVHdRCDe
JmgzNDnmSQ0yLlLqOKWEoyOz272o5+NeSZBHN4Kr46v9jwEYiIj4lDeecKcdpIaY
DKnAwj3JL7cTlJm55wyOoQIH9wrxH7+uDOfvVpmKjhHEcaS7JTOw8QVABiRFyoM/
GhHRrj6HiRw5vXf5vtBkt7MqTP2Au2hd05bU8D7cvq2bjXcehZDnEt2VXxNK1Oa7
xPcO7GizDqImZqzNTYhLhRZctDXzAOM5NGiBlYsoke6BMaCCXRqnNO583u8ej9jH
u2CMjcT6ISEHvhGoxf/1i6A7TSTS+srivXju2AkIOP5DHdefAjWnsijQuXS90dEL
mTGfjMus/Cwlb9dmjrWYLtRHv7tmJFZJZwjOmq82AGcNIQpFwfTY9536VNEKGPSK
XEMdqPiLZEbyzNZcVtuNLkYeApxPh7HrfW3Hj30jVmPNOFW5657DxpdZEatAf/4j
eSr3fY9pcFx62JhXU/iWGtr+F+RxmDGJa1Qzc2lQhLA=
`protect END_PROTECTED
