`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9aMRy6IEPioWlfMhXKp9I9sB5ih5m3dwJvYM1I5uxZ/9ZZDTv0YE6JcNPrfwJQ+1
Abjn5L8NCC73Dwzd2dJQgB7XwKUT1oli6MQa8TLTMsnTIz1Sn0llEi5Y7zNzYDJh
AWfaZVfA8p79LUahZJREbaII+mEL0YGI0X+Xwx9ZDlkBLxZio/zvmoojxAE+04jF
+0qYOOfm4Y3w+GCZa3AkcntYDyhrauqKlBNm0yE4BDhkZbCurOdkyIeoFscWoq9y
otHAs6O9ZPlezRM9wQajKHGsAt+UusbPeD3TSZsvINVmnRJoI2RrX5UHpkwOuDXO
j1UFPkkcXnsu+sRIsc2ZM0xslLm4qZ4O+r5eyudL1Zk30/wKekTngKMxwvJOFwg1
ayYUWHonBSOvuIw+hPkaIkEkJ2jLV9MQqpCcUDatma4ohOVoPBSxEOvkzuF9mLRZ
a9gxxlIrZvdjQUEKNja8PuWUkZpiCEiSn0NVhU4OObc=
`protect END_PROTECTED
