`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/8PJjyfkla94t73SSPvM0Sul/try6nrGHczMMnNVOlTa49jEc7oheN3rm3mVcFwI
SVcGed4VveDUHdlO+kiqYw3LlDy0X5l0N3Iq4EC99nOqqxXjQ42h//LP41/Y/xVx
S2YchAXJbOmCYk5xb5mxEG2wkESlO6TMIICHSvifbHumSttBQ9e2SGGCfeakNVpT
4MBtSCUiDReNKnlF5e2ML+hsQslUF8y45gx8Vt5vfnszyYJ78hK2BKdfxjkh10gn
f04o0JaRjXwafbNBbqYA1KlNq577dQsmKtUQC2nC8jd2/r7DM/7K0w5l165v3vky
2g9WhCa2YdF6pKUZ6RB5qM1w4nYODHmr2j/E0A+G2h2Oy/7UjLEPZCxN2cIDkG/l
FVw9zRCNdIrnshrbPl9rsaps8ffwbzuTTK++23tcmuN0YNBazM+O3xnGM4a3fKAF
Czft4eJq+NiJKVPDgCB/5aRI5N0+3wwUIO+IYKxyiSCU5breipF8HkbT3y/hAcmq
758Y9Fc0Gg91goYp3XlalcAt1GRjfGZ94YIdiMEGypk=
`protect END_PROTECTED
