`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpXYEyaf63atU2POdgUimq5TriZg7ltSy2akhnwQLs6he6ZLFSRC09I0nq+fz7vm
u4SiuzIYhr64va98xhy0YZSP788Tu6dePPc46ShMHN2RoW/pX7YuyUvAtxb4Oqyp
B4ytR7ReqJA+230aYrXIQ7XRYrqdsgBwOKpyZrJ1V9+fPm9ISQwmSwllYitV4YM2
WEKztbCRAcuQvWVRYOYSJ8PfKnuEvUHIq5YyoPXfj41Ho8rhA4M0HTKK1yyZkQw7
DBZI3v2jnvE9meOWCkughKkJ5wyb60MFre9JMIM3mrSZpIe6mpcvXeV9f6d0r1v3
+oDXXUeh3NcSIKvyTA51RuZgcByqp86QmBA217FK49h8Ssm4lgNN+BUQgg9WSjvu
5WDN4yLWRWRTIizcLbG4AJgHP1bhYpIbHHQC+6/O1Xphwwn3kCvpmPyRP+FUxGOP
b6EZ2R7MGZBS0XeFHA/n/lY+kYXOpGELJKnbqHkhWBs=
`protect END_PROTECTED
