`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvLC/szGocWKZFnj2IBQ3HQjTlzYxS11eIqSCOCSVDCbtGDVuirjZkFh29E9Lhtk
3U61itQcLgH9dxvgZ8++/0TOCTzk9fSKLUIN87/75QgqgxbaijquFz9VeTK/DYK6
rN72QCr4iVb6hMxawfewuNdOlUwrOuGjdZIO+J2F/VoYV8IQKiC7qMT2gGrZ0Yfc
rJ9umLiYq97HnbymN7Zpj2Kdk9t6GvD9ZB7VNauCcSZ6iMQjhBjeP0iDAYl/XpYu
LxZHq3gXr3BwvlqIMLddri/O4y8zymemL3K/N7Nt5BkH6cgh0QONQZ75w5gtkw6Z
90Wf6QwBQzIzspM3NTRxOyu1REmz1NxH81L0U/BTah2MF/lBSI3wuBce8VihbdME
Fa2y70aFYDb29SqTGQ7kcwO8cQyRPaKbRf9sEzOvXjr+7WEpTUi7C7ReZv/uT5Yz
3dhFMz4+338zUguTrYVEqFIv4MFFLOrl2M5s2DBGAyzBSdxQh5WpmuD43e/Wv11S
PSwwlsYA991uqx2C7KSyVwn4rmMDqo02YYWWGZ6++rN6EeidU5Jw/u/HMXX4mKvI
qmpD4Kv7grFXQFzWFk0UY8TiecP4VRl05qg6GSuszQbK2yRwFcyA5OSi+TQAhJRx
FOGcfLGS0MeraeMltNbsswYV+aP4uh7N2fGl6bgWdCYkFKj7oYjze/7jgF6Cb2H1
RiJUiJKjiSq59QD39gvBLfOonFmlr5GA2h9Dr4/R3tV6Fb2b0SzM+TzSBW1EdFvb
sS5avHXJPEH++M6R51sLfYj+JeXA/AIHbomWdC8QcYVx/TbYOUKm2C7C6BFFf07B
GU4kNfZ99VFGTtm8sESKjongs1KXoxyBxEtRgQYKhEQIa8oP/2evwm1lQO8UxroB
eOwaSikiTnhyNkpfl8516pJFcT1dK9sdehW3+jfoUhSaR0oD2A5k97UaD8zTMFSU
`protect END_PROTECTED
