`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UC8midxVjAtcd5h2JiZhjtWrTrUUme/nXlgP1YHaiRNCQgyvOg7RM5v9zz0L6N7z
q4GeU+Kbi9EidkBXp9LBCEf4KZlaX+x97r0JvwqQDE83jPlZn6016W1Bx9v5iwGc
u7NHGNCdlmH03Qzlzllsv1sjImm8LUcNHOYLMeMSNGX80o5Rke2LYHZQPMSYYB7o
huWXDRFmtgu8Rl2MjJyDIJJMoxW4N9fIzb+xFdUpGoKtaicJxwbWaJNa/HpbyB5k
/rbsZXtMoteMfluU/ojyqsHpr5BkUbK63ULgfBcuh6H9vNvLUjdgOhpLNDOD9/3R
YfakEjr9JvpzDNdSUdqXSuiZVmx20PjxwpyDM1A/+6Bv1MFH7Z3IutICAilFm/lf
RW3x6J3t10QIByjWrVC9VHCcoIc4PxJ6DnymCKhvkwcABu/AB770EFF1Z/lt3VJy
spNyYgeBq3HEd4/9/lnkeIJbyJd2Ank1qkfHHCvu3QYQ/aROpL5ooM/VpjGNjTjJ
1pL6R9pP35FxK5bOMesZs05ji6jPfaSSPNvefuQHyeH2+hv3ep223QEzqas17dsQ
EGPmqKR4VbzhEE8Btxgs8yhdV/frwl7l/BThzdXqwBQfwzlTy43/xSRsvvPoEpg2
+cD6Ue5Gkz7zwSIvS8P+XYq+1Zvozo4+qU0c3TFa6W0ElexweND1Hje5dGoq66sa
JTotnHe7DMzkv1LmAJ7BZ5oZU7cVJKwh6cTfDBoOFjOpnp5bfDcQtmLwURLg9kVa
VMf1q4EaRtsdUW5Rz14CD9hUzVN6EeEgm1HJayMOeMxu5j/AdGzomOVDxTrHqVP5
SRz6y3T41+glCcMc4Lb1J+/0i7RXfR9+HW2WSJMQFyyOyRUO8AkgrYCmpm6npZOE
BWbHlbAiZeTpfNhBVo9Rol71ZGXtw/nQ7Aqux+8bYQxKpFIBnzI4BEjvbcgVxVkb
NfpN/qz5127is23gbuCiyCC7hQmcB3uk0Ixtc0pVNx34FhrN88gtJ8IKeGUNHG7O
JT098tijILBzuY2vL2ITG6aaY3SpjgFxiJ+bCtkdubO4qgmh8bhemERrU3LFuYoi
QHodW+umgHUG1lq/ixICDn+J7BHCyxD7+2fLlTaSC4scGywjo9JnFF/wR7sMc8CC
y3cqJVjDIGCblm+nHiK1X9TcrgQDp+MRZD+lRYyuvOrus7V1eUBmqDvGJA+pS0Ub
`protect END_PROTECTED
