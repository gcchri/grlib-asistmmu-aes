`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BdQd1GdH4iJeCT9YBDW+5PHTWYLHrGI4K+xrf33nDP7XNF6OKBdzXKSoba7fXcBg
CF7a9d0O/EYndLJerB7XgjymCkrehpUofLwU9ntK/8T1EI0LbmvbY1wri8NsZCIH
21tjlFsgp9gqsW+e8DtIH7qVhS0gO2+Z6PlrEL9wd6QAxr+gc1NZUe7biqXlAIBA
MYQARgYrALdDaAjNGzsUHse1ACRdTE/vSaJdpZ3tTeZ4SNWULN3hvtnpb+iwmisl
Wc5wMIWRovjcSkevEfFgTlbiZQjWUy95mwWUQmh0VommPA5/TZIVh9JgqFUSd0UO
NWXVcc5X6rMGLmXu/MXiKlGljifdpnto4vNUpDyYMCqljoz5fcW019leOYqgHuAh
U/xCqGsfD77sB728YPP1eA==
`protect END_PROTECTED
