`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndLKw//EkfDxHu3N5UoN6FlEtAX8U8WYxuhVpOc+sodYwxY8DANwVGVry/ADIcIO
Pl5+EeYrSJ/hFqnFsIQkZ0m7kV0ShiG990IFhtDgIOWUKFNyYF5Ue6dyGkSdCo0c
r84xasp4+A32ffPpoBvOloFCmM5bc7SYqEBr4t+XIzCK0Hgqlv+x8X4kkKHS+ViS
KtqiIfcp+peCu/VltYH8GbbRkS+jngdd5nc6mAnMI5gigN0DDxL19t58yoY+0o6m
wC3AlTO/vAp+DnC7sq/H39I4tH9mshzyLCKAkNHbkAPYzGjjGCGxBrjpmvgNTIRw
dEoQL9FR+bIEKY9LqtlKUe/KUB4R9XfFZ+LlbYB7D2uv1A4pF4nTkTv4s0iMuWK7
7cDcSZqD/yg9CIFbC0YbrQ6jtEBH2y/Y7Fnbvh/LI1kRATybhwzNIiEYspK+VKeY
eaE5EtX0EpxajigCaXmzOUW3r2XiqsLn9E4j26d88iw=
`protect END_PROTECTED
