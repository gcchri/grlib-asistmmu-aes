`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bNTF5C9PdcuY56eP8yP2cMYzALMCu1kXIDAvgc0ON4aA8YLojTiZUASgsh1/ap6
2tXphhnxV5KOlkHvz2ye3y5MFnWq735r4Y/Gx/tDBHI8arP+6ASFB2ISoX5qJmLr
EId8im8oFL29h4PJCoWCvLGjhmDDOWCxsTneQwAfIrZaDS567k4ByNXmmvnX4vVl
tHr0HQBA72Sk1SBDSelTcyPUxJmdusz5flJHCt7XmOpA9z3VinJP4b8SDwfYrzXO
Rs39xgy3epObrLuY0pMCku8uVLDfNnRWtQNfYOEL6C+z0f9ZLYemtYEDeswnSRlw
hPIyY22m3i35tsv+gbxmsQ==
`protect END_PROTECTED
