`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGaRlTQOJ3c7mL6QqmjApD5Sa+rAtsaYGLy1IY7l2zFcD75e+49jFX74ICOqAyaz
dt78dIYN8obeZMDH1Uxr/UuJUdN0NkBPPXv7426npFZB9INT6I4p7GR6nExCMYCf
5XCzmzDast9QGJhmbeZ0hKZifbu/H/HYSeRzoYmn/T//lxnzBz2PjichwcfW91AR
8PV0skfQb7k8VsYPgtNPpl7nLShIYlIFSi+ezm7sBd2t2XjPiDpEcUTKW4HZHP+q
g/x+Tsn8qPGk1BlENETb4mpIE26XYIQQAZUxEz0cBgqTk9RppZc/3B6xsDTAwlq4
ddjOxz5fRsepLOig3xo1C1RqTDaCj72ECYx+0RxdoxsvvOb7kPMDKQGLWXdWI0fH
T/akk48VFwoMJiV1X8bbjzZfs688mp8jcG9Plrp8pLsNKnXg8hPKWqs7eeKxKgfB
2CosUFtbdCyBJjZfdZnWnjZnNug+JAHnj4o16HQNZAltbZ67MseNMIS3vS6QDcjx
EhuqcoJPN/uCglyQykw/fc+Gk1CkY4k3rfnjFhGBrdM=
`protect END_PROTECTED
