`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CcySggcfCGv4BzGMQU06KIzZk3oxz2uSSEjxq6VpqEIGQsTPiyIP6NRHANOebMP3
tmuvaiC8nhGcP9Bgb+/4uFqFuuGPzmuIszU666kqBtKBzZ5nYR5TFmZhUIMWvo3V
sgqs6o6wJUkHcH0/qjP7PR3MzGb0YRSj4lyUkJ3Q1n7MrjUoBg3HtWLiqBnWK6yg
yz6DlUJq5vvxddwZ3S4yuoM+CyLTKtR9qZpT7b17VtwAU08VTBQfvqK95YXCjGvg
qbMHCZTM3C6Av9uJXxxp592HYTUPnikb8kHvgtwYYIso5uYPisfWiE0R1BXrvCgT
fqpZiL52OVR++ozPgkzfaO6KnpvuCKM4VnvFx1ZzaVu9YziyowWiWyY9JClKAgAb
byxp0FEf1ko9bwwflblSCnOpH1lDf6SbYn/ANMhKKJ+cfdHGs05tPuYbEcEtIEkR
7FsRrpNI4IrDC5Ppj/3gtfDsxvbbsMxFj8RL9LzLo7vLp07JeNPu1lT403nDRXZP
n4rCf+7VOnkDMyaBHH4LqiC4zPXtnIw0mCHY/U8vRRARz8zUo6E5heUqczSmbXMI
sXWu3N0+EWv361D2A3sc9TFEmGNTL04ZKlyLGvWaSnkJjPkVZlOrVCFaIB4utCwz
ypxO2P0+Jw0J4HgDJPKMWvpNpTnvfPqSAGJBlQhmEk4xzZ9FpCYKiYrHu5lLS+lD
oKI0KvxKufilUiZKbdlaWXNreyhyhOZ50J2Kb2wTB3tnJdtGTwO3v2wmhCkqB+xr
FWNKz6plIimIs8V4dVvFH3StdEMUtuxsJo7w79Fd+40CqsknIx/yNVWc6Zr/BkDT
6UHSvV6P4ti306+JMPm3GAwpOJoAlvRv0xa04Gn1zoFK8MUxpLMzTWFYpG0g5Ilc
RAf504b8ps+UZyJblMo3qNaiVIf/pFRmPS+C3+IxhfrBuK0jk2qXU0hx59MHtg2D
T8t+WdY3pyNqsE8iQ18WOwTHIdRKnzi6ygRhNiBQ0dKm8+hoO9eLgBpQP/QdMORW
SojqVvjQlrolQ90a/t7uXLU9IoeGz2JfJUQLRBPXigE=
`protect END_PROTECTED
