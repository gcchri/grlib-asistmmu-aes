`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xLxA8KHrpkTjsomOD0bpKFhfeEg6tWuRR8XlZXTqSGzlykBybhU4+SRHcBu+XiEb
zmicQ0fBEPC9ai+We2n7KARFn2oBpwxMSPEIocwRkSvwDZCPeVw30U3DYxhLMQxH
04QRAbqe8uJZ2E5Zld0rh00A3jlmhqUvqJZ/pZUxxWZEU1ZYsBYZ93NDcA8j7m0M
mCi7oZbRgGX+x+BMTOHRbyzAndjMP0XSPLINRsAScWCBix1sgxpAlIrMWQRV42MA
Ady0pLchFAX5jrISfaV8NpLat6soVTiclAF5lBxiafNVFzZG+j62ymPLuFx3/s1g
1SQ31AqyvLNs8xZKReijFetCt6udy9+CtN32MgSZ8MRJ04srhBFX7qrq+SuBdHDZ
1ezvXeoYo8VrA79DTemvHRuzy4qapGi54dzWAApoPlodZRWHV5hOYrqAhnAxAk0u
egL6UqBEmECQKuef69y91a6Kakc34CkrOLFzk6ET1ej3OSUrN4dD8lm/c7QNzKS3
JVEVm05zf8iDpWKn4Xnk/RRigyyaQleY+Yqbyr5m5VXyCOjWOjaL5Nb+iqm0zPwM
w0TWgNRVTYdfPpEVjiE6MLpF/lkOFhdGQ1vJkaEN4gAvhw2aHJGOhJeJ/ZPHRKF+
iYL7U2R6M9lRa+PDtv7aEagnd5uQhy7NVVvTr8nTSyCfDF6VsrgIQca6MtSKBPJA
pETeoYLVSkDL6WGCUC/ZCio53TXpGnmd/EJCn/z4VjUwH63sSV+k70bMxf3HqOFg
/2D19j/eyFz5sESuoIr7X+SFA2PElESJUORFNH0ufYqIU9P4aOauU9bJFm9KvAvR
HgJ3VYDewx5kUDg4kFbydOdAqIweeou/XoYN2GhMaKPEzDYzLi7iuSZlbDYpBtBO
Mpjq2hwJJ+5jWTXoDfXLyupgSPb7XK87eGac1EQzRUp6k0NBpDfx18ZfQLcAgf+i
`protect END_PROTECTED
