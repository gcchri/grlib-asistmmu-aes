`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wlsxu3CcCSi9Mw2SccRVY8T5RAaGvII1C15GC/kLEzue3ZOuAMIzN7Vsz3Hf2Vg4
Afvzz3oRcHoicbK1ms6tndtDGRiaCLZSA5+GKKSFJAVq/e2LZm5o8eimYOAGarBN
F6hJ+iUOvHKLeKKpePc3PuHrlOJMTkMLhzlgT/hzc3IWLIrRXNmF7uq/0fYf1hSL
pZHnAyeJy7qc5RS578Cx+hKI39ynI73Qk3uScbPgBJc7GiRsy05vrIXgYFddwtQx
dBCxwcFOhgtMY6Wru/xgUFUauS7YPbr8q69FpVyNDDgE+EmxKHELUR3jeDISUEzM
LdJ3VArqsL4on1+zBOsHxnBznIbPY5hYfCX/YZVCy7nNjI+r+IbupP81ZuR1r479
0j4ENARDVA8ejJQbp9+HrqGY/QN5rjHMAhIg4k060Y0cUArdahvLYPlk3rT5dDtI
oYZOe62VB3D3cI9xbtl3w/DmrX71AbhgcqY601ilFmYqCnTPFN34oJSLJZRAJZBE
zIv+kQ9vSjC7KW9Ws7wZ0NBo8nmZIGh1tNtibFnCSiebXIewKec8hhkXu13F3mly
ggpbjUomBchIgSufEXDTE6F39PCcixcgjAim6j9BJhY3/rGUSht2pSXDD9FrRxPg
QJGfNNyFB4DTgdThsL8laRg7yt4aKfZeXMazfMFc5mks4wFm2ZESfZG0L0PgufV1
AohAYvXOHfITqVvtxvzcd4xdTlOx1c+QBeHMW25EfDeuDVtmxxKDzsUex7Xf6BC/
chEdjyKmqMgw9woK9OUhA/tyHi/q59Cls8C/ofk265wtsDprxQVFDOUpA0nDFD1E
uH2N3TTq7CprrwP2WoBixJVlkelz40o9vVOxOcQ6kQFDBUR/FK9W7tN+J/xbrxBe
EGsQDQJpy1Ns9NDTNWWERA==
`protect END_PROTECTED
