`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VF6KD94THnEwacKZCBqTo1+h1Tj81IT2TpB1flEQaz2JjQJFwoQgUXhpsG+AIQns
tnYt8C1+gqRYcxh9SfWlWzEQTXDFFzs8yVb8rbWdi/U2EKTOFTTu2+VY2Fg+OXPH
KWlNJZCozTot/xQYCOXiqG5xkj2eA2KolUZnCZRbfDRi9jaLIxT4edMy8DZoo63B
ikMVzK6amYh7kjS6jVxfjwEBwMFqHoijYfsQijUUx9EEDWYjOdrVzuyAWGW6nonl
srtAZCfwcJvfGisC80i3zwxlN9i1dQZ3VzmUFbQhmFsoZeXaH5GwjYpdUpdHs4uP
9ISyeMyMVWfhYJKwk6gyBtIG8i1tAiXZpMjdQcX3hYKhnRTqHgtVSRxRZPdadSNi
1ju/+nXg2HZIeM701FuN+V9KhtDlzjUjXrWy0nOkjFd/f1Z2eUBTT44lw18ttQ2H
LAXKOuIY+4aN1E2zqfnc6Erf+kcSRiesUy1dH0skAKUBmfnZA5dUs4vTzwgcP92d
34a/zB/jM9ql4svyHZnj9u0Ye3NP084mBq/1rhJLNdhYTXjB+9HyySB50r/eWaK5
dUJ7QvxJ2bePhtZismS7LFFqnHhKeXRz7oyZXPr7S7NzvBODdneYK9C9VTojYKGy
aiq7PfHwQ95NNCz91JjQipfZFokRYLwPvwn0k/9EB3bD9uHhlAhn5PgvrfAQ5rzQ
V9y7FVH/cNw9EDtlXHcL9g==
`protect END_PROTECTED
