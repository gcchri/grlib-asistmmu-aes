`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYHI60nKXRjNbC3JbebXEQj1S8tshLEV6FczaTC0pGInxJUHZa8zqxQRe9C4aNTN
LgLlvy7eTyaxUdHR+MUo3xu1vVdVl+FEzJ5AkKKNg1DhyIJYuPZx3tCtXKaffy7I
GConOD2DZNOM0jaJ3jxTErOJfWaEWxHtotfkyCxy+AI8NsdOxCPvUhuw38FgWYlF
Y7tzf9ssPagRY9PRhjoi/4/EdTCjc6Pqle7MtOS4Joa2S8W511jXufMqYg7y5PYL
EONW2BhEMapzfRFYs3tQKKMFbQMoYkfdC+pFE/GfcH6yrTaKz8G0NoxttCGLuaxx
W15lhkauIHxxfgdPI0HpEHeY5yJAxNdgSBiOFPZkch9QmhRz4oH+Wc6kRrlcnP1M
FpKbANcbGFb3DoqUay5zVWCdXpZX7iV9xIYrmMpd7nObeZecaCL+6cfcu2XslTg9
Zq0sfCUQtQdA//VJAow5da3k2XbMV2rZw40T5IBi4WEvRXPCjJ51UdDurtSpQmBo
K1MderD6ne14zcCK2SvqySeFMSJY4OEF5rmu4d2CyvD4JMzWazCqw4mly/EreQqX
DS4OUh7V+yRZV6lJPDD/7Gme/ZX+ffLlRqDpUpdfSNV1A98uJa1kksJg9xVQ1UJO
QtbDHjsa1vQUwnNsLfdBVEJmirTJjWjPaggFOnWMrw4=
`protect END_PROTECTED
