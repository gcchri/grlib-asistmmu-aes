`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TatMlL/hvlW8hBoLuMXy8KXTmXe8O8pD8GmV4q72qEcAhTwC1GDixIuAzZwRWxqP
JBJOaGHNVd5L0oDZ0CQwtv8MoUKNnzO2yAWCJ+clk0ucA2lfh91o65Tnw7VIspMi
YYgqGqyXWQ+4SAcbVBSDDCSthEtk/eJOJ4eZ5WW+8nmDm4xtGzhpOyFV5Nfzdd+f
H/f4BIDOWsi3aIc+XAUSmV6QcNOPdAkmY7tYqEypbOUtt9Hsg6JCkqYqnN1lHSpP
/riQo4SVQh4cD8qxL+jNxxDwL1Uoi7JaPwrPuakwDjmXi0i/mJsIQVypNwvzzMpP
Rbm06XL4iy7bzoOQ/PAaHn3odAD93UzJyxbYN50J4agV3OczCAvDcHlyQlpJRYpQ
S3n3A7fYpFaXQS+kT/qLm3ACNImJ4lbJgwSzE3fH/P8kWPWSl20w32eNH6+qx4Uo
fHvsES8pUZ+s8d2V6V0iR+YQ1EqJyKJcTrQzSLmQj8as9roPPIrSBtqtBvbJO+fM
S4P4ECrtEJcLAOjFgIgB9Wacf7c87egAr39Vxg8j61W/o9ay9MqSRh0U6VZkYEz2
yrV12E/LvAOZ6k3waTQZQL8AVqvqKK8nZZDoPsXmYAMOoJAw4y/pT3ttHLZvBZVu
+3+DxeMTe/gouAgmHu8Z5JfPCIKoxWQHYAu8uYCTSqP+OjRA4WwbOLji6OqjP78L
MOrUlH5EtFHyOzqcDJO4IazPzRxvSJ8GfChyQvrHZ3VATLy5digtIH0Aoxefcoa4
v5D6icld2aQnZ6b6FrTSW51J0vQOykSqzdwtKn+0W/jkUv3y+sSXpSVeEtW7/QZP
TRHNnWmasUzNoAQwv8YK5XuUpgverPXjGkH/UNcjcGq3CcPmA1zprnoA5unR1NCR
BgkVhjTyPBgdXcsrW74Q7z4QOy1q9rSsDKh1vKRxUal215kcrzLfOxUdfUfOlZ/7
wUOcitUOxsAks0SnyYJ/CRCjpNft0yWiA1hQn+lRNN4dyctf/4ovW+CdPUMtaKgg
vb3hylVDpf7MzxK0/tAo+lx/zbkgllZOW3sKRts+977nxzEnwU2DblbgHxJljeF8
m8M69oi8gB7DFyDsY60AgcZ7rLepEr0yj/DdNXin/AdR0VuWsqfiN7a/lHVibrP0
PstOLWgjcqENtIhboDamtBAuXsxBXYy2ztwU2ULJLjQpjjBMEAXfm33MrBUEkF0q
FJ9dGld57llGtoL4t8iLIjS145bxvKxYFRA+aPCJ50tgaLP0RS3T20GtwLFlUKBO
k5Qy/wVrGh7pKP7HSs/aipJWMOWWR5vTSXRnEd8QXSUD4C2CAOEScxQFGLWQu4D7
WWqN3FBqIE3b7MkdqnheecaZvJwWhrTGS69/s0GI72HYwum4i+eqBO6wR1mYspWs
zdJXxPgvfprllmpVCMcFmX86XAv+tY/OuJOClujs8WpEyKXt9kSSYJGllhTDyp9H
Bw4YCej6E+3wbtzXpeIQxCfIKiW5RYlIKt2vBD+tAXXiWYz3WUrfM5fKWl90/y2n
dxvDtycIJYLIVZoOHbL6BUJ94GMgY1arwwedVWcfjnlLZ0/0ut+30oLArYw44CVk
e089q4DyV6z1I17E5gFyCj0cPiUd4ogRfWAyF1ntCJJ6LXSaRhFA595tyOwsKwOh
HS/dRfWK2KBXzmfpuOn/sKMOQ0F67fUMAtzNuJm6amOJoB6D06NkLVFp7XYQ2nrL
YO2LXBZExJRhE9rvrMYDx7sfprYUYNc2LwQDuN8hg0PsR0iOD+aWbr25EQRnG2br
c1iE/nWOhWhcg+Q6MxNQRtI0svA5xJ2U5awJqJGzj1JDmxxomW+LtnTqyajd0LEY
+1Zaki4OEmLIrmYfHRxmUifZuGUmDPMt1nLGnOibE2Pch+3fseGZqjewE3FxXwly
v0KmM5Ly5w9y4Mvbw7u5aiBrna2VYQA5ml6gS9t+RJTuypTiCMMYGoJmNVNDe9pJ
YAjHHy6qevTju+Na2nxeNdvHyjGdZee40iSyMS1D5/VYJn6zkSXLPi8a+g0gbCgv
V4MomMRQOtMTktoqQfppGbXjXMtyyFz+Zujy++pnBQIqZ2H7CGZCa2KabLk3icJd
OgBf60e7xHDpDJACKFStHgXVhmsWtYDcfUHI6nrSO1cFO1sxioINzAhTSPlPN1SH
8OIUxdY5sV8wmmlRYD+iERwqTMWwa6C5cANT4SCPIpJNAS4erOQUA7yyNgb1I7tQ
mxnoDCj/USxrwxbh8CH/2s9STHvXfGIiI6CUoCvAumGLDoMypwxQxZ7QJbweXfcc
DazhYCwhRReVz2Yo6iJci9kGD3spS/I7hVp6O6TqlRBduu1D3gdH/c7Qi2PkWZbe
+b+upj4R/AyP9ATCLnJKSKB38QZx71KVoTJqVI15KbPX4e3E+o0qXap7miRJiYNr
ymWWRDonfXZaK1+0AUTVf1HlX5Ia/IybZgH0ewrvWOYuqXSZK6FAdC0YUdmyHefr
InolWc+oWHymOCzbPg0LHOHAhVcOxP04OIzNqi3+70wrZ03Y6Fiv287/w0AAd9tH
L+ydnY66ubuHZMQLHOL5GyCwspXI6oTTUPOiI/7pHJ46ODX9FFp0FXsR2aekI3ue
BXbsH6NvRF40P6BAFfjb/b+qoEuJsAOBaES3xicXGGRtJT26GOT0GfXStNv8Gk2F
mcjn5xmiJ6am0FpAQMGJww8JtKwyZnV/Yq6PWg735czWJFj1R0w9YN20S5SQzzdw
CC+2pPTvatkDOWPAFlM4V1btKDK229tPjuVX67snNvXWHWfktGDslf/F5t1ur6jG
0DVsP+FB+tLtHEs4fjfLoAHNcqNEZtMT4N9reZFFn0Q40j6x7xki722nr+jgWxQ2
OlwxLHMbnYhg+PMaGQ4RxlNkiGqQsjJkozDGoLf0gxtIVSZ+3zOlfqicUrmdU/X1
mQwflTsr6QhYihF+j+G622JRKZNmiXz6Id4pDouWGfo0yt4gmXaFshZnkAX+4KeE
YsMmwpuoU+zbEYyOwtIoU7dO3GECWa5dT4QauMV4IoO9Dup2tWWLsOgAA+L0eGLa
ffCJ3Wh53j5p86JWB50Ms2iB+xgGdUVQp082lSyUzZofoi/9sNbeAUMomOKdb6+u
hEuDeb6ofvKQ/23hXcqc1DxUiWqkDI5RvJM8u0d9+bttOxAeQ0WpEb7CqN1oSWcG
lSwtA/6FoAqpY8N+BUrtN7sKl5Sux+Mzdco7a8wKeCR9nw6nWP5HRSCLj2iG7GnY
rCoNhOGYmjYjNDBnONR1evzDRfrvoSnb32l4Bo1RhXtOi9HMpw72yodnwhBAfBjR
rEnm76bxYiaH+7TTmHlhLb/jmhn5I41f+wQ8bLdokHN2fI0KFI4LRPB99oM3KYVl
aCJeOwIYxxJjIb17iZrsT7ifGJjrdR4CCOgCa0O/iz27uJKCreSiPKeosHSAOtCV
I/9cwvr77hNK++N0ibrzGDrN1MdcyH3giGkeXZbRcJSQ9X1PbyRXH0zqgNKZDGgE
iSKkNzI8sqwPKF0abF0RBosc0QGfhFWkgMUbgatk3nQKRov+ZTI+M/qxn/jfvQpk
ziV/7mi4WRpfQzoQrPi854ILUfTmGVkpAEMg1zzlDatOsZoJ22G5oc9QDaM9AM3H
qMQjtfialrOfEIVzTDyXrOx0e2dcctPSTWjdDjqnUy9DeZ5W/tEy3Q6uiMfhBUVs
4XJfgbcgrhYKGf5tVeU78zO19DYnmbIAI6WwiEX5NJtS51/7czLOuBKdpqOzjR23
7yG3hdDuwUCO0ReEkjfuE7NJo/4beWO/4H8cAxQpW9PVkVtNshmE5HRuaoTpvMWV
4eAwO7ZTOwIoinkjat0dHoj9VsVaOYuuDjOUzd+8J37eFP9Bj4Nb9eQ1JkfUkIZ5
c/igqgjRUwl1HGHYDpR6tqlUiMaC9lRw0zkG5DwcnuDubG+/pojY5VsxGiVFZEwW
ufI4KcQByP3MuE/0Nz69ANR1+D+xXTnP7t9CbpzhDmY2m8gxdSU+nCiFb1qTA0aX
4nie0f0/90bzsVeeIVHKidehAw6TRJozqvYG60qjckL9FGUlhI9SSsP6T9NRpEGV
HkmJC+wqkr+1YoA4RrecydgLu40sDdmDrA4077boE8KSKxcZbHnobT+10xHQJkGK
FehKdiSwtLE0hr2QAoAMgswlmlIENZlB365LVObCsi50cLFpYyE9Z5Ry048xg4oH
h3DunIqj96YUvSHP7aJDcNafJ2PD0kOBsd2Pg3YP1Ngx1gvrsiaL3g52ZiKp8G3L
Diea7bEosUsZZcQ7V3quFX4Y/4Vb0eQPPcopplw7bgTIfkXZ16j1GwoG5uCPc/vI
XiIAwqxRuEXCzk31F3hVrD/7E4Vg0sq+S7Vf2kVsekIr2TfJPaOP+edVRnCHEdqk
8egQSoXii1XpJni2eHyFUooRSavhYdYRQOfNljj9ziA28WU9SEs09rTH+H7KvDGH
Ctv4G3yqKBSZNsNvrO/1tkA7VKjRMLJ8iooUiiY6sQrIP0SfLPS0kwe3sWDtTq1f
KpJDcDsZFgA2qz8OwMze8Q7TxP2lB0QQsvUtJqy3GyzkvLdPH1tuwE5v//KUzs+w
LPFJL/zBTQNNfNFQA2VxvcQTA+e9mCFl2yhTEOS2L/VvjTxQtuvWhlfdCW1s8o5z
ZiQ5way/Km7zk5ncdyM014XiMsRx1/IT0JnwDO75K2rUNkJXLPZ+Q2jrATQrMw0r
k4DhESnSOMjpo1gxaJRYeyPr0wzO2xRfp+h0qJyplmJ929scxOhWyvLJdoRm4ZKE
Lnr2cRI7kUXj/1UooGkm9rQXmrUu+DszlaLmOAEafgW83hV5b4/JeRGOC6WvvbuH
ojae4h5WotYe4jIYGdNbC9EKoWy8chqWy54nPl17T48Uh9qt4VxtqKC2RQXLAYyd
ptNqyb0C8ok0JizntL0x6f/P+BgBACkZH6IzJdEiMHzfBWAg0EKj/ZHnFHfNy6LC
M3+O2MZjmurRKajgCoIiCQhyXjpuMENI3qZ9RqPt+PwLS1drDHtgZGkcmWtZuIoB
OcmJbngm9Mk7tBZgQAkE5A1i7ys5iSDBixquvmMUCeWx9i75MYhCH9N0C0nBvQVl
Ipkgdn+7ZD/wLPw3W4Bq/WlOSqVv+xWHB8dhxw3695tnYhoJqONuvaUPE9mVz5fo
fqbCYV0cGhf1+fWFiXyE1qILTcc05hqeWpd3cni4+Ljy0fVHIiv0qABOsTFwCV2P
IUyUqsygSuiX6e+C7g/YqDi5Lf75icSwLBVi3fMugZwwhf/gI18VmkwDsVk0DIu1
javR3GGydTusUbK91cU5Vz3eNECvv9Dg0Zmrc5oWBUqmpNBsDk0xcAyhNPCXwdxf
UULBj7DuPDDXCPjHNabr8a5TKEe9BH2lmuK1nBNScbC7V794k983H8WA2GjBPiAU
a/XnrEwVSh0OSFEXPesnPRLjU+JG37CLNVAgJVCzZwlSNSL/H2G5lpEcede0RkMv
J/1BkZORMnywIgOx22Q1vWbMgd9SXitX3pSYLjix0/R12H4sC/zUfmUaSEPnNzUR
lkhtMKBGDhFYKpgd2ePPkW7GVW04qUUQE+1iYtIWf5z2e74XnecV1Og4i/nUoRCZ
LCEmjImacXZhfPM63rj8evjsAozeduI1fI3e4pbmlckjUejxZqNfJcGrCigDCSqo
70toEWICOjE/Tt08k+1zEvQCjmMt0yPmt9jNVFP5nfOmkIeb5ZiIdyAUWSufabmN
cFk2lbiry09lkMwHOWoziGjV9adEAZJxroXueKwrgpzL12lwTOw6dU1rr9j2K+wE
7cxNJrpIMaA+hCjU6XpxwyReENs77W6jCPyY7e8/IZA+vK2YoYrv8aFKBNGP/3CD
HtZQHXBvdlC9g/e8jydUkIrh962CD4qEACtsFlNdhbox47vsRj8E9Cz2UNEcbnY3
9LMhk/zs1D3dHqFJ6eJtV8ReodVFY3KIywSmidIq2uhgB9oB1a+TLnuG5qHl6gra
0wt+eR6hiPMQvVTMDBRuWIVkgrIZ8LOaGTwIVF6uWWJOIswHXpZ9kJyBbt1uRJ/g
axEMcJx+shscgmxXIpO3ttcdEJGxK5syOn2eFXTYBcbGVAd7tbWCC7ukCCAx+5aR
QoRwTmTwu2lf/d2FzmPYqXFzfDzYvRdf+OavWuLUIH66spoqGRvw7kiaxYo18Z+P
jnZGEPfGih6+74Ado3n9Bs/cb+iJPoGaB9ZXUNx9EQYR0iBxVGCgINtBYxGGYESw
g8EEdZJoWKjgtOEE7VJayk/HZ2FdJek51ptNnC2Hf/BiBK6IYITZx9q5WqCCkO1R
1gezYF1RNNbOlk+9d5SrkoBGrA+x1/Zh0bV8hiYE19pVUMGXnbxGgdDOX2q3h1+6
tS/6mK3uav//iOd1wtZyHTU1fsn+YfGeybZ6lEUvidv9vHTl9gtL9t4we42VXBWt
e3u2wW0PwM78io5oztVdyDLNv+O23VgdYxYiv1h5TVPfC9BoGIX7vUFlrUR+lf9v
dTQxW9tBC2RemF3UFtYILeFiyu7ckERCZfo46ZOSuDOKQ+8Cvajpzh+QgLk1q4QO
8oI8CBPDFE+ijFbhYwj7L3Gcpg1/W+zEXcTWnJF8myFX99xea3yAkQKl1Ll6vdqC
d+dEd0kBol02d2QbITbhs0PIH4U2hCwJ/1UO8686YwFWFo6SYnHR5tZ2vv4j4ZQQ
LMalsqmCXFJsLo37LHfgZcBrVuUh3VLju9b5NB8WuAiZKu/SM9WCbAGwAxdrnoiG
8fX39s3vYpR1bmq8reNVUwCescvMvxegGzOrHI/tWaSnH7+UXqrsVJ1AyQ6HiLTr
BUZ8bJwwWUTDIr95jivcCneZ+mrOcdsCWWIjiOaysoftl0c/tWMvU39jGrvuYHOh
d5JrjmOvpt4Y+81OqXNlnhs21mifLkAXEzC0qOOoE7e6u5CyTGVU/jzN5Rnrf+uN
njkJ9s/mAD6WarH/22bqrcd/GzWZZlqzzJjBwTnuMBbE90QiatLzW3H70+0t2tJN
EWH+U4VY152LJcLyCXbsqo/GXlz4KO3XSMtwEaGcx6MVzDN+ESnvF3ITsnCm8oPO
qyhG+xb9NwxCEnxL9OEqjEQlqGc0r6LwihzF3/r9BvldFlaF/fTysgijHGVy2B/3
X8/BGHjlYOqE5Uy+CoDmwR42DswRAb9g/AxbdNTe8eHPDyLcerSEB+LQaFvBITZ8
F8jMLcHFxH4ZaIeOz7qVC+wESPG5iUQW/epHsJU1c009zs574Xs2D7BRVJcDIQxe
wK4w1Ag/Hiu0vW55LjR2oGbJE2CJU7Tjh0UufCsIKlj6rV5vpKQn9K82Vs5a/BGe
pGwwfMnw5OdJQ5n5x5NHOGUqL6ISsZ+H/EJq4PPKUBBAY+OpAmYPtse4CY7ldMcn
OkuJ9fMRpoVlEUjp8rAVRARyb/u58MrnE4YGeRLF3bcnQivINpxKu/1W+fweY4Sj
fNd5WOUqb+Sac5+izlIH3/ZKI71L5d2iUeRLblrY6iMeAHT1ikrN+GqqN4b1IpXP
4GgIfRBiBTYPrEFL/5Qh3jMgfNHd5KsYBbgu7RnWaHhxeQ64ruGBPuAWCInZAGd5
O5WXtLWZhR6keaoLOYDcAzXrtmceD3RMlE4deKJzuUYUz+XBT3UebiQV6kFl80tJ
WfA3juLy4cdxhUbxfjMskm03Sp0lUUaiYmSv1OH6SU4h80ZWBfigBMmVCnPkOEkw
W2nepYMLqKkGnNZYZD1VzduX4BWfuzoqF7bJKJt7o+us64IU4NuvazVgVC1tU6x3
eMMdYX93h4Lq6q3tPJuXK8RB05MiGBsKvWnX1Fyz1eW2GnZNLk04ulz9ugsUoO96
ic2EN2LHpDw32HbLchO+8RbZyMNSKTEM0NXq+5hm99D+jHFn/JYiL/dL7YopeOiP
PBHkRNDNpMxe9sPo0+wkOZTcSH9pdRT4zyQXzB1QxdscnUuvxQ9ss3IzjDS2/1tC
AGSBo5yyyNOoP6SXpj1M68FE72Rx2uaGeEhc6ptgUAguGeOuyfVlJ/YwGkdNTI6n
8s3mF+tz6MSu8/WzmIeeVzud5FLJmgXYxPbPMTTGUXUce1os5dySw79YX3yBTHBh
00keJeghvW33vfPGVPRGqU8RSvBEfRSd7F5cGhBeRH5rESrARMJBChXbmnPJepWE
P6qsQ+XfVCkBlfis1G0QTMOS6H0EH3ovWMR/BT8rcMzpymCoWHK4tDFPtelTKhXo
0Tu2uZGi5svAfZgMlPLESsGM7xzz6PFBIQnso/z0/JxriaQyAH19RRPuI0M7XTfJ
9VYHcSAw9nvATORsuq74p+trNTxGFvy7MfMVW6HpLR0lsdk0/gIBuNnHkl1LRsR2
TAuhobExq3rF6tacqqlIXmotgB7JBvYPdDzfACEccRk18+XMsMvYFs0rqjLt1Tb4
JJOCUOSiEjYEBp9z4YWDMbIwpZsC5fbXvDgacSFsvUOMwwKEY9fBjbcXaq5vJzQU
xuQvia87/pjw09mCCUKmFSawMxfoHoAgeUa+xf9Nwh2mXgbhhzeFz0bRBGx8iIlL
gBCEQNyLdNXldRjqz4YZ8hiUBd3KxMvEqkAsuEvWAB197n7qcSolt3JIanb7duSh
20UqBdq6WfKADsa4jZde73afEwZd9lCt2utfQ9fsVy7g1VxyXGBSbxef63y3luhh
s9b/Z81M8vhFyouASDJ51guD2TWIX11W5eNEFSCd8dDTGtZiXuSleoNAtUnU0LQ5
vz5B/xV5QJyamD5hcpCuPYtpulG2VYv3kUEUL/j5IM72pwcu+4HfWG78Rij5iKw5
Apo9yPHLBiColB9ZnAIrr8lK5tu61Z+TxbftJ+ciSaomgwf6gFp2pbkNMBpe7DxL
pfJJ3Aq3n/iQ87W11Y1tV+LLvdYaOeGXOOPSCZDtsH2dKYo/H0f2dxohwPw3/VA4
TD3fdcTa5SwVPQ2Qcco4/VLDdWhjtXcSFKWx5V9QW/Mlw6PZ9aSc/mXkqFvshwqv
WNsKNTKaWjMccfhRcTCMwisTtvIeZXfabfM1J3I5kxJVu7cSmg+Twf6xHQ38cpxv
lg/oZHzXvqsS+w7wlkt/esOitQXrSXFvkPrfouE1VrjmW4I5HOHdInuVKG5VB9aC
9nQWeKa4U5rCGEzu6J9e2FVmWVJQfoeKFhVMa09zUlhmELsRa4xNPa86DH8NmnDW
sS1cGAgGNlr61gffsbBfuKZvOA0uU0B4Ddb7jAVxbWMBThiFhjFGmE1d3jdYVwSw
U4/bDWkcTRK7fM3uxo8VzfV086fJttDev7YCwMnJJd0rO8AyU2qcfpSGUafoKtas
tMRQRDsQXSqWpsYWi+wWAzgLzZ7jyH1pt2yci4GHBD5CeCj7bv4qLaGicsim23YO
0663z2hN7p9Z3yAatrP2UUeaaHwtIRQUjhxJh2ZoY9BCrTFadfPmbtuHKlSJQXAw
YGNkOIqPBHQUN/Qqp1TXXh8Nb6oT71ZUARiFllbUF0VF3Ut6JounObbuaLpYd0rF
DsnE6ziXxReCh1Ez62WhiIE03aMuRCR7k32QWj8K+lhZW01pa0u6b97YbYAv8qYp
CV4AxUl9qagavbpqgTBlAmZ/hE6Tkb+ZqNu1bYeNWwXLxvIMZ6hNg2rXDX3sh80C
EzpDYEmZ6d8bPbTbHGuWasnLU93yWap4j/Q+TB1ChGDsii6u/0/Py9ZDnPPu19Z4
Cd3MWE8KCmV2/Usjn6ax67kCGoOWc0TUQBFEXBX9H6eENg/hn/Wf7AXTe3cGpdaK
ougdejQN+6xFtIgubYLUIsPVqtAdu2yDePJSfhgyY2BTyy9bFVrJoZTmFQ2kNHDC
FO82crSjT90z8Pb7j6QmEvNThWtfYqCI+XGcYI48kCNcm9/UNuZYcjgtaEWU/azc
10FGEKQTKrMGhtn4gaAkEasAZZi/XbYPGKqHeIO7qv7jIk5DdVWWcWU23avT+Wkn
nA8sb5PsDYaKiFPcwvE1l8Z90PpcZ3AZDjDaf523nM0aqQbyxt4LktFMWX/Rt04B
VAk2oF+piJ4IdauzLjKu3LVJ0pCVuIM4CWALo0ZdZMs1uNAzMvHLm32N5/1tNzD5
sq91oNBnFore5XKqffaSwazX3a6wem7iTujnpQzCWS0VwHWiseBTCteMCS+Zz8RR
YDNCoRk/z7r2xP3snpASO7b8a0skb2BVxApmoRs6dvuwIqrQf6b8ex4cUVUh/20y
VxdQObrHQf42JcBHdIflXgOXYdeU/tgoucDA7uefbnzXl/q3YGU4QRfrlgnfTpqN
iJJrPoFQwUhnh+69xEHpOODHAGadI2oZg3LFxbCX9tLQ4sGd8/FTUflCX0Gf47Qn
EZLynzSG4SICvL4ACgyhJvJRShu17CRVA9Rp3RWi8nKabQziiA0q6dogFjttPAhV
Zic+7bCfqbUbZjpgZ4uUn20u/zAkMKcKWVOvGdN42YxIC5DGS+NEN9qumEMq0RSE
58pVZZTTvtfJ26hoIS76UURJ86qtzMA82kzVysbnGdH2LBZ0z4t8BCBTD+mGCFik
zTAuYSn389qA24PHfdKTS1rYhhkgasB/YGHTvMds85u0pQE8UEkVew9796oyb0JS
p58FOmajZS+Vn/fn6cTolyJ5Xeiw0kqDGPkCL/xThqhw7WMK5MZ3SUmRnoEeAJqT
dTT6HI2HprquU9g3/4NFlLFNfFlgyDYRTwFnhsC05opaPH6IObmdpt7zgj8HflmC
U/8OrrNkLhFqIpn69d7LjjOxD3pOkGA3pfLjXaMcm2jfdj6UL9ddbxEeJa+iTGwM
NqHCQrz4QR62t7xZhFefYUuanI9YegIhwZpahHnD39MIU6PSy52g4UIOvn/xvddZ
eICjDVUL2A5khdgSk43hfAX7SaUF7PAmBkc+8unrMkVnzsK2YpOgHsY59IDQcexk
IMusrFlCS4lsK/cZjC5WzklhhujA2zhcPI2SjlT1MbS7dy2IGGRHCByc+/tQdlJL
hAMlCqvaX/oU2JAXOiERQg5t/Rylac13Kwyzrjyd/g/JigEnwOOzIQwWP2GVq+mS
9xlosDp+VYr2WgM9VNxjYnOW1P6GrvLzr+0U2EMGD0LBb+p2wGuQgo1dbqUKKDki
b9Kg7SYeUAdMmlxeoNZGe4NTq2eD0aD1lM4OMh8TjZM1ztsC8+g6zNSaWrjSKcwq
jkWbkTZoBf0aSmOeVcRubI2UmzuuHH0ZHPkXFPVFAW4/RZadKqTP/vk8ghqFiPy6
pUdXxu69NNaOMnIY0tJK7n8dMhrRxNtxh67MVzzFD+LQ9geg1iP81jtj+TMFkQPZ
CPPTb5ifSVe/zmhJxIamET6s4rDXezcGALBaN978zqiX7osPdKGiRTMMyx6DcHaX
lZZ/64dj8hWx+phklI7fwnRTDv+1E7/6v0y4MLK0Q8BZHdHpdvQd0cisTIozwbuR
8TW5Ho9Jz2bkoSqI5JrQETBMUVLZZrnFRBt53Bvxa14pwutkXb0K7tIZdgYwHiRi
U+r0Y97kAAUimo/L2ZBKzUjxHYBnMsafN3LZ5cZgMkrD6NOHIqDS1M4QFsU9roDc
/9ivG51jA2SOrWaOZQs1Z4Zqp7V+Vyr4FT2bMGLW9C9o56zmIL3WDOHms0skouW+
1O/6/Ncsze2YMAxqRG7GVdFl2TKs6a1k2mIrbIFJw/+eLGSS+WObHzJGhD4ooCsp
ns4qxst0UV6nO7XXOPK9FJTHCPmE1WgF62uc8VD3oB1ZV6/mND3RhwnKNhsHlHFp
AYsKIkb00prV5BD2xt/pc9WQCF7MoMKoe63LIYhevPkTPA9eWJ43wUZ1zOjAa9IS
8y0RjyP4aMKGWVjYdNp6ZS8p5bOSzJiQbYNd85eQPIuDvFtz/dXsEVbp8rXAbPMn
Wv6DwhlMd9qW61w+CHZnH34bVy8VdX3Eb5dfBWGdhg8pY1jauk7j3/cnOUmvR0mI
47dJrg/+4leY5QHz6xPTsB2M/UPqDWM2BPaDEIEFg6k0f2LC7auqTrnu93A1DkWp
1Ykls6cEEXtigv8gV+3OIslQxrVuEUXftHtDG+HlsAuEa4U3ZCQe+K1qVK9juQHm
l2O28icJHTo4j/eW7CR4TNWUo9M0RnxIqiFgoA9W6dHG4yjkZ0bDKBAk9/p2AxD/
32fFElFw3kgEtWrLt8rVYrg++ZCliEAtXU06jOr0IRuNHQx8r7AH8KRmFUYvbMt9
49YlmdRdIKZd8HYeCm4Y8IE3wPBmmHAuRnvCgW13AoNg7LFQAMP4cx6WtNyHwEAW
McLCmP8gya8WBCAWMnZGmzPl/BpI4HTVDpSIwoNk2xqlS+sfppEGSabYOzzqIpLc
vLJRL2oRdrmvZyuY8Z11MY4JchxuQ6W9qzoF4lhQfcywq5jFWQjoh3WstIYIJQUt
d/DKsCpAvObPyynkQUhfxErtaUcjaWZfhmPAdkhoMj5tmx5wE0aErbEBDTSkAj6g
p4Lkpa9MSEK1ujVMPdEec2zJ7E8B960dm0fmooAY/dwdj6juuZTiuoetWt0BLvKs
IsBo8641mZunZZqLnUtcpuC6C8DWsu9FJecXaGJyemPcKm4Il4CchJ+2dquDhO2k
Hu9PoB6a6vatl/ugxBm7EMH7KkRQqgri4C2bG4QHWxAj5toKvup+wxkP5GRg2shX
H2a5duNkm3KM4X+Yl0fn96DfnH5+jPjF7BWge85rMGwntO6zDTWgUnPJsD5FCjMa
1ZjTNzyn7I4mvexkVdea5X5LMdo0KIgu+7woBYwW0/pMom1o859fEfUGeBhNdPJV
GPp5uCLT1WVK4OZwPxxeYx8agH7ttzrIN1Ys9npkmvd0JVviS0/jndAHVop1m6Jj
SVXJ6cCixsRAPUjsHn3mReK01TT5vUSSnB6/Vvlb5i9TxQ8hG65wZKOqXuy0tvWE
VHLoTUNpgnpXpN6cl8eXSVXntnwhVAZeEpLAWmDZ2v0oRiEZRq7j6nbeYlROBLfI
rofo7/xwLNCWG9lkFx86wbVJwwlxJ94LHmgCObm785SfmE5oEdFZdt3PIH/fAEPj
fENAOFKJinQG9ARJjwZYcgrvD8E3H31XTXjrFDyQBDeF76oOZY+x+KSJe8C758TU
0eaemDzr3liK1WrzMsJWK2KAyzVWw62uY2VPY2ilUCbTd5GAmJ2trk4oz1x0KiB4
YZa2jNXvR+hdYxCxjlHmIQOYY8uoIfLaeeUOYj7gq7n3zFuLZhWDH6Xihx51gpxi
yl5HJAI6xSM7kajuyhPJxKIJy1k7pSv5PjAWaXfKbV+4N4/UJZeCFBYJ/dhTyBzp
65Yf7z3c9X32+Kh8FEE7aEr1+jM1TiNjcu/Qe6whUJjCUw6HzoF6PHjS9+bRUcsU
XYpG7CeK3B0G6asXsx5pKxG6CxhCLIRiBuGsYIqPQz5c8ZGQzTGvZUdVwTfnYtKd
6riaPDdB91Z6l4RZsfp2p7it0xAQK3DS98fwHh488d4xJmu02/5oR9wTeAQDeEwo
V/fyGqqDvJnmw+pmlfs0m25NhBYNlimIyuFPeacSMfNb6Hjg9e7P3Tr15+2focos
eUjSjeIowLOkmU2yorALDa/+GMzcnk8Hcku7K/3n/99UxizR4AEvxn7uxctPWrz+
tH59RVQKp2C5qzCHZ7IBNCNeAgzIAaIT+Klyz7fRCDz+hnoedn9HRu6aZ50dKage
cB5tDKnDPn99+1BChQbjp8oHUdzOwm2HTjtsHhamMuPW/tZTosTy1UvefM5hTtIF
GRNRAqPzOe0kAv2fZ2G3q+7v929bp/4DkduTxAiPyWpfG6IYZqu6Wibk+f2yBSjo
DWiBRZYv7E2zYZIp29oQN3j6og3+xjlWX9XKTZUCTl7ZrUxVK5PUmw3uCJikF+wb
mXAoI66Fv+DBSr3ntrX08jghzIrwDqBpehgj5kCeyxN1QsLkhLSJ0KSvDcQ+fCtS
G1Knn0WDodfs/mTi1emsc3UuPA8FU4hbR21byJD9GYCWLA2m4/oM3IF46C3j5RbH
rM37EjWoxEajQ09l7GUpF3bOgrTcTA/VZDbvA0C2CzhnDd4cMbs5VozpBXrkbnWg
z4HjBfGyAFCtV2h3l12NQPzZ7tQrn8f6GMW2TE+zQt54tN4D1wOQEaSdSiBnycJw
pSgj1//tDVoLEvMaXSA+yqCbGAfhVb1fN8HK9Rxg9d1EfVT+vco0E0sKCC9SSe8B
sRjZYjVE0DBI4AhRhw7vTsjo5EsuAE//1JiqBuL442IwCXzi2dSXSixebuMSAGRQ
yTrJtrp/FI08/adO4Z9u8yNEFvs9uE1hjRRnbVlTCqOP2nARhSmKRnW/pDqG2llg
8Q0ypRIUj0QKsCnXOqWcy0y2dLf51gAwrlgrZqGn0jVkE3cFBReXWrZ03q1kwLiS
ZtQLclR22rjv9/whIp3pcWkjx/ik3x+G49viAKwqDWphEi6VUW5RhwQxXqmWdMIf
gSlrUObt9UsG1k/YRUskeOfJqUOJRDqBkUkv+EVjAn/J97avfg1jCMwW+ZKlDu5v
YD+Ag6AF7VPPnRDSDyza0EnrjmANRsDlWBOo+1QSVGLqiZ8E4xDXbPEcqCz+P1nM
Y8SVtR/CbKJpo6ox0fuvctsXW8eEut1GoS7SGShyluKCEJEqMPRASFXpgxg8KNeX
+U3WriO5CZzFMVc+YTVX/c+fTdQXrWUL/X9XedJmfX1adZK29H2laAzofRYRRbld
SstnonZ3LCMZhvCKtSjX6v9GArJlP0HuvHM0kNbFEMaTgujlO9H9LHK13ch53SW5
WG2fViRm39ol/hpDs4PoZ/7c8qPGoqpHwMidtdq10VbkEQXbXA1VHFBT2nAa4bbX
2ZbGI7TAsWoHXOfCvnSKNonj7ejjxhzXCPzDoTbDHnyjU55cryMPyHwlgY0KCWMV
F+YJmLAojs245IvHDqKFaXoNMITvtZ1s45TfA6S+WHF4z64iaBJdP6xoDdoEn9eZ
2FfLlmcZm8eAKPj6Xc0vw9nIR7aYjnt2ME2Uekpj0MkK3x21Y1gcH6iSUKyYK988
FGYDo0kPnkV40lUwKx43NciYA3ER489cUdUmDISUfrlpWnQYxDXMHqVfnaCpXnG1
78TCUTRwKWufiP+PkBDG2tja9J6oiNDXwvdTFIrgcQxvFMW5pdydImqTGNEf9XdY
9Tk+HXxDw54+tqOYpOWJjNmGt3Ahr95WsGw0au7ZuzRmkKSu4BZecjenXC7j1/8q
RDcQeDMkZRg2X3liDggfcVWOQjABv0yheNDxyS+VtH/42GRoHErQhzKmfGl2taNS
a9K2pQsX27ENx0h38BG61dn7Vq3Vibau7d4hU65EFra00Gom/1aqLdB9GmGF1rxR
rs2GGaX33WM9rTGiHjJnbJjGf4oagzRP7cDys7PNn9VZFK6bGfyN6Qt+XjAZ96Dg
O5dPp+ppj9Slt7xOoD4C/TZotQBu42mH6wo6HWYqu3/Na7ZSLq4gOp4waeEpgQ//
BK7C2TqatNcnVn+3I6rWtwgRG1Mn2I5U85GZhGsH+t2eNeoQZm0PIhCP8nNwaLrA
5WWfex+6z7yjp5qU6Iy0BoDIfkzfnHDVNtHqAIJo90iZ5bQBTw/uNzPwHi+zEOGt
NV13LrhjQQTO1D+Q16mGhe/Kd1wLftcof3PSPpP/sjNTAeEC0kY039ZIxgD1uk++
19sszFELdaWiu5698dkYjhZI2BWoZsMeHVyhfamWhE5B7hbA0hrMQL4/ODjgdkNd
GlM/2QzTv3pJyMs9d+/G20yLOTMuQKVgUZECTHd/6ueNuT7CD/0n0HCCzsyKDSem
BfqemCFwh/x5i5tj8qrLaeXSs/YztHXIA9lfhHTiBDvWlL0LRwA1ifUp0/immbA4
ZirKDqJ0y5TrdEEs1MEHVGKykI+dfIDFuk5WJIJr6VcqbZjnZGPt5j94VZSERLzF
IgN11a2xAvvLzSfytoPk7MIdgAGtTHuoQyOHYmlD312pkIL5LCSknK67ki5s0h2x
OBJfowqhNsqK3mpBj+cvU1XTgkz1LzGiM9LWKMhrUSl2YLFWKMEdUss2wGlByRty
txMCPborprwaVixB1Sq7FoJU2LBgQ4O03wzVQIusfLbcK/NintLFFMJnoEAQ6of4
MH0HUcV9atvNv2rUtrvmSTn7M5l5nnHhZtjVupGS73pRJn6cu72J5oJN3j2fLBut
a9FYl6YryLD9C1dkWg9Wo635pxmM14H/lgIanwTDMkzRwuPMTMnKY43e0fcP+7bu
Hs+QhG/WjvInOrKm6XZa5j8h/bZ8oZwkw73rWhJIDX30zIGw9ouco7IFN57H6R31
plOYryVWRh1hGWnX4P5CQJ3WouWXs4UVZ/4wez9xTVPKZwNcOnVqgwb8+96CVHnJ
uJ+DDLTdxPYG5I+0dBsRA56jahQNDRWWv0nRIW3rjwC/jRw3M/poq9oUze9ikZVw
U5ougHdI2Nei9wNPmDjWmrU9XAVBl4rmLQQSKk0uMEAXQ1/ga2BM4a51MllLT9hs
uvOkcqVMpBG6QpL4Ir9tLEXpuHO04pIueLvWFpfRX+6rSnry+RNynrR18/hYruJW
n4Vga0lBJ57gGzyAJ7ulaPdcV4nUElpCm6sAhqs5oCUR9GFpF2YpKN26BfvIq5tR
iDOHAWSesLV9qRHsZ+oO1SNt01iMy5NL5UjgPSpCLL3tVMnYHoi4diVvoagOeNcG
kZLCqzT+0EEiS1oMhLRCpoGEg/t5bRoZ4OUCQpoRBqe05DSqZmIlwdREWMIagmFe
nruwKGm2SnWRe8qGmlHYaGTUP3Nv+Qw7LkI60Tp7ubqcrIXK0DHBIs0MWjsAizC4
Sp8kAeXEwUtLq4QCKQYqZP09xFbXccheRv9z0Dkwun2afKOUNrKAZ/i4s9zVckoo
9R6bWc9C6WGGijym09UrruoGaWu4MQmXOvsMFL6Q5jp66IMXagrDlruNyGtRd3rM
ZcIvfcD0NJF7o9lLGu8Q1YE6mxF0IcPCHGmI2//tTsQEAUMlZE7DJVzOv5t/B2sC
0G4amw9ExvJFhWb1P4zNfM1UoB6+iPF2Inj+f2IjwvX4+5In4KhzL3DiHysPyEvz
qDjISEZyDkYKpU3aaMZRVJ16OTqoICzjpN0f14lfSUZjl/ttgMUAT9dQb6uwGhjt
ctFj1L2JwZAUvIyvZ/0wbHM+0T63dqDrtk/5MQCOg35C4+I8VomGvMcrz8UzsZHQ
5YTUVXECqSf+y8dLOEPY8dVFkFqLemHHGDUtYKU8qM3yRqAPrWadYnZTBve32lZf
5lJ7HZxfd9h0yQdsIFvcjNjkEDmDmB4MXTwABFE/EKRJTTHOoMug6J8Ip5M5mwpT
i31naZ3TLGzp9i+g1yWtJ8uu+1zQSs9cPc0MvArHH4qeRyrmoGLlt+kV7hUajvf+
vmK6UxL5mRT5pMPUkXRVRrBB13OSU6kNKDqR1QfUpZ3nVmnwID4JCoesagj7LEm9
7ocwBmD6C4E23xOXEWqF6yCKd+hFKEDSOmii8/WWWZMIV4+nfmhmWcI9nVS8JeCP
6h/EJ5q/rBjK3aHVPE+DIWqQWnD7AaIyp7n9C2zZIbxkt8TosLhS9fn4UCHisVx6
5ZjVW4s1uT7n7pQtnIs0kOyF98Jm+8wN4FExBPv8Rmq/yrwfcc3WO1W7h4ecNcf7
4PoMoPltkQRlcGPf2/Gic1OoUqfw+dUX66qSiRA8/9JeTOmkzAdlhLkOwFVwQqmm
0J3gKjqNgwXqDtjHJ2WFaVT8rDK02FsquQZwyO8RpTFKhibZhihHCBFchxByUx/W
+2nwL+SvRSe/ZFvkHtCmGQmNmkAmkd9jOlglaoq51HNcblIeulXYu9uyVBlX0/Wk
8U/YdJVNK7m+mtjz2JsOr6SkF3HxKyo4+Im4Hd3ZLPbGIA76b2F3d21fj225kvDT
t88kI2/E5mzwcqE287M1o7CZI2/Kw37kuGQwQyK0f08UZsfdRjhHtG3XAqtIKeFW
tdgHTdj2LyHRkz6Fr8bIGZ+UgdJRewx63SwsVUi/jpqfkw5kWZTlK+f3baRvgFNK
4JGUJvf07ivlBJ4l/9XbEIxifsU2bikLwsz4x9+Gb8D5MAigfdpWFUOiOKfdqL66
L9fNwG2gW1A7WLMqeJpb+kSzMp/l9aZAXXUggz3Ri9m1DhKkk1j8JtVv8Lh/P31e
RAsE1tWEkH4VBczdTdo+nf+XbdlnWfrpjgTTPfuyFKkm4t0Cf5eOH225hTX2U44J
eqn2P4hIAZZHSitZDSlvtnwRgxKpilsKrZRCLzp3fWTWnBWnqLs+eb0HoFXIRA1O
FxMzRoP4NoV3feyyWpPAogS3FDeNEmZJ7jpaqlq7d0NITzenQZTGOr11MTj3jr7T
6Dolxi0ciAdT9ORsXodA032WlhqJqkXlTmiPt/7UPzKOaBjc8gmNOpkczPEdBE1o
oiryqGFFmeGi/KeWiSpR9sNIkVvXLKSNNdEfcpZjRcSxKKQuaC7AXmO0a1njbhOj
cjnm1lPXpWk8TmTk/poJGUDgXlxX7DaQ2XY6mGDF+bFmU+njtMcFdwpa/YAU0mrI
XY+tQw9fsdvWPD1jNK5J9+79NRQvoaIL7Du+S3Z4d0h/sBRtNjvHHqXYALk8BbG0
72QLvqbK0CuJQW0q3ZflOJ3vAIdI1EeFO2lezfldORvdzLfsz+6gFAjahO3sJRhN
pPPE+FPvqUluHEOmYSr5+a6VbPW8QgtzT6BJVlPzPZREFFGzg5h79VJ/7Vnn0HdI
PFd7AGUmUv3fnfZsoPwG/vk4/VMBrOZ6kX0p52TyhwE43egh0ICko7uvyhvL7807
BMsMbC94I5pOeuEEUJMM84D2LNjNc7dQ3NOE6M+KYDro8f6jxfAuIHyNVFO8EKjX
ZpLZotNQf6ClDBhLcip0xAyljeVi/oZ1aBxx5nDF4VAX8jate8ODSFn27AkCP/VM
T4yrPk2QoK3HmjLLtY5DGiZ2tsPupNtW3wFYjchtsD2B6yj4W/fSodcbSaVWcaTe
KpCXDa3Qks1l+rjAorUe4Eweb6UPtYxNdWgGhiudQ9cT2NL0zZTMCRbDIM5h6UZO
Rkkjzid+RS7fXnZjLeGjvk8ebmKz6SHJle4f4mf2pGOfimGsIt6T4gZrvI0KbE0M
h4ZOHIVDr3/BF1rHfRhF47RFsEoBkFD4MtxK+ktWT+zhTYXqrD829VU/7tJFFRB8
qfyBPUMDUpvRIiv1HlAGUc9lSAs0obbYwA/0E7VmxvEyDjXz+T3EtLUNxhUfN60+
toaSYwgLoPrLiiJWqvpcPjlk0Aa8GlQw6Tj8YkOij5gcQDlEkZ4xBeibxUV7jA04
77omJJS4N5RJKoL94gR/fw==
`protect END_PROTECTED
