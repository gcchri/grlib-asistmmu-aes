`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Q6Lal7i1rn/OTwsqAV5ETQDX4AZ5sqIX8AjqT+g7tLvKsqvEh3fixVuL8JCKU85
RYU/ePnxTaJt0r+E78gwGhgMYtQJZgnuPLmOuZfS4fRtb02q+BvJuGlmA+Ry/l1r
G+wuhc2XWlIxQrjdjZUsLGruKvwrg2iYnI0lYGEzwUBDHQIi4CQlAvWmRazuTr1X
aO6xUgeQy+Gez656E9Ap6hkdCXRdbhx/1S5DKj9EJ2cBHoklxNx4uhhrLyWy19ln
UMzcHhmqY8fxKBIX4kyKjBBWMI28/tlHoRcbXkHJfyYwOlDh9nuou8vmlhZKyvPW
yKaaB2Jjz5hKz/j3azsOTqbXppvv2/MNoCGTYrwLvKIyg8ReAd92rQISPVcY6VLK
qkUtm17hVItyFAdJZppGiWQPyi9yJlbtidJsfHX9eCU=
`protect END_PROTECTED
