`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZJMOBu7YUG08tC0kgurOe2A3nOakhW0a/k9lQ2ZMleEsBoo/2XiRGvPDARpvwzN
B1uCXXHlW+OU/KqmWh5guhvmWpAQHu9P1HFjpvsNJyax0Jw3/68KbXF8etjTBQw2
Vl99jSPCgFXxtpv9w6h/r5v9Pqsg/9+o99gvF/zZqr4Cr9vYK5POvssxlzGlQ2mk
Q/4+JODjaJm9thQdaUMCLB3utAL59INwYXV8+RyLAuHYDoqenZFGcGzgHVUVQVy0
0Y883nO650G511xofTlXwKmNXPCQVZe8wqH8KIn+sfJN1NZjbfCdLsF7APkHE4WW
jpvRDu34OlYE36RBjVIJ4AubRy++bFt8ASpp2CfEzH2VOi7VJMhf/T7c9vmnz9W4
Y0ZtTPW3i0UfaWFTTptsonf7o1dIIgsE+ovAm/eWFy0OS9t7LgmmVF8sYeV1AW0B
UFCwHqvdcSqG7LjfsnMwjsEcBgP33NRHfWaaKPle+1P9fk9v0t+gc7TWLS/hrdh8
Zkzqocbp8P1ynTw+Y/BmePCnePUVlj8KwmUSqUYok+1688353x8lk1hz0PKpaYlW
6Hjj3JUTRmnua6e+DLnvwH1J9hmXgrFfdfp4N3iez85JRcVBsxBcwIP3AnYpQ+Hy
CKV5ljg0xjyrUFSszUPuioZ2wVq0hmXFU5xOgRTfQu5ErPCT12FanDuU6Oz/WCds
TLJVPA+xelfLelmVDBcrEhV8ZMR5UW6dDjqMcyjMrQtI5thRX41jFl7oO/supeRK
NrxtsbS2e2wjno2xZQeYlhz10P1QP2f2U7VHxTLVKxk=
`protect END_PROTECTED
