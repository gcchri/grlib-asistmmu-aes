`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VO0ASs11xxXGPneGSTiTtoc8AymlW/WmD4fmnViaZU0zI8IFY9c40nNTUXSgUIgm
CHkARTczhHKSOs80hRn1LebTlldGACnNTKjAt5430PdCFsFEJJb1TSwaAmgK/lek
Jj2T2FEtD6XjTyjRCxWVPojf+DxcZWmEZdree/YEjmmgRKeC35p5unkbCW261QkP
5S/UR15mruC0/HEi1Rp88HIDsdyNfX8jBf5SeJw03n11I7AfBGfBUl5xxjCiLAGK
BMDRn1BAFu9PDuR3AjHu+NziU3ajJIe0Ekm8Vqswdn+5mB2mfBxeW7MFdRdO4gC4
1wxZNZ3pjIaYXcfgxUesqBI0MddtAPqxXGmwgUNJD1znkRlOJROzz84NCneGhE89
IL0H5tMI2nm7MncKe6dTdFsFu4MPQxSNYorwR590xGxtNrfZS7E1kBkugNdCP3IE
1xWH8PD/0XqXGFFxJU4W2m63HF19eqXbmM3ZRFrtEOsnav7NWgVP6wjNixRMYEIL
`protect END_PROTECTED
