`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kO91TUkMdw36k4Wh8PDql0GbAxnuRNJrF0t1KiIBK0QXnEJNlMhBJgZz0Hzr28Ga
SsGfxNOvvV+hzb5b5KTZrQGcLXf0OJR+JbWGDjTITodMZxJtkU9NfYsaYvh1MNyu
mDIatIA9oPhd56W++izW7iMapVh+IOznopHXj6cM+XNCpg8CJ11MuJbeXSttm4Id
5R3gWAbgfLJxi2uQNgwO3Rsau5g/qBX6JFPVYRzKkZktdEos8dUj0eDVINPI+Ef3
A8/71t/4VimMVQ4mo/7NP8qmdN6FbF9eDfA9RTOKC/QqU2fRxXZhH4EZCHrEg1CJ
ouiiU3qNBARl93hPUgZ4Sv5HHGMjua0FctMP+sVvx9bS7CIjCe+gkw/zdwriVkn9
6XAX+xBwze4Ei/9E2WbYwVaWjXeKHUe4vKQmCd+uB6teSJtWQWwUevZQw5qq4lOQ
`protect END_PROTECTED
