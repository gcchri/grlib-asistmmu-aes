`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mM/Q5T3qD3JrSdTWnuYbw6BLHWgb5FxqJejOAu8I5NGY4MyemJFtIkpBatgdR9tO
6fLDPzRciny0UzhzVRodizOQNkedG1q6dJ3O/TejW4qWK7k854D677AwLIioSIub
9bSBBTmwEmkR/sQHVvuI/MEq9G7sTrSJOE5XnIProCjtI1LLCs2EaewuQuBZfMZF
yWUlVqHukS8jSDU4DI1IWR0Rukdz1U4E7+uF3XLcPoLpXKO181faeq+H+DsdeOR1
B8Ppi2eoYuY2dCERdeGCfQVnjjBK9XDnUZkXkoziQ2smreqJJW5RZR5wmbnyC2TZ
s81979HEaNWuPR5WxQmE1CLLshiVvP1eh1btq38chGPL6t0mY6/7oWds9CZN1ojk
+rxmXc8q0NhvS4XJwqmVMrtQDj6tPxzh6597/RRBTQPPkszb9LBOXApduBwjlzfu
Marre0uGJ6zW4SDrD8nBoISqTU4C87tlp9EbB45eczykmM3YVUShe48lcfC+m/SG
rq8YGr7HEL3cesWsrfMVxPLqcVukKXbo5P0EVJManUDgqqmPdB8Ct6y4P3JIb4Rq
801gVdpoYbBtOWnzomTZc+m3IYTRk0pny3AeA0z9EyJqO5fWfsx7ngkjzecF50JR
p8c2DqpBkXx7N71sLZnWJdmPbqv8nKXvvLOTyOchBGpBTn56xShjMcRTUIelfm41
VcxaU5Z1I11qblS8xu8Hdn2JPyFPhih37hmMVlzkOGLb0DNb8CW08AUEXn2LKD5W
vI2Z6dTI+xfGsN4aVVS16u4JWz89UJzvjsRier/esm7X2JKXOFFE3IuRFwONgDn1
a3rZT3vYTt/XOI4zyqjpLKfLt4ez+pH3X1LEroZPGZ2tyCfX3ZKNosq+MaAo8Cbd
3vSYWWevobz5LDXNxZDXhMtr77chKKE8aPYwhp3apPFjG0fDeM6xLPbI6oIjvYb6
FYerade9z81hjhLpQxJjCpoBGHcDmcvep5u3ArRme/F5Akyt6TTW0kBIjofMyuFW
bYhfBJTBL4dpWRedLNA/zKRfaUdRhVRSK420XioPHY7CJLZGM3v2cO6dhY4FA1Ep
BUEkLZbHFkAzbeidOFnqHdniT4lY2oAVeWkiJw1fntOCJJqfcdi+hFSjJG/r6bNf
4LmSbbBpdGxLUy2/FICD9391iCne0wJnknqL2+hSxwkjbkQICCwIH9IPw6BK51sK
Kfw/CRqel1eBtnbAJFjkNbJ2p+vG2SAMKKnZH4ivcphic1qPUmZ5xhlhohZICM1b
Uaq/uOrSokgCBLlvUXWVBY1eFVSGSxgOBEv1DzexZrEIF9/irzN/M3KImydM7gM/
lK+7t3SdKJ34uEaf0ytmGe5YMJrifjYphXj+vUNbQmfvPx2Hvv8MneMANNL8X7vN
WfI4190RceMuaPUxw/u+SCQ9EevTbD7KfWDpVfIDo4l6j36dzxynswkpKK2u5XD2
rX1Fig+tCH0+PVhtiZfLoDPpIiiTFNi9KRdlCU0V+V5TUpEQEd9QaDLuag+0WaEP
H2FdDBDAbSKG1gLQ9Y5B9VxAgZdvO9I9HSd5LVOxCGagBuX4v+oWRqLdnXhYt0HH
M5zfd7tKuiSd1oWJRk3W1UTsOnfh7+wZjiGvjYDjzdY71unSXTqOLI/Lf9E2NITK
Xwp3JJikE/2Avvwjb5MgWqgt8QTqUGvvfRHI//rjTXzgF0ZwJKVxS7vjtSfjCXnL
CMlZWUwoPxkfR3WWN8a4GT/e8V9zLeb/hFknvbl76fey6CBNxuG7IOnST/ItWXvr
pd0fZQidO38+Hm8PZlx5uWGDZYGvIL0tKRC8lJK1dknL37CW8NhLeIyJ+Jkoh8Mw
HwhiAauwYuhYcJJsCuU+QjYUkGTYOU39PdoP0WDVBrV+kO+A9cWWYGBTagwbPwfm
`protect END_PROTECTED
