`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KTfeaJb0/uxLqgNCKFwMNcp4qaXufJmXX73WIeZmRn3mDUxP9lYVSa5ppUMUxHYi
L/e4EuonI2xXoaV42C1KOl6MBriGg4biMbNZ5hEd+/7ur3y9MYNs59auRM9Law08
oTC6OiWt5Hy0q6mVGKILKYkeOx/uQeDVBHzwrzs3sigMnyLhhyeM2KFhVTxWzikr
dIZxvYEdzIYilG5uxBwVeWPhT0TmknAfI+uIoZIUJc3Ww8Gp6+WzS5PejbRJf5sz
Q3dJmE40oxI7rOKFXTfbJ21jwO/NedEgs30ZKNBQWSm/bgPSLYfjMu+Ar/XHrGva
S6jE/FpOrjZfw6AvwZs6nmQQYT4EL6o7mWWuF7OH0SoAPhRa0i+T/z4BRKH3FUtq
zMSBcXt602u+pm1jtoGN8xpS8Q/RST2pqUBu5VYzjl3ikAaciJt9jNcAQJXutjmo
kmnYrSuxkcu5rB49TQaJR/Xg2T8BJ2Z4K+AZlYEOMkCyn+ytaDbmqV4M4hpK+j9W
IJgjWm5TIvyqlgv1e/UF2D5RBUV9cu53hb3dLsKvUHE6LEnJEBgNl8/CyaMqrwRW
C4kVFspBzG1nx9J4TMP0x7jUkBJfD34hRGrrzEB/5syo4SkIXk53d9LraiyqmMaU
QAehyGYAt5e0CZIOyOe2OA==
`protect END_PROTECTED
