`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m4pQlBO3sqRP0KJMKyCm5H8XUnf+Yjgu6HYjjpIu4zUVO+VDsvKiNCihP0px08pV
fpx1YAhHc9NNMwH7dQf6YWVaNXKwpXhCWV5IyQLlY0bAW1CH2Ya6WHYruYyzdmz/
rjwxKIHAeJEYmXfZUk7rX4GV54WdpL9VInmS7aJ8IWEiOv5vndmIPikg0PTgpp3Q
GiOFoMy75GCH1V0rOTJ44oPHYoA55nTkme5nENd/NaCIjtSWm5AmPs3WWqedRAFR
frm95efzP9d8sBl75mjYFKo5lGoPsI8nyQHUBctIu6cW9DieIMNDrI6wvGyr5x48
x2D7/RB1o3FOPEi2Ac52NMgMacuhH4vxH3pi5eB9+VxNdCLoDCoPVXj2p85S5Q+7
RJm/A0gpMDIuHHQr95z9WIZcukkKlwC1hGZ3ls6gesGoAdx+VomMep4CyppqOdbi
OTj15aYd3MLVwVoJbsLw3InHEXuUDXfObaKNjxl5gqBuPKCkc71qlQSkuXGky/bo
hGMBbVHTFNQWUJTgNuEEtgLhvuxvbwRJMTVA10HsrI2NiZGwZTawxn72raFWkH20
uhfvhN+OsRBcpXGm+r3mkfoc4bumCWB2rwG7AmFHVVxJS3JWj+GZCBiR3+rfNRWz
ANhitOsGOBU4k3Ayo8PQTAnFVhNwpiX9p3+RtFtyyKd/MSoK1PbYMq0m6dz2fuge
9EcDYF2f+emwj5XtSqs0RbFOsNOD8ErUeRtUNU/zrAVu/hW6gSbfJigONAIZnuRI
uK2H2xP3aSE5zOxGZ1qeXUnrQNDQkBDeXKrJ6SqHTV7M5871ZzDlTKOV0efNQ+a9
IuGRnRsgrGM+MTOzGDp2PaytRlcRWu7xmIE9VdkRDM3EcsHT3He1SvMnnyJ7Rpwt
5j25hUV8oPzmCGFU5xsZwJ84ScDvvAakQGvtFuz1PopAPqnwIYZE7nY7NSFkS8ak
i47O6d7YJWIe+TCinJIAqeWlN4IHmBHpb9AjnyjEhx2Hz9J0UZXjlF9Y1wCa9yJQ
KZWy5ztQ4Vjv8THsjfSyZ2K3I+QhyDlTtRLi1OIH8hRBFc+ssgTWSUo9BG8bFcFW
a4r80Bs9nzsr3Vz5sqsQGkhOgBH/Y6XHybddKdtjN4SpdxPZXI4mTQIFtz/tLeVk
co1tXVgCIYPtGit8Q+PTKTlpGRnQ1sd1q7Za6q+CIQyZ1puccxJNfkNqMilljNPf
M1Uz9s3I/acgO4VETPPeb8L9x4SaEfPygtdjXPibZNE5mFt71cs6NqAe5TQJmCUY
UvHNszXi3MXBP003zty/SF9mSz+YSqzWvMBjRH2Zq2/lUz+qvJO8Vn2Z5vU1hXvY
m+gMX5Zk4HB0F3ObwmBd5W0J/xBVy3UeV9+X6VacEF5zg9iDBNGuyiosGBbQrlPp
W5pz73kNTtc7rP2fh0GWzZHRf4JzyDf9q8LHltv7XLChZ2kB4WlHQqw9MkO2DNP+
QN5JYGzzMVFnRTl5R9BhjICzdubMyVSO9SECTBrIJd4fAlol7s3uwcluf2b+4WEU
VSmtA4TGlHOdfXHaxpk5lmD6YUbHp/agR1WnS540CH7QcOgdwUXGHgEFnrtBnO2R
t1NXXfhZnCV4PXRjKO8WiOwI0WCpJV0EfvOwrf9VMFdHwHPt2/Uswpd0NEKY6eEC
Vex5SDuK6Q+ofW6AHeZBw8bjnmN6wlnfkabn6gvSBnI/GzffiqBV9JaU2cg7KCEH
QnNTwDofNvU0m2ssYPwZrfd1qFeczAvd47s+VvSYoEYOPiA7c0IrxxfEyr0kZB7T
IiKP3XLfYGZLFd2IXugxxb2PTUfE+59Mqsy8Ma9GVC/QGEaLFazgrUL4WWutnHov
rpn0XK5P/fdVKMq8QxHhOaLH95V1IdXky18ArjaBDWLllWolAwAI/rOiazLeMKTx
ll3Z1QZJXsThJZStLNG9NEzOKq1LXpu+AaYqoFLm84SKHbCTARJdAsGaChLi3l6X
tqQGsfrMQxxyTpHPGssIZltd2gbhSyNOAlGPObnQFDT9u0nRBQ2ZzFu2mP4bJn8k
Ql8Im3VOEPFzONCin6rQgURsqCf1YKupRmYWA09jSUTj5Vs+Gjq0W8UilrNUujiv
oIYBuvzSUfGdF8ENuTOPawMRgvwrhIegFheu+t3LlYe5mLJ41JMDDWypK3ee7Sv8
zAaookJFiau+3cBOHThYNYuXsdFDXlRda6SDa7CN/6wsV3s/MicwlmYIIQB9M7h1
x1RX7I6RsSI+6XxV8nIlGa/sHWBxNZzU5qLmyxcGe/7gGVxiAg04/XBd8xSl7r88
poIs2rupfZHLNMYuJptt1Q==
`protect END_PROTECTED
