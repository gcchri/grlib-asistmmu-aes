`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h6pxQpcszwV+x8PMk0qV6W8Mw3dhqTw97cc2nXgKwEWEPDuzHlslHBhU8sYrFwBv
HFrM4BzFszsF7GKI1JCUacWtmwlnS2+iQsyeUeifEP12er+aNyay/NojbXids2Au
6TXv0DDXT55ysaJnhi61UFfbkgC1eXWeTPngYzcwJtkvdOesq5nh0hsCnK3jO3Ew
Kt5ImopK6+z62UE2aw2j0zU3FZxzUnI7Znf485Zor4m+K7Y460UNP6r8jU7ofXcS
e1FU3H8HaThGKXmnDs7PZlfC5aC7KQ4uvq2aZWGYIIaz/4GtpVRmplEhxWVyp1Ln
mNbJK+RoSR0GtBI17saaMAsu38bzZvim1EZZHb0RWMO1/ZBK5WmuDJKCF06k8HNU
sYw5JnChgz/f57Ttquzqu8UDoDEuNPUcjRPrpTG+grMx7DBnJFgDQj3DSSsJKUaE
ma4blyde8jVfRFxw5Emxe2Nz4tvCVhChzsFENqtZ14OX/RpYNboezy40ag8aMpFp
R2ijqvcUmNMJLdcTGtHNfv/G17WSsLcwlYpM//5dZtoaLoiI0pJin9tZ1AeFNQnf
Y+tVirMXnyNHsqLreVYKbowftTVFnmmeM8DBG6VlFlpr+tulPn7yrXE+DP/bfv0c
1TTPOG3khrjyRHLwOMdBPLRAKp09sVYD3q1EHGNvNK+MEmLytQd5yMVG9fQiHTls
ulW7xvx1c1GpiMtFumGWU/TnCM334U1LbZcpGNwqsWgLK/0/0qNv5kTlkK6fAPYx
+deBs1uP1Z55h7n04Kp8IMJMjdi7alv/PWNGpcEzyTXAa59/dbFbOYEaO6a3Acuf
L+JBkncuycWTWStgQWvCz+596G93S00/Y+rzbSgXX0ungwmN90dcP0wvmY9WGeHd
fkpaKzPAp+MS//nBYkjOD5bmMdshXRH81JDH5SoUhr+JmO1rK06dJEmkayB64A9D
T3Oq/z7cMJxX5EVTk7MQrlHFpSrz0LDW81eq+EbM7G3K6QZJD6lt4cHBbAFtXYO6
cNjmYknFs5u9ytAdw+bGy15fxUav7Sab4JKnj1F+9jXkarWJIskQEFqHtqP4l8NR
hPzyvBJdGOq9C33D8L894XxFjWqMa9BHDWc8cstEIPCifvydl7pRyUOOGCnjCEqj
jyj78bEsIbqlNVtAqG2VegzXF/fcjvRGRhxwIbYQHogLDtWxYP6hOGJKPrm5/D/S
4ajXXHVFaMLeY4Jz7Ce+YANmadKu4M+fP8nhpSlHrMMr7Ah0rGe/HL4sqd5yaR4s
9kWiujikbTGarAHlU4LE7hJLAE3OynO8my+bcm+7xZ4FH4aI/z0xsWahH0jQi013
Cpj6z+pbKTAIMyH4icQb/diCcD4w1cAXzd1JdnHwwKY5yQECfQbSoRchp0N5REx+
IpmI5jfgMt7ZfvFdLS+B7mJeTBJjye4M0A1SDqVoH+eZj42fU5IOlKQpbsjpy1qK
qMCXp3HJFnZe23AL+I9+zqneAe1H7PFJK/DuKBYFc6BH0ejQ29sfz0TzxxQ5FkCk
fbUuDlg7QpnbZWaZ3BheMJP1mhKHlxeeW6ysHUTBH8P1inLxuFfV/tJyxs4tNMp4
vNjZUoGj8Zwx3/tz9Z6raeWLsecAGnAtTmpjLxMFqBH3GHvm0A9XVqfT2kqzMrz1
EszBrnUTCB39BmioCdU8/6HeMtwnJKkkZ0a8CPTuYX2gd/m6c5gM/j3qNE3uVvPq
lsIr973caQ+eHcaqxQdso5cKNryOSUgk+UDbK4njOAfoEUISTp5O1wImd/x44PHv
QL3MyMLwZMv7A8DfH0gXHFOT6Vqt6/yDygF9U95kwhQA7TOg33ZzF9T/U/S2rv4u
KBZ7L5ArioPmXrrSnffxmM9HJZk5Znvfxag+NESpLQB5dEc2INVZRzs0zk+NQQob
Fm/WrGNcybMn0/fvOXniey7C9//gSakhVGQsAh2jqfmQiIHsrHLqEJ4oCVorz+8Z
yedk0+ESEar1R9EHpi1vXvJ2gOR3YB0olySYHTuMpLdX59DQ0Iry00A//tZGjWAT
htnrziIPSGlwTdP+xuG0HCeCDRgtlSudAid2PFG5/AK46+xce0qu4z5gTQajlrJc
AnUoYWF+CmFJSVFcHIqWt+nzQ0d3S8Fwo9cCtIaZmW9OgcMjvJvagz/xjqh3cJCI
NzNsh8GPwFpRoNUKnqNbZTZIi0R+OpK7tUZlDt9NDTOZmUCnCmLsVq0R0eW/72cv
lrYbBlluFmqHHbV/ynlJJdvPS4Yjw6KI+HSbsP/7M7P1ZYXXBcKLq/BNyEXXVCLx
Rp8MCQWNM3OovPjHQbZ54BEoJYw2ucNP2YbSUT+uT4ord+R/Ww+t6olZjGleocLK
V3AyAHwTeBlJSUlVLFNLJua9UZFj7vDLr9mcVFHB3TEa/M6eCIBdkq7kOUfCmlmE
+qA3CCbiW2DFcM9NlOZA1EqymycgqXOeiWaestvTvQVd0Yn/HR/jS6pQ6DRXuARP
uOceNSipikTpMe+6XSsgg88XeUMcsLLkUhxPebQXPWV8wIc3DjbE6MKeV3ZxyagV
GOqZMX9bkBZ1icFUfcuwUWCNIiE3mhLrimymd2YmNqRvKS0q8OHtPw/qDxmyrXqE
KWm5thi+05IUV1DrsfTTzz1RLh7xtoiGmSStzfSwhzL8gVydb1LsLGlul0q1bIWM
X4crSPn5N3ZzWihR/GX6BsBj/+08bDgzB2ZBnomDDaMx4t/XTCgkGTG53lgGAawh
Rsr9UdMRCXDvJgi2LdpX4Y4tBJK/T5E8l8jGQ68JwLEzXwvNriKTmvNJxgRwwZrP
kRPX5mm0KyoUxXBxHt2AT9/msYILK/YwuvK2uJPRlHD3E/ibql/ZYPx/DbXpEYWc
MxFIR4g+LunvQ1NEI3RsHyWzg9GHS/BQAVDV5Gy5rHy/gjD55iuiTBNVbVemvRWd
1ZUKyNUrlMswOrmSqQl7J/EQh549FfLHT6iLMLco2PsTurAv9mW5uIT5LeV0YnKW
FdwlfwJMFfLatJfX5Ri2pnmS8Ic5JMbaldHTUbwetO4GNVPfHgqx7x8IJWXmfbgB
/QBnZwjCmzkK/tNgiapf5ArTkX7uphiQMWm0zVi1mRx+hmdwCRWwmz1gakcNvm1c
ZaRrb0w9HW/AqYjxlZNu8XSX41oUsZ8k14JlYYwnhK5GCnuQyO8tZ8ws4/NgmVZl
JmeHwUT8DLh8PflAJwh2gJWYxD/gyzZ3P/TJWDq/rU4imLnzRZ3Cq7JfH3dI7SDw
Irxc7cVznSArFIFMeBvYeoWjDcrqeIMcoRm0je0oZrvcwYN1PZEOBaqV01ABdGrN
b1VKQKZwKFDYprOz+GhPIPMED9tE6nJdH/5moeiR6We+3NW30BSXdfUSXU0rMuOv
Tx5XStEqklsLtzKI7cQUXS5pyHYtQv6HkQz6PxhpVN1ZN1Wg6cOeJ6WpuSzgZ/6C
egBwzQiEYlWnzGHA1QF7WTg2MNEckjcT6MO8cUgf5PbYGETzhDPQq5K8UHMuG17p
FagK6IZqQP0HLlmIySnUpGKwQtUUWtWbtJUsp4UR59PJTJr6IoCs6sISd4/aaCIA
yvgiUqP0NjE9jieeQJLjyO+r6BG80w2oWXn6pYgrxYXMX1AuKWN7C6iZSQfDk+6/
rgmIHVKAcP5J+oXa9FEgAJA4EvPgGtwo3Xxq7jlg/CLyH3GNgLIocSmhLrZQkQj6
C+Gh4eZYZ1U97uRLtw2xeX1gwzmhlKHJ5KRQUESIjEKvrWSDqoD7r9L2DU/c6FMe
gxkPCS8dN5KzLghC+TS0YBQPg0mSLkKtNuYdniW0zvCgNiI0PrMa4v3Tdr+dzx8E
QSFfRysmr6yjIL+N/Fne3BqD+u/DvmCWI4eID48W02RtnQltaQC9fwsRw3FBCDeK
DXtyHi3bFxQyGwsAmFI+X9cfPDdWwotN1z8NEr/jB7ABPu8d6PPtNOPmyvSu2rSL
rYbwMezRiK4cQQnPrLL5gi1FS+TloncX3rqdJfy2gn2RlfQahfUkEabuE83OxUEE
AQK62A/mw73DNJ88LGA2wmIGsNv75F9EZDobpmeGUovsehEQWnvp3bQv6rwr1Lja
1e3zPyTSbuh2aATgqqw2DGMnvrX6JbmRF+Mmkw1qDiNjp6n3TBL2fKGcrVKflQxu
FHhcU/zoee3TzwXcGC4FCpq9EeFrDLu+8P1sTi30/AkdE/7/DFdrgFY0AXhKLeLB
LzQHORrHCq+tCb5BeuLeMEHBJY3Wl0qsvDJsPr/Nmqs3tKTDv+6SmEjv5izEXoYF
p6YzRV/ID+wdSoC8XKVUummqHMgYIH4aZ+QYS6g/sO7gwjVAgMauCAbULfJA87SV
xN7Bnk3B7DJXIC07SbBNQOtru+vAqpCqNi9sJhukHIf0cEmVTxvq+6HPDv+BT+fH
34sBUaFmKvR843OtvcuVYjI7Xzy00aSiQk6BzwoP+VUs64rjkqfihDyPUPb4UCZH
ZZcB+FusHYgzI57IDIVyts1/CGQvIMm9TTPdFtM4hn0Luo9nJEoKrvdtH9Ffxnci
1aqarWIT74nNUnedk75ORW9ljc3nYl7LkFY5B1alYuh1YrwjTmQfCcL6aBOy4yLr
lyEVPu4zjhnFLsj2TVPEBAHRKoO+ZDEKIShWXo+PlHb6J3sGMXRWAwGmEK/8hxi8
hIzXM3Rq7dftJkcTAKKKX87onBMPOcSRgsJD8+jxxCH4pooilsx0SFwU0qFLPtAC
j1yEVGjHXMkUJ8J9fUrGLSxdXBRoG+XANAT3w+SCgxhvaWCQSoTUhjKlb5HXHCIa
SDiDPYiIRqktGVG0yQR1CwxMG+QrG9MGErRSx92y286SmWEHRhKjL58jd+ELm2wE
q7JS4q56ioOU4K+8vHBrfO9cXWQwAYVAvFauI3xpAkBtbwORhBMvH9dyFlXSAB+4
iIj5lUBaVKr8qdlz25cbwzHqHew7lAb9D9wS6hzMg22UswKNaOQtm/MWtvaoz5QN
XOmFMaJ+AVfWw80aDt02xLT4nMXFQe4VL3Q+nZTJNpWOaYWMmZwJb4XH1LF0MtVJ
I+j3p9zYrzruw8pf5WVjP5T338GT2bfGMoD56FP+e5AyIIgBav93UmTYvFNkLqZW
JKnmhqIT6PDtB45CgQ2YNkwOvecTMyMYvYGsRhhsst81TzKOFzS/IylD6bUR86t+
n4lv8bBnFw25CGiMQM3CvxZgv2SCx32lXMnQX4R27OPEa2dOjqBM9equloQWwPdf
17s/9VJCHbTorx40VkK7QVJ4mVE6PQrq9lI7v/NSzRAuyOo5dSNlW1nD2iFOdGRL
j/AwPRFEBgECc4xo6/JkivXeDEfshMhIKxp6eOUHmvpf51ljRGwr8TBhL/oBQUyQ
ilMqP8PoOK+yypDtgPz8yXoRtVvpBGQCE19Xb2Z5jsIORBYzYboorNqWLbd2tq+G
XqL3dtcePZHhdM7cs3uj9Zi2fZZDxBRtxpJ9vFIXLtN5tuh0FEXW/WGyhMkPawir
ComXgM4+KJIeGWmuNUbPqKf8z3sYpJdd2FkVswC+4s9lfGD1Xf6eDwuqTqdvPmDP
ymLfviNJemx28Haq9OCm9BSp0d+fAUmtwozV0qak6FNqlruHPX09545DSbih2xc1
CLJ4Ii150tEVInkAnfUzrzGE+R1dTNCs753ngDVAQINQ72PIAq5TAwcGpeQjAy4T
umtvX5uD7W8JBJQY8K70WIJNFTCOSFCzlkfbuS9s+35aReZeJMuSVZSJ9eEafJBe
uQqk+h7qZGPeDlSjAklGQ4kDI5WV0Cc7B4zT82zl9bA6gBrz0sCp8CATNg6dJazZ
VHU0mImqTrEMr+d4GiExXJmBLJe9Tz/HBjAOVFpUGP7pq7MDgu7zfh5q4/Y4rEXU
iehD2iZeQQdLhF1C059xQTZ3nAls5VtdKYY9ZuS+NBvG3C35PLGqCk4xPNmtnZkx
+YqX51L+d1uBuklZDwoy4IEG5txsxhgZpWhB6siKM+5oFccSfs40m0D9BxyzDAmr
6oysX11DnjJwqJADMys6s58nd++9+6nFxb+kVKzEvDJU3TumolOwkRGOoRge3y/b
ubhRuDI57nTrC6q5FosBtZCbh+uXmhFZSlv3r28XqqzSfa9PwS8TN+eRlrvxetRn
zdQhq8SlbIcj9LeoNdsFujxSB1EUoQ0pIjrtCiEcTzrVKpiiYtZ0dPQzuCwlf3An
ni8l8FoF+uaGrsgQ8IRoBuu4FA3QzrXY6cAkB5YkQdd59D2k0Lz5B0gEAi6DFgyN
RIHUkA0QOHZBunIev9XAjMnW/BNPNrJohCQ1WLAXQyM7vF9I6Dt2Vke3wKeuLoFF
KeT2DikAwhDYLrsmvE4dq+BLxN3vnEaPjVbYNAORx/MiA/h+UXRFz5O+eQZqQFhE
KJ/AMjbm0sMRFaguIRFl2ESYBpxaeBAAhlCikHW6zyfrmcc40tI65RCRCp4ktQCd
lkqosV5sPwEaitdUntfPlzsUlVzetjgB5C6NPcrsSs421hhwuSbjY2daKFxOmPV4
O2kLYdm6TakBkehGFAWKAikRnrQFGt/RMtSH20JWWPldm88Ow2rh2F4D8heCUzED
MG+tNxRWe4mIVmnprD1CssltbMdFAvpjW7T8TH3DqhKk7pXkgzgBC/AUU1+uT532
hCD3cwsUDBPbYYIYlgt/RLgbItFvZsklgtiD5/L6b82pROD18eQezPyDalsGBi3J
V2667wFXu95U5ELtnBnzB6eKc7lFP0H60/1Yyrz4H3IjG1nwyi3s79QQWnbFx5P4
32RiOXdjfBL+O4WtEVefxZtnTZGmcbTDwHBEquah3ykHV81s9l1wwrdS7SV3xFVv
BI5cZ+Xj/kRdbMWz+S4oac2MUQIc5iSIeqbo3hzZ1rPfsIlqm47QdnwVJoeqrMmx
f9oqYs+lIycz3EA4gMRO0KkRLEJ5cNredFyakRSNNYApJ83ZO639wRvxHOLpM4lQ
E7APNFh4a1p5FZCK/1bGV6ZfVJYiwxGKW3XlDsxGdaRbiiThXbQRAWwv8wogQsqK
S/pOqlMvRbJ3VSA5xPcIpmJnqD7eaYTAwsYqW3gTHT82DzcWLyCT3VyEc468IFvf
1AhtxxQFljRWhf1eMKtCef2bZj0uaBpoWlmqdW3j21+widSiinr1ZE9Lt9W2zCo4
r8p4BKLs95nhUJjAyAIzhyiUzsY0TYKFZOLABT+1kb15586un7+q+fMavoWRTDA1
FmAKXZAAAHkUUjUutLkB3lmku7xCL/Fl+E+ypaaqpJ2hy+X4eLl3QYfzs139fFPt
LcohdcViK78a2LaIW1wQ5pi6wkWxaVf5DN4TT3+JkyeD2f6f+IHUONAeEl/wHtya
V7HBd+mcH3pOOWiU3OTPgf5o/VpUg4/yVjNBUz+3M1W3eOE70MH5mEdfRtUQdrlj
jSmfpPm+UWXY+jMM675jABUw3y0z4Y9suk0zfa4uVaPHCC07wsDv7SOfD9DQ027U
wyXPQlqLbxig+3MFECbxfGMdZifLBf8T1O6ATXY31J2Gl/ta4TLW9+xfkdHAWiFW
DEcxy21KM6zPA740IuALl8mHabXXyC7TTqy7jRTUlsurUPiFMOXYmnI/OAT+COlM
aeCJrAqZc8zkHo5FpgspAe6muzzz4n9d9pi+QOviV7cn/HLGjItg0F8T13OkOpCX
XEIeMFxPR5UT93ZzdcAnA+fYdlMCI/ZHBIip0Cy4nivZkQnirtzrAnu8cDZYjLZs
MKpPvXE9NwHdJiWrRZZKdlZrgCvNHdnelGKuQbgOyOmlwQQeYcDv0UfIGOPKRijd
1Q7kONHpleY6foB5C3cqWDhNlA59us+/erCS4kzqSqK+rxrd8IpNf1uJJ/RinDkU
Muk/gkTy48zsStB4scbBHtBzlmLasB/eVFAITBLh7XZZPIdlGcRqTDeXLRkSdxSj
iTXFa7d+M9SY3YCw4UaqReXakKfG34siYeI9R9L6NlQfgHks9J9BW8L/1S2CBjO1
l/MafSSGne7M/wKurI4UzLElTn/rTTiQzuk5g+rT3gVnL+S2rTdrrHmnup++LU60
Iswkvo4yeB/hP2sj4EL1dx5KglPN7OBM+v/CCZIv/dewfdnM2uXFEIn2xUAz5Njq
3TOMcQ644ZvOZscF+lZn2+lV8muiWniyMqTReX8z3HHa0MIeV8D6f2DgIyEghGWa
zkh5yR+pTIFdVF0JY+t2+Z3iOwrVclY8aM9Dj+gq1Rjnn+WIri8wzQ+aZ43KAd8N
dsf1+PZ26xijza5XOZKDry4+t3WEQ386AVQnxCeS3JcupcdFzPN4MkilUkJp4DVq
2GMAcECmHYBylmmfSOIBLme7OSTH4FNLFs//f6Bcf/B9nlc9ym2vSJx3jpTwKAgx
99nQ3k99qhYZn4qSjiYz/QFCkdLo8vUuDPslWKa3UOlqrjiuQeYZyu/wGGCNhYc+
DbdZjFYGIQugZkMMqHSE/kb9BYWMjq02p9TcTMusUemgbpV3olWIHq8OZhPmhFKS
d/fnswSY9cFSAhLZde80Udf1FH2lTOnGnYGADnZtxQhnR8W5sN3LaYKVgk9MCqga
gbfHGdWtrTW1Wx5Tjbd+RZPJOE2D8hPmsM6uyohCurj6qRxkUjhCHbY8sx68AeB9
adE9pnvwkUIC0C8pltE6LpFpBOo1o/fT5ZGCw4MKPMhmZtOmuySLrpI+dIcomCT1
+VlDLX1gtTd/3dmBS2HtP9wbJ446SRh7yYjtwUHdpDeQjyEg9Tp10OFyVBHhPZVS
4lELutKc1zQucaZLHtN3TxXqcGboG5XweLgpPW+PcYdFg7IXO3u3XljQ1JU/YTFP
GMLkCSJ06XtkO87zDoyyb1wXyKKg4neSO50kOSXtEYo8JkIabb/V34oXOumzlROJ
QwTKbWiec8obFdFp1DpVjQ8Rpd3vhj8sHyXodUuh8pS8OUFWaQRB/ObI+fmBz956
if/9lVAQsQGncNsXpSMuKOHq1Q8OHgnNaT0Jjqc+Po/LC+GebvWSWp+hCIGl9tlr
pZoebH9qSykB1z8iLm+M4rO257p8mJPaUEynL2wxAoiU8S78SJSIau4Fs21uDh4c
5GS5QU4R9k4b6atlhCeAgmeRepnRSp7BM7OF33jW51dJLipKCjPmfqW/QM8akTt2
B/YkcjnW4NecBBd4KBxhdPfSMUc69sCaRwntFfGo2iZ7eUwbnTv3KZJupgFJTh6i
skYJePC1kOxU8OpeU2W/aj8H30agp/Zln7hzbLWAOGXKXJydP0v9RSwWJDQr1nn7
eLNW6nDombHWvmcSql9EY/dF/kl8YtTCARpxrK47WkTmnMf15hSEW+ORznCey7TS
wGB3r/9QaNhJQxWpCcmDaggeImYyIIAZecNnlUmhrJYdU41BhlVW0ri5/taDIRYu
0eN3J9nC6tx92xxAEvllKmkWFTuee0YUEwWF/iHD2efhkEXkiWlTU3Vor/hHjVRe
TyoCje192fwkIpE8Re5zRzkCzDP41X/ek+TyGuoHtHMcvtmmPR1692uqoAYsfmmq
eG2BQp5D2CQTX67t5vf4O05sVTE8tHlh0gGPa1sbu3vxTa+idKdrHtKARoOgIYef
//zda3QG9jCn6aMBPLTwxoJFRXy/uWkGlX9i+ZSj205h5gmAuDCBceC/zDjUjdxa
7tRgEqsDEr0qD9I3DKdOWQwrcFpfkeSA75N2vZoYccj2X51VvUBPRs8PFJyLH8RV
V48TGqsYLBgdNVCJD6tdnYnltr1zf/C/ugZVoB756kN/9qpBUsQHCse6N8gj7v49
i+IiuSwvoIGCXYhOwSebw624LkICe7fYRSQDKhNwtbFWTZCz+i18yYUNTQGeMzZ5
Rll9TE6NfaOr1yX+mwEnxJSx8utRamZgEznpjVPI/YjsBuqEUofk3pidggKXaZaq
XrpWCCmhicvTQSJ2Rmm1vlw5AhZk2pbEz7z3BVakwW5mEIG3g/u5p33ZPAOFh3ba
atIf7uDtErcYqoo2cZ2RQWEOIQ4GoCVarNfdYe2sVMXyqYwVmh9YtfJxFo607bmJ
t5+6CuM7rRdRmQwO3eJ6cTNZ0QRSfz0Jnps7FHoBYlV912VZ8iJhyOEgnDREDPZq
xuLE4AQJCAYnUzJMxdCCZA==
`protect END_PROTECTED
