`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKwckNCjIQ1nKBrTkFSgkqOly5CaKC/2pgIYkT1QuIuRQ9FanVH+0VFD2JXQcu6r
o7+FRnesD3a96Zain+KhMpOwSrlXd4RFSQEFJ1HdhD2OvaDLPD+Sd2io5JA2XGwT
UOXRaJsAs2ElLxOSsU9HG3gVZsevdOxb1BxDJQfJG15Qb4QKhYT8MgpFKdvAwW8j
vvgKZW0vNIVMIF3pPgLaDR2oHFl5qgiSu8CFwqp6ZnqV/3CvxeIZ0gZaXDigerpl
0lNQffbYeWWw9y8hEM7ZD9kenaosURfmFj8vwxvW+GM434wN4m3dDymFqHKNI+JP
3xDfsYqiKjFELbaVYDC2+3ZdiahdY0ReS7Eir0OinF0uTn1VPoKXcPhleZKrr8Lp
n0wmwDLrphO/ZHjfauJj8ctGaAqYRSNE+rsZAtGw55WZK9DbhCmMrhENg7oAWQ51
bjj108oDGhPY6bznlYBW85J+beNll6KJ9wkQQqYKrhs6ekG80/YvOJTeT/1N4eeH
P+WQ0XIU8XO8GHlMmQ2imnjsBBQuhqDAdSVPDE2hh+aQgI42RlEnhsdKGUd7REkp
jywevOdYTBrHredHUZ7Tz5sNm2SCYZ2+Zbdy/wS/zJNNdq7lZtGokDb9j5WB4ITM
b0033StLITIORl9dH/LA1qGEsGlk/4t81ZVebYBuApc5hPtYZc0T5J6sbpPzZ+4W
Rv0aivKtcNgv/ZDUhttfJKLhX8r6buPLQID9/yV6l4p6rwe9dsttCQBZ2p+kEIa/
jojx1OPLkDqUEZAjfXvU07BlA/PG3AZVeeKhvI/G9R7Opemj6+hkHpu1RUCrlowC
819JYJcXBF207xIsbLMGKe4O40JDVJGLQdK8yTXPD4jmyytOQNCon7FYgTECB0PW
xq9d8Ux4hhuCoi1TjoEyfXP/ocX5m0klKipxe7a9Gc43q6OTepAyaFAtlc3Whtdp
Ph3rQZh7WiOPKQmgnWQEv2xU+MvtKMJ4nM8gnIIH+G5Onn9sJn3OMiUzfNhZb9RU
tqqSlk4nX/A02PLbJ8hVU0j8EC4mWfeQQHNLfeIh5aRe9X+OjlFm2dB7xuPcvQ6i
hIWtR5vZ8iVGE0GDQMBi4MZzakCsfdRi5R4PHWzg3MvwLcJY7cD26gRRKYOAVD5r
hfPQuc+TSwsVgoqTACTB2d/L+IVTfzg6djJJRblCLY7vh9UepZbJAXK/kKDXX4nS
1mZ4OfvBC2ah8N82KwscYXXXbsjhO4lP49DTQwh0n379RAhY89ogtMCrrYNpbMnM
UqHJ+QWAB1SQjGujbC4kepowMvKC4mtR5/2rOXb+ltpTjBAji8fQqtVjJLp5ZtVy
eoDuRqLSs8BXuRyjVs/9EZoi+nx69FpmLjlDKXuzholKmjHJYiGQnwf/owrmXNEa
nOzMWNVwNKb5Xz1nHjbXnqdD5fMejhe92V3hd1GVtrxSw74O6sWS7D7WEDNeTHhC
tiU2TXiyxMnO7Kx/rTXqLDyG3RQFpxPRrwBsD2cssxhDuz5Z010aJvUUn8ArSYBr
akD9f/G3xnNVpC6HMCWat8AiJYrwqr4g7u+KlgeisVhqW41rfjIXpOQjDSzS+FVO
p+Gr7UPX8B8KT9tSnEuYSf252m6LqV1WlAmWOT6k2tli608swI8mn5+kxQJBSfcC
u9YOVu2mYXpKNRtqJN1l+z+10wCrxYInLptMpTEsk1JrjhIQVw89IgtXcim8uLvu
Jku5/XnUzzcb6jM3/aR9W4gFe1W/GX92QgFoFikikRr4e8i4VoeMp/momAIZDWfs
0nYDjm5DAg6VXCjFbmxZfB0RU52cWRHOJ6p1ZM2QDuHmkdxsqsGkasFViOgFF40W
H+EofOi24mrsw0DyMqGUspilVttW46g1Qkw7EYzXnPRBUUeV7sHPLCiqIQE6vfqI
/du1shHAPUuYFVggf8liZ6jn0umHLdYlxlNc3al/mhXHUCGnM1NRTm4XYsUXaDu+
T9ynBI2VnXSiQ1C5P0LHgz8IzPOYDjvenoryrpEEpoUK6+e7XDXpSCS7xvRS5it2
ipk2iRlwf/R09oij/9EyGOsPsVNYNvs3XEJ99UxAiWqSepz6MO256zzkwqd+xt71
wU4OJ+WFSZgV0lunPZig1wk7MUJxA8lRWgDl4oN1Stwt+yzcRxPRqlTsyGzu8u0Y
EleakYkv6EUYQGvxArerDKKeJcwd6QeOy55vyDMFoFesr6Nd2FK1e1+xSik1EQjJ
vVL5TbndoffCi+laI66Fs0swa/Xgoid1XlPn81IhfE8dbJcLUgZxqmNmqp+Lexw3
DYncxf3sJtQ+npfUnZ8cl9kDEIKJlEI/HiJqvVuISEMux8sX2nvXOwiL1e7sdtjB
0m9JmnmAJPGH2gSUefQgisW12eQA9G6G4qvutVl3uE5CVjwa+aX9/g/8dDtWnUOK
Ob1eOswU+SmTXJc+s5JDss2ehAKMiFYwP7a/m41r/vKL2l27v0RUOiyYMO7Oo60i
/Qq9O6LYC7DbJtUVAkIhKIS0K+Pu6KRyvXPGTEREn3339rGJgSLt++lnIpEkmN1g
SA/CXMGLo5XWl5Grhq5UshadytDu0qTY4zrlyVnKZkxAd/puJdXHf6Mck8J6qeFX
Z+s6pCqbWXRop3BKPUuEWUTuJP8RyzlxOmzYjQKcGZyOEH3hjv+YaDsKUP/9XyvT
iF/+Dxjvt3tRjf+e3KuBJsSqCPXcppyPM5nqwfDTLgt1As/UUCN2TaqIP8d5ljJ4
Lti6XIlzqhFnSEaSpgydkXhqQqLR9PAgOKHU/c2mMf8cUswRgOCsQchuvhUcn3m+
hqxSxu7On7NF0hLGteOYSohGucGkEOjHkDrAhkd0OwK2oqSyOrxq/btubWmIIxxg
fANGbWo5JodfsoWLjBAak7WzqsWW1X1uguIwthzIqcPb22s//9x6HK0opvQo0lqP
pqxJ68VISTFjJrp1K1pkqbE0pc9bwDJvkyt1MqUPSkH8EJUYZ/X+neVl/yuj9d55
MwIhqYGmaqi86pyt/+xiHHVNbYPK/Yaa8PPipqtHEp05sRi4LusJWxyk4OJJGlPO
AQAjUn03X75TgH8ycIMkttjmnvLgtF1hfzzoMTN1DUrdLUmU1oyOCbXSV5Bh4/u/
8ceTr14njjFajsUs7yYyg8BIwn3UHwh5qiU3IisroTml+tw76/dTZE2+IVidtZ/t
bMSghFqSyjnDk7MfDNFwQojKm2pSq750Y/70fFvvZZPZjSq9u4hewCSqaEfv8y25
009tSFJMfF+wIjriQvjvzhobj+E8EeHBeDmqH36XH9bhQ9mRbkoLf/2tLvbVXx3U
7PU31FFOduHH3pkpz+seuK/POID56TtQVqzP0Q7cmvxTCReYmQ6j8f9crMrTyErP
EAQI4L9nJ4U8e710rKvbSQcl3UkwdwyLpAvSyD9R2EVR+zVG+jRYZXF+g03BTkwV
P1sr+6TLzkYIAZL0nFTU51S1gRzh+1m2UCcr+hE+oBl7GudFVAQU83Ok/uZRM4Ln
Z9d8m7Kg2U8/AwHnSOKfJIOpvN2vMyFXltPCukUTdNTH4Z6fe2f3f94w3w/bfgdr
LURUGlV0WfhtaTxss6lfUowWDRaXyqYEWIyCX6oxPMjftzVieVrx9hWufqNDD/fZ
+ykQlvILpc9AGM00b+YL1wCzqOP5jUP8xTeAtXPdeVHjnHKly1VcF7EYrmiH1r4v
Wsd8LQ+cEwC90T7COUOLuJV0Vs8SaSOAfnkyMGy1YICWKc//hnW2DK8rYNt/2OqC
FboVtya78XBO5t1Wt+YTxC2G7TrV9vWfEyKuW6JPM57N9rFO5w3QcskiSyFTQbAl
TQeY90NOSxsl6gyPpTgzckaTdug0tnz24Ef+w90kYklZwuBLiR9uxfcBe+Gudy2q
ROpu0gygw7wKWBuk0FHVBnC7JO1uOEXhcJlN4KlwDnNU90DKYhC1UvfN9UMIzjg1
pb108pffqBY4Oa9piwCeLk6qVS+SC2Kl/cu5N4NashymLSeHNJjfJ7vvbBUYXK3R
vEFFgRCc3LlNIHPBz/9JzGn90VOLACIpl1FgmBL5JIk35MRoAWBa6c+mK3+jHZ/r
8p6pNOpZHJ6bFc/UCPEh064icnGL80bVr3LqxnTnOgUvPyHwSVqETy7wg4DU3JSR
88vVt5v3NTT1obXuS9WUOO0zhBckGP/VdGXRrefygQ1skpxcywjV2aDSydRLgAw9
z0nnHHENTRoidSynP+wgm0d9jbDt/d2XvXQ9SV1941wBPEiuc3pIkd8tXlZgBGG+
wvDRc0uu9MZnOXBek9Lc8B6W9xJ2b49Zdr4BFLMZZIaHxq3VwN0p0R/PX04QV1B+
DSBOBjT+rsR6jU925ooAashNVPOUgqtlUZn98Kte/TxJVNgj8ndITYg1MFBEYzqt
ojg3J+jBQllDhZDptqbtxXq9ZHGlsWch+Hcd2DXwHTk7OYNBXZZz+Q5ZwDsuz8yK
xuXd0YTa7CcfIV4AYoDmQDMS6j7e7w1dcGVJiyfjROLC3q28LARdOjPSOk6+Rk1/
DmpYInubUZqTyZ6AZ4UEFl3GFYXsaRw5L6xaMGejP7Wh5AwT3LFeHTvZG3vGF5zU
XQ5jDy0QG4KCZpIO5sqN6N9Tqb41wTPfbKGS9Or4ibqawterSVoXE8boggBSn5X6
kwL5eftlxjUPvoARPMC/Q5KYa8lC2DpLm7atI3uwwpMk0FjIXh1QbN5gKkhX4JqF
IetiQqArFxvwXbGH2CEiIN5i2L7W7hMgHy37FTked+y1VxEDB5HlliKXNqCC1pYv
Cko3GaWppILWCYX5ppaq1UmKFG24FtkARnZGE9MItB+MWrUjVFfEb28Pp1Zu25ah
m/16pg4tfnZVWa8p6GONfGALHyhckRPnaQ6zgPWWIFeUTTMWOJN7ytDXfE9flI/c
dh5mswbHs7htfTKD+SxLy+DSgpXZ8lm7zzR1TUy6l7Kjq2ccToYZNaTQWLJa+dwI
dvfSjuC5YuWtbTrE8XxswJtS6rLQ3tyyRgYQKMVtP7eVS0JAN20e8nkGtRVr0XuI
oG9gU6dDTwR9zTurpBNPNuuVNRuYPB3VBFG686qQ6+SehVQIT6hnwkGZo+U1JI2w
s83L26EE+BoyUZcOldo/mKtXpzL9OKGFbR5rOmKfdZLODNaOgWHHDSDvFtmBdTy0
9xWtEzUP1jhBGD+x0zbdQMzID4Nvpe55uP8CuO+yTmdnH0+OVYhgz+nZRWgeOC59
I9kBPk7kNVXw7c3glrc5ykPrKtd+iBavIoq4s2IB0VS0Cch+3/TBN1Y0OTuc2WWq
zwcw1N8F6SYCzEyIjPYAcccWy3e4OGSWDtzTREasx490wM5OYV/ol3YFeURB4Vee
7lc40aGd2fXFSUlWxkTPANAZxr3eJ9P53sGaiCr+LRsTMenJO4f/Imrf0Y+dOGQg
nlpwuArw429palCKxQ12N8I1qwd4V2xABogTNPOnYnI8AXaLlkvXr1FiBz40hn/a
E5kOKgoLna0CZ4OCbiAC5uDAM8xXX2hq8XOkNPamLquq6ED381yA1tacL25OrVB9
k74+t/HQSVxhXHTb3bVv2ez/SOeuFsl2T6yndTK/uyOVLGKxeXmAJ3arPAoRLdrY
lYUI6UTdSEBX2ImdTLs8ugjH+w/iBCr82MDiUGk7H5E98tceHRuOSOP16eCTHxrS
0LP0qsHx5xN/NxLjctsE+5GyL150mtaxWjGBhWfckFxCl71xChgRJMMgHuBmkOvu
Pr4GHZJAb/5FI9rwROUG5ppsfAxdYci8Gt+EMJQskoB/a1W0ngk2JforJRqJ91mJ
RXBucvoRrhfS4qE6Mvuatq1cVRGK/J3Jbq18vansoEcFgpVUw4QJj3FmNo8apNl4
K8sTVmHM5nT/+rd1WjTT6YBp5Svy53UQ05sHeFHFu4FotpAoReXi+6K4BSS5DSSV
10Lwho0hcOU7aF7UBGeskEwJ1Lm9tT+/cymKZsMeanaVrbuJl0/P/KIxyrv4n/EL
kLvl+F7aBg2elH7oLYwgJ4tSTTBQ3BHusjt164usyBHjnNTfkNKVOeZIhK1IG78V
Qo4YIC14lnIljqFymsrVMs/kmgJotE8sx1rzUry0VXVfDefcoKrly+jTNBPceYQU
7LNDwwuPENOVz2Kfrjh9vb8Bamud8RhlW0Jt5vWy5YiNRNMAKt/AyATKTVsrXVt5
fxL9sJiudoBS8zeo28Okxsows1k3xA9jcak78Gtynd9n2OtDGnl81251Iz2xwYWt
gPijYaDhct3/t+gRgQMBuDdjdhvaoUKzmmIZEjV4WZg5s6X1B9p+F+3S2i0M8Jzh
qiffHtIR27bk4GKUAM5JCx2Tzxqg/mr7LRfSP2lRc5qcgK/jRX6u+xnvVFd1Mfz1
rK1SN0b2X0VJKAsPnmtHPH8wYQn44qNcyyhYR+x8+rLaN48rHryPpPVdhk7kg9vA
3yCwAYKrH7hBmptozTkhfdf7bCt0FUMhk4IL6GnE7t9iC4isDGa63A2N5OAey8NI
V7cwxGNSzg1ORjYYMsB1VKykugO26B3rt4ujl7T5a5HliZG7afBXQIdHmbeba2j3
kIdUK5tzlBXZJP1mF/b8W69E+Ayi9tWONM8XIqzahG9dkRd0dv8NEYF58xngCDfE
IznMN+UYk8aW4O77EndTe7s8P7u+qs0q1MKGUTHRMIIKw9+Wfz0B4f9C6Mvxr1nI
/L6TJcH+eQODiKgss0dRwLntuUqC9cDlYqczxnLkFZFVmw8vKJLIbVawOH6ShQyQ
3k/oEk2gPkBJahpZRCBqeJnI8Dhp4/vOgwLzSUwnbaPyngVKm7n22v0HlUGKMThE
HyfTfbh38nkyunS/0kNeARjsHRzTsF4k8fBNTPWwDJTnPwgXM3xNlADSj/KkMG6O
dUDBgQhMtqvuCelHPjzYkqkoFwydWvIrSWQWr7lsqX9cdL0xV/MjO1r3WS5jPF1a
pGIEnsu07P8/W8iZaH8bHUO7ei38hPRtVN+qOwpPg9CSFW2EaOEC0nZi+fZ9qvt4
uUUXNxunvCtZT4YPavk2cV5oQLjvd8QbV16n3MAu/Q2R8i6UkLWjAQ8mFoS/HPeu
QznSpajBXbgyIS7kJ/BS5n+yZ38+ONNSd0OILXBKnYGCQigOSy5xLvmzsAwfbnYj
e8wyMhCUNTfpm3HfB8SnZ8+QJ0QwC8J6FHUhJkkIK286MOUb6CU1l07h1JNEhBsG
yHDWsLeUj2ViyHpHqjLHPsDYVTNH+wayL/4WhfdJxSGEaf8EaJEeL+f28cEkgHf/
KBrbJiThOKPdFNxhXtTGSU/zGcyS4z5Y4W0foE3k1iH60/OwNMKd50Yk1jxxThp2
Q/yZVe2udnZzWvzYKWcUEKfGVUrAf6nX5aBJwLOK+DxYZxdmb6r4279PzuWGSkae
jOQ7IG7fXHakB94GY843mtfSDdr+7EYBkTjd3kXg1NxBaim00azzxfN7c5h8zd2C
W8mAiv7VmB6pvck4swIUkdOef360vN7DCBwcI+IiXkgk3PLiUgBBhoLbzyoMojOI
ifHEG3Fozz4mOm3OTaWd4HlV0qYax71QO6z7Kdr1QjzY4hzRFPZIS+OFosJ/aZzg
YomEnAJpsxizxxPlPqGmqotieYS2MNHXSAjWN88gk6Vb29tc1tqKUWMgjfhiyNka
co77vg1okuesJ2UHUB5BuoQGgisj8Y/pE1Q7Tiwr02Faj9NkER0NH6OJJlnXBJtg
G3+NlG2rvBELUMSjaYhlXlKlx1g2jRe1hNMj8YT7pt6uEtQgWbUNkBWnvCZyHQhb
F83p9XXiJg1GCtuyX5VNRwgH/ubYfsua7vNgZB+g8YL6YIgXmcGufI9Q524fX/pk
ZuNHFjNa3eQzZvQQjYcvLDeOExtFMpI7zjZ63ssjHOaQDGDatG9JyX9i+YgHoCzw
diAzcoZn3la27G+Zyd9SryW2FDRFgb5/uULR0bETa1yqz4W4F6k8bVMZts/fLWO8
67iwmfFrb2Bvj1yVO09pPXps+5A/RCMD2G7/4OENoBJS6d9jHYC1Bpl9NRylw9qe
TYx7iTH+3WQGwRTRxpyF2vqnHJZiOupr/r8T2KDGwZo0SZHHS/CymlEBj3UW8FEV
UWXYRBgRId9ZX+8AGYDn7uG/xJAB0exgXaedBLKfz7Bc11MnplXumn0vLVUCaSH4
1Czj6zVVpQOi9Lej+FlysyRz6N6jC/uggiiZPXWN5RCl0c3s/Imz4Vuv7ZZKhfAZ
JvpOx/ft0nIiNl2ZaVW+ZD+BdIBcvhbM+xFi8Bzei15WycRyokn6jX1+nNrIjWJV
cGEg6aLOg2SSb82fiNin5EVXBVL+YDgiGiRUslDNN0WFRMl9BpW2HIUKCurk/mrv
mxNC5APN9azzJBRIzm57riiAU3CjirQon8DKWKnif0tOR2zdvH3MSeyyaXYYTXrl
IqshP8AAidu/m4GPEC3F8/tRNv0y0G52x3Kn3OqB57p9B1pcfuPAGwvXvXJshtZY
7jFSSWPY63OAOWQ3bgk/Vio2AJzYWvvlEw54AYe2NDWJEhvvZqXnMTUSS9ZIDUJw
+nrNhJKyGMuL3mQxKFzkoaRrOi5F2wytpdjfZ/qPIFdhXCWu9bvWRdJlljRKIRB+
HXUwtlNWgFpEH4stcsC32Ul3fl9QESGMsmkI4JH3NFC3T4q4SAKBkX94a7AB+lLu
lrEYahN4JJAYROBz10jChMk+ccTl4dE8n9hXeHFUXa21f+Ge0jR2FSzyRP55kZ9a
/ySXX4eR2wnhJDf5nDZz2MRhTsHpNFSUl74x9E37kP5/UDMOZKqt3g7xU8ARU16V
ls8FfvE7TYn21FnTdNN8h2U6YEaAwztsuDiU63wrEuOJbtPm25uhanQakGSQxJH9
4Fa+1+wRfgGWG9WX70WQSCqLX2R2jM/NOOsmjkLNoDeVInGr1OjteDKVnREC836K
772JJEF5LvRQ+B2iI8+xIBadwRS4i91Ke28WOhsMidMlYl0b1cHOklysxemxDHAk
t20IcAFCQT7UWlNK4BqK4UOPie1CX205iWOKHX69N74hWbMOHaYmm1xlItDi1HK3
rfpDZwzHOYtsFKel2P7ReuSW0ksmDOjwac3KbWGb9DrU7B7utveh9pkvSvHsRSbe
ZGGj2bwTTxHu4Ds8yljaca9K8P/NtR5ds41sATj7LQN5xBTvHEaHmqHCgpTljzsj
DYzjQv5qFHgAywouwoNJbYHyMqNSqoq9CMMxdFpOtL6XHKQaIMzqg9/r9MKM8rH7
Y30MSfWxavcDlO3w/oU3u4TI1QTJEms3xQA0ZoL6Kefd+clslBIbMlZzjCOEyeUY
+1AiyMART6JPe5T4UKYY6/Mzl+vZ9mCnqV3++QA3YTkvn2ZUj4i4k2eqgPgLTB4p
mp6Df/DJx7XE6QdfGokjVdtYmd8TYc9YC9eDQyw540dKkzhL5mPzrW+OQacCeL0a
BgolquBorf7V86jUOIUDm8aCTEbXBdekhfqimPiqu1hLSRhe1FK6SnlULwPnsUvx
ynMZZPsPhurJGHYqHXQZ/mPScwSnx8MuLvgI5X1KUG/Az60Ztlltk4iIo3NcN4q/
jOJxgb2bShSU5bMk4Q8vio11rqejvnZEd/qTSNPB0w5xWCWu5+SxwXe8gcLryyCi
9nPBE/hLAbtuXLCiy59Vy4JvpxYv8mWXo3K5zzShA33sKK0U1HWN3vNWl/yh6RFw
osaNdUiJpUBXTMvjZyvYGxN2poREFoxirMHXdpHG5nEj/7sMm9dK5VE2PevGdmc6
3/n8WjEn952bIXSjLtjzME9mkVDk4+CXZuFSlYwWnBIeqb8STrrFV2pORAwraZUt
R7f9NW5/EL+W9Kzkab/UMxws0nyhyFRhtIQj9DuyndLzLQ73Xt8xGt/hNvo2/8ML
H3zUgnW7Jp/yih355UW6tm4v8T19q/15/vNyThPbyqQD77JtlmaXetReXo9DYSA2
L6x8kqXHfKtzRa+4jfTlEJE89xRqCin0uJ5BVtSqGea3sGkjMHS9m+zKwe2sIMXK
7WGLt2RkiJ8wPuGlbZoKlFLfyteofS0JU3Bbp4f/k+eWRxKXzd24VnllWhYkUBKG
pwTAKzuBuiYyv6tVEuSKlgWALUbU1oL7SfBgsNuh5zuiAOgC8PHS4ffLcExzsobg
6/spwwUuor+FO1E6lakmPY91+ALuOWMtmxCnbH0Hm9RR2DnUMyGybqsDim/xsG6a
i9qLrOLwgfTgs1ytL7GYn4vyzGcFkObA8sj4AosQh7ms2OPU0hVtXa6glsTLMTiO
HqbH7ylEb03iP4HhXDM0jkZPtadXnerP4+SMbqqJni4eIXTYDyykAs4cKbl9QjeB
Zcpeg+JVsb3sOzPFaA3QQZnPdc8mebaG4ZkhWY6Y2Uax3gfrcHNmSTc+kAS4JH3g
ehbp1Kl0Ai2N3fz8Fegjp4JAzwzUMpiIZ9bCmmTNNwRjD23/NC92+lHXBVcEBNBu
wfsMT+UFvBA+TSKgkJqaGjxWq7I7N80YQBeRmoRsm7EHoQzpiZUxNnDF8goue9BG
VX4M0KrLL0S/eFkEJVXPFTrDEKr0f0d0lPGOiCeuPNeMlOAzaeMEJoKzeLMNs3Sm
CelS3YiuUuYcGcAwMG0HBf0/SAXi7TI7/2x75rMdsi9X2cXROwVvzlM+EmbdT+Bp
gZd1ixRLP3SbIEi2a8VVvj1eoaWSJuDgdaiDaQCapkLYcVxsizqoG+73jCabnI7w
vwFzvFggrRb8Ohwoi9UBQ2N83O2HTSzYMFN+MwN/l+lybplvo1E6wVe30bOx3TRd
mtBe4wQTgUqZJ+pGySUQHaTV97n3Oz4SWz9QPtNWP8zNRnVUgCfbpdqBQM5jMcp/
BnHzqcxpoDmZ5Y1J6CsAhh6kNNWwjCkL9ILe8m989qKEqYT0513RMGibSLxwk3gu
Df21FHJSL3aZXZcqrpc70OfTBp8QJfALTxVnxIQFRwJF/OCguUyQLrg9f0iuWDd+
h0p374LjVe/itvvY/YmXlCw/n1lRGCBmKM+StMKzRyYcmEcLtNMtjKxXkLtcoTo4
cOjkikk6yrutFmZUV1kxuH66Ev5QBOBd+vTGXzqSV9JqfStFq5jpDiP+2NUa2IBs
JtrCqkFoQejTbzqUd26sDSJb+H7t/mEibiMtJW87WFAIYsuaz6rH3gOmENVXBg20
HoJY+43qKpa2+v7aFlXe9xsCWpjhTrpOhlGDbYCHiX2uOOtovUBr4ChoX0EiEVtv
mOZJvC1WmamTxll0hI2sUZeO777f8neJ4vA/eJ2uQEU1mvfvMECxck400mR45ewZ
ma0uuwWaGHPbL7VoIyi/nQa0PHkKqC7VBv/kbZPMA5GfvEr4JYVuQUezxx2SHCNG
9NiN1B0cE7HNWNMlUQ8VrH9qRISy4ciAwolB4qbkHIpj59J19axyCaP+GO/CAl2u
mNdCOCc5KuQgj1bI0qamc+JouSVCH802YocSQXPOoFeLQRZSH0HUhd8tBvGWOXR2
xMPBYxrTXSnIr6t3GVDynV8sNgdCc/6ypoqw1XpgVFKdAfiFWAtFejy1mJ5karUj
xadJUXeiwtI3ycZ364WuKNvnNrQzSBC7D0wGia6sDasr+ERnFjOEKsJSxG4UWbVg
FxkogVw02j9qd+drtind6d7+weWwH6WpWwrf2ve3wBhODT7GOqV0KXKCjVgqrJ8s
tjLFQqIP/K6UuDwmX0g2Oo8NEgCw7NpEsrU8crDJ1AJh40y5MGUzy4vFVAtVYa0b
a1RRvFaDOyCVWaSKa+KpPD7VilcKQ3I8kL93snkXd3My7M0LicX/rsGwDt/rHGNZ
UJfGqtELjvnznfXOBen4pjwSveBOmRnPvO6bYvpSMuVYojsqRMHbmRhep/uxUZgG
5Ly1pQXl9KXowkgrfR1NNs+fdUj77yC2xIZezqJnmrtdvMshkr/fsVfWOHV3Ahwr
6rl12dRXRB+31ag8lWhFrXvCQJbdL0dDBdsu+YCK+wm4pYED5+I2034eBKDxiLbb
8SCZNTW23qP5jSDOpMTF2MRQ8a0NWXSYPL8zvvzOf2wfETcSfdoKqoYRXlrF69y3
7EqGXxuXw7KtfZ9rsKqmPromL3epY3ZQsI0UIF/NNbmMaW1mIa3qiL6TwwrapEoI
TbbW0+UxXqC2Yf9CW1dnlV/RI4eVbql6vXutcwveb0Ggg1oxU5DX6uAULV0E1hfv
0VTjAX7oLK8vvqga2qVzkDjyM6Dyy9qyiaRoLQEHYT0vweFe9+IKewtoI5O+Rf1C
ZTEynMTXzyO9Oyr/UvwKpUIQ5j55f9bEeD1AxpLjOVueVkWu+en8TCym5WU2nZ4F
z+cCZpFnoTPy+59ERbOyL8EVY4Sl8Uf/R21Znjv2uIkO1ZsmlNli+z+vGkV4K9sy
9VIiKTI94XwRldwlJEQuw4s8AifBp2+CeUJujH0JE8g88zlfinKjsZEMfxGFrWnv
FCBCrfWK+zR7tZWTVCsQZXRLNKlQgGPbekXhyDuaECC+8OcRjVMsp3mJESk+phGN
4bKwuutDvTdfb9CTxPDwHGMjetxoKmFYooRhCHBy2NQPVChwpHPQlMagNwzztddO
rb9Ttp77CTT4jerrZG1iiLa/7LDTsZYids3/s72DbM3Rl3gIx/SSpjNu4dvFCbF0
QJSY4pV5dtPuwFnPgr2W4ub8dMp5057iDxyZmT2kW3TE4vn8eJ3sfMXhwsSG0o1E
44zmtEx3LmTFkF96FdMXp8b/t/l4Tdr+wy98Qw3w7maYtRLjha3OZ8D0N5SE+zK+
LYwR3vuudVqHl5a66GYLGMY2nzO/9uHIJBd3V+BaAJGBN68sbjrCOxY6vxcU0B91
lYW2JpewggKJYz657oZ1JVFiENa1EIpmyFmDYDF2u1uZWhWWdy6hUks95X2+nZhI
BDIQ6pvInq5YoEg/gcFyU7AW+CpUKuk8RoG0StqPj07Hxta0dNSwZGD6FjQ91tBw
MlxGJHH4ncfhUOgMJJ/Xk1QwNmixdWeuryIqxfRmNn8RIO4oZhy8QdiIvx1/Cs/c
/VJSQTjCGgUlymRjQPiNqrpDohlFilgHLcfDhqIF9GtY3hKrZ9TnQIHF/ooID47b
qu3mjhh/Z1cz8m/RaHTly+ufAv4iHY3AGPmP8pOSeKUoUkQBOuCpUboF8QcjrDid
AgP+761IokdiNukNxKh6+SMS1dW7ixIPDaMRrtE/IxdAWd/9TC33x0euIvKUW/RH
wl+PeB2qb9lZ7MUGr4x0BAchzXI8jcpSdZnQGJqe4ts+giPYy3mDQrO+uIXnr5Mu
TqCMULd8dM855CuV7ESjtOwCcv4VP1/eQEbMKtyIkhtOTq45Ufo6zh7datBombEp
sSUY6sULKXjrmTves1fJi6/v5m2LwF/NiTLN8gp1ia9CrlLdHzoZjSww2Mc5mVMs
t7tE1yxO5wIRDft10unYAVh4bk43rNeKrpeGdHnN6ohExjZyxEaxdos5nBl2LNDr
o619LijLPCBq6oKdMbbsvMXAQaAoSpmLjzhc+cabTdelRGt2/T8fJ/1RkSWs+D2d
WaMsX5j1XPh/M6Xxzs71EvxphU/WGgkF+n4tYp/vYYlL9UG/CSAeJgkFBxo7xupX
2lFSJ1+cNV3aZK+W8erzlHINMeMT2nPn1AC6OMF58gXIXTpvlX97vzy+KBd7zky9
K6jtT5fOfW8cZN3Jt17+wQm3Vb5LPXzRTmBN9fi/kUUhx9oa9ROQNnt+uu8PKTlw
m2Xzyd4t+ORjmGk7OSRatplv99AqBRhtHdG0HobSjOj74BBFrlYzUd/fn6HY0P4J
2vlpRQQqth2je3NPL2vaLDuNqEJa6t0Z3o3k4yTog1x5qzTUzZslP6+QGUun/lF9
JKUhRNxRxWAZFwDTC4pIen7+WJvYRLgIEh9MoSwOWv8hPbDuEldpt+4GqjOwENbc
yB/h/oqV9YWZ8pxqSirCdnK9mvfABHvI6dfq8Q0D+qLL3u/1fLhK2cAhPLAWHHqo
+aKUXbjhbC6ycOylJ4Bv/w1fwpaRPA9fydHvwK+XcwynT6WKJkOAakwTqxHfaa8k
nKlWKO/jz7+U5xTl7wmMXgvw2yd2cnwuPZQDVgjZv7lQJNNAqbX0pI8Qi8Cit/yo
nDNQPjkxObyAuWWCCyHpW6TSz6kPH/QTsRrDiZFB6VAKVzItF9F85+nl5V3iEm/q
94vBR7ZD2PlXvHCw3e1y3HDyZVSGagHoUWpp+MIsDX1uvbLsMS/nJltT8bCkh2CE
d1EjpcOUZLfuAsW7DNtmzoKE1JpGZ8iTR42Qljjhuxlr94zTVpcspFKeNtQgE87I
Kx6Qs7KX6Nx5Zm4SKPB4EEDx53uCTxhieStxwjp1PVBUNYoF7v2YnUa8Xzh0nrTQ
rMeeY4p9SghD0MniOLuQ39iLiGBQUa5gR4kaSZFjwvM7QWyJkcx4/7QA2xrbuXo0
U8pTT6+cuep8wGWdX/+vycB6l7diAglQkw4ziw+dmrw0j5AUUBEtJysSLyO6L7/y
c3zWt1LTqKbNhfF+2bfdCYab6bBcLM1/FMQizcIzOG91gxqu3xujKcugIh9V7KVR
ovmr5ZpmBD6edDaewNm2njAn9UEX20gvs3uw1hl99gwz1G8rkNy3/tuFW2JUJ/BW
Tog8nm5WHCUMz52qu31arLUDF4mDbA36TY09lYPXgSkuryy4COqnh465ypvzCfz3
RXlrXLXz1PCmSeZK2T/scZEs04RNrcmhzjVAjCuo4miG/nCE9xu40LLnx7ejN76L
3MVfcAKRmoCwdg+NNYFCznQrcrm9X2odqzs5cGn5GgJx2Mm51pJtjPLA5wXgkqPJ
qH/bC951bJidWstuLD2nxflTK350Dgb38JTcSR7SsxijvO5FugDqnC8MUI5gBTgL
VzK2Qgbxyv4VRVyQK0L4H0/wn3v8vguDv38SYToKKLKrjEBADroFCyHKoKkf6BTk
v0JUtcBCHML4LpAKuvRiUAqC7/PpHIXzZLeYeteSgOzj1Q9FADnXKo5XVOqUc+Zg
ih9iLPnUwXcoJRbWSbiT9I9J+1QyK0ayjLYNjS1SEHDEfWL5ABaLG8RhgLdZ+k3a
448UkwqOty8vIKfgDi01PBOLiNvzdjCiababYdZWytdwsq8of9IWMc/1tBgZpTCk
+jhg1Nu8rstID/UmkC9mB09oNLC68Mv3VScSfWTT2fHyHs/4qJFz8OIgtDireeV2
vAb3byh1gnVJCRttYpYaseFfq8GddbsTksia/wOm6hM8MBIFJw53mVTC0f93HFv9
ylrfET+GGfUmBhWxtuUonu/iCcuUEP6U/dMBEQSTZrCUMbTE9OUUqG0wKPyDkXuY
WK7PlStxw2imxJsN2VT+mSlfbwVXhfqmjLRsf+wzV/xxe85T20agxl6GG7Uz6mZS
orkixHDwS/999hohT6a6tgetIAW14Nh1kRZmUdkUFur4OuxCiSCzto3hiPFmfl8E
p+NrLbMX7GVQcJOXWx0ZIljV2VktbK6eCiGdLR2c90sYQBTJyuYfHzkkKRNfbMC/
EjXUodvqnDm0fG9aoAjT876gYi5w0Gz6ezVTuEAS9NwvsD/JN73+pAg/C6Qm1GRv
omUXV+HLBQ1beMzHUOR/QeV9zga+QtgC1w+cAAmYTfvjTfWZ5jlkKlpQfuP0Z1Vy
oz6ttimIXpYBycRmva8oUkYxbRs57ozFVBNRH//Na5h1yqd75CZB1P80cSXNnmUx
f6p73uhfHIGTFlm679QKOGAdPm/CmcncIc7eq3mTDug2cBvpkeKKu0BOceoYJFSH
f3gemM65em2RLn/tfP8KDv+0yo8umM63PjFpIwHUM5XIqGJWh7I43k8GOqkJ23a0
7tcZR9hjeT5HCfusXVfrsD01mj18lXrUBsPxKTU8rjHqQsItEJRyPBoON5wPKWJ1
Oa+7DhTxiohtvHrcFf7MIt2xY+h8pU06stLdKW6Yt8uFe4uKXiLMVpdS9GE5AJLB
skZlU0AsCES8zQVwrvWjgGwFoBSdy0807FB7m0Aq1Ht7ayqorWDpavVAP8i9DaW5
6e1ghYew74qyWqIOgz2po3HeIo9wicoDT4wXy183SlEJ800vRtbfQWgHSsUsCmqK
OjggiEYe92wSRKrSAD+62hB+hR+HD04QjoukSnyM7xIo3BwyKGR3y4v23fc54KxK
tqYwCn/PM3ikqcHdjV4BagnQCZztDsz9LB+QB3ZQOOBYzBONYuGMjqPqFiWZGtCg
YO4EdlhTMO7Bne+xxHY+njHnfgLuxVr9FvJ+cOBgPDzN4LpU+DCs1S6bSKE0pk5T
vF2SYcWHhuRkoYWpXqvB3kYDofkWZciy7OKrnzD8ry3RWwnfk+J19kRLIRtjC1gu
Rr8SLTWb9vmaaKsRPJmNVEQtwwKTn1bl/LmEMYU0VwFHzeJUs4QDUSzVDxfJrjbl
f3U45cUBoRFqIBJV5K1Mq7+B60lS9VwOdayYvpWC60suK9kRdoK/XF060pQFHd2B
STsLrnkJ007y7IcMQEUmqWCYyi+CcG5EzlNxzaeEYbi/geV6/VZo6t34AV3Bvo7+
T0VL43TI4De0H+fA4UOt1wmXUjUGjQGV0SEKK3H6lIkVwWQfleFFjuTxlLKUF+y0
CS/JTG/d0bIHJoU7rmpwZEZiOQL2pfreKlkNjNPnPW0ERJ5cT0KQWv5D5AaxjgMI
9L9kqEeIsYybsPeDBtlXibJ2FeWOcr5eYbfIj45s8fIgzHHcoqCS26F7VL/CGS+7
BMBb/iWGOsDgrj7xBB8BximYvDHfsbMP5746bEJZjLpHABBM7GbB5iYplU5w0AJ6
TFl1l4vAuQ8kwFokrRlmgXXkh2pUzjIsAGc926pPwj88YUqhNRN4fak8Yx0nD4lx
UTWP1p4RZio60YBcAtE3Id7tVehowvB8h0nbmybLtmf5CaM8nm15g1gPKc+er61K
7ocoZtok8V0U/SSNXXyvvM6wY6OsPc8MB6x4lvAZKr2XLc6TnavmnPzjAjCI3s5d
bb/qSCA2UG+NVQHe2IKRsPxCUBooA2ZBfrc/ewqFwIVB0Qk3XSLK8g+REWuh7nHm
Al77ZrXZfz/HntgTJaTsuTfpN8SjsRc7xv8z4nikWlGSa2wrIMimvC901gCc6RYG
AvI9ASt0AgUgWa/QgoYH7pAi9KyuOoomK4Wnmff7zThRO2957Fn3XEEumAoQRnu4
XORNYjL6aX14h5z7bwci/y+KGHrPU5PckI07bymPPoAednklyPxHVOHXn/rc2UbD
QDCO8i3HW4Y3cQHBOlsVrU3nqP0fPNKUmGtxUU2wtkiEcks9yB29SPtiOK/t35Cg
J96MVpOkgXdc6+JxT9ZDBENaCoD2//1CJrzSo8q+k2FzkK8t5mW+VMljaqVm+gJh
uYTK+ZE+tv0WuaIzsblDr4UHA4gFA3pb0y8m7Vhd1qG/wlv5gMFSFATF1L/l2Hdj
2szBezFgm0eFZbSmgpoyYjcZIwgRIzMGmdCLZBna/T8hNyreJRePLfptI4nXQGOo
g+q+1UzK5MZUZM6B8uF8iQ3zU8wkPPKwm4lez1jvPfsudzeLX+ZnyaRX8wIJY03Z
BDFmgaQ60lGx1Gw2zBEBBWdc7JPRQyK1ZGzTJRGA+k4=
`protect END_PROTECTED
