`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uUCWKdIcdbjP8ehravZKcCTjx+GExX3MYEPjeD86/2oy/N0lvcK6XJBTI64WTHMM
PFb8Areg0NxIpF+goq596Q/h4tytYaHuXAUFa7KpNmyvzFWTPo5y/ukDaBkW3Hkt
jONM83B7Mb8soYxfcDr7bwT5Wa9yZX/oDxIxG7rlsnQqxe1ezGgZSE4akkoUoSHT
aSaG6vDih7tqujmPq42yDwf5EczsZQnIW05vnBB1xOappC5qO2swk7lLAwViYGWU
XRmPtt4LfiFRCOgTV6aH6TEmqA/ntqJf0fmCZKsFlXhTBzZ9q46HcccGwm+UVJKp
gyAA9fZKZOB66lngMeHN69hNdoAlmW5eBuGY0TGWiltOxHjBtztH7eLLgtIPCvZo
VpkN+IqLIND9MHj2qfZxM6uo82NIV3l3GBT9A4g+FNbF9SOOW9JcvsU+HNAHrLQm
wbda/kvE/ifWFiJzbjoaSl0RfKULiTeVY5LGZFS4+44=
`protect END_PROTECTED
