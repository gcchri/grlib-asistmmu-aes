`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XvtnxM/VuaSd3lF3rMYza8JOIOW9lGQ2+RhUHzrwPKFW6iJHo9kBLJVR4Cg3S28g
D696Z0KrBLlV/3WNa0soYDfFMX92oX5q7L1lSP7IBEuD3BelYsEO1IRGqh13Czd4
ILbyqGaTZDQGlzyVA+yhMt8tcYfB8rAyDno/oVUxZ5Rgi8pTzESz8vO/okqv+ZDl
QdKQ4tVHEIMTyrOecTKLc/7FkOd8zgdaN6r8cSKYIvwWiPk4nEqro+dMuz9sw+lj
8x4/FjD5+NfB6xcDfrySngnbV2QXBltaAtY7yg/VT813IwPf4ZEn2XW7ywoYXtxs
/d1USIgP5IuVmkdx52llOKDmPKT3dQsBSA1l0be/XftO3G0B/bExBZG25iZmxSO3
pIEskqapU2igzoBB7XPL1NreoA91AD6vNsB1HZFsFxsG9Pvzd4gIkNPmigcLKUnn
kNa3eMEtS/lrnQL8Zv7ZQw0G5y9lYEihIKEsIxHwh9cuuMGURdT0+WGGtlsznoiz
gLGiZDykupB5CJlit5SiPbcHjxCVqwyXXe5Nt3cjuV3PDEgD5kKKW3t/zDA6/q/0
bX2fx0h/SMuhmP//IDdSmbwz3zshMoBOe/M683uT33M=
`protect END_PROTECTED
