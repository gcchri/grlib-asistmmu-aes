`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rm1OGbZxmjyRPyYPwrIfPciJ8AP9ZwbcY1D3MDMYgnR6zgj6ZByi9PjMnfjZI1bd
anthAAAkSbeLpSRq4wfiLiZxcMRwtUsywcr7WwQKzGBiEjMltje/CYtLUKRbX0UF
uYdQn5aVhedIcqCz08rjgBpLy9VJr2wDCYRSAvp5qCwWqU8FeTqq5GnuS2tWebIu
xYsiL3mXEktzJPsh/g4TT+ab+aCv0JTt7+mbMyzighEPtqAEYTjihCs2OggPWmk+
5vkivjDtdTHiBdvexQguFIqKaNNLTI3dTr4rZpG8HfvbGb4v0PD7QF+F3zZu94Kk
152lYbJZ9NmfR4f1QsvbcA==
`protect END_PROTECTED
