`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ELho+pDF6gnNkEVaWivqjRSogaIxu6QFEtUY0/DXEPck8N8snGJfYcTDnW7E+v22
mtxBvSbVCaic78x+ResAbOHU2b/oRET8SyauGKWXVQjhfmh87BrE/mPpGbya95E+
plfC+K7sqVW4j0+2m7rw73fZM7UOhxGw3AFWV5PSZvCM0HJThVqfTnb0AkYjpHTI
ive1lyNcSphBI8dj+3hqp+L/gjx4bDXujOELrdgtA6D8SfCHItnosrCr+EbqXnNT
aXLUJ6Otrh1w0R4ahUMIVw==
`protect END_PROTECTED
