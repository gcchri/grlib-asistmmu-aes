`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9viQmvMwrVYW1tqnSLP/Fis2fbAh2M98Qu1W/j+ECzkI8xbhMpXmMbOZOfkm1XFd
FfW4zgFoT137zYO7A3nwHXIJE6I4nuE26tix7j00sYejg7ixx91x31aIy3XNMVrS
GChiR92/dPPx1KPMThaxDDXEWsJ9HMB7OPQH3eLLKoxRKGSXyO0r77XsfoHMdjr3
A49g2mbhOQ/bObuCPsJBVPk/jQ9BiAf7rWJav95wuINSOy9fZ/xz33U6itmHMIfM
AyoqUKpDn4JKi1Vs8lbV/eSkqf3wZzgetEn/gp62sA6/n7tP9T+Z1W7X9tjShrqc
TqPY4XsxCzC6ulebKnLbgCOzLxpDukdfifKPiUbz7f0pwnCcRLqBhLKq/c02kMoZ
9maPwzjyQMypJlqsGGSc5l3U1ADqcfV7cze4lnBQVbLOqIf1QlGDzImTe3r7yixd
fJLEl7ioDblLqnNpQyHxRX6V3BjGisUxK8SCtC8hNla+63xnMGgpB+UWBykOc3Vs
uK8CCJU3GrY51lmvNArfoZP7apGF+/2N/v3biNbv2ReuYJMN+ODefPe5pdW5mpyJ
ve2EAfb0lKKViZyRxd9+G5ct/+GqfAAikopr3v3nsKWl3AFj/GtKpghAVrQruJ45
s2M60lQcs7fTwJlmYH7voa3SsSgfScDYjzbgUMpisEf4YOVsNrnsXYTY3XlQm9O+
`protect END_PROTECTED
