`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yozuUaxQ4AmaCn/WkCj6Vvb8mpYN8udRoBy9mCPM2HcTaU3Jh2KQIJM/RcClUhqT
KN7QY2SZOTq26z1LTOqAFHN/Ikju8tH8yto7YMD3+SuwqL4etCFebHneEMg9jVcy
v9eH2rIEiSF/AsIXOtD3M2662j6TInwmdwhXPb2YuJw5Xctqo3fUQsf7NvrCvZUT
W9bB/9JDQN6ddC903uRjV7LrBURtkvwao52aXo76nIjN0YjlmVmFPMKq96HJRrvE
b9YwMVhNuWYfd9/5B5xmZu1VMnZ3jDzbkyp0kOeyV28bZnOJQQxRGGopAUd1f5ee
UT1PM+C/g6ymGU2jQe+RBFd8Y+NCCZGc6snZwG6h9jJiNEJmoLn7FsmMc2KdPaGA
2vLdygpBTm+ChO/SlSZkCuBY+hlewS/YcJMY4blH7Jo=
`protect END_PROTECTED
