`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AA68cqSommKR38llmxDxTJWDrSJxCu5HgHH9oRgmxsQ0W1XbW2aNykNuyuSgY8vR
tFuXNwZV0RXyrqD1lCv4bh/AIro9Y/vQ0y+s7B72e5cQcOk8CGrAEOaASmdoI2QX
4BC2HzkdwcmOs9PBkTOsB3lcyt0MDF8NmfbzmHxASoqk5q0jgcMEB4ougfKHUv4F
7ZEHfkx0wxSTFdhfdFsCjqZ/hoa+Q+a2zU2f+BbKEoK1zrTF97Wgey+JZjijN+cq
J0y4wBvjlSXAySFsWgtboqxKVuaF91txWoNl9Q6WcpcYxgiHuZ7+bjY4SgiEj0OT
FT3i9xz9t0dlwsq1k37Nu9l2VEVfcE4v9yl2ZMl6fuc=
`protect END_PROTECTED
