`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6L+nmlYt3rGn5EosXylDsqlnUe9YtxsrtzfitkFTp4nzIeZsHCMEE4DGQunfCMH
4bN0YsCkC8gpee+mcm7vpko8B3OJH+O9jmuc4TDyF/aRJFNY14O09jgmGDTUCUMP
ESUBBnL07vctf0x3qM21viyJEGY2/TTcT9mpf99vCgF7eqSb+iVZMh6QjCvs3o3Z
5pvDnXliXcL6bbrFJBqdG23Wl/E37lO6P22w4sd6cnOT+Xf8VF+MJbE5mFKDx34B
8pMGdWEiBNyK8IJl+pF6qiiG9eD6jl+WBfKx/NNyaIN5dd6lS3tXonn5SKB6iu79
fQVUE5u9Q63r89dZw53xtIXVNhSF+uY4D+VkS8Eu5pUBdfF1rkddtCFwa4QMVCvk
mhumIAjn6MLaFFdq/AL9J79YIWiy8XTdBvde46vFT703NOeSqDDZxG2dRHJXt3sd
JzDyaFG+qVtJUEYJJO8Gq27bQkxRNhpvkyT5LOlyN6w=
`protect END_PROTECTED
