`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YaTXnvkJdnYXJN/RUwMXIbh3CSvWDiYmg4Kjj4Nl2crxAjQh2uvBxKC0+9LChvw/
nDfG3moAOaoXuWcBa6U+ikYSagn4R8I4q0RV4tf+ZSuvLObREJ4neQ1kRO1f18Gi
dUA4sCgN0rgz61LmZJNRYehhbAzlpOC99zeMVUcLkpb+JHPAYmkEORvZGl2q88Ac
1O1gNTiMN4NZ3XH0kig+gbLa+mDFr+3AOOlSufYO9I6nzeHU5G/wxS2adkG/hbUq
cYBo97QUwEzZqefDoOetKBCoC9ld6tfHHV05rtb1objXVM9kAvoV3Sghn7HKKX5f
8dU8vqWtKe1rwfE5L9CXOxFj5theW3EVbejO4Cv1YBDZuDq//DuMf93JMvY7S9MV
VikOsR8zHIi/pUdiqRyWPCI34vZOzG1d/iRsxKc6fKkYV1yFL1kjF7Hbvid1zJvJ
SheVXvMVb+L8Uym2Nke/aV4FbnGamYnKBQI5muKSNe8UnMuEJU94JA1eqi8D/wQs
68nMHJeKi24sN5IBMcmF/UONc0GRcukxwONf/B9rgvIO02tTgqZ5s/ETMqDS6uq3
qrZ1UQf924t+Eg3othP9vw==
`protect END_PROTECTED
