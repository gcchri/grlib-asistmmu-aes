`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c5Cpg0Qwxs8kiVL60F/rHB0sZUbMbZ7CfvRbE/VsNPvp9HN3TbyoeIXea9CJ44yd
WGo0NvfG1l9HMTC16w+BHdeqXSp8j8QoUqGnEvVhE3D59/ZtoNyArTz3n6LoubK4
WZotXe0N9JPKJ4LtYCqAk5NpnevXkQKc2WaL9mpMLmDMQdFRhIm5XdNJtyhhIdLP
FplFcXq9GuCM0JjQB+4U33/sh0DCBq6x6hdqaXo8UcJru531LbbwWUR8I54JWzKt
tQ7myR6SIZvTcFPDoHl5yw==
`protect END_PROTECTED
