`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlNlzA9aD96irzEfoNj5KzA2UUhXWkkfIfAY6vSEGrbpNWsP2uwrB/XEkh+azsC9
+qPbGkBHoKkplqe9gPFqaowIjj5Zi65fFK3OXROBUh2XrmJ8xsJ1WsyUjSczQSTX
gZ/BekkMaq5TPtFaKNCNQ9JIUOtdFv7dta2Zp6sP56w2pJ/pRMN3z3lQ9GQiq/wI
WdO+NdGU5uJZOrtMl7/AKrx1v1jCAqUklf/xTdpfokFrIX99hxcVq4mDV8bp4OUG
JDolXJ5t50KAyvTOAw/T/Fz2XbvMZoBLZ59RG2ne0sjo8iurM15KQSJy12QyRoGG
P+GRgeyKO7i1s2LoARj2PPRQXfKzgdyfqe+vnvkkDkTywNKQra9DqOCmVfbo+wTw
zPa3TOJfgPP67Cx0fX1lWi3r7OsnQDE9vCPPgT32CJyiQEr24Kn4W+JGyH0jBj8K
40K9iN1O5VQFo1S2YXVrdlt8SOMeSokDNo6HiiRXYHsP8Z9Y4srurawURapds+Ua
0Yni7mcjeSbspd7G8DOYSTYDO9V2rBSSXXibmJ/Yjb7tngilHbTGmf5i9uo8pjfE
7XQEhtP4BcKjVYhTk7fvT8rRvUER/YedRYBJgaSqIuvCiX2AUghzDpBvtMmaVSCn
376vMEVda3UPYo46OflJKzVGKoksFgsMcfyuYmbFWSKV89sb0tHm4x5gUN5jkJVm
60MIET2fZUOTwuEQ2r78CLHMbWaUKry04OfphdcoFszv3LmZYLRJTpxawQCBrV03
DNpRiGI1ZvEnqjEeJWcvmfwcD/dgXyVjW87gdfsh0VOCc5F3SzoOh+ZRLihCb4Jt
LSACS/HzjX62MT3APe8X1gR+ttOJrAP3YL23S/FJOdXCvJ72m9Bvb09aTCg65ovv
T9se15aCn4IRAhw11fk+zRifW7yrtEvtxwll/963CCUMcuQp3oTEsBcgC3D60vAB
6rOmgAcNBrB6Wal32o+1VZGC1OXhU7NOXdctzk05tVteYrSemufnpJMf2zEiOBUG
VtpuT8+DmZYMoKM1onKammgY701IGCB4E0e/ITZz7STOGfPfEzrYuLyl8pcTw/Lc
Ry++RMqT53LL3xPnacmRMXOPO65Lo5LUAHHb7ok/ZWBcfNrxEipbQW7p+mkEIbpU
9xNBfm1s+yXZ14BEMEmA5C+vbvefIjC3O/80tgX5aun5Z6S1vRpsl5uUEWJQFBeb
jEtWTs9aEEuTSKrIN4f38auhSDDmmu9ZhhyvhmoMPKT8E7CY8fgNO3oR2QiGAXUp
gP1vGMRKLYbkbrAHbBdrsjNdNyKCkOSn+tJtK0Vu04WwU0nofBcA9NyV3eKknbWV
qmwGT1zha2MLF85702wZm4cHCb1cI6RoGytiu4l4NWnu1Mqg/gneLcCkZj6vBN53
2SrIAHp1oOpzI//7TWch8GR/vl7HLTw8oe5d7Tt7dSG1fcKetmFoUJs2KTFB3mvZ
DqeJMb/1/pP43cwX6dMO4LccICv1Y7vhRfex3h+RmO6XOJZmEODPd9uHyAuoaZJi
tMxp1OWX2PFdeuqWb0ArGQDeDIc+hrR0xifmsrsTErSwgR2PXeRVE96LVrrVYNVB
1yP5HtK1if1q4bhlMUnHWt5aO/qonecFXWaQgqdq+Y05o4UgYVodJD0qtyMIG88H
eSQ9LU4zi9gPwaLIdByC3FQApraKyEazNd+/c8H559HH2Mxeci01K2Eznwgy7VVl
V/41DvwjIRwo2GauU8VYOTvuY0QgWvYwrExhg4prmbeuxS41Q1KvPVrHDiCyk2i0
ElhfElg19Ud3tQcxpCaJkSN0x3LorwK0oOa4afBFF9kwCJySk3h1EP2arfxoODPv
nm5gYJJjGT0YxQ7V52jyIu0sMj16O1xgUmKLzTl+Kjb20gyrSR47JBqydqz42eVO
AbHxisNkA/13u1/FwndvpQQd+kRrE3Zg9+a8x53KiO/NVp6XwdiynBv6g4o+ELR4
LzfRtzEQ+zFi3l+XaTvlKP291rIbAdLIYh/dMy3uqXQ3qKcdo45LYEAx7ym1owFM
PcZtg+YUReqvI3U8rboNUnZKm4xb0bvsanvNucAcvnX0dUGihn6gjtSHkJ9sWmdo
P1ALS2SP0swI1j9d3nLi1XPqLJWhCgKMxYMNgk4Q/HnNJIn7seNs7WsF5mV52eSK
hPQPTDMa4bEqIslRm64OKnHs1QrN6h75FBfci9RMtLSfdJdMufpOHP+YpqwPej1Y
tY8RgTnwotWifjMRF4PqulyeZHlrRFyEcumU3wwhn9+eiV86SlkRqYic0MB5JwVk
PSGV7a2YLVq+veZ9QuVMt0qb4ueLAyI3QK9cbAZI35FhlcQcHGD05h7ZQh40C3N5
J3Ag64NrZfKf24WbfFG9OwBK+VnMJOZgBaxKtQaQ/5WgCg5rivkwQcWbHri6ztyL
nMogQPP3zhpkqyI/pzNETPTwcQPoN2uhYt9xeWlJfSfrE9xoRQWs6ZAwhULRscIU
s/bfRJGbHGJJpT00ztGZ6LbN37whT+vwY+iqOP2iW7VOhDA4SLL349n+z85tex0h
ibI/eoimvmAoPbxxefBDkr2Y2dw5fZiaDkIuSDsOmQD7o5jKtF8iu156bPl0GWw+
Zxuy951Bicoz3SOTQO8BqhDA3Alg9Dv8kaOiK1whRhrHJAXgN3VAwnweq74BAXzs
B5r8zhSNQTrtwpGeQ4Q3yg==
`protect END_PROTECTED
