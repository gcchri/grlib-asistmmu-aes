`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbOxv8j8ajI/RLCOw45uqTWDSrvGqtkjEY7yGn1l3QNYlEiebIG0ZHpekO4fMKQe
lxTYLylSeVl6UdM8eosVI1y2tqMf/zK6P4WLH1sh0bYm4PupQaKRXqxMck+H83Er
NsdMtzIkkhATNxfDuSIDpSTj/GpcBkTInbzdScmx44I9BF7L3V2g4EzyevInh/rT
Xp7NmUwW30XO6Cu8SzvsU+ljykMVj4Gbd3giupFbqUdbJCpLptWi5ds7UYo3Wok3
vFlUSQ2bPWmT/UbIYXmU016YUeHTRP6gV3VupWYIlLk=
`protect END_PROTECTED
