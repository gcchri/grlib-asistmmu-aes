`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rjvrl4aYB6FnaTilLzRL/Z8tORyV/nzdPPLrEBzLOD8RKuQdzsh6qwk0rLH24ZX1
t1R9DMynlvge871ExmKMw52m6Ij8h4FDOhfZh/1z+yHnc0r6q8bO7FbkcaJxs5aW
W1CslAl/36kDoALgJrsb5eD5l0sGAHE/nAHlurb6lztJ/B5S/Pzi0Tujl7jluu1l
uqRuj2bUZU20tcS/xQJRsEBHXolT7tjxR/YmSo6AFVlHZWS9nZDTSxso7Szc9UZD
9+FC0B7OOqH+eSi3NxmE1QLEqTbLc4rXhg3lTbkLcvLwObFzmtm5C6feho0ayDz2
DBzWEo32YMAQDIQlP/qtUyQdZxwZcTzCQRxXG1y2BFaCOQRpZcvFvIma6qIAjo1X
IdsdAskgtTH+qRpwDpSBgOuM778GboQ15kZTv4cLS4LPusUAcnFX+g1Aob17MOV/
TEvZ9WcO4PQB3otdVEAI//tiMKrQEyp/yQV7lOz4/KLsxjL+eGc30KOfqRIjrxOY
sPPbbMm69cgDJOX6UBksKLOhRQzmtrQpONIFbucDFTMaobAE8cG3ADElJHgkF/Yp
4E9dpnueAFY/5d518FYd0SfNB0xObaynKm9v17CX8oJV2vWlMvJOgTy0z9Tvl3Pn
NiCjfvBRhR+ptGPiNeHKVNZm1YUxJHgRC5qJoF43ouzYDPVoMzm1Xgmq31s528Wc
vaM8tWINVoK7ptcdFIQGxpkCP0DLYwRJl8IKf98fx8YbKCrLUpL9mRNwZEhNrSBN
yPHs+Jaawh53LuDPQdGbU/aLID5qItxPCz2x7evNy1SnEWiFntCy1U3s1Y5VSN2B
PtPwyJYQrWlnnr1FndXV7LKnLRddfrVpH67mfXk2Y6NKT04JrXUFMXfiw3oW4pir
6LjJDeCNxq7fN7jpixowuSQ/moyHMlBBLkfNUeIJiIWHNmZY/S1V1NR0w62QgfS1
d8K82dJLyYhw848+wztmm4ZVTXLPCPQsaD960IqVqhFoBXZv/vlxfonqmDJuC+kG
u14XOpA+S6GoYh4hq8t8CVbTfuCgbFUcD5EQ33R1ez0HqdU9nSa0Ku9jz3JdUvE5
cSfZ5X/y/oAvzHNQpFJZDyjYaBs4f8QiEvfhomAfRtURHztCaGwCyQDMHV+hvau1
qDyj0qp/vcXVeKaZGIPGejSJzbul10QtRI0AxDIbON/Gm27Y+AR7ahJiooaL+hdz
dBkcdZ1zVUcQadi3Xk9VksQrNXWobDbqHn//9alS6BNnqRJVjg8n4W+Ge7yAOwl4
9HpqKRK6gsbgt58QPBphqz46AhujQ2F0qgWk7KqpxxZW49Fc6RxmKK0dsTQJkhBE
vju6rxaVOp4G7MkexFeIp6KoxJJecrxsCzZsyCnrFOh1RvmXYB0SVhHRHw0JAGAg
TF6F2eFuSR0JX+eCUMbp8CjygKM4aYY0tUI5paj6Fe7WQxlAsG/hN4IZs56dR/fV
pikhS23d0R+zIcKK6ufmFxIMZFcG2Axio5+7tyDOQbxQX4pJqfE7cNh2OKTBPxOU
Aiw1nqOnw97WMIq6mFcfOpJtsTVxs2wmORAejEt4CU1XIlPnHZQ64+LobidERp7h
2emCtlscmnOEOL6AUQ1i1RJyzPZvD7II1eYThbg80WnAT9UgC2AfWQpduVcexAaC
gGj7rGI9Aq0JFjN+5B6D/bTaWHio9oVUDWoFlg+cASdBLSUZadx8sPmU0rMn+TTo
6S58ZN1ZOhM3H36EEplA6cQldU/yNdWnjvNQKWN2OE7UWSC8AUuVxj2NdRx6QWLI
FC8TAg5AeJlCWZZ3Yx5bplgtNI1askKcoTdpx3wQFlbwl8+Obx+jATfW+uGAR4X/
cFbIJR6bGj9XPLxn28xbgu8nZYN2DyhCw7x2McuS8nw=
`protect END_PROTECTED
