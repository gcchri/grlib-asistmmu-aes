`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IuYEDbiAFof4FrS5LFUqzyuidSrQbWvMfJXWmJ0Qk6c8SOBRzLljui498vstdnsO
hp/FoSY3DfusfBUEXs6io0GwlkCB0v/WcKz9gaPiG5CAy9CJ3m9qJAAyjTlpv6LD
DLk6A/XAGMpVutxHhV0RaVNA249IIjIngxx7/pN5wALVfFlabDcqofuatIFdvE9H
dTM/BtwvmGqWDt5DlpYJ/byrgOcNIfsPLlDgNPlZpuq9SQnaC/7rKXkPQbFxcxGe
kQwtfEggYIiveghJ/ai8eF8y7CBsnnZEtUEorOUddkoHQrQAf+zFA4teBvhoYjmU
f1z3pM2dQuE+9VhzZVQAK1q0eOBDRe4/JDSaceNr/fa7RVQug9rQ5E2a6aXHJgKO
fvhLTvpeZFwWSJExVhurhIFpDPxhikDX5sLDc0RxAoZVFgtwbJCT9v1tiDwUnygH
4RJT7SI0MKyf6rv7hdD0A1c3+sWVyztwsmSEQrjLJHM=
`protect END_PROTECTED
