`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zpVp0T1ZRL0Q0k7yueusFQK51JkGzH2fEDw+S03cgdD1yqCNtt+ypjR3fjuPm01S
e4pC9lDZ0e1EJP0LzslT9oG9TLenDQXp4q+NccoICSCdZbTddyYcJNMzpm02Zsk2
CRo3ARlANTCXJkP2TEptr3AEBFh+zyRuF+yriGmAEl+EPI6VpMsqVo0YbDTF+qNv
Ji8TjioLRo8OSnA/Ci2pGPep9hqti7xnNf+uOIWhdN1mKFBePjkZxOnHgmQs5xMg
JotH6YCMFpX9OdMwK0EnTXtJgL/Brm98q98j1L8jEEGhmRnilJgyg1CuzFi0PCDO
Z/7nUly/uxxQzMyV4nreKBhyIBibGWFAR4KJRdMvaLwwwnIjnnxWysxHLahTHCFi
e6OX2es1u7GUD/ZGx6pQZwiswEQbdb/EjTnJcxs5Kpw5PObzJWacIrDHPXwWqSsl
Fol5L0u9kn0O7+Iz0nXAQQeLsmHUlKsAh79PCSEnP+3cd7wYJE0rt6391oIkdNV6
nOOrvARJXWIwFelr/qjC8aAdUsDMQMAaMjfCp7MscVSBQ0nTe/4dd4RCRm5ayocX
4XD2A3bcx0AwlA5lFMRlbOxVburY6JrNeShr1Hty++2RYTbRnWBpNMvsyFPm5sCi
FQGCB5ttgvmaW8OEDVv4Myhzr9n/cK0jA8L8a4KZSC40OyqOi+j/EJYHUohD46H2
1P1X7XIZRSkV9lu3joS8KCQCf05W4hTL5FxmMpz++UoZRfhmYouRC1cSBAqpYaws
0APhUqRQ+klI2wNHhRPI4a4BG6dNotvkAL3jV+TvxYwNVOf90qu+siGJKrNlt8HC
TQN1nCNUbpj1dCwfBt29Spg0O8tUzOc/BTe/x4UTmpFhRXLBp6QrydvXKam3HMnM
6IOMIIyhafdAyfxhACJdvCQV6XtsFV35+FinFqx4/aZoOjiQPoDVg/XDm6cU6gFK
GW8Pj00LPenv8Y/MwnO/iSAaKkuHOHe04uUwf0h6K393zBu0CMooASuKTwdRvMpB
eum7NsJqDIlmspbT3wmCm8wLJLVguK7EMmodkiFWHFCbVNgwRlhFXyYPoOvPwLXm
CCflHfWNMkz5MYGU+IUHVahmQ+vFS6iis8blFEvZH/w/xvtUjNyZ78vyOds5TAYA
cQL0SwuXhVH2OzWWPKi+EaO9CUvU33fHyFUMJQOJuYr8vzWgGi4b1AaDgqoukpUX
emmNdXSrgzGQ7WhG1Aox1D9DyTmA9Z7DojK69u5T7e6Ux/N4BvqWspYFu/1lIkb9
`protect END_PROTECTED
