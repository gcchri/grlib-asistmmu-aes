`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6cAQnxayXCpYn3JoMHrMVsEpG9osY46CXnvXqOoiZWwl+mrkIy7n8amOyhrNmYll
N+cwo8pBa80N4hwUkpi8V4z7/TICv0amVKx37LB9Ec7q2dBek/rQcQ5BQMD07jTK
+8Z+0a/3PDmYjdQNf8tnoyjNDwDqjWpTfexn5umtnrXcqP0D2aUqDPdNPWaDzxXM
l+SMwWBKxSNfK6Ofdi1awbe3z65+/aJl5Oo8otHrLJRashObHaLUrPp91DhtwwE/
umqxrB5qJnBrpuG5TXRt8bPrE2KjHr8gMk9LBeuU9/3CB9EkOwr970GGWgTLk9r8
rnTr7khbAX7axA7MQ0dt39I+mGkZ1MbbVJnvdf78UXOPAragK3ovSG1Hn1af2kFi
zmQon8sEqdk2WVNJFPpnZYkSCKTgWy0h5Lbt8k4wCLBiGfxPtKnmJhUEoBKsHNOm
HU9DiO0+zJlddSwvqkaHfCzLWXvjvMVdoCJJEJTztF5iqjdB8+5uBeV+sRBGQDdO
aJoEFUKAfN6/axaQX9BjD8e63VQUXCWPbI4d+r6yNIj35gTaBwpz9QYXnjdIPeop
NcJY1LjjeVoxHH2vyv0xrOp1R218Q1/d6dhz12C131sffQw/yFEmyVXjjyUbvTQJ
VzgQu1hBO4dCcP8ZSH942DEcUeeprSt/67Staizkd1zYrGXKhUlbUUqaBUy33+qc
jX2YxG1B/E18vX4npqO4wf/g/9s7XfQN4R2vQyiFcKxC/nxXcB3z2TTx3J2gfxNo
kFIe2DHW8wH1esOQboWMhNAyyz8snWMACTlGy2mgXN/oZ8lrf7oUM9sAHHuhax6y
mc0x3hk36rfTiQqYcxcXCyiQ3AWij9kJKDnHJE3ZSbp2abJuwIb16bj2ez/0OV1y
1CAaTzA1WgljZT4ngbq/9CwzXlRMdM2hJ7x8jVSrdTxOZkV/PNUfS2zxvHQoBYQU
xIk6Y3sAUxvw1+/WBMcNh9Oe8Siggy9WsfGf/nTtIVOHgAhhfKGAexa2HInttyNM
Odcn8RfDlMgm82r7+AHjA84rp00XiIetu5R4vQ9+zOVaqziJBoR3HD+DkEwZye3+
22ea8wsoeBahNG78ufFfkg/9BXq95Abvs7w+PJ1iVsd/xJlY6ok88gE97YYRbIZ3
CjPm144AiILqAHiW9jJFOU2FYZZSKRPOH+tb5pyEtDdWylOqk//JDw41syP3ZC21
UPmbpp91z5osJQR1ce49rm5Nr+Nyw1sNOthboUmqAufiGn8jMBSPF+lvIBLZ6gxH
0vS/Q1/Bo85rP6ZS6UiZuelYsSchjpxcm2jr9SKk806X3o4Ft11QmtYWUmFSmXMG
3xb6SACC47SljZTYLNnjdxy22KhvHcsjq2qb6bEAjp4RNvwe0eHGgAEZtag/ggox
8batTR33B0ZEKOhCFdMSW8UskNsOlPjkhnxhB+5JRUufvfH7jYHJXufNkcJsBUhT
Tb+87UefbarRteA1nWQCh0VnhnOrIoo1r13dd3MLMs+GZMAZaM8IQd53F8n0OLrl
SXyKEXxlr7P/y+uXxF+3nVzBoaVyBamAk+p5/ZMfRwzj1x3jWvErq9DHbXmGCGZU
rKcEmQoRYIPmIVzXrYd4XZhHKPoT0aRtPSnwyEviKVXyidy19i8y8NYq0UD3yFV5
pe9fQDeHHmRlS+l9uowTttXKTpT01RKsHm9GhnU0hQ1EwY+qwHeF/NYzy9bSy9OH
pr0VM1EZP7MMSh8L2amcxWHJBlWNwBW3fILanYKepcrEQz23dlUtecQB76v89h8e
yBJT4RWqFtzackfe5Bi1bKz2G0lbj2YVCu5dGzU9YpHoEHRSRlVw8e0JUrRSByjv
mWUw3WCUdoiU+GtgTbr3eS5Y/QKOxi2bJsTHmKi2V9ipxy9358YszLAHdxngyGhi
beUNgh0D4c91xmFy1W6fNk5k8tKETytI4GZjID5Q6kaTaleEznxXLW9OUhwmMmDq
dPCwlkAMnjG2iYOeugbKsgyhd4o4g0tsWYUaXmmGwnLFT+jIRRfIYfOecTlRIDSN
nt6ppc4RkBH+Q+VVp40loXSzrUcL7l1QifZJoi6CYCg=
`protect END_PROTECTED
