`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltQ2V2G8BCYwi41akjL+WQL5Ja8Ip5jsG71QvQfnqZOqHTfb9iFaUeTXvcN4KI0D
hCI21gjmIjtmD8O0pUO9/wkgRIt9sWhKORg3LLwGPFVoPsL3xcv8iMHMEFxDJmwh
WHUWzoDGMhUv9AE4sq+/gy/H2RElpPD5iShRx7VZ16SaNuzxFVifyC2jx8SJb6OB
s+s+mgVEK3nA8PB3UXYQpHMNjYrSz7vxxhCkd9jdk6hpdKR2rDy9cgL93ZP1Srgb
gahT+BU/BVJcPHbq9MjKcSOvqciXmOIEaActwV/x51zRQdQnhllUmHECobI2zSV1
sG1VDn72Kp1CdGFxaTd5gzxSWVwOzsmDgYlH75TjNMuAugwQZpV/3mnxj+Xy0BQV
Pvq8T9xX6851ENuezp0h5Xz87mHJXNDe0ijR/J8EO19WK5D2hBvqR+06SkSKuAgP
YtCvuNf+VV1LThLanhp6UgXIXZMpa9tmRa3XtHOvNRLsfjU+/jHskrd2YP5+hSuU
hU3pAJ9cC9Kh/UKwJgsD3kAeGuImdC0u2+XcoibV7Jjlcry2/34nZOQXz8GojAnx
7o9zy72xB9Yb17TopVx+CuYg3/lwoZ4PQeWL2XgZtmitoTPW54A8eLUr8GcR7In0
htG1J5y8n7huXiS5WcdbGjbFuoBuS+UM3KvMP1wsvaORpT/Z+2HcLsLyBNy71Quy
W1uZEw9XXMoyrpAg39ZXdIku2rGVkUgeLGzzb2wK4nveYS8uvgjIL1cF4H3fEmIq
D6jbmm/lKtmVXKGghesOrw==
`protect END_PROTECTED
