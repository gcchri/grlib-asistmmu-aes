`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/XLkucb7zS3RwhFFwjObcFl2Lt03Gg0IqKGznPKhLeiI5mRWyWuVssaEFMiB60S
WlmvfqOB2eErp8Kz5A+szqGzRnzKnYGxb2XYDFEWstC4hEkhacsa0n4f1ecyzNwB
Tyho8UuxWplUjE3jDdv4hT4XC/SngH88xAEQ0HnjAPaQacUjRjQAwBwHbfNLd0wE
jmI/djgLejhReM30LgnvH1GhfjcWKcrc5X49d/wbuJ88hojC+ZmcmiL3Gg9l92H9
dv96Fo+KoVbnOvda1WeHH2Bbzt1p4i7rf2TsJKtnQkFypImOT1P6a+hTiHNjnJZA
/kV5uJM5rZb3dfPUotXyTzjeFDpOU8LCgI6LX8DOCiUZcUVr6M9qs7Y4OBwipMFt
9pIAsuwG+zMgXnGUasxJHvoHC7tFOk1uv3qTIXgkTLstWSgRExnuj1r3Y3kHa4sr
MLwlaosyRErp0I49XfkTqa79cBgcXjgyL+6Qyf8MV6tXxo74bd/rqwBepGsTyGEZ
vYZ/r/ZwshMKmTKgYCWa68C4cWnMjkpoPoKxqt1O/Yy9s7c8zM5XdLwdfR+E39HB
Rdivl6Xu3z+8ZkrqVVsVNx//zKURt+Xx1MBkoLfO0/7hRm3XTV+TeRQ6CFQjddX2
7J1IoHQSKBYinG6s2aG+e7zfncfbkCzF8CDIDes6Cf6CBH2Rdn0RQNAbliOWxpJB
Ia1KtP+bZDuuS5FS/1Y5lubY3gySWla6N8w1Je5ddem+A1mdGa9OxOnGbKA3YjZx
Zx6gkrXx42zqhGbQnLwcCfWDHH11aD2kvrVSYkkWM0qfyn2u7Hr5ZMW/Gj4eR/NV
pTmSlskDYtREB8c7oSvFrZjDdVpWY/5GTTqjroRn6CWnW+V4CNW+//V3r3M9+u+H
t+vmPk7zKByp4TLfu91qij6ojjH02XnoUSB2VwBMtG/vY3uuFXPb9SASSu3wqFD/
OD7ANY4RQVvrKcli7ak4/7dWoJnolUl9iQTl4kIeHhtzEYzZEJER3BuR9cW13mQc
f9e4Tfjg/oo+x2DwULXumSWLezJZUYiwVaAijp/qYOJpLS+egx2YGKIxgXVRt71r
z+gjaIcrcKEQNQvbglfaTJfdzNvm7sG0e/O7Q5WG4R+Pqm8dnpreku6PKaKwifh8
yN2GAmOVovFBAh3vYH+dW9i0ANuNNFPkT1dbBKlgGs1pPRNegET0lCjyZrPe5k5C
oPSYgBWgK5zWqKQ5m2CNjTSBRJUxD8985kzXDzl3ZvnBG6Mf87AUbveW5+Nm7Zc+
ibmptNIFLSlcutMXnXYvQE0gbnBU9qvQCi+MzzJuCCujLvFhv1emgA8s7f6qDiND
q5QSpID4J1AXMIYG0+BnBg4LY+c7/tEMUVhVWofRlvxXwwS2LX7MQev8+Rs5Z+PH
JLi56UuIruTymAtmcXT0xHZNfFging0xRU5p9kSR3cHo3MvMiPvRlhfLpLY7SWi8
ukGcuW/Sd6tAFerowBXBzVMcaGjuIyJh7ahbaeKbDCIO3Zb++4Uzy3RgKgN7ue7z
VWXB/irZjohMskQo4jdOxW00/toGuL1doGviXzFwhXhC4MyoXEL9+1x+B7ejVmTG
WKtQ/1Nad+diIJN2uoJ6h0azRR5VyrpvVx2hwlneWlYAU5jek/+onBVhMgHEmWBx
gUSKrr7bf4+UTkoyupSIZc7uBh4rz7Ek93xEurtjdiX6dDhFWbyV4J7xlx9MPpAt
vvOmAR4ntG7myTbqCCvAz0FUBQgElt4k4pO/nmRu+zQYua5uUThwJF1dVeEqc+AM
WJGqL+ir8LllaS0yhHFqJOHvBcE8W/piQZE5w0xsf6U0iZfKQJrqVyMWYysZ9Utm
8lVfu3lel2FSi6Si0/9vkIQ9USiiiwXRxefatCG18KL0yv1RvmDJ6Unzpj5VvhMx
mnNip1ZKLvmLuE7Od/aqJlY0iDNa7n1HzJEQJ9jm5JXAHA9GXFiriCbA6Jw8YjYY
Ap5lKcrrh09485CwtbfHnJQiUAEfREXMYXJ9NjKHK8/HRB0n07x0s3kCIld30TP2
/Ttls7MuKltxsf9WXbx/4wIqwkB/V1tmOVgDf6onHuZQr3l3oSI5gQqBJ9oJHpZU
a+k/HRr42AX8aH0JWjoLjxYn3a7LcUf0WXQPse804DnXgZLDGjy1uHqK4u4/gmpt
hM7gDVVPNNvS9PB1m/KLpQ==
`protect END_PROTECTED
