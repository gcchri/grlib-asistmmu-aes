`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DIuAyThXxQGEFWtdMpfghmEvXbFSIo5aNTP0SPDfEiU72veIA9WbHR/vabMj4ppS
lq3hiVMiLFBO6P4PzIHsTp4nJ3szWoVlNoHIL78JBRZZLrTxH3Cm3dUww0pWCq+d
Ay7HySxua67iBeHuWyT/qzoXSBOZ7Mf1xffg9GN9PrvDN466tyuieVTaJLq+MyD1
k7jRKyExZP715HVxtUesXDmVYDkTgMVEIDp28AV+XQ2fY8d0L5bWa+AFrWFEzwq2
o78YRUibLtW5ExCOiGZ4SkyYlGfNjWjFPakirf2/4ryEreiunplj3y/kiy8E8iyO
0BjJ71nDsl+UbkpknB/Pe/hF21s0L/n+ZZRWNLUyrccqeCrYvJZnaAKtS+GJecVQ
UShDSJFQOIIr7Bi+ygAgY+yqLptwyk0s5pgldiIPuZvSgNnArcf5x5fD2IWNkJ32
SK2A+QjMyj0rda3mdUgaVE9LdDmY0zSOJhpR+qdoJ2FMInn4Zoe+k+wz7zT3Sg8p
`protect END_PROTECTED
