`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QTKLZ2lnVl7G5Ag+y+gUngY3PVuJ27aBVgxDz1C/y/0KloUuIa0e0JZr5Gud96xN
REHc++q0erlDMQ83uMPlJ1+dsQ4KynlCpFz8uogGUawhX9po7cC1AyDCyBEfA3Qv
6Xc0NIp7BbM42jmJsySYMgIyguiFeUv9HsRqLJLAsLXnUodUPEZJiKJfcEgQsyDR
JpeCEvPkCQVPalycmRgQjU2nRpPDNFUTGIcO/THQEU6nfTbcStZD3XAT5oDTVYvw
IiepkBU0AJl7QvlnrAq2h9BLlBPkbYjAuG6aunyk6ty7mJfitVOjL075CQ+rw3OC
UcdVwjgKw8XojQXnp7tDGma+vzKU9iKINe66oXqWgryDOCLPDIFl1huHswVa8Up+
jDr8RCfEpLRVlduB1H7dLt6SgLFYrW02prLVjwUVxRWf9mbaEraSdggtLpe7IAwP
aULP1jiOHQYFQ/XI/q+G2Ld3tB8leOKUhtQC0fpWkczXkw/WH0c8xnVrbY/15imQ
HY5hFIufF/MTjV8lFw6ecDRI91zM99c70T3TXpEn3PKEBFZHP6djgoutcGhoEYg3
4xs7GwTWXgl2kPmNCEfIlDD1bn6arBcj1QMH+A/S5s8=
`protect END_PROTECTED
