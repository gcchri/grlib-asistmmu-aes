`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AEEU8P4DKL2+e/kl9j9pSrst0G2WuW/a70JZYsyH23F/T3PNUItTA+cJatlpQtf/
JuM+gjZAnPLDK+xS7Z9dds1RwlNITpy5/BdsWSNvrRliGtvAXTkgjQMPwLs6aQkt
XJe4j97m9bYBPiQpJrZAqBVG9xfz2G2+jMuJowM5i7JOkmq2vrVijeEGkVHCLipp
H/LMh55nwPATx6Y+gESGo7/yYLmvqpp+KfobHr6rI8mFV8UlKKrIZKqd+2A69r9I
qeywIqDP7OD6m3gI5LUkuCmWIhxVjgylkfV+Qi1NRBTmgX0aeP7lIpUd9uHi/OBx
LwwsC3M21HHzln6uCDru0tpREJBKC5gLSlkGjv9gCRmJ3jx43vVTETk0ffb/Uq4w
M2asnUtKfpiquwAJFFfaTCHaJXF6EPtdywUnpoYP5kGg5cJyNhHBTyFrks4eVdGX
CP+DWLl652MlRoG49WVhtZxyIMi3DuFYSKqqXUemkO7O29fws/fNElI77thFmJ3I
8swNxovgDF2R5zGQJJhvyVAa8jJvSxO0oUq6WiIRLnCtyR3y+cC1iBZ1N/r6JSrg
7rFMt5YcP99JzwdpNJI0SA==
`protect END_PROTECTED
