`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8LJ4HiNklm7cCPcccXM70JBH1Q9fuBe8zSht3j9lK17FqEYPBaWl251ZcpZsIMRC
HMwBxvvmMiVs2rUJrTccbgYIVyRajoUyOt3z9hhEDQz4bYKrYBp5J2oTXZ/+NIoW
BubD3pIX3ZhWqEdF3exprd+YaoxNzHuZnKsRb4mXSbDGcBrHmvlsxJqvLieIbDIo
hif3oqBcVA//cHwSKAW/yn9h9z85woGWYBbKtWH1eGOBz9+q2/PRRLq7gtRqcamF
LNzXZDgh6pZ1e792Gvvki4KFnrhcVJV5nAIpkjIll5YBiWBAWWsmBGOdDfADoHJn
8H0KEoLOGz4JYroLjGpSj6z/ZfD2aIZSBnae4e6oPiDc3hDtYBBVx3JSCt8Ib26F
CENY6FDoQTKd2XTGwAsPrnj99/mGoQ3mMIZseJ6SM2fCbU+Dfnc/3CvQ6ZG1pCb4
X9b/D6u/CjVk655rNINQ2p1Ss1ywur24QttDbiriqBGz4BuFdPkM9/fPK6qX7x4q
mbBGib8L07hZmmDioamxmJjnn5qAO34QQwH6B+F2cYaXYLH6VFH5F4kSDkT0i66j
XJqp5JbGn5N9KMGICciLJOQnaO1JQsZjDlTcp6NIMdc3yu7zYH6FwWnflW2SwhSH
`protect END_PROTECTED
