`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1t4noRcOLHsCFl980D3E0xz/gGfKKOdMmy3aHPGIT0Fx9hNZtrDqRgWyrNtKNdWS
IqMGFYX3HAGsEHMpCceHaZ9O3eSG+fcbWnDeWaV3668aAXJ8b4SFOys8A7DhsPLP
jK7s0B2xpPYOx2UP6JphvP20jemC1ZhJE5KcrE8eW6xYd5/aLSHS6uP1xrqMFtz/
cDd1UpxDqMxhqAWHfWt30uJFKYO+/bzdC1MypV2hw9rjv788S9KaJsmBvrnyOmm0
A7lexAtEVy8exexffxQw9ogL9gn1j0ABq5lfL5YUQB7tPLBvGQRttZToU5Ooly+n
yBDDfTQfSE+AKGYddFGf87sOcFAXxv+pyYoNqZBe5X6EI0DqpykFKBs19dgX5jIM
WLJ2rvYzuPj8gVxy9/xH2v++KznAXCE3Dv63WgmHyZZ1aLKm7LAsuLFw6vuDv1DQ
8s99LSzwka+syT89mAFFHeYuOU4t2Ia91xewl+Mq117hVsNEK3bJlRT8plH/Oj+o
ghESuv9/hezoC3DSjAajhAawUd9LHl/os25Zsdo93lAxvsObV93+tKUtTqobq6nl
LD8QZGSNsACyiuhimJ0RFqmlLPPFhCk5aI/W3S10Lt9oUsuMaaa/V4v7xBeQf4ol
7K4kQoEfmYCfrU0gRLTDRUFy4R5U7vOsKUih8Y1MYINvlyii6j9aQ+6gvVBrud2G
`protect END_PROTECTED
