`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jIHJEsCUNHuhMurfMsBJ9HbUDhwIRaSh8gYy0jBUgqpyTTdNTqeBTowWaKrlXL+h
qOJK3bLAVFPPgkM29VdFljEheMXNIqqTR3ybbsshocDVOHAD1DTYeNZkMvluUIj8
6E7Dre/Aiq6PRaExWDlVhlU9g6kt56cZjDQohYitVsJYX1EFOHGK1cXfj9kXIpTw
6hXAD94DzsVqCZOW/4WTPUk73KeGghDes9+GUX5YZVTv3QGqI185zSh/Eqo/ek7D
KsSAXunnf2u4TVZPwDX+UNMsz3FQ95NEATQp0TvKpFzGsxDRF7aNXeqCkmE0xgDh
h6s7za/un9t0do9dcv+Zqt9fNhF5kPtcG+jVG92Hjej4zv7AgCUoIarAZfaHmiJU
i52wFU5bS75DGn91vKYT+deZVoFgNx19Umax6Rg18ovRXLw/poy6+wus2Lopsi+5
/xVMM/BI+ggsj9mMp8n/caUskJwPhbsYjslvqu9bWJww0tGCczJiAAZp8cFmz9vj
RzlzBA4Ka2tIsMAAMmLM0qLXi/oTO1O/Pyn1+wox52khKYTIrW8xugInKPfjzCXS
YMvYRZdKquS3qCvrzjSfBVPAtaoHr7td7zGKiS0wvDrRchkBdEMDHkvdItGy8p2s
GQClYoEKJPthy5V/VsuV9A==
`protect END_PROTECTED
