`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4xWSKnA6lSvwu0g2Y11omfq8GZmCRj9PfJJzaTDEltGuT6JS6eUfM+u4GhWY+CF
zTqyk9Al8120i8Ff5JyoJ+NW9ZP2ZNtJhn0YMxj0yul5Sqrcq944nJHYZp2FhZo6
zhFWQDLEIwW0A7r19dnOv68IkUtcn27XNCDrepcPZKswtNC/GbKXcxNd36JuiMBL
n1Nz74EeC8rXuNlH7y9rcR5TaJCp+P53wwoO9aTr4Jyo4HUCCg8afEYZjqwCNU0P
mYWF+LiqNyFmlNSdlcsf0X5lTVK9NlxkNkilTr5/yaCDmWL1rk/Y38edTP9yOn+p
9o2P68hPgkkVNJbFHWj40REwzALFvjysndzBDKRiW8P8qkN1cZLzcMYrIQidHfl4
3O2vl2xowKrxC/lD2bmQI9Sv/xfi+G87Q/WJxv5dAxT2mil6QI+k5vcmHRpneZ7o
PcYRIMias0kuoX6w543IkshLA/MZ2oh9v1CZvnLz4KBbpeubPxtqqy1EmNrHy+lF
UIBn4S4Nqnuy0vsWv2BTmeCOiriEdgCvn5vxegQPoQ+9A1EWh08iX/HAdCWv2onX
JU+9bokR3KeLZ1zVE8p77QbYoRIsYBWAM9XtR+dDErkbNVNiS2JzSZ56+RvR2gpP
xrHk98OAzFGNUlxPm3ekZ6mihXYaAy8VacRhbLh2fBsd0uNYjWeehQYVdFRy1i8F
e00+VSjINP1UB/vwC8YKPpt+sZOMPT9+4JpOVIkyyrDwxPdjp62nOnTxd+Zz+chf
/vv1wmXFn8fj4CwkwmxQq1PEj4Tt5B9EEBgSnXjIzZSrxmjqtXWhcbXQXOWYMYTU
7vzxsgBfsr0vtS6FQEe5YVw1VfIveqXiHjFEUYMhBfyKq6e0UzlNsrn1mSx4lR1o
EMOd1mXnbgGT4hGce2qQeE5Bzzl94pO8IP5gMXUJWPGloULYycBO43hjEjAmXBlr
4jwnuN9rBVI1YVeoePljnvmFDcEtqcGNCBB3D2FHjVYg8u3/WnKJJYSmnD4qvt+q
QS134DehZ0HOPJwxMQ4kUAqKvQ0g1mTnQUofiEtJ0BvAKBEAKfdimAKzUDlL2uIQ
pOnW0RBJ9QhhuAUmzuRnNb9jxTT7zHbun4ys+mlrrdJxktdzws7VLupHl2qmuPAg
EJIpQuu+HhIO00Sf0sgbhwHZstaU41/q5yhKefTGD70DwBOYesXZ54QjKJ81kpu2
VKokifba6AT5TqceZTiZZvRlKt1cplEngyjucGqm/LjDt8bT0c40ZNLDhTyYLleg
LbZF1Z1dAx08DZYesoJo4/o3QJjlzV+KOGFDTx2W43lyjCAJgKbjzQheVKmVSTez
3V3s8rY5AMlNQFgEjwN4M0akNW4Bgu7GEe+DvTohU3aTf1ybHAvQpiems7jdKxtI
VJnbUJBDMpoNlykzAdw5UVQ8PIWyOHPUv/uUF/6WvSPNzFGY0XKWZhUniukbF9T1
HvKZj+zyQ64ic1bWqoGSLJeoByKsjed/A+BHz5oXs5Btu58MJEO+Vwl7fze0n0Qo
X72tO9HLhjxop3eZOQT5wp4FfKvz5nkazXEVBL5YlB3IApE0gleO/t86ZzzJyskU
goQCZcVAQfWmoru+eR0Lq+FSsAgMr9PKVghF5wUVRcHnxGCMBJ9Dn6OsJhQtfd8V
PTHIzxRpInYNADsWY4PcTbsFgbU9ZxEOvd2zG9qPCyM1WKmaJ5PG0jcnIpt7ZlEm
t9zjNHRYYoupj6RRJoo4DYpY9SXXGXh1ZwWmFtX1OdydTcYgrc0OtxqBu9gFnlHd
mXzAORUwu/tIlgiEORdbggcbYG7iBeLfCVcDS/l9at+gROTnF8y7CVD+QxeynXro
jAkw7XIpbkXeGy6Q+7qUJEYPN1CA3yO1iOpQzwx977YPjsH21m8Z6n9aOy/tx4li
dsyoknOKD9qAbOiP2bL9x5A53FGjfIUGg5QlpIA5Ll3DdR3nOqPrba3hG4fZrUKZ
bpZ9nE+BoAY9S6nZrpjO5TK1ioYI3V89ZrPr+eFn1zG7P1PSxxnejDIjPAeSF/Dd
nVs/c15gJcqMtivNhycvug==
`protect END_PROTECTED
