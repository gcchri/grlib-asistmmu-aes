`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WB493qSwk9qBQYomQzTusGA4xheylcoOmU3wEeRy1ZMw3nO6gcd8q4OFqaopi7nD
I9BWS6NOs/4FG18UHgWgVqxxXgPjcBWLfTun/4TDYvNfLKX6/SwCFqQDjZ8hlQeA
uq96hH8iv1tgWWisCPS4dTt6uqOKn/+aGxy82Sc/3zqkVQJ+yYlSoHCHzflBXZfc
wGD1/in9mEJGLtgJjjYgp75JjAJJH/VReJn836UWVulSr1YeO9ZN6hroY73dSWT1
X4nEVvDjgYmMLk0hMsXvG5RiKIXXKRp6jgTiMPU1+f2ym/Yj8ARy4imTSqnta7iy
Gcv4khQ806+BESB9Cv+oyZnMIUWmlgMVNT7w6nmy0wxjgcWMhSqx6yPCa5ciqauP
fHr1wNSEU9wYC3xio6AHODQ2Ks13tBFFfviKTvr6uGWCbTg8K0Be5xaINkSzH/7q
V4oOK/bn9nDlXgyc6E8eDZ+GvMc8qUBs80TCat9l8Jo1JJW9FgDowEt64tDVByCG
7t0iU1niWcd/W83MUfEk+1Vi0ZOY6/qDJUR269fH6RcFyNBuxtaL00ReIj2ynxME
J/mURQddqmPMXrr+lJrUT3hqHUktzlzz3E/y1s6tMwBJa2NdGtroghPINnwfUTOX
QAoOWNGhKm49DK0UyWzKv5SDU7tHkLWiewhaAaVazWDzz9fd6n9whtCn4sxgD8LT
SlFXUkVLakNK12Samyw9WayjzEoUeFtvv3jky6rtzTDbXYVe2H+nuzEYs689ISBP
V4dcWQMd2zBRxP27IOH0dkl6WTuJqaoCeoKvudS7TDe7YAr9mdK2CDYwUY/WPRJa
XMPI14OeDdNPGowvdYM2DbQScQ363jrlVYuhdpiVrheHViWq7FOapIJleGvBIR0x
IN3NFgPcctqq8F9NzUzPLun4cwCKob4t2pKAL8/FDRjpwSJq0DqNld+efzHWA6Yd
pIUfDvVYGMapCkdznyev1cxMcBZ6yLciVOdliGqSdcUveaWzR0B9d2PGJDMOlxki
G4+JQ0LuULGPV801EhJy3NpfzydHrYlAsn0YpqRWNKkDrow3M8Th3bOV2IxgnBnN
qnYp9QtcDvCe1/rUobMeN+mwFQ9FnJeEUPrCNIWvmBv3TK9RQFS/D/RNt0YiFvGN
VJVQHDchNNBDqYIb2rWSFBtTf/rhyeQ091OPSzxc1ayd96tQOI0hisSEXWs5mepJ
FAhZpPkNrESMBx2DjujFXPn879S/AdkhMTz4m7CPKnfswalYz52GVv6H2QoXLhAB
kZq9trwWSWNda9XDQT2HKMbGgQQhv81OuCUXkodJH+lto5oplYaqzLNsILTQxISz
Qo3QMOiAm2YjLALgnYLTnzHq21y+5CayrhN6O6wFylsBGQPenA7nCibW7VKQ46Sr
p/KDrSt6GFBXi7/nXtBzYu/jhyDHyXGKNi+LQm5ZHOrdNnC4tBhAjVRKbwpuPdEx
5O/m5TKV1rt8KB1v8LArxZOdrzkZG7WPPukutdtSaweVToYBfniHoB1LQeKG55u+
iyH4LecIzU2m3NdtSx/fgIROa3Ywz+/BXoasMEiz3z50H9cqV+8LlrmcPT6M7o9z
1XmiNWkvIRWIpHRH1nOgjK1pPmAyw+/V088twuowk8e5pWI/6GULupjmSKYp90Z6
vMDnQk4cYkNHNDi6o3KjXmmV5q/khPJaFqKcLvinLku7oDS5Gm4cLEPYU+wx2t2i
sthk5AuR7fWoAL5EnWud3Q==
`protect END_PROTECTED
