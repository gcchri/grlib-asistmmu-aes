`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0VUQv5eFAtezUpekxPHEKrsei7vw48x6iMOFrjUdFp4wjcTI46e0tfKHgkXBxw2S
1enGsqL6D7LV3eEPzjKDEvyIEYbkywLwT9kwP4HlMoxof3STJRxM3Goe/XPG8OpG
20kiRXHpFLwjUWJTWUo0nXPpv7To6NSvA98hSs68ZaZJg61hn5WC8hisuJrJ1s4z
kkxwnVGlg4v75bD5z5t7hY9YUUDFvO60zLKU9Um4Lhw4Yq8VpeT4JFqFdTG0isFM
Zmx9W1Ju+p8BnOqnEZdJHt5U06N1iRaQsUF0Wl3Mpz3rBBXWQPO3kE5Y/6a8lvtX
a32olg8Rksu44n0MyYhf6l+cj8bVtcqZ2iYYVx4Nxksnf1O8KNAEHjW4+0baOkas
RVZp7AbbVyZ1sVi+o+iJ9bDpsej8vz/+CqQSIkiP1OuaBzbsQchtjOk9ZjlB3486
HkW4xaeh0tbd83HqhkAMXwluvw/1SnTUMHNjBA46z6I=
`protect END_PROTECTED
