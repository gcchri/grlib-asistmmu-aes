`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ErXMK5e9eQLpF78XQQSIHEIsZXtS0wNnQfNW+fAoLpFBZV80rygjAl1bjZTdrOlJ
PfTtZhZtj+VxQlWxpNJGHpdEFkIiGi50CIAQSQTvc+6TH7XtjzoQzvw1suXtSiKQ
WADveK9Yzycu7L8CowGnur4XtHyR5sxZ6zlUaj28lTifb8NNy7uBbxK7c2VSa52K
l9AKv+p8aKF+/tjQFgjGc49rzeXcUl/qKYM15QzbELWV1n15bv3YLI+bAY6vAAzA
7H2vVGtFcvpmd1kxzMH3hw/f0zgtQv67DVLfGt/dUmk=
`protect END_PROTECTED
