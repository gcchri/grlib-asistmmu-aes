`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M78n2LjInDk9oe9ZWlsqeAYi728ZbE4U7NP7Rx9y/qsHVrL/kUQduVQjtfU3dsr0
wVtiYl9cVs9BOtXp8YLV+3YUPtGX+ZqXkA4+jidrvqH2tlQw0r8P1L42El30ldX7
CB8mhgrATYGb4PNM3YGXVfr9rl/FK7XEaEmiGMUAYdzqY1/kGd1XxcvJVlNxwNOu
9qoGMc2eCMQeamX/EIPuKE/fj1vrRgaLd9MV9I3MQj+JPzQNSbz09Gz6SLVnCYEc
2sL3nTfXR+y49Rfv1hX0/EQr/q6HxeD1CMHyJg/v+Z2nouysmmDlVUJ53RogOqvK
m9cQLpCpQUFgWfX2weMMyua8GDXquB5B4Mza2E683L+BFH3SVDGnTCmdVPwa2cYS
11QQgQ7XcBYuTs6VnGWmdEL0ox3tVZ2WsM9l33qqZLlcw7DENHb/ZOnTDhhPpghi
or6ubBkgX/0j/hD2Ikrt10nPxgY851xa3t7E3wZmgXUCItL4DwmViMEcguIXoADl
MYRfs49tTKw+gO8Kk/6STKx+hpjWFeddIBzmk7+jflmZEpYnIGzzXIxZx6fhaDXl
QrUxjcI6LzwOpVFi4aeqhRg2j1tGlgfUsAdbdRn81IXyuZS7PtsnZLNxEytfkKmB
zeVzWc2Jzte0FXgCwsg25Q==
`protect END_PROTECTED
