`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQk3+KII+hnyrLpDoGsYTAHVLtKzFHFIvLSfJWGiGEJ+3jyMS3YOKJFysrywLv56
ifhrEnwUbaTQUewHi4K5oVHSkDEYwoSkXj89cYzZEBWwct7fpbnqLA5FRcWpMXWP
VOh4gyLvSySRvDYv6zUaupkwPQPMw9NeQ1s9Bnc2OjD+5qmgG7IWxAqB0CgmzH5s
ZoryuFX0gOJE2j2A6bkMeNK0cY/9eZP7KVUM7OrkZrykrDnbT4uEH0yitP8JM3IR
ZUMSx7RDZiYs26nJ2V4oCQU+bA5ND1LPDZOSeUDBgMgZ2K0W+pfwDjxTGAbZZzab
h4EP7wK/spyprByZIRduMhHiVoamUjxtQdzzRm69esct8PAO9Re7f+x13VYv3eFQ
85xNbFvR1cEKfnux6L/klh1sn7ybA2fgA82epzIj1gIB2NjJzyEKQ1XlRJFozrxz
52ndS7x0gE3cWBVym+zJm+Xj0Gf8MDIUPtEGVZGQX7z2zQtW65d1Qk2gwZLdN64M
VbjVJfGJ+e2n3xa7k18/6kWIq57U5hvFBmpKPsRTFI/yYSU8KHJDjC5JB+FWeH2M
Ns37OTzbUJQ1Ad5SYRn4PcYslZ5R2R+fu6I/ynzO0EnM+7TMcbMxAYThQRC0ptoT
SgvUgeIFC188uZuVQuFbTWdqF22N1w+jIwhH8YPnOLIQ3kljE/qOcehwe+55Y93b
u+LhRLyAWvLhpVQ+U9aiWvVp5ix0iCauwDkt7K7AzkZX7kYRPu5wsdrlnk14E5yI
/jYh5RAHi0BxDY2cFCkixpkw1sdBbGTnlKvPNBJGp00QfV6QPr42+83+AjPh+qtE
Vn//Q3Upx/9Tko2dmUR/vlrKjwV5uxuzJssXEt540QXslUmfNgr4JJlJzM7O1EKf
7lzFFIcG7XbCOBi0aRcIS7mjbZKS7gdOsqNBarb71Y+XyvDlIh52QPRUeDG/p5gP
lxZcyZUScANcxb05Ij+FJ4I/NtGUeSnFbu6KEWNmzL4NoEbODwrU43//T9CAqXrF
cCtzLgt77aw5ryZ+0gp8To1aL/2x/vyU1k1p31SHD0wBuAVNzKtYYZjv7x8HmS7u
oW9ucK9yt3UW5kUog8GVOXfqIhNiDxZSs0doDjz7qobnGW9FGP07z1PeY6hu9bM/
efWPUkHCtHg2xGwwDdAdAfsorn9AjOHziZBbO1ou75Q=
`protect END_PROTECTED
