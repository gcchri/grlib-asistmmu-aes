`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rVqn/J3mUOpMUPWgu+FEV+GsE78f9geC463JaSlhMTigJWrr/xIdrfD44+hmfWGX
EovJZVAYICQkPg8G3ThbPUrXRqVx9CZhVWrkSjn3E55/AtkCp873W6d++2qaI5Jt
E3aPuhmo6i148A8a84CBCyJ1JgDln/vqQv0P0v56TxLrUiC/puSnTy/CWeDaYvDF
H7C4uZNZAZKthfYll+d7RqVxmFONNEpd0jl3hX/kUBvtZtWEn+nlHwY2S19ysMBA
6roD+L+17PTzOfZE1Dl42GV3JNSTQINZQ2PVBxDw75slJmWIfF3P79rv8hl0j0mV
3jLHOaj+Htgek520GsUpuwi/5j8BV1aZLfoggNdxkygLooTiJQtg+bd0hRXauo4l
0+yq4ElWxadaVUJFqqPrwIotXbUjExzylNpU6sbhJ0L+NLGsN9T1uwjaa6DM03b2
OgndkXJMeqXQ/cSJPGMbPIXor/kfwbCkB1oBJWQyOzWmm8hUx36uJR+sc+6hipYF
Y+gSImbk42tawMiV3WVpsHhjAmWfsZ5iPm9XmpMA71C4Ga/wOrfXQpvmJGWPUcU1
Ox105gxga1igaGYTXYK9H9ssZDLH847Y6ihvW9/Lxhv9V720XUy5R1/H9N+5LfZ0
18TYirG5v7Z6mzPP6l0CZ6Rm9BRjiowvh53pnB2sARrnGx73mx2XS9evCd55m1UV
2e3rWfSOFiyucqpwAP51be3pap1yWTQTSJMMhuHmkz1pAppbHyKucLMlx8WGAKxi
R/dZQ2wSgaGEjKsIM2IwzRqJkvW2t4BUtYAw48gnm8VAXPbp/fCfimC04b0dvKXW
mgwi63PhUjsnVee+uETa438uLVZM5C/MWdjDH4YTZSUWyGq4K415XnQajZW0stui
URHVqrLEtZFP9jYT/fbG6wKrxvreF2rIbVcD2AR0HGKYXGfNr6gFQ6uT/vU86hNV
H2hlU8MRkaPGC9eMyg6l+6TE42nAm35f1f3wYevoqpuzznCqVqePVbixJkYN/DVu
vzUkfJBfQs3zo9cR1+jPtxl1AkCdQ63+ualqVMomPiFCyEyActT48Sm8VJ1ZZD7R
6b0jUwu52d0Gd2lwXcI5gfHKeySjc0m4xYXLnWO7tar6HPgqTVqVCsY0DK8BCCjY
qaBmeVnOWcebQE3QQLUJ+kLgRbE865a3dyfAxhTxjsEWFZ82z0NpFYmVo3rmmHP6
rr57LtJN3GtcOx5OiPff3/TRxEr557/83vFfQpag32JqT+EwVtADhFlw4shmd0Z0
U9UXpGwOz9xfzEsmV+DslS8bPcZP0NXNF0eENUg3kTKn0hPuPzoM8VVo0ZvTnYev
LDP1EzBgUkHrigKoGpJoFeMGhpjQfaNlcnrP2s8zJz2SusavEHxnLdhtpD0oVKdn
mxcMC/886uUv1r2+PvpaZjKnOnfP+4aQ2ZhtccfEQK+ddPgcF1uW9FHodO2d6Od2
VyKYKViClEmwq5wj8em3HtN0EVeFDbA+DoyqkHQ254a+XQoWXRddNSuog2NH3zpK
xYYP7m8P5nljmVJDIYUGzgqRcmOUmEDLpDq8EvNqTF75gSl9Dk7Y2KdUMkDYKI3B
VWCyIVHIYohMd4FZharcFmssJpkV5BdvU7zikX5b2EsG/UWxNKHBwbKlQUnyjR4D
m0OKUQQN6dmC8/S/l/7nuKYnmQe4h6mEBfUmOv+z64gHDfWcDkfWuEnLDxFQF0Mg
bcxzgsLasnGg7L4FOyDQ+KitMlKpD+5LCDZTyTIvELmRE0sZORBNU31+TWCRWycc
9FpQGBqikNw1AU1gXRBvYzx6hSwjIa6MSX8kAORxVztkRZ1h+TeXQqxUi0LXy8fl
VlLv5hV+I6CPJkvmEH5NNhzLjt7Nafe5JCMApdQiBqAm/6ybqXXOSpNSdsStcXjX
vlFPlKxgQddQVEQrJVBWfSpqyyGlcBp6ztp80RTPEAAUNIJOkH8nu/XJDUzcqaYp
utvhUEPy3S6H1ag+BA0THkbr/ZzH3MU8NXvsHfOKTapZ+0yri4eeSkBSR7LhiOBI
4auyhmY8VAHiCzWkNrAt5nkfTnSKFaBJLG2WgrPpnnBZGvD1xwtwY3yoKfrWQK60
9Nx6FPZ3/Qe9QCjkM7axpqTGrDkpPVudr2GH+9o8sZbu/gVHiaFLVR00zabirZNs
X/upQMG99g0ZtJnuP+vpmPcryaosdolCyDPuhTQBtkcJH9TZw/mmzH7V009juCsn
Y2iBYmDqMMoqzKmWvxcmoSf+Ay0kN0kkkczxSDFfNtxWAFpyZEpjpQCh9bzSDPXv
WOHMGch0HUemGp1y5HrhtKtihPULtwNj7RiCfF05/BaLBn803ZwDwDBo1OQehzwh
wVDkki+CdgAkuBNWQ9Gyoa+ilSbspnsZ9peO3na7mkUdEjTA/0WQX5qTKbUEIHhN
ukImmS+sV+5LguvSY4rJx7g+M0NlE3KaxKF25wUXo0ehjDMlyaS7taSe4tlkXLCz
lAwnEYZxC0tHLemEHcdOjEe+G8vgFvoNMaKf7J1WWr4mwtB11Lep03bU+QMHfvAn
NPDH3GgH6hvUBkg06BB1iIgrR2c7By3cHWg4WWMKDKJLsf35JVXLHOTRXcA+Xaaf
6J4R/5ZYxwwWVQD8NLfSWJhufp3DROpN6y4xCPxg2rgERKyMgZQaH4W/3+axcNyI
0yyb2L5EGfZjG02rXTWJHFIyEJEsySKXL+fIcVRRxvALip1L7CCLx6ngRDCXE0q/
t+WqHrvu3jqsqUV66puQVwdBwb0LPA8cL9bQaTOa3sR+mppkpE40JMD8eR4BvxRp
dkYxxu7fTeDuzCdnv4sziE1wrY9y3KV+PwqbG/Lkt29yEHdLPHoMItmjsRDUNsbc
bF2/PTsjuPhxbx01CGywnAw+DwHB5aIXqeImHHRrcob9XUI11ScjBsNhdF/acYZV
d6YU2V1/sWgkfohnKuN1ZC2iljpQBJjvYXOpfjdMLTYOYK/r4DSwpTf5M7PGSLen
GA9k62vQCeGxh9skKF8rc/8q0omIQcwuCYsDQlR5rZpAVTV1jaRwgbviG90NiRML
/Jt8YUKniYl+wNf4E0HUcNr0KN/WrWgzHpgReVnD6Rxq48Lj6RvQMsQyKQPubHsi
8FQKfXA/nb6KpfGognYczFojKsCDAyo0CewDteZSAIvMbFmDbhLOmQGDCE+9m5jo
LQIFDHmnVqS03gPz/pXSnliD0iX9MGza1Bcb9n6Sxbynzkw3Xt1C74d8SL2ofEmD
7ieFEA9x78EE/iXosBUvbY0a9cTekGtvN1kxq+iAAON4ogXDrODQS2l98Z8IntN5
9T9OCkjMqltarNbFv9P9T87H2+YdPT0gjJ1HTobYso/ij1wzTXWQojoxHr28swof
RGI50dUEZZ8bWEH4h/a/uOxlmoGQpJxpJeCQFPw/JUEsNz90g4FcpLIE1521Qv88
Kd/c7Tusoa+Ljej9BLDpjZmkyfhdK8Kwfnm/w3SMz+IeZvn3bXODqeM6FPqG4r6Y
Eu9ejB0ItRoZBgLbS03DGlHVWlfxkStKJc2PmQrlKfkTriezXIdSpKqiYuB48aG6
Q2G55dtEa9vLnDpDntjFQEJcVw72CHylFvZVt57dmNtybNqkh4izA42a+moDACxl
XJQ6sOW3ztgUn9DdIwqRml9umrQ1VKQDY9wKYqpAIKNU4PCqSfJOYQI6rly8Eapm
hsQ4bWEp+LX61BaTWuvxEhBT1H9aXQl+NoJt6WJgAP/vMhcO18L1M3mCsHnPGZVH
AqFZbPZ2YwLS9Om96HiZJQIggPOvb1IECtMAFSyAk/CrkFXTqKBdHfoyOSrF/UV4
847MkObkCOxKFV5bfhFlHEF2EG/OIoyQOCcDD4WVPUxA3SunErZqeVl7gqtfQKvp
C0KhcxLH98PgpVEGeWDC6rAWnJCQwVePqGhBu6ZnpERpUzSZRSvKWPRQ/z+QV5wu
41NspObEIi0WyhGyp52fUf14Bhw5+kQ9ZQwoORep3fKbuC/hSaG/wOefxVzk2Eo7
5ss1lb7IeOqv6GOnRRsRsC3gYEWxf41U6IcFYqSsjesr53uCHBvuG6XdqMwaFS3x
gOkcxC2BjgiknuleNQE/TFHbQcbSpji9OwFjbp6ZO4IdI2XPSFo2moXGcmLrjlZT
4xX4io/bYw9E4vklaT6xIwi6dbkyf4LAEpba1QosCshhGT0IHTvlZKogUHfizpAX
wD9HsY2Xehsrb2E2NloUxcYlRsW3o6ibMdmK8PlNadHdpuFwYX9r38rmzHgSOvpQ
LF48jEto5P/tFzv2nz6P+HCZsMgroSwKtkXoEY1dPwAu7p5BLv5ar/0rWm6vwHvt
qEPXySiAd/HD0/4hIpeYxpEOVFRrHv7uwZ0TSHCcBFqbXjhrQVPGNO98jVw0yqsx
R30x/Kx7XPXbEIpEajg3wukNVo2oDAu9hxgqdwfGLYSk9u2f3C/8doW596fJQwPR
nwp0F9FvvGnv3W/bmjnxL3ip+K2LufKlVue2ulAp6SBMY8ef8XGB92WjzvQSfEHT
sLzuBLSlcMWawE7euDSIKtxTI9JPrt59E2WwqRekmnbuosvVQq9qY+9cuOEC+vL5
CQ8KQGrPuBBlIk9zzKIS4lfHPk7md9DCTuxcpAC4KmY6pyD+Mk/6YcXa1Z3pvlgM
HpwzeFUcjqXCMONpT2DAlGXU+AS8YFDOjKCIVYVHljQl+PoPkLOyOGq7AMzOCAql
JFQjIsW+faqhUCIY0aB4+J8QgQWhmYSxg6VIRa9nhWXgIqXJeSZcHaalhZhfniK9
eM2rtHbsuCWCPpmHxsScpixgLbLfp3CgErLkaXUoX2E+QNJdwIqtbloLEGYAFIP2
bLJVIuv3jjEOBG8QlqTN0XSrwqTg9s3PzqGxJh//pwmKbDBZpZbwKitL4XYk050S
RIdOJnp9qjpscwM0Babqp7RQQBecXLvNCFbMB8yvG2JdW7avmPd6eFZWP55FAN5F
CXasYQBduKX0j6YM9ZDKx4GoSZvCOBptVExQDoHJEebgdHcI1qW3191P6EddS0kk
vam0/qxDEajf4C45moSEPC/wzAWog6PRsjwpVN56p+/w7UzJtz51+Fajs/NhaIto
ocsNmkKM3EInJ/+EWpYj1d8bjdVtdUHG5nDdbgWvQJz0q8mlbYJ4yL2dOtnkuUeO
9F6pU3lhvHJPHc3g6j4D+LhVRc9dcRdxwEgvNZJqIM1dv96ouor1I2L8M5IsjdXn
eHiRLPs6E8h3x6iXxa8h+gCEk0vQOv7uovPzSWVh9G8=
`protect END_PROTECTED
