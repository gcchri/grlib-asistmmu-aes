`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ATIiQXlQV3WXwz+zrsnyazgZHSzmnsRnGvC16oL+kakY4M/7jt6W5r0rFNy6EvGg
LGTDgLtniWkETXFQzofJQ4wQ1t4M2ottv9Wsfg935y6dZS47o2+f40FIfB+dXlmN
EQBHYdyYZVRDpgIyb3mwavY/vVYVGqRHhdiWJQ1kSJ/YytF83Jsw3FZI6wZuLsFf
vKvwczfvZNwTZ6nfPWQVAdDl6AUC3a4dJ/EFUSpnNKwZDx3TLuwFMUjZ+A0Bx+TY
2ZIGGutzxTysY1ox+uh3Bmh2C9y7Mpk7zd66YIoj4Ko=
`protect END_PROTECTED
