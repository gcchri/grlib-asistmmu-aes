`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Suis/spMjt8RXAFCT683ZPse14wX2LheQv/rFKXjtfgtD/afAWyDmoN6hpuoaA/q
YR6jn2igdUrwwfQOEuHaRPX2UPnHY8l4kw9/hYZjPUAwCD8v6oIgJzTB5ZjBSPzR
A8J39rbwdhLrTq5wEh02rSIwm4+8CmgAOwZSrBbrFTTI52G508BGdHadBiAOgaZi
kgiTIbOpfOXELs9wtneVoBVZ4nMyVTs23zGSr/m9g23XRgx8HId7gvpnsd4OhuQu
ZzkftAsqATJO4HcOqA66DVzItRJHNkz/RlaKcJp+D2I=
`protect END_PROTECTED
