`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i78GLU5txC5Z/E7WfBgaNOlGPf9CWOpSovv/wHE00u44trHw7aVPlTNmryPDj66S
kNqH1j0y22jAvi/haZ3XzTgCayQLeEg/u8CNj26A5pDQDABzxEKWWK2YkbmSoTlW
TS8ran2Z6EYZabEy5RW8O7QibTX4KfUpwXCU9tDGS/PhKCQKpVdjJk0Ogep/QSt0
MHtOahCsXokzJtFyIrFkNPBrt5qx5qzgIjqNGs1YpfnoZnuJSLuupowgUTCcEJcl
C1gOyUN7WzRWBzrhx9SdBC1+csVzdy79Heu08WiWGMXWiMjC1c73ZVAdeCjJx8HD
c+gC4hAtxMByObd+tndnAiNA8AnuCpWpkB+PUpyvCHvJQ20VQnSrg3pxlwVcx9FO
lK2zxex+PYX68eZvwps63CZHi8j1ZgSXrAIHQwCQNylEzElWaEcrnuT2JwHfMVRb
tZOxwa8uNgaCYwxyrOwTG4RV2knQNTxaNrSZ0TCwNLHbkkl6GH+FUeJp/knBJqtk
`protect END_PROTECTED
