`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rA6j2nhA6yhlgWXZzhacOgeV2ajmRx892Ga8PysE9JM4oBQBwk4M/0nPjXxh9QgE
oMmHxP8BYId8ImqC3SggCQfBfjEdeC11vsMO/rYSo2SYtCrQp2dmanexMljQQh4U
zPcL2oAR3Y4xf4jbNXIsgpvLwxcf2AfMyJaMK/0UXyiklKf6fKTLrareNWWrCX0S
4D+l4/ipJgKwuSQdSx6v6nqp/SizZQq46kx8/dy/5F6YMZ0EwY2MVn4h9D/HMCtF
LYE+wioj+avlhTWV7RK+Dg4tIfRCceTsWRWE7jX0HEoYYdGs4j9vGSQCPxgaMl//
gu50U4iEVMAe++UYmEoNMbaSVlkqBsZLG9YiB4nyL9bF320TL/Ph4G9DJjyxH8Au
kz8YNFSVJvmJOUgWtLvZcbKVIemOGx6tGGl7OCzarB5ct66AoJCt0HFI7Qv9uLP6
mDTCkTegGHMCIlzKPV/qRBK5rs5IO2yDXbDv0V6/hNMcFDs6CaH09ArpjrJ+Nwi7
4kX6q0L+Lw0NzefAB3iPgA+2ponge8rWxWs+Kf2tlKNwltz7SPAJmHIio8vySI8x
26PyDuUk940NyEZpg1vSF4FsSAy0sw8nS1NrWMRerCqFHZd55saaRxnWw2rzEdZF
`protect END_PROTECTED
