`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhzoAyOK8Sm0dA3sxXjIZUGSU7l1LiKwDnUguL7CPCDvPEg/pTG+uJAiZ/7TrqHD
/OjM6bCc6e/9R/ja7G9oG/kFNSeluD9MR9ZDIuaa3oQJkiKbXlmsg0evufejZgZ2
2PFlaJIEPniljNjeic6jRtE6M7Jdav/PGU4mPT/jG4a8j/Rd0dzXpwWjSfylS80V
DTnuE/J+oPmLUYSVpIJb/Nu0uqHJzV4EFGoJSVjMBBT/1i6uXp6l0fGXFwJd3ttZ
SD9Cm83Ay2oWCjoi1+qJag==
`protect END_PROTECTED
