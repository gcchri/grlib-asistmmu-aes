`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qD7QKQjCj1JO4b13SBr0Nh9NA5YjuE8gpzMxFCxski69xqo+WTNEIVLh5lRcfmxi
hXQE3vSGNzzt4HKnYxWM9lBg12Ek5/Gkf3iN/tZPjmskJKEq7qhhGEXHn60aXxRX
ZowP3SDUxlqTskrXXatl1rn1k1SNPHoZoewygTu4buGbgC1mrewM8MieF3YyY9mk
INiAbhVnkLCNFBd5cmuWWjiFMkkyH4Y549+jJ+NnfKKnOCAsXFGR72r3KwJtb61l
NUMaZOWKninDAfTh35qXG4h1LSCiQvVhQ/keHMgDLtYQy4P5Xzrbqao2k1s3RMoi
mcJ0S6JIaLdcN54gRUZ5Xg==
`protect END_PROTECTED
