`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJWXxVWONRdAEkSX0LnOS625U1fVHBQ3SVNGvAk3UA1bGgyRdOxa2Kr8bloApukx
k6+Q1Ed0beK/g08/2ly3YfY00Fi0setMmuteAA+073J073+7IRBBxX3j6Ec2DKEo
eeh5bsw5+4MNuIdjp4v4PVZm+pe0ZQ3sZ/sCffFsD7SbRowLQHvtF8JdcHHlwCck
3hBt6oIQiFfQJ2HJAVTsq+VK7BZakkwFxG1hoOGd2lMBu13pQtJqhCgu9uZ1Xq/G
Yv6qSIE5QTVhf7RNwpZ6lQ==
`protect END_PROTECTED
