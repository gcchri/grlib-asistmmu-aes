`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nofmAqRuuyajf3n1ks+OsD1LMlFDTwYFOnxLU+sdeocoIdEPJ4HB3hXVBSCMlH+u
S3JnHGikbZQVVl4EJM8L2vJw50b/HDadD+I+YAO5qVoBVLczV+K3sbkHm4BWvRl3
wb5tvhGq6FYj1O3ZUK+Abfr5QPbTDFJoXhof/gkTggiKkL3/PzThwAm2Gjh1U925
38AMs3EsElHzKW9ljVfte8ev+fhwhik/vnUudXblwHcfyB3FjDMd6scbY1b4SxzD
zXCxwMvuVo+iSbHSRFF0qe/dmLyKDTcVrTB8zq1V/vifMb2qUr9R3kKUKdvynJ1r
jSto2Ia8AQ4EuzabtV10f+2hO3XMCG+NSYQR8J0edhrObc8QJmxaRysdKU3ySCFl
6CDtfiAwmV5PKKCsAVT36nCq1l54TYnDN5wC4Ddu8kuO+NqMGSG4iit9n+6xNY3i
FXf8pjTusBMEe4DjAwt0uKCUovDYg6gmy9yoTR4TzdRNAG/6IMTXv7yvQIMZYXGl
3Efy+3i00pBE2en69BounbVvKeVJe5ux8mcu23AP1uElLZPn9cDIg+BKSvjS1yiH
OWV+YOyjSIdzLFXldm+t1lHdQBPjyZJW0+jYJhdbye0Bz4yJKPzI3GfJTqQASQaj
+OwwBi3PXuvdOlMkUGUcChCqx4Rj/D3DG93UI4uwn3l3MjQ8q8xfnq7Os2sTL/TX
4KxzYmn6+Xj7U52So8EsL5v3cIEf6U6gbISq1Jjmk2tjsFXBBNAzoZvITRcJ47Y4
ghcLGJJMmtfdGa8eLtAuyV3GDHkfWM77aRPU/hsC//QkN/CZoiDLXdfnOKDWcWLW
/Dd1KHm8KaXUxlWN+NuUA5BQLjWVXiKjMrsA+BnC967Rd1gi0FK3TLls+TkveoAQ
A6lllMexrGf3OgaizBZ5vrGNFjDnDrK/LTjJfRIZf36LKZV6Vbd37CkBveDFQHKT
EJMYAgh0MSTpBV2bHWQLT8hdTsRuMDvYEOTHVOe8VecVkvLit38WdGUeKTee54G+
3ptmJ1iiJP+6KL8Zbq7C3wQEoPf6AVwx9IhIYeiUSoBh39RLDDWzK0JoUPk1aPX/
hF7n2DaQfqRFWQ5x2JGqUul6M+6FTNhoMEy0HwZXprQGPBWvgiovITYuhUnBCHRC
i0mAlD4YE7ClSuC2CnEA2n8KJP877B0JkB6xqPU9F1NTMHJ3P3oZ29A/Jmfy54nC
wZnXohwUmiW3oo3NNFz9GUI4fSzSCDzBKmvA7BrVPiiTlwwHpeBbBYoCd272k1S8
`protect END_PROTECTED
