`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K74At+8aRe20AxEcjcC1wZCXVyOxDRvHAyfbaxQC+Qvf3hs0NTqLZuKocXPjyLgG
euVG8tmgbIinMDoPqOnfhPVe0IUbB9578dUVswEvw9pxNclD/SRHW/ZF+WW9Bm1A
gHhGK0b5thwdM3KmN37FxzuPWZUTkxJpgpHLBTAV3Y0j8+P/vFQkatl+Ts8t+/W+
Kmix1B7AzqaVahmLSDDrZfE0aPQtWjvLu7iADVulVN2y+FEgzPRC7bh1RAxZsHap
FiPWnyZYc/6OrVRiXnSiKfrAbkQaO4yylm/Vpn3KZk4jfW+87nvpI+Z00FZLlzps
TIUrjRPqYnImgqqdDN96dzUXyHOsArWCB76gtr0KkJOKKr72P49NJPWGJH8bgFMO
trZwrrpXRuJgVesrLSaPWqRwyEegkJdcvxAyQnVntADyJ+lDGF1V7s6TC1relvLq
K5ZDlB7IeGnhC4HIH+ksiNFJmqdlrdc0P69WI0+P33EB+vN/uo00NGc2wrXoT1UA
JsJJXCyhIIXnJgHLbREuwmbvYiMBrMp1m3CpqQ9wKY13BTgShkYQGLZsRsLfWReZ
2i49u9MMw8d3lDm9gpK3RUqycfXccsrHAW1wPnG+7R2b2KxC2OLRwyh5R4YFNUE3
QIXOVoMOAtLZG+AXsLZZABwqhWf+Zf0KRJ9Pq2u4yYeOzFXP7bxCirBZ/r5BBH+N
ZwHzigxFeHSd0Ziuew2W939L3d9JDNJWwIc+1FG6X3/pZ3GcMjHJC26YpQ+JSqyR
xlEqGvCV2SOGc2XICHKPtdk6EQIjlnewPOPRud3ZP8jXqzr40VvT3jz/3KBtLOB/
Zzyz2qnwzRcPdl/5AiwxK0j5ZjDDpKgt+5303H39FpFAOi2yYGJtaLgnvBNT1Fn/
6sXcLFCyq4gP5VddatUp9vvF3xyp7TJImTddpZiY/L7oLVc11XT8Uf/VGPfpOkYt
/QJ8JODo8OT/H9HzikGPNU9YS4GWmh455Xlmsall8eq3Bsi3iZhPL4YLeI+AaNme
mi6Zbz4yqspwtsFBW+Tt/JMFHtAgnewGoBF6403CC/1nunzEqKNaaVZtOuhQQ3fr
bzmfExAxRcUIU1jts3bI8KvgoGsYeOFF6uzIB02loX+d1AgT9gb87hlIxRWVMlFH
BxElbCb8X9wYrlk5GnJpJscBGfLbajy81g4CVvqcAfgmu/5AfvPgYzXg/qm4D5ye
qnL+Ntb+qcFRFoY6U0KiicvmiQbmdBM9FN/I8IU4lBlkRee0HJDVdTj+kks5LCjc
wVeGqYyuZ6qb0YJjH1uu8KvWUJ1MyW7iWqh2X6kxVeYCBMyUv2xPZ/NdZBtjIIFq
1JmOIp2l+f81e7udD3bosj9qj7wxDpc6lKF4Tr4u1YtC2oL7XDPhzItDHr1GKkTZ
DCRQBFo3IudwPLyPrJ0WfvGUCZdNvKDnZLd84QeR8AtmfvE7EIq4oITMGNJqGS3r
Z8eyc0Jh/QWlJUedRg7jE1+x0rcDjBpQ0K+bc/M0By+Sg0DNcWTose1Z0spJQITv
ae97TyWKAgv+OVIdIcD+2+BHteyKWUMWaxr31eSwENONhL//4cPBmgAwZV1Z4mCl
ekoPHapeEizFueen6oOzlhJKAVEAGS3XvOc3bUFsVRBS0E/At92V45xZAW0HyMB+
JpYusNVYB1DeMZ1bc+SdbLVOxVVgnORAtK6P1Yj/75YBnKDzpycGSWexRdTWpLFL
+J3vTDBFyw6EUlU8nj/OXPqYr+A5RZ7sR2dywTh31dLftjdiDiz+DvG8tzV02CE3
S+MKxv8yuZM5xy5nd9aGUXZYWONSmUGnjOPaxPIzbpI6T+48jz4MFemLjiFH4Tux
kW7WE29TSv68YIC+IYvIJ2yx8eUj5KQtbn63qWewk440YR/7A+j3T6p12UCSG9iP
m18ucO8AZcBw6B9nJLU2b4d97HeGyXyyjo+VMFj/2dg9fNyfM7/pICJpXyl9ebjz
f0/CwB6Rdny38T7bWcC/8PpFGLuyXKYDBBN7CfP1e1OZikYvVgu+VqUYnYqcIQvi
4SSDoJHWxsoxa0oE/ERvEP2tB3BwB4aC+Qgl2xiilHmeDQmtBbZnyLicuMyyZLuE
iYJZBtVuLnb0zxfQDar5E7qt8/0e0Kj4bo+jAMM0saN1xkxAd88GgpC5e+AphmoT
SpXVNB0lDtxBDKI/BFjX9hKljU3xYWSY5v26AcNdFd0lcXxM/gGb3O9ao4xhffff
+etlHPqtmOWu/Gse61zagOpHmFJfzi3lWkBpSa8ctDKFhEE01dZ12g1C+zUTUGNK
xDVGAZYJjVHZS86qzpvY/Y9NzC5veRG44jw4a5iw7SVkrxYPhuey2CGLZE8roUwA
lpANfYTO53+FaatytN+os6FoHTddrYvjWB+iwM6F2yZKiJJKTafiwJt59tnNiO5+
`protect END_PROTECTED
