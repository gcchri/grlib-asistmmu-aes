`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQZZQU1k10vHyQxPAWxSrQVNMoLniZ2l5V1JvXaU7lOKVQxZOxQLnLuM0K13TeHA
8D+ncsggN0D9qfvAlx8SH/tZhP0QTGmKOH3mnzk9XZx07smbjNqDJFShYVrLvkFf
xx8k04kNAyN4leDBYHVfbBuS0G4Ad5Q4N3oIssvIGy3PxSfL6+RXqGZOMuK4FK6d
ogiuuKFQdnsjTsol0HsPNhTOtz1y8yeKsS7e1ihrHdnAcmiTdXlrBGnK0meCKknt
4omUdTUiz6tyKTkE8/b7h82O8fWfjuyWmRIVlylCIeBWhYg2iByM871fuy+Gu61e
fVjJOmGFHaV+MYbFCRXeNyZIM/DTGnkmTftWnXlgoK2ZMfJXlC7FuB7iBZzm3fFw
Qk5qUS5FnxWQYr5mf89W9qqmZV/E+i5z0o8sg30ZUl7aq8sVSNcMek6eunJlbGHj
27nszVT340ykXKCbgWQJPVMdkFuKv0RWqWBu8FFBjCWY/avBy7hu+hxFUGe0i16t
o3W9KcXi4Rg3BkpfRvmorf0FEbpqZYM4MUjy7+/VWQqnhnO5LmaP8ZCuEObFOKzT
8Lw9HZGAaZ26RR1Dl1HNp1NWSNGctfGOPrk3rB/+5Y+J8Qo7FjKc+HXxMHojSDjR
JpxXQKtnbhbnzhojzdCxBzfPmnzrEBJrWxgEGMtdfYdmkc8QtJnrw6HlNU17cas3
tLYXdAANJthJ0Pf464Doi4v4h+YqHVs8aPyH24wDlQKwzz2vP7hQeO33rRecE9QX
ezQubWr7XIvj6x0uF5zByi+3zSaj5p6b5RP21MxsfjPU1ldRbore5W8LfwyLZcUx
6MsNKkr8C7RSycJzBSGmwkZYolTJYeEdyhHbE5xGu2O01rnUOR5Au4ewDmQaUBrO
dw1gXruWShjN5UAt7bWT28ykBsPo42p2Ko9b02wDIQvAaUkT/bfTaItBZRz/hmun
LrTsWaFJyBvwvxrtdLoE7CqrSt6rao5T13HWYgQ4Opo/bzrSuHLP4I/rvir0laLD
oUeAtkWRU9RpGHzHku6KRI3Vj5joRxu7jonjiaaHhUQyZUrMbP0t2CRUUYB1Tr6c
jXUPUjM8IqKsTL3pel9hkcq8NcSzPy6NAvKq5wKAIGmtZkMR+Owq6SRv+5J0WUVJ
pAA3c28pD6al0X4oanDklrLCbK2aPjXqrfI2uOMyp1uxIMXVx8uKmPCx1GfGf7GB
iSGgWlbUTlmUz2Pwcb/WhwTz1OES+9+Fc02HOQjPLztlK63Gx+qba7+c+hHux0VX
bdxaycrhms7b402Lo2ZiC64+LjLR0ppxg8q3TdpPtQV8H7gWQEzYs6sExCVJkWTG
bgTSLGC36i+izFmiB++dy93QbBcah7Nh514iSwythxDXYXLHRhPWD03Si9ouVb0i
fUgV1ZpxcsTyfYhz3K4aKVWygLoQ/3HBFsYYHRk0IJ2lpjsQcGxzLIvF+4AJuj5E
7hJ5mcG2CmXUSOhbOObxtFbwL5ch6NNWa+tMh9Xbo5RVzGmBdYZxUNtFfd1PTkoE
WNBBq3owxz1hqctABhznUkh4YJoF4MrhsXvW7QTKyAuiimSQfhTJ6eKegG71SxmH
WmiNLeGWrcclqQeMNFn9ZrbU3XHV9VpsNqI6FKQBJpFAMhsI4/ZDMworpvNra29i
VAkSo9odpjO6oiOquK7JYdKzXHKL2Wc3MIA3tVh9TBnQIqswawuyGFK2ZPss6Xzw
wuiiB1uag9ltR+u0jcIGwn9Gj88uugMhI+C6GV706zv9VEjb6mK48/tK2RUngH7H
o/vUWciVshczGZaHjM0QNR4ZQ9ImFMWDGzFZnTMKmEJOEM+J17+GrdAA7yETnFPw
OOPon9KXEF4n9HgkXlj9dNoYqmkKE2Np3io6/Iz17TDjhb889dLeaInVowGGA7I3
pAy5GpUoBjObeQUhZuFlXNXC4kjkbxpP5Qk4Z1wHcWY5dHGthRkA9b6OZR9fsZY/
LFEDwwTNWO6gkBMu3B2v11hsEYk2mHSQRvXqMIKlkrJKymq/DEUFkM7DabPS2Css
HvumfB6p7FXHm7Ay6jgRq5vlX1N/v8dfVz180m9jBrCZKk8l55hBo9e0cUqa2zwz
Yo5k5Hdq7XHf7cSSO+eTh0b5SavA5Rv4kjfkJIN6yu3udPcOJPVCQnrHTvo3NhZX
FJ7wu9bL9r9oe32Wn2ICI9Zlvgu9oMZ4rVTZjUNnq67Rmok0WVdcjvKxKg9tmhRP
CWGXw/dSq7ADPtwU4hNP/BIrO0NtvmXHOMmRp9ZV76IxqKilgY64vf8XQ6vIuwbK
n7fSsJgDK3AVknCimNbtzb7ewj3QWErGDN7GbCfiUm5kjpM9+ajNCKCvR7+xQugs
h6OeOFIQJow3wUMd/mVq4FFswQbvxdVfibpDCG+vQgyk6PJKllWejaGssggaKgN5
AXxfqSnI28Sh6yDjrSrXfhK76p0Xj5M3Ad/ybRC8//Sys5g4HqSpwkyXWya1XRIn
miEvkDHTXTlW5jt139GVlZggdRzSHHHNq0eMXVoZdh1aBOh/TYe0jkhG0wFyxSAs
ScaikPxOuEK/HnWLpU1vNAaiR6pYHD8Ez0e4DhcXaPfMS5XVDH7U23AOInZpw0MV
O3Wb1c6+71Py6ixInYA5nvNoJvSOg0q/dVwg9x9A/41SYfwtD5vXBkeEIuxAMlQe
5YmG/Pg+Sui+UOYCJeK21wlEI6pEOGmFELcjpGOaHmuZM+/nytCV3TBfRgcSIxkl
zEpAkeotA3wRTTReAJjcFxd3uMlUMwfrzsM6vGRyNWZYOFHsQpE4uBAWlgTO+fcY
z6fqCAAZavDjTAe4FFbz3X/45bbxh+Co/Mle9iyeCuqaOsjVZICqzgmnZyDlsSxH
OnM+K1i60pPZCZsBTIVz3MQ93WASvhKBF7SnOIxleXNSX2ZrqT9Jj5OqXWrhZatj
dn7RgcN4NlhZClwUQWpBrB9/xPWt12DHWGj0bvxdajb9wddODUw7uWHVEb8oZ+eG
aXZqI6VvEBFFE1CEbCMYYB0KYwpMN/kPLVvT9tJ6O4v0C6wcXooE8E57FitaNeTD
+BJJnRWWk3toTjq36LAIi2NPZYGEswITLYu+xF9diAwJv/1wqprbTLUN0wJCubJL
fJJkHJyS0ZNJThUyFRAt93e3bfix8YAK8NmcCXiuYcEjy4uOoLChcCCBF4ixKB/F
nrU32qEXYtVqZ/ZIYzzMQzbNHaD/T2fOeJj6/OqE9y84D5KgzssMJvsfqQ4U7KUT
poQf9BwX+MHgMp9t3bbQv43s+fusOmSp3UurLRKUKR0qrCxwHl9P14hKSdGlNFTO
5bz9jRjginN2khHSK1ilyqL5Ee0tQnuyI7kVse3aAjpzfVhHxUIDG4xhqHYhx53g
DIQk63G66ngobR9f4tmlqDjYOqYhSKvcsyDVOhN/0pNZ0F+E2eXOgqfcJb5Z42v2
KKoa7MH1IrdH4SJHrZNhnK1tq4UGaOTI3CBrQEeU7Dfj340XdaJ5kMK28+jGE/BX
5oZnZWvrzIatMpLGoTQzxHNQnddayebcRJ5gnLuV1pNC0ZGOe2Wb4VyX+FN6hD7t
0aBbiWcO/NZypRktgMQRGKV9E4+QD3edMyw01YKCp+U0HHbLUPNkVlTyAf+i89FQ
jIA/gUfa71isI7+vH16/Riz4JP7l/bUmdNZzpUs2JVJgSvz/U1Omo4csHmu+O80X
RwuRMylvhVJUF9u5RZQmBHXsklID0Vs018y6WrjWgOo/w66Dq9llnGw0+1wHkPb6
/Nfn0+imkA93sdRNVqAJIU8+kD9ru0VbRQz2165/C7ndXYXYalNGkuHhXIMAPlXd
1iYiJ0QDXBs7qcCc5vLxianT5PKAH4AeTvjRE3S/0HJr7NzoZAn6XAbOO17QJ6Qe
RtWe40aV7iSnNL/uhJn3fOsqBPelSzXoXlISfu5E8dY3BuAPQ8qHQV4PTyDOmayX
QnEG+5OqlKOhEga3HF10qqPGJJQeswDNFlfQ5YedaIoKVu0pI5oSb/RSyDWB4nnf
BrkNEvwgvbOETj30u8MH2SGnbjONw59RvZbm67i1rLiIMrw9CNouWI/CmNY7FQFM
UbnB7NtfhVtp+kHEEOLr8oinvHAvsDd2Pg+uJGlJXgrhyFADqMjAC2C+R/GdJhw/
bHxbT7sZD9XrsnNS9cfjer+Z5UKY/QbKlsOm4SQ1SVip0Cs1oUzqfOKptZsWlzej
2+ApJGPI5/covVGIMC+GQ3ees8zGF2qMSv+TCR4kIAeDwndropvGxQARs0oT5fYW
klaFQPF2TdXqGBuBe78kJ5qHSm5O4E62CeQfKZKlvtqFK1rjGueyOaM70Ulp0UYW
fRRU3NWv28QXvhWqwEgC6y4KZM/jzAfXpiPresJoU/pznlUjw/bJzaobGr+v+Fhw
JO91BKw4c3pqOLMD3rrcDcpYYLEK7rteqiOK21d54F9CIjg4nPfyMO525CX+rXRK
phhEBkl4UhMXZuhfCnT32tozz5gXsHbIbMjH7NzVDyRAFfx987ddEDh5YiG0qIke
3nJrFpZt8ELMz/WSHEQbul2+PdacUy5u/+fJwI8T5cpD5yI8FzMGiRxBVVk0NOt4
hk1Zm+X2XXXqQtar9Pjm9O3H09MWGF/8s+2U2s4fLSU09XUrX+WBE2FRm0wrU9TB
qcYuWhL+sHMIweYNvzPpHX3Qg2DzIEf0gikAiq6dWcABNcRD8xhsgZbMRQ2Jswsb
og5LeFAZJUCkpITMq59HVE7FJV63pm8Ixeoy8H1TaEFD3q32HVx5KkPT3Q9jOLwL
HlgQpZPa1/K5KzGLWUOeIO9U6P71sDyduuDQ/6B3UXgJpp2XCer3jt2N7JfldnQ1
3nzNf+DGZ0f7LHQmoMg7ANCvEF22hfGM6DFeD7VK1zdHmWVSxv9V6OlCPDXdNsl/
Zq6XWpbIxNmbxac2EfuzvjS/l/fUbYvSkMemkfDr+btI/La9B3kLyRj/tvSgLVzH
6K5thMY1seEuJ7wXHHCUV+U7S7OemD86VD7XLS+xMwBjX0dgqaGCkmeeHVJ0dORb
uogyBuJceIMf7u+Ia3cxswLEwb47hg/dGDdapZO4+biSMZNaG5pXiOzYN2CT9lWp
Jw46tjgM4PubFlOBrEHsmbkyvGr8yTER00qHkSq7hxRoOJZbHpTDnksfLzuQh0nf
qdk9idBJMJKvy8+kQzv+rQ7wqOcRxSyQiXm7ml0ocfVBVv/0KT11ASRQ/MUzTZv9
Z0GZuNMtQZHW2T0lvTFA0Djab6hSnMIkRUCbiNRSToIBllKikcr+GGIiaVcP10em
oNiolmPJ2uiacHIN/RNRv0g8WX4DncYUcSw4EXFXGdGksO3+7DRsmMgCmPr6Aij5
D0YGN2bUvMh/hT7zizjIUe4mE0hNhvO3XHh2pzUIPip3Nyh4+gM8NzckQlnqRYo8
0sef6GmZ9w2FuAVqwIpg15hfQf0yrmHcUPPO0wJCWsqRdGiJoQIHtYEy9LFP9IfV
yhPXZpvtIKo1pwO2X+XIIDZ3aiS01Ad3AaMs5nHLKhKG8KoiUuikdahzLu4nnMW2
VH3ps9g4DpZY6fDPcuhf3CEflY1dKRbjVuNO7G6l0B+jMQeeWUUt4dAHkNoAym8k
uf1SXYl6C9AHRq7PFwtONVc746Q/a6bT1HqL6NlWVbvZmriOcBQiHWo+fpXQxiWQ
fvnXU4p0USJcHoHb7KW4j6TzrlKWOD0NncogEAMHZ6OtQl/sVgzJyYCzXRxyLAgi
cjWUSBK+p8iP+lwnlUaP9UE56eJCpCC8J3zejB8cWw5CiohDEs8qS+qh3a7qPkZF
MDeeKtCOcWdAfx6oy1bE5i8AeDncgLT4qgS1Bi5DSlG4gPhPsgAfHmqayYxd3Ies
0PkoPQfHUsjFI9u8SMXnD3jTnJ528RtrJuGQeJS2tMe14LMYVzRD/iFHXVUaV3Dw
iqUldLQ/fLjcjuZqBIXBO/p68eEaLL/OpOsZPtBepiiIgW+JNhFaVLkK9vTTJuIH
a9ELnYxmv1F0sXErm2dWDw6Ebwy5HDmAX03BtCahFhkjlRrIX87nlRoRqkvlQAGr
+edyf6Z+0UwEmmXreZlXYa9cK8xiOcBYOYc2k4lV8SHvPHc8IEXKAzEnCxPB6lY7
ao+G0uDnNK5K2j2b576IE62MZH3aEypFYKIZ1HozZ8yWi3zfxPi2VQdBs39oroHj
irT/frd7704BbvrEGwdMEPkA07472QYst6+foKeXOWd94vTndG/L6FfMj7y8NXrU
3SjenLwFWP1HCnKHCI2WKwRR7JeVUuz5GyZAFvUOL031IO3I9XEsZHxeHFtwqRt3
2uPcQFYqgrI1xuoUAHnumARfCbdZ52Yok53HoAoFzI2QFmXPBECV6+Xnir1Yu/gZ
souWQ1Q+5jzMm48RQ5VoPZBhHDuDFGw++kvNKCr52350l4bGiG4PPs/MbL+zUuX8
q2h+L1XffaBCiy7hqKmzYg+oM8ePHaMQik7gp/oU46XiYJ6KuRZSTSSzq3SFPOH+
RsHpx6+fY7Uw2SmRRtSMKJwXKX6DjhSrfaLApqtyF+hhUy8xGS4WoeprwrVLcCI/
DT8dBdvNPOmdPIZjwNa9bLjObXW+QtxG/DNKlcZfTf6/lNvWAmiTFeEt56fgE2Xb
r/EzjpkBU3mQ277I9nxc3pkOReHIJxPLmdpPHLxJrTJYS8tmfPm3yJxa/H69+uIH
mSzotd4PIfAanTkmWd0XSf4BKeSJ3URAYYnYD/IN42HGz56GDB5Z2yPqIfb0hBK3
23BImJj47RET4AgVAcWscJ75dd7BlgKtob4pagAL+DORrNba2PFFgOqnPpF312d9
mN0WKq4/y5U6TVYMBLVSrJuz51j4ZvQYyec0n5lV4uGXQfJEvjunEB+MD3yhAo8g
W7hSMQub7gygPLGa6BGA74y56r7ftV/RMgF1WHjc/5DT5rtPLe1dm/+RvGFIIxBf
ISrnyHDwGmQ6hk81gj7Tm/7WcYAhkrb84eSpxnB73/FMuP59qWMAkJatqE4Ue5xH
8I5AMx/4UpdlLRKv8wXGH02QDdfy2KegMPGxT2kXYoDZ9BX5Jr5ARN77phGls5je
iP2TG6R3PvFvc86Cf9BTM0tJtCh6ymM9hypLslPBq7e6IS1zVGuw4lpXGcrClMHY
3+bhUilzVLhGh4VdlEAZhYLFnPnqA64utoU+TMB8zQ0Q0FP616av+OZNUNp7kb9a
V1+iMG7IvN4/ggUhmvlbCwJSvEslr7B14D+upiZNRmOqaEgt/+jdOzs7hupRhjF5
awlwhPyJ32+HkDDlyl5opCnb0a9sisEqzote75EsUDl9ehUQsE9ytLA2HOUzIhjO
FPghZg6HlR0pShINwYqWBxGPMhkVuJHLwgyLoNQs1ZF16L+WYuJfEvW+xBtlKkQA
sybz1iCtlGLF2H1c2/BCbqAyDqtGxh7kHKv1rzM5zu3CP9Rbs7mAIRB8pD0NQFYW
Kvq/fYjrqSc1Y46BSsdQEiSZBFtlmrlC/xYlncaZnET8EmZqG5559XSHvf7hHQFl
RHiQLQmnny6/bk9om+YG1O2enc4pXeD+ecLW3YE14aJqx9Rt/Fm7sMS27Ps1GZG6
hNZXF5yszoVdHoD2ykTKuXkI3Ch5euMKGVus3TAetZ8qB7Sbs+TEYTJiQMp4Ne+7
dRtKUdrzVcDwuPN3w1ORkenhPztpsVXmjiRPVD9QYqYjCBsBSK+Q0KGvZarXDN/v
4ED4/y7BMMSxAoAfYXsaGzI6+VWxsagKz/ldKgq3lphi+R8X+qwtpglcBp60Tq+W
9E1mxhPEVY4pmu9F8x9dWjFKpkiwxEks2K+rztZYbmnEHNyBFOMMgc0TEik7o94y
rZGEheoi64zObOPI5XWduG0NqqqukAqYRIr/d5KnB+udwXl+ujr/sEot6qQHSczB
aVLz7vJNmUou5S5oHxxbJb61VIm+KlTF5AFYzNLXM6fjtR3OSAELzMi3teDQBYn3
fextWXJINTI6qwRm/7I6qma/PbDTQ6KKf6j8MJZiSyoC88QLaemnKhx3/VviTl6U
+tp1/CsZl1Gzaca9z/1T07dJCkiiI8CTegPIR7ix+VB11dbp6muzNHxUiEVWArt3
DUU3tWTQy++5T49cuLw6S5xaGGJE7rZMq8wUnHYH4oEotigIBD4UpGepK2jGISVR
JTDCzisrYyeiKwwfGCFAG1K/zFeMgKVEQooHpRlDmbVXdobI5DQL5a+oQTlustcc
QnzLg/8bfnoaMChEQU2exrVwlkuB7dK+5WFD9aPZE+E9kEpXSHFFWiuDsW2Juwye
nvgNr69idqRT4IHMVyG1Qvzsg3u6KHIUU5ILmz2s3AQRo+5NspssxRzWgkqXssKc
l+BtDasu5XyitOKT5UzJnlYOFyuM69HYRZjNov+usGPtSjrfcDY5GYaLe07chnjI
4q2pBkWRrV/2Ghld54JhMzFDmDrTszyKeCv3QybvYabAII+U3bAlcnX3vjEoRxbk
rUdUx2ZrMmj7bhNLWtUOs4tvE21mgZMz2pEjWcF3P8aY5lZyjp322kfAuGwaHL/G
gRi/ZNIPv0rnyFqknA4P2toS8MCxCB2y1655rOY2Mhl8imlj5IHuk/NL0I1iutqS
0x2ntBti1MAF/zRyFaGQz7dqoHibQGsPais1Crlo4DKpTFa4ePCetEVxvv4YfEpX
RWnhEG0jvsRNlas1P83VstHdX/eLIMsJat70lI8FEjMHdWVg4b+6BC6i0Nl90ECD
UBUNO2UFLu4QnOxJnQWiDHFZKjurcpn83jNVbkG2cikloqZ9Ky5tC3C7/OhXTjyD
597WmvzBEgdqO9sT9BAVc2plihvuSPP0fMgUz8ioh4eirpLy8t5feroEiMapRfX1
7N1SwRddu1dV8dvTRAMg0OSgBpz2UXIDn0YNcp/g8rROgqPwFB9+H+CQLBTnx0lf
WLWGISUaD6glO8QRgBnpYnxC5J1gz2GaZJMZgF0hxS/1b1vi8Z2bv9MsI/Dvb0fH
o5SyWuT7VnFVL+wh8tKgIQgXRsZvW4G+hKUfGrEt2iOvY8K9HedAzo5G05IF6gie
pd39yT496HSMx0XC+Q2RW2hadh4xFrqpCMTMmpAwxlAFkR5gHAanVcR9kzhqgKiF
JtC6w2ispaTf16g6anzk7dbcwvwbvDUAVe/umu0Nj4KqBK6iQzp1O6NvDDEt5En2
1064Wfy7gow5TL2VD2F9qEcT+odiUYOzAZ6PLDk9/lecAoZUuNzG4kDZlXGNicAJ
0mrzpWQFQ+kff7/JtL/EcPZgBMcrn1gmoGDzfX7RRMl+jOhFbhxeIZyShbpCsQ47
g+IFBRzSC1Ixlw10z/F1K+dmE3xtfgatJQZD6k/TBUTFBt3w3OhRgEdwLtm4gvp0
o/g+Q9f+b4qFiG/EvcDaW7FZOijds9M5d7OQjpn4FKcwyATEYvNWDv3Awl26litq
LnY90Ijhx/7ktOy84rzulX0yjfffdoLNRncJAWBBd5+qLy05mqn0pmQttN+o6a5+
Vo/4ju6IcBW8q/HG1qRQEdjewvI0h4QSxGBy9SlGPD1gPhais70pWitjl0oYOf7W
ysfJkCQ79ta8xYSxkbYu0L+bFVpaGJxNeeRLGqcqvKBTG3h/FGDT0GlCpWJOZ7b5
Y5Z21OaV/yaK0bbioD8NM8fj1kmplbuOVu8dytiEVNqsTRtlJqI0k0CuKABsxd10
cbfM2zDeihQ2yDRcRPa28EntX56mki8ZyRwffiPLDm5FQ11CBidZkPNt+KZPBMay
dM+e7mpAeGvQ8+2pKBRsAZHDADTJDrnDmLsSBhl1nix07xY8i18S2sTC8QEZIAAP
lTbyHXDWi2ZsIptSzNpZmULJKHEbWF3RNtdVsbhMzgeH9QXHlzSn9UqJrwtNZcvf
3AZNMXbmoued7bzFlTlJvE+yi0/Pwi2K2RyGlt/PJGMQqq35gm5gXzDjrNuXzS1g
CRUAT9uMFaS1Vh6gqp8YtMW6W3NJd22iDcTxtvdoDgOZ2x6Pr8udHxOWCU5IIunZ
OZReEiq6b37YA32wFeGMO/r37N2woonGaMFy71Vjz06e985VUaXv3SAlzJ/BeZkJ
ByKtHFW2/YS5qIqTDWVXGOCy1Rt3Dydp5zV9Zuw7od3dk6y5k/c6MxMfUcOt6m5c
1GB9RRk7yMoZDNI0q0Ni9s4pq3QsSEizwugoTsI/cNg4mHgao2QVImqagZz630tF
aaDEm4Jz4gjQjr5o83MqW+hUwQIMSl0SFTFWzTdR70gAWoCoy3JAxwrxFfbRqzlw
PeqnOuRi86jtGCJMJS6rH4QKwm9qb2KoBJfAZoQcyrgc5R8JiQIBRsh3bZww/j0P
LXsvM09ZUq0QUujsZHItKNjci1US+WrsCVIVcN9IjF9jWV7adrmCz+oGJuOO4+d6
lFbkTNpPZL6HawS6DEUNyJgHuYLZ+EyJUiBHcTqJHdoXu2B81ijX/MZAzZaRmEjs
mnaNMSnGj4pMge0XAD3E+XxV/09Kzx5HSnpPB8zxiSOOcXQiYtqoZevJAXY5CM5B
90gtugOOHMjImXJnwkeUnTATapYDrzscGi2je5ws+3py+DNYX+Mrr+zSzxrgrzOF
ACiuG0StTv54UNEuZfGNuiouTqBw2A536JNRMD5nyKtLzQ65q4YXBA8F6ZGOPvPr
HcmEBR+/DR35VJj/V8tMiEnKC7b+3VRY7AJV9ACF+kAI8SOP2MqL7aAw8fHeIwAF
s1s7FAbmlvv/wQ78MwzDWgCdS9boqcMuRS8HNS2U2HTXCvOEvkBAogroBpTQERTd
RX0H+udqIZZmxgE/D0w1aITR02jjUN+rliiI0j94K7pTawGsL5rK+Jab42SRwJxv
85i3ujQjQo5YOvmAyVOQ+KnXndeJxspCsQqpfQglMbLqxTdo16e6sk++2vHTcl31
DeaFVWrRuMsJo5q0EyM3wPxtpgdrdGT7dfCU/SYTJy6y1f6Ybrmy9WgNewYsJMgx
TX6bd3R60toq92B5PS3jV/AJKfwOKzFLMSL6gT8YXHIFNUReObT/SV9KHZ+wODMK
S1AWom3gtdOMy97NeDQQPwUp3BncUTfmGHjillJRHB1fB4Y/pO8I7GhRmWG6KVvA
50Gh9bJc6ev3/lXTodxzVxzH6Fi/euZg6NyzQmZrNv0t6XA4Pb1UP7IgXgXJZ8+E
Ix0yC1hw5ZNsTTL/SWdOguREPO2Dc26uvnM8SmQZpAdVExzIPLbTowxGpumqcaRY
6yV+nlciADokqT9lP86EONLd93aoDP9Nch1y8og1RgwNbluHU72ql1qKWGxiAHJ1
Aa9AEHc/ir/v7k1PazfCCN0+yMu6a4rrM//DAKZ3b1Z3JTArNzfxYpnNJh6ieCsa
rHQQqBKoFXJoAk45RpOCZIDVP3vzR09DANybdPLyZoTYn6ZmN8AjnAVZGu8/hg1S
MOgGq4MU+DMp+FHCGR+Vo/gwujcPIDJqWRzvere0oErpw+lnFxGWk7j407FWofX0
ECfJ8kOKQwHXX3GJpFcqVxPRIaQ2AdknD13Bl6zvFGBXmW45WJPKhulrMw/m5nXT
PtxLbiUDrTNur0V7+2SrnWsYwax4bKp33ogDqfKwxGgGq2qWpgA5KaX9GNxD4Nol
8qAuVx2IqvsVzCL8+9KDgiYyXFG33NPyG+v3Eqoo7oJ5NegN2N6BZtbCbQD4se6w
fXdMmK8e6ceLoeB4VKQQnjeQuhBtRy47RfJb3ejuveCvexZQ1hjfu8k//n1O8Dua
21M2gSQifECsmb/1UsNltJVCpAuT835KRMdb8CxesqBC+ZqsVbuj8Rg79k7+ci+E
hXhqiWk78jTw+6dbW9j5KpxLRSDnNfCfBEI6CZvrFT2ciAOY3C720CbrSbkt9j6K
3kkeA4XbOq1a/zbXPolRKqXG8/zh90IvQk9QG0yv7Nlyq01ERvRxyQGvvtt5yFd6
q7LFh2tMN5gupoa53iu4fd4lvSQ92TAe9IkM0jbzmbjrgktaTo0JBcAklcZv/HNQ
no/IPlRo5gB3Ov70U5BmXMzWvVInhe/MTw80q0JrwF/UBlFuS3yFouuf7aBDHwni
AMhhYQf2tLB/y76nH6ygwW4x8CqNVsieh8Xq5M1ds/yH+TijLDYOJ1itQUeM2E5b
QJojw8AL6Xan3qOihNcqSCrElEQT6NxeAmVifty1gZoMlvRJcSfSx2CwQM1i9Ayo
vSRkeQ9if0+kpm8VQAzeioUynl+fJKbb/nZF4ChzX6N4QMCspY6JrRh8y+8gd9xO
1BHNhPGnotPCJOXRUPSuM/mxlQhKJFBiCwLL13s1b//A8yoE3PCSJbXFCcaQ61wX
UBAOSnVhP+EVE63i+yXZMF0UYANBuiMVWdlnaTPNdVy0J3LKjWxGYrtyBaaQQ9r3
H9VCD+vv6t4ka++0f09Nkv/FxOrM3AAK0HYuNs7cCRQKrIa/pxap5Qoo+k3rx9Fn
NWgEdCAdUf8+ODTPGaRfsdIUjfKFRrjjQ07I79cl1tZYZSC6LW30Ypd5xkUMaWro
XXHSPM9cj9G5Xy3GcRPhK78NPhOA5nQkbr0lmSiCppEWMU4VdilZkWoG5rVykpXI
nuICwIi67bdNKYGs6ioYc7RA1MLRnzDmeOLmiket65oe8duAZ/Bvi7l8d7IZIhfO
7P34zsehYNV5hRBKMDOhd9xEwQNyRdZpy0+HLsv0mTH472VJafCkcbl/UGkXvpXj
4L6V0yaynkQ+/+HlncBxquZe6q3Ads2qTRlDRaCoPan3Iqj2RzCY6jWqeKAPHr8A
7R5p29it3TLv225aS83vXgAQGszk/4yx22z4o0ji8IyEqefH3CpRAIwfIRLLFcQc
HbZyyyuoD6mTdPW8eD0hpor210TCdVJoNqctpmu9fUFkjs05miNWZQyZ63O0eUYT
wLWw+2gxPsm1pz23+stGwJQg2g4+y4UDhCOX5ODxwHhxjZnFQM1bo42Ll+OEF/8/
H1ou+DjkJTkIlb439btuYrmxs7Z9ZQZP/F9wc15g5CCF7fAhZr+koEli63oygZeo
kzljkLDaDOLUXBKWe4mNB/+eMnT4KC5cXU4+zz0osfKv3plhzDe8+8uJj/QNYuVj
KSlxubplpwAJw8+GGxXO/t0fu9BeQvjABR91fb6HsxIogngCmKX3GfEdI2UbX5EL
QUGG5p3Cj1YS0ds2apW8uYEDOi4nVPUULl9wzKQM4sACtENTwCmCzttEQszmnKmB
Q92hmAzBwgNMtHHXaqHHWhWSLURGzSmrY+0ntacHSVn3dlpqxP652sJuWFGAM9CY
YVuZdLMvy0a7nmAIqFeQFiM/ifzMVld26Ae3IHWrl/o8IjJWZovNfw9/n2mWegSd
38UuDxTlat76ISbUUl39QKBvzBUSq5R/6KviwJZNqBxr3rU/cRjRhyz5/OG61ahe
Z7SNtOV6jfCTAjXVFt059wLSuLB6MLtmHIKrBYGzK/hf9B3Z3qg7YvoWVp1dN8Yy
NePEsPBtsHlugKhUANfs+KJjCyQwjYt6dnd8HOShXS97eW/Mt2kagS1wc8MVXFjc
k9N7Qj1jCPQ19p2yMse6r5ceWHqavOvIYWf1ufIOuMAyi8Je7LucNXw8V0Ib8yyc
w9zNW2jPF7FVbj/l0GCeF0AAtYwzmJUrnGbiRuMiuQZQ6cVUgPnWPTFqghrM0aKj
lZVQ8BIpBMstnOO8SAVtBV+o9eKe+DlBblxsONTwAFO+vukGZL0PIvuJoYl0SqKf
MyZJ4jb5OBoctTrpWlIKDQTfIcn4ERXASQsjtKDJBuHnhBV4zNpzz52C0abMxujl
VO9O5G7Gbha9BABnGF3lcHVeV18834mNC/GD0UTMtcjmlfxMeK7YWZz+XJO+SVnB
3lTxUCTaysX45Yes6AfQYgwpmWXkAR8nOM4pS3fnMHrRAWK6u7R/X/DTAeMf37di
/JrhKeNKjw37h2e4yizoa2FJkzjwEpM7crwjsbFX1djhNwVZWOALlCh4pzwP6C7F
Yeu8O4pFV1FiuM5upn9OcUnRsp5n4de3/SqnZXqdal6mM4l/TG9+Qr586mdG60kx
XpFf2Ph2BYljNiEDKVMfSy7VD/1WZNSe9oeoFLD9TkO+g4QlzfjTUm/KjhmJzyGT
EU8VExVbAK2IUV46BV3hIdnEbFt9unt9lzciHZ34syKKuwSRo/Sd7mm414IXD92V
eoFAiK8PDW26rujDDwpTkL5jcy/egoWvSK6EmFL8+vkmNRGC/VtuVQhPYOg0pK9Z
Fej9C3EhwIF0Kwi9zx45ip2fkKcnjZFU4Gz4SDJq6+G1XCx4xn+zl2COD1SAI2E5
BzNyr3fMgcLNisQ/9HMgjurACTNaFCMb/sbZEtW+iBlg+ZYZvTSirDrvH0hqSSmp
QWzTy4gR4MGUc//zroL41ViT+3gLZiW8HqDUriKukzepkhmNt2EFLgnVQHdz6IUZ
EszWbGkJx9/wVrE8TEYBEytr6ZT1tMku5u6xe6jcIJ/ODvFobizC29tU7Q7uKBHl
hQBHWSE/LM0aDHAgHbVkmFST6fuq5lCmoSA25yy863P0eCP9DT2aQOmqHc4xAEp/
4SOSDyJEOsuEu+iw4KEjYG8yrvPfRhTPz7CNJdPH9BFf/YoQOp+VshUXnORb+8EG
GemvcE/cee34L8zf14NnWfDgtH8cn6+cm33cDxzS7bu5YMdGh3aD4wfjtVYnOOCC
dFFJwWtYjruMLl+Q5tHuW9UVadztrsyg9dx8UqfEXZQ24fI5caAHPM5jev80X+8M
QEgV2y2qzrw4QPWgEdoTNkmFW74SVBou9sHia9t5xXExs0OQayT3V0fFLDe0543m
fl0p3yvftZuqcH7ns6IAeyZ1jkIszNCmP615Tu1e3aUVan91c7xaVe3s/Orptf2X
m7qZeC/Icgezlc0C+6206+xi+9u3omeNPC39XsP5kUHcZM/QgUSHXnyS/FY2pHe5
OysWThQkFDOKcjrfMOCWSo0pQ9PmTuVdW5/q6Of1SruvdsFaD738cdzaMu5kCv/L
/1SyDorE6F7RijrRj5CT387Vgpuao2CAPWygfdu8hdAt+vBbtIMVnwdkQX7WNgwn
kSRbRljwixy709UM4og1qotW39GYlUmGEvQTsZ4odkDmNtAt2aJ/tnizPr61dEGp
2lSnos1Q61xAsnN6DwNqG0JhWbwzr44MQlpb0YZci7E7cirJzU88jvkTrjS9lksW
cz7GiQMOyy9OvHqlDplNP4H6hCI9ZycGus5GZgzLHzGDg6/UdfQ7YWVeXmuxxrTm
8QI/nzCgxNlC+OWry1kXV5Ae7Eon4xguCiPP2pT6Pfpbshz408xSvOm+Md/Hwtd9
lT/Gky9i3o/+X9RnkzxFCviJ8+oommfZBvdPk9eiz8CzdBcN7qvoZfvJkj53URPa
12xshQOMwy7MiAzrDD2mRSCSRU/54oZNfOGBZB9wQ9FFC6Sd+FEsA7m+zXJ6MnhW
exi+2czynUGrnRYbs0Z/uvV0bYQk2L6S7fhtIka63W9Huzjhs0wmACwkBMcfb5Ai
GY7jGZUOmYZOmhUCxOv8ZElmNNxod6GhLNc3899x9bmnNwC9A3WCOPr7hiGeGWY1
vNxHTPNfF5IJSX7VfDWjxxACqmORWpJh9xLvcsnUf7nrz4KCS3bmEx77sVyOng2t
7yd72T51eHPxqBtRlOZpnm+K4+QzKb6aOTX1tEj5XPXkA5pJnRcrWc2VB5bhcyLx
sv8p61C79EYvmV3BJBW6kOxBdty8jTB0k2UmAreDefjwFaGnnjcSW7uQ8KGFslQP
evaWSn7gkHy0jxjKmTJHXSZJ0CJJ+ITGm2xs1wHiKr0PejzaqaWNuE9mn+v2Kcwk
Xe80JT6KniebBuu8ibKO7IDYTy5vvI19z8d6XzMj52FVI0i7AMknpVk3X9lV9zDI
SKIqwaHNd0p1sFgcdgjP9RcxwLTAhJ/17qsyV6I9Jlvt/U1oskhhkqYgCyd9g3FZ
E9abtVQkk6KIoWV+1yRScHV81xMLfOstP3JZb4LPkI6M9GeTSppW1tEBJIXgX1uV
A190XlsHMLHoQhj96U9W1ttVST9g/dSiULiFS4D7IS9iQaE9TT/TXqWsgsUO9aPw
EnjpFVgnLGnvXAtJ6/5eC53ICBawX3SJoQSFEcb8GRXa3TxblhVXNffg6TACy2xT
+Hqk4MJmTopy9SMOKozDFykCA6sqSOWALfM7HbSgFPvAH3PhBGeNs1x0HJaPKMei
j+5D2nS6OvOYCMbrG0DFxLw8hE2KLDeCm9qlu31SSAaWkJrihMJolEtmFxGEz6AF
vxD/EWw3ADzBGVYSWhCPdRRA/puzc2EgI3LYDwcCMkuoyocY2q4BRHespjeYs95g
bghzRjdO35oxG+JSa4noOKu3N3zxiYwE6/pV7P9B2w5+u3/9uzZxyRnL0ph4tmpJ
u/fAFLe8uOey38NNcMt81ShbQQnsOXwIXDuBhcgsSXdi6WLVdUrTQMIgMRdQg5GE
+kaR8YwYJ0ZKddkCEAk/HKw4IM/WxtbVMojm7QxiSJ/pxEKNam5gCwRXieZeeVmU
J6CNPkHnMKk6jVv7w8NO7CVftjD5aXmkjVold+odQ9+ArqVAKSTQOY8IUCf6yiLI
OqikDz2ugHVxjCowjxNoPRvpn67PbWtGLE0yYh4N3yaS9qYrCIxO9/a1YUelOaPC
CueM2h5zLDcsg1I8TJ/aaggS6NcZOI7mA1HXfjehk7nkVHwdMp//WK3hPDhPOhSt
zXqLvyktiQUDkpVZOMvFJSEFPa7BPRbLpQuQirH9CKDnmCzoDBl4KXRDKBRyZDQJ
ZhUwTLt7l0p8D44YdUDh/OiDhjGTVLb8q+PIx2HRwGNYcFdm6V1lYfxh4J+Wih9S
6mMr55OpfGz5MST0IPYWd9VaBNmYTia4SOnsvpQ0PNCEzIYPepQUAZ8PeFyZNtSm
Md4knps8JpWeAY2pfk5e9Gvek5imPyYcOK1v3b9+34+uXgHhHgvELzi0zUwItQNo
86rctWK8i++sV0DCTH5MNOBAO0SuAnSRTHuhuAqEma8l9XZmNnSoqdjtxSP0orls
+XqHjtrVsEU8Gr1CZIjngmC1kD1aDL9y9sV9R5Kp5HKf4nmBOqjU4PIzX2p817bd
+ty/9DAri79+O+4nPPjKUaq1gWVk4njsZufEegeMHsD6OEZxaUPdTnbRA5fJZcO8
1eiaqras1tO07nSsgsPplUDryZ+P34sJSwdHBc3r3wkE1xPwPfiJ9o9hMW4pmyVN
bXjtNixX4JjFSzLVm79vvPl8qRve8EhgW+D3ab606C4vHWvaq0qTutn3PgISmrMQ
ma+GwzUT4qd9iDR2w3p4DLhmGJH2XW3A3bTf4lM86RAIUZS7wBVh8NvQoGH55B4N
LFPhjoHOAHxri6OTS8PZwnbbhGcm+KubXsGdO2R0gKd/nEZQrOBuhsLc0yovcDj1
H/j0LsLOjEmite8GUkOhBCbEX4BbQ6AoBnd/d88H12OH8xrUU0FjFQX8yr5G4sMa
+rPU22VRfDLmn1u1vjjG1DbLRbyPATvO8YIbyKsSp2Zm4Sys8sDfsebM1jZeLeis
b6nsoQ+pnMWgfEOG1MA7at/WcrFaaT513R18SljdSRoyRPgB/bBSC2CmxE32uXDx
+A4yjeUVsEj5/+eqqe3PP8sPzRo9KQScPErUmKjnqsd2aOglqHwX6DeB2/aW3Cx2
pwOWr8PINIZbZgQlHxX87W+85Fv5RGk/6nVFDCOXj9Fediao2vj58bwPEj7x7vnB
SrkUeTYAy7sVTN6Y0Wj98VUavT8Itj4U5oT5MXEc9/wH3EeEL3nYGjU9rZTw+zo/
vwa4SmCkAcU7fn5AxV5G2Vs/pwwhqZnw0GB3tLIKA0oOckj2QSno7e0F7/9UEHme
XcaZPDJfthxFxTPyeEkmQUuAq7fL/jmXN+u97j02QOSbjHeMKGKM8PywPuV253R+
4TXDbHhmCiSAZGajc8zgRyix+5Spb/vct8vbr7AkfgoufOfuiRvJ6KyxdjXYk/nF
ghpT+kB8Qv07C9fHNmdZfymdEkzvLCrTeurrQoKWevZxwj5xEYsMflbe4wY0bV9b
E8f93JfWdt9jxpsqgH98Rmcpik+EeqaTd8smubuxPHhlhi9JnYH3XzMu+DlXDfGe
NQH+Ehg2p+ZdOFo7uwVaVana8KUb4ycIh2FPeR+QtauQmNVkbi6P+SVjXkVBqKVB
EyXvKsjnLLwLATu46Ojh+sNdNKkldvmWYoBWJaPaPa5jd7s5JnRv7hHGSAFfBVU1
HVPxOwywxN4Ak3qYL8tWMqfwI6IZ9nDpdvOl+1ShzE/AjKhy7VqkFXXTJJ5sAgJL
Sx+j1CUMUuj+omBBRwqRBLaaBy1m3AvdAawohimCz8pqwKJ+Flr6LzqqkJVD99zj
WcjZzfAPZ/GH3iMIQCVHFxMdaG4niCjGFN8ZtSAWWkLg9fL8sMactsR7YpthJp8z
3WcSYY536eJ3bo+YIAMmNRwo0nVcHoafeONALwFzb/gVTgvjqsgC/k7eKTdXEPFV
VzRAsUdpDErBtnOSqlNOaVgJU9fcv4i9g/uaCQavXM99A7cu5UXZKU/9Prs2lf8P
szHMemu0IrgJX09bp9oU7jFRbTVW1CBuUFi3Y2pOlgARwH4CzmsHbZyRgEGaTWr4
2opAhN4eIoBoYMD+ElAmQJrsOdQljV4EdqM9mgwIl90hyLgE3ibYiLsv6SIY5tMF
ovEWpSO5rtMTWPtdOynfSDbfpLbgGw8SmhDAvERypqShotZkE82QrYIeCZaLCrhM
3AsPBWaXvp/gu7yua0rk93h/h50X8sX2ZWEmN2DmZdwT2EMvHm5Z21VLsRrNRdEa
58G+8XGX0bFUNzeOCy1j0iKdaVUvFtPH53fLcWPzwEcfcTV1skjR+Y7Vri9tdBH/
FqhOxywihSa66ObCh4foWaghKmv5sTMYIh0/LQAFIuKg2xo8ebrBOLIdXPVpmcfh
2Urc1b3qVLhxsCCxeJMhrXvn3zCz2RGvkQc5RS5IYi3G4xU654bxKvkjHQjaXE4+
Yr3Q6ObkhMjcbdiJw1gZkJDtxWIuACkGh5ItzWgHPFB1dPXvB4iKfYaVgDj6/f66
HzkoOs6XLLF16+dLwfmWt+kyGRy/+IzmDCT2BISpQjmAxtBy1pwbhcZx0j3aj3d3
6JfdwKDOqu3vH29/wGTeZmyUEBjb9PXGtvoeBggMC+nTsCDDwWJJWl9/xw5J4Qea
rl5X6CEfzLgf1grfmUI7+YcHPlwNF3ZAXUBjquFXklVje7pOA7V2BSlKeM/n/a48
J3yGWISqK9Hqm+7xtWViCHPcTMxK0gje0kIbmDTdFZzaIsjQrMNJ+bfyfWFVK5Y1
WpoBmLbmdIzKtmaopiazAvroueZ20RQ4Z8SoctRaXykYVX/TMy1HuY9wW7PkrUQb
B4HOf4RtceBHUgBwnr7ag8AUJnsAMQ4MHwiD2Wnbty6xGrrZ5TOOfipGFJyjwNzh
m1GF2mT8JEV/wfvlKe4wEnJuCBQy8VVemmrTVLYG8fC86FdgT9jriZRfqh/OHaFa
x94kNuIDfw2Pzcod8H37fFyn9o3DLFR7H0/ySWB0ivTykkW+IEZYrQoP0AQS7LyZ
d5L0KlpYAKJqix2t+ZKAKCJsR9353HznW4SEu+2UcvKfY56hMAQp2ZE6xP/WchcI
cDK5o2pqQJ4lRWeFWeHGIPLc7jte8HUEaCdi86q2WcjPSiMI8EliPx2+v3Rf6bX2
gJbbWVXGJmbL4I+ONolYeHM4bdmOG4nrGq9RY0cTcIBq+LTXAHUkQVCwjwSO3ybD
+H3yAvmoK1tsTQ85ELpqDJ8997ganHWRirFj/Mat10QLmGrvgPks2rIK+rEQcaiV
WH58V2gL7jmsyFM55s0Q8+30f4Zt9lpf62UtZdVBLJmnVyAy7TJZ5ByRKq4+FREI
82q+rsPSQttS9mlShrJSSL5GY0+uVUnk3ckRdCj7mf1WlEWmOVLk7TAUr1g4M0mA
4D52TbKc/fJnWFm6WY2BtI7v+4wdFL3Uz0hnpfTWDrE0w+UaP9E0qoHbY9B5gpY+
NlYjQC0h0kiMSVQv6yF2TXYH6V7kmOsGVEN3ZNRfTjqAKjTsH0+29EgR+nYNRj1r
03cjwsofNDFNq/fbSAE1WbD1NdaVCcQCGSvJVQftZVm1TmVmJYtdfvI1HCsRZ+/n
sjQvQob+cwdD92dteSCxuvqZdoDlZVdNjeqZrO5nMiRYbZ3BLse0OSEFUw46Fvjh
C37rUGUGzvy1I8weQpn83OBWiyI4r4Do4gSiCNJLWhuv2VavvpnuuEkP1yjPNcOx
BBESVx/1OJP7oW8KV0KAmHZPM7Zxe9ekvH0XzKJfarsbLIYU2XSyKSSZuB+M1g8x
SBsx6cPOp1zZV61/A6zDB8Ah0kAA8atuTQe3XaiEs/PkdabSLL2iztvtu/ETK9KZ
LUMu65xBJXnmffokgN+RjeWcAptzA+kNHsCJfe/KXLx1+4VhcFvt1XduFZT8OHYp
vLL5Q8UYo9L/z5eSNk1sOuLtxaHOlB7uxgfVOmmmDxWjM9K4SXCjQa+eJtG49OjE
Ek4rT6By2+MGMzH7tzzF/YGd8ptKRO7BwyaiOqaHdZR78k/vnBqVN25ZCdvqq/KA
K29d+zNiGLZ2Fuw0MGbOVIHpOj+3fgvNdCv8QDKd0kU3T6e6wyZkgAuxWlfPrN7g
897HgqmSsnasbzXVSs0EWhsm/XFmp2NupnIex1RvZAkpVSlXrmRy/fYzNe50JIpb
wdwAJU9AX+lWAqN3YdEkLucsKHLyUo/h+3gtEugUYpIfYXpHWRF69cbJGM5Nbpsx
esizTEFJaH+qChkAOmF4846CJAV+EsI7UMlYO23Z9+jLpBCWLAdRs4vIRw5sHDSf
660CDeYy5X6XhulTm7QGLi42cEX5MCXnd6V6t3gySyQHW7Mz2SjLqqMebJ1wF3kb
WQE0Dk0rBZT7sQFqQowgtLh+fcaLjKkxq0uCa/IHsWn9JjEE/xHaEyMSCLWwaFTa
9Skh0CPy082xE5Lj4bfitZAN7hFC3B45VipilwcCEZcSIXNTNbdzXDzbD/yRo+bh
nXXmkQKJLXrBcctzPVoAsPsW5aZXmcqlbJRsjhWur/WOwQSjrzBXH0979miBJoPf
F+rxS7tKEQicXdrKQNB+w96iuzdKgpOIk5AWWGCN68/sTZ4VYr0roVjNXa0SEWFf
dgckFHJGdysNf02ekD/GQyh7vASa5ENIvR8rDXDp4A3rtF/qJZSXETdn1yzUw4/s
zB9T0laENI6CNKsDIwPAoBXDyaViq4osUch5VQN5piOX3pB7JJmPC1MU7/RCbMLO
6iqyXo8GcMtPJzpJgPW2MbKDjepG9uKoBhuibrHiPrR9v9vEy9eemyDolUQd+i7g
U0oxXZ/9Wb/ZzAm53s/pO4sSuDJmBkSG2JjCILIZKVQsW5wa2RgcFeVbNq3IBKJu
mALMEOzOI8tJgPJ46xZLGZGqqPjJliqSu8PQZSQ8OxZQblTwmvhWWRlMBMLgY4bu
zjBskBCCNvVNnhhlWVlx7nwIP3EpPESl5SByQp19R0NtH9SPttO0oh/x2IUVHGcQ
nluynA2T7GLvP9J5DhGkUevBTEQe1kyUdGiXJ4gpJhuLmjp0+hff/AGi5zh1WMOK
cFtNYJ7bCq5ibL3J20VP/3ILDnmnTLV+HYh1v7oXKImzk/4yUgZAiGs00AtWPYFv
NC/Dobb7t53eWzyjA+OLwRb8CCqPMlYu/+uDWB2sRKRKhec7Cpl2/Hg7bjYmp/vz
YIOxTYVPyZbA7r7/5xQsdZsF6gvd5X7MlGkdvXdCJSmdbOkiDkJERJ9iDL2+7XT5
C9KqnnjE/6DayHz34CI8Wa9i7ot9cje7/gvFBmn08wHFVlfBlZfCGrBl4JNUmUpL
tmohOYPxY5M2vDGP809F6V8WmNcgCAB9WfxeXcj609PJTS9hyYZuICkQXKI/d2Yz
h/dpLYj3jHnXCQA3AEupnDP62jJDL+NtCpdgLGb/WcKOOR1eC9TklGaCr/2RhH9P
8vWpkWLplKBH8laJouNBS9oPP3qYnWAD3Uw9jfCHvDziLybFg2vCCvC45Nqqr35a
E4GjnsE9ldJmS3xP42sNUPNv+4AohDljy4oleDqlAaoZhuZw1yybm4efromKG/ro
MwPPzQ1GI31rL60DexenSxVahvnipCCj2ZrHuw5v4fnBGvk3R+pHMnaw8ZxrHDl4
ohsh3FLG262TCnpdnUu2IB8poZCIXiN0H2fcxeqq3wFHQBKFQoR+xhv04fRANVEO
WTPRn3qYuNnQkziLMNvAyvgza4eSH2MyPZkWDt4At7Zud/0c9aktvQxQOEKBJj1y
vp4cdSbgDO0CuyzyO48KZ7C4d4SpqSwMydyNqlf/Td9XTnbsRTqya+AF4LwF13It
2SL4nBH7gDNu9tVjlGLTZ25BQhQvzwRGEw7Nmsmz2edjDibuY89dtauVJ7rvZ4qM
O4PWGhVslQBsC14m2/DK/Ud5lXrd5fnTTk+wILG7ivCTaYZpuQEXzg0P1Qh1gSu9
K++DuH3ZlNkIR2nhMMnvcRK+ZJIxEntTrfk0yPuzokmiQom6P//x74BJ0bt+e7kR
DOTppL6k59UGZ3fBv7AUF1OJAUxn4jVmjfCKJpFK3BlH1NqVlAQlkdxoEJaD/ERj
+nzqMYTLgM1+PRftIp1QI/bSbzic4OCO8lXZ3aLUnjR8E3cvLcyN2X9Lnp2uXrM2
1oPFjgjMT5F81AWUeN8l9fEuSssinqfz1K3+hifq+wLfAYVW5aO7h07xuKupZUmy
tBi29/tNubj3wdlQRiGay8iJ3CiK7Q9o4qCb4wAcO1EEEBo6ISewhSeWDN77CYoW
1K88TWJqoxmPZrp4v7gui5XttuaRnG2CDxGMw4yqxYGrbcHHW7/Ez5ByeyBc1HA7
kYgTkkCkt3u/sL3gVE9h33suc9r30rSKlXP2+/vFYiVzcuKFg5sj03x9ICJ36DwA
6xnvbDxrZ5u36pq8y8H4Q9BqnUpPkQN0bWiexgeplrUtqBNflauVZTDROfJUgEcg
t9So5dp2leC62kPIKFF+qt6NEdhb/MrtFZ0b24kr97L3f2tZu3IXqUWkBIvwJ7Ct
qvcWybDYjiH6J3ZPrBUTBjWzf1kKDKG7sZJzCDP/m1KmhgaFZ17ty5QQPsb+tDWr
RFrcGnei7hQQHn1rf18D8utDh430yPCHOwTl0IXK4iKf6GJUMW+jtV7uu3ar0BBd
MO9OARlM7LDA9MdEnbxiOEtlLX9C+BI06y0yapMXFlJqMOpDAW/tA/gkmsI7+Toy
sH0vW1+g16IkMogCWwDhxp8SZlcnfB9TmRJFjLhqTVHvyPtSmkiU0zGhGGID/JKO
RelzDBz4yajnoefhnY5obepyznPC9i7SXckk2DH1gn2PVYQprct7W5rCBi95HYP9
RAs2SVEIHx1HHWE5uuuzWe54PNzZF18Og5I/N81jPoYWp2sr4KHhlZTLZDc5cYdf
aFXq18WVy4jUI6aV9gCNxEAXC/MVZKqgOmM2/hRWibiZPPEIbTRMhMlCRFygCqpA
tpA9PygU8QdMKQcndJpHkGHQtg/KiaQyrljfLWU/qRB/Ks0grVAW9lUt+AOABDes
oFIEoF6r43QbesOKdjY8DPEDYV1bu294Kp4vr3OFpoZ61ygoDZhSWgXvH8J4jMKO
IJGVbJS4lwiVQMer0mqN8p1x4ji5nzwwavKS84PZFFsPXJAokOO9bETDec/oZhJC
att7uY+Tat0c92FJ5bNUoKBTMEEhZDmJo/W6/6A9cE3NUNIgv35HDscWLliuoQ2O
ry/yVEjpxVwpm0U4psGcm0+0rium7iwpsTC+/IUC9it/MMJ85uqIan6dbrGkcRbt
bz24HdfujFy50Sdfsuatx6wM0+ijsg78OdW4Ph0oa/vv/ZeRlJ60bQnW9n/pVD5g
kFXd32mEjOZP0i9Qkvx6ls0VonLmLD6K43twXOuKTBcJHdovMkbEiOuvM/5hDC2q
OccgZPxqewy9u588gF3ol/Mb/aZHumxJwEBeF0IuWUvy9X13LgZIg8WpprZe1SKO
mS40Bfm63YWf32k49tZ0AgmO34Xe7RWrk+Bm0xcV8hFpuHyijfFWkyFi49O1WTHg
mVP2hbllMoKKbkuriqQqzzWtjD98xu9MK/nk23uvKFfwsQDaMDB0ScxyspAmA+AH
wHceAEh22EXNxuv7xTCG2xGHI1x/GGh63b4TYOmzOLd5U9Ibgz7t7vgTtOBaNTaw
MJIXF6+VZwY9R3lvhIib7GCusL5B/PUo/RHzr8fdT0QSZj2k5C6mutD0gutHfSSa
NdaSM7uIJwh9t0uUh+PuFEoq/OfGpdoJGK3RhvtFGNVFJ1G+gAl8dtbcKxZ9lMnz
lHtn4R/AApwT1efyeUNOAc0D8US37Nri8vTr9m6S/GYQlP16GKT3cj+TsqzqfHqS
umD026ONcpIYRDkZKyjCYEDc/+cXVX/YjFO/WKcmdI1zRlStmZVGK2ELZPUz8sQh
0857L5wlSh1scay1bN9tX+C67WFajnfGKLZJbX/zXPRseLxeYem/b7aZP3NVs5d6
9eFjffzlk9SDCQJClM3H/d5EhQiZk6VIZ03OaEt0ck/MK/uVHhdkr4m3pwMDMCbz
DYXG1iGtp9/sN8l6wd4Tpw35gKpd4EHx64wXOFigKMTglFriN5e7PS23CWlFDY51
7TTJqICCNFEcbeHS4FmREC+fbgNHZzPIC+s2i/xjuzTmbFq5ZRtN1LcBGRNVWmDg
3gaxiNth6ghQ3NQQD6pt+28ijIOafaP32wq2voijMOD8at3nPGS9FPULkPnLTp94
SQDyiruXXAGhM1TMq4BJbNfZpAsVO05xnTAfz3S+KjwoLv08qULqP98Cx2tfOgIy
7oVwtEDFpWQfiJkeQyze8magDw0M3Vey4Ve2uM6WJjEqrXun7ia9cZaNVunFWbOA
oZpWPjG+mO7VS7KiwFr66keNtd7N5x38fz23JzMaD1o/oWAK95/P1dEKklQxr4F1
uLrISS6MdLfkxudBrzGNcF3YXfbxDbeJbUzNYOld0SY4NUxuJkbGzg+CpYx26EGh
BgdbolzhTL8xsmEBQ55DUmrxKkpgkG7INkC5b2FogN4vstBgRnqRzB07bF8cs7VW
Ie9D3OyViuRX2yZWlrz1sARx03nC1UzAG72F5r9gBgqZReodwSj+IWDwoeaZHVDq
x6dhWdxI3wl3yRKDwricACPNTjzzYKO1KhbbVw78kZP8n9t1yNzt6iYdyz3SVfRm
qs/qdyb4Fh4uQZvUFb4QEW+z0EPIPKswUvPFOwDH9aphxyizh43E3v50o9wXy5sq
hnh5hsNbQqkaiT5+tpOv6nNZ2iq6lNStm/VzjRppAH0Y+FiIAvoMVj8rhxEbxKtQ
3cGSesRWOiHSPCe0JHON9qHzrYzLes1gKeOwS2cDa/CCcauCYt+LIQTD3aR+cJ22
xskyH8fyt6VYmCf/bTaanPS08MrE4xqpn8Js//AHKAdY50x8zAZrkAtHhc9PmDAz
TuRvbYBCXkoMfcFLDRqSZORbX0NzgaMshFLhdHZj7AH7cwF399GZOsMuLgm/6XPa
3lsv7HUKcDHiCVaGDdNVt9grB2wqwNbjjTNNvmIUp4CZeczg2m/1X2QQfApR7B5q
zlnYi9iYkEJhKhl1ImUX/9KCsob3z84eSqjShdrpjAmRlG4qX/iqzxhFs1c1glPR
KhsFHhdCkHiWzMZcHILuU5JVH2qzW54chqmomt7/Iy0W79PEf2dTwGfvPUad+uAP
IeUOJTFzPmUn1bdQEownu8JOuuB+1msAZhiYbqMbx0a+UhHwDj1ONoJV5kcr//dI
TjjHafUdG5vDjtBtK1M6k9xmjWoLV7mi4Tq6yGsqZJq2lZOw4Rr1hiVeg+elLirV
V7ExOtCcFKJ4qPK2ZOecv0Nzvd3VSXOTp/T3V/UnQP5L/So+Xm81t1Hk+ilYkhcC
W7+9u42igzra+mUFtgJOhJwYDbsQrC15Gw3Y4xgJR+eAX7zMp0Njg66FlnIFfabM
h2c2OjHSwsRCO/fPTJtPI9oUcTlsF1laEtlQqYwQoCBoWhzF3B47QSRLua2Ik56J
sD7/FPjxEgbofagUWEz/GrdZvTyRKFQZq6iklU/DdOWmNXuRrK9vZC65cd65b/Kq
Cz7vwkSGzqd+rJ8tq9OapH9orbM92FlTT5BpVvJktr41GQNlP8UL5mb87KVhDL3/
r+NmfqxpH+DFvBbfaORB2Vfv/1+A9l4lCxW1JU76w1fxANVz/dO35ilh3eS3c3Wf
TkzpNeRUI4Mn74Vy3vDTx4vSN+mA8LxBqxh5m++axvtXTm4RRcQigC9OHBp25W81
ljkjub1AESlZxaNUGmDN8SWpIm5l2lCAiZnGDFM6GVvZwH7uIvZ92WOnxk4im13Y
ouR0T3uKbG0l3BvqozQt9nVU2ziaD/u7rvBgDpLnM0ryQFKcKNzItzo+1uDDgrC8
nYfLH35W8RHPwh/szPUOq+0ECOo4LT5xXssUiN3f/TZB5ChdlF1nJdRF33samyey
Y+TIY+6RDtPkeOoDPtLa/GAXdxhx+mKAq4TM6Gqln8Am91xHIp7h8HiPkVlljNJ/
/32PwfiNXtsaiY/fcE06eX1x9rlIaZUKm1CBnBHPewV/Hk03gIVBH3w4DgalEV4x
mQ2Isjvg+KUCN+Dci9zpb72Bvh82FenkxgBX1U+g2g3AXonfP7nlCI+H/NW3Epjp
ABwHdV4MyZKcZvDFuDS0SuLmYlqX2deSb24Wu31lfT0Fto6Ezx4zNfZ63MszDs0X
oRXpSx5t6mACUGtkxa5dnl5RycCNgDRsU1LICjy2PnaW1HYBqKN+qcKyWg+X5JLj
YVvO/JqjNhyvBW8BRIfjEZPbpyKZJ6hJzDGXG8KBlrMQlzl3JCpG42Szp9fuWO4X
cBci40zd9UWpOsaWBlke4AG7qN3HEYP0e6mJohZNVTmbK3Jf/knSSl1SDJlnoEFm
dm99gha3tmA00u5uICRGyd+wQvBUdyJ/OArG3V8T9GfOn7oVJF6DYtZqDc71vSxN
//akIgCCbMGtEZREIEtfxZKiX2SPeHnRHfqkF2FeD73BbpV0+tSh8u+u1ipvl4jj
gZyZ5GjP46Mtx79reNioGvjVCFOFKtHRNpOl/JP4TBHgZbwi3ym3mg5z1MIlzGL5
Zh+B4mVBGPr6KTZ+Ka7AICYxKC1GKbCNUObg9Y5RjyXeUYJYt240iC4E8w2z9PGB
7sHeXmo0AgkAEixAsG9l2NS51Uy21NE5BMTQhXZd7yqr+Oks6SyoEB1GPta+TcMz
Sy7hqoraePM6m3bRPTbkMd4him6FYgoBdCt8ywyYG6Nw0TPTro5Kb4lCLUS92sf6
+nBqOTyRcrQaooLi3Pyle5JVKyGjA9lEWAaL6WDxjXYc52t7zK9ZPw9xRxzlenwR
gJdRsIn4D8SCJsc/GDgKed96fnV392uK7Y7cFmmHcbShpIgVT7eU2XhpHVVujvCt
PYvCvzsr+71zZSFLs4GfTXPsU8rj4txZKmCiblSqWw2Zl52BS5DTBTKAHPv6jxqZ
BTHWJX5q5cgVO5Urjt7Z87IJ41Oy5ZjRnU5YsxfA1zlof45GxAtw7QocC/bf1Ju3
+NjH+avAcvZiqBEidiXd1od4x5CD5rjNGfFWiu+JlYtwHZ0ZS6PlWvVfwEwJX+97
ao8UyDRKpM8r8EDS78yoNh5oVDQXMHteUlgEDcm2z30rQsIGIzwGcQ5bCc5fRUgg
BwdaRSPnxyirsZgE9t1I7dMJCXY0zJhNrY9Eg4ax3RHEkT9p8CNcDAbUhb4jCpcW
yyP2schPZjyrJUn3dRg6q4BhQkmbEe7gQiafHNwzvIj3X6gegYpy/diWZfmT2LKW
Giroj3842muDBL/zKOON2pD/EXAR1z1WqTSUEm739jkYXGH1uqQ144OdYx0pIKYr
96mQCy1FX7ocB38jutxoy+XW2KzoJU0lO8TsT8peUC7XGcedgI55GL7bwlLh4Pti
QIChYtZcKgyIGDy9kBf9Gm1xt9kRR+t8m6Np83zYz+4haTBjllEPQit6CZiGVWe8
EOucFHK/KiFx0yH52rMtsQdxO4n4v8M8MTzQ0Tf82iw0wkqk3UHdl1dExNVQ0xpk
H/P++JAKI7GJmike7SgdEjZRg9JxkpHiXfDZKNqA1PvsWW9GO5oL8wW0T+rNTB/0
174RjZhKAbFgQQEEA6Z6oynVhP+pkDGL+qMLb+dtG98PJodFjMXoCp51B0UwpMaM
ew4Jz187A0owvAco8jV/VUqjGWpt9Mfc/h2BGaB/i5Ly16uPQi+FJvYTGhDITmSa
9CxEzTNLytgTDgKrcGuSEIgLHOCOjW2tbpiLWZmagRVtr2zWRxKYkCzhR1WdWAsq
36/m3hyG2h5sWx+LgNyqpX2j90EcaTEdsNslDEHLWX6m/Sz18yc7d/5LvK0KWZ2C
QM5ePr/Ojlj7emqrQh2RK0TaKUVml4oZ9pdwWo/bREdq1SQBOn8TDlmX5suQCFEc
Bl5Kz5GQf1gnKIe7/ZFcuuzCAmIoe9z3/9+U7yJd5WmuT9acmigEmB/F333BcXOk
zlOLH6X/oOY/FsHtSuEANZsBqvKO8FSWqhYqTZPkE2yCO5CQXY0Gzvx4jElrpru/
l2i7RvVftnMyq8t0HpkLZz6/7EKuFksL3to57SK2M4ixmvJf+NYAXgolVqN11Obv
KIpp8iqsaiLLtLGjee4ODG+ljNCayfhIkjM/16+BDJH4wNJFYkgnw81b5rIXmwnb
npUgd504tkA52bkNZnvfimbuVPJFIB/BfWwuF6XPz6vdd59LGEHhHHbPynFETAcm
DSus9DxKGGHBZIogR7qz7Fbrv9G69RW8f7n9NYJrfdzq0KE+buW4ogOTWM9lPaC3
vLhRSiSIMCsn63zOwd0INQLWw2qEwOxpOWWGjzltuI9VIjxBq4UNj8uicwyWCP6n
OYpoBPurhGhkwy0BnmO0QksCyW6T5r5B+RsttP6zKyV3W/QEj99PVOTIwt+XWKt+
6tZITIfsjr3lmcRIiRh3ffvfTQxvqw/cvnzpoSTiG5WvzLY2iNnUcabYHypb2uYs
zauGEoigImKrIrMpDno0pf8cI4ij6d+9TyEVGjYR5gpOr6/BcjicQ52TxZLQ8h5x
6H7HrXK1AEflx4Vbvsv3paM1rmbWbKHsPdPdWWbsGz6BafEQQn2PkHqKNDPqQ0na
cm5/lje2zB5WoPMooVK6gD8X1rqecVb+cHyBB8yspHSCD7ZNEqLq9018OVhflwwE
9E/ET/bK8I/QnBvYiffPrLAQTaXsMqzKBj14h/50jUUaS6y2DStOI9NuPWOtvXSf
nepsBFEymkfTxTUFIfwzLVr7ehuKI5U9dEwp27T3ExtKm3AdQS/9VskKIGezKUn9
jw6CXByricvgjOi6OcnBf1gWwuNSq5IgxYTTs7VUKvtsJspqMuvjeJsnym6e7iDR
hh+LCoNGlRjsKFRoFbFA5N9ECUHM1aM3FWjsme89OUFeFMFGliGttT26/Jq6p3JR
MlvVJV0DWhI76ze5LlKLK0IoIECsBlSybnhUrxQ7ZZ1Q/SgjyeHA6GsN9r18kd3l
v93xGhKSKmElwRdnmHkQzh6xAEXPJco5OsTgVpgdx3Kofx4+N37KCBO13oLkOB7I
dcE6/S1DxoD8PC+VenlwfL/RTNAJ18dWGFqwCeIrBRs4hOf8b8IFwc1gPAMWJA0C
vtF71Hct4vtndXiORaZnu9Q/+3JK0FeeN6VMJsfcu1A5yoKZhp6Z7k/d7QZc/hNT
BtBq8YGUHQyOUoKj0Maq3cL7SZiBS7j/i29FSuYg9K2nCtwOIP74ImYQYV5yrBjL
e8Nf984AzkVFhvWGc3yv9m57tY30zb5ZhZh7w43EfMhYdWRZpGWu+QMrFtLz2OEf
wiXK/8ydPKCLAvn4wiOu22JI/RrMC2aMUU1aXkZFQ5koaNJbK7YBhsA5b160TATf
uvxQdkubkqdc0jTR2b+2yKUr6enVvpExp6XRvMFvUbUFlrpSs3j2p3PFZ1Y3bGuQ
WAcP7BPowHfHWkqSE891Qd6Ut5MmlrAGCEYYUc7g6VQKB3qovpXc/WXqaxJBYdJy
ZBUSIlU7xTuiFy5/BEXVfaGB69dgnz+sZ8bj1v4UTZEqBhN7H+g/st3CnyDh97uw
VMZKH1RarNQ31TZz9kTjESwmHXaJDnSw698ZKpj53h1bLzKcQqHgiY4fS9e6SJbD
CBWHTpOqhraVopxwRSghMIh2EJDd5dVgGgzY68KWA7yYjYRC638NCWq9t+IbJT73
25G9OwjOzZkEzYwHDGmgyRvhmXbgrJ50lc/6Pg37RbZJymYnc1ZEBBwgiChlRAVv
cESvfASnjN0cgm5SmRic5l8Jyu6IfxA+EI2uVWwgEqmxONPye5HeOOVGcDD4uyv7
3NlAAAvtAKaVXu8TlqOKzs4ur2ICn+jRHxx98EHHYvDLF1t/gk3zvkz59+kmZ7de
yt1MXOz1i/hg5wszSMfH54k/8LUBkKKBAE4S3g3YcKs0sLxaf61n32foO2wlx22h
FZKa0nLtn3bdGkFi020qPA5jDzzRtBKPtMZ8NbNJS/XFEqGqTTl/roJgxa+4bvMj
QeKeK6vwVIfrbOMu/ikcVbFw5V1w5OTOd9xcdr/5NToa3Zppc6tN1clXFeerwuIs
P/3aplbuRS0yhDvZfTXgYsBHwKBPxK11hOzFrxaMSgIZJ6hi4BTgrCgmOCLojrn5
KWE5TWzmL4O/Jxv7IwOiFv47ZheK00Hnbs9dt8oLWGzw9gG4zBrtNVXZnzSvRESz
GkBM6P8tU58T4xFdC+aixVfRfvEOE7f/IZJInpCmsChQIEkIG/ydEh7aRAX9zDRl
wQ4BB/XhYZmhcfXixjj+BKA0mgQXwnENcN5RXCQMebavmk2GC93qhcUHj3U5qlvc
OyDfxJEcmHbotYtr+AatEWmClLLiZPgdVyxjK7a058++3og9siMRRmR/GGOCh0Bc
zLuAzjwAqEoJhbyzoMFWV2mUu4PFWn+DNMYXOfuajGW9CqyxQp9eLXYVsb4SMWzL
cXgbvvMjTD0+HGfUYUHS01NkoWgYLDMXcqLQuo14GceLiVxoAsc0Gf7a3rdJ0c3w
J8hCmEGVRUE1tm4aP4+hiZZIkvAOkt//JVftEtPPJHyiwlQzEE8bVaHJpDP0Cl+u
hYAlqHn5OyirXj4I9gQPt8MFLaI7F+9W5LGBiYc1xJYxSt6Giy5yFMc3TrxK0mKz
68psLAcIcQ+HSA8ahm/xl5o90KPsv66j3gM9Y8Nmya7XP24IIAzxafCQqwgKniR1
2PW4+LgFC1iGKJD8PGRhPlOqHvE0y9nDe/D5xKdSOPeXkg0VQ+VmkRKVsREZzv5P
72G7ejUTEPZtL/REN/PILNFfmH9znvc4tr1OzEK5yF6urn2+cITIFVhGugPq0Qfs
JfByS/ebUKrbJmG6a9vPf4DdYS7lsMa+idv3XhNvINMcTJh02z7fJU5eWlA0XQdS
foEVxpspA1lZnbsonwuWBjw0fko6XwjoVRU0F0us30/WK3aP2ijip7wnP42Fvv3t
5LFmj1xVof63SooBVP+InpGJ1Ppq2wdKybJr0uAt/1IR8Pphc0JeTq2jcK/XVfjQ
E7ZVobroU2CDwHjXynr3J21XBbRhu9UVmiJs1lnjOoKEuUepDcKiQKNjL7wEXKUS
ZFx1prb9wy7en40GLxRxXiGMqzbenQfiG6lcxl68mWKRILlECvxRv5idGz7mUr2M
WMlR7CnaGisMW8hcT4yk1/yiQIPo3kxmWxFoH3cLqM2PkTLcssxZ35yUElhEFUvJ
K5O6Uup7QAEDKFBudvyIj61ijYFf1FLTNXDxYeBNCMZtw14RJpIbVomT/bGacJwN
NJWXtvR4Q7sc9AFuaJI98EkEcwmqDAZgJP/Dfm28omBZMoflt34yrjxfi7+485qe
XKYoShpb17hrfvVm+RzLU+/QrJ+vDmZRMSANUJRaEXga0ucJH0v/jjFVvJ5qNugX
Peduk3rF/VyRgKDplYSUiux1LtUMEKe6RjwDrJVAV1oodQm+rzs8kwxlhwWzZqvE
nr7ZUPorXfMMSnftiYfOBEnEtJowWpoO3bgmtYtJxTCD0f+uwT/sln3+cijpNMgT
yK769+mFaaSnuSbhzoqi/3utQUoGqWAmoA6KmRRVlFpZCHRPAjXhraj8qpHC2fDE
v75bFB+qrNeuMAYbQqP1CFiW/wiwuToKzYzWbaUk//pJg7K8l8oCQaGSdkTJSvQm
uErS3t0scapPyvtHKRcSXAbL4vHJA7zfvP0zkEVD3Socp5ttUWMAQK4Pi/BVI5mR
JX5Dv0O8loMNC4Fn2TvUbv3nV5s2q/6X3AR0Y5g0lPkv/oCzRWF4PNadBBPp9v3r
It3EtVKYkUObgzw7g0sOKrWXWaZPUQBp0zz6f7PyT2uIaUXoHZG9za8GXDPsotck
zggZccAFkPb0avKTNlDandIB4vXnOOMI1gekUxTlz9wqMUPPM3KBS+nkZCbi+cDH
t39y+W/H312SPFb2TqrNLmK92zQU0gMl0qhDtlyEjoVoNn3PKbi4U2T7MmyQHBTl
fIkuTF+lVl2K52fGrqR+YInQ7I+8c8xlRawhn4rSZ7Dxo2qFaqa+tIEt/a3MJ/rK
CFcxcLk3sJ4jkHLN5dtqStrCm0Le8NeMxRJTzxRqb6nu2L+8MZCa2UM8dR1vLqsj
2kx+m6x8k5ihDop4xEFUq0CSfwpl8e3MAlhZdQbE2BktLYkix7TAaq2N+eROpTak
aM4ISsb6mwa47svRL3D0pqFnaaVAvXuX4YXCQZpiaRUj30ggRgXhr3bv/7cOY04K
uMPHOVL9hYXRb0o5mSphj0Mmgrv0wHf1coUvNa9geTcrb1z4mjivoTGtWXudGkfo
LvSLIEPuSwVWYZ6hvskWgpIytJXXsTigZbDmblBe0pYJXSuuSEZVEZlpCiVjdUrA
V1MAFruOl0K09KHvt0bmAHFDYGNXMnq6bShEwjQYIrB5bA36KPG2EzEp7qfbm9Ey
Aic4ljZJ+eBeWrlPAODLMWgAmKPVY5e+tuETkylms4Lz8vwljHGPGXu5wT9p37VO
oOewuv+8TXUaB+wVkDg3/i5fRIH2Onk4t/h2ZMFf0RZgxeT79nMWCONWo5fIn5xk
UQZ0mURbX/1etlt3GdxPDKsT7L4FrbHx/cTs1LfrCXpPC+BQvrlNxOgznBLlLk3R
1goSZbqi1GpEb1e9eBpbRK4CJItZsOFV54JWlgKilU0IzMQxLVv7LAKQ2tfzU5wb
NEpjtqp4kU3o3cTdf4iAoRM+rXV0sPWcQQyzE0OHmHSKJGxXSGgca6mu1CzRSJAX
rm/q4ZKLH9nlKP065fWTS9LBarramCurzxlwvxvA4H2+z8ooF9pFyTmsD+QbcRwb
8WxsDkwBlbFWMvupaPhgcQtlRiEpzSEETrZhieArxqFbku+mppw7cEeuhRTN0BLD
mhzAaKfoOd7qzVrXZdyBfEAG2joloyoDWeovCITf2ciW302mjEvoRaA9HJb9knll
JXriPb663oVxeVX36Lh+4T+J4GrRgLZNVg0ucHpyAR4/16snwJdwwreeVHdw8h3q
q+oPv54TUJaTtt/xanVbkIP/P152R7TUHaedwJvI/Hbooy1YF16GAK3Myz9v+6RX
aJUZO3q9PMcxBNBdInfBPx8zk2xs9DM7cYm6XaKEBNkCEojtPJPltDxBMnyTTTst
dg05RTDsklv9SKualfbqldWafkolO2AHcAM+H0kWrruTZ99xqp+swMn0REbr4u1R
7e5DVXrSDh4mZVLmCcjF6uqAaaVUu2Mg3igBV3K5dK8XI4K9U8yYoEwoSY/b8jaL
eLw185w/pbizpKdlIepuWUBJzOSrngDAy0XfRFFturOl/El2HcDUFSpuDY1g1mNR
v9yLSzS80Sw/WiBOP+t0fTVyicBRPRy/Jh49vdisGQpgMvbi6PaBmLBm2pMRpfWz
hj+WhlrVgKGH7RLFlcdb5wxFhydaoAyJlAQJH1xK7HJpa4i1wnx1i8oLHiz8RTy1
HUe2vb2/HSCIGI60wygW1AGql5acFNy5nvIfHMoz14e83gbCPlgNFrfmxp3iwKnY
q8Mi5BwmeU8iA+3L772h0Vb0spxFEuNhLmM91TtN0wTzcJRxpEgxmntHqLqC3QAX
y1omx7TfXoVRpqUGjHalJ5rtz7UaHpivvNaqU/g8e6/C1SUgvFr3YVMOZ+JMKnbw
Fk6WbL3HPvljA/Z8Z/EquPZ4hfNoM060+FcLXqLIw4LB3d3sz1YR1syQqF9Tv4dz
ZLFAdYRG/77dXhXTzp1t23SvPn48VgaqYiBaC85g59c8bF5qfE12k+huVxhyCval
0kVExZ4FzX9TfcFlZrKI9Aaz2r47rsFEHAM2W4xcbjO3W9vYz4ExdYgPR2SUaio6
bfOnyGaHGY3byPWPygYbOpnafJS3vSlxO9iU+lDYCMKYjDNYrBPCY6wUrnkMT2DZ
X8ROaeQmxCDHARuczmWR+LrpxYCSsEirr+qZ1InVI2zUaBTe22TqhHEvpbGPiINi
wr+U3WPAWBWw74f5hgWcIJeTcdZzkVbPRcUfrnm6uxMOPd2Khwz5axpYUN14UtC/
IjE/9KrAixm1966Xo63i5xT0SjJlpR8JPTpcVrcsOYW1KFyBAI7FQF3i1upUWOek
prtwGwrCh7mQEcceTR7OaGg6MAV/Joshd+/eUXRFUXl6FGfCD3qeCTE8hTQmb9XV
dv/+2R479c4cqtkH6GyqwxCFjUMAc6d0i0nstYr6p+5ovIxmg4NHFpaig9BwP4Sn
P6NVIkxwJFexzqfhdCfGlK6pCiYCmPp/VBxa/0D9OIgbmH/9H4pm5r7CqXq+6+A5
Aj1ttg2pxfrxdNhSQx1Emalhl28yiryWUulKqE6fhMDJVwj3u4wPbRxPBbY7/JPI
61JqQAkHvOdhya4poDocG/4ylCnVWr7su0Oj/69YaS2Vd7kK/k5qLeAq97V+SVEZ
hUUFrfZ2VNUx84oK9X+muB9FOSlhXbnmUpOycE3xzVcgppnpuQr2DYkR6oybrbJx
etc+oPu6ZII/gDrLVVicGMAAzvVfVNn4PRj1Kv/nct2/AbFvxAxaRa2nk5YEUS5C
ooYXXmlZBm+OF6WhggriE5AfBe+4MCuvlw03ognDXO8bYNJyt3AWTo+9ymcze6pa
N7nQq0k28w7PHLgx8KWLER0oJOhwYVL0l7T9Qrp9/JQlQ1FAkOEDvvWPexg0vINU
whyOoyY0NdXMYwBBtKW8krMvDAw1B0TMvkX+uHCuPjt8gHtkNHrytKVPn3aADlUe
Z4jOS8ozbHtQbRLMD4NFTazKmPFe7D+CCKvkKeBggyZaOs4eXT4u/uWw7CJ4rsYV
1kEAQsy46oeFnFWZ/tynSpwCXKZDOEndHm87K6LvTOrepjoLB8GdDcg+iIXxwHo7
f60nFVdJbN6IZiVAGNBFqno/t5cqKhGo1RWmjFSDt5km5Au1+A9bD3duCDyrdlR+
EVEhoSInr1nfxAL3h9zoOG4t7rMPdKRWkz3jv0CwSTHRNzU297xawr2OzlrO4RzC
LpjJpAAa3s3eRiTG7CuqzvaLFui8YkM9P7QZsOdWjU1GwUC9surcAQ2s4T5cZSYn
oLM5bI3j8+IXO696eaSUIOWDJ7+7tnSL7QqcPznfCReLFSTtsut+rK462wuWad12
agHAJylJK8yE2QYvEI4+qFb/1CscskXJa9VP+z6OirR/lQhcVQHR2iXrmpXTJhGr
OQJv++EuI40YQyu7dmDt6k5lmbvw/iFZAl2F+Moi2ypObmUvtsqwsGr9LM5/9MNV
BXDTOXtEAM2cuwIT3i68X9KaOxJKSwXUWcnWgFrQSEULZbDoNzjP/t9XTrg8qMTY
9HOJ0no4GsZ752QewNVZla2XsALGm3x8N5jVSRcvxM/EAeMez3Rz0uIaZ/b0oWrB
gVSt4hvoMxkEuXou+Rg9cvCIplCdX4uJP+OWEKxL/h3Web5pVyojwe21hu0Cowdp
C/OVkUR0atY9B+aA/8gDdAi0T0UlhsV/GE+CwTUaKT6TDU05bTZFyE7ARPd6fSZF
U0jLLu/e2OIuGm1dbUzSpQqGEig/jjAAzhmUXGUzk6q+2uCV5V4cObljkvvS1uH1
QHbGV567T1VZYlAUTxI22KLwwsdzhJuRhZYRZSiRcuybeuZAbt0RXOajJVfA2E+J
Se0InMgMm5VE/iXsHqnwP8JC9Ga0uLD6abBccdKyu4cSIokKW0N3DIQGhGMsxfFS
QtJudl7YrT3lVIb2UFkzeKjcuxE9eyi9lANG8q1xE88woJWhFPf1PMAjRWv4Y84u
Fgd35cH/zm1YHl8i9mTVFdFQnotVRlUktBWFvd2D52j7UmwO+ndfhHVNiKvXXUlH
Vlx841vFpxucDhmASWZ/xFlnrKa1PCI/APK2/H4mnaEbWPNnyuwNOxwbBEfe2eUp
crZ+4CH8NOZpTdpy/4+FMsqyctC2WMH8SLxH3e/IH9W446kSf6M8fAP1Xa99z6vc
Lc9dvqXO7BG25V1VM9quk78ktiWwbFfpInBzL80QEeRIBxvGc3XEtWliHDh1Fzkx
kxwCDaiESCLd2jY6L1o8QOHh+vj0hOB2l8rY5HNwgNRRC1XdJKuA6/HUGNGM5Sj4
BUYvJszESmhArAtw7lnwXv7ihggCURxAczy3PSydJ/nszGuPAVhnODfWt3kHH0Hk
UxG3rWAOKjaZTv3TiC83MgEW3liYsDkPP2VGzc3FTptlrTSYwdfYzVi0pK84idzh
bpSoyBiJpe5LTjGbtr2nsZKjQ1POonradpUt+VGx7S/vtKQVAPry/GSli8hCJmZF
wm1NAvlP0KaDJKIiFrXAH9fL3katAw+UC0ArF/tIdkPmCEDLli85Ic1Hrqlbr9BR
33DrTo4kvDoNgDCMu8lz+XTON+UQg+gfSU0/wAcskJ/ZoZhOIe4qjDIIkuek+3Ll
Kb+V8zCTRd80ZwLU5hCXwost+Rzrwvcl9lyq+3OswQBLH1jNSJjRT4bddT3FZj2h
qrw0qP3fi0CCJp7llxenevyB1A49SbxohWNLKDpFrKIQCCNVq/YjKHl04QiafxRi
AK/NWHtb5X9lIOB1c2+wosYuP2yDJgpm2Y/njwrFKMCJ8ZNTTMjOjpqoLS/oIkw6
8UNBy6ZGjb7XNjEEgurPAqh9e+CWgUX0nl4nvy/veJi47uS0kzOjW8gnDZG+Vppw
ijJtTDIc+yo8a4vEwGZY6Vl9zqDtwwMtiivCMnEpKYNkRN7XTmBKlYIwogANtZmv
4g3xeSMt8VXxXQbPtI7ZpyXrCp/Hxy+nEr9UzZvmeGL+djEZj1nW0bFUeZxw4e0g
nZq8lgEImsmPyGBK5U+qvw/kseAE0DWRFVXXUnZCJPz8C7VA+F54M1joSgIpCPjH
PLcvWmvJKuOEAdI2P8JHTowsjT/BlnB66zqmikHlqkKl4Bkq/CORU2sJcY5nOM9o
gFnp5sZSxlt8G4HFHbFio752XB/zzVcy3ytLTuwWi6wLNTLtd+B33TVHaJjl9EF/
z3cNyueIbRvgEaHY6RUv2QNjUUmQAta5BUdc0xQmB4xWy2FxOA9aH7Rjyrnbl2HW
VB+hByaRMAp8I1gv//yIRzzOLfdXISqvk9qGJq/RL2ygS+qDJLo6CkarBt5Rh659
6LuEhhMCJNgyhq+VC6aWeN2X0ge4Nzq/eaaA7XzLLUMY2YkS4CeM86G1tq7MGcEx
ABw2didyA4eFxkpeBT2QtjENMMA0ohcoS5Xfue6emjnKMU+gpatXH0/PemVE2fq3
RQK3HHJWXQ2yxNE9mVgulCWmrC9EExNIzH8rzlUYasxbiyVojrhhfRpvqjmcH24L
2D95Eg8nrADFlfAdUs0KS8aild7PnUglQBJCAhJZnjxUuEN1FzzpsZpM6ejh1DXs
TAbyWAFWltyIs7Hsn+jhd7leWt/Cy54BLtaLfCGkR0bnGigmT+ePv37DCSoxHqmm
Y1yGlKTwT3hl4X7W2jtcaecZ7g0BR1JWHdey01FapTdRazgDeT63NjHyYw/RmIsq
kcFqNiG2ATtoC/TatCPqOze9TpBHiBcuoGHKOZpdYdJQ/cKMdNHszQFawg6sXHeR
KTo1/4zxRfWb8uMtpImgjf+TfoTf+Q9XjigqMGB6jHSn4F1VOBDvcGW7KPNl/B+/
DyrJeKTcGR9iu+iPVmvLo8zZ15CrQMKRUCx/Tz32aPQEU7/QBhefnJg87I9SKxq/
gmufAuCdtg1L+FzXTEKJUWFXiQg3QJBx84HJi2ZEEulNJJYSkts1pmvfq7xQzwZR
AVMobrsDJ3MTRtTPf0guzWvObNJV3Myfq8Vkco8PMoeIy98jGOmVzOBQdKDTflD4
psm+6dU2SzZPcYw7lqExAc46uQvfjtnOG4uGzVomCJgioLM92wJGlglysObr1hSx
Pme+w8X++xqmrefdO6yePaMgU+ayi8YUgj8WqVb7Or0bc0lo0N4xzPJKYkE6k9oJ
Xf04iFqhWt/TAb90DHkSer3jvrkj6KIEfjXY11xSpP8Swlp7w7q5zQ6MhYYytdMb
Vh1LjWMSHKb3Qm5X3aunEhAaSSUWODnQlp1kNjL127HNNvBXfZYtjuEskMnUHME3
qfXwmnpLKs0uEU+Mutln41eH4ImxAdoYPT9Rx9rIfS0vtGuO154TLR3MXD0w+GL2
sdUx1FAYpsyB7K2Is576JKyrsk3430ADy/xgqJsfFDATcuu8pCI0exJqhFRjwzt3
AbmixuwBAoHaWiskvazQZIBf+TmDbK+4q0GTaMv3jfjQviMUw9Wa+n0PyElMm8Tp
2e4bAlwztABlnLZ1y3R4F0j62oeMit6aKAGcvpJft0EKlEfh/DlyXojwCWC5hP5T
Y0W791UmtOOvS9brJC9L3rQdBbDXoVskM0ALDT0l2EmOZTt3pGpVkoU2Rmp92CW1
iObOutVEvkDF48OzERlqkWWlACuuPNTByAUP97S8OXTIswaniNNE5uXke0dgU3ol
0W13a5HHJa4Cq7ScTEVs1Aimc1qaGk1vSzVV/lM7SgdML7CpZjRALSVRR2mXXbR/
tN6GQAHRi5ye+vPn0wzu4gh9/e76yDivsSTanMuXHv4Y9Klvs2HTpqbZnqJV3CgU
mV0Mt/2COcI0VWbbmmIZ7mKwWtHzKa1wsTynLuodcIJoqo4XkHfOm6nM3pUqWoIM
rlchjnKPuJYLt+9Y9M4fFt/5Chhj9pmMVUjKfq1QypE9TGLCzKUIJegQIDcaRgfR
PzBkjfKUEKwMRVG1++hMfCteiz17eH/qtP2rIg6t3bGU7i1i5JBV6gqX2QoMsRtj
NKgSfaXf1V4o7MLeL/Zt2G+h+7qBV7iSGzz1/ivXomnr5K2rReAXRzBeKMEYBYqp
ts51aLvddPpX+BL0x9ehZIhNCkTqAeQgOvs8GCdUXoi6HYtaXntUDGYTLbp/Dn8m
Rg7+8OXaFOk8vuepcv60IbN5gpstBwJip4yDFeIZCM55GlnwRQ3frlYqxcKvS3B0
6WbuSwfnW8h6i/PxzBgg5tz1k//XHFfjbE/3S59iiGm6LTpQ2knXesTcMY3lFkPp
hIcw//w2MYky6MbRID1AJnF+bJhTj4DcuKEFKYAOCJMjrBJ66dDM6mDHgY6BdSC9
9p7/FvSJXAa7566g37H/SDp2yM+8aKVg0L5O/ChYK5jZhL41qNkAEsDLjiQCqJNa
gI5p8zarVSw3q34waqqjeQBrkRpDLL4QygWJ32fKPkU+OZ5tVcjNNkp9N71AAq49
awc5+roszvTTr5fUnYEgX28TYzjTvcpX1fDtq8+I8E6hFzGVe56MNPYMucuX7+o7
iGOKWeZCfW1rgCV3ykQli/cUA3Hr0OUFg0YwULwqRwe5MlSVAbEtbF+Wepl83J+4
tz2a5YLdof7LAvRQXCUfRmbo/usFhOLtBB6sZyk1fIYxMx+NmJ8lVDFDpZnoMlND
W7R65bDU/o1fITow32lPlG8fNyPgw/vsATQDoFYfHzAkhu+8AcX9mSQciY0w9ciU
GFshYCfYvcqJO6CjamuJV+DWxfw5y1keZB1fGzQF9uaBPc/BcXV8G+p+62KWCQjk
NaVtjsWhkfI1K1LCdlDdQzY4EF3qVpQkomhtzi8nHgMNPGAC0WcltFxGf/xrMV2Y
NR7Uy7ghowLnX9SndWrcEgfRJfPC5lwNQgAidYU9zH98kur5k7fO+xYJL4WU5wF8
AJubCI2uQwcATYzxzXC7baV6FpCc0rAAbUR2uRIKPSbl9dCY2Hwj/C2LaaLASPmP
AUwDKvr+GUbSbKusci2/6jBTDhg0fZ5zcqBwyMrlYeapo3Q3kWpuQQd3NW7UXEiN
pXy0JHldRTcyd5LX2pjL6+52DDKe+wwt1yUxImmZsENy9Ce2NMjKVUV+ewNGBDOi
ZhYRqYqaRa1AmoovKptvQ37BjgQ0zROjVtlH0Y4cMZh3bEabdV6Em1/2YgJ6ggy8
pFWwsObX1IE/3NXTinAG1yjZ9laEqwrOva34lgRQEVViYN8hDRkYaPusx0Xhpy8r
Wp162eWA7oFq5U5KsFKC8+/G6G+7KrRqwShgndKYyZnzl0oGztV88bnk8ViI8W4r
NBfJ/6fz70T91s3vYUIqFahLsMV94KNN65TTY6k5cUqV2ILZBTDzqg67M50LozQT
IS5igpbwbK+9yy6ofTJM98Yek5D4JWN+buCxKW17e4gDgUdrJyRjD/miXEI5eFIf
EXDN5W9vEFyagikSnI15LhLhyLoF8iDg0GudWuyDj3AIqEdXY3K+iWbqFQlEyPnK
V/mkVMaZ30o2zLRB/h481D87/kQVIQauJAFr6KkkzslyLx1FtNMI1bZJELM8AUch
HoYGuTsr2ByHanM9Fo4oroIY6XafbSmXtwUu5La3O9TRTbjOSOiKtP6DTDS6SYdp
aJRPMQRuJThjPWk348ZV+HFllL1opiE1QhCe1aqinimXRCsPXyMWi4DIeWK6mVGm
J1qJ76tT5RdOlMQp2+IxIIjPXzzu5toJZpe22W+4UEEFjTEj0/52BzMMgbO4Bf6p
8eydpg/qAcQOz+TFlTzuCYeEy2hH+zrgdd5U/l66SDmGyYZgZ4XfmnKDV6R5UGdZ
EUOmKKIQl7mb0W0XIeH7/OGPUY/42WuK83N8JrcDADQq+y4tu/wyO21hmQ07HLwf
PfcK5cZ/pjAJBid5+LBgCTNHU1TniBBAE8IBEFYPNFRe6v+wNExCbmth0NPTXC3I
mpHLHU0w4YmG1omav4pnsa8MR/bGW2rY7j18ia63p0IZU/suUm85WRubI44srxTx
bauH+vjbgLA4ALrvOW54j7nQNUrsZYG4cUCqJfUUdpS46SEceFDYY4vx0skiYcMv
ipz503CikwBIIveyyw8OkGpX5ML44u4jiMiYXjbIr8sSDk/IZlKTqTCqCG950d+Z
ihQOwlIsogtLrvg+Ls+xHGBmx+WAGtrDi3oRYdtjrmI8KEZRPOPCIRkiBBXpNEof
td4Wl54fh7+lx+iEQB161i7646lNzPEQ64MrX/tmMTn0CMsrurot36oMjQQmvn2F
KyiL8G0iPgQgg95aEO/BQxmPNxwmaMbo6z7iPkS4OQCYbwWk+VTUUi4q+/JY0glg
ug/SzETwzAfWttnVfLx0FAiFrDlpRYKkZkt9NzCkfIFMXNtEFjWlvKbIWWSMXtv3
oCrSP64C0WwUeHEAQ7DjBSY5kw2xU/KzEqp4M2f5QwKUX01KTm1w74LXU7inbEeF
qGw3ssWCNPaHhTSNRdZuU2AuQAwF0hvYIcM4GiLzFVA2UkQoWrJnn3QlDAAloxhR
E93Rd0FK0l+LocbBD+BlnJBU/bExnfYHPmS/Vuu3gQpQpX+byN+F3mXGrEklkVbV
lekoUmCqbSIKC3OhqbEnedmDesxlyTddF6wOlS+DhOoWegF10eThR4IhkM74SKWm
DpzWBi+iSjg3yI8rBFXwzI5H2PWTJ+kmyTuPvExpVoeOCjMrMLTwt7F4ajHaDAOz
cQ/qP4zIKy/cs2HRav68o66UqTH7+GN0z8238QHUqAVWupSnt5FMNUypOkDst1yK
cOKXiEe6SscxaBlLErPzJmaJElozESDmXh5YpAJyd7Gjy/mARxi/aPVRhBQC0lo4
qZ1MZbegFw21av/deHORz0VG6Di0WBLD962nu7Cvxooyd2JY6XIAxNYEHj3K4K3/
4YOIzHwKgu81f5HsPD3+uVWflTOvEStVW/3qmxzN2Nn2zscH1qXWA+/UFBbb2IgH
NlEY88THL7vR32Ga0vtIXmmXIbcazuIFTnN9qo8M44DksNUUai0wtkLj6Q468TRV
gwpF2RX3tT3EY2Lv9EyGXNaDtidxuNzEVFaWFeV4Ifwp6OKJkryXlHM9DAc8HZaU
2SiqKIy7BK4/hJeXKrTvXjPruCXx1boyiLiDEnemPrcG7T0thzbWNoN4N6rc+FYR
oZAYqPM/FgBGO1TGiFTaq85lYPRfVWMeziysnXdX5onIq9IVoJuk3NrFytTxXTMo
NONxii4wjJtSBVcJcMCWoKs7N3rFsvH7RgrbRMTQlfnbEhMdsseUb3yJClVW81Eb
RXo4bVplUU7+jQ8VITD9NaKSYQFRZANl1flXXOyGZziIREvdkHUX2xZa4odZecGE
A0H+mJyFdZC9+k3N2iJmVQX+YKDBXuSqXGXQCpV5qerS4krfuuTd4gYfvY+9XsQz
sN/VbKDWmgf86PMYgQ1ww0x7S5bGsKM1uoN6DYELMtlsohxklxgeO0eDnyQXSmyP
g/HtC6dDVBaSKHx1UPuXkP9/mMPguDTN18RaMAd5Yqwrxp8BW47YTduhxIy6lkZ+
CaU4mrPu+w1pjaGy9CyySgGMX/qzxXjO3X1PEaNP7xKwEuXKlFbya7NKBtlMPkJw
ZQ/WqaCQIRboONRlzYKnFhcod9w/1qfZpjoP4ZDias2q1js7R0eR0geSz8WU5nRX
csYVz1ARdo3VEM8+TGsw5WTDx8rzb3mghAxYSyVaqBc1lI5I04kLSoRBZnZ9rOK4
bJvLVOcOqWtIp9O3KRwxjvCe7O68tG30pLJnkd+Aw0xqIyIBGt6KnRSEL4tuCAqR
zG0CvKW+c5MRE1AZ8N9+WrV8S57kigakmHHIqcEcdpaEYJnYdu06P7/JGUnVYN6o
gGx/rmtKoHW4Nn7rd9Pn6iHaR70hdu91i6kqNqYCcEwlnkzVrUes4LDYYL4COhH4
pCny4gfvpbKbW652D/WpR1xwxtUnWQES5uXpamfab/uOrMV53i+kD/cLn3adQ/O+
HxZw097/qhYe0cCBcxtu4i/gx3Lw2V3xfGgeWXvgJMdAcgh1ZBBlmxGR9l6lQX2Z
kuRNAJG+2SUDYzBhSBMxGbKFjlxLY2X+azuQa/kDOtXL2eHK9pvTMm7yehk1uD96
RFLGRwct0wu1ryvnGkOVU0n8Vewx3LabihBbErXV4yFrpL3YA59LJTO8lRe5zOj+
4PUCwgIpRBKffb5uO6E/jQPPKyF9o/JFtc/PjnvV/zRC6Byt32pUSCMjMcXe7WYs
f7spzCt6+LOXoxa+m90AoINUe/x8mC+itQC13rhD5L1RYp9TQqgyX8lzFimZRDM+
Q+SYm8XvKBaehNU5x0fkFQz38xQRwsEXRIr5cDk5pXxlhIohU9G1pfwJTO5iA26T
U0ZNsTyj1wAgo7yQMecQQtJp/ClYnm//oznIbILM6r9OJvwwimX1hIsOTDiuMBjq
b/Da5/KJoKUgBOLdLOo7nVJ5vsXCz8JVycMfA+U1x+lO04AS3ELStXpX2otrB5a1
cqX91WQvyhEp0K9pl0MIQDnLOeTj23JCt9oNHnD8vU+fLYSMc4kmXfwWhcCxuKb0
2q9gPvAUr1Y40tAlYD7cKeqeR4L/jbkuddm5+vx8unX0yKa/0OiRYmJr+zeTRkjp
RTWFNbgE71Yfluwi7Aj8nlua8XP4q6NsEBiFtPRSU/dTakVSThNoEpGkp51xtRX0
iTFfT4vmzQDh6Rf7dLeuiOsIG5MezqcOfN6z2KkFvUCUTD1UrOq0wPKELEmxKNDk
VAAyRdcTGvD5GkwTefVp43+2TDkB4VoPf8Fx/3RxT1DAnbDOSwVfS/VuhqZMIPU7
4c9YRlP4NpGPpWn6S1tTLZSc508QEPYcvDBC8+oqcBa7lwYm75WP0hNpYtdQEbfQ
urwv9NYCCDI7GPFfqMdTeHNymcb9MaMf8JTfX4wEajSVdTj3p0y/Q7mCRzEJRkYr
QZSZIoKCi2fxH2WoOteJwUtl4NErw306I3iHTo1ho7nuKEYdaEUMI87/bSFJHrWf
0pl8uqj95e/gbOerB6OUCmQEuouvTEaXguN/mFfwyAySAO0bY7X2EwMoRO82GOd4
zG5KNCKr4EnB4T3P7Q2lKY02gxZ7jaGsn/h8dANySmBtazmRS8OuvhkaqpHC6nbH
OiQaXOSg3SY8PcVDXY5jjsh8EbV7YT3y2hGVZCk6BC/r+bd1EHzvAf2INkpuSqFl
csRcj5VOsBlg8UFmXifB7Z/XM8PLa4NUYM/BlVaZdtBLNC+94vls6m2876EdHMR0
lTK0K/IfVH6eID11B4+wpmUuwzC2EYTADKV2tCgUwwqRD00bfHPWT4NvvMrBy96Q
FR3pF1PeQkJ1fzm+mG0u6f0UwjM1yCa6W2EMiDtF8ePd9MwpnWBvyAavNCjUuLGm
O4M9vdWVyG7eo20d5xs2FI6z5rWrn305rxQOO9XkTbyYBnnFVCCSP4jB9as7Ph7l
aL6UPu1Jf1alZxuOeeQ+XTcJRbliSZh3zVaL1jN8a5cz4fNH57IL6IgxJk68yoey
nLkjPfi6t3FT0DoCYwuPMNpTWScS8VxhYETEAMT8MO2YMTUpbq51UieuKTGea7ha
BJWRCGEerobDxq/JU0ib4xJ3v39LSPnPhLBT1mOiv2lMFgXAKrybyrcoEmeZiNOY
+lhF8yX6AWP69zntNsoWJ6vC72nV4kaMy0RswReFAwco14qz/Mu7BpoNBOw+5dzd
lx+rfJ6cO5QSQqQJmYRF8uCHTe5dRWFgBZ2rBoXdRWRdz7cwAF5JiaxuwCvqoNWi
fRyMT/b3W9AYAPHCY5BGkWoPnEQW68tBW5RszrD+JIbYl/3XqFKvunnGFs661vK3
m9B56ywxlWwW3pWZuBfH8KVBplX6fn4yleRBcYzg+myMKC35SFdbEmJVns0a/oIY
Ul0ouaDWdYGutNbgGfQJ9jE9aRo1Ss2Uyoqa7kgPVzbtBhN5HFIpp6hMdInmfpCG
iLDsBC4CYqCN7oVnesogrpKR6cg3+l6rZdixgFNA1Cn7pwurVjW5rw5t9sv3HaCd
wwaUwbNwVnxJbVZclofoALK31sX4+lv9KGLDVsGW68QrY39ItEIZTsrCCoW3+fJI
DchEL4s+xP+ZVLqjf+bdM6deWvaD6eS8nBxIyaHgFvEnmU9ChZtq5UQWvIUbnLcW
cPtH99QSYucNqsv7DfD2HQzZnWa3Pix7huMGCoLY6fXJLnXaBqAEnCIcvhG2mkeW
mtNdtoyreHIiq4mWnxJXvZclQDFmsf02M/iH2eRuSSuwQkh08Bv9xXy0xqhVf9Yl
IYz0Y0UrYa7QUxcYoiYPINJ7Jd/0Nb5fA242EEYmlfSSaAuaHaVtgcVRw7fBvvqc
krztZbMhQecm4sQiAMB2zHtvqxrUuh2L9oGAZx2woVF5ZfeFhEPpMzhHFYwE82kX
jXFCigAsI8uNvBdra11iCxi4qBaOfhwd4KNgbKPDNDxoo1xGVoZYGvcnYd29x4CX
LlYjvOnXjrigkBPg7G/WAafLikm9AvYjstPNYF1+nXg1PrU2Fc2efi8P2+8GR8kp
JPcTNQKdyIB5sBE5KSXa4WtutyVhim4Cyt4Yle04LrNHnOL+FjZm1otKvduQbY1J
kn/G24k/qEbK7p7slAIXGz1hZ+aW4PIlQnKxPq71MyJZ583QyYBw9xlAOfcimmmk
f294855T97b9k2+cRH0q3AL2Z7irrHwjdFddvuoqBF7/K/zg39gmO8n+5JPg/2eQ
ZIwfQwMSLptOzScPFruoWAsfile83WZmZCMrKEw5HU5jVO0NR+Qbt7z37pTwupHl
alLSrk0byxqVrcjZvxGvOWUOdGHdEOMI8jf/clk1rbtmaKNNbBoDH3sMr8pk/98h
wtpTxSKBH38hLSj8FIr+e87G8Z5iXxYC0AaeYjpgTokgrz8zCiqoP0OKTjfvRHIG
cV7jSRU5EX9qXdr4AqAZ6xdMY3Pu13RAFTIVjtD/ZbVbQwA7udGbcgObPLL8C5y9
0qBq20RnosamYBSDVNvLD4XKhNsx3WHWrEXOpMSumIe2h3L/KdG51ZCV4ejMnwvH
k7NttdDioUuhDLDRLWWaYAg+xbjjiJXpwaYPPkjXcvulT/Bf2moew/AxtaoHnsaR
mb4K1ZFXhOe7OvJIexK7oXOxIWP9yvaXfrxZVoQUQAnqW/PTdZpuWnEPIitLAPQZ
LPhWPnHQXfr5EJDCuB/X9ftNTct+rsN9neRTUy+VjR6vlbwLO3na1C00PqykLawe
NjWFQ6aEbGe7IJi8ZJ9RLD/D5M4Ql5LK+Qp8VQ3e94qKzbQhrhWcGK7gS3Gch5YB
EjBz8jitoOEE9gQC0udTSDbOrGikFYMg0+McKpEZrJ+m3sGrpDTZW7nRzpHwMsPX
nsyzgniNeLUQhg+8XoFW58DNMaYJHLFX7zTw/YfaPqO738WWJ0otjNjIlNwTWzaW
JChUFc7IaehWTxOgxFQHcl98QTqO73TWD7ctooOaZgS53zd4dT72YCvy8wzZggP+
htPgVyxBNZKv+jDb6uM+fKNTpMH2lHjsrZqr2nnMLxxROTJCHT15iPhnAGkxd5NN
QXHm4szT9ZwWvLP7KjD8A+b52W2ivG3Z308TaK2gsWTzQv5S8c2fULmCfmyDvG+h
V3sKtxb0SKuYK7+rRKm2Rl1PLTJhElbbZXoSIrj6mMU4Dd6wCCXQwF74mFIgBA/I
Bx2gJmkuBk13NzzWR+JGGSjVzR8u0XvCA93SYR0u4XXpZseR/crVjOR41aAuejjz
dSKgNsprtB++nH3bqanBNDkXyyauQx7sQTigtQqGwbXAdfadUtvHzyDUUHMUFZou
kN5mEVVxX6BNtGCPyJihxnBmjAUtbyyZ0qINJk1r3JxfcTHoPd/PvnrmzjVrUpTQ
lf8YIVwXdQ17bmFb8oLwaOqHx7W5WIRaOzBjkxgQFfXUW3IBI4d9ds96i42Cx/ZY
nJjPA0Edoen7jXqK2MAwvLrZZr703M4ZchDeeKV3ZCXDP7gjp4z9veeB2pTW5CDN
UaaS7rpLvkQ4Zywp48Z1PJk+Hd5naGPWvPLnStND0ZUuoQhdBAbEllF8Rg8bwY0N
n4TOgpuoEuf/1cyvnwE/UMAbVG8lN+d/1Xmm2sRF9z2it3z2dlL5L3QNMR5YtgXS
V3998HnYoI5QfS1BGxaochhFcmDUQ2uHqthcKL6dWeWGVZU1C9eQ3vBFe7MzG8te
1kdjo6CyVFcXePqaIKCW13CF9xy4FZ1OOTluSWarncQjLO3/vnfbp4TSFqzuSy/5
/wMJfRFXK4cJBRX60BMgZqCDoJggZKw13MbtyAD+DUQ1pJiYiiFzSfc/JaERdT0o
ZoVvTDQ7whrTQ6/KtrGdXSqw8eU0eqgxWF7up6N9yvCUAQLaqLrVk+Te9K4azlDx
GWcc8+HELK/ZL9aU4qjnMbDa0kTaV1enRCpE0VQ6dZQtXG7ZukLzmVQWyWH/CKz3
y66q8+eVwD7h5s7SO5xB+WhJtzkLTFRUiy/OX82O6AqX9hl5GZZ2oFmCPDgM4EMG
29BsCjl9+AZ2coCH+pBGsXuuFW4bD+HzjC4CxWGE06UkY7lESByJT9sefX7OxdSm
j1WB6Es1SlSFKeK9rzbxI0y0Foh+UxXJ6kQcVTf7FbRN27Xa0umnsyDCrCWGL6QP
NWqery8cRmN0SWI6AJoWwIbucIt9/E2p7ScAA7Vupi4HSLDUoRDWob2//s6H8+Yq
c7eGYo9trXzL62K12CziLRT4m4yeavM8oymLt8pxIqhgzsUaSXnF0yT78GJxxVK+
ueZHGSLL5BQvpazt1uNdw2SAI+YRSYjnWH9H5CCcy7Q7sc/FJL8HqQnJ5CCDC2BL
4VG4XicV4bFgiZZXSHgKi7tKliD/5efas/jaMs+5YHZHwvAfZ5ogrfFtZsA7w3tk
ybbTiZKOryc01smofjeQmSYsNlbCsKydyGx+728ZVE8S6uGlrK2oGHusQhUmTCkn
KMuSWt3xapWye4sDIeMxlwEMI9AKpiaH1uNcbxEv4zFsIq07nye7Qz4KycP+z6JX
M8/NGmynYnbPrC1JnOQFcZRAnIB/SsBjl8bg4nhganTjN4y9tr4gzJl3vnfsfg1H
0IxgB8VRgk3yIZdoE5jLcPz457qyPWyZEqtjyfKLKKajEQXAcv/4ayiX+C2j5SwW
54iZ6Um45lLPVIZZtNeEkXR7UNEwRa6ceWf7GgCL1LX+3KRo+eKQ3reophD34KsG
n9uaFU042gGcGT2e3MrG8TAt2Jbr5FBCddwTA8LjW9hDqDrjNL5I2H8L9BfD7Hei
wxSZaVNibziIQvJ2toBD1Kj9+Zw7RX7BgCEqkjYNo3aUWl7Cbw74w6Bn31CY7NR4
L+sPhXKHK3ek/Hz34BKS+BhuLrbo94JXn2FInjXBNYychDcKewagfxiZICNCvIaP
odSrhQu8lWH2qe+kohxuLPlNG24lujaWb72W+C5ofIex8Aekw/8diJ+ENccl2aF4
VMefSYUqBhbhQ1qu89TqdH0bELefJtgq5eCZTSHZWc7MZzbyUePptcbBWycrOzAE
encR32EB5IGiiyXxOzraG1aLg3Rydydr82iKdKZFIakdFhCeeHEyYkD0Yrzt49VV
oLjc235rSkm2xyb41PjNjbkj2x7d8Stvg1kZgM9AVDUbUjIJEN4eAAyhy5plO8u4
ZY18Lxx6IXDAdZE/tQEi4Rs6tTj5HwsZ9tLkH1316977zriPke8vvj/RX2EK0M/W
SbZZjwl1OiRzMBKNMLcxJxwFgDRoxtYoZe2KxIQmWvhL+RoKuQQw79aQy7lufN5D
NpDuNor0TdRahpyHEyND+3okut+hTNj9Ct+npUfGk7u1JOuNQkousgA8VXuWnpzo
Z3JJC9TkSuVXT6i3y9hrzTyogzMsd5kcF737nTUhBmoI5opRcJN5wh4B8gT5oJRg
1jFIvCT458clXqgYjue0gBOzY0PPW9ITQAk+Ps2c52SEbf+vN8xBOlJr0RBMrjwe
DQrQwdVORdJh73kkSzpAywyyVNzS56/qP11ay10GDTI3X040msA+GefA0p0WO9CE
n26imi2IYT+otpXCY/2dV0XPftXzhnpQQz/kC5qPuEpWTb50hKiALr1hoFWUTTIf
Tv70PvODKx7vTI0VoJhuBcEsF5YWGTU36htvpovblkyCrNk9eEinsYumpWEgArQh
18sDMlzMQwiyTeh93HqCXjGjrVOOcJT9wr88FSzbO8q5TPE5+pa9laYgTMxF9MMP
52/YXepgRLsl0dtsu02bp2N3W1aJ6CqJ9sXWNlgvnX4wNxzgVencV6exf2xQuE6+
fSVUG8WQscJuQkqaJnKHsddDW+WFcTqSAW+qMl/+6+iTmEkegsFhEDM+lGzrDWGI
hfm4Hj73qYfcXzJAys/7mqXu+wnFc9qOOFXNGNCuX6d+tlUYZTovl28lEabwol0g
oRGI3yQ++LExo5j+qylzWvAjYoNGhuG+xKOrkmcSGhnVjAYXAy+FuyERHw+ip3B4
l82pQ20Dx+K1pUXOJKX38fa2lAtOb6Otr+/sHi511EE0Nub2sUkieYssYX/qR5id
7Tx8L4z3q932/1YL6TeTlcZidZSlTM2O0dvhmQIZhg4ugu+49pCu4m+w3BHlYodR
qSz6MVVTPE6BmZAtLVgUUD34MQ/Ohx/gWq58D/QI0utqNilRgrUThls/qdO03rr1
OPtG9CHbn7EMcHaaUTkH2NUPGmgzcRXcXH+0HQil4d1oP2YOLAzJV+OqrsIB226C
OuzxRrjnaV4QQNoFrzxzoqT52N8MX0jFSW+BLkkHMwYOsewcnN1MeT7OcfoBEAuW
hc0MqNc0dZwvxk2Py/Z0scZb+VaaGOj606yDdGPQoF6xR6YOCzgdyCtGin6WMxEd
laO/6F2erIYMFc75Vy6q+olhuAMtQQo20/Y9vhbJ7hiS5qFntkDpVcSmyc7YelcD
+RL5eWfRLzYPNuOFh0ITgu7LoWy4L4WGA0EozUGEawwu7R6KWH7gV/kctBZkLThg
ERz3LcUYWjKjdA86X/Tr05wtB3J/MEu8Xl/bKEPAJC41AEpCZbXIywD2kl3H9umz
Rz3xR/fsO9C3FSsSm5dDFweeiVjvarIJcmRFJJivCD78S7XyeXltVFqF1r0XNCgm
xdlJjYwDwkv4Lvqry4x47qh/ZsU1QwDouye6o07qd3tTZt3yOxK9wF2LkcJzb9BP
16QWqwa9+E5RfsrsTZcqBGZmC0XHulyCkCFE+8f3hyWs0WHNgcZlHuo4hqtiR55P
B/By4gEysoduP8lbT9+JmGiNEEailWX1nLwWtmQTaF2B4KDUdau++qtMRZEAelT/
ojZRCrZQdKwNXHrmqamDi5qPcWraXqBQg1XPJN/Iky4JCSPCe6daF1kI0Xl99vYv
+vRg8KiuNg2heIBD0sXAsmW/pBPoPCMVNjL5O0Itk079o7rQmG1pcjbOYKPjnj2Y
A6nWXxVgQGNo4RvEToULZEGzjLxFXJjSiK1xj0flWa2nM6ybJr4Pizk7/ir9qgLe
h+p0s9WKMpWq3VlnwxB6cBbh0LJHR2iHSxEwPf7/lu693j26UgvBQasQjPdUJnow
Fd1oNTJagU8jYMv+IHxhl5AXTR3sNglh7cQj4hRB9dknKONW+KUXQTDETVUA3fAS
nRulLuw6YWNK5iMpN0xicqtjG92qi6hyUDcOwI2S0aUJaKpJPhSRGMYC8WIR+dgl
b3oF6vWk9F/h0UBZhC1LyxivGWvL+Xlu9Suvg4T/MISmzAJyAwwUaGgohJOKkr3P
tf6Hd+lXKlfbwkwuaGy2rUlOlML3/j89MCWJ0Ec6Yrb0b1n8U9ck1DhxvgIvGJdf
jtvCDIbJstPBnapQBAe2YJQA4dohOt1qq8AoySZ6x6y1w6fYSGtalyx4QRCdJu8O
a+3XxMM3WBOB9L4JkfSZ+hUTT96MtBIOKYMKlteLsZhMZopbSUO/RFrGpwh3/rNN
Wgtinnini5ByBWmPE8//31EHXQeR288iAdWw1OOzwHRnRzj8a87FAsVq0UG2GGSU
SDEsnuxs0jFknh/WRcax4b3d/5jsBgQdWMLdOW5diUaqw/nPnupvq5O/z4e9sYeB
PI3nQZIynYbdGehtStf8V2jCtGyuT1WBBJRpOMJk8vm7GMV5ARLOmmTVk19aw+Ni
kOM/Iai2v29WIpEmGYCmKBEIcV2309XVvGpchMe74WympzlD8LNh2XM5E8p2yunt
mHKKEsgIQOoMk1F/NCQrIYo+xgbIAE+v8OGEGWlMOJgyfyj+pAoOrX9Y1WeStN2e
PSu1k5vudVk6jZbXnLpdbp2cxhcTjh83nRrwm6jxRk1L49zQsIaOJ32Ei+84z4co
Au1abGiWU2LwLFTlI/A8A3jBNrvIZcCdF5xol527eoPQamIvCYy3rb/5jzslu6HE
H4p6FkZUUOlhCnPzhhh5lkWuCUMx0Aux2qSKHpQg9LFcKNHrgHXhhymVjnlXBmhC
ZEh3dQLO/9pH5n++R/0eTBU0Vb44Y3a0Y4Vm6wlEN5gkuRE5pXyYH5SFQ1tKQ5eJ
tPGEDA23M6iaoiRjyiIpJMWYZ2saeprqxUPD0easlVL1hghtpT1LkEgQAATLiRDq
qhX5NN7vtCvXGTdeLX7PYIdFGtRr9HFx4NeKtzIdN29lgNRWus8nkESfuRXSC74b
A686VVi0fFGfPP8sfHhOFvrEGH+yLGltS0lguJKwroGN9vHrdm9L/qzwKtoxkqkN
4YsMtp5fzu+u9w9cgK0MkVR0c49WadPjyf7I/miwGbTdMiACuvLkOXhldA4YWv5R
DJubLFROA7fdgCEehpz9MC1RkQNh9yhucV3bOueul04ZLgfGiaQSi1d9zZNZhQTr
0NqQ8Zk37z6bVUeo47BlskVpSJT5tjQJ2En/PZFLzWlBlwvB0hpWQpT3GxjDWk9A
3keAaSU1+8QnwCj+cWWWlbzJg2aGmJ/HecvU3lS0jBRnTwNuqoCMnnZLtw87WPU/
ikyAJyfCIMxxx2OUvx3TI3piug9OXh7AMmRyHMOtiJunA6sIxvXWAf+Oy6rq+5ir
+ZFPm+tiRiTLRSNB7KUmfsXBQoTnGgvrQM2VY+sPZW4EE9smnxHURd++RF4CmcfH
qMV9K8CyPfB6eqqj5g3feVWrMQC2Sr/T5PhXBmjKdeKyYHykTWp0D7CKlvrSaqVt
JhrmTBnkkOYtsid17a9fLrU6P01dzwtpMeMHfUFju2C8c55/4FQy51KyD+1+GA7v
j1Bk/MTIwCcD1IPCIzwpsCAnAruQZWUZPaT3iEYd6SIexu94bUebQ0f+nnRlTA4d
jnUsJ+WU0HQAsOAUHLjq19EcnSo1BDCj4psQAKaT8wQjgbiif+34iaKfcpeGGR2B
+pCXXmMvJUt8Qg0kT5uiVic6C1kk578DMN0J/MKJRIstqExAjCk2EQMNpGRHyyn1
iqm9pNofS0uNCHNQA1YuFLzpxMYSJGV8z8CXwGajmr1h9JFWm8VzVCQlZoeYNqf8
whyb6Lxa77sy468Qn77MAORR9tYCns2PQZI7iqWMJ0Nm57cRZRxmMIAX8bwyPKnj
KO3lCPiiBupIMcolgzm0AxZmjZ28tEKKmp6CMBAZccuevumKUakycArWIO7VlFN0
p8Y/v/iMfvBxBuWwSIeE/B2WJsw/5iXBqEsdmz0XzXFTAVuZbDxcsZ162U8Eyvne
pTcDxCov1WP7eG4e9R4N5v0cWhocZrockDTpleMAwPgap1Z23Hg4w30lcYql0Xyf
1rNdYHBcu8a/n5P4LvAaR4bxClM8mjEXFo5+mIscJsmEkHycw0Ds9R1dQKHgRoDi
Jh1hWEjkdiUAOk1b99JSr0QfauNsIXrgoPFg1MrPvwKZKO3t14v/caP3OWHfgtew
9iLlJEykRyizzPSKlE3vCMpYeQ4f+GWhiY2uMxDKte6v3tz3lkSx+6yac8qpBqBL
2d7SpKVjz2mzwXK+f0HfWFhVGIHHcWHjj67gKc6PpeZulXAoFmsZWSudKZSVMDX2
GgolECARyB+uBAphau7p4UBPcpo7TGDzv+b+M4kJbrxtRu5oo5NU98p7ugJCpXjt
DI6aA5p9UksG1kzUehGAWW7vkftE3cDMsKlSGT2CQ84ENV3HqSbcvL7HQTon/LXS
ZCp/mWTKSOrmSAuVBwmJqryHtrx769KcOFg6i+ll0oFVHYPiU+35yRQaSHGs+5VJ
8JREe16qeXuhwz3GN0EPiVMs1LD2KaC/uN9PurGtx5Pl/zlq11Ov3uIN9yqtPgK0
ApSgSEW7GuKKq9BFp3tqpBvpN3rnmn84faYOlszrkVaqgo8UabajCJhr3XR0CdyV
I9+90ousA0Y9YZUwIuSpL2fNIe/bTlp6XPmfYqZRCYcM0RWAzwaaUEVf9kLmYt8M
Rd3rLnVNE6Z6TOp6B0zSO47GhnxVOGKanlU7u0/i0OWYpN+iSOBt8n9zMZIs8EP+
PRy/I6XO/KXkCp4NBih2Q8SE5CZ82k+PHoV81FwX2lixoyjtl0VUenNWBTZLFOTa
0F+yg9eDqqY2VpFgEXshZTlyvpLCM50fb5ihRUjncG/vs608JS54Z1Xkz+SxG3QN
QRvkq84888fYaGpIeuW2P6ZCMFo5LlgNve3v0lKpa5h9ikQHTxIT8Zvi0AyZHBY4
Z8vFE1TdNlsc0HSxe7/AQz8BavqVVdEQW0YXc9ViSJ9jfVgkrW5SjsB2g0+aImK3
mZMog+r+pRCgWeoI/3LOOHa2mjKtjLZxQHfcm89nFqLOBdTUqxdqGajqXtFuyS0+
tzFJs4ZSTNW5shdrtUE+eRFEknBt4YdmMLvTgT/H1hn/0B/W1nyUizjdZgdm2C2I
DE9TGx92NJTUV6JiInJBo/PmkdfzillPBOk7Lglaz0tf8SWyyPY3NdbfO+/k6rIt
wMuLoMB2yGOr0EEKO6BYnhoTwb6WuSw6INRMew5WgG+ptu4L4laiYkT2r9CiBwKI
nUjVYRoeOyhNhVYvx0C8dRMKBqrqocLUghB/l1O8qzbGTBpTxh6qyJiWOzNAIsT+
48OMeVDp28hOnTwaZyy8WuLR/knl6H42wl7BIkbSp8wwLseUwl0H933ajj50F/8P
cSc2NMV/qNB4CcaB9NJlfNX1zDfpUnyLynQFcXMmboScG5N45Oq1ZCKXbcAh1Wgy
gZePW3gSGDvKr/1glQxQo/GoURo0gAgmxRPbBM98akBU9qGLsu8CBWbMq2NFK5uk
a179qu7s9YlXYL5ep4aMyDcjk5Yl+9JMr6BcvTNWrpu4Af4AiTAgtFuqTd1lZp8j
jAI60Wu2z1n1ufq4o7LoAzcwrPg9bDfLoyMJ/8IU1w59Bhr0jNbBM35EfUcu+Qbq
SiGqwbrl8g5wodyR3bjkMP4h1pr62IsSufYrAyJVo1lJZrGSfh/bMqVUGNsKcDhr
RTZ7GLuc5xWpxBpVkRrZFyrI5Pb6Vbk/ckD5g1KmzdXpUlm3GacYGVC8EfTTphXl
uesglPEAimjq1awB0+C42cea1gHS+1J9hK080xoUEIAe2A7DHDH02eNuJmBDzE43
OROnHS/uleq+jQgTtGQ7CyTO2jjoYYCC9QgLHvesPawJ9BrOfyDJl1j6wjFpLZCS
pwY5Y5eS9U9Htpall0k9tPz3vnOCf393XneGhe0ZJZeGYz3uCn06rPgAkGeozAZA
gV3+egv9fRmrIJWJEpEfYQ1BiS8w2/T8czAQAc2uSxvxpKPeYMMPtDKZ6Uj/uKwE
NbjTxFmSKiynwZZ/XcDLysi7ARmWvJr0WLW5RtunMq3lw4WV/R3m7Gbz9U7W5rjf
lBoOWnJ186X/P0h+jzySTbjxSVoqexmSq7I3BiunjaP98VzqEXjf0GEqgv7s1Txj
ak8l0XZ/srDQUFxT4V94HKxHYOhT2qNLidjPkdIGdhGuDMXYChmAOZ2dXC3m9UlO
uM7T9QkriHZFQ4rtqY1VGjvswO2wn2eqCvypFN3INSktJ9hfQtdVsWRubaJh52o7
w2LpE/4UcOJJWCkk8VJiZImL2mMDxYILtO4o58e/lGo9zTymoXqFtyrypqa96c/+
kkWa9xnrPNtZvtOu3Y5qnxT361Liq4deQroU9Tn6mgI+I0mnWPqNJpjsR9h8yqmt
xP/bjZBYh+zu7fJ38ApdkOM3ZrSGgUJhDjeciC5L4pXEIR4H45xYNCiMn4mTu1Ri
foHronBGIl9i70flDQbRjB1tyxFOj+LFAg7x9VIRNTSRxCcBrhqbfSM0QQQ1PBG3
806D3NlQvfxP04Cd2Rfzf3DwheaY3kqN5MNbOL0xUUS8ga8NYTy2ebNvfA63sZvd
vpI+pPWdUDPUooWpwU4/V9e48Q42YItK/JeDqH0GpdzfW9q6kxRORkDd4hwn6Eb1
crOQvsIKNe2YE8W1ijiMaX/lLDp6YMM6F3/6bXDO+AOmV+3Y++D3OtkgO3C0FQHF
Fb8AJKMFHGHUyxeTqiHSH6glCOOAWAFQzf348ha8VdgW+gZ62Cr+1TX2pENYMlmt
Cpq9uSSUwAFNdC2olcikMzF0KMbvU397L2nIThoKpiK4RW1NdoyvE/kx2ypy3wGG
qHYP6Da/WQ7ysa0Kfr+9j8297eGmfXhBLQz/EMZHF1yz4hpQe/2ewoT0flerIzHD
j+s2JCeScLtfefULvPTYffa/wTSIpy3tER2gAlUYnboaSOJz76gTKLbW9eCPDy51
DzYAPfjtl6/zNjT+p1MDlnRThftF/DkE5LRjVc9ypTSRMP5fQKSgyPfwBjkPnRVg
ujiGvg+YxB/BvbgD33PbqonuG52CyCo1XEu+48i+K9W32WaoXmIWrh5/32iF1ji/
ufcB39nkk7jyY5cOgZNVd9tGE84jhiOOXJxfEKBfEeEinzBfzXTLmsgFE5bz8gos
SNO7GkVe7uFof1DoAAiuGY5KU6FUQQ22J13IVb+iGlAGRq/9AhvIT3sc2YMXDa13
TFhPB7zcvsEpZvZQqVR9EzEn7jWJvOawwwkFXyrpj5fLLXzDJWr2wuSRHOLdtCld
ecYWxzg5mKkgBRFL943pIOrN8Qbrxt8zj4CIpF35Jqno7/pDnlzCF3KWYDTqZSK3
gNpLLQRB5SxMaQsoQSSTl4LepqeOKgi4qLCNIiv+gFyNENYA45YjFMoWRKsYDRYm
azRptHlWCBqA627ttIjmFtUMxcfz5RPDhh+gQUv01jJSVKZl+OkA5sSOxSePCbSi
lnIBlJciwmv1tdqowsN9W1iH8ksvyH/qv/acm+tI0+syd0YsuIq+s9QM9L2rTvuG
Eiud1hsA9HE4g4Sw3Rrt8HfuTj3iHlje3pZqML02LdNFui/EK7FG9qPfITagvyXX
0m3jeoYDS+C+qNZ03BKl3RW0aNcCxzNG3K2MAvvzidrDlgKhQG3TrdXwSdLhfZNi
Z7kQ2BEZsQ+Ptu89iyHIDhxquU8ZrNW62vXUeYCL6G+dyYAnvwngujbar+0xrdDa
5DX73zCX3tL4rAMwXKbauydpWHUTusbEctKPHYiKHZVKQkRzDOUf4WdrEXJilZuC
nuVKb96voJXv+9BbjlSp5AFAjzUGWP0kizXcZwfaTvNT2GTPOuuVW4mNDpuvd8kE
Fj/WXh8SW6zh4qbxq0+xDhvyKvEqbXO6z63Gg0juLB9pigiZU9P14JCHPWdNCnNx
oFoUkI5e0lPLMMh0EK6IuPIL55ueTj9ujRDCgY76GePVJMXq5Y2p9iBKGp1jfr88
lrmFlmMUef/mwkEvNeoNPH1MjPGXDsvdYPjDMuK/0L3yaXi4J1Z2Mg/1j+jpYOji
2jyC/U1gvZnZAhaEet8wVksOJsiwv0Ci0gjiFyqjE/2QFIpDpvJXLMgPeARvI4A4
Y2kFy4s+A9MSBgtIxAaDWjiKp3cQ7Oz3+tz1YZs5hJRpO3ldppWRkuABZ7r9z4yc
kumIrHyJRA0cHN0BdKpzE/abG8afJWcwGLRaU1Q7N2odxPpVhAsXJzgie9iQEjMf
u9yerZDMHnF0cX5acuC3u4z7t2EuB4Mn2hMazXJ3FxLpqFKgFYZeuube7PRpyFDQ
GGvgMfBQogDn+eFnEOLWpcVmvs+1juGQja9jbARQCeP4VWWqGNm9ozrF4nJQrU8o
jL1LTaL9hGcWDchkjas0lPb1WY53zc00yzabaych9r32JHAKN7PzwpnegfJd15P+
KkmigmswySOESG9TrWf7QmnxniQdUs6wxZkgl81qgk/8kpIC4oMw4jQ5GYBtMBZF
4F26gtUUuxd7KsZ+1w2MFytpKbbPynssTWYYWeJiHwAZy6n4ipmtbwLC1b1wERTP
zRo0ly0UpBPnj+wJZlwx2GJwmRhfRrB0fxgBmhiuqkwNsZUXUsOGKRyazFvTBjxt
gtxvwiQQe5XvwkV7Z+v/juU23KxTyN9+Nrfxj4ZP1sItwihjWeS7XxGkG80PNAdd
SEwzjtApDxz/7UgNnD1oeVv3i6AKeb/FPCTikT2OGpVE+S9lTAnLBW3g1BHNJY0g
YOk6ak8+K6/8YOSR7I//5ojQvHrSqUQbyPFwxYiLG9fcOvvtXQLojVcBD/eEIXru
zJwb8GYyV6XyXEAe9uS2jaUnf3fVf7y9WYQ7EMrVtwdOWdzYLydF3/6ilNCn0zJn
p5R9lIWjWyHSUkrmS64/TfVWiZT7BXh800nHhX241xErsq0k3y5YlMfTpGln8XgI
nmjZqpBNOGdSZ0P/uf2bx9EyE4B8qCEalGcdzAbAynnV/pkjrV3kBzx6vY7LLEa1
2IwC0C+xhBojlit/xk8C1c5Slp1v8ZiI6rbmlBKrZkG0SJXRi1MyOlcGbRDz5Bu2
3j9d/yu8ha3APDmTvGZUTHXeDhLst7NPebTsqLCuP6lyRtUyXSxZuTLjWHUJl1rv
C4MJdmZ5prSfzvHHCKWEoppfg9VUx+XL7z+qkD0T8xxT5cgb62iD3sg0DKrimqht
P6NewMnD5NhNAlFeqfbjWPSBufkFG/C4qk5Y6bd6prAerO+9qTefx+N8ResUwp6C
KPHwREjlSCAGwONWLv8LSFhZQ/YzG1BKmJiXdT49I+GLmjUDvg6slomx9NW1j3nS
MCx4eQmwpjybFzoiCxvYnS6RwL0yagev60SzxarE2TFa0I5acdBMVt6uY1f5Y/M3
uZhzeo/8uRovVOU/K13XB8RjANzkv5RJU18gPcyoGQ77qP7ll4mDP41W5YAjEjRN
urVvIeNO5jkIPuSs0i3MUVjtQv5lL3nbNHr4Zv05Wws+vjrg7oZMg32+Jh6ZfAQk
Qjji7q+RUqOoylYLdquq6n3im/4Re3WKoC/J7rxBTojg3tYpsBmrOM9ewInIgfG6
tHQP42eBZrauE4EZvJMWVQ8it9IalXxp7dd+8C8OSlVaFJT816vwqff/pL320CEz
chnZY4NSmqVWvSZgOtWd5LEidjqHNqobcKKGdDaLXFzONA+N4X5psrEc7Nxkj1RS
zv1eQplP378kJRfSSyOe5FQ8VXWcnAN8trz8QZ+tzk6LjN9YV3n537XjJNiB1NLy
jj/+1QNm1jIjEo81ChxyJmLUQ2Vgi9b/lAIYr1f0KarSmg6JfxtF6/9kC0B9OIkg
81ym/PnCE/yqAKOge7oL8eiASlkgOcr5hUMrUK4AE6if2E4RYktqE9DSYBP6Aa2Z
S4v4jI118QdRvIvsYDiN8GTmJhf/cyFbPeOJtrKJV2IyNoG2foXsGyJglPS4wOti
gt7II/jLS8m5YeRtW9DfW54rFNuj+qfx77yLofOxRZn+Sm7pMGZzlZTtkIhCwyL/
G/bTecD+C/pZksIkrOEMru1Sxi+HIIgklV81lizRT7GSw2+Xdyxyth8IQfp1ETa0
WSTl6kL8iVSn7ZgolUJU+Oq2mwV4FZEEGr5/E2B3o+Nt52y4U5qYLFP0s3Yg0Wds
CRV/8bU42xQwDq4WkFRb1mw/UhBqCwERrHf4QJEx37LAnTZJM6T/tNhw7v1do5dk
joc9lzhnWKngipCyX00DaCZLphGTrpyNf1D4daWdtOWmTi13+WJOXv9SQrJX6zj8
DAGCKbVWT5sVG8aUxowGmudfo429S7htDp5m1D03rbhuqJbUPAOotZa4l18iA5+y
YT0VMVorLCrMSAA+y5kWN1FScCGx5szBL+dA3hSQqjK/DkF83MnHQkUr37sVwBzY
r0IlpxOb44NqoE8FnAtXykalyO52r7aTBL5/1H4gWcVMGBy06YicXaFtdV6gnITd
fgbysKW3oRiW70psIL0NbFFSBNijiDue5NKivErYPRGm4czeGdB/Afp4UcAdX1kx
Y4Te7lv5PTHbeW2dj47JOaglQqS2c3wPlcXHVt7Kc1aKY8xICQy7grp1Br3X2Qee
imalzlar/AZfoP6FOcCRmALMlnw4nwUWmgrARVIkDXEwSSgLE9tAAYFujI99KA1y
noHMDI/luwgVTdRLdalbfB6SdJuURBsN3CFXR0jwdS8P02/ixHfYgmOQLkNSJq8f
pYHSAwayX7DevZWFBDDLEQSvFBZumwUPcnm9zHAmtgZOEer4UoMd249BRInVyiew
OmC7H+GB8gwYVIoRPM8IWjXt7D6xx5o2YUCKPn5VWirXhrWXDgs5oplahy9O8KG8
whF2COFsIEG2PWAQTgttAGuQT6f7AvGXRRtQJg+n46X8unDpCc5AuAcZ/mB/8V15
rO5evmt3a8zXMWthC8I2l8Hc5jwuJKpvpjY/X8Zjr97IRSNROjMcAltiajotH3re
ZUu1w2/AlT6mrh3itfOSscqA1t0sMQMaygVeSQqo8g0iIzwU17SzpmgPomXMf6oI
0zp278UBinpGQ5VB1KeITEeR4DfQ4Ec4BALcia/BM/w4NG9qOOaP7JwNm2as5e/w
JpPCGH4WTxvwAsOQmTnfAwtpN8ofIZCeJGX9l9fV2HnaSjtHfOrE5m2ZGcdyreRC
CJV4iDSgzZf3BeC5GRPJl2qfVusabPbwjCSN/VypQ//rQXT3+QejyHIxlD0yFjP3
0OCFaiUI9UuDssEuc/NKEHxzNKBs+7yLsrAKsGmmoYH+R03uqpqjfgiMZj0mRGtc
KPKHGPyJi9ZA6nDN0zjn9zKMK9SWnr+wvm88O/Jq1A9eSDANz9ZZ0yLywXNK77nT
Z25xPeXZzgAsSxO3RTB0lkN4omqdWUo2YOcmhNeNpZxZQwnP7d2ha2v2zzkfUdiq
O9K3HUK4Cg84dNDf6K9zXiDbaL729jQ1qXbj602/PyrGIO4S06u+yrQfFKbcNXPY
VDQSGDbVM9rywVWZp2dId6LI0pc16BeauztUl6moeFxQnquUQqbYJbAe4ueFSOKz
eUzVWZ1Qd21gfudlTKE5xGXs9d0hqvmPEu22G4v4frmUsMeE7aChcQpqZWuyT5lp
+5JFKlgqQffWBS/J3PzTEzoGvFEjUOgUub0S1EbRdeerZT+Xy9xWfl3gONzcEsTP
b0eOTrAD6PPS4EVIZUy7lXLIdvAJghFwcigAPqd8pl9CAkzQUWdiI+/yNfkmp9OJ
c0KWUd8NqWCZ1HxjMQPcN6WP8oxpwLDeK7rweXBEQ+mHZsag2fHaLW5XgxLwgWsp
QSVKUjGhPpoZVDcnaK7W4r9bfThzpmUAPllJPke8DfRct3WLC2Dmv7RGhcjxE2/4
fcE7u9iQnWH3DizqzMymUNHmSsUFOJTMBGSzzGYOvTWlQzeT5DyANuYioLIMTwMh
COQa5cAu2oKQvMe1nyMBEC4ypWwlCRn8TG3mUM8uPahypczGB7NVuc3NOnJ5i+W0
8aA3nbF5hPewhpEhUtMn7oH7Z7CF+2dXa9ujQMLgbYWEmTt0/1JVVqSxbB6w5Mus
N+LGvBc7Qjc4dMGXftOYB0SB+s8CktXPfJI3Q2Vgz4VDvYSseontHy2tIQpT0G7u
GfAsmtf6pD0gIHcrTbp9l9eAHdRcJjM6UC0TisfdI7aSdxM9YmNpx824xn4zlNQH
ZWdPzF7cBAuT6TQ7weVdhfsqYR9Mrdno28MF1XhE4981W6Mfof+BFG749Ta2zJBF
rjwmX0qGYoZPA0E1aM5tKBIPLDrYjTSs+ZI17vMdv35Lx5OmlcPmvqZYXps/027v
u5XSYc6RKfvdRNUdqSgkXofgefC/+HFF302Bjw/Z7vvILCTbu8b2Jq8Zs4Tf2XYl
VK6KkzoYGKmU41NXRtP8LgqF4S/rN1ygCWDx0Tf+9zhrogen8IlUguGsygtFzTxo
2cywdPh8DiwJAi99zWdbdzE5lkCSQ10yEOxpchf1J62kj2i+YSHOtyxfbAAivsTx
mDzUj6vf+dYLwVHkveuTR+i0Tj4+hGUe5jLtpyTa+cBoe6psTbM2uVGhdXZQY2Ol
hvnkTxsxuaZOHfBkxnu5m9cluLu/3A/n+ZHhYxH7awh/rLC26rN4B9NuuMP4YlOE
MFdhlOite615BK64RFK/TN+5Mh/w6/5A2wy8Vlcl5ArC2U04kcmZUW+tUaXdDdxU
yHxh7X5LGfukPcfd8b+3lkQTVHLrSANw9HkLDc2ICvUswAEyQvOjhIHuR0+8jtW2
K4wm30gmMloUDz0bzqEZBo6hzeWKR+FCr/+Nr5xP6gCXN9YB5uKj26IJR2v0UfD7
Th0pAr1n/mDABWCFAb7BEDw9eeqniOcFqVP+zF8iqW2TkFRXnNoD7P9R2dqv0xon
rN0/WYPiuteSxgaTxwgtLh97H/VkRq5+D8Wii9cuETLMtdlo0XF25dtarIow0XSg
DSCpGraU5dTKKDyyYettNvCv4pUQdIXn16ONNELErOR/Kjk+8pizD69EzvLPCS2l
Qh5Lk2TiouJpP2Offr1asL1FtzTYAKRMOCnrT7bABvNWbRZjPtFaDi0cSyMayyVM
aIdWez0p2gJDIc8UWQsFo2TPl+S55LVfRHAW3S4uXjvpAobFIPSYkhIioHbZPZdL
yXqIG7I+fGo6ezGYzzlqHbCn4/3FHQF3ybe5ZgQLokI6HRcu3PQ+2vqOGZxglT1n
rqTj46nJPIPPl2tSmfLnJWEPEVo+VhglDbNYSHYroiQ3UO12uruDa3JRxQL9C09t
9mG9/wBPGxWNPi4GNxtLW4FqlsXhORLtDhD3AvkpWZ7wbJfDij4zx8tr29xbTLv0
KabI+q8q9DWyi97eDAKdCoh7otEwNToZml/PQXF1+zyJ44pgOpjKdg5l/PH818kj
yyPxNYVK29EPWkycFRhZ5gash4ltGE/mXhJDDdIVZN0UHxnSDfYK1mEIeFrAuUMb
bI5zBoPGKzvtDDScKeFRlGvJxq0/+oPd4x2A0Um7gPprBQ2yRdKJ8+fGP0sjJX+p
pGG1KN3Sh5/jRQTD9C2JOcoNQ8eE8c5awUaScEjJzu6hBkXqa+eDRLy+JQWNzQZP
l+97rZD2CvPmwayxIyOGPnZIj/pKAOaO9aERyantPRm6PQ+M8Cqe3HDMXUW8R0VS
OnPe5JBacHEVUk+m1YeimIIHI/0g2CMX+NPrXStmDzyHyit9YNAo3OY0UEnpXMW1
Oe8rnzL/vrw+q7+Ss8aJCHEeVZk1f+AxhoQ7Dr/yZ9Fz1prn5lxFOIZ/JLIrk29c
4ii/PY/KANpJPDKzwUwj0gy9ZDYI8IS/n0XL0zQsK6V1qFhrVnk5DLlNj3dOIbvh
9waNw+cDb6KfkF3PJP0KvBR2uFqkqBWLufvVdhfnfqu/ny9aYm5g6lnHlF793EHN
DSj1zeAJOEQbbGTlRw0vcrSOK3f67Ga8o1RSCW8oQFbJiEUexTs6mKJvtdFMquxI
4kI3gWtmvCtB7GNGw57ENP0p82Rfu8PCasC+POLvrXACgABUxNJSupYQIzY/lkhD
RsfjHRvC3mjF/sZC7s2skQ8FXt5hB33n9JFUxMNh70r9wp4c3Svuca8CSfQJl3V2
lX1y4qOytjeSPGTQgm8RMhgdVPhN8zJ3XFkfPwXbrhWt8+rzbdfb6DqYwAFYnkdy
GSko5Dpe+U5JQBd33ebMhyr/8jDTNWuUmjBCL30o5krq3KqY5AT6TWwEoBOaJiPW
axEtn+r6bvBbsl0so9VTnqxCG8VvmOJrdAp4v2w/CgoBj3egCJ+h49NrGx9NZx0W
RqLT3Bksh2sU4L8XIHDURa8m9FqekUjH0sJ1n0ZXUrZjrydTbKMWilabWTmUFyxc
11kNfVawdVeADtwfU0JFrZKn6AFdWUevyPYnoCJcYCJHCbib0x3Ezpe+c2jkttCV
DaAyq5lElJl2D3/9tIsZKmbqlb3afR6rBmXJRqy/0IZO3EyxRjPdsemvrhVZhsTi
GYne/9muAnkiZ0caP0Voen487ySzoYH40OEAGXuKAHhzUJk2j48W/DlcWyQkcAgi
qmCJhIx1vv8K9LmRWxrY/XxeaLs/XIfxokoHarvLO4eW/EZgEd+NIGKLDBMhw3lx
NHM2mmSbFL23OjpFYoVf1HRgL+AT43Z1K1waLgGo101h0NcMGHxPaGLuPNrF14l+
khthIwCqOxSFVuOAllGG0/GSvqhxoMia4emREAmi50u/5ByIaykNMVNH6Hq/dD5T
Gm5C5JIXdOPnFL1vz1d4E92tdDq5oaMq5vYxPVYkzg2hsVcZeQ5PMJ3qN6CUOvX3
hcp5TaMj5SV5Pgtd/2gACcSwxP3S6xQG7hNi5sDFEjaRF4bPXflzEi5J/lTkgSdO
EsSIfvy1AKTLX9LPd+ObhflBgrJ13wA7LBNEXd1/+Tk1WGHauxmWiCXXjtljc38G
oRyrgETv0Uv6S+WGXEd+JjDNQqdliMM5lGIjIi+Zxb9z8iVXPeA8cXyDi+D/5yi3
1Or3Y/eS2O8u6KDDXWk5LMHKooi0+BZwwRzDFicjpiqRrsvUUB18mQuoFSEzdqKW
f4XCqkX5ovoALQ8lLH++7RW6sRgT7eBr7Vqh58zlEA2jH9nm7fKcXKukKhWYJ8PA
/wPajezy8EHcw9bY97nx5/WOQGiGDcFD5vNB95LbvaBE2vuCaiBpo2kFv5qG6Q10
oIlyz6/baWu5CMTAus7CnJZuvK5DUzCHZum5XyJqDOL8BHSOugBSTHRZgHZmagtb
mKmnwaRjKeh+AygJHndm1AXFUwnnbR+WlZgbJU2RWWoo43PaNU5eNFQrRIFJXhkw
95junI/SKfp71xpFp6Voch7wyyI9J69/07PqogcUKRBzNMzN8i3oLZQADgKOop6R
UrwKJkq07VOxwRxsT+nlbgzUTRrLltovhfgrisuvd09UwFK1QOVLbVFQA8O/j1XL
a8lSkHg/jeRRrf33IStEg0CEL3BWuidlN/K5IxOrHqmgRgQc6jpXNE7kgMur9XE7
QShw/TNmrVEJQXM385bkl3napNmMsy+wGFI80zo84QI40GHso3q7FC4jJMBkEyof
SWOmoHQWIZrDWY2wTcnQIv4t/KOx3AqQ1BNq8FD6pW8GzweuXcZYrxxccrgjeJ1N
EkWAJjoIVHbt3DnnbFPqK9smqc3ZQtx/heLPAy1jn9x8moEafo/t9LVOLBegm6nh
lWTDhBNGU8XtTa9F4oNda2RhqpfTElw561T8Kco5YmFeC5zoJjMjHIXcwVB+Fa4h
hj42s5USJ8nq3NtEC4g5VY8Tfo3bpgIIp3g+rolmHVien3lAhsc9qeRm7M4VR0f6
atQ8ZbWqdfwLBBmJ0LMS3JwcT1mQ5W2PvR9UX/k/O8mGpLeZ581HtV7hy1Sa4V6p
g0BXmw0yD9DCTAVytx0Px4bxTr9k1HNTubeV3tIe88aIe6aKJXUzrysibhzslS89
ABOX41kyUKg0uqq5JGqkZnX+Kio14Ssx2yJor4Vs/6zkBtaGugIMVbdD0P35VbpI
oQFP3DE3l3fjri87hrWXGo7UZZ775F/IATaz5RSM/c6PfIiWguk/DY5A2Ef0L3gD
3Y7+Uu14qpZMJUDTY9IovDjWFowgwN3TkZI1fNyFpzvO5drEkmvtbxRS41yRwpba
cWY6nTHuZxiR+tB6VQiGbbW6pEBnqu4sak0rsIQ8tW9jlozbPhkrCUwezcBJTb70
JeE+cMuC1Rgqo80UcCVJqxMl48ozstuT+gBnKziAQxzxhgy6+kcIVrgSRGVZryCZ
BLGgeQiU13hSHiutA4gl36JD3xUF+U1JwG3D3Ud08AvjCpgZbh4MKEjdGJnsmIfn
IpJnOvrcaVsHaKtsU9IqME+VNOWenTQMMHVAUa/PLmjhVUlTOqJPqdOZ0t3cOQPp
LCMAaEmlQVul6dUcRRbH3KK2dy2OjcggUujtA+EOEhb/S73NKGKQnwm7P/vHFMDE
Q7ESVVllHEbPcIyzz/Jtgp6ripmvo2BpKGkTuQDMh6IdSFH/DubEKxIEHtMBChlv
IjmzIaciU49O2+mEdCTtyM5cj3ot3CpkNwRbB67brTeWz2YZ3f2Pg1qL8Wc3aiJF
CWYuOOzK2o2JJO/ACJquN/RbPPiYzlD1p8pett2Nje7kpPzVoziCaA/Yrr7v/ER1
u1N3Y5rvVfLlP3o6+HHPlHoiMSZD5eWgTx5MzOQbfXhUBvAmzwUnlulrob/wGiq2
hUQEI3aSryjvnnqtr7S5CYnArs9glBAdqJUMHv0MKJWPci95kLcqKL4SUAzPXKbp
1LDKeL7ElZnfR9r9ZD50cOYF60+OwLcXjp3APMUgdk12VZlICqPFN65IjcNXZi++
XeG8HUlHLR28gYjh188OqZJBk9ZgueOCA41Yldr82htJfMM8Jm9i1yUc67uvMTrf
i0C0LcJKXuinKyJXukES1zWoz6UpqmuT2Q+eALh5xJSdlCZQbRC4EccDiKlJ2RE8
CZ5ViMy94kgHq26uyeDt0sucMJNKu5AXJ70rd5BCdngoe4fQDpMnAFiHJ6kXp84U
rE88FIgdI9btAH0HKYsW0RLixpID2rkXBNyVMEM5MlGUxv62dVKjqCbXM6w2GqeK
usvi8jJZV2iF7ov8NJUWYXJERG6arbL58ktvtoqsuULfjuAtClqCYrzDcaJgj68q
IDmlOmeLyReSH0jvnoImy+goykR2c6KJUBKdn6fPBGVz6VIO2bAdsRV6Sp7M0af4
0dnvy/o/xKcscD+3bzUMyvivqOLPORr2GO8RjCq8Gt+YKV2TDFASfsSC5PS9QVgi
nsCyco0B/16c5jjgKPwecDlv8SxJb+neNAA1L5xTLsGESVNztrW8FINnwL7lDeH9
xoTxfJmILMR+jLzNADO6nK7fqXEjwBcEk9AuDl/e+b+62RKLMhkk2s48Oc/4eYw+
iwp9dHNg05JOB42la7HQrFYKAQiyoVTvwpcZ8ysbykGi6uaHGcUp27J01QZRpCi2
PWWpt+qfijcGnlJrhp2J45zakPFCofMIWW61kUXnxVlG7cgK/BAxUrQh3ge4T5N2
zGgTnEX3yJfooUBMwyBh0ruaXEem8LpZWGJbHjjmTUWwHPxspDBOClYk2GQftV2e
dhAkSG5YphyviA6zcTsF4v1wQrGRmkOYlHw7Rr2iqZ1JD8lzSUV39RxpuRtrBRZn
dNykERXAKsoakGPoMamwQpKH5rpHiDIZ4iNRhpAjIzKi56181oHYGshQvE1ds/Qm
OmEoLoTbkr+eAnkxS/6d2y/t/op0JsG87NzMvUTYWWZHj144/OIYeoo9dzMruRlx
3kJ+oMfOhEV9lZKOmSpAZLKAl1hbvvr2B0wgXiCN8rDZGjviRZdoTjxFTR0f5cIV
stBLA3JN3XZ9t1Zc2+VK1Om3Syvp9SqI2+lAsMisDvCBVxiKQrS9FsKdssq1psBl
1BEl+EbD9L1rRHqy6qlo2ZRowDSvy2Wx8PJwQopMNMGTqJZ1L6OOSvkEm+kOjO6A
AvDSzACLwXbCd49ZCPySfJnyYakCDj1PNdb80kP5b87ql6w0Pg9Ets7hj+pT2P44
c94g82NjFNVYzcFu8PaGH436mhtbYtWXIlKIAHfJ7OpYOKHB6AWRZ0rxWAdTY7yb
mjelFbj8WBQ1supfktxPcEXZnoG9Y98mSH1I6H+ZGAGPg9PkkxR0WpPoU8fzd7lD
A3GGaX8AaKmLjYkROZSN59rA0UfX7TE3T0NkUu4/7A73DodL+gzru+YSLQ1KLunf
vphmRY9/5pOI16a3rxYnKta8jau2Gj6Sf//XSniJwCdEiXjKn2anpUgSOBq+SnTG
0DGxq48LK1Tw2hgihQzw4HKb/+IHd0bbQqXm+WGH9X1kZiv3AjVqltG78ZbNyh2e
/FKgNHrBUw74JH6MzOwlG4wd0si1a44Xu/T9TOYE02M94/reOFo6ioyuOq1zpUMm
xq31wvtHDDtX4xqLMccd1nSXyNSNW8S8qsXg/CC08XclEX0vRM/MSqmDo7HGqbOf
fsW0EMWVhsO/Z68KD/qKj0eenqjXmh8SHq6TTqCtFIoPNwXQMBL6+5sRJcmIQ9eo
f+JkgDZH7igJxZccX90SgxGDBr5O4Mf8jXm5cDU58H02mzPA/4CelAWj8ddMa7Tb
pWyNue6VhHklELBDSpbOW+Ovhw0r9A2HYTHAQplxX14pr6LTeCEQ+MPj53cWVS1k
ZL94dWvXO9wyp4i1z2/4zhkggN4N53kgR6jOzP2H7fnpYwtH4xqs9jTPyYXmSUgb
urjt/7WL1U/xaO/LOhOUM0yu6J76bzmVqBhLnH06vVBMm8bM2t7ZYXIw2eUjgoLM
vaXXdpQ99bChZVIwk+u53bzzcD0cP8qwbDahMivRbR6RrAB+EehvoGLOcK1OddP+
jp6j+3eNuuxyqeRU7t4P22eix8gDAwbVqQc+lcGQoc88UsdXYoDHMimQFCVdLG4s
7vMt9tVZGyBsHwdCwivVNO2JSinGUP9agdOvk5EC2CJqVGLoapelaputDLnNdcEF
purIHQrEhcmUNm7hHzHduyZcs4Ybb4L+JIuI8M5g4pOIdn62T5Vi/RjOlaBTBEwo
pVZ9YCFqtBU3LNFQQ99FDN6HHIwwPit3vXvKTLLO3ywYGuW9MuULNwdJdWnkHYvb
OUIN2fKpXCtMsB6Mxqxk9h/42rqKVxqx93a1xi+Z3ZBV9d241CDkU7sUw0w3MTch
c5YOyI790ZGdpzHtVXY//8C/qCAPXOsrpTYl6a6QOmAem2Wow5Ahx2cT3y83gjo3
Q2LjyPcCUy6DEA8rZ4I+VHtxOePA425f8YsDiVjXOizOC3B86F7hfV8sfNhAbkmZ
vB9DiPPOTh6Kux6NkqUsVdDQex3R9AuWQKfGmA4RrU4VYdETzr24w+bx0tvCSOt8
LqSguxUfRBAN8GFiyA24YqKwglw/JXc8wnt+qhEcBd8nwaW+x/bzXCgtNzUpRnhy
jY7YfxJMRbJSDPPId5rfOqZR2hw8MrI0O8FMEblpPPWf8AF0jau/kJ75awzIssZf
hP4G5kBsn8YU6vPKr6LFzLo2Xn7ygN1+GCim8/pGpD4C1E/rFV6bbt6wxIR0/KCG
BsrFSj7yq39gtT/Uj721tKwi7ImULFLRhDyn9GxuQgjjgnjgVn1PZQiDK4QdQbJL
vWkoM3+hyHD9d4ULff274vEzxjR7OVnYNBzLA6r8dkhZxDcfUrkCUGreTyFVe26E
HMa9B5092vlOQrsstDJjpLp/iVeegpDxosXvDnoWGw9HT5yx+melLMUYv1Yj5PiU
bUJn2ETwkdmGd/wbAtkPpN1sqzDZHTp0mP4pOhztZQcqV0R444ojpsJ69OfavuZy
IsStiMJDjkA7MykIVRzchIzE3gvxo37lBm0kcb+tAFMgCuDY1KDyxVkEv8tKUIKH
Gc3PSPiIUALrlvyGFYUyDwnZswQFd2kvOVxJYIHTQdbQIYAaChniAVdaXcF7U9d3
yg17oNkS0Qq/UxAvhFAUuX6PimC9fU0rNHqW64IJchWKbSSA/rZtUDlW12BJRG8s
qpOP7abi3BF9cH61omX0AM2/Le7GtUN9Ie9RI8z5jkKzXPZORfyjZkGm5J+9bFUM
csw1rI69ZeK93mxp/HXGQ4i6eMEoFyQG2xPMQZAQA9BP6HDIZpcOoDWjXgMEi26s
9zdT8bjDjHfpVz7UFeh/3VwVEINIFdn2G4iTWKHCe2WHS5ArCmzwRxfXwio2r/rA
vAJ+20F+UX7Qb1KLmu+huWLGZqlMp2Vv6MQuO1Re5/2ti+/Mmp51TsQt7nyg6E/k
9Q1jiD+vvpog/jElFLwfwtEnqNzOU01tA0iN8m++GypnemVF2C//lFTv2l/od2jq
oJ6f9Z8O7EeNCX7eooieDmND8taRLoiGz7h5gEH4DudN15NTPM57tTHq2FSNhzSF
w+7nwqLqnDZ8Q9xv3wSyROu2JsDD5AObGVaiaD8QVGCxOAKRXZKdwcyqJ+rkhpCa
m5vRChdfnO5/7cGEA6PKjlRUWCbOCwNKVHhV5L/njtFg8+u0GEyTEDWFbaFlb4ai
x7pUIw2KI/JO/m0GEnMVcsUMnFj4DRqLJWB4WvxJ1V8+P2qq3hiJriyiPbefLzsJ
8ZikNQlWhCTLBdOJFD/gjNQrNoOvkEe0MI9GUZs01lMzQ7p3/+i4fBQi/St97aOc
EjC/n4TePVCwftX+hWXGscwSO8EMEYyPobeE+SvsV40kiMhEGswJkffz371bu7cB
M6ikqa3seIM3SDWTdvhdDox/ef+zD7Nk3hRKYPcVMaCXuGtzYIehgzVHzDIJoKSA
GQP4B6sXD59RbM886ysNBGtjCOGIKSlSs9Wvh9WOYh4Xszb/kf6hwezef1Clh2sk
RxpFQeqOgedouOjEQ1MSfrIpxmeNaOBfDu/Hv6q+4oqg1VRfuMYDVugPsP+iaPV9
b9JZaXBpeYde8S92xgrlPJmLQOQUJfiGWpX98DV9QQFlF/9JWC4j4fqynuj7kScV
dsNWmWNwrCopy6FXud+CZI7rG8jTAkvt4S+n/1Th2sf4dps43h3FSEzKaEBj6+bm
/rj6m2ot5SMmE5CL2RiSx0/3CXoh5fC/jtpm4/zVB40DPDa50rFR2HPa9PoWwCnG
lYNooMT7QVL+4/X+hsDjjrHQOuxuTZ5qbJod0krm+E+cO6gZvrau3vkDa8HSzh4q
BFbog1OUzphzlQJaV7oafLQnMzitJLoB9OgEeTnm3NB3RHlpdskyw6l04lbFawmx
iwID7QLGIPle2D/A9ElUoudPkpZC76NqKo+C6WxgdpdNIQl1dGrVDcguzwkWGXf+
3B4S/nsXkursFPrbi8HIx27DyqDO/h3XXOHWfqxaanuUYOkUEK1++bQb25nsxXkw
74jSAw2LfZRoZXBn4gRAeUGx6G39ppr1ZPmsxlwwk7ZkmmCwahq1a5stOMzRSqjr
NK9zzsu1aFp6OoWr26ctVzNNZDPnQRfPTGfFBbwsiOk38Aa/kOss8v4VDJL7o+yO
sJdG9mAzpGoVqMtrdFd0gMSRvh6FiH1Kp3AP0YAlxryejbyA39hbfF2IQENJwz4A
mY/hijLuHrFqw4pZPvE2CIEj0s1GVXC5ePhKmhP0cdF+0BviL6LC7yUlid5sas/Z
bJ1NErYNhMOJ7t2SU0/AkbAibxkxuzh+ZbBsURqCYkttpH1ey64WRFQY6mO+UghI
rStFRUJVkAZ+PwAuCNA4ciPTuWBoe4rsjdc2dlnyinQR37x5totmf4fPE5higGGO
Rnk0EHCGrRva2uxzGEfzExWvK5x/R7vYi5e5Yi1yD8fMon6jshH8WG8z1tITJmBB
yfBLJTeJtlnV2NtxjALkrERb6eHHMb0g87yN5ATsEtylluq/+liRAio+sCsFBcrO
gmtWoGFX/MygcDS+qleI6gkMty8ePX7FaTaizv62VtXXLNIZ6Gr3UjeopidRWz6A
w0/V/AkyEJF99tKPWbNI7auaVyxASuv5dlWBCKqsCCMqWAN5vZ78UvAvZLJE9A6i
Uq8qjCXW3GE3oVyJ3ST1CPdF79E8HYxYMLg/9qutA0Vye2h+stD5sq7wLQJHzSHj
O95gxqAxpdkaS1G5n5iu+6GMOGXfZ3ywYXIoYIv38d4sLpusPdXGmCaXW7JLZ4Mf
uk48VpbO4XugcDyciYQI/vDb8ZKzEpYZAQ02DtfDiL7SExtBxhXHG3tD+5A6ATS7
wEs1V8KdoWs3Eb4GYjhI/kpBua6Ef9Hi7p/mHhblLVjFtmR1GJJomgZKjGaWjJF5
Aq+kc9PZXPVNe9cbmHb4rarC8O45SKviN5SpickwzHtmnTPgLzcLGoh+9gj1BQ64
wRT1olDTFLa2PPhXZVU2QUmGrto9eB6K2pgFp3OsHCM5g8dlxkvuq3MUR6yI02sY
qpu4cOWuf/UCG2It9wGBHE1LrK81+itcZJ1UuBTz0imgWRbwuTdFHmCaKiTtg5su
Lv1D9uefZy3CspJjW6hMYRGkF37lBAJyAMdU9f+9+OctFDaylNVywFlL6v1IF+T7
O3k8LDV4aiDrDeHjDxDGB1XnVeQLdbXxIZiNDSYFxCtUXjxxdbSmEXK7fU6UrYWq
aAVd0Q+otT0cU6Jw5C9n8X0Cz58xKREG/72Ip+N2CbLyfklsHwcpEAPw40tldOEP
MC2gCSjaYPelYM7PuM0YsN7Hj/S/WhVsIHE88+alP0UIBIfW+yyqNGNejiF01Cmj
msOFb3El5zXEMQV5E3M+l3Hqcuu+lXm/sl8NFkTjwCOqD6D5pWGynqH4xVRF/HCK
r7/yTPtKxuLNrzt6I1REYtmBkcRJWQ1WxRv1wbVujAaoU3ArwouWu5RsEJGBZLup
pV9MFex+hu3TBV0iGOwvUt65FnlFVozrQSjxen3LXPFUhEmcx8lm+2ZJEVZ/fhvN
vf5mWsZHrXSpteF2oNPOWxRUN6iBN1WVnXCsZEMpnfGe9vdZszua74l2IM+TJ8vC
ujKXLG5pwI3VmI4omEBot7CApboh5mOZHtU3x/qGhV2gTaOY3/hHxOsAP+n3gYLz
LDHZm4YKhQiIGZrzJqeMkaYt7Qp2MqLzDbB5GjAZhXDJf3i8Zzdf0ZQrU8voIkam
MfKhVdeKuS8C0kEeRAFo4eHx93LBuwtl5e+dysnbFD7PXsO4YWfB56KHry49aO7l
a0hmSNyigAxgywAWh6aTwiUulmhpmfQSKdMGUIJgNMUYfXUR09gwSFQ7pfOdkHyv
t+v1XUSMHdZrfOdLTpgRHCGMxq841bUYPb32dJIvQlrKQ2I5OZNTW6yxO7OzqNIk
15q3eo0kpTtHtAhd30wjs9K35Q5A+3XwQRSAJjZ1jIdDrKJNy4/U6TTE6Bpk+uxc
CD5LJ3wWsQ26iKY1DWuEF63kCoJWaYbmHtaglCQS6tn0uz6FK+We2pNXVW4fL7lY
FRl0pUM/mRDGCkRdugj3ubOWeJe3wtRgGuJewx2AwvFjiODCNSOav9pBC54TdhoR
rDP/diay5JGr3T+0cDKa0G5Nb8h+B2XET2o11VEyg+IuNiQn+G0yY3eY5uvcUCyt
HeH0HDy3qz37vLnhaa88MTVG/Skvk0sloFGbSYyU17JxZt93suKLWCSalJG/sleb
Qa5YwPyeOOopg4ZCn5PrycGlwiZ9RIyIedafrSnny7H8waY2I53XuKXanrNjx3yt
xSBps+SlVW8atZl435/lzcYP8lwipWHCWYi8PZR9kqu+v6ZHAJ0X4t7AzTgi4jxT
zF7hMAbvEcsB98EKkbTY9cGirpDH/m8UHozxs/pDg2taUjWn78L3ZObsladau9Zl
AROQ/YrmnSWfebVURQpHOiNKIUtFXXAvO7LIFgoK6zWHfPgKwwXunYu7DgxOAyzR
GMvVLQ6uT4E/lGeiq5dMil+JOyyUb2M+AiQC+umkH1oxP6eqRR/8NiqH4TT+iOb2
ZChzpkkoQwPfEm+eJKFSmeoZsf2CE6mHabFsraJLrbdC81ewfmAWdRb/MlowQYNC
eobMjQ328nbnQCDCSifa8kQ3zmDN2K85X46xZAAHLcnPKvP12d6RO7yU4rHHn4Ub
vo09cla6CsBs4UHHzFKkerYZyKXLa0Z3cl6gSWmBY8gjTX+zw6v7YKQI+E5b3k9G
qhJyE47OZcyE1JCXMfmR27uc6fwNet2ejgSkzGHKaUxFnqEsc8v5j84SOkcTMEgp
O+KnWrpr5oM2IP//xIoyRidruvtA/DSGbs247AACGvsbM959QjPVtlN+LPzaWQUl
tXsAPXk3BHRnGFeKKSBSDo5odyWG7QChHGxL3DlA51qZMuhBeaIsAMz1TfMysHIX
h5PkPvIq07viQp8kHU5ca0CFM+eK3qdfxLPFV4ECwAEBc18J1+meXRCwNPtr8/5P
fFVYGtUqx8tMoG3vjm1U3IMk1hzwguTukt0DkMriW/cojdGSyoylg9VTEJgV4sBJ
VW205TQNGFYCSIY4TuZXjjvyKXgcmEsiYN+46+V/CA5j5SZCaMFtpTHmqBKfZBfP
aFV7MvhbkystEc0Z4aYMrQPef7KVeFS2HSFcXxXc4UctDKI7ElPvCuyCmvxZjqeL
1IZSJtOAvg0YYjzYw1tgaeVFSObBijsbbGBF9fEPslCWX1evv2n79LMradi7wXNq
Q1Xe3GYWDtusFpIl/skK3A4HhRlSGPhSVyT7u8MRIEiW+yLCnrak1GIipaVs2Rp6
rLl9Ok1y0aKjelPW9jf9TSt7K2R+XO5MEbXwryPLkMglYTUzlcFW+YeO8xFoIGhL
dLE2ud1bhHIPtZmyv0s+EWm6EPxdl7FgBginVqkiXpNJWqWQyri03+hGEh2cHgyL
eiWoQD1JMnwmqRp4PXbrcbzKE3xgBJrhk4ky41JbRo5DGWdIE1gdH7nSGgw5UF7x
c0esgbl4wzSoseBRbP/urknVX7TqPAYcewRlskWLuXSiF3VvmHE4YXU6Nf16DV8b
aZIDWUDG0ElVXefqXl4ktu1mRozf7j9Bm7oi1e0ymV5vsabOz1ns4LAc2DkpuID4
qYkq1z7BFLQ04zE76GKTgyEYaqGa/zRn0vK/aF4gk+MXigHgFZn8vf9HEQRGBkba
MDP/zT094fdKTLck8++4D6+d4J+zWZw6D5hB5S6YhRjbY1chmSlmMkr5nGi0HrqJ
Fpt7JTQWVYx4wVPNh/t4sPoSVhQrKODYNTbm7kXbLSqPW85wmOwJQuyvtfezEmoq
Xu6rWy5DUAm1n63/2MDn0vWduo6etv9hfZ1W2+Gb5J4Aal4ZpRQCRkDLf/jgNOTQ
qaNE1wTYAkFlAk779DLI02zOfJxG7WljYd+04XhJtYzGzvjibxFAlQH2kwb0F8DV
m/gVfb6zPAqoeH+W8aRC0gfa727Nn7onFWwoZCrcm80uefD0CHZNtmydgSz6/Bdg
FvoxElugPP9IIFIS7Qy8zxTO4EhIqquLOFG1M8teEFXuDfQLVcsnYnmD67Y/F8YD
+IBOHCU4KbRBn2Af9Fz280rR1eePKDu9itgNwqPynio0Wm3hzCWW4/jzhSTrScgf
UIl9mp0K5c3ovxXhsZCvtCzcQQZqm7pWnh0Prs00cA19UPwlzeYIJrXsccXyiSMH
kojX9OH2rBG/8ho2nFlYlPIAGSd1H1AlwzWcH2OL/r1jSyH5qWxext/+OQZXPiyA
6mpHuvR11zYjl/R6R5DEAmN79EldJIBJWeLwlGjfGZnbfAoWM01tWGtaBx7j688e
H4JrVrnAXVg9RQLUXQU3m9dl1kJU2AbUdxQXVIsK2Nyh5akbJk8ExqPksE8AqMif
7h3OEsVGy1WbHvKHAaB0GU8fmU8pdG5TQrKoNOTD7zAahYL0iDzEzQq5xZEibyLq
ZiGEMVYRCw0O6IysEinSACivfIinum5mF7I2YW+ZWARILz1o1lEgtlRbC2AXQO+Q
KU7wLnL21g2JufdMpFojL5iNhQKGWeFWwW1GuFDtQKpnXL2NvfPEs3Onjhkogtz0
bO0rw/XWwfCojojdgEWlLAnaZEYaFkv4nfxodwTjBoKlm++qNodOhZgHAv78e+95
qg9WDjJ9FEc/I2cEH27rv57YrtlF1SZopp8oAdCnOFQsNP7lEv7y9GFJrjRxsEBw
sgD1E7s3ZRJvPoAyUhiWimKiBEHayTZXrIgPXluiKIvNVtkfYNaP0zzhP+2PX8F5
ezrvd5LV10m59OdoHNBBKzS9dv1KcUUootu70JjX+vz1lUc+h0fcxstXyhPfIC/z
7MKFrVg9WX9jOEg+nkBqU1lvFfvV5UwGpfkApj5+DGVQcB/838sGRU316KpJAh82
n/GHWKK/iz7wTxMOPERFOi2wsOIGM/1hag8QI1ZNJgxsDTd7NuOqtrqbOtEjsC+7
uPvR7mr6tzVSSyK/2rDwjLenruGauPjuOUHttPDEniL3ltYp2um1KOuUVKZQTDfn
GjMJevb0V6nV9bx7S9IzkWzv3y9P5PtfDB2CEj8hlL4nO6cgWTPcaeEnbJd44vN4
/2z4lnd1HluvZH4vZuE/YNdLp02dxwmza/A9MCx+5QhVLky5rEqkHFkiXNtr1EEI
COET+Q4wdNMq23nJ4mM0mxMS9XyEHKVfoxXjqLctCQWg8XrGzhwh0ha4t8dLDwW7
Xe8fElX+DBZhWyZN4eogoECfVW/K0KOo3eRLpRMwlIi3uw52UO1oSkIqmm4Y/XHL
NNdwnOLsGfuRi8p9hac33kynvuh3y1l6wVzy00cYuSxyqdZEItvIAvzswafASA2W
F9R1MFFHd8/3WKmJHLLmWbfPyq4qhFB0/UhGTPMsZrVKM5mmPqYgaZp7GSi8pJWm
knOTkPEiTfWTtzO2mI3WfihE5/KhV0jQ9UofEwqxqwG85WkSBVHcTOaDQTLdYT9R
smbB/hiWUBpvPguRnmO+xVzSECbB3Mm2yMCS4fsdqARx/pKsA5ZJj11sfCHDyyjS
zJZacob415kVDjn6YM57b2ZDimxVMbmo/MufW8C/6F5smi60OtRVdcWkjdvNKXK+
cYmcsIIEf6xOvS+hGZUueg4nV8W8aQ44+zQoVt/Or+SPUWuy7MklGLHDafqbdGkY
/lYjr2lRP5v7tsSPASnuFfax9vzqERKaXzg9MHtr6UDI73yLUb0BVlGWOFg+i5VS
otRWt54J2yBR4HLmLe3YZ+2irTbd5UNFLsYG66g2nEDw4e1Zk4VM20cifLag2GMo
T8YzTPjkOuXMik9ZhYcTC7KesXHf5kJIXKmB7uD+GTWpWNqauQL61F4h2lHXhdr8
EOtEpwBso1y4jh6nh4uZYruGN1mTj1yu7twe3Nf1THi8tci2F4UEcYIZmfNowgDg
46qWMee5LqwZID9aWxqXUtEJs/9K4wcDR//Y5RzO2JYW+NiUk5Ti9SgUvrGwHOUr
vnuYZw/kgIPBYZ2dzry7qnp92DqTo6YBetuU1RdGps6S73ahVlGhgiIQ4y6vRf62
yuTE8nylyyCSO6zw7tjhzA5DhvslQx2HVo/TFXSbItKt5Mw2i9pMhWYdG0LNVRP6
thbMHyz80PaAcaAINlD1F/YvijC9udQyTe+dIwrzqL4U/Pmzpvf0qFyfhZa4pvdV
o2VcOTlgvnOc4o6QEQa15MhZ86m+aac4eUgrTSgBZre+DySrEJOrEN3FGiIcBLXk
wWrhxyxe2kSMlpx650sG4lOImsidXCmBw/TV1g2CNh9lFC9I6U0gzbB8xCQg7xfB
wiVd0hA+7rrOEDbxCJ5mJgsBExYOgUhQQOcgzVOa7HlzlGS06+5BfwUSdBwXIjSY
1RD4YdwOov8+BPMNWJ2bISeQ+mX7xRyDL6Vf6zku13eP4Y3M0HFy36l6SBG3ipjo
5Zfi4loF6C6LyP/RxLIClVMT0cKPEPVSbHA4PaOAVPZCmFGB0g88mzYuYTHRlmYc
e64tkiUWFlyNxLQZGNS98cNVGqOkufcGBcZBEVvuY+ITQLWcnzNcw0RMcsqE01JH
qS2rJum8oRMbmuYT68bkUvIvFTtxrTLZ5Do4cKhyD+38LIb/FZno85ZdtCvyIE2f
luaJe3HoBT3I9VJXwpoEUlWaQWYbaUeJWQ06Sew3gOi1GbfMobRXb8gvGFwT6+1Q
AomW9672cZMy6yymAW8YcnWfCIj+4y6hgIS8hTVdtifI6DPFt7cj7zA7IV7ZGDRO
bxq2KXYK7IJ8ZACzQa/jTybhe1TzueLdBHeIyFFVaVb7KOhgK99yU+TCwWgvYYgO
U9C3c7m9LHZdIoF3uSynfrbmrgXGkjL3Czkfe30YShE+7JA7cwhA3aPCp4Yjex5e
4ib9i0kl3aUyq98vwZsEjhxoVBZ5EHaWC5dJyyx0MKn1GAnmyPOZLBsMTbZLQHbs
dBEccNc0bs1Z5WKK+LaBm3baDUEINv11fJEzQgkiZ3LXsABu7eI+IFIlZ1N33KCD
Sz1NhMJYiuEsoHu8KLP7MZHq2QZ4WRr959zKGqlWZxbmT1BEpt8uktiA0gCLyR0/
WJjYegT56j34EnZ2NOLFQdE6P91HBOj0mxED/yR+s92YTcKJ8qczlSucYj/hBsCb
Iu8t+eexN6kR0zxEdf1o82FQMM2kDXv+vCMMUIEwAlqcibE4/p8UUO9Y/wszOTkD
pMC/y/o0fTOat2Eu4VYxBOX4JhQmkODZl5VTlYDlIjVAnS24wnpEEN15uVKUsdoF
2ID90O8lwh6yyaOxvXx3nenA+qs0h3cCGOVeyqlHV44Kekn3hkgA4P4gVgypX9/v
g4YK1K7aCBvHg8aB41EqD/MfxCnvlLDHZ0mBYi7iZcTZk4XgdlTgZnULgGZDulRI
lO8/cImpr47ZDeriits9PjQ4cxSUDloyv08v39KsEXl7MITCZBlm7vQD+K5c7vvS
F2LchSWCrUtDqpV7f/uP7+/C4CZ2Ir9LBlVZlCJe2ARYzbCpx/wBVNwAQf9Y7ANk
LPT1GyKKholk5NN6LLa56sxmHVKnPyYZk7XyuGwTvIE/waMsPpNkRz+CFs7AFPbR
OTGDXQolGxrRbP1tpzt84k++BrpEPy391pBXBKVzSVybsHmsqHxZfPpQdfCLIO3q
0ct4ssdzXiyekrRKyRNRotaRr6if0WQNKkkffv4RiQ5Ruhf44zLScLP5zjaaiEZW
WAnwbad2il8tk8SWq+CUfI3XGG7dESJpy5MSx0Vgu6FCn/bF4IS2+qAOezwhn5Il
6KT3+0dYsEJ7pE7ovJzRVj2wmTYZXxqqPhy5oL4Y5Xin5z9iEymlDVNJ0aoHlgBk
+aIJUkV/NyVVIsJ865KE3YjEldUVLTDbGxFDmQLKZCi/FxMM4Muw7kCgCK31usXU
4N5axYx1deyQx0QlOK3ajaI0ZDs0fAi5KFRKKf5Vnq1EL3L2R19GA6+bJRKm1zpV
WFfoA0719l91nOXXVmQcILabcKaEDAwWKcRdZq0Kj47DsH2wd60L2SQgSQMWklmC
4hgu03WHJeXfiphVdH2w306JJGjA6RQZE6Vhf+vZ86+LaRN+ODJyKhL/nPVoqxNG
YsxovBFAacWJMgxTKutngmCB3oNQQlDIMrc/oWNCJY8G8AS3QwfN/3J2e12FsFv5
2dtipKbmCRv8rpJ0nIRs27EqRb/5vy+5j0vqp5P0BQet2lPjIcw8BuSGylj7FXox
SPfqXVbB7tQdVKTb/p2geS53X7j5m3eD6qaJ0+onWarXQKXZ5yn3M2jP2K9hUy3K
Z7zFNJK14tzShmSa4Ur+/p+U2yLfpMalNea07DoYfZvTD0jEutVzSTYGm6I4v7ow
qPxke2o+AfVWJ+nqr8nZ8e4pYoACcngg/xyk66pNKm4WljX3CM4zYnCFn6/0auzY
rZ10XgwVqJsWuBHns2VsF6DXOkgRRKep9ISY8f4QL53k+Qwf6h9MX2yhm28/wusC
aH7Om0HoTknzwqvJPfV3Of6usRnol1UcM7lGmZKbbQZGGHOAp80YidOC8AzEV35S
oI0eJXxMcVBjkzMOrXB3EnCBui0Cj1hiYMmtZepDgTFuGBmrkmzMsBiw3os/vFwb
FdR6QLVHuLirpyH7R0WaudqwO9YZhHvTeC1ZbIvPYXxP1AhQqwQvudsPr9rsIzj/
q5GOXRzkY0uAJsgThuw6zRGbJipuMzpNlq7u6490RPmrSAxtkNlBjeAvIDgvCRzb
5sNDogHZG52Jous1Dbdl5L+Ga0Cbx0N9uSAn6Zp5DYN8pUSx2hGAGof0vTFwcY8F
QR1WgRe4fFFmYafT+u0sqnqIYr1zbRbWSEXLd0vUOwl/8E74EHjTcZNJ1u/9iliR
AD7P75hx+qTCJJO0XXXdwOlsSrMss4uJ8UiDMDJiNxyan873C5+5Fe4Sx1Oz/c2L
8zJpKYUSayUuE0XSQo80JtWPSWnKJXzjnKGzMvsQf1YsFARwqG7y9xBqbwgI+vr0
M0pvhJgr0b4vwNob2wj+0FLABM8tmE7pm+8czFEm5NxtjLNTyLoj8F2WM8gt2W6+
nyvvCqqpxKt0hzZ2ei+kQMT6tqBwcMgg7dZ81DEm4wxR7vlCD9mXYteFDPJ4WyMi
BIZoUf96rul48l0FsNbT3R/xXtl7uMqY0SDjrhuejMDdl735V57mKLC2PU3fNSdY
+NauORCXnLL8MDpvAjXe/bQrLtZyGMh8dr7w3j5WzAIa3w43cOQ+s88baROnS2s7
xkJ275fOd8hc5pHS/c21UB1jhRJnGmm6Q6DyECamEgmZP7VRQ4Abz4fg3hUAV2Iz
IWtn/bOkx8Q8o+ew+pCBuR+aX8kBdGjUPFlbJGwNYj0ltqlGS4TC9pA7mgFboYkZ
K9pqcozfC1Ctnnu+zK1n1sKeLwKMYRmdc0TxGI+KnY0tqatk+ix1j6k4RNVHt6zX
LuPTo6De+aTm/LldNJMcnKxByhT0mwsZXY2bYEDRO2ZNOKJjB/KHUMsSRuHkxvrN
7Vl3tG9XdOc9hbREfDHJHdY6rTFdnXcDURyVawQcNJ0J0Z21eqIQSGR6yIWywsH4
7n9FrYYCJr/s1PaGJa46BV3LTRgws5aNM08CHpyq0DbNHdFWwSTLw5bWa68ZFW7b
IP8S/AkkeFuMmRqq3oCI1XWgk4DwyrDcfbYEL6PUbjpPsxE41XZ8RiK7+4WzDWa/
tju79MwqNpbHpMGzeAK0ftdxdCwNIb7wAbQ4m1X1+P2iQ7s9oDJAlY+RVMfbFYQ1
iuEAg/goKczKbqP6FIiswIK1L8bnbfPam6lgHmX3ZtAcmBYOlhqK/uuVo0Zul6iZ
EfhGrIkEZR86bGABa7Sl6pFEg4KdNXOAtLxRNhN0CktlqsGs/gGxEhQjUWtI0Nl5
AI1w8atN2HK/NlZDJFUl9kjg/NILJoAsCuk4g4aA52+5shs2Zp/Prbi3sSlRNf/U
pQ1CL5t72g6/zDI1Q+0+RgrZ5LaYD1oGfw99n2jrrZGPQmry3tuWoNIAe0jjmQga
FCmawGi3tebctAROQJY8LkBUrj2bF7t3ZJTtvvpRQSCfbMGDajiyJMKSmcfyC+WP
psbWkBrv/J4Qzk964lNXhTI8qFFl7JqXKAwFjrdeL95dD2ouPjWw5v4znJCOaTyB
Wu+Clsce/bibWGSE4m/O5KRDRcvq6pymrJl6GaJOGuIvN7fC++FV6GKcUyEs9SFu
Z6lxJxWGDnVexHZ4EYazvWoJwEH7qvJgckPUwljAwvAe+UJ2QEX9nZxJ/o8Jk+0M
z1W2wCIYe9K/3WTZMl+yivGweM0NMAh9lXWgLbFhBThPdZhpFD+9FNSQEizmOhac
TU3lq9DJYgdk/sxuHdrB0Mg8O0HO4FR+DOqtom8LQwhHZN7RvvRFbryKT6fo80hc
gUEHlpJuHj7jqbM9vJi7vkev0IlkzZSJoyL+8yGZm29ug5ZYsiv71oaGnCSyv93w
awNVzPx1TmqzfSOEuQYR3pj84W82wgeDK1A55iWyPBKkTA76GNFZAAw8fyE2XnMn
IVYC9mG9mO/lDRHTwo/0aIUpIkghQ4m56n+XQRIXRpA38VhDFdDjIhH8zsYKmwc0
NSwWg8imztSXBRGqzVkoIxZbEm89I2MehPqSehdenxI05+0lnhfmt930R6bxRcSH
9iQ306RBsUOR7ntOD3uT9jo9mDnN9B9xcbnCkTKh/B3lIJ0AHUJCvkJXAPvnoEW7
clXYLvgbEV4XAySkO4zXwcY5cmeh4oVVXS0/66y76CTU2RIjWtZtRvr242WU5JBg
wMlob6PaWgF+5Coxpl2a7DOUOZ/MwQuaV4YqPTyQvdsR8ZvavgdMKUzUweRguGNV
g7U4zDve3r1q9oBQQnaYY9GR90yhR7LAdyQqhEoi+LLH8KGh2b5QvNb36z49Ve+Y
yLEa2km3yj6cky6yG/dZyGkZOFtxWOrvovvTg6H0zS54zaJH+fYyMVrRwbQa5SnL
ed6OpLg9X+1edkVax4xSr0cGK9x+dptqaEBDkVXyXBjr3i/RME2zFJwYvm6051OV
9f8uQSVHxSDDpvNWbuxjgrO67NcQHn2Ga82tMW6tUDj3ex+x7Fg8mMifB2C4yDQ5
6zkvyphc2AUWn+RB0JxW7FjGnYnf6mmkpfASbcpl7f+Xe1Y5JHubVMHuAGZUaX1r
3832TxighKVVJ/GZaplOx+PbtxZeM2UKYL/B7wAFlEXY2jleCmbeJIoEL+TK3mwM
FkGFLDWIdLpVY9qQjsFvgkfcbw4fwwuJvYqGi/j5wzBtXbUH7pJRdhaRTNxLA6UD
APDqE9ejfQl8Q60+BIwPwn5eOl04ReBLAA+d6Sr4pdioPGE4o5pm5MUQSZM/p0I5
iM3YSa8B2sJTR5lsQHWfzXG6JY37wlzSt5oavDOkYZQdAUt8d6puoY92mFlhdAyK
ocCfKyUiomMUIgl80SgsMsp/LWHirODt8wrUTdwAl3Atgs7vPbstPtD8Dosk7Uq/
4fqLlqr4wRntDISUdB5khoFfDSbnaQa3QMg+v1+JENi+byV8IASlS3kuEuqjoXkC
KrjhoUSa4hnHviO1toaL9NgBfJKMdczBA+Bkex0jfevJ9jfkA1pG+MCNFCFVGxVm
PAnXJkF7JU6q9uvbLj9ydZzjIkGAn4CvQ5QhEeJSZR8Mx99XPw68hkJBP6Zqu8MU
EY8ebGroqJgtmGD17B0qXKNv9GlFbbrWIISnyB3xX0Wpt4+qqnUKS2G/g4v77RPb
eolb+VY9UIxfgZQ16vBepOgF2l6PVFspuYYiSCxl4lGQJ6qU6zP58NzOclnMSjtU
+zp/tkZmY/ZubL/LgpKXvhJpP0rn7cOwcYbOsMVGDNnORZ5VTb+Cm4X3TrujHilF
0GEYBtkt+6dSx/C1gwYHTRflmbGzZ8Wt7nPxeG0mnDxNcKam9r5gbaZhK2LirmrV
FLNetfORR4YcaBdc8a3qnP9XUXadJe3JF9fwZmmI0pJQTVxCaXo1MHDq23QwV+Fb
9aGNZL4oxPPcwazFJd2m+vabzOR8XSGb2LJb5++2sBjtoJUqj/m9xz95gPZ2vrl4
Dt+dynGNCXkV7VFOyusCJzYJ8gPym4icSU7EFhDnBmOwBwswL6DjaAzqfZaM0CF3
zw5j05pbiLEgGJnY/wkDzNK4H+p9rSyOyBB3UZ1q490UCzkwphcSy8NFRB9IYn+4
yejtrZb92LCbSa6Fe45NVpDbwMN3GtvdhMfnuQL5bUw1Y+SS1yuhWuwJonVcnpP/
LME20nfLrxAhgdYvN1pFy3SfDt5BVTQTQ0yPXc4fydvA9gRSwG6yPBu5j8xOnyKD
nS1rFXPVc32grRSJZIN1XER1DEcE8O6+39xtWM2DlBprPVubOBfovGsuujUASENw
DzmWC5Ae0MLNY1qWXWPn6zRC2zdg7JaouZrvKsIid6qIH1F1QYEafB4Bhe6mt9pF
OSpqqIwPbrXA+x03OHamlimSL1Ch8A/FhEW8s+zrksnS+fw/IrXfN5F2JTBcdXzj
AnNAnlxwGwoVwm1IQXHAhtTfQQqQwuP21OFWbxJc3kQdWsPG5gMy7EY5TmWTVRVH
Pi+KZl9mmxg0Ocnb3zaMyNGmijRXl1F0EINVaBDUaccISWgMHqEXVlZLKDjEpXRV
bSL5gsCM2eXvPcVB6YO5SAEkYVbeGpaqEwzIYtNK5bQ3Z2wVOHw/rq5Ah6hPdIcG
YGEOHr7ySrFbgWVhfizpSUeel3vE1kElguL37Ydt5c1uTFm70KqCuzuw33NqEFzt
mSVDg6vylUfZGPxAIfFeSkmQhYLHM6/ymZz32OMdStuReW972iF6Xd/OGH3CUgW3
aBTXc2UHlrgab2g6tKRklnjTieQrTWcak4WHERQsKuOZ/ndzs0PfO9wJmJ8L/QzC
djYzRZtyOGXaDaBCyiN1Mrez5QZ3mrWpI5ZjiHbuVGbYNcRInbm3uGXMD8ApFmw5
8A7dyxZOJAfHgeRtWMJH0vAMCRaok+DREs2R5Cp4BPKgkjT5Er5kJ4FCUfQCXrn9
gZxB96wjh7jjsBmyCFvU/oJ6gvo9R+8HvNpZlekUWyTjKA00hs5B1mDJuTz398sx
alrobjUqj+pJ8+8w77oT9PSdGdqtHQ//cfqohMDQihiJqnAgxt1w4uh591aaa5S5
gJ+D7dmbltnZMqKfZF+lp7RjS/fz2kvCVUADpov6srYeLktDoRhiTK7kwfeosm7e
dxVkEWuavNUbbeJIr4el51OmdwxEdsEYZbYxLRSzyaSyRuk2lyPojWM3GBvB9wu8
9+w5zJTq8lkkdH3ugUs6t+oOMqoZo4fV55Df5QXyJ/KSSLji1kcf3rPMCNuTL+qL
vqqI/cwQGl4OfLEO57MAZ2l3mjimml6aYe66+zunMRrVG0BvX6MkGTHByyi6l//1
rbnSDMo1jGKYX2P4XSexZ/CmvhOdh0D70eFbng3+QSsKE+OjGUkNjVB7fMpkkahb
rm+cLMJO+4EiBiX9mFKDtyCIRhcPIGAEpkGQJtzNNVxwxtqQBDQCDjuspq9aoRms
qMt5qqbUPfoDy17BP8jvO7kS7Wm6bCUxtHJap4x0US48O/fSyyIAO3yXumcc+fd9
DQ5RmAEW7MmP89g57Bs4t1cHm34dL21rBt2yD1urwFHc7tf8wn0OLD/kFjrMG99X
mlI+tDiVMxkYvdK5mK9MKbujVfpA1kz1Y7VjA810EgT5zVyiBhcp8utO81bTRj8N
R61tZgVeRiEf1gRr+PBUCgmmQ7XIdRH5Yz5htOBDCartdF3L5/vDtPFQ67242fAt
UtEZS7l/d9DJrtuzer+fMwZhJH6Le/qBoQrsvbTGY2y+XeXMH44Cnn5OIxhx84Mh
JA7lNI1NAF30LKZ2Etkz6t0Dyc+mrbZxWqHBEEnFJEob1wLa4u5LD2uz1Od5El+g
Onp+Bf9ttx2jgmAhmHzF82QTW7VOH4v7N1wPvM1ZbfzKxzMCsZTAb0Wx1ZvC3IUP
TQ2xTcahb8NCsTlY1QkLvF3tD4OoVDUlvyBBLFAJC1zS7lLFLnZLyRucdK170zsr
pydC2OCuDHu4Q0TH14ndeUkvt3Z+Y5qOJaMOwC9B0R0ZS1Ku/2JgSUgBqDC/F9Ye
0aQfxhDL+5U5O8kDwevEi5G0maHwW0U54/Fz5ifR9raoHfF9HdJkP1sq6xwtmXAf
fTDsuvGwjA/aVqHrNnmeNaF4PSrfY3lSzfUdaN5rGYAxQ0tR3N7mQIeIqSzF3JqO
lCqLMr8/vwaCicEm1Qqn31ltoItQo22iomcKHkREh6YSRHcb4hwMEZ9UkX1jJbfA
7fyisaDbH8BNP35cyLl3YNPNLz/UiUbuHacnj7bHITvaTZ3fibMo20inPpAhvIy8
S7ROD/G/dmOQ0TwWJ0XBz9ZMdYuHIcV4WSL8X77soTd6bU01FwGfPqmuoKRfUZDa
CNPlRcxUQ1QoAWFXliozCLjWb0VHYb+O/4CJGUF6hAWL21vIFdZW5rLT8tKkkTXD
tPr2KIT9cZYV0zhrPjkQlLbomXwijEKD+lL3nhMijwnec2zb/we9Dm39IRUCa2pW
qjLI98g7NauACsGW4igW86EEaIa8wQ9hmWSvFA13ivovDDUujVwvKr5MvY+ItRoo
jc1emTfWiLx73mljtzvV5zscWVBEyDq/XZDMsgY01Sn8q/zQ86J1uYFzNmAonPYX
jiEQmCtLS1HGaNzVP3JniyvlZSXNS2MY9RSPfEgGc/cnuY30KX2lBztSl3YYrRPi
oEGyXWKLLsFy1x8pHoOiLNoWqtq3f38LiVE6IYUqGlJ1gaduOw6WM6exr32SdQET
esW2lOFrU9gXKq/MhTy2mlps2pUOrrspmqmcVgjVLhfnOKTD23Bt+3RQqDXPCaeI
RenW/vn7FTXlGNtcZyIb2VHCLnmfx1RqOOT207LMroNK5elH5RFM6zq1dNdN3wLz
6c4CFlDyBjwiANIPGIwLopcKODNiLSkkK7d44L7HKrI9SLWT7eAnEabMJsRZzmtk
Pm86DHWlUx3+ullUxHW/lAFeaUhWmV/zGcrOgsvXWxfGlk/kQcpOzchsTJM2VnOR
yEv0LNq5awZ3LyUawVRyBCcQ0JqBiXNnUcQU9xLIOR4l4plz+trt+pEF7hq4W9kd
DTHwcbyyuYXexsY7f9CvAi3G+1UgVXQ5qmgCUwa840LAfudSh2TKSwa7P4fHJy9t
p9xSU5WelTvASPeYwDPv3V/147eheQi9xK7NHy1F6n28Kdl1BdCpiV12Ndg+B5Ge
sBgh0t/6dU8A+thXWfGBB0j0ue3NbbbOYvr78MHYJiOsVThOADKuLxpLv+IA333y
yO5COLGRGV+bq15K62T2IxnfBCKzJzgi8JfQnQDy4AMW4DORuZZE8FCzcus8Wnc5
z/P6kL+49YI1mC/TFHxJMMLj4gnYPAOJBLRqOQK53+IA5GVlXC2PJZzg4MHhy9F4
0ChPm/dyvO6yl/kbormgKBJbDKEqjYlp01ruBd1HHBzxvi3cG9GqvDCyOypf9lp1
BR7yabWDfYNh8dzj6Cve4oTAMQ0zqUm2SVugefdOmyc4K+ow9EyejMMfoYKrjRbZ
uVlmUSg36FsBZqrqNdb4xJPgLkNk2YLVd0InkJOE0t28t2Pbe6j6H7X5MofO3RTo
Udv3bgYRrRV1kq9UR4CoiFN49jdB6yOY3GyUKxDi6ZujnmO6efWwDsIEeyYDKflk
GQ8WZW39JXCFXRoN6Y3+ecakorb34NEmVyJi18kex4/fr+qn3dJ0yZlBXPnwP9L+
j4GCJqLuof5MklyvASoXsHbyxOnPNrjtA5/G664kfJRlGw09pizbVaAVvSNyFV6c
/9sdQFKnTfB5xQ9cdejS/weL4p3dM/w6Ar/H/JYiIBk6H5mtB/6q//r0wNomosm6
7bFct+GhTF8PdaFD+3GsPubc/rdlUlmSdVmfCjidfBdPyNvpHirBjWPeA7IE5vjz
kBPNv6/1qH1hSS98dW06WcBSdNcxqRM3zKU9ykRREgEaIhehBGPRA3rE8+W8vs8/
KBB51wWU3P8kDUgrjFThdeAsvdtXNo7mpFYBuFrz040G6GkLJNF6eXB6pQSgFEqv
jIQZo/hJ5gpqd+ahUlsTifOR/p7eyBmWE3uCk3kzbsE5vjf8fELiOBAqtFXlSQ87
0+hDJfmUYzDVuiAApFEY0GUvkElsf3WUV17ZP3VCy/RpjTFqXLg0wNBWFMzrwlxx
Miru9htJmWGAOtrT5ThVc3ObEZys69NUqK7mwUhsXAq5QiZ5bZ8BOBUy4nzJDSGs
S26Luk3pEHRWyTnD21idQyguWGGcAA8WIst2LDvIPdExSBRbMc/ZK6jBijjXjBOZ
Epr5KiK+VYbRAN/dbY8PqlZGhWQDDppFpSq9gOmqc4Sz9TJGbQozd1gwVgbv8Zn3
BNJov5Y9gQd1ExJU9LBErdiWcfnr3tN9SOJi3eVuloogIVgaVdaRSoWp+7Wo6/Lk
Co1eOsRpG5jATuJ/em6/zBVd5GiMs9CZK1igvDZe0K/RYowz+H1HascB6Kg91a0r
hPLs1sDm4kBcy3HKSm/LaXFmOh/4e5rm4gdZEY0Rk6U64LabKRIkAExKw6ZoqZFZ
hInPrct4hVT2BoOpMmLR2LbjVU9z4AmVBiDTT3/UZl3GD3iLQ8w6A/+VdiuDZYkE
4b+Sd3KfxBtwc9wj8/+OOpDMCH9N4RJCVMMNVHnAJYGx032uIv2nJhtRYLnuzA6l
JmK8ROWHMVZJ9n3jjPNJMCVFNSbr87cAGixagksEgOW9DqyMqOQutRv8mFpqofWz
PefBbYVzeURLrkjlyUTlvGTJ/sqrkVXXOXgxww1CVikjz1INzS8yxj92Y8122H4J
xYXKDEaBPRX/lB4yZupqLTCiCaXreqAH3q2CimF15RTiWJryY6bmh7UFVydD+4FX
11+Kc0MjbGVF6rSlODcrAeR6sjqsf3Mzrkq5QGArDATUsLE2AM5GIIPKEyq2J9C5
i4lfLT5z/y9GA/C0frt8XKla+XPKNNDR1cg+W5p0RoMb9zRxgrlEIEPMhuTbLvQd
oDNU7FFqcwPNp8yK1oOnhG8WGVL0/nYt53guVQ9Y9tBKZWo9FalnYtMtdVneu/0W
d77lUjNL8S2d6D8FjBotzDQiHvU8MQSH2waii0gKwSz6MfdLADs6MRQbDRsW84zW
YJ4xS2EiybiZTtKwXLGoesT0ljkYvVIo2+JIdKJKWpif939kf7N0sdeN8K0ijoKV
VV/YfHJ+/z8ZPU7liqG/PESAY891YMuNtePzfpNhOk0tdQ4lU51mxjklwqZAHXYy
HPA2QN+TeJl11ZDO/yp8h51YLRcOyaV/hrwg4yvhG0SLHFXEo0r15auersW3UrNv
jnaR8nlH9Pr3O8d8vyuwm1A9ZXSdgdpzC8dJ4gFEHFfGGHFPdFe/hFwTi5Y+dI+D
+cLxBFiiVYhHLGX9+diG9trqDtESC8Biv99bbcoGtqmTWvsZNK4jtWwpahdpJIzA
1VjzQvBoOqkWdW6mqsk1yv793VeXT70qusmU2GTXljvRnfDXcua0JMUKiwEfll5f
Sjw5Nl08XvxsoSbzAPFUR5gZ/xZs92tv65RVAUVReQdJevZxkVZ5+MQaItPh1X8O
iCn6zsO+zlCUEx1ATgznyHgVB8a0lyvk64L08e77YVmpYpWN2gQ5SdzYi8mUkBae
TWofCUGIoPC07WAOWS41FowXDElzFBjZk+iy8i/7C9dsf136yQQaBOD5Zxkwf2fL
3IysdDQuHfXwC6E6zxjUiMNXnBLbXZJ/fps84EFTNkQDd7G/pA0LFRVzAIPDjJdz
N8Pat5hesrHA55Y/7rxvhIMDvqy5p7ruVWbg9gYSEh3E9dpNK4c8+fxoX8jPfr9g
v+3+wOc0w0l4BQZwpUe7nd/53P16UiulBhBr8+yfaX7sAKRilGUdnfI8GlpGOZLy
LfWiN6+AwWOKmLHCSVf1NsPzp7n2G2dMJEMDE8hOdt6IMvx3oLuX924D8z3mWkFU
XdGRPCResb9MND9lkMbdhL1oVYaGF30mOAXosD3PZKdq3QXUeLYrCcAtQI8T8vGz
5TN9Pp3bBSMk4TlG9OiI/QhzCmDb7+pOkJR6T21D4fJ+SMBDgX4ezxBHxoEniJWP
y1JpuylISOpGSIZf++sgQEZG7Cewdl7i/rPt1rWsdNepWn+VUlB0GPSbtTt8iOAH
W6L6e3Y+T+S0kRhUx0IWwBEjmWDT5Mde8uEyK+MylTosN055dv9d3QQcwM005vYw
ux+Q+N5y0m+eavwJ7jB9/lFf6hYvxXOZ1nBIkcNagZbAo8KZ+iV6tmWKUA85ismZ
Gnq+gaA/SSMCAr2PUFE4PbYfk1w2PUTmDqoAvm+OlhTEAvULxE562484VN0Bs42p
czG8XKKJjthgn5Dt5h5vJr/gqF+i4GVdC0IfE19zGYt1Ixejf9uUVYyxrz2X6wk0
1VMpysl2Ru3jHlsfoHzrA/uF0ULBtTAOS7ljjaB2bK0TZK2HGeVhREXNBlWCjt/f
HjZwBy8SE8Ee5PI1Vugxnsbcr+fGZDOgAAjq9DYK7YdGmDQPe2au8XbJL3clxqJW
KzOx0CMmhiA3nr1bGLOMPbPL58xTFct0Ibb45VbUZdBVop3WP6gTPgAyIXsldRYc
WtYyRFGG87yU0us2JoINwNzP23RACt86A9CRU477KVP+6QST9yyIDgc797Bg4eoc
NCKGvrQ9lwXaL5VydBCvFIqqEW0UQsHmxhirCQKccQqGqt68xpJDNBtXTMJxz4jD
UgwlCL5jkrlVzx/apR9wQDTsKwgzbDl8+ao7oWWXXbX5luP/riMXku2uBvpUPxz+
uAGr9lwhKhM2czIDunEtO+rYdRkSVjVsYsvFBzCgMdpn3JLMUpFFEblkugS/2D3o
70a1sNL8aUElJ6BK7/KgR5LHEyq2Qi9DO9kjMkz6kmACWlUV8JVUr6BC2Pza24Tb
bUjBWqcAU7TxtVth6gL2h3hcBkc7zVTYdyweUlyDfeUquyn19Sz9aVpx50f1rKKc
aoEP+FKTa0sIotZ5hRUuy/1MQqLJM3d+PYvSNJNQz5s8rFyC3mch0IEF3SHA7cSp
mRON2GnZtxBMSUfKE1LC72B+sZ7TuN3X38rmndwj9EwOUDA67ezzXdnJFm+bZW/W
41gBolTmo/un7V6nyDXCOeT3F5xZ5/OZCep0efVd0FqWy0Rk0wvnB18bLrdMUJ1e
45c08/Nm+LuO/I8nOUPe+vrYNbsHkNS1pLjFIj5FSflIFCbdhBXYhlOim7YYsLCh
QFn7Kg3SRvIhJ4PsCGlndxRQxNmMCmusxDPCSYhUgrYWX8eJf7ipe3cXMlAdgRV5
tE1ZL6LHhI56ih+QobJQllQ6loG1SlphEvovcsOl2igVFIc499kenSDyvPmBKtK3
mggcPheUO8ejnS+xIf6zfWKUJofxeDKZGAW9X177tO80dX9xm66v5awu0slGqbzy
i7z1tdzpXeVyDpzXvN1QAQRLj7BGES7jafNzKsr+SKP+5CuuWncsuITcd3ZeTxdd
iYNf24J0JpAzL9p8uRoz4tzA1LjRsJY6vNEv+dn4RDWOwthoLxsyFOoNddjnkoxg
Vvl93UwE6isg5hoajAPJze6P44Q19Vi4AsnEbnAcqnacNkYtfo+gWYxuaemDG+Mb
kp0hU+EYn5nNrKyJpxiUqWwRfMwOgRTPpOXI1xyd4hdZnT/o7L1Oy8InjR8wza2X
EUwk4kXCVtxvP8vy1PZsZZ6qFiqAo5h8VeZpv4CgpnnJdKZ8CTc4CQxCvvrEqNFE
m4h1GRiqu9Fqsl26O7UfYRw7S/q/DCr6NfuryanBCB/senGMP4QeM23ZNGu9CvZh
biGN3StpqVLu1Z/On1s3FBljbN2P7LlsBJddtg6k6ahnlaON/9/x7OaE3WaDc3T4
F6qxFv6YVPuVsdIiw2WO7ssIFozSscP143fWyn3SRwEOIURXOGBCSqx3Jx5Tnv/x
z2yEnlXJN0MY9ixrayyb2hog2uddNe7NogAKlLA0nYCsij3ferC/57sourRpZDXO
9VN1GDkwUph5+UKoUk7/erhmkWpW9hbRsGZepoao3CGn36PuWF2rAL3lTRD7dbV0
BZmiVL2l2vlogZdue5SCnJWiLdD2LWC4tE1IDzsOabAks3P2hh0l6a72veRH6huP
Y64rpN+b7Ex8rrxjpFXF3MUMgDmZ7BQYajVBoiR3A3EZDmlmM87l1mOo82lnyS6x
hrix503RYffgVfMezptNPvTnPJmKYLCdYe0cY9GLwceQiJYeHGOuTSbnwF07OYgd
9qASs/KdeZB8qQ55rVIpdk9sWPybUhCzPkIe8zxlBheuBWVW+KiFdB9YiI5wddA0
KDeRkB2oduBTy0w79cwFH3b9OIecDB0zSiracX3DQJbbk1mMFNNlc+2KSfDTpogy
SApVVImIp14wka51+FeNVgdJe9oFBVv2u7ldTYmPzY/DEIdvGtkIR1XIQtSHOJFA
5ygMK5md2aPebGivByZ/P+ZB+S2ZeohV5s1mI2MsyudlTXJTg1o4GWYLPBKvWqkQ
n6OTW16nP+fVLxIubYCTNF6F51qwRJJRytaxB20HOtXVdpOlGRHmwOp/ab+ykjF3
rI4VumrqPqBzgcaNOc1MbnfFx4Fw8f3m1UtyI9xDEjSnYxukdDaUklO7wDOnTYwQ
3kfTiK0Rd0V2reYUf1bXTFSa/m7PgUzQbUMQCfbJhtu7BixJYs1re2yR/i0RpCi5
Jv5RySsah4Ehud2BiLs+eBTI3otjvcVdkk/8BcWf4awJmmiIsbUGUvyQERZGMPIL
zuFITPxbY4o13YENZpzULsqKSVehdKq45htdFwqdAvTboRWg2VYU3AlPAmTKb2OO
HyX6ZwPmNzJTy9MlK6P3YjCr6WfI0BngYDI+M5hxqyBJ/kwE2dMUqGZR/6UUeTao
gaQM+DfmjDV2XpSUuaiMI4bM+B/E51cCg96RRwMxO9SkYsLEtUFEZ9IiW7XEBEaZ
FoMtUKg+7vmux6C1sLQ0FCBrGqRFlSxSUE6fP50vc1+T44VDHJEYKUuqK9JQb6hC
rurpSieLy0iu0QL4h6vd0ul2hH40got1imOKtDFRKlN47m1KGWUaXnA6xZt4SSrZ
cs6ROgrjMKPsNwA+mNWQZCmWVJJK73FMcaG7NNhiz2mfeNh5kZLj5LGs9428YAim
GDFM+3/dXHjLp2oSUFmTUpNRNzu4QWCLKnOlbz6qlJaLNmB35o83H1nhqGanCAO3
tUfGfIeIjJ087pEVTroDP27TiC/pSoXJm1ht7w+NOXqpiBNxl28E8PmO2gUa0ViQ
MnA/PzazJp/R1/kesDoKagfg2u23iSk9EmSpVBs8N93epQk5XaDQUMJe/G1fWliT
o8aPP6jQJwMtt3ItJUFygkSQnQLIHAG+aZDXL3W1f+4U0ecgonW6/AwMr4C7SKR+
ndR/7x0IM7Z7ZhD4Anm6kQj6Z+/uiUQcHr4cpgaMvUhMDcOfskSqm5Cgj0p3snw/
CUMgewCd8Ve714bFyXPXM5gaWnXTHBVLXlJE/+vSbvfnODwad6rrZ2v2RVERjOTA
xJ/VC5JAdAxZ8pqKuxkwQbZiVOODAWp9KoiDbgLlXkI5yNhmepNct+vCrUHk2VS5
x9JyuRSsFjpiGORsTmawr/eLmr0tU+LDMk17TohN6ZQRj87k0RN4LwUZLHnGQT7t
lgGTykA5YlCfQC89jLcrnyrIcn37FyzY8rOZCLCzhi60l/NBpjRph9JUONHGneyu
2B9Eh2Nt4JhHr/3ZIU13ulJlHfqip5Vqs+7NGfqxU+Ilw78Sw+HzRCUtrvYU/mo/
zPad8adWyCV5cWlG7GLTwoznsd2caa3YpQosNOVo1uShMjnhkgOOOTgBCzAyJzqE
xLKlm3ciQf3mSO9TKvpybhM+hSctDTMX7krg9T/p6k4E1/uaARNCQGSzZjsMEluR
4z/3izr0XXWD83Vo1jJtnduXXiAcQbmDXQpKi1fGRZ+Y11tx6q7zSsxpSVw2JtG0
bztbsoipNBBEu/D43T6f1knwWJoi7+TwZ4bdjT++vQc66PidutsSgFWUrMB4C524
a9VcO3u12h3NDl3MEFiScGBmFywPFvc7aKQfl+VLib438QX1J533Oy3L2GuuXJYs
+gAarLqtLYDponjnckrYoDK8Dj0s5LfsF1Rssy5uGiIvXaSHXaNot5f1leIfBxki
HPUw6iklxz13bFEhJ4VZSjcAfgpDcNkDhaPvpEAJRKxCuk7SdmbVj9YMUGSZrcmv
0E3IqUfM6+pRQEdb2xXRrUD9EuXgx1xjbAsYFC224i6/UsXPhus+lk3F7icXscOx
LOlojkj0PfSsNZ2qMaKvMgio6iYR5JcfZNH0FLGNU9VjlM/X9r1chxhal6SHNF2F
sHXI8+s3w1bBHI/mcY607EGcZ0PaASk1djwrxIOABPKavKMxPEd+67GluKIz0MeO
lF8wi4KdpFWbVz01lvrc1k9fN64+ygU/QsWV1E/4AoFIgpO7Y+j8Nf+X41In63fw
EyHVL0YEM6xwTO17JXg3fuXD9xZMGI3hqlSHTeDaW37oMSAzh+LPB6lJoNhbhBT9
Hq1WEvLRsidcFcst22pBJ6/jG9PaSZh+iO2ebeRn29obljrBeTuFjU+7TNZ9KOtY
kfJXzErWJr+iFIPZLPpGHA250o552sQP5Smp1TkkVRORf7Xgl3A4ZlhP6oJJqOnB
+fKqNg1ohunLqFdD7wKjFBbFB2GXLnkpeO14o7CeQ7nIcrY7W6GNewzl2IUIWmrV
JbAWLC+UUu8RQJiwCjs/15iOWI+kzaudYLNKBOX9MliQDBLILdiuDSJTou1G5PzN
Pud0zJyzXTltlbwLlHq9TFf0demQs+ujjhrYjLUwS7bZe55tQmQokc94zFpjxRu7
cjZWmKMHb0HvtTW89cYRojaIXaAFJkdsTKGB8sAtkImf6cUPu0AxVN8e3yegRqLr
eUOOJhiKbOrrSIuwixLcCs9Ri+6b95Or+G9w2L6abMKTgw6xS1c9gxmkB+O/wrJf
LyjnCNAHwHCJNp9SGTwRir2nJ5x60NJbekju2EoycCNIUEbKmxdZ/pWniBIkYuk5
nlAqbOAH8txveFdvDncH+rxevglXaw/ZyefNuCtMo7BhD60Oj1fCSzyfJ457MvgY
w57F789oR4xu2d1alBhFJbtcBu1ucRNYe6ns1EVxZ5WEVFiuVV/XO2zjOMiwVYKJ
C6BA4wEfoiJTV6iX8mleFxPczVXkSfRoot1l5PMx3Ouc2ZUca3RJ+Dt29rPCc6N9
AppjHTvEeMSFno6F/FDBEYCI/s1oODLusMIJd/NDxIw5bxBo3O9BLJh36BmfKAbt
R6eMWf1S1lz1shBUkHbq53fBcTtA7a9n12a/ZrSNVubNzG4i5a7SOB1/OTZKtViQ
/nKKKu4rDDr8NNoMa+lq/zgM1cVeA0j779g2x9tR1gt9ZQngAscZ616kAsAe3rB+
DHIcSXaopXwKsf4DsqRbZ6OlFL1yCEDIvb4pWVDdaxdvcharpe/1kCjZA8Lp3SHi
/0LU21mA9ZyPzvVtxPxCxtjYCaYIcW2dldEjQtUnSFai6SV4RlLb367qo2pR5vWf
AHsLYmdbokLc1XusMna0g8jl5GlESbFQwqqqA/Ylms2bGO6W454N9VLNNiQugTzK
hfGJZ5WU+7FWDPCtIDMuog6Y3waAJ+ne4+M+9UP0XOcXp0uTe+z7/b6+80S2Lm66
nld1Xo2lv9NXRq6GXKoopX3DQjfoZdf3qDSDxIe4KrbvwWnFMc0RlNQXXy7/gE8m
TphBE2jgPHoFEg71R8jZopehbkFIAQX/32QLlWKWHEuXGdxLVaXXgNZWyBOiaFoN
LkSiW3dXLSCwhmIOYKrwyfN0s7RxIdCrvEorS/q1JfAAX7Ap8so/JkqIyTshOkqG
7q6aDhNz7FHhvd+QpdPzVP+d0MY5bt1CRTnVj2nlbPsVs4RRTUKfs6m2Ooz827EC
0q2jNvWZ1gUiOnFZvDOe90nOvfP6uNjrjLO4BggdmeuUY2UwaqsTYqZcUB7EXIkQ
hfWYkqRuD4UpnUvCI8GshGS2NRWFQdm2Tk6CDuueDipO46NvSV8zE5gTC/IBk2eA
SjqoKcZDlfrc7rQqXt2M1XOfcPfIIWiw1SPZonDTdtRjQf8ys5q0EhKLiyXeT26i
UUg0c+ZuWRwDJV02r1eVBlzJhjoMpIiBoFqhwlXD8Y359kCMcjn72z+j0/ULUBSe
u3GJxVPh9c5v3H+QACQJIplMjbY1oSbNCalGY6/VUm6JjpDn2KF09Rh7ybHAej6c
TPStUXt3mkqVaRCyniRarHhPCRxQhh3B2bLS2GhMvXUen8P1p25ZbQTzkEu99ip2
xaxPSA83/bOYXBfAdvXjC8zHm3trSjG5AVmsak1zeJcFA6TlGK/d/N4FvLhpgxzu
8RLWL8bRt1Zm0mWteYAgS2BZaRRrX2fvpZw6Y2PgMFlGhCb9vloL1fkx2OgvM+do
UReS7G/cwYs976azz4DIeDmIDCLFbKCkalEYo09F3jbr7flVHRaQtcDTlnxrl+rL
NKsWG72U6WTnud9bapc6TZpK3hDZD1q7+8nzFrjZp9x170Rj6EqGjDN5ZrvuScma
w+wR12OiygxbA3ocYmm9rNIfqTsWQhIY1ZVfUqrkOeS16CD/Q/9l9QSzXvHcDB3A
E8wissxQt0Ae+bRZ0jSzrERDM/UexBceIz6MQQomoKySFRIzHTVTMM1iRgPhzWKx
D+ZTK+FJ/8d5uwAVqxCKfFTExak8rVvSWa8/VbxEISWt9JUFOaKQ7NAx8fuX7GhA
GP5o+7YcHVXcixhr1T5izXOOaES/41iHeK11pFWis6pxso/8CdxTbMasmeZDsJl4
Xu6/FHh7eFPGyg8MXQbua28sOFMXuoBZH2PZ6rRuAcI5R+ZExc6Oj7cYu58Y5r+y
PS6QaaGPFWh3WTsjsKgtAw9RLocXnAOnOJK/zZGzcFs1oZ49i/GMJJELOBhyImQa
ydf6S56qCreYVUMAaEMfXM7F/hPVxXB0+GVrsA86gp/BpOFVnHbPGgzE0f1uTCjZ
vxUEulPKQvH2r0NjuxmHGVOdue3vBIu1tzPnMpIWaX05J3fcT2eA1cmOvIkzKxjT
9S+yYaEh8xPhHq1imhKn27T4+wXCbb/N4NTUv/z2fRirnf+bLd6Fma2AnrFumyqM
nLsiix7VEMftYqNhL5UPo4io0Yl/L87b6f3MGnmRlP1DSzivshgVDqV2KVgrvsKq
BecWATLnTo3c/61eeUxrJ0Ai1QXAR71nEcoGxy6cFMIlEmCDOMZBQOKsj8bZzQMZ
iOhV6ToWnrhz4e+peIfS8V8S7zCi80mmP8jiP3dHnx38UPIWYLUHykxqnRh41eXL
Zx/NO3fxpuRX0jM6GAdkcOzG4QKmGCpVZ12oAgd6MXVggcXlSlAa5t8vdJ3hnWvW
Xod7JAJIPUXnGFfaIUgERFy6OkoJvogcqogHj75Cdi1nzhUy0xyE1wVbhBJSqe2s
fmBmiyxF/xLTN1yRHLAnnX45JiaY2dE6zTLi9HoEbFO8vvZcAWitaeTsNh5TEwi4
0FI/v4GEsI8GbnhcwBxc09+Nrcp9kk4RrjKBP0g33lUwkPjgKO1HTybESWbXDJ3Q
3xFtxM3oXeW55/cbd2tFvKijHXHFnvz/7ic6H7zbLwlVzHxwEwdJvkn4/FQPrr5d
tlJQcpmJMTp+QWdZLnWAFprmzyEhhfjtkxEOhjYKb20k2PSPTUvGfwV1LjsH7dkE
rJbxYlss7MrKP20R9Y+nYHBM8UovXOUMdb75wHwO29o9+IraajTmZ3GxigTZv1Ko
CxzHxhlOURJ2sl/ViLYDaj5efbr0Zw3cRbA2YkusIC2aR9DZA+kaWx5qb7KkTalx
vAWFHfQ9ZT+CJjB0cjRtYRHIsD5fIq/AOA0A35/9FZx7pooK9RnM6Z1V/3RtzVCP
rJyjBlh1Ab5fzCmtRVRrivRXlnxdHEJXL4vllhKWqmFb0GqTgj68F9U5ANl4RLy+
o/ZnKoN8ApI2031lqvjLcV06cGN3Kuek4M69D5t7okjR4L/DoTvw9iBXJEoLDeqC
K4G9izd1lB5D9VX5svxJwYjZYFw0bv8tMw4PXbtZ+3VrsjXty+Gm/qdTQXnw8iZe
H2nh1HDtfhEcnnPtfcqRa+xTi5wIPOGegi10PMiOl9tpzTqEBa0Ka0wR8slghiPZ
qYWvKyXvIR7B/WOokP+PFoFwIfoyywkEYFfVAEm3hz69c6t7JrL0K07HXYlhjcqj
MljKYaAxFkdNudy4Sv1g8nCEPiFG+77kMY/ndPqn/hXN4luK279dD6WkH02GkmIO
rpQzeIPlDEjpLBFjJzHx5Iev8LN4DNHH+Wn34O3/liXP4/xvHbRo31lL0P9/WGSR
KlsPQBw85+uAiZ7MGGTsZAale7SdiWvhI6eR5n+hNdTSwq8uyVZOF/gpARDmBWId
Ip2lexLUIDrhpmZPcAg5qdrDx5mM2VFoRc8VtTAsp28p3CPZEiKUdcAL6uMa96VN
y3LLrBCi1+a1sR02yadeJQQomdq4414hNcb7T/3UZ4SmHwMS7rqg9UaOR88QmZy8
1lA+226JO5q+IDdH6VIZoh5xb3P4DDAXEz8ixM6bfrlEDcQC/wTLGxvCxcjHKN0k
hAKf+Ezo9pIUYsBdUWYX6sYJ8GuHAmFdXuw9w8v3RL6BWFUF6GCES4cYZ8G83DuA
/dVtpJKAvBMaBndVC3pm3X+OX6jb86cXvNZujs44fPVMJExoZr9V6d88xLgQcSCu
ZTaSlx+6161SYgY3PN+lGPDi8JRxn7Xa8z7JvnVX0AzfDkdr+sNBVPLt4zwRF1uh
6oIupErhOFcfcu1wuDGkQHt7XOjJVQtNIPhaBzil19KuTjm4CwvTYbJFW+Y+hA0J
xcgp+mc9Kfsp7Eq+8rX1z8CEunvW3J+YeEwL6G4WvIxlGzgenBr/loNB+SLgPSnr
V4VHsTanvrPhQXwCi6eGYUhJ1eHGjU+XIQrdhowDjNIFaQJ7WRp2piS1UjyJtyQF
RAA6Z+aCoSZqDaO9N5wtb8SZlZtAoW8g3GbyWXpcGaAMdDVsrX3JszKDF49OU7/A
WM59IW7vZl8LarEGMLrVzda/Ap3ZxxWRjj3nyFUahv0LS2KHiYhTaH8UM/JnKi5h
broSEf5EaPFS/fKrUE1MqFYiWXUGaiDnTQzHcQZTZF24szdia5WUIXmwOUJCCKs4
FrQ/1tgJ6dm8dHp49wVEw12BvKnp0bZidRaEoLmI2rZc7MXbKBS/hxJaQE/wDo60
U7LtHtfv/sUGPRMdeIeExicSQ4LlnqVHg9MzVCekBd6H/N4vPcF1MKUC6Ah6skxY
uEMf9wA4AUG0ZNrXr+AhrW3AgYfqhI+eJxHLbU7C9GAlnyOjKYDq8BgH/Km5s7vZ
DybWC7ZbjDluYWh06v4ryYmoLOQYT//oK1LeH6JZsFPLNX4v6DwvfUB6Itq4GDjv
xI9XW7MM+tw7ADseBwUyT4ungtxE7yMSmL6V1TK4elhzdLaj9D7h04sznOlsPnlf
wpv5FY8xTrIE/utujlx/Jh3QoHAQ8+uuviS3DaQXc8Nx7+EsH9ol+bsxdbYWf9uS
O+pxt3XPuRF32Vqh757Eq/CZ5fu28PG5tmWvT82ivSPLogpqJq6QylPxRyVYetdN
KO0socwbK7xzbviHLXgVcNf7XMXmr2ywN1HNt3Co6MNzsc1RwHbTP5ad/GoIvR1i
htdVJKfXpAoNHO6VrzTti2kWXD/6F8JsLoiYIZCUlMF4TDMpA1eZS5usnQhxyRuK
OLWuexXNB9wKGufHwVdyB07cCo0VM/nIWH215j3I6+gPkDISkrcSsvu8HNaCYZJ+
fKwZhy/4mbtme8pbdp6xO2YyZXmyw8XGtEdSJOq+tOLFkonO9a3HwRE2pdgnv5a7
UZ5/RfNYC4LJIRtrDGRAgtxbK7x2EbHXgLrGQiGlfpwzBuvTlC3xgHt0yRC9YRVS
EOZRMG15GV27A3KOsRV45Z2VZm0V6rlEH7rrutrGeHrhX/B9S4grzjyoaB5zlBdk
YkRREFVJ78x99c4ToDmmJJpPz/BpyIfEQDIXnItn4a53JqQPTJrLrMQR8PteIYwe
6qdWuLTf/DO/JfacKrmNwwsU8EAqRm0teeNFWeotUwyQ9NgKiLKfnlyAKdZMugEU
MZmdQr1OaCIffBJCb4uA/Z4lK/oBUY9SILa2rHgwxJajxC7SEGwUiUsi9bKu+gtt
J+t0asa2AOb515XO3w+aQ2n9zydQj6mytQTOQVdbmY3lmYTEeJ5gMDSjN2hIqmD2
76b/jkxaXo8Q/STVvBrH+vjcjpIflGmfO+nkSi+Uy9tYcOppEklaO3nTgUqBaCcu
ZGIsKbAKuM5RDjsR9o3mO2XG53aNDG5oOWfwtjfiTcPPtcfQmtUl33gduRXNsddo
bgp1rbBVT/i12NBNA6pqQ7Wq3pOEhoN41nXyWg6aaQcNrZxHaYK0EgqtzP6o7nk/
rReJcoYZrgyWHKPMRb4GElPY0J+N5xEvaS5fjBO9VEWalS7DMD/jecgAO8hlxC51
FRxk829x+C4X+itGjuO2Xk1bvgaC/L5tjohgzH8QN2fJhArVmMwdhQXAgLXUrk5S
DmgHnhpS8ZoBU1jTWvgmdgatjUEAQyD40TuIjXeYW4UIyg7VjXYC9hokjIZT8rhw
2J0x8KwSl2GyZfKZR+k8Ot3da9VOJFyh7k+fCZDWy4zFGvm2YWHvzPRltK3cWy58
wJNpmWPCnnHfF9pSV2WYJEFVs4rtpp3pWoWwOIwhJiw2NlQJbVQyfK+lseVmGs91
1B82msaKJMa87gA0fz7lal3VdUbeUX+JixO8/pVH2cP2tfJmFXqxNnfv8u01k2QF
4XBbnnLbdPs6yEYxm2AU6Bf7+5RjFOED8GnWGzSVMWmyk/jZmjZHA2dX89HKgOWd
RDwrCspi5qI2hbiQNQZpsCPzDshXZ2o5C4QXqrsUxzEjoYLLWz4hOMApg4v1Mxdp
LTCLEgUp26W8CP/KmnxKAbHFAIlCfUW6UwUfUtcEs+TDz+Q0+PruRWOVt7Ohjm4d
QpG20rv/MBfPZB9qisrSKfoP4JwUyfn97G6IL292GPN3i+2TQBydn/WGunfGYKCG
OutyaLhHrvHoYjd+MSkGjrTvI5NBvvaPcbTS2Z9zoO1DhwbZRbGGab3t/n3FxIJ6
yWofPhQfgKFzQIx9GXsT/W2JpPrN/La+O/f0e3D+Be6r0UvOKkd3z8Wrt4xgBvUP
n4xal7ppc4dc56bPSEbffkMt9Ypx54kaf45edPL8q+uHJ7oOHDkY3e+xOx3iENQi
Vyc6Yb/8FO+2v7sSbgsQQz6lMFwO4iUQT76vGvoHqIeWdWO0GwW8ZqK7KlV/K15L
EATipg86VFoQiscmJWA4QA9l4Yo5kqUR16pNZ/bompRPl4TtAfttH+75SkWBXhH6
c9W3w/dc5U+98wsd+EKfWKI8N2zg22SnUSZqsE0q1rrTYOCUV+cRIEV8lw+pQ4pq
7bUp0s5SZsy4DLEoFYx9V8DHcjp6dyK0s0x22nZY3RiFfUxI2IQbULBI1bScFrsQ
3+fgeF+F8g0DDZBXktMxbcgnX3RLAipAdBKOagKjmpIB7XA9NwPd3keUzl3pSYVE
0yoKNm94DJ0wtWkzB8V7j5brs0uhLgp64T4Dv/UF6K9qG6dgnGbRIUPcb5mJIY77
FAXUtqwb2bteCVTGy+F1YacFksD0qVULrbvopRd1aeLTniGicQfAEWhMgBt8Rezs
aQorXp4EcfaB4H68DpBKDi6RkYVVVMK3nP3he09y4Hdp3/pEP1IgrsW8nzFMwD8r
5eRbtIFX/s8k7f7lH9GnK/M7lI745RJ9FRd4TkgMeMv52/KQvTBnHGLnjdFhv4bK
ZEGQsNTwMzgaM8lMLgBTuVudleWF0yKXsop9VwnYiQPf4fIjMSvyqzoD3ybXCvg8
F7tsDnyi4018QvXUD0qG+5Iz4ECs1MKqzOyn/AzoIjubW6gOWeOGc8Aqcih39CLD
ds8gDkJRDKDOOEdsMp7MlwOXySHTMQvOka7JCX3YFvgELtcBHElA7tXCOMToPwi3
dk63eYswtHuKJIw5nsHwT50YcWg7TE0F9OeisZu0dpScFQrVsggAHdkMjWXB7NFG
/AGvBN9vu2HFu4dlvAyChfcY3n6MCHNDsUksDsX5UCs0phA51RCTVWb5HHo2aOAG
/eikdOOcOUcvFk6sXH+weNkMbDk7U34tCm8WX3+WAELgFl8nhfQgtYs9s57u/Siz
wTFABOoBZd/n5+VD8M3K+Abb8aZfsdh6M9Lc0EP4TKbnGum1FE3xZtQff6MKIoJh
xxOcsBN8qQXk1kxyx/i9VINctaFlA6AEDV6aqF0Bnsem6PONet+KUbyckXNtXfeJ
D0jC7JCxDzPxwtzBpwa5ub1d8ppN9gIQ6+JoWSepqbQnI6hs61BqNgvEaKSLNbKr
x96tOhzA3mpXs1pHTP0nkMidAKKtVbm2RtlpaZYN85r48v2fE4jaLq6DD8i7ftY8
frFnhC68rjqQll4+HIEWCiFgqGQcarQZDPLMvKh4Bhh+gebU8aEDdPkKSd6a3QkI
ZKNXYhxkOsYgJ7WmAKj4BHkI9g2DigExiuv0Do/MDf+HTT1tXpqJxSJyWkLw5BNT
qKAtQ1pcPkCC49zVqwVmXwO++QtVu5wnVr4IMcfkOzdvoevX/3aH1daX2j1EXYWg
3ZJWEZq6bGuKkZB8tSalKnb0mKFkEdONlEQix1O29k1T4MJwsFNG+l4yPFcsEcqt
MQ9h4BDGPITB1FM4+7nN6vIVILBK47oG5i2rslDFLe/bt+BP222DIbT3087zAt9/
VdzdDjXFHsAbTkZwkVJ+pNris9lXJjKpgYYChNxZ7wHkLWyIfqsJEAxnzsNXEWF2
ujVh9nCFTDoIsuzyGV30OMVVYOz4QPmF5QHku44s3uvfWxDvK7Ad0KzmxpENDwzk
Q6y+2ngWRokgb1KssUQQ6Ol5dScJSdKJYvv5RCotkiszsntUXPxQRBadKKEuIO+z
hCWrJNTb67Ffpw7X9xQHMrxwjBs5stY7FBr25WtLwp7OqY/2IVIPh4p1D5cOPBkh
ZOblG3MSVoq5ptlBhWj9ftucj+cO7pkSGYQPXqhYbdtOkSkr/PQugECFd0d51Y5m
m5HV8BcrdwtRFqR7Zmlc53LNL/TBbiwc7WkRGfDS6v8XRI05xSFzYVjZ5ptmTmad
IiQ+++fl47mJxgxSR77K/Kxz/ghUb7UGvZKVoyDKLPIBMA7B0EuzA/fH0xCVWlkJ
0VqCn6AtjyCfGfjKrp8WkHS7OjNx2HBMzHhoiPTZ5rX3xI+IfyC8eTIIeIIIoRk8
7NwMBUAczRpkt7bpxJhVI9XbsbAmkQdrqiMuLbXv15hKr1ZJgl/Te6LpLEiVB1bn
4HNZfLz3HZ7odwgpLlK3uUHx3SzBjPbDJzYfa92l1ptiDI7psGhcD9me17T7yUOu
gf2MTZyVp4UrficYKhcUaFpIoDH/nBrTpYOIzVopqGBlyAGxs14Y+z8MFlp4oEUZ
E6chm3M1gleLMK92fQf5LlvSx4slwN62BQoEIpdY1cLA7p0G2ivKYiFriHpiMbwY
dLKeAdf5jSr8XZop+xhk2XbNeiJBNb9sXzSSs5adbTmGiiJZkA0KornHgwhsDDTW
j51wnE37LDBsh1g5q/QmNZccWOJYbMEi/2pQNHssTYensU0jH4yWn1MPB19z9eB3
4JmG4f2y3ivJRbnLgU4w+Qt0uoq9foF9lwXWF+jR5Mtpv7GuWLS3Febnx5mujrH+
uwa65MNfQ4A4pBizXiWwUp5rZXagQxNeU6mLMFBMPtwoQUXUEtIZqt4IAsg7bh1b
FW9UCsaridlmCayijbp/PIwxDeFy58080hYukUusRGcheh7Ln8+WCUj1UKHRN5NB
8/zEYeAB5Pz6a8nQjKqq9J6/OnYB4G/xprORWyF67qdErmPXX50c+P/926rRsp6J
EZTdIwhMDaZtpjA9KTqhZ34/Kec9PA7sUmXSUe7xpZnXe3Q3+iZE+l43dR9k+F+R
r99mLH0sHBKoWcrY2Kag7K9b+UooWwBrkr6z+b3irb0o97lMwRua9q0YhGLGdOx9
qPW0eaBH8p2BcIJDMK5J9mLPWGWpsfmBFfUu24t+lrs7NI0JzVsI+WDap9Kx7VNv
LEv/Y6leT34JdysSW8ArovMxaFB3B/w36JYpYLQmXsMz93VcCEW4WZY9uyu/UOlE
vaLXn8+4eB9+MscrZDskLvEAXaaDqJlWopld0zckhmkAEKCkkPuVYQjSaVXpV+Uh
Q8AlNJGR/vIHgL5zrlX3IT7Vi4mEbNM2PeE8NW8zE0UpP2FVxwzPV80x7vav4wqt
QK6zG3DEcWeWOERyR85x31vB0r97Rkp+ARlNSVfGo6tQeJVLGsmzHijSLXjhnlxr
Zu3dV4ktJMvTFb5uXlaE623CN7+BIJJOyLorrxLT8lp2Yly4gP1UqYqPaqSkqIuW
15T2dYIy7dDSJ67gOduIE7t776Ay2m1x8AM3dkrI0sOebO0HjW+i5P7QynnFKjtY
ZzZNIRxElIKdTgWzHB/ZtNT9HMC+kx2Ttb1dAocSXSsVxRktR6Gcr/ZpHqrLfhKB
OtD9H8zosv3rmzeC2m2rksZQJU3yv0qRAz5ROcMl66xhzjc4PM+USL3Z/wzPuDgo
fxtQlo5VQ7bt74J8OwSujwescqZUpw9Qr/wayryty2xPK2RtmzHiybrpyOsGaoBq
B2WRDhJeE5nPlcFYz+wA9h7WEUimVbi3JcelafHipW0+cHG2KOEEmEXBOT5U6YYD
FSKyfhXXu5RVpCT7gJa4HET+vmOXOce0dKFn+NCubadgbnfFVAPGm49oGhpf8C4u
+slcpggUJo/51Rd7NLvlQ4S8pchXHo+/5OOZpFateN7brt1nt1amzzW/Ej316nJ4
AMbTUfELBXVG1Vjv5ahR7il5pejxsZFAwUxdP9wzdApXsxUWwEcpnuVMb4GAbPc9
g1UNckPY+xd5BB5/M5yZw01Jwm3dSezqIQqs1rvm37iu1G4jf+TCvxtCd5Mgfv5C
hm5Aes3RGyVCk36VzyNJlOiMnQr7DmTFJC0qYPwjO4Mq0B768mm8X/NyOyw/qOGz
hF+omPmsWdzNPMBcpA19eZOATEsUGPIxuSv3hTgnE6EMJrh0cxhd96Y/22KBMnta
NL25nTzUWJAwqC75Xo+AfVSMjHV/gznwxRdNwFGsVbPdyjmoo7/B2z0JcpO1q/xV
pwoW5T1pz1TD1hzS018zLJkLtWt55TVKBXlQxcy76Q5hrQu+cilMcoi3lQ4WM4E+
fvQD071VdJtiBCeC8cTZJS/2XyQc0Va7krY+23czp3W6QT7DLEat2A9PagowX62H
Lyf35wrmnoxaQzn49Y1iqjUqheyfZcWF64tVsN8uuMSr2ZMzzWIFUG7Fbc01W8Eh
rPYJqobB68fYCbdvB0sXfqKHr3E5CTpX1T/qHEP9dUjkn6t9XcJNTsKKNyhtL5aF
46/v+C9XHDdxpUCrHpGtxt7Rb/3p23A3UxPCt7LWv04WaqvmuO9Kx7zCxC9vVMXt
k1tc0zkS9MnfIdrsecO/AbRSBDsKQ3pC//jhTLpuDI8YdHvOVE8EDFM553EM2zjw
GsDNFEx1YgnUgN3qTRCDdNZ1zISN4uei6QKDMBKA/aPN/GPFRhRiBoD5bKbOJTEK
VVD/ZaY0brNsPOj4WeiFk0XB9HPI4ZL3HNJL0X96HPrQxSqnUOYKS3XC45jCunxT
HDE0J4cs1nsVr41sVAnnxhNYZYWL9iWtakPOeJg/WHWr0KZqOUwa9py910v+ISvz
J8FH203C7iEzfJqrc5hh3mERpOPR+xvuhhUk7kinm8295jh3azGH8aPi4xQGwgra
G1fOga4Xi45yMSpJDtYj+X8/emq/p2FcEyr0aIiDTiJNJa1p7SzOlBDuE94l9lNb
Hutdc6UdrKOktiGAjla2IDNNm0RgaFMbJNWx+rPnTX2BqL+Uy92oi0/hrVJrPpSx
F2JD2/xzs5AvFEFCEm9imnRrVls/pEFohW5TQHI8M/XDAar6Gw6tvPz7kWR1qZQ0
wNjszTKM0i91gMJMHj8pq8df9sofKZK187UzXdhAnYBmU0lgnK5rfR9SYRnoZ1As
MWEvMMhkzWHwBA1vZ6yV6EXE3epOV87vD3HrCQDHx2BANrvB97jfXBUeodr0/7lC
0XJHGeC9uyLkQLWDLQwdiga+OHjodKaxp1b09aDwZ916Gu7ehEL61WZHIVucfGn0
4vrPauLDBu0yc6jqwdoMAN5nWtn7p8YIvmmNGs/mVRa9G4LGc73AT/guyYrHzHDY
i8x39Ofrw/lubZ2BGBtFhui++aWibZJYTfJHG8gzxVk3ln2OLRfzwSoaKp4N3Wp+
uG1+si0NbYI94AuLFoxxUb4gKqHF8kZ80nFEu7pWJBajYPUG3RjVkUNfu923DjNw
uWR3FilRjz659sduSquN0sga5U+8GYORcvp9cTwHzW/Xpow3n8X/rsF8EpVuftiR
hVGsUCd9JvZ0aBDljDKLUEo+DA/+tJE7U/As6LES9Dje4P8JMOPVIzpuejgD0Y/f
G8x6D5BGMtc0nHQLh7ooq/PS+TlfkKEp+H737uiaF8snYQx5QEoSH1O1v7XmoXYW
7Ln5gT/9ybrwULvl3Yx0Bbvgoal+GJTf84fppTqwafZEDfwall71RlEdxPBEDTh6
83n+Lqu5/ZtGmhI9zsnbF+WAtaEHxdVijsGT+x0zAuMvRHJYtDeuDNAu6Vn2SS+A
fr04kHWebLWruS1chupOcHGHwhmLrTwq+8IMoZ/+ISb0qAtcDDhQXxyr4h266wUT
VVVHvnKcKvF4y1rx3XIFEA407FiDEJ8H01vZjNWiE/IYZ5fSXJF98ZFq6z8CGYIt
F55PkXNrH4DMxwhwMP9TGuwo91418cyfya+WBgz3ntmWNIYFeowgDlOTRRqccdpY
DMPQ/SN3nuX76jozUpBbGaEGt6nMDNlSK3V0KMtPIW/q19mEZ7IGMmEK1s6Zk5Uc
MM8YvoJXRDccVm1vKygjfrzSMaYFf9dE0hPnWIHDA27a5Om9cH5msLh+i8eJiIKF
1fEHggmvNTlC9wYU2m/Hk0cuG4n7HQ0HMcQ3q6Wulw/KUfXEddPsa8g7qyFMKQVQ
NrJ7yWmYF8v8nV3F5347sjMkavsb3+bJbCRjWItpau6hdi1OTDA4QmxJcFhtZm7e
X6v4teu/gcybKbn1eEyzTX1MLWdO7y54PL35S9Ph4oGWCILKrrCtM6S5L8i/5VcQ
JePGNsEEgNodz1PP43beNYIBCBru9SrS8uT7rNHoDE1xL6KYbeAnbxpfxgp9rTz2
xGN3WX/Ibc0ypQZxn4JuLHteWJHb5kSJs/knfFNL2/MJ25tC02H1An2NFEvUrUT8
+fCGE/hUdF2wKsyjXc/CK7L+I18oy0dzXAZcKs/N1bD8DTkXHxSQx6hbjoYUHF0n
vddFUJbqjU3kxTWXI6zJvE7Xr7+CMrWRLmu+eIIUl6SV6YYIn2TKSeKG5GtUuZER
tOeJPRngYcxxPrwTrL+RPWWl2g2+knhlqvNPKPu9dCaZD8Ae8U7ePSswsLi2VPOP
TESWo6d1OGPt/jWG4U8Bdk1JKrr6lmR6G2ZHCEcBVI+RTNSUoL73LN7j1nA7L+gV
/ppMvJNczGMpFCl0pYKbaxYyH8Nz9edQ2UAj+H0oXhE9sFmUhBp2tDI8/pXdMlQ7
C5OW13qnOkysnb8UT0Wdr/qADdUyXdl3c2pLf4GRilMn0L8SycChxZ7QfjN6RF9+
AheZydFyOsyejTSe0QXJD48c14ONscBBCTREVkXv/pQxt5XRrkpj4CSWq5WKaEcN
HcUbu3eA+wcXP9B4mNev1HPdxE5aXmeXpe1WDX3Sz1YZyYWZC+1LXj+nF9TeBBXl
ZKf0xDpCF7OLc69NYldNYR1DssUxjI8tg03VGVODLiwvTNmAIDodzMss6LNwc4rh
+AiDyxJQocJ4zbyAW+e49TljvC4HeospHHIZZhO4r4mgxwNpCCjqM1S2+bfAJh3M
t0l0hJY+xNk2SYOA8t0ZnVnghjZjRF4sa35Pg+xuWGo2JM+gHYS+m21V/2SfT3oj
PNX/LcJvkgQ6HXmgdg+bnTJnYtFIaI2G6UT3N8FowUsEAIAeVbnjSP9/ZBSa6TIB
WlkmknEELcIr8rf0ra/gIpzSVFn0fn6RXOcmS2Ymom7c7MUcx2JWrRvEydcx+b5h
5t1/VlCM54uwxpRFMz+urZ98kAAeW6N19lszBLvIFyNyc6zyvNH7JzLM5xkLROA6
C8Uo2CLrO+U11w/yQUKRrZoalnvo3yW880ACNIGmFZPgZHZaa16wITtteTZzuZPc
dQQgOfqFK7z3KBv27+dnDD/plPChK2h86/kj1EcuGiuuANsCZaMl6ZG/JKtRKK9Q
I1ICROcpDE2qFRpP9MpB80QFqy/0HfrRKJ7GqJsEXhvAwvS3E3xOo+BNmATvYnPS
zdcvvJD9MEd0RNDpcjCr59LGHZR+qX0LTy9Z1xpsszGT1qWzI09Gm9Z81tLNcbhd
994GMq8XhbIVKurSWQuZOhvY8TjTs/YS0XHOm258/d4I8xZvJrvbAFuFIkq3nLtp
o/4Ayu+hLA7nWbKSa4Gv7pU8c4zTAvg0djbuFrd1ntEPu36lXzXaSoUwRPqiNtiy
t5Zh1ZQz6HstJdu6oUri8iMXmfgo0X3ngrxAs4aEPnEA6Um+ln4o7xEEd5MeBh6U
SyM/d8hd+Z4/WRqCewZOMWaO0iuOaUm9bpzV2HvSs5f7cmzf2Dl8AyR6wZWFIDGA
UHxWoTwftVbe4f3LZ428rN7+XCTUpD0o9MpCwxL8VA6zl4ZmfPWD3tTX5Lj4n29T
GnyoUhulhADVMkipBf3jE6VhldcycQqCRrFinmvCMBCN8vHExSaveKUWDMrlvg/L
QAjLEmt0rfy5Xy+VvjEVcZtzBGfVlHAjfEFfpJT8Z4xKhO71AAKGRllpA5+e0DiX
Posvtm/jD7jqqZdDRRAUd5xZyy9v9Oba2V4dnEQVDsN5AQgd5ZJHBEiTV0B2I1Kz
QaNfs/czfWy2ODSjP9wSrSpFd2t1Sr2ztv0hqQqA0nUPCT1gyO/G28K/zQMSxLfC
nyp3GWwT3WgzAI589TffwFBFoMqn/+5ETdgFe91PjqO2XUZdS+YoET6GY3bSaI/e
+wgAO9P+Zf+qjIrjJmGwxqfjsnssdZd2dzDFS3tTZvdPxlVUdP2R4qWKpuj31Ac9
d/j5PR475gLPM6TA3bFBjOTQcOvWQY0378WNhAgrJttQEO08CDoM6cY50GIPmHQ/
QWOi86MRGOalorYLgcD89jT2c6xX41hG/jMaxQpBw6tO8tMp49RYRJDd0ZdGrDOK
ak2O6ji5gklryNRU6FWKms11uiDfyvKhONPiWe3IoUVhSWYqT6UPhJGT71AZIswF
O2XbgrxQZg+2nQOIxbprxIL8KoWASH4N4kwE3dJpzlI/H9/XPlSxf43VZPEnwCeK
3smv5DobSeBYMYD6nFFdWiFbtt17zh6fQz7RHwMGJQlRDRpMlX4jFKZQeS6H+4MH
LmNF/OI/dy0wt76Sti7LRz3tf9APe5DC7iwgJb+bkJROd1/4pu7BJ34CagSmYZ64
0arql8gBtnf8qGlgpw5hKODBq5r+zZAxK7wcACGjHRh7Mqz9RUppxBNxhgHFbohu
HfQGUjQIsgumQtmft+QR4opRbh+SwtAm8C2brdWNRxy8FqbsTG1zs61gj/Fn0hQ7
ODjMekSDcKxkWOEO5bSemq85bZEeDrRPBrz2g+OfYkpnLP4w2mHtoPidjj2N5UKO
ziG6DzaflnLzyNzqR84huPfcusGCQs7bTCWMYWak0WIyiCYb6Y0XMk7ZqUflOa2B
2WDDG5NFRfgmI6oAW+/muB5k7FazPkG/x+qO9MxKM5pm18gVNfSdLNexLWynYFLE
lwYXSn00125y+AbTlzOxaAw/j3loB76TMCE9fDOmIUAEYPtGC4AhVaW8JrNjJaY0
cP55/+ic3mIW7plCS6FMkC48SueC4a6iSV1frVgEGeAQKGFYLyMhupMXujuTLWje
0+H59LLMRmWrUMWU5UvPI7WlpZ8eN39CaUfOB4hfe0tYVOOAWOajDSwiqcQrYsxY
K+ArzMFfYCZ6uNHgCg71D4GzrWE6NZm8M+v4MJ/GmFODnQfh+8v4MwVlXs/mrDKZ
NEl6wgmM+A1qWN830D3NAl5XKjx5nViFfvl/VGV85mz+Bxis4HcF5FYCK886QxOW
S+nQKix7hc0npOV6AfzmiWRYPvZr5YZHXqHgSIUIMIU0DBGZg477FHXOJioaWYo4
TwyFaw6WQbfitFojSd4UPQNfikP+6DXCTq0v1vD2aGG3Qob7XBcqUEULVgI21v9U
7qjPBePHmBsAjNZeYfb/zYYbRMqjojoPcsoeqtNv6hGRzGKG14Vemn34JxZWdiUA
yKNt56E4kyT7LIlpCAhnIb2hIhGOI6rviVQg93nqEk+PMpBObRmdQ+fdGJbyIFU7
GNRUQf5r7RiYDG1W2hb860xrqrVaAifaVgZLthJpj5nvYLgZ6cMRwGSWIiVTpnpq
KdW3T2O7tEOkQKj5bQSoIUeb58moebDbFkPf5QvfoMKot0qfkBvySGIXAr4qTmq3
qOSb7hbCx7gftUzgQqql1S8UOJztbdNg0jAKB8vCxPbRmA5e8nqWaAE3dORdNNHR
8gDf57AsTT5Yuo0G2WH71E39oHVBbwAM+wiEtxc3Vtcy3saJqOSDiHnWriw48KMm
/6DiPtaH5YjbdnK05vvfp0oLYITIbsWZuhRfnIaex857nR6xEwyL0h3g84sDBEbV
oRJNaF2hbXNPjYZyy+2FFwICykeN8GrJR5jH1DUS5DLMIZfCmKm5tssFABmlIrma
NmxRaFw6m1JpAK3f8m3AM92tqky/q1SEK6uDhw9gLJuEMLvneLFHwUUSZ6npfdXh
wcLeyy2H0Uxjq5RbVT9HAwuJK25ceh2mHNMe9dNy36RXH8P1WX8lzc2p2Mp28NLX
vFRFR/hGsN7bK9cSh2BWsZgKmwYxNJw0Tvj2Wxpo9OQn0urq1zLQct0o7nQ/5VcT
TN72GszygOXFod+6BwhcVg1K7gZdu3yvOxPZX3KoChMIBugowJmLbXg90rHhL9ZG
x1qgAunH8sAtY7i8qr5BHk8qf9XBViNe8sOFNV0mye7U9GHG6p1e4NmoHPvXgw+9
Hf7nAWGQ/G1eutIsn6tD6P1+lzN6XwkIC5nxtyH0gnGtQMAjbJ/zuZEB5PW3zKC5
J4mw1aPzYA3XVDFMhTRpY8TxTECchhvByggDLA7li/TKOATMN4lQltceCgPacuM8
iVqyy1XNtEa9OsFjLgxb2zSecsB0XCT3N0cL9EnKOjzUYOn/dtKUzz4GGJTk838b
UB3NoOuVzmcdE0B7nAjalnV8opKE5HW5wnthJNJITwB/YeS6O94JC5sOypRntoaC
D+ebxoPdaATFnn3drxEe7P4Fii1ZRl9xVPtf2Puxs/hmbJ1zRUfse0AYsGYmQ2Kd
DoN4yxUainlDMeFYWKyz600K5j+RSEARo9i+UWCSVvFiH4f3awfnoxkn5Qbv/Xqw
Az17a+Bcd8TlIpI0M7f9sVYj4vVJpAEoDXL5VmkXRRROm0bhO7q/k4lhrh/teA3M
OexCjHg07WoGDxFTB81xCYO609rdxTUX73tCARR3DS60FgJsKRKhavhBmwyeQV/j
Kzv7TjADxGUSWaE3vVNvuZ/R6uJgAbplywAGeE3bR7gyaeCV+9FBb9cvBS9NG8bW
iESgLJvGSjgINRU5ONQ+mohVgKY+OIN1EVH9gHp46eEwhRw+mT7jZ7WH1efguD7q
ciDiDzl8Xxa+Ocxh9ntMgsNSUy8OHRAcxtO1PCAj4L7pD4DS1AudjEbhLuS96j5C
yDPuKISZRdOSLeLZ1b3GJWhlY1J0AQl0hLK3QwZA0V4TVtsa7cbI+TFNFni1h1Zf
mkkjA8/BbNFqrcB315xX8SvLfZwCVRRiczJ8TPAdk5s1Jq6owoA1SItHF5I9sv5b
CMVxc00QQNReXFrygMRwejQafVEqmJY1eleLTv0K9RADTVc8TgDGeqlicZp5+auD
BTceIl+M7qnPHEd1c8Togfy6EF3P9NkPWQmwxHa+JiFOTynEB8zrXEm/w1lLRHdk
paeIRsMP/d8j235eKCyp/+EbOFcDTimWpNgUfM4soIJqZkhPXHNNp+01E63m4+u7
EJ5LkEvIJVL9L01PshezsYJx5F8dFm2b33dXx++kO95f86ntH+bWaFVyrp5Wb1fd
nhv/1tEwnhmWjE+vflu/Aiv5nqq6eqNcS5sM/BRR4qPKfWWDiP5T6IhTW7+9TLL3
c3eG8LPT27+UQy6RyFvp2WEx7QK+TsGT/PKSM4/9vXBfFHi3Hk65gARdBwD377LR
p+Nso2twLcW/rV71mgF1HbBTi3NipJTJjOT9uTEsc93yFl63R+b+5EHYacxgZYth
dh9iYmq91CT6tRmwuZKkqAxHLzS9oUnEplrWA297sgbWDNf3yN1qfqQsoZ0HNwCp
g1ID0FSep02jxsqg9PFtfb9cPqThQqO5NyYypA7pnpmGXLUZnr7uPnRWSo+C5v/H
BaBfUYkT0w64rTk6Pgnsd+YWod7RQsVjJnrY6cell6Wbujc4sWfqqjZOq+wxqLoA
xMPs+Re4bjJAAyM5N85efPc+4zy8mC4kQgDDShE60ermX131BT6/V/uSninOu9XP
s6uXw6/2tZe4C+4F4e9CJKzgjrB5cceN3LTdLsj+Jhwae2C1+XisxXhM2awFw1KK
zoaBhcLCf2Ej/mLiFY9MqiAVTEtARLDTpG5lydITwmbe13bAVLRgSqYkX/97Z+59
2C8if3CpOdJ3sOm5slmVTXGAfY/ozksXCiRdNeu1jWFRP88TcyBDaxbqhhGiu2mb
lNlvDDQU7KzD652PvG+vScE/1SB5RbeMNz6EVah4MsAlWLO4GAg7w85Qd18e6YGb
ABenjRiQFhUumn92zJKulBZjmiERvxVfrWMCBJw2bgQiQkwBbQYjATaGIbncjmt/
aZOyWf5BsM+1bEEJyeRTOZb9CFZPPiwoklb6/f/xaiuB5sVdLxpHiC1b+iLqwkkv
1AmxBIfDJc0/0Us0qwvEuF6xxR8QJWYqHFe9cRMJ045rzcW7+yPB2IP6JIxyklBh
vZoxIY7bL11ODEh7Zedki/2+CdMrX1/cxXul/PxZsvUHEsi4L4SuAB1CwIGpl86c
2eOXaamjEoHukymS3vwpOURbOx9XQ9tnLIqMCJtNrYaIwejjRtcLLh2U+QDx7DY3
w04cy8cTDHVJjbxbu7DAW7Ef9unzzWM5vxoFHeLUdaEiUz75rzlYNJ23U35shdSY
28n40RfRY4BHx6JMxEGzpzhSi7yDFY00AFZZ17mIr5J6eXnEg0k41wjmmYEoVPWP
qGt97cavyymBDWTZyoZU2/5fP+804Ov85L0ekcMajPqVvT8O2svC81+n3XmkUOvl
dY3FB/MATzMSDpGMski3TsIG5Q3rCuhaCg5g07+2dvmGlw8AuMwgrEZ0ijyW45Li
TFRB9sH3ih1yNjcrOJtr1wZSBtFFeHcRGdV9Wl/fJ67vhOgoDG1X1KZRnQQtVV7H
O9DjFWPAHV56CGgk5u7lyBGmPnUXaDKxEvPSvr9+4zXabVvdmomAl5y+gSrCYNhl
ZevwSnLD+VvpkajrFLajebQsOIzwi7QVC7UGhpt+x77fUkVJ+ZBBM4qije40YRV9
ZuEF22AQc+L70ccQxmE1VBLuhp2STZXWcf+Gf9PIKrYI9dJGJNwYRuooZUHAuSaK
nR4IVY5nIO51DKsJQYwafIVi60M+HHMtdqm7xl7tre7qUG1Qg10S+KrMk7fWOs2s
yIlfWE8HV8l0vhkHuIjhinazHzhyg0b3gCMrY7BZOhu6ESRc62cJDM6l3DyYZWU9
JmTiBLchwTFV+TL3KTf/00eVqucZS848SA3EMxckDw7Dc6JwFhv9sPhcRIy/bXLd
t6wjmvBvplWYXbFK+V8zayGYU7FYFUHyHfwtHp+dfuaQCK0MOs+yNU06n4T1W5pf
0b9VdHTmEESJbFmuc+VyxGpp+NLytNj+czuSYvJ41VhjjtErHHiNHgOJ5M/JCrwX
Hnt7SBSLgB7Wom+a++dmNiDLQsG0KJOdAEddbppC7UzvBzNCGJfAQx7qILWFmMSG
HzGWospYaRZlvfsVAorbI6bxfwWoYSJAIZxMHRENDPDCLvp2iC/hstbaUTMVIgeL
8lnymubZfRgLr3KFSZNIjEzCVwMwIXL1E4zabPxeneG3VHLrnNd30yi05iZAkuqA
7Qut+A+RzqxFEh5wh1M4Yt9VqcIaet5ipssS6u4wXFqrENBvlF5QgF182nw+3Wiq
7fzmDfASD8oRBnswrlL50UBMLlFuIyazQwxxRLPJiM7a42dfFchElnl5rA47NZR0
h3hBo8fTPjY0jzSDPAFNCSRtprAVvsJQ3EpPeFFQrOPr8Tv+Tk2rTCFDTKiVuDyT
HijZQxeLLJw2K895I1RniWUehadkh9heJ3KSNDEHllTLtXxfuGuZYTqhQcDRLxBW
8pkyVVBsNqMQg5GaF3u/EuTA7XeUOwj5aMNI6K5TY8bEt5RnMl9YO4JrBQjDg1XP
d8bczPyUy5Pyye7tddyEsDjyf5gtqKwKWmXusBNccXUeDt2Tt0/4evYft9c3OCRr
jxC2lCPpuV7qktDSj4T4PFHKiVuFGZxzxD6LFsF6ia1MmeoA34yGL0/1SALeOKLG
k2QEkJAnuprIdUpnFE7uFHM/pmiH3m2vEeXx7s1JVH8bMq9FT1tWei2DuFgNYN5H
dF1EOQ1nZWslaoDcqCaFvLeY7xsnfGWKMuFZ6ghyrSktnBAE5foFf0glJMD+z4gf
IswuSAI/7lAqLaOFZKj9GMHgyqAIGodmti20p30QwvxeGCSte9XmmFk9jxzpYnv5
Xf+lJ2vTucI2ei2f+wHdK4TCxctpQRPq54f19x6/mHnBmwfQPAScBG0ncLm59b7H
7xHGIo4TRcEoOTMqfyS640Y3U7Loe+JWCnCv0KJm9BNQP82rd8nFWG+IY67RbEsB
4XIXeKrYfk7c7SsLTOfQ6lPZQdbZWqQJLLmDiQA4RbcC7p18Aq9kJ6pd6UV9BbpD
36qj0cbn6dmQOczyfZIUYPwUEo8kbpYsux0SxRuBWxL9lGuEno/66CTW2SqSFXDN
MdaWtIFOjk78t4BMItru9orbalJIpL+d1X2dfNp7TdOUd9Vjgur7mzJ/QVO9nrZK
iQIiO5yM9hXAJRJvF1XznDATd6Wgx59l9qzWx+ivecYetEUppsYd5KRqAGpd+3zx
YDIpkeugO64ha89qYCkreKM9YiJNF2gSkMjZZ/f5gK+E1wZEEQRlLDFP2CxJLzbD
2uiwxv0yxYtkNADpWAz+rRJlxQgTLkl7uOwJ1F7wt2jStlySwYYSv5sCqsPCLidu
hilEtNCkGH/uvNcjRNNxFHuPjEXQh9ql/IBr85SM9hYy2x+/aA2W3xdQnoInzlZJ
1C+y/vfRDd7cmS6Wjm8lfj+qPyUR1tCl8d8nMlB9B9UOPX6tlvDM800Gte/KshZD
5cYuZ2cqxP+6FxrpliPizwkTlYi/Rc3BHkffz81rkMd1mKHrpulGQ8hWcGxfoY05
//ALA+5Bbg5z8vf2GaVG+MneLwqYghOSf5xqovneT2FVzSn/NyrP7Sx8JQfOvIVS
Js7ycWessGZfDbDnuWbKqASULdSHxBRfiZmyKzKXYC0nXHtnODo3ovYIoMdHCqx+
ewxaJXWELaZ1NkKFplU60uFBTy43yHeiSBzVCp3LybMcz1vu0QL0ke6D+9tt8NrF
Xl8oZiQ/Xh0UBXSc5MWcRWzf5IeTBL5S4Bb0MOr6vQz3Gu18IEp16DuxbY0nV6qf
h9N5gaAgDU3msllMkaMRZ2480xLofLnjxtObk4pcq6lKKEsG4DYWc1c/XYqUJjI5
DtWlbV2gGBJ67GYCZ6pLcMfdzqeix0upRdpcbTCes5iTxC4jp1N+0Xh1beEROzzX
Ve0CRJUz5mJXdRouORunD7DzC/QKW/AY+VgHt0hBdUDNC4cocbPUAndbaRWQ5FSE
MtdFsnqrWyQMCI2uYcDbLSTjyyerQUSsnIf+Xhm+RYxbBf5zNGL6RmZ5LzN9AxJK
eIU+XD892cxJr+NPfDbhOPPpwhSg/6KQ4p/m9QM1yAOsgJ3NRoKWj+57/cdhlxak
r9/alLm6y1nBjyfEn/bB8n3dErdrLA6tzXMpl6fXG55vVJJNHJ22A5K2Zmo8r268
5abrTSPZ2oIAE0bA6te7VYBHBCwMEEK2tB7YCA+zh8LyEHZpoCrQHfs9iqBemL5Y
Tiu7fX5a1263o96IqQpor68PuD5cM6EtBlIzJCiYo5KEwplOsAFyE6Ph7I012HpS
y0xGcsHzZnY/dlKxwilzubfIcswIjpDz5SZG05+vK83NmCGhczXOGfaFl1ctbkOF
+ajGvTFUp7G8uleorJLhDTWnxx3+GYI+D+9x63zoVXpNMxn1BmVHNa353mNOwWks
RR4LwmAOcJhM8FPoHvA0Csi2u3lu/vXs5Ih1uKahRMlCqZw3oWatYHVAQ5iUocgR
XIip05gHRAxCiKvLarMQR8y+yWYGGYVwGt+gAsf133cP5sksjbFQ1mp9E/CuCFVE
IDI8yuib+5hnR+KXKFLCJ1K59DVktebnvXH4zRkA4c2sgCXQ8XPcARVxre4XNaDB
A8fuhVeWB61wf6+ISZEmRETBO9D1KU3bdB7vqvwE10KJDw/UTkFX0gSETjlZAl7L
qFcyvawCiti8dnaI4cxrhhblfEqgapH6WEHFtBdLNmkb7ZJt4ht5hlEV8pgZj2eh
+rOsNATTZoQXClTcp+HRmbm3EIFWnDG9ROMv1gJ+YvzW31bEdVcl7B4pLNBpu1oJ
OwF+/aNHFngIRMSPZ3pakQjjf3pj/ApidtVYn+VHfXu7GgctJxrDCBRSf+HXYPxV
Tg2IjwGB3fwNyaMCPzhcnl6Qwgsomv/D+R5P/7tHkUFFkC+gWVaRo9pF3EGtUSmL
KuyY85lbWL1irfxBXFy3safw3GmvblkoPzZNm9eVy6CyQBjDRLVIJlfaeJfH0QDP
BBqhNB7nUl1AdZSXLtK3Qpa4eHFEm+P4JH5hdNBJP8EuMh/hIerqvbA9dEs3KUTd
SrKJoTozSaA6/LuCh4iN07k+0TZgidzMvOJFEyi9wckasfXPj9TJxrKi8HHK657v
1/+Kdtl9n89AH8JXQSRP3V0vZbn4hSjTp8qqo3GmLYlMLDf3gLzP3tliBcIflncg
hgNOsVFNFpBxwrOZBkpo3sIMRX47sBTA0epLXo8jsvgLZCIM0nn/ZGKBTxHXT/Ej
40Mah7rcKp9dPCVqrl/4yjBFrt6lIkZwLHJj77pZQ2FkwmLpeQ5E/DgS3sNZhcOS
G0I2q1g8w0iLLnoa47uFokvWKjTcdFcNSkuQ51AU51zbbSSgaGQv7DLmDk3czc7f
bSkJO8JfeezZe7OnyZzQpFUPQy7/BZF504Z3hEk7Rv7wo9ufy93zcqoB6eEb5Bes
oJupzQI7cjkxOrm6c0zdJ8YMPRIISqehA7pG0KNcMxGLy54FY2Urv93MPD7/7kJU
pqI1Jn5SpFLogRM1i/rDL66gaszVEZDZW1bl9hBCWbKZouKuLdsBY9CAq1OJ2n+V
Kdl4KhZniCks23nreZ8vBNLVi/UYs/g86OlDSsnXUIVDPtagcIwjfuFjRkhon26f
GRK6ByG+gabkNbAmXgUn2Xm4b7qa9lGcVCJU42Go1csVLAkrBWGG46KE4X/9B2An
7VI1zL/68q8THHMvOI7fMVLXgG3tYXdxRbzv1jX9DfHK/FaE9SRdAj0cQEf5MdXd
MGE79J8PPZ+e8qMbd+UAqimxSghMjjR/4b565DrLic75rgGbErjZc4pqO9W9kV7L
6L53TIMweY9bmbMAnpOPA7BKd3baEbMPNMQhhIWZ3sPlC3xv8hcvg1aJntftMk+Y
7y2hKrFRS8OPOUdhUoAwrljQIAPhXx8P5mNaymTHVwFyXczBIzzmkscoKHi2ykC2
0jIh1mNfPUV4ZLFnloJpdmGbkpVrqKnbsLCqbktKEfPvKnKD9Go7lpLT7UlDXU1R
GDFofDxHyhkt5vLS8mXcqJqvs8mVAmkwVnoLIxFg4GNKFscTay4a9NyJOVQFK9Ev
37GoCjR/7ynpkEQCFeAJJxMSfdvPtvhz0CAsW7JLL3X2ahzxnpXiak47sA2Nb+Xu
0yj+2MOggjZknVG7010727U3OKLLXjeuyCfHn7OsN6eu+4rQzgSxnzqZhUF/z1wl
JZXW34oa6CJ+laYx5P8q0H1/xktOyPQFWZvpZNnogT4BgWCTH9ceRHk4s/y9n2hz
Gf/W4B62ibqXSRz67ukQmunamBgujgT9XmuLpSc+tCkrym+XTQwA3KHGLJ+3BkYs
dSLaqomWwJMehRvMTlxKIi6rMhF40yIQIZJElbw2do9yOpAHcSTxIXWcz3YPKKUY
GjSRs7HWFvm+oRHyPmJS7EE4raqQodqeXPkosxVqNF49gFd8vNN3ye1ZJnweAD1A
skYY62GLVxP+h/3Mj+4OsD127z0bK+Qg6woxv9hr8shyL63gWd1E9moNfeYRlRPl
wcB09y+3IWdgSRjcJIsJ5Idf9IsTEIMJSTnmcMuOVmUv9yYPg/z9p8fIpCGRs1nl
CMVCVt0oZ8/um8qh0dyWOz0sjiAVSElKFO9uwc+XolsCtnYYxrAPR59Gh6uvPXFE
ctdInpqYWlArQkvN2RNfDNkeCr8zQlJE8u0HwlPKXbYtfl9LASDBKeRzh67oiwU4
x8+dMqnnRNlCQAgJDqSsB9saYdHlNSNppHV4eLWIZ/rltKls6xzBbs15j6mZWzTM
kX1Nw7iCk0gXhzsBsTr9P/7R3PNxgOW6wShaFwm7BKXaxQyCVgnpy5APkSUc+o/D
Chg6lgf7g2ilQN9X2paR1Ff5VjxJhvxkoRwTS3Tdg/EFe+EmhPI9Fnf7K4Pfc5X4
fwhjUR7SwAKOK9dxbIrFU2EoNeWlYGXQ1OGcPkf5ZAXMXnvrHGwQ1W5UGDOnYVq8
WGpF7rqpStqvReIBZPuu7MCF8nTiNZVITVOJHfNp6LY4MF+7xmFv3LpU32P+k1tO
ZtJQH/hxs9a1hBy0KpIjHwWbIF9vT46ZwdgAalcmf09VPlCdGzT90NaplX2AcUa2
73Pje+0o6238pyUseyTwFOVNDIH7Djhi6ltFkiepdDZ3Ou9u6JP/Mn3w5KwMjCwA
oVb1YsN/rBVhZByWKtqb59KKY8gO6l+l0LX3uDgavNWWmmVECPvyJImbEiVKnS+3
VIKn7HXl1R6vFYRNB8WCSStfG+MtEzlNWRUK0uHjr+0EEtUf9rONkPPue2P6mmnF
/7spA9WCqtPyVtNiDWS6ghiXNqmzG11I3iHPggbBODlnpIwt7UX+dzpFvC1qU/yO
Q2Ux4cmWohkqCfLc9old4DU2apzFugkR/UpaT9zkuzPcYPFAhgr+eno3pFXUuTMk
WL9MzsfXAUMvYFjLjN9bA1jFT4zGnK15UBhz0rT0oFgkndIXf+j9egGGAoLrYNSi
eMPqDJf0T+pqSr3aUdIwF6BZNO67l8trW7RDHWlrdDZ35ONWDtUsr+8V4Rvm+vQY
mvQjbs/ehtROMXtGUvLJAY9BF0qUxBUzRRa66FMdarieXOP3itrnxxwqxifvc2aJ
3R6sVL+IjlJOma+RNgUbSmcnQjLQE1GZ+VRITbvPLb0FeBDfCOUBbt3pGusVcgpR
hV0DCr99i1773117S2wevrFmGm9ME/svUM3q+0NaAQh6Y8my5rDQ7ojmd5qv5FxS
pETt5JW/TKtX6hbaf1P8lRp2287GZQuUx6qO4q66ZLAMHx1AY9PJ6eemZLMEmwVB
Bse4mQdVyjNmcT5l7GKU8yWYNDqrbpIkM4o+AXwxVuyotyFBrgD9mhZkRN0/JbRv
KQPeqwbNG/5xXl1ldpim2WN20px30dxX3lkwVKm/cT3WxlOxAmL+QRpxi4l+/YA3
qtKrKlzYcaOGjywKIo11xUTqkUZgSIMXBDD+KHCIPXbhwerMnhwO8mNcXcz+9cCj
13U31zkZjIJbnNZECfVyOoTl7evMo3c+7WtxQ9ZOdFaT6jZ7VTQp7CqkZTeNHm77
up5CbSz3IL58qLYrH8201uRpNBlWB9yW9tn1tmuTXfkdx5K4ez9N3umBr+Gz+pEB
H6DsKoOBk4O74jpi5FLnZYc9ZkFlhsshXv5pCuyJ1cndOrYdHuvUqDosR/sobDtv
1uH7EoQGNKvj+Dl7hIQfAw0MMiHid5WJHqrcZQROlRdD8BfOJpc9e6qHbF3g/Pfq
uxND+Bi3p0JYWpP3xWZqg/+lMIWWx0Il9dmgYaGH3xApfw6PfxejImSMvM3s3A4/
jt78LAZXxFumDeHHCA98zxkg/FiF+46/dlh1vaAOtvYjbSH5Unc+GDY871waYDBe
+04Zi/8JlWhlqojneiZ2NiF567eVLSSZiqFUbpxRsrE+WzdkA8DBY9Bd/Ps8stHn
IhOt4wfdVhf9I2QagPeevAKYLFatHno2/WnQtmUqV+Fu8CRMb19Ql95htogA3sIw
2ULkdwCVn0rLZyPjMmQCVVbJU8AbljjEi353z9wouW4JQXAhWTXwpOpm9HS79pGr
Z1gvI4brHAT/uyRc0ylPyiyBXcBPnGJtscGYs0B7oUXHOEyYvlPoRHi/L4LKv7Mz
LSSAJAPd+Wqg5nJASbTB8QpJl0J8WKqwjZ9fyRDvcHQO+7anvwPIbr4YIQES5+0C
pdTnoSQ24p3jAcGoH5h2tZ1rFUBKJmOs3XMV/Nv7ibVTgJA7SJGtDFwBKiV+X/ep
o3YN4xTLex1iakmqsNj+Yz8VDUofGy/cC4uzYFzRktXCwT68ywTKiw3qbgW92c4T
DhKQdBRcwCdBR60LEgrIVoc5V3UsEsCnaSFN4IZi+nV0rDBuHPKKOTxqCMEqZ0oz
7Gn/XxrUXmXnhvFP6t5t8PD39SRCi+bYfW1u0hc3WQ2tnUcXLERzBwcvR4dz8Ee8
+H1dWKEmVdV5TRq86A0yJuDF8Smb+m1kMjSiJRf1RllZ9lX5Z//1HCKOJHyLtkAZ
dXKqv8x7PnrjN6BQI+RKcwCF1e4WLipIFy7PrOHNRZUsSih8XzHr1orZ2xBuWsbk
4rOxVCi43EbqEm7nlYLJ+i05aNGfQfejSh+MNSBrd8X1hqvLvkmo7uTj1i3phvAA
N3rCmVTQwH7A/PzuIyicLgV+YdxVkNJFOUr9vyiwtFDyl7E0+XBkJSrPTHy7BGnx
mqPZ/Op8ZuGyaz3gv11iQaxvBKaNgYNUfcNynBtHhQMntVaqCjCayedtWaQgAR0+
GvUje8Kfuoy5VWBky4Y9rFnQu9BaTckfAESC/lcF3SDQWn8T3/KQ4doGMGTYXKuf
HNHr5qJyZfUct9xYcuSNg9NQnMAeHUOyt5M3nbGW5PMKPyUQ11VdXgFkJe2wwZJx
gm0KO8QaEsbTk/QpskCFY6n7Bdy2XGJjDjVVVGkQzRyD/TcKSC1wmY/aEimBmpIN
gauPgtnMF3S23yv9sLfiucNPkU5uhXyezD3K9pSyl7UE/gxBdb/dNvtwO7kI+Riu
VVY7WzUV6HKNidmqjaj276E4VPYy6Y02hMYc9yRVKjEEGIoWrl4CgDhGtFAvUlhD
Mrcs8Z2QB3MKu06jm9RV3r7UFcfsbnjtygkRFu2VQfU/okUNi3uj6Q+e8A8IxaW0
myEYnUzJzTK7n22PXLKRH30rgUlseQsb4+ArHM9zsfpW1wmklOBXb7+5PH2WNSuw
xWMd0PqB4cqaTGlfLVnwDCM9cxRxX8IShNNVhoUsRhIy5+qhnhoJVK9eVYWAxkjm
qd+Q5cuM7PG/PbhEvFf338RZo01M4TtyjScKGTFI/0Xx3tvOJ452x6OW8Wxi+HGg
K5iwfWnFXj56dYtJS7HcujAOgEVJgxtbRr5rtW/0f2p+lPqspBWT8d9H8vINeODm
XW03NxSjA4nhvCIE099DwGo7rIiK0Im6O0MlGo7o6tpdvq3K/HWvSzmTUiJTBVr5
+Nl4hPau4M+07m8XNzO+gHmQf8wg8XVxrXGI+3Ya3ieeRFAiOzBilR4u+g3ay+U3
j8Ah6SyBeBxtTMmQm5LF8No+5SBbHrTE8qKpmweY3ubSwFOsFjMpd6iLJflWOAWI
pNFvCA6rPviNEBu8xv9TqohbK4um6TQOzHfpSUJ+Fb5x7MZTHtFwGp1BNEfQadAT
GCGaMO6VzKkZCeYPQ9BAFGLOtVAV60+OcKFNWTTSJh31ZTgjqoh+ZEKsIE+TYhYZ
BvN/GuSIZ1V+NIAMWvJST9QvH1otKAWiSAoG1Xh9dwGpiFyqwJKGw3fCcygiJSTy
ojix78AHI2Rd2h0Hf7jPktYG0iXY/GPM7zUUtkrgHHy+QGlxk8LK+9kmS9aQJ8Dl
jFVUilhY9etJnCGJYV55ks0wjfrhnsttkbBq+pC2b3IggKi0SPgYKkA9/8LmHuiB
Nqo/aErMTfVopfXCQE/heMwTwn2JcP25fNPKnL3EQCR9GiIPPmuw+1AVveyvfQHN
FKooVaL7auIA8MCyEIqSJKXB2cHDXNhY/KRnQc+MKQsq0rAtZrHOArxdgrtUorQC
VSRmJ7dL2BTU0kzpXM9nKo1YWLAhJMnd6NL7YmBCAYqknhjEAdisu1GIJaE5q+in
x21iygsXsMqC7nhZSYvet4todpi81byBvkt2HvNimySGgIX/rkt4OnxLRlkOZJU0
gGL58GBZtuhYXJVLeh8FVv70mWgtmTbajnpTIs6Xv4fzeonu8xBsc1Vnij74Z5FR
GY1GJeov1TRoS5EStgDl5bbtxt/WShpqPpmhhNcStSgTm27S466i/hj82AzT69/d
Eiqa1wZZsO8cL1VZb1MGMSJHmMr5PVzWhWd9Qt18hQi9Vhfzk7YD+sLYQt2O0aRM
NJVt7BA6S6P/A+a20H6Rg+gblE+D1/i8k0xrxrDkISQHRPP+02TIcIx80D3glVbv
+p/j5054BNgLSxvpafNe5jb4Djb7LEdS7qUXQVbBT7kBL3WdCTM6XnkoN/v/KBne
EccGBHRWeGgDL9x8OU+TJ5b6DCnikDbX7BfmLRKYBalu9pXv6BZEDaDXhjEcqfdW
M9OsRd9wlMuZU786hECuDEaE23D6bmzXjflUiS3sQvVHSWj5uQM3wkVcmPY3pvwk
7fiSSogeyxyeY9IulSVLgc1Nv2jYbCws8oUzO1IJB92aKHTU0mMcsgkmPnq9yhOA
DZO8hwK6dnd4PYilAHJvhUZ7k4rvvISCEEiWSm0a9t+Fkpf86vEE4s+RX2a/ATLT
wjqbMw0S8g/IofdmWlmSAWEwRnMXecbJ/YWw+UVHmUkmkqO6qc2Y9g7iEIxmfbq1
fuiHeMjKtEC3del+ytUpWSRuGsvrgxl0IDnZG79qtG8IObn71uea4MxX8Cp8UEjJ
Qydm+/qiXIxq/JSudhNXpGLqwszStCppKBRCCEbjUa18Duj9Depwn9JVU3ZRqIfW
wUEfOKKHQTOG27SZwZNXV4rjICOs4p65rVk39kc9mWEnTXXcyA92hBnnksNjjjU/
ieZr4maubgPCC+J++bb/nxjsbvnmp+c6Tb0I8PjqqA373jGvbyls3Z6R/vHm4fZC
7jc9nNy/ZSIFb22O5IttI3n3f5R7pi2vzPms7xURBxaSZxkVPT+8UtFtpenSVryk
NbdNg7qeKkFY7WNCkCOBNMho6HeVkl7AzW+EP7vrf533fmMCfeR/WDoIoal39lL/
2KBnZHXwFdiC7QVu6xNkk54k29GzAgbKRmzRnfo8hG6DkIZCrUvzVKYvlqOPcLM1
C1VvIf0Q92Lph+MdQcH9JBP4O2vAYjvSa1lkUDSANsEVMfR5qoBIxCEEbEq7UO9q
cAYRJcSbrTlaExX5Qo2GLp8ZI6JLFrir+dslnJHfdfFjl1hDCUJdxsApFmsKe5Bb
6Nxgfh6bgPgI526X777q74Vmmqn1wIPOU2Rd1CQxyH5kqO4u89c4mlzr6jGb8CjP
WWkD9tmlQCbrEF3p5GmI0E8w+JwD15vXHjkTYTiqNQB5Ty4OFNwARgztcuyYZoGV
gNYrgoz04lXnvLwwHsJt1+tnSmfCeb1WiNBXwIj70vRYs7TjjK8f6Bg3SpXFWVdB
Ivhfv4sCdlZcoNLGcUxpYkGJifTEO93pY84q2u5ZteKJULAJuBVKoXaoQ751vCo6
KW1oKiL+J98+Fr98C0Gds+Bk6h+E9fjpjC3o9pdHxiCJZX1s/CCMn6q+K2IwTc8I
xL4u5seWecSMxIcLEvwsF9ef9jtETWcfRQF5m00oX2h2yU8K3dDTcXObqUE4W9cn
8BwEhVhcgaa2L4mE8615uEjtMB9A9zwWm7eSKg7csn2plL24U5SwM/6BPZ3JPtmz
sus3lpO60JSbO5PfKW3T6OYb3ZMS4GV+GFfj/ckiHubFpHVeEI5n6Rj9ALcUDWO1
e6GK6hzUKXomakYdMtktojZAlfeImSuQT/wEWlnqnbzTUFhsvJ0YUYdb2NotRLsk
SwNzc/wmA68Ss4cc3Ke2oWcegcJR6h2LHPNrNtbQ0XZRTiXuA0dolvCFEm+tB654
Kg3t1MOQTE7rH3po9VvRIbHmR2o87v6/V0KLYgvWe/ipoCbEvA9zszybjV2MRK+x
/6B3kF4diJFGWUczkNBUP/PPtE86efsbDfHR/t4JXvJi4kW8Kk8Sl5oXbr+5dPIc
4VYBTdCDJIwRkh+t7tc+9V2rFG0uMpIgEepx/J03ypxcn10VzmxI0MiD7myTe5Ei
a1L3xcMAJLbwMvUvi2DWaSOyeHFugrCa5YTZgpjDahPEf3X4GaIlbXhO8Ya2QXzq
4mKwuEHvkkDNXt8QZWjex0TMzg3CrY1ouUu5Oj3+cu2fIPZdjNdx6hUsjXuOQXPR
52Y7jheSCrjrazyFrO2UblsbS8oLQTTxR/15ED/9YXvC0xvceEfRR+omsLVPwQE/
fzjmUkdF9lwU556j6KEdFGwn1IDwYY7iJirteSRV4QmjvA3zMnRayhRq2K1AEgRd
s2czf3w8ImmnoVJtGHi+VtN9xzMX33IbVH8CQdxTn4U7YDLQH+CmCwqE1mwbzOUZ
uf7XCo6/6nL6UoExQLb6ownZQUNdd0LRhTaiTfZQu4aBbu86h8h4eQwZHSXZ0ZCV
OAEbEmeHQzeMZKYVVGtiOXFeSYXNB5ZvlDbBeTBBdr25ZgVZ7BZ/G15Sccu8Z2a5
y3TL0nFrOaKniieUoF1iXgU7MaYBhR3BDwkKNFeSUtURu9KX4rSeTudWXPWWjzF+
MpBkSFHQKvgWnwWKe2N7CN2unRbl9JdBgJq2hGjBQ7d2jaruFvT5FHikrqYNhkxa
SbifKfIk/WoJRHgg2FOB3F1vo46I77iMp6T7xgAramFszCLpRZzgTWN3v4lByTsy
tq1pF7JVXj5fz1qV/i7Ri3Ia22u6O86ZM15S3LV2yVh+ipeykcq+li+PiAXkZ19m
XCc62PBNMdzzbznVjGh16ZdG9jMkvkpErrYieRmZ7oa3LOSIUbsF7ls4tK3OjrMn
t3So8fhsa+e+D+4d0RUOM4I730TB+DQEuQwlgwrYUzAI/34vS9Khna2zoBXDHRE2
E3B2TO/2ax++7NnMfDpMqNsq6ciM7wszukNAEBAVTU+QLVh5buaoagF09deq0wTt
YNAIxUaXF8FK3WU0a2NJo6OW1PG+nJ5iaeS4qPiGvDN0ADu4uUoGTU/w2Ff0udnO
PNrPSf9ta3PSAye1hfvJzSCYYfFvTG5HxONzN3Voo9gSb1OygKqwWA1QEO8HjiJw
VtfFwRVcEeYG/KVGKa16fugdILPjGrtVpUDf+FTdolbhtlpAwQRbErzbSFtTQewl
mGCMuYeUeB/rY4EEPzKyTEFrUI+119E9KvDZlQjeOHLNisXniDxo7aR+dwapYu3z
y0iLdKoaUi5zjcoS1yCDeokMjhYnP34E/DTXZheZeJfFP2oSJ/0dUmHhKWOFNuxZ
LUGnwRc9tNJ1TeU2nr9mFpR2GI9K0eIom2ZiWvYT9dRFLXJJWbrXSnQY3vEB1mXL
2LNLlom4QQeOn3KQkC+Hp3dCi8hdz7r9UC5AKyaeXTR+EdcSWwnFnoowEnmIWSsh
ltI80KrDKuQ6f6PQz3dM3PM26B9UrjowlnBNylTK2Eg63W+cqZTQZuvgWa727XbX
tOnCqTa/te8GTAWG6H2LxbNyqt7OMmiZoBtj6kfEmXVEiWp7prR8VZKQ7RnsuKLm
MYDVdGFLKDSls6W4IaxJoHZVN53KFcFox3NtKFhzNdSVacz9eg8FgvRtJP7QwUB+
QR3SZobmnSQHiwweKoh2EZfbWWsTbOI6wl7mZHZqMH3eQ4GB3dB8dsUrLlXXIirR
gd+SBgqeGnkNMJ01yt5sIFITePObaVoTUdAvCdjI1OCaS+EWvOMwoz5LCJQN8YX/
qZEUQbf3lNWROFdwY47uJlF2tCVWqF81aw+AAGKXY2hp5zalTt+hKoD81U3IAsXZ
6sOuhIDT6Cts45KJQXiZ2ubX74ZYibExmN81jgsoIOgHuYlnhrRZ4IHtu+U7EiC5
n/HMphuM5k9sxYQpLFZqVYiemDlENDOd/TS7EXf+/p4tvqtQ5lEIfpTjueHYYJNf
rEGdTNdZOYWF9rcZPX6zHYkUhQCtyo9+u2P9ueR4pbcqA1/6VqvDbQat+9Nqvsve
F5/fW0+ANy7JOD2RowkzPbcrG7EpLtydSLyOpOfYcE3RkxbUkF0Rl88d/h1NjsGA
3B/YkHPAXclCTlfmeS7UNVG651mzs1aoeFbjm1mVUYCjm+SuthOrvm4nrUE1sC3f
rY8VJQpbOTTq6FF3B0veOPKtiO4P1XFtwQTsb0EOaNf3UHpcUyd4VI+zyUqAIhAX
oaEYCTx42eEW0TewVXZobM0+K8gvFpVig2fN4soZzErxqXlngxLy+j8t/zTqmexm
jn4ir+hpeXsgLqPJ6t68NmqzB6uOX5uVA1l8vjmFb/82zgMxjMP7boXX8CaK2I8R
h/t52ISKayxjC8A6F7YPRV2JLr0V8mZ28Dfb3RF9rVnv2w9e2pdirGGllgOoeZMG
bXTbgMM8rGNiBSXAImBk8nWnMUr/jtiOvh+SpW/9hZn5U1nN+l+VrLJaWXWzCLsw
IZH9badUIeoU0l3/EmPDd5P2fUeIsweXOsO+C1IklZ0StbALM3XHg8KdigQRkV/t
eezOB3ewkM7jJUqY2BOnnmfPpnHwoUL9A85zt8y6q4WADys1JA9FfKhDx6vA6Gvy
2ZT8Ond6nPDkKBS0/HoDCIR1ZzGYd7+uIfbN7WuGcZpSnJjwd2f17vcjuE9e9OYb
tZ7pfd/SPentVfCIJwBvltyomBjHQ4ZOB41RrtksTmLOoGzggW4IW/wVK0uuSst+
Nd3hr8b4rBjwidQMij7pItjHiPN8kCTHjrzJiP8YvzqoOljt8BpxJUTalESPNmdQ
SW6tTU4TBzspM8WsKk1UIZAxeg2U1dqY4pjPW2RbbOnkz+6ITsNQsjUnajdGJioq
7TYBpMscQiQy93A9kgsu+HpAWDWCC6zNpFyAuKT7y24SzZhy/Ul8nRBuWBfAwMzm
FJ/J7BvKs+BBcEtVC1c4EbP5paVWPpyTk2LEbHpOfll+T5XahS8qcEBYXVU9gHo7
UHp+q7bcIOI+uGPgpgqKVBm2cTc7wG0mQCC516OhFdneB6uEgISWAM1YgTnwpWbP
rsQ7liXZONPqwE9kqh1lBBhN4aAjk98o/3nD/9UxsDG7zFyky7xOphCbri54FFhS
DSHJvaesLXG8Cuz9/x005tnlcehXDk45bYhVFOS0lgM1lh2AAuU8gr8TsV3zaije
Ua2ucNOpRcfXXKQ91gbNHkFe88TAKo5cuSKk6RTXYQyAW+aCWpg8FkBnYRtJ+vJY
IbRmcNRXcryG4LCiKRzMiY3vHKBHkpxE+VfigceV0+Lr91AoqDd0emeL5SFkw1fE
6rvGrbgHuykB/AfyTUh0CTMsNYdECV6iJ8Jbdakc2fmHKjbMILe+YsVsKKJ36l/I
iRj0VocPbObIVSUxUAKY1lWFJiLeobuyblEhS6DN5EVFZaiXX1fooplxIa9NXH64
/oYyFaEz2ELe3x8FRHQSYPFJnwRqw/7DjsOeu5SiKFnA7TUUa/MpqW/J+EXOCFOs
W1iIYr4zPaqARu1tUMLi4Ni7nSc4Q2kxQSnlk1BzY7am8SDHUifqW3g3EGKt14VJ
R667vFrGbCeRYVeBlhh/4h+Blb5KzTFJ3QpoY0dKyp+wklQD8wMpYAzmKVc4ssRu
dc1E4oUFN3mXzbPNZgIFakmz96NHP5gKXiRRTEKpDCDHxC1q39RzhBvoVdSsJrTA
ieboJcQeip8uZiOay/l62wgrJh7YgYTXkbnkSWYkwtxMzpFTPRloHq/cjTOrUYQp
YPPpkuzvqB1SjuyOOCGJqAz7lkCeRb/aGNffjvUPiehe/rjr66fdvBK0cV16MyXY
fNlSbevl9LHJlWPwMmwXcIT8NMnNX5I9XujZyzwY/lPc8f9W1AtlLvyslZ5mwo8c
lQTCbU5NdMUAOMJe8lIDN2x93K7Ol3M5k1vAhVdjmWyHKjqVLAKdfl92fIrUxvRN
J0jWWiqvxYMNV47hDlmgBP8+S3vzhTyiluPyGKA/qN0ZnP5CCQ6zACnPOML0lts9
R+rPXMKpAeq0oyBVLsO8WjhsYljUoDtadtSPo+nz0sV2Ze1tPuMq9G0/m27yL3wX
a0uzrzi/RwX/nJlQczrsccgGcj+HQg1qIh3ainVoNyATsg48UrBrYGLca2aNilTy
KghchxrI51T4iSjAgyqR1w0xcfY9TUAZRh41HqSFPvJi4X8vFnMz3KTdR2cVwAsK
E/CwWMIgoT9D9wUrP2JgCHRFsBuyluVEapphXvwSwMjnqQn07k9A65p5GgRUH1Wu
/tLP6lZ8r5seDDYjJVX/tdAr0X9EwSrRQxuzmtIaHd9XaSqtFT9J58T9OPq5bkOI
qF/nt009R1endAZJ6KVayhp3d/Y1fkipUs3Q3qlZXl/VLqLL0267c41fLxbt/AwZ
mIN0Eb6EMapgvHmcsmd7gVJXkJWge/x2kSxPUpHL6G7pllQWtBSlhh1wzzskV1uG
qZp3dL/PofwmSA2ybF0BinubPaFBENBd1Uy9i17j9etIm7BByEXU8EMoAURsAbcg
3TkW3O/eWtwtVDnsE/VjCwvUJUtKSVYDyYOMNNx2o7HLH8I4tFhz5Xv1e0/69GDH
mMhASY21fP9uDvEY/kTacpwgtmXn2kbGrmBqiFS5pRPuG1r1/LbHzOWaKiui7ow0
6e71blY5TaQDQ+Vu0+moeEnJ1VhelXENfFxsbdL8D6fESTwULWW15Y0xKw158Lqh
1fNQVBlhAp6x0PmZyR6tM5eY/uQOd1lKnU0CrQA+sNcTijgJIsNnt9bAkppWn7w6
5NDWAB0+/JqcuM1RieNxyMXeIJOTI11sAgWhfTbpk6SuHFDJ9o43t0Ty1Ep6u3Vh
VKGSaUWhG6wesbWJ07u2lBNnJ7ynedMy9fqDWSCRmylSZv8cybcGCZhAf4cuGn80
2trd9uIMhII0LuwMxBKHTvKEGVeo1kGg2X8HkHn47U37a6VkUnubJtoY7yhW0l8Z
MWPl5bTkl38o5oCRl7xtsYFw9uFisjlBz0hvswqhTWxSINGd71A8g4jjpFzp2Gs2
Ye8hx4nqexqLYpeIxYDRfnvCVdETGEHOdxv78/u0TpZzJC9deE9dgn1gICgEmGSx
HSlUHEQ3R0tlw/GAgI1zyD7gWyfROQJyRhMkli6UmWjHtLo+A0GoF5YQbT6SO2YF
n3Zb6i81CgLQwV7Uq1G7OTaEdap4hhsz/VslmQ8lKy56YA04hARxCcvaDQuPltB6
yMUxXbsrs8NaGhUtWHLlGNBU4mZAr1cpcUaZ4lwtEtwpvylhjdlscWFxY6J2/RxR
1A0MSqkOD8h9dzjFTQfJ3W7Tz87/vpOW5c1oXKtGSGw3yilAlyVWkj+irIk4Ht8D
NHHGnoMFxNwbMuErBaTbPPr0pp7/f+NRatfHxxFWMkZpK+yRWzFm3aryOUwcS4Z3
Y/vmiU++mwCZrotr6kakhBzCGajCkxv37JXTQN5zvO7gaJdHVn/BD2WmrwpPTvH2
Ne4qIS0dX/n974MSqMsBVdguvauIel+KmQ4EjV2paJLJ0pQ5NI+jrsiMPpbGq9Ej
MVuC4k2UlG83KmipxgJ06BnxYubtSgbFsDcOgR3tiZkzd6WIEAhRB3QZbtxAxXm4
oeS/GWyhXwLukSyRuR4pZ5e+dVyPmepLoE+8FqaCV/Tzn7nHS44yiIAK7EW9DQLT
9A+Kg0mvk8iMbQKJy9KvVuwSUlsak/6RONC9fECT4fei7/WMBbHOgZ/r2DbWPiw8
YZQe87kj5UdmUf7NlH/7YjxQmCqyEt7P+VX7cxUj+Ivq/skSqzw88JWOtE3uj2WH
DlhDOOWSi+qv3hamHtDNLa+AwyqWIf1tN2O/b5qHeZkzcuCJYNSYhQVctTelioaM
+LBr4kG9/cZ7+Vdx/ewZ7nPNJfNhUNitlGj7OjDrihcgDwshz7dRcVH2SN/iugkP
PSG399Bb7fwNDhxVRaPzvdIX7WhYJ7yTKrWuAIpobIwj3wiXLJoDcHI/XAU7sGEi
znKHwCFpAtnao2OC0mBWj4/E7PLt9hy3gdQmwhUf/2WQqrdiD57wAvca948W13D6
HhoSg+4y8tbWKjt34LHchN5aFUv8zQqS06A2yKpZg85YSAhpzl86ef6TecLZHH/k
QQFdjAvRlvPo/5G5FFbONI0ddjd/mXg7D4AErcDFYwwotiwOWXtYbWsyitTAmvdl
w/gKikautLZ3jGb2is2rdG7mZpZmGRqqdNVrpRF3TZ6vkk08tfPUA12Dt9Uer3dC
AePdWDHqq65kVldP4S0qx69Wl3eMK/qWy4HzBWZ8Ix2VSAuxr4ZkSFYJwavVoMUE
9wyN/lZffXgBq3a3IoS+HS4S9hgRGpKrHI4qsypsV5O5ufFDk8c61XjInq6ZU9OY
SvyMf0DuLWa0ALlfaH7yZcqY7ZjQ+jocPsacQfZZFNX4iiPSXI0JB3a7OWwY0tZa
r4ecYDuXXbUGaRZW7/EtcmT+ODnVSKBFHrygxk9HiwoKQjncVPeRu7GRTJbtUSZc
P9RZGHvjbj3ercYqcncFaL36llUnn6xFfH1vU2187BerXoJ1iIg0PTliVlfoX5en
ReKDXNan0fqcHVctLmgz4A1TlZNUjX/juDW/GQ228de4ObDyM04F+BSodwjaRCAa
T4F/a9Pp3c5nKmKlEko42khuDUqRrc/LtcfBdeKdvK7DADzHoDrQtxStVxiXqEpV
ssApDJvn201oE+ToyDEtNmUsl/8Z8tAzPvAXenqxjhs4ULBfMAqJNGS4GY+I5451
MTk8k6+aO0zjHI/x7NPuMY3I/4w/Z7vrDi5D5etA94KMMd6iEJYg0K9yYRyfoM7q
YbwPyiZNNjCyrdB6yWS8jPLvNhLq83RUJuSMSA+U+ZZbC6DMdE0zs3bm21dgHoRb
hTMDq4Le/EO6AxjUs39IjpEgbTlVGbH4HYpq2VoFCx8JsX9NEwVDD9xx6MoFhQLU
w7+EnLMYSTtQiQm7EV5RbL0YJvYfs3yxSXdP3Ni4eT1eiuK+fXT+v7WxsdpDiizi
/M+Xaecc6AA4g8zI+eSf8k4uYqrI/jLm6t7k+hlXwCIW0xX0VykIChkfznU+HIwQ
nyAhB6Ewl4Rr1LMBUu54hhbIaSnozNxQMfY3nnYsoQjCC70vLTZw3n+KStlUFgRK
ZqQdHkqKnwCiM2nZGAJQ77gtFYUeagdAdQO1sxXGqG4vmatc6TIb73q8EatT7sM4
a4FUPP3DtzfQBVksQsET4OUkN2g8mMeF4XB7CuoOtqtHlxp0pXmrQe3ciLvRqqOj
sS6ZT6i90hnKGQ+qfQ0WHPLCAXFjlCsHply6v2hwMhYCBMI9lmz4BNBchnMquEUd
MhzRuxy57I/Zj/GXH8sd/T2WoYTuWXPM1c/LL3M03Q/wg6Q08Tlqj67kOb8pThEm
d3DaCj2QUDka4HNxIhunDWp1jS4rZhy1sJTuabliYlReW9itzvT9C7/c9mGz0bI9
zXBLUYkmSoVE1abxgRLymp6Dp+fxOMW/HDfbXYBXM0aSWeDlmxQCVAusGUpm6yAe
ZaD8j+8aCpfKlkL+NK3LaMMb7i7JqWeCt1+rvwyBhf1HWc/R0JY0Fuffz2MxVtcd
Ny4Hw0TOY3uHlnBZAdznZPjeCJRl8526fhCM1cxcUQxiQmtHXRJfO3OiQFGqYNdO
ELboRuhpP69GIFvMtD+NsfToUFWGR52mCyyq4Q+TXgCtiAWkOwl+GBiTvbKVqgqk
ZlyPI0t522zk5Et04jKmSH8H1HYPPr49QvmT/EzJ5ex2MLlLfNAN8UeoOUtc+oM3
Eti7wGqQl/P9AUUsEIRE+yHJ+Myo6v3N4a9hcxmGGYZpy2iHZckZi9zh53n0TFGP
/8a6O3qNzyX+smfrU6N0lh48hCnydQaWJS+xhWQ3p92SAglkeSOMSWj3kPYhTkqx
YdMtzgGX0O4V4OdfM5omEWjx6d8wL/WFeJT9mT4sbexmBMsR0K8EBIj2HxnAsAIk
1Y/JekF9OYVVXRltk7Nzs1whyn+rmvVP1TbnISSTPlNyOYD2+BSi8c6K07OYAsgF
r8ScSFTX+ksMNg2TL2rNxEti5Y11JBXA4FBrJGR8fFAaiLQ5DL4jxWAiG2d1Vcmh
VRuyUEA+wze5nd/XTf3OG8Zzj9aAOJbtlY6zvei5Obz9eumBysQzq1ugu7qfC9ke
DxuW4qrimCrd2nKuSf1ahvLVWKGgN7D4LLAmPlxnqWkMkJ+FlyV/aQEmjncarg95
XTy53R51s+qe6WIma0c5WmwxiNVWIjhGDMNxkZ4P2cZjKRKsM0RPO1gZt+XH1R8t
EwslqnwlNvcVCz4UEGC/sZdKxQq+JQRZUQOSb4MnwzZxIsJoVIttA2FSV3D72J8X
NHAJtMd0UL+ulVi3VGmI+Vf1FC3hKrh7ESZdbRkS+OMthpPhQnMAsmnQU2aP+YyK
gVlXH1y4Jx4J9EDNo5EKTHU6shkBT2X8Ca05NcFXUWdDilmdSiSKf1e8eccBOVfk
nDSXOp2opv34v2vy+TIG8QXNP8R6br8Dvp3/kpA3kE0T69ep9AVhQRbJ1E6Ph5si
s1ZeuLIUo8yJRmgOEfY3dcQ73AZDEHtOoEf0sgjClhUFsu4cItqw7w52Z79EELfR
nzhQ17YvTKVwPu82Nym2L1hYpAWkiR3NDaQXoRzLmNJ4vhE9ex2t3hLHcDLPd6ke
S3lEZqxYAdc2+SXvcghDyET8TJzAhJvIhVf+QExofbw6GdiTxT67Iy79YqS/THyD
0nVdf/vl6y0RtwWTnA65MWdn5/rnlCc5PQ2MKADc+wqF8748jTvGAQemeGalua5Z
2NTTV68G2PGTaxd1Ms20kYpU3cchzlXBXxSUK5+SFJfz4vF7pKDi8JXyt0F2tEgB
vwUYhXsP6l3ZUD+VumJuP73irdvTD+mYnKUr7zLZnU3zBQZKtW/raLzEaXg2yl/P
PhuUtFH5WQWbsAUHi9BQRskoV0uvr4fMqHoPI4s0lF8RmckZy61ixs8oUnWsiZNC
l86AfYZriyotHr09Ykgxsm88B23Q9Ef/+i4yw5wpbKswfmAfItAU8JQU1np2ghRo
Wc0QSwy2eeT+G0C072PVQN0dQAD4H0LmlUaNHk5dHYujQxJZgv3Xt2PuX1rXwpCT
bZ3r6OaYtzeHhd/hZJ0/1Oy3b/YkWB9Mp4Bj75yq62H+xZUURtcGmW7d4KWs27Z2
XGCrJW8ZzQdJLSdnYZaJj5wLeTvyjdu5ScSczkuh0kYZrkqUIoJBrCYKx8N9Qkx7
HbkozPomxtVU6KF8FVsyy3ORafj0i7CP0XdFDFtifCm0XKKyMR8svvTPm6qcMqEO
E2UI78TaPeOZ79JclNXevOyoXpX2OigGI2SYWfVqwyIzs7T2Y1AfsqedPdJfiB/K
djb9Mn3nuz7PNCtF/KbrtK7c0ZGoUHsW1xlEtKfKDUuJ5D3JX+bt5Fhn7X1HuG9W
Pr52tPePLRm5k+tNBZax/RcU0MGsRCZM7KoSCxzDR46utIPRz5SnkpQX4eFkUdaO
M7p+QuOJSwSZD9MUnsUi/Rkuon7/Dx5JE0XwoIw1clTvAZN156zdZzxjZ5hd7/2/
lyCHP/r9WexVBK13yET83X4XOQjh5EQkRdI5+1LL8sjxPw9G2bKHPm0axIYDIoaK
6wXzA4FCPTBhzgUDHyTZ/WWHEmPLrr8+Kn6JkhIRwrOrCoSPy9i5X2BPxvfEGyNE
tE+zgo3k+5O7uIqqQGJQSm/6FeykdgjbMKGtddmWIPSSk0yMIQyQ85x2wQIV3otN
5EvVtdFugagdgGXvFzYUtvMfDRn5Lti1A6YRoJDeiQGBI5Ys70nb/vb2enpFhg/j
vGZ2853Sz4WI96K6/DCSRAz1Ci8sjHEDHTuXmQyDrH26Ws3Hh4XIPMLdaBayekm3
myfZu41Q/QBDcULL0GRTYMvvtsvtmXfbX2efT3TR8Zp449WqyHFcurVJoj4HvN2r
KjnJJXTiloIt47duFccCGGe0A77NhfNQLSUrPcqr+4vzCVtmjBDT6QU1wFDlNRim
ITfaCmbJeSVKs+3s8OnUeZSstTsmmzmKOmIPvo1ICF9UrFESzvyO0oairiCOJBpu
xhJJJxeQElo3pLAVE0coxh173FpsHHTQBKgmEXnhJSvn7zdphRDNNOCQ+M4vlKUE
TUj8d7yVF8wsoi4Furokmlm+e7bpo7fSs5e7gc7oBtqbnG4I8OQfemrXtKEsx4I9
a5yGxDBqkrjEcdC+uIxOBQodjSTDy5BT8t0YAc3r+mlsppziG5szrXcIUb/JZCUi
AYJEMAKY1C8NLTQ/LeH2FytB6WKchReMVi7BbUGqegSzbNXjYeSNyPO2BU1MX5jX
7WjT90tVw6eqq0Dwtlfhamr2l+Zy+Azyyn39l0GPqpAkJvDXDzPrQK3nqTs7qTEo
Mkqnb0dm3f6X78K66m4vkUlsfo53Qlq6+w3LexNZKL1G9W4txw4iV3FyLxFEGl3z
yLdeAlu9jXOiSboUEBol8BRjCszb3rMzjLfVXUH0OAezGE7DeCyfAHl10Ulb+oPK
Q2hh54d1k0xYHWI547i2mQlV5III/4WTyQc3/bDUlnACVTXsi6o/WaM0i17Hi5RQ
kY8atl5HjYo+douNAc4GgYKFiwlJu+rGS5jGHGCRxYkn18KtzvIhcfHOXRfOuC6C
6rRx1VqxhEXvuGucdradEoeUpzOELS7qFySjvMA0S55VJhfNiHrDYwlRJVYEHyGk
ERbdOppBxYceC0V3HgsGdiGfvBO+8Wgj/bPUmHS79Y1fsal1FVh8bpHXG1TNt2K4
nH/AXAUJbxwodONi06juFfHqXsY2Tl1U5TyGsUBc1CChDlZ2BR1eRcIFDTLeP5Lx
1eKBrv3TZYfrOWFWn0cD2PB1z5AcjqBy7uLuU23h5NdZya2VVc0/l7Fz8NlkL5Xl
xkwBjoGp5a3C9BNEbqkHxhhWeNhDFhcbhN4bW5gS2c0DAU6tV/3G15tK/HdE9JxL
nnMJYw5EwQx+SjJHAt2AU5CIJe8sHWVFyLMmR0GHgN9n/WSOP7RaQbw6nuOkIlke
/d6C2w3qrumidDQNN2Xp/onoxPih8c05W6u9gtkziGhv6QEWYR1VXSWADsJDF+k8
AaJuEtwYe2zVHuFEOFqIsWQwu9bOQwUJJ2b/mgoaw+AOrwIGypBltMBL6QaiaU2X
KDXI+m0JRNXQD03FdO6ViJp4Er7ib4ddUvhZy/AhYO+GwfCm8HPe44+UD3rXlwf7
kGBvhc2Uj2bkWqJBfUXojzQBEUvuMuVp9RU/s5QoYUkOYhW0IfpxpA6abR941tH6
oH//JGZ+qwZjsy9t0QYaNUiC04ohnkOW0EnbCGfKe7/EPaR8KMKWbs8TevqFlOW3
lPmc6JWDu2JVix5/C4IvEeQB3VxnDq2vpRVjDhK1kF7ZmPSstAjvLjadNRIczEg7
6AZZX1NA9t1b7Nl6yhcnLOxXKuwBoNlSxojPHl03qW64Qt9sOCtfl31psnt+FF5B
8tENyThJNnc8KKURSp7ZrYLiACeKXi43qOiQh2B/BN/qgPH84nu2YLcAzcpKX0Mz
guDKbIVcIdWm67rVdgR6GpxWmOQmF3QxFbKbwOtvO+ZGnlAiPkJskKcLNyiMmbMA
feZB1Iu75chTxdX5OxDz0KkoNOLB4ZQGOLsjXD/WFopm2sMUFNBMmyJ5SaxvLEcA
X38VQnHG0KlVjVIUPWISW/TIDbxv4FFxsRAGKkZdNLvQlnuDppy0eOxPmdyDnhVp
LAbrvNhkpUSHMpmul95JuGCMK3UI5pjrncwBlkvtl+295oGZ+QOP1ySrnsd8Y6He
MhbcOc4wuo1u9iFfmEIw9NRJxcAcGUzm09EJM0OMUoiYsqiHLObK0SMEvTdi03Mo
oE5L/3q6alK4STV/SMrRB0sSUknfEtF/nGwlzH32+am0/dMbim3nM1IqLjw0txS9
XegKZYPx+jMklbEHd4/wnI691i1RTfAkQ8BIYFWtQOu3gMnS5X1cHZkhN0PExstI
mI9X/Qts0Mu6MdJX9ad1th43iD6ZI6ptbd1HUN71Pz/t3dIj/SzwcQvAkXjaZRJY
jirOEHojKMagEyzYgyA55cbpRZgfO7xDkrnUYPRLdtctIHc6ic3MbSC/pN87NyeX
QJNodjnva0thZRjIdlN36/oszR/3QTV8bPOhC8/t0Prk44KdLgp9fb35dt0F+p89
69ubHTUDyYVYQNK99VICh7zLz+UYaFIM+9MQn4ZmDyQUTYMpuyc34ocuWqUikzt3
EcrlhKVSK+Yau8G+/HPK2Q3GzJTtzUV1+VOZwarRcZdhQIUF0KpMLWsZt3Pmy7B8
ZHgiQew6YiFUADa9+dz0pa4pqsrGH1UvHLAe+XIE40Cjxy1h44iJTHuqdXzhb+JV
mihrL5fMMynPlMRcp+BWdHBY/6M56ejIUqPNOC7/RbVNEiqJ6SaULXHkINiDEkK4
U+v+pPnYtSXNE4o/fjv5Wy39I416Dt1fO4pjt4Y4VZHJQxdI0ppZsl4M1pe5VqgB
+b55Aun37dIH4DEklg60YJIdNY83etqtERH0m1r30MAbHfWh3BbB4JEkUsSSgoP1
BbCBw30KTiky1Qvt+ETNs1f3ZIAE1Qw0a+TFR0FTJ09K2qIEiQTaKqwC3Ee+3Kq0
7QiWENUEpy9kdWqF8hUP4buXIEAIzRNmGA26Tsj2bZyOOrRs9yrOS12GaWPofXoc
X8afdlcpu4IVehTBZlp5sN5nvYk2m7dh0mlkAJU90nAjSi64s6FahcMArUXfZ9J1
R+DZfnYkKritmdkHkAVuFo5C28BjhVQIvvD8lsOGsmZwBQd4ViqekXykwkrHkpTY
pSZAyRVFSCOf5WFRd32JrNKBdO3IdCSjqZ24WzXfNIVsucyhBo8QZB5NyFb1WU7D
Kxm3LaMEj1+KBTKKaZcwz8oT+ILM/TLgfrbr+wI+sUaf74sM3Ib5SStCjICVZmn5
g9lYTzcGWxPmAfHHKW9etaUmbrln738mAJvgpRb6qmnInh+ghD6iQ3De1cxJsFoU
5I2dioMCsKY1XdyOQIGasrD5ioQIoOTZvpGlMEi7PELBtzdjlN99JGPs87qMpsN9
7lAUVG4BW7z5PJThlxIu2pNK136x58ISKg15fQyMJwywIyZoLh+czkxNz3CGxGDy
F0QdaGbjUtj62vTL03Om+kih7SXF5MTdXtLDLqznHOOdYLeF593e5uLuQvPt2Suo
flyw8E5biqAzZvgPKh2nv480CH/RsFp4UYz3aYt+X7kNWsxX5m42Ut5eZj4sPeVw
7YnEY8aBkgqL+tz6aJYs4GBjwpRuz32S82miq3hShAL0DLaa2yW6f92CW0xoiGJ4
ZTWKQ70nwQoo2r8+DP+sCIb7AaaoUCoC6+TUbwH/VQ0n1Y3iXK2yuzy752U5DO7m
QGXvlZX2u8okX0UXq4ivx7AlSdX3G43GaC+keb37XP8edokAdIuJ7C6gKF2AMzDN
LNV4k+9Th9smOvOZYGlQZXQQCAz254Nfa87Jqn0CfEgqPYKUCz6dILLiHu9KmTKU
Ol2ojAcD9r95eAKoN5n2q6RCuhRcn+FxyKlt0/2uml+69CrZUI+dcAhaL/XPNyFF
/OWjHpdX3emVszuAbja4GODj8GOFO9Aw3DYP/gLX5p/Ti5LjrLILV9rtLgW+pYgW
NZw+vCXr+ehXUWuPjgODaeivscYuAThZ7Km1i+EF53oG8Fvhf/aupHMj83Fa2cfA
kSqpJPXAXA/lzmZDi3pkODkd8ZZLun3t7CnGoy07DaB/UN9X1e5AvRJI8XeON4lL
WhWgO4mUKC6jxMYjBjvlOnUwjua+iFjvZeBk1hUFUFKUGo6jH4t03zrZHckzoBNo
2DAAIZ7Pa44ZEfEiS4RoxZxxnQSeI6OkeRYinI0zoGdbSULZmXpjEDGro+79LVFS
Yq+YYUzcMnc1vAIV7DN8Iyypeo41yp5FvMn/wMXyu6Iyjqg/GuWo1zn4tlm/vA3a
cv9OExDNPw+9Q1ca3knNx6GPvbJfrwhfEJycL/fZ58NUspMq3mXPZDv43FjzrodY
e+NymNfqWvhzaMukoH471QPapnL6GmaFNs58IhILBC4KuiCNu8uJL363lntP6RpE
G4glMBiJncMIIVxAAwMB28XOE3TR1ffIQos8XbLRD3y6PxT82ItbVwJ0khXCVddJ
tmeDV+YmqA3MiK2TJ1uLQbr86zaxTt8vMegAOiMQ+pxhogiiRHsOUFqx8ag0RmBU
y5NsIiDOaNmZVvgwiZvQGA+QHz6pTsj/1WmF58vev/fSr6qVtgMXghY1mnZ/EfNa
29ALrHMrM4Tf/iagU4VYPS9TNFRBBDcvFRs75qFzI/cyD1BefqOpJ0tdXtONjX3P
UL63m0CbAUfRSa0Geg7TuIdO9WrlPDYJudQsQI9Zx1ZJe1sNasYQurxdjUQKhfrt
f5TXRgPC9I0vYEaoT4cuUcYlMLjGsR1gA+zYR9nxJHJakvkxW2syz6Ds3iMy8MnX
AfzHlneGoNnlOmejerjgZNgL2qxYs9iLHZjc1OehXxhPcW2eu91Vr3a7/no6WiCI
jlytbcWBPGYh5yvlaReB/+172LdJfFNxpVQNWZek3V7eDSXbbb3i2eZPh4bEm0oU
QNMZHVNsrBXqkKSmfa5PYxf3itxA2rbLYW30DVPXJd1Kq6cFHPbUUAurEzBgqc+U
7QGFo29Ld4w2vAgYST3PoTKY5CNmNLAbAeMPzMnrMJEx4BJoC2oymkue/ze4/ThX
4k0I+aO6A586CSL9uBUzuUalbFpGtzx4jGGH9wuVlHWDulvxeziuMBVVfFAKpFUw
L1wwlCBP2W7/FggKMhwtnxgEG+elb5FCk1nlmwlBJhjI1CJigC6ybv/obDTO11eJ
TI4dg/PQwSo0KtOq9gRfCCIti1AHyznjGzj+97pOYBwzrbtm92N5cxaDpx6dzojv
Hn0vPXBONzoYG9foTYDG1t/xdQwvLXrNuMdEZ2HAmQrrSmI+mrU1v15++53UoBxB
5hxAhyxSmRhw5i1M8LyO5AnQ6YTrHAWhwBBkGYzDHpMJk8l34hwaocETS7IfmVjX
uXUCiCshAbqfWeB2WmeqRf/BmR323YgcSXgjkJi2nGpiW5skZq/pDu+GflFanvyf
L/cBafn+sC2lgeLU/QhrKJbZoweX33BSoClu6tKi8cIe9gebMG0PX0S2Uv0F/vlR
X/Vrg1RV5AA0ok27mY9Rv4tAR2++dfXjfqzxgjNLf+iDT7rwEfcVrqB8rfI1Qbue
CW8lAfcmBAzDeU7/3n3zl7sLOHpNBAgL07NjCms0wokL4aU+hNRdZmQWFqZiwlqL
PxiVe1Vny1FwACQJnw0X87kuqUf+Y2G8d89aXu1GXF0qCyPGBY2zn9W5DM/1hZ3Q
HykCMmH7K6WpjpghVmznggcWbAAPvijky8OYs5ZNDW8rnVL56WGowkUhxQHKoBpm
4RwC9ZT6xtzgjrckIIbe2E8z8n476/3WfXBG20qSf3sEb0ZK97enRmiwzp9WFinY
360zz+R7M5d4DSrOzhr14fzwPakcfrBRNJIiYHT+tznb+ETHYWDjg3CVVy1ltsac
PoIwkezkiQPEhl+UKgRXNxJeSCWNI6S9fQECg0wGQnKNVTuevOfHxLwFxm1tkFLc
9zpbsIYofL7fUZgtt4mJOBK3nHX/bf5pAT/2UhSDE3wocUi9MuFgC8YSSI+VOiwM
b7PCEEXyt86U/Vl+S1oy4YtE+9syR1s2C4oEQXrViJMt0OdgkhyG4LQY8A1gA7B6
KIysXrl4H6XYy7AoPpV8AzbzlyuhXb1PoPgnHufDNGDA+/G/fl02DN9qNnVX2pck
Fjm+NjK2MwQC3FSoZE2cCnQTjo4Hlu743MSnQlIzuLGim0kl31d5Yh+NCcUNaXio
UFgEu3670vEX3ugRPv9cM3UJ+CVBV6SqTiiw5UAxw7zITfXGbRlYOmPV9jOZbgKC
u11jtjCDLMh3XPdYvM4WjYCkNlFO9/TB6XE7Ur6Ts0PQWryDeiM0tmcPUxxMAg6t
b93mURCjr+jhcnE5YkGmV9okZMRjx8GevrH+s9EdTBpdoNWveePJ2gdlT1moxNfn
u9niwW436Odyt/uLK1q2ipNCwnS5KvawpfQ5YD5mYjk0AoGwIph2UlSPW4hfcMZW
C54yQrZ32wbXDtr0vGEbybtT4qC1jD6Yn5gkrk0gJ6L4gv1wv7eSzE1+hYKvB/4n
KDvacslInztsBHgkDY2qo6pXoyhMy4M5LgAd/pyZgaOun5cCr1m90AwcDJRBmu96
FO7Tofocqad4JLlB6Ir0n3xa1JEhqcdlqDZHFLpg6W2uwygWtYUd0JPR5qgZC3Dg
RB0kESaS8qQXtYfPJ8EhWfrp+BYWEL+lpWI/DtDVDkqIByD9/9qk5Y4INGkkwJpr
14xzqu3u2QkWsga/gnbIAcZ2pbVU+1JusN4GudwEQjo3FzJ5IivhDijxdwJBeL8A
YTE3kV+iCh7Mxi39AJ1ZoMu5A/TdHiBJGBlM5AbKwI2EbxTxR6UmQJOkB8dzDABN
xWrdITXHhBOKQ+QrE/XsINL93eb1ZaW1EW56J+2b6mJbrcOb013t+jiFABQ7kJQO
nWan33BMDX8TE5iYJRmdAFxb7XgiFw7pIyJJTE2IYPH7mGYJDTKkSk8RJ4mqDB/T
kGZLYf/mEBc29BeyCirghD8DjqkBkAbCmQD8O+2YMUG19/IGI6p9t2GgEQfnrIkH
eNrfMAw+L0QyFNwArgv9bCamz/O8PqQu1Ha1ClGrJ3GopvQk6GafdKfhUjpK1K99
xvEGDib99y9YDb1DxiX56yIDDT1TcFUc0hikeQA+wAbRUXEXylXBHGw+H5jElJCy
jcUWOYCDWIS4rzS4IEISRZ3K85lv7xvTzmVo3/7DXGEoPpbwV/cBMW8EftxctOPM
FoI3BcAT0d/pQ2xVNOG53GPn+TAvoUocd9pwnxV7Tx/Nr9SZI3l6KCs5lAG09UHW
a6kOQdZ9hhaaSdhqltyCinC+ovTYrx8JZdIg0bEWeSVLhsnZVkSdeN1rT+NeU/XQ
EjG/usR9gYzJ2REOK7SPkdomUq9VtW/h852bXx2BDIuWe3g/ekUp08sJIqyjATui
p/55xzhHs9CgJpRbBoN0pdtJMxebfu0WaNqYSKsQq3mGmMkUBuP/wulJ1/nRthsz
7UdBQ0G7re6sbmZQhCsUTltlPCGnHKkuw0/1oHI2NbbOdgKSGZPIqHwXmW/A8UjV
tvi0aOXRpsJg5wtrcEZMYCMo7RoAmMtvDzGB4gbFLLRypYCY7zSgc+TTlr1U9R1S
dIShfRaT7HmQKvPMdgg3bamXbixR3jS4aL4EqMLTwxhq6cODrUeKB2+bat3CgkC5
04xu31kpEl0IInaLeWIxxl81fFAHZN87ODOQvS1Cnz+uuHxHvTmROEBe+IPaBlSb
nxIXeTwvHVQcSYaod0qajHaMsvfN3l964XtaM3oQmkN8+hoo2jZ9mozx4qEuBjHe
f+Fzw1xB5xsGh/LaPhieeiuuH0dcVQqykKFfoy+aaFv37nnos7g/5SlJf8Ps+c4R
KCQSfwYkUaYW0L+clU1vX3P7eUc+SyqFjPe05+tMe0JdpGg9/tqrXH9I2y492vAz
1VMqeeF+llm9DCYu2d3CSMoUJ8WAXU4GJeD9SF7erKMlc/q57g8GHsaANw/hdjRR
xt1aHYKFWyw8ytzbyed0wZJk2ZjZ9rkjGmnl+jAC4U0w/fd7vD5S3uFFvz5AZSVR
9jT/f/Wns/79haVqKAzJEPzy3FIT95iIrgev1LhCGovVUKO9zAL488FsvYFy0jcQ
a91yaaAVaDZ0/BJaI6lkxPFeNY0d77nZ5IUc+r7llSZxVP4wntWrA77Y9ejvHEMr
/ALNwYlrYquS+F/Y3uHS4Fx0ubkZ5UfFgY76T2E3RiJ2xfLOO5XhNk7z6rmVREQY
oUKJj2aavhvvz76CARfuisN5bHjJIaxiWXuIUuveP0w1Z2C47twxVaoybBr07Zg2
MBHHm9TGeZ1/ynApWQQD/H7/LQRgPwvP99PDQpAme9bGsB+jTX0FUbfRvTkii0M8
4/+WkWcBXpFsgdGkEBNu9tVe0462m7iJcugtA0a5bLuKp+BqfoxSztq69N43XOd0
NDcpZl2uCXOW+jxQCDgucC39sxYTKm9Fi5kxI5aoGVM5eHaMNL/dKhQzdXAow93h
1fzY1q0STDL1iR+Knv/HjYXNA8pZFMM+V6oP0M1zLF0w9KMxhzvrLifmJYqZLv4H
YlZDJXp0EylMnlK1v2KSDxPnMg/LgOR7DBaPaVfNgX5MWaSBy3+4NSguO9kMpb8M
kC/6ja/hwlG4UDUR7EaZzhsl6JRXybC7VetDP5cOROQRmW/+GotwSvCwWlufZN8b
zC+rDbDw9XGNDeP/5I8aa+R89o8ZEropy5TREHrA/yPeVs2/Bs56FsjN/EA+pS/3
18/gEuuVpG9POyVX9q5Ecj+4bdUvjpIchf2Ujebn0IdospOKHqNevI+r+q/hvegS
lOYUQL7Wmci3IQc3zdPva8/K6+SYuqWFV4o7vmrWi1qWAAhb+t++Pj9QyHUNH8ut
1Z0SwmVfvGU/3shYYN0XRMDmwSDAxiP17oBo0kzF8dxYXmmfh1U0eV+9j2AP8MSJ
JV16cWlnFtZJu1sOuPF3kOYA5Ox3NSeui2iUxexLSUdw/iXxraEWwoDERbRh1aGn
HiOKCAkPi4uyUtCisqjRp+KiBJIxc9HaKhsjmnHNtea1IuUyobw9ldAN5auFWN8q
VwmkIBXfukdkNi/SlBxpiW1jitHVDb2aFbJimSVdqRLj/xBRLrFMvv89U5B/aVYg
8KqrP1yeK19JLy74366JD88z7ZGVoEa3phBTZXOCYN4MBpauvJUkWoUs+vUvWMsW
og5i9crcu7dXGIzK987s6sgyjdiz0/l5+qyZyfbO24hXwBShVxB6LaA5690+Snzm
HxyGbVPlv0OTdRylVRUdbCh/+IrhFlIePkb4lbg1G1SacZ1sGaHCNOhlf0CcPq/k
t9VuvQL0j2LD616vtHXuPsPcc6EI3iuyXspMOBpdDyf6R1BTqMSFKm7Yyby5+ga2
I4FKqugGwaoVCqr6HILBTFvOkDpWNIb3enpC2fcGXAgunhFi9jPaM18posto5n3E
a8lK91pCOUXvo10kwC9pxunjuPMQbxIudNfA7Tcnh+F/kKKS68QI7MKrfUjutKFl
PUJlm/7lf5ZudZfwJPbturQwDPWqq1TKKVuxH2f7FrjczRSWd0dEra7Wo2P45cMl
Cm1uq2k5eJXDFdSdEYrrEEFwIRh3la7H7/+ZM4MLDCF4V+4ite8h0JUAnxWNDz3H
3tWtlxfVVVTpR0Ngs/yYU0sMKkuSQQPhQta4U+Un+Boa9r7amDRE3hCTjHH0oe0X
55DckoQCVY9hW7AiCmulZK0T0ajQp79JivwDgYs81oLtVOwT+IwiIgLL5Mybjpcm
FyM+saPXctBlEVf4B0o0dm9gYV4qTt+k7qBquwrt2jnkvKAwSQ5qzBCIWtQpQg3K
V7zbm7c2zz32SzlUCGO9Hl2UkAdVNhBk2OYJO+AKIBeMaC6b6cG7chSc+BotKRj7
bs362uG4BJJCR+8F6QWLVZ3/Q2U2CQFEuYFK6zFy56CrMX2mzpi76fuIRJTms6V6
L5H9EyyM5PYZb0RyPs7lPPEcQqznkbLiSrFjl+KxeA20f0/KQXVrmbVB0P7fjl82
J64h3MJYyL7kmTrVMfNUAl7ZsR8apPZSK41/+p8+JtP5nbW4SB3ihudt+n9gtKMQ
ua/7jt4CNDYtEoOCfFcatux3VDaRHu0CuPy8woEOtijSZAGBanlkQCNzX2WMCod/
UiD+FUOJye7MIOYYxKU0Rbz/WQ9xn6WmPKsKpQq29EbQiWtHkhClgHM6IbHPvf3w
RdvZ+vchXNANaMIVT/D4Oh1XrV/EyI58CWbazAmUmWjSsYtLPhpKCEj9lY6E2KGK
YIrKHV4h0yDb1AzL/P3DA7dYBahz2fCwv887MIq3xWtwfzWU7Ip0ouMWOrg7olqT
fechhH4bU8KWBZllfSNX3amqeo1rQ8e/p19P9H8xaJKRPAglKo/nnWqvanv392Ib
J53XOmxuGKKiiFKsD4H7rBea+fFclVclGdIvRFchgQFOYP+j5lOFOU6ksiqoFrdj
AYlKZa1rDmrqV4A+z1ZX0QLvke3T3SUnJxcXhqGVNSjnzxlpSgfl1aOFX8P24SDi
xbG3g9Cz1JUg8m+jJQfzr+IrSiV+0AvSxaW9U7O3yLrK8s07XVsIbIteqNyqUDfo
Z698Tc871H8uokkR+TkkA0CXYY6by99MSFn6MBIAR3YeSq+gE3H9nWWVKA0o2n6L
HxUR5cvKsp9TVL+npP/Y3gPiwyo12ltX7JlToYNtGpppmGuT8C1+XW7+aIUR9WkC
WJzAblhZ8X+FMhdc3LydyDsB/hiy/NDMADewVPF8cFqx58OqSw2Y4DBOkSBJ/q0z
FZUZU8Ah5yTZqNJgiRYws+fMF1B+97sS0+BOmnjt3YUzjg7feP7aDP87pCG2/les
W2SvHJ9sAWwwLMlXTxYrOuVpLDcievRSLUwnJ0ZDV01aV4BTN8s9VFdq6Ko3WY3n
6eXD8a/9x3pAxa7MSCaYAIIRDP/pbIZsKRGfG1DAFR42OFDfAA+1L+YvfPttvwae
QpL4hmDl5x5dIWPouB+XPkuwJgg6UfwVLEbEKJNn9Qd3dIHh78RXYvqjfcGvvP0c
CUWAE+VkVu6gzC762xSf1EA+hgmd9DYZpujUeeo/CTH/S7KtzPtH6wap0w4WsAeQ
S0jsS4Y2KQAKWmE6SbQ4fXxTnfDNWwEbWOrgstK8OAthut25NV8DFAmmOSlgooox
kybT7Vtbuj3gG8ULwsHZySPmA1whK7WrUU2XGV6lcp1Wh+ZW+SCshfl+Xa/we0ry
433q6alK/AZ+pha5XGN3Fv9FZYko6CjqWg+fPycCESRm7oZvJOiLah0Vf73QYZyd
22oK93irdd/PvsNEchrvmhee9scvMGm2f3rn/yBr5xbFiegSMSGL+V58wu1Vq7Vd
vCXi0oV6ObHIA0SzmhtdvuV/rU3YaZTRzXnzPl9MQpbIkHX9oEPmdietW789DNsX
Ufx2ASNs2uvMy94h7iNPBugbSYvWZWZYSj1+JuSkoehwi2wLcq1mLnW1/I/LvSVv
mIL2Ly4KO+WaPomkp20UzeYknOR63/barZUtoTpt4mv9yIHw4DM2ixRZfuF1mP1e
N+5Nl2xMGIESSXmqPIiHN4QSrexG7jLufT4tzW9JBXZLb+wN/LhWxF4NBJiz03Ui
0I4s2Nfi4Dz6FJ8Vsl+1Jti8Cl9KmAKTUIeoc9NVVcJH9nueg0vGeIG4TBw7rx9z
mDdqjl6yaYceRjuvxaXIeglcnWU5I8W6dTNMft+AG9shfKXxDl2+10wgCEy2I2G1
+486dxAjtwa00uPACHqFOKbKOm3Di+Id7HmCaq8rkV6zMKYFS+gESZ/FyM9mqqqF
Pveuy/2jwIJyU9AaF70jbgH/ouF+AEdkz0Ob9FuhmK5MGAa0GS0m689hsJPnTUCk
XSk6R12VuKSIQws9+Cwz+IQdddWsYFe2/QMdtSQrGiWn9V2AE1PyJJNBiRrjeHZx
bwt88X50JwcaIqv6kSpkYSQpw020Nk1/jbCraNLolDMSLT+V/PyoefYetQsb6dXn
8vK1YHMwW6r4HsyZonVbrjRZBj6TA1yvOu6x5sBGNaFVc7MfCrgtmJH87CEau5g5
/hH5RmkPRDLHwtdN1JemUt7ML8BQJtsaaVFV3zCGLRVwnU5cASy/jue2g6csJm5H
sqN2I3QIZCeMKFp63h5aPVGVfZmACzD9eMVb+/b2w9cU+DjyEMhQQW6VZAXn7KR9
1jvx8RgrmkZz/HC8WA78MiNOwGEBca+fQDv+zWSPe3gimHA1cVaMMxo7bRjTz59P
YXbpQpVUeiaq2G+FMp4FljDnd1+xzfNddaSUI4tQ2uxnzkB5X3n/iR/+p3cNPIiI
rXcv+dT1IPPowSpCsPl/oEufvzTJ8RVEbLbS7ZA3cPjB8FxeVOgLbaPfs6JBq3i1
wNZqtcS5E8ds0Cj21gyCL/AVwWN/W0SZolKc3HQHkN5119HOVXuP13Mr5WQRIUhr
YXzDT9ua9reiJlXIKUTHHSPjPIjl76DWPpV5XJfd+x1o81r12dE9LyY+3OuUhlKZ
fB/Dm7/uPWzVUoL/5dzOShqi4VdZil1jwrfcqAo53vmPwcISNkyS0+trbfk7Zf90
xncF3x5UrwnRZjRIubptX8yXd5j0IHl6s3r+S1c6v7t1Xk2HEuYyK5IrSuugGRzE
yuHfGbDZO9r6U4QpKdWOQ8yuDjD4PKWTJhSyfRMFTBZWZbR5cqjsHn1I3Cnm78Qf
FZeAhfvzwh93O0sP6cAFo+v/OIlbUUcb6jSxsb3dkCn4lnQoDV60ki5X5EIdEdF6
QP3ayzyM+pf9u0xNcGGzLRf6gfRbU0HwS0QvVOHJC5BphK2IeTUoCMZGEYfyHfyH
L3AQaOBvEFlzUWeZYxCPX1GYWclIMcKuyrFjOmzS4YkmVb+0zLLbhN6KaBAGq9o0
Qg8/RbIXOVROBLk3FaWRr1g7niy9kCmJ6fA+DWcx7F+ycdpqXPdaJ1um275m0ew2
1odJVy48kcJ5gRhIMKmS8J5abYTcVOHiu5foizywKS/wtKTUm6LIWS8Ff5vTdFHz
9jBNvs0G7drPQzBefVwDzXaoFKcCz4TYYzNpdDAWw8qsJHx2517OjYA/MbhnLj5z
PDhsoyI/sJ8wucJdcjE9Iw5Yg03vi4LAPgi30zWDE5jYK/lRt5+06fLolU99D+ds
KVNgdfPuvT4f/DxqWjh4ZDL1sPGj3T4EYUsg25st8nO+Eqqtdx52rVziwTV27viR
a6vTp3szIe0fwkcVrbPsx7I/pr9urc2x0Aj+7GFWV8zYcH5OjzSVtEY4AzmuhxMk
FWCEl7E66qIYMd5E46XhBdJBhpHi7vMMjzqdnGFKsZCRZ0seLEzj8lafLV58vbjX
IuUvfamnfDohWaV/2aEixE4DNJtfiehcj0MUB/85nOUPIdmiAMakk6ra65BwSFDD
nOUAqK7nZTy3Dmwbeb4iSpRAYKrZl7AxKwhWWpixm3lkipRxl2pMUPDv/4/CbSvf
3upv2KmzK3/iqKgDETqvJLgOqdJAFWb+yylqEGkcpzQa6Xjmu3yND9gwpz0szIDZ
XdlUbBiCinPgSjHXDirkjYhmnV15kppiF1YvItKRhWif91dV7OSXU9ZAFhvTeeMW
3wktnRTxUoB+/A0N8g59H2yH2ju4qofBxBp5HNXNYgQg550PG3nOfdOmgmKvThIf
SgjuyLMy7dlbCE+z+dfOiC53j9V0Qi8nkzbRZ+q2SP70klpGPBZ271KoSScfpz7M
7WUyrWNkWTHbR9EXbK44hmZPFwUuB5XgjfLqQGLKu+KSzawk8DbgQCMGjW7ai/oE
6GBtgpnhtN2vQuWXoy6JV1re2l9BZlO1SICGtwpvsjXrm5pAqoL1jRa37U/Smb0g
Q27mTq+JO0thHvu0h6+q72I7cUugQJn7CB5C4ctjj/0saYvCVeZ1jRjfg4kUrnO6
u8Ypz2NDuNmnW5dMBJrdBwC9t8qs8LIKDFGpfbjtW/xK9rshWUH9CdNh+8b932VG
fTEN7ZL9rWhC6SrD/PIH1Zs4zHwQEED8no7uw37DEctfRMXbj1whayH2uBeKaARY
hcBbG0zBhoa/Yl19zfsBOZVdT7EALONUYwzn2oeW9rjc1YEogfo3XRfIRgVZTvFh
FSMBA0ew7pVxI5I4e+6gFxybx3ymnOQjSFbkvBUzX2QsxmNuDz3vjKzwYR++kTzS
gaFgFSYb1ZToB6U6QopJMLwQwoKssdzsrgAF4jtq1mY/rcgDRHm/FEUgFi25VR4z
fIS5hRIp4+bno0A1b/MfpH1cTEBN0M6Mce/zTA8Z7OzQq3BXUd9pnVKh9i2I1hmM
kFzM5u0y7NntdmEFx4kvF2FKymDf0bddGbCQ+yMH5rEtZsahze5yvGOzNWmxs1Te
Y8IY/Q+hXZBVzbHzSnKQ/QnmR1z+f1T+/WIhvIwzxN2thf9zJ4NzirmdBlB3/iqG
po+YhhxR7/5JX1MgxpFS8H8RKh17mdY0WZ2z6Stl7ZnnkJKW99QG6XH3VyZ4EwdX
zxjqgwkN087fHeYQ+0xUbNite37jC+3uL1xcRAcODR8oe0Sh7tVQFvF84efn4glv
NBrmzEYHc7EzhaGBi0dJBshSPYtwLjuSfUzY/gQl71eDYD1BYww/g1jrUNcIILPj
MaGzpn4adpxF5kA3AofGtD/sKWhzCKjayq4Ms1nV+0AThsFwPRM8tDMJWKW+/jLP
j27bY1Ah0AQWFbhA9/ZUUScvMxn5VS13cD9mrtjLHzsaGTgZ1hLx5Bo8weklHmut
yISiXyI8jZE7yx4zxlasHqo+M01mUG6KK2F9ozkg1V8UccKU7/+YkXcXxjL4w202
WakZA9XZCI/++hTLKyBjh8CwdZ5wgq+H6P3aaBp7LOIuT5payiWBLgNyLjJJTklR
WsALYolEGAmCdT65e1OwtLzUr5MUE8fbxX78wgUVc6d9qivwoOLYv8LCG8rn3Cee
sKs9p3GXS6+NSayd7rKfVnbepO73PVIMA11Yry9rWkstcwIERzsILstukLCAATVO
vlTrYx5Ngc0k/ZRFTmbIewxgRFKXXOC/85NMc+fOe0m01OlEo+v4LkgEzoGk/+ey
IwbagCyTRQNKwE4xEuoAmqOfVuXu2YWVzuNnXUbrDaM0emCcK+O7+75cHkg8wMVD
Oym7KgYX4Yd+rYBogHuKXUe/C6EYTXBCLhcb2Zrck6mwkzHDQoXEhoQFnm8tIxOH
rp2SeHd6hz/NQ06bU+iidW+uaniptfwSIc/zJtZ3h0goIPYWRrXXclKUn5k/0dNh
NL/lJwi84cbgUjtFcO6XqzWsE3qQZq8ICPthvy7MvuHXnUN5FCtAnUMz3Y15Abn+
sqsD5+jBgjg2J+4ZxAG6oUyF3hn/mRB2/BWzSPGTmGpniKum05tSpml4V1HE7PBh
IknMFF1A3dNXbqcLlgZpnIPAPhDFMIlDSqLowNlYyvlt8kG6/LQ3HC6qpLvFOAWI
6AlrG6usX8oeQ0b5ySnB75bIJx7c9QljKq4YXYqG/QqslazOzzHZEvpGSaKfKToh
IsNsUNRQEwk0SQQWRXR8vNLkGhDcOR73WD14M7f5PRxf81B5cE3/XUKWk3KPjZcB
AiccRCRRnUEwztFHxHF+t8WOhXtAgE2QuGGDeY7Jw6u/UYTDtOOAkNgH6Lu3XP27
ekDz+ClMY0PPBvy4nwL3qd8kP91zeX0i05BXpMqslfNvvIMvNfmqEFA+fhS9X0Ic
nxY0OjTBfQSP0JWd3D66gMav/MnBIIvQSbq+GRyGlTIhlqfh0dw5d5Zm7Vbdebsg
f0Pjq0cZGvFzoKBNyy52qeB+2xUDoUeQQwSTM5m1+smmwdCEjUHbnEjiSqVa1Nev
KEaTn9VwmfAfCNg1uEVz67b5PlDsPv58EWQe/V0ecyJDuVTA3lgJxNVVkx8ltgRm
609odl3SfTGmRNz2IXwPtNFu4cs1B9e24LlrqaHJQsDaik2FJWEFaFyGvCwHe18q
43WHz7b++8L4yu/ycPAq5h6D3CJstRXna1ZtBK4U/vUHBugbh6fVlilNRP0t6x/k
Tly/roTCvYzxgmj7A2TcYSn445A1Xf/wh4lhF6//S6z8UqK5O5+N4VgizwYmhYE2
8JWe2NT4+vFitRcM9Cf62xqiLfoLppaFTfoaFt8EJjy5GZrlo0tGZHs/9XhesxU+
te4b3KuceyDZocoiKvWw4StmOAqzmoFQhDRu0RRw0AB/i0tAscZnAXjMur36b570
Duez4QEXkk0W10iCeM8P//CQdpawVOod5HWSloqlNAoUCmwyd4aBkIwVvt9b7sIP
VCmETenIaVx7bADYZfiisO36tcP7IN+j6NItCkjg3NnQpsuaIogr5y1U645iiGlW
6bqYcDDUcBUmYZRYVaSCkuolHG7byizxjZebpzsHaFV/ogJk/33Vc0WW1ladXv9u
q53nynKZuQGvOAIcl4TnwG1RRttj3X73iBSONN9yACZeOtj7e31sw7V0Qt9F2+ke
Paa3NYSb9oR8vBnRTWtUmxHiiE1Mdkeqw7IfMdtDjKiHZ98G3BfnYn9wwfHImZW/
xua87NRE3/mPbEF56UUTKH5bI7RtLAeKyFDjbqJpHFXCbPPP6EU0j/XI+5Hyl/Ba
/nrHf0dX1KR+JeK7nh/TPZez/7T2T+dB4JTZY2a5cFkFgpJxbHL9WHbNr3MLMczF
tMETl03PU87lRT7l2NPUcYPpmTNO6UbuJ9cB8LFWweiohbMZc4R6DLFD3SOdWwjk
ZpdsnVTdl1Y04t3fP7ucQSTZ+PQt/6jCpJ7to8qne84KSgpgBBGfWhj3ERgi5KUJ
fCOwBpvetDVrVwjxT9ODW2KKu5zl2GIX6O4dB6dHU6UIoE5Y1B1aiRw3lZE9Zn14
qYT52EcuDHjidLk3JnAD32LiDOw8NjnxvKscMGHGFFPDBf4dKCeuDkccRKULkHix
BEcGJ+YgCmgVckKOnycKefzdGmAdhe0lvJJcbPIdDQoPErxOFm7kMtCDVXSK/YXR
YRd4viDLaebhVyvz0ofeZ4VphR+HfIz9OdZ+iWB9iErCVs8IoveO+9pi/bnoWf1V
NeywEWpFh0V2rBWV73NJOu8BJptCD21B0aNUGl/kCUZl/lSOr86gp8YTF8/vbo8Y
NykXxOgtGta1HMlNTbJ9hEVwvHR3Jso+lj3RDpnwJy72LQNN9rCe/YM+I/8W4ltM
4fEgJADVHMvwJiNgZ3feiF+4s0w3fWvTLbJXKA8SwVWaRdBoD5B+oJOJEON279Ty
I1BuUYNejNcQ7Fxaz2BTNk+52qvSzPeCt8kbetd8By9Z0eaLa9KgX4onMJfHG+hD
VuNSlaT4FWoTyOgQKXDG/oXG+xLOu1A7zU4Igcjp82GIdTHMNTdetMSvvrK7p6y4
3p93pXMDspxfSudKgQ1/oqOwJWw6FMbjDXP6g7LfDgcws/bDGFGRSqDNGlmqSAfq
sW1JoPC0/NjEC8TiyeANMZSnnNq+6ci7a9Tb/E8RHIenFsNZPAa3jpndCGiz2ljl
8GcSM60YcuFq/yc8mcHoKvrSKaWnR/rs597LSKFK73uGuekWw1BKERckzxKTWB8b
fngbt5rHb2GzgESmFPTYe3CsyGElD4m0Z5CSUhjRN6qh9BUBJBK7awXELlFRRpQU
C4JmspGSPw+2RJ/85ckJ6frDckaooZ7rfQ8d/u8PMKD3VqrakKx+K4uskGzFOcEI
m4r/EsoORFkoWjxMEubS4yFWM8jvMMjc9bDfXdiTPKaA5sQCANGvS2m2XEWqxMW8
DMeBSLwCMrXbb7wIzxiCxtHTRMmhHbJRRpbbj4vHjJK97GkXWKmVKL4tHGd7WrF1
mzgr4pjmrje5JoZMtQOM6TNYfu/uz8EqRkNvbTYdjBn2TZ/z7LckrXezDe7C3siJ
Yk3KW2/xAzATkviRdQxZcusKsUbxZkG4A8tKyQxeNpC7AoIyoIShRqex9B3NgJkC
IppBi1qLZ+qNzjybzBg3jeRg6OfpvQ619yDAm1pDrS7KvqKTS6SuyyNI0I15cigE
lihX1necjJpscW9W5VunUMDhROf2jNB7lA0Zfw6sfdckzd5n2j56zTGMrycLGT5d
8J+D6S9ceAPDvhBS4a0GaqsVIhRYsMzBDp2ZfYA7wTiNG5z7/SDzaAxBIinqWhPf
GkFPZ8/EmQb0gxdYXYHqlEAKYCG9Ojbym/01PtNjDqO8DWwv9GvK1r3Ym36icxdK
XulT+Oud4iPJve6gYm3eiySO5gb2wpRnVj3H1zAAmSfkmgUZeWF7jFsQB9c9c1A5
+a/X0h8SvzqIYbvj0oIH8aYNc5OPsFdMpgA4ATNy9oOS70MaFVdr/QDn7fTeQ0Ui
OirUGbE4yRRRmDKgUCwuul6EsRDS5ReJS9bx03D4If/O3wSa2C5hZuank9LtT4WW
KyIDeAgJyJrfT1tAUL506g==
`protect END_PROTECTED
