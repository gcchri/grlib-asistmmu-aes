`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
feVuTzv0EDqurhhQfQaZqS/ww4Vsy8zfXHano+QTlldVbq6QwuxktW7E3KF0/l9J
ImohSDuXzIJlSZ0KKNzPdhNheVZn31GXnozR9jdutJFHTXyRiq58N5tHqfA0AdMI
J3VFY26/KdrCqwMzWyh9ErAVyBbSrOYhAfd8MGMzdP3uNladjk7YeRj3rGyXCRGf
31qdg5n4nVVk6lzx3k04ymzmMNK1/oUB+eDgsitzdrvDBN6AO2fq6j6UYesL4EYP
Ng1h4iu0lDSd24kvXLTW535cmNrqs9oSpn4INFvQoo6NTaabr3JiQUUvgt/C1ifw
WTKFbIf1QRtnAIFe3sxJwQf1+ofez9XBlDcg91caKdxyTn7kExqkErAiCd4J/W2Z
mBThj8zQggbIkt8kKMTGMA==
`protect END_PROTECTED
