`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XE3djDXMdK8ScdqLHYEWOVnz9EpIJ+DvnDsjOAvtEAY93QvxI0mN5NnbOUA0s/eS
GTqgEVwAUjne20qD3mPCgZO/YW/sIgEl5Z5ELOr0wP40338uh/NrEv/UWsVW27tK
xq7w3BpuOSpvgjgvHRQrNuAFaALD/105rW5Dy4+JmZkCiSJwVgRS0cKhazlaN8Sr
MLyor+dJ3byg/htHfOKskGCffLu3TeZaDhy3TkbMcY+xdkz2BUd5gmaxG4mVgf89
9MVzS7LI94urLCFJSFLAEqTP1ek3b/2gek/StDAq8954iS05M9NHFdUhcjqlgO01
hACfkL9I2Q8qJc6yKu9pL58q3mO9uy1+YjGoTR6k4u27BwPefmqH1LFfS0wrM5sV
VugINTIB5wuRQf7dV1mZnkVEMl5Ip5WB88wb7i0nfyAHCNb7c4a6t5YTt3fpNvbN
UTZ3jWboKSRlmA4FUuPo5EPu9CPyMyiUR9GHX1pMthse8K4QS647HNQQlLw/+TTV
NYPtVRmLbrjOy9jMbIM22XC8P2/9ToFV1WgzT5qpWjU1dQyY32DxLo/qTP122qOB
hoFc8ZFtM7L9tQKfy1SEEmApeQyCZn+mwSLV2gqG6JlwK680Wb2N1A5+sPu2xSCc
5njHuqNLRh+zEBXg4yBq3c+ozttGVq7OreU+0nYSWSAI8+viO1Eo4ZddqtnNSbb+
XiDc8/MFPv1/Qz3ziuWZ+YBRjsNSv1kjMnCxkTMhiyY=
`protect END_PROTECTED
