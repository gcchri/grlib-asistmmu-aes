`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXgHqI+oovvT+Dw6d4VzFkslwf8aqsRkiLBxAZlLGobrgjz1fOdR790m9/trT28Y
9x0bfiINMEgtGcWGNkHxd4Bd7b4nxZLAuGl2XnEdm0/TwXXDUu6ZeqtzoF3vHGSo
LLbLVvivUtqiH19KmuFTgodySFnM7Ixez6nFNWTTUZ0T70ozkxUQJApLZtKVkZiz
kLDrhutvdmdj/vOAg4i8CdcXF+Kg62N0k8mrf7CuFXQXGUHue6zLX7zaFbICuAGq
NFCUwsknUrRCAyeuUtRPIsB6V1nCiwuV03n5nSnab0DS0JCXsonap9MDokGbi/ga
trfwjsCctblg7/k/JUGzWO9CCQMZeKEz4i9JgdYX7h+lLzCQZKFRIa1U1kEpqslS
2/WcOkKI5KYsTcsSNxemHJPmoAJzGQFTaFJL7BYu0eL8YpA4kETH7Dk2pPH2XMV4
RbgLkP1ZLivXXKpi7SIQk0Sm8zSchXk9cFU5RkEGh1r1PBdqWRW5HAYJRmG9/8mA
mZViIq6AwGQq2ajaTinJXM+VaNG9MjofnWlUshBBpPaYP+aRwxloq+aXpzWlrmXa
j1LMJiD4OwnK2/AKxwX//BhuYZp+MhQ4QM/D/X8SgAkrPBW8NrIBqR/B025T6PBy
3wBt4jz/TjiS+iBWPL4wTRmE4yoItWL9hZqyiiYWhdelSGoVBu+wnvx/GW5aSKy+
7izrt8UJYEZLZXPDbZYUafn3aORurJq2tGcOg5Dj66x/DCFFryCGmm4igJKlJJ5V
8Aw1SQyYDhmIudhA2o81+GCw+ZLJR57REIZvXF7UcIjojnAnDzNFU0vdgGoR7kBu
ShjR/FI7mpcuzFHbIRlauw==
`protect END_PROTECTED
