`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jT792YWKndZb2CJoFMhE13825jwpCnKzzzzMW0naviYqkQRvsJgeMpp+RnR8g+d/
H7ATgrYoavxIkJABHcnal1N2PCWfddEOCzuGlTxjA35AfmlBlRoNqY6jCRoJ1jXU
MSU/JBR1CkK1es3CtJ++kewRX4TZjuLOrqg0BPkZvqAo1XQXDwwSNryF6qmNToDj
f8gCy79hY7u3aBu76atmWNVx9AQGRRvkCgRs+Yq3fHAYh0AOnTTgYV5ZakQXR0r6
HVBEfexqUZix/fc4EEobtuKmzPvkbbShdGEhUpGNkJoGJ1V2QUoyfPYN7Gzasjw3
sQkmmE+LP380wWJ9xAiuvX/cxQvXGn369DOaajHS8Tx5JeFrV5JoRn7r3eeztMHV
FrGYMAAQSf+7H6cXJESNCZVr3iqXk+6u2s4R53kMU+eJk8mloeYVJHPxmMK1U3rJ
x2EkLIvYAmnzmiPkRFh4EjX4FheDrtvLksoKz9n6EKQ=
`protect END_PROTECTED
