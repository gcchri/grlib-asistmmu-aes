`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMGL6QHStoS/s72B91Suhw7d2NW84XLJjnzOlZxNxYRIn0/8j11RooO+MBtHJ58j
mF3JgChgaV8chqhyD/RDQ7HTs8fSi4Xiuo7zEtOGu1nBv4d6hKxdZ/2PNabXXAAp
YSi5ismHMTcOIr8cFVfyx1wPaoYiyxWVbe17c24e2SQ/vUw34owdwXGhmf1ZUu/2
dERywd9akBqxffJvcXYFgpyRbDokoGX4JH7GAHUgjrfOhAypK0aiu09GsEht+Axi
j8IoNZtlaHzE92VR6C+R+7fzPAS0H/dUNwrW1oNOVp9kA8d1HVH16oswEq+OUZqh
roFl9fdqK6n7lwsUuAeeGKxHsVIYyvLkHwGQmeyKn/EZ6MeQWnRT0FIi6Gk76WZ+
vt7EX+Ly5pB69Cu89mI1BfrHDKz4HqsyHkSRpVDkeXrUcKyn/PS2lDJOWmqHNbom
qR+kYa52HpPSfDS89YsDPRytUGYFxZElVnoY7vUMNWz/tQ1qcXk90Fg7F9SCC9JK
Tvj08fGCfD2VYOou4V+rda2f56fmnFqe7KkGbnWo+sxRUM+037VP0Hn1xLlm017w
0ELDzXKLOHqEqvGg8r2HBQ==
`protect END_PROTECTED
