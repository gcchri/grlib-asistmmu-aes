`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oP5/FgjrIVorNI5DcqPulD70GgmHp6ayYHu/J31YZuoWm5kPqxsuYmpV2IZ4zoBf
hBQhGjePI5cZTbclGjurdv5xmc03iBPVb+ltnaDut8HCc/7BW0VABj6+1WVy8YK7
ghSG5pSqgacGItpsr1G93kOGOg4m5QOGGuPqRD0TzfK9Klm9V4rijmi7gm39ucXd
JA1bQ7dhPM8BEy9anlkjKyLJI3GLPeIh4W1i5ryjJMNqhNZ2sU9gozinZU7/2E0G
8+e+gTjcqkVSes3UoIRLTIMVKxmfJaSisYTs71rs5AYue7u8aFw3B/vYbV0FykGZ
52q/lA8WiNZX5qcr85I4uoXRpVoQQ9w805la9ZZGHm6bRRTlzZK8MuXXc4OzcpFO
CE4ebNV7wqYrbmxPQZ08jUJtybko2NjM7kiIu4h0wYpQqikmoz1H0djWwrcuWBRP
gn+ylo7gMjgPRf7lA3rSzkPvFV8ByEIb+SSM0bO0iOYUr/crUxZBBhM2UiNLO7jz
kATD1dnMwLDwEGq96RayS5Sr7WhSfDLPRoHxiMaB1UvW7SDMbOyZf83xgNlYf4pF
gPn2ZPZtVLkBva6SSiHt7RdAP2EQ/xaml1/U84jJOG3Bn8k1AqagxoqyRxQU9jZc
WVO571hc5EYwN261QFCU0B8jUOLUFciAbWv0hiythv2yS0bj2oEVD+SKBG5oGi39
6TkGnFME95VqX3V4PWWPTeGCO5TLziehKy2LtT6CGEkuobUxGZJpR3ucNKUU/Jwc
9DIqKqvNCQb7+UCsCuho6boZi2tbswLJ61yMiiX9ISRigFc2xftV6MdsFLyXVKs0
zC9TpuDnBn9UcBVmiMUiKR0/67mhpzU3Rsa0GNojo2/enCQbRD1hFh/i/EmEH4kr
b5p5Hs7ShitPp11po8/JzuVFU0Xu96SQHxCP/mGCD/l1789daIroajru2rn0tziu
S542TwL2oAaXQGja2J+QNOOY+FZx15xWID3163BYRHfPNE7DftyISF+W0rHIDJRT
A3prOS0PR8i1mq6INgUoHXBBq+SyWhtBOZ6+bE/gbP5XRqJWrcABJ4yWwNMkaG2G
FgZCduA9qdnDnHDad4B/OgHQDxb/lp9jIuOFkNYPC1asdhAoS1M9lHmPQuXrD6vG
It6Rfe+zimKiGeBecfoBqFzmobAn6zXPDwo/456jPig+BbHcUkYJ3dRxeLB8U64u
tAZtxlglIUNc9XTjTxTHaA==
`protect END_PROTECTED
