`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lvm0e1DQMyxGalW298j5YJe9cIrebZiPMKQuHXW6Ue6A9Rjp8oLAsC3PQYRimwLc
Xme0O8rHyWQZP3pgBeIEwLqGq6PKRCGZilYKgW6WFTlXmMc5k+qWWFr3dXYrtgL/
lCb4YgE37P6BE/pNn0unIUXTVCbMZ0/gJ0QZVmubVrB4Icn6gaQ/V/77dmlELZfL
WQW9u9eV/JsDcCUNZa3GzWQVtGgYSmS8wHoewS5cLpw61md4vf5t5fHeO4GCZSxH
wkBBZQvHeGlDIFqeKaCZ8v4Tr1ZENaDvOAk7aajX/zg=
`protect END_PROTECTED
