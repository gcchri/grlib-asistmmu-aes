`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RACuKzX8bkFklkehneMk/wQq4K254ihGGv9528lMxMevAIZ5V91XPqVv1nBF18aN
nZFc5S3BECxa1IYhuKhtjS4kQiOUJFPrh0CM+oZYY5sEOZZ0gPI3yzRBDMzKXSlv
VpUm5mtgwOhXEDX1YQV57OPUkAY8XlKOhVO1qnrWMf72lwwvI5DFoPzWmyeea98y
gwR5IHVxshqtNHAf3TnaTvXvC3y0vEdQwlmxPWt3O0MS2RTBoYvmD+ffADpGzXAc
ukyvDQnIhtHh2IPofk0PGF5sLu5Jise875oXzxsWz1V+aiZ5YZn4Tlb5prTTWRt/
hth4QQpVOAK3NdkbpRHU7zSDia7PWyBdQn3c90gYqzMAbVSJeXebwKTO3VlKjlsc
B+M5HJCkJiOHC9CqPLzfGTwLvejc9aOCSS+Ik4IkQBqwnrLgmDi3iEQs+NNBJ73U
yPMwCO/t9OR2yPj+nwyom69w5ZqmlsL+iUIQloWKBSjajzIXBvv4MmSKAyf7Pvb+
w258JcgjgFWMPFXODLLtte2/hHVRhrY4ZIphGoIsuNtkx1aEvibv0xWcZnC/MRsw
4lWtC7ghPDsY0B1g8wbMxvQASMpOKbr2zvAgzGqQMuvCzuMsQPAYK0ZEs5sKynwu
KPH7aexYZPmhEDK3x8gv4zPm46TgA2xxPhpszB4CDlpA6npXfqCIxVtDnqFd16ah
Xiee8WR37pyMz5ODSBlw6ORhS/VHp4DqnNa3EMjXpzU=
`protect END_PROTECTED
