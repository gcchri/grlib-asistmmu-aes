`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Z1JGnvyVxyFi9EOj4H/FP1/8COOzxIRxDVNw0Xirmct0sBVWO26b+QDLPrSK7vU
ewtJp4xuK4r3fng/7iRsLmlmrGxsNr2RuYp5YO2quoJlMOfhZUkMqUqibTRCXSmj
yEh7+pMG1hBRBRRUItQNMbXm2LFXccu8orV9OYwjTf2Si/1+s+tvRCIKrMbNxwW7
Sqk1Zma8MVN+tKqptRhfm+1qLPNXytek8ouDupGRlX8oGAsrQmeQOpGabPjigpeP
eygwtvvFSvIIYjBachCxtt9TmVFAXAkl3Q/hzMvZGqHb6QeDODue28t38RSetPn0
WbV2ERHvuh4zQ0Wlrd0K459FqMqba/L7OwmQTMoiBG7UvIbhAegvgeL3IycFk5WL
JNs3iF4aZLp8yMF7AX9V53soku4VjfkEuWkSnKYomYTS/ZXvhBg3CAHV3U7azt3p
O2FPbnM+Ks6BdezRGEhR1tdyYT05vOrJ6fx7VGBa7QtnI0+6VoN5uU/BqOncBFDD
9x1R64TKzAbwJPqnkOU+9huIwHdmsdl0USF6lASbxWl+ff0Td64dNVnvbrcyvp3Y
A0LtA8fb4zW5Td1pu1i6HGJUBxlWw8sxJJ5CMCSfaMuygceVCKbjuD5Ds8m4kpDd
71w6Cmi8nFhR46gBBum9Sw==
`protect END_PROTECTED
