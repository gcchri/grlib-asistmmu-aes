`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nKu2Kvp/uCVJGCbSslrZ8vrYkDgVbgkG4T3cJESrBPCJrxZEdY79R1DvdAIhddmF
w+sQ9nJjcXqNoksfekk+6mVCu+6W36atZWMenxCfEyHcSQ2o8rydTyru06VK1Vzz
8ZlQ9nI88udRUL13B2+jm2E+N3X7kv9GqnXw873jqg5umRk5vomGVnRPX2+hD4D0
MuxnVj+a3oVhcxyo3Cbd4XszGTzmBSzuNEwcL8s7mdgLcdNoZlGGdXAfZwhkMjTs
IfkL7WYWyw0QS44aaIEjUmqU7E0vs6tQI2JBZWEMs7/qP4H6BEwcsxuUn0xqDScn
VnrCiPQTEA6IMeXJvF0q8Taqne7g+F/FJ8ZKFBePVaLLB2b+sn4pCgdhtIBzzPjV
ZDwFjrYn3RzzVgOD7FFVxFmdrTXkChp9ahUelNlWnRO6Uqn1kIxfIFW5HFvYfgib
DmoPfW0X+Xp0TMFUn2lTYzDg3ga1h4dwfzEMcJ55Mmkck36gdpgBQklToslQ1QS9
LRkncpjcS1IsJb6MdPoBym9okrlmSR3lCGEEVfb3l1p8nfkLs7MV3EKyg2Ffg+7m
gk3wBpWujJ0jWAI6kj146vgW74xanKrRGWuMPRHW0faeZ+cO/N0yodqf58H7dHBA
lA2p0aAQ5PQ6GlgmSXj85OAH9m0V+3oQlpQuLb3kXT6iCJe8QxrOqJdNZcURz4b4
CFRprf6w/OXUpUycO35V5y2N++tMUGKLvdQE3x/YFspRPWbcWwPk5iV3CCfbUbeX
2gZJepF8EQkDccDrOvBuUjXSZorH8yBb5O79WzvLuD0QLTuOFyXJFJ+o5YeVZn7Z
bu6OjexDeTiXHVMdh0RoGJcZHsaI/hzGhX2X/WW+kUikUl1JUOjo1YH05dpPqZIG
2FA2yzPc8vfrQv4fokMTWQ58KmFTFi8NQghqNIJFNcu1qr4H0Q+joKcb7PMAdPHI
`protect END_PROTECTED
