`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fsXBoO/jVbxQ/NgcRLUCjtw7ccaqNW+iue31/Y9lghK9eoJnpi8y9OD+af3lzG5s
iSH9Car8sNvJ2LZGOGjiswIKBzG3WYeb9/ROeT9ahgAomGaZ5cXTF/v4CnHtJLhl
OQdkP8/hpFYeW5CQeKZtfr6I0NN9AefILDJbO4ReOxcmdP4FNLnhgck0SlHSN1vz
yj0iDYFo91Hv7dXc+AeAQuTBJK1RjJBexqKQWyrJVuWNKtaX7oXGwWNopuYA4tzF
eMGnEOSh7LWZcXUFMlAfccTxHVzpwRpO/eFBQGMTZFAGQEOfGmswnc/H/yRsBmaB
WMF5dfZu6iqF4N9EsL1axZ1s/Gz6/Q8C3g2JrWLLwnz6vvTQAl6TIAuR+osC8Hgv
NNPaCrIpPrIL4sYlfWl0lrfLZUuTo1NoEvw0jvDyX2jGpDh0XIEGLrtkSUcV4gpI
oa62EmB0c9Ypnq342olrJ0VoUQbBpABcm+nvBLktySj5ZnagMgDCVEM8U+IC1TbP
WmhaACUAvdbHeViaM9mHSghFmP/xHw84si4Y++97/u2XybZuWmeQxXqdS/Ony4O7
R7N+v8XIsEQZ7Gksj9UqVA==
`protect END_PROTECTED
