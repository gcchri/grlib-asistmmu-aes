`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXpFrvbRd6MITVc68S5crmoe6C7SSrZLwQS46WsSXWFaXFs4rT5s/fZACHprPU/t
KvARUoEor74hg5P0JGUPCNNV0eNrHjHiIgwQhMsyphsIRkBqChTSeW+0MWv2DHPS
ndjX/17t9cY6jmxUquKqOjDstQzqS9nhKW+aFFPOcXLcxPiuJOAkCHp+lzBqQjMW
cutafTfE7cEV9MPMklt9TGpaYC3vRobL0Ha/5iu/gHBfNZt7f4FZ8ms0dSKKGIet
yZKE8OokAhl1FO/pARCu+/PWGc+mvYT556sQ5s1u6flU8lbR6qQDctGunegOb7LW
IuM5n6rw51J29LEtEVfreNwCkyjwG2QOFD0b/zlzxPf2sFfoga/0QVllgBlBao/p
VC1VRuNlNSZD6IW6/E4Tg0qaQOdBuaGo5U1LfIWEMWlnaT4+ACZlqpTjVrt2fYCy
gIIHmHj8Zsls33nhM8+fXppLn70c5T8J1AhFMXHNuGCYoxCD+VXOLmfbqZriYISA
gZEZV7sN6woglmpxv1XYyUNp2mFq9+Tx2C/a3kwfOTVmTvOIgyELJFG7OxaY58jT
E5xq0q7PMuIGu67kFkziDkrJXz6qA2ONAtmyZmlg0nKSL3P/Viz1W0/sLDt2PPpp
2ZvaoHFXzbWvp5exgCYUAv2jQtsM0C3GsNxsmVtFXc25h4fjxiVjKsqQKz0Ikr+B
tixJMhNZfH6kdy5WuG8a4Ujww5R57NZUd7hPPiI4cTtOssB7K7GiWAs2czo/6i0Z
P2PckenyLAjs8cAI9YE/vUrewjpR2Lk1YS82WfdMX0oxLn2jVKgenr/IPIjp3rvb
2Z1Bxt6uirnphjCA2QK0gta2mLVUxHcKVH433oUX2Ctzg134WpT/mj3JW4K/pVFM
Dq2UM9DK3G5vV9IDwxghNrmKYmuaQDXGckcqsMbykuZiEDnp1+uIxphutlXyM1pB
x58hjw6R+pAwF84CQfXXvUpXtmyJwu0/Qp8C45yZ5Nopm4FfGlQC6+8CSajHCpca
tQaCQI+SSG8QAGX0mL9aQeybK05R1PW8RIWDb1TH5/D/DaD30KNfNTobrR3Fszve
uDzb9R28dai94bScnJz4w/7hZ+qR1HNTqn/4QJ+NN/De6sTwLYF3HfzXencqDlxm
`protect END_PROTECTED
