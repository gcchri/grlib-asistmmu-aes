`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjiT/LnkSBPTADoEIIe18vas4URgilTv75FCWLBYflWYBnoo0mMK/853FSO2q8mr
I3rSROh9YaPlrKeb4tRkdEtgstBQRFgRsCbzjIsoQ18TLxUhIHCFDifq0njeqiQY
plmwSGPqVCeT4Qs/DbL8D6phX++HQPxDLmxAsJ52QpFzhu5o3jYwPy4GorFuJbWc
AnoH39OXYGOUJvyihhbV/AMkSFqx7X+5SQXXVpoMuaHZ9lstOLmw7EizNM28bAxQ
td1Pk8vgvSECNdE89MCf4+yWqZr5uo9dWqwe0iCJOh8XW8zzLLGetU5WYEaUMC9N
QtdfKKSycQFTnYlvImJCXuRP6kIbrMBD/oFWR5i9nvO64sbUIiwtaBDQNtSKu18P
Oimic6xKDAxSZBCehIgPB6u8nID7+GyiNDz1b6oMEPn6H1LqAeguiwSRZLSOhcNm
qmfipG5Ct0eq/VIiVl5+pbGgYjalmqCqQMhD8noLQNtnwDQlDaIXUMYz9WDEshWg
tSlUVmnsNGaIii8E+CbxDQZSwolvz7Xp+rpwYpYGtoYGI2MPCj8p7DVJtdaaJOpR
Hk2zufBVCjqjV/PHQW4ODXmJbKjrrOuZ5I04KSwA9WlpIpafJCTdC9USc5KtLW6R
qFjikcXvE2+1SXH8vkWZRYmRi4hesU58pd89bjMrboPPHemCChecycOkpTMTyMvi
drRsZh9vdCyrYz5LLHhwPoP7Df/EGCu23FDF5hK+tTgZjE7ZjvFweMVAJdNnWwfq
csP+Nx/moHz1fokp2+7dDh13GqmuDRzR6sYs0ACbVNf8gxy/Pju/LYKSDsgEHMyP
q1R7pBKw2C/uKa17xxM/apGc1Uful93RCudMod6vStfNyOeA+9DVYaH5F1zAO+M5
6cZ5e9n1JG9qDbpioZm/O5rOHIwwnybbYfsI2p+QUVTlQ9m47Yk0LGKtqjL63SBO
Nm0ipvxBZ2KvKO83ttr9UtWBecg+c6UKPXZoHU9EhjsOkG3ptZ3c7YFIH9sst7Lm
oLcFtjCqkdiCIGUkQg4hJIPwnA/Bn7ZPw1Hq1hvmNC5CbeLXQQoDQXraswNDEXEn
TQVFkAlxwYo9NYh3OX1cxblXN+hMoGRYoqQxKSVuYWRrKSRkfKr4W+4OdgjBVmAy
kZRUyL/bmyBC2cPSxN+xZpAd8mJjLg8B7s14e1GhIxJcyT+RL+qg4hSoCA45EQb9
bXkJSdLqsLl+yNs4yHh0ub8SmwjiY8WbmW8H0aimATregGoqE7HVD6poxzuTZSBi
XjM5ADA/VddAVoicQnqMU3T38cf8r6xeOYxy91WqZn9o1TPLiZEV4rPBx/aFD120
Z/OjmLw3DWRA4OKnp0j+nKsTh4E3T/xWkCJS9nXPfFetiJd+xkZ1U9WZFpy+JzSX
gLOTaIY45zTkf/kTZ8zrSeVvfH5ppWQDUKnxrmxW12XtfzYmUP5sVC6rR5BfxxO6
/RPFXXdbJU8YezcOj/cLD6Ku0iTqWt1Tenr5foztDgpw+dvUOLK8e5+iqGOxDgJO
86gl5SDx2ZfwUGt++WWqvPgWCzuGCj5HPSqLfDSrCYZk3YvBqQTbuek6mbUCpZKh
aUgj3Mp4a2boqDoB2TVeZm4JXvnIzqA3RzuTJNszsXqFyJSAyFnRqOze+rD91t6q
gQ+exHcNBC1slsEbybNSjssYXtGKlPMUkvUWij7dS34SmDOj/8egNKC9mtFMyx5A
LVncxISfoiYOjUv7H8Ernxb6YZbml2iWoZlp6mCuak6+4H24LfvQLnI7EqIfyA9J
IueHDyOSN19dmiduLF3ODb+xo06YNnaM66uuwocgpBowsDknmHW8ICeZvBgXOY0c
oRWQZoGzeLWXI6h6qCZ1n1RQROisRyjOITKher9V5D4LQJGiqqMp+8QsLAvDdVdy
Voaw6mPL8KhcWixoh/xMNRDcDKPbq3R+CAKuyRXm+B/IC9sEWjr0tE80fEmARPho
BW5DW0g20sy+UbFZ1CoH91auurT9xfvESllCSVMjhJu0vUuJhF6/49yCLtG3X5ny
mhWgINKDNSxkUqIsnnTRWNY+652IRPfpNsk7hAS7i/umoEkPN0NUdlWQndzCS5mk
2yGTPf5ugS7Zk7a64Ur+yH+tKwQGIA0LEhTrByOFUI4fPT1E8f5kloU+8YRHuJrS
oeUdJwB3jiWR+DdU9h+e3kHC+fMb3o6YpnbNczRj91lt8T/Z3kuVwSI8mnWrbw5o
jFEuRPWEzycwN7j/mEvXF6tqgshtL4ENJBOvtLKIO+cOkIlo+ulW31nTa7JFzckd
NZKzVbFu2xzhDPYFy4KUwaAh1zQZwKOQu+0hLEL2d4j3fijBcQA1k3bctySclczE
Ox8zDsWNIdLCAvZ9aD3KDh5M3L6pfNdtBK0ICU75BegAfLIKfAeIKotT56HVeEg7
SRkIthojJwoRnj83h5QBYkTSKbCkGHvKRyMRT2Jhqd6qKwF9PRTVege+U9OKVg2H
P8bREWO+82zSwmGn3u5h9g1nvBbGasReX876w5vH9gpimUECP6ijBJh0wtshMwYY
g+o7LYp9scd4/EUTrCt2r5Syt8qtAWLAj6D8xu3aB4WHKJASRq5CMuRtZjTCjQPr
GhDmH1AZWDChIrRthLRhtjWLuWus7dlq2tSQ/Ni5bhJiNohvLu+qtwrG2Va/d0MI
SvoS8WsVZxfnY9h2sYBs3m9KaxC0+eHRlxGJP4lgHmfHF3R3hdeYhRJeyG5Binxh
nlH4/HqIDY4dKbJh4/KWk4Ughmod42ZQyUbaz4MyRov9rBfvF8JX94F/T8Smeqb2
oT8pQAl/10lIS32Uwcuzqha8jNbRtVB/iXBXeA1OPLTwHpgCUkYI4mYEZ2Bmk2ut
XfzJbK2/k78wkrfO4kWqx0Vk/Md8Bb1yLP+EqUKDMu/iBBPmBD0f1m1DDr8KkCQc
Eo6YNjBpkSCxCVGHGcty0YQ7t6IUhT6wOyquO5o0h1+Bo3qZyAfJKcP9OTE3+DsH
oxccWSDb/svxksOmcbSvJpbuU75UdQj3guh6PmXsrsXPW5HNssMABjrOdVPC5MSB
M0wDNASs15tFgqFAhj3IUkZHgIDJtnnuXW4ZKW6dEs/OKLK9CC/2uUaCiG4GHKvh
jcN4PaTARsne44VIbRHd1eQHBLGt/idfDb8/eG1r2UKgYw96YPc5MRpYY4USx9uS
1QdPcXWOBKjuAh+UzJHoNcY/1kQ2oxMi9Zc9Rt2POGRvis+O2Ie83dYrXMjYaQlu
xtwUbFIHWzlP4po8XR6DsTZp9ThrMlGu+ovnW/vYSiHPYXhH8gtnDhXn/wQl6RTQ
bafsP2m8RaSZEqgFCCduOvMdkVtdCh+pJS0Jg+Re+IshdvLyY8ARvuTj/+M2/0QW
`protect END_PROTECTED
