`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zJIc//1gf74crTzooGb6vnQcD+g2VgVv6927r1RNNhhQtTvNEhZ+c0CVZuRoq74
uTpXxqQ28GSOBU2vzCKGH7JKf6fk6JtLzVOOB4ezPdzbinwciEfGj4gFTGLWFRif
vCLuCPToCgFSnxkpbOkLHrWWz3oenIIwy5e1nQfotPVUtFJk0RuyiSapoMdujAC8
QWtb+VJwd9sKXi9RFL5XNb9rW5wUfWOYSahasRhXglR1/1bhJvjcYc/l4pYJMBtq
HkrS7ABPClNzf+qA7pseK7WxF9w4wvSFHMMYKXm1Vhr2gHmFzwX41SY0z36uPwb4
amk1xqjyDfpZmisJdvX0gljAMePBDyfuHSnY8m5IxuIjkT895vidUXfUMOEFFtaK
NV3bCcSa9Swc2PwJ+A1HkrOPipBe40LhBKE69Ckm9YyGc2vWOIMs8fAThPE5LTiX
4WPndXBzi3vaCSA4XK1Obynxwyhi1dchLNT3YbFR9npoBIs/LEWy+SGmxm1Zk754
/cSJZjZUv7OmN0wzfMhaZQ==
`protect END_PROTECTED
