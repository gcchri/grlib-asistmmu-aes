`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
loWoBtIePI5A0KNn6btobNTcHEg7huvOhqalvODdlL+yuS5Z5FR0azP8dZIWEJC1
z2lTxIJ9xl+qilaM7flZopl6k/2fnHPrMNsyw2UUpcG1MxLIkfVL0c7zYiuRrCzF
RxIT1bjSsSMedDhNfLy82TgRo2ii3+3fdKssLYw1jHP4eRmalCW0MhIzQJ0lvvGe
i/iog80B3VmwaGPM+z7ZzpuBJMV9t5hzz0/X4kiaIW+V+NbpakhfPAkQGzlABfHY
YEW0KRvbTjwD1U3yiJb/oGdfpnQJV+aJ+BfCMBfDjywZPNBPB0rFJUvaW+uVUFuf
`protect END_PROTECTED
