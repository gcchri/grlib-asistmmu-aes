`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2IzewfQSNcOre6AukOdYYd0TVjDcA4CkG2TErAi76vVPqguV5elt+QyHIU2jNvTj
BoZazAulk/z3NTzQZY9NF8wLtSeeiY63RcZ6gG7nKMsKi1/JF1At2sw6WfYbPea7
xAnm4Zh97Bs/7GQWlFpHJHu9MEh8Ij6aFASDlMYHb8ChbNr9nB3XK0Zi2GqUIJ58
SNoyB9OcXIkYpWIxN4nJROilN6IULXtOLfBQkOnKLd7wSMf77f+Mhx2iOgIyxbd+
p+KCqrTQulgZ8D699xN3D126ibJ+4o/2rI5qPnqShZNry+UU3OJxsKdeEf6fhCp5
ZujH+kjkgl+f9+6t+1wP7U9O50tjWh21I0Cy08zApdyNKHQIyXV9839DtB9z0UxM
CqNjt89GV0TLO6juwwiHGMJ8pXnwLl02gt3q588xaHKEjLrWfSkcruplwcQWH4ZF
OidGJZJpp8v9SYnPv4j5FnQEJ/Al2MYOcVYmfXVaQuYTCpQC0kFg3vJwJiMNXnkz
mjXIXun2PrxSmy9VD21njMNCoQVhuVtkAp9I8ztwVZYeUAxnoLkbu/J+oFp01lfl
k79jgb8EijEKNgLGOyMA/zwAVxeO3XFwp6Z0ZdhpvFtxmHmyqRp/f2wIJIZlJ5sh
Ze2TZvwNE6PQYwK/yQLVBI+E2eWzyq9da/V9+U0jw4HvPZBOdTTeChnTwoclV7Xb
JlQFmXgocNe+7GX3xh/MqS2Cy8y4DrsD3CiiBGqnjNVi81fLML9sM0s1Lg4PJIdE
qNBbSZxb3KG4DjGQJNYEf0PK+5/d46ZI3VJvoj+n3kahE3n4oX1L12YQJPQpiFAu
X9LxMac+JqhZdGs+sbeEfEznhyFz1TWZXNBp8Ms9zzstOkqUOgGtHLGxLOpUnaE7
G6Zfq1NDJtcCgRjj+EDll97PO+Q9s7I0AOhI2qDGqqNble+k3h5R+acbD72DR7+U
sVsXe67n1guR/Or8jD3nYqtVTiYVYHU4bAFS0adsdfYF742Y/hj85wRnKx+87B5I
wVXLj406rPgNtwOS/iRuMDX1x7P7kDXNuYDtXkVwXghCWJy69tL6kPDbQ23pa1at
lySKCYZo8DLlfRDepZSbQZ2jHvl/tU6uKY0NWIgoq03pkRYnqbln85hpHncmSSZO
PXxY7yIy+fKAUz4FH1CroRxpaFh82hd2iagYaNDuS21UzZ7Npo2sJO8iLIuRTGhH
LGW7zT2dN7ngl/xHioHF6LvJ+PhxUqLYynm8joJNKGhrI+QcY/sUrloRGUtBMltP
X17iJvUv1mS5wdj+OQxr8N3WFqfwtyDnQAqcn1pgpvz/k3dchzEmWND48IwWia9p
xSMBCmew+F68+vQ4zUNhovzcy5iB+B6QO7bdip429sgJG2rd5N0kRIjI/n6WVjAA
BM7G9bzpajpIGYXIjQb5cRjOt25J4zp4RHiTl1Jet5yad4uTyWJj3X8oX28w+svQ
xv8rE7CpIaGF0gFZkcLMEqdn1S3DAz7N4+0rao9Om5rhEDKl0eISQRRbbyyz8I7R
`protect END_PROTECTED
