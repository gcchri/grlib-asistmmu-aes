`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kn5J2y3eGhR9NIKxKAS+aEshrlqRfk+bN6/Z4xuRqEnKHz0PtsIFvm6at/MHKxr0
iDJ6cQ5IzA7EtY4df12A6h53jkaIof352hBQ+V55N0hy62Jx09udRjyKZRkgWTSu
ZMNRKZsIkkxzl8nttOcgCT5ZfXX4AekQvWF4VyQ19XDwqtFzBfpniHiKxSFZcpB9
Zslc3iwyX8A9aIrJtBvtfMcSC8Arr6KQnMTj/aRymqdYfDm+0RhsOZxjSJ1TJ2yi
WyMyRzhYMdpzi20ohdyZRPM1+PNWaOXJzKJhcALU3UPogzFbdbcgXDUnVVj721XD
8/H2QpO9wBhuOwUsE5yWH9oBvGfHcY3aQ6HoE6V9/3Ww7SexOof+59IPSpYxfQi9
PFdV0xSGvk8eD3hlgEcQJOnxkcPMDRKlMDEUiQrCi+DtixTEv9pd8mKHkTb4hmeI
vN/Oj0/rcKE+5BpwnmVcOKZG50n86H2xqduYYmNG0kgXGb36sTCIPFsKE9go6nth
u/Vf1eD0YfyYD+waigmFAcalqoJdTEAm++eI6y6N5jCTmq1GBisJuaqf6Kn3Fww9
GykJrGEzvXLxAOAfSiDljVjabGqPKiW50GiD+QD4wONi6UPTqvrX/XH+7DDLD+2B
/AXmpWjUMHZI/zJHrX05gA==
`protect END_PROTECTED
