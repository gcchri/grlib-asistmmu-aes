`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcBC0Zgxe7/iwFURIzDKGpb9vNd/k49+aE2LZcyU/94S/ioa44hbkjsV8IjbJSSD
J5+IY2nkl89vpnoWm+gLqfUlc5UcuvEJBbXCERuoxwMMvOFvL/0ooHaiOflpKTZm
u9gCcqEKJgdx0ytccDd44pPdprReUXqzsyA8mMRrqlbFxkP9fSCB28jM5QGI29BS
Se6ovsy33TZjriTuZqiexd+Ser59FH8j4nVO0E6MymKzWAjk06Tf94ntRv0ypRCl
2bcrJtuCOQJTT1qgQTuuPg4PECLeoAUmNqcCHSY/UtL4BQoT3sJzbAJjDzbClrjy
WI5d8o3CNm+Cg6hdlhGnNumSxvplZdv00ZwrQPxSymosNFcWggG1mHfsQbyEEPHC
7ULnakQ1YGF0a6I9uiZI787kuJ109CP3ZT3KbpUpu++T2XdJ2+vDJv6iZK4sqfcX
FmIHVqUCOLT8x7lrJREafwT2XGP65YE5xz5l8G1a69PfhSccCpkYv7fnWS6FFFd8
SAGCblJzQ6Mb3lLxHI4V+FxKFpbSdlbNWUOFU5NcDifkY3HPSz69EjM7Z+2mBVgh
LDMHsILJK/uv9RY5ADblyRiHs/TFwWVv5uZ5aXnHlb74bmlDNXMvKOpzel7ZY1pz
`protect END_PROTECTED
