`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3BTTRXP/Cn3/J9vymFn1A1MNPVO6Sc9Hoee+QzM9ssRlFLbpjXpN/X5tNcpde8DQ
wsrDMPwrrF9qnRq3ZZGBLvNQoFsR1/oQcEmhSr4UBEJDgye/DnUvaw/pLCLAnmq7
pBcRbbjthNG30Al6p9d1MC+fBTuowRZXjv2KJb5ZTSy5ekN+4A9DDkhKL5j8wuLh
nbpoctKKkeRiheIYWJXKEUrYnJQWyY6LqlZqS4tvIFhlJe7V7SWcJwiRLVOjPCJ/
FQc/yeGsLyOENhLFHIvXwglJ7FBoEcvVo30XNfEmC840EVpiNJGjvpHGAiPaxIM2
flY0CBIOQsRxphCJA3n9wNj/Uq1PnAAxL+pHEgp7fQEY1ytS4l0DJS0WxSaMXo1a
RV+VrmCF3yX1wvf1LFJ5663yoTfVQvdNzzyoLhPXDzbRZL/JpGGqczd4/B3CPKus
nuVntDpVHP9DNKAQzST+r+FrvCzZFmHrPCx/8jHG1OqonIKgobwfTv9EBs2YO6zv
BdeshT5t+Ws4jV0IPwPCxwO6ENiDOd0qhzPD8Dcb3XbFJKqQLFuBsBbaFvvhZXXD
D5z42byojqr4nOpJGHOwrmKTm6jgNZZ/P7t1EYPOyqLE5RARbyYQc4emKdLJ2VSK
7aRJYFweb6y6NLN8tIVSYLL2qcKZsJd98DZKaMo84/XO2RHcPtZ0i3omZ9ESgev3
/B1qdS8COSoOm1FF2+DdNiaRC2ZDY97MWMuBP9DhItukSo0zXMbSfA0CRcAMypo0
nWrwsaINV7tKNb+8VjSlMLtrHOeqdYelrk3BPozPvnQaZayL0COS/8PzDIXyty48
1RiMxXcqPx4Cw4MVnZMWkqPgxzqsCTQtYuQcwrZzYagg486qD/w8oJ6+rMe7tzyq
Y0C/mgoBMiNYZZZVpNo03avilPfme/JiOJwL6IdCVI+CrXhnTUZxFHWOJs8+JCe5
wNSCxSuO83NQExo9YRP4Ydr0kFfoAxuyXscrA9kKaly4Doy2Dzt7bGbSspo2T48/
XgQEzFyH7HB6BrtUKoGOzh6DWVQweJ1zPa85M1foUF0=
`protect END_PROTECTED
