`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmDjK7gLQiQUZlvGOYTjM2cyz7p1WK+0AiFx+ALyPPadM78x8NjllFBnqrug8gA8
jbtchZdKNE4C10L770XqDiz0riuhshJFfDKAPI8TOND0HrV+GcSWATfb69F/d3C/
Za3VEwCm3uzSEpuaco3di9eytovfClU2fQoKIy2mHLYmNcFnohI9v/WyuISJ8wbf
VQXmVUPK690fSzYQXHCiDh2p2CmFexDIP5BWFVUSgn4lJPdbpNCXnagdzWa+FJUV
1/CFVgeUcC+mRzuEZBrZhWQPe8hiiwasHHexe/z3HU3T4C3x4U36l2If5YLs4dof
DE8VqUKcneIhSYZegp0IwKD6GZ3QJBzjZoGnNvN6AAPDc7J3+9BvgDHXasHrbRtg
uoGlW1U73raG1TJ62vqtoNMwGqyzRrS/lbAnu6+MYSOrBhRPMHSq/fOYfPeU+bPI
BACY/Ym7a085rP1/VJxBF3tvT+XyY3yyzYBFwg733RMXMsc8PgSCRwd7uj3kvm8C
Fms3J9cM4Ztoa1hNbA+UP6RvdgAqMx74wQI+osWuS6w=
`protect END_PROTECTED
