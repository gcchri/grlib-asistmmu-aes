`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XOwx05A6GlTtVQL7ZGaomBHzYcCXfI2DRzKqNdRv2R8+9W0+lrwBCOVFgVlgPYa/
TyqYQgPwwAvlHlZDLuPiaul9tUtRQ289tZOvtW6gitLk7y3gKRVGssO1dKuheNTH
bDKzotGbq9gv9BIolkd74o75l4ClxVdR/MVgdcsNEzOrtjoF8EnbBFjSCtoiL6QL
g6X6rmwMHTkaQ35lyWU0O0+plMWnlrpR9FGekDzU87MXnKssYkgOCR+2W/6uWmJW
WjTuxiadENJgCa6Zfx/crURvIwgCldhnuW4yjzi5GkjXfFlGzsYGL7GORnM+UKS+
Nrev+vk5vwuXxuI7yKvHrix1XAUo2Qb2HX1zHuwYkW9DXD8ZSRy9krP3vhOXbaUb
uJIPQX57a4YHCrnDFRbZP1IYe1KtGwkCcrkG6aNRnu5MTy2ClVPmKqA8syXoYaTo
s1nJ9RXbiXR6KixfvW/jg+rV1fMXkPF/pX+rdLW7oIp8fDltY+P6OzICcT9+xPkl
aOK2LJDvuIFOUx0Reu/DCzW8EzPevJVTxNPkSIEJWOcsNeWagtES8r6lNOkBnEbI
UPKZWL76KSiROwYbFjPKTc4YBjcPk7gu/FZEoXUb0nRVDEQOa7bh6Rmr3bDelv43
TG8njwnZRMZ1arp/MVaCyrrOHMW9548zvrEA2Brn4Q1LG5el5lM/f/V0cympAxlR
ICSJ3EApvJDHQCuPHHah0kQOkFBaV6H2cMvn+4GwBSyqwmAgA/BW+Btk+qNatko/
kjcKXgWlfnX6MNMimxG+GF/Bbyv/DoLoV/CUdNkyN1rXJxnk8T2Mo+ah++7/YpZm
q4LKlc3hQZNzlclbXQaT9GFfCkIaA1TGs7F/jXF9bf0S5sNcJdGDnJ5+fYU0Mt4b
5+tWkFSQAtFh3aRnE53E4Fbu3zTOfe0A55748VkMJh3tjZIO5ruE8OHvXikTqCxO
3+lzZKnQM5uUBarqStYoJhd4F+Cf++HV+jaBvO8RruU=
`protect END_PROTECTED
