`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kE/xWBwPPNYfgTNhvDHwNe5K25wvu8sdBFJSkinQKnKBEHM5UsXNXzrewCTMwIGT
koqWlc6UNovOJTS8g3mRhFOa/P3YpIggA1sIcQ5c83JvS2X27GTEEjeD9CCEVBMo
s4+WqWr9X0IZvXgwsKrhDbHq9AJEgkV7r3ZCHhLynmPtpnwkPFLrAmQF8ex7wTyH
2ZTu4LJHmRb7K2Dp5CzBdoqHndkLRJW62HdSvTPtuia16mt/eecFXD3NZFB3TDBs
Ab8caXo7ShHrDlMAqoP4hfcaQ+9iEawqMIj25xickmLnw+LRG9QSMrlZV5N8tNYq
W+MjZ9p2HtEf2srSQDp01QAs9+R1D5RKL+JvToB7+6E8r4CMTt7MDogCsY61CitE
kbCiblXbLnISyiaWQOvn8173hg307ZTnATzxNFSF2UxrJ4HZjQm77L1JGsZg3sGF
`protect END_PROTECTED
