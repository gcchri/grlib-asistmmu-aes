`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G1tvGcOEfAyAsIZMIMm0UdA+iSpvehdAh+oi16johCFyqAqvK/kUvdjcpuGcvO8o
1OKWZhZAorm+T9Yqg7GdFyvheOXS7vbRqW3TweMu6gkM1anyPNBw2Gi8+1sLgEEh
SL2E2WG4YNna1O08pOeE3bomU5/Z/C+LF9b98xpUA3Y65L7u+QNj1blAkVndBoEv
2BMwyLoKTObcAeQuHQaQL34P71tTw1Iobcr4m06E7+6axPU5y3/t35WJfE8hGWHE
Vb69Ke6HV4q2yrskS2/p1IXZAqiZJ4uma2pIusJdEpbc5Cxqqjqh66o9vmlYWTWE
BZ1Kw8x+RijOIlAzIVAI4DE01Wf7udoc8bPOd/0mYuFCcdSWv0slDi4BdAR9mzXG
Px28p2lHxWW77JaX4O+zSEeWRWIwO/lgh0INqF3oCM/HhXRQ46QbYOAzUWtKYSIz
utoeZV6mnaLMuB7CiHmDDroNZkNsAeSnkF92AtyFO9sM1wlVe+WpCaqKeQNJb1bD
`protect END_PROTECTED
