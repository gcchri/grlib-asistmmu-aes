`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwJ9iwG8KjPAyDMfUeNKFL/rt9ZjLfeOiM3kb7VvxYzMBayuqo/VKM3WMCOWexfc
5IuCEEW1KTC7i+33LKr60E79TASshnBJnS2GKC7SGeCg52O6kYxMUk37NkymUcae
7Y7Dtmbph+dfgwKJZqOBMJni45yThUTNEuE5NJCPldBKjTE3WOV6Hi37nCDpAF+I
lmp2witvZmJbZTrMNX0zTXqm7Y/IOm8Fxu6kQuM4hlTufuMOWF1m9Fy55xmBYgZx
8Fo9TPS2AHxKB5lTrJxqqD1GaH3qZ4uGoeCNe4bhyYS7DHVnFnK9gfRMiKZz/N7M
dO28fyIqlK96AdAdFpBuCITWjWMolo56pHEEoGbHriNl+pQO5hBl/vgbJBK4WWKV
y/etnwLtCSRwhr/iFG1sBcVV6IBEhEqD9EHLzc+LRscTnaWcDHPmlXoG/uYs7TQQ
5r2puXhXuaxybrdK34JW9yFb5RohNbU1C6PJUTPIK4/KOxJyhzJSFvKU5PlOYFhN
iUe0Tqaq1KzOFOGJv1WKG4Ota6KgHCI72qi8QQIycsW+uLP4BoIq7pdtZkCYet1X
7u268nE4nRgXk1dFCXHpSX0pSfPgSo0uPEQua0axoPo3ttPU5zzXVmpuW76EKoy0
bGtpLkfS2qpEfa0eOFOaZ/VBay1m+OXsRSG2Pw8wSP4fCtSIwKRIMxkPUiqVkf46
caYCgL5Zv5OJ8T4yQLCBu8AlrZFnHuv/2nuVGb+MSLBwxd3qABmjWcCxurE9uUpu
sZqqTXz7B+zfFy9ZVbqO7PiE3NrA4x2MZBffEPp1uFnqVikhPCbpQiFp6fnvTckR
548+pfR7iSIELjQZFpmIK4xEs2zlb5HobP8dqIcQxjmD9RoSS/K/zfnumui6MF4T
J6XbqaAi6dy7ZOBsnMHjWpeP2gGFE4F2zTU2T+cjr8q2hnhPVne0VS2AbURh1Ahd
`protect END_PROTECTED
