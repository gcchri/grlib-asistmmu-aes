`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
++xPHN53uFfTnB46P5djmNg1N9oq5QkHrobN/GLf1vx5yZsoGLYp82rRBsCFGi22
sT9L05Z1Rl4jAJmg3/hJ02euyy6z6U8v8tw8z7xiuzBXcD+Na89rN7cu+dJw8SQr
LVIuLv7KGfyQOhF6RDNa6250v9dddqTZz1xqbTu/MP/F8n9yAfLs2h+HuN/2iiuW
H7rI+7DWRYjvAqN7eiQwlwslZI1hneEYsB1D/Y5OMRi9myghokM+qLijmQ4uuxO0
Z4NbYOuRvMfP2nurDKR7TVBQOgLpRUjiUgOpOLdKRAaAod9Ij22PWq0nCF3/6DyG
hcKbm+tbHQQi6hOXJOAkvG9obKfthYdIrezNjMcpujGIrZflnvC/wMLivWNJGZg5
0oeNTinqwaF5XtgHQ582x+S3E+G4Qq/TXbSza9m7a6UogrXx0RZgjz4HmavXX75j
XTW0JJkrUV8e5LSjWV/GHmHPjj30pKZnJFvbMBdxYznkJj0PnuxexwyNs4gAEaEq
bxq+xrtrjpos0I/SjKwlIw==
`protect END_PROTECTED
