`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNgYnCA2nwOuY3WANc/bYnV7KiCp4cGDvcjS6sxu6NsTyyeSO2RKEeBIxgxt1yqD
7BEKfIOQ1DmKk9zFKagALgdyOMn7OD/zJivAndkptQ/GtkXwiLD6LHj9CmibNlxS
YTgmCvoUYRlVPjK5jAi5NeCKpZg/I7BRTKzksufm/L8X18M4BDCIuFMpnSeqzOjj
2RF/OuadD7XSC9oRa93hqxlL+9jludNJWBTqFFTi4VDqHOKzSCcDMcmvk6XI1+Jp
99kAUCoEVg/HdCJLIS7gOg6fAC8/fc5KdNcew9+zFDWetXQ/qG9Tm2rCcQaEzlWm
lnDd40Pnpz92lqp4oIeWinsCevjsaZzqWHZggp0eNqNQv+a9+BXE29LDrVRKxJpO
d3S5Twvik8l85Ufznm7+Unhlh4zjwHi2Oj6MSEW6GcTtlnJyNRJfM48WAFDF1iWS
`protect END_PROTECTED
