`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hu1CI7Lv1y67SWXfzvN7to1y48AlETRJliEs1cyKVn7itoII/XuamSrVxpCSIapg
s82hrfbViAHWYZRmb223bPX3vp8vUePeFlob2gf4uPryGax1fo3sA9HuTA2uxcno
XJK9mptjZGHMvo/NxsxOpemHcDLAb/z4UcV/dtF4jfw/53TvbDNWlhA1L8gxO/80
gsTuF8X5VhIa3ObqgxoTpaM5NKzXDCzLY2AOJSAW2awh8vsC+t+hvuPOw1O5GFe/
oBqFpVeRHyR1YcSL8LMwx7iOnXLbrSDoqWxLGBXE8YzAvghwL2RdsUhQ41GD2qh3
zmCS9xto0JuHIS40BFwSPed4ij7ym5jyunJmeQPPZxuKF9ELn3lUt2g2TPynfkCv
Q7sMKLMEtYKxtptZCsHMXdzxRE01PpHZIpvAgZ1IwlM4PBJaAZSEy2kGMzwo8Drn
N5+fKfJiEipePwB4ivpOAV/BNWPVn2y0oH2WQhP5a8s2jHHpmd0DauADsloAbMwC
auc6Xeb2PB8oUTrIlbQBigt+KwqCFQnI/kSGYzqENM7NHqzD+ZqAb+VhStLWwmQD
`protect END_PROTECTED
