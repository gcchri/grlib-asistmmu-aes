`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aYEmzY+rH4OdeeHH9j4QhH1El7GgmWIHNQZlYNkINgvTogLYAaQbkLZXRUZIzTQ8
mIO843ccMFczvjiW1Gh3q3dRroCyExup893hic/YYgRRSlslOUWZsSNknoUJ20kL
SFSYka+C6p4ytInUuCWcHWtwEQJQcjzfI78OP7S7aKuhwUdxrHc55ly9GqKvuRV6
RabbpvPtFqXnH/puyHalMLh9mkl5Hr9eDTFSsToS9449zxnCQ/ZJmBzQEYyE8gzg
QwceiZ9TG1dduUIT9y5OfPeQkqJ5Id2unW4B1UHQuuAhJUgGr9gJI8tBkko77kON
MVUiJoFRc/N6buyMcLcDkA==
`protect END_PROTECTED
