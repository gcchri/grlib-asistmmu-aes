`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pKjEORy9j2orOGb58nuDOPnctjU/0xpsf0RKgwU45gPa8ot/u2yvHCFtjU1zXZM
9+b6oRsdJExGtHkEs+Sbx9kblMss7kheJShp77BZQTzVaMVsZN6/ylqvm6UzqYZf
cF0N9F2lBlZC0PZMyhETvjeyoQCta2zj3p2p79MzKzcPrAQDlKNY1nMIHGLcTED8
+/EyaCCGt/Kntooj7q7A0GtgjG2PbgKhLIJgZ/9G0sHlQOJGJc+ye2pRRr5TG4lr
3utTfjTeeE/sYax/2wmyMzKkzb5Q2Gyl0XGkuahxDxUbCqw8bAVB5av2Fqqvs3S1
Klv3kKDLGwZOhCPKTYfKuxa/Do0Z6gL3zhJhNVZuCRT7xtqKBCvuMfX2fRcir0LQ
koAr/dseScPpBcq0EewkBCQbM/MLzhSS1c1wJWRVMjv0jczQ2GPNrMZf6gqvaWst
wjDnJQ2bqlJx6OchULJfGs7JZZ719Igor4vJ32b0Dob4H03AvhtOlQj0kRNjkrqh
bEjggVhzIP2LlDrhlAxhYuO4ylfr40jgKnfEH3QL8t272m295PL6amiKozzeQUZ+
qMOXzz9mHU2SLJ3utO6eWoO3qy0WfNVVOXLqLbP0l4UYyzxADioAVp0mn7ZsHo8A
aO4IC4ABioo6YVQjKiocY2XjKrdHoFysJW9pxE673S1BZVlMgatSGZ5UqxQUfaas
cwzRKhw4yxxU3/2ZABu9P2JlBKQKHzt4pH3SUpgJYSuvmI6Tn+DMT0o0P6EoFgY4
VA4oejPnWVnxxGtplegEhjLEoaAa9P+EXGhlIAEq2I9N7LVTT0nVm3py+OlxNF+M
`protect END_PROTECTED
