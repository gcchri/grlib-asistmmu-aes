`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bajlozFIKLTyDm1JIeV/IqW6v97zc7T5RPZ+Z/LIpuA+gSq4wJV/rKTveNTdkKbV
aqdFcx1uxNFZHaZlNbldx1yAR+C7k9gE6wOzI4SK3YUHv3lC2J1hKNGNqXkIrDjw
O3CwDSUSbifkM8Q6bwSVbMXHM8c5/SM1pg9/9xdAXvJB7IVagkCqdAaQgq9DHRRj
Ct6Pe6I54tVycEFDcBO16taBfTG6M9hTe65uI3ee6Zrtvz8QWRAPQyzJnTN4q1xp
+KwZsuaRPvjC4jM4Kp+PLktI2zva26flip/Yah5JFYH8dtYkiH+GgjqCkhv2eTHE
lQ2UBZaIuZsufYR5JEJvdf43iV7eqOQNgBFowu2cRFx8WICo0Ny+aeuZFNq3xyVC
mJV90cgt5jKIFPYZrkIKyGvD7yIzYmFBbYUG+NCeRoOGyXboku1dBC+BYYtwbDHm
HOuZ8CxMd4m2hCOrc7Z4EABMyPRixHnfiCLb4NzQOXFeD1ZXndhnYtH7ky9w1MSV
R8pImAsk4YIb4kSCo9sg8IS/Zkc2BCkooTTQRVTF2RPNUm1cLl9lcrR5333AiMtV
bbmHUy6hQy3NgiRS7my2XQ==
`protect END_PROTECTED
