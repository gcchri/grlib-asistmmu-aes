`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HODkVtMTgPqzLfgpxpUjRtcWf4XhAZIjI2NfCajvmzjZHvPM8uXfniKQz8JsP7Nt
N+r3y2SQw4kn1j8DXnOyJ7hDsUYuPV8bMoD1jpBNHHOP7PcXuPnsRhoFk75nzLPT
10RILwe4/O8G16uJ09KRhs3qlEZNF4UVu4QqtwRDQ1MfnmdAjTkZ1lxI3U9AOPFP
IdabsSAhxJDb0oBemOF08aXSOTDAl6LQ27BnxpMHgHimBhhbNjSpPeYXkBkc6zTK
xMYNENa3Cq+SiynkCUferr0kbnbH5d7TawoKqc17aTxrEg/I5xLgyObZBZoRgxHl
1PJhbchvWXaSaQIU8kaZ/nHEYK551p7gJGi9UryO0+0JQPiV0ZYEPHuFf7uXZim7
/KKTguzOOXBA89/PZ8yVqqpyY/gTEwrlqjbO6qDZYOmC+Zs2jwKox1G09Xkr6CT4
olO6NUsGLCIa2AUwouU4xDNBSAQo9pf0lwCbd0iwvJj5UOEEtMO6FA0APXHIOl6a
`protect END_PROTECTED
