`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r4zGxtwi+YQOBc7c+ArqX9i0uGgXAvAo6OGUmP/zM86RlswLS3C5eMlljcAkd7KC
Vj1Gm3TtRRvHtdLJHthuWmRi9u7EyqgqGFNUFl2d6niCY/KBuIbWT2aDYOXaLMXk
13XcyKdJigYOucDvMjCvMBdxaOxwFsCxbfSe3sKRaup/xoV7HWP0fPknwHEUzSnB
yyveyldUxpBSPl6RLUdGGsVV0AZ9CFHs1XXujAxzfRAgeffvPhCV6tCvtqIzrmg5
l+PKvGPHtiH0/B46h7PFjZIIXdSPj63HB4jiXMgJk5F22jYQjK4tosdOOaFtfFqi
MULNEY0OEvcZBAg/np2U9g==
`protect END_PROTECTED
