`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZrPDe9uzUKTVsXtKGUODUKXDBcRV/c0N73loFhhh0ytrXTlvqI/o8m2pIR3oKJn
DHeizltityZYr9J5pEic4ke/jGO1KO4isIHJU2I0JfAtlMLKu/hXNQaQ2BUnFgpz
UhgS3CCrxTqLxPyn8kHvduF9phM/n4ICuOORwClE1xdLRsb92CPHZcfy+cYS7id3
j/MS4d62GwyVeJWe3I/jopv9BS1H5GVNPR+qWl+DvLIqolvyrmA5cwSFK++qecVi
F6v4AkUrDJwq7G8vyPBqTasChHY3g433QqEZN2Vs0OhlpdpLGFHM1IE96o19qGIk
BBMStMbcKJ51E9uVzCwapdfS356w/KyQdmg+xnFS2lsj+ueVcD11xhZwf1zqvZI6
T0XHLkwwUqYmFcpmSVF0OT64t1CygD6eSQhgI1l79leC3Asua/D0r5irYSr+Nsob
q3j/nrduwTtEUMSD4rzR7j8uWvWExuygV4agLtOClpMqmWiU6YWUMi1uoZ+Dio8T
RpDIz9jN0l8oEP8R18KF0E8kcCTHLxnwQlGSxvFWj+GQJOHIpfJ3Uz5hS2YGnAV/
qji+CW4sCz1nAmpwqA/8zgo1KU/18uqcg4udRntn11VJdSv65rpLpH2T1TC/m9r4
figFUE+7OdkTE4yrWldZp7GaYW2Ci6p5E8T6TgaNgFPrZCp0fd3QvQ+0mpQKbfJK
tBBqoPKBjhNA+MjAMItqydOAAMNmZ4QqQMbTFa3any7psvN7mm2cA3+A8vzpn2z6
z824d1zdf8ryMhIyy7+nc1RqoMxK1OAG2RRpRxIEe9qWKfxhMSwPk1sNo9l17fok
VtJSdz6moLnKSDAR9C9YSpkoEkQZDsFPZBzGfy91+Gkb6cZ+cAdI2v4bgIlL6FbE
kOTWu3cGv0wwaJ76U2EzBUKpEXYQdakSsNwHUE3aoZgWLX06qeX5I7lJJHnDMbiK
aVvmLviKFbqg1tDS8/+U5JK/ER7LcIegqNF28xHKJfhX2VFb5NPU7W8aA0GoeTMR
5xptKLfaEv4BQlO058IX+WKHgI0SSTzsw/7cDXgDkx/cz05k4HJSXfNSWtcTRZnQ
x9fka//1/pSB/n7RDcdRvy5iU0VWnIbmd0+yQmNutaRoSo0kwnbv/nZx/xbBP3FK
fPa5uisRMTQKC5d6AY1YZhHrq3fk8+h2pE/hTwk8TPHSADkVrxgv4WV6TGkwLmHw
mhui8AysOA0cs3xpT4lQ32Aizf32oSiNYFSvawIZSFOxLAU+uWLMsNJ2ZiKmKkXf
VvKNYca0EqdI+akIj+EKEZ1jybt65+5reB0uF32GWLVsPa/gR3g7uyF63AOR8+Uk
f9BeakA2f9s9hnfCKhmB0lN9xi/6QiEBToiCdG+iJgHmvKgdXOm2qIF9homZvIMF
qEOXXs96Ken9SLXViFEq8W5ZafVYm85YKCQwlsY01InCP9nttHPKO/sN30h7gZiy
zTrOlVFwK1bCwCAU9ZH5F4LBetUEl29heCbhHIomRxotSZQw/bySvBL1TgUAe/2i
SvVh64BMw+m33P+WdFVZlBUtj+3sadXTYFnIYuOsSgjpovVS9V4byyHHxT6tmxxf
jp5Q+zZ9f+7eLBdzVdbCvIEMJOqhNwBSuXgOIVgem2X9xy/a2/8mjifERF5illUr
5oUsxgSHtNhi0H5TNEEQnm7IavR/ouV+VU7m8wG8apsKF5StvWEoRHZMqv2xKK7U
rAHd9bZs3JUjrL2ezSfEPQVbNBIvIL9I9X4Wk4FvE24QgSp1Tb5TlezYPqcDI6jf
nY9iCYc/JwdcWJZ0jUc1xmTkkDWjvpSoKIfbHFqAk1l/nwkQ6RCMqs7g7eMolM2t
0WzWa9u1cOAKkbk7GbDcJMGNVGf5rc6/H6oOPICPTmMdaKJWdQCMLZLAP/CizTWp
mJUnpj4PMVjgcbowZCZbVQB3DNPkwUgzDDYkBDn/NdwzeQW/QLEJr2cOOpjMUSui
ySfgpXyCg0dHqhNEoRWCjAakCU79/t8zXkxKZqFNZY520XND6FE4SBESWUS/aZqx
gPC8orR+h0mMZha6zMriSdfugob+BSobnZaR63u9u2AHR6H4s37yvKV8cEirFp6o
xKehXnf3rUYL2fvLTiOGlJ8Ar+qoATmm61gv83EB2mjb6WDbsl5PUJsWM5N87TdS
gYX7vCcoDwPAhv7YXSMCE01bGrh3vwy7IfhTDuDkdoOV45oQsk3L8bLbM79GxTpr
W606htCFtY1AELnecoHZ606jL6k0pU2JnPZyTM7oUvJxgtkB7kmBZVgUzy7xYXBf
YhdLjCizAGH0Vnb3vYcp8g2peptSMtxn0PVjo710SiElPmKpBChEdcm68fDAEFjw
nYfqfQCRSARjbT7INbdP+VzO0ZjYmC4RAiENgSte01hBuweLG1YzIEd2kQh4VZRD
mJlLygU9WsiAba840TUYXkPhX7tCMhPheg9+lSp7m+jjOdbN+dhLf294uAC8wR10
qrDG6fIEm58KMJke6lf5++tNX8ss8iKHLdJwfIU2NWZMKMq/5ma+oA0ZRHuw4PZv
4DkSG26sFKgYDbPfgB5fMPcgaPSiXd9MW0VCkbTAYhUQ2VTY3IKGNe1GtvhWMpJE
+zQRTUPFk0KBJmO+nj05oFiDr8EhpSqRYj+vPT9u4FbNlGUf74JXUg1zeG5JFPbN
Qm1LyRvpukw5tAd4Vw9eIoOSL38eVEaE0ttuUvo9WVrlSTZ0vFYNMTQ3s9nN4w3e
Hvlu07/VMFdcheLX2OmdLFaoiGCdL/lhBXv9vvlHwysclgVrmGSz4Ud7XELXia7a
qcvDTifKS99x/Y1DyAj1FgCkTUqyENYNAQaQc1V5+L0xxXHUMgMsuS8F5NCLc6Y0
TwKYdaUxpGUtX0Kelph3OuhGTNRn9ZnwY549KX22031JTU4f78+EUnATat4NBj1u
eK+4jItJVMz+lC+lmsy5Q049sHrRb4tILw3eSlDA+CU9VHv6gFmVwDW2QgTtSIsv
qN2W9nbx8pyap8tYdh1no9x9uOyWUjLPKiqFlt3MaOtBqkIWLFZqFVgQvzw1cjZk
kpOs9XA2xMB+39sGQlrutUGoHkq+lv4Uwc6Jq/AkWxgKPAID+hWrXHihrjivScfc
/BhZHU0beFJg3fwp5x77SmD2soBJxlvyhRC/SVIs1bpyVvkXJYiEII4/2NBxCAy4
Vv9se/y0G1dGsQdN0SJtJnAClCcUoWVls3osgKCvJgCdjtXr7eKehaHYtYF4drWd
ieIwkpwaXTP2z1uYIEc3up+Tf8sKSJkNu2dZzohHinHBfaxLSbtO5B0j6GDcWEMx
Cs9DWuLfmsDFuGgCHA42r5hl8yf30wKyXhibWEXOQ72wNrZg+zZIuK/Iykd3Stti
p6H1Vx4OKj4fvGiieWjVMJAFhxzIarFxZZfLdupeKEgf7CTqv8/uFy+GjRyF3B2G
QS47IjC43nUB8AoDF5qfBWw2fjGOcnsCQFLM3GwRGJkmrOCCyYcqHpen82PtZjmC
cJjvugmMauN9Gt9wL+tYwA7e4C89J4+4bJYboTwWMDMB/NGx6yw/DHsIj8UAjmG+
XzXvUDPYZ4ybD7aJ5qgTIz6WWPyWU1PEdts6QRyvM7qgvEjMAj81I4nI/cr7W4L9
47KWC3lts2gTurvBQ0R1SV/5wuzyJISS6gevvlaWd1kVG/soxLc6R9IT4GTWfLIu
UedRIHzphc4yuO7P2vK4Pu5wrMCSNNTRjvmkJr6eI+xR2e4wVUinlYYq/eTj52Eo
WjcLwdlY5ePQH+4tCSlfkI7rAWXbfsEcW1i4A89P9a3yLPm5nF/rwK/7OKlnKFPx
m1cwq30JxL+4Iq4JzSzVrgpuI4svvog3yEqGbum7qB5fq65RH4lB7yg9F3MqQKsb
OH6nK8kFteSdGsO/xUaOnQmjbeyJLvvveniDXG6VRbfgjGlsXoNr3pztIWhA08Qj
LaxZWP/L5tIihO0I+O1BlGBeA5W0pRiS1OgdY6wHEAGfNizXVS5KyYj+vb+X7X5L
FseXJu1caUqcVY9ek0kOEBloCmfWiJ0SLjC8AqC+CjJ0+AXj9ZEORcWLC8v9Lfvc
r9dXDiGeoPWVIdvDcvRNc0Id3PzMGznCBtwbframggICDSWdf6c8ikJMu1nkmZ/s
`protect END_PROTECTED
