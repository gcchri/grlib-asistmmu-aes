`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S0d7b1k5GLjtakkHuZr0Ke6mYiEmY2esDgE/ZaaAGOdqbJaCGOq1DxfGLENr3wmK
pX/Nz1uUbHvgyzhEb7q6TPI/SkhvQDNrw/cn5iP055wAoo4Qp46e+oFQkhrGvuvy
7jpFMdTp4b0pCqO2eJifLKVZuVBqLKp4ZPeQJwFAL0Xer1I1yrLMMZb07ZHkcGIx
5OR2Efcd1ikaEB1dPoI0uScA2r2NkqMPi0+o+av4viVwmy3QMeoz4Y6DYxyxBOa+
SdTMcei8AZnPXwtTkOS2JipxrMlZH5heJjhGFsH6qQoFpIlGbsU2M0JwAVZOXzGT
69Ef2Hv0zzpIBXvcaoAXvGC9A0IcZspp1vEkCgbopiHkcDje2ac6TUdDh9xowOyA
R67LnrxvGOyNT/omXIZ3V5lQtNgcEudrok4B9K2j+5pN8Cns/j/8eS16eDx0mbin
TMV2T5cJnIDh0hMOIIqMA5tL1LugVJ8MqILNn8j9ltAGpcbpLQhnMc4Y7Hm3T/BY
/DWl7OgSpGKbIFftoaxVybI0u8mQaKag+OLc/bqxrsufdXRR1X2PrcxtXH1Itobc
V9a9v7hn1Z5ONWlv3EXwTlET4EIYBoLBxCWIWN2MSSQHcMMB2dIOxbspATiy6sAE
w7cs2rP+0L2mnyFuUw49POvEu7pUmR+URMp3z/LyCdBJA6Xh8MA0flXk2R9MUJes
OARFEijyEon1BDJX0LTfKQPOStigtN2KC2ASUdjK1jvr/QQs02VbTBloZBcZ+S5/
P6E4Q2HmbBRzuTw9EnhMoNrARuTJgY4l1i3uXCeNRsjBza/klPAFNw+SFHqPW21X
foNgebIAKc+nomBx8RWK6JqTXM+dTKjgAQbTQQhmOzkG9FW59r3awdzP1SLudZ//
LG56Osx+HvELTIXkWrmn+5cOKy5ekvNlfX+WFFUD5XRaaD469J2L/RAAtnhi33Yc
XDgHiA26oX9Ky5p03j1qiFAI9Uzg+Tf0W43ApyMaOTMd4enqLkeqE6NgpGZBSa2O
JYgLIiTCAPTSGJKwMC7sunMxC+1NB6WR1ujsHDKP1JZLlpDfW9Tl8SvKy4tDhksY
q25VrZ7ydZkCOWO8YDHSSUDDvl5jjotAzweoca8lYFanYuyfg3Q7vH3+g3STgrJg
PhweEFIbfJNWCOSEdHi9w89cls8fOI7DR7woqFLA72//9YYU+qyWIQsbUsUt5Gh0
DkECT7LkOwfqjcfmXtxSp6OuClWrGYfKVm9yFG4LzgRFw6wGIajR/9rJGwjEOOv+
CsaDAhBHt36oSnwHqL/1ljL0Uu+0wwFemWZhSSfi8tBwX5/6IdGprlTmMGwkjZK/
YH/pu4qa76Oq83cF1TNOKR1DaGcBfWbKHvzCSvSxr8sXVRNz01bU84yFQwNc84Dr
DapZOvGz3zzS1DrGcO3M1VIHKPdRSISktCnQ+E+f4wwWzJY+Pkbc6C498Vypaf+/
DEQOpn2C6uAvP9ZeZ/cJvS6Gf3UKYoKZ4BIZKb/w7CqfXRqrjdRCoHqiG6aUbPtR
QBGIlo5NIcy/gH/oT53W8YFITdIrLftwriaheSGAQqq+CE95OHqVuy6VxyTnKhut
`protect END_PROTECTED
