`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ngDTQYDxAVLMU00/lMtjPbHQkIq1H0EzzYQtaZI5Yn+7AXIQx8gYVWZBN4Ynso2
ZRvMBipZxfxV0pCvpTijAq0B/IkoVjXoj9zYxISzPOjNLmWEora0eCiVJnXyNQYY
ljH+GVcaBygxH6OpN5g/CnSnTVnBDiFfQjJMs3doJbfGKQDy7jiR0Dczrpx+AOUI
aenCUnHSpTcuCmSTQoNURpn4EBVcBJ4z0gyXm7ABc/DFOw6AfBIeZhUeC6De9SL4
dNNIFyIzP2datE6dz9gBU1xxsY9ZSAV829YVOEnk1LSuBF7ZeaVNUIPU5TaEch2Y
0NK7GxS8JwHI1I6LM9cns5P5GR54hCPAaCRKa5fBCYr16JHru1K5mkQ83uhoT+2D
IfdSGdx4kTHCf7uo3I61iQ==
`protect END_PROTECTED
