`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ejej5zogOkBOd8mR6rr0xYzjsBp44gpVhftRka0l92ZtBIit6teQ2ur6ceOGJPTD
gjpvqDX+MuvzYH6oXlX1wHDtMqWD6qHw0oHR7o8bx+Bgsbd5aDVK0bXwzo46blb3
KBu8/gUNK6MK/5EGjGPnl/Ig8Vzz2/uDDh93PTenArA/YYgrsLf4xmi7P8/nMRR6
D1OSFdGVe+6s7FyKWy9cirvqYViCFEndLP/XyyzW+Z4onyrCrQ2wNc+lOTfsCQCy
HSuSFe0ekrgxU0WNQ8Zzlf2MQ3vzac/EwbU5WfZY9fHk32X+4YYBHMTYITRjVraM
ULdSMlMqD2r+fu2gaGrV9kwi98T1cq3lhAMyufgNiTLO8uwrQQSz024f6NiUC8F9
ZYUooHa2UCCEJwoMRtfCpxQbYkxDhpmpWk60mKsWaUBSC4yG8RQHUbeM4tL2wdiI
ynr1+BUvFxldmaZGrePATYGlZDlq2Iut0mvJOVk6zWB0vY4Ixi5iXZaqqG0t7CK5
P5pTk4CdsEuNFaiOIR5ivujjT8nrhWg1wG+9MYY5h952eqOB/kBgj2Nxfl1mnBlf
ID3BZOt/duknCr7HrqfesHzSR76i1NPA6FfLwJFIj1duTGrF92GrS/+3DGSq6Zjd
L0CIwWvMTsqJNrLV92q9BsZ/KCBsTdqkPNOCYC5KzNKNW4h5pU1bEU5pXxJ5I1uD
D6VZPU76LIhZU080ztuBl1+fplFD+/RMkAgcrmq4omEgoWuiePtVZZddRIJ4QHhR
`protect END_PROTECTED
