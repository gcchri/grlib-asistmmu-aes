`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBPpYQnvTZvA+8K3LBfuycH/YN2TFcR1fdiOhwwhPbzFq5XXFnsctxP7Fu7qs8M0
rc3C0gVQHDh9Bf0lWb2J7lnVRyigY70Z95RPBy9IT7koMtv+fXz9j7Sn9u7JbRL7
03u+pxOoJ+qGF2DnFYROdKwLAtTq2ZWAna5RmOOPvVxG8ydPLEj8GUiD5kxQCtaG
yOTKt7EL9yaJHVtCDJaAfps4Dl4dpFcjDS5+o6MdHun6kqGy7/U8VLJyoPBpf3qV
FWBJE2RcntadARDYYyNdp/CznzAOuJ89pZ/69bP8e6vGob5zoO1PJb5ctDmyfVEu
WQDK8mJaaiOzjLjfJ3JyIDGnAztaP97Q/S3fR19k2VCeR6OwzcrIt2vQwGg0Yszx
WrQvQMJWx0RO67g+MEMA30FgLR7GGG8r0klqzyd9LI6FMBH+HuYLoInlFXndoWQW
801Ncfbi5X3oVyquYw9foyAOE+3YdwJEWZOr2MSEDalnuSwFnAjVLq+0+gv2qLsM
roSvquaZcpzx/t9qR8jLzdRko5B3s8qISDOELVlhVIE+jKlehYDACh1YFMWdDo3d
o3v7C+rPFv2lL1UKM++WrU3zULGhEZIDIIUG4CZKhhtNd24m5T/V73QSo3qeI3uK
ACQm8hAJmjcoRJuZE2GSzM6NS61YbWwymxeYbVuH3FQdivs8V4UI+yg0fTFv7upv
g4YyCU992t5BGMju4oQhdnUvWdWE1M9BrHI46dy8PTf3+eCQn2xWfOttxYcIhFAU
lTSZpYID1/Z+464NG6q2+gCErcKyJ9MDqBbRE41wMO3ar0j3QNsNC4i+QghnMQg4
TyRi3nIEUWxowa2D2JVlaaTfklZievBG4cRWP4n+Zfxq+LMBYq8enzLykcDvxQlZ
raAfOhFMXVKyuo2TkfvEJHi/oKoszin7Tje+NiUyJ+M=
`protect END_PROTECTED
