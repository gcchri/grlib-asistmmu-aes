`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FsVoU688Z2XG96EbsqR78EVT1Zu685BZkcTinhjVayZ0CHGkeowks2KSPwfQo/Pe
idXTh7Qe5/+tfnMghe7U78zdEfW8FRXn0+ugvIiFyXc5TwSqUXd0slFLwPCI/DQt
bZ//fzZeYLyMSZgoyd0Aoee1/J14LBalXE/RUTBU19rKxSZvPwqMfKNY0QPm30SW
6Mc4oCimKVRx+FET+jNWd0RETVtwLgW2aSK4OBEbsUX/MwPuj32VTm1hDwbiOsEl
eFo3aqu/q4AhbzrDBWmG2AF5+V+QElDymIJBav5A3wVb62tTQiW2uvRHrluvs474
`protect END_PROTECTED
