`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X2lTBwLleTVO8Ya1EZywEkciN5hQcuV6OVcpWJQWtnycITFX0tN2u8AeN6fQYGXK
sPiLY6yYvEgRntIht7z7+km4yyH9XlmKyoGvT+R4ZN5uzHr+mAMUfwq3MSBiQGvf
95AibxpaYy2bEyY2Fje3L+McfJwGkoQBoJkbtESl60VTHmnZR4kTrbs2iVKsYzq5
o1jv1L3qU1KBZ6/Hc4WVuzD/zYJh0zpWEEpbp4jzdT4R4KQQuhH8DXUYSclQOwP8
H3AtaaqBjvku7Ki9nI32RVOGPntCY8afVPDnG8vmgy1b/jFrsp/E0ZO5BXu1F/wI
EI0U6Z1sG5U9oR5mEmns6TRbsggLYFdQQGawOgCgyXnWVshjLQRO7h3zADrKUrk2
yedrykUyp8zN5DoY1Xzz0459T4YXPwWbuBPgPbDGhlsKxPm865s95WqXRKbRa5g6
UIlwrJYX2O3BV8UEwNKUQ5oXz3mqS4kSaUVAoXge4WY=
`protect END_PROTECTED
