`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0xyrSSp3OMdnWIqBeZeOTt2U3w7zIVSmZFX0xkG02xfbEeyNjK91ZLySPVq7gvWA
ekHooe+WKE9llAvBeYGBmyRc4+u4eD+Y+33NRFwM0/Sn///KXpZsFZMfyT70cEhV
2+1alJd7y9iosW//Z3IARsVTNpkpIermVvVTt3v6aTWJPZ+J5gVzXuLEhwNoiX/H
Og7UcFy3Y++eBHXFW/T0cct4GCLWHgTkQxZjKOnP6/2SUKEePC12he6ZXst3fakt
7ieBhvrQJK4Us4U++DaFCAL5J4s31mkL6X62hDoDN5CFziu0v6V/e/C+HfjLxLZ1
9Rv722MkieeUN6imzjAFdyYc19mDFE/FsuTsp08Yqt33UrNL0ufRSGaldUIgnhJw
PjLKZH3Vsmmy+MRCegLrbk3MeeYx1uDvFby1wqOxHaAO5QgvvGqO9cAMyhFlXxpY
kWNrie1mOBYmIPhPZD7TNSNwLAXLbxkrmLJ8SiZ0RX8E2gWCKMH/ErUGGK5bID3R
faduzOMGiwID22GcqHSUpabujzfmJoWRVtjJgis3oKJiU6KHC6WphAXu+WSuwb8c
3wMpw5d1YpRuaHsJdIWbgZiIv+1feyw7TUEPJTIH8en9WHnYkyCDhIzvWtDrq/Nn
SNvx8Vag2tA7SJIcwWncVXPGvT45UfrJPsSJmhqm9sMP82KXbDnh29b56URcNVlB
h5EXSTuLe6D+nE4Cbvxgiq3lb8H70XTOh2lU97/LsV20vSeteUSQOMCT7Chfp4Bw
ALglhYgRBVcQqGZgN4mYt6UDH0+gdNZqZNJpcPVVdHaw2YnKaNCrqQzkbNnypW9s
HTfBNPk9CMYojIOhVZ2SN/beYiUl+dUiADRWIfeVJcD7KWAahZtxqXqFlXYENayt
iCuiEaQgf6wjiu2r7PsKYT2+CfvSzLldoqRGUclQ3E2kVDHvxU8eFkPTMxw+1whi
iljlS01xGylS9YexzXc7UqTWYjtFxPr7B9G48kHsaFTpPfqDBPQsAeifWhk2p9YH
xZ+eu9TkBtQzeX1l9KBL4bYLmJ2836J6vkIDGdkE8eA5evKPPk9OU1fK2Dhq+rl3
KPxIr+umaYd/ruOgcNZ4YIg58aVkTMRaJuf1M+OqCW2gGuzfOZ2Vef/18Mn1S9H2
9fUU1+/Tsf6oZZn8xjO7qGbYLdNyAuZcO8qCPUu7d7FvhUvYK0vewdoUl2D+DZm2
34n+Y2lZ6H7gvi5UmryC/jvU18RKeV1p0RBNHYjtAZsFgSOhiNHfkRMsz3moXkkj
hzHDkr5JcSNtkv2hfobWKwuDi1VXAchFKNH12xKuKw7lFvSgjQs63FbwbecEmx3Z
kikaPZtFScXMfVn9zfcnD8KSSER/no4FzsSdHtnMcwYCBZha93oJNj6LHWIVG/pi
jJIF8drMtEnkNZdNI9UFrLcdfm2VmQc6S6QJ79Nlq6d/zeDxA0WvI7p3ygeCXD+e
gy9mx1sL+hh4/ZhlJHDP2EPM3Qgk4BmG2XEh84jNbWetVRPCQfVlpHtOr9EQYlv4
MAnaPVKnSJNsPacNGQ4ulZqwk7XcDLrhgG+zKxxqG0mTu8D6JllZT/6ige0GhyEc
FzFC4hqDl0aOdsHMqQt6k+5TlspFFhvoX4emCm6Swlol0mOymXcgdcvtEIbT/wel
cI0o5CdR0r96sAts4I2id7bHaTplQGYBFQMZ/A/JInhW/jyEjUnqGdvx7yRWrxfl
Vi3N6gX0hYBb2e5DX3XP1Y3FopNr/xMPUF9FqP4QzvXIg4YS1Bh5qZlZnSTzRol6
u59mmTiH976H6lhLicMEhcN+wFo0Ak1pJRJOcG2Q+lwczod7tqtDudkxQSSho513
O5ndxWfCRpX2BaQFVDS6PKZS4t/o3D5txSTtom8ZcoVwb0ZwfQ2XOXRGZfxn44JX
u6gQ42llMTCq9SeZYsdZWeRBsuwvmivnVpnlRmHpfpDXFHCzmZfki4jvoQ9+KvEh
nkzdeQ7slVg8zxDEX+Si4qX2st3ezGBVypNGm9iMux9ffoAXFmygA/tXDYjXh9xD
aXz0zpCg132JXAMg04V+OUdxdi+74jtjdbH8Psx0rCtmflHHiK/iUA2DeWYA3/iC
Iy5daSAgCEsLg+JUrIhBVrWQkQL1ANuJxELSr3ZyInKvFTgl4mZr9XzJNzbYS1vY
KCjWTNh8HvD3tqc1imBKnggn7Siq/Gh6czANRneuH23W0u8bE3TiYr4ia1hLkJjJ
`protect END_PROTECTED
