`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixceEu739Fx/BvZZ94r8M0Mkfonp4L48x2BPsw3WNUKHSfCvbTdmc/P5dZDdrVY5
y0gBgJrdlcM+xOF9cEcEnzjAu3WpyonSJwkwQcrs1hpzHcLoEWSUrfCrkg1KIv7s
APG11R0SUKpXJrIN3PHQ5UI0nQWLO/rgMsQBCofBBbCpB78TKxlZfyMnsROnPsCJ
fjkjzmB2L8yUGrqob8XI3YhGtidtoIFrwoK/jZvAUauWu+fSgUfP0f/8KF90uqoM
InjlLLi6jmjSWyHCc3E+gMXLLY3qhksrPbGssVrGH1RXYvmXQtji2VaoCjDOihm3
wOdgrX+wxe9u8zuld7XSIsg6pQuNorcs9rC4Kmf2k3S4be89Nw3Kh6MbVPze96lL
10i7M0+OCXDv8dmKKStPJyzkQEUWELIxj3SvS95c48U9yKo48BmipQWzfqhcO84G
5yqbGTIQFysLGAt5OB6xK5IkL+413QG4bfGfwHp1ZLV/e0KZL54tXlUbTWla1c56
QXvzypvPtVby5r9Twa3ZgFxLqRIbNN2EJYHrvTflvw1ldCBI7AACtd2A869BEzZ4
R+7DNvVKdUyiKnr1srU08wcIgn6YpJ1jwW4uLi1JeuYdErsaIrR2R5eTS/F1/lJd
6GrKqo3DBGcD18Lgg/xH6ND4Y2MjoSZZcxCtsI5puWjC7g7zhl7gT6aGC27h/DSI
GPr0i6foerF3YQ1Zw7dnYa+PAZQ6ldi8724NYfv4kjDNWK5AIYn0BVnbN2dL0tX/
`protect END_PROTECTED
