`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l95o9ADr8U9oaAMQTzst7Lu6PxeIfelTvuvpsMWa4+Jjfz8AUv0EOvXOvuQvWujQ
j0AdJhUMev3OMkd0XnhzN2lQNvweZqsEZOoVCzL8LsdSntDCMLaSct39mDfaEt8+
VbYMsnBdsOXrjT6npNQa0qvrKFNv6jRQRBwVKonqpYXVFf9gC9sXb8Hx/yfYsOoi
3b9L7lM53Zio+GELBLPn2SavPsRBdZmqg+sSf5ipXJkPsI9BpH6koN9pOhD8R7EI
OqqeDPDaw+MoTY1gc2isQggK74zvIM4KoANOnRTeprM=
`protect END_PROTECTED
