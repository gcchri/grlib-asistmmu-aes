`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fo9Zx0DNBgWcTIGQuVLWFRkCDWjpEm6yXunsevJ0wxzcorHOIkdSIiUv7zYShQzB
wJbIAjX3MieRGZEh2qAIaK2ZK6wEM+6Oq+mUt1ufEwbRPDaXEaZ03KYHBzG+mmnV
JMICYU8TpfwDRKE/+OF1w7Cqy9ayKg+Aoo8yuAOeqqEDV4U28pIgVps8y5jixX8w
bB+wf7aZQ0vgKi0XU6MY4KiyrlZ/aAz2kdnCCF6ZAwfYp6kNW6RFO3vs4qsnoqfV
GOXm8PmXrYPO+732dprD8WVbLOPRq2tcz7/9S//CeOtVgE4BgA61XJh4Pnb81h95
urC7w0si2jrNoOidXKHypCCowMuaEbhR/y0BQieY8DBqH/0JigWtBANVi6Zy+Piu
59yjsxranxTojXPb5Utl48kERMBnY1VoN/72Ktb+Fl74mRyLdZOzWvlL5Bf52/0N
`protect END_PROTECTED
