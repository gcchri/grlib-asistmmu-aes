`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHJAW2TIRHoDWu4rGaJfwPThKFY+iDXzQXXm1LR55BJtgBKW+dky41XV3G1iBRV2
iNQ/ptejLmGpFr3ZZpUEAWc+1ADTXZYE7YIymvLvB8HbqiPs8ZsQTTe3sEa2ZRiS
Jj67PxUxYKTclwGmfgJKNOR2FxUbb5ss0RUfm7K20Q0pmjo+B50bzEjkxQyTjxJI
Yu1m1Dq3w31E32HNmfkiopXEr9y3L4FoIdL0Dlu6eG62Cqp6Dc0cC0IG8xux1k6T
UbFHhS95GsACwT+mvopyiC8HLaIKP2J+E1j7R9CLSl4MD5WhkMiT47Ad0HLEyAl7
998mRseTHbwXR7GJQVZ03dNcBA/YmQMTi80PbIwWqeoVUL0lGsKPs5JqbjJNi1ey
GquN3jgwVRurHbrC+f8uY++MWuGG+eO+41no8/PS8kY=
`protect END_PROTECTED
