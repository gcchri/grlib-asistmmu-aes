`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+jQVo9s0+YT9lN9jWAEHwFBEcGm7h8gW6Mvqtfpr+dTDRGvb+0FrPFdxje/zHd+6
UT995j0896hsbXjfhkpwLpdh1VKRJ/RttZ8ksG0iIJbNWjMRfawFZir8xYVlzwvQ
1q0HjMgsqjZ5CpYg8+GwDOUFZa4rHPqrgvgSxcZdZnSOaxWRBpgBLBkk+us/EpRv
XKueXG3ZNXhe+FhFgnRwbLGwJyZua2ORRjqkSmmn2osIFLXZrbwQZOPhKDs53c4K
yz90TAbBeDvg2otpRGHsFKsOtbqWVAFzgB36m+FWxDnxPX8vWwzSQrdUb14cFB3X
ChmGq3jl/J/NK0M02ZPYdCXYjD1MQfvknTgeA7kbXnDZf/tPWZQa9YwQf4AgFlg+
vbkIrfF1R+91e0WA+GCASnEIq68ENZgOAZpPoASecAJ9Mn7eKcal41eGXMeWowau
dUOKwMF3B4LWd1oPVIhMfZahGakwo+5w4sVVq9W6My2O16z5ezsTUewl/aOiFIsG
T34P3ffQtyHg8SnohznENQUzplH+2jK3m8ESAeOcOwPAJBQnmIJIRpQX81jUKOqU
CIiTjtouh+rfVd62FeBFQSCR14rq2omat4ecQUOtwusZg1AYEMGGOKAJ70Lu2NP7
Zj93Uy2BKvyyS9p9WXXIVA==
`protect END_PROTECTED
