`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nLk37InyDMaJqKMANOoVqTriRpYEql9TW2vGZybrVxb6D4g+87aWKlzAZnyZWWX
XnEdM2iTtprpvHnPPQJGYSLvWQeG+B5TAYHOhTMLTszKAFzE68LWgMtLjT/KsfZD
6g7gz2ICQFRr/DQzZlvVJWGTv21uF3uGbIfNuVfKwVBcBXG+CS6nRYdpgKARMu2G
wy+Zp8Mx6tZ9XiwjPd01sVqgCpCqTwSCPwyhOWioujDD2zE0ihUTFe3Egkj7mit+
U6F/1KQxdrvt8iy/3fwtqqYv7TLbBe/tZjlwcvt8Wi//twY6IWytIl9HWQZaQQjs
RgqaC+EcHv+HB2DnLiA9DQhVrkTZpMemGJhflWVjER4EDeBODHIZuHg0V3n9bwVA
N2jRrIGmw3EtTx8KWKPPgoRk218aBcDYToMSMmRfloHYT9MOQW1gfkGW8C4Nj6rv
zEoAGfx7k5PoNuLCKqQsG8jlrxT9D+cLQCfpw75uguTAlec0rdDfYsmPTuW1t0bS
PRlER+ro6xnWJXKEVh0903FGnR2HzTHUoL6Mk2GYcVdb4a6evICVZqGPcp23uz64
Y4IfaTF/rX0FKpHD428g5fRj8xTeZ8cr3cEeBiLIYuWThgt0ntRWKvaO6fIaCYwi
AHy57ssIeOPy3Wp/e1IsQj1NWP7Penykww8V/arudk1+e0+x3DR6MDbTSbhZvgPL
OWuFRUE7sZ25HBKO7uhGDQ==
`protect END_PROTECTED
