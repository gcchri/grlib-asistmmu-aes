`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmQfFiEoZuTGtVahy0+SEWdDAf/pYhtvqCq6St6ad3TCJnrKeSHUgdG+3ita52Lc
MTcKtGIxdt5sXDvErngBH4PDwmxRVnnvvgZLj/Nw4GU2d+ojyS7Q2r6XF+OvaD3G
nUldIpR9FDBOvA4kLdORiKBOgIyUeoKdn0EwSb5er7UW0DXe45LiPU8NeK2jf2pD
S3jbwjdSpJNbApMxjl1v78xvhFRWIFRrdobDspaK8dO89a9K8je6pLJEwfr1pDOr
2BbrO/DtCoScRDCV4dB7HC7f8XR71cSrOQsVeUYxwEdn6Im8VwkZ27Z891LKc1Y+
8XdLqVHeY6JNs8lwBN2tanlqOGywe1odhIN/g6iOL16GenfF5FJ5TD54popmY/9o
4/FU3Q8OPnxh6W+8Dbf7Mx7TWuGmpFNTFqe68GMsjdLOzgn6+BTUZ/gWJ/Xcajdw
BGQ7B43+oQuQb1SN6ybABLdkQEnwq4YYP/q8g+9yXv0=
`protect END_PROTECTED
