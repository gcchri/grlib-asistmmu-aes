`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M/84xaoCRthlTRGQZKUntQxvCyEh6UHHyFBfKN0YUQaBzpj/POeQNwYbNYrQasNg
bvoqaVpH4O3msqshA1+SAVbdMQhDwQH8sKvzhVfBnIxFxYLUNgHkGPYD8sr5DtWW
v9hGX/DVfzzsZ4kQY6idG4LEE4Uo6Xg+N5ycACK9PamQviX8fO8gP7yzSqmH8nvj
ymR18JmzqwtFMtDbridpQ0qfTDHesDZlZ1Ym4iT1vHoHbndYc4bppQJ/9wx4OLbo
8ykblckfmvzBuhtJlUktvqEmelzaQI1tZePFvoiYJqWqQfazTmeDyCLHcjVyB7BV
lGSliLhY1Urys88H8Npj5X3ph5Onsq5gALIkbD3oarl85hoVPyfd26vxjuKeHIdH
vpdN6TGPL0hBACnlaMg8WO4iUGjw2vpGj+bkBAp1ety2zuqo0KqHh1+dT6ETdgtB
xwUKYJ5Biv7oEnn+HPQ1nTeUroKuAziDl5C3CYub4SsxKmuzau8GawLQAzwXRuQY
f91UYlA3tsdRjUM04yVKiPhzPuEkHLYvqvnHFynktWkkouANwF0SYVBfoPBxWcoY
e9rGTFRi7Jt2h17PwBoPqUkZnKOBhq87ltut5UAZ6KAmMDegpfjtpFr6B3OUtPkO
b2crGxk329EYgAU6OFsSe8u0uXQOpJjI7qteU1ikFYsE8qPV5QyTNdtIMztc4DFA
Hz5X6sdEhDY1Q0+JegA7oy2BkE4WeS/n61KqqufeUk0YcmjJjeRwO0qqgZ0I9sBQ
QlwpXZUJ0y3e7Sznoxa8OXjg2LjVuPuCGQeWt0kKeudpIcF4QT4xdIDB5FjEW9Pi
0nkwYpY/dsKyOj/cUBAwnUn0S9xCdvJPabZY1O/mun8/mwbenadeaHnkAk/9i9n7
cTPt4wC3mveemrki90VSmdHblSfMVz70T1XjOcVb9G39WyRCKIz5LXEOIhb/T9p+
o8bsSq5Z85q9AdaI6p4H62pt4CMBipABv2w00Zrke6jt8HNblH1/ljVdxWQTL5mw
GvOV8nH8UgwLDAcLndECp+nWxxDIWX5t8UJRzGHObU4yuFW6aeFRVR8nMhUgDiNa
pcbdq58omhOA/kerxgJPPNn/DdsPxEcyUJ3lot++qsoq4ftKLzklQfckLxeht2Lw
4UN83p5HlpB4Pq+wWFYjeEPzZcEx7CtGlGGI1gnAXOWihnng/N8o2sCHLdxQMM4/
IjsjxST3THnuAuPLY+g3lGZNksPfvIWUGg9L8SaKx5CSuvismFkTpsBbmhTJqUT1
m4Qts8RYaHSuqTEaju+oc7XVOJO6NSIrCnbGHN+v+Zg=
`protect END_PROTECTED
