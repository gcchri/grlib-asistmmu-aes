`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EuafZZueT/LGIPJRsJzocn1wsZJKGHrDQ0wz/i6/Lgp10/Po6wFZSrWiIfHunITK
WTt1dkAUxsthN8i9ooBO8qMsGQqRZil7UtmjmlC0ndgU8C/wTrlbjp/1QZqg4aJj
psXP4hWw0C1yHRV5hbfAQZDxx7OvLSeN1zOpSj5/T+1ZJgI3r9mLv/TS+JcUtMeW
VJDLKZ1miOTaoLycfowowzQ7pL4XO+5niWqOxnOpomdWGHFJf7qY/5aZHfxjEyX0
GvfCZ7+qOuf6vEovV52q4t1MPzFf2Ih7oNdwJMw/ztZ6GGqKGH7EKlvYBxpJ5TN2
CKEiEvruNreU+JrMbAGaN8YINLQebu5H00aJgQNcLtnCBEtFhtE4tCeo6xFu0oC5
sZeNQd/FDuAuonqy95E3M1Og10OglFDMh2dlncAimR+7cS7MteJ3csmNoFEbRY1T
oL9N578Y7M9896eyPuNYnnKCgF6LZH4l8VC+MAlP0f5QfjZ32YzTYNACCAX8+P5b
dp6KzCTRhSv1yYjqCEoXFin7i2kP0zteWiOTYcOwScdK3zK8zbRasKcyfWf2J2YA
YGLHfAQqVE7RZJEchIk/J9rfqhHLAVQPTVcm8Xk2lveT+6Y6D9320N40gl7xuqVJ
fXEkOCjwrX8cFe2HL9YCNqRipcfwmpZd8P/Ij7V21x4tQecAPdzOCHnqhp3C3mWy
GAZmVZuEBjWe8x2YPv1iwNXamfyOtWpcI7Otnc4f7qUWN7vWDsp1W82vmZVeK7Wi
F9MVGVvyCTx6vO+X3jFYFNczwRGqxPdMordIikhuDww3fDwZfS8JtG1S+ThjhZ0G
W6IEjDt6nRsLe77Y/eiqZHLgLkd2iijVtMu5a6AyMh5Sd6rs9QhxUwScCYGD9UWx
LN9DdOyua+qggogwf7dMZqwZ+2t58KiStfKRNQUbXYuXeLXL0/+9eKb9oekf61+l
GR+tfzmfbmQ1q4fN1jFzNaSRon3XwB+VlzO35Ml400pKiDgPtEZ0mTzPlIOIHfYw
+JR8d15msLhT6Wh2ZuFlKhKI2gs8AV7FYUT3JVpG0JmKseGr88Xz8k8ET1a0J9w1
8o0/czSLmvsi5fbf9PBhvVCfnVZCVRc8k5Vshbp3cjAmQyV1JlC327o6TQ4JwxFB
QvE6K1gIK69i1WaRmX8Axc3na77wwmzmXP8UjIGuWg0MNSxMMipe/k1Dw67LoOxK
4VNX2raScEkCoGNN9Laeu7CCPUxK9wRJ1nAJ2ZmaykJ3wb/VexLwBJ1NO8MJu5Yr
vFSIL5IKVDWPUXhPeCazkd/m+EIUtMsEeJRaMHAOcQXBFvYXLdnCtONDEnceuZXe
dB2hDSGywiec8BDmHrBHJCBhjtPKkgiTEFBEJ212M3HkPAsuSytGmvK6kHW1Kdhi
ky2R1NEiPoh+1/yFWL7t4YWZyYWgWgffNdLXWLNMNAdrR27qrAMB4EKMblnKHYVE
o3SMOFa8klhgC55dymJ/SwjO9nQXxQBq9KQ9gYHctMFAWphNLXRhDOr6AkJVN4td
/FkIVFS1Ub+cilfC2e6I2twkFZVrS3zOHhgx4uRZRAkRV00sib2gwep19LpCKrjM
i4DkhERNiq4j+ly/O2WaD7twVJCuKqFWxzRmAQQubeOe5DoH29AShC1oKsTSBDAk
b5Y6he/CNlcE9MijvA/kr9vb4Xv1Bajt0AZyrguvW7RQQ0ERU3dJQ4gJ0NdI4ndn
zwmiqA7tngoKC+UrqUX9y3k+ICJBZv/yhtQ5ihC5LJZaRQQRSRtEg3GcbVtCLdio
UlpOuAYytRMDvnpf94Si1OwqcE5FWR5ld70T02cAtL5NKWG1e3zFe0d8OlUhnukF
qmdZfvspdpQWue40BOj2aj0KtsJsfup6KW5sAd3her4t4M3tZ4cwToMQa/+KX0Yx
D6rMW7O3NQ9mw/qiCy2QlKMcO9RYzZhk+1FuvvANWVSiBYUQF/4v6X5tDugYsfz6
CB+LKYod6H36oNnDVGXwiv+vKEOCwbc6mijQs45x4tuW12kI4eevB7Ev5jN4FPDc
ThykCfY5o9x5Xa+9PUUOgWL4qmibr3/1+aDC8UB39ktKu4h3g1kaS5uveZxZjWGo
PHbIcwtp3EA6I6CGG2bWqA0xUWgWePardNxUC2GyC0dQqITVfV+OYlkB3h0ihL/V
ME0aVsnIR9GQOXeBUpo02OtSxcEX8dmUqvTEH5Flnzwgy/B7CVcodmagY8t61yrn
mSpeX3jucPZZ5a2vbCnU4Vx8nmKtGSn06/3hqGLFt/J/zp+SdfQ0hFP+CE+oziRm
pspgsER3Abh36cu6oyDDMQTffui9sZbjjv42yl1n2tQVrCjWRfL0Yy2IwNiQfkTE
ByDhJI9W/TJtcv7+rtZ7Ge/VpiOZ4nora8JkbP9UsPoQOILN3ap7MBsx6mBMiJSV
7zcoZWoLhrcyJuWpeY6YkhhS3qzkjMAdb2Xwde40Actv5xKrj8hq6lXO7zdZBQU0
UJbzR6JeyAqVsxuI2kdb2uGdm+IIQHOXz7h6UCKO4bj9VjwRaL+JNnC6QallHxeN
UpglLIpvz9tFyCJIo3zUN3UBoqskEmj7pBAWStemPGwZJdA5mm5sK5dfnnPnN2vH
6cXyCuwkQHjxkeL1PuNiSVGFYRoQjoycgqtNnN7taeOnGY0DGMcMZXtjKbqFzD0Q
LaDQ9+VRI7ZR/pgdcq50Z9Eh8mAdKSWTo349flji3MWiMQPOsbKpF/Z2FlB5O3PZ
ruw8jilpQgw4U4iCf40XEWe9ijurqSZ3b+Eb3uWENJn2iJ8MiIy5TGbJPhUjuYCl
9Da+UXG7Zl3kyX/o/OC+Vekz2VCFYALkVSdUJr5G9xc3YwdqBa4zL7t/otqIBJwU
7xt9hShiqP31sxq0lrGZvbjoiGg8jPz7WInou7Tl34YN+bxSwSvu1J2g49wYmF3C
QX8pL4ON+4CL95zdHe+ggQbb1MOVtLbCE7ajy1bsrg5cMy/+TtLhkcizLNCxX1Ja
kJ+ehbz31FNvxKfTwl/CUHo8JVgBu6mmlKf8aFKEJa3GrquFWaKT+7DzySWXmiEF
ZFZaZdgILNve1fwZZvppXZx+Pv4GDpDnsAIUad4P8bmnUtbTcmjuFLFPGOfTJcRM
HDDo8A1P7T+z5vcPAO8/iWpyURUW4WMT7malgadZRb5pndad3ltBpcVs7EKCWSfb
8g/b1pGXJeX+SrbfxEIUzsN+a5sg0KDf+c2pCrcPoEsHYmy37X0ZLP3cqnZCqCSf
lYucE3+oNA2a0bhUeA8jJjUj56f+eOXysFXcmNeKZW3yOKU8PAoeQRAOwB+y4sE4
8t5vv5UhCTj9tCPkUspbTWgfu6xdHzs4uGfjxEEY1AnG5Jsf4ltdyFByhPtL8Q1Y
CX1Bpza5VU5jdXUhO0AP+/tR6UlrGoNqXH+RwxsK1Fyb73oTGbQlzljoVdal5PAM
`protect END_PROTECTED
