`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FX2yiwAvVQKrMLBDh0zigun3Xj2p/IUdwYcoFLgNHwM6/x3s2FLD4ukDL/gfUIHN
0GPS4zp92B2yHOZ+jz33G/gBPsqVVanamizJsX8XlUME0FKOXYOi3QDg8mcE5b6i
MiPreKQ2qS7TN5BljAkSO3Q6q6PPpohe2yfokOpMmMFnEgaLAh382i9ATn3EYYi9
+B/RGSCVtQZMwu+Lu/HONG+QKXIH3p7L7QdzIyUvHbtc4RTazR7LXv62gUdrH1xZ
N3ScjMPuFcqwyXJSUowN+aK4m9ni9XxKR85/UwFSuUYrrczuP0NiGpo9La2on4uj
9D7lixo99JcKaKvAvETpbN1OzturVJ60t+m6VGgNVLly5866WlqlS/02RriC6v4u
HdpWT6izo6yz1lAqLFJMfXfUutXqXAfLrY9IfGnf2ZZEl37jMxl6nAlvQ4Ub6i/e
cj9QvGWpPEI1Jc8bWhkzs/7wjcTBZ4OgpkPP/jU/vPvss+05298S1U/Hy6l9I3vD
eCwbR+NMAftSE9euZi/paJtuUHM6PieCXmQVBAfc2vgTHXBWuw8GRQG2FQqZgKB2
5mpOO03yw9txFoWgukOqtnmDavUy0ZUKlBVybHOb/N2hu3FR91AJwW1+KTBWP4wh
pcH1tcRvNJOlc6qDvOcBI2xUyuizesqnNGT3Rt6hnnqfoJb3YycQVWJwXD29td1i
AYLA7jmg2HrRH9eqqTVZ2xfuEno2pLNMoaS+DiTJ/ivY5HNmt536D4BM9pKyDNxX
LFrM3JIlz8guBEUaFvY+jo3RunOhhcSVrFh3KuZWuSNsZ6FK3v2PlHyU4xQy9HmA
L2PqHZVocjsKJkZrTWvs9CeX6qcFVnwZ5+AeTXxbU+UdnlTyT6wGou6rn/dmWAmI
bW08QcEALMHQw0ghECtxogi1UaGfjVaUyHyDDDZtPPH4mulqtP+F6Zl6Nvw9ph0m
0s+1Tf5O/V15z7MtKicjLMpT21d7zW546fSRVmmt/4IRpiWBYzy9DUVb0amCeJ/F
1ShSbDRa+zSRENvfBLcA/91X8Phx+A/q3ALJ3iCqEhk3l73GDKK2fTzukeDPOIfD
TbDIX2CtrIdhHGCDMxZht/aWRQ7oSUJ/H/jysb6tbSx2fSbNen30kA+UsAxXjNUa
cfL1kKjRLJKXhDWRw15nRJ2k7Gb6Z9NoLS9E4OE2P0cEIhRsVcT48VwVTBOJD3h5
U8W6bQbOsxtx4IrgSDVPF1GwGEMN+LbB4zzoNz2MxuY=
`protect END_PROTECTED
