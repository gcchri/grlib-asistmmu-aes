`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pjEz00ESZvzcYFrY23nUVI5KzS5iNDhu79hBhTaq4mKNbCdlmE0Rh1GT9rsp30K
/C+uNGbplW37NhNHya0XvPI3DKm5mMZXCmIg0ZnklTmBOdKBq7uYvdR8kAEGPYXW
SHh18gbRzS0lWKGoPYa49kwwzWOyjb+w5ItBFW7Rz+DHxN3bOnZeIM9Sp6IexOAR
GO3XhfdcfkzIx9XBsLfh5SKCh7Nu0jTqgQtogBGZ+JZJRDwQKabcv6imx3lAUKtW
c62hhPGTxB3Y4rp98ZQHLZIHxlf5FaqZiPNT8mG9xTfDDSptpPkVaKtOHwaEBc+V
TXO35fGK1UBvXlUG4AW+Stp5jrvd4PMXpYszJAqXbUcyCtkOrORUPU40rnENwyb4
HXjR9yR0KpzgXkWCXF3pcYM5gLYz6vG3VhRsjWIP/8xvGgZkz5w1CA3hVq4B+6wq
9IQf6yx2OjP8nZltd0z0GU+ufWRJOwu/brdIDQEAmJfE1DLoq9hW/1tY7KFJ0DAo
vDeBou2A5ZLW3ePy8u7ajdujlFkMO5xa7If2+WvFXvYkhVQPZx8YCWIzsI164eSZ
Lh2v9pci+eK9WU0bzyySpnE3PrdpF2E6zODUWJJgRGRMXwpw9QYvBR/wlOrrVyao
T6DIJThOGqkgpCiSfBTHjVS8L8z7yJZDjnh9i+nGuOf0GRK+MHUj1qOEoU40roSc
`protect END_PROTECTED
