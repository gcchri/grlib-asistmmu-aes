`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R53iFbs/ak0hxWZue9HOMJWBfsJHGxIUGRM9PiPSLPRkxJ3hpkARPN4SHbhVmvgk
p/Lo1Bgfd7/sl0FsM6NO2aUXMDQnE6CZq/YAIuscxgwiQvYXkhZjC4gto01FsYG7
4Om1nFBOuiuO9AqyXoN8893DDGMBzs94NJXWwZ64SNY/vfkitiNU3bJDpcxVswIu
miYl6M/QJJUKgyEA3SUrr9DcW/HGkMrJRcSA0rzC6MQDE6j4zkzRP++Q9G/ZzYS3
ZnLveN8gkcJhnmpUh1+2ZFWQwmc6v6ySE9WNuJwVCLgs2KMS8KulKhJ/9wuXTY2D
QiVNh3e+xbd4T1nmukB9VjXCPv7pX2GZ54vmQ/LxqsXDhMylqxuApDFcB8M0uqAQ
SuFHltajzWkpbSB3mGfkWWNWyBzWK5mkp9r5kEMZpw5b1ITtPmHO4VULAkEQrjET
aGKuym+ltuKn1jH7fXH3dkrMg1uxlQFRcIoL9sKlD1gczhc3RsrWOtTC5GG9Fx7h
Qww3myOFRFFoU+tiv5OCLpBvXfTbxDgnRwO+dxFlV62fQ8uxSSPC5EYxdmyXGq8+
z3jvv4MTRQlAE7dn25hHeFcWWrN2wgvNWfAGi4QGRO9KiwphB6xu8SyWwNA9FZRu
ZynNHQ+ho1lj3EBKP6xD5b8teKAzgCu5RsTolZZWgnZwFdeJDxOnane/QyAtUh4j
GjQFguKzOnsGGcJhcn467CSLgjXvXiPA4QE6h40LclwT5wKtYzQAYyOBc8Xn3y7p
fVeYYYn2QWIAoTV1Gl8+wLbKoWzIvk8eFMMmVJATeChs5VRwuyrxLEM7a+L9p9B6
3x+bafwGJ62es3sOT/xbScaSta16w0CieeiWs7E6aGzyYsFpMROHrPmqB7enhBr4
i0Mv79/ekQESK5oOJOzOsiUSAcnAD9pBKQzVN83Ff73P2PcL7dScB3SpwxbozZAu
glkjealicNanFSQId2+V6vYlSiXVa/u33Vp5MqTCYasqPvFyMkuDXfwKVgxJjVgC
AgNOOVMke/R31h4ok2criE1TuaO3SBvI07EKh87vhwkfBnnN+Yv5enhpX6EIlBLd
ZQYiiT2V8IkOaHRs1q2RDg==
`protect END_PROTECTED
