`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RGoZkrrAcFF67Md7qX4gs6J6G1Z40gqAhdbtlMjUYTAdALDRkhhsrK+Loo491Pv
FldLukPQNldqVDclkSkO0I703L1cOcYd7EVAUO4powvayW8hmlI9mmuff3SsHjNh
zf5OXrKoLAU8vM4/99N6A5ub1tEJS5ZRlos3+9UR8Sl96l3jrWMzpOWTBUdLsoxo
LudSVliFiHPAvhixnGOKBVNs9R+JGEa4vIL5QRos9gA/NWjVD7JHfpCVW/pgllbj
I/vbq5b995m+JMWxtOpgIsBuKUFeZOdjX4rs2ZQbTnZo1hqIeGE2r5wJ+0zJoKZ6
eMpJAPN2NK2KUg0aXCBOfMaw/Xn9VkHES+j2x5R0wATjidBW5iTf3yxGdfdWmeIZ
ydB95uQTpB9SctjQ2zA+s0lkqcR78JwfgMzqAWlCrJ2P6ct0iFwc3NAVZOyi8Kry
RXyEsOX4YkdcsFcnAzv9y4xYDacfzbgFBIHxBdKWGkM96tP2Xz7FwwRzy0cwINzf
vFSD4fcqr+9FTgjRXBvJ/KYmWqlEIKZaXnSGVUc0ZDG1cd6GpEm+ij4i4vYQ6fZ5
CTXcC1ho1+9oeJlk5Bp0FanZQh/qwtI9zhKE6bp14gyLPlSIbgOGlav6ltTqn908
PU1TvsSQ1qP5KgLwCq6MGsT/ZyR8l0ys810b74lfZcscotoT4hfqTf2ZrqXIo47P
NUsn333A7gLCmTkiYhkJCALsYH/rU+Ac97ALPRIi7+vSOFkBpKZupQ6MlTCWyDtz
TR+9vr6gCO06PDFfgaRHV/ihIMGBuIZWHg1yxkg5CF0gi9aoiDyI2vZHv7xIjDO5
HSkzPIrLmJNxRbTGqL+/nnCYXJW6Ef6d2RJC6QAHYSYDn0s5Kf4+F77b3sr+XwZB
xzaklb3LzcT7PCJ+q8wa40BDD8EF+ympUtngFxhNZempPiXbYmpmb0yvPpBTYVq7
ACDjz445sXyWbIpFob07vwMwyrj58l+MnsIyrEPjvFswJaan9cWl8aHzlaP2VmVy
BKY+ZMR69qzGcGeNVHp0JLVQBGpO8ojHyO+G7h2EaPXaqDm0KIU1sYohlIX7aJf0
KoETJ1ITPNJIRcpFNgsXCo0gHSZdIbU2VmjUmhG8VnDFI63So17JzVfl1elXCAUr
/b1w/AVGfGuXM+RC1yqbFVAO/p/E1K8//Sbym2Yh+Izk0g29cnC4jsbTGVET3mJ7
YZ6tJqYRoy4v5nvvIh4il9MTmVo3XIZpqHcGfpyTUr7XwGBt5DXyAenPNlX1agoi
BLKRE7RI70XuHWSKKgkMGF+THDNU3kADGz1BZXJwAG3c+sYeera/mgFVHgj7v4ZX
6U3himEqFrmrAADGVvVT3PXuP5xrvZPQd6ZHonRlYl8q0/By38EdFu4+/27vJxJI
fFVwPW/tPtaWo3xdoNfz5E8jh+vn91/qXYRbX7+SRuCE7/PTjx/xnIPKQe/NR3hE
vNz2uy3NJI+pwnobPlkPDnOigKRQEH6zuJ4ZfOXDwIAaERCxy92ASRq5dLuM5qqT
UoJWa8YNHtiMEcN5E4uuBPXhoymifJ9PddJkJ6LC56sRVti/krywuVlfIXVJhWaG
UKdM74TTxm3Gh4QhlzPkHXve5/LJSsDAbETkWAUvqaCEwGB1KE/FieH/9YjWgjUZ
M4B2DF1V7zLr9TntoxXBgRJgn/B35F+ck9N7auB4E2uQQENx2BNl0hGx1ZMawJ0u
3grbX16NpTnbBuU4C1i4tjq8YpJlIV9J4Yn98XarNNJk/7oajrxvKS5g3ZeL+txJ
ZPHtI6YQcCF3J/V2eBvx+JKDxJKudOox/bfV7xYReXgZC0FtQ1LlRyPLHXsp5ut5
PPAuqARAiQkKC1YgROxC9bRVEd+/1RDQI8UcEfuiVHQis/5IvaKbzElRxGzxHOYz
NAK1sxVh3gXe1zqbMH86wLB1hvqHTCKxbcewLMc3SsQ+CE/VlE1r0zz/c1eMGxnh
oO5mPdlaHP3dEe/+T2bHKpwoI7o5DH9ym+8sGELR0A21pLTeIyLP1XTQVARGRqgV
2Uw6357AMwMao1GlE09373NVoCCH3bnb+fBPE8M6MhBpjfcgLg++DD7jLS1gQe4c
`protect END_PROTECTED
