`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vU2PGBZPI4m/ex5o7Y7VIAeHfRhrorbr345RGdrGZwNMfWQFqkCLIs9TfpZHM2z
Z3wn+wqCiIU8RDQuyWFqiPgwWog52Fu/WNIUPGdSXoUrxQoLKBTTLXmcPSRbsMc3
t7AzBxf28OEctvXwgDeTNoqLln0KGqrjv8W8iAnrvdVjccIoORvmxnZIqL70TYyl
TpF4SbM285JVKHAH0xDfRNXnj/jxU18FB8xgmvhxENS+X0SMf3A8FDtQeZaCo294
ZhAW/5XQN0X7c55kCg0kT4nlYWMMyC8vyshGFiNN6XaVv0Woza+4nCzw1SUnhKje
ywiBLKEGU3+0XbEePpYHWvNrVYwIXKktqBvP6j+5HsK/e2SGxep2sBhQjrQY79m2
jQCZbUT8kdNfuyeYZzpR5R3/XpeG17GdZDbulCzBy4rqJS4L7bITOfuYqQaSlDMt
gw5vukrol6gACtm1gWZvCfSLT9H3Jadf8vwor3feH/pSsRuK1OSinZMG342ZRf55
qhe9TOIQJq6ssjDeh6YSCBvV6EdtIXJHbWtE010CIRa1BSdjN+C72prDCABFsOj2
yjzmahJn2GSs52FvUUoiaxtR7RB9/QqqbBD0NwDELzDbrAluKIzPW1I06ZJNUgJJ
U0AkimlMQQYGmsUjQlCxgs5JQhN8awbT/tBJuYIgXqWBqJK9pRXtvBnBIkWANbZr
M3icKxm6e3ZRTeopdR3wJXNHRKZ6mS7qpNkw5a7P6GDMhpvNlTOzi41EunSaZ/rU
sAuQm7u737pc8wJxSxfog6Y69Dv5EMxCmaJ7uzTaSw4cK/PKSFrTdXTDTiAXMo/G
2Lb6zjANf7gAzcXadLTbtEvhLmoFkan0T+x2ENWB4M4tngqQpb/1hZa15EiCbhp9
GpriFum5bK3netiAqGgRvzSSUoic2XwmUrbqjzLEJQGCW8ay/8piZu/Ch524p43X
0Rpe9Gpbd1TVRRlKkp58jheht+Crik+EX/UnCr457wVXv5uH7ZuzfUxtv/LBTMli
k1KF4OFhilyIEex//N9Xevm4h54CXbG1zzGxmY1G/gJYVIoQ1Wgx0WkSTiY7wydi
1xlITotUbdjTfPD+hwK3qK5DWlKmXqdhV+sqOds1OYnB7KP9BAbAowNvC9LdD6VE
iqqq7WfK6azc+4GOVE/SYADqev/2k2nCCMPmW3p3hbOUKaavsUHNUP/DoIIiOuvI
amr6j4bFOYjRagW4TknXm2SGv3i9/P5KnuoQ+iMkwm4MrFenvnxn9ZHFrIWVo7zt
u5bYlunImty3p5ZEoTn1LZtDBAXLNDAvONPug9QUIf6gLXmv1w1Ha0cNquJKch2a
dXn0Y8Z8bW/29oW5GIfmMcDPtrCxCChujFdavQH7s5zFHLVX1LjeAaSIv5bBE5g0
FnuslnMXEaORtvnFMiTUFkC8P8C38zaDck7ZTW291GjBnaX7XUCzXImeUysE22dG
4spIIzhc7rjNkFK0/vjeuu/WPceK9U1WmeTx4tNnaMX5HHIZlRR8QqWvwNWIxzB4
oPo1LSnELuhwFm/JLxwhJm8u9Ft37QXQJH+GB2PoGsVFafpKbMcq39hnCOrX/Pvm
wX5yXvapcY95bNfm8X1RWrCiQDC1BdFHTEwz7LfGd/Q=
`protect END_PROTECTED
