`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahWWJn1lFsFJylB5f4X0kJQ78muxPFacAGVz/LVJtCRoBhsQb9qc05wSUppoFvZe
ECH+vRVBUCaTUOy61aTQrV77dxAv5KJT8UZUQcpAn5XMCCecZKF25KqpvJUGy8ag
bOwYLZxPs6faVOxjoCBm1tojxLPuyIB+MUMy8FlLlAOtmcRjqCWbN1oPYBVbDPkv
TDqH41Voys1chUsLuz1YpvHzcTlZKZV1l78KwWm1aEV3cxmMlJtQscHCV9QWv2lh
j7jOAZVKvQyo01+UNnjNcMcF87+D/yRlBz5O9QIklYffs0PlluoM3GejJRydGbXf
bqUW76jJB09WvauXZDWPpjmmVZ1494cptHuZpxKZE6386S6mm2f2QyYyRk8/WcI/
2vpD3gv1b5wUq+VfuRmgF+EtAAD/UiJHgAQUvH6xQFPqyerwZ7J42xfBUkQ0YBqa
a4MrXUKQIrIOIJrw+5iBS2JNI/uhDmvzOV9eAJDCv5237FQCqEBRpEJpXAvmjsEi
5oxigeIeIz1M5/kqSDZbY9RSV+cjASu71VnjuQ61IeufTd8k/86zWffBmBU9Mzhm
J5MQpenNhL0ItxbVT/Jfct0qdekv8BOH2G6FEjtaqsK5k7Q1JwgtgI16qI2PRFu0
fxt/wy8ZxcYmkSUZyusF1a9/aNb1nMnY/tybp5pGUcapAP32fu6088T0CAKF4JJM
fwOk3p/muxBmqWw7p/uaUZAsQbIWHfmdowtHId1CuK48AZWcpASzSLM8Z56Dsw+F
G6Xk/hVoTkhhmIB/dmmY+wTPpFGrfqrLv+HWFnPRh7HN+djZna214MAuJnrxYxzK
rzZoT/McrYgXKIKtxO8s7S+Mfxx5AjN9XWCtX+3301jyIw6hvFsiJWGFuEjGech2
oGaDDQj47GkObfYrbrshPU/espbXTUI8RiLE5kywOH8=
`protect END_PROTECTED
