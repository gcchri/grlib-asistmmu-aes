`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tqdwqI0JWy9vVYwGevWIrKDkdBDnDmEO9dK/Sdw8K5EO/2Cg+BNE+CXVewJLMjOk
imZ+k7zFQh4P1TYfLdSolvFRrlUwBHgdmsyqy5ttMIKwvSLxgM6tp/Ou3rOdByfd
cP5GU/vYpX6GQ6lDPVXWc/FOFNY7/UaB48UbpLrrcUNbuYWLveKdM9jqlInlKhHa
Zo8KvqDlogUMiv9v4gi9zfMevOrogX7Q/JUpwcLZ8GKO8xnCrL10BKvxbgiDIWTC
hcHReCvhbRZPXMCSO7U76U76YD1HhdAtkpjzWIidarlzSimOk8BrVSYX39jx8eBa
HGSWsTDfms0OZkyi0r0CFt2Zg/BEYpZSHtj5QZL0Fevq4/zdP1lEycQV5HUNM35w
MxDsoTva8vuw/6LC9UET3QQqptoLNojNeGGHf7vtWvWw6ZTN024Ebo119oYBCn4t
OWpOP208mhyWfLQicxAg+RAElP4bgdZwTgME/doUGZZ7Li2RbkI3Vm1W0ydHlyI+
2RBfiVfnRKgbRCo0hcgp9n2/+l0Q7NcXIUZtgls0sy1a0rb85UVKf5t0JTg2RvRF
2ymIcvZ60vXZYPemBSgWZA==
`protect END_PROTECTED
