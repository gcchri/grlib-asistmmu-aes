`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XnaSz8NnA3PtPZHzRkFym5BiuFT8XZuqOTdux1GZQYtQjqwThgSyp/USoF/UaChL
/KBHaD18Yld8E2wtpSuuYYZGw/wq1C6LhjFCCYuB+RzzHtsFcRVUTV59Bi1DpPuq
PQ35zUEgStHaJyWnReVZ6qTZSVoZcacGxMq/iMh3whN95GhVo+P3Le9S+jWW6ElJ
qvd/b8aRwuh6BmROrjjgkRKLIj6a5I7yTMePNYaZCn2fRswYVjHMuz6Iz1ehCkdl
kT5Alqq5IDd5s7dJCIdZnOKzR8dm0prBBCDRn0+IWNDbU51DAO+kL5GSiPzVhd3y
GDahLQhPSeofymdyaM7gPydGwan8yN0wwnUMczXbz4wj+tymGt513oewUI/nx2Nn
IASus7DlRB9GUrVY649qP+sMLzB6neSLYUi5QGkaiEJ9q7USMlQqqztXDnr86J9m
n0qf6YTu9JjFr3OhvwKhwMbcyM3B19L0cNMi1g1OsVg=
`protect END_PROTECTED
