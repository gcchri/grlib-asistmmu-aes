`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvx2EjHUnIqTp7xSvZMJLg5BX153L1b2V33YaTF+dxubaqbYepq8qeYmR/TkohdA
tyIqiTa07qBxUo87LaOoWzy1ZUkKnPzRTaXw1eymmFG68GUDX+611nHnKxs/0Qy1
K9DWBbwF3BIL1VyXuzvIVsSaHnRfU0/uKBm2tJkDQzVWLImmu813n3KXPywn23+B
hHQxxJ+M0l2jpLh2PPUKnw7qDigRBImPrXFdFdJxqH5O2jdbsRPDM11hyaIiMMYE
fgNXCX+eEAiYgkdtXLd42/zvc8fciw7G55OQ7Cun1d+4wsi+KYdEGIOimlCq9ZxX
AfCWRM0YLj1VhmiLdlI4Gw==
`protect END_PROTECTED
