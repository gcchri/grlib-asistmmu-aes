`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HwzGHwpJRfDfjrNHfZDbob/enFLiW7UwX/rxeSYXrV6u0tA3H8ayUjnu7gfVEang
V36sWeiXNVzE0fpSfKD8INA9uyMwY3mPReBXSkY6j93jIpAX7INpg9Cd+3+5WdpP
b+atM0sKrlQFaWReMSA5dBOgaXcc6eLUWXVsMSUm1AGoIr6/QAhIbK/g1899FBgT
HP/aSukt4OSuppI2fxon7qDasWIphaMs+CbDnG7cDg7enxOQkofnp42kFziCepPt
M6dCHfG052dBx//+8GGoDF/SiUU3pxFBS/1N1MZ8APKgfJfvHJtW8v6Hu8K27t2v
fA+MZhOVea9q12uYpy50R/ghhuWZKgfcyBxx8OsKAIFrtXI6xvvOr9OTtNn97/nN
YUpjFsI+nuidnjOULp6sPTisGLX2aRRERk69u71CP9eJ9E8xMKPaoiDCbNLhxJye
`protect END_PROTECTED
