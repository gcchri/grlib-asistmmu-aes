`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yl6H/bX3U6g/GeegiNWWcQs90Hk7SwFLh4PwTX6ahmNyaiL23261CHm5ptjh0Sde
zGacXcSRPa1JmjYx+ceOmwaoIMOgHAhFTV7hoF89R2jRNpK9PQZOgpwd1DsphBTU
vf3I8LhnMuRkDseXY+Olp4v39EyAvOuvEPC8C+2qtn3VrxguQqeMizN4l1Fe2XWf
lj0qiMT+LprXqkpTejiOPAbv3ayuLwz/E0MhcGnp+WLyfjvsHmitB5PA8yo143pp
IQhaT3A7/BORZbMLJfIfk9j92WMFsli6Cx1DzIvWftwiYk0T5NNWuU92HC7W/USU
WrfqMNNMeIrd2fpqQ91EPUnaZJeVdl9kQCkCtTICBnqU+YjHocHf4gmRnGvFfp6V
IdpqvVrzjZAMRhvu5v1vSEmrlHpsTHqCdX+s4wdOEo9lij6AaeKWw//+E0EMHe8e
1Q5kyVFH+OBcamlNEpWxhaUUF7DmjFNvaJssQb9fjt3kKUgWB0uKf6l0OTAXeX9M
`protect END_PROTECTED
