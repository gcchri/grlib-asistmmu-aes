`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zglijbJ7XelgBJy4YGjtv3kodt5jhOmt36nZ5+gloP1OBpZlwpORyP5UvbaSbqJt
FECyx9sKvw3rWG8VM+IkHLAOGp3r9PlvlrJZJo3vxhDF4BDdezGsmxLLSLUHPY0v
6XzEPgyGg8g9VwaGZID9PL0BuhsQvpujCTK33JHE1H+6UmXdyxNgGIFFAyTL7ojE
r37evcioPQilkn9Exvt/N8i7PEYOTr6/ukKppwxoXI3GS3h4s5hdUhoKPfB4ustj
GTBddVvOZzg+XW39DkU7y4zysCJhwPEShtq4rY0uUHtmr3snJnBdilRkZQdeiNPA
W6AudbPf2yjkLOs4YSNkuNUp64uRGSnEalzBUCRkUoWSeCfXxIYKrJAVDZt66UdE
gD+PcdyrW2RYoBFRCksx2j/NBIbl7IZXjB/5OWpOK2J+brjRBHqQPMOyeCEq2NG9
`protect END_PROTECTED
