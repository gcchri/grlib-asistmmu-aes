`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qgR1NpHwMNwXp+6OqT/y8EQn+JXOLd6+cbFcVXEhgZB4naqVSRyEgy/zmxd+5USb
16xlw4vV10WnKNcCcjd8laAgg42cey6cTmXdzLt3+kraudyFQ2hMjaXKDZ72dkbS
3vY7xzO/Y64t1YfodGjDiLHDNKtHmyaYjLo84Xcqbt6o4t7P1HOiqxoLwy8XD3yQ
DtiR1nK+ydMLmlYO2CltP22dDtm4PRun/RWz0GX+GbaXP29bZmw3tV5qVjIWbQEE
k1fqGMxbwljYPjrxVOOX8A==
`protect END_PROTECTED
