`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6aNTxI10IRv/uYpS85b/v/yeQQ5LobjuB4wZJgTmDcIPzF1Rs5yAC1za6KqjVruB
Wq+tJOXuHZk8A+QeB8AuKVypZrmj5Fq0d6fldneC6Hrn5DnW5MGHcpc9YenmfrIX
lgqUUvA0Eo+Z7xitciASruAsjoZjl+q5/3EIQnwcGSw+uY828fKp31rTfH7v60uN
ThVLqirYs4BGGEpjIfDfXYyKvoi5Kdoa3UnE3HVk6DMsDdlxvd5ZwQYJNmLWdZnm
R/cSidhJT9WIRBdEM4HYGD7e8VHIGZHUrcxBuT9qBzdRDQwYw5n8P1q417dGchEI
Irto6WpB7xp932z7ekI8CyG5VP0YVACQmo1bGMHwlJ8SblzwV20wlTyEn7lKBMiQ
dyuXVpOfIE2FxV4wV6yeaABoP3ekCPfr7eASY17eo3G42s1fjv5xw2VFs7L/A4Cu
pX7q+St+NLRK8/6skxuRhgx+uYyE5vcKYZnQf5iUFXFQB35uIPX8NnW3AXtaTQg7
`protect END_PROTECTED
