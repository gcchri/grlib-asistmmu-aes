`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FkFZi5h2UGi0ksdsrU1/PGdWX+6reYEAob0YRAGczPsywIMfcl1SrYTt78MoEeRN
HHfRA6N6DGCm6P9U8ceIMjxBNzNpzwwt6+LRgDi5mSC4VSSp4vOqE/kFgXFn1ijC
8g/Q/x96Z3Aj8tK8t0gvW7XrRxeThqcK/Jr0C7hUvYuulDGB9Yx9OxXuG3ykcXOh
DB1w3tYlU8oc6DKWSDSekxZBe+Fniq7l0buxkRqLgCS+r9RAaHHS0FMVrs8rO5KW
b9ZI9HRxfA3qv4rCtfZ7DKYr7kfsAy/p9Z6xKwy3AZdn+kYnllct4eL8x5ZaMaGq
gqIvOn71Vab5PTOuMpzHdyuX6qNJLEwTh3pviI2dvFNdWFM3bz8VJzMilK1MUC7M
iddPfIJ7+rfDThUZ7vjRkSwMWp06pR3HmnEkZjHfnra9LvqJr6y9dIf5HFn0Ch3g
u0/pXSnVf5Dp+bSs569sKejOgZX+hFVYdlPYqFTGM5+9PDvBWypiaFl41RQxsgz/
`protect END_PROTECTED
