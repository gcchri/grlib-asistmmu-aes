`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aNljnLzfoYo76DCCD0JEV8AWlMaVVMwq+yNMPsDP7gP495EXUpFewUgSnKgMzFQn
TzSTnO0Q5AjhGhDWsMr2plNq7keU/5O9TZTD9NozBmrrDDXnlK6Z5edyMfD3w6Y8
Cy10NNJ6KMA4bc9X8Ks3BJfOBGFO9bRqHMWiVTEiul/pDP/0LlYv/eVeqWX4HJB2
0QiG0/mmoThTo9mgTdyxQ6t6jOyBCBEToXXh4y+oxE7AweXMYQyd3De5XSH4A8Ul
/AUrXCusqp1c82gY0uZVcDSvDAOiTpFHPQ9cPOenM8IR8tEPArOceGLOIdw4mBsG
fyC/AftVD/++Sxc6sxTZx3C1mObHB17tpwcTTMq0ZZFtwcnZDbvfB8rixHbOnpgq
GmfPt0qzni0UQjigP+DEhri6TehH4iXKTEFLclEB4Ye8vFqsuEYgCGS5gYl65xNO
RkiafDU/9npi3KvK1wzgjZW7OiNg00eqYOq17xmqrVt1yWxEjDsAJzYjNRj15/ae
pWLHOIgXv23m+kO42tPlRCT+pi+QuEvBV99lRovd4/Fojizvybb1WXiXVJz6L3JH
121VdyYyMS3rZabvCQCMVA==
`protect END_PROTECTED
