`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Drby4BUO25GFr7+jo9NbQn/BW0ZAImFnlHesiTJBjB14JMLkegEGcdIZWnBQ+YFk
FV0rji9HTf+bI8R8X0xJEJ7G9v1z4gDpc3RhAQxLbcKpBhBJmUQYgbcMpTpuRF6y
M443uhg/PsoqmUe61CPOXk+eZSRxad2PjRvESZF/yJK0FJcTfMeWucBaRjOi0t1H
dVrqpNtXWtv6FjKeNn2WUGkDvTYhPG/V9cw6838/eC7myt0ZgSPlTHVqD7U1o1r8
aMTFSAtFuPh4Jz59HiPvprFTs5rgCbKHzfm1vJdcJmAto3jDKlxExloA+b6aLU34
QihdBryeAX5rKoDTd9nNsAP9TsmehgP+dquvCiMxSBbzG3+EKXz629J71bqssp9G
TJHUshoEmgUpan6xwaTVr0qHceSxJXCmVGp4tbBx7Sro01r5XCYbHDnUdTTe5MW7
vm0TSxHSaypIp0NrCkpJ3Xx2vK19pxtE5+ShLmQAVfrUb3ZRMrTa9G/noEVRCnjy
cEfkapPEV8uXmpxVuReDeyEkxdyJRPx2MK/dVVJjuYOefOc8ziycHlIh345LMJ3/
tNRWlVjbs1pM01OABKzkSKLvCTjadpMe7ZGmaBa5ATs0cjFikyOHouKAQrbrRGuD
igHxbX9Yvzjv7I4WdWK/iBz9go1nm3s51QW3ZN6+A+UJWJfnECEiWXFQOX6781wF
M/AP3amhi5FW0/+lt5g0ANh45jCJ2Qm29uPgPpJY6CT6idEszNh3ATAm8kXh4pIp
tHUGLLXaSj393LjykUvwTC3XShmM+7nuvBnIVNKtp8h1TNpwddmK9A8252UsZFtM
3p+AS0qMDUd/f6WYoB8ZlpGZjowJIIVsfZJLrRX2RBOw/W+SgGsQHYBolWlosayV
6JYtk+TRVdg7KkDaQpareDKnwGfO+PDHp/X/HvZocR4VITPjDne03sXiJF43hP5+
HjUw6pen+Uvhk7CbLB/binfxIqIzpt0mnc9eZIcWlPdSVyVbLQ1IOyI3fLxwXvkf
8hwhzc6KJDcJDKJBrhy5H/QB0K0vCIAmqRx92Wspm1e0T0WVKixrmBjRat0yMYJM
YlQXmtkW0YHCdZNBEYC1gXBzPMX1iugA5bZQnfCnUL5K2+NVg83PmAHKpBgaGI/+
`protect END_PROTECTED
