`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3jDcmMEqmow11vK2yYJeACJHGGtdudjiabTlAip6IMlb28Xm78rX4P8gJAnFuMV
LcngvrznQ69/AeE7mX8ZlwEmHWNyh66OquXY1A6EZkG90TYtIDtf7w+RgLeY4F2Y
1ssqM/1u3jqM9JBvtvoov2qQbjeVv+5j4dJgAq+HtcR/Awew8v8wr4h73GgkvqtF
Ru8rKmHoT6RExyh6qLNVDEjvRopPzxlsroZBwhRCNJbX5gqlLOh7uokYLIv2pega
7HNpRf0YEzfBIwEIHC58gqQ9JRLBAsB3hie8I/nohDVrxJTwRBqiTRAPStiWhN80
LFIxWeWFYgcld39yyOB0eHKZGb4wZXMz1qOektdddqVjVKj+wpMGBccRsAdTGE/0
FxqCYit/Elkb0ob+DK1XNQ==
`protect END_PROTECTED
