`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sQSXcq+t7FjratI7V1KOx7OHrsiNNiF7vxzWWx3eaBTQmn2nfGb/r3GsJeORZr8T
N+hKp5JlWqN4eY5guFYxB5aP6w1JO5PMm51j02gmk8A9q0tEVxSPaJVtrscg0x3b
a6alMa9D+3SDUWF/t1dNWmoerwGlZ9qIa8KTpBSSLl5HDxxl2CibPZ5XuJHgiiby
jie7PFRmJ5vdAbYQtwfEZmjhqDSYc9T3udIaWp89050l0tqgbPtrbiAJ6QKBn7Uy
EDSpd+q7+Ekc62MXSW0n8c7NwNT0WTnIT6sUfruvfPa2x8VWT3j68s3pRtreGYLy
8EWd9DORvP0T3Nm46plvo3QJ3aSX8RTEGWkmqlqDAVlVBJKMKWa9TwmFEnwdULbK
K/ssI71YmLhFut00C/e4m5YDrCpOu5IVbNqfb303MxsOvHu3+tFluCmBuK6y9gSo
OuKkrknBmXWPSK7XbMt/V1u+brxH7v2DIAol9Ah/DTwxW8hk8GNeKwcq3ZVFdctp
+nPdNwPibxhPl54sWJutcX8LrOaAm3bTaIVd1yFHZ0/gLvmP+Yvuj5HcC0/ITluq
RQ+sDDhl1bo6uBA7Bh9ZkZkTY8Sy/LTBSNhrWNA6eTeoJkIs1ZJKadWA9l3760mu
QU9RdUnFfiZBA/tS4K0FZLE1w1VTzfPk2/zmwEK/60P9l3dl8UWTeMAlLCM4M7uE
deWbB1YoUdsQeYdYl26nK/Btft3tQmHXOOz2Ux7K7Letcsut/nxRSIT6wQq5Cb0e
NUx60KshA3LTYDcq9gpQu5dwrhN4Ui9X0lkH1xDq/jbjk+IAxmUeqcDGfh2OKLWg
wiIiBjciibtbxuw3+8beHiuIJwubC3g5NL64J3nJCyNZyhtHXuQmDDFGwAtugOpx
jWwUgGVOHizLgTYaHQhHIT8fkK5a0vf++6LldmQtGABHg7wMqdChekVADfNT6DUm
96Y4z1zr+E6ozU3eeGaZhOCGGpOPPWps9VjpwZxXeQwd72tX0kWVYXrHo1QvRx7z
shefeCtD51SbdpEo/ztyCoZDBXcZJdXaMKdEjbVFZP48qNzb4x1gFTOw5yuBv3F3
927xCzqo973v7VCUZXaTIRBTUD4TU77B4F0//Gjk4FS2k0XPb93b68oJwJAA3OAB
qRB/h+KjvvJYyV7NLQiMPWONpJXYUh3/YifMSCVOiGxPWK4PMQN/V23mJlR9HwG7
GTAJ1aJv+AuHhWp4Eqxk1ux8M5OJNnVsBRy4sZ32I8WxdnUiCzU7+ugpyRvcZjDu
cg/kEA1kwYfeWzaHFTp2vFaiQZ+pjsSD60RR9zIq67gIN6OUhjJknolcb2uLnMi3
1LejRXJBeXbVVhvAN7UYr0RLBlmiPuDxNdlaECHKD20C1zB8gBRlD7//sfelgfmN
06ojcinwGE9tHJXO/mMWE1Tyxchn9lBHAr0Wtvcc0ww12sXxiFgxVEBKLFMrui4G
/Mo73Vs1FM76v/cLyWGRtkEPoWwg+tzLU2Eu9g+Tl6zV1lTQZaaZr/lRRrfRS51V
aiJnPvDTBvN6f8TCMx7gIaJSoy5svrvkexvtghnd+kvg1oeeaGEZibA4a3D1rRee
05foIuD4XwU/incjsLP23tVVsNcqIXcXV6eQC7v218c23ph4LakwZ4no+0vYwzYT
3qihXwsQDBYVcSd2YTK1EuLt9MMuwKp96kG7LlE2cffWNe91Hv4VoYsg3flsZ1jN
1doAlQarIPvK+/G0lSgImphhC0WIIqSaBbbTD7y1PvS16k2DK/SaYCVGfFyXQawc
Yavo/UWhlxXqwOo4Xj5WGnTDhcw9yYO5p7FLzoGtNmc3LeIj4FCZWCjJqEvNPIlY
aA7zkJ6P2KVXQ72QsgdxL/AU7KST/hOsgiw/Gr0+q/r59tQfwtOcSq1gTFe+yALw
3rr7XYLz/4IEVIjLuz+jjRE6Xhrb6cWndql/gYwsjWFVewVkM5G9m5VBnY4M8hed
NZ2HbZP5cJ7a9PyifCW2ba8bvEMihAU9Imkfy0iGonTY8e1P6mjYTWySK+GXL1Oj
FYLJLQTMioChE0mLQfD6oPThUUi8rahHzSHHONZKGxUsgjQtCXptKsmzNSbCi2vn
fbg2JzCJBoW8+gMip6nRoQeGcpp8LuGGdPUvdAD8qAufKhOOED4RL/7EPv9He8Dc
XHIzTfZNrV7eOGlT7VQrGZFrIQNB/MvN+ylzXoJe2f2WcW04YzPFtWs/Mmmass2M
OaadEO0B0pi+Z63fyeRlFeto5XLEjMx6sBhFwgTNkSYivJNyRqpqtVpGGNQEnGr3
k5hhBYsN7yFRGEhuCRmtKv4Vv6Hbf3RXtjhv6MdjssG4Ai0MlwzbcJ8bPR2+L+gm
0knhLcT+Mc2V+EzckqKOnwRB3TG4+Tbvl0+IxZnoLadQiFe+hSXek1oBj1u3F2M0
hCFnU2IvU10MqrU1qrvhubgxE3R07laDyNO7SDoSYBcUyJX2c2xi/wItNjTVqb5y
yqvQmYFJIiWh+bmHZPOlj9bDInEMUrI1wfefPk1mNxvsaP+XAjOhDfpvHJvXc8M6
Boqix3yLJQK9By/q2dvhdEcQTe2+IuuxHVwiNMsSmr+b6GnEN/5HHIzNlY22PPmD
Nm4fH9ZEc/oHxisj23yaNyMZg0Db/JWbS+qgzd+OyRnwsJve6yo3Pd8m5r/lQIWY
c2tEzM6wkJVrqBCJRwuIpYUo2pd5iMFd366KnRnJ7GFryIcd/XhG7wT7UUCEI2aD
F/BQifsgHM/C1e/RxXs8C9qsdrBb7zg2XrFMrAJvIwHt9vElg6yuwnB1D7k+S7f3
jWQRC6guJrBiRzpKtMTZ367Uahs0mdfiyiX1nnqb+3R5i9UT/XUoDEV8Vr4O7TRU
KRnn9zEIsxFeeWbySLK/P4ecVTzlhJl0gZ2rorkFmtAlQ7clvIgQ2BJnxntlAtNv
hnxU8cb25N2tLkG06DJQtJ34elmRf9OB4SMhbo5zaMrmLq3RH41s5bbE1h3gjEAb
Jz4LKfG0g6etCQbN8lH8E+x61UQjHcDYNYeTyi+HV/O+O/onMz6MUXgh5BE8Mt1T
2e+GolGWO5Edn5JZ1SPIeNfZTeJ4HKgtVKxvOVXBzxykXYzoGOsxRBi6aMOkyV6D
42T/mJDC5lWhm4jl7ljhobcKp4Hm/XmsXUq32Rr8P+sNBzRWoF43lJaceOIxBO+g
9VjZR6ZoEsZrA+WkiAZ4Yq8WOp6pEW8fsS1shcPKyAB4VNQPcUzhTL26C54QZ4y3
vzPF+7vNMHsL5SRrR96PR+EXXAuC4sIQ2xT6Gdwsk66l3bcD/PdQlPzjYPSzSIJB
PVr2IFYx/UOBR+wXBpkgBjUIjHMxjgCTH+Yvdcf8TOMDtzzTXlUSgUR6oiEAkCsd
MtOXRt80xXKnIxvI6bcey0d/kq1TxamcZHoUsMrPRs4fFtAEIKnNmhzs+IbB3XLo
jb3LUw8T6RC4PzqGTdaTSu+Rqc7T+SsQzCZm6gQPMGE9oFMOBGzCQMkBOBdjS2ES
TQWq0hUjWB2TOcbzqcKhcSPl2c/l6xrTP/4drmKDgLTAVLz0+/6imkpwYL4+rQtB
tUe2dsQhzDs4NKE5XruDyxoi+Ca5+WI9SD+I679lpzrQ1TawlJTxySh5SExWF37G
+rYzt1v0cDYWyUcNkUY82txE+JQaOa8gCNXMhvNxdJo4Ox5XDnz8/fy3FzIDiVVO
HqheZ4hhiyzSsEC2IB036iHAeTjOWc286O5REz5VueyMHPox6PplHp1KCu/fw+tK
Cbgc46DzSAMGohkcfoFUpbQz9Z6xYU9XbQ4XKF2WfhA2CaOKgDLEyw3xS/isfqF8
qHWwQJ3AOpXuyWkLyky4JKNFgkTrZPbsj54fy9DbVHIcdFjkyTXa7u+5cklTtCr7
Rwt2885vQ/NMjJU/dZYNxtvoZOFnTSlu7xFzWBsW2SftzZVpsIZ6pMmfm5prdq9B
5yudiCrGkFqYoD2/Om/C/ZeCnegWiQZCchJG2BFJKcjsK8e4s0BKp6EPOdNYdvT2
kNpIHY+mr5klGicsKfY8SW41Swe3/4CSM1DR8XEA9XuwI2e4bMcyrgyFXVP/ezh7
kES57n4sLKQ7plr8IiPZfpXD2t3xS5tH06jNnXM4Rk0TYr/hpwip+nxWFZPjV5Lx
dBgkfUa2tDr/byoMrI9K9UUonl3I+R47ItleR9PPi5l9noDeZj5uPnreNHAL4ekH
O51HIxWCheM70+2u5kRfAd4zddnRn/D58k7aQhBNh/rqqCled0CpmquJsAgiJXZN
vXOddMD6LUBECclC2rs/THn8Hywzbyxry0MkhKjplYrWa27aY6XaJwpNwLIqsQcN
/F0wbgRwiiTlcW/LHKy4NEsYsbHG9rkrpwn5p5/iw8bBKiz56Rn3W2GWGA73hbvq
ug/Ef5IM4bdhgMQP6LqioFIQsMdcvwqMHjjkeWXJSLRZAqZ6LP4DgayDHoeuUdrp
sWLcvgOcpcrZUqDF1M9gc7dLfzmOi8Be6kxMC3DEYTTf/MZoqP1h7KbzVl3rrLOQ
1khnGyCzsLYiejcwU6WLzFDviPoa/6KpRYM0CkFpoc1HiY5o1WJVTwh4Eu47CxXm
XmcoxNQcjyO9REmK0uPErPe7hMBWrcwWi8y0+7NY6gQ9pnVnBb7xwOvbDT6b6t5V
SDjZr2+GsLYJo02hBeJHoqRTinR68VJIpknVATlNQU4hcEwsVB7oWVmwjLYJnBih
XFb1pSHjZSC33g/ugPYB2NXUmie2Uk5EK0LS59mQY9J0zbByqFbn6PueFZ5lX+D8
iiKe6HnwsGZF1vXREwJ5tAlw1Bb6ONTLGtMvrltm/42bP7Zh6QPSqxVx8qPVwW2H
9gBcpt8gBAac8VViPMqCmo2/QSHjgvNdQyHAI8rAuDoWmVkZnnie/yvfzirEHaOu
kb3EciQqNC2gKcbuH57Bva9j12qX1ZrKFW4iAAGiCHXIoBzibXuae9a5aEXozbW3
utd5Wgr2J3gqdE2kDjFemRlFNv3gvWItCOGspxs8ieG1vcOzrD1e2FCHd0AKlY+o
n3OUcsuojK59yFmJg5yowK3zrF1uOoXAkSx3igO8gkdODoh2xHHItcudky/f7lbf
b8GrOjkSMvXAfbbrKRzoR98dfBk3zuPT396UOtj33AXNfJqFxfYtOHV8uj7TtY+g
yGkYbzUAyYslhkclaVv7pZzHJZdoeiRCxylG5NB4ZEw5XRHBqTq/R6gzbyWmMJEp
z1wTdj8TBG3ZeK99Oi0reemm9SgH2qrcRrEzF53t8Wjeof2jgs2+j3/1J4jdrH1I
CRuX+88dhoyr6aOGGjI5coZGA4NZGv2ddGH2EKfylFZ72TheIA6ocKMrBMb5RPTQ
2rc1A3fcvzpRBHEBNBLUn99hpWQ9E4U7m/glvwFH1jUmy7UhOkQU/oqeWQclaaLK
Hri/QSqKXZJRg0tp8dTlHakTYi1lgMxXql6dwVVlyzmxE8nlqQ2Fs3uWk97xuuXz
Qm4ikDEoTkBJ+HsinuqK1fK+qvXnIZEyzepyIIkNbEX0Gn3jwzHlSdHuZXWX8IMg
HNYV0JyANiwfz32ecVlkVG+8HKomnOQ4EkBQXQmWSoR4WD0JaoALlnn0cB1tKYia
gzYFbuW1HHTQKbdUaWNJ7jbuucpfV/zJ9KZ0H5DRuOSevSzFKhQdc8o0rgB8Db92
8LwKygTakEdwAVDYhU7AeFuzCaM+hg8hovZk4QT39FnBPCsv/N0r0yMHOinHfsni
0EgS9KEQMGg5Sfe7OdmKWGRA/Vutdsawa6azc4P50nGRSnmtKQBLZA5jPQr6MM5n
itjeiCUx87RwzDnWVSwOKoyK4a2eWLiAlmHPVX7SJruskMpk7uqocgWBNzryREvC
1ycv3AJ52e395rTGAnPu8PaDAstWTE6PX6PGO6igRPvCOtyLCiMw4Kseh5X7medt
1ZNHSlxozEOrit3sWr7u0uJA4GwHP9w/FRo7Df53FyC/Jl1DsUotsqNu/sBTEo/5
xRfixzixuVwyOltu8kxisvM4Ui3IN5n/B3HRFzioR9NKeXFG4rfNnoGATgsCAxVJ
JlYRkvAHeIEmQvTs7a3J23EArKmohpTie/l60X5+3ECK/8FqdK5b71XVPzWBY+9L
pLK1Xd0u+xV2+qZC6XFlXRdMBnTPbCl+6o2vGLNF/7fXTeY5SiihB8QKSVgHld9x
jQiyy+y816KfQxqn6njwhs7eg0fWNRs6OgAxa78xF/TzgwM0VXJ54/PytZF0zhdq
8OXN3gT1qyu6Qif++XJIvMpYnMnblT5pHBN0utrg5CKVvKw21Tv7zgZvle5IPafH
nWNr4W37FzIEvaGKoin/cXPOG4W+MqueKEkEm3JBDueayyM5TA6bvsQGTKBnBodg
iS3UwOEC7Kv7xNOSPrVWLiFPIlfkgUAPAejcsr7QJ+6kTskynjj92ZguhDp2y1/V
GB8ySUoHs6GDV0df0XdA1T7gy/Ue2lpXOAxTEdbA10Q8GMFr+lW6+rURkwjAJFAZ
EHB++7XurXoYf/fOZLIgv3jV1Kqm1F8DhMol+34u+apO1GbgH1DlYIZ5/RXJXFH/
pMMn8VM7p8am/B3+4rw0mTjSvFfYdyzGsaEqDgBFyP3HxjTrqbwGVPpx9KtaGeaK
BRG7RyJEDFlCooP92QtShqoCJwXobCkZyV7l8oiDuKD8yYYGNGHeQz/0WASXO0qp
O6gSU7FL5FO8rOhRND8qH+F8A2lTZjZsLcWyx4uvDLBWWD+hQWUNaji5FMhluZB1
XvYexIdmzFzY/bR7cYqGauKsu1eZteSo0zuLZ9+R9hqXX/TOy8kiiMcJ1fcJAVSw
GSx6mnqqiIhbnLfvQsqgbOpTZMIrEB/sD38yuzfO6zsrVfC/arMsivzJFhnke4jE
fjV2mHHOtpNf3gu1QK4pwzqrEkjbt7sh7exrvp1mMA2VBw3LdwCy6uvsENYLir9u
ruZcn8MtekVQGpQO+ebaZyO9+FSf73PKnPrG1cBNPxWC/BqoPhllpLWcrfXyTz+q
M7CVLxWGZq2nmz1xsbSyVcGtjN0y3Jkv0pIqY8Ubq/AK8r6JaZhcQao7m9H8MMYv
h8OmIXKO3E4eiDkB+6Q2hzsFY47JbJj7loOjG+5TNTzuC4ouSPE6jaE4Gz1TCsBg
6gn5/LZ7tXkg4egvy1YvZh61axhKOgRcXmC9ZUdmjFHUDs46GPi5fEponAi0l3tZ
n20U1YXcH33lXgPHTXNE+iQoC4a1ZKKKYO+xl3IzPwWzSmSDtQdvNtJZKPqrIVvl
hk25jRP9YNdG34pD1TA47h01P71vnelEU9A0p3vWooQox7/W3yPzoSEDC06Leo9z
UOpur+92+WRVmHfQUrCrP+e9dc/+o67qRlvYDzWLAz7s8NVrinS9ZKhmEAXHPLxL
OX+jZYJTUIj5GKqJxibQd4PfxEt1CjMXCRwbttnih3r/DcRtees/qZQ/Ng+s2Sbw
N/T1nLzQCHFo1CTzreK4/Yi42FfAe7fVbKna+/+AL0+m9EmB6rl9KcRcd8Dlv82q
XW7/CTXulzIT6Pm+TGcQkcaezoVaaD7AecZI7Bhwn6xWEHnCxIeUgCVeEbzQ0l4b
VE3BjH8dXxqJ9d+d2tBCrqhLpqXhdrCutMMpOTwZnbipRaZ0oMbou2k9BIzm+Li2
2ghp9SjD+o/kRzQ8ErcYGMtZLhoxKTFbskOOt04q3SoeZ09rUu00i/hjYCpwfxG5
vSrxqy2KktLJw7CgANrAlEkRg0WCh91uMSYUc3/zy37EZxh6NsVJwUxrXAHj++3p
iSY/jB+/hs0CFhDn2snHZDIaFfnhx3N5tVxN47/ZZ7XWq8nhT1zgcg4s05p9xw8B
GUk7Y/+37z4N9CEPUuPGt7k6N+K7e766pijdE/vKGffjynWd7YlLWywILhiR5d0p
bl0iQjQODT6vbv0MoLLgmWT6nQmfGs64fbPP/6NBf8ezynKNS+UfnjmTA7hkVBhT
yG5t8cqGM5dvmyBAr3kxjyYT9XpIuA96jP862TZKN2kht5alE1AjQ7SSZ+L138wg
No5qKp5t/UQkUGjR7ql4+3x3XhiAiF1LH6eX1UgbBCghasmueAaPya2yErgc5gj5
xvN0itXzgTjqa4XMJiRNKnPW1I7+ajdFTOsD5frV+wUNALJ0upKUBYr8VDMRgRj0
By4FHd6o3EVCMVBeTZaHFqgxv1UNjG09zRlL9ngaZBZMVu+qxNhanKzsEcJOIlPe
yoknXJkZGwJPBYmHuov2nzsukNfBbw+HdZaQ7TH6z2+YhYNGWadruD/I1pgqN4k9
vRJ+CInhAIPwioVkbzgkEFsxD/MiWyPIk53UhDVVdpi/659JbIS7t8CwUEikQSGO
9vcQAiyh64HmuP7LTofUoL8lwPS1NNSJULO98IZg8oTmND3JYluXDteN/6yIz9Zp
uGGQ/n8ABnVRUVVRDIejcg5rr+bmxHDBgYkQfhGE24AMfh1A3JxLkioEVs/FaPzw
zweLyYAy2blcinQkC9SkGRp3zGe/LaF9NcYIL4F47XnJ5kGhUiq9YOToKYLeX4r/
ufwNJcnSkQH92h50W6KphE76Tffcf3I3oh2tIaAPmvh8ABF6b4f7DnWOgHaok2rY
lA5I7ccmyF2a6vSft45NuLo+1ec6dmrYTRsrTs5NnjXZhLl2XFkO37I8E8ZMZplg
QzbSw2F4IcHmY36FO7gLHHLyQ66neH5Ah+rcv39a433MVcm2fwbA398kx8ns/LhH
tC11ve0PbN1Y74/DhsXIOsJZRXMWQTmxo3Xpos7My0HWJrkn/4z7/+13amB/P3X/
WOKQmsjtZ8MYRxYTmm4JiUqda68m6e90fthNiPIMV7y03L7f6VBYMCIHQcAvw0jF
EHkf1sWPK5o+H4Hyn6johOOIUo1qFy2MGDpgtiYJb9YoZQJ+uFABjuqqkYLXR/se
pnQEjnMQsDsSHDKHRe4L8M3KDJz6Z9rIU7Q2fEzlnb0/bVQblk5az3VhI88SdLqn
+tq0sRZlXEwsxSGQF8QMwFHXDRur8oAKGEJnale2giroDSFyI7ZJrHWPo/IgRHjt
ZaHx7EmEWRP/gB14KCamYB4Zr1Oi+4qPPwUniSt97IMEeYiNPP8TayPD/9T2n27f
TEYSu3BHnsPBqxDUePEXTprLvwjl01UOG1xXyyVhaPVUk/Zrxo9+Ax4k8Xw190/2
j9PBBaaPNdR5fgGsen2xjd4wIszg5HfUfkp37CUJRzzKm8KABjpmHTzIkhVjht28
FlQOt1DyuQhm/6ijw/D7vOKg0fumfHa7oDgCmikrCAbY3uwXgEetTnKmGsHLpPft
uX3ItDz5qn+8I6PSuHnRoBBsr0MV3Fuagax6yVB93FlT6vhqFSx51O5B6DWnJmTN
B/EgmFIMGYH/srNXr7Ni/MCciWm9paPXtPfmTXOAf4j89LJ1cQK/h3ATz2ueH8rQ
2bpOymff2GwJox81YxfV8Zti827L8Fjv5qbbvhJmEfVlPZbslJTTvTf8g9mVfn+X
2RcIE3QAaDj7K/WZVdv7auKALV1Z/4GGCTjtCurS1gJuNNeXWe4yVBN0qAwxNny3
du/YVKPuPxvItR3q4W+RH8bmoPQyVYFeHIHRv7Yfz01Qi/1x8XHDg8fMikeni3GQ
5uc4ynYS15SNy0ukvJOJdpXiX4dNlsOUpQsfGpoSPNrK+Uxxz98Vqxwh4DYdydBV
iJZ65Lp/T/+Lg1B7+bJWnxkDYdceCMjFwA4e4g5qtkmZkKInysCCoqGwmdUYduWB
e6gU+arR07Zdp3SBpk06IK1xUtMk4YEcvS7I+whNGW9RRQyNvtpjanbHMriZX4Rz
JHhmsGAMrT9bWuDmmehFEnNQOd3BkYj0gRtCqmidOdPQlgSonMLuOjXh/5c5fiDI
5iHATX1KsB1ksD3kfHGZtyv3z0Pj5Qvn+lB9PW2WX67XebvQxr8xWrvOeTMtgaVO
cNC+/Hj/hayFEl4x3sKKpIAJEqvqEfelbgAoWW+3smOzaFDzuU7u0eio7CLWCbEj
ICMr6Zv6akIeiWXwGC/fDMwMt6EIAgKujO2NAn5BFebv1JG7YBNFlszV12TPgqgb
aj1rc3eLLGXcLSUdRgSRvoz7eROscsfq5q7wdHd/jJNkNLEQ2Sgt4w1hFSk/0XPT
0nFppIzJg5/ljLANk3Eklk4F3fkAvuUtO3gV/POcbM/Knk6Fb2GkArV07TL5EvwM
xSvp+9ZrGV1ljCDy9jO0okTxjUgP3Wj1RjTwdTfK/JLheAcF403WOSevkjBRrQfz
i5z6yDm1GDdpyU8E99lgaQyj4DBXX3rGeuPPkCLWtOAHd9y9Zvzn6gdEZqF6qspK
3detneKNA6xSwqVdT06ejdclHbG4KGkdIbCp6YKEc4xYaNFBarMINW+oI0kCWdsv
BqUXeCg40wxx4Fs5HalA8/Xz/yyYruOylQOloTFRm8P1V0FgEEc9XSjdsO2Mvrw/
pMY+Ud3oACV33RU8YkH4sPOot57ZJJq/e7HUyTCwjWbcjPcLCNRx3ArqbT1Uypck
qMHPdU2s/1AWyTsQdil2MzhbOC6ciHsFFRmvztd2xG3cbGY/YFTYn8jP4tsdjaS/
9UDnShfcxUN/hVhPU2VhqnHXV8L/EroeNawjYdcJYEnICjlijM9ClelhRN8yTg2M
3mgFp7wlWlcLBlJf2TpiksIFv5STHV85aOiAr5+jIJRS4J1TJEseWLrkiLtwPQWj
ypm8ZEILAPQIo69ltVo744wKuukaomWECBma2Q41RBiYoRiz2VFj6PI2EPOc6tWw
YEeJCWY+dWumsNObyWdthrK53l39Wy6wxrKu9TnexvSoH3VXuwZ8uNCUNnPM9YSd
tnKKAy5l5xH1WRTdPn4xKzpc9r1Lt9LWcz93x/N8Yi8DEKgWx1U1r33JtoYvBxLR
6y/J+pgBXwWK1k8bB+7TuCoxVLYRDuDej9waXkRRtSkA3tOSccmHdJe2atDQmLZM
1olauL8Gz5F61HrNLGMpgSSLvQUudbEmBbQRdqFhiHHbdpkhUODs8MSlTIS3PpWy
b10kZctYbY8y+tldT+x1eM+Drz3nTy1vaCcDKS4kgTJPYqLfIWs5C9trnc/96Gk6
It+bmbYOSCE/5h2+MZFXtqE4wm+xCwbpNJkJo7Ls32zIfEU5Zxbwlb35K+f2/o9u
WEGFJ4tcjeiNN5r5Ylj09+MSPkHtP/3zhq4VKs6b2VT5+BKIkSN6grJ497XqU/ti
GgJKyW6WkXbzA0CVpy0w9gTlGz+8bfCadlM54TQQdsG475lB+F94F0/PmeUxNqoY
uUmMmuQkvBWetb1LJ8KHmOvgNQrfMU5Y5EGQVO6Hg1cbNzGlNVtdpJzKhFX1JKZy
Z813nnrb51RfUa5Xnfo3r0QOLH59CcXsUCDY9fJTrON1CstxlGwnu1huHgdl7o0Y
AoQz4wXiXD9BLtTQ8msysqHpOTaBKs/gwirqIXcdXmlzxhBN3Ck9XYmYhemOl8H9
l5fqy/Swj8BF1BhZJLxCx6Ahs5sf+IXhLkThaYyQTIcUa06FYS8f7P7TAxyap6JD
2T+SaK7uLpFl0LeUmTwMyhGPdDxW3juVi0n0CKSebip+dX414ZhV0daSNDJa+hMp
cXlxaJZHo4VUHXkcpaQ0QLh2iQDck8JyzKC1qB3DLwlMOB0C3oy356P1rz2TBKBi
hf0f3nGaMW8XlfnZFJrX8Vt4NEiHkBWHL57SRjT2ZnWfKWJ5jHGajHbQ3qSmvUeb
me2JAdyqHaYwjXfpx4fHUfVJnhgyW2CZ1oXHmtufp5pAnYgvmTA+FZZeY8rF6wcQ
zTeAu/BX/tEj1kfcpLqHeQzDfDQwA7FRNjQyiqWQj4c12NScHp4zSJwW3rMPU9th
7eDPZspfq01bg0yB0sZHg95+MrymnzLHbVqOTiX4L4uPSYKrZyCcSFZJhL1wAuE7
AbwqjD32OLOR8FrVgGId9Z4qAATdP1aMPTbhiBnf9CX407tcOJB+m1gr0MM6vr2e
B9tbnfAPoxmNHT2FaDZOyfAa8XIAo0Tcxx8htda9n4nZ0VsartKDQAIPJGGsX8xc
hfCNN4LV5/3NQURJBqAy6dkjXAy+0qI42K+rYp+s3qfy1c2Rj8eG5KuOujM9/eNb
kr+kh3dgfJa88iQLGOTGy/jL//poTx/54WHlZNIz54gsklNXm0t3vc/p8TzCrTEz
txO6gD7qlnIIk+6Ryrzzjo0C8QHnHFRyVBrLiADRzaTESVM4ydIZYylR+1R41FQu
HX8k+IBTUcC+FxmhLOuuOrUOlmFdPlS8sW0O1sH3S5tm6UXfHuk4xOCd8s3f2GME
ompy2N8/+G2w1tjY58JqwEQE9+dcT19VrWNR1YLbvjeGubd9vIyp7dk+SojwqUY4
TJa97AXchQJt73ms9hPGoSrgkOCotprCG1x4Mw/YAmRihl0NRS/t/r3GUDNVU8R0
0v9uADvc76pwsqby0DoSewr5UB68O0KihnGwbaDcWYnETXxXB0WsJ2qAe11Rjq39
cnhDlvtB2Sn/eq17DXJrpTykvTUHCo+GBAeNY3L0HYlHnsg39gwJeoLkgolaKJa1
qBNZiprNJK93ZlEQoOzQCquOGmiDYY39J7+sMXWHIyjqVv2GzDzdoxlXYeFMAIhx
rB7IWM6RQSsY0f2leiQ1SE9IXrwZBdJjQEyDToUDbG0wJz9AOMumfIeW1tj6Z0F+
DMndF3CC/2yvrHcz8hlZXtKVBB2PLRuhj25c2nQwb4JlI3k92moXaDXaR6/UtvI1
w1TqU8WMbp/3AgfAciUPEdPGyzRv3EOqj5RIHgKRJkKH7bLPoITZY/OStOLw5Rjr
1QurWVJwZpmbBGeWQRcT26SFT/TzD+BhghYBk4LIjrsaGnVvrgzaN5oNqY3MbNVb
KtJAlK4b1XJe7I9seConr9Sm8FNWh+JwQOCEDiKDqPEnLUMqI9uGBhbGv2ZLn/7G
5Rv0m6H3qY1fAaejRJk/pLIDcut1WYDtWTbX/4bcI7rXctPJAmN7F5RbA/NN0/15
Tt7/8W6lxnNstYVErwWbH3jztQQ7n7xPKpqiomV7sircmDdiwj6F568niwG2qo9R
d3uXQfxJzLPPL6fT53zjxqnRfBF9125m5/pjBOOCCgtu8UxcWC7/aacDHDTS+MRw
/Q99BwdzCsRBZxh4LTXXbUZ4CbrLfJHhpgKSYSGtXYTH4W+ncQ0cPsNQ/ndpLwia
/r/FifTelfeBmY8VFKWmzpaIQqKFWIrYJcyVS7Hb9jYwNRmWQanujT22YrliAuYs
gQ+ogjcxdce0vvGCRSFhdXt3wywrPFRsTZs2gnyBkIqyXx2BOTS79HjiIzmvghj3
LLqNMtOPV8RDeYKhF3nBpGTl7oVeORaXVq71eGXy8qvSiAUN/auGzLUYhiGELqhF
Kx884kVkGxYlxa2TMg+h+y3Za4tQBbD3Yqm82wGzag14d/a8bYTinUlxJR9WYlCp
7TRmeFe564c86epFtS2LzZ58RVhonZ1PIf7NOrFLx6lIEDQNP4p6iqWUUO37pnBt
3cVcOndZ8w9d2c4UDIbAOaj8hbVaFonKToHDqZh/GFSKBRVo/m1ei+PhN24x1vvq
ntIjoucVnNlSwL5ib4md63bZmDSYhDl7iEf8Sn/+Iw3+RwXICxknnvmYXYHTw0BG
tuzMpLMVc11xbY083WBXer1MsJwghnUlojv+gaUDocnijtLWs+6/8su4XlkwI6RT
bpqzRrj4saYQ6iQlHkV1sytZG+r4wgGAeuP2nEcvkxZutXWyC2Y6iKYoBmTbkGxA
+q23dAW8tT+qc0BYkTWCbM1FZHzRCsAGXypr6TkbRu1rSABMNcHNYZiTJ8k+ngAm
yDrkI0DEN3KeEiGaHepWsmhoYtbDDd7aTNxXwFvubeMdFIt8BoAyIgkkJH4q1Y9t
h4TjkpKmzV/3sjZSHlNyX2Phy1HSdZCyfbHm9blxuXAdLk5OJwSC9ZMFocHFRqG7
fiXxqpmZrPELvfOQNIma9aFRWxc0K8dlV+ucDfKyvi5noa39Ln9gaIZpOB6jP4bF
ymm1YohZc6d4Y5MS90pbMJ9jKDOqPSnMNSudEuUh+uHfi/TAAtMY/vt6kd/e+Dko
vAWHIEeq0HquPP/a1ycUKyt8nb0QpE2awlEWYcULRrPWIDHbSCXkLs6puGqPRr+5
/95bivN7/BNGz+9YzqA3noX6H8H/MAyyoaPlSMvzeiU2HRSYwc6X1/mzG/WxfBXL
MnEtdhvSXHg8lglKQOdm+mLukG2XIUZW+INde/Whe0KuSOrn70a15tHj72AY4tt4
HHbOgJJcOFH+QgBUsztT2SF69kNE9DeBHXhiXoV+4Jw27eaYDJGqbsZ3kbMdJo/S
aQYxYh1t/OMhZSiCmfJu932tPHZvGOs6d6oqj/Rr2YjdOBv1ZT2U0xNYHIsPMW52
w4oH87KyI+nOnLrmgyX+iebnzg94/ZPuIgH0Gc6GLqYfqy8x5++ZcVIkjnobJo+F
mXorNn3nL5pgFGjKq5y/WGtCVLGkHtbrkBYm9h/13IVChuRUO8GM4CcF3DUGcW/m
OTiCJlg7eNW98Wai4/iVoU2mv7Kbu4QiGJVR2Fz8FYW88+sF1kYDYSrAJGHU/3bd
aLVz7SEqmMt1tPyTv8YcUh0VIOTFU2qGs2li/6P7rBcqGsTFuDF2SW/x5kINTyeN
F/EFk7RZut6Hl6RmHt6cI7R2YQXWHbluNJ3qugY88JRtboF6o+pg2+cSeDxtHlP8
MtcjHGKnIss9MdRSjivnfapGfD7kkmQ+/inbDbNnZ/JsswPVqHP2fIqkxvdkWve1
P7PCwtTPHEnBnw7Z2UIkdYvlXsvqSkNE5UNLJkjhzWlsc4BDlLaCwC8F2S5mDzL6
/RMTcjGVAb9l1is0wiN5bYM/q4EaCPSTF9AcHdr0LDHyw8imScXkytdSvqjtGPAb
NZhfoQNTUNmFYexJRaRZS/NcspAF6Yr1lN5hZXvKaTXvlEYrK5YPMbfgzNFt8zZz
O/L51XUip45cLIQbTnAh35QPCBHg7MchyAJOhP0wmOPGuAKa9ZVgkA2z90H3ck0Q
CQ+eRcoLCvOHv8T3FpWCFRRlZFZ51RAISM1i3ITFJda0e/xHuLMq8Cx1Jn3LhGRG
8AVODHsaibcSMwF+PEnC3g1qejG5bpCKyF/aqt2kO88mnVL4Bt9opNDLKUOs95P9
tvb70zO+Xdv54EHZQ1sfahFqvaIocu7CphEXrbIbXrWYqTqR/P47IH8WjyRSrXPD
QByB8IhwlSOXH+CL4tK5OaPOJ5L+k7sxIzckyesBJyhSQDNqFNW2mqDLhyo3deNU
7OVAQ3duPBlljeYIeSlBFuYaEhmrC+ZU2bmEU7jHOmsiP9jD7Sl86YASdPKNFyE0
QxGuoXowGenqppSe5l+h6+8z2GX2OLq3x+CY3hYO2MI12DVLWuUuN8J7G7Wr9rwY
Y76lkfskF/zbZriq/II77DyWYqyMQm+uDC+kFiUgUnj98fTFui2978l0SkzgrHyY
Q+3Ar5hsB6DXl+AmTdCOIJ5eQcLCyuy3Qo0IpIdMDqCMvfimLGSQJRxOFpNJ1mq4
/gFKVIGq7F4cytsfQjocgScKmJsyH54GoZ7hcw4zSmRNRXOwBQrv0vAUADUYknva
imsHPkRjJg6bpe0zHwqp4iM8EbdwnWZUEIRMYCxIjvkhHJOFQ5N1T/sCfoz6ESi1
ONEwHOuk/zKrrgS59FOgT/hBx/xblGzmigJ/r+pp3bYc5CAivkvboMWG1WQM0dUy
5VRychiH3dixoms6Qiv83JMabUorswlz+kXTq5ajRjIU9Cjl5vNgAJnuRKL80ap+
MOnfiTHk+TkJvODRhcCIi3Z5Dpy/I3xjdWieTrFmepHLAZtGPivRzNAHDpL2b1o+
SjjHAe3QrWe/MG2+05klXn2+ykw2/noy0hPkHUQUOgRYqEkivdaTQYFIyiaL6YGt
jxSKmYntG05ad79VfciOPFz8Iew3n64kBbYd6lDdoeD5sCNY3XuhKgHv9nWJnY2v
3+HGZAOwTB/sYwX1f1C+umTM0lMg9d7hFu7EnteK7VpBBx+ewSrRDfyXGuUfS5T3
1szhs02CRsp1Bfu9DoqzsY32decP7b3ohJG1Ul775L3poAv8UR5A+pggOeQUzR+E
xyu/whYtvgU8xlu/8KGCw9qcw76C62EM/EExrb8FA/SmqKDb1uOkqMMqVIxptYNS
o7Bc/WpEidwwWgyk2sbqfAw6lswzkfGD8HwstkPL0TgDLnQHEbuLGUtCCGAdDU9O
RpsBscCKaoZf3lcAMylRgFuJta9burPPV3nvvc2KKkSC64/RuULVHx75e4erCmjH
RyWFYB+LQ6Q+8vw5ufhddssetVn92xZV46J7GPsKhLj/mwGJyMMtGAh/3mZmGTRb
+hcawCMnI3+ivjUkrueaEkQ9sbUcGza8eXXXhwJ5FfgjYcYqb8Ip/I95Yu1mhHpv
RHzc9gP2wLfdrIomLq6+rnjjwomQCpLykB4KKbpJ6lDKGiBzpGt/KpNjQIcGwftN
ma5ShhNr79uBngHYSeOkxlC0HnzCF4gk28QazAiVg8lo7Vz0bSrfYukQLZ9zcp5e
UUJPD7g4FeQB1OeL9q9KHmqieWyYrojjVZjx60ssU1HAVTMZQ3V4agVjxgY91YvG
PG2OcuBVXiZs8nGDUU7THHJFsWMRHIGKYHPeSN+zDxgQawBF71jwxCLc2unLNKJE
n9uc1vOSYn08+mYrqpnhaeHr7RKX8x1gP8c9noOXAxgupEwPdgMdJJYLg2LY1OQ3
N03ck61dua0ok4vtnln/HnNZB7L8GuN71tMwN19Y9+2+h1zlYpYS6DnkWl44Q6+T
dOPirjR2hKhcD/tqMlLh1qGNqeqpFX6aGc3j7vvCuACC96trvANwtUPBrlYjnmxB
9zeNQIYdrDKm2U42ulJVFtigr8/bniyM/1MQ1PohvqqPTXeKOPUH29kIt9lOYSBj
Hx4eqGy0vap3Sjvm9OKOOK6bTT3e3AOGA6lipXEtuhdfM9Srd3SyP1hrdWBqLdyx
x4hwE/Turp3dj2i0J64nj2y5tWCwo7I9q81jkVUOWNMj4MQzfP/6c5Zg+VCChlQl
jXiqau7Qd/hr2iKwyvH6P6HVQOrifRnMcXYX2nZ3UokgWQa0a7cIsgweGZQPVKAk
EICnAc+UYs5Zieg5kh8lx8TSgI+JZ00lRYbf7Y8WDzAT4ZXFUm5DybF7jL5M+y5n
jnTckOmpanaaXH/j8sHrnz70LFPvAbE3xQQlo2T6P7i/fjz3nNxjZRyhLN1eevxD
rNCgpOBjXQNQgiJloN+yxORnjZlJ18RpmTdTT33ZGWyw2qrsCqr0jwypvK96BvyK
zhaMgh8qT6X6OEjgnAUk+TBNm6xi8ARapliuJb3lLS1heaePXeRnUqvGCQ7qvD3Y
QW2seMBhE12Vn/GuH1TRyiBgrlI49xHoNdC41YTMDScOrp1kjY7qezaoTg49NdFz
y7kS+yVwDiATqGhmoouINyU79asaW8pXul40KZW15BSQW1q+m7oE97b3DAWhNTpQ
ktI6lZWdSJbi78Xq7drLnAoxT02uLiobtRNiOk+/+EzVX4PLuUvrM0twncRaELli
zq0zMkwD9Yb4U8sQnImqVAEauCwe2LLRRnPzt5DcokON5xE+rW+Q+740b0DmHJTG
lKONlSInDZmsXB2e/QBwbR9hTd5fQSezUiSxhKPnC5MyF+5dIs4zJYOEMStmetl4
GcGbY2s0EXpVidmyibtl0dSKXDg0Zv6og6cLCJAZxY8xq9t8gY69JVIrD932S/Nc
OgW4vH/F1xi4iRivgfUO/nfjtiVg6/a3MY2/LlI1Y6x5Jntm/4y5WaHLw/U0EOZg
0Qkkj1xFrlSlrNtg2P+YzjWl39sd9lZmsmyd+lonDO3kFCx4TVvVmWMEBFOsYPtZ
pD6IVlsAiGnHmoKTWmdztg==
`protect END_PROTECTED
