`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1uO8SExjrIT6LZMEGKNT+xbgL4ZblvSIUr5hIU6eCMFpjny02ymMWbCjFqkDbqIZ
wbjNYDnHZXM2uB781VGmo6Fi4mj0vMOPnIEicvw8fW8mVnAyWhoBxZSWaIUb7E5r
D/DBAbu45mt+alM7Tj2ILqIq0I+Fms/NkYJHQJLrmYs3b2F0Gv4BqCBvJttdnTJV
RqHA8vdFRJFVzDTg83VkO9JE4uYdGTKtRToCb7nioDTCK//dIu3AoKOOeiKpYvCH
sFCrFR0em8UGb1D1FIfWcrSn7Bovo5JCt+GiatJa3ehLNY1dPNc/RJhg2GCY30ZR
4KIalZQzYAiJcbjwp4hgKrzV7XF9kTgDu/QBD55BfLSJiBBg5SPgHPPxW7YcSeU0
iKb0RL23p3TiYLiLrxyGzMCAQ3xyiI0ptNhYGyCy/MNpmX8ec22EcxDkdPmxqVCV
gxfM1i8RZqUK9QCaSSShA9LbAzOwWrZnjBWWTvWPW5ClaKOA/fXjZV82JtTBpsYl
k52KNlvrUOAOHgA+n3nCj7LSaWKbtoFwn6Pmf5fby0Squg2+U+ZWFtAvATmp+QnJ
gko4DN6x94o6VtSruZVPVNtdhljsuTZ0THhmMeex7QMltpe9s8Cg/PdtLYfMZYG3
T9qawq9u5+T981WxVBZ7GSoey0yUL5JnE4MNmXP1OdJxJrYhNuyg76whup1ik+B3
Zg5H2vouo/ILFWSKFE4iGS1YJsxsCylFp20qiO7Sr/CD7rwTZpNZo5kcjigXj53z
JTG0X6zGXTLHvk02etewhA==
`protect END_PROTECTED
