`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sxEz7/sSmrf0oUrKmb4714Jm04PBOW4UTk+68E4/fJGuoKjw3YKWHPmUc+mIkWGD
Lifkjkh8lp/hZjWoj4nuOZFhIIulqEPigybI/P3U7l/n0ikrbaDC0RWsZMbD2Jh6
xJgRar7FJ0rcJt87dRRBhsNyz4+zaFkkyF6K+QaTDQMPmEohrLyPl+vEn9FWV2AN
Ep+8WpbJhou71iudpfd2dA6QSd6KxxMkBeU6if2f9eME3RYcfpV5e5+g0otoKLK6
uBG2fQttqZ7TXafAe8vqLEhQrUB6UrzxV8/T69Grlja0pPfrhcsL9UMX+a6kQ1m0
8TGjdStefsjOSa0yLe0OfsdIFsBFPggiqUNv+D8km1UPIOugb14bJtIp5leg6taB
NheB5B/Ssaga3SB8PsNidVNCbkxTFffdclNduTgrFf05a288sg+jzqfJjBt7KO15
m0Ch09WGxKinnXBpdVE9bGKoo3gpdhcE6hQ9hXRuhc5aP29YY7iMmH8ydKq/j6MU
hvipUZpjJt8dpIYdL3oa5yf5bY422oE+lcoGpX76ACbMEAfpWtoGJDujQX9gJrIV
S0rQaZs8VsvDVl0YIQLc1/Fjiz97pD4TbIvkmqX6FRVYQDXphwoBlCzCpQQsm53T
zt9BQdOGhWG0qjXwhhCsEQ==
`protect END_PROTECTED
