`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lhs0ZrfAZlDI8tgVl3c0YL198REzo2Z6SADbxvZR9MOXJGKSed/BBXA+7LvHVGJh
fCdPCgtdy41fgEstiG8Z+eUVX/g49Rlx1jPcKBd62V9xEZ8DObmh88Vvcy51XAF1
XcrydfjNljPBYtaeDlitbj3lMoFQYFOL13rSoMsNZuKK+u0DDlNKq/kEeIGF0pnD
cF2PLxPYu6Qri2t8MFm1QIatBbX9u0Vp2KTvkBM5zag8avTvlSUyOcD+7/zo8K/w
yLvbGkGvkpN+Z+dkcB3gG49Ht4IyoEVkKZX9SHnJvlzSiFcj6tspW+Yfrl9lRPEQ
VyNCgBrm/AfSPU+ooSrvJ4ddSlE7z5LHTrdTzLvL0PFLrEbacViai1AqNwshja75
Q/0eRnmpANHrrgm4XWARdbV/1Lw5YLt3SZOOGK5m4VpCjU+gNDuUBfnoaICXYqDr
XzXRIr+t1jGxr8Z7Dfb0WxAwAssqoG2zrNv4NjZrT/CMbT7gCaG1xLndOHCz6lPJ
As8hS0P38W6uGixPmWxSLa+oxogqDy9cehJHoeJvfOgZIQZHe213W2DVhUsiIqTT
ZkuM5HoWxGW/VVzcgJgRjavrgHq/F+q4dYjEe3c7qpeLzpWF3pjf/T4LYcBEgHLL
nezdE3ikmU8tMGEOBHF5yWHmsR1edlciX/H3vlwACKyC30qE9jjRruwzti1YOixu
tg+xbOgD/0fLQy2u4yMPb+kDGMKqnxgEKfdxRSz0FS5ouM6NFuB5RMgMlJDs1ao+
zypv8UrE2hnZ+HrKh/6fX5WZ9XQBndSOxWdqXPoDidQoqKzfjuDSz1jXm22GcOvK
evI2k2dru20/qI8JnA+NNbP71ejFcLj2lxsmDac37GVAHP1+8aLv/7L2s/ROCcrn
VEkR6lzIqYUe2I1Wwt6mgHTqoM/5k944ZEe6rg35E5z/YuA0w0wtsOPZYowFJTd8
XHg3qAEvKm66jl6r2Dtig/WwTqZ9K3f+FOh/fnwvvttxPAatfdLgB6GnucWyrYvM
cE8l8xbW/UN4Nx5XgpGLU6+4cmYEEuxRM/JPQ3mc84tcovSK7ZY+YwHXX92ccwDC
t385LuKg/C0zk4DyxCVenivDb0j1/VuY2VHoOEWeU62MnNhgfdiYda5af1d6h1Z3
7DF7yjLAhCwmrFG5GRwLokGsKiEp0n0ULNI31WGbvo1Q5zT7hNxXeiuenaL11/6E
hSp3vF7xuHe4A5cF/j6FjP7E8SAwRNzh8V2AHdNTCO3IUrr1TJZkEB+bv8zQp1JD
Zl6g4jegCgMqF/MGNZIVQHzPDtITD/MySQQWafAeyYGA/lS6qwMbhIZsEnmqK12c
ECPIlWxygNsiMO5HQcGQXkJhRvVfxqNF+6R2BH29zeJM9rZ9o/AGog5FWVjBp+7/
7fxCkOuiNL1trlYJ9YLdFuJjiki0qo25sPocQaylS0xV9fh8EZQZ3FZJwlqlpmQH
TG4seSDcxzOPLYjL2u8LDOQRHBM4sZyAp0K8QLPS+iyZHRmpY4L/8Fr0XkHf4l4f
uBbXBUOa226Rd7XS6JPBp8GGCIE5shVElgVT+FPextxrwICUCd83luLMBkxNLBvy
bb9X9YKpS44vlOGOGE84tQCMmILLAR9pPVr91NSPxgJWs6iBIIdb9ovTwqB6b/6I
ucXvE7WNFUjUd/jmghN6Qg6jUzXTuvIQ9JKUL5aUTrB9zk7jj7i3q/BhM0WMs1AF
NXKAm16F26CgLwhi6zmbfs5u0QfsawRdnBnFOrMQ4J4EqJ/ppFM0NMmipFDXu36B
8hP7WuWj+/LlDBt8wSrZOtZuVfBt/xvBFWL7iG7AsJFsxAjBQuzv6lx3BfY/XIAn
TYDb9B44lx4YZytGFfTLX1oppL8ezlE7rWJ046Xz+rQZl2LR7PETSFTnl8IXxCYU
cKA3Bw+KOChJIK+ucP0+J6QbFUf2QrjDKjwuKzADa0fDyLaarx+ATdTUH5UF1IOH
njcx7FiSn63dE/BIWifNcu0If0kWQkia4V4enTlZkKdbbrp2iy5iZx6PZj/V3sNu
gr/MCIOwwlRPL3VDFf93w/BcHMJvhMGpbmomRSUSz2oj261XOIyHyc3Yn0ZxmmoQ
IeFSxX+ybxsekdjlWrpVpXYU7oDrly5HqEho94tgJP5WZTFMDE79LspCNNRSCZSM
2Itl/h/efXd6jBpmlqPdhudRMIE/SxxpCIvpnS/TuJzPONg+g9O0GsgfGX6meXFL
bKYXDkCvnuvCjUtsDm5jkbetKOEjX5VZC/KKxkL+/zM4bJlX/Z1UjfYnSNKEU089
/p5K86dAFdDT7VHSCBVooFsEVCFGv2LcN+YPAbFQr8/zVqe2VBEwFY1n5bQZMPH3
/8AV/qPM3cEWlh/ZvPh+FKxlfp+WAY4qJJbLj6PJeMUyohjJ7Hkx2VptvWyx7DfY
TxkBBF24bS0KXUgQpTLRveTsikoLNElWrNoGMvKT2pbmkFmzxgqP764zT3STPCIs
xMAhYzxtuh0m4drW4hXOYZKKO+1loxKCIFS8pha+AIZPqCbXQDzQuz40DsiSHN1i
oP0aQ4sx0Q1ZU+GJyYC4bvxP13bmkCeBN1omixCetwPGVdz1Uux5HnbFxkr1sLmy
ipC4v4ZUEq3tdkXZgA+DunU+DuKpQM1P4+KfihXag8rPE6bcXMueKbX3CORWlSl+
Q1Uu0zJSYpuq+hKKBLw+5lI4Q3lE2sk0Twkxhj9NMK8FIZo9kUb/kvlNZ180CsgJ
yVIXQJBq73/PoHk5upvpYAd5a1RVH9DnDcQSbVeu9nhgdI0Xse2+UVCDHm1qnGWR
77mw8WBBuK+dpENurKNzyWG8JXKr+rY14iFWoHJkkG064KAa6VXg5jyu0sMhUB6f
1LlhKgoDwGYLR2kKm0I/qo58wdXSZEuBockukCxmqqzx7u+VftzmeluUkOFIP7iB
oPpr5FK0p2LNFxVaib7yOTfZ+jv/kXX8ELmekXT3q8WXTfoJt94sKRUchano5cgN
AnLAz9XfSOKcKteX9KqlWa6GyN6lgyTap6rQW2v/oI38mB9ZUfzXJ/tagVAWZqf5
r13OuQfm/i5W74ZeNwRma4aliHxgoekfHbfL/dDTxdEAoAxTWJ1QXZ5vQBBhHKbS
DQArtmhfPOCLmo9PAuc7CpPlwgj3bu/angAaRiaD1CUpU6BE7H1znTook7D6ePYg
ThU/CzwDJG1GEz+mULsD60cX1cv7KlLBsyXDFqaaT6DgQaGdw0p740jzOZdPBaGf
ug9wJY16WD43jGkEVXchZyURxYFAo22uH6CCa/lvUcr8P2w8UKYtzelmgIDCrdnI
9UELH8u8W6szIsDx4PF6j0hAcV6Dg5wu1pHpDXr9IlQfIaB8/TFTRpBbGd9Rwc6D
8OR9co8Gyujjl0qa0IqmjCCe0aSF6p46qXGqSk1w8qeqeEwKZC10I4nEkLIQPfKQ
z37RMQ+13waZBw59qy1RpqxjZIKAntnBtySictHeg/R75xxtq5iJidHU29tayMXz
82E4zXaWzU26jXfGFfdcYa4j83zD8mFjtKwegpzvP0Gxov+48Dk1z+t0anlGKxFq
VkCQu0CMLdurhlDkx2dhMefCw9/oRC7bzDmeFpoYWS5wd5bKQKawoTuFeQUo7VNA
SztvoPTlo+8NhqOXi6TsDnESoN2OWQQ3t0uPeCSF/Ijmyui7RqMuyfyTwp7lDdlW
y9N2vbnyuR+hKopHDa1xVp1uvwj9symSeaU3q/9f1Tgk7cKtWmkRFkP01GNzfM3z
5cbfZ890ew85z8L+9Y5PVWRpdWPt74rMq6/DNBiFu4o9nfV1p4OmA4z1B5qnbTYk
gf5vBEOHpxVO1ZnD2Ykusic9M+e9dPkewhO0T+3VM24JEIraQ+8LCTZAnDchkTsG
NK9TWYJmUhktzufGzkfpFOA6V1kgC3x4SeRxvXeWVWeWGJVQwmrfcyTJSpYSmsgV
dlsVz+IlWhfqNTtEOiywZzyCVqr9aFb1X4CjqqcI+gFcY7lcJ+k8MDtlPl2uYGHJ
4zixVymy/ReTNXpOhTiD6LUHoJ99+ePNsM8iCeNaFZLxkzNSHMVsE0p6LBrmdV49
Mf9h0barOQtPRYXMnmz9VlpMa/08xxCKftxLKQXKaxlHqoiNQ3UR/DVPUzrqtkCj
xuuogqNr0CN4LuIYbTWsx9ASU0CPU9D+IYa1q8ILYCYJ91tiXs3jQNkficvIwSjw
Ex4XzbcMLLXBspDHGTqNV6k8JaPx8rbz+Gv2sHMD1wiCvg1ESirywSegOAC3Fa4p
0AQ08b2+w/ldk5kSxtp8bpb8K1CKRd+oOcWYRYzAq9BrC5gONBEzjnF0/E7CwJRI
5LSW77WRS3lZETvq5ZZHeXcY2g1NWhUAmp8O0tgalD2t/8RQ6jfoaMZrRSms4Hwh
8NnkWRGlNj/G1h3Ss8zJYx+QSpLZ0PLTcKoENtM/IKrqRO8zOdzs8iLFFhaeczDw
NmwxDcl1aDML+VgKUzBih4mv4nvmkuIbelG89BG9lrlfSyjdWgyJfkKxCX3+U/Kj
7vUvE28EGKExLWafCyUGxEjBFSoq7S1G4erPSWDmKBk0vO6qnFzqo9aZ45mvp0pv
EQeWT16hqXEcnohP7ZIyHm72zyyTpfrUtu5l6bGxyBZAJ50+Dld4Ro9mKXw3aRG0
Fjz2iGOQ4QFMC1S6mTWnIeeR4sGPJvY95DldG7o4lz61S/+8YMjr8oZVL3R6IYhS
5k//WHufGEd3P5XmWoeU0/GmfG6X8/vXUtR+d3hrsGNTpsG4Fm3Bh2BfEWNEH08w
QYW1XbNDUMmDnP41jK93dBC1u8L+ok8Jn3/qExkdxN9jj6fKZnrZfM2QI3ZYGr/r
F+hxCly4THrkeY84J+t6nhytMMtVe65BPy0UQ5K8VuPb5XmHIFVC3CQE8sJEuECT
2MdP6Upkg5603FKSbcjSs7P95snDmRUJXg1vFXJiq8G2j0wCKHJ37dH3RMqxx5+p
O9mRNZaq9NfYCNSyKCJ1NzVnLov7iizFPYPUxv8K8Kvr8zTMCaa6Pg5QTACYByr9
vU46EWRUk1L2C8XxkGwqHZ0fsobnyJsZFrB+s7K3lGVDFzTx/CoKXiCTTRMdI9E+
JxioOv8RrUHb5rWd7E6GP06vKjBigr3Vk4ZVP8IqiXpmb02KjDsE1tK1IlvdWP5E
/TWFydiJ2SPcsEUxVvslMN5E2MUTGL6wZI4hIk2RMr1wmurMAJuBbtD39b9/YpR/
Tv6SZe6zTvlt3oU9TY5ZqcKMMui5o5mcE+TlN8FDAjIdlUB7DOFUZNfdXJrRadmb
djFY+Ol+n58DVfoQRVr0luvHbnLAvL14uieT9MYnYuYv+qXKQTrPcZKzqNqxrpmu
e9IGKg9IuWqzV4l5be9i3iH5iST7KdJtow5EPgMoF2eXq0Yfs5s/5AqMW6Y+4iLK
G8Evz9x5l0oOt49DyUu0E1iDuW4twc6L6N+74GDtcvIZjI7m0p7Kv+RNKaEm8dIg
Xydi/filKpTvzmwReX0k6M8dCKq4yWGclrNdAVeMTn6Krsl9T9Kv27UbtkEeNUQ3
gBW329iSgw7cl/SHDIeeHAcuZtAAtVEHA3qrwfTgvqhynojuWvjxOkvibNE/hIdO
emQezyr3XdHuSSkJuUNIfsJ1SBN+J/ZjopPbQlmfmOqv8lx0Tn0m4UQ3hHWDKx4b
bzFZRSODHLPNed+yntMef4U/goAh9sLV67T/GvM3mEU78S0BDlOJBrYD+DDPj9nx
ezuiPOZtj8gK5/63I1bNInqF1sZdwGV2GuwuwTIxeT20tJ+EZ55uKdJYs2UOu7up
kLDEPZ4bLrbsGHVW5NsWrG0GzVH7AoWa70BQJzdAupabMDwgq/Htr+lzDz0wZ+nh
LFfiF3Ir7r3BTj/AwWdIIpZuj+cjmdS4jRrcSWc67aqmd5SS/E93l3/wT1RpDEB3
xCn/2j0mL1tSPwa23yClslSOB8z+wyLOURzVbXh7E9kbLbVvQhwNb4ACwVGCtC95
48fYLiyQ1sveUs/nNhqPuGG/5W4Kufc9esQxuZ4GgFPj/rjjgaK61EAGB6P5kIBL
PLLrkymq1WGwLuqG0Q2MSPPouHmNOVi38KEETV0TEUkX75GVHpqEVAZxpPivZbPx
tpm5QoFBV+HgSlwxnXcd5GcA7b/H5DaI8YZEzBYJ4FgGrbgd3MYkW0Na8Tad6X3E
6cjVmZCX9+YXP0hKblW5oE1Qhtzz1kHljCvLwHXZEjahRO2VxHNy3Y74i3ETlMGg
2wInu5LwxOKp6FG6bQnEtnEbLZdM0ySIuKCu1ArLjVfPJ/TO259sO604vUC+k7ol
fJb1yknShBX8aBoLYv1vY2u52ml4c7kit3NJx+W7jq34m7iaoEWChoRmrKnYcKkT
EX/yHOvMzd8sy+oESqWWjSHcQzxETqKVxRZYcVYsamFBTtOmNjIl6C1BSkYxV0vo
8AK/BIvWtalUSeM7vwkdXaIOInq6rNP5UI2ALadioMfFuVSxb5o2eT/HQ1UX/Voy
mEDmPGfFowOuIZCm9TGAHReKYMqalegrfCPf+7c4T3ujsap/YH/o7oiaBBlNAL44
l9yR2KxIPixyXJSbMJCx3ykoG0shrWhGVp6s571mtXQAsFXVg3gkaOQmW39Nm2he
AfmqjpTDtQOdwtKzcyOWZBdpGgvNRodGZWcy6yuM2OO2VfIrCWczjJjQGBDaH5Bu
hGjSYy4HXp8l3F4zawx6PBduql5BCJejEA4qt+MV+dUE5RyEYBkp4eFYDeEKAB6d
BXkCXmuWIR2sf//m/bLTtgiHKtd5dUh+Hh9aODE1R1J47c51aj/wi7GdffKkVNYV
9qDIfKi2KMxDj4MNdJFSrC+bdI3TRwdPVqtm0mtHg7RVUpuKN5gErlXqIpOUUKF5
HwHz1LS/OUxFXlMkT+RoG06qhhZtTs+Y4swc7crt0bnQX3/oBS33F1bIXWn3ZzIf
drAs2pJGIKb1G8p/8kYKz1CwCfEJXfgSnYK/iKhxSfsvuXu60EOCaD0/RV7rVWxy
FYkFATieTCYNfhVaGPGa6AHbOXCDB+qcgZMlEG2bS5z2MnNRS1PieowKEgQKgwO5
hOgsJz8cORuu6chryCAcF8oM/iMOBHa6Km/nijn22rQIv5R4X1Zok+T1g71dPx6D
pcTPyBbtGFkbkA3x8rCr5q/pHGy9FRMgHjKtNBShhUD+FC0l8HZhnGFQ/hMOLU2B
5UgIKurz1YHGgVtWArQnCRvzxHt9ntFtfaFRGnvaLxn7yqTSFUfctGsL4XJqaDcl
ngFz2NtKlv2Y+34UnGFWVers6GWeWK4U2rI5ZjxPUS9i6PwQlKDGoqk/8vXzXgyt
iC8270SpsaiCqveUaeBR+c9jsnDxpJjvvbRGB9ork1Kvowa8DkU8l2Q+fOLVVZtT
SNE42w11f4OgulV5gx48y35dV9E6HULQY+EPXUdZAvXVvSgnsoOTKk74WycNbMc4
0gg6iQriYMM9DeD7NTOL7WrVw8p25vTGmJc1WMcOT7U8E+nTCvO6UUTecv6rLCS8
hIijX0QgV5AIXeM7UVxwfQYfLbvll7iAynUflKFYV6am6ViVj+1cq9S1sxiYafJK
oPCn6nFxu5WOiyiKyLilQ2k3KVkN32CqRauq4XVcFa1rmVlhaHJQbWrirZwr9c1A
pAiRvyTHu7xLh8fmMwKss02nEu7IvgaOmm7SM7jzc5lfNM9rHgkz3MSik4GfsltQ
Vt21b3WrFo1Hry9V0ZSz6rrUjAqP1MxgdBq7znIMZ28QjjLgb9/ntZwFinFnn9QY
4kXBI5OdKDz2y1L1lzdgssrKpcZJIywORNBvieL1VMqvY7X6OD36EJsX5qzC9Xzu
ekvR6+Sxxom2IlLZkPmR+x3FrP/xtqe/5JgSsEE1OQRDPD03rJoHFwoDD7kJpExn
6N3ASYH+oI2dLySX7r6xurtaO3I0XtvVQm0DhAsATAQ2SwOsqAhtqOgOlGWGvbEA
mu2eIyMlyYpoLn2Foikscn/JJkls1yarJxR9ZkjvMA2NM9E+kXzmGeSWkG/UWrdi
bAPZeT5xlSzfdlNRA7aKKDdGW6+eTx44+ipXDUb4MIoQ+XzCle2IOYd8Q7cRkaBY
jltJ4L7OcXX94Cc+blVBj3BuzE5FlWRjeRPBtHHBeTlZ7yXNhTDkpXXODymdTge3
AxLh62z1X/ivTIrnShteY4GyGJ1BXCiUd6jv4l8n4lwpEPljdqIFImc4J1arB69c
vcMbnzoUCf8uZGTDoSsvK3mfmbJncjsTY7Cd/HySFguUClZaVcuZ8JSL4f+kurBA
9h6mBv7X2wOLMC2SVH7pEKj6L0e623ZpcSoZ2h0J+d6i7X8Pz+31M7tipoOqyHtH
NPLCkZFzkWUQ/JN9NPe9liYYwX2waf44S3m66yzrT8Ibu/mKHAa5UazFluAY4Fqd
7WD1OwhzqJWWq0PInA3Cph13upLYNFwv35PjcxMTRHzURJJCV2FShfQtF9AOl3AO
zOLrKbHurv6YwfRatipO/Um77n60xfc9YmilcV8rhsNkqVSsA7FsrH+HlplRtjwm
dty5DsklH3pz5eUC81iDIK5NgJyuz6Xe9fBqx+BpSgWxnIxNUoyNNlXW64JPBsiu
3K+WOeIEqD2FnNe66gEeHfOpe131ydLs/yqJ1R+k6Ukzp+cXEabQWzEkBGk6oMqL
e86SEyObzn2ulKkME+TyBD9a34Er2lmN4WlCLUHiOFBPhaIMdY9vNeO64qK5VADw
CVgL0U2iZX77/Xuz/KJoGjD9154vsLw1JXloyMo9kwpmHP36P4YVw8Gd15sW0KwC
PMvPB1BXRl7p5c2l5A3tZJAPc0a9HaMe05W61Fn2XxzJ+knp9Ycu5G6xlciRdok8
wDVATIhbV81QJq2CCAHX9Npo3l2tX6tr3p8qlcUOpbRQ76H7q/cv5uFuh8NnC3Zu
Fo4mGxP9oAtc9TNVApgiEtkBeC/lGuenGwNmytzlfmANym5PDopcdPFOGPLZyZO/
M6qibWgyp5BVs7FiC9cQJEY/h0QvgAncO4RZOeB9SyHD+t7DlGA/sW9RU91nJR5T
f0a7Fp5HzJlCJZzBAubzdT5meF4C5lHePv7gVM8vjiFy0AhiorklS40+D+SDVM5c
aYIlCngX+JVocxopBSNcCHwtlNBI6KjeiPAU95RMJWF+iwACkSQapJiRy2EefEYs
ek8ylLEdT07c5D3k+Jhlyj9Ej8A+Na7DC8XKa++VyVwfCrGC/xYbraWzNHJrDBn6
DSZqPGN8sWeVwG+AG+HZQN4+mneXoqPJ5YqoNDRK4oDFBU+J/EUpUV7W3yWuDplN
yg6aW7azb/THwtCGyYa13A9WH7/XDbkvEBHFL19fhxdrgBRNgRmmXxivDMU5PlSi
InKoAcvDe1DiXlio+w3BNF+2q18NNs0VAqOSJqKZAjXxvw7fe9Al29i2rybwVT+G
LV/Ai1ytAR+yDu5jzBZyN6E3tyd9Rd0IK17aHGAXLUkYTXpEv1Ird0XNtjk8fwO3
IiawOni1AsBmt6wBxG+A3rdT+f+akzmdevOZLPnRWMgjZUXLHvTPizTCxWAv01sg
Dgi3tJQ5nCyaf2DGJrszL7OicFED4F78++VYcljBCg4jVGKSDZEXguIi37/ijDUx
Gh2JzafRHZNKtpTRleJUKW5MB8ZW0IqFr0NryV7B97ZGrJmMFVtrlg/B3wToSlHc
BwwDx/RIEgA3yIffsRg6yerEBoepIVw8sqaDOrd50VqTT2hnIW1uZMvVUkdWTrd6
9+30jw/cYRQnWnh0+RWB3G9uM10v1ML61uO2BywhUvhm4i2ahegj5bDqct/O7bPd
iIS7beZ2yA5SDhEDhHMRjwZ+tBNmXWjnC28Cei8S5NlTS9YLVhEXb+qiJcj1meaQ
iUT9IeXdScEn3+XghCeVafIi8SNnoo3ychDFPc+GIrfnCDHj8zhA7IVU19YGAc3V
3cXU8GABhmKOdeeohBXHaupl1OoERve+5swBqMU9MDDf9YKADLSgMTobQoRQms8l
NcMgnjlbxZR+9OkqANTxOx81TWdpKOmahsgFCjBfUK2xU8+QLXufx9N0vLlqwCpH
mcIUzwO2G43rUxEuGphrMxWyIGm7GBW/NaTnCZWbzGiV3JVWNGwX8GO6XnMqH3i+
TgUq10Wq223f4SWGC7q3STH1Ye+dzb/X0NvYguO+hCmGrjqhDlxnQl1fuSiMSydf
1D5qB0kcLm27G9rv/IW6FBAMC7/2Vqtk5O7SPBqcLTP9kzRPTqacPtoyeXVDDDd8
lzoN/hFEhQRDQqHlwqoOglfYFaQZgkKhhNkpidbfBLT6Mi3vN9bO5MhnF/vqW3Pk
/9qL3sGWXi/h9HTxCtnJsjGUaxgPdnXHJRPSaJM8tCiZQqxywZ1n14QySR7MuAOx
HNSE/EBfcBpqSwBMn/drgsnLaVrIPUBDWdCN4Q4m/LOzWxODbVHT+IYaIS1vkvkc
/l4sHZa8QiU1K0WdPbF+1uvnNH0qrh5H0eWLq4AQNvrWKQPNxow+/zVe1syy/Ku9
/HyO2ICDS1KJl9p3t074gC8OqKz9Fe2uPtKINdgLrI3I3N69VDH6gd0SYv1dSTpn
hEt2VcCHcTrhrOw54Lc8N++h2hksK0ZYHB/cUzivb2m049E14otoR4kV+KEt9jFy
zerpXtspG3P2jmo/oS+XGwub84jLcGkz0S48s4EAJLdMXGjt/5MAAzNWyrMAcfBv
RiGoXH6hMKgSGakCl11o5gL9wblQta1JjZD9z/x5oOLsg0yoc60kb/Jh7BuXbFdG
+bpkmvGTmzpuBW+B2xK1ympOZROJAzYmaNDV9wCfUcRhCGV8pagmoHgmuXXKrsEL
Ku78CZpvs5c9l2g9yWrWmvUfUiLQdnIUAaQlccX4biOpFzLSNt/2vLZRWUFPwoK0
W3fPp4DxwOty+sBUQWll7lA4XSS0skGZ8BiPKHh4bByKgHanOvssE8QujpNWC47R
HjqxP6CwVhMoPJPyU22Kbnb3Z2Fb+9c801mCwLjEmotiFM3pACCHkQP9+h3MRA2J
O6GuEVZgfSICbydFo1XhOOAtbnCXxgmVS1Kd2m/7y2o1F5eCaEmltgxv1uLSFce6
eMFJFZxjVf4Ogt7SUlrxXlIPcvK47+m4Y0ao57WbNfj8396B4S8torYISCEb2WaU
2t+Hxmb3rENjGL7OQcj4itHY70+9tsAFxyByztp8DrHh1yLarXJ0ufirz/cKLF6W
tTD7jUUgvTHccD4RZne4IvXeNfg3taSdmnDtj5TYevFaOwPUuu+lPPqpM2SBHc81
MiqHFeZGqnU4jzXEoGDf92vNjMisNw7vAgv7Qv+A55UiLtjuMY2wr0Gdv3aj/Uev
Yqr9EZF7r55cZ7LsK20gtg8/ZzEXl144g+n1Ruortzju5nXDgYn3SXHe6TFWW3Xo
mEhPF3LGv+WieMPjL11afddyavugEQ+vT2kEdNL+MmKV0yrl9BrW8p2U5q346WzC
++pTMq3oPSyVhySCet9kCJ5grINqvm7UUXLvwx1z08n0Zpaz+WkcWKU295A+KHqO
Z7338XB3qpzCcXqtErQbNxe3FmNP+S4F+EQBWzr6/BRrAlaEnd5cGjgwIcHwOzxW
19zXHKwc34Iex1WlHBRSUvUZSof85bsbOu0vicIBk7OJV7z6SFoJlM2jhskNvqPk
VwDRzgjyQf7K84PmDhcpP7Qkoo+x+vii+a1DyqsnR28Cve6XPOQM+eFEZu2w7SIZ
HLyH89/eedg7e+mKirBY/d9ok+2YepjgpyciiIHsJ7uEqI3CS2w+2TbMZCgju2AG
XuMfRo84ZcpgOO5anG7VD53zpQwuX7hrxvxKMrYM3DRldKaSVWJDJU1wpX+xVHeV
z0N6rvB8+CoF5dRGR9jGsClXrVzIJhke0/Uzjh4laxzFProYlwcXt0WgvsPBcE45
L4h80SV4heQSl69ldYCsR313ALKIchYbWKW2tk5xQBRViguv0nhmMaoUN5ywDt7L
34FmDKHt1wek7lpzlQ8ZlXQ2hWTArsKcBN8Dx/28kUoQ5GfpDRT0tjqA0h18veng
Yw42SthP0iQJW/B/75CUscYmnNbgVqBSf5/EkRfn2SOpnEzNXVtPLfRmJpDMM1Bm
0qKsKkovw0TuS4Sxg3vND3dvdojgp5k+2dLulI0txA7AVyAs1XTjeeLMKPsWKi9z
B7XA6IS08s+Aw2QlEOdXhWNw63M0umkzGSvqYW5U288AOIM7AdzDS1NppQr41Xvs
GTP68byzOc9JXbbEHSQ1Bnu1vU9lLVjsZmS7YFr+6B75SKK1lqMDiqcToNcGkgvt
BYJebwfzoGDRHO0beD43mIZjVDnfOSXJOdL1kfaGno1J4F6ce2F61DGknMpIM3dA
fwdgz6YLDHoz5MMf15JUueS0y1ajTMWByS0ihUrVNd8IQxujAcxgarjJR8NFgsOd
xB4xVRCEPCzqhQe+LdthaqigS3FbwG3EwMAzlOoz/7BEJvMuF2zVbnnblVNWmlRL
4QomEiXjRp9HNzoEx6FAlA8RVJVPjERIsEsBdPo3j85l9iEnDzVWZkfJnuIgOEK0
YE9R25L68kJ2Na79r+e6kbk/kRmX+2xVaEuQn4WwYhsQtF1jx2CFKs2P/UpQ+uTG
7RXHXQAF7fHjfo1VyLuH6LG1HyxmSwI+T/uIQdkivKBq0XzZW63iEMY60uZRKi7j
nDm1q+Oy09cSu5ua6OpwbL9vbkUwwfGGMYkWMub6E6U8bOIWj1NAH2VNbOv/+M6y
eYYS9Q10+mGMFeWrVD5Ez6WZUbEXtcoOZonK00EaA3aByYR4qQoHEpES/4NSQQAN
X+Gz7TU91DiniVhBRkL9R+6T4i9xHtPZjiMR7JrbfbsMLsCs4Z15zPQJaOc2DFvJ
nTw8pqo9ENxcIvmlEOcHmB8Y8IxmvJUZdCc1BZ++PzWYIseLnKzAauOqqGEhAxKG
lF+dw/dQB5WPJi6xIzT6MzuNfQvRDkYuG43etjSoNa0lbsWSRgxVC732gXpKgPxJ
iCKMsWJ21hN9B2l04/iHJz4rjX+CsmMcDydB7MwAB8XGAiINrcWgNPhjYkQeRQsF
eXDQ9+8yZiEAgfIqNwIg7mlcF8F0kl6REGZ6TmLrX0OHs2H2BELEYvBm6jWxg46J
/x3zXSVORJZ1pUNZuO++Uc9OfuVM6Ds4FqpI7U+LEJD4uDsu/fodIoedfTTis7Rg
CjCSjmiI991BUWhIvJFIP6UhysU33QV3NOgovt0d5fiVgnAdDcJifW37963dOfdP
6YFWDat4iBeIfeqsObLJd0OLPirq96E/mktfsfmwcObp/dkVSkV02/GJi3dsXX4z
92zqKnCg1EQIz0pxmoFNa28w0kaVOpWYNMs7zcTIz9dU5RW1DAc97wEDqG7c/Xc2
o8I+tE6WteBMx5ZkL0Wy4dhflemfH6GAwcfUfExqdfkWoLsMY6VU0FqfMSrh+rIZ
oGkY6y2Pkkc9VXH1888EX2xidf0ns2kfXl0VJxNbNIvl+7NqAH8DT0VTjva+7TNW
BclmUIufea4D+kBmrBZZGmaXJsekBP3y5bNGDSIvzkLF+poGI47nXxBYOzt8ACwr
Um9TPDvDVL33xXsk1F8vQBf8seBJByv1tIXCBJsVQ+Z77yQCzhVaL4KWBkmLkDiM
aY+rCw8inGqp04TDauhjol1GaeAom0xC0ZMqlNf5s67qJ71e84YwVoyuu63YAk8G
UfWol7nKXQ72O5EW9efNjW7SeB8LdwLykuw7vrtkyYc+LT47FrD28By5ROCAiBlM
iq7TAjX6xZfmWnHmVptenTgiSRU/boCtI1X5Tswvz9Qkf5ZcI7GxlrAp4Ka8s3W+
WoRlyc13eYHgZ4WIpsccOAQj3unO91kFKRXnjhBuhXYzjIyjU2vQRp2C8k+6HRYQ
IPW/2Sc9YKgp6ypK8sznFSTTGhBkDBZq0dSOAXJv5SM24t/wgcsfgme2e/9p3WAd
bcK0lfjHEZEWbH5d8q9y3GDb1ovYiQN77Gv01K2Vw+mQXE2SNHU5OZKJ8Tym66rT
69nM3YgnpQkUtYaurCWRNserkwVBKXJP1pJ+xiUlsfEWTOnlWiUYIo3UYHCeH2yZ
NufKOfff5fHNlAwGLmy5nA57nshKlvWDST8IT6EWFI4mGHgB6INlEUOUjrBOi4U6
yeN7aXg5Ov5RWYWIUi1fxPMcg/Vet1FozTn3B69gbdseOPlEbkveHhsDJkEm6M+C
piNKrCB7zJ/c59I+E7mRJt1UGr6VxRAYo3niEl3WeMMACI4nUdVqLHzbRSeiQVC2
XNrlWEn6KSwdkSE7Xomv8B95nPJU12MC5sb2O/kfeBVZ7qoDUfu+aKWZwEOcRMpC
fTDMMedildm6htdyyxpKOphtWLjVGdv/0TRXUQEnF3O7Cl0u/TofMR0GNiVxZJbO
rMtkcyRxFNs7VEfjeWKdPIYX5ea1qk0JfHRdWJ3d8b50rZNz9f/ZQ6ryviW84Uhi
Iluuy2997D49LviTEgg1p4OvmjqLd2bqecwS1IDw/h4cuDKmKAJRZJMNpNJOx2Eb
dKfqvHIGMNwaBtKXv5gX5QPzQ8Ek67P3GIVM1/njvtOesTBHjoQlUGMLwunDV+Kf
x35nWW0c/m6HObdDJhQJ1nfdSe/W6wFADv1ZpuHlMRoLc3k8+orBdHKfu+h8+yDU
+vx6vl/bVegxH4cGroE1gOqw1mFUA4YfnZ5m+rB65fcpGyNp8rAnGmyzwoebRTmS
PSry71/i6kD2wBaAQi/UKP3niMSyb1fRWmrxf8E/kSSbhikjdhEXyoW/kC5ijlg/
Ho1aXaB0wrVzjD12h3u7bE9NOEeyWcq5T1HSrXuDTxtcafCdRsClbKjeLELzaonK
PWV/I7mRIUtehNC7P8+HD8oMpn67zFjtzQ2Cw+133IwRWYAioOakCycGnKw5iuCv
VN3X+NNBpFXQlTvAfW3WuQW4+sxToJJtwJahpPJCN8vWgGBx+mgXQXZbcYa6HIDQ
eUVwTuxoesyT80jbBWQAOiMQUQ+4u4a+aQ+FZIJYHLdnkHNyRnaXx1Mlweb00lr8
3uPL+IOA29atTEPqgi+vMDEOB9DJUfCkJ+rBYbRCz/VYDnOXXIFF7IMu0jc1rwov
emUBlI0ATXSgWYoqSYIDYMcjjfgDCt9PrmW096pHa8lMTqOdBeiuyMHOOijLXYVu
6ahfYsJpOPNSyVLfJPmde3fZRtugO9mnT1MIVCsHkEUKbdDVUD6hOHJ7BKbRFrJc
WCMAqWePXtx0Q87lWPATtPgpVss+Yt6fzIp4El7P6DYbJDDa3eIsU/Hz0bjfQ/qa
5x+gM0C4b73Sv5tgPaheL+yi47jKXZ1y9RFpQbJJpNSTbAKhlWjPLuzriMP1uTNf
RD2m6QhtXJoJvPmjnU8ZnhiBwQekdZvSEt0fSWlbN+F4gXVGE9E+wnBm5/iyII8X
8c+6h4HylKTKAYfUoSes7hnBDk8DR3x/+5KQX0tJLKQKxpztOn+NoyYpTj6Z9cY1
dYFRPSsihxLZ/WtiPW/gfeWHIGH1QZ97japmmZTgP+ozL2mhvMlxFEWd0sEuIbNT
NyerfgCLjr7ghENAtOauAy9PBTnShUamhiQEIh8z+hmABhnKyuDAYqOecVYqj7St
WYIQo5lghY+HhADcrjt+RxnCFrTUDtL+xMUjwik4JATyQa9JMqxZzys2qA2AcHXu
RXeqjIyXca8wa61D9cmVAFLHwl3q0tuBypAwibSDdnbVCT5mFbrsoKqJIsTUV2nx
s9sRjJenKyoT/dzSGkb4JIUYA/GdRXxLhtpwRy9o8psgYyAPXFpohUr9Vdjgu/uE
GHxyTgYD8hOaclFlvZ/iUZY/PhtWT6+LJaf5WbUvqu5ydKzDsJMNOZs7J0pLco64
D1fRS++UFcWi9PykozuylphheaMk+gYHSIsRysGC1zCAxO/ZWZcGYLqE5r+fGqW2
k/RkhMnaF7fe2O9b07hM9FyuODnGeK8Ssam+2Rc+vMIUYkBY9tFhy+189sLMxDT6
odiKYyqB+P77+M7L1jMIZ5DLq8Y02bXabwUA/OcNXmGmNt+jSSu6CNm1gu482Mqb
pIQTOj/rfber+SfV+TexaE5WWgxdCWN9U5Ju6E/2PSD2WpXGBNaq6B80D4SXMqtr
MO1nZGjSqQiKp5AFAL2zkzJfLPN1IiqEeNBtEOPurwK2KJq5HJ5THT/g4XW1MNUo
U8ApgDNqfQNQNeH9ptJtLe0cXFXeOpc95bBcOWdZR4lf+QPvlbrUTTdh0ECQwRli
rt31ByL3mAHDIwnRYHs5y4pcMZ+V0eCNnKtUBKsBL7nd5jTOK6esbJXf/m5T3xSh
CBJjm+TmYtMLKY3FM/WUkbC7seuntQMrcpWJPTZ+7+tChgMVE6wJnDbSepg1148s
QzxqPIPjPpMF/NFI8DNLMwvI3y135D2j/U69hipQY2LD1utUh45oR5YurthUNFBj
FTGIl+0Tx9lL7lJ7ShvcI4xpU5CDgY9/cFackXjwSJM4T2dn01jKjLz/aB8DLB5l
u9yGcCnNp9FI6Ozb0mtS11SxG2hfG/fqUMoheFKrRZaPLNfg432WeBiq33yMKpc+
X/pNWkdXrPGMMoOom/nLTmnfsjQep7B8W292fiNNq8uC3oK0f5RzXKviq1rKXrRq
nzcdvlvHKKJQ8QF55cDQcxKmS+0bm+LKptMgH3IE5RnCVm5qNH/TQXBQZUpxeN5E
kdK/MJRoodmGXC3wdjNcKGHbntn7iIrlxlz7opAdo9CcgY0xFlEV5CK8MsvDJj5E
3SJVYh5oZfUNJ7SchU01kKXupg1AEyFSjBRBOcwcvMa80iCEEqD+MgGkE5xEDlCB
7etwFP8svSGSsJPK9n9wjizGCGj/6BsQWg6Q6PduyygP1bmRzBcXuB2UVzcaR95d
gWP4h3EyOxAhXilY9ARM9e0p8Ej8AuFZrGft9XgR/lExpdD079iyzQzbjKDmpyXn
d2dZJJRq2PuDxlA44rGZuesosCcnkF2JmEUHSJ2Dfqzzs718l4e2xMWXA3GiN2U0
Vb+e+GtQ59eGxLp4FKPL9juLLeFAa6z6ScrvKDs/H8bOXIaY1vPed7aAoSDczPnp
QBMSsdCD7zsM+WG18Kdk+4w6ikSU/cTSq4dVEh5NpgbK68FijsfuoBMi4aFLR7hh
3jXuAHwoOv+UjIKdlTUs8Lm8ioiYUnvhEI/AJxyw6nOmt8qMZyhRcp30cDGdQQxS
+EDv+oSApyoW3n4Wf8QqDnaLvziJbulwOfAWUxkYgHZMUtoalDb/QgqpoldXMa9U
jpnscUhHCBYGfD9Kwud6XcWNvUi+0Prd9KdnV7QVnyHwicfMYD70CjK2WHL/lbZD
vqQwFMHF5Z4qsWvq5SWLkaTzFcXIcY16DiouYwpMglejl3WXcGP3GqmkmsnOAxSh
m1N9s4mF8VpW22DxUfU2uVbFpZVJ3bPh9wTYyemNE0D0r8YeT5Re4p/NNd5KtGGz
Bu2WAWysSwRdr+fGpR4MYaAzmQcCaGQs9xorHOqhJTDoXfuYB2hoU6vtVw0sQpYc
xGvmy9GoZcWddSuK0scypL+fE7XrRKO5fgMqYOKXp/D1PxXWK4uPF6z6cd4i9BgN
HST9dAWNe4eRha3+SExjRy0ygBqwxF/pfHyr7h7mUOTCTAfbnfJouNagsc5ydLQY
pXH1/SW7jO/VH0Fnwhpq1p20D/fCYj3VDEHYbT6aheGGdE1SLgLPDceX89hJHqLd
rnzhHDnoeJRrYLvAFETO3bFk4ziA0BUZg+5OlwS7yhqHe0tbuA4cUyjrMiRVkcY4
i6RPGqDBHSX/wA5Lnzsseo21Kbxnhgf3DUnlDG3pcgYcdVzyS/qQAk+K5yHVSpY8
PE9NUnovEPpbJdf6OmjvadeOIrrFqa70VZTZligQwdzgOP1Ufub3MY8wuX/fIQ9U
SMXVKMbIR/qjeg2QRA+EtFrf4r27C3NZaoxkd1Q2mjIKkfSVTTZLW1LNAXA4LwvB
g4HEOlnsLLge2k32va0oaebdTXVBseW2pXkkQWW8rZ8pwqYC4bkxBYk5qw5UWiYF
rme1LtyaPmi7ujql82iZu+vkb9zAJYxtPoqJ44HRmFZzypIpJyT7mvisIilxL2Yj
fySDTiCzRglurYbe+wT/6q4KBEdsuMOeeEZaaW2gor3ch3MmbvBjWoNqAMrVE3sl
+SjOeIH7kB+QF1so+9xwt+4PpJ60jGg+R193ZSAq8yY0lMmpda+336UeejaBJ2lF
+8BQajs2vawazTieuLltQedXU76PhH4vNEvjeBqcH6IrT9uiLXYJMDHUxE7n0Kaf
PJHN9iCR9GEVRRRwxk4p0klLnJm9T/pKKa0RxKj48JC4J9I39pjvg8tCrSlIJDkZ
Ce5pFXHy3aPkcUH0QOWwRrMDasxNu01L+AQi1TfpAHAP5HmMUriLRtIbKomPk85k
Pr4AiZ4aj4/3X0K6lLVkVmaEd0jEdUqpFT3ZCGMzRogXU79zgiMhM1EPxXuWqXGQ
DpvfoWc0t38JZmEfqQSocm0vjUz8nmKwfJzed36t4EevRZLLxCTuDOAF33Z2Q0A9
uTNfoEAvJ2GYVtCusHVG8xKSgKu/JsOap+JSNRPBBT+hR9k9R53oWwl5I6LDwA8f
HpDBbminV1+qZp8sanxDUbgBvaaTsVVWxNV+R5w18vQk/kSmXASJA0gWD+1J83+/
bqitBkAItwm138sothSCt4bclTDvyU0AYKERs6Hkk45bmzDpn+Tml5/TR9ne5kkc
UKR5PHN0I7iHwcfJYSj0bQ/vnnBamN+rAt1Vp3teso0jD7iEvwXK8G3MQSFsDMOy
IxuDMiWSbg3MkWEnlpksOmMpROWJi7SldQbmnPn6tP+QKYAZcVwZeZ/iVJ6yQ3Zi
+YN0qFjqA+vPtOXwL1lkAaLQfJk/6AP447pttIAUwe5BXKrxq7BCm+4lSIJH9UCS
sEGzUrr49rwt74lB2KZI+tvd1oa8+Eofsth/jG1M/Kz20DAW+PmpuxCw0PK5jnBr
dhzyg1Lm81WkxtDmx7+nSFjPKHVhWg9dZqhFPmGy8GaM+VyUiNCG21IfCN4ZHt57
4Bl0x5nx6ImDVSS21BcP4Ua6njQO6gINsn5o9EQQ6AROdbB+5uvJ/jWBwh7+vrdc
NLl9WRJ6zNzb46jmHq+hpRheDktmDh6Wi2XCyfwxkFSFZ2QZu5mTezwmMAwcOAYO
gNjDUCkaxYIrtHYW0XrmBHohUJAZN1pI8phD4Eilc1/mQP6SH/UvzLAWsMAkmjxU
tGqlxiaE1a3PZ7A0HKu9ZZuVDPkDUgnK9D0K7AZ3U4zelGWEuRVJvCUFIkzwKcUG
5Ju4PeAwonW6RocTmQIY49BHW9K+Ezn2Umy/bW6cOBwvMy+DHgen4BxawaHMUHo/
2N4dUaD3F13kRxJLUQ9FrynP+yrYMOS4r45txDcM1SlxxWsNBYM3xkn1qDmxmSu1
TogUlkm78nm2qdjNcarPqmdmA9vYFfqITZkphluShQrvUXMSLRpj1/WCt2uhSI2g
mOnImTCFYTa1iaMzLbjOQsVM2Jd6fbd6OjsDFUyjQpuuOuzS1neYWyhmJ9dCU79K
AF06chZemCYuMRqtG32t6dXUtrrtNUdfv5GEf9FqvM8Q7A38LgO3wjsOCNRuXOEp
wEFPuufqDJ7i2ULdabU5sO8n1XotquI8QO/av7hfeQs1wgVp9mqQczE7LMvxov3T
NwjXSTOTgZNL8LO4roy+jEvQnvPVqwKQHKja+OVUkkuIcUmFId6Y9uloaWta6QqJ
fBATsvU3Ro7jCSsMBqb/9+yCZ4MpxSgCFhu1kSQQ/7UUczdTwJK6pJ2lzLf6UpUQ
YwXn0npcVak3doYr5nFMzFjdqEVHLCN5B84grts7A5tiH29fjpIGypGQYD6xOEE4
D2+/YSCvRUqZHKCNpvSzNKGasvfotEnqSTcG7l/5LVCwa+OUGQEPT+WiQYw3L8+n
mthz12CppQr/NXAf1pOkfbzOYGNHFW3vIxZ5fy99HIlHJSrlzYs6gml6vg9zkIiu
q4yKUD/yyrcEzRoPhp1lUK9gF7esO0Ww/AzSbjTeUffW9ksvrkFezKMm0ZM6YJOs
c0ox4Ipl5DCrJDE+Qtnv/cSLwwz72QmDyCSnRi+bKXgfe2U6YJ99qZRaV5xe95kR
bFgoLffFwzLzR4O407kbq/oRzrzHPZ5UfktPZPB5c5HMo4Dkdw8gzo+YB1stYeeE
q4+TPDUsyndwCBG1Jr+IeJZ9do9dz5mr6nNaW6GaijUKyrcvTJnVcCGxuxr23Z1A
v2PKPLDCggT5+9RAYgezFoQKDqhLoj2ILJPFnUZ793ALNIgJGXec3IfbYjFFXfM/
UiPk362UjKtymGRQn5bcRtbCdoTpUaI2R+rv1x95jCQ9vouJRZk0OAb938a9HSkd
3iB102vKyJm9rZI9nmHja48qR76lpMW+pEaRpXpevsFcD96LEN2bkicnHRCXlySJ
1dOfQ4eOtVxnlcZtQCEEzw9xwXZxL2MtCHyYVV9F43LVUTMQMGxAM4O1NciEPmIi
uS66OCQKPAimh0+r2siKCYChlaATLo+ZiwA7AbUqfkFl/Yjk0GTeL704fQThUkzj
uDdOrwzrGS3d1h0DlXokqc+h2sTOnY9G5RtvqpD1DPmDqcLTQ7c8xm5Ln074WOIl
r24XQSocMThdJB3h60SiQ8KWnTZ3bbZNW4ja2x7FdFVDGiFm4/ucZLFVseZ8EAMu
UvQJouKZZxEmmX9BCb9dAcVPXLxIKPlQ61u2CM3kjQlExzLCY6MuHTv6huO9XohQ
vJdYWtAIiZSYBA7UCxjIvPA8wfe89z+Dz/WXlvYv0pChMK6Rse28H6elr4MyOOt7
pwI7tYLLGL4H3n5g085Ev8obp2NQPZwNEfNYXsyZXB+/pQQ8/C84srDb4MGlIpVZ
sFO770FSgFKIvTCjOevIIVm+QMAe2l90Tz5zfZnadNUer283ReL2Ntq6xYOc2g/9
6CCMuyBqsXWgidAX2MfQ1roB7MY8w9T7r2iFdViEZsPfZMNBXhwNw+01ZUTNbWjr
sZhkv3HaDWXugk56xZpLqDEsrXXBsmYGpPyTeharnjLvH2FWalTdQfRxIpamJBz9
jbMXshzaXg+6I5+0t2A90tT0bWxQb9+GTcZxgHDA/sggozTFyk1eiofxQZOgOH0l
acLq1ywBC9/MMcZBGQrw0A62FEiJGkougQn+0st6mHMu++W6wmp/GHAfy8YWtEcO
6bln/97QWaUFIJGXlUy53p59gEZJWq8IPq1jHKOgsis95CHXTs6wS+gSoP9ubJ90
3Pt2gUT7IOmwqY5UrqlxCUbIPjB6/++SWwftw0BVAHTHOfYfg/GX/rmRV5zEDczh
LxGGAzCyDp3r3sjumOn3eJbXrlRk5uRew9VgBHJvkDdyn8bxx001s5/feCmr6oFG
XaUiAOEN/ITQHZ3CZBh84iUKrGRqbgZ47+OUts9ZbB1WNyvN5um5PhWh7sPGtGsR
u7iJny/QAq88wf6lz39SBzjXoDYFQKotuhk1U9N1rMq8lQAkWElADIVZY80OGiVV
JuhYjQA1o9xbU7/7mDyzbBBT9j0WB7G+Mwcdfq7YAgZmGM+4hKhn0B9ZgapsOipg
4ypKPE787nvY6q/6jZl6nGj+Ht1/OE5v1nOiANAO6Ib/L8zKuVr84K0hAfxsYnLU
vKRgmKNnRFvFCiQj9CwRduL1NA8SjPXS+JzZeD1oi32rng5xvJTvo5QIUAwAZSyr
U7Jas0zjD/m7pTe7SAyJqHPQjXpZXkW4yoSgmYBu+kJB9xIBieV64LTTQ5vvbojy
PX2Eb/1O6wCsNMbhvBC9OnZgy4VRO88hFfVNwI2wC4zku1575FUP5VO4pQ+0HYBW
DEzbMhNfKgMglYpgpqauAnwKA6Cj3W6ZGkjUhzMPahjRRuqybn+5hsi6se58b7b3
Vg4IQW5BpzVpiqI1IY1Gl4DMRmHN6zHcLiD6GRSIJ/YzBp8civZwKEa+uk/pbzir
bBGxI1ecidMk+4okR1mLCDf8mw4XqMo2XIAG29jd+VvbMGI+TNa2cOIAFMF6OVWy
Amu9t30TYtKF6jSrBpVkVD/C+cCJ3asRHWGotk6jnUvNJ8tU/XXVXmKccqgi5y2n
4zj3Hg6L1KjMer9Z9yn0PABXbl4dVCPvzI6hckEtfGMu9VfUhl6wyOyGhvReRmtw
iLUzNMrQigJ9AFg+0x15CrssSqbBX0IYVoybK6zNWEraOhk5NVpwulSYCRK2DW1W
Qpbx0EPLIPGTidwp+CT9AtifULDJzva/O1goZBO+BxeZ9wsxlnC51PEoQO88IuqD
SZP9iib92L0qYClI3nw0LkiLhbgqzAne9Io8DOOnJxk6sUvzDr9ISBsaJ2w2AbnI
EeP95eigyHabsV8sy6loP5yHSDWGjz4SpqFFKcp7H+3NTcrHE5Jq96sShbt/gWpD
fiK2zxIjLj6/MhKkAv4nJzfrHsJ50+NIaE0o/Zyqwc87xOwS4oOZ7hzFK8G+scsI
Z9j00csGbseV1oWzb9OxTXf6OR28gk+tfv5ywwttrGmcdSMkRNAJuGi5Bh6FvsRm
klCT8DyO+kSTbhMJ8u1gi9Y65MGQ5pDzbo9UTzF/CfEUPfuG5RY2iVBJRw0lXRhU
cydW/e09LGFz8Bwm2zSbpeyFCjsHaV8SoLlwl1iVpQOapzvZY5O45hDiDH8LwK9L
+WCx56ToFNal8Moom0hOHkPZCxARMdwS+MNvJDjnupNXtnQd8hj8oASdL6NI1W9k
LTfNVqANsaZd5g9Bb3KQ60IER4IneGFxl5Wn3gkp6+u4X3PIvY1seJbSx0xuXZ78
qtjqFlLFcOmHMn8N1Xhket9JAYR5hwQE7rnMp1AevfVh02B2Qm9AiqT58NJbfmDa
sYl8Xi3TM2f2NdYCVdoXTDaYEV/owWS0bl7t7vpie4EgRAGsCeRYZTmB+CgReE/0
eTwskzYPDqzHvxHAWPkBZBg2/+t1O6JuQfNazmy+BN6fvA2Lh47yt3lxIwOc0hU0
EbMQUIQEm2jVZJd86piC8qm63o1qosQfqXRB3xLhHWrGA9i+6K3W5i4Qy7ELu+9K
EM6fvnYr133PCZn+i/MAm+1EfgzOHJ9tBo71KoMOIGc9QeKuqazkDZQHNhBtpZU/
sZ+lqPrZz9P+Myqt/912iwsAghe6M1UgwlXnfbmIosUIwiDkzNth4a6LfUjyNewR
V16LmFuj18PXlNwrgLFJG9KClDRT0wEGGxoarR8QtZohWkXC05QQR3x1FIDCZBo2
Ke8wWvl+2up4uIp7AP8dtwdk0nuxuvZ4sAp7u7++32RXjI9Ffjrj/se53ziIyOzk
o63qYxNVe5Fb9wrcJVTUbGjT5yOzRXg/3vK+DL382ejRYam2CuMy2Hn65vRG8jti
qNO+ZDTcz0AkGA/YwpSkyWs3IsvWhvcCbX0xgR6t55vcSHZjBO7G5WNsUa3u8VZi
KKJmrDo1UvCGwjWLF8554Db1OarG7fCCBxgIm0vXkvKnwuawCYxpiz1SbtTd7rWU
mb2C4FWlJ3zfdu44F280eQrUoqjHTQpUcy4W0wQd+LxNShM1cJwI1YYOHKIu17Rg
Ip9ZOpMJ6TW00/39UVashFizaHwxicqTyPkveo+r/0YCo1sQgA/qXtNldmf12PQW
tcprrYW0xyk5KjMwEsSxkLKKW+YltuuQc8RlkNI+HGeOnSgY4OzBEfdBIW+1SQvf
FoGqDMSn6/9o1M+BcdsA1zB5+ADpjefvnG03sUHuwpNHWbPQAvWAjbC2aUiCkMzE
1jRubGiep4l/ZciGsUJe688ZXwpuCiiH6pmounfqtpiL1IADx/TMK1BdiR9Tzjjx
f8kmhKm2cbWfYVSpxkBybgznrY/23mF9u7NyqxY5+qzSFVtnypA9dXFFzjqbN00a
j6xZQPH+IcTCqX5vVTwvekyhq27aFF9YsMk1yH81XBD5o3+5fBu527+uERFBW5M4
wUzcDWTPGB9jwvwNKeO8gdU6BILw0jCTw/FxrNmIfcp/Tt2xFk4O6fDFdOPGltPm
VO8I71BMHUAj65BIsFO+34ojb38lfxCdz6eivbRk8LljIABacebbsi4Av97a+7V5
Fp1I0IyqtO1tW/0i23pPjMhd/16RGvoiMJbo6UoPoSIgP6cXjvx7MzgL7JL3UMNY
MJTdOWPYE+f1eZY2B/yv7+1CQ0ov+KvSuAsQGa5hKUAEyue8JxpbxVRUGfGuLshn
eGI9n8FozUuip1KYxHiDc0ODNwJyyhy5KTu7twQMuBaQEi80iiTF59chQZKElhVS
mG5OtOl4dEM54Mc2K3/Cohgud9MZLcXBn+Ihzt8RmkwWKXvZGIRFtXdy5mNujDvh
Z3dqNVBx8q0IThljQd0el+T2DixdmXh8HFBFXZjVOePqAeHc8Y2qIVOf2mrkjbkW
8Uhr0r8oX67Q9bPWnMUiNiME9F7zQrFP7SJjJjXXLLpImDTbDa7Nm0PUoWpa0cS1
s/tDXMqvZD1zSVL66hT+paffFL7dupUL33gVOwabZ7clGBPCZf7WzRaS/sfBhw6J
C1vGRKOHPlFTzaDZxDSsd8lKz1YdY8hEfgknh364cLepFunRyqHhpQAmTC0FbRwQ
PjRkQy64+yvccfSjWYPpKl6gu8m9rF3rJ0Q9e/DiG/OiD7rDsVpxQHcd84q4s9pN
eDgCQgMtQXPx83H7bRiC6cmYJ4YCZGDLxSdCFuinJbJf8STVL0fyhty0v7ZbWjkb
2GYvqVuVk4LPJW6F60VBIUyNEEKZeS5c9SiZ7TM66FMNT638Xt0IZtHgSyDnT+XQ
YYVkqsqizxoJzDuWCRBtGEnwlcl8qfKfAT0mn/KXXzy9DbSOQfHIYqP00ZD0V6mb
j6iGCYlQUMKVfelylcUT8PwcbcNEri7ZD6ju0YJ08gcI66tUMjDNPld3w0xjCImN
zo7zw4xmHNjQNKXpnjO3u+ohha+fmJdz4Xom5l+GGwip/lYl3Jhz2a+h+NVkazSy
4QCX8B/SRstxmr6hn/rWE320ibtz+gy8JY7ubXlPKUePFwbxMI7ZWPlFi+BDOOSA
yqV85aKjHhTXvOV8U0g3cIM+GI6MC6RtJiIWJYLnb+CYNg6UlIr9dvkjMf92aAvx
IjwpIxct+a5x9OW9T/EzmixZwIork8n0JgujwXrypP+PgAF4QnXdwHDGH8dIb4o3
Xb/g4DnbzaDej+G9E2xeWAilpxAQE8eoDqjRAL2LqIOmfUOHylyYK+d9zJvAgMZK
UY/64q5q7P+666Z64PHqahqOlLC2VNoqDjWjC+7r0RvzqSZU2tTYobgGcy3NxpZJ
jeNcN+6AweY3BlmFU/XdYwSFrYlRmsFjOUdNTDB1kAqCJ2k2bUKy2a6OhlB07ELK
tLDn1+KuQGLHJ71WojWI0mBduOqjFXDNxhwbo/2XzbCut7d+TKK9Ze8X0TcXXlDV
zOmsMhW8GIOxXGTZ5sGVR2wDX+glpVxv3voYYIMfWhAmM5hkp2DqGc5bERVY+arv
+3BxuWxjLy2qIkKZFvj8x85hZPvjB80Xnl5QPZIclJaPPtCsVWH7R4wrpWEebxg/
nQcSjl3EGX/xaLddHXD3CK3ZKDe6qpy8/zTs6AEc+cQeMgbiqyfTjNtkdtnBoU1q
Da6ANs53T5JCSIZ5tnXrkn2Is9zK9qpiPeliIAy2tI3NaQp4m/NKzK5bX0FJL/RI
eEsgE9vk+wIhiXN2EHl9SMod1wmc3vV0J48l9IQnWDO+4UW+xAP9hy3YLJPBu3+b
lndoKSFzwBgotXmKxJCKHeynMpr1Nt9PQ6rHAJIZP0cEC1eifdgOEIp3a798ER5t
Pur36OeHVIUljnFJ8Bznzih0J+RdFph9zaVEhMYRGU9zLcdk5pjryohCa7mVu25F
G3cGlYXsj6VUn8EBF56llRjTYiIG/4ygnm+1JpBty4cWWf2/WZwE10xt0xGoRwn/
FvyRFvBzA61qaKVsxiwrA2PkOypppvcST9ng+WAoZ0FqW52+6kPCOMsoNPAlhsg1
44aOt7llUK9myt758wElz9PGJqxju2DdvCcCMijiRXmvBfLUxeLs5k9X4WzxVsjb
nPDrViJ8kwaoF22JX2NbEHkyU6h6K2uHbFV0V7CTgII9E5a6yWXTtyNkd/tS8cJO
OY1A4/9KLyyQrjC9lpUqClIPBg2wT1iAWhcacuSumHpg8Mgxzuar1DFit48+aX/E
zjSwoj4mCLrUhSB7oQdw6aWfhmoU1JCuRCpabZ7kB1A1po4TDFXzkPEHdOpYO8tT
R1MZeGzUXdBMefFTLN9/vbnzeOGnt6kTEVUWrtDMhDUTBb2aMeHFsslmsQPx4C8b
dL7pr27q14imsbJr+KGfX6s55vXVKUEOhdZMQiNjeOlObKwxhSeTqqFrrq0o+uZQ
AgVyg/EnJ63I4dOg2j/EAWqWhyZdS2Ad+POn6kGpyGQ8G1zO8LPBN6mDbiXcPWPj
XN8moouKcafDV/ZuBT+vuH7b4NwnpYqx2C5fxJmYrFSPxoUL+6VOC8H2v+vo4jDY
swX0tIlgP3Rd2zc/VbAdMCUbqpOoGDRghvoOoBZ5I5c/Mc783XceMAgucpo4Pi9L
qICvIwi9G+UtMIeA/gTS8mfGOlhUyEasWWvgvsaH5RdKS3Cb5tF+gRNXOuM4/v6i
cgjOpb3HuXLR6piJ7hnH2lz5MpYfyB7qvI+MgRcWFgIDmFs0VM7KTnAqyCc7NRJ+
b6z7Rf+bdKT4qQ9UYaydwWUV46Gd3dyuhIQr20QkagiYTHfZ/n3tWBUEnSr4OayA
f+CFbhkJMDPfS55r15ybuOXrjNBIdOs7B52RDCGDfot8Vib+N44FE8v/OIEvzgV4
DXRR4PYDpb0d7b9sVrLMnIezx19Milmyq6dCSNznYWBBeDGtBJUOnBzW3fqNodyn
mWcloiaI2lbLXsnII0yUtPDRYviPwOXH74n+QtrmKb+NEWDAPmy6jmBvVrhQQLiQ
KywuPxOk1OqFVux92gsiI7ZftDG+H8B+mb+GNAbrwL01uJYbYBMqun4kx0VI4JJi
LoUDmgx0zCLP4hjeua4oNIQuq7Zn/dJqSYpFCbxKhPMQZWLCTkx3WGvZegX/JfhB
+xnqOtCXMuH48AjMsmFKDbaI90O0LOFWbVYqd7wXUeRt0puPNKmylmB98l0faAJj
a7CS4OznKl8wvK9C82v8POizAmJHOjwRnC1c2j3NNoT4TlSekDFnVdLXe+/TvoKn
lsB5an+iwmq5x+/32WMA0IPzXdWiPMhEwGBHh98Kf5BNuxk/KsPKOpa4LLp0dypP
5MzLB4doj+ypqKP71g5XxJN7N872hatgq+WhgRiwAguSgNQExaC1qNV2vqVYcFfi
o0tbO78d7CP73qXDyjkoNiGJ4SoxRcyPsnkBVry2bh3bnY1q/KUBoQOJAD/WrogU
+enUB/sEMMqcUO0+5rC61eWbmN78TVYEAb/i+DpTOPGjKHaseJrTkNE9fTQPfE9w
X9cgF4DyFpvnw5oLt/cfaK2HxLIepFQIMHOy2B7wViM3oAYIfi6PRYbmAtEHy6HG
qtJeTjFoniZ1B7i+2Nhm4nW5ijw1s62FnyPEGoIapfbdbZrM9uvI9a/aM/9yD1IZ
/20jrog/gSoM5bSJA0wWVRfsuWzxFXWvpWcSPFioT7ntuvip4QYR2E8z5I+wD5pD
FdMsm7CRiAEO0oP9gM4VV72SLYZt1Evun2oua/d/S8JiFoDBx6z1nWMtimYJ3cGN
flER7mpiLXTvRuXPpf/BsoRnpq1npQKOHkBRjwiz6WM5hvRKOAvB1ZPr+i+M22KW
5j0IQX6EOex9dNC5JoP9H9vQp0amIBW5wfrp0kDRytTPHTWA3DQfm/ZTl4PrYCx9
+ArjY5U/YK//4lmLfj6WjXKLehla7C+3QbmjxLrto4RkcOYuj2tIjZ9KXkcrg1ne
AAGzL3w5rcoITi6YmOAd25uOo6WdxHOoF4DBd5huTZQBBUqhiY+jh2w0rYP3JWjE
c43t4/1/7/86Ovi6TO3ALoF+ElUl69XmcnKMdmKnSO2TBg23Aw07fEDkIGTVyB4i
Ck1aM5GhxL4tzqXWeP8CQJzKfr7MsepScLreTC6mJpHwGSHntVl/suge6/euNMMX
r6Fw+e+iJyErGBNEOFhgmLK73kbhXR+hC0j1jitcCMqmXqlwVhrnL2SAo6EB1+C0
F99YHiyE7bhnbK26gSlsJmXGZ1jWAOu87/tVCs9+D6oK5MfJniwFKWv6EAfUeB3Y
M0GScGkJNH1M7nm++Ifbzi5rV+6C/6b9OtxQ+rPaWKQ+RiivP0+loXJn2OLMD0vu
4QfNcmVdaQxqrybf9eGEP7bAqFW/nhYCyLBDicycYKcT+ci1HM+0kHtXD8r09TKa
e3fxnKVZkDPmnOXbikzN731EgxY9SixOeBC5mLPsoIoz4q+oihgkqDtOtKoFgN2I
rUl6lwEypgJUW1IZAGWHQuNJ4M6YoRSzO1b2Out5m6mb25nA/Uc1I92lRkWO8eku
uo1o/t6YZ+fXVo2Zp36jaEQbKt+APsOlRlLAcG0Q2ZWbPBUM6x/b9b70qXrt65vC
1VremdLyjHdevKBwDGhXs80b0Co0CJYr0t8wdy21L77oCKNtAXIoP9NemPIZuKIo
XjENQLNObYc4Gllqh0br0GY7Co+akTUZ9HqIhFACcU7iz+ide+pRywO9RFX2RR57
A7Dp193Jh0pHuJ5toSJZjRJ4IcqMDikiNRpOzAxOUBkmG0dU8WgG5EwzD9e6lpQy
fwqnk9yJkH8J97ui9PXtF11sUl5c3nkCf2zN9bGxwaaVmPjLPmaVxnNJ9BbyA1BB
hRGImVj0J/0kfrMMn1BFkDjNEELlZI2RPDaFVrwwB4UouyHGwI/lxa7N+5s12GTb
iuj/VtIJyQkc9ABmjPr+9DJRKpuRtjaH+KF/x6qqsXnjsaWA8xF1lSVt6XMUoh9q
PpjYy8i2caPwTo8otXV4bNDfUjSyddiJThB1iT4mfbjHm1KNG8YlMBQapfkYwnbq
Hb3CHnxKvP+a2rNLWLZoE7IGySj9F1KGXydmokLux9hWcktarydzjEsvO5lAfPdL
R/7Mxmp2/0FOP1htBSPbnkkRDU9dP0urYtUB6mwpi61RkGqn42tPImTWhcqYY68B
F/nWk2470ciyVxLt/tcrhELZZXoYUzvaohICPeLF3SDjqUrbkWJ2nUYa/92gKz7T
gbgfmLiA1vMI0lQ/WtLsiZ2E9EGP0TgIRmZiQBJlW9uMueRudYhnu1S+5mZLRyen
zWBtFK2NPE8+kmsJ1bGHKwjydRhv4nFMH37V4U1rEr4Bf+SrKKYnOigovBicd9iy
nkJk9u9d8l1XI7wDK0XNjGIJU/PVUqF5lCLGlJXyYHQmdcJeP5GR9eIn5zZUrRBH
Pe6Ywk+Z1tXmC3a4NVASgbsCILyimSFLtuUwqynI6si7K1tWswTDmedTg1fc8uTq
7s8r7/k612VKYOtWGZauS72sdRi3Pg2FriXmleLjaXbPtDH30quO5HRRPsXk82uq
a6auosqNfu848bPfv3Grv+7OggTz8RPmr5X0uEnodxEIQAlN8xaXopbeFlw+DHiS
QmU4uog0E8xUWyLkFvIRmBHi5a5P/+AmEzkv0OYvh76zjthFe34veboqrFs3SDu8
Q8jHB+fACfvGnLw9r6o+u1S+9A94aeyDqUq9Cwd9cnQrX3Hq49aSpDc8lx+cgUZC
6UzZQEAOXXRvabpvRdugL+4I6uaVmTGlLQfj0wthZ9AHuFig2MPLxK/K2moPTyTV
icTKlDZJOzEGwwARmkezBqvb8ewhMJwSabbxAGnbBh/Wu6uFa0Am/jUx/Qdbn3as
brzfRN5GCXrAfEq/55lV24Imy8t9v+LYhUjVL1Raah1LnbuaNMfOK5qnLZ3MsfW3
SceNxGZ01Hg/TItMCa8HotIRf7rfqB/cWq6Qv2neHcvGfi1tOqiHZl/1lFEhPAVU
7md1N0eFGckWuMCLkhsUtCHqY8a9be4xvPV1kHrMIZ3x1z2KSkPkhktBe5R3k0gw
es7RtOrpvd92Mxx0Uuxp0ttF0AblpIg9SEQZtehMjPqR31SUVAzJwlTHf+X7o2iV
LFAT1vF0EX8o2Z0MSQvcz4+as26DlDozP/LLrQCfGmDYFvOY/ENJDe6EffkEoVc0
9OEELdAsm4AwXGr2qZJFi0WGcxpQePh3wun5ghb2e/OdnySPtCi3n94QsuPt6yhY
CWE0TEXT9f6yUgeprSIRmbMNhEhF0ZKiao8euEX0cLlCxhuOOF7ngUz36bQPb1KF
IbriJfKw+O3j+MEZOs/WBJfgAIurzZNUXOj07KpLB15/8ulnazRPbZOBRtWDj60p
2h3705v51JCRf95IcuR1p9LjL04nqVLWdCfixz2Ipuya4gC18rODOoEMgtohaZ8v
uqOVaVOyRquxlug57XemtTK+6DYKvgOcTF1VPGEDXtN29mwlzNQnWIDFFH/+HaqY
ufDIlu9zdPMFnYtAOlutBan9pN/vN+GS/q9e/gVIU4zhcX8g5lokiZdBnehuGkaZ
cknh2XXU4e8/DYWtxsbNF9g9UZ02j+gMkSaqiIx4WXKruBqmbAo+T+eCD/gBE2j6
f5aupSdqIU9QSpT6yZsbQ8owlpvD7mtXihRr+R33YhKq7jqlmhyu/KaUHc4dVrFy
bZNZQ8VBYy2dF/Raw0jtSVqd6V5i+4h4uK3NxNbnV7Y+C0x0P4i5aGWUlA6qeXdT
wxY9nXDJTvToBIc43MWL3ZnHaMiDQggs8Cdq8CCfAli+eI9mYY12wqXQl8UUxFze
mBip70uPYf6OuXF+zY0/QWG66l5kDpDUOZT6O005g5Nq4Jaa6CneayXHJvoM2lSS
7VWquSni3zcFQSOHu1bk835S8OshXJp11qEvzXcje/WQZNx6KkCFsDhVIeUReJ/R
9ajScK8k8SjHgI5onylpP5y0FRD84Z+Amj5zcXN6zi+0YufRt1FVCjBpnXeCZ0wP
zLYx+PP89f3GJL5MHAwkShM/TZ9oS7d7YReViKmPttdP8Uvy2wtypEgBuOBMDNrx
n4+buN6v8Rt5GFc9re5C9oybEWd99goNMCsxhxGVGvawZiSVTjzcxGs/ehrk47Ee
amSCqWpqjS5S0SwYz0THQfwleQVzHDHNlfhr0RR7O53CVOLSAKtZTSqKN7u6fz32
YBS8NTitOnX2e4GZ6xZe5E6XPmtIusPk37lXkzpZ1md4khgt3feFsPNpjYwCZl4c
S54kok8ehLMxKnJURiWqkcYRK65houaEXqkiL/etLaCpslmLxjxfkqLoUPw+GcsF
1g0Gex5P3KLtWgcl/7sWdpjRtVOxmU/aeB4w5MeIA1JFQlnCIEB37I5c8uGh8A7s
aRVWW702eOnfzjdBbbx4AqWHQghuASnDWXfWFRGbQbJQiiz7jVJc3hXo7MtY0lNX
6X33qqaI1C7xJNdjY4q1YhGNGvgFcsHWGiWjOTAWfGGLdlLKlcVghDXLPZeKx/gp
y7R+QYyX8COKwIAIVJgfxvPFKq8+GhBgi/LNajbU2ANe+gMzOt1+dJB3C8ZQyBbe
XPSfzEfOjEB8ORCvtLuSOEvrbVypqOeewJqJHjPbB4EeA9O7Vinb+zqG7CzKYDEY
Z1y2fPHr6agLzRqMLRmSZtJCb784keXkc/iCRsgCcFCDcaVAcvTkcjjqCjlahMAO
swrGC2lett/QiC6quwCVYGEHRtS62uH5POvUrcjfZ3RrOQsEf1+Bm5AO5vmlWGf0
5M4242jsO6AL33+FusMWaVB9G9cox9IvSDyMF858PEx0RF6OVDNix4Vs6JTJtTdO
HOaHpK4c7B74dk/Gm9MRInmcW8TDSjiykjEwosrMFgnwzV+VFFlhWHzmnFQGSi+c
80slDStq1/tTexi9IH0yVnhpQWqpMKczME2T1icdQ4Pdt+wM0biIxebdwmGeELYh
jG/uxGSIQQLKTEUqaw3uBVTVfoLdEJd3+Ak2GlcrCpqs+LuMRwk+lrMaUR9nb3pi
Rf1vwPPS2QaDAr6wC09lgUN9QqgUuci7TLplFyqjmZvImLxlnKTjvjzJ8WYMVjGd
W8Npj9xpHyvJjzlH0GNVM4YXTKoZ/RzOHflbY7jEkhrhewsoSeqKt9clmKho30dE
4EWOorvxeRI5QypLKGDw/ery59wuaqcCDOEee9uMAgBKFp7WdST4+JaT2mnz34sw
kdGL9lzP4vUbcjst2e/PpsNSVAspWePMvKcKTwwFZJ0Zheiv6xGFEfvnSI+yBVlu
ucLmfoReA3jZPAPRkWM7QSpTupffJmZXXJafpckbORC9N+q9D0Hf/VpJ411T9ZP/
gtiEo3mMc1dYc8OQOSKjxt/VRPD+7HHbGAxVdvss3dv7kF4vIfzBtgb+mbyiFA67
xpELLeO+Lqmpsl6k1CuOSUAv6O4EBlv9r+X+1gJ1ar0zMhQBs7m2nEsiIsU8qTSb
kCp6L4zbbsaUzYaXj5VYU0F/FvjmS+lT9qZIP+2PVqhDD9uOXG8KIaLpqyZaEQ2W
QGAZzprK+Nec8F/6pCJyzxEbkdsjfVrKIvJ61QGIXMmol6kv7kWG+gcXFADxprJI
fc/etPC44RwamBPCkqlHZ3hvq8uTMpr8OVdJA7Yy/TPgm4JN4VnnFXjJJ2RiU1jf
fQrPdjpG6AtmlBQ2k2LQOeJwt9KQDaCLQkLOLUidD9uvuDZckSsSOZvztMvzPAeZ
mvXftNOgOWhTu0wU/ZyN5vB7JO5goDoeiPJsaCCqZWPLISBqkgMBQ0uV3BffTPVe
7ZVtENPfJM4lr/T4TbhCrVOvZ6Sfo7wzdp2EuT1BCW0QjyuQA7BhIm5+or1zutMf
zMKK2oN9tMePzy3FPjIHjsbDPurN6JmHyagxWTZnWOlIDhTNDt+ZTGB2uEidn+hy
HWi8QHZiES6VfIJmXhq5Ryxg70MXdXy4mG85b1mKvfBFLUNvHu+Vxh2LjsF5g2c8
Assc79AckU3qEs6xpz87IktlnSRT+R09AJugOZoroCQLa8Z/QueC0fgg+BDkeY/c
8o1I8awsBZdppxF4oZtqEYTQN/rzxypyknnEPDvXnC/8gaUq4//XHy6gGmGz6KAy
0zs+5KoUqjbIIU0sb6T0hG+aBSS6TDa2tZqF3ZPLnVXiVTFPFSlAGloWrdGG9tz3
Q+SC3INGlcY5Xa73gzaXtdAT7XOqZUKfibnusFhmdTSun2NBU6Q6hFx9wSIoamCZ
1x9yixnqrSmIZ7ZhfSEoYbvgESeuu5hbbdWlZcYEIcMTF7w7LPfst2QHXxgA8DBn
DVtPa/EMooxqCmmy5tVwwb80WLRCl9KsP8nCvZPFZ/xdNOtSJgM8eIJ5fT8Q6Le8
oRWphI/17x0GY4PARTzhYN112HNwp9dPB4u0V+IClHMOC3ncinOcCtS8n6dYygR7
Kb8Nk9OMPjPbNtyYq1wsVoDkspg4YV5wc5j3z9NuVvi1bqB7yrNzsFlbPNa9uRk8
9Z2VWYn0O0tiCnv+2YHgvLzCt+jfrKQRM36tDivPFuIK31/yZCTw/d+NWw+8bozh
LAtTK93dk8/tMzfp7tPvVBO79fDqmfEnExFhYcnkl7sqdIAJHRsgiKXtdMg9yG9R
VhVcNUgYmNvUe1JIrCyoaqm/8GaoVe453HLL7FWOUWhAbf6rf53jWrgbUpjH9m2C
xD52scvynHMWCXc6H6IVn6ccSQZ8j60QNUjGIeWnPP637yE3LRpxspaxSyrUrT+B
VYcvwQNcexn3ht5Oc+Tob91iKs0/Znq+qCssnqOpWpE8QfhBOjGO4ryHlFGO0uN0
BBQLVg19UpkzjlUjQhhc7B9k3xECqcStM6yQh0P8HQIGf57pP/aes+DLdo22MJ+g
l+5wWJ92+N8Yxpu1RLZs/XxBK8zIhuroOnLye2KvWFBMml1u1cHk4MOsTdqlyrwz
OzGn821MHSdyFSRbkUSTmvH5M0D2Iu2J+z2y68jq80SFbBsXqYpkjM73opvmUdrk
QqCyWcFkiWqneqtTnfbrgSkVrcWIXXAU+zmLkurho/OkY5DusnrC/fyRp50X61Qj
e4St0I0WpDUTuvi9kMGBEMKFp0bm2pljgbBc9GjCJ/CnSHKsiyt3LhxlObazJS5J
rgFN1UMxAPgda6culM8fCnaiB7UQP4ZAiCWKZo5Wea6EvocDKoSW48OYS23gH+Pv
PmW6zJh/eXt0RiDBhdK2aaWicASXjNixDRgNgUZDMizHGNiGDDkovIOrjzlf1M87
ZwK98/3CR3yZj3Dn00s3EL0ltNp3mhtO0Eurt6EvE6ZkNm3hIRgwVMZRQ/BHZ6EX
YEnVM0Q6jjWVpLfhgPhmXExc9x/W//VOip+Gmn/UevBjCgCq/+Bm98+auDIeGAIp
Uh4yGHet5G6fTG4bDCkvwcoJfMUKW4yJ+lSrlBrs62LBLiTK8r18smr6yeGIxioM
NTIfwP4/myHfhFMPswEEQPY4XtX+ZPb0sULer2HXcmxm8VexZhhphUxkd3kZExKf
X1jfCd2JBOvUooQVT6PZwQduAUdYyrBk3Wk2qOYpWeyNhtGiuzJxIMSAuklxSl4O
B7nnrbsMYpzcOLxHcNBlQ8IejSf+1ljx8LCGie/7BqoHnMqE9OxW6Wkkjb1YyYiV
1qDQA91msJRurjSQp/AynAR/3aWoXUJN4M72+tOFR3zpGH9xrJZPo106CfWhtqlm
pqRnh8uRNqbGBQjQsAkjqm2EIkuPnKQy/ApHNdSTWLH954FtWmUGwXsL2BHR0Gcn
iHmgQwPFAjVRxztjGBEJAA356hjBf8BGh4lMFNey8p+/H2CXvYH8JbZrDo04IAh7
1kXSmpEUviHGiksOQNABINV5bd/3SsMbJ30KKHC/+0HRKdwPUJZx4Yp65JvN4UGZ
aD0L6cb1KpHeDwn1pIyyt5xTh//2MJg/cD0C21uIHs7bjDdT497OdJpoPDLDwYmQ
GVXmEazWXdbvznUA8+AyyHA1zZXikw0Ev+/30WFtoyxFo08cfJb3hfh4PEVAw2RB
xAzGMtRCGojVq+yENUEkrmVnUEyfrpTGlFOnerIN8ywD1CMMaPtIZYSkKjShUvXE
kIFnWB/k2PNxA6xZ5GSRlrgwgjWS6rVGDfxrY30//rn+pJsHXfhKOSIlCZZ+8jyz
R6QbeFYKqnWLKQipBYSsJudu3MSGGADtR2X/+8WmBGScI/udoloGDtdhavNajdHF
/A7aetjWN3fh+KWKl5ftaIzJYyzd57oRDou0+m5dwH7DGW06pdmrCXNXk/4HhxFX
wdGHH4Bpnge4w12pSMMWaa8/1qlsLfmrGVheHpTvemXgiWbHcojqUvTYFYhUxQPt
Ztj8Bem5ioskjmo/5F7e0aVzI+ovonZ8reMnX15C5CBJYVmnnaimmMUrWgLrEte2
7oN8DQ0R4L3D7zoKfRbYZjfM5xzNnTA1VT2gmKrgxM26nfrggEXfDUjWiEYLjCnP
SMXxf38pMUP1OygIIhYbzyFRErDzVQWczTT1gE4wMkYZamVXy8qhxBx53Gwnnpb6
mb9wnWkTH649q4xVe2w48lv6HMmELiG57kqh5dDvDZgzEu7SNdEKRDTe/9lmjpSg
5nNKt7kCA5PHv5VTOOuFI5uIU3et/Hsm99BY3dPzYeJjvyThsAT/sMoi7DgR30Of
yC4qKpJDeP+CTwz4sKY0hwX++hEzbJW8BGix1Qsr2DE+5UO+7mDPY5LeOtfaKTTN
q5crb3AtWpXrd8WBDK8LWX2jBVVik3SxB142oJPsIGcoGbU3JXOQvcJbjrn9/tJv
qFWsTLZO1gTdTqDCYirWfMyCdxI0G/VA0YccTRjBmJ+DGrTJl8+527qBjiDP4rLr
iZ3cvPL6Gvq40XnVCLVx+ta2BvmAyOkwmVTw1I4pCwOrRU1FMp6oatwUjaqHR18u
ABQ7z7GV4e6Ksk0QJz84UeFYIYn+BEvI4yfGAxaYh7fEueaH96E9fa5O7nrtYJaF
6s7smbNEDzH6+aJgDpVOXtY7A0fNk8toaZwct5AygLB8INBXpVCOlDKhAcSLlB7k
n67sYs5tdStseO6wllsuCRveVra2R8CQNePlRnkCLWzeCcXXZvppotCEsKooCuzW
Nn1uHxXAj91Az01pQ+JFfnuUjPanjtFAvXvBiekK0qPkTrmQdrlcL7QofFplXsQP
JCYblyPQb0TVymVRCvf4UlGPt5QrTayispLK8BGXJ++XpNYc2ZSe+fXkf7tMznR4
VPdUFUQHozHfFLPEtW5y8EN7MqcK+TJO7DJZmHIPEFTbxVKsMa0n2zMaVVfenmP3
W6gSAfNUGa1l629r0cF6uCzPOP3C9aC5JsmseNDStwDwlPzZec/uhylLXT/Sgv7P
dZU+nU6voaEdiSImX9eHgbn10Xu/00J1z92ZWBgL9lNynl35QJ1LriqPTZ/J6xd2
0H6JR/YHXxBGaurk9/hRr59kJ/otaPSF/g09cytLEmUU/rxG1r8IFv7M+LqkHpIK
v200EPKJFGsji8Qke/mkqnFiLsLqXFCKEhCr9EHTd8C9Udbt0pf5bNfrC8SJ6Q5L
u50EGMGPDnkZ2MM19E8+HqvR/x0NdnCKb9WCodUxo3mvoWqxW0cl6uVqMZap2lPR
hkY1Ln2/c3/4022RX8sxL+chCkhvDOFr9mRsQmHJ0LkRKKT4q+xoon8XqeE71ICp
Hgg9HVAfcgiYWhYhs9jn/ZWSXak6u6Z/hxSRlUdf7Xt3VRXZD82kowAAlDY3s6iq
L7H43Q76Vyu+JUxhl80/Kha71ACEIO//EXm4bqFPpjhUaw9E+TMVV2ArwycE8Rnk
KLht+gLsM8DyLPNnbc/YoNoAQp5j1hU2ZqA8Hs+11AuavRFpWE9L/lCXIUaJWRCf
IYdkhUt/QdSyci3HBGSISw6ZqXH2p+eHJkSXB0zcBL7dgzJadjiM6nrhDx89dk/0
VESz0UJEgiCC9JkMst7NS9sWc9Jbd03J9qrnkwY+4pQp4ZVOYdKnOgFCnKFU0UE9
NJoy+6cd1XnVtELgzSyj9vxanfv/espiUveZmFwninchJiTmfgsvo8MS84j740K5
+xNonjiAYLCGwvuhkUB02nIvEq4tTagKqijUBr3jZu9qiPc3NScjWEDKZeJGlBze
fpMZlywV0KGP4+ulPlfxQA8FvS4amRxP4WwTz+3jW5ZQ+YXnDeofrON3JouX65vB
Pd55ou5iMKkGrS55szwOJytCcIu0c1ZD9MfuwzUNWVM5xed+fr03UbIE1l9f5ak4
eC0rlaXqynywO/XtyCILEV5vHOlsZHc3zqLEfn3b64GGiA7R6rs+EKY/uAxgJFLj
NK1jODqCWlcVLnKdH4VqzGpd/eYay2N29MeBvRF0yhHtSJG3aoinl5osRBeUQyWz
p0gL7wq/i/9tWZBkglx1b/wdW5LonqFSnCkKmOif53RoOp734PUB2DrPvePC0pEM
snMAEZwwXtyMKpvucAKskxgozs4oCpuOO5NTxkN9xXqoxxrNwr+ihcTsRv4bvKHu
3mivLFbm+hqo8o1nheIiIOGiq4Lxfk31B23DNKtVFsHyUiEXuLBvqsjlKXrsa15F
MwNLc+w6N5dZdRHrlj2oK45KfOIOKldeh12ZlDAfV/nwchkH6/UJN/k1/XAUZ/Cb
WbHKc7E0kOJbDN/Hp5fOO05yOxxQATVUnVH8Nk9L/8CvmjsxjPUvkZWHw9fg0qd7
qt1ghtqNA5ORUEeUTQ32MqESZVjQ1JpfrUwoJJDOt8q6Gn9OlxlOCCrc8oUWBGw9
yRbCZ1sfGDpQMib+LBYA3G5c+m0LiVcXyxOVW2v4mjIecw807Qs96VJDyKZurPYU
q6AijsD+6EiOrjeYxgEK/JPhivMEuPs2CoOv0FVnNbdbburwU4mrm38olLWdzW9A
bu/UE1Pe0VFvYQigTHd7B5w4disdrulMVFnt3FBhysz5+cmHp00v3gXahko+N3WK
8VMAio40yqRlPpocbCo7djEydIpVxzyTp5y32uu3j5MXH/+bG9+tIpoCNFmb/uNk
K3ppRCxFdVeWCFvdHvoWWwopwDBRtRg1IbeT+znqe+Nb/Xh0POXBaCUAGQtVqj4L
Kp4EdBbERgcNLJcRo4uPfs+jWBCU8UEx2eAnETuFpnm6eNLQdSj005DlBQzbMzs+
YJ9f+aRLX+N48pSaZn8Ns6GKIwg/liBjZzCYGqbbb5ozTaftOsXOa8iDpvLYbofX
9XtriM0LJw3KOTiB1EAOHtHjhXMadpNkHvUjgJJrozfCdca+UdnT40AFPhTOGXDU
eVUs2QKmemXG8s7hXmRkMs9ACLvjdCA3/xbFraxxYQ8CYMHnGoufpNl4+Sqy4Vgk
phei2dMP1x7o3N8JS5YB8ubtDvgI3qpFgvLzEOByCMevw7YqvDMjjwhRlZdGLT8S
IVVuYpDKL+joqX4VJ8oCWjnt3daXjguz5CkCVuL/EjyNso3se8lkAlrNdzOrTGeo
nBpo6JaNm3Y4tUGEHp7oP9hyVYLWyp9/v/4WQp7myVHjkQgf0FuZskEAaDEXijdc
0fyZCJopY+e/v7YZYFhnTSa7ZczLFnZRc7oHWRY0Hk2UlolYNXDFyUfIpnALkEDh
kFBn70zC8KcXqW3HQtGaEZEFll4LYQfVLqkvfsPCRVKJzZ5VcvPMMw+DlfFBc4Hp
d2/XqCw6Yoy27ET4prozWeARJFALlU8JLy36MTI7mNJhBAVSOsCrJVj8BefRrcnb
j9UbsqYPYuf9FnlopF+bCCt1RipXEBtfp1ASbEodYQ/5SRfnq7qncqtuu/5VY0ol
16dajiGjbOwAXR2uOf9dSJkhuRwd+FHzJ0LjAmjc2HMarMLon1q8iTNjcBd0HWEK
vpdmQlB1/JHbAwP6m/LTlkM4H+3Fdk6lDdnAvVLU2hYsjV8FM7Zu3DqFJc2T6L+p
uprSg/7jsomnqCB3zqzCV/YLmYWmuPsWGyMAsc5JVPt/FUu58tJa30Stpvd8Cl4o
XUAXg6CDoBBdoPQLDNTnk0+1o1B8hv+39mGmMxISLKNxDfEKq4gqIDuVNbkQ0y35
GkloU/t0OMtS1OatCa3Logz36g6i/D4VX3lQD0UBHQlGZHEga62WcBgvhmvoO+bo
fLad0rbUdBqgFsYI0RrYEzkItaF63WCQh4dV0RIr5RGZ7Rw1yMl1QeOs2K7VJbhN
c0MaeHt4j1bkpnhE6dRBvwvbXPi7iRvRZlQNCUfdSWgo1mrbHrC9bMIuVFpvVGud
lXNdEUGhNaDatgPzN6iOtEenMeDXQSzFvHxEtALUVR+31DPB4HsiSAUSwJQP+izw
l7jE9JObxps/u4fALf05nTvjpziF0zadCRk1nrZMoLcINguR1yJHvbO5dpWMO/8v
X47ntCqvQSYhMP3smCsB854jv8L43ozp1H+sFgVk5z5ktQJcYgg+OcbiLqPh3lWm
OhGVM7ykz8MdHghBpfz5qjGCoRwKoeVV1rHKMF54HwdHfNAf4VXc5CEoQ5++bjLJ
1+uZEGAYTGiiya1364rPgu3Kh2w/VvnbmWafJZTSN22DQXwl6wudX96Y6jlZgg/R
4n3w8xhCkjJiCNg8EcNCv3TI066Jyb6eiRWQiXT1mSVsEP2lqPBvl4X5G2DYVNOh
slw7EQQma/IJeCASq1RlYbzRcxZmbTCnlkqOgB/opuLnSw3q+nA/URQzymJr8Mwo
AsHWQcpu3FpsqzxsqP7eHp1QbN1Bg7gLKUNsMWd7bQgNczlADWNaenhRu2nfABda
nApzK2RHR1ZYBUDJVNc0I2/FEN+b4uL8qystiGrLkZixDzlBjHQv7O6JuQfVyFoc
i5CGrMRBacY0kWhviCsQMzg4pwmQL1PSFuwPCM542Ph74P5Ai9ikI2THmELsgtkc
rbhTpidoOUmIKcrvi4lCPgroLQHefg2VkGwy0Kvn6XP3jd/CPDEgpIAowRoV/JK1
5qfDL2+VFePq9T2O0wc6cZN1PiupHhircG6OHNMDViSS3w4rqW5fR3KvvWx8MXDB
JGMt4fkiP2MM+7nwTk9lloZ3sBsbBgvP1Pnd9PUo4t/SHfGsmXrN389MHe97tmBQ
ISd1rKvNe2C0rgVc7dycCW7ntwnU2yLrns75AbSBST8Zbld2uef+dfOoppxXIScv
rMKhYp/zwyyOZdG5pzIKFKpD76A6/F8ZRIlR1vnxVwvBhkm8IsDGUV19gUR6Xbye
gymS3PDXuEVjIembKwi3UjhDRZLuAdooc9fiihtnlWFTQvud8Xir7J9pO5vCHa9Z
WdP+l+YXP2Mjs4oy2NW2TT9EdYRS2i1Az9YD3cfDLErsSOho8gycLTqD92kbY98j
z/DGPGM07yfJsRpqjA7YTrJ2UF/l2H55wIKQC+BMQQKBaYap/OxSBlqm0fmi9dGV
yg/fWGD7Pt91q3KY25F83xF63lmhvOY4Ij+lkkuYiNfTtTPmTaOapXV8LEQcohPB
VNU5yF3GTpSz6OnjZUMzOxuYqmWorWwhS7PWrgaEolZ/Vl/e36xYgOHQUkroeONW
4e+KW1ooxVndXmBKpzgXhObc5u0068GRozKvTxQrOqtulDSWDksj5CagRQl4nxKp
aOXsddYzQH3ysg3z7JtanLxBMO2DN+Y/PNsZ0G+BeP+FdcorG413J6d2rhho0zW1
hIfwQ8kHTaOnuAhwMdt56Kb7+UotLkuYpDtXadu29/6LtC9xqz6+WzinbNTKMF2U
L9kbtiFPPMjwlO4h3pEGS0V8AW97HJyhqAYz1/PiZ9ivzG5hTGaMxjgKNKXjs4cp
8irXl45d7mEZ0UCNfA6zsBVjPd9UNMxzWGqI6f9euZDLTXtbOD8to2GvPdpL/ci5
wsGP91u54CeI1gOVc1E6UeqSM24ZN8tiLb8a1hnsr0AbIVYeH3i3cOfRnm78LVHA
2qixb+pyZYuN0337WiagdzFKrNRVN0E4HC+xrEcfYJ3Cj2G6jCtyO+9Kv2KkkXBJ
feOcu1nMWTS3jpFjeRukFdkVzMmBzhV0AAAe7pEAkOhk5BE5fgpNzI+y6uM/3Kyn
Ihmi9QkeMtgwW1SA4N0Z4LfKJfjzYNo1OCGXlV7/KM2HZlyZHRwIY3f5fBdZ9RJr
pohCRCe0Y3qCDi5iZp0Im67trl4R1swLLl/6sLNWds/qkpEH8lf3HwwcgewnJXaj
wfrV7EnhvXVueF5W0KEclvlPRFEbD6bk1f34h8p9nh5jMX56oJlPld1D+BAvxP/x
Fcl/Zw19gFNv66XuwUi7xGMtEqbTZwirZxXzksxB767vQS4ekzfajkyfj9ltUPr4
TtZG6j73xHSlPeQHRci6w/30wwzAkqA1J/eZsS1BtFQoNBHtfuLYzbx4YnLkdDlY
qCw/H243oCOdHXRCgwhF8cUIIKTgC01tuU8OtpLktF+Ibgw3mOpFSIClNwlm0+ED
hYw48dvuaPeo3cKGEMYEjP2l4mT5DRGAqH72ErsERvGeO3rpwhyC3E3uTr9hPBJc
j0aFJaR3XMduYuv/LmxCKz+mTO6FaIvMEh8eZiwyhRl0mfAbqXDD+PZHnKdHURED
gstS9pI+80DHzVHyg+YpMrlOf0GuWe0qwVpDznkv0jALt3q5iMRDENmFzkV5ggRK
1bgZDyufmsLapEYkHaYEVDSQyiiMJfChtUBHncgwnz41hzmT5ehCV6IFJDo9h4Wh
6YAQNsz2zgV7q8DK9GpB6u+UL72mDKp88YKeo5Xo+JZlf/0AE6SOqCplyqx99qye
n9ZFgKfXvOcpl3qJW0TVCN9p0G1VDcnIdu8hng88rDVROvSqDxoS0dRqAWTbc8lh
TG/6HO0GoR6B6QWbMKS0CoDlqQlMyTU1BvfH6jp5cbEhmv2i/jWAQQf40PZyRcXR
v1BLSuAEqDOtbrg/+cKXEZMdKwC72zyhubW/c5fokW//fJFDwyfb5xd8LkK8XN5n
apPLQihBqWDSGNxW1vYCM7nuep3arEdzQEW40ABAEmh73qLoZlX5CzK/Zo1cq2Vu
cUodheu1WDsms08/UNKIuqTEuLyOoGuQPj4NcYPPsoLKAzzMiu412qmGrvxoo4Qf
zOItubE8mUgE3S3GjjvFZ8HRlxDG1f+CHPZb07d+EtpC8cQRH0GyXJ6wLlrgBDv2
rBKW4XWvGLMQj40mhWb69CZE+0oI0TjlehjCk0RK2kcasH02tX4WFUlwNbw+HUCt
o+XsY3IlA470A7p/cDnjPDuoipWafr5LW/cPAeVB4bnqfnloD+sbiLTtuyMpzplE
N3x/MXc7o0syqL54ePqyCgoeyWpnXoaF1cMNJUon14hBDmAkKcbn7PrtjReMzoU6
wLGvx3YcXplRAQ+LPFrbMp00PF/acrRqGELugALUn9XfjNYi1Zsv66dA3yZ5/pLH
mmV2j5h/3tpwoHWfCl+h5uAmeJftOkBTKhnhtaDqqNXWB/+86nal5Nyr+Zm4+uta
RrO02AEMzGuJafBBk0RSAXsRhRQCzury9q145xYc8lMnUlmQboLdOmpYVeleKkIE
FI/QYzmgZBTzZyKm4WW/wcxW9nKPeCzvWDZYHFQWz/+/PnTPss4RnBBelkWbbuSk
b9mAJzC5EMEqExnhTJ1y5W8V/kc7Kh4scj0rJzcGIovLoCH+5x4fLlBYd4rhQ6W4
6bCDMGPiDj6maFqsSlMwXTisDozmX6wAR4ChlxOi1W0L+daxCtMrfvQA7CvJowUm
TN11qAMW2uXgXzUgQ6+P0WF7DTk1C7Hl7Mu64ufj7SuuVUKHyQs2+GqdeqnBLSkg
kdWp5XLg0JwsnhwVS1UDc9XjzJR8939W96IJadQG2LnXHs2mf+L774GRPEp4VoLW
xUFaZntJAJM5PA39PLxgSSHAuzizYDVorPICY2aLvReSAPPV2aj9x1IHhexScBp7
WPi2V4xdrOYemjO+Qr/+WQSkJMmLuvWOMJ85wcu7cwtuXGFVa07KXd+MvPk2wX5w
YOT6lqKnfoq14PBQrBsxI2ktgw/X58yvP+LUL2mCuWpew5nTggCYEPNrgJ1wO+0q
s3HYBdAL9RvAQ1uxfTS+ER8deRuhoqvuS5AcoYzP3i5/sebfXSLXBdm8XzEPGX2o
A8/u+gOIK5+mT6fSk4SHyK0Vu365K0y01flD9tXTaKwjqD0dPgnpYewXt4tDtyug
/cNbeCct82JDGdzjeGNX1eJluOjyOMZWD53AjF9l4dxZN46FzyjE349N23vCCL3w
KnDLL9NxRGZpYPdYn255mgPWRMXvDhf5C9Ofh6zfiWbIO/vR/e6Z07kRpUcLgrEO
aBaC3dQikEX+fGofOKfAWSYpeuGC9DqNv4z+TJ0M/jROJxr8jNFpMVVcsjN/dqJc
PfQIrjUgqMHJuNnI/YhyoBDMr0kkaRhNHqf2LQp/SrvjlMKff9Ak5SfkpksmZ9en
CsVlMZcGykPfdOS1IcRR9NYfLQK72ur8dPQJikXsck2nOIG9Wj8VduL9uvXtEvdi
KgQwTipgAsen7PuCLEV+xXZf4m1VJ1dYeO2eYXwPfs3OV2ue8WC1o3uTvcgAVdgW
AMksZ7HO2GIhzV2kSzuf0pszb2nznCuq6WeV6lkSi1ic4g0bvkALKcUEcNqstQfM
mHECEHs74+u3qZCokKlUNPcjQqVr6NRSHM22DI0MfHl+Qm8OBxgxT8WpBbMW0hy6
0hSs41+OUZ4Uzv69md1WgF3pu5XjG06Gk1a/dysDnPRch5Mp6omPYoNEyftcrJGE
ZOOx8DJ2ahaea1bQL4a2weQYuLHZPRJmzt+zZ+v7OjA2w5T3RVusT3YcioCd19EU
dTNXDJJeTbbTDjDf++gDlEhUYxBYn0AcYoG3QqnrLDnXtGdz/ZF5EQQUh6ckU3KA
NrUNln/4j8nwAIn0Qq20I7DKLmBDH5M9f1idTcygGsVEGrHYJ9I5dW1oVYDHCpa5
KKbmUcv71BSdQYDe7EUBRCn1XXH9BKiczMAVfvUdUnEGA0ON7oAoHicgCW5vtnGP
2k5WtjndkHT6EM4IuuOcfDQ9R7x5uL/pxSS0xzrHJNSeoHEmEtCApGDerxtF4xJw
UrlU98QOU0chfp16HtNNtMKQWqEbZHhhm+2uaqHu8RbmvYKvr9+diSrdBKCat7bZ
zp2ZC4QxDyOJ+Yw18SXA/8H7KmH7X1nnhqdfKgItreTiIcHkf9dfvCMRjhTVTBQH
t4dazFVIkwhFgiADu0CmohVeNu4FDrvzoqcc1OCT4oChrlF+rMbSMZJT+PC+yunx
SNLaI1skTV+0cEzGge+J91cfAeUFs2SAwQlqwBOI7dq62hq3n/t81UGfOfWwJUGS
BS0SuqIo/F4oNyUvSfBjteHiVc8QvQkT/MnkuxoB+AaTb1XDAqjGnvShgASmI3jD
s1RcC4hBLzajvQ+egWctfYLPjDD3ZCCOEPLftiB8lRNO21N05ES6z40E8Co/PN+O
Ndb0kTqh1cUUa4o+GWG+JYEafXk+hxGrIqp9BppG9vMRrBNrnZAZV9i9BUhosP8d
/TCXA+gxuAXlk6LAvW4CsV+8fhQLcQlO4NyLHEHrhgunL0nxCYCCoCV5u3m5efIc
V6Xf6Tsgra/0DNdACSrzwq+EAzfXGU+M4oKLZQB7hzW/j4XtQGh7a5FfoS/Ptu8A
i6YFUDG9NA6WrsAHzerFr2fqu2iDZBv49FgXQqvuR2jRsOZ5XZsk/IH+zsTR12dU
f8qm7S/Hiext87RtxiYZ7UoXwXYYUhY9SBGNyku/Y28xF+WFfMeYim2xGgjnmWir
zc6rEXAWRDTe1cbHr0TV0GqrhLlnWS19M5VGQF4/I8MVwv1cPHcOFRHDsQS0SDge
AiqcBkt273pDotesLGKGMv8rC2H5lyCZrb5HMamjDGowJ74Y+E/qQk7pStzaUEbh
Cu6++XbiPGj9fFqi9fisgU4TYFfhKTlNjQ9kAj6SX2d4wVEUzPCi0gIcEe7fU0m7
2VXam4fpqhVBWlhHrepkMomytWowFDDZo7p6KnUmLhSPEpatZGe7GJ+DJE0hnWTd
eHSrHwD7DQHTGqhzaF5AYmgGHR7ux+RNByGDKEgpoI1uHvYJLe0+bJcRHq4FXy9S
zhi8Zal04oW9Jqz1vJsf9yQBhviu0sZT768kK6zaA5jMYRIvWj2+NWAFcJJqlrFV
2cZeq71TN63xK7xxx31Q5u8d3yJrTeWsFnw5DQH7fR6hIic76MRHCq8qZWEB0gzF
DgGfovNAGyBPEFZYyBzXR8ilWahLReb4lmIqxBWL+jjEpoVIZn+g6/pPB/Gg0jVA
70MFanuHY/qstWmkrMNNAUFuJ0iyBKPX1rprQK3do3D7ODwIrmDqVszZRZKrx6ES
sREVBSk0ribrU+EyRMC95DX9DF8PNeGNjYL3c4zYtti6aKxyEq4dSV7YxhRREBeJ
KXY8PdUXgRnjPzqUyUVHafuUnngXwTbpi2dakyIdOolkdfdgU3ZCCVz2wam3MUeD
lOXlwbmtp0IDMB1HXMENAa8WNRrcIs7gSBm8iFXoZRet8Y2K9M0ybyqTok4z2tbQ
hcOM3SYyNM2AQ+QKACuw04RfNFwDEFN8rYafFQ+IXMdyj7yb/8n6olIoLQZs6Qeq
EgEy9Tof0DnUStFcf/Kf+yrqUv11adV03BLKQML/GqEr9V6RoFF30NWQTM0LLDlM
iX2LjD/gX3huACy4JasazaDARdLFDfUhft9l+egeuDbdpLMAfbVyaUy1zqD+AXF+
ay0tgl0Op9sEMFGWJOK2CveDXJd+gkG7AFUd+KJIt3MYG95LOS98MpwUR18s4IvW
PLJP9X6DhwCHXD4/i24n4RUcThvMSKAEo5qdRB6VxqPK4FPrj+SO0YMWUGjAYyHJ
x6NoAjB1zI6IP6gx7yoUs7QU6vx+EqQBu3PjQWJKnnBdApg5MgWoI3Y9hJ49CThU
chh+2q9tg27N18vnTu9XApnhvdoqwCUEtMOLTvz5SVGcMPCbhAnWpolyyHy3lfXg
A/76qNbYe1up2hph2Cp6Tp02xKiKkl5R/MhLDbgdM4GnP6I8Kl2wFAuO8wezxJHD
Dkx1tc8WKPg/NSq4l2ipDbMERh/+WkHcOwky7npIbI4Q5Vi7s6MhrjSTlkxnijLM
spAgumzrgC21PTR7QWOZsbx53G6UvWMWSG4GR091z+p+c4pohKRwiwm8qaNOBVHd
aTh+QKG62QXnHoHCMgDYdM29iScVldn7elQQEB2aFck0s+DISIxRBhzAqRUG6s96
KnHEhxMFXS305KcjBxGV1S7MPDvlb0oMWjA1lnnLp0OAm6WZ1/TT1rKcWWfwAOhG
hyQ9ONp8U+4+dleQL1jz4vhFhZmepp/TOhBd0GgEORN1EyKDfJN383dxMtUloBsf
xm4TXnBNY9MMpTbJ1pDTc6O6ECBN4GjbgojFl6tTR9utYcL+sM4DicjFxuN4opO0
6meSE4BGRJJgqfFTRPcBAjNCTdYWFFNzqROh8GhR+G2PT8jWk2B4DNBMg7pHbkLP
1lmWFygf6O+4AyxEWicmmYZ1l8U+L5f/ZjFvZml9PgdSsHqs5mRyB2AMqVU7oju4
zCOJanzIplOl+ONl+xItZ1eJ+a7gmIe6Q7FzM+VGzWLhWQMImNvWZkolYKeDLjgm
fhtHjtYh/F18KPP27GxU3bpk8GHDmLxDA0Fj9+xKSgNlhdPCMK8nOuEvG8ZYpwgL
qD0p8ARgvLFHs6NEZwtG/UNawVSS1pRHxTy6Clo5LQmvDxfq/JHJRf6qAjb4JuK9
IOj/YgJShmUtBYFnQIJl9wmVgKJlvUPYhR0VMTHCW78rnzd9WbOqGee17WA+dCeh
8vbl8ge3RXtJjpxJhAsAw20qkwEwxQAlCUsoVo7aL6JrQCZfZqL4bALSaPRopKw/
OYxjPWE0hpeMnJStt9sgkTI1KzKgVtBtIWrnp6dtu1oq2RgR7SWuEQi9rqJNsTEq
4XX49PSwTZ+BERxmLFWFujKodxURiR/hk6gzCRxnZGG6cH1F9qBlaONYM3d6g5UW
CmdNMSaFy03zLB8ml87+1nMkUyxwjcovXoBhkaNYD0muqybk6uvjBsEPZUXb9U2X
aUcIgDIDMVqLZIauu+Ze86utoDQGfTPB89BckfMIUpYUCGw3yeonv0HYYgj4bytH
zrhZtASv1Rrz0Bxi5zagYWA3KNpimuoaNlM+MEw7kvowEawRg7MXjKG365CGLFCL
Bhd7Nt8ZvadqI2/flfhDHj/CrbKm9WUHc/CRim1vUhHmsFNMr7kxtwX7kSDgTy2X
dY/uJvkosywmieudJVzur8pFKooIHLziVFNqM5fXgEmUA2ARo05eSLDlP3CbgUYW
TDC2D+Svj0O/HhgxOJNyK+0mlofayeaaHGZELev0NBIE5yW+euVbGpv/BbLEzer6
6Ss8KYiQeubCp0EITIbMCDSiWHMVOWIM1JsxLGEx8TeY7kIOBo5z0cMBoZ4LW5k3
q8/eE5hIqMZchqsq6bh76hP0z0Gt/fd1SrakxqqEyDzrO/2p0frQ4rzLA8c2Ti8G
2nRznO9KqiPKYhqws3ZTdOPQcLZDKh88dPXKz90tZQg91vxU+warko+NIZEZONCI
tKgjhkFicmqtIg4VOJ4nWVfs+gkBY5at3ye2HuNUOPVG5qI7rMtkgaeLg4QFjGPX
L1GEA9TTotufMaa/crvL6zMYriCdek0sqCnrpA4ETZBZdFt/Jjij2YKx+70KSm6M
JUNAM+32rtmOszsd8yhBqjdFdkAdwuha9m48GnKpC/nuJQqZubs5hieAemDLwqz6
Eq9lIwcPxd38pQYfUOefUyPHHKxCemKZlAbzBhIgjRfsamOxbwp8gl848/H/oxVN
b50fQscudRNE3+AHN1AB8PVLZEzdkzAdDk8aGMfO4k81i5u1n0+WGmYlCsYu2bKt
RQi6JRY7BaAvlbi/hRuWgqSKb8TOsFxDLHz8lWWIs2gq6AbgJ6CbQ0EW9owOIHmY
qRt9WlBr3pKNZMHOWfxkCnSS3Qnds0nf8W/t3I70Nhz0qhhUKEXgWfxW7urkbp4R
x+YhUm9+Cu1jQySPbiMUPVc/wmuEYs4eGaN0gujkAcqgCa+4kvd59a3cFA1OMA7i
Qh4Hj0SpQkz0w8pCUzC+lJyrdqXXrzQUoulmKHrav2SzA47m7whQtWZCAaDR6L09
7luSxufmzsjr4naAHtrVWi3TTMsl5lHQ55kOrnVo0jArXYGPm3/XRkxTnG2VKqB3
bUzJiC6Q33IGh9LH3/L8lP4s9alxa4MfXCvGHzLeSLhMxhyfOYLjeJM6apycKv+a
Imv7q3WyI4eQCFFhgdIwThOOvKgGrUc+M51Mro+HdEt9S0fHx4R0JX4pyrnxDvt0
8tiFvO3QCcDEJtEOcRm8tv7vOUiiM0MvX7RpcGKi+HLCjGq74xM3vLx225qpYcgi
+MuzH9DNHVA/VSNIP9J+ViUhSsNGea9eKDNOEafnKfrXz1EMJBkFYpigA9KnoJ+N
1e4AyPecvKJh/L/rmhke9j5gXEr2sE5K4R3dQp1xstP36KmB4NfgcDGC/4IOSkfZ
Sy8Z3BylDy+cG4JEiSgw0YP8el6dmetBRD4v5udpceKd9Dg38zT3hQ0txP15aJfS
mo2Y9QCrFCoBexTRbOsL07XR0E9//h58EcqdiQDZSRxtS5Y6Cm+73E1qbe/qtuSI
/xe0bTQXlfP+9USlc1urSwHhD2rrwfEWQgU9IQ5jj1yon5QH4sv+B7VyVb5G44xc
YKml6sSh6kl+L/+OEuBCYLfVQiaav9qZtOE/Z51+d43V1bQAtRKVS8zpgp5gpBTQ
LfsGpwnMyDjnMoCStnCrplEWEodmIdkb8k0dx6arpKSnIu/ZldDEnFS055Pq88VB
8PrcKBeKqgTJhoIqABridYXKonYDyGni0bvTv+1LKnnEAXwbDe0RxgsP7JKcri2o
eUQ05Pj8fZl75+wUbjcx1xYSmpgSO71k3QaAiC5zmxPC4c5dY2WurzCVwfjpOnyo
xXEp3F9SzmEb3HfTvSS9NoNk+Fy0nDRDdVKMc331oGLvRt95PMSa2EPOcmpegvz+
hPZCmS/B7gnMbxNi8xWPjc6QEplwseXF0Kj/GoSM/k1rgp36KF5xEfcbkm0r6Zoy
0+/PMmY5TSEHlwB4Lbf6A2fdJrXNqabJEdtc6t0O8Ge1KsRDlfBGijXIl3pMBj9P
6MdU4qk1ec9hldVMiXFxfR02PbZVmlMvLmzb8vvM4FEjVnBL0SujEgQL1TOzYCbO
JkbBtY2MJH9+wTK5hD1ySJS5nrNaeQIYBFndPZhRYIKrFnEUD4u6mM/GfZbJ+LLz
AzPju3dqaXobmZiW/WdM5EaR9LeG6wf/hQS5JJa//qPoREhQ9Oo+NmA+R+w5IkgK
VCRZvLdmKVuCbEQYXtPGOgpVUyt0WiyHgT4FATmHNRvF7rb7j7FFh2cIOaMyfVO1
w1mSN2QFnHvkeLS7uZLMNUdOe4dJ21pwRzeUL/UrmJ2uMEFFf3M5wY1EjuerrhPI
FucchRLrSEPKxaQAQ0K+7uQYuViBKgxqLcIfjHGvXJTd+qs6rWz8s3BnjeiVMoCO
+f7NT82HxsiW3CL6STVSoU0Xxfr4Hbr9amiv1mhBaFwZr23loTQUbuCt7OXuyswY
Rk8IFQq1xzsX4rK+KUky8ndBfi/Rba5NgNPnJaZ4Y76YxA3/Oyfh1J2e6Sw5Q8Bp
jyqtE+vjBsosstnGtQ8zEfFrwf11/Wy3IPXVIxj6KGAVSs/cWKAcqr5ACWeg2ccL
WQGUtZ1Rto/5gLHPIIM/KOZbU/A6REesBi0H0w3REFYSrfHA44X5Q67IrLQ02pwl
nzlsFbE/rn/UkUEM4Mve1uUi9DsH6tBSxSgtChFO1/bKLIFbcYSA+na8Fmh0pG7m
avPJi6gI9FZujx4bOUgSyNZNvnrmeKdaLHgnWPm4aSS4lKvNNZDyP7eGcnIvk77G
A+4HzLDI1C74grRTKOxsop9bdrZlTPM1vUoZIJ1pwMXf4kC8xTF4iOZwpG2SUn3F
XOblD/Vh3qsO8txS1MFUsqBCfVCHqeKmDnyExF8epHIaGyHGEEGIZC7ZAjriQvOx
4XqNoNVQJou1YGmc23HTC4Nfd/WJDvAx7hMeQ3KvV0wUd3qWKEn3+pkpIFs5pZpN
iwp5zLXlrv5h3WOY9V06UU74rUv2IvZnSeIH7FgdQIDUyvB1CWC1b4pxZJ9M9Jl/
YbZWjSKITo1O+NpzbzgiXcl4N/kzKbIb0DfY++wDO4bMR9mDLiYxmBBFW39HESF9
jPPTmzry0olK8Ba4+j5aJsPVJAiz6TzbLyj2IaQ8AifU0zQ1e4uFs2LTv6KnPp/r
C3oc+1J29L2a4fuNgSlC9OsegSBSv0KS6RtR/xd0CVkA2fBEMLuUXrx3T92vuZlw
vnpW75hlW+hbJ/6AevwMX+SZRQvHMDmGZGKqZfBJ/ujPWyMjyLjCbfIdEByqa15u
wv4HY0AnSATabh5PBjulNueiNRhxVheyRqpqWj8kfcM/7acnINrfgeCdQqNteatw
/2XzRjGaSrAzef3qCFK/z7khJv4t5/nxU21bSVphUa6YiMEmI3iWBZ+q96zzRXBs
z+baahaNzX1TCr0GQwSCJbg7t2ORi64jq41b4Us0yey0JkBIin3Qq++unGAkCz28
RNPC6omYeYUPVNN9+lJuRFK0eBvSGEj6e5PsAUM6Q2Uh/n6y1YLbJPuST7JDv9BS
Nt8vmj+cS0DfMHFBHOyQJMBBoN4EA5eDNVf1rAg0ovq9IkbDVEAcAhd19J9jj7kN
qudaVMWNAghWd95GQ6G4Ebnj1kc/uGvqwm6y+qpbd9y62J3q7118iR8gnwXJkLPJ
QWpa6GroBj1RIQYhj5S8mrdUBrfmrLwrN6t4aNJEAIYeh1XESCMmwNnP3Hko8/UK
ySslv1GYO5H4C98lag94i9pfTpGjg7eqmeKMH5q0sVcgF7Hg9pLqAtbchUp1yyPg
Bl6UhktdLNzIZeMvSgsMZT5aZHMBvwvJID518KhG7WOKd8lIGEiR6Npg+KQOpnDT
jEV5K9hUafNlkLTf2yaN+yeLk0D6IyDAoRaGlKXBOMr3++Sk+bUPiI8uy/rJrD3+
zEmc90QCAq+xKjqLlJ1C/iwJbYDObTENCYTG/wAPEyqWaTvG2a2kZfBCqv26U5hp
gh+cU5Je7TeOWYHIAVUlEcWceTO9F6KTMZ4tgztnMlonnxzaeDSrDRAiLcxmfyws
FPsenHzyd4IPLMNK/yHxfOPjP0UZFTw37Xr+vZEhYssxtVO+SMxV6x4ezadlpAxM
BlUxTj/5Qj+tC0XS6XgdQ72NPqkKsfVNlXsJk6vzpg0l3OZ++QnuG1pXlpZSBzns
lVraOLgnkEMXWwTukdJZ7vqNUm6vCF964djzK/IaZcRGkLLAFEtVHYaIFP5AWLQi
EwWcqHi6dZsbMGgzGK7gsfTsG2k4P5WaCxx0TTzMlg1Uxn81cEVvjyKXFWSXQziV
xZ56phLgqUgqeBcp8CxbnLLm5mP6Rx6ylV4qXn1JAa8IxOIHrf43UU3jxeR5t+GD
nDm4eTRdU8EicW5OyAdt3aFO+hPcvbYSDL99z9L+hBQhyKaFwT61A/JTLRTQKhrd
J0PjFmQmAc3ieFkx1AuHtzs2dUDNMToDQ3qOoSUbnDtIcQulsra65tb2Yj+b4jjh
HlDdcp3vQEtpbuucexvfb6Jid1g3+kcTRatvkdjRbjgGKcU3ZXDxh+bw/TUCs6Bx
devylLSwYvDBC69xM2hwpuvPb5YATpbtra6cp1wvxM82ujI8xFpCI1P4rkgSTQbm
DBN1DaF+3IIXxyqK14PO0AfYnvbYTBdx3NG577QYKfRAciA/g1UhF5a7D4fvmuMD
jNFkWycKfknhEWyTHp2RKXCwJlOVqhRRATAfbCHmkliIdJzZuPD+ge266ngOQBGH
ONuvkHwNb5CQZwWMmOkeLfNNeuU0nm7WCHuyymMSS+GWqhYwAnE+Il97cmuvbgvK
gbon31tCWmupw77tNggtwcZX3Hq/h3mgsXYuegqxjlPvvJfskw99NJmtPDX0HPLT
RjLWzK/uLCu9WySpidZrAhgoivfvKeHuscKyJ4FBgRpNwmYnnn7drt9l5b41nbZ4
XxZ2Yy9ADZb1ZjTFxMvop9zpkKzxLE9QM9BZLwUiH7kEZxF34gzCqJzh8R2i2MNl
I3tMduOUn+YVvcg0LFpIUhslQQDfZ2vhdwngX040zB0tRrLtp9E7EDAAF4MYUy/c
+339dmjXaFfjpawxxNCpp369sssP58zVWCmwAxeDGTTlEX2Mh+PU/YnJKOle4ATm
eQgnkht0fPlO113hGp5ZHD5wyyCAqXK/V1dNAjfzDmsKKquN9YtIB2Lmm1A8uUDR
WGOq9OqhydKTAeHpukhU4hx6mjkYzPrxmhzRmRRQKGZyvHfRZVXw2t5mB0lRBVuU
S1EI6zIelc3KlXApvRf/yqsklwJESilo5acOFw2KHoArC7BKBCcv7TXXWKHqZN29
S3m+4NeUKGcdYVgkub8LaZgkSnMiuG6G5WhxyHG5OWJyFS0xcVqEQObcB0KHrAmd
QxuUI65nhsnt3X1rVzXEygPAdZaqvMEyX3925DQg5TvDECRYgW5ptrxTuRDEfo0+
NY9uCZJEDmLPB0q3uN5mNDlIl2vcY0A5bznrYT3DGDqwuvlfDE7wEZ1GEZII5r0b
/kIAG67xyREzslIMqqTTXTB7lWsZd/lEal3TqSFONwIrVE7Ueh+6nYcXBC/+G6ME
/PLNZpb62SIjlfmMjP4SxBnsBtKf6v14tNK7MypaspOMZz3nKSjcbcKq1H4j3RA0
Mir/ybuXh5EGs9Zk//6h9ygq0vJvegOfSpK5A+t7W6/YTMsjw0y1IvORVlusnaNH
ruODIuWpVHZj65rdosKSsZ7VGvfBjHuMrKR5xbmlCXKA6zGSaO5kwrck4vaIk7uf
+X5GV1t89IQ8gKxT+kCIs0NrxBIPnDAr0iX2ngKbCwV2stGHvrbTihPJDe+5/Ecj
1E/7DZHCBme5YT7ktPdWVfXoPePJq28pMoRAmA2jOuuMJojWtw/zDEREBid/ASTz
LxJYb242JuoQFyxVCWfI9kIUbq6Rf05ty6qXXZb+fZlW7+Ar502HPd9WUD+q7dUg
z3o79ZVh58krPZhyLim9jvgCBDZbV5vXHBCNeW82iwIrkCMswxcuVEDFtLpV9S+m
2uXaT/NIe1+Ajxs7m4CjYWj22t5oPi7eEI4Y8+Ing1KL1rF0J4bSO1WNRAM2rK1N
IFlFPkzhnd7rj2FLs3inJMcFpJ1yE9acsF9bbDMy8lfrCXziPlwp5VnP3eUaA/Kw
QLxnm2p0Ent/hEIc3A8iygli8VHv4g4Zyi21LmiNE1pxtplKrTQVpLXoUZL4H91n
USUAP4g5cBM+BnIFvlC2ab5EdL647QjekC61RXFbPiLe0As57CEmJojLGjG8bhQi
c1vPWSW32tskbtusRroOByWIYO/DPPd9vX66LJaWZn7egoZQHPYbASGLLD+mG6JE
V2E3FCURyF7srrSTwkva00545IHDVdiqHZmk1Cd6+dhsnKCIhIjsikRPGKqsl+MH
tJydpsggF94UgDK86vPgk144wJmwByPiAvvQfPq+9gsYWyDidG+5BnNGwMNA7oUv
xfHYBrLHZ/Ph/cuw+EUXRpi4U/KRKsp8aXLsqHD3jEW/kJJHPsRlTlbbLjKOm3s5
9iwUGVIS4B0mAjtkPfgm25QMx6bJYaJqPOCq+Gs9f4SCrkVypW22g1LhpMsamyNj
p4x2bN+rl06nC0O+v2PHrT9sFUn8zxlhL/JO8/dYQffeUI4n/DVCyDlDEXxEugJP
0V1HwIIerTRwCl49XmCIL5aCTFxsVxt09xz+1aSZQg2oxoj5VGGu6a8Ztcs8xaVU
KuyUgN5NKc3j5ieMuk5sGJ2kpH/De4nBbxfwpBYqWF9BxCm+5fe675PbCs30djrb
nMi4o6Pf+INi9Tr6BBs2S0d7UZKZY2RSy/jTi7Yo8US//WJR/XWrehFoah5OYI7h
FSc3XgM0JWkqm5NYqeGHDVs/LjaDc2JmxPp2ZgcfjWgUpO1J7/cINE/JwIt3jjWt
pvA4TnEFXgf9kmPBB2IG8dmZl4DLS3iNIGV76UgBYRYRoq5bSxDrnSP9wkWQWeiY
UhZDkvdbxigopK/YEc+eCcOOoMohDNGqYWKqpmzmTVRz+CzoZDqWuMw83K5sJmFo
yvYi/1kzY63OcTbHrEJokpytjRlc17D9/YzdNCi5Tband96s4yCQt2Vgulzxcx15
A4O3zJs2DYS3DVbnEfazts0eQ0wjqo0YJXsyRbR6xaAZ4m7l2hburpn0KStjcJ/e
sGsVnLmApwcr9M2//JS5GfWf1pGX9giNN7PSAs8ZPueC86x5CCtnw/y80cu4zWE9
/7dBWVNBjbgsII5QCSn481vb0nGARxrfjIcHOySTGgpjm0PYLgDgPXJnM/AA1U/A
5LhdVIe4KtfxjOy+vj1uo4aPb9//apy1Gk3ZV004PgiPX0YvmNaiUFENFPH4ovel
ZOxJpOQF7qjQK4PiMn1nicRvG6JZ/CtC8tetMKbqPQZwhg/dslUWiU8vxo2eb4u2
HwjEL1yeYJ1Fapc9UgA749njvywvkY2fxOylKWMo1qVK846uQwKMpA9ZBujEZuql
dlJdWfTQ+hrIVltHRiKDWUwZjZCaVl6VE17Gi63r0zkN8rU+VDBkGiuSBON0Jn18
sFCR6aI/erdiya5VuDA3ODGUknlPyEEqt0G8jCuje55FLtNi/0raJjbDvkFdsyNJ
ybwNrhgNK3a7dIcWwND/evl9R4MzrMnu/GQf1dDBtFJMeQg8CEeHlfWEL0RwWfc5
Fu1UNMqMMp1aEffI0L1I512o5hMTqw92/IK05ZujjXYGd3NH975h2/uPCK8XKmso
sbghK2lh3WIF2llPlXd9xyD6B38X7KWYurU0KGVX0RQfKA8ET8ucIDsgs/Q9OcFf
xKOfIO3GfnH5bfUyTBGwQWdoHVx3AByfDMX6GxZZsfF1JbWXpq9qP+AFkij7MSx3
n8d+4mfLhj4XEEv1tvGC9bSuZb4rFbt9FV543JvPmLAAK7toG91Nqvz7Vp5NNftk
Fu4PsYYXbru0N1yz9GO9o02YiMH5yG9k8RNE6r/fNQ+QJQHWufrUG9p/I/yhfpIQ
+dIWreICeeADOt7Q07h1JBRJmTsEksrB6yGpN05GtIt8kWUM/dObGc7RBlYHCSm4
y3AhUrG5gM+hSdlDdBpg0uZISTwTW19MCsm7huk0GRsacPMvf+siQYIy6iwnayxJ
KVGiBE82xd/n5Q9difn8jvEfo9O8ojbGQRrbGBctXKVAUm/Hixc57WRH5GhqBGnO
r407byYuqdqGSe2/D403loBfhbIoFLpcJiLMkU+n8HGRWL+o0D7REhGy1tzD1rxP
gDP4HTNbcBFhxl88gm/MAD8/N6OjXzeVidt59tMKSx9kEdKbwK72wnT+HYnzAeSc
f8AAdjit8OKrWD0XE5VSnNvlmR1xmdopG+UXXhPJzj/lMMT99yGdkwC357qvdu5f
vtPRXTKcQ7onxhxdUNiq6U0ETPB2MTliCkdrk4zghRGpbj3AifNR7sBHtkMhdupS
aoGUFf4rd+IJW7tzS7XzCVLUSoNoni/6vG+pBJLpgz25z9fRgvUeFeOZARkJvEn5
e9Xf4PcWxUQ6YaZ0c4MH/bW/tVHgmnLIcKihrPT8JM6uj8sHyBzs831q2oO8Rowd
X13NMZLaPV77q1wWdgmuNduyg1qQ9QHpNeOYHCdnmUme7lJYRydNo57QOJ39EMjW
fJ71K3qBh7O8qMU9Rku7tD8ydw2Jnhxirg9tiZuNEQmApwcSG5ArYCEqQoR3D18s
aBDxJseQrd+B3NANsEq2twbRnpBQGt4aqUCyu8aLweUlg9R6RikitpQT4W/Qrp3B
6FGbm3zTpb8z29WAoRTVRqFCGfe0FWpyjIS55weaf3R+5QMwm9HpQdyRX9VcenvK
q4zs8GBCFdU96ppoFQvDCZLeUMndJifNOc3X15ZY1BxVbStpEIjK7M+iU1KexMY8
86IJE5RZEmTfVSZS3LSpp6FwDT3HdqR3wk9g8CXoko26Uv+may5I8NmexBOb4kZr
hwW4VWnj9L8TnXM/HAChUcwzopzUiun6E4xpMu0fOPS9JHHv51wPKMEqpyMvNciw
ZPvPipcUMmOYPrMjKcQ2uuTz7kcGcx4VjpUf6ND+bww9p54HrpXbrYpSdLdOnWsC
E87HjpvkJan059WhV5XDL0vVMipC3+yxWjmJLFPP/SBa4mTiPxswA6bVYbFsN2Xf
dKkrw9se0TWOFrZt2O+BYw8pU4TvpJ2odidmC+FmGF8dKM4XuFuKZPJT4ooZx+yP
IFGvrGpswQa04FYEMLM8dHB/tvXMyhms9QQ3utmo04RjeMBmMxMKeDn2tJ87wzeL
zgQ+nXkKArSZDEGqVHMrsKNewglMAsUIkrQMuoN16naA7aTgYkTUNTN6eFIELZkc
CNq3/qGYygMLwrhGwZOQHt8JH7nxIIHzAetEuJSom2eJ2vorxTAu2keUbtLfcRK1
m3O3Y0Wq6BvyP8qzZP+XGCMr4lekz3ws/vF8HQ76k8GGpyoV69AnkPJJerDz9KqU
Cs6HmNHQuhM5lSYjHtRoKN8zCU+B+wzvGDS2Tz3jumqSzR1xU1ue814E/tm5UYj/
0GpWS6LR0oV3j7M2BTpot7Vv1qSM7feyUiVgjQ63xEiIt6zgjFmUm7aWK0aqYkMS
k/BTM5Eq1fw6TNqylZvOYS6QQmeZ3DiQnXsrlPPqh8XbazV5oX8hwLqSKsoy1f7w
u3YrS+1izmkQ8hJbeUEJSL2o7O3S1W9BYLsiHCRw66eNhDj+ne/4K+UUBOOW/g43
11FoaxcRyCWeGNZkM8LWhG/aN5UaawyHg+k9fMb9mnhmMz1LmeD750r2GHsYP91Q
xWXWbdA2E2HB3u+/NhAk+n9oSH5OnAhSFMZKyGFuGj5UnxLKU4pfuxkaqQ5RFxu3
L3sYv0Bk3sPn0kFsky5FYj2anpK62K3Bzco+7WUmQztHV4WRIaR2OFHKU+t/Xtoo
djMd+jC0ao4Q/i+hEiX1Mx8TQwmBQoUaHLnjWXXe32pmO6CwxTLCfn2wfz3dlbDk
juwUm9KSttnzjUm+nYVkKcP7N+jUCFQOP/voLOzoiDWl4KrHVlGB46Ph3RRoYHfR
Ydy1p+FXN6fakSFSGne5w3B+uVYz6FVpuN7ivz4PGWIdg6P8/bwfy3SAsWOfotg2
khd5S+RNoqYh++vkMhF518sbim2ghn6iaK0GTd6jpHBqQ/tyviqFtsDO+Mlke7W3
skC+ZyxaVpjc+w5y2ZnYOPcxgE9oBuPYMFWLyoFOlcKR3ZwZMExV8KQHUH5uAU7O
5IqsquFIp9rIcRb/cKeLnfNGhYBVA/CHgBvNgRJ9iZA+O1g55H4DBqhk2hzwTmW5
9mD6LrGsdu3EZjele76GjZWT9pWVNwbcE38ZHirP8hAZCvihbnnv//rOnDvyMrYs
YSntthguHFHH6tDKjQEfOX1svXB55a1yWNj7pOwABmI+dckzGI+igeU8BKkN2du7
7lXRylkrbMV2t4YCtwGWd2mDzOkr/pKCuBLLjLbDWCjel7Zd64MVq84KMr1+sDmG
wmlvCXWzcT0oNz9cYvVGiuxRpS7OLxiV48yfLB6vHKyyilUPZlwCgu2rTGmsv/Lh
DKw+Fn6XSzVBoqLe+iV53rJWQJP+E6NTiES8GfT5NKcQY9/wXn0FAOnpMy/em3Yq
dKMH/7CiNj3VhOPLY+hJGKXP47eNDQ8bmVLuPIm0gNH+iZWkxnfUqZvtIc+CWA6z
IazPZoUbk+IoxS69AE7SjbnkuvCsk5UKAgC6FCdAwEkfK/rxJFBIeMO2bwYQikM9
AsBPJs74NXdi6iwLsSKhlR/8nHVQMZA2O9DGmAbyix9/aGgdmrWHHaDqqCE9iybT
dNkCDckgzr+X/K0ev07RDJuzQLUO8CBoeDLtdP9NZ/tYyqLKCNIMy4+XGIZoacxp
1+MjyXUAZ4V/jO++IGxxm88z+liu2C6d2ULB0aPVlfTNx0fEe16MhCMRdEnT5TnI
QW1jZinD6DWAHBFt93IMXp5XP2yisYZNeycpE3M+7Z8oOlGdZ+Rjd3U7QOiEMsdR
70rf9zqKzAefwdicsIBi+LAZgJPh9OBk7VgEqCPQibw7PoQ1qymH47T4Vm+pH0CH
wMG3beA7kTKRIpfIEtGw4QyRzGduLVgmueb/TNQuKlVUoOIcrQwh0Tp+mVAIQUdu
PRFJ6B9lIjbB7PdIRtFEnTxWInrLT2I2cHTUlRcf4tyyMwMNRa877Zwui2q1+a+/
ne+DYk1vVNzO9iyMxZKthDKysrEWHRUsxd3POeglbGw5HDjMZ+EHwkPIG1Z9wg4u
OJPdL+WmNhxhV5VVLR8K0Cb/whuCBelA14EgeD1uRmPfZ9xOIgLcCzVtR6O855wg
sdVuem1IJ5G4NLdVsqohHLI6jUZ3+UHO3fvmfMzSXe+k4ok/9l5Sf4qJC3TI0f3i
YCf82sLpKf8gXt6CcUGyEYfx5cfyYtMPCPeirupv9NOk9iDmSIjpLbhog68zCUBk
Ytnitf2cWBDzYEi4u/kOe7GcY7y/4B44dENXRrrXXLil8Fcl02ufPj80b3XYZnQ3
edP3hgD02bOq7c31yAGX5jNZ5wx/BFb6Z4DsuYgpjpBzIN2VWU/on3zNjbjOG4lM
YU0flRPiSpLjxixUG0/Xs7OGOaEGJBQLSEzMUW950Bh+uZHOHa1HN2A5g1K11OlP
WCgb17I1gz9h11+U6Xm/4YkwZUNM/cTjzQWndGzHaBl534iAVtSBss8GyVZHG2vj
D2KUELULcf4N+ONH9cjTXsypSkoHBR/15UiCybjh8XgDJVb0FMOyyc1vVApHWG8g
wApKOIm4wXZxHMhfVrVFzH/dgQNAVUcP5EOAtm4IWBwxjxDsDhwxwU0M6dyqvQ/K
S74ePPSsKCGQ5qx4X6bcYTQ8F5rc+Oum6AzxRqeCoPfRM8RWNY4hOZKuMmZeZpC8
2eJlp4hx4MJ4cc49M9k2DExws1DR8UmXGv7rg+ROZ3s0IfC/nAgYKqDBWZk2QBge
mlMZGkotaKv7PmzpGvWQHgKN5wekkyh4EovPdBcEHqVadJ5JZW8a52uRRxlsHd6o
g5xvoCLTRts+PwsYMm0nrABMiu1Dv8wyvzi4JlvrJtVxSdX5nPZdTM8NIAgpDe+B
8Ch9E7JYETuKX/DWn3b2BcMwX3LMKrnl2tHQcdLFwIbLuLuoptcFA0hkSMBc9CDC
AO2blhuF3EOEkWOy/p7FkfrPFMznJMJ0bZGeqE52qzQ1s4ee8W9V7DI/jzZfTwme
Q5nhCcMywUxL/5v/zDPgaOym59DzrOu6azFS30akc+gX79+jsuQ1t6i8HTWuZWyL
d0DJZFWVicth3PfrlmUOU8pjA5ShtfuKQJEJIy/d4PfIFjVYQUQdhek3JmP+vUv5
l3Uq9jd3j1iHuucIYsEAO9J5BzaP6wPVlUT8vwabFVs0Ek1jyB1Xt3r+YqgYGM7M
8p0Nh7yKxL+2gqe3VT86iag1S7mq5iZD8hnXczfpdNPwpwYNDxkTdRvP/qiqpT9B
eU66EKTxRDM/l5/zBfdFhiDVDrcoTVZoV5q2HG6hpD0XxHE3ds0ewYPJc0e1e8Bu
zN7OQcUd6Q+67rgFR875DfUVxtdrM06v83eXXcGMLduGoA4DsYCiDHuAg5RRvJ/r
fKrCtAyzRgEWQgYU4sfRCbyCBmtAhOVSAzGHFhU35kM4d9oo2DcJzTCwN2v3RZue
HzLxIoDIKWYxPO55pzDzf18So5HeMQWDvewS6UchHxKWDPZYhTdeu+zKuFpz7sUQ
F7i6r9b0pD53HNY8r/4/QwmRfDzaWk22Qw+T8lAuLGRV89kQBUmZ4M63sa8qtYI8
+BvBPo1I4BjES9wC+Vdzu/LJJD+8j9UON/v+7zB65xZ2qkFiiQtyxwUOwGh0aVwl
ED8d00BE+Np0+Hk755VcU02OioK3ugKp4tOGU51YNLnHb+5ugIA/3JAUfJL6y75M
IzDfuw9MhSQmGN7B+u0CFRXeZSe8lwvfOB9cZhcIb11XQloUtMylEGGjodnkbg/y
ujtjdka0XI4sfKbCKD4dgbit3RTvjco7qg3gMw9CbM7haA5MOkbJJzKrU7T8o2QI
2zBXb5cjiyv700WooPh+dG5HD5MhD20Hsr+w6FzHc6gb/O4cq9+FxcUNGmX1Pn+l
dQRXhz8qbE579Bey6UNPKgEMoz2Duw0JY4/wr/Xg59qeuwcZn1cmh/5X7c8SUT7D
oEKOLo/Wxi2EvMTGVpBXW8Nkb0J9UtD85dk9O+pJwsmWzp61J1ZM72W0c3MYnXVT
ckxtdodI6CIIi8YwB2NO/heIQMIJbWtEycwLvRM9sEUbqSuQt1ripLkSYAeHdJal
Xuw9AVPRZ0KpuNol2PP0mo+C761xSsEbyTxcvrqtNVfy+zlJSIw+Lf0pesP4lh2O
G1mm2+WFfmOSWP3JWJcC+OPK9Wjq595ILdNMTdEmNOE+j3AtsCaR6bGTNTiUrJad
2uaftzm6KYkyEjZrN51GLA/3uYjKS6hbXzB81PI+z5c2AlE2+JFIrXioXDRE/g7t
iM3TBGqyjq8FoiGpfUw96MVsqnlU0pFAa7ikbUBKtxzS1/GwaMsnTLmlCg3mikyP
4DF/yEX9GwBrdN+0rd6ydCGpv9oRMo5dtvWvulqx4waWRnOuH3IvIXSKm6SEhX90
J9sEMFfnS2Vph5PzZ9wiYIDmbUwLkSGHLJiuR/eORJQd8twk/Rh444zxxnBhL7xv
tQ4Wt0zXayGdlELUJ0Fu3lwlMwZf9p6kzxLlAYP9x3CZUoXp+4/rBWwEdukSwSql
FJgB6VoBVwQ4qzXThZzhOsyCWzZwzRheMpG+j/pcK6W3cMXhO6mcUp2dMmlHYhqv
OLyOF8gZ6iwGwsvfB+xf7IORJhBU7gcETBdn2UT8LNXFQPRYjZXZK+0/WsK0aWKQ
VQL5sCAhlxT/X1ueHHXr3sC63qQH7DxjGejKyxcL68ZvxuiTuZx/5vfH60LD+T5p
59B8vdUHXIsNaV5dKzUmWKvHOumK/SvLj41jMYoaD1Jxgj5kQUPpyjfTw5gDoXQ4
MUeQ39597vGLs7VGGrfvo6FO2/gxxfid8jLKpqU7t49cXS7AdDsmHYckGg98+Hjh
343vNTEZdsuOWiqcbQsox0ofaqYugd6iNghyz+yr8n1YAOcOzPFb3WE9DAL/so9a
OnMwpEGj6KkOuA3rdnm/O2f5G3TpBeKWx5eMbbgP1qH81/XGrejJDxNdBt0O6ThD
Kp2H8P/F9MOegoWvZIVt5QZVZ6sZMNaKF50STBdWhTfqpvZLpBww/xL4p6Zr2yzk
yqpUlut8BtIlOfWnNtDXHbJ3Qp2qvYonaSEtN1ux60zrQUEpv/vS9HT5yDMzveJX
EcwKU1aYECR9QlHPU//vDWcKfwwF1rxrF1rBmpJogo4Bt76T9XnW4poj3LLy469j
Ky6tUc08uTqNRnFJPvC2zTiz90v13XwVfVtw/znDB9oXrCOsvgpfy+d/dzwaVOQu
gIQ6JONw2M590mc7hLKjuay5ExI7Zew173uPFB3xPmo8mXjH6/KyEi0fFNecrz9H
OPxrHXWqyMZu6dJF3ngJg91MO3wgwdqzR3+1crH/N241IQNUPY29XC3kUYvNkfZ7
0hhSpG1nFdv8sEYhATKakHseDb1hg7NiF1Cn3xqzQMZTX4zdXNMZbVSBvhxfmD8j
rwwOcG9MYIubbdkYIMi3n/WzMJzFHGAOuluP49/rHTFmWlV7uM16S4lJQP33U5+W
r++izV1bkyR4e4AeBcmQpv8oWnSXvafDDtbBnSnbmAfHXlx+YXzeC3U50auZLPT2
jUoA8S+cKzqg+A2P3Y0BIV7bdqUDMgwvBCbmHiTsx8RymIryZm6urxB4e6A9cnpe
2FcERZPFbz4le47+fPY3BIqhY6LKS/46DYl7nh9dVu6/n3yE6E0p2ymhbjmq2oTo
xxZWfkZy69cGhQiRSBDzgQQORYJUo5wg2Da0y0wFLjL1HlzzyOn45vhyza/GG3f9
YQTPok0rWe1GSbsArnPj4Z1rYiXeJriOQOch+cRIt5RTXQOwD/Mfzngxy0s942hm
yK2ibqhkgOv/bf5cmi9j1ktm+MrWq/bxwiRg2Cu2FXC+j3/qkEAdVCTH39JMPx1f
d7r/sferOX4Jh5AZW2Srp15ETveXrDgRQS8A2+sG7QBg7kXwilCPTiVI9vrTcnKH
8GRc4K60oDRRi9zdeHXgAmab6yWcn8KfsaZaxVPiLPajEEwC6uaAvjBFxh37z42h
PxlhXyo4vvACGQ72sM2RUk3TpXC7L/Ur2R3L9aiPPQDacMmxZpqxoLGJgDcAh/+S
kAWcQI94m2OOnvNp1L0B8IdACfW9aXqXl6j4u1OPrC40Pmypt1SaQ1t5Nw7yb6CO
5ocgQCZAMVHPAqTUnVsbvZCvBqm+2xnsrCnuQF2SBM6FGMB8ECGC1QPD1NOnH6rb
briUs1AEZ7m07ZaVfE0HRlYi4UdTmCJ6PCVcUYgVNqYnG8IAEyyU3p/CDXMLdyUx
8xuul4o5POkXTqCdQ0Vdb0TXyU15j3ccIj0Lm2cQnJ33Xbz1FCMlaeT4Y+lj0eqS
WSgXdzb+IN92+bLYAXZ1hOHl0j4tkkZDSiNJRhKGFmasXO61EoBFFNmadgvaJSvW
2HYi4mGy2CSGEBdLM3EqNmWCodV8cUjZc5D/JyWGS/6nH18oLtqaWya80bCrd/Id
AZ3k0G+T31/7QB0twx3aLLwY9l9w76WS76v0DNI31JSYO0Fp7UyGugdK3czw49zm
/lTWdx26DehdU+WSsLuhliTOQjoF1jvy+WV9pz3Vm+jlAg6IFL5rSwLCNF2xLCH/
/FlNloAsSMr4n4zoiHoQI3DdL2iEC4F4Z5ue+KHyXVokkJJ9BhI7wWIm8KI8v8oh
0gvaolHKRtHmVV1Ja2jCn8zTqhs8X6NtsyyB7zZcoxRiRZ8aotnMKKt9rixCMhD5
EVMtJo1jmSPea/SdZju0lxj/Pav02ZwH1zFM5ybOMw0+v4tuyTZNoUgEINITq5iE
ORgPJduJV2lgVzRyHVJ3pvaUI9Ysb++AxKm6jqKkAZ7EQ2wRulBRFSVqnySsQYi1
57Wxf2QVi560zRR4c931g/0utBplzuFMiHvfP7UiIxUNSVHbFxuClgDWYHu23YpL
3ctXh6cqgcKUKsWwR3U0uwbHtveI2/MgpG/I4N5GTmTlPNIzWYX7t5ZnhPKcUikG
lwANbgp16E+nLRkhS9jrSVUXbi01SNhncm16zUXK1Ao2YJk1GrYeJm9i5B0Jx39i
MS4A0vbr5kK/4a0mXV/BCtoswFyTIdiJY8K1lnJJN30tG+YDSHCgHq3YnzKgo4je
BWpmd2jOEEebPMtpUaWZfsEQZ8V2xdXULxhF252FQimDL2vWsmB3nfGe1SVoW1qK
lF+IuIntZnNzplQ8L6QNq2dgcEZW0Dd5P41IOV2efsT+70P/+0/cSVLM2W5q3eR5
zb+OXQGQ5O0vNGx+67cK6x4d6oPXgtHSZuC9Mk7dOrAO9Mi4z1DlsYQevl0JtFA9
mEppMwbjJD9Btt1poZ69MikNW36Jn5kPoD60OxFZ8uG9kV/1HIwMI9j983AVkdEH
NbpTWO2M1l1gDWQnfoKSqMmejTSCMBjySkmKf4ggvTiAotQ98b7DIeNPrHNGrZRN
WwSvOMu0Z4I3sf8qPJHy2S6T0d5utQYFNddq7SoypbjvulQ97tIsDqe738Nxwx2+
PILjRoyXfmGtfUwbRsTreALRXvFLEgksK0k+HBUK/ESME1djHZNtQGmGavIBo566
nif04b8LbqFEqtlcNvpmzQubAGAJaym9gkWNmn/bFHmK0C40YaD0dHlxGXQ+OLa7
h+sgyw5k7Pfl9S8aRsmfUCaESjsAJ6KCcYCCC03s9DL1kGi95sDLQ1DveYNhDbOA
yyJh49RJUJdPy9DXeayxToGJlsbZjERHaqay7vJDCShFQLhtJOMR1oiS9c+RRElF
eDPw0QqUasTLibokUz0ajTgAj5UfnDUHctnHJO+vvpxxbmi+xdgaqK1/gfiH0WIY
OXVXH2Zt+VFNDVskZCc0l0SGPg195s181SBAp2pWQx+stJaY0riwoyCUw9VyoqA3
J/RJX41A/4otexwfGilgR+zK2GdkkraSyYbWzysvlT690vXHAd5lM9i9CI02iv7B
0ew19P32LWsPdGyerLw7wwHKdbm5YtGXE0yskf9P73Z30HtOA4T2uMdSyd3rey5+
lpKA0lJuA2JO5bHUhNdGkl44/wsaSgL2yJOFXuixOJABVgIVahUwoZ4NDFY6pZ3N
1Ub5I+wuiBBNKNFrnbdIHZoTtCNXdQ781jkM4f4V5j4I8csppI+5DCm2vebFpJu0
UoUQEOGelTOS7Hrn0NYIXkc3uwymjaU3457V+8PDs7ZGzXcGOK6/iXp9DZhN0iNc
wGO0P3csN6dTI5UVUYTfw03A746gkuYjFJKNkJA2JW/LpQ9WChQlO6efZWlvggeH
z2HpsT3JIZk46Bu578qcnW5SWeqOAyLxX8wgK+g+pYYCDUoraKChxA/NT/frczDD
Rnb9hEfx6UqZjde9ygbWkOH0+uI55grNh7fXlbIvfab33vvIo/j6NxXrbe+GTteD
2A5XtS+235jrj4001wx/jBLrTYz1p7wK8q1e6ds1v0kG6JR1TP8sWFRv9kzmX2RM
YhqSSexHjS+N/KPF29pmSAYhsuidHQI9TeZ6u3tGvcGellL5d+Dc44Hgy+uYikDv
ybptxXvi60gZF8ZNzg6ADe/rxJMkJ4cyMt+Bql9U/vLhAPGBfezi8FmQaQlAiPEY
fMBBUvzS1OwcgVJoE8kYwstATDWL+JA/stpXOFKhOKqicsML1S0M9YGWGiRC9cse
eqCJvdqse8OGXAV7VGXv0BMZB3uiE+8GHIrrJZNszjVAPiTyprhFYWQ1+pYrXLw2
jdn97F6yoEMD8sSH0dSmXq0zZLBKN9gJJhzU3f0brZhOnV/BhgBeqsK+FA0/6ybV
v1x9oIuZMM4d3OimWLlgbVTN0fFWOrWVnG+c+WjDkSi0xt9tDM8hO5+FStbb/4ja
A4XjbDTIVMTgeCC7zaeWUgK6TUlxzpPAg/4Q7MO5TG6lWShF4ZHeWmJ920exTdDt
dPmiOZe8A1D7W3CVOUjz8oGqpQd9d3exNr40df0obLbMuYo/9hj5dq2i8pFBdQJb
at/saiD/BnwKQeyLqoEbQOI1UbvSTLIP29sahP3ET3FuHaWLwtKd5j3FJFHZipQw
eHyuM5XKIyf98aCdzznmqZCGnmiRPr4VB9XQQDLEGlXRv1oOYV58YksWhvCEnLai
HuMFBP27STm2Hu4JLB1uJAlI3oec7vFZ+hEausThUswII3F8kS6RXgEoGDvCopzW
yfiIYaCzSXLKhUOlP9tyU4kG14cZqduU2k75CelfCk4cxGroFwaDdWrfXRAcCyPA
H3snGUJI+flBh5z4Pg95RqpWh/ha2TTbdtapiuG4Wu+pWPRxbYo+j6UWgdxRJSeA
UBf36Fw05qwlpmcxllefQiT2rmVYHJVJkG5gxhQjix+CAjdljXkcF7sdB/s6VP8s
c5BECD/153GD2H0RobsrZ3ZKNYxooO3ykDyJJFW3717YA7Ty9Uc76EddNr0ObmwU
IauwzWmD4ZfdgZMw3plPNDliljdqkkRCh33GTgCcz/1/T8ZxNuc+Q1ZmYtVvcFVs
5flxK58CvRSIHa7gLPdeFvqWblgzvphMY1btJI8P8GJwfmD+nSKOEmZVo+HXkxr6
7m58WThBp6HrnSbIPotm7NJIApnlHcnG2V7tD3IyLARvbWOiQcbjTj8h8KlWyJwK
3H2Dugx99y+6SpsH5DFQ8nATeCnwzhCOlmK/l4fWhfRkJo+6cCCpmR3XNrblB756
Wk+KKs3vcYyHb3Lw9NPLE/4GcNaDchH34xrEzkpCJTvzfz2qF9TuX8zM3xFemgeJ
dPfGlriSfNtmHLX7uMaBU1CBdyJQCYkX4DBELH1hXLL6xyVNJGKVU5NSr6Am+lUa
RBHyBe7uOJ5Zc0J6WhE+03+zYUGQ+PU6vBngCMJ70iyDsLE80VklUNS5UUEZLMEo
eX9dgRvDHLM2DpX5lhw/BxyT7LRHk/CvF++ehZWl3lhX5+HNiUOksY6AxU5U8wEm
plkSsEs4yOpZPmOVGFMh9bYXIXc9I5oY2VSXJOCDwA1HyCDKC2mlUoknwEF9tVHi
czocYLqtdCsvGQGxNAaekWncWYKjPkQ8GC31tRkKShpwd79s9naKEHo0l+LVOXtq
ZPIoAnzuH6BvhIgnagdd+kmp1FrQv/EXTWCWrx6C8N/L5ivGTYX78ideqhxTRvIZ
zDMKv8W1GpYDTXMCwt1psuWB9guzT62pwmIZl5XeSJVL/LWcsRVeQ7UdmTZ6vxpZ
CGQhZjdaP/tG7j26LB5VjQmvsFrDsycEV6aleNd/SWa9xjIuy3z4/8hSxSlD1J46
FIwybqP2I0HLN+oXKhjpy2akgHdEfqsXB93pDB7e0v4XX+MmKzgOWD5kl6uL4Ail
/jIH4htdzZRFTxaTBxqDLD6CW43FwkZFBYaJbPHCErWM8b1K3pDGnBmpetyPIgsr
15xQ2wGLnJUNJfzoXJXhBwLWb0EgBqOmbXVd87TqwAMKIvfysLS+hZtgMoFyPxpc
kj0InGH4s0S/wRSsZWUTAnw3jD0AO86379/YUsXGtQeI3Qalg5q70OTDlIMEmBO3
JuqNbGf+bcSoRIAxxEDkEBwJUzL8VxtaD2Y6Jne+9J4MuVuywTM9TeVPyWF0dZvH
LuNq0aG5YWSVNdMzXRRWYldzR3MrUnQ1YKeVjtsLtcGfghXYt1ITBmQwdSURm4Od
uJ2DhuJ07zTKVSGIntko6ZxmrgRL7A40bWdGfcgvuGRaZewHf5s/il8ZaGjgnTs7
9lghiDTgNzx7AmnwRg+zHppzR6J7bvwgVqQ2El43NY913Nc66/aOC7YTpgIcoLNG
tNAVnJsDWGClLro0DsTRPutW0oGhHJK7VW/T/FiDPT/62MKCohdBbFGNio9o6LXt
+AdfndIPMlI+vtTifggDBakT3xlFcLlM8qyXek2jRZKGe5lvFbR45BbjnVwDGevs
hAB3l6yA5cfZQ8g7P2eqtXPMUqwrEKimupnEc8FBJky6zOoGFVB3yyZurwmdmjWp
Pmy6DqLWsQ42grMHRf8z2QUl15nLDw1DonG79PewLcc432SuQe553nNd98cBDC5l
zU2D4XbF12U5zW26hRinRyZFGHgUdZSzvDg3UOsAF84DVHvV2BmQw+fq2Sc8bkLU
m7QpuIR/6zKYTm+yDKW5mAErHKTLGJNJp03Ow5XFvf6/m0QZr5lFPAgqyCxBBOhF
/j48lEaSKs/N23yj8nnR5DOy4wCojwd61PqekzICk0HzPWfZA+7V8En0gQTWyv8j
6JUolSKeAgZCyYlyOP476CuuFBs0OfAb/lVPe8P4DTHOHmbpwDyah/K86Hfib2hm
pjl4W8S0LK9RgWcIxcVm1Zl6r/HfHkJrlfX/fWPKlaCCPTOGngay6FP2SE/3ZZMT
hxTxpXi9JG2QLQr1hYnIqKBZz0HI/X+R6WhdpdSKSXYfSKs5nlpEz3+6iW5XxITy
KOpldC4WgQp1qXMXPcDw9S7Hbt/HOPMP3ThFVubbmTlxOtGNjCOLEtaGvXxGzyIm
NePBGQT8uwy7IRmh2jjhMzcLDja+pZyaU4zdu5AkzJrYQF+craPmCNWAqzK1+o0M
sX12k4vM+V8a3Sf+nlindYOOnQMTr9N+OJlcyER4GIqOuqXA1LDUA6qQOwAQwBOd
h+aWBWPC3DeIecMWGvXAIKXxw6HfrZkQI2u70XX3yWBTDQWaZBaMJHAjcNOnFkXV
O3DSwyC/TB3NzcUt27y9rs09/3odeW9NyFKpI9s0CMkwRa/8OHmk8sYb54//brR8
imZ1eRGClhauWlgEiMvYQDPb7x06cHvgLLaOy/Wb9+9fwGjUp7leM8zGdXWh76Yl
/UVZiSpWAZXHh1R18cvHhvnue5FHzVVpqakdjHJ8FvdOCx513guTnewxkiXFX0qt
+6plN+xR0R00artsvYPq6fsdop61xkv4kj7LaeNkGTqHZtxLwgWiO7aUnC+lg+ax
SqFMJrXRUzx3CQyaMPmUBNf02b/AudFOndzCN2m3u8Ti+VpT1et5Jpvs+X/oCb6S
+FD20h52k/e+S6etQ4ncHkNrecAeIs1DLeN2zILnxp+aI31jfYiVMQEisPIguWk3
clyd3/NuD8xcSOLtXKss6OqzrX1Lmyw0xlE0WyFSy2zZSTpfducYw/U0cH+C5RsY
nxB4GSzN+YTlBMqpjVKYzAMidisgZdJVWFCQ6k47fvd2AYpGD/vA/NCgpzFM30qC
gtmFeA8dmkz+Z0bY++SJgbjKWnK+hI3Mvf4WsBj0h+ynWerVD7c92JC3t5VZBPAQ
gd9qacWJltAEX/HvGO1BDypNDkX514+w9fpfV1qfpUWjOD4Ik8zWs27iIEo7x/l7
DX6v+K1uDN9qTfK2KJZd3GO4dvgJ+3AgZc61O/74yZI=
`protect END_PROTECTED
