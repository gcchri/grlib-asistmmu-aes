`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IfUzepFYK/KKAVmjBu8iq9MKLN14rlx45KKoAwdau1z/QMJBN3e2XHuxP6XTP2gj
97SPrMX8P/s07LIlezhnRNvv7t4q3I+alE2a8LMP7ruVWpDaG+MhHOTz2jHWepGa
Oya3YZ8XAGASzjKQC/dKx84FK7R1hje57R76kWZHNIwLHMBASNEIrJAJ7GEs8csQ
7VKdGELo8Zwjcz4ng2sNM08toCKpOjwwJ1o9nInC9AranBmTxxnsOMXctNn0I0Gr
0uO29eM3rmb3TgXwubbZXw0KDYtphLq1U+Kgn6vc9CkIBY75meIJq+udM9eyXHVe
3YhaRQqrOAJJYWfc2ifZ1acQN+1gk10agGHNX+gR0BHlgSvrqsTXh2wtryrxv70F
k2/G2xnoB49caeyGOuO7n6hMbfpphQTmjLHmRe7JabTdGUWbDWxnCeuxyodFSrxi
0BUdQvjKc7jB16Q6WvDNOHY17Aa0AenrmaeJ/I4Dqcxfk41lk1KiglU4EFKIr/Dj
21CEHWB2VxPC2I48lz+q33q2NH5RnEZ4QIj4qr3ctHFa+qYw7s2+mRWpWssJWoUh
6HlCTq1WdL5LFRTN4g5hljC/1kL76sm4fjNY6kqHEl6X9MJsfzw3cLvSAVDjG1xw
EeiNTK03wDRWltBU8qH3bsf73JaDCzvEDj9/zQ3Eb1yUHnzryFSKUXFebWy6nn8G
Ep0LSlVoZSa11xNcEf+SBtHMtc6FqnhXs7HMk+qBkIBOtRuKe09CxPzqS3nFn66+
rC8C5W2VYDavGUIkKOAU10D94ft7cJhqG4tRUYG+j5yW6SIj1uKKj30w8j4LrX8s
lf8bMJUZX3dSzrO1IrMbFH5nsZHocATq3tD1NpsuXWIsCs9KpO+BV4KVrXig+MNb
OHbEbt/zuRq251ZOXHMqKvHsds1YMoRDkD4FFLLD/oHI5aaRpuV576s+ckcjkl+i
KFx2e2y3IuRyYqdy5pZogwXf9UZyUpmtCWeYgZMNiqpBGz8fDUboiaMDzLgnYyD3
OI0Zo5psQmCleefiHoAu0ddeGzWOfFpQP170JkeKRYtHodMF9kd6axfeRQEn4bMY
a3XwbK3wjgAUGhdD4b5WqK2n5gQROfKHEGGBA6O0fO8/weCwx1zwqyxSqRhj9p7j
Dt5IY3fq5F4lGBHkBDAGEhXX08q7ehWNB37JHdn4ZppzNtj3eYcMouBOYKN3bQ9I
qwo7QPEbKS37LAaEDCGbeo2H8jooVttlbMWgdS0opmGA6+e/yDMZq5ZKrRp8zi2V
LXdcoDhYMikP/fNXAO92zrQ25oDivdl+XFZFsGJc1R5ngVlWYUJUtVN4r13IZpWD
pZKNAd0BvW2klDDISpNu5jT/2LaYZhZgDovwUMvZfpHEzKAllNPJ985Zr3R+WW7C
nSwaQ8S98ZgNHGF4S5flOp8dkFXF055VzPNgQDgKN4KIzq1byEo+cP6gJ0aVllhr
hzdWWo0D6KwA6vuIZnNUxVory0Q4PlEVlKosotl4gmvE0R/3XED+vhFQyWtrvmPN
q0rkdSLwC6iVWXEpouwa8J2UatnIHNq2T3s4s8YGEe8vxnBPBZCxY6mDFJ+zzpgt
4XnGwBL5Nylo5vuib6oIWE0y6til2E89k0JpwqvuHKVNNPnpq7U6d+PW8a3PV2lM
4+3T/pj+FlG7OPwHEoU5EiprXnuC/bmhkFsydp9KduAUZs1wfXaIOvYGKsMMlldO
lE8DKURhg3ZOaBmFwT3ZjKUK7VmaSFSpxuPJFvLym9Q+V7Eva4j6wqAhzWNhody7
VcFUHICzgwsiMUMOQe14JAb5DUd6XXJDR+SvH+vbNT/F5B+3CyDgS0m7UQo/oUk2
aU1WbI3psbERuHPSVCKKWU+uLCaM327O3CGqpU+Ob4eSYDIoTEYxwUS3xPj0qA3Q
jOc4po6/3dWBY/AMre/Bxe6Cy7LRtovVWLbtTa6gnhe9DlzxJ3q6DFalh0VEkJSN
OKkZOJz1JezxjdrlMfYp6lnfwSwy3OGimIkCOK+L3CiyPdB7tjoHQ/mQP6uOjBUH
suCx8Y3G80gKfbyjGZ1+TOCckJn9sB3Xt3sbzmUEPtRLPklTjAL5c7FRwl9mWqw8
FqLLl8VJQwC/O2/8mpEt4XuQCtpTQj9EPLY53L6o9d8HUe7ONw4tm7auC8t3HJ6D
j7c0rEu2O7gG8j9YDM5Zgf8X4yc5gbtNqWICAxpGTeO6OJr9TZRDGm/OkHAm1Xpp
dx3FSmCzUzU5mATKwdJlv4hbxenTcmLszsC249N49Ha5qhSEb3x5pZw0MQc1Xcje
8Kl2WwFEcPhk/hicnZOZlXFBRiUDPbzP1n5cF7IENKPE9oLMBGB6oJGUg6n4Cmct
U9SOI7dctil3b866N7qjWHGtAVr/qZ+qi0FUrAUu0tk820cKqm8Qw9h0ZxVHNYZC
H5Yt9msZzpwUM8qpS2zpSVMd++b6YPfuzryLxIKLluF/zHV62BkC9XQBTLpu9jeM
P6gmy28FY6R6V1EfPqDynfZa8kM/0TNQxgB0eDXteWDVMotSovV31+BJtMnErXBn
KwIa2YYOrpMysx4s0W3cNiTgsFNw282CuNVehc0rtL6kLWtOGo+NmYG/NpICE1oP
AntcjxGErUnHZ3q+vV/ssWv2Buy0nJCTb0Uolg4c5q8oPEeVB0W9D8HPZ7l49RDv
XOD2T4FtmK1ZjX6aQSntzftz5c8EHrQhMClY/BLAAL69224VWOOrcMsWf6VvC6Jz
rwQ/Mc7r423QQ3HsSlA+dGtiZWrXtN5Yp5pl8ceDFcuzuvIv3RCqZrJJjDEnB7lj
iy7LNKpefbM7AAugzGQ/2VvWqhFdFWSIlTyTazoQmQjwZAp52wLeHMYs4dJuELJ1
ETskVR+17jyLy13cBmSqk+SD1JeQdlroUA2PbL3DMk03ZB3OVjTlSk9k3i6rgR7E
6FJd95YDrKRRiDNQdD2zl3nqtMnkCD0YVD1sOVkBv3n+66nZU7JWfuI+vc6lRJ5G
BZPs9cA073htrfKEJMQi8Vz5l5aG2gyvX3mPPQPJBxm0Uz72L28L/c7y+sramB/9
pK76yas5bywZA+5JpGponqChyPdtBmWyOYwyKZKuNPm8PIMHnXEnn1fj9ODfW4SK
fHOxFBVyqEocES8LgDTuAV77PICwieG45hzZ9JyOJpviFuKRBg+xuVO+h+kbOt9k
4cxA0rOAdKblAscpdgiWfVOo99EWPtyrwwki4Zt3yEz27PsRubWYEEnH6uP+P1dK
S1SypeMGtT5UYNxQoK7bYOG8OVyiIbIAuWFvOb1KzFUo4GmDkMDU/ZpHkd2HBZqb
5b+4niq843mpm7seb39HjlI94TQeoz3kRBJ9mQ2WTK+XwSo1bWWbnV4JjEZcR145
KeDzdweFJd1Ujcf7jrfs7IKLO2Pk1yC2ND/5wv+z/V36UCglMkKaI7cL25CcYiwN
YgETtP/rWPQ8r7Dz8XXRY8EYTQqfvzznpcTcZKk7zUks3101mhflXUl3hKBtGwUS
zmmgLXi8bYSSThbKPufAbNTjr8oYuCj+kuRnVjk8hmm8eao45YyT5iDylMQUw0CW
xp23Ydvj6vVp9LuCjfXeyorFK3S9vrr0prXAORKI1Y1E/GQBqMXOND8O5DRObNRm
J1akWaJaMLJ1SALONJKYC0R6G6eKN0xX5gG3R/pG2L7ICuqdsrJty6LKDFqRAAZ0
szMvQTjGZQHRqKls2/inL5Kcawr94K20PrBCVKyh9jJUzYHfYGX3w/krrLSfYMqf
GgiKUxzbmd2Kfn7KGdkm7lGmVNHEOJhJPdqGB8UsbSBEhyDt6mFHqAsfhXWjzJj5
GSqOsUbAckXqZnqdJatoIt4pzniFHkxALSHZ8ejPUjtAMNPTSY2EmzMtjyCsT8ty
Nh6QcYQVpU2gQ3/7UMKqwzoMpL1VvVXKU2jYrqgP20Yz9SqXXN8s0MCBZ7zZXcpT
E6XfFVJw7U2suEPo7QQusecpiJFPDwZ/gM06QVi1S7K+CfzcC4nbT4ajZpt4f9Al
6sbaf+ZQXRDjSBMaU/AGX2N2rwyqvYmZHfosh2aDopetAG5qJOrcDX+ba2StEVep
AHN7TnoHW09yvlAss6iuF24l1YKh7PPbT6ZoRNy3VkL6JAkGmdCmWXhJfdWXNswF
hKIUETzfzPXoP/amxLmI38WG3EIuvPY/I80EaI5xDs087PXk7j4/POuV9izvK0PN
AbuDNKZN0bCWlhv3WOUTFAdkauYpbHHtRQ4AdySSMlaxqNP/gd3fwqeTMDkMsbML
jmOy5EWhicy09SWdUekMorbnaz1QLgtx/cEfPJ0V/+s=
`protect END_PROTECTED
