`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHLDk4KAxrDTs7nfUAsG6y2IhwQbwcBqH78MUY0+ZDpkS1TGUQsmOZKWIJuNO8vM
vNnor7TL0G1o5h+TPIpb80kf/6wUXm/YP/v4FyYXadCqMOhScktIzeoO17ileTC9
BHKt61CCbGOO2o8al/MXstBEkwo14hcC1keSLzxzpDL+VYMVhsaP2n9Vn88EP6LE
aAe33QFixWe/QUbtYEOK92ONUHbeNJ6RRgIBdXap+Yv90rdKHPKTfW26anxuuojx
Z8LPmqylecyo1Qp7k3XSNPE+j7Sq56kEkZ93/X9MN/EfmnZvArVxDGDvWJToJr8y
owbjj3ITvxA/dW7IjiMUAQMZRoWc5hq/eOauWzV52am2GoM7bw+UK7M4eAxTbvUq
/tcnl0XHZjo/KxwGu+C95/zHy2Y/pZYx+wbW938QcI0=
`protect END_PROTECTED
