`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4WDx7ASrC+cXc2oA47T+arrsfWzjVT1MPiQ7m5RZInOSr/JBPTJRpTbXVC5BGWt
w6eLdwY1RAY+hc3pG1J/pLGBggfT+OY7s8PTVQaXVakAd2vUY0WFvO/bSllRv8nh
wLKl4e4zlSoX2gPn6BfwXM+C5nhjaSYeutCxjlcIGzw6VDOGNFKadrZfuN4+s43B
6t0m23lmJ+YPynyyMzs5WNiU+5fGy4NEe3FexsBcHddmSwaiBh+9kEDBlh7WA4fQ
O5ZOvPjCtwkhDdnL85kQA77QC2p1b1K1qJzLOGSpZVcKfmY0cbxzrUWm0xluW2Nr
2g776m770hrENjTPcsHiB20y2hOW1xoYcGNo/iXdq/xIRGVuHDhMCQPfEIslHVCZ
`protect END_PROTECTED
