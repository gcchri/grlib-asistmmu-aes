`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s0gROWgWxfsPX+7sEi7pWsEAlsdLZeFvJneUD8WINd0niCm0h3x4ERGONa+v7yJo
8duFvuBcGcsxl4sMfoYvP6MXgSOzRzRpHQ58E5j70e01OL+btw1GVjkT5mq4qb+I
hdYwGIZcarTtSN1D2XaeEZpmf7BWFzjDq9MpIa7k9M6r9XoUVf36FGWJ9qcMPRny
F6T9NGH3c7bCwqa8hITPjwBKrjuKpVlFzOurOR4ZBImQyNgi6VYWpihrXuZcxRL2
fcVFUCecAGGRosH3s0H5g9B4SMx/7YhOfE05jXHZRCBDmps/SJaP8r79/umF4fFZ
Z3BtBLnfZmqzS29CAjoJy92FQvlQB0gdMQJEkgbvkHthwyGWYve4J3kbuTDbuLRr
7y6PODjy12fhxLThe2zywIBYMMgjfx+x08Kbbp1BGVvfKCX738JzEKie7omHUHOV
GdQWBXgMnKTyIUxfR8+7z2WmwqIDH+WoN0EOskjbqiXbenBW1Zs9xQ5nF0A0Wvog
M2xrsNL7mimy7Y1rLZPjbCfsOO02u88VAmqQZixr+pZsXSzzwzKRcimTCZE/sD+L
NdJfWPxUc/F6jxzB0Y2OBy59oDI4+YNE3ZHehMkNJQvSVGjQ1Cb8FwnwAPYBE8To
ni255If0+WFVEeDxHENnDPi4yTZJ4olpONNds1dbCKpJ8YAsYMcB5XBxw+3auB9j
2p61bcf//Y03Kfm2/9XZUuzw5EbnAMuogMz94u4bnIM=
`protect END_PROTECTED
