`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jg+WepdfS7HgdXn7koRIlZ9paYYsX0Jmv35DcK3KC6qnJn5hcmvH8Mqz11pHRQ4T
uSk6Aq4HnXkcaJm/jSY0g1hcUnm7LTPPWtoKF3bSHH0npBXTayMDvtxAmlju00/E
n2yekQlskQGo603BDc6yG+hqODrle2kvZZqlXtuiv8gfSYnbBwwBsi6wp3HTDpKl
IUSPYiJisPLyhM+MFLUVTEK3lWBuLkmQmhS1eNQTBheUOOC1guusBPlt0OLIHhDT
lheBPtzxhfg2Oqp9OxFDa8+5EEo1I4z4PLwpEVtzDmuB/gtQgOjwJdfvf2e4F+Hm
tmN5M+sxYMlt9wvOQEGmQVc41zZvPT8bVOTEcRaVzLQpt3ZNKqXKMIK4mgqVYm4b
FVZPnUhDpTTYAVCuX5LdSxL/EMsiTe/ycygcjNc2Y97+COnFl7/0MlL3FdENBQgm
GybHFWagWn+UjEmak28HmeBa2EqJhbvrzUKuJwciJX5pDRG9YwbN08G9igMetwZS
GYYVkDuynVXf9D9r483Dqau9Rpcr3QI5GKiWgu5WsPGLGvEwcvpSOWzBKlu6ZoXW
F6wTKdFQDLi/sK89TWVy8Sol/4cxRSi1pV01yqfamLFJ0gvZXwud2pfdRHl5gNd0
Ouvs/89KaBAAoj66uyIMdsKGwkrZdDK7BAHY4b5UVIWgxeSHQpG/Dnp9ZpbHlhe5
DTtcX6DXr6pZXngA8igKIz4P9FV8hZHi6GZVSPKruDccpGe4zZT+o5KPRRbgKu2i
7W74vwswCCQz8jlguAL5urcRdNA26Wprr/tyuMHSMyW75oscoCXjdCF3YPKfKCb/
Rl7qnVZ+tcZeMyMwODpXijuExmMHpSaCHPgYc0Utckvt1t3lRWx4a8Mn54yZD0nw
M5Aby/+uCH57MC3bPwc99CzkrAIItgNOXE3aHDWnnbOJO1+dYLzMKzEzSdI/3Bu1
FONndpdsvpls5SKH2xGzk1TCqQ3Vk41u+TRzeAi18H2TaMmze9wjxBzU/Jep8529
jCa8J+Yt1BfVISEyKGnphGEDOLr41n91rgjV3F94HGBIP+OqiElecloR65cIuGO+
ppcQguUA46vjLPZ0cSLyO2/rnBcSabJq0vcHRDG1NC1swsz1DFIgZXZk7r5hMxzf
rpeqCuWMMbet3IMAgXwFPcU8AxsofgLAng1tht1ocZsX9z8dn6WtxAdGZ8pHg2jn
nAwNykALqVs2imi+7YZwuhkd6noEOIfN0/lnUqmjFq2BuF2xG4hhMyayhpKjoT6t
nar9V/i5ya/j5Dnqts7f4mjhOP32xJRLgptMKaU5gZgAD+CXVV9l52cLlPlyANJQ
PyCz6+W6onCVEQShMZeSqjwfzH4idotWdilp1UUy1PSJISYWR3rHbwTtg8Ry/pGi
wlu8lrDBIdVOEwIyVju0B4DqaedLqXLrc0BBRQPRm8qWLcEH41HZ9sdJaq70udJC
Y8nIPcXgT98FwUj1Dl0/5MR6rBLA3NX5yaoVKx873ff46t9zpLfIM30wolamj2mj
WWrEDaiLSGRboRfGcPQMYeD3Z57XVgvb8KKHiXqGiquGlgVanEuVzEKmErkQnmRO
WzLDt0A4AeJVClk0vNYLga6EIBGaF/804EnIz33e42Kkgv6cKTN1D7EvR42FGy5V
SEuXAZhKx+/hzKhImlQvNzGw8064PdHJ9+ZlJJ+lHgHVcoEdRt1Tfsc6M191kJE6
WXMeosicrELQr2c+RRHqXaAfReIoDIKe+oQVMGjkzEAaXB1z4njJKtRlGuDSsLBq
yghv8cwK13pTO4Nd7EwaQIjueBuMMbc7Zwz0XWGJVxDipqL2PmQbehFcO20sui8A
sNEY+W44B13vrhgG0cQC66xlPLZw0B/rZ8siDd2xNGFP8aBdqZMmtjb1HMFD/MCb
n+iWEMLx2hUH4xivT8blIXukKeRCietNfRS5MOhZxG68P9+A/uYvz2xbUtVBiSHt
Y7bQCClO+llxBGFUo+QHYVEHOiIDCE3WRIgDMf0MqULuH46xA+oQIu8udRwVs9Q2
q4MmkSu6jq3CWmCZ2pzeQlOeBC249BTrn4ywnsLW7JNlPI9ImLuQTflzCCSh/VV8
h7mPZq9SwnFYF6pGghzKAbszvpkKJzmqGNNENQDMALvtnHOHUvm1Rg0m6/5QH/+Q
PrKYuX/Xkl4a2IcI9yzObcZznzLD3moabVYGiI7P6aDFSP3gB1IvS5H969NuZZre
cNm40AmYpSWG6B8besCRh1p84PDsZDP2toMcyxrURaIMNVIP9DQcOcFnH65MxSct
XFYf5LoeEWw+GpjqfTyAZLC7T6fUeL0wFi25r88dUBeJpAI0XDpw/PXG9q++9Hob
qFEIvq9rGQOzdfLpsrGy/PMCt5dg7FAy8sjZWUJrAMWm0ogx2PsTZDnlfM7Wp1Nr
vpxWTaFy6CRjznQRmn7cJ4wU/po7i816pjieE08eAdhiPz+xmKkTTc+c5atbMEP1
jl6P7M47TakfOG9obRZyKa2ZqpoAEsa/SavxLaDA6VIcasp0jPNPndUuwHetCqbw
tb75BzWVwM9xFu4YFkcr/9WlrMuH/yGbnTiCTUUfdvbDMB7jHBfLz/xsKkxmyTKa
jZEZ5o00r3tP90uiEjqPDIYjsuqab+G2w65AiEKJpjz6d/H4d6aEE5vn+GvAVSAg
C1Ho8bp4Oh1qr3Rv7m7qbuAwlU87WFpN0ciplJA3dT+8XMUf6db4lCLv7+RnPydS
82Gti3ZJW9WUgrHrGxKK+g==
`protect END_PROTECTED
