`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5SyNyeKkjGSkNws9Ob0cwt9Y70rcufhLUJjHINW3MO9CuunsmdcLAqp8RiiXuJKU
bk+vn6Kqa3PJoCnmy4Cyck/QmcqYnOmnAvQvEGYq0R+v2CcjkU6f5fUOS1uIYNgN
k//U/SsQNYrt1iXIUfU5EqfNn3ZuJNPFPUUQOUvSE0vAEncTBA3nRxGSdV0VlqaM
n59/+aNKaxDrtgN1DWaABcgBBMQHx579d1S/GzSNjwjq4xeAYVz/CGVhOx0rEJ4t
iN6j5rHGGjUrchdJbwv83M/4Axa02dMefOr+gD0Hrc53GEUvFn89e7uAEq2mAoLF
WnNUWfcwK0Rq2KOEED7lAEHCPiNrJcReeUokRPA188dITDzPc/ti6bTMAi/48Wcu
T1ZzGZ5fBypXFml+HwERTL6DrO9gf9OftBnRKccSTnF0ZLw01OWjAIDASYgGv8nC
59d3HxYNuddUQg3DlJxDXxkawohjvzIeAK6BXN6XtfVo2RA6L6WCZnoy7/josFQc
PRPyblzmTzfrl56qQfMhLnSMpnEVXPO8eJSIgBF1kcxjDcdc2Dubnq4CjAvOM4Gy
h+jWxn1kGRiwcx7Jgh4cBuFAvHnPcKfC+d29G405izsDyia4+Qdtnq4fTcxPhIHV
keQ+5sBplkNT5hMHGMB2TOzx1/2HmiPUP2QlKs28IfN0VcLZm7zjzV9/otXLWYYa
2VfolR7jtgFrJbrZpE601PJuhxnFBI86ALZJXxDgv/hHBz7i7uylflKgbs/2hBoJ
E9kpclAUhJ/7wW3MG1jNOwuUAKD9z8VLpAt1zLY2/6lJMD0JAy5khgCxRQ+sfHKw
ngCd9zQqalcLPBZuBQ/+e/A6uN4R7NE5dUUnSr5GMiMpzpepw8NoLZaM1rvXQnhx
M7AVRq9O9p40Uh7Pk71gBKW1AJ2SoImtuSbQvkjLoT7PtVb86KaRWeHZUSY1r87H
xx2FJMF/5pfO5QWWQk5z0o0v2SyGZZFAXTpz+bch/y98zhokuOUt4O+vHm7dh03c
2AnXOCWM9aIfSPmE9dTOzhHYvw5CI+coEa/KrUFVXvgBTN4p4zHn1+ESinGmF62l
jagjxJ/A+JcZsuxK4vacTJ4c6TA11hAasZ9JwbOOxY6dShATg+YiVQmQagMMmxRO
vEcYFREsIsGCHnQGcFizU3uRnEBj9z1NOEe54dhnl1TpdYkzZ/iUo1w58oxGu1+m
rIhOpL/exWYb7+ytcesO1Rm9pMN4oD/jIp70UMQbIziZ5is9HpLvdvMukYJWhaMm
sjzOc+3XHTluTGnaspTKLnOkO9xZwwZl94c4UbFQMhPCW4GXrEJk86DUN5S7oGXp
8Gj1iJb02wUWVQlTA32cqeA2veN0szsP5FpgUPJcQQsjsT8OMyLV7OQ5ZV9xJ6u0
Vmp6n+2kNYM0VqGrPGuiv0WSuDQqWOhD4y21VcDSAo4+3VEgTqe0LqUZ51/vZso9
ng+1UYJvuKxJY1gPrEDmcy7WxkbgDH9lwXACUMjucpz2KGNCwEIcU3FwE4fsMqBG
vc3UFZxQc3WlOknbh0hIZoUaSgPHwcJcuHuv6PU1jW8dDYHA2cF1ohT8tT24oRP1
Fl5U79mOG+o7O7UUH6b4a12U9r8GWnEdbHfat0I/APcWJHCV2on2/aL0X+pMoYz4
UWkm2g6A1M9xVAzZhsoUPH0+6V/TYSKfXm7PjtgHw/M9uitOYniB1JaufDowkES4
04/rTypkpYX/mY1pBxqCakfkzKnW2cifdotzoQx9P2ZJHfFsyG53SanS3yvYmaTX
IjMXe6/OPBRsOC0LCVKK+nwo3OKUxrpqzMbzaYcvNddGuecEB2VZ20TNdFZSF5pt
Ml+g3FB0t8QlWXLvKuip7VTNdD/edZ1o4Kc+cwlt6MXr/Ijo5lM7YRzbfy+rSrOb
t08A8KBxHHGxADAafrYJIyZklJEz9Hhz387V4NwQHElQUfQucXx5/kXz/W+Qv59A
1anYzlIugfERKo5/yrTReqKAhZ4yQ63Tdp68ff8efMO2gkoviOkR6G1lz7f5MwAW
mXB7odDO3uWaN3Nkc67HPQFnYjYsaaAgypLhom1LGYMlJz3xqrBS3E5k1EYcXEX0
Qi8DC2C4QxqnvjTHscIrxW4JN0hSrNjuiiIMTxfaTGAmi7N84zW03gFj95S5YREI
kJXFJHRn3S3+BXnX38CVjP6Ty55qNCW9xY7z2RLS24g=
`protect END_PROTECTED
