`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jsv83fRx8eMLK8iMIXm/k4PT5FMvfTpHfLU96a8b/3kHoY3SO3fu1uJBeEkHD1kf
iaOgnthtTPzRUkTbCubYFJv/LZC99iuYeIBMFTK61AZa+WxiCpFVfff5xil9VyTl
CUd7M0H4crlkotXjKu535uiaWf3B+YfWPqPCtS0BrfjXv7cSpaNLIbc75QxXme9V
WkX8Tu4hORAKjITKKPFTOz9hbG+ZTWjZUSogXnrjalMWOLqiciXVuG0mWy9JD17U
uemuIJavxdNmNHViAhSMEzgBCWWDhswv2L73938EhOzYM0IC0HqyqnGqj8IyQ/DU
2LF8HOBuoeduicVQ6r7JCd0YaHpCU6azbSGMO+tLFjxwto+LsxKyuKjMqKesz5Vw
Obtj3CbZrQmqFh/L42epDGEidEqQkmqy1vBsDisdMqwZKwyaEnCNqLj9aJuH2I2G
KCB8y17tUfBSx3/U0T9M0q9lb26UZV7M53vNB6U2JNeFBC7sd7tSw00hYU++YTHP
dLcSwiYgBmjv9+1yhB6OMTTLRW6nm+vwklWMb3hdemOOlqZyAdxrEbtIzfhvzvdn
4Dkh4FsnUlJRvTlFtKrmJfxZ8MUdhDx4ZE+aLeht4Uxa7WSf5r/wum+7XkL+g58b
17yLJAoDRarRmDV3EFfg6CKamK1xhmtjkaSUv26Uutw=
`protect END_PROTECTED
