`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twv7RaP65OdVlH3vfb4gZ+aRBJM/REFhjnNEDW1yJlVpiEcwAlfI7ztzMkfV44E5
ftj/W+ffyE6J2oETEWo3Q1GL64dsGJm9Wvf7vlVuCAtFXrh3rN+Ca8QolkhImhUR
bljJRUMywvAk6GHx3f//PXFsBa9RDKSXuOR4OrnI7qjzG+994gnL2YI82FwpBmUq
bTt+7i0doVV4GtOB98ffjKtcBsk950Lqk9IrHZ3kYGXYnErJFh9ryRCRU1Vnuqv1
OQHYZaQTgxTm7vw0Sn7GpsCYAakw9Hdh+gXVoyw5me/n7H5kjNwBJAWzD1qZoGgw
SxGzrWyROWzVyw+BXLNU3zVdHiIuktHP/0HbbH0JEl64QqN4TvLZFXeJsARNEtaH
wfCDocYGQRU7GsGIdVark7RysJNbRP8uUanc6HzhJF1dsrqCxXQ8b/a49gu1qiE3
70Uai/fIi5Lys2DV1ylVpyyDTCmGJ6M0sG8a/iIXDTy1Kr7I/eJcG4kFPQTRYVvu
uAXSJqcSBaqqJNU92D++pJwyzuSryHRjiH/sPJCsnckJrJ+0sLYDVX5kfwOLe7F7
rjJNCdPehBt8pI4+qfHaHV6Szwnt8+0bh6G4ukJRUKjG+M055fPbpuw1FXGVQByQ
cE3Icpyk19IQku6ociXGXwzDfH+xNbntddQM0OfZM/vEIgY+H5MfZlVDjCz6WP3i
djl8Z2ZELkhF1kXGeaRua8hjpSToehe88h/ZEXFTEMbqppbizBQ5YDaKSYQrxfw8
eVQYa2z1zjN9hgVHFEEg5MHXEio8TDdSKYid5P+fPIl39WvswYLGbwPIgNPp5rTS
ouhjw5980f00vkA1Ot1f+EE7SUNM7b7JoQV0vdxhb9T2uHtbz1zVODjLd9lHd1U3
/JZWCcfLJpr8XfT7YZ8zNt4ESmYmIUK7p/m8nMQJM5MKdD/lyHSrdcZa2hADFnMF
8auk7+N4Cr+LFWdN3+GlZlXLdxsK7tBvh1sUbiq1oi6v0owDW3jxzoyELGj5FHvE
4yAYxAadanpAmWPIQ2MXS9uqib2q8T5CmlU3L7emd/Imaxegu3JU9u9jW0WAcgUl
pgKpAcl1VR0rlwIIdh0uXulDUYxlsHzhsgwAnbVgydy2HCZ2n4KLZKYhcl+Andv8
RnyBxgTrZrsaKfY5bn2lYxGBEwPRCLsVSHKoH0zNehG9AfVCIq0/0LzNbeetL+Z2
ZrTMIoEmwRqNkCeAA6WjtfWjqb5ebe6D4MFcAxnRfwptEdvKewNvQBK2vnLwidoC
vghQxUk31Qep7ZJ23FXT+LwOoqteBNh+EfFw5vINL2OXxeRY5BLqBn/uk/6oxy1S
rOYochfHlpqZ40CI4aTGD5KJqW5HSglcNleermkg8aJLXwkSFnUypfviT0Li6xIM
efCbFFeBDr6Duqn4Nv7B3aiEZGj8tssaGQ586TTTGUBhs/4+xwQT1dk9WJu1pNHw
jNVwIa/zC05hPNDy1Mz3pEOmlX4d84ex8OHCngzsXp+eijBl4Zq5QAlnQJhm2fZ5
sPg2xzCk0zx1J6j5l8TFeGT/XCeLayTmp9UzyBBC5DMfVx7X5XHy+8uDiY9uDsm4
SBPDGVcqJIMxxvQbraNyWZE1KIWF6GxFZNJdGAJF1t+tLWxUgkaCp5iLG1FgUom/
i5ttet2uL9A6Nm3K3Y/CBT9MFst8+y569aO1S0BBDn2PBJSawgyOKcjDg6ExARte
LaWWt7PFw7euCE4XCw+ZfjV02uA7bWH0ar1UZIWRgrFsqLasPjXgcPMOmaLuGikH
7uOVL6RB6XGbO8Ctlj6/8mNs9tvYru6MqYyuSDQBmmZw8tvFsaLy+Q30kLArm82Y
Nv0B93G2cr5W+rmgc3Z4hB9iPyMqAT9BcpbsIaJFmVySD+vRrUsnCtjudRnTJMG0
BLxKZjZpLXO5FbBviYf4fz4OllTPFzfHnamieGtsq2S7pSJmM3QJMKV7R6HRW15q
YJ4qIhS57EJdVnTHJyU4bAsBsUi/P73ZWThmSBojEOjn0/bvsxNoKbBGfIHTyeZS
MxkgOnF8Wawk/sTCEmfK/wtAkPE437/tdaJFwv55zOUJ397g63XfE3wcMHHljZrw
N7DMe00bvu7tWslTNvmrjuCIGe/VWSbg/peTkuQUHy/fJIkODkxqAk10v1wRBkBd
40oeWhQ+9IyhqXCyQPmR3bR3JCzMaIAOWF7d3ZZZCkkROPfLCsePbTMP1MGX9JPk
8+qPn+lFYgq8mygCTryQhb8X8Cel34FN76I+/1ciICOxwpPNpxEv1qKJcDckaW+K
1SUYzB1mwemTtRl0eU+Bd0uz/yxJ3Yhb9iFviCA8ntN9eQTIMHm+It/W0SGMdSMS
fVNlpDb2xsQYOAN9Nj49x6/UM29fUJL/4tcYbVi2mTgdWlHrvj/VMAHOWSrg6eXM
OWtQsX4wlO02h21jvi1Oc5ZoTlXHck2tH8/mGROGxmliBRtL5ciQ7CjfU2Z0b+xt
lvdKscoI+GMlyuGzzhmrP4bhvTX5Ckp0WPCRGxPa/vNyUl4zT3ve4/oY0xjwDrH9
Jqj1rbHWNBqiR6uQiNRpdE3jsoDECqNYB+GB4/3bcVT3gRUQnaGOQimBXwGgqZVI
pk5AlfTkfsx03fENumjpNxwWt+gsZxD61KiLf5oaJPTDandAemkKwY+O/UFv8WJ9
eYpbW2LO132IVJqNIjmhKxlQ3d3WLA7Z7seQf5H6atKLBiUOSKhvnqM/5TdU6Dfi
oOHS5VwY2eBO0rvKqm/QYUpdchbplBZRVMZQhceuSlswhx5GGv3oMCW1aPZJ22Fb
yoJ2Gj2lHxEAy8343DL2wbDYSyCYdqUM6uJ+4cUCNSLdHad90Rj2JApalnTNg8uU
JMBC3FwgPlojtxHD9LVHqQgEDjBYvDpPEHc+pEpcP3/cS1gIbrzLk4qnBYhGOBiv
nRtDpaxN0b0fiUObokRDh5/entMgmPX1bmX8SiKlg6Uo0TiN/iPm7TgSknApBPBt
yUMbw/qXFofy8tDpfXoSbOp/ZVJ7CSaKDi7ZdUBxFaFYoeYK1nXit1FRK9tRwkrn
z6j7AWUhK2a2zHSNKQ8NaxZtgF/QhAZPx0rUG9bITxIvZwuAItBOABG1sGC3qU9V
ZIS4es573c6SU5hLXk4DBWG7E1CnhZF/+R23INWhQd7cH8vNBiBtrwmio99olFYT
/qnnFrIdwBnRvHgozWl2cnjA8Nb6quXgUdJYiAWJ87Nh1g+yBFrpsTE4rz/XpgWP
1O763wRG53iGE7N14lov1XtDlJbMMoZTiZPUiyW2AIUzqoxnBiczsM+PW0d0tMgU
0/oW/0NYcLa6+aWksOy2qMPpBhw+RbR7I3iRDQe4+Eqi8Q4eZpjkHOGzvkdl9ZGw
PzeOE+8NFCkUAbh1zOb5mSmxGE5z3/EvU4jNwPYfdCDcbpJ1WXgXaocXky1zKLRH
fQ3NQoJyl/HswFq4JkQwQccFKlVFpKsq1u8JBzcTn+5gHFkp6sBLlHsP19wYXz04
sNdhPDoYjaHzNkxEl185LCZ3dPU9GFsM2EWjaUUuJV7kRBFLSjf9/44N/3cTIT0g
5U7+wMoR53rWL/UsjDyUkempCZaqitVu9xlZFX8WU4peXFJ9K6bkdNdJxqhONYJp
gr1PvAt15jr+Ga10EVJHAY+BvKoHd1Z16oay+UYeyjyAeKpveVlSznF2YT6Eoz7C
s1VhMMms4L0edQ1ozUNWgbtYfojtuLnsjvc86TS9c4sU/vphCd9xCIT2gb2Z55Q9
03E7aJTzM5ykQoPWS919JkR3K3BgC6X4Gfzh6IipSEJ1dvV6dXLIUl3IrEBMdBBN
UQDLSgfliBn6+gsssSLOuSDGo4JKrVx5TMkkoDPMyiRI1uAbgljL7J/5zpSyK/rh
esLz2+phyEU0FqFYeY2URmfvjfYv/A4K9S7SI1BKWrejnLfz08jYcDRdvb3ew8ta
mME4VpvdvIgqoB9svnhJZf3sFLefSjprRMgGVf1bknhBC6sBtKAGUYBH7se7aXxw
dQQz96IQQ+g1QsbegHTr0eKtaDE1kgw35D1jz1+dv5M/67xj0y04lf0wXSSkdGuN
RT0uEKncZ6ElXfuJGGwbQE51d6viCTxgSaqlgz4qh/pkdDns3yDpTgQa+bnl4jsl
FQf+zlb5pQwP7DaDOioRKgk1eSDxFCFMgpLNYge32wbv2nLAUmuaxPeIdcdkwYHP
7rfQporFDq36MOzNESDVePPTORNye7XjjglPFZjT8MzXpN/Wr6fPc3B+JuFnhRrt
y3b3BUmC112OoFbHG1tesmV2UE1gNSB0IyBLGiCJ3wHQgRaY4Nrz67+cmJ9i6775
oFlVLXlQ7NYddOMG2EKWEgpqMGpTodbo0rmNIio53orAQ8tArqNlBhI6/chMYA0S
vop1pOzibX4ieHt5MtT8A3ohPJuemo9oG2/Q2PGoB7WNdwgpU8S+Hz9NxQvT9llC
wSsMcMmfteEUyvHYXTbk7qFFUpl9tURBiv5f/GYyveEiWp+L+vRv9rrijEiEGfdG
EdM+sRBkR1FuUMUH7e2p6vE39dCrOQsoUKZv62RnZUEAgMD7AfMZnq4X8XB0Y8wn
FVLE9jbxHMN0Kwtc7QMxiXiqNBBR2yoGTgGlsnWin21K/uQjcQY/yr57o6x9ePDG
D4av6pTddfoTqQM08xyTlVC3oQbAdnwagOPk4zDaK2gicYJC8K0h45C9avhInx7O
ZUVLoaRtMpNoVYdahxQVAodcUyvQKj99VeH1WZRjZ2y94/qrueojY5GVMF12Q87T
r9/m9QaAtV21CwAn7X+h7xzzwpSwFFyIhn8fYS6zy+S+h6IcC6wDuVwI1iJah/Kq
Tv7FwUqYmjtMMsTcDj3PjGULnwAoNnUL1sc8m57fDPdoqqWsvwoF3omkZE0olvjI
wZRkfQCStL+kVTO9eCRtMlBcA2ZL4XCEqZ+GFvr7V5vRuA00UpYpdXRpPfTfZbcm
f1ZkKVW13plWloc8fhLXJTtlW7LqGoZFK9QPKhg0fjsVNwa1/N6swmD69k7AGw6V
pDfttMxbHhSjp8skxigjgpxtbOrtEhrfWbhLdRDKrqirgRPVW5AbS+kPWueNDzXl
JY7k2FJKAt/LtMdy5pSeJvsB6bpU3KfdwNcwAwXVmXPCagADAkZe2H17OE18bONF
8csnHuqREPETSxM8EQFWOQMrlLoYWrS72+5g47YJx0BsukUi4b37GFOX5VT8aB0U
wnemdixAmWLwvO8qkN1uRm2qYpuKClIon0rr/FAO47f5vwwpWtVW95hOew+CaPAg
JvWxnIFJIQMmJUJRKiTvly9johw4u9SPThVPUcw7SqfkfKSpBXC+HqS7vQfFzl+K
Atd37/YDtTb3HuqiZQQRaUahAn/akAzmeOSQz4UiKabdZxNJrZoFhxM64m/KEbeg
cMDCh5PUCHSiz+P8+FyjIahirAy+wbSSgQox8f75j4ORgwSh3XbpboH536AM6UQj
cVFLXpFA2sAfhN7qBinRQUZmqsJRD6/+dHOO3Ml9uCnT2P4F+joRNTsRFb2znsoz
ovO76niWIxIMR6R6utntbY707IBM55QKuLwHTOj4SLjQ40Rj28+X9e7AhcBjIrPw
f/gy1esvrfrkV46R0B+QIWtuYRM59cdaRnOs+0WXHjAS9J6kSlJ6Jdp6JKFinLjb
9VcL9SI7CuWjEpWcvCD1aZwHaqaE4GGJAIHHI+eJy99P85SkrBbExo+RiNo6p3Pl
3X4KWRlgmxlb5KmJYpcGLAiPVdQ2yq4V9GXSGZW2f7AX4HN5Dr77tRr6mxP00aTr
oMSXHgFTVP4h4Zk8IVk+sSWvOioe0gEC5ahdHH9/o8luSBcdAaU79EmgaMDLu4SY
CrqI2pJ5wZoNVTrI8/Cj5HILIXdEpUaEW+4WjPk9GWPqucyY8pt8OKH7Dtwvk60I
E/1xJh0Ol+dQtgEmPNX5UqxAhm4T8YhiOl7huN7g45BOdxNmSwCYnK0sSe69SpPJ
O2gj/tYFVf2BksfB9e32DhJ7vSYDCC/xC7Lyesf6dGqPR4kzSgb2W9m/Va9txyRg
HPvQpvzjpURlOE+gSHL6z3t7GWbgj/IbUFKov9aOnzzDW9tbz0Jq1GQSnSOExDll
oObNpNoiObPj4mO1RjDpUfDnmmRZjiii2+ctQP1EKVDPryuQYm6mvHVlK+KNoQlX
yLGD2iwd4CER/Io7IGkCsaUEp1Bot3G8IAL1+dGyaVyeFhc+VaBm76MRfM4ubeoB
9yV85/M/hv5AE5AMyXDGvdLUb0VVOBMgf+isw69PusybFFvL31C1k+mQ1peOFcE/
D9JQ7sidza8CKi6Lw/flL19dv2NGkzqUQGXpTSrIAeV87biTtG/YruzCq07UByGf
9DnTDwUd2OYtYWPYkQiDrUeIE9XKpFt3VTm3fqZY7yBQcXpt6uFFFH127xEX7grl
hJfYtOAyPohBURShtL1XXGQvFtlTP9nPhf102RQH42xEkhhwE0YBpvI2oxmipNZV
Xje7yn/0iun3axOxrBBOPwK+/3U9UM4a7Ttbd0meqG19xUQnMnnFHmu2rKmMnWfS
LiYu3aFyCiM3F17CRJSJfDjQnUS1JCEejftryYfe+SpezUrJAQmjCHoXsfQcIKSn
OuqMJhjiyrRCx2fiEtpfS2apHAsrJPxGfuq8i4UOclhUE4sz0R+0yg4klKFd3Mbp
N1DQYs4Z8zNc7zas3ovv0nm9kLTbcj+J9wAs6B6sJU6BI6/sKSeXIocASSJnfZVG
31qO6OW0OmjqUowTxxAoCO4q647YmMDNAcXGHU/5AUb/H7tbNKLfHWDiS38KkdoL
kcVPQBHbrq4KMKHF9PF9vHGSWbxY9YOk0gxZKRhqX2RTNFToHFl8ojmUkLaGj1BQ
Y2bcfcuODOWQfR+XZOI3xERF8v0f9+UjCeSXY2hEfYuPRd0EKSyiYVTU2sT3pyo5
Gzcc/0fNk9fzsmvQKd2ZEJxpHZc+/bvBbbhD9PteWLNYgSvXOZ94pVHWjFic9VZl
LMnm/Vo5TAt8bjjMBy1t9IxnNu99Z0f6hfqi/TiwJn7p3rEHPudZIl8uNZDdOngM
A8M8uJEtm51d6m47xlFV03PDjn/RIwoDtQ33Ci9HXQ8YYn4Itd9j/xpAMaodtNqR
oqlIIK8aeNbQCFI0aJ2Ffwka8Bzwf8+Hx5HiNmOz5heusbwSNAcoXZ1RDxo/B6ov
/XT+enAUSzjdp8AnTFF6hTK313nUU+EBhv2DwC3e4VRJ+1pjcY4c9JQVuoL8YwWz
SzctMdRHjT0ai0m1jrZsSwOPza+dvEsN4tNBpLEjvOzfZxGNX8Rw0vKYxYGS6fTz
B9iBdbNeU+iGNgP0VvkI4rEaZtqTE3w4qK20SOnOwakl63v+n13dSF/Ydqeba3eV
8d11lbzBzf8V1MG96Dss12nJIhUjg4KEjvVOGOg/nlxF53WkEPRsR8/QCPqmhtlf
NEhFJzdbRb5wr8WGsoM/Ey8GLx0k/JYxRg9IThSZOVpJzoP4C/yTAEQOEC5bnbUu
ImicmFrLtU139vklLeAMfdovD5EVun9hXpYgNBnhMpYbd5ZT2zBzsaTtFkbxiHS6
Vf4Ujjes1wmipAvjVGlHqZw0WVJX3wzjPZYrdugQ/rYn08ZMfbyxs1WYT//w880n
kzbz4x9SKz3NPoecuW7AC7mhQPMcvb8DmQJX/OwCfOouxPa9q4Q17rtEl+Ziywu/
i6mtKTt+xXgA5UWmrJZflVMx2EGNEoqWzHjQdIQI6PLM6DZ+tcAbzEmW9CyqdAaC
QtErte7rFy+mrYms/q5GiVPAIAAceo6rw9DH3B0289ceFb3KJsAQh3b+TyNSbLfK
VT1LG2yRBPdulnfJONLWom02gv/YpS0v1F0nbYnh5LkXQlsB/awndARG2bKhjI8M
pejzaCkXEBDb8UohigkHIcbRMzCmAj8Vbo4ONfBiNFFVR0XMRFhGY6vIvSHZJNCx
ww+6oAjYWl04EGOdqROO9mv7Z7CJYg3++pqxTlDg3/oHaO2h3/wTyG2S3GzO+c0a
gHcTC9c8Xjyxf+gkfT0SzCUXEg9CvaM6GTpFHZxjwGaZbfIXdO9+A3sJ1nnhBR1K
N31fJ2TGmUsSjWwahQEXfEq0r00OfwZ7PEg2XkXbGN/QfWyrK8fOMxf/qaerlou5
5M6Ai7YOCu1qPS6DOicXhz6rIdySA6eKx5Jy+ZnrrZHlrfFHmXrfkAZwUAvQ6P7w
9FlrR3ROVenfNbAKkrLuslwxxlVzUYVvX0vdOLS1/tBRnlcjbU3cLzy6oTWJAwpG
NtUGD8mtp36+5GwKNG+j7680mxJnl4cCZskaadodtlG62UR4JyssU3W8EyM8bUZc
Zaf+EpHXUSW9UAVYI2xNIJNQMVYwHO5d/XTSFTjbnMuga+fvGs5HEIIEwAQhttso
JynwuZSXx8IhOpt7lkiWwhFRq5eGn6OZVd9vBH4VJPFWiF35O+QdqUuMfRMT1gYh
`protect END_PROTECTED
