`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kh79vBp5apE3kc8VGMTvJV2E37RzDjREQplV5DiWozsKqZk5udfQyTF+CqHZJ10z
ELq4bs1fK8DjhSvp2Pal07nU7j2ofGX7OKevCjZcfV4LmshvtuCAuuDIqSTA58Rf
ZH2c/0XvNiXtJh2jDJmXr32kVWg+7Xi2KSTCw2tE/lo5e3WObHrO34uKuZYVB9Ty
rNpFFmG2RaxV/RI1oLIJUXWSdGwiheBrQLGtAkglDOfR/i9AaGKrhCloTIBwpbr+
I3oaHUYou1UcCFiOobYlyMO7qnnGqRFPh8HCEZ9hMgfaFSuNWZejsnkLsNvmWCOI
yJ1g7TNyjZjLmf2eCCAct+keoiYTfkgsFPnAT0xbQUDfpO1pLS9yNU8Pu2MCCcF/
cx0A0G7L5q7GKq6OopQGHn+Neqg1r4V7yWxECD/fsZXn+D5qdl1O6zmKs4v1RSMv
Pa6WSVOURWJcyvCOFEu7TBGdpci1bF61HAbpqQdjfwpUE7g9jDTo7+eW1QxUH0b9
jq0+uuaAUv4mDirBoFHslEP5ubzc0CNH1x96k1qEXlmA4R2ejBrwfdMK93ypo367
7aDDuoR6juHEbHNNmp+IU7Wue63/kbSpZBEWuP0vmRXiwmPVYUXwHh+HJH/7uAxr
mpl84XH4AaeaIYSKjEuyJzk5YVkgp+/y8OEcjyT9JARkE+UTqFgVbS4B97ylH+18
m7eWCZLT7kXt/jytJsUM7N7k130EkE7nePugkwNq++7/uSs1tM/zDXW/7IIbTuKx
zBJ4ITtl/6YTuq2AmoXAB3L1yPy0//Reev8dqverm8b7m+O7GIkozjun0MIHdA0H
Rcmc9SJSqPYSX4ROhzBMARjz2AK1Q1jIEw7BT34+NCK17wUMIWat9mo9Ma1i/mtM
+A1W/a0Uo+6iOitPjEROYf7u9cyQE56KUrf80nyQI74GNxRxcZkqfMHh+uqdyBFp
/fiVt+22+4nJwfuIjEWHq8J4xdkgenFiaYmYXGcBGByhJ0ngfkH14oIAfnaazRgo
L4DuPQBTME5Pz+LBwTmFA5Y0UhkwtipeT8CrMszFmct+ZUy43uw47yo1Ve0sIll6
lW5QZfNEpZDttk8B3GggEjenjEZ5AbuzrbUfU1XxtKfqOt78HZgc5/DZcNFp+/uP
QGFaB45CxRUVmI6Rqv5ovRxbgvpOt6iNP7ASjdAFbAi6KeRDzKyzSDeoyq7GTWba
OUmwIsAq7ubi2zWBX9Q2FLQNGVw5Nw1UdenTL9vbhb3wTEcC04fSDVogwAO5yLcc
sWAz9ZyoWX2c2aHamSSOl7cOhCZ/KA1C9+psZKSCepREzcJuukapsdm0qGfXmdV9
uDdU1+lLK3/hd+kzNEMS3TPY0CgSzN1oXREwhr2ztUFPTeRKmbmDPsnu98mWauhY
DqlAYW7ggpokvItUTDTIRS6cfaGJ7mJUc9D8/CXqssojgZLNQYYk/soKRKMwhFBM
ihIerP2uLpm+JBG+KVlvliDBRdFxdJkNJqgMcAzQAmWjQQI9z4G5t8TYErP0SE3t
/k6h4ojHc2ZJVEzJC9YPvjI24rt1RV+iC1UEOqknnkHRuQrpZ6s8oMUVEjnYA6pm
zlauHAbQc6voMrG0zugRM+uSV5W66nN3XRFEif8fTY9u9x+OXvw+/QUmHW0DUoGr
xSGDzuQzujlcH30Hng5T3eBk9ZMGGEtlyDmQupWoadMo6NnygazCmVZCUy9uPKgQ
P07eL7H+0kLToQGOCDt8NTLn880eG0jyineO0ZFiWGDFZF3KWXHXJMJ91OlOcb9k
uDhsSdAF0GROJbWpLlyvUaSubCum4POyh9gEwnSuD2qYm4kKDB9Fsf1ENNIebPuN
ARbiaH3BPNdE4XNsO+XnjwowFuYLyYyK2cYTrUHeNguB5qbOBK9ofAPPdkhb+1a7
QmeAgoZkVhdOJqo6fpa/LcbfP5NA3MSTG9ZxPD3+kxANui2YjapQLhYM4rD/Eypd
zZw7NwVePcRyuj/o8xRXVatRv2a/D+ZjXwuSFwnUxPyQENTSTnNt76SYSj6uQsgF
5CpWlJjDTguFvEq2TKJEVxJXoMwUNTcXY82AVqDoKYuGbsLgqp9CIKO1Ag6dn4UN
LgRMM2sDnGwqjintmoRBXMrdsCVHxMWiQIoQn8no3zlDeZ6ptHKT4OaFtDp7CUrU
THHrkzF6Np5aXATvEamGXA5AyjR9a9+kZMQeLFyVe6uboj3NKUQkQfjg8iSmi3fV
Jj7AS+LT4qj4jrIWqYuH6eyCKuyy09EHy6uDrJfxq5Nv4LvdecN1Y2+iJMdnu4R0
ecdtglIAcGjF9jIQ45oKecempF4MhPNPYtN3I7Ws1yDfork5b+eeiQUKghLX4Yfu
H7DMwNIVo8rNMB/mAvPdqd1SYHN1EH9UHOkETKLdkZjUz2xlY3bRTW8wxJKSrY/Q
w5j6hRVdGXPw20AK7g/0T9hOE9grjXGjBCUyIbieH7zwcsnNLUkn/aXLXPiTjktm
9VnhoaOeeR56bvyKOwzOfWI8kVoyE+9x4nTXXAR+HTGsca+/wxIRN7iAO9yFAhGx
ozH+63NXSqgBEY2Le5mhkQUueTIYWomlscBqepOGikllc2umoazFTubToGVqy4vD
igFzf7xmo2I0xaK49MT5UAbgVBiDx+6SFTcdvDx+KfJ0ieba4To1yw8KG32U8N+X
23Kw+N9wPkJxrcPhghaUjXqJYjzrRym2N0TLGM42/GAhpNJIKpXYDfNgeqyAQVb+
CGT8Tq+dPvXlzElqvg+eLwdAFipZpf2bHP4Nt8Krhuc0W9aKy0qRpEgGBeBT9AdW
asNmj7n9WgysifrS2tzVldjpY76UA3RJLVQoNc1DFIVSC4CjWHh7lARi5CUT2s2D
yvwa3ehetgDeRSVtMzpg5MRvPDf7Ba0p86XTgrj0MUE9y7UVBYMdc4IoK5H/FruD
b7nt748iblqPGJmIcRyQyFv/YqSAcDgo+3FrYGpnPp8Q5cf+JrZTi0xo8ZYgKbR3
BNsYYdxMkkfsKk9uh0rfrK4rKV2ANKYeS+Z1Iy0msh8UWsAdr13PGDheaPBcQExl
Lsf5aXj5RZ3g3EaBsgsNtJ2s0xfcpm6XaC2G9N0L9z3g4PH5qcEzgOfabe4ZDy+I
3ixRiSzJkGkeZcMy1zKYF4G+kyQwl6xF4MoXCYRjgcZTXkBLVCOigDvKbMnIfdzk
4p3fZsqNFNFQ93KuaArIX9WlV+ebXV2BlBTCRrzeMDZ7gKQN3jiZ+r4vmXtE/sxy
8bvxLRVqiyGEn1ixQBG/nIYGv4Dk/sj0Xsi1LyVOwq45W9s2ewWztGoHiuKI7+Z2
TZkRClj5W9EiMeNRmKTFXO5dYzFhSIKACVUfWVWkY12SFvE7/xsDWgfVe1cIZWsz
ozpSpLpQPTkRdrsRIlUJR3NSiWIZHHlDiYZJDTLz1dn8muqLqGorGbqQeb2R/neO
h8BDxPT2Zkq+z5urvnLGujxczvu+aSDueLhyFKo/ouTulC/ljQSkEvpPiX0gmMjE
8pd3YiMjr8g7JUEb0ags6FyfrGPhRosRjZSZCkidNJ3dtSXZxSiUy5sd0cxzLFmC
op2wDErOIQM3GNjdgoJuwDThkvvtROfzSHSxEI53ape+doUVPzLFZSmxXpnqaH34
WEI911gaadXJu+UnWlQcbWhIPDy0XIty1O1P0tL3yWFZxbanaRIApVGMya3bv6AJ
oyA4SNflHtKJfAbj9PC4N2R6P4WV0tJ7sOAIRCmTqJEyC+VMxGjrCIONOYyZDOlj
hp70/Cbt01t0/KPW0DTBoBMotjhjjqO5wmAu86Rzsmt/Y7QONy7jE5Od639+lc8p
r8ni/13jjnqYJk873/LU2ug09aO/A6UA7qGQ4RzD/B3b2nXZw9IU7QvFUHOEbuAt
b4Obb9P0iOHsAIKt+4YtOmedoK6Giiv+LRo9jDX6rRai4vGDoAv/pc67JQe/tmf4
isnSQ2LPpH/7RtLEKkxKZtIzBNSrlcACUDuKPPW4yYte0bmlIbp2Xx5tUOszP1TE
XOCl6usJixUFE8JvpAEUzdxEa/clOA3guVgwBXmUKuU+Ipdf0oa5U6BSpXhiB92q
y9eLXskxDmcXz6zL7HtJpb1iCo9RMzkxZ4T6KRQLzJG0c7CjoBWnbvGrdRihFSxX
c9FIaJZ/DRIDqJfpckqXojFErL4QKlDLUyf7eCejcKpjASaz1EP54JlLW7pPC09w
NVCCT11RlJB85SAoEqSh4pS+TQDfTeJx301pEvlrAWZegvqk+0EgEoaCKWevJB0Z
NfA9IuR3Mmls51d0wjwWap7cmTBx7KwrIfJXHxNx791onGP1FRf4bJL67bV8xuzg
0NqBSfkydcQT2MIvYbevkx9Sm5s+s/SCJ4KyfvnK0i8hrttSWDEQ8Vk60dmrGayl
gSXJPVmDeZnl2grv2KsDDT703LFo+iGapYEjR6utDbRdhZxYUCNDaNK986Qla5Qm
O/W8qckqgj/WlGJp8ZKVV/ieqFomK++liOV3cL+CGtzgS/Yv1l6wVDiPeEzTS9Su
C884IKyEF0bgfmYAzQ66VTvL7TrUrlYr5J8rU/1WA7Kr8P4kCpgdVcJuCNLE+30t
o0HZBZmluaCHHydAiIlZhz2rv56Gek2xq+72Ciuh1snUjEe8n+OjpXSx+vEHx922
LG0lAiBtfC6/52mvSlQevO3xZNYEyAwSZqQQDRG9eGefPoRBtpBAAWhHHsY1w7Ac
o0tNbVGrBnq0by6nThHpRUxA+CQu+cJCpzf12Ogdkmk48YQUCBh7eoDkCuhOpEzg
9u/Uwe88B0c9bRtEMDBGsSVelt47GdaJ0Wz73rial1KnOO9lIqHIXjzwy1ob4G0v
uCrzOJi/DY/E50PF41xRsTMMlqIo4J4YhFNlVt5ZqYpCSDk1BQwk+T5Z1vPuElau
k653s7eHmuoMUL48i48m/EJkrtVH+eprG7uLMHhQrFQy+uEk9felBx1nl6jDO7Qd
MlbvMgRNYO+Z5O/A2+OQ/+wKZCUhR2VpiIHIWKAncL4XSJj2lKedSs5pVlA9i3Wz
/RN3BzsWhhswJiflDQa6nnROxkBgS+QMcucCrXFD4jJvlWN1FNL3PyoIyU7DTMhf
XhajoE30iAaZuKRUz/M1SeCBIKi3LPzqUXvMpZgjVJP0P4gp/0rG5gM1MzWtF5eS
Ysmpq/i465+08Or3CMmb+0jn7KXkwoVLLJtrOFyCzKUANYN61ZG9uJ2dYgaKSubp
mL3a6/qP29bKQUIhYBw2vOBv1sZ1Q5c7S/jv3JIGjyIUH65fMAqckhvQ5KMuc2Ce
vOFoGc+2oMqhwnHZGrqQGOrcZXOHUl9Vi9RK48hjfRGDi4OVYzKRd9VaBpmFWOKt
9R+vchr7vZNVlQ6YElH5DPD/3Pfj6wMEZtKzoUcev6l13xakP6De34YCkgPZ95hg
nopsRGINrNZARtPVLSI+mZiojeiQcc6fA2PhdR0q8oVEz8rBsvfsNVCYprAWEo5B
N9YSyzV69xOZWOF4osoebDxeE+Sc+GR7MV5VdtpWbqKUdEYikSJUjZB1H+YXastL
ONIACFaAEttoelDQkfJVVKJbwgjeDhBLbGey5vevOMaf/cRmM+k0gtoIj+Lwhiv/
32jssIGp9gdlJorsk7b7gi7ULozAeaeQuQnfqlWRsArurM+mqmNmEMfU/y18Pq/5
yG3Pv+AVoZNdC8WsMDLnHAsT9UYntc9EiB9m0F0gtgsvrNnfFteANX/iUW+pETYa
YW4gkWmTSGFeRUDY9PZvzsCsvAy73T/5Kdxbf4x4L9rgN80kSBjjQN9ffL1j6rx3
3nWxZzE/jV9GjCVKhpMsnS38PlIIu/8/qV6/Z5uCVlLFsqBt734JFzGzg5PHEW4p
lpMbVtlmHPJg+bcMr2c81V0EQzEKUPCw/ABCtQklgjF4KGA6WoVQSnZmYJ8K4aF3
cY6T1TbTXB1p6fj5G4esPv2eR3dI6b9A9d57Q6B3SBP0vMXkK8lOhpKE40mM52WA
9iykfIyMCzGmkdFZlymTiiww0RfsYyqHVCqBuLBps9cV9ZfueE3i/WuWZjVhVJjB
cbouqJWYVatEaLgpdlxB/L+vhfRIcfIg/avD8B90CfF2J75R08sVoOb19fQI4BAw
YnIyXQmFveaSQGfCxHkasUinpF3w9CNVFmBwbSuQqzFpHp2hBik5o5DNnX/SrCM5
hKpH52VqrrrO1HeMpzry1Ak5pS8lvNzVMpB9BLlLRtY25cawkPaWV8CTImxH+8ic
xq2Wi27VPIZimShqQrY5HiRkQvWUnrfQ7Y1aIVV87vlE7q4s8RNAq4SWa3JISGa+
wLnCek576DWVNi5QJ9vMXjVIyOJKSbMqRhNBb18dbtDvVwd5oDd2Ths1p831AFmE
8XvOeQFsQeowZMyR0ain/RLnsa1wvNkJHAJ+6sG297gm6PLwdh6yXutUqj3SX5gd
guklIPgiET2k8UwUYp+7CzzDHI5FlT/Oa/GQEHLHadbAQTSCVIbZ8CQG5BiloCxV
Nuox33Eg0iu7pST9Hx93rvF6xCoBhtiGdhUbE4PY/qXv/C4CLWOt2b7H2otrgdcT
0w/+hKzXQ+5914eYShuDance/qUJQpOVIMmT0JRJHvfYsXEvDWfiWk7iYLgvhqob
AaY/DR9077Wx40h7yewtw8yfjc4Xhi7Cg15Na+IzpDU9pyk57pm5XL7Qlnkw8b46
vaC7uHs2jXv5geyy2X3o4+WoUMZZk1pllNMNlD2ULVtfnCBspQDlpQUSxIWFAqnP
8FhbWxqZFdsLIUOVeH2hP7IQwuoWW3/cfG+nVWfwNDbnl16tqMa6ftKnrfK2G9BH
AMkW5YEyalQKLqF9gMKgZ65kdb+98ZLKHALzesAu75fFvs6d7XsWXjWvqrNYNRBb
EJfNw9q9XJ66TZzRhrEU/T/OtiSFttdjRMVzn11eeWA3jYATFCKxkwmieGoO/O9B
ZaHp87pu0h2Qj9pySGVuno3qmKy9GkAK3hySJk3ZVjdUYzn7T2aLquCIRV9O1E2Y
zDGH+pQM+GgwxKSjXbAurk0dhpQLNkE+ii56OgBamb1rX+illdMDV5PNlfzhkMp0
7LPWgI/zoomUINEjxH6OcevwwufoLeZUo6TVP8y9QzX9lzFqBs/0iCMLRIE/u93Z
LyNHzhPK/hAjTj5zJneZWMhkQpuvcrcgnI6AtliKyUXBhO8ks5C7o2/NGeYEvMSx
EZjTLV3Q5j02vsfCm0DJrBaAb9LHbfVWXwcATsojZGzWC8GpYYegAo3/2/uZ9I8T
K2fWxvh3h24Dd2O1OxGFVGPXKe3uBeSAPejTaWEtx0Dns+F7dlPUuoPjGKQBJ7AG
cFA+oXTVC6VTXiRjEsa7v+Vja8msSZlXtAB0Nig8xH2GX6gGuEJlHSfOiJpXOjYB
F5sv6pVZSeQvq7/eEwGMwCCcBuDEBfLpm1OpNF0XSUalsW+GCT5WjpSZRwWCwJBW
98i1xNJJ2t4CivBrMERCoDCf3CeCoNS5jd77sBuEBmVsFshc2YrwkhvoJTUbxdd5
C62OfZvu4LkuTFwcmhdj4KBHOYNgtXJOPUcFoZCDIA1Ia3XWQ9SPrLcZUS3TwVOz
UCioh1Z4iv/hLbn9EUuy7rikJfamoe9+8nxMNNRxEL6mTa/XGgUV5GUm/rjhysTd
Nd1Gjjz0fRSck2+POUhAHmw9Fjurej3VTr/cofQcCAnW20Y2ueHgS/pYenPMQfBM
uNuuWTN56Ijtm2H2tKLUr4CGVX4rtEl0qYRSEcNRopL2GkVcFP0dt+pMDlQMgx62
G58KNB3DmUwq1bD2I6/Hto8K5ZakFNVPbDqcoahhrDr+gmlBN/JQ2VHK37lxEsDN
9Di8q0AqRMrPATgAB1O1T08x0EOtEsGf8HptJQWlEDDGtfl1lGc1xk3a9efYIjNz
9E0OrK+zG+uJrkxGGRnupByrsqDKYmKDeAYhN6Rrza0Bpjxb9SwWqfacFbmGgCNa
rSX6vuESv6JM5+NbAMFL3gbOO6AeDaQ0Ds1oy18XTJQTIKaUysCrJwHTqIRVOZu4
ISLbEqjX1Xu8Cc9YBEKnhwBsJvHFQjYcSw67GVs3NMZgxj63FxyIfOJRJtQEp6AC
4Pu/mZVXxsFRMBqjbfOwMYsWSapiYu8/E3HRMtIS4FmOJ0zs+4AtNfRi6O1dDGZJ
V+obmbwuOa7L0WBYOxY2t5M2935LQBZDFLwWBB5UOls2TYSpRro1n6j53tmGbmA/
5ZexgGaJ9+rDzEP64ZSFyROrpi2A7d0inBqP3K9QYegBYRLV8ogHkjKh7vPQxsqC
RUYXi4sCbubzUQi8eL6z/YTgze+qMew9bZPBCBmC5gFWTPEN92UaBwhJbw8R9VOL
Jd78OSxzJWUViPOSZedGAGEXujuLymx4NFgO7u9kDlWrFhbg6X0pZBG4vCqVhb+C
TvjgfW2/Hw2AIngDFskwgFVbOfTxxySWWo2DH7pyef52ZNSAoC5mHpOxvXBjv4RO
oU+7qg8HR1fwEU6hdbP3V3VWJGEOR6cO4dt8H2D6B2NiV5ilRA+FSzMYTYDYCy/d
V8ebzBZyjGS2dqyMc7Umr80esPGjalO3wa8HOOiwuNS8GlNf6gk9IyonWr0dSEgm
54PLwZAPHGHG/EQOjRlQ/UeHF555ml7w9pZM4WkK1gEzDeK9yPPIcdbnkGCy4+sY
5eQvU+znf7QkqT66BN5npudjBsODXaSS7Bl4GxKmsU7rRLNjDGMhInkIuDOl8nHY
SSPFBCuvp77FIPN6vD+tBK18O/AStFuj5jLha6OjNdH0QCaAYUvnFgCTGbEywZFh
67dYt2EaOMYUgiUcp+9bI8HtmDku9XtzDExWAj9BueC9pBYwt77iWW/M6P4lbrgI
LcxOSYsF0bFGv1c/2+uqX7nIxyz9cfNrIGdZml3kkTKlZXHmuMjtyFgwiqQQZJAk
v1ewaolrBgWXWeccVUy9c02+GlJbO+N+JdQ5lFG1Q6UFS4I4q6gi58Jv9SFU8edb
kD+CKvVvjOY1vEeLLmnqI8XOtmd69ZLz8FB6wuXCQ9SoMhHo5ysIOhDUYKKTkYpq
vozXhTgeBpjYJAwHfQkdZaV0xQcg3K4xs5Qn/huByysVzGQsBc4UsRZeFYvqfV5F
i0ywJLVDI/9w0rANYnRD9AfWRRImNgnoum+eAzPK2uG+TstPVCr5mxG93rcJ+BZl
fhr3c7ynIQtRy01BepbNciEqE5gIr9rsqELnJzwJF1nbbtubxjle66XvwAQgtUOV
Z1ptapmNGMKUUhPyiWnPV7/NTV3r+MuIht23f4PriTf1D6A5yLI7kSFIaQAOhi19
nczvGeDV1bxrWfvfFegUlulabe5x78fYkJtt+bdfUE2T7sldBj5tix1qM8YMB+W3
yY65wRHLxm41vlxGySRW6Zl9mrDjvW5Ey0JEXiVCdAAyt4mCx1ntrCIIu9m7ZOjW
LJDRdjwwBhZWLg/FMmHc5JgrIF1WPXCG4bCUfPg5wrqTTU79E31IGjjFrHeik1Pj
Q7YP0VNaALjHewyFlFqXqK0g5MvmOAmZfwqSvjTN4xR2fClh4VzpbheWdbqrs8lf
m7pthfBPV2jKqA2CK52mXHqYtK6AasATHnvJoeAUcut27uLoFmzHWxr74thV+sxC
vxZEGuktjh+oXpmpkMCx5c3rqbUOwvl7GNsXpRXUo7av6nGM7CpHnxk3HQm01qYe
VSkJKx0JkZuLDAXusll8IKp3Cg3f/LiQ5PWel9QXVK5yADpmiEM4rr5rQuE+pGga
4krfcj07UqUbz0oeWRpqbrCrjCoV30p5THkCJ1TdELlBuZioifG8hgwG6BL6gQaB
fpTnZnYpg/8g9p6+wvH+sI4/iR1joeRw88pbmZA+sVL5pKhPj/JhT/fUNoVXsiYS
nfumbr/ghdr/yZJacWfqrxp5s+yD5IbTZI/oBoQ7FXCUmIBp3yvltLxWkqahptdy
+cou6c2eS3Sxn1DUXbzwJlkWgu4NRZWXB7q6tCTQ+3io+FjJz5yueMtgMkRrR6fz
NWKiBwSfOQYWkp2FnrN6nYy1KjKSsCHhmzJWUW0OZHY3P8GdH4VhIrMVxl/mD0f8
jjx4iaK2tI2Ih3XzpNKgk7cuEzixYo3gvO0Og3YpSFMvjEbCEENZovA3VXtI4xBf
c1eEc0bYBIzwpXpHVMN5yGchowCPALIauEf9MaL+CdJvEB2ycQS1cVaquh3XautI
hdyDDGDPUMQCIoarx3/kczvhO6tDm05oTtaEX7PhiQfXtTo8UeA0pBA8NpjKeM4J
SIxFZ51waLBghlNQEIhDeOPwa4zy8W8Cauf/KbNOoOorXHqExJz1QJm4PoOrrVOX
yHv07ub9LVOlgWhADm9+h82/3kePkxD55zxxrIWYRsAMLcYIlWxPOr38c3usa+wO
lYhprtV+EXvPFFC445QDSjVWBD5ZANd0SsuGDsqHjVhITQWB3YDGFBDmPp2iy6zl
r98xv7BJwXCuglkla61J2qx32WN1ZuXPsV7Piq7e/HnqvqxmtUXY66AC3Ta2Daok
oIvBmr7uTT2rGG1qIo9pFT2eBHYq2xWAL7I0iIxckGJywaUt7KtNJKtqnWZRqDCZ
yPSoTrVOYXWfoBJ1wsPeQQbseFVMTD741qgzU5T1ay45NovgXwd2g2lQmUBFJPZD
ZNoMndW/Xlqp338iLu6o3ddiMcMGhfHOBjpJINMRl5VyKuhEvETxxOLSwXEnZYgp
OlFyxk6tuSCFRGZt5WPnrH5MxqTjwJOmc26Xxa9Q3MBgE2eNWiG94bk7lQHCSK0l
W+Jpm6YpUOzSoEYGjukg7cU8Gr+1W82bPD0Ja6gyfACL8h0j8Fmtiw4vQEriKeXY
+goz0k98X0dzxNHkHwo3inIROim8Tz3iwhIxIEmF5e9q91uJNc37rixDa8+VhQbV
kWsjH/JxILcD8DmXFZplMzReooZNZD9sirsJf0uTQbVzGpGC4i1k7f+ICpCu6Zt/
e/ft+gaS7SP7DJJeUmGa8G/9EFpubgM/2AB1/RYQIJMN/owN9ZubYimvNJ78qOD2
YoKPlJKc/Grl90CpeBtDm2RWYNSliUpQzeqk+48nGCK2Xy+Nm+aXHghaQ33LjX4b
rTGJ0QsbHX3o1mUINJNnll35liQatBvXiIagyi/RenhnsMbF2AlNWfXDAFnqc8l2
g5oKw1wqXQ2pnFMciJx+Tu5kG5C9Qz8Cwn7eQLsSh8/SCzNjtdn9bwdsdkivX4OX
M2efH967BJyrN2Mz8AIbOO4w1R/ZFNgT2xMcUuwulGkHFI2yfsTYHOt+TnIGjdnr
TWdFus/msDxq5Cw868lILld9t2VLLc6t2sDMLBLaGi9CdwH7ziF+Zde8Uhe955Fa
YU6UrOrHY0oUOfNMWr4o22z/PItvOM+d45c4SPw5s/NWBKceYLdivg8H+r83sdNt
xQ9mdkKdmjo72r4qTocw3xq3XLiNC54U+6uDYdr+WAftCQTxpgaNVeFm6u8YEntn
1wjaDVR9Mslb8RzZX/Sm53tnmMMGXZmeNuP9rL3WOSLtsevXOYL+NZFrtY9AVOXu
llVWDPB5FcHuUEN7v7F57O+XeNwxna9fc/3F8eCvmxznyyix9D61BK5sL97vJzwS
d+ON/28VgrjA0q77Zjd57Xh+UMBkGzwqjNPYy000gCn/29P9hDZg9A6SFCpgiysi
7SyPb1HrRuIfVJ/xII/VZ6lLz0ALelUPo2xaBAbAvjiGv2rXDbj6dOCeAtcuDY3W
pX/76WXfNkx8MVHIObj/RmYgTC8NdyBzx9fc5LZ/fXN7Zr9l72oAjXR4QwdXbU+D
jrmKReeFHPXz7rL85WpS9vDNRbv2Y2jCk7796NEWldEEKnRLpqWGkDfN8gKENcjY
OHFAHU0D4EhX7cLK7n3XVEgks6jezvsbVXX3zGkt1WHC1XHXqMHPyzzsSs9oMJTL
M2ilq7JPcA4y9Zkw0T6fsACYR6Mx6aZ3Fo400f8+y0JgkG9or5kGJik7uDgtedDt
jPmysS2iFldMEvtEc838UijL02cFbjOWysTX2Q/kJRWzzNrkEC8ZllMcIZsdco1O
ySIT924FrBZEe9sPI16WpmRaNfPWDknsRyStyUqBvIbmWmo3I1hagYxkDXl640Qi
6EEnYvXog+O+jllMkXYhH7s3bLG/EeW86OF2kpfwGGRPzLNL3Qc8RxHpnDh3HdXL
CiJ3ahbxW5KV4e9DFzmImRxB06ilrx8zHdiDKr4idIOFTfioB3ztBh/NQMWjCDur
SiuAkxpOznx4UjQF/QyQ4Bw2mAAoLDKE2wBs875P+gKJwFKRp6OeN7SPXxwG6icz
ueyN40qqiDh+I0jSoE9WORZ8LPpB80mSA5st9tGg7C4Z+UCxHUIE3bvrOmQU1tw3
tNG2GuS0LzMZBgX72s+vmSIpCUvCiOvFy0m55nE5MNrFB0M3EAlwR8xlSAQF99Ow
ezLFB3p8JlnI4niSELDYHDu9BQj0dFex/JibD/BPh1NmJvPvv3H3rNvB3h9aR/co
ILX2n/N/fxnavOcXA9/8ZlHJ63Mx7A/seu8OKeIKKLejYHQs5nxAkVOcnmBc5msg
pipYWvpobtgEKsuD897fmGAu34EjByB5iTOs+VAec6+ZEbW1mlV3LGJAaNX/bLa5
69pe2giqnhThdUojM8VgwYKYN9P0gJlBF1i4f1tq1/gD9gY8lnGLpDcxu8EXV4Cg
r1r+eqAaiHd7cnAVJpEarsNfjOpSon6Z+7wZLlcUQeuBEWdqX/htIfHol7MFKWMH
BnX9zPk8//N89ZY8R7IGOgGrkN/c2dxww98gPe4FQ1/xNAe+Si7LAO9QG0zBqoiz
1WkBAN7Aujc6g5k5I4piWmnqTxAfgiXkCWJYRTNGMvG+rOQ7Rne4v32bM5juSbHo
dPKQx1GXUP+87nixz3MQDmFjiwqeEbvcpHUGQORlJRo5AJswVQfKIullUOw3pgBC
KCvByRTF5GpyTxQUq9zyfz0e5OzUjDRzNPsLs85lwfxHB9kfHKYPOiFuYKMyGz96
T2coiLOPZZtR3/uN8whW+wufHbIhA736J3Yj4SDJ/IvJ9Wmuv+hLw+uEp1OdxjJi
do4HNxb859J0X9b2t9+cfHEG1f5JWC/LKHlWhsduht3P8WsuuIBaX458I10sCQFI
kxx6R8XB9apwTEsRfM18B/PWcup4yvGt7PXMfbKMjEZxf1zdccUduEH6rtICC5Va
8s+9CAHOPVcIFnahielT4CKD2FBjpuapG49HZWgqLmxrv/+yGXjFBfn9fjllh/tb
/0ix9UvOC8qlu6D0u81i/wG5sgUE888O8TA5YwjC8VkKfvo7D9BG9stlhWefMZ6a
DKYIDvkskt88DV9U+hVtn7DUpVIfsxGujwVgKDkXs9NIrmtTB+OCzmKoYruHYL7S
eCru2+cLuWxV8glRc1LR7sdrZJ7F+N//mlmzgWOAwG/YkfBh4HWCFWSV8ttOGj3A
miZT139r4NC3yVfmB9JwKgULIOzIs+dCdP4WJuIZf0K+nD7wHLkYktAQ5Ob2rObY
LHMZZj2qmzVoJ0KKMwJhB+VwdHtg0YSiRjviP5ocnEaklUFOExT6nKqpA6kbo4PQ
1PV8rp2zeKvi+/ZsxxGmjFd7p6cqoIJ/UPEihHAsv2EUybUNAIrRt6mIamvMqEuA
TAyixmyZFA1yqYCM45IQ2rQHlEx4xzieqkAYcZORGfX96ZVatF3oB+aOAovwugAy
WRNxkgk9pZoidcTwjH4eio5shezOYppSGy1vHcUAN5FTgCdME5ce331Fpem4qdu2
e4Jdqy0XKNyroB5Fk+kCQo6Z/NXVI8e2XZ2kcQtDwpiXkC4lBzyZ8lKSV5vW5YMe
s+o5C8CcQpnC1Ie3zlmZHGuB0c7jgCWyU+KpKVl/rH546Z7l3quA3Wn8RVPUuGw5
WobKos3FgBUH505FUzJWY9X9XKrtm1zKiB0w3sxx35q2Q0kSa09fVQVoc8hmuBKr
LuRetdlRQshfloETThIPR6WZy81GGjM9IVWQbYX6mz/rGWINdJaBZSHYlHkyT0jG
Qhtl+QiTu590JnalZvrarIFmAPeRUbfzubZDYzOtaGduNX36239U1yKSDz29E0VM
v7xsWcs8pf0Uo68lJP0punvJcfDqValGMh4S4dBWlpT5HSqJCrqDtpEf33bsBgNz
LNPk0pL6m6P4N5vhNw8KKRRNPy8Q68FOAjiaBPaS6ZHsuGeE5xTFmKoIm1X948uz
osNPKvWrqX3+lc9TwffZmSGHsz6nezydVGhUHWNquHga9FjQh2DdFYAjgC21H9Le
Wphcx2Il6UZJ2f5f/t09w73u23Fr9sxETr2GS+brXHQSX61wKAJcmIFoN+qYxE+R
y/t7NqzIwi99+rHpVrpW0GgfTJIf1Tq8HmW4o90ICd2+PhJ38cq0YE7EFiGvFlp9
NVhkjSNdAErB3rcAHarT0yjLuLDKhSy630Kd5YTKSJlYlc4mYHZycOQYLDHc8XM2
ptsI/RfVXHPlXGYrVlCrAlWLVapoyIho4MxNKrW1VYPadIjXCHNZn2KjVe3TwDUK
tzoVgR3XGCkOUAJUj0JKauEzFYtMTi70i/hbRYD5vom/txPQtRgLRDlgwgCg6IAX
CoFadrqm4xLfyEf7T7p9YsMWzudne4kVTin+oVk6fJwvNjWR2zBUvLfNtdqxOF7V
dhCwmEKQgsjI6H8Dr9o1Eug57ClU0HKXjoDKI8ZVQvdgPOyPU+J84UGC7YDV1zq2
Zz9ku+02LIJR7cEwkW7bUYEWMpGh+BGx22c3OJCXgMpkb1iBttOuVlOvNH20j3JT
b6PafurpzuzTGnvQ63eUHN2e97ot+tjCghGikouORL+lVY/nMik6aVVavs2r6x1x
eZKU08F/c4ZD4AMLfIxPnHf5T+/DzF1ICJiTxWAuSMhGpWt8ycNjJKW4Oc3k7fGa
KM8eUasmaCb6exmb48+C8HYYaCbfj7AS03jdpqgua1lUpdRkplRxIAy7QWDMbXuD
CVsZtfsU/Hl7ZmMXV4h8NVVsSHQfchRUc1iwQRO1xecjLDJk6po/bQ0nks16bONq
bWUIfBV0ivYXiIWRcjfvq0co3gr9It/K7odNtVTaI+z9vjzzcEwIzeWrJnS3fD5n
4Z7dW5x5ecFLxJIDs6cyTRV0mSDGfek2Be1poi+3hOSz38hk+ucnahwsDoRy4xbn
ySl/YVTJ8X1mHTWkKlS63LkhRmvVyfKRRC6STDQsvTa+2UsWX/K0qPf8pDT48r5o
rp4MoHZWZJHHdTEijJwycdYUU9dbPB5KgzIGoVTyPwEekt2c30XO0jda+X4U/b3R
1hW+4KRE8UTIBk4HWT1YXEdMxvUB+KhFHu4tCpWqPy5xwwbKZ8Ln1dhuc5gub2Sw
ZMyuKWSwcJC/qzVmCK0jkJOmWv++GUV+qaNLAzfTbutf9lJEo9/Gr84VT55AIMBu
QSuPCHdrrB9j5n1y0LdTCHtQ1kdgWPWeYce0KBNmBKOTmFSTpbiPYmGkqosTXt3N
Og9g9aV85Iv6io2iTry0YsWjH/aFuoMChpJ/vqSyXUdo3E3gisS9TzwSrvpCiwq9
27PLGxrYcLsXeofv4pkbypjalmDtaRklzFa6yw0i3bdU/4rhkz9fRwTLoGLJGqYf
BnZKBmHAPnEKSK2VmH7Ug4MS3NsFKQk93x4QlXlGsCtd5Xv5P/8fGTZ0LRIlwrEl
UjnhxuHG4A8r7yZgrxr67gNxDGFpp+THca0HPQOH0OLJm3bqIv1Fpft8hhTTKdBk
AwTLgdStBqgK2HNtGIuKDRmvqR03SwsZjDoeogZ3p2qaF5HOgVsBT4uUssvYMcro
E/N/LTBpomsxnOshZ59feKo+9RUq0K9JFjkPoOkOwjnxgyxYr3irn9jOk2ygiKXb
TUHYTx4LNX0IK594zptER7IuEpTn4pMQ80LV0EsqPi2fPffnIerPR/+HsmnEXR4U
1pn1Y/jHtSdqTsSaVtefGIaGS6aUaT99AkJOGJ+wfGZLssLoioFb5DYdrr1hnEdV
hmf4XrlRqq/tV9xnTK7ZRVFbE4WcCxOEyYIfAxYcLbo//N7BBpbc9QHXNM2klyvw
LdkHiZa2pHMiFyPdO9XDhMlIPd6I5D1u01VR+qlhVdaIQbBqRoBThNtAAHkFFxCX
GWFa9C8DNBhhDKqgIWeZftc6FSKQrPhpjLUblsbsie65/FI0JNJ3rIqgMq1x9U/q
4Lxmj9IE/OiuQkXe29vI172sQTioWw72odrkI0Qn6rtLzkD+XLeYtLn17m/5uS0d
dajAvKaoAUwgDqT0MkV3il994fHl03O0+Vzps10gsIPSXvoPypJ63aPNg/6pJkaF
CaCioYVMWkm0Q+PFvu8wU//VTSves1velXdTs005+ywttBFz2JHhFNm4PNOPc8qO
Ogr46LpbutJczsvguOevmMnqgeKDo/OIm8mbdBjTWMCix2JeWuKi8F6gQxz7Bgby
5XOIS6VlPSRJUm6z1LEFBTpvw1BHfoVdym+Ow//oxTVA2if16iO7/i3+EyPVosrp
vOPNsHeyQCWCFVhermu+xiYYKgTfECvUcF1R6t1rIt+vMQRoKmNpjb6XApoY/FkI
QN5xNUBBQGMn+d4PN0eNmPhQOKiM722fBWxY3/ggId7fLe818ina09mbnnVmvvE1
EG9uHg5skmxBtHuvkpTmMcb7+9vPKgcxbZAYm4t84KK+8mkKJJ1l1BYgXXbP43Ib
9yxI5PdtP/mw3a2OZJqGH2TJW2WYOn+8olPuyBYaCXqmLcDjAyyjFMG0A7pyF61q
zuY7bw1nooPxPiOmKDDh3piPJKxP9vkSbGZw1ePRidaKGnYY3eba+RY1mthHTrDb
IZMB1sBzO4+aoUWidqEMt+gtknEd1msQGurE8N2Ei+Yw+0mUmfTw4qJACGulOGG5
jONv2LJ+iRzphVLuv8cezx3bX1SbCvhyfRdGIl/jVYV60/Zux25jydlWERf0OkyB
hMmbN49v3TXbWrfabxPmEqoTwAo62mHYSEU3hblK1KyI2drsyjis6oR29BncQZRu
RhO5yMBpBS5K/K3qsIzD7PAAPaILEcEjmeshI/5AJD562+GL/ZPcJpJKXTuKExqz
Cn0ivu1YPmquuRnz/K/U6mVNvcsA16wtfI0bcTSnEPVJcVqKk/RFd8f0bOJf6mjZ
ZpaMVe62xbAtvV/CS7UPVE7/Y95kkP6ahWW26pQrt6x+3wl1Ib9YTV9K5ijuzZJh
awt31nPHQvF2KEYZi0Yw31x0+vqcGMkr4bG7nRG89SgWxYuQXCi08oTget/JTL1O
6plZ8x8URby+rLHoiLk268B36dXFU6zmk27e5X/R5AGhHn+7b2ahIIy5jIOt1L88
behvW31U1q38b3OR668qx/1LmcZoXX6oB2WdaROMgSG6Cyjycsyw847nkS4wNuWt
w9dpgZZxQqpApCE8mMuyggXsMyYyAQ/jDoE22wfcf8HalrYZTbuz4ZlPCPsjNN1r
l7Ej+DRazvG3HFoHbAXWbApFi1h8wkCwmr0fMLo/vn/qGzPotnIvud2l/6QK2JSo
UXHMS2F5kWtVq8uRjg5TjGcwNClOwKFMuypHakDxbgdiLu+TIQlAM6fbmTMgNEmi
nlKCjL1zBaLca4wAb88me6vuQ7WcKxAr9Qcq3+u6y/I1Ym0tvS7CG82+Mi+KJMeg
NWZHkCtMZ6m+hZWrDTXRaUdqYNKZBtmSSQqWcUAWiosOT4WuG9LOjZN8LL+eQ6yo
N2cu/FKh3AQ6zRYoSrAhdtOPWs+DrY45f8PQ6wf9GvUR1S4/t0HRPraHem8Gn9aS
abwEObOe9ZA/H3IxslR+FGWyVyygb1DaUgd8IAlJ6n6QaK19tpjkUC0tUsY8SPCR
n2XndT0RecLvwMdo64Zvm2/s2rk8uHelA5RDI8/jwSGpHQJOcrAOk3+/vyul7ZWL
XUIbZnTMvTd7pIkKyiq9ZiZQUU2COjfPlAZfoIltbMhO8LIDsbjukdOO8LJ7fRzU
502sSD5Pt/Rgp+/SSw381ioQmtzlO7qBgsxfRFy9eL3vl7VpeQVvS0WNLcE7rOGP
W9tk2+gOOb1gk+9Y78MjXrlPlck4rVB2j71MW9Xrbx0Da8znTZIk8Vmp1WruMW8L
PzmX09uiVdJQsVyTk6ysbqVFKVFYhz8NCYcLJVAE0HLSyu7RUaltajCY5GBd5kG2
4EeywXe3thvjaHagGFH9UGykiI45JXu7U9pNDbZ+BYl1IoR2fSPequjPnUcwMKl3
gdqB04ZvBM85uSej6trA6FUpHbWgWvmVGNSJVyp827KkInmdYsP4z6eOD9ftNI9o
7pZc//8+TrFg7dLbh/V05hfpB3DD0kYxRcSWAlDYWYKVaSQcrL3adQAu84c0OkSZ
3OL12hvWZQoDiwiyfFEi6hHXdUge1SzQcU4MeJcqtB4eUbt8J3BumQodEWBd9x2V
fLL/9sYq8JCubuPZv9RlCoybiYztaYOcX0ccQGDn5FwQ/wrrsb+QQyFhd96McbxD
YYkREDwDURXitcJLEhHD0rkcB/UIHe4PJ6KoM+sH+VQTGmCz0aRVz9STl2EHVpxf
A/pYLEUppW39t04t9CU/jHbPqzwbX34+X8oLZ7XrmPMhDsCddUZcvcKPiS6rl97H
Z7W2HhECI/bCglZs6065I8kNpYIsmSpdgfk+9+yo0NO6cqrgxYE3vuTIHupmBZbh
wlPDgd6fDFdbazhVyOCsvQmEfvqxlMz8+o6yf9hMZ+v7UWxkcPPm1sFVc24jgcrL
0N85yjLnOwjkkaLMlKy0SykTkZNHWVQjuAsOESQ5QTQWl5BLDcgud3jmY0KOdkEa
NufDxOzO0JoplPi8ed3kEjqohXMZ6jqkWyTR6ZbvdiOGG1U0AqZNZFQ+tr09FAwA
XiyaFWB65dWtxHzEjCeYpSpfOvOWvoHFus9Pr9fQwIk6O9itQQ49juTRsgjqilMq
6PZVvSPV2GfcQYOPMxT9eor0rRDlguhtuyivm418oAms5DQkz41xb/MUAoBLbp/6
MocLUbFMzKKP/KTGO61X0Pd0LpEWQ5YzfkkvZLvhv3HpLW7ueloH5mTkpj7+nUGt
NGzON75LbeYlgeT8CzKgUlAZ7C7sKY2CLIYaDcct1iIuoJsBPN4EfnGbb0ofDCAY
Ut78Q4mxzIQFdBAgH7AkiPPqmiykdM3C8XhjSSHGZlMAdGIJlG1I3kTP2W4YmQ4z
8Z6f7sEkID+FHDRYjv1RCS0LYyBznp1bNPLxIJ8LCXIvKxRJlRSID+OBzKURCq2r
PRw23bAqY2YFBDWR1f20UslDMdGPxCxoz2I6U9chg3JcuH9dWWdY7blE1+pePK1x
H5KPveZsYkurNOOJx+K1elBHlVjchj5ripGkJ2Y3KrqKvg/9GSm/JKV86yTBAZy4
h/o3wwlQvydFoQfJvsGWYAJxHjrB7ydLSo0jhcm4SL6jmkNq5UPuqDnbFxjWoIp9
UvB+LJO1cL61AapcyDpG+ylG5UZbeKH7EwWLDLHNHgQ28GD/feoX7Hi9KiKNE/gQ
KVWS2Bmtyb6vf8pP3QJKn0pvyVqddKseCYUkFz1v+aRtGUpz1BicKD3xe4nSpRJP
9y24CDz3US37/jyMVnkVcAR1VU72uhCkA27nLwA7NV/3goF1dcXIK1cwkkPCloFw
yF4f34iJ+h2fBII+hK5vSV01s9nKqEAkSu/nIwAVm5mQ0tNuRys4cKTFEWHy0Wkd
c8Ldnjhc972a8VfvB+lQWoyLEr4q4WzDRF7ChmaE0DMrLVMXiuJvSPSd/WVNhbgi
Ed0cBUA+eYQ1DcMoadKsTUZBeAkMBnl8c6/dhaTSwD+GKLjmBL4N0wgFDoSKvu1F
XJfQCDkvwGKUY7FmGfVhL3ao+k25+7cJmLZhQIqWnggVScagMvoyFg8AL4QsiHSS
EwCkNaFTvCdwgNJc0bOkFd8af3G0vz/slzDOouRCoGHqTVXh0vGPBYWr+Fu+PVCc
3ZYRFrM1K7YFbtENFRMOSIRvaGtp3sG1t3T9E/VFcX52smuD6RY2qHfjd4VBsT0b
sOJapxoGY+xJc7cxqQj+084EoaS2bwqQmPrfU+HJ/TI1Wk86vHTAj0TPp/wOy7Tf
lH8/0aqLcEjSaS5pt2huTFP1i6ZScUa4FrufJav3TijGAinWxhprGnNSC4tQ3Mro
o+hTl5Y0ryic6yj8GKkWCT4G36RXdk8vSaWhDPJOzCSqbOhsgZ6wAAJYmN04G/0y
MrDcN/T76YiWAbfI5b3sxvyVpJ2cHo1GhkOusMNX3Dxu8B36AZxnWw4iBj+eZm39
NBXHJvNFChYaVww4sRuMWvdi7qiWi0S1QyjJCR/YYVpHs+sVKT5TGK4+CvlsTXxs
g1BufYhdEhntKX8q2rkUA/Hu8Ub8GXsPrDZxRgQXljBIYB9R7tD2yNld5NR9A4JZ
ukAayYGdHqTD2GG6ptpm1d7eeLlcPASlxyrN3UpNcXv7le/f0ubcA5jJ3JrRNBic
RLSUxgEyBhRu67nwim/mthwT8sUh/ud+XFmbOzPucX+2Ts1JHIlGgZ9wlZbPNLlv
wwpDymh66YGWixFejuR8YLW2oNdQszA7IYQCh6D5Wwa2bTIdr8ljcHD6ScMoWQw5
s/HhkECSr8CP0jh0J+SR7V8BpQJtFkZPs+vD//f2oi99uX32dEpPS5d0yuuARqkD
CzrhWtv0HH9K47ZxaP6nurfCV2PAoQL4JhYM1x+TOBkcEuUh4m8tClMvTowA3dLM
psDsfblk8OtsTRF/Kh3tPBYBbTqKKlS1LMeqC5V4iaTSi3SKmQvlocy2F2duiXnJ
VsX71KSvWXzBJmpTvG6wfPJwA+uUuLBHdFdmUGo5hiOdlHG+Itfxnt38tTKfHnux
4s145NVybgO9d/gH4q3Zz9fwSCkCyyRx6/msHc2aB9kq75r2xhZKna/SoITA0zvr
g005NUSTPLqN8nfH81GHIUXEu3YtK0PncBmGwRcZ3dOjKLxNBaqLzIqvKFpmXa3Y
ncmoMvx8BDDNBvUqYoC8kDjj4lXunM6UCxax7tRQFmOK9SM9AWuJ0bUHUiVEAOXQ
7TMi2ZebGDRSSIpAG5fDxz8xBd/bYiCTz8ujq39FBPw2KrR6YjTGp2eg2wr2bn54
4Uey/v0GWn7xz0V5zpj+jQgitmoPQPprESDZCSjk9VYiJmOxPWH1qc0RLwbNnroa
En3l9u6Z3bK8sciCyO4+RKSpSSDF23dAvaVA/n6DL6sbMZ1TxJE45WKy844HgazI
PvgbEVGr+P+2eIkAEzjlE1Ztd9AkdxlhV6tF8TikSkQSkKFhvLR62Wg5cGySMG0L
er4+HKvPR7KXMsKw+aKrstICsTRv7cJ2S11GIYgyKM+CeHH0YQ3cTB+7ys8Pt9Jn
6xr10shug+ET0zeEwQA68Ut8R2Nt7Aj9tCBhAjpKZFwAlggBbn6We2NuGmWZDRvj
7MHEhgo+Yo4mF5ih7m0N/uXHZGp7VUBC/g+TP6eO0r2VMbwRFAJlMI4/QYNekEHE
UjsDwfQL/sLxtWawckgX56/oYV9crrj8upikzmQo0uDFDL+Bfs6k4h6uW3UXsoEN
hi0Dkbuz9EFUMj/m7obaVrdsJWDbEf3SypfkmvEolGwiAedThsiMyID/2kb01UX5
ve8w7SEYBOr8MuDH+/Eo9TXV95u5iEH4LIWa477bNHJTw28NCe4Ia0K0FAzw1IGV
ti53RVZQYZ2jyr47EVZVnQiHg/F1h/o92bzt62sICOznwuQh6qhDLAFOxRlxSwGS
EMZcGBO/tqkFUaJ9qnLFMDgVAaluzCwe2v7tp3fZHZCk61Xqp8BPDhij1g76S/l1
5K0YCBWiShULke+UmLH9Drox865gAF4hhg1YIA8nVcENga25yCLCTsmDI0g/Haqt
VEIxwbRALwU4teq6zzhkJgD1AWZLxxnexx9AsRJ7kfRQKJoH5fW59dp2iHoLe8aG
mZpoIcnpDn1weUIdq7K3queMjnp4+HKLY/tydGQ+Rtt8/ISwj427BGAmYjO0vBYA
KHllI+GDJOgQpgPL7C5ovxF1MiRHmXZsTV9GJ6k17ZvmIsaleGNELqI/xBBepeOl
u84YPoBdkKpHCiqeXhFyIvELXeHmfa0XUpdFVQzakFwINahPcK5x9KObjtFk6Nd9
0/4EzSZp3yRdEaJ+s8B6qZ9UHk1xezaFt6t7J2UM41DyMSX4bJZ1iC4RtJEXdinP
YWAXFIx+vscboSTB/ZjCp9iWYnIAZI/lRfu4SAiF+tkxvgmp90bHkrQ2t0uuck8r
wBZbild6Z6ZQ2p5MOmGUHVccKgjsiTO8VM6lMHy9Qt66rqqWjCw77ndkQW/QVZO2
GnK3NvvHnLhg8jM2eYuHk1my24BOV3DJj0cP3GUzRSwPKGHbIaRf4omLAIG2MHvk
DDY6yTMRep8XWUUeG4mEYQ4bE3q2XMj0LJyngI3Y3d/vBZR/XiybBvl9L3B10zfD
r7fASjfvMxhFDgIULZNzXins3v1rvG+eghw2oWy/hQqY2SRBMwNQXHit9qWPwHwg
Bdd3hYxLk4jtbc9n9i+RPDtQ6NtjByFfSmQskCjKqjy+badexoCcktqw+6ldTC1C
/JsmKS/ia6xfBbMzHG5HdmjKaH0K2x4/Uh+SAkm7ZWNHAduDaVSWI43BCgbqVuwx
8WXCWtGF2ctgZWYsfuzYT4C4cYL3ZDL6PfJ7XhFZhexf8/pdVa4uS3WR6mdzsjLS
B3Ou5yWPjo6qdeg01FrkR5ULCzr1hYIwusrXMObIRd6rdOpUiewNldNXbjWYAZpE
7NPWeE6KfAH41IqLJSDrj4lI0SJEkBxkpuDHaz0BO+DMB/I4D5SqpMqt9S5ncLD2
cn31/GoqhsbHhVne4JJ5TCqtB2KntBiJx+4f9sj2o1X+tyINbxJ8jl6LY8mtVuZn
CQIIgYYDYnAvrbuOdGqrtAI6bfh7xB7XJeVY0hDBHWr8AZzzBGDq4+niCmgev2dB
auQQWv0sNYtwOKlgo42mx1ZtYFj9M/CsgQVC6+jWp5XiaQHWCzuV8izGFse7FmqQ
UokO67AXpcuLD6x20psbEFzs4S6oWJFwqXJYeALKlEYKfS4dq0v9DGAmliymWrtC
h1Jr0Hq/TD/OscDElZyd4H2WR4Q9nSO4aVEc7lmvUEZAaadcxSYDqaRX16aT6itz
IWkTef3AhGh71CGsV7WvALjLR0HbV7N+j8WUoba57ObDN+2CpHcnGQ/pnWYfD94N
+qB80jrwe46ThGK8YPvb5q/ylzWwuOup/J6MO/VXO4fLGhCv9l22SAOwNT2Dx9Um
tHIdGX29HuGMVnKUaCVMTXc/2/KC+ykzvZOqKJ6vDVPR3G4pvIXkvU6yEL0+Bsa5
K3UX/mfKgFNdlwZ8TCb3+a9YeYYEqLUxeiZPg3Y9/nh84jIwbr3/eRGhRy5tVA4b
+50qZA5WMlkROUK+WWqkVpwcHFqdJXE0WHyYArvabU3ALKSUgujeP3NOzXYPnLCT
K1acfXoRa2qTTWXsW7yN5PGZ4QUveEUM4INtt1AwWDVaWj/aDds7ksnyeTOqfV5A
VLPs8zCyVfjSr/gKoMEDItJgmG/aAROXYd1xsw6ZuSnVSj1YXnvd2fjot1orLzxg
qpk1i3cBLo1WuM+pdn7YxarxKrwJ67ylvSZmteXI/J3FwwlgnVoQJlSBLJOYThgg
edxfbopEnkSaTitkU5hokUd82Rtj7oy93GQWQ3zQhEMUnvE+sCAEtj+KIVDx2+ZK
GJ6B638GMQZw6ifCdUZUh0sUe0jnmPNHZD1XvuAJGLIGVKqKZu1cw0Fcc+avEiPN
lyjhs+n/Nwpsoa9KuCPQZK01YhY6FXI0dU96pgOAmkh5yPcvqdPXN+01Bg1CLeFR
gIbqOOydq20drZUF+lKqAsPTt9nTDEIMomaQd99y+rqZKgzjL4UDTcaCABD3Runs
oQphrKI2wQGp3A9ZBGrIYnzFPMewtD/ZccTXkK50mvQ7sHEcSrkWPXRk4doB2wTq
aRigyRDOmiqEAekVcKe7ZBZ5abf7e8J8I/WjPEAQGZ852orN/p1FYPVnGS/n4z3L
u/jBu2nFiiMujde7mysXqPCMg2EyWAejGw+SPcwpyqsvwknTleBZYisf5SLwQUNf
MfHRknxYMk6aFTUmQe72LpSlgN+hXIYAFsSpg1se9sHmW5lG2hh9pfas76cxtLx0
pHu136wMF0E6Z7whg0AD9aO5i8cw2B/FFYHV9wVX9VOaomdJquj6d0FW8As8IP0Y
0v1f6pExMDWjU9eyb5ujnopq1rjbj7qqHKQy+7A+n1IoNw//smlQqHdeefEM46Iy
hRXeoTcgFCRgi2WBQ07tmMW0yGDzhbUGbtbWLo3o36sSiF6u9JHzey7kediImjwf
20u1ZzHEyxOF8DQnVuiD/kDT5PGwfj4YGeULvpwH5CqAjOI4Ui/6JYbcOCLBUR2j
iOtC/ByMZqxP2kqelurwTS9sItMI5YHzyS1VZceCw7JtTmAMj8gPuJowNRTqYmoq
6gDv9vrO6rn8BtTuLYImbyhETA25PMuaHrjkOE/lYXCLz/0vo2nZR8SCBYxBHtVU
LkURUVqNujI9IZbCvxgs7W1vV3Iap668AUPy732dpWsezXJ4vBoy423Pnai33de7
4wKjAf7vWbAJM3dDRK+fo4TNksLTgHSjBBLcaVUNsR79fqFpG/WdAojZiWWXvRPr
fcoJuBOZSlcNE+zmf6xXK+09oU7ysWdZ7d6QsSQVQTbF8xXbRG+w5waxUXYkAhIM
S3FIKtP0vqUaBMNvuDo/xhbVoNWQOUwAZPSXibsKU01ICO70/Pdcz3tBIXillwiV
jfed999XCAnxIUK307DQ0+dCYH4BrvPaaNDk8kZlAcbD+GZidR2OtZebgy/N5bdd
nMvZeWgxN6pefPLqi4vqqNm8pEFNaBVzdp8bYRF0KVXiVN/+YRbcS56H6EO7P4xP
FFtL4Tdc4Sl8JSQZ2AiPek5rZiZ+stXmdGnhaRNbgKCwSXkLW8xtvdzkE9sgmgPB
+KurG0pUZHCzDXvMXCeAmPi9RqZzD/9epJTh7tJReIozdShC5Nkd2tBTedxu0Y+Y
OCldY8tqHGsnlx6YawR1oTj6CvHVfhRkzWMRfOQWPEFQaaR4/Lh9xExyH43jlWIT
sM/+UIYthYKlK450G+1aP2KnXBvRtkj4iairrKJ0THqJC7dim71U8cJTwIhzOl2p
se5+4UcntosLuY8PG4CIR2iGUJFvSEu4LGbyKx0EH54vpaxnHZ8EEsdZDJHyyj7K
5mxk4jOfSlWO9Y0fw/vfvQedYLrSxdIC4wAsPioOPJmJakDseMibyYz0CXqUV0Bm
+kbjlUGqTOMabW2pMxlEX7o3iayS5Usnb1Ic3l+GJEunc625AJswvEPl0DU+B0Gq
RINVssHS6w6UcjxCsihRFK5SolYMtxBMIJVFqcEGjKDPlcuJ3V3Frl8fHGz8HXU5
46aV42UVfWZoCdwNqakzmYnjh1r/D8d6n1ocgGareeD9GcjmibdyOx/mmkEfIjQk
eocMtTBPWRwN9+u/gZ6Si7H8EWRKh/04enVgFi5W9v3IwguBAaS+yyNVAmbiCNO5
Se+vMNf4OvIzvbeSBFJz6uVqpbS5G5dQKx+7afffqBDAp98b49oqK6Te9jKwRtua
PHoIJOFWACEqd3Qx8EaneMwmDsg3YBQQh34ItTgdX1CM80aN7to+WeqaOzZ9+kWZ
HJqCnviWBctRg2g9wUpe4mTO5Tu0K+M+LJP2xYtyzCERvVn9eSzKx219+e2a2RuL
34UTi0P7KQcgg2+ORGOVW7Krd7DmBGvO0oUPAY+ZNdus0mbaIbLGbDIZRtwghiR7
wpZi28X1FMGbGafeV04A4eLAFH/tBvzinhXi/zW+CkqA50i40JC3qbeDgwcr2gNF
v9JCX7XOHTXfaVi9k/PgGkzI69Yzqn5sLWMY2wHnjmtt6Drrw5SE6B5+DIMkhti7
q98Eg825Z05tUrcsBqAt/rGcCf/ukF8INC/ejFB/C+GEREr14zPdF1sXgPhQDr0S
iQT/fLiBf1uPtRPQ6mCXINs68UMMU9c7/LJE8uHcmY3VsvhFNr/dGGWy0owniDUV
36YdLMr448VnDymE23KjAnoG7H4Wdl5IaQ3GLbdZyvvzUJlDa/rNyjc1afLXFReS
kfNJkT6O1ld8yJwm07Hj4eOGj+vC6oZHwkVPilABh5C1nSYS5/u73HGgiL5Ke0Rn
yD0yB4JfeQbc9flOhHjmvgVpSqtPP0FiS85E/Ssd9nO48mpPZOvt+zUz/C/ECZD8
ZrJOOscfjK3AcqXDzCFf6o3gUHCWqpJEWiN/XD4IzXw8jx5wjHcxdlr7pBxrvYFU
DF14MzgJCU3ApgSwDHFivkw7zuGwrNrfe6n0frMNSd2VNurI6ycX2Lee7ih+NX6F
KK9OQ+1+0/9GqfJ/U0stYRJNxKZQZ/3icgA2RDnZLEnsNgdXdH/uj5Q2VIc2aBZF
RoineovIqXlVRjay1wj/fEgvNeC6mgrLSUI4YJ5qui33MRIIRpGdpzrJj/uzcAgi
0Ga+mgfbmyy09FrrNiPAXWGL2r66FR/yB0T3fsya2DsXYrtqT+YStzjdeFrIy7qe
+9tfCopJx/VAu4h2sKDJrS2kNVkOK8pVqXcwdus0jIfQOK94Gaq08W+qUJeET33U
SIIQXme3yAUYPWCER02WAKgwnhKui4u91kNcInnvBlXRpuxjlkttRncotPA+qvg3
UHmee5a4VRPOOrVHLw0FUoCx/yXlZdisg6Ho7VBL2d9W5Ho7PKGlKbZmxQjZ6aRD
4Vb3sH5IFSReXcXx7vc/IrZC3KAlzs/X8Re7yXwOcOjCbnla2CT9slRB7PxOPR8T
jYjw71HnMubhLwrPAmMhzyppztgHMPH27NGrrXE04R1QVF2O6y684K/Vyzn02X5h
+hGubZCdCUuUXHFfpva8GOHaWYjAJ3j1yQYKn2ThRrWqxKLqV/pBraagZuhjORQQ
4P72eGWDBe6DN8TiiwZfmjEOclj9825P5CD5jP7h1/Z5OSezHr5j0UM55nLYri34
uW0INoc1AxXUr9yBBPYti6/tltCZ3kp3sNjEax5Ve+9WBv/d8U2CdkAa6j8OKKbk
hGHrhHT/gZbpd3fwe4bMdaJWUf1hlOY8vH8kUHfUx2Gy83H0r70b+vbvziLgYxhw
yXAiMEmUgTR15modTF/ipogIe9/KSUZ9lH5cx1R2TkYSARS8JIn7Usf1PctghTuG
gJ0Ve1LQ0iJ7xLB5PyiQPgEkypBrFW2Z3WMlnLmYwY/iYfkPl8E998Q3OGZdWRXh
psyqBtN/eSVHPQuX65cgDnLiljm0Il5r3JjLSYf8FRVIe1QDih//ANAGosxg/a44
V2ZT2KO+qGs7dWJfJqh61rztVrZso5uR7Pv5q3z3iqabAT9uUuyo4zZjs3lNcEQz
JohgUwDlwXSOrWqB4pCDh5rFc3zr640Y/tpjwM+3wIK46xO7baqa087/BFr982P8
kaDdArMBq6HBsDe5ehRFhspiRSH9ZL5hjmp02bW2sWpKDvFRQaVcJa8bWCkj7cPU
QujTy8cOFEaRU9ljOzElcTm1Pzyh8Cw3QgElOEjyzXPE8jrp/TbQcob1jjwiWEti
BNxG5evctze0g04pkzPQ7HJAVV4N2jz5+mqOjDe/vVNgaCMDhYoobzCmygfAHqik
UBlDa529jWlU7boZfLQfZg+yeLf9Farh9UhMUozGJS6MeckRtSJk+YrC6nwV3l7T
AnFGgpdtWgZT/QyXand7xw4xcQGoDgVI2CbXMKGBSfP8mZGNEahD/oeYz6kgltlE
zuAWoH0UI8nYq+hEUk7nwJ1IF5GGtSXYA2750UvVSuhpkHjuIqyRLTiqZKLTLjuU
/7nD8ArYO5PyloSnJSL5jVDn8NcQuD24OmF7DkqWmeX13b8HCTEVjaz7JjuhLT2Y
ehycxxakG1YW8K2HOxaISVATzn9LeTj8puZr0kYmLcrYGFss/VYxFeVbJhe5gcxl
9zNkYYiRv50RRiJbeq9L5SqFTJQDZLSThzAvXUnxIIstMuM8psrhDQBYv+2Q21N6
ilJlQk46Ilq8l65tlmMVvRJLq0SAIV2gped2UV9WFlCEIYQqL0yXS5dhBaPStoes
vTkb0gud/Gc9oxpY//GI0oBDGs4O8r0x01lXH8sTsBgDpsXIO5LnjIgSXZZLf+H1
SqlMe4lfJFcYE4eH8EHpBcHXryqSxdketjKo5Y7Dz9alTjd0NxPxtbAg6UnJyHin
rmB1PEY/bBaMpMj0kV47huT1Cbj7hodWflnoeQWlHyR2o/edOuflovFeMCFKdkGr
4o4EpUARBVYYtEK8V+yOQ1yvSKp7CYuw5jtNTA/un6TUXVP1ac9PpVTjW+MZ3p//
sunOZOwDan0Iw5wVZkWQmi2ZMdbS9pGku34fADwbpcS8k2B1652jhtkSb2L72c+Q
+N6zZF7JR365jayHHzIx4oPB7XEmN8wQ3XVQ2O5BVxlX9jU0xpx00LJ1ICKYBRzm
Gj58549u53bgjo+lN0zlyFieK0EFgr1YkCL3qhIxioARRQKYcGD4wWuCAPJb5DrY
hmyi9oYvfhrN7Nyq/Y0mGpJylnQwZN1MS4tA0VVuYXouxd7CLT5Eum4y4ZwUSMAg
pigR+mWSwjFbIEoeOhrBvzrJA05t2rTXWni4YbEinVew02M8+xzZA91wOC1UX5dR
lfuRFhWCZqPlTwBJPvDmnTW+kleq1HMnSEh20w20+XNg5SAUZfxMIN4ycVWCHfVz
ZaMwr0kesjVijIqsLVaOnQ2VzPA0TxIjtNIDK8/KX7/E/g8/LAI3iYuXnagVyFO7
xKl7leY1Etybfbq0BTQwBa7bugw/+1C5AivTlnR07Fm4jsi7VFSJFOjozpNtLb0J
WH44rEiIkpsrH9E9wNje9sbxIA4qF8FPTbg4Q7UcEz63cPEs58zEryuCcu8HJi+F
smUVkk+AdYKowQpdXGCuaQiJEz77oG8XGbwvixwYVxvrZPeuJgVQ7yh9YK3hH+39
/B3GEfhEVyEOdi8SIwyjFcqufFcntg0ZRA5XldwH+rRJ91d4beANXm6vu+bpJVST
H4EPA5orRNjPWcOMdMUaoi+HgpyIFJnv8s6uvwQJlVUUf86D9pOTiFOgWXdra8jF
elIHWyaUrSoxU7F97+lkaqc0/LP7GM68SUaFmxUnuiXIyQD85BCe6moLDGBGmH8e
ZStNO4q2n5PXD4c9nZculPLgFPSVvGfTZCVq7holNVObxp2WLIiAJTrCn/c3G4e4
xlz8N5IyCkOriVk1tHGJZLNHzDrO9p+z6OA0yBVTOrwjwFHVfAg2ju3jkXY9pgJ2
9YZtIxPpxBHITo2wMgDoieoImwp9mGYMcHUb0nq52pwKdl8QMH06N2iTcO2kYorN
qqMLKs16ht5mVww1/Spv04Pz1wM7C/umjwMDTAubAyYmtpitZayBzYMX1WL1YGjE
2LA87VTrGCIT7wbb1IQk7Q2677VoTeT7yeavR0bMDBWY+XqbPNjrYJJcuoedqKdL
ZijiPd5j8hV1D40xU23Fx3j/dg84E6ZGBXKJI3EkYOIU55/OD9s2fxqtzjVAlQFT
ATXKUXA/Wbo/56KBlHc6VRVZky/lMhMGWqPo6QbpvHqLLhY8P6nlbf+s5Q9Omls6
y1Ag5M19iPXatlR8nVJV55NRQ87BqzJEhy2zCUzW7TOv3WaP7czF2s6QdOzAor9n
/odce65Ur4FU2IZvCi8gu+mBReT/M1pOqefJ1uwYw34icbB1A9OQcFbBNIDDUYE6
sNRI2YgqOz7kwXn2DxSkHz6fPzTRy7lS+GljG8Ota5yQsAl52eIcTusoR5q96Hog
cpmFTp9ymkhlqoZI0W6G8e/yenpaoRkYWOjevW47V0t3NBfJN3KgmN9ga0+QYjN6
hrk/CjCYkLTMBNcCrvDXneUr4zqC4NMT8P33SwUl0wk9Gy0V2EpZUvJO7mOO/mgL
Q441ET5NxX96xZRDRYUvEUmNHqKQPqetmGysW8ZLJDN+8fw7LeV6o9rKbljqCjwl
OlheIfc1+Ch0peU+Qz3hHUDZedEGWTAKcBxW4PcAvkT9R0bf2AAUetLG+B8+21xE
k0Pn2fDjcy0MbHep8SjS6q2DxH8L+NO9nEMZ186XBfSGALNZPZRD/Rf88TmxW1e2
jfGZBhnARtZjLrMlk2fkrkAdKcJ1Ln+FuVyWe/tWD3v5r7PfqEZcrMFMTdclIlPj
qUS/sXC48FkPg/JliVkoD7UrGcyqxzFbV3Zbm/ij3QmIiv0bZGqCq3GzgvmCiOcy
x4jN8NQr9ztjuuo+B9keUjhdLH9XwEepyJuQV6La0iUZmb7FOMquPyfxUpwszgmR
MJ1KEU4NmGbUIEBg5zB7iRbVRxZDYqtV5D4K2LdftTlXFtynZFElLLRb9lpkKtI6
mKXSmCW3bgNbtsmFNpY3OKDFtYBJ6NL8NEGZlVhHC5OXCSrHh9GnQnTvVGKLRAmK
xqUydOY3uT2ZB40txCM+3Ry/CFOVeRLGBJZ6K7h/9TpucuTw+3XjW6cM5B8yxbgF
bppB4iEU3D2j+Lp3Sst8WH0j+b5xmJK+LvEQkFj1jUNwaVIIUK87mfLt8PGZZ2AU
6gwzs5EWufva/k5rqZ+y4zCMleQUiZLY1bWvXYUczUb7dQql+yosrXJPFVhf/Al3
79ppnhgODM5vWxFAD84TfeDWPQ7Ae15H1ZQCN5rCoU6RD2Dc29nivRrBEVtRWSnt
3XZ/AEesmsg+M1oB0Ax++ct0Jm4xUpBPAFBRHoUPiwM1dAZgP266p8wGCLhHK2GX
ErPJomp4T6rZQklPe3JdNz4s8PJsJKSgB3sF7s1u864co8tGrpoHI2JCwkil0zx5
QU81DvtlGjIEjKv9/ycpwCLjUJgwUXGfZJvwwNc9L4OJlKljOcr58vJO7pAI/k+E
LZiqSgP8BHxVzu17fssq77zRZ26sGfMT6an/Dak0Pf1G2CDiUr8NuhVSd2rmPJx5
vu0Q+km7b3ItYugqJrISdLs50lypHHeuMp+5ORxSX61QIvzQ7hlZexPrwq7IL2X2
zZMG6pxJPy0iPyOiMW2+kN9a8QMgPf7uHPp39I617MxPKSNGGn6SYnmh4UW3jOge
bhnD4JW2BzH7wYqS3r4zUIcnUgmkNPMTRMXCTGo7vzSEV5Ez5e4bLMeEruTdeoEI
ViyJ+/5/dy9ybVkdWrLy7NQgi2NvmW4RL5LrbSkpgdb1fhhwnSHkoeA9jmOKmeqd
dLaHygNzhsdg2pCQjMS84obxQUlwgJC/6bj99G5vbQBt7DUr2CKV7YDVx6aedsqE
+TAxMu/ZCT1BegSqVbfUh7sNwi6PF2Rr3cXHecBTCP9RmqQa1UAVaMJQdqHxZsK2
xNJ7N9u4a1pJnYA/gdUFZ00gziQIaoflYM9aODaHySpc14difgSkGcZCVWAcKECc
lwFGgSSOs43F727svxIItQ+jU0gJ9KR296lPy5qx6/17IlbRqq0wp+hGJ0+AesKI
7XRSEvX1N4mmgtxSY/LXKjW2LPst7QEquQqae3L9bmnAgDDlUPMMNUx2c83kabBP
pdfMx0YPPo/JoZ2I8FfHcw9Z/SCk4WlUWlMPCQH5yhHjNSuRf48utcRNS0wuFFXu
6Nue4v5CXIcgR+WsGOWxu3IUAZ7zPzLEsLlncq4m6uh9mYNhuRJ1apqMkAuOdaPj
an0UikLAHB1w8pHejd0GiqpDiZQOff0Sm4bZuzrMxr2v7vkoeHLKfA/vVdwK7/oN
EDx6WV4kThb7BDcIH3sDRbXqZ0N+Ayz77fvqLpjf+BCYIRBW9QcRv5uXL/LImuvB
ZTLgR8bOyYwQMVoJS+KIez+FqwpTZFv4G8aa07i7fshbFo0Tf6S4HJ1579n/izn7
Y0kmd0tkDOgfeVCFlO0i97djvBaySB7sxyKg1RjXvvQ2AAlo6bMyiVDt+h/Y30hI
w0At901NFlpiauPA//Zp711IYyz073xkpmDA8xKB31Gw/EeP3LVojTCM93xx2R5p
MIsVaWQNcybueQZbhKRPLlTwKwE7zQ/ozSk85DSZK+XsiwvH64MAnxOKFZoMZKcv
LZKtDb3nNW/5ej2OHjGFmxxivzv/6iZVsGUaCZjrTF9rbCrJjg6shAJC2cPcmbAV
Yq/XcpIieXXgVopti5jWsCXEcpz23w8uztVBdT2JQ5bNIIGo/zdYYnD9JgI40Cw/
ryRDxspzrzCzEj/3WgtPHqwS3ThOWSab//VmIjDmdc0kajtHoFNKmZMkcY4AVf8i
DDk+WCruQ5VqKfTfnFZqvxRFeWxFXBrXo1HPL0S2mlmuGJ1Cf/TgGxUQ9zRAUsWB
BmiZwps+TJ4UFig8rlqeFunQh4dcRov80xDShjrZxXyPe7Fb6E14udrieof8oRxL
`protect END_PROTECTED
