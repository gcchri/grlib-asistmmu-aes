`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d6gD+wAM8nwvyHF6d5dG+2ziqKm1VfFsd6OoaIO9dhp+1NlO49KwORFL8qqRobG7
LMwktLsUxwrORMualjrkjLS98ZLjoY5b2SkF3ueWPH51I2e7qfB2ZyXTJ1mFA+7n
8cxwJdlFavdMDqOs9GRSufNwtrUspnX45p4Ap10R7FCyWqr/qwZGmyEpq4h46ybj
GNQvRIjaFmZUSjHwsSpU9Ao7Ljemavi/Oc1M4DSQZNZa82JD6a5QIvhQYcVAOXR3
jHYzV+EvQYi3N9A3DSWpqg==
`protect END_PROTECTED
