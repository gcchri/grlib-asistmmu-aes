`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7VFPyBujEvsHbh4vM9ao3Yeg7hXJrAJULkVFvqW1CVZcMKVqIEmISOss8B5foNg
JTOwC2ms6YhABC7K5Wzh5EQcc1lErp+0mRTThF4/SP8YwQnXjgJVhfLyNT3/Nzpq
VtYxKcwtvEBWl7JdvTru26MIyOqdo6L5x/sMxoK6RGIO1yZ9VSHNzgHYnsf8JTnt
4x8HVW3EQprGRyJ+j+Jw/miUUBmM3inap6sJXTyfPT8olpKQCAU9t9cr7QGRKTCk
LWje8Z+effrBy6/zgaYMz5EX8GLn0cu6uti99QL/GHRrTgFpnkZQIO0KqxPlmtzO
jscG6SD1X6WxaganplvvxV8v0Q5ADNtAFaDqJtJ1ZQ+1WF8zKBQ/dTfr77b/Pt5r
`protect END_PROTECTED
