`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SP+swPeV1zJRiftX2JibmvMyGjExvsQYQaFdhY5kWCWxCVfvWMefOa+xjjaWrRyw
YP59A4HbVc/YFgOaWchn8jH9r0gRV0I7HUGus/8qINUQMwUMh0wnWWSwzfsd/3QN
j6v6y6EuJ5oOJhbtCnfcNxrUIheX5q+IJ6y0XZ7nRDtD2MVG/B0/mbszI1RvLfNW
+TVsh/127qSCU8fS6EpJjv4ErkuhjKcEzYVe3YHIyGFoAPEsf+Gmc1SwydqYKozQ
0QqVLMokPPpG2xGwB1rrDmfgEKaIEbE3/H9VAAoWDRQNQ2ffE8CzwBkjlHlozCde
hUbxDNE4dQoOtAZ4/Zk/4A0KCm8AX+VZ4P4dP9tKhabYiVkRSAYE3pD2Mp5ZzQ6f
w9QgrXClGnpNp2rc7BTzmzH7pmmi40BUbaoqdi7KaAIlS2SNpplz/q7cXSyXzbCy
nN4zEU/Qwzy2phhdj8qAPuNSxWDpLGc3SbK0Ym30PpUWxhOi4ukFRk9tqHy69ATb
uskUmE6S6dsh+MLi58zB9ZyUTXjQcoetjz+UtATARJttpYfQL/CDEy0O7dDjuZt2
0G5ONKeaLSim2p6STo1Bf4xOcNOuDKB3cI3hAZFy/ZKszc+oaxcQnlbQrF5l4xUV
HpTOEMJUnJXhbvpX4X0UZEXrMsqhbSbh3TNnEkOQ7vgAUceAm4L6/CxGXMZ1PaYf
mUT/6wgX6l+ZqioynVIwagVWcREEwu+TkxuX8+6k3bZkwwazUxMSGkCrBRyUsWaa
dY+Q4IreW1/t6jMbwrzfY4H8wecuP/KfbxOG/xNnhTIHBQRkJzGiMuwQxZ40h5Rj
AXG3mdcpVfRvY2c89ncNOc3xE/L5E6Kuy6GSHys9jLWZnqLsxAYA+hL5T3kfcjco
BqEIBwJlgrswzFhi4Oy/McG/0xn+pXObyaicc37YzIbYI2XvOi3zr0c78p2UUuAk
mGAfl5RHiF1qA1tihViyJt3SlIJE4OF+tAHvFNcWJ1h7Ye6cab4QYpgLBBEIvj2J
bkC6EPniR1O/5tlMiZsq+0ZvzkZVFnu4RGd5aySFzGnJRWOk+u1S1mSOFNgcCeM3
AThQ6KODNFyI6g6ca1iR7P2pqghS79fiDtmQAyjSdFztBHeKZjcIGCx1BLMLOXjR
Z1UmxlKbuTEiiO7PGs75lSCrhvBDZR4aB/9Feal610eULbSqKVS7CaXkqiqhVlej
8ezy/okwwhVhfocY2gWqo6qFYO84h44dROMF2n8JNEt+0kSHnah9WYXhCXsuAE9L
Bymn4YtutZFgEqGqm0X7AqQzbwTuR3u9XCIpDUhXSgrRi4ZOtNgqmxFAmFtxDYrr
16J4U46//nE/zoeHhW8rzAWF5nAykHwcdpePV+FCr1/08yi5FDBP9rDmanD9mHHA
`protect END_PROTECTED
