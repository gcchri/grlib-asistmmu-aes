`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7kRscY3PNCyrWaMsJxTiAabmMJ9fueRof1uW9sRZhxdWekmA9BQyym0FK92LzQRE
trlarLFh57j22nGl/2oBuXMte6Nk9LtEFsOZIQxdF50DwFNrYPIWWCMhEpAJb20R
e1Wp//+wgVtFAdEwd0V9ux+IF4mbemdLuaBunIAaYzAyl2CJCijva1Et+aBFQyxI
Ckw3XeXzHlXI6HzQzREL+q2LMCoSp7wqHSm3fdb1dha7KzHnWTpzW7/9TXVlYD8R
rd87KHlnku1DIxF9/9TYQ3T9/nPIS+xzu1rw2aCAfD2SVQyIYE9J32GjWogkpfPo
GwhwGp5KZlkBlwjsyLQYaJ918vnTh0IJkO/G/Z6Vt9pxND4oBWuov1lYHn1ruKfY
rtqi5I3XSoGEeK3B2zy9aM1ehGPH+lbgQRJpEK18wJnorAQBvIV2qAibcccd8cqu
p0UHlqJd2mFz1iHkleNJ0uotZqoTLkux/ineyfkPOMYTbr7BucsZ/KgVkTKeEGue
`protect END_PROTECTED
