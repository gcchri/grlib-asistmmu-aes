`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkmxwKJMb91hCgSezFauBFnmHw7Pd+WgMUzOY9GY85eRpLW/t1WbDMtABcJXKrcj
WK8RD4PbznFJ4gP+z+RpFI0PMBIGqcnirvgQ8HvJDDc+ggGUKb6c2kIJMzwgX+Gg
wNsrVEQyBYIGpmRsoWjVO7JV7EmwGyixG3xp9N6pdFBpxFgOJXGANcsGtkNhBMY2
5ODTZE7Csh6U6pLKsYZgpPn7xXpa/JtsTleWGfpid3358o6rFTDbv15TCx8ckkZa
KeQhodLc1PErO+u9dGpqxdtQYUODyAT9eWVe4jgoyQYVF4D4yVFusTpOXzVaqBO6
5CjVTb/rfe6Ga4hDdK7yhx8rthIJyKkhR8inDDdUltVuiiboOwP2nZwtSyNPKvkA
2pMvRN2X3DEFlxWa8g6kN1n9BcJrM2+YMaZ27fB7Q6xULoekIlOzmqluKJSoWQha
Rncx14qfmIFLaP/5QUthmadZJxXJU08PuqZHFqxvj8QC98JGjln6lTX3Vy7hapw6
Dj2j9MQX8jd/+kQNcarYm85Onao8Pjz+YK1WYp9WAZXWG6I+D/qRhrdfvgcwk5z8
9jnXmM0UgFZAsPBXrcfeAi9AU4vK073Fhs6V84GbrUswejQ1bdAPOSv+a779rlGj
wRNzwdK2HFTYyxBXWtxyxWzw3TW1/CIPRknaMtTuDB7fX2xpNgJ0p3Mlc/WMlxaN
yV4TokXDFU8ZnwjqMGdC7u+sgPWFoPATKfeS4PbEGU7hcNMILOabarwS4r2CMIFA
ucRwkBKm2fnFiGnxOrMwxYYLt0weTUaJ7lwVNCa3qQgNoC8mQUHz4PS8pARnOmEa
cLpadhl24GwCijERdkIgvehmR3/W32sOEUiSxmeyMhIb1Ae4JypHYMCNsFpjVvqY
eahuArhTNxq+fvA9WGTkSv5C85GL7l/8DulgmnsmMswDZ0Fq6t4LQLGysVGu/63F
+qudVkX/nyss5O5h9Yq6SQN3jkEzW/oe1Q2njin2ErTIjIcMWo8Mc3k2F+0oitS9
RqyH+cdhufHUc4HsGXd5H3h/T8/IopF8aMv530amZpORjVC8bgz8AO027Ys0e8kv
PncNkHckN/6CRbLpQib1NJ4vu3jaA1oXfn5nGoCtcs2K4vbrXfmVDOGd9RMUGPam
mRW7h4HzSDT3+LSkq52Z2BAvpc53No0zoHS6d31jGK6tBMrIa9T9UX0qJKoMmh+0
QOIWGorfo02SveCxcGw4Awri7ycIjJ7rt76A3rckARKdFmrW95CB8vVny1Fv29d+
Vv+MVRsX3GeBcP9AZx1atqGA5uvTO6MN9iRHrAeRr9uJQMDkubfl5MWWRR396etW
DCDXFs8F85aOZ6VAoMl9SV9eLW5/FpZdFI0I5x5NSaW2av0SmWcAbhuQFq1WNTZr
jVSOJJaHJfNp7oSAL0UU3T9uBJR2c91PeZMKbq4mYEaWYMSTVFqc3qOU+5Ope5GA
AzQdSjmcXuDyF7Yyh+Uiwh0bHUh6DNW9kuy7S2PQfHE4KGS9dx254yRWHqoB+xca
73BTKB7JMCzePyqRW6P62C0SRC+XZSom7z5EC7H+cqf4ALr6gfO9eJOY7gkxq8+v
DOlOgNWDdLH0AdJkpwwQMMUGHzSRh+5lmKDebu8LVUkctJwBl/UkVCWvHxhncFR+
8MGyjhBywzEXe+6ul5io4qiG3OhhE+UKvhKL0/urKfuWmZB9tKgSgqZJUvUt+FRe
chw5xgyOI3oy146ipAowJFFrGGp2Yi++nO1fZH38YyiHIq3eQW8N8bYzebKRMtmr
Xr0nUmIQHPZTn4Xm+714aRORYUKxC5xEeZ1hLVQ0I4LRprH08NJTxcf27Ae7Ib/t
8fqX4D/8DTupFIAVlaTUBLGol74jqwsxx4fA/fkGyG+A7cu5kfrlCEFV1s7u92VR
uKQ4V0m1m3md2vEwQQdHLS7z5Y9jV9MEsv8sX9Uh6e0R9OSUrGq7N9Pw3FolpN5W
7QdRkmNric8lLsXJXhyRBrpvlHE6wsgWdDoAGN5enrIn1YhJsKU7t4oc8aYRnQJg
HbS6iVR7gVLRzZIdhd6DnXGfzXEtcjTs/D+bbqZGN6p7SStO76vXk3TSHksu6V58
QBSeo42bNh6rHGaFYvwmNXHPAaJ7Mqf2ZdNXOq/PPrKc99p5l/ezSBWeL3bsloNH
ZJ3+gMfq3lK6PyFqmdqGZJGiz9GOUVYQvwnuGcp9gCj0c9ZOr9zZMJcCYtJWxJNS
RmijINCj6IAwJ1Ar/Fqehdv3MARuCYDRcYf2Pva/MQoStRfXnoX5NYQ8VRi57nBF
R6afN/LBykzyJ7z9VnnJWK6Cz30pFcCo7cgu0Ie3WAAWpYPHG6Gc7l+8i3ViBL5H
+dDN9Uz/BU2QtmqDLh7VYe57lZVqqaavlrOiq4m04BiejnwLP7/N2PlOA0T787p2
N3u6RiNiktLoFSm4z0XXzxBUBklnNr+Nt7moyt65lP0TOdz5ey5K9GAVDxbGNBKy
pxTVkx5rm51AS8zR/x2oWbwgOdwCa3boOkMnJbaeaxvPyb1etHhqZ5btP6NEzijZ
eFSa8P9iCNTRBuPaLlYls+EIg/FKkhxMqxkBjedR0Ni3t/rw/p2et6DPLG/P0WQT
PUSHPmHC3HBdsAqYGlxDqkFeHmHNEvjvTaiVBR2gAPTYs9wGJSA/381Z9BRiL0fO
+MM0tnW4F73/kZxSZ/P4iHwKaMAlkoi6iwCWSJ+mp0esAdHF6EV8YpJZ2CVEQWtC
OQZmVsIFcx/Hx5GpQFeNdCd99bUXMncUTQ1vuwHlPx3B2T78TBRwFzScbpdIEC6Y
/floTTy2AfTscOgn6RxCVVLtbLh49E0dV5bdWIt9HYFPCE64kpzwEJx4sx+hNkxM
xYsjrH88uKJSsn++KUbvICguNr1HIFc5jr1k/Gde5y2w6/09WBHQ3BdkgHLn5uqK
NBVfZnfZXlkOULAapdsS+RVAVh6gG2DghvsDQEc6fgzR8uTC1AGa/kbg1T577kYy
yCyNEjK5wDeb1NA6sX7J6nQVowF+CVI60pGeOltD6LzZ8YrqAEkdcA5m3mR4oY8K
EKQFdzrzSfghfivZfCXMwPe4s/rCM+tALALo7zujyob+aETteRVJrI8vd+0l+f9y
`protect END_PROTECTED
