`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l85Jc8Qz2YKbDWVk9NoeJ9TfYrOZJpeRGU1g/e7fKxnEthBUUXlK3C/59qBu1avs
/oNyJT9MimnDSn4rzRHimhSr9PNw0qAxCQqWRBxs/UCW+WSyqRKtyzc8VkDkYhGn
52VlVFGDyvtgswB27AQWPU3hLoSRlvAPxUaiA7Tv+pZ6LeKrOxghvp0QmB235EvI
ByF1WvN4d3OU76e6AEZiDkx6PA1YdqP64ee7ugJb/8+PHZ48MsN2xFVR5PsqXDFE
Y8+hSE/9a87BGo2JJYOA2uSheGs9VAfCokt29j+sYzALipplKPXc7PlM7DVLgf/s
ojDa3tmZ6hx485ac1Jl7+dd+XJXtY/U25ABTnX8pvSJ3IM5SsuGd/YldG5N0tGLj
is9qorqU/U5/viBgiPKulSbwWvKGO67l0eWwrFDv9bslRe6X6qpX2J7OUROS0j4V
f6CFD5UVENscKu5GqFCv7pW5F9jh1okWfKjo5qguRgU=
`protect END_PROTECTED
