`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/h+aOWQ6Kea0wwFvhMKQZOJtRZDmChUG4XvTSP2h84cd880FwkM0YSJfUGvGB9y
Q6itLxNW6KbHc4FUlP4Fw5JMUTByssCGtnrwzFSTw2fI/+5Ayo9o3TBP153ih4KY
agoe0kxXYaXJDDeJi5yymV/WfA8ynElYdtNqH1VWeSbUy8Q7PJEEyeC2CHXgpZph
9sY1QgueAEmK6fNkkiTzFPG+XNJTrEm0i0N1H6GQDTVg6xU3MO8u++u7VcpSLNmq
1JcOAZSV91clGkejMMtqvGYU6Q5RaR9ZxU6jZ7JTm7loSo5Ql+UqjP+1fsHBg02M
FoXaxlgJ6kL5fhRJu6CCljqsdqJSvArr3rdUghPTUCdZsunvnysHevz6yUskzefX
oZ1vJxwtBy7klJ3xMDfMD5Neg7EdtAxo4ORDI51OI3lF35qR0ZLYtpUnSMIsBp3q
x0APCSeG4pz2wiuAHnI7TJ8Ui/zGanxBBscu20gu/A8Ppna+nngTGwvx9Eep0vaN
pJVikvYCBvUD54cejZY9ZMS9UKblaasdg/yXXnd3DtQ9J6HK895BNxsZFdiBR80d
hvV9LB3ckp34wAfjX+qmQFMV3A7IlUYytBucb3m/VCNOM/kSbuRlHom6GbEC03WD
OeuUeTXUTVxrdy2ZqJoIRtzevyApflIUky7tjp7kduXdN54xePSQPd3DuQ1vD/bL
IdzsWcR4vlkFtMNsPDDTXhv3aqTdyo1DzoSGYdf6EGU=
`protect END_PROTECTED
