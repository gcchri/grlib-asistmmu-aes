`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0EKzv5j11eWZbXSQSBj3EjrvQy5yAkpEzwgGwIlWv9ZIQrHFDHttEmeU5ynaTQ3
E1GjNReAGESAG2R1BSI0+mMlJw5Na5XGGX4NbxcZ8bInHHGmTtv4Fqqa+Sx43zU5
6ZiAgOcgQ2jcLJq3HpJvqW9qGLpgoL0gOaICce4nY1mKKUxE+YcCa2FPrQjYM8CC
GO0vdBBYBobxN8QiKpaZF1zalNHowChVN2DwZwTy9z8nfG53RrQxIGcSSv0jYYVA
`protect END_PROTECTED
