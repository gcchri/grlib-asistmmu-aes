`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVxSc3xQE7kcwdfjxfdd2gjb3aiQDm6fG3L/5Hi6kguE3tPc9vhh6iqGrxN8IdWp
no48wou2Ca+qo1DjJ8b7ZKBFKcDOztZwUQ5cEbvTfQj+F0XlUIIbf8uBODuqAMtc
I3fJgcZ4KnMw0i/aglNp/PSpNBhChvzYf1c0j2zU9wdqPYpbRMu8wslttbREz2z/
4FF3tx/VqLSAK5G/jqvH2BEH2MhE4gKI0l/q2VOU/N4xsRXnXgTz2hh+j3AtEsrU
+7VJogg2usvVrzB2rMjL3bu4lc9kbfZGyWJ2Is/KCmLMp/hseoGq5meUXbHEE32T
cM51UMSbeC3dy70KFZrh2nTAb6Aue7C8CGA5dbd/IKy0k/xerhejc+ScFXkda6Ek
DTwRC0MJ2MCLZsywEJL5UVBc0pt93CL554Ekv3IdMpHwWYDfXnFd1UYZKv3608Zw
asXfteP/Dv8Ouv8HFWEvgbAbthibiTV/RUjjC8rU3lmL4v2WwjQsQ4PMNainrxfT
+JU9d2FvXsG8pqimf8cxo+tDcFuevhQ40yYEEsEeQDLoX2K0OjuT3mpDd3ZVK1R2
zCyKZuF1e2kPXrmFnLEtFl4qq5mFezvwi6v8+TVIZdl06KkbXDPGDqqRc0zBD1tT
zMJMB/wOQfewjHmSY7ihTJs3pIo6eMeRTCQ2mhSOvUVXyKpXsbsqVQRx3ckddLeL
1cCUuzv45DGdK7Yjt7sESkcdbhvbOGeo4i76hoNxxd7DIJPMZZJPZQkxbdB108Ya
iVL+FxdOBOGKBNrHdJw5deUl+LqcDx0WBG8vEUkblIUsAPgzzzYKvI81+VZCqaDN
wogdUUfw2X/IaiUgDg0rWZEPKahtr4GNswR4oV48nZH3AAvX5iYJ6L+TaTtc2bzf
uguiWxRvUMTxmGw9ALFNmbyhPvQl4LeqIajNHrRDR7d7UpggIt4dkCanWEkEz6Nh
trokLyDgsGJ8mmNkiY+yy6/Uc7vb+cWDVBuGT5fTMP7FxIAefM2DBLkJtO1U+kHa
VbPa6FsnxBEzrTNTMbXwF6gpbhwmUJ8ZFv6G8x02+PTCYUFqOv0GdiDOT7l+sOXr
9R+G7siGqUw+YOedGTxzBuPJ7dYHb47xQvzRbr79mlC5/VMHdypfEXCwEhVdAtSQ
QXfdb7Od+zx+nV8Bp5yc9PSgZlPmVlTeywnk2NFeYNDIcLxRd7WdYiKkAXS8OfSt
l4FG9I08lowW4m6WXFIYhHZ6/bbzeC7b67GLqpDSY54=
`protect END_PROTECTED
