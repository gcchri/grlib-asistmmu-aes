`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/eyi6jOE4Jyvr5zvhelviu889dx2HBgw0+UgTr05kFd7Ifk3mlxq4Xt2wUo4W6We
GtSOtPWUobUhhEUWYBhGed+70Si8liQzpk5BN6eMw2OquI+OvArN01aECFU8R7JH
iorg8h29g1ZmpATE1TXkw61eno/OhlZKWY/h2P2lEdDUxrmTjCb0cM9CZi/RRw9K
zhlGfowuMPrk589Vr++KYqBku3X/lY9xpvLFPDqDhZk3l6sS5hYGwI7/dRBiCU+Q
gD2fLi5MpO/iMBAL9YATu5Do2d73/Sy3c3EjkRWS6q2n0QDWhVM492bgr+OrorRc
KIh+uoqr+QOwzGRwAvRlsBpENbyTjfEURJaTcbo2/l+qhDgWZCM9dtF46b5QvURE
kShP+urMXQOBLF4tdzgZ4K5USw4Tohn8Z1WSEV9PEqA=
`protect END_PROTECTED
