`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lEXInRLG7StSxddj0qTtPLF27B6AsVc3rjeRLWjffNlJMGUCdzKNa6looFQhnt2A
XVWl/j/eCcKkXIUkKMFa8XUKW4Vdy0mshbD9WRCooyKV5Cn8JSKvOjCFwbtf0rU0
0FKdR1cgh30//g3bud5yLQli/HyftrmfJre+56TK/SBCICq1N5F4sG8IN/WKxW8y
hQE57MKNd/bAbR08hBpaFeLN8QaBaBfCond9p/P3zELwe6cIvey9qSICtXjFseli
e+oH9NS6LDQmLM9rhx1tIcaxPmhuhmtlwRmMOVVjesVejXCepIiedYrnfRcywBvm
`protect END_PROTECTED
