`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TgTsiTJQ3V7nO8VKA58D4LDh+Mn72Tbk3ll+ASyjyBQKUvv3bcH1uYFI0RuiFljH
eDPvAEEbWajtVdkrQopitbd1Aa9mSN6Ld5Qnl6flGBa+yLCOqekfyf6S3bkabQkl
Wph48SsXGBmgJwPtmmiV9gAGbYHlNI8Ets+p9PznASNK9QywnD3R5GSTCx2wl/83
K16AXCabg1rL96bsRXboYTxzJ5vMLQpiYpNLKHapKEpG8r/VqXI7U5tvCBqOoDfB
8mBk+YgBCqryPcp4zSj9ue2Uj+tl7Jomm2LaWO/s1lRSi+CCvs5hUkCYfQTEY242
OjbhP/z/B4GIJWMLaopgLPhxQ28pxUFfu7xdsvWnxiy8Lt6AD+qW8obh7s3YKDq+
Nez5tigEuOAI3tnBSCcRf80oq1clQOZWGSF8ihR2jB/04QrHTrFcd9PoKHCp4MmL
YN0ZkPmZ3lTxU8Q2wRQqXbSXEWCD0p52ILKze5qkz5QNVSGNbC0x7WyZCAKNmSeT
vzB202UyYrvj6eHL91hgvZdLTIb62ONJuHoVXPlvGMVX4QS50n41/VrKY0xice4C
RJcm2tdDvQPryxaECAFX9QSiDmKT+mZ4q+QvNSx7x86fUFn6h4bLB1mnBJtqGGRH
ffQVc+F0sU2REHViwTwkg1IT19K+zjuoFe3esjVqKTb8wU4rbrzI82FJjDCOdmFf
sc7STOEoigHndNwKP9YGuRPJuOcGExOAQscuxAkuN97zXnwT1SiuXV/RiOiUXkCt
MuzkRSOI61WW2DM2G5q2ehVnGTbRetcBxuTlSpyROewA9Efys+34UW9bMpJKTT2j
ioaL3o83DbiQnb9TRMgL3COeaGkOchR3Pk/A8h7xF6jfnZ4UIxZGB1hvG4b0oBYG
7KMBFDJf/iDjEF9jYwL7wpHHx9Hxap6mFqK/63oCcGmOC73MAb6AQ/EMwxFKhIsu
ZuLHQbksq9B19f/6xhZwOpXKTlfGO5tG3dcvu40d0nrjZ+kUJBWXn2EoeVKRbE1L
rJ/KhUUiGO9fg/n7CIjnmjkQnnYKGyoE4UgfwcYdkAXzDfciO17lUiGA2CNqOlwL
KnHythMjFgOv41EOWjb80SynDamcrb3+zbMkw2NUPx6Ds6s4r9sPedvOt3XeqS/V
t7+KIm/uGYOQ2FJl7DAjsF0WbOxLCfZYPM8YzLVGoNjDx9QRQ4aED0hLU+oxiyfI
D4GAO9p3aDO2zKO1itAlcAT87oiJXh1YZgHwXyHxgq6hETy7J7U1W+VVBvJt7FTm
sX5zh5dv0Qvs69JnnCeleyZAiYKfNVUirJiNZxiSIc1bGTT8EIVoZC9vAmjl5C8j
MnomSFwa26Wy6jr3NO3HQNdkZ5GYC9Q0t2L8611SR09KWVrXaRQVCGJbLEDjSxoo
BFqjD1Sw1P2lu+VgogjUUVaMOR0dh3naD4OHnORHIeSY9HtvCcild/goYwwJu5zt
a+sDwj2prgNpGLpMVoE/oNQzHtJbJlWESLtn6OKvDE4iieoaE4iMPsuZkpf1khPX
PgUnukgMDPOmNiCdLl9RSyjFcmFfzOVZd6PcZxX+sgTYluvW8j0yWEiDO+HErnV2
h0xOZCkoPey5UdrLE8+YkabD88orLFfoZ9u7AvzgH/uOz+iYoCKTroXu5eAeH+mK
bidx5GGu7+1Cv/A9enPcz49H0sn9h+QsGy4V+OQU3WG7uj8n1EQO2/vHyuu+u2nz
TGYEvEahnO/KJsCWsClPIR7/do6sy6tH44eauHajCoANt5E5+5oJqi3ttT+1/Viq
nobHa2jH3kKeWmFwBYdrr9AgggiHEuKokiHg4Nv2RG17fZu13REvPA6o3gg6IoCI
FP+CMuY162gkOagSUHfQpmJkSKSst8RYacd+HUdzFOqGFb+iHrnZWrARZr3XNjK1
Qx+F6c7gDAmpu+Jyz7ky03a0l60xe19hhUWZoPrCKEuswRMSnbX6REsE+B1SIV4z
kN81VlqBxoVotez22YopJmZXr76EJQpXDtNkZSYePZSmjSF7mLJ1qyzVTsLgJLRF
s/79cT4K/Pf/7oHqSM7jt91autRyWE/A/obvUlt5hSjOe6Pa0sO758H9q4/gsNsr
/QXga/+2UiaJ1vJYBf3RLL3SUvvm/lgzof/5i6QYDdD0u84Ni1PobZ8ITF0ofw+Z
sfrIHW7VfuVxV1FdpD5w7pX6yqF6w+/t7CnGckQYRHtFlLXkQfqFsu2NQe4NjGOA
3H0JK1GDxquIcq/8XlzetEoSst7yIj1fktX7YlX+M1qWZ+2mFJLKAtdOv/rlQxWR
E+Qw8CiRDDk6SY3AkFx42DlqS6IZkPLB6g7y+AEOFM3agSEpbb8ehFb2suwSqnnO
7W/IKs4gYugHCx5haKmoiVq9JpLfvOUaZB8hoPmQXQcKObx7nZQAaCG3v1CiIVYs
ACiC58oR2KwPcs+mrb3bb47z495gdhxucHw78AbZxTbIBAMb5Kl/WLYO+/fwV1pR
A9qb4g02CEwG28G/Znn9a5OjAoYlobZGpmAHCVGtzjgFuTV+gNxt+kCF63J8V8sj
dQmhoK6PvtIFontGl2cRFzLnYn9YV4FnJcSG7JY9nquqLSUKrsK0DFJAz7+nCcNz
rIpaEePYFL71UoBH+kgcvcgFHNx3oL1uVePjQZ7KT11jAwOdqnoSE/xL/yFlJT0n
Wfb81xbsamtF/wbCm4tXv/FA1+oHFI1oYIGtYlND4ym2IBk8o3uRwntjT0NZwO6O
4c50jnJPBvr2OV7Co43ta5l1zuTdlJbD/ghYNLXJbyQKvlnEFR7uVaH1QWFCi+EC
rIK9K8tPmMGUOJZ7hQZtKkWyemye9lfsQfqZgC/KHCB83onAr+q1FMxXEzDffLWO
JFWmzAwhAjSkXkan56rf8Pwl7ypeSpmiaKS+Nh+5/G3KAsJPR9jm3d0MJlJEjPXy
rP8xjkhKJWqyrO+8wFCXUWVax3dVuUzBTwQJlJdPOPrfQYGHnyfoH+RzwclU4lyC
3kGlwyVVXBHUMg2s6LRNxY8SXKYQz28h/ia/JSXUU7iS8due6HOulp7LHRbeG2j9
2P6EhXcei5WFL5bKhE1WoAV3Z8+t7S5r9Fok0K3Eyu0gqHe6KGboFvukmzbQ/GLG
SZCr0nyuUhFDJ8rdY2s9Pdc3MS4FCHlp97E/6XwcSowoVwkerPyhnGNaEFJJwJ4U
zFLCG4jHHlE5CsxTZSQs7Q1l8o3X9YKn/BEkSiTU/gGuU1nlTYQflf0T0SaeVEQE
0DF33iJBX3MWGOTAqRuHxrmG+hnPqbw4WSymNd+Sdkfzl4MVq04RZQac//ycCFKu
lveMidqUAS9q02u0XjzLfH8ZNfbevD5NFMHk1IRec+heyA9ZDljJi/suOn2iGX9K
8ZLvRiD1Es+lhFget6jrFmanAiJ6CdTNEyUJPldlBhVDExFD12RzN9M+njBCty2e
U3sS4VQlmnjQvGpfTz3NrQi4iNT/WL/WzTX2+k7R9ehRdZfGDLP3SFuc6w27/ULz
X0BVk9MjF+b6EHT3LXo7aK5hjqJj/3jG2y2Hj3+1coGxLC9mPCpAZStd1khjnR+3
UAtszkenhX12Ozj9P60qlj+gX48U2neRoRoRICxeeVAtYKRjPceLN/61HmJv6doM
aac2edRZ3u636UpNW6hrSlUxMl+fJZDDkO7GaOwdWIVJSWXyj7vRMyc35vkY1kIf
yyvl5wlqlVdUk7iXE4FTdpjxjtPm0dghvnTmcXgoVJqEFXhOrfhQHa+NcrF4YGNt
TLpBET+3H8Jc9aK0s2uSc+dB8UTbo0q2JYBCcvXMWBrRgWfa4Ph1I+Xmi9YvSyTQ
b/OVER5Aw3M3PpwIxWGxDGHoi5xHT4pnIp8TY8r8qp35tFgG5XJ9fKA4JMwOFCVU
+mI88AL1c8YTub8oPsDWgQ==
`protect END_PROTECTED
