`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vLxWRFJCiZZlpSTPFHUF2xrMQ1J7jQs5CDzfub3QGkfEgLq7XAoh03kFG6OKYG9k
ztz8zo+U0wU8uFAyLw7Qiwa9kpi7uTfn4GqPTX1OeJlrvHjoCQFf4/lhPfXNH1fk
x+4dyqKydTN7C8KOebgZ6uTbAuWmYsBRPkcIg2zWwqC60RqzYLejyBfIfAYiBLgI
Uodu7DPZzg9ObjP2igLSqq8fHIcYLnxUq5/KjaudS94cNcJramcoVuMkwm2Roe/k
bazPJnpOkWCcDujQZOSoQ2SZRpFCIb8B1s8wiJc5EGuuprN5LonKptApwm61+4ZK
hBIsk6klNiGQ3WADj7MDniRBXaFFQehblLvLfqFIrqw5lDQXY2nqtFdfRT920+zz
pJHJD9a1Ep+xrEpzJU7yWDjd2/BiURKqa1hpPMTrjlV1smopbyzDjd6PV+U38gub
aLJOWz+loIYU+dMXQ/y+FQ==
`protect END_PROTECTED
