`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vuR5oUwkRa/OKDqz7/dziQEIP/iwa0Uu/K1VuPA3SJcUFfGGMYYE9du0AyUfsQ0b
ZxbBwD16ROkzTCikW+8T7HR6gxQff962/R7HBLlC8sdrF6g/YATtzaJR6TdrwBTn
9CaWgHFHN7XM+MMZU/qrJCF+LJ69gg6dGDY10H8U5dX/2dbfkBNbq53CL0lT4kS3
TqQF5tWroBb9lpKvyVIVTj4xBJC4NSGlb5lEd2oD27cS7VUkW9Hj+c8XS2eoFMY2
BF/I+mR7sNHURqGEPrk9m/PJ9sbeydmca4GOQHe2z6wfA8McCfAFU7qPC/C3IzFM
k+UeiBtOB2yqnHUiDARGEKxYeXCAKrTTylKr9WSSr3s0jJGVV9147zYenHaYiXou
t/P4zvRrSGCSBJzwQHrDASkc4pXRVo1weKY2gAxdUbbsHedmWjmxshc1uI18hq2w
R6M392pluwB+26gxwTCkRxKmxXzZvoncJNqQha5dn7D2USHB9FFs08Qu6KGxmO3L
+s6yX2BJpAuwMkRWUsi64jPIhLC8nFQA0nDNqhPrhMRio90c+XWDWjCVxAXNTnlN
+0xBMRddZlNveSQ+AppakAHCh5+vqyi3Zvrp8zLIvfKP51ufPOnpBbApG2v26TLt
GjufwKWguobgp4CJTYY/I3rGA1tOkKvxnDwDUhrsMyUF7vDncS9FTJvWZSIbMYVp
192TPUcK790iRCpGFcnCaDCoc2SJ3go8eZBCS7tz4LSA4PawVh8pPfBS62dcdhWO
ZnXQPNZ/SRPrNUrPV/gkeS+uysPLCxwZH4OORBjNsbl0F/SPRA4XCbHsR87CkCuI
GIktGJL6Yo2Wi0WHL7o/KHQ1F8SGQsGSqq9/ZxI2MwC6pYdUqSP1qyGFDkd4e4X3
rJZzhnIrMiUIF80xj7As36e0ZCqioF7WYfQsMkTf1WPVPC3dKEJkkRhXAnFQlZa3
zFZBPgRjqQ02QPOZQ6UOF2YcSl2MhhkYoT8WMCPT9YM9yHkmylYAAe0fXQOJjBPL
zu6q2/3kZl4zkvVU3PNp5sjYaEfYFzv9DJ3NxZLymrWBfdSjpnj0LvLGyzN78Pg4
EX8q3LWIvG/NgaSzy9A+eAcSVxpioCEkcgY2G8RlOXiGDngGlWDpdC4if6Q98xuc
w+tT4dFlT2J+XIpalMBa4tna+h3qqYBSurvzuz29AcrgRwn5kwCg0/9aSWZUVigN
q0ncZVHVYmSfirUcK+PIIPRIvcjl0pc8KwFC+cxlWmpgu0ZBWWHBI5pq7VlvI9eE
1pWi3bVg/tboMZpjzXvP+3VKT+oTVCKJ2hLt2e3nRGVAo3bkjYeSY9UOWlBmiR0r
Pzx/8dDzUpidyj/29igVTWtDUoFPnSc0ysJvFha8I8L8KQc0qq2l/ioiZYzDDR1r
Dwh2+VCR46N7az4PX23VaELJxcIdYW81uvRFfH2cciHF+hZryrjV2Ha1g2DtnXe2
l7sOIl1EnLOymH7DhG7NSKtKjhqKRQix0nmBevxLeD5Z0kcSIhoiu6WTNntzwczn
oL90fFHb69xDoiWa5aWexbgZOxB5gmqPBUXLNiMs+kPERKtmOJfXheUttycxyb0d
ZcnYj+OZEY27MtxaJOj8kguXLh5DfUIDHL40hE72jeIAg76hbjlcd63UHbQaZ9QX
a3LvA7Fnw1Pvmlw/0M705/q2bcY/WNDEKCMruFh/b1ghpg2FLiFGoHsXqenZPr9q
W4eRgnhK7uVG8JjZc8lOjjrT38Yhdbg28SeOrLqXumNQF9rHkaj+5v2laGDn9O3N
fjSstQjy4WoovGGJIclX+OgQ0GGZv0Jje2gyQNTKi8BTqYlF7j6JWsnJeeVEiy20
m1Msjz6BkG0tLoqLUJazZrxIzxVRIvssL7YWHnWUkzX4lBoCtq8IZIeF0S0Y9T6s
kvuF6LCFbbDBb7DZoOUrS+78VSBm0ECALlN/LG5J/LXy03efqJ+/5UZ8jP6DmKf8
Z7r1Vme0nXYnZUTna+FCRAn4jFQIBS5VH1cHcotSmZYNF6IGf/gISEUhzT88rv0Z
TzpkrsuD1G2bH2aKq8NgrnfEVCTxXOujD8AFmK4vwLKlWfb6SSG2/BI5aBE1Cy74
Z31EVEbMWqjpPqpBTS2SMtpLQWUsJ9VFfOEiLCrzQTJLC2P2tnQf3yUTL2Vr3jLa
temRF5a3QxP6hE5wgsxrKFbnXy539y1/hdGvh6ZBHOQcJJMuMFuypVbHi54Gbk8B
N8SpXNDwGL3JzkaJJ352WNFvrCzgT0wg5ougTIYEGkwj41VaJ321aj0OjPkkb2WP
//OLoyT1YSqclopulwXs4pXnPoUTCXFfVt9MlQ4e2YLmRoU/WeyWMXrDfVSZie/C
L3dFYzsyBnYzyZZt7fQgvXKZuky13M9rvsSSR0Onx/eWNI6xrBHKisopImhsHKqw
cJZMGwbJyjKoGY4Wxx/vJj8DbrszmakrTatdMGBzxAM0pWjkgDuA5y0AYF6nrA+g
c2Bad3mW4Z05M/DpXOtCl28aNeSewojfVm8d8GEQUlVDfmh494L9mldnQkavDudJ
t0J0iDq8FaevOXKuIByaFZFvS2OQbwW49VkEt569zAYHnNYxalUBdMbUD3sQqgpD
QIR/UmZKPfdDPoaZrKJgYM5MNBY9yuYsyDhN/XX2cPFJx6QEY1uJE73aG7/sxH8u
qnBPW54zaCn3YSiEn2p9T1Js+oKzfU82ANqmg+vtQ/KjbBQzBJTFQPdOsWQD75sr
B9M2GcJ6QlgGn41K2ZDJbGzawmkLxyRND30apl3ozuajyCsMGB06NjhpD41fZLp2
e5dz5oZ9H4/RXRvfKlEh2CBR+fCGEy0EdL640K/XZlS+nxQn3D8qut1Yh5eNzme0
vzl0P1llgoqC6TGXvS4MZyzWj1tUG8AnS7OwhNJIEwLIaJjpDvE+VIO+btvOxRKz
aafSOv5ewWvKVkcy+Urp7kY5o5JyUlM9fSACe3+fgTmVaC9Dea92LVFZKkX9pYA5
R3b9w/9wIymb05ZNNmnumU2c3LZ0+177LmOnVR85ZXpkn/Z/A4HaIZy0A7SCjHjE
JKTryhu8ONfkzIsmah6k8oOf7nr1DwTpaTGr1erE7kxNkbUsU/vsYNQD5s1TrlOX
BOgyYfyXSipXdqJzSjsLsRucN5m42yCcN2psCzKZW5uNZ9XfC0NAQ8guHwHtLUN9
2RQInmFEKG7nqMYXAg/HvL6JsfzNdZcdcR/zIdn8QmABLID0dnNPh3pcrBt8i6BR
UP4duoXsskzW2y2AEiNq+dF6WH8H5brydIkvVRtfjj46geaGiijnYzeU1OZqrk9Q
aJ9dUehiSF90o1hfnHB5dNjZ+cAc5VFEDB+u0j1O5rcUKI4AyP1cavl0fw2yd5lh
GJpE4J5r4VBT1tNBgFJXM690X+BYxPTqqefkjjsy29/S3hipBFM2+Jz+2ceUJT0+
Hh2gHoBAERwL108Bc4kPHmfczVOPZ5ZoFwcG5hyto5vXGUIvW9H2ZDpjjqlrwe1A
BkTP/sfg0N7DyhHM+F7AmX4/xWRt9SX+G//QRGNI7+S9EmQpihJfDWWo2BmI1iqb
`protect END_PROTECTED
