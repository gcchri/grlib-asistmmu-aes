`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MRtuOupitiYJUyhCfifMxJSffl373V4RRogtuAOB4BcLZqYcI/aGfLZHclD+VFv0
Gt5HVGEPzJKNbJ25I4DwtbBxNlzt2gU5kNeX3IxrvdUQrLHOq/scA4AoxvC8YUw6
4kpfEx0wqrgIy6bccIt4RcahQr6qyUwMXMzQfVJSSDyK1vKUZQVXKjLoP42veowa
VwbUxXOh+hR344HJ+EODu596/ZKrHhysiCuEbv/Z67unXxt9zQYLHQrTQ+W10b+t
C63xjecvAuOeRHMBTwbv8sXI7/06PzCogA0Yud4y6AulV9ApKvbtpsKN42QirUxo
do5wNG0quuH8rsmWLV+qT0N45Ay8ArnKB+kNsmnH5a65b5jMYs1yRkLYb+SubYGv
LWsQnRhcBXGTPeF9FZFi4A==
`protect END_PROTECTED
