`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FT0Xq75q3N89eVSvyau6ENJDYPrCbxU5vByG+H9S/Mro9jrdHiG0nB7rDuPSm6ex
bZL3dr+zZbXlyKoAKSNDaxajqCGdUbeRDhm8LaCGN2ZTZIZ0a/aebm/CfNHqLozs
EguzUDWwzwsLWcc/SErLpczSxizaUaOcs4zTK5MQOpuXrx9jUvJ/O0bknP1bynom
zrH4bEvnNCXTGGIlo2IyU4odgpU8AUVs6lkKgbg68QfICwHEdeJIlo102q70nd+N
52TPNBTqzCOtuSLmDtkaB0eMfUpEzMIEcOhXC6EUld0o+ZlipL/mXD9FV+PHX7Sc
cZLP6SNAhEIoboyB7ZA+ygNT+dLXTv/0Ii2nCgFWtccy8jsi+WglBoxSJe45IAR4
P/5uzy2eUNowvUOtjFS/IiLkDXAkOOiydFWe9SvUpmrLS8Spd68UJukQB2NThcdS
VkVQlSUc/nuZ4J+BDrB6fqKjmT0ixy56WHK3dbq9DnXsVa4yKrRe7ji9wquddwgE
ZqhIsSqZdEyxS13y3a6FkX0mJBBU4AmLCZbydO1ZHoNXqb+pII84kXeFJuv1Kt33
cMWG9JYtHpWQge1zGnuv2TZ9Tw8LMjSuWA+jd1oneqtnR3DAZ0Gb9k2HHBxTP/mG
kxgKF6EUKIBNEfjrG2NgXIwzSSqcw6SvuFR/Re5Yg2EUKHHYwKSdfZPx2FjN1Uhf
+t1LVPEMnn2k1Hxs5vcWcr7JfT7BbnNjfPbVPf6KQKNvD+gheHhFIf4ql1uSufG6
rkbJYhYojhrRMc/wSjYaJRLOgBZFfCliNlwnOoGdWSpmNNFUMrSN60xvI5PQXSta
YbQmM3maaNhtzeOQIBkQEqSXyqjhw5e4Nie5jEvZu0mZeTPb6FMWB/GSs50zz/Lb
5JDYWbk7+QvDX24h2+4a1qkkLfaohtAPulGYwT6eiejSlaE55Bk8tpzEaN/WJX+P
TstBhRjnpA/ZIWh7fSWBVBc+lcIKSTKA+ghHxEJf2MuZ9VqqvsqElPVGfJ+dkFxw
kMVsOjMOYwscJvRB+ZrcPf8JkxUbkeSR566QHbkn5j/rSJRu176gqzIRxmQFgV4p
ox0UeeBG+HjUT/NcWKR2gc7yoZzn/HSjSCBsq/PURAmdVCSBseReWuFfKgDEbqWr
yAzcVunohAkMBZ2k64m215LGyQucusYFLGgs7xDZqQEn/agXKghFcTATV1paSyGx
xizLhN/xbS7N6pjQtm1C7Ure1vXaho82RI9dMdxWHnZjDOWr0dJiJuiBTaYIV4Dk
zrWkeOTxFmrZk3dS4hyONWp4FctS4Pfv5O3m2W2XI1oFShsWvpK6s0PwfL2KQigj
3pHCk2isHSa5CVZMDMazXx4gXxJYPFYBDX406rnSoW37wjB52WEsHjLVQ/f1jCLB
48ibRUKWsZ/OZo/qt/SIzOydZ5Jhk9Px0HioBuvDoslxLUMZ8XvwEqOOlyow8Yu3
G1TcIQz6k58RdM5n4t/bLr2MVn/1oGV1QZPRtAfXegedpO6Rq1o98SkLmP0Fsd6o
kP/fIEZXIr4ZaS4kmh+0opuc42SC26FtseLLq2zdJIP2rxq+RhasslUo+dztqyvX
L6UEh2wo08axjW4jjOYmfA5Fvnioe2r2rsBjCu/5aKokiPjwWTzYw7gj81tpVGa5
XYvpZvs46ql4g315Yx5ZoGnNNK8keLSDQ0j/hsdaELzZKczl8VWHFqscXwVLP/4+
`protect END_PROTECTED
