`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQlIDrdvHvBt+TyE2gION6fePiJ+GPiHbRckPJEDJZ3LpcFSNmJYqSFD4vGQl8CK
C8CyvqlqIRb+IbNvfz/olg2AckRkvL5s9RMPuTV92nT6SbuPTiC83sPpUURetJyH
EjEqHycMJENOsLAJ1HEd+1wWQDeUedqbUiJg5mbH0OGo2+TV5SjiN/cQTYW2Cq9j
clNa6SkGhkS2Jdfgxr8jTdMIxa/RE3323LyU4tdNEEGpbdddBufGVxsQRSZ7cznE
I8F3HEH/mXPmzjiUOqwHkj/K5rFSiE6IyasGTxWFt8HgaeIZjHMLOAbdk9bzrEw5
A0+rhClRFCXnEQdkbhVWrQ1HjbAYUr2w4/hk23uKLV88x2SWBsLJc+81WyjEcoLS
lq1UxTc4pbX1FUN2kkqlw9XGmazTwS1rdyMtfAN3E9MVduMAxjPUTfdEsrSeN9lY
17crgjZ/sh/p2jTjRCNZGqy5wjWmCrnRmBqvXomGnsBejYitJa6DXg7SgdYOEhIc
EGObRi8JPEhSHL78PdjoD+82IG/gRsDlVMYNmf9KLWuhwonUqsffSi67KN0vdA8O
iZO/ecgiexxkpwgaKlN9y10Mjms+k6VDKOSckIxost8=
`protect END_PROTECTED
