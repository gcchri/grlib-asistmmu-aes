`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+gEwYA7kKi0MrUwNX0Mv5S0wCM5rMXiPnfkaImCXk39OwqiEwnCmHBWp8piVDBu
gJxFMNecuwipKDLJ4fxdDpUs9vIDqu5lLAKEisNQdwjMFbD4QZGEPM8WVcTEIsh9
hevxBLwwZ52dm/stkE/f0hplGMQU6mg20sZnCscLqlIR49CU5yNrIVGeiv23WFHZ
epy7t00Q6FACO4DEFKoj7107d43i2+rkdUYOuDLbfIOFvLY3sOS2JMgKk1/Pel3V
VzhtMEyrUk0hsZEksp6LYAP2FtQoE74UU8Bm0GxkxNnLf3Blzo9EJPkFo2sE+CG6
FPc84aw408VV245Z+nWbR+moKlh7KBdGuznbLYOS7xwKOezukkMGegFPxVJDIunL
W2oX658qwcA8m1Kc9xIo8RhRj9SBXb1LnL3VQZDBS5HQYXTyJXx0/iTe/h9zW85A
9xhnyOgyYdSOAKFGmrwgE+mhLxU1UvjR5K6Byvh9qD20Y3ui9HyG5BHXHd6JSQ++
0NMqUvBZ4+DjrtMCngf1H0dX3fHcZ8DqEVAlFSXVrDlfHEz7ytUNtCLDF9B/aJqB
xr/DZkDCz1YxiXIvNwC72tHNd2wa2318rdpj7HJCzQQQxjxkPR1POs37pX8c8JU+
UaCVyaCAY7ZLHtk45yO6/ucF36KY8FAVlZDDveEEixuKaWGtRgZnS0A/U87i5b59
5rfHPBv8uKF8ahHP9UuTr5eb8KHg/775dFlDW3rsvsllipmf1O5isAfHo1OnjPRi
C49YKN12GIMmAK/CUJIjopBcYPBm3F1GgQkvnQGmka34CI/Mgfeq5ICCKfyI4tJE
l5w6oNjq7gfv9RWaxJeVu2+9gTkZzkATd++k54J7F2Z5aljd8QQVzfMo8LETFwtV
aUTWEkB50jzzyEk/p2Ocg1O/JKU7rSotyaM/nd4s0l6/d62pPxYOCSFwMmIUJe9G
STarJKAJ6yC0q+/aQgpIxXhVk3H+XU8M3z0P8ogSPf6Rz0qHdpEWaPsly9vEFXN0
V+A5ZC8GD4E5FdbJXRHRk6zug3W2n5r6f+zYGGACUvC9tZwsYzbWmxfb4fu5BRQC
a9Gf+yg8z2TVG41NmHSy8kaNtaoSdjS+p9zzr06dgqveDaE/SRt/A00mOE4HJuo9
Im8lE7yuNubGMASNySVmCbSU5D0heaXQVk33qleTYtzHGrITBMDhyQlLq3ixCku8
zwn5s/CJGreOTHkIEjZ95EXkQsobW6+J83rrbbizzvsXt+JXPzKp5Vktp+FlJOQb
4XYCnly6B8xkOVHxEmmeB8gtub9Fy5gWZeVw4bqCrkgQO2P26vebvS6+X2mdgjqi
xEHG3rTlzJD5VwXX8p5ToTTCdXVTRBNHUNvXdhVRHcOTXwUbsJ2LuYhmn5JBm0TO
fkCJgRCZPSlUoT//C/+s/BzvOS9m4sbDQVEZFouFcvWEnbZ472oe+ZdJMQdNbHlq
56EHfWrx3BlFQm/lxPsLjLvmRniV6tIYMjiZOIyb9tA2J0T47s27nIWPjk03ulO+
TJq9t5PgZqlCG1Is1P4lShW1/Vrj7HneQru/Ll2/udcFG7q02UCD9yu0sQhOtdVY
LbQpPScKQMOdvuZOUda73I6mdIpwlkeZExm8a4InetAVWW/DGJqXuYsbXLgQqs9I
nVGGWZm7uawudwA8gNdfwikcBnURvgOpdUm7frIeRJWgeROhzSo4PWLhoQGME2Hz
7j9f1FEOZmMj5K9T93JHTYd42nDug7RGct1CXPJX+DyR1KQRXSOy2JmbEhCiWVvF
TOfnRO7PX0gIe0uVaGVcv/vnKoht+vhpeMdkTYYy+XVF2PbZZXT7FAXOuDoUsU03
iEPpGrAtbeZTdmpgzaeROAkrPRTcA1MP5r+oiUjbNcWDuZiRRUp2BVFz33VkOExL
VrhrigAFBPlBeYk84X+KLdDu4tsAwI1+CnTZTDxKZ3hd9gRQpAXrVjXx1unZpRFn
PeHofKxm9upefD71VV7Fl8fiQGjt+xa5pZ+4uTYNdB+qAXQNKn41knOa84s4lggK
5hXu0L0HEIgflsNyGF1svOKgHCwe9bp2mBhvMoZscDXIgPWXgU8OkomsmBp5XT5X
d4LiKlQkIhEFSi7h8Az3GgLNZS/z/LvdofsDCguVVeaMrLgOPMcXkxyCRwZ7IdWu
4vd0zbiofFVSrPxf03zUFPSH3V5wAKlo91hQzB9Lu8YUWzurQyEK0nP9hmD0408V
r0O39JWUDnr0e4gf+cu2QInOemg382jvOefWpKWjw4usRj61c877Uj3gUPT1ZxAM
UnoTknzjLNPs+FrWymy/35oXtJv7G4sviDbIf8+sW33F6gqlV0uzXcmjNaBfC5Tn
EiWHR+0E/XzVINylgfQj94F77tfycuqwVZrbYK8exuVY7/b0FGUVIQSs4ba7Qs0w
NkxDHWVqkXnz2m9Xh9lFP2v6jEMk2j17rW/ao5/ZGVqJydDJ6onVJHtuiGN/Q19j
p9cLIxMu4Waw434LjOi05hEJQ7TSxCjZXwgxE9SWaEJIU5kTqD6LLk8Okspl6AF7
PfjBZL6k6w8ZXDcFmcYWsM5gntH5MJayXum+Excf3blXUoIhCD3QjhH70jTToF9H
0Ldgka68xJhY+XTtB49kTLzmzfi/kt3DARIjW4qXXPPveXxr4hjYWF7Gak152PMF
YpBZ7RqUf3MDxfQCuA5YXSfl6PH4X5qsGmPDXfgQDCRV7OvRbo89+w9/OeYXr+mS
ycF5IWm7mptLWqiHIE+2eyf6X2THZZj1nQ7yzhBNo0Wm1CPISozomQuG6qtrF9+K
XcolrqoME9lKu8gksitmO7GUyNJ8QM3zGOhnig5Zzbyn1SZWlP7kiSPKgTkEEocy
TuoN5N22EoLKOylruoVsDGtOG9QFq9YaSbCttp+f8Vdo4lX+s446wdD4X0dIgp1D
aDabp9iIqkWkyiciLSDwVeYvjR74N1kR1gb3lUYBrDBUwpQ8pnxpKL6sXZ6x4Iys
wwlgkxEhL26lH55lsI5RRLHUUuEYLX4++nGn31hLqjXEGXb6KFkX4EJZ/0mINHxU
41NVgBvsmhWrb7YdsNrUJ2T2x3qu3V3Pkqk/yT7sZQeQ/VV/aIczOknJAit5vL0T
yasjxAmb883V7jftn85DE2pMD1Xi+Epwki0Jmr50wM0tk3y4TjWQn5wuFFo5zw8c
+XO1UJLovIptqJi8awZMM5JPvEmdm4KNoUw98fxPqHKVM10HLHRmQZEJ82eEJu75
4uU5ZlmusqBZv8NGbAVnT+q8NZ5wbtUrHGcsfREIoPTYPltwT2cDi67mU4B+K5/p
Sys7iccEyGHz3C1zotQoIFRZlc06Gf9aCn/S7A9xeMgu7appg3ci9SoHjOG0D4ra
ZNkWR1lCufUEkyebdE8vXpuQxarwJ4xFE28nI1F+PpxG2aKlF7vDVIxdFSvm0nYm
Zxz8dK1jnLoL+YwaNpcf5woaWMMYi/2GbU/ByKQcxfIOWveEFvNMJhOIDa+oXXEc
QQk81d8g3WsgBrJt2o6n+gNJly/n+fn4JNZ+wZ31kNxxHsErWOqLv5fAeMfc3iwX
ln6zOuOwiSZHiikWQa0l2kOcCJJrt2T687TZeQzfMmo85wDzwZ5Fzt6Pl9YaxFJT
Jerd1d+wshdAVweaviwYgoH1ZG9c+gtGysPCSGvhbemFRpq9UFjjuwqZPCnK3s7c
w1hs+8XwOBQNTBKsgZeGwxLmiTl+fvnwHXN+Ihei8TcAgQLYtg4qk40324MBkNSc
IAce/jrHVPn0LJiGCfWHF1QVw7zkzpjv7X+GqE9K6AhM1cwe1CsZiHT4bIACbT7k
Ce65aP+8N7LSmKUrPhWIGxu5N5iKDSKk3wETexrjrkrIBHOPCj95UlYTVpmQ/Ja6
Lz+TzJ+v97yDqk0/nQVfhk/PCl7+6ozBmbr4/HwGZULNSQ597l6dvvq9eMglGneX
S9Moza6P04PL+uTbA/O3GFzgqIcQELzqpHdayiyRvwZ2YLJuHn11N7bU/59J4ne/
GqAJAKEcjaNutaLXmIhWdRsk7U7xyr/N5U5Hw41ygkDdzsQGmhT/onjcoNiojy69
vDOlAwF6+Dic8aJvjkEFBow3YhgB+3+9cwX7hCEXQpdHvNJaFFttnL36vHX1XbO8
ifQCCbuYXdhF4bMcfDqF7JC/eFBEvZkx/GqbbHWp75h/Kmm7p1GnMECp1etSt8bU
QtAEDgS3iUSpYTHJaOHciImh1ITN0a59UYeqbydBgaRE2MDtB7KFDCo3EUSU3vtE
`protect END_PROTECTED
