`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UjGxxGbvVmGVeEVbfqb6aKNie235Of3Dzf4ZTwA5Q4tLw0+KR3oNpkVNmVjnChae
ks/ySMU/UYyV5g4GT563YpV3il9UrSwfRKYHRwgW1Z1oJxG6M15X95fxQYPYlNDM
gBVRgtghR1hSauDpIKTb46CM6tj9Lua1xk+wLXH9aGC2sO7URJsBDOvvXlAbTVIl
VWLQQP4t+G6nhFKvj50m8WStjdkcpMHXmNoaSyIxWaJaCGmXxCprJIiJxDJWPMaE
kiDWl0E/EJdVHK/wxRb26A==
`protect END_PROTECTED
