`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lE1zygFJyVIPwSaAtOlEowiH1nQaz04/0qmPuGugDECcKfhUVeMJ7syV2ewj3rMq
USouJ/KoebhX+2lPYBHxa0f2XynBlx7JAXg1YWV9ndn/LAG8QVtJsCtMeBu0x7+p
NTRVKwVNPh8NPO5U0EQlCUFJQdVl6yg4vEnjZJSLvD7z3XvOmo1AXGQvcVQL0Z+/
hJ8C4DQJ6bOTCohrqHGz5BHVze3W17RJ4l6CHTqITrTqf17Lwb0M6nZ3OhfIXlJp
Jab4BhpCKG3SzUhCaGac4ZnbCxOoctfcZA4MCoUdfbmrFyV0Gik5j4a4mfqW6h4d
rSMOJqGxv4C5sUO+W5RIzVq0+X8HFRvOcOut/tQsBblVQaJLMthi/7nAtbYHrJdT
qYhyi+j1EDfz24spFFq2YUhCDy12TSJq/vogE58N8D5+wBQOZ6z0Fv8kwWPjAFrV
4vOzzmjHlPvFcPDBa3RFaN/1lcZtpFosJkuU8zYrpJM4jwzUlFDei0uz0p4WfX3O
8nDOLX5Csi5uHoU1ynbnNexydgxSBV6Rhykd2oICSs5UQz6WTjcGNBd+2bcoNhcB
ZH8WRdaaWVLPT9U2M5DkIjU9GKiY3q67NV/9kVwkqJYp4xfGAbyjeugdsqLMklOq
csmkN9ln65IAGBqa13kRtqdxKkcTFapx8DpqFkzWxBxR+Ujn2w4OguPz8WUy5gZv
XDuMdsx7qDLgV8BBAcFlINmrFkk0AqPt0Rgrd9CcohLhgeowIRgQcQVYqQY5cL04
KTHpIf+aRezlY/OicSQrBlGHohi6IoYWhYNsxaw94fIZ94IlvAe+NjfSQc76Oyz4
b8JS6+jx5GvcrFBvMucmf8i4yIpdC3FWgfuDh2cEs5D026TgkWeKwuBl/jiZD0DX
vKXibMlKTXSP0NzoK7rfC1a3yshAjXB1OHodsso4A1E8aZXnUDU1RVbfHi5W5mkw
AcV5QSBwJwuE0Nwv8zB9P27XkfZch5OvVhTrkoPMi1FYemxOTYBQH9NJfm9YM/H0
6ptM090aU+AjlG1gCzd1WhGE6la+DSkElBeFLkgVcHUSJnXG2jAxJkZkxXTJlElq
mUnLjw3zBUobYcJlQJh8PxrXXo/iqNZCfE4G7kXpKd8CHXmP6cBqCwPU+RePJC3x
kqJzpn0DH1AP1kU9VoeAZ//8atHO+/yIMDSsybxARBI/oxQtM0XGtI2OdaIufEEC
9Ndx9ZwQX7NhhS7yhxuE7iXw99RFRXsfUlgie8pPa420sMJRnG8IVIwgfW9HcuY+
mXlC9xq3LzzSlLWxGwBxYky3TWs6K5TYCxyhJbw4/VE4L/sWrqkee1HypvAX8VL2
sjgMma/tYbW+R9RGoybuRq34aGWZnxLKT/GVIoxD735zh5UjsjHFmZjGyzs7xuT/
q5Phn5OmMLEeB3DxETIkgt17jnTOlBo64ZPMIYxCA2wF2JuNamuEwI+lboGVE3id
AJdwAorgyBwLnuIgCJVAfzyzG8yhgn1qj9mFh5jWlF6lqwspEQdkTJF8o5wa2wCk
FBU3elu/BJFn4kz9r/7YgxXZfQuT7EIGLJxDuUKYM9KpzZJ849PQXs/H8v5HvELD
zybc9yAl1dmZMqSnLcEFNrcuezHP7HGjuXj4dNgO2inpG/xN9rlKIbpqsF1iaUQ6
1l9IAHGI/FGrV2QwW5sPiB1jvxRw2wj/2D9chjMMuCBjXcvw4FBfC2kFOJc60kun
EGgggthiA6iEMxLmEOyT1w==
`protect END_PROTECTED
