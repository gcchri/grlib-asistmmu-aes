`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r7oMvPB56BiaT3DsMED8LDrnU2iUWQu/993F9Xufr/2VJtb114Ui2iIAN1C6rwsX
tWY5Ajf/Q6hNWb3JmZXmlHIRnxqZ9reu1fUYOkMgTJn/oHD2wwvB1iHpxhJhVpCL
sbcWIdYivFBphkpDjgd5whCnLigu+NqefiE0t28ETcVCqVAMSL5Rc1Zt1ZDDRoAc
ESf0plga9S5dYSJYP8tpX/CXY3nuf9McXy+N8sE3vh4+Xeh6wcE0tpvItnxQmEuv
j8v3jJpLA0xOX9cd3gnq4uMWRjvDq2eFPIWRLpY9YyjmIIN9gdYblmzuVe4OcMLr
n8uaWoSohqc2cR+7sgPjqA==
`protect END_PROTECTED
