`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
btvk1ydQHrm4gdJ+ihTw7AvlwXq0vLoCb4RFSVx6M1ugjzehfMm0I7jmaEVFlc/T
leuha8hNuhJwhD/CO1NX0AegugLZi3BGJ+tBjGrMhKYjBilzUkV2/uDHqDXSAhmd
HeGWiJ0gVaNIUtU9nr05XJNCdcEc5l1oOkCzdFKWNjZ1vaVZJgmWKAdP83n9cOEh
9A+RB23RaLldWXfKDEkmxF5CqyQ/eR6yVw2jDVBlDbGNc2uRp5FvQtkq99QvsXzC
5clmIw3+avehuyhWSrQ3O4no0JLGPiLs2TznF82ir5sGC/6tQa3jerNoqn/YVCMV
8i78sUgUWEORxrX8nI8sx+K2IOceMN+q8mj6OBaYuBEJzxCUMUzsH1KoKFQWZDEP
JsxRqyQs7EBmdIk1+EvlV4XO/rl+944Rg85NUXXMkMuaz3XV6MNuIY+xPaHqRrGf
y+vKSiGY25IWpnFla/inrpTCyQRymvprGliwvnA3jyCQO2VoUGShX244udHP4v/d
5QZ1HItvtEaTOFF9+6n4yI+F4KVJVq2B/MM/JWLs8RSJfzyfA9MC81dBl5hbVmNF
0RPfLzydUmomp/AtVhMYTg==
`protect END_PROTECTED
