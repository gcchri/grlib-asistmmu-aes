`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
awtEy/6p73izFJWz4CUwhD3OpdItRq7x9kec2kasbFL9VIHXRmHQsauLihgV1L62
1KDcnkIGwueZHY8gZ5PIOt/AvE090dQR4gc5iawFuWqRcLHxyshoEP/tiZRCc3q3
pCvnDcikXcKdNAK4/5S3wQIGNQzmyzLI7y6jnszhTRApvVv4cJAa0Jn9ltrlkozG
fb4B/BUMJEqfcReq5Dj/IU+aM6beUuiLE/jc0wmTQwgYI120I59KaKDj2pOeKFyi
5nbGPqNKLf74qbQpLC82vQt386+cwn5KCGjmEZTOH97DI+X9UY4wFUpmu8cH2MMJ
fqcmtpi5KgSV9TZpCF5SrWM1DgbYQbwA9PsVRSU+GtjF7DkhDMYzQpr6LNyVAX1I
k3coIXLAWcJUX/83H8Dji9T1MoIPbbxB0XW2S0aAlFruLjkPIJK3YFWHXojINH/6
bkHC4yBbn+V+3gdI13b8PH+WtXe/vviPoxSii0pBE5kEij1cdYbbSx75brTPTtOr
v77fGoDpUKgPW9QKjTld94ItPZHhZ0nUp499Ep4v1Pk7OSATSrtRMOnQgS6yW2Fi
KlukL4y5d1kLw6lqDl4OCT6MN0c7lDKZCweBD9wuny8qMq0lazgnYcLdvPO1I3GA
tQyq3MaIvA4++qEQwpiZXCHH7gd8hvuUjuo7+flTZbZY8ftpV+3blyGSxN4DRX5i
5RsoZYnYpx65A3DftpCLbw==
`protect END_PROTECTED
