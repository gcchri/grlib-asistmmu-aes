`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xlwutipIcqEpT/kIi8uHls0ouxWN5unJM3u1SXwzSpZDyniViZhjjnHnpGEsGJiN
beR6EOW92bpTzArx06W+a2judElP3spdesGBCjftULUCu+XB7ErB1vWCca71nO0E
Xfd3Je0U5YipU7NvbZP2DmTp0LWWmSMHR6DcrWuL3Dr88Bzfuherhx2HhpbgCObl
yU/uL6ja+PRU/ZFZBo9yNzqBu90LrKZI3HpB7osQfrnjOqDjQ++eu6JHEU9cOvQ5
CYgrgiOpAznfWMPGIqZbjdEfWRRbb3l7RmfaKOnE1GapthFAG/auSTaGzAZ8SFLC
+Bw6u4+WcKxx+jGIudYYSPVsxquOnfLAEmku1vTZ/VLo553R0zWqQBVql/TD7fm9
XdtaQhA9ZSlC0eIIggIf+R4/nR565ncNfGyrGAtoxX71qCqxIyYuYiRN+D4hsDIx
fXChMgdgjaImkuMYXCkT3crc1Tmi7HzLIAXPZrVSzQ7Zn8vDdz/XlU71MJ6L7am/
G7xMbFxtGV1s/lv62MTEM4g9ca/cGSw1EVEDpGRf+oJjcKcPqHJt/mNVFXdhHRxW
S1LbOElOc18HaW8kj2KXL9UDfg/WjoWtstGni1UTOYDiLC1dUxTiZ8CfhC8ei2NN
dDqWFQxr4+8RUJqiki9rag==
`protect END_PROTECTED
