`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFWUzCUw0z9sGV3sgWDsWS5ylJajZNmWR6ORuSLrl1MDgaTVAQgZqiGYMVHjAHaR
7x4r9ikBkk4qiORe91G05NF+NsGzsUTGgtdWdGl7L964KeVYxnJDL2I+kypq0ILa
KtO/1pkEiWm47tWpLif4rvNZ6gduYYFFVaja6ujvBXnpaaNnHq1oP5eVdoPKI7Dq
J5jxEF+PdAQws6PY2FiJ/2+BMILMU1iJ0uLKs8Tk3fF4VrrdIXjbWYtWYoLoaJ83
7Q5EdD5MkgEuQ0zLDfnH//2n6Hjca+IwQDo8oo4pNZfNPbZ6WVywvzpXcPlpfikZ
a15qwijww2GXfgUK6HptXVsundQssVMJ0+VkR1RzykRyAaPVVDNUf7D691EysI55
egCin2BmOIcMD/rSSEH2+aY/VeMD3EMBZBqiiqfZi6/mOBMGBYNE37rvlUDAkUa+
MV0G7dF6EAGuwnP6EG/o6Zj60sJJWJ81cipigpYR4QhW0DKXaDcyj2MOlil50a+t
cogFgXbOv7BwPG/jylBIh8MSNgB4ni6iBKPJrGMZjumFZRntm4+71rpPfiMClbIf
Dd/zCEvSdlzwpjFqxCGesJQSPgi98E8PddE1hUqfcp+gL55bV1OPqNYB3MOsUmwD
6aCgeBDL6wJ9zD5kogf2F+IXZ3o4UlUIlWmvXmUFJjQBJqJSFrZtPQ+7ggb3pR+Y
nstLChFT3lpgmtBhwuAJtg==
`protect END_PROTECTED
