`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kkjv+CKXTLJ/PipkmTfYXa5ecmDSnbzLjAWMQdHo/bN46zEBaagcrJN53kf3ij2d
tIgsUFV+iva0LqxHija2Q1BDnGvxDNnYnemZrN3UFodOtn8jd5rwBJ8nKlZipQ4j
mPooOuUk1ByMORiGNtv+b7ferEfg1GxePwq9hXFgXL8OzblhznaHZiuhbUH01U0a
1eUqUCUtVl5YsOEWd+nzRUkwwVZD/clYW32NRAad7V1Mf995t0msCWXcsa3Iblv/
Vyh0R7ibOZnBNfovufocVDSo+c6EWpZMYLArHmMzx/wDruQTot8X/93BV575NhDh
shKrq6oMexAM4e5lUyqSk4NVnpeBei2mFXkQ9X4jfL1qtEnCiE82OlkeR9wTwCOv
yPR8aqZfUPqpQY6ntEH29ZcFTldJUbU5/WmGAaogWXpu7dCDFpCLjAVdDdsFAyAC
Cx+AXsl7Jo5wcD0hqnopz45FELC25aCQFvKzwdc1IuLsap0G6P/iZ1JwLGo3EbLU
ml+4qY3pdQuBlZ2RPXR+3b0F2Ypf2GaaekW+pLS0DXL3D9DPFlV0+NLfZ0rmQxeq
N1e20gzrVNu0aAX4Mj8Lx8pFx9OS2kXAwofjtL57omY=
`protect END_PROTECTED
