`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WvT6R129Sh23Zyk990213lQc41Dg9lsljJ0reLhXVE8YxpDkd5Bo+DOIOlkUh89i
gJPBbjCltKNsGttzlMpFsbvnGbcO6lx42lD2I/ixBMH0jwiOsxTPQF56ewWzdqDV
i1TFZ0cV/RcWFoXm6Kustpv/TUPQpTgNoFfzOldimgbardDBU6VY7y+M+uu4zSic
h/R2kS5Z+etI1x9PzX0TL/k5RQ07nIYXCJLSrh6UU3c7J4Gqrv33GmEVyTMp7ilq
nuL/CSR4RjGXnDEOQvDLUlB13IbAnGCeMKhj4bqAB1qzUyZbLD86scLszx/H7fCD
peN7CmMCyTA3NLy1B+UgYRaQ0/1F4LJ9cjWZg982HKVlk/miRV2bgfQHkC4yJUFz
MCJIYQQvgX65qxpNARBAZbLmZBth1EcpS3GxNNGsiP4=
`protect END_PROTECTED
