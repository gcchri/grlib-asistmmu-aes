`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NyOS/0s2u27vQN8z5Ywp0RogoF5b3Me8RmhE26ChthgKbTvqejgN1/nJqSR94Gyw
NYbxqFsl1zgR4EdiPVJYJKEZMrit834x7lAUrFyNm7PzR/pUROej6oTt6xRsg6E3
DzH9zXmch3epLZul8ahjs18Vm0m4CSf8b1mg8ictRX1vSjzpB4PNc0VAr/GVGiyr
r7FvzvB3s3iIdnQWA2elJqccZxPb4mP0Ekb2Pa6FpFjPmx6Sgl9XLnhAnHPc/NP7
ja87RMed9JRfn0imE0RJPlhbxAQW0b7my14asqOyqJCBBlM15rhtSgclhoG7KunB
PtfkUhTxfeCS4la45NojdCRsQiL67esqpEy6F+sv8j8tVapAttRHTyUbfp3qY+7B
wNQGP4YafwwhPyPK7V7ijCSLU1YeT5ukROgerYfEQpR3Hn1uDuzZTwLRBYlS+He1
SgP7R9OPfClGHTC+DK2Tekwn/OSA+ZJDHaIP3Dp1VKG2Do52I9uQOSxHoNc9VTWj
5BBfqiOGPYDVjHdXKZLrLGkZd33HROuh3p9CEyuNnzWlkF+OLW3/NtUd+vL/jEfC
h5URX+WOsq4JAp95YLVkeheIIqQFAvhBt90H6dDvxc6kQCBToQmER/iN5DseNyu9
X4dNi/ukbun+/wg5zpOYyA==
`protect END_PROTECTED
