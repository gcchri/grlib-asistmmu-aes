`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOIZ2QQ8zFo2xcE+duRVX+LkiuDCX0IM+q1w0ic/IqGT76ff0HtipW4Jw9PsK1qV
2gX0vNQFJy3dlMprTKvZGEgvsm2WJ4Ae9ccFqewgE+I3oqzP7wW+9nK63zvTPdZm
RPKKhaCDZ+2oZCZTkQK/HOaI4W2QRK1EPKftdvcLCWy/48BvBGuil6HcaLgZ4R1I
tZPZWb1fef3Yo3pPY1r5QtuRKtPZ2JXXZWAavvHpbB7HnJeUUhpzdk1ZbOlH7+uT
qWTyMIHFO0JbXCLOR1p4cjtAsZPD30f9HaZZGPwSfPlf9sIITJS5EVi1/cuKiHhy
Hk9CTmQnR+f812RvBWcBoNhDLx98WF/a7nbi6c9nLEtydbgwTBaKkkYqb2p9nhkO
hYj17rqD1Od4GyVNd8rSVCZgRAGfNV4acRHb3UOt3+ouIFIUS2R199QEpl4yIY4R
g1lqgDPg+dQzCIAKgGO+3tPJ7gCiAYroUD3Ny3BtLE41laAY9qc8M31jzjaErn7c
Th+nni/Ub4SCt/VLMIZC0hHkq8an7r5g+zEAvkqZ9AIkMK4jZ2ztO5bK+K3KfdTw
Sz0sgFJktKvQNtnzZcuwkVoUzt4at6avUzgg2JSbw1D31yrJyIOVm0e0FMBlrAIQ
Nizf+27rLt+91+JX6h1yj243+aRQOewuMQjkqBOw2lsneNMMFZqS7646Jbw/3Qyh
pHXCBiDFbaw5/Lnu/9aifi0HGeVo5U3r+LhP8g05Y/ve23MvVCyYo00kdecrK31H
3EKaX6wpVspR2DX6Wj+EGOJ3OanutxiNnOoIT6lMTAozwXyQtmhtWeV0gsQrpnLI
TZWdREF9jMmNlt6uTjji++tipg+d5HImpFxOgoK2gV4QWd+HEZQWDHxxINykch6V
SvEsOERAafkbfMJ30qppol0MkHrhzhqL5BFfk/l3nb48IiauEYJgiy4k9u/eBmCQ
RVxzz19gvZOgD7Pm5wWBWlV0k3Mi9lyCanFWuZXrZ/hRuWfcINEgpMAK80zAE69L
VTg+sO6Iyet3YDoKspBjcAm93oble5aw7j0xNuGX0gi9SHYvffBCQmPjoCWfNTum
S4rRhaZlfLzoMc9saAqe+VtqayUrTFogQZ4NS/YF2OR3eQ++4eQDJGOwCKPW4ipg
mwW4/1dTPVyzq6kxqXmDQ7MwS/l9M2qqk0oP3t45QXjN7h9rGA4asg0ZVq/ZW8tB
12vGrfyPR+sWaNJyvSuPkaBs7PZOPvAEYe+StSkePIXHuOyJ1qCE6pDVKbRmx2dE
`protect END_PROTECTED
