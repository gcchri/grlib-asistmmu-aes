`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aZ/n6ECi77owXwcHUfVVEXLNaG2PIVJQ/ugYpTl32LhBB/wuz4HELKVKVgYKEDXj
ObJN1p0qhYLXQDgjq6riCdSUeebJ/gWw2J9d7ECshJTniEJ6MzIpxeSsTdLifAjU
24al+BktrTFW7TrNhzyZe85CmXrQL+z0Iz7SjTR52R5P5vi81xVHZ31o2cfiBpAW
5NpzRI3iFrj5BYRXZ7KOPSE+/4gLAeTurQYPe6Toi0WbCVNiR+nD/o7c1Tao7eIH
Ob7gaX+bO1g2QVWh3Ff5S9K+zt2kd0YXmTt0YoW6GIVrw/+YXArHxqod1iECDogs
RWEw6bfWcw3YwxjAMJIWIBCqdHSEjH65anWHJDvim7C66bvnjx4Cq5KCcXwOAzBz
MNQdiMHSKpMfP6GWWpVGWexnUg6I1O9cNjWv1v8K1pMF+WrruCImDnwhmnSUyU7/
R2UysXOQRQDyg60BQDmYHOn3ZWAHWQtiDsrfx7TMStKvFfW/G1Y9zMBqDNXTh3jD
ec5PB5BI7iYArU/mah256Ql4EqkoawSvNGRmjb4zMtEulBr86HZa3ODqzkCjASrN
UmC0+4wYwlCm+WklQNV5aCvnqJwvYkByxlOP+dWVt9d2sbtn9XiYQcCYVRpX5Uat
Lij201PfcPQx7B8Y+nxLJEuHMwDa4LuBenHzci6FuCYjtohLCv/bSzEMgAF8YC2E
e00PzzjctHXg8rDNJ/q0FpKA7c1iZXOJg4UShoorRIMwmI7t3NVjy3iFrof/NErq
T3iBez4QOYmg9MqM661y8i8qtZgv2o1mcD9nxiJEEdLLNXBcXC6sBmdEjFemTtRc
jMh3oqcLPC1n2u/hA8kUYONcX0C706QR/HoCjD7vZ6Sx2TEgDJm7XNItCQb1zPGX
/eFppvS5PA/TgtjxdslTSL+BU4LYfZRaB7ntHOm2wxVhKijdqbuDtjoclI6xT/Yb
jIZVVw5O1XyrPzN9vUhcGtvkC4x1b9cJWRova/vDBIJWJ3Mxk0ogF2P0AOpdq5I5
RQTeWMdNgthADwG2PoLGz69pzvt7wDk1NYl/soWXNBYbbuC+TDvcNXqcLwTUFi9o
Ylgax+F5zwR/lIX75FmSUbRqiI7fm2fmNvIEejY3+g7toCQsiFnKchYqkLB7GeWE
GVl86WrusPnf0SPMFcM2z/MMXJl718V98mILi+lcoOhoTzjKB4aOLXu10VjjsfAa
sb8eiI9uLyf/rBqOKvqcIq2FuedfPfdHG20iK2C2LuY+gTlfyA4PhKOnW5V42FCa
`protect END_PROTECTED
