`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VY7B05DczvU/xjBpJ+KUkYNV/1PVf/KvVJWQ5xfWEKgvY4WHjvFt6qt7fCfSg7PA
cu4v3exnsw3lk2HauUi5Cvi0t0XApm0dBlja4v4AXObbiIC1IGexmskGomIPfjwy
R9ST84Zfb330Ea7yDqZKgkcAdHPEQJKMlTq8pznD1SjTCntmzTGk8VIuwue5OYVw
NiZus8EibQ/M5jiELxr/fulreCtwpobQTvdaekRyQO/tEyH5+cjY0/nYd3Mt09gn
5U7m0Ya4ebq8CJDwgRCiAXd/Ee0LKEBulMPzJ7OiddIcvO4AhI6wpZDXo2YMnkMx
XbTIamnaucX3DIki5+rdzwe698B7OAeQccJUlG0e5YdHPeIMo/6QPcejxPsEGpuE
tW03GCKAKEzOPwtNPnZcp4h4vyBawkVsbvEWZ8ephokypw03/i7k8yPFxD/M96uc
mmsY3D2xcUqa9c8ZxT8JcAI7m0bjRyDnovqBL84/CZW5klsGV7hoqxS02gNCR0xT
yC/K8fUn/obmPSkx4CfonuXxKTrSAZOmDfFkpfrorGTZA8E7xPQAwG2tO8eV7PFL
q7JQiQlIj8BBKOQJtpEOjZBrPhyviK79UyOHqL1D5CJQGrK6EzA7WB9p21M5DYN/
lr1toxayeoqLHw3pQIPuSgbROISzwVmasXUxkGXTtfIZci6PjxSfImj+3YMp3kNL
kS+7mhgxA7Uv4pUN8ziEIwa8xmvuI9EurLhSwUoKiwg=
`protect END_PROTECTED
