`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDxoPxYH6DR5L4cWcSJfqCzLK/2IBTvKyKO3D0wIlkbkxP9HupU6Ng6uKnKx7d47
KPt7egKeIrGlfDjAKnK+GmChE+FTOlQfLs94C29OhS6gsTR7eUugdkOWrIIDNpqc
wiEkwajfG9oH+ma9nj35MwoCWBiS1gg3fGQHkdnTzkpqtwh/jR7MDHzbyyTRjNHB
MaVVhGVYU43G4X9pbSSfElzPHgjPKJ9+zvpI4MVBKM79VWYrW5avpM1fF1KE7Ia1
WAYPKpHEwPv592xopq7wWd2dw0HmhtaZawl/lZYT3eX2EW8tGMV7asmkB8d38u+j
TimC5cVoW/w9IU+ao3zq1UuRm28lCpY6hRjVw0DAaXea3hy0G7n1JqxHN/aqJxpS
KHFNm82Z58SGzA6OnoVeFRFzGBLmscHhCeyEbY3FqiTUFak/lJ+dbFF7eTKv7DL6
uhUUs4lSTR6cbq4LPoz7RoJTlaEhFhUdeu+BppviCu3J1iwOzUVoXXIr4dxQhrnn
uA7fJZ7RcLAvsgdYFOe8afvKvJJzbkcT2ZKoWzoUG4ZstQ8Rtmu9MyAGHvsGxWwr
SHxxFErTwj9wZjxSzjFsBbXlgvaTr8fcd4XTjuyOtPa26QcEVWYOu/LjkLfMXcAn
B47V9aLRMMvIdhMMTdftmdPPj1bgBs182PoVCCjtNm0hSkdA9Es80LAlT3mHlcCr
B3Pg0WCRnQxay2veYelqJ570jNb01uurMbe2GL9Q5WEcFwamP/JmuNqyvH4ADe7O
5/4iWNv7BdavnvBPOOVyrzs3+o7CFxD7D4TlsREnwriP9qz4dOLBZZdGxCG8vG1x
ta9tBYy8/C53Jj6MOR5TvJg/R7LU/WEmSJNYawQDp5C2dNLjBEw1kDVPwua8+fX2
53o//6b4sfsab0l5eyrj3PaiwKfKLBKsYNOXq0CKt1Gw3EV5tH95BWdwBKHYoOTy
LL1JYoKNgzsF5mOvKHmqLSLfbQ50xbGMHlBvYM/cGYvMus/QO14gh8an7EOuEg+f
bQaMnoXAuljdghw5jsu2pOwXWw+DZbiuIUugHS36ABgygO5Z5e1ccu5M9A9p0uX1
sWcKcELU419X9lCbboRPhcO7fS86ppqronk/kabfXLjR2D600+RLDjPfIAtKBTES
OlONmRR65oH68gfRbr7MRhQTw5q5whuCMm0Ul/pjOsJ2g8kB5NmmSkSr9+mdSC5c
Fwy9DAC4D/2AfBY41OXxKxKmC6p5zvKGplIK/Utj5ToWf7NzZJOBnh48qLDuXepk
vfBDwol+Zj8IJFWw/P8qIo6IpxVTQ3vHdGzdcRu8bdFGcjjbd1AINPBSJ/JI7wcY
iNvvyLszo2kisyAcLbIzT4gqP+I7nYXGh9nod36rQqLkcHIrho5RjnaMisT9SAr5
r2CK9Gm1dCwelZoxdgBP07hnB3Jf6Vi95vzWVDjY87ls85qi8V73sjojg7doFYCc
vdHW2LpiyDDuLeL6OsBtccLcgfN59syD29QNJD2SpDjBWYXzZvZCEaGdj5UMP7T/
p9asQ0R2DXy9h1WHr3Tyog/IjXxMzMlFOv/zLqehMa1W2et9YYCWylxANzd9F+W9
+j5OX+VaamkEpY5HPKwvch8/Vrae80RalG9EUtX0mxulS89KpC35cQQxeQp7LixV
+rvbbU/IHlSvqwWtczA6XXhxK3LDEEqj8W/GEITy+G0MwhSVeTYPAv5oude7AbVr
x79otna7G7KEHHmFb9frvpgxf0Bwf8Yg+W1KSXjJzeHR5+oYYV1nzYVXdsT99/g5
FA7nF6ZbSXRSW7VZnsv+/4LyPU8Tm1KZ/6KvjcZfB2lqcB6NOxb7Fo4snHHn73LX
ui3liTHESKGxlj0aiDQeteS1QEW5j4jBtgXmMgNrYddVTcFJzcJgouchGVEN+Dsh
G9IK9mnsKy9y2yF0jbUho1zs4IvusDGIJhn4D8Oo6u7oubuBv3yYalcLthh3PguQ
AfN1LUaAbdVw02LiRdP2Wkeos+11auddPrmY5SEdX5qtLG1ah+HVyKNroEgfjSs9
Rk1XtUS3usCceDlb1haI3MXmAwMm0IRi+ewrjjCnL4W61FqS31qTzLLA2/Szxvhq
arW806/EEAbVyjYZlo5bb6IdfFWp93Nop4CGbpDSeL1N9CGaL/hU5Xzh8hi2RDbA
F4WVpNaYWtC11BxCDsoWJ95/l5F5DIBXTgDpgc+DWjur+u7Pk19H/UUs2Cu8B1iw
ayx0qfpBAmQr3d101Qie4tBkSx6Q+G/iuYXpw7KOr2ISFSthMh65aheeM1a+q7Q/
rJLVQuVUu9TkR+eAqR33sqxg5SaOFlN/lfZbXNXzsRMNWA7M0lo0v2GDVyKfJvFE
MdSQFlcWa7iLfK3kzlVmJs1ceGh/8uah0xJQZ7sUrOE2y+1XxFDp/2/uiGPVrMv+
FoRyhlq5nfeBH7NVmRSFcnk03RjwvoOpAicga+uUKi05ZpH7jMDq4rCql+7NldvP
nPbGVPqT7WW9z2gc0gnCiH/YILgXDDcXjr/AKtODyamtA/t3Wj0s0PJtqhAyLakN
0KUBQ/0TVTRR/3F39Hj+qmM36aIyVQcJMiwm9Xjzzp2sxk2krizhlA5acBVWTJZk
G+RChPsWaif19VLFW0VxC6Ch88qOEDidTvsr1I7GtaO5Sb9SFAMnIcYyJDaCHT7C
nYBIHtYo1YK436XCnO2MRWvWZW13aV37DdT3ZstLWkezHpoDIOaxhoL9fDANhAjS
t7djXaSs1gIjThIsLZSwhnaq8qb+NKOFgm3n/qOyhVU9DMf5gvdxiXBf2JtMyY1w
PM5Q8a0t+ZaAZlejtf2alPQddOM53pykdiE1UI7B25O3eIsdsFUbhFahlA6XKqgs
COvxrhggFIN6dVfD3WrB7i7Cn3rFOX1VH/dfnDokRB5u4KuruP91OuPVzdnE/HA7
MDvkJ3QP6aJLDdZ3aFifKt96Cc7qVurs5//PAZ2r1HiGTmk0HYU/o3nT2qRCVmS9
8hNhxEz3fPa6Rh8DUxLtMG7KEwnMpAwZPvNR/7gagtDvNdyJqG9UQQGOWi2Vlp11
t05o8SjAZt4+7/SFKYxujc4pIle8SwnRIz06jKjulaMbOYnkb28t4KaUA335JYRt
c2AULZm+6efodLjEMy6bpun8SnYWXH6RoQIWsyYFrjYq8zHkTvRPHGdbFtRIp1VF
s8kbSz/HwxJaocy03xBfQ1aeOwq2QauIZG+NmVGJ+yljs9sVMOYkIVZ71z7tcWVK
BT0NlM0sfRiv+Az99A1Qw3K+64xkzyBExVxM8g/1ed3h4HgOyoPNDG6yB9skIAkI
kv1wh329gXc5NmI+tjiZ9GeTil/h3kEi2FFUhYP3NdcgRL1uDDKPn3tN0hTZAvKQ
LWVbpjncQnVvjq1XDnQjlOPH2XfkbjmVDJEJ10G4VYPS0b5VWf3l0v2sju+ldKMd
v3fD5wUdJQbwATW69BjsknDeJTO7OgyZwKXSWsUELi7rhYhiabjjjmJIETwEJmQ+
1jYzYO9uhdQDlWAcT0r8lWzk6g5NCGd1Gsd0vjSjg3wz6oD3XifOA7HD7oU79Nz9
BjlNzRuO7UfLVvnsll3szdCzHUm6ek17w73UqmBpA4GZHBBZVbo6mMWr0WDyq6nx
bBq/fUROxKg26vW3Khoq2hFnwVMN5qDVPB4UgI1vh7NlYNi9Zi4kBtHpGr3oNNbY
TF1D0KMWxfWP0tIeSJUkQkpaJH1fsXUH9vYW0l3UlZqLrVOFm1bJbs6SRaGCrqZc
Kxd3iflru9gwnttv4/3IG/KZQcwhUoar5vFBiDHGrdfwH6Xb2RWDuzwxplgjwI8V
fYsHHKvIJSyOOHF2OngK5dp3t2pP6DYyvUj6S31MaKmQkRgcHA+oN6bK2CevG0Nk
i43GqM69ZOza31IEy+3wKHFefvVBeWc2tljC/PJGGAaQZyttXi8hj1uy+XapxGSR
MVrgBpKRI01nAXnpsvhmOxywxor1YSs+Lg+oKBh3cBGGXgYOLPzb+Od/NkatnugH
5+u/E2qeayQLGbdmuVpW3QfI9ODJVq5lT94D+w/mCsZhq5gNXTymtCMkqMM6JLdE
zUQBDPK+VSqVVzrrL0vSEUY4dbioWH7xi7TFHKetpCaDUH7keGhYplVqV6ePadeu
8zRD+aOIJksIerUxUVxxujqgz0jxRY4ZRvw8CRRgEE3/FmXJUxrIqsrxdseobFo7
4ybFUtWXSsUZooZ5ra4VRJ8Ah/2097rWc3b+qOjPxlb6MI/7anK0ctuw4jjQ2QBy
nEBUDY9ozpPEBCsMKoYj6doHMlOZsCA+9GNn1izIJAjlOaoB1xeV6DvdzL+A0f86
b1tn293rnYwh+l1gYADyq4vRl4TswKm6MjHGrEfEWOFQvFC/S9hgJYX80aS+sMhK
mG+QxVcJ6H82Vvc4OP1RtxhJ5CovdlsWj+GxUJunKVxIkkZHc5lXiHos0GaGrk/K
KEg0lxtiT1Rzy/3tuoh7gGUIdMRdx9gyjhdFPv4izJPGGSdX6lf4oBL58H8FvKXn
wXW63SX+CZAJRwdTGwRw2R719ZqASFvIROP6XWQ9WPxB2iar6TIJpZrDoY8DU21p
YSghJLFGjJQFDAn7F0Rq+H35kTwy9PkpaVyh6/zmDSbjA1LsHTMps8uEZ15bsv3f
S+FQRmS2LFT2qMI6l7CiEGTCmW9F95/xWqCPlIxUUx2qnsu2giJgdPp4W79qpcVF
g6cGKkhcAXqjTsCkIXuDdJTff/vVKp8iNz+9POfUDAH+fPNSvcEPs3/ezQsO0evb
BVGq0P4fwlKB8JcLTE5ec9DpyDrYIfHGheA7hHusNnGjxvgwGd0kL25SVoCDz4uh
HovUhM2mTcCEmsxP1v3ZkLDFjOHsnX4XHT2ozS5edKheR1tK62gylFtUL1fi8S46
rh6Q2/wlSPFhMIfLTgrdrNj7VzaxMqSOmNLSpKlRGahVePMYgPF7NlYdTn04T3Zb
9Kj6hT2+gn0wDLe/pfmKPmfp0D79ggreul1sGMwCLUE/1CoJMvpYm76/689o9+Ha
mP8YMZLoMQiF0loEjRp5AyZSzkiXuMjVUCkeb0dtBYlkn5fcL5PM/VYCwmDav2O6
y1KG1JJiwMD6lfwuvrOQNPbZjNLP5Bkfw5+zrvutDpp5i+sZH3Sq3crEoeQViMO8
hEo1vJg142wsh0FA1CemS+f88PfMHR77GMrg7gwjWBrXIdS2ZkZwAoYjq0BccPcY
JqYaZJSe2mYp2XlIHlu0RWgMLXAj0fqtLCXcMw5Yt6CBAK3LaK7iHlm8Qye7rwct
j1XOg2k6WPbtPitgx2/l9uRKXUzw//6HrETYw2b9/GCKL7P/4QTzOpOuRhEGczt+
iMFPFqYcYEL4ZjrYNWkbZD38wjBQoCe7G4FmEISiBAbgOa5nwUO7WkHTJAb0JknA
WHK7Vj6lgFxReqBnbcDSeeCnavPRrCf6ZQn1kVEA2leDGBGz9jMuzXqto4rpAM/6
TSVsIDON35q+MllfJ9LAJG5Pno7rRzStM8Hh3sXGRhYfuLIuEBY0aViAw0Nkc7Gg
o8iFQoFBv2gTaMjcS6zA8TDw6/SOik/Rm/uD0jNlEpY7hfFh41naEIrDTwdk44e0
pFCosKNZ+dTAjZQOqMOykxRPeeKuj1tl6redp+F/+I54TAdRvaaHSYETP8QF8kU3
SCFRWpOAqhDDJot983FKcFA7teQElfdl+pycb47GGKU3PYtu8EW+FAFwpH65KQ/o
S1WfYVhZYvDsp0laQckP+C3I7I0fBdaAxX7dyvnpgoRI2ySR7D6fo3rJ0HmK3PB5
6Gvk44R1tsyjYAZKa/MhfZpzlKtJJrBiwXtkjiWe5darp7GICl/EgkDMcYCmzHRp
K2on1kQ2xySb2aVFoNcolxmNIG6uyqSK809uCU7kntMHu9kb3ntx1TE9hD6EIqmL
FIvzdp8NLluwscgUDAVXZhrYl6jyEGydQPCPHuw5LOWoU4HTuBvQUMWZ1qkbh5ol
fbV3mC576iBNEOWIelN1o0HuOLwrDzQRv/jlT2IMJ6TA87ct5SVmIx3rpWjOcnrD
C3fJDgfawMyNiJ3qwNDCZoQSDOL1CfPfGyUSQFeaeThdJmJRsg5oWY2/xBUW9TEM
0J4b4g5NA7YgiYDQPeoYOKEoZHdZvh7RmH7qOB6hnrMtMVDLCFbUzdpQEg1Y+bUt
vCPYJwQOao159NgbL0kouE+9Ho8Uy5Q8KtOUkBfRtKP9ZQuSQG0ZtNthCuNVvH9C
ZJrDpyEbWdt3jWGASu5mf7bqzCzUyP6LkeDLQJxq5hpcUn9q+DipyqEby0jcvTxV
UZpEVRb5VVU3S+09o0N37cmVqaKvT5KUqV9nB71V+EO39jMDe5MxnF3WEcJV7iSQ
RdFwjliWrsgdK+aOoAAQNeAoP6IGUfTTkOWlZpX/XollGFY6BVbXO2AtnUhLQITh
OCmHoXvw1l+0kDj3fmZSdsXHcQYhrARBcEQYXpKRW7jUu1mg/UwBKDxVF/g5neRT
T71WwnXAaCnxf9Iqj3io4jLGWaEC5IKGmJcbknGcpwiDZkcG3oTM8ibeXveo2mfI
wudPLllSzncMKIJTBTk5Eqo6l9nkUIKZXJOgCTCKP6TY9wB9+LCwi2WFHjg2NN4z
O3+vIXNlAvFpTpPnSX4CqrG8JA1osoVXELwHWGuB04Ird6nGQbhMQ8MRQNJ1y1gX
7XVdKqez7d54eIBawMtYTSU+0UFr7iejOxdMCyijRCNu/gdONHk3GEhpxeq/RZe6
ZVEbcghrfOAFmPTNgy2uYUwaqSqvog9s7zVcCR+ZJ6IVYYKNkCqlTQ6dDTwW5krg
0MDS8QGLliywtaMhIcUEaif7PeSLoQftTwAty0YE+wAu7V6YyHZQu+1OPDf/VlZY
ZqaLpOtruQiuM/f0ZDPwR5oT01AJoU4PruzxGJxiR6E737z0vAJ5lq5I8kQMmZi4
G8u3M9ZtC8b6VBV5EPR6AJkjbro8dwNNS8P2nXximNqGmPcUJP4NvgXHo5wiefzU
QtMEuZGVvX07hBhlBsV+NKDLtxwoqLQTsahGT7eKQ884aHPLbsqtj20oyT1X4gxR
0VlFHjvmaeThLqagSJo5O7sV/PkozglRrwpiOodcyJlBRohUgY1mf1BqU0hj9WgZ
ZTirlt61Nm7pyHXYdhnG3A51dpS6gVgT8PeseyLEgxWotIIZLr30Tspjk09Z7CjA
RI3NWPWvOB3Uj5S2Vdp4o0ioqo+2g3S2mF1jX1G6YWxf2zekale37gegI0JrzhJp
eDwDQ7qcJgc88v8+GnOfcbhleKwzl4+R1RWnqrLJMMirMNMglQyVvS3V3ntsIZA0
90B1B7PqfZcqUhWMl6owYWZfw6mWGpHMDUFBupg39YgWMmvjKuH+JiASAfme2mrG
WRGLBtW4zTORcpu8oNNvTDv5DmrHnFYspmQ+QT8h3Ugk0jeATSkw4VBSCzpCj3Dl
x5iE2b9KiIn8yRBMuOITuiuIhxZeg2/z/rsRXbCUmV98EOBeeu3silBlV3tQAQRE
okZzqdowD9LuZOmAZJQOE59JSJ1tQWZHllPkrE1RLf38+1qQN+I0G9XLzDLDOoug
eb8EcZspUlYnOHJ151Ot4SqWdDzr2f49ipgPFJtQpKOPHIFRDQXXe7uZNWcdi4xz
X35og5dpISJnRpIW6e4YZUq0Qap2nZ8LtsMXvbDEWC9q/Xensux6fQhjajUlszIn
ldhs6EqbeqsMRP9/4fNYb5b9lGCiUAUrnM9K4vq2Ei16Xzs3V6x36dU1Es9zul+q
KA5nHabCssNVtsb2MxmxxUEKSo74y1VKxThbSHIREQh+ElK6QDubpycGo5TDgJSN
oSRt9zKKoYvw3z5EMaK5uNMz4HvLjh87FN42JFCvF3XmRaX0EVcj88RR9OzcH2o0
yjC4jF+IBvZi3ZCDqRKpsah8pbnDqWINfFAr3iyn5S5sTedeVkiuFvwnCay/nW0X
1xwENjgYZSO4G85om6O0ASVe4chREsE9//CuV5L7Sa26Y5H65/5hM1aes+IN3nTW
HR4fpyYP06umpgzvom8ZqyvUGQJZqyWQ7Ptnt1HTC9Fu6ubQ8/F03+jvzFzNcHsQ
X1B8pgO6Ym9epjaK3qFZmBkN7OA2j7ouPYpwuSfolw60iSibvSbDsbct2/UoLzyJ
sONSaXBVoglvEya3PnGm8IGEcKcxrou1oSauGuI+NgQDEQRPQuSDkvWsb8wmsMcy
UAxxSDJEvVBpwJWIw/jHxfm1sQnBOuEwQQkqiEHDy//XRRuVW1HedV3vndZjFYPf
71K5Y32DiE+sHVS2SiVKEUtdGUjBHnTgd+Kk36yR8lbjB9RZam1YR5ne8TX6zeET
7JvSpuMWBv2G4lG8NeR2u7lQKkR24SUkE9PwcLwYw2ARbcypt7b77Dm5SKF9gMJy
6jKqQVglmIpEuHFwuTaMYE2eT9AMOFhE/GKT1VOpJo1jKOIU9QknjjMLduLvSgnS
tpI8ujDbOVa5fHJqjYxX5hrFqPmQ2QdgoXePv+hCAmu/AgYM+JFte3YuoRVxkrcK
5QOGwivZZ/78va4O33hRJAm9dpOu+k9BFJppObjVol9l2RqW5MYugSiQ7MselxCu
so6vAJ8STdEqg3WLg/W2wdUdrtjO7+wJoBIx7h4/a+Cw/UiLn/ycIjxVkpbt+4NU
urhY6RzH753fnUdN/UPYKn4+dueyevITnA6oDUbbIO6EWaNsl9kGRi89AkwvZgvl
5gGwW317dJ+gC47gz2Azp3iTNBJJtrC+lQZBhmS/hvfEx7aR7lry5reGGqevaw18
fWHUzFmMbvjqAD+LseOpZgtos4lgZXydt+Q+8EnlxDLeDt3x09s+jTwU+KyEHHsb
sOio7Wad/PQQk2zutwqXBKZNWxxWT79RpfpP6iRCfkVuc/XKLsqsQ9cdloKYaHnv
EB8K3rHGhFlKe8s6yjBGSEHQdGCSznQdzmnIswGtNdaJwbn8hPOkRQOr6UlHbJ3b
AVjq+cTuW0oaZEUVGgrpITVf24SidH00E9UBqkGsfSzU5LZ69jctV9gRWLTU1Jeb
d7kMc3xu5f5phHTKEutlZ7mPqOpBKdzjar5hYX4jcLBdwZnMkHTSmqEJF0vUaSeM
zOD6nwX5X0UNJ5fOAQFRvwc/dR+sEaxQ4VI20TZqXhwHMsQy0e3+3yVNJGSNEjfq
T4ScTZafDFJwRwMzZwKfqdbaqGILh1wyqPumDBuJ42um2D1wdQzhd5rmULpxxpVU
MNNP5q3CrIzixSAa0OzdDsbhdVpr43Qv1CaUmbGkAtcRxSlsCuI1liCQDI+9TYde
f0sn1nbucJlEW9VCkweGGyuIkqKrCslZ+H768qjbB3eUP09BP9FqidbI69v4Tv/E
AOUE78sQePsNppATvjampNG9kJn/THhcq5H2W5+8OHNDFkTgZZTNjI6lSrNU91gg
DCRxZo8/AWFP1zkado4LkzO6rkOy7Ai8mj+S/bhKU+b4YQTtqb8FgHTbWrhbgpPc
ln2wdcnAbL8IDQy/DvcG3J066p9N8ZKyJ3m9mEzqOJqRoXklkfJkrE8meA59fIEM
Pc7Y9x+0k96v6uhrJehw8mkGChWErnKPa2RCyS/FBxDIn0dTVxQhny8WpQSg7+xY
KwtJKxn1EDK51hHQqDlHf+TWVJXjdAwA3UfqHhFenTnP3SWbMyehS55NQJO+FaRf
qGOAvXDhZ8n/CZ6BaIl6atOer2EvnwB8+Zd4r3gHsezr3w3VNEEdpfph4zIHxBHA
EDpEjPb7D9RmshP7kGCxUoF9uWxYH8+QfgDefTedAsCVEHL+ptU4AcatkB6eV+Mb
zXY77b7PVzxXqnHjebFTNeOMPQf8Zb5w8g+EcoWg/snYrRwKSR1K7/oGnWt8teP2
qUy/VuRQ42UQhvbQ8kAfxVWiY2jcj9SXny5mBZ2/4OdVJrM2OzDAQ4PVLxJtILsP
iI1LpRT76mccluIiRfnD60tCoCPpYNmKMK5yWCbhXA+jxBNnSBgeZFlW7K3/dR8r
LsVq90OQzgBvghXaOx52DSpNkA05Ys9o0gynZGgtkuFkrccKlf+gOdHWa2AHEbJo
NtUxNMA1MDH+zgK/MmDvKiUHx5nUBDShDZvOMYoYmZmH2UiUnuFkJPwKv8jQ0LJt
ao/XVJiQVnuP2TxNSj90S2PYAE4grCei+YoqLUGrhRCORyxiBdB3teHuRAPMY+hn
Z+Sri/l7jOHwwCE/q3+R+qiOCSwrIwz9NMxs2rOuTuQvOD9b00edImssMNSNQs6I
crpE07XcUHwOaQQZp6f2liDzwkO0JHzTmBTJsSdp9QTlKliR9LFNRLF5ca+Ew896
go/5J+7ORnhVrmUYalIZ3too+uVziT+zOB8SoIMZvAndElmJEXkXfJCbnUqEcR65
dqkWKQocOf0WJ+WJc7ouYGtFBuwQpgK0jXXhxpOCYH86N8VaWPm/VOPdzkIf80BM
z/hs4UWS8eYfbD4dgPVSaCVoWoZAQB8JLRY0oQen6r0i79y18osuU7AAbYpQ+th9
Zyrg1Vt6kbAGGzL4uBo7qOrRmwpg0ID4cYuZ9z3+A+5gh51GLd5t/Adw5PL7Y0S7
+yZMcExdvznfphNLn6bG4TH6THrgZ2Ei+ppJO/WDVgCVnV+XHjzvE3e8s3szTNcF
tUanDqh7aZ+jKbPNaDx+ptrZP4Qs+qN7TVmXaX5tU4Jmd/RzkUFGmoMPLXLz8DNj
k9r6/ipM4Mi6ih0XR0bjIPpESS0TIbyNHOZWjS4IMB/+1lrLSnqInfh/jEJ8ib90
VlO3eJIjiYTef5nhmAMI0jLAD0SPtI2NsYMWU6C5FOD1vthgrJyFQYHJQ9G8cnDX
axNdltlb7WDsEhg6OBpn6Jc8FAkSSg7WWt9+HMZ3wU5h3ExMenHGQpHwI2XW/uaS
Eg/4jQ2DLoKaqnsiXznWzyQgqYpUu49FZrtAMyh1bo4dl899P2eKBduVGufJNBce
QwIbv+PRnJe8iJ4XV/NxRdwovXNPM1j14YmgAiDPr4fG3N1neY12CTv++jhSvoOf
vxbdffx3h7aXISbkwFLvWgPFulFcpfWiUrbJ+VKmo7zz41T7VD1OHQVWGA6oQDt1
KYKIzQVp28SfMcUrGQF0BlXxN8agBYxWve2nRb2GDg/5biUY33UJlrGr91ODWFFt
2r82VPrDq6V+bIl07GXjeusRPp7v81cXYgzAfwDq1AWVerlKnlqnDcK8FgfbkVv5
ZIlmTuZlCnGgqE5G8A/6wAv3wmtriMp4r3O0dCtl4DPjUMZuNB/+HeTQ7ypATcc+
0U1lMLjpCEP5KsydzDwDze5X8l4jSHQpPo1y4SrSe8H43C3+cHlhkPjuHykN0kwd
yCiIEiu5C8fjllPhtfZi+a79YqmSrJ16P9Bbj74aklGRDis79qB9tDzvFPYajA7b
s/y6HRD0lVO3mTx/WagOv8q5V9EXAF7DZkDev9A36abDu636AP0UnhKsnbkO4OVp
3GzrdWnUq+oFO5G/p1a/h4b2rwFPFhcGaTmkJob7KeCfJ8k/fTw2lpj/yl0vJOPX
fEqGUIBUWD7iYAtzfmALSAx/BV+dJGOJlHqoPYLOlbTy1i4GWzCnZ2TscA/d2Gfx
VY2mjgUxutaobdTnvTccNtj0oI13mpqecMzP/TeztUVLfJeFEfvpd166y3PfKoKo
Ih9/QBAL/S8h4111H+MaCevQlyvqpM72rD0rOAncPJHBRjVXPTJMEx8FXMZAc9FY
g7+lIKxc2S3PCA3YcjwMB9/5tWWpunmNo6wPbXDSyvoOSZOBqVyXMD+K0cNZMkxn
I1GUyeeKsbZ5DQOUB6GjIpZR6WkoS829pvHOaH3oN8hCr8icZU5Ovtub4rQLOBbt
uOyYyA4TGdnjK3yZOvi7+ZYyb0wlRomGtvEZr+24ZnIBfiub3Rn4h5G84LmZfYg5
j9rrd8UH4g6Q5V5ZkdRX4vWBpbLshEUrt6IAgcZzTygy/md32v6FMsLV3mY3go4k
zypDCEsg0us0G20uHEl2XFVlAGchqzZfwXcY3+o9RoqycHEsC9sx3Bj6JsIpOd7k
FWXcogbVjo9rzJpomuwhvMR+cjux5KTnwOIHZwfOHFmvHE4L1CjPSiQKnYviWx0L
PmDtzYeRO+euiCI87ZXWmQmmomkota1jtuvA1HwUuqKRYlReMH1B/FJGXXA7NLDl
pDoXXC9yFni3fAOP5QSmzdZEajePkZEioPz3onwRylrAhcXZ8qNUhuUMi0VSosVD
LMBZi9lh6zAwtw2MIxYCZSeLHjILvhxvLAUF2sC30do1iGNc3/MISkJfgk9ymTwO
iduP9Ev4iY67ht5UvX8kFw3xxCTkeMot9hJV60vbLcLLshJBD+kQ0IVYXzaYVAWK
W5hping42PVK8GnrLG6/2XFYg8C0+528N/2Z0OaRM6MtEczfxKvsWnsquJ7NbC0p
wAkpDz75WsjFAsXyXvD2wOM308IlSAFrtobN88Uq5jYaM4gdcjAmfzuhSfE1Uy5R
sirxPdwE069dmzBm9OcM41BaChj3U8/JLjUTuAilm7JNhvMi/2mM0NWfuf/+l//f
AOyV5FugKqeu7C0KMHCG+cil5Bu+3DvlRHbElfQnr5r1uhCo83BFKh9LpKFv4QNM
HggSew4ZyPvKKqeqM9u8WINuBWwL/w9+II52znQJSuNqFIVoK9urkvyXownE1gBx
hMsT8Ie2gKtT4+CHyCnU7AtIP9iF2mbrG67BCJdfRgUEZ8qaOKcoHkydhNiPpJpa
/9WcUMlmEk21iJ9MbzFJrUSnJxYlJfi+sTNftrf2uXYWDaxvNt3CjvZfKXVLoD4u
N/PgA+Vdx4BQPdM3oyp+gQMnh9k14g/x8Fz+euW4w8xSTK9YrVObzBP0wkIPT0mh
lT7GeHWbeZqQ0b1evv8I+4iTjzvP3Y1UAR1HZt1aG/yTGwcovJ+mbd6JylLjeRdg
mcJ7HpD+7neDQSJTugWsHbfMJpre7i9bzAnT11/TMvh6iVYiqQcI6skHuw7zZX1Q
8mSdXVtrNlWSmFu0T8GKaRjCVvFQdgbYanuMW9JL3RzqNmC14nN6YUtJo6S//zcy
ILKpxlQ2VCr9+1XN13Nm6BZq1UWrl0+42z/w0aFZDO8=
`protect END_PROTECTED
