`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W7Wy1zi6fUMVnKUveKIwcMyJ6sB1BxXtnAE1fFge//IdighJ6HD8T/61TF9YDxy1
1HVxyCkA7GS/npfbP5pb82xMmiUcbE5ITReKpWm3CIOe8PPEGFh52ZGw0LNd0NQQ
oA+RfuuTjxr/JPVzQD3gfVe+ay3OPRj/TEN8qSEeOYj1cc8i0xdus7cOCzzUILfo
QxVfpbUVz5EZllAu4x4SUvSjFW8Ng4ytIsIfXFOXlJuOXAYPt/YJryzi4Fs5iLK+
I5CKQ3PRLtiA3MPe0nOpuZDNd3Azfyfdu4rHjfBRai+TPYsevZZFX9oyRLUYgpD3
fMfQG6XTH9Qqv/OsA8NLp5rUo8GSGXjEhScwF4IwMPviVx8iof5BfENiT8KF4HVa
3RKI6T9KpfDu2GBKpH8k9WQiT51q2HKBSl/GHBCrgbPSjxyYPHqmRDRky0d0V6x8
0Ujd7sVa0V3w0Z+S+K5oHLjWLUGhBuU3w6f8Oj/TdYG0nqbRnfAJ6ytxgUlEs6qk
HhQwmLPPX4xcrP6qm3QHWqxN1o8QksPyJan94pnVuS0/WRBwDjGBG30QjJrtWBJc
dax4q28eiY1j4mXvqEy6SxOP6ituYy3/lULzmTljSIdNt6PiGkY4OuK2QbwYoirj
JB6VVhUmkXucflpekjic8RFBBM2/dLwIX8f1tyzefQQT9RoZyyIffxJN2KO/6mR8
YJYnmMBIQ3AESsFawBc1Hh1deTGLMkEhIw1eYi0cnDxo6vTaXssNRuHhLWXJ91W8
aoqADzEz71YX3sB6hWuhH8JVV67M6aI2Db9tQm6zZRM=
`protect END_PROTECTED
