`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IF4mBjeaSP4tH7bPQSeU50Vi4o3FoH70bR4kwspa1W62WcFlMdaX+Baaf6ke0y8Q
52U3HkAY5TKExXLKRuYGUIn5lJPYwCYzLSnFCWHgDqmYL/SUIC4bo/CfGHyKA17s
yKCvCKWTorLECCrWuklNqIuCI6HvjPGisDbBGsq2uDbUZzhXgdC8UW9XaCMkr60u
cFANex8RIR+M1lh6xgFjv9j19pGzlzCX4n3nkhSvgcbVYTt2yonmb+5jdwDN+iyh
7eM+Pe/bni26phyX3N9jPm/V+I5I2xMhYrNcnWfEu8f37MoEPagNEjzABm8gffml
YEsPkmSWBRkCi0vKkqMAUveS1nyd3QSdfQ32rZNO35mram2C0u+FblY07q5zuEfy
OvSJQsw1ef8KZI17tOPDT4E4OVsmpvlsrmGVPI0jNGWjlBP6Yq1vh2ojuhjsbF5E
WscjIdjNvXMpq6MPNohWPQrPzjBQtAEb7Id71Ud2Choe3/YBb2BhUflBE/ipkUX+
Yh1g1jpR53YmSMO/85sEmMzZZFTQsHCJ1sVgRjG6/EX3n/xVo7/SE0RWF8q13Lbg
w8jTcKjvgpkCu7znGgDIVE8SmWo2CKCySP+NB22cEQ6caWNaaJ5tiIxMBzsJKxo5
lQDbM+AIDPEZC3BkbIN+Wn1W8CS2OnEQ2BHcdUBnfmw1m9unZeLGfY942ud17sWa
osFo79gUPQ/zuB1wXYC04zkOwODuz6fTiql7aPGwenk7Cln451jfJ6e9k/JsoMu7
rW0ieKDudIxViOmhEdRokRjh9W26Ecrh7WZMs+qod8NQMy62k3HILnVQyUcKqCKF
9wB3KDOpTOeyB5+8rWq2rz023z8UeVa/Aja6s9xGbtA+Bd8qWQEzMoPPV9wigJ5g
0rSFOcv6eWzMOGcmoW3state0JTc5I2syNkjkHaPP6lpcdw6JYMUX7gV1oRx3Mmb
`protect END_PROTECTED
