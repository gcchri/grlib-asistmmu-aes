`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yuVvYyWbiaQv07Z9vLqBz0eUGz/9WBWPufeHvH/Vc3Aavme7JTWrIdSbyZA3ok1f
Z38h6bd/PqurX1sqgE3fFmumbhT0rP3gADt7KFzxgpgV0nHrTkK9ETFbWrJ7DSgj
CsRolw+Pcfm1CMy8AREoxRjE2g8gazuitt8X7Cmvlx4DL3xNBUk+M/Ug8RCM+PcB
fwWxvkivGQYS9sY4c+g6pxSlRZgmaXVMPyEvgTYW/NMaUWgBXdlIPisQb5GDpkmi
rz+qc+yCNRIRT/4Gkq8hp7cD9Pwic+CJdwctgVJt8Gp/1n+kwoGiC09j91qSWaIs
xVHXkZXUh2peH4INg62u4quNKoFcSaRr6XxFxfR/sQtlMjxvepveZzBvzTph6tBN
3lYW2Ko29I5e4I8CGlgq0xMxbxP4K8Tn0oZ5agWBe8Yq1i2r8GS1251zoVhq11rV
bNYBOMIKvQSiMzE/srPOjsoXrjQkWU6BMvZRtxzxTdde3hQmwc9dJsOF/u9UebZq
SOdwEqf7EcWpyM7e9qFrvQexaCkI1fMSGE6m9GjgOMq0XU7W0DgkJAqJ/I8Lo8Wh
fnGTQihf5OUX4hdfZNUatyXbPIGhX1flvFf8/A9SrH9KlQxWbmlewWK+sesK0ypI
vUEzqsU6Md3k21RN3MdbjU21StY2c7pqdSi0jbqbeeAp8yiH0YmbRzFORdsBsuSE
CMyGIz7bCQW3RT4yBtiZYqJ6iBuEEeERS0wz/S/DQzIzfxvIlzCfUUvCXwAn+lVo
8ItYFV9maei1rzWM5hKOGM5/MFNc5xn8jkW//fl3Oaw7kzbXlJqWNei4aTbuRJ5I
Wm6ybc2tQCWT4Ywfq70i12HP475NLBEdqBEHLUcP1iKUiKW1X53eCpAWJSb1Kj8g
w94GQhYrTmmC+8hZWu2XG9zkox7mGzcocJJNDPJrrxkldOhdnl7LViM3RNfeNgTq
WZ22dzPQTfpkTwc/8j8ovhPNE6g9v9VYj4bxPoNtjjn0t3kPL1I1BhynGmB5A6Tn
7FY47PpUNx45ZzWyF9GELXIdT9Y0lej3qDrpF0biVdPnGpPyPD7LQHf+9LLw0lWx
UDh2WwhXfieKry6rF7uirOz8oo/8tHkasQH5LyR9FaOt9NHVDIj8YfUgWO86jo3n
S6T3lSMbTY6m+1fpI2YKffx7p8W3Y1XE3PeNQ2HVR53yYFA0mlOXHLaVJJ+ngbip
RP3aeDqkIcuAC/El4pCoIgjCeeowuyS6We5i7q+5wIzsKUuh/yQqQNKKeVAH3+x6
I/mW3MF/sk8rViE7PrUehDkaUBjAOjElyIweNE9BK/wA7Q4jtS2TOik5HAdNtchn
7TSOUdNK8WwGx4I1mn0ZanyrczQu/HopOKFOfCjfxnAACCDZ2mzbZ91kdQWEo1ZD
n66sok4s/KE5iFC4jrnLOUGXl389VwEL9HpR5zwfFbXQShxH3WOJ+V/6DnasbjRD
gWWdx3LArog+EYQX/CK3HXdZsmn3VvrnRKy7ZZIwSENOshzbMCLWNRUJpTeZp6mt
/1yi0Hdn62A76todWhO/fYL8Y+gtOyjzK1ZcDpjbQljy8J8MbTeEF/MZryFyaZ+s
BIS4G2itR/z6tlbncZ1AZXkk/8vwOUoq/giI7IijrvH1zv9/NuHOr8rVsRZZQaLQ
BhIVvwylyTAnQxpXhNq7ruZFXX6EzF0sVDjaIRHiAAjD1cb0yKY1kd4akf3Qy2Ig
oGV3u2bBTADGN2ssjcQxvZ/hss3arGE5DwRsYNe2XPuaTnzVcfI7LN5T9Doedtas
AvGym3YIm9qbexRfEIAV4hGw/gvFmNZuuKB+OFYuaVzB5hg7s9O51DTYrQJ2qzi/
7wwg/mX7GHBRDMkisevHwX11IhdwOwHbUKPspPY7tC2SrCLUw9MbbOYM9X6eIYCZ
tIdecStL6cV4tm2V1F3lu7CDteJYhZ39KaW0PXB6Q5VM+PKIC5hNJRNjOUDj80P8
NU3Zho6GD1lDyj3jilQymoOdhKl/01rCfg+a8yZzqXS/PHtsbU1JXCqlzVY0tPjx
M5fUqsYrxHYkagZBlSGRKTmOJUQGBpOq7y/PUpu5nc+OiDJCqAA/z6qaDjKsIkeL
zxQKC4/h46hRfcXJR3g/qxhdVqlE8KlW4UPpu6hwe57xniFoZruRiG3zVstyjsc3
pIPaAAvg+jzVbLoFr/YDfIXhKzbwZ/XqixAqLSOsImv4QWH3nMiul7snK4P1HWnZ
gl/njwO7mGwUyY1aCJBGo5ftyyjecUBbXX+MEiGKc4f+pTB0Hqnlz7fEqG94yQS2
2LRGmOqQOW7zR+o5RriW2rzqoxhanV28uXWCvUCqWC/+Mo554xxXKHadY2G21ShG
cq7U6R3NQIZ3b8ppRdH0C+5zb1rhfC0LWxrZac/U6i2uw9PDl30by+MZvVXT6F/j
iDHHVbNQETFaAvMkwxp+3Jsq2xJ7VgiNvr2F/PS4jlDSSZt0BZsT58t5KXk3vxY/
H0NooOTpsHRSMU4bIRM9CWAb9S5MtA9zx6m0GVJk8WNDZDzaMd5n+CCnDNS53euC
2BehPvoE0QE6H32gGztfZBFR60+pICKC6CvIybXgLM3a8w/smU6OnlFlJQrHDbiQ
RK4k1evHc/mxiUd04sVgPux7s3HQGv93qseIvknOqDXzc49n76gUURKw2WTRUBn7
GoSgtJO/LJNuaXT88BEq/jP/C0L/ud8Z+Ufqb2QqeksoQhE7rmh6nSltoE4w8i7P
B8cP1/LfwqlhC6zJP0/kUE+9jfk/BAGtEQVafEdAsefLhrcf7T76id0FV3yMurW9
/Zrf5KZn2T1ZZelnwV/X7I71/dwK/4ZPqTrdE99+D1r7CYPF1t3jDB9SZWLeqKcD
YkYPX1CLTWKOT43tyLAHI1wcyzwNpYEtiQsv7mBB3pjLzojiuyda6el4BKv6SGSr
`protect END_PROTECTED
