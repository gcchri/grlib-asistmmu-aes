`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAtLR9GjkubRePEOiW3qCCIqeJf9t1OAzsAs3TRLA3doWanykUgqsd7kjE/f3Swa
mk3I7iOpomnxF5I81VdFKRXwd41yfwPVjZ9IR8WbHSY+bMPXVAcu7gP/hupIy0af
i/bnIt9Js9CCpSTAYrvJr5DW3JRyFY0XYrXbjueAwViJCF1I5P15z/vqDNygTpeZ
kq9BNcYlfkv1SWquLQK6UpMS/6la9HswojUDMtARHrT+YrD8RTsLihV9lPQojwMA
1KhjH8eFZsw/LXROPR9iOSfXTeWKrUoozS9y2g5pfe94wUMo0xuKHedIN7PfenaV
KHkNliLXSylacrnuNG51fs6KXaCLXf67sOXDiDre9g+wayWmgLxKAzaDgxOmeZQP
Hp1RjkoE4fV9qZ9yF7ulBQ==
`protect END_PROTECTED
