`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Quy8JXv3qAgoGNDE2VqAuWJk+6yvoFJk+UFxS/bQN/yczMW/uaBgGmlodyK1GrCQ
HkxdgQAfkGiY717U5Hx8l4LnmqZcs9R5yMl+yka5HauWuFYip1K2B+9ckfoVLEXH
TEvmbq0Qh1cSViCJj/fx1Pm55HgWLHleDt9xIzFxMu/vBa42NmnmDJDulJteWUpr
UtmyePDMbSSc1EF3qYGJaP2NlUekee6UogwhfjsJtIXYrHlcXoGMof22YA7zMhJ3
PaYhDdyKaosuUGlyRLVbjD0RWoUS/uDKnsiPNdQdv033SOb9dQuMTfuJXdQ008yf
PJd7hQp7T8hymND7CQqCzGBebpWyN+FSMXb6HJpDxapVrRfcnSMidJJQSIcu8hDL
nEzC+oSvcaHmvbvjaJFJfgIB8PM+DK/tyKECMj9WUaB1kNvu+/N2ddh0H7TY3CLX
QiL0PGBo3fFq8CQOittv714nE1KlHe1bSnSTYE+44v9H09KfUhbfDNAjVFOqMRtz
`protect END_PROTECTED
