`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGgRGHVBBOb6XzLlG78NQ4LfTmFDQ61ep1hEQ5v4wRezHNqr89l8empgLdKK+rla
ZMv69l4K7J76XxHZI3UIUPiLMwF19CZUpvVKMctCi0EzZzal8I9NGnxMw0wNrfp0
ZvdEyCX+Gj/qMZdHJxhsNVgEv/StOyAxno50QHBb32RdBReUzNx74GyAYMSjHZEZ
mg1ODxr9MWCwmoZw6/WhGh0vw6DjzKtJtyUgLzaE51zbw00dWGgPrLIiqM7foAH0
kvsXGpii1LCMAQBiIq9LpDFQ6Yagh+m5VqwMVJ/yxdI8Ns+6je8YOnbh3Knhn5mI
nXlQb7dRQUGbTW3frAtatlpCm9tsbrZ3p4fvseCsDQEaS6uxilrbNuBi6CK8JMt9
TBAIfotK2cBIG69bLmiAwtEbYPbvC6PswjAmpbU/WPQwzW9L+bFcJaGbErr4geBL
`protect END_PROTECTED
