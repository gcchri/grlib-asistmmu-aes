`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VrzrwB4acRZrR1DfGMZtKP8LQtUPFh7r1Vk6IanyH5K01qF+7CbqH08HaDkzf1rc
CtfKaKPNULOVgaxWDb/+vu6XAM3u4av3/95Zec3TJpSKjAAfH/e8PqvuvSkn5Rgh
SdY82WMTcV4gJJXBltAVowuDtdW/IqUzFBdkqmnd5qD1Ldm0R7CTRgVLnHJhfjHl
/O5pdl9cFcapYxO1dWp2nrlqDEeMH8oqmwo4eUPek1X4G8h8zyND2pfgD7uAdzw4
MdHO4FxunxV2F/0H2+xb5UGzB1XpCtRNtkkEUIOnNNz17XIx2tP1MPuuNvjxECWa
O3cUUgaumONDSNz/efgko+ELhKL0PoPeMm56Nndppb9oC+VyUWQYb+MeanJ00/dQ
`protect END_PROTECTED
