`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0nUtFnTSs+Se7cW0gm1W4glyFY5oFl25vBiY49RQnZsPEcqpbTE0TtRMR5cSyXY5
AAKJJakL0DJfaPBIcHbE9t6kXHufxYGPzli59UjqLB0ZjNPVjcvmRa4+P02ZzUYG
BXM59IXiDIR/dYDCw+nVMt/xDCcQSUinNdQTOm34GtzkkYRdFdVZXyu4ZdS0ZNSm
bW+nc9FAF430Kr/2xqFmASBciKlMdaKGr7kAKsNxL9q35+kw6hI181uF+AEUw3gK
CwDy+sW0WjZcFFv0SJRRo1/1K3SWlLNZOfSgrBhln2IEYck/a8ga0lS6UkDAMai5
Wm9m6qbnHSi2FWcF4kruEcjfRPke3z0W/09/mWMMXz3mjRxZgzHCMPuB73TSCMuG
rudqmlLS9GlfDkKtBze/KJVtQynWZEybrC14zYLkGEpyVh97l9s9FHi3XtPNS313
2aSlehpcra8Nj2peb80coSYTjj4Ras9RVmycpxkdR7F3p/Zt43Hixb2fhCVAMfql
8dvx67XBsZAxszXCfxq3j4o9s2/Eqf8bl1NT5CLjTKjWZvjcLFHXrLUIpCUlB3KL
M7mBeG4rAgCW5r0H2aGEx1hE6vBEJD8OifwdFDVKv6VLpZ9Mw9HO+Eb6cfOK/SBR
voUTl3kxldJCMxh55PUXIebe1woGig7IpwcnjoXJG8MGZimvtAVG97a6Twot1vAs
E7NFSA32Gfq2eAXbXzuiucdW3aURpNcfpwrVAPcwMIZ2VTFOvS/FWYYQ0RkaMcPo
XxoTQVjfltqbDBSeLPuG61udYVZSLMIy1XVmbwhiQHD/1oqSUZW/zbmERHh7Ws3T
EavsQPW26a7RStRaRssVHMWOMOp6jIgejTB1d716fbEVzYv6pJlVsfYfRaetUzwX
H02Wl1zBwYnJzQZmj21g5dkynERwzsp0QzZOrBQO4hjE/oiDGCFw/pdjTaqv6efV
Vgo4ocTjkzPiRxOcwUDcex60GLvGaEJmatdokQ123Py6HVMWYBZ4oNKPVJiettt7
NM9FA96z33jQfIOKrGNF1Oa0tSfNbVw3er5W4/o3aG7gIJK00uJOuvkPOfWVl9NA
x6aVwbvkgn/9okKi6is5WQ6MPY+enn02kJsAy9XuBfGARLEwr8sZ0Fu9OUYW6sDh
o8wZqXxI6fgXer/p2Q+DKP26ePGDsJ2R+yXgzzy3UZWnElQzWHbfJXkN424iS2XF
kgDN1LQroo6e1f2aKN7MGtIVH1sw4POKaWaONvjqxfG9dBL8BnfYikSRJDVb63Kl
1Gibw/LGd7yVNHeybO2lmF27xL03hGDp+FIZFU2Mk+7F6STx3MtoxO4MkL3mpPFd
m3RtTbxAzhbomFTB+1yI5Dm7N1cMOhncXJc9vEupTticF7dL08OURNCKRRRAwO74
HjK7KVe+yrv42sj5flO2dt5/pcRWAO+dZ7ws1I+ssCDlI7BNyAnZxSCA4oKm4Jc5
6a8srHhjxrvQslN/OV8JFhU+XFD7b+Ezmrt5qrhrM3lD/c0nQBga11p9PgxH1UlK
A/J4fA3viUlZwwkD+a+8Ckn+esbUPGSddgtA8ApbHfsYx7G0Jw1cBycBclDWMvR7
SMphx+ycroex/L2FsxteSTLV+ndIghAzGFk0gGfKw8exAl2455DIkE3AYrFVvS4E
Vfmjf5J9M3HgkDABQK+b1Ec535xxNBND1lHU+XekPiIDPIfSlOK1UcvnQ9a5CWMI
3HVRkzp3AqNG/zOADQfk9YqrHgwLVUGNun1qzciZEFkjY1NgNq/pWZDcIkK2DJWY
hjBxyXhq2cbvyz/OBsfNC/HcJpKbEnmGzJ0Ldefu77PidaVaq4Vn/3RbNmSFSdX7
a0p5FIuqSxckaCJORoohLWNQFXtyjTM3z/jPJIia+pV/1NtUkgosF+cHfuYB+q1K
OYOH39zOSELzhnkGOIdAEW5GUZrilAyG+DcCpBb+nXyJqSG6IJKnS0Py/70cjPYF
6gQC+1YsUfBMucl8ccmbQLGBncCu2fFi2HVYZ7iV/IA67kqgIQuTv/roIixrVFHb
cWDNEtv64WxKcG4BO0QCJurM4qZGTkR8rjjBnlDqGkLBW4dHLkOQ4ozl6hlTPUXN
SXonsclRG5GLaShw+DaNxIeokpG3eL9adqIp5B0ck0Ivnods9peugwDjjrj1igS+
gia6i81H7Ybmz+gScxaAhCInL06+ApTWmtl/+1RAhKSDZ/i9VU4l2r4RJxaaAhvj
vzyrATOKzj7UR84noy3FK/BVnMgkjqPkGUM43/959VHlgwImMu8w3CAtjacY5gb1
tJVM2fxaRO+PWNQtZF8jAgGPUM638ukOLcQ+DwBzvf4TpEM8YOrJ7gzvgRgD3PJA
ALyRfgcomKEh6EE53XOjyB6bx1dVOUDmsWe8jdR5dzUz2sP69KEJm+WB09eH1pId
WRSCnwlVXYH1O8Zr1OoNvFBSWgh30V+feeGiMFTuCcTmd7yypBkUx6hJq1/J33MO
LBTqdZ4slw/cHeK3eB2mk4JvYTQ8Z2tsDzfw62sX4RCnqc0JrcI44+9YCqIRUiPv
BdWdJXazsxVNY7hFHq6A7H060x9caCfHbx0+dA0GOPH0cNoJ1OtpuJCWCKI8DwNx
P3X9PPMFUswdkFqFhmOugCsrqKIR9j2LoBj1z+2X8YXLqT0YTPhYV3Ak4C2Bg429
PyQOrziJxcNm/Jdcztv96g==
`protect END_PROTECTED
