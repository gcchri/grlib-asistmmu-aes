`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HdvhmGNwg7qIXf71qHWF3fMv3MwwMPK+i8nPbDJKXSCiaqlj7gzAzmlKexUToZZ
ep+fOrlZ3qnpu53/HqxdDmMhFs7n7azgwRXh0w3HbpDYP4cB+oq7ryn5wY+9Yglb
IJv5slC3HIS165vrJTS2B4Es9qaH9fXHYYdWP7hN7NdNou0n9wQIgLbyOPjTAAK4
TaxZsJWuyiHrjPitxVBsBc6hzaMGa4Tn2ntDcEj3zLGQf8FaKqYiKjO9ozci4Jta
buN4a+pqxkm3N/mTa0nrmklHJBGcukl2/cU+90goMtrpQl1lG13+gFfc2RC5zCc7
9qm+0dcotU5KyiLyRIbyh7Dz5KkQuMSJqGR8s9VSKOBJgdan3SKXVS6B10j63kHq
F7u9uz4XQprN/dIzdSJ4CLYFFVRNngmlCg5wos2B4dLbLGP7A2LlDgHnWeelhB06
OQZkKCtsVNtjO3RSuQ7SLsWF/aWnD23LlNtuJSy8ZqM=
`protect END_PROTECTED
