`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7d6GqHutVfAmsRRy6M3KouKbMj/HHtrxsVrbgIPSl0cNkSS64GT4XXSGf5RYtLtK
1FjhZKPUTVaYJFNutIpOkoANfrkPdOkM+DYee1OYBW2PpUT/gDPPoWgzWKxYgyLc
+hVWnqCwCfF2hexmcy/Eue+ncN1cFmx26q2DaWnl9UL7wLUivOPTeTZoF+C0QLr9
clcRNL+ZHIVNf+4kZmttdemiABWuZHw4RUaFf5HHC8fD6BYfUm3veAXn8NBkgg3n
g+TGlUKQr8jA8DAjJjvG5Nrdzr73QJe15j/pYpwRKo3T9Doe2adeVbfMawAQEEPh
C/CaKZUfQTi1eTRwduwuts3Jlu2F6wBCZzxpPpDmrZY+tudQD2Am9Xypa8+pg8OO
BM8hAy/2MjtgMW5sbTeL/ADXYe6ZJg9W5e5qdxgIITpZ/RGqzl6quhcMnwh2AnHZ
rUjc5sfrbs8mPeWbz08C7XFnKeqYMYkrmxsT1+J5/g3gkdaVluviF/EPtSn+T54K
3a9gt5Rw4pYhMUagXaqLi2sJoqf0PYXWm9KbrNU8Uz6uCWX+wRM7ESaXjtiHyF1m
1G8GwoC0fWlO+Md+PEgoULLKL3ggi+4tPugCDuJ8A/8=
`protect END_PROTECTED
