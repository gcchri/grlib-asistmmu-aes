`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsGVNMVa08dj9mL/mtE11vTIQyNLPPvzKBayEs4Unnm10Rb2D9tM0P7dnCnViR+G
WZVvl3F5O0G+9KEPNOdIG23Yr1fYneczKfbwy0egCqxr9FFeu9IKwTd7KpYubKd5
oeJzGOTjOKRZz+sorAy6wFAtSWdsGY8TiytX1Fmi50+EJgJAbsnG8KfZGIsdssCA
ZhEo4xvwzpuchc9mjlnt6s+HGSNnhWUalQTYBKW5w56iGYLMr+ehTcvBN0CIyVDL
viYDMyHKfx4zoT9NU9QC+9AWRkGIHguPGzKc03NRcYyZ0KXll4CMHiudKjir8oo0
3jkyqjc+8x/ITXCRGan+eaHcZfrRG+sMrgz8u+z+SDR0gqBwAhQGKov4Ub14KiMH
9nFVyYtZ3wULUdlvzYAShiJWPXLjWuEJGdn0ToUWO68jepdQ7hQhF4ZMtWiIDPsR
S1iy4QSWip6U7a5HWYG8U5SNesM09V3pMfe4m0A/LKEErOL+PGhkGAwMq/6Qp7QP
`protect END_PROTECTED
