`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u1g2XUWAs/BTUiKjBV5lNMa5dK8c8qDnLplId/46pV4gHJiGP8MM044g1tuLXhmV
bmnhPsGX+Zun9McGQ0rOEk7E9KO0o7YVLUiNS3A1kq44sigo+Vu8iXIYXolM0o81
8PMWml7exwAn2JkoMxGJSH9bzkK5EZ/LgivI4FyuPIJDFtTA7LQacNVoCw89h12h
HidO8IWZ7ggO9EP1M+B1xOFU2L6uqk2lw5hKogrdu4K0wfA3VAB/EDUM9lPXatLZ
sXL6Ige/wPLr9P5RgI+7GT06LE84RbqWzLsHQIocyhs6PAuz7JNFYhxgirCNMeLp
keQnd68DMtSfDdHSKKqIs+SV0QnUk34jJaBpdAX8qCPaIrMUjgca6lkcOhBl8M4J
RXZIj3aD1uIYnTUsKjowjW1xuQ3Z+OmRj3KYEfL0tF4=
`protect END_PROTECTED
