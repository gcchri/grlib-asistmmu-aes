`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJbfk1tgjE+A5FoaR5X63hdw45mcmDZqvJUTSypeVo4t5QdhYDpFqtVgQvCUBwv2
7yckj3rYZwhs33falJioRchv8sEKJ420/A6m3xJH6yB01ol/bN5SNSW9oWFTd5eB
oz5Lyunm5W9EnsjzcUfxphgHtIvje7ZoDwPeY2M89mRHv6TWmjm3L50+82oGz2Fa
DjhT023G0/puc+mtnr+r8g7c2Dw95dgP6wOR3+9Ombn3wQmQHhOhbOM3n6/0J6mz
5aPjoak4hn7KHFErrCMkN+rsFRQBgt2jgb8qK1+1t4NvOtQtIy2ZFo5obZk617lF
s1RjRfnufrj7DcTP9JuE5einPeMuq+LI58cqAUbGO361qnVZDg9T7PGBCVO9Qp8B
OoExtY+fXt/ui/PeyurVptCj6YAA0qNmAqF6IPr6g7MG/+NkfaJG1vBjx5WtCg7v
U1tf9ioks1JhDcKcS2YsZBpuqo3zwHuvl5YKbnY/k7Nu9Ty0uV1hBIVV+Ko5UmWY
MfIRGH6RTfK2uZxoCADYUvSYyYuhbrpQ4y6BRWO+o4DV8FG2WXEOGrxSWzqhC/2c
eJqb67AEz8RQBlqk7WVXxGXfAJRXX8UNMx3aYWTuwSX4O329QR/kQMEs8D05XFgv
wxibNWMNxR9yt0dhFBS37lzoIiKOVOasiuarvyIVmqY2J4XTXwZaOd8BY3P+3Ie0
k+KOLlYJsUABfrRmjT3calZdgA96wexx7nxo+SIjRvFpQcL9S7rLS9zAvHOMwLqT
SRM6fWdyAKQHrSvFc1ahS6Oy9ZNEU+KOhhY+XufL4FoKYnY7Jw+VQYUn8TUWZBgS
MxT+/aBV+4B1PpId4zL+n+CUmJ/O4NcKmYqLbR1ZbeUppEyGRE2TMV8M0BkRMqkg
U6KyrwStCqFp8aZLjnHJr96mzZPahvuI0ofFWW5/sXbKktU+BX/3MrdQVaPgKm4o
4nSWp2V70PpymHqxJ9l5EQDPBcMBkryj1jOD4lFHJhZdKxRINwYVZRJ2V0UAwJLR
gtrUnr5Qf9tgPJSggq8VF4OTLlQmRouUWmVNL91TsZBfTOcWCOkHblT2kYULqLMm
pkQInQul1Jh3lpU473g40hCbcCIN6VPxyOqVCbIsC/wGtZJws7nRg4XcltRuDB/x
aMvF7AAcSUMcQsS6uXgKw0FqKPZ9nqRdAsRyqdi8DxiZPiL0PJd/spV1NloHjS/y
pK9l/QqLN8T2jPaNeP1uhH25cea4T7PIUrIDcMpGFR1Q/9hIBKsusa1WQ9mymYpw
nFwdgz1JRLyetitNPD/BOIfLLlkhMLb7ohYGyHbbSje3f1bLRzY7nl00GGl3pSb1
dQdrm+0vHuLEV0PBDYegH1N9277ZEN2Pz3ldWbgr7oYYdaIl9eddB0sR4Cv0MHfO
sIiVNSzzFZx7p43yivzbm/4MRPp2QHGYcTLPDWagzhISFr7hZs/5/VoME1rwMrlA
VZP89KGJ3moEsAesw1YxSlssuRAJoLqhgu+8J7QzyMVp9HEv2wHp063afVYa3ecw
xv49ygu7YILm58eIIvPSf0utoUCWDp2fKKw6tkmD33H71C69TB2q+qPoRFN2OLq0
SwpP2KrnniaoFjifi3xFCubOBChzD8eF8HA//t/6UhPHPh6bYCTFmro+56YJQc+6
cDxplpow9NkyH5IMR5mKd0i4Y6UkO7/2qqO4Q7u0urRZCyhHztEgj85fkMbyiSKQ
DEJECeI7qjOsEb534gXrV571GykHN36uBnZL1OShS04Ovatc/q723LouLs/Th1Cc
665Occvssk6ILr7Ielc/TA1MU9gurQpIlRWNV8RZz9tm/l9QjS2ZnH/0JIntalYC
uGWIiX2eKJnamCSpk66zWqqqn0FpFRC6g9ebL2STDwFaRJ/imDYzo/G8QGIzmMzt
yxUsoZmo4iSVkYGs8UeddzSTwK+0rNcF+THVXi/PJYxzsKJAd5PQ//JJqg0l1D9w
uvOv4aOlJ/vTELY5U1Xf4QxnwmbYu3Xr9+7SDcRy6HDUDMjoFx8Wn8ymUAepdm52
KCUMd0PRa8ejvXgEGlLmcp48Ilp7WtX6NTDSg7jTmxq02reCfB3UqXksdKnFpwO8
U13HdrPsuHwf+/KpchxTUCdcOVNhbdH+ATyrWyZCP/NYx3eDg3VXI4gMYU9JyXEw
jF7/UXX+wX8Gd+PPce+U/3CD6ZU0x6sdlck+Y/CTO8SN7SI06Hu9QX0WldyGHKrO
VO5O9qoygquT2uvkYoMVo5O6qbQixgzZCHfGgi7z0qZrEMYuqMPOaoeEJ4fq9/FR
OcYiktrU0Q7u0l5gS8mI5NpZuMzVMjiPghg3WLQPjuQBtu3EP9U4ef0GMnprqEHR
RyIdrSq0wP9AQeVAGhsfrLXSAGY4utxL2uwLCnpBoTDjXmAQfmv6E9tEjas307xa
C1G1glbfyXGL1CgZj16ebyRd9aikcfjV0qmzgTdNs9sebIIKUo99Svr5iS1fUFeh
LrA0WM8ZHTTPBGA5/rM4rY4dsQynrS9Kj4WWtIbfFC/JO45CJbL3QEuE6Ct6KftQ
eNS331f5NB2jY+N7SKlcSyqyKhlptxWU7CXsjWe6h5/80lUbGzu+SjaHepFuUFX3
08BTFrpZL5TftOUZ7l+RK0MIBwqK6s69w9HDxV4ItfRR4FmBFiL+/x6vzSvp3IlC
99KDkIC5i+vJpYDGYLHQTN20CDvaj3fA8gAqLQOAu7VSoJjQYVTTdbuKUCCTtSPn
9edGN+bmYqRz31wDH+VyOD03+4PNdFab/v3+4PRuhPhNbHx5+HD0a0AQ48zmHx8E
X7zp0cCAw4n6jS6ydR9f4iYqv36f1ESSD3fnZcP+ZLntDt4YfMzTSFqcvHIQU8OV
TGLAathrbn5S+0poBTpkessvdk3ROjb4FfYvgK/mfVuiz9lcCshkZgdiZvyko9ko
aqlXQr/uAqSRk0zIweGGV5N9EN3+ppmtGTiAKeEtxlys6QIwACeTVuQ7pTddaBos
FdkusMRJTuPXbuxTNxyY2KBRKTAXiCcwxWhwhGqYHgGdFRe9WM2EErCXPCVX/FzD
PvO5v0lr85/JeQHGd1LHOu16Bv3vhCmLR8uwD2HBfmv0h1d/0M3h5n06zKrWiHcu
NHyVBSJtxMVyw8SIxbjF49L+cvBGP6gR19KkxwjlWup7hhY7okaH+LogsaWSrCAS
oSy/+Rc19qvQUdAqZnp3hwXsxnhB7Qj2bIfrElQ81RZFOsZJ8/1FpKoy9roIKMJW
hJCWWoEYHaXo2tD9p/BFcTeaA3vVgt8XV/6h3amdbN/FnEPdVKBTREbhwse5EvfV
X2vtpS5q3Mo8frwQr/u9dgFD1Mmf+eWRSdzJLB/Fww83bOsEacZGI2u/3t/+jjK0
C26w0Sj+Ql9KRcL/HqqWUNABZ5lfXcyR2ZI3ribgQG3qOBcOPcf7eObaBD6+oHuw
/RfjRZA7h/mRLnXZ5fp1RHgNscLnY0YmqWCLk0wMUoYY+mfSPUNBP4A3NgKdmi1q
0pR2Ul065El90uemTExaswpLZt3ypSF6da/kXwk6LcG+uM+PqitMTICblm2x+96r
jLwEVZ9xcfG8GOp/i7sTnGrn5qHc4uxSENHArFVIH1Nkmp4alexMAvpKHHlxL1NV
GB/9ViaigiXdGVw0X+Y3G7Rdl6lYoLug47sLJFTYqWiWt66KB8fWS55pw/uQp5r3
s5sj+epLtQoXbgIuuS3bBAhX54u9+WWB9A0u19A+6GbhbtCmyOr4sSJV+i4OEPqM
7kLWfahnMGHt1FauQgRKUZoZ52eC6hadmsIdELEdvJDufTP6PSXAjQiqtrRJMTK5
coDUo8h54G8Q9PGyI6wQTPRR+Aj89GID4JoJE0C48gBMJca+1MlenQyAZ5rzWTPP
WQPWDHhrMj2Klh7eA9EzMpPRRaix+C8cEaiab+bUgGWmBP6IIONiwIan+RYW5m7x
uX97/Q4XhHFbnqGICSkYk/7hLqzjPXOel0dULmfoXiV28jS/DCynL0Lv9yuBswFr
u6toNLHDahpqfn/+Ld+ofmZyaUtkPMAh1Mo3jroFadJlRr8mp0bIAnTMMX5fWgjX
/ztYBlFmJAWdy7puBAO+xnyrk241ugvgr6URzr0h8N4v2w9cmFkfzdmlugU/ZFmR
GgaoRkF0Q+AdaByZ4WOke8pCbDozyCMkn5GkhhJUqdDFYutXGd4dgOwz7G/psWjK
1BxmxPm9o32VFcuydCMB6jwXBP41Z+En5KA5cf+JSuW+vKwTpw7vrDe+nROPun+2
gGg1UxmOjykmeIfK5l+EAW+wbV63+WPNvEICGaNjL/AI0HioSOKp4BetFjGDA/tc
cfXfYVZXlgdnEveMSQ14wqcuFXr9FIefT0pwVY6Us9lT+TfWiWIqGzQwF/7Cb2HR
Oi7w523nn+Hq638Euc9X3dMZpS28DNbDAe3kCiQJqeNXVkYVOxiTTbXeVLS6ZF53
MlRwpSs7vWW5ccBOs4HQOAeUdc09LbOCPP6fXKn/8oqiKhgjxtLDPfoSVa5kt9Tp
C21l3wBQSHQaEPliceA5XpFrXqgsfH8gVKHTNnaNnhODyQgORHWPVb0MiP1lu4JO
GX+By7Ro55ijjfK0tsEdETuTRkcMVi20g651dpewtyx7KR+tCjO6+8fxaGYKsVv+
RwIQK9FvuK8bprUpcAYZN53OedNBn/YHzrKtsKZLMRsageZjAbopWIwbIhjggpxW
+0oHZPPWH2i+dF5jYdr8IK3/QOV62Cd4PB7XaR5tl8845mvQAq67d/P5gRP/XwhR
WOji63snNp2pZwPVZoNWaRiQM5g4Zcz2tmHN5rJvMK4j/PNq7RM+HaNn/sTWFYTl
vFAILyBAC2hfXC3Elz8ODfTqnPhR1eQ+pcVYHUXEmc9NwteROolpIm7iNlQqErIt
zuwJyEn9fgQ/3KujvM6wya88m5KdI8IWuOpYVWX+bN0pGXGYvVt0UCTYvvpM580N
vhPuiLGSVmhLblXLr0dwscDehZ/LimihtSu0vRNpfZ9Gg1JeaJf+FsAsFDmHbgyP
jQDI1o9TF6RMOHuVMBRTlCo/QG+7lc6j5oAn3IPSTij5k9eRufnc8erhbygO4IHt
/u+tUfhGcdguMyxidAimzqS/ZDadhzQxd+q8Xn5UsUac5K4zZ3BK/LfMQQnxMUNZ
habaFCkiUVN9eeuvEy93WATXsF/hGiy33yvFyeJF4qn59xy9w2SqpktSDL4y5Cal
u+AK39QaaUZ5C4lPemweG64pmNAzmtV38RihpcM10B2Q7ePpg0p9l/ZWt2XWKw9z
qNeXDCCYCdpxsGq3hYoggLp8/lDgwWc7KTsTNgHwtF/c7tdTuTWSD745CzjXhvRz
jdgfquMn6s3cIgWo4fF2w70RR6EnlOjAhHrVzTv6S+ux54d7CMgLtho4VvGxSgH4
a8e/WHxQpTuw043gGoAxwI+4V8LEgDPSPi1YbC/1nyaclQhtWzsgc324J+WWM6Hh
sAX4kYk9AORjeAGzwqTDuw7hRg0MwbJWUrKmAHOuYJhQMV5HeHAdfSRuH7o4o6LE
JlbKWvpHtKLkyVoulfpnO8a50YHx9lNy/vdLW6vbt7dLCDzui2ewD3y6firHT2GE
CuIEjg6ySBEPLIKxNM4tpAAR+fw+JigTTKx8chIPNWjHmbDKMB3TSTaMvFzFKSwR
mpnPAxeLRbc895X5HEQRstAKrWZYAX5Y3+19cb6pHAsgXgD0jx1swr1aGB4LyDQA
LoyYJ40XIa51pXfiMDoX2MgluchZA1u1lQCpJ9pWYpIG+MraX17iItDU2YCdV+/n
BmUCIZ+L0nNxrHaqde7vbgzHMpvTZl0ujL4YD/jvayLeJvyqdtTKlFkty1nE5ptJ
e0JXb49PTE8Ti/IKrBbZbCXOGuTYqohrB/NyfYLxtrE8lz+bTKCks+rjUsSN1DsE
EhauSAkibzv8xD0gyJ+6dQB3C9ksUv4XGyeK4rZ3mFMuyWlBmji5SuEuB89uk1OM
wPmOGcgdcHBing6qkEWCmTVdJxNVZPukigawrHOyKu16HeetjdN+1JINLTRAr6Rg
UbIMBN/Le5MuTmMtP1UJ5FbW+bKYtIr5PE08D6uQsBQcRAHaAAFsdlHwLNnayDTp
8GmkH39PbU12gbZFPoHPOCOJ+quHz6GNRDMveg3onnLDrAKW6FeiDo3iF/X/fM4v
Rx01UEwMDk/1Qo8I1ngNpNNhbVmaCWgt+jZ10NGsuLo1s7qBLbKsGstcODbkpmQr
qzC9D16uVdlkCw5f4u5oubkpHfesOJ7HLLxqvqAbJBaI+0+wVjBJnh3eREeCfk1+
aLhXL/F5Kuj7d3Tsj2sOHyJjHzupG672VXZD/74Kr88ps2fqUzMRLHgvv5w1+l7K
+5yPgUXYtsFiWDkIIa9nlo0mW2U8WWwj9jvPFGyvFT+MrkfcRO6jlY+22aWCemVH
hB4sRSzZq1/GWsTLR0xuUbgaB5N23rb+NDddZ46G1i2uHvCfmBswXfKDLPeR4am5
or49JRVKrH9cEoyqTgRiuyoY9HDPKrYLECQFtjeJxPhXVSmJBoshw7klRUw9O0ac
mB4H5Z6BntIQSnR+QpVFfJtrWJCyHsiVKcPPKnuB7HwY9X1HrmcNuuf/0k3GKx6m
kUOLZvJftksbhdDPF3vddy4lJ3ZMR2v+vKhrDp+hkAK8jmO8i1sEWSJ2uU/kpkgE
wEA3H+dxQwZl3e4raqNfzgfp+Nc58dYkX7Uv0ulmKAAG0N4fHPmw1yYS0aYlgIw2
ER4/FIsLoVQAoRWj9IgqaafDaIrJvlNV0sBkpLrk09HmA+qFYJluMNeX7rGU+h1b
F6j9NWT96h30zyPVaZ0KLMXcKMr0sWzDGJtSSoOOZDhOZaDHMXKnJCaFio2my1wn
+Vdp0FJuec3Qhh48iRe5jexVt8vXIQYXJDLiMeKxTzFfMzx7MUpHzcT6uau9ATDr
bB7agXUnzg7h85TwpRROSYsG6K4l+FisdZTMXOsRXhMO9+oUwkHBZ2HzIgYneUhv
oZES4It5tyCW39/dAA1/n55+YSQmHJRoJVIsM0kL+jeODGL63kwoXrfBrE/N1wcD
DF6hLE+e8vYONS8Xm3aoxRLT/FEWxG/mwqs0vOT9OAJ09Tms5PnNXrp2Tk0WnEJc
k0SOf5Ixk/MLhwdrmt46GCSKjv08BtJTqNmhJD8Gwz1P3ln1l1CfUbdnJSSm3wMG
rGsElIuC/KA89Rkby8Z8NqRO/tN10/jQIcbf9GqoLJKOos2HvQQsQNbmCwamqFEg
s3/Kw7/1wQD/cQ0IWgaJP1FQnP/CK3LCd6ZYlFLJ01Tgdl12+iOfR9zTxt/2YSYk
cigMRjeimvuE7MofzseGKHG3xp2cpb2t8HHipd9Z0wadBL41Xg2uJ4EghA95Mwz3
Nq/FVk+9NpgWbNFiSMmFIWQG7Y+bOI0ic8QCifZTj7kE3Hls63P9TKoRPH64F3Wl
Xc5spyuMTaa2TYIevgXE1ZpFangVgCFO1igLfpjNbbrJdzH1oTkjN9XgOlQSx0DO
IYXTIpkBLVS/YzWIlo9EoxhxeETpA24rLPVEg7YPyrsX+ZZUHEQR7j5ItlXG8Fgx
cW3MqgqPG0AeQjRFfEZGrRp7qUy7zkd9W0zmFyFZq0NWYBFJwu6A/MC0gKOIyqsQ
YlwQc/xdagWyX3ab/ynZ7rwpZ3r/PzByvtR+feOHOzHNV+EsXRQ7PUR5VQWQWIOD
90Zc+a8tXsm7EK5nP/N5jYgIVYe2YhkGRUClSlCD0NFNCi5855o2P4mUHMZc584C
NXZYIplz0x68r4HhrskFouwdM3DS07wFQsEsPtBRa2l+XU/oVuSPkEEIhNv84g8k
3nhBv0WOXvKypzEiZv6PSppvwETMeLWpXGzpCWj2mwy6d+HOt82XlSnaOvQ0QH9e
B8ox4AR+kUncQDi2VIfLpnKhtnPg8YgiEebYrPbmmSVHecyHAVuYG+cI9TGO4vkq
1EryQyrisyfbJ4SCnd7hCrViGgPH9V3r8FUlcdYy9W1vznPhDWP6lCyVDZc9VNfZ
0OboRG7L185Sovl+OcwxGOa8dNS2PkQqg+aF57pKHVWidp4KkWFCPI5T5W1T98+A
PpdeQZmyTrzQkPFrgb2JPlGw1Oz4u2TpkTAn6Itkubx+fWsId3Ip7qCL8xEDHTJz
1mXDADLe2uYIYBQ+Q5lAqn9tVQhWcURPixehmTrB0d/btPKPCigRH136Gg5maiDS
32Qm26ydx804LZHLvEMCaZJbVf47rzH9xZQyXDVBdlkucMDTfmPPNB/LnssKS/pT
xVDMpY2Pz1nTObFltGY2vLPqQBx3UTnHR40mvhao9+OFJFS77RJPd9ybWV/cUEsY
gNWgOaWUg1L7Ks1fiGY/acgUev5CUqp+ZkCcJui+9Ew/9h9mL/Lh689aOxd9i7Dc
ZhVph3hj814nbytNF9DPPTu1t2WlDkhjw6kDlsdt+zLMzSg99NlRYT7BWlXE1NbE
8KQCeQEEQJp1O6Z33UBSOoNFcZNRsLrB+O3RhiYoXAbB/LVg7UcngHdzubbQx+c+
gv5Yy8xL2ErTpv0Of+7CQWjnfMwmLdSLdDGVt/6Dv62Pu8+3ejiUlsSIaz7mlLAk
7zEYJvY+YrQFdkIrXF3ZsD8CVUQrlgui2nO2ebRlcKgdOdNpkHP6PB+BV1gix9sX
f0tHTSrLV4qSJM/cEk/M9FRVebAGBRSUEunW0kttswZpqXANlu1KALNJ8DSyzsrr
RaoVU0yu9hVEYf18eytBxrGfJnsasJiSCT9xQIUhNz0y0uYzQPE8nYX2SsRp+VOl
jW5urnniKjS/UP2VpJtojaOC6tlR3R0x859CXK4+u9WvzrfdaDGEjQtXDQsNXu+D
s2Xcn0uhm/BKY2Yr1uXT91iiDr5WNh8Qe/ZxbCh35Ia0p6ZSVpAFExsgORWYZwV6
YsEdYF3Xub7zOArh5LF+Qb+H102aa91pbDazz53TjqV+pNIgmTtyN5Dc9rESH+kT
B62gfqoCFFSrUtn1vRtyoY9rFlJqCEiTCXDEQ4o6kh0zuiCKaMlnMaOUZvkVY2kW
InJ8uzgqd3yItcCr4c0Bbpz28m0z3qPrmqK4gzEpubg7bdROF7ABebn3m5OPEJmt
wC21CznOSNEdOgPnGiJeF7dKiq01IA7qfZ1ul2CjzFwgmIpG/fjQJzjldiAW3b7s
ik6BChg1T9rPMehvOBJyIHjbKVSVyAERM2WpHaapsoV1X4xWVvlDM3XLeYPBin8b
IuTTE46l1AkouO4Qf1ygwPmDurg0McyKevFzQaDBzKNx3Lgr78fqVXs1BzhDXyfU
2XDxHhlFx767U7u4x+xzh9yXe/Vf87Cc7LaeVycsNX6uKzYBVKyBbg7+CRJpjgry
XuiQbIKRNaNByKuUVqjM4AFmH4KA7AU9WlajI/CZJydGgJyHn1TCC/p8LrjN3B0N
Icm9Gi3d01FaSvi4r6Mu7B2vknMEB6zNtNMp7nrsTjuH2hnEpTzOUQDY8xoRJ5C2
rWNpIblOTaBGyq8X4RRN4mPgjPhU+L4EOqfaS2TzIdlP6kWoSxdoxwMtBlGRbGo5
l8xj3DP3R087H7kxI1StLl5wvQfNma6vIiki2+AeXLzznd3qj6f6/zilD3md/0vq
mFiK562gMKFxweI6RNb1SqxFxMf2rrV7t1e4nSwppLS8O5omYEP2NB0yP2JpxqdA
rdu8p0AVVHZShJ9Zn59NOuaVANqbgYgfT8Q76+SU4aVI64rSltCj17x5NGut8Ow5
b0bEwC8UoXCpKDJ9NmshHlLdd3eUlQIrWPrv9ZZ1+CUIN/yulmbl5F43f3RZ06wd
Mkkm2zUsNUf6eOqvRQTqWvVIvSWPomqrUrRYctNytIm+LhQ5oBse8GYJD0LHYgQM
XrXLMcYV/k2hriu09Fr0mVPtb4XT+6RkV4kNOCi2ofo9SCK7JmkcBgU87AyN0Ax4
0duyuSykKPE2/RUqQxHyBvh9wIwEhxK4anyld5rum1gro/YmUl50pX629AMLEUyq
CIyhrVoXbQyiclHWey9ycm3BgGgoDzVby7R946b+9xPMOlZOXU2Tnf7/UCgusiep
gRCBQUthb+vJspjMZBtuEfAbZNM2zkKOsop10+sh4A0oOVX+BZTArqFcVSQkkqTb
+1JC+uccB7iPFqmqTwNE+iW9yO8Vpy4lZ7961zuZ/5SqZQkZIWIxV2mYBeVYL9JS
THEBlHW1MYzYinvsTEPwm54xsesJbWcnWhy2Cl0q+gk0EGzf14uqmKvLN9wRSCii
nxk7j7kAkANh4sUVMbr2FyA1dnurKrPw7t2KuYvSmAIQD/c6tU1i/ad7s/8KQhOH
5DiHXpOYVOJybovjI1UK6I7fTN6ckCBBO/WJYaommEzTpOpVst+TE3i3oaOw3CFN
RFEE1lxr9IA/+oYzAiSOFt2riyOR/09JDJQRQKoY57dlQfadaG+SDdCZFFJZUsfx
991zZ9OsFIX0bqzFIif3BuvpKBPLeHSosIveu+TCyohYAc/CKL0k9Rk7oTbn1nDS
EW/Mq2SjXUWJH1XoUDpJpQOT0A5wjPbd3id6kYxtC7R0J5n/n+YG5skdrqiM5LnZ
Um4ZP+kYxe9A7IEX4/7DcWupVyyYEtqGm3GMq7zZP0P3camYC8k6rb4CozXZ/3Kp
BxiLx4XXja1LRKjW1Do0M7s05rIPPWREb2ZUZlp22+XbqkeZWTIZe/4NRPS7QJUn
pya5kzc7NWwmGVEN8n5sXcQ5X49PbGR3aYQc3QWAWtbpXnGUg8lAZELzDMfmxKV7
NcpgR4vRSlzeuqI8jJwecw5rdSIjWRJJic7i1UxQ/fFsmIFsrQ1m5Cz+YgJHl70M
hq+ue1/QtSYUuooO+8YEwabv5sZxtXc4s9KCDdPiZYvJQc3glgFLW3r+jiYZxCCo
rRh/umnYWiMlOTm+JMRXR3B/nBh0soQL6hQNM+H8vYn+Z/WT+VDDPK55Aa7yiw9j
nnCmG6ksSzTNPSQvGf+B+icNhKuD2BSjirKieHNctHAg5LpSf8XaI29mbDgRXLuo
WYTkfFDWnVcoehRBrqQK4iWMDfuNZXzjeC1iAr5E9qdMUUov6eXL34q7ItEThI0q
prlEQ/JV3A7b8g8zwXxtKdy9M3Bdzj6HGIErZ5ZzNiunchC2zDnE4aRX7r9hbA+z
jd6YdyA0SvyVB3FQ0AFUnNJdG4eh5OTtklJZNNi5VV/2FBbNe8O178lpWTrR8qVt
S8Yw0/ZVP6DEDvPcbGhENvFLISl9/YS0oGFJ04pWUPFF9YKdRtVXNm6KNN/rcxHu
vi5GMh7HkvalJCgQWe1PzHJ2g63Q8FGqyRWPhXHo6EjWawfmK9pq3XxrDhC1QBhx
Z2vYkEO1FYJSF67FJAhdMqp8tpDipXa0K3JN0fb4hG3LPWVOEd8RwcbAxye+DVG8
hqmRDSgTI4bbZoOxisGMSxLCLrZvmvMP9c5hzAO9D04MZzIKDASL/g2nrjvSnR42
VQK4pRaaeC8bEFXn9RjKLNkYxfLw8nbMITGWa9WsRjmyNGtfs/S3nrfVmPGDJ+ZF
Cd0IIJ0L16CXblEiMDL6wpxA8XZgAzPoOCEP+N1QuF7gwlncV7XBCn3pnqklN4Vt
YTPyeW9hC9+WPPd41NxHHA4K3JF6aHNDu6jQbzW11NM/3nNqFX8EhsElQR6JibkC
/2TerBngMpHS1wkii1+TFlPCBC47JMCp9R4GARmf2griTN7eAfjZjMVgR5Al95hN
NY4GejjLxq75JzAerg4BwnyW5F940gZykzX0nqnX/xcJ0pkAY35xcTrmT9izHZGb
IYz2xlPzaEBz8HSiLK8AEOHIcHF6I50dNZIOx6HLLPDbqAgBU1xbciDAlw9945F8
+xTaZC0fQkw8CJ/A4xuhFsJIuzF6gEh3XP1Qz/pY/EwCK3Z322OoqrSqaYksR87r
WWrVeK3zivEuIeUgiJFPcmiJcL+rHtoe3dcA7OE1s+bVJSqsxJ7j9XSOYfZ0aSg/
ZOvZ2wSKH4aQ+t2Onk2ta5X7f4Pw/oSNiu6Er2phjz0nPvO3HrZSVZU+CpUkJZEz
V8GoJPfLqcWEc7Ah7y22EQDp6R7f48PqEFvWsxeOhFh3a1ml900O0mUv5vl9pg3L
fn3GxQfiCc/9TR0eGoQ+7Wc/zvjUFY7QA9Kux/8OD/5Z0+jB4hAdRyVf7y7D1XNM
68f0NLv8N3QZY1TiOZWmn5SCm8hZIQ9ejJA8r3mduWUc0ZNAGv4HMqFH9yLthZTP
HRAygMQTHNPPSLV35dM5NGTKRRHubBoljXSHWVc73zyk6GwRnJQWHTpV2sJuTuvr
NAiu1zZtLAytxrIo7ABiupoDmUtwXdJqymm+8JPOcSmsDJ0s9HTHJFVLwvB3F/fR
FZBSwIbnJokMCkY0yb/yARIW8nP+ioKDSs4MDptTSaU/uZMtHCTMoXXTKY+mzw4R
pKsJM8tOHYRUUq52lSnyL9ih6MEC/yosYfvw5cUAbOPoBYu2ng9BDSvSn72Azi+B
O3/E3DoplM5xN8ySwwxJQYfqO/RWAzOqj+eHtU4ur7Rv/7qAVu3ChCc/ylGEraXs
bl4NkWmFBj/bUzI9H0fo+g0P5zp+yd8afNz9ezzheDdmL60DwUCbCEyOn4NDFOiE
mmAVBb7MeVfI6D9uww6e3zZ/hHn52MO2Oqs9MhqRILLYlNfeO65K7GxNnLvgtOXl
Te+uL/FQ3a4ZCvNRDBub4igWGAdK8eUhIYiOoyv6jt3QsuoiwGaWYZDP+MxkX8kf
HZm97JM63e+ilPcX+VN9HyvIfI3r6pmUIusjrlwen8IWF4uPftiiD+QfrlLCLZw2
wWjave6/FqRn+e20xZJxyrlrg1Q25pLZCRj9bpJiMo6vN/fDCZ6DFErVUCgUDWo4
Ba2kNN8nBN7ArnKrbQ8D2EG0J8qUzVJ0cmCi3ao3qQldgDyJjPzW04pFQPJP2Qxq
Djn3b2bIjZcJubToU+bYiIuPDFjMQtxQYEhBUZNOa3fMyv/2hdU4DpD+2K4sP0uU
VXuPT1j1rao7prueJP95tBQ5t8ajhsESknzL+26X9CJry43iLKbxTtRq+QnXqu5X
aqMWT+A/kh9Cx0vGa5/d/gDcuvIfi7rxsbYyjhsXMVzFHKb6V+p+0zTmM4+HH8ed
kdL9/6jwZnW4NVFePvhXJmIy1dPS0vIMGWP1KE0N4UIyyDPgc5yzJcwUOIYcqtxC
BNsJGLugL0iALbCIZR2qtKE58GJPxxgWRXPcsNUVSrE9Ss+VtvR2BFXL7AdmRMbe
UdLNIvINHFJOAYfGz7wZZBnQUfIxfdGCWF9RtYys5eX7ynUaVHQng5YDwxU/zO33
/t/QV9CyC7dgg9I76hq7CR+CwbX94tVFONUBSiCPu+yHjTYPLa9sWIG6wlZvsT5C
zs7YWE05YRVXUfv8+unT/sk735KoFwWxQrBJYOKhkWuN/ECvGPrG5k3VLw3ueQPv
nxGcynOlRiL6gkUN75D94CPRRWMWpN8rPZGoUWRCGHOXQFxb2RxI/vRALmmwHpVl
W25J3/iZ+w9I2Q3SwasfM2x7hJm1MkteUvSuk5PmaV9lzF50CxTWTI/d7AyJhCK5
Fle9SKlr+3teLGcEGRj1PcysjOSDDHB+05DQZ9JvbGNlUpS4S4fbxApvtDEEx8jZ
XSfXog+T2Y1IET6dsjYgSJqzior1ruWPAvYtlKl8x1LS6GqBDyaYQUbJdvyWOsZ6
kGGaFboRY1EfxxJf7ZiC/kvf7p7ieXg+KsAt0jCB7A8YIBQ6OyHSzTqDMHcXICyz
qR0i4YmBFKaKV86SCARcxD3w6zxvHNMaPZf7tH1txm1mgZwzbjiTVHgTuFdJaiX5
PxX4UaiWlMMitTQ0fmjEZKd4AnjLOfmk0aJHaeUv8rpSkvoPtgXdewLpp+1/W9Jz
/5s6bxiBaMMLS1PFjpezFYoupY1CKXE6ifWwebrJrz6ekVWnJuI1Yb7TdFt8VOmm
Flk1ENgrvmwdwM4aQjAEtfKx0Q32cBILKs/couh/vAs0ZFxa+qBgsYqxnOG0MN0R
KoWZI37tPiYRMDdyiOMfbE+WtCHeHR87zwM4ALj4z9aMP2hEcXFinTpb9nEkXtH2
XDMXwFMJsvwKyVSEKsjuCjuG2B+m5vO2irY81cZVp0uJ+4Z1FYhc0mGu7FxTeb/3
IaQy+7HPBCSNpKtkLj4/rfOmuiU0FTgmkk9biZLMOr1pIDrJ6UP7h7edZG8bF1sJ
czhBHnADUNPnRotsdQ+QWtJkJJmMEUl3lhEN4zws/CnJfNXZ53K0oCrQHfnoMmPb
1daIvV9ODDa/+w2N0TgxLaQCqHWKWKIA92YtGDJo2bry8YWZveGMwu1FFi6eUwj/
vJNFb6TPsNocAcoTlX/BBjAqgQawoTCuBM1DVnhaTsRNdndjPM9pfQ4E7vEq2Cok
dYmILhluBcDDJQTqVSvG4V5fe6GYaiV389cNv6uP3CSL4NDrmc9WRCZ3Y5EZP++d
yAtxQO6d8Na45azGqhwdJ5FGBT+owqnTm7YuTZqKvU6cNlb6AmUA8Lp4sNmo7yxu
+cksAz7P9KBQ2jo+ic3Id/5ba6/7AzsBls4pDIfmbfboZFSIme0wVZ7imtYK6/y7
U9ErkMGW/9kxio6bZTWPtKU+31BB0L3afSpQZ82NS1ZfmoGC3rbQkQRJwn8ES1Qf
KNi83ZQHIGXbOVuo2pXDxL5+dk71azXGK5NNcMCo7H1fTbnRimsplki3kCr6xxIF
XAft8iL2+Dsr0jUzxBcK1ttmvElzNTwp30cw9PjZg8OzQ62F4rLYCMjYL/F56j/a
dGMnyjXge0et0KFRw7zrDmrZmL6+t7XB1eOgDzCqBPoj8Ok49KXuPO7h3mKegVwU
FrqwqCaycSeQVtnI0IPkPn/NfeZXMv0M3khtETt9RD5JLJEZWe5MGi+fks1cb8mv
ogWrrt3DHnr32t3XREWVYPefYUD4NEcjqmtGEoqMkBtqQU9KmQyMWZ+OXkLsWh1m
pFq5O+Iig26w4ewL+ce/lux0MeZfhuxYs8Epq9XCeS+/zvEt9ltubv1RpC4zmDEr
V6ozbgN0t0fipfmsmpOuKSD1BhcoBwRE4cQBXL9sz1ahGUxNmqxyUU31i5CauvOr
0IJ+85+KqSpQ1X+usx5J91gT86SyRPETFaV9Vd/2RGVxL4fDdVOlHEipSruxqKn6
KgNcLU5DTyLesblBr7xKU5h9fmRVvdRf/v0s8+en2H7Uc/jithEQFPWF/zbRCNAp
R2GjEZtL8u/Udrw+E7Ol32VrrNxWr9wjSiyynekjBvbE+YXrA5hg2JgpMykuz/mr
dfdb5eVNyCNTjzfLxk4a27sLWMO12R3HzW5+5dum0h4IesbRF/KJNxjU1Dy6QYP6
OlsDJWgNUEiF33B1L7DEM5RMlSmeBKqjx8KXqrA5FbQRmD0+HicVDzCjyNZyY49t
PsI88WjcPDQNhBARirHrBeV509QGKnG5JVHMDXRD7V9SskKLPONpCs5uRIrskZe8
m63gDkZFf2PMFuyd1XkZrfv1uVVv7spdA7o6s+BdgAp2d91tiuPjC/Dg2rlQJVVF
U6OAFnwruvvsC3J8PnGKnEQ2Aug3zJB9DPUlsiBXcGcHqbkoUROFC4s0MXyOOi5m
Bd3FB8AsOFfVNrchiyCoekgkouOplTnkJE3qJWiSYn/bw3UIYhUeojtdOXGvLvh5
PaQwqNpGqUgi+vmRHdfWUyBNxk9zqiM/8MORjyvdFdDLMkQ1BK+R31FfykoATJVQ
f9DTkKafItjY4IH8Qz8JUwZOpvXlzhbHVSM4z6Qs/EkuRY6cT++UY5VVLlvV7XT6
Bl1AEElqSyr2fp2AsVbJZSkGIWYB9jrWnyTPPqNW7XIc2ZVMDHJVk06QswcnJE/E
gDEhXy51L8pQge42Z6d0zArGKHHFAzJ/9fRrBxo17e8hJtAzuGJBkM6Gki87T4bL
ZtrAqqTfQkoCnA7Zn42nNUz4+fVNy0pRVap5jWDhjUua3EOhskXBQ6C49gByIuec
DmqwepZN9CQk9owHDE1FH6AQB7VHznLpsqXmkrCSXApHB+vj0mKSR9EI+wZ8SOyi
P3HyeCIs+G3toLRA1WBuZZsr0D6U+XQFS50/EKmCeJlPYu3RRK/h/yKHYOBWbDBH
MCHji1AmYIezCRdRgjNRLv/ftjLSBmtukttvz2+jf3wLXPp8YorzJYx2f72Tw6oY
7veurdqcsB0HfxRRhIXZCGVlS1nveZ9k/CmK+hYc3Mu3duqjzMZ8uKJA205Y3s7H
gMY8WFQgENL2P4h40gZvPKiNeiFnwmglU5GX31TZZwjvtdvrd867qNludVT1/V59
pW7gtYN27LMYUtzyJtCTT8cRjNNYUOEX3F1B2xEs7e3ZaHfM9JqIw9JNiu/ga38s
/VCN+Jf6mRQOm+jIueB6eLqitHUc2ipqOhOxgJh7JbDSMa2NGTCF0dgFv0hSIzHf
aJUWE/871KNEiZ9GA5TSESTUuK+PPIjr2EvFU3vgyDEZhvq3YUhcZ4QBIlORVLns
G5ZlI+oEmciPRi+qhnivL0He3OBWOrCBNDln4ueNcdC2vNi9bSK3r9rU5+VMWGAt
amwfH38tUj1Fj5bYfBJRVSW8eDyW5UE+QE6zEtTTRTielRxCCIBeZtXB5kjefOVI
LsTtA8f9YDSEq7QGc5/GDcdmqGJls/+fW3hfSne9b1zFLez2hrKhAsSAY+gyzwy5
5wd1MLEcxSmLDcM2bQbxAjYwSBnfy3ma8LpUc++b05JCGQNV+4rQ35tIkZgIXE4a
frVajrFeMcUQZgb5KMxq8VLjj1qrGPTn+Cbya5LKmBwNoLtju8FyXawjFMD8mdfQ
vlpa/X0q+n8Vho4YqF+EyGjbUn+J8mDUz+XLQIAUMbH1B41165JKIHszOCxanR54
DlOqOG0bbkIQ85JRZkZDQ1Tng8Bs9CAMhagf83vpAQKUDKYEaXvuqj+YPRDeJiyS
n5i3u/soPVLukqDUITxQGtuFxNECseC2EOO31JIx8gdBkkA6DI2NE2ktDsbePTSm
SOyJ0h4UAA9PHWUHRFh5OiRBSNm9NNzUy9xbPT3N1lfZWKuBGOiI+ce6Wm465k7R
LdSOvqlUfb/m8gLAYJpqqfZ6kbS0wCHwXlOUNEjft3khBUk+qr391yBt3X92SYiY
4kbQJwhwRFE+GOaH4EyztJtAo1yWFHkjj6yBHW5dSm+yNFXcfWV423YK1+kVjoDy
upBT6Hv9A2ulmDz1qzaPRmBU76ttWvmB9FnoHzSOT3RC6gn7qKYjlbQMxu88D3Dz
B1mKF8v50qblzK43NrFYSjUEgzi/EL2c7EL3lFpaqygC8WEtKVm06dAPf/pBTGYL
2WOqbzBGWqXQ9uTWP/M5yTxXSStysxwo81FK9pbYJ0LzH+Zg2gLkP2ZDFIeY0Bzh
s5H30AzOP7fZctCtJJ7HKHkaNfsH8CjgJaiWbsjPIDKrVIZq6K7gyVy2InhAASkY
3ufWTkgf01+OcT5GiYsUXUEMXGK/slG8oiLXsTF43r5EthUneMbPV+6ixFY4YGme
oDgTAWHMC1P+KAgpYmqYGtduPkl5sj7pP49for0fs9MQ8KxDIPxGSVRF1Gz/3wFv
FGG3G61LihGcT2PiR+ZP7X7WdJz0sEBhlxgm1M94aTHUDaCft5OblMMpAdhoC166
6iJcgqHVyPdntRZol9Y2OIxoEqeJftAKq6Py0iRDc9j8TX5otnzFz3hWcf+uygNt
zMXnutgta8yu4S/Nc4/LttM3hSxHit67cOd0vjzh69NcJ84C8YaNQlluZqt6gzHv
2uAqplsc2dQ5P0K3oB/B2/Z53wWbvIfBhj/hYFeOG4GeqXJHVJcT5AsJdQlJAajM
+s/f+iRuJY3PayEO2+/K7MTGMIcbjn1XgsvsdVST2UaFp+pTsnx6ltNVDSCGOClH
zDglh3hKWaUlvOO90QIHbXIHkOLXgH394WoPbobGO44QUTbPlw+sk++DhOqnNsmZ
nqe1WtCcf+HXJ2PyJjJFZEu1q2ha9lRK2JoZy8lRWlaGH2yAxt4cNwmiG6y8L5nc
bUz5dDdyj8ATOab13twGjqkomj+Wrr9OXfsI9jSyynu4+srGfgCG1k0re1Tde9eR
50LR8KAl8QZs7ALjn93sZuIdfJhTAAmopXWsb88kMCQ8UAZ1K4wD5d5QRUGeZVZN
QNCGQwx1rbdjG4E86fNRFgjciAEZtERqb+81WIhSOMYSp6NElxH64No1UXLuhaNo
O2LeDCZcoFnm2n9rl3KueKe+m+f/EN5nuz4PhjVKP/l8a5zRnrb6TbXI3vvcqktb
FMUYK115ut0zaRcAhNJ+sZzBV/K9s3CxZxUWo5tVhLhRQNhrCdXKFW4FTBGSaBq4
qqjcdmXPX7Ek1YnVD6xBCymAypVbtbEyOKmuRHEWdf9K9vHEngRsSGWD2ua+dSYf
PduMnnptbOhdEt4qQWWOiX+SoCWxDjVSp9SomdYCK7AjxzwqDM36uVuu+Tx1XsjW
FiW7HIZQEdkdSLueA3SRt8Cf0Tf+TEdo3PjcdONc8iXBfY4btL5fNrIwko59hP7Y
oVmqChB330JCSY+/rX4mDhlxQSKzA0Fzu/o+8ZRJbI30ZjVeKaO74JNNCTZq+Noo
HnQgB58XWdrf2TtI1SBLa8Xy5Zv7MHPMml1JHrjADDQI8CR0gn9bzfjrr8G7sNY3
f2wRW3FWgcuLbPB7d4xbXWg8ugZ5EALIvNhCE+B2vmyUKCBb42vxc0N/4aujKLFP
uBut0VpcjZIw42R596YOg3c2DvylsOUZPZV3vh1l8LkKrd7eh+fRGeynHrx5/vYF
Hzr0X68lZDVGh+YqPONFJN1pW4GPAl8DRi2XyOv4xD91B/EvH6rfKVp0sZkxvFBC
6r9iaxLqcXJ8w36nTizw4y9KB1JBv9YA4we5tlpr6iNeDvNS69JF3fRbRSFhNpIf
sLN3NO/Do6cdhJ4zArqd60Iu8987io2ZeiUtuO4Q7bDMrfMvo2grpINARYb30pn7
oAJJrIzy0N5JyrnxGbubN8U0MxEWWR/KN6vrpKf49hi8h4tPpO8Ir3ak9ySSHS6n
cjm3vEYXpnjfeAq/iLNwEpP3T2Z/swqSlK5bB0Jdd1CMqz2ib4dRH1Hpsjf9O+nc
R26bBKC1jTw1iWpSbx85UQfNwPGdS5/XqQGQNeooiVW2pAO+AWV6T0XqjEPcBn47
obx180UfG8TakPs4jc3sjomWaxieT7QtZtBTGK4VgmGhuTLzNAoTUMm4IFTjvFmR
uBC7E4cFjaTGeHOxXqD5I+3Cvyz0vlM3vJQ93hfrdoTLvUrb+nztv++BqTMGOBJQ
bjZFwzjnlcqSg1Gq7+qQVbctRrfAkgYZlIlt0sY4IdsMmlIF/r941eOglZG2OSBt
DlcV34ETmtBZRP7zIavylEFJ7e9Qr9EXUq2zQUGDeWUe/GQQRluGI1rNqZmpE9fM
Uckro/LRgW4U7UMfEmEQHjo2S9VfrArgXLFF9t/HVW6jKDw2YU1U2BOtJAaguUDD
IYQAvVfpK26qVuIMtwiUdO3FuUvL7YFj7xNBRmbmlZcgbUPRMgs6U3XWfliZyZtt
BMF9wGpHWJpPLx07wFP3C1l2k6+NaGRBmI8mRVDGNf/Mqnyb8PKm1UWR92Gi/huO
1qXRviR6iPxdDf/DGaLjlqe1LaJMHznUgnbEXOvv4fMVZZVg7e2+SXRdk5ix62Nx
MMaB3nTJOKL7u2l6UOl1LHqUMXO0uSh1haM22q9ZBr2e78uXYjgye2xppOdEckX0
8i9VhgEywb5zAMfq3GGpWJEi7jLa4jSGaxZD6jX5JGauZD9LgfttZbzHjbdPNVHl
QB/j0NeLTj2ImzUks6gdRMjY5uVM/144U2erSce1Tk/qW12/8ycc+KUOvjJATKrE
sxo/MmDSVg1XsyzPtD6+17toGhW5yNQzewCcrJeEFZjMu6poDwR4bDy17bas+GcX
AM9dQitFS3T8XWWpwTnocc2XOei40+li3ty2tAdvyHtsOcpX64Km3ZHAonavrYdW
e06dEVgSU0/TOkr3KrlQi1WjoH4/6PEx5aNZ8gSy++qBipPXvJTLXx6Zy1Uc37CR
jyLL55YifRTI4jy+7UY1t8I/ArE1DeUHPUdkE8eugzcCDSEG0lcYc4okDQl+/Nyh
rUB+GWeBDjU+zpa8F7QelXLEPOVJr+RB2fy8WDsO8o3MldQOFrgxSG0egc/Gd6OY
jjUdnT1Bvv1UqTfo7P41FejZ9B976skZ2iZX6m9bcprjgFiLnmD54MjSawUXFEfA
44RRLLDCMRfwdD4Zu1Xm87scZK9JXZCX8jIvQa/JkgYM/vf2XHXWeyjbMduMGyae
0IQeVagEU6F2ybfjWFkEkslglmB3BH4f6ko8hUU8SRwJEiPfMN8OUb82Q7eLIOeg
8RPt+QmGvlO0g5aKhHl0fBB4QsLwopcGrGpy3o2SA7CQ1BnrGShZzRmsqvzmjp3S
w/AkBRICaBxmgVTeu8xUCNJawAnbACMY2hqTowZlDWQXKUKddf7f455toPqLvosF
T2l/Bj1ko+q6ELqv/kv9RV1AWGjFTAlgiyCeD1Sv1X6Nq1jVa+DvoW2wknV7/T0C
5N80CSx/3IOg+cdCKDWzGmbfwK4uI0mV+Lcj9njUr/BodLh9n8dTPHUStEylA10r
KELJOnK/3F7n4Jid9AAknmnTygRVeN3voSp36suAvxO2+++3xn56XJ1UM6BfyMTq
GIwn7hMqiuKNEt6WLM7OCsvOwKNrMtOglkRqRRvD1jaSDmMbQ8/ccAQqR5Av11rS
mrR0gZ2zZAo5IRV9JD1wGJeYditSOEKaYZamF9wrRV9f+LEqK7H/qzb5U+o1jZDF
yNC+Ksh0i/CA8nm8MUzx4uuZ5JP56ACKw22ytCk7L6eWQ+AEw/M6yHCaUAO0kc8H
7F2m+x7LeTJ0mWPKbSvIFbwePpOmz8DUIVyFd/pP2yx3O+t9se8G+LSCW2ilzuY2
AOuseD/7T3UqS2O5HFDG7/7LBmgroWpCrzakMxHSHQoPYgxtIkx3b2UVulaCOI8E
dSEtWTvK4e3ywd5Ljvj0vawfPGSUIfmA8MCK//xkTwkBa5gxhVHPN+sUOlz7FIis
PhpbW9yGtikyK89ufgLmBRx7jQiptae9URrJ+mXoS8lzZOPk6Mc6gmHfg9Y0nLGE
N0jKgFz5k5D05eSrpAbfKYxmCM8RXrkbZt09Lp9b9Xy41T0AperKEOevfQfMGNRM
l/c0b8VBFsdYVyXG3qD3ke+w85Xxk9uHchG85u3rQnCbi00Dy/pCejcJYu2Cqz45
9XG55jqzfQqYQCHdlqAYj5flwpCanq6e3i8w52n9VFKmjBL2LF2cPN+Js6Vhd3L2
o2oM8wePVxiRkhMZDFklk+hEdioxnGWirPLP3SNRrVNvQT87x5pbgp9PQOzh3b6U
6+TxUCjNo1kk32qRpoExtm0dHPvWd8vuTC1bvQwiX13ZINnqi0w0cQJxv1Ul6FXN
ezjQXMhS3oJyUccHMJ/PkSLC52DpK58R9NZAcfGNGhkmLitWNdrVUa7fXpMD9iK2
E0gjfyXufXSTp3c5YeV65COe1GDf8vML1Uj3Eq5vtQRfJOMTKSWHUJ/hxWs4qiwu
Vvq30MfdaViR26F21KADe0yDMVgMBExT8E5yEFU/O9A3smZ/W4HLiqmuLtLKpR2/
fj4BDQjHfM+hjInAZryNQxK6r+Tt+R30wBZDr9hjnli9ADw7zAVHsyKZk1AGEumg
VvsfF6Ig6wfvofvGWDu7goElopsdTvLaBljHDsGvnzpl8YAouwwgO64ihpXMTaKk
7vGOJoX0K/ZadVYqBmUKZUscjUhnE8Hb1kNfYrMS7sF7sMPjozuYH0Dal9J1LF7Z
WncCIdrkvtCJpA6Oviu59YDgds9T9Wo642+0K1Uj6mbV7iIXhIg2DDu311if6z+s
9HqdINHfiLbKkZaD96xXtWvVf8ER5vheJchvegwqXG5p99FjXp0Us0goNPpRrML4
2unt36320UuzCf+5DCgGGjLhSpMMU6MwZomZn3FrkiA5pJL0BbbDB2faH6nrA5Kj
EtnZryXrlBj+PRTVGnBnl+ADB44RnhfpLd6SFx8k/9Gbb85tESs76zuCuhJpzJgK
BtGv2UghnLdXPadO+j5CTeggvBmH7tsU3vkPsnsTjo0UYitovkLQlYrIdMyAwNHW
1PMwLVv/bRsoQqmJuo5h7e/VrS/nfEeuVAyzTEf9/TK64p0C7eQVXgvZylIyuQTg
bunqdMsJriHCkk2Cs3hV7+VBcOUBHraXA1TmUkT4Yxc6GZEdT6vm0kGJES866tuN
OViRXbcErysUZZLyi26GCmR/wlCscTWhyvjip4p6S9n1ZYKwB9x8L3f0USuzqnl/
zlAP+MBKDRXUQAXD8TJmivoCnPyU06WoEGqGO38N3IdhK61aE1ATCLrYVo8GyiiI
4FWAUXTosoHx7gRCCNd2U3nwUDGLs2evjoBrsw6P1dbmSqXmNtkt9gMCi1skbpMz
/8qDGzWv4tCNaTI0YVVyu/7MdjZ1DObAD2dbae8A1hPiOQeiaAZUVu2nzHxFEH/h
h4PGOktnUgmKLzBI/JCjeAQTGyRPj4ssXJ0PimynV3m/+ZoQxWSc/5KUMNSXAZqn
HSNjnpUZp46w+jF7gIXdcLekvQoeYNNUHbBWBwtAd0vsnfFFw4S/pBmPGyOc3TnL
G5Lf60yeVQTZWfbkWX3Kip2yyVx0bATvarIEE6u88VXqaDo8ZLNFM3jf26DKQWvn
AqQrxoEFQFs6Ky7dpsYNzdRnBxjKfy2YyWb+SgO8Cr0N3ivsylaFsCi8KEbYOY0M
+x8B5qjop2rAyAEzXiVOl93bptPMuuIowpkCU0QUQiJnoPa1vvNsv6Fl+TDO3cXv
afq4L60ZjInFcvX95bAhRR7FkE1ICFX66oxeXsEZpQ6+ZatAqOe3R5EBsmwaBFB8
LBVPFostbKJeA3P7bKPSy56uBuLLHwwu2czSOcKlCz5I7nXSnGE2NAN1BBAF3Otd
mTjSir2vetDJo2PfX4oq+oLKGElHDtPIp9dAWpW5xqjVIEbRYyKKCYEFaEk4dhFM
pR7OF4mP6RZI9V9fksZ0H72MG7aPdQ32fOB8WwvMUXiWGeM/VGirJMiF95odOtaZ
1D+CO3oCBd5JAQDFNBdiY+DET1NSZZxlG2NKlQfbYsyrajOMgrzm+fa2tqTwSbbt
uyubg3DrG9yvaHpxed3a5aOA++FCeEdQXg6P34wsDZal8HGVeINh2nPHgjWKCTAf
0dpg1OiqM3j+1N1kT7SzNUpkYQOTnr5qF+poJpYa6niotyU3j4EAkJ9u3XAFOda4
S5m3kGnQ1GNIRi4ipyzx9eOxsNGO7gOUVNiA5mAeox09xvw07QEFOpWXlduwyV6C
+pFbWBPGSu1xh+yL2/TJTC0S1ye+Box33HXl7epghoZZg2mP2KelYZ7PN7wcmXbH
0zD5YfLrVfREkK1Z9S5RS9Zvid60pUNbH9lUHNzFjJzp/o9234GjrIq6ZfCWGV9H
McvI4lIODG9sgmSJlAmWjZkn6DUSuUrA0bV0f8JTutpklFQJMp+DP7FqF0xWd2QS
y4p2hGgzGIS8NINS32FtwQOtee4A7n9Hjtw+QWYd1rTwm3aeux/EFgBjl/VxdkA+
RLVuQbt+h6zWq/JFN9wanzi5Wl/mmaN2aVLyAXQL232VxBvC7cCAJWA/H5TV23V1
11/UPv4oP5xX4aEZ7D2cPeutc6ydo9oBxxGShwmQr0xKxWtAw9WqsXy7diEcasgQ
Gq5hizqtKNKRH1BDwwKqrRGej46RcMTT2vSyAUxiOv1X3IYuWUfSepwW1xz8GtWn
ROtWAx4XtaCcVtSrZOcgOZmhxIqFK4jlPzS8hnnrLqDVJjeqYFnAeh0pPaVPOtAP
8mf5D/lCOxYvkNrWjD62xHDiO0s3855dsTvRgl6E3U2xWz6c5SUZOy3TfsCv+K85
JmNCIJpOdAf8djyXDi2+cgvwDxmlwYYJ1xBP3Jei2bpCiQNNpfn9NGo/+hvQLxYu
CmJ1RuNUSL5mqqHrmf1P7A31zvYOg10G6Q41XqJl50T55IiAxiCNiY/zMuti82pR
OsoR8ZA5veLJQ2a+RZDx8VDm72odksqV5AFaZj1g7ETcF5EUjifAHFSS36MvvyA/
uOBoVu54Da3Y2WRk0xz+ZOpCEN9womHzgA/FdJXZuMI9wOYbwKIEGwSV+qRVZ67d
U6h09YegagEJwrlyqhHNMcf61NbQZv9onNNnNKLi2e5T41KhR6A0I1ZYKVTAJ46Y
ycMNXnZKiOYWJ/bYqL6LSyW12BhMonV2nujgFjBGCmJ+HpLza6v2moiATiJ1tpFN
FNKTXzrsWiFoYcrWvvnCEw388LXIdmMvzL6sNda6tTb/Fp/KmokLp1ZkRuskq205
wHBcvsuTfaI8I5ZCgRNtKcabpWzf7ek3R9IU1G95MSq3eNDwKErOk1DkdMjVh8bK
FLqN56SdtwHtLx2PVYlLOswBvlCM6YkZsfJAViVLP3zGJFPOFLt/MXMKq0ApyHgN
Hyn5/lNqpRdpieEANl4tFeqqAEJYlGVka17zDQCS3p9AnkJxlife79H2K/VFLVqo
X8tjYC45TfwbtUSTqscKZOsAu4L9coujuL+6SCUpyFs1eDplLbD5KrI9FCyesRVA
wSv5pzZiEyqtRKAEY3a3X1gq/CwctFMCVfFXi3QVZ8qm8wANbQji38RR/FxtUlzv
VxTAjJYo4MjnLuaEQUQqYta2KSczs6I8W+puWGtZLGyHYyHBEHWFu6uPTk31VXhK
LPFpdFILBJ/kgFX8dNcqAvFyewsLosCylhvzAzQfvG+Hlm40KJA1s9Gc09zhNydO
y3RdfbHD+SmfNm/OKjess2hDqznJaGmJZvLCx4r9WzT/mk4OafpFYvKtwCrk2EJt
9W42qcYpge1UFgR3Y9B20Bti2vtTuvm9Y4d+Q8WAb/AFSLa4TsqZcPw0ma79EaEX
U4b3sXuNE1atkOoDmvRXuavYYMX2bulr0r83faauKMeBDiKlc0QxPXhPj9hlDiow
tqKDeoPp7h8q8BnlFzRdvHTBx8c0SthcCPTzGIZjGoACBj2rDy7ZpPRpqaWzDMZI
be7Vl7WTLjd++Zr9VOnAuSxivf/XinpqChp12UdhQsLm6SRC/ip6sedoBjN1fp28
zBYt3sLj71lFW8O16T4M/AzoRljPSKbjQeMFD1aVtCh8EVxVLh4gGm8DPTyClLPN
kxkVTlfaQ/46M8C4Uoz+F1F7LZPKVLHw2YydPTvvcy0N+90ewBpwZ06uK/3SJi5U
9+ccGV2k0Tk54rkOuoIj6XO1M9nIPGj+OKUVMdxqIXpKSv527hNqooyT22DcP2oj
gd9khYM7xSSB+SHPdlxtFce+sNstRfkDJzaCAaXVDu00EgCkFSnoe9ELAEYOqziA
qt5e/FhxSp+8x90EgWlYAN65WHVCsY7ANiBr9sRR/KfUemk5U/LJaPvFOfKiF+g/
VJjy8Dl4SUlGq839FE08qJR75V+qgg8/4CIfSL6VjtLbj36ogcS5bLbY9phHOrP3
9oHa9WdB+khEp/yVXJbTmpvqfrp6RVC/+DTnLYfFllzc8IrHBXl1G+DaxcCnW8p8
hEIBjpwR1T59sl6Rt2X4/6a4036u+MWYP3BUZ2xW0B18p9+Q8H2J+RheaQG8fCoP
by0XqvzLrqEP/rSh05tlGzPe8YSkKwHXxT+tSL2Y09OPCiI9UE7s8laESlEJmQv6
vaI9QLlsaONnRj9VNrH49iYQzmPvfGjf7lCAp5NTbupczTmDcetHixrWTQeXHg8O
8Jg0YIcdoEMU5pYAq73/mO0VzaCMvNU4KUcqSwpaYxvkh55EdMwPtaoD3Go5cscz
92qR01bOJGPN2bACg8E0Ix32ZE7IvTrG7obpirXImDwedahi4Li98kOg6yZOsRhF
cxPwqoJg9hPpQjGLkll7Du2CHEXLkvTaMEKnztqn+9jtyU2IB03DJUxo9oYx3GTT
T4CKPGVblyFT70dtprD6auBONI45Hc0TMX8nvjv5ls6z2cpKNfnr/sTf5yKWQwxF
YRKEwRaQQHvMw7JzcGdtvB6ktJ1+HRAtbjVfDV6uWOKnDLiOBW1X//C+hQjUl/0p
oJiuLJErt5Q948g1AY5yClDY5lakToFG96iHJMKSIpzH6C3N/RvVwrL9NNxQzpeN
SuPdTUkZ5cS3tZhp1xnOLWWOEp1FxG9wQ+ALoj+fikQXXCkqMdNfc9W7GecSMeur
otAJZiIxv6vsIch+pqzWZr8Hg/SaSZQru6MNuOszTw7UnucOO+cvgJrFIwAFTPSs
nsP56uUfH3/IxMLkVd5x0kU6PY3yNWllL3wIq1r5Qcs12TvOVZ4kvUsWeuVY5uT4
Kev+MZJ53x0WNVp30AmYLQlKT6rYLcG9q9qYKIIUcO+3K6Fk6xnGhGq5iML4fY5f
56+sgl3cW/73xj5zQQ8Kk1y8PWL9l7yanfMxEU74DX7cSGDBWOjNZKy2t61XUxdp
KzZ8hbiueMfuWWTGG1YuR4N6Iq2FOSIn29rqkhhPslxJIhjB0PAAjU7RIb2nvrds
LNF+YZRCOI1G5b3hR680iZmjbZqPO/eVJEARdo3HPK1W+VDgHsbfT+k/QEQurW9Z
LDBC/BRKb5p7GF4csFOAxd5beK4CRyBvvOrfwqkQiOhxuYLz9AusrzrmGMTe7u2R
SQwYe+pQ/OWemo/mZwHc1NPDoRCUatnVqlxHrjYzfyqVQM+Zs6eLC4Ublelj+zRB
+jvF76BCoqTEmG1EvGJsd58TaDvxaBI1KvknDL7IARPAimBcDmjjt39veL9YzQVP
Yomqh0v2PofXCQgPT3ad+uCp44qfYLOSfDUjgxWx0YKO5mEojS0orF2WaIagu6VL
d4H1aOjJ0us5MBELeFvcfgN8kUHz9gOrtR72fp0rMjWUvOs3UkLagdtIPqWduogv
HDVYDUxSyNxD0ayQePhxos5UnvAGpkseczsM11+z12whI/2jXgJ+1A5qbD9OIl6j
QvxA5fou0tql7i1yp1PM+QnLibAAvQy1SmobcFLRTVDDQU9W9rpsp6mJzW26M8CP
KJmAS1PybAMCe0r+Zy96JyBjeY+e+jPzu0T4Rza+jI0HMCp+LiKueARqjC0jwXnv
S8rCrdH0+Q/T1mUVePZmZNVh/0LdZBkaiYDvfUfamBELDSDyyZflMZ2Rf7gGSOUU
0onhatrPFmsHVw68q8K7NZcu/7j5aqsMQO2D5zhGSnxIM3AnheUwvAx7Ix+NMh8M
Qi0I4+1i1kAkLHtE+TFsWeFKj2oeoh8GKpqlaGPxL+/s+6Dg39wkLlUjDoWxtsbj
OmDurpp1gxKhV5jvZpIVZ5b3N0w0c+8/Ev32y/oyTmBmMiNKOHgjkyBoZQ3AQ8jJ
qc0k1PyH4NQ8wqPVgAIVlRLRGEzRTTvCoupjSKUKLaQzsRGMk5f16MThhunwWSbh
cZCy74GA1QK+TV2gNjcgp2Iwp2bqz92kfljo4kDg/3V4N2PFz4D4ufXI/E1Fx1vf
0ifROle72MPpTBhhEZU3oaJUQSO+R+aaB2OL3uqDxUXlGcNYMqzaE3dVtF6o3lMZ
afLWsiVhK2DHxFt/IkQTYPoTwWe06URtSzM33Od2vDVMALXiRkRkDlcCmHHh6c/J
bApKd0FdjdG8ZU5M2Ws9eEWUjrVzskSiwCrbTnzeCAXP772Jy+bpl9cyfNsenwqz
rBYP4jpxiX29hFL+Cf8iU6ntoFrbJQqiy8ne/9/7eHz/Y0iuZqgUQKABJYmroe6c
t4bWiKoYsH/CYRT7VmDBrq3prfiJNmrnt5yKr/MWWfJ+P8lSDV3tdZ4L7LOnhOQD
v9PuAsmuILe0TCdCaI42smmeiai03QPFmT3VrghgvilQpfNF8JZ9DQ202+QNQbpP
/g1iOI+Y3MiLLxQBnNKHqKKXO4kFWz1aqISD0lFnQmBG7Ygkmsdbn8U0ZUChmtFH
U7zNLZomWto2si83LgCHW/LRVcqeIV2gM5S+ZvqFrfxMD4XPqJFos7SSv0hhYs2t
mIq5xyxMyjrh2F1Xq+4LeI/yUsYqdTS51vy8lFcnJ3Nas9nAPXobnrxEQOV67S4S
lOBv2sdZXH1ez9S1ZMmYRc8rti1bbEYWTXJw7O9+AO7NMEwazn6pAEE86Ld1lcUj
v+d8rqqg0CO9n9ou59r/+lCOwPCtlRzyNFBpFIHONJRIIiS5H/YJe3BWMHlaTqqR
BqAzOFIsEN2oactBWoLWJNd6DKyDrAjARp796kxNmwR4uj7QssKgNfAvbfOuZ5JD
z0/aJyfCuOjFMMT3oPgP0qpnQJ7TqCm2jEUKu0GtSsndVK2y41tSr3YMNsIuYlcF
6jtNrLnlfrEFANEjwAXiNFm/VwlMSP+lYOdO/TB5W7g+l9zge1ZnYy7xsHMLd/lc
6sPQc5vBYiYQivD9sLmDmQ20fqeONjUGRsUmfOOAguJMT8cgKCcdyPGWiTSWflh3
qKUkKyK3gIvqehK2kAXYdGlX4dTiQ36G8M4FdgP8IJ15MsM9dZbajs5qCaLhO8Mr
3sBVCFFseWUwyiDsMUsuBA4LJ4Ho6BxVPdT2Cd0ZGklsXBF8XWQ4exC7R04K+FOn
iTXETdCXO22YU03AbwvGK+fp/V7AvCRBDdZdWA6V9B7I0clqW/6f7I3syYLznZEZ
3MfPXrsNElGod9CMZzp4P6yOfla+6wIGTqMV89P2VYGUDZm0M2uoGR+dKnbfvEOl
UnB234ZhPBuyIPPb0s/F+PLTXBXjc/P5hsOwywMQp91N749J1iZTQrPlE8f7mec+
LOXgLazusbEN/h/so0LK5horc3cz7oWn8WFaNHu3+WbN3shXDNLu7zSVr3bHM0sC
mNtopne1TsFEy5DFbHiYmMZNpA8EgQZqtq+sbCdSFWv2NMDuPmweNFRYdbowgBEG
li+t0V++p46tKAmtbE874qPKf29GQ7nkyKwgFnfwGsGQyl9XbUSZuVWIL+RKsvqZ
ArONPq45wH4A/7/NnLXyG6tlLt37cBdbeX+FC2oY764T8+aWofzpxUryeKJujEbJ
eo++jmqC5d9Hc9wL1wA0sRIUukAtaMSV7vJx4zBjLp9vXKL/560SxCtnAQ6tYdWz
7WG+mH2W63mvivE9IB2EtiyTlRK++LzAT2K6E9UodpsnuNYsJ1hqDM1ECemoJq7b
NXZBZkhwCyGd3jHaDrJu+nKGo7gDbTsu2IQai8HJPOe+iVUWXcco3IB3Ob/M8JyC
IVNo2Ix0rRhIxqhWQw0GgPFSOGIzd+KjZxOVydyMRpP7NarJc3DW0JH5a9FolFH/
r0/x4syhy7iZpEE6D3cCfhZihn0f0x5fDmST5O3h8LyAQbkZvwV7a++dNIZl4Mxr
HZ9zPn4vCwn3SK7DlMs+c56OUcxSpOF392eCoF6iKWruL0vQbwN9W2q2NGbjcZFA
BqogSnHG3BLmP9r2vSN/uLtFeYa0iwobuYJcJtyFGB731ZFtepL4TiuL4ALkYQHs
p0gB7NaUpMTJ0uZMsHUvwavXSJuSPumCIMxWRgfgd5zGlGVD4tfoSo6RjL+wwIug
g+NcxD7FdFasmY7qHXsCyJa4g49QZ9aVQSnEA0GlgClMM8eM7+kPsBZB/1jLpxUe
s/klQnPz9X/SAzzFYaJTtn0/i1J5ED8z34l02fzrIoQkLh75fxxV1aL3WcqCTVK9
TK5+QWPiZADIaPnH98E3dpy5T94nMiF/0+502xvwkG/V6OG+sshY6K+ZDBkCw2iU
zQq/g0KOjuKMWIB/fDhwq9FSXPHd6QmwBdObqh1CZ5uXu2wJNk1O9tvGUP7d2iPI
eHSwMrvn3rocaObQMkORjupHDRklo46PNHlhmlhQ7aZUfIlJrQY+LSTkmaapBP5d
wTTTWfRA+oShL0U4QpSCxcxMWpo/NgemNCi6uRcHA493A/WcZ+biILvK95p32PXO
2eR6FKRIMYnZn7ZCVeJ/vJXW7ohBwg6wRyjGCgcFlJq/+acN+unowsP/PukxNR4D
9VKXzgvI0e911Fp6pJR4g4yAf50gF37M+NgPMfQa4ANEhpyGGhuAfYcK8wwpHFIN
ZZNtvyZnWLRGM4elCM80FNIjF5unKb5OL0zR9P6+/DkgPCTXsiZ9fSgGuTVMHgfl
fNdgMq5ivMMF8UJ6FI0VrwPtElYyXPDca+HpQvsOUp0ZCB87BBka9Oo7kkwLpM4d
ZQRCKFGAEDytdqbq/jPy9TI9u8Q36pZflndvR/VHRYNGCDUQE5o+WOhRC5G1MUgY
KmpOXYxlPH9Qq1N41MsA8p0oXO5Ck9iM2bwEzHyn/fOkepBS5J9dSR2QpjG6Ghd5
zU0subpUNrkZMwE6pY6t0egnRtyL4wTyY6VarGq+vGHLUlfr1iP5pGTU4DWpeVLH
J3J90GONbQAcfUinjQqcvD8sMVQ4tnueAIHAsBGJWpRL1l32h0gVgNT2LRgn2AeV
22xD7Mj7DOLUh3+2cercJOvrW2yuYMNR0ZOcVV4T8ulr/ebQpdTTInfXBAdGPrRF
7uYcAipCV2fsFQFonQrP/o5RkoIoOGLo8FXae9GsaRGKVGRNNKR7WSHjzfnc1jFz
01krIWbkPKVYU2j7XwMoCeaoR3gGdVuSr+uAsSReZJLvNgR7kcHJ4BMxC9aZQX5n
h5AjHfq34YnDVhl+1i378jDu5O1IIMq1k16w999cteqzcsf1qMk9Ay2leMw5djTK
joYUyePeAFoiLG4Lt9VqsiARkI+HZZlx5vIfk2vlVfJbqQEQo7bH9/gQcvyzuYeU
Cp/w8+fCRRfwD/DPYxQkGtouqVX1kOmppDwipLC8Fx3TzoKm/fXsBA9J/AIJEGqT
XZryjusMZLjVkhA5nM3SWG6WXLsfD3yoGyTM0GWmTEiH8u09V9oGWKXvLP6BsMJ8
aJDzy2zTUJOPg77MkDvq/IciBp62hyM78wPoLarrAE/2F/HL/Ubxj3kro7BM17IL
A8DkfXitqu4/si+s2nR4wxeyKVGtstVqu0wN0zCObCl6mos11VTlpenWzHI0bwVh
XvQdzUjN8ZhpwRb6oyssg3XfxQR6gZNfjqhwBja6kZcjONiEu6sopqIkxZv8b/zG
xiRBc/BkRPMbRejO6WwzSbIbXqCMJjT6JhHtEEAxYoCbdfD75tr684Ss4Z4fyWmh
A1co/r4ocMv14qpKDX3+sbtaQ8EXkLpZUKSRE7IUNCWnIK1eYiXhN+7EN3YZ0jxW
oUXwesswghwPauej5Ypurry/CGb611ccbazZaEYDnq66CiUiUehr/gtVBeKxLGRm
9Lt8g2l9CKrxr7H+kV9NvnQsYLGUxed7ffwHvrIqLyYimOlrM99gtZy9jp38U8kV
7wkTJTkUnLt8nH/LVA9KU0O8bi0DfchCiKG9yES9YRtOoW65mqOrsNArPvslRhH8
02FxLRZVnOC7pGVXW4sUNtme0O0eCZc9rdwgYJKEY59ClYI3oz/+SLFtLOfwF1wP
/DGpHKQ79ze7s4r/yI4/f0dzLjBVZCF2k2F2XKtWutXH1A7RmfrJetq3mTPjHGtY
pddbT4DK6bDFQxPnO+oogJ0jYeOJiJGi1zGNgEk7Tf0C8lSLwyoKPrDJ0B1vdEZD
AYvdAUKoj/h+rawzRqNrErARbRuwOUAqrz1mhjp0C9+Xdo6q85NlloykfbFHvTAW
294bsX8DnjH1GUS0vaJSny0A25g4iGZvbf3lbdhg6wzyDtPrXl2WtYvWsW6Pbcmr
LltCB/eqQlP2sek2uPqGvIr1RqPqcP1K/VhV+4sVyj4QPX04tF9SE/goKd4ukmTg
5daQn/WKNU/ujOOkZ9/Qx+Dq1ZP17k30YABnI3YZLJ2lpTDBRgaEkNVAG0jVBSTp
ygJEdtA04I3KYfBLTy3uVyQKyBY93HpDiHi8nGXpAJCfNyuQh6B2XS3NBLpLGGuf
rJlleJ/BqsxuJSZO3oYvODO5W/UGalSuCgepLD5HeeQU56/kZ6uwDON5VXF7th5m
yqk+qAZsQzdkR0AmkrfkzRN2ZcMiQfRTy4HICvZ6ZgOOrC9U/oRLrqcXGumVjP1z
odrA+HSLQfBy+xnkEaTpHxZZlDj8nNwy61U7Z5FqckW3aYa62y4+1BURycBN/KVu
OaEto3VfwWrCxvSX8Bz4aPcL587sRzvRHmFQPwMOVZeUuCxED8QvJyyHQpZTHbPG
9WtcFI/Rgk7sUFnM/1AdwUMEitXtXfAokkVJ9sm7UxGVlM6My5e4PyHh5EoLrT52
aCgykCaqEhlEaYWw5s0g7Y6xputTThiHjTZZA2eAG1R+nH6oM2TT6bm0yHAfoMu9
dd4ziYh56xyAX95cTtsymtC+W9jGktlpGXJepX+/sqR/As2fzGusSxcmU4U89BoK
6nXqAWQQlsjuXRFJgFsiPELYo9hJy5Wq5wBbN4m7BzuvihIAy4FKM9QmUnWZ44qr
SnKMsE5kaTiUGNVyB/clp/Dw1FARdujEf+d9EWgygyvjKpCOuhseBDx7WKuKjpks
o2onFcFurFrXsz1E85Ai62TEcgEQl56K4taPcTZ0npJsy4757QOntIoOWRE1aVuy
YafIEJt1IhE5xc239NSjBKofVOxHWIjpgbyL7Q7On2Cs/6QsBFpvwg4Lt5u2zi34
TU5AvXzus/H6PyZ5bQ83C8Vm/KPcZd+mgmruZAx8b8TICOXzEDXwnXwhWPXmu+9G
iiorqnigaI7Ur1WxINIg2G33St532cxPeH2CUAqQ6qtIFpRkRTomnzLFJ2CiW2e5
8qRqrs3WBDvSelMcsRxkTZDJaICFSlgaBPjOP5BTcZMgLxyQjm+hSCWHT0GhkUa8
62LOnj95nOOYXHHIfMki17meDmxI4lFtOf6kJhV4sYgLy904BWnXI9fkExC0O/oy
2YsrR1nwatHxjtF733XWYzF+NWylinlaBakiyNaddQo6koqQo616ZTXCV6vE08Yk
fBqNMXn3/pwI0iTONneVhsZaK5J1O5f7tvMw/HawmD042+r3Fz1bbIFhPW9B5IQ8
bPJeNC7mzsdw10v4Am0mExriVH0TEzbLh3CMCI2jDsCflUAIpFyH6ryN7aW2QLNW
XvRQmvk4xzD3Cj2/QuCFzB3fKryoWxp8f6Uu+16HnvHN12tuc1Sm4QvKuONBIfuW
cAMIjzGMs1FBvTb9SpvmSxHHv2wA0pVKTmzWCn0CEcmdzbzvgDQVrAkqFMna6FVL
TYMh2dhAdmKGkXNgTwH4dNyvDlYHZxBJ6Vf7wzslaHm1gn5mRO1c96P5etYRa5jd
OhKEBIrmFHVQorU5WVbYgKp9vuf4oPXS3NIwh8C8afzU8MnsbOHf1hrNakXrSKsa
A6DmuqfSvKuhlprfjBfyoXv33lA3qaY53gvhCoPo6L7TSmotG4NW5LY4mY/YFF93
iiCrKK6fzdjt/n7bzKuiHtMZruY79M6LauGQsjWVGWNMx7UDm070yExj+y1gH4AL
x/lOxk8C/Gq9b4I7pQRsxqwSMrUajznRrQ05t/FUFv/pdleshtija1IUs6fZy3ek
AENbiVZ8QfpNOreLffNSi1PVAUgVaLaA9N6GN2kNHKcAsmZGj3690TJDA/+Hl6Av
pVKKi0c9mBH8S5ZZdykkB1hd3RaGxTln8n28g2I9cPFeCpZciv2YIaCqBhVFljT1
41zNuCO+s53wJ9aW7MA1jiBmsDkO9c6RS7mJ5dZIUBZpjFT8RIaZvaJuLPfZrUWY
6rQGJ4+UN2Mw6TmAvJdq8rXAp5eqEhyZ21/8qX0FMyg1+pZMdTkPRb//cQuesydv
dwyrrjY+8wRNV5WpnWVnDpMVADhmYk5+u6lAyubEFRO2EiOgTFpBjscDYek+8KNI
oASWrxJ6UPnUfD8YISKlvwkmqbNwQpXcc5Al8wURV5HFziMfu1q6g80rKnqWlT8V
MPzwwJ1uTZdKdcpImsmLHGwRIO8+MCGdpG3t9xfVrry9p52Y6Cz8ivf4dOQcqPOb
YSZIi0XdUBvWezp9HWoYimeQYXugp5OFEVJwSP4P2I8X4LOCb8RDAjkRVVQdnc/s
Oh7i+SbCbWIhwejhvxLUHFBFIPkHAh9LWft6BWIev/xZDyO69NC1Fs39lMwNlqCH
7ZVGlBlI0OL9oAgU9uILhxpkq/cOxTnvBE1PTZi8P5VjiSyb5tx7Z0WBYlgCLQPV
shjGkMLiCQoJqfwWFiyjzvicZpQAoXFBNOsL8Pib9tOm0AniRJbERuyEkQfuvAOx
Ja73kv2nO0dNF6G3FfMIx19658E8ECtAOEwq2lXloe+nHhXJUrsMMgf4H7Lqxohm
UXYU9qcMahvea9tt0FVfXSqitO+yNFtiejeYMzqnwM/CvrxswboXTS9Sr2IppPqB
+uzIskK2RJb7BlWEwZYPwHXzgnD1+w4mL9/txNiZZ/DFNDmeW5YtOCVjfgs4or8G
wqSTwXHkVMfcin5PfD3ouS+1d8EopkvnI6USayjckk/+x0k+s/XzvJqOp7YjlgoH
hH16wbsPu3o6xf4vN+jsEk5oywB2cWNbJvMy92teP1Ym8VEvtAAVqJOu7nf+TchC
TUo5GlWiCc4hQZjQLZvK3zdrIPHLRZndKRSvRf5rfrurN612DGhb99YGQU5r/aFy
VMSBwjhuEJ+T/manKAIE9yugd9rPADjrwdnt1FaPAyq2GOpTRffnOC50yiLGRp4L
+xPocjpFlsDBTJBKerMhrtkANb6DRA7yvKT22hQ5v9Ed7EPxuwSILys2+E75gxEW
7abWBJ9K7OILLPXC4bNueKSdk31ae5DjxhjEDGb0pBwYohGy6ePrYvMvbkmZd8Wg
ogPJUeBRduSLx7kpyLAVpJg0kNgI3EMWRGDTwJO4Sx0SxYIAsmHA4cncSJz25HGA
QuA+1+uTGE/LdmyvOd3dl02BLVb8w9sykbDB/Q1866ByRtwdy9+Az8gMXHaI+BxG
VaXGlJnMgWFxNGWGD0paKBPX1VppjVUJ0C5hKsuXCDeusBPsrZ6ZSjsYiGquA+13
5SBfnDgJdXzbPhdzRo9W4AHVv8+3ZgGjsFIBvfFiwSG1A/33Y4qmIx/IgvbEnwsF
sRvGTRV09rDgIrJShM+17cImBGguiwB5L7Kog5Xc7f3LRe4mde6BHhrYt9H0Kh/d
MQvF5mCLRWCn/2Cjem8Y0UHFY8WZO45ZVyGyUCR/bSKhrlfciOPjwqAbQ68eHzIB
grm4YMkHJzBmkp9WIVUkLucx0DiEe1pMOW3r/5XjF0Eje29s5y57OZhbh191lcgE
MWp8w6kPUf69KOFu73YduJ/dD53jdHkMliA6V/BpMPQu8txv/Gg5eNYX6OqnnSfd
ZmFpbKQmtxlxUUFQ7/Io9UY3iWeBNL6e4DF8B/rZGFsg1+Sppbz0aQ7lkwBys2oS
7+yFNXbV5JzHEXqlmH8qwGG7uIb/WEqhFObwinLvKijg3MgYzDaWYuFX2TBI9CNN
LrUBxWqQOfp8b1HcN6mLTPGg0kCh5Z4xs8j1bs602YsYdexQ1O+YuSzG1lzAZQUI
sdj/WavetcRGFgoQOwH6u/yoAzopeAOZpMJvuQp/BEPxh5kZ/pPM2RVBde+yj68F
5Ab98Q1BZfDu3FHyDlwDdYLpFKHqCJZGKYzJK9Uk5/LFxdI+iHWMcCJ1VllOoRgD
8vw40NrYBydCndl0hl1dAHiCHcECGHIEjXnxxr3FEOTVqrkdbZAm8DlVaN6sRUNm
mmuQIkoYAMVgHY3Y12G06D8LF48pdyQQQJ2GIV/8s6x0k3ikFrtoQiVAeifaBOL4
JBN12dt6tBrthW5n8RrgzzNqZUFnOg01Jyzm+E8pjSQMaR6cNp+eBWQHOXY1qzL7
MoHbhXI+NU/gNvxlC5kDG6ARLfoPE2MTjwM/mtoqT3d0xo9BQ2MLwEFw2FYja6X3
cF+jgmDlyoafpW6PmyGauYFmZB7RcoS3nizmZkKgUKB+d4cDjDgX2OMJCpIf8Kdl
Aj2tLIkHzE7v6uBsTxf+epq2eoFQDeJhHH8XCcoiuYSesDI7LvFyY3Gvtvs9XxQ7
wnt6tEwyVUkCtwzM5G2Xo2liaLAGYhPnRCqGYt72AHr7VBoTLRgZRd8i4SkkRKD7
BvvfraX1DqZ/6E9fIzIvxgFALiC4TIo1dOzOnFKSD+JUDVF+0S3XIuMKYQMpu7Xa
Y/kkph4FnWGsSedfrBeELB6epf3Ik0ty8HJOe1ScVixv8fBgLbrUiDPv3Yq5C451
riZefPNH7DVVgYuPIOifAVwy1dwc6muXOWgn0cWy1Fnr7s5iu7+KDZeEim2I3H/b
qCxVlSrcAd4WZ2XSRK+JeL7e7/o6pwXsn0vd4Wizb4lfr18pIqUIwPDJcAUUxFxj
0pMkEwiHhB9BILJxB7+5PITZv4vQ1Pzr0JMpmm029cBtYBQj+pIxSSJxQGWG0k2G
Thor0S00btHEEg63KyDFT5cCAKH8SWO1HwSezKYuxXmVAebjPVruydyXk7u6LWHQ
uJ9ds+4lieKV6QxUq2JRI1Ql0zhjwb/r2Rfx7jGO2wY4xCB59n6prBDWZiWfM2Cs
neBQRjgoQOXuCYuutmTmISLnbYOAxhpsdV5M/Oo2kZgyoCiLAsYkOWxHaJ/VwpHY
0QYDPPlIhP2ISAE47ThBtmmzJfJEMFC0fxll5qyRZwYXN1ZOHVMtauoZKff+5KVg
rOwHE5/wII2E+PFZQbT4XN+AlEVA2C6qDLS6KvcwasQusZ+A5BdwiaJb0rRc5obn
G5o7RCimbeLl6xaFNL/WDedF/r/iRNe1GG6b6WWP/5NS4Py4KaHCV7J3SWNa6+j/
YZOfY2oxV9N0E7Y9Pm6GyjO9+BRkfk/WRsVhwcXEvirGJ1IDwRSQZgQB4hOQDrqX
Fbwhr34XtdC/Qc2VOieBbsz9HhwueaT9j5vDxNw/auCH97c3Yn+8hnf0gUNxQTHf
F06NNOAM+pkfY6MC5Ko5Mycl3TnTIF14l5w61szAwGKnPmxOh4vrm9rxwYunFqPE
JLPeqmsD/qYZZFWGT4/WrH7VUfjIq+ZY24RRIr8uCKqLovoZjfMH+53xIerTwR+2
rWj0WF0CLDrUwHAausH4y4llxkdiZR/QExgy41MbgIc50j72K1/hCfhspmF2txL9
scNULv9I2nD5SpBvGb//1yBDZvaGL6eGPVMI5m2uzCI2nT9JqSGNEiJTMaZazV/P
sXJcCj6oxnnr5mWankA8RXmtWtwyerjhc6p/SadAKuyLjkco1EwHd+xOZLGvVOMl
GE67zCgOg6y47I/VGQnWRLHN97qLvfsCsuxTXuu/Qfy1KfwN09ofaMWDWCFu9CAC
eaonpGINaL4CtA1qpewB2o4NaV/r5qbv/LxUh7kgdHacQwtKCCJy5kOW97Ds1Euf
TUaSZ+FokXLuBOzGfBRcm9x4atQ/PFkDCfdix4BJj2qRn6okeW098kPIiBFmHfrk
hkAqx9umSrLlQ8CAcVsjJOMoyNPveQ+9z6z6urH4/ysn1QsaJHkDZkvz5TVLt6AK
SGW49avvQs3E3YMKmtosrYbITPxvPsXOAUTeKvMKDV0GPAHblPqB+7/Nsr79Dxxh
H0x1zEk/Bitdo7TSoDmwg6wODGPyEwH2xTX2jnUbfQiL/tSX50oyU92fJjEo+Qs+
7vxQw4GEYf7YYJ0zimQLcvJC1dzZjfzUoWOPo8eNVIJ26VYCXbsD8F8LCZjsskBF
FFIg5v0ptQds6Z5dBUQRPUx3AqRHHK9JgCW7SvvY5XLCGbRCdKbmBJgGq2bueQif
Zj8IvIZpkD5WF9uSCLquGCCkb232/VXOOspc+1gHjjnmxF1wbyoN92BTnpWLtfgo
XC90W7qf+LRVIK9mJMh2v3l6EjE2qB0vlFOS7GWEGcdpZBOrtAe1cyjaenZxAzSu
LTd77tFiZNUzoIJzf4fP2PqM9MEKIf6zdUc1TsoCa4eJHjGJKsX1b2dMxfRnWpkX
EeCKX3NQTV/pli5/JbeLSdlZttsJYvCgpGeumH/hlsxSCrkglpdQZ95+hjHmMJuI
yjbCIly0KUR1WPlMcC4ISDwWx2dJAYdzgUUvkJNXjUajAYB/GMfZwQ8j3StCk/YB
q70jXFFbMF38EN6dr9py4AK/hEVi3666DkwWD9LiksaWC1to8kQ5RMxe93DpuEhs
nEZi4tUtJeO7OnXK9RvxMtbauHklWljSpkXICohTkUhG9ecyFZHDnnAC0ECo+Ahz
VgXb9XpBxCmqOqdsIitdBeJtSWgy4ZW9GtZ+F50SSbAUjvFYXEg6g54hzuk7OMIR
qz2GVy9SupFTo62d3eT1TfBPkCfb+3rVoXHC3pOICw2h4RqG/GqIeHyLwf3JGyfI
xxWpY9OaKDHWjHfp3W08ZamMA7yETF5TjNYgsQOIoLIopg/b/BN4QJLNmIatssmA
TBEDmQbU9lfEO03OqNmfoGjISpa4lzzAoTK4S8Eww6Ya81P2RGICK758e9ZuGVUO
4tyop1zL9pvppiYM6S3SQBvI/0AzaZvFymX9EvvuEeQzIEECqRG8RZlhXjKWWtlX
TDs+fGY22OKETSjBFkkYOI9cTlhthdkFnv8QoJKMuOfnuxLEbE0ADwq59xz3YiVe
dvdRxJGLaA49ElKqeOhlCgTsT6EUHg7PXJL9n0ZnV5gaGjqEz/bgYy8zF2TxUkOD
YvHEIzK9AtF/D8SiPv9Om9DcKq9qi5HHLHpaki2lmGeAOvvmxsXw+Ts8Uw6p/Bld
ErraK/rf33SIcJup4tQVQl+ugW/WF8Mu5paHbsMeTRSOgUrPWcYanqWu+qDtEyPX
IUEWDOwMyPx+SgkaxjXt4IfGV5FaB4pAe8VPB8NA5RgMn3lLNL9xR3Ft/nDvaM01
la6/uS0c701NOOgXt9cvj+Yr23UhSOLXv9koz7TVLZakh2fIWm0KT2/VS/sZEWmV
pFGkJaYLAwOqBuU2Z9XqN4Kh8/1JwlOQTPLLsj2yTDrOQ7cGyoIDFl/Cp8TpB8Gr
tXL6L9EP4Qvpz26NsNpvT+XTOImlCfXcESKBGikXv+koRloegfbo8Ire+V6rvESI
u+ngYKkYIpiNphsgOs2PgS4Hh18hzgcmyH8rzPs6M+fSNwYVXKmrZ3yDcFFPx9bh
IcfSod7shORsLXTLbskuWUF+8rLRqXFUz62f1bK2HUGwFIVSFRA912+5m3QuU3bW
ND/RWQe/CruHH9ooE5jsoRL8hLUt22bFy0OGhQGYYWfWMyuN6BMbJ+/MlrkPgnqr
thAMlXyR8GBO/ohIHBkpj2QgTmWeEqKLAOc08OqMv+kfe7NDHGlIycSM6BRmMDYy
jy0xd/QyUP4VxdULGMWCDiOiG/kq4x7rdOQOtiwU7WNHA6SsVeOg8mvdOYm8rT8n
0j5SJNSb2Juh17+x4J3I8VA/zxEOYd2xRogL0GDQJfDEIJkcw7nT1/LMIY8WIxGJ
UmcXC8iZMKfIVi4XJy8RAmvtZOoxSR62pLaAY8WjFHDS7wt/x3VKcrgguM692Vi3
JJXAqv5qhB472ARiu4O8uA0eGe5WWE8+GQPaN9lFi7eSpNWqAgVjbu17hlZuS9mZ
IlSgrClcet5Jecs8uQztxC5ZNStjh7QKnYlHzu8jc9KCSE5ph1/+h/1YtKdljEp6
vaVufmhuRt9O86ypbMY41oD3jMFFd7CQ1jj64XGZSGzpeBuNM/d4tHMW1+ZesH6I
cwo7xBFd6KaBmAyr8aWKaYlxuACO+4MAI2IP7aymdohkuK3X1KFOV4yrF4weo7va
gCpICh+coDkNPNy8g2tobD7JyBQkth84j0kUmJZdnbGJyY4Ru5MmBwAL/Z/ZDZtK
8mGo2pWCUYPWufIwX5q5woJax/umAa2iy0C191hVtVNLD+rbxn7m17Qcglp3OXjr
oNmFoda55iYb0eL5IO3sNJTUeyPyJo3YyhiosfqjVFmWta6RPTqYw8/bk62vi4Sp
QA0qXRWb0M6ukj268eI/rbh6f/w5abaHRPomGAVVL3ewc+RgrGuPSWYmSZJcB5U0
oKrSXzRB9YOKiFGAkEI588MDlCTViBWCCaLOnwnA895WE4seezhL+vlWiWDf9Dl2
Eavo68XoWXAvgvdEsy+pFENuDpUBH9Alg8Ke8XYKNVvLgL0hVRswKq9dnvv+8vzN
jxwTeSCOlBInGnVstIhj+D/Qem7zTynj4sP2XEV3bczvJusm308u3iNUiNkkEq1y
TA693VG2l0sFzgYF4U2CV7tpE72Rl6nlddEBnUDnTZGhFpgxR2tEIwgFqSBWkvmm
9gD0iTteAj3JjsWVjsjtp1fZQxVMIvpKWiiugLcuQVmuZND9PhPTzjMzNBbecvbV
8WjDicfimqq3yQq4L8us8QNR9qtLxLqHcxGCjEhDzIgnZ6URuMse45MoH4aINDvP
AB8Q/g8VV4SScEzvWY0QgberODhmIlYoax1acq/V65/A/uVtJkamqK7EmTkRZRv9
M+V7MY+YUC9+761zuLN9PLXE29pOXjv1/Gw0Mird6Z5/Aa4IC7r9it5HgPRSeipU
oC5bP7LJDqAwH18FEkafcMUUlXk9hN1MKiipIHpXrPnkbKVhLuZVW+tZaWuJqDcr
bFE6cWIFpXz1uzYCMHWxk1KpjJq3WNDxa58LozaFcYQ1DT6esQRSeSWpkFp6qc7K
1POG4kkiZB7bA0vQk2EN43jzkalxnJn/B8gHBhjRe70MdG1Tx2tWC9bkylzA8Bmr
o21uWJInvvfkwbkgEusmcbZUCeeMrsT7jwoO7LWNtFYH3X2Yz8WqirbjVawzcz+S
oTbw30S/fEOJXYS3ElmR2AOUEcXP2WTG/P8nuXoUFlmZxHn0H2ImGi0T1CKS2kdw
55YcSgN5CcW+4NwGOluHBamSqNNbkSKg5+QNgyjJ9S5mXGzvyjUMUFis9cZWjewi
7b21I//1sCvtcxbzj2lfoSfIn4pisxF44pnHzG56BFjHRi0h571q6OM2ePueLFWn
8Ur545WPwkISlDid1dV1CDut7rBXC8DmrKeryk2Q38bcDboyIEqGaV8tf8D12hJr
/+tfg1VbtAQnJR7nt25N+bUymz0sGu6pN+UamCl5VJSzw1DkLFkUp8FQkel6BUaG
/Kl3YcJvTYXxo/rusTyE6px38K7vA0FYyHU3GEl3mpI1esgjCCW/u86yeHWEtB7l
8bzTrN9aeSMJcTPKUipuHF7+YJrcZC4j/SflZ/e57afpBJQtE2hHp2jyc63lkokS
J9rHKr2hOUsARfELz5hpLowzrdjsUHqEiYa6Czbinft6ye3z5ao9UT/LqH+p+ZM9
uUNy+uBSoyq5tAdEqwD8em72yGuNGuT3VPUq7cv9gNwMnPfGSl/E6Pbxsysv1d38
JwXchPn7bT1V16gkTBpaZZaWnACc83jbBDeCAudOQkZz/CZuq+ppJP+vUrBjPSUl
TvG3/g9tJFcq0XL7l4kee82vOeN1Wel5it/sDKsZ/DvXsFwMyfOTOc8nmHk6UHll
ZlSy3DAUFJ3xpzghX6Mgw6CTtQxUFCNF7f9/4yi8OWLytI6lpwip2osym1Gdb8aO
8WntS5deRjaUNDwI/v9dfRMSkUaW+yPFoH7VQ+O/N4oMpO4723Z6e7FYiKNR3N/R
vj6ul9xKYARGutuJkL7MTZf1uMeA/Y20AydcN7Vnu6fYS9H8NvxBRvLL7hiqIhaC
R9h4vZyUDQLMnRe8H8AtO58FFvRRCAYFSwgW/9DvUY2/HlLsNl85VtyLEyD/Gu8A
7HRyrYLH08oagcU2mngWoNkxGMzGHrB8xu1SaPvL2PUBauYmR3+fLM9BiEyJKCVj
o/m4JfcOZU+4Hgdp/4KZDGaHT8aIi7X0f2Wjtg90eQgcXeMNeiSVjVRyIX6O583L
FJ/0Zm+0BAFI80RshFxXsmmXdQS4OJbpXEfY9JtJVW7UCyd2FxmoYMG03ZozWap8
VceGKPxIUYARgLkl4bljdudzSYMaKQ6V4Ao91pvrSOiDIyavBXVL+kNuBxZjylfo
0pdUHiZt14xjcDzYU3+FNu1RePorAGec4x8YK7ZOt6PhtVP5C2Pk24hFdasxMMkS
ZAjN5ARKcaOBPL20Me77SRnEEKLKhCIih/a03VDEqkuL2BNQggf4VRiVQ0fNTIu4
uf702B3+2mJxSIyYSFy07smLTIt5kfuZXxjawlpXELsyd5ncWHlQe43Aky/koFo3
WsHfmjE1u9XOxTcwzwy1bgSyHGO1cqkMSN0dgAbTi+OzAz+CzdZyPPwuM4ObwkQU
b+ar13x79ndINM4A6Jy7aqdWN52QiIan2wg9QXoOMKqPSIbG0nRzyfHBuEBl0C2M
3Wqrr2S88vriKFG+tDN+lW/kncPEZeuzwe3IpY4/HS0iAM1L+631q8V3qUKMwnP4
ZYrQcQwZnnAWFQ16nASzdHfTaMXeWjcGLqrgbR7FZ0MZZgx9Q5S/h4TAOeIL1XmH
Kikx4ed6YPS7GkQStB8+r+ohdjD4LdR2niKm8hKQ5iAV2iyCHhhKSKKDUYDfpNsx
YqZAOUQ3eYvU1LDITUUIcgmFoG7FpZHFEHqBys4PaxDvphH5eOiPoDU5w7G1QyFx
LaD+U7WzErDzOWkizzjsqVBbcdDNdQsck1pyfrSNjFfPPM1De+N/czqh8I2/bqo2
Rjte+wqZCwaz8FMmDS+lGQi9Y/pbQtwavg5OJ7amu9CVymCAOpzEx1eMWKjPl7Ue
EqB2iwOPVa4/cmT3QwPEjes/00GEU+oEOZtIP/hEAY/6q8vx7ejVjlUbTVQu3i8U
n+lBlssS+nNwY9JyoaoLQepD5Jd4zlu5vtHhJlFJ78qeZ0oeJ76wv58UnBoTXGjx
YMUtIEVCyq4o2WDABD1czxYLf60wTBYW4obQXjE8BGW3obkjBdzOrtfh8yKkKw4b
Q3aTGKBA6mPI5XytQ+PEwOoUbN1gvqRkR+mFefy+w+nALUKVXW/sDpf3Gqv0mXIp
+7953GZh2MkuECM6dZpyLeUS8V77z0zkCofuvDDmoeKD9Ko9GCgt+pqyN3pAAX5w
EKAfK+ghJwzEFmxs86dknQ==
`protect END_PROTECTED
