`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmbCmAhXG/X0IF+UzqONRkShhCo/YdS2/9U/5rTcIPWn31hGxIbaYF5NHHctvVXx
eU7Fs6F3WrWKjbvVNGpghXn2GUzx5EwbLjqMf4iEUR9b3ChHRZakHjEAqstQTLAI
qVTrEP+QUMHKBgFoYurWfMiTv9ODp+lyqDjx4QGFSTDXMj7YME8+mDdBDcF2LOLI
56ONJU+H6WTJfeOzG9xTWdfb5FCJma7kh2tm+4rYtmLUEu0/BS9WEzFUK1NF/f7p
41G4SCn+hKMt7n/hIre9VWAQqaH2f9bkxYcXo99h+Oc=
`protect END_PROTECTED
