`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+iHyjtRNm+QVuNFO0Wtm1zaONgxudSgMo+7N2ymh7NeDbn1dvp/dH21dko5zXKG
WVQGH1N74GJSDICXRxB23c96UxaL9ADaSurIgiVNA/jcDjs8V+flbQ32pID48tXB
f6pbs5oM1GU0KlqKGOa0TvPNCzUFhqAHd35bah//PwE+tuDJzsTJ2DXX+TY90FZT
7JD27vKQgo6V0kWo5eV+8DCHLW7A38VE0uGxSAIluZTi1MEzxZsdLKBImQB/jr8u
+BuCs8KYtDNOgJMZDptjKfI/ipGXkMwZNxZIoHSq9W6xdYWGxzfyfNpGdFa0zXH8
u22ylCv5t3+v8255LhEW9COX0OdGgcC37sA7pJvjlLEuV2rKLF200w+hmlml9Tm0
Xse/BSb4wrxop4L/V3EiRZgg62721ayPE5Tp6f5+fMIbjx+U95VhMiBnDYZmqT85
HWTq1IYL6Awy36YaN1tgAjd5YlKJw5cG7v2pzYKYk3biJ4hRGs9Hs+mEeP4xBNSU
q8VJjhxVpxqHGcG4b/Ngw4KFcvGYNiKz8XRk5lBRoNpfxNdJFn/YCADll8WL0hLg
nsmPkJSBLs7ckQlvVSpW0g==
`protect END_PROTECTED
