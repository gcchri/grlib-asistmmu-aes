`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JOcei/WsZS6+4se8W9bRYP5QHg7DXh1WQcv9MEgpPk9yUYu/mMkeG0+HqQHKrvdd
D1LNByM/B4LCn2LuhdhmTlZL8u/NoCRxbDl0q6wWjqy8zTU339RNLyng4qGFNdlY
QcZWSKYgqN5TB209HrcFM9OfJ6UpYTQ2BiHcFKBnDLxl1j4EBA0RPoi9QQV46QQa
c7VxVtg1YiOZTz8ct2dRTz/W7eLJnrw/00ccQdXnpTOBTK5FFrugyoqL8w00tzRH
mj5f0kXWLjXsoyTqO1j1700ihVh5sJuBh9UYKO4uAQ90EiePY/1H4qVdscTt5xMF
6tKg4Alj2BfQJgeplwn2CoY0oFkyqobD1GPqcpYSI3hjWqCf/VDzfYOozztEQ5G8
PwJZPpZE9CJ8GWrZVpaNqtJZPUVc1JmvzUwLsnfVaS+ZVVcr7TvTA0UO5PHszptu
UgndfLpL9kCkAhHN2L/YWRk/rsIPARQ52SfU8iCWClJQEjHtUZLlp1VPxYpLjy3r
lNmE4KH5i07+r4Rcd8vDD7pr03PuidwQ5PSe8ozpg3ua4Y7LeCecxYaS/k324iZ7
1M1hkNYrvJCJ02v0sreCmUM3+/eP4HrFZP/QTBd5bbrXMQZStyYNcgUY9Rkpmrp0
LZZ85nK2rpPI+Hc8uXdtwA==
`protect END_PROTECTED
