`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0X0dct0UbZiOj49Krka439DKtCFXsqOMX9b0VuNOmOViVFWCHT5ibgWhjQz7JoDc
RBzJcJp/QYs3qOPjYeYa7yTxeJRb1doDAmvU4yyIk6p716oKQ4aQSy4C0g5W8gqy
v7cHj2Q6b/g/8YOxyio9ajulZGums/2yuJ+c0GRvUf01zQL6LA3mFCYQvTdTFapu
qpsHMvpJ8PyMoYBubTXrlOCmUcJfcEr9h8Nh+X2j2zxFbUOk/6sz+xUXmIjI5Xw+
j5BYFlfuV3L/6WEhKx/1TyhycpOLfzpv6uvIcakNidv5XBkDWnyiHN7PWkzsfAoY
ZcNVLjoYvF1EMbXmQEhJlKjW7RUXrPvM6yDvtW0f2Q/fUHZL5FNMTQG8AnaSb6yD
baS/pm423/SQfxQ5vAwAdrp+8lZ7qxANlEmaTG6VjeTe8ZlwEESostBquYKKnIOo
hIorBCWWRoQmZ2t9TksiAURXotinlElsSUVkTFAPIc4fuM6xO3SQRXZHVs6pds58
xZMxYLkI0SGmwOuaITEJNV5adHDlW8EpJtLyQ95OZ+dgvvWTbhCRSNLnoEuZCgDP
ZFTFJ8AQNSVJbs7CD5b3cmfuWHfs8uUXtxq+RlRBLmaCxE9jh/VtfmQqNo1wKX+Y
ZcDzh22Cud+9qspVt/Ssq74b3s2w2VALrofdT19m0jDrVVldOHZgQ/UUk600zIOd
KzX++5g3jUXE5cpfzlTpJ+sNaLoMjB1mrnUpbFhDZzT0jEnRql1dOiLhA3/OiHjy
To/tVu33pZ4gCLwcyO925X8De3qgcF+od8FA72BUDjXRrcZj2eS3dWxmmlZ2IDdY
vbzRwIHAQaUARVQIOo4En/n2Wv3m4UnANYw7sB16qvD90jWxZR/5D5D07qPJVO9a
TBzmjKSG8FWgdtALIEhW6XIxFniyLT3K3ji54OyLZyQFTt+P4YVIK0cEwyU7vWrs
DbSoIermVkQBsVk/n8Pk/Ealb0m7Opb5Wrms4PJN+PtE83/zioDC4tg+NXWDU2E6
XHKPHQvttG2eRSHAS57KSpdXxeQ7cRoLZjpIU09w1WC+WDSTxzg1eDr5FkVK661g
LNPUnC6rO28boZTF/k1F0BWSAVctjguqNI4dNuRpB14EMI4jaQBaRSVgBtqSQD9n
VoEemGp7Tu0Cvj6OEmI0gAk9/yIzsLSo4K2m3Gh2CNZjWljj7nEMlXVIO1UEkfnv
fE6NbwoFAXmc1F8bzMAlgndvd4Xm93aZcV3z03Bik/MuI92aAiIit/WVeoSMywv+
A3M83y4WBcffyuOVxXNmXOnx79qm8TLYzL2A2mrSjEXFiRaX685vSN+/0E8cN3QZ
K19xEGHaEuxZKkSDFen04DTH7o7zT0iY7uNAUSATOb3J4LIs+ALMniVEPKRZ650b
1VkmTroQ5L6VsCwox8gc7pRGFr8wYlUh39I+NhV7k8F6tNW0hdSgR1kkOIJ372Sq
APGqJ4f2gdfy74ADiJtLG1eTEXwoYYflFkg5YHP2U5laDQgPmCRUXc0m54nnrdsc
klcZR557Pc9SAjQhGXjqtLulDb7xbORLW6DJ8KCPAL8KBXbpj1agcIfr/NQAVaBx
X7zbtAnn65wIr2PdQmoD3YCpuhOmwtx1Bfpk40xSulLo9vk3x+cB5g4DjAMfC16O
x8vr7fpbEVXgbTiGwz53Vv+Gp+ZbhDIpqtUfR/6GAOv4s10uwxb1TVihl3uF8xjE
ZR62oxnnpw2KMWC2PoMse962PV0XMdN0ZSNxuqC6BdJQMLNrMpxRvYqqDWY14Xg6
M6k3WHVENxGFxBNKyHWB0htdDp1IESUj8hi9O6gCZ6LDSF41UiE6vOqWSbzAS0e1
jcUzjAlmxEMJ9fyhErfZqq4FjJBystoDKgdNCg6ylqWdK3M8P5HV9YngK0IfVzKD
gtqkwdMbFa/WijwQ69I0pVQs1lIejt6fLdOZ+hzk88oSMIj5Jd+5aDpqTPfgJL0/
/XSTaYvPjZ78+q7UH4y5Z2aegVqBYeBZ4G0ksMEqobubPhy2607Z2nrYTQ1iM9lF
d4DpLKTMbLyPNH9EaqSFq3PvjBFmMI1ApqXaRqOTMPWaf0fbcOeTjMEAXVmK8gZ7
lUWekBQQmGe6nIH7mhC+vEfXfpxbZtF0aSx0OKtIBDGT/08vNj0s6/dIbCsRI8qi
NZXkcV+XGywF4o0FGLF5Xbkc7dRfA2s0uhNZviYIJJjhgan+nZDq3Vba+viM+2Zn
4Q8MvCOQVHDBaK3qrWA97RXMkBWYe720S4Ac3F7d26vY0pyEyEHCOksae9PjOXGa
OksByUwhGCyCD8EZIVC3sPPLtBc0nQsJVPFAtD8BtAXrbPJD4yWeMzuPxLub5kBU
vwJCcv281JQlpx2OgzfwOcpxzYpqeY+UmOMSsDwSK56CFE6YT3BXzk7baE8Ff0oR
OM0P/DEcGq9E/AzSqs+tqG44FVX4t5dGKXH/ZPC8CEi5V8W2q0U5XI4e0QvV+k+/
DaA157ddudezzO9A5VNXCDqYmf3Fo1nC5CgJF4SD939aVLBQRRMp3hmG2KWOZtuY
vHiI73LVCbajysCxJK1Ypizcb5xWWaMGZXMfBEnZf4GpywwBA0z6j8uASOU3nEyL
GadL2cRjhQchuA9616uNx8aCiydnwhw0tGO6MXDIgyXIBxNLA1WbpCz/rhMbhqEg
f4EF71fNeYiAK+P4swRGv13UR3jsREkBcEqQxBz7IulXqm9NxvlR0Cq8QWajXE6b
4SALPVMb5qBDyA6Ue4P03v0xG6E37UVEXsPuFuc0emCb++RL8e4T5rfvq9n56BmQ
qXrqChIM6GAHGSo9SFOZRtx6uZOP5WzY19XHOgUP+73pOtZIJvpLKTvLx0OZS5s8
5sP/blHZioEmcxJxIolIm0MHsRrUXlRAB9SJJPyIMN94UcKAu7gf78/QxejmBPoA
pocFXWeT1tL2TkOsYgB7rCV/OdH0ADbWhQ+9Kh4cJ6QIAht4Nas5yWHbiWHHGX7I
DF8XM+SsH2QIlSAlrkzz045kcRit+6xwtIb3kVmd97KV3wdZWQiVXY/WvcsmFr8W
6jhUK6beKxd8swMQAxZLQsY98dxHiJ8Ltvdgp7sivYQ1BU+5FQcEvEGYDetUuMUv
zEp6E8Zv2bNYGbUeWkH68EDThNnnxcH130LPYyHisq6Ot4UchUOUjmW30a9fYkh7
dfkKf/2KDQAWLlxiLU1xWMI/i5LYumM1KA/PJeJdlxbXYA5C6AIAX7a7c9ZKtjOt
+CpJKgwZrkSEU9o1/RTKNjfHcUCdkgJkd2YfoQs3pRnja3DhLL27RftGAXtZ/yTz
GvajQzfE0cknJWAeVgjkPYmz+eQu0YbLZSTA2Nir4fmCBGHu7sQvARmcSlHft2tw
Oureak6vrHpaShwUpQgMzFqYFdxCYB8FlxD/KlIy1i4My4somtXFd1iVJWVJzvRb
eUYHCB0cQU25vqGTSobK+0emX2Rdw2i+f4kxay1pCDnoUSA4s/88mGv2bRyHYINi
slu+M4ZrwYneZrC+GTlu7SScahovEp+q3yoHrOTO3cKrvSHqXelSUB43OIHmmX1I
+hpH32rqdmh8E/h1rDrhse2xocdOTnJyPfORaoR+tQI1VtCbl51gwGdReUEC+2sO
y2KvW6Tl5AGcMnIplfeerosaGze6I8yW6UPXKmaOGn2cmT7BTiawNxoDuqD36MsT
XOd0vBj7JY2ERpL99oj/CeTzJf7/1yO5s4sQU7I0m4DtFwlg1/aYuJ5zusBwR4Ul
qJYvz4tFAMsbnl//dFhdfiwTQLEdfizPxNDqt6uYLoktZznSRTwRMPJH5dGpnX+V
7TQTf5qmbq2mmgerkIQ+Y/d0LkntCzOU0huWHl/zzC62fDLWFimZ7qhJGyiAUVds
BjqCcn9ttLQqByxOH2arkrWlsQWPdxwx3DV5jsI1oGDjHGLaFsUAodSstWTUFO1i
ksW0BaX9SrhZIHDm2vYiU5DeTA8ssd/gfIlg9nw2FFXYkAEa9JROGOoTKg6e1yaO
HcxOVdCBNLHJN3gseGmwYgOFUUscHXTGDgBvvnjUtY/4u1gJ6EkIBqLvzsvFUXxF
z3w4J4OO8n34OdYF3RRSCFb9MGHWIl8rJOO9EgSJSucFhUNAeP3iYvnTqTJcnTrG
Cor3CbnzM8BiXRPBYmvxvcnWCpyV/rmjMIieGjZAx8G1xJ2UKKiH7MO0BeFq9Fif
Hh+NxcyprxGMSV0+tO/Y9y7dUN08Pf+9pQepl0Si7uTifCdiEQsv0kP/u5XtTeGD
25Cs+WwBWt2biqQM//WDPLPW6DZxWTGrSPTF43QrZQI8Ao8AjATvmdTeaLR6XiAL
c0MaQxwIXn90AHe79WWfKDJUSEq1wYlVx19aDmsHJXDPML0B1oXh2Se6FbjM+AIl
zjnZWSb7gBfilVA7rbWVhLAUmcYFxsmGAA5DRiaKxZ7TOtX0CCsm3QrZ+PBxV9Mz
vTJFxeMZPHqdXyUvjhXDh/vEF1KuLlHTuoNx0d2+ido8fWv7Rx+chxtxH5SzwFsB
6o4BLc/tzlHYi0Arqu8lMG+cQVSQQL70YGd9TBtnXo1mjSzNAy/aomu3Yv8xn7bN
xKNrTgAtXJXLio7cLKLGeq4C2fYb9LsJH+hvdXxZwsE92pLVY5OeDx0kCYWHYsFZ
JeBSRTz3z1fnLE0aBNQ36Z5mIXevxh5bJtB4Uj4R1fZ1apKLqqDChN8kknbbDxr5
poyEeRcqSvGDi3CrfJAxLKjfQh3zAJEcSPepGl1634pyN/Rl8HmXQ9qfm0XcUpGJ
JQj43C5ZsFI+P+Qd1ak/+EZI9x4kMQs+SrNpve2Jym27YdR0bstoOCxLL0cd9rbZ
ezengyBD3DBAAlNxbrGgj1WkyO8ZHWLR2PCeDKvO5ErWjYHhrhovmpRgxmpeKo6o
ejVxFYt+l0vXz1iUGHkLHbkjmrGIGVAGlfSClMniQixDHE1E2/ma2zl5P0gIHael
TV10tlVK8ZjnVumGEj6Fsrhpib/bZpIJQv2Gm3e59Q+vgUSfo5B3IRuB2dZxoc2B
DN0qPJSagUknqUyMr1BxDtccYK85vCcIwy6ZmP2xlozelWDAUL5RNdHyFv8btm4L
DejVYL2SCE7Xnbx9pKwX4v8nnMs0wHPyFXw29qGbA4sqP/BkL6UWqkV+VODLuPbF
JxST5yFE05puGxWJLNfRp8cR37g3xlK4yn1gZ+73gYu3f7hkxixBp/EoXrmrC9vo
9J7HyspV3ZlTnhwjvRoT6oimmQsRZdjMlm2cHD28UY6oa8g9WVtpd43mnc023aRR
slnq1REKOPCQZoQibwNcttTHo4izRI+Z+d0PGx14dng+IDClx6bko8OThi1OgL4w
YxJe5Qm1po8oszki34oPjqO6Twa7aejlGWjjVpnUSSBYWfMuv++8a9D3oPRfHy/R
ws/HbSnZtTJUcF6Rld3QkeaLCYDsRGJHMqk1llh/mSujzUkgrDdniCR8OZjSAMe0
576rk7Ps17qM4LMCGQKtmHDH5y6l/7C3BAwZCxRZhPG4dBjYTPsfL8VogtclXMdH
vdCX0yK+xaptJ5th4zsAAL0lHnTARtGQNZPpVIOfv4W5f9/5iKv90c1jpKNfVE5o
6F8B9Ht9ilBeJYR8+leNErbhqUxw7CK3N9ZDQON/YUL0nHx3ACGIAc7+yyWZ5zr4
FApPh3qMB/8l8NKT3FkggqDNRTTq7F5NMIiXuen7ZHemn/sasN/UDm5CKL5x79d5
0HsSc24Gy4/CTVY0mESYkOUpfJ2oYa5BLFctcYe/WU5oJOGfc9t7sHbSOSHymSXS
9V0xAWDW2SQhyMayX6QOYysPJ6FD8E8iIOlADm+pME5w4lCM6DQe974YeICgZ4G8
Jl7gIk0Csj35s6WTAch7LoC4m65t0Oo3u7pGgg/Xe33cqxF70QgK3gjB4bUHZbWU
TRqRs2AQmu7H68YVq2ipmEnln8Ea2FT/MHzSxaGDr/tmFs74kVKDzeFQkAPrSJYk
4CBjGbC8A/NA11dKLl9gesPXWg9kyEXsxEVB2yI4Pj1EKOibjOWtUMLmXrJsOZlP
9Nkvecac2dENsh+8uas75KPU1roTasgBV/O5vE4nWXh5fP18DnOQrH+wI3d9kgUx
ifkRDDhbG1Wsydt4CCwqFmBGKipM87stCd2CFxWiS/gtTC41qTcaEWCsmZ1C1yLU
LTEdYFgq8BEtKzthw1MantkPvb9XMG61BFyaHnU+tgyAE+mlfkmp4UTUxjw4ufp0
HlJR5trNi1lh0MuadulFhSdpHhJPLYPv1mXIRlUCICOEDK1ynaWTdcS+A1gvryrd
Ml9fQYXUnLPTbu/sFPtLNnxY+aZ8awFBX/9D6CI1dxd6gl1i3BKHOy0vwaKOEIPg
rhv+vsQKJY5YLrpH8DznxblyZ8PjIOpelggOLArZfJytLJlRyF/eA7hbGtpiiJZW
9QtOTL4fDJNBsQEAiM/t9nFRyvjzf3hjIAnW6IDZ0LT974X2JgTpGV+cC4wAKW50
GuVFNUJ9pfceSA0DhLlRrau2H7ZvtUEGxrhVHmTDiAJoGvCSU96Yo/XOpGAkhBIi
RB2adpZB6Qe2PU/WPUPS5kRwme7EuuU4gJFENUkm1YNL5+Qkz3xFwE0hgu+5MBdy
mBY8njhlHRMwBfq+McWQesaIcmI7fVhdOauD21ApIAYu+po+qmgfHrn05twEXaJ4
cLDfFblHjyuLy3Rp1m1hnBjCP1+LuWh+yE6LJEuuaGGHkv8xfKyxj8PxaqqC6FWR
LAjcptfqunpSsM9ajmP5UmtYTb3giepCGx4632A9A20T6IF9+EqQhqo9cWCdme6V
JGSvkx/UJsXCcM2alGPWK/7RrYsu6Fz6F/9YDcl507K4AsumLivbHVapfqKTaOaF
HFzpCNHWsMJu4038D509YX4YZWxYFqY4TqH2Bpd+7n40J/UtLCh80bRAua2l0mur
PpL0dyVLHBDZlu9+rSfBFFXiVLL4KCDhDl6OubKqz/L97+SnH2vPSL5XmnSkzKDB
u9LZZqxEBUyRWY4Bwo6K83O0IcziN5RtqmpyEfpCiepTmgH97N1qesVjB8A7h/I4
fPBJ6k86C/IC3idVZuZAKlSByl8MRI7SKyzWO/sEngnnaL6UsoR9Q6d9jVvn3oao
p3com6ilC5b63oKFVGBt2jnMOMvBBO18va9+1Ny//rxk9XNHHwJTvev/BKKtMSdQ
f9FR4qZ2/l9jlLuLXRpfRkxqKPuQ9CPorA1oog+uHg3WV0zWGwcrPuCh+9CSNbLO
UhkVqrzhI1hmXhM4zDO0qAhCt62pd6QmMPnKDvd0D48DpSICceVXMIo5bqEKfb+/
ULwewX4nPlPvrOl32ZxT6M850gFHZYNOBGeeFovI/ahNuX390ZyTf1SSTTpVJDa0
Qq6t2/Cia8/QG7ZUyyIO30aJMTUBrGNMeKUggRcxQ7OBoZwc0cfMUXprnE50W1zP
eihml/LeoN8Qh0dcBZg8JXMtci8278GDHj/GQEjL6RH35blggFTVNmkfR8CUWCj/
DEA1+tulWWv/xq9PXYpNdQTInMVZw2h2bJ8knqPCks6d+2xZ77vA9mFq+TLZi1oT
OlToE8db3EpfeN1Spyrs6WN9AnKIDwfWbpmLpaC1jNO55jiMPgHfr8ER+R1RQbDr
Ub7bOh4fTOaQlwM0QRrlYrW+S8KkvFA0r9E8sNfRCjEuw3hb44GyaLvP6WACKVNS
TxDKY+xWhlMxX0/zN1L3p9hBbzhBbV7kDFvMhwMKZ2PQjDztSuK3AEDdmW3zVP9C
QjGilU70fawJD6LvRKc5BYOlAPGUycPZjzu19Xneyi4z9sl/1b7VgUFQ62eYyONQ
o9ZCjMY4tvinm1DvO9bBPJLkfgbOtvAIjaJzgxCkkclbdv/1af4rafjlIMjj+MTA
8Lcrc7VVsfmLpW2TMPx3QfOaBWYnuRzkDpVhqfVo0jP++yJRv7cTen1y2XvBr7hi
FywoMFBHXeoRnBVbByDvmnB8bZl5aXJ6sxQ1eKkU25/lt7SjzNpMQhmtFPQDzHv8
qByWKIy/aGmwsrKle8Ey/ViA5cly8PCNIsnFBLHeas8nn5ucViR1MLy5Uz/jHh2Q
o+NsvvUgVduSsxCTn+BKRor3LvUD+0pwtnp7NVfJJKJNgGP0juzCNPb8pySE5fR8
i21rcp6/g0jhXnsWDEpKFuLEumY0f/2pvJyk7/Y7SM2NSiKmKHDVix4oIaw3y3TK
DQOX/j9knTDmUAY6FJ1SOUh9p3MYmekxlR/rbJXfqP/2nVJkMKfJZ7SqrCOzKQwQ
4Tt3d9hNjT5/TIHi25YmcPuO/TcOqEjVjXiqHDA0FbKTIW1ctBb5VnMcpjc92GO6
4d16DkMPSiLdLnGUwkMGDWRos4ix9yXHlhwME8hlXRNZZYpRcjwJcrioMmsGD0yH
BNTzsduZjHsPmh7QmBykr3C4dEkZdYU+Lh5UpjT3yxuN7KAb/XeuIqtVDxhbVUeW
0DO3H0ydw+9pTLBkgsbdmI9aRjyB35EHp7oOtlnyzvg6hD4FDGFnkeFUhYynbe5F
w3yKmRQgQxgfVT9mxx/mX1XlXlDP3jBM0m7jz7LjeuvUtUTGpK7flxBgHyWLoyn7
j5EVZomaf9/KpACGY/ia/AZXCS+tVJ7Zsc/M8PeBduVM4sf3Y12cL6agDDZH4xxx
C0MTnDnCSFOhUnhTsnLVQ+AKOOWtXc/7sd99SVAQHPw5Uw+krfZKh6QbLFBlVMIh
2UaQMSlV7whCNJa1SVSdtikpE1tHgV4VshZSV6IK0NDqEOhswriXgPIS8SL4VSmE
wLeVcUgyZt1RYpyWwBm430dDFC8ejRTAubP3Dddki55i8DFrfTbIHMBTjVraMO9/
czHqnI+UTu5gcyXo/EOskDqaZQyLX9gWztZfdstojFr9XlcaJbW8T5RcJNiROv0u
8x/7MPt2xvcs1q+RIqCbO8HfVJ2CJkb4MAUb/wrqwfuJvEJ6rgVKbBQh4gOdB+GU
VIpGIi/kStjuOHmfjOXPB1Rr0G5scY4lEcNcxaJ78djKj0pUHLzPcHfL8tGWQIvP
FrAf/lNaYhToe5YKT6k6+AV7Aq2wsqUfbAs+JEw0VP/fuoKYt6gBoQWWNXjK/uUs
vqzoaIEc51oyQ1t0MDvNTcM/8j5aN2yA/88An/rHDSjBGq/nz1E7SYzkP3cEXUPG
Px5R7vCr8lXEDMHEipN5DzbsFIs5zsu8uI6DUXgzzHGre/IkQSDq4VUqnTin4V9z
3bFV7iFtbe3z5r/tPzaj1itTpIfTVqYPGlS+ufMcmXVB4+GpsZ9GLvyNFP0QWdfV
aqFhVCZuHhpm12AGRAG1he9p3j1jNs9CCQkKDH19Zi7CJATt2aRQxjJeoQqbghLR
RrwPfkJQ4fnvTOB6I8Q5HdpgCK9tkqvfCxkVBGRr4d73X68e9rNkDx92IN4uzI+B
y/g3w+GqsSoVWF5zoBeQoxPPl8ZJuqm0LBwmnwWw2tCHS7U4u2Y5l6GS8UUYdFkc
UyApvhYM/Ge1nsGkcKRWvxKTmSMZm5+TNUlu7474KNhugmca15CO08Aa1hW0SEav
Jov+wFoXx6t9BDWkLEoOcLf6lm8GxMxsSdGs0lqI9RCA61PUDJJ0IfMxryLPlueS
gRaHbq1+wdG3C/EKfqaNqReeHux8SJOxgLagrrGUSsSryswwWiMb1RLJ1XAA/yQN
Se0rT5p0GrPiGtkd7qqUn8R+1/UkVuZwU48zuOP0i4tGo4GCslL1AQLt5+TZNKg9
IDmzMDSnJIxoqWPzFPXcgCljzKbJInvrFf81Qa+/8/mw7L89VJ0UlW/R3i42bD5j
M/SiRe+x9Sv0fQdezcgyb+UcPbDX0HAZU1LcSE3nV0gtlp2H1HlBvx470X5Bztsb
s+MsKyiUKgeD2XcoxHhP/8Dys/041vh7Lhb30t/tPlPuy7qdJdldZwrcD6FV7BTO
O7JkwyGnBhd5CXr/5/OnNRKahzRKisO3/GKfeobC8x64LsjQ8dMMFubrZXKdj0vl
KrPUu041RN9hEOhJeFFBI7G1Kua0WzGIxSRr92FFggjWmmCk1MTn6mEEAc9XYCVh
5zdIHSasoibCdiI0dFp3KWw84KYlI7/ex/tr1NPjsVTZtxu4db4pufY8NVOrZWOn
Iuu3uWyswtiLBlgPJgxPWyWJfv4iReuZmH1B2AVC/1RsoBsStuN42+mN0LnlIomD
MsB65qA4cCHssp2QPU+hwF7R5NyWDvGouszejaF2kycAeDCbFauvEbGdafd59ABA
pPpOYFOQF8lx3ZwLgMly/j6YvgIzLp4zIOh2GTjRrHQJtnACzw5VjW6t51KAnwGJ
BkeOSK8xwO+u20nObHOSg2x1gk7zDvX6vAnPJX2EC5U+Zg2zGU1EgHur28ytpFDy
X8pd9BEQUHO0kNtNSCHsT4dEAhmwAsejayGGZ5Ds6GyOonLAEO/oHM/D3o0d4qC1
a7Tnaz8YNHbuI1jVSSYJmAOBV8mThaOY6sMixWmF6VLGDLanf7tZAptariGKbUT3
mLKqmBl4NG2AYn2M5DtZYJP8l+E0XRsy46BqbyHT88xg3kWTjw9TYXi8KBkaNKcb
VPPiNp/MC4XU2KnJQou6AqTOPuXvxlMdTnDbMWA1lE5PBatQtuM8thgMN+vgRLFA
H6xdhMVKpD7RCKt2wjeeQAqX7GnyYDpLF7uEmGPLMl6uVk5d/NSg4ZuZrkD7l3UD
WICzbJ/P7oGjvgirC86GUbmW/xbURYQUc2AkiH2S3j95FfiP4yZ7p/HX2MkAJ/dh
ZC3vCxvXpZjo45Lstjp57upsO/mXtJMVqmfwPBy/AmZ+4iJylc7Gd+XCMAV/3S9n
SnEUcSmPJ6+CYjg+j4XAF/aIvcWeGdj0Ixaa/Lp7C89/10BRwkd3B96KtqfPmz0P
2JwSJc7DEozwOEkXJa77vOy78EcNWA5C3KVWAtC2whkiExUAsmrgCpNE94x95jsG
WSkNtEAHZHkRtIjkdvhqknySgjHlzqVWY79I28lk5rmoktxAGTGHMul0oYfywbKg
0g8M7q/zkbUo2G0JyAXAo7dW+mMYqaawnsMBGyI1OXCH6c+/GduI4JZ8/TFdanWU
SjP7rh/H4rBj9R1IHJxuyc1tl98ugE3AW84p2l+LL68Zv6Y5AjpfbJR7X7tioOdG
AImOKYJsV5nsCjC3kpHPom6HfXD0ggUPsMOQ+l5405rEDwEAtnpx2aeCgr+61ZGs
R4jQ+B/DB661x4Dwc/aK+d1u3Ux/5gookMYDu6hWeziKnjLKH7v0plLbUcDp0dyj
SO/whjx0TsB0YXSzvCRXSDnNimqJcPg3xjh4N//faG+TkpXaNRhHNcP1nM0CNoVj
ntzElxnDC/ANrptfxs0+9VQxRMxNWwB9LgHTWLt6SkemA6HTPYJRG1mT4ZrzGxrg
1Y1CVySMwSB1K4mwx4sVXJ+24gq48KjqLVfC7XqnaQLHa8Iz9wfbK4XRO6o2jL2d
ncjIUQ0wp324lI52zcp1pX7fauXXR25sr6O/1qt3i9q79Zeavegh/CT1Dk5M4h+j
rVz/fPK2dQY6/thYF1j6yWDwZEBhYHY8a5oysRH1qVwvlE3Sw954Y32QDSoKS+iX
mLaW9jqLPSBZloLF9W6Og6+QzvfQ4m7yEifaFjyJKXpylT0nvJVpNqNkypITt/k1
UP1Zn+S8573TTpz3HeHAmCmBZdvfZaeuojlMSmdVP5SUyF5ekCDNyQmuSz7gxTPQ
1P578fmqf8hAQqZzIc+LXxQ9O+S5NB3Fh+whryGnVcMztMeuoyVlze4tQQjSspkf
3JsQRx5RjpJUa/UuEa3Rh8mI/+RM40L4SWNQX4VABjXNqo1PhKoGKf9uM9cksHCN
viQkZIyhMwq6sJnarTkpUBu7gvB8liVso/Uo+eprcciKj6fk2zsIFaSQe0MC2zW7
kqmGX9ORL4nbkb3cEqxV78vIpcbnZFcQR7QjATYjsSw59uLNWP7dxt4Ciag/9lGF
BB42FnvGR0ZMlCBvLNuw9B7kTkK9N0gChaKNq05HKOPlSVf3nh9LGXqHHjaDixdF
3+wMpiOL/KrgPFXlW400IeQNxXviZdtPELe0kfv3HvrwzxYhLpw3zAUZGfxjmnX7
qVcnyX6bT7GfnZYhg6jHTh5ARYKgC1Xe/fc0JKVd98bwxZDihurafJ6GJwzJiA5b
VCtTnJfopj6N+dEc0t9rZ8G97rE/vwhssBdAGddV1+KmaVXbE002VJqV7EExltKk
w2ame/1DisWXE1SdPtyXJdFOgAP7h/wbH4Dfw/3h57L0bl9toxsHX+nHJnkMAu5u
3hDaFAUJLHe5ZdWf6pqlwCnl5lzs276UcnpYhn7wDCznZjKlbTrlg9igeMmpR3Sa
TeKOgQmZkaT6W1jSZTxt4rn4Qr5b4etULy+Wc8QYdwWMfiKmVM3odMsxCKogPNGH
UmhP55F+4V/y8E/LzCYoDL3l8psCFQrR2kub+fsW3XjvB1fGfstGzI64mIWn94si
3q0Q4kChZmlX5YxXAgJFKy3Nxcg0HBLBLrOT1lSowbEdOIRccr1Km0udhvq+GLiC
TMbzPZmtWnkrt3iIW694CO4c1a3ZuZ3Qn0fIVp3mmPMyhhCfzA9nRyhDKjjGDA5j
8G9igpJMaQs8VjpLm/81zO1ebLaaBRsuRodxfERzIso8p+TYPditXM2MC4NyhxlL
xKGCABTv6WCkVMJR//gWbhi317av0z6JLIZqMSLrIR+s3TywpGQw1ZuvCtyB1F+3
K0XsH4HAryGlPWcFE/e8nwrkrae07S0bLVC1fBPDD9o6NXxJhs89tgL2POH7iF2s
3o18pyKWqHBpKPqMJ5FgIxNqeMkMAbVEmR32sQLnyV6urOQILZRsEAsVG4mKGUPj
4yWU4GVGKwxOEycJgzkBZ3eeiLBnQ4DFie3A0QnICugtzkfn8+xiZEJYD6I3VWYQ
fdIT3xcjb+2RENvVjgTxQgLE+TAzRBkddP9axsWXVy/XlCiNDPUgmr4Yfx9LChjt
hZA4KWJwaQv9nXR5LhyEwJxJmi0xCs0FaSa+SSbf2euZH9O8iv1ftjth3nSwt+mr
rmYe/OYlJ12vARvRxTmA5EGCco8ElKUq4aceH0TDS5AK3lTBqHIzmAoJrykhfo9Y
VTWek4POd1FMSXPOas0BucCVdLl6eqALfC2X2/foVLY1vfHuWFovs+Xpw52n+ijm
Tf2EqLVioe8T2bAYUkboS8EN8G1gcX9yqmWFksppqLfTGAfsV6hTWFqvLePRi4Js
VNjVMvReTvUzF+UVQd8m4+isHxRzDIImximhDvVkwcE6Kt/Pfjnw7Amw9qLjU9wA
O554z89Ai2as/oqvGGuqRwPcoAShZlrqTEhSoLZXP+R4fzKefNEfzosHZ2dSg0kk
FOswtv9N6b9Ughbp00xAifcePLkovDJmLVOt9fxtlzlYX17uP+XeFxKNKJV5gkuR
eBXk3mmXvTOfasWnz0YB2lCcLn6td39B6ZwyGAbYtMOxo2TFbc6egimErx3woR/4
bqEp2LFfVsYlQeIrso4ohDkAZy2cFGU/Nt2zbG5eC/NpBj031WmFRD+S5VXzg8Nl
+4QuD7BBpbhMrD+ZubsCSThnNfBXK0o/1+MA6elJob9lzP9TDzAKSB3Ix9OJV8j6
jgYv10jJMtH2auP9nEj4rm8zLo/GhQj9Jq7ZEKPuN5ATg+72mwS5fT3kr4qQinDR
etM6pH7cNB2ZsjSACVYJ9ZLUqCrbFQKvp/vf0WPa2lT38xpaKwpfgGV1KTgKTky3
egsWxhU7FxijHWn7Zn6Hk+6Bg/76c9mAa7xAd7uwR/ySl+mEjtlCI8CiOJ3m3UcG
XJI2PX4gvCGcJYjVSVSpS55QD6RwXDpcxgv9lt7nSrXfcSRM2dXZnvdnkU/3fRI4
2f+9Q84cFgIomWNjkZ9/VR9uQZPR39e4JGxntU38iw1EOyEEztwLz6+d79yRKRzH
ENZnfqjbOijIgL1JUz/1mJ6NIc1pOOKTacAaqy5bK47TXqVvDVej1BqHjjpgQBP2
tY8SWk9uZ7iqpGt+jvPMvJU6GNg2btqrA/HBsOOggQ/rLPek2WHitu8lcPRWf/be
QhIRI9CDReBYELg/6s/CPQ5TUUpi5rSE1OnEVDWAC9V2x6zK/f+mO17DwDw3gyh1
zz4QIXt971pkd/I6f+f2T+KL4N6HcbJLfnNR9Ebl5f0n3dl5+VrVHiZVHJLszUhC
b7mrWt9usjsqdogRdhvKzUxCxpcdko1AeiYRN2i10Lnn+ALbTckEt/JsrsB2oj8B
JUzBTlbN/e535QcPuUV/umph2X2iynSBpiawVF4GQQCfionA7SDOgOdMi5CI0hc2
i077TfonrVcfHUcj7hJgcaye4hD1P8bn/E3H3FsBFUvY91oe7zlyUUCJLZVhZSTA
mDcyjOHa40V43S8g/R2C+CygGZYLF36FDbsJa/EGgpvnsSt1llLmha5wRpQHPxv6
MVq+DImpKNPN/9kWbFJhm13JC2sRQkYPfLT5rh8Y6oZ84RVod9njGkqZOeQtm3y2
DpKWt70BeIMLWBmGJ247fu3oWs3tCHerK23v+VPEMz+PYhsDnhh0yhumh7SRwKbW
Jur4dLMW3Wn0ODKMB7QrNf/SzYNw3GB+iwipgV9ncBigph35Ef0OoBMwqUXVJlzL
GfU0yA25gc76Sb9ewUFnrOKObHK6I3rh0LFlwNOnIdMv+qU0pEY7gD/dpt9VSVRm
IUAFMBJCeeHwEaygxqqO2rQSidXvpq+2mRzKW/hL7VHvTnhMOV3snTs93HDZNX3H
/8dyDGtkEFr7gIs2nx3bDpjli9ngsltYzppwrQ+wxO/g7UFgKu47+qlng35RGvH8
KAbW5+QcgLiUDU2BhOXmy1EqNv6Wn8DNxoGedhNkSWrW0ku0bnW8iZ+zzOYbQxes
xc3rRJN3x33z3cefb4Y+XqtTVEQLJGM9VlFxfKAsp4j34wjhrYoP1f8ROF7xM7vL
EgDHXVpv71aI1DhGX/tV5VDL1zrxq3ToCGFX7yV9O8L+lTmBSsbYK5Wv7dEZ7fag
MMwJfeBnb/AoEOjxMROsWtAS3TaJvVZZERTHSTRMv9Qxb4X0gjY+l6wMHLpibrRS
D035seHlWNV9Utd9yjWPS7/+CY8+CG1hsCYKh6tl7cuwlOb5f28ixm3zr0KsH/gB
BNkXts6L75mioSMmECUXUbLhvQoT3+Qa/a9nKNCHv0bpyOm6rh+JzeN/ymhELeZD
fDbPTQmtGsOXLfB9A4zkOFFY08FFZnAizsw2hKS19+zVjsQ1qWkwkab5boyKxezf
V7HSMRceOmbTWtkN5qMzI1Z5/1MBsFLwHm0TtvcU8FDeKG9CPQhI5y3NZo9pZvBk
W2ceaY+YGqWaJT3J8U2GxOxL2AaM4pgd5rQaFv2zZ1/elwk+JYLOmgStY7KHyTgX
0wIP4oR96ih9oiaQBxbWhsnRNb6Ek/UaAx0Hk9SBEdjgkqABznzu7MwTwZp7HHLD
3sY+5cwkNgqtRglSqJ6+eVtHe+WydSbNgq3+Nv7K9HzARNXYUZpts0ySDxSSbH9Q
y7jgwEvRmPyrlf+e0GiCeGTDe1m6nDjgtj2slWFltPlcoch6cGHbJisu5tOHByPF
OpbdCbO5+xTVBnID5PkVUotqIrp5Dmq076Int6Lld1PM5w1G/znZmkuIjvc0kDRc
irFha/xVN97VH3wdXLlA2+Axt0pgqT3vvRsyN9QGz9tdnq/AgLlU/iosShwG33jU
7UKqFKdPZnRUzB503hunERKzYQTtqFhlh6ksYBxFJIMJUTZ7UaXyFaw/yrOnYrKR
X8dRtvMumCirpNI83gOFI9ofcyMyjHsh9XvHTIdRvAtv8y1IgpKWcFS/461/Y+iu
6hnS2MWvydo+J/vONC9fka2YUWGGfqhHvrCM/vkR0wdhOgXxOl07sl+rmFL4tQwB
yFUxS10qzk87xVh39BF/p6DkClNrriQyK42IkgUm/0RMJ9GL1E3+K7ylmQ8pvcC3
Bg3h7qqn0sCP4W7WiKSlFwXBs6zzRqdoNv8YhgSUeFWZRdSyBi91Ss1cTAsRdXu0
NgkQf9QwE8f/7qNQzv6kPe0uuWS0PDNhDhGUfWvU4V0BuiDzgdRp5uGLgd9hKBkj
AeBHf75+grFX5HqegKUyPp8kBij6mDQVN1uKSD5ShQgK7j0b/McVnqSG2wkEAI81
T/OyY1P1b86JFjD91HkfJxodWkFYHNlUnQc3I1oiwV2tkuYDbaUf4BveiL/qppXq
6bLp9KH3sxKg38fapPQ40AdxTva4tIZ3VOlM2BZhqZguCr3SB6dSHD0tICR83NN2
8uoaOvv1wtnQohNBPqmyXIavKYWRNmrD9wqtji2sm6fxMUMK6r9k7tkF2nDg73rN
YrPqlSDBDJQUnLJ8GY8EpVzgR7Np2Z7KH5ip4QvygW31v5J70+9ld1F7cW4JAi0S
z55RmQg1DFJt6EWswlB6mzIMVoydYTmykqB1wUINeS3epR2IrMoGsB+Ohce+aEE9
nWR438gwf3YS9yxoKHCoYFRW4e2DjMJI85uxfdyGnMg7ZvJjilJTQBN+iNbhCbYo
7zjyerhyofO3EueLP2ib0+6uayB4HFwB5m0ZaPhIFKRjYXsIc5fu+pWDbZoIF3uX
eWfQB3SNeWmT5gkrPGRyj6mkydueSwV+NQrTEMUswo21CNfkQ87m90976VijSirf
uJlSrBHyVFzI1yhwieaxU0N3CkmawklHwP/ehB7fz2RFKhD2z5b85OF9J/RWu7IW
hESeHfFyQci30TqjNiDKtUhbSWdtSD56KSGMD20ojCYnE2a9Ui8iqtnmImZ9JVZz
CQKil7nrYdGA7rXGPOh3g4bVbwfLBQImnsNC+a2/IZ7J+Ae/+bGMcBGGFBxvVXj5
BkbFmNGEVNkm9y5gWDMu7GrWJwMPyHpR5Y3CUIefYvBQUtrIcXx/zyz8WvlGBk9g
RDIc1QnlMMXJwqhRpf4iLyN+ue+LhZ6498WKwW2WX9lwYRWeB1gQcWDJua0jNGZ/
T+1yVU5S2G54SBfg9Ko8LT3PjO9HzF6iyYFOuQ2Xq7hidBDkN/prp/twspfBmNWl
rK8mV3sjZivoc3K7IlQxs5y9wtvtABMnUV9il88V2yCimYrtFSbgrddHAzIeiI9/
XKHGpzdjS7sIX+SiHdlDLhbKAiV4i7c+UCd8pPpGNWgRtdw05BE4gu0olMuusdkU
EpujBlt4GNHZYdU9TLb6Dic1gRUO3jdAPP0eFPWhwB34zFtWv12ir+spTGc/Psw0
5MxMeWyV+IjYKDJTxGuPVTAZgF7vGkyY2N1iTJvvCEou/9eRzp3MW1PNc6ig4FiP
lBcxy1GvG2WSADAhuI+oP3qxfZjo95K35i1t7zH1xwpfokGifoFLSC9PqJ3ecjs8
3AT9rzFcaC5KMQrqQi4wTV4G0k69BEv22IMS3ZdL8Zetu1GiI2bcqELvM5gzTdge
P2bopkfx1AAeovgWDkAL773nMSTtRKiYiYbplv40FDBBxeQ0MaPJgK/QzDccdG7P
l+V9vjUu2LF5dWjFRcHodjlmZpTjAUDH87sKZ1tcA7C7frIDD2bT65n9pGggkJB1
KVV3jdHwdk17ps74pATyZnqhT6oop6aIjV5FTCoUixu2LYf5x4Pdirrr5W94eIu+
bRT0Mkc9N9vf1xyCWPoLHIOCBycJgK8oE4BAyQDvPpdDyqi8bM3nh286Hd387XJR
Sr72B/z1K+2DcmeJNxl8msqNMAUHCsQJ+tQuOlaPXBwcA58QXPP9eDSoc9GaZ3ls
1AsPpzWw72yg2LOLq88ThIuWeJYoFJcKEB85QItiA3Q7+LPa9sgVUztpDsW7WMxM
xAS5mXLrc95B99hWcLCTtGu0fjAZQT4vQkrUR/uN9eYynkviwCHd41pT9gihNZed
NsQqcqzlpsp7rBTE8eurvypshQ9M/GUGLk55DpjW0X5DJVsGPva7r9xQkY+aOS9O
+3IUkSQv7o7Hjm4KdHf5h+G4bjGq2a1R0ktMPzUUvk87zCPmr98u3EFNO0GETo3d
S7oekwftd/jYMUbbtuXc8895HYExSHM/kD2AmTNJ+ONeiBqEr3P07pv5edgdaf9Q
HLmuxj8jogMWjXe4+2QteTLD+QhSp7EmBdds88qOptY9NZtSXLWhE1ZUGXvlw1sr
DMdxUiwJN5Y965MdCfBMb1AIzvR4/oU9xXXQwXrxozcKSKhrMorBeU8Fgdb8GJXA
9HDB7Z5DT1owm/VtsGilwOIW7f8ZBGPNUL9X35nCbhu93UDQl+3itfXGr+kjfsT/
9s9+Ou7zuSYp2Dgb/g0hDMFKzOnIsh7QhtysLzhaJWSeNVX7V7jdojSn2d3Y8bYG
4ob1TrXvGeqcEcMeqkIyLsA7M880EDGVhYcFrqsWnNxInaUMyY1WW5ZRJts6Sp3B
Zh+8wA5yxdF3cEvIdrurGHlbY6m55RO98kqfpS0n4Y/m8n/afHlbiiv815pKWWCo
n0Jgx5ZzOg6M8MK7TXWJcPKjATiSpfaH+EhqkoiiCNQhGJ5kOUpz//sZ+FblBABJ
+ZWc908tcQTwGgTNtYlty+zmhOFgRQBAzM2jSW/smsmIukDWd1DlzCWMeaREjbdp
KcyNxVE+GfJF2o6oIm/vBqDMpFjIyFoB9x/hJhAbReTkQMFeC6bzx6aTd1x0Q+oD
2fHNH29RFhhH7MBvPerDWP93NiKrRt0BLvaxx0Xb1O0Og8/Ar8F5e0TLN3L3xrsU
Yn6zXvlAGjqB0jTOcU7LJMyQB+ldXAbBrRhjSVg6rhgcBgFt2adzLiJfHB7O02uz
2ILf5eX/zvZrMVkXeyXVfCB/wzUJZWABfQYJNjxRLWFxbYxwssMWh1qGw69d6Sxr
TqHCGUA4SGy7EXKIBwSs4xkuvqIRlBKPE/RoOlHLP0S4yZRs8zSgYMigE7b5T2JY
etJNHI29FnplWMAME8XsQcmUvWE8cpydrpse+royfZlsNvk1oDC7s3OS+MNsaL19
I2VVpc9bYDiGthXfTKEsMvR8jD2GcXteHpe2cNQgPipGhpycNeKmZOWI+0ssetRu
cm6uDPY6EK94wgdmEd6lRM8z1GvyllPt+R+CJeg8B4MgE4HpeV3mv/gefg/WlhdE
SkS9htR74TG1GBZo5dsJish7lMr7190EY+8QR8TtP5c9WKQs4u5HzKMxmBP4n/TO
57M6K0MRVayngoAPgHfMMFOxXCn4flmvkicCOz64YjZFz/ZZ4GFCEtCDtEItzBmy
vzuiv8IEuH+sontUMQgNOmGS5ijzrXauR5I/jZfoUVUsL9TJ3lZyiZJdkrwTf+yE
T/3g4huf9x9foRKZSDlgPKer2H+AJUFb3fKj3Q+8oALcHAzrWz3Z3l24evKWw0yE
t5Oa0Y8r2zshH5lzpKbGMb+0QNQXzls/JmTvleuBu75EsDVQCMWHQAg34S/mOSZ2
n5TLHyKGgwilL/RhDbwQVVLshbqFVo9ZZ5FLov4WbBcxXCpQWwjo2w84yfQKgTen
AHQa1bkV2Prct2K4CuD2Rgfd+eXqruVXixhp+RnTxJAXPJxPIAh72Wg3nZIezhAo
+bSiKQUKNEqGVHYD5eb9/LR+YY9cQLCM+cxgCAcFjwiKD2c9/vYOKVAd22EfgWSw
Gh9IPWvwcMErd68Rt7GrdEkXaR6uZTDGMiPEr7XioF2IqDt3gQVPf62LaOvmRZiW
BosDFE/S8dKJOcnO/zK3OG+jy/0yqilNz602sEqDhYmekKc7Quc4yqRMzwdlxLEk
F4dCyAW6ZtlKiMP/u0Hgye1KvlJV2VXizj/7l5qhbo95cc/MyVVDxHKJ0Dm197XH
Tgu01+OPdqx8pfI77eOcEeMfUWaLCzX7ZL47CdTgtxNtlLUiaJ6V0KrR17U3e5s5
OVWoi5jVKgaxXFUDnY18IxWXaPW0dTakHG6kYpoKQUW35E45MgoQGTeI1lQtDkGL
b95swj49KEb5xd0KWuMypo3QzhFa39DGxOOcEMa6CSwKkwDeXHt2mcMpNQgF9jZi
d5/elWhxApi+uxVSpip6HO9WMpUVSImya2TqUrYKK281wj//7KOl7TNTCooEenJd
UF4JpxKi2Rshrh+vPNgMC2rl24hJbw20uDJvGGRDZ7rLoLndPty4dmePLFqB7yLw
8K7JbXrrbxI5D99uDkqLk1FI41CGQJZN1Hm/rwxzJaTBP6A3NwpV2YLnDogY/PYM
pxSRSgJ3cwbBE1072Tpdbnm6P73XPgLvB6Xhkfwr++V+Xku0+Md6zgH3f7YNBWja
QetqzNVtitYG4p2bk8hfct3TFyNXh7OhlGwGA/KQpTXOXQk2//OyHwjrsrUtV3Lv
LMfRRfbd0K2fwyfvxX4Oakb22BSu5bFhubsDwu56bljoJmEkHhKV604SdFgChadg
YX4aRswc5i1XYayjjKlk5tpxq6LnFzTd7L4Za/YTUm3Xt5Mt7pQCw9Bfa9Z/fnvy
EqLCN72nPpV5diwf1ESLsinarziZ1xTi4xLyMUDRGnqkYcjNveQCcjnWneQcQQNc
q0cVQOdWvQ7KB3qadNrezX5wba5plhUz5G/c7sQZu2+B0pP7n51oYnGr7rQQx0j0
TdWkK4QcqDIhzyuiJNMVwaZAcTLr+o+18bSVvkJ5bI1zq/SbK2QUBqO1U9ekQ3RF
Asp2eVnNfwR0fuxO/12Aava9C+GVUtQvCc2Nz0nbreg8CpJxE2FXtOtO4LWHv5Mc
RuCAvd7TYS3YlVimisLbf7mfdBoqUkVkl7AckBUY0GBN9u4DJPDpfAeIb4sOUfpT
X7dItPh9yaWm831Fasi9o3g40la8yAxAAzKfcFLAgwtzOxONZtYSwn1pS0AHAR5I
w6u0hiIyYiaWQFfaHOhInsVMv/4vq4yr3DUyQAaj/8/g/mmw0yuCYAbrJwYEFHkM
Y+wLa1TeffeLzsAV71mqFdIn68uEN8G1DMYg++D1rMZSiGjKmYnX1hlollLPPg84
+kIWRGL9drXOO2Q4odULPHgo+5nhwrbLNHfoZNlVSMqW0zXo08HFTbGSRhlLtAiu
VNf0/JXuhBeyOS+BVe8ByF3Gadehgq2r257hWzdvDLB1JIcoMchzE5Z4QjVqUJbF
xq53QqsMP6wBdVksB+I5Q/38KO1tSNgA8HhvA33Aw7HDjssSYQ8bVTdxZiZKoi6h
u+SvR6RrxPFCHXg/YHAqdigubx1CAZUudlHYj9i/G8xycUik8ZV9dmCR2mYN4Vea
nulk96rRExUrDlAGIIfHg65FXBtj4FDe8nQQR8W3T5UwIrqe13rwMeNAkuzVANWK
Nr3QAjKB6x8jg2+oE+xlmsu/YgjxpFQoX2ISoBRkdx1Fy4r8najiJ7TFIRm6Nbiu
yIxMmU9zqTx2P3Wid/SL9iZnUzvSM5sTJkZucwOyQpZOoBEFrcZz2kAYOqNIs6+1
kSrBhaI8H5I8DiB6Y/CUIkgb/TBonHxOyWAh05uTYQG42ZBX+kE6ueGeW+aRY3xz
W4TYEyVNAjpHkAVuOGadU2GduuR8sCSkzvAHBvNJIUhbJeu5T+vE2RObeqcQjSEO
IuH4BcaznVCdGRUVGHITGcabUnl40Sqi5r2+lr0MdcMuGltMwMo3R7Aifud2CM93
sFoWbv93IGJzuCdGzmjWXakmJvP0tSTASS6DpRx9R2jF7BdBPKbdAVEPdqO91Yve
SZMUzyLQzO+yRs+DPz5jfU7fg/NtHezKBPYv6cEeqoAFOADLVgslWZX0gWnBeb8p
YUnShyzyVWF2ZX9kK123qbS9xKCUaQ8k2EepcOIrplCB9hO5kNXHn0TlhntatKkd
o1VwpXYwH14WMKg+/RE27EBHi7xfJVw3S4f6MtDlYFMS0RxjFCnI1qo6cx7nzwRz
NdGlQzgnUnWoh4noYP3LCRp0Dd6IQpjBPmRcc7DsqdqoGl70Ko0XceuBBjrMOVt2
wgeMHH2UDyA7dNCIYBGwAYNQALg2Qcqkmdvfwbv6jn905XUHIi8c5Vrf+XA8psOS
eQ85kpzJV0fNBDmWOHGTBBEjCsSsgaZEcfrPG9Wkeu4y9/eGQ4ySrzeRYJlkxjjA
t9jefpY6nUxkRel8bBaONJE1HLdfefKKUiB/sZtFXoY6GX5KJqfxqKvoS5dKXHX8
J130gA1IPtoat3dQSm1cxjF/fG3bdWj2MCrAef4goqdrsQhrtuUPw1uDEGkT7iNJ
0GnSWEZp8VYVhKsGKLr0Ydu0HJiQYq4UorEowHXP3iCO6XGYWbeRB9TaanoNMmjo
D5PrtXnXzqei3YQ1P8WzNNzE/Gip0JOcLTtgyEf1SfING8UZb8tvFeZrP6r8oBj/
xW3yfOhoQvJTJw17jISsViB2yE30Pxg5FUCbeX+yHygmKU/Raq5K7AzTHsemNMEe
H6ZUbt6WGgBZGVe/7kCvlMct0U8KPH45hToy3exlpGVXK9/4fidovHcxzludAIbv
rY2ypQY0XxYrjAHS/G7+83I7Mu38M2DHT2kPvCaBMQT1MUz1q4a2dUWkoBHE2X3m
cs2rpoqWMOlaKZ2q27bgJ2l2Cfym95gDy1nsw9hY+ixTv4tDS2RX1yl0aJjXA+Ms
nLG8Kxrx6ulibtCJeiZzD3kKQ8HxLhNxVwUrMdT/uDXb2Nv4dx8plG8ROb7wFm9z
nLZhquyyuCVZd1uHrE6BKHclwt7JkrN31o978T+Q/z80m7qWbSXzjHtqRjIg5CKP
Axh4NpsGBfUgY/+W/BgnaOllmroPR5sQoxIYUOGz5HkdboTKb6zoUZMHaTkj5az1
SKWVsLjCCskzJl7AqV6pJfnmhToGmZ8MOaHZn23LTZ0bIQDq6wgjajVPRO3sksim
mF/7/dlpHcmSoxxv5C8y4skz0T+e6TTT71QRi22tOkbsiGog0moW0wXuat9jwfLz
q4GbrFS9WG3noMT399NsfI4Vmyrt7egIxhrDI6VVoPVvya5Jv+gxHt/yta6N9Okk
zfl8l98Oxdv0RF/+vZ4ROsWknK31DEGGeliLJEuPMeEw+TOoMz5EtNDsguZy1C0m
VAmEERjJ4rac+BYzdmhaCBGHA2ZhEnsLgLz0Oa5NQK1z6EE9Sq8FDyD8/+GmugZ7
dYrtiKmzP591gE8y/CQdO5L5WXtw3qe1uB9l6Ndj/SWlf4t4BsEUQw32W+mUGeAW
HDiYGaw4jOMuBw096NHtdo15D5HLJY4EWFh+CU7VwuqohjhgARfAB1spTI42UNnF
mmTW9zUMLrtNtf226Ke5akm00zDbDdsEAgBKdK2MpLPL1xYh7MWj/TMzkp1sdMUs
h1gP6nQoZ4Bc+nTrjIqAFfjDQFZ+2HlYMuCXHI77k2QxjBLrMq1QsUPaJdDGAEjQ
cnMA3LPQBqjJDOFld1Lhd5QcscWXPjK5vZDR9XTn4PLMMSDSSK0T2udklzyJEb+d
wu+bmvspXgXFhbdFwZDeVrWamuQbQQtdMOkhFtY1wHSFGc+N7FFydDt1y3BTBNbK
jF58Yw1BEJJnvvhrzZzOy0aZgMf8w5SJJAejdDErXuzAU+umhx94OfRcIq+xQaDv
hTdoQAqNShcCDLeK19vWQj5tO4uea+tfl+lMtJD9zDqsXqMAxa9cUat+olYVndKi
SpGc+W65rSJpJIRVns0ithC0yTwzr91hvod/Hhde5GhgMt+HZED2MFlVo/wETV8u
gSifUZZAIry3con+noo390mEnpWUxq/CRC0NUler/Nm1gmqkxHnZauKqq9TNRl82
Rcemq2463zXfBMrw3G9HaGDj7K0+MPVckoFZ2aQsFRu1KD1+yhGKEXvmDSl/WQVR
SJAE4BQ2Ec6Wrk4Vl23nVKwq9msOcW3oTMFTQruuOknZR3GRZ0rdQiFwaHpVhaRX
p8WbiujrJ5wUKWgLhZodTPvxzWs38CnUQAGMFURw+Bp6goZ57nuw59osfcDtOe50
NB2qV9CU8j4sc9rO6RV2D0k/xCHChfz4GR82Zqjo4mMi854/6gD/JJ+E8lHs4UCr
HBEAKBPguuE2cu8HuwQSIi8ABHvCCUvrbWWHX/IVzja3SX5E+lsX2waG29UauOQn
bmQdrFPDjlKp5w7oZKhmpalpPW3tnEkciFuExT1t0eMXuQEn731YMaiiosfVzbSQ
+oM/kGylVXsnVM55KPh7ahq4Q7oRfoTTYSFFbV1KH5U54GVttX9fjapDU5bdq5LV
ppqiqrEsv+IX+UvXCE3b0XekjqncRdOIUdEyFD71I353Bgg12fZKXLvChLwaygaE
j6Igf1T5pprF/PM69wJX4CuCI9fsPCWR52QDXPc0xq0uGXJO5sn8yBpDQhQQt8zh
PrHqLg27VyOlPW7wQagwgxf2VAylVKrWHJ5KHFPvUMIpWRx1D28baXCN8gicJZyL
MFQ8Ue1wpMVC2LHmiNFVguj0m8zGwkWSdroeAXFVc2ZCEYIfpkUwfmfh2w5TJC5n
J1X2HWkNydqu01/MGSVcwa1vAbre/VY5nC9oq2WvgprbLUJBG0w5XCZmeTwsnG9f
u4E54IClVEAJxmFnCTth1roz5fgal5Du/loyfu2+ZW36GRXYvteNafYdmBAReqhy
f+Yup8KbjhlgwvUQGqBzZNqXec4p201RFWCAmjwgXY49jTY0gN0dQxRiRraTJ+GA
H5s/r3YKAbD1ChlaYKu1y9anoY2BOKKJKFQtyhGdbaAhVZm4aQqbaGwIwdy140OI
6+yjkGr8vhLt+937qFXVrhp2Q7qtgVaaT25YQoRq48frPgHeKeoM+fwVf9aQU7F5
1Q0VRIXJE9oF5kGpMI0pwF/Fr8sGIsqFZ+BfvAXL2pqbSFz4mWxdApTBjGAwTLqP
/wh8lgA9qmfUwMnwfo2pIqdhP+9Phxhv5dJX0w2t4w5pjcj5kYwFP+tP5QWLnIEh
0SQj384bq+JW11Vczpjp9mNIwFmsUs4P/30H6w2CRIgJ9Yb/fxn9Ia0wEXRtmBQ+
eJNrqcomMs/dNR0euITDDaaNY3ypIKXLaZ4jTJWf5lxUofTD+fgbjHAJkC0hXn23
MMUGdYSAR25TczEu4/5nt4vK4rcfPlgRq/1L5ra3ZytWzcL+xJvpGGaY5zIkkMez
LZXQ7ZV1M7Itr5y0wZfseis6tosCqa9vG9KOxpltpWG9ZoBt/5swIjPHOwG8Y1Ux
6qTYyunOjkL8MBxmrjWTw9AybmWxw3r1EsIdaOSDdjqCXM7wLK9PUoW48rDOR+VX
H85Sa+RQra/jKTw+cmwaB92KVpqEIZcSW3WLpvb2XO5atL/4hS5tFhY1qB243Dp0
YwP5IrCyIJ5ukWqMspOKvFnqvU+c23sw+ErhPQ861q/HGyg73P2sH6zb40WmbIsQ
b6QrOgQra+13umW3uuDUCQpDZkXH7ADnoy3yrlSD+AOqmOqDB3U0a73uOE9MMkgO
2R+SS8tDkJeA0zQpparjBMyYkrQ8Rs4R1bSgn4BB4Nsk+FLPhZCap8cb7mGwSiPW
HgrVBM1TTD83tJSy+sA6EXWcdnTSE/l03HvGjGgRP8464N6M6FJzI0A85bSN/tBq
z6VEwdOduaa97VEvNTGazj46WBFwYaKoWCQ71WVXG7Fu5QTWFSG8vQBmDV8XfkQH
k0kTfXuZjX9y1bw0gFiVPf5Zg/TN17jqFalD3Eket6mHBn2gWGaVdMTb5XTjLSMf
Z8TOE8jzxqJnw9M62ysWSOwhYKwA1/nlzPSxWRzzM7OqnBk1klyqJX9NGFeGporQ
+JxF9WGKFN6q8JO06NBjuNfJJphl5suJ2JAvzGsEmcKE6S/AZehWr0BgYnhomHZE
XAGWbjmNZrcHAEi/G8J2f2uASZS7H/1v+M0Qzp65L8Yb/mI1YP6NfEHxu5iUxKck
9DKN90kJNS6pz1Bfd3tuWz4d7Rwu9HRHJeDZCh1oYuUjHPslkO7sJvdNw3V62u/o
DhV+10CmDZQOMPfsXxdKPT6RX13/loqq3NSgBuHsCOOD9updeVOFMcs5Tny24QZl
HkpX5ZeTkh2QaPLP4uUbvCSgGn4APdPlHoFVIMXTsfYvcfmhCp/WBK5iL5CS7hjd
KNd8dex1lc6Va+D1zsWxk9OWz/eoAAQoa85HGg+IqbxvheHyz1S5vaMu2X4We0fJ
aq2Y9g+aOQLpyu/edhKDWT8lPpuYfYgu8Vap2P8WPYhOkcZh7V695tSIJjtphCwg
d3OPJktz1mqNBIjXCIYrjxvAejtT1TOsgKi7/jY31UXi+iItXZdADxjFN8D/nJ91
k5skM71LwPR5ouIVkN9Vi0ZjsGnVWUVs6d6u70sREZOMk+KEy20J7M/Ew1zVTYsU
nKTQW1hcUPXjil4oNV/HfARKjl2B3Qceb2+zvwKIBlq4pujCaWe/bKgJaKlrLkGx
00tLdx/mFUTWviG9L3rEGHZTUpINwgyd89/AsULrpGYgfrpagLqpma7/JD3zhTQ0
pHEjqV/l6HQNgzl/q/Yk+Awu/1KvlL+aCjYijzyK9MCj8chaFaGUTdMKsy1xDbhi
U9fmf4Nf2yDB/sF1IeK/xxH+5RYIah1yblXJNMEtRRjsvTAvpgCbjCtZL2jsZ/P6
wWwY1tw0NKvLzcrxsNYxTXAs5n3LUZJPOfdHJNZOXaFgCReHWBMrcORlhxSiOZjt
GcOieWbaNEUof2gzLvD/BPo23tDI37WJeDtLHPEW8l/VcwfMaUu/09glMgMcs7q7
2b2DGI18fnA+pLaqq3JBOF47zmi0kLZ9CxWuLOfM8i8CiOslCpRX+veQPgHyUASx
G1tqpF0Ck5gqISQ4SRS1h50xbNv9SQgI6Z20iIOEnvpPkmTlWqaSTahvZi2CzqF1
VsTV5ZzFKFSOqeYzFIhIbGUs/hh1R4u8xQ+2fmVqmceuv+VQZ0s0w6VqUM6bIWtQ
D7oboiEqf+IqWeXwpmrqYtZsA27i1zhjfK05yIVaXk1u/hZxw/AmT9iHtDhQX4Qf
iLgJdAdlKYMEFs52Lz2+IaL8IdT/ijzO7TKD0yqK7BSiAobG0klpvdmXhfRBcAn2
jBX7TT/xQ0Hgl36+LEYtbzhp+etzt9+edaRu8azftiU1/yhYna6CNXyJ0FN+E6dj
JZXpVIKm4Ja+L/b9VyBInVOVCvlXv0KuMM6dIIQDhfQVgE+h/lrPzxKOkxHyQHg7
Mo681JP5QH+r0GSBCvLmPoatGUvge4AvSHOMeLGzhoJ4IAM9Nc15HUh4FVkuh+vQ
nvf+HlwVCbDy3xW82yKiV50hILPELlrBY2GY6v+UCBnCOwVzC4wPCOYLqbz2bkDo
GW7mTVDhSeV2xr5CVsDgs7aSnZrzWKy1tshRW/+oiEJy9w3jqF4YUs+3v5/GOxzD
FwoCq6QrE+fDlpaPdbzWlR6gqXFTiksg0S9x7aYfc7Q4gFlFKOykKuAGDIxyqiCo
6o12jBPuAN/t7TuryRLX6ExwvjvM2rOTryBO+ht+q5XRwjGhnQmEFzDw5Rn62xjt
NkDA/HjVH5rovGXA8N9xoBYzRPNxgkgYnKjTrE4cwWuV1UFg8RSnENWKMT/qZajU
7Iw9TzffZhi+ZOLhNFw8WPegu251LrL7YGhGfCIJKqwWIbGKbURBaOO+mOpgFymr
gONXOAzzO7dSSXg5Ef5WXOo8BME09BcUmgtKODv/9btvO/m1BLtPsBYqkN7x86t/
IaV7Ng1F5Sv3g6+eJvmNN0tGsOCuKv/gCC3ARrdVI7HGgrzgune5ufR+FwJnfPwo
7penmFkmaNvWGSVUw3/BQUsLRUgSEP2hqzQVp6tsHqT7eh0ilyJ3y7mDQP7cfKOw
/ABRR00mmrknFfZLPUoaO0qkUvGd+cZkq9x+M4DDEhhc2K5yhO+WArWyP8yLeb4R
8HKo4xFqKVlz7pyXKYqRRR4KP3f/zFSCCpooZrxqB21/25M8RI1dIVoxoElA5VU4
QMxyqyu8JtaeRL3JC+7ztA4BkWPcsv36tK0UsCc0pVhZ/8n7zKGYO9j9bUK9ovoW
2Ra5+cM7dAvS51W6B3N80spfruTtu/5UXg7Gsjpj8v/PbouCYJ2DtTDRp18orA6y
waJJiEx04uZ2J1oj47z+I7v9lq9VIkvOmfbpX/YJpUtG4yBW6BNj9nxCqOXJ2YtV
8Za0Mqz9dQTviL8UQXHEzzn4g/n3LYmV2ONraJ3ljlX2SokSTKEALRo0tLE25yft
1kFL1T6+2RLD+dpPK1brESigt2cz5xZx7nl5T9tsrfL29rQTII5d2jGtkOMgE3Os
vfuEV4mOY5oDEMcBWQnckF2ByNnWi9pTR6PBSNQP3YGOJz5e8EedEWJ3hw6ROZaJ
vbeERfMspV3ZpWIViOrP+5tlx9/0I1EtWrBaNpVKs2XwAZfNGa4CJl1JHuGrllKZ
7+HuKDTXeii/j5WsAJkcvJN9UMsONI3m1O4qRN8bkin32VGui38exhK0CPoNYWxj
enR2s7xm+fmCzieKYmGoD1SWrELFpR+oqsijtFojk1GW3jVnazPVggKg6aBUJn4T
V8f2yx8LF9jg7hHr0kl8xFdxedeTd4JqevvuHUQDZe8gwRNWiOhBMjKuqovr5fbg
XnCueOkyZXoIZt8nGDc0G9/m9DVY+V0Fr817QaEyci6ZIvE8MtY/Po6J0UIbJi9v
/dVtvoY6YBzwgrSomChT/5rKP/9OnFPn0FIh6bqhUp/Eyjgt9jsHQutYMEFBCMEj
qVnlrDUkOgrQJfe+1Z0irtNRptj19E9570huIB3JCzQJKdVtCK+niOMu9Mk4+X0w
BH/dfMF9DioaGd9CwKrldKObxIv1ifuh/WUHhsFchmLWK2v4s61+HcgUKfR5vmAq
ngKJrctXe5KZ7cPLZzYI1f/jysjgS26QBk7dRMkiMwUDIylT7/cwGH3oLThgN+6U
Zes29TpwJCNUyTjf8pQrEYBImpRH5+TTAzDdkw4p62CJZuqg3C7qlNXAadgXonES
F6ijmwbwfjb/8HpWQ7kg2Me4H9xY5gfZC/PJNrIhmEIAdESRInsZMiz2PHBhCvjq
eg/H07ozNkxUnWfD6xwQqonoIZLbHq1qzT/ePnmJGOh7YUu7JfkWKUkpOibUr3Uy
HLCRsl4WiFaN42mg0BalRJe/XvnXwpYbGyhGsWl3TPbItAmPOC3XpYbZyvIEF5IA
I7g79XHfAKDcePJ0FEI0iRdfezuowp0eAO1xXvKK6BP26jASSMquUF6DaPaVE+SE
u59XQmmVsMt8ekwaTLD/iCZrpp6p9kOXlNzlWwA7FX0qLXMZe7X5Nq/kmJEPe+Fq
wlG3vVWbXsmkafcAOoptsEsTlNk4inyTLfK1joVYRdKyaEG94t+wP35qtPjZFQzL
3vOUhzR4ok09FKqrHgH/B49aB8PToHw/FSr7hY50wF/y+y8A6g09kyOLdaaub7Xn
MtohxVQHAPAKG6pepz3VySuQcynJFv9Jdw5dDlSqSQ21JCSZFRuAaVGlP3oPMsmS
TK9+nXqrAKjmyj6cCIFmAFFbQyunFdjZc1ZxQvXXYL6vzKGOu7sEwyGDM8UyPxSK
D/OolCYA3YTi/R1MAGAjD1mSjglXWfzf+7d4f4I6RXnDu3075wIyDhzZ2Cptqlos
KdaVBKvbwHO6r17pmONCXk+cLG61RHrFuLuPetjNlYtskqNhFUlXUHOIU+U+LdkO
9YwcGGpAXGZJ+UX952FxtkWGcUiFAmgm41DET7vK6Rp8c8wqjUyve+lNGV2/aSIw
FwL8LSACjbLGDNk6BhMwK7gEyhbToD1VgX5dNOFzB6zdE6Z+C6GISP0wpEdSkI1O
+8x/jrWTmEwcWChhOolVI1FFEpLP/19VA3tQSlUW1JPFBkllnQnd27l+1qPT7bBL
t2nPxkLpX1rJJl3uGTtrPa1fEQvZBk3IfDpqVBzjIv0mUnmhZhLFsqnZUNV00LXn
wHTFsktaFm3tak6B13uOgedQZ9iBGCWqyeEV62hLKeidFVrDlFs+rvUYXQpRso+W
AM/KKtrUPrm6MQFZcBDYo3gDGQObAX+vaPZqNcc+zeMII29nODHUcy4ljQ5VNgOW
8kTp0lyaOFttOZgVCc0dqE0A9FAPFRe9ceInX6RnnDPh2gauXAZhtTz202HlDc0+
kR6NoFf2Xht9huXsi6DetkoSxooQoYE34Rrd8AuRDAkvXiEwBC5WIzfJuqV+ZJ2g
o1BWc8alMdAOsHezzaykE4PeLIGqsa94K2qL/xAf09+OeFvcNvMPVfS8MV4Po4iv
NhPGwGn2qY2lLe6FqutIK7+g1LP3lnnZMt/QcBL8BYCsM3hf10p2d6cqqYMVAkoB
/ldmIL/4oYoHWJ+WtdajT4ApdVOZUIHWonSxff8piLAUSTxRgLstCu6BOx7K6iHe
ttvbD1IE4VA0oFQVDlCHuaII1eYIcdf3MqsQxQWGPFPdgnsBCDRup61hWqfMp/pi
6YGY4hSyHV0qQate+VGzU2xbUHoieKxvNj0Rp9uBO0CL99G7H3nFxskdl/yBRuJC
muH9PArrPr5XKajuQlzs9B/Cgs6O8MY9vKNpKakRy4CO70FfyDUHg804YLjP0gdJ
r/tKMQJfP2AzYvMLmn8R3vCHWnYACEEwmKEKAKKE93h/b2Ps6Q/lyuSA6ntgk01K
0FrkL7l8x1VleweB9A344Uhs3S0opfcs2DQmzUE6tQbaObBN4tF+rEow66XDIz8y
gYbPDITYQMaGKItg6BAD6OonLvNL7dAs7JyYpxJCvBh9LRiE0RNXF2vFW6UGmGe1
UZBISNcnj9zfjvTQ60Dlcvhq+HaTlb5fEjAhchW6+Fjx6R0k6melyJZowk3VnBBG
rRrjXZRk/ftsmTfubqVAjN6JNfEiNDwtzqERChyiOYPSQ9LotKp3QChwaIcgNgV9
hnoDl0Tmjjs3qy2sGiPPJVfFhvuCjbbY9vpJeFYSXgsMA376tZxbpfgXyQQbrwRM
31RNU/i4Z2mgNdIW41s6zijeY3T0/FtMt+O21kv8oT2BWkv+Y631wagIKOc8Xn/j
al7NzD+vLcMMUThUSxYJEk+nj9w7nNStTPnBnmHXE62yE/U03vo2ZJQipXF8biLq
e/z89rczco9gVauPtVBK9qvceqsCIXmaqwB4kGgJ09Fgm2rDPNZE8l7PVVkqneEo
Y/bHsB5BuUr5nqAqSS+YZLF9FfBAK7SIdkHUbnTc3UXZXhi1MgjAb58sLi/BFqiZ
7eNuzSW+wPVXayp0Bvosy+/xwXksKpqxEV9h/0fwlvSVT3LVjROppel2lpJDqRI2
f/6Pt+5D8XMpUNLtZy5I/IXhelkPVh40BRhxRw0661dt8rBATcrT2bMjY9eJwMK3
YiKJlQ6ZBdoK/CF/KUcuRHaW3R0BxYnsDvFa+KB3tD276t8M9c3GxcysAjJZI4oA
rjB/QzP5kvEax42QNpCtJeRkpsQTOqaZ1v6c81lxTZY9yyGlofse7soiUGM7oxB4
sInFuD60n+tNTKQSXciBeEvc9Fr0VXRZIby/O4+iyc87e8zpu/xvzsV0QHG3kePh
oOpuaUMBZIvHvXqcsx4yozsGxbItVO3ScomtFvyAYnKJAukHI0gR8Hx01I3zpXJf
mqAFxLolC8i53Tvj4VtvRAvhILwCfzpRZkfOTTM/SsCT0NBZimep0ssAbMWRxE7i
CQtSV9M2Rg1PHw4r9dJBXXS+H8r9lsuN7n4I48j7Goe3aMx2Wht4SZxjBjT01TOd
E4za1sciT+jWhypSLqpufTaJHW5QEzTfuEI8fUW+yqXUv4tHb7PyIIAXt9ukC/yV
VI/Im1nYUr47o0EUwOlWqcuNuLJPpiiZ10G4bVymVA4TGPBLWuICDjeHHqZZVGOv
8ngH8oCxQ2lJr6xgqh0njbG404E0+m1IEzbjODTmjy69O0iHm3xzGFJr8NDPsDJo
zaWkDfVmKYrIEXEqndC53VroLTQpEPrwlptLCZD9EuIzJMuIwc5S8Ao/YjvbEMhL
6QphQJzgMhqSvdtltbXtlTxSK4Hkc2IheJEyZWJKP5l8pIxzEqHh3ZNl0ofo8UUt
0kIw02wwzCT8tVxOwNbZe4VHDGiBfOUuEHzTmOJfN3bkAMIugF58US/1AgCTl1OE
tiTKTw+tAkinmrbuG+KsZU+QnYyH9kmvdODloV2EfLhdaDdEVnABAgXzt6pAoKBd
oOkO39ZDysJ/cveHd2QSZmlTcGjyTVqZQ4RyVG89KbpFq5Nq3F0mXGZYeRTnI8ol
AvgH3du9azvn/evH+BVbqUlTedKRiCg1FqKqMLI73MwbhFkjK9E4z5yMI+qyFOP9
upUhbeZn+um+2j/AVbQJ7HpR3rkoik5C+i83ThjZAXT2a0xfndGCMHocFAcc1aM7
MfBXxa3OTfDIuD5J2dr6D0fDZ0R18xmFAS8xnwisx6iTWxhx1/joIVaJhLsny2G3
QtD778Y5NRiBeCwlexMqC0gRKAvjQvwL5ZEAcpQjxWTqufGHuoPtJx4P+vPhbg3M
Jnv88x2QyfAwnzBxpDelgEINcuDPWULIbeqWe6yw8YyCpP4f0d+lWQ/IhcpMdc8j
KjjUlUKe1a1thsUy2ep6Jcc6Gd9EEF1Py442w91H+XspXS873avcMblzrCXjxzbK
ioC7Bj5l5vfb0l6XxRXM1F8BYpsmB/NTQedPPCoAU/4oKguZpGrpp2TRdmhjepUe
IgHgjWEygK6bWFEf0Iox0TqufweHmS5JCGEzTZZoHP1gbMrt7FIywJ8Iy+pfV0J/
jjvBEosQFF6qMOzGKWPICv7yRBvVD58PpJfQ4YeCOTeAuY0AqXnvUNTH2jBrp/tf
PvvN4nXZ2hi8lDsoYZvYdquaT+EswttvgKNCjMfMRFYVjqZWBtZeL0ivcYF2ATLL
FQPttuWv8zOQQUE5kRAoH4dWbT47YxBgFVtJpPWBDvWyC1LBTRUlcUVrCntFIWLD
aI6UEG8toTOR0X9nx6jyDLHkv09S0yEwB0NlZ6tcUg+Qw62/lSumIRJ9awIdEFM6
TThAd2Y/dI4jDT4i1KYXtBDh6OG+n/5qjvVDErN9YYVN4WYiFAgtqyfvPjtpbEGU
fpPLluAe/xklwal4GLZ6Rao8kfcSJFZwEw3mQ15gCyofhUEAAijipKqK+9ZTYmAa
dcyWY+H/5l7NLHy9wsE7Iqbj/ODw92TPlJC96nOwA4tL8EwfarXjHy/l64tOyycC
N41Vy/1Dzc3frJKVw6v0V+pL/mt1qzkekCeW8tBJze4150QCebrqQk467g/axHnC
LIz2LRkBgDMF+MRnN/RIzKH4aOtKnUVMJxbraJd5ALBF2AQpXc3SP+hTmm9Y3qmN
5OsZ5ZfkOyB5hkSZnX9NUBw2Wz3npIMEP6XzfIFwWgrQhSrL2IeJBZ3Qjk/8ZRya
5oBxsbfEak92BDssWAcYVc/DrPwMdRb+QUDqgs7/qBpdgxyvPhNC9mjzuTYznvqA
YpQ40ZeUpDiDJEZCeB31v1wgXW82NTlv99MNuqAt8uMHbiv12gjej+l5OWKMrcst
/+Iturtu66YYqHiCDm+aZi+SYxUSgzXaeAYWeninJN9Z6DmSsvacCrwS691z5JtQ
4Hestr0O9FEnqRoiMzuPju91q+ztEEnvjidKMDvkg4g60jHz++zZ8nt9fHH8qWOl
nfdszTmeC9+qZouR4PxNUviMY6MWGLNxk89Kl5JVYsDObgac5OLyOZ4HWgfyOVXT
SjRV3gYHflIUbLJgJyVGRFlm6X6CvsjQAk4cN4sFNQl3THaOVBi7Mr72vihdOMIQ
4rx8g9DTA5ny2BYWXkXAzHE54ns8NjiwRRLjewgToWKzljvqQxCb9/ZT678/Kx4+
JFRT9zpdgSzH0nXN1hvEsNCkK/oKCS7rD2BLY1jwJGaT1mSa9f/ct/Zuu3+jR8XO
agO0kORENIKYsc5zLQAE/vSxtrfU8wuku32z5hIjAKnUHUVUK3dsalZctwBYCXAA
zkF98VNSw9DGJKroJAtW1aR6cLfXJ7GBdvxRgDWAvWICz+iTsisJsQzoOGkmMbwa
87Del8ho1HQkouON/dtM2Sbnx2j4M4Me9SEpNcAnA+lxykiFLyCT5vqfUbOBqSNF
Yo85T0gw7dTHDCkWxStaAuoOGwCEyyPVqVIWJfBaaD3mN+D6Phg++wK/gctuQlBh
R0uqejuUUuiKhDQyjQsMSnYxmf8zraPfgOTIJmJVYQ+DF2+opM4UUJ7oDrVwkeKz
f5Qc+oQaDwNZG1LzRISnnsC9XOC2X40cE8tfxf6JUCt6ZZ+NOQJjihGyeZxSSocb
CU2eEwMkkr5XrvAEmnUJnXyQMOtmzvlad6Nb9/QdC+vy9UCnkurnSQDMgqlKAVgC
G/rpA96JQQdb0Vx/MSURHEKDosHUyNaIzAn7dHDRsQn7AmcI400LbdgJW/5pRMup
gZG0GxVM4GcsJwNwySfgZECmivhd+F7zbG57kENFRwWFfBpC0JLr2CfQQCIqsnGm
ZVSSaPiUCtdyJyIQinU/TtO7Lda+qiuJqLRzKeVsUurLhJVmHCtOEmIx1CZN9Qls
/pwmIzFal1gYoRkL1xGyKlzQ9rtqlkAjMGH7oJiN5c9hB8JKZEPGOOxfx/KVFLJ+
8I8Ua6GYonJkROuMsz/88sWqFadSeFqCMp2vcz/tTvUwB6ku3UiQ1k5d9ddi71wN
xBDsD/ZAyIyvdW2afvapAOONWqCGw7Do/BDCJLUjYUyvuK9wZx01E5GmMxrlveVt
rX7xnNbXwIiaVQyYIlnuSZ51Cp6EJ5qd68gHLHHb7EXbWuL0clho3ukhjxonahug
9n0bUGcpSKaWJzk7PblCt3XAlnX+ORs3uwB0buuATt3MtH+SpjQVz05go4WcXROx
Ua4IN9MIxD7h10YPHxEKPd8WOEVTwhrVTgcakV0XXiZ9ICchxaE6Wj7/xDalbkE9
PFRaXduFpUqrBgOhHUGW8jk24h4y1F726foqOKR+f4eq9zf3BFv0HRWAAizrxnC8
DamruSFFtabZFtsA8RqAicwbvhxwwxAXSioV5UeHD+HlTr95waRd5F58JohYMloX
K3ioTBlprN7Jy+N6XZqLhZ6NstVyEPiP+2Oa2yv6Ur1edYTaYX+U9L5PnclIitqp
I7LbI9PhX/fET52hJoBZPEKuehlm4a3LW1czEMwjQm/3lmfMEjXPqECIML5a7PPQ
WJ1OGLuVt3PTj2qEuRkCu/c++PoTAkmoPk0sL6SthyMo9a/x+Fb5b/Qui1N0uXsV
LQJnMUO8qBV1BmGR8rP9ybBsV9O2mOT+68XuOA9KYvWSMiKIN+x/e6k1SxtDMIet
55fn4hw/zg61nO8uxuT3nGKGUVeiO/g9gYzdt0h+l3d9A09fKX/iABSThzSGICNp
tT6FtkpZDUXVuSWY3l5t6bqESJk7WzLKMra3QzHY4FjmIsrWW0dPJxCB/PJU2uB5
YPZCN8VvFqGiz1Rvxy4WoqB/h+z0uoK4aic42jDlQRMs2hk/Cv4C+d+bYXnsFPCn
vFycbXHVXB3RKWSoJMjBOqe2oEx8/x/V0Bzo13Wpqu6UQTMSaHRnKALk42c+Kquz
6GmAgc1IWSVV5KYvfBPyXIgwkSmisjaglmy5h/N0UjuI3mGmfjWEnMA+vRliBbZF
SbNokr9kpwBylHPGCh5GhAkaG/ZcCdDPJWAsd4KDYbvMEspb6Cg25V/5EJ66dU0U
zp4l+zB0KWmne4bmZpKn78tZ49OeWM5yE0QIv9wYmYM8LE/BExuPB8cR78qi2l+z
oWYaRGuUj/AqIBGytTQUBRbUb10pUCnoQChUhyO5Dx+Sc77eZvrlRSi1R4TbV6gp
qnaQUs+H6OiTwUXOzBDN8+A3FgsUuN5yh7GNSj+ukQI5dgVQWKfXn6rDvnTFMDT1
8vr8LeR2CgqAnh2sJzR7A2+WouJj8DOLJled+JAKZ8buF3tR2OpSBd0VmXpSVDgb
`protect END_PROTECTED
