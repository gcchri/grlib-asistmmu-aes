`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQ3Cj8cNEduKegoJTEQZdcdZGg88Y6jvdReW2UxuDoD1UAYwulbRX0hru5K/cigP
xofyLxizkpTX4P/NY+kLXvnq4kKyTcIFRSvGz5UW9hUJ8hchR2chfexl/uxMLPGq
HNDXzBKS+9GsDlR5pukRDaF95ZSPZlYgb3Yf7J8lYMRHJa0Wcp5dLBhOhlP24jWo
u2OCvY6vMk3aBI/LcxNU5ccZIFz3dmg/RqvZZEkKF7c2en8nZfuGOBs41ttuqzDj
sqnMHYo306gTXXBiFKc5l9Cmgydl4z0oDNNX8kdQlK6Y3Ls+QskSn8JpzlJmVV/V
c1auGuULp9AF8DtT73imqzUR+R3Syr2Yf3QKfoKm6g9VcXQ6J1yfcTPD8+u7QTce
cc2ZKJxk3ds++iaLOIQvh+dVXeHB+XAW7Em7MXe9/ynMIDwKuo24BssWXhq4yhax
Okh/opwQelNgVr51295BUORoDIiI4Nf93949mJmeGusNWw3ISXaQYGx6IkCY7L+i
oEmWfG8iYC+gyAznwlJOQkzef/I4wvPvQQGlQBJXo9QOwcXuRTKUwdk/sEnY/g0i
LmU9nyiu7l2ZU6zQZ7r196BMBdN9s30DJ5NGMuvgiVGBB9xAQCCyc0HirUMN9eoQ
7UMqfUB5Adef3hEYWQeoWgtmrfYheKpIDl8Gkxp0+/jpfvFHs9BrZSlnzmqwi412
`protect END_PROTECTED
