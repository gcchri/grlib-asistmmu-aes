`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iyAkJJOnhSoxt1M/U7SPj4qJ8+fDqY0DWaV2NMjsa+efErnGzwMphrpTJNUT2WYP
5utpdzAZZVTtt66MZkQzJsOpFTawyxeFrfb7UibXaeHoWNPZDoNLFzxN9WrjsBwm
UaoC/U2WXTO4+nHDrQzLnV/9A2ITIwDTlcmXyrCEySEhyktUEC34zRwdgru6p7rr
1wyXjBLWuxxpLEJQkq1TJSqRrGfMWddNHj8RX8fiU2gyEnDujU9SBZyUWD8RsQdC
3qhAaiQMdFNv+gpSPi1j5a8uRPgdr6rjAmo2EhmWg92+oRSovs2yFvnTGB1m45Xg
DQlVEDGr5fPcbDbzOkKDxP+xigc0/6nn5zpqzfu8e0eQ5GbpJfftss1ETVlerLQj
4+snQAucwVwnsp+36RHR4XcOUBvBn8JkNwZJx00xKJ01fClX3jX4TZmO3pOl2a/m
M9mJnikUEg+KFWrfB2yFYQBQIfqBfp4OqIsLbj067IBFOaTXhOZLBllzCccKXumu
+nIGZwcV9HuQntkSHkCisxzDFkb9Vme1hPHuTfidnDWDnPDp2tQRaoCNYNLuetGQ
wWXfgJjTecQY0DxrUb+WUxNYHJvnwbhEbZ2MUFqC4CQhXNyT1b+OaXqSNO3q0tHt
t7aETIKXwRQmJBjImbsxUdFLVV6N/rS4KP3qlSpO3GglSr+9+oBqVobV3mLdrR8c
TuNiCyP+u0ulQO6y8KwPng==
`protect END_PROTECTED
