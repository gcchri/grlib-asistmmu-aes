`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZM/GtlxyWTS72H6hGWEDviOs4LVV1vvm1JJZqwD0Hf0w6AofY2jH6q+9SS9c5R8
6w01NmXS8izIgPkgT5im+soVmYT5apf+gUOJCO5p3WFk/aQsjIjl6GCaYx/oiLHX
POXb68HuNv7WEjlczP2zsIHxhVRZuHFow8/6mj6tjQd6+2wwknAqN2/ESrKuFn+3
ZxQD4mz2mjueofKtPXh83cFks4/Z2w7j0Jg1uGw45w8JKePk+6GrIg3FUebsgOw1
Pik4yT/+xArJ97Jzsg6aMQC20C5/AQuNESVbICUt7tA7rbg7GEtOJOpiCaj2rszd
N8DD2v1MEsODVRbU/ttg7L9vmYQL4utDlMMg8J2SqM1gH91JSZ0TQ0SdN5Uu4reW
`protect END_PROTECTED
