`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+AWJoDDM7JvTBGZ1LsRSfjZN0u2XxlbsGfYU049YMJEoP6oOgtbGOUyCNFptBlx
ZWV5/ni3ltwYnfBqwNZ4UyWw8Pg91Ed1TqkAaqQIcoNqDlBgwOKJl+Tdsgoc1G3k
iqP9tbTM/OQQ3gKDcI66sUcGktlvfSfPfayX1wgbFGW9/rYh4pwcQpX3K3acd7uu
BzZbqR56RFSSRtm8awUww4/KlXdwtaNprfe6eGWtQqi7oTweL0H8izCZD6OcCM5n
r+vRNl33c+u/AyCpARFCK38vfS1cQYPh/su/dHg3bVx6zkjm5Pg0VeLvL30BT5mE
HAOY5EiUPPajls/82Zam4HeKJaYOJ263E25EDHhP7gmB8WBJ5iTt981YSbOOve00
kDHfrbvxiiq+fd9HILBForZ4bwEmpeIe13MSzjZXLjJnorwn0CKscZRLdFOBQMQw
6HIHXjB+VEeYCTn2uEGo+5+cAzT7a/oWCO2Zd+VjujC4ZC9gfxSuxRX7QXC6LGYr
`protect END_PROTECTED
