`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AMtW1MB0DQO3ljtkLqE6vlS2fhellQ/IjM2Ukh9wAIpBLFOVcqwXwjddkymvbtrm
RF4+Pxe9BEnNFPbFggZDriDRhNtxeJ7sI/GNI/7N4Q+w6tLkkcp8jn/ZiLMW+MEA
KaXVd051LVCW9E5rnP3DPmyHA3uZ3MWw3oEXUwGrlAsb+u+/lVGbpDT5ZDak9EmJ
s/FqOAIpHleNiOl0MnpJHV6YxTDzKtD5NF1jz/Z8Bj8X+/t9Jk6D4onra5n5WXKK
SA/NjZx3pAB2jM+eh0AQ5D7rC2HSydPWT5LEsfXgvmkYIgYg3IuPTXVhs1jkren3
TN9LzhTsbDkFdroYtjJxsZDzi63EP6zjmojvJT0PKzKhhaJi7EEHFV5r0Jx1VYdk
GiTz/eUT6xOqnlFG3EFOWF9z3IkzCHe3krElt/rjfXIyU9B2IAkJdLuqTHIlKUXp
EE+jNhzJf644xmgnAWVnkoGN1c6gw368r1QvoYwS63R4omZaxqkKIsmifx6W14sl
ORplnb5BZDiALWZdrLHNymFsw/Npkx84GXZ6RS+e/stYlXCqFF1eMi5jkoAYF3Cd
2mY9bMLIwvRxazBX5wgNXCJVsnNGsRM0fWfT2ou2Bn5QVP4tcTLViPhfH9DGmLjK
h2vuswc4AvEaatektSTB9DVOdLOZnpqUWdua9DShgM9eEgab3m43K4bx3WNVGbvs
6DirTkLVnaKnpq75xQg+A1yI3eCYvWlWzz2b0enfzCR8Ptj+4S1fHQVox0ukn/9F
6QzXYx5Rn2+lT69Ph2ZTf1NO0aD0TF69yPwCPFfE3gbLY4ADOcWqXh5+8pROUmn+
sz0rx21U/rn8rUDUP0bDlQAvSRjuBn4mqmx2UOEW+wFwETpwWFLjZA1mPsLlNxaa
EuDiFzLOJ4A+tGz+QmhckwfLkQwBMe1ganmGAryu1JvJdTC4cvIGLkUtXxQXKbYq
F4s9WT0jgbW/ilNRf77roPmZQdwLGsEzg1TC9eEYfQccUOOc0p5FeYHoV/vX5LXU
uqPetiE61mdbTiSnUjQYVV+5r3T1BoxT3mc8BzprmM6LhAnLXi7cYW6/iN9M+1Fu
7ltEqeCLN38PFfGOpGaubdi0zQYPpxp5a6avBb0hkaR6z//YKRICTXX0i4+o4TzU
GGHN2aDyQbG+zgMYLfVltCxZ3M0nl/iPGEUBM9gv0kLqb2QHS4wxc/P4gHlqDj0s
GBMHQOnogLvnwrR4P23kel9R0j8aP39ftliDJvKaz3cz2w5bbBPbLSC8pXdnc7YR
BqqOZ20x15GogaWGT4IGV2j7j8sbePG+ZCCdv++C6hzkzBVWlm2C+hLsxA0KaVz/
r4AXT6DGTZvLQPxm7GZyiu82dWLiSkqLE2UeDWn0nf6ZyVAV/vk39BcV3fvV7uAM
mkOgZJwq6ZHr2f4aNCD3EbUhPMADJbCsRENhlsB4vxCjVjx2jaN4uwzaOw9A83S9
e1oFw+6FYrYe7GyRKYbPyHQ+NEY3hI5fy6ilINoppTeoRR3zPBfrWAQDQLqaQ/7C
8yLe5eMdnfV/g3ssbHXusicQU072JupvZoc2m0nzpgUm+EtRKgq7nSnVDkwqUv2i
6FfMerkblLuytdmIXo9ixS2EplJiMajJrQr0YI67m9UBgPqpAKC+2FuQvvaoctP9
voXUPrhDPnZicDDhsAIALtLGNOBhPzct9rVVeWAPJeFfnUBmF+u/sTG41bOiFzNv
XoJpMWn7om5ngFWxXDz2fe1V2gwkUZMw6icrhst4VczFHcpTYkfKBxYRME/9V8bO
evHIQLxtPFqpNoZFpU9Sobk2oVoafTjQrk9EKXwX6+1mQXp8RyGhTh0hvvTSV7G6
/J2x2PH+ToTZ4hM/G+mnvX4ZuQc34DWhEFcKUN6o3xhOevTFv/VrdgB7pT65SRiz
yIE68CsrkmZQaBNdLEonnz2ZYW6M+suFYsN+s7W0YuRAp9idUeFQdLZlVX9HxfPq
U9TTzbEN997IkaOL/Q+uaMCPIMDBTrKP1HHcdj70uK99l+IPwLOfSyQHMpwjxFNx
xNdaJBOSc7MQzrPS+afN8T5q+EysBs4rRZaf5QDd5QroiKRWdIA7sTTDiI33A0Gv
Y8romSY3WhP5+nlTqGzSmGWIhgnf5wckrsfVC7CMJrAm5j+NRynnX3h+sc2204cR
VV8gdEzQNfZnOyXvZdwvN+izHIhLSNReKBeQly8sIikaBG48yJ3+4YmVBrv5401y
LnT+lzO/Z9l9puGU6iubdA==
`protect END_PROTECTED
