`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Zz2S5AcbesxsmfJj7KZXSR7Xi3FAR6PXFu8hFvrkMxqojZLSSOn8xFmHe46S1w6
GtSGHIpACDpWbXS+sv/PEQNu2p7eed+uHiMjJl+3yTSpA1+zplxKWaaHzZ6oQu+g
U7oc+Nj2cQ3fYh2nH6EnyArcEqUQVctM/s3VFImwtvRC1rD/OMBem9ymhXDMBNDR
iVMmyuRU/h6ibxOr4AiBg4bPB0rUez42PruKPHMOX3Ir1re4foTEjagVuLSoMOBc
4e4SICqIYcKmy69/1mzfa0t2tZxOln7uSrgdAEFDB2Um4jY4ryJgqzvlT437bngE
Q7KdhhB4mUYPxYNc+7VWk9+FNlZJypQTzX5pV9qYV2wypvPyDT6/W+qjM1vi9LKf
wf9y1AAgOytvHDFE4VqFCE/MZ77BtT6MQo7gFbbMv0r6pxuqqvkVw7SykuBSUR4F
fHhak+L1A3KWD/ohkNXy8Q==
`protect END_PROTECTED
