`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVabzzmkrg8jackyAvrfkMAPU3kqA+BvjH0VYWtNP3vd47PurGXJyLX5ksTP5bLs
sBycqUZb1od4/LpzotM7Ek45nW17309MSwrkr7wunux8YBtak/TuxnhzeQUQ6Udl
Y9V3nT7ZTECi0nbFt15dW0U73P1jBkWV2cDGW9u/SDMq+B9Wis0/+IJhivnq8WFI
0ScFKk26FcZG7yMff+W0eq84qYLrqIgZpwerBDPklXX4h/6rIM9LyZPhy+blOrOw
oZszcd4UPGcZvggSCNCv03TITI4SCuI17+Lce+7/2DO+QICeUyqs3UUWUnNvKten
81Y536mmEBBnWGUKsKNSrANzB43KW6IabkD2cKwGD6h5OyaDZqnuGtd3eYDE1wfT
gxj/wN4U9vzvCp82FQO4oqGanTR4YgomK9uPow8ZL9FWqecGW2489bjDbZgullHW
0Qtrn3vh2OkoYWiTjGpadsiI0795HEk87tOw7wyoPtRAkD24A5MCKijJAkIkQLgK
VDQA+3V2Ki1361YgDwD4CcV5IKNbQVKaSCa9BsM9CxoMncjs1WDikHxiYrF7x6nw
h1AyXV/bUhXuC2TrI802ASo6iJqARjnTP8cKwVn9pMpDg5NiOERVAxcmMWk1Mryy
43q2Of9XMZVowmdzmsadaZRSi7wp517PcS2STE5VOhQ1bhoQl+b7T6XLlzHDKZry
fBlbbrXr5YQ3BfZTQ8K/QZWxTh1iFZU1MNd2vRYhlZQzoTlqEt1Lng/KTWqYmHBy
z7passKchdzGL0OwWXiVsFgxDef3LlE9WILrdEHdxvliXUDHnPSaM++etATwn01c
/GTreoWPaKKbzDQDnmdrSQ==
`protect END_PROTECTED
