`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kO9tHv4ZDdHxDShqZnFM4rbdEGP4j75wZL1h3JoaRHjNqrwZzPJi7E8GQjJ4WNms
MS0G6XZScgaQqNChDvYSAL7zHgzom7C9xJhnKMa8f9Xz/61PdLOaJISQNKsPcXLA
PuolTV3zJ88TBikCLtXos3hU1OIsW95K/8r3aSpFI+lfvNXgWKA11sz5K8of3MM6
M5s31akb163i5sBYDteLouEdPV6+EoCRp3LnIJtmzvs0MF2S6D/nuhrb9bYvqbWJ
CrPYtGUoilVYCeCffEUp5FTkBjRRC9xeTrntMInW0oEeAbyaJB1Qg+svCI8gFMsG
EQ7Ht60PsWdTGoD8+DV/iw==
`protect END_PROTECTED
