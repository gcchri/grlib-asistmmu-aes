`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjlIAAfTlF2ALtG2Tfu/rPz8vq3pUEL+prvXmYDz79RbKl9UedqzprfLqWhX/ESD
lenmIN/2r2keaSIrk/UPlzWCWcfPD8WAagNfh3e3LCzslq4C2aqmWl1rpNPqjo41
9EimxVVzXRqtlm86Bqs9jQ/l4R+LL+8GSBCd7vu6rItury+AmEVvwNm1LlWNBcHt
juty7hkWNbueGvE2JKMsfdUS3iaCT1Kp8V6FGRtoTUGHzbErGpaLOJ1guKhPuBfe
tR0yWV2Q/eaQ1L2VmdLs2UX0O1qqsDEzJ2G6P4ruuT6WZGPxwrraBHQJRxx/zyds
+pIc9O6zJcvLX+zXJHkFTl68r2/8y+ckw0Q05h7F/AfoXdlGQet53/EqvT+qHBER
P0LQPx4MINN1exrrfxXdIw4tmkc7Es0iXnd2cTTjjlV8HEkLfU8ZeQyIHMBkLZuC
TA01FW7l0ndXRdfqiXIOmj9XSaEgzdOFDO0bpR5cDfxpMK6u3lP0XUAkOvnIfN+u
bvZwVr+HSSm/yDykWrWHh73rgR04WGwluy2f2NrMLknYUh3Bw98r0G4GWpIkw+Gu
`protect END_PROTECTED
