`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+eNB2+YGEwZwOqwsztfezyBZi7bZa5zDt+6klyk2FYApcV3KVluG1e/Y1wKoMmko
98yCNNrmhSgMi5NejSBs+ZJcwuJfV0T7XgRkm3gPA43iyua38y5dZJRbO437l4QX
oLHAyQZet/o2l6PVY9JXevH2eM/9mTXX5sPz/sIOwMID5j6CKBXEqFGxOrLFyDFs
heFtKp3wZnZ4bxb+wtJChvdpx0UFmVnHilb4ADpqM0uekSWqkP+UYUSo8toDL2oe
Y/N0ldVllZLZPvC/3TF1/Y9WTT/uQsm1JxNLjq6XrfP+AoQX5CWwFQRw6SLHOC4G
G+FKK4Rqeg0mVyCmhJ47gWVHSb7PgKjLBiSBSUxRWvMT1SE6rmqh9k0NNc9dwMe6
EmEaxCxppa6qz0Z0oeURxiH8V72atPX2pc1X5ipniJbIr4c4vB2ugS4i1Fe7NRgg
oHEgwSNFMTyATMxrwiZClZxcmx1xcXkL+qQ3+xh3X7kIdRrJJ+Gjo6u9+GWUUkm6
NKxSWH9LA/UclkUSCriwhEGLap0/96BhNf9yrwSNyVtWcU9yDUJeqY2WaaWZ+6jP
kTUkcxMHOPF6tm5XKJPSKUNywQOYAispx6gcXjC+1hjR5PsViS4osqLtPQ76ZQYy
HJAQoms5YZ+HVHRGeyyUiTENpTJ6NoSqgm5UjJ5JMnj4rUcSboygwXL7VB61/GIr
mmy9jQLfr8Vbge/lLgf5EvaAT+cBr7aWGO+L2jKfmyldezxfyZduy9iC4FpS8m+q
CxOkgtUk1EE0g8mw+49PEu+fAAEr+uJaTAyVFUhVML8=
`protect END_PROTECTED
