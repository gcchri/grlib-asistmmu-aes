`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ABfuUUg5CfKK20iDdX1RvoV/XJpdRs43T9s2ynUGTGTyqf0rIJzvDUgBdHhgZ9l0
b2tZBQjb6dZ7bDh+8hQOfuWn6BQr86G3JEJX7kQCjUAmiLuwHpZfmiTLWJySR75d
9n/v/gUcavsTC3FJT7LK1vKqw5T4cRo5Inw68vLYoMFtJueOasgIZGKWBead+TGO
l2irgxZNTKH/Wein9aBQ5Ch3dzdDsxnBKHcjL94G6thAtnklgDTWopc9JYlZNHfS
tI3m/xX1/eUxSMwjrmpnk3QQz1iv7E5fnZSJfRBWScjnRe0gz90glUW8qOqUGImA
76behJf5gstVjitIduVfZKBifzDeH4O8b8rHvyLX46GPnIT0EDyZNuddZmknIAjW
sXbi9zAcXuQGNniu3dHfBA==
`protect END_PROTECTED
