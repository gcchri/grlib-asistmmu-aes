`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JpIq5g04ypf8OMC/CD49y5Y74882GupLxdlpHpCTRelCLBBsFRvZCFfFCT/7abNK
DkEy+GaKyHX2FyTyL/zM0tqmAAzUgEv1FJTN7N7XcbRNlN83Nu6oY2yJu/ovX34j
eYk8p2jIBwpp+2VzBEAsy+bSCRZIL6dWjPbQ6dZmr+IQCsobZ3JN1nGezSrs/fje
Sw7hq9fdl7IF73vPg+3XQXvSKKLEb1N4+d78yESguzXLrlRnegoinrIO+xnopf79
Bs/J+U1ztE3ReozqxBP0kMaUcFMR//gtMsaWPGHjd+LyzRycQmjfjKwU7Hj+MoE5
`protect END_PROTECTED
