`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPmjJbM8JnW9suVxLRxINcgneEkJ+cTxAzD89APcvjqv4XZ1A3aSEihPJwvZOWON
qMTiiZF9Ceiyp76D6b2a50/ZwAjrDKposmA7MqLzb3Y0deIMk12QCAZKebWRyUVh
hIdatxiUhXrfGlzUP62C62gzyh5uR9ep49GMGwFghgvWiZcPMLuc93GpcATnxThG
QvbfqgBKtM7hYQ6bU4NjWjdR1Vwoq0FtwhSmOvMp+fQbZtJl7R44Sw8RbHBu+1Df
3KaNod9Q53alESi9JWqPXNoI8fYcP0BL2wsz4ThwB9s=
`protect END_PROTECTED
