`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YTFasjW9h/wMxw/QaXHZ75AWoXxwfuA0X2yddiGGaPE0iSzfMQP4+ndeSHnKcSf
iDNduT4ncLdnlYhrfmMa2LHfVWInaKCP7xn6QAvUmhWHxJH2zEzBXjETARWyKrPN
1dhQQAKWnLgdGitM1gA6/31XVy9rouNeyEdgsyOoKqVAUwL96ozrHkP2EMO9phCE
Oq1XrpNDLLlOImcCLwOWCNx+I9WJN/cumIFUKq5B4AXGd0BorB89XSKCu2Vf9rf9
M7UNKjp39lVkh5u+ryWpzyJ0OJbQeONH/gpyQJXscCLn6CL9/2a6OcSDi1HYfShx
yAJScCPToYwcfsItE3dhlaOGw3lFiccLC59FLyw4CInS7qlBe1w1AEvioib1kp/J
lmcLtmD9BG8NF7L8NKFbp2nFdZaTqt0iUKr9wEmmlD6woKLU63hxubp4boFVb8WJ
FjBCAXoqSZ3uKeMnIddSuUm9k36Bl/YA3C12sO8tn2ytqdwOtLRwH2wlu09LjM2k
5o1KI962Ps4uzOHbJHhB+g5WYR5CKpKYA/RqawJa966kKsieUI2wKNLLi5aX0/fW
eOS1D5u/2tCFjuvD5+Ri+yCchs2PYSzLLceqof8xfwkaWO82N+UHkn2ARgQr/PJR
tW6heU4X9706aN/2qqw98I9MgorFwjDEiStzGACnSS/FyKV3nRVyVKCodVmAG8TQ
QbrPQceoOy7Hq7WjzZ8z3imbs2sI7CYXuHDgk/+vgjcA7jRisBGnfcP2/DGj0XuQ
nADeETnT5oKu4jQ5ksKEmzXyudrfWm2xEEMy0/1IMKY+ZZGFix5bAEniHaviRmF/
tHbxUvuAhnTXtIIfqJ+HjoPpccvqJbAczEXJPOqFmwcnQrMG6kKS5S9UI82PRvSS
miKMmoYISaaXJ+A31FHGnXNVelrj2mWcg+rBWWFVO8MBCM5C6Fm8jt825CRvRdQJ
KyhGgdo9PULbgU/+oEMsqdfwTelgFrwpU3izfy66Ob+vrA5IX3NXNkmn4DtUPGaI
+n8fBMh7fbRiMJc66DSiyyvPvF9/pd9WH+8bl9McRDmRlqv0sA2i1xbd9MwAwvwd
5bqq6kyMKMEPuK7rHzkuaVVRM00vuZO2ZAidutrmjD3J6+JneQCySDcr04g16tSA
MBzoWNnsxRj+TUQZj3gRVd4dykhDYV80sD0j30B3fMMQoYQxAmgquanBc07e0MHA
/uvMPqSAWDR53GOA/h1WMu95XCcnCbEaMQYeXv65juecoX0gKW4DJ/6ISYNZSW9g
nwygpgL5+sTXNvLhWyaI8TAqlFd/v3KWHFWP/VOEDWsecyOQ8t8zjLTM+eQT8VWB
vE42qd9vh61xBTM+QRpFOgdFJch99vX92/+tMa+tFDB2sfwoeq/weiPC4FiHvUkS
4a9yMx47aHQH5r+jFqBBzwdjvhkNIKhDCRQPDymCFIHcvixDG+P14WqoDeh7tCpL
6ZM/IS2q2uLtlCiD2ZOQX+DnStgbHbRd3r70F91Ppff0MxC5GA1bStoRp562cW2j
ROQ29BUNGbKQPc7KnJ9L/0yToNpNXj/8YUt8Du3WytjJtoPcuEbF8S9dJjG41Jal
Ph0hlUBpKZZ7+hBaRL/YCbOzrP+zj05j58f8kFp4ZRPEF+NnGklkI1vfiZcSLcMl
uJSzSjwy0z1IBsWf8/NmU1sQKEjv2lTV78ct2KvxYwzEHRcZ/jxkPfT+7fMaPGX3
L6rvqWaiIoMZMXnhmx5uLWL3HTZvRkM5XHNy6MBf/Hk+Z0TADY3I84u9tc3dehfr
feyBAv9ZMBzNg/180Np8LZZUk1i+nmktoCSyNlUqxsvLVXXHXfvtndlq8vLl3ufa
9PQ1cVxXbUpcM6OBOrFf3lOU5yofz9At5uyA7aom8mcnObSzibGfs6nLbIPxY59R
iw1On/QjiTZcsQMhCstzeUqSj/EDzF2qIp7g56nFyOLF2G7W4IqJLn/YkFY47fG1
c2o5Np06s5wzj7dXkD9+z7td2fQeKxVrrkP+IQMmizF5nbwWHuVoc02mGZaXR4fI
LndaaaWp827F6Tv76Dm/niYLFG2mNGU45Gy5WlAAjyBlMrEVLXKn+8BQKHs8gHyu
BktfWkYuRSUO8X74Dvzc+hxZa6NA/vIclkTRAoUFyqVbAAsnFiwqksoWe8SU7/CU
cP5+5jMUnhZSUm8xHpRkr1Hj4J0jiDD4R9xVSmM2EQCnKGP9CQmqGBH1eqhMTGHc
3yD7Ge58XDC4/jYJPBkOGzqG+1L2u56qyWPJ4sdutMA=
`protect END_PROTECTED
