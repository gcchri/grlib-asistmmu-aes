`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WW5mRqkDrjTOiyzd6GU/wnlKBhqy9dt0KG2z8ItpIMP6AK5KtEkVkzCp9uZQuh2g
7fofVZWqLS1dumIdqCViorAp+4mr8xlNGAcOadEYHlJ5An4lHCKLo61eF7GxEgkL
kCC6wvxozAnf7xZWtAZJCyaUq8xrJZBFYlkWC2lQsL9ljQW72XIDgq1p2cJ7bIuh
rO0+SNEfWooBtD+M+He5mz+rzhJPIbCgYSXTaQUGHPYEuqflDCV869zuFl7kDq5t
K4ozmlIFW+rPtv8On53OaqA+GmxW88naD6SyTdELlsfRl6d9qKCG/ovZ7f9xARE7
fsagoVLUKriZBBjlo0TYCOrpUAeVIABtSDc1kpT+FKc=
`protect END_PROTECTED
