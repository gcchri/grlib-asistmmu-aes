`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8v/UeBZnrPriref0hJAgSg75wxkg+jPdYfnQCNVJuvxzW5pl68onQuNrcacifZks
C0RoOXN5mDoq5EjCaKMWOU5pW1cjpKBgUr2cIuBe/NJy8uri2bOeXMx5ei5UnLYr
JR9XhFYy8Z30qCAsAV0y1V9BaCSe1nov+eeawB2M67LtHwvFDKIxv9ZlElbkV1UI
5NcnxXuURmGfRatmNMpt39X/64nm7pViGA+kizxRTGTFWxA0nkggp0cNXptbXPtm
/6P3FxHs4CdEw71u8q4te9ga77bMfXML96lKPIiIWgR3NDGCkSgb6T3lcxcsrEHp
E0qOIgu6UvsOtGZFMSTwLyCNv9yFvdYh7w/l5vE8Eyeu6ntbscbAbE/Pw+kveV5n
ntRNwmnVPqR0ELOLz4GwFyM3l8EXzE/2UOq+ezZHv7Y=
`protect END_PROTECTED
