`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yU/vINlKpruTXKXg4gmuoGuQR/mN2nzSuQj/FY+NYJ1EleYhOizPgPKAkzBIQHtt
ZkUt5guW/LyQayw37Ab/9E/chZyjDtKoPBmHjKcL16IrILn5GV+jXDVchUTYrX8E
IVEogyCCbfP+u9aUAySQZxkovA2F+NaE/18suxkjbm/hPjv8mSCy/Rt4DMUGuuXf
CA7OtV1wzo4spFq63Q1/xVWCffI0uym6lYk2KlBjl5ss2eK/CO0dymXj3M6uqV/7
7KvwNOLqYccKqrnPqmlhX5kCjQleYcxC+HXkhbCjskE+DvTl/5xj7sapOSLsvsH8
pntuEdtBi4bQWU8tLKnKeJHZZoRbBlWTLm0GYnjYVtb9ubQ8mRndtYBG9lANmXQu
UmkWm/0CBd2RYYLsHtmFiR2vCHhsyIB7naLVAovbi8/SdyGdT5vHOeUhjHN/EyWt
FwtroygOOKK+3vBfZCRBlMOKFlVvhYn2wQfZQ689nHN2+uqdm7EThkUW1pJB1kGd
C3gdBTtZUq3ak1pF2YUY22JOtr0Qcerb6TpVcC/xV8IoyYCGC4DJ3oNqiPr3NKss
X5SUVgBCCoK7W9GMYHmZ2lY30ucudZIm4jaTsoalTxhKRbPXXfrggxw+AAzga+M9
ra9jJbRPYKoha/xzTXC8Ri0IkOaKzh0Kw3vzR2xMRISxdi4nx6ODPxBKFEiGs2aD
CnQlkMBA6oyr/fUNbnY6yXqoEPbwVkRWFfZx8tNSt7+DWyp6hqWdWhQ9L/ELqO8K
XoAXxolzlgFKCArxwsSwVHALuIj4ItGVz5ihsqurKA3stufIqOddFAADcxgrj+e7
RX/WmX5RyRVV8mDnJr1BhXCm6fwqL3R7sldVCij1QzwoF9x3ct/CKBVhYsIvuO5x
Op3bVZqJEJz7GvRW7t8uFBikW4gwPZrTJsHplvbPmvMIdxL7lJlObhELt3Q5GHZW
I53qxIR2B1DCeOwRPvITQT7QhxpnrM5M6hTmD/xYq6vIozY39t7QGkhcwR1IwHAS
ngxNqPisMa7gq21AJJnXFpzUIuQchtXislltw8JpaLMVeQmoeGboypm5Po28MLrc
RWiiKGXjwFmiGdvmr0ZJiPI7w4XwJ+7hTWVkv5RCkU7l9sKzcwCtSzHM+4Alnlff
gB/Bvyor+n/nsWHjE+lnfrkm5qwnKbBaO0pgel6LzadnL8eWX3yS9p+VF/T7RHix
mMwlYZXT9UuA1q7+peyLx9I1CraKjwspyCyVPjM4B/OvAXqhNOob6H3L2ZPthnWo
qZ0oPxcAT/lzJOgm94Viek1K2L8rahgHN84Iz9Vo/gMVgLMZ6sNHR5QjoTQUa58O
mDWIpgMVXmjzlW/2eLF6zpfRUFTgi153IEChobSAQExwl9DZO2hJfS0UFoC13gOT
2yAQ/sS/u6/RjeEAxFDS0+Qhh66SYkXYUQaGakZS4gHxu3one1xbXu6VFr81uQ/Z
ZHBL85SmI5hN0cZDTa2FOpztzVYMxGd+7OdICqnx6XgvW9/ncRJQEOdFdCCGRKqY
wt/iEth/v5yavD8UsIl2Bk1G4RuvE1AVZ+X9w50hvgYLvfWUE4qR4reZHEk/lihA
O2a9D5GI6up8iOr/TXhPNGL+FIe3qZGItx0aCABh8RRecC4I/lHumYqKTJzyoWzm
CqJHSmdzUT2EZYsFBwMcZrB3LhNZEkq42sXaIrGzfO03wQpO4Z7FepuGK+qFtM9i
Z+h3LGNvgSmAJSQzzIJh8D65X10uH63m3LNwNzL3esALUlLFjtkZ/AytCdoq0AbL
tzG7sSNgvegftqIY6ei/+zC9c5JKJ2Ju12gEHP53evPbujZ3C4qYl1iJniFhMQex
hOn049wO1Jl1yPpJCKPzCpInzSSyBUqA+Uo9vrZtOpDggrKPLNb5advXmc2WuC/5
jFjyBcbGIKqYXwuu2XG0PVp1jcoXj8QAxLpYeXsJlCUieZhfVgpHmfuMxDQrCvbW
TF36TCsXuGb/5nvRxWNx2gfzwy0iibuf9F7k0t1c6MQ9CGz+yrnC4n9lI+x45oib
wpRi4qK+7d//lieNUpxvZnl252wPP6DorlRsTkgxWUb7BoqdcXWSg+wS5ppOIbpi
xhB9piIOgeMbNS2KziLTKIBTNrlE8AQpWtN0EpanAtaIKLCK7Xlum0BS5IgR4tLv
cKoYtXkcqO7kvg2xquFCylOs+FxY2UeZDW77L+jT3o3wrNNRLQ7ehFqgYY11cbD+
7pqqOvwpsOIeXM3t84nzCK7jd5vdQn3Ta3NhO4jrv+pYpxPxO6y5ry+NX9I7hmBl
FsM+EbVRKt+orfb3LaKL4tRk2wbT7S1eygxUJC3DdqQ7uneyKEuw3tOEYOqxBbIq
R364/ls8Fq2CZBhzRkbvBx+JxqPEwUct4R/QqIYm1fOdLrf+oBdxo9crEyVcPdQo
F2eaGTnpJBBjByqncTvdL340m88g56zQ3OdFi742UG3rfDz47Pug0C1oTemScwv5
H8DQ8A22kT0DN/ZG6GCHZg==
`protect END_PROTECTED
