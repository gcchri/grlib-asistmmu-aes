`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j5atlHbssKj8+F9FygTLpBVYrxe5gAcYuXm7m+VRRbSnQrykJ5i3uBpNdgpSaqQR
W+BtUJ2/15g5v/Mqa1DAq+gcMqFhICaIYY/njIpYXd9aGvOJCj9KekXduLObnIpr
0gnHehlBOR7duSYRO8fk7Ov+fTqMTxknIMmrvnE7KlmZGGf5VI9bZjpJhMe8xA+D
QUIllMxZBfgLahecMnJkbjqUmiEVfCoy5hi5tf8UL9aJeY8MzIHRzfMW0HssZrpL
H+Av46+FJ7RVchUyJo6eURDjwMOj6fKP7fP3KtesVuMNxnwZgrPSX7FauqRTnd4R
P8OPIIsOdawGuOPkS/FLCyPjDJ1xuqWLbUSbv4EqwOyTfgOqFpMNWT6awO42jIwD
9AzVsY1Dx5beo6l4g7Zwso1f/2Hh9PC9N21qtoQ/7pECdHZ2REi2f9QuddyO+c/C
dGekk1F2PazszIAuVJYAzdpNVmhp6vSiI/lCO97apIUlHu/4nessNF6e9UG44DIs
8Tktf8lY2Kj7u2x/PYCF45XpbR4pgftIo6BiaJlla1cVqaFANcixUTop/Mw5I4wM
UkqWkXCIK6hu/mkYKXuWEfCGldb6ImA8jqF6GfpJFxmtO0Cyeh3AWdvs3cDZOxoL
XAzfIbvJeY6X2M/Rozv82yVVS+4qlB6KmY7OW1yoFfK7oPO6HbSqfhJ5Wwz6d1BU
qfy3ZRnq5iLqho9cjD/HGw==
`protect END_PROTECTED
