`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fiZzRJzflb3dB4I/9HhXN6amynaMQOJkl1E0kV7ZE+IxkAhfuhfOumhEVZY+sHkn
90sGTH77JDc1vc22+uNtvLhOKg6WWUr13AJAFw30DurSZrSj+LGMcquCxd2RDPBt
d5xu/knTfWe1qcEEKzmiK/DraYpz2Osunx1YSJHYVZGs5JIfis6lVxEkJNc4b10a
jdMKScK53fTCSQdjrpLhwnuYCk7WN/HXIxNJcunt6QShoWfXWJ2u1olaNJqCNRRh
Fm1xmJ/M0lvTeAmvuA1IrC/G1ybllz/id5Xun1Becls=
`protect END_PROTECTED
