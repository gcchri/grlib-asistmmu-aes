`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L2obENKfsEQ2fpBqtYlWcGdyvrXF+AKHf40GYPzI2U0SjMjhUjBCtRURgcgdM41Y
jfDCRIEbPKdFJddnPqSkzc5YEtzYW8s5F6DmymaVGFuN2RU+hwFilsYQEatKPooJ
Kzg1iA+++oPfulFX/+psOuDwakEJg7hb5r9mzSHm3uakVxLsgc+PyyiOteiSsw2f
EUuBaLC20CCx5+A+6Hypoo+sE2HhcGNMGHhggwNNjcAJL99vD+ovkOIGyS2IMW+O
WcGHBWUgC/ZDJp0lLevjgOobwQedKhiv2/rprppv3hLc5XR5Y2FJnmaCu3LqSyAd
x52GwwLmaGZFve//0nEPmg==
`protect END_PROTECTED
