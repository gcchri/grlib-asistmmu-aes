`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mhptcii6vE8tEQHKUPNTbKkCghz1ygvpsvz6Ndox/12da1Tg31XAIc1E2j2JRW5M
UhvbbK+UOQablvxgEO41nLBxdqNdgzMtdQ3npUNBmqwfqGuYfrxPjZRA8LWBGVG0
VASKp1XwI3XFCDooeQXIZTYXSuQrU2eAPcFgZLRa4JIpM+VKWO0SX2iAdWsvdVvH
HAX5tqmUl+2W8y/ateVDpeiYCZJLbDHniPuhgpcKBg5it2l91vlbqqjirmG00c6m
Uqs4/Pxe0jlvBaxAb61Pc3EdcOGgi9g40aat9UWiK9oy7oU2nM27McnXqwkmmfH+
xHuP0CZxWnbGhD78AXFMxrCn087A5gdVwIi75kO6WlgRy4Zq5LKDsFU+hj36bgLL
gFXX6jewoAL+3SNUSWoXxIl77P1QSSd6ikVTQTQqaEuxgSXInPsXnHW+ub/fTsXJ
aBuzAIi58n4gWAYLGjzJAjtlRyihqkGV41viODr3KZSFCGgIqbcLFcrpGkhmzcvj
w+dXUOfNjIEE1QUPsW40IGQHwEU01tXvM9+BmQBYHFKQSCCVrZuuzzaTAlGLdoMP
6O/L0MFtLZllYm9utxk6dvO50QhrXa8NoTUDdY1Cy6gJDProryP8YHD8RDuDr4Qo
xDGkvuHX+NeJA1G+3tJgt4WykbPTb/4btBMBe8wbMN1jUEYvuUQBJYVGdn0SWH1Q
lE9TtG0AnFjThHc4ABo3vMzyntCm373hpL/N1j7+4sclRljPa6KlhhDEnJ0vnxaC
yoERcjkQP50cdlc5isr6jr6FhfutRYxUtViqmTOcLijdsGhlL/Y+505HWbenxGcE
uWEEgi5ouYi7fwygx3nkyEAB/n8FLGGm/TEpvq+++38IQePdUwdZXbf68B8Hn+un
ZRvHbdmit/FcfUNmUx6SLNOUtw3ImtIR7x41gHmLngPHWEO+B6GpqbjxelxAc4L8
ru32wufof0To7vKHtbVN/hoJjnvvhRddSIDU/SUQ3nXKaI9SPfLi0eOqBUNpJDEL
NXOQ3L1OTs05Hn2bE1u8GZa2aIJoAC2jw5oukXM1ptQ4wVY7NtA2CQZ1e+5N9lL0
sXnulvxpmEjMkgevPNJ46jYiwkzvkzLH2Y9W6YdJho73+cMh2KUaxkomsKSUONBo
Jv2mSlMtF3PVJMog5a3MJsoBDKlZmVWHXeq/r3FCbvS+4C/ukVE/mUQrzuVosPZ4
iCvVYFZXBdAWdY1lloCrqXTn/TtKZpBXpEFQGrYMrkilxqbIcultwahT3Z7a+xqJ
qa3Cw1ESqNNG/Sor0knCXJGFG5/rZ+hfo5xw06lZugE2X74/fI9XFo/DJn4mimh4
ZgxeuTBDsFQ9QnNLpMq4U3pM+rMK2dUkNsBOAvjHlHpnEb5Rgvk1Psqd1F31D2Z+
tzBZbYuohF4m0Kyzdog5EgzKiO06bFuQNO3N8OLh8uMNE0o4J3jeYcHbeUfJgqDs
Z1/c0jomRWhKzanodD+LDAKdxwpUAqU+fgUBnTkiH5MEcVGJrIaIeUjZTvNVYty8
3SEAJVq+rCPLmsVsugMxy1GHS6s0omh2G+9oMI03ic0Y6GOcbXeHtc/LRTkwnhIP
rakU4zfXzNmy4LpYLEUinPO9t9IQMEBapFtELS6weflbywRHfuqSJ+/NIoHxUz+h
/o8X2rqMNyL66t6E9PVIaPLIrKoQlisGmcEJO4ZALk7t5PSsudDW1AN0QhTxZdT9
pRXOxkNDHv3mRiuuv7yVjOnBKGrpdk0lCVRPVTxOl5E7u30wMAckHKEd5zxzFBAo
HXIMP5tyASaQP6YTqZTovMskzpWQadzFdAgYuOseDtCRVjO+/nsLzvRyD0P4cVUO
v7jsnhFN0hjOP/NJe2EI/CEMfOzMm2NKcHuDBUMMUD+yriPxIj27K7o6tE4Ipr1W
4ge/VYgBaEsFk/ku0VXvfFxHs0zZP/Ub64JHYUjrMaIM48HgL1YnTRie0G/7XMd4
ib/cvAvlaJHuO+XN871+kUbNDi3gsOh0163S8htC6Uc=
`protect END_PROTECTED
