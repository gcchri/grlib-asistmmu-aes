`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F3imnC/Y6nbvG87fl5P18tcjx3340jxa/Bu3X4nTp2Ne92ibd5Q3L63IH1skjaFa
VSCY8H5zajD/ES3LdU6EUYCBfPCsFWMmyLR6BvEKr8fjuNRYSKJygp+7fSflAEPm
vTGGYatCx1GLQsTvqXssbaOoelu8/jSe6Rsw5vztYI4fFJeQ+aFQPh3jOfONFcuG
UNRtSeNsVTJIDRf2k/v2PbR/ff+Si1zcG8BM4X6GFFW3TFQRHQHvpoP3MX/IbuSc
3yMJsJ3+PSJZbI9hXB8CEZ1Un3NwkcHn5LQXxZXnvzYHYWTyQbsdbDRHOIDPzlHJ
Jzja/VAxU0/Pn6aIhzI0gkOrfD2sZKCpfGIEeT+rolVRlyrWOCMkavSzQzALQ+qq
fqGpNqPyERUcPZxKlAagAyNOSoX/i3Qx7vB6AHmTNjQAXSgL6nmvj7MH+tPfF0xW
9qWL3btzWooL4yLbbmRZfQ==
`protect END_PROTECTED
