`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VtImFiqF+8d64NFQD5YiMUOgb2jZJGVAvmyqcoTHPHb3f+0BS2Gou7jsxB5PpiM+
+k13nsrMDmX55dId3oUL0m3XHZ9nUdt1GVy1cQbTA1vLRko6fU3k/nSXvDbIvgs0
MGr8Ve1mBtGKrRy3OEATIJBdx8W6d94fewzEamjTt1gj6krFigdftaZShLiaWPR8
3lJhmy81brUNw4OkWn69j+WGJiom1UijIkHucKg7LMOaCgihPlzpyKKJccwMLT+L
GoC3BdE+6clqfldAHXyRzrACK4g9d97x++AA37n0LroPPzjMafvC0+I2XSSyEbF4
f8xQ0khOCQyvX6VQWvaAJej38YiVjADGXmKvj7Lp01AKKZaCcsSv+JdfWjn/1cTX
NFfPep2/KFL2DvFMHi8Ok9FdQSFopcnXw5tKJeSyWBMeXzwOg8amozFLSqE2mHwO
1AqQSuw3tYolJgaHnKal2NF6X7KOgbV+FW7kNS18SCbqvi/iNs02ilRxsgy9colo
WWiXl5VfJbLwQpxPCWe9XQMSbLVmseKdn8WxulFSOFKqiL6z8F/7t4jNcMUNkCvZ
qJPOCl1Y6QxLA/PHEN7fkQbD7gt69V9T4SLkzsrG10noNhzRfNvhSCNLiNRrwvbA
/cj6z7CHIz7tOfb5FvWPmZ0xYu0dws3BIiPYSHFJOhMoGKI7q05D9wIR9MlLpxSX
jxAEGIJPq8NSNMjy8lagJbGv7A0x5LEflC4ICohmAok3j5XK5sQ4y6b6mKA2IKuf
hcH3rWPDpFVwvlddUtzgS1KtI00ds9DpxmO3aeWgpvlS26YcrZYw0TB2rx0pHSD+
UYCKemGeDU+N91efw91zeGoMAQ/cEPioCxHpT8Dn1IPmW/eilDXZUHuiN/JXZAHV
fOVqzp4zP6vNyFdmq0B6voPUGisttDNQR+VwQr2iGiDrwhH786W4yS9A+me/bUr1
bM7xdJLutoKEWOsaMwpEyi6lubfzFMeyHzGVqQhXLMv3/cwm3a9jGzMZQcm49n+t
DiE5CjJSd8Fb6wOE6pj2vmXKBng6uhln0fkr2cuc6dS9ZSpU1JZAbhanoqlKgv7X
x4OFxclXvflxHvftWbZ6LpfL6LelvqcL7Ww8hQhO8Wr1WRvQf04i3xlPyohi7unG
y0T0LnvLpp7bpzTv+w1Ijh1Dmls3mPaJUAbCZ+u2YDEjOlpL8ncCYuedLo0Kx86t
H7FIyWuDAXnX2sPdbUkEfg==
`protect END_PROTECTED
