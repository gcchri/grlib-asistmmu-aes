`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EL+1D40MABfYonFWEm79gdb52ER4xGXyRp+7La5E4j3DKX8dXE/30BM3zxGHXYQa
uIhcdKjeDK2GUJ3hDakocm+w1i18qJuh+2gEaR/46TNcK+mbGBnMluVH5IQyk89N
RWzktQ6oVSi9RqGj6n2jBGTUaLd8y9NAG9qZMxiQvBkPV+w4SUTmgaeN5n9vod/f
zXH0Zox1wIU554Lg7rIMJbznkXHYUk7+f+ZMvgw4ZRqiFOXrq1x8Y07Tzn3HX/xE
LBuZv51g3R0jcng5tG+69LFoUxoQFCQtvC18dD0m94zxqbwTMA5cH5HqZaPsJQHr
2mxh28ONa0U6QskR7Z4H/BEgnrMPoNE0gSvJ/jWv4YM51IxakxIa1MzlSm0S1U8s
9w4Kfvt9UkYJl9rBBAdHSOhJevnkDVcurfbPgWaKiAaL4WuYD/XrWV/oQqAXAj2t
8LQeTD5Tj9TJ/tDrkKmdEt3zlwP1VjYnhKm1QVbc+HvdbG2jX9uxrUBOCciOWyby
gIIF+Vy2oDtsOK3GvYKiSjsPI56K6brg/xnSM0JEDA/6gnL8w7TPgoh9mAORpKWU
1lUrk8m1JOQ1F87yeMiCNYvU5SX6zXGT8yQVadI+ZNZAt/iMzEt5pq/9LLSHlsaF
X6ypajg9jloFn9J9V9iAmjB5q0+KqvGFsyV6GWQhkqmCdJgZPbsyINTG4J0SWS+3
/QSQ2358Ful/daFWjA8XJfhjUnvv4O4N37c1sJtaU/s5PUMb9wlNokt/nxAZYevB
3PDxqibvJmyLFzHHgoGH3A==
`protect END_PROTECTED
