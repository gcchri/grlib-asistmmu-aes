`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPmCPKvcEnEwD08XKbdoyn8yWZPsq3CJbIsx050MZEE/Y6jxBm2uv5Z0ZsQeLttd
MqEm9yC/MOn09G2sC3X1NS0AX5mA8LI0rhiB+qc0Gv+KypFRN0MZezeJ07krBfZu
W6rdxYowgWmpCcy9EVPv4Qaq73IflUMNwtCeMWV6mdGdkO9I2ZxdsZhGN/bLXL1a
k8SfCQb/JWFXeRNcytPtv2X24WbWlizl7OhsbKxjsSBRVDF80Ff8neMPDSNGMuz2
mNgz5TAZ8ICodUcghZpU/4E9TxWAwhRRSihzuFElciWRZjTAKiH/9JEj6PHxK9UU
ZByDy0W27GVZiJ/ox1yQlzipRw2v/LFfKeM1zkYxDiA+6R9b3gBXxzIQj4bel/Hc
gwWIg8mHh2+DkQ/fOtcYWn/ZGQDaHmEwZNBBeO4oa56Y+sjZXw5rlNxijpl12fCK
ftYl7NbMI5B+Z+MhM9j8ay+4MAsILJQf+pUWTlez15wbm3tF827YRZIDm6syiT2q
1PvMNOplYC3/4Useh6GCqsCkjC+OkEKXNOSEK0LPt8GrRryjzdpDdQN1VJAtf6bj
7VTcDgPV9adFjyXL4SxyvP+CAernKitfJh8FdOWm9WRgWf25Fp9oVsOYSq3dAcDs
woHgQUlsWgPTzv6VFsJ+xpjBt501tWSxXPowxyhRIVCB5Bb6acIH5isH7Yhb2xPG
6t2xBrk4p7PJQuRPN3mNUdTxs6gVnL9fBhlAYnMWe7rrFrV12GaY7hr8vK/9owOZ
dtOtwxuHK2PPAMKn/bAx3ArbgGAalCaSmL+HtYTO81NXPmXOErFX6H74DXWAb1rs
hiEbx2QAnlQ2ofzkxEDXkB3+vpFb67dcYkBKabgTYbg=
`protect END_PROTECTED
