`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MfSkVbUC76Y+LnilI2xXSBq7pGK4wECOm1CDwWCzl/9EYFdHXX+pVW1qZRBVc2KJ
eqhwLFTQkuvM35+cNMtEIiCht4cNXDKuJSPIHszcJZPNwNXLZDaazijwD/Tx9Rtq
uW5kaXQRyGK3XHJOP5RnPAvq4vfEF+u28PfoY5VS3NLHJqL1q0Cl3am34jF9fANB
dYL6mWcDOFlrvbQAi1C3mXuyTeYypT5zaWx8UPgUH5l++rkzjxDESPjARNXBcvHQ
ZlQOqJdYz0sH5gPHsjESnxCLufBm1zlyYJeMnJV45o2Ae2fF2J3m6tk2WmeSsO6N
McB66pOp1UpR/f849PGZrN3eP53gJYEFVAr6HZALB54Ci0aSQL5UySQwWL0a4iBJ
cHGPrdkhN1eFbzpUKA6vAXtZcFr9/x5NyO7XoYAuBy6jmePCvcNZFhNUTnqn2evJ
4E6jyMDe5p0RI+RW72JsV20nDiuBiz6yN2h7STx5w64wTyP3zogFJ7KUUYNvHp/e
3dKrmel9htPatUc+3wDwyfRfJnhNm+xnL+knjNxzhCohFGnKJxCMWcVa3Y7HuCVe
kBlQIt+/hoCwW3gGqDbCdeCCFOVCw31rLt84cbaT2KM2YYqx4kQAofldTzFJ9m7/
T96nxGcTqGGugEF5DIDsR4QC5SmyDiLnQ9rHJPgI0Y7N2l6CCEdi3Otxztuy/WJB
E+9xB+rko9oJPXFUe2qAHIC0Gt3drtuUBPEjNAA9jIrjqZOWcSW+hAWPxmCdAT0h
002qfQDgrT3kfeAgO5YszWl9IAm54XK1LLYG0XCNugFcH70urr3zAyJ0C0XMnPCv
OC5WSPn5jhS08yMlpxxa8ij3vf8SkGWmCD0hW3SOuR0XS0s8ptYBFrUUDtdX8d29
9WU9ACFYlYfiaNKjrU7NX8jMc1bz1Z0TCUjaoG8+nY849Tmf9s0hUN9N3GeL+e2b
TjTggKeQCZkLOI/MOzicHzOyR/yFkp+AL1nglEQFhN2SAVrnO7W9hthl7c4AZsTt
qUYc4XnOd7mwlKA/9tH4r9NDtJfZSGwPvKqIoHNbOyy3f20YakhL4/xLOzcNPNbD
2+AEoKsbBu28m6GCTbJe46fwmMBKO+rjzheCw7eMbv7IHH+vf6tI9HFI44MJqJ7E
ou0XX99CPeDPPNk0flrLXwH4tfiyGNJYMi/g0stbPTuK/Z22JBAM66LCyiVzqFhC
K1x2wVEd85MrmJ35HGmziwTYP6EHpxTEcA948DrUlBhkpbpklJZvlG1h5WavAES0
Qcj80bbtl/Nr0WtbghC4/cko+t/UFH9z+WEDJKUP0XJ48Yolger33yAe/1xDckPX
MV6th6iTPfOi1za03M41bYwuIHfrK3czeUsMN+i7PvpUWGwxROcTWj1uIx1LrZj+
ewjwVklBK148EOicy8EkVHb/V0n/eQB1uTGUIgLPp7oXgFvAev5d6wr3MSaWcw4T
c7IYCNq6qgT9zU2BwD2qUAxV6lmxXlcL+WBs0H26yN6BB51HhrHJTkmMH48JJRoY
x0+qlCOShPh02JG9Pw7E59MkX5ahF9KRcvnKppiHMXktXkaoNsjCa9TmsymEmoyX
UBiLuqAt064Mkv+bEJnA/FDgFYBO4MOILRQLzKfnok0BwyanpuVQVxA1C2fHoxV+
J40XvlzXqDVm1q5ZoY8kcDXSdb4JMRJiIgzI2rvtR5BviC1t+1VLW/xfp4h772fm
JV0g1+oLprVJ/OLZfyRBZTicMKcX7/r0zT1mX86FTfX/dTCBrysNTLIMlsQP4Ns8
xt/aSCddAaS02pjNmA5rrSfaCcgGnHEJyxX6QdAJLgBW0GvHR5MtZYs3ABZa8wNd
5LoidpfSBgskYhFnROjL3LnYcLee8jtjLp7tlB9hln71ON+vGLgZTHQ7mj9fJcrR
nCs8hrik8++kDRnzImrwK5ygqoOxbvs8B6xmeshwOMgqTRN0pS5beFbHRCnBSV9d
p3CohmUbNjd50dgE5syintiKOIu0Mx273O7xWbYL1yLWntFUoty3LueHDfnVqd+7
Vzw0BnBHn6B99MY6xqDAFfrsZ2n76wR1HKMK6/NzEi2RUc9QuOZIYDl5gcFPtNHf
yKx80ALC3M44UDPip0ybzX0fSU2hfcJK5BE3Cf1fIXYm3uS/8+UryN4OjZo51Ukt
PWgZG3pPcpU7U7qKIFriGZWpp4ZER0PoR/ucS94gDUAOTEduOZfMrvUI5x8HFV5u
uIpS6j5fJMKzkhJ9uGIjzLujkMGXTah5P3lWRiy0Ne8XWHQiOqcWQ+N/pl01ce+m
czeHeFzOpX77ck8wVN2OO31/xHezIe8BmH7opdzgcp1D71xD0Th2l6QkwGMepvbZ
3hO7rd0FjDgt+RpoNL/nOpP8NPtiGWBy6QqPlsTpqUmKEEhMTjP8QVgibLMD0kuK
FlsgaOGDP+dPubk1GYsgmTLdH6F0nyK0IKarmjpjW0mNRxgdsAKZ+G5oKPUSIcMu
rqlV/MaSjtvPNOdifHcmamuOdgw13pdZ+JjbhEwzcB6V9MdqY5IHYlH8lFDhowcS
9Exx1AfQVTwbXCU1Iqki7nmPVgEMJxNHONgp9TItRtP+0HUTmFVlC6lbO30JuYKH
WzFR7dKO0KYMMywt+sxmhtpcmCc7H+dhEtGeovx/u+myNePNQwneThSR0tdGONXM
ZQgLzisb4NqQJ95blqr/QWJxp+gdrq9060J4yLVhihLS6nT3WO4abiyb9CMx8rMs
pGXJtp2WdZL6/ltOO6uqGGPUFDJ5C91T+553SFZqZoCKafA7ldftMWz9Gf9KflQG
5DWi27gFou9mmvRk/pVrQ3N1sb8HrpUAnGeZ/zbQhOWBc2lWYq/A8Fva/QPp1OwC
w6lD1sHZDqgVrXKEGP6j/zpl8R7D7bdIzeYiJ0lgAsKUNXo4/70b6kLFzATeZfFJ
XVQkTgGcrKsRuHoT+ztFfKZnYvrOZpxydjvKbu6LEM13c3OGGpITtwaCDV7AvJ54
bnkqu+3z652psZgfwXt6slNXRiomA3Uj/N0LSyEXWIqrfXJ9Uy5OMO+Vn1hp+YV7
K5MLckP0DTbc88vfuGIicrDRi2O+y9D2aCovjTKKypyjibGTEPn6ngUflMk5zcQf
DCcRs5JvMfjSXwyV1yxrNJ7XQ/ZhDRjH3OaZvlwK5JPMUrrLxucl3XFd3ffSVTf/
VsTf6XcWHpvVH8kF9kKPGBH9lK2NOVKB4YnodzbBjkmXQRy4p6ZNGHUzaTWEeX7p
SeRe6Dtag25XBBCrtj7bBsPfxXp1svki//b4h1nOcW1XqUCJ35apFRiGBrX+9YDd
FcgLSLWy6aoZEyv6hdHbk8yMc7nFHFEXDx5oSMNcexabMMIxKH2eiy70wp7xWlqD
Edh8R1wBpBoC0gS+gB4JDmT3dISi9UpdenzBvROZA5Q0DfsVdRN7b3byvrY2dqHA
ghvH/noVmmpUx2Mj7eKBikICwdVe7aYNYxjUhpiPehGDGUr715bcf83B++RTza3A
0N+lNMeFR1OEaQxQyc4AM6i0rhkJKU3WwlnRNI1B2xGvGIpfLSIBCNxXrsWWZ90T
c1MH8Y2ob5W9v9xSEnAjRCVDpOgQpVz2o50e1ZNaIlhfRfF88Uztz6rSG6nPz778
ftIisbTqzQX62YDGPiqcXJ54gVcELODD58feNDSt/SPsnfzcDBzHAANj4GjiOwJY
7ZSzMTOii8yXwT0dLyk2h7kmgd33U9EP33JqGalQYJHdv3xlprB1MIfklPwDnbQQ
Cb6nY/GTPPKqP0GEntXWE++4miJ7uR6VpqH3OY6LEpmHQk1l2C50oiwM0F0+Gnu3
C0V3b0duPu1M22vKDJ2QllUk4bVZQI9/8g/hjkg4rxcEn8PNeX1UPLfIqHtl74EX
B4+ZNXumwKWowMrhDTfPxUT9ANAGjAt0UnZAF7bRk1c49wVXAXVcx6NdukUNjCtQ
gIzq3XgSeXobk4wTKAa1FGIQp3sFoQOXUVLPgOTFKPPz9zbDAnOOWLQ4spb4AnFB
uxsybGNRz/zyYCpGupfP8aM/WMoEXTxPeTxv4wK64C+2+JzNNnhn8zx7hS2a8s8I
BmsTkZ5Ea8QLUC8LjpBpC5kSvE24CScHbbbKovr6yfiGUKAU7ZiVHIyayvn8txfG
5BDAY9G3WUIWO0FgjNDSh3CVb1mYxmT7ZrxBEBX4LRM0xBSdK2xq4rqH3jfnVBZZ
M9ejj+on4lfWSYPrPqQAn/AntoRtXx8JbuBQNLtaRIUHCO4hShQjBfCDjAdazE+f
7utveYSzQccp52NMWsbm9hJPT2Y+Z6Q+lnQbKMEzDkHTN6u4WfgZjHo9zdFWr6ss
s2hwv7EdxmZksZI3WE5/lue1mDJoRLSSxEqfBi4RLSV7P9MUZ085Lj2sDIPW8u8P
MkIgMMlPkYtvk4NokaUtdqgXSCfHUHmkrRzdrygcLxDR2ASEpKtEQJfWloSyQtN9
A7su4PH8eoDstXODnpMOO+ZBaoyXwIIK01V7S7IkghVXUH9oQ5FvbLz0dX1LhJNc
+XESohrN98JxeTd92FkfDxETSmmuMxSRqyvnaAR/0xeCEanLl5LXa4oGVLNpuyeW
LYu+o1COearjyTElA/g6Vc/F10g8wyaCjtmrWGIOjqcIi8EHqNbl8tBtI9coBwew
p6oe/jf+m4fZanZLmEe7M26kmu16k9JdBVjrMKWqjQNHdD0CwFGfjFO0LTzT0h6N
1/DjQBYMzacthTnzsl84oQHJ1QVOXrV9eu4h2CFWfZlqSOYCNVjd5Vu57y7z8XBg
p1zimxOQXUBTOaUEkmUOdHghYUmK5SjODjEkjCqTbroLZ7EG8teZY/Wid2d1eXpp
OReQrciCMdUmWtEBiCWfntBk8arOx92iagvNJmVA1DiasvgzpIaAxelGK7DN5NR5
WaPHa2izqWuVs4SQGRZ0PLwBkRLUT2mG+xgwkhpv6eEG4YNBM0IgstUN7av3sRiI
HKSKVinNblt4Tw7jzPlB4fyeIm2vfjQhJhcsH6vkOiSIjbMm9NWiyvgO8fiBRHX9
`protect END_PROTECTED
