`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cKi1qE+b0b4lls2+bm/FqAR5vuRmY9KKacnJK4KdID8b+X3ypgXZIXcz94/+ZnDw
3Jm63GWj+wPWb6qd2fATnHQim7EN6nZQZjUkfhiWlnWagUZFWYZE0x5av5MKgKwA
MUlfGxcbElCajOX3zfUBri/12j//VXtqqNUg2xqgfmgu8cDCgE1FC46dguMDFqBc
5/qin7XNYyl+AFkbwQWYfJzIU/qaousshEOuUq9XTxtr8pyFikbu4vRMr2OdfPyh
`protect END_PROTECTED
