`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4KjK5qsNPbtCQvJnhDIVUTgGWbHfbcec6CO5sNJK7TpZQeZKDVTCfeti3HEXBWo
dpDMmMKN40kvIQQpEnVloecHrzT6Ycub34DSyMyJptY638ZjpyrhroRoqJ5h8xd2
ZTMrxlPRCNVMO1hNbBMgSe/7tw8CFlmPPpNIzeIQmUUpVt++8njaVg3qwaCTcIxr
3PpXdxduZPg9v4gnshPAQcK5gjISJvAkVU/BC7VTuDxSpCNoxk6d4hUlXSH1Zmnr
Ymya4ReFgS3nutB6borsjCvDqWrLuE2QefSBP34tIcQ=
`protect END_PROTECTED
