`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1i18qLCbWu9kaV+LVh7YEIHf52hslR1QauZOG/mTJSsppqpSfaFuHZm1y5iSzst9
B5upHidwrzCR7BxZYcRO6+qDNTGOnT1xu5YrTBMjobf0HsjXRFYaMU7ZsX7YdK0i
XF0oW5f+SFssK5MIfBdBib97jQg/J89WGaA9O4PiV2Jg3Ydt7UdtgvLBAykZqeYm
VJfYhPVuxVsCwtwPNfDQ6hKd/vQaKZQog15bin65UtOSVuY408U0ow3s4wZtDc/t
yGVVuJHQHahm7trL53lm6YxJZD0fKRNleI8KaoeKMdg=
`protect END_PROTECTED
