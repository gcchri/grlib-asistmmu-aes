`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CbZAWE64HmoW0tyS/Wc0bzG4LpVKjP1uNE0+VK8WbR7foNCSpa4wF9HlD2zGOpcP
UZbUfqQ3ackr0tZthYO96DwPCEpQMXQWlK3J/GhyaYkJpeU6y5n9aqtbTY3TW5hy
oz+6WkHE6rhV499gLZ5SCu6tHFYZTl37SzTu82OUv5bf1+4VUEqpEvmv0yDnw9Zt
1DUFuHBJ+dVuUE0R3SQnisTGBkd1LhJn9e9Uk1/BAi+1U9Tgh8uPnkCyWG3U+W51
CrvYMZ6yD8WbnBaGjxWY1uEf/+Zs3K+l57SHAaGDtIPLZp0YSoCPKXMLJ1beTtOA
vptobDHPGBed1oni6YeDaF6KF3v+zbXBgxMko1piEWIYlbjeFY9tlpspUyMmdwaa
FtAyy0T9mE3yAqE1WvrKHD2dzucirng0HxeZeNzf+ro=
`protect END_PROTECTED
