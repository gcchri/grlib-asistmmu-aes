`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M4AYy6dxKlwTLlKi164/n2IMt7tVf1TjwMt2ZnB90Sz7Huxg1VqFwsOPsSTVjPE
YjiW691srQClanSH6qswZ4lYmhOPOckixfd4BrNk3DkvEoma5DPdne2ZhWTVhC26
H84egG8jYZG7Q5pnx+2nd9IoM3H/KceFMxMNZXV38wFZTaDHhoJmjokbMho50gSF
HDk8mwsYN4O5yjp06vkYYGtlv+P321Hiazd6Lme7OCiabJmCDbgFd9anniveXmCU
TD2ClPpSDtjkmQEIJzUvpuxMJWZpMz602+7vxPOesooI1hmLetzRO6xC9LH0ZhiB
Vk4C6S+4sXWuEBX8pqT3ORUEecKEnidizADkJmH0Vk7VcwuQ5IcZTzxBNySbwgLX
OapB/O0631b9bWsEm9+pPh7CwfaWeFyGiYAMO0wF+cJOtD0L2tA92srfzDAKg8bw
seLnKxoQ5DujJLlfl8Ev2aGzSq/kyPfSnflaiLa+/LAmhHOGLs33sy9caMkJYLjf
SU/p6i77ayqYUR7zkNUwsMZM9qBjrYpg5alzyhAd5Y0w+xwSsBwrJyQRU1/zY2va
2+qhibosrzi8P+TAcxJpGMOImYg0FziudSNrZy3RY0eg7uZhH+cR+FQQxs8RONAp
33VppgWPuQ9H7XXG/GZ1WYVRreOlytKs8a6QY7KPjSmrtwxe3tBDUDHP/RourLo7
VXDcNiCbUi83mzaW5vBs456vsGeJmjbO0XHJPFJXwRV2VSvubLauqgsKkqNgwfxt
Epy6WzHityv4tu3128SLMDBdA0GyI6SHjR3Jc5EhaVM12tQy4PuYR7g0wYCC9Exc
cBebVb3xGKNYxRp6xFrI6SYuK3/bT3MI+cJfQf3jMdLgqy6HLbKT053ZYnT2zD+E
qSnjfcrH0YL9En6oZnatayiTP8LOlQnvaZqa9H5yMDRGY7xWnJGzVPbZ/E2DpcKb
dQ38Hs4wY0OSgsWCgPwKqEiqrs/BXLZinprwy/LCJxnSChLsBhm+06ZqRMtpVwmc
5aHayjsScDASQs9YkSuvDFIEK8KZpy2Hq9FK1dB70cREYsYgTN+7gWjpaOoZFgLf
09+XT8/lQEEtFFQIZZRwR73I+Iwi2l8Ori4jmGOKekvYekCx78r5+G4yCM1p7d3I
vOs1NIA/Sq6Ta1k0ojgnxAz2stGMV3yXVSir61Gopzsxaaf1MlQzMRJETMZL7lHr
`protect END_PROTECTED
