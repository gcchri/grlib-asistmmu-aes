`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdirXrWg+3TCoGD9i+Mc/Xpnu8Wm3U1al41Q3p8SzV/27w1yki3MZMT8Sz4zQESB
dFOWUoapAtL2NZTBXPhbwxti3maSjVQWNnXq9FMFVp6rUjkhZ7AjmT6sDihZ8M3/
90pNf5AQDhasp9FxMBkq2LK8fM76p1BFARJs3JNUl0QdYNJserG72P7AzED89Fvk
cPpM+rH/t0XisCkLFKpwyLCaFHgCz7dKz1kz6xyrG7jeehNldjr7TJkoYJAySlOs
BaS/qYZHRR4z2VoFKyUK51gEGWT/Y3FOF0PnfM16L5cnR3gpSI2+ZS7DMJYhKPvR
qQhfs+oLlC6yc9I+8F2tcXloyURcG1jNeP1a2TfX24DFP0tIrIYnEiul3jnxNEry
MAlw585k9XPXvu4BPB8jllur4CEJXTY5xqWdk7Ii0q2HvugBqyGEk5+eH4A+Z8i6
pQba0ATOZDRJcRY97UceaONW/LhvooKuZFO94EeNjMId9L/QPYabFxgzXTDQQL4d
+7lozSFNkGubATq9emgAHcvAxDi+4jQ+sIjSoRoa0QIxhQsIYXSYsNWiJK0R1m/5
mRPd/nmwKeOwUf6E1+FbE51PVm+R9vVgM72h+yBkrcN2WHdwxFcoCRK7v1bIJpCA
3uGyoSLaRLYkem+2WzHmNJ/PRdl8906Bayx6bqXhECm29/qv0LcZiimMpYhOsSKo
NIk13A2hfKK6VzRgVSaf5peUwIGEw2gGQm1OBOyrb2UM1MjmGIc5ajoc5ssWnVnk
dE7a+HJ0v3+DENJ7xFYBILpZNaXLe8o6/KcAA7J9g2zIrbNaLHC0DYjSaKd6tQTp
PfDjeGnE+P2ljhc5sQ4ueotjWuvt03HkRu4zD0QFe2p2/iOc63akIlpCEVsXkGaB
CE/CEpdHxudQULSCvKfTrkYxzr2/8BSYe6oqy/HnuQzRBw7N/D2svaT+4R6Ys/ZF
6MEEY/9Q/n61SrgMEoxa6mAYmFWNH7JJscF1Tdk1W7c2YOFHpDLK9jp5zavGYk7S
kB5P7sX/cU+Q/cbsL2fHaBEVsJlqP347V1NKJyrVztwMJxxw80a56PoEYepb/j8L
eOxg5eby4bztEOT1rSizWHOu0nHpxKw9O1mGR2n+ECeI9yimI4hndg/YrsA4DxpT
kopt4csOPjKgyvNb99oMUMOFUzEMNSrtyF3NW0Q20LF3DpYphaKW1yaK0y1GM+v1
x/sLcvNRVNxMcXikywlBuuCo+MpgcAwAFD22ZKucZeIPsnMP9tHt35ZAt2EcmWtF
VjKnyBPGUHsnDEaCz/sctHJ57LMYV3VR+lnI+Y6wmIYTDduVVE5hmqrFYQwmAQSv
PUIcr6AUfxOElx1ks2b99HR1KAGyx7e26xyGr7IIsXaEGdjbGBfbVs0usE14ueQL
SWZZv+A0P22r/RaaZ8HF8+zXB3yevw58zwzi2nDXczyStCfnwzEK95NHQD4J0Yu6
4al7XoHX2Nm6nNg8cZXmYKhIz/WdmJBB7wlgZ1p6u3Yb6W6jUdB/UFtwWdUfVa+a
Xz8E0JEfnvQl8Dc6erNFu2lO/hJ32xn0Vhu0lgmCm7d5OOxuZmZFGyQbOem3GvA7
OoGt0aTZ5ya+WcOFgqPAP2ggq8c8fKDgqge/DP+FQVOQKvsAS/RXaDt1kgghR436
lk4pkqgFeK/HxMFPZ8bKqSlIEpmSNI0IK7rkYDl8AU2rmA8ykS5pCFSCGhTWfVnD
QCQPhbuF+Jer5uyLmJOX3ozo9QYb95K3Gmda+E36UuOB7tiuChtfhu4KRVqT9NjW
huXqIGjRJy4mtZZzgdYDJqCeneq5Z1260DqTGtFkFxl2POLU8jwRJH9ckvlcDZd7
01I3e8LFt8uzY3y27A7mYcf6ys8CahJ8KCarKT5TNdYyYv9eaqZxkDb3bwBcPNsJ
t/MruyzeJDvyyUFJjuOfrbSLjy1qmY20bKvgHjljidLHI50PHgNQPccJKobfmOBb
vFW/PfHkBrCKrkOfFuCq4qW7R+2jZwCgGuieAbqVDfGocTRsIf0uoYweYYQ+Bb1+
nzbyVyDjNqXyTw+5DuuPS24ON8Kto1IpJu7mOT/ixGOCoowwYsxVI0sLkdC2qVyn
Ni0KYG36n0ODdsQ8xFokpt1M0jlm+/CfyQfSgLp7TsItktrVbfjcLQEfrSJGko1G
25Zbg2xrTQeENqqMzfWiQr1JssqHeKs1SHBuhX9+aD4HjLSWLV4yCo6oONbJGyeW
1eEA6G/mp1J9cHdSQHizi4hdJqWRYI2quMEDOFC+xegTh3ZylJio9/ZUOV6fGv5a
c6bLZg62LCxUzFCN0f3NVTpX6oZKpT3iyaqgU7JlcjgEYPdnSrIjij6hYzz4ctfP
rBem5T+s/D52q9Ws/p4gj0ixSrgGQN330ECCFGTjFagIZK6T5ajmoD+6z30iUzlJ
c89ns64akLDbHVD1vc6VD1lB5DSA7EDQHb1JUb0P/8McTuIGz2qkfW9yLafCFJ+u
AjdEDgRp+ptW08hr7PadeoyV6CkST9uPas+1jJPSdNtpKEbjFmFKru5awqPpVjT6
Nhv234LTdovFFpRqvbokgRuYGHdbCxL42GY0PeiaWNC6gerXjSHzh6yJeFJTKodA
xLwW6BdRrSngoHlKmvTggXIc/5RbH4bCdp/HSCBJLr3AOt0HwmPQlsuEObALAuRm
YOWgH+ubEZxz1J5t7WL7eLWP5kDNEJmgtpEK71o3D5A=
`protect END_PROTECTED
