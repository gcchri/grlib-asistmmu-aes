`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JIZAM/0/WDUVUEBwMHuIey/k9B0ZbiwpERNYyIU6UDGXdd0hDVvjTWbTqH2HCDK
pRHsDo1s6BOG0FeRyafvWxFlDU4JkC0m/nipldXKdLEmUoSj/fODyn7+W2FeC3wL
pb0ZRpcVtvNDaDYTU07Sw6Gppy/ulVEiDO7P2fBBOwT2s5oKY0WafrqTw9FrT3Mu
zzeoO7eQQ3GmL88lX5rWxnsvHMYMhr8pFSBGhHpziiHCGScC0dteqqVdcXFAPyeg
p9BTs74+ah0yaN++NoOLGUIIohqAOXTDdqeQ6zN8ADcW9DHbLX18zZ1Ok0xDpsdp
Cw0UphVXoGaQKXpOd1kJ7nJA98ycDE6nBpEHqDwxHnf2BKjACy0bPr0+/nCudUnt
TsVWb+LyOf83XcVu8X5cPfxLW4kUTa1x78Q3j4uCWElRXWCJetP2YEz/1BK9AitK
2baRIGr4VpFE1tFmAwEaLWiFNQ1H7G1FInoMxE5TfDtz8aw9aK7WuE7wTyZP84Gv
OPf2UneGQq62eVslPwwJB4WJI/5gjW1jwQ2CZR3dJm/CyiTABgIfSPsVxt2/7xql
QEiVezcV+YTvSUBX6U6CXsRFZQQMpA7NQOlEW0dU2QLK1RTvLs9JYD633/p0WJNe
9hWjmQj4RmKHhoyiBT2It77uCj4XoAOfyQRf3k1RJqGnrNKOqOYHutGCy1w/e7Pt
XFzVfexEX7ePMBgHrF/0Zez23+PZAKYAXUKVpsH4Xns=
`protect END_PROTECTED
