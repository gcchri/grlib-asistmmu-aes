`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MX9hooLJoJM/vxbR8jHwq14krb4CdxoTyP/D1Oflxu1JFKkUXloCnKEFNhMHC4aS
4ro/ZRxFaUsl52lzgyLZmPDl88ba4C5bBjav/LdOaYGMtwcEyReA88uw5Bt26Zkp
pWzJ4q/OKS7YpW+jIF0slGjbA80mO8M5a/VN5h8aCOOisxrxx1AsQblZU5HHVv+T
sHEJe/vcB7XiUuAko+vJOMZl/Q28K1AHL2/G1mGNhaRZH8OkaCApFBaBPaiqQCGI
sBekGMJqGm6bNQwaZbjEJbidkrD7/n9kGElCGjaby7/7FQBGPhkFqltk5UiZd/UL
oj/G4x8Z4mahlrPuSNKPgjMtdOdmPpJJa9pulLxi2obnz5T75+7PGIEFG1N4QoxZ
pQ34IJrc/vli8g3KDkUjO3PiT2v6UETgdpS1fJw7hWZrXeP30w/RWsiepx9LPXBw
uoEC7koaF5MQf2yVgDmHC+YEMJz0shcJWA8L5uvLo8eR5ClWTiwe2DCPFqMsKw4/
DWvwuINPplMh1okqgdU8AlI2/efh9YC6YHPejLl5tOl1rEtg4PZwY/DYc5dJFmzE
/QbM1tlYZLIp0ibHzezSa6rNZ59jNUglrqWROqbIz4vR3/RWOnhbd6yBKP89M5iq
HqsEl7nFBfIbQlNJJXl0R5IfMMzUBtLmTKpo3Dsn3RqqKqj0DsjWsxMGS8KARNQK
SZFeekTToM3MKNtj5ahPDa0qo6Djthh0EHi7YmNGC1YGJxiu6UERwVsKXwt/8DTH
7R80FJBlXbdZXqwQb+igS9ctFa4xEKmW8e57F6iPoMj7UAXoOX0EkrUXjgliMovA
0zEvf2W3pGIlVCK6ZdRR2gQCCXneajMu2CpGq6f2Yngisde2gVyptudMDYfRGkr6
2zrjKdMIZG4r13BYgiwNEMo/Z6dyHtANqjAO6g+g7f3tQZEpD8vKn2ecuS0ZrQ8l
gU6yc0S343M9EmycqD5Pra4N/UAwUnH1yX74pwRedBitEBZ48AoTkxJpZ29WCPgc
dNg3TzkiiznWtX5WEPvUQ4ZvGmjoXYApQxNj77kCMsBEl3TBwV81sAvs3OlV8JrJ
AJ+KbMcOffOS64MJDeUqa88HfZhA/hd6KSYBhIMAI2A4Hm2Iu6dZOyooGchYVM31
HJIHcTAlW9Q5lsEtHlfbIdoURUMVU2xhMhcVSNXl7w2KDLSGSIy4skM1TZdJMpMw
yQWAxYx9jm7pM+RsJaHZELYJHYSmf3bGkYlGr6o2aHcNF2b8pQb17ihAZOrserKk
FGvOl1E0QalDvVZS18KRje9RGIDek3ExcTCST40x0If3eAkoNF8G4af6f5Rih3Oy
YzoQsuxpkAbVrLZxjd7tL+iRUlc7lwzpd/y+hotiZtCfSYMOu/RxwHx0OQBODpoK
kX9E7QJX94LS4nG37DrprO0MFNFHFZeiGXNCujn+1ynh1D+8F6epYCdIUBJhC3W1
HuH+j/EvgBoPYm1CoUmkifrpRtMr/NhMBRRcvFdjHSVlMh+F8tUOByolAGeJSNMl
HSMOtwTjhVuhTK+HxEy7C2oVyAB5RlAuPoAthyX4wHfTyLSSoBAgpvEGqnj/cU3I
eChj9r7TiUtviKx8vLPrfKi//vVuwpQ+C2kNzHPqYQlguLynTVaGpi8rb9q+qR26
Fxv52Rahqa9xX04SahHDe2C/I1ZLAQYcVxmL6LM7FLJtG5SJ0YNVf8zRo/Xmznvc
rjhCjGmHSnKDdEp790NaYw/Eu4NSd4+J8dkKtD6JJLzcSDWmneF6G0wDfpat4+TB
5eqnzH9xavxNT1ZXofIq3bJ5Cd8hxJEX4+qCtAsp+2FxDfTDYKyIbGJ4JNIT0NOM
RAQnvzyHBIWwsNXya8H1vWq+3AcYZ+FBUWCAIxYGKSxEYUDG9l8VizKhwUiYGk+h
`protect END_PROTECTED
