`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aCtUcBCpBYlS2U2Ihbi6iU4LBpZwqO9BuoiCdt6W7k5oyEXLvHeq4MtzRD7+tyWu
OUvny6+CQjrjS6MkRFvspSt0Xwxrbs1L+PwAxGCjB1zepTmUR6GSQhMw7+eSBuT2
1AiZHzYCRjp8Tx3CMZPEhQ2gB4NKJ9ikVMxlzxL9OwLxmvgTHcDqkBxQu9IbWxR2
Me08zMombZcs6BhDJQQMljWilClNT5WYoKZG9cEJRxf4Sc3lMsQui+4Yd/NT2jfW
KQh7yGzf+EpJo0mXYaiSnQ==
`protect END_PROTECTED
