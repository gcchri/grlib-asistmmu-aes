`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N/x7m0q5VuEj6r4gkBPSjQFQSqFdSbrz6U33x6KH/aPDsaPm+UPtjmAejC2PNHnj
MmcoO0iuDRFA1cvbcVcWcz9g7aTbIWC2dXYAne7WTsTCIYJ2iXuH3G5tXgiTPKMN
uwidBqegV6AHSVlJWE6UJwE9I/J2I64DnS+y4DtDCbLAJdVDZVealuuH+M2NNIy+
aMPCJfarD6eI/sVlGVJZjvmnZuL55K751Z/eXtLxARf6aqtX2YnmaaChC2ZdeiK1
y1SEdH8uciChzrHvBJzXGZ7Edb6vCn+uhKDuC9ImGgqa1CT9teJ005bfDHKoUZDg
PeaT8i1M6058feJhiyUiQ2JmL9jsmAkQa5c0JLE51udwPgNjlGaZ8+BoTh4d7ZS/
SRCvph35B3Ls7EayLnSg8qpiB+LBMDtd6Qlzes3Stxe6njcueCgTmyOFAXqNjmTd
csR+gdsfDqaMvmQl2bbGqbYJuCvjsFljQvaKp0GsUK1JgNG8C7fMBwgis733Fot9
Z9zW9oH6scNJ8kwLeBh8ck3TVn1kuH0OWAmkDH1oUk9N3PEJsKyp9A2sGmsM22Ac
eOvzHeyds49+5+OaPSH9GPo5/4S4wPYmEBBuShvZQHk1AbV8PC5s7Guj50sRPFkf
jY64pBWYoZIhvI6sMp2A/TzprRTcKz/WynUePVN4y3uR9SjA0RLnTJhNTQT9KxKS
5S201A1YAPzQnNLz4kazHNbwPP+Rn/iF4XyAKa+DMjRGn5fzf2t/SXNImC+AKWHP
yn5Hn/Bo0zT7iotayhB0ByPvoLRibaOWyVl5+6optPUOAaY42ZdmwP29zft+4ofJ
Qt8d8PPu7WosA+7LBr5L8IL6EKY7KX4jGLizZYwu6X9P/E94GALK/ff9egwBciIk
t4aVI0rH2fWUOQnOZmoEhohL7HLDOJuwEzTN579YvGK78RL1zADXa0w0IZfSqMsE
LSV3Boru8HZDji5Hx5pe56B3fp5bRtmzp6HK2BmfRG52SxWvYsmS/5arB8FVtg+J
1CvoULLUfUOitUqrvRSQoLEzDTGObICVZGTBbgzXpOUO6Scb7BOBhwUuQSadBDr3
e/l5mhvjS6naKXG8kC52hUBLNwPbI0Z0fI/ls+i+eRWddrqLUNcyypCshyBGH0IG
sunims/fBVl1hVTMycN5rh1qfLUjduapdCouKVnvdmYDF3TjNQsVrqhpMoRQlVXw
IpPxQIWXCHK6nTIqCIN5+z57Q5Iq2GoX0LwoC+F2lORbYhrRRlcJ7mz7q/SLNpw2
tDsV6UvQK286gw6FQUcjzyJyLfv8YXpf+1mB0+Gio3545SvtL7J6kPeZWEBiTkqv
NiYKVSiccRTVqbLEhBbhJjULSSZSgALLqy4NLecS1LawseWso2vG5SIRomD2YhD2
CtidKgPdH39aYCiFnbiUCIHm+EFxU9leqGwS5atjbkALDyf7hUpjgO8yLLp2zH5C
SWhsQUI/eMKnShR/vPw+XPlaMJaxyDdvEGATz+hbXlYI2aI+wUzg+Xxoc8SR3PoC
wctms+2xA6u+PKRXHWJVDIwX1mCMBmZVqjMmrztTGSUEs0uwtVcfIYHHKoVi+YQc
Xb4BwdSzXQ9lBOj9XOjAuhqT5teOE6j+FYmnJ3qEnrp7lJfoIu1ORb8kqNBovqLr
rBJLhwcu/4702bSTr9BoXuMsUUaQttJoga4ZAo35R+mi5HMPcN/GAcK88uf3rcEL
Qgpn/zKMa88rv4pLrEw4H8djrgZ4n/qYvNYGlFcRJZ5YNjHkkd0DUOdn4DdrTAW5
UKhDCUIG2ZEwxF1cPt/7edkcA3zELoS7nW8uFGMYt6OmVuUMpBLek0Q91xG9mCt2
aQkyLKN0RDdzAvL4sBO0/4q/GrEvW6t+6gzhH2G3a9VJcgwNJAilw0jDxpKvYr09
GUxubLhQXMmu/Rdr/00+nE8Anxgr0Ubl1w1IIm3lQOuTECLTu3I5Mk96v91+uuo7
XYStbGkKjObL384LH9+3KbRsfEPRlPoITtzzvEwTdS4wkBAArWyZoLub3ATqchcp
eUTWuQBPqLGtVEbaIYJW9nTKX7lO4T6G8yEdMsApRRJjG4OLrR+YLNsMkiBYAi08
tG4OhJQ3fgYP4s4hf1Q3r2QpoiDijbuKG7K+JGq74QqzoKP8dyY0QNtp4MRsbVlA
hRCrZa/Nx1SzcAdfPmIy1edfGT78wLSQuupyXgKaIezt6dzU31qqHzD0q3r2prn/
JQEvBDkOjADPbS46ZaaZn7lbsHtJ/gJAogoROi/rIDNIeJ7lLlSmgw7S+BIh6ByW
ZvgXG3pbvVjhbSQUzuDMNa+VIdFMUQIxaTTsh+WkWSreINSxGgKRckVBLBwxIckG
Otz6uv7b1ngOMdDhOr9ZPNYY4OVOsIrmXZCabUJszDfoUf5X1UuTMXSChI/nKDkw
AEMk+a657S955j724zpvowzTA/oZ6+MVv6+gnI/QazVyZ6PfPkzJLji1q4U0vWwS
2HomX7VPe+icGOy4vI8VZY+AHygo75SHnKx0mgZbuoXioi8bFYmM9DWH+5mnOTwk
Sflr/Ugf6PM+cQsv38NDDLUTaLwLnSnyrXu8qY8rMkxX+af5cmTyt8AwESrOotiC
1r1LBS5/gQQuCh3dv6mdXb3RQoVcRna6d3WySojXrLsiDeueH1qKnbIvw4jat4kA
s0Hurwve7N0ih2DU7ROkx/QhEYj5B71v3MUzWXErK8M+5Nd6j9+LJq2cTU1gxOM2
5oEU88nu656jifOHh80Sw0kKpv501+3in3MBbE/uRCKWskw335EbPpD6ldZ9NfXy
6D7Ex2PgD/TiaYvzPQjYYnFu8fr7Rdh8xYg7UbqL1QuQZv01TSdIFuOL60XHXEPm
wWPSWJzGe5mGclxQ+eeHJ4c2mL4ZfDNVTFYmpKqvZmT8ueN+kb0q6DAg48fqbecE
x2OS2lINY0FexPB2SiN5yuHlgkQtpt7IlUFRvUAp8eGPz/R4NadkuJWGRRnWHMIP
p6Q5D2Z0GlZdB+HgOQHFoVhUKCBSQwhof8iJu/nKIgEOJYwDhXGjOdqnpfkfFkqW
rlt1dSWBGemlTQwC9LNwBxAGJKCWoV9CGIYNdePnSyCR3dnxBx+hWsCrEsrADizq
Ph15bgblLbhsMKiyFXcA+Ge98UcV8LaGRc5Q1kydM0ZC1NpXlQzIBA8mvNEZfma8
VYf0vRefvGTjBuvXJTiED+XskJ/DpmK59C9ol8Px+sc37CsR6vPiu93FELYWqxGf
Z9ymVO1SQVyCI9KDn/NGuLxIjPIna9MNhAVA6bGoF6cE3IR214qOljTVSrhsqn+2
q4NTlFosaB43ZD7p6iiviG5aJfo4cBtmYO+t1Xlb/t0XFfnEHK2dYwIQhDrNLHwV
FtOHu/DJy+tgMSch5vtd7EByoxvX5vvXPxhFjTMauEGpwYuZVnGibLFtS/MfnjDr
yA/9u9Dth5uK86TWjhT+ZH9dfCxG0sNCU/2W1t3lxvCAu3KDqLMpD7aY1T4kEx3b
YgA5/9gozVUZraBAt+uUBFNbVFd5LyxyoxhDbXAYjCft6PcVCOLv/8Dl+13XmO/X
gbay0W5OGIEPTBsK3qOL6IlLhXL8bpZrdP4NPLa2FkitjOaZuTxXCJBMpdIh+tfZ
kz56bdir2CnaTSMV6hm4kRl6B6cmEWrlVWdvFYIgAq4mveXVfEU9y91ZEUEjeGaL
BpcouGNMoSKKZkBHlTCKm45GEkRl52P7yEirs2ljBwtNxngLQV/axA3S+JmnDUWC
pVKG4DfnkkGJZcGvLthqseJBraggbISK0lS5MrpgUUKeA/j74UmVuPhopJjkTh6C
7cKcRF/XqxCwl334jWqyaS8ZrQEc9S043VqWJrntXmkE8j//N45zeAtvBcEVgqaW
/eomYIpHrEV5u3cC8rz+paue2BZEvdAaOYgrjwkD2SMxucXzNGObt+3Z5ekSjMib
A382ZkWSe2fFhFF7LylFztLwiuNqiVh856zi24bHveVRCFSFbJL0MGVCymC7r2v5
Q314NQWGOH4CyLkpaQoKcBZRUttOhpw10/86RtddQDEvc+8fnrj1R4CWLIt1+Sgh
uEkEgBnnunKQjx/rXE6Uz5LIgZWMrZe2tJ6G4B6IGWXaMfH9I3TxmMaHMmAUK4nd
kfMKFNf1GxydqOLGQnZvQ9gDOtuR4TWQrjLzZ5fdmAZjkujt+TMHOOQYhGq2xGDw
IqzHDHdCcMiAw/3hCiL+wNzaRk6/uIcGp0MIdAZk6wS+soWUszK+aEwKU0wOU02Z
PA5u+BUpc5Qiy7QmApJiiTEp23/KNP+pGo7lpQmaoatjYN/TMNinuBFVqw6WUKE0
rUE14UF4UWXoWBH4tafxRm3YJIW35P0fPkcsFdXwXbhDWqDBudhJBKNd/Col/DCl
4sOSa36K48TkM3cyIqXdRy3CpZ9l/x0YmerzOr8TVQhL0p1NglJgfB304n9Y1E81
PW0hhXFcK3mQttaaBfgerpKO0ulRMnJUFF1iMdwCieGhbrigHFGGEgI6Anb1h6Ia
u3izOfbiL/HA2Q9wlsrVdbdIlIlZxXYClaJxrtiiy7SAQKUIDH4zHrLHAFtVc1/c
I94PjyqjnEMCmASTdZvsaHMmTQ4ElZIT63OZIpnjITMBh9jvCHQGkUA49bvky/Do
dGvBNaBPLNGlRCwj3fO1ntadTCBTjBeJZyAu3aANsfEGeqA06QW2SqxQSvwDnkjb
9vu5pbyCf6OKhUhZdDHAdY0hCzib4m2+C6VpJHoAQxKhbENQYjzMGUaEvEg5FwY/
PB0UiInjCYThNyoIXahvH14op8PdTXNFsrkp1yRm6U4kRTvqQ/VEf3yXLZVgqxWu
234G74iEwAGH61ha+SxB8Ar5lLm+ClILHJ/wlqMAGDBS95V5iVhXBItxBXd3Qr6d
1s+k4Ahp0m5c1RO4znNh2ar2wqmflqsDoTQbgkVpKriw/SW7D3hiSQzS+7FEnqPi
x7pDpeXhP2akzv1oVtEJC3g+tXPE0k85NjzohzagnP5H0KeTYiCOXSbbRHplL6TL
ieEFR2S6enAtHuAH/IlHXx3fyVB8wLQsNsmK8rSRUIYoYU0kxZYjPsfLMXTGrSSt
fw7nHScxt29EuL+V5u/wBxj9KHZXsmeHuomaO1ki2dIsMBfaqYOOJpHrVwyixdaW
SHLeTDPuZ26FNVS5IA4T82tqkvnrkkg1FbOuVd0nXoEobn0b96L/cesGYBuOj6ZZ
i31w0TroeCnhB8y0JC16rTwHDe7D9t5YdE3zLvGLNjW+cK+BBKOfjxIUEMfyCCda
FDEBKjkpZJGW81lHxDum8LtwGVEbxt1DQ5Iy4cFNpoi4Td4bgKf2DcjPLU+HNMIL
LbKmpKS/8BjhQltyYuMHErbDqxvvPJNRdd0b1lCu5kBP+PvFLS43ybCPNHIfoaoW
RXEaajNHmOyfMiaGrYWsh8OrbUt7v9OJ4xEAku+DsNilj++WcuvDsQ9RMcW3crDv
G6dRKhE/uQFKnDtskir5j/doPiAQnmI+K1o3Jki9wtmajAIZmU3J1I6Lkjps1YQz
m17o/8j7CcEU6SZ1vzL8nH5JnW1JYuSpT2dCXmnpZlKlUwbffAMxjhQXVzVXL5N7
k7YJbYwS4Aa7BHcirwPiUHXTpw5yh8RhG0+9IKShUs9YAND7AgQjY43bRxQ9L+qj
8Od7oIqFQVfZUvTZYV9g5NK9pU5Bj6OqgJ26PfAWgRxxeCFlHPLxWQH/TlsyEcwJ
PXB4rkhR0ZJRdjip84EefBUAp7viUKcSsFge7/YD0SmQslZinykjJDrWv/QNtxUp
RHt9Nbs60XbCRaUP5mzquk2W47cm/6J5q+/iD6du+te4Icl7tY2oAfAEayegzDgz
HRJEPJFbjCiWcvIFFIADkosF3fNbCSO9yO/ZeykkJibHi6Gzo1LUZQSelE7dHkyE
C9lNgTwqi67uhHHn298LibIlAZ/x9pNCNqcX01oXx+oIS2vuGruJoU6WIL0cG/2n
HWXFjnDgOXhPdgaleq6vw+eG2p4F2Fkt5JEEVxUbwPFuky5qkf9Sxa6jpbwhWDfL
GGJt/DfNjz5Nl/wiJlr/nCiquJ3O0NbXAuTg+wj3WbDB/hUZSo4Tt1r3hHC7Ya2X
x0kUtnpU92pC5Vsh6C+gNZO5OFcv4S6P9ax9LUkpkmApkonbhD+2yFK2nCtu6rYG
cbzgV4wCdhIy6b6pKztZCZrtO0mDXHJAOsGbGiT0dDEZ6KSPacqR3yKOXesdPx/M
1/K5ZQDleDMFqIXhHjTxOJyTomH6+NZoVe3/GWkAG1wIc/455uB9dxnQgthUzCoa
gbaZFkMG2/3vyZs7kgjxAHtmzNwDDEcZPky0qyxAJaRYDcJy4caAwI5MY4zG6yk3
YHUxa6F3oetn0qGMr48hogHEdyPXHKlZi6JTnSRQhZvAqEeIU3kzxajW13WOuIkh
LIVvhtw/A6/OLvPf8OGbdZcQd/4EWUOQP4IQt0aSBSQYYEGw53OHGPEDEPjc5PZn
Nvm0gTE2gQ3r7rh+bb/w2KzmaJ7kuAvoP8NAHkHueX3mufG499b29/OF6Yt7kP7M
thgvAe2zQlhSj5MmrmZ0lx6f6syiHl8tdnEg++tWq5T8u5SCoxuyUQbMQHql/Iyx
7uAnIo2O+aIHOgtkH+Q2HPZI1lZ2bH1HMSngXDe799dH4PERUtiU5yPtiqzeGWOf
+X/lIIr5RiPkOmaz2N2e2y2ryJhNrgHizHWizNnVSkji/O+T0yyFRcoEWx6HsHne
exYTw6fp8V1iqh3K4XfA5xs+C0GCbooKG6TWf/eo5HgYuTuC1u834rx30fa8ri+e
H5s+vFHtEjiTCl47TyN83P9nEfsFqMBkK5POWBjKx/urfCXgtR5UFV9hAO7gTTZP
erOLi/zPk8PvRohWBzZb6C1PlpVGTJ+kIeiOoDiM5IxnqFB0K7/5Y/NZOwzestsK
0Q4z0AglP+Lw6yFI9VPtJBrPTpBww0n/ZzkvhgQ/lTI2bfc7JJHEPHQbyaSFy8k0
eORMLuVzP4pZAvEYB701MY7XGhzGfpislQK3mL/HWbBz+GbRGTYIxLtaF1TZ41qa
jEG4Tepxnu4WpQ2ck8cVT5gJm7DUytYdTW17oC0jLhcqcuJ5xmG8bkw7Gkcljb4e
39NLrhBaw7ugGrMmdinIs2tr59glLoS3VIJVXFaG6AcrSY7CpIbKtoQgt/05UdSQ
65zMSDshSa3bZJJo2+8dKNnJd8HDhNWB1Hf2nexwJtEuAP2OOlKqqLexI23vIbHA
mp6Ek07g+VrB0X6SXDdT0HTB9eyZtXIhhsjXbUYhU1JOPo/qlIkOtfURwb1GRNTs
/RqrEZEixI+rt7azrkCBGNcNNfBhf4R2uYEgAkgsYGFjzaHArOGhKUKdZ38pCNZR
FTa9S3YIyg2nHqWA9mNZ8Z/nu7Y2h+3XpdBf2KK0cTxvlHwlkec/DqJH2kQiPXmm
qKWLlq2dS+wuSLyDDSt8e8QVqJ4t76ZNikiUxPClFxReWqEFIxT8ipgTJDHt+PbJ
bvNQT3AuZtx7KTa3k6Km+7XnWZ9dYTbzlSI3MiPVZpiPgyOkImOwMeHs9gBGa4Ev
5sobz4EwhyGYaS8RMaeFRG5g81ZLLCs0MKSMVlMlYNthC+0rVMqK1XqkjvLoarlA
n1WnbI3t9C/u/QdUVdNKXPScDb42WkqCya3cKsQh3bF/TIM/sw6+XWMLwm6UnRLZ
6Hw2KxMhs80n9X0dMbuzS1W81dNzpLUnbsYtqpRm4+W6pJ2naPU/B5O1UozhKCfu
mr7joDFm6pM1E/CFxbmJ5wtK6s5GS85bKjQogFw0D01ywbJQ12umCvmJfDJgWdx2
7/fiRnlvyBcf+hC6O4CTdYzbFebWmd5c7y7wFWTTvDclQ9fRdV/X5+mjMBXlDjIp
lN9bIaxS7QHeTlHrbY6j0+ECVKHnsj/WwQdfb+yXmKsQiYi5z3zj49AGF9ikkTb6
cLh78wfpwf1omFt6x1lMzKuP/DPQehywPqNKb5MZKhkrdKFqITWpBrJW3CwUzvGN
fz/S1+Q58chs2RFctwEViELHV6IhZ3iH9SEHifAY59avf7jRQ27F8se+QQ96R1lO
omNAwutMhjhFyNk8RzQD76e3mTiN43v8p44oMC0acCpsmU+KPwhqrdg9x8k9U6tz
i4f3pub/kKEgrf0EZ3FvPyW/AdbwnWEcLqc8IuZWR4mMxNJJYUzG9i1NshgMouwc
EHvzh3yijT/mJRQ44b9ZDa3R3eVUvl+3OkoPaVw8jVxdVhnVhKy/rq4VWyhRRcXe
Rq6VJPZQK6gO+6BUNLqx2ogQb9fA5eGb7wvyTRQugfW7//tqDTdp+M4IUD2cszVJ
w+bLyO/td7TYoSe7LOoaeUqh6JQ1vbDR0s0StbLKg2RYjxtshDo+rLwHoD5IxVc+
NtB4t+OjdY+pllee13fufclmFexKNAOqkG55kHuUfRZitztAExlRP1ixDmHOK7lO
/s9cq75qiHvK6G+TF1w5jGD/yPSE6MnyHWvW84ZmpJsj47Eg/Nn0vOr951mXCgp/
XPhh6KCpbRhggwb1Wvqg1OEphWi9zDn84ww9hWuaGJyJWfeArfskz+HP4xk2uO+d
jwwx9IsnO2LcFV9UQvjyLxY1AKAhro33vPP8qaBc2dDM37Y7IOLFvR94ITpnZYZM
LuBQB/v75RxQ+7A45sAzkCf5yciepNh6ievh99Ux6icvWQ6ZaHXkF0xvuLhln9GL
t6/nTHxwwts4DbQQHgHTkxgxRqEM6ZczDHCGImVgC6b8a08kW1BXqsOLNo7P6KMB
VIEWVzBmkKU/8Jts0onLMXhdo97uojzWgLyt2kFM5s6nM1tnTIjepgInA1AbUoty
0rMiaBiHsabuAsQmh4TyKj/V6v/tpHbWAecAlb8HAqTWl/pcQmW1nrsAZ1eYDh2O
U/vb0vEjBoi+s3s3lo8MTAce2NoVN/DDdIWCh6ZsOG/Zdi5vJrM96NuglNDMxYRy
h2Yuhg+YXt61Jfp5vfJto8KToQklpQDbMhxIV7a9Vtnq8scIxCUanc699pWDY4Xh
UsYqUNIIlJf4AW8DeKmi0GjozYSWfzeNruNL/aUBV+lAYola5mkH8Uy1/6tUnJgq
+ewTmQP6WWK4EROpKsq2lbTUVU6+5kGpLgLXXjapqA2Y4ScuHTYwTTrj3F+3XNSR
99z0yDp8TX1G5gnV467RAIGrXEACbOkuwM38hmORWl22CewsaOFGE0ENt6d/kDG6
ncCST9jYzE84N+DSKj+k3i0W9lnVSZyVb7lCAHmcBsT3sMjVMtx+eDPTc7g3t8zG
oQXmoDhGQxOU1g6cRpbm4Ar87MasC2ktAu05JLHkBgcIsXqb96SyvmBaytN6mQTo
0gMKoveFW4g/aI3flHWLhcqvk5/Tg7GEofMfWqqD5sLdOc6awZ9R01L51Svjpnml
wiDDqOLIMKvdnl5kNJq0o0UuYeWF/o+uWWhLzmLDp8s6wGjrQWnFjYbImyDB0tV1
+BBlB28MU+KPGaqcJp8GbX8Keg3/gpvZIgTTPdKPyMO2ua44Kd55jrjssZclAKME
1Z2DDbmVKtQ4PAni7AyZYFP90Kz1p+sNkLcAkZk25EcM0kLsBhno6Szu13oojek9
TvhaA4kCZfhzqiOnSmPBnkhesYCQzDCQPKIhO/r//AZYPf0GxZxzIs3KqwJw7CX3
0qgHb/BXBDW1tb/O5WTJ7WVAI2soX0l7eOBrhL+sy/P9MtEtp+TM3r9duzPAXE0e
e3IHM/RgKU+Y7YQSE/UsTL5dwwHM61IFEUgHo7e3xfp3pzK7d0Sq5zq3s3B5H9zW
GVDDDURwo+/RW5m0i37/euFQAwzTbz/LTqztClVMpWhXZG6b4+xGdXflqvcxbefX
C/BxmW8yRJI/VoZl42+B68tB4XsGq8rnvoasZeVJbyPt1m7LtKgdpyLLJumkq4U5
5hc0GFQCpoBW9KXEuIax/V87Z6z/QXxwdgqyq8NXzTt1Gc17ioLGNc0+0gplOic4
N2S77XDIWS/gyWJmOXNTytXGd/t1NTL/HyBZTPKmbRUUD/xCkgMoMtOY2eaySv8e
GXLOhgybojSEIiaeyVLRD4/whpkrLidlX+Ksl9v5FQl4S/bpZt3Qr0mh8MFglR7Y
nqrGtYhRA1Q+R7flzYEDsHCCt+f5gdeIAhtzPXD5Bq90lj11i8BHmGuaJUuGmyGw
/tUo44Fi8ALR6hBKhW20DsAGMM/L3Re9Vu/X76B8NfIvw149JDzABkiscTXZq8kj
E9h5XFKQOTdHOShtRiIwcDZlD1tkgLw2oEJRIiDjf/ETUEj5SsRJCKbVG5pv43fu
fyEc7+0jIugpZLKkmEiYfnNtvY2ZmKYyIP1NNojDM+UM7C7caY6uC6Iw+XHnfaGY
8VNCgybDK4LlXSIin7Y40JoLWZq6EEqk8fQPH1QavnwP2BUGzrck/odbx63BBgli
cKlu6GUjqkfpBrrVzTlp7fH73T0v0ie1QZfyF33/aTa+cjAbbyUDDK5cVhdiVDmQ
1WmY3NI6YyDdSsGeb627gJN2Zy2uA9qq8IMLdlxwadqGzq80eu26HVZ+LqCSB8Ni
4jwF8mcbb1qytDtycHhlNk32o+P4NeVsulEfA8kX978V/87YpXdTjpFMbbs8w7GI
A6IRxDFU5hNL5+RntssbU3yzXcub5i8waf0I3VdFzOsXXqehGR09Mo2A1LFLCMHF
Nhx/CJ+lryUXBUyghCXEKKQAIZI9C/v3lTIihjDfJQzW7qmhXGI3iL9bZhSfdu/x
+xzF0P3z1eKbTlaPkwMarhfjRqlfcvKDoXYu34OwH25+Ue4C1LjPYdA2llOLtBBT
qrsSbvdp6+0MguTjaXFPiQ2H3+itzCAsx5KWZMrlj8yoqmI330b1feyE+yDED9CI
yz/0bbsGw+oJvfSU7koUTTGjO3dqNX0BPMCfFBZ5rt7x0OJ5pKsLAoRT6/67uSa5
2QBZHz2zaI6yMsG0GWWD3aQqt4H5a5HBGJKgvuNH6wSL618Ce41TrZWM/PoDIOb+
uuc73Cc1CRR7Cul/d7xgZW38kjsctpCYwtK1uPsCUjkKo3N5laKnsg5WP786UKjr
GTZ1rcEKsQ7KDhMvcR4l9uOKHzqjfvfkwyG+jogKRBjrbSO62UrSw4zwhIIqt+4K
MUBmgdOsRzHdlbsbA1L2//e8Ue18kTTk3bRsdsEtfTkHhgkCyMaK9yNtl0djLTbn
++qXSPWM6Eu1JAsz3VsBL6Y1IHmC14pKpVvVtdJnW4378wj/YvojIkVx5YrC0mJ0
+CSYxjHn9RI48TNcEIF8e4Vm6ATj+eeJp/XY9rVxvmRaNJipvkf6UlDFU1LED0u8
Jeohbt182GZCkj3UXQ16tFB8/LEt5KY459LL32F8nliWnmpIRcHEjHRFkg2rxn3N
kTz/S0B2uI7Z7pq37801VmQUM4lzTHFCoq7/NzJuO2PhN2nz2gWSZt5viWtXGCTB
l0WcDTks+baHsqkQpQ/4CWfvD05bTOC7NNL1OXOr31WiTp8NJiLB43sGk8w1i/4S
Tsa0ohZodutTqhUJk04mJSB65DrlUAHcYlKe1rXX6hPrPsutiIt29IFFLDLN+zIO
avbRRdDO8Ix+TYJV+KERlLtJn+cb7arZLtYOL6gGHNCOQunr4fLEYEnjieI5P3Bz
8GY5ZYIG0KXd0X29euchAzLsby2yP7foPgGo1VvrmTLynUoyLYSTNzx+iWtCcXXG
WeLcyK3PC85P/wgFWP3r20yY276NLFZaTamcvdyL9XkBpw/a90NeYuB1l2IRp3r/
BO75s7tsms918aQ7pyuCzrOBFsShnjxDdWVaSz9930+J2ag5z4k+3M371pHtXVyI
mJ8WGMSG6dJex8ihzqXYPOhLllSJlHaRPfK8qNAoIf5PS/yOnjchM58O4gKzjvHl
/8RwIbprRq2YDMoTfzJLGvFciQGVZ8l9nreZuEwUGOhZA26kayVeNUCjnRk4SXRp
EOu0g4MZzH7Tz3IcxS5XCx6xo90J3hSeauIlHIfIiV5oRej7d0GQArMfoPv/Lhfy
RJfc8ue7wXpOQ0pIFXV5quEEe0MjnaUUsqfAmjrmEcUvg0smk3KbMtAZZ4Eflv+1
6qlZgL76lFO7qZvKsi05wFeDcP+ndQK166QzhxkwFk1t+xHuh++qA6NQ2Z2eIcQJ
ogtcc+dHS2yRHDq8qF8uI6yjyOwgjf41Fnk8kekO7sp2MFBYR+r64MFQ89o8pYFo
gWww4QJI56BCCXwgpKhlrz5LboBoMVAI+lzjpAhVOV1s8QBi0CzL7Tfu2tnwg8tZ
r6rH2dsYABo+DQ/v+HfklsHcKHxqScuSDgSBa5+vQLwwPjXIev4OqXzOa8Lg0rir
smtFeoZtPVT9Z+KY2pUe3JrJkRfal6+0ZmPBSm/bIVtx0pnp5cNeC6ggDGRVUz98
B9H8HrCf/lVNzZGT+rFwD7wDZ7fpu87oe5MN3ArhW2ISXoWsG+/zb1pzjFRA1i5F
ws9C8a4kn5BCIeK0OS77SOZc0EP9EFCJ4JPacIlM8+bFYwe1EkI5nlGIPcaRfu8s
b193OqTBEAypHAfSDXhzoMMjYGJeQIDbDbQg+ZpV0y7h0D+B2edDp7poKz05gzzC
AeHuuVU3v5ywuQF/yiqO69vF9asW3mwjuFasMui3AaSOBBFKg7IGxg5XYxmF1gfY
lAc+gcTZhs2XTdg4JQaTkPTqO9GDTO10ss++80AV7Wq4/59tEWqHi3DTmBBxVF5/
peY2A/ZeHezuu6v0K4d2c1zUTeorDX+y++3RMqfQs8WXiG6rmEC/+SnjNIYJH40z
CuDxou2PVPA8CIughE1N/EHn89civ/KNXc/k5GamjUjgBR586IdD2nj9Rc78PJmS
nKwR9bl6TSf9hawXM0Nr3Qbyyx5aRxNy0maDyIBdIDBAZjWLPCcWZEcyfTBj//zJ
SMwAgDkdeyBk0AUvvVfZ/+I2CF8etff1bkiXRLBWH5cSVGYaax6zlojLILxWxogU
ee08NBoycB0XnxdG9XmbC2LgdVf78P6f8rE8M49Kprgv6L6A9dr3AEiKNTcftaN/
qQFMPvmp+ERCzsMUPmsH91YmFIs0hMlpBZwh4n4WFezu1We04GmXQg5bQPhGFtUC
bW2neibbO7TnHj7PvpzqEKS6Wfp2aXi5pyXvaqz+hGxwc9FWHZwrfOoPp1YAt9Jo
Q9d68DOwaOcOrV2Mjco3mxkY/g6SOcqw/XX2Idatsu3etlxygfajoQf8GsZkeM8R
jtoTyOhEVBlJ4ECue3/YRTkzCap+c+gNHUNVRyTNKn1ZY5V8/qR1XxkS78lFc2m2
/CQ0Q+xIyteFIRvrejBGc+dPPZ3QIZvuLlcMkUea6YOpbyuM760wX3VUMVm53wTj
FGnF3mEtGEQvBcvxrJ3yvgtxFbIL1JzkQWDNy0B8XizDXWi6xgKUZfe0u0MuwSIM
ZWg3jaTKLvJrT+UPoR8i3h3rWJrYT4gkZmtSyUer+Ys6UvTvr8yeHJ5UaRemMvn7
KkmclVNDoYIncIv5znmCYi8ccK6B0McmHp2WFhLKI7bVE24H28R4VBpILSOmBBEf
+8jOeiHlyKcr3BpoIEdMm2uaexjEXpLQF+VkfxMWmmh6q3Lqzrn3jjpwQC60THqw
U3hFgq5eTmMzuOJEwLp54P9nfpF8IQ5Gowoiv6bD7bnYf41TPstuv8J91zwC+cFf
/SkQdPuO/Xhmn4ja1KpjPpVtLah46J67TN5GFMY4F2Dd1/4AIxVPX7z8/cDdtK5J
x9TfYfCzaomV4SshPGWlyY6m5RwJNsBQ7lqpE2Yypk8lEhP9gQmwd5fYCMqGKG6F
CcYTtYJCbkY5IAPjuGe6nQSKtZ4GOGwiXJIxy4B5j+DocBxg/Whh8p6GlF6TuDLx
h14W8cvH/4CELmD0AEK7xme3rhY6e9SHWIHuMTg/ato/lUBjdne/Z5uMiSNWa/Jn
oahANmmJycHbMBbrviLGGmWyYcWI1vp10hA+t5TB1b7Hnt9xhWVM88eLMtwuA5TO
QQ+Sv0bTr8/XM5WvUp1bERxRz4C3d9e+kgLs+Yyhnaia4CwBdow2VStAA4SpXlKK
fNJm7EV9/SHB4b6xGKBi1GJAazFH+MQRUlftnQDrNPUoGyXPkdUKcbcGjnRmZW9w
+7LUDw9RR4skSka36QTWWM4AEat/7SKrAYow4sejoL918r8OEPmWdWHdQo6xm0p8
jbRrlXOEKvvybf86enL1Hw8WFXbOlCVPOczyjdUUvn3PVTm0IJtU59VkNAOyPAOv
KLjuOUO5aldd5OFQ/Ny59ct2HAOifU66O24b0c+0UI61DftmqIBrGHJV5eBUIczT
gWvP2uHl0HxwZJaR31IdiQG0TGcgdEgTpOuxHMBesHp6nYf58jzF8YDfo4rY0U5H
WQ1alAvyYsclbYciARV7BoM1ICyqjzCYCJYSMDtby/U5Q9q28g13HyE4A898p+Vf
BkjPKhTebkeoMPQNP+keKzMRoeoj7qAknarX3y+aQby4L87lwfC1LjGSJifnCo44
pOB9A3GRJkBxjY2C6hPcZlDhmDJZW0fr7m+vLHEhw2K0VH4T/mPN8oTHk7ptN+VH
TRNUJ1gBoGB2rHFS9FOQNbtOGEzFvWmCobC1Ane6b+kW5QP6AI0p+uJHGjhv/E5v
BhnbuLYTfuQuxyXawWFSsx3l3snRx8zGRvDgPOmrhh5vszt8gLh+3pE9QVO1MWzc
x0y51Uk2h6i2k4zq7BDEWylWGPgfWpqLpI3A/0MQ3q99JKrHDz6iDYxJNG8EAg0/
+I3obOARzD+GjOgof+kaUuwfma+/KQdWEglznJgElTmDi6ZFjUZUDyUu4y5DQ/5l
0E4hHlmein18wB37Ng4t4ufv9PYRI7OMdJVs3/pS403wyA2GidhSF81o+qFN/RXS
ynXQnfaLdbrv2vDH3ol23fCsOU4VXcCGYzpwqXLvQo0bkVaa1Lr9iVbf7jud6jCp
G2gP6epg+D0UulMAm3TZNGa/6rQNzGyCUBVpSjDVM4L84TGOb2UAffHXrM2w45yp
StuM50mt3b/YdxFeRQhRPDvoslY+MUc+Gbc8nYFuT0IbiFYSMyGP0AEMEqO0axmL
s9zKjLMWPn37s/vZ9nBkUgqJt+hlTj862I46mQqxhPCQIXABsh3pQ9U1yvVQReWx
fgxbyA/cqR//1bMjj27QgwNOrG7d80sSjVPhhlP1ap54STRy3uFriVHlncB3Gz8H
KTFtUgaUonq/OEAPZ06qw76tNm5im2WnzERC0BqZJolVtyVmUJjmuCd9k+Q9ZsVz
E+Y5HBIawwtCoBS62ksJk8UUtduAc20HdSvzpnzPHw67IeXB4IUV7TwyjQg+CCi2
wVxYaudPYSWpvhjMsZLOytx3YOKr2bnVO88cE5tP4vNMt90DxZVbgZmsDtVlNlh6
Or6dEdcMpZJhgr+JZbN8Vb/UzsWjvOpf69WIkNKHqqtqiAjJM5fKInnH8LRrsHsg
WNWhZRO1pW7KV9+lVpAfYzZB9gU7CuzzZFvg51v+pJ0IPhO2f18UCL8hbPtoNowS
ZENIutcPhZkOq3oTKAszByZQECuU/nGbtLIe4kJS2qCXhIRs9YDhUBYuKSKw0JE3
ixz51ibfSn37xkfKgSFQ07y3jLi7DO17EVGLa/lviFAnWbdxPFqsgPRzJ+GES/3p
HKQR44K4zTBv2CTa/gAmc9qhD2g0n5O9fT8NZef+F1AcBbszTs+fofB7ESfn57QS
hZdkOmgw0LUjfeQn6CcaNK5iAO9febdY/7GpABpVLGAe6Nm1sanISFTA3+oWDRh0
KBWRUot+aw9AbqtBLTRbCxKh4dBBO7ZqtAPHg4q1+aQ5so/PLDbxFcigCEN+jJ0j
ez0t4HN1zpXAw3MK2JwbW1ixIxlZjN8RdczKsMEnqipigpK4vCDuPuWloE31SqMV
I6Cya7UnjFKzaJINfXS3+vecnRYyiYZbP0+sg4yRNhOoI6ua7rX0qcGo7IA0AvF2
3MYjbwv7b01FTZLc9BMQx5+Koj/mSBObEcT5SzekzB/FRKlKJumW23xNbI6Im3Hz
r3UQ3As9wpW89RDcLtXyK//OQmUdv1Jv65Vh6c3dXNA/vl9sGQa2m8e/IwHtnTsR
lwR1DVD4T/qDPGc1fHuU5YZoyU+GB5DhdZU12XI+eETpbe5B0xvm4j9p0afHLDBD
COqV97A2oEiGK/CAzMRZDOp1wkVf8EEYzlt7eIN/w1hXgbcZTyXfCrcLdrO+RC9S
hlhwV0VNiEgleNKP575Hz1yHeWGHEhGHcGB5H1/Meu5AP1LvMSGatRONXUs8vXVj
i8JZhRv5xghLo1JeZJ/HoKOM+JjlaYO0MIndfi45ZZuDHkm8B45yLHxuYw8hgzk2
LIp6FnuEl4lOr9Vpen/Q2OululH4GYmTVH7QcApiKdetjrQEjOoez9aLaVSXI/OY
ariBZatsNzuJCm7sLOhx6xzkcXw1qes0RMmnTyviAwGIYs6U76qWdvtGWBuhWUqt
j4KSyLmvBDOUSQECOLCfZaqQMD8XY+qnYiLsuGxEpHVpx2IPmtUeIYww67f8nPLc
DREFovsqBf5bp5H01YhhHLZCCSr7hhAwXd6GbjE+faVgHM9kR1CPRd+AU6Kl2qyt
c7hbtdkH9i1Vd+9miUSsjDLfYPCLxUSi6W+q+SrCIC2aSav0ZeHljhbdiMib9I+7
fha8HsUWPly+o5Vjz9I9xzn0hWHY+YiXuHTupIBKVEOFZKbFViuH1bphSBFPCiwy
puJSZ4rZKCob3dr7cQ0OOp55Fj3kuVPOx00SdxTriG39+s8gqfOXmMjCgI0IK7ub
7TvaYH2QvPfMcF1cbRZ88LA2+uhguKfGlusRArTF7RuU2DN5ta1H8RoUUhRE6TU7
bJVdJLjxi0iIw0la3SQrT8RBJCp2bevF497W2HLa1+qVW4UfdJ/a+7YPr9vJ9xat
WecvEOkVzgj0v9KwEDjEIMm4BbOKB0UPih3I+hfc3RhyQHFx2MqKsjIrCfvSo4WS
+eALEvHCFm3Tzl8xar42T9qgzd5eyPJYejH1eOzhd0az0Gtu3N7oZSB2n6qgyR7v
FhY7iSmnXNCMdM8K1Ghla7f1WBndjUiGw1AjwIoWU9NYndLeIin8QngYIDKu9YPZ
g6DErO96RoA0MnyA1IEBNYN2GgcD9X2T3wuAyiHnXuVYAuhxzdyOom8ZBQUwaRAU
knqiCjakaIMxLoCpQhnkyqct4Z4ll/ScmE+GzDEEYMrEWEu8Y5sytX88xmu6WNbg
vU0yjYZdWMjMlOhVG4ZHIRvZTNg73zlUbYzeF23QCl2HB832MCxSo77/gRRD1XCx
E8OeJadU4NF0DklRKvD6InNxbgp6K2n7E6CFcnjjbg2CQsz7CoiMI+VunQ5Ou7GT
oKDJvvqhwHrfUUB616PAz18Dcln02/DbV+FOjY6N9fYZfF2JTadY5PF4uOvhCAtz
DjA002wPtlw/JX2qKNWtN2+YOVkPHXuekqa6gT6u52MLoqqly0k/A6BUNelWRSl6
MSy+OxhMCyvYTHyZGjh3hPpzkfqQg1NQATmaUk1jEbJBJX/245TRAfkd1zwGK+cK
v5nXS/aaei/cCHR/EFNlqY5fC9eX1xQxiJdRLPrqQaegAt/foYFcHg9+atCW8ds+
kAfuJGoXEAAQn9+V2RXk/TccN4voE4qYvXFph95mWRSJYp1//b76/w/v+UELKg5Q
OyQekpRsiZNPFRCODakB69FghjkgRGXqD2Bb1GCrjocSgiogSXa78mebA+3z3m6p
YUiwJBjUdfSQCQiYEkk433GHyBR1h/PpeaXPL/D6tcxZ2EhVpZlv+b+2grS0GdsG
3UMLFQpe7HNuZnWpiKTXVNx+ltZQ8D0DUsOUDIxpcMnckCYoWzdSaGvl0y31Fs2F
ijm3chiqO4Zv1hGE1/GeGnZCqMDzmv/NsmO6ouya80sv9YVjzo26OQVWrThDmqss
JvvnevK0wp0HTdOkOGBgjl4rXnfoS5dBPwaJRVoIVCxebLrX5AvCmiYbe6mzXkZZ
sHjS+EZfopJS8X8ZzTJR/cEi2O/gfSu1a2xZ0NB0Un8YeZLoa/2koowQmiaItPZj
2fCGg3PQuQrwZY5r5m5uHhwRFjgFjNj2fPcJPfjm6DX1UEVzrXGufY99166utXxk
pNjhHpKUsMxwliCDJ/zZXu5Y60A6fwU9Wik7k2WAUL67vyd6BhpyXxwXA+rL00av
1wgrWMBGlSnWnAx+trL7+P5F6dmGxWk3pu4tIPmDnqxH+4djvrQ4Ocbf6tdhPpPL
Je2LqoMkJAow/TETfbSm01FRyBr0c4yytJfZvGQhlYe99vRdxwAJY71EgfMVGY8f
YwpHy1W/SyRq+6fQLxrQ40CKsxmGELRgCC5NMu61wNQYifbNBdcygsQntQQ7hWVd
djXUdBH4msDWqYIBgIahnf+KLjD9nf7TW27+AXkNCLIqv/TsMh+2fyLq3TqXqHhZ
8uFG/zDxwy1HMrtLeVQDBedwpapthL11VP49EnxI85H7fg8j6GroxMl3CpJNb/Fj
aTyCU55ehM/cJl9ag5Fy/3ESz5FRHTOtrkwSd1wzXfODpv17heu4F11XopfJze1X
Y6iTvYlXwAz7DF7hcC730ikDfV+eicJty+yAINUZt1CA9uTHWqdj40HfZL7Mxphz
wXv08d7SlmDsOdkymRrAIcoOqxyV2zgH4yNA5YC2ariayhhOOdSIZW4Rw4QjAvyE
avD7NxVpva+mQWBrlBJE0fLSdxRLQfU4FBSGS8c+VLFxAGalQxK1e1IVaA3cWA17
7NDO/6G6KJ0knnjcx0uAkV72LnywKDUVoC4pnLKTh7dxjcVtFPV5hz+NevjUx75y
XRRcA3c8djMUurp2Nwdz99hOkrk5zYQXnQ/ZgZxGJIQaYGePctM0zHj0jImhVR7B
xU9/qgG4M4EvyT01PpguQ1XRoTMZ1VUAFe5Nyx1+4rnRv54KAj+vROTGPU60t9cs
RgAlDsJ9MLWs28NgkO70IPu+9G6VMOAHADtnO2r+vw6PN5xWxYaHrSBMZ2V8Z/8z
NEOkfsCQ7dUbYnl476X9oJgv2V292hyggpxVU2ORCCpEdbQefAODwyYyYkbYoM5p
iVJwrdMSVh3ME/Sz2EY6UhWLp7O5Qcvjh6PWry98N1N7MDvVwdWZEulIYWTLGJDH
T95VAUntbP5iYGv/G2i0MFu9+ygROqCDKk5VM0VT07NhWcGd3SjwefmfUOeBL//E
mss5C8vOkUwACs+sn5SFaMX4NihhIl9+fkfuz5oYDLhHeYEOdm6e2czC7E/XL23d
Lgj2SADbIDmUvD+Xib33fekIJlgrPirsl8zb4jROee9T0sGyXeO7SIJ0EeJHs/m1
QDDSj/3KlLTq6O07NQpYr6adwiNG+rBTS76Nizq39Eypy9+SThHd3dksx/RUjyu0
PoRQNmiKuxlh5OYdToGZThz1yYeTF6sfI5K3f2H7545rl+K2BxMcr8DukPoVcjXj
6sOgBQ+0gOnvkSXIDQDvfYSw/3Xo33Y/sbTqoO2FEYW/dv1OkK2MrLiaftFocG/N
gu+Jd9V7Ei5wVApRwqcfL/RqRzRSMRnLpOsKuKU+N/5//DYwuxNkDoCrENJSKvn5
ce85mc6lNg2KdOPeqCHIY+ekjlvr1Hrwau77JaHWqKicqCWqRnJSEBotqLDpV8jO
jmeBI503kbCNI2xOpA2hPiZk1keb2gIoAic40BYPtarEJHCDInIQIohAszrYP6hz
ZnS1AjjYZO5x2MpO3ydEG7OxNYEGbxJxUGqj8YFLLBOTuLzEYNprxWTetFdxoHo2
A+p2AyPeMm/UYiPetaDOyjc251pQJu8oF+boUW1SLra6H39bXmM9J+/VlmgAfVUW
T4XLNcylRF9E06icarYXgBjs7QtNyn4Lf3xU5fJL2nqc/cmFvV4skDkeynG2mZLg
ejfzlRInPme1UvKvy8j2QZmTSCtaUViBqvmKVycqWhHwAk+YvddfjqQftDklM0/o
pB87uOSQxwE/LdxVod/dKrUCcN60O8WLzE1kHpIj6ZR4v6nCwpyq52ZEuRk2RFkP
yY6Q1VaXr0ibVadiR8s9wtd4aFsNWxL3EBgrmKRBA3tzCMGUKSOC7Zjv82rxDtbA
xffQBY4j7Kvtm8NlBaSHqthBtj9J84+Zlu2k0/3EGFqrXjwjaLG9zdF5gEA8hdzZ
W+re4QIuS8v4Wzav9/cWniBZD9w2bm8wkFN4KE2edJVrnZ9f2QMpL9v8bpq1jBO2
0df5/hPfLSxyWq1yORLSs0ShxbwESY1GgFRnhaWkwHBaLswvp5zRstd3G6ZadBhs
nSaHTi2lzcte1Bacucuhggn1m5CIxJodMPa177pZDw/VOHAdA40pXED5MdSyJT2y
pvI/dqnNyTPI8Ym7RpiDyydvOc6FyE4lK5Ql80SB3StWivCwG4o8ZvVDy/UUUc8F
1oSxitbW76hbMQFcPDsuoMGoGYHr52txhHjyPaUACOSouEqcTXidrqKSFm91HLTj
U6eIBxwqQS4ir30uhBxnrLgftkztf4UCRJP5ovBAATLv335FyFPTYYkMv0DvnUby
R/hAxE26/ZK92MRD1t9dqfC51anmr2RZxPkrctf87D/sez6J69QEN39b2rxByP2X
BlXcZQFaK/SHQlN1DwitdDWVAnLMWBnZ+d2InuVc7D0F+MDLehaO+nCel34nD+nt
gjXu28DiUiLe4sTgOO5/3DNogIJnGHGuJVkigFLKtxsCXinzWzRB0kTaXn/V6e/+
MOoShTYQmpvF1tqVy/i3nSLyF0L5ceXRBDUPioiNN+ZSx8RWtcIAUFCIAd309+XG
U0l76YyPdkrhSb+MSqXzBzQ4ddQFgua1PASo/Fzd4D/1XwkT0g+6DZE+k/oK4x+m
PnPV8pBAu8er6TCBtnxUY91UaOI3dRVlqClWHV1fbw7EDr4YGXFPUH8vbnkehQqk
bm/IczNd57GHRa84Dv8iuhcbylnhqkYzTCdfC519ShUP4SL50SKsmmDiTe96zqqr
MTQDzBsy3eKGC26gYskrpplADklUjZ1sTRZkv6WXo3pXJnyVzJaHhV6p7FiWovC2
S0twyptWiRrsujzNekqQvTeXUSIUXRz2nJulLTc4kMpH03iGg3sVloig8Zk0z6qA
KO9XFhj/wdQXp9FWfHIhiA8fpBniwdkaJjQ4ifNnnJykPY+z+YmLF+enkn/guvzR
4Jkwl3Y/zeT5gTgixk29YVFu/0xn05archbv3iJY8+94BYGmpFzrmtJ8m71pfh9A
RI/+u6dmWcs36n+6RfmNJcNNTlPk+JKHsLfpJq9JCkF9EhQKl5RhjMNW2cUD5mLR
AQ70iZxvUN5mQI35wjCBCXsNajNqNzlYmtIUMAzSNRqH2redkcOVbVhh1RIyISaZ
PaAaPhjd1M2Di/XILfuyTIJf4Wnbgs9gpmem52a2bYfSJtBywJyiEYrVnbqbDrvu
CAz0NX35E5394hKCLzxpolxrwuy3XA8r/P1OuozLLkxTnD6GPvRgRQt88Xy9FmTX
IfF14UroNlF63PwLYfxjhzhF1GBzs+u4IRrUDFm4qEln/z99RXl7XXJbAR0VFrRg
6rRYNGGFrQTycV/sInyKoIc04Uo+d4+CRbScTKjsGMABfR/4DuZ3XreHz6TFzZef
Ze3DAsyKhCeylvPlPMsKI7h4AV/y5HbPJwJ2M+e0yln67AaWxGsZMB96hhfqM9H6
v4Q81ecTLcwGRuw+5qEybvIgFsKtooZjXqU3rbuxrS5bY74mjFveWMJ5AGmc9GOI
tH9bk8kJSG0E9pNkrZ4JeR8Aepaod4pxtZm7x8YyB8GiAaQVqH6QZpTVBB03WHnL
cvVfUVK0r/8SzxmBV3jWDoEZoRg86aU6qY5c1/OHkZzZsS8mocexN6Vtm8Tka/1i
zTItiFE7wtish07zQlExZdP36N9wC2qMBM4Pp4bx9vOwERDWf3Y4kFw7nE+/GziD
0ORZZH9pSyHNLvrBC5r+UWm366lIrINH2yWOlAO1Do8MCjlb988dY34CrA+rh2ic
4Xjxwejd2AMWKE7KAxN5EZkI9mZTCjjdcvf/ynKnlrMCh6+DgyADLdh1rEFuzQLc
sff3EEZ+jk51wGBP4W4eI9iSlORS94SWXbuGRj5bt83jiJMC5NGefJWY9KBEpb9V
hpdE1wrFlhNF9RncbkCdeBe4ZbggZ//6EAvEb7fhTB4kaaWID84c4diPpp1RztqJ
DUz+tLtlloEQOlm9CoZ4yQcieaDxvZ+85hz5PgRjDMlHU3u3VyaW/Msd9UTLhO0/
GY1oV5vE+g6+cUNHqM9026dOw472C0zuZuCbaIlSWG8cacqO/7C1o73z0g/stFLJ
S07c1V1DCn3aiYKWRzALkC0dGZioZgugbew3lh3niKL57ssANoZwOtsYBZVnqdzW
r4j3n8eiaiMqmh1OmS8eh76nlMb64lvUydGXsScGecOPCWR6W6WOoduo5mtFWXna
YJ4o7zzqMYbvbsWiRHoH1lCBhE2CCaiKY+5TePTmRAJWEHyGrVlH6BXL/sx46sXn
lcqmcarD2/Hzlet0WGcGoicDHFhF49M4cfJY3zWslup4Qz83tnY7fDH+OL4b51i1
3rMDW5vH5Z38+hmWItrFnPi0/VLq1cM0MahuhLx478Hw5PqhCE6SDYQ3//8B++vr
SRvXOXgT9RhEIZn+ERA3cdUHimz7Cs9hpwLdSnKuHZfq9CM4QGBkxwMgdAmCq0Ml
ByMzgvDqi4YzwSDt6cLWZymqiSD/YYmx/N08szpc2MEg2OH5RcfJa1P2v/lbTxMg
OdK8HEWi+jI3kC5DPjXP+cDqxECngw3+wIxKEKe3OpXJjaCD52ov+Nl3FQoZQs5P
IKSQ3Bsy2asa97Sq1gUZJ1QavUeQCmwut5YmkXDJqGrte5xyFF/RXfDDm0O1Rc6o
xR3mfhhf1Sz7iEEloX9zfkuw3VIA5fCjdFTEr9MQ1Rxjp3zhYFh8/j6SK6svGl/0
PujHHax6RGVPxBPIzEPEM/q+jLp5DFvLaUsfnS3F90hEe600EkGpxWedzRuuiU+Y
s0E2oiIaH1+3VWo+NiD3ydvTmJujqjg1npL+Twxl4q4AnlX+EGgZ09UAR6XRFfXa
xAnJ+1hCjscb9+nq9b5m3ry0XPigP5o2AYnNpXHdGRcZim6Ac6EbH6CGia5Xhlps
KkUCR2jnSVVSWwgGaJCkAF7in25AG65X/0rLlIRlkxFK9XXXMHWs818/2Q5rf4Fi
Cv35zOrksUwl0HyrlHYDiNxPHVrbMS5zdVhamqsAiw0TStnREd33HlmqWBFU/zwr
c9JUlKNXOyoLum9j7UMLazOEfP1PmM9ySKEkE22VQ7FdpYQ9Spl/EXhNzcOg9ZtF
TmGDzPUgrYNQjpbe2Ik3ZAIUEKnLqIg1uHub7d60FqVBzp/sPsOukeN6lhVt4ITX
CF4rRGBotbU7+sNA+6MKWCimbJ9YV9OhBbyMaLg+L/Bp9QPLyFNRp6DdTWEHkJJk
ocAlllya1NDnVVEGHAdD5T01mdDlfd+SI5eUuMyW/4Z+oWciW+DYPs88uDqMCJfM
k6a8TWP0V7kV8LLsg53eHIXqqbck5Jz9kLxRiRtxxtPwxNivwuJMUBGkJnUBF4oA
BvmpYHGDI4k+Hm+kt/LAvpnMu7xQnTgqNvIjZuxk1uvLVWjmck3u9YpQc3PDtFHW
JQLSoBR1thbHrrVplHXAepPURh7M3AMU3k4nenLHc79xorAnYoEtIxB7zRKVY2Kw
x1l2bPFDb9dEx1duqsLCBTxqyaNt1PjwuPFza5Chk/OQLPx5p3V+r7HOCe0VZP8E
QfC0Gs7XSp6HPetl4U4Av/2MVhPetNqJJk+jeicm9S7RTNj55HU6Mdj1tG80ZrNj
Yi2jq2pcJ3xb0AyXV1aETWfg+VM2IYODOSXRubwZN/DfDK8R8wMqEzIylN/rrz6s
xmcHLMJreKWdGpobl5yoSl1heYdAQr2kFAMCZr5oBttfGY2Qsv6JNvJSjYx1yXzb
z8HP/dIqhyO5cpzA5Sd4TuJSEbwl4P7RamCeTJ5bo/R9xRHEaUygYmwOobFvc/j8
V5QCtgw/qr2dWEhI90rx4wRvaEekiZ8Z3gjpML74Jkq6iv2OyPgMqoFzXqt2Pi6F
uKq6qlywxIBPNYek0AIsVnz5v4tAI//UN0LLujBZdkJPyvFfJoXmAP0Cc0jRty+8
fiDKx3aW+746tnu/DDpJn0sBOquILiKjJSn3Nj4WUDny66adxWZvrzsrWuXcdQOv
eQDl+XEmrOlshwaPevGcwqsWy44Y2NJeqs3OX+xbXgo3YAmDMZD/53i60EwaWkFv
5FlKsbARX3mEiywuMKe202cvIz+LKf4ewLjEdz4b2BEEr+sm4jKNFFsgWsbHpLIs
UwFRftJtid6RJGpgZt8vhXgjsGmbfku6cJpIVaTiTldHgOe2BxV0Fg6XI+WRMZnu
4B0gpUQAp8exddNNPpeRQ0HxOl6E1aeKWh+GIKAu2kZDDjs6cxnl/hZ6epfc7BEn
9W+1+EfyfxzmZYwY7cU8HOp7iBScZenpxD8asaUKasDAEgOnRyWhj4ZyYwKtuXl/
zpYA87BMuhuXmz2PbVoCE+KM31K0+7eNPaXZ2w4/l3wXEcR3cBhLwVxzr51tqv4l
bD6CFGKkEBN/2rlZvYj8OtWXGM4pJHUfUUNlsBXOOfAEpAV6KRePyxB+rWkex3DP
jCOBcykDCzSSKd9JXVuSVclnFB9AkfI6qr4wwMLwfdiUlNUrABOlZCRav7H6QCTi
Es1pJgmku0mvhaIJVP4nsXllE8tVM6cbXHcJ/4GXgFPre3f1VJg7zf7CrVua/5XO
HfUAcPJzHdW1iQVjVLTvGcRlWSoS8HzU3zDPFP69rryEEu9rci1PQpnpqXwM7tve
EFnT4kusdJCWsMlE6N5LjKIukQf2zZo+fda0N6ZVbUOL5Uoj770aKVhMTtak3bX/
jFufml6i07RO5cyOq7K+IaxqTSPOhBr0Q6/qzUnwyD/4tCNm/yFuxK7AnqMFlF5a
uaHRZGNz3zP/LW1c7rSUPjvLP+5iQzjiI4glBUME9vgyudARyFC3QsYp/sZ5r47l
/g8AR1BzCVW2FuBYZ4UE3LYTSGpj6AXNBTkMDEC52oL4zYexcKM7Bego/uW2CA1N
DbaKh9hfhJLncn3whS1UFXAmkB1kU32hXX6RuQ2rdM17FAN1cPkxwlVPmpOkLqlE
nI0KZnoTQh/bd8Dby7GaR51Qgtb6ku9NPbzZm09cwAS21IRjy5yOD+OOrqh2R0Cg
5silw3lDWqt8XZuA/Cz/lVmHHHHnvFu6QhiiBvNW0DiGxkMM8bJ9GombGhB0cCje
Zh7li8+QHyoqMWmwwmdyxD3RC7x8rhewHVLJNlyrBFHudE+RURby6+OAl7ufh8PW
WgxiupSCb6Q2a/ZEqyOfEnepbLnR5yas0EYzkJfvqy3Fu/TWWBb/390yfPhmkMQn
LMmfT9uwIUVACxaxeYDZCl3CA6PKKQ7fl19w5FZxhi8ZEyDoz6qIEA12pzE58zpx
Xx5S/zWH1jzb+sNCQ+3u2K5t47wBvBilJiL1psV7wV4qfpnCb7CFiz4cEQLf9Lfu
KA02XQteFxYkiFfgdZ3tHrrZh7XQ30lf1wqLyLho3FCqxOCQrl+OlEveIJ9q+8zR
Jg67rv8cCgceTccpYJVwTJ1fo0dROeH8TZl/FM1MiP6229bQ980crCdGb78N1IdB
VBAK3ij/Rq7DpXRnli7T/fR+q7n2Dr92944J8JHf5Yv14Maqg6xkDtgXpA7c+cIm
3FI+YQyW5mz06Drjjmzs3ovV3eYjYRIK0azzpQFHxK123EdSPEM4chpT6HAUshZq
qkqyb2PDyrm9RzTT92MAEciwbguvKIogFtAv02jHCfymsgonfG9h7AXBwTueuiHY
0b+FhMUv4ioaSE5HCwqwHUiPxsYh/33eejd9MtKJPXkMmIaxYeanlz/z7rB5VMr0
Osq2flI8/nfflUH+1mE0xEUD5GbdA9CWzZObOcqEE583U4RJECubUzjycrSaSqPy
ybyYgTXbs3UM7kQGo4PSwQahrigAXADrSVn9rsddlHzTorxcGdY4I7M40FH2GBxx
7xrtknC6XRGA0oLNtTK7uvlko+3QaQ2JiViQ0NMgxitoWmjuKCDuHgPKm7PpHFPQ
10wifggKuSHrg30fuEVQeT03dLiRXTxeQULXC4gWByDwSg3IyurtRdCcQ5fMH+sn
RbLVO/LTeelaDi6TupjAFC6Mu9yP4UXto7HokNB6uJu+gYgHo5vVBPrj1UntxYlN
y6hcoeYg660ioQcU8ACuVC/kY6hGfm5/ufFxONXWovkY3RLxQ0hYrrTxgz5RvTF1
WQL5qypROCVHW5Z9h7jJmckIbzmwTTD7ruqLDS2Dsf+u8aZpAHCp6dQQwxIgCYYi
ErAQKyD4eZ8559AeyxnjT7F69FxqjN/lo1no08mUcUtC9vzHDCioqsc1FaslmR5k
aVP/NX9lyZ0x6ZkNC8bhXrrjU3SuMjTPLWyhlKd+i7V3FaFc9yMHED2c7xaUbBbW
L3RwIkppnvPShh2r3FCGQe+IBboM5rUsB+esPp974mJjjihIRJKedJURknIEC/HC
N0on0C86XqqKDAo6JhHSEY/0QlSrhx+v1GLWW0zrH4FzmYd0aIe3yU6w+zTTKJ8M
xD57C236zIvXklQs9UU12MQDwhvzKPpRw95mX8QcB9btcKoXFLXfQl7ULsgn36zM
tSnzIQBIftYkcwNWtDtQJL8GUT1oio1p7etDU7mxFYD0wYUepSO9y1pwjCBC3eGe
DAyUmUGZeLkk7u1HI1CjdYmow37Wk7WQz+GhPhdevqlPqAPDTp3vnLkntmFkm6FJ
oshLOACLY0dcKyEAt7WeP0NnbGvD9baqkL+0WrTeMvSEnLPN2TDBYyd7GTuj3F5+
hzRzUbVSju2IUXS9q01PARBopxIvTQ/XKM/9gYXVA7O2NiF1Eqrf54RvCria18G8
HLMgH8iCXggW70gqhcjs2reM1sJLRgxVDPaCX9EFK8+mr9RPSoTvTk95aKY1SHOx
LLG304DYEyC5cJmvlHdM+HoQomp7CUPVgAvAhJnkp3BkRPqZbvALi4Oe6zJHAmzZ
onOLzkDceBFeDT7yCWcFOSFmn+Qj/6CiNtBzp70pufB0DyE0fnKe7q2YEKRm3lBM
5Wt2iPwyuTc9W9+ahtQrgJ6IVfWDUNN/UV//mcyg6G5kF945WSP5qj0a2RfYgIq8
0oIRAQl3Aa1Q36wGlbYh5TKg1ByEw1reqUNiXfo9z6ptagUyn9YByJCs0DWxcDUQ
CutWB7OCKcEK8Ar4ajNe0b82SG/nPfkOmdX6CS2hMm7IgqyKeT19DDfmmV3bt1//
F+R5fn3gnjGKRS5If7Fn7JWsQW9pLo23OgLMyXIiSDbhJH+/QbLGCOcGBUerrq3l
zc0SbEn37MIRRnZH1srNpGVvAI/kl2zfNYz3DYleuDAcHxjevCY5+8XgJQQZMU2G
m2B10b7yXNjlEvefPuiHh+sZLyQeuJzNybI0klfxd9hGdVs1yykNQ+GebwncdOwz
iQLXGwtZ0lBLEHAQJxeIg/qAITWVoM8atD/ulvEzgZNKpHA7FGaYxcXg/R9BMqTl
hYwY92rwccKdl8Py4ZXXN4FXDrQMxvQaTUed/bE/dpQKRbWAzyYhQfCJiXycZn5q
0VqTS9/35N3140ta4GLMdinGfoDMl2QlKver7oItagPE6r6YIBTSqUh5XzXSKkkh
R8obTtCzB9rqqJNQCQZwu4gm2xqkd9NYeXWNqRGITeCbSAOPiWNY+Lflrd1jNuov
yRJaXSZPZ9QwPwNeNoX4s/Sh8LhlwKbmvJgF0urSHaMo4uC4yGm8wa2nkefsPZ7s
o/NZC/iXKv2O3Oo1p6lXtG/CssOB8WlUfB8xDeW+gA5foTgDfJdCLXsQgaOA0V5E
kl43VN2hX1/MllNNi1bEJqD2SJdiycrmhXLSgLnWWBy6o+s4M/scTH1527QLlICo
+tfeYhInegdWCemafI1XND7hRR99mcu8w7ZaA8vipNM4tv55kfSuy2HE0LDt+2v2
lEPWqR3bMN34wQLqRVs+rKFJAahWkAjHeHAZY+7372ZHOYTC/3EPWNpOd25+rNzf
EROfYtyZUC4FWpFoijz7rqXBouIiCV9A9mogaQu52hpr7OWtsr3gc/uoAn2OBbPI
BFWP8H5HijcrURC2ShC9jZj2TWBLHxjpBEIBSD6PPPs2aqSBg+okoqyaYDR7QdAp
VxTA8AwdwtneuwjDTXrVg41a6JdS6rDn3C5yxfNTurMytdrENAMOVPRoc+0o7ml4
dNWEmR/4v5+9Z7RXexeVBJqOuCkOOx23ItaEGLKcvwIK2vekgx+2C4nEMiez1fLJ
VITQbUEKcZCc49+eQiy/+BTGspXZIi7U208k994wMT6Wu4DSCbRokNECPUSnLAJ4
JCDk1aGP9USXT17+djxl9rYqjmFkDOYqMayt+C4mbuCH/xRjszTC5ByiC3T8lL4a
WqknFEPg2F7XM2EUZIGj9NDUWrAAocilNZkZqx8w9LEEPf41EWOEZGh1/xkaKJlA
WGp0FoHlX1P6DX5/HqJAjnCs/3cStvJiGRnGGqU9kxVauvpTWepsmIN7M/S9MRrR
CpSjd3/qTUSGL7++cGsmZJQmp19/MdMGUwlGJCFWjCrL2ghSSYmrcljYQm+L01C+
xgfrBVcM8X/f0IUAh8AsTabuC8aK5n10nB445+TvLUaQlSTw1MnZehmdR5IISi4R
u7c2VePeaTVZPDOoyDUjKyi0frOTqoSjuIIq53F45WCxGYDvRdCNiQr/gLCsgt0d
QtklGDXBgudZutQ9yA2pSsQ2b8L3gZjlDA7Eow6/GMEQ2roYYwjXwaGWhuGY6L53
VeXle2ds0cqlkisQVjB3h6n2P8Dpu/buRqqc/sSeRftHMIpr47TQtTPI8ZPYCf7k
vZLYeArrLaAvI0W+B7ow0ygsVsv9iPveq1Gn8xVViKw0Cds27eNYaq0KgDkqmnqD
MIAMgxJbofvx1dcRvZ5WTYQeTRfR+/7V/aEjjLfykd3TTQ0OO/tUTYupuXCnYC+D
JB3vhJlDPPgBGgGtKX/ff78ClVCYIZp8GftmyT5If4Gz7E2Us5Q5wp9d1JP1rXv9
E/mBVlxk/SOEH3P7LhNrFPT1Zn185oNYF/GZcoaoL1TbruMFRNgR0Mw9N+Q9bD8g
XRr6l0yokRxIS5QqDVIRLQguEx+s44CmlTL4sU9UzJhpeEFsZJA2tMEqvtDMyvTP
qNy9nlqu23iVy4M5vhNosN0qKeFeRsISzVzQcG9MJW4AXqhN3UOJxMq6MwaQ/xVL
1eUzFBvvAix8/by2OORBlqPawTK1TScQzL6lNe/qIIucOgYvovDeciubxrOMvSFr
X9y861DwS/m4sBLSFs18ZY0YoiQipaekp0h3OKwFKlsXym41r6NPJpRPAEvy/qhb
iSeci4meeWkG5KPpVESg49lTIqa7+XGAYJbqWj20ag2+XKeLTGbuALzfyAIuyJ52
uVXgYC0EC504dSSgpiXOlEqnQe+QSBT7mnD7vUtJY7uf6WvrbEWBkcovmrLTb4V3
pKG8jtUSRHU0q4VpPiC+Bl41kBzPhwH4+F+Qe4QPtJV7eKSsRgzOYj6J6mGUhHbo
JopNPYimMD8AG5p3OWxJShMhtojLSITMvVw1l21cnzTF2p6Vo33sWUr2n9teH1IE
6UKG97KdSoc3jOES3FDCnoaRlpaPfobghLSGqH/pGQMAKzViV/pSqjNWYrxibgaB
9SSxse3Ent5rY6vZeT15bBh8zQ8LHXpFj1EHfg+fvejFsTsCkF1Tf888ibmS9u7p
u1D9A6IyexptkJZ/gV/ElWwhOf3trDZClcRPXaB2HBrFbRcDjQdfAlNPLuPA1tbL
9XLL+PeUXWTkgpAkTvmLvFcWx9Jyv7zIjzcQN2X0DHJ53fFvjx9Q9jGXQf2zLAyO
NDwKaBxJMzZh2hsM4SflEV3HRDqn4hk+4guky87KmXppVZXNQoodZroLV60ajerc
`protect END_PROTECTED
