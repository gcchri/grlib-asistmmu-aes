`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8iMO47VYklGPCO4ScgMTqDDYMTUnyoIZyH3iObERIhUy3GO9VGMRzuDIaD/EtA5x
MUqst2ntrkApyKkOEMmGhKyGeszzuwHLzOhCdgcIPbsTVGHzlE3Rl0I4DvxMIkaV
h9GhJet9NmTDfZhLT2lfmnptlbC3zTjF3tEXf1uQJZgRu2r864/VJiUD58lAk+th
p/qU6aqhbYrUnEJXFbR+cgqV7nN2Ypf0Djwp5DFOPtW4nvqTWZ9a9GIjxJOrRGm7
76/vglr02DQwXTwFuryy2mXa4h0FfmLZZS+SVOi5V7z08KzyeuELqAlG9u/2sNFx
YMCWSAR5fpUskQXbz/u5Rm/KLHssS2i0TwXKSwcCThxWZXpKB6vDkjYSSP8lu4M4
PFEbfXX3rXO8j0XF+U07jdV0A0MptcCpZIEiAs8MB/GTXyjQtKO2aLepDM1HXnYf
VXJqE+Q17cbAvYXxLAf9Cq8uOppTqMkc4UoAxDRY4VJyMk4Xsk+C6if04og6kqET
mKXVhehwep8ZiiCAw8yxAUWDRNol7WJNCsIwNYTmQqoTFySBZmt7eWV9t+bY/WWE
r+5/tHQ/YWNSggSmXW/JDW4ZLuwXwwB7Lcua8W2dXMrh0fI8nGourux+k3zD354r
`protect END_PROTECTED
