`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82pJ7Wkid82BsX9g1CQ82sXDdo4+OMWFTB9un0rf7EXL/Ch5sQJB2gTN5SuHmq6X
6sfPzKPdT1cAFztiFobJDOsuNQt6mWp9y3iqoKmzvzV870+6BvDwgtdh8Z1iN66R
ErfnX/zW8m699em+dFJrWCay/prM2+AOPyDL1ayzB/Ce1RuJlvtZMzMQnuOqRiBq
KOz6Bee05F6W9gGClp/dNnP/dt51J3bcK1DhpfIQzqq5ooO4dJYfvF32RuSKGrCS
ANAQAHLLU4YDT1fjCwG0NevsqOb1jjqGelx/eA0T10CvI9Rs5Qs0MJmlalFkLij8
cfdQW9/xvf3PC6OMClglHVgMSnzI5fhUgWk/QWPzDJKBNPGle4ndbNmGcxbBnqff
pr4P9NAb2sLJLbgra3MFYmx4QkPPiaMxpDZ0T+E0eUJKa7QAYyMrOxM+eG877wPw
oZmma+Vtjc6+loBglH2nBUXW7XKJ2vvbifH591tGgjBX8LKcoQFX86Urdvtaujvs
7xx1D7b/uYhzfJPE9E+2RtNe3TS57VSA/0hl0FbzBmF5zPpfeoC+Hfx6TmfXnuKc
H737rgi6eB36J5NJ8nJaj41OsU5CfSN0Qa/P+TDcLvcUYo+LdZXSEBBOlmF2okPw
26LgNRjnAnRA0+zVXDzf6pdI1J6cDPj5p4AcxAsJHbaMH5TujNcCqqezHhQt37pt
zxs0vtNBgBsIN5VoXytw0jH+V2CNGTGb3J5aXCuPWfmtPnTMD0knLvpGjxfQFB0Z
EQNjpy/I1pbLzNDxAO9+r8b5IH41Gha0SVnpqhdUHz6BF4NDmpz+YrH4EBUs2Djy
WwdnwJFKZTsrlIwYVbAxgmkqw5bLlMnNlTB3eIpwkdyKZiZl1AsKqAYLV9hI9hWU
UvDZlEr8zi062s0ivJzbnJsg66xiREkJYGPb2GfrHJkjcCchjeek+m6AxTMklUZz
khSvPWskyk710wcIia5PdGTp0Hq5eGQkgvMwDHRuFtzjAbewwC9yTGfJgrpuR5nr
dXlgCo6Shlcejlh2PcYwJuCzyH/7uHWoD+zCruYW0iATNJp9/Y9yknfhhLn2MSJ4
KwQIaszq/YItuSg0EOR5psMeGRo5XQqw8WRDomt9rHiXEsMFe2aTZpPWNBHWBMWM
+jMMP/UPU2R5sYpFTsWXBKbEjF27ZscBjFf11Ir8oEVd81aDtEeZXhI/ZLkTIypS
0ClTBwbucUjpKBJ2iD7vm1ZHzCaCWB28tv8wxJgDn/2b0+GyU/95Thz4rOCO99zk
7YCGket2vZj1aN9XFtU0Kat/6p7XIDxW6QEpcNP7EAFTVT/ic9iKL3Q6Y97Q7NCY
IwlzEDlW8JFm33InFwL9Ub8lJ7Ztx/nXExtJV+z1k8WXu6IrJC8bELWNF9BjvmLq
gcpIKz0YAL9CA0irVqcfVXbBNisioJSvleH71tPVP11rDxvLiJRRKe7epZqMkduD
+TW3NtRadvgdlcyJ0GBSlOXW84PSLBv8o7P7J9AdkxUtM4zp2OykBi52XPYcpXmm
re0Vs3Gl9UKP5KNhFattqCeH3ocfCEpXha4HoP1fOihIcXfLbgJCSJjP3oZwoFOz
GjaMOi6UjfwdYEB6aNBSP7/XXEamdZXn/AmxW4v2zmDi6t+YacIFLiKfy3SLTcvO
pT+nsF+XdZ6P9ntlmPNo/F8XnkW4LpuF5LJYz+AW79AAv2W5+Gx6TGSi2Td0QCvr
TrSPadmkuntEgg/E9ZSH0LkoyqzaEMxGVH29383PacJWegJwARIRH7ReVqVknkm3
MvfuCgNF8TyrAfRG5pfGTBNhoX66okD2H+9FnUmbhyA5rKElQkAQxGhsfYqfI291
38y7OvFXVJhhzGpKc5WzZ2rwRL8MIli5Y83yjSHLBRw9NEpQLcoKPwe3HrQQ7mZc
//mPb0Swu3YEgKToudbmTo20Xib2IbLrnzdw8Mu2t//sEm7ZQH0TWST27aGD/7Ol
db8NVj8nKNyiVMhOlq/Ty99ZsydoX6SgvEFmNOzLrqMxr5xvLvWMR5E8XMe4JZCg
+4y4th9h8L9BUVAJ497yy2/LUSrir+6cwCS1pZmZ8StKGs14W5vT4WSsuyK3JVYQ
kFmv6hbuvibibbUXSkVpMYEOBpArKCIPmSOatS9BV2qMgzn601m16g8dO8jp9waK
vCa852Hh3rE6Ikow6suo/EXoLRbB+77XbXho8ns/hlPjY/8e2rM+m/hSBfTmW4Zo
wtbRv/5Zdy2qbTNshz3IVXpiQIN+0lDowKHOTX2iLSfkNi6fzLRE1EzCyPtMuxqC
5rF2RQZNDgqVfUbtfwy7WwrOV3k4WLc1zOqw2hfBeSXGbJBfbJbay0nmH6t+qaPG
qwZDmGLoABIkRLFF3Xr6OhTAy+EoXyOvBhXRDMuJJWa67zOoDlcAtCEIZ5SMeqHp
asl4VOvUFCUdA8qt72juWSYQKiPMdE75jyuVMcrq+JgPwIk4MhzFqSLgIaXPyPWX
5MSqmBetdjueeeDQu+KMO0M79qcSVINV5bye6E04FjOgu+WDF0CqqiKfwju4SlE9
I23pUWDx048NDrBUCJtx+BJRlQg7YSdOD6wxWVLTt1SxEaAE8tnPsOnGU9bEJV/U
myCw4bNu5UwUQUlG8oRFMpcAC2MDqM/BrzfRXZINHGu7QpBzoAo3+Jmcq8HpAWdV
INRaQImWcgzZRnxF2B2P+FgYC0/awehpygl8oWdYMsfNFAPA+spiDh/f43B/ocFQ
3StkMBvFt1MtfGi25KAyLjATf3RZUw0PwymFvD5g9Cw7MLdmScERPi+EeK7X5E4o
lv8s0WzjyWDHQGHLgBVtWCD4XkthMCDzTboqBgNw/8bragzDcyQAaW1ndCKMbuHU
CK1fKU9Da7JnI3Wj+E0rmzfbmYGZGYA0qsXyhSLsgz7X086eyctzvR9/4NVLbBdA
//Sok2box8rts48vnxqprzLjt7tENmjNSjDmHxhhsu5mk4sYMoBsZzLvKAHezllC
uvPqlLfzbVKhbFjQkrvpgUH/uadTBHgpL/7k6rbLJg4SW/+SVCpFmtdZVL2bfKPS
RbEQV2NAQkse8H9s9aOGnC4mVj6U57Y4u0xMVtnvG1mhzcHYVfeooYxSEopApeTg
jJ/17FqVk+9qtPl2i7UglS7LexniHEupaiZZm2lupIWfbFwMzWyLfLankfoqsS56
8xo4ojJyeaFaYlNNlgHiZZjTfUqNvkQ67pmRXxfMpcJQH4T6EpVt9cxis1jy2kvc
Ti3KveOqeYiR47N6Cfh+FCthtnk/ucT82sJN+hPierB+FbbavsvtDYvSg6q3qWnS
Xr5b29EDg/MyTNgrfGJsQRKRQt/QBZWLZ7hm9XsOGkydHOFrxLNoVr8c6Ec13i0A
THJVkv2Wv9f328IAaSaVaQ==
`protect END_PROTECTED
