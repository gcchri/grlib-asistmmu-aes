`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RBvOExObgHGVC/Dt/9cB1QNfKb0qysj+TlB6pz7AjgMOsdl9f0ShOiBimvOJh/8i
YKLOaxL5AfX3+dF3ZI0u8aEA2b8UCjsJWRI9Bh/+OxPVHZzJwNHpNyjTdfrgKg8L
gX9ueVJG4tQsOtk0UpnmvK7EwlYHYPZKJ8GyBhj9tNCAwwdTIRrGtLQno6LW7v2w
q+l6ner9IFTj3P+nuwchWOHVeRs5RRNKoz63/TOX/0hU6Zw0nXb/U/67XdJngfgh
N6n9zq3gI6YJjDF8R66WseOlROxeh88qiQfrfcR+NfJvxM3F+206syMe/F4VJV6X
0CYWikQB+aRqKoh7E6iDYjuybPRVd7JwJerHFZkiV4kd9tUBAsat4TI8Hn2el5xZ
RB4UsN3jeU1fwGMCYln/JA4lWSeAU6L/GOmrSj5MgXu1Wrl1LW9KZH8/7mWZ5kVR
HGa0ISF2v0kK9yAnn2hdSZ5z2ckausOoTcwfnMNoHi0LGLYpzcexGxtmYc3udKsS
`protect END_PROTECTED
