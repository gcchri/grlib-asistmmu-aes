`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
byNnWh/q3qvFencyn3dy1f/XBV7rY5/Y46009YUDc4HFJsy3NfUeqduhQetC2CAs
NLiYgt/Lsxg+U74/ms+y2xw3+0j4ppigSDoJb5pbs5oyIxslSm/7+s0bM4J16UPW
X2tcGLztsGhs2gFFlmR3AvHZq4dvrRdWu5c50Ee/VTI9+3RMdMadC4veDwnb1JBO
La31vqsnZXiPXPpOc2whBz2lp6mGVHQDqBoEP2q4u8ywUpnS9S5eb4l2sQh4V4mU
KWEYIFX1ywAzSr0WZikLDjp7I9rhn/5+h+f1aJS33WwRUVyWjF3ZanRoaXyVhnBb
Jgk3BP+pHMYRQyMPoZfxJA54tPpRZ/PFxkwxIun4e8X9kk+YYqvJwUTKCtUKPbIO
`protect END_PROTECTED
