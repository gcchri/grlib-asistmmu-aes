`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EElRvKuFCm8aEUzjQWrbsXuLEPCG3RVt0uzRwU6MdQE425YNm6GzN/ZKixHCmdp9
BMNOLVkDjhDoBIRDNYyhXQhQhUps/HFxRo63vB0bHKfSBYRmupPgTKc5OCtnJwAd
Q227iZMuQPERQsac8+gMboi25en3SyE7Pl7cluRqyI4ANx9E1OXeBoXnPC0N74h9
3RSfKYm2ZNhRbRMNDSjXB7KHoWlypdMRTqi3fhTPy48bAc12d4G93AP19o+qw5Uv
K9OGlCxEw2uk2N63uxZ8yw==
`protect END_PROTECTED
