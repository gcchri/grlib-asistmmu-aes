`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tPobvKL7lrFccz95q33+b18cyzYyDzKuYgySa+KO/6gmCwNyI87Js7psZUP79yhO
N8OGdDc6A2VwDEsYKqYTvKN0Bo2/6ULcG2MgZClv40Sl9gMcakq245+Wc7crMaio
Jlhkh7mnK5UNShpcHgPjsf4fNQ+W99DyspmwAeZQMq8qKRmI/nHgTvlsmz2Xpox7
0V6iK9prDcIF1n5nDBRes2A+omfcl3ikENb4bVUELryo12SBMtoYP1INdI05SuxK
pnRnEZytNFKUq8g1o9djl9e2sj8dmR70BU8EHQ/kUckegQwTf5Oe/8zvqA4D1B+L
1pWYexQiA9rfPf9N1QLZgH3suwMgePccaXVRo6Mz9z1bz5ZAS2LoseFRS94dvXDI
GVrJ8VJv+zAHieS/nQs0jcECU3eA2/QylyzDbKVqAxN+SqdFXUJoQ/7yIPo45XXr
egwkId5in+PY05bGmA2tsjx4yBEa3QHsBGuxRwagyTc9mpzF2M0gTHU7v4Eu+h/J
CpnKPs72WXjAWjGj/lO9GMkTWVKT9TmkzUV5jJVwYj7vqiB2hVHLQUNNToVsz2Ab
utQJE++PpUZDc+cIoMaQ6ioaAP9Fx3UVg80nkmsoWodc/N9wkwk2PZa2lPg3gRl6
WI6a6NOCFGJEGAnLlR3LEtk0py9EupKWap8NKxa7DeZyG4ayCimhylktX5quHsx1
UPma9SWAk3wW4Aud7o9F7crBU5vtqFqex7cIZ19pDjPvgYO+j1ioTzVTYlJI0kPA
s7EjRIfNh0BZj1ALhz3/4Hj3OK0rEIBicC4pUdSWmqUEXVXWP6r7zsq1RLFDw8KS
ZqiX5W5oPfW4s32DSmfk7Q==
`protect END_PROTECTED
