`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mSEvuD7VCPo5J2wJ448tUkp+h0GaG8on9IaNB8+4+LCYmCnpSwJ9wDLjFrF4bKI5
kWED2Yxw4sPILzJYu/E7PZdIXmDnNqtGmlMge8IN2pHmKgiHd1JDXEgCJE629mSV
pwlyrgtUqTCKB5OvUsLP89l18F7DyOuseQYoblZIhioBbDV1whxivB3SJbOXfbhk
fTkMYOcVFtoRnp2e8yU91ePByMciGkzZZ+acD8n5n4P6Vhi0sdCghI9fvd6GPXfT
n4MtRc5uUeyoFXFYi6sactf3ntIh03krLRgCB4mpW9B6qVp0tBQOqghzzPj8K2Dx
EWqvYzwCrFH8YgxlKLgQiavNp0fBcerY4cSMboyrCN6DWjwlJeUacmDYSR0Fffjv
vehPiwJ3YFO6NfhnRvao8/8XFaP6V/L97B6Jui6IoXp6Ud9bvILVwZ2RL+SJocy+
oi9M4yZ2ZmTsWeTUqxqsDAI2az7PY1KwMZyqFPu7bU+HbKDWnccEOBYFJTMoKNmH
iLYalHsNQ9M/bmVMznUw08dZbQNMJxQ4c7h9WaxRdno5y+7MKeZpF76nK8rSFLCg
ZCn9CcCNVptnsB3qT3n8UlMbDV1BZ40LhNGvj74cjeVf7QCOeYoZ0cO4mMcnQDhL
hv40AFVzc5wpYdB1WRAaE7fH64gmEvhmsYUgRxNbcvA=
`protect END_PROTECTED
