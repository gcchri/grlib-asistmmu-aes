`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LC4r1RYvTQRwYsU7hLQUU2EIOcG38FuudmBUCuXskb4+oo07CsqKG45X+Zusz4cv
Av96Z0dLAECK1oa5/yKCRv+V/COwycXVvjZ5Mb133AK2BSx2Xsak1TyQHAIKOCV9
24tgdBmvsLt0IIjw2w/RGaljhTx/+2xERC67qPkaO4SGIidBayO+oVZ/nei/GlBR
9XPVoarTVdu3COI7Rn47LIHPa7nlhHuXUjrpD6OdmHFpa00cbucz1FLVDvsBZsRf
6CWkKKeJ18ThQdvXjFDCenErHOY8HRYQPtrsctjf10nSrA6Ni4iNXr6CmifQJhNe
b1Wu2qJsXL8Hz49664Wk8TkrNzkYaK7mNEqn9An5vCgDc0DHYKmqd4etFQ4s6wPk
Fmgr9tmHZcfysk8mA/Ph8wbbDIDxy5/N9pwAkC9AaLiWD/P54sKuOU8NBFzHsZM2
aFVRIyMycKxYRCOR+wi9NdcFRT3hf8UkJYvhvhc8/xWLTWu+Yq34CVtvSaiyZsbR
vJYgQwrPqrIaBJ3Wwah/B52rwbXaK3bTPx/V8hP6lKu3J2DoBZE3rb+QOptIgcqr
4Yzw7O9wATFAjzFB9s0WRZSzEw9hZEPbhS7aLIxAEIjXaQNpIOn8RIwScp4T0Op7
NPqy6fcrVFA573HAlshglxmbOQ0Z/nrW7baHPmzxQdZRgLALbjgwbDA8aaHKLL1T
+HlWIUYJO4Z4K6n68A7p/yFzOdkhQsREcnX7Do9Nt4DMerY/DvjNXV8kU0Bz+Ave
Wm4ZlOwjyEsK21y4C4EXLdrt5QmgMP4OlLREDmaBCoY7kwEA6T0voiYVnDlPfouz
Gx470yscBIngzaq+mAGwqNpZISvVwmDLVxRRFZWIoC/a0ycwO/oxv7Wsmyr40zuL
NHpKrdKslHSareElBBkiDQb2fXhvOuf/2tEIw93D4vXk5W8nc5le695urMAkDyVY
/cQ76KXx7BYqsuBP/i5l2rAk77ZpyiMGGBRY66Uo/t2JEIaqOaGyGQerOYqD0myo
Gu1oPqZDZGXsCTa1NY88XdTt1VATFu0PBflSC5vMhloE2yJWX+xGk5d+V1rdhQO1
nF75YE6IwHi5A4nV6yC08tcRgEw4Weqy20HElgqXoPXTXW+aWIKCEHo57p98Ym+y
tSSHdeI/RaqYkGkm55Tglv4mXcx6lkud3nruTO+ylWKGMyluy6PtlUJg+XoEM9FX
A95bsbQHRop3ZSKBpqVprXvrukV9KI0s4LMrSs1vbl/iruQIpyAbfWy/1TRo7FfJ
fG55rMIOMkgOUUiSGAzGOkTA2MUOGTyo5K7kFK0BL4HQCsp6AtAhycbmEaTlhaT/
gMxSkqJphjYSmEYaL7ArkkTT3mkdqDsYB2aO4QNR5IHkWt4t5yn7MXf+SBGVbAv8
4Ze5L92SlXJHB1lpjNo0QfFmfZtVbzSX7sS9WhRcWk26pyw1eHDIgp9Qu075KLUE
Q/e7sQmi1tCYTUw1fIpmBYBJRI++RmCw/gncns3gNxzn5+Wr4QcXwDjqQBT1yHEL
dVST6NLD+WutMvrkJDTPZKk64gUyPUsRVhX5OG8PkeHZCGa7NIFQLRGW5LiVkDRg
W3tYBcVh6ptIemKksqkVr55N3oW5LYKfEQ1PFXkpEk3lVcKkc2ny/3r9R0mxEc5R
GLBGNQ4VprcUm266BpUcVsOVUhmOo7f1vKqmhJl6qVMQZzzhbvTGxsY53CG9FVJG
AYMsv815jfuNWw06i5XH/0WlV/WVNZSw5UkEbuzaC0XyA9CH9tJVO1+2D/LgCnL6
ZeIwdLANsL1j9IZfFIKZH+1ytqDd0Gmo+BKyutzer6GS7Fz7M6f3LS0qx6iK4zkh
BKoieUp6VDVZZPVAf3r68oNDmo7EbfjK5ir46RIQvj43/SMXDbL0Dyz1Y9IS/Vif
VwAwUu0cgKyxADxVJJudwcwiE/w4vUc1PJbCDF8sKp9MU7ieBIABMLcf8d/XSuH6
rs3zJLQUakcNi0ammcX31YAgy4u9DWitNxLRE5Pu/cOPov5z/I9LwWJ+SyRmMAWP
20HhuW6+MQds5DrkcQTgHv4zn5kCuraTaO9F2yjntpAQKX5gTeGCANAMcBfq/blH
`protect END_PROTECTED
