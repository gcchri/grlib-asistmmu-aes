`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2oVwkGIWUT8KEEwTx3u7fCz1mLHjzZihU21JRa/ZnEbIQNY5AHNOaPbTuTPfhUqs
L1X9Lsk8PyE5EloZ4KAczV0m66R5UEzoF2asLeAaKLxCbK1QomxSPlUkhU88gVF1
8MxF5YsHVbqTHnUuhspVLgCle+gHiLoWTUjfiXiil6syCSO6eDv5SjCAdrJ6a+fe
RWPEopeCC9MX7V7XGTyZsIhDATNzThCNJlB8KJROqwQWjoPwGz6fq4khNhhpx3iJ
48nKzgdkBPidKLhrVMhSr27V+0XtzrPhiROQnxvbWsoCg4sLNlGOHW01tLVH9kSN
/QUl2u0sJI0mOI3L7LwfI4uGhXt625+PT2dmMU76RTKNfX8XIZBZtm9HCgAByQQJ
6VFu10wL6ga4X+rRYenfUgdphoO7bz7Ew66wS9tF+q1ZIkxlGy63eKxX5VRp3WkD
sFbU624NJpAGkBDK6nIviDhmvs2H3b//sJZRCdT8FRgJCtzPyQNBKr73DlEPNmHI
I22NMDyPme5/v+O3PeTnt7KNtu17oGk7kUFmIpKt9Nj2s83+m3+1ajiN6Oj8EikV
sBtFI1m79RPVuC+uwLPs6i+HLFUrby24W2I17TjAv/cWpe+/MdMZWAOmyQtzKy8g
uP2YUHYzI4AbZiB3VOUpkQ==
`protect END_PROTECTED
