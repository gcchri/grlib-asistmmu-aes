`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sZFZY0z3qGz5DXWcP0aLGOg7i29gwuXbXS+8OcDiKzpqWzxUnStC58i/J4Yay83t
J3VSeB3U1FTCUxQLZKKvFuoPOxLSIlXERwMGZqoOuqDy6JUBjEhKbm8qvwu+iNeD
N033WRFI9y6klV+rviG38Ml+20xFC7vpEmXC431dBd6jz/WkXPLe66tq2ewvCYTj
ha8dUTK23eVjaIuXREFc18UB78y5JYowc62Cu9MxYGwZ69IBrjW1KT382+GrqFxW
4SBK0WbqdnzhmoT8IBx37Bj7lql96irX0KXR4pPfDQ+bXxVAWuAB7SVrKk4h7WUC
D1uYk2J4hIaFZOvMDB93AxclSig9bv3yer3czjvhG1Y5WjUUiuI+7NKh5ySwGvgM
jJyt14ZKxJzbq8sK+Bh9zFDNr3NQ1FgVHuCg7fl3zhk=
`protect END_PROTECTED
