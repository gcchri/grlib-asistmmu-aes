`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cb7DiXKyDYNP0sxILp4eR0epjRWbuSHIHEbl/A29Wp6eU1tW956cdSPSsq93X8VK
CajMKhr6yBD3jnnBBkWz0vcUR8B4hu7x1tNFTHZrF/4YGLQ3l0LXM0zjCnYd8N8G
/b2My5nCgWD6mSmphYSXWSi1c9eqWx1Lp02jjWeMw1pAmf5OVYIjvxkV0+hTL3xr
Bu/6o7qMSo32KnsD521+1CJq9hCbxzQkU7vEX1dbRT4MNbWG4Zce2YAVoJBSgAIq
nMybZfDXNsUdXTA17H8ifKGi7oKOriJ3wGqbMclHiJdUqJa8mO7mCTZRydK68hxZ
2vZfxPGe1CuFqb0BfBX+F9BCwVNjGzTIyEC/5DtuQ69N83ephOONq02bLzJbFscQ
7mvOgJHOdGX/cewkOEousM+VVhFwOhjN6n9Kish+TE3eHdFLvi9G3CNyqjtmpkQ2
NrZiUw23l+i20bhXTDnMhjz+lZryRY8MZOA7PTtL4De3wdSWiRaDfWQiUG+NS8iW
WVbQVF8fcSS0oU3sm60Iw/fkMs+UPuOaoXnI93y8obeX3tqRX0eYNiSMSdrr/Loh
5HxwfWWnH5m2uuBoBxFzMzkj9DoF8QH0wnJZJ/gfLr28D35HoGzJ5HxpGAtcOdlN
yXuEulRFyItdAU9jQe2omi610DZIxQ4d8xC/tClHh10MClFOIHFsp3Kd0DNAGABf
Vu4w9Udxl8PDnQd6LAzHgQt4DgWwkYnOMhHlKYyow0JuFz+LrxAMPcJwfDSEdl/u
jx1WcJnE8r2GLUZcoMx80sNXaCnHg06jS5McJgATTWOiCNzoJaRt6XhCW54yhGXC
Z6Fb821Fr33tq6lH2x/gHZI7tNCNqENmS7Pxgwzoj9Rp1SN/QHPlY6En0PLhcKbU
c5dfP01UbUx4j/J9g/vH7sEEHcX3KHV9hYgDjGOxUzD3dyWpu9clUn7J7ZbZfPEm
eyDizUKy3R7x8jqYOVF/ZjBvj396SZozSsCYsgDI+ZKOtkQFBLLtbH/HNt5vrd4Z
c70GA05bk0tDcO3kd7YKC6d505W8yGEh0A71Iax5X1oHgJh381mJ6E8mdSQuKt8n
dQ3ct7w4XtgbPUwCD18MAuASpQgs8dKp/0kpo63DdPF4riatyk6q0W4dkQpiOdVn
1oLKu76hxzv3V0RgpKZmPmQroUnm6IHBi+BjCoIGIpQzIY2dJmMcneBL6j+xsXxk
8euiaiW+YPXJ98sH1b/9teokcFjcWX3EAnAQN5DPicINA/jWRHgq3029bdyQhyal
G/wEmp3woNZOWiITOP3B5M0lzBYoX9feylgU8XJL4Qi/5vH018/vQia3G7jSLRUg
7dqGRu897Qu4DBBZG5fJcFtoyJi+l4yCgWHsNki/9PuU6YAMtngvVEpHShA8pkdY
YEpKiooV6ndVCZg0469IRSFKhmEk0LtW8SeVN3hx8XJvIPzVma//R+JCUqOrKb6F
GDSeY76lUEWHRZPjyHHKakqaE6/3KHYihPYGLEkhQKcVndBpN+WNa3yT6M7E702d
e8W5yx6CuBIs5Mpf45TujXOO3RHbSbUvgcU/Qqkxgkc6kvwysdNiiEa3dMzNXtn2
GMR4zuuv6IBG3o9Sub1cUSCuS8mjbaSDA+7Qra8sXmLl5xiiTZCFThVFc35sRL/S
vpC/sfLH4Q8dWGqGPgHfwAZOayGiGN6Mdd97Tl71xiLu3wAmMBfjjrT5Sjnht7U6
o0/xiGhzFdPTvRXJG4+3UjrSqGKeD9kpzqIA/zjkmsYFYU096wGLTw3c1K2YMfkj
rrpkKM1qeMnjv5us2UGA5oc464oY5yoP0AyWvg9dyTzTqvDh4w9v1A4qosAp2RT/
vXDU70nISpT8aJ1aSeVEEHnNJiue78wglQaSTilD1IttwEOcMJjffGjs+ZwxdvLE
68+w7EvEMCB1dfXNcPqnCt67SBmhP7qJsOvg13wu2m6wAkYUVRXXFu/M2lwzuGLW
HIQLrM8heHWUkR4ccazFaLgkAefGsNQd4LU+smcO5O92Bt57brG0QE0Qxdmmae0H
k0/43jawR9UPHOKZtgZMhB/jvs2NIKyz8+uZOaZMBzIOnGQS8PPMmmB/ANag97rc
JHOaMuSEB8nt4hMAlU84AHfF1VJC8n1OIlRd2ed+9Heydf2PwSh/cha1cSfDvXK4
c4vy/q0Z7T7PGnY4M8llZZ5X9slGAG3swXz47cheRg19WVyZH0vnK0f23Fy087Eg
vGslKMp3LtIh6XODbr/EhLytaZMQcQTUGfi4bRCTnk3e3AVKzz3vEt7/Bn3887/i
xbOWoKGwEYalawTccRQUczD3fC3hJriDrFXkOMtzZI4NAacBuOFYLMMIZgK2gRAm
diA3SPGpH4tH25VzxHYNDJAQYZpu+/l//ZAPq2VRCuI6F2low5L7K/u0eNfKeJRP
WWlpujUFYpthAOu54Y+VVJ5juMpJ9jTxps5iDAqWZtkMi2eE3T9N34sqEtQSiQJd
DkA6COvjouNpuQsJ5F09iQ/I4Umm8C7qCwccsCy3rfOd/ROFcQEiYJANvjmtYYej
IG6ZJx/EQJrDdYIglhqJJRN2FHwTveo7wiXfqKM6DYRLIf8Q8avIf66LYlLznR7n
NJoQF5lHWxiuISGKRR3T5vAQV0MinMHs6Gnb+dSYyJfXhr9jLOS326AwElWX0+26
Zb+hDvPPSaLlUEHyhMOS3qwAsHZQW4FIcS8QwCrPN278rzSoWMfblnsYqVeK/AH9
E9STWNzwDuxZJx4nsz6X4OTk74x1dhin08OJlvJeKKAp0/2A9fWml1m8PRfcZV4B
fz0Dz+cf53v8E6F0X9rCq9XH7DVjze2qS9zcqG1oOx60p/SkEl0U/i9pq+5CrYzc
+vv2W9RvP7uVT5L/gAKKVwlZgRHQNMC5XFtF8P++4jGBaGZgzfjVMzCjrWwKiAlq
5ZLti7vF6Dl6Jhb88OOdzvsLdF09UgvgMBUNScMd8VQUrPigYm7VbHC2EwD2zaNs
nQ2VwgQrHpdMhP2al6ruzQM5XGQLHxH3JvgyeuGSbC2Ee8B8ZmOKSK6PrQVYRyH5
XdIv8iJgA+ub6gelpA3WN7g84AuYS9juUFKRM1Vyaf8NrEqO7BmxAv2iJZm8qYsw
y1bUbFYjF7ltJgkt0AMAzFRMyocJl6E6JohkpxkJkf5aMVLHGC2kxKASR6ESx4Jp
j6CRkRdZX8XB9I3s0x2878Pj1ZNi9f5spwEdstDA7HgAw3VCff3OEK0Uur8A/jPy
BM3SRastVYWnKGYYyrfGzzuST38jS7R2wWg1iOJkOzRVK/kuXFB7H8SLeaHEFSrT
Ia6Rokic5mO1g65B7+XLGQ6g7Nlx8hBen6zJFbosKI04bX8DJuN1MLvhZY/kqPjO
bhpoNgfe+quyXRXRoEvdHCV5AjBrYLiJvCtJiVt7wb0SW4Tp8Yv9K2xidZTps6FG
+yuaMWnwqnVQINwqcIeeN/F1QVk3w0O4PmcFWLpjmWw4fqCf55gOEl+6WaHXRAep
rTX/gfoZNGBPcnXvyvlcLFavhNKIXPmetHnaS9NBVfncodV2F9NQg/47SaVgUY+e
eWxm/rdkqKtQR3Mr5azf9uz41Eq5uIF+xcyR1wNiKlX9QMBik96my8dG4WDqRVj7
rNHB2SEgRn6jBJQRLoHKRvhJOI+YgZwch+kdzVHuBXPRwZGOCYBhOHN6EZJy1muC
LT9SF3BRmJ+ilBuP6W3tJ9j8xZunrSM0FQiAlPv9pCTwf/xg6iJE3wLDWQ8CNMMd
dRH6dcEtyOZugbNEaqVgxLf00EpyjRvdrD4r6aeTY1AliE4YXLqT/OxchTQ3XQkk
1kkcZmw/7lz5wBPaYigVCw/lx2x84TEpySRsKSVHt1EOarcl3iRDrZuoNmUUM0x+
iI0Y50tODCOlaqj+hqhozsWZ+FXAvOngnzFeJbcj34msmuQ7C/Q+wehakOEyTyiH
Mj2mtNK6ig0xNeYXUEWNgdZue3eSYT+qkxBLMCiF6Om9d1WURR2iASP9gaLqtYTG
FDtPrhoNvRyT2FTI59yV2HTt+Ch1hB5HXG0c7HNBIgS+YxP9Sl61Xa8xzoRb0blu
Q2NEiuwqP/QNYGHobwMNfVA+5pzyF2QEf03bc2wTzrT0EhV4+VyzF8jK4MX5c9mT
juVRPuRyhot8600saPoX9L6lBF8fY/ObADXP/DIEiBwiN/LskviA1Y4P9Ejx4Ubp
Bu6FOiBMKJG5fx9w/xxxGDiAePjwoss5Vitn8IhHuSK1WcIqkR2hKGINthE2YaXb
fRKCEE9kD3e1abYbVGNhCDyQ3aSIf4NxxfIDWHB+UOgVXmOb16sK/UcbRcQJtbT5
EBJT3Brv3IBRvyGXdlPGqlxv/u+O2PIdrHFCXQCQCumdi3gF6MfDJrI08M51ibFI
JTFb0Kj3mWNaBrxoUnAZXKpUDr2c7PaSIP56NpWAi5iTsPkpzwk/LL+pFLLLMSap
kYx334DqdzBNcj/FKyWUvUXjfgz2hiCPIbOKiLw6RRx6B0SZlthUqJb+Bfe9cJMr
e9kxkj3IhV2WRYD3sLo0aSBk/UHGBf7gm6Z8C9P04h3u6uCnPH5LXhzjUdHIT0pX
Y5wxT4ABCrhxPofzEoP9YAVc/vD2i6lZv15jEi1wsXGCska2MHoI+/LDMzCUMcwc
hwSh8hYw7ykKPmlm2xjMxBvFONmIqLIzGNn7TyqBlja1rmrpcknh31iyKyRD6HRp
fbv+j9IJCHrE81SaewmGgahRLJK5cME2lzqBrcQB3eNXbe5glALBEF7J/fbAzhgK
E59aX+f+FQxDVDHUgLMkQdgpW3lalCBFfSSlwtFFmSC2j/JmQE2jnG1BvQ9V964C
BUxowFBHAb3qeeSAuNd3m728i5F0TY+I88BydD9cz9dq31XCDopr29NPP8ZKyNmy
MEmcqPjOsYF0l8iRHaU6DIDBLihMyLDE4dfd/mPTAbjEiLO60qvEMXJhEu33F3eb
BDsf2j16aYCnM1toan2s1ZvcEeACZ+vf1MEgZayBzE7vUtjfuCY9b7FgyfVeAmyi
uAd97E/mc9oH7Bh/5di8c063/xZpwerAtqoR8/Z2y1k6qrAKEgfsWmUyEns3wE1U
QwzFng9E9cFXzUlKp5NNvfiu4HA6Vy1RqF4YDHcf/yoQ2sq7T8gL9jcNFuRDx1R+
hOro0FbiDIr6pUGaiVoqVDUl6lDwHHCqKqOPpxEoQG+SFRl1AI4rcm16LX1YEs4v
rDXmjbewIX8iNLzGjsE5fr/tS1keu2NpZMp27uwrYpbSWkjGNszKcdZAQP14UlPB
GWwae3Xksn6kEgXEYT4+AtMHO6VT4I7KDX1SzxRNbPkTUoqqpkRV6OBV8QGRVEuF
c3LjPTRVLuxQJ7IXX72+12qFzVpXVEWYdxgBSZZOy7xhCosYpNlebTB60MGZgwg3
4VIHBLu8EGSja7H1rrMw0sZNJFUuHDjFqDy9YnUzNopeyR2H5QYsRjTGzCVJC6+7
x7l+++WPkSvRW6T614s/5X8h+Z2O4TrCTzkDKHUIpZq0M0l3csnLfFqpccnONgdW
vY6UxQ0BAyGPEU8ykJSvS7xXJvgfsGhVAeHoDkhSXhLHGk5WZLaL9kGe1Dtd2uQ+
FjT6rm4RxLRFTSDa2qZ8DUUzIqrl6JvQIFvFe1sq4Rx/IRIJQH+FAYi8/zGHWGLq
1Vr46MaWqtU1SUtx0DNblsfXQWizi+EizwDoZBJII2vEtIj69BERUuiEynHf87a5
IHEcLTE9NY9vkzQ+Nrpm8pla02+S4FOpPSI2o3SIz44moWhXQEXkVHPsYemVZRTp
KCXDNzOR2IhIor05uU3WO/uRRTwkrZAPIXgrohoIKO38jtDVMPp1eIz8aZbm0bm7
AwQhrqg/UakS+g34OEw19HwMZM774LOhtFYyZCQ7s8an6Es65KGbWhrpgNe9luQE
K5hlDj5CPz06SLyRBGzMynNPK87CAEZfkulg5u8AfGyGjVryBxEGT2XuVqxJ5hEo
Vl/efmoMMsbJxgkBQyoh8TO2p0v57RYiJ0+IxoK4WBP4zA6bDZt7fH3wgsXFMI5m
CevOE6nwKOsqcLhJTl00NReBQbclKzw17D7sUVYgLGYv+HTKfYfLRhxOhjTGpFJb
ijpbnvh7OnuobJyx8gT8cOMdZVck7FjL54fpZJV9rnvWqKZU5WfmlDtD4tuMrGGA
zoJRIAjtA9BUpt6tk93yMAjinU3EmmrBg8SsuMY3FH4C8h0rq/v92cnwHsZJ3Fgg
xIUPPkAVBpzxGMWfKBfFj0dXsU9knARc+veN9171xU3h3qG+UiFyuZxAhffJ/Umc
D7GLOkXRYagRBb82a1omgjLjoS1mU9HKEK7py+msRusq7h1ub1AGx3hrYfmpucF8
Bot1HelqG7Aa3wOlKbaia2VV93tjU/4f7ILINSafc+/maHsB7slJZZ/4nPDtvnVu
FvUS1dr2J8SekSwnUPP2jCO6iqCX3RAGxLg0JyfdNmL7PCQ3fm2e1O3QOWVGUCEO
Ax9rBSAZfs1tq447nMMGfd5sep/YrwY+iJUiWXGM/sXn7WUm7hhz/fAD9oMzZlmb
GZSsWuXWtsV0m3gwVc8d4ZD0UDqesMp46xwjRCuD16Vo0jOkKny3JjHhsIYRwNXC
I+EQMZ4f9C77R4oQ6wbNue61hyWJ/V6QW3n9X1KkRt+yzhfFcVkS1l2AwJaXu88O
oc1oyxGhRwwzRz9akLmcCSLg8+41NJOk9iJkB0bYgdEEAGEpmHa1HvspxCafUsKQ
tqCr4hfvDG+oruSWDgN/9iuIU2Gw0lCqiULAgMWWnn9LB0aIHOIVtEzkjzMQ6bY9
vuC2iNjyxvh8bUOdgfULAM+4wkYx7X0t229YFJCh3HK4u+etMvkJ3wO7Py8+lN7z
8oBNGAioWh+HraI0OpbUiZLMDzE51hwIWiRaGJIBVMTlIXtnyRqe23lBKEL8AAvJ
YO9NWYyGrqU7KGo0XWRt/8+Kb5ImXRDegiQvx9T/M6G3cBZdMAchkShmO7wQvpJH
z/980ubE1OJk6A8Q1fLRrv/R9oEh3U3AiZzj0RuMbwaM8LMVD57NrlYidP1BVJwF
rvqLj0pdN5xePI6MTHx0eJBSnB3EjheF1w0OGfv6/804r5pPHFGaDWn8yziLcYpY
x7YFRc6VzWpi1tf5tphoIjwANMmgs6nOcYAlsXmMljJI8mB5zNkX6tcbCikse874
CVR/F5pEN+Ar1xBs5CSU0BTxht5dwl5DUulEdf0nFqEYtQFnGH//1EEvkMYOaMYf
8L8WNZoC+w4W3lQ21+SJ0FEdYSvCw1x+SYQOtXyy2rV3lov74+STcAbFLEeIqS4a
KMqKy7mPehAUOoHMQseHQf75cXhNb4a/GroAA1OENEFIBP2tUB5f7CPEhkNRpsBa
am2YYc86MUQw5Ewqj4wjfgpPrz/4HRc6yUZLnIX5qI1xmuP2sN5hI8AYzg+DKu5i
aHxhAqb/rqhfpeTSmduzdeg30RxrRA8yJeIQuAaKErQWQuWnic9Il/EU4XIUoTLh
EI0Cyht1Hi+12+lVqECZsIrbpZYjrT/owO7LYLupoFQSOJbthMQZM5qDhEv/hq4p
z1aCcCMsHAY/COYSXFjgrapLEzySjQRLZ1hSu8ZrINzGAadssIhgIPsq/AtxyNa7
1rd8Wh86+fgBwgl16J1/0+q2f35d9exbakqiPz/lqJqMUMeg351ilRCHIaizucMN
j20l6x/ZhCZ5wZHacOLO7mc9+TJ8SZtHmIqg+hJ/XpGhxk7rbgMRcbVuTcrjlv6I
pGRl8zIDV/Yes9RmzH09Iw==
`protect END_PROTECTED
