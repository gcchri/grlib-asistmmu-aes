`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B8AgfneZXKDjQRNBjfb8vC9Rsn60gyLcWwo6oSTV1fTQuJV40/Ay75JD1Fjhq/dW
R0o1o4tOfswWuwH5+JIOj23ogozd+GDpDyg0GPrpOM88ldfcgJIzd7WHIw2TlEUO
2Q01wOlCdaTrtRvpms1iEAxUSKcIBgkUejBvuRQh1A2vcRI0TzK+9+94ZM+9ucmH
vuhRvb4ilHf03vQu3XYp3eiDj1K4mVHX6iDN/gii24TEBkJGko+9t2BN3WgvETD3
arTBDe8tOhh5Y56oX9b/+AVKHf71dxE4VFWgi66UGbKIJpXcIC5xwc9IEtF2RKfF
cF4G0HTWVqef5gIJcb89kA9gc0v70CxC2hF/o3aXEr4XTghowm1Xp9My92/LifK5
RutUav9003v69T71D6bQMTfHqag4fDgtWrQRIKQPLHWFWKX+HI3ZB3TwQZ7r8U+V
XoEkxLjpCFslJy9HOz4FCTRKCJC//RrozczxuxHBirdO8lPY7hVu52/bOIRkuopb
ELc5KuI6IO+Gm6l43KBkg7Onb7Q1YUowndXCkUvpauVFtNE3KzBQA6iQ7WOzfy/h
vzdyahjT69SaykllQ206PPZdLScuccXdtkuqWAw/WZgOfnh3Qw9zL7b5HxjWrhFj
UgfIuEughRVsAkb/u2FOBg==
`protect END_PROTECTED
