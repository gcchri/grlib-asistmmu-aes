`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSD1BKgtaPzMoBlidqoc/DNqEKZMVg5mbFz5HLHn3QXqk9hYgDw8RUWb+W/EvVCb
6nDo0bbGtdSlk65H/FDRUxhVxhB0D7DUbSazePJM4XYoF5J1LV+8VgVnWBvaRlwH
J6a9wcqO5EjGm5f/579vfQ/LYCtPIjHcCJjiDlNGoR8Fru0NdZS4FB1s/SvbasPG
LLHYCzEamyYjnpemL0ysgNXnOnCCj3w5RcOPQbdWJ4+ERjCfoWjsvSk7PxXCkmsw
JUC6aST6tMBQW1ayWdzQIxtjhpzzNWKG9PiDNhPA0lnZ/nFNQeXxa5j2Vpxb040b
UOR2t/mVDDFn8ingqDbP5yAoKTSZFPSeDbJsKvc6m2YiEquXv4Mxyqz0D22jFfWc
v2EtzXwCRJzkAk6w2TqTvVDIipTzAtDrU8T3AhdQM4JN+vz4vw8IYEzDixZfcgX6
fxMNYmY9zugW5FGy/C5Sgdic0JRT3TAgtd2j7tZjlPOK1CCq3CQlA3XMrvf9dAl6
bZiABqb1zd4w2adn+9ua/oXdWSw4O3FuIW6miqwyYHPV4pgqCOHM6Uuok+1zVuGV
DcjtkS2/nmxc4VeQe/tlsb4AGR5wPKxQY4LNUvRrc7j6XMy7B8KNPH/pAzwcHnxT
2a/4KuA0mm/TaAaYM+3d9woEFD+hhehlnxFpjqW8nGo=
`protect END_PROTECTED
