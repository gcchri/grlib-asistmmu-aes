`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nbQ8IXne4WjpLf8qe1JzoMIlGemLlmNLLYWvLkYZQ5Vreaa/pHCge3bQ2hV9vkZC
vPWlc4KIkm54B6gTYXEIGoyzvbM7WD7/1vJuti7WTBXXuAEU2ZVsyLopRwVGIzZW
tU9hw/Vo2TljwCF87odAKPlLLZMTcL4pbHUA98HUGNGbgnenklByHPCwnD66yBtY
qGMsmqbtozdy83IWoc6NFvCnlAzWxpqnmcMCJP1btXBv1qfVmYggXxM9vbl0zSI4
hInlJjdqPqLSzEHFWx8fgQ==
`protect END_PROTECTED
