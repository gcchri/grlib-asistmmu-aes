`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neiwBgVKxX6vrnobmpmANmI4AyeAv8DmYE9x+Nt+EqncljONYx8nyaQfyFWOThRj
drJohHa2V0vBJOH/0Og8MdZSKkHX9HKnQV98SWkPZUDWUz36qlTliLZ0AB4FyhA9
DLJWURkD2LNgUCIzbe5FP1F49BhlVWxMIbHCyoG76aSPLs3+dZp9Ewgb7PnC/i47
lMkD8QxmUzv+l+GHzch3GhmRBHX2fhCrKbmQWQBcOMh7gFAECCX1WnJ341SBne/+
qZDn9OB7wK/B/nGzNLxzT5+TCwLhptaYoLmZVUFFSEz2XuJSQ6G3EN/p+iuWLB91
uDt2fow/2dwURDWzc4+Z2kEfEpDglatqKAPDz/s7+9pYKoL5dVbd+ZbkEMKdYz8C
O/uHuN66QGoRIXSuZiChSYwwDwNmWEyX7AiofgDwWcHFLj1wDoBDP5KydiLw37EO
QuV3Aa01/HcJrLNJZzItwMyFKWfk7hb4e5YK2d9cSSg=
`protect END_PROTECTED
