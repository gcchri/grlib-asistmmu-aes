`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKekdTP1B1V3A1BCmDzPwsdd80o7652/081vVGePQxFcuwWi5f0Dn6YRKILIGh0c
O+cqO8Vc13Gy/wn+c7HY2Aq0rc1WWiFAAeUNxlCvAHnD5DK90kGehkDN3cgxKmJe
ZWn/LfcwJYEoE771jZzh6MMDIM9f9LRSZmZCCT168Iw1ZVQMb0rZuZ6+kP9tuT0X
rDkO5AQAVZ+u/qAlkaJphGTS49jY4CL9aU6kp4AmdeYGas6xkWpFQwsP84LPBxyS
`protect END_PROTECTED
