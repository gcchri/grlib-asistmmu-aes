`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1n+wnEoL2pfe4swtYjC2GQdG8SyfVFUNdirHY2uPXCAjjhFnwPdTn2lntANt7Tw
EqhlfjxSaarUQpvxx6QzlgordCi4APS66rsWnJHoYa18gMBGFBlBF/CuzWh2xjr5
tMsC9Mwi9SCFp+AMaVV+mabjQM1VqJIgd4arQhr3D6Fe3CfovTvHFWkeFwcRS3JU
IA5bPo82RAkvUyAFFxgAIg5G8XBp8hzsjF78X/DdjQSOWHUBM7u9HZ6LkQxWZXHb
`protect END_PROTECTED
