`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6tj/IBCZADQ4GwQMJlcEgekvVehpzb+CKXlyB0dBqbCZpxTwned+iOyhGZHrAjF
y0p813iAVYD5TdfBqlOMPlX8DsNGEB1/RJxhLPAghTQnb93Eo4Y8ITAcRbYk+3Ku
bqD35VHCxpmFJqQktvnH0g5RHh6av5SblXu219udTT5njtVrMNxgWTr0wULRqYlK
IBD4VRPESqf9ntUksAbXZKBBVgXLYFfQS0tSJir/VK+5XArOG/8jKXM+9T/LCi9D
csqFgCzjlEqVy2LeGR9X++IzBfjvp3mudegqSIVVQmuAkNv/E6fZSxaWUfr6fovt
QzeJeq1P+VpbBsg6lCLZX00PBi39wigQhljsuKQvwKfkMD8uWWO5tG89A0auXZVX
14o7P1RHNsCM9bnUDYx4ynp3vDFYoEDlVSttHBdgmHloAhjCpySVMJ30sRW1Lbz2
JZHmKGj11XuO72z+x5lWRufu7eBc5A7W80hFz1978JJ2zeHh3d7Gnec10oHt/K1k
+r/MvHj3nAo7shTk4m+S8SNaP8mDyGEXJIe/XX8prgGaxUPpC/FaOXdp09esEbPR
KpCqSg+wW55t5A8c4SXd+eiw07VgPzf+AbSq3/KFpR6PRjJSojbcSIrnENEJdOjB
hazr2hMxm6bpU/AJRotrGLs/T7xzW68CyCpBdb7pSyh8h8sN4K+AR3MPnJZBsKnC
hQ8uem0V0UVCWb9OR/WZLZhB96nBXcRjBzDcLsA9NOk4XfKwnAUQP95U9C+nUD8o
gvCq/3hZ5O4ie4G99DH+sL0X9GMQgwnVCsyqQlJAf88ntpRwvlLee/vwKlcawont
0lkb2WSXZmLcVpTfBHcy4jDpBKSaooa2cVsoaP/WCaZdLncphfXsxc3CPwHlrUZ7
9VKORIBA8BwJ4of7YctOBbX7cLaddZON/eHBJCcDBfhrzsYe4dyrNYX0VRtTjo0v
WI0ljCswBPKGMc+SZ5gojWX9girqCJEhq/UQgbB/j71rCiY0XwR8wBte0j5bzmMp
zc6BRTYkuW4X7uJ3ZSbcmOE2/yZv/OGpelUJ1X/Ko8X7Iuj3ToBjCsx0PtqDGCJr
TzOOJ0Ys8Dv8tfmpeOHAoh7TcXQ7fPj+svE+v+NGsBe+mrzgOSpvvARglX9UKVS1
Yt37nb/A9Zn7wabRkOQfZ8S0l9LoktDGcbygc3kmc3WDZuiVuV5amZfdY4gN4qqE
Bx30uQG09ZzpX8nhF375x7jvXNHYlL/erdn8wTiNB+PMwJNONbgr1VmDDhNyrqA3
L1Kchpx4P1GqaEf1sr1kBecaNWtrn5o2EP2o9+A4DKPim5X7Ot8lIVhMnlaqs5gV
UAEIamsC34pAshfP0eqtpQ==
`protect END_PROTECTED
