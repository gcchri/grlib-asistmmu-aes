`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fJFKyLTwvhwIAogd7U8tZBYwht/3K1EY0R3DEb82GwUlf7tJgZJhEp8vxRU7rTBA
Im356FCMvFdi2XEgZvLCXS9evxh9ak3wrgFxlKXuBNrXWEObbCyY5pv+1WVZiojW
yZb69GoZa1z9zqpa+ri4W6dO5+qcTBBvg50xTA//LoKTNKw+I+etGArmW1fOv6QG
uShGGoq02Uzak1PpOoPfCCvz8S7tUo6Vgb4Az5hi8Dmt46S9svvx0RRE9ipcp4F4
3Fil6HrYzoOwJXz4at+JtKLzGXWEaglVozYLx0Bh5pgRJNcPyyg2F9MTtojeK9YS
9q+qJpCIwRqFgrM8kdvScv0O/wtjznWc5ObQf+E/rVhero9HkhrMwH1D9dcotM15
avuelPbzE2ro0fRO1XSqhvOJAtR+uYbOpNMLiOaSX3Ot2VWhaPrissiixSUbL9ft
0vU4eOjPdRuVYhw16Hx3XAbBj0l0bYTmZSJ3yWoGbAc0RgcPyehhlPPVvwVA12rH
Qs/29969JL2R/1zMzGsopOfSiZCT8isQXBV+FmncdpR/n3EpzAtYihTvThIQ/HY1
M0To2K6iRFCZTAvaZ/BKJ5lf8YxxFEnhstb10A3NYhgoSvFv+vOjVx1RQw7/fNt9
SJKMmf+PifrKOpGzho2xDXKKBNxa0q6ofAu8FTh91lKkS8jCmuIoxIV1MRapeGlk
eo8ArPEf1mu068trY2fYkS03gtH4G9/tOBkHZTyxnp0=
`protect END_PROTECTED
