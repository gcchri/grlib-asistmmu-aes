`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6JsA0U69uZtbLl0FBC6IbL3oamShAyy9gq55TrWcoMOusj7IWP5zypY0uMKCfQWL
w3WxLx+FtR4ariR6/SBuBYAoSRj6Vi253iNPMY6+EVXHdTvC6mtgMuuw/LCvj/Pb
1udTZWLtuZAgF864+bR9XHArAuDN1/rksrg95T9Ejj+3xshlJRp+v4q1aKKfT4Xu
bbz2AeKRLhxc/Rox39NC4MBNaLemz9TYfFVgZMXiJWl+VvF3LFtEhiY7jlCkFiep
RIeDUTlLigWnpJ098hqvX47W+5EheJShWUDnzdYxsZ1N2OjH8j3ToW1bCv6DOlJ8
h8sVqCSja+Me+/KxhKTIpM42XxEYTHTJVJVJ+x1k+gPUuPZFl9oenI/vvQjGTgZm
6OC8BB9P4j2koOS7LK3j8Q==
`protect END_PROTECTED
