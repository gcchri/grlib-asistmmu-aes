`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zy1fXNyrtjLa7RFk9b4e3fJjQ+yI5wuABzqt6LP4xy2TmbmIDktx8sbHojrLH4TJ
AvlF6Uq0kToSS1dv+GcDUrj1DcRQ2yhrTc5q00BbAvC9oAI038Wa/g+uHyYUo66S
hs1G3t3KHCW/hftQkr8Orx611zCSDIGBOetbLXeNsejwik62S3YkrftR9v1UlVPd
HSel5lY8P5uR6nJd4mksRvOXJAt2KqQhNv1HZmJOAC84KcKL5bdi5+u7Y+gaiYhU
yEIplzFVrahRlliwu98mE6qE2Czb/6acH7kDzSgn5iX68KTjXR6JsRVwLxZl9tyV
`protect END_PROTECTED
