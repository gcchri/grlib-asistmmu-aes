`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3aZQ6PkN0uc6LChYkVjEuXW5SkLP4Sz2OmoVdUeoDOrUfBZ17a6udPm+GjGGK1d8
eXiWf39+6Gwx9jdHCzFaru7tQQIm+zHJnTpKd1J6CffYoTMzgoHeyIMfxuHMiKpC
dhw+2avqCqNRQ1wfnx5s9+kxW7WZiclcDAse/lJPlV3X/H3JW0fF3ima8qycGcLa
t5iIsGisZkwHE6AwdSGnOkBvDI3TKE37YRBWAeiTSgCz7v3fxtqb4rDu0JO9vAU2
8I0A/6QE7dtncf3IcVWleOUEBl/IbzGtRSaMyH3qJLp/Z/rqeOm/Hkq4PYAtD5Ab
Nvr8MjaodNg1IdOKXbIJ5qVR/pli6PM6CkvIczDAAykMOWJRlubrVPyGMaYzhCs2
3vaBYFJUV51gyc9J96C4Qm+IM9YvnqgfDsoE4aHIv3v+Pmm8jKaqbBB3TFCCHCWv
7dMdZN0wwr3BMD0Q7xIGZjferbOOHzMFMNHzZM18qs06TfWMHj3sNh2SyJMv6LQv
G6HLfkGgLGgE0ZWyY3RhN+0UEw92nf7mhJQ4YhvWzlnoOymulWVQw5AhhcD+EJ3W
yuxGgqX1W/gZRkpj687DXrcLA2Z4t6uR+Tg4UHeW9+RgxcNYVGZQ3wI0KiBlmigI
o+wOqQznHgp/r5I1Jes/gN8HOzTMUdHTn6nEdxuquVClFjryukH1rti/tiM6v3IO
a7cXeMp9E8Pmq7GL9kafXVXRZ51a7V82Vaci+mVWM6eq9vZQezdiuq+Or50M++0o
EBbRKy2q54DgjB+NMGSFvsV8E6jzeB+6xTjZDv4wfFkn3ZKrLEFKFs1j27eHyKoN
hUrL5kvFS0l4jmZvPG9v+hs0vx25KrydtJ6ZrzYA6aSX6sg653CIfgRtftA2J/LR
glMLUtQG5/B/ZJ1WTNlqwTFvMva90g3SahVBodVw175W51+FcPO+ovyFZ3pEQePc
WPI2qY73UwAtygBoNXkYOxyRhbqFLojrmyWLaayxf4v9yTAVkgLWYG3ee4gHaNA0
95ifxxN7RMK17l5aSQD/CXCp143gdszu0d6xXf35i3N2VXrs/YkzfMklzMRDnFWN
N/AwR3nyQY/ChV77f/7MJvUDJxPVq+TGXJC6kajRwrfQ6aQ9Q6TEE8y8jBJrQ7//
04tpj6QxfrBGXAZEYplrw9chIlKA+LMiywv+eahOSvWtUmaFwHxzW5//Tr497YDK
jyqPe7sJjMDNO6fl85qE/7Xwe2NOVavTA0RK/Pa5JoruE0bi1Hko0BSlUi0SIoY/
zBJpLBAkJGjO5zwtwOgwmXwqlik13JaQ5oUXadhMxI1G0xOmdp6zmXMPpstVLQvX
7SzKFlJTj5HzQEo59lsSTPkCIj7wWRq8XaR+DBl4P6/5QABdj8seqEN5d0uhf7Ce
szf1BjQTCwr9RNjgsVYAUj3A6pEBCaCOZPlhmOnn970u6JyQttfJpPzIrn367Xhk
rm+y3K2zEYAUewmRpFqIBuu5W0Trwk27m2PWiLVR6l8r1p9kyt4HbYsIhI10RaQt
`protect END_PROTECTED
