`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xb4m5aF6dpPDLdhxMIJnfj6t6CHrp68KSEqJPUVmhuP1dOC7gc5CwXRm7ARn05bg
v7rMi0I8FUx1IL2cpiS8aUqxVRPe30HCdoGKWVSguJz0gaie36ltCxi6Bh8ysFum
Q1EtydDGFYG1pdNMuEj10GKvhCJnmgukoi2+ziCSPUH+7qQCCFO0hKBCzII+M6N4
Twz+C0waS+w9WItnHtoPO6D4R3TwNR8dFj9BBy+wkAlSAOMuOYVPVoVwdYSqoa+C
YYN49tCmPI/vgcSZx7poJxMVMtihPDd0d2iwknhWs8YjWc6Sj2gQs7Ox0Qq60wqo
NZFa1Fmt41ZdsVM0e3Wc+MDYtbyH11MRZBqSqGt59Jq3A0emFGDk5v5ai8j0Stp1
oWW6ZucJpKRU/Zis7XUuYOt1Kn76HtyH0CDsbx51OsPhomYXJZ+5UuOQHiJ0Sk2J
Jz242JCYbzviUl9I18+EcFhUMHntlziZOa23l3Fa/gtsJMGqJIqDhwToEt3TOj7d
4RLlcIchFLTSdcpxj/LrGowYElX5fYg+o0Ie4miqdg/lDz53820cAdMDsod07Mo+
Lq+hZ3o8PQuFTZ8dfPqEgdo/gNTetxLlAZGkhBHIi19YZPiuVd68KuDoXTWg8NBS
iJfIJpewI1taZnDrDN4AqdLghpl3doONe92DrYoncF26d99gNnPjKic1Srbrpq3s
0fjUUhjp77MVGuXnn4z3DINVDTcpKbs8yCLehR/C3+yVJTc4Zheu+rBPp4RWBxXb
95VwyuezFMe676wG3OCGV+tfnYWZ0Y8v2//9h3qh+q/8UzTb+/1XYs6ArJ1wz+EK
Pu7fJ8dbRqxkMy2EEnsMTNDEHU2WPLS44S/cx2256S0J4HR8i7cXA8AuLIc/Wm8j
OZ5uxb2CGS5X16+p4kX5SRDWWT+mGob8KWzJVNVYD0gMC75O/dbgbp4ppPWVH5ud
CxZE9XXJ8b5yJatS8Zg4CSnZFl/XPwLzQ1nXi+IPpr6FeTZF0FHup3DFG/bgIb/i
X576ablqfWgTZ6PknQ9m7CZFXsS5hEW26+or8LE4ZyKYuAMSm6+Pv4wsXeG8+swG
60AkuAoZwz1MjdvHpqqnuEVXDOeYuib1BW3XW044ewW9l9GAzr2roQkz9ZMqtnl5
487ncs0k9KXzxP7Oxnm3TeZTbYaom22akzSL/JJg832bjvny+zzZSCfGQkkhVQJH
UWCR7aZHLJ5U7/U8EVgKvg21e3i8wAUfnyd8b1e21j0CysHtV+5M5r+L2r4JBqDi
T78cFV8WUTpgyoatqYd0hsPuhjjggfoxHMNXdPfdnMa9cL0GVOUL46q8EqhbofmU
LK9BkxWS4xjnrUIxVWN8KJzW8a3iXJx3flpSpzuMt0p8vLBS7OuEXO3ZFGQ2/v5+
BcQAZAVWY6uOUMcKcxYXIQm7RjVE06pQ3QcgY+T/ZAm7FzyGgTmB82Fh1zCfpGJj
bsUEiLFHwfaVy8/5rnk3aK5jIpBlex+KHq0K04aIGkeG2BZL9IiDq1Jr2iPr9gzl
/hjJutDv65YPayQ5xpMO9Ro7R9CAuDfVOxAGFjms1lxa0FPZbGX4cFnuRrJueVb2
EAACQQQx/b1j7zmz3xSmOv9QEMZPrzY8uT3DbSv6O1WKdnanMSJDoECaYCXYOnfu
2lNJ5LmCBDBa6NNoO69xz0bCLPvi7ErZqD+AX2xjFMK9J9yCgJ+6Lyk/+IMabC4J
1X5ijXMl0rd61ZmpLW3NN2jPr/o0WwlyP2DgumwoEWY=
`protect END_PROTECTED
