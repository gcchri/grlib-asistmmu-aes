`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uxSG0IoZ/3nDK0b6aL7d23173KlNcJxgSxNdaZpDqKGGldv0J0S6RrttAld7TErH
WFrjCtKwM/NM3m5uiluxjnlK40hA2reI2p1yPIf/FfyooQNeecOxv6UKGMMQkDsj
Ve/OexMjq66wW3AG74UGA+13x0FBvBGsNFl6N8wYQRd95rz1dusMw9eBDq8v99+L
3IEeJr7H8FwcIY2+vHzFWdAkkF/dRijXfMiNQTTtsnqondXSk+jh82rVdltMU0VR
Vh3aBvlbwwtIzgxhoN8IhLP5mviDLjjIPnuVT/5ABZtC0pbbqpJ00EvBPXgJMicO
wrt1zUveuM9nqtNXXxQ7l+QQg8JfPpWgpZurRChV5v7ohyCxyFqUKW/PXVOD6Ltz
aBnqqUXInNXSGRRp9XpK18vGMqXj59yMRzvGi1wQeeI7C8yzj+bGblEMXOLWsae7
Ec0BursgBH/UCjxk3J0tHPS0ASMF0u2Hx5t77QsRPpKLT14oCM5rELTaUcWZPiVv
Ow4lQUnStDyaWRG4jnrwSJc0o8iZgKu80GGNgZoxc/Mvh2++X4Y7XgMjQ3IZrVmU
wNNa8sCeXV5cTyE8Uvi3sUF4fEb38HY/36A/nMsYftN84N85cOU8Ri7CJxMUldqU
fmRxs+EgqNoKMXMiqufxWjGtDKquGBh+6itYRYHcYPrt2+NPgEWsVMAosJxMENHk
0cUIp0DDtYyG2HJlOunGRfe9J/V42jjxw2rSuMWD8CUZGK6IWSYsM1CS3iH7DC9V
sNSDlvE5k7qyV6IDscOccgzIq5NV/lrwHWeg0gXVLIRbKjiqJ+KMkLRtWyPORP9Z
yUW/F18XA+LOWsimsWi0uxBCYsb0K9NDA5GVj6KTtcS11TW+V0QgWEzWDWZXHnOv
oDcyTDHcqtXocBCt1fZLk4tn6wBfKHjtN8byXmxKB+9Mn8eXzLnzjXywQM+Wrj+L
V8fGHUBsO/+ZEf7zQKG1Z7EsT4OB7uzg7aMlzh/69Inb07sHBrQ/ThJWZngGHv91
QHGWFrCU4bJqtO3JISKzlktT3vjaD1gos2OCsKbbz5JeQFrlXtVWES+xvuRbrGRt
cgPJg1H8nUYoVfOzOnoHbh0G/r4RURju4HTRZnp+fH/RwSyFpJPpwOO0W1/SJMIu
RksAI7jVLp0MlLFdN5V/bYIYbND4OJc5eakirAA8X4ZSdouudjCBACSPXQ7gebU8
cO7w4KV41AEhOdBUfPGJLTAs3qRcWYb6IPAJQiMze5nKtg/yM3+IHIgy6SRTQvuo
iWeNWHZwP8gR45x4vM49F+wWOCkgmAK1US72CaIQG0JoQhF9THeT5carmBWjfHch
K10vmlZ3c8EZNSJLUMrqKBr32C/KJWI7BEe3b/AxeKs=
`protect END_PROTECTED
