`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCLcdsnMMMvMRpKw+O9V1TcPiVkd5KHh6FiG5gAs/JzorVIAMaTQci/BxtQoUPVE
zHwKAwO+efrAMsaYmOEZhVPNgWbjCLAYpbGPj4tUZ7b8BRrOow0Le8g2tA3glo8w
4Kpe0IGNvHKurQDh33u4saSkK5KqxXeIxKivPuf2oE6zxgfAsCVryZwAT2baTVlk
LddFq62aERSolvUHAZNvsIxR3XDh1fsVCOgi7rYaCUBeWlI2hun3S7zTe1NseGLr
iE9v38Bl2rpx5LWKk4KZSNIlLuuDF3F5L1U1UqHCdNSvWuRuHHyhokecKOBGdmSW
FuBnxi9Wr/f9pK0S2akinCROMPE5OYKlxzhc30jF9eUnCjWNx9ZPQe6dFCpyTO58
oivslM5VYi6JX9OLAmAOV1rguItnb3pgrzqKzDTpbQNJaGvoIO1UWfvNMSQU6P4J
zn7rw3WZNJFPKPSMQGIFKCR8NkE89UOwkXqIwVAxK0ox2ouDEepEqFKxingfwh5O
HXTL0gv9xxnSFxjCGPKid1MqtK1K6vAle9B35Dh+IyZmMDoa/MYSaQOL7wo/ChJN
Tes9zgSsde7aM87Urv5TKaLq7193FaBS7FfagRF1mbEv25wn6xsG581/Faa/mVD8
dKT/1JTiQC+K8BK2MAcaAXHjgXudUOQklCWZjXuUfn3Unxq6XgMSenLApz5wkpS3
`protect END_PROTECTED
