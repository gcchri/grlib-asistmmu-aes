`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t5VzXzsSxwEWn8rFCmvN6qleXYfdhETMgmT7N07ixzYajrmifgb6xgaSEW3VJBLL
h+H2CksER+OGsgsUazwS+HLsDGv5lQZZjYRaaSx80Ut3FMpzBVikKbPD/camwmzp
a8ns5+elSxv5p0tvgPWxkelqf0fU8Otlnext3p0rClCdhBjsN8DSvJryRG0oCMCS
ZddivamZljUn0Ndv4R+vR5AKawNRRQ2lTqHQm7NyOMJR/ueplOuFYClmULLueR/U
nJadaME1y5nTw5NRmbF5ybVC6S5UoPPskIBZxnXE92YhvuceNi7znwe+4boGGUXO
rRwGSy7low72S5ZhzYLcTA==
`protect END_PROTECTED
