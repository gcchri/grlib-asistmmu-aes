`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z2hVP+27U2JoDIqzVVHMCRoyiBfdpbVT2Yn1x6NGfrF86PcPk5Y2o0vBgAtbfQ5D
rl+CjuJqYkNsJshrhnCLS489m8GE22cHaHrtaAF6Y5QqUwLRArjsK1oTq2Qgnigq
3QgoC1D5gNJ0Il8XLPEwgc4PzUYHyEp8+fOoSuhBn8SFyryD+8kLHqN33fGEa1W9
y9xPNgAlONYKM3TuroL4ze4bUdlxY8g+v4EhMt8MAcWUj+2CYZZ/POxMNje/Nsbz
M7Ya9re8o+bz5cQ5UINTH5+/gVOUPES/N7IuKlWPfodvgHPmsrVbc+C8TAN1l5Jw
KE76ghL1b7v2Z9NN7ZUPvciNRtQixb9OiwJojxLvIKyN8gya1keqeFhyXC/1E3K7
tQ1zWax/AT21/lNKgwJsRA==
`protect END_PROTECTED
