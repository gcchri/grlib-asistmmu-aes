`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOaZPt9mPMxILkIaJBk+gEYvXuvrKpM0NXmx58EkPc5sNDIGHMCMxsjXoEtL/dCM
tOfCpPJ8yKup9vCNJPct8ALZTV257qbGF0Z/hC/8vpoyZELqSDkWGa+yQjcxYiPE
J3xeCXbNEh4sKQCCMwK+S1DQhk1z+qPZsE2USxNdvToLvdyuc3lGn42cK+4frv0g
sSFSbLwC995VoQQZpr0O7YoYZkkUjf6zLCMDaNmY2mf4FyXap1/TtMASxncK6LcI
2582wiXVWYXgScISqwAymUGdGXCC/onwR2TbW4/IKgHOVorud6CJ5lhuBzC9IyMO
cf9sOD5EOGrakKkHYfrnMRav/PJTCFJ0PlfuPcDEQdHXRfMMy7uwTLuQqkp648tB
z6kFW4Mm91X/U55LSTN0ctrcFcxcWjzhcfk8VBeH9Lg7QJ6+iqU2VSJqdq+Sum4d
i4WgYIWtucpv1GbRZdeS/BDm+uGoB3uK5cXBEVVKkXahMo8biHepkRkOVvgd2CUc
uUm38QLrV37+BM540e3SuPUhEymz3MLG5K04VgpMz2WCywEukhqfnAkpHxthC1XZ
0siLAJyjgN/ApP42dxPAus4oH7Da/dlqXfMp/6/Z5JHDa/bVL4dOhd+4K2xxNXsi
61N5uWVtQQ03ZJ8z5ouhe65jbqEIpL7qDBQ2BG3x8npdtci358L5etAdFkrdMrnK
j6KweOUexd4IAiPqMAlsmYCE+zILw3YZKOj2jdKTIXrWGBHAVGNzBD1nHvuHVRG3
mNiIEyZpyN+VU0k9xZF/n2SHroRyantSjynnkr2jBd0+cWnS+Vw1MOWyDBIpYIgS
0bToGfg1yX+miWdV+JvbmrGOE8JQTmr8Apu3zYBQgCTPRD4csK0SPtyJFee67nrp
6ahNoa6lPCURinwozreNyF5dXI+h+ei/9o9oBt/TOj24dCcPcMJaTqpSvT8EdjSj
gCyGm8DuK1m2YngR8+VtuhLBfOsmhaV0jWvuKg3EQRuZbfVN0UZOTjthOWZovh26
ixxcPqHloUubvFbnGUHWx9mXPt82O7jZiznN4MVoJJ3fwp7ueo0N1S29ElNPgGbo
67E75P+AcmTg8KSMUUCS5Fg60lXCaTNrZ+3hXeZzXQ0gzV0wm2zQKkhW49pN7UUE
39EpPebxdx+NAQ6rDykFd0pLov7hB8tgPM3b6/iE0qHYi+Hp5R6EcQ9SK1dRG2/1
ujo6YjJkgoEEt++xafuOI6Biiab1/ASggJVyKKkqvGQauyZjg1YyWKk98QQxhCzt
QLZenD6201vNCWb7M2fQyCHHWxz25BrLuRQOJ1IjKpLCMRigEAw6AQW+0f0MEoUe
UnkdeDJAxDqn1JTXVfHitqwujs3ut+oi0FWZL27VMHVagZ4l34IWh64NgTJP5ddy
1Xops5tLkiHwvFSQ7AnUHcI94qRsMeQ142wmhbWyugn0/28UEC7kajpDgFeZzOxa
akkRo8RGVc1aBuYzRuh19kj1Ag/jjBvZyX9zcGF6aan/1hvNsQJFh4LiIRmOc6PL
m6dAkdR0D3tOwmV3UAdmo2bNoGw5sWbuZsSuQWQ/8GPYLM4Ep/Oz69upGwi8iBqI
5XC7Da4Ot1JRynwSUfoLiFbVlLxjianKSPIZ2LZXP4Re7ni0MxGub2r/Z3p7pnAn
3ojo0lUqYuV1xvgi5AdvEe6HTB00BYX1+VyYzlM2yYeiUY1ylfJp+JTecVrLNF5g
WaEr3XWd6KggUOMpcbgp2peClpeBti9UcU6IfsgzAeMqOgveiA3gjDtkbGRSfrxF
GD31KD5K+yi8z7xRHAy37J9Bf0uQBds3Tsiy9wgydlFfAC3askjT/j1bWxui+C3I
uNMCD3gHix69QfKgHC9/8PNdGxd6JMjJdnNZFEypUKmx7Hq/ZS8GgAs2VnNCafXf
edXDO0OzYlSmDusZ7fU9cGqTPr0qg/GUsf8025xU1q6BERU5AooTvMvQDMbOOXXZ
mSCDQXxURESKF0PZFcUWcKXaxcP6DySSfY4x7KUqGMLpkVFLEYCBr3D2RERzfAAs
TaP9UJ9cijjAJwux/1HtEHeA5yH7RRqHWpghDQKYtA4SOqTJVK8GkIDs+CCVsPyM
NYOdURjXkM577+s2mUE907LXxlIUI6uLaoPYE3cQrYd5ELIJFT5S9GuN05Yq6Yns
JeXOFDztMrSF07TekEJ9KpXsiHqyFu7meBvnf+ARwaW1xutySxvTF1sQ+baieKF4
p6fX9MUIzxSUF6hMafB0R9l8VnVqLUuo7/R28lWYjLASb7cE/fUisF8PSlo8qnXT
5XipPD1enFSZXbpnYKy944Y7vfUWGEbCnowXIiGvELwhgaGY2OxINy6rYzrrZV6C
b8vf2JTNEx+/tj48Oos1gnFaGUmfa6HywdPQl+J16yakS1bB7ts2uEQvy+3Oogvs
vRwcyAKoa5tmRvbL0GR/Lr9kpBbjZfKt/jumispJnZT41CyLV+ODgf33U9KfCG+S
OsfcwUnQSheddhYkwjueSrVAnjIWtocrdySafkT4AACKtc7VHjGGe9l2e4lEQKll
BmqsDyrmjRwigdMEtn56QqFXO2amfYZPZMbPjzFcUv8DCld6j8qe6iV8FVVOKDNR
EgotOFrwlGkBDG+sYAcK8SOs54lH+hwgUtTjdE1PNs44hFomWX4hNARwBF51OlH/
hfctRr6YEZl4u0+sp80h+yvpad8R10dLWmPLofJDicD4hpUFNXHE/buQiFh+KNPr
+W5/2AZzQENn7iQi0DPqgvEX2WgIVwO1vcQX3cpTLKrJNZ82gcdJDxFODQhm53ty
GaRwGQkbGgUyC8yHSfXneD9TqTFud8G5Zty2LDauwWmzx4mgsf71NWM2BPcGUpWB
NRH2NgHASEfxJflEUSo3huLMLIwrHTi2yjEnxfCzrWpSTf7axIAvIMs6CX9sVZlb
TG32aw4wU8CVZ4F9O7VaNlZHMxSk7l5osR37c+8lhO6qDSaRq7VJy+MxPBlZFhr7
I/0eBt93z0ODiY56SXJovbFECiO2Kfi31dRCIDT4JsHW9DlQZmci9sdYBfay8wEA
IwbPSjLHLCKJzmOennv0p+tMv3II9SOqr8XNd9WN3Iov9MRVinIvYy6aa9nkyqei
WkxkTQJOqbJMduvdtO/BMStQq+2hBJonlschBQ+J2GiPzL0T7l4cpH8rvIcWBt7E
S70VGAp2aK5dd29Om1g+1I9AAab5+mS/NUMkhyKQ83ZJGH59+cp7u4DhIRA6EylG
paHwV+VRcH2vdwnvoSldUSQkQ+qbVWZaky7XDem5LnFc95o0LAkYjvauMTWGpHqy
CM+WcRpA1+gPmMWkaZqsNAs09OHl0d3T0jp6vZEYx59F5mcPIso9MpkFk6QIWNn2
pF1V0vCt3fSDXTinCRFVsCKnovOPeBfOawSCeArVQgZ6fc0ueHdV80TEDt5AD6lv
xvWiQtCO5cFLWOi7MOsaygOWBBlbjxfyuzeGsDom+pEfDNTuwnK1BXhV+lsZ6cfs
No1yx+X57dvAUN9KcCV+HDuyvFaFVyYsjVh3AuAmr9VoKiBXZ9iY4ubgdHlHAy/G
8hAfmsS2m8iAl4aRwV1ldl7ECHf1Tu5sJHdbNFuHIpFnn1oR/t29dezM5aYuxw1Z
/MA0Phg+c1IdB3jMWSC2E70nO5dTczfwLcVOolRTOZ6XQ0IljjsILDzGEwV0DBTe
bfKpTQTjhcdMSvTR/qicNiEMUSK0WZtLXiH0NhYit9bWp2t+iEWTXUoqIKtzuB9j
pbB/xSNYmlTSvfwU991xKn4jdMTb4Cr1qH//2QIt1cAuyFrIt4VRPnEMiPjpEub9
crUDwg0zMgE+TBTuSxpv4Yc6aBOv+kcF09V7Cp4CVa62MFOfysiTUmgp20tSJ1j4
32hnCESMv198iBEE/Z4X42sdmSqy6R3cvG+q534fqu7ybtQxbg+Ec8TlUDHDfqAi
EzeKpm/tbvJDRwrgHK3WATebowc4gevqBle7u7Hj9sNrpFbbND+XtEsQ+E4EfuYL
oVBhVwglbO3T1ir81t7EXb3WWJh417C9TWCFotZyLxEFk34DaBmskZvJp3EEDWRy
f8RsBDlHhax0nwhMJKPecVn4/G/tYeWXuk0MTMe/hmRBxsGsxrer4cKrwSE8Vyj7
YEErz0UrHF0YtBXSAyUAEd/r65B92tTeEnGToz/wliwF7Og70PPRPxcnHpaAeSKM
xg3k1O5vn5uO75pUHPDmr3WJT81/xd/wtrc8mqNOapM61rCqVy9rI0udE9nxTxFR
4hH0PwqpeNK7K1O1Qx8ESjakwLlh6oBI6og0KYJnxdfv/cJqlTiwLXDugCk2PLNj
Y130iiq6uKINPwd67H2ut+XzFdvVoosEqGGtbZmgED+0t2WbKgXJbxTWm54XGOfv
1nnBO1KLqLKKJiG1Fj+abaN5DFdo4NVFUZHcmcelG/zHRoJCRFFV9wIZ9iePSneR
Hk9yAGp8leMoJQksImIDDWFdWvnO0bgpCQB1Qmoj3E+shsjokbkqEnlfhywuoDbL
iSiU6jvqPlxm8kqW7vxOITQvpzcuAcoYKBgOEakqzZtPvxYsQgtPLI2U/2d4k8ow
yr01vqHPW8gQuLB7FWpIFzgkC815SI5q782XFMvYRQKjXma6XKzmv0fnWUNgF0rc
3aNHAx0/o7LEHlWc2KILe/0nsh9LTxkoXJsa8bqnMTDXzQWhtIUIH50bvggBNVvu
SVOOJwHJqzaAqOFRYVceZ5afzTaSwVRTiKfyxdgHozeKFi/QkW8c+ZMzhNq+ANq/
y0fUmA6QMZJsNPz+qek4qDJx+L+hQxsamOBfOs+r+JYRXLEfZJ4JBBtKTrZUc5zw
rK+bNVEQSRkzmMeD8P93BXVe1qO5ZH9fHrCOAtmDOZWYQ/9WgQteP0+UuNgsyYz1
CjkVouwgUtlUf73DPe0boCqi6QMX/eAGu5+4Irbq9mwJeOXMk/Atc3khP6+bYyTu
MZvJQHXiydJGo9AGm6tnlMw2av8VjCC/hyUb0jcdzbEc/GL/RVIaLJm88YrQOJYq
rhc9Lz+nq9MfAKYOBUKWzITV2o9wKhR3XZETvtLk/PYSNmsOtDTfRwOxM7bC5zfL
FT3SHeQXofju+wGjno58Jm0SOAuYF+UTbIdpC0ocshBxYS5QP/owBAG2pB6j96pH
adZN/EjcXeMWct/Sgf062y+IwKsL1ZugKR5W1hH0CLUj2U8M6TUxCnamRxlkQhi2
wwcDum9vQU3q7b0CFSMb2o9mqPnJShMbPS00gK4jZKmOENS2mg4HCwruSx1HNfjF
X+/PGqeBKkAJ8SOcXKptkatGiYvzSrt3bs1fYawJV7jXopMya0lVQsURlMNoTFlY
j6+Ils7XFqJPBI/yxjpUFsjQx4EjKCBgDDaQHD6iJvTS2U2FrDO6y1zG/N3iaSLi
dWFio2L7KO6iNODEbBJWbxXgTM8nqzvOQRiQNWuUGhi6ow3gYTYcKSgTJ3b10rVL
HzLfjy5n77PrEBadnc5V1nxqRIaNv2n3ixZQA9HiKZP12QgvwDN+Ha+W7m/iO4F+
SsPJ3X7vMFrM0qfWRuyx24h680SDHrxy5p+1M6RAawjZP/sJJqxS8az5cceoPfgn
wZKoPMbQfREXVQeijGn5xnsqHZhXMPJgzQ+cBz00Wx7QXx1xla1HVEf3JYhsLtcn
iCn0kAfr39ciPTQptyvk+IFnuk05CIegNfDud2bfEFDvLXuDlvxHK67SIGywEC+4
G6GXCxM2mJio+Wuay0thZwpfz7ad/0dcgL8/wf3iquhHYxyHrUmKyqxhWW8qs7V6
Oj1Nc6uX9mv5cUEscvazC/mjuFlcWEAsIei7Nrwa87yFOIHTY/02/l1zJV4RZJWw
ZZ/a3SJEXA1/LWmAWbKvhGI6YhnW5XDLkv6T1alyGEl6RnmBiVNl/Yb4dW7SIYMo
EpnpEhRKygGaWc229g+594zA7CnixWq5JNgjv9/TyWvMukh1El3UKdOWxLFts0h6
`protect END_PROTECTED
