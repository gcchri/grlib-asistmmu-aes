`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/H0c4HSl5dUTAaCe6Yju6n/7hXnVdZRDMAgRdan1hSNcso9vpeuY3k2eqmVz3Zy
G9+B6c+kyKQW9UCQUseJQZvtNKJOVhN5fidHlFw/ovIUWPKXo2af+ZCJSw6JGbQp
xH2FLDMqg1kd3otDaFO1af9dNPx2+Uvh6f8ke4PqjYZPByMNj5Hh5etZmIHXfzIb
1R35HFaEqqUgWWnwDMEJb60JP0TxElxowPpAJwwl3mH8P+dCwN5aFF1exGtpqBI8
3HibgnFW77XfXxq8iE3Cjl0ncQkfYrIgEDTjYHPNleW++71v2Bb0Gw6H367u1Eoo
KUUe0H+QQyk39KB0B4tmSn1xJ5u+2JMBdrtAaX9Rm4FkHUVNhFeoa+IFMsy2/fdT
yx6v1RjNEdokCOLJPDSf4Kz4Q9H6RUuD3NggkZ+TFFaeNFa2MBMQb/w7Ss4ig3BK
0OZWFSdezoL4Sfhud3ni5tR/Clto0SQUc6p2P2jtaFTX8ksyaR1bFlLINFgTW+AN
wYA5qlGVE1MnRwYTpFuFSyYoyQkeSPLmJoUQ+SQ6c+Lad046tuiHD1a/f3gQuFp9
hMmp5g4XkmzGsVnm8IVV1bDLb7cy+Gcbjq930ttBklEkmD2pt7B+Eq9qpE6jJtyx
EiV4M5wsz2bzn2qbfRfZjDqJ3VtubPSsRibth+r2sv/IAnjaj0+zJzFkgWZxLYVd
nlbR7HqGaSfZPn/P4UBgkYpX9MdTGywBeqjw7Ssh/GSj2kjOy76RbmnkR0KUDpoO
NHbHwrWFZRxNebcQ88PgZnIUdtEABDLTvhaA3xdSbfkRfdBXoxLAmIqay+SUp48/
OOn9U2bRamWw4tpZrdnNcSiBZMMLxZ5q/mMik8yIPF8=
`protect END_PROTECTED
