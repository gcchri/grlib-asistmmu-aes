`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eKS8kF4RMvduRA2yDaWtKPsxS5IiR+ls1z3R544Oi7xVCz7v727sgvHQcNQvWdxl
YlKbd8d2p1IJZP+qazfXLc7yXqJ10FBF+z3NX45dt7UaoRn8THFcszBUz9CxCdpR
+0yYP2CKIwYtFiIPqLmzegXjjPR678SAwzz7b4a50RpQz02A8CZ8EVJvK+hbJ6s+
uSe4La5bepXJ1qrcCLkhXoVUM4KoLnOPkRB1w0U9Vew2cNTxID3JCrD4aSLZCmg/
K95NHz+RZrjSB1CPJmaAMw==
`protect END_PROTECTED
