`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QBpVYcC+++q2GVufgmd60bWKe8fXqWmcaynmfCOAyRNDy/SWPxfUTGQECqY92brJ
yHFVOO0w8MW0mSqDYIoI6xJrVooY5fSs2lmzLMdpiMvrSekHvRDNGBhHwvVGr9K2
+Qy2GZyHLc4PVAjT+JZzekK9r9W7ffCDeSgv995nIl9mo06P/UtHeuvOMDa4Orqn
fP/Ld8l6Btf6vu9J9qrSDnNUhF3kAb483Vl2+Y6YmjwmMU4BbGLRiyVcqfjwdG3c
HFzTsmIvp9h4FK9LzAlM+SLU01o/suYkJzrvnUA2Oj6HxtewGDvxycTjyKlAaiXo
1FTmWhJyhQXQhcaoZO77lsZkwMdoPZCzxfP4TQb1DtilqMPjaphqnzcmZr8m0IgJ
jDowMXLEGgTxlUgaxeaNudAn1t7ysCqwkWvPJyMQUNfAfmL4LKEwcdvkJSABmxEB
1b07W/73y2wKKxPOeA+F6cXnrZw5q4uPvb6+dp/QI2AVOkiDpqC2gP2w9BCMAIS4
ps9HDR76j3IDLYD86UwdgeLlLHVd4zrEh8loQRVUMH2KOIzirXMZ4qB2wdo+YbWY
gnKLiLKFvbXCHZg2jA7hwRf2QaS/SQDrc7Sxf0FINRtB9/lm6X6GhLbG8bunoZah
yucTkH80qzjwVqm+iNfFBnLK59IbcudR3fEhotTarcTnyDm5XcQiVjPzGBNXzy+p
`protect END_PROTECTED
