`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uTWdgmISHE9Yg1vXD/glfEVCL3bb8Lgcsls+HfMBHV3TZhSO5uVIAMuQcnSVTlZH
6SKg0JxizNDpjAgide56nweh4bWE0By47b084n5y1TxcfSJVRL3QU2Tkca+bthBa
uMevye/HR7WfDwU0/7RnuEWcDNEYG7fVxSbCl2U2l7yQBcWf5gBWKyREf6lY8sXL
5oqGaBDnSXUlUaKkfBQftCxPS3VySumsoaQlqUuBHOYzr7vMWRrJhppvCdqRWPUn
NE/WQV+2bE5NoyBAT3qs0/ta1br+S9ap4FXiSexQ5jCB81Ec05fc41xZG5jbcS+A
O3C7mOucinlcdCO5+T7CA4Qay1T04nFywqPZJuenMHLVAQ9NfxCK8hA6/au+fv23
jVQ3uJOAQWQR7Aw7jbKeoib5gtuCc3nFI+xCsWCRAWxJO6XgNfyQexS/1izSdbBX
6Fcg9Ns7Xg5XvuMzwC6a2gj6hDROyzyjV3yomyqzEJvix17SFOCfRY2a0kK1nitk
`protect END_PROTECTED
