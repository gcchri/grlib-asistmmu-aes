`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiwPm3e6Udn+SdRevV0FyAzzVv4lUajBrGleBLUDQUTjAksDUID3f9CvX1HcKDOT
5T0cnjZY8/rqVuGtkr8zLRDqmUquyKWt8nQ+c+A5eWDJDXCXkHIxU5XSmplr1r5o
Glo1vhOT8X9InKnKxYTIL6zMUhW5WeIO9bHfhE9zo8YXeGXspOhFv8Rczb2UgemH
tMMfc20earOOlqDTR+LX/xU9vYUFnDJZzrRnfoxwCigBO5PNWoiwCi/kr/1831W3
ZLDC5G6aG6lu3G3vsJEI0gv5980L1Nk0gGRrNGz18xqHCLYbaNJW8q2cJE3AmhTX
ivfL0nGCaNlSufgdeZ+5EVuGjx+r1wJKRguuybW6urTBlaxRvPRUuAr6utZkQerX
Za/Le43a8Vi/+l0u4to/7sJ4BBPdHPIyjJTt0cL5rCeTQUhRR7UnM0Zx6fysYfyO
Tc9jzPMyC40+EShsVS4An+///pomtlS/Vsr64X7rpoiRx5zFQlpouyGajQe+cpfj
`protect END_PROTECTED
