`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fSGhcrdjEKHhvGitTvA1K+I1FbXUJCPAGqR8g3SRnH2NooUvbPSu0DZ/ceZe7Yit
AVCY98cosi5oDPXvtqDk3it/E23VoiTOu6TXw2TRjxWNzE6dPdVGJlm+Y9We0nE5
cxXL/3dGMjZqNvrGYyyX1kqhgPTnoy0B+OVeKLmqGb/zpt3I0qP8hSVURBbTu5GG
i3NHUQLo3JKRZRrll3rG9zvDk9S2GhfYn/fZ9Pf+G0Lj3f8cf7l3Hz5xLjAMKnnB
mEexCnRAaS6o72v2pDi9/yn3xHgHfHWpYOdmL0uMHn3kGnfTLW6M+YNOLRFdRogz
1uyQAzaTPxRDMndS3ImDR/uQMxD/96nZWzKlvfSUNJKYE1UlFC+wjqAlHp/oZV1J
Q5e5GoFmKXqMrLP1/dht/UCbGM9CmnNLq9InYBUMzGIQhdJN/wvJ+iGsd+JqL7Tr
Q6x6OWSGXXXva0RUjqUlVXE7GdFFKOAcxSAw4lASOQE=
`protect END_PROTECTED
