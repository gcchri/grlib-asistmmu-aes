`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ST7oSdZ41uRM6sgtKmadzSVAQg20Y6yTZI3eIjU71zIys8IfgVVow4Cf7VOaige
oTY4RAvmvqcl8wSGDRCc/OZ4flE2/Khcgq7opXXtFn68L4gG0NTPPfDUN0G0zB9L
V1XX8vIOIU76/HWf7RQtAO6LXpKS8JuMZImX4VPtigghsYZccT5PeD8XBui6Xz+G
C9nPe6nXMYrBRLEgPmY3qBhk6tsk29rsV4InbFg+JVGDv7TmRUO+nGDbP3MhIQcW
gZWPhXw3LLp5WRGFKodP//Y20EamcapjK0CU5r1uaICHsKWBOzcJXZvOGAdyxSTp
xGeHY22/Gs31R8sQIoZc33v+DcGufbvERSp2pAmFnDbu+q42Zqj2QjGSwZ5sA1lB
+35b6XpmM+1kqk3A8SnBtLlv1W9xV3eqApI6LKbvY1Y=
`protect END_PROTECTED
