`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
utJY5w6ecaLpP6qszyDKy0fUf++ROM6IraawxIsaCu7YH33By1LZ3NSd2YkDBRMX
p+b89uamLkaoVAV8IzrnsfKuNAxy2jlvC+xzOHvTLugvZK7jQgGLauLW1WLdjd6W
GHSVGssegfzGRSbL9r6DxUEskqdqYVwMe411ru6hVOhbvZYzigdINdOJ8CKFV/2h
bT9GM56UPrKU80+a9V4Aea3+cqgIv5gNW22iPHxQHD16Ch+tdP9mBUQQDZ8CHmuN
CGRStLVGMLo7xrJY8CcRZqhJu6yuk8j39AHaZvROKtWFM3rIiFVIWZVjyn3zvaTG
jSg+6gwF5m3XvsUkWGjnxSoSk6t9szjbHIdFGKGcJ+WgHAIS7Gjv2jlBPscFj5iO
ij+IFD72v61oYD7CkiJjlq3WZUTdFjEW8FmK7nio7wvfpGGtLXriliRUxq1+2cOs
YrUwpJO8VcqiW7342hLqzvh93KZJ3rq3tG2OSk5xQ1LWQDRKIcWdT+KCcTihyl3w
9NZuS5zMsap9+8DKCKHu4i/0Ax91KyrJ2BBzdEj16mxKAkC4pHBc3a+/AvBPrcoO
pcf3AgZixGtzSN2UJsiRIlXA/EaFr9JO2flwnhqEZD66g8HA19q0lcs4EXD54wtl
7J3AyZ3iJIMY3BT47tYlO2h7SH4di59XOxi4zP5H3RqBlLD2AmRfIk8QPECvDekU
IBjynGvcUMeZVHf233U5HuAmkq9jZzm9+u+YvXEZSGU5BSSBY4i6eI8RIeBuAm1U
CAoHoKsvhnyyGSvvPbPd85OdFk1Y+1oDDnLjy4L+lNTYhXQKvU6vz068dCV8jo8n
KjUBf71bgl14EkWQTmPWW/bhvPc0wJHGfaBW9hMAmvJawqZu4aNBCdW6+2dq403b
ZJTxZLj306z/ktA/Y2VUFUUMqABRiek8HvK/L5KZSwRG9WUz/BbFiyRe141HHZ+q
`protect END_PROTECTED
