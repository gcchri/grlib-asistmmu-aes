`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PhwgtmnIeffdsx3d2Sl4u2MwooOmIyidmMw5daOsGedKyiNnUsMahsUwewUUb0hm
QvUO0molx3Bp0YNoPLE/RHKyk1JRAI+9VEtOJ0TZHLTLcaB7HYOovPOtjdue0kSm
dB0Sofo1rtHPWgAMXUHISJbxWnxZiXqmbbgpfiV3uANVbxFj9JdpTYyy1MyEOpQQ
UVAIX3q66h7tC/68nTemhcNb0JVwNC4skUNrGtR1m8AfJV0BBPVd44sKO1VyZ91N
pLZSZT9EpAehccadmLhTCNGbVtl3EM0zh9jFlhvWghi4UWLuoasAXvbnkdCJspNw
hIHoluJISICROI6IOwJdrH3WCmYogP4ZM6tBRJjLhRzVku+EmERXItqPuDCEyT+A
q01jCJA0ePRdpEq1PY76GnB9l/FTwKlylD4HE4YXHYLcFTQvrRGNMQ97guBIhc+G
+ppM+GfBKOT8WsCgLyRxciw8CbmoKfTX8smcWDz5QJU=
`protect END_PROTECTED
