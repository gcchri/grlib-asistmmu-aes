`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zgn/WPvGLrqzbjGSPQGw+3k6JtmY/q25OKg4OF+kQbLOm8azo1suAksV0ceDYNwN
TZlUoa/8RbJCUfC7GE4aoYZCpqEnLXJK4RUyarM4tkPsQwN+h1TSZ5UkGvXDlHOU
hCHZKuxW9vdIJSm4i6wBBnIN1xNAKdbUFqJiOHsmuOMRiMCxS5EeImXfoScz6pU/
x1HbwUDAKcjMesJ0HpdmdtbeumE9MAdcEc80Hi9SeBesuLKEw/uwMbggNxWAzcmz
CJVMN3k4ritFT+tQSbHluts693gWsaYV4wrcU7JNX3+Aw5K0ob94BAc7fJJebar7
YtM212ZCbk4qaUn5uFqESzVilsTE80KL27Xn71eOWynwvYr21sXVH6iwoyDUjpmJ
dEtGbMBOA805ewQ3OEXJuA==
`protect END_PROTECTED
