`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BnG9QmrBxxAvufXoohutIdUeydvqUWwp6bzWjIALiJ3lPO8W4MPniAdUwsAbX5Fk
9rzQHWlln0YzHOZr66ZmwhmStvjmsyHAr5u7CFLf0Nel7g1p5zamxhqP/fDAhe0a
z1b5Y5tV/rAAj+gwAHUzsD5Eo5EH8GbVbJeEbN+ONe+pUGdHHv30C1inCJ9rceM8
XOkM01Uk5UJGoWkz+6W3C34Mw0ZwF/mFczsd/11LYKdOFOTMFEDiGI184SAlm+tl
eWDYpiAthcX/M4q+ZEen7spFlcIel5GqPL4vkSAu3xhos+lBimsaTgF2lq9pivj6
mlDL1/sxwoCQT7vs2j2xd7KpD6M+SB5hMCbbIJW+/nNltJGhQWH5LCCnNM5wVznI
j8OQaID60yVkAbnt2yXPRL3jgZ3fMy4P25g01sUVuSNJNlgvdeWfF9eXdyi2UdxL
36f4Y4UoDudMmpy/iRIKFVB0WVrA3fi71/wOg7RFwxB6wwcG2pHW79hVeeWQv9xQ
zINGGmVz8zAGnh5UWAgG8NK8/ft+dc0cJBsPrSf2bJclOjCblFH1q/h4r7zxMkpr
xtFozBrfaRsQWhQmOsEVI2f3g1xDoYyL6j18gUfov3E=
`protect END_PROTECTED
