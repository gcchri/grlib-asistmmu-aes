`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDaTcijhhirisbNbp3pbDyXRcBU72caGVQMRvAXr3aBTWtbLX763J0TOLRcaaWhK
a5h5Q/R/VUDhNx1keOxGfId4G2bdYjeUmHYeYQI7zRO8peqEY3Nws1tkBPsfkrKz
FtEahvXrcLQwrnwLc3xZciIoz8uO5ww82c7aNXhbuT9qWZik+tPraV3JHQQ3CizV
bWvING1VpRUsNlsTjAwrrp22CDf219Qd0BiV+iMbKymlRJKjm6gaV2wPNFWRAWNX
QLbUVElTQO5CJo8HqF8d6SJ2TMn15B+uSccdr5HKaucdY4ZMuKPdLrjSJTY2Xshb
3O4Ncaj5YN6jKvAOz6SfzurtTy5JarPeHZXopoVS3u+5TzO34CCNyZ+DTXS8ZUVH
9HTF1CZpElEDGdd8yUFBlwbyc1kvX4VdW35ygvaTqHdIPT4BH7FDOyZgT5/nEgBD
Ozsgr4n819Dhv1qiYnK+NKpdiACCtQ5wuCisHNFLKWyVjckuMGsVEbEzoJ87NIvB
qPur/Z4M1xDWzHtumZuFp8iKNZda1KaAjVJ+3pmwm0vkr2I9ekqVjXxFMRWJRmgs
iibjPyJ1kw3DeNS9CzKE0tNTREnMmz4zdpQ48nylYNO4sym4tJKWA9EA1KCLQeNW
xuLO00AfiXbdPfzegPeNrHR7nWDI/qJooBs64rOnit6UJO30AS23ytARCOtZ5TOE
9JwDH7+mpMCb127H3VyndUwbyRtd3Qb1yLEOAkWsYfJqGf7JrrWU48QUh0Nj39b0
7PFZUJaL79d2gZs7WgRIbOB0gI+5zTOs+sW2oBfXzWvxE0TKBr3OhHAgvRybu88l
uZ6kMS9+MMLtZla6FvXNMiRL5TC480+z92qtB3Ejua8Ek9XsLxtKx1rH5tdls1zY
gjulknsHQO3KdXoqCcYkssRma2pwcV9HlQ7vjRLJfcJItqdWY5ptAAKjUU72zuuP
ORQHFOp/803BFc5EOGRelkR+uvV2nqIgQ+5DwcawurkaA11V/AfDYHCX6TEAaSUR
kVAC0ZFw3tltLnmHndcaM8uKn0RO9faZT2pHDpmkzFlqk8Ez9DwO4IYARxBefe9u
2yJ/1n9yVz3DJBnXzVPFg3/HgnbRvuOoyPaW5Vzm3wg7LPcl3WA03PoaWbzYuZIw
1KvIgHitkYa3IcFW0mHeiL9Hg48CsWX7As8A6HpsGe9DZyjGHs5ElcK/mujvUZDr
ehW62/aqlxqc6YSI4Y8RF9d0VyLF3JsI/UShkB/TIKEmuBBLO8uMgKkbAFIjIXoC
I7xxYnrKJ8MAj1Eh+rl7/5Kx3gIri2Jn0v7PKf6JJqaMR1gJ5/A8ujiHq9XHWshv
H3FMvVfI4VYywlGbCg5ARtQ4RpjZgQjqz1blQOKwisZiqrsb+Y9vFFzVcGEtLo9Q
5T7lY65KFmnB1FhAq+6GC4bgY9YwR94FIZnYxwbA4DFo+TK01nX/DraLjbBtpQ4/
TRnCkIif6yCNwClGgDw/q35bH8vtOutWNPSwR1dEHcMvR1sjA7lc6DFrpHzlC8uv
eQBlAqhtI9ajxhzkV60yTp/MI0lD2ub3tCq7p56hpUyE7p3sy5cdViKCd8TYsYpj
1pbrpIX85RZbaZaKlxM2HlFNcrKIpHa4U6buU45r0M2Yid12k3jy57ffXXSjU1Pn
ibdCUb91XAZlWc7If39TTmNSy+PUr/1S7wvr0YVKTB2ObuWiIEvB/h/WZjSbe3k0
meM+dfIAOFX0aoYzEtlEoWY/fYflfwZZhtb1BXHQDyWhTNcCVWrutfCLglSKWM1Q
Od6TaKB1fHcfdRZiCLGxLaD10sLMFw6U6bojXzyB9htmObD++5woo9pU55PqR0l0
DB3vwWTkK432zLJFEeVmycyeMIyuLmeOnVRmoVKCKf18SuDAvXqvIP7NqwXvhFoi
RbzqjH8TpXn0anaZzy61h4tVxwybnTSu8OiltyeFsJlhJmR3Y5G3WReZx1sUbs6E
yQSrbuWCInieYIDb6R/1YSYfiojkM5MvoTO7wTd8Xzb2LEsYQdLBCdWuHPoNNSWE
K16fddaA3jIcbBzoH7bCuQ==
`protect END_PROTECTED
