`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ayithxp+Kd7J9I/8cDY49+bM3F1Fjjj1EHesU9dHhiBN6zyJaeH3J7ldY74cdMKs
8RySBXHtwpXwA6uqSucLX7jPN678mEXqGB4Y7ZtpC4zh6jLyJ9l04WqLIahRbuXq
dpj7+VCKZhMzxSYaV9ALKdwq+Ct0G2CApAcsEINOqGepkNZdYVZekJS0yP7e4eDi
h0lKIjRnF8nGj7CL5Ul85us8J55qK7VoYI3kvJaIo/7JhFiTR3SySxTJY+Tms1Vg
cRXBX1cbcvid65z86ZSq4Qm4CQGmzVQfscz293urTOaU51c2Ih6qlSteJtWwfhXu
sCCKCbrvyxHR+FG09SSLBhX4ZYvSuz998aruLvhOO4VE+YnnqoV/d30aXm3ZioGK
71VwAbS1Q+lRWjUi1c7i7/09WtwJiFtNgliysa/+2ll27vkrdHH2Y6di/MPzVhke
3cGoK7zCrHacH0S3fGzwg5y4U9iTIxPjJ1GRs2mU7ZwG55bDARhHFww7WrHWhiP8
K+qISHqrB22nSBJNSGb9Mz59Yrg2mSy1OXmpH9rsNmRPlnMEdlGupvTlOYRlE/Md
lL/g2o9HnYcktCv+wWMH3Hd0hNrdbcsMlHd71zAt2o5JHItgNp6esd1pg351lveN
EhHgsbnvHPH2hjib4cO5b6yrmGuTyTCzO6Dy/4XQWNozW0d8zLiw6dBSoG3OAyDa
oNox7uTojoLQgQqB8V+2nZmeo2dPDy3NyTbQIcOKUgdCvAldym+MzCWRfEylU3/e
+J3M2YOe0VOQFyr5YCAZ41W/3A6Tsr/Yw2KBgpFe+l6Zdg9qvqjJdnjrH7UyJxgD
VboxlZRJxTUCdWsDttHjX6AjG6JK5RRXE6/xL/zYlr4l4vlBAHgX5dcBWS4nnnlm
GbWafJCeV/G4ICl74SQ1jRNYhzdzA4aICAK2W0Mad0jsV9je13Wq9F5uEwh71d9C
qiqzREMa1mXIPDnr2h+46mhO/d3C8yvL+cCa7yY04O4A2N7ZZkPUz1YABLKhLpNP
LLIpd2eeCLPsT8IMwCJ8wURWe+s8e0GNwz5Ly8NWkeUl7K53ymP1FoWWbD1T6SOQ
bzIuGNvnWk1EzxlMq905DmSiWt17t/didIT6es85K/jwyjjZ+aDYqGGOH7fNr8UO
MMVVrmAFY4CfyXhxXlWhsapVqxn8yDt0s2fn1+03uyqGbj9mzRwkW6l3eAFiC6yg
CYfRTvQHe6Z4iPuEO3KzUA==
`protect END_PROTECTED
