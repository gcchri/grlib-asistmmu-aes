`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YcpI9KMLO7b9a8numIkVtvY9+8KsglFyha+xzt1qqWNYBoS0VQUQd0zmoLp3Jj26
WFKLItsDongh18qGkwPHW/4I5gLxqeJySyG5NzXGbdQHZOWqrv1nds564c4yARkF
lxOp7jFoAUFSRdFVpYgUeV8kysWfJBpCWwrp8/fwH6vGbuvmfjELA92V12LYFvxa
n7cdE82MW74JDKHtI3RIbmFGKq91jTwVDv4aSe7sLwmWQJ5DPpBzB6rtdTYQawAN
trFLk28hs46MxUa96d4uE1sJhZ3WtJ5ca/epoEhrlpoC7tHF3xmGBGuL45xgUwY2
g9QyccYoCuQFp3LwzB71U0KlSMUjU22a2pCUVJV5aSJbIUHeWCqQKNkZ+cwrOYw2
pjizaKXvDcehESL4VfCzPjo17u4YFgyqB4+KuxmYtxi2nuCbQWlROFI5tk0Js36w
UGI4VZZYoz/GzAfchvs2Qw==
`protect END_PROTECTED
