`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ubfs0mXXQ5MrN8TF1rPepHnihAva2oOtWl1+52J95i9RV2cNYpCgPXBhMnJoOSep
XLfCvPH4xP7Px3eMQ+0Z+/QFZ7A8r9GeKHzggLcUo5sOYLtGUoQmCP31J3rB6TE/
WUN4f9QUuRXKLuBU8SSS8XIuDoxDnkLKej77Da065D6M6AFHhofblVcDljwBDCsk
g9Z+akjWTiKbyY8vMaLbvgS12eRDtqMhm1coV2aUVs0AMwS5WLj9JXL1M2VqvV5H
TINWOnbwLycZwMRK+rvnUg==
`protect END_PROTECTED
