`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8W8O41sApP/vK+5ARJY6KTs7fNY5zYGaFvwxCpEiv4NVDCmCtfSQjpfX2TdT9pBf
8qjN1QAaEsrFuru6u8HhJxTwCpFOaZ0veN5csycFVtTUiB9Qnlurk6/Mo2PBtYla
JGYR3RRQTkcvwBH5agkSuH7OwU1HvuXWkRHH5EmC6VkfVbtq2aDcjAuWbIBX8HYc
nKj7iVjz4x1RdJ08Gox+7VmJWKlFx9P4oSNSR29Ctgrtipfl/cTQiCa23A4+qpLI
xypFleOAQzyAxJyFYu9fw4EWDmoDxOZcuJbEcE1Q4cPAE6PY9Sk+n6BdyO/uWf8u
UoVuzqboUxrdvZDtBRTpgBqbv8kgh+kH/9jRTUprgiKx2NKwrEIOvbWc0MIAPYoG
QrMmf5HVJmJxgRrAUA1/uq4e9+/dgmPsl6aPrKc4XA0rdHEWGEgoAV1orP6PxBiK
9xbfPxPcIEdivY2HF2ct4uJ81gFFGGm20086DT8mo/n5DIKHFRAAQjb4oD7v5R1p
MGBwpGSA1ze+V+fUtDIYEwssciW/Dmktuth7YPIAhZzwKFEHYVBnDcHVDYhiVoeo
FngQrwaCkh1zrC00yH12WYBJ5dwfagL5zPg0aupylZFuVOzsUV9rzcVv/6FZZSTO
ASNeO0QB7r246aNNxI2xLisP7qXYpDCaom7e6cWVD70zLq/w9IAdpEWtLnVpF7kH
IQ/a2AkYsKgYRUOF9bYo3m/PzbArcuiVwc9eCZAHjNZiU5vGztryGVsoxW3KxJq6
LR2n5oO2OPDcXcjtfb/rRNmI3sDH31gU6XwymN5o1H0tdt3WVmmpNOSbfRS8sjpz
EahBHprzDDqYHO4IeLmVsv9XikqwWGDAYXqqoTZ0hK39ddGYuvKWpzUIjJuWWs8Y
VkDRJdUA3VZ94YYfaMKBPBu9nSeuF/rbvx3EP6QhzQZq94NJvkLbA1k/dv8HJMvS
`protect END_PROTECTED
