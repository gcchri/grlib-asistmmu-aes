`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1p0riCozdu4KuwL+saxMz5sIIZ4WSq3TNT9uagvFAKL5FMYLjBVSK0rnaWR36ui
PFYxS8pTv8QKauy5dvS/MTVHrcB/xkX/VOA/QZVARTKwCEtOMlLPTONzk686nOqG
3deRtKHnbpme7rmc4OAdsUJ7PZGHP1VBQXilIIPYgzqXTtf9Dzl66Vp4IUFXzHYK
+eHpXS6fxVgu7hPGHNqrMhyd/0bs5gHAo48QrqS2iG18lxYMMObjf3OYUXzE0hnV
eN46WCreIXANhskqH/8uq3FuhZr64ooU964HWoGYFQVxfKbmGhxBaLnW1B9dh/ZT
WZ2ZrvizAG5E8XtRY8nPkxW9/zyBo2QmH/1ODdNanoU1v5PcDnvER9ZR5lq9+Ros
`protect END_PROTECTED
