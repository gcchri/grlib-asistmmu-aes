`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N6Q3SkG938Qhb5Oig6qde0/5Cuis191J4atTNQRLNlIZdr9RlG+SR7UB78gSFHBL
QeMLtPhigg+0aiCyFdM93dID0Tyw3QqmTyVlRMwHYqD4fGtyyHHcBmVmt6BfKbT/
aArZimFVZqPfDAlipQmZuZKvEQd90yoFvdM2xkOK2DyHRbQfOTmoZeaNWvKOmkG7
HHgS1Ym+CFLeTze0RXUxbeXS0zqojDEXICwFKjiBJQBFgdTWtE+zjO8uKzTMlPKs
khtUxVH+slltmQWEC1DcuuO/Ma/oqh3o/7T0JepA76e37rqlU9fpSgp1+nwaZRuJ
73EsV16hBO/0pBdPufjv3yBV4SdcR52Z74KQ74C6S9oSZNYgHyQ998iTwl81CX2f
AoxF5qfYjqndb3LylFAttSSMdmUU+vfvVruScMMRn4E=
`protect END_PROTECTED
