`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hKiVzgBbz+nbEddLZ6H8FgE0hDwWbaq9FhZPG/npGaXYpBAXnyO/feEE8zfJy4Jd
HbUhA+3AbwBtS26B5sVYBLW11XRtjVHXbWf25GgIpbmKeE3KgPkr7hFpjAZiplUj
q0qYPZHyGBBb84JK+zOVSKZgW1gtW9BjInXaU7/4kygZ5KPVe3pGTPUeW9yG0CDH
t6YlYHqz2yxr5hG8e2u9E7Uq9VDVw6nLLwDuLvsESWY0hYH4z3pglVIyur0Y244N
s4WYOol/i4DEEo3jEfXTc3BxkH3xFBoQFuwq2haEE34mdzIA3n282tP2TCe6AmSU
jTwQkVyWrmAxLqh1Hzk7Ko28q/AMHsfqhtKmV2O+zERcAlDTBw0Pa3VbF3OjNFFi
F6ZqEj8kipSOUXpV70y3Y9aPWJbNDaSgp/DN5Nj1qL665rvUsFnmfY3W7nB7vzLj
GH7/yaeYl9v6wSNesWbnd51yayVG5e5Q2GomyqDi/AxjdoyhClwPlGTFZZ9Q8vMD
Rwn9j+AV9we6XOLENC8geCB40kj7R/zNAzjV3Pap7rUieSPRl3ASOCmXdGTuvkb/
Ri0lRccROctETPFVJoPvqew5d8QZ15dBHsR0iZwnUoEexmwJNQw5UaCSaHEYzugA
imnGk37/shPcRSXiJDrO4N/zlyeTb1VYwxsfPtNW51vfBv9Xpak72ZTwyTTxrPan
azAN1VYFboHZkCkpCOFYWyOJDYpzCtxLzNtw7m5+5x2PKK9JAabY46sYvJ7apPeK
xSsnkuaCp+4AnV/SZgDTO0PXvT4PRwnCwjGTGQ6P7iMYeH4VSb0T3x1kC7pDknvw
aTE7zMDysDvkUEfgI0DxxsrjB12NqyyS/B3mn9qbd8qyYaf5ovqFh33xr1q7Ydho
CZpousprTGeaSqQI8fNURt5B2DaYJBGKWoUa9C7Y1a8Nut77WONZe/fw6BD6ElTS
5izDkH1FLunMOsjZeoUK8pk7DRcs2az6O06MZuMmdd4QBZ7SkQPSrTihfOeKTg7O
loALPSorkkjeXnkXjwlG6hA6o3mDR8foSlr35DBAoBYKeTCrty3KyfZVWnIg7XFE
B3iBsbrxOBRVBdmb+mwr/YBt9Ytmpy5gAF7j6asqE/I+ZqAEp/oq0V02j52Jbpxj
yrPTTJNVpxoaYuISr7wvm45Bu347CYjawUBBEUR1NUN3zFlcKd3R8Vwk/+54UBic
y0qLEGJ9KFu6dBz8dH56gLqrvXJXLCablBBA1cKjD/gzS1Y/lPhOexu6f+LD8civ
QFjNVcoshgfLw3G0clM5a/Wn2veccufwX6fLWgev5ayLWnsHpU1TxqOyzEGv7oCv
67fGUDnYlUMTZmbOT7Q9khD88whgwEjubLLXRSJ4N0jU62Mhi/qnRyk1esfDno6j
l7diAJeqQ6UYS+vM+9uvlScIss+yY3X7hsJfE8714xfn9QgarkF37Qu/sJJCNfbu
lmauxsAaC/n5T2oVu4s/896d/NuBTU3nYPFAbCDP/d6dGgxJI4zjqwh4yQ8BS8wb
Z7V3ynVHkiIemLra+a1UtQkWP1eXEpGgfp+S2osqpYF8iVJ03B1DPUE1TCQ0vcsM
J6QSryue4EaVG4Gaz8au9AbvTFOO/nC7J71dNlFCkkjrDTFU0f02K6ZSBr3VLsj8
`protect END_PROTECTED
