`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHTNFgLZK29u1pF0+RUZVZv9KYsZSLCbCIyFjfJH/K01h5zQ7fTCvlCwRhTk1fa9
Pv/XhacSy2zSZqa4ZlHOrcctie9wZ/cwcyt1fzsyASaG/+azFQC4T3MVRXCTI8Uo
UqxD0Ucq7hnpaaI0GqRiGGmcZJ2JR9aytgi2rOpAR36d9VaSZeuGpLUMvrtHtZAR
Vqz5ApMTz6fXwkvsxN0fEoyJCy8TDKnYszhrRpC8chm7T+LYu+9jLBsPD2ec+fFg
OZLqhDtv8lSkdSw7hAv+DufD4UHUuhEYKliGZMoXUvw+NZev8GHStaU7nKlqFKgX
FBbgizysMVE0sPlUsid2JlHtobHNGjrZxGrAnzQI+2t4QlrTHNINNP53KjZzFtZd
td/AP/7PUg+qCdnoc7sXjMONuhot4hywyQDyZwV4Vgvpo4PNKtaIgMZ2eNx0PSAg
mKgFaU3BaybtvbkDvxQOsbZPdFp0pzbxq7pNL9w4YZfNdBiTGWuYefsFqgf5Z39D
NIchMik9fcytF8ee1RZbIau3UFpD8aNLL0vZscrow/xKMfvKqpCKTa0b/swm38W7
5GZgdM53mSDMLXqoICW3XzPRN/+QI76NOq1gewjbpPHea2vatfD/xkXf+qZhE61B
/isq2dtlqamAY8QisVTrZLm/C4zrHsMq7OzwJBD5DWg=
`protect END_PROTECTED
