`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KBLNdcdeu7ivwOjMSBTcq4xkmoeQEytGYn8tHiG1gBhz9y4m05wY/GNLotTGDFlv
jO+0hVwt8EfYVowjYqKKgJn5ErStH9DI+e81+A/k6Qr+i82mlXl2GJMEE6ulVDid
RW1u7YsHkaLm6N/LaDSqGHeNYJtwCZEgk/Gu3O2jwrWjMSCyjcSmB1TEc5+Yjgbm
zTza23FSfHbdW7l05rW6OjQ32qd0GGi8KMg0UQo0npRpQMtmsIXklNdkLOG6VK+V
ODQ0zG/wRiGZtP6duVWulpw4QAVS1bVXITeW9jPBegj0UKGj3calTmECu29vJC91
ftUPTutiTYGMxFV5OyabYMlqwNPZHbubRa0OJMKzeJ/doEcb0+VyUUzFz89d1iNx
yCEUviQcD6O5kHIT28UlImPTecaagFDvyb1XY5BsknTYlZp5d1/aqsHfkQSNtbya
9V2ddAzgE94OsntyfhqiHJ2T2rc3OukJXferv1ZD0WDgtMPxBVgboLQXxT5yllz4
DtJKDpPuRp76abmHQbtHauC3/PSd7dIFDbv82rFLdKVRWys0tSdY/aabi8cuND7i
Xd6y/v4hwUebLnBbHNqWOP+Fp4f6wgJYPz/KMcmTIOaO6kUCPuAGpmUf39k2l8il
cH1ZPWR/0KJTUcyQCLV5rt4Dk4X22YaQ9kozo7qoAiTioA1//esSnsBuTe56uizq
EDpKlFYDd87n7c5QUg+/lSLh6tHPDamTPkZ9GGPvTEHblHtwgiPB6Jj7+8SArD2Z
0HBxlBgNEyC6Z9eEfn5sTFrFt/fQwYajSyxig5/csma2u6E9uxldXLI3+j0dHW6K
7yUNJiM49CE9s/yxEAFRI9drsS97XDQvjYrmdI0sH8mgNAwqfFiQ2xNvNQ8a7Ykg
FXr+PsRq/7pT6O6XOobc2X3JwLM3ELsTWtIPmkVdQpD2oMFeJyqZu9/XFslQjPBQ
hNKny7ZEguMYRta4Q/9WtAccWztcRnyE3NJUO7HQlb0G5so/YaYHKoXTQLEzGRnQ
KQMs3isyc7Jm6xTol+FBls8CPG8zank3N2TsTmZV2EEdBZToec+HqVa4kDo1j9cK
bb144Q/x61wg0nUaudMwkAk49b5f0T8TY9nv0m48pthXCZa5G3iRhg36Hm995b7P
Ueh93Kq8LxldBr/8AbVHLKh8V464xoaDgZbagS81gUxH2HUo7GbYqF26sbmEo2GK
Z0MKrO38LQOib3xqoV0kDS1dNZz7KDU/rg1RqYeV8a5jQDAVTAiA+kqhujMkvZ8D
29nlNWth4nFnEjOrdEjZusJyVS5PXFCta0GqvXN8CW1HdNx4kthfMaYqnDDeb1Ks
b68UKhS5IOKxWoa1OU/95RiktpSfw6Jdjo1SNP1c5Wwbt9VjPzeTan5bDhZSA5Jv
WmH0xzDVER2OOJT1ZwgaHl8+oRaTETYorOrD8qAxLWjkGHDFRVXceacAug97BL4s
8u7h8WnYXPx9ojiPzIOXWSYwu1g+rYTMovfhPaeVwrTs7b9rAcflGlg4SFxrwRhC
jcDbILnkY9TmUFwmB7WxeXV0BGa8fsQcRbi0vOptLJMZ6Y1UiYrFhxsYY4aL7pqu
iXj1Bux8aj7eJ9Hk98g/HQ0P+c5r16/XCxhZx0diH2E2dqXRwqLqrDJNRzzyWv8R
lJEzmgoQgyZtqOyC3qyAMQB9R0PhTd1TwknGdJdKmcZjqcgQDDU0jhquyK5ZPI3p
7Y0rbPUK/g/ZCMjuSxw6E/Dvz2KydZj5iiHUsWPEDlf7EkN/em1T4/T0Tq/f1xi8
1tme2KNx3dqPRR3j/NoWYS1j/eBM7YeRcFEE+NDys1XIMPlMsERuJCzONp4HtjDN
+UeP/+4JyK/UmVW+enu2VQ/1aHXuR01VB9WwgrxR7C3GN9ePbk0nrAVSZ62fasGu
DrYbdjKDZmtAyMYspxjTJnyq0Wppz5ocP+ryvc+vNUpHzz5syauYAwxcmzaB93IX
YS6OPQF6lm6imXnB3GBRSxM9c/PpnpEyvh65bwpYTcp3LPJOOEjVd2LOFk4/YuVn
1gA1efcoN8VZvwYKioszjZZQ0xX3kbBEUcm5nfFOKwIbPprD5hbDmIAKr2KOnJbh
V2KfpLaMF1GlntIDySaF3BIOyUaWBcFz+w4DC+WnrDa7BNTHapM6C4arYSgg2QJb
BKdMZBn+2u3taV5qMAgdCyERxo2NSlbIu850urSxgMUd/4emEvz/3g4APiZ06qS0
CrpeArrJGfHmNBxXfTCgb+GB9yOs1yu90dhZ1HBQG+fxve634YTNRKi/ASkn9lMw
y3ittEAHBSZ3RSnQJcsfz4Ggf8AskFWXJtlG9IgFFPG2uiMpfopenP3kZG1iEdNG
R94vxVswxIWO+2oWUan3xyruIPPbyhN7mZYynnRX7VHBcPHHNYXzaLA2zRQq1wOJ
+X90xYfI5WtgYJkVvzLG/b1O/LJ2xq/Ndk4tCQlVk9fs8FUbHQb3+6M7/y9pVo3D
VBF3MuqmKpgFK8CWw0S+O3zCNDYY7CntwWXr6ydwgHX1a+DZre+Vfrm1xSrzo3fT
gqWFS/OZF3AIYjPwvG46VloQ8YoH+Vpy6avsYzUb9W+KKTVPT8xGiSp1daS/rpzC
2iyiKCRzNf0MdP/ak/J8Tpp6/AHH6JIYUezQI9Z2yGzAqEFI4QP/H0rfIvRnn6Tq
Img8Kkg4Frgm5CFfT7NWWMd674kVQxMNygG2T5x4wrjP2Xt/W3oLGk/SUXe8XQxT
iqA/4vwIGBd/NxXZkN0mC3iGQ8/Oba3i0LgmMLLaot6uI5Jf5ZIuGYvre/pLE0Xj
O0OUozCXATipWgqqqrqZwZNvv6Ow7JvZ/qBIdFYRFmEfJ+3O8yzrECPWUfLjZetE
/t3WOEOWAdMpJWVw/vLg1CPbHQJRg/5eqAuShUsf2ZeevPwws7KssoK6KJKuLN/v
tzQ036xjSCCG/XSaerL08ApBc7a/IhKxwlHwZWL8KwT7CEzN8/LxDHb0ANrkcu94
+LwLvn/SCr+iMEYeKjqk63b9XsvIdfhFwSNFqHoPxlj6c33pN3KtoDzm7eL62GoY
YYtDEZDahewGfyw1MWbLOC3gs3j3FqnYDm5JRXaXUDNMUXzXe3cQ6GB9H51HLWGE
KDMr3ttk48Mzc+HhvViJ0UCUZh4rr/p/Q8AqHLyzXa8uwdavzY7SUuPiqaK7mpBf
KNhriqZU1nTy2aXz4hRLfon7jS8WBQpPcia73qYCvCMNFbj6LayEoaRJbP7v4oZ0
U/DeMM3NN5VKLZFD6IgKJejyioFhZl03v21OFNRJDvcGAnUyoONXx7LLgmJt7Wuo
AGK9uvqTf9LfNcu64Wm6XtVU8yPQYzIpVNXmulKIOvyLgU4SAmITfQzyxkfQkm9V
JNRtXliCOd9gFUuBBzmLIC/fwD8WMBiStFiMaCLe3YcS30aJPKq74zGLQCcwmR4y
kvTWgKd3J50wIDIi+CE+0D0JkHOx0y/sDF0Pij/7e268RSzsmRFz1bBr/FKao/XO
Oglmxyq/czHtqQluach5Ql9/cY7RkVWDdPWx2bUX3iJDQk9/BNQZHvoCsEK12/kt
CxlbiV+PyiIZWK+M7Zn2skLIC/2pYUeih1VpCOAl1vARJk14h2b6n7tmG78CZ/e/
ruzFKhBCyjDiXYCMs6yoiTebNBjU4DteOflgNQzpSj6cdI0S6RYuqmN8iFjgUZKC
28KqbjRk9EWKGYoek26cIvArKYqfX0ho5pnmENXP7SuPkKofy5CqlNzrTViHOs6X
ovM6HA7wp0wuvQVtlOJgVIuBz6JZuwuNS+biUQVlrxNSVLNZu0kUq7yj1Or9/ZIM
jnKv5PK8zX+WqNJ9QuR+ah5pmqW2GyNg2rEPzYOMZKOSQt64h8phqcNiSI8RFGNb
wIA0ugTQDbADObmxrXsJtsrZKb99MIlUjbzK7ldF8KOMo1VAtOaRIbv/uhqFoIf+
c0E3iSQ8G5RPXXlcpqW9LaeorcOJUmJERldwRmbFXTSNT7l1iIvNET7dhcbs+8jU
KIs1/+As7GvCL5VKw2eQKZ/fIpmUiN0YaJvZXoXoEcNAe/4u9ho51/ObGiIsor4W
3SCg7SG3+/LHzyxj8QmKVK1xCKFnzLBuHtdnnMO01gSztHiYWng0yoaMqlChtb6e
jF4lmqNOK8l0NoyDVGxQ5s+B/YGLCPE49IWIKrGYtLwQ6nN/BkFQUuCmFeZUQfXx
hIXeiQRFyAkCNAopyrr7PcWwhlOdAybHxjdyeGnCEbUcxVs5c500q5CgKmA1c1UK
H2/eDbkY0ENR5/xGaR5tvGko84bkXENPKK+Tg9LWwpUk2jFzWc4OdvwVMQTG2A+F
TJqMFacl8xH9NAJUn8Bxc0i38v02sLl/6792c6zBCKaHeNtueoZxh3yun/KHbhaT
I8btTrinHae5HNyoxIbCDOZGyd9+K9WYVgS0U43R/PE7aWCWTw+YBd1RDsS64lSr
9Hj+RhPoAXkUQFu9RmBACxThRhINmbDNc8xDawL+SPcWt/DmDtcRgCEBDfXIVbo5
ozvvx8zLfd0wNwsKPfhBKqvYAHnFif2nWAX7hPo4O5xFIyLHUwEirkjPKyF318DS
1Ly0N92DfYVfDc9pggb0lQoHvQmMdtMLzoOU0HkU5lMZP0ZnXoIfGPKuXxxUnfHk
Bj+fNppoIPjX214vVy+g5AEXnJu4HkYz9OxxO3H92Kee/QrlVd/uCXrROHf129ze
/5tEJj2hLHi1xO7orWGL6CK8/vRIh3e6uZGGOB+Cb6CbIAWSn8jATYWfXPXdLTAr
smsfeFLQ8nBAGDFh4KeQDHQWGh8CP9zC7vKzHmfomZBRBwCuuAmRRa/jkHViCEH8
xoC6khVTOVS5m/ptBZpmfc5vwqGxO4QKZjpfNJPvPhXqNUF96mHYF435ZargqqQ3
CYco7RwQ0DbGJWfdFhvT7xaXJTzCMMPgXMrw8UQLXUl22gMRFxBUpHmzRQiQLW3W
V0+742nMnybog+RsMThsGZIGnyna0k2LZyzSW2RMEICqaAL9+jwvl+Y/5W9sIo4z
TnFy2oXdoaYjoDdxtNCjAXTL4sfcwjpHKodps2ozkAXAgx/Va5/aJwvqpLDvS7Xy
2wJvEVN4ZKiEG3KFTcwA6MpIv1CkOkqeJuCANdaAgFG5lhX8EwLYLACuV+ql2iXC
3pTEQDbZ98eb2aQlkl9lzIeOFwjtIv5yfbe+H7TDX9XN4zXjn/rQZhAy4+/inFDG
lFVxloenEVCLj/hBLY/CAWgq1XtnXL2w2WYCUukxdL1sN+pjz4YJz94RJWx9Ic/L
Wl8w3HI947XJZPcMmTS9oDQdNtDHB+qIkrVUnpTbEOl4u47yfUl/3asTRg1SwSaM
Ha9o19smQ+h6O8CXfklUPaa+zEF10lXRC2akKJQh/d54wy8dQGIBcZrX1CMznKPL
DTyC5nNI0/+unTXYtGFTflcJwfUPs7pMNVFHkAV0zv2ffnb8swWe2DRL4NJeo3HM
9YSlGPP4T0zHptOYqudDowfGlW9HhCBF5OaOMJk/+iY=
`protect END_PROTECTED
