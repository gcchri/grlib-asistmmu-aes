`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R01e1SuWymHMLW5eN0Fcq8+5fAOtgpufzLVMraUktxdL//LMIfjSn0BNLgbeDCkh
XP2JUafhL11trWssxxu8TsSh43nGanHl69hjFNqHMXPkzm/ytm19Vu3gCEren0iR
5Kdn1aG/pSa0b0Gwb14rQwmQEteglq+j99hNtUqZISyfolNKGXDCD1KIvlb0Du2x
kuxZtBsp/5vP7C+WJUGEvH5LK/wVfuWesW+rMMr1Vi2ZXHNfRsEF+AdxreF+cRpK
WFYwOqa3fV16clFggmCy4NhDwScA7Eo5Ru9ZAxwagPThq7pVKkyowCYtoAyxIG8n
KJ+8gAhWmZGUoMs4WzFX9AL3waarLuWxHDdpvIiNZMztUZA/ClvVWrb9AajoTLF1
srlIG77CNdQOOE07HHFxWQOPTLu6EMucYMMpBXk+alnOIPGG05YRPomDWfDhsZfa
SglRyQPL4GpPmMGm/pn2EEtqaSdqEwFmTDByG8D79rsZ5DgHA+I76P2vm6ZUGf21
VrMxQnRyF6xAFg8kay3uP0R0mVbudl3JGOLFXC/0027IlckoqHCyEiy/mk0tvbj0
sbAf6FQ8YxF7g51jcrarhieN57FZLoEBXFNr3zbsatkJJ7C/Qbnp8M7rI8wdMm7P
aAJbU7XyW2XkLO2NVOgBxp8+9FE+DRhkXUB4SnKatF5YHfJ50URSGMWtppQVv5v+
WsG5ww0eTZEyNAMxzBSGcMRlJiD1eOMqu3asHIqDOzgi9MhUPp0eVMR8Kg+3VprJ
YcaZZWc8JZuy7MyYC8pA+E/kV6bGSHnLjw1tkmJEZSK89upFIwiGvj3B0xALoYCp
ToBLDqjlRcufWts3EuPPYhgd+tbcVciojW3/jFyIsQjKXmS4BAIqCr8KcioS4kIW
LA8bhfp78Z+6PNYeAxjy970gpdhBwZe7Oad4aE+41hfjz38maUXqjIYaQpRkXvqL
`protect END_PROTECTED
