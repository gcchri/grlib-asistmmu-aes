`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
re/R/Q385FOvEEk5WsDCfw3oqGG4evSmTi0OpLIUKNE9QeKhcOVM0YStGPUgSf+g
GtoJZwANC+HQ2DOysUovX7bfWwIwZWK19wddqT4tf6V99f6iKbqVanbdiDGENi6G
64StsLjYiddtP/EdacCinAcS3+9uJ6ZY9HrGBOm/vFFJhS8+v2SkfguiU4c0SaOZ
wBUSUunAWEcWFAnZ5sbSO5dDCnep8uvLa4D5KVu1G0AJPl8e0mOhoxxRpGX3MHu4
mYJ5GjG6GAHgHFFp+xzKLFJ+CAx0L3159nlb8X1uW2M=
`protect END_PROTECTED
