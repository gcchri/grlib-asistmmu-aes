`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ecJFc1GrGFSwey3hQdIwxcJWfvIgbRzcIHHL2W58RqVyx81kXuSHl7RDnjv6CFKK
sL8akZ9EazUuKinYqJySsIpTqPhR15zuzyJiNhQJH8CbCBR4dwgALZUgKsWNrf9X
h6Bi8CbEgaQ6CbjQPXC0n8kSOLeoQgPOo3pR8O/4eEc4ZMubBlh2kZQveoJlcvWg
oZL7fbK2ePkXVZKylwBjAQ2xRzaO+9j/IpS8M09tUsEffqRBBDsAKuVYKnUQ8/SW
5KDDRX6o6RGeB710qla/RkV6X9PbUbe9p6vLits+Yu8yjl7y8UKIwdwO86hJzchA
alkheCyZTVsFGdxJKt1EkQnenzWXJaVYsi6pdME3vkRzqYOZ586OZ40iF4wf3Byq
vWGBHjksvzmZN59JjNy4PQdf7eaoCjd4O9E4xWMeBOkRR2ZzM4PS2iYhUJfwxgHE
uAXO/NSu/5pqrgJoDzKdgw==
`protect END_PROTECTED
