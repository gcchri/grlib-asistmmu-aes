`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ArrORUpIyInZnpGmpl5Il0MSzF4VqMXaK80KBtLN48ZYZ7gVXS2o5taV1kfm5cp3
l5TNw0aDd7mCWtItqsMMmNyBsn3wiAfjLnNgX/TMYvh10TDNwMaH/UvAtI+gSi98
ArLRyrOq1oiq7+Vr3CD4Mfeeo58TKVHeOg4Ukgm2+X3o077jxqeJmVbMHfjD2VNz
FrSwh8efXBaBLu7qNj93bpAVJ3qvPSUMEiZmmsfL1Lknc9sgQ2Gx/bTZDQFZUstK
0tYyZU/kpP61urYx+8jsEQ==
`protect END_PROTECTED
