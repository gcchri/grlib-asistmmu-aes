`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UwiTo5q6He4hl4jcEYJjhUt4C3Z7glyzpIAdYzA6wnnzZrQDKCNWQ0uqKKS+M7cQ
Tnf4OlTG2ClQkYZS0RPAFpAO3cK0oIpGCeHIASXL6iUYko7PGsZJ/Q9kjbeF7QjW
t0/fje+hgHJE+N7hjZY+IjFpZqW7PvfTHeUqmJdWU1i8xl/rvtPu5priwv2eut8m
K4PiuNgrtg0ITd1xLP2gmY4uNbXdGk0q28qH4am6LJX5h1hIkrd+zLcWbyuVdzRe
WDsB6HWARh3DaHlFai4CTLB7yswg3yG0+99KRmvtyqDdNAQ9PqU5wxWpE4W3Rb08
LE9JlK5nPsg7p+iiqSE5EiSB6JMKW/3S1f0rn2wSum5D4UUSrnlSo6eh1NhH+e80
TIZ6jSDHhLzu0L/jL9V44ajYCC9ma5M59iuuY+UyexGHybQu5mhxN3GtXmZOAHHK
mwETRtsaKw7yx1lybxtCZu+qADrZBUtwtIARTdlB1OCnQ/WhdIxbzAru9Z8rlMQY
`protect END_PROTECTED
