`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AClM5tswCV30XLiGa7PygBveZlvNDHEdPLiCT7SSYyYZb3CnIXLmZa10b5qXldUk
qF43+vYyw8oLVhPynVVZAKkVjL/JgOUQOJby/IwfUREnZOJXy2T13BcbYaunCAaf
ViRL5xEodW841SPBuKXSA7nJG5mjZsPSKForxr6X8PhALxkbGhvDqdiOtEXn5upt
uhMJR1Zxsy2pn2faA6VeQo+qyZgehxfzpy5o5YXDVo1VrAGmK/LgOlWs3aunLAdq
hX3kjmV8L01rOBt4JohbjcZFepOzrrbu3l/WCvw+SrzXPzEaXCoWd2CjgPwXOWtn
Dqcyuwss+KCmgQg7cdQHkooOPTQF2fIHlV2jeLSr3LEoJScDFbsfR34WTxpe/CJB
5Ezaeh0KBShUf6+VW/L1hqQP+Zdd0Hmi5Tga6HO7EUKgH0c9ulE1TMIE5m1t6K4M
Bcrt9Zhr2QbewO3spbMzk/y0v+aa4FfxoHqWiqWEZeAqT9CZTRzOKBm14qLXpj2M
`protect END_PROTECTED
