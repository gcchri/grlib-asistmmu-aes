`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bf0bBizezRbUdtwsieca3CRNgCgHUQjcpJoRIJeCxQLtc4zj5Z+DhZEXRkeNBDA
hi3Qebrv0Qttc27eArItahelb7nM1xTLeZW9pzKLuU6a4SD+2zWjJyqmkcUYxtVt
KWgwTR/J+p8cxVcbtnsW7CWEZQVK/zHBytpHCvG4U6Pwmg1n7pn3TNk/f4yewCu6
M+HY6q4QcrwUwV+uJjNda0fUA3qjbuP0i3t5fyeSS9S+biI59tsE9yM/og9j8xjd
61QfEuvJaROtp5+UCLNm+JhRdsr+PtekwYtmPIrcYiGlRku8T8x4iyzlH0fIy8+Y
4C7HYqllEi4LC0t4rN498QV/Nu3bnhXjvYj1YbOFzOwGnwVqqH1+j5FJ8zGDsGoo
8du7K/Ye5KHxWB1LHyFXPXOEOOPqdJ0BAjELoaExiUpz5RWlNK4897b9oSWqstXe
cHHfa+BsG77kt5K2tNuHmHHopygnM3t2fdd1syRp3ZAGcaW4eHgF6jcmWzkPNV4o
OEMBtlDiL27jO1o/GCXSY8zcHv4MjA9FU1PpB5veZneaCuTb1tLrbn/raZ7hquc3
ApBD68ISRbX9/lb87nhi0PUaOI7f8jKu6DR5ku1BN8wQXVSarr8nTzu9xIluJb6z
lliKUZfXFVpkoNJwv751O1p/zpoq1psCyo6nZV8pMH6ycDt6QYmi2wzg96HYNK1r
6P0DPsY91KqcNnfuF5QT70OGPjdsUkbc8AXnIgdBqNZrHZDDL0NKLrwVmA/U9Ir5
W/LNFeFlEyCfgN8oeHbS52JeCFAs1vvustsMcR99i7xSxOvUO15Rn0Bvz7Rh6F0k
+cWFAK436iCX5ELr8utTugllZ0MpMFcE2qol59NikEIdj5EInCErEipDq2TszjpI
kftm+lsv92AkNNcc3TuP2YpV8pkHGyMzJQIOWHEC+yKGbN9ZMOfgO3LabUBEzcgC
i9s1RwZKzYXabdTo+a0wSD6iP3pBsffISjRDSmywNvPiXUOysg2WSBS7TLAEWZ0f
ZOxiCGEwE7tmBYtPWNw6uS4QbZoydfuRDDeDruSmvDX4qwNi790cYMtqGiVfs/KI
GnatmUpu5HM+ilByigfnDZq8+EBmpbErurKZ632kjWSzcZAWywczex7KjIXSK6fb
Bp7CZuEqz3f5Wmh2XrdvQK2I3P2ECyxiq9l3FQWDy2gcRpR4nckRcygd2jlXAl0n
suG80NAIwJcxRkDeTdtZlD6/thQJiE732VIFjRR6CrnrGwpadBrnuTTeTmiUAAV8
ddpHf41n3gI5m6Lk4Buao5Hhl3eKd4yNOIrNsnNeUi2lRU9yTAOaPIpv8cvDDd4n
stih+MmKO3GgH3mnX2QDhpOKCdS8+qtQRik3b2Do8BT+JkkeM8u1waiWv+ohfMym
G3rLto3oBDtBELuBKvTaiP4ihOqEx2DgXMqmCLm0TuKGwE/ap6/faAT7wKOrPOTQ
6ZJsbuCR5mPu4Lkpdv+Ycu12N0OsDigsVNcWIJgAgwE1otxd7prb3txSNS9yyXYJ
21+ODQ0YzOD82YkrQSPuPE7k5zsTWZdP5nYeJXTSonHgle84cBvWDmg2gEQUEQvk
TGvetWhxrhOkNL6h6zjSicLMp2RssxTQ33HH/OO1lIF/m5VTgJNrZRJhjZHzQJrS
a2gly+e9InserHgZl0dlN/rUm5CeRO6Kv3Q8rV9Vm53tBap0UxGmvidqQbWCFRAA
psogG1OuY3FXWCL1uGHb71C08oWrZFs9I6Rig019gM8rCmQ1EbZs+enVDYokOTER
6e7XVBILfkw830ilCPHpkPeRlkFthHHVEUObys6xFmxmSL07IeIatDp6bg45fbkA
GT0DArr9ALxHsX0l3b7aAx6omdKr9kFSKFYWFou0XD3r4A1N+nDnDCzZCZ2ldWnv
Pfn7Z4Wnm/xuxkV7haqAGHcpNRisrvD72IwUdsXJANmeYBUg5pYXfWCTSfQxz2HQ
geeJZuQZ4K6s2jelRf9qxjTaKOAcstTiiv5JJWfE0SOBZTn4VIu2EfwpEqQbpZ3z
qbZHsKYXKKvvjesgFMx7czbdNdDx+8QhDVJm8/RTNjYMW9wT8sGW8PfO6ErsqSBP
qBUE4oTaq5oMOrmVm6HB0URXx9v1aW1Yrm3WqQx54lmRqWpVWKP+wcrOUrX4JUr1
vjTrS5dDzYDPY3/JXUD3OSGXj8xSZmzpqJeKt25fmoSUbUsFi9EnLqymi5M8fcRy
pjEUVsc0Q/F+UrD/7QdzZit13F7DuCp3Iuypi3Zt7TkZL7yGTcZqYkQVSPScp288
/eu9mPBtSNwEI8bBVJXw27qHPLbMoI04DjoX0a2WZP214aP5cSP8gzqvLM++2Eye
AEBxnFFqsRPi/PuvEz+FC2MusvJSW3d1Lo0Cm+L+EpJawohE1kj6Yl/YI1STmgCT
`protect END_PROTECTED
