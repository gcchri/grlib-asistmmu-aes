`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yrCR4usEsJbgcHALOVq7IO7damn/IPvyKgUX0tHoj+D4cmZyhcC24FP6Kv1oOG9X
aR65UA5HZ3hB3jUTs+127FYB40M931AsLvC5mfP/9mFyfggpnZc09rU9Oj0pLAQk
I/Vzz4gkCvpgk3QJVMHIaDeH4nyLBA3GHG2RoROke++QJeDEMGMPtW6IubcKPTa2
N6yLddyevNDbgS02UtESXoM9aNsMjI0BX3brZ0lAxy2dK1m60nsdun0RAu/hQRVT
X0WxJxzXjAdsJ7RN7eDQwAdt+lyRYHjtKvj5M69TbrTwBcaU5iT7oTKo5PedMs0p
DVWwnxmY39tIRjW4Ra00749bwjUukuWAXy657A4/hzr336qQr+6eaXX8ru1tR1He
`protect END_PROTECTED
