`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O4LMXyioWT+fQTf0YkW5e+6hdjztlO+zOSojQDOAkcV6w1eLGOxL3OBzxvMhMuF0
EuNw0ANRRBnzpE5N2ULydr73gnSF8KwGfPit24cX0i9S8t59YMYgF81C+xbs3L/O
0Rqp1pgfJGIOV8PEw7XGi8UnDlCKhWbjebafTYQFNl5mCuDuKMf/QSS+22hdlFA8
OdkyHHWpqZSxs4W3I0OhIGcc2/Ic6vRuEV5SLKuzVqsMFbh625CtL9jy2zNQCN4M
gjZ4QKlEOvGLHb3Qwe62rEI5Cy4pCkqFA3qteX0Bxemle2OHzymkN7HAxSEtO8xX
a+k+p32sj2ydfd1Ny6wnvZnYFuWJYWF8c7ijuyQT33Dm1Z9v+Kk7HzLx8emqEiCy
O2f8iusvpmg2ACAp8T6ATJ/Ccny7vqto/c4bm6ZGgEgWzSjDLxdTcHSaSRYbJwjL
`protect END_PROTECTED
