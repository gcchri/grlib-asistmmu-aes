`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HDvJBjxH3guYH3mb/NMrDCdIZ2PuCslWEveKznDClFHRn/iXRx5ZJ/gG2MZ5QRSb
c9wE4C4WikLuuh1vsWVGG9rPaCp6hXUBqSv/cJoYzfA1V8XlBEcEQeRqp7BYTP2H
xVeMal5vRZD8gSiWlNz+d1/HItHiifxPDuyXYCMDcWfavikrgHRG7/A/m05l4MaG
wWzO21aAZDl10igdyJQlJttefG+4K/79gmZfRIMNhmz7jTLcUkmrq96155NIo7On
hlpnCkOh115GUYZt26I3OoQkA6l0qFAnTpvtkgISVduJMDY1pLkCGoP1EqvStliT
CQ9qO88FSjvXv9kp97tbEzuAG7hcLgX0Q7YV6vq8rM0w2dyeQbsSQo/QL77xT4QQ
0BMjk1kI0yhy6Ln4Iq9VKg==
`protect END_PROTECTED
