`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqGomzI6jF5a/MkNFzFZFQ6jN7qE6oO7BmbTnegDRpB+AufnQFCHDxKDvXbigC6n
gdXAbopcVray9sIA016gK+wnJXUSLVd6Qeo/DLewbaoFZ/XIQLx2hZs1O2tOMCcB
KLPNdWmGfnq/8fQ6HQb5flE+GEX3oPZhPH4XyuqLvmGFn250E12Ng6euy235NoZk
VhDu7KvnOroU0uSwG1YG8a9UcEbi6KtSC/kXXlMu73HiAXwf1JMcQY7QLSKxR6+7
lRcUAbTxoRe06Ts9jG2nHNL+fZzRK58OBX2QajmXGxmpbKlHDe+QEv3VJRNZX9sT
GHhOd4VIwkVCI+6343Icnw==
`protect END_PROTECTED
