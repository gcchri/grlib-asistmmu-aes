`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+QgkEVc/U3lrMxRo1XJF2xxtBJDIkOkwlxkwWylMy6uVSMIUtQvYZbXJ9WTzXUb
49/6M7DUt2jim6GdsFXfGMMihMI1ZfwLEQt9EDqJooacwWS3Y5XrMkcyRQWJuSco
VUiOHAtDzlxH5xeol/SjhY7g7/swuZiKTHXhofFY8CS5Wi9TqpThFpSrUVYqZ+7+
i5M2x4jgYHwbXMV0VjiSU8AJFECuT+19ItBornGF+NrJsWiDwypZVQFjlaWKyVrj
vw6M0Bv91S/eIAr0BuKeaFt8Ye1wkzOX4yYSpK3MtRbJy6ExxeGLNP9eHpzBVTQK
f9NcNg/cXRHeysWsfpuzIelX/17uzVRyzmFsKPv0E73og8NqGdQ9rWa8VfUeAdWh
l6x2zwF0gxPmCX1jAAhl4g==
`protect END_PROTECTED
