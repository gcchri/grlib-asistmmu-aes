`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8gokXhlxoYbau/3na7pa8cwZ1IChayCpnuZbhMRm4TogZ/YQ2r52leVRrFpaNsc
QPg1sCGCIqwqOVNN3mnOQTWnfL2a7k7r2/3pGh7D8hPtB3aBhntgWto4WOgFsQ0F
hiPT1v3zuohdhX5Rd9MDsN5HVkk/QvBfbV5ZJEcGdykt2QJok2MXacsvR/KPcRoc
LO8yGWM7HSV7nfhzTOjtWAP+4dGPbfwCVJwCdjd3CiAGyEXQyw8l9xw5isdEpCaO
Wgf2nAfTr0fzdXlTV5cTG+gE/YELCihF4bWl2fx97ebaWCCV0/bZJEbgKLttJl/V
9mdVyFHjWNZAua6c0pRAgesBOQg4Z99Ct1Ey5urHgm9Q1pKwyXk2dycZp3peZBSP
338iHRR0TNZn/K+hubKMXx7vMIs1pwXsYUpp82UvHdP/w8f84YUvdVl5igQjISxb
R22ZeJtpN/E1ZZf6w6XrKmfQnQ5JpO0zKQXJ4QEM9rRwForq91OgOBTe+JVs/cpj
gOpdaJ7e76gnztMKN+QHbyvL1pxTr8B26ccn3FRg6djQOnkaX1m0y0CApNmLLMkt
Iag4wUiNthoeXXrmATAPlrXk7gb0HofOssBO2dfNQxVzglSZwlCRGdi8hhiWzJNd
zsCaxHzK31nvlQwI/4DCwk5x72PMKOE7LH81RNTcUAjfjdMLNaztuB3yGXQzdjfj
AANQdgiugKiTjKEHY6Xd0nda+uP2vraLAS8rkx7yXRhLHrgDaaXvnsCN9GUmfkQl
sikMRmbKNCaS14As9JwWROFekYNtuYNa+fzcpbt6HERm+l/ytxz4WcTtidbF9MHN
Vrs2ZxPhUkZCpUy+uuwrGf2o5y5SAn2/ICKtFpOrqTsO+LRUzn9kbqSurwR2p/VK
OXZp+6VYIB31lvwW2RsOniTvKU6TBVXOl5jz0nGzJNGWAjbArVIVg98TpLo7iLX3
pq7qj+pLvPntW0CkW36kop914JUf8alXykrcjcCHgl6pxd39QVlLXqcDIWVsYZ1E
IOh6YSk7BBVEqfs+F0gtbrB6GQhCDzG7O6fNsWvbhZEblTihGxlkW9O1ZJ+cXmTK
ek0iBceHN5fv6ZBB0x3eLMOYhLrVcBJmJYNhMPh6dPjm+WnSVkk+41L58ySFG1X8
fuwNxWJrsKkCqlOGLHz6sADDozhvLNFFylu9JGy8XtuPuChs3aw64P6YNaSFGH2Z
79G3r4tZgRBm95PRQ6loF1jND4IMZXMg9GJj56YBpfJftDVVOGFN68BS0+6usA/e
rL5nAtozgu6FnJsalNKN2Si+ZyqLg5juYz/+f8blw1CQJaNt9jEZT3GdN9y7vujN
e5CL2ErE35bz+EJLIp7p++Zo7YxsQbhPrY9mIFpjkAhdQk1i5fi6UYbOWcyuD/pC
w+k6spNHTIv6E34fIvqfZOmfj0tnEtg/uh94jidhP/26rpH2cyKbvcvjIvHDnLHx
`protect END_PROTECTED
