`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9CiRAZ96gwAdXyMfSLT7Wmn59PYZg9LqNhaUFFQnvSMStRRyyzGnw8cBBNDqqIOk
cqRH3eEVBdhXYLrBaR1hzv/xdMh/QUzT1yVEP9Kz+Rl86bn80LUnFvlJXl9fCARP
b0J65m5Ee/qP0OU0idOJzSUgmbNbFJgi0opk8NBYEQrvDAkUXeT2t1179eGCD603
n+7fFFl6IibJT+Pto+HySw+ByW2yPrtaGLTQRqkj2ljCo2LOnEBSiSfIK0a5IXFO
3dfKzbxJd2/dyU0y6Ff2HxbIwG2vdxYMl3KYIgkYUIrAhWg1qsP1A1v5bTF29Xzb
xC9/vf5alGcLc2R7LfpOknMHRG5DtNEPrW2Tlw8cWb7UF218ekt2CmAz9Ufhqx/c
zs15ocqtsnaiwGgCEb44MUTl42sxqUhJ/76hZ+YbGXXLc0y7VvPLuPIBEkHbcoCc
QbfpLf9gTHcefiTUWGaQS6XaIxldq1d8/yMDg6oZVVrklekt8qalTJjhHLRmWFlC
wE7fYPBr3jQn9NjTARtiVFrahDUeUnrUL/quT8KGLUGnCcKPSoD77PPAAd9SZxqj
Cwx2gLFNaKgO4qSAvKGD+kCetLuemUjnSdp+anbfFq8ATBjgyVQIvgttTHCCuycr
dxT2oFZs5qWCUIsDTSDppemReYuSE/n1EOZkU0mC/Xv/d+ebKWxyHLmkx6ce5bSL
ov3iLDW1pUrI2SS+p1Vjj6zcqZCKSHjamws3ctK/kQ4=
`protect END_PROTECTED
