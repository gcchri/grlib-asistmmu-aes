`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1FUpzZkCkEvbS9M6a6f+k9jxLL/kX0mavyc9ocroluUhZeLFiniR3vdpS1e4JQWm
tCBkDRRw60I1lHnFKQDQgn96yq/dfl0zZgswYxhGTSaPSLZx4FjYusJRkDjf4HT8
lLR/iT8dWsu47hF4ZDmjxaBnKccq3kJZb+zcHkzRbiW/mGegMbIaxgnD//9Ou9c3
CbeClevKvqppPZM7pAnG5WvFilH3kwk+9nhfT2OpF5XxbCmivK7QJdxZAQRjr2Cs
ky3oKfGb6Nt5FGAsRIBSsd3SKkCGwDttPewTdNiR+sU0tKGTxkcuIDqoeRGhgOMB
`protect END_PROTECTED
