`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tvi5iNc3QOvUVlv0ZHCH8+0rILNd9fLEU7Vcg5PjtpXncU5ok/bOEaRThXWPF47C
F4ozKh/RsB6y5ADNjYBF8f2lB9VJezHwTCGqDbqtRwEQdbjX0Ci/th4d/1rzWOpX
OikOkZQRUgnPbG7RKs5BuqXE/1IPOQrffBSXJ2xpq/gYWMwwnWSu+D+CPOwh33jr
gQbzlIOnj9bSW7KsXxy35mrl+cpPCDVn9UNSWHrNsrdDOz4vCILU1o587rDwfaER
CweUG9fg5VtjKgSJvrOgIJrLvZjguu1VzkX0Ewl8UJgEVH3Whz+iTYmCBOVWq6TF
hPIx/QFYJz6ONm3vkebLa5gaIufmv8xm0ZuC5yQ0IRdOBAThqbSdsOh4ZMoy72n2
pNS5FwPlT7vM5bb3AgN89x8QYXBA8oKX/6fB1zRE7txj9O1BtW3fjS0Dysm4ZHk3
hHX8m3yMjDQEeyPD7llWcuEzp/kZdxRif5CUuK6CC3CVsoh453kFvdAoQgc1H+wc
fUXaXZdxBiyx8pdlAr2BGxU/ZeKZnswmyc9+N6QxNwBJ6PrQG6YPGTNjHPn/Oc3n
M4Ufb7Q6x56ytj3GI/76Q12gKHATo65RWbejyeePu8WuSRyrvCoI3DQ/WVSte9mv
5Zn2EyKG7fHHapsw9OE+JQ1NWDAq9i7itBjOiyrxnx/Y83LvAhvVHyGVxTdFU3eg
RN3bET1eS/uHYek8MfYJyROrenT8iaSZku73k0jNiz1feM61x6nz2hRw25gZtVu1
zWBPDkUotQf2u2UvKWumgenh1WEVpcIhi6guce3n7HgeEhNgkoL10nXO41yDsn9e
p94EhudmVAwVMSdt6DYrKLc+2gVfiijABSPtOxy240nn0AMrM8oYHDP4xpkf+qW6
+bMAzE+cKXyQyX5Wfkxg6mCZxCnwyoXp+csK0rknPW2ursfS9ZE+rVUnhgHYsZdd
bJcU+Pn7ETrshrKPpEDjT9LYnLxHI+lEcHjRl/aZLXqx1NbXPP8XayuQotkGimgj
W7jn3ZGYKKpJF2X8RYbdP81M/7oAkApO/i6B+H50lEGaV90ng5viq0tGKzSW8kxF
3mvaBjZ4fS//Y/IH7jR0v7A/0D/KB3NlQ6EOudFcb9BbJwmy+qDE5VWwYoMEImYJ
0nTdh7Nfo2TcYkVVLcnigEqdiODOMEJZAStUUK3yLpJU38iyrQLZ7Nmxq4LVekrm
J8o/iqrSYnZLHMirMMHUlLmETGaKz0GKK3qnhZqqQ5EiwLG5Pmg54MefKkbhGcgS
60oc1N5jbPvbyuF6UYT6McDRMW4XhjeeUQ7iTjrioqomk7o0Q82FafyxOOpN8a0Y
ucOZRwa2EZdwBXCRghoDQPspEGQ4KADXObHb3E3RfAC/WpBD3lz32J8pViw3s6MN
ogLB3RbNDKM6eBsioETJU02rT7GZ6DQqC8mSDOm3+6RQ/fArz20L9WbrERhal4Kb
5lCahZVcEcQ1fG4mp2E3fmiTWe0jeOnr1oz0+xdyV8L1DCSAGJsCT7Pjta9ZgtJ/
YHqn4/1liOkdvI1bWGWWhcIEEh0YBw09ygK9YggOi9SmVRvrcSi8WDoxj1Jq9f1K
a3DpCXVPKh+88pDv6KsliErTA5WirV+EFE2qCn3P8QL6m2Dlk4yBUpFZea5Iu0kc
EwtgCh/M9NhVktfYfI66u6PywgzHcY1APjehF0wwqQDBpqFdP7+gwXC4XyibkLtN
FPQJ/7ILk5ieWjPRgvTXTSCjM0MGNAqDmqqiScIgYhhErFJFA7ReRB9d/q63ZP7/
jPVpC34z95UNvFhfJ3hMqP5ye379Q9+kmBytwJ5UMjgbacM/qDsONi7nP+z7P3Cz
mZ7NGspGRwc/Xla1swOtC/3Kq/0OZ1mMH1LUydxwA8I=
`protect END_PROTECTED
