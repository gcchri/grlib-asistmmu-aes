`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gdgp3uF6yEn01VM2SlCRhnngluTOsOwLBHf+DX+m9b1Y8VCxfu8IZYOhypYWKeYJ
6rLpcUT9lNrtrPZoXxL6gnyymIAgleFhVvQNHds1sHVSjHdLCP+czlS4gc977Zdb
Era5Z3OcUBPU+CX6B6PwItpEY9t+7t8T3ZB4D7DkJ4zmrjgNbfzZb1LYjqObEGyn
eXU6NUQMIBrfr7NXTlJe63+kgJ0PHSHJDfnGfwBDaJPin1XxHacMLWJIzHJIubfz
Ut1GiLGB3HGjvLCkNUD82tB/N+4Lj5g8nYyit7qVnOUc00U0LRXlcmqVWv6OpV15
293nWvI+OUaBF9fE/+BQ/PkQsNSQy10k3PlsEHt5JkIsBujgIJXUZ6KZYQrxVHI1
VVbiPjVJW/L4VSHWAkAAUP7oaNKf6QXGZhryTW/DoqS1nN4TE12m3BvesnKIZ1wO
pWVZLcL6/QT6Y5L7QmeHcH4yiFq2JMZ2SUMxLnX3dSr4YmaCQBrME36oNy6Tgmbe
q1bZ3/COlBQJ99SqIc8S2H83LActHMgpC8WZN+t/5/k=
`protect END_PROTECTED
