`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5r5P1L0Ob49LUuPev0esEL/IU4x45owgQNiaI+kdwgT8X8SHXgG3U/vGTSrpqkf9
7ZzkEmXseVFq86ycbxcdjTX8W2F2TF3zgV7PWHhpwFr014V4FboubBrEP+W/gDCG
xHWrZa+p8RrkEBMEm6mojxfCXA/leWPVhQU8vR/41oPGmI8qLe9FdX6Es/13pRM/
LWK4pzCIiskPTUvaLkMJUsBHL/Acvjs5pUjl5deKH2KDWTd6vZHROSH1O+mIWCvB
dBHb8RSvdqlmvGjT0q2QkO6MHL1lkKF+H7LTl0wC1VoIKepal/1kimKjHnBrGz8t
mTFPp/fxM3kzUGHUZCFEkv4SsVTd9haCoFd3wm+toLREW+XmnEFoxOxENZjWPZb8
uUIQyThlmrV5ra4AhqxDk+LmYFc6YaR2qabYw+jcObOcAIYnPXAw4U9rIqsaBddL
AM3SCZI9UCNG9NJcA+jtA4WwDF3XfCVx8v8tHHnEtS6AZ00R+YyCMyh8osAXE0sM
QGddnRAIJXSt3d0jnhl1GEeHLPkkAzVr9ROCsuiYI9k3rVIKi/Y6vQvvjk4do40E
86s63iwYh7EXsrKodwT8CP4b7HeVss2gU01IbPOpcp6L4Uz4WpjB0ye0Y/pSOhTW
KhxiuCS0KvUg0aHgDC6Yr/d6DIXvxQDRPoZkRQkYoEAa4X4QslXFYP9jo/jVEARJ
ef72f5WDlxxf93kSQa0tmv+vVTYNKIZW5FbVNlE8UXGPi8tSYQQqba2UW9YazCV2
a/PrIgv7oaMIrftEVM9KL3VSHX8PlyjLL5y1vRLXbfXhfSw08KOrxHvNCKPCo8ul
186U4N2k+qpcKucxX5Yos9Z7EH8j5YvQhkrwAqCy6UXXhjOKNjjllhWlRhHJtEqY
sSGjs2gTnI2ITjvg2A0QWVEGqb/IUHF/g3Ygwz1lXA7HivGo+cVTWsPk7zDYFGHj
5cP4BCkG6Q5kEU3T0wNiwdb2qAojM0mI6dE/KqePHTl2DhrBHJH8KGBjWqhAhQpK
PvAxnx7xtrXM6NVT84Mj/Qzy16SnS9vvU4A3oYu9en3VYMyB3Uv7T7BsccaqgyZP
/xSJk4xohFsH3A17LV17jdtSfRWbX/O5Pa0c49a5zQK/oHeqcL78dW9r3qwbp1Pl
cUZ5ef8xeWd9Mfx7/vBv4iXmQs7sJYtnhPGX/Ss9f6zmrXmrYTkTplQBpvDjan5A
D5fpR7HZ4RBiLQew6tTglKjleyMOFU/hBPAGFsujOghYfb23DYDkh/U/loh1aiCD
WD3w5pRWYNNzdFxXov/Y0R9kpATEXZr3gpIUUiFKCQ76lL/KuXmDrvVnYWnFKg8f
A0FMiUmtMSHY0FyFx2hHMgMVslzVlDt59MV9CFuKHWX8YSwygiOf3NANWG2Hh4yN
JfI5g12hLoUevqhkZfBOcJAmLXHqHCKBbOJMldKNqv7m4eB2noyqCAv7rNYr7Qdi
WfvulwOWHQ3dc1ET8rek6sWSBcvUk+yj9hlo7S4gANp+pyO0LZTD4JklkilcfvIF
sA12gJmR1Wk/kE1hKUGk/DyE+rZsHc9ZRY6VejxhtCNF7HV8yuqEXxZ5dmQPamjc
hYvjIWN1ExqY+kL2gDKdkVBz6lrjCnZxWPc1vevWgzCw1ItFlIIz+9uOSefym4P+
4Oak4TJhIjYw+483mshCHXGGHXf6V4H5sta+YloR/7fEnbOgBhMsWJlHpkoIfqnK
6H2pI0mLr2PaJPzBamw1Qm1Q9PAgCd+suza5AzN61YuSlcU1sSmepOgxmgFoItfo
8oxqFMKX0vTFXfzqE5v8JQp0ATmaBv8zm3fg0rMm+2I2zlYQ3PP6n1bw4qPBKKxJ
K4S2FR8HyTj7Z2jRTgX2dXsDHXSx2wjzzEVXwbdaAN5d8UvIgxUEoTB+ujkNPVou
4Aqqvr1vQ7nKdrioplM0IYxQHRRZtofwchBsv+/8de+GkmBxseDknAt1GK1o9jl9
K1T60Azsyzcsq1JVVAi92uhl3LSSH4Mkq2B6ARC7U1xhPo2IXlKU68awUmPrSb1V
Q3Ro28oiZV4/FwUY70Xfww==
`protect END_PROTECTED
