`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WlgH1OZs6D3AarJCOhvyBp2qj4TY9Fyq0PejFGSZXQtPUf4d9f4CokbMdvNfJ9Kc
/lqH7Ime+jgDznDREtua+P9ca/VFXDh0L3e+xGuTegjrtdjRfewAr8Zwo3/O/jSO
o/1IxO+5W7DiIE9Xs+P3uVSAc5KtNyYl8bPde/gcPY1b/EFnEaTWKzSKPtN7/QxF
EmnUMHP4TU46a958Ts9MPWG7ACPIjS/XeWtst90Dq/vL65yu/2+TbzsxX3njxqgC
uXpQ7uJDIcDzXqTnpVBnLC2vduVS6JYIvbT8NSG8m8E=
`protect END_PROTECTED
