`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mOilUXM2PvVP2y0LjgoXfWOGC8sLS7loBfpjxxCUlIRAw2WcAzSYNWRYuZhfxiFP
M1qRdNuXrEpMkSj5qoyqpFmDDtk8mj+b+yPEGcmXUURDYs+zYzuuO5M9+y6wvLBc
S9XJXx7O+TFXCCUD9WjA/lVh1sUQlmhxchDF3qNmgMXcDEqLaQGYKEy8FwP67ncV
u1kPfxxdeSfv2qBOxd9dEQK0z1xFEElU5hTDLbi90xhjip+hrccOo2T5PqYFUSZA
CBOOyCBGCwwxpWv4f4sBwcz1Qxxy/LvEJOx+yBgI4coKndr1mtn7bq/iFQ0UmMKe
kTlS0krnhAm6mXtYw7SWHN3OvDBi8h/Rpc3do7B/lgvmnAQwt+DaGlj3Hn/Un5mD
kV0wMpupCj50112pTugym4LVUQ+FmUd/epalpUh/G692Shbq2aeUjSeMCgQ9gIPI
sNDDjD5VR4v5KU6RwUFM70rN3BxD9G8fNNYyZHuGqsBnvqANeTEfvjCIFY2hH7zN
`protect END_PROTECTED
