`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+RS624AbkpsHHtfJ+DGAxgocxfj58r8QeSwxnz64qzcwy8njcwKHs/ZaJqfvodu
DATudV+Z86y3WDrXN84kAKQH4OX7bXlK51EUbVT/Hb8cM9WezJHkr1n4TGzb38aK
4aqZSsvfPSW2p8kiOHlT3VErkHFRHEJxzTjVl99pnqFZKa5f94H48RCi57P/R5DX
FDQ5hW1q+RPSspdeUsb5uR97Vl+L8UznPyDEJ0K+iewlFKqAuUO8E6TenmS7sL3K
Ee8od+5xXR0Zvg/lBR8IwFKRoFATws+B/JDFFpMgITTbhtUf7+iQPm+Js/TE+iXN
SSIa1uP3hKLIXJ4PY62LEbfgcsAblcbVpVviueaCrLNHByBlUzAvgTWppMs98EVJ
aLdU9/RHcPAitEqvVu19Ybp250XhJ4Ike1OEuDxS7omyZbwUEBfRK7Xk+5Kimmr3
PZ7oVemdgjXgt5RuVt04FjVtzJWn92/eCms/d/Ym3XSJ3UhgCyxut8Ug0dMxt85D
QenabBzPmXAYM397m3O49GbPzK5dpUW3eZW2vr8TugkRgzqi0gidrZDGYI/Spmly
33hEERYC482/2AMD8eP5SXl+UTsq1ajinrBnYMknWBbBx867TFjLrRQ5F6lcPyvC
H7wJG71pxos3O6Jk4+lP0K19L5wlWkJDr6yksa2mSJU=
`protect END_PROTECTED
