`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6v2kJKJ3BiRYeVbfctkGmSlbvbR4UToyi2b/YqwUqtxRVyxMmoqSMZvDvh4fOtN
4mBPCj3EEw6S0s50i2Qv4WMoMlxxpMho6qV667M7igf9kNHBSPWdcIAldmYCcAZk
CXpPFLoz4cxnL3vRigt/4xTG3AKcPxYGb7neq13hb53hHrOlkQbVyQ9BqA40Ql4h
5uJdxpMtCM5fnmpJcnHc3S+urbXab6JDwZcs2AOa78ncwW4M3vqYgp1dwRPDUnIy
xht9igx41DqgY/Wb8Eh3CFWS73rWlRuPHjgnX+jRLHdM82p2KTExpOk/1aEBI/gb
Clpub32Qb7FgWteSs7JnQXCYYcCFVy3Y6fF/QwGiRMRcr+b8mlZynKtSvro67xf0
de0qdhKAOK+fbYFjvMvWs3634lW9FrG7yeAWBm5MVkxzlz3nGLXDTLHGBbWBbiJL
jXowJxc2QSVCYpXeybtKHfxsgmbFVMfuyxBC3kwUDsAJoN2x12kUS0hyF7oQ4lx+
N1Cs4YhXKg2BSI3iFCymuh6W2Vv3DYml0PNoy/ZjJoYfmw3StLsW/LYkNb7d65w0
Z+KuroPALeN5FlFHqQNEfLxCzCGfTlmgKsjMnrLoLb26Ue5lD/TYe+IJu6i+yNOw
sB9FiwEC6JZrl4cWXQ67p4vuE2xJQTn/N24cFBQRJRZ/OMgpzFSmXqCX94UPol3/
zyWSUh7e/sJq2VLX0dCdl2X5Lu6vYVWHSHcuQmiSVauBOZo09kNAit47gImWe8xZ
moQmQVeslxVN57CQaV3eFMIz9SoSG0a7cRxvGFzeTvHQuoC10X9CjaiJtFdIVTFs
GhVxD6/skXd9b/qLtMR2VW+NBGc4ap2KLI1YsePAL7Ec5GYI2StRiYtL/UMKE77P
OaQJ/C8ctemCFNhbo0VKJFg9vceEtD/bexvEzQvmgXHuW+Odl8GQCo7b/PV6sz9N
DeBnEe2pwbqyTgdDmaAhLYDoS8Ap8Rlkh+qOuEnPHXBPSfzdozFWGC1jf9dpKDfJ
FqXCJp88XwicI/u79jPQr1Qtthzbo4qCksflSKI+qW8HbWGMvzP27cq9DexThvPS
kQMoIztkE9Jsk2RpL4k03Mx8rCDRJ3di4gA3gtAeAa5u2H+T+SRG5PK6IUGLIxcx
rFd68kZ4FQUv5hRTRRb9A/M1aejnJ/2kaFJK2rrFe54/1Fb82Eu67dZSvP244cJu
Am+XibsFdZDEkQJDiR8T9OQDR+7/0q/fYLdev6cg9+zghU0i1os0+Iq1cSiUY+p2
oo+0+KirgyPGzxf6WzHqFqTlEsvFoVrMpulLqXQEb0ek+S7LqWluUm7/laIwPEm/
6ti5dQO9ytkZPT1ZrQGdaN3pla4PQ1yL3luSxg91gsYib9Tf+T+fZ9v8n612m5f/
3PEUkBFdQD8kzNTkaWggAshH5Qufqc5dA+VhZ9C9cQ+/7jrT+wISuDSVjHXvhwQ2
QkTSyDH5SCz1IWrgHSM4C04WPz2KMVXGpfkd+Uiz+GpnqF4fGJaYa1w767H5kxt/
BXzU7gSmVg2mWL0A3GTGUWh3D2XssnqfqoZ1BR8iDX1bOB1aQ+i1nkv6YEshIkKP
cKTxdJIEWtXQLT77S0u4UCbgJWdANaROw3q2GKVPkpG1ioo+n7iiTiT6elY8VrQL
KEoDCxW1nBlejf482U4aa4UWtBOFDFPBJUjcKZwln0vSKZ3geEJp8jQvsKY1dL7p
WWkKHvz5AFuLPLGcMX8AU7nwK/va268+XdezXARFtDcC+dok6GWIYOzr+U4svZFV
uqM6zJNDlzw9em3HYpEAIcu4evj1hzJthWHqVCW4HiGCLGNSdQbrxDhCQFgftWGP
KMmy1AtQM0G3hUIDS8CA//CootKHgtPwcSuVIUf2MC0nqUHlTKTMaukyf4y8M14L
lTRPwYipCHD2r5TpcGznDIXdV3skClJz5z2N4mslxsS0yQYdhaRIZYgyBVqmp9GU
TUH1qF42SHJGSx1Mqau5SUvQ/l+Whc7YUncyBRXhO6b9G8ibakgpY9IOdUf5GB3B
3fq67JHJ/NXJ9sPO2Dcjxfv5EWpyO3FobyyD2Xg3Vs2HNvf9Cgp+toLkp6972EjJ
/BWfRj2t761awgrclcb5DpasbM/zMUfFsn9krHwbKl0Rm9C1/3bQ58KDQqF9tOQV
LB5EAU0RBIiYcZHfMLefE63IxPyZtFGF2A2BE22eQ2xOeA3n6YUTyyh239WVXmGi
QBzuJGUbsi/VHww1B/u2C7zdi7ebURM/29A3NdWuEvhPmbfJ8I/FxsBssqyZsT6G
6jE4amVoRy22lNbb8q+cQWd7KTvmOSt0WctpFVrbGPdAtFTXHUqB5cFML2LL9Ts/
hkO72FYlekp98XQZ9I82t+daw+LwThKUD3/h6TJ8JWy8qUjwW0Oco1R/NhrZrRKC
wu8En1i/oAdtQu/NCUrZ1nkwJzC74YVBNGGWGW7/pnzfKPm89csrBmcj/VKtLu2F
Z4fW+2WTOtU1q2jTgq5bpQbw7S79sJvz32W1bYw09Al0oyNFxwCJwMqpUF3j6tUN
Xq0E152iA51qW32IH5uVigdfJ3PdK793bHlS6MPHRrsWf4DJXn7lmib/PE+1RBIq
n82uElrQXeYJdHFfoz5q/ZIHRn8sCKfZgwTaJ9X3DXyICWXM2YlzBCR6QX4frHHI
ibrpRp/mkYsQGxLybebeACwcZS+gCZFaLl1WpJTHSpzIIfH4MAjKNMSS7K2h71bf
LYYDUg52WgWnB1bg4uFDALyPm332MfFOJKlaCDJWn092KrtlkX17Glcdhy6y1MWh
vpLa+QAS9V8R9vcmajedi4r3k6icN3ha18UoVC3L6SxcOBpu9eAVz2aA++SfRe2e
2vkoI8b8YgZrCNyhwtma/n16gGu1PFM+Hy0QR8SCu+ik4gRqBK0quqhR+wRKI5VY
Z5Z4K0ojJFC2+QxJNg8qHbVx1dRfzGjbKvN76jA7hfsdfKSGn8KNBajEJdDKIlvT
WV2gSJpw39FFx4gk07ZmvfLR1toLl532udsyr1QCZQIfZ+Wbh//KjnKpbUpsZdG4
EF0NdB6tlQmwn8OGNXSyKDkZ+uNLijIjlX5lfRSbVhRsxQCN9QuTkM2TF5dM3jbu
2ENZWF3o4iCvKWJtcbUW4q0wzBf7hPNKJvcwYlNvgq6/7VhCNEXp2ouk9XGolHYa
5/ihAUWxGRaL3Nl1kBsKaRX7MJARkTYcTurPC63L5wnebb+/W4Q5OHeESRlDwvqa
529+Jfa8GZoCFUQaD7SBY2BCTNnohnC6iNk8u3JFSXU/Yv1fUS8EtSoGgI20khJA
OG7T3kl7AdBl6f2d83Bu1j3vaTQ95ldHkWZM4WABwGsC8f2A93DSyUlBTf/998Cu
cTeJ6L4X8jK4GL//ysvYqLQfOJC7SgG2z4+uKDc1Gfk557KQ9zmiHwab9fmER7r0
BEDIw++CKxeGSSchS5Z1Ok/nWcJiqfM5a7LbHjH9nZnvSfjRnM4qHGHNc9WdGg7y
aHqZYsR1RK9wCBHoam1upDHOFmGmBTbu5QFErdC0mK7AgT33HYNMabHaknlSBhIn
oJYJW5/EP2a7pH6hDxWgE503R9jhV8IRwcUlZTjjpCVWF7D7AdiJCEWR2/H5S1JT
xLUiQOg9TnbjR4wtxZ4/nsUYlnLXSWOm8oUTqgJA0jTs+XVmsuf8XX7zU0oPeMPr
VDEPeGCKb/8VWpwKQjXbEgy5Sc3U35VVqItbQ3NAihyRVgAAIkXbfq7D0us7y6is
n6ByRmnxcNkDHI6Fqufnqmyi2wwJLHpZofdF1jyehaBV4XqUxNodL1UVKNJ1WBIW
8ZQtdxOMAnV5576A+h6ezcuVkQjwvI7MhgN/L53l8pCC/IFX/BjO1+EyodYUb2tR
f+0XN9vu63/dmLk+REecW1D4AAqy9BNv+d7SCYyLVStnkAIFFF4anJJNLR8BH22r
/0G1kon841uZQzutOeyxaOeWPMAq1NRIQlcnwHaCVKnySzuYVkkr9VPuxX/N81S9
NZfFYsIeo4fHbGpc6kukPyc8dqrc9ucD4j7CXriC4aAMJUOiJBPoRm3woe7uogkC
6/1aawhuAVKoY9wptkbg1l/XwOG1+nuN4TRlh3z+2BeCS0M/ZvIYeWh6TozBymF1
syiEVK5sipLzMoP0Sow2vqWEArpZ9OcWWXMzQAGi1uuRTBOjZgN864dW+ehhUMAg
6ZnO1Z4nTQyDBXBDMQLzry+M+RPUcSLj9Ql1lktnlLpFE4t3N/LvOL1pfmtBPckh
zbYHxI4/neRcVZlNAc7qbhTMPiFmJNn6+bhKM9qac8Xhs4yNtWYzLscG8O7QjY/3
m6wTDbcYkapv6hz/8t5I5Zp4ohSbbgz+XDS/6h/6yDCPzSICVtjKFZ4foxUxd1RK
W30ZvCFfwMRKCSsmGWl/jsf6MGbVItnnTkmh0lt2ymipkGIH/19Rguxxomn6rVcf
SftlOCyZ8EwgDKvq9ginHSZ32M4bPrvCJLWO395VRrPrj2xmXCjD73UToJPXElTz
lxC63V5bqkYXS8zDyDzEpzH5nWkMEhMySJ93bHcd6Riq42SvXxTrhKkaTaCnwRcP
g2Qc9asoe1fdYeL3FtWTkQe4R1RqfS6wbr9BNES3X/7InsOEVu7Via4BW7qzScEB
yjSZnsCFi+Qwt6g218bHEzaDPSc1s9704DCSMtSpDfmML+mvI30JhFZyVqJNwwR/
72m8zAaK2IqnXTOoqa675ZQop9QwCZkJNaJOkN2ebe5Th6r9MJQum6yoYr3eL6Sa
qZjbGQgLhldWwmzxgVr+dl83yzDIkB3yfaJVE25YOsdOtYpkQBL8UfhON0mZ2U7a
MtJpJLrR6+woRPEq9gF5+nZ1znC3kCcXJ9zMaMJcG1E/ftuiNhLnc0OMlGB+u9UU
5kCUBQcXROu8d4X+/dOyJrzUPgvxhen0nQFwbxeL8fXenT49GiYx67vciRfh4GBO
6rtvnkO80goWzm3V731NS26D6JBBAANCFf14Ay7eTEnqJEg7Yt/Eb7CJJtRpwlSb
nKDfYRNgH/xcVCp+uHDN+6pfc+X+Rzh95mZKjIg2VLuolu8ilD+g3CI6GccJ5gMc
iWn6Vj4akTfCJt9YHLIsW1Ia8/taPV/coudHdRcAfjpv61g/cDYp0cl8L5gh21yy
4gkMJSj7AVMik5dH71ASV5XtS6mUJjD6yWCfMs+D3Y2smMr4bypMZXsnHiejvV8C
aZlxGIwESukICZtA7wqBmc7S+neel23f+1JqM0jYb9+W3OSd/fjOOr7NZQbdu8eZ
zV+QPUWijlbdf/XhCgDsV9uu1zEnNs3bCBCcKjUO0VxH0I14l+/oBQiBSFPUbJmd
GFznFvfhDcUksjYX0PAsYhlOn15ZisS7jhUYVzjCuIFZJjXJhvJxwK6neoRvZc9w
7/q1O53CBo8ip/b+K+uXtGE+ldP0dpi8R9NQ5ILklipxD6JdejOlOmYl6qquIXZw
PDkp8E6QaUzI4sjNHRMx48QX7LCgS9Tpsrjb/JGWbya2NnkXQZQ86hx9rQHc4+56
HbAGvqCsB7AZkskn7cCrFhPytpBFCp973pCHD+QBnDA9OlivAxX3jSzel7dxCk1s
1xMc+UG1pzobb6HMeJLnaL4YzAlFOIBID5adhtkUFRnd93K6u0gzMGhtmXEyl98G
JNummCd/ga8NePJBAuDpmx92XPcuGrs4FpPVMEj6G97vgzO0n2A+iyc/bMmKFNbP
RX6tQuXvBxn+9i47FQwXKCfhFm84VEsFH9YmPRQSnKf2ns/PdrJ/SikYygjYa1o0
iek7rv6g/fewuL3TVZ/GYDDyrjmckBDZ+rZT3q04PcyV1+7PN+mopQxKn0TF6ubf
LwMpXRLugDgqtpsDwHOpXaPV6dG8zlBLQALUlD25W4Y8m7zIL43Y3du9d/EXnDdB
n1uEcI1dp04RGuv1saQYfkfK6cPDkJG4NnPRE3cAW5gtzPnZQNFvL5r9SqSnX3C1
wfNEAGs6os+KEdh6sWMa80YzUtFRUdxk34uqrPl9enEmqnDN/pEAWtOyWJwAD8WS
4+k2QthYWLNsgP9XDkydnVFiF5NVlRZ6E6wfR6l0p8ejgdtQqXx9L1Ed2UoWbYPu
u8duHryaRxjKNP5LnIHTrwyjA/1y2pudyNhEkpYRL8RxbnkEllD6sHbMGy2AEqk4
tzMpv4D32sd+5CJ7DA5hvTl22R1afnJbSoxlV/JIsHVACv00qwNWkjYkVLjrz3y1
2OB3s/W7fAlm78IgOKU0Qeb9pf3krt14KVunYL5TkwgPa1tcnwSb8j+qQerbXAv7
q0dUrZdvIKK8A6/H9cRxVNnmnFBBloNcRgWz6xY0dTYPebe5Dh9zAq4EEcPWrgLV
69dhkVVmkecIQxhuFoHQcOnqDD+CvcFa69Fp47W8LLkVNxLXcE7PS67bw2XcOdfh
SX7w6UbAdcExj79NLxjldBbL5ajIaPXrGwm72bxGVnkRZj77W5ZQUzHYlZjD135o
gRpnlWMWws8GxV1gB1hsfDO+K4TzjpigcRDNuT+XxsVUFwzTNgDkYQKJ9sD8szQE
McBKcrKbsnW2ymErF53UStX0WsjlwzJCxK32+gGbYxO8QceBItrwjThV52rtObX2
tl4lk3YD3+FGZg1onHQ7Y97ocWIiaisBYq2YVd7NtMw1PGL+BF/7NFPI/p2+5YWc
dtZOE4yLAAjbEMv/b/FmDsveQRE83B3J25pr/zNNuWXkyK9NeU6JxmvcqJHSlyIc
ddRBO3Oea30YNlMiapqNaQuyxwIPQcJpReFsU+Chbd3mGeBGdNFTBnqcWgenpLl4
QnZ1CQF3XIX9Tzeu+KZCUmGZCU8YHZQuHt757Mk+5t2IFVJ+z14u2UR/QoKDh2/a
UGeGUUH8ZRBMIycBAsHMOcHV9NA/IxrMmai4HFno7wP8u9C7qxbvkzgUf9fcoC8Z
B9M0Vvh/EMpNF89ioUfTNVnn2sKxcP2jO3IQ+sm0qh/krYimfX51KSLCR/uvQOrV
p/PJpb4ES9sQFQeQP6RnqNDCAm9xQ2GE01qPzl7O0KP1C+F2fJPhzqUtbjDVfHtH
+B+U4NdxNIEYVCXS9BcSXEHh9ud2rMe/cLn0yjOu9xYSR/TosH+0Z29can6pL9r0
HzTWE0krriNCT/syQtOIZybLIl3a1NbfWDbf15HmbBUpYw9K70whU+wpbhiE0rMN
IMSJKSssYHB5tmIoX5Dx4cLrEvtQL/yzNP8uAyrUyPK8+L4I3SALzoxO9pGHhi8g
3voNGjDPNGeajZLCI2eZbAH+HaHQUBUu61/cpVhuBdcW4ceQ0VN/r8CqYib8Ysoy
9VnIJz0PKnUXkOOCdwThDv3M09zaQBKT0PP6sIYtQ8qtMRtfJo3NiGWfZCMknnE+
erZrh7IFnS5Fij1LsEvTMO9LiUJYdHjg2aGRFeYnZyF8VfLnZDC40P2Y+oJ125t3
tFYbxCzdgQq0/EdlXXaIfl3aEjCzasK66LsEV/SWVni9fUkfPOtjIc3eczj8YUnw
pHlyop8c+jVUYvPxtO+OF0j9466S6LGBHvDP+7z3rQv35bXv3A9X5ucCpv9iGCWs
ijn5Ur1zgMprWbooWuTwJWE/VquYobRuhLR7k1T5HN2P/skqLPbKCU5vXi9T7BwY
s3UbKPJX9y3FVjnjziSobLt2qHA3CWqlh7Kh307OutSYSSpAUzaNswfhuxJ/47mQ
2TLO1498z7WCVnD7Lp2UsztEDpprcRF4Fl2OlveJ+rVeSctgeW79JffI7tIIgk/3
msBp6oLxG3J+G/KwqQpY/IoMx73DLJ53vrapOwOFCOx5XSOgnNBG4vAhi18Xd30I
FZ88D6jUGVOjw9Fq0J3PaPrnv8uOGsV2selArKwYKlS7oyO30Zx9kxgfk3e9e0yj
m23KULq0c42NU5BRtX7OeCLy6XhDKQ87AY5lAIZquA45+oC0AcZqKWyain9U2ONF
x+X44B79E9tqg2eR/CZX3M+5peu/eQ6zs1DOPYa2sbvNwUEUmCpZwO49AuT8nmEj
qVePXEHMDB9OvmWvYhqKnlScYjsNjVdIcNT5nS089cesikMNqXypyk1XNCP0u0i5
rs+yjPdUtsSUOX7RSR9r1GcwAvsb+OGKRxCSOAHOUesjJB53n1FcrWrfg+3isNnK
PoIcvacJQn90/nR5siunuioDRQxs2KNH6NQUhOB7XNicF7lW30j3NEtnQGEwBb7d
66L7I5eb/oT0njC0InRw/4U1NZxbDvtpK0dywGzgxa6jvmqtY3WNMVYWh7KFFKXI
ZCDe8PiP0+aoT7w0T8CYi16eDwE+va4ewfCU38nQfJ4iwPnCtrJufvmcpZ1eVHbU
TB8Yi0oqQ64vMZLj8g87g029n7JJTa09P2TSoPDUwv8lLrLRKo7iWnaN9XdDC0Lk
X8p38ZbnJcqkF316bLv71qUWCxOqIqD1ZLbooPO46SctL9ojTPfASRLq43qZclHX
oHy385OJ+k0k7otktuOMtA/A4P5bgz0uFvHtfNpU/HinsvXD/4htOxSbfFs70DsB
KgJJEadBx8RRsq/HRRGi46B5d9HqZYSpnP3junPEw78PSBF3c1UuMKvynqsHge75
Tp/YfMSsA1bUNEaTwz5wFPk7A04JGhNfWA9K0n3L3/dkvhxiJi+zwBNrJl02ft+q
vS3CCXvX1Z3JwtxEV4rf0bobQ+Il1qfQcepYDgCnVk0hFJMzkMetB41Ol7BU+Kcn
XoYp7FoSJGOVQNqCo8R97S+tIM67pr+EjIxpTAaN9kp0gdgXPE3Yn/pKHB/YiSBj
jJ9tEsWI49kYzchw5gSqCd9zXbZ9x9bqrqhlhkjObpqQla7xLhSiuSY4tZ/3xFGo
iPWBr0FfpWqGCFflAP9rJshah7/wEjKql6gVEHcQ8uTe7f2SGBK2dE9qeJgC0CET
lHdnUpqA+ryxodMmMd4a+rmiz0YXwEbGtnwu3oTKtu/f4QbQjzBlM7j77U92vj2w
legrp3mBSXl+5na49SgB+2qjyyAGKfTD7tIi5GZ8971Wvupe805bk3hR1oLI2HgA
6ryjiwasu+f1vHBaeBebu+uWXCaZfG7YAioOF97/azKXZQj77zEWBF6EVoVwrvJ6
6ZRYPdXWCmF+snIid8/aj18JazS3ivObQfqqaMq2eImdnmr8WnZPXdqORjvK9MYT
axGk7yhCtaZxqA8dM/aysysk4a5USVhH2St+81RrOiApGGJHEgESdwjVzjIJeogP
j2Cb7dMcUiMrK7KuwUsymHhI5jN2Hhe7/qU4R7EzQgIcV+ow8suiS6RbYIQhXPCm
YuOixSJcsGM9CdCQ6kma0ReX1PFM3wReTPO54DvUC2KaLU74MAccup2c3J7i18Qk
Bt2+VZiOefuIlkguBnx6a/2uSvWSIsF4+fH7AEwJUNDcSpJupJ0aWEcB8mDWEMo8
XgTm2k1nmIxDR3P5/kRe5ZxgfOdpWN3pYNEYDEwsvaCXpAaQ+GlH3qbO7R4p3Gpj
rhZ+B+L65t2ToJSVGNmMOnTeddiGbt7ZIhEcTcPWFSDoujNBzEFD5DAkFL9/JWKO
sruJIhE+Bi5B6B9wwyPaAxMgwyymb3TaiNV9/ThldyM7GyNnziT3Q4La0hdbytX2
F9SLXsGF/LfjZTigBoK3BrVxDcAovm6EWgmRv7DJvWYG06wyZv94mrNWDDVzg7L2
Hz4Q57G2t0BPORfyXROZ6CzR4+jlupaFQ8SEZXP5N3qjF56CfS4VD3zSjrAPBRMM
23Y9QMDXOLbFzG6bBPTqR0GkM9FSXP+erOTodotGBa+bPBXKMRsEpS+dV/dgi5ZB
YibYKPeQaN3vjhFdja44b6bQHua0OPJz2aTOJgux0SGzhDUxwtj6GPoFPxxKvX0e
H845XZ0JGBBJOahOdsVyUWgmu/QOk28F5N4TVgxlaLm2SdOldTHUZEOPBGI8rzhK
zSMIxgDRpLhHqWFm93lWIeMWiIbH6itAUBpHENYedIYcWUIfGOBzKnwVaPFn79aR
Oy3li7GVvjQ0W+IvD4z+XEAilAanEkasTutZ2oY1/PhQXc9JdJymlviBUrhkRgVy
LEJlv3zQh4QhqmUauC7eG2aXHQE59XcQMG9KUr3hB1FjOcW/fyudhQU74850hokw
jj2UTbsqX6SI0xucG2icp1JH2ak50FOuAUQwaU13U6USdiePcyBbfzz1l1j7ivqT
me4SywiCAxPoGJeyYSiIDmUNP+PwH0LSMUtlPHmhubUr5A94Uwa5+IaOg1wgUIEP
NShhk1wloqILm/6/RoR2EAgfMPburoTmd/LjWTRHpWFxpRG9lx1uhZtWM8N4mFfg
0XzAdVnfZr/7A8qf4NQen+Q1YpGiVki6aT28QE7qkg6xOre6gwTvAgDg79qQH1st
r7Lmfwwh9SvjRJUfcIuGOSMzQHUlSpnUqwPRfXrf9zxKPEh3Oaq9i4FEt+eJAJJS
NGsi+3ovtYc1y0fJLi9U6v3sX+smiJV9tvR9TRNi8TLuPidNmOcaZ4OrmdFURhk8
MdeCrxn/8vVb/SmUpJvNR5kmwkO0mI2elhvbr7frSBTFyZRwrngavcszE/A4EIc9
k3F0sADvDXiK608Uu3GvCWNn+Od5QGLV2TWKFw4Q0BX2wzgY9YTdjfCFjco8Ex31
WbyQd0VFi88ApsGgOfFBR8ou8Stl1AcsukZhZIgz3rRTyOYX9j6+14bCWyWM9W94
VTN4Dg0nG9F0BEjgw4xySicp9rtV9nVJecHP2oFy4ysjG3oJf5MKjPCRbo19IHAg
NiB1EY1trae1o3eX7OCYVtQeEJMW267XdzSziowbNm/MPdgeGCv+rnj98tPYE8li
87ReNT4zspu13wtGQHA64nGFejivo1UWY1cYvIOdmr15yNnR6/lEEf5XYH5gRQI9
NN85prCKpKBKV+3m0Eo4OAxS6/yEQrn7+c3DhwgO6BJxtUpLCYFalcXQQ3IWZVqr
DNipZUmQ1l5o/HKvo9jPfcfO/wxtOl6LZCR6qI3ELDOIzZMYDvrH5wcNuUzh2Hi3
ehAAvK1SN+eRLcheVcTwkMMd7tka2J1cOkgX9H2WJhpKbKaAN6Fhl5zHlJlwX5/T
p98bisS+63N/pXw60ETKNhqqyu9t9waehSWamxdcXCwJmscGN2NwuVlRHFKgkq6m
XjoH+y0sCQDnq3UTmh6Xvv+7dlwKSh759RH5bxEpooJbWGig/lfSFOTl93SXHApM
XjFemyaMeb1dDM4YXE3IruGdHvUOjNCCi6k3IECQ893MJxTIBhMHYjjDQHziROe9
PO62yfpD2yj08+XJdOsdE2/Q72w65ezZXYHkOpmfxZaIdJqDAsvRik0rse2jA1RG
kLBloHsrUXH5iwiYpEMXxw8WAM+qy5EZ2I/e//+FrYEUwh7BqyWxbp7FnkAmczcl
3I0bsr2GY4aVvIfJlaOHfr0MjJqlxDAAO/LqILYfscfnbTsM4ZWNcXd3UnHzlzsy
xOmU85r6qwp6g5xkCK4LEqifVXoAoymHPY2A7cfGuHpxNTsdaZ4KFRYrwpey6zeU
h6Z6Vc6kVJbPETa3mjSCFbm7enZmB53nceqolZEJgAwHtuEJJCWWf+21izSkN2Vq
DFC9h0D/zUKLtbvb+bX6F4UmrqLUlpPU4gBKVqMX0jUoK8ya0eb5vBKwJnxsDabo
0ZoLQaoebl6T6I9mwomroT488oDSubRsvQ2YIa2YmKMuGNIsji8+MGhwxuTBsPQq
bA0DPwntmYc13mOPImwKAMyKI+Z8bpH0MF0tAE2E8fIBBrXPuhdBSMsTOjIgbwKC
XvTWHUwgVaaLlmWpvSdafObmLw5/sLIFHyWjHvId8mpLnyGa4wDYdyl2Na5T29OH
mBSpF998oCsiONOIJdM+q9dCjgGQNTwTUY90sttkjxl5uj8jHvVSKsDhqiACqqIE
17QuAyDS7SBrsI0a94vtmDhLww4BBcN1qWcT2s+jrjColyHZsGYfETuNyzTdcQyS
ZZs9V5xDH2f4T6t9L1gd1h/zqDDZnbamTnpEkvOoVG00Nf37WS2piOHy4shSUXwf
DMVE7+RBeZAbJUWCuiQNhudtyrDR6eBBRFI3GmiCQtFoFcXUPADa/FBKKICKgpWE
V109Dh19RmpC2CZlIKf10D7nuoXyf79UEPJ3amHzQQctt7FONy84Z7xS2/0zP+Yy
r4TyLKnDIRvQCtpgAKd2OSVCHnJBk2W0dXT7QdkNBTeI6WZ7XmBqhettCeBPsqtm
m0QzWvat2xQ8rrDRjggbIpHyNmlSNbAsrOOQ4Cz6fBPMHqsPIgBZXfiYBHggCfIF
ehFGZPqVT0FJmW7r4XCj+m8iZXQRcmnp/Xo8nyzczD4Lsg/F3s3i/klAoCUgk/Pc
9qAnqIIidd7dqEoq2rBKZFB0rCzV0cE998Rvt2orTHX+DRO/zpUsM0M/8B/B0gBH
HC2e9Tk3Avhiy4bI2IhEta1flsZX4luEaqapXRFeiYalsAhRBQMnhn5LqkdHYaCv
wA511TdQg3FvFbAZ+BGjfnFuCrwiUgorZXWjwIweZhMkLAcaOiMDC4THag7ymy0r
29YOCA2FE8QNYwunRdu+WF7JRryupVhgZpcZq7Ckvq+caQxgRMIkLqaKQuehDhIt
nyLQIFTCDSyQRxd3OJ1E+cvNunseprpekaYSlKdqx6mUj/nkOe+y0R6t3QXHJ0w0
SeCkdDBkWCxKkVZ9d1wvxXgSjMlfiKZ6qcq1teC9Mvy9uYj58GE2rwgLM9HQkBNe
Ol7LQ64WM1N5A7402nBno5XQo0q1rmS8TqaIOqVvFhM4oLW19Pr5TbBRXfIOcxCH
svBAxDvuCDiDbWL5vzHkKL6R0TCu45lm+HcGmovaUf4jUzK+im4e8kc2uSoaPGyF
xjO//OJbOv6j5Jh0BpqEjKq8YRhXniE1e3XMspaDZouUnqnnZec7xPTUgHIK2WYo
zs2PZG/k7qAgifnn3db4YAC1zoXXFVKUwY+4Ubii9wMMu2/k5+IkgVxJtxMDtgx1
tF4ffVt5sHD60jbJvdkfEkDzKwP7kRSTD2g+ANsIyZcMhDBQzljeMfH5VfQ7EjZG
IQlqVI1Cf4xVdnn+2obb7f6BHh7RX20oBRnI8QDdFLvY3tveVvflkl82vg/WRwcX
MtaRvc5WeVNDlZ+LeawSVqqV7QJL7P+BtIpwFP2NvbBEGJDiRriJYPbn0/L9/A3Q
V3zERxQ3WoTKVvBybEiUbQf+ogDfPNIZPfRVCUQXoEzn0iRS7tsuKjUo7FXWQmn5
l4SGls809unybRt9Q7l2CgAUdpxB1YtaQVMWozOg8lw8+28KnVbbpFLVZSjI2K0H
gUa9Hzk9lgwAPhow6f2J7x7ZJgvuYkQMdp18DFq4xiAEsjGFGWfxJC5ufwlgzj4Z
Em4T4099mzndQIrJklpYEGm+R3mZTDv7VAybkp71TmjkRuLrf3nCXToRCKKw9Q4p
BXPxpfAV7Q30QprCP8w4c/24Mfb5+VmH8/vm5onmogXbWudeLziGeXDQAl7CcgLl
yZZRx3YjWV7PpCMD/pbeQeIzlvU/riMsRe8KoDV9ABBoLBNNAsMbMDLE2CBXG4jo
tVD+TBjTW/DMXNRdlP/CMxrjUsAGVPotMOVjlntF4bjHGI7jXVHXnfEHsHOaQgWn
1ooKSi/nvsRxx4aAe7cMqGRCbQftQFOwIdk+yLiDZMw0MUZSd83oO7eFn2JfyeyC
fF7yEIZNwCPmRAIWe+glTzU8Ghh1XnXL8wI4rxOv5lJzM5utXwtTKJ3W1gjNaNGY
jyKy/i6T2RWAyVonpQanbK8U7iF7DYmCpf8xMPGltjwd0kKSrl2iisJfx5+lYxxh
K77Gpa1AbTWA2wmpVPaGcl+2dzbVYg4GSisqcNg/Z6zrjgF4Ac31e8uOdr/Gm+M2
JeiOPE8Bqh6mEh9ij+U20nmvsXnofzljec2/OG337KIvLJ5o3Ke1e6v2pxMUB47W
oMzbRKGXB7Khpl32bvHqeOeWwX3fOYybY4MYKHUQT0kIKrsD/k0B2xcyC1mdLkZM
7KXcGW3oxRVm0m1cf4CoJA5biTOFlmKIhqlWBx+Pptbw4AGxuDWEgc4uLzOgJOQ8
8smEnSePw4umBBiJYFIGbRUC1vBpaqEKqj3470DuOQCnkcwqPbvLMGYHul0BrHSC
Cn2eLsF9qOmiRLeGpwAWR4oY7Lsx+4Dsc7kzxio+Q7H1kHQi8lYaHL0Qz8lt/OTk
PB3Ctat+QOOtCBjKFh9XtL/RGagGYQP7AIc180rrWsJo73/6FvLVB5at+Io9l4RQ
ayMJ5s9+7QS2E+DT93yTzfmsOIBKPZZnY0hWBYoGtvTV9q+nOnyUsY74ae2FzuIU
reR94VIJj3GqRrPq90CnzfD0feZoEOUP432bSQGi+nMB3h/bLPoNpbsROScUitEs
vrO+iiAkuOIPBssXvldSkBhTwTtCHHyEoJfS01kAO+McuUG0cSD+b6X0N1apopb0
2me4837Bv3C5xMIGiju4lY71DnJ3GoR6fFXFlMLeV2yfZ/CQisOlGgq7BYRId4v+
mbDLrau5RFT2V1KkKrUWe0dUoPrv25xjKJjJDPuSeYQIaVtWs9NBnrrtNDtykaJv
7OMTBcy/uzTn3VSPDIfJRKQWkmuOElptP//+1jScWs9cW+h1onz6z9BsOWkw03CE
kMtKUH+vSZP3cnGLnRXoElqhpqoxSVtx1WB9hUUDM85XcQ61ZojOdrDmneweLsCO
nHzFCU3v6CIFerFvDB0bYglRXcLLJbnegXeZWgfrHcBozh753fMjLK24BYL/L/ET
VyjxL/4QvEKlH0cZa9NkryMu9trNqu0Kfx9J7fhVKvtBLDTbSfmutKncOelDG9K8
1P/VvLdWFU7P7O9XSzgd13/vSWBbWs4ynZRJuAbghzkHZAy0MxW3/9bP7rw+JsYd
khV2c4Dob7E+koJ4jIb+xxoOtVj3CgPnG7LzsEudKXOEt0KpzmOFCsukenQUzQCZ
Z21+Th//alXImT4RqU5gF5nXMBQzl41dfqneturr7w3mQ2KlzpoZk7p08L/WDINy
V5hCk9It5OhCYF4QNheFueXjVDqvJrvDy2e+R5kWTlGA3o3W70/eP3eWym2RvFHw
JVwPICCjFPef216YT7YWu9EjVHLC1TA04rHWuAhPJw+/3dKFmIrfl0gMAcpYmhEH
eQv/8ecNskv7GJyEU375BZbsm6UQxZFtvtrKUEhKi7xD8anLr5PtHdm29G0myIKx
cCYj8u89nf350c2o4xHpx70qv+HGrtLckInIYjenU2uWFRfSkYIPZv0x4KNExbPe
6kSMF0IrZKVTJunvQNYjXTbMeXpoCEHxB+qGYsZJHarDbGenX9ogoUoSRcdH84sv
GvdCSvnnG7DvDvMFLCEdC+4GJZMqpMz09q7xrt9XSpN3jPDGgUTO36a5TdQisu9F
18shyNS22T6R24g7h2/X7qwd/g672k0eASd/XTDiEJ9tAbFV7NAPiFJseTJgWGFh
RBmg1ks9mq1q9lhVftFdynF7t8OoFQKQruWcIsUt636znCU73XKSFTkyBVAmOpac
dM+Zf7q5o4g6KP+xWMZSXfWyWs1NgCwiZKUBR+sZ3rjFOkFnUIUQU97Q10fpLkEB
h2PBDpJh7tBek9Vsw7kP7eUOniw96/0vCksGX2OQ0EJ4+4I2nE+dn3y6emQoE4Gg
FdJS6lCCq6mDZ0XfQudJ6r56bDa3akqlhF7OoKd1EjjkEn+j13QZ3FvCm+czaBjG
vxzlDWcA++jSQksyW4+13drvDx6lRevDyKJIdJBzoGVSI/sqBKJTkTxxzd4dDFtG
VusFsdWaeLvz0sFuJQ3I3RpJePJUDs66Foab8FOAnswWn66MHaZKmlSIaWSOGTHU
Bc1zUQvVW+eLpGlVj41k8Arq2Uae+UPoOA1qEJ8lr7iavDTwL5zpsn6WvtPg4xZJ
2WZGTXGMuQbLcrcNDej/3ozNiUDf3LZujaGHikhJPefva02UpMfBR7qenxM9uwp9
v2+OT0DH66Voeaiz+e2ywGTT2uxhl6tKBbSOlolr9A2ApE0CD5xzUwuvhTz/wnvL
Gw/tX6c02Wo9UJnq/oG6lmiLNT399/kI6/mpqnQgepctaXa/S+zeKKAzWWSgXyg9
F4gLNaB2Dh6K3IwQzLpzt6wKP5N3CxEaRO9JwCKxSurEjhy7sQZcN081Dc6FhZAp
/PGlSL6ciEje9LiQ+GZzFkGQFTZY/fac39FoGbuRvKyER0x6fXBv16Za1mw+BCKd
+5AnFU9xusFuCWQSum6f9LgLSX4WpHUeYGOk7kcAeWMXUuJRFbUvA9AAHmz6rS4/
s6VLcepraWOrnduomEHilZ8JLtEp5kb5jdChvnj7WWEBTd5QB/rGQCnMbNLmqHAL
80xsrDwwCskPc4XK2qYkMJzrNXSRxTD2nc25E4/cDpUmeuI9WccE6izDeY5gMIX+
U/1G1LkibeM/iRKhr37jQzlyQEX/2cySncuMxv05k7lxb6do8rhDyRWCJps1Hd8N
x1/cWz1KF2Q5fuROWYULUjJilHOojM6XbqM+NBrQw26/cDYOG+sR6WXDwS3xiFjt
loOZyDQcLND6IPwnWQYtF5yzJZB2lA7GxFH2ibpWPZB0lC3uc0BY+reZKeBbR5uk
3xCLzBpZAXWJHMe53XdmaswmnJbnc/y0WL0YfU8w3URAy4hgIneYWP8qpUgdolb4
frWhIGk6e/RGrLsb9mj15z+v++AET1wXE1FA5mKWuj/nwaHNqk/0vQglZdpe5JjD
RgTFPDHT0rquB4guJabWY92MPM7XPafG0/i39oPmAf4Yrsh/0K3KH8FGlY9ziUhi
llpv8wuySG3KzkyxnL9wdQoLnjkne2dAbMtWo8zVmr+9VF4qSpIqkIx4srRicFwW
Njrwcsi3UBpTXCYWpuwSYt8JYBy8okcXhxmfalqGrXx9zBp6DaraGSo0O2cxwUWt
qgyPzWqrID36+OtFRsl0Gud1ttO9u9tOL43hyxL33Sv1m7GMUCdupn25cLufqegN
VzkejJH7Cf5eksUKOPEfCzNZciN2GAVRyHsoybvcNILicok1VcEsa7rzrfzo/g7C
wfy3dvoUgPS0Mnf1FDnv3l+z6QKJebm81ZUI3aMtRti73vlvAx0A9y/jt8+65FY9
Ctvov2xaw139EC22F6GJeVsG/btBOnflaA1QnVHewWkjc/IPIMDCEgWfxCPeUyG7
W9GGuyrL5V3kxNip09fGVTBGDmWtGD4yXlLkiqXw/TExPGoqZwVZocTJI/dzKtdX
avQ5BkP1xLmEzWLEpESZM3OS+gDdlXzs6EutnS9dnkiY70nIuuDYnLgZaSnXW7QW
jxR+Wc5m4fSj9Zr/cFh4pyTthmGdFtHyDN1pmY5r/vWqSYBhhCsck7RdLW6TgOSU
opTSmVi1Qm6uv9O/e/WnrKW/ZsZ/XuHvbeHPWOaEdhOXp9U9tro0scToNVh056Q8
C3XsDpGkHMhdyt0+wpdWywBErea3BpqqqZrS30v5AAH8ZBM4GJKL1XvgOoMzo4gK
o9rSGqxZESCtjOMfP6q3Jawn6bqCOWrW7oTGyI7uo7gsXhgrSTn9Vq9ykMrg8uRT
nLPgzTTjYTBHEG6610ALH2C2nbu1Tgpnh6MBQoT9eS7jWVZpPZ3e6piHA5/z2SdJ
Y1sYH9s7wB4JjHE4LiwkXyKFnxQ0HFcSId5WSJKCL0GgujuILECK+ueHlIW91sZ0
OqP8jjcqC3ykFKYdRX5bkQkSOcqlvI+4vuBtynTW3PhXhftNt2kMtG/Jh/cCxsAQ
34uV8UBh/IosFWjhL9r/9Ur/b5+H8JuXt6oM0wuCVthdmxlh7abtZA6sZKsVtHKP
+1Zk+4SzTXKeOtwWk7mbXaerwaZU53sOPb49gHFmPCTB1nhqgNPf95al/QADzYs5
DIrh4DxtdRJNqbJ0MihAOqjnSv72ZZE1OzmVSKzAtNgLf8kfGOaJh2QJEsbOX5+J
YNa0f+6ltx2pmW3gAlJ5iKPKNHAfCZV897zq/ANSI3kr0/cSfGW9ufHQO6q/EueQ
btD4gD7p/tSPYmVeTCbpqB0c0+9fMdhwMkXMcCwV2NkpsvjKHmh1ShpaX+ZMe7Z9
R1ATMoyxejqP/r9MJS5o/rU8O7JmlXKEatWcWtos3AchEKA6uFLIeVccQa7v/Gey
mMcCgw4JA+3sJ70HZ+0nMz3gs968Hwc7JsnLQXHWfOz7jR6kY3YprQNfI9SKLCey
GpLbHIOP5dV5uhYJlBqnKZ1zjjQhGjq7RemElUYMf3O/uBjowd6xuqrVZsEHswnN
7OH2wdhlL2gQ/2gtfPCkpdah9NhXejDbcUVu3cttLI22tjoeuMBupPyejMsOcgpp
wncJBkw3uvg/pd0m0N4Dvv72IqfTCEoKqHOEALEjShvtmkwfs7wk8vUDDfaspHgI
kGk5a58aq/XSnXHd1Ci1lllYD8pbsM9OG6dOKDUpj3Zn0Ha3jcxZdnpxpVVYfhwH
jALJYZtPxKSUQGJPteqFHUuPia4NTA6Aj1sUhH0ssYZp8r2m9tJkBYZOWCJx5XZQ
LQ7wUYGJM1/ryICetFb8zr0YkCfLHuGWnKqaexA6gOZfScSAx8SxcTTrLy0eBCPx
+P2Z+IYL3j4HfFV8Ll9nI6rMRd+Nyaqtzy9pG4sqsCM1gZSDix4zGEuMql+XE697
P1copMoT/y8N2/LPMKp9JNwEtx1AS60F61Lgw3gN1/Xbfkh6+gRJ8WHHxIHhXGIc
IivN6D3xXPmQSRcqp2lOBkdFXEB27il0jYj9KJz8QoNIQY7T9qVFL9h8rgWaL0Rz
pocbMSnyylYke3ErHQFagGRVkGwDNEi8yJxoXwxI2rBwL0b7uoBhDfJ5uJrcRO0p
wv/JRHouZhNjlFgEQryXsmg3rgQSH6L2zVQKNjuqbXHzellzaJWrPyxD4JpdgO6j
UAj2DNtV56czghIUBGNjprZ+QxylFhyYmjuCS7sVIw6OvA0yvoV+UJaoE8lc1/dd
vSFTx9sjPc/ZM+arpiKHPunKd/5pHB2UF3QaRdonggCG1H42bMkKDDGQgm8r2W8h
sl/G3yK3uHoTVhkFWdLK1y/Z/2XZGC2fN+uUPlMj7pp66rUn5NzOu0dSy3ODthiP
cG89HWTdy18X3bNi1k4IF3pm8y+RD1hU91jnhF5uezrh5/VvmszrozGUYk90o88Z
90vW7m1+83dxXDLic0T0qZ7b868JyGDoSZiGnHARtOtZoxlwVRcvMLbs8aTkg8/j
`protect END_PROTECTED
