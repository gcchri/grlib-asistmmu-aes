`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j7Jj1MixarvornuV9XcaARNLrOqu4fvZLcY+Uu7kfLP4Q/6dcEgz4fgjsGczmCQp
vJQqDEPEP2G7W03iOEJTjC2flbOOJArlUqTUgjoQ8zJ4sNFNahzMBJmuQQFqpIHU
As5yW2rLNsGc1vszyNapGD8C94MFgotC7wJN8cyPcrrIaqOZ+Hr7juvJYyNymtO2
hH7dGoMdlHeznJRGZC/WQ8tBYvk/PQjfR9e7JZ6xgtPEPr2cnXO/DyCe8OQ4NDGb
4O5a1diwB7lK/Fzc+H8WMPXpswNxx9+V1il1cMD/+C/+9DaZtS3lwZl1jC5ywffZ
J6/iUodOB5yQvCmKzgGw7P3emgrhqM6d3aGtPiJVdDWZ4ut/6uUkPCH14OtGS+sq
9YBU5YuAGT1FXvGH8vZoFDpfzSaSZpSfOaRvW0whviGfB0kxTqtB4VKEimTWpge3
xpRmOI9kZ1NNkhHINb4mCfteSQTSyBieyQLm7BGXZZt1KWALFpysAWJqpI5VqWtR
Vs5cHWZ/3GEWUcHvk901O8OBbt7+H6t//83fDyKorzG8vik0m/g2LVoRl0WBD6fB
AJi+xUDVjy+mtfp2vis0YjCLBICVzZbkI9J7osLjBGApchDL2fBp3fj/XWeyUZO4
Z7IBc2EKUL0emmkwBNb5XXPHyI0eJ5yHEtOzaA84PdzBlG78L4MREK4ECutokUbd
efIa7sqoACEteUsVQOkYhxsB9qBQJY6yXIiIOk2DvneaNWsGH2GzLMuUpgqiP7uV
`protect END_PROTECTED
