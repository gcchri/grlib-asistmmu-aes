`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7feA4XcY5urANKfDW4PHeWSUqjXgZh+uqffkBTsTgym8TYil15eA0p5YePCs5l9t
gjI3j3OIkh8YJe0dtUW9LKQaamJ8DsyPWRcz6oAuwsjNq2uV8GhsG6DX4WvGAYkI
GBbz3Edr3aWIzdnnuNm9yzzrVef3TgWUZvc2vTfVMDFC8S1GlvGKRVMmFHOWVB5g
sO7uw/0ZhlYq9RtBcODoUw8CyH0YlFv7LIjREmIKiOy37P2wDouwWhvyqC02YyY7
`protect END_PROTECTED
