`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FUCXd47JrL9Z6ay82lrFGIbp/Jrhugit+xeevrgXTAUsYaAM/GiE2infH3DxxHdZ
Us2k8oLS9HXpj/7h9UViXlN2k1h82rfaIu854MjTPIPmGCvlqYEIwB5XxPvZMUMm
mh+2Oogbb/zQTK/uLA+qSsqFqdrAYOWtc5jCCge+1JqvExEaCOBf6y12MoO+Aygr
KJbDIrM2o7yUMSwuRYXnVE8mTYgh+h4MGF64Bz79QM8v9RNWT8lGey3cwhU2LptS
SL2zOnBF8/1EHXKnhVv28TtCF/HF5gG/b81pq9dKJerXkLBLDxT3S+dDI0cYe+Y/
9ZbPH3F2eTblk0YmelzR68ZodS7wsP96UthfUkYxHw5CrRUxU6Fz914Np5K1PKEC
BDjuC3xR0m4gnEUC1zr0E2/bo37ijnUayOrmA+wHvm8HKfAjHAjjhrTqxai95xt1
RX/ZbIb0DzRGFK1pb1STe+G5oX3xkVTDNsdhDOcnQFoE/Y+lxX3WCoZM0Gs4XRhu
`protect END_PROTECTED
