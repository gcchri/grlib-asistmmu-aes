`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5A5hW+tu6pgAhZpMMrg2OUkGwIhcG3QB6i457fJodCfLT8FogLIf9RR4M97esJN
bt3RvGahQhdH2ZsZWKvoanKrK5YX9GywnydM0NFyqkpS1YfwXefEXt+tmXt78h0t
2YddmNjTZU5zM3BJGN2h8NVINwrKyv9w48svDBQ5D+rrm323proTsAIvUyexewbA
WRDyVfwg6PvvcS4H/U8dp1Om0KWQX5Un9UXWbq49GFyaumzxYg5MsjvChs7jw48g
Vd4wl9unJURzk9Fl0g682FnMCEVQRLMoaEWWEvwpMzuKmfloMMRHOIHC9YMIBGfL
T5LmJetgGST5yS3i7UqQ0w==
`protect END_PROTECTED
