`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4g5sHQQwEE01fIIQhmfisorzXJtu07GSSXS5QuLaS+2fa4whGymJuMsTeTVShS1M
AVMsxkspfjNqFZIRmuJlY3WudDziGf8K9tLTiSvt58KFjwoFqjgsoo5d04BldBEc
Z5RKgZXvNIuf1f82gF6W3RVkYOtI0xCc8TQ/GlE3DFydpqGRFeZv8jTDXXEauNz9
CsylapVjQ75igU/5ZSjPzQp5hpgNeZD8JGad8HsGEcoBIpDYJtiN/Wjg8bRhhZ+U
27sYH0K4TtHmr3fJmx/j0+gXpwXfI5BvQvP/ggkaxlC8IGGjLhv86Mik+mWd2/Y0
2d3ZYvS9+bghbvdnHzBEUe9fEL4PEZvlAG6FZGBkWJyPY4Sv5+y8SXnyIqprOe5h
pFTfjxZ11OR28Zitss9NYlel1cT6Al3OdNLVxE+UkVkRI0Qt6OOSgjFzbgu2fEAn
Mot+5cliAlz7nZF28lIX7Ky/OMzG/sLss6i0fjzt1qooec3ubjZKHTJxr9stgLmZ
k18HAwxmeEEBLQ8dx65lIKjzRXEbzGLFB7kVfZM7C320pTv0ndwoY+BNeBCUzpOI
OF+pq5SV6kH60fWLB/jIIb5eSDJv4NE7164xUw/uoIGmuQ/lJj2Zpsdr7X4vCslT
JRu6bNBtRkZJlzn+4CLSmxcVH5DDaWKvqXxLta56ThU=
`protect END_PROTECTED
