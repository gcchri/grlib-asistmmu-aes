`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lA2K6gGlRGClXqoyg6uzTv0cJNfRa+81FNhQGpXfY/E/EfCY+9GzEPVx+touopot
oGa611HfHEEMkn8HeioIvrOFn1hutk33R3hLRwaIRW0i7KT8nd6AIvOgIIj183jI
gRzOFinAVRM+dE4Y04rRDXwBK48/PUWx9oBkH4EmJwkaPIXvkIH7FvuMaAw4S+AU
0lOSHKFKfX6ZbPYhy5DVxpkkB2P0eUQVE6jmzZJnI1dlq6EJr8k1Bn048ZIOI33E
9jhCvRvYQDYKToARxCznS0bgoaIPhIZfGCLGSn5Doj3OAmfwXpacqFYYqFvKnmQV
tc34r3gFp+qmNDfGWv2sa2m9ILGAkOmm2dLMYPHLBzQIgY/c/OVBKmw75XgVL2Fl
YoKrn7Ov1txoPxsHo/313bzt0PaTfk2VnjxXTTznwBCIuux/EdeYfOlAldEjUhb0
VgAfF8f9rRs0nOcKotmUvwlbzR6Wlel/PuXs2vV/+UE=
`protect END_PROTECTED
