`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCWyGsjTlxBO/OuzGtw8RNUo6S8wAxvJ0/UQvytxo9kk9moAbnEOKHN4k3p1dhTc
TVn6CWG5knWuOjvoyGuTNLP+B94Iylw9yQahU4is18Xybll7zubQWoufdirawOvs
Mq+8/QVqJ+eYPobX6OcZ0Pqp3XPL60Vo9qqW2/fkgoKT/XI96V9IalH+Meoq3QRo
mdCPC/ulG0xiYDEcgDiGzWhE74+F/8KePFzUCyYE9ps/tNkjOvQgRIpM0Z+gTpBq
ciGDoKGWKeZPltVOCf+8vBAgMpk0PXqOuzHZ72k/OYvfbKnAu3QS40kDOPvo0Gow
eneIVqEVggHYYUAoFUoQm+dIRMeDVtZAUKrd2AtKHCqk+hr53b3ghAlVlf8rCV5V
LHcIMKNW7G2a02fGwYzbQH01nEbMfXnwHsg9Kos8jZvIBjgX2qRKY14ujVvrpSVP
XEZSgW+lf4vzHelFtm2t3dQTmjtpOTSoIPRJj1sAFxatKGFNJVQikxK/d0JMgIKV
`protect END_PROTECTED
