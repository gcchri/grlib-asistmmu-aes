`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XI5mfenO0y5WXdSy2J/FPyeDzJki+ig/V2wqTeDbMh89BLUgYVyiChowkS/irtrM
5afolnSK+5uZw2Zv8rH1BSbhxFXYIFBFm1F/nR1q5dN7x7k8kp/ayS94VC9PbUM6
fmGpbLV3laSyOzsGWjnb0oPAyL0G6hHK4T5dAa5rbxsb7VIWkrrKTVnzR56h9GcE
kgtzro6Ars79+U4R+lG5nIfCPGGkz6mv8OnkCEtAvy1bYYv5Tn67L9GHS5xctS8K
rm47jGxOTfNwM6WB/AG0PNNRZsashIMxSIgR412fkGkRROfg3VeohLW3o1yo/yVF
pyEJsLV+lsO+UmhkT4pdP2YakRQo+OQmJP2K4cQPqPXjzZfVfuhPAd1JXnlCwOTZ
Dsgw9orQpOluzr3ZpvHSgs5FWr2bPUM0HBKJuW8AYH6YJhklxO5Ou5AXMkzDrcf4
Ts8mmGUbSr6xX15ni5czWiIKEP0Hc6PXqHYUiNWcyJxLJgWqE3zEI4n7yYtnQDHK
Z5Y0nPBvdlDniYM5YG041cFo91ehcO++FqVgVRexz5VXPzvmWADzBQ915ibwZ6n9
W6ie7iEzWp1GAuyIWSSg4/lLxt43FyseyRpNEJqs4No=
`protect END_PROTECTED
