`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vynozya+s25gkGZVkIwabTczLNFblXVvgumDkqTa/nEKuzhEsg1kG2x5HgfZ42oV
j1hu/HXhpWDYv5BlQnjPWlq1CBisLfH7UIqGCI7Q5FYPLFKAa9xkpRKOaNyjho7I
NkxX09D7vCUDztDqtK2NPeSSAGOYemRG6gPWCrhC9/8BCME7RAPrF5GL8vRzziz9
5wKxN/lSFbMr7d/24CTBrx+F8KYOZfNiYb9OyMXTRfw1djIXSMEL7jcSxzUZ3IgT
mlNGrk6BnXqcbiIeRicSc6ehDWXC48UirIxzjRE/d0h1SmyjmdAFB1WRamspv5YD
HnWdGWqF4HIxp5RgFl+XhZZAdeougSp8Zz+gXU+JFzLeksbU09jSy8lLpo0gRDrd
1Ndnp30fc/TxP963+Taq42Hk2fgFlmkhKrk0NJ7VsVDGockXmo23jnBpr2sh8iLV
KXSBoZGC3BDNqmF29QW+iB7qekUR0NQ4vjXCH4x9WX8Jva3YajqvtVxRttOmRHCD
`protect END_PROTECTED
