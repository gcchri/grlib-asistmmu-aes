`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8IxK105bnkOpctkI02OXgghCxDixMcvEZoYvveqZU1pOypVBkeCfn+Pz7/sKpje
RgrPSLXJkq0T/d2Wg7EGrK+3stOh5pyDDhMb9doIMhbD+O1/SZXKfOpch25ARAho
Wwtqofm1Bw4J1zyo86Hc+OxPKVIboEe+049NO7cN105VmJ0+AeIf4pP0eXaqBWFo
tqbcv4oOut8pJPxMDT6X3gQ5bq7hPI9isH6ezA9U7Mx2FYUbbObMurSDxsGx4zmI
xTiHN4knVL4RnrBb+YoEg0aKzdcHOeC4RtxMjpWoEI3l9iLiVcG0mPDWEyAd82be
mdeqYM+UXjuZ3w0zBh7mG0Rv8Cidxfg/IliOHi5qTsg=
`protect END_PROTECTED
