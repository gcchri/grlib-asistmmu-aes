`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IjSXv/xvoniESikMCCyf5vHE7ioC2ghgZxOdAxob7O7FsfiXGwVFdlMlo1/VroDE
k+kDRaRrwGYYOucXRCen6RPfY5U8WgmUJNLJce9Iwbf335YIP0tICFoTPUEsx/iE
KDNbjoG6YZxPunIQs0eeUGIoorh3W2MCM8DZn70QUTkPdlY3AXvCOxQm+vuyg7Ck
b8q+lbX7sIWILgWyD9e/qzgbaRz+ApptC1V1YCHQKJfApHPzgvecT6hCwqUQQCXq
/WyUCcBtWpNchjrYIblJMa/0/6jf/AbXPK/ziou+STW6Tt5CyJ0H2DCL3WJQzof6
0+MVgC1g/4NVcMaqn1tIrphn1goIdY5/rJtHvEUIbpxo2Vckg1HH+NuJVFfWmG0v
Z42JKtwFO/iefZs7XPCrlEbF1j/yhIjy2cfP+mb0TSA4VROcAl+ElbUcwty+Jg40
H6B3c+8Tco+H1Uww/C5HKw==
`protect END_PROTECTED
