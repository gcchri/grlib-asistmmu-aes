`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qw5BzqgzFQPrMtOvzYRj/rn5zyOBIjaTXuykNawlnT9e/gFVEMan/6BRw4qP52om
GgSn9TRAq7Jq2buRic1yW6YpJDTq+uJlqvkdvA9VcnXVqgmwh75+GrmHuLc2d0YZ
Gj/H5FMy3v1JTlkOp+f/5f712cn6/PTaW2REYlBuW/NMDBW3a6JU61MNS8O7EfcP
OBBZNHVELnQKEY1bjZQJ2gyaHV8rzHgdiKVBU0DdXHXavFzRtfqNyyq3tGqOSXGD
qtZTNOHmXDM5M3vFRNY+eCkuSGU6hS/ygdJ+o3sKBX2yueBQmdzCFi5PSeaYsffX
//vNLk8pVTyu5gvphhdV+moqxGTSBZ72OiOet4+stOt/xYz9fHTuK9jqKzuNmB0h
yXxfG4oFHBO5gyiktoFvA7blTMlOYE2s60qx+ujQZxDrsvWfkVMsb1wxvHYcFSP1
RpdwOgFj2vP62JQ7yVxEhHvLBagZ3hIbUt/+zn3cx0aUnAcF+vMI1lkEvIt5Z16H
Yy1Aq36O8uO9Kle9Pnk0XUN/hNpEmYSeafbHyKVYg4M=
`protect END_PROTECTED
