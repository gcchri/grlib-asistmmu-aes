`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7DtVMvISXnNr0QIC8GN4bP7uJb0orb/jVYJbRa09y0zFIpVY6RlpvEdfThiOPSLZ
keqMoX2Mgp1aUqcGltv/0gxHWlf7PkiasVAmTu7H20EAToPnnOG4zDu8U0u45W8X
hJjJZEzcYycp7P78PQaG/zUDEFUuFVAitdBzqQzX692Lv8Cp5qiK6+Xpstsq0lKW
ZeQ8fo8cq1SgECFhIdD4jXSrooUHZDRnKcTTl56nMXZ6QCXcnPNUzeBgiixVcJM5
3aMJX+wSCJtjirXy15S9Boe/L6juH2Org+OyxKGtsiC/krGhouHRbILED9IaTr95
gDH1zbzGwOXtxIPA97cerdab4B8GLT5u0isyrfHaI5wK3GwY+Pw2cZ6/EpANKQ53
KFA+Lv/gc2L2eTU6c5Y1pPc5fZrwc5dd8oJ/bCOiYF7XLYMeREimE/cuszJZPsr4
jqXQGSg6KTL9igOn2uPtamhmDrPWTYWD+cmBHeGRmLeKPYdFGCR+Rd+GsM+PgVVJ
mG4m3FJwflJj/UG779M4gV8qyCH7M2rWVvwjERm7R9ZG1NMiE5Bgr8ZRa1fZTA8a
TCyTbZ82qbRV92tbragXv8IrKeklvsJZ2nz2LGJkYchi6+bok9u54l4oj6OVUi4Y
lnul6/uPTZliChnQCjjnfw5yUUz4Gq5PwnjRfGTo+e73CBjx0LIgXnZsLgW5f8jK
84anzpglnORFWUYBcuO4jGI2xAUo4nOPt5gTunJhgdji3R3L4MJwiwO8t66xvXhH
PFf6MGVEXbRfUQ35+j55jP49hd2A5B1bMJAyb7hi6a2NMw3EcH1mHeAVA+zYd8D4
msxTicJI1vDvTATG1wo5bUcLpXGKnJ4lW47CzMUhidc+FfwaPKPQnuNF7MDycOl6
l0kpp5wVvCK6l30ntdo/Ok9ivucNpHsjBOm0BO0RljA7ILKtBlufIl/yuz3kE9lB
Tio/NdcR5EE8xaT3J68S7a/qyGiBIs7hqXfFydM6mIaxq/h7fkVJYF5oPyX0WxNX
vSthELUYcMBoPJecqzU0HZAK+xSE3J1EPvBDVyp5tffAEt8QaX1aMFioVTWWOZqz
CqwZzYi8ytQqR6KICvqXpcKwPuIRvGq1o0tX4I3HYL4PvjfMY0Q3jfLdrMmVPMVS
KM5gbya8R2tTDMuDcVKYj9y6mhkzVEMFlWxN/0gtMImG7PKncwmogU3DVIm17xdg
BzRT/PF7j3ZkGerogVyJkf8c4uQH6jMdVZtN6+oGhpnFUEiTTP0zTjq7Rl3jCR+m
UX6F2tmvKsQtwMAlqBd1lT0rwhiZEa+5S/3nPrJO/b6CiENFiHgI8smLuMFyXf38
OTh83tpm+QsT1WULaiOGfVBtfvwW9AKaDqr9Kf2lflutTf8n0IOoLAJk8CQOIGON
Q28zUzScpsovZBYSTi8H3SADWqOmdTohmYH/Q+5BYF5Wvt/BzQl7jtfEIrLCMMtN
1oMD1QMxaSteKo13hOc+3hH4hAhOrWZHnOO4Ysnr861vxhpvZMZvQjFm/ZJVrzSK
4zCK3OVq8Z1d1z0daPAAkIR14Y029JjozFJLMf9Z7tesR/+A5m4deyIyHlAg3FKE
z6W/cBbuL2ybQqbTu+IweAQ4Vmep0vt66LBw2uwjUw0rOdOvTA+YPDttsFc5PuXc
EQq1LerTw1szC9bw2gjpytOQbTqcKNN3gW98JA2zbK3/wT52jLH49v0AbTNlXPV6
HT5WRjR0gcQDfHKA5VTh2U4LZ7T+s2kmwNKAag3vLGWilhaZZKX1eRFyqNVjG8uN
mNX+inzTVLYGplk1nWiSLLMaJl96EmMHBiRkF/N3s8AXQ+hdbDgtK1/WwKr5VDmH
bvJS9oWsVdJJpJGx25tBzGjL+pEE2COUNe3jNhHQJPTIWgnA41HI6K34HjATlaSq
3uvUR0UiImjBKNaFlRCO2NKGWJ1c3qbSJ11cyfpfWhvND6wiYQWQuNZ2AHHqtDlq
uqxzxn6gV0UPLg2+Gi3QpogygtOhRqTjLiDALobpWW6E4k42mJH2MwoZ7EfoJQqi
VyZFG9oNng3YDSuIjKJAKIrxW97LvaLOYTvI9uJLZGL3VSnSGtjl2C1BnTNa0Muz
+GsaI6jhpTisQrygeMiAMMD1SiSRcM6JCkY0jHe3Dba+teBF8zPU8zp+IDppWxlr
GeqawBdqbzre3YxLPT46Rf2CbKZm1EU9sI8FVQVIUu00dojUz58+WxvGUOOSxYUk
t8ku78CniWZ0vQjeKOzNvB+yzipcZcSk3b8SxUPj89nDpvWVReS3ut/o6WIPDchy
PdNx4tKBAS8QrDppjW0rYqeI3sRS7qE/PF0Xfp3cVqrg/zhpiSi8ec7RJS2s/Gzr
NDqK8dE7qPD93/8mMCWyeUxqN+lUlrHG6OZIPL/woqJ36yda4gW0TaS/gyu9A++9
k4mCl64OUuUjDaeGdbCvcKmZmPvYjn63Ak4K1y33dGr+fs3aTd31T/FNufZivtKu
K6Gd+AmLOsDVkp4wi1CExpBTpy5/aFYm77jwXQdEanGB1mv7s/j1tAKKlNccNxGq
NhzzyvSyHsdVqXfu7QRiEaNINmkhMfDeb53a+SjJF3TuM4MUlAUe1WWC6WIk1yRe
kG7c1CDJkKLEYXIuE4SXPS9ISbqUMlqy+yU90E6GZvgmNSxIsvrzrKcoV92TlV1Q
5HJt4sc6KrS65C2hj/QNw5pqRVq+sWwCqp9DoZj2UQ5Xrlsq+YDXZZZHVGUxZt25
R0pxmHT85YufMx9wLUo7DWt7Gz7eFAPqDNF7miCyzk+dr5nijc7poz9IGMFi9fg/
i/pu7PylDn0L9UsW+MSmKvQFXv5zJAOmwFpJ5hFDUWZsY19t7Z45f5wdNNtdDODs
LZJuSN8irq2SFDcqk9z7qZiVduwjgpy/NSVlShTRDyKP/32vgyh01LTf25CBt1eM
1FO4jSguDU7SjjD8dafG4mE4cyGlxuMrTN2MdWu8psUMhNP9Pw7BsGg+/ziV+3FR
2Mi6iufiziN+8mbyTRL6kPUMhbpEfhfAET4q8apwpFGv2kjI1w0B3egODQE4vTua
ZpKfAo6G/6H/SvfX5bKy1pkWlpKodcOGbYmH10Yn2pJptSrnC7p8VZQI4Szm0q9t
pDvOEiBvWYWpypneCi62CwGfSfN/0XqOziu2lZDegbYDbZEZ3pn1y/DukjRO3j13
0E07qE6moojMmXcDjk9zRt9DK85h/bRmpdkdmAMs49dkg8ncQh7JWBOrcpWokHbI
bgiYAi963vlhD5Wh2XmqTEreNargLyOz4+XgE5hngCum3Hz++8xU3vjm37DEjrSs
haU/pkgSFEC/UL9+3/fRhibnZPENdzkP59IyRUZjpyI3ApuOcGBgUDxYsKGWxfz2
l7A6z/h5ZgdQ0uZQe8J3uKpuufVEsS83x/gFwOwwmXChF8Pe6/F8bpK4bEKD/uv1
EZAxx/NG/MymI/k1Z5dKbRle+bp64GL4rj4q/0c0KIuPY2PXSHjokYCkEejY6fNn
E5NfQOYS4AGr75ESbhYLhp4lNlUi4HpTiVHCKzkoy8IsWoCXOnI/Bdk0Tc6plboG
IOHB5qgiQ7T5lhRLnaWUbXPCYoudJcsnhVpCgqfyVCftw9rqGuvinxPl5VaaIcDn
soAmsSODPmzrwgIh87gjzdgOZX/dQKmhPEI09l8ebcHFbwMkwPaycrVPt6bx2ovT
A0m6limUe+tHEbXxkK2YUnQ6MTyQgRl4GrqYzZINvTl8qdEQ3hBUNc/nN+KGpv2v
tMPeP2KnQGNpM8wS3Xec9Hl2qUmN4y2mltjQJSZpQylg4jXUQgUqiulqPOul/h0q
aSDCtM++82GRJrVwBi8WDslqePyY8e7e7NchSGwLHTtuPNXdxSeGUiffIosdEti8
rAOZQ7nEgWx8AnpqamhcEmaLs8fwOCvxKAdlve8u/BdTxpVGBUq5m4ziY0YuxaYW
ebjp0r/4Gl8MOy/OMhFJ7Znohlb8uOcDVnef2FZ2xznMDh1m0Z80Gq9ZXVTeVYTD
bHQigOjptrAA9T+McrgCZuO9zX9UKv7fBfWBkg6oJmBbW4H/o1y//sPT6od6W+ng
q2QOF3tFHWgabQpBlELtnXxcGMbKqJJUhkJmVoKOqjFDgEz/ZYLam+CK2iuCvC6M
7J2YV7Tj23XDO0pNQ+Brvg8tHxY9A9ukLr8g3OBQpYe8iZF7DaNCywzSxgV5nGhu
T8eUCNocKoTPbRp+kReCIIAlZUTGGKbs/l73jfFP4v3nt5CECC+a2nWld3bejrXU
HxuP+0skwO82Y11RA3illbOjCzY++lzUMPRXhAwfQavQ4TtgA3jEX0+XxoF2GN/H
LFNoU6C/Z3JT+oMgy48yrdSwDCG9VNSNFOcONshtyN4lCVklfI77EFIUouZJUi7C
zPJftgkkvKclqGy3VTKO2Q==
`protect END_PROTECTED
