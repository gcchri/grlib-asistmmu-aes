`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MWXAZi4EryqGC4i0Gt0JN5f/Im8ldkWbUQ66Y5wnYetuVss+zem8lr2QnYbSQN3v
9ljzrqF8NWW/SIsAvSwXa+lAchDTN0HzHxcldVuC61sDZ0AjtrBag4vD3YAZLuNe
TbozK69bZNJVHTfbOUnPVanlFf557zAFYIVqVCROEmtXE81krHLYOXw2Oxgd0YTR
6ngFrrBT+JYfJnG8dtAVV/LkVlEk7Qt1JqreingogV3jMixU3salC3HvDnqLb+Ij
YJT9ilKzlk9lCRUHgKAWenyUsHezkv4skOAyFoKsD6F+bR10QId8ZBx6j3SyyQ6z
rfXuT7npAgxTexUX2cm3Sr9TKGmz55/XVoKlKk53W84=
`protect END_PROTECTED
