`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R61c0lQCoVCzGnQpnLWTO5Kq66r8Z883PwQrCgrjd0Gx4Sxdx0ncHt46a/erTH94
f/Q+8oqUeO1RU3UUYyDU0ejdvUUNBP73d5BHawMf+IAgc0wyKO6pQ34D0ahi3Fos
ExnxzCpSUIdSIPxlr1FqskGNh3WcA/lZ73np8lfcCLuQXWvYEybwYrOQooOmTmXY
n6W4Kh5ySSnWQI4cECW5GFI6EXKjSpUOaKoFTOdCu1XVD3GdApGXWup4b8mQI2Lz
S/MIGc2V//vSpvi+Fr+oUbfnBdUD1PnDmxmjJnUm+Q6SBeMVFLJbcpvWFb+H4a4V
8KUzZy/mm3UF7/v8d5ciGR0h0Cp2ViPqFixPoXMo24XfKjHCp1qABCfua44hFQez
6OCskL9HJtpAlmg2sWSycCeUC4HS6vgbMJk2rxx0nD11bkHTM5jxzd+Jav7PpccB
5J6LVdmVjMkb4u2ETmw+WET69ywPcPCvMCvxwLi8h54=
`protect END_PROTECTED
