`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f89TAihwV12Botg1Tg0prJZ3Fg+/EaoZPTptLqP9M09nb6zoDwxVqW5BLdYRcB34
th1sOBXpzQA0/1z/mEh9Fs4uc20k5FToDhTocf5kHOVCQkZWV/SLkj74+mhezzPm
bI2fI5phRDo8x4YJ60x6kBbDiMG7Mb4riFK1EyC0BtE28Lduo7hGbcm4eTInCIN4
T6t3svSo8wiaWeqPpvZimVVKGGyfbHlX1bYOx/JS/Le0h7uvkX/KRB3URDR84IqN
6hfdPO+T2oAUW+RH6WgkeOmhoZO0GJv8xMCFCh3G4x61g2mb5s6HAcsbQrhRAfT+
sQ3Wfxlf/E2Aesi7nhl+N9SrVSbkTVMTBWH1/OMg9ks78qvsOLhNZUIYBq/6jbZp
JNZOaHc29FoX2u+VdXzi7BePjrv8I5xMzLOK9kJta/u6Q8WwfGwihA7M5nkozRRe
`protect END_PROTECTED
