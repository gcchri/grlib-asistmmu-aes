`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4KC2+FCV1TSaiQz7UbB8Y+ytv89qheQIYtDvD6+NolKZP7YxxvfBmHmBZOGC4hip
oGBEKjnZLJpBHb5itBCwb3vkZzJ/X6oxvvyRl3sa11NDeGGZMlZEFE5VRGcndkiy
WBJOPn/BRPw8N7GACs7B2XUFO/EhL76PkM5IRupKP1hCd7sj43TNcP497XPKwSF0
JmEEH+YUHHS5kXlDk5vd7E2bIRHDRh44aXXUqtZTbFrHBk66BUlH8goq+9bq2g5w
PL0lUC+EgjyDdg7WlJExax65DgLfV7LwkrjM4mqEKk7fpnjQdRtgGhOZzugaqPS6
jRj9aQ1Lku6QwcAPwHItmg1MK0ABrr3HlhALgZdp7crYqJTJn/3zWcu2UwmnQZ6i
Q0Tejbo0+yjiGB8D6NmW9UQdc5fv2Au5a2Bjot+byNAGNFpf/2cMYlG2MMga39YA
Jm8KqsOyfWCGQOg6uULowpq6jxVMCOyDITrk6rJ6kr/l8Nkq1C6CoVaNZKmiaIxS
xTVzbw4caEOY2Ltuo1Q/ESuwJYH0o4jcLwe425JGj92POwacjOkWJ8JKgzE4XhIc
ltAiPZzLQCvlCTxZFdmviPdBnQxGELqMjLoacVbg+5QngBsza1uqjbEuvfpZoQ/D
fx0wn56E+OS4DopMBtfFIxb3F9ilm8JIMH3Y+aVpP+h0DZTGUEj50EEUzgX4HX5B
zxYiIjet+AnurEK70TGOuuBKYQsKuRpsmdTyEbpnmVCepGgmFLA50kiiLZDB0Ky4
aMIpbusmiDcyd0pgQ9ia8akXRYNuvYJ3lLmtxnzB4Vi1Ekqa4ALXwvCPjM5gndjA
VsgXKnOkdDU+DG8v0fmcMlK/A8A+qyUUhdP5/7QLI5+uAQyuTXPnvdTF6AIBoRBg
qFUgb5rWjZKqutXnKCZv2MTK/Ny3EmpA1w5/RX40xQAFFEV4znngAhEEmHjC3xJ2
pPR8d7D7XmVn/D5Ls1oTfmgTbZ8wZiur2PJH4wWFL+vIzdNIkHSmLcj56bdpApM0
NZkCIPgbzRkpSGkEMDw2l6MEvMLR2hGe0jmCgEDKw6bUh9mMNoKqkbNJiVSlwnWb
5ZfobpQqJMmTiFJxOOeweK51enuBPzes0zPt/nsLNaxM77dTmClVNCEh8f53Cw3C
agPDf/pCVb7XeTpFtWA2NFHu+Gyiw4NjpgfnNvC91bJtRi3fMGxmmr4iyblQSwKv
/SIqamYwZcsjKuZdCxHV4WbqptNaissDiK7FjHervvJLQBHcqV6AR2K/0NfGzBd2
sF8uAJSFrqWOVTg/BBTFHrR0Ntrv77qY/1KFZgLZpZBl0Rpbygnxfqwsj+NvcATA
k2XDThQ3BOc9m37awVo00+bz6w/5kOSPvnzUTSFG17/iZ7UgDZfQJ4TpfOHVg8qd
A2Mh0Xy5aKKaCL+S7rGq6M8IaXfDdolPFz/+HofjqZHom08VASHaq/OsVZdTvwQx
lUtQrdYiQKmVY4mijOYrp09BZK+lGfAH7RjNJFeHz/VUWReFs07Hyae8G8OVTVoC
jNHjGgbwAIz2xAXPJnN2Da0v4q92cV8XHzEDsql3N2biZoCvbkyEkKfUoa835sAo
EbLTeh/PFi60yJruXCTb14VKKJhf6zYevrNQwUH+5ERhlxaksiV5cNaYG7c5B9WR
MvQyE03ZSQc06zSlzgeeVlYCR0aySyff2ga9XxUBmrmZvX8HD7pjx9gBi7+pyJOK
xv1yl0oaKKlXVibjQYdu8xc5zkY80ZL648t3oHdRWUrVSK/RT1CBYQhf4aHWITJZ
DyQa9yBeY/FTAXrxLBcKyb/lrg+L4b/1XrZLBw7hmA00VZY1SLwN/8V3k+8BP0Kv
uW4zwX+cp8VJgu+cVauIV8schhhMmqc313+NXqn68dmn6vWSnMC1rgVBzJtOnw6q
l3T40cOrfV6eutBdahMY8v/IuI+ZW3LwuEtYJNaHxlgfU6JrefEKFqJbzlugJcqV
dDNUzdR+D+oTnowpdnFJKI/lKYcGfEmZ0taVIUjXiGbs5Mg/6wEPG8+Pg6F+z2n3
dNUhM0mVVjusFDGti6BlWncMRh478acIZXN+o3MuZrYYnRNdMne5Ah2SpfA8tBaz
3tPNFznJS5eDcK3YiMt/4W46Gzun+eFERQ0REFe7okUERcZNi35FKlHITo4cGNeF
VWZ+eVXRUX6349jx894wUVU0Qfgpz+2M7D4nJ157QulJcqyES398feHMHO1KeZMr
AtuYI7KGUSDTwgm+pIsyusEhlEWJEmspEQ0VL82ZinYfVgZ8lTtORisGwI1QR7Lk
tOdWuhsn9SCjL6Ux58X40S0qrTe6fBU3PBmjhiR+5InCJwIXklryLrNthTLuEx0i
LpaDgV+htHdRPPl++Y186jguqxq8nV0MJzqgn1+RW5hUDHRoYvq+bNeq2uREKFu/
FZ+RGALcbq2Xm/jFeK89fqepMfEZKJdOLkZxXXsjHR5CPoZQY1uhGMqxEJK258sA
Q7SNuuyvA3nHqEP2LeDt1kIZ8GwawdvsKlmKqoH29c/Q7LjV18u7/c3EqEdxvHoE
cEswf5uo0+oLnwz2kYNuyVfxjg/UjNS5exx63MsNtbWtr4WsPoDmTq3vTB6nMMai
tRS3KY3Lrern90zpFgZjFN5FEeaZ/AUb19HVPcDryZs0TiENqneQuYAWcNtXD16u
IyXqdDZoM3BhZgo/wGG5lo6MjcdsQr9YeWQwlmrcFhbcILn27d4N+x4fM3Vpi3O4
4gaf6wmGycLeJ66fLVsRJQ==
`protect END_PROTECTED
