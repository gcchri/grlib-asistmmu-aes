`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pWQhpwGAhC+E7l5aia1ve0Ll/KwAD7UkGrGurpc9a/jiV+GyZ6nNTYpqgrvIk0ne
zDAKmrxF6HdxvzA3hMn+N1vK1wtYvQsS80k4y3deBvtTrAs571MVcHeU5++IjIY+
K/X4YZgLhKmnuD1zqzWcVjpJT6q6jxJvR4DqLZ7mafEYEHsimNa7HvGu1xyUZjQ0
rQkMeI4DOWl8s5Ct7tUk/4nZkUEhWbApmmVjmp8tOmaK9/4iH33RTKjZr70QkYcy
yUBh7EpS6/4lkVfiP7FveKRsaQhlE71KBNHZlPi9VajyPZTJs5amkMk+aEqxS2i1
U7iehdLlOury1XMbBzps+cuBqkymU1RPwZwvcTAm+vdFF85kFuNfnKvajobpyFg4
iv4Mo8bbTKeOvsW17Jn4I6NgOZFehDe/bPNEFNTLZqHHmQYcdl2sh1ABVJ77274T
RIBS/cpJblwFjnDvLVbRLBB8gcXh04I0sbl9+JvrkRWF1tZnfi9RRPOF37Skz6FG
`protect END_PROTECTED
