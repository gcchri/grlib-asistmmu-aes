`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FvBxOfzhjJDKgrV+EuADe1CVP8tW/NA4oR7OeD1O46/lwCf7Swc4wLNpCUBlngnM
uUGNDWNbc8JXDpLDvsygkowBfDrAmvc9p7stBBNHtjeaJgJvbtnlVWgLOyASmJk4
XNf0wMcW0OKsu7OhH6bz0bqaeNQ00pTReM8hBA2tVBgTZX3S2UnzhCnlaa9Gapbc
x5mbVKEptfhhUViNBSHrfuuc4bxBeNTUanXtJ7/7AnivrzOyr552ZRnH36J46PNa
Z8ofBZ3Rk8Sl5PHmVibBS7sZUI8wCBP6RgCd3KWz5u9VFt2kZA9xWHaeadEZ93YJ
T4uUpob31YmX0u0anlMF2OnL2+EeuuT8LH0/cv5FxkFf3tqpn4ZTM1KuTKpHSb9r
3XEc6Zjrx3VUc5h3BtXo23T9VS69sLg/4cg/Ldh3c704tZKaFDYqbTIR8GQUdz9l
xDtMXNdy3CEkfKzxZqwX7IA2TrJ89KHfyuVzYEqU8XiKLjnq7GmziH84HrJSbhKs
8AuXrt/Jic/F/Z/zOkMspntNmTb2CqY4QZYwN0kW8GAcKROcaI05E+rWEBAss+2b
AxC8cxzcSWXmcgRYFbXR/gm36BQJL3/JtxjDS9of6jZ9utN0dc2JXNprW8zKaSV3
e6u+JVvXP8VSQQ4gwiwN5RCegti/CjKNkCCAUBOPQF1IkV8Xwe+G5XDf89rcp2AC
hQIGQMco0h6UlTBn7pvHIbOp7WccZMf2cwXtyPx+p4FhFyeCIhU7BPSfIZdKSyAL
pOvuYsDYh7q/8ENUOJ3YzPVwAOAMYd/hYcjawXThoA5vuYjWNCvGvlCZK7xH8YgA
kYmu8deYuaYWW8OLa3iAFJIfB1jWbQmS1XL2+9et113Xi7qI31wrCk643uVpLkIT
1Pb6uUZ8kxMOVtBQejViAdgExL8ZH6boeVZWXvM1iHizujL5kqE9oslw5/FoHsc+
`protect END_PROTECTED
