`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DQd85Z/rn09fIC7+fW4J1BUyG6ozkrWIrtsQlUwd+lq5u6FzVBeNWc13lgJz1Hrd
KUdesmOIJU0GrYqvvTE5jFEOKHXvyOvQlyVn7xb27CmzDdNuTC1RrHNGlooamOwL
M8zMLFKCYrcCb/fdLcxGX6DsD2NZOPZVU3BZagNw7ohCQPOML0CU4rXtv2h4pesh
q++GTYPgAuYw/6DPHTuRw7zjYEYxVZN1ge/4mbItGY1qYXnws+DL9JBZ5u4J2IxF
WJTZRa8ieNWrxxBc1G5Pbx3Iukkt1/T85XDxgI1xYUcTUeF0Kxh7X2PGjpmU3qkT
GyR5ZCiKj59Cj334Yx0VpY7XHVuVewpdfQHIx+KJpeBGXyRsI7wE6Q9gM77mzLWU
W75eFQ0dYnX8+0+YnPPlOeHx5SVcPS+WXsFXfpORr1hcMwLCdg5nWc1hgiwd1Cg+
OnykICopQEhmH8HtPgL9oSS1/PxnwqixXx67uLB+81BH/9HyHQiONeMI/HJiT4ZN
Nww5Orfbj1xe7HlbifQH7Ek/xXMtRnumNp7K7SXStK/YQ1zB+AEqQ2up4dLoNogv
zpex2OYlsES0ebw8n/0nPg+A5LjekhPgw5RzBF7gelrP1kyrC/hUomi2LbSsyRnM
qsnXx4KDyb57Yt+D83f1wzXTKA8YWqogcmecMPf7xXGsYzKGEnzcqCPmH+hynPT5
s4T475dREPe2W8kPNWXLfWWvAdyZ45UmxEHo628TdAP0UOVmW1npACBwDKI2txNe
`protect END_PROTECTED
