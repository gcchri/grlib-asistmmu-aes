`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qjy3H29lyGnRHQuD3huIOmk/afIZmcr2nnGyGqdgdUukls8vRMwe44dZJi73p+zj
vfReyvuak6PYDZ5H0Rua7ODv31IyPds3gRMDf7fxcckKhlSa8fIRb007eklp3TgU
C7IBuEfL7IlJmoJshTaih9SlCP6MaTBpPgmCV3J45gu10zkQBBCnqKL6GuvcNiBN
RPVrc+LcfebD9Rs2LNTuJvVV66gsC3Lc+1ExykzPateG3yvSif4ui0rmEgVAaNnk
Q96KeDGL2tfU1mGCNy/1MsaCGd1zyEPMoJHUWdHZSCj1Vxm9VvE5Kj2k+aRF6wAO
wfg/OO+zTI3nhWz2Wl8YgrrGuCK8N30+lb0F4WYz7jKrvVKSpiIpcsDi8sKT3sSd
EgaU1mKxRsmkAS/gnLskh2lS6bw+C82hyuFwAq778tO2JLyj4VsziXgrMMjzuHqM
EHk6QqxO5VW4v3t6ySwFV7rr+YSaClF5PUVjljklPMSsfbDxDppoKCjLNVDIusyZ
Sp/6jKg06z4d2hAbO2BM+6nhJTFoY5x4jOCqhqIHywZ4/WgwnVt4XIipuOwgnNFD
5rNKzDcKOYeZvKSQfAxDtXLxUu1MMVlNmTjfhBvSqxnS67dghkyCWWAlKO5DanyG
+kMNhLTkAzV8y2VuTHBsYNAFIPLxpOvzVtbs1tiACc3Bl+pLEbI5j8UDMdBX4/P7
eYusLVSO7iM8zzOl5ybxJu0RNaxb7rOa2oH5+iOYz1zoapXNQ/goAZJgBO7l/TvQ
4g1MSxMMBh+cYTIqST9NqPbYjtaAcbcnx4ZhUK15tVz6ccR3KX6kzROJzwPAm9rp
Q5S6KPb4obY94vFmoSb92Ug5s6vJWsUmIxLzNgHJhMaUSWXbPtgdGJx1BfkggRk1
rH0PdMUwLY+dn+b5qp7/UySbnMedg70B+but/FHMtEXV7tA0zjX4C1dAViM4vQRm
eTRZHcMhgax7ccUO6xeiqy9YNA06tx2hlUO4Pzq3mRjXu/xGi2OEOHGqkTpCNM1d
5osIQ5NVFG96I7i6UjD/7nsgxNEJkWMpeEmsAkTJOCtizgzyrDshF8mbK4Gk4q6P
Okkz7ZOSktGoy7N+JLVtCcaHNIFSf4GLlJDX2HCuVvKhvmR/z5EtxI8okHqye+HZ
P7Ty4AYUcNZkeuXHrnODQ+ETu19EJTEyt01CwxKqh+lpp2ecbs+bK4+KyX7CRkH2
KA67wtVhJ6aCa37VTmTkJZldlvfmCZC5KkQ3NXEHS5LwJ/A48qqgfYDiK17vxb1V
67saR/H0aKZjHq3rYBgo/jv0f/e5PgW3Mnuwfb2wH8cttebjj3HM+wcx56rBCjBF
WYH4Vvsq6fZLmG1bbUrk/A+cncirJvYco+OKK3HbBgl8y+nAOpesITzaDFF/gJcp
VFAFl4kqLFjChNR/PpfxEm+4tVof8HeI0DncRws0wk4+wZU2aNEuYXBlkBFTnJVP
q0a2mcjBog1m41D9sAYpLuE9gtpLSRsGiMaJcore15BNzwyY8zecGjdSfzQ3mZWW
ZhUtd3oEzDKxxbk4vWO9uknsihGcO1/jNN4FnQh0YV8PWek+BQuwJ1UBY+GdscZs
6YNLV4VnpbT5e+Yo4mZqEhoOmBMX4inwuF7MRpFPQ1/FpGfCm2mZx5eX5oipQHhc
7nHgqqR4QS/Sq5g4gW+wbbhI7GB+USyxafG+WVheEc5pErIA2bKMJBwFOsGPfogU
BS/n/7oqsxEaMMASmh5vpBzdZnFIy2+nkM0dAVFzPYBxcalPZNWezNE17LMbqiAY
z9NJozWXHIMPUuRYdB+1O10vSfmZTHDXq1qWVKgcacEwuqpNnIa/fUhzbuKXsBGf
VKNviwecQLMCS0j7Hkgn9HuzqTxv6gI+q+zfEXe+M9I7fN7Y6H5bsGMupzrMpNy2
oAfx6fP80HjZRbUzu67TsiNbdGeTbwfcD+g1kr49nqYZXa/nWZFJ3Tr0VuygnoI+
7u5iGTNQRRBPQ9rxY42jZo+WJ7FJEl99ipsuB0WkzWTGLZpHvAm90HamO3qpO5WZ
9N04fPIQLl+QeYQytR1ME2uBxWNhazeewwFROicymkxk83YlZeHqNcWMuDWv89kZ
vQdXrkeCbajPhMh43j7GowY1q4hFpGYMhkKA2lpaF+bVlZ26xuzFOxDZxdfsHNKc
Q9g9tGTBvC2uTSg8Q0N8qvPOmkNPez2Vf96b6t4tVeOAfkPdandLwXq7IGWxEonX
cLTKXMQl7iDNomxj0bbwmn/rBgGYfev+ns4fKlxupSgWNBEmFk3nzAUWWfxSRCDs
I6ZAFhWKmhZwkfkbxeVZQlpo0nnrnIE+pxeRffwsWz7yixs3I+ToCRDqEmXu8klN
FcKyKe1BkGzs4aco7QV7pfQ0QV4hcQ9Q1gZYo38Hv9oGy4FnBpCt263ng9f45JRA
PzGRqW0i4u3+t/uPwb0ZCpadux/kvjQnTAsrD5SkmZSgDOqGq5aJi7N8PGAdI+US
1twsfqGbKMe0eRM3kb2iw6Eh0ZfDTZ0BW+vs+02UsGH2V+o2ORaWqSuTZplWhYGW
I0zFOCfLNy8ooI5AXvNNHHisoDCT226gsXfOHE1fBX3NaDv7FrLgrxx10dJB9kNg
Tt9B/TFDvNuDPLLAKi3ta3TNUR5y1LJavctpPIZ9gax3WEVL3el+clHRIcQoQ/XZ
eCE7zMCNB7++TtqeGUG+M3frnAEUIaoe5CEoaJephSzbl+9asaxG4wCPpuW3zNVa
PtzNa2XVygGvMzlF2mpu4Thck3uLRHV5WCEsIdj0wOPK8XNcSHHhFomuqsZBEAYk
S/OQi/VF4sZ0YXdKW8bXQQBkdjHuL1tK19kptj+70M4kRS04fbAaKZt6IpPmzBAo
HPv96wdSgBrKFt8OqMCiEdIZ65xcFqHfovwe0w/4tqV7ZPCCfXQcb9IXZPt9MoJd
mCrP+Ow3xI0YZ4liDpK/C+Ol1uAOEkozL8uU1oGI4hTN8SgAYAHgGYHSGV4OA0IE
FLf+AHw1S8C0QEBBJfrhy9pzTDrnXf9exMDMmX7kuksddIJxfMMmQ9H9Oiiqp3hn
0XpSGY9gS4PEEY+JORcSzmAi7czq1h4fTYo9l0ci8SaW9n4hd8ie7PDtvAaluQw2
PVZsOiWK4mggAqO8WcH7Vpu2aBvSRrdHsNkGOTcbQDfFG0XJGXiP1GeQbVRlHJR0
mhyZSXTSR/+Wp9GxUJ33//jz2PxwRQmr9kzCe/a64DC+Lgh3cOUqUHgEBsz24pBv
gPqYk2xMRUmQUN5uzucZa8pXHpXRVgkfoXDIYGu70aoLSZCMXv9i7gxserwEMF1R
vp4VS+Fc4zp5P1D1uxl8XCiNSUIdMdMiN69nJpqlMgWmudeIjbDKWdagAYWmu0EJ
mJSNX/kmWvLq3kH9FByEDb0o+BxqrizyF5ecoDuhiJFO0rnExpnJYoQwOWr7Mlj8
kg42lM8u8FgBVDNLkIHLr9SfvGxZoMSVQH8MT8ukekzHs+9k3AU2xVA22mXepAIW
wuWqrziRomwkN3TtmHvxP19SdSSYbk2npkU4N94Land19RUkheahYJPZTLNh9ITf
12iYgLtYScC2ztQNiJH5lElGLgUacLHF3FFkhlz7IhgPRUazsv3DGB5tFiVNEzoR
Qu4wKcRrFxNEgppc7LQWUK6mmPyIopknUjHJIFL7MXIFnwxqfZ78beoZaamrJcbt
vcCr4fVIG+5EW1D9hdnFhI4umuDLUMoB+4tQEdwr0Lv0VMnyq6/PVyToUH48sjht
6Gb0NLnZPyvSvdNc+M4JeOkKvvDLc2mxjcfsFtGeoIdwqGQRkFzR1fzlLS2XZ8FI
DtNXYz2AFFd/zbVTwjTcRx6z6gBwSN721GxJ6VzMqRc7vvA7tVNiAQ5mYDc80PEc
c+EFvXDeRU5aNaCJxPTzUkdu1qz1/mCPck03oErPHTgKSrrYyV4CWj6gR/OK63T/
S2qmR8HKGH5/B2JYjO05C1JX3a2x3XjG2YTl2Se3i8yI6VorRAH2Ee5vQTxh1dgD
knV+1lT+qSNji5O3ytz42BkYR+RQxxUT4MPdxF+ZGf8mcw/8NHxJuD8hcwTM735j
dZXieYPOaI9V3f7z2f6oplm6fJZ7JTXjFiA7KjEnZ+Ly1gQngLgb7mC+ZNsIiyNX
9Gh76UzgFwhjHJnK9nnYHLHlKabqrzCY9LnNdsZ1lmipddIknB2iTUOiVCCw8/AP
dui6rXN+g31xOS8qRHecEhClLlnzYmjERHHsfITIZk77XhuVsiayW+RBd0BUJYX2
jg2Zuh5aE/ru2DwNP4wPHDfOigQfp9Uv2QZnExljVq9nn8SbSZSRx9I0qhMpHm7+
JjBzMPtfbJeTa5Gd5DuOX68xrff/Y0xggCZbicbXLbyS6zqmNSv8ogYAOtUHCKvr
joItObQ2k6b2iyjUEIqgXQmHR6WUnpQoXlQFjK/hYiyyv+z5sbsVDld27QHK1dvM
Y/Nml6+1BZgoNkYStKThP+OBfCO873Cbq/FdnMz/CV6xOuh2aFSaTMkgoFevcU5y
X0mWyIHlqTHISWcC6Ir1prKTnGjcSf/HSPqHvkNvC4HdW+D1ojvqkSQScqcpl1d3
hjKPnkSB07GYOjYnoBPyiYrFZV2H0F/wfMm+iG6/6EBvvbGjtW6xkH8ONXeMAJRx
tP8rYud9FQgQvPlzd27At+sCW+4+ge884ndMN2Np+r3oPaXLYEO2Q089bWA2IuOX
tXjHRuwNRyQ4u1no4fgVSDOK11y86oyKow3RiLYTmCy8ts8AkXrpbuwsOz5dzPUh
QfB85KtWsWRIMABtL32nyZelQ9srINTp77pBNY9fyczTJzLkVZyJW5q2A2Al445H
X26ifmz/2ID8tG8arp7kvh4ywmkzwFz+SGxbzNGItE9G9rylQfooz+kqtrsAciIP
9Lna5paoylCCLUEKB885l3DdmqZkmHgO5wW+aKBuumdOMFZnBKPcMGDK3ljasMAB
RonCyfY+x8+UKBY/PRwVOTzJcuCde8KU6P1t4rqCwL6Q0Jw0jiwXXIfkWKynXZtP
1fpFVEWVViuLttSU1CtbpObWU0ZFS7+hG4iZGARkgBYeOGCeYVPyi1SlvXHgBbR2
bzqxgJBBGn7V1HDs4kZTQ6vYwJVnAzpIF5LPSkqmkZVTx10jdF7u99OIMtwlN7dU
UpgDYqoRm4sxupAPGn95k7ovTzNlZg9DAPo5aOvDw60sC/+utjujTuVVMOGy/8ac
pXUcIucjM12wI95Fzb2YbRmDcs1MswjCszEGrfym4NAAm6V+ooW5+dJyuDcdHLqG
kfXtLay4X30wueJT8rVl0jBVNmbtsD7yyeVkmVrVr6SgydvCgfszyrGwDIYLYHOl
8ig9ei205SghoNCwHrXbTohfZW1kl8JFxUuhqS/P9+hQ7g8rye82aD9i/P1jKK/a
Kg0zJINfdlTEwNoqKPSnLSzksjJbx68QELSLJEhlBReYhQX630vFQJk+JEAdAmvd
HSWElA00aap5DykjOzC9sHqjR+K5KaHdp2MmUFlarlop20Fyo5GU1XinfjJxy7if
9JrVAG7CWOh/tA5ZTZofMeyyOOww4JDoMz1TcAXBYHWdFquKnztvYq5UUHuU6+bb
Ohv897TgYn7s/7KQacRDctbb4GKVuwOMtB5JVBoRhuqHCOoDIFOEEh88cYTNYIUy
+z90w/RXt1rNNOq9GcBM/QSrcn+rqZUi/SLoXpJp62XCmlyEQNKo5b8y+n0xyTBt
1owaZdjvdp5t6ao0HQIMYgBihe1tOV10RLGqIGleBeNpy5uFPEqEkEpGdlXCx5St
ZFS++34SW8hxNBhjDZ9Z3ZYn87l/W8S4EQXyQ1C+QXV2DVKX7/GsJplox21X5xIX
fxQTKZBSxoI1htVjFt7HynizsN7o0R2KFNQfzblVatLuQHTK+/u2YbGcyN/49WOe
Sf1XfD/a6RZ8OlcEiGuXs18qw4nTatLZCkl4Jj6kaD8YPxa4O4fpZM/PB24rQ13U
+QBXNhLOHUTR5QF+0lHZ0Rk8quyQ7TVTihffGp6VYGhyAN0qy7f5OpGDpCW5ETv3
6BxRmoyFgz44waSLdfUzvBb1CPsJBRirm0yDtz09A01wG5B0AJ5ijOeGsmU345pC
jo8dNibahaX87bdh2BbudLGZLp2GYTes98pgyZzBfnJv26jIun7bDH/AWbaCL6aJ
7XDqCl4M7s8r+Oa2H4rm1fV/pnGlA7altYoY+a1WAacSoXuUfXc6kqHd43qcEfn3
4WQbFTNRwLBn959/+u4ue/qwoGujOteniMddQNqmDV/FvPc+UASZsCxjMmxazEc2
HyNyj99pvAnxQ62hs6OnE7MWRTZWjNDpjsURfRX3rIT5e7XUD5TIOocmdM49fgki
31Rf3KcmlWRUNN2Mn7WVV6n0tKEmEB40HgliiqGeYK+P0JZvQxixJLUdqljmHS2E
XETJIVHMCRETo+500Lh4GHX8QzACk/P+dcbxwqzinyLkJ/5VhDIkbEku5hu5OE+S
0EPgNM1N1cGIqR8wgwGDZlfUM9JSsQyZPi0SrHeSx7nMweR9AwD3hO48iWqa5K0/
FK3xWByivO0eQU9eJe+qCt7dtbji0QUhp50zvx2m786rxgHHvclOQ3BEQRmOoxMj
Fu6hm8ZyqM6l5+PX8epH0WBADM6A/tSpcD5vcReI1Decqg8QLMnwrRbeH3OS2ci1
Go+iKkRn4S693JdN1ozhNCKZPpSbZS8eYuJytuil+iN4CVpa3O3c23mxQHmaQCmn
pKqBMNwAkevjmsYRtBZvhAM9CP4OAF38tjeolxGoNFbi8bc119YVgzRCDJlYU2iD
6rY7e7AKtQNpECLxTNYokGrVuZsvmp8WRCwvwOg76iNuNTqdVEhc51UEoLSatSiT
/GFvE1zBpYG4laU6IXKN/z9M2l2P2vVDXCaU52ztEC51Th16dGurNIwuUsV8AVJv
ZJcXgbFEiKE018+B67L9nCFZngWcgYZjRlj0S8D5YAHudkrOoHfURWidBTM5A89t
6M37uFw6YmPT7laH4UQwVNS2Bx+sid+ZJEu+KEDr4zMM+aZ4U1Noxd6ud61RA89W
wMD82oF9jdzPJEgFsJ5zauSws6gdKe3/fhNPeu97dtqni5RnAZ5V7Vdi9qEeARWr
PV0MzWpJCnVuPF5ksinlKB7AzzXr92OnY6IgyynUJcUnwtN/tRkQLG7MFsDiuFbp
Sd+YgQbnAI3i4Ju6vpVsRSQJox9laWP5KFkMrvt61C65fpEkHkEdYnsfVhYysqyA
iCgEVMmo2mkXjyM3AMvkWJb+nJ9re4n36LXgZoIidbUWPSuD6zItjVI1a4ibKK5R
PRBFI04bE0L1DKHcjYaSLHUR5r0+VPLSlt9nYcD07OpYikpaLeo9L6T3x6hkH5pE
Fqz9+sPKaC7fYYYQhSbvPirHVYK8FhkHzWn1o++ydOZUrwunSDa3NYq+rjkXxvEJ
Yz+jeY7UjYo5r3hmpzFjgDN3hY9zIUAxRnLNROH+NW7puNWePbJngLxoflb7J7ab
IHd8pXr4Y4aPdW1EoINepof7mtcBFS6R0gH4xsQSsgq7h1uijMZqEsC8FqSO3SkK
BkgC41v4eyf378nY9VGXv/KZyGDPxpp/PmCb3teD8/4fL5sBbDWDnfwsb5xO+HgI
tQfAULJasTQe3QYanDDkuI2unjRAEYNNFTPGWf5hfuTKcmYvVkPwiOhfUMANANZM
Zm9l3mNzrrTP3DxhcuFZqLiJuEKJwLJhwSmpIq/RjSfXdg2VHVeYPlEUJVBC3RSU
xEzPqT8tHv2rPEyxx9c+kCkv4YGEkK4Tr6osZmyUWvPGHmRCqFDj8RDoaI+5IrcC
0F2XnyepdXI7Yck9wmviBd+f4W1qkZ5RiiutbkDhPCY/bpiS/2HxYQ7EGVTeRo/q
mqFrfdW4k8VBM5A2bliZzIR/MI4X9M8GzncaXxVMnjzR4nFzNuvXTE6deTOCyaai
DVIorpbBiPD551KXGQ4wpAOi217JjKS3oHclawDQhNPdDsOTako2ZVD3lYk3HJmn
/hdPzPkV36u/88CiYCSkKfOodSMte/c2vywX8W7+e2J6cxGjJQ3IoAVMJDNAe9a+
SegfR2oH6tgP9RyBy7ObCwl+A4pIxs0TlKxdVDTUkwBemyMyAwzr5139p6D85aAk
9PHeZkgcwq9zS88nlc8IuF5A0K9zNWvIDV6iE0eqkUqi3knb5DwhPnChB0nJnm3Z
OJjVaJsxvXwGPGDrvMvWs24Gues2qpMrL+Ct5W7XP1m3NfcqXgI/3nhvFfhnLg3o
cTkBZ9V9YqhR4QW6q02J//OH/KDZAqQ67MAlfYqwG5J5Dr0dD7otBSfd1huUyKf7
EWS5fK0W6rXhbiUQU2y8ZNgfFeZBDm6VT+/m0S2WPImaCEPeM9nF9bpY6wXhocMP
bPRJ+/chLSGGiAaDRKZ7Dv4ShdOF1911+bdTYUaD5P1SEyenyFlrVDVIPByNG3fw
J/mFLgXGJm/aDd+wgntr81Ft9txtwa1odvrGuhTl5TJl+qkL2XiMMOP25ZPYCvyl
paQZCV68yAFH0r34qEMfK3LOPefnWyCv1MAvIJyNwgMsKOkDDl7tm3calNGFpkiW
6DyTP2sengdkQ77wO5tdt9TenWEIr8xuBClGlKafd2Djgc+6avhFJpN1NEA1v8uI
ItmwDD8B0OBp3xCjdvLxrfkO9W+bAotTxyXxd7kJ2xaxiPJhc5RfDPynwGeV9wrR
eML9ZZUn3LTYrKSEYdFEcWwU86mo3PvgCTJsY+7MZSYBM+BqH4yTGLMMtzouK7OZ
x0OygFaKftLZKK0Wiyu2ldFvqNOIFqP5PufyHdZiPkfvy9IdXGbBanUMvW8bMUlS
0K3i4ql5rTiCAuHy8IaCDFrcdg6kz/D2hf5YcMyuia9g/EKJ3Gdo1S/mh54PpzwN
`protect END_PROTECTED
