`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOrdrO3O+C9QehxzkvJ0cXgHclMSFlYolhEBh/yV0oi/l1JEiCbEBDc+DZVhEX8f
2ef5ZvoRJq26CBi71GTr3iVIZOouDxWsJYb+4wAqmLvw9CXZZfjoTu4cJckp+mGe
Gr3a+VCeCaNZD1/RMowFf+ZhjPFuB32p51Oaw/EC1miSTEVCagx0HQSAivwuQ7Vn
ayuUkR8m52FCSSTDZGiLyS3Rn3rNZwl+ThZhV4tIzLslW+YutcPR4hKH+AeAVBJW
F8jRIPO4x/Gl6pU1atz48DVghtDnCqDli7aceHy9nL3nhth8WDK7AUjRc7GRlBJK
I9mCGdlKiBiQdDT0RhFjzUzfssOOXxn8rxJngMvEXggsDajqh9c/590O5FZK0nF+
SH3VYaFH2Z139oCNh9EqxG/o1M3yrLIU9cZ7+SoCAGLWkyG5Gnr/aVbOfITK9k+V
iBGMRucC5i9b2yk2pMMN/RQ9lJdahnUzEX+79xzWy3XsNV2v4usCr369IPpPLPhb
`protect END_PROTECTED
