`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X4fcA1U7PiY79P4rV6/tE9WBeEblU07o562GmETuSjiEFqfliDwRvtcqE6pbvoTw
nkFzvxsWU9ZzMSvqz58fDPb5xqqxpMEsmKs7ua8VRGld5qj6KHidSStLW28lqifG
mCUtkHRSNJgAZsjR3pA1PhGZ8wqrmEFsKD4IaAY+KPpFrc9jjAfazBr7Ho9eJ/yU
IWnuoroRG1LRbo7NUVE6oTX0f1lZz5e7+6cMNZyFcRastMarkhSjY3hltGVO38lp
g23dhwhjHhpnHrxzS9Lecl4WIpf1QLxN8EZCiB6HQZGtebjZb2pIrIwgCHv9erT2
870dTdant3vC23lbF/3WHCWngoSkK51TN9BhnmWTrFOLzGado26oMD85b/4Ru66K
2zTuNnXD+/fikMVBIM/QufFEEUzDjxuWqQnFF3BL3nL/im22o3NN5hqxYFlW9vWQ
`protect END_PROTECTED
