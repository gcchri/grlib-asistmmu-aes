`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kBtwSiFqMgIsniaTAq4M4cOiKgnivVBPYYe4BBMXkaUKhkQXTQoj1v9uCLTuwTV1
UzVfCQw1w1LN+pBu7PPwpbDabZBIeiKulkTOeUqGX58JrsjiTtIvt7HuuTEdGEPN
GvsncNM2vOX4gcdnYeYqu65m+UeN4xnOfKrlr6tIcNKhNazGfKNDOBxNEPi5caxl
DEn4FPv8qp56hoQbZaFtBBri7/G4DLn3OYj5fL+9qRJtbouGCt89NkFaSao3PTak
KiZdI6xAI1V82BzdI/fwMFz49FX9p1039hhp6K18x0T2WLBTyOk7aR/kClsHghzf
9lEKSTkAtkcq4QWPs5sX+dqqyex9jBqKbu8zMhGlP99NXNSXHpJUZsMuRTeSvSQ8
CzpfqlwJ5wGjYU4mp/rEGQ==
`protect END_PROTECTED
