`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vUjbcet5Cg+WhFucof2EBdbpCI9ckaPpTogGe0FniKYirRNttGzmssl0BMJeKf/0
GvwjT/rG/sgCrQ4/jowbcQjqUBE4sZZJMVYaaz9jDk231gruh6ER4kx5piq9lYOa
OZFCamjl/qsqZBlWFqjtzGCnmzFmmfNfRdQGq2PHtk6NSf1yF7jmTcPauXRHYcIJ
m4353796XfIzzzqHxkDTuNVHysOBLHwvrxwLkuDV8sPlO1RquDlgDHTMj1E9Ii1L
aijU4L/qu006rKpJSANZ8ATfI+JG9uHvETsc2XrlMvKBvATfNEaX46wFyqSF0C6x
TRwrWJMGt+Qn9JZq449SoBYE3RYDB6mShVDBpmW2FTnPcQj05r8Glf9ZurtwkOcD
bPMmUDOwgXvZXSC9XlRiL16BasC9qO5U8wxNyPicYjex0d4QPIzJ2ASqIt5a0lCc
hHmGeW6EGtpggAIKxYLeSo/8vRrwrgSMhhiR9yrHTV0P9Aw+bCjAZxW8MdLMJWZ/
ahoFoSpbdPD/VQa0Zrs+Eapw9gP9QSrnuuPfKfju6BRboWFb6BQmKiL2ZhAOLUZY
964BIN8eLneKENV/kmsAPRd4nJFCOim2Pm6cJ8qaSYiD/DqFUxwTme3NpsflPr+c
n/BCv5J8x984g5HlszMqY2RHgTa6RufXSsazkSUrmg0v3GfYYqF+j7/XRrt+dzSg
GXEJ4tDMdtVP2+V/nyDPg0NVracKej3Xs23nYk7tE5ihmEQwDmZOByIsVRh3t0Ir
G5G7TX+LdVha5LiUVKW4F2HV4DDnIAlQbh7C8zg9K0J8BtiIekjpZrWX9dEFwHCD
`protect END_PROTECTED
