`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPKFxcTTR29+FBNc5TPCsdiW21leUviTAMg3N/ECYx3twW2HuJt/CbRvmOcnSnYq
9CeojT41V9FEVrZPb6iRUv7vjWIUeNxNPxKKjE30vL6oHVLKTVA5+w4kKDPdKiFF
JFDZ7eim+D78NCN/zIP6iCgeXCKOOP7yRvJ+M9GFc/KJY30fqvfHQb1wt6ZaQT/c
H9NHGpvVCIjWSCcFVxZTxbYDmQUZ8NZm3wjIAZuCoRgfvBvEEYgiyn4R9+5Qz5Rl
wJblOR4baDdYMyasfDD1/EMNvKXNEao/ca13CCb24ugnTEfPb7Z8L5ee9DyyJSIR
NsZoXIylRsXMLuBjMHKhQuvpdhNjFIFj9Hvu7wVFfCbH3+PIZ2XKAFdHpsFl/osn
2+m4aFwIbYkxY3X+9BMbSJOfkFiOSWcVdSYv5VeYvrV/HzQ/qlEHJ+msQst/xWdX
EvwmJeqs5KFUAsAGwTISxcC4aHR532FSPbC5r9ZpyED+/RerKFQd353kICqP+5SC
rkgrbTsSa2OpQnouxsjkTeDxo/BllRNbQnrrF5o1kq3lQkMwMXfYlEHv+6f4HAYO
v9jLvJShhaBsB3FQd3FnkPxlNRmkGxwDmF8iKhTZwdChJm6WZAzeLod5npPiG8y+
TtYj0EguSkE3hqrICw4WmXmcMoDe1k/xktqpYyGe2hJxXtiZXbnFpqh7bPWOHT6d
ltgHQB6doeKKtIWx4jDDT2HdJb9jkUDfKwDCd/YTgc2HcAX1DMWb31lDBpS4NSbt
nszXwLKO7rLXyXRDHL3ahI+RnHA+OHFuDYKVb2fTgzbTnwGr+IxiktxJT5THgn5Z
O8SlcItinrcvgDzOIeGT6976TQGu6q2wE7CFUxOfuVfNg1kj9R+R2UUpR1cauMKg
o/4FtSml/N8xMu/fsRAwkyf4heS61x2SL6a1z7LWqnYD4ufa8xCN1fnWnFbY3iBE
QNJ1XpF7RRFKtNZ1QtCsBKnrZOt30wNKGv4JveXBBA193FVv5/tl9OCWm+uJi/U2
avOmZQxyaunXxuFaLjgEibbSHfdLldST5tn2JM4QGITp/xLJx2lIMesM55EMf9jx
+anzOP9j/GoTxIBoOeZwDQJpxPdKpst30Ao1gND0AzdBObwF6GKxl38q+Sm2Jpos
RWtxvLwC5cd7Zxc2MHcp/cN8Qy9CraYpO7AFz6LSBAI9Cni3qWxzmwJj6Yngshxe
7mJC4DCW0Ua3FqrlaKC0pmFozXabhiBcsgFXaufJynJQNP3dRe0QkkJJ/2V1Y5xR
SZjbyFWjnvmVrJKe4NZanTLnFYhLGp+Fg2VM++xW5s/nRq9nLErT7c/l+SKbn+X6
OfOTpVmxvgNdgcH6WPIjENF3Tsl+mOIiCz5szb3O+UUTPZHPcPRI0oKTtt+B/5Rl
bsJZH1wG6i0p/LLc6VAEcxgN7fyp+UnxBWj5MqJQ0gK7lgWbxZtkeblB2jAbtz2m
jCkdnJBLZB0kYsCK01TlxFVDx/X8l6Zy9zioy8Cizjg=
`protect END_PROTECTED
