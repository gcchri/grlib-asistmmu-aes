`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1txwvg27pHrut1jwH++NnzVQM55tFC6Ob98W8m2ErUBlyjUXGxiajj13UJVIv1qg
yGeEkzvn3XJYsuLM75T+GH3CSIezL+CmPCgAMXFQ3ENG/yCoOWpaF/swY9QOyAWH
nvp2GjV00DZl9DZAhCEKyTJOigOPd2rOQoQK1PfkENq+6XjKnIgCbU1Td3Tb3g8q
tYss8bgazqUaggDbGqa7XD1rntbLXItv+235i27gAeSA+q9EGtKC2n3yzaN1vBpQ
DUh2QAVkmqfTqmAEODqDg9vSs0nXWZXW6dBZSgh435+qQCyTNWVpX/CPWEHvg5Hl
kq7c6x6uNqa7jNNJ41w9YDT+QqesNPsgfzgJ0eHnMsreH8N9/OjxYJSKeNBGTNmy
s4Gi/tVkUTRzpce/i4r+Xuw/9Ec+A1x9ObFCiYlB5q/mhLJ5Qi1uRHHcR1YeubiI
IoFuF7FRD4nBGe8rV/tDPlqUObaHMoHdhxq+JXxIILOTP5eNXgtf0ON+z0U1/CwQ
JjQjEAPZctjgYwiODfGN/YTPUbvJWSom4DqlqpsrIa/Z8oAnStukyOMucETpi3Qt
NmB88UHq9ENEd9Qk4qAvLVl4ZZJ+tk8ig9wlQTTVmZK3f1Hjav50kpJ+HAMHS0n5
aQTMySRCDktIKh97sjbLLiAw0pxvMuXYXglF6zdkLO1Wk2dUsxYmM46xC6XzN6vc
h/bfYlxYRX6GZ1f7pavwdA==
`protect END_PROTECTED
