`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9qsTs+nAVkOO/iAy5DVVcgTyv5qkjCsvwgQXuDqYKNTnW5Q9UoHFm+fGzmL5bm2K
3HDhnUyd2dPwM7vorZG8L+aE/m6eO3Xw4nbxiYXdHvHIRzMTEUqq4pgDyKatKNyR
wJDBydexWGQz99PaHvAg91A8k5qHuGn0KR/r1OdGLZVcci53Oqfq4F0nBO9Dl3wH
nGBO5uqUVTfLTvnxpSyzZKlcyBvEqScyV88zedK5EfrdCtf22kJ12DhM15UzFYkD
diu5HmZsngSWiCzwDEDcFxFiBVB6aTpCqRdwD5+bQnf9+uHiodN32nNnKYLcdlry
r8JyVw3H5RoW7rmfBiMPzkPjsK+mj6H+D4k5dbTVYK2DFfEzqLUN3R8K4XMOgQ5U
nkSr9NRGpoYy7Og8ZTXrWyWGqsA7eDDeEXSBGNtwTOAPCIldV9OROrEUnkLop8ev
lpnh9fUwO7b1jRKj5Fqo12u3MY9DBAN0hlg/ChEShu26QhtIYvl2P7RThdVC15LH
bfdeXjlVfvwDvcBa0wxrA91KYPmobp5xbB+GU6VXaa+EvLWSdVVVo+8a2x6vAqpI
HR2xy5GB4zh9VzdopMec8nv8q8RlOoYrrf2y2jvfGv2X0SIdGZMaLazi1VYLr3Dq
/+RukYYV0T4NJc292582o1IW1eF5ncmjlPVrAOrTK+3Qher1N6EXDF5AQ2r0coHc
G6RMEOr0bXvrwCdi5NRaely6iUtyCbrrBr0tYmsoHLmnUZPA7ieDxx8brM3wRajF
5JdOQbt3GVu1herI/022xvl3rBDUP7O/ujkrbdmQCFypIMDbeGQ7LFagdMIx2tzF
8i61NR93gSH3iCnJkhsoCnbUSHzxOqq7yqGW1T1hKp0UOQeKbwfIFP22LKiIXAr+
syQjdp5l/2u0x4o7/mrw9YJ6jCFPZ7CEN04lfdQNiqlQcJdDhKzTuUR9stAfI0WG
hm6dIXd6n1ccfiO3eEMNVHa3kpUk5X6s/mln3/Fw8vrt+dnoOtzYJVDpTK7EDPHt
82xiW/DhV3SmOMG2AZFAchVezAMSv05ZO61uEQDd6bQd5NWjFoOivSEoc3Sfciz3
`protect END_PROTECTED
