`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zw7NL4IV5AVfFkoCOjaFkeHjFlPSlSjLglx4r45+qfGVpOCHUBfaLhiYdr1QudJb
BOgJJQkkgB0HsGF3rr3SeDvRmRahIDpbUUmWOL9R8PeVGmeUsLCa4rGm5qr0kPH1
/tkkbbNtB/qVkf4Kb3uhFsgjPsrwNcptzzv0HDQnBnd6B6apRCSJKtt5pslhUfzB
/Q+quoUagMfCOwQjbPT+644blzz2hc51jGr6IynJm/u1JCp1/hZxS8k3Fd67GeIh
OAqVhg5aCAkDek1GzrkRCvyeBM/vJ0uNI7c1ka7vcVD9LN5tBSIjwAyh4GWZ1KL5
o2/wrk0J3opI5CnagErIaisvom0dxHwoB7qWtQgl9+g4QIzTu/14/hOTjMTHI45i
hJnpaKvBxBA9yo2bk6SLTAji31105yufvhwEah8DuOJxAvU/QV1jLwjaooB7n5zu
Vj7BbwfArVXPAKTicqM+d8t8AYkNxd6f7Fy69MrV2GxVX0tlNzZePYmGOWMUxhSP
`protect END_PROTECTED
