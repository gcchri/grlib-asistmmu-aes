`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6zmJII/4SP6SjwW9ZEJWVey939x+Aavx/BTHNae/6/7WmYWx2tbauUFtGxsvgJw
eAURTQv3sczikdhUy2RC/LYk1qEI4F/DxWNSdQ7aTZRYo254t7c2Z6ot6G+8tRyb
VH96EEiPIcxsFjXjGMZR52DmcyCxQFTtZFvrokiwBLP9IJOXc36PghzJKfL1DY+b
CUJCtN9BbYCECXfsXgnd0OTjdkfcbSrDGVDaCcyGbjQxQ2Px1zvxJa2QfI/DJO6g
4/zkSEz5PsG/kfGLFrnYJIE8c4S84gETBFmghwmy0bMwhgE7X+9TRX9/af4sKsXf
9T1F/NHOmZ77SUhZqWma/2TvkXB/1rgOLwvth6z3Cr5Y2Hw5vhWej6Jpm0Fma5eA
30L+UuZqWKPgktCeMkKpEs1+9gUycoGOMfNVh4Kjm10CYdw7bEMp4yChndtC75Lt
RPHPJUU/mFfw5AjLionPY0BM7QdeVMFq2ekP/Ozml7LFGB7stn6jHBvLc+CmoVi7
aI7c4QgH2r2zjbxxGDy4R7CarHP/19yNMnQ5AdHs54Cvur9D+brAKmQx/01XRjV0
EE8pkO8vH2F9sIYH2CKaJfIFsCEqhmHuxw3nLIBNYWaH6jBRBCCW+ysK3cAaneVE
GF3JHBU4X0mCcBlqdu5DZg==
`protect END_PROTECTED
