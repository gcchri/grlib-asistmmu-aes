`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/YmpCQfY+eTmMZA3hkrYP8cQRPCBB6tZ8VzrzmelUcLptvPfRGVkTaS9h4OIaFK
ZkEC8ycUKe3+7iuSSB5gRjn8LZdrs6bb/X7xml85V+fHKw8D2T3N5C9UMOM1/KiA
0rNMrL6spDgha4s8K2xeBFfhiLQcpxx+G5uDQF3EkVKsvBsGz9Q44p2ta5GP4dBi
OIQ4t6mMWQbr8X2KOiOZqykAsJEtOwzYn5jO2g4eUISX0oF0VNLF0tr3dGWU9lZ8
Mhu85ei8v6CRIU/jGjQ1xqUT5v/sekPbFTFMLTOOTdPcEk5BMXRWviev03Gq9Rd1
qsLs3mWZn9jD05gIP5vwYeYn7lVSUTmhS+z/SyL+/tXrnCchbsfpyNa5XFZQeS7Q
Whtrt1bWh2PZWrqLQHaeNa5RWorYslSRS/+U8lrA/T5tAy0Bzp4ji3oxfSxNrQ1h
Af+7gFjp426INWDm7X/X2ow3RU5hpgRAZOqwt3IaL+Ijluo4cn2hB8I4t11uxgOW
KaP/9lqgvo2WLallWqXd5pHIdUA5gjgChZ0Jev3QXxXjor4rsaKUD5GuM83S16bf
/xNQmAx1fuKxD4NsD8ZzgEu0glYqZsWqW1lYeZiGPuk=
`protect END_PROTECTED
