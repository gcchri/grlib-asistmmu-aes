`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kE9yV/iu/DlNqt3fnzJ+8Hi7CQmyiPN1JVC8pD4ncyfkzK/4UgW6K7+Blz8mrl35
gWqfANedQ4pDzoKFxCr9fwEjCOSvPz8y526kfmyyA7u3udnCqrBjv3UTJNAyqpwX
0dzlxzzaewffD1LwAEAHZD2Qg5P0j4XJBA6SqPbRdDdcUZWoeOoiR8ZkEeP249gB
jNB5HvzMRwunv3n+FB2ltenOwO8TARe1pfBQHMowl481adV+VG4pC26LMY/erklM
SpxKYPJCUokS2nh1GiUPKzXvO0wzOLj755ncE+ey5iECJ4KT2CxyDjD1myc2VO2K
NYRqF/i2fJB+XDs/15orsEq4eW+TvUnIQ0vzPM4fgqbzUQHRq/whbPOfrWtdJ9Nu
iCV38W1clueu/7ur9EZLPCvNi8UPh7m1wiGYKSYREZ1XBHSP8ylbAnYx8b1fo3j3
qQzAsHMODPcAFrhIlxd9BagK7GB26kZ8T3SuAinELgwN7n/BoeKRS+ppZUpmHYg8
mfZDwX6HTJJI9hXcKx80zC6BlM9OVNw2rJwkdbCXSRonao0dyW5RMSJqGMgFAnqv
GAzSGHzJbEpNP5IZBb/2vqtOM5MurtPgPZ3GFuunSV4=
`protect END_PROTECTED
