`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BsD0YbJOrj6BffAzQxb56diJAFbvl/7N3G6Um6R3mHhXWKWUK2ZTZHhf2ZN53nmM
GWSpDPhRK7NnkRtbPq4Tx1gAPbH/8TEgGm0JUtjn7/t3DwdudV1vf9Se3x8y4ice
DX3x95Eaub28mrpEhno6j7za4bHKPcnFZc5g4h2ee99n2/lBtw10KXBhsxGllAQt
2u9ctuyP6UYEYMV7PRiszQE6zPEhAV2KsFnum9T8HhYWiuXU/2LCJpWi4HxpZEe3
UEjc6pGtalhfHg/Yyk+PvWH/CPoKJbHVL50ESKcDq0kcbwvNC+pEak7fMpScFFlw
f9j+u5hP+Pnp8bSymMVAIEUPgx/G9VMPTwqgcIu5OYsWouSgMLTIdSfRsO5ZIHVH
EpHDNbtrZKIMOqbDCRHmD6gHv2niM5y0xAweAnrEkzpcyGEXgz7MQWcRae4ZWjle
AyFn91Hl/QAiN+TOPujbW2duI/2JtNumi1H2ryIZ8oIi1lVgE3T1RvYfZM1zyIMU
dlAGNCqlmXnfviIEoIxh/tL/qJLTkB4zeDOEyqJRcUy+8aIbTHizHE3+VCOqXL5x
TAfNgQ+gGoSVAO0BMl3rfw==
`protect END_PROTECTED
