`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HegnDFFvPAPCnF4abrq+FZLxEC8TGUeccFVpIrSKnPQE3Y5O9wr0abu7bJP9PKnY
HxuLsdlvgWGrK7hxuk7X70siDcrdHDtog1sjr8HtDD4Ugp8AJcLznhEYv7Uwpify
2Kibl1a8Nrbo+G8fkEthlZCL54pAOGaM32CxH4ULOx/QJdvf6Bbfae6tJEdEXfg0
TcG7l25oWJ4Uc2ByYI1AKTJDlf11WhUJOiDR380zAb0k3scle2PAcEOz98MjsosE
A13aTcgUwHZ+8ObLS7YrefO3loFjJUBeoQYiur10vNE6ARwr+X8ZBqD4lQJfFQMQ
MxKsG3uEi2uniLxkKNthFmv0R70MdJ85Xxt9/zJdHVIUwYREl4fIWBwTmDT7l0FB
IdvcS24h5bQaxmnkH5X6PQ==
`protect END_PROTECTED
