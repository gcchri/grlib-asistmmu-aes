`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wupMfsvkTQKkDI1Wya9WgzWaSametaAm7w7tKzsZX0XnecFCsze7dTI/aG8tPTgk
7/NwJw7HRwjMhlr9yU/1ZjVSdkIMJDGnW8WT7r8RP0xVnW6ojlSXvWziKx8cKMyW
DFYwHsgf02oI7DHyS/FYXFJWUaZStKw9FxTIo2OzWCohB+suFavFFMd3U+C3prvZ
+mTFpP1O60y+04Ed3QYzSunAU4JG0tXecOwDgnFntH657zldL1S9qKOqAcCV172j
c9xv2wmMhEdDPtDf/TCn+wSg9NbZV367YI2lj0VcNCBNva2gstUbCyBjy+tDh5yV
rKI4DV4IntAch6Xb3JigiSDW4ibL/A1+7c4AQpq8CxLh52/XyHoL9O68HysQ4Y/s
ucWHRJSLdvv3+Mx4SU8ToBxkj7GpYNA79/Mr6Cq1v9HxC71V/ziijoC9B1x/9rgh
b9DEKybq74TfG7gUIVwi5PAsPAQVJrdelhH5oVlxJXka8m+XLEei47W3ZooFWTv7
IqWVKedpA7NwYeWkJA2r5kyyUxbCgMqgTy3Zuoi33D+sn6KAj1+7FWKlW4X6+V73
C+MmFAg6LVTa8D0E8Njv6E0snEOYlzB8bi5TOL9rN1+4aho1Py30iUubwe0VgygU
a+HwytOsggpNvoLVRF82meAmW7E8omZEhxUtng9U378=
`protect END_PROTECTED
