`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUY3Y4zfZj6Jeo88dRbMXrdPWR8AlxfV8KCu3sk+2Uwv/EYauM2okO5srF+B6X/9
X7czS1f9sONmDdsCdFdvShm2Ni6+CuWhFkDkz1SIUMophpT0ANmbu0W6qSEHZ19i
VfpsmNA80G3ypm7mRPzbuN5X414XfzvFOJLIvsGbjZQXhu8T/p86iy8pW6yqwHnM
ee3ZzefAT73E7xGLOtNGdyRv2CgOOut2pa9iiposeBXGnkL1fBzpx2Wg8C7lse2B
TydOpoO9sXaqQ8GhrW+gojp+NNlJzqsjF4EbHlty6+/VvsrtotlZ7eHSiJpaz1Sa
hoHS9+hUyy5xZuXbbF420kJaWsvKH9ljpH4KzKeACTGjJARefWzhYu5UJNnNaIB4
V0pQEHsIM2tFHGcdQD7dDKNVnAzhtvH5HBPz4rVwWOYkXklQYxRVd2aTVgKtw2nA
DQ2gNGzKnohvtjLJNRtgwN7dse7VDcRqz+sQRAAgwEAvZzrHsI8t24QrBy1g5Enm
6lNROqdMClPQXFXmEMBEGqXWWZNOy6+lbqh76Lh6UoVIdiyITUTM6i7HFCWECFs6
+Ujej2ubQKYxGQX1ViaHNovslaNPy/IKoeniILZ3QVf1MhMFPUiisYzhSP5wTPGj
p/FhZzhQ6Epe1Rhg4n555DPcLj8I8xyVufuAJAVXz4N8uEbjBu3PywVLEQ566zXa
CKzQK9oGRgmWUA3tnMGqgeARwa9W3a2FZ0+ORvZBHbLiosq/cOJMqMVrIYAsW78c
Yp+oa8HGE9w1aksO2qx8QNDGUquMfuN8UltYz9wTX9vQSB5ZJZK5uLixMWiqjljW
a+mBCM5ofOWxi67fWLM6x9Tnjt9peZjuat5A/OihJ6mOkpfqqru8gQ/TcSOnlDNj
vI1gR++TIMsyoByz3RHXsvCcBMsHsHkiMcCKjAB7RTmrVhm3rFQHin48KIb30a5O
`protect END_PROTECTED
