`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xf7V8OSafLPQnQw1NiVdDgdH6M9PyJ6EzzOHhp0qq5YISfCk/xV0XY5lj0pBZrlF
m5vQrdbIXww1bSFJzGy9wQfy6o7Uh2zRskpGYwvObVyLU2xpGf7o9eJx047/54CZ
rLYDOV5Pcvi8gGsV7XuknadVaQhB+01U5rWQt7ulXNOnt27Uy+3Mp+oDueKl8yGY
9DtOrF567dtlIW5PIEy19mUi2Fg0k2kmcYrsDYUtqcRVuhbPGOFxy4ivfmGx7rcd
ekDCa33w39u/qsJq0aeaD8xBL3oKK99N0SL6IR9vHeiy794LiMwZG3GAKGHbAxWE
svd6uoJ2J7m+UvogQu//J+dQ/WQ1+Hje3zt7cCnW1tQpLPp1fd9d6WtBp16qStU2
LZpz/3OpU20I/1N3pKSOVA771iz78ewoB82kG4TGoRatadfjCyF5qRvJzEfMsU23
bLjUwI+duK6BSoKfT/rq6BISl4IraTZnNJMcihwuv1h+riFBlVpSvusi7Xi67RgW
`protect END_PROTECTED
