`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYQM+2dkSMjKVCpzWF41FWMP6Y01cgZA/7aRFZAZmXgFAVSTmwlDingvuwUowb8I
nT4AMHscXKlUQQ80wqzKEm+i/Q8rKlZv2gRE+/oOronROunhcdke7HY+CPjJNxFZ
eeMtuQMMGwD+jzRMQLhBbLN0Xya3HUEkWlpuym/rvoe+LvSj3HBz/cDLg+2NQYYo
MWwA+ojQ2ROkxpPQGwb9SZhwFJ0pTm381ermZukjvkIc58uDTT4WS0X8ItKkk/BE
7FqRVFjvnzy1owdPicWpT6yUEe+BERJfr1RAd+nB37zSwOMKk4fA51hU/pfbesEh
`protect END_PROTECTED
