`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQdtmhPwraCS0sKlVcf+RmfMd8u3T4gFJQ2o5UVRorD+JU4fST2qK8+eqBM2BRPY
fKeBEQFql/wzuU2QuS1+SWHl4Ub/DaHybcr74WQPYb6FDjK5sS877rK7FqaQ638K
3O7xaeMGA4vgppDKiEuxTaaEfvseN0ItYRhmgD6hetdAUiXPgeaOhPAky5pN+q+f
HrwnUjN0aR+o8zAR1A8+DuwP9qEin+HNsW14IsekmvFCcsXvhHwuxXM93MJs7CUY
bG1Xc/AH8xnQzVSzrz5CJvJcIb5uwndoO4TbQhODKz0ptcmF2Fs41jlbt5gwQYmP
RQs1XPTFOpodsTZ6nfQaSu8a0Fj34cbDpiSceTPTdo/dnWf3hoT/i26sWIQDmQXB
B8e4+Gj7vQUjXis6awfipY6IZBWkzrMNZqi6PkkLDmpUMvmD8QzsvzXA6/3LuHof
66/5o8qdIqasMg98EN9cGMTISroumNd0EBZB/4hsnJ4VmBMz2crhOa9BwIsGXMs3
6XEdXlq4U7xtu7UaY9vm5U+Sv+MBctoHYbPSF20PjRGl37PVf9/BjhVgg4UXk1wU
4LtNZd4ga4uqYoSRa/JW28vIeW+JojG/L3WY5GlVbZtBN/wif0I1OFxjGfDEBhwN
jiKXO+Ev8SBqmTUMju35tGoEjyYIfR2YAIhqIeO73U+gOsnd25M/a6Eizw+GVTnC
V2Nbx5OTiGv05aTbDU6fyWxL07P5qFHCfZGtYZ8UVHLko6Ba/o2w/3RJpNpv1xpM
`protect END_PROTECTED
