`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c69TmhypRGNA0UUxUq42nu/z76OncHABcpVwelrMCXk3IrruW6dsE6zqeYEsRldl
pBmlMsQy8VlnJx2otBbgVpPSIIZeqNZnPo6NNmGWazvNCRHa7Q42pwVeO8ck0QVy
K+3S2ATtphH1ZHEh3t9nsWPr8zoj32QnJ+yyZi2fRJt2PWjwdUhJpwbSPDQiee7K
lfmpLkKxdAON+7COuPynxsFCxneL2LHJk4RbBKNgjgdZRL5lKXwvm0f8NLEmVqSl
fXmW0+AspWtH4CAw5ZGnh1KS/jZf/Cjnv3xlMqaeHvpUTYO/i+Pr8Sui25z8RSqs
LWNolzCWVNHf9ud5ZJ74vfof/TcrbV4KVgpAzhRFI9qvJVn0MTyKl4upe061eQq9
KYx1ii44gCguq+nzWpuAr8Ex+UTouD+vVL5rI4OkCiSz8RdKMEjxyeCPMGWw2Co9
osKYAOhJTIfyvOFH44VFGddU5alFAjqD3IsOtomW4IwlEXEzCSWKUzghyBTc25RP
d9fWo8M+dS3vN0qSD/l9nUNDTwCaWBgXAWqUZK0gMcvRbj7mZVecvHetoj72zp1a
yh35EtPzz/SVbi/663YvnoohV7GbuUmrQA8ZFL0w0r8=
`protect END_PROTECTED
