`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eo/9MLIXcCI60W8I7iXKr0t9RujPjhIQFLzcVkFaivUA3LHEZJwV7hEQ3pLze8cK
oxEPUTzmTM4uTAOCtH8pIVRAbt9WmLF8Ruo8Fg2BxTGMO2CHOmZZdj55GBooVnj+
Z/0jsiHEBGmSPwBVM1dgOkWNNRkcWEeGkQ9ra3vIFSENez+hRFhmiL0Ae/rcr326
vlk7d2xGP7hAEnFNyFDKmWtbA4/PzxypWRkF1LazuMXDHwTIRT71EGMBfWUXL75x
+EbDzzisiddvIbdkg6rIP+hwzgMmQpR4ZzpqT1NXSD/U05bK+91WH7ibyOvaVDhl
m4zrdy6iWh3/KY1PwbEGofM8nkroKeNBUBXnkWegCAsYDhnK4w5Ko2qDP29L2SDG
ICAzjzhZLGuXO6O+T+lmVluCGVVnN22oYLStF27oqHZvNgOffdLnXcGaHwqjRF3x
CdEVHIpQusXFpAGSvaTK/uyETaWn81HC003MfJ73NXJ05ZJcCseZrbX7grqTqdy2
7Gvq3A6850O/BZ8lAiCkWN/RICyKbbuB5A6KnVdu4qNyzPFJAii6OGUrdPdERni/
4XikMo+pXcwqA3z+VY7d1E0vlWpXSkULUj7cOZxTFxYSgKWcy4dYtRII/d6iAf0t
p9j9pB1Z4qJPexOUDJPvMVrV720P3gHsI8kcJOeh8EPOFyG2ddDB08hcUyiW+hyE
XTi9E0JQ7Wpnmts30J6ax2A3Xa/B0orRcsmLRpSHwnmd0e2GP4grXk9txgwPByCV
KA9zvVOFg5GhkpuPcDImVvlxzId7m4tNpV4/loxiJxyrt9wByROstDuuqTgFySkp
SMcWo5uBtPRBfQen712xmiq7pT7AXiS/iw0QlWN5VItnfzAS0YevQBgV77c9LMcV
jtZyj0mNOHrSpxcx3dr/J9Mf7/TelRxwuOH7bailyCydWTuSV2tW6+vp5+pglUC/
`protect END_PROTECTED
