`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LIoA0Es1ngHLUYlE9klHdr5P1pVlaYljb7+95pa04BMWDaQp+Uzvq2PMc2NsAe04
pv8erUqGXmKGNNzbqnAwzgWnmxVA/0OWc3sMXKU1La5Uq2V1igTbj5rMbOo1wGKn
Dnry5efNvKMIZ2mb9yW32lqOmfNxZkk29EwJV+tpH1NEJIi1xu3GHFM/Qwww/kCM
s/QgWXc35yqL9hqk9Epe27xFuwOfj0IlZ3UTvDf5Xscz7vCiHn3bDnanYSbTyea+
O9GrfOQ+UsqpGq9JmH9kT8XcPIxzAg4hHWqmjtbaYMYirS7WKJ0Z6glVz/8IF6/O
a0Ls/KwZOXTVx+PIN57zloyqQsv4RRdeDBHroWRtdUag0lcLy3Acb/C4UrtESZ4W
IV6rtLtKImodTbLWpBf0LWQsiWCgXi2H0lUcayOeN4S0+n06pjZcWY5zYHfPg3x7
frFpBRJ7R2Z3f4VpvT2RwwLQ98dKA8yXR/JrhYrjbEGURWP3sLTgsSD910CE/c0T
sEwjAgGEiPDlMxVkW3GZKythUiYEj7RmnpOFMP/qD3TfcmOEoHD4UvVAkVYRhe5M
Q7JVcyaWU440uAuO7j626g/yujwKSMX9twr1dLHbOxx5CLi1yoJ05xkw5mSkijjZ
RnXweJinNimQbtWqfY7WJ+gyPF52n1FS/xAVBlxF0ysr6ESm8CfOKEw7q2QOKy66
kffZ+lYjqzWirVy9FbPJVq605+i2TM+tONNuTkT5xGkRNuTw1c3Br15MPamnEsio
VOBmQl7dhU0cB+TgyUDTSCpb0GnXwPZDyvp+j4ZD+AwfACbkqlEf4OP0xc5Kw61W
igd8R8MwpU+r8HHkqBZBnFWSC8P2mvHoPGf7EoLSUppUV+zvnfVKj8o7tLTje7Xv
lkYvqtd2n+3xDU4h5MOZUJTPIe/VZsEBKwG2aSREloSMELZEjUU2bHdmSI1uvEk5
xHtpIiKg2OOHjIkIyO2OxuwM95zidN+TB+bP3uqT/dgISuAyASzZO3lFf34xSX00
09eMCmUk7QEZVBe7hnNH0HMYgt6Sn0CSyo+OVgOfB8wlLlmQFHHqODrkkkCLPuPu
`protect END_PROTECTED
