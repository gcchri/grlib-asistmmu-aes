`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
awTk5O8MjkUavS19cTcZ90w808ezByzgO27kOH7PtDVeuuOq2uAuV2nTmVTYHRhm
Bckfe+u6IEH6qhqrmdV19i9WgUGH1TIWHdSN0IFXXTIYp2O8pxuVBkFOABk5JYw2
B7Rs+6gIWWJmkvoeVaNfpXBz7dpZY+vRhsIs23dYDO7DRTZ8I2uFjEvAkUdD3OAe
/G+93a8uhwSdZHC0BS+NF/OMrEBLDHqFja6wjFTaIZxSUb46g9iL6hKQozjPN4SB
E5L6YexpXpk+Fb/poDDf6SdoQ2NmSOlHNaXKmm7Y+QxdVw2hSWpJY7GsidybVUyS
BlLFXhkTJiQLpa3a30uBe5E4ouj/C79+TC+pXBaijY8BYee/68TQR9ZdrfZ0RDAP
cQ0PLbYrmzk7nXspucoSeeshcsYdYV2CVULsXxIOOBYQkJX/8rEbrlnv0FtVFXmv
HDrnO1ljI3v9q6Yi0EQwlI5rrBj0WFqN/EtDDbo/XPqXH75+BQVjdPCEV8thNpSe
+XWMYUn6CFNWu4DW2Lm7Om5MrSj5B3wk8kFfCB144UIwSTmUrvjyMR+x/t8qRfjX
fZySWCbkvtYoujokNbHUM5uzk373GiMMnjL2dkzbwzg/l4p5p9DZL3cjw0BaBWgQ
s2fULO+KTMQVoj0e1dIvg45SW5hRAHQgmFIbV5c5t2zm/ETsU1Dz25kmheyR63fl
LdcqR8k68/IiePavRfZ5QOQ+LI2vztpWHzbO090Ho7/YJDtzVXUlz7o5qEPjXODd
8Y8WrvqV751pLqKhgl97/VRtvj6n09Uo1aVA+461cz2Z9HOYd7ZSmLYTUxC8MUV6
gSn2fQMPAcak0COOhWKLhCjfi6klqxm0olKLhOoL1WE0YSHMyFC64wFvdhEMaoe6
D5XE5lRXEN5zMYADnJXNFYEA0QFbHtXiGc1SyQj2qi6+qKBzzb6D9X3R2yJ4Cwd6
yuzzKVDUtZsRdN1VIbf9+QwAR/vLhoQYo8lNjBfYQmmW1qhxAo7f4g+rtoRCCIx7
EP6X4d2V/Gn4XilVH1ROksSuCWs5m+/ZSdg3DnGi91fvTokMNZe9I0tBJMDF+4Gw
sUfno2xQny20NtkJjw95FYj7Udz92arnmLgvKKobOaE4xX3INazC3+HMXh9Q/M7t
znkzgoIQpBgLHzc4BNRTycTlBhme/dlY1nPY9Or6zH5RAUCMo1Ms9Aqa/gO43xVb
4GDtJz4JTASS74pwLpHf4u9n/JkytzE1xPKY4SPThY44II7RbyDL84E4cuJzH3jp
jqChCLt553/3H0EGW3TFIR0g+OUJ/V/6qMAyjNQO3gR0J8zyTR8qKWYRlQ99gB0P
dS8Q7rDhyUd4seSzRjvdS3jIVhG2m2Et+g3pT5IU25rwz7J6rt4WxA2bU3e6nYo4
b6a9kMb0myi5XAKL39X1PlUZilRkjGYcrfbdQ/4y/nTpq61Lg6f8SrelwGYTrOhf
5iFOpYn+Ke1D7bymYgOVvEL25XAzWRzXMkJr7ZKNa8Cxn2/Pjpf5EPdkNKSamhRA
hJNMdybtcfgahwzJgeGb+HlH/B4NhaoDi+ZlXvHeTyWGh2kUkWDP1p9Pl9pSlL02
OYTUjtoIJxABDCDlF83JK5sR2USn/PB367AJV4Jyo5ALYI+aVUFWYi6gAELkecwK
oxjZDFXWGW4SY98+fQr8evQVi3+0k/QmsRSSxxIy+cVZJn/T3KtN+PT2MDkFG8fX
IOIElQUenaEgCThroPXmTQjmXsSsJFffy8B0R7eY3M/aQmvKUgfhN7009NWt8ofu
r1JZ1jQX2p79QpPntcHot7e8AcATgqBhwscoVrxs2d6FmLlA2EGwMRmZYgA7SH2P
/uBbnmdBvAny7IXYxBY6ftB7+KJTwDpSxPgisqZGPv/Rn9bcwXhZb0tgH7Iaabnn
Z5epuat9SDTy7nJJptkyzgrT10OFFiJfIZO7MFxg7qpi54zmcpIW1xEK/YhJscTQ
QfXjxaD2A1eGdxyjQfecv+yWBkOZO5ZJp6m3Q5ME+mRoCK3vsMC3jcAieuJrm/XU
v4SoWXGIe/N1SVQl+E/okdRMwwPjRmTwS1JGxaW6SFoROfUI3xUsInuuGiMzxsxb
EXI9JsRUT66UhX6NtI78a5FUPi95WLA/zU8SmmPQquE2pWc10JPUo/0i7qN6YeU0
oVQ2lnu7tgbL8TqL/4DfYdMyh5NOREWfYl60vF5tEaFwmLOI+49NzJWAxu6qJj6S
r5U/b1d1ov2LnlHaddn5qAB98CWM0Fz5Z5ggQIa7gKerixx8UoKtqicwgJJGwjOX
e+ErokquQjOiJkQPbUVbIu2czmZHQgS77aZBNXcI+O2Ryjt2rxv8lQhvjF0yMV/9
Sgex7/qbDFTg5hNwMCCDzkQJ/a9Cts1PPsd1ZLppgUNPnQnk3rb5I02Vm75jATZ+
pf/dE4SHbvOpSrTPgdnraFOR/LIsPZxTMZoKMX+9px+jWGcVT1rbAOY2FFabeiNv
Hwd7kmQ9siJNmRexvcHAP6EFfLg+zNs5R6zVvjsjn+L2vxQSBrR1lujOX0cEROlv
ZAy7WczyYa9VG9W88mJRuQWHBR64BM3gJfqW8/8KugjlRMIJHoqfYd54cN6ByjYs
EVmw+HUW8dAzR0HQp91S576qdopkXTIrwObuLAaTg3Pwv29WP7rOeYh6P1x9esjA
E5MIsTaih+MLOFqjDNupDW6Hol5zgAkAwLbq+NmrdAJqevTzpAAM06ExZi6YETIv
7K47sMQ/jzQj4nqxWJiIb0sWGyurh5Zx2/Dy51SqLwVXt2+2Xvc5pyasJapN6sfL
hcvdO7F7wOf29YPytinyS4weRbQF0aCUC00RIMcFuGsAMT01FrOMvN/q7MC03htS
wBUuYkRqZELSsjV81x0Xd/iiQp8HwY986dNdobJwrB+JUex8yP0Txks0ndDmDBjZ
LW4eMMbq/TcQEO5tCqaLPmbm3OZv7exsRGQDFClxO9khhqkS4/9AurLd3IfkoQEK
H0+QFU3qRcKIsL1kGxQqb1jns4DHie6t2g+9NwtzjqLq3s1XmSX3Pr99tBiSIp5d
NBU0Xa48Ha97MBAFgQn+DOun1AVBfZrgnpInyOzP9urfxUpGEm8ExAjSfcbP6Zp6
6QvU3osvEsbLfcmEG5uZxsli1p7FykL0KhujmdsdzSkrwOgg6w7s0qnj4MoXM+yT
ggvzR9bulBT81LRa8VClSQtEAUZxazHjqqkU7JjUOgE2wcAQytw1FAw+sThbBWeP
U5BpRBDw4tRVVSMEaVweV+z2A1aVDxOfvXDkv8GNyG20MxG6iMI8v/eKN75TSr99
oKeieG6Pg3068xC3UivMcGOmr1IN5TKHX5a6lcJeHJltsoPqUdc3gJaJfjF4hCsN
GCSCHmHZ8C0m0fg/55nXl8yQcnaIJcVZtZIrtSg6GpOLc/qOSlMHWc1DakgS5l25
0ThO0jAGxYd07Q29UgkoGHp/oW1isC6Mb19yAGS7bslz1J0Rmk2eKZ3iC4WIkNJG
ZA4i0SnrxMq49oFVbH9y/5mP/UHEajlye6f3PQwVZPmVhu4apm3ved1hRZxcobG4
g3htGykryHvYlipnb7qfDGYpOHzVcHW8VpSy0Vb23ZzU8IQaFkXfdtuu8aY5YoI6
Y8qBcWIB/cxaMFIYPnjRgzVWmCHGw2DwxYH+3tEuXB44YUdz9qUzkGpq21EQmhdB
YzPoaEZFs9cEbFeMyuA4oMjKkwex64rq6Q39ERVcX4xlTEmt/w91Nm1kWBEXj2Xj
gFsGprNCvB/J85pJ+8LnuIjvfj2tkX8u9BjQse0dlDs0UiLuKmNemIfBBn/JepSS
/sahqN914Z2csTljXAIJmnuAh7Tx1uURt6tpZpy/FqoI/1uPS+vrFbW/Y2NZKBXt
lanv04jaFUlE6EU7KUSZg7hyar6q2iQvD0DfZsc2PySMVd+/DlFJu/9vs2uTZHG/
pEtCcdUeBftrSs8BgCw/kO9TE/T6B4Go9kLCElI8JypLciIgcHu3vL2Uk8s8Terz
MdUo2iRVUDI5mkMoCxF3DviD4byt1jH1if7sv+4R4Tl1sgL4RWvZWIyibtdSbnoK
VBngxLqao73yUiuQXvk/AEm/002jKOUZH9+qgqt05g1Ss5XhQP12M3dcwLh7I3t3
zKxTtlF0rokpAzs+a3Py1IcVmAWoVXLPubPwKL2jg1tf4hgca9KlhcYMUkke66P1
0cbDW12afRugd7MmHPot57vi5yV/A2WEhon+j1xs8Ics47yVuDpyQU+vd51hhcHi
qPzWgGEmyo+JPwIQNmTDs7338z+ZD/aXU4WkNj7N1R5SqbRzhfQFR+V8oY5Kgqo4
C3hBOtTPP4U5aVvdm/OiS85t6d8MoRh5Ks7zHWp8/AiUQOylhZzhJTUp1KnBB7II
gcb6anpTOXAgXohMldw12FHMrHsi0lO0vZ9he/5hWfvHe+x4jSCx/aK0wNFOg6H4
Rn7qEbOCpGewpUa5/evj+GFoGnP4FDdo4Wl1jI7svds0Y86iui9t5GUqC68i9Zdu
03nhrtWNmwa9lLmZlkXUl7WfPKZPqAJvWBF2AFhnfYSNxabv61YDK4oZKeZWRJtU
Sd3DE5uvee6gDOBNs5MolgkwQOI43z0ylXlmgPZuLDiB3typB+nyBgMyd4PZbVFl
bqYp/+vpwesTKtPvaaROl0wa+lphibA/sE+38v9B2UDhtoum94IyXRzvAsBNHikR
QsRxfVHyB6IrR8Yd2+txJrTqC9SjtJiBhawgZRDf7cwjQmweLs3ToiupX/Dq/i7C
TPox2crQX23zgv2BjVe1G6R4DU9WXO7skX9BFLq7hl5yJBh7M3BnLabI2/3pX851
P2xYpe0+7pfb5hIz2Gc8j9Cj4kMvQxKCvNB9w8hfGI+xalqfqKD0kf9S6DTCVOr4
yKKbpnQJ6AbUPFoytzQCq1IjStZLmYZFW7J+HtlYaGuE437eZGdYUA5NuPEimiBL
gyAMMDX9Nr39F3P2Xi6EZT4grLik8lOhwogbO4LxWw8R4iKVnpfXWjL7iWz2z/UN
/pIUXoDz5elUX8+CWHGtKkSL5teF/w18dTLJeiYqssD/F5/QxtKSyNP+cLvEnQFB
zHb2WCwXXFBbgyVwVjCYMZom05q2JmDL9FPX2jGeUCM7AO1SnRBapHcXIX3Kyvgx
keeBQ6G7103e4GCbiDkzf94otIqFeWX2w40rSiotkZrJ/8utBZNTRohP6ROOjHSP
jc/Erzsc0V22nFGxkUuGZ2Z1BlbWLxA1LtPUd84gpnmH1ctXfHVFBz5tWYbDC8lo
lMe3bHArhc90YITAVZL2hlpT2/eTRR011yoZSaCPedHd4/9FGl6LoCw6gsba7+OY
ATFiYocwJnYUANiik1QOALhVJYpdeDjETFwL110aCL3Mxi+KeitVy/8Zg++8vcVQ
8fYHHRO2xwCgsyhH/NCQbiFEsvb6pnF+4Z5GIJPd8qhtgY2e0DrTyAo3DdiwpJuC
zY5jib8ZOWyifHrpwzzVJPlWD8u8CPbiuh43p6qcBV/tJ8m3pWKdVSvmDkVSwsDG
sBCZvCIbFgtZDvtWgKHo3qKytV62l2NSwLiuvWnRQ7NcIiBpTzkhMKGjxzRlL30N
UIa3Hz1YpKnCYgy7oOICgN/Kl1Nb5m/j3upAbfrFU0OG1Q5TR5ZhK+7hVilESesc
8frFknGY8LcxO6LHaV+ME0spnXCrUqc+xEuLwHbiBRf97t69EgxgBbJt1dZHoedc
YE/TMhChK82T/41C65khxpipuewXSlnXAWHXYipqF/8lFZbrmd2AzyyJFxUstSGJ
IpOgsJGOdT03r+wAaT1ny7UhLQq6KZkQVlyKXoctP2eWojzEojx9tckXzfM8p+Xq
Cgqg9KWSdcekenj+ZXi5hrePcCg+CH6e2biMu9K5Fbvuy0iH/pMikZlc1ywfoJgk
eatnHNdY7c8ympRMjthxm9LkdYkYhSafgQk2ynig05oV4vs/QYiqaBIbJ/xkbiMh
4Fo0lGN4Eb2n6uIUlt5CtfAY56w+vTmrupxZg02HLdA3lLRbgLxihDLD87G576eH
KG4p4bWWoqWOtRrLc44FAKqSOrUgsaDARUuhiEdRp1OfDjyV6aivvWCX/iiFNJNb
2VhSrrLosR4DRhPwCqrF+dHoApfo1subTZ/HACVpXun3tptheWwu6mzZpF8lyF1O
rXd6fABKQ6dzqnaTy1xZONfP4XPBaZ++aG8tpGxMh/25p4T7UwJIsUx8JlwzHB6y
uc/KD4ga5Gw2+cN//uB8RpB78d6nOW9foe2Nw72rOyuq5ok1KXOZ6HFQiv3Et3fE
qTOl/bRSLaNchRFzZ34IFzGHgm+32/ufsEHE/XUXvMTI0JE25CVAdS8idT27RMSd
KTwAg+nYMWNUY6bABoQbCASZf3F/8fDVnsbxIGn6yUfIDwENzCNZKXE142hVZf5Z
Mu5lvsil+yh7ySRYDoeU4rNRFsWmo2dACw0tQZtm3aEBwvxnvTKnZZA2d4w8ncWp
Eu/8ipz+dvJBcOcH7aAuZMUpBW7EpIjY6XaUbpF20zQP0ewriwyPZlvLQG9EbXLc
NU9VophaHKoWku7r1c7AcZdFQLJvTA0/xcUqZTCxGvwSkqdrPdZQ7oX5EITjx9AB
fYwgBMCP6k+3wodjd2tfYGUoEctfNUC/oUCwWnLPWp9QXvv6DC6or/9vWQXeVA9h
+SG1GXPUD/dy55v0oc+ujWhVgi1GjNLflrqr3Ed/xj+VBv80pyGD1mC6f0KMMsYi
YW6y4fKY0ssPNIZ6NUIMEHwDtfD/UpX8v0O8uRxvmgubSI7XNMNGvkQw7Gk5qStk
rle/0GBBAJoq/+ig8O8bdPZsMT0YmTlgHyvJScA55vNHx5ZrjaASuaYhtZz3w7sx
keFv0HIbp1liwUfK9qJKin8qfLYEJcPjQG8QgLpeKQCl/0teoeSthwyDf5RROqCh
hUfJo+Qq4qaLlqOp50bdvMB7rBGtW8pJsXWArq8l6jOVJ4Pu2IUksVDY4xGoyIkx
jv7Wc17rwub7wB8ybqFIJ0z+5GUM6fNV4IvUqZVi7fB902LHgcHOvDiJObsvPMje
JGAhTDe4C/63f9+PE+h7vmme3kKwCaRcOyc8iB6TJ/UR0yjIS69hPbOTgfxWdazR
7lozy6IP8GRKMU0vV4dIehGtt/iQynS50yVUVyZpo53qSgcBBTAuPT0rEAuTJWBu
LXt78L/SdfdYHUId7c2uvpGPEuFTfdDh8bG0dYdkIhgJC+h8pT0HSg0dWJPMzjzU
Kclisw0NirpAg7+4HCsJv/Wmay2fFqbZXm7y9VYpoYkTfT66DYg3hLG16eo/pNFc
lBOfwJDmvLRnLdMz/Sryd+gHkVNdyXNH4DuuLI/GIAJ6LY83HDrR0ITrKwSQ2fjA
/t2DKg/IxLLvh/5162E7IZ0QLMXfFaQEnjPN28ceR6lqDmcueLzR7OFWiLNTVoRN
zLT/eMPo/knfwhcE2W1fvTVXR6tm9EehdVaqQ9OwBgQcKcPCKusltfty4oCY97tf
7J1BWlnHcBR2kTQDhPQfCj0mFTHfMDDBmuz5d0vlnF/8Wm8LoOfgohDOTv4FVCMW
RLGDWr7w+o6LTIJwlbsA3ae9DpPqrpWEtbVzNshBK04z5AiKGRaypAbX+Wg8omPG
RX9SiAhXdQZPW7nVZd88a+Ik/lSoy8qEwTKaJe/LeS4xCbN1dWE7cUdg5+97pKK+
muriZhl4g+OkxKPAYnT+b+klU05KMLQNHQwBwUWi3/v0jBYFrdEfEmsui3ka8JNs
RLqz+pyBe3SLOfbFHNDnNDDTPiCy6TrYcCpWDBA7zqIbQcxANIT3Yhs4SqWhbkDW
rodnxmg0Ot4/UpL6IL7Y6/oVmZNxK52zoQP5o6NZeHNSgOSRuI9W/MbHC+b/aHa/
AGzakW7ySMckL54653IcqyoMMWbyQ+3F81bm5wigqsx+F6KayVFBT4Ju7Q0jYZbB
/CTtGfUcwiUTynIlqx23pqJm3qWAOT6BdYsb3++t173YGZ4vK5NN8irI43K79aFv
DXYKK9PpmiL/yAqDQVjek7ZpRxEsiFJ2YF94+Sujudnr1l0/V/4653i/gAeRGpd9
EJhnx59gujsv+HPOWQMfZ3k5SE8/F8VBLI08T4SNo6KKt+ejMnGwR5zx4JVOa4HD
1uWFxnq0EiUVcUwDR7EYrm5b7cnLPu21kb2qttYnY1OtQ9dYEJlW2byDD7UigxiC
7Spl+JlzjnKE7/oO5noDsq2WSq1sQfIgLfbuFFoQIZZ3Zrh/41BIhgj49o4dRtKo
NduuJUo90ECZEOWZw4setWk/DLZbVfvQeWLXSMm+bRgUA1fvnEZxks1BV2XQp+ZR
wh8wgtSMwbYYkzvezYps/uxGFfbvQYi1HQp2V+aKI9f7FBbAABT8wb/4noCuUgnB
SkZ2snml/iM6oEM0FPRzNtQoVINcWnqRW3kUw1gOIVz1VOjesbwEA7BvOwNg4vqo
g9UFfIhwBKeEZhh+I1j6vzicROe5Uamk1TH1Ri9krilSxDw8jczXY3tvwBRxVRdG
xPR/6KlqyoS7o5wCvohMMvAKd2sN4m2LBnTp2ncytyzGyhLoWXgmtBXwLrfo85MI
VWfZw8xzFQXQh2Y0L8bqpH0k2LZmmVq5EgyXQmSLoOYRQL/zkC6u4dA+gF+QOpiE
sLOKO4xzjhF9tedWxnc80lK4N2rPs8znXZtcfRppWyG2DhmeDCiNzBpLwuJP91hq
4nfFUbADT29xWi5+O1yOHKKKdpqJfq+zbiz9DuancJD0babtkssRzh+Gky+CTGDc
Q7PXmoiavt4RYbkw0192et2SbsIHQPGMeBFmrrQfMvliYRvZ1XbitYn8pRRrim+4
lYV6aaT7b1Y3AbtAxPXeeLrUaqhAYi2FHukwdJE/Ksccwrz/qLYqPWatMh9rwQ3R
qVfwRaKeEpp848nm2D5kj42pLO3QVeyYHcJN62n6nsVIGVkbHtSmjofp/aZY1sBN
qlJLQ2cCWCx+5jml0SNZPxKFNIlfbzKLrmPgwje7xh6nLkDDijAQgSRuT8frF77u
BY31dqsv4SOdH2d10qJu+dz5KMv1BW23qlbIzYaCVOTJFrQwMux8aiyBdG4h102Q
1Q5ZlhVsYrVVpMIUXOC1Zmt0GzpJD79QcN9bzSQt09gkapFeekNC9uUFxQfLPxq5
mi3Tb8ImpLx6RjmnAlTz6iHf7RXvm+06sJQdNctHctCmFFhP4H0WLPh4FuUOSUo7
7s+ReBQv+YgTVxTjIPPvAMGRUdKycvUFH8GGiVkouYz93PoOkFXNn0CSg2f1pSzN
zfQgkcP7TfWgwEWdN6GYrAj+UJJs84OMNqo8owtD/SBCG7/vI8TR+AwPwhRGxyOu
dHay2X6AKkgB+PimqZCZHYe2hxmQTj258BsOFhmMZ5mO7pf0p+GtXw07a1Tc0YBp
hyVItUgHzzQs4CKnzTPLZVtaxkkemONMMpVcN2Z1TG8KlUFvUE+UvPct3AbQC7Nh
Q2Y+7LeFvJMiAdY4FjTBLPTl8V+MrH7et6WcRhNkKPo1gYj5+XRLlM7/pcy/QRAs
slwXKDvEhLdVmTPM3OFP8NGTB1m2Nwln2TRP+H2qjG2wzum5iz0OI4Wl6HwILwgF
6o1rRfexyvW4wNqBByLSpTFyX6Q9Hn7EiTtPthHvv3+Dd6tMgAvAtGvoq+IjMgST
flesLKB4ziKz5g2uenS8/zJcMFS+8qGOJ+IMePvQYbskHyLy7odV5TMGolQi/LQl
pm94ipA1x2HWp4ppBqe5bB1err4q1fMW0t0Mj8zqxAg1RVx2dlRDe143CGjev2MU
TrBEjoORmFvnHCiPjV3kdXHs+FfOEKtydyk4UCBN6aPavaK2wzuPm5hem/cq0Zby
dEbw08SoaS4r62zq1GmSQG74iDkXI9u+E29HuMNvLafL231Kqro0a3c5Q60NFkhE
U5gaIHrMVQ8KbGYr4mnKptQOxF8fIhjM1duDGkrkFS20Et7RJwZ/MzqDRnjKPcRt
/Vqgv3ml8xzCN3TOqnkSXCeMjm5b4IsS+sw/hjSNpLbFLvNKbM+vpMdxnQAwbZhK
tUpcc5kyPSqN7OVzQyf1CeqjheX8kvypIrrc8YAKPP2CxyxppLyGnq6VQRVkhEmB
5B1CBd/JCzecmk+EsO3OtMNMj9slRXcdzpq0R5l448zlFW7coYhdcuaz+LrDQkii
MgCO3JKb0Mdzma1PdvN9a6hqB5+5DeCTbagu0eWtgK8XWEErZJi7mLv/d5CqcdWZ
NGtAmjbHLZ6eN+yOHCIUPyrLdi50DwXlhhNPlzLuieen91fPdNJdEE+gMigFNPbY
JqkgTZmKc+JN4p2+aJHWEx68yqz6xir0eRW6l11dDitoNrddJ5bWHnTNPP3qSG0m
mo1HuAmJBxR9/5wUAZxPD5SOpcEqLdR+I68dGSgh9B/1y6oiXodksNbtm2VsB7nk
8yCQ/UYFl0Lg5Nhd90IiJQRAwgBOA9CLBb8PuKqpdUG7WP4QeNnzx42ISjuKGn12
VHvJhWwQi6GkrGwHZkSQuvj1bhAIH1J8yeNhanBSG3mKDEikkT5v9ZzhDowaAU5s
Kwdmdq/a38K4KUHKbqVlVjP9cbq5r/tHlwm4L+amFqL2NWQUp5AOn9YLffuxPtwS
4Yxse6uTcdBJonVl6mKnP/9HU+wAomfi9SVxvrJm085Fr/ZlMqTWYCIcuzNvYwId
aKsxAYTvJCXCM4v6wprlT3IgHKct6E5XZth32sM4OEZOBqPl7aw8cQdYj9dnn3UO
U7zZ72RJbGKRGzv3AA4dxUk1kpQ0aUpB+gDRmXi3CJtvcKI1WshZd9N4T0BpabYG
F5vfvuGaD3LlaZaEH2niU6vf/XNc4HvxivHfK+iAERvLNmnACRnQyJZgpi/sP8dZ
G1Huh8ko0REdpCFNRsKBXyfj6Yq4bpiTK+6hx5csld7kj0TT391b2Y+967LBjpzG
mC9T1b8N2hKgyz6D90xZlaA6dzbAnv5hwlcpnpIoUZLUWrYSB0dztlWp11otMlRE
kY+aQcXUxvs9//T774w2qmPdt49qo/m5S5XbPKmq4gHZm3ejLa5vSWnAD82jvkWt
tkpFV2T3NSIZpbI6Kzq/tIRgpLHxveGIq9JnF6pFy1z8nioEDjXxmYA1os3vScOI
ZS3W1OM4dQUHIsahgnlA7GKSXZvNRYTpDBhRSPEka8tv86QmRbfWPnyFKSXqtsxl
ANgxPHMQ48PyCco8dSztRUVzQkI9ibZ4cieK/mOhrNVA/ySz8NcxPDWPRbpRyrOL
FrKzwyeiyGfgVPiK91AVgBxbndRRHCUo6rCwSx72JCSuS+7vlEe+knLZDgIHXpcB
FKewAeXTsvruj/KcBLSSzOeU8Jdl1NinIUs3VVFJLY/8MA4Yni2GE9jROgGJ1aAJ
5p2VfIMN2PM5NUcnzIWaEmdjq7ErfGy+1apDWhIJYS9n/YfNdns5jxAXBnLsa4DK
nCwjSLiHmiRI335iC0HI1v+95vWQkYQWfo04LnSmObCqd5tKaZdx2RI8DWswbDGJ
+yxbhSEyscjaQ+Jb8pSR6dq7HrMf7xytzmRebkjFDIPnhgHhC10O1VIZrss0Wqxo
C3RR90TBDlqF9Mf/Woxy82H1fYQw1gLPhnUpJ4Ddl/TVfxbgv+Ah6y9vAC6SVj2x
hsO/b4UdYWf9kxqYltaiHklVCSwDqc8LGQ41Jsw/WKicy64Dz5IS7dEjG9WEJaDn
MghTElEWcek5D4K7DtiC+e4TWmqZ3a7rvOvdi6JfDgM9TC9Wrd3ZtFa5Vbt89LAn
2HZoIwHro3YYkuNlM2Im1mdcZdAYepbB7afyDKj3+C7dNqyNgIb7wMHBjCo4H1NA
0fe757nfG2CS9mn0BNJl6388kZ8Ed+wqCEEngINrH++mUCgBjq5N56E0Il7FCdqv
jyRXNE/MPnv79uYiu1Gv+9QEgJHwgoVpOtBANWmH7D2KtN0C1KRpPkhV+e2GANda
R1NL2OWFmJcVL75V9dbMZsQ0QpUMUXZ7X+4bb002i+Sug0qHEu9U6NYgdqGq12gX
K7GQYUfa0auLxVs93TrSiXswZAjdtwijqVgwqLVnoIERUQ1b1yDM9jGOrE+tQVv2
7Gk/loSg+mNueQc8zhecBLVlc0KNehpg3H3zcgHY0JBaJ6v1QXCivElhJ0L1sYsd
xzo+zz2O+WNX5Q2X+OgJnG7fCO2rVndTwpcaRiO4loCqkC24VuIwYQbxM7xnLQ3w
fnExZEWUO5wpY1TmUM1t+OTzEXHdBhFrzkW0nfjjMKIg8SO9aTC/JKGzjUaPjxAq
/GVWPsrGvBZTWc3Wo8y2ANwo1diF90s5jlkvGsDm/tLd4MPdVVctSvyHhZIJHJw/
N1y9N3FhffajqkC/GWOQrqSlQDSPi7y0SNPEEWyvH6cZoxPZOt3sbFkQMX38nIMt
N/TWUFhTn5MUmXtg6mLMQwKORMja+mc87mXqnRpHvLqHj3Ac1fGQV1IRIczJQaAZ
lazYwxt1ttiSQPv01VZ/XoMfpOjF2kQPU/kqaLsCtiILxRuYGBxW2RiVmO5Py2vo
iFnkZ4dndCglLQyWwgHsvs70pk40ECbef6Zzt7iga4ZxztanAuU6b+1r0DtNenUW
4SgdwG6b0GVwUkE1LJToHC+QAnvjkECq+XZZMPFifM49FD7ShcBd/yNlEcZd6k/y
yvcg4jpwO1VhUR3eEUVLQFYOp3LZCtxXg65keieQakgDuPYt4qY+JbYzy8DSJDFw
DDUw6EOZSJUdlB88P/vUeqk4vMByi+lVZA3K0qcXoQaj4Hnmvh9kvGaQzdmnVuQ/
rtd5CT1cxJm+9bP8BUeCKnsDKz27i+CZZv1VbOmhKcawbBmh+AToP4j7CkO3bIDJ
+MBc1Ksmp0gT1u9dduViCr00NBzPOz0p2HWjPeHwuZtR9GCfI525iqBIUdX+re4P
kLHzmhoZSmeVoYKjtDJ5Bz5Vev3iFqrzPngMdVFOY2zrmPOoxj10G8yZs2vOxL1L
mDVwbZctm+RnLKcGzXbiXsgz4wf5PTfpN0qurZJP6lMHEihNJ61qJrIzhwvsbwaq
yzxvd/GRj/873WJUkaoVZ7uJosv92fBsTYpMAwUH4PSDu6lMQqrbB5+UMyScWJdM
/jSy029H8kr2VlO6E4g76YxIx+RIOcMyVthHpvooyl1ZZwX7QWo1qAFppqZeYT/S
JbFCSflWuzMvZm28snvXphjhkRlsltzTAaTJmmM5fZSeYryk7XwA+FcvTbqGrn+N
Xgbe0W087ZWCxnrXnNeowOoHRCjk4GosV73HqTrB7+L23oIMge/g55JfJzl8bJ2O
pZkBv0jSZO6c5j0JCo+agY9NduT8XG5E1dVKGo6Waz5be8u8Ld+LdwgsuGwGvV9M
ckTrXNdaurktj5T75gn9P6hX/+5W74Md+Tcizwhl2JT1QeVrdKKyMv9ilesfHOpe
kGYRX9f/KRA54sOOjvt9cn3y/HIgLdIUhFunCcXVopCVENktcByqP2RRTwIU08tw
tAttA2rEvRdtdQusaXIQoGxZlSe+SzF6JITsQDjmzbrGSMRHtGqbsM5qHzPhB8sZ
oFTMU3HfO64Q01++10lHxtm7YiMv4cPBWN/+eGvwTUehElW3BfTXSVCecPFi7BM8
qjnC4iWMS5VoI65N7zhDyNB+Yblif93Itzf0jNU3rAyPDHHWjEWxifugZ2L07Tkd
T6PLAWQeQj3rr6eYblkgIOPTmn1vxpu7Qk+uNjgMOr24hKJ1cLqPczr9nUDcjVY8
v/tvTYZ5/SW4ePz0FYROOYsb+vC3d2+EST49P2wnZWnzwl9bp/zQVMcK91HPPXkY
GWnI2aFrsp3rkV5RGTk0z4ynCiPINCX6uDk9Bxm0VofV7NLrxHoQQsnD2S4tv2fu
tI8y+ASm87HLuoyVSVHPIGd8fM6YeFtwzAPOhPlW6Zv88lQjdcc9uT7ct17AXA0f
L7rrSkfJCIb33EQqvEnoDjyAWYnrD4v6IvYGC3+dgDjRycPJxKhaqJ/hn8AL/bOK
uTPkOHBQPv8OwHeGUOAVhB9OheZAYnDiT6SN/Zsq0uqqWguNNoRnXJEeizbTilKe
CsocGpyvaC0h+4OeToNPgnaBn4FW6sWPpQZ9eCcPzEanwMSsfaJ8nVQUtxFNtVBg
okO8Hdh7EnGAc1ZG1jlZFinr1NEb6dGt3zgdKHpl0+5rDB+g/uVnDnnQgyeBTMYL
44yMJIQvlDZutqPo/q3lOwFADisp8YZXSZD326ztquomQyCilAg7+ijmmqVMJdvn
kOwJnSIMT5K6CcPgpgvKUT1+TviPCzuz3ehGpF+9cdH+ZWlnTaB70qCh+7605Te7
hnSIfRIjsYHPvYBJpKU3+UC62wXjYptdQL0TsWdeJYGYuObjBc9ImAYT3TesyQE8
LP99GcemA9ialKQwDFDqKw0QTYSaV5eegM+N5DG1HqWMtyGSTq104SrmXe8hkdtY
L8QY9zUOGy4fbERuggFcn+lO9Kydvo6Mn9RHF2Yj/OGS/OMU/3JMPi59VNv3VBXK
PwiSiwiOTiMkX7IW58vCUzhmuad8fyf8Bv1szkWIpnMe5jRB0zqiMqjvCPvjyUVL
gwKT8IyLXEl6HEM/24WBLAYrDFOH2KwPKSaRbV1eRYp9Sigd8Dr/ryrbxT30Bmuf
oeXGHaUty9Rio/Q9QALcrWgpHGupwX5RHQfAtfDyjJ1PyX9DZhXRVQyAlqpUX89N
qMLoHpqXrXTO7PfLCXl9o/LFGXKghi3j1Tp8uVIfer54ZqEY1qN4lilKEBIXFVD9
9/tgz3c/bDGINRGULUPNikn3an/P+Wn20yno9RwKlz3AZUQemBU960Xk8ul80vTy
vtKVifUQ1aPfQi6egzobOVdPENGWl8Vsezch07dC68OXFnl1nLfzv2CElzWlWrfW
bZTo3FD0ATTheBnsvodwTm9HimnnyBEssJM+PLKBrerxBe7dVEznGFHL/ZJ1IfGr
SUhSPuRYmrp9gAhsf68XBvMTu9ANXv5ABnGR2gfCGwvKKwqOJWGM0/pOYB20GxPj
NAynOeuQIBaTcjHlnvKnypDHv4uflRdo76dtAkV0nAl03dZn4s8GGafEiR0JcNck
buF8nbfwDvu2K76k6YshXoiph/veMGU9U0viuAt8BXMb4M6frmkWeD5Ad7VdC/Bu
3mSzf079BVLpJDgciFCf6NxCsqyrheCowgU9p1cy/CsLv3U9lfwQ4b3MSU07/FXm
CoDoA8cTyrriqRms0pUeeFZsneJbGbalHLhDSGO83r9i+v+kj3ksNEGD7Qi31uhH
hrjZ27H12HnGNv/pLis5nQz//HX/TSYvent66gwj6gcyfhJ4qh/07hSRnPw8neMV
3USzXXlULPpRG1LcH7C0J5yV86DoI6LpDC5zYZ/dnztUCXp0STPHks87+sTPXV1m
8QREWnfAMlKJt/U8+9zdrliCUcJVEUVsNJqkkFx5jbvbizUa4c9sCmEvKPKzzDtZ
bX3HeHo4FHLPTs5PdUqyfdwYkOKfKMQyXOzjfk5uOdPIGL4aQ9EKaZ1gluXETCiU
j9Rdx0iRBy/uOPoSqGB7DLVSZmv9qLDlj2QBcW0pGhgDcWV8eqhyt9SbjRsXdfV/
9fLih1HtaPDjRFjFoV84JXJt94peS5JqG3ELuLOyaMWg8efoFM44SoX8d8GXk+xA
dMLMzs1enfcmnJGXwmSTNE3TXMs6EvR+masDm8XTpFXXDwZMHa/u2iwvki4ckdZt
5CV35FpAW/xPabtMiMmdpbPHvNDJGc42ZGvemnuJZXE7kHNveXUX5LY6PpqvEM10
AQ2evmBIJ+0Cg4+Rtv3X5/llsUnBTROSml8vPoarzSafKjhqhwwTWfm7Vg+UKaeU
HA/9sEva7Fo7M+mbE5xLzCw6Bm/WoZSba9dP21RELOAJ+XVhflDGWuKepd/f8wcV
K3g00POZcB/b4WALgF0ocAnSbPDjS9STdFzoaLwLz9OMS5BebiVwM4FAK1P2EgGN
WkTTFuc/nlfw6kt2JLC2tfbxcghWlRraQYQ+ZRmNzhgslFDRSs8gaUqG1Wptu+Ov
ed3cPkAmfMyMxqtF+Bs4y9XEVpkNThXTguEvJU3LIvCuhtTGhMEq0e02y1GVPLQl
YsJqqBiSwbLJwAjCZwKQun4ljUJHAN+HcX8f90pHK4qvax+bpRIvbgkmVpYmbqEs
SFviZTg3tD1nKBOK6Dt0JZRVRSAe8oH98T5SBFAGkWJwZ8fw6cF/1dkdC1FawRgU
kCRmD28jQ0DZpvlXIKcqfLSOT4EqAS3KrhIW0AkaIXZIct3fh1uk8GK0ZF8orIut
l8H1sefeOWf/xI10GhEWk1lPUueKOqa2URHSUcGvQX42Ia8Omscvf9zMoNK5mV/M
z5ZFUiqvuvvEE8p+Y1BV22JSAVvS+A29AEyJ7uq5ebK+vRxe8XtUTwsA6YmsKld4
AR4fDW76FiSwRArXJ0wFdZS9asisTQPEX1KtAFX+CPpMAMxnBDCENclpWXR6+0eP
dJH+5347Fm7eKZ38vWKSZgqdAvW1ggxQ85pA2mecDEgiUOtP9UDu5BCbS6HEHNNi
t9BqcXjTlu4YvJCt3/Un7os49Vmg5DKnjmNoJ6mnqa5SsYzZkMs+0SIOQsZUP9Y7
WAdiZzjaV48osleT2fVbR1bfhtfDkdLkryYhFKhHJyfc1NS5GTMfxrHwFxhJnJXL
CQxcq95R+so8SykWLDUi8oDwPWRSG9lykSJl7Axdl7XyrCuWR+5VlV7b4C4zF8Hg
uiuxzw8j6S+ACHhdkya8mMrrPtg6D9DCQOs9koMlxnQ35h6gbUJ7TUzk2YtldX/N
MchcUAoqHiFzN2pA6Jb/g9hm2neb5wxfEdPynsmc1/jrSSl5bXGtG30k7eVGY5aW
AHigw08MfFHrhnyI466MJH31csc8WKEMSkSOO2aJafbK3il/mSqA7L+/IJI00Bwh
SxrtkXPns/0OKTF7YwjNevLNhx8xoo167sgNzUcVx5L2hJRLl3FMBPyMTRH8ADxu
yYG/C3abDpLjxqutuNgZ+jLmLSixiElijY7n/W1aWikrZdAYMs4WGYat4U0TtnRf
yVpafvpKx3ueoth0c48zkPS4ewX/ne+uRkTI++HxzYOONa2AQhmry4SsNZyS7MpI
XXyHdMY+Dy24g3gotCbnuII5o/WAONcjHsfky9NwFrLVuyCKxY1FUSGeBYPQsJ0l
/Vm9YJEFP9ivUpqJKB5MDd+50kSMOd22zr2e/HtTzcM3Xipf6vBCrstKCL4PVje0
K0gXjgwdxs8Mof+5ZzobWpAXYrKtnxBGdb8wqxraOxGca5dfKRLI/aTFWkU49d1L
m3qi1TeRn2gWZvC5FB+hEO4rzAFzWRma9bTrBOGjGfmxz+lcIFllcIMpIuN/oB5L
JwsqwcJhNiggD+cezkGtytjpbmjDAnR2xz5jJYpVs5NUa1RAgwGyg9rGoPnwNJ00
X/y0rzmkXNktKKIYD4D7T9QRgfEVKZ0yCpdHq0jczOfck2lKPbqckvy1+zbpPlOy
oUf9SsIEnW0HphOs4Tw8qnAnhanG4irI+SOY4R2VIF5uEiBo9xmMRzKV5tn8Pgdb
Gwh9x28IXoSV87N1M8ZBUxnDbFg5ZqxViY/0GMxpF9ICu/A1evoNoaR97niZZvMk
bzVrtuUmPftS238JOs2c1r67FB8oTwXUqEbsOXQGFkeuSpzHoIz5WOKcWGsX9hfp
/7hdK3KvAYLItvoyNhaVbu54v35ptlWKDEIsvD14H7x6zYJPVndqpOmrvuMLVQ4h
koHltUipgbBtLBHaMxaq2DB5vyRoFScE3xrSmuoADZfL8JvC3kEIAX+VltAPGI+p
AWcpwRIQac2WdW1t5MOsxLuD0AUYZDHAHF8Al91EpzQDM2h53FfZWbBUp6QYTlP2
9Qbp0JI4PpgXSWeRN7JIVaWiAUkcmHkym+Wps0xjDCnEw2FTIYcqPR3952K5waU5
MRajTQ+zvyCosF37viQsCggLywexQcAhgGkFd5/O3jaoc7vtL4R8gGkhDunBxr1a
cJoA5YuK4m1WlbQx7sco4UlgX3DKqfrz0WouHKJU8FgjSa+YkHBdx0IyVb4+gbyZ
DMdhBEcwd1ylc5LmBnd8XX2W0uQE2/YlmGqSY7OIYQJH1jpK2nrP7ojfy1utm1d4
cCcpxbGPWp66HjE0d51dM04E7rW7TYT4RjAZzN+uFoOjMnSIEl3EEj9gUo0NSYB0
4FzEWgDRlD1nXavDuupE4XEWauUYHE+m2ajUjSHfCuwRZcSh7wzCc2D9H28rYywd
9dbXmklqwoXQe64uthYn5nRApMMYik+OmmxzFNxyTgG6rNMbghuxZUsh1qcTz8s9
a2pCmkawfFuvLuiXImn4seX315VEnHYZ4frKiTEaqNmlp1drTveuWuUm0CgW/kV9
GY0iUBsBZpnrYPj0yeMg9WR7pb6+GyLK2X7R50ODIHjI7q/CprsHnu4aSp8ERjTB
yT9hzy1Tj3W4Ca5NC5386CD7/rhPlNgxfBrHRxmuxp1rkPH/tqWLdqeNbvpB2aw/
Pb/qliokZHCNPyzYRezK1d5Txms1ecAvaYUvbsPhcV6V4Rz0brxaAPr62TSbMdxh
eyzxgll7A9aZRVizqg0rm1+ws7KZejeeWi86LMe7HQX8vVdr2UIcIs/b1fhkZX32
NIj61CfTHzIOiR4Ocb3TkzOUHGdfJ9L0LF2dbl/SETdROb6TA9KqrhQIzl5tUAYK
0JhjT6OcQgat2m891TFkCaPEJaTKeFZeksKEZR5Tk94QZ857dYqy/ZGUNjozQaKp
IBuT10u1ffdRlsz8wurAX3tJzx4ZwqzQ1krLa8LSJaTfbb+TBoP3zEk98F0CdV/T
gDkLFWhXkDveltfktTizQezptFZGs/nU/nTUL5R1A5qJXoCh/ZJBqXz7CU4R7dRZ
2NAUEQXzwMGB7FvqvuFpbMAE5K2+zkxcBh5UnJ36JUlqXBe+70/QTt9VbBUKI+Vl
lIzexN47ydn/Wgq+FU7z3m9TgI0Bk701wuE2ekXwo8/HGH/JunEkhoXoxHGTit/x
JJLtUs1AAXFAa/sWAPUa+NhswOUS+VRNGzmpN9dVvGPOwJDjrrqgmk6FdLcmuS3J
QaDzhdB26dQb9N6PMOtr8xpqEmJMtWGCsJOxFNdXRLNG4iItfy80BnTxFpE73whV
TeNE+cdq8WTvMJPwLy54Btqr7SuZNYfZ/ozPzOuoo/ydsVDUCBI8tcA6mS30k/D3
DxatB3ZE5h8gU6BgGIynglA+inchHiJZYn4wg0Wlsssa/wYT33bLdljmCzugEuua
vvuC5eV/xg9IUwdhD5hrtPePVVeUUixdXBIYTy1/rNmvxNRz2C/Y40bdcxgkxHDe
F3m/XVx3DHZPDMhkSNHCYMJZWtg6v/SmIvCGfW/wvokuOphwOX3paFCijaFyBWxz
YVGFtbRO4nlOf/bi8pLawPHjd+ZIKVCNJ+n2hxgjcJpmUh1pQGsumAE6J8UqyTPU
Fn+BofVB5nZZeTO9w3BlbgrKcEHnv1qeajXqyF1v5RWKrfb+snuT87HOgj5vMAPI
Df9dlaAWeP7oCJN1zZP1XfH0zYLBKF8kf3NNYyv87/AEfont9sSVZm3gf9e3PlVh
hgATSEJJ0j6YJ0E9pNCMoKyR9v+lFWFaBULX4L2dmq3ngFrp76de59ZiFsWpal8k
1H0XvUSp3EfiWHq+aZK1wTEeLu4KqvdN6gGxmjF0I+xcgrVuFm0Ezd/1qH/iyFSB
J0wb5fNrckYGlWRaaOiwixDUhl4pDaYKZoeZI1GiDEALV3nXqW8nXE7Qe8rAUI93
Hx0CARyxNmPoa/Sm7OEcUoFN2ttOj7wuHKqYQ0XIdaXxGtWyCgvu4aEeWwhgOftS
hgoYLeJtFr8r4Ay3DeeevlITCoRJn5KJAkLpwJbFpuPCTcStLgqJwtWsnRuX1HRY
vGdKI4AL+vga+zQRUoFAhqafQxAurGzQElUtvsna2TPE7ChvE79OOXVbSGuiRFiV
Ga7uliJpOpedwOCNM/Gh7VMuhhzJqbvAwKfdMxvtkal3lQcaHmINMvJSgtva0vdc
NBTIJVVlUpLOP+pZCr73b0K1yshXhj5ElDscg5x6fd99qARr0/H89DSxlaRsR/Gg
TM9Z0mfM6wrGOYgXakvqHUioAGok8voc/VBM+9n6b2BSLlMcFt3mKg/gF324rILx
oDZaNb9upEvUdiqpEjfXwsyqylFNXPfow5LTdwDhweSob9O6nx+5lKtAfB9KkJQB
Bw5/lLeM1DHYjPEJl5s8BIcRAjniuaToWHO00e0YUegxihZS3Dnnyr3ZEpqungSD
/n3FbCMRRWFNw6VCEJ6sWf39vxSv/9/EDWVFvoS3fQbqWx95GwRECx92T/FG2zFD
sI6v8p5sO6Hbo71jvGEAegaSVWd3+yX6GAt0D4RVzulU5Vwo23dwO6Tsbuj1J3op
yKcEZ3Ug+LTiqXE0IVMY8bWNOONSc24l0vGm1o85Q00gkNIqIY1w/Ud2TAX9mB7k
bPBJQXxxXPch1gGbXx6icv30Xk661phdqOd+HIZ8rFt5eTEM2hOthTui0ST3I45b
Airc+XrNZhjPPxcJBQisxWP7J4eZWoeNxoeas8609+00cJK9vW8adAYK65MyY4u0
FhhtOXDWpV9ecNqbfzr9gHfeE8Yzp/Ra6benZnam4XrZ84KmaTI61ELFrUIGfKWm
1+oyzyLukAAk2L5/yCuIs45+pA4+5luvAUhhKt/2MKIChajMF6tSBNOaeaTAwTnB
uf/NgvVNDsOpFej/VvyF/U5cysvTp5GuEHk/U2AKR3FAwlv9GVXRbjOvDe3e5vlt
O5iFlTK4AdSObB7N1f4J9wQbqSr8FjqnN2Ye6Ni9S4Hkx2rY0slo0qzn9nX5Lsch
q4iopvpudv1y3zAzY06NoLBbq5F/JdxUesecSbPv8JXlyjDfOf7w71KEkEdwQzGO
2P2aN50zqSEaSfeY7Bqy6bCYK6ilkugzb86VypeKWuyBJYHmk/NKsWDfufQ6yMDH
/ojI6IRIJQ09vlo3PIjTtp+ONkPbyMq5vgqudcVrcqNPE6TKEkPqWXRUq5FAWEDR
t8q0reuc/KcSNTHG6m9F5bYtJR5oHPUkNxec8MdHuj2NzzaMzlPJP5HJfhppd7xf
sg5Euzer4uDqJ4VF1rjpfTjZbR3R0/p2xnjrMFMOpf7pXgb4eDaqECStwHmi5p0X
UrlifLWmqi5xYBcVcJnc8aCrPCXmJ1e4C8G+nbFc25sAGuEZs2kJkimxU29oUuTB
Hx4U+YHmJOwO0fzjo9HyX52cmssLDq6V10jxL4wbBZTDttjfSnn5KsUt561zzzuP
lB+Z/cFFhlL80FSMVsWtdYGttNQqQpBas3MYz/3U1re+mCA1CWCPOMyHZf9V+icS
ScPSBgIpX9/PKXzZDuFC1jFCSv63jAnPOiykibjqU7wVD3BtrX+Xq8Bll77Sre9f
4uYPmByiu+fL4pOVTc0FZ0uVoNSXmc4yRTTa3AXzjlFQf0OPIBNsJop4mpTXKRiC
+Sg7KEOMLVs7SuYnuiaVfTOFyBV4SOxOJU5Er4lQ/+tMlzmaqvWAPi09Rypy6+Ah
f6HDA2OTJoJgtu9K/Rrt3WUGp2+T+WJdnb8RU29TDsn/FQylR/hDIfDfA9xekGNI
qmnuA3PqS5o3ykJl2KtJzB0EhEphy0n0z5k51WCt0KQFriedehMQUmrqVR3S7bcx
cK8ymr7pI0xNUi3vGYWP5XuJFoK2vUg6URDCtYgLb3hfwrc1yzGE/qejXQccGBZG
61Z5TZIk8nQkvfGc8Z1xA3Z3+cf60OR0vB8h1pe+FzlkoeLFoueLR+G+cFZFgZ4/
c9xlISBOw7dezMVrn3cZhP/hymI79HaxK7bUV7rWhrN5kyRGO2LL4hUoQR/MGJXd
jA3+7i25lkun6BKd6LewwMOsXYBTB8dOH5QExzsywDiPIL7yTSli0lomxf8RJGLf
oSUnMEUIJujwXHgMvEvUujU2Kd/Fu8KLPbEW3fiOQNUjXtTmizPKVhHYDxGHAJ+/
0CODVrdtwdR+qHeQ3zS1M6tNxhOs52Lgm8oXjbxeAhSjLdWhz9Yug9wAaLSCrETf
vI79FUPo2HyQyNglKVleU1F79MVSCCspZ93ygNUktkWEHhjcgnaGT+J6W2VGv3aj
lFjmXpoALAa1dKqUzuYFltpMHlVTrOiCi+QvwL2+X25phdsH41p/YoUGbZz4RhLI
iaR2ATZ4tFwkb0WX5iKxWZydiufWqb29mALq9SPEVHioZAX2yB6WMy5wjiT5pQti
/6qmjTzDDazdTReoGgE5yNJJFeWJhVhjkfBRTuQJBZtB3LnJOdN7VpRlsFoqomap
OTi3f+EUNXr0ecrbTqBlFLkiCRLgtt/G8iNDGJptYldbanAbPHPcrXDbgbh/RxJo
djJOtkU6KfVB+wLXxDe0MzyPoX3OuqEMkUXJ/5zTEyjGgKeJqK6/Ow3pUGbjd+0t
C2nzR3e7M78n0Ll8y0ARrXSE6eOeHPGGoo0TeUsa4veU9up2zSk0If0U0yApvTgW
uRZfg0AjSFiWWjv0LXHP4dGh4JEmLjNnsCfE6Z37VVOfCbbZJvnJwGWFwlP2C/WF
0O6r4OcjekcsqHTbUY1wFeZWekac4zHBG8+zltSwS8RYiYPAW3cLXSUEDmVjtkr7
h7M1rYxBm9EmwyODBbOp2u3PZJbhVP3hwLX33wSW2RP3EbJv0xhWiAsa+QtuPigw
ZRhc3FBmrHnLWP8aYohiUupxUN4Q5tuww83eERukex0q27wyR7w7mdnEfrInPYdn
oMuxqlzOYlJ71xeyrBeNAWrroeW3RFE9WTjjEEn/8n8X8orZuEZrOhSa9GGDkReZ
MJDkwclVAp/cTLRS6Mkx08VP6gs+2iG/ax2mVDzkyt5f4I2ZcIdBG0UR5U+HEHlJ
wAuWKaqLpXLDl0ss728wYmdSTXsaDztnXIS3SxVvsp1d9rha2ik0M9ly6DrPF0Qd
uEzPTT0dp5qBc22brd8evaCYV4KbbrZrbVxzvsWIYWTDu0yur9e2WWgw5ozNvlXI
GQuAJyLGW4mYmGON/CR6tuf+YeD8qyKVapHXwbb04O967DHCZVFV85XO20rxNVq7
Uyv8BytSeOoD6BoNIxm6DO7GAJgxMzbau5O37T0/tKV4U4FnrFJ76JTS7WQ5Pxst
oa2nVGY+TD631/46NIosWyhlXTF/7Wx5de212paSOGs5stHkYyXYgea2xSIz3M14
PZu8MIlnBgyl1z3aHY8mEkYjtAu9knuzapk2Ix28ebHkqS77E/9Uk3TawwixZUvZ
Me9fXiVu7YEteLmyVuhyunTnN5Eb1JfjG0Lr6MrIgnyG/7K4NG61B6eHyl/HIzQW
zPwtR/aEITZdfhJMUmFCrFoJDpTcOO6UyrrfsP7MzAsIwsEKqSpCMUAbKotS4MUz
rVCp671uABAQkzQFJ/3h98DBAZcEPqYp6C3RVgNZj2CaNVY6ZRLeWlpu3KOHtJxB
M4/xMh41y3HOOqeI1jpkW+EFvmc/L1bKMS4g1rg6Z+syb8ig0SjdR/nFf79Gteje
CcgM2thPIyv+CzGEStyd88zqwX3QWhjXS5g5qk+6esXeBTTb9rTM96XyjqBgOJA0
nBib3Z/EWkqaZzi01E85cO9yxtKxmin/bNsEa3PRfH2UyWUpPQPvq2BPLy6fnJfb
c8Zz0dwyhFq7OIXZCdULQzsJAP+jMoFym2h4FXJS7/Ej3W4DFrbywT40Lp7PVlb+
lQGAv2KoLWwwDAwvOyK0SdjrPlLh5yNC4MvNbWuk7W5T5PlEhuBNkUMegBedBsS5
9BqiAlmyiQk2Tj9ZF1OctRfuHQG4YUgtASsq4gyTeFchDLvejJp2LI2EnGK1JwPG
Q6ZweYA5MeBse91b01/hMJyjybtOdEVZAKFg8Uf0vqNtp8OBZKJ5jumzTDbmx3uO
G11UoR2gLK2rOvIWYvJPCpketm4B3UrV/l/AgIXvqqImxgfDEZgyzot86vcAYsVk
2dLelSZKEEmVlBg8Pz89KMviJttEu1OyyREtfb5TJxaN3jA/Z8J+zeIiD2WmPd+n
gDMCkk5gbOWlahvs8sxtF5QNOtSzITsawanpEvJ4prEzyB/+1YUQK4/Ea5FOaWlF
0XgO2P70dYHtlBagMCouH8qv6ErL22Y5fQWODMIIGqj5JSSojPyYro7ECLiAmYH6
8nwI7tNGBCYOX10J/1il35LhhF059aCZvhTgekPg4fsMUyS+Rme79pwx0dFS18jK
7aqsE4TO+JFvDQ449dQv4DhJugbZ53UzQL94XGwnDLluLoAy3HeTlMn8XjlgDFQt
Kl/XnuKlEDIHt2po1AU4YriK1nQVp/1JXf0/StzWiG2FeTuvvwz8HcEVR0rlPCFY
Gj8ONY5DWsw/1osOWks/bR+2pyjcrruajvvNxbr4Mxmj6wj0OgXKHL6RcAcVKkeG
5eWwDduTJgz9MYYRGy1LFaUVoCg+Uz9GrG7iLGhlcTKq1mgPc9rs+l7OOsKMsvE7
Dx7uq1aAI61caa5atj2geuy4YPge9EJWHrZXRw9TuS28RMRGwZEupDjw5UFZx/2a
5CGI4UWheGl5GNE5TrVFGTTf0LpMOuXJiFJmextlnXPBru8eBnYg3avmYuDigrLp
JuNd51WAoa8bxdDWNBfKpi5O6+0J4E4gVTOX/5YDABv/fK6PwLpWaLT3RAm1FRTi
KC7pO7+yaaJ1EvIOnqHSVnuSB3ynLHjaCRZLhP8GJ8b4BqttzKUR7BH7JFhFniMm
2wmkOH8CgnHq0QPXVIFPcVMX9TcVMeeX2yiow/EB5Og6NBxL4VtbLLPrXCg7Bc9L
0d6xt8EuD6qz/3SjFKByORbd+0XRXyrbPA1bJCx2DVRi7a/eV2I0QbcTQ/EWFk4l
Jml5qhbplSqeJyFc0vBC6wRTy4PUZX3OdDp5LhnyVhuDOI/GBjliaAwpV4CqRCjE
4f2cwpML/efq5PO6fb6NmSao61KHNbfRm2GD3dNcgwad7ZHl+awBURI3RIxlLkcc
mEYUjTNlqQCia3TZ1jX+p9dWxnv6LH27rHNn+AdNvv3uobq5S3w3jAqccD8pJ/cf
W1klO5sqOAHlUJKrTxQXQ3DQ/DHXyI3l0l8dhOeyXeTC00vE9aF0f7ItqRPRFoNx
s/GYjNN+m8wKwJDp9wPwBcGAztrISW+5WPBBuRcOzPszV+WeitAU3DU452NW/jTT
UJPPG4MN9+uHOOSQy3Od5vAXQjeSr47GtTPduf5qweeWFvlFrNFFivHJ18rZlq92
+afY63mMcPC2TtWmkLzCxjijZMQPjbW8kq+J08NP1/teDCtCtoaF90PGwJMpquqe
EIHK9nS2Qcy59zvukq1j0ffCyjW6Ouomxaa1gej5TvqICCIDzsg2oZszb2HtJQ7e
WXyeHMMN9SleAPRK2SYOa67/rrnphv3bB0Ou7CN/TCt/a+Jh3d6mI6DO5Q9MysKv
ey/iGeSNetE9IOFsNqXMIevxpnmr9uTHHyDszwutC+eU+JJJJHiX5s6hsznwb3J7
P2b3lzSKwzxT0eABth3lHzJ8o69b3h79xG6z16M6VmJQ1z68oSIbGygHsGwU4Sr8
zX3pOBqGpnI7vGhDAxzmcy5W2sJfeD2Ehm66UejrvXzIOJcFvCUanrsl3ztwjdyp
y0lYrRnb7C7qN86kEob4AbJgfBwsvluAlWXJvgGhVk7qsx0O5KLVDwVG4izFB27C
qaR+Ax9exWyMb2Ih4s+KlQHxAB1V8uaHz/GhmnNDj9kyCpml5A0hePf97ZBL7+cS
7PllsRGSGUGIFGVP2E3duZIzRVQGhF9lWTLZBObXLIJ4ypQ8f0ik/Kj9yAfRdag6
0s1Lg0TjacFKUXfzY1Z18rd55l4mao2f6NZHPAj9iOzQUBpQl1iYc6AwWMMMquql
TPdzm3J8qsraQgRjiCvTCvW+X92xulHB5CNTYI9yNiKTLlWTPRnJmJK59jeyZsgd
Icqfa2ZQTM4ZxhgS12rKwHsHfEuvvBE2qJnBpRwVqjN4UfwwVnukcsJ/u0UfSQ4j
KHTLVaRJJRxWksSE5tqECSbq9mPG0XVRGD4lUnjBb73gGRP4vQvc4fwGWpue9XyP
3ZJuUycymYjBcX05rJUXYDAxbJmjdAWuSzMazgk3TtLaVIhXykQikafyfoOcQ0Xb
b/X7JDibSd7UWKNRcLkJcNedYsPDT1wTkN5hKi4eRcRl1fuazZybrLkvBigPMWfu
ZmPvgIYjxv6pIvMNETLY0UDNXm9SRHO6i1aXv5qPJVFy8JW9+Yx+LGUnZfybmqCF
N/3ffa0T4dURViBJaRdURmA753g33mlT9khQtRnOypRXIduhpszSvFIpZvhNYZQS
7Nbh/iw+W+q84NFAC0ofBWqZqU89lqh1zpTnATzDmATs+PGrZlnuXmQ3n6BjvH9V
PqlrBSBSq7+QNyMrsDXnfkwfF6RJpPuSArnHF92wnyvODkRTh0bDzvnAdQTE4Som
cli11oHoXKsWp7RuVOndQvRrgFWfzaLKnmPZ4Xz2uxmju+zsCBHjwm2gnrQx7fMq
Um3Aqohv73vb0Wzy8aH9Dp2HnL7C0Gdt7KWrkjwNhv+3r9XoZBchwiG++SfMNcHP
6j5GKw01a80N7n5nqgVog9ZZRlM1RC6ebK3dpMsh7AjTmRUyQxdLndm2VuV/P/Ig
1JCuIaPHW5gSn06eIQ4yTdoeqp+LlZAacoC9r5vZFgr0egh97v9ZjbVO5vkdtMey
PAVvg+MXJgdHOvvW0tbwQfwSCfQlnMoosodqF35FV8ZinDqlPRk5534O0OjBllUl
ybuvl4o88VxCZW/SwdoHXh4mfTAPka643WOSo1+4d9NsK5PaLphxaNBmUgHzsFw8
fUX/aW7TDTZ/V0KNTacXbVq8ijDV3NpbHPGsbX9OA+ZNSmGFoM73jI9wVaAl/9U3
EqDNMMeqyQ2V5AkCWQdo8KrljgvEnwwqqrRFGs+ia08jjm1pIIBCaVSHmWzimwZH
U1ooH8XRjyrogo/0YeByfz2WTkAAPKg4IyUXy69Qv7ytWLKjxdM+AJ7l3scrztZ8
nZ5dfiRZUga92Jk/zkF5tOjf0UIZyJrEOpIbwgiJ0ANUpSo54obIF2+EBwpuMXNN
2ZqfOlKV5ijJ9G5HAC5VH3vbK/SZjdncOz7Sjk2GdojqKlwSfCNQtNTfi4PGi87Y
i6SVLYwVvo8YiNv9/lfnWLe5hP/LVtbCqke20icCvzNGKXxsMgYpyWuOZJTlQFH7
qRw8pKh/VpENFK3RRgn84p92vC9qkgdBhsnPDgaB2xhgLMc5Gyxdor4ofYwHzphh
JizqVwYkmEnfVZ9KmDQpncsxciaZJxdnk9k7H0C31RmIwLbgs4UfsA5DieIaI4ei
sfvT3GL4sH4xgLKcszVooLqrmTXtDTIDWmd5v+yK82hpnnoet0AqvI9M+DgodrDW
WS/f5jpqNN2j7GoeCY8Xbosx+N1iW/aEOjXRFYKucrNXTnqymwzmwQtpI259iaBD
DSAeMl72LGnzkBxd4BXL0oxfjeilp0VuoCpmItAvlfShZER8iqRJq0dirhmarGdA
C6pT+pu/xVQIKeY9N1rOP7n/JIIMygcprZ2+n7AwBTDLomTm32WBSnmpsg6prxQ0
f7uuJQ/YB+1nuaFhG5kDejkK6h7BR562EEKrNsHbtKdQK1Obxyj7nd1knUuwcYKz
F654ic8fQSJB5+qNDKJfAh5cNbcE/EhqR4IqtPg66JkQZZN3bK/1HnanI+sscl5j
hIefKyfN4Qo10Tde8pxgwoyxKQXzTuFB7QiW/QoWf8F7nkK3qQA7M/Ie61HyLD2P
kZc4nYmprsWUnmiew2RNSjYvqnwmwV6URmzFBs65PbhcIoUI7EuqOWrMh+Ny9aiH
/Ih/ynCFKoKjxscg2cgnutFkuEdoiP2M4Irf+VROwbrpoD5Sl/LYaUX/wUVOp1Jz
yhtG1iMu8rEqYcR3WtNK6VqygzNPvtazEaMqwnfkswy6+C4vLH2/F+yM8mBMZsXc
U1BXjTWaPpQwL1WpV/jwrfUAlfqV+JmWjk/iuYfgDLRkZf/d0MTqtZjcDMZaKjZx
Lkc8IvcbeA5xjumC18wfgcuolT3StWwKgwuAjgzqF52hLiJ3ZlLsYASvFZrekQb8
FixnZTjHHTrr4cw1BpQU2TS/3mrGU1eOlyxaISSrz7Z5TNnMSVLyXk/jUgPeJBYm
RUy+Z0u+3hvwHhYTPCEYq5n5QfD6VAu+BXAkU45tj8hoVCUlMfaGtj4T4Eacng/i
mTGJGOFHvsK5i++O2Gl4GB66pcMato9pqZkt9zD7MKDP0yuF27fUy+Dry2e6v5+N
XF6me2QL11YTbjfWGP0waXA7pjxfRhZF4uZ+02evoPfYdneopSgyLimFgaWg68+8
1CScq57FPU5zWUlmylySddShwN2jEbkIqPK/AJaqgodsS94HXhHMMDeLH11hgnzf
UL0gh7RC91IhNyUKqFT6SRpJI2HP4bawEzf8TYOttMI9smVFE92Jp7OJS0aEof43
QNyZjv709QT9TzzZbwXqJoBjOaBPQBR2nIQEV6HMKVpf7BpwTxUTUdiAyhjVBRKJ
dGqrcurqCn7g2ahK5QQuWD6j9HWBFJsvRUeSoghmmikLDtwkWJxWjG+3BZgav/Jn
4X8u90/kiP8ZhuWY1m88CBxf9xlwcdwW9LPiiTujD6UFEdTdfCaadnXdgKR7Ovdo
dFnay6TBxcQVdDLw/YnlMAs/3O8tJe0o59isQZm7R7M5ZR/4R4OaFfpi/RMx/Bul
htJ9632AU4HxZlp5AxLOtTpKxUB/PqeI2q3k32kbODT/RNObLzGCOgxGxNBZB+11
cmcB+5YPiNMCjzFiu8QzaDn3bq9i9F0rLVbo3tV2XV0EZMq1ByXFAcmxWHpAcRja
DWHhWwJJ0ua9cq27+PQqT+YBhswaQn3pRapxvKeQBw8wNcZehdeVxuCD5AY2NdQ5
oqkf3XY/8K/j6p1LFmBY2SlG31rmWKBwrMZn/gTB8shUjprLqFDLmqdWVP3Q0Kui
n0dlWRiPGG4IxE5DEPmjsLAZckhXlkGy8v/JY4Up6xYzDAvzMfGGV7TUN0drMzxw
JFY33MFbkLeGewJhBAmIg49/tp1JgOPsePkoVVrufcIcSqeZHDoPY90l6sJ37/OX
UZ3B1LdGzYDGNGMsejHa9gTzYjx1yrpimSutjP+5DTab2UwQD+V/qPjxpSAGL7Om
jyTvnyKw8mmAe/xgoVWyAIM8BPQtANsq5OYHYQyUXSb91h+alMXl0wo8+pP8KVms
2muwCiJ3on8r8EJxc/NwxU8ac+7gDEyY93bKHhkqzR9FXvlQBeJwAlsF8WHC/bSi
3SwtS+r3xgC3MI/UFEkW/o356njOVyWVlLrWkEWTPfiS1Y4kVrPUEX0KmQAK+e+k
gKiKa3uCNsga48Aoc0j4mNzZVWXqLQSCkvnBfhfufAatB3cOxEJmhMdJPLVzFVBa
Vk5JkAh1Ozy7MCpoRpDCcLjHNjXMQNuz2LbGhDJVPqmhO5DqOuT+r5EReWyE++lp
a+dDmUWg1nyeZq2L4b+Zpu7jsbDQrDpqB4ExglZ1TUWcGBsxt78vkpctoNpX5+bA
l6Pjv5JrzNKaHbo5LzBXae69Frpxpe+DnEGXF+GLLoWTrHjqjB+Z4J0tf7fXInFY
84wdJfLA+fAfw0+ZVu8n3EyQ/2loN7V2aWzpm5/vnTrL/LYdSZmb9yjAnbxXmFya
qsDKICFXsvylTXQDvAbrsVG3Hmjqa/zYaWC6w2MiRApxN1fh4LLHMzndtjuxUhQ8
UsTEVgQOhd46+ln0S9uPOsfkeDUY31jXxzp3Wo0LfQe/eIihQK9GpB2g2OZAHA5y
S+W3VMlP5FMCU05WoyThTyHRzmyDjdfpIn5XZWlDiHmAlwMcNVaiIOmDZNaj9zrp
iqR6m96wNYTwkfMPrJ9ldJDynrFF/+vr7nwWGsYBtjDYVuO6AzbalXhfTcp8iNrB
pXe8lsb4qr7M0nQUDKJ1OVwbL1zMT3kQ0zA1UeoVLh+Fwl4BU5wKxQqaWuv0LBvw
nJ14bDltr7f+fpo4pbW7vkm9fR5PADzA6Ozgef/2/JjMhjnLI0JE64bI75MtCCHa
jrmXiOikKsExS+z014dK66kpVSYzhXGDArds8/BVJaJbXHRQtygdkE8W6RRvL1zX
lV+F3RNXE9/1kyJNlw8qi0LInRwiKRawrq2G/NLVRD0j7NUtMEKN/BDgHoPKQy6V
85qU4JPyhx0AqfbcrE99Ej+Sktz09+lFlHOscmc4nuZCsB0UWawfOMPsJW3fWNzI
0/XQXWGTryf6NVeGjJMexg0L44g0aVRAfvdS1LhLTAF5b1Jckbj0Hu/ctx6gFoKB
LhDgNmOcpdwDc11ByGhQxF+c2h0PNAJc2Jd0omM6Fr3szEAwEnLV9Jg1fLobWzMf
IeCH5d0QWYg9wdwzAMsLoD2+sBcgTBIn42sTT24eJs3gI1veOdTE7/0r415il9qf
ge9/TnUWGs7IUsAF+1qJaxAQDnDhsVyOG7xYzo0xesHuvi4n0Era0cLw2p2kmB4c
jzBYctQhj6Da1VppaMTLKqbgJXxgO/nkmBaaakfAZ9YpMr3ZjH7M9JRs88CvnxjM
q4xX4AIM969OPn35Sl4l4b5/TAFK/xG8TsYg0kq5O2ZOvOAwQiiBpW+4py2K4AcF
40dE2ZE7Ib0EEFD7CyBNf9m2oh7wzXHR/QJOmrhIuoitfKjoikIB0TOXUq/s6GXY
RQju0MkXDaAJWqXudCP8NE1IRA2e7CVlM9pPFE/Ay8zUvs4Ysma/RTjlDhti6fTo
61iYgnXqIWxRPzhWYFKlkDUDCGkOB8/sV0KgduupWQHpMg2cG0mzApK2lq2efspD
gcXfOIPZKvb/zkStUWeDPpqYYGCRugtR+RJ7v/i+wouv+fk9rHuKAtG4yEE3n+D4
Q7rvTgs5YEq9mRk7z46X4nVgjQbTvJxMnTW/eSu7MWUP6tcwfm8+8fKKVCN78ucn
/PuliDXi1QLHxyS3GwDFkQw1Gme1sqo5huNK0PYVxYxi5Xa1SzzeuTZtP+MfvMFf
rjLF433951MU/ZnqP8oBAZ55IzqTF4VYLD+lVKrI57BS1Bqso+80OGZeenRYKYqz
YrjlgPrSMs+yGekvDH1jT6UMqiA4zVIOpzklhvOykQpRIl9QlYLM+pn0+M4+GGgN
Ddc8sgNC/dcmGlc6oBbYqk/fAL1sM0ZjAaE8rYZOpSTJHi+VzH4D3kcnOPN5KHMq
VFMTgGtxspH3m+v7d+++m/UaZQjorsYPAVu5zGsr9eaidhH8liTQ5kDFrtL1BYLf
uCLAf5ArFLzfgFnpd9e0VbRE5FlBD6ptPN02cf8RWHayKlz5Z5HDzxuYcfFkILjF
3dpeA9DtgJ8uCden436jZ02pYd1TpeAO8n/I2bigH7ILx/nfxSLVteF7CapgH6fv
CiO2ugTTTYomrfErvM6c0RPK165ior2Nb/Asl1ivpcU/b9llAHu6fmoOhCEUN/wt
f2luup5qzuVU/vXebepQqC9fzyi0vBtVFrwOynK5Q8sZ93TqIdzStrJavfXyFt81
K5Dri7YL6Z14WfGilt4uHlORAcT3zNgBc2+hVnudV4qqIaFam6NuKH1QUIEtheRw
XomSFLAU8c6MEmdK48XcjKB6UojRnHHo/1Yqy9qqMPIwCDwtQ3heZiMEtS0QtrEZ
bPtFyGBeRgWmNQJVSZ6fL6HTDZ9qSzNuJ5wZUi20fviSfYPo0G514izuo/Jbo62z
iofAHP/zOtC0j8hAXP9r9I8I4JRhwSO+lnwFcP+1xDEGfaDjPmTfDUKydmwT86GH
CmKwfFaib0/9OCE9xjnoRgJjLC9+8ut9Gpc0XOgTJv5PJ3rN1vJtIXu6cHZOfVqG
LEPsXEA3ucqJGDt29G1xsRhHicPWDKVLHVH16uiluDmftAPa6qiF8jVRnJgcwF6V
LsN+vZeatjp2JF/jtgrsuRwmFCxjKn2J9Hrr9sPge8V6f5p4ZAq7PDdu37pMYHMx
xfh+B+0FpbpSw9+9j+Z0A8nsO1mHe8lV4unf9TucBrG3a4764aXR3zzF97o9DIpN
vmeV3ESsCree74UxmHhvr7/fS9ad+7SNyRrGu93p6dpHFLjkjLE4UnV0w93MTzZN
KNHQ9qFUVcWP0ePeZo+jkf5nA+Wt3QbWGcncjfoXduWgHmqKeUlMxVlq7jpoz+RW
wdZbFbXLQGH+rtDqx4pRHns1sg8WTM5SZI97tDsDeAnBEhROm7pEQjnOcGraL74r
yu7rfFQ0VSPBVl9KMzjX9FpnzVIunWZS61GEOVKX/L5yNmFx7g2F9FrrsAB81DRo
Ljm0njrPnEaOCiZUOEiut9UCnjWYuruU6sbdNSjs51KwqOMF1uDG+I5KAB16fevy
gW9TbaJAku4gvjsgkkw+f7o4KDosRUCM3WbxtLIN3Rbb8d1zvkNc1MzwdW3osxxn
gCsdQH9SyDcMHZYeK2qk/ujeSQwkdFVcVkjIpNFFTeih/14DWQWxmApy8XSYFqYr
5RjlvN6QGs9giZiyjP8+9/AIJTUIQgdHpQAI0S9UcjnwXmqMe/ZmSrRdw8hKe9If
uQlCKgAxT/UBmTRzr46kkdzQKdkI4D8HDkSVWp61X54nokvQVtrc8tstznUzYyCw
ahi4+VnaQbGdEbu/WRvs6Fmw2lKoeGr1ezTUe6iKmKp/Ie4zU3a1Y79SEQsVU8Wy
x/yG4JvVln2QgS/hhFsV3VoN477NNhHm+XjYVkrjRqRgxQ+fq3NzSbl8pIpXEcSX
2d+V5hOy2t5IRIm/EOXWRYZZZQMyKclyyTq0C/osT/vCgOgaHlwaonK5vG8adnzt
ysNMNE5jxKGXDeamW26DvkzKZ6VPuq2GfEfw1o+El2xYgtB47ocO1Mgi9PnuZ/ah
+TPfUW/v3Ttzu1AuY+SBJ3Owp8K/gmB9tKDf2mh72npXuAxK/oBqVaB83hcb8BG7
C2OO6QkfBTh95aTFD6CVE0MGFU5fEtRLTmFP8NPEAZHPBLUGE8vMl7o/hY2kTzcg
COBa+mfEW3tgog268Heg51in9apj2HRQxAzd1M69KIfBQZbUjt7l2ax4zDqASlrn
1YyquMEnpuqZbH/ziNEWFFZsoj3ajvkz6QCOs/yjvedi3yKVy4KnXWWGoNVqXpas
Bccvnmi0hrWr/dz5A+zPs8ItFzsoJ+4ANOmlQHmj2W+wIsGCV57oytOkoqwOmMmN
eqY8Y1CFBhE7le4HsMaqY268pG4IZZ3vmgXswplkbejE9ywR30usEBFQHCJS0S13
pLE642qIk6F07/T6kPrHsz4Tk+/k8PaoSPlugHmdbENE0O6L5HPpA6PkqIlL0k9B
zJ/Z2t+3ncvC5mYNc5RE0Zu7UYyFH98+HuYGGv4tHivVUwkoUrVJf/0AiuXAJNBg
8BXxx+VG1sj1XGHzArmRsRT5SV2R+mHhXwxXYWQWeIYD0+QTpGYz9LkoIKF9lzjS
/sABcOHnZ819xOuW10Qy8CqLvrIC4EfYQBPiCC6DC1OYg883fEItbYdvGYceSCZU
xVosbqTceW+2Z1TrL+RsgL+iWP3da2YR8dLTKLTPbKUq28II0YaOjKUbrIP5EPZ4
UcKqDZToAqxwkX0PeM2wJexBFCpCCGcbHyz05+YWA8D2qBXEuJquTZTcs/iRW0BK
7utbOgA4rJUAgWGYouC0KWoE5Ma7Z9SDsTxxXMYS2Ihq+fImElYr4ByuqSH1FYsS
gEpkj56wiypCcQYqbNFx4rhWVZl9xi2yGBpYWDMOj8tFnsQhyhsfpbE5dcrhc2K4
O53+TrUgQg+EgGiBgX1G9qo27pZG1/RX0lAl1Xn3BTB4jrwuVbCG1APgS+OPM5LU
iJEtLN97borDtG5+llI8JgfMOHtULcQl/Hf/4FCZ5qBywcsRBkZiAks344Q/GqyJ
H8zgsN5Kcmbcd4ZLC/DgrmNtf+s+V9e8oQyUJQX/b60uCjKqoULoXAo2vhaAza36
a4YdQms+uV2qK6iXW0/rw+TYxg3gnoTUTrLRhRubpjhfzWIQqeW3SBZChlWq1NI5
PdgQjYyvlODcKvyiiTT9Ptx9q+DX9uQiJ2wZvv47ymzJoDPH0HMdbem1im50uXVK
FrUS4pC/TgZDdNeffrE49rg8trey+R57YNdcamycOsCt5DwpaeKuRgP6FdRR4i4r
xUQkgkC1EJn51ei4JCNgAlMfd415f55gfrOiXBU779kg5EL+ezyGSvyOEWcK2/qF
JlG/EaoqwdFU6xNThX+28tb3jIEeM/T1Y3RinSDVCDsjC+0+8yFKG6Qmpw/BdXqL
eV59pUy5IUU/vjKADEhKPMmg7VOV0nnXr7/0wNzwI+11L2tOQlyEA5mlMnU6pgeu
SW+CWWLvfW4ycqEOZPJX+rrTI516Tv0Xp8Ln3xW+MBa5pdHdsfwKbsu7L9NvSizE
Poz8hY/T9Zpk6paEa8Zw6nYIW273SLw8/RINlhz1bm2M94e8eGQMchIgueXqvxzU
xvAHNDvVzFwN3mPBV5v4asRIXoJC3jMUihxaCNVkBIMznJabjIcHJKyASd2Siu24
xjadbyF+dUEVTUrWUlJ/TB3oEV0yERrGbRGoPZbz4CVhX8AQarQqSt4Mc5dc2Xsq
0saAEAuxFKmYK0nVJkZ2dv8cz4nSrcm2wuHyfyWoDcCyUYX3xsz+5drLIUZN15jO
zLdN/WPInn0uadS08Oi8U0LNR/SxQVPnZgWP91otl82EuJgOob76+FoUFLAKKypu
u8JWnuXXYNPQEDtWh3ftn3keSRB9rK97HMqY9W9gQRSNiKzhWy9JkcWRFH5AkpTG
ssw6IyC4Eguco3jL2PR40DXph5jJV01Nl/QGhzF/QhkTZguJ887F2Wr7SJK28YMN
uYZvdWhMM3XHX6HxHygR6ShSfteDhVYSKKzvg3NxcgMsu3l08KezAy7ZHcvNRafM
VGvesBOaezsFH9pBUkVN+13XTtI7ttS0NKoO5ve4fN7Aqks1YsSWGum8yi/NtjLc
W9Mn4Ob7v4urKr7gI7X3kJuiB1w4FWX0Wvim1n6Q921czZCjKDxVW0xciAvc11TV
kNRfCP5GxB8bKi0JTNeIC71EO+RiNsmpBt9FN210uw5xSkotA2cdezl+G4Ie7E+x
Ft0pojlG7nEvgFUNNZ/Xfsiw+9hS6xy5rrjjr0fpYBhuxJx/0/bHszWyy64DO3k2
keMi0wxwamOrkn0r1bLOVmk1PnFD1aWY946otbArAMKesEwzjGXXjDdZ85hjsCRO
OsXuyPFLJj3h611j2D3wQBOXrmBy4upimMSj8Tpun4pDxfECnaRLqqDbqwXSDaeP
dSjMO2rl+nMdyu8PA+qrZSdOFKHCdxqOAeNLkVbyKJiqJU8NMEpYGKz0myrT1SG3
TmTG5gp9evu3JDS5GxnRl/2/Ye4FWWbess2+SroFU9YbUwIjlbe1OB5DNqzZAipH
yBO6NezPHJQhAXWU2mhlMXXTyEOPP2z1UyHLxSD6Zhs+uCa/p0UEB9XyXUqGYjC+
wwQLYu/uswA/n1gOOTl7b7w3C8PaOASItyk4mqh5GIIs9//3IeGL0h595V9jYYKC
hXYgNIOhWT20+dYWzXuhA4vUOQnMgQ9gfsS1rc0NIerITPpaK34ZBNFa3rlXDkeP
BAAQrSRTwZ9OXqGuBshJo2o0JO5moQPUEWzB6z7UB2DGHDtw+4chvAKunLynUChh
R85BZ/w4y9cjYSmLdN1Ygrh+jbJw/mYNLYrTwWCrupQ9DluH/JpcrVGnXXzd9qxF
jCMvO4aJ8UoUWs3R2++zEUAU9sYxki89KxnzvYSObaXFdT0vPr7ncftgnEglAzWo
atCxzD4TR4932bvF9JQUh9p1T4tl8xXJkSGvqYjHvIgQKKL+/8rExLh26I00FUmX
rScA7ZpUkLAgQrC/CKTwbFEA4WFSgHluI+EIS5rPVAL5WTMKgIgkwGnDPuhj004L
QZFCCUFaswp0TugYNbDvHPfCzD0AEYr4DP8ybAVquhxDGyFY5+1pVcfnD1YMJFxz
z7DcEYpm67AKrAY+JekCzN5fLMTOyqV7mReSD3pT6teLjZQJZ+mFfZwX18mgFwsx
muat25OTbWcsYiJNHZtP0XbK/fn1fObTBnCQoXnpgdkptGcpD9Ua1VmrK/rJP0EK
1rW6AtoK2qW4Dh4bWGxLR+QZGFDj3/dFz2kw34Y8HT5n/mgAOdJ177T0u/5wEcDs
SIXrZsQgdPaVuDwCesVZHMgRMqDpT1IBDTgrDUcUKC6uaOGPEcDpBIoRIocTiuG8
brpXqoJpNE68bwQ17QHIYsujA0GZBCuLStoL3Skczqd81O1X4QA0i1BhZbp/GZta
SkgKoDRn+lXhnMQVr8isXtBmUWcbDsCz+yGu3pZI/UwGFl9kassSHa0sj0cgIgG9
QGH2TxA6okTO/V1c3DFN0mkH7fY9DwzPkTEovLRuW2ctC24+V7bMyxAznCjsbfwo
roLt2D0gaSn1R5yMvckGWEZScqUCBR891gYYblhDqD4Fi+nbT9J13dcZwLXM/GS5
/AtSiOALL32tmgDyP9hi/odg0Q/6RK5aCbPjm/CqHmBUQ8Zi2p3lBqOdYa41avVF
cm6m+0yl7xps1Wd3SY537eKmgPseHlqisSxphK0EJqQA0IlUTVYHL+RTulEMJObG
8zY410RuJYiJHpnuephghXUf1tKbhpzHJJs7UCNSEx6tS9JcI4F0+tUCzgQdC+Lk
gLJ+ogqItDMlj9la868NjxJUHS0NqbK1EcR1L4cVSF4PEeDNA9Chux6KA/sVHENG
pBKNPXYugrzDqn5CplVHKKUc6ujrkN1s1ykTAAaidl9oqTDWtTnnVOlt9CHgQ34z
EdeRNQyXEjQlDGR2MjEYaD7DcrWE0XeWKtdFrGPaqTobBstFIB01u+3woYgCGKX2
1n0fDfd3YAZDTOZz2ztb1SVMVYKmB8Zh+SlNBqEtX1KpPvwViJEi/Ef+Hj2laX60
jTAWBN/OX6H43FX/urjbGYIMHTXCYnfSN0CWY+mvD06R2nZb+g+zzSCd4NBNl8Zg
k+EJScLHxSA/3Ho2Cc0h2BITWuwWhxrYfD8WP5D3Zw3zptVJOQPIrzorDFefbvfp
MGP6zbjyOSwRkfYqHdPhXhf+U9BTqznrs4DTUXfKkjqwLJwLlTrniFC3HScN+gls
LRMJedfh+bK7MRIGwnNUHkE9Bwzy5qJ9QRZCfQRP2qhh35O0g6H5Y57qB9vsb37O
qaruBJMr3OndkXmIxGQF/Oj0wg83J4sxlF3LOu5aGuqVxVHAM8OijGeR5wjPYgLC
Tp5ozIxD+YzrZy47I6NMzhGzD7OzxMJOszKO+cl5YYYNVJUQO50ZAxzVMXHKw0/l
RyL/wnKGrXStEZ1MWKg79Yt5dK6QRNHEIPHYfipy8ODaAW3cGw0/JErHU/uP2Zvt
1bsnxwRnki0aem6NehLl3PLCcD4wrVZLTZnwCm/rwZKzYdeHhH1UXNC2NKPQhVKv
LMc98T4LO90TDbdtrLQ396/lq+f1+5Gvk7xf02Jk0OKoi+nmS8NRXu8DhaO+8rVn
0a9fDNDSjICOHLvYR6GfdlsLFi6/XT/fLiM3W2yJzfASJ1hA4V506SKwYTAeTSB3
LvgeqqfbaLYtv3L73os3DBsEZcIyUiZ9Fna0bMopuTCjWgH2Qt5LS1F0yc+E/9lN
+ogKngPkJEjZu6mElMMKdKw+LwCH8Ny5moWD6mOgTtqQS8x6JRQsRXeC0VnMe2o2
kmGjaAOZ6RKqBDipu2j4yMI8Eu8dHrnn/p8UH4IS3amPc2riQWs27BpnJ16T3Lim
Q4N6fAqyc5e35GoygS1ryk8HKGBJuYenap0PyYcLuPohYs5xnDCFIAmO2xyNeoBG
dgH05h1frG7WeMMmnyGNokM0uzP5urjZwsvKznsIew4UrbzbHRSWOHAfTlqQEhT3
AHmbNuNr+0WDYtZTsWQG6zfyeXsnlWaHuTIpMkB4d0Q+5XhLpt5Vq8vYMt8gtJD8
quoUdnaMzb14Bveh3TOg9jze5bLXf6z1RBFXBaRBbTbPq56jYFc8QsIXoMSixIWI
CnJbcx/y2tnvxEuu1KveL6eaU60xb3CtEiOLv0BCrsqtantKsjzCJ9liImMhRZiF
xIicAfnUz49Wl2+GmY/6BTCUkct2xHUEyJ/Ouag3nYHpT5BEHcg/451P9GSDVhsw
RqbCCbal/ugML1o9EOYQX/i1sY3w43DIjZ10F4hsFeFg/XzgIGiSmQOEfhCIP0gI
/0nL2aifvATVobsAqkAi4vUNYZZr2VhcUBc/HdFUWKcZDrNyWm6oqU9Qdk3B0j9F
2C6c/Dcwg3PZqBQ9r4Un2dyCnVITAuiDcqK6LS7JW4pUxP46RAwZe9CsVXJqNyL5
P7clx+s7BZWJHGOJBXb8qof6Ae4aHhGpum4zf8CrngGcPJ0Pa0eCZplcpfnH0Gf3
U4PdAC/XenU2juBS3Rs7DynQQt3ioO+DwCrOnVLChtai1lgDCUU0danp9fzx9a07
u7QDBn9n7PeBgCOpJj+lMLf4uhPu71VHbz0Md/xUMoaVLXZtYGPZznVdlvIknO0H
wddJ/EKHSEllJOqLpyj3WPTjUMEYtCtKIUzMR6UudklTJS3w/w3Y61TpOZtnRQbW
UK/OHXBevkS8G5f7ThbkMOFocGwOQaORyxUPcaCS0CaJ1WLN+0+F1/JFeo2KOx/z
k5iyHesLb17F9TxB1q6NIpKEHOfUSm9qamdwjYdkMEvHIAie8MxctfP7hr3pIroA
dQxL06la/yizYLSscT+Th+OlTb6infFx7VzWzxAP9KQ2ckAesnp0Vmej9Cqyw7wP
h3WsVKtM54zuUV4ZlQDgObQExQRUeavszkzZt5ODU/OjlKDrAIhT8Tcz3o2kegQx
McxJ5H/7ju9mCetYm4hdU4UGkEw513jY9KD53+Vn1abpbDKcrnHFjzI37vVEyWSb
+LOw2Jo4jTra10/O9VAsh0n8d6GOXNavPULA+1vOouDRGYcpMrXzQRpXHYsSiJrq
YXD6oWkDwPGYx00j08xaznHGhIU8dqbi+Pj4OS+ZMAt0bPAOkLUMC/vy6npr7pHA
9GDqVxXKkqwv6X+Gi+IBVDEvFD2Q+ORQrYEopFk2yKqNYWYVVtgiR+Zp642BUs49
H9DrBzPQ2B9ZJwG23wIic+yi8Y6jMoUCKyt+pxHNDNZ8RzugSMqy5K49H/bIxZc9
rGyMoVf6ufy+UA2kG638WhIMkkJKMHOpbkoZYP3BUioygwbiaPUpHb1c3sPuLFFr
uzpUkJws7NglmzwyxHO3O8jkAp+TrgBlNC3cDOuSsSVSNXv/f5XVm23WnhKiUxP3
outocpMl/gQwmxTs88A85ndS7tBZWS3GP0sjJX+3pEZiqY4RMpxmALnhtFCn5ERd
a8Hre2Eu+W8I4+Ld5ftoyCPQY65d8g7oiIZJGUcGds09vIk4rvSFRhqlD5gzQha9
QS9nV/QMt4MDeBfesFY/He7qtG8qUbLppyTy+p5FHrEMNT5SVVoGnoh8KTqBlBKi
w4OwZJ89kKD9WAARRyPBnQwK4yo6BkTte0VtHaYjkameO86QLM0kzALnXKfaGWgT
qz1ZmwsjoT9aYZDn/Rq5NNz0yOlGU3Czqk6UNHj9rV5gqlzdtLi5czcNl0E1i2nW
RnYsQ0Gqt1yKGMKe/PiO5HTBVozkSKRTsGVyG7Rox9vCYHc96/61fupEOhmkTV8s
2e41cBjEylWJI4/T4hhA9lJQUPFR6/gadtmabkdrnaC7YJSMvunvom0F3Hj38tI8
rUg7cI9AAeaxJBQblo6RrVCbBB3dWgLaQbfO+aYd4pNyH1SAojlax2BeurEMlWr7
MLOFsKYC1fakzAWJIhOGRLz/YFfV0gMAkROViqGsgKFXRavFNSt1bjiDEGu3E9Y0
863niShlp4iNTN11XhYJ5tCG+HdfmcBk/KXQObGeIhnQAF89CdoKHPoXZXSBwlW6
QbZVw0Zd/9pdYGQAwZjHYhdeaY4aop14DQmJOyVhgIwA+MSG1DCfKuX7bxSpoGSJ
0CnoOj2D9Eed1dwFcgZvhvH8h8nbc+9gdnmjk43VXxOBFPkv9J7+0FvWXPwmfEgD
MWqwhX/vrgCuhogLrJ572ktt7bHcMhBSmREgC66+7Y9pksRwosOsH1G8FeN9xoVW
PG+3VUWo9tSU8tCNO9jeHcxR1lZlIa7ZZtQnzkCPMWG5T6nw46uijHAKif2DpUBd
xqmPH6/R2H5IAf3xXIcbdh8Z/fl5Sf/1gxWjGZ07bxdH7wVYb82VRbCDhQU1Hc3T
xNgc/rDwNUBE9aX3FXxyKqL9LgKj5Og4hALvi2Wabk412BhutU7aSiYWZFGx6hkm
ELQdkCY2I/hJI3eQ9NTVKONs2ILQV8eisEUyqjT1m+ixPQqRFiPYIynisWEkgLHq
xZtTWF45gDGHHUtL32Z9FaSYp9Vr5lJj4j9Q987E9GQj70KYhorc+VqB5UAF+RdE
vRDFCzwIBiMnQBsaqSK+mOEh3GeJTQ1qOYQOkqWUu50LnouaTLpn6wcepq2JXLpC
WhEnfQ+VRKkhK3dS/pixkUOEgRpPLuhRTfc+YPt+2U1RiPLuqaFSG6GDNWh2zZ85
AXRrg75+zreC/FzRiVKe7BW2IIPv1gaF6nCnQ1b2I1OvFiFQdNk/jJyFt7lzT8Ne
V5T6tFmB2gVdhPCi6XTJOeay7yj7XnMGV9lj3x29u4G0O/Z421wva+81KXBlpuJw
eie8Fz385CI6v6K95K/RmyI4sTlufmxgcKfYa+/38ASyhAJ7jz1FuHUJGUVP/8bM
qA+L3Cf+nnIj1WRZglX8j8wKnla8Zv7wG49mqdVKSABx5fj/rQGUIzwZDtpACv26
6MuGRHBtETiV04jivSjTCNkPHjhMiV/cndMYHpJrGI8zg9rGmAD8+ekQrswgJd55
pMQ5J90NWREZH3C7b9SDZ8skvQBtvlyVJnYGwgITMTF6CMcmnOhvQqKTIxf1GsBJ
KeyPxNSwfgdPMeHPcDSvFroukfI9DTrHsaXkEX5ncaCBv4ujspaUX56oYP8pDF8u
1ybG6Ed9wLRNJ6dpgDeUDGq3Ri58D0ktSKWXfOV6/KbVOdSgIuOW443knScFOYo8
xKZEKse3w8yqi0DFDOPLXnIME9e3xrZVhyNeFBxN+4dDVhn0RdDCU+A2fKHGxCxi
mDCnLxH7T6dCys7aDmhxzSinDn6nKAo/bXtnal9C12fWIcnbBzqpn3+OeFPcZlDh
bHHpM/EezUz4UeWiAGWhMk/796UuSou6piCV700/6flnAo+isk8Se7nnT37V0N1/
Xr9BsY7Efwy4+3E8fVTC7IlxF5619MLCUYCFH0fhMmlGoLWSvmuZon6J2FW4WFkU
qkTIub7XHPahvenUypLWxDkufddzDLEGpZ//64QJAK0RhizICfjAwjw1Xx8IdYph
aqhp50pE0TF29bhYH8IF78O81VZ1P+FzupWvRrfn9/S+sXg6z2LscoZ24+pL8nao
jWtT3qIs96FWGFodNG6LDghWMJl3eoxCWS1heABaYN4Kf3MI8KMLDwbz2b+dl+XO
gb38zTLMrqJ9rvXm1uQgyjQFHxHhMDHsGrfUXhHLZ/kUlKAiTYbxEUXossyDEpxF
fW6g9NvOgqU0ZkgzAKAB3CRfNzkw1hfYgy/Ibu5PAHKo4knjADqg0TEvyzal6uF2
35d6MEsJe5xsit7OeX+t4C9NtCv07gSJmQZnDLT8h71TKv+Y3vd63QDkF3nK+s9B
hU+a94rOu1+LuhMrBF4Ci2+PDoBc2efOt0GjMbJMG/f4PP6Ix2dq/vb7EFY4VzKw
DLVq+unfGzMwdFNdYo1pwFCTqP5gQ7Gmt4h8a2Q9oNgQ4AoK0m/XIfXcz2b40956
+iFfPAFuO+zAf7rOp02vKtplZunaiXsN5rlA91HGUmiNuBpk7vs5lqdEx2PojQuk
J5YPYTFZs+pHB5ogOKTgE8c7isxlHoEGrqAaVGNnK8vqWNRpbUgGcrP2267DVQJe
jzKIeZ0ED/HJEpRR4qYhLA1yrdza/aKYaBVv+CzLWYQTOAp7Rn0Ue/A/ZO/pcnWo
sAfi52IRfKCQgZEYAHuvjvwhWSlQxQO0kUfI4OTmFLl1f6N7clzpy04cAERwg+ZT
fRqd2I5Lh/q8kcNOq37Qp6K9hAYRsMGAf3l33xDc9EyoGmRAReorzr8c17RULcR9
oyPuHM9Za7LFYTXXezbJEP11EktNsUMBS93QDdP0Zi9A23S3yR+4obLcXQ8Hm3JM
PBsjMvR0Drl1cyjXv5lwF9KKQ7ckuAYDi3yMG2V8G+AgCBcmBSih+19DP1uBTLLO
dMSmTVc0EgV8n878dp1p18KQJ4xJa2N+eC2Slj0BGwJPwYaLsoWuib99FPFX0KkN
eve/TXqXt/6m6aO/lhSrGCyNdfUNynYKVcTmfcvn6eSEiUVcgINQx56JZQfHexzm
OEi2fndlKQIJRyK2qawwEVS0nQP9DiENXb6yPjVgb+3siN1xs437/IMLgudgZafn
eK65eoKRVDZeajDlkvUQM9TopaxQ2rNvJUr+YBB0ymh5HVrhgOYiizmIr0Ik0mJZ
DaOlq2qYFshpgZQ62I7J5QGgM/nN8UCwxpHEpJtydCucHPIzgh2S8b+h4fiH0UUP
kE3s8wj0gzEUAk7OkH6XPYiFPOVahExNV2zZteql2ce/MFavKqhegxlaKo5OAKKh
Z9mOhSqkhgDt8dYdYWMmKTed+hPhXKQWY1nDRaHIlTkldtsAfBhA7v1si+GYRypv
bTBSed/gTMUW+Xw/9ho5MW7IvbSkxDBc9Ztolva6gvB0OZRUuLPbZtTcaRHCVXzg
B2Pp5qt8u4c+gmFKK5E/yTJUx7voXZ8hQEd7pqE5VyrNVw7thytCnslk+/kQcL3a
z+iwsqgcXGOVY3Bt6QL2rCcBszZlkfiBc2PZbLzfd2xgdxX/DAbi0G1D85+DjA3d
ju/P5XUCptzgvtYTlWnEQpUX7hbdBnb80RSS9EZwf06ZZUX2D2BNJ+wDn0P9iR17
85rnRAHIEdXbQNOOV/Gkmd0t64HXXA48m3RTpoDT9AzuHPnSZzJyMHQAbgpZSW67
KBb4REI5lusP/m8xWoSLnQRAihoH7kPFStXCfGkvSErkovfTe6oDFa1EZXWiS2dS
aWEbdHIe0u+qkNqwgUFlbEUQ/hDJI44Yo39i6Pla8rPQ70MOqm4GNtGlnKDSCXsH
BbQfVICpQCwtyhiMr4cv2Oi8o7TByCrHsFgabQx+wjR+SyOlVaZLbGmtoLJUBl7w
qLa80RIRBnR4b8vcuQdbuylKKVRBf66Pi0kz2cnalraq4PHdpXLZbdAvqnzc3gE6
YcaLerpHhQfe39nu0ta6VpdK1FIDDIHT838gUUW8lSLh9mLR/ER8s6m59GIUBRoK
F1hlKhRwYyM1Znq81D7nPkfelT9wFFNt5xc4xNyMILAddAxAn6qq+zZALd8F0Jyq
78P7hvw86rfTHDbflq2TJGboFrh44xUAKkmsT5JDfcfjyS/m1iT8wanMokCEwQxi
Cwo4YWYQbViE/Pi5p1qW6PYdUE+amHopni1Gc3ky1PwhbqpcNN418WoZbTBr7Cia
x8qMMJuP3hJr+y3/LSTMY4fnaGVd273v0kPTml/27Ehb0yEvsdqnu0ZRxDgPKgcg
suqUucvU5VMy6/0K/3X8/lP1w75oTwN4jDbVCM4UBjyQP1k6/rzou6wG48PdyFsc
LC7mZrtFKXnxqJ1J0Puwk7KcWje2mwlHIGtabtiZDSYvk/+jh00XNbI6M0TN7OLt
sXR6duikwQ4oyvI+ytDcQcoWctKQ/X0JofOLYh4lwooHiOr6+Y6umvXplWyG9MgS
rRWbJLVvvK+qJIXp6Jf4rrayih2TofU+BEKiKKKgD/fuqu1jTnG3Tsx3igwPdr0x
Fw85tukf0grkC6pxaLcqwHiQxALyAQv68xplCfTr2CKakY/4rzaJkX+ezBmL686d
Ik6Qc58wMkT2cBVZsEC++cuomEhZ0UrBx4G290hp68xLbwtVjQJECoqM3bqBGiOj
VSsmaOsD3vnnJExGpKSb2px2ju738BAU3rk+Ir+gjGBRhJY12POh3qS0fajO6tDI
bPNQS85UBF8ih5wLutbMCW5ncYVbWXLHgK4DutcfMwZDfeiIJ+fAO99mLUGZL+r/
MsIMMy9lrY/vogZlNwItbbGIVhkpcAhwq04a4/Ant4Yrxb0TDlMgTESLet+Kspsh
SMW46wE5aeUFjO+SBlYJ/uNF88490y83SNEsDV8ZRy1q/qdxwARqjSDkmlvB9LXT
FZ72e+3Tf4iHb73bKIhnvh94N015uXzadC3gPOssjGwHQ8irt5jzrP/saEPquz+M
Cw6kF4pr5bHeblhSL4eiaZzThDFnn5i+vc4NZnnkHHa7lSs/rKFj4SmyOpw5WeuV
XV6gnC2yUEujaHCAOG9kjXVuSL/hwmhSI889fAOGyD4KiwkLFYWYT/umW16sfW2/
krob8yOkg1exjFR8kv+mqDhSGXY0hqJ7+CuOOSByFiSKbs2xEVyhKC+JSBSWrPZB
Gxe2IarBaBT+BdX98zdAflBV1C8Yvt26Ehl8DO5h1+DWCi8l3ILQYNNcLSOT4nCJ
8aAKhOWkKCMKBPFYHPgDmK2tALXJTHXb7VoudhZYFLuPCkeYd0FhfvVsPYH4GBnc
9hdnHeXhQ37bNtkW44DzLUs6uI+f4HegQilZBsGb5b0MKNA6xhPUCPg8D9micUUG
0oMZ3ACEdW+avPL+N4jGAXhJCJEXYcpA4oUbv0AhpkpFaLFkTYYKhe7N95QuiSGh
GFMqGjTpjngw5rBTeGfa24MmoUBLoVRuE0bxBn9fZa4m/htyBYI2KooRKF1jrFPp
A/B+YQWTQpxCk1X0nRlkHm0HXGGYb2uR3DBvvj+bbRWuBq6X05QLeQ94HyHPFysn
L6Wi5kTkXwiXWsq/jeBuzYprcfvBw5/PKfUqRMehytlevd2mOEoKNpo2iERPTlrp
QHjo+70JI9siCdBM0wWe3/VaC1pg80J4+E0hl2msi2LEYG1bT7oxPb0kzg9neIUh
oBa3W1K0A0TA7QclGG30RhIm+pEGSSNOjLEPPX3opvGJub3ZDRua8XrJeqys1xg2
mwKbei5z0HpHwdK6HMjmtu13Nq3xYO3p1/0SZXvNXQCH9FPHnQDJaEpqj8l34RLQ
v1WiORdx7QWCri5bOnRy6YdKd7055hJRNVB6aAq0TUg9VJyXELRtiBcu+69Jkyfs
Sdx++Ibi+uE/cQ2ReZY3GDUsct+PsEsUarNVLGa0BIqus5JVA9gHAcZht0uj2sRO
vXOHKTE0Ws7/v21SkJtxmOC2r/DFcS7H2nU6WXobOE+2PwZQUeaUbP8PPdKQYg5x
3eZQy0AvYl1W0TQCy/nhKVy2CBjWMSLv6IKpllkUD6G65JVcB4JGsE48QJJ2C80u
/fPukF+tOlo7/GiTe3WuQq/7b9KWFBOUnqFcA5uzAIfpSpMt5TkutpdcDqMXZPe8
e5EOITED2CCfYl3gQPH05fQDQmZo1tHiptBbgHwf0zzeTG92YZEdTPsLJvEerjiy
7gu0maUn3uE1RhSMXISXvH8YmC4n0XPze88N6gOb5Tsw+zEMgWdbU3mMoB1RK4kv
xXJeoTyHjtSDOeowW3jrj02LeODpmGw2h4UfCZisR6bnBbmYzb/0DLNdlCCaKVxo
sKuVHC+drsiZak125UIS7Q9eiMv5zghkOqpDfNkmrY5wnAgwNmMB4BHqCWtX9ixt
6KWu1SNpfDHcu2Mfo/S8Qdb9QHBY94Uj/tgqBGW6uboVEx3/ZubTsE4WjnEX+GSI
950eFXFR6V9lEvtKRvbkG4xzn7rTLZeQbjiLQHEm6g25Zb56dhzAVvdAFVC5kEba
kSaUGMUsebakSvWclNz4gFAFUrsIBCd0ckE+vSG462XpiQhKCXvDX6Tk9KVNRndk
82yncrC+zMV8n7ry+/qLhdciTFehjK5cKjsprKXYd0fqhc+6+fV5ICAm0MEaNdBg
bYPKZpd/2AiGm2ufzJQf2sV1CL1WPNy6eFWfC9UXeLDo3yWCwupGtFnouDaFtjwy
kn7y/iKb944xs0YRI4eHbutEzJ/AyXW7OnNtFX0LC4hJ5bbq9yy1fz/26sfDBUmx
zneXPubM7utiWcAtvZ1aOy6ryudNPp3OnugypFnV923Yh4KStGHF3RyuljWawhl4
i4ag0pdLRkeoCTQa/phC3LOmd2balymrUxnl7wR78BSE5m8Gi0lxL0QVVrFPVtme
OqF3qp5POuDq7HqlPJDG7oS/qCBYeX144WJ++jqv6AMsDVdMB7o2wGzGRM6qyM+i
gd02y+ZhnzjhalRuVhlB4w6fEykFWDrqEzvnP56uviHa9e7mqyf0ipT40NcEXRyG
QhAk5BLgiSfAvMiTQWnbKa3ubqxPmLFVbyo6sQza/UXV6evFPMBrlaDBazQQoZU8
HgPnazhHt0sNll8xk/WMbPdC0FcPuV8u3y962shEKrOxZTs+ZiwfhowfBCjBHUNq
B8nWuzb1kWD9KP2wGRCeJuNXG8Ld1EJtiEgZWDczGbQOPMgDU5DpxkwzG8sYNrap
W9Nfys+BmQOpq5UGo8j2GbJ8UWu1KOOo4soJAHDswslmdIz+sKz7zZ4JM0/ejpQA
3kZUqZkWkm2cnSNDY5cbRzSFUVdGYEtMc34yJdsNxchbsx1kokpzXchZmT2TyVHF
/l87wZZM4O1XijBTms72iI4gBUklXut0DWf25KKlNElq5EJXdTPoVXMY5s8GwR16
35n3/r5YftOTBbQhoP4xvufpM8rVa/CaScbNPhmmdPa/87bckcJR69n7shQU1o0i
KIPm8vfPAjFr28P7bxkJmVRM2E1u2E21OooWM3BxahuVOCgMEY+ZM2EaACVEPi1D
jL0zC0MEtcC4KakpXOPxuDZ9oLNJCORNpPUxH0bNCHKFZdcMWqabn0Shb3AujlZc
kt5NmxN5VhBgaOlIkJd5fXWUi4gaedJ9lIFZjfeNfKbdQPfu+vYIjy0bITJtt+Rz
Wy22xZJoH2vykNBr6zVb3PXN/Pe7XiQE9J0E/HvHo4QhqNqi366Uq41iYdX90/qD
U1lwTYH4CmuFY4b2Iln3VKv36RP9TH0fe6RFSdMqbXW5TBcimiGWmT2PJpJHImsn
s5wfIcAytVZRE3MBTiKUrQMJ6g8RI7ST1pzM/IZRWYZxxNmqNLe/Dx74vekdrwB5
K3Ia7JSgDBAQsQAU81HyxsmQZMgEbttWgQ5CgYUw1IIdPqkfy8wzyfuJBRqJ4e/i
9yUjsWR3x4jUzwUgw01zTeCeT//SQogcAmutFoyB6MOnrC5LmzVQPpWQEEhKxcVh
gdQ9mBV1f/V/7fCuqdhMIiYmp1fCV8Y7sdpCbXFPxtcUIyJrj6vsT5Ep3gPbW/2c
EjgvF/dbEsIJJFmQAe6bIwYO2P6q3AnF1tfG1f89iSj5USAY3moiZ72BGbp26bO1
72pDKHVcOC0FgbltJ9uofeEimi2v34IkwVcZAfODGB/uRDbA8FMtGCE7EQq88x3D
qDmtTIMNs0hitSPoLRdV2Z3dyOLkNuFepDHi5FJXtUG7xD0DYPl1N6IvQvabqrkN
QlIC0+4ztUTqUFZe25W4+zjEGAkMbt80ixtpGb9gXFIPr7nCn/vErB2fZmXql/0j
TWfLDbKp/b+kABEroqz5/YxwguWQ0QFA0ehHGSXUfjR08w42KgDJ4pvFE5kP/kIi
QhkY2X2K3R6jgOolRRqGUIO9Zj0OWZVBS6nS5qwHkNpKBG6kGu16lK15bCE7mIvR
sAmo1bQx2UgH49Hj5RAkV5zJItSe3snDkMIEMlRLT6OpGpmoMSc5owCLUa5hs1iA
1R8e/uQqP2G/xAtzk+SzimRJVTFRpIzaCdKhntStV9kKjuRQw9Y4aHnX9w9OIhIR
Bd1tJou39j0YYTl262h8XUwXx8SYp1s6vPzb5uS+slaLtAorIHuNCTMHXnhrQDZp
3gwIYV3XhVVuKkzldLqhf1uHKrH3qVgVW0+rxvPr+lDolnuUulAWQOMg90QUU1mc
uwjIBh39MVwTYNUh4C0eNkbHyt0uSnYdCnIvkTaCz9hyFZ9KrmFcYHRybj6HCWJT
8u5Cztb8N9VnQJFRtzfL+mWHncfaSMZsx9T92RqpaJ46pyCCwfEQ6KXXmdxBbb4m
kOjhCNovhAlNwjNLA8Cgv6jCIJqMxNdaiiAl5Vtrc1KW/d2xn/KzO6tIxQwcSz+0
s9JjNQH4u7eGxW3CkixvYOD8QsVz6QJmy/5ezWXmRx9fVw+YhFqZNW6rs3rQiImJ
lfAQAxLiey7Zi1SWwnZvGgVqyAiavl/aJexd4dTCRO51ACezWu21IrFcBjr9a5+A
pWh4cWZXQdteqAG2HziwFy9EBzYCUa4RpsxR36dw9kvuilvJpKgAlPd73jo6WBZk
kRsN0fn0Bc+cWJILV6hkkL1aO2aN0hNv8WaYC+DnHsOblpn0SUeTjyN3UMlP/KmG
PvvnFbVUCi3TdjY3XBFlJFuA82SxsuVMWjHYidGdSYQmnXTKZe6asaL25PUMlyCm
8KBSobDW2nNfn1cv9HIDKjANY90GQYLvSZdfeTx5q7eueWLfNTL/VyQuvnlU5aEW
/uBBypa9ujyQwNsRD1urF2fvjnnvE2TChXmPYlNn4/ODffXneQ4t03NyhI4ZXtWF
IpjWe/23JXmB9+mAghUHiCXDG9lpQgZrJbK/jiVdgsPLH7/v7Y855C38hvt8UAib
ptniOqR8dxBWjQiGdUTESu39Ur943c5FVvm08JBF1bYeEZ4dnZ7BsWcsO4WnapXF
p2GFU8WlxL/11hf+bj0wmvVfbtQkIhCuKZf8d3fVazoUQCPivlOhxZj1dBmrwDbP
ogekKXSgAb30uIVYXR3/EzMXC0BAo+/3L89FBnqJ5At845z9HwkHn1REZiXMxK+f
Wbuk2da5zRj0fs8S3DLGEliSzIJDvKnal268DqHjZR4uOJ5gxqZTgwin4vcrJBhi
S/nxJ2YKCjIURyI8hb5ypKFCamqUJW1lYDCDKPDPOc5P94CbDPLyyl9AqC17Wtb+
rIhkKGhlsFXzb1TcTxkUaJWgkFQZtfoO28pTmKFgrgEj+1FUtWGX4hvwWgWLbm+e
hhBPMBQR+A00KDnwFyvQ6fIVfqnoPow/20H8o2weHkTFd0wgy0zVP0hDABO1VnN1
5OvOTF8Guh+RBOxbeJDVhXTGiCTyBSt/V3ZhhBhmCe1pSVQPgiVHGJPpp49vPFw3
gQ2nkNe/FCBsLIQizdjzQToSdGvXTKlAFo88WM+LuJG8YW7oqPpS3KzI4SfmdDDR
jVEttqrKBKtK0Tri7urY0k+6ab8CO3+7YLzimo4V+p7fd3gyy8sPSUlUomLlD2/n
5RX6ePVrA0WJkKSL/DEWJT9t5oLqWxHavgcObjfsxO1xJmqgvLgLrI7fXKQMPUDM
yvXYmV+S3LsKlfKjNH1pZs1djC+w4akMi1Ao1K7uXXfU3Ax8aw9ovqmidjdjPP2c
BxX5OGDdNHFuyFLKQlaaIhPHspvwYFnHq8dg0fO4TcCe0Ll2ez6HsX8OHZ+VgiT9
qMM159rWzrgKVrQle9UBnbghVgCwb4DlJPVCtgPGGgEd5ygVk63PFmbrFB4eLot3
iV0bZRnuBGrK9/D0tqEnKcC7Ry38HA5riJ91TqDG/TCDmbHcQhQzDOvlBzZ8C/eh
IN0XMMm/j8jg1qTDYA8awlac71NE4fUQV//AqFmPnWNiZ2kVNJ9tQLlSzhl/i/OB
H5iyYAA9/40CCu6LR26e1wn3fyjd9mgq2lMWSDSkacAVUywa0KMY2h0dKVIxQIUV
pNsbctVCZzpcUyico6oAVrB0jT1FOlD/h2NHxDl7jpPVhPI552CD+X5tGcnaqsNs
zSl4bvaH9Gc/c/915EAyYXh4Cs5rKt9BpLjcNenvs2ya9pm1vU4NmOxHqyrwv9ci
UHtNBBQeBqGvqf1KvGmPGLnshlxcD2Hy6v8xKWwv9cvyy2KwQkHzNjqATKVuvLlu
i92DY4TKfVT9Xq4FERuy+Fk5bulRHBrnef6jaZljacOVgk/Oay01qipPQujzQLwO
kvssExfZZkNvJTX9gEQh2CSzFfn05SXdozaXhtfu8wrrZnoTlfJty+FUX9mB4gGZ
etarvEcQMtvg9P26Q0FfyDk4oJLss/Gp4vJXaxLNVT8A3iR1n7UaFx8qTftPUWSd
P9ca62KwRspvssku+BPEmLvSHzZiRXP8YevRBXO18YyHCVNXv85C+DH7x/c+hrM/
ShYfpsrXHEhmvrf3FSZDXUrGHwUayQu4E8cIicNfs2ANPI5AJJgyDMoaGC+S6Vnb
KoX22ZeqSHRv8StJ+jliF8aEqVW07PgxtPCr2mjXv5NcLPxsjt8cJBOjKFt4tY5M
EkZdWmLttMROxYocHIJM6FMKo0k7J1HWsW/ur9H6BOm0GPev6+fnChI05TCqrI7V
twSeDWSEVSFdlrNFWo27Q6Hc8TZWBx61yzKMtxw6lFPtzFpz1p6Idm+Ab6i9AXcu
YvErqukVFh/T+Pq+p1Z6NhGZuKMbcyUzlgIKT2ablVOOVxm7DEpEUA+NPGmKnApc
QqQQrAKB+lUIToE0ZURnMayQ5q3rKAs3PcZORP/XEVCTbn6pHQFVqBF4UcZmNv78
4brZ/MBODtgIqhtUSoXTf8FqWRQNEJHc2sxiWiipUdP+7CHXTwlJMZTBgBFJ9rwT
73MNUxeerfT5wHfOCWF+CeDbLDYeBqXc81nb8CT0CGYJ9Q07sxdDQ3rgNpWfIIIW
eci5aanMUNUm7dF7Fn0V4Tn+uRXMNvxjsoKbt6rL8JkL2i4MyOevDQCplJUkjPy4
C7hthHAIpwMA0OiYZayBGwr4aX9Bostf9UqSOxPVRTvuiY4VqYsBpCN68kpomTUc
qW7aHk+GayUKiD/J0sTNLD7f9HokpACuocFAxdoZucCY2uQ7yUQGJ+SzOvdOKQ22
78n9kJ99aSY1om8Qcfwib1u8ZnQGbHG/gh5WVTjLEv5Hbi8P2E/fhnl2OWitXCPU
lhDDPkN7A6QoJV9YngpYfagdVeUOBhoUkPoccx69x5haU8uyndwvLxHlT/BXoEkW
nT9HUIMLTQVSG9GkbKfL6yiGAJ+td7BQgEAdUR+oSqqN1kMnkXJsR0z3HuQO9ApU
vRBzxD/SO+mHqkGAXJTEOQTxQ7qke2StZbeS/7a5WMDOcQL/exmRAQwG9cSafPF/
SUDdKIKs1wXF47mo2Y8jUwUFjnp6btt16H644nWd/0brPJGbkIlFIAqvMsofMTjD
G3Rumw36CdXwFG5UhqoXF8n5L8FLL04GnUCJs0ypwb7FWJV5roWulGjv03pg88Ji
jAOkdmEoByDVXxyavB9zu9Y26vpKozMAzzaR8pcT8CH/w/Js6PIciNEKQSKRLpIE
fU/S0zGmKKnMl2SBvITBypQXiRHDUXLUPCGnOPDDU1imPRr4kVFWjZD/yUytB+N0
1K+xirtfqID0YaiOCFdD0pqQa6TupQW/dE7TQX6GKI9I4+CQpxXvV3XOUitFhfVL
DMB0zecgeHuMsoqt7M3e2/NSpkxugDSN8rUggDtantMxSptC8EHxq8OBz2FzuXNm
kldXI8Fc5Adc3oZDDOn76e+qjZYxG7Le7mP6jvoT11yxTtJ31i2T4qGKVBSv2tFP
LTTeQKYzAs9CHKPdILqZmqEkx6vk10Hv/HIrsbOtmkLDfC0nXr40qeNJpXbVHzSL
5q3gofdRTyKUvmby1F7+7639ISfXYrHxkEznEozNRyMHR+9+WrKebQA9LXqnJiEt
RKVrjgrHNytyCIs4qnk7Y/P8dqctBtAP+r5NN+UtfWPupAq8IcLputyCeVfsaXuP
SeA1J1nmsCDh0NI+dNcCvmhkw0sD5f9yOR+2OeN3HK/fFy++kFPOKXUh/bX5jD4N
KydcOm3Mbk4eDQp5y8FYw9NoiRJ+3WlDZhbsW7YEEN5HXLWW2w8WVj3EsqwKPceX
Yg2Pr0mZV++kpPcY5vam0YVvzoVaq5zvxeaZ8YYdAst/4umeG8AJjnGVfGAP7LNe
KEI1avDVnurb2Q1cn5IWkYmNIWo8d0lE+BeVODHr0TzUsJnpuIcFJxwJtMRxWvBF
z6eAMX7NvasmZsagaOvBadAFMAldaCydeCDv7oZ6z8UNQQbCnFQ4zA55G4Usl/mv
n86Y16uEEzhDlUnguWdzZs4+KKf0wpRHZQBtAw61eE2zamE3yIKNKRBw+n91Ba7Q
uTUCKn8SIq6aFrj4fgq5ZZHM0hH8CC96IxMcjGmj0bH5PBLYlpKkIEy8dk8Tc3rF
C69xLjZ77gwAoFuqWauB7Dn9VEpq2qYST9zYf14UIsg4SS2cLbmQdigTPZff6DNL
90r6xA7kMl7jIv03FwHmoqXt4K9W1GReh2b97WsymDFRZoGZAmPZAwr+iGDsB+zr
Gv2G7a8s2zKza2z+bz8eYdkvXxBxWmQrv9hDNMjA06Uz1TGNIF1kWoGPR0F+14hc
tVrA5XA8WnUNF57w5RRnniqAv+aJ7JSUEOrQlUyer9on77xNsrnIBPMPF+83KN2/
wqcM6HEJ7jGnMGJ4UenCt2nXpi1HT1GvyQetu3s8QyILOPKFhnz1uyZy59039Xpo
ThC/S4GGVSRYG6qgjO+Oh4GFUerxJEt8Q+t0hJbYT55CQayA8DXaeuOLfM/ge8xH
yMLnlChz+5W30AnLny6u2iqcOTfEYHyIe89znasFErTkTm9Wg+NRWwXWsb43Rcfj
J86g+JxxE8DzBXpsaeF7xjtTpUIh7a2s5cHyrSCuZ80gaIVoOfNpYw4HEIWbDe5a
39fFdELZqaYmkm23CkOIDUBfxRvpbBt2DVFy00CdZ6VdE1Iq4roQ4uuAuaksOKX/
xUzCdKvq+fA9ZQeGNu0PgskDjr5S9qKlnXixO2ZQJJxuAsSLbeZ5bh8X1TOXonqr
jQw5qCuIFoNj7cID+eU2DQsJnANe9R8cbl8hm6yytr5CwicZqC8GdDByorF7q9Mi
BiMqqFg4mhJHXxJnft8TFleBjMRMo8bMFZW0icXVG5nFXM6NyhTLtUqAEfBrkCmi
tykeDBJhEPDU4i0Y6XRXErV2mqC4r6Pwa2Vg1cmb44lYvh7ETwOdiOCfiJc12kIj
854aEjkK72C37jMiDMIzDneCdJL+/GlC7o/YgYXVIx6npQDKZUgbzN1FP6dExV6b
QrRO4+gRIG/cpmtI36MUyL5UsnvwrX1zsba/EKwSIRgt4KvbpgmGc5csXzbf/kz6
osAJ/RZQL9OjTXo+dQIKen6LRZWnPbtC3+wEM0O9MNNd/XfxKZq7GHV2yRf9a6V5
PYVunzrtxtNEOYlURMwEiQhIA7OUoANSIfdVWaohDT278xQK+PxAGl+xfuCauX0j
YNV1oQcKxIcqW2cOezNxDkBPtnUj0FZrqB1l03DNOYaIfbr4mZs+hyQH9tIM3Gdq
mqAAm8m8fgJqmow3inZhyckEWW/Mj2PXRD7qfLqlgiihH5jtNcFNz/s+Ih6WuZW3
WCgJ76853eN6+TDBf5JreUY8h9I4JUKvNBYKiGrsL/3v+NEWqm22+ePSlyDE5RFk
HupDo7U3piOvfjXbGXzGRMAE0ah25D97K/4/EWWMc7Ud8MsVT+98O2ekakZgfhPD
BeMB+b170xnmjQ+qHtC+G3x52CkRV2tsBwAgGs2pSN8m77pwuR3D5QjFr+yXvylQ
d825kR4CHZrgTs5gaijTIM/h6aEIviuNHtZ10jO4NF0pYrZ6zz3VzljaP8PTia3V
9JX2ed5xl09d37gOpLaqeY+wHIeqc+hIZFRFpzpeoJGGvOEC95oV77L+JcKWnhhe
uyN5EESkrsruHPcHVVJts/tMrcqAYlUdZteClcKSED3A9n7OgfxhERePP1rkXQV0
46xEQqEdlxoXRz4GbIQsKExBU+qqzia0EgOZb5yrkhCWq1wOnk7mIapu4Iftfrna
d3tSoqYQK57g23XZlmbZa9FU4yecFcnKQ7x3Q1E5JksKhxw01Qa0WWqKaBzujsnM
vN2RQuR5wcToqLe479lDBb7kgye4nojcxI1PnuxhDuu/E5PsABkIC9lZAVBeaOfs
wQRnyczD1b35Np1vYAco83IG9V5fnucWzoFtjOERAiPBF7bzy76O+ys6k3Mh8bTd
/uQrvKIpzb7Prk9wk0e/N/kOnNs6hFlV1pk8B3cRUuz7ebSJajn290C2h+yg2cpe
Vvrz+bbqY5GX2YwOL3rQQ67KQn6ydf/5y2Fl3wcbcrUH0LLIWe0Mi4MBEqI4KB0W
j0ckUNLsAoz0I2taOm7rzjOP37MPFPGVlL7vCabg/DN1bd6ZWiKCs9w48YnIKZEu
0lSac7J2o2jTZoJ7MpRuRwfTKBclDsyBNCqrsZR2U0aC0R+Jz7P/4CazF85OCzxy
u6iN1cza0nPglJxtK7DIwlYO5bmOtGZSGPOOmiMWCjdofLxj2pA/Xlitp8+e+GRJ
3rEvy3Ug6q53dTx2n8Z/TVgQDWltmqrQFnyvRs4giSFHw4ZWdjWC977x/mNvaTBi
yF4HNOJCmBeYwgzpbBD2XTVh67Cx7uXyPUgKWbcMWZLdrN9U/Ug0GYCotQ0/MIfb
nVNEjRZu1LR5uYVy/JpOARwZqjdiDsDZXNpqrbomEefn/G2gNs6piYHhz2/xOhYh
oK3MT3vWvmXHXkZf7DMJSEdtI3yV9YZYyZZeItQmbmdmsjTEIQK+pb2pIua4wLYM
TptTDsHnIvDRKSsr6zxfN2HplMMTaKeXaAP8DuiPR6SsVfage5UAFne9KXVgowAF
CpAJj7Rh/eBDPgE2v3s07QNE9/zZM9fSX0szjRwDdcY1W1mhTVLoc7JtKN2FlvYD
oX8FI3926Nx7VwT3CueKVdBywCgilXpgYASOoU+xPjMvfNO1ZTksVrV7vCVXGcUa
QAmdNW2er17orbObDQ/CSfo68pkxkIK8qPotH1HUCyYZ7N2m2QJyzvGCo63gkXDd
j4dHTsO5F8eu9HDQieoS8ln+bFcgIZDfFUvkVAs0LhCkuSQWQWv3fEyBjfH+I0w6
z+Inj47Juv7y12h4io/ROKCXF2lXHMdaws2oE43j57l4V8cuGVU+35gjVLs639Ka
Flx3K+kEGOVREE6xohnqXJ0MW8yo5lg07pDZYxYnChFY96DfpD3VoJFeNXkMCjCy
YFImIaYG16njCoWfEPzwViVWxTmo3T0IszIm8EgC1sdH7rxRVid0DqYqj2280u3I
5gA79alT72+i3aEWQnK81n91vzIES1PgIDOkYKU9heh90z3bM17LPGaz56Utu8Xg
MYNDdoGxbAYy6rHlFlz6FHpZ7EZ6Q/OlNC+YSp7AwCImOOckzQYT6GgAZOFJ4M/b
EgmVwHmQhXQDOA1K21waTjKlzHzs9rbZqwdEhvPO3BJzqEphGTUAeT2htjCLyDKT
mx1ZzTNiMYxTn3R02wwrUlJYLBsGp8tFUzBmovcNwRKnBI1I6uzgWBy2CsucUV6q
7pqrml7i4+txOU5xDHu5TbympPN5/iVsSkCmvB2/jQszfLhHIoBpb3d3PoDD74Rw
pZWiwPGm9lEb4okeEQF/H4iW9YI+OWVmnDtKRjrq/FXH5RURajA00Vv27K8ns006
oU8bNjGVf2OT9Qu8kl/V7td6AD011mnLYig/TZLuRbT5fWxGVSR6Dl1r2eFSpF+c
WjguGW/Yifh2lWTFV3hJCOs4UwO04btFpNcM9W7tgVtW+2RzRc4Cvv0TTQPjtBKp
Myt3G5BdvojoBpfVivM1eeTxGzHKqTu5OJFDhBIncg/AJ1iRyNchOSu6jVsMqZ+H
F2AGrU4QnfjuwivEuqSvX/VAFVbtLF5ub+Fp2o4OuIognO5PXrYhZaZQ+nSHJsXk
ZtsPO2GYgxE/7LgolPFrR+mii0ASbRKPlw50m5izr/2q5UFQSl7iPMoUMWwEtAon
r5OxjExf3X6dy0ROpB45OEqmYxsE3mhaueWiG/KVmvLt1lpUErRN8cx962RDQrHA
MQyo8vRQ9uquoNZ71dTuebCxrnFJ1TfGPBxzcmAR28WE8+6r5AcdsZyxqDD3GQlY
GQEW2sVh9xmQebOOE6LRIMPJTB7ecnZaUuZBA8tQToycR09YFaX0jAydf9CicOuY
dktLLgUTMkYgDRKP6SSYtZ3tAI8uF/hY9MhXjxWqdXGETMloGojaPNpqG74Ficxz
G/yKLiYxbTkzaxR2im6m4h4Tuz17vGnyCFPrZsYCTsT+7lKB0Vv69oybFNtboQWV
ScZazgp+67D7xWT+G7dVRjvYbxnyo68rXfG47Qz9PiGTjCMEUrrj7AJdfJ8ymWYx
VtYsOFmn8L27IoG0pd0J9S6IvMxVb0yV6AJDGXTIWn5q2RTBQmYXV24yXrXbyiua
K2fMUcYtpgqdr5LJ/8r/rqIhaLssFL3Zv3Y6iOpKRnElxYL16O8IlOCPsRrj1K6i
jGZttLCPQPvCrTMyNW/NzpmwPPL9r1KjDNdfsTs35wndajctooe8HIW6zRRLEGGT
/g9kpBCNB5Ix6ibnek5U/weFCYeMAFNVqQymK/FYorMavtrvb28Ea4ebx/ABdUgq
0D8p75jZU6Mww52jCF0b7u0Q/Sg6tfyauLKqTyOX6uiEQ3FVF+4uTmReAxSY5C7K
KxmvYND4JQrT9j2r2lyhGtJ1W/oxnJ+KwHWf4kFlLS6wEjncMjumjYo1+cuXVc27
/UAK9QGW5I2tlnHNpJFC6ySB22/jzTP+fDlN0CbGXbEmMfNMCgiZeE2jEPRbYohe
SUK2fiZNN7MdAVP2K+A4cf6QvpYZ1mHffS8PMjtHMCXAtwKgYSIee4akOhMoeKxI
OlZHlURCaFIlba+gNHKLyAgTAoRFc2qAv/BRVLIZ7BtvLTUNA9QWQqNKpa4qHpvu
hioX4rv0MgxNG9L8oJaPCzVFY1cf+o75R3LLk8tPcZxhi+pXYf048Zo2UfYSOcNR
Onqwhhg7MdrYvg1pr/QzEygMfGAPox2EZgftFQCSNnyed++q5Sn2wn+FB7CCUtZI
U3ZNmQuwQ5DWtxM+tk9mMv7xPuSlTL2Zqbt1BJtzQLu2UGL89iC3mVPxP63Edc4g
Q7Pc6VXF1KomD2+aqSM6AmIj4DqaQmCtkNM1T1eKCvuUt/pzcNZXlL8G+yRV2kMd
bxNfvcjIF0liddqRf7m0IdL6lErZAPGoTgyxn67O7NNlcmOMol5aL7DabsYIM/sp
FXjXA7l5ZLwcKQs7ItH1oB5KFaabFHnGmfMEd/TJ9aqKG8vFMoTwYphP5fMcaC0j
EJVXJDknvgKBb/SkgM0S1Xi0uHoNlng/jwyuB6+m0bllpk8pCmei0f0LexmZUE54
KEd6hD+AGQuXaXhxB2tZvLiyv/3sbcKgRQEaYZP8coTmMDHZ7hkRbSiVRCbNEmf2
5qVgD9aoJbZXD+AUBn2dKxMHJWdZoW5E/zWRjA2sYIrg2Wyvz2rk8KX5U2OY/YUr
1b40sj51gRII3o19d2+KeaoBMFpUdMNgS6D/t7aRC8WqPZqP83fBX/JTkRWAIid7
6bL1r2RzRcArme1hzhTS1hF1sHiFEG8kbzz/r9Fw6crHrW0ZGU89R4aGBVtWZttg
Pf4Co+iQaSPP9Mj7RetDTp823+bC2SpCr28+Gpq4GcybPHsRKvHTfTA7xnJvtexX
lNR9jG6vJUABRjzA+XH2KeCS9BJGbkf4YY4/ebHKcJcJRMc/IywUDkVGUO86nXMZ
4qnegP0PkFqU0gA8+TeMoZFnRzmtfrZV6av2m2tza7A1z/Z9Asxi8AV7Vw7F/qVv
O6FD2k/CE54ybxkEHdgO1qgh1SigAxMMMU65dh/toHmIzCByZax/YuFxJqEiMZ2q
UIMGiDOSKfLilZvRG4fKO0oKIXn/uDfd9MQ8YYHmGhBq9T8imwed9fNo++ahc6Op
PHpxhlFXfONcNZEPhQ69qpeFiByYjIBy2gQ4C/THByEYiYhi+aingZigp60ObT7K
x6tMsJCfJfb6mwR0bZFggSMyXuAQrpEs3jQifHbLaKqiiwg2q/qF3CMarExzMqxG
yv/ai0N1/ekJerKJOkZZHoX6sDwkXUd7x6haqQpjaPconPNzd8s2niSejAtb9Atg
riV1u/v9OX60yl6RX9VvNkF666pYS4Ue+L2U66MV1CJ1ZLUjjJ0vnHp0hWNTTwH6
F15lHfDaMGAfzbLJvy9ELVjsxtR1m6SeHDF4215D8GnooG3t+r4+zD8ljmlNeuY1
mnny3jlzlRM1qt1UOCdaxtafg5zC8I8LdF91voumQMdpzAuHewoO2/0tV+Kwh0G6
d7K3kZe4qk0eSfn/WkqP3CCIO/mH6kDB1NUVEJ9Opf0YLSQT5So+M4z3fOLa1juV
AGIM/Ajif8HguGsY8w8x9GGz3DYDdlz3qsNPM6WC4eL80joMyDiew7j2wCxsMuXi
YWBOisPCR4woXpH3YqeK7lXVAdf45LiUebS3JtszKmI/oFG+o1rMutDSt+8W0DBt
Zw6klNKfbHVcTTswcChgOlvGImdtBWMJZn0HiT4iYpC0d34xGcCuMi2UVwfcMIaZ
gdTfqxT+podNQi0UpC9XIQ1Aw+jY33npaopgHZ7Kppzau5AbxmumDf0VbA69HJA8
jEfbY4o5YG/SwzBy4KALGcVNtKMAcMno3MGNF2CZvPoHzuQfXEnG0a4sADeZMs61
0t/XcJdFZrDgf6fqfFZihNwpVpMTK1Ovrr17LylBM7WQXHo2zp3zWUfuhmToBLNR
NidrX2w3leWL+1q3WdPZ60DWdF1E6RqqKL8KYvhVD9EKqnvLkLSJ6JCqrt+l6Ens
UkriUWVpBHhwRq4BCnpOfTFlvx87miGFp0+EzDUyJA5yOzfH3wZPm6NBy8/gqblA
Ez2kOUrMsOhqSjLWtRHYK8Ef5MwqkL5s+IZAo/0u/WAku9yqUHlAqsSqXNRJvvw6
AMt1IAxi8idRjgPrZOvrNHgxukcNP/VTdR74CyXwOAch27/OgKNrUxYRCQHG5pwz
y+ZHo4K8VgptwIsOVFVTTHUnH2DFcyoK9kACC65qvXljF4LRgFj5r7p12uJ82sc7
hHqElNdIyJh2OBF5uRvfVtzMbYdZtSVFyoM3X3o8ABSwzQMZGmNhDEqNmrWKoASM
l5zwPj94nja45RJIfcUTGJ7i+BKz8HFAPADq0ioUt5jZvzJFxKp6YjyuTRdRaJ2d
+CfJAIG6UNf8Ek87l2oFUqSKUPAqDUjpQl5h+tC+HPPBV8JCyV2APU93ZEMRl23h
IAAD1QIX2RzvDrmDeplRFzrvLCOoD27Zd7HOLKZ4yVVXZIx+vKh6PHYL2P6yrXxL
G3tsGXnzc3isR/TerzkOl/Bd5M5OWFGtV+HkKycb4gZagvxQgGE9TFvZ2Uktlc/0
43Lbt43i4WBfGd9ORxu30NheUOPaN33hwY3xGCy/DXgzKnsVRuvFNmEL+/NbmMar
v8PNaMZAS07D3TILHUo/ZjzO/X8c27L/Qu8ZeknsJwiK/rzztagiY6wFh6cgw15C
Z2f9MQmNCwJ/yxcZ63b8P8bFRc8J/SeWt86LSvaWtEJhDaF6cF7ri2pnYRzu6Pig
WO9QJ8KtZ9HYRZ3OE/Zk3Wruu59UuxJNF80uLMQ89NA8uM1+1Ga4G29yf+WC7R3i
yuABRqA8a9POywceSkdSTAoB6QV5viXs2wtMEOqJwGKqRltCIY28HbQ5susoZCG7
+h+up2WoTq6Bt8/f3ifcY6Thfcr2BhDpIDRX7AEhng+4M02kPlCEc5KGWSNlkR9F
KIxEtLhRQddBD4ID+Vvr2qxKhoqqBnGP9TcWjo21Qv3YVBgvyhS0QZSov9/mEAsO
WH7Vkzej+Bi5q6kFuzs50MnKO6Y1T1Si9zXbrpz7GxzRgnq0pNmk+r5333+iBjis
k8otFjpuJZ+nSIFsRTgJqVzoJoJTjfZoAv9RhIeRth7o8ybVi5DqrALZHMWP5pdQ
bemXPwUUdJUQgcosC8mpOKXcRuN9V4qh14Lh1JCsGaxb94gbaSFHa4ARufTldoUS
jMX/8EBo3Ow7MrNAmi8itS2rfNqA0HDp8tIQtsHnwC7TalbHfC6eOGIHrTrXza3y
M4rTLaMWtOqrGv8Mx0M0Iqg6YjPG+nCEFQcvi7K0wgWvJntrJIW7SlIpjlxfpAKZ
vqFgOYKADaJSawbk2hJKx1S5Pc5cJdJ1XybpQUZdckb62SVd5ZbjCWDD5u0ljT4Z
PrARW+kIswoe32bW8N8RgBlQYNSyBDOgtq3QmRT0yCgZIROC7HhrtQbxrVG7vqia
9km3uC7QB7soJow8EhnpPMx5CzrFK8dTaT2DhtecDA9++6sIAvpA3f+oNbrz7EZH
jofU8P9M3OI/752+OGa/Tpkc86Wjs7eMeVkJ5xKZHkbnG5M4Jkim8eGbQIA7yiD8
jOqfUVXu7MYtwNCpiCqwKkbRacYHbIwD0MWQh0FOKNZKf6uzsarOsOmr+BVaFn6C
JjCZYHyQvu/WIw3W31rOOb3ElwVasg+7nBzrR0y5zpjXlhCko7QrRPekS4DRo2Lu
wJLDszufVwIAbPlVMqElWYRCseD9dnsDmCeI7BDPStZ6lmQxKNDKoOIqJRxuZJGt
dQO8874cEOAPV2yIsrhhdXmKyK0WSbYBGQDAOuN43UJ1VODFGUXV3T4OpJ1nJH+C
IHRQ6R8pCmPSyHYyHAcBLylBY50q/lipOr/yR1wGzZ7jX5e8veF/4HWJ96Tl9yUT
VUoPdx4TX3tqHvpR89CtGcrje1gMKBcxeHT9FIo7b8NY6VzjXtcJi55K8N2FvG/3
VeTDaU7GT3Rv8MC1rcT1iYbIEoB8hg8PBvEYQgCvsjhF49C+3FDYACCfabJUelLW
DySdlDfbuii82VQdYOmHsRQIW06X0OOputKan8BbJD/FR/CoYe9PUzgkO77i9xdf
DY49ex8ymJVuIrjJHvClNWG8wObI7mQWQJP1gIdMNlgQye8ElAQvKKeEBC6jbpTH
3o8PrgyJQm3LQ+JckCzxJ+E1PLPIXgK60Pvv1B7feLOcvXrgRbfux1VMZOh/y8vM
Tuki5OaONLaClwf7hr7oPfUs+pBuNmxvptsA7lOBIPbMdS/25p7yqOcvx+U1kKW0
/itbbdk0bvn2ddDe+rZf37serYWwXSZwg/PmJLVdHAV4XgaMj5qkUfcC1A5W+ZB5
RyeXeDxnB1YpZgVfB+JGRMBRaHA4ENBqCVSxgZWBK3fLV1DbC/nk742Yz7tnaOhT
iCkna9tsk73H5IgVbIBpIKP/hoDrYXtA3tf27cZod/SqoPo3dKHYBYfSNgmNxlN1
bSYW4GMjFMnG+hgDZpACtweDOUCdijHDhiIQ7bHQJ/j8G5TXqQ07PEncU4OipT0Z
AYrIlCSssJqDRsszn1l6zRG5c/2rleEDcvyh/I82X6SCHw7HnQCSJuquAxF8MSCo
2GA4/5CunMuSJ9o5hGFLhpIihXXKb9KslAbjue21e3r8r53gApbGvpgpwmOoKAAB
5tTN30K0TriV0b/vxs/e09y/aZsIgoCW2bDTf/iI2jW6fY2+1CfbnYBYlG4CjHJn
m48uM+5kJdDdC8tOxpQu53QjRg74D8DVDCrslyg1cMaKCVTLLYXR4gKMBq5xoKf4
x8Xx5YjPnbglp/Fk2FdliTwDtF0NTF/xhWlMU1P1YH0UZ3J1Q4N8XsXJpDSjH+Kr
A+R4I/Ld6AwDW+Fxn+n0at1MczJnnvrfvdmFqKRwsrTCm8QwnF3tu6AJjA6gsoj5
FQlRc7gvd3FkZMPS1U+sViqtzjV80ihEwT0yr47kk2+I1pqdR9ydkGBAz7u8QFNe
nOsjWZmC03+uFvsW11tcvd2iSpvslpRAAb/NpJDCw8FTPmcZ/XGXShHuE9pCcZdW
dHAbcW4z9PhIn9sg72wtZteK/kgMHM4rNAtldXSZTTU+rOk2bxbbSRr1x05poobd
ji7AUn5Wbg1mY7JIbpg3dncOf3xM+m/ctselddps8aTfFQcAw2dmXzmG4tS7Rhot
PWAg/Tz+ZcE8qf2lBBRwPStijbvwvsJ3q497TWcdJXz7VBRGFjCtTp/ihgxtp27/
DZyzH1TTiTXGp3qKS7iYDxI4PAa/1k9It4N7no7/H3mJueBuB3qT7Cc8KCpk792d
/JcV/evtSjoXUQwRjGFHzJ/9HmfsOaHOnlXT4Y8YzPPvGe8MRk1mFhvIBQimnih/
66AT0HAO/n0EbAgx9PkvDg9yb3DJeDqRjnaRJAGuEZQsrch0hSB5ZhUaoTwK64Mq
8w56pfbM6BpeXYEQXYt0VkgCR8wW9F9/D9j5mGtkcUcLx9aWf5J/6+dAPLn+a0GD
2c+pN+jMFSGh5FIlfedBcorL/dOJfuEKlOTLFWmp2ZL1i7lWGa21EwsGWO4OFuws
G9Ys7/MZjZmtIzKyPgg8gftA9yc+mA+/yQJiLUG+0qEnpbDEVTBlMwZXUUAWhMLc
ULo4UVt7g6HNT47UlserMgYiAwu2Mnf8CqEUXGMQJgyzVKL3jpMnfhmrN4kYhqzS
kog64GaB78Hv7ZHT1iV2DO0F1LSALN0a5dUQZkpSUTmIvVV+bRKZrNFmMPrbbAbh
3r/HzZzATblbknKYF6kdaLF3cQcukHBhdpuvC0vwjxY5sf0lhxU6s3xF18Uex+py
oTJHoFb4XW4FyARh0XetECwfNcGqFBbhEV5L854Z9qoNUMiIPUlEnEOmIQ7eBUtt
cH7cdng0f0pSYVRZX6SnMvkvOKDH+ND1mCmAanYoQMsJgC4dVngE8C1TwZAdJfDh
c4NMi0Gf1i9UlRIygh4yG6MDvcq6MOjKSBHptk+6WUVc8orZEMVHcfEqXaAtB1zt
CM49R2MBgLg5gi9HgjrhOjJ/nwiBM71jmyfQC1Et1VCE+CKs46lUJMfmbzTjc5NH
9cenG8yfYeG85EFYUH3eSPap0kEg7P9hEkPJc0umuKMKMorairFmt1F84W1MMZOD
n1eZGd4a4Ub26Faqq7G/llQ8HggwaDIA5vJ5rHTMqiOyVNape68vYe5LodFz4kiX
vovRiEzQ2GXQOLvIxZ6DIVyK/rD2s/Q4b2/4V8vNdMIhiPdx48AbWFtRwFUzeFOZ
p7eNhdCE+oNQfsoYDWAl5ly9kS3TZOTdfFJlxpDtlipl69rs8Fqv+vVJeuhUqNvN
ftVcni4Xaa0pXfJVDnZiMmR3OMaPL8NDMAS3VpkETlMB/26nzTym/oZZQqjOR3PA
Qfhxj3L+J3w0uo/Xb0WxwfYkwQ/rx6Ga1vDQ1KMOOdgbqFZ4mwZELl5cmW3C88pf
z173vuBwfREBOpZCGIA1VVse3QLRkV6lxD0KKAxNUTrRJ/To0Q/hiaVfX+qH7pD2
BEbmPCzGlaLsMFKSYiTYpSnTPR+/36UqgYYXJDKeIwj+gDqarK4BRzBHweoDqW02
6L6duxIuUNrLaKAbUBOqNd5K0R16yvltGKpGbkn6D5+0TIQ5CN5gwBxMOb654yY8
BPGuJRUt5EvjzSxKMCD4vjwyRj5DXHWKLkY6opltlpcpQqdGFcF10pMS42dPdBtP
KecRNxhEADmUvgrbPRhV775MVu3S0xSka5vBw34Srd/qfIkWL4LYQ1dP1JGKfyjR
RjYLtn7+0qOt8ywmB39y2NIDeAd0z+5wM0xi+yx7WsJlFlSKSeutS2Ewrvd+4/ek
cQYmM0ZpJVuNfF0xYbrdk4WDmmud5+vXj9m/iHC6yKHGGl/LPw+H9LyDt8rbTNHP
pYoeRgkMG7NI9MvRtKBoPLFMjw30vYeNsRfFlZuwSANX2d5GN+U8VfCUxCNyqjiq
U2N+1qOYB176GrSHQNZvzEco9LCJ+cIuNRE8W2oLT5Rr0b/RQYjE6POFMlbhpmu9
kap3rq2C491PZKxUhwD9QmGngfuyNj6TQMN8cQLz3PXldkmYdRy6cUHXwYt6qXDC
DgomUZj8WUc8e3oxJ6WQZkP6jedgZN1GhGX3r71keVRdqkY5zEOGRAZG2mjGLUWY
lKC1Ue91zPtYTf79flVRkMe8qCiocZpvwKuW8lZMf2Gme+gzI+CANRjO1kH1UX+A
CG0WgEPDu/7JQIm7RtqCg1CV327Z1deCstZPeiYbsbC2WwJozmPq14wHhGaY6Obm
4oR0Po4rN6qzpEgp2IUyDxjV+PiRfGeDIZWdi36DfroVRu2BvVDYfHCNYms3Nh4I
7RezN6F1cL4X0L1k+/iogCTUACWZJXejTQayQJfzd79JRp+K8UCYN/Lt0Lr2mPLb
qmaNSvidkAXB+tRhHe3jRT0EmGaMJR5N4T/52UmEvTo+P4V0eoFNQiyvf8KuzFcz
jcKMn1cylfoReCMnmgbPdpsfSerkb54tA4s3LWX2y5lRQip3Kl6YCyUbm5raIcok
Bknj07xHnjk39x9jLxuJmW0nNDqI+zQVxKMzW6i9ifvEVb4bgKJnSL4th3W3kyx3
VFhnv1ysQOHi8tNxXUYqA8nm9ZeT4KPJ+zLbYoCEO1OmGv3qag9nLfxSvOGv7AXu
CRjRQdXqaRzHT39XatELsu/b3dKsLBEJ+V7+6jzQn3vb1FEvC2XPEbyYFlVvx14M
DAfZceQp/DX3oO/f6eCnnudx1/bBjLSwRSV+lXmP94ZJVZO7A+pkr44tUIYcYWDJ
F24Tcq7lmGuUwfFsjysGcJyJ8sr9PSqGGsvehb2ooQQS76S0ObK1ItcAQqLk6o9y
PurBTBOE/97yu+Y/f3Jfjl0QHPQBV3iJlta7QxwvcvsUCN7d4DfjE4oNXVTspONl
i3544td38p13Aaak+OAbELNMHfluqTtpR/0fhSnC/unYIUA6Atdo3k/qPA562yuE
/yVwM6XLWnEnq3E0n3RfpkGyaXcvP8PO3R8lokN89TJrj/CsAGPLMj/+SY9naVHZ
OvypSdEqFH5oMqnSvWl5EkXkyjVTnJs7Q7YuqsqrzdAg1K5gAPWslWDHnZlx+er2
LrpQcgEODY02EsyZHu6Zqd56SQ9P2N2VabhQTNjjaIGJqbEgvq8eeq/ozAhedJ5J
zOkz1iKpxKGXDdhrYltQJyUBoLncdLLJPG5LNwNE1hNWnvHVtdh2jO35f2qIZa/f
CN3I3SP0wUOTTkw97qArDMdcJBdsx3w+A+5l+lOexp24W/0qmhYh0tVUg1/WmzHD
xgFNeVbyLrXWIYQUHxWRHcxe78MIoCYbVEd1SWJNxA3zTiW06CcxCt5dpMIkmgQu
Ryv2G40DQSE9bAz0WOHsSoih+8xXJyyT7ylXxBLH8S9hqD+j4YkxNfzaVWo6BpV7
LaxsyTlz0kaJXELm6HX+YbgJnHBeJSrLUPlwdolaFsRoHxMFswfJtwN0VXlGv+W9
Vb/Iv0NcV7UaVHYD0Pw/jzlt2kZPr1K9LZZgPPjcPxkCL04r22m+uqmV18escS0+
RNG8gxufWy5HgC+PimXWSNI5BD+ZVy5g8r8foPOuYtP0kBOSAsP2/4bZU8w50riW
ZYXEJGdD9ZyRqqu8GnJVZSYmxseZ/5r+gvRgnzih4oU8QpwN5RCcqV3LGW8k9T9a
r8W+EqLiey5uGuAzzMWUY3jpqsBYhDIfCzGB2v8Z7fug0EegFS/tvIVMB32vWRjR
W5vHNId+qlYdRB8V6A24hLRA9T8wu4Jn+ytjkD55/HKDLu4uhuMtauvbiXg3Js0i
6F3uW7rzrz2NlUvuhwzeekDCZhhkYFzMglOR8FDNzZg5uHLc90P1YMY722LKWJDd
1UEhaptgQmYbm38mxwHRmBukRHWakR3KJg/NU4NTxIwYqmVy4si53kGUb3OxOIzO
faudAvI4bTE/fneR9xPNnA7fk78vRz3pT9NwiAX6MDJjlJIZmuEmd2XBAtuNwZNN
Kw7g6YjSOkItU7uxENP57b1nh0x+4+r5RG71TGM8dLsJTHRcZQskavdaoNf7HgFi
iZ265L6pJl6kNwx/FR8WE7C5Itj+H3gdMnyxjRGPhOne8FX/mX98TZNmihQoqLQr
Ky6jpGVuB0T0I1M98iC3QNm9wBr/Nt3fYxT9R6bWD0AIDM0oh6A9+BoQGazAOzbb
Z+hBGwk5Ow+M9RHhzMPrS6+/YCaRES7iSbT0gKeNd+NL5WixyMFyWPOIjG9fT1L5
1VaJWkbOLDw+hTZrQhogYERVLbTtnVYNqJHBGwmXbbxINNhecRtQyznlp/cNKJ54
dl0cYDpTWU0hp9JH7xBY0NgB3ul6TvB4KISLEPeJrTLsMmVYdm2D8xjZbgZhSzuk
by0FmhyryG1O0hXTBPexfzD+Sbg74hcwd28omEDv7A+f7DuISHerfEA+bJgXsvVF
W2ZnuNAzzo/H5qN2kIWljHYhxkOXjoeINiTViKf9ke5IquT58a5JwWgIrEeCc5H5
2XqF0Xp31mbXu4IpAGCdD3EVlGeduGNhCUFADPAWzTMF8rGMYWq94ienuSbjSmtP
YgMLF2BnDPN9wHrXYpGFgBBJSVDdUQWX0AFtoPjAs/tl5zME/0z42/tYRGOzbS9Z
2dYrpP80EtGejPvcZHvX6EmKND2EHtormJ0u4oDmA9rY/NKYAqIapbtMXTM1Gjk4
/L+q5zVT20yuL7wrss0S/+k22GBk+vqabOpGIuLBdpkQ1WLAKQpen83yjjsAvwEW
+oDDqKG6kJAOKF5FO17Fyif2hVhtaxQnLp1LPc7wxZDEBHGQ0WQvNagQ1VwLcr9r
1Wt8C0w2d+RyroOgKypW02EFD96GdfM06gHifBGSFkIgyPW7NiS0nCTaJ719ZOYg
fQ72mrXBaQP2uDgj/OhF2fEmvocj/6iHZBRvLhz1Nuv3I7OUUXQ34k/i9QAe7wdh
oA618FKe2CHXtSt30Z+WlA7uq/0UJVOzjP7mk5js9dn93V1PgWdKb7h1vk7/9Lvp
LdCJJvzetkiYSMmIzF3RZ9HMnUGj/rysqukHafTmVW8AAO8vnSRXMlSm7nC58/vg
MGOdj05zQeltBTovjzeD60HIbs1az//+tw9Iof5jLLLpCo6xnPx2x7DlxiZRMzDT
X4OKHY2T+wrdovm2SlvlUjhZwh5cu0UdxREYkXrSaEEpH4Ke5ZCxv/BSObDZmQkb
PkNfi/kajkhRqT56YXyWtEGLgNe4Er4clMaKW4bVVrEgBTWXEFspa6zdw3hVqAsA
IP2W7SRb5GXNAYaaAqLk655XmXFOSPe8AQxSITS0HgrJyIaCz0unFfsbFuHx8uUv
jpai/iQGKJFhQ8O+FocojIXc8jKgl6tDVJjtOJe8663oAxzjRj5GBm5xpGffpmhG
WOWQHQ3sQtfxYbd/FPFJdnTvSxmOXyV1Rs5I4kHOSpM4plDcYXWTgGcz4As+mcjO
iXPeTiW2jjLMtuErgpIXaoVywmAdnFbj93SoFEFCV9IdrfS7kViFhZiuJOb12zL5
M4IqZE8dM7NIAZZggtpWqsRvZBEWh5eSwK93uMQ2/cmSv4oGOp/VQnU+f6I+Kwqb
KCCwCS4LHZ64sbS0EM8PVmiPp8ncxFrjTKQDbtCNCbbj5oy7QF1znANIjN2HXAvt
E/J62rNMSRQ77PvSJNh9IPKGrk2nKTxHPbzDZbl/Jl3cmifwGXZvr5LwsjVBfNDc
tmkmfqTXiWXRhQp0JKbUVBe1FxUBRnaUvPon/Yb+cUW2E591g0lG01nly4hKOASO
kFAxpLnyDQGUXXlKVpwTbmtTJ6otdxbt09Y6zLMgSXPbGIh3dwEAFMdA+qVsfkls
tVISsp3JJMJABnGqb5lfIm00S7PnkMF5ivNFcXTwXUKTZu1UDrnBjBn2su1Duzpz
th0/X3dZ1MMcl1/ZkgPuWzFCLmPaclyVyomJ1aY41ttJ9s2Q7qtUV+ACrOQ0WK23
3yvmSMQTyJs+nUrHckFGDROfqyd9XPUr8t6Mqw+F245lZkH8Sg0DYLzFPfkICVO5
L7gVXhRCOfYXGHBt10R4qtYlqBcqJL1EKWsZygbWdwHWXddjIEJe0q0tCvojUfR8
Qx6kYcSzKS/sjLKBDb6gUwFaq8Wj5thBbwmswZ5wFBSe5pdSsPwLWse/b19pIQzF
r5nHymwbaG2/iIuTsfS5eoMyonsjdpNNZHg+X3ZyDIR7ZUHGOyFMOPLCdcRQ5CKs
td+cjaooC3P4j4OZdjgGYWsBOuRfxUa2KZwS8TKwF1RM2FxNkMhue7jrIxsmFFqJ
MYhTYlTkrn8AnUNT0bXkQ5ms/0RHYGi976h3c/bfhmcAoOf3IZrf57gT3/znLpT3
2defb3p9EcQB970uyV2xi02hsxxCzzxyKuDy9ilk8nrXILKrOug189hQ4oHnaVxJ
h1Or11kZpaNoFZOilSrx5rK5hSpHskOgogabXmN6aDocIAXGN5VnGC9ptrBAUp0X
eT61wvA2R6s1EFg3MRJYDeX5XDVKlIvEUncszk8GimJ/4MVDtRxRR158hUQsDwmy
EnqWOZJsRXSqwi/MqYFJyn9fiXY0p4DrH0mcbiLcSKt6sQ2kxsySAx3HYc6AFZxO
xEvMGzkBlzrVY5yWzTH1V4bwGZbGMWHuNMpUnNTUZfHlYF2TPPwLg4WUhM7FoNup
kKJ2/WNtUB8d1difidxpLUfi/LSfgRB0pZukxTbHfCVeWf3g6uNBCNebPyUcmrA+
Wvus+E3mlK8evzntfS6N5dWHTl2VOUP7BgdaG/UwxBN8wCP/MjqntH9rb01pXqMN
G3ArLfUuIA/bPXYbJLl1NVTs+j3nBlVARmbN4cRKp6HcOLgH6OxFrw5GAb3MlVjs
E00nKkWHX5A7kkJ4SzIHfrrwGMuAl0tno++IWnBcMCClUZ2aIfhEjIdNwbtm+zKu
jLcL10Z2Okvh5QtVSISWlUMi7IKNicxr+XFyDj1fsLlSCNR05bjZWR5dItYrFkOA
99kzV+w1OtMSbBkOYrfatklQjHI61oTTrHksXmPdOsug5c9TfDKQx0CQ2guEuLGO
rtPCmHCb9ZZC9Uz6rYhTzjf4FjlSDFLKw3uTi0T6Af9uEPP/8y+dAGHIGtNdNRph
SOEnFX710woCl6RpEgJmAp4H5Ti4CFp6VXd3AT4LYqe8ftSkjQY7uDj0jOpV1Iq0
u6tJJ3NJ7lVtbeIvwCAee+u1xnHrI25tvrog10TURjyC9lrXVn5Q0BZSO7XSJzpZ
DNkYa3xkheHHJewK+c5+2nTimKNfOe6khGlwHSEh51HnaFUVKK2RxgUaYo/kmbg3
ykiQRN0umkjcdaSa3/p88lsCOTR4T6KiOZQXaHXKK3DGaLdzIM4CTlRjFuJVbKLP
AOWaZ5xh/YpAw4rjkzn1Y54NeJ4g0tjYBxPZp358/CZPokku2vk4gRhYWlZ+odJD
meHSdfMQEDyQUI0Auu+FDPz3LbcX3EqtdJ6s076jXHrNzKQ8uTIbSXyn8No44dcY
lAUKSIAuFKz6NbtmuBlE2E59iY8zcSZTl8sM/5ENYqEf+wXWoGKz+v+MI4l5Twfx
63fKNSzVIIN2fH4I+9nMIBX8NjRkQOPcRPSWrQh7M1l5dA7PndIiys3DE0hH+/D6
llUI3Zd7HV7LuyW5VPkT3ZLHdyydHgAcs9peeGU/ciyPsklCCihxBeNiAn0i4dTI
0XFlhduCQnc9srkZnaUh0QMYma56tts61xgfJSAwmobTG+iN0Y86KuDln9H2F7o+
Str7iIAsfB2BGBdVWMnl4AXyyEDNnuA0bktQu4FKjxRhHV5n+6vcOsHQ8OtQ9XqL
dcXobgpb0x9+3epObpXJWZoq9ZKVDQ3NgqdT5ps7bhLSyZ/x1BeFHtIH58CBKHML
cT0puLS0ojRqCGeRFuVN49ku01NzZb72X2t+VU3Ex+Z+eA7iGMxqli56ycIitwGn
ttV75Rz2/Km+Oyg1Rcj4yAkwwTWW4jmh0A8rFVSJACAp6NVBjFVaZ/A9anh2iCBk
AJwa5mwPgVBfxY8Z8j7aGTPwo4wrIBC01tcWF8SX7TNajjSMHeXiv901OxpDkrVk
mirI+OPaEDzrGpMYcEQHS6dV1QmWzyunlrnYYggu8e7TpG0ONe+//s2WTzTG3znk
I7o6PqHWX3IzcMWOO6mLd7CkCeHnmfcmcJDFMvLXOFWAE/9BFxMfcVYrOApSRgPP
kWp/L612O0kzHvsUhDRxqcTfMyMg//wFFYswsYlmrDTPYLkdBdZjtFSg+9I2jRLu
cIvn3/hDNOdtC5co+nhoGX7HzvlGnocS5rA7Cs8CwJTstSDOTscogC7uJYfogw6s
LI+eI7RnkHO0diJBp6zSB/WWyvrmgyrDkrLZfTuUip6FGQDIQ4q578WiSJIfcF2h
rAOqUGvqlATDW+f8r/v0R21ukmDLYolEvp7vytnqjixaXGJkkFwKpKsuVvOaWA9/
+DB/nJ3UlYWWiQKlidRa5s7qrxBL8bq/bgDRWlYC3nHdkCXhy3VbG/Gd1WlmPO2Y
0zIqOcbh2+m5imgWx+vfEUiOKS+bClxf2Oxm45lUAUfU7ygsvGQ135mnIAqrMin8
1oAAwyc7UdCRC9BP4wpYd0lIrHAAi73jDW3zQNDdbY1tovvnP4XKNYPrafMyb7il
VmrSlqU71KR+TBgC8kb9iLKlWbRZr/5sjOuXNwqIUSRzxGBblZwsckoKFJcmxyZA
ZxPSNGZjbKIf/fK5ep/TJgtAop4gyKhLkF8XFmgv0vdqEPHS4gfmBDO79NIzpGeK
dvSAT0QaEINvRMqb8eW85RhLdbNokOhqe13MhbPNQHDWnbv7D4ORGCWVRzl94mad
6cNwrSIZ8vOOfqGoCeWHkNcn3dJ4AvCC3g+bgPN4EErFchcontBb6PQZxK5GZMZX
UJ3XfHIyCUMvZrEFiNuB9kuk/w3pNK8avNzZjLfL8kxeV/O9cGZgAcaZVEbXmmh7
3X1PfjpXwjus337WIMkh4H9eQoPldGDr0b5XjAWYV/vTsRYr3aaMNyeD6MCeYbVO
keKpxGTEHqvLCC2YhbJeb1lTsk7Xhz6s/iVMSG/2ttBrkxqK7tFTLtysLW4vJ7i7
lm4xhx+oAodvomM9FknDGvl1Coh5rKDnX7VEnwakKTPnVA1QWH/grSn4IhrtHfOw
nJNnI8NO8Cs7Y4A9rvw0gfnKk62Ycl3ILa3uN76LdYKGe1645zRnH9ocMTKEBUEA
eMgF5N+0UW+ujd5ZanURYCwnA2SVGhFr027DuIR86TQWzc0j0Q86gBVg8ko9ZbDc
k0NBvI70KSVmwIjSadEf8OujQcy8BO/FpF825x5JWywnoiOF5lePPGfyp5PCVaqm
oWKeS7e966hWXmlI7AZjyXpTAgu86z77BeLPtCpKpq8KgSk/wVvLwGSQByTj4yNo
IxzCMaCq3t3Zr+yCNOuLKYpdQI9JCl1fux49bbrhCeM+bk+n6kB/Sj13zdBSIaI7
fxnJe+n/3vFyQH9P+o/cxh7LTT5XKhJkTo7RRI3euySb/GvyKP8FMpw6X3oZk6GI
ZlbxJ8BdLcyALC2sQo4eyX2Vreu2dZ7r46zNLVdpj0ilEvdiHOd2GI5p1cFjMh46
INJd0yZj8CAJjfhTiX7+Q9ldNekGe70jL8awWF3+52Q6ng23wsyE1yXqM9YLLQ7e
WYo1/gFGIacDRxE3Lv8jmshH2TabWCvn5thizIhtk4HwqOvdfViuzQxt6qhYp43s
fewU13jqxQjKJwQckF0UY90myMPqILPredUBp0u+7zR226h1VBuKQw0scxuNXyD5
sB/8CSxtEpeqBU3Zre//ysJ0lLoquV2i7C1bIWro9bFW0nYr4quvdpoiPjcz+2Eq
k0zrb2OI9rqJ/MX8TgB/TDQJIVbyfthnFPgD3kI0pJOZgM2ueC1KCU6CXjcNFiFp
WjCE7pnySqQHj3KPGplV8Jc4hjbG2T9akx+W0Hg2bqwQv0faJ7FTxotKbfKkNX9Z
/rduhMVRopHB3PQ56D7F19fLP+tImlv4jcSzpvLUdT91sm38SYuuT5vQwbGBqxo1
IRCooQjDz0XLYSU3sT2Q9f3Ep5nfWLN8VfRgEcmz+0bWF2GxhTfhmc3lOOAnJwhU
y2U9zV8wxwlaSwBYHNhe9FKn1JB73wX/2M+E1vvPCEPRz2GJ8Df5LjAv3OAzW3PY
OfzwBxqMN80ng8VcUzPYCi2loFq5oWP7pfgnTHI5WLteS3gsYGCa2wL4/dhJYRwv
FjRg8wXLrBmp3099Ech6G6mdXssIG1VKDSM7HXm4oQZlR+0O8XLlOq5tVxd2OIt2
6bPH8LRv/uWMZ3C3ZlGFDFPtPnps0TKmcwnbKwln3m4XRAUE/qkQOgGfmNHs1hsx
uGra6qN+oWSj0FDWUU4IgK6Rom8HNXhh9x8ByZG7TTbcCF5SG7gf9/R16Oavr+qQ
F8LokbOik0zuGZEN+VvJZLZYTDy836uiJQmPIzD4r74OljAyuh3jny1WmMwhrKaK
qgq2clUu5x1dKYZrHcg5nWVhiv4XDc3tgiGWh2sh7jgEe632+kDCUo/aLecv/f5D
b1c1UzK+/E07Bcwit886y9zWjvb9wZnRleruWyjTCSDmDfw7WoxGDHEePPSBs2hP
0+cFGvdgR7xWzdboMXVh1fSKo832WkpYLPUgwOB0ufm1OxAoj0MMRNxJoqhHyWi0
Hq9IVfGZHnCUjigth6zQjsKUkT8x5wRh3Kw7qPQak3S2iDGO94tL1FfnZYpwvhis
q01iQawh0Yp+y+8rrosA2LKEK4ClUQ8FNgUf2n2TaTPP23o7M7ZDNLAFFUzNRtft
ULNyYjISOxY0L4CBzTJ7mcHbcbWf9BThJG0qJTYRBLxh/c7EFBXptFb1Avcv97R0
XjbrQc6SPG4f/Dh658nreGJCIgsH6vq6aHtV+kOeZ46PedOmRjgMPp6rvZLsc1ss
2TYZD0gNvAUPJkFNuYL+0rMD2KytnnkCoAxCKMAtl0xE+lnkLc2lrqspcZGBvO6v
9r4nUeIpr5rlHOriiliN0uA4c14SznuwDeg4A67xLvbXgrVxBDUYWzcfrX2FT6E6
G25F5hczhn+xLhwWZWEXPKyDsksrlb/4xi2mOmaGem1z7oNLWfOgUqdWfabPo741
hLxJEVFcSvIm9sTQMtcl+g0ZEibBnw31o+WwkdgEgdg1uidw99hr+LbDsC+LWjmO
U92FiuOKU/s/9u3y6sjx3ij+1uS+A3Cp6p/JU6oFgYFN57kiZ6Kqb85ZDbAicI3u
FtV4jQDgfiIPRf18twB4pZCEwxTwJ2aQY3rgWbU7yg4HRJ64Rk0KA6xufBkAlPUB
Ao4aohTPY9V2aMmtvGnjtt4cPffrdLGQQpifmRNmEN83EoKrqPuTzckph+Ek9C+j
ZJgY0CiteFwTF1+7MNbV7abIelSBzohX73p923auKXdZlF0oRoeeObAUh4ZPVP90
OGdl2vWS8ZYcXbdFc+7RsHqIqlxWZUUrYX7LrBr2q5Iavrg1oW27fTOB19lFJ2NM
6RAhqrFZFUL+6wGZoVypLweDMcY4zTw8Bpf/qhM+PiEqduJ+m5Ivq0MbgLX2ZzXI
F3ol/zw3aiQuxtCQZ39omWtgfRQnt6ARbcCQco+KgmCazb9IJLRVRROTVX3Bl7ac
031zqkB+EewrEw9GnhzAdvfMHHI6bOA5b92aJ+cNgswvcWHsj/clRMfIHqFfKKBu
A9y2J9xm2ndKAd7BM8/ZPnlXNd8WBk3Nir1+arO4x8hk6TCqXV+56JUHT2V45gxh
+vOgMaodwVUpd0Uq8yEyQQGF02/j58hTC8kDNP5JQI+WAiXCqeGU2yWw5W5tMGgt
OzaFcRLgBeDAyjdNMnj1XlUD13sIjfpAU/gKKI3hvHZXMIl9btsSe4iFmyoY/f6q
j5VqOZwwAQDiNKDvgqPxRAspmVJFPcQEMs/U6FEffLrj5dOP1ZV2ZfXduR1+XZTv
2rvpDbX9zdrCOFUA3IpNZKDoWQvm4EEvQ+BWaSe3UumSB4NzwgWvttsEU1uHidVQ
uewSF91vUQYLLK+Hy8mpnCGnCaVLqbBlyU7MjH+QXwh2MSdg/ZN5wms6obo96L8B
kpdNkteZnxVMZsDHw88GNGLV8dwywBoQ7wlSaO1Bk5WVdSos2DZw6qECHtOuxuQu
9zvfcnJMCB30xtKktIDuvlLrP3An0BuUl7ul/YjprLARLJ4rI2gob/GMeWO+XheZ
efDa7D9g+mcGwrpw1G+VR6DynPZDuI704d+k1MjZY9qwVxrIg6dXZS+r8VSdM1b6
oQf3/YrtKMwsyhgYdlptdUUmJeY0k93vKfWfsCSNMWLVQoaCIlKcw41lryEEnL5Y
ExePM0AcwGvFdC/uKlJM16AnhGAMpn7W7TMXtXSyyjarfOBH6kZugMUfIz/ERt3v
2hbaphEq28lqlr1oQiiTUVljm0qUta935+c5YrtVxQU/plVYJ1mw9iAcfQuAhEWN
Ek+4+Jro3bTbkaUYtcrkCQgWPkz/avDppf03HmTdFq+QYYN9A2LquIp07evNFSN4
6REWTAC7D/RD2TrUPnbcOAWJEaB+ygHBlfLLx/gNtdZlTYc95o4Mm9iq+3oYQNiq
jTKSyCidwg/9M4JU7KWjWBG5ul2x3Pkr/9ntP2AawSiPQJMyX7aAuatD4Q+m2SxO
C0z/nJxvMUl06U2lVg3xwLUMW5cFODSXLR3YO5OfjbthW7yShVfjKUgaF79ZtJCj
EduIk1zuTyfmgVLbKt3q2yYskTk363L1zZYJAiqEwDJW46b+rj95hA/xrInTSna9
6ibpNz6DtQEwH0Yraz3ujDdgjmS0iDREkAVjqM4UGJnlMuP+sdG+RIgEWrF3LvQw
n9OnNC5/sLJ9ojc+cJ4Iey/x0IvALPSuc3iJdSjnwVOZd6Nb2WKC2DlVaj1649Ai
dWXHrl3nFB5k81uUOngpEwlKRZIFFL4n8EnA8zsi3TtjsK0K2xaEe/rH0oCxFeDW
rqNvUBsGUgFZl9GSl4L6fMwyiDPR1w+oyw37fYimlUC5SexcPQG8fTGm6JENbT48
XlvH/gxF2dEbh+A+EgKPjwBG7GXs/X8cjjhICdDZHd79AKvPFNE6sb4PoGdtL64Q
XRxACCgZSJsxfuEmoW7T7FwsMsO0WORU0BMKrRGlWX7yBI9JRxwONPKseO9ioaz1
AdgUt2X77o9VbFC9YNX4wCbRfsjMxiWpE9qMNkHJ1OWZfdu1l1NQUHqxXjW9AOlA
+JK1i5el9rPPnm9szGBAJxXobZuWLYFpqlF0qdl6UdRNPLzt8ncJ8ZH7rTPFqKkC
Oo85dNz7uIX3tKvBVTk5AG6Jb+Zkqs8YZozfNsS6ADTD6P8E96wafd+sh95sN2Wq
wCSiaESIuaWf6MIS5Vbsp1S2njc8tSHNoCnYR9uSAalkLWmmI0/oGbdpl/Ofl/T/
3NOzKfuObpN8jL0eZKMEYaa92Jj76EBUtLTOvmvzhOr/3IPjNz3DzzJeRQhWADHz
mYxzmhpkkI122tFotcyvB+O/gBwnAVDyAAM3XMx6TXpIdtShZpd1WLPC5PhuPgju
vNjC7qOfJOEUE1fvChPhglUeqO75J5RUCgDkkQTs4mdm9U5MXs2XQcb3t6WcUvVb
OnUYpB7sUBN2PspWbcqx3R1QIKfBzZ02qKHcDs/y+SDPzDKUwxpmWjPrnvLbSaJ+
oMrS+kp9YguYuAQkqSnr9nDR+houhfy6jZ7ke5J4r3Y+cEbVfy9SdXnzN9JJmHb0
fwJ7fq13fv+gyna09109VtXkLfbST7snld6VO+Ik0k2y11laPACsUZlvAFrWD0bJ
WnZ/SJ/eOUI52YuxM7AK8TFibBVqQ/l9wcYI+VgByE4Nh+UIYiRXL6wlpLTxMsfH
0lC2oreZppnfyTuO46AAz5y9DOkAlh/9eyL2VrQEZ+YOG0TJ92JvmEhxIqgzp5X4
Yhasd6RyjDpc42uWZhgiEotXyVek80pPVdn6tJY4U1rdBFsjnGc03hA+a3C1+ase
qz4tzF/9QRvxnPcb1/3UwAS8XKSWy9CkxSc1fcZ9fwb/WkOZ1bfDI4RdCdL7X2Gl
GaavmVw8vAArmmwbH/guxiCC3l6ZAKV0mkxMFMNWBllU5U1H5sdeDPl1BfawEuxG
NyF9cdEI44QHUknIydLpmTvfPpkiNjLzTAfa0R3h5QnGcgXODfG47Ug0PVyMl+9v
wRrloomWlqOgIxBQQ0MUh+BDWPBZI7WkZi0lDuSVsDqO/7NF6c0JRLehPzn3eABt
a7Q30k22Q71U1z/F9M1+kQPn20pQZBGiu11tRq9uesh+tZQZaixR3PNwbn9lIUhx
ZwdGmogKOyQOkPsfrJQcChNiQKv66/CgX9GkRlxR2YCdP2SWE0XEqOgveecooNBg
HXi0jzuY+yE19+QcD8O7bDBO5dkspAScPu5pMtfPTnTgOsRIRmxfFvtTt5HVa89O
P7xEYFwEgt2/sYiy9rgegOIj6phVc8laK+3RM1IX9aMrVqg7WfA5ZpFvU7HEcrSo
s5Yf9mWVUA6SdggOghEv1S69INwT8Pa4Ht+oeJk733jMvSS12SjPOOJNXXSOgWnK
VaWzPWQo3qzkyO6fB7I2qipiivkr8n06p9CbP7MMRMM1455bE80QV8HxU0rJUuxn
Ip8v9XzIW4LA8Y5M4KiDt3EvJRSuTopoJ46CzD5k4rHw9juIYly2ugh58dXjJVEh
3NXLAJUaTH3V5x2oltUInPAzUf+C9rmZ2vyb4H9dgLXcjamPl7ug2HV65MR+PPVA
MzIVIEBtJUSy0UGkxJq9oZ3BVl6/Hux9nNQCbX4GZCBPZXnlFu/7/5+25UCdLOqs
uF1/ni360LzRSUC+2JJsJLdH/chh5toijA/ir+PisWWXmlPbKAftYPp3Xd8iEWL0
wDo4iQzzOa0VZD0riKzXRkf68f0O0lei/vHMU12EAndto6HtWZ33DXqGvCMhsVzJ
WY+W538c5sdLzZ20V4CzV0puZNQGlsQOnyPrF9pfXGczW2PuctlzZvrdryHdR/BG
aww3oNL5dDOFhItD/kNqgTnb92lhE/YhBi+d2JSCpkazsC6z3VWeOfE2vD1EuMD/
B6Tl0K6vgGmGXKvvlDJal/nQ77bx9vtTeym+jsKlr9lT+NFuSGAt5NUSnotI3jp+
SDIfrijxT4rBnd0BOxm6nl/UDAwHZoubsbsG2F2GE2CgqJsDVv0mzuAwZPU9mhqU
vlYgzwT3pEBdIK5NsOWEnGUaKWQW7WB86Uj76Gzed3QZWytsOD6elr0gxY4M8aFb
MDX4OSaVWC0E+Ba3C3x7qThD/I4D9YS6RWHPR4UCBl8eGkhvaeOORnkAxOj/xomT
ii60gLXbCl/EKxFI/9K5OEWO9GxmRQq9gc86YcFNuNJ206aN38UzjGarEY1Lu/X2
D7iLyhiR1RzABhB2n8Sdr4kG4y9zDtD6R51eG77+4khLyKRoh++L/gMuO4oD/Df5
uPeV4wpl585zwTlY45XLGkCh8UGhkN+aLW4bc5hYY0VT8BrvUhhW93laCfzI6qI7
+WZQAnXGedng3V07ly+XjVWGKUZ+boEaYkvls9Hh14Q6bsqs5lFRBc4w4ayrMCP4
VcOzhBpkWyIUowp1jul8OrNGZisYJM0OyMMlUznOB2CWE/jpuw9uJNzjaYIOMswX
b9xbWmtQ51+DknV9wRzWd+Xb52W5HbbUnQ3Z37cb3qdMyrPcg5IATkTbFS5J5cFK
YGFYwLVoRTHlgGZ+rRAoHMp88k6QsVgAgh2TpfLhZLqe0Oq+z3uGeEb0hp7kJKWW
udjrEQYib7ZoJgcT24d5/h4CC9RcSpifJy7yt8wwb12k6TCf8SZ247TLLblyPSte
ECMkojL7z/pOw7UX15WwsIwZhpJV2ZRaJRttMgrk33sNt4lyrN8m+DwRf4E0z/Ho
wLkTmLx9qxInJ/7Wo++BMkApZFGdiKc940b4TTWKjgDm2PnQ39gorSxY5fzTYEGO
IfodtI1WR/Iy6UMYt0r/LIzy7e4Y2kI1kD6iRolnp7jklnuCs4KoCsQLDQ7Fy4XJ
W4wiVslA0rv/NR3rxTqMjat33ZViuqYMBnFgwSOFQtSuKpnpashOjYV5uGl+53RP
jxIFH2ivycO4AJCqkhz1pNPmGrWSPZFK1ffq3R4lyA36qEWhkADGHwLrUzdmhUO6
o5TEBTslPgBamfCErXAwkt/4oyiAXte7G/QEUykNcw3aXl/Re8y56rGtmQBQRU/U
LxW3ieaDOexOnN8KQ06nV90sIFembnwTLQt5G6ARvuUoMG24UZSNJ0VLiU+1nVtm
ofhaZRly5BuSkRkqJ2A+WGO4UtETRT2ohdejChmagKr6HQN8Q1hj1Tu48kDHFo3k
u4DE4qtmweKu6nGnl/VNCbKkosNrgbl/ZaRRlSWvJ0C4Ti86xuIXQkOjVJ424Wre
LRlDuuLNK4atoAIaQXeLMQK+yBGDtVtM9SER9jPoAgj3W4aLDYTC/YFXvivrYyy5
JCX/D5hZ/3GuuybNmFyblwXnlZdsZDIoFeqbR8bxSI32P6QFiGqI7Vfl8Z+gJ17+
A+nr6ksGPdrKCICKo8VsOD96uq2KJRIgLP7C7SMysFNloVMFTZ9yp70M6rfU3030
/vw+vSa0hWu0ujCR5XyqEBfV4rZ4O5tEBjCuCigU8dh76EEAzqKDjOF95237S7+m
Qfalm9nfhg0gRzN7gSDy6YIjjl+hjy6zkdyo0wNhpe2HFeFTYim+SjZix4nZCtQE
TGHjv4rSTVV7QiBuTu69jm/XmwYwrfce0ZNOWNCzkDxEBk2VwwILYAMh8DXxmZD/
oDQbsNWXlUs0dYj+gNPd7oODr+hglMxTYGKvs3atPDDlFjFHqmPYIt0HVcltQTun
J6gwgpSWzthJAuXiaLEUeVJBsnGqhtLZyCXn+67wJk42EPC8t7US95dGfxT+G1GX
okIHTiL42hoNKoMEV6v6LQZG0NzTzvUsp2OADEpIUmkBXNq/Q0nrdGXkP95btBM6
NGEpSlM0GJjyhWHvnUxAfKetxNdeioX8XlM9Wo7mS7NumaTvZQ9qwQVXumolfd0E
au6Zj0nBRtGpPr46thuG4oMYvQjSI6Cf1bNnHSJMhE8WdP4EOCA9WFLeyfgwVN2p
jqUvOvPJ3PL6qq+5IKMSN+CBEs5+q/qVmDvGC4aBubkf2sLuLp748m4yXK6BKw/o
3FI/qJLq5BiS75arz9dA0W72MaIR8dsv70KQR3SJO7KUB9zuTgkuVIumDq/vAwZf
buWWGCM6Apq5KPMypqTGbWEa2yqQJnw69YfEkLij2asEXeeTBw+lE7vKY/qTU8dJ
tLPXWTghqLr/+uz83XZ2cRk8bMTTPbSLylcu2tIQ/+urxR5jZ+NAtXOmf3vnsQzh
kPLjxGPqVoG/yCKmWtug6jr07LliYMr+8TA5rW/7x12bwrykPpdFO2E4vBVisNEu
EU9166XQCg4HIBOsw/JYfuSLVEelSFKBSf6BQafa/WRLk7Z31lH5NxOQwq0NsMte
LZkA4k24J2UIpj6E7PLVGFWGHHF3DzXyJfvyYymOAo2/dNMzyFQoUbVGvqMYbRZh
DS7JkMGvaZzmk3qVM/rVc723YdjKOaKJYnfH6eLLU+yXW2bC+kUzMe3GXwtjjwqX
GoAlJ3rmOKdiB/iGU/fc/DcceDLj+9BIWRD90ufJmFh9J+cw5qUFdsvKVHAvrkDK
EeF7PlW7Ex5YyGRiwLJothe4+vSa6TonYqr+osiNHSTFHczVgDpRvNr/O94eZ3fY
PJ4XC+FoPB70xQLdOc4lkaG3o84R9FaVq/5qdpi59+E8OaoOVidYiOAcP4M8MsWr
F9RbzUcfwW+oYx48qbHvj7BWC52kVSSrimpRMxcS7Gl4wVLlEDei2KWKeB3ruDDc
Jhfg4ScAHx+rj+/TsqE3ROnWjKHNhHz7Z5UIhIOFHDRvtu0Akpi9mUkB8DkUb5+z
ywEXWu2LCogngevTko6pj6H9UBeAxZjUQM8cRbN3mjZrNo+nV2igfxu/kNt6yUpQ
crhgYiyyawfAEwul/iiqemz1nr8N4wh6TG5VCq7KBkv04j/aGeOgrA8hQdX/aSh1
6DlicfhoSEjkTIFaEHI2+4jz2nFLvcm91r0mV//1953HZCuJWy66n6H2H87w6dB3
O5H9aEkkh9L5Yl6VB8zrp9ldWaY4e51dYkLdDkWQVrMVchYu7nQnM0cl9VRlPZfn
P7VU5HphhTLREuteCgrpJjSXe6fr8pXwEhMUS9wS+L5x1iKcSAsuUFj1YKg1wdCO
p4QAIlfoEhXUdlUY5za9jc98/PVZO6Z/LcSVsla5SyT/9Gtcnw1L1WoppFWT9Dqb
aBYsPeh/7GqnltcRLHpGM6QcgEeJO/Hi10cEgoqzAELxpeS9joZgVCEanewf7Inx
9GB1zuuP9F4SzMUb2mlWL1CEe1/MKLGMR2WN3eTRmPuYeb8apoc5kKzYv6dm31LO
Dymli4e2x773hMQQvBisi5LQ/Q6qLd1mfI05NDFASlCRDSXUSx7uXi25ElZWPk9d
ldnwfxshQ0gahPM40kjrwfmxHVORLKHZF3RP0NWjJhi4im6Hr5LhvKx4f9SshFJq
QVkhyHqFYsrhLC6fmGb4ARmk5HlH/MtMA9VRwQoMlzesS39Wn0nH1Htyb3epN7qO
VSRIUji0tuOJE9DS+rrXJ5ProBn5Tua415ov4Zoo497erWJMSrd/CFyeotGtYv8z
WEQYJlTYMU23CUvt6NbTJfAfQeYTnVajwtxMSPD5FcYaYU0TmTCKmOEpZ+vUL963
cRWM/F4+Wa5kzSy8p2qwNOlQmoT1oZxveGPnRYsbRXWhejs4AgE4mrnqNYCTNUjx
VdKG3UEnEC+9UxoD4XECmDVNOGA4++HTM8kVrqwJFnrKzYBFN2NprfxXfWVokeTB
NHM0H62SPOfIoJ3KVll4AUu6fM6bG4RSG5LBz4HVUGYisSTHgb/NbFQeHuS6wQul
A6+IRKf+E+ikgZEzhnssYSGeksicW0RvDu4HILGySjQWfN9PuwQibTtMAPT2WX97
HQsMW79GlLWhWAaRRhltObe9QQFfXPwOJXpEh5JnKgdXeCCcuEDfPhwoYiGoI0mE
6iADEh6MRAsLC35CYJpmNuEXfonDXpTYSU6EC0jsn8FSy7oY7hvb5cPxapoKyclK
5wg35CFWkHcIXcHUSJO2KFflwqiVvJonpYf+QIRDnzQoLpfNWjzeAmvYWigjVXCb
hQ/ttMnxEQwhY8tQRnjjkJjsqjxnFbboguRvFn/wAkDoq560i8TkE/9geI6JTGH3
geF9uJTGYRsDQOBw+OdOmvdYVdhQZOTOlLO0nnjVTyRMk9uYwQfMwX9kBGAKAeGM
KbK/vgrCzEL5xkPVJl4kOclFRMIyVAxXqBkLKzm+eQCa8ITPayJ2z8q1o0Fwsbt9
hFDRS5XO1eKA+8MAoAPabDJE2vrkm5GbU+hWgAqFXGjL0t1WW5FNS8BY3MpIQsKb
bQHPZeb71tZpDIYs10GliCXEGj+ARQS3/fKN6Xy6AM7wtWDX2YsJmgbgFsXMDsLJ
qwYbWao9NYZTxxf+m3UNdoXWRl1uHQIspvRr1DDf5q7TTJWNBNcZ1vLlr2jRbVA/
atuDldoB/3XJrvCNA2bFOCXOofft7pKlXm4jTeGeahbdYgpKLdQ5Cg0YkenLg9eT
QaujzXpAEwIzNt+n+y2Bok5X1YAcpr18UkWhdwx5tRFPRg9h++2c9wiVRsFiN2BT
856yt0n034oVf2VqfTPwMjikeFFwRQ0KyjdelnmywlTHQzhAIXn0jQMVXEaPsT6u
0885YYH/7faaultF5nnXHBVR1VV1q6FW8gxfm24inMMaU5GdaelcnLoXhgK9O9kR
P3ZIXcwCOVqcDhorKAAWNSs7kQONf2QUxyLYhjTs3JCL8TyK3ik5kXefhOEZB9k7
7ceGbJuuc4KUqp0ZSVe8poXat/5+d/Yz5vcBuARA9TRCcLpd8SmRSvpEdzIk4Etk
pw1xoumUjXXtpVPMPsaLWetkBUqAs7DvR2/TKVb2D0u9MvM2s4P6DmCG1kRVDQnY
FTT3BH55EvBqgz8KIWkPScXiU9o42lfASsj8QrNL0uyTGLcp7bi9AVEgeCWIeV0B
jnnjRcPguQPFnrYZGCyvix+h98KNTG5bfqKLhAM0+OeP1uVMFqaKSZubV8IrVjo7
eTMuE8BRhotW9hEJpeDqfjKyJcWM7NUQ/x8Yz7SfEamXQxkW1ksie4XEJvUQurxn
mXpKArGJP9JOWiyKv4IdbRqyIleG31eRBYdNBOx0JvWDwlor93qUt1ft3z7xobaj
UWRqcLlncjIV9sLsZtyAlmX8qRSfvkGL6OfJb7SD3K6DET/q7WKnm4CZbahclbxr
0MfvpvkstD4WnAA3F6AONgcBsEAU7rwFQRYfwuJbGJbaVDHyLOwNt4pWKpiaerr2
td28b2DEqGW7lcBFQ/vSk/OfbrfHlG6JVkZ+xphjNKkWpCThtkC1WnV+Q9RMeoSo
lP3HOpBnqitl3suIV5aFaOKE/mH19TGK14lnH0P5HQvXWve+IUqyfBNDI7PqzNTa
Qwlw67c0CR126Lg4V7GmLbBSFKpXyvmACjM+A3C2/5kOXsUN9maKwBBylXDyJUmM
dT4tN7iEnWmeZai4efV8Cy0QOOURHkbmRK02coPZrlaWCr9F1TQEuKLsUP3jJHvS
YCdm0tjIhyRXAqwiOZD7GZiuc9LC82/6Rls7YdQXkNBM94xr2i9nQ4A4OUUysf/9
atXxlrtCfTUPjscVgSoidgOSLGmSYd0ZaMwlhxiIqQkb5KiaJGdGyh7Z8y5gj6Za
amiS7icnpW71yZCIcJ8KZrUO0jhlsh9PAIY5Pfh4oEt9B5wdhTQCZGwB3WhJWOwJ
txRhhx3ClF0EKQjqYLA32MRbbYFuTH1hSO+0mu2GlhGiDeRG0yts2p4aUkQUX1u9
WyF5M9IJvUUSQYM61foB7rmSKJKCD6bxERMNGLsYWDsNx14aSiN7uzlDujVanX3/
MDaF3nldEBMINDapdheEHtL5ADc2ZUNLmm8hNRMWW9jLkvt5JyQqJEsMUVs1qk8y
QyRN4/9ldWqWCxlsmM16ytfoLq6xPqrcUIBfGMoB3w213Bzwd7/eQHJb5PcJeI+W
R+LBK6m0Rui81bVys2WXOsbn8d90hzAWkPw2vHzsZTXKEcvueO6ouaK5bHF5PQEH
h4XXwlX0EhE1NOzOiS1idm8Me1JKKN8nvjs0JSjhv07xullyovz2Ao9ooJQMmHZi
bTX1xTv9hq0O5tSqBchrtv4g0KZg949ayvbdl4FU3H+CiW8uL0YOHofwjvlInae+
B3H9gD9O2cWKJeZGa833fN6WyS8rHTYBfcTMv6xQ5y30FB7wytcb/+8OBmgZylxp
CjIznQmCxAIinDkGzpR/6YuaduNL8f+GgW/omsGq8lf2VKtuDsKheTnBBPU0JWYd
Akh6UP17W5llHQPhAlp2Y/mpNKKmRplgkEI93/zwsSWB+yRwTLuTf7Mv46fOa7wW
NKWucacCQoiw9jU87zKFHwapyf8TnhZa2T+lQ15koJuXcS2INOuUbhs2gR/gSn7z
adYDoI4vgsWhNWs4Lv6sVU7p3sQlOk3Psi6r3+G0+Kv0LYrySr3if4lECEa6KAnI
9c5Crz7ngj9zvve02dcplOGH2C3LSJpVL1fgD9HYPwaQRpnZDj7jvU1O5n8t7b46
NQCO6TIge0tE/wR8XQQATk5kWdnOXZ2cAcTsbM3jQTHq6vHefAZQeKdROViresXA
j/RUi/L1YtPkE8lgUG/ZffjvwIBC/CQk3vFE2FRuVhaODvq6Kb8kzjP/vkrps4++
reAHPp76fJ/cFa7WmUf93Bu8IuqeVADdS9fHr4Qe96igNRZ47bFtD1A7RjO8Qnfy
PhHFz6e+RQ/6KrHeZPrZfhwVU3XQCrtpPXJN7xS8QOqhEn/J4EuxGnv/C/cQ5FN5
VHusWzOUeAbLIzeCf3rnGfuYgC9yYANeudmH5wH+tVZLxg4+pqGM9Aqsid6QwpdY
YgEN7rnbn44gWU3OqPrOR+BOflsOo2GyiNaPTcJoy8r/a0/NlGwb+w++jZhQq5HK
xDzt7ONnJQ5iQDBTuwkgE6BXtc/JOi/cgb4lkaNMShh7DUTFAdskmIIr6o5Zp/7Q
AVkVSe/+n0Zt7qyhmikhWI/Uop2fB3EqGvuRlSz6dBgdCbc/b1EVkhLyozEFPs2Q
vI/4KTY3aNpjmm3PyaF7h0IAEK8hCZioVtI81D5tOhU+ktcqE1YJenatHzp75NTU
XkqT3kDkcKL9aDrVHyQj+kf92T2OcA6GEbJWWKAC/MF8ahLnUQj71w136ZkR5yQs
U6InU27I43TjVi5bsstF7BCREWJFPbDCTws84sSTd6632Vxfx+p8BJVaaXWek+O1
5WD9VZo6xY/v74wtCp7Mga6PFdbLhs+3iT++dU7/gPN9b+jWI7iK/ew/nT8AJ0SC
3uONCPOv/cFgB9JVCX0pamaHiTcdsUVLnhBqX+beWUhp5dbbEdL2uQQvq+m3uNBJ
46mDuoVOV4J3Ul3RNITkh842sQIXsgGuBlveGKfEn9JBgPD8G0bouDcz7XkzI0g3
9/6A4ZTnPzpVWKBahQvlkBQVlfQ7jo6NOPu+wDomw2YexVxHBeQleQjHljhHNwgj
Wa2iIda3cmbSRVGlqePUm2e7YZuepDnV7OxuxxPH0BljWSvMhWJAf6dAgpB7TD46
temHZ4cfduovrRo9Z9AL71GKRT7MJSaNZ20mwW4a/elBIQ9h4eaVrqC5I0FjUBvb
7v0B8BEDh+Hrie8A5t2shUAOzbjGPZkZTIe44I9SnJoOtbdsqjORijgwTGasNV5U
pVhoHdSoh9GotIiCfrWuJzV5dd4kV+kzdG+ywKrJE8r7N5aR6GER0k+ZAWbuRD9W
s8uZ5Uco6JuLK8MrMoyT3uPgKWmA07ykLMXDu+R5+3kfOdAgEs4Ao46d97HrF3gc
UZVuOgCulXkI8cFIYI7wRlRXkN19tBR1g0D9nuIE3F8/Y+97FUji0lvEDplAlpWe
ynPndSZiZe4wa2xl/Ob1mQyUcjnMvu+EQq6PUCx4SgabSmNg+Tq8Httr0BOp2Fbs
ZEjPddD2LIpMsnMQvEa4BHt4/cWwMHsYQ1p92uQZo66nkOiplKVsi0mO097EZ8xK
ftv8EpY86u5L29zTJcAR9cqP3nAxOBC8s7S49yEL+raWEy908Dqtf1vGHgeb973j
cDrNg9IhHuIYwrJBnVMoGpXHGRJ15cidbdxDEWyc3DCwPICIIvzkSeX5+feTXUMR
HvqX1YwudNb8wjIyOyLKldThRfd909i5+uW7WbdRqe/ClnO8mCHu53vJeOvnxKvk
2Hd6GoId00zVls9d6LXiT9IlzyS7ZNf3fL2TYyhE8PKEyEIfeI6xn3dgTvz+/JcS
xI6F8WfNBGvBbaOl68RnSLc3Fpxb+8D+Ks/84jy0hxlDO/6STRZpbRzRCDWI/BXR
wATGzBQTpOEc+xsfb8ORbaPr55VijoSWRJQ6WtA5vZcNpzJeVpBnRSRCYSg7Y6oq
Kpwcyo6WwKUASXe6DNzZchMxHNffDccUSNpmq3B7ozICsxzpmUgG6B7UvRt/HoSC
yy1eecMuGpXJ8PkgOmL9PHKvhKqg8pOOk+ZUb37tLBqyx2OUz1V1IbY4A7YVCocl
aWLXghbUteDCQm34ak2rWUmAqDtG9qW3KaR/7QkyixJsxkxlWceuGBBM/MCPu0kM
oKWGXlN9yVWhtjhdXm9dFi3wyAkpjsWjWFoZxfA8WB2W5zekxcoLFEe4ICWB1ikH
zQqTGnjZ6UgRSJKVxL8kQL9vHcUCMLADvW9jC+UboFXYhb3/ZCFIEtbuXm/fxkP7
5epmnfvdwXyYJYxT2uU6aKxGmbbb+nYvk9URQnGZeaejgwds92PYLcwa8F4bpTio
OmuWbNjf/pqRULJWyP0h65LXE5HF0SZq/Lxq+SmpgSMYaiOlOKtNX1txK7wWq317
0EDEZvcXdjcf7wfWWrDrGXSm19VovQ1yEgFWImR/dxtl6OeCR9MGyKc+Yws+v6hr
rUphTDO7dEqrQ4vpRAeuCQpQxyOXMuwzQPYHUffK2ds/O6T5HRgHzopN3kDTBqyB
OtvyTKPUXXCMNx3Mz7rGaDYALwRbrTNRAI1uiE2hD+EltcVlyxMgUclGuc6kVuGG
HZ9eNh+v7BIcZeOR+5zr1mQXwK1Wqw5sf/UWZBldDRbV8rMil2ojG0mxY8KjAwQ/
7Ds1NYAn9lhYWpFotcDFpcIXKpKL0e7QfOdXA4lB3N71HVABbUzyiFzNuRebut4s
g75Xq41R1x0evRXcA+zQ2IyciO4ajk+GHut4Or2E1MHKb9N7QIJrnriKZszJirby
XM8qMpVuuFYyFLzLTlpIYODrTLQTmneKnPJwC5lT5tEhAPHAHweikbzRzvCScSvq
3sT8zXGZ+PKvGaBEbMck9UNsQgFrIlDgftOw1Efsr/u9SP3Et/1LvbxFrdWA9458
47LIiL93FhWp5To44vMb836R/paIreUqsdJeDVTllFlMfTNhohwDcVeQ8/BnIxXd
qSbhO+/ALHNIMg+Mu9zp5ZfsOCF0+GOxH99qV1i1Gwp7Juyn6IApljEvEoAdUUYU
w6ngAUz1PzKP294Q9utM8qduUfckNT2LOBpqmMhh/BEl4MKTQzu9Uwe/NnFPpjVK
SyFp3ez3ns1s2zTPQ6dfGEIualLpphVsEZgMFUNbIQL/L5QHcpc7ww+5Q40VdyqF
Y06fhXX9uZij/cvsuzb4m0F+sAOwKDn8ThC5cPq2ZruLv9iA9OzacRR30gZFwBS0
+eAhf8XhTGtBQNx+i/b8QOCWZaj7/45cKd0zkSvlyznuS6UDqhWiehAeE0UH6d2d
jyy5sDj8NejUHZHd5gqwac9ceylcciwI8hdnRlAO+0TlV9BDURFJ4BdNLe4I5m1a
uJbF9PbR0ILk/CAE02GyBscbKLsLk0A0H2jmmt0v1jXvb23S3f6jG2ZFARg+hM50
1W7UERcORYG8C72rLamVIYqGrudSujBv+JZ97QfDrfAxiGOT2KCmVL6yvJtHZQuO
4n6zOn56B+MttnCQXZxqtvhQdjUFRN/AxY3+va4NnuTsZhIOwXkbNkrVcdzZ+W1u
odcqm+oV4D3oIFDhZjvKHSQ4r2nLkN+TT3yisMwdC07bnoOis6nJaPU86UMoQuCT
VbdvOu3j9NGuJAotVpuCVL/0+5MGGBD17Bplh9xi7p0R54DtUb+S19eFvh6zx2hn
hVoTn9G11mDp5+zef4r+6GKHNtmW+sjYji/0p4H/C/e9soXjwEOD2r02HuLqB2FN
nsz7CNqgW186xAw7nImVhA/cnhPNplbFQwiTcQ09j/UjAkvnS92AcLEsEC0aBxqi
IXUt8+jETHS+P8u8t7MYsov+OL4lVl2vzWPXBnpCBPy/6brlz4ZRhErWmC9rRL8c
KdgRyWzgbDFJfH2VytHi9kk4u4ts86CsCCakKf4qCFpTHqqhVu6io5jsqlA62BvJ
oQJNUsUtAnDf8HQuPcD17+T/v0BeenqgxiNlB92IRCBP8hXBcrsoQOzfqx6Wyopd
T3wwFYy5o4qVEjU7wA4cE8MsAaSaHMSWOA7UfyDa/ykank+tzqvOOLoB0T6Loiqr
UxFIbO9AYDPkRfCP3dgAeJ1ILt/mtxOt//DrANg7migdRjCtUtGIyczpRRRpX/pP
xu7cnigl5Ni0BM9psTp7cbGFs1RR0cQuuGb/L6yuE5xkcHOlcIFADOCbJJzGBmI0
ftUkkNnZ7VqIeid9VDU9uahdSxzfDbV2YtAUcpdy+WjZW7b0XA5fsHdQIEJenQbT
0EbxIbMU/qi8j64JDGlbnsOFXjjOhGnDYA9uVwv0n5o1ZKXIrDVBY083a81EVwF3
aK5qJyMxk6WARIi/I7uDegm+fZXzZB6gNLoDjAK9aswvFPvVnTscvuXLKM+AyH1d
MTL97SYRGJcrkqkg1B8A1+gpLed0PIF34il9oTZtZfPS8OIp/F7UcfkTVW1M3GsX
2mSsLaG5vqNy86TWpfGxYnsbqVIGtUwUO3nzWBADY8WrQrbvV5PLe6P0/F1KkQIK
1Az+itP+FZibw9JneZsRf6PVB9EYZ+ki8wNG7BsKP/hJ3qbJsGhA7+ULB1tmVrUO
y9vcG7BWS9MQALAUpnxhtkku9OZXLPJHSMv4rTA3bcyo8mQ0PUbgG/Ud9X5P5/ko
+VkHfw15iLLciomnm6SFYqPfqrDYH1LDe9rb62pCfbIq0u89JNPxviJgYCmtTAzx
e3IbXlHfNy0uCLCmbU7uQsVx46oEd42Dkb4fZg8GaebLTlYn2wxtX9ExMyw7BTtJ
hRgTM8SGh7WeeQqIkCYfzbi+3MvGAxyK4b/ISpX60uu6B4uXEOXuHjBTjmW78HRP
oqdpOBpEXSKMiT8XMARMwX7e7l7KO+8lE0XRqPVFSqV0ya6gYsk6/2nvz81Dw4pv
Xk3y4ksifshn+k7KFcAZPi73GpU325B1Wqg5EJE+u6TlGMvFsNYB2VK3okmWVkz7
UalHsB5QfzxD6MTGjN5PDcMQ10SFCUZTPvisldyjFr8FiXcMffJlsOHKFVHLwjGm
Ci8Pa3ZqGwYjcf0zKk+5thlYy78XwYE6pVwdq3E/mVBXSi+xLBa/b/J9I0ac3cYs
o+BNcdRA8nLtc0VRdN7mTiVhlVCsQKzd+1bzlYfeUy/eL36nRNOuYDyCAGPKb0uk
slUYiP58AhDoeitv1ltEGDzDaP/s+NDxMHtPwOhOYstobcfbCR3p1qf7/tvaZm9M
reqQRl5eR/INd8VPwGXIYrewEIxPgRjE+dqsIVgf4y27H4y3dCniLRKSuUy0dfjM
fz8pCHGyTscUrjSa8jg4fwj8AFYrXB6iTynrnYr0ZFqYu6CsTCJ/HCw/hvTXqsEu
ctwoZiPllYBGxBOSNAjtQsmQFcgA9KVBW9KIdAgvnH6g4EwLyRCLehPL5WyIdAjA
+2D40HGlMD7cY6H6eJpVgMOsHCSJ9a0tDl4w7MCWnTiYJ2AZQaKm/a4iRp86I1Ae
dYV63kl1BlEygZ1mU82hZ7AK1AMrZ/mtcySGYDnDRl+nUR7K9eOmbK/BuSISpN8W
etXirP0/0bV+Y2WrKZUSjztLbOsvXO5F7eCVQx0PBXWjJH462KZKn65OB1g7/5df
3gz61qlKwIVIeoECeeH5Gf04yNwGqUIZBt945H1ncf43vfoOyhxBmamDmadpBhSU
HpLd39tt0IlJXrK8y2ap625tH2iy3XPLiqyfFkRZlu71u6W8wUowkOFcnk6bODyd
sOSog8pfTyRdEmiLvWhWY9xDNCQiDxq5g2GXZ7JfMGxf4YMjfZkvdFwwnIF8KnWq
P3FC8fzMLARI6clZSwpUkxubjg3cVy3ZkkLk/QiUVgMXuD1qirD4G0jgv7de4DxU
94w6ih2S+g4+RDv+T+BLgCHF/T0c+HntaQMz891qQMkYGx7ipQmpzjZECMc7QDCq
lCGldGlKvHborEsNVEBUdgMax/49T2U90NJPzZ1vrrZT89U2SGpcemgoJXyhGEJP
sfmv1D+6AjtZSL6m9pURZ6srS266QOB1BmEEGjam/DU9ag4/vmUtW1JZBwN/4VkV
XchTw2XC2rwBLpN8DLHXkti4m8/vqhOm8D7YrSJSELBHLGiyA79phZh7umaMEitr
yK29WmQZ/tBLDFBADjoFSFvUY82Fz+Wnitd06+EUaIYPicsjTVfEKpTFkyTc8fGb
9Zy93BjWygxqTecBWqZWZ+if9w23mvGFXd+vDinPemRfqeZyYoGkqM9g9xsyDXBR
9gSFpJehQ30YudDaCXJrpu68WyvJX/79/WKuy3NUGve6TYnPTOmNAzYHGJX9tbV9
ZlKyYj40i3gukRSC3/jdnEyMS1i5C+P6rn0CaY9ELF5h/9nk/RRYv2ZpUAR9DfQw
qb7rpoJtqrZhVOn86cNxc9/QuBD58UkDVIg253bJAtIBsZ0BAikXKxaBCSRNUIWf
UawBUFWZnd6KetJah5BJgouTHicH8Va3/wyB3JrT0j6rP4ia+NcCYOktBNO5fMNT
2GdQmK+By39/hj7/AW+EnjV7L0fjId5v9s6AsSLNTkWq+Kn+wKjYXOlxT5SddeCl
maqn0h64WJKAHIY30OoKzOyXWesFchMEZUBs628vYwjh8eetHmNkDJfgo+GN/GR4
CJJUscO1Kyrw3/emIoig9zcSlSVzrJLcx0PhePUbOjhu4/1vUhmq5y/rHb2cjZT7
AdKYNYBO8cpq7ai4phXmFmnM4hZp43OTNrCBCuDatJd9vLcPoyJpuavj+5U15mM1
jut1hww5nacyp/n5EjtnEt3nMlt0qPf00e+aIOL5xOcWAeK6hn4Hl/AWrsqnJXoV
RbmP1yiuZC+U0nAKaPsl4pXDY/bFj+YtXpubarBxwDPLjD1lXKiyFFJucCHx44KA
uMYlBCOKCDPgusXc9jG1wYfzDJJNqPjcbjnPMdAkBuZgvjcRFUTMcC1omj2TAyLY
Smeor1giJVRCnXqFlPfOO+OeRr122yQWPqqj5VEA3sqL8T92K98+ADWrqMxjkoVQ
lQfmk8Ssxw1v30SYzE5NdqwHOBj6huuSOyRxOTST9+9KOGZ9laIEsloq25vByEL7
JOnwoAIR8QocOpiTzo5xFJgxBWREoI35NDFlPoVloifqwKc+n4kG2vkMJ8VNoLNb
22+YRWl9DCLNqS371zsjQsxXFJaa4whmgsDxlWCwabEXabGnebZ2Sf4w7V5qCgdi
YADKRc/kKomZ7FJk5ga4htHSUSI0EZrV23M7aGbWQMORhfHlcWkg86SXGJumvg71
2SYZn4xJW33wzYS5RR2lN/8iVSv/Gj4+wEFKUmd9dPINzHUmMjliY3/5KxGGgqas
2DZ752Mebo6ouM6I6GYoCPbYyBTjHTW0I1N6qoMyGzL2ZxDWMyD2WuAzdtGuTZyT
g1AYlVYfULkb2O/m44RjqStMaDv9M2/BNUDH8ke6LL/PGwBviQy4pUT7SKj+Ztex
XdweJ+yIX/FOq4GonhrrkOvMMeSjGxxcW/aSnJyv85UyQdWoR4TBWtEJ3hYMIQmC
reYQUEe9IbLoR2hZohesRGwIclpv8EOqcnQjFE5sqdzCDS1t7En5CoiZnu5NfJ9D
kOBebvrw6MgU1lYL7kyZcU0bvf9S9NIMH1bZJFNI5GxGDuiBtH4Trh14zMrXEzoE
mb78B6yyKVvfYtKrPQbrkID2uvISv5Q2WhUSfz3rGC4bXFjkKSrxA/gK4TwbN2yL
xtN8FQR08SBnNyQmm/R5yL9dDIH64DQ6kjtJCKJ56hxZKRgOfwmQdG8s21T60UxP
p2W7cLZLq+2FI/wVgABYFzy99MS6TuYRUdyVX4pI0TFHTSNo2yBgdXH8dW/KCDes
Lf06BXYaPSVWmJ5IN8QhwpUMimzNHAuzHV0j33+OT6Sulow8Fbg4yjG87rcwnuDY
Tgvkk2nwGPUHHyC1dz2q6m8tjTxGyCIxCPseEtGBOrjZX7sb4GTdj5nhdoRy8E7Q
ocGFtZB7bKy5ahryOvwO/A/UKm/khBgB5ZnozAhfDzlMiTbSbq+3ndv16heyy6qV
P8EP+2wBjBoehZoYb7j43T8OJCi7cFKJ5d3zFD3xd3O+nH69EdOrLLpMQedodZSZ
ytGIx4a0DUAQCc16yfcfUTOxP46f0Y+FwiiIy3jZ6XejkQ7M3WlKpdJ4vJ8Vwb3b
QP8ArRgagWKJ80qGyJE1nReLBIoYagezsOION9hgkYqXeJhT9kpqmeCxH5UL4K94
dSdaqtNhMnhW5JW/Q6Bmw1AYVuFHku7tVW4JLO4Cw1K45eRqFf0d/KtgM7XJ3GNe
XbtjgBISlzBKwF4/A8UwTOAWAyHv3NYIvNSyi4R7HpRazmeE1duks63yHt6NziHP
EfX2c5Bu/PXDBqMWIYtSRgyQ+uwd8yxDzmm07izDoODeJCwm9I+0FbYXz5l5YlYL
3giCsKHvD+aHY6tDG1NfdXNWXrr1hBMat4y+DvP7k8/lf0vX6ArXfmJLPFhbESD/
PxMKrABzEe4yHQJR7wOQBD5zytoJjtHHPaLppCLZex3iyrQybZMRhkuEqTca0n8V
ZvUYvvVyFwl1Z2cejanQ5ML95/R4tVkw2AiuizapEW7FVSLCMTKTHtBVhi5bZapD
kTWj7wz46eQ/E+Vdq08RHFgNwNBqTLrYKdU8PuG7NkEu64yOjg7ZkzCMJUujwYnp
Py9DllxQi/w70DXSNBOd4AP/qfaal7gaqTByN3iEeq8S72mDqqM0kWPIjpZPy5jE
mkjyIsV4MsWjhrFd/UWNrH9UG7tC7M3Nuy3fX/OhwT4LhssaXVc3FWqeX6WxctWm
S5I8XRahcLJd8A6NUEfbIrikZkEPHONIO5YGAXb1Y3OmpAFfI6HL/EMS+hl8Z/OP
kR5F25o8/KOFjAsJN0dyClqwAbOapTMs688hb85B4BhYM68ZgBJAwwntY0qp6TTQ
zDvdHcciyO2f6kTTLcmcuzEf+Ivgmy8qbd4izH1DY51SFrWGi+64rq02AGiRXRU1
c7c+W2EIOfxrRA8F6MPA77evCB01eDTbHoDcZUbvne3FuW0f9Yyl6Xlj9z2kAcOo
e2iiNYRKZd/aKNtJL+iJ7x8mMPvsuirftWyiHLQFABitHjXIE0+RoNv2ERcCRHi1
gI7kyKs5QGL0xPxf0dTjr7QsiU0Kzo1RAsEomf9KX7wqvPbabsMvCqXWchZ7h8Cc
8eBeSuhUr2y0ql7T03HhCiFpGVYORq/wLb0TnuxggAkUdX/DYauzmV1LvaF8OrFX
UR7eLqEZvIYzymKxVzYwZHZp+LnmhFl3IizyN6y0veEYX1tEeWpmAIGuiFWgeo6S
5fEh5PA2HQGPxHDHmzO4KSpbHKEUKsbhegrTBrSFWY8tbQkDHck21If8YmBJm//T
ghUZfQ7T9fIQn2rRRD36j8UMqmCI3I9CTqQLbYK5YfjR4Tdq7mqKHCIwn/rKtGX6
mt6mDT/xsUTHgLpHwRK/TSt+By7xBIxaqMXlaonC+J6w7lYfub8ASseG+qq77whG
fFgca5Its4MGUIcv20A79n9Y2Ia3jzHeLFpI5TzPOTyObaz4vtMakqSxMtDNH45I
bdSUMBStLiJPdgqcVls8Sxu00io3XVJCaZ9MXTTXQWzmfMYIB9YpJVfbncRfGQKB
GyMyppCKUANyhM54hQc97vW0z2EIEc/7tEE7wMrJNPzX1S0iJmP3OeSMkQ208Ruk
WKDBoyqvx7knsE1vutqvTR1c3lZ0/rG1vYBQ2BjBKU9ABG2BwjbMaABu6DibkjDy
+2ord7KvN0XgbdybjCzuEXlogyv8eRB1+L6ZlH4rNlPegaYa1hVBlXE5MfTGg5/V
2zwUIJ+VygW/ST+kz7tEA/YjZA9lSpOrfn9aMPqJx1edBIkmHj/I7NV5g7gvsr4q
/K3lAZxOYk063nNjg7GUZxYfnJCYiK5MOC9FObGaFqUScwItAhHlqTxipoX5J59t
NCaeZZzJ9aWNLLroIawW9sUS9dKnCjaEW3TT3TDmTVlAAKaUWaYxj33mVZkZqFvt
xkOZgR7bYUkezdc9cQOsp3IPnL3z7tPApxrAoxlww5988fkDZwwsgu9HDUHhXT4M
twHoQ+3f98kACOmrkUC6mVPOxfgPo0j1Y+9tRMVGcCqA9B1JsYAylZ0NBQHu5ygi
YexTC45DoJDfTseUNCdkRG+PKehgDn0zGkTUoKMW681VvDvj37U+vaSqgNEnKEYA
wXdHiXLLAo7IM+6o1xzlRAMTV5GLy224QUKaSRToEztXBLzBv6h3QgwGJ7oUoQMq
luUwcYVxnzAl7R78GphERPz+5WvDNUsePyYcOJ1+XKsV0PJBvSJ+uglOyX9GMYqj
M+5pVCYpKfAJZ/q3xw+up4vBvpz1hsmG6szEIf6VqPZKbmsjVT46/E48BDstqpXs
6OI0IHpl521pLBEheZHerL1gSrkJMU0LiR+3avu+jzwC+hRENQnGL4BWZCpGHtyz
B8TFOqmuts8rNCtI41spw73gw7/XLIn1Ynxvc+0BlB98kF92Ec9bUpkp2WUdN9z0
9yzHsvAvii8i9xubmhH/cSZEKTqA2JM2ZghV4x1lH8lqcH8Ui2/AclCicQDMDugi
dZlGQh5H0pl9B7oKuWHfhAcUz2dGCVC9Z1hrMDMLaXHRWJmsGkOQ8NBFUMSXz/MR
/RNj+InQT1L9vka/XU8NtNmvQoBRdrtGI4lSclWnDElFJfFN+aUe7uAYsbECazaJ
kpAssgDXy2KJQfnE5Aa9/gxt1niODMA0zvGiKusQR7uzGVmM2oLOkD37HV4Oi5sZ
tnEl4oGFWsUJ3y+O2YH/+9ygFrKFJ+PDUNSLa8J6u4CxQ4eCx+8yz86PCCZtpgdu
xmmVAS2xQI5/Yp/K/p2kNu3Yp+QUFeG+byqITyP783gzhkpRqFRzdPj7xWXBnPFD
xYpkX9QfSGYztkJPM8h+OZMNBaTfuAuZYjLJe6r5uRqC1XGeXaKH0TOPLgZwZ2c6
j3mK4Rfl7uV3wUomabWA/w6ZPLiKsgyNjB7h2PYQMKhC85+sBqK3dkyUHSg8qrsn
VPMy6r7lM6BygucWj8qITzLPgYhMGbT9iU7M+OLcoLJUpQs+vFEKqXqf7ZZxHURu
OTYjgdija9v9hw/9pM5rixDCdOGJjHvUkRFs6uGFr1HEaSOmZNwutZ/JmIEcvS4+
PQZFSHQ1PmTh2X4+sIoxQdMzjf+uEZqkfm3/uQcpXeC9uiKdB3488Brdfjm5PI4f
1cqnsSRlRSCO4ePH/UqHPhFWIL1YAGwwiOrlc93ZMqv4HwYXNduu9REz95QEv81a
hCtIugXMvNCJ07/ZQLIaefcj+egGVZtOinb/zHo9JScpPnFQJAo10KvJDebw56Vb
L3BhLA6WjJRdCCNoJLiilKmoyO3lUvobAsU1pDCqHUg2pYs86Mj6HJdkNCEzFrsF
U/mLWIB8wZlf64zxogzD1fOcI0wNFg62eTdzwsEKGhUDaSANmIMB0hBYF0yHGR4e
J/R1va8UbmMOCGbwffYeJe3Vo/r7hH/kUDWQWLEwM6YE2N2EzHp9coD8BHXzRBFs
l3BZH4AkFQ6u9eqvySfEl6Z9JerU6evxi/BCxjNwIbzsmCxmflb+aoiQSOl8Xkgr
0YDc/A3JXGpJjIwpPs0bKPYuAdk+0NPuPMTOFqmS8A3sJjy0DYZ0vbOmBIZxNlyR
exrRcdxZdYOzj19pweWWHSqkF0Kgh5fDjwqhSZWBsB73YeCRQTjcJEB56ucjvlrg
96qWI4MKMV8Y4cJtR8GqZU1qohP6pvK90cvTNfA0YjuF/71yNZNE4kQR4pDf6eDy
WdsGLYQ+Dbt4yNQGC1HQpHagShR4ikLwz9HP2y2E5qdUIACllP0UNTY6GboOapJa
SJLaOuH3x6UG3Drs2dqOVE1NVzFH4IhcJ0dTdcGTacZ8vsf0k02s/1/VvUyNhr0R
4cJxatsci2C2rP35M722JdU4z20HunQQ3FhS+3ZNN+h8V3Boj51GowYxzJnkV2Tg
FEpWLa03I+Uz4A8GiydngAQqPWiNSeNx/AGZ8yxGjJQmN8UgyiaCiak/UIl5oNk1
034fEeWNNh/9NX2DKEZer26tnW76T3fZJ6MUKEJ4CaoaI9fholtKY94UzLKz9Q0p
lvlvno0Kl0v+8A+QQpyGQ+RxMDljY2Ul1tsqfP5DwBsWhdHICJTrkxcZOaTvDtkl
iR5Wc5yYbvgA/ZAnrWTFubq6Ac7df4EYljjfHRJ5YSFd4W3OoNSIhwfLb9JMafVa
F5j+qGrceX7vPE3FSrtud444mA7E4PNH9LAX2WHkHnKFlj+S3J2PUZ25mIhwGxzO
CJiPE8qFpYE7uy3lJeOtnU2Ul22IyT+VZk0clds7i2Ycf8Pm+WwCutTqKZ3FCzgX
sEvZkzOQppubLxQeku39YaEl886MGSwehmrVsIBrO2FeqkxSMd6K1T9yhwk1aGjJ
U8bBgoQBQzkLocsix5E8R08dhZS4sMnFF0DMuVLrwBo2LpBVxHXUNDXmfPHUwoFF
Ff4z/JESpkdkqKMmSlj+iNajK4uEVcJ0CVFMfaFOeyf1bKY84OenX7k6zjVC5dl+
y/H/WQHu5S+XJ6ZsgNeekOxz/ZtYSVKQ52WsCuYyZyaS4EEACov+jg4zINCh2Etx
rzWUQ7I5ez1mcnrRzJP8Xj6SaZTrKaWi9b0ALz7TSkzU3IpJELjn06GwQtbqGTXa
9h62ufeabaUX80NUcplTaa+qXNz3TAkwGiuCoJk+Syc+mpVDLr3/Pj7O2N6fX1cO
r6ku2b0dZ05op5YTZGPnmW4mR2n/1BrM2G0xRXOAQS4RkQ7JDhoXTdpP3U3FNkZH
4+V+cxVG9CKC5ePekhOlKxpV1J1LZUG6tBFB68uMOSmTIa3eokLNJbyymdkLNEzn
m+FsPlkFYA0+ZfhWlDIbXWlfcxhCYb22d7RLHOXkoq8n9qaxIhAIGzuxkyO3pFWf
n0InZMdcLv+n1EBHusygbICj50I+u+88C/Ds6F3HZRrIQQigC/BRzFRR/eQ1MoId
6PKZjYzYt5TMCYkjzODm9ytKkSXO0fRXpE1ypDJQdLHpK0BkTHCMRCVInrsVnSzR
BU08aN31O+z9dJbGwPSRNjGLW6ncmZI3uhLGQsZpiEnxntoAODllEx5mYl+++U8h
+RVqos3+Eq1gF5eJ2u7F6flJo1Yy9Wn0o2nDVIdV07UeSLN9Z7DOcoQiiV2+dK1a
0WwqyzEx8O7bIZq2+BoaJGFMU2lj4Se+0tFNfOk+/UxgnHHd6R9z4FZ96Je2L9a7
Ti45zb/ln9PRbP50m8NVzxNej7olmk+wvRG1K7tqaBCV5nYIMEqIEQ/0/h3IXo/k
9LGc4v6IbscPTLB+hVRZadq8xBTPPPwrTJYunhYhJ1j7jS4CqOukEC2tBY7w2YMB
q9ECZNzqL9/m4hS+HaIQt+Yid2vdSULDwd8E55Y3EcpjG0r2VZrn66LL3/UCOcSh
LwqVKQnO3n1DBkSTcQrQ42zcx+0gTzlcTSb/wjz6KSa6c2tgGG3qEqLc5CNULN9h
os5xBl+QlwDOZ9Z+Riu3NEAy07wKGG213Ts9K/q/XtA6IAy+M9vbOouOTvCLvaNR
aCeZk+ncW9zLCYcAazYASN9NQV8fPeojHlwomGH9hfRSuvcxzKrR4nPOjVJdltZk
sQatsil3p+gCFcyakxmd6jAy3v0p5OAhfFZ+OWRtSUGqDuCTqLkKh7f+SdDYOX9E
nedCtGyqw9haKJPbMl03XFCCxpzB0Hdjc9fOubBrGofVUXFBgLjBhhWuiWHZy5uF
VS+Ks4D84o2LJ2VhFXxfMk3ASGeugOgPiryaChaM5C78SNubKX6m5SSQtqjf+0W1
ShjnOfg9Gi25c/oGHaRX0zHFnwRFtIzo+4lYPUfl6yamDyG+DvczPToOO1IGeDkx
zWWYeYEInRQQ/Aj2J1vUMt9XaWxQjvQpP1N3RghtqwDfTou/VLN+OXtkc67XELMT
YOqy+Wg9YN+I/WeBEW8FLM4LRaASvr95YQ3t9Xhxxp2K7tev0uV+QnjSWd+3SgAH
iAodZwyEbNESmHoCINFSyhqnr6zq/cOI6Z+VAOOJFwqt3vy0WuRYzisoWJnN+v7+
FIUWj1xkhCCwMMwLStLR6Yuw9a9Z8yAnzXgexZk6/OUCuMzNMVoXpY6PAGykTrvl
ZM1hmX7EenNwyx4a+ESOF/hdl0FJ5P6QQFT3p2OpWG2fk6tS0NvZ2ZcgOBc80gxr
H1O4Mp/oV/6OgsnyJMGt7w0Uf+5jzBCuuvKKeYXvs2HIBB+gj5rj9qqBPdYmp1rM
4T/g1GqyQwuvXvu2jiCTNhgwgMKloZaH0tcC6m6y+mHGyDFp1HGXAKNyE9e9Lo9X
pLkxUBGF6HAuCYqDYMZBFcqQY8KttNccZcmcCFGIx8JWD61oK6rjjpakDqFfsQQY
RkPNsbtnfbdxzSCkxLq1qbBqcvCX5TShxCJvhtVQCQuESsBZwbbPToHbBYZPs2ft
ZZuDqA8eYm2oy1ToYIzRa3jKlBrm6JZXn5oyt1Mvw5ZsRs4PMNbaLRY0cecahJiE
a5Sm5MvrTCL6FwRjXtdpsb1l/mzDmfbCyYvT+5KPJODu+Dc1mWDB9v7EHBLlatoW
nChVssdsGooOLodXo5PqvTGSei8n3VDVgSqH46DXcgiPq4m678St59eNRmikY8mW
z06i7pm4IryP/c87Yc1fkl9tep9uyrtUHwxVKbUYFldJSQYFnD4JZ7X2jPKxmO7i
TBDzgdbxObD6vOr4ijAMeSepFEREDEYMWnhYHm4ZBHni53QtTHzkc20jSMmUIVp+
aW5a+z3kzUzSiEY7XNlpc48qzZBemEizqPKVAyjv7rA=
`protect END_PROTECTED
