`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uC9cvndAfewEa0bKmI6kD2si2lS4tXPM4QUqlVgdMBwiMHHrU3TniJuVlddfpt5o
wv8dSdqu8cBZVQxFDtb2e4WAN7BpvF19FbB0BDu6wqSUvIvR7f30VAisR/HVNWPw
JsJvbsSPcZHUQiHD3U+gmO8H+gs+T/9fWFk3XdqzEm4oeTDSnVyh1eH+udgClLgA
ADAWe2r8/WPBzWgWAq1b2jykKy6kkEfbwcBsx4viU1QpJ0N4ZiFIR0DH4u6uliqj
OTa054oeapDLini3VOkweoF9Q9ImFW2iccOO45/KiIu/x6GdMVSHr8jP8W0m2pMy
uJM5RcwPddBaZl65p9c+f0P+XbiaJEBfJcm9tmdpms9r79MBxh9PZA+/4sykKgcm
amVG/wsz5tbKwaJgjStT7nAFc3APrSqqGKXSD9jnVxDcBKbgxtGOJY7o4iD+jdIf
nTVBAd2uXa2O5YRybnJA3zPuinEyig/5I5r8VPbbh6XuTIr9vBbxOgxEycZakOFc
vrDOQpN9By5WePQFpoxaA0gYmfh39w6cAoSjMXZTl9lmxSPluVcV/pwR5oXjNEyz
pYMSeGFzxXRuSrHuli5kTsgglumc695KMKZjG4RmjZnAr9CCKmMqPPh2ABVcZKUB
zluG0LnDsJOL2Qr31E40zEvO90MGBEekqlcfVen2qs6Ksnw+Mfe3sHi+N2RgpmqF
L/K953fN6AErQRJwdz1FhS3Ocf6ukUgAT3o81cjxiW8z7mrOIoBPDX6sa0dVWywJ
6mRp3wt0gr3x8mHHomrGypfsdUFF8REvNfH60o6vbGxEcsgYcMfsmFqH4z0dgBuq
evMzNjAva77ey4EhASyKAVHeyRsP/XMpA7dWmXbnPJtP1Vef9w/fkKtv+tZvT2YU
GRr25N0Bz9Lr46zp/MyyzqaJk3AIl3X8e7JkUFTtdGJiDRjv798TVV6r98ClbSwy
tJcLMjRZClkvXS71XKev3iinLYdG3UUNMcwyLjSe8qLeyjT8fu6ctIMOD7rXKRFg
O/3w3UcEKHBCYIjqRMiD8MKRbpIuHHDpnOlswffm2bYxxE2yfGQeqEYlo5Xejaig
HDlAJWSvYpYwyqyFBp+7QpQmPdWvYJVVRMhrzRfjJ+dlOh+oLJjZaVIfghwUhJna
XwSqHvHTK/BWeoygKnkjVgvLFJdjW9ZTS5EEnV/XnWckvjsOkKW/7jaR6Cn84Xw1
WqnCYgNwKzg1zBIGxr3m2Z19bDxDTJ5MLhW2HKDehRcB0SMsyBZHKmQKSr7cVbLr
E6GsCYw+wUBdCVw+ugjALoo0ojfuteRt0N7XftUVwnhnuUc2Cxxt/aGNGqrhcrFB
jkleg+rEtTh+HVL0TTJEtvzCgbF+UGYaY1p/5oWnFKRjxbM/EdNvhoVOTtha1HSh
M2jPpjQ/bQ1nn7E4IwECXQQItRUs3KSv0xOoQa+PE+x8JjuXAqoJQyW5RuU5KwOB
swcVdbvNpGNiSpuFHv+pOROllh+YJxV48RQ1hBkZRDJMcTKteZINZ472lQx7bZm0
BQjmtq78FcZ0G+surg8hUoKskgwwtXwli3uLIgEFWeN+7p26CTQJPiHzWNyf1gyk
`protect END_PROTECTED
