`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0p4G0k1Q/KdQZvNHawcLVmM7lb8rE3483u3H/KDwL4GmLhi8YIZzDqUdr770cvlV
n5zHS61MNlDWQtTvVSn3RTz5FQT2IJDlW2tL9JEQZcLAqECp/d5m0apQnLJxSLp6
SUctsVRkDIuANDBc6VLo+P6f2iEL297DdUzf+4T5WNDw+ArYW2wR+YTjBaQYH/Ld
taR6nRk+/LrofsPODz6QMbXxWKcyu0cI/tmaGmbI4zzR8HHtCWc44bqQRUUsXQ+0
ezZKAMmFvtE1+dN6nrdT66IJDK6IS7IOCsUaKCS9ZPB/FmS1iXyI75NfIjXMQUoy
kvNTnEOi5lQo5TeWya1SNUd54BRS+QOdbC4uhOMQE5EOAnrK3a8pxKcXSebXkeZu
1jAkQx0wBoxAEJ60n/Sb/K9nI/3CSDYomyY8MpWbjK39Pkmb1QbmlOs6VYHEwiCO
o7RHKKWc9pQZDkLPOw0ROCzA5rRlARQzuN0W3lPTsR9nrBhmyKI/VFNMhHvawRVe
eeT1PK7lU2ATQncjPmXy5CNIhy0GJIL4VEeqcSTWObieXq3VEdiWLE1GOCRpdxiu
Kkk0I596SU3RhKnS00drGqmUGh3ppPACEqBCR4Ln3Y6244KviFNP6jKp1nY0UAWu
N0PoQpse+2y8gla4EQWmPL6iJ6K4BBx4ywveMShyuDALdtdD7ei9tHthy+m4vUk+
GbzJc8yDvNvEhjM3y+nvVdzVFdfFbYz2pBgSRYf6ORhZJhNTkrhC6pBUcPEA2Fee
Rfe0y6V/Qsj02hVFOd4MaKHWgudVjkL543WJCmXlTktUMBxD1fgxZ3mI0R7B5nkP
CoMxcz+aDWLR9AMe91b+Dqh1EBY4ARslbamXxy9eWkZABF4xTYYFpLs24Ax3JrdA
vJk9sj1yKwYtgQ+8SdorgcTyubK48pVEcUPighEWGj+a8uVotyTS/+DeCGGKzTHi
g1B7Va2xFw5hXaYpoIMA3yxsrb3+Rp3wbdY/uuRHHpLD7ZGvjNUmLFzsju3Lue2Z
ab/4gIXjc+YZd/d63APNLt/U+cu3hWh5bLcj9uK9KLJsZcUv0aUWxikdwm9GoR/H
hpTa7LkF5DdgKhW0hgju1c6dmLoFR+Cndw2z2IpKj7pqzvRPIBt5tvmgPDYRSJTs
HsPqP1Q344n1BcDaqDK8rtQRcKSAtZ4nk8GP00MMNQuWWbVeKCLIP118MQHILjpD
1oenSQTxx3T7P3tvgPRuuScpx60U9MdLm60lYYJWb+sR8Oiz9ukHnqV7uDNvBI0W
oFDWOJgpkZRCyfZSKPDLmAsQwQD0Ld2IhdXSGUbXFGGnqkiAIiFJfapS9RteBOWa
P4xg/Y8yyKU2mTAlPAVtx+mxJ9OatZuUuND3tgNZ5M0jQOZfrCwrCBzdfcZ8xg48
z0w4GkQrxIvFRc5Ni/ppkviSNbRcJlZ+WC9+3A8IVDx18b8rMGUUt2NOY4mZ+X63
KPtY/BSdkPSrcnIH8tL+fhaiHS38cR+bwmb67G6X/KrR3bxNIKTJbtAsGaaseJ8Q
dESFZfxQ4IkVhA9eH9n+dhzU7ax0BsXGdGaVWVjQAkXWN5vwVJfbU99qbPzgH/dU
8NJmOeCyBaAJxgHXnLgXNy4TLbdELRqy5XKh3nP693bMKbojZX01/6xevUgEn5F4
vqzGctXbb5QmN+ZhWt0W+15cVPQnx0RGc/F9CV5OhCNAaMen12UKw8jyU7Hkq2tZ
QU5TyXspPo3KThRu53hFDQVpuoSaRibBesmFYpIGDNtnucBiX84rNZE+sTSxmsOP
u2oSEbOOKn2YErNYVn6kM1XQc4GbI6Y3nVZBF5ikuAdFYwVS546v3xWwcZx/D+rg
5QJBKQpdpov0fo1lXUjToMAoYgRiqx0tOWWpBkg4rtNHYsB/TA86+Eu9BxMVlmFU
5qrje5yqwSgWZOjs8yc7E3j2ShSkU2DWgiDgF2OsE95fEkC/TqiUKhHtQRyetdJz
`protect END_PROTECTED
