`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FRtwnztBlDtxgiwAAltP/lOb0v7JpeAREe4tz57cLUyPrNQJuWk0K4fXkdJD6WEO
afEvcKztZOcVGQRz6xUb004ZyCLbczE7iDl9J7udTcII3Aj0R5JawyT0LLrjqh6K
x2bvIFlOhcp5uMpVZ2nhKe73UfHT49/Rv9CPFfH1q4TD0IyP4I0zwpsq2rumxg2Y
MqVKcRSF6WZcPwZyurHkFf0+hxG8MNfFzz/2k3yKaKEEzirxLgiXrecFGmFN2zlc
yDmSnj+fs9efZ72d1URK5OB3qj1pwxX1Mztw6+CetWJi7Ds7EMaoKM5dhV3AEOEC
sgT/ge37Efs+VexnOt+X6f7KAl7Qpc88NbzBmJhVWk2pfF6e0hCwGU3Wx5oGtR3r
YwHrIlpHLwQ9SQ8mD18rh3tmj4i85FOQJMGPYN36UXKti35A9PvWN/oN3YrZ01B0
yx5UO91OvtM3l1/IOqoMOTZkV7nkWS9mbXfLjXd89y10yjxk+1UlFcUjhN+8pana
KQeDeq5tyt53OGX/edD2zoLzdhABsaWnvDiFPVX+cc9IqVHkNBVkuOhj9LrFXEQD
weQNA8vh1uVX6NQo26/pftXLxP4isZrEolwSURUTp1mzAfQ6G0tOp6g2s7ve/HRz
nV1+tBhdSoivMCDL5Mq4w4cSenvq8h7Iz496Mgdjlk55ST6T5UeP7wtFuHuVwkSa
pT8RL/hnRs/5Ic+xkalEYkiiQRbZ6pVefsjtTbTT0NxyILLwdSOxpN+MdYymTy+D
6mIEMya2K3eg26joNQDoGbSiSFe9KnfK8ZZJyBjmkLRwWo+ZmnE+7FF5rHc+KZkd
YLe04cSsSKU5K2xL+fvBgCbxgbsMRmkHDGGIzvvynLpnIbRabksXQauBJ8ecVwwH
BDVkQALz2AE6+IWXv0Ut//aW1RcG/NN05tG36pbBHyONEafWwFfBPW1CdhX4SE24
CUpl//AGp255bMXEy0T+2x0gzZaoO5NvLFJepLp6+1rIDa4aPFX6CeA5C+ERT7D3
Run3JUj7HdRVibz5m/ABFJ0MkRAVUk09b7yVDouvQFpAb5T+Mtl+H9aKQ9ZbB4rO
G1wg7eOyqrhTh4MBlCXfhChRwBXUdDybobVFmTkTK1RzTJrkShMlLXG3BdeXzcIM
N9aoxZhBy9FARWLhXCQbuOzKL5R30Nz9hloPW5fUemBKUab00FDVcDnP6z+bezfQ
UR2NT40PvCBFj4McHV9D47/Hi8CVbfvE56rQDv5qIfU5EBS/VEKymmSSjCAzChCj
5cuA0QwCUgNxo5+B5anyzrGj4PvUqaCW8VKlYyN9BPrAR6kdryWJ2rlouAzwEhJy
`protect END_PROTECTED
