`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2IGkD7eU8B60IICvfg/Tnyo+qs88tRHRKN4YRNvtSo7twVuvKvxmw9w3c0f3oAOI
rsV+zt/CPwOSJNKHSQWpkg+YywIwhHpUFq4DzydUCwuMDFqdIbhknWTRvKMVaY7v
Ofp+l8bQc0fZHKo3dZb9W51oIYkorpC5jRpVhfI93PQkDqUFSvmBZLEvtZmderOs
LE2I99eCG4fryzIUIWfVQnbWRy4YlDtvJSOUliMSGDtEWlyWcd0ubc0bO0bF3tx5
Djo95P/A53ZIAmmQsjlTpYVJ0BGMKLKlQdBSKwCrh8qUJgftWyH5uiJMwiY7j7W9
LsFNx0NN4gkuwY/IGKWxvvys9YbTk9y1f7ozJi8/yzkhSMDV2RZiRkZ+akDTMft9
xd4UH41vK8OI2PxhLqH/k1VHgGLBwl5YBl1GyDULN8lhu0NNcsC01rLl2y5e0g8R
n4gGON3PXc+Ob667vJemcyjtIICdNiJf4ZQfOkPb4PUkcsE0bPOfJdc5pQZS32Ea
ZOqi2qtK9G7p9v1MZqzmkLIm8y/Gth9/7Xput0yvK5uwn3reU957JKOggpfxcDMJ
CU0jAJqH0TP694PdW6BEyhOKPclsyis6r9pHQFd1roD9kMa7dyOoetzTHttEt47h
20r0K539tglNGX121Nc/7SN7+PDN6gniDCjyMikVb3wDKQUSBy4GmROP7z55riAj
IHlsOCWSpBoW3NoL7opGjSal3R1OhgA852pungfXClvwbqeolWy1xWkIFljYns9u
hBz++VTZpKOIdxxzTFTYk1ykgWJHPxqOu//VbfVgu1jQ/ckGnyUA8fZrzvNZyI4h
NxGu/frOqL9dUN3xgMsKKhaGjWr6DjO7V7itAHJ5GFt7Ef4zidMOkvqnWNnBeFyV
S7ezOSOGqcEeGkgQ1zSPSIxWTAnRp8b/rsxV8tz8NZYYbFSTIs1ezHhLUlRuGj6k
GVbSl0PFIsYFIc/42yWB3mOozEwzAboaVpj7H6t5c76l6BvyKDchEivfw+1brVI2
`protect END_PROTECTED
