`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zmw3GDvDayr7HB7zRTAHFLL0n0BMcXdxaMrGg/jgLn9Y9Gif8SscaZvQY86G6Jyy
7aLJWUKCnh64yw8qGwvyMB8OmtFk3y2y1ER4ZkrsAF/cEgffoxBHMs056qMbUht7
LfALuA5Ui4oujhhAE2ArSJ1uQtmGgqaQ0zOpSlRCB1WhGamJ2udc4osAmyIPGlBs
YS7RlZh+zegYSkqNwuOTLhbMdy6x9yr+iPSsUFHTWXXGcpXEqDRo0XY8iBhrtnqd
Qx2sW9UKV5VJjQ7KKZ5uOJl2L7aHosl6qLDFa6Ip94I9sOzPOH7+n/6ImiJZL4Iz
Il3h/8pqrlho3xvCFtBJMrsZ2ocW8q/BmCtmsjqz6SKXv3DAKgc/ZTUbmQJDH7xC
PrZ1hBHul7etnUu9bOjV48lkKpeNHGsJ7c4pkVrj25dD/n25HKCm7UMlS3Hq9ju2
41VzaYU33+Cubvs60QNb5gI3Sp124qTVu/ZT0beksCxr0pNNqqaijZUAZHef2IXH
nT0QBrs+OaRtZO8cSdJIixGSzFv9oe9StBwDCTZ8Er+5M3MoHlOQJTQy3yZR57ep
KFqFpM+edLUHcCnrVGVBrz/EBv0TLiqYc8lLxZ5ipXQFDfygLJ/L3O2syaE3qcKO
UVmE8g44zxSnsVvcyO527oTJY3M3yLM185r/5QqpadfLCt6z7o47kdu8Uh+gs8AM
cIWSIxFCuuEtIjNNZ6jAmn0F1tz0RIPlrw/HgoaGQ2QAX28rER3++rBZt96mG6uy
`protect END_PROTECTED
