`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AqhtlNFYsxfAMr+pQxPvVE3C4mWEaciYzw169U3v94BlbZuhqzm/M0dr8HBwF7iQ
CXCLwDIuQ7PiOjnaId03pEswFHPeJjRQeVT672xPYVb167WVxPuDvkU7yMPYdUzA
zJBXoD/OACl7WEFDfWCUZQ1yEX1vBCv7MVdx1tiH8/Cqqj+11UrhkiJMlrl21HXx
yk64yKN/vJ8CarWCch8gXuTwnOH9LUzB4DD2vxXyCoLyAIKGygyWdtjGnAU8/mE6
GyraLh8WSubxNRDKATq8pRVFCR/2B54j6Q11zgnleOqcycDdL9u/va4qSTXajS1z
xkspcUk3QcHcoI2qtdUtsgBg//ur/NoH6FHq/evcZgUhyvb8PYw9pUcLZvjKeUvB
hTvYj6rTNwuRQL7Z7gK5H3x5MWL24j0aRP+tteJC1MZk5bdukXVEINhdao7CSFfU
O8oez573IKFzUQllG93oFcgFwGTeHq6SmlmXy6645NaCTmn5QWGFYyANI3aGW0Rl
2/scYMRYk65FSmNrIQFvSgOwQEaqMngPqEsargwPF3ELy8j+LjZJZbWL72m40rPw
z6lG8omGq3USZCJFBB7PZ8wT5/F9nltZfb24Tz3kAIyAEYYGRO86bu9CT4aOJiCb
ejP901DrPpZAWaSUxf7yHY86e9yyDXi16MW0I2yF+bt5Ag2sLZEtOBHlilbGOhpR
9NVw8A29asikG9dsjvcS1Lf4Vv2yeYbYBun9d1sBtPjd50RddTz+Z3RgfmS5zMNF
kfxPo2RmsAW+xYwprHnjczoPl9lc9sKKX3eKAB/pH3kd8V4Q7Kq0n1lcZFSRUlTL
xqIT1KXNv8MqCoQA1q8gGXIjCFyDXLzuM1syG+0LK/whGW/6EJO492AK+TOBXgr7
QSCybqWwZsL0XPOEOhzm4qhbclpL4YjLxhtg7RLoC8wyuOuv0MCh72hZ88gNYgq2
/5OF/mR5bB3DgijKHNcaRq2di/C/i+tx8AY36qkXEG1StegBKyyElEOkyVf0wspW
OiZ1XP3h7StSVVkjAvqgI0nicmEl7V5s7CLCwnOJnuS53BnzcOJe4Mxu1qke9gpD
PT7i9delWb8ciRsoe6JDlLMoQcQNG85pBAH5D9OAIuniueCeu3JPXfKEYmb+nJmX
54pn1ovV34UFgaqW0Z2UmQnr8GZvpgpNdOXBonQFL1XoECiC8977b0OfF9HgRxWT
O3kkvqMITf0dXWFqVyMOUqsSH1FI39e5iNCs4Zsxh16ngVsnOwCWRVd7m3pz6yMl
oWWCtCD+s4Cf8wuVY1mqdTkIsx3U6d6/04kTYlra+qkwS2MUkUCy+ADZmGloCFO1
JMU8fWmqesOYm/MdYuOyGtNprBazS3d0BtfeW0yt8DyVaPyggxNls4OEs0Yu41fI
M8oYUtlZY5/6kLV/gBRieGmtu/08F2THDsy8TNC4r6MgnSIhm2//QMpmdqLjQQlF
Pls5+0k8dNfxuz+rDiPz+f7mlTpHkgjs0ALNcvlg+JM7zdJSuNhYnHU8FVDLlkUc
rrhgz+UC6rxpb4rtT9b8q5TloayeM52hMR4Xa3RY5NENe8Z9GtBHOsr9vG4HRevd
lAcsTaKHp7ZqxELG94OoOFzeL3D4AsdSSFZqzT6eAwcB4iXAps5Ez1af8yn4jlea
vK68OHosKiP7kWu7Cxmi8fh+OFN5b6TRacxEI+pUSTjmbH5mPY/EHxh/Poe1LHuL
xdfyV2qzG6JejZsvdfYZBCf6XeFQcGmh0KBK3q3AAyT2xw3BdVWNBUhbEnpWDTuG
yrVVTVYlC98NNzOZ3pGpyhyvr3mrmjSOYVadNf+YHMFhewmLNriJr17k7+6PFpm+
fzKRq3c0dyS49EWVZwl7FHoCQCjQzHq9GibMRltR9v8Q74V95cOn6nxrYV8QsDLN
zqGKihFoFF1rBapCtJvYtw4iCFlRxuKGTxI5T8BP85wA4Jb+vqlv9gtc0SyhjESS
bKw/5uB1EW5aG1gk358c/pqmUYF/96dghDRg51l8ETxrGofuCZuk/F5fHV0o4vXr
2PLx2Em3OWDrnavDRzeRI89HxATBi28+iObGS6aGl24=
`protect END_PROTECTED
