`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d/nmFa6mLZvHcLfjd41RoasqT/uTKMo2FZhZzMvHpuCpyg5l6MMx12ST1K8Wj8Rp
2O2+LZn1+ffvyShf2sO+9hmhBLCQSfqgJeU5xzpZWVua7sXqqbLLugyWqG7j70Xu
8IT0t8s/f/B8GFmwslMHVgU+4nVQ23QVwH5fHUnKatFKDVgToy5/Ilhfaj2ZJDqy
ykFugrkByOduSOcLOa2BRN7PZOI7GKlX4ELMBoGk5FpIwVnR0XT4pQJzlc1iFFVF
rNS/FgK7nD5u5j8eN3tA0bl96H+Zq8TE5scSiIkOx8t21oHxl+allWEhshio87iS
uavSMofOGRIzTSSmIrzbIJlUeU3bj81edFZr6y6ZEi5aUGFQH3lwv45bDdlZkduG
C1+K2rsL+G44wriUGuV/imN2GIeJFOMk68ObtA/tz/QEmyo680AbIZr6lQl+FLaK
o00DBHXR3LaX5qyQ+HHpt22kDonEDcqQkHLarUj/Ml4FSt0KhUJgppEX6g/m/ExN
OwlzIqkz0dQ0afRpCn0iXaZoEk9mSsuuv51ORgUgz7I2dP8lXzEfPgpH9cw7UbRX
035/ltAcZuU3y0DviDyZDvBKscsNyvIXqsGgfj3XcxLOgKQFx+pcHG1gBYK5P02O
qtlCdopaYOzU2YMOuyje3sonHz+m7PpNrkkhZus2Qw6Z8g4y4Zj6ybBDTS2OUTir
df7DSyf2JF7jKZk6vSIu8nzz7ZcAvYn5kLiPJ01DlwKxFAactwtVv0P/2OYBavPE
6KlYEkGr0JFQkM30Q+GbdWISG+k9jqcZf9Lr6R6bBbBIYUbPJbWHCQegkF/eEgNy
truySF6jT6e2ksEeS1S6wO6QQMcjla40t0WRodka+tHG5sDHM0/oARXv6DrFnXxt
DcJe4Yl5UlEodrZDeWZadv9NXO/VtaTASSJQ2Bs5ejIVbgE6mTidd/8yfu/2Y0VI
G9I7PV6xtNaRiwsONmQxa6jXHaScvKtmT/1/IyYCjOU2JVk2oQiZEgMhjHjQfs7w
NtcwhWd1yIl7hgaM4aBTVwUBUXl8SstIOsdhup3foPVPMUzgGid15Qnm2GRi8LqW
w34NRvoohBoQF1i4quggxWGompL5GpqFh+dRqo+B9G6qZdlb4NQPfivygi4qIoNW
WpxcKnOD5vpJwgQJh2UrZ3WgpTTvG+IPjFDpMwTLMJRUrGtroI+eW2hvyunapkqp
/0mZxmgJSS56irSAHFFij0Y/D8uNfaCT4u1ufPEiqe3L9dz25r2a1Xy4hMIekiJu
PuMJQGuA/sRCrdB5J5QA95Ao4/Y8GQxh3KHvxn5L3ohtSSuyRw1ULRZgL3ePDVxU
vqwumtse9e94/erzjrpJHG9EmxHvMbIXEDJVjm+T9h3zInlmSxa2lKfYj+1BSpDd
aphTrwYKbCdhhmntWQYvOTsssU0YqkcGfkjOcA87wNrr7FSJej8tLo6k8UVnxQZQ
vj4P2KvXy2zffLhZDYE0V+Ozshq+NR4/Nzzf0Xluk5/6bxhgK2rMfROsyIuFrB+8
DnPAOLS/e3KH4OYbFoLr3H0qrWGMoBAx4EkRyYzuydMwsnID4vj+AJ74wtf+CJJk
cgvTSjmJcSrpd9EWeeiY6Dx+8m80BWkTszyeh2hFdzCJDo690EiEKCucnO7oSzAi
c1PGOIh7gKBU0SUOx11hK12oXpDGArWWgqSiH2nvDwAf1ycA2prBbrQdg36NbAAM
bGSThavuoU94HR2mSy4TDcbfQ2HU1HqXnFWyQuSqbj2ijmjrZMOmWTa+pnRiCoC1
B1b0RVeRxdzNbEYrKfARgf8Mr0jXdwMVgOIxSmQQsSOfkP/3n0fDIkrKq1cap/Rd
zkWzV0kUNgMuW8wgukvt/rLLMl48fj86/WPZcM1v83wF6VA6EbzgnVI0CfI5Nbpy
Bqmy+E6HzsA9riJVub/YlJjvnvpyr84qi4gHCGdYyIzQwJmlIidUicZTwh42hrYx
1tY14FotKeZIYgPXkqgH5YoFCqId/2/ww4lXeyVihPBJO83lxSnvOqGab3aDOXDW
FgxCl/DW5FVcLy3xhG1VoYHVA3V1/tSRSTnLlvqeVvAU5TCO6ZO1pY76VZf0ZeCK
D0vjfgXdAh6e8IFRR9PZG8mSMJkd+iV9JlYMm/ofx7QoKsLqgrMocv0SVKOMeKb2
HsuXaUC3Ddkuk85XNHLMlU4+3iHZxUWyfOjRV2cAytKDOWlYPvCahcs13Xea3qtU
RrXVgopqZQm0xsk/y9imnGXDQB1gQoaAW7qnW2eHaavWx8koESN+qoaes4z/najc
/KhJ3V8pg1WtLZSNKHuqESuz4+xY3J6FSvKFA+8rHU52KfwqGP5knm2+v2QgUjMp
HnC64Mw5CH4UPiJWXjVhQJYv+OzQ9lrQMpjfhTrwG1fMzSBfRSNVr03GMiTzBMO2
tqZwTfIrWwAmyI0cqc89Ip4sVXHR8J3bq65JS2dB1lnujhue6aYpANXDWHjCxcOd
tFKC9CoVnpr9Rt8VXtYpCyER/hQu/UbmIdbYVL5+CNTpXSY5F5tIev3w69G1VOM3
ZItlbWLdYakUa5Z0FYbJVzAgBy3mGE+MIiqvaeMDXWP8bQogoyqvqhZz7Afiqzqf
0VHb2onGEnzOoJzaEJ505HS966db7qRIJE3vYOw4TD3MUnNfMRSO1MJ0t33oPjD2
jr5UnFeo3dcVq8VK5k0xAwYMIn6PmSTmIREpvKefWIvxfaCjJe1ChjC3x7q0uRCV
0tqg7iast4PmHwYc18O2WkkUUFpiC7C0qXtMea4fk9z3yLhYjiAdMBz+T0wUdpGy
2S9UtPiONKsBWlogwZO6SJ2VlcDfT2rEvOU+hpnFvWCz5pzIs2qq4nkNG8aottbY
fH4EeClpjcIFSJFluWJcjRkcVvrAtW9HZwUSunQJtjOWSd89YhA0T6COFLMExXvb
Q1guPDWm0OHh/LTQBDbBHlQXUyxMQ+K0XS5mMQiG4MtAPVcURHiYMKPGmTDxv8Uz
fmoZCY2VbVGnInVSNlfqDpb5TSRt0fdfX/qbJWXMJwnhxueGbXZ4ydBpdG4skY3C
gnTCR24LWE9ThpgqWUlL5MHhWsq2OYXJK0wt+3GuvNkYoqLfeemdt7FG8EP0I4l1
ILX0ZkUgh9B2WFSTWpZODkR00QMuH4G1Z7M/LCrPY74Ab2UVgpcYBbRNKPNSrgNC
Fx0K9C7/+NdY4AHINAlNiUAe3paeypMPrS+s493RIWSCkKocWYbRW2xV+mCMHkaT
TBcXBns0q8ofQNvKYu2F6dbAT8PdayLeTu7IJmVaOkoU3qMYdaeSkGaNGj+rIohs
bLSnbDZ7W4zGEZiJo3c6BpDs8xJMlXeQBQkscHGuiO2UlkAmNy0IVqvSLlr8W9dB
vSU2zzMaa3JDRIyp4/Sp67M56t/OFMOLQI4JZnpYLRkiueF+2NZ9MxbPjuAH9jZy
Qp1EHGO0BEDh7ZLr82+6tTeHNryIJpFK4d0P0wPqOfrmk6NEtxjOHKgHWvMEkp8z
iIkX8dzZUbNHoJHXoKA1pW5eS+sbyIR3O3MdAd/Vte7z+DqlizalhOgSXCAuzchH
Q/gx1ckjiqoTmiJwatPMzPXC31q4wpn28EoINQdl7ipIQXBsMO8IJPkTh68YrQZu
WBwlAy1Btk3DRmY2s4OW1dxBb136SxSNalmyWV72NI7QxR6ctM+BNzq902ilQZYF
c+S2lwcYGkKiSEfUYX+ofHz6lTOf2ZebczbqDVXrCpPInOeGqj8+Yy/jMvuOJLkc
IvMejnIKWq14BRPfg2Zbr/P/9HuPgwTKVC1/lLfLqujZv13vduNadU+RRDt/U+z5
h9e1lgfxo4lRB8rX7IHk0PTcpenvO0irP95fe/Gzd/EOXsyiS32pajqLrsoZRolZ
kTt3dzQvAjztBZ0UmN5Sj4fpHRPGf/8oeOadimKEcqsqcxKLcv/Pra3N1k9RMm6o
Ij1vtC20FrUbY9Us7UM8YBwqBNz+BN8DLidgKLjr9lgwDhO9LXJaKvlmeD95nQt+
LjlO0z/t0ZWjfmOqWRvXKWo84A9jpPl+hiDF925EMC+WD9g7OEd3G07JVxevQbXs
5yT8qMBkiT24n72CdcvlT8kP6PZCypr+1YIoUHlbW1x6os0TJ4q8sRVQV0viozqh
nbuCsRpyC8trEK1DLmnv9hyKeywV8i1/IEcHixbSmf7QRDkqttofMWoXikSn4r1E
KxBmW91n0nKnCwhhSbfnet21xPeCpFIsf+gfd6/HmhY9j5B9sOIyKrqp0truIQl6
jFKn9Hre2IkyEGl2qMiFHYfoZLzr8M3ydoG15cbJZgENGnC+hQ0hEvrE/zd5ZOu7
Y8t2Ys7toX1t1zYrkZIUiG8ww+5yLUjbd4OtmEjvoUDycqFnTmSVRGPqY+Rb4hgs
H96v0+O1BxXd5W3mwS7Csb0YaB6gmcSkTGd/56pg2E5GlzAmWsDUo6xsUWYbGisu
GfArqN/PCO60SIth75pvtwXkkHKnxpj6aDjpposJ0X6hNYq4S/5XvB2Y5K5jGX6f
PQXRn6p9cKoNU58DmaY85qt5WA8Qn+1KcfKmPrPcO93ps7kxhBQ4gZTWdO5r7U01
mBiGvnvH3+Ujvbb7Kday7+Cn3+pwx5ubSvuwBYGHQkBRxO+uJayKaagl0R64vuAM
He+PBrfBfmpz1Slk8/XuLZs4bYhMFXUwGDMRB3ddsqtomHbsaxCVfw2sA72+5SgU
2O3uxdQiCENEQ/R1YPe8hQw/tn8ulfcwZ5Fza0PXlX2k0u891Lv26tL32631UIfz
DUN/DBRVB92yl6JmfS7Y2oYZ3aGdIWEymWlGmvTtRR01MX48M8rwrqO+siJ+fnlU
i9EaI23NhQlpniR234M68vXBZoFSvzGlwR1AuoPKl/5igSx2R4pm7erpHYygmn62
4lf0Tbs1FFKriPfkTsb+0LB53N0Zj589BvwXSiaqHAuwByfiYj4z4Kw5OJ3DsiTr
SGGGh4K3WgE0cfGKnlpLU6pnvjiMKTH9BwiGaMdAHFTcdFKCZdSnNTRwBFudr5Qn
z7mHUXUeO90W2VhsjaRddl3sBKtZVDAQM3k9ghIEsEYvim4ZKcroKd2yVogxu6wD
hyooGZ2BcAK9q+MYwC4KgZ0KPMQZKDSggHiddWsCfZJdsDj/8b2KrnDRr9Wm3Zzb
cR8HnvmZlj6wPAP28lDvbS8FI/WGs8NzdeNsYXaX8mgVlXn/bUzhiq3cBGNLSDdi
iiUMRTsF2UcSZI4nhHMpsPzCaZ1e/EV1cHfKKIUIQfOXilF0TWK5hO806jFyZcde
jXtqhh8YFZl6JHyijka6tEYPp4yzGxb3rR3s+1o7nTTG/3pb4xAiABv7V0aYUtj3
Ww3XO/ok0ek4WVnUjok+zN1bzzKCO/JTctsgwJdreXiUR/ksAkvNBaJD21LQvzUX
/AyDAk5OkhD9B1RPCoEEwJrjscUY8LzOAVvkLiC1n/gHubYxhzVDFq13h/Jd6WSr
T9FPMFzswq7hdV8meN2WIgkr04NXPquWH6br3ajgarInDqWDj8kGDBbISEVV8A8D
+7yeFzD05I7KzhMSFdp88CKNdbhodRzorfPbPPgUf/M+u/yNX3o+2Y46x1TC48YI
khGjLWU17WLcyLdt9aEZS2K+SvHZ6gceoo91VGbyg7vN76slKi5eGUqlrTiYbNiL
4vLpcho9ioDT98f6gsHqsBjqvMUVtAA4FbxqApubn206ot5KyKzSNx17Kpic3fkU
IX/h1RvRlZ+NslfEb/WlizYD/H9fNeGR1ea+Fumg4eOqlpXemUSV7d9Y1Avt4fD9
LFLBWnzsfNaXMdN/AFI0Z/im38pS0WEfU/CV0Gk7qKWAjIotXXa2/nnsOO6sIDBY
HjDAWUw3gDT/zZUpR3NWn8o4AsBHnIO6ItQIh9vqIrX6Ln8CoZ3zyILomGuFNOzW
37FBFTzVoPkpjRwVGdrSf/x9OYmkVuX7EZ9P/5927e+S05bxnfiP8dymCr8u9kjt
ycnrI7r950wkMczL60hoZ5LrI62HdKa6JgZ1KgDWW71GKpm/dG47gNsjWJAx8C1u
hbnycL9LpJSQCMmV37Rq6h3wkbj/pESZ5UtNmIeT3+bvtJQciYofXsy3vvhdJeQl
F6QNbRNEDgXW/SOtKY21e3p2OZGcz3bmF3zwEoclTCO3QMFrnkuxExNVFDPYl0HB
3M2sZUE3M5ZEQqZ+rrFaf45Oi2Z3D3cFfdNt2z6AicMdrykzHcfJEQLDUK7pNRuy
n/Pktg1B0aaXrgl5WLX+Y2XoaRYDqs/R+NYIx7qLv+XkFL3b0j9nQeQs0Qv3/VFw
2CjveQH/h2f+WcokpC4qf6PWwb6vcdIvfwb7FwJm9b7rSJBJCLDyzrjinXYTc7iP
aLAGDKoUXZtkx1w/w+byfySv/ggX452CoaDhV4T9I6ujwPRysc3ep1fNQMmXJ2Vn
qBtyZkqH22n95dhNVI+mgOzB6hHRQgy6ySeEfBIQ0NXko4HECYOdmU9Mll7sNrrx
iUDES9xvSctrGt8F1EEy54C6JvZRZHU5O38BY8Xc1N0ohE8cODU5wXPl17U8AVIh
FbJamX/keMunoS/wLigKA2+qu1Rgf5J3zJfiluBhhXr8Odk9dmvlymFhrE7XaYnK
x4rnoIXgSR5uXEsjPsvJew/nXz+orPTeL13GCBlLXdKPHdj6QK7f1TiaV6PPHm2F
KqvwanV6Qu94sMO5VE0j1s9Oz8rkSVxDKT2B8ryI82UIWstK4TP8jigiIYaLjeCY
kYRM68DJEFNAYQ9sJH8j78oxCHu15+1oIkuwj1kO4LXsjoixK9PloeaET9MfXGtc
za5DOAWIYARVcI5BN8g6KlXm15oYa2V2+K1zmw5LVfoxcgYeB+AJ4WZ3QhTR9Fak
7UAedriw0KWWrCDEbSAiyCYc114z3QDvUTvRoOhRyHRDMDG5nbrgBC+L7Yt9GHeN
QWdtoLDl4/GIqDXcSvb9j7oxZSzPnP4ccUjvyzT0P53ka4lo0mFaPA+enjOSIU22
GCHY2f9uu5wbCyNPrUwLjcRGmlb6bjsoz9SivNeXCJcmw3t/Uayjnp6A1MM/z7Pq
Ns9I83rrujVfeI2n9lOaeh9QZ9gNTzSBVvmu6qoVrYD41WF86yLJG0HjA5LZhhK7
n18zQ9xL83L/BSy4U7km9uQhVBEXyo1IkX8f/CGBWT1xBBT8Fu8JtntlGFDFqaN7
6hLZ61Hux1PIcWOmMm4egVYVIW5FXHTwTGEparFU54isE1EkT2chydcC2RC+dLrE
l2dbC01IvFc5yCQdMnEYrJgGNFK1eTfRDjfigFyFYCy8R+aCyV2mjFm+VNZ56lw4
nLZPKC9PXKBbk8Z6wMAL+xYePSD34CqGhUQAVgcvsETb8Fo9Mcm+TKJCNBCCr7UG
sA2xBMNANdc5x+yj7yfouclIB+2V/q1BlKXmeNaaTXg0BoRTZHRCoFYs7mS/MQnp
1q96b35roc06T8QbcphFZZSmCGzwpHTyFbWXVa39phGaMQbCLPDbyvGRESaajOcJ
ofsu4Fw2lS/kpGO6ZLEY0tJgCHrYqZGhwzOLvYmlWY+onAuSnvm5P3I9UmotpSmQ
XO3r95lcdhfZMDU4VwzbyONrcWvIYDxqD1fDtJdpHUpESxH/CA9B5lHcthP+cS1g
EB1XbU3X017QtVKJCsfc8FbHFO2sRJcB4hlyYxBKUTG98DIGU5i80iY+ElCelDqQ
ljwQNq/lXvuN8HQ7CCywiJZzYBneHxD9cxgfsYqAIchmd3eS/mmmokj47q1pqb6Y
Qo0c+vIgU4baGloZZyHC0cw8RamkJH2itFPxFkVBP1V+9bzQnana57VjAh134gLg
C/Kh4l7aXxJ/kbdUIkaxxTKVOTi6MiL4eZIMqgmtyxf+qx11JpykSxqjuSeS4Q+X
IxhpW64kWpERI4fTAAziCUjU8sl+c/LaJIe5J9Nt7K/xIbDIfa5oumsRAi8UWwUt
5jxr/o07S12p/uxNtrWKeEvFdhEQXsCAo92elo/gCDF20L0TtUCUwCqu3oc/8WYN
0B+Ele4SQOD+yIDG39Hy7eDuXys3kbG6ik/mQk0qIwNU7/uZhM5KNRMsQLVUM02G
3l+0CTz/C63aEtAanYlIkoW0C3wLgs2p1wpVIMn6kEr8i2dOJsVOOkvHvHzKH9Y/
tNMVGSXQJM+1t3YJZF3Ql633F4/GYmjO8skcPI4fR4/4tw+8969kSRhDFUWwKuvC
Rh7eYdCdzTY5z/gKS94uhxQowEthNlqnnaZwMAJywlrukihctKVGGB0dLwmRQqsW
meBt1DRqRruOlNAGpik/WkXfUWoUMP1fN3+JZtO5c7RJWznX6GzvhzE7Hg77Wym7
RT+ZDNw020shM6W9VsM1dSl5A6URyWYFNyrSosDGlE0VmySpz+ZXsA5GlAXfI3rM
FFPQi65rMVvd3JiX5DFB0r2FXTF2xgnhZ37rkYkscz2EZXFFDdI3wMFJN4IjqxpS
q0PHmkOwKNGad0GByRJ370pJGo0hB8uQuigxxGCsbeZadQqcpZ9gL6U0nR6HB+Yc
AMRXS8xwbopLJjVK/C1mkR9f5p5EPNxM2UaxXfMrOS+kVk3+REdA1puWcKiTFlNX
TbKIbVGKkxFmJczmFRDsBSNG0LfpoT1CdKCB5Jqqc5q3OREgPWh7gankwqCwSmY+
H4rVgrbb+ogHwMWUzxxcVjjVyCqkICKuY8h4TRUgC6raq+GW52FFlURstvDLVCVc
85zRGO7fmc8+tJwACIxcTXS11l7fcr+p6tLgto65Qkgxibcb6ubFsU4DhqHZsgkP
piDq8s3WgfTnm8H4QLhJVtn6dMepiECzseO97x/lhM3VdLQBGftEtEFYj8WJSIFp
RjwkuhtqHORp0ZJg+IHVa/LLWHKWaR/Y2mj/bQqchqU4gte3xIpBx9I/MSv6P//9
Ul9ndVf9/CEM1t3WJ5cT58PNhhfJUVNopu8UhuVApHUFcJQguMHfwjgrb4vpg8aX
lt9z2Dz4NH6oJfNqxxoGtBE1/kPrBuBX+s2e09L+7/QyNeeYK/1LIH6WI1RbvWQg
+Ch3NzCVIYE5JF9BxVIIVeltrdbzK6P4dPJn2++1zGGFgz1pDUR/rljq5VW44jU4
SPiDs6hdBzjUukPMtz6G3HwqySHBzproWJXOq455yYgOsSDHo1FcdWaLYeRz9cD9
vjU9okrW05Dqm6gZ3RVSi2sGXUnLlYfZoi0fUv/eov9WhjjgPJdQPG8CGHdJ3oaE
yL/QiRCQ0zXSra8G4/hweCX9Vt8f7iMIZylRjpPRceH/YRaDVTYNTIQNaFDm8OoJ
d4l3yd+WHYY0I6U76N5oyEsnp6n5NcJXcIvKPuW6DautPinZXkl6w/HWaoZuV9vR
lvDKu+cCCISjg+86uDQuFoxw7+cBfc/Tm7QYtM370nzsfmg+0PzQmWvphTjI66LO
KY29qD9dThWRygXxxzF90wnMa8ZHB7YVP9Ps9y0WQLrA517tE3QG6Pp5YAi63E34
U3KgcQjE7KxzUneRHDp2OFYDFkViuhdC88kvh44kloB0Ls3E9s0JdFUG3PhZaD+d
OQglW6NqgK9FSiP8nq7081xR2KGvRlVDb/8PjmT8769bUmNqc9exhriLiE6f6TCM
ogkqFgqCyUIbz4Wl4a8B5meBeoEdA+MlRDSxKddmOBvDkAzP0CD/GBdt1EkVxuDB
sV6+VPfkQliQoZdswghfZyKhcu5vK2Z+t/olgGmKxtFMr0PZPczRAKL7X1FS2Xcj
4VITfc354Pz4CWr4qoPLhf2rRJ9WCw5kJ/zjJV4eWh6f0YkCTP9HNycygwKepoTZ
+vmmb8Y0RNT0vKhRcIblnw8SUrZEmXPkzfnpbfjYIN1te4zyYFJ2SpMynTm4OT56
6+8ndFlCJcQh579qysNi7lpAEbPYWciXWyLbUu/0RiqbOIgYXmxVgvAmXLlwvzFu
X+x59471kiJ76Gj6hjIkvr4Y8Wr9gTMI3na7iA6/aGVMnd4q0tFr/42VJ9WeVDZW
E/I9xWiw6ty44jM7G6c0oWKQ0jMSc7e4HcPuM6z01knoqwO7aGaATc57oxprJ6aF
7zWdkKKY6tIymw2rfSLcuj62JBaimocLBQ6CU5TBI2kMQCi+ypdOK8BJkkuiyDPG
Pu+Rn7jvZ+SvABUy2io0//AhzxNeKJkHt2BKbB5n68RexwgHp5yZhPZGd6J5ifLo
XkTlV0bjuxkdNZvCn0OqyCafPYmf8UhaQhn6mQb6eXeNODgbnb3oOzwOKowB0vFI
gIeO+ic+p8aLhBQLHL0czKqKFp6DaChz+/sxMVkQQzpjPmdpdzqeWD5yDmrfKIFP
OFaKn45UqLTkelnZPYxWpPqvIoYaIiCpBMrAeYUfuYty7yYOOWNOgvDxzNifiRSi
/xBgmioBHpHyajxhZAK9E+ARdIRWXlKHaRrh6jPO+d0gf1xKaFuwPctd1hwvMQlt
YEDCeUk1ytOkvk63c3LHU8F9b7we+uvs36MKrzyvgb7zDLHRdDOs7YuKPrjb2/0S
s6aCi/swJpd3PIUPO0tE5NW4UWclIkbWskv5jQ4dC7HZA65M7f4xZlCq0o+Lpec0
NixaO+OPPEVwsf41kNJcb78MKo6DDJM4BFonDajDKJPxeMERWK4D5IkZxPqKnL5Y
4jY2jhf6j13gLBXH0nC3MPKBR3HdvmD+gNAuW+/AYLvsDdapz7CTbovZhGj7Sf/f
x7edx9RS4pcnZ3hA9RkRFWd8t2a/DaYvSMvIm2vc7GAvps8S7cSw0b96z3Sso5j3
WGH13EWwQoAeBd+UywvHVFmzMQcgwqG7hc6vmBnr6KYs37gqb51BSDzE5flT7IYR
uI0rmoi+tFSmrjL6UEsjxR2S3FmapTjktzb40EUsyPC3qC8t01Q7ffuO598YlCDj
dWoRcHZRiC1EVLrZ3IlEjJqxpxutd7F25jRNs8SPho9/YjXTKLoZTLpByZMUAHYP
CjMh3F1pNAxT1RBLDdlHyciogKMOtFItMxmwQbfJosrHrZRcleNaBqOJm31kDWLH
1CmMHV015rz59N6VsY0IagewyX5u/RGCq69UdVcCQyTmTWsktw/yNmA2RSDRgd4g
xyLz6uYcr81qsxE3Dgea/9Akewe4ibRkAIY012qTFbzjcFEqayhJSqtStqoyIu8J
hfQCX/zjeu0wql7CXcsmtxgL0cKa9+GwEIafF3/0h4B6Uq/0LqoJRzl7/YaRq4vb
NQuRr2tsqlKI6Rre/vdvAj0mJIHrBj4nfxD7E+WAbnFB0Pd1zF/eRAyJPEhAFjwq
JGgyC6aXHLaTvpKozzTZzAMT2PAFDV1U9SRMLZFxDsGL1QzVZMDFWC+dXnoecno6
CNvm+g8DlDQOzCNqzb4bUgyl0I5XZsVXbhbtG4pkv6BqZj8xPpv56SVMPGqrO+C1
dfTtO9vkT+WSSLdOXrBbwHH6mCSjzqa4Iq0Sc+9ZN259Kh5vH3QRj95fTHjQ4muA
DXx45MT6bQenPoC4WKyyLNTw9MidcBbuAqhBDyaWv7yp41fspH1WSPoCh/3qZ68T
D6DIFBDoT7QYEiEqSs9gBocrMp2lAf2E9jnBiZJjGMk6FuZ6+LHNJt//WZvEx+1T
idMkAQoIcQ+J5/UZiQgVHfp3sr7gvl70Mi6aJd6yxPu4ulBZpLMbF81wzCxWiwFG
0BDy/25sSl/RIl9Hm02jWVD6d4or9hB4GyLYS8qQtD8T9calSmPQMkXccO59AX4b
cwCmQ0V4pVlMSH74IeCwm6aCLu9+avj/fzOZ8zF7FK+UzBGYDVomjjutImdvDZ/k
Z9grV5HGJEsrIAJfWLesb89gfKSiyfTiGoO5b8Rue9dXxLTTn7cPbH5CDxWDwKa9
ndTfAMfaQX3bw3lQrzKfLgeFZMCTqV1osRzONJLUuB9hbVYNPBbFjE2NOxlifWI9
dTr0v5/v6xjF06w/RxntqPnqKUgjHe3+XI7SlKG0WEP6QaKDwlFyOh7W3fIg/Dg7
/Ru9TRXWz7y+XH/xhzyIbWTUUB5auddV+m5tjpAklByhJU5WLZdSgNaDQz2LH9jq
axNRrmPwLX2DHXtfabOACWpuFC0gGcLQBuHP8EyiAKPlPggfy2MtLnMAXpM+e9pi
i1yGh0NENIqBry8ddx7vjCjcoAspwzGujAPQxpZYcPZ4i1U1xqURYPyVozCavEJW
nobo/V00iI4gLjRa3lTeAI9go++YENKqdWB9DKUgzfXvokPhWS18Gzfefu1uEJKC
NOe4khQSIUWS2MhSzgMnsV0iVyaiMfgYFn+lqYGaQbuhRjDIyjlwU7EWg25xNBzx
O3zK15P/TzJGwzrWQqg8myQ0RwR/e3++0sR1Ms2DD7BnZx8U8SOcKV+0onboCvMu
pai/4H8Uii60c48QV3tgpRz1Ix6I2O6AIMUHzTd1mG666jA/x6sXtOq6XEcu2R9A
TOn6rWg1y+2Nur9brdu22RhvyiunwfPiPsRENOcVh8LRWhckz6UFYNshMLa/L6lJ
ouykcCaOpY3zVMrHcO2fOKPlO1BCid6eZm2z4geVsd5ymLj0IQS/yNz5jylarsTK
8cPd4eXLHaGT5vxbYbqaioYSV6SeYJDlawNJ5QiD1OOZ5ErQsEE58VNLGpCsKc2e
LpqzYucDfuBNpnC6wL+5q0W8FdEIrjyt1seyrNCn6091gpmop+Ow1H+J3KX91Cd/
/QUFl0n1aiRq/Sp1/E7F25Us+aOmE6yff2KjfhmG/5+ATWcddKoqP1k+7lX3Nf16
elaSlJ+bKLSt7M945F9wlEgr8IqlW+d+awu7nyrpmV8O9LxgzhJ01DRZKvizIE3U
9MxXnQxqIQr52kA1GYAtmraaQtMSoKOokpNlsqjq8Z2/iYMEhx3nD10ZBg2k9HU9
Jcv4RBJNvCmr6YLeGk5VOuz07nXODYU6p6sGCi/FMIkCcjSY0I09o3SZ+WTefqUm
03mt4jqh5ERpzArs/jjpRm9RHynoV7685BTHEvTI+6Wst5LiSa+xCKPyTHYNFseq
YJzNQ36XG7B2t/cOf0ddI4h5m503MzfH065DShwHnz3l24g8WRfMaERC2K1ADwtE
dkFof1jT4gj1R+PFv5vQaqJHp2dP7scHl6QjWCSskwm126d5xjhclqMbDf8t8YCO
lPiNc68ww4Gqq3WjixhOeWUGqxYNguI6BB9S+ZPqZb8ZFFmlVJxYkM2LFSzSrM8A
mxxI34VSqUpO2Z32vnL/64IKrRciMHv/lQDH9FnhjG3kGDUuRI/W5HvMPaTPbdRD
Bk5s9wSVsntq6wcqV65Uh2j2z8u2XUvVrlCY0EIGt/uBrVLzcNAecAJzIsj1trn4
lZYjyIuCbSHtQ3X5piRAVv5qFaxwsEo7w05Qn8CLl5IU86WxWgNnIltr5jDHMEVI
c0Fhl2udlHtYNdu2gqO70RTyZfQquuWTduGEhfCdJW3rLlhZ1pWlXaylgVYRixie
KtGfEGtJJeZ8eXcqsclq4M6mOFRm6kCIOkofqn20eDWarJsLqkqVvvyuCBCcTqOP
I/RnpMmGR0jWZZJ4uddXZCFbjjUYpDWNWHVILd0YtS66p7GVtiX8TzIKtdgfzu48
vbkko+BKBTogAg7xp+x1APCR18iKdOulfLgGjmZd6vB+JeiIxbYFU6cjgeTwAWCB
kDuNXEWZMqZBwi04eJUsEAY3Vstvw0xDokhGTYUeMT4Ro97qlyh8m4qdiydFWEY5
ShV1Ri8xOdJ3fcE48sG5O9qLWPhwwh0APZGE9GDUxbJBt3rlPBrUZ9L2awPdBAUI
tj3lV73YEgh5wvPwaejr8UmmWUbQrid+GJC+s9hdVQ0TwAXDkNx/SbGYE31pdueS
zscfpsVZv6T0ZXwPyXEEqKpEFfGgVO/lGN1hRbj5uDDp0lC8U6xvD+8ue3okOcU2
ASbO0jI2BVFJ2ptviGUnIyquUyh5DXdnwLA6hjpQtCPbzy5rF0AhSiGtRN3Rw7md
J9Sz7vDWp4P84BclHf25wXLlBTaSrrobXLEETroggLhyTOhe/8nS141Hpmna6c6t
Z5sIYqyJ6oTnxkjAPWFA0TKvBKsvpXmawqhfMvw3YXVo3J7pKZe+HMHP1QI3XWLf
/uQ/lzwUvfFUqTBaTMA1U0AZYujNxCpkm6xpBtD3uYEKXlvnk8M2rPIEvgO0dY/U
PBeH0unAmK1w7P/ASpeVGL+Gnphlfp/X3GJJc3y/jdWXzYnQSzSRrKCwdHMKEG3y
eLk60ngflQx19+kcXHyYywr4um7YC0N8yf09EH8dFuPl9Y+Fq2fGQRSGRSTI8NxF
VXx+P3oIKVctgThrJuQzZPp5Drbsd2Hzik7FgaW0zqTxeZ5gAVtVIt5YpImbEkoD
mfm7QCGU1Xm+Ng7bzR68tC3n5XRAKP8ZUXMGKa2DIc34J10+tVy8b5BBhmwG1AD9
Yyz84ae4z+lynsBatS1Y4iznwvxkIuskFrEa9REJVUiA5/HD+jaq+U/WY3VUXC7Z
PAV4VHsawtUJNVknf20Zzv1OYTiAFsYrE557A3PD50CUwrdzIWNIK9+Ihp8FVuKQ
Fq22yJODQBuN+3/yZEV3jm3X4bbsg+AugoLgh0yA7KflBKZM4RRhVxxaEGRw6TsP
axx1rNbA36lPloaDvIO+T9o0DUI2syDUevZt+BtKsCYQ/JNRjVyaW3Zyk4CExjSL
xPkHFDoEIX3O6sZgZdmJl01ZMVDJf5Ey1tYIIGtWdPX0pMmEmYKBJYLX9ik3Y0Q6
/stoR/n2auEBWoTuiuisGhGfF9M6GO2KL0Z+mv1On9t37SeZ1NFda7m58r/P2sLu
5CHoAYW+zPbVBs0QnAmp4eVq7VqdlF4ixFdDq6YLS7XuchapduOmjyDV0eac6tXG
nLssmXXmSCFaK39RVCYcU9ExTiaW2+NzRvKVZXcbe32y/AYv8lmOmp7I8tePt4id
fnVccqG60XUvinqWfz2aXwL5OFg0rjr2srku+8UpkUCvbm9EF+qPxrFo3O1faZ92
fVzNFo79nbfF77BmGlrGOmohopvaFf7E67XvcWoxXHZT0XBeRLzrvG3BBX2L90SO
ggkFqdmxpVtWT5HIdf/MHAfuFAjhMhQ3716UjZ9OyFyt6l9XKXlmsyaz42ZYf91g
sA45ogva8b7fwo3clLh0pEP1YHAInkBRBQa8qS7dh7ROXDT+bHlpjf53AkozoH1T
4r5KHSjXIaCCSLe6greYI7477m5yruWpZ8wMMLVMXC0HxkZAup8bIuhSOGlNqz5h
vPpHWlLrbpVsqWdMndSt2T5PTnd7grbHw4feFH+Xzeb/lpSj/X7aiv6L9GT2ndYE
42oP4Qa2oy/5QRM6YWXMPHtsyRQb/72jqgZhRsP2ThoxxkdD9s1pfwGZW42Qj/IO
Qfq2uHW7ZSD1bCSe/CbWlurV66HL2EC2wKj5KlLRfwJU8RcIBuxzL9IryEL329+f
ogo/AYHgoErCk9qg4xAxSeiBT+bHvm7h9gWOyMFH3L6UzJHRB2BipuXyYoNxYepx
Im0cNZl4LS5HaSXc1NIkWmoUEufL5On3Q0rQvtWf7xVJNZYLBo0qHMZMvqgq2qiv
g2OZTheJwJwhxdnGJbtO2PjxPM1MKCEAdOmgJnwcd2eeG8E3Gf5uqPcruXJTOHwY
G3v4qSEqtaBjhIsD/qWIcqLB7iOwnFw3DwxFHubg1qSrYPm01MO+oNF6Ps63Or3V
d6SwRGeP6ibdkKHnLDs1E/6KgK/6zoWSFzu6syMyWRS9XyUKxDoXk5c0xT1z+zq5
uRNnltT28UbnFmgCPerTrdCy4ajQgMz4k5k49xdgI8B+1ChcJpSP+kiTeBpvQ5L8
a4lyUrEg9LYPXX3d1f1poPICKSC5/H1P9zsSgt16cGA0IJEPfRWwxG7q7fT752cN
7VsZgKltu7GzePx+GLguTpeuiSxDFmV7a2VFViPNfGGfxbaJ3p/O7rPLxX6DhGMc
VgfSl/DyjUCMnviEhM1OTezklLDsYKa4I9L/xn9MHvigZrk36BL0G7KTlA4L33XO
Xt6Etz8lkz26GUWOBZO6IvpAMkDciASNmOwe9dgEAW4nmtZ0P+7oOqu30mRd/cVF
0BuMDAiHKJ+7DN96WHTIm+W1+kxBnsmMc4Uwgn7oQwzaXIhpSvH2KktQhkI00mCF
6gHBTa4/VXkKkw0WUKJ++jS+6D+CmKHC0xq4rBEOxIQgM1kb7TTnPx2rT8Bh1PnD
NAZuXhFFoFV2kQTF3tXEJW4shL77wSsmao/49dzo233la3HuWkK7kK1z6f0UUieC
EOWE3K07M1Vu+HEYiQ63jThkJioXFO4SGA5go6UHVcGandMsG0zyJFueJd31SPg8
56PGLLwJTNh7QQ8Dg1Tj21e0wbulF5OVit2w6av3CR2Irg2+pNPA1u9FS+Tm5K9e
9sAVu/B7ANrcinChHQUg5nLakzAWsEmPz6FyoijHUDCLrgY7BijwVgkSqOmPaIPb
eCHNUJOrXjONxOFxvLlI1H4ABc+kipVOLDMYbQKtkMrITiSaAW3yCLiQ/lKh7aup
D32P925OBmjy7YxxrAZfmacEfc/Cb4QVG0AXn73mRaGISmK+Y4LzDFW3IB2UaUeX
1ALaVLD5MSfefeOJNzfeWidlOSfVXQrPwTnzayHobgTblCVtJdqa4t4wgjUCHL3U
xUlJvztxHy6phQD9jymcfcNTJC2whigQUg8S2P2/ujitaibzRD/BHxdwkC13dlTt
tFpxNDzbMcBGrXlDH0KyrkRR2TgutqpwmnvcwvjrCtMKK3O691t4R0KKstybuWku
0AdXhz/rARCsepYpJY+MIkWjpecU3pzCoYyy4eems4V7kI5vRqlvG6x9yRbwoM8Z
8ZoPKecnjwhzgT2TnosU6+7UAsQPsriBMG9knZb8rqUlhGB2QOrvev40ypL6BLas
NgXKlkjucyBgNCufLNYhuxNMgSMTgcxiK/hku6W9v6i6K3E6K6qYCm3GJBO4clqg
NJ9aeGX9FHH8ub/tLJuN8zMsmPsQmWX6lcRHHyB+SxYXTSFhRRF483YhEAF1kG8O
xqowY42qc1jAI8mHxu1kJxluXHOeyfH8Dh9aY8yYEiLtwlHCIdeyWBos/VTsANfA
fypudy+NPKCCQSJABg+BJdJv4A+D7TNFcCE5L5m9LQwVNM9km+H5Z65gC6YW7EKh
Yh/QnTuCWhayHvqSHS5Z5ADINTDQschSgeFOH1Z24MWDLFUuFqtlDXBrubzkEQZ0
oyv7TDjduLqx4ejz8w+r1fwVUTWOxkQmm8HFW1he3FJSYSNSMA+gVus1fWLrth0T
ELQJo0XQbRAbaISZey1oxR+pllgACOraspri0kQn5ZzDYXGAZ7QqsQ1U0UPUm9Gs
gz7+o35GeBHRHUJJMKnyGvEmhiOQ//Cm08RuVrrokYPOAMXjjSCJBZ8JwcC+FydG
3YrexTJk4FCwiWMrpsNzoNtHHseC0L2SheA471+BFXcC5rQMlqFNLa2fGKgzdGcI
NR3l9Jb148G1zYAwHJ3jM2GAEGhrQtPY10xd3UvYL3p/ayDMznA+knTALgudd2bN
OdwIne7xp4O8wfZKrPx8P2X0HaKaNR+7/EKgNzhnUX77czuCJvNnH1/jevFV6CKP
bBzTFY+o884e3xrsI7UF4OByLwE24iYcQBqkIF5vKH9LdfPS/SbGMJ1tSpPsn8OW
usoB7a7JfFwGqZ7rI96tTagVe0HLqVgwcybouJlzmUK3QcZFoz1+c0d8RSzVuvpf
MTqiFqpa486nQ6Rzqx4tQekXkWtA4bOKlkrHzo2L10jfX3r7l/VcKejSOW5Es1Xc
xgP8BTk/oLoQYTVYVfWaxkDZ7WYbvkKDy+GRierGpgTcbycbVPjbG/ovsn0HWLpM
VQK0SfD6BCiBYSXxQ+QI8cMIjX2requs9z96TqrS7+pjdQCD0wn696bebPBE57Gf
CztqUOl+LdajItmtBf/r/SAi3ckUN1g+S4eB7zinEG9DatxzLZOInJC2n38xTC8P
+8nU1IofhRL7etjXxKmNQyVvsbcBHK+hx39jh75JkZIL9J3m7ytXrocN3K2S8JZc
unYZ29+M2/CZF6nLYxCPG32Pdcn2U0Cu6fzTUb56PHx8fvf6WYKYOXZu2HsmKz0L
Ehud07560MzpmEK59PYH/SfnAZjSq0+1naXKiSL0vJDhPzBa9wkuDJgmfk8hGiYi
t1reDw/ABe9W4gT5mvyH8RvypPC2fR6kME9DOWEyc10xc6xpAfaw9qOj57RzwHWx
Ocsl3X/RMu6/xlPpS3bMvTA7+/RiZ6TxBjb7RmflDqf0ArggUwOehU2D6FVN+JSM
DA/fBXIl6MW75faHr9Zf0nXVL+eDr2D02cw5s4wePASRyjBZgq387yeE/hDlUgqH
e0VXj+5GtFqQm8T3hNgnsGeZZdH+Ex0SqCaFwqNn0hqqW1+l8l9rQtPCBj7rviWY
s1OFas2+htH8lKGXYcyvSj1rXrulID4Qudm6NO8A5opBdSbhxubxHUY1B8I6/fCH
jboxiDxIxHd1U3aiR3Gzj7umri4Pj8jWbMFnshX3kbCdq460e/p3P7PFsTODJiq4
wdpUMgBGPCGkuDTh7+dAuz9SQrED4IElqePDHmUYxLiCovBbmv/biUidSMDasOSt
NXbaY9nOHcgZ3zvBZTvk85ks4NjV8eh4GMX3klMJ9Sg1Ya1W4Gl+shXLVUyaEbvr
US7H9hSWpmpeMFQlXnloH4yf+ugDsi1cGY000K/5d8od3a41gmeLiYkhJY+W46A0
v9HH7WffKsqr0iU5bGd0lEqWp0vIFEpIpULpTen5PK8O8Tb/1VCtaCK7SYuFsHnK
gnRKuRN4oc+P9Xt8Q39rBt5J0M1AghH2Lzq/65OCab2Q/7+0eg8r/vwilz1SimsR
eAxav0/ffn8BbYyto/pzNlv2AWkVlqtKEK7nmxdw6ZO4gejII6GZgJC1oyWLvCyd
MGksEz+X7YtTJ90mO0MXmQKfQlz1sMUNsRh6BoTubsLEuX66t+1YOSj7vxjRspDt
HdWRvcXoJnK1iL2PqaL8SdIxI3QcrbZLCG8+jA6iu77u5Qo4YCL7q3An/2z2C9dJ
yJPg2DBjwW/Wv9PQQkHB1EslVJ2FNY6vLfv9VnaPPGUrfQdtIzVbphK90AHpamEC
uABxhUFZH92rMuTOmA2hoO9cotseIOCQzDz9rXkQdp9HAFEeqCsLQ1xsMKk7uMeI
lqcElVqqtz3sn5LxUbpfJOQg+8Hjmx7+YAInf35HKIJ8pHMbapZwyulK8yYvVJG5
/5K3JqNaJCAzaa8hRZvkQhYT23sNX0mCAFljiwEJKuKFP7+it4b0TGMQDamlgntD
BnPzZov5rSsBr9FYQniT/9i4Y3gX5hv+mlaQ4dk+9Z7pxBLb1A52KMIATZte2X5R
AvlGryduh8G59hqGrmW7ViP8arnwgrJXqOh2r1FT2oZ/lVL2J7qqwURVR4LQWuxb
kaTUgR5JXM4pPBHXYUACi2k0CRzqK7E7O6Rtq7tf8O52BP/wzUvOo9FboWYlIckN
IoCvFbPI8xO8a04tyPDYe68rXTY8cRwLRYIaxHtnnGoAq6alasfUCnpIidGkoPqm
aua7VOfjwg/1gzAj300wLaGTxbnZoIhdBDgLOQaj1TpNKA4NAul8l9DDXgWN9frm
JWqfSPil4frcxfc0SqnXy4KqVE4RnPRYP7HPOVHDeWTv1OOXaEbnV4ny6pKFKPc5
OcT1ZqyIEc+rc7AI+DRzinXgqSZ4piCyZFX0TEDuqL5DtbBshH5yo3hkRHLyFap4
ym0AU0lJxCFUv01ROshtrwnCAzvdIiEE48oc7Qhe15euund63XkiKQYmDwU9EqeR
X1uvHaCjrZ8WpJya4sI4Aefc6Ygtaf3zjF+N2s0kCOrxYZmG97WnWpbIizWCAAoC
Ichq7fyoLQbBrAf6DcHO4Gu9kITWRruIQtOAER1UHHux95V9FtVkV73h3zMBD5eL
lxKpPdA0uZO8GYn3S9424VTSnqRGsnIQnJHrC/8JTPuB30KlB5cY8llWZrRjga1j
OvfcWS9RYYGhpNRFvmZa64OYYUdXF3HomntlmZvvGMiwdcMh62opiLkIeKZZRuY2
2qhqMmpDu3KmSjB2YxdoMjfh60I5NATdh704xM9xVwhRQ99ftRDYCt3kNtf+N61+
YW622nucFp9Ug35miu253I4c6nfN0MOm58+M3/bQ2aEZrcX7dOhgR33IQUTyp96O
2JbaNr8NfG/VtHWRoHGhyRFAGPIHZxPVjrJ0C8yLXnOn0W7Yo5sYTAW3MzvS5htS
e3mG2QyWhdl9A9xtXmul1FCtqOqWDRkfaf9Zu24yVyf2QWaOoLVU/nu2aH68xZgG
LmJAU54VuarmHVHluO9L9g2tMJcZpht8UkkAoBMfMSPZR+Np6JExZ7CBPJpurcAi
S2hEaUof39aeyIhXYfXEjHXaBRFaAcvTCcbT8A9zQgN1CS99NZpJKIBov4YX8dmZ
7DGnc3aA0aRl/Xcitd4+rbGVGoeFHyhQ54PH/UPCPDZ6k5qDsuSdidPi6xpC1ezQ
gtqvjJJqmOfdyLRI2y6ztuf7Xzh9bTXL+DvPnHGdvAyLLWg3JMbUFDR4/wbOVmCe
Vm7vtVYA7/k7VtLq8Z0+a8hP3++G/wYbpT1r6W70zh61zMBMeqZcbyXJtrM5oWPN
h/Pls4eJW9GG9QBd1XKM7oBQ98zfNORvW3+hwFhj73BrTRwP0vPWOi1i1LwMDPEv
UVaosXwLBNvtWvnctB/vKIDDRJDxiiubASexR3wBPe7Z/PC3Ovdf22d7Qs/U0mPV
U/mceAirJgl+AOZ7SG6pVF9YQbdb5czUn6zLtJJLtBWmC48QfEyKpkgPKaQ33C1C
li8dMwSvv4HYL5ZVY6TJWwN3MrtaAw6ht2t93aQJrkw4mpJaFkzxV8oOfJWj923S
6InGtzGwy6UTU3NTjdwz+w1Juq8jeeM75EFz+mf52nMylNDZKuCKMUOOSefhtp+O
ysJ/B5dbbamvQr1iihcpiEw/OB6XfuYwJuYo21KyC3fXKw3x6CKZHeuzTyVEWwEr
4Q+vxS0wtXHyRatp28C8FzVBurwBEo+Vt7YLE6VW6uezs3b8FDuKyKQxWteAyLRi
IzP1NUG+kV766hb/nHe2RRqV6/RqRdcejww0Yl1CZIxKerh5W41cIXrW+Mdcd2p7
mmQVBBjdpeRPud7cHVMNwdrWkzuX8FBKb6Sbp70wRlrNdYOJIw6DJeNtrdDRGh1Y
UV+FXlt/VqKBBEQfT1qI/GzZCbEN0bDG2rHcJUr0yJWsqC5QUUJf7iyJiMAMDkpW
WBNmrv67sj0jhBjCgPZLx/jllA/M0NpJ7fdj3lXStsUrnROCRof2IF4LY7iClAUs
2rmHN9KH+zra98VoWBVA7DGcmJOiU8AgyiCbPNy7lr11C9SsiUD17Hmm2yN+R1Z6
zzcdje8gZkX1cSZmfofd3HdOfpWhFmpHvWatvqmCYD+/xl+DJlr59ReSu3/3Qwtm
ErwQL8gI3p14Ad7hKaSJpZHm8vtAUmM0dlmMRtCQFI9frSL/PkwbB9gvJa6CSVky
IxRv/QULir1iB9BOdmThYcr+WXr+XLmpkSxdOdMvKmh7pmuNL9Lz5tTBQznFmCtD
Qnj2szwNPouvNuewyXssBjP4hRxfBGwOGwRYvz9GsqkOx1K+rginCdRghsHTxPNK
7jFklT4Nwg3yzKe7qBV3qnkIObPKWQXxxFYnTBcm6Z7VK9KdWMJ5duxG7/1wuG8J
4Q5a2udewsCNmIL90QiHb/cOhJV94Hayu/WEzhUc0Dh8rQribedlIBjfGpUz6Lyy
h/2zl9IHNsp5yFzSOAQdTuMevr9mjUq8TUy+ba7cBBiZw89o/cXIYENdgBZzK7xx
3xO+fYbDFnxoPH9uauj5js+9XZQCLKJQxexEH8ouk3RnOJwX+FqjN5dWB0UJtzD+
YA0F6zX23eYn6IY1cvbV1Lm+YCLmabeAf/pZhsYnlyabKYuQa8juWPu7//rwbh4G
mw/Peg9WLlk91QPVfOq+dLIagkEuW4FqWNy4QcQeXBuNMJq4CNDKt5Uyb6blu9sT
9LJotRsw6OoOfOFJrmPQio/WTQkKKvQBvRFrVy1TMy1hekBRBNvdqiHjB/gfXAlP
k+PdAwEu0qNdvSaXW/eogvD7YorpwuWu/pxHJdxlKX15O1ZSkQnbVkboNqgAkqm2
T4SWGulpRwYrIc+BdpudahvuRTEXJ8blFFdEjuYTsXNFcgE4g3nbrHoBp3BJTxBQ
Xkr+tJyjgkT/OJJP9HfeGRIJY1nAu1nE+GCxl/SzJz2ZVmufB/MUvdfdBEfQZQeB
tel2nVPY7sdi5yR861851Y6ZrgLt5wWKMcG2tjk+vWjRPEP6Vo21FL3i4I+470lG
FgYgp/j4eG45UsycjsDoFyrnLPlGLNqHi5xWCETcTPLnhWouE8apYUZFvkwXH5OR
HylbnWSozTjApFjBCli/odp2TUTf0z32FtKGLulkzf7DDSHA8YXQLL+CdzrP2pLZ
MF6bTJbf8/2JYpsl2VD0IC/kIUOrm4MAqkFUXuuvM98zt4etFmu8cS/7ZNuQskUs
62eYYlV7A36QIgG22wTeP+V72uDodrN2Rlfu3YlZxbeRTRUNPZQPAOhRMY7ssRDc
F+khoyNDJ/Z5jEwb6YcEKKuy5D42qfAhr7UYWjXbrCywli4Kzfn9Pkk8P/7F82R4
9T2NK7J4aJU8wjiNwmqXTU45JnUqZl//j/ghx82qhADW3FPbsVx7dIxAwbrcO1vK
g8vx8MOxo3TB4ycFlvSRWpkO0j/CB+X2N9Hfxi81tUFfkxlOPA2CZsn/C+wWDDhO
SF2bhFeIub5J7qFLpnAu72Cyf24STCbA3jyedfWOPc53W99UMmbeOqGOO2IHdviG
VNHitTw+F9UZDXGxRR0BZjT6vsx1yH8NqCGcvzTc0aMRn7MBm57lnotlMiKxF534
HPpyulTj5qXFuoeCesdsfxXk99+b/hYUyM6aay7S2WFnD6r6IY0ltDW9hsRE1M5Z
wRJYuq/lSJ1NT61VzHfsXEm12+/GaT0kUaXnivG8zNr82qepH+HFQChcM0uifL+1
UL8AGLoXtE2OFsMbNSXgQ3u8CEej7XjYzrAJzwmw0LfbYL/DDRy+flTT7N+XEFWh
MeHPJ/9CEs9TJblMikSWJvBGOJnXLqsIz8op3X8AcDlcz6s0S99h4ILIjVaNbukY
yS91eL4ipj9BYomCQOwC5sbJu11HZFuysh5NyTeyFDwkU3wJ/zpJ9orhebETXH9d
SqsDLPNo4vECS2M2zwXYBFb9WFVfXcIHQZISaOlRUuLocmlblhC74gGU7+rjVPpg
T4ImGQhiiOhRXKh1n1wHgd6QTKcBkUASuA0Fj7nnASSe4J2m8qv5JzOA2oSS2K6+
/OrzIpP9EZwebxE2HBpN/i4b+65cszQu4hfdPAI83MADzB67ESdc+1KgcaS8/pM7
je0p8Cf630tZ2viyxhdT6/uQzBUzGT146T+S22toLAGryYnky+nFok5C3AHxgXPV
2nMk0fel0qIbOTHjOIK6p+0+QKhVQWmjsVRhYq/x/MIrJ5/MEEsdPB3rdIgtvNPD
q5mCn6HMxJUJruM1ux7kmL3Q7eB6TUXlA7nsSw80hB2zpxyRFmgDsxeJaMrYX09Z
9HlNusXWHEx+qeW+0PfzZGcmvV96MtttrfXbPTj57wvFU3LlvT/4hrmNYx8j9dGy
2iJzRPWUtB4XtUkohGl08bQTrF7WeCbLlfawf1Yht6H2oN/ycrERs442Qcu9btNv
lAeea78qZ1LDwyVbpfie9suHQzBfQxTNIcagxh150XItQC+p4mYMyZWnm/HrCRKV
XGj/lmrGkfqdTwqsGnhWjifFOoXY9gVRY6O/ExRZ0AYSwXj4OV0RWiluwUA+RWmT
/jzGpB9cDABbWBc4qmIqH0/s+CcmuMgdsiU0Gc80Of5NeInO4zA16BsT7LE3BFKr
Yk/6t9bBUEscq75OAVHb3MWJpIfkZcFm5q9cksq4IISgO10BcoNW2erbqyxzj9qh
Yu+Rf7xbgB9D4Tw+tWeFp6kb9E9ZDnnSB+7ACuuU5H9cWSQum6Fmz1heGAmQxgW6
0XcuROOycAMf6hFRAsysU1yOrhqZJ3bM74ongvbIzn9jMyfm3fLLaU3fEZVM9TeX
KUZI6okA5TuEUDgdhFoMxY9JcEU2YkYJLmkcgjMZURJSoa5GC0ZGrGbgwBNVwD9R
6UYH71sgMMoS+rn58t7zk8rWUJd6+GNS3s/h2p0MsEnzQjPkmT70wbpfZD2KoGYC
5R8x9nilR33X7lVMjpemGyuyYeqOl21CC0xAV/Si71qNzOlouTyLFZjMO5w1xTXq
eZlxMcdzccGsWepXH+3sjCMYH8cCCnlgyBpeeyWMM/AhggqKSbmQ1jK48AzlFc1W
+bqii9p4Mxg/APOFwXf1m/EaYDm1914R4hOdy6EstAXhOxLPXF/YyXhVijxC2ePZ
cEwqyieFKaKmctfjupByzQLKtkXIufOSa85fCRHD+0OsLCwigTNjk0lh/yyMTZT3
WQcijrceLQtcrxNgFuuOMOBYAWqGYtflY8SlpUOUcmZtSQM36AQEG6KkmI1g5gdA
pEsFsiTBI95VVRQ0YMJCaUUj66nk6MDxG9sQ2qz1aH+P0VXH0d7JgEOJnZl+bnFS
73Y/wpO+kCs9nBgVwWPc3p3QVAQP+EiTgX6/Kxvj9ZSnX2i9IU2VjoFUvqZ3gLGg
YLnX3I/VQ45XKMaLcZNQIl07jb+exY7IP/baduXmb3ApGTr+7OU4VlJukkl2jzfO
ANbmvYz05pXVfmNvPourSbbtBsnGXDbZLcP7hWDmaVoEYp5dwU314BkUjcgFklmx
Nqm6sGlChCtvuJdPLNiXf6HYGMuoS7HzKuI7uL/DbBEPUHGoPb3IUz7c/mlonbYn
QosuGnVU64I29P/yVYirqkSYMqLvQpscDDSjDziq1VdZFP7k2a6TrK4BYVGvh/sI
KQ/Rciyf7/3FIBRR/iOV+5wNwQWrYaJewERNCTpwvM0DTgXol2WV+C1/J/otSPoh
zBSEd0dSlncmrxl8z+eN6Q80J1yjl6rZAE8HDJJ8oEV6YD5IU3VIT+owBdTyMv+O
xBTq80yw8TEJoJxQzBNN3s2PgInVgcwqpr3DNqJVzlMioG4+mjvzrCLdoPzUXM3q
xjPzSNqP+4lVKDrMRsZblgEBH7r5vsy+N30YZQPunmlWc0gVqr7sgxMzIBRlDHme
nowc911IQ2khvJ2SfAzi/wTpjkqEU7eNncGoir3KZ/1zm2bkxTJSsd3suzCkYSQN
Ryp7c0axc86e5wN8iv41wYthJIOJsZd2cze6aMn16xPln0+uyySytaXMPzo0GUOh
FXgftIwT5PKpG5aRWwCbhGg8dZrZSdTsGVNVuacMJ+fbYIEOjxzWtYgD/x8YT1Co
CsUK6G5ErtzDciWfkVCUD8Z0yjK6QiqekDBM8IL/yQ7rWs19q2a78/4ns0ZUlXGP
gp8QZ1OvsK4hoLdDo85PRDEJ4dehY0xaHldfIQv4iSDbJKhuP51v+GNoQcVYUTZf
5qBuMbu3M2G3jiZnLlDeVggDksBRNfMih1Ng3QeP2wDVBM/5DQ+SCyBzzv1BuVjT
piPVEg6EH2GA774Qi+GE2TQXBvECnMALhdiZPbCygusi50AOtoQrDJX9mPp7V0GM
+wI7qpyzTz/XWLCwHYqLqAIt0qVeikxgj/31vu+54yVMKVm2+BeV0gka1UsRG2HF
uB7XxkaE1pKIaYuDyCmIgyN85u1VMhPHFwho8EdqVsWBV1V7bgALnkMRCnQfqPIP
tB5Z8IIPhbIOxhl2hex2QxiSj5fbM5bHTEGTl2JLxeNPdQiYN7X5Xx1LrhWbesrG
PUCNc7Xk/rjh8wF3gPAwlZKsGKSDCJPCFFLikNzO7tddOLC5tjdri/2vHM7nxHW8
1cXWYpJ4cYYnzwmmFP6gNcQLYal15sa4FOQwhpslBE+T9FnWBOxDiQqcPs3b7mGK
4jjEMyDN5jC/Nbzv4sdNJMNgo1xPtJFhPUyhluI+UVCT2lKD7+4vJYEgpefujbMr
YFTND/haG3Ui0LByEGyNQrTjcEyBQ0dIEavl/bIHu9GTEekCoAG4Qv/JVjwLWQtH
OysqJkkguTjlG8IYGtiwyzt7lEihqB/x0WJql1R0+j8s+doP5uT+lNJTEzw4cj2i
GUEJTaNgLFolFJgiB5gTjkWJG/tfeOQCeR9o5TLEwDZk4DzGqLNOIpXafrmccLJ+
6J1vUUbZuMmBTlX+QX11o6dze7HxTpsd5eDkg2QMgHhlWEXV6FHb9sDSlQIJKA4L
P1E56Naa7KQ112DV4m0VWJXrGW0ON4CIL3B+eYDWxpXscOUbE4Nb+5R+ydNcdmk5
DOZMr/3ItP2ytnYod4t7wbtASP1yx4s6lvS/PlWazCo32q0uJ6FLR8ALAXR7a0wt
Ga3qsIG0ytLmRygFIO5nlfZRx5ONiHbU3KN9I7/zmwrp4GCqDNSI+B5TEHOnrE2Q
Zmw21viKAru2kEbpOjMyAmJ3/BFFBUPnadAxwBPL4Gy/B0nmMMnFQza+HW2jcN5m
v8gFjevHQCn0AIZhk50YnPEZeo/NrNNJV46mKUvuitYsGD/Cl5tvkblH2eEwIoiY
uvBh1QnoyBB13U3pjZ59JqrP4TqKqutXB1xKqSbeKH+3toBYP4m5aveEbaMOM9d6
L+l+Vi+uly8jwAmf5s/zXFUFFJqrbbO/ZXwJgCIXMOYqFonVYCswg2DzDZagNrDk
goXLDBhdaubJAy5bbDl50g52UUsNTHRF4M3UyV6C1N8r43sSfDEp9zHtRBwNRTBT
P+f7Ib1oYbvVEhabM35pwpKHV5ocou7Sc1o8SrGNKuj7JvcsxLOFaybUflTEP3Qr
nPD6AyxLO8y6v+35L74Wgm7gV8YEXRHsT4u5SGDvlac3MWBz5AuaULLVxCm7qP4l
Yv2DnxeAgKqaHSrwsgB3DYuj0Fu3Gseh8cuBw2E5fH3qoUgpB/MGJembR09o3epy
w5LS1xB6JPvjKniF95g1qY1+zgMbBm52SoOrTy1Nm5TiiAN1b2qIg3puLjOhueo5
Pax2bFpycscIDS9VVt/1QkUIme2aV2WXln4+z4hdZNPHpel+947mShrqnQLpIsOc
Wd9WrjccWQcwzy6qozYG8IdrR0E479+pxX/hQuBRwLojJtvUf6YKCPRdykybzvHi
vO5QC9jPopToItJGBQg0PE3O2Cfb/8tMTjq1by8fEhjaTwPggw66B5uUszWIUcXf
4XeCxN0JpDRVHQ1uReoV+xEqoHZ1ms2+1PCGyABfm9EQQAVTl1JTjeGtu8yJdUfc
4eQ9MZFmSsZ5dcnPiyHrlPahtoo74u7OtsqUMF0bTooOPTE3W05/PXt7DIwdrJ7h
ERhOOutezHMZwYE+cRFtJ0iXg6PVsIQvrvy63ILTABMxXjedk6n9Dv3hSNE37kTO
Eeo/YtIdTxtrHYeoFV1rFngLwreXCJ5O9H7G5nlN2FO8lAWqz975/iPSfEuPnpb2
ct2m6VgYmsJeVgeLZZp2yQmM84+h1SB1l5c1fK6ZWB4PD5QhVf6LO0bGAcImoN84
Pp4lNX7tdZLXmI/J/oH7/s9uOOcRReT4RLY0q7b20oxVIMCSXlZI6dtunHN/PKlh
wxUY39LLTprkZkS1XUxC04HonzmAHSp7R9E6CSjxnX21LHQn3b4+6eZX2Ftt/t8n
tfn4tkShFqGMJ/jujyqcQqLJONWLFQMDqLCA529p2Q9VisJ1LAu18hmBNChi1PsW
AtvkAjK5DLLstQfJYxfWzoHgCX2SjSriXduw33uHKgHSJf/Vx0Rw7F89H3YZ0Qtt
j6IX1bdUeHyQ+xpFKa2TFXVYJCGmwqvWjHFhygdhgpXqGczyq0/8rfj4f6q3oSf/
ayI7E8SLB8hWx8NIid27y+OGRiW0it4jDPJor3ASu82H4g+8Mnr4l5wPkOHb273c
CKsMMMW3dpWvF5bcpb6r+p3qFNsTganT7ZnAFXVNtADVAZ+a1JZrT64AGJpKTPO+
ZhOXbY+x2VbBl9aDyTsbOU+4uzmylIckL04jeIrUYWCtDm+RBlK5FfuEgIunIJoR
+QojuGJuXpCY+Fo8EMctOsnUomCD/T42MRd+406uSD9a+vCGhLnmK94ZYaaaarYF
9MlHwmn99OrHrFF7klbeZoWXl5Cz0W00YAV8N5RoZlD88ThpxiZFrlPyXCS0Zd+M
f5Nh4u/PX9rFWXVLfPMb1XXdtVuX3DSuSgdFszsfkmM9lJn7qUQOGGpLXSxgtCU5
HSUJgb7ZSKO2/yiki3QTmVSANNY/lJKIfl9VkHokpPEKDcxyw7NK8fFqSuim8zfl
+sMlC7wHC9PFimJNJ+Va3lquGVNBB1WkkL/OvqblhpYAV6RFBC+8xpUwCit5vqik
EnY0D9bgMClyZyY1uzL6FIJjsJpKSxDXrUuQg2ubOU0TDtmMjX9rnu5z95gsLpOh
zC7TY3YTRsq5rJUowH+qK0SoKA2DqdXPNQFNa5VfVnFpdcnS8Xc/2s5MB1RhAPHJ
aqRKlx1vEhuxT7spI3QYHi9/VzoQhx2lftix5vkVEGDekPJlBLnjRtXv63Y7uLHi
fYkDz5Fl6PftpSHWT6OE7rZN1GaQ98XeqYxWVDv9/O/TikMfjOmlI8zN7+Nm1lCW
6Q2PBNkYUV0u9N/rE1MXpzMVvJF9rxPaTgxrgv0wr9r/O+HpBvYBG0cjNQXs7RkY
CfF66TuNc/tC64qk5XdWWeQpIyk5g4U5DiW+/JHyIYfuQeI+jd6lNTx5Srz9Dsmx
TKXDn6kJ94WnxvF2jW40pgyACOnW4Km10i+ioZig77GZrfYb4Yf6KWjDYekwTYkA
PDm2rsA00RGBJSWYSWOVaJHB1nm7Xoc4z3ModqmR4XROw/8wiiWi6SVRY/3MnOzo
NruyGMQ2OYGLIgOYhSFLJDZR49uts8OuBcZ6943RhDV2biZDyF09avPYzGdsPiHS
j+D8Qi5+WJL9wGLorLoUQGpPJdl8zm4eOWUeBZgxeNVERvcjj76wvA+N6+B6DC/N
Alh2IcYfQYovJv8/sKtTPncQ3QTg/Q/us4l0qwCkBDeK4I9X5Wnpx5HvMRY0ZuUI
FXszuW++Z5LDue5o7omqx1EBxZrpm4MdziqN7MDGQDVfrQIJM8jrUY+VdXVOM4E9
MNj6M8K1H+mx4gEA4Whrt9t89RfKRG6NiP3prK37E6VwHgyo97NhXDMJXJcROL3z
DtFR7JfBQYfCFUb6+MEvd0NObuzx4y61QdVTBt1q0n3g90O/6bbeK0zLKHWtfEA1
ZdSzDhpwG6dUPkcpcBnpALD5tS8+7xRyQNuEc6fv+NdU5k+DevlO4cunxLGirE7y
C3qIi81/bFbiNnvYuepOi99eua9JcmNa0avOjuSyllEFIT4CqgiVTyOIY0DD9pQX
iFmbyt8HIiSWcU/sPoqe9QOVzS06Gs1GYvZDTvaKPU+R7eg9lMb6JLPyf/NHg6GK
6ETMB28bXP4tABFEhuoLV2lv6wY/32ITk+IR/yLKFeAj9VW5yi7fIa2yhrvVHIXr
G88yFtTVT0wdQTKjkGT9ZthhpHh2uSv6NVS090r1LC+taH/YxYBm811ckzReRk4Q
HJKEF5dNZQI4KRdLYz4hxsJxVAAHxeqQF4eRJ3wEvXxcKSS6aJ/bduZjfB1jhvyL
hocMYUfaK1cb+VyLUQ/YHnYPV7ogRe3OV7OFcNTJOs+hSq52MTFEMxa29dF3Syli
lAHcyntHgYvzKznPnTCjeAWfBQwXdXBa6I8zBLNti62LWQGL8EcwARGCfVsimLBN
TvQl87bdgbcfBu4iaJfQKMaPzCwIYkzeHXO+ewgoRAYLiUFvDqYnHTy69Q7ncTBA
ejsNBkOPqiNyHUgpPSbsyyletQ3assmoQ+X9nKb0WXL4yAXMI+sOSAbCNA7+lzeC
YSPkF26nHVHiYNYEOfFWsrqZTPz8n72tz/geaBCzyTPe15oNf5iKnAee0oV6KASC
P1njQ9F9qiVo/fBZ0no0j7Od4k8MC/gHGSwoFVdQNBzzwelGb4ewNABBWx77/PLd
QtIX19I6FCCLkqN8alzncN8RG1geUgJAR4j9eAZ4PM1rgBPKMWVEN039ru9PWYqR
TNCJVKxBTx9ySTUXFr0CABMkS8CJQzQy6TkoJMW3m8EFnZXnjI9s1aXZk8A7KVR+
xYHn7dyaSSpULeStmJWUzwSxLdHWAKA7n7xBjnhbAd67BkBHH5IWqSYVG55Eh4o1
WjKV0xe4DPRdceCbyowVaucKxLVA6W8hspTRYDxRqkzuuUKCmGE5GzoBUuX2XnHp
LZrKqNLUX1kP6zy30KuBEp+XXzClvb/EY474YAC9rg+beIMwfaWsSKtB1Fv3mccC
DrbI4a0O4G2q8qiIENrl0a6Nn4DoJ30X7ULndCvPXTMuv45Gr5dc+OhqcLJ3fqGO
af1vPL6pjJVDq6hZWmN1EfhenOrhFWqAeUE4cpFEO/gerBXyD+Qsmbvlj2PQW/Ug
ilTpzFCwSVLpp4aWfUq9bSO2gyf1MRc4UqdLngNy7CoFnuI5w/PE1Dg7q6CbrZik
ftCBPVxMpXqE95C9pOrvx2U0/CPbDswpyGj4mbEQTS3wAYhK5WBLK1l2FbkIqkVU
XCSf5vPM2F+C0FTaKbK8RC+nCNwZvTsaEY1rExSnK+ols02oz6gDFx4eGoGMOsh1
ZhX3PKRlZo/0QbGk/L3guLbe6PsEi7TtJ2lg9b8ddxOXpTwrr8yT1Y1o9KxHAf4P
rKPy/CZX1Qn6RUpyQz8QxYcdWbCV5/ZRtdxJNuQEU7K5JwtBktucD+vKLocHbQ5J
ACcLtO0Bz/QjDpzAHE8M2FlDJJHpatROr8gggSQ3/n5x+9Nyt0t4+0/DuBVlO55L
GpDM2/9Lth+i7QEzbedz3Zput5xsKhItBXAgglE7JZOr7kitYo79/jfslkM+4N/n
Ss2vOw8TZHvPTaR8pFlSyc+5qXbAQHdDu8UCFnL+qj24pPJ3etFQBzwUSTQ0aLnH
k7RRWQBk1mELudwbtmAzL3iVWzocEpd8gyVz5160WueEamAqnSu5vL/AUomZbiF5
yMoxpc4Dvlk2GxqDAUs6Oy3xeGKqbU4FoUEpID9u62gNa7bwo39dTj45ANXz8ob9
TSfvSoZ9x76rhG+LdbL0RneaK0FoRrMll7onN45BGS61vnBNuJZoxYwx+5q+fDJ8
1418ccoGZ2doKB1gYebayobrEVBp6WvjU/bhnVg6eEja5zGp9sUKFfUDfOxpvqgD
nEaW6c8N4RDkAHsPQlRk86L+qcLe75O+nIgSSEXDtxzCoRHR8XwqfuXDhWEr7/Ti
iS7Gj0qNoG5Qexj7J8l+yN0Kcf3Jfg8s10Gut/4P2iG3j24Se90nmEfUKv9HLiFk
G/aXdJmTTpL7QDsuzClPfF40ZsIdjGQGL59kgcNYMZ3+B6yIdc22+RshNdG4jNaM
7oZIz6zNSujzjzlFS6RtUWxmOCfckZgWDjNeY1Tx33ADGbsEJKFsWCpSt80ms57f
W4wxb6ggSZHwtilBwIu4mupYT2rT1Byi7hv5BAlR5Ah0vF8jlbX2mq5EYJ+UrGfe
29nerjW+cBOmbJH2HAuSIjCwGSdO8nUWeeuHmpP6yj0RvGGAWVtAsqYJSHecOX9r
U+cTmVQHJg2g70fUGryc3TdMM0+syobBJrgKF/TihZdV/i1aC4F160DtN+vKCMkO
O47cpYXmWABmDJxnjQprdtayyuMCvQAZWUpg5/EiDzFwhLjIjyyfjxijoCrzn7Fw
qv5ImYBhdpV5WERq3iDdltSsGYqXA2gvWCWm+tpV26fSfuIgWrpE9+J2Ox8SF8pL
hWRlWuLFfAloMFpJgQVSy6mOs+fBvuphjj/ErpvmJXK5SwdW7bPrVAeCYnbdJKZP
rAbwqTrkJ/vsRPosxP0gfy7v3wHP8hTnvdWAm0yBu09VHAfyN2VSBVz/7dAKN0gm
Ub5BgtoHv0tA+cwUQ8Hy2Nzj4AuHYv98xrMsH3fPzdH6YB2Q+pe+JWiK7rw9322S
8lYOQeNHbTJObP8q/8d7KeyYbSDDXjXwYCd6APDB8a0ILTbD1xE4XfNMQTEDFNCl
Dj6CfKeEr03+8qWHngufefaAGv34EWMWrC0rJ8RDZnpzYIOqY0+7zWt6uzDJsxoH
Yl/xxEKYHnXYAIqBmEzG5a5u3ukHZY/wMkKALPQgPWjtb6u7zV4moWa7oJUHFcY3
NCmVrdzRaLS17Ajm5iH+EY3xLVrqmxcYq/5dUQOKxE6LoNIvFHaH1DYL6y6uJUag
aD05hlL/XTJM+CnXUSf+Hq7m4kxsmEs3dPPb6dwpF9J7zrRSPdrMbY4/fDBdIskf
sznnNW2RIGdSRPRWKqIs6ZPQFyqEcz8k9Sk4WS9hPiUqDDAAmTNjOW7GrIuTU4c5
Qq4iwrCjzWDtsSNlJ+hX6hw2h9+K7WsOiKG8IW5qArOF8RQ2EAOIH+Te0FyLu6MI
cE9UGQ5udeY6IIvHEtcws83NXKKYSQjKl6nMjxSR3sKJOFvLBw/S+jpW2ixoTiw8
Qn0pmWZ0BIymWPTKrKr8sMRIsHoWIQhPib7+pFBAaj2KkV+gJ19KEwfXv6oY2vGU
NdfB7rtYzUOtpIr8CK82mvUMqSk9ReJEaHkqpiDnSBMmFBG3Fd2o3sdSEwzc7Pbg
nTZL9bFwbhCrMvybjL7PkxualUTLuDPnplCnDVEp6GXyhwpeEsraFjoH+6UP9Ea+
ah1bN1db80gbE1nJMnrzgrQpvJIiPeWuJg6Yexp7ABSW0V8Fa6GkpSSttbZtUsMH
e9sYScXuXqI1ydTm04RoMwakMVN3yrzs78+Lxla01/mZcHt33EtQVQbMMMIby3pt
XwVgNDvAwcbjekL969ynRNqBS8xSm7pSSdFi6CyEqe3kvSIPTo69aXNNfKLkbvZg
RR/oPoDArZLqtrGLee7udLVgKlcOzgJ/qmR6jriTHU6/9NK5cVaIEbwX57ZkOj44
2dRTkUDYLz8W6lp5oc+sh2avJSFRA9WFhsRABqJTqbkSVF2xsAXCV39ffr6NeWKr
8Z4yVrfGusPpzfJh5HtagSqZkAzfzfcJchKiDWQSiu4pnfi7DP3kMG/E7+hsJ4Cn
iAVHYAouOaD9X63TuF653ZcBW6eg5EZyn4DpsFOroh6jetk/RzIbmZLFy3WPiMbU
5IinRGwx+1Hjw+IdKYJvK8OkzzMpyhjdBxwZmEXKfBkeOU2iEx0CaCoG5XeazfLP
+/z+2BW4r7aXkUXJ6rc2HvjZB7RVO2YsBwp84uLM4LHAxlKPynvwERDMR1TCY+Hg
yeDoPTi1ZcbHgddG8c74czseceEuv/JXwETN6/AgNZ8WcmFGL5gb94dylwqoA5Qk
dIcjoxB2TVdhl0RawVuhDH9AJlBdCQ9ZFcfRpEiOZ2sWcZmeifVqo5hf61OuA8wU
5gYvzxILwx2lwHte6oBtQ+v2dvBSn8/NlhIBi3/vk1WK8/bKg02oH2Kiwzadz3Pw
/omWjWVMZuilv004aSs5CoJItv9L7VMsfIJlSN89ry75srvfjvXlQBW04R0MCmUr
SvjjFywsW8ZcPpp2ndGSRDx5V+Ql2ZcQaLJwNZmVfZM4O4exkmUcPKFsawdWXGKL
WVIU3MSoQyQpcYciVg1Asn8nGc95cO8YndY/n8IxQvi+mieF/7rtcApKvXDFr65O
0wdqUOx3p9YaIV/DUy5k6/DQl2Qz7gH5GUHMK3LOzhEeSIYqhsACT2Fogj49cJXH
kV+/0S4+U6vD/kwPNKIV/Gam4hqg5xqu898WbY9Z/Wo0lDXdIZz2bDYHA2C7XA5T
KFstyqhGujpDsRfos1L4+0mkgJ58tG0FHGAJ6q4lrwwUpjH7bdpjfyMWfU1Xr3mm
tOEudKqlVEPfIPSpsG/x72pvVzCI9suUJYzZCE4EcW8gl1hpQWZcZFrXdyAcvkg1
TVAqDsMyxh/1MyChT7zWav9Bob5oCPAv/f800CZBN196OttxZKMk8vkGqZydHga7
0KFSjwTex8RJa2cgeVljBOBIe12teterdlUO85tNLoQxsZLYvH3HGPzpb4ZhjxAL
zTgVO+bcRiue9l05t9766X0iZ0cJU4YGk+jkXRsO7rqTx0MUiXUelUEgCFwRfR3r
mKJVeDNBOGc9n9Sj01xVmu4t3ym3Ov8hrmdtr7iTPFlqUhs00IyX9AoKiCIt9xqC
VlcLw+m/en1T/f9IppZzsrCTfpy0hlJLKZsQUpgKZvQEuqJkdCCL2PNuS4bePhSQ
TWMXVLs2zccyIX/a5JAg38Msgwp7uIU4a+6aN8OgND72L47xYuDJfslcsxlLbnam
oCA6Pff1BKHALuf8jBbO91brdo9l7+rlcWKYV5cj+Z2XxqXccOt64uzENV/5bOUS
zULf7Nf8fXixO2W9+PE5BekVUANQvp26g36YCvvDyIMZAHpnZOGYCDGodXu2Xj9U
m8nVMgZ/P3gZErCfStrKv7NldUILsdkdCO6xpQlJCDaeLoMipFGiKeZ3dcOENJvU
scdvzv46tE/fYIzVQM0ZNvzL3x/lgS8xI8lwDhtHH0hlpEGADWkupQa3/l+gse/7
+beuyKe5PPBBq0o5UtCZUTM/F2rDvgvST29hSPmr4e2ufWQ3/yk4QePK11ZRHzy9
vNbzVhFTMr6V/MaWKNF7hRMmOt5L9hm49GHaQYgxu/ePDRGwewhDV0m6n3L17NHG
xdKH007/QbGShHoOWKJbE13cMzDNYVVPXeXIVpKQm0ncpBWs2rSbssRIzf+I0wdf
oFuDVJREtQy9YXn4izzzhv1/TFAkF0OoY15NnbX+RrL4cZyN+54p+qRqCZrH7pzw
PvvFbgHiWY5hsADaBJCSyAzPOEGojnQO7/bT+9QfgUi9yR15rAfr8bHMIzkpUO8d
pvZjom1eh9egEcZoQ0q65DRqH4LPIVRWCiKLVBFXGNN/LC98qn16mGCvwe+fx48B
SeBSxieHUm83m34046/J1xOFZ1S6PyONKq83xPDKnVoSmqVqCN981hsekpSnob18
viWq0UY2TImt7+XkDjXsQiOra3rvngl33VlessNmNpuMPGrbxphJ3eqJzq7dy7bU
g+Nr1URorHY9wDA/d8hUxt3xDs20lhy5/KWcM6sPgDEQjeUQrDBjM7rj0ZsP+vt5
1XFgoIUKHLF5XTKhhjPf/KIZvRCRQ4c2ueaIu4Di+fp/EwDojNW3htGoDTkB71Q9
PinNSctFVjWYWQ8xPNyRsSzcDzLMEg7/xW5RHUKG52MpEiDMTTuYWSn/Iq8j20G9
t/rGBKztFeQAIgBbPNR8BmsM7rdP96g9/i2RcfOQ7L3HDBV31IqUSITWLfgKGnBA
pmd8Q5JOPj5N0zW8re/w2HjvYaGkvRe5CkiO3RDPMPPRCHaSLimZkaBB+2JrIfqA
uiE+iUZMV4vWw/UdFvqnAHGmLzze6RAf1hyGiaW9Um9o8cVrRtVLXBOXSZxzg1ch
OR0bimC7dod4ZB7ZVgiCdorDTiyABTDp44XrrvkpkW3tpxz0Ksp2yNn3DK1r8xqa
cKKbCfqkYsacpWrc4dhtYoGD2/j8lDqfrzN8S4AQE10BWMKYWuPzaNZVxNJshEHf
U0YFVcIsFqV/mHXkhOAftBiRCYAkLpMttXpu7xVYaDIEernmxDspmPphv5VvE9EK
CR8VogVqIJw9Omu6NZ3OVRPvqrvfaLv2W5I6qX5GoqsJ1STozH84O/TZQb3ag+8d
+aYrZOotO0tvdrWAJGa9DztigC/oalBY6PF7brDzUTN31aRwPubQTgDoT/7nuNeV
JaMB26wjigvhpcZw78weYGeMNjzuPNGh7jb9EBtVv6/K3Vr9tF3hjGAYKBrhatXU
ilT6tVjL3rqcsTz+Ie71j/4PfUUBINmnvjGo53HqAoSVCQykkMQg8uFeHhZSlGDX
RH2r58Nb0ezXKohWz2S+XcwB2Nlq08CHCi1megkRywPX7TN9BNYlAGMw1LhqQ3uZ
QHfNPZjv2EbAt6kdJ2txdbcYV96dDoqIdot/lr8K6eYklavpNae+lIYytsz8i8dB
OZBeG93Ofiyj4c8fbXsZgoGgDjlC67XhPhwjhrA2vhc2Ffed9mHXvN4SAXapCUaE
+vzPKAUzudWeItgbQbOG5l4MC+j47nI6GsjMcUIK6z16e96qK/kzyGcYYJfKn7NW
6g++8GciRx4e0T4h7egy5qnncJ1dfC4NYziw0TBcNDf9ROxxyNq0HjsAUwbfDqnM
cvTFgttaMHVwGa3Bh502N+9wwpXHejL8TvWgnNSeJQxvh4XE9LMR7gvEM9A4G3qG
8xqPBh42BYvHYmOxMQodJASCo7Z16dxteVyHVSayPA2frx5Ka2JSH+EBkSdE9js1
vnCiOUObBdFioOejY59gWtpbrYqJF/d2ema6BsoEpFHVemJ31rNmBQSVRZCDTetw
E/6PF49PerknJKOc3vyc+SqYlrRdX62puqc7ilbaGaqzOZOdWrwTd5cwjX04EwdJ
6Uwn8gVlIx3OGGF9Jg16Zxvd2ZdXrFMYm5ltg8lF64LE8K3tJFwNe6eFZuPriJ+v
jpoMU5ne8Y8Sap1zenqBxRDJ6dYnZJayNwIG6vXEwEUMOT5XCa40Ko4FIvVDO2k2
E2jbvaLkdED0RsyF7m1+U/4fpBSvi2gn6CuEKG6GqJCNxsUHqTYiWpOWqYwh1xO6
BAZwLnHaRbLVAFl9xhzrdRVwbkE3iPUULBlJlKtt4aN3ZMu7P3FiPswg6toJ5aEi
DiDtxi5y9zDA4Pi5j4NvVED8iJl/89Sc5Dn3KhOnhOsjeGU++8OksRkNk7q0P8lY
Ht5aex3A8Kmbm65bTlDugqMCq5D0Hti4aEpM+8yWwFMebTB0wZYqJ/zarR5OYm6D
CMDEmKzYhnrN/kV7znGdBS+kb/tsBq9m44ltuxickORFhc9vVYoq4qT9R06lGeSt
qgNnoX5C89XmfYWmMjBah1I5NrIM/gl7bj9IytRXtjPr6HHK0KUMAfBTMEi9FvY2
kbudnuDgS+oCw3EtXprPF0b33R++OnKG7mU3BE3ExOONfuUiKa9hELhEUzN5MAOK
fNOUC3hnPJ3QL+f8VtoXKWnWbm625qSHsRCPj1ArTVnImswqfb+lTnb10PtQnkSo
FOJ+g8Q6L2nO4KYNsBB36RiqfZ76k4Ycdm2twyKmhI7mdLvE1XAPSb4V3tLmngx3
MG00aDLUyR3lRPwlGliapYVd6uU6Qk+WLfP0N4G34l1ruIwLq1ewAfoq1xnJSrvX
PHArk8rxXiFuOv8NEx8K3WZZKm2NtwxMwi4ZrweYquG4zEgpfxoJ/c+vL4X/OW2S
2htowV109bWgtk05UHXVEjvCb52NNzZ1w5BallfF6/StXA7gwKJ8NXony3szTRlE
4dYnMa9guDR9HHuRQgEK4RYrQSSARXxu9Xtu0UV5B5d825SE+kb54H2FUZaGF3dZ
+M6QVcDBwwaxglXxVBv6QQuxCPuEfwbcN5zsJWom1eCvtXLiaa/f0w5FTU3Og0AA
4sw1RQMZJzJt1lKmPb939Yt7c/8q4fSilO/rkTel+USeZdmQZg3JBtUROJIlskUD
VOxwabMQSmIkfnd/e3cu2zeYCMc9ScFWiSI7NJRzFEL40HZFF7MeFKx6T0q+Crld
wFhwKt9kYgRtv5gjjFieqJdsGIHyJCVLKTdBXuGZbstS5KICrmI9woladOQ1LbZQ
YtW3ABlL18FrMsUnKkexU3cmzl0T3x1PVt2gqOR3hQzt+CKVDAV9yNDlyl50FOt8
QeNDrfV2sG7GmSpAHyVtYFHTlW2xrkKG1kq+XiZLcR2GgzFgWrDIOvi0gReE3BDP
PB7cumYPPBG5d/e05yUw6aXp3bvObW86O0HKmky+0wIO48g1LxtShYtCJhnayEUx
HVEAc7tgI61WjzCa/v/HBLFkRjlxRRj3A0+8iIjup/Fw7nfiw4+5Gd1GS32UkuBg
63UcjLKKvvxyiOyeX479LlKNfn4mCL/dLinGzbNDzffMK7hzzRdKxiJXZI3lc3Xd
VHndpvQbkMcG/FQEwby/6rgCnwypsDm8coeUaBmPJselRnYSzH1R9vC4r5nuxC8D
Sxz2fDKPBq+Yg/c8l+wHcbJNBFmY6p4dP9CIRZ8/w3CwTdkb/5NnYJvEuylPd075
DFeIr26MKLZJSa7XD/c3Gg+lGf+yq2hYbSLxDyWgbGg63qJynKXPH5FtbuZv9jgP
8LXNcH8aTUT0WHSjgorbpyL515DtCK4+HrUd4iHX9++P6F9yMWdVduH6rxwsmye1
BvczL6yttGxu0bjg143Uc3G8ZxaHiOMtJNfWsV2+J7e+xhA1caYeu7wNAFtNqWsW
hmoh+MxAKbYKfWQm6MIxFVcsssS1l20SEglCa6E8zIJ3eSglc3SKs5F+UJx2eAHk
vrGqSIN26+A74WC7Feg+mJqRLdbAI23r5yPrvbV405HqXiitZMiUPgbWJKHIk6Kt
kkB+9bv+W1tNc2oYBvGOgy2rtBy72dNLfGiGBljWsl5WfycYrwSeAs567tXCnmM3
par7fWTK6jNpBJn/esAi234khsPsOxOhZbTp/QMEZvJ/VqH350qS1WejE/OsE5BO
Rkq1G6X9HuBxNbkKbhdl06joVZazwx0FVtOPUrkrz7muzgDL/O8KYBscKdm4vjcJ
newjt7JbO52ASdTKbiarqYSXrYXvZ0ek57n/x8P0AnJHCX0D2CMA4/mcTNjI3qFa
qHts1ZPJyedmyvPZkMswgUQau9fWUc4HJYJtihNqNapNQAkEo/bOKQa0ZiF1oayK
QLVThcgrIGZJoEnojItvAKGKaqrPChL/0MhtSA9u6NqcYuui8qx8nu2LCequZKRT
KtIpgEE08QXK1GX9hDrFc6i8IJRSptAY2CsqCboLz1qxnMsGpkzAVhzc7IsSrOmg
LCvP30XRzYC2ug+bPkURFMQzIww5Z92tdIdbsznzr+ZEpSdF/p0OvauyXWx5/No4
0g1wTbG5kiNI9qCeHl76qHMScl95YskN2tMPppn29ao0VFgRHUdv8DOuN4IZu5jL
KYTaIMWX31d6LTqBdCdmC3NkWs4sCZGRGgnMXmKmf6MLg+v/pXqOx/CEJzL56CXt
Dq9mTSv7bBhHw9pFUHhFldvZ79EhLDjs6Cj0gIuaJ27bOn2hWRS6pQ33uZm8CQVk
quJjwmudoeJI6vOVZzp4Gn7NmqREPJo7GdBjCSCaPADNM4xRBuFQH1J0F+85H7f9
CWSwSXZ5liwcj4A/TfgkTCzkcbbMrFDfnuV3dB7co05fUyvgcr3I6SadwhNCvjDZ
rnwtT/pLZwWG5cgomQWCL3Z83/hqdHnSFoYrSAcRbSRRhWHFRge7y4KXvi+wTFRX
1RZbaOGzUoRqMSRCnKNp+xV7OdVDsDgZ+5EWeUTwK3wdKrv0YYwDC7vz3rwjUzYZ
mAIp9IMYLzLynFdLmAnzxnvZDV/ZXcqc/6F5K9kUeZsB6HninAaKqz5gNbwfLzh7
GNMvxhabN4oM2Q3vdDdV4bQB3eB9HxkG4wlS+RXagKKOOfP5BOR8kcPobJu70yuw
+tqy0mDsRta45H3UGfU8kQdz/tUShA8ZiOe0fH0fOplKEuWIpmPOnwXQdl7jT5Tg
nQKFno28TI1wxKHhflkO7M3UV2n17G1xRo2byZfgR2uT35bnWmcGD1LwG/AhSg/8
V1dNmRoFhtHDkr4qSfggstgRja321YuygboFxREx0LQneHE4rXzw3I2pjAmypJ2y
2MOyrrMVnneBO4QGKUeacsx9IjXv4qbI9eAoG01BiJObwsEzQesjl+FuM/bkTVNA
fXuJRJJqeFfTWAq4I3C8Q5ZZ5TMvmszqFYIRCu8AGc4woQRpwABNoSltwVGRA1+O
OSwEh9OnzIrGcLkURR1JlfHDD2oN7UAu5CtMs3tr4YPfSxX4Waduf/a4R7MpfFQ9
DNzsApcsX3pCEGwUKmSWX4xjINJzQMJ1pC61RVz/0lrZgozXjq1tBRBJ42/HWSnX
ucCv+eldlebPg4ikPpYLFaFMmCsFI/Hx812FGzv++tfccxPF/owf0VQt2N+RCLS6
+yDkkowLSpWq1IpSix5DcHEkD18qBbdkTkCjId6IIPK3gjgVlkaCzFnmMtwxNoOV
BVjBpqOxHp3GGnHcH2KXjSpr/cZx5zkkrKDe3wFrK0YasMHpVVljOh3qOz+HH1gK
TX0Jfd0wHZrCL+l3T4jis2mRK+tFfeoFwzPzSinpdfwT9HIphUHYEsWNj9aWnzB7
AnihHI02UPdXdK3DyD5r4abHpDl2/RL83x/IJKtFQO1kc/jKVpL7dAgOtxmxVpc7
jI7VDk3OZccQ2dZsgBuT2XT53zaCxTmBYife0c6K0/dLRoODNcschujwsNdkrLNP
EpJo5muGeAhZOr1eTJWsTts1Y6o/J1Y06DvoHAhaZrgo/Vf9pKi6F1HC1bLDPizk
CzuCiMHca6jySVffh4wDLtvUxjGy82h9xED7RGcKQGR8BSm3G95u2ImdaZOdEw0g
qpzQPcX0yFogTH25YoflV0h8c0EYK6H4MWsGj29PeQ84lO2FZr0Mh7TaeaxEeQNw
FstIaSK1sM6ZdMptVgcGrdtNEyYFbOIt6da2jKSdJOMIyBQ3X+9bKhhxnSr4NJCJ
HG5ojwgLW8tjSdl/nEHUmUJjzz1a67ezu2p1OAmaftWpYQNaBezp+a1I9RT4OXSq
LbN/UQY3oViGdZO7K6D8iipJxTupsX2nrTCTuaDyYdSZWv6kmVY3E0tjNfqJ5Ewh
T4DXKCEvPycst3mkHqWl3yx3B3f6l659/S/FZcSVD3s+uEUcg/jYltfYQKMEWmfF
XYE3E491JdhwipmTdlxMaC2OEorsr62iv50t8ckvuWoEH1cUh4KtBk0w57akjOL5
UQQjD9d9oLNh6fe7P47Mrg80pm1JBh6PNOPGtMUkNNDZeoyseWCJKUEFTlgaNRU5
rY7ujzJFc8IKwiDmv8p248UhSQVjB6rt/ObcHQ1/wVSfmGfI9lBSGBL4K46g9jPr
veRvqMM1XaYtVSD7gZCuIHStryuDiqZxXH26Sf3YfsvKMG0SI+/EgIjWLBxqYvt4
K6l/UstsaT5QOXgrtPu2Vtg31RgF1pBuHRWA/cVtAYNnslEPv0dz+NsjBKYOAduu
yRT88zioaD3klKZ3WqoYO+Lyx/cJipf2RYym9qrKkvu1o3o19vtrE4hanEtOoEMp
f/U5R2awanfj8BUbmx/ITbLeCDcimXvnwMQqoPPa0o+1mhXxavs80TqlOuNJm/kg
/934QDiG7iJOMUCghQUUb6a7QsxgN+/xESgO6vaQ+ls=
`protect END_PROTECTED
