`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/Gavq8IszK3Nl3RX8TJzjtKMWYlxhM/fNUS5S4GWsu7LzDAfBsRYPI7Op9EY4fp
njpqEoC7B4EDOxYe8HCaNqiLCYKgrL0nRkfnRLaX4p8mJDyvQhJlEiNcxixOg/At
F5yPPlbNLjLGRyMdL7F1jUeYiTX163cFRRfJ7SOQLE0YY7zX7EcLDt1yfkjOc+rP
HgUpQ9GdjK7VwHffSkSRoCZR4RUdwYnoocPP9b6DQpN+3P13E4ERQiR8Ln76AanV
3j7yk8H4WD1o9ypsS3krpg==
`protect END_PROTECTED
