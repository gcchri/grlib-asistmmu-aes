`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xVPMhHTCdCNmfP9ATq2xZDxxfzNtwhdZ9TCqnGqvAkjoVA589MolQ/vgZMrCse/o
+ESUxqDVDcs4WJVmUvL3q4s0EktGqItXQHZAp7q3QmhlHB4N0KcRMwzlrozWpcXu
9Gk+6Jk9CuY7ro9Spk7gj+MP0Knf4OZvbgr3IDs/j2RmneQelZuq8BvPG+I96rVj
tvg17FBMa/jr1/7ko2jveL0H6NcutbboN/ApHfB8BiP8LOSYal6esXntownDWWTp
bHFW4Tp9Keugjq8vTZVJqaR8rib2p3WMTquAW25ue/Ti+8O3G91AYL8FzHoKKf0T
NznRIFlKFM6E6/3iwpN+Dn+V6et1KxSifp/FuMlRNBO+/WlUQq/7D/VpGU3zQdvA
XZ3zIE85ecDJzJSsv95zwg==
`protect END_PROTECTED
