`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
41wUF1Df6FGmMXyzlsrp6JvlMXmd5/C4yqEfAKwQGTBIWPdOE5Kuia9PGSZDwT2n
bu8jRQE6XAIIaqH81H0BQPSAl6yN9/k9pgr9XBbNNhZLsfdjma0NQaTH2GYgwmTt
1QCIXbdvUhdnoJX9mPJSvCrX76XpuWedUW/P7U3oysMt6oIKc9qzfWlczfIpJiYl
NMuPmTJttJ67IQEcK4gtdjfLxHKqa803JOZzE1bczEXxsqutt2kM5MZquATWOpD8
4aR2Ibojjx8u2LMzkI2tlOj9j7nyOl2gHddnevwxup7InWsO0gOMEhHYf+sjArHe
hW2VMwWcUBChnIPEjG7XQ67N0ivTP+s4ZbPy9V/mIyc2nCQIJPekSHcaOnGEngh3
MwCPFCLMXUMFwys3qGnpopRkqqrnqWBpRyBJnFJQ2yneYslcEM918Br8I9U1a0Sq
zzlP/C9pWrhilm84Ztbo501DXjvqbjwBYsNRskvJJ4pFVUytAK4iBrGCRKUYZ1WL
`protect END_PROTECTED
