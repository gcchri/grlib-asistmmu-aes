`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KTs/PFtlBJDz9zT3fiNibi8JxPEusJzhB7seevDQfv+VPbUaXy2muYfxzf5ZsrnO
GL3wewaYtgwwB/Ius1YR2CDkKaWrndswGcb6L/XdiTyURC121BXe7zTcZYc4nlOn
F4zS0jAtVn2lQKNHukE42tFk5Zr+JMOaSJxI9OGWKp4/IOEsJAeBC4hGe8M/8e/L
DmmLPd+BAMqcGUy3qP8w+KeReeZH770XEnMVAL+CgPd4INdhsBhNj7gICWqOQ7h6
aJVVspC1XAxaAe2PdNOgnw==
`protect END_PROTECTED
