`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4pY6f90RmPZpvX8eEY5m7XKW5MMOac7Sg0vhGlmCLfddbW+c9ZRi+l7CZ+i8ljL
DvW4yN9vZHXJAdAjhXuPVtmdZcrvP+DLhlVccXyGDz7+Q5c/Genyi5ZF5k77yc0d
q8unC5EExiVBxwHPvHVLp2VpRgoHo7uQHG7Wet+/LND8ifhpNTLc/3xnwMwUCS0w
bbflsVfIV3KUcWcTwwZCnvTabfnkqRAaKk3WQOTCM1h8L8bJx+r2A7cpy+Cz1DPy
5C4KAyTBg0UEtEk6Xx8aI+e461DDeBt3FpaystfRsz24nUpaQH9nANB4fb0Owe8X
jDGdZfLWgbQ/fOCOj+sYkPfA4FXj0HMUcc7ILVHDp1re+By253ora8y0Ld0P2CfQ
yaDSoGdta8w+zwtFByJue2iZV/GcBdpvzAvzXcutcG2K2kaeOXNQtgzAlO/PtzD6
U511eXOesDvuqiQS7yDf9M/lQWY3daPceZVZKM1u5bWN1SUYyMW26WfrjPT+gPNv
Rnx8istrvI2vOMrN2aRcZPqrDlNqfNLFgjKqWiglQgAbeEew8nWTyrlzAQiUfLYG
bryGEAS+/HmyHeGDG/AaKZbiUX9n8xkCC+nCsNFEhmq5SlX0B7d16EAEwiS3Lc4X
fZvkJDv3YQXCfWPARdwdGYBFDR3EjF1xaOfsrileVT9pVMFAKDclm6OoVM1KVaVn
Zww5UibFsMXzTdggk8ZVRsCK/Cm8DnR9q6iqOgzVf9QdDOvVmKU7p62r7bwSYOXS
/qBTMHR3kJnAXWPHuUKMmF1L85QrgJ/245bDXA+j/9DCPWPC2hEm5dKckXCV2PcI
+DQ7AvWXBz8j9y2kPBjeqENCKMYpp582CLBtWpaiW81SJg8UDsDNoszKRq8SgAJm
c57MSSKi7Bhcdpn3leGwePSKpAQWW9trGNh6vUlrAus4xRhPzyfYqodAOnc4BRhB
bD1MLnWcnghWkOmdM4QlJxTIQkG22jFsA8a8NZagrKRPdYNghyPx32mmTG9uFAO1
ZFt4F8YUSo0uZJQQDjRMu7eXTVwt5YpPyLrF1C+eTPh1nRXMwnVwaQmF0CewkzcN
ahOs50vXIEGXHRo2JRLqhqJwZAkjQ5W81TBhNSXMUG/NX8pah4GmO4QtaGZkJu9F
Wj2AVZcCPFbGcd6MFzZHvO74LAMLykbMCwxvyHqNacGlHtCCZ7PvCw+xBJBCn+Oh
2BQ9rB1YA2SxR7VUOFs6JrMFh7SdMk5Z0rOOXRqUWWI=
`protect END_PROTECTED
