`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+6Xgwrk0VxDtcUtUTYSmMMUrZ8SL/A3eNiAFGqW09PCq/DiCq0pwX9yRqgjhpGH
hQoq+sJrQ4FtwzlwAmHF4dXkeXSdQLffN/1PoA2CYps8TKKz9Z3sx5ppmfMDB8cZ
DdDwsj6w+H8WQduYm5HttBcT7dnM/ub4jsTTzi3odxQtBqNUgj2A+aGk48b7kfm3
tLAdTeBE4s+1PqO1tJFtHOeqBV+Fmdo6IfOXq2C+Yruwi5HtqbVQNYLR6DT+u3gx
qmCq6o7rQkxeKpv9m6e1UEWT8sIBQ6EgTn1oLXPWERO6K4xs9bKUWqwXh9fEMeOO
yGhx+ISITk3D70nCXUHL158b8nm0aCkVqzoXEWIHpoBSxQsM8oUO1yPx5RIOOGGo
Zk1JedOTl+MZdd+cUHQkd5q6JcX0sQBwc9yGFuFEDjvfdSNvLCN6o4o5JXuGALPD
jNyGVzuw2eyboCeg6cN3wFEw43gKaCim4pZ8Uc90WcBltOxJY4qk+Cw5M/2dlasb
xPV1b8CDiorXQ3PtgSQel80CwWGI7lThf+9696yImN7oJn0JZstBHqFmnRBcvi2Y
pf40BPEVj+5s93kCnmdNwQTp9rF78KdQbrJ5q1GdIcEMSS8u7sWAaDK4BMRwBZ8p
NL0xh58BMt7YomeqCbvheLiz1OlgcFciNyD0WhL06ibCx6LlOBZYuCXsbCpo22vA
s0PJ29YVSA3KXbaBUASdXANKIOB22s/T8DhVby46YdTaDZnUAUP1uJmaPUPwL3y1
K1ZlLWLQlOve4NbI4hD207+bl2+VnT89//OtkXi1GWHnPIfhmUhj2L09nHwiOmMg
M+w3UX112pJI4dfzpfsGx7W7RK1rLf/atODCokBzDj8CmjT1xdznoMgiARNIB+Cl
U0ljOsqc2lsc7l73ZDTslCizjxyC9qInGzWF712dZT2i+Z6vMgLH9EmW6+IwEYbr
BjWW9JOvtNS11ayH+9j4cl7Pr2QNH8uQFv7sa4gvuf0PyQe12HXk2rBCfOo9b2nI
cLmyVGHPdlIV+QkRSRciDExs8BgF5kYPQVEXGD/9t9duCwcj9tLQyhiJsx5Lcae1
cy63uYX6qrqPOGlWtiG0+5Wizv0bbK2tnJegzVTjRyQYJHTL+xdowqzEn/KqNWIC
KxPXPjwI9jWgDYF9lrR4jG3ElWK0xLKAXeSo9OBIl4ggym8YEtpHdYjreZYP2eoN
PxFkzvNSE1wSyZfaRkOzdZN2SHbRItj5ogAHeEAEkSqgYiaX8U/qlFqM2ud2fDLv
kE2bF0sLwzeR1R8H/W7K+fECdwqqz3urahpscJpnK4Ce3erEA8+4EAXKHmK9JCIX
wRwRWbgPJ1dMBRE7m+CSf3hRPMRyHFhx+qsC1oHRdgg1+fevrBbrKj1sODG5bhiY
HwayEHkNUrN+SrKHoKzkMAVepLyQIQAfr7VgDrOT1X/k+FjMFAuAidJx1rirq84L
Z+iTpNf4RGERavX5KbHhMzIpf9s8LMxI4f6anpjkvWY6ShbuNzRNb4QN+ZSVNUHP
zoWu8+hOygqtdZqWaaQJ/14Zbgz6AE51UsIC53J61ht1EKF0FAS1hL3RA293GW4i
kyc8gCIOmr+gRitY3akWnGofpK2KIvl/+JHT3lBX3GTzGRbUOv9FDTxkyKPNXcSO
69XH0g74s7ZhVFymr9DWJjTSxNgShx2yJzMbovFgA53TgenlE4hsXGoPjEsHO5gk
Swe61PY10FdG82r7IPAu4+DeG1gea4QnANvpXAmFX6w+bi8uDeCBgzSr03OzcfC4
eYo1FMPuXxAW+edBAUWiGkix32IkflpiC7Son4YHykl2UEIM0IsbkwBE5tjHojMc
GEX+340mEJDpEATlALq2LWVLocV3OtEsWfx6jmttykOp31xpZLlQ/mcNPKNASemj
aQx37+79LprtxtuuqbbIEERh1UZX0V70u9NGtCq93le//ZvViYCRoDVES9FNSgsY
4idvfoFVBxPF7VrStigXkuS3+PzyRy2BkNFSvfyLSq4oIx9dzRcifN+EEpIPcwNP
9hlQb8MkmdurWwasrpWgj8aZYHnVMup6EmeTy7FRojUjKbT2nl+llnMjwkdnZFJ3
pv2HFDDsksPGm4HjAHg8m6g7jvI4kAPPwRzHdKiEkjLttFmPtVQ/w4AXAWek7BRh
/awymuZH4PIK6AqZQ73JJnHQf8JHOf1C/IIdBcp3RfcWVYYraNDZ2YwNnRqwbVhF
2ZX8mdowPuJ53tpcmg4PF2rqcvouNsvhrC0ItizNSuoSGGqeD++qMRV/Rhs46fte
fNf3L+9UAuKu8cepEvHJSdZsf5y7amnNiuK5jPzLTJMOdcCd4/GAUAN8HLNNiQ7b
PT+TtByC02b/aMiAJrSP+DKoryJzTd/awdZKiPN3ab7mJC+xCgeQJVMS1/ZFXu69
Yo/v4tJDUyVdCLaejaGHDfFpEfT9+ooehIXFc4M+QJL6DfDcJ62pbPEXDV2RlOUc
bAj5CosM51nXELRfkA19CCi4AB6WcmHEQsf42H6Y1X/ogzr2CNpL+WKkOn86RaoL
94DWVMy0lKL3OTMLf63e2FCiweDGe9+z/o0/zfiqfBihbmD2vUl/MGZIAa7i2asK
Xf8qNXxEpil0VF5ono4p8MwOH2woQ5jHrki0NMggNx1xiiGaoewwB5zNUxMM6FER
9fyyjk6Vd7G/57p6ocV/orXO5c/bhnpTWAh28FvAU0KS1D4ATi2haWA43LA9pcOR
wTPaifunGc2FdA3jXsfeDrzHZKcYHWsy/nDd2MymdENDQG0OVWwcRV4M82z+amVr
sV6tYdfeUn0aYItCa1x56CB6LXbbMhmNcxHWSr5XFwNDEK+mDDXJljQOtVLffRsp
5J5UTMoN6/ctNeDbNG/7RnWLDPyEabn8KT8B8HYlK0czEATWKNIq/geuQO+kOrPj
J7wkVXVoEtaQk1VC/lLgEOylvM25MS+54kYtPzI8Asz8h5DWhA58WWsqGVajTC/B
kE5RDPBuBIlSnt/LCXW+zhMZtXRZysqvE2/GzLyCsak3yye/tKrKRPIEVnN+I8Y7
+gqy1DlX7u2MvbCdy4wKD3zt32+BCjMdKCLqF/y4ivTap5OX69V6mqlnQh5D39Zm
VwLt19zV372PIuBx+URQklYPD3EzdahcPCA1DWkdmDyP8npmyicDLdU2gTK+wABp
enxyWnBsmHnw9K1AtQpjVWL4kGyfolig9pmrDsKyIRAlHanDJHf9svXQ0IPuTlL7
AHRfoLq5XGaB/Q3qnIKVMn0BUeiq9QqJXawuXZ28V1/GdYS33yzzbk2LsemZwDVA
KYy6MmbIDSrp6sCZMe75guGdrgaGQOXnVIvxxIqruyNlN2hs1VqMS30SMuoSkLcr
jo33G7S7gv6OwIwASxcJzbp0jNL9/sY29G4WnvflV/lrPSMhUOj2PTjPdozHd9+P
yeHTMrqnE7y6y98d4hImEy2xq3BnkG7KyZF9Npy35KtFY0McHPWwK8N1C++poRQ4
b2FOsCFaYtwTFx6/MVbOorXNor7+RlVW7JKdBkbXBuSKC4QEZBkPQB6aeX/EOm+t
p8cs3M8UOY4qeUSj+01hnemwukuFx+RtNNE1DuJZmThkWhC4LfPCLKAutVZWQaUA
7HZo4GlsUFZ25N5z+BuKTgEf6uQHd84cWv7VyMs+36axPtPQjRTCYie5IXh1zl6Z
Z5CM+JKafMVO0M4EPSP9eXziRl/mbIWFv7b3fyr83/zjPlu4gFp6CzApLZkRBH8w
ElYXr5/zB6/lt0znP1sBLMeigyEuQXclkxDkuPFK6k0Qp/lfRsIBsWXMzmI5KfVl
kz8nnNeUnE10Bon1Odaecax8hyK/U2kZlTJRG6sBKvn9ByYmKfnETbNLQiuvkmDD
0e8VomeO+RBySWq8mTVOY2mrAt/LjARct5k+yxLCXEZg3SO0yw0g1R+SIOoXZZvP
6J6n28IbkKWqTFBzI/UYC5hcNNWAP52uC6GTSNVFO11qXkaxWwo/oaHdETfY3hVH
T4LWlGNb8V5YGrOnxhkIKjAcyyJmQJemV6GBVHxNelNvAzjIHxOkkP5KLIyPftUB
DhF4lQVryGurSdrTvmjKIAmIN+7xnP/DOG6fStZHIv0wLbWhJGkLIBGrW5emmY4b
2cL35FO8Q3j8YY7ovxghNZ2WASM0wYu/n8RKCoPJC4s06Q4SuHjlD7M5luXevLQx
JGt9zsGJnO9uQWHKNCncSAD2gNmlCxecL3lt5Q4OYEGrBOZ40EoHQ+tmzfZJzz7u
OWzzXNZGbpHRgOidosla6a9gdDY5a3IdY94veOkxcyio12S5D5gC708lXmhiKqSD
DQjg76WIBC0gpZq7VrUgMqTkUHyFQKHGgYAYCvMDLLoUAcVBMUf6wd78AXW9jtTr
cjgTXNqZqGdlFVWAuZhMYOEbOrq2iNXK7Cl+6FqbdPxgyirQw3Rw1XSUpNwsLnGH
SxYWZjoOY7UbhGhUdayVQqAizO0sW3pKLVRwj6gXiWo/rmWsjvm9rYfaKW8zIchN
BQwehQJ8Ek/gD48aPaVaPb48RTnxv/ETQ2HX9OZTA24jnbF/vOh+5rcs5s8CtPRr
X2HVgp70W3DsEpps8WR/qyLSh8VgC34tUpVHkLUTCjGtQOqAXOgnSninNdsULdhf
KsY0psIZj/EqWJ3LNTIN62xPoPDEXfsWMfDLdJzcUQGQQaYAf3fccjzzt2dX0Pnx
ReG3eCmvLgmJAPgbAuHdTr5xjoGdiew8/7fI+lcTAvy3tdwOWq0/a6UNRpDc1uLz
TD7S5SEe8UsPXBe7nd1n/A==
`protect END_PROTECTED
