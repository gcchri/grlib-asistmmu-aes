`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kO6BDjAnejMAus1d+IaqFUsm29D/kZ/hbNgQy15GLhO2DbTOk2oaTWdFaLmAgZMO
MC16TdzBpsNRJIiee/AbsYYiZdXFQPdIEgT117kMZCYhlBHgBYadG+mNPCwlbJYC
5z7utN7s0Mziyz0p1aF7TJycBvENElqatxVgAucivseCNot7j/PTHJ1gLd4mGvPG
1+tbapz2SHA0XKXEv59eq/x+Vte0YRcEd3TaeAUGNd/4u5xo84FH4IVCgg80NEGk
Rltk/9azJe6qEnjHEbFdLlm8q4leXH5zLM0j0eYjmgdpl325mMC0uuh+RmMggSgY
zSJZU9fn94tVXW7VpucWsl7Y1JXcm3ekbfpf0ZJA9NeLHvlfa9bKGN4T8DY76OYy
uF/lfd3jTda49AyOvoVNuBmkHrxHIdBbuZczoBCwTmp+IIPAoVcdC1yJKnPwnRUm
9cF7g7dKXhg47WmMjrHkf/bWGXJMlvo75DDhj5Dff8v64LUSuM0UMDJ/oJo6H+i6
SKBtCSnlHr+VDK86bOX+JXqZKgORew7Gnuu6UUBf575ScelKnS0QzEAZludDRVXN
OLBvbLiLp4vT8KM1mlusHpSf/a3/+l9N42LidPpeJvLbSLG+nAw+jnipZCSJgv6I
JjSElAGJYtbWHLDN+7we06vNd2kAyxbAegB4QR7DqCOiz9kyhD/9EVnTluLVaR0k
nS8tLKJoEASO9Fq6TQLF1wapMyPAGRpGh9L+Xl2D85gkALIVWv39JQlZ9VgKJ1Vi
rq+8nsW4UAZWPYQ3BWXz8l1vMd5L2xSOJilTXUeFy3akaT6Y+teihWwxgXsULjCp
wDzModOn13ct9SwU+x90dyYDCUlC+V9dKF04111jgQtTs//qtUIEqZJ/crTlhoNs
0iexIugyTOd0cjD9IygcwYPNcb5v9fMdD2cLD2+pBBPm84dfcd9YU7dLn+nRcm6z
T9Ttt1nNg1fHr1/btSfwCU0ecJtdGiQQkfGSUcSa1+WXYdwx1On9t/8h+/eKMxjI
gqY7+xfseGsm84H08vkXng==
`protect END_PROTECTED
