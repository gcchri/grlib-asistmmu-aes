`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1eU5GyQVx6zC0F7ciBHT9nocVOGstIVgGKyhVlj5E75LytPoXx7YTan3foSTVDL6
DYR9/Aade/9zqZ4xNNeI2oZGtwIX64p+PPg4ZrwmBgW2A90tntpefIbrV+rtSGds
se6th3XoCr4HmIuuUiJcmJOXAC9wM8r9HLj47dhNaeRn5HhnQjhhdlQEYdz691gI
5x+LDTQh2DqEwLmQVg25C/VPw0t+MX3TbY6/MQIKFp81UtkfdqfS78QFgbFpqzG2
eFgZWfzl1iwvnETBdi+twAM8FUp7zBED+u6crp1pYZ6faFr1nHWgPt27AnaoyEg/
t1v8xgZiwjxEqtvcGH946hwjD1BGxBoj5qwexUcyuiysqE6+4L63qxcss7TYxMC2
nrKv/DtJpqKt8WhZd+zBcw==
`protect END_PROTECTED
