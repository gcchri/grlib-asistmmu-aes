`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YnSoUMOqp+hFGQGqdtnfxXlRk5Hv4nMRDMsc6b2S4kJ6s4WykaLlx5iArET8yjdl
FMX7qsA6kW8Ffv+Ba56jKmNr08NiWM/KkwqTpHO7sGQ6/1e2apxj478Wm9A4MgO5
yQMKN5rxN8qcFvvjGC9Hc+fGDY4c2DsHBgUc9MrHNcJeePWMr3feg8hV7XjU7T7+
1GOJKRNu8WqHuflyEiIyHA+R24NUHnGaR4uVeS36JrBThTH0P45nbexFZrnB+2kM
LGpE6Ut9h0iB6QnOjs1PJjvKPP4tp5q/ZIR/LAA7cGmcyY6f7h7/kcbvqrlqgaUl
1SeCA6k7TotCA/jG7d5Z6JJF55PIb0c/PIHoaB6Y9KpJ+6imvVzRienQacAxLHWB
6mfLMEdjkfInB+iM7S7n/n2pMLXqUdDwc9ZwkxYVyWgTYxKgrfWhgeV3yMm31Lt8
vJgOVV0dLNdnUDxrFgh/33vjQiCvJ1muJfgm0MdXjIuH/1FjDlTA7Dlfwauq9VMp
/2DoRqo0fHx+JVUn70ZRJtF7Bbrc89FNfaFx4JZgHlPTTlkqtNRrZ7k+91ENxgxD
Nro6fcfAXqi1/BeTQKYRwA/CO5EKGJmXX5HnCFHooOQpKYfcJPZhH5E8YW8njFlt
lAgCEbz0e8ZYLpltmIgOt+VR8R+9Iit6/+QWULoDG9i1MmYJ8Gn2+L2i1Ecrt8bR
+YemqsJXTTLuAgRLTl2WrA==
`protect END_PROTECTED
