`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
il5cZTQlQdqMYEq8N82f47vrYSgVIJGsdcNAT2xONeqzFIBQtPJBJlj398ibI8XB
Qz9AgL1sMTMcLoTGRYXxaQpyZQiOoJRRlKk2DOvQHQrsSXFKIP1wgeFvYn3xYJy/
JptNMlQdjmVrUaVAwzAYFw78nEmlCOpceAtGox/agNyo2qZAL89o6zUWrUWBbR8G
0bTG0VsFNdH7SZwqM58qUmIaEHUK07vVREiGCp3/rX1MuysdxZuCZKI99S5XLqhd
5XKZ9i68/4hiwiGclJ8SJvqCf8cFgHHmCVRhgkZXxIkSHk2lZIeWKtRTrXrCNZmp
jAEv7fXcGomf61U7+JcMkeElKDbJ2YWx2xli3U0sj9qP38nfuKoPCLPreQN5pCH1
Tr+Lv0qQPreiTCMzlYGQERYE8v4LuxCbmuhRek9MTwGhEp2dTVg2zEsdcJh+GpQX
KiSvYLC5/R5Se1IQPeq6mYTI1WC1+JVlIh3WFhN2lg4Z3RDChG70wvTvfjddQ1Ta
WjeUSfwVU5m1S3HEERq/O1+GvuV2SslB9Z4bslrAJuhWYz2ZdLwlwQoDS2YpUKx0
Atjg7bA5+uGgB6Pu3xEE1zrR4If5XOzbBLyG7nUOAmMdMQnTqCitG48/B2hZwRjY
Qm98F9qBPjrbV5F0TIGV+20eJ+pc00c8SrmxcTtwM50NgvlIGDUB5og4LFTA/JEb
U0CDlJVM1ty08MXJquZYtQ==
`protect END_PROTECTED
