`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NmNkUXr9fa6q8a+fUvs6BGQIvhr70CgaP5KSEUAoeLy3XEXWof1mMLv6Oighf0m3
Bm9h2G1PIfW2GzY7RkvKrz/Cxcr8u452u+8tzPj1nN8JDj6MjQ2uv/9D/6DI7zgn
21jYOxMS31Y3uC/9mPc2UjwwsI2o0lAqKgpwx4snzJqVjf8VXyVm5RT/rxFq/wOa
pkrGF3XuPZ56+3evdxToq5Px/r48SulBIwpxWBOKbOvhJF8E5BkXNVPMf00g6uY0
7OOERosCLJOv7EU4jEE0bqO4J7LGyt+DQEyi+jV9us8lIbaJIZaprNlCdhwa7NvN
WK74d2xAKLKn35S2vP/u2WxWNI8aGW5Co4o0Dt0/jUu4RSmiunm3xjYLaMrYoc7t
z6bDruUrzZSOh+h/c6ekh+s3hZf9bHyXKDHJhb/mg8lqhftE3xboaTkGtBfllAfo
uvvZpK+2BW7Z1uFPx19bbzzRtBlPiENYNdnVfeVhfV3iuL0IEziRMgAHR3V1oQqX
T0aBILYnzOKazwUS7WHFotjqruoCjfBy/G/VgTDntunkiiD41YrwO3bescN4uG/0
aJyLfdmkK+QPT1KjMwlwv3q+zPG1QD3+Fh7fnIo+C48T/hLTrPzgNPLcMvi858A1
JePBzl02YJiODMOG7y6SKzVcdDOE5Kz80XlOMXn7aPVBaP3x+Kir3Q88RVBMypMi
uq0W+5Ijiur9fHUUpzgcEtNahxtSQmCDHmo6W/WLKquwaoL2jg2STC9xWxEDBHaF
Jb+EuoPBcUkl9q+uiQLWQvxxSwebJbi7XlC7lQzFiNNvPszPOhHFDvCh0MKWqvX0
FyxpkRbtPZGNs/mA4nFGejPdwqab+hSJnfl1DGiWWvuVdq9q/5xp4g7ncG1g7CzB
TWk8POq4Lahzk5qrAOnURv3EFOAhh8Ra+6/2RgI3fT4oe4SPdVACQSgXeRTvNiZT
+VTISjhSDiO4E4mr0BV6MFzxAqMw9jJ0gSozceklT5ZwUQh8CAUGTZpof8b1gT0/
pR6LZtFbkHdibASEjOXqjXeuDiuEtDr48y/Zp5RHLKqvN52A9AYlTYJ0ra7xxEoS
6cHK1NzDYrcg37awMv4sh5izzqzJNUhHvDUjCoysFDs5jKY3YUrV72CWubo6jD9J
5QQDPVoAbe8bctNfzs6l7KgmAPkL6X5rb+z8m0X9ysUP9kscN/NNdn5vH1QhseSS
AAwZWYnNWUbb4GXTBaowcn22UoOxowLYXOF3k7sQSBDd/GG6vneZAGWpQC1IAwCJ
bfoOWsz2skxBthbjSoCZRSxpi4v2LUbT+WSYyOghQ562jgkYt2JK6wcSATvf8kzt
nEgJ5/jdgsVZ+LCW74FkacMus1TjrVPFrhIEtK3y7LFk31rXgoubA2qz+Gg2uCAC
z2bR3cXUYjpdROyLvARmE+lKDu86nAqHZhrUcNeBTKOMTyCXtteWkb6YOaluNsHU
7pA5Zb/VqYdZJbZgZHRUVDs8HCklhMp3xiNfq6enalni+NuOK41WNEFPWp8EzyXP
v3c63HMoGVz4kCgp115DLh4p+wG83Lpqol1/GTaDG+EuRJ+du1+F4LanDKwKHb1d
LePVtrj+jcOCtjQBNH3BAuEp9KVhMw89DwxLh6HJzgnksTVETpYhuNO4+7lwmwG1
ffuGaIAg0e3jxPtbMmmQBM14VeFFhk3jUdyRGBMegZWdcaXhDA6+qkMA1ys3PX+g
ADBFAnJ22p2JjP9tkcwX+DMbCfeGisRebdORd5r3BX30/yunUKhEk7Xd6+rm9aDT
Q3QYzqaK982aSCB/EvGJh98pntyW852ZWkNfDCLbhX07Qx1qhpJvrUCG5ZwzhUQs
sFPK4E6RUYyc9UDXsu9B/2nj0iqeQMHPB8HYB+xBDeXuq+iCR2vBnRe/0mOTwRrn
vPpGe9N/GymQjHHtMtIBv+c86Ul6ifYhjhRSMPk3D4JBZ6lta/FcoPltQe0C1Q7i
NHLRNSgqrveg/u9jeJeMktB8XCm0C/CH4ScOmrNKGE03p0IgE2rgd1UmhW3BVo2I
4xiN3KncSKjhbSzFYarIO+NFDnmUjk+38JB4CxqNchunSqW+epEm136biFcgHBmx
Yxm+/p4bjpxo4Lzi2MIb+ncsevZpHGnrmshuz5c8tmKCSefBiriM8tmqMJEePSPn
w8vXAYWgOtjLpsANC/L3/r2m3w4eVBbRVuewg6FrrH0I9nwrPPtpm3VZBNIJxkoA
QzPuvwtnGX1AQKa19Z0gh2rkj0N9/rSZWlrgGXX9MnPUR+npQgk6Zz4HRBJ4Uif8
YSyEsVrEvHzlzLv4ofxg5xckQ40QwPOudLSy1IXa8ev8BJvGnoQidzImK+6XvYeH
muxxTYL3csqAcB7OOkTcAiNtlPzaY+HuUT6mGk9lUhI4KtwvtzeYD5oH8JPVGK+z
yLWLlLJG67cYQtYbx3+WpuNgnbaiANvbEqd/iPzQVF+DOCw5to1iZwXRBcpdTSeh
WaqA0gPy6VWgIfVBvxX/+Q8mZrpj43To+eWJSqHdxDmLhDu2p4Ybiy7veAT35tS9
BJKYPAYkQEW1r8rlywy5xqXnkH2mr0e3xeeopaf31jOPOX9Va2myqcbhrp7KhO5c
`protect END_PROTECTED
