`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufNvddtxs6qaTFJzf9Q6gDbjwSsEIQPRN2Pt92dRqrcxKFQrEO/f+oD10/xbHav3
SMwVvNM0Abv6UkwnrDHHpyJrPm5YxwsAj7u2k/mMUL4cEfoPdffYnYRd4k9HUiHd
prJGKNg6BXrqkk5X+XLMZ7GXKdcUb3l2BvRUStfbGPx+1Ew9QtYNWp39+Gs+Db7D
MWO8XBu/yTuE2FN5TX5nXfhYwE4F+a32HFKcOMtg7qFFjo/197e48BSyLYZemTSC
4J1kkrxJyxMmiDk3e11Moxqi5oE64d0P/QwWTy8QJYjYao0J3zYliFxb/C0SciSP
nrlZxXSgKRVqNFkz1S2BYvvnPFANgUnQzmY2/2piDRJF5Ru/2a7r+dUlv88+qzXA
lb1Fcu1QGR9jFnsKR3ycblLWr032lAqZw+IL1k/nNNn17CpY3ucODgv2nIwlbFbQ
iqWmklKzlRbGDuP8fXiXNgbv0ko0drP6jP3daogqLURS4fCG4DtM1QWr37aHojVE
94kAXlZfrxvlwaYF7JfuCMTGgEPlH7Ig8J9UtrfH3L0HuectE5dBUQvy/GhLAr60
FyYT0rckX8PPjkqf4CNLhrq4ccOBtD6qHWQZTE75p/MfkjqDd4ek7V8AZBCYQccQ
3L6ATEPUOTQhXbE44/RC8YDq8UOXYOUOD0qwLbZaRbpLAZsMywHJcRMjfy05YC95
tE8YrVPGnKGbPk4PmKYwhdkv3g0/MgnqvqvEKC4vSYt9hoBx39OF9It9oMoLsNSX
MZfJk5lzVKHY0xdU4xPVTA==
`protect END_PROTECTED
