`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DbRrxQhwXm0kH32RH2DExNzDGNyFHyfzXOMDIr8HXKo14tzxnQVAw1nhNZdCuAQ3
UraVgE+98Y936zIIG0Aon+qKIZVBcMz6MPlgo2NKRxNEs4P6KUW14loXY6Go0Kau
BHQUo9QeyZM2VhSa/daNZ/3RPXuhGgy0Fs7mInC8+IpC8m5nWCD1nRk+xkP4SqmD
cdMxVBuiCry3z/vd8i6llkwQG94YtJvpvWiagA1y1K1dLW/B+aSlt3ntDeiF0+QG
mKG6R2Tj0/3BXnciREc5Uvvknxq0Z/wZ4+p/S1rtdSpHmyupbWqgtfgkrM5Dgipz
iGYdn629CfB06SSodNUYm2GuwTYjYhsiVh2oPtbw7rptMPn1GCng6P7zC/2FGsWl
YiYB20Ughy+kiInJHxupe3bM3AV3u8CwBfu7TxRgzoRhVSZ/z2rsf9UEuiAKSQFU
SWe5aUIJ7Oy38CAXnzhhi+O02ErBTLvus8lLivPC4pI7BiZs5WCjgrTGP8Q9vzFi
yovBghUmLkPgKDfhQyZxfvTS9YIpBSg5ksfeLFIxtz8lG6pzRs7ET3w0DstA08By
0gJR5p4Lzv6itabUgUVMGZHUWOwnwnDcEudRi1AUt4ifaQ3rK1o/886/8+8C4Cxe
ufcKGog/JZbCXTt9pXgghQ==
`protect END_PROTECTED
