`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KYdS0SyvJczxxMTRCgHXMKHtTgNWRdMJNeavqNZHS5BISQ8Ed53svQstyg4OKpGL
u7HPOfx6hPFHI2QEhpKTJo+TqON5iVH2+F67rH33nvE73s1eqpalA70g1xb3rvO1
YQI74jwnEpxpYK4rI4LrImAj5dm/uy8oLwsnsXypDXIkm1SmtjsvRNd+IPGo3ozY
Z43u5i/m5LCN2pUXC73p8yJsVi7Qp3i0Mo5AF3ivo7ASDufOWV5TqgxMEr/9Nyuj
uIIpUK0g7/U8OJQeNWOvM+AEpfIthSNAWDnoJRfLoUPDUpvwE29hp+jmFotgAnBT
5WN4RUSaHd/9xXKVhr3zu9gihifOP3bx6LwmD4HDxjScQW6WBxMw5tEBzn9qQeTY
0UxqcppFPzgsuKLHEdg/hoQMTvAWVE21zMTDXqZ10bEPZZSfiuTHVYC8CZhitIU+
ql745iEGnZpMkvEttZrhZEuC716rxHZr7o3ZwAuVqh2BmWAGLgt4JqXj0uGpSKjm
`protect END_PROTECTED
