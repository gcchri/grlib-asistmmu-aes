`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vvnFwpbbWH8VaVRACHMoEHP7g1CHpt1OGxqDfDono8nrOE1wAiRu9Q21co5YYrI7
B1/ujprYeNLowk8U4ZwxsUo/Gy4vYarS5kKF5nNgss1WXJvZn06HIPHCHq3OXvzR
Od//5iY/q7TJIQtRMAYMgVV6NXKg7KCKIIxrVNG/q8eg5Ynlexdvj3tYC596mv5l
oKUrZuTCFqnSWbqpoIJ9Jj1BW19Zg4qz6RRyWWjQ2XKxKQRj+j7G0m4iwRu+7w/H
rHrZxQytD3PswN9bxZYl3lwCOT3+PJzuS0f6qTLgocKiDSYz34N12r6mM73xFja9
dnHQy6+Yjcuhhlx61QVHpvkLqUV+ohe8KU0vY1oNIFcpdYWtkOk1MSA9g3fmbrl9
ip1oGeQ86VejQw//R4MGGKK5wIGEZeMeOlqlANtGn/y21rH3Fa5GP7bYii021g29
Op+Qk9z3HbKkGOhKxZcEj7BR91D87wEb3v7i7OPysP8PiLbItzadNJrN/WPw9Zb6
hLjDAdWtzsAtCayp/MRIbxb28R/i/dL7ND5BJrC0+z816uZlAxOmDZhUKXZ97YkZ
jEkCt2nQuNV5n6fFUL/ZXjqHrvSssox5VcT1D8OCOkhHFLYLXFtLitXeCD9rxRtB
A6NJDV6g+3Z/ibuyUWb3/Q==
`protect END_PROTECTED
