`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGOekaqGshADhkjNmNNuCDs1ygeW23y2zGh8rT5/E18admvd/F+CjX0YpMzO6GPg
XackFZfN3rxrpMAs0jHiOd87p0lmdricB7S7k6sIOQkn0fq1JIWCP56t60ixPo+n
XoJ7tdH/jN0irlE4QBmhjry1fHHkP404AoC5SnA30xNE4N+HTrulbVj1baXPKBce
MNhVvl1P6ZVfnzUiCJMabsUtM+G0xgw7zI9CY1c36oApd9A2Tee55E0nruO615lN
U7eKjfq/nSWBOSQFm228d8zc+SxyPze8/u1dvPK0X3/c0W6u80OK6K1Gl650VkP5
d26N5xETnMsAdgJqZ/WfhC4RAKRLxKTc5kLPq28cRztrLaylTSD0sfbtHgxD/wPF
kQaMDTWY/FA3R7uM+TsPzMR8b0VOtet3dxQB9BMmcw/A7rHYETDf8QgNPUss+PVN
Tw7GxoZmRBfeyO+hKWrcaKjOTBbkfVpngjeLJ6tZsbBzeo9t6yzAeKU3wXGl9CGI
XP7vdxL/mnVilW71JWQV4YdJQhwBovRl2PBAugMPiTY=
`protect END_PROTECTED
