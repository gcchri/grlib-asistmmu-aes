`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4nkQ50DBuLssuVgq5tL+3v+L9IVV0ovTO436pcIzJtnpd2hiaBz6qiOrM7I7XYff
q/MtOAHwJEeFoSWTqF2Ur+OVqhCm5ugQWAE5T5K5nnarZ/68AHN4JMdNonqcv4MQ
+PhJIqxy3galW8+OkVkPkGXNI6hCFoSuNja53HbCY1TZLxc3bUDHE9nq1lvSmeb8
OUDjX++2+VC/ySLSRGs/lJB/sWihMMXO2NxPcq0oab+uB8zwZRYbpPHUn3YJKuqW
k3IggA2kCRB2drbhUffI1l/ORgzyGyCMzgc9AYXL7hfY3DdBjsYKvHsju0Gr+4h8
0LWw0qai64FyKEX2DabkXTUfP7DEPVrzm8FQOaqsmIuDTPJCGmGnyam2XSgeh7Rg
9gK7Q1rt4YW6wrJBrtfhbY9JaebtKpiF1ToRpOSG7Bcket/H7cX4oVlY7MWnBdMK
D2kbxmeuojq7ZxGOvhgtT357KINK485qRsMDgWYYdePw25rOHngAfOq0HgVO4vno
aoBDCmF9q9lZyy3mJT5762xbr/bIzpyQauMBDgGeL6+Y893IYwLR49Ri7/VvN2K8
20UnBCUfclQrsFp7XKFkTZDy8puVcofdBHxJKEloHkhEiXLtxg4nIseeRNYcExXp
t/VrnmN4W7MUnTtWxl+Vge40X5IkTJn0umajfhB5MzhKJN0F7sac3eeiIMdngD8j
6A6iJwvj1KqdYPHSddhTHZocHTxvOO7D7VbM/l1G/wtWr80WYOvkOXetfup4OlA2
nKH1kYeP0nDm8dH2zBDodql9JgGlkx4vHV5xZibo8qeMRGnIH1xYt9LuZQD7JnXQ
kxh85LUF0GWWn8ooLL0T/SqIiOpN1F58j0vi7M/eEK2DGJT3EAiZ8OAZpav9HbSf
gJeQZvtwlRAs/xLgwtMVpfbQOV28pL5BJyizH2LR+HpQkVojNs3AajAKqbmXoEBR
afljmtr/y99ykQ4jDs/rafwvbdg+jMzU4kGbwbFASaG8kDJ+fFpaQ48Oeh8jsrQ1
ngbw6QNSzjTUBUgKGxApARyMBgEi3sS3P+VWlIprOe+UR1i12+rswzLybmmkgbkV
kqqsqcP6l31owZagJwBho2AM2mTXBoN2fF3ScpGVu3ao0yOn/qADfkmrmI7rsoBm
jkrqdaiWJibWbDd5BL0oHE6vFTb4HBUby1TlYU9DHhwRj35vURel7pR3puX+E2DL
IU9Xc/idogNEPWzCf7Kq4TE5OCvpw4HuTk47Q1Sfb+vLESHZQDxY5bqmKBXZL4z7
B8uhaHIGWbtt2qNLFoi9R+Xp2254tfrMWY0EOnHrnuiBrt2Cuy9hHJreURoS65Bn
24SeM8Mm4WvdzfLM3FcvgreULdkIsH/TkKyQZFNq5jCm/2toB39mr/2bCvs5icmO
3GYhnh0A69lz2AWjCgGIlUfWaYsFkL9Mm1MBJEnv6r5sIw/ybWIG8oahlQJeJT1s
3Tl7V2cN33h8nr+05t88eXpZl5Lvn3z52DNvF5vy51LlBJCL4leVrLB/3ME55nS+
YJMtHIjXJpqWZoWuDXUaHe7873H8F5EUN2SvjXeL58WpkwKP5pU9qqS268LiSXIL
kEHjaqm65Gpw6pBD7QM7tTS6+bLOMdXnzTcaxmb7h6MRTj1MMuRfbNjaB3fF45gj
jr9un0arMkMLMZrPO/11Nn/+NwDGtJiXlgu1mF4XDs5r9ZikOYjTol/iX8FP4Ij1
oF4P56buDuHCzdk6NLiTS5WNAB0CpXDYK5XbP3SierCqT/sTICAuFUyevMGesyb/
8P1OKxYAlnNYtipIW1eFmtDGWVVB4+9IvPVNj5W6mwHxICKUUz1xZn1jd64Rb0Ou
SxsNjzHx9o7gMZyfUnjuJ9WqfTIE2YifhEkfGzxO5y2LFRUkSOjvBT94sbXrY6g9
5am4L0V6g17pH6k2zvEJ0zww9a3BXqZU9lrjI6SbAVCkDwNbjx7f/rEUZkBF0mTF
/YylKLuxXSnqAeV2RDrhdnRBEbYHEfLg7y5vGbQcKz2XsqdTEE3NeqSgoEm1HNuP
wHgojXdUj3yZF7rrkSyk+bVrzcVx6uMJAUAGuqnAG3tppCKqmh91OHwhi+H8kj7M
9/SUET/k3iuH0uIMQKOPMhX8S9RXPP/A8HF4jNeqzWMu8/Snw5TvH5IVdGm49ihw
1wknYamTVowbduV+5CEe7pHJjK6+Uwm04czfl9GSH3611OaeVf4c4GEFJiPP0/xv
WHN7PX+fvXwF3NAjpb0E8fLYyN76LNmgOFezLa7KD5w4AvbDqWs9vJ/wSPdQl8t/
Tg4n2zCBEG8qAOraPK33n6O4ML1YAidWbVgpYHV/mD83VK+XCoCUtNVpZVe73Fts
tE6OVzreLp1Z4CYrrsa62P+F2wCLXC+Wr1jiTaDigy7NJ/voBwYB0KXtfvfWliHo
0bOF8l1WfzwxD4we85BQmIr67EgJ4gkTBy5ssmqtcmsL0imk1xQdlDtF3IShEls+
1dl0jIEysv5t/q/KMST7tbma+Mz2SpHX6bY10wYIRVSxxtLpD4srwVOInw34du9R
zNrxDeraRKgcSeeyscdH9yglXvxfcys6qMyp12+g1tdTUTp5bUc7VA2vNpB8y+ji
kkdNdX6/xShKAnNJGCKW7w==
`protect END_PROTECTED
