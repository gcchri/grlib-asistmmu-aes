`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+6g122W3WT3PTRFwg5fpPfsCh+WcPz/Fv95XkzHaPpTps7noaHYPJYSUSzBqH4+
KzB50fvTpeBiomNqwryZrvdtLXd09UsbSNPm0qhH1AgjSyGB6V62jiXk2K0wM/4U
bE2eORJBRB7rnvMDItJH+t/iyygWIDe66TenPHHsdNuP5usqPxye1WLYwt7eaY2b
u/Z4XecjDxd//we0HyItXlMKa7HpRvPyDORIuxXQdasqcQA6J6mp4iwMF4khtKFO
8n3thiOAHLCLEevvr2zrnqyyjCBi+Gr/tP2z/nZxCKE=
`protect END_PROTECTED
