`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j3HecqjLSE9cjXJU3w2tS6ieW2m8JkSQ6zf5cIuF6o+8fOKsqXLeiacPdrRapJoh
3hl+zSNQ/SO943aNePXsFlCI1Djhj9qZxBkFFEgSThlRhHRhUz9BtjCHnU8fd7k5
UWJ36RsV+n5umwPbomzt97KtRPMJFUEreDhTppz2PV9laZiOQOy2JSWU3zFf4dBm
+yapYhNp9Tj0sUWkj6BBBkvb+Cmz35Asp1LufmBDeN0k2U+vDkBpDvoob9XyC0gh
6Wzm3UqK2dRWyd0nE5hHowfpY6JfKNix5SJQUG2NpaSxR8pFqOJniXux6h/HveAT
3gGpNasHaE8eC8C7aGfFA699yrS/T4LLhlAE+ue38lLOI+CfBStUSyKYNM+bycE+
`protect END_PROTECTED
