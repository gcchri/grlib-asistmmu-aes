`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iKyE3hZfSyTiJPJA6vtdBtAMnpD1Sz+ePtQzFoQCSBiyfh3SjKkXOpej9PAwzNqf
sEQHiLwtQpHKdsGewpvZIGBQCMeR6rMgxUv4foZlqerhY8VjLCK92g9SXQd+J+GU
MzhVrXiQAI/GTP3UE2+vmtxRi5lY5UyUJp7aMJtSYP/uTHn1IK4aqia3VSDlx462
qh2wd5V3exWTLkkjnEgNywzmEMoFqCNkAKKsNrX3Flv/IAApm5S7fMato12GbiJm
4HCp+w+Lu16XC9v70GzuGPo7YIxP65stSC8fsRUidpL7igFsdSv7JbknhSBJNcJ+
Hiz7++63qjcGYsWQPs/Q8GSJ0+6xVR5uVNSsCgKqxTKXrJhXMlDJiMozxisEl959
YZNcHRrHRHh7qGsgu8P9nNahDRXw5zwzFW0LsOEmN/v0sbMSJlWXT6L/cfJwpXnC
EkL0EUhuOqV9LQUJZI839/tfuMFvZGDWJeFFMYDk2cZbgOfg+zzEQW8Wiro1qCqS
3sEDbjDB+pLqgnG9+2tmIGO6m8LxeuDTw5DOtH8BNcTNQYzTgirZ1KXpz3g5FBtE
yvYyLZLGjb7C5AlMQC1wOGLn0TmWEcHHfnyRe8k3Hmmrs7Js3+xVnAfUCu1+09us
oJPcRj8O1qnmLm90L3YSRe+UqF9l+9VGkXnqvgIVH1ZvLRxWZFxMkF0aaccRqmgR
bzcdZjzmbaQDDFuuXv0V2xA3tbF+WJJbXN2G3giQi9s0iNM2XAnX+pAi+kCviNDf
9l55mzNlAPNMK3YZsGRHKMFvCI+DjV2iOQ/zxovXUuPavxKIQtsUF8K+w15Ztz95
RWlaidaVhA4mUE/fi5ZI1xj2gkBzlVRhQyGB/QwvYPds/JHis0LvWFp/NpzrL1dZ
Dpq1PiSAvPborwOpefNo0qzKuA3ld86dJeHBoOyFcnL0fV5nViCfXNExzEmLtHpH
fZlahdl2o618fOckguTNNRpC0/aG4Lt/ozE39t9V1E/GlShbkHbpR8rVukP6sWNm
XS/4ExF9p2FK8yMPS1McEK5usstSmEnUixEZHFyuTim2QbDOk+qZJu8a8PxaA1EY
ooX0UOxhJidNXQYQ4fiA59f9Y4DoAw+PRsvXbY+Az7YMnDG71AmW6tpW8GiXJp36
BMqIgpNPsT0kHuDVmVNr6MeMiNql9bGLLNHoW3H76COrruYJETKbeIr0IqgY7Sys
C8DBEAB0/rg+pUK9wYuJ1SD8gykDYcdok6HnLh9xgunEyuYWxmlGMF0YY0LNgCg4
chzizsFO47K+531uZ/opfpis/q4isPGoE2dl1A73VdpHTJeLMqFWErllOmOgeSrj
TKJk88X+uUAT++PLfyfPYqROx2DMrIpbRQV4M8yPwEAgEc3AeX7ySMSxUuQtWMF8
jXNOXcQ03mUvyBgVl8Wd/9HcdsUTympiOj07TS1BxtzzrqDLYGkjtR6MkxvXM53h
c06O5EkFt/FzAZ4OEKYEdGZsuCaFwMJ6MVIJiK+yMHU/qnkkIsWGQmvDVX7ZzDwi
mk6pBxa+68lI/EVs777IRYfwGMaRE7lFFRLd8f9YZ4HuBGGHncQRHE0l9p4QECTI
39yGo+eyVJ32dY9/qTk6G01ci54eAhW3TtAUIOrVjC20EurFze0Y7Q4xgdjOK903
67Ck1G37oOsQbmaEmfD6ez/8EsPNppLQpkAPNaS3Ap1MWNbbk30wgJfhWY8+fQEI
23GLxJEgrEfmaegqn6U3JY9BVRzSYe/Xi+Fb0kcL3s8mUs3kYuVxaSlwEM1zWG7R
D80fHX9mtis7j0nOm/sWJDsjG17VUtqlt84rsIGQ9fUQOuXqpLTpP88z46tPirjD
0PPpCEwQGIxKEa9KdJEPkkfzHunaCyEpwRN5geXrxBBumTilwCDu5Dvfn8WFpXqP
Wx09Ub1lUmR8qKSY0lZ0Mm1D99QfqRcnvi2Tu3jFt+WbaFbWe8CRJuyGWjivdmL8
r14NPByirk4f9GBicTTXbFIVr+QxK7vy9M2e6kr4SQj1YDHDX+8HO0vT46Dyo+XQ
Bj8fYSqkeVhv9SdC0tAtZp1sJTtdKiObGxxfeMdp6Zv9J4g12CxioX9lgdih86il
Lr2HhKEhb4c21zPz+NsDwx/SVgQljd6YKuIxhrcaffJMKrY1HWvWY2F/f74YmZiJ
sFxqdaqtvZ8gzXBismGDxO3yx1TF14b5nCViOdE+7akOUHrcgfuuGuizHEEbsDi0
ppjzBCYZoQV+YdOc3R9r5YfNC8s6Gyw68mHBtEjSbBHlkqjFlRjZ292OF53lokv7
DBbKBqO2LHp6BxOMMQE/2+n/4aGn8q05ByQ9cNoS/4zrqSw6SC32BP4E3aPIe2Dy
IHMCJdFQJDugqr7GKLX/WfAu5KUNzq08zs6bSL2LoDGoAZtC8t72uz6h9QY9lhQq
iPECLtrsjbNmr+bC6pfA0orEJSC5LTCtKUCbeLdQsE1Hb+m3DLIKjyuD1HSX4VtK
BXEeuoIScLRAn6RC3wUkQO5aXH5KT6waSQbacAXB+rfdxhUeSy7b10Xl4Gf7TfCu
86l3DgjciWTfCtw5Dr0VatPJX9rPU1l/DnGP5OWnszWb1AkyEsW+piix5y6NjX9t
`protect END_PROTECTED
