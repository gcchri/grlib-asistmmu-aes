`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZEXqtvQwomNKpUng6q54R5cy3UrlVscqr+7g6wUU6uCKlFWlzHDN6Cb9iW0u9tSb
JEaVXVXROY7m5gpyNHades/+effzVyG+7NCqN39l0VQQ0rTkNIGn1nf7m3pI13qq
hq363PvALnddtE3CaC0w3OXr7CimSvOtUcJRV6s6EyTh+yuVteFidIwG3fYdX/4w
lJjXCu+5qvzP6j71VKtkLgWwriw6abaw0V+XAlAXjDIa6X8TdUD7AoWGDRF3eonL
BEr+d62y8Pvj12NZ2WfJpB0YWUxkHtr3Bpz3GGA35/vUyC+W0BfjKd2fDm8+opA0
mJiSJKDuvU3Cl+9s7eraLXaOU7ElgZTtMDXRILVtKl5hMLtmS3stGf8KPnbRciB1
Ezfl9CIRuOl7sJd5VQRgt1vtwPDbqQZOpwCtYpoD6os8/jx2wLoF7jHVb1VSq7w+
+vqhtbNzJ+PdZaekK1r1AJMrZQMUqRd/jvTnyE+8F/ZDCLvmeLcnwERfeb3+s56L
`protect END_PROTECTED
