`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HzGN1XPojeMxDVp19iYTNqfCmv0LOSYJjU5T55eTF1PV8jxOPbedxV0psnmpjzbg
mbwgux4IL/XPVwrQ6K0DW66xAIUUKGBLnd5rk4FxrssWGsIOP+qQB+l9Wx3sv/WJ
1dHAdwxAh75nPGj9r/kdptV/+gVCskp5R+nPlxac0HumU58m9W5GvHCgeDjSaxHc
wgu6VTRz+A3rgE/g+LhHX1Mcnazf1TINK6/Db4PFBoJVnIx+9D1bI5dwvSra3HTu
MOwXE5JaybUdO7MJbjSkwjkeTuwa54u4vdpXu5H6SylWzmZu44Gkh7OsN2HVkz25
hlUKrcB4fpfm7f140JMA2k4OMqjlUlmCQ7OWiaPiB5F2G4FvCbrTBlvRcaLA6Kbg
fJ845k/6msniQvjgeagyKU4OHRokaMNIrjLdEWHdnpkpPIifCy2UJDMYgqyRoSMd
ckUr8NPUr5/ot5pQSIVakYIn8r/9Z+b2S62rwGVHhPO6DWzLZwpW8jpOg0sZozzX
8DH0ryZXezOtr7D7RFq2BegAc+8vpzMb2BUqUTAkQfbR0zv8CQ9Ol9kChgnmDpuw
Be4lmcwEXYfqM/VBHxoRCt0DeLsfLF+GRip7ca/AJlPmeCzEZiBYrq38Cz+xiwox
ZAj3Uk0S4/okzxV9r8unaXv7D+uHTsn1tKy1RzfAHJIZihlk7JdMtPxmVUCpIFfI
Umd4hXVxWEGq4/6ww/c2x24MFw8GTezXNRzsGyD6Nbv8qGVuauPcI3OIqtKQMSwM
/F8SpoCWyBwWB6KOXgHnTAfwY5k1cV0BlOy+Klfvw44eEjYqqDehcH05xZHLpLeX
Svby/1iEAkGLp5atC8J+vbrGsLfrqDx686fjxl7BSBngd95vrO21dxhTSKS9/no9
7qqVAHMzUOwC6e1IMDWQcMTkeSdeIzeC3t4zdk3DbmKaQW62UbgMRCUALv02glwQ
SZp4La8FNQ9K4PSnLUNtk3stu+P/QaqZExjofLKgAN8SPodt9KOuqOQKKkLX3E76
B8yF+8smDt8B15sz8VohAPliSeXoCL57RMKpX7IOibKUwKsSi2Xx+wIfdn+pysFM
BWCSGBdCM2GJtMKZnagae91QAZ45dPmR3yNcz3dl1Q2yVU52PBsdfXTwqER3IHFI
UBQEJHxsDDGx0V4r2iDD6M9yoTPvD0tKAOvs9GKux+DgLBTeHfCqMt7YIjgETHWg
7cY8HRRClcBoHXTIVP6UXw==
`protect END_PROTECTED
