`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xQjzK7oY2jgj61TMhY7NL/tnIl4Wd7CU5/4y9GNr5XxkF+wrpseibv/8UO7wSVG
fLSl0VOpLhp/kqpui6v3HgNVKSqgQvh6ekqnzPgvtSSO8kL9oB1ov06xkKXT5I9m
JGWqcQN75DPbnLvBnEN9Mg1pv/EnURnOG9CT0uzlWfz4Y7l6kJ4Mk2p9DFe2de27
WVxfWoplmyQwrHGEU1D5VNJBTI8+2EaK6AC3F5jvk+b5k2DBwGPQl1RCRNqMrPyx
`protect END_PROTECTED
