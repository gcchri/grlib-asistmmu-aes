`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/ZahFzJydrSVrx+U/91goPXNI0MkDfQHFMKs2STUfj40i/k+9aWRIliDKbpZfV4
hcczGnEe4mTOF7nYa2aquK92Tp5GvkX5herp0be5P9qzy4J7KP8zJT1q2bPABs6q
KiejGBEoHfsPWA0xiMLR6ROaHR9wqhoZU2T2IUYD8bYXXERS5smBhfFLY4ib8o0v
hR6siqMI0TaEF1Rj/1vv5L0uo1TRKjK57IYWUnr6AM3Ga3D/P5KFuUBLZle+7rQv
pfvp6axrudRW/heXyjlreRKMdMwK/nt0lQLfPIT//CIoXLeNcYVviUGKMsUPvcbW
NzjehXWJ3kGx5FyrrGl+G/NcdctRwyfFaKf3sc8qz1TKfD5cJ8Kn1GXKrfD2jc1e
iQhuHxcmKimWjChPbEp6g6kL0L1i7joIO/zKqJWO18BAvSerjj4e3QR0KtI1HoBk
tpNYdzctDHnxd0b8akN+EIlRuRTaKjjr+KztYx14LLWekuL/6JF5bARwtFiCQmaX
fI9gxNeBwu2U8PKNQ4G9uAeGRADbbQCMt+y2dbU3yzqzIeq7HC33anRNJlI9FJbL
9vzec8yl/4xQ7H2xIJx3YVH0SadUFeb8LpImyR1wiZyncQahgTsNNL5tbM/PLdtQ
xH+MeqAsZBwcDlDM4X4T3q/Dcmp+s5CqxXTDw0we+TmZ0KjA1pLmeo+PuK8rP+c3
SE/EVB66PgBJbbZW5TGaTThGgn+spqpLee0IQ8jtJUyR6321pQsSLypv9qdEViOQ
fSdhQ46p6WO9kL5VFipRS29wFV+iOx7u4ZNrf8PbuLhWyLm6+02MeG0UNKGLERMT
EXhndSHW+TCMx288TUdEugV2g4LytEC2nhDSz426SIzUVeNSoglWKLZ7QbMyZ3O9
lz6VGpUzADjpGV5rpkvuyCyqiXMcT2tPiUDyO5E0ijPh5KL1rjyCW7dJ+PlEB2Gi
lgzU4eFxV3Ko6VvDaswkPHf348Y7SccJQO2VmnJYVzvj1VSz8qbgh/nNxh4j96a0
4y78nERgd2dKQUhDc912r/96in0SbIvrc07vURkQ943xgqXX8oUWscn7YzY8/b7H
7HpKsgmZltgAP9c+tyyqNBAhtrTdEnF/zmPu+bAgi9x4Z5kGXm9jBS/2PlPoNTN4
FjeZLYOThEWhnZ/Qj3CqVmR6yUlquMEtZTF+gjpKWYg6JWacciCArBeCq5ZWZK9b
OLoZadMAjqhp2nIuJz4k3Ffkqvrd7e6/ndWEj15aFg5xGDFtR/VioB5dRktu7pIO
e/gbcaDC9AQv7a/EJHwJW089SRdKIunzVqKuQ7Eyafm8SAjZiF5Je/b8lmBUnDeh
4vqEpDwpkP5M5rvVXJb9fL4Nkg5/qoAgd2iwDXn+ApgpOreo8WGynfc4C3uY75xh
RiPwTylq39fC5Mso/tBUvoZTRVSUGX1oFMSCbVp8M54pGrQtzYPBornPzSC/hVDo
oj2Sf0qRXkoDsrXhEuFYZjXZ246lVQFcW5n32DzFAqyFWKtxzBsrJIZCRKRADMtK
7MsiRS1qYglnM7HxJtK2xhFZr4iofuKMP0On3aFu1nr8u7KKDazFbwSojomiUr6i
/Jw2ndnLvxI4YVqFgKKEUCDBl1KVKv1Mi4sh70iEfaHyWu67Tz9+2bSTqm5TpED3
73My35MwAdbTBegjyBod8yHVo1kWlqUfajd6DdSaBGy0NBrbb9muiQ6fTz1IqmwG
tUaHd9i8D6MQwGlbXyQlxQj3syFdvjiHNhF2xT5rfv73OYSf/gtpec0Y8mw/IUyZ
y//WZ0dm0HJkdrLq99z+GfPAVgQfjKDDIhV7dd5Kwb/m0G//mhlKyFzjq8kgARkP
1PrUw4nSq/7xrURHA1YUBMsnVB4zyGJn6Z57jXnMLtckvb5jvyor5/Vx7LrxTT8v
IofOuPeTv0Sd4CxD8zbTMDoxzD+lPg455AvZzSlpmkCI7NAkwNhO3Xie3X2d1BiC
xT7WDYuK35K7Lne0QWVCMC5Z0E/8mdBNPUv/qOydVMhnbLo06OIAas536DV3Vb1c
ejnIbr4QTMvHEdchtGEHihnXfepujXd6Tu9bwfnGScJyxBYeHzUAmwQmsuHcuZFv
nooNEimnrX4cOZKOQ23Cmf67Cl11WRYjXYGFNNGzTZp6+zWhavc+d3GTN/wn7YKx
oKa0PZFpPezuCBEvXmcSYJyupn5mZ1IUy3Ffuhf4wGOvr7J7gII+TWoGVmK2aHgZ
DkgdMkAwew0YmmYK4TSI5hHwzPMeOJfDYR6c0ro9i6UZ5JPH+GmtrIiXCHsw7esV
2+1H4h/MRRpKYGMmr3j63bXQnxiZ8JezWMZ2sgDpU37DdrH204sqdHayj0Pafrzz
6Z7fs+rEFioKSiX1nnvqkQ1t1tX7ME0WeshhxhXUQx2TQ1wgpiKIxVO5pxuA2zt4
d5Vz43XhtwyDqjt0zYkSXatwp8baN+fRY33O7qjxkly0zYiIRiEmeHGQgvB6JPtM
by0gn1pWXyUTgpj+FKN3YQMUNZBm0OOK8Ii4Dj3xeizEykLeVcibRuglngilqZyI
nQZP13F1urbl6FkdQ/vu41KfguWCnd0woQ6h6IrU7ote0ajLXhJc2zgzbEeNLC0C
G95K+QIXJkPIErTw0JQHSkiGFOkJAghNAansxo/taJsDge4yn0h8JQE6hylQbf8H
WWI/gE92DwvuY8SwDkXbgn6LFM+nKcud+EURB1boq3YZCDXP9Eq5o912hAT520cN
IfC6RlYqKjAO8Ic+JtBFDDNxFEwAWegBfes48FkVppyIw+KJx8HHwUtqzLF6trie
zJSqPgPET6NZ5Cv8iAjeJVH9lpTS0VnAPeG4wvHeKk5Z1BbGAR+/avhIlrps/hcg
ks6mA0lUvSeRlP5jysXfrZVj/S+IgPbMYB6CZ1MJ4qsSp1v5sXMPJt0tSkeP4S5c
StEtlFiqwo4++t6OxJil+IhQ6in3Ng99ARt/1spo58tzX/iQY4Z1YVpdRK+uqUNc
XbkD3WBKfjg7g/1zhySkEVxzYOQhdWO+fgDzu4HeXqimpjcl9ygy+SJshTcpT7tx
4FmzRI1hPMa6nfBmWyyNW1unnL7/l0LeQyCkiCxBIASEkdJYSZv0MJ8ay8LqnRSn
yFOslhis0uWIRfiPjLAlM2VULyXwitjGF1kYBawwX0vaisfDjQQVm5COBDG8P87a
x1wh/n4Tv/mUMa2Qao57EO96z45LGp5q7VXJqxgS42IQ88rxnIZqsqQCPHPCoC6u
pVLePlee+Sf/mWDqpMeEHGJxsmPz9zspAnYpmnmYTWaGJZtLuIV4HDibMXhw2xKU
k2Q0qXT+TXjtYDxADNkGwILJFZXs/dKYVddWrvj4WNpsItjmRLRczYdmCq2U6zI6
fpQ9kxzr83O0Pn+M7AgoaR8niq6KPyWUCAbJoJMcBLHeExoPkekgX9nouohN0N6l
3Mc4rIl0ETZSJDwE+RvA3xCA6U3UVetYJjWk9a+PkIRxyncMEmkx61ak7jqgceAu
UQT2sOAkBuqJLLbOxST1OevFCOefr16EYCoHuZjeS+j406+cp7LExaLtaSPOiFpO
tIN+aYo8p+F+wbrCQnhKuf1EqryFbJvBpC8ciVVqbb8jWcedYUlTh7K5TGd8BLzr
mk/UqGElJ8jJMm1Wsjg1A6xOT2dGnO5pO+RPVgp0YRAQTq/WlEei55AWNwj2ZeOR
AEg1VajCbvaXih89HXgrE3/6hAutSvmBVx4hzXpGFRxEV+o0ORaXgYQMXRpOLFf5
HpXMUWIuJj0DzOnao8Nu9uYWh3nbzgaR44C1yQfVcQVLZxkxioZl2cc5cfIS6TrL
PjH4W0XaOuB3iyNVX/x9WGcHr6EoWI9Qwl0cpNxd+q6DV5tSr2gxiB/f672CgSR6
yMV4EtbTuzs06vmSO60M+iuZ6R1wm1U1sp104gEcza7DmXY3XZTqPdk8YIQhnVyp
XmG96YWQn7O4RC7alSTHgIqnGq9nM6oQs9pN4XCjVtaGSSIGUG3UzAlA1pYABz9s
QPjud2WpJwKW1xV68Hz56iXd0TBhUXT/+VfrMl8DUZvs1WbXQmIi4aca9OdHIJSU
e/9LSr6SaJV4SPSPek/xtgEAnF7+S6nL0TaH5giHcEO3d8FV5kIb58jg5uHpFVak
1MVtRLFOadHDAuWaGZFoAYad0BubZl7AigjwvQRMAdk=
`protect END_PROTECTED
