`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fI0+BcBZ1HURp+Jcid8OH/Leyrw1lBbnaMcsjKLqP+YTiw3vOxj411NYMuuzAjEj
AUa4oyTb2gwUgBdrveU+9kQpgpBQPOuxev3V/qcLvIMppzd7AvL1OEaLKjXGza/4
YOwtFkmSVgoz+diXYMegIB7A9thnCXj2owDPFkQKQUgbxFRvkfbJWfd4tyUPqUep
Lc9vw6heD9ne59Ak7jSf9LLfmBqmwNahVJ1nw0kGEAAqIeRdximD5LgsGmwoIrCd
RmTYPc9lX2OppG6RIwzG/u6RwdCFOAFI6IPdGIM3eDkw+r/Ul1RsT3NL5DiqhS/G
VW9OVf52SRVeZ2OtpMnZlxkhMuPp9evjhOs4//Pw2lw=
`protect END_PROTECTED
