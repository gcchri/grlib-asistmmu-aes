`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7KRTHyPBPMs3sseqDBUDcOl0KveOOYpCdTn5oOQ6QrXtphK64jA62vEmyosTlAS
SS0qbSNL126GIDTtQIjxKS93IE7mkAw75qf6gT8NiopHRyd7LvVypp5KXvXGfpYl
+g9FDgxiVuwxApiDXY9NK4KNGe/vvCWBY43Gp/D54ULTHjwgTwXsR02pEIB+KKOW
0VwbjV5ZULsUmZEwXu2TXhD40v6eDd+UU9Vp+4lB1vRljzbc6/0JuvQIKA5MZvQs
4xE45IbTc7WFHLfRfiHmyvrwUWo+ERv55HKB1CuKfiQLOIUCl80uJMtMFUE5K4Bg
t6+Dos3l8re5XqRFaVRAQ/G4+AESwzRqVEzEIJ+6U+jQiyk2woW7QiBSHWn6gS2V
VGMnZwlbtGwYLKWKMhuZ/5lnme4GWxKUlkDkqlGiVu4aksbcsrbAd2H75tY59fZo
bjomU6JOX8jDTVgZN9DjQp06hchvtlwtTAZrPrUR0ter9ngAfkbHyxuSLjTO0aCg
DLC780WUGdOZz1g4DgeeOQ==
`protect END_PROTECTED
