`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWY3YrKQrFLwMZdBRtlzxGKC2Rr07JOZmAq/ScYLIYNMteXBhJDgy2Yogvy8+So0
OCEAaVidieepwv5MIkOUF8LNWuzsqYRFtg6b9CTJeiLTbNdiyPlgzG62hMUPmCPy
6ET3MJHfAgd0o2mK18yTO/8efRLhMEurBGLANqZW/B4OS2ZKSB4g40aYXn7xJVYV
MSA9VLrv+EaXJZd9s1ioEr7pi8PKBYG4YaPaP14JtRAOQARqGvEdPVLDm8c0RQV3
iou7P+9mpIu91CCihrda2hF4bn753OIQ40U5B0FLqiI+owpdr02DHRihf6e5uyVW
9/VqtV8mXt9HbN/4Pb7ZvHXWe3BP06kFvyBRTNGZ455kuZZBjsZI99F8GgnGIo2E
TTH2xXFdDPbOu+KJfBROLzi8H+EO/MIIeDTiFWQHsB/4PINtCCTWC5fy6wIBwuoX
3ip77HDlDTagj7fjm9KyyCzCwZeS4ciqQaTmw/Xsc522Y1x0oh2FpkGwxv39c/9L
aVk7h4ZsbAzvibQiHKXorgrSS5Lq8IZJbFl0awZFsKkBF4qnn34SOdWMNfCRfdlx
ZA6TPthJosZMbMVF/FzL8RoXAhNVYhSoiTLCofAvM8MFLJwFPABhVe6uYCJCkeZ3
+d4Swxx/E2mVZDhYt4OBjxorvdxgxEhRa0Lb+1060gxApuc0SRfh2WHF5D73Tcjr
DT/ZALA5DzARMbxrFrZ8UaLndQY28THne5kngYWBjWPj+xzgzARw9nfxwOIzZFzD
sH8vApsFqZtqDtkk2LGWvoju4xoGnrlPEwJNOmdFLzpq47NQSKb+2niG6th00/+8
JftwqrIohnxFxhMglr3sq3B5Bq7HTeswmbd1dRA5cNDi5JqDhA/FnsypTxb+pwos
mhdVw8j+ao/hzrVprGik1Q==
`protect END_PROTECTED
