`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9bHOGuy7wbYPt2+VJKAdCX2uXuDyvAfemE9Bd6AVG1JfvwfzoOTb5FHHOlmWaOS
xdNRdbTRivfJKwNuE0UPmjSYELQnjWCXS5TJ3tyVQNw9DbJDFbPzKh9KayqEV59b
HAaeUsjEeQmoeY2dH1VjM7dHkzAWAVxwK8k1tdJlUHF6HnBWo8V91waGd2xDdJw/
u7bsDcZ9zwnUbbjf0BdqHUqciqVPVv41VkpmUJxdsltiXN0yZLBzO/UPDIqkGmHQ
yUqlcS9/YAAMaEkzm1ukuOuOj4lRMrJ+o4efVjHpD8xsfNoGeQDEjwdyx0CfK3wS
Uu1Gn4P2tBqvMcVR7BuyAgiseojJClgXGi5cKZY9HXjq83EMvJecL9Kb3wiLLYj9
jNNK/1WCjbiCjnMQobA0ts/XUkX3rNbY8CgibHCNFX4GijI1JulJBUwVCp8cuV4I
SBqXzy5Eytm3aQWg2s6Oe3FiTD41m4VHVVwhYgK7ys8cQdg9izRIkSJztgrdsWj0
NfnTe6i12ijMA0y42x9dxB3K45GPz2GXRCVaHP3E/4MCahPdBXRV0gChvOOV2/+m
B7Wo/kBngX1GI6csXti4uNpjMA2Mwi0DZCHRqWWxD1a02Dh6RvmXMvvBt/X1j4CZ
NeV/MSpqGOnR8MGHotzPjaNpsxga3sqE5/Js7k6Qy0jn0ht26cc90RmF8ZdqaDGW
zExnJJG4shf6RPUdLJY69cm21O8/ZSo2gU/LKBqCnk5JpDtNYlrcAEy8tcQu8YYm
g8xuko+8bLqCNp+Htng8VgDUJ7vbHoWs5ld+lh0B7J8isAGGmtfGsW5aUkgwxpd5
cGkaNxTd0eldr2MQnTtme1Dn1j0pD5ONlfzVjVQlESoRtGrt58LVvJpwsUK+g08+
VTTdLRBt5uVyE0IdcHHqKnqpifh5vPJ74ZijMD67+9pZl9xhoAEWZD2JKPZ2ZjF8
F+6kreOJ8DTuDrluiH+TwnjirhOohLJl9AlcdShnQBEFEnwwX12t+FrGilLg661A
9qkWY+/0FuCzXD46z/v5FHa8V7uN193eSHgvEK5eSklyPKWhoFvn/i74rWfb7duD
FzR0JQS+5KXO2y/5tT0IVhRmuP0g1f4ZCYfDyristNXurO7pbDJD2wWplFRav3W0
er5l0DSqTew/fiqcuK0XteeymeLMWDHmp1NbIDdpw9Lhly8DuutDSyw48bCuoVC6
XOkyTr3Nj42rImfjQ3Y/oqEhjmwVL9BFZ7+EvjYm0yqZuSB6BZiYafB/C0ooBx+l
6gmTbWJc/Tp4K9opPQKtk9jeDM3UG1BGaHEX9PeCc2fe4DyHlfpJO5pcFtifasL9
LvlznYtMkMqwY7WP/qt6aH97MiFD2UwaRDA3OmLVkXkeo08T7d0bylTYHpT2azWC
aA7sffpzUTlnarSuITQC85UqaNBxvU9QQb7YULXHN+rsekwpH0uy2R4ZYPVGSpn6
vEfZa2TwKxQ/CWnu6wJdXkD3VO0Qxc9Y16ymQqKRlLeDJ2c421F7N5RmQMw6kUxa
IUqxNdNJHJdpBkqMdNMEAea4Vy+oEHHyROElfCdZwrYgDSfQyIh7Eb1PDdtw/+zw
zgdi/LeAD9Y9Ad2QTAK0rp7nYreTdcS8W9WThueiwO1Lr9AOTPv1BeORbBlq5e5f
1y7+VyYxAYHdHhD7kI8dxUJgFgJaS4W9ItMZlt3zBcM+fiFyvcLp7a5EjEVFPYni
p2FnAvnn+rDWTaXsx31sJ+HmeMwINUcizgzCBCLeisKG+/usGEiatahs3KQzrWhT
fVwFA2+Fz6q7eBYVGo5knxaCMZs+wSWuQd3D/zfmLVLoMpC0vCHvQP1hEHOBnKQn
Ob9tvzchhtX7oSqnzM1z8i9hzU6TnmTrh1CVF9/gymYP+ss8o1rhIaMK0V9BDAih
MiB3ZC9ZFzdqLa1eNDBlJ/CO8wR2gRAmWzDSLv3WRaQEZcssTQkCtjdkD/WGbmv4
BJovcWKOvmuUCWKVXpgMT9biGtx+0vK+9SZrCU50/pHRzD2G6tACbZh7N4kC7DZX
ogWvkQbhPw8ynbvie5YjQGrhc2IEoJIPs/aYUWH9d9vE0zGiJvk/8IL9Z/5CORRP
StzuB+UjlwsbjXqw4P1/9TP8r0QfI+akg+yyKDV+2UABFL3+yzXIaf6T1503mYEl
1F5vUXuTVHTYQC57zeTMsXdyPAGILwHC6QslSbGmKB5WYsk+fYG5PjI+7eBY9gWB
gSPjCS3gD0mH3Bm2229I0MbiLD1JX+CcJJqb0RHNyHhivKAiuajw1hocXitMjlIb
cWXDNk7XriKa4yfVAV2HBftYrT1hy49K1gvct6cYRxZHu7sKHqSTBlfSbcdEN1wL
vQKsdkEvnyxlHND1Ow8/e1yMCix932/Tfdn1fAF0TmSuCkbyEWohuDc4e4nEfeeI
TQ5m/z/oZSi31MzfFmNrb3NNl/7V15t8ZTXmwExvTC3G3EAmvTpfZS3zE3LgZ2VR
xMBM3kaCghjbOTUHEFZrymt96LMFH3gycuRGUpoB+IwzZTV9Hi3UaiJBe8Xfy9r7
`protect END_PROTECTED
