`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zvi5X8AiNLEoFKvbU5SI1cBKo1Aht+TE+j3+IAFyJZ0PeiOI/c84gVxR7bjZrcL
52mHYdkb+VYCQDpqOeMq2pEX0vdk5Xp1FDRW5SC6+bULVB6KYkokioG/2JEoro1T
HGvEQqP0b6AFg2wVZi4BgIVd8ZR5c+idOuawA6YjvCVenaenYHOFw6xITDOwciHk
Iv0DUcnEJm0PeuSp/9sHEXuOIdK0919LVUqVkyKZStEiQJDADQmrHsbZo56pOQiR
BxJ7pNkdRq/c99NJ46ojVQ==
`protect END_PROTECTED
