`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ei+pHWSVRo2gk86Jk8MC5gefdleivxBWuFyNE3wDJXPPWEveDEUIszr7M/35cqcM
FXmqWoZemdp6gGnJzrapS1aeXlxcY2EYbytUI5IkhLH5IUK2CPchaCXvjztGcTmb
81XDKxdHV3nZwnhb1uytGkGONPE6IDFGv0NoF32M/qM94fIwzl3xdRrZ1JASXKgL
1Z8iuw9Pkf++i9I1JWVDa2W+qENHbEYVjX4gr1VHwxhWdLYqMRMJ5nj4ktrbDlyR
3jngPk2mmNdxj7/Mhwzg6rsIf0zf3Ub3u3DxR8uOjW8WrsOXei0PgeHm7Tvrd5Fn
coCQjjGMdORYa+62ICFbkL/Xbfza5NaULGtqvIW2vVxKzX77X/FzCRfsLsW64Xgc
poGRZF5TZAjARw2+Cvz1aA==
`protect END_PROTECTED
