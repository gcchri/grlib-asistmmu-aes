`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FCuCOvaH+aIY5N7CRwDbUvsa5JAQk6bomSTiReGJrBHJkbg8gYObHX657yifFbo0
mcsxS1NrhmYAqtWrG0XUwpbK3OT7/8Af9vwroq7VJGQZ7W6mzOqKvlPlxLzJQgZU
nXx8IOVRhEyNQ1mhByW4YGCliM10ynfgLpOMQPdSyClMecd3jhCBkh3Yi+IlkKij
8wwE7rOoHBkLtzMMwDHycCdle7vS6bfTjhxHXZzYkNJyWi92gk1OAWONGMUlf8z8
1TY+uLh7OBv7V+aMbWveoAecw4NM/S4ipxQNZj8ZvaL3MeloFOnBjzLEJbb5CrAS
Wga8gr2Sr3zXH/ZV43IKSp0kZLIwVBzEfj2SavCP76M3r2Fc5ENMjzInXFR4V+yu
CXG3cEvxld7ItkwkpZwyYJj1PrHRI43/N3SkYeK/ktLNSpSm1Cy8ouKjrFuvL54I
IK635vNMJaeafwSdpjhme+1la2I6XfixdIa+gihvy7RK+zEPBsAkBQYalsVi8hog
Wyq3pwpJvrNGJ0yegRXvfw==
`protect END_PROTECTED
