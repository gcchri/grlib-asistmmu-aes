`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRa78Fewe3MnTYSsl+H4Ay9Xlxz26uMKAEXWvFRTlDz5jagDERIjnhJkOrxZlbFn
s8jyyA414bFZGiyrqqLCys3x4aSm1VYkDCuiAeBVAynhpVaDcutiItO4tGFt5YbF
VcLxxSbxW/R/7IlBi9DaqYDxDwLNPwFE+ZBC6MKbDn22EulB9dSjssITaWDJY8YJ
YF17TldYbnq8H8GV/W+0gghQW+zNZaWIvS6ws4GojWFLFKa0pW/FcvfBPzs3Jgul
C2ASKAeeMxJBzyjSkSXFPN3UTCzpbi444l5tM0zZnDVlR2IUOr4ONKXPJ7EfVufN
YdQb4vw1CZMx5RaOvzT23KEr8GpZGGlkz7IIp/zpLbJ0DdMIRWyxWFKHmW3zi6oH
8nEMp0WJNH2qShrBJcJFChdGcWRHupc6GFBwA8Mdcc+e9V0qVJCwnafwLYywxmLg
NmQfVwTFrbygzLDHa/QyBJC+Injse+rjrjbYyrF4u1HLP40hfg++NiiJsLRYTpUG
DpWsTa8r8yQ0HnbhgWLOlumM+AQdGPqXqpWF75LV3Enk04E8yNsRvFfhYXrLH5Mz
ED1ea2wlZY6WzqibcaCnpYFGbRICEPnymv1VmgEGjw0YZSDyicrPqGd/DmuVaAB2
T1lj3fgsPY1b9bQLP/HkxoSsLLYXnZiLAp+sjNTuzKuf9dgnDFSOiP8itGsPoKq5
gmSPefCM+BcKAjgQ3rpJbwRj9NA8L0Ko82oLS5ecYDKYhPfuoR5aZapf8+7DDDo1
bdcAXCxhIJ23JraJIK9NKShV6Tqb9FPEbPOOcE/G2S35qdqaFhfZcT5bRptFyHYo
3emYkwUqLhmfdginS1W4dMb6jBQTdiCgbbd1A6k2o02okBu3lT7cqURInFPZv1vJ
8d0X70NSc06n4y1X11VisddmZpthAuXm9Ki5h7lnUrs9l+8rbcE5Sud5XATrSAAa
SvyMxagenRiKpCe/P9croi8cK7ExHKhg68Aq0aw8CiOqw35PN59SOP+rLUWLSPmp
k083C835ZTB+naYnOgybuAniCWeOSHXIyk7/kMH9ZaiYuJ08GyPB8T55PoQZYDOt
S/Tq9MOaa7l33AO3oAOg66057JtZ10P6/x3JC650PxBLZTO9eVvGB07+QdyuvSUQ
5DGOxPzxyZMXntDZTkXKRUdfHCf6GjW6ks6zPPsouIevF/QGiz6RKWeeB2k7cU9v
4PVn4p/Y/O8z8zBRVVUdDpYZoDYhOOg+In1OJHQ2NFeSICRujbLSHnsweWlDwwce
P2zMzrCV+KHbLKPiyq78qg6kNxwpdHFCHDMc61PGZTSm+bk5kfXGuVrKPWfIdv1W
JiqEMBy75spaWVpMDZ1dNlgPMFLq77m/6srDu0Svhkaklwx8tkOJmsQWs2cnNjzE
sMMoyMdA12C0O4jR/LHB16b9MtxTmeJ2tBePOonhz2jDF7Trihly899FUoPpdbJ4
y8oquWluH042roeTeQMxk9YZkjio9XckKdnpuAaQD89rsYnlHq4yq9MSds2MPoRc
rAQBi33WcGZWibth2yu2C3/07aFHQ7deCwPoHWML845+yBC00D9IMTzG/4OJcwVI
fvm4sEypE4EFC+CUh28XMHlR3Ngt/G6xizC11lLzEmGwfcK4swGsNr/LtA/zUalR
rBY3FdDTuqVfXbzA1Tgyy8N7QY+wPQCOMAKso4ESLoF5frwZmKvtjfMaIScGoCx6
w338EiVfgiMVJF0N6/iETGQPCFHDl+BFjdYjkMoSmq+qwUuqcsY5+sVhllmlTl6p
Ygq7NSo7QONm2iHju7MkSSOf4T/9tkkdBhuvICLezmJSMm29MHZOrfCMXjZ2IL37
6Nozq7/AD4GQusLICbQr/3MmY22axhDxb6LcZZSOU3oOMPWXPz2GHDHxBupbEzCX
fQyObPWliqLb6MBJ7doD2FEntrwpDEa6lHDHTdI2DW2EnzLQE2Ms+JHY6Chd3fvW
Uvpl10nlZuSwb/NGRIazgMftlXCWW/TkGzHOFBmLAN+8dw9rlG0MyiwyGG2Ew1CA
`protect END_PROTECTED
