`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rUBQwRp2EGiN2CGvOUNgFvNd18qTCaogZo268EBP/AUHaDObUmXtpP6SmGyEKyrN
X8IyVJ+gTUMTza2R/MX4wPi5sZL7UeL0jRZ7DEIcojr2gr6GFd6/TgPKPch2/vvO
/0Wa9CcqXsEz8SgfYFFQq06zcQ8AirX1wDivazQZT5z0dGfwak23EbW0d+ySMQ5M
oD2ZZ45DHv+325Ya0LPnwxcZyyNNe1XtJF7yUE79pdkSLB7K7izpsJthAmBaF5Q7
/hPC6HGhSbn+SQMA07a0NvwwHCgP78g9cV7WzBPpwLmC7zG2GxAcRjyw+uUvS+Pj
R29LGgoMIRmqnb0NBa3OFSP1kqKGH/9IxG3tXO4UF8/DDEXptE/g+3jYM13sPJfV
m82d8uG3XVxngN50k0LsqlkGNHv5SbauNPEyx1TgMn+Wgwsk81UPgDytwn1KKOOx
`protect END_PROTECTED
