`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aXR3FzUt780KRZj0mIKpqQheRpXB8BqRsoOEPY5KdVAplbsxAlkE8Pgzn0x5yYQv
BenSGqiLkkAVNDohXqVwKI9W5tN/ETqc3eornJXEUKkRBU5MpKnNSdBxIKCzm42u
9CSX3e+RSy7xkaNfk90n+mxHIylM6NR1vZeH5R5i2OBPivtSxvf0l/PAbP3rZJlu
tQBN6h6DdO6M4Vje+sN2FwR4Kz5iIUpytRwb0nC3ABF+8H+0VH1+jMQ45MGPtbwK
uJi1lWwTVOb2qN7uqSDXEd7P03pHvKriQ7k0uGVrZeT3t/v6iuVkkNLfzKmEyo0M
oapYpW/so73j/Ma2YdY5c44rNUgUrlRPsf8XKA/e0ogdOH4n4osEnxLWFO1frPbU
sTM4km5AgT/YizykrZPR63CqjVp7dDhuj3LS4Lm53bLIWu2uj4uiAEWHJmHEeNlO
CItW29jSFEpDMJEaNblVtFXReuLmwd9huyBcAIFQVEY=
`protect END_PROTECTED
