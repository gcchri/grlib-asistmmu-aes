`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UViqZOJvPgp7pzaGR8eEOwd2Sft3sZaHVdIoit1kwF1u/YQicbX0CViQkZRtdKAG
qMahBMJZJghn25/I63ttfuTQiTtSjEWvX7IFY+D8OTfgsTCV9y2aS9cr32+HlJ2H
bOcS0gdVTYPIFuefT8LYVa9P2H8E54rlA0flvCaQE1ZSbxJGYwCUDXNwu+a5oWqP
P6yhYYtiUJ1oZsh1brR5v3eY07+JwyCKdvBaV2Rub2kD9+/qi8gcieEFmm9ZHdN1
l9T5p6NQXAD2uKIwodbus2CdgPcg+G1QKiTV33IgKgzbX02ceA7vCBetM1vimTEZ
VZcDryfMN+rWi1viMTDDBacKvqBPnEXjUR+rYd9y6t0cnpXfT5pXtXwSug/d4Tjq
G0zQIWyer0Hx6NC7aeK89IUkJ2/ga5Zp3hc4C2oh9ptTNWZQEihA44lyMSu+XV7b
a9SXiBFaGkj8thd6hRo8UJ2rr4A1Sj4L17aiKlznacHBZ5mVOulPa8rXgEWnm35l
uYus+NjgUFagEIiW7AvfR3UDfPWLjFI5pqIldyZSOZY3cIeIAHRURO5N3QRTsd5j
pR4e6eankA4v1kdJrmh52NfbQfDAd9eYRaSzP3aAVFnyDwjJ5NLlnGVsDSrQpe4W
FSD2mLVPm+JTf/B2H9ybof0qg3cdJGl8Kw+S1F5NxRYEMsc1u2ZG/WvCHZh//rfq
vEn313dLWFt+MzCfnJ3+3PJmIymntbyCRDybteFhvl8jcFRKhR84jfCf6oOnBfmk
s7SrvuwPzZCH/63RaQBcHj31Lnuar9b8OHEI5Ry1bwktA0zvMrDPyItDCQf3A//A
gqMzn8CpgHeczpxS+XsM5gf0TqLUw7583gjodJ+Hz5EC4Eo1L78xFMWqVMoBiPmB
haEqsxIR+BhVBCJIBkRUTo9pJKPMHdmEyAUnw+Bn/cfdLKaShWgSrtbOP0ds1Q2D
sLUYq9HbC6qiySsLzmdtQw==
`protect END_PROTECTED
