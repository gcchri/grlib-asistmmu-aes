`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8J2ZZml+dp6q9knIwAhm2JO8/tUlUL8H9cGEgK4EyUom9kW2veuenR9/v58tselb
FvHEerMA6XQBq6evg2TtwfILknTMTXN6S8O1ZuShNLgVEqoKO8V45cIhoPFZ4CnR
49d2elBYEQXjHfofDqXqwu8vRQm3cKlLqHuvlB2JRKwzArELW6do51DM/d6pjRJV
9RmWWQV3IT56YKiFud/lmJHOnnSM7PMURXo6o1soop0vu9hxbLWHhKwv/Qxzdej4
zwcvH9nUjyHVeNY1VuX9ZlTpjnfXEgYYLtsXlGccB14jdiaKU9QR+Il7C/4vPs3C
zHCPET7z06f/KSWmxYcSYpMzgmq1nJzPy0hZ0ethyAj/X2qJuk5bLUXs7SnpH+Xd
DnZXqsJq4tajAUevIydJAbTcGqd6LRphR16vjpTKXniX6blWMVOCKAVniNkxzNCb
LF3KNiQWHUm/SE31VNH4wOu55/H+WK64XgN1tLPY70HKmpz9cg6VMS1poSwIAMYV
qfacbCoGMcb+yS2yyQmHXxH3J6FGPe8GOamBWscIDKoAYzg1zrFELsGSZltYdwEn
wU4g4JeQdUAunKByKpCuhW48luMf/9P5kl4OQb6O8g7q+mKfMoeQSNUDLZddBnat
Y4xz8jAp8qy6PBLs2xO5CaYcNh7xqN68XhYv7PI6wet2gTzTiInuow7KM7Qrq+/x
q0zgsumP3WmFw+AU6a3DwEmIYqahi8KeEC9APUCyFXemieOm3oN2kAkO2W9MGUf8
uj5IEVVErJrAJKdrbiwwFuSQKYhWDpGSFL8dMvYgOJusWIYMBrcJQ3HAKxmP6X/X
zpc2Ih+s1yH8oStfRhNiFtK9/rDt4RWBWgnPPhxkahrtWY1pFausIwWCd+zrUUQu
K8n/sfJBHlk3seAdo6XSePVDJqta4jjOdRooYrvJWDHg22HBW9Fj3A5PHYKyYcVW
oHZNcGZCJyiXxsOvT1psxzRyLX7UaDV5+I69E62ZiJBX0zzw2+1I7LNE2mk4U2hx
g7Q/dd7PaUniX7k5SKBBNvZxHmg2pS3AhTgrWh1kv/l/eKElPHh/05GIEZnI4r3x
HWFPxXFaMAN1Nh830Z4Kof02vRimeLdLvxc6builYrNNORlqxgD29OssYUVZg1g4
sUpC5cOdMgNGVm0ci9NnF92VDMxyHu8+jYSAMPv28w2UOfu2s77allfW8eoSUDtR
a49CJjLzIPpxuaCGHNGn94n9549PYqvr+6VGlBp83Zu+b697KsHCPh/fl5ayPnAK
P2ZTGlzeyCZPUb2BQrGePNTB9niT+G0Ul9vDTwWnsLrpF8GXgZULXSOjKN9ZxkAG
0vS7CQ0lbYRzl12DCzwYSNLDJrLB+qK1XULVetf432L4nWTyFHG1FfEs1EySqwcD
X+O9AJ0xr8juJFlZFMPNzFjyApp3mVKni/aRn6uCO7zpvCyKO1cfO+qTXW+sWD6D
V8fbSxUy2BcB2G+zVYX5PekArCv2pJb3ZJZd8QZ+hKiRvBnq8nxAGi4s7xC2tCRE
gffnuB7GRLDpdclt9HyhMu0hEhTGDqSQuhJHXqDXnbgJBqTAkd7v5sM+7vc/0a9z
AjUvmt9ORuuAT80ftD8IpJ4rHaGiZki7vjAEiOTGnApeYpn9KYfYjA8s5wsPr872
Yr7l/KniRqC+mUDwgFIkWUCOXBENWaRVCGpPLHUAABXxG2iYbAq2x8+uBXOZ8soU
/bEjAnyxn2OIYQiM3h0oJSjlHM4/JDbUO4ud8T23GxEk7unrvHlgXSK6uucquam4
D+VPtJQq6d7OALbBhcsAcD7/xo9WMQE67ANn2W/YDP/GL8wsC0bnwEvA3NfhNkdy
LYLHLzAN587yeUpykG3ZkIB6GSyPoanDwOhdNSFSjipdc28hWNBVjTfVtCgZnox7
ChnblR5aRV3a/K+v164is4AEz+TEyGu0qdFx748dlYORuE8NEAtpvnmv+kiHhTw0
uH3jVUMMlIYSnHZXGl3iYlbLoxyT4bskD+ZqXL67I/mbfqEFYhIAahdTEaOW/4j8
MJxA1z3jKrdHuMaSdRW9c9H2PQm8v1tZG0fyevE03Cg2uIcH0gVimAy8RvIE7kr0
qw3002qOaO+xGCvU5OBggnn6yIsPv9IJRKzv1h+zyatSsczlnPZJig9OdzDAV94Z
gPHLO44+YZ9t8Xx3pr9LVnweUMzm8nE4bCrg/BoEYiC6DZxLbKvL54jI3jovWxam
T9LtJtsVwN26Km6sZEf02QzJRGQ7XV95JAiNZ5gjPgM2r7GocSSRT46NeXO6J0Az
f4XIee/zLCOmzsaL/7mlqWUPylmLgGZ+x1Ms/A8gqto4Y/lhqD+LZnaK78xzKEAu
Gq9LDDs6WwtdedMFHI3SD4vhTQK6kQUv7c3W7u/IMqZ2eoXFZ1BpE+uQdYh8oyb9
L4a3FomGPPKz9khUs82DIJ57aNz5uViNc6YL0nWLe5WtOfrP0SpDENqqu5ZEjZDm
imQYQNS/qmjhWNfWEmzu5jywk7expLJtaMw7U7TOzkTZOeqiRrNxOPnkGYEowxh+
5bQ++l7g5jx+zclP7bv7WBjj0+GD+JzffDIBmfgi2cXQsGiQPMQ/GbkIGwTfN6cZ
VJPTCfIQWpWFX5KjgDGLpwiDeaN4mgEWM2X57Gj9Wd9vDTo4vgDOgIsR4GQFOiWH
lw6bkwtgix2L5FJoQWjV9Q06c2CcfQMTV9xIH4nGkT03eAzUSAgdvasqCUzbk50Z
husgqFruVBiJZt5kP5IVkcDL8sH4dNhsD501K7gc6WyinoIQeKKodw+W46Wq7d/i
TK8WSo5DPQFqdvtVthW0S/xdVD89/MyTDSVLHYu/Az0=
`protect END_PROTECTED
