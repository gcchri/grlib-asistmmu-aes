`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BND0T5qG8HEDlKxvlGtbtpc3Zy+eIbastIzIPVVk+SJ/4azKW7S5jzCu8wuExVZz
Maqt5SHmtiOZeSUvoJi2Bx4tPIEr1H7oHZ+j9ft7HhfE3pIOqgtQnpskR4Ie8xET
Z/HPbZo/LS3jIWMC4Zb8Wa4uX1YgBmGtaAUrqxeHthaOw09kqL56h4vVElb/r4C7
01TbVO6o8jP2Nz+YdtdUGwu5dBIJM1wASc870HHEoRQ+Ppq9V2Gzu9DojXO2JNcd
xsQsYeH9cZE9KHT1M3Z5NWqkFkRD9RFbAkesCZYB/2Tx0YqkqE+e5S0384dM2opp
0snodCC5Dzg+LiAzZ+ePNA==
`protect END_PROTECTED
