`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1ePiUulOPjggCMZxjzbkdKVovIYOP8kMdZFi23imm+3s0EYqW39+VrfAYffU3hD
rlDJhVapyMRwIhF6PlPXcv9CYcqlhBoDjzebYgYQOvVQJVQkhHhCezKabJdgg8qW
ALcxsijmIqcfrfoV8R4GfuJaKmOR9yoOqLkWsrTYfi2Lrbmz/onKSAtGBxGOFQex
FyByvTXaLvq/cqNkENikw2p0ozDCThR1UTd/K2orUekmiv1uj08DBdoFoLrdgAfW
AvbBL2I9dlWq/99zrfRyCeMocMZ49y5kkQr94kZVQnDssQDGOx4oISZzK1JDMhzb
Ekm4vS7voVdcnoS7/lUSvEDXmeoTBmi9Pn/rOmwVZlnTfJOcLFJxZzUYh1SZ7dgO
lL4IK0E8GtAgGOMVn6e8ey+BdzPLsi7TZEgcMeU4IIVvxwwqG+8Vt86O7bVZhl1H
Na0Wnh6yPlp7f2RYFvY6qg==
`protect END_PROTECTED
