`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K057qWLT6HBCUeR+O0IMWyWyQM3DXxFyTJa0h3XvxxoI2k26VL8ob1C4ubepJ2rk
LN/2wDECHsMp3fB2ULmLw6sPbNlXPgUAjp8Czm92+jW1C3jux70Uk88D9M50RU/q
kLhINCB/tTfn4DW/EhVU2bkJUi37CRt2zyzx38UoazZir8aqxj9ouvWDD2CvnXTf
EcZD2WL1eXLnFIjiPj1A+3y30ty61c+ruILgDCXM6KYa7uVfhd3emIjjIsjxjb8f
JDi4iPuk4A2gjtLKfE+fDuqddPMeR0raSN1Do6RZhQNi8cJ2ODlc/pacoEH3krPH
g1nvMHVmUKqBWQTeL+dZLUFQ+xQS8KUI+msVeHAW5uQ=
`protect END_PROTECTED
