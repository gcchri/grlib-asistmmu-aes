`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6q+QebkuJv/l3HdB4UxT892ldk9rUOsKKaYQVV+rhO7gJzWjvTjRbtYkFZAt7jAa
fQUQwNHTjickwTwnZMaXuS95PHkPW1VJ75EmdZ80zrdR8C1VNPv3cGFy2/sBWhPm
iTUCDT2z4S3+gynstE6mJZfZnlYelC1TZ8n5bvEYrbTaTvHH2GUBfMGal4dGFBHw
eoHP6n9vQ/mbTgZHtbYN8a9kebNXJ9hPHyZ9o039DwoFWNHRbIYIHM7HAc0LKoa2
6v84yl/Y5oW36SFMrW7fwc0cGBwobDhCH9aJ3gCJ7NlQydaCPl34JCTabX1+hFb4
y61aA9SUXuoC/oaCEnhhebWu5sS9c7rSuncRUJy3j3v0+H0o+BTRDdvn8e2VPcqn
UwuCT/efMMDPKraOq2CMUZgDlh0zrXRKgMVeKbe5ShSz49+t0XtXGMi9HeDkC4VA
nuQxCjbXMdpe4KoQqYHdZhVf/atzOTOqdY46L3pnNcVpHCz5H5Q3BezddGuoHJ3w
7LOCr2lHKm/7VWH0UseF2LlOypkQgQ6eLUeXjEhD8rhhxV9RkHdjSi4ImYk+Vuvf
47TGZCPVdlYa99Hu/tQXcvPboHVrfRD9ERCQUW7FZPYINsDEhmEyTS1NKe0wC6Pa
jV/vHYuwiib+IMHw1Vio6v7iMSQh+kiUoy3pnsZbYE22yXQI55nC5DL+soHS+mtt
JuVmAOdJhZqVm4QXqTOTGpiCw8otxBltnNFutOh/XmyfTqTLgsmi1nPQIPuf/WDh
reTRZRcmJ9KEKTaSbb8yqTsjPkg8c9prauxaSdbcEt98tAG1uAzZQ2T1VgacxY23
W1Xo3maanVHXbi7p/t7L7cualM00AL4jGMk+Y6NVN6LqDMgtO7+JV9ejMXgLLi1a
TcvtUA7w7+kMTDUYG3OBGc/ZFOdhdrHBI5ona1XhG1TletRXADDLpKvfBsw73l0t
3B6WaG+cgeTUlzPEv+f0LclvpY4M2+63fClGTzhWJ1Xn3I81ZQvbrWh4l7o0mBMc
oRoxJvIX3iPte1VE81dFIQ==
`protect END_PROTECTED
