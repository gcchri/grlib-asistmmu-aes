`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wsamtNrVHgEit4IpAsjSyq4FM5aKOrbxpwcAZ3QrB+jpp9pkZO7RmyxZaJBIlGJ9
iibm3tjwr+kF4d0tCVf3SwcS/ew7VAKUmep+ZH5ZRzrCjaMarKKOCxVkIZpMrH9o
Xw5xMNJPWJ6nZNlMc6xWxFIBxCzhPhKpTavSzz+skw2diMVkmHuOoDjFwmGbGRVT
ZPOUkyr9T6uiBZqwnGyY7gsn+IhUDYP6QoZM13EQHykyaT0AUFppg2wH441Ydmz5
n8WYXBh0PLx6ifY71sUhjRINi7px8v2UcqujO+jaSBSQp/4tfooEff7StMt0d34F
J+G1xvtyKKeiSVoFK+sQ8UIgf4vxxlrRi2vn0GloWARn8PZJRLxsh04Nuy7LFVoV
5exODYFcEQiot/qrjgfE6A==
`protect END_PROTECTED
