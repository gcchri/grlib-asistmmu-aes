`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CcKEgU4B0owCgjI82IYvceaVqiHdfJnhDGfH2LvnKZOY8ZNdKphSVKvZBJyaC34u
DHGxdgxTAqxpRaa/EDcDTpvcC1oF/AgicdnNBlfiyjJw45SzywpFO1llQZykVeHh
XlHqk2BuKl7iLo3+a60ApS8rn+Km+BSdbCc8OOfzdzVtiIk2Xnib1azJVa9nPCLT
SGiaRHKu5FRMKdlNEFaAemZKcOR4VEVMHWiCwbDZEvE52leNGi0Iaz2UYX3xMSU+
K8NU/iuqyfyO5CXkUZ9P76k9qJ3sb/1bB4ubmK6a2/k=
`protect END_PROTECTED
