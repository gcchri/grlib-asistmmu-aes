`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yEcxkX+9pSQMq8ALWJMaYEo/Vsobuza05uF0l9bsZnnZ4+fHxtLFaOunUcKEuwfc
tic6MPi957LdiOySynAlkQp82XWglMReedEM6Off8yR+bcIdhoYSRJbmtos7Xng6
lpkpQflR6LAiD+vDN79WHbRpOue0NZ5G3SNnUB+v2j3jrTUKujAr4b9SKyF9P6kW
jl71+DSqWLPWbu63EfzoWTXI73pWTYCR7KIW1wjfhOqVBppqlXZW0vMXIx/4iZ5t
pLMkJXF6R2u40arBQpC4sGRNsGEzI5TqmVKRDVCfeuqG8jJw6n8VYKvxQPZ1xkDQ
psMIocnuR4eeUmV+VYjrHHPP/mLJitQtQZUk8mAlkPxVS+8PAb1Y8b+TqZhPUa3I
R69OzA/xVN/sCpZr3SrcWmtFUjE3fO11R6D3whb3DDt74dwecrs1k5TesfF6U9Rc
0tdSwKb+nm/klQ4tCHVrzw6Q7851t7NmvBeZzjTm/IUPv5fbH115LLtMsow3IiBs
Y7FsrLv4YwRtciIGnfQkPVpOwn8nth753cTZ+gRNcCliHc8eyeIiKbwM3EoGxMCE
FaVY6lNATQKDl05mYME/g9iKvWJi97DadXTC8yXiLCE=
`protect END_PROTECTED
