`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bm81CazkSGfbr+iv+eQWemKVxs1PJ7LnlHGYLTclbH5k+/YUViCjuP7rLSLBcK37
kJ+v86K61iuzzi7uH025sYjW6p+A/lqhKHgIkFN2YpvVUOYGXyIwogYKAjXFGJjF
LgqbvdCozWElyRk05bdhdk2T53FbATqTn2WJ1A6wAXzPLYiAMkLZhoVtBQhIg7lv
OlXNb8BAHdMNtYiFJTVzyesAbfH+Rzdtg/tX5/9/i5zcBNvacGAr/UYIB6yrGc+o
X404UMBzDmrPkbddeWvRkeWekiW005puUHFqZsMkWIdNtcj+kEMZz8Y1cqap63Gu
ymI0NodxRdqadBaGVoCy1Hz99d9xkpCBfeGjBi5HVeFcTwVos6h715GOOHHOnu7u
xUz3fgKX7v3dQzHsfbLoXBIBjHRksLXIO+LF+AYy7gJ1kBh4IM4sGTlz6QctJngX
YOnBWCjP1cM2xNn6qgxbomZipCp0uoKiE8HdtTkdS94oLi57oo5xHyFTyjW0pgao
WYcq6NbwWwlVqUafjdYua5L0rhRJD9wMY2StF9cVvB9yAejte8XIRwXShD/MMec7
xW3N16L0jVVu2bhUWqcCHw==
`protect END_PROTECTED
