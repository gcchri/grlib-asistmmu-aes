`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BA85BiY2tc4i4JfDHNKfWYW5OIYacoVlRYAb6Kk+wmD8Ga2OGimyHe3jFTSRcrya
76uFNl7zae+7lNU8/Aqqex6MqGjLD0wl42u/98dh7OlOqWuhbotRdmbJ3LgSFr8n
l/l7yYVQYrW82qWx9Lfo/Ij+RpAZteciTh2bblcT3lr9XpP1qQbKD54tvksB2s5W
ZVbQtvme8EdsegqXSob4QwnDGgleqtkjBbK10XI5K9m1QGrgIpfAdhslTtAavZ6e
84KINy6q0aMAzNc2o8vCHk71ronl8SqUcP6Ou0iVWFO7sfwuAD8DeYjBQe+NW8uN
Xw2c1ZUvqqXM6qMAjMYLPBJ5Jg8S9H5O754AtIDP604AhGI1e+ZzaeiwWSV6lW+B
rQe0lIAmWBPWlixmgGiZns+drwwq+5xmwvOTeM4SxQYES8UTJO3QIWZYbEISLnPg
yjS1HUSZPKaSh3swm6iN71Pgi/BpfcCWcMgd+7iTtburlRgNyaKrU/555FZ2qAbF
UUwjCD9A+2mdkGz7mbSqdgT3Bbfc/MALFBg0WHPKFZxop2En2L15YiDSVeCaC/gW
aoG6mNg1rMP2k1f3chnlAKQq5JqnbXDmwb/L9nyJ5CN6Yx9hmJn/PK4i0akM35wQ
JkdFjGVZpZbRIJGxvmsS0XXlIQasJjCXtVdU5AprOW81VqbCtnEZMP5kMMBe3B4F
xZGsmGOzTOAms8lJwtrxSYq/PgtVBc8oz4YQMhMbycdnsFnVXCeN1blxg2LzAkk6
EpKHgqCWANtkExRv1KCK44QFFC4ixarzV8AH0yE2h39vaj4neq3glavTFvAVgrRc
iZNJyC7LoAEq48qBKxsBckxBeGgALC0URPQKnektH+ZycOdE/U4angdstcrTJAz7
`protect END_PROTECTED
