`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kovivb6Hk+ASXKQ1TJPFRA2mkYhsVjeFSU+wu38m9s1TMBBYWQRExAPp9QeomKQR
cFTdKZ6j64QslMUsBRHNoKtWVW2tApeLlj4RNYZPTQ0dKaoRfGr+Mrv8XSt1dpd/
Eo2V9FDm49y0ASzu4x+2+IIQVgME5cUwiq1edyRGtaxwq3AZ/B6LgXSQc8SD2jOr
8S3qmaLN3qnLy5usRujBtK3UvvkFPdvKQDv1rP7dAnU4P0gRnMITaGnE4d/RwOZX
7NNc23wwkkcLIDj4G2vXNGJjrHuX1UpwtII7Of5R4yE=
`protect END_PROTECTED
