`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aSg15W+hoU2KMrkFbvIkWxd/gXi7r63uCuS1gRYufnD/8oV0wZoxPJ5d5FOWYEp7
umWj4fcbnBdzRCGzM+sKlkYgziH+67xABGNRMVgy/M6H9tBdrnKcyNwGO//pvb1j
e8sbhYnF2DmA/z1yVpBmfjnc8HYEXVj5scDowOSEnKQCw5HQbvpf5xkQM9+pJGfz
ivo3U0C0YonM7sVCMcs2DzTehBELly5oa3LjODg+T2Y/aQJ/oRY1XAGoIVjPUYeP
b7zC1kMPljYsivERwu4YwTWmcn3y7LbhsXa3FSgrd1kqrdWrCnI6gKR0xsHpZ1MZ
vdezjgFcK7d7yElCmxv6QPFyq7tTihNmz8vYeItMkzVLi+V1uwyFjQ6MnfvOODZD
pmF+OuVsGRPX7uKUhTph+L8/pZ+lIVH/0xOf0+/37Nnzn2QAy2jq0rlVqzDchO5V
Tv+DX0BHW77xu8UIUq2Xut1wJnlDiJpEu2hr8tNFSOqHibdN6sozqOLlP4PXh+GA
wSb2t0GnTQDEoIKL5ZlxvZqlp5BmS3BvPwUA8KKXQflxQgN6UMG6H6G/iiKtFWdB
gI2c8hXDeOk2RGmqQGQiNkXIGxBJmpd930m5Kv5X+9XgnFk3eo1lMOB5nxkbrtw1
B/JyjE5Wgdrviq2l7OvCxOqrPEvcD8g/9Jxtbm7LKcV1dDk6u4z6Girx3Ze2bMoo
Mla4ZLwsjT73Tzp7B6R0KZwlxeYSj/oHVI9voC0BJxSZ7X6zI/+EAUuAKvDrsk9d
`protect END_PROTECTED
