`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWNZLMjmCXPkN+AH8GGpYAoNalpXsRbpEm09H40zPGmF2Hq3ECo86SX52SUZpgsf
Lp4lyiDC7xRtHVjeME9ndEATXPU+9kBlYZsvYUDA4tj1FP1LMJkg6iDobzBUfitm
p/AvAxN1UedSb0Txr1TEj0hJPtOHTkNty+S3JFjbw4v/4ryMTncK8i+0OUAJgnZ3
cGqFLqDrrfRIPe/TWg1/wKjVmH1pHTAAD2tgTnET0CQZ0UzSyMr+gtY7Vw3mmdOS
FD2PJmtQEyyToSZxA8IUjHNX3FAxdTihhlFi7o/9hYqqmA2JIR6kci6rmgz+KckY
9ctPB0FL9+K+6pZdHrQdEQO2H+pJH7dTN0zxYlgAjqfpIuwX5to0839897MUHRas
b5ouYJQxVT5/Y/dZ58Yv6HF1hM3RjEtlvdaK3j5T9oJ+kAMagRfkymST/Z2wbv/A
r0t4cD9JuoC/O6bCFFjnbtoj3KAujjuin54tnlyDjOI=
`protect END_PROTECTED
