`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xlHoZzHpmY0qqmDqDWzvx221qQQOPqFwNoVPt1LQw4rQP5x14xBHSwXbe874GPft
kwDNPCkUFLIhl9zxQ+sIHi6CUwYZs2HmSSYx14iQV2FPG+blCVPFMcgZ+jAiUUQB
hgK4cUoY+I3ZOM5kJdxpqxJ1Ex0UCaCynwb6ImB5LG9pMv9BbK/spn43+cYUUjrO
amkCp6wU89F4t4qQjB0zQTBbZV5PD/gKhohS6mJEfZHN+k3/D8UBHN03QgsidsfO
DIMIkFPZrxCVNytCZljEozf1LkvvYhOIBEYYk4GPPxFuj/zwXQ2C724e9yfxVm/B
Ddkk1RPvs38Z+1jkydPMIL8bJ7/Ta7eedx1/vnRXVZgB5YTvp5QV0KyOKXK73uJH
NhGyZambsapb1zqgHjTh6ieyHl16b82FqPGnqLS0jxtGCNU+m9+PPT9du1DBw5UG
gzYlS+eIZkO6B3cAUXdEhUrODZPhR1GIgF8ogNJuBaT7yHsbTf+NNd1LL9uyndre
upv746yPoMDs+kjU8z7HgjvuQJdOpw9asVszD54yblbDBSi9NcAWPTUyfMPlTS0h
QIUt1NYF+Nxb5sSVESz2y1I0yN/WgTMgyHxSH13evi/ZHoDBdu7/uAuLUJKF5sM7
j63BH8kxnm/X2R7mx0eEVFooILkDvq1i57PLYADpq7XkegelzLjTH+fhSjF1hppC
O+ZzbBQXyVw0Dq7PsuUTg1+KUGimgIa11PvcgpvKVSvzrcjzGqXDqppzzIr8BE2P
rjXcs/W0WnN/Q5Z7idVSuQ==
`protect END_PROTECTED
