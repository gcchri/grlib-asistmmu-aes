`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1fWP6irMY3KOR4EpMLIj25njCo+7ym99TG8F2e80Int4Rq0myiEAYMVsigpw6fT
Nzhnf4ZfTNULOIkXpRZG653yhNDzTdmdlHGc54iLkNwddc+jOee4mXCq55aK/+oD
FYvSghlBWFFzB5fzAgmlaT4oqXYjn9j3MP6zxS5MbKJ9MYnMwaYHlkmkgEGZNdvF
xVTuu//T5XCdjXEuOhqTUkKgWLZmJhtHQPOjDm+rQjbeMnzfJjTCKNaROt7vlcAg
cuubZnZ/MO8j+ludIX8MHvzBaAbgg8kG3A2Y9JVHZf+1+VwiJzHOmw3Yy7iHJB6P
+OKYxvVP5zQTnGqlWhZFamsew7qB9Nq9UWnxHOZglfhAQZ1MQOv7OoRLdJEjsaAV
9mBolu44nWQo5UtLD4uJhEntkBe5l9gZCUgiDQYLbaLpzKFL8wcsHiLSLj7NfE+i
b81cOYpmtBpjKwU8ztOTpakIHfbXUUmFqzB1fgktrW7KGNvmDMMLa3zNEBczqF12
VnriVO9eQxkdw7004lKW1Sv6APCbh/g1Zy5Gy6au1ZadCIl0m7lJYv+9NoEqMdBJ
irzV2CFMmpUUx2gKqh3tnaxs8GqDmSMl+/UqqX0zG0pelvWW0vBxnbjL7RdQp2bJ
tXZ3p9+bGEVaTRQzmTQok5wE8Bz6O33/Lrqpbwkg/0SXSZ4oq10WO42Da4quli7v
`protect END_PROTECTED
