`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
leuRbyYKNuP4avnC67AR/HwOSZ/4bu0ohZzVyUpNOJxvJCugDDeoKbTTSEcLG/J5
JKRXoV9ewrwivFqrLJn32g24HkQONsphFfc7eKPPYih7mplfuH9u8oCkf/Yf8EKl
nGuFskK7c2O+kKoAqcYhfqVYaAb5krGmnjQdTfeE0Ci95Bpmu1QPMFqjAI1/IhMt
deR0tvf5KHFCZaoJF0heri0oGs5fMMxux8pcialBkov5ZkV1kBhO1x5VaYSMhvO2
YWshoV630pAxWVRHCoz/7yoIS5M/gMtnGwWSTRejdq0znchKr/OhXiaHqsIzpqIL
n05sR8pc06l+7FoUjEd7dcbGwYwW7UcySPgH9kljKsL7z86L3oRnbqAgPqlPGs5w
P0uBXtiBXADyfHQZIM16BN8r/lc00ZNSsjTT8cZcBZShcI6WBEPy246pgKfw/SbK
Epf4ea7o8I3dZ0Xddnuhw8Y73F6edOH4Kin6ow1UTExNOn40asPA15YOeg1VvDWd
2jp43ajkrjXCPIoyrasdMygTqu66iOb7YU9PnEdVmwvFQnhPve+lnIKFSGCa6gfr
MbjzbS/LpCbmEbPpRNiGP9D3MMEDEslpr+kPIGrVITd04oFiBizVckA0bl4ZSXU/
FutO855Y8asIWU5PeOdkrOkUr3bwCIkUKYt0+jvBGHvfxFrPQoTXun0XyzjGBEB3
kS38OPKPSaReNhurWJVvB61Zt0WZ5IjHsDuh9oSzw0T4UvJB9JkwK0Fxxdl7G1SW
qcOREbx16Pvsy9W2iJKN+V/1ROeJWsv3JAKnSaDt5h01/LIX9bT9wLZYMI/k83Et
qwbtMRDCxnLjBOZCKpfNFMvxOYsi/InS1O4n8kxmdRn1Vo4fWo+APRkir2+3OQgy
Zv8sR/6B8gO/EFnYh/lDX+gCXBTt0TIoBak8lH4/P1DM0T3UCfG0K0xR4KLPIGDL
7hUqpw4vTg6ab5iaoLHyi8OQD32cU6Rv++umjJo3S8XDBCXyrJT06QGdNC6yWGfh
Bd7gBxNHEdMc5hpM2i1yc24rO7J3TIOtninOk873SlExT/10+XsaD+YsY5PUwSjJ
iRu1a5iasL4Ixs0rxufiOr2WYMZtrXOCxUDxQr4QryNwF4ILSGNeVUoRatQ1N3zV
BqJQyfCh+6Os5dQ5g/SyWjx37NWuPnlAd37f8di5H5S8UVrpTWpB+ybQSGzB97e1
hpPleuODb+m3XMN521MYak4FfIl4PI2FozFDSNZMLKlUaf0BJQSUsx0emP7W0CXe
Js+Nn2zMbveDG7L7gmQUFH2xIuj27JRWGY7F0pAjlpu1lOPkKwkshipN5d7zVvHu
aPLmW0iQNJYktI2V7v85dqU8VxxiH7TN6OwoFPKzAK6wDbtylYLPZXlBXJWB8dAX
7b6XyyFzi1+Cf3ishTlYDenHNbY9qQj9tbX52f2ms2iJwZt7wDFwdZWyF+XRglLf
5ith2m1Pt7w0iuR05x6MfDWgJZIBNEcakODdwCvjMMGaHGHNakpqW+KEeY6TOA7v
PKavZcoEf85cehe76CjmYsFTuR1YI44smaeT4EVwGNrmRzDonI/dR838BR+XvK87
OTOW95CG0zLdtGPxrKTosFoKUiXyEw5Kxulw2jNyNv4JnTpXcKTEwf1TaLNqEEpK
LxGwWejoI18fvGX6g5gxfAbZvKTEzeeJBELl++9eBHcezeM1+i2qMZJLcrWxY6b8
I6e3PNhDrfZVLnoaWsGUWp9M+9JfXQJraYVItvBRgMuaHaaqY2HuXFa9M2eN6Xwi
RFIydoB2W9PPWKiw/O5zoPu8GvRw1Tjhtpxd5sBSqQoh573xLQz/PMSAYiR3SIE1
UPffPWX2/sPC+M0kBQGj56XcpJFJzcfqHIHfKa7RTRKL7o2iCibHooGcEaFGVQ3b
qlkBD3kxuFYyButuKsb12praWSn2sWDKgX+V7FEFvesvN8Zjs2N7IG5+x7WYhxhb
ywm5zJgB+sYb2KPzYV7KRu/PhNXxkELNC00jFaZrYWCVZfllBswYBsphIOqBYzx4
kad0ZMgkUBV5rSB5x/0bcPOLe5ktc4K+PtOAjeoQ3rYozvXv5kdSz4OMfa4a+Xjv
zB80v912tkt1kcudHQat643ZF6HOm+z4fqeE9ScSGPwXGtLiG/y9B2qY8/DVaAEb
IBTMHKM3F0OoymGcLmrMtkQRSDmnQlPlqe5ukpC8En0sNadWO3M0kkK3DXRsNgAW
kdhADfKWSgYvODFRQ4+zTX8bfvE9sgP7Taah2GVkiUeBmNcBP5Is5cNbcmP71ufr
T2JzDlJvZW+nhF6W6wHyaJBuWgNccxlQM/xK6FspqkwF2CAuBrlKiZG1FSmD9lp1
+GeCbylFXz8LhZjTblrZ3Eh2ef8jbNh6kcIuwWiF5CzQh0J2c9ZfklqhU7v6BCaR
1+NC+EZzK5rqRAqYHIDDrK91D/tfcK62+CGYukHacgp6lWS3SEveHM7ymDxrudGx
h8nj0Hm7y+twsvQgoPlnencRjRK10it4WDMoqhFhtEU8oida/4M1/dzh5hqwTj+X
DoRxbt36+rHUk/kgOb2HR2tSq/bxiA50zssTxSaqbWP/NColbB2d63g98u2Y6Ice
sQpN/pk5bHyHwKlBATdxnrJ+9qcNkJwIymjJUQUCbvO1BQyI3wsBh9UhWL9FdYUq
eIgvVQBng3fwKFQwi2Og3I/4sUMbchqoEfbVjtPLemr2UMsNODIwiqgXzTSmEJen
xXt5jw+vKaRxzTt7iDKKG+s5QfwSncL0V4NrISPKam5EQ1hVRZv8Qzjb1bVjD6S/
kGwAIJkRu1YbceeMVS8KIn3ze0kRS6DxToZMBW7PhKE7pM7KQasQ1DXEmrQ3CdQT
S+wzwDQUfhSlyztA1kW/NTWffLtM3yLlVdIT0V2zUlXfoAo/ZBub/cVl8M3qavXX
iaKiv5GPvg44SxqPyfLG2jIcrfSKLF2Ec7Z/OlAm3Ri9UJG5F9fH5aF2ToGmwchc
W/48kxaN5jriqGbZDNqwXRD1dtCuoTjaIiC29RiAvtlJDaEBI6argmUwz9MHwcrc
UkeX6rGHZKCaXl6XcZn/4bAp8+HZvc5RydJuoEBiqMOG6FzCRkZRXHGwRVr7l7Bz
nIBDX+xZkCFZVIdCWUPbGjaDrhjnL2jiNBz5nMLVZBN/wRvbv0UbivripKcx2FOs
lbE6gX6KvhT23lgE+TOn9wF4r3zsINy/mQpTzyMFuo1s5Otj94TCiGUSE4UQHTAf
4TOJ+1f8xhhEyFHhQmyt8duAcFHlffMsAeGoDwnh3ZccmYjiEye7u4/YHklKv8xW
B0eZJ4Vxnk2QdqIuanuyvaY3RFNRsAmLdPtCU4YPb51jMNHmzKptJRY7qd5DSpI1
JZeWUbVYs+OXMxs/r4eCE/ncYOXXY3zgd+uCfLOnWa0UwTJDwtKlcCZ6kXeeYzEx
a0FwVaCKEnAPQRpntF8qRtCDcaPk8bKk+QdsD+TRp5Oe7xFepvt2Sv8UhF3OdfvJ
ZNSn1eyM7r6eFEIin8iJl9BlbotmJoeE6MbsiOljx8puJSfA+vT+OvFsYFJXeo48
9UU1zIdqCp5tYjQ0IqA7qgAVjxJiq/28n65Rw5tsufi4IMgpaECURTenKjWojJdK
KGt2bvkBfqyL8WLm6bjA1m4Xxy8h3r5nhbCPKuFNX1RkyU80rVU4/h8AKXmcuZi9
Y8bO9VFHPRL8upMfiiKcxknKGP7DmItKM8EZ5Q3gms6VAmGnt7FkFuZ5CqEHyYac
T/7YytYTJoYLCa7WyD29aPevap4DBU1OSYQGxhy8uUwfoE3EdlUhW/djmqqBCEmN
o4nIkdFmrLvRLFBfWyG1+8eYNKaLqmIabjZhB0oUnxSJxI5ALZMcMBy5m3sT10ks
a+gxhFYw42coKlBXQAMeeNrwIteYBPTVCL6EvKu1/Kr6LK+mwftkdVf4oURooK7J
zUpN6PmBDSfNB6djZ8Kib1OVxzanseGX5zu+tIR+ipFMShoINk6sTyn2ZQFslLhi
FxIlv5taFuzYLhTeszioEmaGT3IW0UDixNy2lT4b3L6SojGt9jj+NCFJP/raXTQr
5/MEdDZooVdnzPs9s2WaljDGHVhpWXNnm+J8SpPuqtgiIoQr5Yv3m7UDf06FXfs0
52gEmnCHHfwaFr4iaAbFoTU3nsw0jUI0t9tYEZjRn8ai9XZdNnnqOTOqe8IiTw6t
mdSPayVLisKYnCTrNG1v94ygatgpgWvjqlETNy8KTV0TF1kVFQqctM8TuFgFibCH
3oNZICQd7J/Vi/ufSxzmklpU5e5Q168SgZ05R6FFYh7UlU1jQt3vuKvlVk7kJh2u
jRDBCJDrcos8ZpHMJ8ys+rRBrWTMVS+VPDDjolEV27ZXKq3toDbQVH+BpkohVy40
Mm7LQAdicwnr6EFU5K2Mbbtm5z4WpD+cBO/NXSDKqezKBlBc8HSlTP5SlbOFw5y0
gaFUL5BqvnVa7iIyzmYI2jAhPfSAcfwqoBlwHXk7UdCVIKGD8JFamEdAs48/Mhw5
3P0Kb/S/z9XkqQ+s19r8UOu6UOQFp/nJPVf47VJZkL1sBkaICNo8yowrUHmcmpF5
Ie7IIl647TzxDhF1E+S/tJp/KKI9Xj1hyoXus3CsEOze6LgRSMZXTYKsU4B/+F76
95KbglYABpI05Wu/aBO9MQX7wnD7zVtfR3itwnhDsWyC+r6tRAZyspbktAbaRF/Z
ffXlN0MKRALulkIDN47tDqv2TVFG8bfQ8GWDjf4Mtt2b2aSCq2bUsQwIzxHUsV21
F/3rAoetLzDkW7mHvJHZKLMLqFZm/mzJllWTL0P/QQNYa2BdX00XeS4YwZNZ+Lru
B7nX9FP/Mlp2NjSusMxnSwwLerH2Ro+velL9JK7nIj5t8VMFmQK+lcLp1z/OeVJh
4Flu8tyQmd42yH2YIi1SRlv3cBGZ9nLFG4HhfKhIW2J/xUOzL3lImai7lJlWG9kD
zXBHZXyrch1/uRf1sOaceghx7kLiNe7gvkeKHsfdipAcqtmBR2+BzZPesN6iL+TZ
r63fLYpJ5+dYlWw9KDF0NxXm9csooTcLwdMZXRs/ujODUCfQuC11HTNCBr9yXA4W
JEnkFnBdjgCFBMfAEUKfKkwwSuuj2dh9Bwiyo88iKPkoB9opJ4eSYnStrtofBSCx
VekhcSFZgLGxYHoXK1pBT/BLEtiJU4tSKTMqQfHb59jUFybZTJkRVjM6HVaZ94oQ
IoqQoZJ6u/OynijgA2hgnvTezdkCdAC1cydzBVckYhbRJSbfJs25C71rQkA4Yl1a
MjdQDnLh/6bKyLMgjh/ulVNpV49Ka4WIiZ9+TUi7ZjWCl9ukqH119KEmb+4KVZYy
4UQCfGoYD2Goj0Avq+0nEImJ8rQHoB81MUI/Qv4vu+uo7jDoEIIJY5OAdbOdUUNp
sy2WMqQxsOkaRKGuhkJYNAlGfGsI2ukOPGx8FwuOcGT3Ra7PIakoYgvIHaelMff1
/g8vyVLAgJsrnEKwnsfw/KdIy8j8qn2RO/vyviB11VotcpmsjRqi10yW0ETSMS0A
SiZOGuOLF6xBwCsVPtprfDxCmAS9lZToPOpvRM1VsW6dusl4BtoSi6xpZ8JMQoQt
XrZ3c3c9MLIpvstc1aYZxRmv6XYEsclVJrIgdtuPI8RKWQtkyoh/hkUiPV/NyTKJ
b+If/IKPeO018ZTZInd27DE1BqGm8gCRAke4Ioxi8ZHoBn+/18RbBjvoHnws6oBB
0R0WwMf2x227C7WiIyvSSFw1IODQ/0wsb/oKU/8K8q81C37VHYXx+UdTp0Ch2zRR
wlMBeuAda3x4NGy50awqT3g//fimoZy0of94QzT8eOFEPnjp9awt3NQY5+EJgK4d
VxLM+F2XsoiiWDUltkMSafH1CV4T27ac/8JdfN6IpybUIQVddy9o8GL4dzpnlqpq
IHT3cUGm+oHwgQ4DfpIIXghoXTCVP6hwxKsP/NI74Ivt5GuVVEafPX4BUYmGkdq+
59c6+DVpC5YXUMKyCznbSf8y6mTWpX3YgCjjqw7KlHmQoplfc/AoBDB5yPo+hve3
7sDhwHELppET3MwoKqq6rG0KdAjqrxNr1Rob8hMXJ8IUmuVqMJ1B1zInDwAQNCZP
mVjX1z6o8PSi+Qh4QP5rJfZ9GDHOvG2p2CigUu68nJ+RYwGL5l40lo8LiecRkagi
X0HQcUhils5IYHNUDKQimBNhwK3aL1Qx28UmQeGABJ+mLjDXS7IjWwkRyoE+GWyq
EQmtOg+DWWhA5D9EauuJ31cQ1PIKjKjga2RiViGZyHyA+6toGc2nVgpYjHaASZNu
x89xCPiTjkVsem6JtnhonhXCJxOKaN03+HF75Qju4ucqHWPDDhDq6LZZBDMk+qXn
hJEyIt2RSQU4hEpw1ZN3MMytT1mms8XM4HAcENo/9Oj4Aa8zoawEqyp8UCWugE+f
fSPmCENCEzgKXedGry11Qp9HovNSJpAPoZQshfn2lzg5u7TauezCa7PLdtgvB+hX
TM57kUFMJLAZe5NOx6LevLUMdoC0yupl61z3kmn5z8RClLy+HHsQ3CEEvsruUTI1
kn3IGpGmG5WSetjIhM+SXL4MOE/tdC7EnANnDd5CaerLmVRMFg/rs+7MpxE3LYcR
7NGN+Df+nxXV1N0BMP19/pZnc3wh3FvBOB6N+rpkxjFVo/kU4uRRZkjjrflmu/tC
zQsuFvqJtkvqMSsQIHkfjLkjYI30m80MzUM7GAfGi1W+14GE74HHRubg3k4yGFZo
M9FjIKp+Vev4H+S5F4n2Bnd0mjyfZCr71Hh108rBReybKC7xetgIhDZ+OPb3evfz
B2K91VfX0uUa8bvhP3vw66kAnXph7hTrz1iK2tnZ5IEFrnQwn+AosFfcw+m9Lmeu
toP5HcJYRGvcW4FLwbxthKbKdt0hFFiI4uAYZBKuZogWp8Dl/PrldhYpcL9DZGdp
IhdHauW/konondIxijOjzwa7JCitZPzSl/xYuDat9aCh0yx9ljNRWNyR6E/KmwYX
D8mO1s8FJgCpv8BlcEk7j6+/jByoWRwLkx9unZ9gtntc8dxVsVCTc1gZ7qNu0FG2
QlWgLsFmpIxryesQHMG7C+XfGCGPqnXEBCkeM8G7oHR1bJmiEl38bhQ7CqbTzhvZ
XSOydLi7VrU4EWk7tR9ncGC7IYNIKEh/TNfjoaiV0Qiw6r2LyY/Q2UvSI80Mpczt
qf4Hw9NnDqWSyqlN1+phf3yExREQStEm1FHBF0SK0Z4g1OYAGEvr0J6/WzANA/kg
tyjnr1r1IYDxuCD02EgWUgn1cNXxOjuvC0bWpFz2J5EczUCsMrYJ9H8bx7cYO+e9
yO5AF0c3XSCqR7WBcd7QFNxh50pjt/1ztE/yMz5wSzd0mfyHgqHE+n6N3e1fDn//
pNdp9oDidvjLdJ2IEG25SrFjcU/Oeuo4t4lCgrK4b6gczEnE1KvZgECnXjPlDTpy
6VTP17dB1svUq49yj0sHIiQfvxMgZa3J6rSoE6zimrGYVYGoYz/J+UQ9j1ulROXw
cVbRpAvmnLKFJUtgS2FbMgErlCk/gO6NkYooMQboWtBaziUmuJMamck5DB12b4uz
gfKlgikTA1LGnTIarT/yXu7Sa7r97P0LQ7cN/0iwMvcQOoL63qQ4yGg7WuMgimCt
LQ4EMAZNroWc65JC0U/UDtwdtKBVK8mdqYv1+7HMAaSz1j70zsAuUCozg7qi2Ak0
6dYvHt10PMNkCtstxBi9YA6oc55Wu/JQhKdubypkRfXSV6YASlPCFOPBSH2xYUdl
22+sXN2/xA9KxJF79RkGLdE8GUdlFT43SfDi1LuxxTVbt6Hv/GiyUHzCxErguWeB
LX9ACFvKwP/CeZNu724d0wNGx5+sm0677Jl+az0qMxIDSLg2DJANGWaLKaEj4Fiy
qgOjo687BOMpKrXG9z9wvm5WW2VLL00bag7g5iVifptkDXM896QMgJKZAlwoadA1
7TcmZw184Kq46rtNl8p+Lud0cl0+egDlG655+5CIXs2buejqU5VdiGFgqsXWBMKk
jaZz3tt5JU8IxEbraEH11gXWaubH/vxlvK1huR8ACWWGsMU1lUkEpsUtWxOCtIpc
HpKV1BC9XxE31mFriWtTQ80Hv359CshwDy59W/K2f7KWdFn0JMAqpnVxvVFsCoYV
+WtbnyF9nTiJ9w2TwnxM+mvEu6NyWfQe9w4WIORtT2I+rxwQzCGq75BXgHldCSgg
c0BpQPGYNYG5I6Vhsqe2u/ohz1vtk3MStE2GGWhlZbs/E4Z2ddoSOoImPcEffoQc
H5h1OBAnevA81fskD6Hyf9/FY5Kup2egt1oc5EvPs3gc8sMBRJPXqJMzNXak62wu
Nya3T1sjI0LfcME4ESXS467CBRd9hZMX1G4iMZGHShghgec9cU7NpeANUf5OsEEm
6BZO3q/MkD72IgQb5cR0vnsAA09HhUDTua0eellJkRruJtayc3P1LqeN1QKTVcfI
mL9eqloBEdZzEGohL8CXXMonMhDOO9vr6kPAUQCBbEBURlz1Nz5Eh5QXwvO3hGSp
FY8A2r4MAxvde8j8qZGjbRYp6Yo/KMQjnY8xZqJGE/E8IJ93/A7V9IZ2lAqL1zHt
elDr+iJMIE8qE2f6FL/ClZm6bbFR1Ko3Phjd2l+lqsBmFZND+Rr8zzPIzdrVI1k1
L0mDcYTaqaahCZdyDEo21nOfqlUh/vRvv5ojLK3ysIGbX5b5JECPy1LDM6Y+992U
9pf5jfTZPlE+45GtBmX2szPhkhp9FrIj+WZEZYNlDZGMIX8zkMzDDZ7QaI86ag0B
dhEULXenguuPWUpwDPR78+x4SpEPOdbRtleV7R8mQtw82B2uk577mIjS42II0dru
kzGYnnUsgxDdqSOWcGgRrjaouHMA0AylntEUebAA3EUjapuU10p41BvJnM7F0rxp
KCqQBrS+2I5TzR7nQg21j/oxiCd03kxUnX+vtoxzmPxjVti0sste4NpT3GmnWEgn
sdKq64HP5IlOkylnHUUgeeW8A5+HFyuF/Yk3rrBrtbtlR1R4/cwB9goc2KInVwxC
kE6CDDAREFsUMVyEf+3d2Evuuvbl1fmvCznm49aOeQAve9E1TFEwv2HYqja3C8MF
GnUWEJ9x/9o6cLxjMds6AioTBJjgA8s9hXqMgafmE1VmY1XuMYhjyn6dIlmh5600
FcgFz4B+z/eX0tH+IXFNgN2ltc9arB917IchFKZ3mkN0+eiCpdVwFvUKP1rxFUZG
pMiIcpPCLt3icoQI4S46TIGek/K9Fe2V8My7LX7ISWWwMUhTI6Q48h3GWIL9pJSd
2dlpAgXf4ESUkvS66hQJS8aI5BAmvQnzZNatvgd0+f1X6Eoqw62Hg8VZ8Pa3WT5V
d0ungcUSgRNnEvZm/Tq9MP33ttw4bV2ZL5L/MeCydf/pBXQLH3jeWFmHwk4g4WVb
vj+lUSze3mXg14YTjrztA6rfZj6Z9X8/xyUvVlPTK6ol7nB4jQhtSuvyr1H4NBsh
BxzQw2bzEb2Ze1cJO+XXYeWyQUkwUh1qjy/VWAM3f5Exwg6xsmAvCo3GLHmSX+Sm
OUmtTVw61rD+N91d5fxtsfJek2gjBp9/xRPXFGN1IEvDM6AlXQw/5/ccbmmkLwJ+
Saekqeu2+JTXrtvhkWmGV0BKbaVtP1QYq4w87fvM3zDMA87wabCNv5jex/Gq+e6r
FxgWbmjfptPEiE2pHV4fTxYcdi4Ou+GApCWKjFQ1yuyRn57Zy67CraI0rvo95v3U
5Z2Ty0RL4KD2bSZSBXoRIWa12BvP1D4ueokkq9cq9SMLoY3n6+M3uBTJA27Bz9xk
zVhPpsF0d5o2YzdfIMgGg5BTgiSUOeMNqIHoI7Ur8F/bVj4vYGHKC7S4LUlKiRE3
siBsx/zkhczN2QtB3tqC9gBHLE2r8uWj37GJGKcUrDiUWgb6qifkGQ+C82pK+TRu
Ur8IXMOCMreGCiTrgeOmV11Iiz1gAApFtcl7dG52+aMbNWRp3yeu2mynIzwmuJHU
oI7xnAljm9jLD7Liu13AuRopsYn9BygV3gaqWzObb+kXCTj3HZereOHJD0Pvtvzo
GMkm5shqVmf4hlRuAa4MnQ==
`protect END_PROTECTED
