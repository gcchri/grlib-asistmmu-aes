`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jeADF4TBGZyj774jU8zpSRDnmqLEbTjdmwa5nxAdr9XVyLHIqCFU0IqzjXCGrYFl
0H6mgIIacM+fSI6JHNJI6VPWYyCprbu3W23BNUavqAisYUZbZ8Ll33gTjODWs4Q1
MK19Y9s1CaMe8keFlDQV0dQKyT/RVmtzM43jfmL6eg3yKQ5GKhJJ+o/snGoZiyU+
tKdSq0cXOQ9NMIfaBJbVppeNQD5O5/U2huLXw1ck4QFyokiOt9iTNsrAYunyS5XY
kSI0pyegkzjRrFdVwefO8A==
`protect END_PROTECTED
