`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bKBKQOVbhZBdsnzS/0PBOAMrIkgLWLsHhqnebyTMU1tEdMHdp2TWsRjUbD3wey0i
okl03tnblwvI5l9uGuNvr2+u2+uhGIiF1ATI95N0TE10i9mq05m6QyaIJLdoMIXf
86pBrGncWrR8oQ/prWPconxpq9xtckPBC7eEyodo/lixmGEGx/cyiVqkz33aN0ms
o5VbRwvlCIWLkQx+3yO5Z0vFTyv4pUASIwOKFth/7O2REIsWwVQJAF49sPDGRLVZ
a/vdHLkkE2IOowxi29VuBm3JPsQ37qgIasF13m1VKE3NJwSBCzX4YzXO9rRiQDtE
a8l1u0GK0aPISqGeLG3D61JylCwQAaZs9F4YsUpTtBofrHT8/pH38sivEuZrTCXw
FPhQVj+qfBm2mbo8Ijze4Su8LVra2YwOckgLv6zHe7yUt6inrQEx0eeplD1o1RCb
9ShUSPYbQyDl47R9JLt3vG9RGjUDqXTHiUwbU6t4pTAdV01v/qxWWpTayXT+JxvB
bsolTyBdTjPx5S6SnU84UAjim9ku760EAEvTvc65Dq4Ak92tQKSgSO6TRVc2ybKR
BCfJ4YXmvIRDsMq0Ad0nnd/5WKUKuv9jrBhUVEnGikP/VpHwapvIdSnl18sqp6f5
LukqpnpmOT93tjAI1cIcxI4ja+EOzw3Ih5w1EERiuog1DJbZu9EvFXQAurG9jav1
DVD93yg7NG99vr6JVGaQykIwa+CYigUsTjr8awORan/ceLQkDk1VN5C4adyjuREH
KeBNYPtw4JJBanAqSW/6FFyrglIWuPnjZuFJPMFhUxBQ/j9IwQZNTkmccRRtifvD
n5xJfIsZrWwNoC61AMxWHA==
`protect END_PROTECTED
