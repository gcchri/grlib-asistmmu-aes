`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pljDL8EA0olKMSrnEcQNPc4Gdt74H+JUWBw/iLSrYBY1b3U9zQDzz3uIC9P1NC13
Herlx7/l57KjQGaNjaGeObPv4yYtbiqdnLzaUrcCy6aSymY0ea+Op4r5gHF6s+wF
Bo3luesqltT0arRxhB3n93DGHo/qK6ZiZnxSbo7p3Ch+dyA0fgghRTpdGYqN81nJ
3oWWRpzZDDa4kTgCHuf5K2N0oawbphn/FwaaL0HezRogXqCvbfeuFS7eAEEsEtpT
GeFoNX7zvXVCkiZNgaBPWA==
`protect END_PROTECTED
