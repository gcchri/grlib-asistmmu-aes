`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SCafxg8SlSWyY9ym6yvs6t3WeOcnacX23qAnH50AbUyfDZFUR84FmsUoGQFHCxT3
/09wnW6m6/OmIiLXAuisB4U//RUnGNj7IigjVw1s87fLPnvXYBrIpnzhakDdGi1l
LiNJcY6CjiREz4h6hUY5tUmyuy+GENZ2fom9lAZH0KmSlr66R1Z5WmM/WiV1icM9
ngk1mJRvpfPn6CeG6F2nb8x5kAXB8Gp0sbbnM/YXJ0kUOCwKxxHTXxjWSEmoYgfY
NYw4i2jvvNyAoxRyjldF7ql0j61D4VQnU7wJPSsRXPlIBrR7HQ3/fHa08cG5HCRw
DCXpLqnpSUbBGyc4KIor7HAZlTqP6QMMwoQtZNlNX++Jt6ADFsIBTf2jIRHioLwJ
hZ0Lpp3//jLrMIgWTv85xQSAFWX6aXB8mjoIyIJpfGKFtyWt/p+/FBbZxANCC8hX
DHpONsY6su3VokBYUuUmRnfE+f2Ignxv6m1UqUvIU0jVtMXWw8mkTE4IniPP+IJK
2TQO9al9MjwFVxhJr3QYk22vFaN8TX3wn9LOp+pC/DVfXcHT7R8Ak7admW8dIR90
cx78qyxVz7nKn2htRePiQqK20L0fWpF6k6Pts7kBo5IqBSkYbMZtS1h7EWmhvBUc
e//3BXZMGqzGxdpcswHJIw==
`protect END_PROTECTED
