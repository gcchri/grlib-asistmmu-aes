`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFnw7H4z7XdH83FIxjKslghdP5kfP83vE7DTdrZQMiRCs2Uk+aqWNXYdILFaM9kt
tF332OIzzTmAZIQ9Tn2H1aQYRUaLFGN6IJ0V9AUHLtC+cUt0AIBPtbjbxFi78HwA
Fvw/PK45JL53JCIxx4UfOugNFixFSa49n+h77AKN822weAEOr+W9VpqkUy10jwUf
GB7SVTRSPPkmuY4D0Z0QkNFMsGd5wLe6fOVhQpPgYNWWBEMZEIDt75IEcgMpSAwX
aueNPm22S3Ephrk/PthokQs9yCuBlXzRSvSQ+kKmfwtgimI7+/sS8DUg9OXA69FN
Eq5OLPdcF2/mN/aqtnJu7IRtA9AzyiJn0dMEfxqQSFUIPTL8wkIFEqH9ya6vA1Pc
2nrXj647pC9D7zz06V27oziSvp+ZZ3bldluq1aI68dlMOjN3Jec0O36uxNvUyMaf
WoTkQ754/N043R7oWE/RprQ/mNnP6PeChVUszCZknrA=
`protect END_PROTECTED
