`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9XkhlQr8UvycxXBmGAe/2kNrJ+nJtXThQVpz/ofr0yeC/Ow8blCNonP6i/LOWy1i
J1P8+60jqqPhMC1ksKYXo1qN6qZiVbl/QxVzwwwW4vDRKyY8txwpAq9sJYjoWzAk
KeSF/aV6b2hXtah5UORs1FJHZTvU8mXHSSlK5K9kuchMij9hmCI3hAPn5Bq+KshX
DXqxoT52Ea10OqvcMUNH95uFXL3UEOe7hgoZJltZjy9RB0/rRXuAlZdxxIEzEaMu
aoB5r8wsu0qO3svlAltu/KzKV+a/3W0zgE1XtjgdqqXZ5SXvP/eMCgyD2JLUpJro
RAa0+3wOeUvYmIv3Jao6Ix+aHdOvJPZVUFr3MNbdJAoiP72pCamHk+zlcB1ERGAm
8ETPA8H9kX6cJEMgtj9u5vXLW+UDV5HOPZ4O4GUcnnXihxsCw4yMaz5C2iaTwwNp
`protect END_PROTECTED
