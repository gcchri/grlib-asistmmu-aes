`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iLNLrTEgMC+4kzz1JuevmjDrmXnbiviL1O5Fdd92qR/ElTXq4ddwizlV9uKg8Vtr
WAQZ5wrxyri7q2q+rZS2Rklq0RVcVXBjKqmnuZ8DEi9z6dAHeG2xcwUr/Xa+J8Iz
rhTI+21yMfnaE7qTzxS/wME6f+KOMjbgqeZ2QWVljOC5beS+s8gtd5aWPvbQCZKK
qbuLwNdjBKpKTieIjwRnibscr3ZvFI9doLCHiLt3LSvZ/zHjtcEZmHW70VqoD1KL
LgTfYnXtP8w6Qxvsq9SKSI6MDWkM+iA8znJkl/u8yRgFlFTUIJ4zlqzYe5do6qq9
dD3a2+TeBdX+DNGDYTYMLKRdXQCql7XUPI78ngBx91DHo7/qLjnKSEP5KY9oaPd8
8GYurIwFO+6hmNvJYzK8VBztuROhYhgvVEKHRsdnDzd9pytW0tEw94+vQt2OvZEX
a+gZoc1wnlIp3VZ2C/YBfgxatGwWB3MaUYNVdStmGSI=
`protect END_PROTECTED
