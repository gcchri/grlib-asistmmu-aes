`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2NIiX502KIOBrQOVDjWuAsUuJqyBmKnRpnxeliQCheGCn8rg/z1yWrbC3uxLEKhU
qbNFKC245+PqkmZLV5JFn7eYOgflpLh1AINdK+MQbaRV0YdkO9F7KXjMXV3Ok66P
jVfZEv08AY2QLSlD3rxntrynMl7WIiboTR8PQB1Pk/xp49CMBnXUtSSwNrug3pbA
H4F4NMWhXjIFRA68TYh6lOsbslB7h+CUXaVp16TZz4/BXm54NFadK0hCOv7iyj7i
Qf2AtRgHMBFykZe2nGoml/kHYZ2C3s+nS7OeIDV8ZVL7ME/cJ6bCuW3ULmQ+/n1o
Xu/Q3vVAGNvvJgpgk1/9FT9B9BytYUXLsIP5HHFyh/0d67xsETGQiThJULEikL1h
lm7X2ZgT0zIt4GjWxS2+uHxIG/aoYJefb4OZSsPQdfEdmQ6kjhsO0mkgx711To/u
iUqaeAFGAE49UmNyCt48cr63Xt6YiyuHAbqv5MCywURJ+/Hw4j2G14dVTuuJEexM
Qw7AW6016ADBeq7pQVKvSV7+6gvlOCa0u+IoTnu4lPaUHeQVLmSncM0VXkfY/pvU
rabax8YRuV+MCaib4gs/tAcPCrxX4DbWqY0kY7PK1vNX83SarHLGcX2acdbhcaQA
zj9ltWtiqFU95v/7skZKzn2ecScEeyPz1y4jVOT+QIfixkHv7bKsCgJ+Bj0USETP
R1OHzMtgEr4sx5Cyr0o2aCWIx9XoDmdz7TaNiTfsQjY=
`protect END_PROTECTED
