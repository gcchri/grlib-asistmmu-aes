`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wetcj63YBDztEJ4VIN9Acn06FnMJ9t2NHRd79julANQilAV/vTt90hWZB4AKYAz1
dH84aYX9xlEmqPP6D0NrQ9ANcQcAFAYH+qZ48YHD5h4RLoydIOBNdG3cO5dliHCf
n5g5DgXh6NIaMmC5gFT7YkreYXZgrY3GDMdFFozU58V7MIAT7vS53hm8DmucOE9t
L29Rr4R27gf06yLMgFl+4RT78b90B+pP+bOY4EBk3tC9PgfOnMwhhAr6jkT68ufg
eXaHP8MonVBg/+V2lYqoWPY4842ZC0x5g0+ee1eaKkusTclsatdT4Btm6Gkyq1Eg
fpXdz1QzkBSbaukv5BAYRUTUIFw2KM753n8ji8GSw1GnQgXQNMoZVbYn/p+gQJkI
wbyclO2BVMS+kR+twj340tuAXIc/fhmuk1X6166qqdqyarJb8meq/MzSh5Ug6hBn
7Wdp9Vg6npRWzX7DDcuE2BdaQ6WlpnwQTcB5sZE7oPwHsiPppXhLoNDElX95m03F
bnhN4NxM+tta9KAbLbziV/nihMapdM5j9IyhfpA6wHVn1YLwaN/gd8VQ3ccR6AVU
Cy/vVLuF3gBn4M+m8NJnaHhgb3jS7xC/Yo+VYs4P9/g/RxWCP0iVjob+ef+i2Jd7
Yk8uHcOCiJ3k/SrYJupFyB9M7wp3BYcb074FNfzai8tSSrmdqKzATaKGO1hPNEDF
AhjNupb6GNSahnbA3vO/6RyNqeNy7aA84IPrdmoUGQ4nufgw5kfvn5EQpSjDoEi3
/r6SWpPl5GW8j/k6yZjsx02E7snn4v8wW6380RE7lRn59Ov7wJ9u33+JUjKnFL+/
6Edtp0RvjReR7Y8ErOrh3q3q7hhmlKb5LIOM0g7TuKUMg6eF5ICN8sDPsLa65tkb
y4qkIvB76kVPw5lcKcgBMU2DIG80gQL0GNhUvjGQ4xLVJV4oecgTOFgrS74xc4/E
XY2AtDyXXzghCs9TdwqOcqiaopmw0Yhby4w5MR8a6/rA6t7bX+NEhflJrRkIW+Qk
7c+yHhDkN0xg+lL4ZvoEQjHvC2SZz0Rx3TAG4PpuMBBpozRUWon9ioPv0YBifTiF
N5EdnmmH9NVv7lu5W/09D+t0UJBse0KQdN7rBbU27SmNQzoSBzp4hFUsYvtpU0k3
Zh22iZbLcmwwPeein7hERzcLH17w/Qc7ux9mc/a6DnH67KFU2og6o71759PbBx0A
qermJVhGKYiNUwdOGI3+JppQ0LL3UYvb8qEhUF9i5LEnZ05OA1OfaL71F6zSlyzC
Ju5EUzx6dCHlyZsSqbovLEOOBJWgWCOdEmm6sLd0bLx+ClIasU4t6NWIovbkfnqW
Q3XSTjaj+vi1TsXNulKW/hMkVGPH17WHoqQEfLf5eDTFCdafSlg4NdMsMZM2j26B
dTR8GsW3dA1CtBwLJgwQgvj2HxzrfXItNu+EJgYKdGAuEpSBPHbntXyPjGLuA0sy
2+PfiKsVlHXub0wRkwxTcO2gZGS4zZg8ao+Pi1xNI5g=
`protect END_PROTECTED
