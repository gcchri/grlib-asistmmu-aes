`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNBxLyzSAk2fVKEEtBgZ4DJw81qiuFn5scdwTjFUj4stbqtCyn5ZWEC93zX8yIdB
U0FOq6rDEk7zCLSxR2fxvTgBixYstvsWl5dqBUWwNJJ6es7/R+RSaktW/t89dlQS
IlAs69T8QI50RiNMp5gChu8EOqvBOuvrgtBQ4bT3bDmKtG13+uPVh1oilPcN0ppO
09wZd+DqyvaRU364irUttqA9zIMCNW64rtBeWcqwNqmEaYwEYLRtEJ4+EKkrkwx7
+u1CrkOE0EyprMPXIiO9Icpk0fKIsJLIIYnOo3I6RPgRT+JLzEDzkKYzIYBgCEdG
ob3+Q1zEpnV3Ok05N5xwOhIZJMRe07Xv42oqn8bsVhZMZhOXkBC8+BP44soIFvdr
sagvsbbKX5d9JO9PlwonFXFP9skhTGJXfjgDTRJYSjdCoTpvCiTOsO2eNANeEmPC
KbHiaVyOXsB9R/uVtMAbznuTbWWJknu7a9fY9IVQmilpjoyh3jPyrYNc23l+0dXG
+mz8HZEZl9XoElTHAdMrzFZlrjw+XU2l+2Db1QkmqluJueXYAkTKg1QYJ0dHNxwK
rqFrEYO6I++Uewex5/5j5g1SzdNp3i9HXw3A8djJ/lf9WUHKZfs34lqZKjbKoGbG
fpEAyZq+fUDLepJroC4ioMJakt+aqG7whZcry7x8VRDB/mxUvWGLH/EgJid+MXul
i7J0tfjGTSGvtFFunuvqethYArGtLUQa4/3nU/b6mvitUDeFvi4AOjPDH1NeUZx1
a+7aV9CfsyD0zM1hjPtk315iRVUbcfVUZCRSRJjH8UFvp/6Y/IinE2JGiSQ4HRdl
5HC7lk4dDQKU/R7lr3BsTFG+m7KMoE/fMb8TwX5fFTAdKGtES5O7fDE9VfLl8PKi
V0/bM1CPDJH6aAYyW3ZTtWKhTsXlXJMP+dx4Lk4AAi84ZNqG0XVJEYF0VpNIh84l
COW4D6TFSDEU7ExfFtEsr+mxILXHybhl0b8lpcJTZiEOa8NpMaqHewBd1OgN1+o1
vKxeyLBNUbJSyX8UugZpE3U4TMBh8E3Egt7pjmbJtCucGf/loXaTbbNBMY1VOOEb
/aDlYN+hxQYzJl7Z3yRcjmi09rG0U4DnrcADtKDk+ahdVFqqFzzwPdZvFaNimL4t
oJbiYmaTB2hZKQrmnrSAkjmBZ5OHs+8NaulCk9zm2tTidRXiD/a7+n587JKgO6pq
bTSc228NJXL2iNxfst7Fm9Po3UvZ0MRbNu7m/8MTbxsNVXN3J9IUErfO5nhwA2m0
4L5UEzOqR4ZDoKT7rgSSxw34z6JfhA9ELaf+WF8fk9PTsRMYkRbnVQgrsbLl3l72
kd9cU304dJO8B+G1C4VW+iE1b8P4x5vi4F5hVFt40FlB29DWNvgAJ1zxtVGdju0U
lSZLCwF6lYYk88oiQEy5lc/GbQdvokSDGbH1N+zAd4K11d/AAchbcD8pFfsnIpvL
ofrR5XW3ADWosUFq9oVZk6DVb2DqT5+yZMipA1/tYV6mHiNVssd0gHo/NlxanOro
+c0BhskdmgddKTTIGUAlfoBgELgW0o6IDFVSB7DB54Jr//61cY6T7a8zMl5oSNq7
7fG1PXp1Evjn3eiXJsnI1A0FcnpruajKy3SkfPrDa0Ka80HyEvhMkJq0mDgGtgAJ
+jbt314zL2ug+5IGGiYxIcKkoQ4Eo9y6baqKviG9SazyPfuqrquA3u94ycSg9Svg
mp83k/Fsm0tHBL6nRz1cnYymv9yQ8UiEALiDdQH9bRRY9dtM7yeWh0mLPTdSmcxr
lRAhVMRGqH0lCMsLVzrgr5lXSMVSkrHD35nEAQVBja7iJctByY60sS+ERqXG7Ssq
u5ICG2TWWFzEzb8QmDvP5cn/KWbUMGp5tEIUdfUOWEtDmNqCkCdXbmx5JseRA4yU
Y3LojP4ydWToUnTca1/ksy2kLwus8NmVAZ1+ImGlOuPUL9Ou1H1pdtOeaWzagBP3
GlUpaJBLouhx5Zen+wam55oAQHs6WUyKvhLP5UzhZ1tVopdvIJ5WK0ZKkCPwbguQ
AFl0FIavasnBVof+WPuaLGLlpmqaekq7vE4JheKTciG+gDk0ovDnR/W+a9E2hcNB
Bs0s/h4YmNdMJDwna+Hbxv6gxDGzvxkyFv0WqDFvmNU=
`protect END_PROTECTED
