`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HUK0CGizDbwH6cYY8Q3JG/XpgqelWXiI+vrBUtIuRsWwQiH597xF/YGJnd8RxnO
w+5xrY6x0jYFK9aEa8Ioi4JxaoKbttn+L3Cg63c69otxCjPbEs6CaMIhHVGnT5Ku
Rs4ywD3D3NF2AAm7NDPxrBLC7Gx9rN+4OVouHMl4W9iq4o5G46Gkq03Ew1DgWyKG
8SI08/U77hFHXqfMQq5mW9jT+QfFZE4yshbeXdd8Mpxaoh7KoQXjzVNdBpKRtMBl
bJ2EodZWKymkz7MpmJZ1ESZkKL19pTpX5QwfBqBU9ZiBezA2kceuaRXRqWGYnvDj
XW+2QxSi05neHyZWtPWA7cmuqhhDIlVx1khJHhrVCNDHXA6KzT53nf1xbGwe79xf
4SOXAFAqaqHplpteP39TStoiRVGnFN7s3gk7Ek6HpEaxaZEBMPy4HhG+3NjLGl5F
OErtdFeIF77l8dlGCQ5bJvuJIvVI0rd8BBuVs2L7rfyxMBq175cwQvCmb59H2u18
v/mLqjE8f+TYzOJJFXLJezOsVk0zYSWypO805hKtO4XTc5ZIrjIDXK/K8Qi60Gt5
swdrU7mxL8bNQRqQKM3zXMlEn53upZRUVgoU1SAl+pdoJdaTeKkyYHWUf/K5zRbX
nu2rfjinEB8Io/jfqHzUOmhN1h2aDJdyEo52ga9IXb6ispWdPUI35FN0JMxDbBke
q4JYtOedmIixqxEygoPav/sIFFwm6xMkdkSZHYE/OXkQoKpd0emML4FC3Y/K5Zt1
k55A/L0U/Qtr2rTs3QBUAPFfzgzK0/x/sypiVQSxaMLOv+BOoEaPKoB3sUHQxjNW
QQSCx5t0Jrl4JRrOOvvsB9p2v/p/t8+hD1YpUWw9woBkHRZ6jNxn6SgtsDM7ONLg
8PAXHp2gUDbMwrZoyMwF+5kWt/pc5EtJkQMmkTD6SfCTWoNMN+9GLRAWdp2vW+ft
5A2p+HGhOmiqpQlOJIEPpUUlKMc0QCsiCb+WDIvRPxnBZqp6B4MkHpv/CIOctIAF
PPNb+T8LBlNqcl3DJQ41hI0R6KAyPSdjGk9RzEtyIAR70085dYotP0524RUieNZV
qEMyNmaH4NDV7wbXvFEM0/poYeU6jX5t6xL+ARY3CeA207wS3P6F5y6eB0j6gV22
iN0lz4qafD9v8OFMFTaknt61MNRG4XplqKd1lORV7mCrQdYncy1D0w8+DteCSgkt
kL3jUArjWoMLseGu/zt2bxHD3VZffGyI2F3VOGeacrmLzek5zGAIxejF4aLmTKXE
kc+wkSCBwPRdMyzR/uCrAw7JjY4GCZYw00B++K4iaokEGDMhk0ysFvGgm+0phX56
Nor84xSF2GjaQChN387DNKFE3yQQSBwQGmjbQY0uvv/yqejUkMOiIMRdezjtdcnj
EyISQSk4Y0fdakjentVoeOjj9weyotRbd0CTikv1YWiJ3JCvkGDZwiQIzgyAN2rQ
yLmrGEnKkLVf63Tr8XsYki4VxExjZ+hOYLt8mKCdO1VHw5vPsoCE3yWg/92wulbp
MRyuOEmyPspQ0FtxDShlU3GvnQnA688j+Dgo4N/n9tnK38h2bGgxA6oWVGIgIOVK
Yc+KOYX+QACBYznl8nmRJTWNoMmxrvOQ5t6IqoHBn4518WOuSWcYBRA2nMLAuWfA
dZNKGthzmtOBV5Nqvyf5t3vqvCJyEhJvwZtpmFU3cAR4d/NpoiuIPpWojtkXo4GM
71j7JRY50mGfo58DHoZlZ8FY2hhO/VYpJCndnAhVTCX7pL+5IVbxHceObGNIJZpG
IVE+WXxY+uBv7l26k7QGTZyvZyZG2rot4Cs+dCSMHTG3C/lfYwwNVW5EQdYfvlaZ
FnvroM+hrkW12QDrNAHwSlIBkik7kDYpCtVEsQeE1YT7LliVXJ/mt3aItx/MLvMf
/V/cQfKIoRKhUMebTpaKSY49jdQMnypL1E13nkSFJhWjpVgYLAX5w1JooW8HBH29
oWrKFjgQOQ0iL886U5MOjbv4eCuiv9JNTV81T4PYybBAPg2oX2xJZSQNn2G0pcoU
KLnXZ95CclCj4fIMMsTGogB6jCmDDLgkP4ixV4MrJz/kmUGPamwZoo0zvywi7oJt
bMPrnRIBjK533MIvNOBSoOF12N4i7CwmdFG4T+KraArLzrAkhWqmJ67+31iVvd9+
lMFEo+c545eLYuNddiGKWMUgSeNomcf2Aqqv4+jGjTVvLlHS3M7KmYogXPKXjdTV
XtTcME1QNdrw1eNJbC+CRGuc1o5veQpvcWbzdYXMyWU=
`protect END_PROTECTED
