`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IpecpSeJMy8rVMJLOMbnPT8xJtsOB9f3XFqonCCPR1t0/jqfgB9wTMdfywB64sR5
df3tXpyC3MtiTotj2G56CAnU00rPFh5kILqvl9e8i5yTcPRDV0RRMBHbcIw0IorT
v0INZRxBo87g7loY568U3gAUBFW0fNj4/0dWJXQlBGoS5rIQ82V21+MtGauBqs2B
jOP+jH6uJuxFjWLOCXZapcuFXker/AAx/gkuDaedfLBFze4W21kZTh0TUrH8e6nc
QBic3EKB3s/7icbdddKXGUAHUhIKXqCJoT9UDf78Ga9APMgitx8YD1lvk90DxcPe
MhyNV2amQvQatB4WAcQXKpMyW2hfBPliyV0Lhe4soOcagSjh6zTIDuCJMymE9wLk
Xp/akHVs8Y3duJYVdSFHTgo72pmLNX57IBskO1uLU1VANTDa+lnzE3uShPbfnKZq
Bq6ZCzwHNOAz0U14vmY4ujlJruXLNP7o88eko6ChhBNlK8hoTY5fMphVt61/XH/2
`protect END_PROTECTED
