`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KhsYrO5AGxCuP5/GskezWL+THql8fF9k1kSCIheBLocCJeYr0vf7406WGq7CSB2M
WzB2KHGuKR7jkjNEP0pHcUY6ePZKUMpkdwbUqrtbS0YbDkbP6QEqJ7ZowvRDX/dW
XJjyB7Sb9X4ZXOKIlNNNk0NOLG0AYRY8gfqd9/xoEtQzCFzKdkotgWoNgSejWp7G
WvgHED/t1R+m1F8N08SGag3Es2r3N8+CAvpezu55fqhyUYUlxd0BCWSkdJHCfYKL
PZxXWhgG6WLDNk0GvZNU1Upnvj57mTMvjkQDo8Ydwf3x8eMFD6b9K47XKWXx2yWc
japqr8KMTPmqekPt1n6Pa6MDuWo9dRPRKd9GBrxu/apMysIF72/ZzjXPhWGR9lrg
XusWeX2Vzvmc8cwZU4t1aBb1q9trqROnWeSvVydtLRMG3Wso6PYXU2O2LaXl/SUt
32bWTzPAvrRCEXKtgYeOb6Xy8AK5OCtB+1P+Sz0umPnTTNAzvUP/L9Cgjj07a1cw
ckcGENW9W28yZzbvDb+Wr1D339XkTAdUDyUj1MhcnmbY/eo0Zt7M6j00m65PKw6W
3WAF5NdsEODDHJPuse/O8CyTJohCZ3PTJTc5hU+rx/7PUAsHmN06bv0fqHck8HfC
CYUVutVIoZai8Dc8iJI0xRuvcc88XRqTYBue6JQEBZRF+3vE6MeS34Hf/WQvx96V
a4JgwDKKwC9bXV7sjjU5hRHVF+OuixBpl4QOV1t9KVdAqNecIm/RZy7GJPl2tpBj
h5uk/Sl2XIkATYPxWrJkaclLOR1hOEwL+Jp8JEYWao6ZvHfDYslkhlG0j04ev7Cl
xRIdDXzd69H3A8gzi5/PAkw3flSSDiXZbSSxWu4KnZ7rpCmipAe8oeCndoawYVNb
FXj/q+KixslRnZ6DLCJR1ctAPLMlBFFP8qMsSyqk/F66fWO6e7hhR/BwX9btn7S1
M2qyiyKyBLBj900MgZo371vZbia41H38NUBGUvwN07g9J3Znz0mYTGzMaulUink4
plu25WlRO6D34aEeK7JPbM3AzRSuA0Cq+R5x/viUIcwJkraG9YBFbpq4rR/H77Qw
54Zqnx6GTgnMa9/n7CUQLx92tlhD756fZDGdG6HLbW1Tidcv/q5yXTZY6dTFoy+U
LV95beulg3kwjVvxUq1hebk82kfFavO4wLbnrY5U9bbLrCINO1fGUmJPnDLmkrk0
qQZx0cKO29HpEstFkxaQ0VhX5mto6x/qHieTApE180h7gJtGeBLdYVFgzrX4DbsD
+PJxkMOAqJJc1CQ4Ee/HP3CqEPXV5FRbKKQ6hZvHoeLfL15PqI/YernPzcRQqg9y
dgqvBUVtonSb+BlHbnQ0ku+H3BYQ9Zk3mgjVW7TdqM8vAA2Leo1vznieE5Uc7DDn
DBMmzEDZBhXTUJN1VY8olujeBmGn+6HJLTU8klpoYbz2MLvp2lp6PKHyk5PprqGV
BbaB6qLJuytpG+JIGWwTZFDyAse+pbpyECVTSoBx4nq6K2s1JkrslQWBAF8odjkx
74iiifEnweiV2ZfAoEdZD9mqmFpLy2rfzuOA0qv/b6nhQYjL1ocArVV+zbrU+T8D
m/Pc+W0PG4Dm9/n3ts+YwqbKdz7c2j6NajgrJq58UDBuRJJv6OKHne81tCTVkbia
AA2A60E4dbZrv9LM+gcnZXYYwEwIV04wlYUD7MM+3fh8hA3DqJmAwy2tBNzQvrjy
sV5dghZ5cNgZvf22/23oDLbmolHLpHaOO5iKurqxLC8riZ61PWcGCIf4GInluYLg
/Jfk71uBBJDzfxopwO8MaNUrqPAYAL0K1FAGg2DsBcFN8Fz75xm4cxyX/WjCPfrQ
EtGwghnD+UlLeNFspbR0shTxcqlqysUVZup8ApIUzh0gkz291ZrfhcEpzpTSg2mm
O5uDI7Bsv4EeLc1lJNHk2meg8Q3eUvkJCiy4Krz/e5xSHVdL/dhrcPSAGR/m/38O
yNy0/7pUSkrigdoSCPyAtfDm4vqB2I1VjOVd0ViyJhxGTHcPhB3M/WnDRHG7Ld3Y
1SVu7n2bHeStOPKw/N3iQk66rQVPsquPthcYSrylcZ55vLA7zRwl+JWS2zekNTl9
EfOOxrJKMpRcV4FvT/o6OQvcy29oBw0r4fawla+Gk3OCb7CPFvkmg4e7cuo0F5ix
jYhWUH2/sQwmFNcJnOQAMbS0foKpPB4SyeWXyFzRFSiVX5GjBRCfULR5RKTfxPRO
TXP6bKezi9MN9OTdSn5Q+M3eem7XOfo8Joh9wSQeTiJv5mH7t3pg67jPe0/B4xrd
iqpeuiW7olyItX1RjVWDzxTc7+OC5YAovaC20Kb1MwFgVMhoFjqlzj6fm4Oyg7NJ
86lSZ5ox+ecHypQfQpnQsFgOV5/8p2J6gc0EXN7Qr9RZ1GCDXhZxoNtQRdnDJKZs
UJArjtmppLaJm6eSTonEwHUJmsf12rLktlSHonQdVlSOPetbqVizIqYWMGTkQJVI
swvNBh/97jxq3jGJNGE/NMkDKhGkJzMegSf/qYcslER+VrQOWf1PeJLiNd1Ziw5f
ABPd/i4b4oYd3I5YHt7pdgvQgFX4FjHfBhgtVrXgB8bYvwozcyVWFcKXIpEG3hEP
l4hTxj0d/EcBCc/PyyBEvYfSo2x7CYohvrdm3nfpy4HzXqQzN4pA9S9tZhMlWFAt
mGoRLnWdZilDD6KPd+xDB0n0fKr9bPDTL5bBRPLNasgrbjTE9K+5euI6ZUuY3E0v
6O8vm1ALflN1GifVlwptBaaHYTgCmxt4xQO6UVbefhszyrXgUXz+lph3t1mkY0A8
S7MVvtpFGqGetoW+SNlO+sPCO57sFs6teeky3kT3y/o4pqpL8pSrWTxmmYgF0b8r
xg8kSAY0tZq6QD2ZzLdLnSXro1pqei6ciDcHevoVxy1WauHQ+hOXOhVd9cHDFYcT
Lb6f+VtHfi9Ov1gUCzt0F+1T8Ysd+POS3U7OqHYeKfPcCTuAPpQGCbd6AKfDWDoK
`protect END_PROTECTED
