`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pH7l+w5Dd4KwZmV5EINzZAkpNLcHLDp6JjRQmyoFgP11s0R1HnLKV+QKAAxj/qmk
q+sboLDNyqThCTkCTVnkNyX/v2+BV8sRR/UmtzB0NpZl3dzBOPvcYWV76o196/BT
Z4SDN8y+LjUkMgpUtoKqBP1tSVzXVzf+JElSc2G9Nb9qh/kGxhdGSdWXCfBhdrAN
v+ts87+HZha7lUcunOgAMBOcTWuSU2HOShRxvCJDwC7RGipdYkpprV2fmWvKMZWU
mO+9tbWDw4sgSm1l9lLSYxBEbVXRJYK3gOb5fJQsd+ZG+/rU0GLlTmsYzAXOkvvC
7BJwnVP8mDbLntBk411sQSsll0xa34r1ODgqEc/lh/1qYfzolJcsz+9l5Si189ai
vkBDAB0lG/ALWd2AnmZJdiEtJl0N1graz79BkAxaxOpKgAJgn/D1TJH4JTICcK4a
xn2Ku5dKH0E84iUY8m/lbf2aswRLPKhxZtztAGGml48=
`protect END_PROTECTED
