`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Lv1sU9fLvTl0Aq08mP4QKTQtiAu5NzMzTlLgz+5uGUszxxFu6Nr9sxy9ctrQX3L
94mB+YSrUqicRcKscaV6x4lqe/h9R5KDUUgMilscSwZ+6tCyuxkOgwD/pMczTwHX
9JH7NmUhbftP9KAXYNkfoWbo+QGhPvh4XQsRjvXP0z6lfq3BfzldQbNRZPo2ZxJf
uZ7QGd4wM8p9fMl8OO4yqVzvV+EkbYC4MSELy4DKuwPYqJp3vTYDbDFKaVli+fJ/
cYi+jVo2UTdVnQte46OQhqY8YapJ+tjrvDwnfyeujwaTvJY11qL+kNR14BNzWUKV
LOfPQFF5T0COfvW27IuZa8BezryGc2xJpqRI4VArlQu9IiOi+u/RVsijUmtvliAK
dseJUBNIn44aS7Fy4jNp8mc7rsAcw5EeTCttyIBKe4xP+7bIekSeqASw7YaJoWGT
eOcOPNq/pLfOYwHCuR3KSje3C+xu2a93mqmYkrU5G93uo235eOAwKn6Wh4UW5Z9F
/ZLCX3Oe8V0mMlbDch6Xj+SbTeCxuXPiZ56NxuDFHUvC37gSBE2ADhLk2MeskTZa
uS5m234oJQilpA1QfQ77NGiXhgJt/VtLvJYvAOGUXNEh0Sh84P/Tn0s5PekuUBZ/
HL4j5HacgQcqwpMwGVLSQhGsTaDZ8PUaQpCiEpVVBgn77xJzV6S/GTH9vsm5imKC
61+th6eRVahqWG6hEXEDyA3cwcl+CUF6u3JA8wifWBGrGIVmtp+w4jdDX3wiQmJt
+CIHa+fPy8PjaQ+/8HNUk8c6RXBkbSJKMRt5k7f4zw/SDhTEo8LghLk0v6VoRUJL
z7+dFrHUquPljfs9LamzQ8V1xanYLsm/vsqeOuFCld22Ay53TxiEW5NAZoBT9g5H
KphcghU18lTGAiOk7MbrFTMwPc07B61viOLRjlax+sc=
`protect END_PROTECTED
