`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oKKtgmryPVHNmwdrSQgL6u2SQ33D7nBgpwwpF9ZqtnvJYhbyNNlobu9HAgUcJFJ9
v0KOEo54YKnK8tmHEmmYquZWnOCkYCdKcktFKXeLoAUW9DMgjELcWRlO/yEKqI5R
IpHak1uIsZLYDF+3sDHAgeT9zNKYpgH8g6g6wuyeIIQDM+DGcPCkrpsbVTnV2ELZ
AuUxsxaNRsneOhpAJzX11V6/PVJEkZPTMJO3gUzBzF9snIX0Yt1vhYvheJZU1J4b
Ef1goKBaXxGj7dlkM32aiqheLY4ep+1Gq3USs0Who9F1a6fCZzh6wRYIXgZk3gV4
OydvGeuVy/rLbY0LDk4exRUG+W3nWEjifP8UadLVrteqXl3ubFilA2S3Nh9+IX7+
CU2we53d4w7jjdrElKTcHCA44CNOS4YFkm+tCczifty3HsuR1Vb8oAB+Y08Gywcp
ziGUSqU1A/mEM+skYRmFT9qE800MK3iKiLGTU+mtRFeH/EJGtvHn8yrwKXTJM9M6
Llqq8Ydw9iqyso9dVUk5mT9XnSs7wk9pT2gj3bB6MpAxCTPchD4k9d0v6zuiUSxG
Pty4MwQRhWTAaeXYPpsnKLeeH4L7D7bC4QPAb5IVaEchz4SJ36vKJWN94MdQB/JU
IpJUDsGLcMbX7E8MmL0q49Ri6Uhu+xHg8rJ5iOGguUd4diiQSurj/5NXq8KMJyGW
Bd/T2zbtdt1EQS8hXf+Q8LPUTD62JZCKrmOZ3CmYBykZGyJ/67b7LYmngF6muyRq
mn1pG0fvDj9MufyKh2FwLj0eYaXfSZclLrH1stKFABDc8eYJ5nYRAqA8xRy5QWBX
kDOTXKSZidutpPedMBHb/68k3yqMyA0IkTlCA+tJvNlUFqpvI52gWXwnhA9mFrI4
wJQrdI4FGrTUuwbPMowKRe0PMZzA39fW5S9UVsYaePhl+W1KplwGntf/Hdx12bOK
Cww+2/yablAsHRMbcWWlKeOfY3OlINToIPSnTCooVAo+kkizbQ7wJmH5hBeE1nm0
3jZjnLSVFylJ6219VremGLXgk/ur1Znpkqkcf3OE9Y4jTGRISxCRvLFUPdqVVMe8
g2M7hWFvDLgr075EkY5GNDuEZnFzZnsthub3F5GjyYMnm/fPA15VWO8zkvHDX7/W
6ktFQUm1jEJiMeUWwZLLeApXum/a/d6q07CpRJFHI/X6VOdvDMDcyD4Jd7dC8WDE
SHGMiyZ9DqGouAvI75Lnf0ZDAP0ryxWFkNpGJwaIdHXY6jy7FZnoLXstOo3MvyoX
OzZO4OiBJt+jbDxO66qQuJWwevy3mm9UkCSWKBdpKDCRMP/RJuXXiwnhY2b1IYZE
ciHGEwAWX5snKuuJsafHlD75kL+DblSMRH8CvBqwu2E=
`protect END_PROTECTED
