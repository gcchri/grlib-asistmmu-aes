`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzKKKbia8pBHwpKO+Mx6mXVq54h/DefbFJdY7Tgl9Slz718+rGvrfaDu6J9xoyzi
sWG6AZ+gORlqk93n/yExg57KY7Gmhs8QaK4Da5LoKL2PchxlHfnkDOB4F0/sGSNS
Y6EizVTkLvLm7QdfF94k6wiBhGt2DPXT2FhI9l/2JQyijOFJZcmg8E/r1xMNRDcj
nH1YVMjRrYui1LS173VeGaUWZXG10EG7joTEap4/JLT788cXHujLnj/gcw9FmA7B
xyUYn3xSa+V2eAgVlFYNRk0i7nXwGwgM++HzkdnwJwxWQtHuB+bOFFNL0rdMuXaS
T+bbr9dVsHVFaWyeBnMVo6jVn4T2zVAVO0hE1y6bxEiOvu97iKvGfvYsZprRRmJj
kIY46pJ/8UaoGV+7pMK+a/DsNpB4RBKlltAvQdZUnJx9ZwnN4kD911kTPPPHgMGV
GZd2rSobHa9P/4xXUTI0UMTQhPgg48oDHA05DOGJ5edhhEbnC6eV2x2Ssf1D6J0C
SulyIbruxkS02NoZlY1JxT6F72DvM6lGXnRW5GCj3uB7ZmlDHITWefvDB65Ots+H
Y3mmvSuCa18gnYn820E2t/ux7M0VT6ur7Q9IIS2kM1PwTqzh7ag6l8vTRfa1w8TZ
m9MeaiwGW+Ss/zKjS36zLgAX6TxMGVfRihW20OOtpHhyHoxnaRX5gz7Vi9bgbuJ1
s5P9gLaeU3K8RGLTgIKpfHkkltoCzg0Vn6OLxQBROpHkmxc2md3SUykPrv8Hpjoq
dt3FvtmqQGvzA8V4f1bIiq40eWQfAuj8b6SmnCUgN+29CsJLJ+tUtWysMBDCSEbt
4bx6eNzBtfS223MV3u1h7rhmHtpeL210LwUSD2av5DlByxIUgqTqQQVtZADqstQM
zxKCRLL8UeMD/3R5RELshasdZDLg72L5yipqkkAV/PyNvQWu7maLwvOzSlvsEJvo
Rgba23jh0VlWAPiSlNo1PXtjeDem8Qxa9A6GZTEiplzpLcGlUeZTcxUF6WBtfuWc
SU3CKF0MH+AGh3iwOu+re/lnGLNcCdU0/VpCZxFKrPk8u4nEzEVimjdxxTJoDvdX
M5FYh5ivriLEeDyPu/uzBITwhK3NlafUf5xdkzri1c+elUZD4RyMvbxleCUi6agR
aDcPCKqWhIGVnNrm4bhzrYLp0GBcKGpEqnA0woXaWUbjvZIKJm4M4pq+buLQkrjL
CgjUSasWBuUJOJ27vZzW9YfH+3LBudiSqA+Atagnbtg=
`protect END_PROTECTED
