`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2LcdYsLvXt3YCDIcovZRhhuLg7uECDPfJEWX62QKHrUjLJ6tcFV6wJOqYj4Iy1RW
RmtwPCQviwccbAR94y3ey9CqVp3X6y8TCRDVJa3BPAOubB6jvJTCHHuGosUUCyCE
e2y6CJzEnSBic/ChrlMfES+PlgIa7TRs8c3o854jk6d1VpxpVo0z8BxnGexpoflN
4TfdgEJ0wGbpScWLxalIQF3mlcDPebQBAFBYe/BBTTP1pw1LyV9QWQ7xhMNgOQ1d
CMSBZkRtEW8nKZ+c9Td0kYJrTbsTM/yP4uMewyBrZTRLF2V7DDAQDI2Kl4wyzrSl
HxJjJDYrpoCy5mnd6o1u8ObfBgUAP7X5B3r8sElIvliEJA1Op0NEz30Zwqaf4VZg
PCXwQmjabUP8HMU0vQp5jadxF0IHUGwzvrNLft/3vk4Hk6HnoKr3MpEWuUU9qUKa
91+HuNU0NP86/nx8Ccdr/5j0oLBm/xP/XIelOscZT/J/uVGPinUSHeze421BOxTQ
LGvElYrCYiEnM0Orw6RAfYvc5KY/Kj6qpTn/pQiP6xOS0q6np+q5uyuCbntF4uX8
ksu/bWAlf1Pd4x1lTkkPjGqb6Aq9m+Uc3TSkKbCwYte0X6WwPneDV9GI2zK9B8Na
B8zxGydR2ytQuTBXC+vacPDlXZlCkU3rlPZJpt3mkTESjULmY7rKGTNe4DufbScp
WqinDm6BD4iSOQ46vaT3zsSh7TjwU1pwMK2PPwCA2tGDo9kO38VNqmA54PY2lcYB
+PNtEZrtMF+W8i55GC5tLq+IJQBJTc3/ar4exfGkBnh6RCBLEdjcO9KDtmdnzmFH
5NAmkTLVUnqLqgTS293ag3R/SlCMUmnwuP8muDh49I1/fhC6Xc/gzviuXCuNu6eU
MELUQ4WDsju9Not805BLn7ncZwAncTnN3SdIUpC8ADDtmsD7gpKAW+A+crShu+dt
FgYg9pPqtSZs40vx0Y7lMpH5blg2LNvvLhCe2mwf9N4wPY49SOgplbZ6E5jRhKtp
giONK7GQyqvuKVNdxbfRq0Yg00w7RbOp3TnbwUqkg6XV+XMDKlE8k8ODn0qeQjEB
ZxnCT97rgmn352pYb/x8dQ1HOIzVi5mhV7VNOKk80lnNfQBIYQvQHXDrWCdVfTSa
lOSzUSznmWZnWDIsa/9809gGRm0UKQMKJQYg1kdGOFuCYzzHvlSZ2bmC4L68fxfv
PXy+Hgw2hOysXSPsaBVJW3uz5Tb9gNCm2K1ir3CffEyVUU+8pBVj2mbmY9+b4eId
KBsVIGoJkjJwiFhrMGB6nQKlsupcBxspJk1sBxHIzXjPZMGY/kbxkuNYH30Q12py
1beR7CW++mrQlPP6FcPmtUbFXOsq9Ca6RPXsYV711kNhQOvz6wXkyU+1+ZBeHwuY
s8YtCB5Zc2MHKSQITBoW0jHU6tQ0cbp8zNBzicm8SMtbeUABCrgt9EV60ncNO5u/
aLP1cYDa947KUEL7jiSysorRxTGTVAVHRlJqwdKn14XvutwZAi4fJFyoKlmbTv/k
oCD5fb7o7YUC9w4JjdAu+187Jc0wRvHlV4oLfQZqR/JwkzztEM40eGQBvVVJLxwE
7dzaO6U0m921ani+d5DE3VnQLmmPB0VHTK/ZqczzDDIHe2BcQEhnzwFRR18P7fdy
HX7hDnTfWulaJYNeeT8tQ2rTL1nUkwvSTicS6ZwAjmZbhTsybOqHItWx3LLPZPkq
5HHnUzftD9ewPnzH6O4BEhWHME/EqHONL0SexdgSCY0XYMIbUBTUq5mZLiYqHTyA
Px9V66ywwFEB5G3je4+NqHyTiARaka6v4/RVz2QraWgSC/9G6Vc1plpfOsMBMKPG
GRZJFEHH7iLCSZPQQqK003uu31yKhGz10MsARp29/zgxK++9qAra5D6OKb+Qzyxz
IGR7hQTEpd9mgmYZ/ywhORSrlcjGXzvJ2Xnr7/4FjhmNS/M0hFr5bgJB3xTh5fhT
gX9RvPBTYSu4VQO02jpcZ0oHLYkO41Hbry9oIdRp+PoJoJLsShlxSx4ta+MHAtz5
00GzbCtmmFKo0cxIQmODEnLZSMZycq3hbR2xNRVoV7PfhukcxINH1WO2YKwX5tHR
q7XetqBdfWiMVHYyoxlsMCuG+/Bko9dg+eBRqRYYJ3alGdCo/najdreGYOBW5PEd
8Z0i++d9FmSLCXpDzQsszgjZG8CrxrVTKUy+vN4w9S+om/Snt3ufPURBYmi7Y851
ijsud1WvWx+tjb/EtYtFynJkeh6H3fq2nEms60/UCG6slBIZ8YaFh36ssi9fr6Qz
8kgJS9wetF0CdNsvPboMDD8VZmM9MF0reprzqKTvcY7UbqP91yr4HzTMf8HAAdrj
eMKKutNhXiZwUZjK6iG3m0IbPiQtxsG/nFuQ5RRjaM1GY49o15EvEXDPsbBakBJZ
OszW4Uq6bwbIZolDZN6Ro9I2Y1mDtUrPEWsSe0P0C4Fn+61S//1y32fwgf01ZYRG
Vocgl0hJC4Xj3uj6jFLdriN333tKsRbLDb9bpkOSGEij5SX6y0u5iQ3JRQgOP7Cj
rOFqQ383HYxLSt79NICvjucWw4EEocG6YJDpKt/xcu9yLJ2niFSQ8TjTopJsJUJn
oRusURzMgmquo13y67v8jaojiofJQJINhmv7pKNSPWa5REoegkC6fXnAwUQ4RciZ
iAap0FYZSCbU4aguxEPmM0z4RRaijGhvI60R3kct9cFmdw+sdCiIgf2UAsGgvVJl
ZVKcnZ8YQmprIjFfA37liCRtpGwXu5NSTjo1MRGOlYGtJJkzSuTmAL7wsrJaUI6G
3KDcx+r+pBFnn03csiGgWIgbZTWJcHdrQF1C9yWqD7u7tELWwzoZncwDW0bUWCw8
lZnFacinlmRJQbgJSXfkZB8k8MHdkTfpDscLXPwavq3VpmR76wW2+8p34i46ME8b
mVbZfmcvKG+v61Crsb/BdiVBMyGDhpXHGSfkKarDbn7aB/gMbyaogOGne1J8VI2V
HIXrJ3A74pN5RVTcat9MV1Hp/nmnWki0j6FNrZZtIaM23y5RIJLFtR7Xfqci0swE
RwxBhAuEfaLpt9rhAC8vYdeI/3uhJ0thsw73ggFg1InwUQ1LQm4K7ch4/uDTSX5f
6tuTdW2dwkmPTfohfeEArqCD/Slw8qWLF+V61X7kwZoTiRbnLgryehLu+pbC/2ib
Q3l2/AHpRdRjtildYOZoHHFdXVEisH8bp0cE9hX/eVIaH3elDMBNYLHIutSdCBF4
7zPMRTbtZ0ZBaEqHu4SfT5YLq4LQT8bsg4f3O2bDjhitEuxUL6OndeLNSWkbnZxn
hTMJXTHwRujwZN+0ToqjzPIGaVP9GtZ/BefwQ6suVLXGbudlce01ToX5TH9x8Tq8
iIxMikE3dU73bioq8ca4VFBBQs3YZeimjBqXJzeLboZJFKwbGGqfGz0wQzKWeacE
uyNbpTx6CBJuk2ZcLIEUFeAEMB1UwA065v7Rx1dzhHXcbE5hzfmtvGaGy0Ss5DCt
Y8vtwB8/7LBaY1RmaTBndqq3UAjUvwwOqdO/Co9ShPqbF68Cf4FzFzfUTsjBvFha
DV+3JQvREF2vuf8gMc/ifOPXctV14xGR7AbadAXumMKSYR0/AuEW/YwhuqqTeA87
6NrMTKLgUQtRFUITCy0u+lXA/lbRmVzNAFoc+jykoIvJB+BUnmN5x97FwkQw+TAW
a720lEf4t7DcQmrTZMcerDmOWeKGA2EoR69UZZrW/6nQp6JSDMdFDG8cXL0UqDn3
8l2RGLrfThRbzxrs0504K8GuEtjMv6PKqoWhfU+Gzy8gM2vA3804T+cjQ6de/hLU
DCR+rmFkF22ueo66K21qJwYbpquAUXcs1Ulu+Ea1kEFNMxFOaX8Nb0yw1gusqt4+
GSbFCll/2F59O9Q6oBjCscFCrOyclQ7fpt/f2Pszm59xJjFn5OJyPKphVj5+XNzi
/3azhv5ERrcmp08lMdu000eadu8iE9cq/Ct6WSL+MCxAFK8nnFxRZQ7AYdOJfDn7
u+H0sCITcalBHWTpUeloCr4XPyKIB13KJ5jc3vk2cfGJc/PJEmwWtnh8NZS1SdCq
f2sVRhw5JPJyVRog7s/7dkDDvUBLx/GVGQYpM1m/KuPxNqaE+E9mqkAoiv01eJ+/
VQV2hGa+osI71rux4S/mXtfxmTl6d2qq6Ou3JHaYQAtog3WzdAUpB4Wjo26KtAl8
JDFYageJLSny/bXp+7tf2vGW78CUZCccDX9QFEwK3t/1jh3RlWeDkjbkJqvmMWxm
9w7bDaWi2oZKJiKlPK7vEGT53OOck7NVJSQo/5BMblm1nbkMrLGr3DPbCHeCRbPW
8dCHpEMxF9cdWGW7eu+LHvMrqUNn2aScmXC5PcTCAwgEQlPJmymEfRSJMGxQ/n9G
47AguoJZAxojd+piI63lZnzeWY6fxAD0TtXUlP5R57tqfDnD293+6J6rZ0+8FedS
AC6eK/Y+Etzk+knT/2Fgf4rvTDZhbxEvYoTttBVTEisRl+vcG83gLuMIEbCITGNN
h8MZ4uTSDLfNtR/ciFABzg==
`protect END_PROTECTED
