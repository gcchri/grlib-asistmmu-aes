`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5JhP9KQrCHGIHcJSU0AUlGGyUF6MloVlM2xDc62qTE9DE5szvTNY/d0nxxpZ+l3
DLQG3+U6z9mu987x/UHzzvwKmAY832ouNa10Ebo3sduY7CKMP+LCHoKJVGQm0Eez
MhVwT4gStyt5+SlDeW8RdWsfDHHf9ImZ8/wgeeDKLWdNMJM5XFi59nuwq1myapcC
cKSR3NuqlJBJsdRUBHhE8TsCWCiY1TwpHMHdexpN7hYS8SSBBZtPRrSima7hwbwo
yncHG1DHJTcLiBxU//v+OPdlbA5ci8miE4FcpeS2g0sGsIECpB+FCw7wY1FoHksp
Ix8eB+K1dJLPd27ToPvZBe9uwVOoA5nvs2VwXKHhqoAz1P5yuolc2vtZd+DolzTr
VsuSYzbJ6/4ElVuO+f4BUlsvBCZ39bqScOPmq/yOwYJ8gsbSHVRKluROJcdXLUpA
0ztNxRo1jFpM1dcCzugS0n4sku/yXz+Rwk85BMygxvOrSHe0GPAvyBHzSV1KLg9e
YxsUvy55GsQM0t100JR+C777tqm63o8EcU8P6LaHa0TcU5OqOBacGxSvUyL+O88p
AE1vBLmVq4WzvEAyYiIVByKZkLC5uLalfA6oBrZWmascgBRC6AOm2JiBXzlrlWgz
sLtxZqJ/El/o6TdK1Sccvw==
`protect END_PROTECTED
