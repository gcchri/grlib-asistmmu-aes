`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MgKpW4Oi6isIRY47SHqPMji1TTV2K2opTzS1O7nzoNTUl4gm+kdXWhNT7JpANjdn
51tS5lJR7a5ixxIpmn3MXUiSxSyUtOFft3zzvZ2/SCNcAEscnYveoZvYybJAoXYp
89qHuf06VRat00gKcae/Sm9oMGgE3GI86k5y7+OuwNhsucMRwmR3tjYIArNNeXAd
RnXN3LKXEe2SRVnU/zhj+xC44JPfgpihcOYbBrJ1Dcvd8GpU1ejGynUxkBvnoId/
kQlZUmdtGaEyFCs8JgCLoFP28uxef9ky+nsgsxscr04LcBNxbbB8nxnTG5nDgW0x
Ru1iQncokSzATJ11yIejo0syLaYQ96LoYtreFBWBhsKctO80l1pMCpAHWVB14G7h
JL6Jv8LSb4SOgyZcymONiA==
`protect END_PROTECTED
