`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6iiAOtiuyjFis0OyFCbrQ+Bv3QZhYKxFi8Iasl/v/ex1l9h7EOgRtljEqHNiiFP
t1y76UpAejWjxlnaDUyE7dyzqn/9hywk0myhYLAYF7vpAcXtvAsgmwfVpdClRHVw
CdMM0yZFkhSDKFP8CbN2m+dE9zPLhh6VoDt0t0oARpV+IZQ5UecfJXMmTnZ4F+mA
Eg5Hctc+fKcY+I9VQSiNd6cQLW0wxfxZJd6m05leH+0fWHXvIroZNTUl3LuhYwfD
YsgPf6medMOJtc03RGKgUkQVPRUGcIRVnoLVo7E3X4Ir/0hN47fdBL9pCdwgG0tV
PwngmG6EcPHbtdpJSojGy7XK9SO7Hv8lfUar4BR3pgQaIvKThJazBN3+um8e0ZWb
KQilzJC9t5PdA5/33kgtEoMtmAmzlYgDQ2H3eQJFKaI=
`protect END_PROTECTED
