`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IoceUTkO2WlezdGyoCsQenKdy21jKIlDW2yYXGLCJDK8aAHz78oIL7oINNliTaEw
dSsY+h4RUrfPJ1hM/7J2DQ4DMp5vtQa3TlXf71SP4gz50UEOxBt4tmbnGKWym+ha
kBeC/aYF9yXYaiQAu+zwj95pTLZjyuaTf4iHKg3xD27wZHZAX2Y7OUnl4UDS67G2
2nlQWGFRPZRIkJF14NLbUKG1nn4JgMqQ7AIzVnP4AM82mCQWZxdy1QXcOPpx9Cl5
QkBL2huhXZCAvB6v+b3tAD2dE7/DWtAsoAZWcv14vzDHEPIHtUXCvt+TALur3mFZ
N34JRk7X195TfJD6vhMkQB3hdZPB3OqDPBYWEhfSIjPR/oIBdd9sZUxf2gQTa+mB
a3zFqU+2GlR7fTUUAtDahuLFKtn5S5OErGEIckMuXhcZ3gddUWljeAy7HjSrtVK3
t6YzFE4wUaOZH+rg7EA1TcNT7SgYH68uA60+YS/KAa83PiuWC7tkG/3J2PvReMSk
dGFQlSkNO9x7OweUqeRbhlMJgE/7iycNKe18+h+OZs/Q8b+8wfVzwV4i/tpNkCl5
j4QhWC36l4GV5zY0BSUsy9b5uqE+rhRUkkaCLlm1xcH+LTlq6oQ4cmvnp6BiGVeQ
/eyAu7zfPGcL0owWpy0osNdc53A+fKBuG2X4A9vZJI9/2Bi7dTRGya2RhFVyrzpv
4//n9jL5Vv0A9jAXrfv1bY1BPt5HMZQzQFsjmtFfWpeNhwSQVebEwooveQRwOT9u
igBbI9Zy9N3loS9U2AgU3+RWcXkliYRMDf1PSm8PCCcF3sBKdUkSxVMXDL4jhHwK
fXjxL16cruBWGGj7Sch/Fiq5ao8nufQa7IaLOBGSnWBq8oZlSrtEwT9MdoJOIHrV
C7J980B2sxBwxPzQ3Gn7F6GOsf6IiAHp2O0w903qIUgOREEViXl82iZWTGHUQAhU
4PawX+Vx2RG+aRd0Hun+VwlR8q6TvRycWaiphPiAhrvmNAq4O+B4yt9o7cBG8esF
4tGe5oMgl6lFihyji4ydLq4h6Nt8CMmAczE/n9eBpiKGRS1tWkpCakdcXI4nwYNg
Zkqnye0t+ZxDvBBnedDVkBRvPr3uH7OqHsfGTRmcDEMLZeNsSlRu2TPx51EF9ewD
c6okFjUyvEKgkyt08KxLus9baftuD+ImDz5YPrZNfvc4RwQ23IPpA9AfevOfkGA6
sLmu4fAov8AgzjwjkU8X+za7esu+BxGZ2dOUWbdoQ4NvMHARXr0AQBJX4ciXV2mx
WQr4nefgPFioLtB0KnoS8WYP4sgzyc+lUWJlMeZVa4VL5TL++rmTojjIadJlvXYP
BCuDMae2EPUdln/Oct+QszLzbEeXXtLSRJePg0jYacIf4Fy8sS4FQXknGLE7XDG3
BfgdoTxgS1bk6f7YCLvf7xn6iSCK8ULivlgruXJ8sZ0V4qg9HZz3N33OsZbfdq9u
gz0v/k91kkScXif2q8Bt2/MGkrw09vnehJ8V88Kofk2MR0mlmxbCyea+vWd1tvSx
fQfQdJWIi8UeugUHncz2UIN3emTTQNI7P449eOho6YpLgkrIfssGDaCIN5K4TSw2
7uPEG01ZjcexljyY4QIBJUflj8HBEHUehLjHYdIbGHSLVgn7jLSYjglnE6YHJRgH
fDNG1dASO2IEYyaKUK2G1pS+8Cr+H0mSX+ZiyMNf1VCLYLdiT9o65palAUpqDNzh
RIZFhMBtQAgwm2m8nF8iF4grjIcdNe7VzWHcVRI63erqLvrJQQPG5sFFDs+tCWGo
J2fTyRGSdg1mzKJFFP4l/9HtrKPXgL1Hua3jjzSb+V01L6gyX2EwU+XhffKrCG0m
Jeuvndi6kO45iiVFktOQh8hbnaNX8b1W87JaoKq+BIoUzPuA97ztwO7u+KNvjMbq
ov+Wdf54zNf4CVtO95Rhow==
`protect END_PROTECTED
