`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kDsp6cc/J60xbOAsHoJu9mduTj8BzM+hea1jEB3ij9ugzgeKftTNPVt74BT43l6E
ghfcXtTMaJYM5GWoemgg3bYlmzzhHCmDzKQXVYVp71pIHQUaY4qz+TQoJLWdSh/G
M4ENC3Tefg+mbC/2MRS6QxdyCm2/x16frbv9bM6hGW5h9FmCrlYbywaAyUM0u4L6
9NikOxJHZqmQgSpdk2CDC2JXFl/BFIqba3BY22ptfrA+P1bAWyllhZvs+VdIq5JC
MiG8CMgzNu/4TMRN49gwUkmNs0/4+jKOE9nv7fEq1dKUKGoI3PLrPwusS1pZpR8U
fQB6sd8Un9TnEgA2kQHSGz5viq0gMm2aZ71n3R/J2VZygKuLWXfekHjptX94qUGV
FINGKqCM/kEOROcfSufMFsR6TrS1ycAZXdyF1+qKxWLVZe0BAcc7jjvB6EV/vU5A
TewHdmOq9+9lzT/srqLVwTM0IK0plkgJnXNK4YmQShIDdExcFiUy94MtCDwE8yw7
Dd57Xzx5xL1x7NCXIT/CGgD8AWe7y6LoRaDN3YW3w9Tp+VY4VLHB7tnK13/+jFzT
gMJdBcy8ufK4vffxfyCwXfOsCA4Pz9tXoIdmK3VqDxVwUxwx63VVY4xsyF1lO55N
RxYwJyygAoBL1rqlDeFvSXrCoOgkvJVddJNxq4XX35c9knE+D1y1zzOHpMkd7kYI
LZ/O/9JTkpJvxCh5L2q9C1B249PwN0qD2pu4G+0yn5kz2gWTyPVwZI9DqmKQAenL
eXCLcQKDvCasfjh1QegG+afv8I+bmjDr2NzE3Xib3WL5k4IzARBtgCJALpTR7cqi
xugVIDzZ4CgDslR914LIAomtKRKv89QGlMY3l46Quo7099OKiNs5/2vh9QrebacZ
rZaXz4QBg1QAGfAgy8wRJdORCgLz8v3FszzPl0eCPdAYCHDV2n8yTz13FOrU1Tgv
+hhVl9M2zJ/xK8B7Hl0RhAxl3L9Th7WrdMW6P+gQEi3wHn+3ytoSKXmh/726j7d1
xfF94jqsj/jDqb/vQ+DjyxamiKROhkDQ5X/Hwc6uCuCLlkAxy9eN/WAP65E0+IHj
TKWXl6ibgI1lqyHPP2E6aCyS7Q/LkiTxIc2I4y8M9X+SFsWiy1FrTyYBv/N1WnRE
7NMydCY4kSmlkfZ6pon3g5OtWOotVc9IdqkC2zrj+6ARdrnqIApXQPCjocQVUPAh
5Xdj/Y6PbSO2/eBtiZVn2OsrEC4ch5aKNcOcT466d02Tc/xahmm8I1Gj11Zropsn
ZQVf1U8UBtjvGKAMyjFDgAqrYLLhvu0BZwDmwclXBib4n+/mAIU4D7+RWzEThzQd
2meAFX4KEh+SL+wD2xzPVItZ2D8xWmHII40VxX8ZEJbj7BlpSp+DCSUqTgzZw5vy
arGfmW528K7eB4A/eekR4Ry2q0SC+q2uly6xUb5PF5gQkyBTA9GNBYMWkjBEGuXH
FDw+jotnHLB6WC3Z3aGvtXZpdET/r2dcQs6ZQfRHkC0m3J0pPB1h76diK5Pxki0D
UbopBXYC0iwZqDWWHbj6Fpu35dU8solnxnNALSn/IQV11b36xFK/huC1Hlsynko4
82F8isiNaxwCCzSckXOl2JjOLUBC60MfRWRO4CL6lcm4wW+zLh4iXY/fHBf0bOT/
AHgddXZyTzY1leNuKLSZlfINAnNuAX73F5B297qvQ0WD4tDmG1sb4o4CB468xEas
ERTDJB19Qxwn+dHSwn/mi8XfH7cS3q9GSnKx1+2SGp3H93+OL82feHM82iATCnwe
UYFLkNbFboz/9gu8ZIxnnqLfNva7rgCnsrn4mzN22TqAcR9UqxHas5SAwLnoN15Y
Kk8pqTNZb5xBK1w2vwtUeuEYjX5mPhTyWbkEBAaDi3PlpSPujT3/FRs9wVOFLpE2
glsLG/VEfR0m5odxTAdfZ4Y7Q2g87Mn8wm1GQg8jKWXp8ZctUw4UykW7D7O5bgWj
ukW7Z3jf/hS8IXN/1KatLTD9JOUCUE5IeXWiTLbL4u2kCaNP1GD4n6a459o6w2Zo
r7wALO/XU8ORnDGY3XtZNvUduMGtu1K978Ufy2mo0xYn3KRc15yIRMyhnU9aBmuW
FwVOOFX56bXR8qZ4rguldG6pZYt95OiCVbhUfjPDit2OUTOlMfE4j2fq41yHg9CH
Z4NtezXDfNn7+AkAVgC9vki52AYKeNHUGDqr1/zMybrPiqWA3g93iJxK8YRPGLQz
Ztv8kb8NJThvaEh9BBOptxPfaqELPTFxRyrV/rI4J1c7XySHwFd1FGTWC1WWR3UU
QELKaZ1Jt0jheoH2E1jwIXmuOAmmHly66B1T/9N1wz7/inLoPPC/aBI3MC4CZ+rp
XPv6y3Wwujq1kgLRQGjonrwk8E7qSpZ4fLLJMieJDnWVl2nL5pbDWGBbkY9F/2+h
/V2Lfsb/9aBgnTrWUqGoF3GR0or6u6fguXMlvbf5V3Fo7cgRIeaIIe/ilbihi5OS
eNGg7o8tQp/Tli6WOzPgwJeREn7MvuJ2C6WYqCo3P+LNPF1WzGycNhjaf7Tf93rt
f/biuNMl3FsMeRBwmXMrYsbCBbyiqxC6YLQdJGc7e6Rw9BIJTQJ6kTEuxR1BP7sJ
Zl0b5nJnIo2Q5obRfC4z04QIu2Jnf89+1FF5knpjw0dFKfO2rU+/r3BGLhtOynw2
Z1oKZEeXSo9A8p2PFNhmv7HTEoJoQe8hNBRdIIYq26pc6/h15eS6Imz+FI1BRJDf
vO+aIYrDyQABrhcVTuUIMwJ2fJXn2H9qklZbU3bLa6p3+TYhe17I1M4BVIEA3MMd
z0+sjzEOKVbgUcCi0LXP6vj6ZtHbIlKB461j2MwyZ4wDaBfs4lpzYfjCFR9AQ43A
tCzmUDw3imF4lQbEzYN2+VcUICy6XjC9yiOD21hdj/Zu1KjWZmz9Y286pouNcY/l
T8v3BD+s/xMDiqyaGFT/cj32c5KKQfYqT5rJz7+Syi3nfV2Mzi2olM83i7JndXpv
oiz6cxdNq681AhlXfKv8bz2aBIut3nal/JZ1nKb4MPqGxTZH3kAfZpQPeV70dqzI
zXjqlbmegC8AQeASt9OwaU6r0lMGHPQkXrfEcr9V9GPW4+yI2rS09HkZsIGX97ak
qbxUsWUG0Zfeg5ZtQi/WvnWA1J+f2Iab4a6h3zy2W7Y1I45tTfx59V1CaV3d3iml
c+2gsvhqFJ4iPMzrKj7aY463CC40WTBFC3G4zl1P1IT+1pzRsp+aeqKYWIDemtKe
9bLVEX+G5kRU1wSATj1I6l13lkwADMd8WGSTUaVTgC34qm9sGuIQlFGy2zUI3KgK
iZFGOBssdd8mACxMGoJCRLEw9OD1pJ8YB2glk2e5ojlxnIui+mbXc+jpPHeOE+nc
HHnM2ycMcnGJoBqEiNzDFyJgHq338Lz02K5LhrHoSbiUpbak2etvE09aZqFOJuUr
W5oFrduLm2MhEI2mCYCMM/JhjOb/Xp5UdSD7jduujAkgwwdJuk3BdpwRSniWfVbs
gCOq0Zt66ASRrh2zPh63C7fCgM07LEcXnCdVznQXVslPIuLNBFeftExeVJLPTcKW
0zKOeM9TNVnUsZA+YtByjWrO5NCDg95J2V1NwYy5o74BFXC7/6S5KXBqxkz6LrBr
A4nsEDsh/LmuyHpHX3OtIrB2Psf3CmBWPi/YTUnPL0SutO9gkIp3iD40e0Tl2p0P
qc11lzPq/kRjWFd83MWWZI/l3sZBO3BpZOUnBuNwOPUJeBBmsT4Pa+FI5YQXL+dQ
emg/rtPZqLdC/5YtAiReb3hxVeEVMP4M7unW7v2LFPKlWUIYN8MUiaazTvxiyqUT
muD0QFypbIRwdKAFCR84t5a2mV5HMsCekkr83zyB5TLCYyIlDfIrcNXTPkyxebrN
fkA8GEl/rL+RgWNUv2pOeiVMApr6POMO/AWUi8SbDElJYDPr/5PXM3FAAEfL9Xxi
vHrxcomkt2JkhMzEPurTiTmBIP6N4m/pvuVD79KLxVLbWC5mhx8tx6iJZHQ/HaA9
ol5nyixUpPFLRHeXQeXn3HAxt7Q4qK12sWjZuWN/inAmkpbwmtn+slAa3ID9Adqw
KR2VL2Yb9KSJrvG+BuaU0AF71mQ8mWT4v9cQ+DB9gytQqKbDcwpZVMdxFL4GMdDZ
EEx96hd6PdS1150IDZC+2KQplY9+ZdRTqng/46VtcPfI8LRmAjQfl/8MF4ukLT9y
ZxLeBbsD6P7S1FYMNz4+9DrKJSLNAOufFz8hDtPmOi0Vs203zXxaCXFIZtWGglBG
z2OM7KGTeErMGertobMbDFh18D/P8oER5lG8RLl0JkFdNTs5eIh10cpyMwqFPlvr
1nCQmzVu/PkxBiSmKySfebN9/Vo/On3erCvGXxyIirHUdC8iHo3zMNkNBNqOXss2
WZYjhM3G7gou2X5yA7zqJaEmUsZhLAQNKH9qFrn64oAlhWOktKmXZ99eQSNX19cu
oti06U/HwScgVc0hwn9FR6eSTogRV3p+CbgDbRSQ4kM9H0DUrnQ8pjmwc0O/75++
fHDcqAQ9JMwHrvL5/8EmJJEmeFejX7TLi0+MdscL789jiPTE4CrNwG8OYSkCcyA3
4Nf0qsqytGhZyWwpi0//CvrGYoztrc5FQltqtQpz8mzbHj9IIkI7IOnpdPZpERRe
IGrvevxIKhOYvNIcBqpXVODf2NyhkhZBO9/scXmW4UVxXez8nk/wW7EhUldCbg8n
ma9estjH4QxJmRIQuP1cN0cQbg8IQHSwUWI3JHF9QqjwjoZtpVA4srMm/K/ozBVl
B28KxOGEMK1aP0Fbfy2aA/cqkqWFuaIWS1It0MssMAnFMtGfkfPVqLv1qyHNV+kI
VlnlY50YwvTTTCve55QobYDkh65MnUz7Gvwi+zBVTZw=
`protect END_PROTECTED
