`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sz14cfrjOfngkQpMG1Av9AcRZDHNOnvCg7ANstHT1rRIQ9XLmG2zpiCASbcm3B+X
iY+M/uXJWaxFhSUudyHl74zrYWN8ZR2Ct/WFETvv9tUCTkezOSkQQ6AgpJGHgek6
k0DHSOOXP/qsTXMiskFk1C5wGKRN7c0eAy+2bTrASOlBpmqa8v1BOg1ypmDse52r
g7lSbReKTTmgJ1V6nEKtzodDsC6YhmDfEjtWCEcsUniEsHDgYxzzpdeOqL6wR/mX
lSMD8oDQ4hYfA2jXzst7gSBb7EkyOtIS5wkm1loyGo9HqQzrTXvxk1iVkQaeEad0
1TZ0tYQoGPbebghT5JWlpreStB4aahn9IbpDCkpXGdbzfkdasI85vPB2iZobDGcx
kWvY/9pWoXIqCLyxzLXV8jYuDgR/RzSkUuSsafyTQLkr4i3G1rdn/O2fVFVqxth1
rPpU0HhYgI4NvxXGFQf91r92YHpeEPN6ntUwUQMnjU17jKuGKojnF2A2dQ+NsTQH
5jFwBK9fBMmTJiE8rK/WtQseyB9jSf3sGAm9TlNQCvcDP8GgOQmdLnXleHDr9ZQ8
vs+pUk4JuzftOi1AV33Sz5TuMMpd+QSAelhCBJVNrrA4DIZFK94Dwq3Z4aRM5Xrb
ATArvZTY92cMtMQk+5/j6WpuumWv/YswiUtrhp1ol40IQg0mBqkaiV6qXB7+CveH
n0A/rZr+YRwybT7KOjSldb5hEMEVtchqN6Z0MPoPsPoXyozBK1OnZCwXVyIAvP/A
kYumA7oY9IE9N9e9U2aK9ZaOBpYdgnNrC0o1FiM64/RpQDNxlpV6L/7pnE2ZylsM
58Po9SC6po37jd84RUCz8asB3SbXwM1O7a9xeJIdMydxMCHxkwmCNmBqo/+tLd8u
6XkpGyeCgeslriM8H9IQFSbx1BtEmXA1LgbxLPATl0QJLSbEiI2MUBxujjAx9O2O
EKWk2NDB66SUm7NrNhDUZBzCfFY/ANXd/wd7T8/QGJJNRLdrvwXrrC6nb7p4lDR4
C65lDkdHpatW0nLS9Jm8hOjxtcr7fI91eA7ISSwZ9WU3DmWHkMzQHh/HbPJ0PRCU
N7krVEPMVyXgSU9YXLGculWMpjcRb/0PiNQ3b/6tnwsN/NarElFemKngN8zF+CQh
Dx2ZAKo5IFFtZI5eMHhkR0U90sDTWckyLlA/509YL2StlDnOuRdR9yRA4eEEhljb
CQr06qdcI7QOTICrmJbDqfrsLYXvQkMGsqsJwtlhMNJsG2lyPfq8x8rBB1LZiucy
ApVIFwz/fhCGDdYuSyLH2PCnxa66NreomH0pPRVg8pBQYhskOhzLr+b8MqZ7JZoQ
AqLGVysnTxmJF4RXFgTQFoVVs/OyhJc6nt5IBhwAsRBZkpCQEA+/697UUc6TVe06
dsT770SoseCj/RQxC/ryD33mEY4tyC+IONkoZrAc66fjaHqdLzOhkfJEIqocSQNk
rIUJ6S6D6jhoRnXUE9AZVpRbIMfIzDPl5M2OfW6Yl3aOpLFeFbsXPV6NwQgzrl7N
WlnVa7RSzq9kzKLff2M85wmapnC1/UueO+tDirjAnhKgkDeA4lcvhfN1CVG/VMi9
UO+KvveJ+0U6bo+1hcyzRgjQoJegciI8PuOcx7n3Z4Nk5PKnRm51FlJ5K8nBk2g1
LyCmgtg9adOCGOxSHUpCFQtVU5eXb60YOKP3608n3ylL5/yNTSZfY6Q44YD3lgex
CJ3A4KP1kroOey5tGMgeKHGUQHhP9gFgsuS29JyBednp7+0S4ejOullb186Nfntf
cDpqpX5+UsQQPVtqv20r04o7wdKYnJcVFZLV5tGeDXQXRDW+NH/lXfR8jnL7VXJ8
AlP4Jkw4GxAY5ZKPVMkZExzeOHxt+imbipbrts5XydEGZqfRXgq1528fO050Lj+/
/UterdD0Iz85nbeO3F3+PtZHebHlZL8ConzvPQn+MqeTCLj2iPAOgKwYUT+dOJuE
BVHHSKrxSoujJUIU0l0pomj/WMcXBrmEuVZdEMqvSb5rquksiuM8XcAvZdEjPDly
OPWCAjU5kYaihk0SE2jIqyXtWtT5UOj1SgEbVuJGndTZxz9pUDccmGls4ZVCQRuV
U8U0TUCv9Wwz0ibd8mHIv2ohTZrfqcL8w9ilYMuDuDVcCK+WiQltLZfkv9/ESccb
R4Dy5pYNQPXde1SPqz2cf/CG57Rge+enWa9HgErhdox8vSrq7ega2Z768VqVaFmZ
qsAGbSPpxd5ADpXJBMsRq5Ds1UHZ4QPQVp7k9PvJAttLTb6Smuib0yvyTu/PD31w
c44EvPoaiurlRpcp4nsp7Kl6PCCJDnD5NjyvurDvND7nmfpS4ZGMeftQhyB8Lnc0
IcFC2MPybFJnPcfE2YYIVH6UWme5uSnVpttkNYBXyIH1ClRU/ANznDiSs+s+em/h
J71qHp7GAcadUgIQaD+3gd1LU0UXAikSwKds10cGSPOjh6+i6ET9B8VbkSejbH2R
6ZqD4PrrvX5wnugZY1iOm8XHDXW9uWPjps9c5HTYgtGmuE8uJW7R7aDYKbIuOPwy
MQW2/pfyXhI456reBAERLachcdJgbpdK0d6FVPV2HKkR2uMRpzmIcBWwagqAL3ov
Pp+7GrWjllT2kmXsrbOxAxNf9T40I61qJ9Qkxh/fBKnT7ZZTvi16032SCyZmgmtj
+oMyjhyPvNdknOWZjRy95vXv1penWCJjPzPtdqb3lhnnpWVdguE/NzQNLE2sPzZC
qKPMlhJDN8h26Y3Cq3KvYJFp814iOX9sAGB8VgWHJA9Gf5CH3/S06ZYcp2pUrgEU
vb8kWMoHp5paERDeI68ihf7ZJeLYHOIWBqY6TlSzmA0+oqDCILujLIuXvu3x95Qm
J9Mw2ELzAKtmgGVWOtgYJ84OadugTJ+VsREm+P0oc/JaNom5QMldIWrcWwJ/KzRa
NiCnbLq/kiySYvaExgZMe5nz363Fr27X6bjyvRHEGGOmoecBrtJ2Y3EMYVXPahjU
0s6keBJxT6Ro+ZdLc+9QWK6R3Hr9TeRYfqLlHw2H0zqgiOnkcrh0bQBWfxVfDxIq
4Ls5EYUxBNcf21vzcHIPuOue5mTR+E8pHdjkRnUo9WztTvAErPC4K9fofmSYXxoq
luc8Sox0iLogVWf3RAUGgALKoHUWX22GFQg6zJefmir9WKpI32oESkpPdVS+qVhA
OAzS8+xscruRenbQGgoJLn92XGygDvKlIETjW1BUtB+YNTPajp4wIC7Rnc6/1Y4W
FXAL5G1UO1xCRC2FIV0XI+FOavhx1Ghu52/TYrlExodFveNoe8+56VQs2Fjek74k
9wDf2HK9+jRYrQ9zRHGml98YSFJvMFXL+jy/Gw32+VE17Wt3Gl41UD4tLh/1Nk/d
ABo9VrEojPDUk/5K3oXjT3cBkqDJZT8dQuy1iaDRZ3a5zOEG2ZasNBdJ10+SkUN+
mixZId2SC/C+kntTZBE6NvSIDduSqhoWgjRhbVtbT0xE+kwJIMybF6N+xOG5nys/
XVZwaw3SMdFUPJh10pOw+vp3VJCT2uqQeG0uhOOiWPRkT4L1GH1GoifYJenAz6N3
MI2wjAAkJv2MW2urrJY490uHc6gRuOcb9VUPkmFgsAjVLCx0iwsjNwToIIGn3Hee
tp02drR9BRQevi+aycKSfjOaUAKGIYR/BgC7gPWyzroWkiT4hmWgn6UjrQOKvnCi
WHGIcvct60VuTVG39cCdU7jrl2JuEZY9RaXw+1Uq7yuFoUqK4u1oVzzRjVmr0ZiL
v9grIyTd4q6FqQy1D4TZ/H0du5irX3Z6vWeio6VoZuKdlcXB+3h+E+MHlUWS9ZlN
j1eTShIFuPr4dz6AAErxfrUvNH/OabUGomDVmf4T0F0wo4f1xGv4wVG9TM/XJgjC
tJ/Tf+vXCGQhlgLrGpTJpIEWIYWcbQhsFmfnkAmAItKhuWn+XLhztOXb+GI0RNi8
PApuL9it+CNZHdPL4qNxl8SCAGZ9FtUSvB6Yhuurr7cvSvECvfIarZZ1opKIHXyB
vu9m8hrTmB5rSje2JnVCI2xMcH5uSXbO2oMGb+4pCr076Bf54fdVwC5M58q+4G+B
Wu6pCLIuyzAgIgy5kJ1zHRRYBiDzZx6hMv9C/QNaftpoZFbNCXfbp/+UA0zb9QxA
wgdIYF+Bh5JNaHJ304mO2B0+9Tb5OcpXXOm3uQC0NKgyNyBSGHeph8042sMdJWET
sSbza4XZI2ifkTSYovcLCcGRxo5d0TAw0WLerpqOtb5Bk1VWScaczMBj92adWhqv
X/J3WGor951rnzAj7+nLy20m/jkzdmB1H6siYeJi08pX7KUTZcY1hJ0EKjyggxYb
5dO1Bf5EgaQPAnOAwD25BguiPM0WzsaXjqsWJ79eyjYqxh8z6SleCMqDYXjRMRWJ
qV2qpZ3+kiN15RanhTIkJcSx49+l7KyK3lyO5H31M8IAu4BxxXz/xH/4/r3b8jDO
J/WAL29/+jxxbVOlM5NJ0V/2rCxIt70HUUUGpaaQgUysUoZFskDVdwWqPrWY76vD
MIgR7Zh/8nGZm+mldWZgMqteJzpTmFY5OhMoGxgP7u+9bmfO6XpQJ/GCaS6YG6Yo
WVCyF1KV/k6LAIXA3+fUUrPSnOBZQ8Vu0Edb6j9q6jUiW+OwQUk8ZGvHBf9/NgfN
CnF5LJM2BOZtPoW4TjolwVGMSvHguwkQnEl/unQgq8ezsisUFtG8vgx0UoPICgqS
mA6Umxuc0RZbYnTCdfS8qUUL4IuwySg6NwARqP+NHRxa9FbXvln8ctkSmtdTanGj
HYcfy6fh/H7WF2a5iWdXSG1129stWIVpryoeO+79MVkeRWs7wwq3NNFZ2eDDChJI
WsGtVycD8IbmJmRo8U4sVBtHQFMEYyjgdbMTEjzwVd1ojBe4uya6bOy+mXOCObf+
Zt8dLr98SpWnPnROVRVaFKoNLLmFsy7dovomGDKwX5cmzTc7l6owFY2KDa8XmFJD
yyKSXP/1mrXXqbnGp79xuRB10B8BTT6Dorpxcyc8qhoMY4/K3knEmJmppnOY+rl6
IaiYY9eLF3SeydEff/QUQay7xzLsWKeecpgKqmHs1LIhd60y5E2sVS+fVm3fohFz
Qlw3JVZctCdvWqGkjcWBfAhO2gQitbapunMgPaAqlNOahclEycs5erCACdNgbvCM
4jJjTKnjzOG37k5w6cdv16iATF1Q36yzB+wo8675NVn0McfITqgJ57dKeiQ2SWvA
cVQg8Q4N/kaK4Oa8cuiAo7E5nHTlHUZtx8QSLzT4c7VmoeZkK4CBoOf3/UZ1M3Gy
2WwNrRf3sT5pRmO+q1eWB39LkXxoPqkME1EvuhGMEtmSLAVQeKz51HltIaAqoaMJ
dSKa2QTAAk0fklRwto35DgTf9hKA99+/5E00hMg3n9xXNyIR1Gm8jb8OwhvsXaHl
hIAoDZZbviCGhmw/trzVH+xxsv2fSDiZA+GTo0QCv/shzvZOR8lEiHsZqbpwNf9T
ZjzkcxSBM9R6qcr7jhByP9JEODceuA58yDsqutE3p8NKpDdJuA+goOUNmGJz8v3o
56mIDtV/uhfM9tQ4xrKhW5dtxw4VZDTTt4vA6kotOEMKHMBiISiJmodjemAQ/oHH
UXSbyrQ3Amnd2S2bH1jltRwKxxqkInk6sL8U9IWK0aTONE/c6RNHFvE9IQXbdPg8
U3VxJynhgBe3x0cH7z+Yvu7YMZhCiKJuzqaVKFcHJFSsLO6UMgA6rtcy1fqtiayu
lGkXwov+QvtIJuOIOO5x5/9z2grP6c2FceUUA5CbJ74lXZvb0E3es9zigLjDA6bF
c5mxpgabbJeT5G8eWLClLpXD68xfl4j7OnYKTwaaoIDM/WzboKaGfYdsCNZQZ5up
udOQkm33rKNaIgMVCQGm+gncj15mBeVHHG6f7ULazAp2T/olcf7qKj9mhgUToc2V
0Sl8OSFQ23S6f8sjF7ouUMI16E5q54hsqIs/N497rV5e/K5C1hYgcEilO2fcFZBk
UTIbBzKieydUhtGg/t+fqceP5a/4oFWM2JmzOgvbHKMlVBLT+MVrMDBjkA4BK9q4
TBASqMV33TChyXtleI76F8SHcBoETe8tAuy5yX5ofFkgb+dii+RachwUkGjA9d2K
QBnV2Lpc4zkW1cKXOGzaiQzLLTBx2WwpMUS0/yn43Hlu/RTCx/RGVducqSAgueA8
gkY1fh5CEAUdwp3pi9r0yipeMcgXmu8jvLI4UPRat6E+/D7vP0xN82FDzcwgPJbX
/5Of1cReaGEGAtHOCzqtiPZgoux3ML4awAlUMewoSkY1SeZV/Qg4Z6w2HS7e1gPk
koZDDkI/R9Q8oIU8gvuxE95DES1c6TazRn43d5393LelS5628WTbEuOgVVUDEgeo
4fyKn52JX/qDc6uTUk0Kj+Uk3PBPrcb5h1MXUFD4RVSfQyupguoWtcUwo4D/1ZKG
IR+DO1BUJMVufeiYrD63/eQ5aOxQ9Zbar71QQkCTXgNRrpE7WIg2sj5x7gefqI18
84DywtNKs/qL9MjvIug8W3kaHoMUlT+QsFDK4NY4YgsX8/gKmLwGrEgrQO0TZ/eg
mEOXRSPkXEoA3NQWj/mtDZhGEo47xU0pMD6gFIJ8pnFq1Qu7eKukzljxpaa7M0fC
VHOaKUkzSrZXFVZZKwYAzXOYUFvbZKJuEY8VAfwG0ci24t9yuSdmtWWWTpLFsHvx
ZUSGWj0RmM19ka0Yu7va/SDebeA7LKsUkI6sCTp4aPc3+NDLadUb6hs3CABXm22V
CcxBFwaL7+LpO7RbKNtp8nqRH3NOuVAV5k/ustPLAe/FxTKSVoyld3uh0LGSelF1
I/0WVRJaIqbLoyhFNq1feWwVX/MI0XbDei38x8MbR3Cs4RQDKjj7G8VytDTR+8tg
SsntIa5Fsb0z5CygBDHbD0Jj/gVcJxetnHyc/M0UsGO2otcXvcGwvONiZB8lnBE7
OwyqM7xeHgumPrRAT/0C8Nha5lB5ugwmKMT+hBm7EO3Insn8H2b1xgSad0ykHK14
V1IVFD8MA5gAHBCDmoL1VK7OW7vCSMTcmeG1SRsk3to+wKI+g+jeAATlYr+b5BM5
R6Avh+O0ODqKDF+mfVjYe11Lzmn9wVA17Wl83jXoPpmmuSwI7Iq/7zLXPUCcZn8x
Ok9qobzoUlRFr0llHV9vRFNg5Nm3drQDtqddrPfisqeRbLgreRbFFD6cS3u7msuu
BmOF9DMNIZWMTWmtnm164uptNVPIbUYyznlRQFt1ALWUC2ENcdOp50M+hS+aYhu9
dHcmbOU9z1pG6DdE5CIolGLxICzELfd4dQ7BfZUIZJflFUnmuGgxLT5wm/FV8SjR
5u5+Y30Q0lXxJuVKq03fLBrhX+Uj7ws/oaOHGsoV0pv/U+EkNJAdNnoFtWpivTJI
ah+Wb3kN9dI/QUjHzIC9Q4UccUXrHdHKp7gmA4IHv+W6aGLWLu87Q26rsxUQ3vRA
A537dIaUpUCh0Zf3MsX20IwJoqiw4T6eGiviWL0heVx+JdBQTpK2UaM2D3XLiFM3
j9afG5yqcdOLrS9K9psDvLQhHrUaiV2pvVtdBPF0EVn8VVxAzRhYF8INwge7LlNk
lEaOPX2eY3AR3nXknnSKeY85Ph9Sl2O/oPYYhZByjo+GDYK9KUYPJ2sNreQnO7DR
OU8BJt/3rWxyLsP40+ZLfkVrWM+U+O7cw9vatBo39JiVDfX0Akc4JwvEGa/0qnuj
WyE6fL+IoSJ4mYqxQuo+yuny1HsMMnjDVzlTZNMjb9rk0MwPH+Xb2g3lGjNdQGC4
35HN6TdVY3jdpb4S3ynaLe5icqhuVPlJdoBaJlOG0pMXclQnvcFqxb+MFRsa4Z8s
JYI/DANGlsGI8gRfAPWgpmvvlW3QkUAkvHmQc72QdbVLQq6/3SDbip9Qh9kyM8L9
qK9J74P+vSnaAeh27vCiVSfyYWtkqdz6uzQr0wSGY75lJDhzEEPv4JLadGMRApID
s27Ck+OGsn9D+wPReqhEUf9bx7TR3P/68ExrqFb41WJQEx8Fdv0xzPZg/X86u8Py
BeTWp0EtRBCbh/DKxmF6aRvoP+CfHBzzhf5OUf9xqZZ1olnWDASLdWpDyfLPyame
ieQm2h58cDb4JbTF0pdp88JZ1UDn0Dif5PLoSzjffOTYEFsFWQnwQau99lx1DysE
8amcCjBs8z3UqzLhYntA5UPq6c06EGfNg4rL3O/dv93GVxVwKhman1IpAD+Obhy7
q+l21da1I++z+7M+Rsu94F8TA/rIyLEBl12gadV7TY4Gc3JMFm9vkkxTP1hkL6LD
3XpN576v2TJTz+/H3CeLxjVtDaLCtISUs0viIIuFL5Y+/+Enh1AR+UcFmhjjFnSb
9CKBLwTSLhn/UorIfUDiUgG0Z7SQSQ5cdglrkzX0+H5K5sqKH7WdQqJFTnQt4YeF
DJtQ943y63RXWojGMqdoOPRSz1VBSkcHtoTKJeI5jgdEItIMV/9ViNRgziakdLZ+
lYX7hOkKoCLM1r/ZakAO4sindbb6DBLaGDnPyRahmpWNU9sH2fmeAUIRsvXIHzN0
2YG+RYHeEse+R1bcaUB4zh9LwFOksVLM4zfzinG+GgCXGg67sb2vuoeIQmVkVohK
QYEOArfIAzVUJQG19VN6XGoy7Qu4OY4o7VDVEfqwpJkhQ86lkxEUWvYOEIKqhzPY
pK7qm2gKGrs2GirP3SoU1WL6Tv69sCT2v88IWxLRpxLabGTtS/ykYO6gEzU/UyQJ
LAarhfgU8LiGCgjaln4+Tp5r0+3xcBZn5nR899bPBo/Q7hoAiNQF0oDAH5FZIiLd
HGOvv4G0k11ANGQzvHyfViE+u0eUo5KaO1G14r6s6EPC8xhcLGzE96UNkO2NupRA
PbvN9ucw3xqd2tslyqUSorVfdVFlBx4Z8eGlD6TgnVECx9J+CrwFhtU29S2Pb+4H
8MVd++2N0xuqMg+X4PQdmoxLCB+9nYci+r3zuNdfr6+O58FeiVVQI+VtjfJLiW28
FzJb6wATluIv/fyP9Ts0Ua4MKnGm+TTrIJrH4mKxHiiuGI5MuNvnb4mRbcdY1c+E
6s8LbzB1MN+AI+XbAsFjeYy5aUo7E1tbe61zigLJNJ8Z/ul3w4JamgEPtTV6Md2T
0BYR8HsElC5ipCiO6C+8RhZNhm2VTM+S3Mt8NlviwxnreY0qOwSdpniDYe1cIuXS
OAIZQ6pIHBYP+/BuukPqrzmDO1TygITJaHyZeYYWb43En2UZ/whEAfNc/SubjP2p
8CsQvsPHBvFzkvKKQ8+9de0eP/ppuudqxgJVu3ykU7b36mgQutStPxjlAL0EMbcg
JxTKDS+prDgidSVzqqQVObN3JlpY2wmaFqKo4j6a7WlDr7FVkxu/q6tFE5xGUIyj
Y/L/A3WuHn+m0/7MmjBluZVT8caYToOHtjC1L6oSDBo+VeTZWQpyjLA648Et577n
OXMlvaPucppyvjiEfp/oZFXcYYEitnOb/gArwHUhCoHGTlaQe0n/sFN0FUFaav0r
doGqUMZo+kr7BVW3Fb7d6v76VhVzO/pFOztcj+rMS7LPfDEnGV+GqZL30qGdndzr
LH0CwLjPQf1QAVb9Tbm09tSgaav11KP274pZNGjSC9INVihzHcCAl+eMBJB7VsYg
4iIPw/PwTCwrkNPaoocyqmWUjM7TKwupOQt5UcgcHQryj+fiyI/O9euLKgXVJysb
PTyU8z2j5/7OVDl8ZDvcyG+zva50jx8nSv576hN96aj8i5Y9qKqouH6RLbN/K7Z6
CcOifgr3Ev8GlBxwDoVJv2INnh5T4G9njf0zBx+nqs4QLJtD3k2zZsUEoYqaDxF4
WbjDjkXcCcwLwiu4Wifs8vUHZZ0viiQZbRQiKw+BYGdS4J0kJ8r1jtkbibh/qNA4
2P1q1XI3z5n81Ga9Hs3fAZzDGJPDuwNWwSJaeBLIawGYvhr9eLvGwMx7FsUkVA7D
YhQxmRa23h301Hlbx5kFzwoBOKP6g793uLwHx0S24//mIZvoQcVsHg8m8zNgNUdu
7k9M+qVuXeOgitqogMioXLrg59MbF4PbpZk89jZC98rj2FO4iBaqTKc09xMMzlQr
CVHJon04ywag0IfKFSFBiNEO/yQsH4u5dys/J15XERmCG/xQ13YlqMXoIYGh5Dnx
7QJiizL1RTBw1dL3CyvbYg/EJX74motY0zAIGMx8RQ9zvfwu1RvGH2BObZd2EHG5
dGg33M4tJ2xwKcDod/Dzqt87prsUevxuhuMW5jP7ENnH/E75NmxRczks1cmT8M75
jyS6XS5gJ/y22XC5yy6yjw4FHCvlaIub1XHqQmKD2Ma3TdbzkXidUuTg2kpWi7xm
GNulbV/CQLdxk0RPI/M7Fy5s8h8ON5dV6jsaVkyIGPQ=
`protect END_PROTECTED
