`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZ9fJJFux1DwgJrSZ/9mT4qiE+Snnb2y67F5MTMZ045fLaJjyJSoMjFkqJGC/Yzm
+JvsCt/pRI56FWLh7oZXinuXgCqZQKZyXPrjI1DsCbiz8Hk38kvNbor9AoJ/92HJ
nq8qfMFQhLYbPxk4MH6W1KLhEYFsjYMqwR2XYGMlM+sk6twODPaprEcZbTLu7a4H
s1NaLWAWggFEXioYUDGP+I5YJUy1mlLVldXw4yjq1tbbxmsGB4ZHF01A4rRP0jUQ
+DX4sI4f8FlHCfctXAwH8AiQxzmNeCAEoagIzeLrsrPXL86xHb0PWyfwEzsUC1qN
j6lRoUaODxIKJ4EFJrAI0MgeZAAB6BjiO95NmPCfI37oljdvrmLBi9oU+nr788ZS
BzTeWUz7l0vXd6shI7RteEb+k3RJ3f5NXQ0ys3Vmy9mamXAaLl3OLCTuf0xdonpK
daBpub9M2U+7686zfC8iXZWACuZu+PsMCvCq3ne42mAmuQNimx/PuLG8aq+m0++L
usFS+5TPn6Q9g5kLfCQ5F0orrOhBQPUMbMYQrYJPaKYdTf2aAYFPYgm6HAgNU/LK
8gsB2VpfsCRU6Gfh5AgGz7ECLKj1rfkmIacW+CW0wDBZxBFGIVhF/IF6SbSmEsmS
SgcLaP1JNAnFnwU8cqbG4DJBpDKUcaE2HRQrCygtFmb8DJhPcJs1SqUPk14Pl1Bt
p0w1D0U1CTZmSDArEJ8IlhG1LyQZNWrvP9QbPFStFmVCnA/OofHB2eU2buQ6n93i
h+QEe6s7QdCmKzSZWpqYDIK1K+FEhlovGMcIU4ABsSCrwi+2xy+/e6QhSBYL29Q6
EhEV8HkNFM1dZ15cTAUiNqgTQBq/zfQKYpPKYTgZC5Ssznjj8KnjNkp4gWw1T+ph
XiHGLgQWJqSLTI2Ihu3OiBj1RzUuZzbQbtc/qtzIPAeLxlkIQ9OI51cp+VXiERGR
rare4LaTM3wUaQ8eErgK/rT2I4I+ghEv39sz0glwnYyC2S2llUy3TOD/2hmvKadb
CPpFoZBdLD/MWcbFZHptFsGu99EHzGGkJcxc47SAtnlxOH9wtMBnAUmEnVzOfM6T
z0uPaLsp1wddtRaWiUUvJmA2UINlCM6GSwXk78giB8EsfcxC93IBZzUZLciCK1Bf
armMepflyd4nCRTBUH3oqtQn4i7845feq1fLIVtkt2PaYJiQMKE1cC/ggpeDEasd
lJXhSk0DwEeUap4y39tGEbQvJRYN4tdIArgoQw92PdsNocHf30g4ZclaYJ5jA+1e
3U1V4JwK9iTj/1C60CjifxNG86THB05+hENkjA4dAF31trXwOBF7rW75GADvmC6I
DDx4B8bBESdbz6uXmDEcVOIWq3oFhpHZQDntpntzQeEjF6l5x/+xaa0Uo8NasPru
rBQo4IjVGGKRw6kZU96L5ySStDTMPHWrMxw8UNKx28fcV6NmUkU47VIsl75OuIlb
SsxRi30cQ3uiFEX/2jph74X+VQjgQF0OWEihDLpCoHzBPKBGsWO7cPXzpGBSeKcb
QnBDD6/zUWdmKmbhHzcC8JZQgc1msvn6MhAYso2VqHOPmDuLsd/Z+PKKKVDNDfSB
xX0LEmEy5Xhgtq3A2CVCee+PwHsKfZWJQTFNe5o5AxISJZq3wVO2+G3zOSEFpETq
+v8NBnsAnRm8M3lqxj6B47gyw1W+kqwFjIK3tHzsic0gAEslZd5ZC0oGCF9jzuWw
FaXCZaaMAVRonBPXgvPNSCczRwxwzb/eoqNgxWwBarVBThsJGP7ak6hBmscNxszj
r4a3m0oyKfEeOjH0aCIZeRmPflnKPCtRd9KI/Wa2VIF9Xzb21MK1FFyL2QCvhy7q
inmmR5T8+KPAB8iR6bu9kiEpFdc1CtDyLERNdqAJDFrVs20Ej+1mrpeGZxXcgBGN
02TZ58I+zsWWI40W3QJ1n84rIx0/+V0Iw/msthKV9leQFw7tgyWbHGW+62nWhlqx
6EE8TkhEtMBYSOuQlwiJAB+UUR+Wi9NNNcuh4fx7J8VVa3e4B1nQ/DyMHKX77rBf
WuT0sRpS97ciBdIllYLYur+41DeEugJLzlmNBJy3LL6XXk0QSJUeoaqhLVmGpAVp
wBzQEaeNw90x/8+hjuodJ5s1LNMCd4/h4vSAPQXWSLISo9AYtZ2MTPGODphiB2Zz
T59eri1VgIlRxHZZkbqNtg/M3SMhC40oC/Z3uTbdVfkGS+VZ/vkY3AgQ5/x+239J
9dpsOjBwPNpVQI5gh1lIKTMqPv/hEkerVuA/pznEaBB27c5COj+M4H3DU2TDGT12
nSAY9+we/dP6UO2M3Gj+8FcxjDVtPlMP2y1pz6u5r50QighuuoDGOiPclGAmZaMN
sCMuPFFviK7GFmrLmJpJ+QEUIx32jn5Fk9waOubuD2JrN4JQqkYke9bklDQxMoOj
1v88s2P43RXtEkVbu7Ugrz6j29cBcVbMA4zkmEpN1QnSdtOTlnJcKUSUxC9dKi22
SgNHZqScHF9WPpZ8T4Sjke6OcH5lyT4CLVkrJD3qdCnzxQXVHg/kLgM7cBsWn/M+
UOTJwiuh1U/wFD/v145mNgaGArRWZBhKek5Kyn9V7G0ZuVZtm+EBz9eLlvxziIpy
kWrqP/av5fL8tZ8TW7VSY4qjRdmF3tRQpFhFn294LtwqgMrfCB3Mid0R+zr5SSkG
VDaUBeh69xgV4IwXD+x/GCcnA+j+7L38hT/tHmdG9ZrJg/QAy7sgRtYgbCtgdjy+
NZNvR6p97Dam2HnyHYemPSG5pUD2AkItT2dhH3rNjryG7pmdQmcX2lroU6G1pe92
`protect END_PROTECTED
