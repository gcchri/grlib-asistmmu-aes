`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yuAbOmZUi0SEv61ZoGGSv8leE0GeqWD/dXeLMXF8T8DjNZiyvQBnBa5yojNlTeX8
cthozwYdiQX/4DxmheTI+iLwGExnDaApf3h8ZRASJbFp4Jm02P8e6GM5vAvtWwIN
OiE36xWNLT68aq3WsK3mu+OFk9ZfdYfEGZ8YMoeSpJ5nSYZpfxP2dkm/m9RO/4gs
d9ARoAQ7EU0ZasLV+MfdY/uslojiVYs3BkZmYA3RH35bkt9yC3p8wKp5VdJR9Mxr
63lY8apauSoosVtLgmYv2YHlQG8Jw9EgQmnVNVvuQjnc2uCZs6p2iRDO48U+qP3y
BeJUZ6scDN7AOgQfKT6HqyRxWKvQSGsvFeBbI9///Gdnz9Qy9+dEXenyZ7v1aBto
sJh4+vBrzhGGsJNwIi+4Zi1tP7w3j1FaLSn58yz1VCKnc5aP3qd+Ru7iReKZDO46
vv/sDwB46YgJMX3gxvdEErF+42vtg3psRW9GlbJj4E98vyDlk9+YZgVdrG3Izca4
x1Xpv7mUR8M6h9zoYY+6KtftPuuUbpVE3Gyy4Z3C6Rh6CuN5ArOtgDqoVP5QJGku
ykJb8+exT5M52MQnxjQ1NCeyp1Oyl9GtzZeM1n6YpgtSaSAozj8wtkp1jy1FTYPy
6lTTsyu26i1hK/bm0OohQA==
`protect END_PROTECTED
