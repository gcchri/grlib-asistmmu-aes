`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v81YCLDdarmO5EQMujjlxq3A/ytw6XwmRd0xSWLcrJu1un+DnAWGV0esso5YnOrI
EZXgwR+jgqKGK8hfQ6+oGuqZ1/EY5l6Tkz5kkwjsQxB3vIJBoYeXVji1M+YHeFwD
iJ/3B0o1oIofkIuFsg9I1GZLXA+atO4lJUw51DAcyg2gWlMgwLMmDL69XQLV8QRw
cv5FyBmCwl7Bqrg7NzOXkXxA2yZmoExcq9oP+Q3H410W3X8fuEwXARKeGLTMW0UJ
g9U4WzhjZwFK0yRaqWeyakOi/MBqWbJn3XARVgkJ/R9fYv7pQPksshbcEulne+OF
KgbXuv8Iz0OlbMc+uckaZEHI+pPKhLPAzlvQ1hZ7+Za6I5Ou7TwDysTlaSurIbdn
e0goz0UeQJzqB3fiWeCfFtCI2dDgpU1+BATHjSASBj6irnUK+EH7mf73PnZIflBU
Aptr7AuP7MPpnmoOhWa471L/ULKQSTRMWXYnlc6KhvhiTIvA2B+AEdqIJn80N2Vy
39i/lgZOHIAg6F5X8xkKI9e/cPpGVM2la/5Gcz+aU+8TlpCPYDfX3IjZEV6ZEagE
`protect END_PROTECTED
