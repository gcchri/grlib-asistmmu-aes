`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PN9cGT6qPCSKTagMOBMI34MSabrbwPkaN0D/C3TlvgWoz5FSJZfDbXxhL9xDHQR1
pd6wZUU+jTyLK20skfagT8hVwSN6SYxrLLn8iiDFnMu7FZHyLgVRgsaLYROHhjIH
QFuE0nG+oQU+ncyQomZlc8ag97KQcwf+vmN5eil0TgIPnuIREUCLxTUgyTWJJ4Er
8KAwh5hLmoOeIPIj5Zty+ma76cFYwSmvrIuYPr+EKbFYTXeGHruIxaKESPuOyBy9
nCKhUjy9FtFp4o5DxbLN/JcBDs5STfJBLOaZpqqQClSUp2phXVTPL1P4T6t/3+I2
Ic2oSy9zmbpGBbEhQC8p3ptyd8jYHZzgPYMy5ir1JvX67uXgCgZ+JNH09zhsZ5hv
SmIkaRn9ffnVQi+Ct/yLeyeZz2UR1O3TE54vSymOg4Q=
`protect END_PROTECTED
