`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fwnocUsyt3IsTG1xEvb46zjEQzXpAK+mTgonA+MuNIvq9iIfijqOEehFog6LuhF
9lqsVK/uf/fjFyw+/egkxGsSbrIJctdKpJLA2jkiKjIMbD0m2relyF1X0ZJbOnZd
hiWiqhe9kt4osDM6XI3VStF2wnXGGdLa5t1a8k3ypuilXRaIWfErjxEX02UymDG1
QZXQ8hO9TCPQRz/SdgmUt+dT4yBgCCqn5pQRMxgZr77+13nqo8hP2stV/DC/QHP7
j5UJ7T/55ciafPn19dfqhCHn8Ga3riwcKVd6Ul7fUFiRpkXQ+AGNSEM4GDwnRLyF
0Qf+MAvEr9oWeH16OZqJh+h4y41f1qwF47Utffv2ThVmCVAJmeZ/+9rTWRtOSz3o
FSvxEjhDROHIcDgCZfcCxFItPNaL4yyMDcrOMm9/1HGZnflnG50Z++OOSl86vejb
i3d79AY1QgGEI0RT0EkzL6bdIDIRTorq/9KxdU/Jnzd6F9zujYC459wcngw08fRn
WXzSSjxPwXy6RIEyhPq+xmCXqxGrWBgMLs62kgf5kJ/I9wnS7zbyA1hYZqhQV94Y
DNfh4gZ6Hp7AcoaeD/IDXQ==
`protect END_PROTECTED
