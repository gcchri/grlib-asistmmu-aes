`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EVzeOz5dMVSaS/TQdSD0b5fLidM+BhDZfeyho41HLtI9pnjC/ZAj3VoBIF7j0ozD
E/1visJO6w17m/vcvJN5F4Qe5csZZwQ/q9Xw3ZDD/Cc9TMRNGIXGI6bhC6jYXvk8
rP5xqtgs8nDJhZ/sl+arxolHT5DBBSmwxpD5YPY3qzr7ZUvzPUqL1Ar3tE/t4cba
6MV1Gk3vQefLbTwxAtnjiGixMSky7UvgBNvcN6SwTGkbAqpPxj/+qAKkPMwizvFh
Ck+vIt3T9e+3jdy83jUrDQ==
`protect END_PROTECTED
