`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ykhadd+Hwyo5tdNWpX37Zxi1rLjkQ+hNsI0c/F3Ns2kweABWMtvTCmhlmSsCmmiZ
+fCOJzMu/uLhmb95BhKGrV0dM1e8F+GKLZz5Cy+W64ZoS4CVww3c9mLEevMJoszH
fygy0pb0l3G7EX+L8VZ4+X1TmfJjCNcWWQaB7asyNu8BOfpqNxjlAfwRsUJIlUCk
pshkoyGH+DN8pDd4poDYCYQACSK2jVCyQRfMi3IawKjHV4b6WJF6tTcLz6qwcvd5
PDVGj5imsFLe4hZvmUV6reiCdL5VsK+uUm9P5Xn4ilDqZe3CEhkFrQsyvGOpklEN
oOMoxKxhqv/H1JLNaYBWzzuY6jMoJxw+9UgfrCF2JwQ+N1RA7pHR3W+CDLzWerVo
3iYn8yw8krdDW1d5GjCrcg==
`protect END_PROTECTED
