`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
05dPahQU/1hgxWvjChavsQ8XDDb05wjl9NP4JfhBLpKz58ytd8eT4ZDof+cz4jOz
3ZqIKGqbB7HChynbAa/kEXTEfi95zF83V8OsWchwItmhA+AaZnbLFZVi9s12+3w2
+fjANN7ADwo1gE/bgtLFJiRxSwUIPgv2edPpiyZbpPxO5FHlWg129m9IiLjp8/7y
l5BQaFJr3FYDfhXjNXNdgQ3PldtKVzagdJfonBFgSnutOr1cHVDb1Uzzq3ZxJk4x
`protect END_PROTECTED
