`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q0f0wZPZ9n9SpiYAeQww/7WLLAnH1pz5LcBkGO3iJUF98fVUOOqN36J73qIisneU
1MN8Qa0401bT5z7tBYTCosrgDEAMsZxgmUhkne9JroDBUkmE7H5XFqjMUffVycp8
vUzeVnkNM1um95OUw63AoKDqmFP7hOM0lCM/c8Y4UsOOo/kZDBefQaNtu4lcxtAD
GChTUpV1Bb3iJUhvBQDJdZUkhvCHm6V5W9Tv0Tg9WTNMjQhGv/3GSv3Udag6C7tE
pLfkiZ1oxqT65bzo9juWlp+LYJP2PgLCfpoT5QGu2jr1GU7tQcNANE/0UCS7me7h
TGMxJ61OtEEv9es+nUARO2Qti6wcszqPNehH1fCa4RmHOJ8TkeskyvjoCqvX98lj
AnZuIlOE9Hp7986JDfHk/mfazZBA6Cv5q2In43LY6v0wgrZ/igZt9OpzpEumygH9
`protect END_PROTECTED
