`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgOPVVqvnepzJx88kMOf6N8L6Sdfmt9swoHJ39pEWXkaQ0qXo6np/kqbtYgpc6at
x6oxnODTk71d+IxF/5/Q4668AbOynln6DfevaMaROljaRxzGYiTxm46gsSyVX1Y2
KC+jdzHyCfI8D0BLR9fSflSVQzn//CP0NZQCElTOZjZHplKG1QaAvOGWS8zJ3mYh
d/n/HAi/A/1o6HoV2BWxg/76U+kGTVb9MhstB6Rvrql3NDE73EH3X4+aA4EssOhx
DBrnKRwpI1tcHdY+3VBhubmOF67tYckqiJ2ueAp/gPDn7fJ4PcQSZgzXopqmRuOe
RLav2lMxxqw99YJo/ZTY/HOk41ECI4QIuYK25EMloiuyvDeTu3B71dPN2yTQvNvj
o+l6DtU1XXYElUliKn+2Yf8arr9V74sDiKfotQik+cJ2vE+fZOVwOOXGr6UjnWlH
5t6kNH/sXcKPMQZrpnEmqtUQHBrDslLdo1mfyLR+qCU=
`protect END_PROTECTED
