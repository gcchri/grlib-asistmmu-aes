`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAXKg885snShHxSaNooITkJ9v2vTQq+M1bA27QGE0MFGVXDfn54Ufx9bdM/IBF2F
wUTALArWuy0b+412Cj/gEUjInC3bx0C8Xk8RNh4gUfKIGlsevSSpQlLAxrs9hIUz
uxjImZtgB3Gn1P5fWY6J7pDBYDK+84XokfLOZLOyExUUh7DtN3DGpYYED66eg/pO
jf3N93+LyaZns5WSbN8sAcE4/5/HFuzFrhv78wXB9UNcT89XZuyftZQjleeoOoRz
/1ebjk7G2wNLTsP8WcaOxzZTwt4Z+jhisyLF2LutYDG1GtzJTIVIVhl+bavQyAy6
PjG7bW+Z1ucWHpbTNwnfiqWUDh6KPGcuwuv2zuFzjGmeytFTUShcCz/oXk1/80Zy
uC7FVXDmUhL9wpb+zJjxLscIO0b5Hapff3qzVAmJEjx7jngszyg8hZLEIrcn2PcU
OeSKbwTrYYC0ASBH03qNkVgzr7l3V3fDc+nb94pgSZq8bl8bqrpX2ooTounXVlrm
tUh6n25huzRtaqIf4U79uy0TvOSQRZt+hdiknBGBvXV7rdYAmMTb/vZfF+rtbBG8
BPRE1flo1eGoYLFpgw0NmrCxwtE8j3VeSSL87VBROU0Litgyfu1xqs37OKaOy1Hx
v7oAjIfH1pUjjiPUvCeJdISQ+Ae3Vr/d1QEBJRcCrE/HlpDAqHHm70p3kCck16dn
Dy6TWSVT72V/efch12GOvRyj7zBPpL8jTkDkriXkGFVNvSk7ncmmfnNbUzMEppyG
RVQp5CA0mWLKegOePygxD8wAZRNIF1zkJeqtuxsRXE/0PG7I0hbqebcZA5eij2FG
bMPyli+rKtOUhKQsQyLf4hZyzazIDDTx54svcu9MJDDR3pmAGPz/uZjNkFHqZqsW
OcVSq9vhk22QBTgZSpEbvR8XV/OrL3/Vw/zXlKvCoiGihKL92QwxA1KEy++9AD+y
JzO6/u60zIVrtRDrN5itxOzBgJK0HBcatxU4Cro+lv5r0o2ov9mUYic07uOxDylq
L0ydQczQtnZreJZNI9WQonpsOap9H+i9aoi3lnSrNO1Q7bDL/nzKQ+mJD24kQ4iJ
XItYzQ6sPcFMukz3GkFZpDL0OyETTSY6jtt/x4imIqVDtMLTkyfP4qeBk3xvsTsF
sR8b1u+fp63X2yhpZKpMlMY85pqNvvDPdJ5nFvSwe4ADcPwwXxBNdCDd3HBKCv+g
p0NBYkiDuEGneNwfCi3qKA/UURPbWBrrDFqYOhgwAihgomKrLxLOrLWW/rVtxIWn
wkCC4s4Q8hwbXjkd85h6dWFpr5APm7QRBsVTWprdu/OUaEeetKK/0+mNQqeLc1yD
hzlTG1lU+YAQhwAoKAxGO0IZ4e/3fLfWMKgwM8krbI3awoUsGEmhfApcNwqaOlNj
jmaIdNl45G8w3wn+974ZWUI4DpcfLcXrakPt4ptc5D7FpiRo7PqDqvMEzbjcHE4d
tlFHaJQaEgJvaWPsDBVPWtWvpvEI4RyXuuokN/zZw2TQhj5ksTHCA+gA1vV+6G6N
QWdPMQVNpJ1m9Xca/OPsbgWRFUf4KUE1xontib4lygSzMkRPdSrn1REAbyAtNib3
eTRFOCoRva5WgiSOt70g6BdECadOzRfKwFzEmm+RXaUgdYnkGML74JQveTXa2S+w
xJ3r+AMEiDABHKqvsItPz5Lfk/+qd5ZErVONsclahAFtALXiJpq2gK9VnZnaYBrt
Cbe2o/8C+H4vRMcYiCi+P21iHpepNNjWN8b7AdrdwXTsQCRizEUN8/hjjwQ5dtLP
rOyfK2AwbbkDTW+csE7yHafw08QJFUaj5PVl6Mdk/E9lHrQGcqC3b6Ju7BCHyQT2
MhvQx+Fs+U67BBjCi6hwddJPfRDO9o6Mhcqi2Gin/wgCKpmiGYUXXWkWv/DYHMFq
0Na1Ix3JVP5IVu+vnWHW938vS4Q2KzFW/uW4qOScnDGbKRHSQq4nLmUkI6i8S5mB
Bkd6o2SOjqHjRxGxJJchtUSsEv1pB7doLmlmPRNJNfs5RYNx3vZ1VReOAYChSQJQ
guL2R7uyH787WE2UCgfG09iq7VHMRrXqxhFslkA4cZ0FlxSz8BdZOdw5t7B+Y2in
vyV0bCzWbpW6vAj47nHvebsR2lhXQoXz4AJp5LcfxO7wXXeWdRa91oUtLbT0KnMh
BducCrV4uD/bl6axhuf1NwlRtiLEhIx5bqSYzh9ej6pu4ElxkF9o4uD4whbmtcoB
dh8EWGwfcguzfXryorZnUtbuxCcIq7vsxJoKnS9N8XzkJapCng8QSLy6wSLZFaVd
7PxIrE7L5vSvJLxY+z+tfa8T/EJ/K4htNJOR1AqxiU+AM9cB6cCu2Y8/9NFfwBDh
JjQrPhZIMrGTq/DECwVxwCb24kRBk+/6T5iRjXlPXZDwX3fnF4ERrNT2+aYGD5KP
8WxAzTpvfEeC410EzGf0Ev/61I9iG/ki3miN3+cW8Eb/ukd5+Y+7NlOJBent+QyB
k8sq/0nSRnd/HJDhbCGCTmz63gAopx9bH5dkWALrL/4P1PZPJQowAJ4cGw6ioeef
jLpXQ4AOUEcrYDGteYtdj7VYD76zkr7E8Y7+/1BiCLH5spkEAqZ0ij3WcAL18p2J
PTDrZP29Qv6VO5l1fndW4Uwtd5RCLEXMEdNVa684DUb9cyvHgSeCO8j3L/5KxGFg
+eg7F/g43SF8ZE0vnIqZ41WKQAUVpVuhAu/4JRJJyNHlW1xDKTcBwPjdbRY5K9Hw
svUbJLLkSauMXktQ3HUZtjKlpe50IDAAJr0/Mprp3YNqZAztFkDfdCgUIijGMtob
Hg9SI+uB3SQh7tmiawTJz3pfNqYymEX4A9cnQggB2Q1WaBtn+lPvALcpmuYei0yc
KeX07f/Bj3DR8fZA0oKRvSBjphJfrfS+Zx2VxN5vz+/O4Wh6fwzHcKtukI0hntyz
b6/lTP5a9HkzTqTpMqLFD8lzU8TQweCtmR6xMKPQte5olOQnkISn2kDzU7Lsp+hL
KbsxRTc1R+pQZsWfx5h9MRfAtzRbY+CKu5D14ZDE0BJ8d16pPw9R+NUeRjJZoxhW
5hSCD6vvyVBJOep9HHZH/z+Eh/IoEsNDWeT5dXxG6bMAXCjQMmJXmufunlcVpnam
np11ZOPQ2QZxPfabGXKquxCJV1zv045C0tr9M5pIDHdgYqhL5NGViY8QXZYPxpE7
VK7pHM1/0S5jj2rXlYQX4ztkBoneUr5cEKHjuwc67OAtXA29KuwgvX77sy7Qf3b+
vSAHmmBpbJqAKJrxpLuA3NhQSRy8JGDtzPHHXwLtOu20hk8tES7+z644c8J8M9HX
Kj2SkgNGdDbfq2xavtTFveGJKXOGcU27A48eXmhtTI7FWRtvPpdR3RbNmkWnfbgH
F6fiw58UmHOozcP4/ahqdecIiP9n1Ea2kkcHAON3260KC1mm/vCn+kI4BBbU23Um
dreOCxsE4IAuGByT7D57fAltMq++LyHE5qW+QdvyAitfhBwNnA7lmBPF+E5O0jqO
G7dWBLNYEBd9MqCSmwDiWqmMRpvCg0OCwh3reBM5yJIXR59hDcdEHqIWchnon633
zzkCV0vd2Z68JHWzcgb+fSQhd6mee9spO8LsWr8gv8+NH/HM8ysBeUAXH/x0oZ01
P5rZY3xMPOli+dQ8lnGCm5tzTzGn6zARV4Vk6NzkRBc4kX5Ew8c6STFv2IWYkpn5
69tyUfwIfkvZxykSuAwka9S2sJX/i1xlZ5NVS8vUYjNUKCWqyjCkH1gDtG2P30Cw
xpCuK/HV4tnazk57lKarqTd2AEL1XoxH+8KjFXGn/YOlHeQ41tFv20FQqbX793hF
52FQzvRgyhzA72qCQHgcgUlzqlu92b1IsbBQXAxeN15T+7t8DGmDzBJ34XAWXrF5
IoK60TjDQ4UtsA3l7mFF5kHkyJuUFL5aMVli/gdvLV7sUjxkJYUoMtsZra/nIV5W
L+ZAsh/EqLbwKxo5BSACQzaXOBzZPjjz8nb3PBkolUe6WBy6pyRs8i0sRBPYlsqw
gtLoyNBDQTJ89a2Pb5GrqStXgWO0z31pHjgJFVYMug5nOMh8PkEnxz5tGS8qk7Og
iart73Q+yXEwu6s49gA5iQFhPtvAMIDPstpC29Wkmpa8F/X1yaEIT7PUsjuwRYF7
l/4D7ZgKSktNEP7oiIpJqjPePLEln2cGCNFlsHE+L0aToVK3JpZOAJ4XMIvgCCdy
Gr6tfR/BuYS96RTJcz3PKmm5Oj/VDv+OfalX+REuyiRVKookd0Z2hZT1aEhut8pP
vSoz0EIqiUC3XABOtEP8GiZyAFBnTIGk23JUxRNVChDaBZiaTrV9p48RS+Klz+0d
oEECXZihoWUkYrkROBtPY87fkjEIUvFwIWdOGNhscPEdPdxcNBHU3OIIBmlWU/XO
k1La2TW7a/8zYk6RLvCDecYBW6QkIzhvBmo0Nc17yRgbAF5fCMIHTdW1oNXnkYU5
b9I/xWRQEHiYohe5JjxMwLEomWhZMNzlJvhDgzlhFRPqoy7QCJx4Q+L0Oz/mmVFl
PTzpdMuoIyX6AdEhbZfapfAKC9DrZkHKicA9nVoTNE9AnzXATaK0P5DbSlHVC4Gp
EXhPvD+LZxSHQg6ZNoQehQVDOExG78OEbFh2RRB8IsoNI5mRh0hzPhRf+GvWII80
n8wV+ORupfCywieq0Qw5OHCSw6Iy3FWJZ1pRZ6oR3ep4eLNZvDGCsbHtU3cHIVu4
fbb62YEr5ymzVw8kFLS74Q33AjMFa0/aSPipGzx+WoktQiHpHn9YBbUN8Pz6Lv37
MMxrip/KGRDlbgkdHGKGd1ofTSFfkJH32XQB2/AxKrgbGSl7iwFS2vWeGAQ1+/gG
xz9r4siHeKf9BXIyVNPRqjVcjSNKfnfofEyjMFJY3Wv0AXAgjPR7TYZZvffF8i/k
gjQvS1s76d+nYA9grj5aj5bjvXlv5RMPYKwatpoXgF25D9r1gp+WNRyjwDTCPqwW
zM07zZG3CYsUQiNLGceIsT2RA5x5EiAv8uOY2w1yuNYeEhov0BanLx7QffRQYhND
MOnhueJ3y/gW6JUWn9eWxg+M7rc6sKxo3i5TRBriDJpVNAdMsbUGXREmmh6iFTzw
5ZOVk0D6zVC+g40w/XTkSNHye3p696L51a0K3Y7te+ZXfPl5GnecsKrGX/zdfpxu
XBdedF6afnJHkdL2WCX/osISRQngD/S9MZIbx0IfsplAICyL1aONieVWEM8ak5Cv
wZFTaZNFpNnCeYigpIWMk9cYPqt5EQZNgylIJmjvERZnxcAWtwZ0RNBfAVeMLWbt
BZIzh8dy/kvvW3a5acStT24ArsFtHyWzJ269w1TXUVj1aztJdIQ7Ahovp9jizS0o
AyRwXi+mh0VXx3PaRNmaA+7z3h9Tq58nj6lyYYaNOMgKXd4szHxZpKr1+Jk7BC8I
DQUu68+XWEkBoAVrE/aajfWrZz0LnHU9xFbuBKxS5Pbs0yQUvFIyXlbfnLvF+iv4
jogXuuAwG+RXd+x0WQ+4Adz9IJBLEEmxRRScRUiAsDGcpvAAFBY1XoKcIX5ltdvz
1mWEVZ6Lok2qRDp+dHhwjcExErsAex0Ct10x6w2KWCt+m1XktNu+6cF1UWSMsBx2
MVJqzp9+6vcHasI1tSdE6cQXTKZMfA87Q1GG00KxF2VB1rPgS1VRod7ntQV59W7z
bRoOA0mGsRQfZX/KhLW/f8z8XEcJ3WQ8uHZxKAPqI70syyBw8qsMa9wNJh0YDnCp
qe2XN7d1Ffne45wQ98Wfi8Dxdv9vfOIUcbE98UZSv0B4KKwvmNflfn6W75+5uh4E
BGgnNP+Hh5tWDS6p1WvmdBG2S/SB52gPO67CAIFIUBHaoLRPqpe7vgEBVLEaNorP
8/pFda7QHw09tmiIx0CrksW1U9+3Ih0MINxliw/9p0KOik2QqLa3F3jNb7+/KJBW
GieGCG+OFwbgJ9q4QBGF22j7OE8Pr7EXEx9sWIsVFUNkf7V3sAkZl4kxPZjfcmVa
/bUCYoDu9kMbI6u8mWoYdw==
`protect END_PROTECTED
