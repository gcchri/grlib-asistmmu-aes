`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTVxSzvD+8RuLUqq12PJ670Y0fyT1IyCMSWtcDt9G67RN3ru3Zvry9nblX+gJP3Z
9RTKgIcEP6quRwt4pkLrdoP4t0RQhJuCqmohj8+a3OQH9acEg57fRpQXhSlz9Mq7
Yfjgq+5jPtLaRF++b7YBrzPWWUIwocxjwUiVvi+i3l9Irz5yUk/4I2dG7ojwpvFX
rilRzflpNWtF/2kZiXkoWiTkAQdqOTbMyChLliiDCuB1KNaj3jwb7qwS2UyJDHHE
staGgIElQBrkUaB7+IOWhay6F+ba7WE0XVQL8AzzA20OOq6XuOQjRNAfxThtbE5e
W8+3GGwnIR6DbZ2Z8psDkyH1P40J6vGl3HoPcXi/QWNIN7gs0AhfUt8pJENgKXYx
ZeewQKW7nnWcBBe0iZY4iyjuLh3SXuWesxRb0ETVLR1iSWqr9kbtqO8RhH2V9yma
718VfWAULgQKcu6IGxK2oK4HjaUvPUrj+NOL3wETIx1LEHX2vK3VjORNEgH8P9m4
hpU4g+iF6IkNxFjOfAm624+54AMj8RdKbBsxYVN+kwJKbFLkfehiA6xYc8KZCOSE
juNqqh2jub120Sz1+Ym73sK9Eo+353lp3hypydTD9Bl/kUx5lzD066JPf1oxtWIF
EOhdYE5GtXpjd1fQ0nK6LODglTpVEidBvA/DnGXUhcASkDl8Pz1t/PxNiitdhFhL
vnNBcwPnFTFRoaFvztqBn1Wa3gnBJ++nxu/WUzzzowJ3uAU867pK7R9vAW9+LEla
Jb095VsXOig00bdpubEdMFzw+2SAwbCYzOMqc9QEUWo=
`protect END_PROTECTED
