`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Ndsj+2M7BNgDJneFhYopd6rEVKXj9xADLJyQIpZY3uvP55Frf6RnsfUDjc14U5l
QAmcXEybOqoEV5IRxLD0dnZKxyYDusJwZN7b82ni9wCtaLCH1K8pAy+2rhTLUBQz
G3hIOf2pSrlCIxdzXY/3TdfnHskx2mxpMTuWKxRODg4BczBSoFb5EE3nNLX50Ez0
5QCzgtUU6O0Rbyv6/Etp+lX+LEwzytySE5PoAQ0MocOMCsUjTHlS5kN+uKpiVFcv
kLbeiBtIu9mkssb1mfI6NC6d7hOR9A78pYPDUQufE3kkk8dZkqEQXdRW1Rt/p8vH
JpFb2TzYLlB7BpMM2tHvaBazza7ca3xvFThsGJYdKQ2TWITkgp1C1MrZqLPTFn+k
0FdrMntUp9j28fRmxMZeue3pBXMi8DLUmJkI8ivz6V6+iM1GICRu7er6bLS2Xbyn
ZNRx5CrVBGpituMtr6WLxMEOh54aFSNeRnmFbav0WfsAJ2VjL3WKy14xsByVibk0
JTMY+ajjVtzcLyK8itjxYKOQ10JJqUWu7BkNLV0iLjHTquI3k0cEtrsNhbZ7xdaH
2IWSfXtoN3/1sfesvgrptsCbBVbq6PSSLL6ibbe24GHT0JSeQghJXgQi7hgQ2zYU
lPN0o9x/6nWN77VJBZQoYTxI7njjYqCX2P81BEalBmM=
`protect END_PROTECTED
