`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fypPQBYlLbHO1YN97XbfIXvYVGvXac3jnLjOz19Jy0zBtBvdiNsk7a78Qr2PyV9G
/GihoXT+VvFJ8B8atZexA9mb8R5DyaHYTOMgr68wPkiatbDujgA/57u2aHnHLXvp
gbvLySFF3QsnImJ52pIoYeqRqDLp24f7+hFqNQMzka8r+9dyMRldVvVe9NiFkLp3
t+VDasCi1bgwHXllO/zFKzg2jsHv3VK6T9u9zGv54JeFOWV2Jd0yxHALx3wPQRvt
fKt044pWfNwDPV/GagV6blQDhaIXxUx3j8/0YGgYT5BhI4rqTHRxBY2cwIABiZdV
TM6JhTd3uigZr3TWZ+BkrY1aLiJQNES+HE9PXxlPxRE9aXMpHBZat5KCH6fHdStd
ObPqvlGQC5qFgIqK1VHISSWRFc3O3q0q3pbGhg8/XBlczXnigzWn1f6Yd/PsD8N/
cUBevLb+zA9W1MUrUMobkMr8EGgsqLeHC7fvObbjHwYjtSEAAX92Ry1lxS/+AZpM
jhKob8NSPiBQz0b7wc6LGCIRRcyVVqe1XHR0t8AedvH/tGFrcGC+cSxSzwi6UDHi
`protect END_PROTECTED
