`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E+YBKEEBrXcSqtJXOAaAuWP9k6c43a0bSlb1RP5UHDuetg8aRIvtDiTUzqYqUyo7
csWfcLcDYE7j8D27E+mKlAxRSLd3xebipKgjDQyb3Zbv/lOz0d3sCkVWkkGfprIX
vCnnt0r4F3g9P1WWsyGsVWVyDiRYGEne9OxF6zpurcfAElUeDB0GTL6HJs47/fmy
J6F9EwD8kOrZ9O5+M9mcFfOOWk1Z5LuY22Xegyzk0HPuD5BhzvUI+7x6UW6UC6lk
Ykt3ucZcPdH2QHo0ztmplx2qJyjS5/bM/O+6X6mB8snC6EWnbQhifosHGOf0r0S+
rpgHl5fppPEZjgDL3YNTC7a80xlbWFA+rfh8yHNH3d043QPub1/dPgeyi2xKToOC
ecE4YbEAOpEsaSnOS4pWrqpV6WqbxmujJtkRv7tJcxvgMneoStOFGlc/9r7cRN8t
JeXugb/9iAxG+7SzJwoE6Tj6pIPlmXzINyw9OfNn1SJjAP2mT9x+x2nD9ZEq3nco
93y/vld6qNOlj9Lc22TvlN2JQ1ulAdrEmrAnE3Fu3tilg6LtWy9uRnVPeLo+tBPw
7SuZSM0eiKNL9UuBgQppQA==
`protect END_PROTECTED
