`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9l9nLhto/9Z6vuG/HZ0gRPYzgrOb6HqSpuN+FTf2d59st636caE5yUGjmKkS245
SEu7GMNak0bW0PztVgC1oUxK/O5w+JGQGJos5FBlinm+PSN7H+nop6Fm7oBr3UPy
IrJzw/l/UUKHe9gqzGP6HaoqxuHgEUHkYhFDNoznGyzH+SSXipfi3U5U3xM879II
nOU5heRLltAPcHGnqonz7ekBF0JANRsTU22LnJJCw1AGuM5c5Uwgnrj7kUqzbgJA
TQsBsyrEOW74ugUKdREJ1g==
`protect END_PROTECTED
