`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9qWQN0RWEAfuMXvnZOnyA4STOD+FiZSAzU2kgoWMxvG2heI5jrc4avJ9KKKlZC44
6I/IvVynqtDioZS3+iHFTVNX7EFJOwgQ7xdeJuFrR5y5sZ3Bl7j35baSjZWNF+P5
fog0QEqOlhzk+YFjFojMm8jI3lOZo2p3yelTqjk/l9CXxxSY/F8rtRgY2hfoCURA
UeAjj4WSsAAFZB+EjP3vIO6iqZaurTn98mFMCn0icdaSyoHylBr7eiFgbiIZ28W2
k2lyFLpIykE0o+v+dYl+fypBFPM7c4+y0TonyvrWPQ5lbkYrkYMR9uZztUZbmh24
tATRHbD+u2hCBnuksLMEldzpdzyOVg/noPYRRMFuFtNzZQc75aprBTUPFebigWNS
86OuPbgVaqW5VhJibJkBpygSs3LIO64VatPfY+AQ5Qk=
`protect END_PROTECTED
