`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+iLDayAUvCw53joN74v2IRIhI2K2mGt3NpYJbzA1xExG9mGb+Xj7b3Oj6u6og3gA
7OtxkaUXsgnjdeX+Fe2d1rxRzYbX96RiBkx4fafruLHlgYIul5LSuxUnTkj+WJ9s
O4USJBD62m0XKHc2+0TZHNgwVq9BDT2qEZOI8S7/HqxziEbp2/wlSLMZae/mhiTf
zSVXsCDi7n9I4xMUHFrRpfOyQBjeLmicusMvSkz9mRgTvUr0JW4oBpp+sOOqRtN2
jd4ka1cJAaf+PaVg1qdh6ROvlto3LUaKEwksqVDxfc3ueL7JcKIuZyNVHfDR5klO
nDkmr6Scu0/4TQ578CVKqEQeCv84CzTfHiSqmMe9WnhY1yLc61wyN/warx+SLWyK
SX4vyv+bT/48E69czhvax3huxPUJtIUW3j7wedjEBlmHxlQ8RAukUqEZJYym5aCy
D9os2Hm1aJB7cbEMKXylTiyGNXbJdzSzl89pDXRif9wY0Ra8bAAoC73oS9WWalLA
IBeZPbzgI4z06jbz/TJqMjKBKxby9wBwOv/8jNSYYVrdcSF/QdjSkbIz9Own+pJa
WjcOp0IvOQGeBDVL/D7ITjTtqSN/QCdUxeoa0JXO+IyjN+nS7fNjDzsZOYfM4bks
tzY5US/wa5Y3USe9FJygCCA468lIhbbOvkVLoc7IoCuzYH5nD9EoYIvEgCHNOagn
1oFr2hPR0vPSEaNUP4/BGRBXQewKQh2RuVncW/4rhn9pk/EB4DNovdr91F087M8G
Y+q+QqGYba3zmNO3Jsb10P/Qyr0WlmFXEf8GZ5UGqbdwj/EhoRqUu6RjB2Ld/o8U
1bEkdt8i168hLWb286FB9Jl9zMQxphwyu+8FchoCZyS1wsLWeS7+lgTy2BPkuJHK
DDzKWNg31MSBlYHzPC9RVEMc05V3dU+2wFwr77+ZTgZThg1Pr3LhYUU3oiP/E4P8
0E543DgXjax7g+MgxVXo2ZPOCVcYEFYS2QKRW9TcditKInK+g7Ua5t+79EQDVnIu
gYsFUzT0f77tS8+EOezRTdq1Aeq0e3NqIT6dkCCp4Wb9X8VqCLDzQQZkBdjcVzv/
duUfrntoUMwcduav46kaqOIUCr+huPfpyKwS+RlCCgyaUnUfDK6wPmkXbp/62oep
xv/r5QWdS9gDS990b1jKKhsPmhE2P0JrIzm3OjqHVVN3fFxL76yBtaXng/ynKPNI
Jioaf5Oo998gFqKzyigEEv8fGTO/Yz4CN3dq/yaFnQ2026V1HTTWJEVFg6rQ6kRL
KLLWMwv974sF8rmMUjqBbriK8aZBDUuuLLymWo0BTPeXfK5mg1e11gROMeG5TjfU
Z1u0uGDYku7Uc66lVGIzJV3ziHmDHX1Hvfq8Nv9TNclCyafB/feCMlO1PmqRJ4Bs
QUoXaXG/Etd6OJ14pWzJh8zz6ayatn2wMjXVts7tQ+0zojh7D/Icp7OIjDQDqRTi
FJWFi6N/eq9viNfUZktWs6o5LN8yJyaNQEOnvoujBzu01o02OhyDXtBBAZ1adNYF
Xi7T6H+CSfF6dCjL0TkxKqRBCDuYOQwzsclBbTkoMIXyX0MaTUHRPbBnWDVlqDj/
qNWG9u0LEkWsfpMniWsg+MXf7hL2abFnPEkPm6ggWtTLMiZ7nsY1FiCaXGHRmPl7
5bDglTqPYL5AYOdOSqxS4IXTdPIHI100XiZa9bhSP3wyM4P54U2OgyofExNEQlWE
g27lzwTJR783osT4F1qKJ0SfXI5y29UPXp7MWM8wYJ4WDlYhcuHUz9BxguKvFKam
TIi5TUDU4LueSgpqWhArlYmdrOCh2ruEzXaOqXGrs+IkZZpqB6d8fr6pMSDZE59/
oAm0mzkLwzxWkHKmTTkN3PeoCH45Kc9RSF4bOVdnpsY4gGLicLAQlmOv5pPuEfi2
iCu7sxTnI+opb5LyzhKdPYpVPF3Tgq9CCX0JORH2903D2NX1Hsmye+p4klcRfgIK
EokNdJjFsRSctDVZDoAxZraxRWQsPrJsOIF16/egjdbnpC/C7JW3wXsFXWndP2WS
mlcISZ7Kjt1nDP/a0+BzDkkotxx607+/AxJDQyGfvNDLbKI1SbhT8zI7rVQ0I5CA
rrKmjYmlTY1XDzDnyaXjHJIf5S5lLQpGu4YePfQFjxloudoE7W7k49FzA3BenIQK
3vfeT67o3dxO5RxAG58v6GmN1Aiu1od2r/dhtNLklDUTa5Rnk/zwN5jgRVrS1D8l
luvaFFw/ZT1vHQdu8g726PWLlb/zRJOIIo19BdwaYAfvmHYjEbz5eoNEfEMDz8EE
jxKNL0qNGJVJhLadfv7dRGSfMA/Q7hUkK01Mo6oTp5WYdTjWqjFYUvO7rE8nT7kl
s/GuQ7HuQ66MbkZoROyc9fFz8xzKRdWHuDHVXG97IYF14YU4PosM701IX3CB52bM
PBthRTzxtGQ1tAMiEX8N8TYNJceFMty98FxWEjuXzTIjyjGGqEgNdXfnfDAWOuSy
o/f1dQxrxb5cBgQCRNDx5YDAC0OuXjamIiEj6dHetaoiJDgQK1JhMA8x6mqOumsf
6je8PYjZguUhTSadiZviIoE+zFLiIpx+WOHfvoa3af/5VOtVb4KwEjrwPo7NvXXA
B81TLixZdGdCJNncAI3c35VA5hmQfBxxrI3IXGrF5dWBSYon+nd5MKcx8lyLIfw5
3+XTdsUtbblaBXWDOgrFoDM7qRFm8Og1EnrFUjMtKj6idhQmPDxpmeGEBmKQzXul
8O1mp8EAuJIdJv+TYxt6XADY8L5KP4/jjXSnuw0feTaTh/IrB9zOOAlYlXsIuKqI
Ng/f6FPDvpHDSWyNumjpJJmQB/VrDEdq3hjx9qsHxjl4cBpEzGCyIJgATGyiTjbs
ZwU9SXStpWzSbHhaUqS2B2nDIzjNXYuk76bGYJ0/p/qS4Y7ac5EiBEbru3j8uLdB
E+lQh8d+oXiHrzaNZR486co3cb6iEdsqju1SARxshO7EG3MAtAkRoTgyU2FXmB8I
DY+apJ/MtTdSJgYWU5xLAVc73cDcTG7663cUcLgMdOUjOwCP3AjH/0CZfO2vRgaQ
79mvvGtvEb40CU9pu5S2g8xJQHewEVp8ziVUDjyaVgWW7k0ehkiso3PD5Z4BgP/X
oAr7JitqCyWZFqNCjfpd376I6lbmm64dyGKISgaA5CgiKpBHhZLwYaY5BfmhY1Wu
tdU6V5OM/FSxQw0b6W1EwWQFQFyouZvzeS7rzb5bO9mdj4f3+oIJz28P4sFR8S0/
85TJsxaQ8SFLZKJswuEur1bjxs8MJMYxxRZiIZCA3hIbSGAdsoI4LRYM8e2aLZW9
+MRsq4LP20at50ftRkFB5mNCGLnFP6/yedHlC3p8V86CpdFPI5nJERjJc6JP2Fv9
oTT5Fl6zo5wASZMSvMZb1a2t0F+3AE+yLWBpV0Gr2dxftDbzXCbPb1rlG1s4aY14
SaImij/LaaBNZPkMZFplKUHt6MFLlg5qT7sXKWRTKaAMq/sEdezWQZ+5fQACvLLx
BrDeaPPwPstPISylKKLSjXZvQ1suvlFLfYmcoZiQ+NlIxnuYExVHxgyfaNvcipNd
TByYK+tk1lenQGiC9XJWWXlka04YnxbQwcohkbKupNWL4BJkMrX9hGGwpb/EigLM
m1rpZDgVosb2an0uKGHFsVd9Y8pJTe0PkW/85KALVNTd5Soq51Qea+P44ksyTraw
q8nvSf1JSKMA8CsSen760fb84yrzA/+ElPof7SGItZvJ5Jy1jS2fOtyX6PPceP9K
HcTLya5tbGdyWccOKPjNekBSvkTo9Q2mnqgBhjbLyHZIezXQyEzbxOe/SW7cHXaZ
Gbc5ziI/ZpLxo7m+CtgM8A==
`protect END_PROTECTED
