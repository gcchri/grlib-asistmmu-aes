`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FXQ2h0FHRDcRWujhqa+EwXTJI2XIgUra+OMRX4eoS6CJXV1H/xun/GwibLcUqJos
2TM7yOp2zeM2coJ/ca4b2ip/zhYNHNiHFuMjs0z4aWAgHQWnUPuRyzwprAYh5gvy
HJ+qu7Nvg6jQrfBimu9c5neeqSpNfedE+vfT2V1rK1/iARSjY8C1rUYcX+VcN5wb
R5ZEweVp744CBgcR5QmtBdRkx9f0rQtFt1aczTKkNU92rcWIWhpe7nhCfhvQnFly
leN+jKy9kfEs5ogjteDU3IMLXXS8gjQ7fnEi+2G5GD018wcKC0pL+vk9oL5gZJnG
lrP7fCUrSulsarHqWoAoxHhs0e3oZv9v2fyBPImghWCFijqgkeX4W6Y1GGDTDp/0
pGGEIle4t0VswHjqeTDtwwANWekj4XR+YeigsYCNoYRmCZ93WFUkCJ2bcwRhZcWt
nj7bmMs6tf6yvwXjbRPOhUcogFKBsacDyhaOMNneq+KbylNkfiwI1qCtnHhHREtQ
XSy048dKa+sqGICOmvGvriX/bfOTPLI/ASXMyAtoaMn3tlvV/7eDYtTT5BjEOS48
RzikTDWkvFziUPKu4loiUkBxEgqwOeKklZ9IWKjuPwrEa8M2UxE1qKfNYHrhRwqA
8QKlngz/guLmdLKQ8Vu8xj0xrXYs9JtAXRysC+i2NidLDjPZq2MLetM04QdY5ppv
dCe+0cqcWI+Ocd9MeG68zyOYD6XRcMkON/Ci8SVtP+7A0EdgOmjqxIq6gaagMMFT
`protect END_PROTECTED
