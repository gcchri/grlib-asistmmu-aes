`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRLRfwzj/pEKHEd2x+xni8cuiSrPH9u8GzxYs9Arleezy19PsVgp8aFZRypBjuQ0
2WcWpFvnJ524bpAvJptYvRCgXpLTaikvv/2hxwklRdBO51WB/U9yRiTshXVdLIlf
GC9a+sxJtkbdf7v/UL6zKaZ2HNkAzLrQ0gdvZYqaZXxad0xt/HrSkYB8ooyu8YsH
LEgO2TBed/SIM4uWvOWhUPCqC4rs661RVHkzcqP2Ff9D9Eb1n+Jv6Ec48R59IcCt
8tEzU2EX/swoU557nXfNiqLuizkyo4QI2EDDPNoLaFSkyUbBEQKNppVlxjgIzbnQ
gKLAYW+wC7L0Rt+Fny87jYFhUhIBf1k242k7WyMeEEln03kasRoMxDY4H7vo2PID
3KJS7RTuuKQa0HJOfSoBx0V21kq/mO75FQJYLkwtZLcQ1c5sKNV2cttTzVIoSAkU
CGAFAbl4LmF3TBTsVayggu9a2YcO7g+lTY7FDdpXi3llkMzJWA+IGlPJluDIzu3s
0YRH8QjiaXQAChK40QV0w5ol1vib/e7yUBjKIIivFS8mXs5noNkW6AwXXve5RfzO
jQR9bW4srtWZC/IM0qZv/Z4bF46ntlgdQjRKcNjhGokpMhgwxLPicjjHl3L7OytM
b5Ts7HRqPWDnsPCpeaq2HdjEvJElODCwmYyOpoLr5J2Piqkk1z7eeCl7ZxruWfw2
RAVyZrD8GH/ZDcRnar7sh2CZ5vjjOxyJIr/P8U1vCaoS2e9HoFxxNisyrnCTVzwN
SMsJ4ubFytAmQZVZ5+Eh0DRLQkEVM8WXGb/fc552YP7YyvfehN3H/ZSZHjBFmxDb
r7qanG/iM6Z97IMGn16FqCDFmIffBHSSbWoTkxWfYLF5S6lHfHSyrLAyvC/BD8Ig
h/toj4HeA0My4MlsYtQNr0eQnIRkOfTlycUkWWH0ToZBPLhIsKSYMUFC+LfTLa2F
CpQADaqh2lDWhPObUvuyZk/q+7lSwuoPltYGxYl2hKqR+018akr/bVGGBBiip3lV
BDL2TsmHTadhcvXKNNnadleg9C6XdDvD9pxIbNCCHCRcyNrJhlTmaMiFbnpdsIvx
Xs+5yuuAVsW4GSAz608Eq/q3B+ejFXYWYoUPzCUkgG1F+9At8UPCenti5lBPVY6R
/K9uY5kjfXUGtFaVGSOVYgRRIj9uSkUkGMjLYd/x03dCW2FM0VdhFjLO3HjS4y4Y
GHV+W33nLYQmWhr3MvznDa825cTSJK3X1Us/KkLWoJSNUrOansfEIpVnmVtDJstM
6womd2CiQhKe7f8Y3i21KwmmU5exSq1ViEBo7ugQQModaut7LEAggKYCYHwJpxGY
FN8cvrYhmLGDVvVPoBs3aecSzb+5t2EjiPgv/mW/RPM0hIB4ffRuIbUxS1d0iBB0
gisaTXrYErhNWq1OWYFrsveyLjOINcUfDspK8glxoTt/vilKigBltfUo8pIZVpUt
BXQMs6dRL0tWaKue81qQXH+kfxIWCZqVp+yJgDMFKm2pKrp7M6kCz5BqiA2GD26A
d0L7OfSLWZbaAuw46Vl2XYHTCBPjFyqcv3KvMuaHVf5cW7xHxhwdKaGts5cUppU0
iZXwph1I9+89wIUQGopEp4mc5KTLZFZywGoRt+hZoC4uuUkGnhs6hEMnTP5OeoHi
mQheZ8GIKty48nMqmCYLTSNKgLw4EIs4Zx9V5hPSrig8HmZtfWelJ8KLXT35v6cB
AUiEd4annUSydXg9wEzPgA==
`protect END_PROTECTED
