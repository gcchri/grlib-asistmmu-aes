`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3x42sJxVLQhrGDHwuP14Piex1wBrK9FwKk58gzkTjjKxK+i/SvG6349sIHonO5fT
RfAOu9XN01h7Tu7ntoyOudSGgI+iHQmRAdmHtdGjoXLbOp+umwvSNZCHwdeEFlwh
/wmFoVFe4OTMazwE0pfwb8NBBn1VxFVoeVQ5gNrRNPZQDQxqw/1BioLYBRQj0sed
Y6cdYjwJow0Dv7oTz3GqnFkz6UVW/NRakIZ8tDdav7uPn2iB0nr/vdmAFemmTjD6
H5gWhlEIXGvzHNwYYG58265ZWlKAum3bgO5r/YPK5WCZjBbGsHnVVUA4G7fiY5DU
Dr2hvhKBQnF01af/1WVQBEn5ByK7a5GpLCe7nyas7tKO9pbDwMw2XOULQz4AuVXV
o13MCldkjmDNNY1w7VIJXVZewkVLqrZYOytxWY2RLBXA2xO9oRRAMI6hEljNSd49
4XDSNInror3dwVcxh7CDowrjxlE38yax4wQVoWYcL0Rg92ZGAcG7GuyZ9y8au6ju
`protect END_PROTECTED
