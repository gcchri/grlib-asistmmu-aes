`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sneQqNXjbnv/fsweOwamqFYWkhK9kk5TrN438QLQwMu5fH96KZkvqnrfw62ivt9u
WCO6wblyHL6jsBz2AIFNjaRbvfNiXjVyRx8aYaBUbs67DRDSBxY2Pyhlx1HVDJPM
ohGkN9TlHquO7H3EaAEqjw4j0MCUBBeIZt5bUKT3XrwBDnmpau0wIwCDWnc9SaoK
tTsDkiD6MYWwgO9wiBbCpykDPOMAfOw9yl6xQtpIduSL6nRsKtbcgGji+8PHntSu
EnOC2Of++Bv0C4+cU7I+IJM1Kcc9dP3jofGCdi8oVGKP68zKCERlZByt7r9QTJ2e
`protect END_PROTECTED
