`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HGI1UcfKfJmJO0bdvtot4/5ofIKm9727+nEORMx3GbzYbvB3vch93cQ+S5gw/PsZ
bIRsuFoFi4wIqghU8gycfn0xrn6ooHqM1WlL4HFOzuqDQiJEluUpceIjxPjRYDK0
XZyOt391AojTHScXlxJhbbtee6iuxVibhadB6TtU64VYDjiOnQR943WgZfvOxMFN
SjlMtfMbE1cyLKjmlm1eS+Xn8fkx81hzo1l0+iKHuIpmT9fDugoS2FMjlmiSMopU
yFMxrqlisowgK0NA7l1OxtEvSbYSG86zcSr7mB5WpAAfC3F2iLO0oALp8kujPfgC
MBoPAk7SwSsYHUgVmceAvubikXz7uAq8WQ5CGGBFKz+IIis09b8U6gaubllyNC9j
024JrJLsKyX/MwJNupPGa1VI2b7WCns7nJuPabRIgaGOWYyhA7Em1io75Q1k06Us
8ZxdZpMXjEuesm7yMcO64gAJlWdUnzlwap97/EjTb7/eUSn0FPRc5VC+Qw1UpE/Z
xZYpPAjjf+xH6kg9mUVlHMil8P5btcGYTeER+keMbwZ4WvKWlNmkEZeK1N+XVTKW
U8DBZ8yzzZvmL3LbLImkB+WgByRmb+iNOLKMEIxWD7yhy9juAQKwW/X0qUE11RYz
1W5oMmfW+bC/Z13dgXl3oEsy/UvU9GhLrzkcErJhbhBaHRTe+0nZ98HP0ckzGJlq
`protect END_PROTECTED
