`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
di0+UeXVRhCXu+i4rmnaV1EHdIcip9TLoUf9AFpyhFNsA9mFnoxiyoSGs0j1RaRH
X8JpOk5X8HiysVPdKXUrL+XTw8PtnLUAL6XTZMsd4GCCG5BY8uND8oCuNCDVWuSU
pguwkov+05LfYn2XbyQpi81nwz5DHd9yhrRh/dDjppfjrrXOxyTppkfhRuA5SLBp
5UOC68VmlSkLryQ8JKfXFwsnSe+zz7e69SmX3sj874JRAZX9CHXfdb5z1n8VaK5i
5fZutDWgebzy0Z5uNzz1HPDGQ3d8Lvf9JeW1v5CjFChxMfZkBWMV1uNfg1Bz4GKa
xmYznOGPgwUU8L1+SatPc58Ih0pEq1uaD19d5Niyw2TCUo8oFSQ4yXjzoZQjdTx9
8703OMHQVulWfkK8qByHZHB21NhzTyhccXqpQRa4sM2wC4ZJOe8Q3bPG1wEZB5Cy
rgMSKq/NcJMX+jD5TnqeV0NV/Dbjg8hIIkNADwSmtyc=
`protect END_PROTECTED
