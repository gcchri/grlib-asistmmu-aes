`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hsBn3g1fGMuh2adp97qwGx+00sYMHQC9771V8swzgLXo3b/vPsK4zJD44qm/sIU6
vpxJoxPakMOWYjl407++DsaZx6juV81RbP8ACUI0C/9l/x/1zT3/IzAeVazM+aa5
xGhyWLisyqafgaM15iCqi6FsU5pGylEh7w1JQdbYqJkMwbfAGUva1bbELaeMOB/d
NUVt1+hqpLjhmiiWRIx/fT15NjuQZPWLFcCriXFQzkZuGUvhcAfOatsHTRhvxzzQ
mZeh75Me/QnPUlWKGL1KZRRJQhB3iOXKUg/K0Aq0LotYtg6/Lz90SvLUkv5lmaPX
aAlfycpdtYNcUUwMD7OvAMF96Lkn6kG5r4tGqinJXMHLXOfGEfqZIdNqt6607KLN
xMzP7FKCMCtfPmoW+ODfcmGgeTM+4+8A/5sDV60ap6dVPjdxuFDN8jsPxVmlLC38
PzIHo3ts8enFiJwTt8uwJtHsoFI3S499mPFKTpUJkim34gvUsSJ0wPrZ44hYohUa
xcaaad7iua4DxLVLs3znIxYopBsi47QYDJmUg+3oRilbKePavvA0CNT+sGACNQNS
Av+bkqEYd0UO/PvKtwGJ02ejN7XezCkawgaCpPcJZB53RTpTf3tnuBVb4H3klCq5
7c9NsvmTbdLn1T6pmO0vy0+C4kzK5zawFktXIByiwpKrZj+HIoXcmtUdRNIkRQNH
/DuMOKxyfhWHg2HUtbkUUfTNhOGszFId2Xm8T7F0L3b9BYmnV/aQmVYn2MCsNwj6
zjtwEJDx4xzxoyY4VBoMcSyK/8U5TjXEsW2a2HKVZQ/6AZnUKMxQr5+RI3tLCFCI
ee/JICk3n2ZT6ixIyZ1OFUEe+PQi08wyNOV7D6kE3vyAe1E3C4aWl4zxCz6d4CuH
7Trv0m0kBxcWwpO8uG+RMIuM/xIM+KLiZWvVBSiPKmZx4wjwrzHHjpoFvwXEtUwr
IrdXvqr20iEKPMnrnBlScWNF+aXTl0VTLy5gGlBxgkUMTd26sM1QPXYyDnJcdTKy
/szk4QLLrw/zJeiuUOtjXKO5bFB34tq9td4f57maJpe8V3cuVmh9jwBYwG00Yhb6
5beFUjmOEu3SmlRfh4bagQljPfbEvbqhQuoGtwudeOsVz16PSaIeDGWfV27/hPS5
nANb/4xYiYCBN+FF+ztzJaCogGn8ckcCNXIKHmxCUckza+8ez9cECwIGLYTYWp+a
J3jf5WPRLuWg2GK3lZavxvHUXp3YInpvL8AFUF9saA/e7KXErohzL30rMQSv1hzz
u689d6t5dYwTllGOqtt14u7GuVGw3TBXy/E+WR6U2wsvtkrs5LC0UyQfTRC6olU9
rjN+rM8tEcbyYGehAwrPTJCxg2J9hRH2jyS3S/hI32rL7fo/UbVE54lmFXuuWKDq
xcK3v1VbC5bVNQAH3CNvtjxoKOxU5afbrZhfG/jVEENXrNhgF5S03006ILz6mDcy
xHi7uU3qfNHpLzApI3AaE/DO17kRRMCMGmXqJgRZcAwuf41KvVkQLMQSHFz+Vudi
zzHf7Iq7uHHTHiri1hPnb1Xt9ykyfRS/WuYtBA3v2JJwmqeMFPHX0TFGSyh0b5HB
zHKj3C3McQJ2vXLJisGgFu41yc8v7M4ztHrX87Q9tgKv9pB3opYJ5ylxH/as6mGb
LCT7rkJP4hUIZ7ap45cQH5DB5pOzyoDif9hYaGBMpn/ggr9/TtTAbI8B9wfdhEJ+
yohZuwDsHcrcRE73C9lACS5egNXc6b6N2uosYOgY0KV+eu8kErHK0XRZB3xnOnMS
zNTCP90Rs3sTX0hZ6cY/Ay+6kueDlckkHqBnmeCiCJ/0IE6HwTGG2lXy+IdMMPWC
PDnVY1Ts0I2/rHalnB4J/tYeMZkAciP2zRFOVFyMx0zSzQvlXfz3mTq1SkcYFaP2
dzGSFrPdTXvjlrf6oFfQcGYNsO+8luwqJ6F1O3Nq29lMcDbO0XxAHe/B0MNe3XiG
mycOkJXbn5z9gZQm0SeN5JQDUWmyTz7pjIXmB+waYBW8EJKeFgv0aq3FRzfew/2V
JgfFE8KuIDn2GP7YAWw1ciyHPB7Qjb4k4sc2bBnow3oTuUanKzkdhcioZQO4SkwZ
UcXHVnPu1F/qbhxsBYOxL4b9yMIzzm3PF2+WFs200Uv3vC5BRizty5NvaGNkVpX1
5Kj373eHdfwHJMeztPvq6KuCefRy8mFESnq8yPtnvKnVWUL3JMRSLyno2eVzOIxJ
7VAh3XAXBK2oraguXontSjG7Z2nDd7dOav7EZl1u8Nw1m/fe4FqDbUinHfPmRxP3
wfYFOs7eIxOPBygZBgNuVs9jilz1K7ixNWbR4cu22CaqDKprZ1t1RT/BJoyfwbyQ
qZL/OmlDGKP26OwY0bWecJlklW001d7Jx+M8rvLJScHIs0XTxb70zPwIjpDtgHQB
+G3v4Pu+MqqhOUk4TjAI1eqXMbyyW1DxEPvo3xMsXgIL2NH0vPMxSjePpHsbErDh
T6JvEuAI7Im2ti8bMlDYRm8Vad41nBYC1ag+BQVNT7Qb+zk5uZJWvAhYgFMVC7/y
PzWjt7Fd6rbPuQE2nA6c0M0WhIg3zO2R7zGXqdGESzMZeW7Cbprm/GN1mdllPAsq
Pl32Xz2xgnKIQlrgvhtpfzgptIifPbwRW0R1vw8AB4cTxIZdQAdPzR/8FYySoqzR
CgP0E34RkxJ0V2l8Rv5t2JZcxLvyMDWl8bpKyRDwQTI/+WCHwLrm6cwry1Wr1E0T
P1GL6Q6uQqy3Mv3Gacr9rhdiDzuS2GpFaOEU95fiHRfsJ+Mmpmj+s4ZRthE5eput
FLsG0MDlcYpcf26favUqz6U+QzN5eqtaMJ/rOqK+5io9LM7+/13GW8Jt6J2DXust
/Z47xEajpklJH3zuexWzoea1sWL8WUiHh/o0WDfpzVEXUXBqYrjzf+FmfqfHWCiP
pZYP6OyiFsDEs4+acNjxyp2zq14e44zf1xmCclG7J8Dg/RaA9CDUx0XK/Bv7DXeh
K0rZTUG4GST+pRe5A6uY6EuHb8fTb1pzKLHkfDP6s2PANuHYYcgg/HZlErsr6c4V
0uxd8CCcnGFu55kBXNwuc16ZLcnOsapMe178j+9PTB66e0OHZFvo8M+++8OXZL+x
+5ROU/oqlOz/SHh4NQRSpOBu4UaksFGFbr9rTOlkJoGK0hDG1vTaU9/ud50oMHh5
DT9tzFeBtbmT7ZVL/nWroXfuT1jlWsWtsLflkLWcyyZK/3pbK7pYi2kykXHKFbSZ
YYiSBReyNjRLvPvc4fqeYNQme6QNLKk0T3HwmvO942wIZk15ORoSEu99DgaBV17b
YxsCTl3EOWKJd2sqmqobpqKu2xAwXmmfDwzDbrICQTHzY0cc4A9W1g/lE0YIF5dX
UYWw3deBfCdClyJeEo/YucRsRralVTLBzLOheSY5LZ3gqMBNZznZKemTwkcQwOq7
RmusJ8shMqkbq3pgGfDJ4KWIJZy8x6cLARxuFztHM4nVamxr4W3d9AG6NYVhNMQb
LJhVcXLT25RawFXWY+HK5n+ibzqa20Vb4ZBmDVfihLNtXFvDGAk6NgHNrwqjBQXP
7heCn7sQ0HHe5KaeU0a2teCmAwL6rwmXlpgN3KL5hQy1EhWfwWdrDQHS96603uOp
pOPy/wvVDkxI7ZEmke+INIencserKgcyJF9x1sDbbctCjHfBRTYPy+eQ8o8Bm2M4
gzWTL4RNl54Jiba/6B+dZkRd92f09HG2zvsuEIhZR7hPWswnagVFqePpOhZAbsDZ
u3A20CFgEL6llZSninutaCuWzLDODv3/0ReDTLph1Wl2DZ3cs54FWHPNptWld2b4
t5l/7zK+2VzwzlO1f1Ope85vCUrLynB8iNQtjD0yE+jQa/qIBYQPaydNETSxcmId
+rjCuPQCnWpsv65/kftUcfUkAyFXl2HU8fgD9RU7Mtp2oOsEl2sV25qRDiON5Oy5
2yX3xfg3jiU94FKMGLKWwaHn70TtgAEongrXeDrXyTHUInzXlq/TQlL8GKHXvZQh
ks/ioXuMSwrvwpfY5KJy9d9tjLog+CbsVTWXSvb1d4pv5FpAFMjIpsM9oQ1fJfL2
g2WmN2uz0RplT+qvWvAQ7Z/ycs1n/w5v4HbDFe7htgPMPzc9mSMfZu0mIrCaTICS
rg3S08N41OjXgyVMl4zActEWu/uu6BW/YXJkmY0cwkju0jJWoU3nuP0Oj8hXXfnc
8oNpmTHchqujRoz1fOfxz91PdCZsMf8I6IZNGUe8NdC70glyfvRKSqnWfT1GwXVt
FLQQkugyHCULxV50HAb5I+S+7vV+sMOPTXcotN3K2e9bpLNtvjdX8gouh5XDwThh
N5HoLH/X1JBsAGSpz+0jBH+flmgk/xFceJm4AezaG51ln2y3rAdoJugzefGMkSOR
00FC//ar5B4aRURNCcDHkX4pm4Ckf9PoQvQ1FZrvuwzAN/1cson58G+b073EK9ou
3bJIn3E1TotIk/pGMtZfabyKfNsv+CfKm39CsUKDD+2s0wroT6hJ59G4hdrz5Wwh
VFI+9NQX6q9cO3fxDO5Joztgv+mU+HZcagc+uk0CxbALbXIPsLc4yiF8i0uMejTt
edPJ03Zb1fiqCxI+4SYu8ZieRwBZqKUiS6sN6Be0RWxBx+T/FtElUFN8KH2l/ox/
et4boLRZHAKRplN49QBZDlC6EShZij5r8oX4LTDJ0mOaKBkZC4pnzNBXT99l9S+d
jikfgiwo6N+/5uqLhIRvYchhCtkew4dWJg+GyxQMWwuvl7dCICRq0e6oyVF7Uetz
Mz5Kl+Us/DuDMXGUKTZuXSIWYoTVA96NT3fWaOxmW49chZOSnDZIAHIzwX3QJLG1
UZJKEEWsUWx79qs9pCPhhUTngt8QjFJVdQ524AD0ZDf9A5dDpi7cpq8MknyPByIx
yd9vg2eSab+Z/JSiX9VZtcanfzpRiTcJNkKVHyxd5myyJnTeU2y22/bCVywSJPuj
eeje2ena5HgwMGi/KDgkZKUSN5l/t/kc5J3aXsM5z4X00S8rfHzluHcegdGvD3u4
KmZwSPwTANus4GdIF+J36phQWMrCDTs3mfcEvIr9P0jsPmvNu65zGeRbA/XUpf8I
iwYl6cL2CMPpnr8uA2XSgJaBPlFkqJByMYjdzdZFV8sFGEJBEhtMeKBX9CK22wLS
Vz59Wb+PJhQYfdvBdN+hztZcZXzZtX+JbRERMiv4xdBgofS0WbBa4zkLtDQQqlCM
lYfXXqybdMCCSK1ZeNgFE9WF8DH5UkC9GjJ1EmRXxpSiaxfa/4J+9FKqmgnEWWE7
Iv8IQyPZ8+FWpUU3bWix+MaCZ3ea2h8JhRP8KMSB1zFVlgnfz5DGk2H2myiEmswi
rCVlUE6soNv4lH6Wk0c+2RC0xFPWzvQVE19VG+iT3oJyNYn4/nGBrd1WnOAvceD/
CxrZrgFv6iRRjyOOih118RCOtMcajhf2BlxiG+5XJ15sERxVkNitIk93RIfDP6Wx
OEL/5cnLuRQeP51whefCJlk94Se5HsDCzQMzUltc+/OkTVBueMYGzSqIOwPcciwe
ivzR5JCsGAeAwATHjTmCT4yNrhoWeD02S1Egwsne8S7HyBXmcRJmDwkNNq2ZX/1Q
e8E+dWbE2e/5cUcK8Wit9uCg0zZaposX5Xuto+ALU436zLNomET0egWjPOKMLPvl
BrnKm5YQtCitGeYn5uMewq6U1L2J3Q+nA6AsbwmPbMi9E5HB/6cTm6MRP4/dAA0c
rwLd5GpofPdQKk+zC1f/RIeJhqLcemVdvfcIKRCQG0hFCPwvSZurkMePvG2WzU2W
MjRRzD0G3r2WlpU8nYfBEKsfTm3dNWBkybDXFnswm5Ww+nvQIiP7r+XKyrEY+qFu
wW2/9+KB0X0Q0X4S3urIUWCnaUDfYJBKqEwiaiKP5oEB6NkfJOfMoKkR9sc1tRPq
TDUBdWSUtinX1tW7s8oEmg9VhyALWpNZyQKXIZYdRi2N1l12VBHjUJiAhodnjjbA
ZrD9OakwL4VZtONoGnooWzoJRuY6IpNl1f9DHtQwE87I+Ppf6H6fI5BPUf/EgdYO
ufLx2XOlaidGecYKzCKuzhLcrdO/gH5sSUpjrSvgGfdtHLQAQWbkcFioOI1xgbGZ
TQ/MLmu0BAPuqyUXDqmqPtAYjvAPzXU1iPxKQQS3WmXME8MEVOP3G3VEhR8dJyHO
okpQXhl10dDWC8JfFOf+O1iReJgBqQ7nBgf7vTOAW+Dhx4FhZaDwj+4ABmKn2y0c
aQrNbOIpH0odv8MSjHeO7mSJbcg54G6Xgku98eoRRV/MLNI9T2FjNlCGe234mHeR
/gI2Bbk8JVnJJ4vabe7ei/xpHsa2I5CP+dEd1h69O1aLTxga6JLh0oBTGEBlr3PI
dIxsoOSDuUJ3rDzxMTkZIIKfBcl/eO84dBkohkk9EbKo5ccD0AL7+vptF5k+EOYK
euhCyTo1dmYU/GRYjfvtYH5om2lC2pQ2WKKibC+IAMV0fugDE/6rWoXI0H/71GbT
g8UP89zF6wYDq9aRNBcjBIbmtRLrIE6T1Jn7jmiy/b2WuBms90zNwpP/zTw+Vc/j
g1irZJSzaMan18at9mWJH4xQ/RrbYG8hR/kMRox6pS7KkkrU0p5nQli/wILYaydk
Mp4lCJkG2dn7vhChp+Z2Lxcq0Uk+q2uvye0/aNnMFYCP2LyWezftPxtp9gOsRzcW
NPvWAYApDg/hh4nn670VyD2lsBEiQHXecSwcjyu3+SBtYDNKJRioiyNmyHv6KgYF
h79hdeDq8CL+05Bkwbb8xBaTL7wT9AogbOlwLIBOJ0vrXeQ9Q3e6gnjF18sobuvf
z2jExYzRZKuv24nNzWB/N0uyEu0nwQqP7kRikLAwzhjDlL7Fvj/s6jrD5BoSSTY5
DOKAFiB0zHMvokApeHga37Q7CqWdM4qJQ2tR6NfB6yA6BQsBiTj2llGOp/8dZ7F4
/LtPww9xCV6fMIMgcdcbPh6VJkkWpLJLeoDJzzCRIQO1FO8tbz3Ketgtb23utYeK
BtRb3EJMmWytLj8I1MBFffd5S+ZUT3Hp0ZiX8rL4Q9PD8v+vSvFUnv7KmDhTMrPS
TVV1qHq1MkRHRYa2ZAn9ubsN1930EWW5fyam3QuXqaZXtLB/b/cl12kbnE6nXpI0
Hx3ygG5bjpJhMifse+Qc8f0yV9GcsJhoo/64hKCvvWjoPIwChHgoWLY3NWmNXWsK
wdkygijn2srvw0cZ+N1eXIWzVaheQkVhXhCPKafzd0QyZAfUZKMhbIilLoqqSbn9
ui2vzWZcdFy+BlKTJ1dFTDgQTcecFA8XWAAha7tGDcJzykip4Yx66yszo7CZti8a
E2wZKRiCEMpHzao/6VYw3/A3fEo7Rjbre91Ea2/NedPBVdGT+QbCkMxAKKonHefB
WCclSe+ZFi2Z3gOmgvtYiguhM0Bkj8L9kBfqKeAP56onfBxzGEnQ3BHHd/6tVB9x
qUlfsmlfH/IrjW8Y/ZbYpqSBlt3H9pNIOxDPnzqmF39zJx88lO5gXnDKxr/WNMZr
wvMB4DaoNXCVyOKbXpvSOrWIYTPVmAhbatI31i+r/X2NhTTE1O8PCvn3SuqQADw2
dnub8DuoGcftFKtIhx3w8fIA9xJgWbSddoTm2VawfmG529evyW/PDun3T4F4s9Bk
QmNneNveHWp9eZhxapI7BIDb+gHEuerQmRfVAsY+E3gP5GZnGZEx/WYq1w6PCnrI
ymrSIvjVFVXbLExXVePTldc0MgOAwwY2pf/8qzChJWIMy2x4BVu/9TVuQJSf/TF7
+FROLRazId8sQVwDIxTyce8CVPBtId0EfZzPRVnGjZIzkQLIglgbg8SehU7Xx+dv
GmL8asfMFTZtXlkYW7cnvjWYB78yqedVSGYkF7FqC8CNm3ZGD4V6+dSuvR1UbXo/
ETgRHJFj0Z2hK7/BET8TTBVx2BMDWhHRhvOckKKdQqk39W4bYnUJPHgNg5+fatY+
8T9oRUG5fMqjG0vMQwiOSVSBcgrmr4UHB1oSOmkGBbrxzPIUA+Vj42Qh+Kj3c4ku
Ms112DllQk4L+OjekP2ZES7QZXQiLtYQ3ysLBBJ8RmFPrqwS/Pvz4X8tvMzYHdn4
yKdPYuFZV3E8obBxacUhcc8VJytmVTMVJp5ePRWAVE4I+GaJQ/SRM9Oj6/f8nAXY
juWuEwH0oZ2avylm4Ce4sqI19tJECD9mVhlzD6ttJK6RuI24WWVOZ04mT3hwg6TV
z4BQMMOWJfQ8tJkAGQ5u3DUcewNSAolMIAVr+5P9vj5MwnatVr+n/QhKTZdKMXqT
JgAcciTCh9DCLR221Mr5aZKs0QAIKEEZ+DdW/kzD6iW0vJrURIWcoG29MnORu5YN
1FqIircSsdFlPQqSOBu0+qKJ0D84+vVkI5PJnmAR2dmDBYW/QQo7FwoGOMjL5lJ7
wYhmkgV3C3qggj4y5+fyp/zYj3uQtQXj7u7YVWi4v2tbKkQy+uqXynINMIRW24qI
Gt8NeGMQmXcLT4Snqk5dz5t/Fgmge0v8dErEPvv18NqGbeTSKblAqGOezCBtFl+y
dOXAN971qt65xx8XD+iB8GD/UCSnuaCa/erxiKi2F8ii16LbM+E8SZDZcQ7MkyGX
ziyIPjjbJwyIfwI3uHIwNkgAHZA/a67tXpcVrLENPWgrzdxNTGzPaOrtsG99QLgT
m9wMLBUkYlkfzYuX+BYzK4XHVVBsymw4uI+lHEDUwWiqcSqwdP3Q6Hck1hAX2IHP
QtazcEJERh9ubooH/bruC9qCbcvDbujGJEHR258pwfH8aj6INwjvlbsK2bk4sJcU
oTxdDiZylzKapWYi5oQjQtNcyThVQjm/l4McO863G6pSCkkdouPgHpQ/nsMOyFPx
xWvsJMk5ISTOHmx56YhKCtVEd+sgPIhbESB92o0+qKKM1rSIT+sT2BFgvT5BqWiL
PNHq5kjBzLxiZdBTPv80nP6o2dqP8VblGbQjVUVSYqurwgaLCen4GVarlLqZa5Pp
MMpaP0poubp7X5FhrTFkhGJ4iwNsxSoroOF8X6D2FSc2ZWY8UodXkJpW/QujR1OA
eD0iCyTm0ln9Q5uszHYDHmp7VIEkbMzn/TgsDMcc7oNzXLfVOxQ+bUD4iWFiimMu
VkSJkOxum43YVJOFZh3tp8kdQ39tk5dvV/6/JDln97tunq0abPg1ykY+rSu2do6c
gpANxb1IpprZmjoBnuhuarRcgoxmO4g6qUs4/Ve99tFkZ1IPBUf6hhzidvMPuh87
GhPD0r1s44mbG0wwg1dImvTTRoPIZO7cuHV/RvnSlnNPhN2iJT4vnLEiNYY+8IMZ
QuwO+KzEiWiLDjVCt+DoMPQy7kkWj8NUU9auFzlCIlJBejH8Y1J45MnQof/vxBQ3
SwefjCOK++7XIQ5gUv5NA3OiAk31kSdI75axvdNN7A/KpxkZ7D7Zo1LRLbimLUDp
lnunb00ae5fXAz7Hjp2jCK7v7QuL5Y8D2jMSiyQy4eIQvLLFrtePxapikvWSIagl
7wOSnTwUFKgvZBbC4hoAYd3Ln8NprO+d0H8svlxOy9oeH9svB3Ngf1TP7OAAodJb
fz01qYof97yowiTQgnx1Ffc6UftfKRBl5Pt5pTBicDMFFfwYYGwXRvFqkbXP4m0f
LKZJLOgWB516uNbrKYxbRVJFBxWnDeVvYiGGqhxWoUDwdFXCj/klutlG/MU1WDQs
U3ptiJta2y2UX61Ojqnov7LIYFi9aPJ+cl0YCu6MiObYieAVZgEycbb/4YX/fI9z
RNYbnfwhml3CpEBM8vCZSfeOhxcQx9ZOx+NYtWpQ0dmJkmxrwdSWRcz8QhkuVs/H
FxzjqGr85gd9+3H8fouiPBAjk0t17TUl7+1unTjeVhppPdxBO6xMwpnZ6Do1zs2i
ZRCTczuDMcb5XPHWUWayO3USK4QX4/Q1KNa2wrzIgUJpxyk24PmDyhuqfR/R65wx
AYiExzkZBKZJZVrYZeqIkBT0o1F+KI+X/qeMl563bi2Oqst80+qA4rejn6mg0gVr
H0hr+X5ihB92lvB7WlsRDdDphCmaUQsPFtwJhfg9eAZ0a+a5xqcq9wAy21ChOPsN
kUcsimqNkYRyoS+0nh8ySP/ZK9osq/o1NH1kPwsL5RGgb6rKbqBDvJU5YYZFOw9p
KyAlteugCnm2390oz2dXXVBx0/ekpIWtM6VUjvhIyHBQeqfCqlEq+Z9jVNCpu1Tk
Tqks1Eh0Kcm1+ZxibEVYKiFjEMFc9/1CiF310ZBxbtEEnxBpBa117cU1SvEFuieA
9sfvIy+5F6PT8yhV/Gmx20wyCFW1W+UnR6k8z381xCGnPm5Ggx6/FCu0KEJ6XLPU
wD7VBG62xRwOnYTPg/rbW5ZW9Dh5M5HXelL64vvmgWDbR5YSN7XTDbrkwb3ididm
6aLs2pHQilkDtM47wOWou3pQPr5cXjZzgu7Xy6/2iSqfLMEnux7rItbhup8hqVul
HxT77RZigWHaa8cp0/U9HKPQ+1xL/YPuqdFnte+utmxR0kUo36MQVZYZIUszn2Ud
Tlz1jZyuEtjDU69iNdTZdiXBT4XAPXKBhifdsL2Xapp1im2r+Z6CckibMn7e2GzV
pa90BouK1gkZET6tv6PJDo+idOScz3CNosUxMylCdwWmSm1rJT3fIhE/CXEQQ13Z
hgITPoA0bJ3v4hwIq+/LUyH4voo37k4qWiOuymgReoPNFy+lHZUR8YmPRk12Dxru
64u76wcXoSBEruQhl4Xgq103dEJqn1QnV1AIh/eBS4lpySrsXyKn5RcLZGvfJhmN
re0gZQM/OUj6Xcjg+2zN2zbbT+CvSwSbyfY1wozpDM6Z44o8UReX178wlv5D+Lxs
HgTPzDv/WwQ4I0GeDIKW7q+q0xBEN/cIIdPLGuGH10GQ0K1m3kpwYG80+rbZ0D2O
kzFHvqrb7RKoxI+HEinKefgENl5w4Lk+NPONGxvuCBmbvpNDMTNDT50vNFzt4UCw
6eVxOyBrfI9AEj1X3+DR2nIpkk7V2Btdu95kZ1/gUpvxZW8zXtCSu7AjrG19wyb7
R2845yMQTlyvuiow63tni442x+Fl/7QXy/6o5Mez6RNtDYFpViFZaQcgLmpgOgeG
6ToCDKjgTJPg+L1L2R3FmOTY8hSVRK/zlyy/ld6PEqaPrFugBBxJDKGGImFk1xAm
2rcs5wpEuZEh9ZcMidHnnvY4/JZMi6/ZE4fssSr8QIYz486aa/hrrCKPhvlKk6Rb
tGVlayge3Xmy5ZPSmZD2fLu8uJHKHKUNO0zOWNMy92cIbJLQh/qMpiwjQky+I1yn
wkn7ZK8CPB+q8khCnXvj+LpBzHKQasgd+uepHY6wJ6vWzcDDjjeLLrVv7AcYqIAl
tvKXgQWEg3Y8Hzu3+l5tFqtuWGNAxd75mMbLDm/gnqIFpL8EJfRla7BEXuNcz0kO
f7Bi8UNY8p3tD/uBxuxAEx0dVArlKariAt4J8lMlkYEz3Lc0EuJ50JUERajVEe7Z
oXEGJG5FP/05ORyb+16N3xH93SwzDJmZ9TaCee7ZzdP5DeCHKevzYBRqeW6548pZ
vZm+ppe60pQG2ugCCNwQD7Md7oxvir4XFQOPqF5Ydz7xIWnD6tcSYVZycCA4tm9f
hpEP+zX9RsSst/4GB16SE+4/Gvv8AzTLD3kRSKIIuz7phESL40zLVAAkANnkiWQw
1h9hqRluUC97hKb3f4UtsntP2H7CVQU4oKF6owvAqdHS50L4zX1jEqIUXwnSsbHl
cuEUeJYgYopzD3q/6dgDi3dLi0HkniYPH8I+rfUQfhTid/eliCobqQg1vTlplZMw
o/zWcVf596gRZJy3YyHNF4Vsiz+RQ8b9tW4sj3N5ojgB+ny+VXqXWUZAHBMlqu68
gRvE+j2T80uY7vtvm8EHlnf20bk/aGl0uyQvmzwtz1TMS1ngyGnLIJJk4ApDxs7U
AA7JDRNC/OKczcLZT2PQ/UPlGp7JCsOHb9BPZvXWW00ZZqYKOFQwUafeT+N33+hb
jGns4v9XI9H1SXmSE7IYyi6adsg3fjndSrPnzePCga/rOqsmGXY/isWP1yG9k+OT
4K//UISEa7kjLNCcVRXmFyMZM6dfO0nCiogXsfSlbtcSv+7w7y4TjpDiepeo9Xzt
xmL7e8oZVN7yUemkh8EBhCEXx+79yD3UkK5HJtP9gH+vklqRJ2Sipcw7pnfjQz4J
05xrvzQj14X+Ubhz4NutoI4/TSJDOi0amdCr0xyMs40AHLDuD3wtVS0KkJtEbg6q
e4d+uN5gqpdtyj34O1TPpgwMtmDqFUcbhw6zTk9OdiNWPubczv2+PlNMGr2DIole
kfQS8SI7c0WCGturlZIRKBhQgFm5NdXxrHSAvOXJcIoSczV8T9j3SEWYed5YdS+G
1lt3bBEiTTsT9vCSZ2Kv1pw9PV6b5ms2U3JByeiyy3HYMx7m1fgug0yGMTJqmaZF
9yCmYFNFXh59VVnsMue+TOyzQxEGZiKDl+vik7xi3TmHCk8ZotlgPx4IXpPzSgzP
MpFgqrg9t/REBPAkTSwjSA4BdJ4qyKXkN957Sg7Poj8kNbYh17iJhyvVpFAp3q3v
P4nAAfSHksyzrZCK9A2TYPnWULqOQHEM5LPc/iYFkBteUznGLUlbobe1Z7m1d77x
i3qR9TTRYDlvQuv04ZWkJEE87SZEdVy0jUB0zzHW7jFtKBmlrAm1KEHQv0mOtxXL
7Qzfgppvmu5ZprNUmjRxP+f5j/0NWQpBRsHD05Rfv1S1fUxeZZLQGYhp2dH+xel+
g83Sb8YkcMFRXRg0OD6EU44cmbdy+wakVJrLyU8DYputukgnMs06Sks4x0jAQIVI
mQ0H4Ouqjjq7+I9mGP+cxUVAR2PyrwCDImGaHzir4vQ7wnnH8tPSffxzqXWZN+to
xtHy9R0NxBbINSiyonZzzly+XdT56kedDyRA6+Kuwkewi3vbeQpa3fZao6JmpLjg
lvJ07ZSaZ3+3Nk9gR2udOy0e2m88BHdHcWhq3i9MoLtUh355u3m5Fs3afBHWg45X
qH5dr6Suw47VxvX5fTl1k03TbJh4SpJN1/+7uFyI7tXaM+S6fWWTTYkmqv8yXTKx
fA+eRnjmxkhHu6d45mMtGPTpmR105xypru7EUHzx4dIsHXIcMq0sU1Sd/UIPtB9N
Au9JAEF/0YHPmkFgUx4zUN3bFm5UTkRrk8t4vQaeDEi87wv6HxGjrbu7fxCMFINh
F0Kf3tEcHvJtJQEGrkwgzRn/KrhDlk3g2gavgZXAVBZz8MJfmbEQ4dTLRlHOlD0+
EhTdf2o/FJod4mMeYvX0lqIt4imOvXjnr3bFYmVMXjlwr3pUOppm5wWANS01eECi
AxWIz02mlpPqf/Q0T9M+UBeaT1oO1pe2twipT1XFuS2JPbSA+vw/5H9C+27so4YL
srHwMP1J6yu5upIk8Vu6l7nnJZPanoTao3bftp4Ourcp6cET6OfF7IEhUKG1hfZs
nHtAOEr3JiyCI9lyEsUeTFrUsIbfhoHqpg/Dp1W19rv3A3UTZwaDnLgJUeZzd7GJ
n0vED84kZmWXWn1UnC4rQtauZmmiTF0DxHZxw3QMzz7J0SoCIxOyKWCeHTsrwM0b
XT4niensJ1thxfiz9jwJmP6KlICMiv12kv6GUAaYqiVhAz5O/iuTO7tFEzNeYD4P
+3WYd3XvMuQwsrnz5dP0pVx77RM2mO8YEsUnlGosjxBUWV5nRawqEfa11FF7M2un
nmxKi99u9sVKCbqAGANyd545mWQarEs9yVp2Bq2hDyHUIs4HIwhuk4Gbq45MhOJz
ucc5oiDrWpz552RMoM7hwW0YWUJCdFbATOt5aqc9T8+TVfFRtDQ1nFsfBF+Lc42r
p3cic7STLWCZ0qfeZfzhTJGIV8TEGaJa7pC8oL9K2JXhi4ZFmizk4RpM9cIL2q9h
myK3u8o8CsLozdJ77W2kuHDRw8XKXgDKd++WKfhEQJsTCkd6lthm9zo9+MPeLpfR
mRD1gTvvm8J2oKvbTM+Vpyp+nmKf8NgR1+vCNjzfF1I4uC3qjOrQhTKPmli6WiI1
9HC62UFIP8Ve1w2uBRRAAn+/Yh164mzc+aQ/iCNF4wTT6bjXBavadrYyazFBl4oa
5YTG/ohIWPq1rasipqwf9lT7mqq59UjoLpDomiFT2/gw+lGaGiZc/UEhcxG3eXSK
kvMMJSQvChRh6t1AxgHcxPenMQo1oMcvgRFt2MpnvbGu27Ba8Y08812+qdUzj3VV
4csDRsUlNC956oNy6M4/W2u2XR2/OQQSX9GG2CyenLhC4hGKhmVAtIwB3CjsZryS
dG/haJA2vciExLkwbVGCtRE0JyJPzrnNmMNuYbw9+FBe5xZvhhyMrQFXMHhlOZHy
bq6U89GJQW+tR12zsDM1LubnFYNjslx4IMNabD77g9XzwUqJjNvOobmbps1zz97D
85cw/gSVNDwaFVJw8IYvqbfTiVAgpcMuaYHnZh3gqinRThnmMWRrxRk6m8gMrshD
aIVI0b4h2bc9taIoD/4GvBgXeWU11ZsGs/NrdcMO2RzvC8vv+xOal8H48wI14VO5
RCye/erhGmZpBJYTf5KpHQB89t/lc2O57Qumky3ZR3jh0RKpzI8N/HvCZvePaZtF
QfFJPitSetIMVEjh9f+V8tTSh//daokmjf2a3+Creo0wMeOpqTNwMAjp6IEUCX6S
xSjngCcl/XjHA6Rrpsege+S6VeNB/BxFMeahGRaz6OT9J9a391juS7RFX4i3H5hx
nyKQASqRql9iZiiEcWd/7m+ssBTU/fXX5GHl4wfbX7U/q4rohdWURVKIYOXegTR0
DeYgBG+4xzpKiD0VHPvg+4XLaGCKmMaQKx91XJbkZMCoH6H6pHi1gB931fqL1epL
somvpNnIgVrxipDX3UE8iVySQRab7kD5RVASVWgVb8YOkr7rmSkGc9hgaoaHPfKn
3N/GjqTvdEN0nrVHa7/UqfRR08DX9VGUzZpH/BI+tw+c00js6tJevwWS9AfKBGoE
jomDtBs6RWJhvhtJLT2f5RDp9Mq55DEHdqYPWPAEshsx+R4pTWwA1QpsYShtZGZm
0/zXY3rE3PCOzmIDXpsrDn+2KXArOA0Md8kur2v5o1MNNcUd/Bt7Zt4JAbSdrMoB
6luSLET09ELAhDNZw955dc5Fry0xm70ANak6yFGfU+wYiwtZXkW3/PKz8t/0YZPi
9lXlU4yLMNXeUleUD2xmy/ISBoxsJgYzo0LnmNRcCt6RKI+9eLd1U9yQ83qiSi5C
/DK5QiSgGXxiVt8ShWPP2GXAIIZiFQeiBQnwMx4V9ODaQal1TXW92vUJkUpcNEls
jXDu55CYbz5r4lVdRq2jyU583zA8z50S2jGPISobgN78yL/axz4rsyCx6+f/aQoZ
PWOtV1GKTKmNmhaLtxBOnf8/zrCyGrRBNDmjeBKY/hGfgGJ81D6O2/AzeZwqoEHd
MrygrpMeEntcsSV81mfmB/IYDxG6voIZp2CzfL5MZOzGz5hCHAOkOQ4IU5XdlQix
eF9eWpGw/per5YA9jEFN4WhSyiuoLdQSwhxe9iI8GJ2WIXuKYXsQ8gy2iXFmKZMZ
VzP0q8nCn1hlTIIg/JXHstwpx99XGH06LXtin4Qku9uqUzYB07cd4pNwg/kgV9D/
rX0bj3AilIEJuaSOcFGzxl3rnb64YOPZt6Om2vbi3l+wMNJ/SQAj/fHggzrmjs1W
y4ohCAVcNdCErmaV18xCE8ylp/LgFIWvCWAhYU0JLB4Q77RS4rSVtoG2JVVja4Ma
nl03YUrNukWT2dZkULxkRlbC+BM5k96rFO3TFEVKa2wjgaJe2HjCQzqJ1st96qXk
y+jJ5LZD/EozbRRR4dBp/YGzF/u+vExNG4urtpUFV6pZK+Fa842d/JR8DczAW48t
VrpJDSfLSsqQl+vO8/+GAUvVLG1IkukYkRDbozYDPyvQp2dKQxIuQNA7Ebzs6Fdm
YKnzIAZtT1RFfbiArV1fvd7LFQkFPERUBjC5fwYe8gEGpfigWkLLhwvS+A2wDOFP
0EG2zUIi8vgJafcIJyBMbBVXX3RDSB5NkltC6Pucg8Zug9PwVpxP2nnqWdX/W2BN
t6M2KrPptUQ0krH059KxtqD9sdbaMsbcVxK7etDrJBntqdVsSwYQeNLOzq3XD79G
xzUYN8zuMbVLRHGNWtdR9psbkWYq4ZgJqjdLLdlWUAayoJfxgQVuxWsV/t7AubC6
WmCihZgpKL7fFKicZCoGUsQklhE/DoL1EY/sZCRPVyZ0e6gYotVwGSIsJFUQgGk0
w2SJOen+U8B6Ux3gCE9wgcKInwVREhvmQKEnH1iMaOQFDeImvAE2V67xyzzdOAAZ
qO+kCOIzxAWXItulWm2a1oQ9tMVPc2Pd3WmRVpnr1nn3U5yfGqNa8boDjIcUp7ND
rUyIh346YwofxL7gTn0kr8goyMQRgu6bbt9f0XHG4Q1IgMDCaO3zkBWjxefodmkb
RS/F32yWM981MPQiCeKcyqEU94XKo+eOaHmDtnvuX30WThGXuCAKJ6fv+g0nTcgL
nC/o9WebjCEIiK1LlNlZGU+TBgBRPD0UL1yhwGGRHbNubYumVqFEHUeKT7iS9gN9
Hm1FDcWnFgR/u0BqjUjtXekiGcN0X0RwyRkTmUb3l1WycLa2Qvv/UxnZNr2rDRfs
GMsx25DsibJy3LpCJ/xTTCxuVC2ITxgOEfvcuB1kzwejwKqww0svj1qUjGiIerAq
J7hg9dCJsQH33QnwL/nMPfJJ91W2+pVfHpRcjR/O7wIsbsDDWoZqoo37a5AvKWK4
JV1yVNXv9+Yi/8+N8HxSO+WIQhse0AwrNKTP+q5RfOj5t/gDhpKptCe/IdG0yLQj
Ct4T1V+kx0nuR8s4GCv5zLpieZ2put/Z/YtNyQpL4CHrjOWisatUZpwZK5u0YA1r
wMPkyAwM5djre6UMRqlmp8N3rpht9PpzLKqQp/7vBUrt4jGMGZUayTwbN/w41qMb
pmg5W5OLnXPQnzNYIPxQmw9DbaedaqV1AW07AtivWibHAtQVREpU+LXepk8Y9xG1
UEOl7xKc4QcNMrF24ZCilsfSCPkriFNRSO3AMs3dqtwnQgMw126jRwiu5aBWjIXt
a7BigjFJCIjHqur7lfWzPsLLc/AB9yoGffDtuiDMQ5S2CA0fGwFUqqgJd+cDgUBl
afbQea4xlqM5CBw0CzpTf6RN19FfSn8QXFDQz4oAICa9MlY6bH3UtxR4ib0cqJn5
LoPF6uZILus2+h4TmZhiNvLJ6IpkPfunqSpftTNVb68ZOS11FOoVNFk9kXZRjDYO
TCQf4sUaos9QLEwr8mxl7mofRN1Xu8wJb+/bhB36owxlFCCRUS3Yt/7V0+ksNDsO
q54xl8wPN2PtmhAL9UTJrfv3Un/M82EqYz0NWw49M6Ig17TPTG5iqR27IcPiC5hF
fwKTeuQij/BT7EaL9R8U6E3CmjxX38I9HuCWUvdbsQtUUzlM5a5Zcwx2juZRUKaY
PdyQX58vuI+Y66PQYbK2e0EtkQ/Vhkz3TPuDJ7140w10OodmMwxIW0liYQFRGzaD
BM9dEfaVJEkDqTmleGx2Vlx5PUEjjn6kRGnkN1tB+K3Ad/ywigda2PNE7lk2PCON
pgKWfKsMANHmeGNfqOYoY5cb/QtqxmqT0VtlcqhYScUFJ52faf5TplU7qVZob3cH
1STX+VMe2tV/MvR0zL5CeYsO+PvKM335c2RPrdKx+fENTfYwFSO/Yz8wqblY8fb9
Y7iFAZ7w6RABO2YFaYA3nraPaDTHdU+92/cgstXxEae7QlOfHl0X5QDiloc8Jhm+
7rR/a4M5fl28Y5cQBwnfc7KMNaIkBNWdD2YZ+bu4FTsTdhz1owcG0SpS10jWkkkB
MQDZgf625OvyYiu3CmFdi4uJZPSXzALwEE+4yoDoMiG83rQO5Y8pnfbZ2myuGc45
iW4i7kAmnuwgsPjqIpQ/9X1QaxE0FR4bs8P8vOJD1sH4a3YQlGpUNc66V+/AoIIZ
X8cEGPcI+KVnvvqKxm3HxsaZ2pdUSiZtJRhTHFJlLN/YrGAXoyFP59CH6DKy3dO9
UrcHGZTIQ9hjQYHoL2ug9+5aFXzRG2mHO4g30gs+1+vR30qDIdSJi60b6aSNlzZQ
SOXbLKJ8zEr4p23dTiOuuSf8Ug+FSjJLBkbIdLw1sNeG1+toy0GJKhB67uMiAe+k
PLa3tgRhgVFs8TuMe5P4s0nQgHkSe08lX51mcmK+yLKTn/AbBzZXI/yqLUx2uGk0
Ui7NGh9ann/lt4mFhRdv72ntZTCirAyKFasvCbNuQ1Y9KEgEqEGG//UfqxFhaIva
VjGrYFdV016yobdO/2oE/SgHDkTPbTffnTGh2d4Y27zc967xv+Xm51sPZldFQpuw
d6NnIpRfmXvnEL8kPOETCZ+bjlQRQDeG+qMyca3Hntq1GwFOtNs8JY9RcyMGC/Hv
FHngByZpSV3Nsf66hPC7EFCk+IDT9jkWz58T5ov97g0Z7dEcYQpVU+7ynnZfKs9S
PAVsBeKTd44LDco7u6v+LZuVnm7NebBqS7H2268zwdxjsNkIyxrWHln/NAsJtoXT
IIiqPUEKHwkkKYUY2TneaCwTK+U15m1qOwKCsv/mH19Vm/NYYvoelkUGf43PGOJL
1AXcCMoGUjfXuTNkM9y9dlmerCqv4CUgoBM3/Nt4BxYbl7z2EPo9xQLlazF2b2M9
I1ijuS44CJTuMwvsfuTrqVoQphH5TqfGuXxPEm5U+h0s2uB9Nu95Gp1T7YJmNV8n
EwoBjwjArhfGuaNCTZGh97tC/HBAljt/drjwIqjzP/19chc2Sz8gKT09Zkbl7tEI
eJb6zEDk12A0oGABpszdM+J0tMS7ocA8sy2nXpQabjAQ9mJb6NHOBLE7InmCAWYx
jiBisRFv0ExzBA2/Loi1NsXYDFrq6jMTr36TFc+6O3luQLdYuBF8bMMu+ONRifF0
hF9Fo1arwwrxkJzV00BEoxDj1dgI8r2HNZi3q/Qgo58HA6BzL8RLvl3IrLLEATlT
IUfIj4bjnbYeBx5+ljFal1JqqA/eElQLGb3FjmbL+ZvwAQ+i1w1x+scbD479AJ2X
43lyb/Zxqijr4uDClsNPgvL4s2bbs4yBitgkcbRpf88pK4+E3UUFRfiMHBEyRJX9
WtOfd0GnKqqDRALWCoRExfN1zEiu0liyFVWVlTBsOBd1/i3BEt54mGm3LG4H8ewH
O1sVY5r05i/+dbAzyLvPVac0LC9UkMrM34REU2jZ9VR92pM6fDB0nnnN2mAc73rw
lGoxnoQsL1nmNLsXu69mL4+MRHCoXvjeoGx7Kcy6yC/hApWT4t7K/y3WorHZPWX9
M3SUbbB/pIvba1/ZC9RRxGWQgNApgC/yWYd7R5JnC1YK4KkffYli4C7LzQBfWxpg
cqU08BsBK3IqW9dHV8zi7y9nuYnz/f0D6BxF+P/+/wDFTwOVE5i7Niyewl2uUNss
5uWjFNMjUTi7FRjxzoS4Gbb4zZZ1Ki4mv+JUMtLGMiVH5VLTLsGpiqPCU2SYO/SB
HlGKTa58E0TnSmaEwBxb12TG0O7o1pmBIAkGZZ5Z7c/Leu4hwPmXn3miMfvudIf+
dFroe9rFKVFKjRb/pY4PeouYjmoQlaPL5y3pZiB4CZJTlKPBuwy050Bm4xRPdqb6
/AOGjrQ0ImK/wjuuWNNvZQzwefcYCD7bIbbujvq5zE/ENP2XgTCF5YKIJ9UMd9Nv
L4KdSGne5FuTbDAAbKeVghKziRr3uhlA6NlzNEW0mx6h4+uJckrRIPSVQSqBUj0l
RjGhR8An1wGaesIRRyVWlbTJ4ImAGQ3az7MVl+fPXm6t+JNF1cCzDAtpDPtYJpvD
4uS9zUy7kf/A5DaTA+Jp9PXoJ70lkQdt1fKPNpCHKO4QQ5RQT14Aq8tCPrJa1SlL
7A5CMuOSaqz7LDp8cpJhmwuZ7PM11J6bONfbtUfT3uXafZV0v/x6odTIqWqLlyxr
5qk1Frrf691L2E/5P8g1TiY30eV1j8HL6+cjhUAtWT06DL/sr0UQX5rIReM4gKfn
yVGDyg5HVmF8Rq85g5xruYaMEkED+n914h0Y/qLlVJ04Lweyuu8XzxYtS43Rf5DC
x5tPRjj/wv3RClL7SYAj5EGC3vE+eZTKyW4GNBOM2MJ/NoOR0e2mnPGATsfIOQ5M
MrrMTDTh4RSAK6FHyueOpFrP8Fs6XTmUcIRDDSLzVEFZbBIfdEHoe+YS1BZYLdH6
Ucq3RFQJ6CBEy3F0aafhKLy4NM7BCD3AyLdRb83qghyqBAD6VCy7kCDP6VO5esaK
bJKyx5o8tnLd3IzVnwdcLqy4+7migwkkLnOPaop0iW0AS6r4wYB0qptKdqXXiMOD
k3eZQ2G0FAS4tASaW68EP7iiJVfo0nU4Yq4Yn1AAkfnvmJjOHzefpXkp5MF9DQ4B
r8D3LuRV3a9kWkFFe0+7ci2w6WIqU5ocwQHlHsOtyCIV8eaOltCq1ZRBVc24I3L6
LahCJvxnpDdgiJkTDAUpb9E48MzHu/bu4tV85ChSDcUUAjYGej9o/D7w9UbK6NhY
X95qde6ZmLuXO/Zlw6azXLAuqz9UfNFZPXUQcwKOYPuuHoVl45ryTB7Y0lSz1u6l
w/14R1EyfBPh2iWNDXg96HOh9i6dj34w9Jo1R5eNABALN/bph+0bBmn1tKSzQwnh
X7WCrkz+00ZFPItLv6wqkq5nxhACSmFS1BU/qw7A0v1alrefebb0J3x0ss0UtMWE
QnjqVjrSguunwVrHF3wqg3rLhcvsLY/0yRIyE/Oou31tS2+NrzQV45wVVd5jU3lZ
3a3mucmLQAcgl8yBRY8fqYEikVVgI7dtHkD1PX2gfGJ8JwyjzWq/5GcaJm1HxIY9
4Cnhxe/JD27Ih99CSnnZvvCd+bZCEj5HUmY67Kw/nM0jveWhOpPxs32POMuFUn20
R7CdqFyfUdVmBrHc9hiaFcJlFPZjcxCnvYB8HcXhhZ+2HSlJKhgdd4sj2j/vygJK
e/QV4W3mZdJMGra/RCIxLDVGwepvRc9BN60JEgDOj/RYNtcYb+17DaR8dDyuefq1
81cTKG/wCeYfJ/oAABhNXdCjQi7rbYwK0CNuIjAWdfi/Z8xVWX9IYeEfnF/yrPSd
Twaazs2Uwi1MGVm43bnu/Qhv4C1PVUA7R98SGA97gMqUjVLWvnJCIlVnOCzB0BNO
lNbHua4bc3l+kSUNNR8Pf/2E5uOLdabw0MlbYwZcmiVIMWsSObDF3SMToaZnDdJU
cXulsgbN5IkoCDCjGb7LVqT+hm37/v6NDDCWh1a+Qo3XHyXTU9p6Z4hPS8uZzhTM
JUJKazb95/95GzRLS+NbINCHe9V2sv5GituQfc9BfDK3svrtLOhM4gwYaZjzzQBT
Qg6kW0JClA17pTbie1cOwVskm9+iGD3jSvNXpSaEj6BQzPeJucqK95ATcbPAdbYp
i4eeQTbfDwqIXQ3f32o/VZ9H0O60p7mvFfPRjXlqQQ2mPikIafl7iw4cSILyztee
frXxq8F/NVVvgCVlFk9zcf2+ziWqxh8bEV0VUbyfK19zSNlb/OQLShcmcfHrrf/i
15vbtubz+846WZAKQcEicojNP35n2Hiz/agAAtEbml8+JVbvKj6QQfRs16ghf8ev
BzLhO24ZKsY3oBL7BTqLy1syi63JdX3fk4/jG7pyh+otdhNqysZ0bBAU3GZFmy1v
cfC9kpmTxTRuToNMuKzRZJxhWFUEcNMNfrzdgmzsDAJQ0OFl/QiJbFt8EWibfran
dKkh8o1N0T26RKIPIP7NHVeKiRykPiIk0cZpvZ//KgK56xVXPEqxaIxPLN5YgsF6
VXeCYKWvRkTnoIPaS5u8rLeVipQvtEE+gqLdNnMv1VD/wG+YUfYs6aeOvdBZ68Cd
hSbX3SgJdVeFLrn/bX2l6CJvAC3MKLgykXUF2bzT/WFBNSsYYTq5EDixxz62MqwH
UMhLnjFJ3mzZFvrxKQBNSk3CPChaN0mWeZoJoxS7WX/Ue/FgdrKydF0FnTmoGP6X
68YdvfSUfOOQfrX3clJ3+gxESElbH86Xm279TtPOoJJLj+3CiLTmCB3kGBKNmV5v
XuVZL5ZIPrSy2gsZgGh6LKyMovfc8De6kYxNy9Yk5Vyd0XBccbqS+vk+rxiJ+ygM
tF6rpi9XxE+WmhHhy9zrn+0pB8jEF/NUSPE57qCH5i/YwKa6wgZji9MVbQVJbsN/
npOGjhwxg+SnvW7NUq5IKB2xcyzrvGX2/RruS5F+zBYe7uJFQyd56rc+DmMpkJnl
hv/3XUOgP7y+jksE8z1HNnIe0VbWWyfi8WNpXFsfhyKjAb3sFa2ey3eZiCb9Caqv
yG/5Rg9nX5FWOszX8/rZxZ6WaW9gJ1cJPslgAT136H0BUPcBum00jfeevIUogjpz
KEjhK97QGUN33kefNfKJhV8Yi6A/CmeOcOwQ2zVWZws8Dg8fl5YUtPX2Q2eMXF3g
p/F8fG4WFhL8quAYAoFZSXv7p7OXoW0lXqFx31IYGbZ4hbb1k7dYrOdUhXUOWHxb
Ml4wmBsZ00sQ+T03KQK6FO5GShI11dDJ2fDaHLdoRlc8O222gebeQgd9M9cRjaAy
IbySdU3AOqIpHG8UCZR2fMZOk+n3jan3ubCSvhW3EvhvKx5ebw4XV7Xidqo3wQw/
8+ghl4Jzc/WPMrfzzHksN1R9+2sjyF+QUHjzgZc2CemYRqhCBmrDHNf4dNZ43uyA
wEuSFIHm6eKcw1XdBgvJan0Nq51y5L2+ZyHxbbmkMrRGBfGn8guSkwcEA7StfRgv
ETHowdU81tUF8VYGJu1ESX5kqbn8s/8SoS2UN14MJq9Lrmm9SY3GbuSnDjUHL9xy
L7l2gQIoGt8+OpXRn8BedSooGJaXJoWjt85BRy8B14i6eGBbGKqWTAwblcApcZlr
1fZm9KPd5in/kn3ZrOHiuD5EommcBTHYUR7f7wM2q7A9NSQsG8rzvhReB8XOu8tN
jAU7RsUmtFC7dTIjQU9yFKl8nn15XBqtUXjURHRmSmL2iegUpeE3+BmQUQJGPLUl
zNJwQZKQgW7yujc6RaIPhC3ED6i1w90PSsFLzGHceouAqxK6Y2trH5NXiCmMfg7R
2rw+Jo9HgNpgBgcJ4aBukC+IGXg1SsJ2Z5U0J2YQBKOnAvanT6XyxTMmE8U+dAcZ
i2wz+J9XKAUZKnMjF3Pyek9mfWW6TkDVF8AxumFOl4Dfb7LkYqOvUOmB4ECN0Ird
TlQwe1xEjcRj1/MelJ0kY1gnGxndVkrP+Hy7sQW0kD6ft2u6wJuS5nwSyz0mmr1p
aYsiewcaKs6ZfAbc/oGqRObl2cVQdKMSHP/0oC2X2+d6DhqHfPYLgYIl318PZZq4
cieAz83KjERFSJLQO1ClYgZjusShvI53myV11x82+pi7kYwriLQ0u7Bm74DEA33b
+Z2Hy84ONWThBTnh/1KUadYmaeBMIv+zKDg/AUYAC12LJm5sWdSw7a0u5c/QORLu
bS4DUB1Q9J5tA0MWe60eBHmU5DIS/zojXXgXb3t+ModqjX6bFz9oI09+4rlR7VWl
ggMuxpV914jtFiBjG3i228i0fuaX1Xz9gD8NjsNNGhclU5wxUHHc0ICfajox3ckq
kE41GA4mE5xfYuZVal1Kw0wR68mO4GVGuHw5trSt2Tbnlf22ZdaaCD4EzUps3Ylw
u8xP6c7HndumbsNTl9Z1jtVveZM3mVZVjmJbGxVrbC48sIaNzdiOyjvzPXsGQwIx
uDM+aVIT5jLcFLyzgpzJUAqpLf9A+KX6dIVDBleVmyqXxXhVzfPmVKoPtikzijct
xmUvUNc6uLr2KYGnSJvknarlYVkNkGpVXXZl1cqFZRQruoFYaluKDRXkYdkOash3
pkx87T14TIdY/MBcFq2H+xvjbNzd047KahmCgVAgKcMN3pvGWPXyGuyhpM67MVUa
nzV9F+VH9aPCwxTc87Y9iBjRi2YKwNzGV3eB4OqaN1Zb+4F7lxYBRTZYln3GTsQ8
yhSDcVSQdFDAklmvDwlHd/03ENUzu6bZOCQwJiNlZC6Somk70gTSSowxLVOteD5O
zWVLdusKf2CA10x3qElPYdQdP2zIPNFhJeRIVioyeQxGF/2PhrszdA8pY00THTVY
ahNbhtcsygZUI4naDawNNMCCv7DzL5Knm13vaHmZnGxM94nemWKzT3ufSxml2xlr
tbcyy2t4s6p9oh6G+izjv7oMkcmfzG7tmD/HUm0HUBBvUp+jolJtKV5ETKrZErNW
sO+FjiTJGyIOLkM4gcyb8zPIE38C/ZfTMmWYPHgVUSWQ58lhiQ5iFRt64RdVAu9n
UbY/CPXcyrRGhKae/h8qsIxDULSqeU+RXgMD4WzaHnehdgLuCecn6CKVcoU11S5B
GGGyPEBuQ0KkfrpFFqcn8iI+I0d6uInMTBCfgKoAAF2CDF7jJfkeni82X4hkWM9t
QFx2GDntoX83cKUBa1V8r3UfTtpoiI8p4cTOma5FW4Auo2L5l7kYCj0VMrg9yQpc
dwMnlEcEeKkhlZi5a9eens2IhiFu1UhYL9Et5abBFc92zCyoIiUY8DcZJfAiQWSI
s3G8cnjKscLfwcYZQ6YiUuqp/D3tEaQhRSS0+UGK/0R0atYiNpBXV4imC+fzJKHS
bq8LiXM5mxIbeDI94TPMHrQDvgN72ahr7RF9KHHQQ+uo9ejdavmHNHyNz57e86gX
xtWhBn0qHVRU7S2tDWAEHSuGLz+MeC+NTQq/kcp3VCc+xY9CyzWzJK9VYJGIo/aO
uvWR9s4A6U6cnJByxZmhPM/ja+8GBgu2/XJEChJ0C/SGaWlrPmbMvh1bVfG1N76y
Xs2/7pIwURUYIlpsyVFQQIQobuHSWOeNmusdoofqyMU2MzdVNVaQ/blw9lKn1uQZ
P6N6ZdY7C5N0jfsKK21l08rqHXibY1cpgj0iR7Ge/jBuwZI+mk4+Ep/VIHsXn9LW
51w2eJDtfDCltIhctNkIwhpFp/FZP6EDzWewo4SdSL2mjQBhPRGEnKmxpZq5gr/D
qH3C+hmGk1Oqb1y9YdZwaRzoeO7rhsk8ilo8WqHXZLqqAkh8Y2xOnK1Nd9HwXbJj
TPoA1r/j/8CnsFaf0Lujetv+V9bS7MMoEIlFL1WkCfC0485AoztNloqIo/TxInSk
Qia6r25mg6axTR8L3P2TFOBMbRYFIU4QctQ4sm7m7ZpTwIMF597pz+ffXE5IOEzb
oBgqt7RiauQftHIcQPslOPFYqISAAgInMusERRUJHuq2Wv1LyOKiiwqqLLVHTj96
0w/BC+y2Bm83CPhxt7NW7MeCNplyPRkn3zLW9ht1HeCajXlD67buJPZVTj4KXKZo
8fVPKxe73TXz/5fY9Qb87SYc1zdQft0IalrBI3HpeN5qgA/tWl6xuvwsHmgkQ39A
MPTmZImtcPvW9MHQBGf0xUtrfWxw0Mnbae2ySv1OdUZXuLa9v8cDbMYcWQLTGDjo
RGSqKVhZaS/tAYLAoMoe3arcl9hiCsHcyc5/Tuu1t1gmpFsIxs4GbAl66qh36/ZB
BhKxOE9Qt3NlUKTKfk6KzeFnN6z6D5tEs3pZyiSH56OxPhls5zuCvxrev/k9iq/f
UXWAqor+XrTbtgi84Ory5dqFHZgegYo7PnxbgNyNpx8l8mD6KqcVHP0zFC0Sb3Pf
Glc9eYQk/GxiL1mDeMs1UAcAYwoBCSdQGhoT2+DJp1grnZR94y4oNcB0Xmban8G8
lR29QUnA+E1JhtXq7q3N/XdJDCOafICYCGGp855k2UT5qsunWuPYNSdT2C7Hq0gu
xooFh1YOfszKufsq9vhTG3FRBC9TNnWE4Ggus2fyMdMkXUn8kxpkC0K58N3a7KQM
zx6DFQDBrbioUSSulEbhcqoPXFNJle/t6mvWJk1hz6LKU8sNaXFbtX6ja4FoCqgx
ZRnJtpWtIOnxrCkJPhSfXA2PVKxsgrcUmR7xv1O3v8xS1ra/OvavHM5yw0JFa5MW
6e+UohhrvkSMWLIncj74LfigTAAd0ykqKV7vVyvuUbglX0wIPsM4IGzSzujREik8
hdKzQq1xT+r9G0oN3dqkDSJGrMuBhXC8scIviO+ylsx4QSP1E35JG+i0B0vmCwaz
6GFN4yBGMx8cZsgkufLnLaESNAcJoGlfcY4oGigj9mynqjmfO0iJdkRc8eeyCJaf
JNzxTRz7slR1bBQWJDBnVOVqAmw7DO1FAtX+Lpp7BTZgQHw8tJpE/2koXYh1Dxn7
0LzUNx4XtNuPhy/UitnuK/oVw2mVt37NCWoqsDUMsHo6d1DyqisSNylDK3BFdjqU
HdUcG3Qmk1o/DlpxfpTdCme62+s9/YniakgB45+n+EkfqRAdTstla7rbhHwhcNxN
yGsHjRAGQxasAaT0wkaOrPTgXJ2ob/SDxQpqJZrmgdGgDlkwEZ+06yIH9FH46QMJ
q3q2KUEkWmqjD4H40wqvPatuxRnsVpGG8uaJB/rtPW25RfOC9WUoCHuy8nvCYN2D
VATTj20QON2Qe1/NvQ4K/0qbzS+YCrdFy864TPttEMo+WnYArJcmiWM0GoFf3Hrl
Lzg7XCF39vjDEg7G3CWgRZ4QsDWu93VBaz0WAo/KnaNdy1OMAStTmvovFtK1g5kD
XnAX/1L9H7suf+rsBcCEM4Du0W9GADDZ4KmIZ8uzyIM9QzfvoEaCkpAhXHR8xGED
QUiV8lKC5ziYcOvmjN9vmeNpNV9I3imaU3cgC7Vdq5ZEzFy5ie3pB97cqCyygtS+
NcKrFOZERciv3cqEHiK1C6mZvL2RPfhbOzOpRSfj3Ttkn/i5qP0PU8mR0wotFvkS
bXHlVjfMAi1yUnoppyOdlm5i6Dwvkyaa1soNK7kXv0okYsr54M7mWnVidEAOc+dI
K4LOoqiaAYs49IeohneBc6uilhYZEtBVDUGiMfnowPoR6aQtTEQgiGcui9OxXnJm
cPknioxbRU7v1sKGnMn4Bb7pKpBFOtFcTZZBurLZku88YOvtdHCs9bnQENiY4P4L
fYvqr208EOS6Rm3lOaC64ef79uVYYdkEXPHX17dSmXf3GdQR3Y/O5TjAk1FetwhR
dyL4s3iEVTYDlXLbvRlu4HgvcLP7lx2vCbGgG+ju72m12tkriRT+dAjeLHQfRUIj
/D3BXFBuNuSTXFhktwPM+K5WTUk5Ivpy+pT89zdZXyUUzHnsgYdP+R8eEV2M7ft1
jYje94bBxLSq7yxB+N9CeonOtHeP5i8ThAM0/HIYS/kCtFrR4ebZ14777QuqvnQE
OW589UI7SjgHYUTliZMmtj4iGUSnlFBmqiUYuJIOOGp6ZwxWWyBVa8rgLYFoLCHd
dcoUE+IKzzLwxszGAfqTGu6Kpfc27Nv4hHJGn3NSVTPkaaIHxe65S1RkA9RBqNnM
Z/J8etokwytNBB2J//gfPpR9wJf0udkOfSzBB0yrt1VKRsvadCa4o+R4nwTv4LmV
evLI/u3WfefNpAWA4dmHHTDi8j5KTtbdY7e2utF9H7z6X/+RUHtyGv857BEOHlLr
3hvv4Ur2LIE/aZLFt22EGMonlgENPq4jFSnPPmOpFYmVPzwuhzqs0+xiEvEpCF6Q
85La6kiw7I5KXam16OiNYgNF9ryY+RHV8PUp4TjG00jSDXiyVTjeqatRUl5kfdyp
IYSnvdKlZ+XDhxBf0OLoq/krlUi6/H78seNmdxOdE4gm5IRUeg3yDVXPrnYq4EgS
NdT9M8QA00eeSrhMshzLGrKpv/y3XGv92AABIj+WJb6DIF9yORe4AZ9ERzOOAuhe
bxY/V5sPj/x7yUToPVNDpcuBby/ev3OJt+PJTGa+pdCZOu7BiDOX1/9Lck1/2Mlq
m6+GX0MgG5IsJKdlmofeA5qv1QOjgZbf8R6ltjAc/MaEP68mgvZcA13+bZQFYpvj
lvksQgPoGtwlWvTDAPRjKg3OvLapPzkRENp1DL6f3HKN3e+bCRnf85e7SoaOKD5f
30ifpPIpHY5sDfBr4BYhLd+lOe8gCaxJLHJ8wCzKhOTrIh5MJs95cHAAq/5Tl8VY
V6nnSz41y1V+51/TnSJO5ORmY0EkcpQUs5ZgkSLqfT8knxJzlhiGko+IcuDqy4oQ
EyZayczH+B61f3RuypTOgano2Zx3MkuZ5V2qF9UC9244todsho0ZurKMTvj/SDPq
s6Q/bPpkEsZNOMvIkh4gduLsUJrFPr8PsMzIlkDSKrwN6gD+tBE1jgktKy5YHU5y
jieRU2ULaSAo3JCOPv/+m9I7CRY233YOPZ7DPhbF4mZoJE3gSViLY9ooZdDjg3oh
swBCIw02qRLFJZwzl9scYFK+FhL8z4wYzKmRI6+QGGk6M7Jl2bqdnanMjW7calzb
pmGFM627yPKGDESSMUKZoQWzcS9Y0USu1hJBo/1LxvP2iJkiQxA9Bd6jU7oqjMcR
V3yVheIh4Ms7LvzB9v0paxqt3qYvD67neHKmgk3rE1TAvTz1thXF7rBTMqU9f98B
g9bqlgwbu8fq7PuH8d8TuQXZQVSNfv3fsQtvOBOrv3oc4PkhG+wns01zh6N28jW7
2ytJDkhkUQENseSJ7OEXOjoOTPiFH+g8/2NlvvEUh8dbPW/O9VGNSRhDA5lmDm0j
9g2BSQiRBF4g+J8o1tiG+Qzou1vhk4PPaZc2bqHKSDgZNKCPTYmv0DGQPzUR1t3K
MLMsQAZfadyHLHcDqj9keDY8SRKeZOggp7HA2WA1Wgv2xj9tSQUIyxuNvp44gOrX
oMpNGQr2EMQ7KZK8On5TS6e4YQbtSjmEWPXRlcDw+7kLZy2UetX8B1dnrp+yUyyz
xbaXsc3QvqBDeF5zDXcwAG85q250Qf437xMF723Vuy5YDc1eCzbkbt3X13M8LaSm
zMhNSaImy6RMeh+pak3Nxwd1V213ZJHnpPVgdYvtj/cO3G2MF8sRVRLtZVWDbZ+D
rK/g3OyhG5SQ2IrhrQ/UvSk42WGM65QTWkmQMmz0+C+2OkRL7KMkMWIM6f6871E+
k68/ocrKgloLe5Br1b57TbGPuTYZsKa8ewixxgKTgLy6sYIIcD50qD79mYdWstks
A7tItVCv50IgjYjTh5uy+0jvfA/tiDL6FXX/udHXkFK2kDqrPfX7VHENZikN5Tk3
6iXZePXNmJ+4MjpwoDV37LTq+d+wOEjxToGzL7SFOna/vAwjMXIAnvGDnCzMzrP3
kT9QHYpdMGlRWDeVCOXBb7OnGctZKPtup72BnYHS/5NEG2v8jbJNKyJJ45HGZ0fW
RK3AFtptn+ZObK4wVKgO3jlysQc1CKkFPKSG+Bh2ffgRrxcpgZCBSzDEiQI+Tsz1
OfCQWlTG/xRCD5U1vCGx4NbFhPFfki6jRjKdEVDuDsjdh9Ig/XrTnJm5QOzwBY4X
+Ta3sQ7rKD6G61hg70QC+Zny3PsrbkQX63njT4cpfWoEzYcwz/e9jPS7b4eGia5i
j2a+us/Xgm8DcFyG5r6aNM6ld9V939ERely6pSYzLqC7AY4wGmU1menCneG1uVmY
WTjSSmX9dT3Xb8pjiFcy23Zc+kkqpaqLaKxuVHXIDG0OTDthgN5TDDEkXMc+XZs5
iyKrfmx9HIy/ZSVMXy0YzRNP+PnwNYqaWkHtfs6d6GOkM2E7z7P/KRpjJ7SYVkps
PsIGoxZkddsf7/nLUwcpYr8Nx1hS94rhrUK6kLjxf6KWGqLIkO/gzpK1KfgVylDf
qBlPItBT6FtunMFQa3uVH1FajTUYzpyQQK8V1a0C8jcKtdLvuJBsP42afsBuBs8u
uJnemAJQi8bY1X2zN2ZM03tb51v6e4iENW1lXsJGEdWidY+nzfBj4dufoiih+KP6
KWC5hBcIGV0Xt+2HVXAjvx5o4dprMhhUSIItWGwyILLGJ4nXB0B6XDTTGHzlRvY/
aoswtFYIaU9qoRxtLXepcRG+IDgbWfxP96V+Q5l1hbtUTT4NhNzL2Vi8rSDJ43nR
uUUgOPSVJ6UN0CZrgUs42TnnkUrcVieu5edZAlbdmJIW1od7nFHNKAlKd+QCc+He
I3PdA74pJIq2GItCYr1f+eaQKh2QaKR3XshV+NSRFbO1jOB6iQawXx9MrON8is5E
jRkfATSM+rkVm0CSSqZP/E2bW4CM/BwywN3+9BHWvgE9IUwp5XsJ0k6FOsprMaG8
8Q+tRw/o4+v6PeGJjZmVNTAmIwR3PqMN+StoB8L8nRLUW5oLf01r5XCocPqfkUPr
pHAkLXeJBu7ojwy2+BBH6ePrm8uYJT9ZtIW+ZeGaxX5iAMGDmWVdByA7AAiIzJl0
qcQ0S9PHiZWbrbwZw5nMIQ1yl3JWNXt72ceaAm4lQkNspOICfsXAEazbxLoVQNJy
PgNcRS8N6qgerRCF/7mwYiRMsVv9sINOnzqGKIcvW4fEGMAj69s8JU0cR/6pKmhz
E3a5IyCLGchlrwPdrVwJ7yoeuYt+56GwQzfBJdVJrHjJZACR4MqbLrFzBWAmzaVN
+fX8mGknzZpxZ/PtvRDpLpGGNasmW3S4IiF8nn4L1c+E7QNZ9fPGEWAQ9Zgvly1b
NHOKvKPy87wLHStCZrDqEDwFknO0icuCivgV2c0IDlWgZgTnpzaAtoUvBIvzDc+6
x71wIUlFlemaKEdJmPm7mFcoLHFKVpX7bskBUjapM2SY+HZDlqUGv83LvPMRkGaN
syGFjG1SOmCdNNi2Rkdfa3/Uius9KVmlZ5kzeqMytHsOK9FjHzfZxxEa/NXaF0E3
HUpH0HkDIRfKjJY0Zgxz/AUWqZ6JmKs8HcOTgjWvtAxuTuFDnSTH4FD9OEdhxmwt
EdpAnAxw/Nf8iZFGFcmNFJTY/VO6ngdvhw52L/U6kD6g2CBvM4EHMIP3FpGleVqb
3on98ZL8KI+sHwDHtg2rZA6r0kqesfwYRlZnkHtEDQUTM8TM/yQrKGl5hrCcaIYp
45tmObi9Bjt+31DP+ZDYNn+WE1oJLX26AFn0fNfmDmQ0/rfDBCM5+fmMXXfNKjgI
xcn2HLeN+mSb0fb95Z/z7S27OhdiHXB5WNeFa58wqn+skGjWMi4ic6hEWyAr7Bvw
Kr36D8aMS2AfXAVK2qalzfDJQfKlSMaeSw3lBxLsliOZNGRJkLxE9Tt5tKRBXGlL
yfdjNOfHev9nNBKP6SnKNh/GANM0eqZOuttFogCO/SIdYhNr7Wah93XlYpts9cIx
Dm3FzzUF1qXU8KxHBqHDedUArFkCaoleIjoKvs+oHo4LsSp5+OFb0RVlgBRa1w3y
ArOEpGgfTOcjQWKGNTvXuLvWNU3LJ8MDYbeb+x882QkfH9v4NlOwiLrpa/d/UrUh
GPEUVO1ObCAamFVbrScekwJjOX6HYlZpPRsNK/09hzJNr2rwRh7VLI9SxASluoV2
oIt79dVO/N5GZt47oTLVIodF/3K/p6yXhOFTLeBNgOxVp1lXvLZRwzQH8MdxuiGo
quddLOWZsJXfNQyjQR1qo/9NMi9soSdP9uJayNsE0TM/j0Ti2EaqfEDkR6Oaa9Uc
z8atohn0hEzTIAIY903Qx3CDJY00cwxtT1I8zi0ESQnBMKvBE5bGNy83Xhok2wMz
sp1K/fbPlXoXgoum4hdJSHRSEGCTW99/VXjiPKS17oBaf7g6j9rPNYllwLgshdj/
CkTItErqYrQtsS9WyA26NvMyc5Va8lHeR5EsMGgAdwypeghpPQxHLLZpXdWjZY6S
yjiQxQDpa/1FrEZB3CZE6+4qbWBTxo6VKGfnt2cb/x8MGa4CWhfwC99+ePWUTNMq
tNT6LIX2Psme1Wdxwi8kf0gnH7hL4jdOL61a7L1xdgn6IK3P7Udpe/U7DOMLqmux
0WuVfc4BtwEp2NyrXoD18vR1iUhUuh4daQpmGGYbqR1BTaOGsv5KDX9+U/9cPOOH
BmyNS1ZjA1LGb7wMxoFiLDt2EKk/KP+JSE5adhwgq0ekechIn66eugGvRz7FFQws
Ycc32nL0JWM9KSHUL8MgwPxgI46TvALM8OwnRv3JfNA5FLNoK6hBJxGlIuPOan9Z
nAsqP0TpWWDZ+H+A8xhj6lTMo+K+vIDk5ECv7188gZa0+P4eXliVrJpHObOODs7c
n6nGVPv5ScAXGZcskEMKMWwaCpO95Qa6WMLYo4/1RsKq8J+1i3En0nI23BD4fVvV
c+fD86MJpU+X8pl+XmmtGzvXxyxW2ggGv1x7gYSwill7d0RDRrt9fkByEM5dC5oJ
RQeOaRfHsCeIgSqaiOq/0aG2pSMHzM0Y/PxXbSQ7EPcsu0PqlORTnskUEzielgcp
LjRCSahO4Xc3hRPYDq9zKMaNTMlpGUAXu+A8ihuR+pTl7gwRGvEls1O5gTDooTvc
mtNdXyLrOY97YUPPcxNB0/0fDcqBxdh7flAjKWcY4jndw5NTmC5Yu3yDMEaUgMOT
1R7Ct609rgxpQJWCg2W+J9BkaeIhqyCvBeQ2I4vVNeT7gWOLL6j41AEx77dewvgp
DDg57PszXk7Ub9JMu4n2HRb4NZ54ykq4CnGRcTjFJsjLylWSvcD0qHSabfLI8lNQ
P6/pu4zHlo6C2h5Ycmq2H/EQefcD3Rz5rG7GGBp4JrADRnDkZhJQD4UOtR891RJF
QtB836WC7S6bu8eaIFodg249cnHNCXJXJvnKM65XaIXIfFwmFel2o90o09YZvGMO
PPDTS/fT3F7q6nlrY9XrDkfo9epLocpvUETB8lY+63FKOaTK93aOtcfZWMP2rseu
UTAPE9/ACQZzrL/pcfsy3BtNTRTfWs2T3WB++LJh3DH4FpoVAHsoVOu+R88qyKLV
JKh/wx5wxhafMFfA5G2FaSAlWkSXvY27DOmn3SzhhpjDv9II6V0UwcHT5XI0wo+h
LgyVjotgaKqvRVCGhLJMXnAvNUHGlbjHPisJMSU55dB0aH7WXBMnSGj0+bbh8lyz
CESi4VOYtCY2LKOJl3w02zasXvMLnDbMYKb1CuxrtxjLi+t5kfvlf5yLfyufLFIM
uhkaWFhN8rJQoSDg18OXoYyLxqZTdeO1M8zCTj/gfnZNoGLir4xVpj4YGqDQpZf6
WKbItL3l24DfXSytk4B0LHwbDqezxgRiseIsRq0j6CTs/6DXBkU+EOcCwLT+TecL
VX5nmfpWALYBKQSBr93dfbBustiXl4YfzJwhaNMttqBBxoJNdjfOl69jSd8yF/Xy
oZSKEF/6F6a/vA5JUsa/r1e46kOK7IjP53RxKUAqlU/ip8LfNIUGWvRMoyRswBqz
JPx9EVtbtjD0lqq9Irmf8caz9R/M6emStm+2XRpunZWvSF5EdqEshUOxO+B9VfpR
btox/HWhR1Q3KL92MfCclv3GVnSwMHpN/bgIndxbuNDKI50IYrhODEncGFiVxAby
3Npn5gmXePq2vlzntjMNsWfJopy4i3JRGBiUtivR8pPXb5SXRCf7xH9rwpPRiCra
8Jp7N7pIQcG9kreuFTFM3jd2By6RnEEtIxNtpFwqyK6GiwBR6ts3kVc2y+SZiT2L
AT6JstVC0bcHiG6YmZLx7va+6aN9k8dW6iw0YD67SnlqwI7wDxLgRQRJj/Uxlm7l
KaZ8bQQ0DmnhZQfMjfHTYMeLaaE/Ti22EKiGGv0kY714ZUjpMVDJT/yCaFVlL2fN
88swaeCcfTb9vVlHSJwunn3VU7ZR0ai4yULhqGTTEFefipxZHYP9vc+TKRGB4lct
WR1QRAB5qlEs63Yvrvr7tCE0q4wqU8vGvNiOpotnwzeycvhtYcuHOpkFPlEZ1WcO
W7IZvgLOSVd69BhTpI3hcFix/QsZuzNhl+jPNtVjV0qJNU1NyZZdKNE9hm0pf6rU
6QUxjsZ5N6sbfNXwFkc/zu5oFCzC0jHlFm2drpQgFeBNtq2qQbw8Y91K84k5xJhB
Jkj6C8b748aquxJLQvl6BamSiubtbcWjaTaDNuSInbLUwx/sV9RAQVI1BH7oQp6A
HfFPkiiU89kIk8bM2aPDFkzngeDxaVGv/tvphl6ACx4flMqNy3I39e/n2V5wbKp+
giM1Nogvz6A86KcD4B/Hsdj6JYGd7d0vJAJ5XCEYdy+fLBEm9HUF6GOTV4GUePzi
LidmRVx6+KvUZnvPHlNufwFkhJHxLpbCAyQaA3Ipn2HLE8eyh6VVNy1Y612A+Yo5
mUXrCo41+mORU6RRCiE9V9+JYYf41Mv2JRPTNuZtQxYvSq1ex2dgdnbecXMo0QUu
v7wwPgghnvAr5KtBh4dw4NtypqrcQ01JxYqdPahiocpPDcqWcQEPlH1aI1Oo4Ssk
kDXVeqyqtbBZpmhmJmQgXUTupc5QVCgkcs7fuin3I+qDErBb2bTeZszY3zCYt4BJ
QGhf0iM/h61MoJVImz2KIIjnmN7sLS5Sf4uHj+/yBZPRMmnpVR9ELYxPtIBJckN7
1qIkgz+P4D/IIieiyq5see2gzalXGmY1XZzwBcjWdX35KBRiNYzZMB/WUvEsVsAL
436vJGrt449/lnLKfLPGmIfUIkmm//M/mlxi2bh3aP6IVaUtl7b8l9xxmiJmtTS6
cnf/4f/li35DhLOxlE0ZarLnKQr4CIwz8UBwZmZGvPE+BsjJP918wPFcsLuKFrzx
Tfa9Cr3VKuKIsFkqeXs6I3CXvM4B4LRSLbk0E78tHRUzC+mH1IT9PweT89rucVUx
gYY/7UVolT45q3HmSK9J6h6T2D2KPdzihJ/To86rxedQsqidXMQU7AFSvGt1an8R
6mjUWsNDgV7oQRDnUk91B7gSbMHRNGjRHbERtiWTkUNSEa9Ntj5wA8IvzyEO+AxY
JINDvHTL8pAUu67oqSeI8f4YdHRb4JHS1UU3RmB8Q0Wf7G7ZEq3kf/vQsTfIBDUP
Ea9W+vUOSeMHjVOows8lFYaDFUE0kAQOjgCWmsyoZibh3xDBsOvoD7uS9sQroMEY
/2zwk3BDmYV3SrcEkLfY3jH/olOXKJ/ItyhDmiaXYO9vpWQYZs5m/O9i4qtSIBOP
hhQT3vRCVpSOQ01kwx3+AI0/j2VmveC+ACDY9/ntNqVGYiL8IxlTis2uhkSsCkLm
hztS4CvgLsM/pCg+O9cD3NJqCya7BStuODP0dMydw7bDwpu5QPwiNj3oqubFZdBh
RuftmvgMzKAb00ZGl8kNjFJSzeE3/Rv1nn6uqYJ0GgOecEQBdvsMpma5atcFj4vM
AOM3Bdr67HOnE8wkFkOSVHlMHrhCV9pdPehNPHd+EuMoUNRoF/W5rC50AJFS5Q8x
VKiYewKjl9sZag+rWkM5fGOnAjlig5ywYeWUQ37rGz2LPieVKEFaHyC/JL/NlHGX
ADBMKyxcQUdL6svQwK4JHtg8XwWMPKOndcf9EzvmsOii51KwD+gYWaIpyig/iuxB
p37pKwEgc40aV92dV1MRb3kfXE/prak7Y1gWM50LGJeNRgOiNTuy8rv/Kt2HU6X/
bLSrCHcaqEcA455oaNCMCdU4xwyRgBl10sXa4W4fJUu0F2p0xX5GahB4EHPL3Ozl
A6U5nyWo+yjIEkVmrFQbZHJI2vRhuHQSefTmm0Mz+43JZTUAzCLWiTQ1+i5Olo76
dVZHv1A2J+TYEN7xIZG61PNNFCjX6AWZuGOcRDgBjysvw5VIh+LgKgKGIx9lSyco
AqOxAxz0SkLnUrd++l96131R0gtBHUOo/dMF4eUSjNSqoAxDb4+gwc8c14ToBOlX
k/uuu0b2b5ech0lNNcMntRoKuqX0Z0SzaNkIrmELr5x5vDaeBcpa4aHuj1LBxpc7
UmNFJ9aRopSOoHlRXCQrDeqEsaD5dc2Qruf6V72lo8wCt5a7RUCcq04seE+81jg2
5rUQ7D4GC/DabNnwAoMXNXDGNJJ+Lhgbc20JFyTwNSIpbqiNkxN6hAl0i1LvyhAl
UXYtBWJyc1XrBZtcO+TnoPCr36+WMaLXTTC4ICzE60Ed3ea5oxyz4PD5RgMWA2ok
K24bMkdK1rIy1FhwbSr2hdUAHgS3Ycp536Jw2yqzz22oN937yMKHUiJigurbdf8i
bSJbaLSh9G8/+aE64VV/sXwpsYWBaIbw8z+Qlsd13bbm8qSotHlo2kI/pAv7FoC/
i4m04co4yCXLqvD2aKhrSmeZctPbv8Dib/lE1Cs+cbf/UFUdL7HSeEM+//wmQ0Tm
QJ2oEfdsTEbSHh22ZFL4kCAGYKb5bvttt5h3tT8Sv20QvIbyNlz1FOgKC79FUrZ5
+UN9u/wPvF8N6h+KuV4NtIFsu7PQjOfQ5Fnc/KthuH5PRO4ro26DUW4ypBDnOEKy
oymqyElNSHvv4X8i5yINsfV7cwCvgdR26KbgzONt3E4sCDUIZxApPr2DoEusg0S/
u10CVirVEydl5BYaBHv7j+YM86juhnKjykCFiiPTORdBVVTKr345Kn1u1NbQz+t8
xGtP+jgIH4BtUpSNKiRDTPsGGkDSbRoNrqwJYx5n1Oa26T9Wr1oIa70MhlyqAEwm
1iUmpusqIAvTRJnwJmkqfUpioPrcnpR9hK5kkxVTnPySGfl7bHo7WPWSA/dV7vG0
huy1TwkDeQGET1A9FXOdPmEPYOMy4DppWws83baSB8vnnIZ6wmC5JaGNCtRK2MNs
YkKqBdA+r6FnP0KmHPFr+dmUgN6f6biy5PJY/gjgZqrk3N5MffrUwgWGZWLtIwi5
8UFLJNaz0LskGnkVspDsgbBgb/j+kzHRUakwY/fJnYIBsjQdnIVsmnKB7G2RZgid
133MXwW7r7vBp9ET2fqK1E5489XbgremuNY25zQTTt+8DLAY2C2FW2KgFA3MWzCX
6Td2BshiU6OX/FA4CcKWWjHxO/gNwk+df4josqnpPN3llQqxTEWRAN9Fs/UxL8eY
CsqVWIKhflmFdf2PElm0OR8BTDlH60hn2c9vpj1l+DRE2Dxqiw/K5uM1HuHMXTyL
L8A+2/5dRtQuGBkv7O3VVsEoIB5HxtlQZAVmXyT+lS6Y8B2N3wr5k1nicjOXzn/T
BGkl89h9z8TYnPBCoCPWD/AujOAzfYoq4s9kq2SxctjtrrorXiwwY/LdHe3xHMHr
cPI5+cbsyi4d3wQVjhCFH6Tw5qv+G7016kfIBSghLgfmXYdUsbykcMUFygDjFKXC
C+7avMZNRW4hblk3P1qnMrBmWLgvB0wOLUoy6lXp/KEsdlpG3QanOvYFhsFD8drR
QJ/EcQQp2JAX+heyYEvBUKezJUVg85/aJF0eArIA0g7QNOyjeWGlDZz+OdxYy48L
FyXo0w9jAlRmz4T0O/ZiSTekPiZMAPDzjMuuFrnNVmIUZsbDnmImCERbBxY8nwcL
Gi4WAxs3MROUCeJ++fDkmbOy2T159+Q/vAb0ElzdGqEULYSGpO248r1lbQou+JwG
uq5q/RMtlxk/Q71O4XEAyVxWRzYMZ2Uj1fmAdLqX+CJMK65tH4jvgmkStKLW50FX
w4PZ5o6DLHTb8NPwBFWQxdtwXrCKyQBX+QP9ZOlrACHShi3HtqnR4DUIbYKx7QV2
NYukbyAbDLSjxOMaJD2DBHSCnX5gdMPjko+0APiEMUvjq6NYfOBp8v3eQOzOOO10
BypYbRpud93X8+wsD29pUvK4Fku0C3hEPHd3sFIzsj95NEwEQaomO9J6hzzOT1fb
5WxGA09oAfI4pxpoaPRE7ykmhV21ZzAubzP5k8zZTXgYTYk9+2OGakMDlPXrBP0L
NiC38oSRmwTdUKCm02DrXxvhO1EDU1sc+S4eQHQOFBXQ2y8wFtYASqpNiwgcVxFm
ggFjC5xUQD9jk0/z4s64t0lOhtOeeP4yBeSZCjsJXr0VSnIbIMTaH86kwFbQye3q
U1/QgUaeFgiTL9wag+XjSUpTxSbUbkpWxWC4LcEJzlXnUxybY8lWUuiF5aOdTIxo
HfgphLM9Qf7NmrzdWflzH9fRLjgPUxXq1QKvoQ5dCv7w+7KQPswDxO08UdCWy/6y
Z+0Xn3YddFM1lyYBqjupZ3tt978PA06S67o2SzyfXRkIZYVpXQz0M0LDNaWE7SKm
PiAPMg4IzwS3v0KSmDAzNzAaf9k0JYvIwjjzajEoHEgJnFSqE/ekDg3z4ElWv6o7
bYK8+aavbt/byR9zEgnE5WkzIv12OVdEDc1mKstg2WDg4NDM0pBvQ/wK2hIuYa16
J965Qg+PiK4Bo47xzx31iFghcmnsupziuEqb9AwRBkobuhXA8UrKLgGZ5H7HEHYa
OKjMTAgcF2Spt0KdqS8rRC6NpP1J+8qltLu+QjZR/2/kMk+Z46lmK3LaC2zv6LLU
phwThytbHL+U4v7yqqznLZ5PuUYOuLC6F+7sPTwUXKUJxd+5HzbAGs4nPngQ72vS
/xnkpLWsq3IJuVCvtoWJ9VHMDOgjbZ95tY8c5KfbI+TgshgdDCNNYoFeQxjVsKva
CLWYwlv8JKSVaXv4t9v//KxC9LoLc4I/X1+Za6gRKANbll25px+e+XqbaU0KuE02
fxJWVPd6P7B/NQfTdOxpWR4nPrdAIJOCYVKedz8YggcrrkRdM/B9EQSc2zP0wf1N
uK5/m/pOCUtkIU/iAV5pw/8TlrMovjj0Qwg/uuMbOku+vEXypT9lTcO8sUANX8H/
w/ciZCQOe4Qc8R4iolxBMdjPZZW20zPg5SwIZDYLQpkN2eZRnXD+8WEgC9CiVeCz
tK8tlUjdnHnIg+Hlop6TzAMpfygnEQl4GFHNuDeDJahoWchSA+TUZsr9b0dpjNsk
Jtla9ixMt8BtaVFFbb4GYZQbGCYKhMUjnhIfg46lIT1tVQzv278RAMRFUnCTrVb9
ATjHdxGtB5MUEGNxKDSpiaQggF7j64Ct7T1ekXhQcvXlMeMT2Gfp8W31Sz3b4nmr
fhQDIYC2QxdkIf9R6sLWVVWlIPu/u8fAhi+3bE5F8xXSqmCYLSCLaifJDVOUIFfA
oZpLMNP203KWq/EHBXxOrZM8tmHdKaZSZVyzmd7HRnzo8i5+dCPjVd1QdpSE+jQh
d8s4Vg8OKBkx1O7AfzidlYt8gTUMhFlJWmvByto3DgxR+GW56GmexzSVM3pauQpH
F6gUDRcbPy4irIlwAmpil/IJjjfrfYzgIahLegxVz9rL0JG7vEcJeaMYbbCDIvkT
Ql5EaU/OPXhW/eZcXuqdCUzxS7TVdg41MSIMOJ8HimnGBvsCfx+/R3jnOCNTgxYN
+wYwI6i2b/x3wPB4ufBuL1qdAS/hh1Ci1/rkUrRPVdkTQtdWSIzII37rJctO6vOF
ARoVqESBaSnDDae1fMALC/XXCqN6JNlKht+OUd41A1j4U3g4YzUBnqzrG4Sx1vUP
I7crvJU/QkIsPkwdLWlWp85GVQoL54Km28iI8XlYoH3a3cRZvvmHOrrWiNlLY1dr
kRg5mg8YPBqn4IM98WsvMXAj3GcDsoT1bh01SeH89diScWenZ31hZRDhqWuzDv9m
QcsBRUFmGImVWkO1TCJEsP8f6RRPMYAbf8R/zHKUejk9lMa4xSmqO5mtFMx2Bd2x
9ZJvWs3ydk6y5c0AteS+BrUg4IK9d1Kk6PW/hijGHGjECM3FZDAfmnOz2WiBemit
2YqOSRBAfgiID+VBFXXyMilKmSMhczpssOudt4gKGFfK6peNeZg4hTq79ml8ngEf
MkM/pSr41h0OiqmKPQ//Fgq/inq6wsUYbLg99eFAohRoerSBGbp7KSFJlVJ7E+ZE
w1DnB8+N0F9rAIWS0EWvnsWmP4UrTA1hV0JyABW7Zk5NAxib+BxRtW3ggs9aG86W
QJ1y9zaL1ehXZvQLgL7pIIWoHFY1tTttMvUj6wDVWERL03znzNT5cL6rxfZePctF
yiUqOaasljlOIkAcHuU9KLwn5FSZseFMjwbyNHjOLsc3emEOw6uxoGKDNIggCul+
Cnv+H1ALZWd1Ew0UF8Mm8a7BdL3zPEpOpYV3WnZycx24X6SFXLox2i6i6TSXuwzF
HVfLq/fGR6J5UrWNgiEp8O3H1AoqJypgR91/dF6xb+eFB1fuctkOwUauEfvSlOAS
ri/vBSwRuFfUGQhm88oJt1+nQGISQU83oPuLLx/tqNjsGdhQSdPaXxQ9CJh5zuia
0+OHN293zYz+iBKkpYejSMnopiqahvHo0OJV81AVf3zS8GO1dgMzv8ExV78seew8
Cf+9g/L4NSynSVlNd/Sp77iBSy9wf5SnFYiy1ESPJQefQBsnszAL6pjJ+WcY6xkt
h96C5OZ1dzIwYG0aMyi7CivCAxegAj1brQUv7eDjTNTh0yaxYdgov1sIK0tn7elL
poH745TctRlh/QKu7tMh0DVBuKda8kp89E6biiCHjdVbQ8Mv95UmViGv7UqbfdKq
iKOCju4ng4HzYBj07VuErTi/QNSOkxbeleABlKX40Zcj1vzQ/KcL6O/yi4381Sbf
/U361KasYGLykvY/dlVr/UjarzM49I1LgTvN8/049s6ABcXotD8PSBnp4GlmWhXu
UrwGYtslvHYA10kgg+FaOo9U+i4VQD9gAqWpzZL8fNzCf1azsg7o90MtmOTraZqm
iVN9DSygEJjXgNcZ3MulK6NLCY7iK1WihkWf/+p+7G/K5OrzXuhifXpczgja2Nar
IGrvj3BWJ/V4UaYzr11hx4gsycbcH4mB1FnFSki7iTlykP3Bh5nRHP86iX07DMyv
P9NYqzQ5qJEc7vKpjqKrNajo5c6p9DJ5RY4+yg2EF0qYs66IWz3vaFCL4sGHiXuD
NH8tLo8uN6A9jbIf2XXVGgFjqfrFyzrjck2YdMHD6nGhrIN8WSqjJfDUMLBjXxvW
vv7EGuIN1fHhd8PSRRWrEu6n0ArFUyNyWuofpbQMYX0TyqA4hac9zNKYyuirSAxK
GN5SC/mPVzc+vQmw1lDM70dbOKkKhtcxvHly2ITs9e0lE6hw95sp0mqkTEJ9EkSz
bPuJ9fwRsYv3bWJf8HJczvPXXk/ZKIA+E/1t8iwqo19UJKd6ZIqH/nWVX6e8Fsp1
CfYE+9fbQEn4t4W/TQqTZCbpVbGZLz0r8pVE17Wj6cFXwnhklnRPKOiLqDxIRmAZ
GbYqU708pX+5NECdVTHdLSzIZ3K0IWtVmsmN6U/UM51XARfrgMeY2rBgsen2iUOV
/xzba2SC81aIFPd7jZM63WkHU2AcRKt0dafbAvL0ZwQdAtt49bS29SRlWy0tE2wy
Z3ckMcb7/+maHepRKuYdFa/LAPMmiGorUdgRbSJAzfYwb1dEec947Bu7i3qgyBnW
31BaBU9O+h2WFl2XaDXsU+iZeT9yMe1180pIKZQbXXXuzGrBGikGV/L2lhf4EXn8
JkwYBgSfq7rUKA0wFCf5J5P9s69AYKYV5NrUzjIv0XmWpbitojNxmu07IyhGYc2O
YbVDI7CxsVLHNvhwcKftkJe1lXtPVMYPo46eOkKzJR/4tfj9QxJ3gelvB1Z2KDrR
9slBT2JvNgZmcW82Rn1lzx8yO+1bwEyIX9IUgINm7prL/YlmK44/nYuc0LrN1Nb9
AO/pbkgbgv/iSRL9wWR3Or1WwQ4qBfC6CYokRl3ZCQdn6V8Cm7I/9xpNjlLdkRtR
wUbzVXNsnFdAVzIU5Xy7/76nofwNjnVfNgmF3zcQOfyGdgaamiP6QO5W/JYCmGQI
kqKuuh8qTqbZXLrRRyt2ahUfNAMOSUmuECtPQMQ/u4NBkw+L/+cG/VpzcZax3/Rw
b8qHoXEK/w4hwpftmr+1ZcRsFqRXe7uuKLcXBxnDYxSTJPCyPNRl8lDuzuX5qZzv
XrOZY4gC4Ga+8+fvewmNR/cOCFQCNSmUcYqE4XDCb3IL82tWVu6U7sWfYcjH5V69
w8MxMgX4QYMeSJk00D855BEbhKMYkbAMCADZv39mjcNlZKPYekEaCn6/UCB4xRJu
a9loFEN+FPEjQjd+q0XRe4PnugFsuFsQFoUtDYaUewoHwpTZDi6oa43o8obCgm6Z
rdTLFx2JxKvxhKG+wUpRLAzERt8kjO54wIKJy6pq7GJllIE94do/XEzRpihKeF1j
KQSOYA/BG8RDkYPJR2wuYVLkeKkVbPKl7Ft+J5OMas5YNJoeM8JlpZi6p7xf+TdH
tK24nG7WUrN0HRPkrmeH3vTEKRb7xxtAkz85cRKuToWaH0GIARVPS/PbOtbmteKs
QhsLlya7VoP3RM6yc2Qt2LivDMnHkYKIUY+aZ541QN5vI64fc32jRRf3R+wRzpvT
fAIM75E262dK6hOWIrUpDBdnSICWstMajvTuxGTHNE5GYWzQ/apWrkxo2jBcisy0
3a0RpOs4JMp+Am7RC5fCieto0PDNpct4Cj7lGKVKsxPfr7Wts0vT7VzwgOGd+GLT
lXostajFgsoFez4/ttgowg5Mk30/fy3I1X5hnM2pwqnlWFR2sKRA/POlPrjZFOwN
xCgOEw1aBzMx217dWQ6AASfIhYaVtZ25+XUuyaR18GWUVt17ZOf/yRmaeS3iOMyi
26lrX/zl+9FZK/+te/tavjb62EQMej5XDjzujgSn27AQ6mmjJqatFt0PlvG2v2zr
Q9cdBysREA+rmDtQpqlPzO2FvzKg4UcV0FPi772QbWvCaui7B34dD47tfti3yZVg
qf/K/lO9nN1DFoMnd1jsPiGo08AjaBzbV0lNKPJL753BQm+LgzI2vnL8W7cbZe1S
2tJiLHmVDNi1vSPkDFOVcTApYJtW5l5kZiYdQTuC3bmCIzdeQyzkZRkxj5vGZEXt
2Nmb7oC2PMyOm7SNboBBXcZQLWPX5rRq2HTJGfxqhAxfHpVEkP3Lp1vSN+pBBfqL
nfjERcvrkMSs4/xMSTJnlGSfMKaJmIbsnRo+4ORHopSvEp6aCWGDQIDdvQR8W8mr
ezWVLfgDzwpXrxylWfJToqVEgL0+UYjJPGxbr0GWUxzzjpgvADL5IAWu+ozT1muW
UdxMQmb78zsCrfbWhrxqxnC7H53j/BQDniNnhwV8IzmVizf3YgdHF5cO9+6TvluU
+4twEaUqkpxuvwHuo+SSHOud4wbnrRULtKTbSju7o/CBoDKJEmV2FiOYoDOwuHZG
MNlLrIR3P6OTcA45GWM6tuXvaclVpXrE2Ge/I3/XL/NvHEu43ufdwcWYtFMtMRzO
+V2mlGG4tY7xayDhqlMH72wbBrJPgtU2Ln7ridz0IY5AnqkK8hbnYSBBIhpLqDgm
ZPoDarXZfIiak31oBb9+YQQdogEH9PdCccSyd3u0oXWmzmZFNZMoAwlqFhJYlNcK
rz0lxZraSZMk8ONxnf7Wi7Ek3+glDYkDU63yvpfsbyXCL2l2/Yv2ky2y0d/Jyvpi
aemEnYgFuVGC+N6yd1FfDHCkjoV1u0TmVxSgj0BexrQNpY8oGser05imnsqdWRyr
UmBF1tyhcOMLCBsGui7pdez3WvALhjH9EpCZ+Tgd8uembVJJhNupPnmedJ9Q+f14
wG31cGTA6MehoWiKwwE9iRlv+vJArXxlSwBRUhqQbaf1645sGqPKwVw7ZxZpPxzO
u0jJ/6HqfgaXRvYTf2O499ct7nmkraV1mJmbY1FDzLCFGEqxIdsc8DdjGwqWgE/P
RXGH8xmolLD/F6TmDTOZBCALAK9rl2KXuQbNRC4pPqk/LeBObKdJqBcmM4Ta/PQS
7RbQVatOOniMH2heXTcuHt3i7Pvu+8JbDLqiLFhEJ/ROe32pAEVh7GwR897kktWl
J+PMXKCfoJInW4Qd+sfH6J6l9ZYErwnxV0xmrOzX++6KUYHHF76aYIPnJ0w4rT5D
aLy6szkhcy/kTj7U3kbzGfak9LWmwL9Ppqqi31wwxNy6+b0sD/3TuPfuMElG34lP
XPU4WUqj4iNqQ8/3zH91om3A1CN5ad0+D//jbnbs1CM3hB2aiqiPz/VB4+1XwkxR
YlRkVeKFJhy4vLK2PJ/RKBVXnptEfnWrWaZHodAvqP2WCdSlyfPSggDKARbVO4ap
dItC5toAT1JM6WkWauDFRhCo7QkSkdrhXN3Sw67HCm8Q9F6LA25lJrTjoF2udUHI
pj9GjGeW9rmCUKzq6eDd7fbCqC96tE18F5CxrrjDRz9U5Jos0Le3p6SnTTFScswi
edWd5bUKjpiZQEkxuQlbkAJBCcb4BfDDs+TBRgCzIrEGi8FnexTdZhZVRSaLw4TX
PLae8AMwmoogmoq1JDvg9KoKnr8dkZZfrM22YzCIa34pRRZ8/NmhgL9ORUVTWXK3
G40kVKgoZm+4tMKLq4S86fHgt1mPokQJjlw52gR9AyA1WLM8Mv6dGhiHXZ7uKWEI
m+hZ9c+KIOl3OX6J+sX0S9dsihuDjm/JKDeqCpKyEPrJ3J06/3du4GUgu0hNtujr
d9QALGNrwUOgrbAEVj7Z0UkM1yRn/aMUNlZz49gkyyv+avoBL9Jcd/LKE+PQpnGx
MZc2VBxbgfiTXbq9B34y/K5JELezt7gRhfB26io1GQQb2I/jzT3K65u++8n68u8L
vmL2PIU9n1PeCjrfmlFeBozRtVtyBH3RNQWUwsOiq4+xxr61z8K+cyGsn+1xYviM
1kDoUUbJdLZ3HTDy6XUSTwecyXb35dPQ1vGq4i8XRmIOI/ey5fAG6bx+5C1nlS+T
mNNx9e4ZZjUgmGGEljCBLpG+0m9rlR8GX16rQ+dksn+YLx+dUm7IY5YcGbaQy9hy
iWOnDv2LsHNBFvfSEoGMYuXI+SMWurqlH/SGQh+PgsZrrUN9aGFYyMJ37Vow/jqC
sMZ4g2PEm027KrEjJRz5aiDI78D4/JvDgr42Yct5WLbljuev5TMkcZDhUX3j4mNf
O4p1Rkr4e/Y3j5huRW8GXn6Q9J3D+pmxrDpyILpr3AXUjCyA1Jq1OHX/vKu1f5wP
RFihzEEm0LtYDh2SGyYGU/bVBbsCGE0tvWhszPLlaS7E6MIqtroHwxlwOCYuLF0B
indFJEMGJ/68suqwVlmIFL9dJeJu6JDEdq3dSYJI87Laj3QJlRAz4bH5StHWmwC0
0bHcWeZnVyZm1M4MrR1FjgEig+vlAQ8psDOpmSdAyb1Rjcp/7tLxe6vnckRsYa3/
yRwk79qr3b/lr0S3ix+Rfi873gThQQZKnNoi2zjJ1CVbG6W9GKO174vXiO4vK50G
ZCTTw8pJgmF0/A7dwnz7TTFwe+eglJTvFjJSJ184/D8had0KI7Qci6I9JkbSCBzD
EWu1xgOkH/ad38XkKD2U6ngTu6k9YzhaYpoG46k68Xy68HuLH2wLZA3YY7h9BckA
MPh1/LD8xawqC+LTaRBoiOjAl85us/diqIMfZ4L85FKdyX6CBEXFNYA1OQEY+AXO
rIQz7J9JQti7yFP2hhap+JV33Buug/tHrN9TNqI9wRbOyxUEZEdtYYzPe3owP2UY
8JHGoL3DfCVkzLMnlrdu3Fz49fOW3lmTzABSQubiFeUcd93aEhDkA5MuNYII4mfd
0pcDa6YKD+YPAfxmR2ZHGWh1yZCxQjRig5woUO+PpxjCHFTMTtOIJzjy6u1r4ZWn
Xc9CKRYG8VbgR0O9YoDQ70Z9RVWC/9vRCthfWQTMcHVrE7CG1xWNAC0kJXEbKI++
Y3SoOhsQu3tVQL03fhlPwS78ivWZpo+7eMs9qBcOwGLy7R6WvzgcFYT3NdEA4INO
QiXIXGFkVWiBjcox3I2nz8/InusCR0/4ougUHP++x7JkO0ZLc1GQnA7ZFI2tC1vh
+y8Z3jpKyryQ0n7uMfXq0L7xuXXF0wQpW1//+bMPHSDULEHEp8KYIZ92iHINPoDG
uudJ3ZsQp3YCLrEJBMmU5EbNBjR4V/oWHIS73Yy+4c3MffOlnPLLASV+Q0+ZJ3To
ht9aYOf6ltfTrJty6bqej5ULmWLJxQptLamoakhEZz3+q7jOW/uOw3kf2GlRT9sT
vwiBeyQO2j3AuVb4y6FS+1lnq/CBBPAhK9YQR3Cv6UAQ0Ysb80JPd1gMWeo/6thT
d059MGYQZgcUaZ2EH1H1JlF+ELUnZ8ic+5WGjm2UWJuhd6MC17ZtFwRDlJA112zq
cZ1dDymtXR3vH8WuWBF9rgVjjvgD7sXmAqut9iSDrIQrRmILrlK82ncFYz86bMeq
YowYYeqXA1v4sTIOQyxSvTfxrehvwX+IIKV/41238ifvI5OJEZz7cLShEk0L9CWQ
lYjjN7rtW87sl11xUKxfOgj1C9OnyGeDOBgMs5KqIvQxkG4rgemOulW2odXdrOXo
T26xcaAdBNZt4Jrd5dKK/PL9aRv0WDqiid0lf6J0n8bleL+6Db7+ZpocQgWmAtyS
DDv31MPinw/ZMipmFbkjf2qNOITPTnR9NH8fWLwUZVK1zZFZKWyokECLWGzJdudl
bH6Rbu2wUD9FOiEWEVG8Qajl/SeWVOQfVyoVZSId526zy9GEw5Q6rmxwj6mO6h9g
PJ0FeDa/GaDAXlZB86+pmSN61jbIRoTjhjhcK6pdHlWk4CzP/67b1oNH/P/cZ6fF
7GLQUhCuppCgw+3leA6xxhxEdr8jsokTJZ8n+rfQ6PXKv3AcA9rTg0WKaJXNZ9UG
uwZJpy+/nTNqITS+tGg2Ycqi3Orqb71g2OyLx4YphK0BX+0KUcw1i4eDrLnyPVR5
07qdea596fyrCchMvHmAjwPCio0HBFOQSdUEqh6hCEZyx+WP6+urmPB0HdU9ecno
HKDn6YW/F00OaGn1Dpwo73FTLZ6B9WHUotIQOvh54LTAKdltq0yhlVIoTS/GE/2z
CJIzX0dlV8BxNU9HjDLODHIDcKC90Uxn25JrxhHWrOXQkWgRqVl86VIX6WOEFMep
8LzgM/bmFkWg67E0oxz2YEBnoOh69vG9T8ejOHT3gQH/maljZmg+D8dREf3sP11e
tM7VtsMPKbGdDf9kVDI5yBXugAAf8FaN4uEFcku3IKuC2YQsXUEX9HK/qf9VUKUx
ZDYKzxlgoC5wfjUoDJXoy22vKfsDyGY/l3fedaMyM8+fOThH/ofompiwL2eRJEZZ
lt4+y73wMEFR6PGGxuMCzQ/Dt/A95ZE7MXNpID3jaOUs0QFU7yxIScWRGbfHz1J5
5A2z3nVgpWcKGbgxVwGbVS/SmnudJFVhEhcun8l7W2OHJ+e8Ep2X7Yj0sNkrGorj
1cLFudTJytodLIv9py09KclnZJuk9uhq4NSpwf9q9jzscRYn1xf7rK4tZGXMagy4
ZhhwxTbR9uqYfOA3+/1migKcxytinPaXWFsbqO1iN6NbVyr98SOpY0BrHqJNEdoP
XgNzf3f0e/pCTtEaRo3HcDBhB3ao3xQoGZdIhVjtkHBvwGplXpk52Y8/kZJZDYdA
YiLGb4abc4HuCQSGkTBz9J7TDSIoDRiEasLFXwPhFEWJm70sYzIDGzEemAAlMARv
orK9c8y8GFnvPsbGvpXnO8UsMBbKVwHmzjOEw5sx3mvxnxV0ZMIFoSZZQ3Ql2Yed
+ymxiY1pvaPXuHtqYHWexPdcryuJETyXVkcWHyVgR5KB2bgMUuAentXIEHg5j4j3
jgnzwLzAKZMg2kfHoCyQP9I/YRQ5ECn0WtBMDcCmVaEqzfmTYq6FXrprCtFh8q0M
xkEstaRvWQHsUBnh4AkGCtXyTnkEiYPOLsleavX/EzOlQjDuldErwUBGamZbnm23
FPnQXPr4Z7i2/nALXqxEKwdYBymvTC2yTGkxKOuRJb4SQ1eEx54T2t47GaN76UxX
pV8riQwkla+kNjfvZKOCLL8OtbjOJzf14yZDXznQ7ldjxGLAPf2t7ZS4d4fVZEE9
U1wnWE1FOKQRRj1/XUF8+dvZv7yMKJcnHuA5P64k67C1fyP1gM4GRUuAajESh9yo
ynVeBz0HqRhZepNgOYjsmLoebIRGU7rbn7iX7FqKayFxeH55J4vfs4QXGahA75Pv
xFPxcPP3SrMa18P01Wim+owJHPQ4EXF9buIjZG523M3DnxzZJ3/yQ82sIGjlYsI1
SCUBJJDDWZgvCF97F3Gr1IUp+qTaVbiAuiLd1riPZiOC6o+b5MZW90Ibey8Ora1L
ZbmC3r0ImLrOIIpH8zvH7LHB8MCD6I2/582l5bL8qh55hwOVCIyl9PaxU3X8mwAq
loOZu405RhChldAriR5WnkdN55YiauGxfZLtgJP1R5u/qqCSIqDh1C6CyP8RhPEo
9iqC4cS2Rl4K7UHiHc3h5fHgiEiwdOPqaWzkdUyojGv9v4u3H+2PA+M+xw5FqnA4
hr32UKL6tBXKBCaY1dMMOB4ZJOwsuUDY5Lv5rVrH2GDs8kWOIBLBkTki3xFv3TB5
q2SWUSwKd0yl2/BGd+g9tFY+THgeYYK0Te2dBVCmPeLoVc1cmgBuZVbINfjuIOef
J/+0q7BXb2YcLc0/amF5QmWnFz7t8zE//bA9ab/ql/y2Yrx1hKzpUrLxdlYiTkEP
LKjEoQl1dSS6eijzX6Y3AM7/WjsJuYkLPuW7963G08bxJ+7T3kzlFmK+m9adLsAM
oHFvh4KYHX+rjbqAvRsGUsSU+V91Dq5onRmRZeWpDAfZqNpxv5N1jEA3P4JAWbld
S98w2nQToT3qh5Hn8EivhBrXxTIMsAWsLxMQ7oFoK3yFMxzEjKog2197Wp/fzF03
1dKBxQQ8/2bUPahoU7h62kq/0bvPntX9heP2+2heAS1E9h4uXSiR8H3Pa45KJ9am
WSnmkr/H89qGKjljx5xXQylVgruMmv1gaea2ec5YuErGAHuUuaOs/ShZjdte6j+G
afdAcYSe29edG+0iq/44FFbGpAuxZ6Cc2SU+Fy9KWEZFG6p1s3RN/l5Ie1ctv3OF
NMCjZ+PqkQg/NboJKbSQQ48MRJBJiT0JI73rnvzCtmU43Q2Ey8pzGEmVgcbkBq+A
nbEqkrpV7bSipyJFbg3aX9MO4tGyvNpTS++CNid+s/Kw6eCxKaQgFKdauY26wJkL
7bQHxE3skkcb+c990kT7iAUgMBWOSCRFOObKwnsf5ifZzhww+ir2rnyRuMMDMxH3
XpAko0sCwuCfxic5ysBCke6wyJKGqAWf/lAB70mB0ysL5QlAKjpmBNHPPZ9wbnhw
1bXAh7UndKYFvZvETWdrm0J1zjbAb6/UknJ/9oCEKBsNuoJ5AJBrXHGXtPEPYYGz
LM5fKrXrB5eX4SFxmrTfZ8EeilNe2JRp4zQl6jYcHbtQ76h63AcXgcBOfHw6di3L
OJrC8MFEoUSM5o+wLzSMZurv66GwOrJyGPKO7z9jfeXqIEsAZanLEluVdX+JwZnj
RoNZa2a5tRXXoAtbvHsJYL7KEKOR7BKV5cN+robrNWfZGsyhnb2PHk9Yp3Dnaxd/
o4/ZyYF06TuGobtlDLuncnlkxox7l9gOUcaSwejCC0NKP2ZLZnw+kdyRSvvKezXx
WbU9in6a+k+pU6aEs9qxrA3yMEGsPp3nmopBkcdxCSN43q3Owoc0L50pZIESR9mg
telv80nU82ezpHMN9QLHXjRCZZ/rTHHcMYP1GtVzqlGWVbC1l5U066ZVnFF66pAm
3LJkwIg7E0p8igvjfSed8Sq66+nIcejOf19ckJYBE6kxly8PVW0oV2uVHrONe0Tl
dE6hd/IMgJgDpVd49SLybojblsY1DyBiQQ+jrxfxTZ6lVaiYFAzn1XfheuR8u3tx
YpbNGb7qet0U9j1lqdwKtmD2bFRojkpjfcDcT4JqqD3YhUp8D11/RjLaayUNvhOB
g47qHhcDOF34x/wMntpXJJNxf1uR/GVkOhjeGVoK6pjsaN9h2c9E09YoReeveQgO
xEKazvZcJfEW+fQA9OWYT1GEh5yE/dicxyfAkM0p5Bk8PZd6BCGFx6b1R8UcEFAO
NBqSUr130N6etbF3a2P/+a69fXV00404Zb6cz/S1AWiiRVfzWJJOTLlxUqR5/c6k
laQUks7XdCyjxvG84ZzlnM0femLWf7zgloV/B+n4VYer3YXcn7MWQ87DY++yPKOa
ikD1mszg+bmqYM+mwPRf3MaTVwcwssUu5prEhP60ZaPxk65AZAz90jv+SA/pkjv7
au+mO0GFV57DysgnnODMej2L8/qBjnTKZ9Kmm1/L9j3ZClR/RTxdUYp8SFJ5tWOB
NZb957nU2olzU413lZWR3VGCn4+GOLmwRuDBwuG+z+hTQbjU2er/pP3S9a+0Rn6e
A1nonmlEl2r9m2hD2inn9Ld/gpt2Ze0EOJVg+3ATM68Ge+POkO7LO76Bd58FdZUd
t8Gva9pa9aPNKtcU+5epFezrtx8+7tXhFbG5/yIH0OI5vckzlyxv6L+2Z6Hmb6St
9pNyR2P+AYP/x18v8iaG1k3M9UZv02oFD7rYbdeYCBcn2zMctILHPMEODD22dTZa
L0H1uqyVupBA1WOHUqBy8MsDUneGP43zyrbdmLdMoQNZB+3ygwaxQelA/dym9BX3
XCbkNA4m9HTHzyQg/Lvoy0pVuBeGcg15PEwMYyC2sj2uf4t6LE0Y3YTmHYC4egH1
tqbkpNbcZIN+JBfB2qWdXEZMMNoGKpZVy2jBM64TmDq/bkf0ZDcXdKVW9us+rj7P
5duj1aEI7Vke15ZT95GpVL/cLPxoQ5srHh2L2Yu7ociFiO0jZlFY+72P1lxcOZqg
Ool6NByodP0qO3p2j/ic4NYl/VRi6KaNMsaV97r4MG1svU9zV6kn2+JI9IMdNvut
HTAN10OdAKNN4lZsx25ahXTroBenXJaq+0uA3pXUL2pHwxzRT5ih/dV40r1ZoX5H
UV/mwWpapMMsWVwh20Kpff/6bhBfPttvD2l1qZ2bYaFjynr1COaXUQ2K3M5CalsX
c+UhGtPCwx4uxQktdqj6ruULXDe5isE+/cIguY2N8VdgOX4eDulO4tmbc8Zdzyry
gWI8dAobb/SzEBHzx9cHOODvgy4wSHwbWP1P+o/pX/tEfnjyjWg/tNixg9YSdOwG
Fqf1abH4t/LxU1yEChxrSMmwzFsXzEcvMqCC6NQBH7oSWJz0r/auTPa9HWVlvba0
mAlWeWokfm0o11yMeh+RwjUKqNtnNmkZd3+MzlITkalfZ7iQuKYE68XjhS6ZMbW+
5mQaJ5vs8nh88BrZQbInIAsxwFydTxbZnYO4h0adry1pHVnOade1JCvehBOAs7Qy
bvoBWfh0z/E4gxPpRphG3fq36zGLCv3m80yLhP4A1ZelFuOVza/QKP33K+AW34FH
zzq/suuKFg4B0d0XxGm3Or48UtljTcpmZ/7tKApmqez6c2vIbOnEE2cSnj/IlfeH
qGD8OIc3i3muLy2sbm8bJGHXwyx+coxlvkmM7cK62wKbRFz6NkDkSUJJHrkgIn4a
QFpAWeXAKTOWgU542YnnKNygTSNG+ja88DNu77f3xG5pygYqvxstC1LMTBL4tvyv
MFrYEX2sgGaxEGo7ouDg7O4kxiwMQrWeDWoIdhHlDQH5cCqgyh3OnEusExx5LaZO
wnfZZ4svgs5kbKEoOVrYpOlX6LtQCcvO4JDcTv5ycBTuprKaL0HcbIQIVUIYfITs
rztL4PlNQPg0taA0XYIF64MTPiDmRyLJa2by1AEl6XHE9kPbwucLX7dd5so7HWaB
/zZSjFvJbf036vUpjSD6O4gOIcB+ESWkG7vtyUr90WMCzJ/gxvejTxqMUbDixsIZ
vsb24rkLmHzB4Pyldaw7vRCxujL/MUZjmnWcBX9XdnQ55zbx0RxpKIEVNpYcvjw3
FRqqoKJZrez10b0mdAA+v220k93mPEzG8UAdjf3HPYsvun0xT3uI4IjjyYtwztTG
CUlNSjeyv0IQa7xK7g+deprxTCVa1JXBgTndG8LSMSHGvj+mNCbwQSxK0HCLn9vY
l0ttWESUGsyxFHJp47U0OBWKd9S/EtZA8vz0D3YvigznAKhJg5xQfpPlJWc8U5hp
QRnJyXkNS04MeCwUHmxL3hidcbXjvR6kS2jqEl/j4tJCx/FpYovfgTsXEW1H5rIH
m/FoEOB+/qiOXmZji+iRwZTVWOcSDEpLqpARRPLPcIYK+GqW9rxEQSa9Q8MG0Oko
rw3fZnwq9msE3q6CxRLesiWfTuBwQW2bdQXc6PVMdQbibQlK6T/gLWtY9g+yr/oo
ybr8hZ7dTge0GluDgqlIodvVg8v2JRilFw9IawYCMUFm1Mz3ckr4e2UGe1G/Sion
krlbe/+Bjf1U73PY8Q4sPOTuG755WascXUTt+QFha9jM1OvV3B6tLuJNEdjbnOWE
s9GRsdY2aQXcAWi02T14sH263yl+SALjuVuyqqCk1yWb41GXHyWQDHI9bWa3c0/T
Toj2KcI/vMxCLGYV20U4Zbl/SEtKt/k1ooJ0UrQm7YSQDLEll3LRgPSqqlVfxGrc
MMNFoeEk/1F4uNYwm4/LOIJxNeiHYFFxcVOvaVCPB+R/FRbu7fZiv0yRj9vxRuWy
5nq+gaQX62vvo/g7NkgaGJ2HZvYgTA/X1zB2WfO2VPY5kASxqE0VKy7LxgdHH88P
ipw/RFNjtP03wbVoIH6VlTh3QjGu809ARvPA9YCl5Iahz8JzSYy+EwH6HuvfOEjD
3aR2XnL8dN80KvWBZ8wVvuAgcOv5ly1CqR6OlC8ZUGS9Q/MvV+6W0myKWv+R36fm
ZObWaL+W8MTxuZpH/I5Jj4Pk0K4RcdgSn0yDb35QfltOWi4otzDIw4nL0hubhOpz
SDwWCBtx5p5CeoSZceWckqpQ3fwE9ow4W5VhGZIBw9mzNTbJv9LX5OzqDzfu2s4t
J9IC0pSy0JDADHh8NBQ58yLd7/f6ZMq0LCVs+gix55+rGiFZWv4kxvm1TQxPETZH
15oFJiA8f6hFem+7+eCCMyxj9ZYocox1zNNPZzq32pSOAeAwA4oS4PSvjrRMWs4A
LaxsdaFHvnunSmgSxhRXmgga/piUmcooDwT8dyyZolB3OBMFIvZvZxmx7lwEF5BO
mRmkUg6lNLf1f9SJYkVNMzJYlnmIh485Tlryp7F8qpkwXb8J6GWllfr06VUBzqD7
IypXuMVRs+CUnYWn1GmdIHfBaI59izf3qsEl9gE/UWzxtL+7ZFPBNBFdw3WIT6Ss
YGRUtN/Qk2SfO35/nxeQDYs0QVEtdm/K33Fduq4zGjNgYYGXh5ArEKvs5n2mWjJ6
204u2QrOd4nMmDi8iEV1irh18A1APtkXCScPqdNbQ8vLy2yV0/kFbsBFcGFwU5sr
tt6gKbRlKTasKUQ2CxvXepdLiL7iWp1efnPzD8ibdGaGYRXmp90jtgQPlejkxzra
nc5W1zUKKsb5v0URG0LooYIyur1bHCMHOVVeM7MZkjb17cAFSeynhbBbfSJJlkyl
85yRKRZuZXvlTy/r7+/1bveSi6vtvXLPWZ6adBGRmM5LtA8cnQmJX4x85BFE2+Gb
T6nPBmniKyQhQ4Ep1rS6vnaYmMUKwd+b4AY1jskR0dlEeyqZAhQNZkYE+l8sOnba
oNWTq3gFFsmX844jC6Dq59PSSXPc7y41ShBhiCW+OV8E/vbw3D06/0aG/uvTgUYO
4cOHljN6sFhadSIR9buwPHGLpxQHjNMO3TRW1l0y1WSf8EIUkl2pFH9t0C4UsKgk
35AvWIfiBcE5XhkT4K2mHAJeNtofxkAEi5SGnWBXT4uBYdTHckQ2mBgFXzsusrBe
tpQ+PdPjfcWE0zx1dbWVXre6GOvtVbOH7s9kuffVZQqQfzpdRcPY8Nc+crmuZWe2
Y1Hf6lzFaDaVZAPNNV1xxOs77nq7NKpTQoi3yh/q9IEh4nzbzUlpTAxIHFfLRQrA
6LmdXS+3b5sSgofFq/tx3h6i/sRhbvbhhJnp2Gr1+rcAG097w6Gip4uO+C3ahJih
O1+ynVZJtGb+Wams3H/mG4piNcd19CY0s/LwwIZ+7uTCqqfdPPgUxHNNzkg6N3qQ
SZvzfEUdHBK5gJclKDC7Fpwu2ao4QpK40HWlKjdU3LtVGPEfOAlomzWd+MwqkZcG
+DEB8oF8KAA8KO+Vd4RaQkobvGD/2mBOlB42kZwDVkHmmeAQX2uEHydSiI0X1mcx
7EhpNuLbggiTJjk06PgQPbLcHVaFq/JSEQoJo+0t8DwOGRVPzkh28UVEJmm9IOFL
9XcSn487B9qo1/SGxll0703PPHV8dTMmoa+OsntWDp3ZM/76NT/xxlD+edswM5Xg
/fDb8pHfXzd4AIDQzsrP1u+fsYlmBZ2sWPkV6AQTA6XTli8w8Hpl9X5iKEoK9ged
CH7p+Fg5Pgc5x0JK9PGmmnznqoVYqqkVXASE8KV4FoNQ5Je6my4+FobNvDqm83To
jhfMMbja/dxUiQfAPHoj6zVQa1uSvA+jXQE32DWeklblhmZHrcP2ADsrpm2ke3VQ
CZkv1QvDMdLA6H5AuHgLJ3AWrGv8YqHItLQxqMyxojY6susvD3avxKsDUTjzfyOX
i0c8ds6iFq999Ig/Aa/CZo4XzMLs9QeRoL8v59SBbNtXyJ2JipKXaCM4EMDp7Zqb
2hDsKBYD6BJLZmxmjn7iiEMgHqMrpY43jpC1WoX47Ye5I9xdmc4T/vFKBuu3Mwta
eyxjfjp+PLVRCjTVf6B9GjLyOKJ198OwNQhqj7x5jigsDkS0hRfSxX2UzRwWWLLj
BneldXnf45nlZPHzdsXIJJTS3QUSMikyDhn5rUIohxYeD52rh8sZX3Sm4QRqGGOm
w+dncrSUBE06M9N18zOjZo3ZRekmb/KZpxs9yAjlCBc3/7wrZsfcc0RUNmSw4lJL
+VpV6QV9fsW+fYP3vgZPaoX4ChxuirBPKGCPkzOKh8A4rQmjdaUSPrJBlwh3KFLO
HQ5NMwgec4/92HyH+wn24K+KIHVZaLoGYjcSYwJOQT1NgpnnXwHIQ9NlFNcBYF4A
yDKRtbWzs3LfVSVlv6n5/Qmejn+xIEkkyhyQYFQvY6C0V5Qt+arKKCJC9ybYAlxr
dC8da9fNAewRBofALKnfj/G4siZA6C76dZ3b261MOCXug2zjj5OhtK9SojrZcUFk
0cellqGze0A3ud2h84X9mszDV8/n8pCh2MIVwuNbpoF8LjnaQ6Yfzwte7JbsWBRC
61YcvrcIRhVWT3VK7OG5kxkCSlrhzz0tD1Ob4bW1f7k+z0xitrLgvKqrXKGw6SX2
nN5JTZMQMmutTqP60x+qNxaoadPYwXr3zk5csSIU0+QlmblsS+PgxQkxI8/b019n
ebJATKtMRDXTHFeHR90yb2W+2G9rVkon9XoHb6cqRRfH9hLKcJavA1ymmQ+Lx22k
B7NnscexS5CUzlvy0teE2K+gJG66CHC0aUDfjF7HhMtLcNdH6ZIZPYJ574rljH5e
+pRS6wZ/0VNQ82nQQgcFjLqE4bPBHxo2UWQqR/VtvGJKBsBm7L5ESpJEwdDCf3gw
4RrcDr2GNEFGb+ovO3SN6waGBN/0r7oTYCN12teCL6UNRR5tROBq2CsGp/4kP91k
TY6NaS44ZUtrxpOYgU2ngXfiL8ncy2OyTIJOfIr2NpMXs9zhR5zauSpeYBjNVlTC
rSLFIT814NVq9SaYXb1XQKc8K5V+uGThYjOQcoG+6FcT/VyOiZF+rhgEzZD+ap3U
KOeWeCNr1+mTZB/KTQ+8fPQhjNP1EESRDP5MCgyrQckcK7oV+1Z6yg+5U7GCPjxH
8bA7kIwudgwnbOUIFdXGJAaDHZ2aaWOsSztLhbKYuWwLzvrur4xAMPSyaSvqXIn0
e2wp0Y+xGtReH5qZ306HJXephcBfRE1WtFy8TsfHIgdBnhYIHG2jnT9xOsJC1KlL
iEJ9ZhhJp8VzMcvSlDass68BWIafLMYcqfP6Vo0NMOoO8TyqY/CcalH9AqxBqSZ0
AXkVjb8ue07XEYmFr1xjl2fYKZ8qhCRYwDPA/Z7u1BxPtiY6gRZSMVnRk7fhyD5W
/hBgt9VjGqve2IM2DbGMGx8wmV6Bfqx4gJ8vH+8dHSQgmlpRsfjR7j5Dhpx6ayo8
JiGXA3miHPBHJU1Mc3C5nY3VyOmdyw1VNJFGADkQTjwtKZMYuepu1mRtPpSIor4G
Li5Ayegw+nV3KuwMD/qw7+ISJeuSnXi71eviwO74+YWkJ3BWi59sMfYXwbx5vONz
+LYpmnit9rj/iHLDbb6YyUvHkBP6v79xm9uPsjjyddvJoXHHic3IK21UHN9eDNYs
8KmFCImpvZg7w2/7aZE7a7J/qRBWo6UBeEDpLyLmM+E5EAHg7cX3sVidlbNeIWuV
DicMu2Cc6N4O+o305/0pWYcKBjZiNIeXtFw6FCCn9hxxZFLr9Y/7shAED7QUKDf1
OAWVyjjJNqBwPbsvr9+OGpNq6xSjj1lxKTOdxN38TYyD6S04z6ttJAYwqg2Ek+Uz
c/i2JuOMQcHHIfuEgy+k0xat4TElWFxfei9auhJDPsWF/81Wxmc0RHx91pkEF6BN
nqObXKgxr/YKTmiolrx1sQC1RHangOrIEgIugon2Kd8Y7xW/pBhYSt+AJnma2yJN
GRjpK8SAHe7foq4YC2Cf4tKOOTrwvPTLQAaUob89+wFHFcMVwyEryy3oOJrbw81N
EgTTIl0TF7oeR38gJszxU8ua+tKATUFkcV7vBGvl8Sn6JP4zvKEc6bLeMibj7VAr
2eAxeeom3WrKG+aoHGOz7s0+bhRUkeTcEx3JDCGtIMX65qRNR0vsGB+ogXPaSsTG
rP7HDW0kY6bXkQzT8N88y/9xevhMDu+qARglhL56SQaBzpw9p+W3DhXvIZWrYdiD
7NuQL4WJ3Al7hmXhlWoFDNShWhH4UN5OGWPW59IsFgLdmfBuJE6XNwx4h1mPGYDe
eGJ6cgykkH6h35G7i/INZGYpuZnoUju17QegmNEe/xzGLtjOrH47CyjJcg7wE9gp
Hx95n1lbJuMjcEJ95+eQLpgJWfgmEV+VJUc0lFITssjrQZxECj29yK+wpjQHREWG
POWzq1A0vc69jY3H0JLJhCivwsbdr4a9ABI+5Z7KLrvipd+1/yOXDGQYxuyLVgJB
4EmD5jDyCGooXKdHeco/z2Un/Msn+WETFncDVSF/RlIrSmaULWppIzsvHUPRlrgk
/UhkE9pTicNgfU3RBUnquXsPH21u4NAKDY/7cBEtEpe/I0V2HOiFJc8Cd9vlOyDj
shqPt3eNswu/3KskDKBqRGRNczqX/ldp8w2oXjqP9kBzz+Tp65QIYyg7aNp7b0p0
5Dwn+lmNzw3ELTNyegtRoZR0DFU1a0FGjT5StOVSVs521KPJfI901pBLb+iNZaG7
vQ9ISqPQHwrY5sY904Fy/Nkkzxl9w72nr26TALnaz5WzxHzGVyISrA684NGbXafA
L9LhGUYY/tU56OD7ZtDGGOU6Z3AA1M44qQGX4fCxgqiplNCiS6KNirRRIVyQDnNW
FADyA+45djixGChkbzfPWzpguXoeLDat/N+Vu2OgJW3vOQmX40YQBdfl/AJ0dWcp
ey/TTIfG5Hj0rrw5pVupywoTbxiUehy8L/8CRgc8LxHlKO+7OFcbpqjGckgG0ibF
97dwQMe7sawMFEhjxuCHEg2V89ylM+S3NHR2AQI8dQxT3RzWyA61BdzhEwGfhdvN
tB9l/f7IcwO2fxM1E+6lKYGndJ8pxw1uZCKA7gnJg+IlU8z+ktGWaUML5tgAUEqg
6MnQwAHZlOIKSD84BUuQXbkv0nat/vdMqX4oZzulDVhhBiEMd+AF1N2kEYt/+0Id
T6r1n0KxFKBB9fZaTtMH7P3p75cCshAu+dkAz9eVRwBvSubYbtD3UbLuGFkV6k18
FqMXTBl7FrhU1ukca2ppwpl6Wp4H0Eqi+jX8GFze7U/bd2MR0L4iHrQULPZP1E/6
Uc/MJhM7oThnBHUhD8RPi6XLPKY2+D3XDBVWuRvEuJY7D8OnciiKTLYbTDiSo0qM
EdkU0CDwcFUhWrACM9RXSaw0YsL+oRGwt0z67wD3aSwwFX/WmYLHM8u+HFVtKXam
8zrvRIOA+eqUsyENg9ZMYEKmZ4c+Zd96FjGc3sOUxP0PMJ2P9GjD5aGbD4jxJBH7
9iO52plnvqeOInkBSa5nYetCnaXF3HTBc0pam30F+oJ5JG+EfNnflHdgzx2+j1W+
spvwfqKQLZbA7E4kpwi4Z5YVcNm5MdYNEwVAEhayFlX9zHv4omPrUeyqfwOkM1h9
gNHaK45dlTDzpYAu3uIAjMBXVW7brsfkYyKQxtTuO2GH7CvsyJm8F2SeBMA2I8s/
9r5lNXgDig1XKCFwJr2No6D2TUNoQTfh1Z2Ki9DLZvLjMIGsCx5f0yi9rY7BNkyd
mbd+qU5ygPugym3A947SShXXdl0KjOBmSdIMM6bEgHWe7FTwqjDZxfzLh6SZ85BN
jiHlA6pFi3Wg4WG4UzsSxVwzI/R/8/qNm+Xr3rNk/lhy0ZUsxQe7QqbG4l39S1DA
JiTQUHISQ3qC9mn17yFWcEZfdvzkgYNndKNcz7gvGbLGYmd25rEUpmK8OVMm2dfn
k4kIJk9RFbaIfxiMRuUkpJolncPAZw/Y1t8QOcJJttytrLRKoWd98oUFBxe8PJBK
EUpyzFCg1R3GlF0iKUH7DK7jZkrbQK4M/2wdml91+c/87zyedCrUVdKVia4Vbnxr
2dTAW4tmkaqPpZU8gvUgFY0BiX4ncGKsswhYhXntypI97boi+bHlp8Go7BXD/BLo
VX224svpJmHf13f7ZTR7qaGyVQ1jT57i6Yfju98ffIIRy9Zl3cf0oVLYSyzAuaFW
FuiPzofPz6i2UEnDPDfVVyGgtyENIUn2dNO2F9FJbOm7sZIl4BJ94/mOyvotgOIu
VTh8+G+pUlxhYLvjHj7ViokEdMNbWB+byuvd2JHfGzZ4ycVpXOpmhck3WhRg7VpH
D4dWttlv5mX8re/325iLXs6tXRkmoomt6/K+AND/E4sX6gv/qb8vr5lTNmYP8+/3
ma+Fpewg+mwvnhHvIGVEgWVagm4kuIURGos26rJFDEwjJel2hZ06S7PJBV3kzfg8
ttOWvBGf+K/QV0Bui2pxN8KL4pShd50zDL2OM+Rb3iSOhwH7BzMpXVGfxsQX+44m
xxacYR65SYesC/sMZrEkGIlLMxRvkccaTwOBMh+1z5xbs+uMWjnvFMACpYSwMw9N
Aw1JtHChxh/LURZAU2+lL+9LkGW2dSM/JkuVedMTqcGQ1rocHe34Bb5AafpCk3Qx
N79lZ/su16ZIQLTq0fMnMD5i3SyrIM+AgaOSF3mhLaLVYuClt3gp5Wp8R/NED6sf
iu9eSifI6kQ0V3k9sNexRvlhq16Tl8RE0JMEklpfhpP2ylRivCg3beIE7AgfZHrf
qD8fXrYodvf6YamTXs0vXH+2eC7Eze9k+FcGDsNRRx9+ecPn8HFlafKloCjZgt34
xylWjNhvPdypDufvmrk1h7QmGux4+uH6H/CqpZZQkD3yi9YnKncxaR816Ol2Rb9f
QU1uy6y9JRQiznATZjtfa2YHGxw9gbWTkuxnKH1pcBCssqs/DsTQdJpGOMcfHDcJ
AXQhYQqpMZiWEQcqUlp40GkGjiJTCCjYBvW006yleb+P3OKIXtNVJmB7WrREXJBC
9G2atc0y5UeGbf0GXrsgyGRzpJs7O25/jeKYiYYmb6UxfIOpb5/BbcsibUBKWWn8
aKiAeUYdYuhuQSOZnwNGme8FZXQPVqlxsa18DiTc7DZj1zIBgPJsIsV694mCbiQ6
Xt3yEKdzX9GhZR3hNeEdGgGTk/UU8weEVzhhuttvPhSLYfqnPWyngW2tD+7VAUAi
mybvIelZM/VJCqm+RpP+xEmWEA0z3wCCWRJMbNrk8aW5XvMrxG06WJWMItomN7lA
MkzRDn/Qw7X0MPWgFKEvPfiBxLwBNiTVJMXaioYcT/1H79ft5b24f/lRrl7yab6n
ByIZNY/aFgfbozPPvtcyOwuJZBIsI3JzPoJVJh3P625L003ShbP4b7EsCVinYfUD
yGbpZXFKYh+u7dUc2xo5mcotdUn9qcHWUmpWXjSjDRiCEsBQszz9JbE9zFdIIb1x
6O02N8kDhGlAPoMVjKfH1adfbCXgdUDTjfEJDr4LAIinoZshX1dvcJON/MuRBlmE
t/EavfMQAGNc0V0eA0uiaKUtjmodlS1fCU8ixy5pV2JJoM4Z7Kmxtj6WdaqJ3hE6
iwBM8jS0PQAdb7oXDu3lX2DBiBOGDnQiXdNyUKh+zubF9+xA/IqKb4Mf6lV5lGLl
KNehqnpuOQaLTsgGmbbtGHORi/3njpMoDj+zPLjFsj97/5J7fuYV+Guwfbll5dDt
favYq1t+1KFHPGMW9hwByA2QeYzlFR9xxSRXAsidrbiJnl50h750QbL1Kh9cyLV7
cPvvuPq7ww0xIw0UXIXb2qgv2a+v297dl0lwUdMc+eluU2D7jexMuh8UGrzujl1I
gSfcR2jurfR/wExLLR8AnedTA8zQNuAQg0Mkfds7vJxfyzTFRL3pF76f83w0x6Ew
n6I803DXe81rVoytBcVTDQTrhnFBRBi9UDfhJK0vK/7mckSynZ7LCSkfelLFkSJ9
9zvdZE9V57khFAR8Rpk5oXhGL2Mc1Qr6mXl5mvprO6ToxLrNcV2X8cpx7ebVtvol
zvGiJeTsOzHXBbVE/6mEd2mxExbc4lApoEGlFgyOoAxzNsM3QpDo7XuyrozCZMyJ
JSNKb2EC7mIyEqfzGeyGggzV6UujQ2cs0qNUoK2a817qX6zbfMiSvd3RDt1usc6X
HJ9YxwxwYpH7+bYzrq54OaWyjupZIrW85wyPhwQKYIzaWdts/Y50y+BK0D+2m+pu
XSgjsrTrP3Tam/RDbl38aazccMkzGBDQ3UiWBATB65h3B7yJScBxFAhw4/vyTYXQ
Lh/P+q5Hsvgbu98NAp5FUmeggc7IvoR6R+BfYbstBGQGxA8SOwCzgpeu/GG8j/y8
ILta+vmZt/QTypJnUTwdH/S15PLEDr1dkTM9KREjmDTop19SrRs/NJKZPwXOZkII
JDPVAlK1keD5qxbNI4JaaJ/93DYSbNEqN0Kt1VVaoGcNBMMXkvwfndUQbS4b5psm
0Ndk8B2mq+65gvLFGCyZKtc/PRRPZ0BnoUp7vWeyd3FsicGc1A1K3MXR/qv0CbGk
XTmDKfTHJtYzmig7xZa69aAEV13tKdTSUbLaq6vUWQ8++izMwI4xdjccHDwdBgjq
MaW/ECUHFmYQzrkCPEx05wtscwj5bDj4zN9orTpIcHIa4yKTGI+ryHVcm2pyYOOk
m4f559ATOnAvVFwk54GhumOEtFFKt8YeBLfoj0ukDhJimMt86VU6hbRNJFce88aD
8RFY97+Ys0nJFbXJ1YrFh4qHg6E26YfkiAKEBhUhrPMMWLzns7S7zk7VaRFdUGLr
mQisl/6OxIx1EeRUNuutXsYg+r+W2QqVlaYCkKM3G8TQ+QmFOmnqbJGrOggma5KX
HNLaebeJBNgIJcAedp+ehfz1Hba6WZKHIqkBI/vAnrRem4VEie+DMJ3wfVu3WhbW
oN3NJQziCEY0Sd2D3LPXTNiYcLS+/GY7EA6udM6VJMT9HxpldUk+2p0Z1Ft51Kt6
UQguJIA2hvPdFKITsEVYhv4BMU/pzc48HW+Ot5N2ZVn0yocZo30LYe1Uqctmdghr
HgkTkGYMN8nbFMtYbQPV2mKJM9JaWle9MuH/ndFr5LUVrB/1Sz/Xb3VdGoEqinb+
sS+P8iRR6/yjBYGUQCQAtneL6/9Dbxv5ImeVx/qfAAB2ee43/drKehe/+Kdu8g+B
ULaSqSwamA+jwfCG3DgeZOgZKouEHyPoKlFYcGwxm3D+8Y+faH6rienUdv9VbZ1i
LzLa2DhkRG7UEbY2RPQEsu+Dc9Cge3oqyb7KN2AXnaP+1GNbDS7nQ7oDbS/aG2M+
1cK4/lNcITe9R2mlLYFj4f0qmSxzqQf/ulthslKlvvFHKPbMOehlRyyCtwj1bU1E
IK+1vmnLt3aQ9ZnSBYYdnh4qjkxJ0oewPYcbQr7Y+6fSc0wZ3NsD5BVqurSM58Nc
yITBWyztYdhY9Hi0sRfegBreEMLYy9MZ60+Hy+xRWpSK0gc3A5WMEzItuc3sYSUv
FbvpdlzVVDbJVCWiGaWz+ah65MLam3yYR0/op7sWe5LP3QY+jtNQ2vwNzGRW+9LK
Hz6dhfru78+tisrjZtdojTmC+bfsRORSUF4tdYoJaw6NcyBm9VvycGEHiCZ6qUu/
VrQGxZyelbtn6BujI2wTAiUkbIkqesNAtWUnw3CFCxwK/ekVdt9UAbBpPLSZ6NB4
kdzWmQvuZPYDX2iqZftTv149TzRjVYNj1C4IcWLKI9T7vdGA3xU5kLcv4ah346J9
VRv5XMoZtXUcviietyNptRIl5WlzAyHvlFGTXOcHJRECiX/Ss/VrQN/6r9Uo3JOt
aMvJJqqIPVF7BE+51eXDRV6dtVDg8mwEEI13q1abrEuNiUEQR7Fv58OGJpZ7mGwh
YvmtEprWVMEj0kGdhFxDqICpkDGNl2Ny8F4pUORH+wuvq25qXMvVlekZpCXTm1qJ
oVzg7kfNsn8CIS0AB9XWcbCE1zt+EyBE2xH2vs38UcMEZ6MrnXvioCGp8uaWdqsP
25+OBppI8C4ChM2xMNz9msK1Yc65cNpPjtm4pMyAxYVjzUAQ1M6frgXjnfbTURYU
BVSt86TJdwR7WpQ9/rqN0E4y/mjSkpL9FLU07gQp9QOD5w5TaVV5bFuu2DeSH/L9
Lc3lB6ruVOyCu/JeFtFE0L8xo9xhtvlJIguVcvXIDpPe9vNPqTcDqzPCoYHP3SnH
4xZ5VEeUPE4IvI5p9OcrnFPsyKb/up+3A/f3j7gwwrFOitTD7OndT3wFysiuY5P/
J7te+egiDg0YiaoaxcUYWP8PZ6XJq7G0MA+2Vw6yP6/IeDINiSUz2kAmbz2K9KW9
3Ag6D8Fi2QV64otyEw8i/GF0g04BljaI84UiN6tREtal7xM9J8viImb8ks9YSbcj
mgOGXRWSDKfVuX0BaZ1mfa9DdOyeXYghpa8khrcgJ9AENl8Non/MI5k9rC8oM0CR
5uZtp3aKQ7CcvMI2cZJZ/xkwRvLA/do2J5M0v+EXGdtPyGGk32up4Z+ewt2ox1M+
oVCBZkRgeGNMv/e2I+UlZt3DZQbQIjgv06NOyk7SHmk7KXzO7lIRgekUbQybCQmS
R3ONIWl2WtKdu4hKcPFZrTQfn+aH+bKGEaFZ7P/d9C4W4LdCkxJ3yKxXOH6Qk25M
EtvEmTIuoXKbZEWmVmnXdU2aVe70rEV5awJS59NfWWzP4fHL3VcH6XSQeDHSwGEE
nQSP/ZfHtCVrATkKZgSRVQ8jv9AiM5A2SYx1gg6xR56nCm3lbKwGa7Gg6wa+gY5A
VJDSG77nZ2Qasq7mwnP/8UiB1oN+ysH3cDBOMUMjhZPhHpahQBddS6xzbRax9asV
lsuDIfp7QuNZw48ZicW0ch43bOPQ9wdSuDw/x9Tksv12eb9Xn4REn67JS0LfYOjC
kyzB3xcTCTnP+Tpl5gEMtCM8gwWnu9jfF9Y85IxOyU0IC5zmCUZTclmJffFSr5tN
ImzARxJGXsjGm9SWDc19eUkpERz4VrBl6XlnOFK8jSPebFlSkwE+hyV4o25p23zB
ZtBUIAtL92FrJoLD2nHTFrgYqkwGKXMj/i7AR6aOx6ac5JwpI5HvxTgsSCpxAssa
qHK+JMFOFDg1IpDjVUHbt9TUkfgt+tRJ3ekEK/XS8UgjzP+aBUUYj4KiD6u3jjxW
PQa/bZNMoLFAa0DTBSKMhI9LGe5+zuoLGhLZWhVq+q5lJUVtsV2x3JxfzLn0yGYG
C8iVItaIgZceRjVbyYIPuPY7ltZCfWEh8vyPu/ZEPAjLEjuLSd25UvutU3SgYoVa
TKqI1VWINCeTcsRNC3VYzg==
`protect END_PROTECTED
