`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwKXseJvNn+9s16btUvPhn6CCUBIfEbO2bpUTYZPRUP3xnYsbnPvTklt1JqgOeXJ
fu9h2QRjtkOEv+L3sKJUVrWq8pFKnqhFXVZIE+i2m9jdNm0UVekx3RWPuEjVv9BE
6Z42oOeKnOP2zE/GwH5Tqouhdvzqz/ioLUA1NSx0uK0vlh7o6ZQgTBr1Sx3rEroq
1ZQkqukRrg6cPhTlBvfTlTadoruMMl4pC7CT1wCY6glOaMN89DEw6f1ChaPh5i7U
aJDPZ7yDEIGv7bAT9lykIiaa9IyLm/ST4zOF8JqZbkBHKfw0LcYJHtH6sjuoCBlT
yrCaANRkZwMFQn8uk8NQdHQskC8f8UVkcZdUdpwDtd7MghaQsNpQC4acNAIvHdOZ
KzIr1DG39HZY/uHTjfzQ3unhXOShQbwjwhjWHczH/FMFnn0sGyTSMKC1Npqx4RD6
pmv155NJ1oRjay5gaw5DDFaXpMvXzaNW67nPkqCgo64AQFMcPZ3F0mz4T04HDVGG
hZsGin253UAGTtjQe7CWr6LbPvvVS96T8xarH+axMGQ=
`protect END_PROTECTED
