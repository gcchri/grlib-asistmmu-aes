`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
23Bvel9sBsU7RNm275dwxrANSqfyuw4HODTE2zF1SnvuDZUdwBWUCg5/Z1zmd0oF
j/qQBP377WadSuqYA8UZtMCswJYX+XHddWdsNY208RqCqltjJKmSyTLKPa5yErMf
K/nGUfUW9sS2rhWZrJxkjMcA1Ehc5Vt++YEd7kwQuo0pmQ5aYn/7FLBTt/OEEdr1
91q1aCXEt2wLIOilNfEjm6Uj/CAhA2yCTn6g5KD5TuX2VM+iXuDdsZkVT1jGaXA1
EE1D8G1RvgxdfeqFc9Hrfbf2wO3z0XxTBnY+R1dX++onbxdhmm3A8Qh2ouy8iN3R
jZqAiJJ/QDGS2Bez7/J/D8MnNFMypWgknEbiiBk1yzJC5FqZ/LRzkHbvhz3U/9M4
4l9a1C256zGcouZMc2bowSDNd/yt9t+aN/Qy2my63YnZOtGvED80m97ouzYtaiWv
o749LLmqDiFCVnuv5G6SQB9fHck0QE9lUJJ7phxt2t2tcqnUbqdtFbgrJTMACSjU
`protect END_PROTECTED
