`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVRJnDdeWYzA8EJWbsVL/z+CEOJ7lpNYVSc8ToGPPf80+OseGbsRO2cbYr1Ffji0
pvsKcj/Sdgnkl+zKF1eEZnYRYByhWjgTRfrN1vPemnInhyrbCWeAOecudbeuQ0KQ
FBiCe87WHF/Di9xQ/mi1Ld5BApt0ODGlxzrX/KSrNZL4VbEDiPiKtyg+yOqOFBcd
jSvHn7eFbRb7CjebkSvBcAU2Y1MRl/kr3zpXklGLXDzZjorhtPW/UY/ynltdt+X2
1zllDtGhdItIRdd/TdkLcMJH3dAtN67brkX6BD/8Gj/tcVdJw5jaK39X9g54BJib
rHbwPWMEmTEcv9qqoI3caYBhu5NxXDUNNpNvTNWnbAOnoLherbtgwCwv9pM3XfHP
ZbbC6Ly5LvHKNILu4Pyum32bVuKo5Y9PSf8Vd29n0w9e4d+1y6vv5s0ssoEFmNEW
N342hcJRL5OxUHvc+Wer28sJG1aeqL0CIMXLmkthAC5fsfiR0YOwCiqAO2pXpAdO
jt8iJ3u6N4cnhV0cf/M9sH3AWYZnv3iS8XQIMSEqxANcENDzOV/XjCwz02xh/26J
P99TWwZ+wqxYCeAl58Quve9tntUT83ja6xj7bdbFw4ZGGu+J+kX5ld7tAYXLAsDt
RiLMOBc7/VVIt5hgzqc+wmYpwHESWYUZ+PXA/Y20hOO/mFPr0LhCDbgGOXgT99gi
`protect END_PROTECTED
