`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xddxrmJCZd/mb9+QoSOawNxboLLh85sTs9umrp4Lwh6Y+z5BPVzNncXTaOcAot51
ks+fG9Ce2Z/bZ3AHsIRoZmGg7v8amN7uJzURZpVlUUfHH0qtru3Y8roVSAgmVVsm
t3rm5XFMqHGlI75qo50/WSFAElW04w0tkmsNOyt9Tum3qi+R6t9jCiGYvsuVDBZs
ZMtzJHtjJtcnwSxsFrpj++EzfjM3Kr3fFCNa/HFNWZGL/J2souEPH+nz4la10YYm
WsnbW0XaGLynkUBdLLoQOO0fM9TUZ/04VkgN4Cvg3k9kGwWraE1qhPBifOToxorb
DwIbz1+677rz3iDR52fFo2AdiFUtX2wdrKzxyhFLb6s3OS8gVnAdi06joWQctXbT
VT/yWuSLx6YUVUsnaWCfEA==
`protect END_PROTECTED
