`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wf+dHiSpiUYaj98apMEe92EcTCGXBNAXW29F2BzAgpqHgC14SW7xMeiM75wxdaqr
1vYXA8Wmu76S+Ok2j1LRrbxmRnuVBw7jzZjUB3TW8BvJ6xil3TU0eCS9c8exGW12
xgd8XadBlQNRTBQUDxNalW2Bf78zclx3QL5tdDPjWxU2EGQD6pkjqc+v9Un/mXjC
Y8BRa7jyzmv7Ij4WKeYavTjiU1/iM7IBINdDdEOggX2BbMg2+AnueYpzn5NmqTHR
aeCGo7ldijMcAEv8oBdGBUu4XOp5P8wZaqTpZ5YmJn6kbEwJMdlWEw2KQXl6NZWV
5TVyz9sNxAveM1jk5m8nLx9Hnz/2WGYLMVQEq3/p1MyJc3W5FNI+Zt5gukuJlmLZ
IitSwYgUjWBugWkHcU+K3x64ZXNNK/oYGK0zqf9MTWYLfyKNoNR/m1Lts43rezsd
x90KHIW4wY67ez8BOQoPuAqR9uTPW68T5VljUzhQaUucmPXTOD5z8hlkroyICcTT
rgPqe/Afh36/WcrJs2CkbAEL/FRQsecmGDa8n7xRG20lIpDUSJ+idpgD9twwl66y
6mvsL3ZMHsleJqz7Nvwsgz1TlkD+P5V2JFBsviZNmVHHp9SDiagW7n2EZunI0+rQ
gJid9OCL8zL1FG0TAT3gk4ygUgJUjj42Q6ojtT6dV0RDSquu5dfvb8Xx9ZRh9OjM
FW3IP0qbU8mNf+wDh7poeAMacqJQ25cVkXrrV0cu3XWwpmiugwyrq67pA51dF1eO
Tnl1fu1lzQe/CQYmtdx4KTzN7akA1FkZJ6+FN6Y8b7bna3yDztqasuc2RfeCGQ5E
UEQsO45L5hvwXnTiSzeKi9hzHrrBvBy5VIGfUP+mjBfkxMLkzbprl4z/OVa0qMcZ
yEn1T9ETsTlO4AZa91OsZzqWJ1kjpbLuuzcWjExOQk/JDPW1uaWhfQbDLCwvfqaf
cMn+8FaiJOR9XG+ebWdmJO79FWq5rLRGcTcNHhS3/ey0gq6NX1CkY/RecTN228+s
kx+ITJl6nBJcgNKJWNg+b0+iukWmjr/FxgK6VwhZ8VycBHiPLsBt7Lktce4o9ebk
ASejbeP4x0CMX6o1sZZja/QJLC4D1KvQVDaFpaf9u5D5SeSpN0l/vMfWXYYWatG9
DEBr++bfWmvQIYGqtgOPrw+hZunyLPq8p28E8fn1oERCJT1AJ4xU+ew4ysL0UB5P
Vi4d9rmH4982kHymML5WQkiyXpzvV/9AY7fyuRLWPLYVs1tOjDQw08EI69Mh+eNy
/zj95r3SpPea9v2FKJ7MslUhMwRXeGhtvx+f8PkLwY3ujXQGdnO16LcmWBE6bNfH
Te6AB8sQx8Y3IUnWdtNQnklQ+DbAyc59p2Ij8tgk1t7yaTVx3WSj1NNBK8LGHPCe
`protect END_PROTECTED
