`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wrJFZAyt0YXzwhW3aS6ynLYY+B+BkD7cZcHDjpe0hIGlON3NIkXrrJyCACKE2sA
WFJIbncXG5i9AOBaYCB/YLxlAidoiII/vkmxVPXhr8xx8eMf/wpcQ6ZPB4RuEjic
DymwYoffsufHKoEWveoCtFKNKGf7VObd9rm90jxjXmFqIOs9Zu8h+OoqG1SgmvJG
9EJ4L6T/4O/XRAsXqtXwwacawLZhYSrp62yTPzrSaJP/akFf2ibjRHDTuN/9Piqy
HfnPFQdtJZ77ynhtFWzF208DOXDoluhmTnUOqBJrtY3lsuCaaivYbPza/kGlqIch
odZgmRwh72NDcRmaLI3uwUHeHoUYx6oF0AB8oKMq9W6Uh5YYxw55ZOW0qYb2ydSn
dReQzqI9m0uPndc+1KLZnLeWM1RoXO0OF8s0F/4SBqq6goujLJk6+1e+n7ZgEq8C
`protect END_PROTECTED
