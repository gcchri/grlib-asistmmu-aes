`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TvPd5n/82Z6S2hNtYkMp7aYqVXPPZ/Rq0ir/7L2p/kPF/5nIt4N2d2U9VCYsPSpV
9rB5xbQlzUOGYQu+yheZbCogYIuMQxRlJFfgmj421MvDJOMMt93dofDH9zZHBtxU
kQJqK71ezdh2nPHIWUmFXScM+yaCUadXxC9eeBYj5bSoQF3KsHmBI8KC5q5MPtbI
cvxzHAQalyMPiW3im2rL/C4BHAVXbT2BahJ6FMohLWZlC9gLXwoCfrs91Er9yhkt
4VoJvsNT+5bleEyDqJJIQH2RT6ESmoZS5rEwcAItOEO3wbb7faVzhEbxZDIs6vpd
mXEo18Pb/XcUTLnEmJBbCn25y2rvUkA005alKu3KSLZPpw4LDtVjR0a9/7La7gLg
yc4V05KAZgjs8M7ou5ZUzA==
`protect END_PROTECTED
