`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dAGPSjoVmKeAl8eP5hjoEKV60FUCoTm8xB04BbqhmicvxpDfHHZAlcUiC+adjc4l
jf524u2n4GDYXWzMqdPM2MKME2dwlof6t+RDoeu2ulcUJ+JVHOJqawVnY1zNcDOc
KD8U66Lic+ytlxi/NJhIORXkCnPYiJ1tzPFy0iNisSqely56zEdXg7TzRdctlDnw
57OP/+X7RZmxwL+Ag9+8gs/yNmKdK6zIX/Ax8qbcp70Og0XcOKLELM4vNUSY3Xkl
HS5kFnJHtbD4c747CSuR69WkGX7y4F71GmBPVenH5POUKdQJh5fVNm0zGkw/DRR+
jWhp4KfAlJTaYNAbv+fMYEdTX9w5w4u4qz5AfOxRHCLXKwTqm55Wv4ZKH88Z9Kc2
+L6qjL6J9AXYq2l2RiXsQGetm8jDZekp7TmtVulaDplMA98CI0Yuo+r/exdevTYS
efvKVA0jSafOiCvXpgpTSJp2qV1hvLtplbFfPFUdOTat/f6Py/W/wqQIioDm++N2
0IQfpn7E0Mw3ONAlliX/eEQTvVUUQw7zzFLTpaZHVyNUo9eGDqZfDwccaHV32Sx5
`protect END_PROTECTED
