`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IsNEc7a7zNjw9KTdJB9l+a4ImGY7Icpt14o9KhKBlG2+siK19Vt60Rn3+TWz4jdK
rcXMj2H+tbtOga6HEDhwuNoSNztlqTNvHrt71jBvRxz8lxC3bU44Rn1/s5pUzzuA
vhMEfeQ9GN0HeX3orPW2puwxDq3w2kiOlAMSlOrX9WSzoYdhxBdsn5BNtxeF5g+H
4jfOI97cmZVfBhDmaqME94vnQg3mb24AsBaJl/TsB79i+vvNR5gnVtQANDhi4LUu
zFUZ9h4hW3q91+g4LSJ4T31P5LqJdLeuO+uxSembnBU/9MOxS0zv4KD1efuMqnDB
Jxss12Zgi3AKiKU7AV9CiTnb0hfABwMClqaEysV2EcvQUbFm1Ov/kI3I+HmW3gSr
QNg17sciE47fXG3ets6VLXbXcuyfPVrLl8g9I8QN4TlLkSfbb/U0wk86TH0c6aWs
syQibTHVZynbcYt2aP22Jf7UA7fQtqoKZU4iv3UXdR2NYAMq7mT0JEOef8P8acKV
`protect END_PROTECTED
