`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tgEcvOCY8BYPn5iHPDnXeXLNNuW0ZIPjhjCZgeV8CnkceZcmIl8TCtnv741CzDr4
ZnceWWk6AnFKK83OoCcv2BzdOPIzeBlAa7WYCWwn4QhMOK7o7LFIqjdZk37l7UJT
9AgsuneSRPtaTfVuG/cdpwxqxYhvzWD4x+hdSVLHWtozkkjpZ1ZmE6n6/5w6TrLe
DBxhNVs9g5GO97mLnjsbAulAWNIENgnyO0+dODzv3zgQAamnGkj5voF1worLBP+d
3Ewo4F6NTEflUtXehmUO3vH3ayEhtogOvXRgSROcpQdLONUXuXRM1q9MVQ+ZitqT
xHciCohYjI6tGvXtJzOEBBn5CYqTWWHAKvXlUBRuSsSITWBb40ls7vPtskoyrqZX
SpALrAQ4jNozhGIkfFpZh0svTEuzhquUGYPENC/UXZTJCzICKtAe9S4hGbPgYK37
7IDzL/gcGZ/gl8EWn8xxPxDNvgsJX/0KUek6hq7y2YFROusBDlX4xXNeOANJP3JI
8vcYRF3yQb1z+FcuJx1f/3jFswm6SS28tRM1+x62OsjuCO6vsNyJQlRgGDBth3Dt
PSirELb7nQVDTn3QFsqiNAhnv+/g1pjLk2b+NhdEU98pkTCbH5Xca60nHJIkWy5c
qSLobQfqaFJ6m46z/SnVQOrIHWjRCuOpD8SNmP+xaYuX/V4UfLs6tFz9V0LplCXC
wvbo7v2Tqr0BT2eGoDfkKgGRRiydSnRFP3k573XsfTuePCJ8jhyi6NOb2+ssIxU9
UUQpnR9eGEvnLjmApJCFF7nEfIW4mCAVmCiUN8g//+nofIVLT11NpqJ/zMBG9rKs
6tlzDgXTxsWSCauzqzaCOW9r2n2+LlFdgQXx3NZBeSKKgeCRDBa4r7j8h+d4RvH+
KbMFCcfogOn4vx62vYFnYySpWHV0dJxFWhdt7930HlYr3/MZJ+RJ3U87wBHQAv59
en5ZuitA0ks8aNucYmZcYEvG9mudkSrOmNOPgJ5hlT1hh7frBK0T6Y5LLU9Hdqeu
`protect END_PROTECTED
