`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJrSJ0Ndi+FFicjtiQQdCu2mcB1anjeQagNuCNhJxmbWel6Jg/M7nXq1vTGkCI1f
kpeLBafQsTIcgdVQWFJ1z7SiLYqz/SNiPkzl2thEwv+fn1d/G4zLV7RlcdRTHNMk
6anm5aCK0SbqHO2Z+rZYNO5F0x0Bis5Ul82dpFMhdYWTduby5HX3OY4LuRTHKEXJ
SoHLIDEjtD6DJtyJZwXwaFtuHExcWV+t8G8KB6fpJ16kl6Xj1Ih8UdLlxrLxcj7m
GupQeKfTXlYZFnI5EMp0Wzkpn2r/7rEIslBUcCT0fMfJO27NZljZ8mSmdkTBnILT
lpanDFxpfFPFH5DoEnLoeYuIjmWAu5kr3DF8TKonk7MshSc3bgeOyflt3T/YE6lD
`protect END_PROTECTED
