`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ynqf5DfR9BM1J7yq0uufDnccC+kWIr5iPeMasebCn1ndQ8LOacTsjlkkI3fLloiO
PelEeDBkspbPuwz7noTgtIFx31MWXAt+ve0K0oupyO95y09cuVlpIwmBZgPdM0qj
9McVj4jZVW99P409hlaSueoZwpCFbVZRbSr+ZQ6sh12hldrSaeiYrr4KCEnbJWMq
Zz8HW6HS2m8lepQTb0EhnnIK3d5uLyrUnQu5vzgJbGygGhllVc+E47W+LZblXf5R
NsyikLuwrmSO7emITW/jOy1b2yP3lmxaVLC5Yfyrgu6CM4rpvESWmKO3IQPALUFY
ljxvyfm19yT/dKLt4lDeXw==
`protect END_PROTECTED
