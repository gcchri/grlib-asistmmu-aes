`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viFnthzUJyV4XmcvEL0B27D6yqfdG19lgRuLvPeYdXpsbjN5z8t5hLO4n93Lbaqm
+nwfefrIHaet2ZyXwm9Y2FRzkuscfBVk+mfs6tRfM6glmGstaKAgJ/dpToKHQNLd
JDcYj/NMXohAyEYxVcpVZhyEPF4oibTDXEdL9qxfkAOzZ1QvQwj2KEuhXJGIs7ME
8icWoJsQ7ADi7a1WPoDRqv4k01MzQVXJT4Ii+hDirrZJTWe4fHasGdt+CHNvcztK
O70XB8eBlNJcp2nA+Ba4DuIimHzXSL0H6QGFvMuOyTE9tUmJuR0hRdys1OBo552t
iv52hYqxIfkgLwQsTL1ioIFWOkY5fZvObtN+L2JUP4WmDFQ5AGALpz+HbHcNH4aJ
G/SPRCD29c4tzy5RfD782wysMEgfjecbeXhTO8E6pd8rngoREAZdXRlQKFcHCPnd
Tv6ghJIsfxGlYbx0NRJ6Fo6dzpsI9ag/Hz8GuryQHOy47BEBXkggqaBFdOA161aU
XlfdhhyY9WcBz7B6qAsg125AyZGpnrBEDPWoPjepx2umKOZHhabLH/kLN6/ok/LQ
fhbHQilj+PmaSPAnyJYDD3h9Y2WKz1jsECKsJV+GCSBHlRK/O5lEZAwgO4g+RY0j
2QxCqZ7TTy2v/rhDFkYOZxAUO92yNOzkCxFPDKGn3QWyLoMpkKg4LKPgAKCuNo82
NiJLUfCyHQIw2n65UINLFTPDC4gOMGmUAxvCfGamVx8u6DXylxQu5cFvjeYu0oD6
KJCIsO1etWnksIVzzIdiKWfAaZcK/HAAnaOouaWib+F8fAGeVLtYjVtdNUGKpOd0
xIphGWn8tjKa5cf1Gzot7ftnIiCh8wNgMzuI87tQt/oIKcs04EbB+UVLQ10ryAl7
OSslniAgbbXXUHTLshlhjJjIuxztdb35gXVcMmuutmA0cYM2fHhGyDFcGoH07r00
otsZhtNeJ9JtWfcFPujsHu90wzda8p1LyJbvQCUmQebiB0gqg/K1xn2G9EnPTgy0
Yp/Vmh3FHAUlSOZOI/nzF92ICScRW/NpP9EHLACFfz57E4o4MokzU//O68bFSO9G
sIY6l9V6jPNMUugcGZiv9l2R4RG7YmGyNIYoQmRMafm4eawlPSh4bWUsrxUgQFtM
DT34QNFOOJhjbydhBvhbi5TRvJ1TJslNQJVpdRIeKyMNLVP140fBFbWVE8MtpX3U
qXL9cxZX9rGbWNEsCUaWCDK2nWRWycZalaRRXEF8IkOkhcHaOlOs7Se0huBXBtZq
IDfrWrUHysmxLo73QtM08ktXMdxACs7L6NlgB3HhAJXc2zbK6zKZ1u9NoS4zhcUm
aYyUlxfX1zKPSrayPacURkzc3b5IxZRf9fc0cYyJs8twq8ruIf1yfYjR6Mpon9Tj
8Gj9FhOw7Y1wZQBmoWhBq/14WbQH6b1WqkFyYF8DqzGALSyK4n+Me2uczRWVeayx
dcpTeEf1LJsDvSjZx11vLxxrD/eWdITHAVg996wLSBFCbygenwNcexF+R2CyS+cW
IHjSES80Htzk6rsHElZZoZImRyQGNNBRcSo0T5wjOQUEZglNqmPF829Oxis3MOTJ
oRJ3QnnMvfghdCXsKoQXyadgCq+cyDfAAr4cyU+vRBGat+hANH39fTum57nhM82o
QZy7yMIqFPYXj7+NuvbaakJzCE+ElHA2wyYK7VpTvQ6gvqYcgO5GGcnUFhN7jF0G
976kCZLMxpCcLMj9AUJCZCwQHGV0K2l6Kn6zHBNAp4R4YnB4P/CnSlNSXzsVRjOC
aSGFWC+0aQ0oEp4GGeNt6fjyTpQ9oW3M5n0KxDAZPWjfxPE469eiQF7fqHGlbQ5N
jU16jOrKtrrK57yJkRuahYaLo/7vGrbJ0+dPyLDO1et4/FdRB8g60znKPa7jTygS
d0j2vDE8UnlfDpY9uJExEL0tzBL0aIsLDRyv60XxT33Bt022S0uFAriIQLNpd7U4
6X0GAioviDt2YJtqa92+aEr7k/gO7E9JGrfn5OehG0qdGHF6+obtaRmUJ1JfkF/Y
baBLjf0rfKgVGsonYgXYkL8SFgEsmPRTomQK9oJVubiFbZn6wgnhlEPhDy2u01Os
84/ZvCBar55GPjHRWmEE9sehIgLHgEX4MIjjwbZ5oWtY5NIndo++CpFIfB+ftFrF
iInkC7AB5JQ8MM6Mhzxp5yDI4D8Z1K4xke3cxGtmweR+XwFtim9I68EBZNRWW57d
O3d7O0HEfVvPNSXQi5p64aQq1BJ1CPJIPLtSzadVEmgMzTlDDnXlnGwwgVQ8b7av
tLCOVzq5jROkRw8Okgxp9l+KSf5Zbk59wgUwRtX1O2kEeMB00mit2h/vKOI8roVL
jIQKI3sx4IGiQ9cPqzNnTfdAJI0NAjylFtCjRV+2/4u7gv3HO6msVvRgZOGrqiIg
5phQ8eNb1QeE30vyCnWM2E0PCRxHijli/UKzhbF5/OJ7pNBcJHtHP1joeyhNJDCn
5mmcAHPH2ox/uD0j1KLSdbEfwLKQKB84iaaI7Pp1WPQ2NNweQv0YMjYHzA8rQMQ0
XN0AYjwhl0CeksqkKGG9yZesDHVPPv/Xiqzx87p8JFIUR27o4becGgAj5t63bGMZ
dAe5G/AUYlMMoEFqSzEfXj5BMU5RRfsTx5uORlPJiBzj8cFfBOH+r4WOyN6n2unn
p++i07H7pnETrGr2kzDA2Q6okeMYS99MF68Hntzwo/CiZobs5DY7vxxx5WA7cm5d
3md5xAEzTrA67tXBMMR6JF/wkYIQwFXPLJa48e/tkpFvmHAPmdWMy5l6cR2W46ih
dIpVpXUFc9LNUTZ9bkB+ziZX1LDHZksLwu+v9yPKQDrOs4FYnmxT6Vgt1CYyKGHv
K/uGi1cYhBcy3yGT8Y3qnTFpdpYuIKT0TZX1lcFq8+ra9GivAJwrKvBkUtleRGi+
7DafbAmJoDvycu1npfYkK7u5dwbru1TAm4eYbPfpA4fwZkc+dSmtextSv5dXXt5k
YW+YeM+flElBRR3W1XVtZ4bgoXsgzkG+vxZLsGp/QwpignpDHIrET5MEJK18P4L3
PQNyyM9r6c8tgye0T0Wwqzy6QfvAv4OKhveaH1cnDVTVIxoghyxZa8dqBSZH6D5M
/w6M7XXsk+0iLWpSYh8NB58cACuK0l4USevRKW9NPX+xU/sSxu9dTVBLSVHIq304
5bmEyoL6+jAp8p67PuwK/YyA8BGA1Xq6b9UPqbaf0pcrJuvB7V2HpkxIoFv1MZjP
YmaQ1f0eUiURni+TZCLC8rYzMALWG5BI3m2gJI/QwZ78CYeHVDBgHngcYMysoSka
SX/9IGL/z/rghFNKa3TO2Cz/rR4twdDjrGbP31xZwVrETkYTr09GajK/ZsWcsK8t
uJcu2Iq7kI8mqWAwUzpIdKYPvlkDp8arO837rt2U2LDNcoGwLoAw8/Ufar2XsLwT
sgxRpwmLarNW3wuDHqqE4jrE3Hu8rV79GPjadeR77t4hWqU4rmwLUXarWzKregqN
BTw093XLYrYWloUc6J6CLLw/c+EZqTOhvRlRmzZkz8Dp+BdBvh1Uogb7ZuhONaNI
koGHw0m9pP9QuN2CVoprHd3afBoQSD0gPpEl57JbRuIHJBuczC8ZWDpzAqZh04ZA
zbQGA88sohIKeqG0h5YduTqAMir6rc9HFDiq5VkLbesWu3bPLe3sMf2g/5ed0AHO
M23HQd//JvL1GvUploKMoqkcl2Pmc+UhSkLZ8/ti/K9WV5CfHM0m9XtMpRuvc8V0
UfkH5N/p/MLEUUGWBCkVo7IXyKjk2NwduSdChjiN1pM13KhLnDNhcqyhVeSJEPgJ
mMfhabxDgXPAPvfZdVqFcvY/hRlsthzqc33aYlrW2Gb6mgZi40cFr6ltLdJjTQpq
Zrmh9rmEUCyhxkN+XKXIBNlGQ1+9CJx7ksTXOpDOqcKBRBJUp0VTfVhZC1a46DJl
sGV189d67q2fZ0oIQgN7gKcOZk34glpAuVwEk1pAB3N15ItULk3YpCfqZ9uc9MoX
8u+gvFGiBC8W1j0suJxHOFoW5lkrEEEinfF7smL8JecO9wm8DO0ZAl+DqYdSVLIk
e6mERoxEaU6j9rByb+5soSa2vExYbx9XjtE2xupP7UnoDQ4SGnPR4LmxDIlPPQ80
JZrXDZhPNGx9UsyDvGEifu4T/4nJQrFuZ2xb9AsWztC19kZjAL3FFGxBRSazzZW7
ql23GUy3Q2HSFM9ugzy8nltenfcCHQVHZTiWmbYCQiac2ruTQItdEu8XIzZLNT9K
+7s7ceEe/q4vaAcxhPhoE/uMAzLC9Tc3AhBiaLzV98I6PyE7kc8Lb8er9DIDz27H
mNWQfkHTnQAx4ytYFW3Xz9pc05TV5AMJvHzTaNV2BfiF9ql1wxhLJo9Pdwu0FvNt
8jEX7Pqr/vQrcR9K/ZLi8UCzgxwEHQZhcc4RfkyngWlyWAxczUuWUbm7Mhb1nD72
FzbTJCazPVnLH+MjttT1aS2QpqSV4NGR1oz4ScnV+LBbvaJ3knnXRJiYKClxFqoy
K7kUtAjBG4cnwI1Lql/3QkC8HQFW26iYvL4n0wt3XiN2VcYVQ36tiAjg2ikjKVZW
7WdGrAcKSoFEJ42Sks5n8fyJloi/JcyjLYpsw1uSu993e5uW/eR+dRowZp3q5JYE
FNluGKjVfb32NheJYvOFvmrChIjrjoB2EYnZrBn0gm6hzu8ADNyUKtJiRpx0HS/D
CG4X2fWpWd8cd1UsOsL9mP1/qzpuyuhlgmaImmDRiVVx2PPxRGHRAUKw4Oozwh7L
yabdcB5bxBtn4L2i/GdoanS6+kQkZeP8Rq/kJO3CQ7Ny+qbpbMDE77XB19NCLLUE
r2+jwAQaJPFqT6BNxYSCdESbfk3inHZsc/K9DS6EqSG6PZpnVw5grVm2+MVzip/G
fr3VV7c21WVD+C1Eg68/TgKuO1e2LaTnd/Dpt185NfHq0vqm6F3qvd3KNeGixYbJ
WQrGq1dLiI+Ux8armBVO5oPHBSzeRhwYIFd7/1WJ/BvTBu991+XErW6rrzUJijkI
S4eCxqebLScQL2izpn1u5o3SoGvu3DUjHO+fVPlYVFi1g+gdjRLJlT3yO9MPqPSx
/G17xudaXXhnfBPzHempi+OlqLoxB+7Ssekz8feDddq2sEp/+ylt11z6iS0AHAA+
/uxsI+Ck0k3Sh3QCBkjdtekZzLTAY2tCvgWRt2Nk9XJ8v5PeJxmomH4aU0ZdQQQ4
ygLtBKmhJgPjfpZ7HdX8pDa3eW+rsTe4P8P+0P28cjGrbe+6D+JzkXpEFO14CuYX
0RDXjdz3Nw98JUwi5DeYxj4BnLyM3n6h3toG0hS6jadjE5g/milNF4UZ/N1uycdv
WQSN9lhU3J90j0AP/uvrs0wQaSzKgOX+ACbFr3/FrYv/1IaWF/8jluvvI9pMIy2r
3sf5jXvaf1qjrcJYe5Nk27KV5QgE+LgBAvm5nZGTc94o8m4aRTwgN5bRKc2vyzjE
tOgPafBGOUhKCSVljkuOyW2L9rY7jJqQE8bW036caf3aPGlMH4KusA19ocrFlzY9
lb3xvK2B7qY9U5C67J5PlV5ygNlcT6gHOkoEpGhu2QjIQfU7EQmXino2Hz8mYbwL
OP00JJCFxKN2saaxEIpI1ui329ZSpWQKHiyxXSrbrQTeKM6+E53ETP7gN7RbwUDg
fSXDLwPiaGyCtb2qcFC+1n2dJqFjij8Xa/VBRfjKSaWDNo/Y0A8GYmgVTzUNa8GM
WLa3yZ6z0WlTUvdYdzB7TiuxxW7CjSI/0Z/dWF1/4FHUfyXmcHnI41eWeKNcXKpk
SQdyjE80v6Ont6HE+Qz7D1M6y1HKPaIe9ZjeieGof6bgIQLLvm5FiXHqdSSjEIwU
ofIvTbXV8Ejckw+huIrL+3eB18Hhal8QATms2xY8dtR+jV31QwC1sWbXWUeEgOK0
`protect END_PROTECTED
