`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jXgvfjy23hegPYEE5Ph3ObXoogYBLNMcZ9hkXTOcsu/Ee3pCl+ajHkLeEj13vXZR
z+3Cms5/3IheicLd2b9rX6UOXTmEipSS1dVWOK01TW1s7skCtss/SfI6hJFp30Y7
YO4e4eB+2XJZHJ/5ppMcnQ1tdiLmF37QI52mtlAk0PFJPTKO34DZzaGHKHIsnbiJ
M2oUJCJoSGczi0PUzQMHT9WXj9Nj/XafvXKdmLEzIfhs0n5dEaQ/3rMB2zzxKJVe
s9X+peBBl80j3pV/4NkaJ5c7N5fCbWZRESbZiDBAE4SfnoHirfP0OElV0FWF3l/7
fbD7/60X/kf7LQDhktK1JAHPF9N4wWgk6yJVmSO/UlrdYw2ex7X41KvNqJU+qsTZ
BMD1nmzP7n9ZUSA1N4jsdVKdFMYrAh5DJ2dkVA9FRvggoRgI4lmkJTH7rHGzGZgq
6ZJGiaKJUDm78hBpfRNZKPR8LDI4tfXDSjsmQDlKHSnezszgggvkDf/du7w49UDa
oePcnm+lWQGWOa5ocUSsKmfECOHuZHMqqxLVXuB68FWCU55K3yP+FFSMlxhape2Q
6MZVZ43qI0WyBf9mMT3w0LtEMpyTdQqhqxiwCsq3/vqkr403V59Cqfd85xAQFdYV
J71lWO3OsF6CGP73i1F8Yu38JUv7LFac2Phd/J35QoD5sEsFX83AJTwyIjG1NNOa
OIBEwNtSNwOCv6IVWRIWo3WfnTYSOR1ZEPc1U+nkgpiZi553R98jCS6amOnmPtUH
`protect END_PROTECTED
