`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wE1fBpXtth1otgk0LcZU9R94/lNmdMDAtbl0Ps1HKRbx3+nN2Z5V8JuAbik0PPLn
q4P+T88LeVDGgzV7y6UDTH8rEL/EOUvRPLtHItzcuXi6vVOAmFq8jQl93uX+aLET
3imQNR8zU5fMoGW4w5qRp/NHNcP26OilmoqtQil1IAuIeE0qfILrtScLFx2qF2Kg
ceb2k441nIlxnA4EEM/hVDSIszgzrlBWk5uuJjOv0xRZkFzdLRCDjaLgujWfjW8e
Mfe3N+/COMzCRTlw1HriDaAQLIhD4qwgRywy3VbVN24Fjh/ncDH8SP4mU9KZU5eA
IqrU8uSwhTvgAmv12LjSj41b1Qfi7F08y3vNTXYpbfZzQLWxqdk+nKWyKiUn/WtB
3EECwonLUSLt/YNP2b2wvvqkkSFRD2BuaLyi256DVlQ=
`protect END_PROTECTED
