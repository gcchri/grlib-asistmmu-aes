`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISdlannkqdsmFvnxs2cf/uSMGTVk4OpgqptwkgXbyuNR2DvpVL3LdRXScZNRHRw1
GRf42NxKui7ZwIehCLiRKllvONknp69CgybteLDoHkm1WTjs9zYOiENT+bPybrAg
hUP4eNwZCfiXg9taFnq8HHP5gdFovhIYt2UviE61QlTKFApIANxgm1oloWwYZvGB
wJUqmAH+Jhk1P9zB1jyZESBrVk+TuGRnHMnJF0YZiPS5FfTKEwSGgPF03DwZB63w
7AwNrMgjEEctYAsB9qDgbeXB+Y4uuAmjIAkRSV4zBCLJNkiCp4srvJebA1JHZ8sr
zh9dJvbbK3/w+Q1iKdQaoOjEvASvYBEaI6dmpJQCb9IUCSKekMfCco77WEP1OGyi
CcOs/5QGd2pjA4ZuRSF4HdrhwQ7DGnYaEOsvAXjz5gmW5v3bQUCTIlP+qgALhix2
ZGStQmVupV+tCE0Kwyp4S3WQaXdwc8HbVOnVoRgNpOpHEL6XalaRDuT2zQleX8vh
vHQsKmgq1Dti/0Cwg1E8OVP0v8cCw+IlEba5ZgT/Mr3KB8RBf3f17NwF6SDBBwW6
MF0e4ZJCpqncOHHceeb74OzLB1Lk8qx+4ovvEU5gEQ5rfiBRtwecb70raTgvsGdX
7elA6/4xa6Fsms21dRWgO0q16CfszXY08VAa2YTOZMECWqh2jTfJqNV8j64kDZCJ
PoeP/OjT2JtzKUzRTxQoqgJobwhv4fqKrVf6QrhNd+sFTJ30q15tjNZ50hb2a1hT
zGmH/z5CvQy0TefRhnFrTRocxxgEthreskfU5MZpVYN+o6JQlFdPvqVfThSbuu6N
5juY2TvJf6+aW5S+hmgnt/ktc7cBb4ooRez+tx8xzPK1wHLg88MQVzOSExFle0jg
Ufs981mfJfgwY2+27ng0VowMUnUR8g9QnzBXDBc7zIhHNeZ48EGlDwhw50WHSv29
39Pz6jWuc47CTyraLieRRwmlJGopC7Lpnv6yVQ0yG/whR62qSVnqV9l3osljmF8g
/aIVtygQSRZJtdwvPx/xUNZqOTq5C9O//jgWPqmQoflk3XJgKQGPXPPoMUxuR06L
VGotAuyHQc2nSIZgRS4wRTe6JF0192dVwVTAiEwoRy/K8Lv6BN8WekeIYh8FPrHk
hNkvOBYLcFhAlBQp9WW6wGnPUZkxjSd67rwfDxc4wqRI6IEdLNCJLU5JPTlNgH8y
AHtwOECPW5I2pt6sfRhEsGioVNsmQCiiqqD9aSiDGonjZDHoCOkyrjwjRtxFJUQt
nZ+Pql3g72GYO8HYszcd8tynr8Pg+D/FFmmTtTLj/x8haMY2nmTuJAdknnUMNchf
yvA79bd/zUSjpArVGpjyv4g//EawbhECP63Ah2nMLQDbIudZGGMdpiVezSZmpKe6
O03x5K2sUaKjsUN8e+1Y+YBUOjwhTyR4XVq9ZEquq910j972p3jNXo1qzXCr7FL7
jE8tEO75+Iq/vWdF1nqZrb2lT3JUZIU3STSFYnzioAEQukY8PK+bRKuoiJpOOH6M
cd6H2QGWUi7e01fXf4fy4A0fZ1Ty25AFwunaget0z86aVywwMK90/r35vl1Vw/qj
J2eF6fevvlDCX5QH1osN8Ewyap/BDlosxrNmn3VBz6b9zx+5leRgRzkcRFF8CMPh
pIPXZgXxANnpNxHjbHnlwrf5QRMGEhaF1VBJid9g3GGLTXtCvDln8BL7JeRtlBRx
5vYG7lukLdPvqXx6aATLo+eaRSBgtpSdSndqEsGqhoF6FJ4y1FgSF7Hkt0xPXgIB
ck9esCb9o54FRH4Bo8kumE73AlM8qArEMPiUcTqfpxxflyQ1SOHHI6QcbRS5xC2m
ghN9+8RYqDaaUEYWuW66+s3dSoNoWV/l9PBnFRvBJtWMXPFAeTBepi4noTDqYCvz
jDZofr+BHYGBTOgJTlzRMRYCuPYhkhdBTSEVxoChdU1DTCiRQQi5IFBduw256pC9
4b24I0ptesePFYV0dtsilQ4AJ/vmIVl1caTkNLYfM8KWkJ4eTJ2YcBXVzvX60aIv
VKYjiR2qlsoduD3gHHYuCq8jaJqIFOP7UIGkpwFPqMz8z5r3cRiavEPKToF/zGQy
yf/TxTgV2Rf6i5F8yrDup3HQmdGCX/QbvVQhChC09hbrLmQdnI49umpH2IsF8ahB
9ObykAikh6bBn9ktE0h8YbAZSkacFgpmn3F9WT9FhlVt5EmAAaTr7lKjYs7GOufT
qo0K5q/1k8cShsdWYzzqgFlAosoCAwLl9EO8njEza5BHvHTUxNTr2mnM3YhtBNO7
FpaWBUNnYL/xeW1Jvxt05m751Vc3fvykJAuOA2ysK3vN/eSqAi3dIgtj3aTTWihM
P+t6maHo/Ne+SzfEajCT2Yc80DY2NOAlCgOvX9noZwXavVMo5ZgU7pblVqhMHGCQ
faFaVAsX8W2axl0nSeP4t/cXWNqFmgvX0O34KEe/2fhlgTXI2NAMEbHWkLDnsA5Q
9XccPTUax42TMei6b1TSwnd2vQ4PhS6HUAxOOByJtXl8Vt4K9PZ529zXDtWw2XIJ
cE0+wF2opZS1DXvNvYJ8Ce2DLJlSwDX/ifAZRR2bUG9Ur+ixTLyIHLtrsC3HeAJO
FCgBOYZqpKzisPfIvnd2EFoXjIoXaTyhHdyQ3YHkTds97fOYJdMiVIac84yQE5mj
h+40JB4Vmybm9wWm/+wiOhOKU0RPUCWwzRMpiq0SEJcJuQezTJNDuonbF0yLD1sm
8jB9Snl72CnnW80qNxXjOdKHcqgiM7I4zK1fklqDsdHVNZSSCEIA+Y5Oq0lOdQwi
7aEDHfIv8SnJxeTzsSTfKSkYy3PYZOflnePkMrEFRNK1Ijc2kVHdCfxYfgiu+h/3
Difj0QABi1cZ7gp4LE8FbEZfo7EcxAKtplBglsBEnqL2euw0NwWKIHTPqP/W2vZ4
FngoPYnuwnGxVMaU+XqaFS7Er85y+LAkWnbBW1BjkdAIiK+lQvoZyD28JGI1mIYm
LCSyZAX0pZW9J2TT5OUvXsMH5MDn/QfDcGafaqhtxN7QwLlFiyn8O+Ja9f0rrOWn
aQzXFY7UJDOzA6zRptt9m8HrYB8jDX4wsE/HHjAY4bo7WDwqp0RFM/PtdIWm+ii1
1k2sOtdRx5lWWOiEOlf6VrLF4bgSPsTuGq42DH18kw6srwf1NRu5oQwc6neA3zCX
D2LpRbx8W/T7SH+bUBMOM9OsPZEL/JpxjRfACiC3wOm4rB2p2LypYfkt7um4+xDU
PjvpDFJqmCCmq8vtKO/+E1LLLMtEeK5ts6JpwLTuKSrqb6vsSaEJLhlJ5RC7gypR
Uj1jA5XG4XHF2rIQloE5pztnaeFB4jRRqLsauIJNa+gPQ22Ngkkc2ap2YOX+YEAK
XXmCg0rMjv0Wp4RKP1x3hpqfkOKvI3canQhPwg5AWlkApQe+au4FmKUVdVjWMHaY
DOkty9wAoPxXks7WPTvxC77OAHe9oZkyUpdY7+IwTtGkL2CScg1/FCEZvSOgrvZi
08aQ6JEPjIiqYe/DdNheH1x9f5I/I+ZGhM604JFBW3sK3t0n+EHwXGFixC1bmR+Y
k0CCwQwAY9MMsGXXj+a/OK7LmnWsfHzSDePEPyIfIWq4PNngrhN3KdFR0gKuXow2
HI0ed1oRIxA2PHrYS3s3AqkYWKOivfK3dCUQ3rb/ghvuH37hw/2WkqzIse9oiVxv
IXCSPlA0qvBE1QjuwPvEymElz8B6589hG5JDR9igVVyVThp1oBC7rRkewOhL7IOC
3crj331B8VSvtQankVF7+lK2S92ozUJxbdX7Tb4mjKwqnv9q2k4yKUgJU6Ytkqp+
RObmqNXT8WB5qNgILfiLHfpMzGtFp4JvrPq6cVTCB7o5bdfh8Swr2tRn+mi9Et99
YsIpjHn8GPEAlWNfSWgM4PlLnhWWHTKrSfKEGKyRMFIoFIjkL0opyTa0o8eJpfbw
l642uSRus4hMNaZf5oeeKexJzlhq/HcKCwaIaUCnpgs5glkWk0BeZA5dV0ChJjvE
hsO4M3yaelQvmsd1faKDpRL4RCl7Wue4puGLBjkYE5p9Zo5RJkkkbumymFTduCZJ
Qg3+duQuTVdLUhOMqz8nVFeXU0KmtcQ8kpNECjTtEs5fdlw/zeb1rqY6iu1A2HyP
XLKGZFYlukZf8w0nTfPfe6+2PpoHVRVgRF0WXerb2l5F+jlYqsT5NdDWHhpDcs9s
984WhuKXMdF7kdVvKKYFH5pI9xtvxMr36OOm9CNg3xwK65ANQeS5pYTA1U5aYrKS
s1LQ2b7tu17N7/obCm+zmiiXJeXS6amHWXXZmFnV31waGebHg4JbyXqRO82u/YWa
GS5bUnhpAjXhYH9ysw2MC89/VSUw9DnQWfRvdupRamXKhEoBcpRhohC2X71rYxHr
50YDVu/woZZQSXmpLyy0PLJya7vcamEOcsZNjBLFc2AQRQW58P+pn1g1fFST+RQY
BBw4WIwifCvrSIbNa7VjHq5DvDZf9ts8h1d299d2eEo+W1nNhXq42F6PLhi1OW4d
FWa9oB1pzGAXIKTZ1q8QhGczJjCX0m3ZcgF+H+CkBS63FRWyQs0hduihcpKU/qK9
VlCVxKndNNkmr8b5ahwJf2MkUcl8Ihj/RUWcfj2X+Awu7srsLkINXKhXul3zmUSn
MatSUi31/v+5tfQ/xFs+2NhkGXpi0awfogenZsCPr8X0ujSwgHU8glr3QpWbHj8Y
FMizOQRkkP86xA1vGDe2MhG46SXR6IlkL4XlN31rIv+XyOL6y81MHUVWKOg+KXSO
Pu+x/4dk+853WvXlv1ijpgpGsOnkuqv2CXubHjeEc1NnUKfGTHSTy9ojJB4ei3cR
SIzRmnKe/aYneur4aMUyWV/G0jtXxY6LExty/aG6j+DDtyvFvc6V71pd/xx9iFKO
bWg7rRwBAMAP8JJC5jRyINiCTVNmUErpzoN68plNMwfK7TEKDIlWj6gyOI1UBXt9
IQIeLS5pvy5gdqMzc4ifZ3XO6HgvZ1apKb5CcNDmqtyEOn0+vXV3rkSWH5v+Y2V/
7xHhvR+27y1Eb0hS36u0Tvvs/cNtvQe59M2NUppH8OM=
`protect END_PROTECTED
