`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeDOyacUJJyejJeL4Tpy8yZ7AnpfGK93DxYxRGw5Ni/U/SnrWQA851s1sGW61io5
q/uHBTJy3M48PVzyETDZqHNjQHK5JkP9FtKEa5L1Cv9n47kzZAp2CZD/JrDARMsi
srz+RaGZgm6DuHu0nbBL/xibU5E+EwMIW9g34Cm76biKxaic2V+i7mPRe1dFv1vn
4KwE9wpc7502k1ZVPG/7+4Hy3gKN8j1xamc0pLDEqko9ERUnzMA1Z/+9PIxv7eQg
Pc3d4D0e9SaAqTpXYspta643pFib0PSFAR6q+gBTuNlAaVEmOqaBouTI+ENTnv94
WuJkAq/CPXE2MuMgScV+vS8prFum1jGUB77y/xHRjd2osYrUYbroiJycOASfHJ51
ahm9tU0nNKfEpWTjzacYyFM9dPlj50uQ7JzFWq2di5dq1R27KhEFmgQbbbY1YsvT
lQoSRkvtGgPqk39n6awSTW1GCcT26EOJCZuhwWARgSM=
`protect END_PROTECTED
