`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDTddf9v9lsNBcSx62FKQEIeEj9Bp26w1gOdKokjJYny/dGlnf4dIaNiTQUajiX5
vHmr5kV4bTcP5QOmYFfQ29//9VhEuxBVdkTH06R1y2BqFUwUNf+kEg5IFyq5CHm2
BRHxd8PKT7quqDCfn7zgBHZ3JMUovPhS4KkGO1FvorT8dPKPRnte6VAT+UmnWKdm
kBtZY4XPXzsgvJjGaHOpBpJMaRT5rC9pWlqNjCoOsFzYEjL7KltvrceukuF4LxM+
4SvjYAxid86kHPg6PoeiNgv3Prj8KFdQIC84kTw+CYAb+hIsrYnlewu3DIiyfmoP
A48Jdv3jwDcUXSd/+ahQRwjURpVptSkBOxyYYPt3M5b/Iqu//s9hqixcs9zbwc7c
ur4H84A2FNoaJg4dCBfLOb2WeVsEKIf9Rc33eXSv5B26FBZKK74clWUCOwxePuqt
1bk52uH7ZAgHLo2vHpbJI0A90fO4dzx+QFQd17wxVSaQ80efYhP7RUl1cN6v/cgW
B8bnAX7Aw1nN3P1MpBQEvR+9bETobtOVgEIr7geSAAvKFm7UpawAtxpMDyxjn9cT
YkHEUWzwU2dNFj/lc8zZnreCicV+tMl+HiDRFiyQ1J6IVCmmoZo2btKQNE7YRmha
NjgQ/wJgXnl1anw++nHrgJxTkaHRZG8cHn7t2jh7LzGbem7oEbZ7AblMBzXzv51A
2LdGu5VShU4kCgZDfdj1NNDXdfYTWRgohMokc9SrSF/PFGC57takaIsN5nxY/eLe
zZfik4KbJYQ0qfwdiQVi5hyxOsogCqrpyxTtM70xQbJZ5LMI0I8+WInYLenzguMW
pU0VANgg+rraLoq8cQnlRVWRPg7odBFazLj1KmQKE1OljO4bD3nF3A8qzXDpBR3b
Ks6PfiGClwxzuuwZHJkaRJEs3jbuLA5gWFgorDH+YtlOQfVlAOeByqeZp/YM6hIA
9OSsPQ+2tT5/3f1NXSVcS/eBCBvCcfUCfDSLz1lv03pLgn6b0kwM4DcJWdK7JXAE
bNHiVVW4uvJchRLp15nohzqguiMvTunY6NSLx+5qYAX3z69Cfi9rz+gwNkaE5x8w
m9V0C8/onRNiIBZqg0w1ghxKdTQPvZvafW42o32YNx5TTdYg3HP01TXOmp2GIsxb
4qotLpb22D8skKgqK4Ii9IOcOYCQXBdkEfI8VoGHierArLziJT5411+ft6ptbfj1
1LF7lP7PpGhejSXL57cfecUxkN8wYphIRuL8CHpSGMhzBA5eMqp7ZIwm1cdvVDyy
MjzOTjkZBvijIvjtf/6Xaz/cMYXUJXLSLrPJAPfbTRP6VB33+0XX56PcnIa3YQos
XntuixGWFC44Ijpu71af6mzIDMB0gAqeIYpMYfFXrVBwjnYfrpYrsqXvu4pxnh9m
wiMWgkogCIq6y02+fddGy8cM3As3gpLt4f64kINy8kTVl4pekfQ+d5G05nVzSFY3
chLYaR/bN9eE56BVfSSKSpmv7MG85wbqc6k506nhTWFJuAFJrWY1y40naX0NbQrK
EUJAKtbKhRObw/7UzFQEf49grzxGgGj1e7ckJnGCQ/3Lu3BLTidH3MeYYSoWBejh
g5mrbPbkgyeBkMsYfXCcssJrY2RX1r2z1fyrLsgISYzLTIQ7bG+4DlsT8aAPYFUh
2UwJ2FLadqzgzrzpidV+obgDD/G4ykXoAwfIjuQGynJKDHcgNDL+PpyzL8VfJJcz
sV+tdHvee+qgjjWyx2nXv7DoP8/1TmO7LEeWe9iMo5wl+1RpSR14YzQZ5zaDGKY0
SLjLR2R3GEvGr7TpPLGO6NBncGj/wfVwBsJ2m/u8spxWnpDs5K/w6sfMUHwDTxfP
1KjMBd5ipx/dpDsE5a1NppC9xxoII5KG5+kKnFzruuIFfgQBG9lF03KRDLJZ1vgd
77jCgJueXcc7PVUgGYhQYT7nofwWkIfmyvA9NXl8lY3oUwZhThv3JAnYp+/DAfib
mj+axaA2QrHYYwqqJRzN7vjMW8UwsS4aYiFKaTByRCQsQkbabCGHdx76f/hLCt+n
/oqewJFVvLxlv7HqxEAzFUiWKR0wTMnGcrv/ZXOv+Fx++UtgrXKiuh4Bm8J8lFBr
UtkU4v90FDSVlAFYAyQHCxydQvenxG4eCYrTLMFwQAF+UC0hfkLQXvk99QNFMGVo
iz9yqkpUjX0406FaV4A3NpECE6ENdhHkH0qZijzJ62JTSLV/MNQh/oBkscgB2R/4
SBY327J+ZwOA7K1QOuvm4jtPAhCrFGbMg1N2/0cmFgiPuzrPdmxWCib9LHEt/24N
4MvDnYEWfuo86d5czC3CRvu01kCF7XzeDEJs/NJBZkBbaVwF3ojYZ96g1lvQRFvc
2UZ50Dkn6/toQaGWwuf41cZgWH2eTfCNiWM8xi+y10PZkRmmG5Cnf0Wd4g5sEgwN
dTfjJUokAZeD6PR6evBamnkDOqXKTtYB/nrTS4Wdm0bZ3A+ZKFGoaUttukyeqlzD
YPa4i63PXYg0kbo+oAyukKWWNXvQUHvi0FyddGeETqJeDgtd+N+w9H0YwROEsK06
nDu9HeOOyPU5fSwZFg4NnQVfUjxZPFsikH91S6RPId36+yqth8yYMhQ3n4yGTiQM
teRKnC1Z+3nbeGkENVgvvPZRPGSKmHT2S4MrSSoTNoFiWw7DUcEXbpEK8ZmpTyU8
zWZj6249mC7xjtzuhZw8MzO4zA09PHKCPqFr2vORREad63OraSVAkAAIaEZ4FXJQ
bbnJhenVZol8ey6D+GxzGxDh6/w9WAz8F/Hmcic10ILlqxTcTAb2v41bGUD1MguL
`protect END_PROTECTED
