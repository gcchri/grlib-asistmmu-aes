`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/SpVLFOqIVAxQw4ePkiiRk6CeSb+gUH+0xm7hg1JwhNDXceggdoJEwhIFepOXqoT
S67xDxueOLfO8DQNdI0gC6C5HO1nGhl5/xXsTdRHBQ8PW3p3omP1zN9A3xORavQw
NZMAL3vnxlganTizXNILE+flpbKtpaDcEqaVCPPfHpCKwvrAsgxkqbcxQRDqqh9C
DGjuICf1Tr+jhFoBkDwR+f5Ivr9TN5T7/OndFVthPJ4=
`protect END_PROTECTED
