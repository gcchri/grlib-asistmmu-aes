`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
81yQQSsh/ZXlgRNE3jrKcee/irOKm1K2d1nkmb25RnYQ5DXR7Dkj8vV5Utk9X++s
4l0xkuEdaE4HWcY4zmMfwWenpw+0oT8mJST0MRiomCB1MIeBPXZR+X8b7AsZK7ha
QQUzIEApJ/dfILWsSGBeiMJCZ8t5rt4iQmmC1Vbs9iTq59One5B1FQz2Qi3sOq+A
SNsKvdnRwBV/6Pfi0wIim9zPj6AiiASNQwx1wINlJdB3UvO3EuLALQf1MTxJ3T7I
yeuXEAbDahSS9orgjYAhHgcrc68O/DzUnFLbLQhGQX/tkDBljOVOSrqubXxbWojE
W9thjumd8YTrSzM6hBWeuPo29AsH6525BVbfWAeJa8kaKH4pUz8+yNBIER5HpxmD
3U4eFVoPs+1y2e3DZ7F/gmH4FKbHxX3le6VRw9lFN7lJh2mZBfimpGJUVVBUajmh
OQ54qbZTu15X8trAbS1ETrD0MirWi1hQCZIyPnQD6ZyUcf/7Fa1kdgj4xNEOxf8X
l+RZLfFUKhY8BFEePHFLTC4TpAJAosEV117VF8cn409cqd71UeQv8UPBz1rw8vCw
S174ZWJghBBYumIwa8w9O4Eji4MgEsUw1lAOnPA6VAAl8GNgceM4lBg7ab2o0Vfc
3WeYTOwZffYUS+etBpWdAJ57uzhnsi3mJmfLVZgqiWDvSH44yQH8W9zlR8cWj1hH
go7irga7TIUAKM49u/Jg2hFDsqFaUIPPnPJoat/wfX9Hb3ElTUHgCZo2aMPmlw6g
uMorFWiUQVckS3c34tUvoZSCSn4HOsVE0vV58Nhl+ZF6va1I0XpBy9LXAWxSvx8e
0/Fp74jyVfthrFH/IKcLrpaJOpePYIOa/GeN3cFYqSvkuLYOki9z9fkhaSEkvT5Z
CRjBKFS/ZMQqhISxxeL3U3V1hJAG7wJ9Mfha9ZSWVoEDxi4v2PSHY58HsLDH3zPf
ZLViVrig08OTDOuHEobTPuJhouSUTcxCFSTev+hBJlBsqiD3vzQXAfeK1iOfcRw8
eskOzeYtFAQqkrFkYs0ccwnQ9mN70XxEY5SJoz3VnO7aHT1pkfiwh4Po1m4X0fCF
OGuEDjraHhNmFYcxTEQY2r7jJ2QpMbJZrgh7MPwQpoBI7y2AOwXikV6//YRd1bHR
Tr4j0lo7W6Bns/62uBLIshJyjUVVzXZ8diwOTtKEmBxexGUZKdapTKznvZlQdAIN
aUwzYpfP128nAqniqZao4tRgxr/u4pzF9Rboxh1pLqABF8ypn9NqrWeocrI7NQ+n
PHHzQSK3qAZ6OKC1oX+34HYERpPaegQxNavtuwXWtbHR8PZqz4FD6eF+g9JJXsU2
EN2x75ZW5qBmw/DPe/ZDVpc4PsbBSdemHdkMA3MxQ2iqM3dTUzKKGHdf4lwwpNWQ
LOwLTIRTkV6q6GkL/josR8M7NjjFAK4aZKJAtGtpk2qii5O5Iyl499RKE2krtqwa
njtgCUZ2s4Zgp007DDR9B4tOky5RcUhz/DhIwxdM7LhcFXtvLFHOFlJ5BnrSKggX
FUJeWShySOLJbOP8U7UArqLQfe0uI+GjWqcFHXCg9VOeMJsgGivy+siADlSUJKfp
sDAD/abkdOKag4t0ltw8qBRzwNyLXY5GvM0fC3VSToXjezeX04nunncgRK4khCNM
0xdC/RitUCg7at+WE7Ax6gF4Ae7jP5KG+JZkqY9MaByuDFH755ybx4l1ocZ/N/vp
5rGzuqzNKVuZjf0ME5vPay9AjcZhz+nZZ4rLork7NLMwCRp7nck/IoRY6t6n0HeF
35VCje+b2JDcWhTSJIqOjNtkVUK2BZXHpowNIcx5ddkeTO6kkxlnmUs86AocAaW7
f8/s/zgvStletWwgHKhx3OSCDIDqU/4QvdIkLGtnVQrtNDYOIBpZYgEYL+k9V7GE
xXYyBxP1Vszs/xQg3BfduXLe4z183qlI0NRiQXq+5kgtQOB9Q+i6N0ye4qHvk4bq
ps3IYG5Wv0lczkVlozZ+7mpYzCgGgqa5Dwrj5Y4sTg6HmjaCfIp+pElCPFlklXI/
26k5Ose7m7cHMwlhUHIohZsjTSbGJs3CWETyuVMQFcyaJbldD5FRccEDMI4sGbdn
yPdhXwfwKjTX85eGWxZS6I40XtXPb86bNQYpPJD7SALlqg7BtcKySWx9D5M4Wu6r
8bcmasRBDYq5K7RD1dly78oe5Z5bdMiHyAQKQICGXQ7mNDqepiG1vpFGXDNjKGP3
SEqAJEXUwGwk65YLom0WzrJ79b45E6efz0IKBlJM4gN3jNIKW+S/O1mK4IKPVLQ5
PYoFlx9UXJYOvJorfazwA5Cbl6jOby6MXV454sqbJmJvW3F991PIlDwFrX/BykGB
E4nd0HaHKswIbfmlgezMdGyNpNPs7v+qI2ebQAxQ3iKCBoLXNLrPnXriqPIBTiyW
DoTbeNPrqhvAw0W2Bzfas1byslpEC+Q1yhy/Nxj4lv0R978Z4YcJKVeQxGZeMEjA
Ek09/D7AG2ZCHWhXqCOm5EaWgzcpqrexeTeNc1ARnj8QFDFW1iR86ZDtGLBCrN9+
6C4PVDggno8zIDM3TCNRjCFG/2F82IzriTI4sPw1FJEaplNr8WJrUCCSTXyoLfUS
GG2URrKeZJ10qhQs4ApfBfK32tv08SugU4MK2tOGZ38ccHq3B2ag5hjozvAM913g
SjU0PylsqLMHu1ZfndIfdm5mW0wqV46lVFJWwhTW5kHJC5E2oRWWNqr+Vj+BHKgl
VxuJ4nzzM33+s1dfZOQ1QdDIpFo79aZpuo5irszj+8KmNyGQ3Cp859GUGOm/Ep3q
ssiYWyn16muTHbWMDFjjcUwGWWkLc9eZXmMpATphoUvRyzzKJgdrtxdPVTvccfi8
FVc8hKeBH2C9UDvGsOF2RS64/mc4pwkYMkoLAmpr05zNZwULcx03rXwer1gBmB0q
N+BnKAXI0E7b2Hr0WSHvJkBS2yPuk2EnMMQ9KgmKuCks3LcZ0TPNLgRYOONachxI
roNmihKbk/8gvWWeht00bqTINOkazFiDh7UYNOUq7istf33GJtbbV0EyCyGar0at
mlKjJa3epP2ponmfHFWHhnq3bmegtQlgwQtAcuVqIjx6d1gceomJLz2NhNCtaVfC
d7K2X++ikPOmKx6L0eOQwdxwFcKhee5ZxzkIDSWnwtD8bpXiFqPer6kcwwNKdkc/
UM8XR1VKWnsIs15sZtv5mBMTXt8S7SKnwk+zoxUlnXZENHdFtyOcQwMyYMqPU7NV
Jwu3Kix96+EbsS+yo1FZz8stRyKTWFgqqvCELIEFKUD2l7cJhXZXh5mpDveC36SC
HOjWk360b2E7HC57NXgV3p9gg0iJS9AiP7DVPWyXl47YdsNYO7HzEP87eNACLKQR
ksMYetHjWKesaW09xx8WIsl16l0zNdOqcOe5rwyWwDqqRZtl9PB/wg4Kj5RM798z
JHCcH4Mf/ezdo5DIH2jexgYkZP5aBny9lU5KbMwxmGZIQe5Z9RtmOlurm9xqMA7I
uETxaAD6Ov632/O2A1x6sJVPol1p6aUtLNtLwbV65nbyFfnTPeNx20giKngDqmtj
enxEVNkE8khkn2Ir3dOmCscsa6DjSM+Q4vAxLaOAL8uPKdrn7LKrNRyHxmjrFyw5
GmOVAkQJlaEE3HirxWPTHdFJ2B1PX5e9Kv5jWm9yOa9P71o8+iTxG4xfwuvFCbu1
Q0/Sj8jeK5BvDTlzksAYmvXT5gTuJwqUEJQ/Hwya1Skg5vQr+A15nPyH4bqdYcG/
MCzuOlFDL2bnQPrT7//hApmmNYFUUpITVFBj0nEpF3XneS6zozZEy+tRo1HnBHJG
7f8VtlWBu9TKyQKjLFLpK2wp3HwqFTwPvNOnsYpCXKXluRycF2K3bA5rTboJGhcU
ySqisKqulIc5qNxNBUFp2lCpnn6u7iJRXAG+v08nfGvUM9gAXPDfPX05+hWYOtzV
IF6oLvhrMnqBiC4i/KbnLAb92s6g+VbgSEv2dY2Nor3Ds9QHgS3lDui0lNNoNQ/n
ujMGUeBHfC/x/opqcw3URvRG3wJvmV48EphLUaAWa6IZbvcIVRHFJKTcOBOZnuR5
BnVh9EC5hfAf4z15+V4WUyIk81v1msgMJHbfteEDfyLsr0WDa7HyIyDTwmSoY3dG
vAnxIa/ZALNTezV1kIJ4l8Z+PdkZRZuOzkGRU1Qh3OILY666rsPkwGodR36LP8cw
ZeW1/4NuacZaLeUcKzgapg0g5zLh96WR9ukRziAlHzOhv9oS3jzSBN89XCXTpkBM
VtTCQFDUr7XwADYOF/xj1iQ8SpFIANXQmznZAekdjt46dgsMeBAJeZVwBLYnQS2i
TBJeXgXTM32MLypgrEv/a3Yx1oy4WBjTFc2uAsuUjk+lCBr2PT6w17f9uL16xpj2
E5WlvMK11RuvjPyh4/o7d6RN0cFaDvpN3yuRuxE3nQJ9m8/bJb3X6LIqAj1utZdk
0opPz4Muf4MlxoQukW7D+oxnEApNtbyKFRazS+sAnJ0hPRbwOj+YkdboVsnDVJxJ
g+ThwUJlpBUMjX8FnsgM2WRBGi9Zl3aFfU1ceQ4rYbQBdWQXnLBMgqpwIlmWLTrn
W2wPWRmGYk6x8YB3Yn2RnS+uof5Iz+0Ppr9ThkGntkjeEcNsY2DcnQxgqfMAY1I1
gCdrT4tPC731MJW/MksxFNeXltW2nZZPq/PN0EaJvjJsCkOPq+MYBE9jCJ5DMpAz
E1TwukPljZ4wMX5bRhgYz6M1ZSfY1TY0NDxmLV0kR7DIz7QNEVl63cDSJOGYDOYS
xa/eNQCLecqDgBFAoBs/4Fbha6HHZL1XpGU3ZSmlwtwpRlpL/g52TKpURetK/QaE
jEU/JwXiWVSGPIbYdf1qZa+AgoIFVW4DC/9zqvggpM3VHzLVrBSmXVnyqYd9qsww
dhjUNlI1CmQqwLWbCevRJI+Z8eCSIbbCd/o4wwdyhna/8N5uojtjzMDdmWMQhJ8j
lGj+JjybBSPTdwA4BN3/4CzrLjD1A/l6BfTYDOEIcF7EZdOSxLRxdY7BqQGYbbhQ
Niimcs87rc2G306+fSAelvQ4+uCDKr46mmInjYL1YZTuAqOP4CilL+ozQhbLwUaV
QR/TQK/+ZUj68DpaNckPKkhiBxhxcT4jyhk6U+LAmtCrYs7Au9sqt/XC6ijome1X
WSyTpYdjIpOXws7zYmwPj3q7Hupp3uhrTnceUTGo/PyaLay81h9gm5Ye1vWQLkKL
d+UGEom6eTJKLUhXLeeX8giVC/hNZUmNTLo6qTgE/D64UdLHKUGfTL7eO19NYXw6
wYAP99cPb0GofvfEr1F4ztS76MNyD3wSQ+EN+F9zeKLrf0Y413mAw1wmukahbhPD
sGULylzgfLnOshVHtdR+U2X6ajRj+NeIgayFfedwoD9u3AFUIrtl8VeS99e8SqCb
6RkDTnVcGPzlLCE22da57FlIOde924NL10Zm9yiXp9XWhpji4iZeYzyjZg2qnTl2
TNGtQ+w755jUOoPbFhW9x+RjB8LzVR5UArGPL3ltt8o6kkn01QPteM/JUbDxeggC
3TRA3smvfvTMTh0fa/k9gPD/ObAtQBeW7iyk9qq89KUxsgevqBURmRqa6DK4CV+E
H28rg9VAuFMN3YkmbUQ9EBZNotohT0chZgPnoK8pRU2ERkMTP4dA1QixtQgZzQ62
F0ppA+Zp2mqNwPVLVGqXLAGAj85CMi7c6BGE40dQwWmuC7OXhCnvfyQZIHpFaz87
8K98bMNRAO1aP0tx7TjVAchEExOphzNbCQce0T9cedWesplcqgXP1Qd1HsZB1X2R
BY6wkliey0ablC2/sHD9Tm02qMPS7ynZSMU5k6JMwWTm5aQcZ8hvhF6w0xmwFpve
mjXc3M78LFuIB56UhOhei2mnI+k5Mprs0LtonlEcZ7U=
`protect END_PROTECTED
