`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OMhy2bADT1/SGcQJFlRVvtJK78uvcn7m+bYeayXR1iX7Ib+PtxkRS/54A8nbV72c
Ad17V1DuiNcxftwXexThnTf5OHZ8BO3lo2iP/whrItsJq6UC5gb/C1nvzvQY472O
s8hUZyA1CSfgvMIPy8+fFdhwtM6UF4KY4RJlkIuWi6H8jzbDOOo/4aMJc27Mlus/
78DbzmRXyIp3ecbZNj2GzSPuTT3laxsRAO6e66JzJ9jx4x8oLrNHb0mjSyvAflVl
UUvaYsGLCdDb0pGQ6Ue39cPDC6n0tEt+wYR1d94UMwxKtUWL/nxc7ZLJZuFQNBrD
0oMma7KaApzjU/6LIWOw2qpz+Y84gBdTKQ55JDwWX/d5Z/OQpMwWEv2S9n+ww3yX
RzySTi6NbppdlHWVPcR9kUNNvDC7rLDZfwrzkpzO4JTF5eWThIY9ALw+jqjUG4vI
EHrc4MFO9AweHbGfpEjRw3P9iQFxvoCW2VNIGAQRash/1LQx6s9nr5HAL6hJz95a
dnbLwlzF9awI+Pk4u6U68kD53LM6f+Kq0OqttK7LHDkdNDmJuEvC2qqvIN0cEZBt
lxDtpDa2hW1rZXLwdURuPMOM7GZMTDQlT6lmE0ie40bVK8b/e0xmy1YPSkgY5chH
jO6N1g5DO47HJfq2rIIMqrDZszQ/yeB2zYpPfsgQnfU=
`protect END_PROTECTED
