`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9lt5XZLBn2ITH1Db5CcN/Cp27d48CxN+hH6iJmpaefQtYQq3+J0Q3ZloiUHM0Nvt
OXEXsL5ss1pwIoTilFCS2FezqqYpMV7q9W+y5xrcy4jTP1Gh2YLEzF+/AabQFWov
B1a/iCncFCtr1G6/ePFeekWEKHgpdfUMzqpFz+KwaQ0ukCW46V6ykuoMf+Az8C4C
Bep0rl98QNiOUutmQWsV2Oyc4y7PlCL0UDJ3tTOPAMj0jsEw1Oq+EPjPzJQd9ac/
fS3213OK6bKDj4xvWGCFqsoQmvAubTHUekKxrdnl+SuPLw6Uu8EB8zbbhxZrmmCP
pJZpOlYiq70+M7g/n0e2+hDJfrYaVjAcMJpDfRnT9IpF4FpEZsKupP1eeU5VX2IB
z6xNhR1PnmAKWUFU8Kjs7kQFmC5cOpPLBHoVWjMsxulEieSzIfBx383u1qUZmHHB
CCPLxLWxve46xF8He8PcPoCivKz5JeMGjaZMBvWupb2yN5EOra8M4NErZyFJcRFl
epuD4UoZlqmZO+UPxjqZmSf6LbE6CXsGAqvzBEEoy6Mcg97HtTAl0Us8kzMgiopI
eMLUFt3AYpuEH5WmzlVcu9X4guzp3/0206qczhIlexPoICfTCANIXfP61p6vUz2l
wyHJemrXMKUM5AW9sK7LyS44gXAhq5oxpVLPHfhcw61NEITnibHgW0P1kPxacxLV
/1enIfpqQbADqN6UAVFIV5AAtm4eKDLPW+4SL4sbow7h4ZW5oCdDM8jlUcEKv1K/
Gfub0zGTLFUZykkhnJY7ag==
`protect END_PROTECTED
