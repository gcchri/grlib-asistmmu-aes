`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRccP00gUgEkiHRXjypgAXxBsvFxHCN87yR0deXt/jTKFFwiaK5GkOYxuVWd/2uq
hUzJny/5LdeaGnkZDwzsKeS6N9ichBqYRDdgGJ8gLnYf+ASbXvJihmvUQ95bJrMo
sZveJgkDFkPZk6x31vqEC4GPJ+ewW5iN9EO6imp3upqmrdfzN7d+iylZbTYNm6xT
dMuzPSWDsgAN9uanHdjQtpk3OrM/zxS34tQkB/hUkoVi7ojuwlo867cqZH4QA2+0
5KMQwmFWPgojjKmVQ5aEyuhkfMRl3LBX6/WDcdui4oE82qTOaogriqbEARxBO33i
qtjJNUOwJDNtVqhGD6PoZb48/aLn0JHHTrjS4SrL2fHM2UHBtIlusUqt5IretM+S
fnS15+RmyjBAbz1S8JQVqk0S7Pfz33yWSfzhFoWHOx9/t2I5p16YroBdXgDRWg5J
`protect END_PROTECTED
