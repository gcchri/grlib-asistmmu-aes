`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78ACs5m4pyP5NG0/HR48cSzBF8wbunlymmCyPyyqJ725JvZjUAulr3y/yQr7sARQ
u95swS9qPqOSwravL83wajsDuqaHGxzGPcC3woWLnQLucMnvDXWRZrVa7ovz1qgx
ciH8sXUIgnAv/ITjjCzeFITUu4AXAZmmccY3OXnFyfvSQjcn69fJ/s7qWjw2hc1T
XpC4Ny1y4uObZkUAjhflORFvGuBm6H/z+AlEwpxZDmikQupHVC1TpNFDybgAFDvR
kyck0knrBkEKgUn2RKNmozyZ8l/EqHY7VAunT7WNYLWVxIXx/xx4M2ZiPVzGdRXm
XN6J3yjfEr96O9c+7YMZ7dhhOX3PHlGRdXoW5WUmn9hlFgJ6Gxr2kQ/91NG7JM18
NOVa9+Uiy1nnNEYS0VdMrRWz/6MNWMJ+KVAfbqcunx/nC9vXX5cp5G9gHXuWKCXQ
Ml6AC8zNHYLk1eVEMQhYa6iGxAM4RJdWE9jLoYa42Lg4tnoqHtv9nYre5x8m9qP5
`protect END_PROTECTED
