`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7j4vxuu6qIgJTbDlb0NmMFd/FN2XFRdpKkkLCcvKfOiadTt3eIRQuy8O2O+3DTmc
tbtjZkkCGMJggB0A6g3lfX5JXSHqDmTTqzUPDsjxtN4xehRsoW/w49PpfKgMr7ss
oR4cR6xe5kRUTmmn3G84d7heYtwzHoIS2bSlbA4s8PZavUuKi63YeFWxb6I+Px+N
j677jiCLuNLlQmQDleTQhOBPxZgTnKtrIlZI1Kc3oOWoA5Vq2qHBMh0VJZotQXWk
4X5ucUo6ogULgumV0u0h2Kt6hD0UAMPV2o65N15ald1yblwJKgrqvLHo0PiQ/WTO
5bdvdTGgiKAYlrxKlptgUfF3JoZK5YTtnF4y16BBlL8MPwGvftfti+Dc8HR4lph2
r8HAnhzov1Vvd8z0SfSdr6jtazHJTPPD26v9TK732qn0Ca3+XBbXedW5KFz+hFWp
1C5OITwNMgQjhf8wKYEI0cOSqUZEW6nvBquSnrj0Sv2JkM512SmACZhYkSBsNbWj
dodxlu8rLsoeauotjIqtBgwb3pPq9K6ASVqo0sGW1QWkHVh0A5wla5OZ9wZ/32bk
UxjiombF2oI4TYlP+yqcZSdj2OxL7ghBqMoYf8ujsO6SSmWmVOwJqZRoKtTqPlve
/PBBg34Qx4pMhVnCO2kT2g==
`protect END_PROTECTED
