`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5FTP4XMPApUQtdQ7qQRIHwrjhdWykG0JgNIvhOcGqQJQesosOtXakKbcziOV/tki
SdfaP1omhhGbUn5ohVmgdYWVLVksv2WkWhMYwxLs1OybauIb9dgPimprm2UDmMBU
gaf/H1Z7XlJtAgIOduWJmqNDPxhvODqoCJgXt7dYwcY6eVFsanP9r8t1U4fGFUDg
0UqP1mVZceDFurPdxEqU3/ZcnDpIVTIZBMEy0zYmgzjA8qi4Yhe86OYTOYKxXXP9
frn/On6j0wFsp8Xv84760oTV3RcYUWvqtkiuiucdJ4wgdLqCc8La0Vlttgfe18HA
JnQmYEJ08I9JkjGQfAw1cJZPMkML/1/svFXIVLEGcH6H093WaY9Utrld/gA5LZOH
zHB6r5Y6rEafSRWqs3wFvya9NXNDmD5nQhlDw/qF8kXgWHuoF7g1W3mYwn4pqLVX
iuSrhWQcMIDvhZTfnIIlmVd5TWvmPxi28xOLgV5eOxBzm1qokDSMFIypmmTcNRuv
kIIB18YvxmK4Zv7JP5LuVkoV79lqnS3ClcMtkvLfoBwcZsRpKz3K+ScnE/A58hNY
IJ96wBdOqrp2AvuD8D12jVQZ3vKpnXLAF8Ycdad16AN6sc3JyKepu/G1/K+0dsf7
shNCOujwmUUr9g12knWteEtfnXOg75otg8vHWq1UN8rI31n8Tg3Oqr+vf35kuuqN
uteAXkey2HX4HGDGH9slf6CIKHDGVaLeNlYkQC+lVaVhvLsEyaNp90e83FE7Y2Be
85/Vc924QIBrTwJmEoCUlw==
`protect END_PROTECTED
