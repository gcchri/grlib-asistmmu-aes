`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3wtPShsDnU98VxpsAS8alQNJdRMhjZ+lGhdSlGqW1um/LsvdWj8gOE2F1/4+Kny6
HzkDW9Iue//X0sNEAy3QO8lyFCAE7IVSoTcisAAMcKlGqaQsHoOeGJdGNTBBe51B
0b2SzfP9rvD1jrvgOvYbrX5DQHpcMeIuZOXCDEfocjvtdITdev84cdG1mXpeRwoj
VpRbHMYOBw8TU6rM7hnctg==
`protect END_PROTECTED
