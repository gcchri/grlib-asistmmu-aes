`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHVfelxADTEj3huA9DBhfHJ91oG62Vv4VXmn2x1aeFkytO0gLgpyDnEalGg5noXG
FFNFth6vOeEFQz/IeswKW95F0xRYf23DPAnYIM3lsf1YrElsz38/04y3CtUBmQsY
5o7CKL6ZbhGd2Z5hHepIxtI/yZEjUxA41STxEJwjeXrpci1T/pMCSLdtqvnjcSbP
aY2ZCODgUzjLXQgCn6bhMzgV/sF8oogoGSV+NqDujLN5uWEQWCV/rmGOTGBcvBFO
1msj2uEXidB8Vc1nZ0RtVhuoQC/Po7RDX+Tprm21d0HPgh3ei+Pnu/dp1PQTy1S5
nv+AT1lorOmP3GSBMa+WOGEz2rws2d91OXTpXEtMuHsiD2U96YlTumjjbDEvpjYe
HbJNTMjqS1ICdZrD8v6Eo6xOQumE9kg61isFeAaLpRk8Jm4/1dUpfrOs1TrkVN60
9FVh/xXdziibKM2k/sSqeRM6Pz9spKyzDTda9IHMJB1umcBEvWGM+zMtopkIiWzG
8KmSxB/PJMkd0TXaw/3PG1MKfX4l987IapDW2Ilvq4W7R2+o5pV9CGl4XW7Vyt5U
+7nasjzRE5tyWynMkKuIbQ==
`protect END_PROTECTED
