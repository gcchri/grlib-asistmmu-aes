`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWOFHOV855azQGbE7hJ9clJj1DEu1zQc5cbc+3JlW5gwPgZO2y0u2/TwvqQER0kn
TPJ8JuJXGYdKc+i9yUMKX7LbGPPlWD1qMNrzgv0KWqJ1XyrJ6vOSMGp9WCuagcie
mRs5xDYgg/NqIBPPz0RkjKjskIhyChQmnhGet8vR8ScoLBEESyq6uavUEyCl0mp5
Kr5xDNuPNW+UPY+MCn9018D4F0zC6U7Pzlpg6edo1d3ifmKTKvie8zmDIvNwxror
NPJ9XrQ2TbUL8waz4CQath15xsHcANr6nuhneY6KZt8/HDXFk356UjYB8rt3pfih
u80Viwyd8UloW+Nnvp2xRr4bOpArUOmhCbRY71PygVFX5I8WfzBw48bbTe91lH/i
Tz42XXIaJyYIymA4FgFi+aaMmO4UhGCoAZQuIRlNHf/wW+N63smapE8Oy7Z7DJmr
h10wed2RJFPDe8FeK2eqMyswbHpk97oNcWJwoBMA0ieYeKif6273jBQPKHgCOt1R
Q536hf9/64c8ulIFnYKY5NtHmLfBQFCebrOz0hDdvqUeiOJjFn6t0yy+PJBDTNxn
2TvxglmyKKjK3qX6O++NtzIVvt+7CABydTHRKjnBXSROKdB6Ffj4LtCQK4vrVaei
VsT+RqS1YW8Cg26pngRlivkQ1fsL4hPDF1CcEhyKn70b9w9XQesGbsMB3LcOsdpo
++NOzTuc4w5caQsYhsi1hjeYjOqP7sGdfEWD0Tp7scQS+9BT24eh646QYSOyf9Sz
G9dsE1ouoRKRX9I8dDAZHfAfmhOJ/UACmXbecsJfIJCMlrWX4rAXhGCyJFOdNf7W
6XvC51dGPDFUjg3bq6AVu/MzH+WCWhqjkOcgeI3HYFstU1j4U7z0//RtIG2NVQs8
JJxf/GywGqaaE0xYzHir0aju9+DyxC3dWvWI4ZBMAixGK3351VgplrpjGxHxkUMf
wvLbq7F3T9Q/kIOaqYsReMTndZRPHWGyvmdfN4PSYdLkZQOKd1MXKOd93PEPOTvF
NCdC4PJyFXULrBc9mpKWrMTqxMmvj4Joy1kIyx34+67d0fMLW2Y/ZHDNlg3FsSJd
cUhcpu2ZCI0tz26ejqLFl6gAthH3jZo7Q1bRyqhT8iXh3Vi8K5Kr5vQCZ9AeXLIC
yScFdcW6kiAIrkQV6rpfSPKUS3HvqVpDKkbbftWG4TGwV5HZEmSkP5n6BUZv/I6j
Y3r4u5+PoIUfztKIOx0ehBTml05I779oBLbWXsW07jB8RSZLYdNCMaf8lviFU3dO
V94n+lRVYTKwt7U+YODtZ5RkKNKayVVo2JPgowzqEW8=
`protect END_PROTECTED
