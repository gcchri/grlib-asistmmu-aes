`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06Y4zSyerXcuRxbh+jKTKAGXmm4EWJoe+D/0uvtymH16G/qB2XyaXlpAeSQUiLI0
NPlVawyCxha0k5/8I678e3R9tg7Vb7cRQzkyH3xD5A45QUNgSyulvm4ypih8iVP0
TIUsMKFYzq2RGEv70rOM5/eE8yjKvzMN8YxdYWu+RFaeZx4cWEIM2VHxScvhJ4Vt
4njUyYzhHNhzezuNAupcXyncFr34oe7i9L6MiYjqwZn3Ej2/uUMoay0wCWY/KPZq
1WPvZTUg05p7RXA2iadKvXyzHyULYNI4yJNqImwoHnu7ssuijZSv0veH+xvy6Cr7
`protect END_PROTECTED
