`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWOWGiLYuDAc/cIfjdQPpH6PKgrzHQJUlNvCjYhorTW0HXKCCUlkEGlks+a1Vdd7
ochnLbQ0u3/EKlTAKWSdVZyxzZv89Sh4IiadGY5DCRALXT/nAtNxMCoPdKqneGDN
CwDE/FR6eMw/MCHafJNg4gzMIAkyHcd3qLGZ5mZsA212eUfNwrQ9jNLV97AD9VSc
BDM5yvVEBXxa4ocHv3kJLiNr5um4NKQu1GPTRWn1ZMhJfH+n90MBXN96dIcXB+hB
TUzlj2i26R/0rb3FIcW4/E+8Sspog/y3itkRA7dGXmFsWcztQyVEB0F41C74Zubs
RfeKC0W5UoW5YAsQZB5c2dj4tptV2Md2igKvwAyVOaLBQFLofWDIKks3/oBthjQs
`protect END_PROTECTED
