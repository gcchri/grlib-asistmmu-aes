`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k5JJx+TGcrKRc9EEuwl7cQRvaIPCF5f2KSdE6pCf+Tv3p331KedAZBHmtGhZvP5W
+SFDp80Me4vzn60FQAJvLWrCczkfK8QGbQJfSLVP67TS4ojHLsTNTaQp/DlaAZ06
ukS2w5k0b0MO8p1VSlJK8LgWs1x7LyNdDa+OZwRQDzJeStbGuunyNWAfbWRGqyAd
hK4tM3y1pQQ1mAXR16yPYB82uapnOsdyeOyXP8JBFOC96kl4h1TFCP0BpLZ+VKmp
WxroNrdqiSo5Ufhv22h/H2/T4KeDxhYEPFTN7q3zgyijBop9hI6t1QMjUoZJQiJk
rvXmJhoXd3rOBmhCFiVxowvVun/3tm+QvEMAPKXqHk66SRH5HjK/G1L4KeLkE5hl
5U6YnVjidcvBnPKVeokzCAGisonVtIzf7mnIbhfaZFTtLcGIvc95L6f40uLiC21P
`protect END_PROTECTED
