`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2S/um9NQFPCFgryFPkdxrhD3g/ShW++vVuG88s3OPtrZh8+SA2iauFtXiLu62qN
gquTeoyKpwvdzQp1B1RVJ2qEPa8+T2cGuwRn4Izz+YfQJDvFGcqFgoGvAdWenVD8
G92Ji53M02UiLRYYBkttDtRi+EZuSVu7kw1AvNQ0FnLAhUo4/J5F1BbA+wtRta+c
/pyGTLs9WlxXr+VEFN8McJo9o/d6tYRnJwLBMTHRVVbPTb+LNlFL5IF9IRk/aSQK
9PmYyNTiLQXzZYi+p1AQxK0lVrvhcW7w+wd7V5vOiiS4iM8rqJbCBMbxTpPz2pz+
Me5jt4jUsYAUWrPwCE+p6h/6Eu8r59x1cKtFEQaG3wZkPhQt/yPrg4snUeyF3Czp
/rr1PU7x1RQ96F2ODl7uhDKJdKg6I5hcMhiOWD+kjEs=
`protect END_PROTECTED
