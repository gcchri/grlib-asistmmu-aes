`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0JENTeYjQJbGe6pjejBA/jZ0joMfLduRfUB5d+KPghZN9HAUl/WKLxyrUGXysLKB
7/FxHLCWK1g3swqNxBppvEB33S/q8I8rx3/KqQEH+TRyqushIi1C4T9ZTsxD0rhY
6i8xB0ODyALTu9TBTtTaKNrulHp35qy/FRVzSQ0/9y0IIzceE7zKsZVPLBFLQrJ0
d0TgQ88cDoddul8y1NiD+/qmSLR5OToVpDNdOCgKj88rq6Dafxar8JfzXmDEzW8w
YTfn/mal6uxB2z5SGroAoJBX4PF3qodTntQQW9ccZSmCJqj1dnh4pGsqxXiReON5
WJxKv+T7NW0A6v0dHJsmF+IXO1MyFMbV+5oqA+BDFjmvQVNHNCk+AjIU2L8EriAM
igNO6EWks/iXobZGAwJ/bg==
`protect END_PROTECTED
