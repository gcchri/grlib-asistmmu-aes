`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e0Zv/m+aobUZjq5I3dJ65ud3Z4d7Vng9c0rFxJa5619V5ihXg5Ope03rgJO5eazy
J2WZa1hCaKIrvbHtbBQ0qXD/OeIrSxIb0VSDJHQqIhJggoL5oUtOLqo2f9KjMb3k
t9wujur12U0gXPQbdKumbur++EpZY/GaAWqiSLcsVdCN9o9gMxonhLExTaIhp3Xu
EKIxlZg50HDHRTdhLaaGqiHXb9sMww0jyLEa/k/tKBxhFANRV8IpFPWxZvMEUDth
ZEVszel7O2P3f2cuEkD4yOPWdYWtZnAQ1vw2XzzrFnmsyyNhcxRjShtKkKvooO/B
q1cwKUBeWPgkeER/AI09MZfhgwpdF69vPVtwHlxhzaTdNYqgKcKqas4eU5mOppGK
JmQTOKXOg7Vq/fOSx++rhPt6R/l5ERpDwWOk7r5ckE3TZ8nzF1cBdQB+es0Y+Myc
`protect END_PROTECTED
