`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZF3w1ook5AlhvaW1Ln2NGaW4aHYS001R9vZHKJXtnn6tYYh4wttptzctXWyzdPAn
UcdrS3vVaesNYCMQ627Mvw/I5lm7rlMaqpL1UmgL+rZ4kntb3oZwAFQPc/kb8E/m
coEEtV5K/IfWdFPJzB/hW282zNvpjrzcHReMj97Kbce2jgzA1+nUEzl6FICWWjGz
dl5W5yNfTTIdBogMsip7LPz+rbsi8nmHR7mHNcVp1Rzv84BfMVfU//jl6qQUwY1x
2QYz0dAsvfrVjL8R1YEyau05y5n7HeiEnZbYelX2AzzQmcjSDQZBkA5gARYido7n
KPCztocjA04J/nzh5iEtQ9j4Hu6u7elumBlnkSb3Xttm1jEtq4jQi7AdOyn4mEjX
lbbbx5momLrrmMvVcz6fsSon1wqXM904jfI7Y53IWOCsiKuc45BaNUzON62SzvxI
E4Glwla+4Vqedw5VMGlHCvkbY2FsAQwslhO6lqRr8R7AtbvOnnOSwl6A/BmbYUCG
S9cfAcAkkxruwNLB6SNB8ZiFD1wQBFftvEkfFr0eYu/Ha2n58VUAP4K8dW7CicBP
7zLqvxiTrHkNyENCBbbBI0y28CB68uWZUEz9aU8UxU1jMWqkUsQAA8gp8opKk86G
IXFA9GoKzcCrzuBJH5s0hGn1//S9gmQBvD2PYFmbTHFuWT89qhdFOiIPAQt36hg6
WqVHrpYoxpsL0HN0e76Zq/7bxPLb2JJKS9DnklN4FNhb7jKlN8/R0PktsRwSfrS6
qAjxJ4Os+YP37uby+/4Q6yABhNVRJwbh96QUpnyXdlFalxJ4dQ3uNVf7dnGA0bPS
ZR1UEEyD9oearsygh3cRbBRTTUYTqZoYhKZUsd4rH0X63SWYTvAoLs4LuW1dNfqD
xp3OadYzOFsTLX41R4tRM+pzuXFvpMTfYfbyvPlNUrBfcAyoEgZMn7Ag9UF0c2n7
aHJhzrJNZAaJR6by3Bwv33hLKMpYqe0Kj+/EIWGT4W9Lr/+j/swAU0tFs/iBCScH
4ieBWTtTL6KAKwOsfxQWiqHR6V0WMxioMZz9B4WTEnziN0863E7i9SSwEp1Fagl2
yldaI7WmvoEyZnbTMPAiLQLaZ84jia7RyyJ6pBPk8wmOzuMdRVP4yFoOBtEJ8rUN
3vUvPOcS1g4K77Pw5cxdP+8nRh8jT80ESV8Rtx2lHMZCmzctIsTJTjk5tHvK7YXM
Hs/dRyl2wJfZE+uwOK6AktYNpnMosyINIS4lcX58l0iTw1ecgDgEScHqQRoIVWOw
8pW8plSQBkQqrzzKom1zQNe1G0wHRCX7Uqt3w2XEV4DfPpTxXHfufBpePQriD7oO
7DmxR+1Gk+6jMUsL+cAVsNuIekJ9mT+BiPAMf8wQrc211iYpCI+C+fueepJMwLcQ
TS1SzFoHFihEzS2WndK7Pw==
`protect END_PROTECTED
