`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODZHnuTFXIL4DtIJbQZMSb+2XdieDbRZKTXfHBPCvs5n7EMJDd13vbxKCb2UDvqt
sm/B3uMlReqBuL5HSf7lIRYTiOtL2ALEwPMy51t28O/xmpLoXvfEpaBc9mbsaOGB
jB7fZBjODJTVPqHdCPCYvuKF21aGeol8vsbV4IwOtbxsC3hw6XU1pp8lleNgOFN8
TU4hlV6XnSjqmAm5fcauFJFFFrDK1jk7a1fAoBaQ8foAjPLVUZuH6W1gwNpasjb7
L0j4Ss88TBc9ZgOvza+QmT5UDSjJbMl6FZXWVeCBM1FgdLXI5OhRtD6K7LL6nGag
uYlv5URgk/gZxbvyj4OSp+4KJax08cH1ob668AGqAhzN4Vh05aaQbS+StBf2kW7j
kwZT1FNb+7H4Xn68+W74iON2VOEWjQjCxyUxfQVQXg3Y8NLv9K06+1ABYCExKREH
p0D47sWsnPRg1kxvCKRLPg==
`protect END_PROTECTED
