`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JEUwDUo1QqeKDfjRHPryYaxL4w8Uqv4kgECHU+UewVegzXm6B3T0hQKHccA3Hz77
ONpECUNF47nw5zJf0Q/xeU2gzwYklu+gs0kCQoiOHbygb9Wr+wqQOkiUUcWMgs/n
+BWpcCXu0GAZe6u2yrTmFMhZgHptHunRWrSb9uJa4zk8Cold/YxKdnw/U3XCWftg
VxHJkGPvvxHJ4W7nxa1lPgtTHCuzLKXnyYqhi+PaWEhspjFF25FdyrGomNjmFM0V
9//Zi7Qgo2xf96VgZ2b3eBXPOIW4G9kDS3k+QWXoJ58tbFXOM/8ubapToABUkavB
p1lu/AR3ksGKcjb+rkMz1YVikaCquG0x9cvtthmywnz3Te5tpA7KnUo2oULQNrcF
chEzvqi+dNxQGXLd88nhDbwBEv6IpLFdX7GnVKWFr5iO7EQL1y7puXR47y1tcAN0
yLq7dg3rf/mgzKx01BHdOsNI80VJJj9ehcYEOOGTG2lnLny18dI+xAhrXnopiLW1
Nv6fas+SUsDdi86yfB17LrWhGDJVQiP19WtIEdZfucwGflvg8zrSlq/6Uw0Q5DTG
ZigRyPnVWK9vAYKtAcIzE4RmtVsaSB+hHGc6lOm09B5BbG3FgtFcxNrt7tV9dMZ6
M9XxNY+IKlNgzcNP4+al6/ccJuNmchmoam7rPf9q7tLNq13xX04osHTb+4wpNl/Y
gh80hufrFXGCoEJBch9Lvobw1Ps5QGxDLXP+R4yyFECNLHXDzChHKq2ZUHJhpssE
Qxet4icCdFZaH2RGW2m8CfWPaMLx3Bp3gmcp2ULWLG/yNQi+GR+Kf7wh+JSVFvT5
JxrSTvHqqT2HFYIa3GU2wKWQ1aCOVa5KfKdc4mpDlaFlKmp6LrIG4hrU1+JJ2t75
bhJSCAMMWdncYYtZm3HtmKXBEUzDdWmnArqcZQac2Ac7GzEeqKXTtTyAPKOFpVNK
Q7mnMbXhj73RfaEg5bqyc+i+DoH+P8uQLTdpSZGJfC4QzUY+AkDFYXPbHgVd5wit
M1aIDV5eRkcD1e5EZW7AxQNAPr8Lm63gxKWSYFEOs0FNodv6aYvwm/gBmgFWYSb9
ZqU2CEc9qFmSSWzjg86pzKKbsbVsxb1o3HoAQKjbT1at0A2gLeDktYoI4UVgsSRR
6s7nrBnqFcZy/gImAj6DWssbvv/ee3/2fiDm/uyYLnx06hfviUKFxFkLNW6l/CSA
Aoiab3C2xnhw86Db7pl6ikm4bTKzg2M7hcq9XsjF5fZ/LMy/hHVKNLGBstHg6iRP
VcM5cPCMi7rdjaEiD/jTOFDoPlVjsp6vqtNApRLFn1pY2MA61IiyflOlWNFzIxSq
rvZSpvpxIoAAb3Bld83tIgspNFkQf9LzhGnjrH2qNy8fYbcmJ2IbTdfsXbjMb/3r
ERtCEhqs7DbjMSPnLWL5GqiRBBvgDaN69PDhi1bJuPcI9ksZuQmKB48ht4MbR+Pn
wGIWx7XNDbAGLzbfMa8YSnlDFlhIt230W6h/edgaUemLuqCzsiDFhwbZeepftRA7
FOEXK1+Sentf0zSQglxWW2LuG/y+qgpDF2w0c14dUmUYR95AvvNr51aeeEkRwrYY
1xjqtInTMBFGwmMZuFiQ+pQMHChLr8t7200+jjIKgdvsS0/Ba1WOgKamHqvHaeED
HWWkVqKIYlYx2kpILuxd2fKh6d2pUhe26IoTRXrS65FJj/8oavPajMn+krXo+QZ0
pqMZ+9wWpeASI94kt7Bc8B2UHMQpL5kq/9umRJV90U9u3QsdqJ1va4qEJ0z/9o0Z
aLlP6ri7mNKQGbOO91VTc36xvi9hWpsZYcIkZSBOemvnZHcdS1hLY3umeT5Y/9hs
3woP0T/g8fDQkd7ufNYbxn8jd7m9vuMaxv/ZCoJvEj6verk5EjUcqZQ3M+GQ8GPS
t3V/Q8SxtkoYiNNrXwi60ali/9LJ9ONDKGkjQU+dMlVvLhX6O/sX3jWb2q6ZH7vc
+yr7hfKOr6KeZpW9OuKZ8PJriWsCEGIXb4kDmSaK66Eua0W3PmjIPk3yJK5htGM2
cArIhAfMYHBew0zq/1yQlG6bbY1v5PF2TTvdxeyk9zRZX4IJSJM6aLAtmduESKav
6LgyWqeAWs6pf2pxrAqzoQzv1VYfLw9QaOBACnSCPYyaMCBigEpY3567Et769xuq
yV/m3bTj/VVsnJZN0/93WlEBEE00fLop6l/k4oRy2oxOxfBwik+ayRPCDGRCtOf6
LxYZNTSfbWszDk359Q2RBvmMFTarPz6QVpR89PMXRUObUnKkfzo38JyF46Vodf4w
+zY9MQEaj2fj1Kd5DorPK3mdMl8UpQIjsFeUsuMkGmBPjKhcDAGKQhesznu6PSJH
esrCVsPrfKUxD/0x29o3aOMZtOYULpu1BOEBVhsqieGWnQn8TjZZVh+ucqCU9ot9
rF8ETT9PKZSj7fn7IyyVdXAMGkysi98g6Rbt6DHyvYO3ukJ1nyN/GHqzFkNQKqQn
/qorA0wfC1pgt9q62BHrvYEpY5bC7qriooYnLwynSexZbNoe02bmphUkBmCWhxDq
2PyaFZ/FDFPl7vCu81rYE2uwZ6iALzLxm1RyCAAd1v3MY5GFGShsWYuUUycvuIF8
EYQkmQsKkgivWbtcmLyawkhNTe1meoZJpitapvTN2wivh+3hapapYsB5xi2MSFwD
+SKuhhN5TEKF7C4gmWde85/oK9CPHlUnI5i7lNvKUTVeQz4MexLSXO4ok3FnM4Zp
hZD6jShiRwiH8UFmP3J0WNZdwG/yM+myPsTdX7ilSvAx1Kx4w78o3NyEYXt7ECXJ
MnSQ4M0AA5AE4D3C5x5iL4myVeAtqBiSVhAX4V0j60fIZERftY5yIeAzR5x7h0tc
9G+5aGJ04YNopWRZvA1tTUW7DbOevS8sa7S+cB1DwYj25nb9vhkKQDA5d29+n82e
g64V5NkOxxfo5zcUoKA3eDkRVHFah5ILHUZLvcPC15PtZsQL1AP582teOx9i8bhN
n3wM804i/ugTZFpZNExJLQjwNsPh46xmxvh3fF823Yvduf0NpI+p+XDFv4Y6KxQd
qnU8yYPP2iDh8W8RmpkOVAikulBA4tWre6teDzB8+6b3sCkVfcpcmPkWvKQ7VOJ7
jw/rT4LzHgu4LrYqscXTS22phJarRAC6Kv074xCmUXhPbqULQmdBhVLZaKnIpKR/
+wgAVmTBwbf8TAn8x8DiX6rLx8Js52nQ+zvcrvFmwMyHq1nlCPE2pSj+RleX2mmF
fEKlft3Jw4LxNMLWQJRNoa8tjyQR/DMV26D5R7/ZJHGnYFSKDcQEEG5g16h8YQs4
K1wdvwRfYr5zf4I338dWhf7/y/pKa6GpM1FLUwB9hIXZV5wKGi9fQoEaK5uhhUaq
ZCZrwngx1D5cy8W0oQ4RI826rHdnkIhzZi/Jf6TwykoI8uztsTeSheJFQ3MktiBA
HRUoqFvxtqXG6LxGat2AguUCxxphc1cRh20uOzJjSkcSscHLqjt0Yj2QHCQSLlNt
TW4EW/Oto37IexXs6uchz7aXD7Br/3JbJbw+pKo6uoJeHxql2Q1o+4CPQp4yic+L
HbTWCEEQjAVygEsnyolWQn7F7gmUuLh8FsNtEwG1XNc/hFj90NRyvUkEf5+t0wrR
vmb5JHfFUR3XX9fg7IN8A1QQbVlAi4I9mHSKkMY5/71uLksl3MzTwcVi5m6JbDwZ
EfpFr8en1aqNhl164h0h1Nc8nsckjKRM8AWbZemUEfV1rtr74gJXR26JatcKeaz3
MHtI3pZen53m2LVhaWWmu74mDuIajniFEK6T4Txg2Coq47JWNPyw6WeuyFaU7aMy
5TrE58J4PUpdCh/d4BsFaMdn3YxnHE/JbYMCRPYYe4DU+G3lvgGOlw+OLVUjfH4+
XzyozOCK4l74mgQ6srNiRHriuBkM6/iq7No8YCEV7pgYw4AjgfprPQFo8Z0XaXZt
DJ1J4rTWkGQbeKqdfNU7THlx+k8/+pbuiVOgauTCJFT7H1QGFIW1STTj3PbxDpSz
+B4xEgA2igpK5t4ShJAjsaZmAVSnHIX7hRe53Prju68HEc1MER9Asi6QWti1U0Sf
KvZ5PAoUugKyQwbyHQ5jU+y7Hiys99UAqxsyonSZn9kYqsFhTtXtkiK+HMg+NHkC
kD35OomLs7qHtBD6py7YYp0PiJHJ4i/TTedAquVhF22afefgAoBz79681p48TOuv
+CLBDXsg89JIqgReSfY3jHh8+O2wElN1RC9cXLxBHZoN1EukLE+CgLTMMDTvdC9n
fiWkBDX09Hsw38BWScxeXKZR8/1FtW0iUTwcscq1YeQFCWDHUQQcT3ooaf548lWI
Ur4qg+SpTG2ypSZ+8whx+uWr6IIT10UC+05ZAMZ2ImP9tmwTRMHjxdhcb4Ugi3na
GpyYI5LE4E3F+GY91yMQ3L29xu6n8aNwOhhg2bJZdsPD+V83rcZF7LW0Y77I+A7G
/Ywxl2ynQIG5+10zF+lxK/PT3R68pxFiXrLWKvP/r36pFDKuKvsO/YZTeSciyj8w
pe76cko1z+DlgKDtWuXQe5KJtDvBZLFg+Usk3Xlr50E7MKpLN5BIwW37VQXkOkdD
Cqn5siCKw9pujnTKN4QcfB6A5eo9q+D4Jfpxj7M19ghKaj/L4eF0atuzbrKYiT5u
dKBKSOHUfKLmEcvHScsPB9CW0v5JXNWfdaZLBPLLCMne2sAMGeyA0hGJsrifyCRr
Bk6UhrJwEo/fZqmY3pLgWpwSV7a1olvgSieWkDvRhvcNaLC+j5ogWn7C6aLmxUg7
StfZ55QmLCQorrukkazZJQh1kr1VVxLAixXAg77G9r7GXQaQucRvuhQCFlcHYJ4j
d5/4PooULrwb9mbn9WGOSaRTAERXAfMvw+uHQuLiZAmGoaUPIbdKQOkVSMw6CmL+
UFb/miYNswkNqvDzSZOf8vEcuyZNS7x3pxtd/eY6s/J+DvhLUrlk4tzAteEPcSn/
dzpbIJhKK3TyQ7uGl/UUdwQaFFebB5358ZDdfV7M+aovyugNb09VcL0Kg1vaoEdQ
xJ3nJmvSQgqu7GiOCUt76DgYTwLXXwOKE0yiczyTR4qaPWlHUN3g8KpY/c2bYtth
Qh2iGJS+Djo7MrL3MdcFClkKEELd09Uid0RAl9IXk4Da4WOqxBcMqtIgloITcoB1
ZakopNXirLNqLl5BsGMh4JLeWVyebF7zQzWO4TXSM7631AkPPMx/1GfWmUQcwLFl
DArf18Zc8yNhI4t3uGWHxAsY05QJRVefstQd4bG5x1VBow1T5D5xDPlVzHSkNq6X
subMVhQNPxOpq7itZGSLiJrqR8B9/1ehtdGbKx478VaVab3cgsOTfjzzwbVaPI8j
icpOPJ+Icd6JaVQFtmV1odLBpj0HG8Ji1jfb8zG7htNyXA2ql69vdHwvHYtzN7iN
L0DvCOocdMCoUG+o3cF7oKkDLmNv48J8ieLWfCwcIawjM6mUGwRTeWun+621CvHc
/MGKLrYp2jgBCHhtr7FI0MwITTbkcBic8s7grphH2eDhqvhyWioOf7EnlXlc4yja
XNcuMhqUMY0v/GfyJRpql/wi88anrVZ1IPpy+/Fl4tQq0O4lqVW7wDUhyGS+JIA3
0OI7EgsdB4DlcCXCWKpoiFPV8Pv0b1kOTkdm/EM57WaLUv1V5aKlLZDfCh5XsKKu
gh24wIV3+nPqhN26ucx/u9+FMRWv+4TtvlBeHevUDr4tABIfq6LOclEjZLbh8KvQ
jSr2VmtP/1nKMkd7dA0hbQBn72/cTi+kE8EgREPAnWP9Z45u3zocV7xD+ndMFGZ/
8bmtW4uj32TZ4eMW/1zs44lTne9THy/G+6/7jlMuXPj9I8VBBrCHSPq6GWl7QkjK
nN5IqnOQwl5NAwpsCa66EM5SO6Cdjq9sirOiExuNOJJXKFD7jJ9aXTnvFvl/Yxgv
gWU3R54gCdiHI+Bp6JEiz7Ft0GdOHQQ5lpMkp7yreVOBpWxHBpVGVtXiwDX10Cn0
u+zJ7wyWGusaKv/po/dtP/ZDgt9ZuZUyV1k1nrR1cz760PF6b4NWumvGOTBoCEzC
SGmieVw81ODJyUNB5yc1am74Xx7d/92zk/NT8HQAsqscvtTih4wJI27NwIh1l9RK
qxIuxQgIwT85sIykt5mcD2cR7okhK/j8nJx+kPCh4fM4ZUDOpry9G4hCgsDbBE4Z
/ckpshxBdtDqtk4C6W5xwxrEmcFkstoA6mEFXn+0gsxXxdpGB2bNANJCWVd1rCCp
vtO4RH18Ra0oM4QJxbOXcr0rBXeawLauemG4POpTLfMk6nTGZXg19XqQxY4h+y2z
4Ql5K/9JUEDAQ5Spodp+AbHeiQiUfAX0C+rFZqhaWX8h0pf5kiaHrQ2rZVGwjU0d
5y/hONh1zYM7kW0lVEE5AbQyndeFnnb8nhm/BlH3hf7IJik5/WaInbrYa+5q00r6
/Sn1CMqbWeaCKXavPYxQxyrxd/ZywIFtjXhtwyS0+DAkZgh+A54n6VHbw5gMF09i
OnNs0eexsbZbpqOLKT5jljWjWDYEUQqrjAFsqFjW2gSEb60l+m++H4Mkpw33YXzC
kAuTpfpYkNi1aVygF77jXnmt3lHKdfhqjRr5VNzjQcqDiDPcWjdkE0PeIiWnbFKs
JoG0gcU8u6nM2X5RsKGZdhklGkTRK0hkHR5gxVflOXL0r0bZ/ly79EG6L0nAod+l
ceEtaQN9GgAKzw+/tPVkdfeiGvddja9zBUZst/7J6DAnuyNbzg7hlsSH1sPDaelk
N8YVQvvADos8Wnr7NWfsYQvkJ1uQri5awi5X9gP0oB1YXwEkjBHtiSOPbp1e0GK4
6yhvUngaoWYACGih/1Jq4i8lVLzB9vXaWyubwoHvLWxVEHvCHCYiCX3bffjoa9U8
i73H6Fzeyp1XYvU7FnXrIhBoD1VCRt6CJn+2wgCpBTxwYvpj/UobqQiuWydBjo2l
qdNNpH04iBeLmI0jg/tAqUAINlvf6eeVQLMJkPmvQrtXfwWRuPnl3McxuEFAe/Io
0BgrEt48H5QXECYymvrk52jpqh+HsuoPiOvlxuzLDdKqWSca63MsQxn4KApHcfHn
ws47UN/5wyYddP/TlZywAK/fNrFERXZcouyxbyJJsOD+wxlIUsqTb7Pez1DnO0dW
RZ1M6Ks6VjA7XL+C99zxTJntsJwH9/fAM34f7zr8lrYqr3mwSR5F0vQSsF73Y+Pj
n+ZHuagEb09+g7364FwOMMUBByJoHTiYPQUkvWBz9+NUwcYtHtGHE/TSlhOIp9fx
E9zXKyKBWjhlKX868ktWvG1TpXFV5P/IY122xoJuIW85PjxLUJ6imMcy5rZ/e5qu
ssu5lqxJnGvomABP72dKHjpP6/8geLXV0B5WRiwFG3ztSGntA3FXZDxZFstRyq90
MTZCa+GFU4X8K4if9hBIxEwIPfwLFRJshvK+n/IsItw8d5mTQw/aJxcPLME9i27/
BBanDnuyrxrSpAJoHhUqfcaul6OW/3EekB9n4fNnxSr1kL8Rw1SZkc4n76o4/Oz7
uwt/o3K05mUH8+kmHs1gV0Ql99FCGtGXG61sDmXxFV1dWpxXR4Qe/W1GcaX+AhRX
51eSGWEK5B3EJ/APBHF0NgdasJcv2mipFpJ08/fdXmcFd1xoD5yX5WcaRkuVIhrd
fLim3MhMQbKlLlbKX6llsS9llk0+BDS1J+usOzUilJBCaDl9jwz6ur/bfFaHMG8K
Cxg99byctjQ0xdCYcTuU8PKnMCuuHYpcyfdTbG+JjQpnXL40cyjEpwa1pDQKSpBF
M6fwUcL5AQNBNnwn7xQU2wtDFkfwoJ3cgr2iqOFv7vvBq6W1zVx6BwwzM4U3H8ln
XDgn5aob5AAYNKKf1smaKRhMlw2OIhNUJ0zh4cghJKq6L+QNvA7gSwWPZEqqFnDc
+dBWvUK6u5Zt2dKBEowdrspG0gNkfrWfFipAJCu8Ao/xD4KM5unjKutSi3gqVSZ/
xQFXtiu47Nk6eFynhYf/9xnz/CF0p/ar7iCHyyT6u+k9yCgXRZAy0T8otictK7V1
hdQ9sYoBJRkUTdqUJfl2Aa+L32cXmXkv8Y47muZ9XVGK0O/Pu9Ga+QHqNQXI1LtW
gon3Jm4cFCjDVpoSumLD9YkPCiaPZH7eQA+LcNegtPxTwrDesdbIce/XOBZznbP3
AjB0D9OGNEZzp+l8Rkike/FQ5L/lFbEqdppoW7n50Q3/d6ahG9hW4NFsJjKTQjn3
aRDzKtCtVQ3OoFiAMLMS6hD03TctqfkW7lKLQIAb8B9LCY5K8zKxDJTmNGPiYch+
OH39qC7Hefr9raZNXh1O9iuaOQO3UHtfwRVgGIaqIiSipGpuCqbsTR77Q83daQbg
3NOZtR5p9zgJ92LxZX11uGs/mQ6/nDnY135EBQfvdr/2tETiv+1kxn2VVwcCricQ
9VoAeJHSUSs4vWhIW3lA58JA+rCsNQ+xQ2rX7qC5bGW8S+hJulp96N7uB6HMSi3d
QuR4mjikkwqctLNSPLee3h8qsdsG51GgOxGrLUH6cf7VXBERZSO0nx3TKRDffCRz
ZKNLVPtkPMRk8rUXa5l9aDgMLd9yVYJkAS4e7Y+FrSr+9uCoj1fu8hrlQqOYFDkb
ofZWto4CZr1uUCUZEhjT6XpjOCXSsWz+F7Xn/AL2lxTb/xcv0Q6teOeN11e61Y0L
4P1c0yEfaXbD7qCnqPqol42Gi2WyDsBn7+PJuThtmog+4IUu5lsYApf2esAW4QYG
lvmzeCRh7ZD/0SvTILk5Hnz0FX7CxLE59SXlQfEK9MI30EA1Zas4XpNLQKmA3ptD
RJVXeb2SVblPR5TpAhETrqLXpeBMJwgOXd8tvMS/qcREZVD736b5TYyOjbKyo18i
686xvcTS/zWKYqvJqtD8gNRsLiXjGcvsafAtJQVJwKfD3BUIDIT37wZXD8DG3HPV
Ew1t9ITJSQl53JSB5UGRemLOye7xdax8/rs3YjCUSiMz5wb9UBsJBaVWnkuH4f6W
Yfj6y2eX4R487Y4tvQkkJ/BvjFfkTL3jnhnC5C7HpeaaTHl9wIrCIexZ5iG5yAyH
ZoA5vFO9ONMrxzPn6pj7ousKcqvKYCgwyKBXN0/PnkV9sV1ROE1upp9CC0LsHmbL
X6fI0+uag5pvI4H2U9cHdnoeyz1fmOerME07rmFwcemovCC9iU5ojtfR/CcH4kbZ
tdOoqW+A6Z6A8r9+rLe1QLKkwZcy470DrkBhX95xdR1aa0z/rCG0yBSp+zbIecpz
sdz/0Sod3N5Wj/bBIpKpuJmrcgItXhVpJfJeVS5Kdcwnot/3fxBKdt2aUL0k02lg
W+DGyO85BAyqaCS9BKcP+FulDmMTQqpmRkbsMipwy536of09tWP2bWwjJC4+kF8M
hCp8eFt9SZDyRaU5sO9jduJIWyi9zBqULZ161qa+ekm0R7I8oVlugK3U8pfBZfMK
vH6bSQVT0UQquJWNWqa6vkePsY/ssC+WvV8cscZmWCNy1rOqNHBGb2UkFflrWpaH
UZLIA4FwGoMlnhwhYKpJal+eKHtXYndXqva6U4bxLcfU9DXP7WPTHyCVH/ZceIQa
6iaEmPuG5A/9BWycdobOvttd/JSr7viJg6H6h8QNkK3xo3UZ5I7MYs4h4C7HuuYu
pH9uiHMq/OieWLhaapnJU9E/JOgFeFPbRIJ5AmFakoHB7qJJTb5cQAedoW6OwsQo
oI5QxhtpSR75k9cunAuPy9heju3ofPLBI0aRcvdE04C81c80BkEBkXSTqEArtkxm
heexxlGHV6CDzGNvIJiairal5QGVOzFInxuTt150kgSTNeoNgZhtR7LOrc4dR/q9
7ogyLvXORErJkUbqGemlebX/LlDTG/HrMX+k/17A9pk4XoJGID7jP6xrXJwSkRTf
yhYLJywjR5ANr5+5xMcZf6AHCYdXToL2XOlkjkIz5gzh4skseYu7DgNKiaLU6aHu
rFH5NzRokwZ7MEqx42jFHmPip46GQdRE7VL4O4z0wlc9nvbSyY16GU08mzUNzTix
diRcuhazTEPvQ2q4KQ3LKQRotEhgzDyWHSbyKRpHvTqadFKlWJ0JalmpkG4eaFOL
uyqIVnAEMWNYeiWc/ZJb4pdaa8Q8OOvf+wH+Jvb9tqI7Z5m1XDKxpUVFUapIYBS4
/3gsgaA8X4Ko6ZVdoa/8AjuVfPgACK1tmkJVr9WvSvUFmYEIbGqIiv5yKTyP4gyS
QIT5ZciudRxDZtHnBizYA6XTMVu2dEOB92zeuyanyuCiMIGWSOE7qcvB2WZOevF+
7COBe4eKLaUj94CJAWEj8s6ih3T8kUZ9ap4byFKrs6ncaeyS2RirgPD27h7wlQ8k
jZeIBV0DBDyuIjw4ovQXkkW6I+39xNz2AY1aXfv6XjcXgzb94lx9oLSvs55BJ2m8
7KK1sa2qGyyIoHhNoWFc3K/nOOaegpZuPa/YbsahboYfMFhyZ1hqy1XXmOW3SMud
JaKFXxw0xh+YK6HBrgGOtT0sw4oBQe3OQnbyv131tKZIMVWRYhfUmXUp7AgIJJ1h
Gj2aw4haKcjX3xvN5uZN57zpULEzUUKBe0cokaReSYUj4K6xYPIrOHKcklf0VB7E
ki5Qza+/eS5HBrCSL1h0vfgBMRNCMRyj6A59s46lMHBNXw2NXTbANQTD0FI57H8r
0UReVzHNS2Uhwukc2CorJD5tt/snf3fLr6uLVGBGVQAuYdPbvaZPcoe/5mlQHTnR
v74yl3aAWFHL4HW8Dk+HI55o9/h9O5V53VsyNP8dCeDKSfkqVRPWsjALapuGw3Xh
seLo4pmUAkc1bctxry0TFcZZcBKK8MFNcwRGH5r+UoQoj2/JA+sen3POaJDkK+aj
u7adQteCTqWG3mx96n1Yb9cxfB/o5S55fyTVS1NN7vrMahp6nXEDzUi1HWoAg8Yj
jU9nJoopN7E3NasnrU/z2ZvQkoegRTM8xrFEmFhSM92u4fhu4TCvi90RMk2e3Lrz
UPAPk5KoRRPguglss94NpkMuqi/N7S2xbTsScte+68MTzuq0ZFRssftvMGAWtD7l
pVj+kSid1ST0417Z79rYNkn7qHiv2gMNRaqEQ2yim1iPWa9gLnqvbZtJtXD/qlyH
xzbb/I+W2QTX1BBFated+r4MnlQTb0xp5rfaAvO9Rrh/4KjZmEi6qSDI5WEbElbl
R+YfI9O/jXJUq+yV3Tp3RSrmEOLE+99YDZNFHfEP7dm0gr1ojOcYfScmxu7+xJD0
8uif5vzwlvcXwAKuPf8RnCiPtIYbVQDrt0E2pIbzDmm9IyJ3EctM1Ed6CPdieTfV
8Bo1lxnFCU6V/X+MTj6pPKgDh2ElGImXshbf4fGcA1PoJ6LaLWAbY6CAgDrlmfXc
wkkkuwTgTwW+733WCtODVcm6OqJE/kdW+prQ8lyTpiZUlyCmLAk6zL3q8evmNS/f
rkInzNevX+g0G9/syHl/+wgxU6+Y/r891Olq7Ebou/bP9JjU2lzia+neiPg4WrUX
tjxbNmzKbe0SH9J6wpF3YWGuSYaa24OpuxIoTJTAiF/DXAEwxO7QKkyagyB0Img3
yIs6a4TVPopxH1wLlll2D7NpNQLB2xIwTGb2A4eaZbnnbNh2G3rDrIQfDac+IMuU
YTHuydtwpc0INYG3kfOyXzk/39hUCQvapfXWg6mbJYRYbceIS9HGmoxn9vNYa2/R
MBKM7MQGJfLsBOECxsM4HsV86NHeTut/mvPDRcdFkhZlVUECtNGoLFVJ4h5kwdhC
/hqfOqFH8UDE60yaFF5RWmo2e2G0PumEfvidRB5E8LpSMNrjeeWHOgyzBLUzMvFF
g8hZkQCoT0xOrsBI5xC7gT57gvsLEtuYF/VdOaZYmPGGsvI7DLkLzq9ama02Tz/h
2RsN/ykZy+Uub+igYkViNUptvdPY/jsjupyCah75mKg1Mo5A4ab5jjlnAR+fZ1aB
x/P+1sJMon/YElBWUCVLjOhmcK74JT/3WM6Mu6FvKpFn4BEyLVbDPJHdE4ibG2KK
5tWGWbxtFfRCb264CQIo4XFaa1NumH2w0md6IKtCH7ROfLHqPoEIt95RSbhkzuWy
xWmlDevhDy5f13uPW9uUGNpeuNAO8XURHAOOJsTgwMxGrekfPwzFAiVDtkklaCvA
NXQ8Le3+APnA6BSPRS729JQnuell8vle+z9qgQdvbbrFWX2fI/1olkDsubUDVE2/
mtVQW9H5YluOONK5r5IHew5CpnMrjiDjWNQJIAmHEieppWvOgEOh8D3O/Uwa720k
ZcfcOA8jcoi7HYyvZT9WCBhfnyVxlpF14ftcn6DfG3GdKYgEV8txNdyhiGOuQcMr
pOOzRUEkcKxEiQdFrZx6TBSx9rbsqAJhrUbJ+u2c+jI5PPGNEd+6OjvU+tE9hEwJ
AGRIIfIlR/tTDFBLmuXCjHxvstCeUScNMtq/44LyEwSF/WSkG9DWmwrsKIWBOSRv
PaybldNdu1mHWGqD7LNI3R66AP4eBMhDtI1UzYVrbxRAyu33inAwXu4TwDj4zuIq
nfsxXcpVY6iGvTC8y0BViAd30w4e58V6ECUByZCF2/vyCf7KN5YKxiYF4HSbjMEb
j7kXocNf4pJl93SWzHdVoAwxUzP/YeYI2jj7etB2/34yWMlE9LWJTLKaEUChXCCM
0ofGI+82GxtV608DqLyisjo+L3fln3cd1MPWsSCysYtMELL/CCL9hM8om38smvNQ
c9qh3/TG5vyRns2GBZlUAOqtVg/I0jBlAehHGRnMpz8mI8/e8vG9iuL7Gonljo5G
n7s8NreVA6cFxtqQ38LKJAwHWCt/SIAPh7whwreFkhuCEFPz8nvB4XfdttMo1jTo
7JLtoCA3T+VcHMxE00KDVsgJDCEdhq8eu0ZhNeV6PBAOeKusp3RQjSZG9VAdq00L
HioajRVrSXeqkEf2f5jtYoBkVPAYfWjfV0TH6EfubjicrqJSjVfLkapyLPRpzjCa
B8HfDMDDdDmlSPSF+FDlHM7QMnePtQOl26cu+o5ZtO1++eVRiGlBshOQBI1inKJE
yxRuFaMGvXpaHc2UB1IK3ohrxjDjsnB/M5hugk6nYZFgRI9NidHWeofTAKOTVSro
SI7qtacoMESwsN7K9fN4PtRJIoWokjXOQbHv7+Agm5DeZDElkDQyzi68zyf8hDgp
fvRJGxAAR8domvsVIa8NXeUtSo4pBBYguwrk3QSRBgIemASmEdjhg7gXkqkCFt90
4ZtCNsya1OsGbX8Y2TEXG1gZbcrc81Tz4i0a4PUAO5v5aeLTj/tcJ2ffez5tGLv6
vl0rtTw5EhRcnW+ZyQXXxFqxmH760wlnP1NWVvlr5lpYC2aq8uhQ4VYGy8S43/yc
nW8zU0HAB/kmCrGRri1jrUj8FblHn/dfVoZDsu83pmXcOQ8SzEDgOrxLX3BXAUxa
4adtRE2vhEOd35Ua+O2u7uNikngRX04VKHblunmTW2A2n7qgHO/4Xw5ci0SHcBNT
ydMB72oMD0M63lsBriitREFj18pBjEaIWL2UMFsAqgOkDA4uGiM/5ftsiS2fDVG7
Tv/GsyI7XLaIU8wSc/Scma95uMGFe8MC+dZT8pj52YrwhrJLxOspQ9qnOVHqcQsi
ipD9CL9QC+gk1Ii8semh4dTdQ6ses2DZfHNH7N7OdW1JVfzBg4fddaizkGBvGKVP
YXj4SgVy/fNDhvVhjB4JkjG+RDE/hXPddSiIsSmQH/IHw6dLwGKhEc72cGK2LNEG
VIREChvyhMEbK8gRBuimKkr/SD2aR/1oOMzNZ2VroWYP1winwo57gYPSSl4Nfo5X
/kMmKzN+6wFeF1dbs0rHyqwiCMOD5/SLnTsyH/nfLlfeN6eAtpzUtGCOxdzn5DVA
v8jMbjRzYvPWYB7+AdMR6ZhOps+ZlHW2SvlOdfFY2kFD2904J/Tu5HtbENhQa3t9
psqpAN1+lfofvajwCzvxAsn3kSa+hJyKFHarL5JQ3NYb0DfkEVsXNeUnt8aHtNrf
FrmtpqOdc+07//GAITlj7oCFj0UkqYo3TNgXHvfT+kegjNnTbcQj/qjMqu1hKhs3
W2xdCsVuzDXRzDKF+toE4zQA6b4w7OmS4WWHKEvBqs7l3R/I3R9tLuTIMFLtE4Jx
ac7WC554fc2FEjFYq08ar3ZStvtzFaeae8Cx8Df619cs+GCEmG59MjxRh0hylry+
E+VjBIh37OHiS6zhs8KioTQsKLc0exLS9tYmQIot0OgKPk7SVCzXz2z7+v4xbTkx
itk1Mhrh+u3BVmPm3OD0m42SHXwSkDNF3xymUYOvkETJmYF05PanyllWEiVAtNxV
KBhZEWpTDDhakAjynYfqUnQNCQ3S+Fu/ChUMFCAsEi6hMShANuhuxXS3tUj+2iHW
jnP/CPcXeS38yX4+PTvoK6iECC7zAeZxQ8Be56wFnDCstx/sHB/GiSGyYm1T0uSK
uRHY9EL1NAkPWtIr+JEzUbQ7oQwR4S/wvrPsJZRpUtWpwDIfE/hCUeXMX69wgaPU
DokfvUfyQJ19LGvKVSqve+C7wO20tHlvKMNquzJz0eteZeu+zMp9ziXTsAnxXdWK
k8yusN8yhlBc8mUllmVu7gEdLrdzB0jS7a9o0AHqKWgn8BRcGsxOJhFbkpJi/9DL
9QmUx0NbhXWIPF529J13izEhBNDhe1BQoj/16WJA1aLaFjmn37sL2O+pGJp4MIMP
xRKUdVDv2N4NPViSK+WlSdRDF1GoGW4vghwAU94xwO1roUNpxCtizyEtB3oFo/It
eZvA6n3fj9Nlxd5xEuSpRfu/yadNUsTLVOBgjUurbnmDDY6pteR6bfnuJO4IdKx1
aCzGNCBzpYgKKzgVCnsgvA5iI1k3jf8W5bxJSv1r62NPJrcQjmTofiNNFhlOyGHx
55EG3k93kZHjbgZhttzZme5l35oFlIOsm+yWkMFcUGQ3PC57pGBgLgX/cJsJ72+q
/Pgwg0xXuWamW6+/YtVVGkhpgl05Tu/IwYQKFh9ceEhcrb/yBFvNDFVXmGg8ZvXa
RDqobGS3MmLqDaJO4jBQUfEBo8TrIeugHLiTaK4uJrAS2YTAWOe3CHllACVZL0a+
Z430AT3Y0ywWhB151jcNPShpjIOfoHxXeX6Zsi6yTua59Jo2n6GUZOOYKFG4bgGS
wWYTIovBldBichJuAUqVyYcUjf/RtQ9nW/PM+y22SPElxPc9FhTMHnz9Wb4YJ2GH
fMFHYwMQryPyCMwwjl9Gh9gBnQvB59wj3xK5g/POn22lmHBSmsNqtwF/drthAD5s
tXl1Uo1kl80jzJvgsF9+Iy2tn4UZ2zI3C94uSg1vdZCxDlKH/beEPaEF0sxb+l+D
esnlYGnjOBtXiHgm3cMB29aimfJzY+XoAZZiO47E6+CGesd5UPY99hLDPqieIEvg
KK1DjHYOQC+2vME/YcbtNMF1GvYK6bgD0w9uy5aOYC+mxzcdzBQohJCzo3ITsROb
IgHskWHlLWYVzYTUsy69xqPEGJa3vc3U8KmEH0pn7HKCqET9OIq3haMMpsiCNTuX
iVby7r6F+fsboQyqOfQ3a8Lyn30zTsQpmT6vQ/6O7QVgxUotFpm8pTyVanUiccg+
FwNArtP4dsqJsndEY+kNd1br6urzjllx3XlYJFjlxgifT/kNUp4Uy1G4xQuiLmH7
c98/n150iZC4j3aRa1rjUXqhF4loxyZQgwk3ICVOINnNAdcxndTOeUYAV/SytIlr
jskfy7MvLmj0vlIfj8o00R0iR7buF5l5t1RAishFODPwTZvxbYq3LCUa3IJqwnSE
/i2NPFfxDYZK/uqN4ZYqIiaBs+Ejz+qKfawqI3D4fqAM8jjucaLayFhYFb6fLZ/O
B6FsI6WW4UnRDhXgoW3Kuf6uU0+kUYdhqRvEQ25FTTrxrxOR+d/4NtWkIBpUt+Vv
8DLorv/C9sFPqYw8ICTPmVbsfkhpN3dN6FgJ62K+abODw5kYD5w+n9diGtdWEPyr
re4uX9H6Bn4ZfYxkk1BfUd3KIZT83grCoFC/WLs3AQ3Jk9udxbkLHrenMiExI3yu
MLdpwfhC/aWtrZLm+n21LxBXKEPSw3qDJNhU5cijAzStH1kujl8oE7AHmEj6O3sL
bSVK+UuKHk9sS7sQMZfB7aC2kgCyl/Ee6Flv/ndFF6wqzt3fozR0aSd1zWSVSvp6
ExwlfF2XfY4T2URYMOOSDEwHc+j90YEwQ2hA9yHzfkuckF8aLQOmc/qrXpF0PWGx
XDZdHeIT1qUiL3VYqGCICAztw5uNeaMnJND5TRs8RqVLRLgq/XQT4oNF4agiQcPU
GJ3UcmbDhaILW86YjKu9+BNMpYyppPCujtJOcRVQUbq3gD19g92SzWAxvh9oUghP
2xV1V6QqdktafPPbHeLJd30j3O+OTVBcYyDhPil8ZjIzATPAiwdT0aLGYlgh5lzJ
XTFi3/i+1MjlkvHlFAx+s1rd0A81FMlfmeZzl54pUBL4sQaB6szorC6NvjdDMt1E
fbTJXqWixeyIHniJM6yfOUrsdfB6YBG/tvto8sz5VRyeIo7MD67sfl6Fgx4MffQo
HEC4nMIe/yfxdcGD4nK8l+XdRwn0yGbFGv/olbN9L1YAoYvB4JdPrwHrkhu7Z9gW
qaLteOlG8l0OJV64PQv+eo+DT2WDwHuYaUImzoBk7KMCTZy3ie2zn3Df24sdMXXY
0TUUKxg1OT3ziuDYKJIswNyvKAJ9NpL+wMpY5p3u2IaWrrKcYDr22aEKi05Q4tDu
//a34Kswd+n6dxG+bwpIZI8cblaZvpdxKDZ14mMAddhqibRKgtT/Yk43z/PxjHO7
5Sx17ZsrzDKSdKeW8+8Lb8wleTJQ9yrNM96EV8ekMua8vSEo2X4p9Y67Ps+NnDNr
yndHKL+zp7IN7HL7dLpUNT5eUJ0o6QjRXzXotBFzX0/583MzMnPf/kOQKbYeG2VK
Idi5ScErwP9dItx9Xke8PEcLjSLJNyP4Zun10bEiQ0Br2liAMIro1ZrLrJp3VVvU
p5jMXmNUNrfuUXd2FiM4SdJuWuRQ/jbRWqdt/ItG2iBHaVdA6w7GrNzwx+X/pFYY
shCt+/s60d9uxYlREhew3pyW5GFysvhEHyMxrR+T6+Pg8tw1A5H4xmvSWYgQyk3S
kb+CnJhxDrrVm+HMSLlKc0dBFVCiZpWnnEh7nCc1YxUW8tcRCDHTrGhXnDJlzIGU
+TDZisA4rxrZTx1sxZJE2QHYYlA0QvEAtRU+e1EQ20OYsWRQi3L5y3cBv9UHmfIa
1Ziqoiwqb/inUtyTuiYQiEER6+l5jJXBMr5VT7h4UKfEpHWk6LMnlh8TRG3XniXQ
4JoLJ4VVl0Nny8iJkG+vF4j8LPgHrdnGArf+gIN3QuJ1V2v/LVpozaJKSFkipGbm
jwN6O/qwU+1Pt+ZE3liOVufvt0KOAe32w7eQe6WlzmQlML/q8F5OYGAvZDBcYr+d
0M4VneCz6niBF95gVabV6K2/KHGg/yFYzpr8984GdWfOXVUAFS6Ehk84wRLZCX0p
uK7/Esqn127/tdt18+bKsbIuwKFLugHwlgNmYueO/gUmr6YCPyJIHbaTzfUdOuRP
CGzDmQeoJAbuXob5hujBvl9TnLxxfIZ9zu852kuAjK4KtHQ+jutxNeML8pgry4cJ
e1gGESbGKJgcOQ76XmCfEJRTLwMhcYTEyO3w5u/POAj97SAKDn1bUxHG7FqMQuBC
OdqKiiMpOHoZRS/YZZFN8SOa482d8pOiaNFC5EWoeIykevsjFXhai972WJ4pJKir
W2EzKs4Z4lZUarvHv+Gq/heAeifFxL5gKRjGaX0nIW1pOK3l/3bEDX2P547JEgMD
aK3VpHPpUMZix8n5fy0buoIY9QkpASJr9oJ7A4js+Xmk+sEwHAf7dDuQ88UNRTAR
DJpvoaRXFS7cQHgwLsJFvRuaEQxWsiJJzAg6sfvRiy/IwceJjKXOZfIyP8nCfPN1
Rrb2k4I3WJKuZhUZXL0oKX2Fsu7zbaSlVTCCdvQENH+VbUiQwRbfz81nhu151nYn
YxiskQHQxrsspOLM+z15uvZFlpG4wrZu6bmREAuDgITiwp8nfzgUusT41wFA6weK
F827dg1sPWCpN6uRcQsKjD5b7ByQMmN+MfvatpLiMleiMsnPk4md1SfDTjfW1vGh
SDsBgAETqNxMzQNn71RrrFj5GdAeppVdF3iE7C0n9vKLju4T1bqN2sveVHuyQLWS
kZeV5hF3HHguRMpSRa58WAfHmbAgJ+RDCZARQb49E7xDFfcTe6sBtk2jiB2NreAr
6U3m8aWYVX+vWkh2DTIIOzpDNG833j3FhlGtx/YmjfsO8HvZnNhu6C7HhOI2PJ+g
0BaLSSTnw3o+XNky8Pih5IYt6xMa/VGq0X25emsqhXWKsNNX7xNCKjnhwuefc6E8
eL3dtoWo/NHlaGTZchkCzQR4FULSyF8STvvU6A35ce4loiQSthoZl2iWuD/mMu9A
aZyF4Kz06VGhL/jsqFtprLXxkgDYL8ySsxT1rtslLWAYJM45xVuFliBVyZkOo6/v
e2ICvNdNsm3OeiKVE0b3Tv9RqixXJtmtJJHvIvBEaj0nxEtDooMT6bVwcV0K4V0u
5/tZvZo3GmKXjBUcCs0dWFHMnaYrJKoPSPOSEKbQ02Ehh/PkGRRqONSgbmZwBvCl
dGsVYzKP3OE+1/TiLGoTWUzSVkjt1+6u1Kmay5zaEXKxyaw3wU/gLuF3c/Fb4TGH
kFO/+XSSB3V4ZbOpmUyK0EtaeUUyzw6KM6P7OFq3v/c9nHqqfvX4LxJHE2m/x2Wr
0xGhQ/1aUHpXYV1ZEklEGd3KnaGyVh1A28Cm1RPuvwSTUEUxXzF7EIMuKqoCTjBr
/HD8dh5SQ417/oGwjqqhjKAEPJ/dCAm5+MjCOnvWFxmECC9fGkGgl/jT66mO3ilR
Ci3aj+NBMvjUi2y23OX1AnkLOVluV+g8GDE3MVGLVyu34RUI/h/DvRe9rDXN34y5
rpZQDlRqUWKByIyQPmiJS4Fptks1gQt5IntWkCRL+PUybk3daLM91fEptEMEb/mJ
vQaqrxPMlsfw37CTDBdNHIgNIz8HJLPC+JLmv5wev9t3e8b8W1LnTKfKSRHV7FmL
Az8fm7j4wmLOLv5Elawm0FdQgxi3cyxSy3Jt3Uj+WzC244JkWNmjw9csU3bqoaRj
++A1Nr+MvMv6Gv13pHFDx/hKKBfp9yCwxv8iIN9rbIDIDZryLsVl1IKyTBIBZgvI
0EAlhX47hhoIonm3kTjLi+CJPJN1srmEKO8bMA2mzWQYQFpTYUAZlqoySClnSclU
Pi6QDCPxP/O4aXRAHX8Tdg3+MdWyNtqA7oEzU7v8o+4+Yg2z5oQ5k7aTe8xRAM1J
rzmGA9I0YaGN5S36VUzmZkPXzL8RwgOcFvXyjog8atNJrsFCZPIfwpaJY1cAj8HX
CeIfPoFrBVVHyolAclCdh1ixFjnNiu3BaB2HDRnAYGAOuU96xYWEKHdCjvHH2QlK
YRd6srqqUk55Dax9DqXcQxsg3z+3ljyK3DrW4FuGrW/ZnOFkJaozcAEPDR+t4JrI
oNmmgOYe5dO/TFxvpGyDEOKztciJDA6SNffn4ZRm6kHmLLduQIQLGRN2AVfHqQuX
fDsbyCx2KHQa1wI1M07yFl7MrGkvgVCU/SV0LdwTCk7gdS1vGVo4jqyqLcN2S4TN
THvfFpvPivKSrutMZGnT7NuVanfdYZBQRkqQcwFHFx/j6b1SoUg9X4DOAI2Mz84C
x2OTHiziHWz+b4a4YHXq9W2qZ7roTEhbb80eGTFTlxc4yAlKGdpZWjPbntzlvvo5
vNb7Ylxbk0Rshq4n8oAf5uggynRbIw/3fTVXB017t4izGn07J5OtSZj0u9WZ7Zbc
0mvF/hrNs8D98SHw8HvF9MXlAyh6rxcs6eP4ScQnln17KkJkMq7B2O3qI0o9aLeC
JrYjskIk8O7v1M3AwjIIpC+ln1jxyQ87+Bv5Q2NChOK3mvUvVwdBLaFpHvYhF1bU
l9yG9jAAL0JyfuXpCbc0CM7KUIgcMpNdJiui2OXyHE7HMFm4QLGQu6i47dc7D+y0
raMxqTo7IMyQwY0g9dv5Jcg8rRs80tSJw4GeJcafW3/5UlYZiAHkWbOE9roQc79S
V3azdaeVeabekIC9uO4uGbkmmwSGeUoq1SPaVqlzpHF9f9Fa6cYjcksmP8vbAtpG
FVrBOv+f+gjxME2x46rTmGIW9imHyeE67TwjemtV/Qo/NoPNBYmFId7F+0ET2LcP
XAdd91UUaJc1+rI9S8bKQ4/1ledpFVlCAfANSVxOGMCKGBUNQBZRdqMiRWPXPffd
PLmtyY53RdRiiOUTIZUiOD/kPZFUwYBfyFUG3vcxEYQMaZL9DseQe138Wdw2SIbx
qHA/FDKHI7QUgAocLVSIvECEV/qJsdADuo3Tsw0PNwN35/EWXP55+cqAuYzS6g6R
WqDuYBjVjyphoDJDSa0nQie/SIChn455DXC/9X+A0z9AuYzCGVfZJODzvxknq9uW
fo3nO2E9397Nnmye3i4c2pNOSqzgf8/bJb5FidGmYHquZ269yBM5ZbuVlYry8E26
uztQ5vCRcK510uDpuAwY6YNHeEROv08RAGe6HqVnVMr46Vxy3ZfpE0dtm8puxjUV
BeTnn307ZHn8Uux2ET2Kp0elB32O3EgZtLqmO9G/HmoKoQIodrYTvG9jUkk9jTLl
9CgV88waKWHCPISnBaQrAacg1ii/upPBafUZ2RGeco53VOTP4EssdglvV2yEWwFK
9aRrmZ8uXOlPnxz2KarKynICbkxHFEIjx3bXNTeUajhOfAIhEyZKiSTclDnDWWmA
RQTu0V9SpiVXi5Qtly/kQqSF/R0jbCpQ1u8NNfWOw/4Rd8PmBnXtyOXBZ4zUUcQ5
BtTHqvLUlfiFUdEVhl6G/boiVBZmY24uzh2WXNBNWZN5gCNY4J4/r9a122P+ECAA
Kp4GCHoUc3LJMQBYqFq2sJI25mF3f92sI1/PkBSWDNUpdYfXiHcNCcLNw1rAmNik
XwCKBICLoVWGoL2b0gcgbNnriQX5lWwaiERSmG/9T2zr/Cp474sHXcTlKhEb7GbS
7+tlHwblg1X00zvhpDZrgS4c1fhm+UahgPohBosoaOa+haE+A64FdKKePVoD4qx6
wYeA1qYZNn77H1JuAGI62zDhpfNsyEyQgAn2s7Ii/NQewrhfZD8X28YPyzSN3sIo
ulaFSFVHH6FpDsynLjPiw7i0quLw0OH5NSvjGmdQF3RINlTBDE+Yvy9nN484txEn
n7TPT207312Cm6bVXYW6DGhXivAwtaxl5DegrXvGc86rOE0rVC1km5Pj07LjsAhm
VGjPcD1kp9jkZmvTVFROYpCbhbzpE2lY3KN9VV8gFavpmsSX46FKAgFy14MOljoU
lpu2bOhfq+DfiI84RDMs2bfwchBVOAsfa3HBfAC1BlKkUfDHDVKWZnDgwRT9Fcr6
qoWMaApZSacA9fh18Oxy80A/5CQn38xqePxO7P1NPup+Pj6fFY6gM1frVjWALWdv
7hhjQH7bSMH8RMglHS4j/6Uq4l5qopWg95EF6c2v9IKoZ227fQQoMRZpSGgDbJUF
jnDTS8fi7uMaBLWRxY8g9UA2AynLkyyRWjCzdOgoVM6b3Gnjn7NNiMn4jjstmf1P
hIgBniiTE3M7V95eR91g0fKYtnFxFvgIrWNNEbs8tSbEy2VHaCak8hxXwbA9UyB/
jBQY65PVoVEIzLfdd1JQ09rb6XAI47KKXKdHqcmmzGJDciB+RVzguzCxGphaCGUw
wKu0fLXuSvpYduGZUgPclHhBep0ThnSsRr0s/HQ4aq9wzmyJossa4jYiZUjHPZ3a
WDYNDM9WvkLD5YIUTimSrpcES4SFcNPuYFwjDqqGZvpcAh+AYpZkad2M9y1Ogs0F
3NhY7iyCGoLESy9i0KXGgYwzvlMBWuEpTp2la6ui1TRvyoSz/W561BxQCRMm+39I
eFiZ6EoTOKIBJ+MmXcjVIug40oEmmM1DjuaG/yu/yyLU3G5N80hCGI27Ih6zdlot
IAZXwlNnxJlr0UYTuQ/huBo2VsmwN5LnAO+e8VFar8tu9YQQrM8SPWm4IwMKxMb/
M6HChx/IR3YFgPeV3YSgdXUBFfk7Af0rvP1ZiAHLcM/6mBnW4u7FskwMqDNYmQEn
2u4OTZR41IqCFimMlcyNCejSBa9+phEellZUdUl1XDCZJzIjT/sE+0IY3QXbtEOZ
V0WiYIl2rLtUgKH6b66LFU48jGDKpERDak0aAcmbZ2Cf8MuJTUCkMb1tkN78EIM4
KWSJ5hwtAaW0l1Sf5TdM+UdQXAGURlCdo7UA4ZZuf2+Hrxe0Z+C2wDhV6zkreqRB
E7Em9qO32pywv/9CqZYHNU7FHMINBmR8Z9DvwfFYHQPvJHHdHG1MgLN+VO+QGlsf
05YgY4QHW19DwGQjYfXwGKuy19+vfnc7SkWGtMF/naavo7bnL49sbsCH99KRJwdp
9nboUweQz2qrD6Ajz6Ze/h5y7R0VF3GvwGCNW46A56ZGVA0xcF9eiGkTGCvW22hJ
m8pxdkS3UAE3pvioUggPQ7N1ALBHVm5dezIWAxutZK8/WWBW5T5YNHVhB1Oqv9mk
5CpZPS0TPPnAwIrLqsbfAs+r89wVQGGsM2cuA0PaGzjbflDDIBIB4bJm1uHfyEnl
KFizj1p25lTXoi17SFemjBeiZ+kNtBKqNhLpqabMoOjqFUlKt1z+2WrsI7NtfD6Z
hEhjk4pFzIvmqqu1YKhd28YR/5jLZLUJAXyhw199yaflAvSGWeuCHRbDxTuUnjL9
JxWTZgnZJMNt94mnjyMqW1RqfzxrS+o0LAs6UbFBA25QaHymFXhFI2eGsfW8g+96
Y7nSmfle33+5qv9UqH38BGrV5Om6GXrDkigwj6ILhMpy01bDJsHFiSsFTBrj0Ll3
mYPmt1drztjYkUc0Gsh6TMu/BjBnL0sD4kclRHK4iDYVb25lYFuI74Yj9yDtAFo1
q1Bu0E7Z5SxPdW+YYwjBcZfrF14Tx/IFqDZhxlxBbKLZBJLbDDoZ5wjHYZaVIKZ+
+cjQnUBDD0tSNyGPP4pUG1eDxkMsWGyrA0FHPpyO+L6y88Z8+UAPTSeVeNeqYZjO
OgsW07BnbRLiMcK7FAVzTTJ8SeIRZC/i+ZqFCPC6h8Q9Q9wZmIqSt8yXMYNmcWin
ATFP+nNsUpVGvzFI7I6sXDD+2KmdAzPhPOV5ZaeUSgbCjbBdhb9t1f7eCjUBCjGf
udG5M2UfysZK0y0E93dg8xgxVktIdb/SlSBBoNcI8FS4p+6XYCtO43xqi9zhTJFs
0KFEWt3gPEUmk/pD55i3/azvywiX47KyBTz7a6PcgfZvAdr7uVrrRpoblDdTISdh
vHRrGrWrmJUIJGw7f4cq5P4Ien5ywbxNgyti1I9zbNDBdIv5neiH5EIgk9xlpLQ2
laNI2l8jpEcLNNry/pNzSMa5cvlUQhIEtUaiAp/9Xe9sDz4bxJ/gBIdWdlEEXqAW
6hMHqrKoznpxiS7aBW2VdUXA4wibDdTPZYo9PvgDy+qJs5q8TXaORpE3p9YtV1p7
xO+8EcqxroH4mqCgwvnL28kp+EwpGUcK3vh0X+JCPwki0WBnFF2GirGowJ8Psi7a
lAjhjL5yKa4b50mdiGoKVjgHE1qbh7HctqIWl1k1cfjYc+xbCxNZTqEo6+Bn68/B
+BF6+b+CdAn61G64K3dwDDW5JVCUA/rtIGwiHLvDHojNo563v9BsHV3dJl7LGS1Y
VzDG49SbVDdAnhS2PmPRIQfAIyqS3kGJNt+RGFpzHYjOOSwoVkR8PWGbDI9j3X2B
MVBjRwSWhgfSUqbJi44nDXI+zimlaG0LWX++fEeB3ywxQBaoSAlN0aPbvoH5IDNS
TQ2DtI5zXfh+YJq8dl8R7AgRldwEUN3bNkohCSt8NNp2RQoR1gU0jlXGI528i8It
AlRXoAnKsK41LmdeyKmlFHh8F7Kpr9Nr1S+S3sOhgY8ktaA8gTUQ7rLF3+epGz/1
lSPdzRLeipJ7jMd6vNhxMZcV4c2G3PhHtxE/NOuEYOSr10NuXiGEGj2iIzeuwzPJ
yhP71Q7DJu2IOyXPRzBgiC2nndzziy9fNEaiFw0hdH6+lvCxcTdZobf5giUlp31P
aAuPKhmLzr1cqlJic05RAThVcmKMpvi/hFOBvF3cz8DykNvFtD8eRhBTBGUKSWp8
51QPedB8pTaHHljTGmoPtGHmADTtp2Ce+qJrY74uzug2hkmGyivkpKi64Q6cyeJI
jDJ0duEtmA44W0wFJe69FpwWN7cxHrLfEeJz8B8UTzmtWZVuFvfjRFe54cKsujMN
Mlt3o2h816QP9Y9PClgtkw52nhocZhPehKIcRzK+x9gtziFKyp7lP+HdyfHdM0zT
XZS0s0gUEyCHZsG64LQjXi3tmzEQm2Bxskf3RJvYo17Zb5rzV+kWGogEEkIN1BzG
V2BKaZIZbZlNDq6Ple9r7YW7yWwcOFHSXALFsjlHDkGrom6s0XOdSdyLzmLFqVvM
Wg90QfB7osXlUi2d5aww96uCoBuQpieIE8/xqaYy+eBqGyiUiA1CzxotNVjwGtiL
x4XpplqD9jjY2eeXjjvfY4SWvRPcAuy2V0aYVzWh9gpkScme2K/AnQ7LB49m6SKz
4WX7RmgRrjKmMGW7KMwriJ9PFRrmi5UK70xBISp+8dicGo4q37mGQlRxBTADQnLW
tmxQSt3YsoD8khJjGyGAPptDDxHek+spivHdXwloZGLtr+O2r1xMaS6i+AO03POo
zUsHgiVa3EeduCZKYOzE3wJ2VEkA23DpSWLHhVACbMRo8HssMG2K45HMvkHsZrPl
lPV32PxaM53idHFoLZagQ2a8W+XxYtI8Z4noKcbEkaYccCKfRyDVTDA0XQ02l7CQ
8KDz8/cBcfcMCX/ek+x21uf9FAYATJ8/TlinO18nFBAxd3TzW2Kiujs4xjrsdsJq
ADfAUPaEpaNdXo/Sq6xwnExvrgvMCdjcNhpalV8+fZhpB06JBDBFRp7gjF5iU8XB
6JbcFR6iDROnLOu3yj/DkOHZXvfojgp+hW+IMRaQBWpPrytQqumMKg4KpMgjtsxg
oOJpQp9bTrYcaUIQiTPbtgcb1xhRVfIbczeey4+jhshTQa3FxMQk6IPLFt89hSOM
TdfA/FupAwcC/Fe/AnoPAp/m031mTiWfFyupzyiJTuW9fsWYLiBqPAlCayJ7KsS/
ViBg5HCV96Q5/0L4fPtToaqcT1D9GrZpPvucsV7C92ahbpaURZ/6QBxTa7dv3+KF
4hDml05tjdfjOO7mUujb9lUXAAKbx3vmDPBJ7wwntrYE9dfZ0/lEslqg7IKWKlTD
L0fxsew4OPzdYlWogXNaSrmoJW4JyyvLS5BwzHx+HyojJuKu767MKJ4pnxJFoOub
qx/Dab9YiTx3o3a58cOFKYufbvJ66OiNenZZhBa9ZccSe38UNDcu0gZsW11HUOGG
D0+pa9biAjB3alIAfaQpWa5Is5wiRZT7FoOR76zKrEoTW7JrPJfeFDUk5QaFZlV/
tWrP65Ql7prnIGlFv+wFkabxND9wM+kXEDNl0u73mIiNgXZJoK3mAe1/XYCJhKKW
p5ZyhBbaD0l3f1ylOHVKo4wkPiufUtkcoZCw1nDXdmbTYOllmjBiSTiyH3JAaQpK
3dy99WKUWR2MaU1EOFUD3jdeuml1J1yHgWbDHxrWhZtZDez6pXwf+igS5imyIR08
UFDwKLM7guel8dBQVemvmBjB0ERto2I9lWK1jID6IW13j5mEOuUiwdjEsFd6iGVz
37spjLf6jaNsz6W3aFCQdMqE1XabtN4Lt0cmqx2obVCqcKnLS72hSgzXq4TUtQzJ
NR9jMgmHIh+HH9xAyGLkwG+9x2SjQanfJ/8Tr6p/JaY2YcwDd03HbQDpTz+4A+AR
w6nlmLMJl68P0TTPikdFo7JrWe7MQ/8O6dyFX/mK+PdpDK/kvcjSvmI9QIPhH73u
hHGzkBQD85hQ6H4IloDLXHG4O4Otv0uxjYJOr2YVj7lDggucO4SsgWPe+DCAui6Q
slsfHktR5Vyeeg9BTPfgSM4pYq8AKOPpjN/qdbJLj8pZi/H3SO3z0SBaPWk9NldU
vrutri5He8S/tSZ/L/dsL9zwnaFYy9+DIhnTivq8IpRVOs6E5SczO6y8RWQnVLor
xWVah8dQPSwNpW9BY7L5fEZHtUw5Vw3lm3FmJbglBOrT7d+qzoFGJKfTLR0pkRz7
MH52tBzCLiHuAGi5DVdAnuXA8cPr7bbKRQbI89UhmzcpZcZ5zUahac+4xSYiA8XW
KIB0+9RyKEWEddymJswKMjDaMOfdXr121Hf6f65rBKzS4TjPxIduUrPHhNs+GmEd
xs+Att7O4xgWa60L13gzCgnpUKAgfbln6dmIgZp/PFyQJ1MzY28bm+rMBDln/41R
YIC5FpPavkr+3HlquU5G0DR0AYNycVH3XVespFnfLS185vjYaF61Pzsud2b+oTzw
P6L8cMNQq6XgP+em/wpYwzcHqD+pPmq63Y5d4eEnFEVlR8hfDQELzgjOdOBjIRfC
GNwQLEXPwYBPNodGtrBduubLU8ZBc7+AgEFtkZ99ZiTsnGwneHxOCuTFrgTqCSTs
Gm4R5MRPoNFqlN0dr3/tMZOJ448taOXiz6KXKqkHNxe159fmEXaT08Snya0coz2l
412Xl32idACZGQX3Dk/HDYSso/Ekh0e1tROwUIR4Ub5WJVczHTphbDMsi0GpIfX+
xI/dRp7P27l0YZ99YyB6h7iQe0nsAM67xaNQJTouBqUGGQEsVx3SRAFZTq4kX3Cu
BfQTAFz3lcLwwXCTjPaa+fD4F1NbDpubs9Q5XhwFXYcw0WVr3ivMzQkS00JQQels
WXwBKhaE18NX5rbLMcwOzmJxkjsdfg0ScsOSyszLHdSAG0+RfbZ8OotAQLkB/1vy
10+z3OrSUm0oZ3dNYlSRNkHTSdpcszHUfrtkheZUr58YWVAnn4BCB2upP0wsy+fw
CQaFLLmsy9viOVha2K6K+IiCie+MGONiUSvM32CQwO0PT5FZsRrt6oyZqCSqH15X
PT1/qjxsDq1aO8dj5ojo/DgokoFXwKc+x6VMVgk2W7IIbV37VlfufBudhQLintYu
qgIr7of8FQkw+q+K6Z+wnTzuYkjoaodCbqpfZp4+tTsn0brjQ+KStDfd2xeIajzw
sqXpFB2rY6OI3lNb14QJZF5CclJqtqwaLNDfThBdzP4lRnftAHPLdjtHSOrUT4SX
ydBBcp5ncCvA/GAvKgDn8u4WC493ujxF63LTQanGWFbTOQ9MKmD8Nn4VE323F1Nl
Irnwh6nSoF65MplwiAOnOYZ/wJzOLlucGEWD07PVrP6VM0N7YJ9+d/JWAwR89FC4
h5OVLh+LPRAXyfM/ydwWSGi+4+AtNM/BOU0nUVDJV8N05HqeP1kY2CTbiIBwej5u
1gJOZqhrAYCg/pYH4GNWEyd+4qy+C5KSW+vBAxkhWclFJ5U7Wl5C1MaeWcDGcPNF
E5mJkcy2A2Me4Cv6LTB4RDNPSTvJhc3Z8YWPZh02//TuDV+Pa9VeCP1ZpbW9wNf1
tF41EMg4UGlQRbAeQefvlBmgucmq46q9N1x9nPzqC2nuhUe5hAMZw8owKxhElx/h
bHXGYhY1G2RQnrrapglhhU/wORMGLWrqd+BtrESo5+02OfxBM0YZbF64Qg1+Z4jp
rQ7QFHaw/2uZ4Y1tO4z6qn6y/HLroZBFfO5jFH7XeUVaUh3N7ubVtbK9MRT3ErSD
+2O3yW/5tLdQfIYCWL0X+OHT5oxDJkWHTi/qJJtKV/3/NvriMGVN8KVtThHrSlC6
ZbUlL6LMshHjSzHVbzs/Ye0nLVVchYYWPYWL/1v12RszTn2/n6LStRY2j6o2HBDz
fQ2Xa7ikbd9Q5INikiQx7566X2H+3gpbDawRKwm07OuYkwN10HKdq4js6N4z3Sl5
BeOKL+08ZyyKOwepHjnF4E8OMcJCaa88wUwadqkwAI3en5F69MeW5qDgepQRkNC9
aPMaQFJRi3lw9wuA6yv9JiwxdlY2sdyuNwNlQHZ1+CjXP0iNelXsH7zY3vJQgcTu
TxUWzWRmLAAmDoP2DEtWGrkaW3bvN2zgAGuTQaMoGF4WDfAKZyqG15anZleZaTcR
9UXzdUmR2PQw/hnACGfxFlrB/odFv+p/fIet4deb9/LgfeX4zLDJMqTxwVA7pKbo
DyY38Xdb6BcdD7HgmKduLcv7bwtMOW2ISVGbZ4jUnJenYqLOVFhdYuG4J1T08tPM
aq6rM1yem8IrolSspel0JbpjZpafnWOabheAyMm3UU0H5MUwdmiwbV2/hMjqhJe+
01NMYQG9jknyAw+DrDe7QeLuEhS8nG+cdPuRl2j6tv3kC05Ls5cKLZcQLvMkZ393
t3rznUUz8Q0Xar/KgxHB0ECik2qTF3XAAmcZdj8t3YzKniLzLX+5vUJZy6IW1qgS
eYfGVAAZJCWhhySdt9TOE3zwkduU4uDikKt8CYUOQFMZnRyFSRz34XIrc8w70cUk
wvICpi/Azz7bp/+Kdn6BGMXZWjRDRKfFm4o62drQOK3WhwfEqpGBJjL+GZlMUkKZ
+26u6IJFmTZZObiMolmcY1Jt7TuLU5C+8Sa9qxVaS5w2pJ2lpM/5OzMSYEklgEoB
4LNpWZxelNi3bJ8O690JRrbW6FoYwwBI9SF2fGWuGieJi5asDX+ShzekTkYuX8oz
vBjJSXDVkz8PlY4/uZEPaSzy45jlxKfvPF5Y7s/stmQeCYx2qRcaSDEB4c0e/OUH
/wlutSEK2sMyyxs4HP/PO/cIo30CmlwmnrklYjaRKypexN9nAZWIuChQVF3fFXwd
jwVxDKOFkk4R18tqgKV2NKj25STWYrsvzHJJorvwk2B0IUuhzEEuJIrV6KD6H2qz
hhwvaDSj+ITXVGw0ZCMvzqxYIKWbTOKK6LA5IX8zgRJ901PPYkn8T0nOumGvRTJ8
Zf2yFECLAwk9nB6ZqXOq8re802KYzp2DWSgHbTVlBOLEBZT/i57+E2TTjr952ku2
XgMmG5IkgvejZbrJoEKP/T7hjbibVGRb+e1862p6M44ftv4Pt/adEA54ltVAB95t
diqLjk6sipG2xqa8QSmkAray5XS6tF2pLV+lzK8psE+WpCEA9n6ES3ZgROaiz6IN
EPp1ZQ9JhiaLaxYlQ5G6wfClRaLZeltgoq4q2587ROaaldOKeTVFbUcXv7tVUYLT
M4cHQGwPLOJK+OBEXjIHVcTb3fcEHWuacKXYmsX0X1RgFOnEIzIt+y3F0dRZp6QW
Jlb6wfbPd5b295jF6Ajf55Ka1Mqqf586zJ1pW7FqvzNWWm0ZwyjbKRgtLniuYKPz
V6xBUR3JAWuUCLA8MO48ltMi+oISoiyEJ+0BKie8L7d7MOmQSLVSDlzVn/DoDsDB
am/Fr6dl+jKPxq68t1UUJIoxIcYo/YaLjQ/gXnbkSyTT/TYvInmO+GEiYlE+clbj
60MplkEle2n7w2YBYMUVOm3NMvb2qWhlzozDZfH1c0g/O4sEjmKJxua6alIkpG5b
IZpn8GSA7TR5bnW+nmEq3vK2rJ/I22TNCKiQf5ALKynDb8H0gWwjqxrRmUNbhwvc
xc6mmdZmFY/TI9pFovmGWvn3sH5ZmOtIeHtQjHLXY9uBUTrXiQkV8KEUFURnKSO4
9qbF+/fRWvF2pj6kzwsdffxVYqQ/wCceXArEjNxZiIAx/+h55RocQybcnCXAgsYA
1v80zIKodbZddpyHdQojjex/9h/UFea1OvI3boAgzfT1gBB4DhivfE1RTmL85EMw
W6K/WP47DgZ/T0coM7Yf/01Vriimh2Q7+JUJinEatUC8xairtvGb0w4sg0t4pglk
rc/1jF3PnA5GNXXSL0kRl8Rq6U/ga8W0EK66bdHuJxoSBaYgr7dYZUe6JhE5sk+9
JP1m3MbPU9ugpceDlTVERYtuZrxVnKEx/vkZ2Nht6zB6VSHQ3Fa5HtRJ5WZ+BADV
Xxd4LBiP+21o3R+6A9cDvB8jHyybU61m+WTUVoRsPdR3tF4h8gdXM0fPg2dzT4k2
3K989Stx2vGYNnWN1GcnJmSpQXProTUK79j7Ij95rK+bELa2hvMpr+8l41afyHpT
aGy0/K8/2j44ILyPw15ck9R1ccIWn+lWdJmZsb6feu88Z5VMujfoZsw+KGJaeS+v
nozZMTUHqAgsl4Mc2tmlPq9Lb4TmRmqkNuEH9uHhN0b4rLpXq2RaAcmRWxnCAKa4
Ym1Z6fABapVwf7SOrDPM+S7XBSBHKQrlHm+ZquPdmWT3nnT0vORFed3maYHDnZPZ
wsJLNkSeMose/eMpQSxve0v51nYJIG66DMwCTrXLNa2Lat7VcuJKHV9Mt+9WAfMt
RqQX4PNt7p9a3tyonBsAQalZ2HGsI39DimM28dxaWD6ge+18SJDp+r315WuKGam9
hU4SkIT7L2HhHUSazc5LPilvT9ehrQyPECwzJIWAvR8++LD4YDsVJ56ho20+/Caa
GFeZ8ciGaGytwTIB6N3tdSq6WlzlN+Ary7ZplUO3diN4UMcdUzbyRiAUCjn8FJHx
X44l0b7bzEbkljWEbqzNYzavG+hyAYiHoo7jd9aLabpNKx67Gzztk95oEYio1zqq
jTDBRKtFBtX6W6wkcxuSKIjzE6HGZlVHnbIy0HXC4LKD1SgNAAF96cXRjdzEjFrl
Nq/WTnhMIeSjYyrFoBtSBGcV5H8E1uMDQS4SIp6B23ApisXy7VH4lHIsdovfHY32
hmBL2DYI5nim152XX73DN4Icf2H2q5esxdfXIUkNa02d+ZGDGYSfK6ibZ7eUNHms
oH8qJ8Rpcc/3oPaIlVdrg2ZVd9XzHU2a7k5idnk4Pe96hUEVn1EfYW/5ntBXmkIt
SaL/WDcnbySK6Q/eig+3kk80esqMjlHupHq1JTs8U848qnIDBC5vo6Wa+MCM8YuL
Mki7joIFysXQgj/wUN+EoMwEzDDIBnjDRXblDhsIKLbkHQtRwMvrAYAaUEki1Ie2
m4wJ9oixOx1NaAMpPvhzQ1xUonyV3NdJkQAuQyEGqWGB8HSXZg7AFuacNsSDRc3C
cJ6gmjKcAnKNHiZTma/Cq5+awRaP8G8yQpFnQS3hI3TPAkSGidUSXjn9EmM9xknE
l1ZXqVFR3aUapTtxpwJJqUFeYrnYroB623ZS9RZTn4TFydc+ozmPEZSteIwKznJx
NGAR/XYPB4w7AbXre+m6jsMeVOx5eRZe5T7TV7C39Cj+6DiHoF8yYjFPssB9ydkN
8KNVAoXN5IVydXBJHoLk2RDISWG9ulxTkkASKVLsK1hw4Bor5nmQTeCS66wKHIz/
m6kw3/9zdRqfUzAvsa3c/we4zRZts6geH8uY9ScWKFcFKgFdJTamQQQ13YIn3M3d
Q2BsXAJtFxxBOuUWTk9ZVdFXX2G6TPZ7BnbTo1H3IWUu4LG+XVAag8pqfdOCwsLj
1du35RAw81dNa9QZXjxz0mnjAxAsjBgYGUH5aBvb9A1iZYSD8WfNw7k9iCyg4yXJ
FOb4q5TgF1vb6FU7fIsUrqcUMEYBgbuU4QKP5yKoVW2J2StJbcxnDx23nico3fPw
R6tdLcSLNQ+YpOgBSpNvKQOLG/iI1J7hCTgVZUTGVCLhgkQhkKkXEMawzo31fJVJ
jpD1m+PM3mffHTW9/MmtOc7JFwy7cLuhsdC029ItQv2unBihPFfrfnrfqd244KSd
MbmjViQ9mkz7JOfiZE97IyBBSm9ga2JA6dy52eETrZEZ/S65g40vMijYRe+ztUv3
9TvUBPGnLSsWtfX/0toZV5uuZIFrWqEiy4g2kZKDDt0w9dHJVpWge02kUb5YCgqz
vkhUz0IeudGWUrCUZig8o+PIgexCpgNpFBzrC6kg/XZDc3aTUtORKm3EibmzI3+j
ttwEbf2prmr5uDoCe1/zHHyAhhjRqDNeboHkxSwtbvXJJxUG8yF2qfHRR6ziHILf
7AlXfWmryOCYi8ZkCREkQZPsKKzIJMhYCBjs1X3sarR3JPqxv1jxCfe7D19HzVjb
Xxvz6w729a21N1JXYXbc1f1Up/juMp90WZiPm7QqRh6OjLn8NwEEnZvSk9pKz1Db
/fwYuAk5IR9NotgJism11fZ0sOfkevwgA4cWXDhiPtRfJ9cAu9Vr96RIxlSqTy21
4akONEPBdfc95lDPxmz3O/viW1NycJJHbTfMIkeI6MLjnaI4BWefxDV544Uc/YCd
kjhjhFUEdoDiCcB0DhfQL8WJSx6wLxUzPMYlw/8IWVIgfcPVpO2PYf4OM7Ilqy8e
zTyGXA7lg/1Rcjad1B+QYW9BLzarOTebUuckAWUzjS0jHQwtu4B+dHTmWv+DBxI/
zBh1qUMdjl41b+lHUxM3ggzqZBe+svh6ssNl/FMysPXtBXZHx2eVEVm10p5ExuJo
hMV0x4wnBWvi/p++dhrr0IlZuS1RZgN0/O5/+vf/gEmoNllwXJXIiNl5rFHtReiy
jliEvryLG5ND87C7TIBiJGwuP5BBpWTrpXucPYcP3gt/KLb9jckF0PYNwEI2D7hc
TcvUU5yrhX40p0JMLsAor4QNpZONfiYjynTCuJNc/Rl/Pn0RrVp6lpFnqwP61JlZ
5l6Xt5TV7NaehkGIMhFLeZ/jZbs4ooCpHUrCj1llITAIrzCziDB15hPDXDTib2Ao
NMzIMxrBgjHm58d9eFQuafem5oS1im7nb72TTQUrcQI9Trf7jlC32/Se2C9tmPTq
qwBoUdTaU++uj2H7Oi8HkFzl7U/nF9zb6aa+Ho3iREaHABwxX9eqGMHeOlx2nYwW
lqM+QiO3PkSGpc3IGheWA9ygNVAiWSLVIFaoynAL++5el4+QgvxXEDH5/Un9pmo1
b9H9PLeaaEAEaDpYobpfF6+/AgqUWwxUFe09Jjch79fgi3Wig7E8P3vGLRhwxLnE
ZDEcTpk6MI1DllD8RcsNlojow7SRCa3vQVBUrW5gKtcJxvuvGZbIcsnsp6No3G7p
PK80FLKH/ww/i0xTIt1upgoYtmZJ5Q51y2RZu2M1VPzH7sgsmRd7Py/HZRM6/hOD
BrGMNYy1S39PXibxbjJohfP9yim4BjvXa5ET0bnMM5kzAdU98eCnGr+pG/hIcbUS
ELDbjUHO6CsTT9BMZ3ya+vbDqNzrD1r4JwKCVzaKjPwTRPHYOnv7yd+QBosBNlvK
grEcX6LFYCBKa2dVS8f7j9dBEi+gPIa8kQgVYHcoLPG8Wduc0kkO7DI4RC49p8ce
oXkEMvjv9Hc/99KYdgSYtzbdt/FoQogAuY1OD44KbMwBm8gIxhEjTnfXxJy1OH3B
TtJoeCNwhzcCvyz4iyKuzP/qIaPrxmSmASm4qhLTIsmxWpMUC0cRIUGupVWZYIQ8
cW2PQejDjvKpcRlfs9XqnVTY5Xl2CL2TSBcS6nIBMO+iomHMFYCNX0/GH3NNE0dZ
/MlBzKDD9K6zaeTTZYHrUo8P0LnmLusQVB55ihwyely5c0U8SI9OS3Mgz08Q0myg
CIJoLPWlkRWP9fHu1T80StxneGBIRxrNsx/vH32tNDj+FVr3MkXQS8L9dSv3kz34
WmnBCAvizx5dsWZJv/pVdDeUPHq1hfEY+HY+8c5AmUnUBV4OVLywMwA7rOslVyxG
E6B7JF5kKxv06KXzKQnUSXslVt+Z75zyFcB2re3psumf/OOAy4i0RWRllXWQdk1f
MLggdUpc+snAkI23ENYLdyfS0oTkPX+6JWC1lJXGzRmkPsdU4PEOcpIPWVDUu8Jr
zN3aHn7Z6Gs3e2u6Fm4CM0tov/XJXcv3KqjyeWxodVVpiJIVQcGP4BHZFBX6/HfW
3p+hu8UTBcv7tdpAYKrUAtRhoEvNVqyHGBqzWkn+Eju+SPVVYzNS383COCT+tr+M
r2NSgV2Iko2+Wr0hj8rTzu4rT38WtxHDIzo+o40U/BzBVrDcJil3QRplAu535XRK
87VTrIhmKyEwD1wnsWBb5owFSDoFWVnd6LntXNEav8YmMxKVon6Q6pggEpZAGWe+
15Tf4XN+suqH3foMv7yJ5NQekDjzhJ6+fhnpm0lCbf+TO2DAPSA/+w10xOP6C5bb
Gfh0G0zFH4WiFejpu1QOkVoRok5eEF8Aue6Cx/u1U+XqQ4ArWHdsxrXkHiRZ6au+
STzGvJtC5OHqnFszJKh9BILCE4l3Bs5/Z9pUjIYaGEbKoizP1KPoIsZCmCp99Ebl
XNkCcaPVJGYxjLfW4qyYSVks5w1+/R1Do6SBkGq+DXbOESNC7jaqT1HKIWsRRIdh
pVJVITnxP3N2YS/DNY8m5bWU8hea5Pd2POchPvR769lEIrsa5aJscpYdJFwJb7YL
jNq0mjAZkmZyS3WDaB+6wxaqaUE+1F14NFELb/DAXjSsL5IOCruQVKUpDk8T6SCj
dV6rYbiVKRf0++e8r5bQJWPln5cg6auwtEhawos5rHoTjYwqFSXJjhBsXjvKcgT2
uDKD0h28H66NFYEafKJ7rzPs1Mzf9EeU06PlZoTg/JbJVSI7O2oKjL4MLtL7d0A0
gw7ezw/Y0vN5XeOl9Af640pcGoEMlIyp1+Wy3Es0tOiC8rDYiFe+52cNdAP8FTE7
d5SvfpgQ7jTxAY8B8IHvJefG9QulAKmE8pidQr3AnYZyjSKg0Qda2jeduum/NacP
RmGR7KfWt9lxVsICBmVLRb4vRIQvM/NOwI/7xfdc4fXrOOLz2U+/rXxrY8o9TNct
fSDnF1hJWI50ov+oyvPhAlch+SPueYa62UPFMiYJa3qYNPb3FwyFRP+TAPnFrvDn
vmDYyAmIN4PS4LCBvyEPYKIoiarb76p7MST9gfi//S9Q4HOi1NHD1BPOLtnodJxI
mmdIVOumj8ApklF1AwoXSMxzL/ySQ2L6cmMm3RPKqRP3WeNu6FTwUyfN/ymb/0VX
P7E8DFrL2Xv8dFgg4hue3tYRwIIleXGDeUnaJTqPc8CNXYeYI4Ctrj0AtC49usjJ
aNehJDdlmfDPu3AQr60P4H1I1eKy4qwuwgXmHSkygYpMK2QZnEHx3JgfJGZx41+F
0Z1/YMsDJq5JzvPonGa2LZTeNLZo5s/EwbpcIKXvmFs4vm1CdsM3CujdQB6REtP4
vsv/dTsTi60c8WmtrWVil95AzZlOhsmbllUxAIuGNZJUznck3/396O57lPa39T7I
PTIuFfK57eANn3+bKnzTQLRjhh6gjvHU3+SfSLJzHjuC982Y+i2WvJThCHqVKmT5
mRGx3oz7WsDa5LL21ZxogJEuJknhYDzPyysC71NK8SOazi4t1sEKJ/MJ/oiji1TL
IZVFfI+Y/c7ffT4LYyb5xLQwC5VOndcelyUGqUcyXnbxujle0B+trldLRoweD4XY
qObhFbZZjmuZi9S+t7HUqUh6GPCfjQPlzcIqMRZKOLx6zMB27AOLJ3zs94VezWXW
o8r3aeW3yCS2/+MJb7XyFEvXuqLy9XyhMKAYfU0XrpJZCmga79XDj42iEv75UW8L
FlXd14MD/qaHJKGoCcQP+Khihuyruty9Sbvq9eiCxxRH/SFCDHCUH4Gc4U6ZzBdF
rBo5CgOqjBE18tmA9maFdZeepE3TxcxLzLHwzN2js3uR3rv3VVja+7sFYCTk5G5A
tIjtZH0zCCIYIPyNUcDWma48Kkhg8zThYuU40OmyKqNnVaQyTl33jMkR49GVczfU
R1no02sfmSEeWkNOYrbz42LgBBeHwGpM2NqaLI9q1eGSwKZMsp3nfx0l9W3r2YN4
KJuoC5PjjXJRZouKyXpE7S4v9GmsxFECdyi/kpMB4T9M9dt6ifW1iIUNKSig9lZe
8kewqHVCdg3zCZpGTnrIohDxYydITvf3HubPpMp36+nnKzvILH1hCCY9eNZXOelG
xULk5KPIVvRlEvf/q5cgPfESnFP377VVFDn7D0CxsnuS8tzPG0+1oVrXFuvYWCNj
iWArxI2FWeLS9aAeZOr4bOEfzS5UakcKwY9gCTi7Dw1YmpHb4I1wtY7Hu+MI3dZT
1fa5eMumBBSBrNsMONZ7cr0D9W+hADOE3XUxZ0OXyQ5NbW3QqM0MIzLUPtqIUqwu
cNx+NvhKpx5YjCEb2L8TndO9N+BWS1AoaYJkoE0K58taAPrOMurCmF2snBqX2ltp
I0InWYhH/cYKabhXs6lWhsa6IlZX+6GGj0acn4TXG/vlJqVIY4B58/xkcWJXCug5
Jzs2xibD1TUjsjEquWzfuBaj12PadBMLhcmuOZmxgHY3RBtnUl+uUMvdm67Gtgr1
PX5KqC9yLjE0T4mfcHDU5/82kgumo6hZTfhzSLOuD8xt6KgQzUDuwjgQaXgHUA8B
/HHAxafPeqH3x07EKIJrxHbd0/DzQw9OdTk+45S4euyCRsReSUlp9QnEQzDfOODJ
KBGeAmo9uFlJC7iUKxLJMUO+aMBnRLIPk7dpfmkfUl5Se9x9zmjyd0yYSk/p3lbL
3wlEpzM9hXCn6mkwCGIu4WYmQh5aQLSw6/uoh7TtBDhAKqSkZ1S1SZhVSIVRjWsW
06F1lmam3bDXpQexCVGB/+wv32fdTweWjOpp2uKwVmOx330i0WJEphVwG7N03CiJ
c4z5V1mv1D67kCeEVKz9oR7ePlkMI743J/Ffu+Xv8kqyb79uuTrB2NkxRdfKpuk4
GEGJCmhVX9hbROwLQCZ6+qB2u26EbsJF/oz36KcYsMZOVDJF+kteNp9RQBIanFVI
llFs2pre4H8XwUcq0TD4qfmyLZpEZOunKDgySeAO5CrVHy4omVr+RZtasV3dDCjo
TFvzb0ZliME3b6aJ2eQDaNoSIcFGxuXWOYN34zc9Jq+LSDRdaxlNowe7quBOp2q0
u0smyQgLpUOAdxX9XPc76m3qKLJSAvbQ9tOsS6uvRL6wEJne3X+elyJbcwEh5by7
o5/VUgV96x1zMouWlS77sxhJRhFnCgJCxd1d8FPL3XLWXFSWWm34nSa0XeorG3X/
x5BNT+gGysI88b3/U7u4CnofAiGuI66gEws2bl1ESve+TFPI+4lfydXr8eTzGnIp
YAz1tHlk30kiefl3w0rDi+h8wOZknV2kPUVY1ujloBputGuEj9yTL8sh8nzZ38vU
wAQVLyJoAU8icsuorLVWsG/guXFY7Tqpjdb+UpWDSMjrXIVhB56+YN24ghdt3LCS
vfBsU1OMnU6k2r2hmQ/McdEKmdqSO6Onj0kN6m5EKoFrH+Nz6TfsR7EFQgAA0+PF
7w9Lzq1wSvi9zrzt1XBfBoLdnE2Yes3nlrx9lgsZLRii+Lr8VrHTJzUFmFFH+5RJ
oxeSjWrx8xCB6QNINOgnzVQ8gmdxW/vb6jeLjOMZpNjUEvQoelIT3nGggGOCAGyD
/DcBVrMD/uvn4FWjrdyoPIxUMzRg8OmztV9/S0uQYdwPA5MMOT9poN5nglg/0P4O
zktGUQRm4bd6iV50zbWkCSJ06GPD1TtAB8rS9J8GRBjzNgO9F+O76A4CxkV9D2xR
EUtVN85OtvMNUKu7JH5sPGE3LZoG4q5FXkZ5k3XqKvb8AOnCaAZr78t6XwhNrGOw
CkVX0ZggoSXTzUwNL9AGf3mq3aUptYFcU1HhMrgtQ+RRrfWZZd35ZJVqX5W6D0vR
5b4aOzYvPZwqfI7Ge+rH5EVQfrZd4tbCDCs0qgpUoAXKSIGKeAetSSuuOWbCO9uo
tQdCE2TDExU4nKsBCJTh2vyGrTy0vGGdKP5OD969l4s=
`protect END_PROTECTED
