`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wZmoGfDov/6wjEYGMHfheUiHZDu+ne5sCmumH6u/JnglCdRuehfvW9D7DFNL/AhT
VvOPg5rkBd7nb8mcOPf5KlRb6gQ0B8+5YVQA+L7++3ruz++oroHg8egg7FqQpQEu
IGENfNR1YZDv2K5elptctkxTNRqfpKDPLB2Y0Jh9rfD8wbWq7k3F3418bpCoRnl6
S58JtrtWVYeyB8L8yMfsu8fQQFqH5BXKXElzp/y2NKiRsQn5GE0yWkeym+aatpV2
ZnaVxCcbpUPxXjGE2KwzrQhDAechBptB+uq2t7FWyEC62BDHKJT/gCll1hqKBxQr
+YBmIHa6ObcDUlpqb2WR+Q==
`protect END_PROTECTED
