`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTWLc8RoPUO/4idMprBBV/Z6yZ9VO84l6T60DAmcjd0RKomAK00k+KIeF3mbbhqg
OllIIySBz1wOGVbGqpbove8EinsCRH2SYZZzZy0A1U38PhiSY8Q9md1ROkvoCB9a
MVzY0oJvQJCxVEox4qpa8c8qJo37lCRUVjzQPl/5S8MU57G2cT+Lkkr0wKMAri5J
vhjOeL95327IbNBj0WI7JDRogp+p1G5hxy2/IIW46/FaCPY/SajJ4zpdy40SzAlg
3htt8qndNOv9Gnz6IcI/LBTYjfloDyaOfxG7hSi75k39ft500IzqfSepLcy4mJhE
6ZZh8GySybkFL5++otHBgDWZaMr6qPKFgWAiRwbs/GvYtYJrYWnHPbuMY17y6Xh+
4QJB4ldDQLMvNPXhqbxxg9/fxu0UsJYM/+Csm1S5vjK9CUtJFmitpCfdtn7dMLxR
avdi2kCaM3urwQqmUKbOyMDB1brqWj7N5lZHC4RMhBej2fWHZxN1stuHNoyvw+fU
dpoKyPFeQHlEw4c1wrxthWJX/Z5iK6v5TtkCsSHEdCI+IdFyGNFGh0wKXG3gFEw+
`protect END_PROTECTED
