`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4LYLI2w9aauVtGn0Pq7juTylSxQnHOghZ+L6UsH050hhAO8FO/gCRD2VsPHkV8D
FHBRd81FAYsObGPKtzYcp2fgFe6IXlKRrgZCH+WgE11Poz2H2/KOdOtSVSebh6qr
TvoY8DCJxO6h+rqpufiM8QTm4LvJ3YM5pZrtvH15HD6M9EtPOt5lvhXdNABClRWW
tEgDuvCCLm6FxYHKKdxJFizSy4Log+1Lu8kialnSwE4RapmTA9vJ/63a+eCxltBw
f97C6a6V0jZoNX7cZ8uGo0iZNWlJ9P66l/yM6quLG3i2zisCLOwbo5m4xLBK7bSk
gUXjWb93WQqOEKu/Bn60t5Hqay0pFhUhYW1Xfhu30uwI7WLuogzYszTMlSEF6jLi
sNjWBz6fBgDpEDwAa4m2oo7Wg5ZaDrcsscLCa6aO20+p2W1sXWsqxC+g+23Kul/8
3lfvVz/dvWnxyy/EctMXioAmlDOJ2wYyPV37GC9tD2k=
`protect END_PROTECTED
