`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ek8AMKT6CGGaiD3oM/Ah8RwnukTnwdWzKq1hVFh8CgoSOIm5nIYOqR0h+G7VYs9r
7AqDIoiMUxxgDPKYY9sCVWZTjz79qfb1Hn2rm56KEBbBnRJznoEwLHXsL591fUim
X1MP3i0YF2Nf1ML9sUN+T+F+gbtcd6kDQaS+2qBotC4ivxCTfGEB1AI9JYinquj6
HsEmPW/TUnS9MHFQS7J/qvwoJYtu+qKtrC/vtRQCBXhDVPL30RgQq0hg5Bgtd2pK
LYgkyzphYIFyJY6CQJBl/lC30NLp73TkGG9BBMlsIDMUkCLDX71OeuQYw80ScpUx
qWAeQjJp2ML6BwrQKkZZ+w==
`protect END_PROTECTED
