`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F8JVCh7XqlZr9mb5RD9ZhaV++YS0NfFOVmTxTt2kSaebDqvlUIU/pjVm8o0UHd5u
P2JmnBp1qd/59acP3Oz5+Qcm4Pkbn2TdNSW48csUk5zARQHhilGRInboBoD0T2sh
QI2uB2+jO3AbMh4gSCZiPJqb3XISoZ4UEQxv0nlDn/quZzl3Ws3495DVPjhvCslw
Vs4YyA1MrQJVxgkfF28HW+xPRWRnVmspxf4qXgyf7gfKo46NBI1Xh2d8u514CkSk
nnKwtYxNgA4KOPEemLSVtcwAGFBt+93qVqp6Empz/ToZLfEKeG/wSY0ELkA2e0wB
sh7Vz/ISAfxrH67pXX2E3OgRD+R+scduy77InRvH8LU/uK4ObrTu2G3kze2qFC7L
Oa+8leHuh1qxphAwCr+rz3BSwk58gd+idNiJQ88M6pkJT42tgZk6QNAT42IRFbJB
nxCGEwyutnqPiQa6eledJ+n51mIPusvBpYUgrMZYuqgVAjxSaYpO/6RQE9kVawnd
BY+1ea/1Ko6jgba1Hr1yyN3Q5OcIaaObxhF6ItEIugalglBCEJBqOthmZgoRWmZb
Urr6bMUoljb/gzzmzJV8wZi1wVXTYM4miecDB6FMZeamwIcsw6yEbR7YI/IxihVY
BeNyLcuQY/6B8PJEfr2o+IsJSnNtbB6DvOFVZ94AJw949YsNFBxEUiHL6B8ZhRSS
ofnW1xM7nvQQZcKFtHm6ec1QKovR5as7uompjuF+Bpe2TBj24e4QX390HADamPgW
jMBMTEHy3Bu7t7FjpkYdaxgqtdK9IC9LW6HpgrNM+BtgaY3D/3k+ZXoFc1Q32Btq
7yVX55hUTZI9WMtXNygsZxYajg6C0LE2BicFbEdIBUtUIGEEw068FVxJZXQmWoDm
pkjt4KFqEFftxKAHm8++GtPLt/ZEzQVN9YQitT8+H1dMioCTEvDe9GA+AoVrXXrN
7xkPWYuOw3QvL8kJqfHt01lx4B+PIu5nmmXUg16GXaaf9OIRXaQ8sUDx6mU7CQA5
yfxv+LvfgAvTGEduTHIIsPiln5B92/3CI+wpPFvkryfq6MYpT4WeLaoNKPAmaKR0
vBCvozmTwkaV4AEJn55jbKAwWuvigkihnPs984QQptf6VzOdME9Dw94WN0GhkI5B
1OQKfF3kj492OLBBPRNY9PZavbSAW3qT8tw3Y+HsdLiZqkA2uwHoTwdyboFp+srY
bBK+PT9juWPxilfwuKplZinQG8sWA9eK2ULecBFyNqrgyYtSWQ4l+5/bgvBbBYlM
y0hUeP6swxAAyNMSUEiDnPl3aiyGo65TJaT43+1h+Y/16C7Bo2wAdssj0XvTQRzT
iwvFq6OHv8EWhPc3Xx19hu+haPjXfd7muObv2KETOmvxHnz6LOvYDGwqgE1XGshN
HChQp7gSoIl7vt1wkqtc5ArTrbsC9Xvg6A5cKJEkx8FRWZNDgz6rtbJAztUvP7sb
COMePSZ8EGKmrEGkCtBr/XF9gEj8F+wJMyB5u0LfOcPHgksBvbsSo6TN/rnRXQGf
qiHlchDC1ruqcnVrBZzHWFWGrW1iOFyO72ouH6aZ+99w1T4AKTTBDGyxc70T+0PV
sGKUA3HRupZihPZVcV/OiyIQ8BFxzCqPviQXLmgAD23glGto3TqIkbFQrxOaC0NG
uwbqShEgD5VTBgH7PSlAtDFDyCGPw4PjgTenWydmfKZJu/7KE52h2vyl4JG2y6wQ
qrJ6xqqebVm6wwxF6eQ0uXZnwjI+eBb6BCtgX5PCuHrtBEvnv3AED5yZOfZt3LIS
xhIk2/AadDYbt09tG8beLl1N/8GDc9MO19CL5yCItlCjyQecXK7juvbyssxjXkJs
uO3pgxvZRBPU4SUZxpzDIfhVgAyNlC4bZX5PGkl4NsSrQzbMUCz7fPOgJL4OflUc
6UZYa0Cf7uHbe2Fe8abMpa0bhVNYIoUAuqC1yxL6J9jrajoIIJQEgBwMSt9RdR3R
`protect END_PROTECTED
