`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8YHL8/TRVvizqA+Y1vuXoE0sZl1QBX6lypMjseEdeK1yS1aRDYi7K4sEkJjB5gtE
NGugIWotJK8pzstiZ/sezoztRaSZjbX/uuDn/qXe0dTwP5CPgTSRJpzKZgsX6TPO
l9iZLETtz22SFNhO0uwvjuqeU3FNPpN9FLxqEhsdUHz58Ah0FbjQ3Sme2q5CkoQm
HY72b4kdmlAxpKlZgUixo9m4rI8XD8QEFZAcxAZjDitqRMLBsoI7XUVIAIGBuktt
Pjvqf6aBWJX85dfIJIki8ogJF/b8IT9JTVCw0OmFUpcP/hMoi68PZj3Zo2rqxWU6
oFN0TMsZZSK3llS3dUcLv1wYgYnh4QFgT4bGGOk5i9egt2br77myiJ5mqDoVybpU
lgUxTUH3aiwN9C8+23R+08CLCFhTNuW7grQdipQCbyWVrOSeOra6qIV/4fwwL1JU
aT5xI1tV3j99ci5sYcUKNCWEUlImWzwwCje60TBjzHc=
`protect END_PROTECTED
