`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9Kt/9n4WRHV/FlXujZ6CrkAKUxErU7Ju9//JRYPK2Gb5TguDQZOrj32PlkFKt8a
j65aN/eQmHy/tS4GgAK4QmxEjty1qhcswsbnnkiXhlMJRp2WrKpCWQBDCqytxhyc
+72iUtydb+mo0+kocST9RHqPphZluAsa53i8gOwAwtje0yadyeNBUYpJwHsYzv6l
ATrBg42yogH0sE6pZAK0ZO25WkjDSYvfDW0kbxwMmKOmcj0+Q1D0nh4LxfeTl4ZB
QT1ok0HYyzWQONhe+I9iVQLvdaOQuma2HGrNAgpA+teQEdk2tM7yXhK1VslAY7Hn
F9dXwDuy7AjKLRPlG91pgfQZ0U5ABJjCd2U9jnGHpw+xArHMoQXU5F4SnyANjnVP
e8aHg1vg6j5QD5EdiwR6zCRbsd3FZsY/aw0gsfhNJE2xcoQiWfen/K//SA1Nglq/
TRyYSMgawUfrljJeTLw/LmenRFloO8QL9acXJlN0eQ1k29Q7c0sk3dvkpU+zYIgE
g4hqvHA/cL+jOXRx2qM2GRzG98FPJhj45AY+9w2jI7QiMKeKyEfCJibSlpYC0aI3
vuhYidVS1uBBeF3ZahvVNk1NFVhS3HCXEym5tlhQAx2w2K51e05IKXgfT59eNxYJ
WPkCVXqbQs6vwJkhAGh+qbCJjkyuHzAJV8daE9AzLPhtgldfTV1UJjjuWNcO98Z+
t/KIt+h0rdMoTSClp3vmeRO59wwwz+ry3tstaDEs/avZhJE1DN+v2EKnrhxIIPN4
vWsvyM7XEA/2o/y69z/E90edyhsUeJnO0Y6FojqeWSdvqVa04dbaVEdDMqmai4gO
6l5OVeO7cltBvH3kc+OM1Q/l5P8JkYLjSD29wMSPgwzTqp9BpHTYo51gXoLQP8cK
CAHUVyj/QwA87FkMZWvAiPYt1yorgwGQSCWuhDtc9EzziHZR+7bqMJdS8iJxLzCw
RmCzlJs6Z2nxvepW0g+lMbSs1AB171jVVl/OJMY+3kPjRpYDxq33GNVPvYmrfCX0
nQlfhJW1OUeeVWok59HCz/AV0+1nP2m7EamjeG6d9+VsVz1ptLaZjmv2KRgv5OaN
bA9yX6MZIVlZ/5leG2trN2/tiy3NW8UFOZVr51aaPFSjpWO5nho/LvyjCSx+2AOQ
OGh8cAWnO56brAl8qaF4s5pWaxNt4tkqkbBwY4pODVbjgLpcDFAb4D0Tigv+jYqc
jk6sCjLvYUnugwzMvnZyyJoMWIsPCWiF5uIhEElP/H9IhGSt6iwf7M+43OVRBcIJ
8OEoBPqPLoDiYO5aGDM8R12juvavAr47aR0Y0Mi/Tc7vkI+H0f9GBDm9ntC9QnCn
kg9gKw5MSieaEOA5sWR5/tFGmTvxgcSDfyCyvFSs7jbACz86IIMqTWA3W/8sJE96
FGORi1Ba3eokj1lkqKO31X6xhCfD13CTo/vbJ1nDT9M=
`protect END_PROTECTED
