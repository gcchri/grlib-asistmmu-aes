`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j8ikq5RBAzyVo/ljqKX06jl08phb3dQgN3dsecR43AYsCDAOhWw2jKueC/QbmyRQ
xNVFElccd6gylmTZRgM0U3gRou8S1O6iRR0L6xiuvuSB3xTKXJNvg999ZEjfFIMx
mTwSsWOQgbhA1/IGuZGTKjYHTHP17by7u21XINt6NLZ4Ljuq4uJq9oyTG0nyTVwK
L4WQa7l0BfsKQdX9BcFitfc9AJsFSlPET3GMXwmqXVzP1PAi8q5fHqTd9m6Wf9M0
iI/b/wtrCzghxQofkdlesFPtEWRtomUnXYPKiXRhbnVOdshOWgdmELpGIf3/pcA+
uqm9KoVP1ThqwvMhkWMkAlabnKvJ8Xg/02gHRrflI8vByczBy1VdmvAgbSyP8nLz
haM24Vo7i6up6Xl6ALtubpRFQFtd4byZmY77SFt0hqRl6cAnPlIVWSCA4HYbojUs
boyiC9jgtofYKEiw0SEhMI4xuOOzn4jEMKel651ZMzoP3iCtl1cfAwXeTC1QvrT3
6DzYGTcxHEE+2FZO5rYt0yRj/H5nRPcG2eqZYkD50qws3UmZF/UbwZilogIL4NQz
Xz0Q0f4uqcJGpaCrH12rr0zOPg7qtjkVVLW2FodiKsFbRINBLXF/YvqFgtojJKKC
6CmiAY1R7OPkU4DGUUi7XJmTNb6QJW6xjTPAOdii4q8xzD2qZAjE4yRU1nR0iqpZ
RbDwAVrtBQ1E7ZNstCPjn2J+Ya+MevA78QRoTS8Yy0u048GpzbTJiiEp8JiK3Ad3
amiWfYFhJ28RRfiqPosAXaCxG1NQpNj7zSgIXgiwEsgSDOtoHydGCYgEfk2WqziE
DtXOKA6ySHEsIJs5ERT3aUP48RdYhoy8BAUg6+561AgNTXD/WAOvinMR2+mreC8M
yXBmv1S58U+fr3KaOwpSDvrDcEy7Ss1kx9dveOP+frO1D69GrSo1Wm298ePps2UI
hhhGdmA6NTf0lLhRrEMzgJzXVv5kdKfdyvtLug1RMONx9v4WqcpmZAuk4xbnoITv
pFqis6fQqPX6EIIcTDEh3MTCEFPJHbXiBzem5+9QPVOGq39bxFN4SixiVA++YUEx
WLw1Qy3lJBeHk+LgsK3OLrajo438L7lym+3k+8cruWoumU/fdGTn//vCmAomI+HB
8WF5W1qESjwI3dews+PtvfID09vI9Tq69BA8LVh08cIJCU150lO1Bq+xxlB3dv6P
ctCRHLU0DoV34KebGdeaPlQqwFAvf4LnvggMEEr2mg7ZTBQCdFpMIOZIMDU1iWvW
RYom8bdPawg+vbizG9o80pVo/haDjeA9f4ct/IzEgOGNeJLUZS++jHH64uv9Evdr
/FlWre9iskR7WJaKgwYE+DhXx2gsCeNB9TWG+G87u1ZHFUm4JnO6jm+ttbwNNqNm
4/SHo5y4oCc8X9UbdnYeaBXy2kehkdPTqYFCxJEdT7hlubDBa/va/fCmsZnmMKu0
/S0mh94BKf0IVV45zh2d7Kn7OID8qbbLdviNSkDirTDZmB9veoUcUz3eYsyLdpTg
1AHlXNAAARjIiZBFQRVEap/W7HFkQAnMzt0yhnuB9TB/bpUbZF8tVCM3ZfsVP15O
YcddYMhrFJDBbo+kRj0GQ19vGqsBNvCrH4GNZawPPC4SFS4KuS8ojI4VJNfmwSrN
Xa0jflS4KpmGqfqZ471x8RiBTrty1dmORp0h0rv43seNXlDmhOt1/5nz348mvo57
GnkQnnVJGdsydWxry+Zcxd/yNpw5MCtNWXjiRQoWZwpqeTd3Ujjwg1vlAUlLOpl9
eg+qfIPDyXRgkcXxmQb9iim5y9wmsyNJNTojRJ8vJrsr68ZFU56RcFzyLYOHC+nd
VrLNFAYLg8N4PDX+OWP2E/fa0E6PsA+8R3gB22S6YoKVQ2Tha8ORqbpPkUBMhQIK
CFCaysi6sU61nLN7dpAudKLwYRMuVchby9cGkQmJCXtPvdb2Rvotxbm0q4Kj8HPo
RAileEuVfd1TDpzPvjdZT3OC60J2AQuMV5L6TgP6XX4/g92ViRUz8o8efovaSiUU
bLzIoFyuA602VAbDIkGcWyMWybnKjv8/rPjfXrtS46g=
`protect END_PROTECTED
