`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F1VA+PiqUsUUayiKTYoCcaLIKn8ZoXiUalnmGavgm0Ss7blbxBAmePuZz3S8rAgH
7QWXjTPY3FWO5wsql7SGnCaIQxUNvoggOU9r8K17qm+1yTNOP0W/M2CistbcE8EY
MCyiLPNpU9qfGsVCqOOuVE1Bqc8unt33fgZc8618S8TXshVYbpAb57hLJ+UXtTFB
VQ/7/G8/5b0iJzd+gGDNiS2BiKOpZJQ0BiFa9HY/5oo3Y7kNNlsbvzJfTR9c+mUv
Z07spFcRgNQlhk/Er+ElTn4ZWlSfyI/5gHSZHl2XzC6H7t8V41kdDaR9a+hfO5Il
DE8VMIAaVW9G8mEQbnTAKYdf6jxAVZt+j6hpLe1qBQWZz1wwHXwQd2Q29PEOoMN3
mP12QvciZMrjZ+pO8eDszPBQl8MtwVoq1QfJcXW1XPa/aNS/Miz7GemnefVC4OKB
r5gap/O5wbng71Kv08rEFZqi5tmCWSO9+YYj4usXeEIhwW7gZvrsrfErVKWnmEP3
kl+OB99RoETfGEBYOnRgcvG3D1N19zUsW7orK1TNPydivfZfPqoIRqhTzH+DoAXP
/gS8xlGEnC1RsGvqmkh793Wc1UJVkq7gBt1MMezQ440pdIsFQbmiwYqpCyhr7Gpw
I2e1yGiZQ64j61RvwwwPohOx1IUbJFAgVzVoqTUqxX3kLwumEc6nShtz/XCtc5Dw
ViSo4IQN21ZDUIZkJEpBYWlLAkZbLO4FD2p6LDi1/b3T6wFTVlEujrj3wzt0PUyg
0/+fbqsGPVkFcFg8MZeO5vTlMs99/C92UmKOaV/njqYV/SFAoNEp230N+ZtOvzGw
ttckO+bEl1qP08+VhJ8zcIY9POvSeGYM1vU23X5Rrrppph96RVvHdEVBX5Le4BEm
A2wR6QnZVJyMPjjfyGvtt0YOCHkLwXCtrKO9h38wYc7rpt6WCLFXJmay4OYb65rc
vVL23+oBq/l7zLJ7uwIa4TWK4tD0mn5Bd1aQ2te3dqs=
`protect END_PROTECTED
