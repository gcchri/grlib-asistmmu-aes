`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+JmM+sJM/g86ofB++ho2xYtjsrnGddj5y2vLyWqvDDQp25KTyIdYEyjCCi7i3Uo
33VWeSDiWvmEp90RdvGQxqtzDEsBZrGAU7WWbGF49lLSeMBQUT9WS0IDX5OsfKd+
s9s+x8EproQ5c+v9e/SPV4dH3OWliplIHGijuqkM3prdSMKF5phsrmzzGBPthZHj
n+3tXLeSHhlTZ79GRFf+fw96sL32/bQG83wBRyGcjycLHKt9bnpvLL9QBBZdlPtX
dyNCFGvUTWCh6QZujCINjB25Gi2XBaTlZOUtzKY4EiLkvWx4Jfpa1iMIOVECVk0v
Rzu3JDVLz8mvD8KzWHGMfxWCbq2hEJ5oyTyMYf48K9CwIME5VEIEpkc6FDKgoTYy
KzU3cxkET3WakXDV4eyeO3Fi04nlcSXCsmOf6SJsxAOwGKx2iBLoJp5q/IJtSH3R
NFSTsBujRzSRo/Z3u2wFVRPJccxxf1S6bUtsJdH9+FWNSJ52V1z8flZpgGuzwtMq
2c4FaVcIeFdXOlkxiHxboYGcuWV4HizgiqXmwtZONa5mS4kBkChoR2Rh8voTWGdP
efjClCXQpXkgOd2GG8wDlOEwx+vrPmu46R6bvH8aVRBTUXLt7T2O2JjJuPW9Ou8d
EvHJ6OOLvyJLVY0RhT/orY0p90CS9L4CRTpGyLs1bwlazKYfFtNbkoNJ8Lo5QbE6
AtRQhDzofu8IR9gGbQiEbrTrVs1c4hGvuI3Vvl2OI4dCjo7oc08tV6CLYUQND61f
6bHV7hc8ohYI+SFHY0vzqIBiC4aK/tImcC95baDZ9W0Ei2/knIQ4eKA6l+4jhrok
NrINXjfyAPXNaxKEsYGdfXgW/R8Rqe1bqa++KGXWvHiV/9DFb7oE7VjjP1+rppu0
2bf9GgVFwXTgWfPYWdBgfvDnEHA9Uw1PBOczRSkBP5lzhYvZozgw758fH4ll8d7f
x35bUqG8ld+2WsFbIZiK+i3zrWLH//Zb8ofYelM5DfGhPIzPi5xrMS46dOoQMJzp
SHDnLNQIAqf4OuFrPMaByB4lO73TmRywix+c/1yfkfr9Yw5by3XgnzV9dV8/Zaa4
DQG6HcCK5BQFlp6FdZUADgu1YyauvX24SDf9BUbEZYBJWf8TnVqOIJFNBd79eKU1
Ugl0qyHTaQmNAPyzp96lwO5hXibLsf6O6zSFTAKzagmxBoBfxI0ygSjsXhFbB19L
6ThoyyHDvx3arN04lYdbNhopSlC9cd3YT/2MuDTcQ7kBGz7BT6UW5tTWik0YSE/q
5o6HVx71mBhzDAQkp0HFOfsAXuxND1dydLg7BME+/anBMmpgHHfbjBbcLQNAy41k
d5gF2A954Lo+LoyeaVDPP+aDVIiGlWNyjWp8gyFIPBhk8221bKmmIJqzcU1+x0Ef
GEH7k5lrnkryg2W057ysR3o2e5GnIVN9kSLBjXQVJhWC54/8ohJdgUAyo1MShbmZ
57d9Up95PfI6IviO1uv+MScMbkomZspyByQiu+GMIppV7ipW9AmEMJtVZtfe/dUd
4HT6N8blQJMqTBM/gRaQChxUWEIg4uS0evqzrB37LDZrx3piZQOunlSwmk3HxTEy
JWlbPB34WotktD7MvATlpua5P1HSUd4bqs9gl7Rr9iJ4pHTIgghDpeMHlq1OgPHz
bfh2zY2HE3d+lKQCGbByJZ22UFFoQNLe9e4zTXoQOA4j4aDnse/DdpXGs4LH6Haq
BuDSeK/FrPDD5jEn/B9qDFVqFcI0iDM+LuIP3DecCtSf2rUe4u4KGqIvSF4NfA/h
QZnradtWtTLVaApmN7zmTSlN5PPUBupM5hkssYeLgvCDWUQBTHK7ejnoesLni4Cm
q1m1m7xMYaXNMcIpQOuCz3mwjps7B4uZY1XDLBTp9SLrKI0PhcGSjH20MnEbdhwz
cEGwOV6/XucmivC2mUdzSV0ULemMAoWk9PxQW2l+yICNI8U8KllVTrNr7XieHUWA
ltGPXmmlUxSfbQcf6/Ys/0GMXUr50Kr4PtJRH/c1VpLioyAUuGxuUHsWrFLfIe6i
8EV51KiXCyeeaAoANBkFJlyfHYyK5dE4jYfQs9fvMQd9E/Aj32kw6jOdiKtyD3TR
VJ7OYrNFzkpjxXDPw27Vi6kIRS6z3Tw9IncpstcCeXyIL6dp2kFzFyaUv62sKnha
BUTcq+J8JlkQDS0BJkax1kv/HPy+kib/buQaY4FgEk1x3qpwys8LbSwipeWp8dAS
KSyXmB5gaT9EOXaj1uQ2UMBFAYaBUAXzDPR4k8HrP5tUyDzO0x5ew7nfRBut8ulN
gs//0KoFg5aGqHM78wBgZ2SGCiS7j27qV2i8cw3xAI54gJDpLvUu1Z4YvpPkZog7
OGY/NVDNK4Qa1LG20K+7XHjZeHMfAJ+NNizY9gsxqyJ5qsUmVJtop6gowkDodP6K
4ohM8vFL4kGARfm/c7TMiAmz4IAi04dpScNVbrKDLkMfifx3/FgcuYjEgJ9PQhI0
pnLMsK27vMZRlxVasgAshW1w9NkZHSH9gsGgojwgJYoVndTLrNPvCH/FwNhE3gnl
lwB474S1xOKMQwfUKJMRlQy9kn4irA+fac0Bnz6mpE6xtP1Jlc1QSlwn3X1uKAYI
aJeb+o6aQZ9VXs8OKSp7EmAtMxTKvQdtAXD83wFzTFL5Xq644Nb2c0C6BTLtzhQe
Bs5Nm6W9PLUdZ47LIUlxpN8gxD3cB4UrE+KEH73i2Q/UNaKAf7/FkQGFhWDKNfeL
VFdq+Ue7mnG98ZHB/+NcRjU1I2rdcBQiQHYo8rdq1dpcHZJhvl4GgPr5tzP+LNZ1
unnmjGWpelJ3praPjmbLgaqtl/UnM6X3h72Vry2hctaCkPQ0zEcfNtVnl9GzBFWq
bKQS48UahQsWf+m778i+nxmwb95fClY54HPzg88qRXwZRLmNhQgCB+i53IRpjWIG
lXAUEg8loKrUM62xTvkSqWFMhoH8fhaLdp3IOrZmUg3yFUbZdna0g8llTyx0uDZa
PStnXfABE/muk79oneN3Ebw0vRlNhTZBBZex+l9Q+xb9z+r7EWrIuycKrxGApB2O
UiA39abgMbN/mEakZjCW5rm0mZRJvB4ZoRhuV0X54zryIgV/x62GdowvVi8EVEmR
bl38f5Eon6uxukvTjvTplXR4Ta7f1reVIFp9Zg8BWuBFs9PVonWLhDL4UzR4g1EA
mvzOnxiaWZayg7elwM5J5yNUBJuxRnM0+PZMTJirGkkNj+EpuH83cKVixpdsfWP/
i7aJQez9aeufsFZL6SE8r0gJ+5S7q2+ilg3CS/2Qaa1DrAnbZI4BqTKwnn9fGMZK
K9QEHrkecafn8AKQoJfcQxD9LxrWptvT9pJqy95oOsjyPUoDzos3I2MVB7iba/3B
tq9uZq2uEC8bkF9bFQp/a/widcQ1Yx/x7IlOBiAW1nwR/YwBpj7cqhw4D4Or+4tA
DHhbVd2WNuLyNGtz1Of/+Cwat3v+esPwGtg9Bl2yLtYIZoMr+f7sCl9adf5TJ4Q1
OnsAzfB3QNyjwQyJDyiBm9iUL8TizOvPqICtfWcpDWpHV+uV5G3GA3HgA+5ZZp5r
AiThof3LUzwD1ddFUatsPIhx94A8lqIfjIe/5B1Un/tuOn6oOc3X6CEkhubEuxPh
2mTpNBCKesmUGJXtuZoH1A7rPFEzwosEFKCANmCqhlp07gWS9t1cbSjog7xvBXWk
+8jilfg8Zf/X3FoxG59HLccl+15Zjzx+akT7ufeFsSP9oSwMSLk0+MnH9KH5Pty3
IWrymn/6R19pCAQuLmpu5cVESXjLS4U8E2sL8xidqvsUUKMCG9c6YFXwpl1qeTPK
ycKBYKEYvyiiJAafpcRyKBo+SabfgQgX7td2KIcrxHZ6J9qZxp+rLENGX7ylNmbc
FcRXi16Q7saDTtuSCFd4QU5KAWufu8lxDJv/DeJ+3nLBu3MI6HW3aysa8Oh+l3RX
PuaOWsEEqsikbThXa7v664wtlPmADAu0Spl720Zj0WEVLjFD22E51BRNnmlbpiZa
pTzny+LqV/8l11dwMYf9Mq7IcbToHDrb0F1IUH5htxd9lAtSuA5gKPTGuTUOwRBQ
LlTX4JFnlS90wQM/5G+SeD9GcSOZs11E9TixjXcDDcaxQB5p+IryaIvcbgeG9xL5
yKFPLYZGtGYUDUfV1ohNtczd9TovyLxdvcb8gtRSKiB5OZIGpxFX0lf2/nEkMU/X
Q6SMG7VlV7AVtVicLaMql54ayzZRTWVbe1pyylf3bPUfLocjbsC3b44/qBwvRG/l
cAghfhC3497OE2wAbhJIffV1ADoOxCIdOD6aZjY+L+lK/nqwZ76V6bmqM6HHGwQP
OyQ55QCe1bshnNXqOFlZKDUsDzcLXjOZKRNaZ0PReZH+d5uTxSw/gHFu9PwzmD5Q
vniZCSVDkTnkpuUeHIzKK35XwwCcMuUCrmwlanuMrIVj2qdr1omXzvdkntno2G5o
7LRI5KQZ5DFM9VuAsUXeWt2A7zScQUnxInPwcaVPYQfG6zMW7iN3AB4qcAnfNIxU
onKoQ/PTfV/5DEour7K6RbuFpb/9oNKViy09eDcVTQGTl60xYJQtmVzlXhAdp6UE
vULXFShPnbN0cS/V+sUhEVmbOUKQH22j9MY+VkpbfhPSbENR8oky2KtOhT/4KHP7
y7IJbMDYsmQEqnv3psAW06EIpCDmwu6BvU8LMRs7msgGPADE/KGlHAcPoOz9Z1J2
9PrTRka6qcMh5ek/Dl2V+fDNCxA2099x68CCsXkI3T+RC3NSI+vm1y7BcKr/BQmk
2qv4I0DBgWcmE0YGcxf+WPovb6rNdLF0pxz4R+B+NF+QSIfXpOq+kodMciR8D0NQ
/ZqIK9QW/lvE3UwAoqaKyN2VY0+nOX0auHkGmUnbQAR0gdYIuiblQQw0ZK3NbCqK
8eHtzNAuZM08E+FRsUNt/6kBV055KFJrdtqlwmLxVvmQjX75nyJXML2lBNUgBPnZ
G9WWXicwhhmboHWX3AcF3UxRWXMPMB8gxXCN+ytz2OBXtOb2r+uneF1NiMyHJNNN
PUgS6z3bUGVTvk0eYnWDl082OO6sD1kZkzbZz6b2amgZcd64nOiA8qkZz/YCRjXi
vClpO2pue0nK8AWlVO0WKlE/zNNBC57o79D7d/iJ+f8oVEhj7pYNYho3oK8+1hbA
hyfTmhOFiBnPEE39uuZ0SaeEwy1dBrsZoOHsrEQ4QIjYVHy+KoolB4Ht3RqVBl+M
dnZdERSjTEXxd4u2XI/R7+Mhe7u5IGA99mORzGvUen5WuiMdOA16Utm4XAwqf7fl
aowK5Cv+8yVvptUNKsq55nTsYAuRPR/ewevWSw9YlEpB1El8O7MQ3QigngISOE1M
ZmUsBQTxYWrGls7KqVvICsYOdt0tGP/Qmv3QSiBIx6/m+Q6c2bwCOQfD0Q16mOty
nZF1LjDQ4ErW3/WHHALdMcKPTbBRDwufx5p51tag/gGOuPy9joswllNAOu2xWEsq
yWuGiOSdJbQ6hAaV5XWXA6Heivv5M/AJByu1ocWnef8ajc+apBcpj1hNFi2DNhns
B4UFdsM00ukcPLiSxgrM8SLErU7S1PU5WNG6V9BMp6/coeMZwn6R6fiQN5eewdYq
90opYvZ4jWrsKMernaQmlByNdl7emYjdgEsF/HvaMLFE0VoBQhOoFiU154+t8uJw
CEXk8CbcZplj80V6avNl8sNArmSz4CcyUQIWM1currzDa6vh5gFKIOqtIkJDXsFo
99BE40+Ll9JUBXKkxaiQD/IdyHOJYBcGbpS+MydIXzyrexzD2miE9Ke2Zcoo/uZE
tW8Qa3Q4s7TPRryqVfN4YDeYG2v/UC1b/WYhf3fyZK9tuFYlSMGBIGWWuRUCBcrg
NFZx8R/JCw/SCBwM6IpC5v2Fb1rc4CKRfsmRgz06YcGs/KXTLuRUeAX6o55IjBqj
WpY4wm5woirfivcbxo7scn64r2Qjw2jcMURL/YMfcB5VRuUcxnCzQQUP1Czv5Q8+
cphyNDWgXnVp99GeRAbgwTjV4+hewOiErNIeWUjWcLKR52KW0mgZM6GBClGfpD5Y
6WlD6yUGqoYx14F+RyjpLX73sLCZSIp6aKJOQOpD62zyIIRqiMiyeOfpR+VxHnup
CAa+e/pNMCD3yTiJ/xSySFqW+NDgLEV/EzfevBC1F+syDgufQDE44BFxGzkoXRCM
fIthzZQezBSN0Ttb9zSlwcCMiCO87SJL0+aDbspR3wDlPAmnziWxkKJZZuH2VRTC
3ECfmagm6uk5W/gdcM69kB/fCzi6OAIOOUolvmWCMNg=
`protect END_PROTECTED
