`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDxcIKp2gY8AqVA86+iHRdKgJPhJNUCksqzcMtLv3WYxn6ub7QcHBxSSi6ECwBBD
95240+MBmZeZItD/pPOCgpk0YIPy8AKW8keOuwbCv76uTUYNFWX2JdfF9K+AA02S
nRATUecsbT8iBBcVItSOE6qTdzz2ASPiFwv6DhUHYON5KHffbjy0RG7WIE/D5qJS
PToc1YjfzJc/+DAYi9KoXcCmP2u1D74u2vKkx4CDBwn631NceOSjNKAkHw6mHixA
6rVkmJs+Nzf/ChgLg2+Kanta8NfYlc54TTLcBEkrA80pJS8Wbxn40qHX+E8y3Fde
SXkR2O/xiwjOHX+gBUtwla5jqZE0PUz6pQO6pIAwPbU=
`protect END_PROTECTED
