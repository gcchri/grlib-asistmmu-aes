`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MnqnNmFGgSL25WlOEh+1ZSktmcvQiupdqFPvHwTwx8K565P9hf03FdtH4U2rl14K
Rf1VcveBC25h2X9JfWY+LTVUUw+FWm+izpaAMH0MA2UwbnIsWtdI50Z1cMqu9F8N
PHKta4jAmdrVHBH9nSrZTPFhv7XHBVVWfzUNkFKB1nV+4N932TutC0T/fUE16J6G
26HHhkgSwcxV1Wbe4SfzEF/ImM020hCHW6QGiJhT4NCNaUt9ef4dPDDekB64aKc5
fVhyc62s1txVxcBeG66zUQ==
`protect END_PROTECTED
