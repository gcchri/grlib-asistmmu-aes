`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCMniB84Pzlbo61/5zx0bsfOz9x6MQVcR7E7n18QTF46w+T+/YKyxWdoI1bEYinF
uNfc2AelTsmFAsb03zuY0tnv9mABMEBKSpppK5n5XBkZAfxQ2N7NH1SQOn3dOgkx
hSjMTtdYBVYsOCNUsPY8BeRe6lLa1ogH3RafBqnSk3YpndAdPORC5IMTvLMFBN7q
P9cjGPxKMLkPXfGXs096DO3z0rU3odlUaNAeKJQ7J77+IdnDIO6gx7R1CujuEzE7
RsMoZrxYYLEcrdbwK8c0YLejus85Ija9Xc70A6/EElnAmr/jR4ettXr+epGnKKOU
X8zy5bveEDKZIYUXvpqZun6p58Q2tCIzXStW74YxFYm13VqarMxjMRWwf6QLew14
YMDbDOPukb6nme8lRs3SyvR/hSkjAhZpruWYOYbc6ZF84tMYtLLM/oOj+gFE4Kh9
7DIDJq53a+U1VPOaTZ4o85rgJKmfjVy5ypR0XjvYgh2GYwARx5UIkWtbr7AYOaUn
`protect END_PROTECTED
