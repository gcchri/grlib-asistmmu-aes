`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWZVwvNIyGgCcjOlo/e7rnicwNqFWPoEZsZcg9YSXgpsIJ62vle0HDocbdHB3dbM
if7rtLSbWDRyhv+CazVVfBYUSh3kg0tMaYjqVbkvHGgGbwFoHP4eQ9P27lTL4VYC
ZENvkQD7JfEKSn5/54zQqkXBnkTYWKIUUVgu3PMN0dDV2cIvHpW/SixV49Klo5ET
3Ljr5uV5sRucN99mPYpujjGl6gjtiuxJ2dLqwNLcfrnCUFYtwt2x3Hya94YFRVuQ
I3Kmp36liNQXiBTiuri4tw==
`protect END_PROTECTED
