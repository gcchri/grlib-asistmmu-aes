`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQ0KQbV9v7dcz7HAhGs9sMH2cvnx/uurlsgNAFLrdWTgTiV7VANhEeQbTT+3spXn
nxoqJdc8aH0h/kuGyahyZDHcM/gZcJyZxSyGT18KmB0T/DCNFBAOiC+ywoIgfae0
q3ktnnCVGjSeyqXvA3CunIaUO5j+u7r5LQwjLOFW2WKmmiMSR8DFqCaLdnLfCpHS
7lZHuti0RR79OWXTjBQDGLFOglUw3CTRZUPK+L/mtadjuNSXxUjXxctx+Jps8jVg
4Jcwg+cJ7OldQcLxXr7D4J91L2maG2vb0L7dlpOmOSnyIiPb1b2x/AUaXPRovndR
ghRYkms17ZWHMBr2Qz/PEhNbJI1HycUQ8B0jJGScl2+HjVCC+kjbefhuG8NSmYaN
gJTJ/8MFyi0+KnhT/CZo7HVJlDblWrPCkrH6ceN758ebUxIkRDIUyxHELgDN3qjW
4bFDh68LicLOhmjPj3XO5MrFV7ILsIfIbJwCDB8DNnpaQGKUzfiJNMMOk8shCpl4
eQMJN58CDjAnlCwLYFbsfNzpfCjP4NNLYhG44hWpaoGyURJPyp64BkICNofl3K1D
7Rb16RuxcGXDqPu9NF2WamNB87pt+oFDSlzBVj7Pb0GOso/pVOIHrwvz/OXr5LPi
yp+jsDZqabSRRoaxE0ikBJS/1B3uJSF+i/MZ7TjhdlUwf+B7JJxef/XcjfVMKxrQ
WKMkp7kZ5skiQMFcFtZKbysgpPGRwjNgPORWyyivukv1OWq/cH94+3Wg2GDdjY+H
/BTe7CCY9y8HEl0qztWUQEOq7Io3U6Pl3ROtPp7k0aEIyP7ipvHps1I9BCXs6/eY
ifKcLbN8GWg5cm5Xh0oJPrG6mkX9G/upvoFS0AFrmwBOYi1YsJJwigEN+/Z1CQvA
XiUcVMfBb873RqWKMV5VQ8V9v37b/UiH/DqA4H2l3ekY0SRFgQdml99oeNjhh0K9
Oma8Zb8S9mEzksh17AvTWQ==
`protect END_PROTECTED
