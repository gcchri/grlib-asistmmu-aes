`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ewexpVNVI966eYIi31sHN64qxoDzOo6z8xoVOAO7KQRKgs30KIyckQXyxblrVcgH
oBfgnfAlOPBGCdIVTJO2WvVh8qu4GIy+vyABf++1O5JGysgWOSgNDakyODCoQdzR
JZ+Wl+iR3dPtSc+kXKir2TIhcMVU5NrzL5GpunTMBR/4iauXpM7z5sNRcK55Yryx
YQ7aGCUgjYjrBU1UUIUIWmK0ed2qw1nKi6L//UCFUBWcW6en6w4Uq8DKAUdL5AAf
1nlFCpuAetLKqVCDaJRmOpzX9ywRgVXH+sbGupbIoRYwBy0rYhyYTxt+3yjyGLYi
o8hQbbTImK2QIQcHtri6Ulqk04noQZCi+eG4PzkR/QIRzU+ty73+HbaWjWImwCUu
5YFLgYao9mTZqHSggbQ2MzZPtw/bpBphMHsDv8WA2u9EsjVpy9KHHFvtrXKox13z
mxoUvBbUeiNnSaUCfh7dxbZZJWH70i58jymowN60O0ie86/ZDpqFaMGE+eIRX0BR
W7xGMMjdXQ7p0Kc6QAQUXemH/8nGJY6DoI9psNrKueHFyDb01g+EcydH+jUP05ec
1hGiCWdvZH3jPXyRmWpDTbCVNototcw6UZF+QtBBLPz1TU3+3IRF/pGWDCc+cETy
SrWgolyb3A2fvZu0WXuX9Q==
`protect END_PROTECTED
