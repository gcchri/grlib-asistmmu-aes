`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tebnPpvHRgj/cPpLeTqVeP4Dm/UGNGgWfRyeZrTy4F6QeDBBjsivc9qIyTSDaU1F
kl7K1XiGJGGSAl9Svl/AwND6ykr4NNfCQlCqQ59cVDGtlDoZPDipsjgIve4LjiHO
7271Dib8+ynzQuONbgD1z5ol1by3ApQODlhpwKltsgogeMj3wEcKO7ceGaKoyEGc
5KcYzTOEGnis5n5GLYh2YkqH1z6MDgmPMxQBQUFYytnVGTlZbCZ1OirQ9/RcXdUS
SI2PYepsjvfflkzl3eZD9fTDd9Trd7BP+FjJLZuSs5Unn9x3q22/8AVvQx90+oIj
YbdcQc8xsU8aq3tW8YNVPfZxnZ759mjmpi7Qv0QN58d+AnlAcLgd/B9mSggF7xMP
rVn/s6duy6/p+q7JakJ535KbU/JxAwOelWAB7GLW7VXH1mKq2mvywA53AuNaB+nD
+7ImlNDODGL17G956NhrBXXCv886kr/z/Mt4gfW4c+oLGzcLyrJrs/q2wV2nimf8
INNx52+rkot1wzVAEF4hyyF2Y/3vQbEE/gMx4kS4eH3L8j55WwXJx4PUAc6fF+BQ
8rr9gFbq3byaYYbvxKCgUBpSGP8jZApgoRRm7lpRqcHkvXpBS2E/m3sjR4w/clSo
aa3ubcX7P/9csaKg51QGVUVEErZSe6hB7ZBw74HgElwbcujLTbKtO2s9ygjeOU7Q
oE3WQbG3qnHq1jXl0XcYNfZBZxSbDn/8Ai+2GJ1P/NSLJ+NdHkye3HYoIqAY8Pkw
6dhY8jglV8Cz2rXZUmLcFA==
`protect END_PROTECTED
