`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pgx3XyrhnXiLLlBIdIOE/Pi6pR4Rz441wZD9W6KixqLWbzd8qbZgepo+ADkLEBN
qzHoBB9ovgRzDVDYg2wWiUjvzuLAVL13lNNWkIOSFgqP4DianTy7fDUEPlOi22VX
W0/aKN55orkgqhZf9F00jBSDj9tAW8Y4Gi604CGzxGxBwkj/jWNlou5ohnQKXHV+
K0+I6pjQnEhbnTa/IDV5vTPP5L2SeFECJw38d2wfmqDkzgP/Mta0/3cC7K4eW096
KA5cz1K0nHido9fhMR/ntqUjfZ5nTtjXxxN7qLM23ozIB30k5kA4GAVxecxX1tPv
aHjXgUwowAqQmJNxaXZAZA==
`protect END_PROTECTED
