`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XYVTEIxK8GXQgSPPDxABvXZzSyVBiZqCiSflczZnvKk6UGq2upAmmiSnA7TAUZp4
Ghv3eGvqMpHR9BeP3Y7k46rJnEKxYYI4cnbAqKza1zEtGrzwN+c1lERl9WPC3qqq
6nu5DaW1r/CN7I4t3McBtnIvjeW51Km4Vei/vpgwNs5EOkyYjX+kjROK6BQYe7RN
EuKkuY2rgRF11QcGMjFD4fEYnokLf+AC3N6tpQtRXmEeLz1iUK2H6T0IN7KlFQZh
fmb2YoqQCO/Cvps5DdZpBLhqlJGxpa3Hm9RAkZLcaVYFjLcujIV0kBaae3k1To8z
51dSkeXB+ELPETYc4amRBfEGGNX/nftbQGM/8KzcUVbx87vFMNRMhmSoahyJ1qoU
4RqY5FapXvRK+kjYbku6JidmgUchhOXDOYXps3M3J6QCRruW78DrPn2x36QzMdPs
+6P44dfVHjL7MpkGa1A8rOzgkKzdUCv6CQOjEKCWIk95Oyc4ouTLwrRpBx6kvFfZ
5DI5vfJQsNeOXmVWzByyR+/h/i2N9ciKkm2YVFor+vfoh/wQJKO/fD0Ni16uM1jt
tzelwUlxhO/ZiUwpOVGtG8ToHmFikChvEzQihKkh5zK8WCWVS45Rh5y7B5XJJRtE
Vwo8TDfFs7mfwLiIPziDCJrLTfZXtlGDgzklQvZIJRJL2drw8wvGgIr8zodRs/2T
`protect END_PROTECTED
