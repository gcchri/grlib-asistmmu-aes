`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+fLd03f1a5mUDStltoGe9IhXhDNlM+VslIvDGj5BhQLgkmmLj3fnGZN51kG4uyH
RgbPPShj339ozay3h+1RzW2xwwFCIZ1J9AYXbzxlF6apNgsfgiSFpXRO0ESdOqRr
xAGbA8p3L8G8JPkHfyFjqytNcmI62PwneSN+TLGAIPpJJu4XvmZN52uZW7ctJmJd
0/bBL37GMEbii8SV8geDXGunI9u1sVfZhh0uD+TOBZjbGW+fU1snmOPoex6jaMa1
2ZmhHkL3EN2kxSnxsb2IO4GNBYJ1RyCogt/qMfFTteTjVlFb6vnV1+aZDONzrhf/
ckTLhnC62bM3xJZ3hoLs9ViERguSWuZ/e0+3UM96vRY=
`protect END_PROTECTED
