`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5yG26yZsj4UWwqxm8KCFfsN+lk3GrkEqcOz2m+MTR7fUPvZpbvcTYLUUaoVh0cmN
fsEDLNS0AEN9KYqzXXE70Fe4a4YXJYC3rqsniTy1rBjga+agqVxHrAKouUYUAR4p
NvxwPxmAuUtHUBAUNvTRg0KwhlZMxwj9+dYQBXUiLwF10l+EVbHw6FaeDVR7Hs4O
nYObb9Mpc6R+uMJbs5wyMywE8iCCA2P0T5geRpLXQ3FTXc5oJ4cHbgBk4XfOdTDF
Qlx6H7u3hQzA2yxEKjps2qOqbbMsfUqRFNWAsxCm7ON7qfSk7RlVRE2nRrOHiJxY
sTA1E3lQiV8Tkwtwh+jIPUMVE4LfllOvV7z0x5GsztWNEijpzTtRXZC9I8pKZ3YN
ubVKSCuh7CYYJ3+djYYhJzCTVm7j+2gs9ir39u95VWImfAT0lCfIbE7w5P2XPHKg
vXx+36H/rTRfhEWm+XBpTLbFKB9gHRDx1sCGz635q4M917Sqng59tNZiU7DzSxQC
L+MPx5VVM2D5nDsjQTgIrC15vmWOyntPNbuiraoCDQXkNO8WRGfLXbYepvToG5AJ
3aDllaIMSrI6hANzP0SHEad/JcxNFU+r2RsRBgaXZk0Q6rZOVxzfcw66XooSbL8x
uZjLcy9Wk4j0WtEb6TgBQcc9FdgT9Xzc9I0DKaYmMh39G0CyFPqMklP5gOYkBImg
+OBeNgqJLpbxvWltNLdHbs3YgaQ2qebEPWcy024eTotJmvKx+1knOSUOAXCXI1cD
j+/X5ShLMZXJcNuaonlhbkqDrQrEX8y3hzRCQaI3nKBf+RdLcBgZ4VafDRlAy6X/
QcZHEZnmzCbuTB2YAIh7vkflWvHbusfGFYTkMQdAHk2CTCoKGBZgBTWXkag2iruF
N7ll6JFExJl9Vq+X5P2uc1blc7oQKVHaX59nBnqrCwWRZ/Dk+anovGnUEVi59Zt3
`protect END_PROTECTED
