`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCxwTLGaoFZxmkVkpH/XQt1Z/wrW6EUBmNxLWDkm2wYaqYun1ZjV6/4EWZnzll8L
shxdFABRU7fbh3DGjrXOza05qFBSk9sBjFFD9QMqAQMoGxpXck4iSnZPNM4dnAyc
W8fJfCnBiFZsrg7ikgTMG2RbL2R3ck4kA+UICpPJWizmYbf4tGccL3wKk2pML7U4
oBBhDVbWrANVM38tztkQhcm/NMosfeONr738z6XVQwaIKKYVQc5kAgfW6RHJLNlV
k2pLdpi3ecsTQMw0/048ruUWLGvJysHN52kdrNfx+weD1cwVTpHX2kcnCqNKRZpR
cGACJemJJqEp7PyryDPmztN2xYixIDUi6dBWyqxOTunmfwJRnDyONfE5AlZKHAqa
jz70ysrsp01O1jymw4j71xZBCFzuuu+6llbWNNzE8iLxcPzx3FdRIff9H+vha1WY
FogDKddrEv36v4+vUAD1yFGOIKFdmqCbwduoVzq0veR/9bs+NAhK0QCSN7mc64OW
rmD+CB3OUGdVy3M2Xd7yzljIxCDBew0wUead9QHX1/bocJbI5SpOSqQ3yNEXBnym
DxleAjwHhwVd/RRfPzKtP4Wkn3I8ca5iXTUcTcPjDJf7wV4HsXGetP28HtFWhzPL
OdIBzCGiFrOJXuTPR7Yb7N/oxskjkpARDIa9gR4hI/CAHw1Q6AqvH79lKfnwOwZE
4//BjDwhOj1nvwUtOrDhaQ8Pl+Wg8fAAr+NpHccGF4w9zAN00apj43EdpUWMPh/x
F9oXJi0TmFIQqe27oLA14xyzM//gOLvK8AP0tZAQ37liHZlZRl5MLJzwJKUuOrQN
3grp5/Kj7JGlqaJWFHvsmeDEBGo+okhS7n1cdygC6xDCNduVmIgj8wS9ule9zS+g
v/DeFUDPmlD2xSmKKnPfKQ==
`protect END_PROTECTED
