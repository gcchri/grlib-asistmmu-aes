`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
im46nRmh/4+UV6B0imUX7G+hN2HbeNLKJBPUaisFqAF+CxssSjJotYE5YvK7jRNz
h6WI9aJqkVmJV7JX5fKS4vJqGLROHBq7faRzzeiDickIQUU1vZilvYJYfkJPiMgR
BdJO2BGiEXr+JqOEB8Sc89C/EwXtQX6gXvFXptkQRftttFK7Zc1gffjmRm1fTJNS
jamd/CBOcuFWbq5YIG9u8NYtq8X/J1PfZ70POBtbksAtVrQFAYj9W11ZjKING/N9
wv3BKziJ6c+g5+6Uk2L/wxErJdDHNlF5f8TBnsuJXdFu79+ApSHiPGawSH7WUZMd
pO+Jrm9rUAsyuSBsBrCTS7BHx/7HMIbPCvZrgnSAPdW//0VlBrlI1F2IEB+GsQtA
fOOPUmPkCdtgDsVGohXhOuO0J1J2C+QP4+/YbB5+cx2Zh58OjIm9GoVBzrT+Xjmr
liVTEvmBYZJt2m3uzDC0ihBT4zmi4aFg5GHFO9TqnjtAaeWV2v6+1pj1nhkBeKgU
nUZ9aServc9z5xPs6EQVariFXfoXhNNHEkTtkbUy2YbQCM41D8/Hh0qrEihv1AxJ
61PNDKpttHeYBqPDAUClToH4Cy1n7eaMcytiErwBObo=
`protect END_PROTECTED
