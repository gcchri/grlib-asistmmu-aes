`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kv1Pjnp8WLZqhCD0Ivhy+Js5Hptzf8a+fuiF4b3GlpW3OoRVfAFWtxRieCkWWhYI
C1vbetqljHu/zSrP2Dm83y2XVXgBpW7dv9wiG00lN0oU+BAbCt70MpuwRYB83XRk
sn5vI3veHJaplz5lkAbpckRFa8i1tuv+qJNzFAai8Sxvx+T56k9JZUxFTSnTn1FW
n7zKkY/FAW3RHqJkGDMj62SCAp8wAmoRrgRmyKKxopM/Sch6nqxn0sNnUQE8nMN4
NCs6WzqTFzr9BGqLY3vR324RIN6bi7jDZ7cacH42KhTNi8l2VhtJNdrLtTqsmCBY
t8Gu94AtFZTCZHpIeFHoipTbUd3WXBEQErbUdShUaryJDOt/qqyXvnINXGKeT3oZ
BirJbTOIDKShokfanNu0SA==
`protect END_PROTECTED
