`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1B6Px5x4r5T7w0sxccMaEJiqfCIPYQoYxiB2YpLl8+/tY2gcE+xsq/57nSJkPv0+
OcUtG1NdYR94KopUQMRQXpb4tjJpYKaOmYSCIDusKMSkpTbSiVktfq06QkHIV8AY
ILvG9tAYnJ4RHv1xpWgmjrWc1HYzTK5aaaICVicnlFKusH3BwKTDLQ8wJg0Tgwbi
rm5kfLQO8vRrU/ICIKjzckhFrnaZ/sqMk0Z0OANR85AISYq4tbWW/J4kEr5V8buK
pPK5yc7qZ1TMHtURMX99Gt5FBpVoy0tMZ9pXHYF5fJdYjfG4mPPa0sMMT15m/C63
c2EUGD75jO2yiXjangYmGC39fL2sgdhUa9jaziMWKkXLS1zvANKX86Or3BMDUxi3
14flLTkgmBuSnNIR82+DIBUxmRwrm9Gu39iMgGvQQCje16JscgW1LQgYSmyLxz9+
7LfbWrnNnaWk4zE76Y/SXpJnbu8t/5mUpyaE5F6KtnLtg2pzqV48UIB5W62tO9h9
2kP953Z/IP8PL1Ack9qy7Y+LgZabxnZhEGEjMULvstM7ivupsHUsUqYhXAhV3IEE
hMkKs7qYjRB36bOLamuKd3NxQC+Ngw4MbpsiG/b6sxxESb075RDlzux+WTSuG2gp
XdqrJ+gAVXZCLrH+VPenx1Sth2C7GCPYhpBDZzEFveW494U1AibK0Bj7fbyre1dY
NbdwfCFBhjsuuAHUe+AFtjTg6L2U7HeLIPupElY3vJmQUu9Ge8cN/3jQ019suRub
hzLUGFoGVBJZrio83qkmit1wM4GHVCG/8n3k0U7mW69y5hMNip/8VVu13x+wG3Uw
AaMEvh5XLw653VW5kLSCLxPhaIQJmha+GD0lbr1zofGfoHEUjZ4bFgISo7LrPB6c
2NYloR+pzY6wlIr0a6fPTnfXtJshTqg8Fjj0wHB4GDEghFMXb6UxDYZViqlVo7Ws
Tq2eXRhxCrlJTuXZd+Y2PqZ6ZadbURvHdh+i9++vyeEltGoyqiZuRBuJM9M1FI0l
lRS/9kf3LIG03BhJsM/9qZG08exrx1PWt11RQLv6NjarlcfD96gBwxIw3FAe0RgJ
acCmzXsUNgT2Dy3m3xw8z9bSJuczedLVzgFUcA0zq7WHnqzD3r3MEGRGnIAr+R4b
`protect END_PROTECTED
