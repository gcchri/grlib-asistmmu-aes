`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4JntHnWfcAGH3b9ZRN34qLUTVqWYf70B79tUCU7U1P4a0TrrS3MdIrqoZQ39rvlw
nyUguImux1k7oTcwhr+3rpYHc2/8O3wKRoYB/lOPH5ugF234xmNzbcWCR52mgKqE
s5bgM/1r7lxGRbonLAbFOVUcblXJiIIqVr91YTBgJ4tkan4I61oW42mfspuUQGwA
rVWVm2YeACCdwnfSZerdf5YSI3SaIHurGHfgM4xQp/TolfZRtHpfSAO6URfc7C9H
kuR4qBCzFxa65gtoktH+GqUuqCAPOFNN1T4iuLOxM+B20BlHKcaCtyoySRpH/eZT
5OWgdY1m8vIagZppL0ZI/w4Tiedtt2DNKCqmCRKGNdOFruGj4i56+N+YAANBrYp3
nERRE9AqI8lhpAcuuNx2WfWSKJTXtsMRLa3LKRNF7ONAPiaX0HDy92dNDO2OhqLs
ijYN3V8sDuF3JhuRpl9y/znDNBnfAAl9z/yL+5l8fsjM6F+pRFuYt0FK7RyRuDw9
9xUop+tux6zVKwSVPRau5jniPRx7jhpufyazyuqZzw8k8oC7G0S20hH++d4fj6Fx
I2yLwMxIFn0vnE9LgtNtjdpC55ElAU3R6JN3P5alBRtqm3fyeBDVhClthxDd+pWv
gcBPmk1K19YZOBOeu2LOQN8bK6hRj2CBGxLe4bgs8GP4EqtrIsPsBALnRL+UTWFS
804rsV+lVF/51irTrz6rHg==
`protect END_PROTECTED
