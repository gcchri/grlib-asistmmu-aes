`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6s4KI60dNoX9yK/ELAAxRUFEZaLTrd3I5TDStxrCPmrrqygo/2zMy7tDGVQZhnk
3TKZEhAcSFjhNowZtS/KvitZwIGLK8sbXpmrV3ZV+3FeGwYPzlHmnztrEdrzdsqf
GxCS0M6QhfdQtkOgThl74gxclUzckuktrjp6K0hMBi1YUXDz0DNo+qKBHnu7Uyw+
8gxnOnVTxT+roXt8dde3ykFOjI7UcTUx7dxcGhykk1jsCL8dH2vM7Y2rlkk4K+vI
PZFah4M+Y4W8pWIcAEsZ6WsuBWMMXQvcXpT53cVTmaEtD2xkXHw9XhJFijV4Vguk
6bSAa0fzyyJrkthKw075qxVV/gG/mJeL8ngD6naoVd0xIMRZBZP7Y/+PG0xlBgpE
vKny2QE6GF0EG9vR2WrY9XkYE1+sCWOASc6rvlHgoYXaBLsVABSmdEuXjFvUlf8/
PM6o8Kkj1wyY5DBv4q9TPUH8v183x90IsCIoiIPcjWpF557X66SZwl7cJbV07Oc9
p8xuzatxpp1P+WS6ecHQNQnnYYiTfeRXxwrAmFGU8siOjqEbKaFty2Vr1zB2XUxH
sxcfSM86eAnZwNPTbzglK5zmwwOrTuPICX41Nk3nJGbwdAhXdpEGBlWcEpJ4PBLa
PhAFDhKbWM9/94gmWuaQnYCQlzzf2dL6TM8rWaIF9m/icLfvpQGfw6yhTe1HUpn9
Ivbvhrhr9bey4srwz2fyD7nOM/92An4dQQzDewfph1MFOFW4Yo/sSas4hB5554Uv
HKZ/OOHTDb57j9vhCK/ISfiN0JlKb0QSl1BBNk+fKPsEtKIr8ru9M5waxowjmPPK
JRihtqzZefRZbhj11OMQO9ET9IjkEupoDWvxa6R6R0RvxXi2nLAy0bgiqjNcK9By
DgAZovd9xB5x5oEVJZJt4jVhFOcAKOBQkleitYY8UGppzqtz55lFO0mhbx7fp5VR
baLT5TAFwFuz3Fo+rdto/jKKw+Vjy+dW2wSLxtYZWyVg7GC9+cbyzGN/fWKwuIKv
b3MqJr0nZpXb7Ian78h+ToMdS1UD57yaeRGf6NecVk9qR6SJK6AgDOT4I44WGYja
hpCJuuQUqES5NxOn86diylT2eXuwsKy+6hUp7eHkoSQQ4ECUCAtmyw2wpJ4rXCxt
PHtjJdNJgs9cbpm8cAJp330uP4iyKHbt+5eGptFUNFf/SmL42wj+qbj368ViqG7r
W4grPk86n5mpv8tEZFHW/AdugT5d8XnVVPSCWedePerFDWaYrftIrtNH3laq2GxJ
sxLzhI7ay7+W6YZA6bJPLz7tGcSPBrTAusFL6yhzuWxnlLrVgsShwFNVJ5ZTDzCx
fweRDGlbBecdGbjXtt2HrupOUJWm1j+nOfFw2u75nYMQuIYpmn2M9WjHyQdX8ri0
K74GrZGi7OZQgyRI3W50PQqisNraX2DNpFZ64cqLV9hYNtibjbKIvtgk5GiKvqaz
pgdl3fEsqDr/nHKyCU47Q4qGVXi9Cc60JvmwgUQOeiLYBI1zRQKrXoVoBAURDrVi
zz/cwLtCcOONQN/Dw6pMWhfVT5Pmxuk0CYc8W3d1orvSSsW7LmV2nAC2/Vi/hEgG
baciwXzO0b0IrFQZK/BSl/LXVZRe3OAtJ7BryYJMZAWkJvT8+4eP4vDZdDJ+akAs
tIxaao+50SPfep70vtzjZn+wlxS9x7AOJKyhZIn9GDdD0L4Ue4Lsv/bBoCSG9hi2
YiiCdEoNWgbWMCa9cbgCtWk6Ckc3oT18x6QCyICfTQ8GS3+dvVi6LL1NKzmA726Q
1iad8FA7E3hx0BTStyBoAgFnQE8fSmmgxN9Djp6OiJb0Bjomj2z7bvyq4W74CQfT
EZtQxRmbr4n1FPYpd29Tph5yZSf8B/0wJb8IZAnA1vmykqZJ7M3RzyyuOGCehalu
u6563mPRJ59Uz+Te+5WsHplJ/mjk4jLcGssDpMQc+p5Chg/NOqNvhERWsdPts3JC
MEG6Qb/lzKpeND77EGsEpqe0m3bGMhSIOQ1XudHmRqNAcqAnP74GEd0CKAaqT1/Z
ajUGNQmIhNpi7HA3yXaxOOLsKehZJjMUGleWKreBk4OAAF4S5eQ4dOhLRAdh6VAY
tOkILbaSNWXefJcQeQio4JNMdD2wtufsus5MlXEP0P3Duv4AVkjhNHOMokNi68XN
RTXjqgYfWpsmPMZkgxlptY2CtEqtfDSyLvt7Zs5V4Yx0ERWa/rOQt6UC5YN0ZUGD
Unbh5gxt+EPhrFSgs21cRweyqYuUVeNgdUXErfrbnjLoCyOTc8K4jw1BSnQWTFg+
HCY8h7VkqqGBTSQOtQ6uhPsqed8Lbppdb6p/I7pdQ5j0yYb2WWqE1R7Poz0/NYsu
s5+SAVjj7886T8lTUDwLC/fOzJRL9eid2sNTMrBouc+5KFOaAkYTfVy6eZFaVIVu
Z3kG5k8Z/eMubs/NKWmy5xrCkDO5Jr3qLoppGAU41gxURFMROPxSfB3sS09+bTYM
BcedXFVD6wA6buvrlJ7sDGEVVp4ifd7O/lWosBSbYzMXoWYTGr3tvOX9OueXSnSM
qawwYdLjOvwlSugQCfTV7HrS4UAjxmQsbjIHsNZTPhWh66ddWjghXsXoeh8rxE4S
C8WX9dDC7WRiy8uWcTqYr4Wctnxkhu5yFH9efHEIHBlsxTMgPgcd3yEqt0vEDYh4
RzYKJzFvDREPqkbGDQVE9hDiygrv26vc0rbKTHisnHci6dNzw54/k9H5CpnvVuD5
Bn7NdLuyYwIYD77JZKGeakQPfMFfCH2bOq30fK/LOIx0teQDI9l7HqvdaLfHFE2E
NnXClfviIoqjntG2dp/8Tw2aMs9UnhFohVHzoFy2vv/jP9M6BPOei8/9JnOwKebA
rNlsS6R1gS1etos0z9SKI5eusIbJTOlU5X0BEmP+luAtvlP4FnbRNlfiT6vQA5YG
h8wfMNQWjDbTjOIUqV735ONtyDNcWhc4Dy85RVQCp0FEVvnvfq3B6iUZi8M96sfu
B4IY+Dd7pysUDoud4nnF7YD/vw6p5O4uNq0x/ZRVSqrLDufrkWqU81+z+JBqQeZD
4MMUC3Q+fsq9B39knVJaWNll3xT96q8esuygjupZ0QYpQt0KZin+FHLmr8wMNX85
e44kMK5d50tJUgk8Gc3nxO2YABbdQv7Wb86ckeuB8GU/EeLoPmWPn2NJuxTqo/es
Sm9P4Qjd1G9KebcFj8h28SgoA81HC6d5u6tx2BXNQbL8aqro4b769pLxfVC0eibg
gntONkWVI+aWLk85ZnQorS3aZI20tMpbKP2pggwWXdZu/jBmKvOqKmUv97ikhZlU
jBPG8tX7Wq944ehAT+8lX851UuTPHZ4IFPZZ5x6yU/waQbl3f+9wBPoBDKTqdNHj
vcoYh9kjAidIg2k0nVgBtjt+xCB0O/EW/a7c2nc9e/98Ee+QbA/JwCdoxq7PBOnQ
pq6lIbZ6tBSFCvntUDeVRb9vcMZzasJX8NwXJeYEu3MAevDKNnGmGm32h6N+71GM
xIhSSz+OTnkH9AdmjCpORkeB9d71afscDFOZDbnWGoS7zZkjXVKlk/THseRjLauZ
hNobSUuUd75uuK4aK/P+Fx/E4I37+qwH9Vl7eZuHxsJGSWmLZBFlcTwZ/PoN+J2u
KFybFeLA67wa/9ZD+Ib9j5A0xYGm8EYyxmpvu3p/l5qXPWfrBGiDiYllcCkM5So7
YebcEl3/xaisMhfA5gCLiHFyfbUEHYPJq8YUzevYwUx6wDKKsVLXeC1VBYHqv7W0
XY8578HGDrorMgYN9qjkFMOVH/oXUlnznJtnI4uGzC/7Xpus69mAZTjJh5YEm1+5
ycS8gfH/2hpWYhBHBv6z0K30AcK+Ad7UxCSlO/IOlOLufDn2z4E7DsjWhjanulSh
8+TaoGE/RsR/3iTy/8IVIZNi2d7wYaDrIRDa/FPwIMw9LoZgMC2Z+2+1+HDf/4s+
PJR34d9MZgd/5i796JoV2mR5NeS0pu9wtA+8kYCJhrrrUyNScWuHSXl1MTNGPtxV
n/pDJCPXHAx7/MGWKKYuCWLJSq5GKJnu8eS80oBqg4URq3A5+xhExI3o8aUZSdwm
UyOcbsmpxKoVNRfEeivQG0WMzRNoeIsFr5AYyvqZGx3O0n51Cma9gP+w/BOmjIkI
tRgGBMv14DnpAk9oLuxVPpvya1eMfYS64GYjmgMx8iv2r45ucQH7UJpstKEQzWkL
ZE4FkETnL6CsdzJLorVa04lw0S5T74X2R6WWLnVkc81pQNHdbcSC5dAMJkLuX0+n
IciS+MaHjsT61g8vG2XfyYKL3MdQhAAAMUHSB5c39Ck6sH7MPJ8tqIVBqITJn2K9
gLnLtyy035+53n92Y3YgLlUGKksORfz7HpI2o+jW462OoX1b8Z0i0wVLzXyJVqN2
45UBau1bu9nnLkPFxe130KgDdV+1uJNdbqtze90b4C/M4eT8hC9+lSsz3GlsY/jj
IroVWTWVDvrhq+VLv9Pcc4jKapvZeDOQTPEu6wasqzIfEBH1TEiNGs81awR3caWF
kVW0THHjD6Mvosa3//7tKgQjJFh6xU5R8MSFGmptEErOttad2+byD1v+p4xhc6K6
uFKpjDxLEYxdRsqPOHFtxfhOuw8/GlMipymV27erDeYenRFVgYHhxUi2SigKEuKF
uIxirhZcXb0kyV6Zwb5BgwCiaW1RJOozfGpbJX7xEzo7DnAfKYECDySAEa0zQyzY
QH4PX0VztZReX1G4VpmDOsx/US9LdL0Eg7rv96M6KT9EHTuqHhkJe2+hUPeWk84l
M85XqJjfM+kOURVmM8Q4BYTeWjV74x7/61Y5ll2GHoODfggBMsDF1r0BVjI8+i7O
sIXUAqZPZqIcGeHZkXPoF8HdWhaceP3QQ5yLTssMVKADKZu9I1LhPok5nEX455Ua
wK/zMiWcvshvcA/DqUpe/4nufXIg6l/UYyMx0TKnz7LkDEIndeT7XGTHwek3zGvr
2ldp9jkU+JhXkKEpzaF63vqZGVoIIhV5ped4CHWfosMPXyMFD6dGh80zMRmnLIbY
qqdlehtUNPgNctc/uKuIg93w4m1HCZn0n0929/hSsTZuhhJyEZ/bAJPG1ca+GLdf
HzHKc+IyDP3exfShjv+Qz1qJwUmh4wJAMTxESSHyhMbJgkBcfGgpIUSM3UgRCBqI
zTCKwK0kKZ2EeGvNShTrvivsEdKDGYTXle05QbjGiBTYQJcNcnlS/Ix4Adehqbco
SY6O9zDGqDuKuwuavLGtOhxl32giESQLe16yPDySQvM=
`protect END_PROTECTED
