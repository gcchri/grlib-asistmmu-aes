`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zkeilFc33yfjFU76OP7+b5H8A7R2c2tZDuMcd3eZMaunfXGNlghC4ILk2PL45IYN
Bu8bIdZFjUfM8doKyPkZgXI7y2HNjR3W8+xiDscW4vfSot87gOzypRcUECPwgjVk
IR7CpwRv93GCUQqy3zoCtjgIZ2kmPqqPXrHJUR7V1QbWDlNFvmeJWbkm16i4Zyf0
zk76JNjPNHlCOIl0Dz8ESTQ+oLfGJEYykfEVjNui5xUs4V7vyGAuwKyUUGZMIl68
ISrSE9lcUfJ0icYE+HQnCek+dMLtTaiULVHUHAuYXfRRXJBlnCVdlNPc17RShgqz
0CGxrwX3Wc60tWbcIqkJXjzZwK+HTXcEpNgW25XoqE3i7d61colhxmp5HRpyaxOL
BvDOR9b+YmoFJkvOXqjB6XTwdS0BC5JkykppQc29pNbb9/OQUQB3EkwtOntocyGA
`protect END_PROTECTED
