`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ePt7tX0gfiNV7qxFZPx82NS7e5AxJ3GmPoJtIdWP0jU1a6F73DLhmQC7jNTI5rL
X7J6RlwePcgFhnmprcIc1MARNfWmmHZlIa1BV9MblCDZR/6t98RBN/cbKjcYSfG/
GfhxwDE5zhIkPHwF1kQ3h14rH2M0sBhsLpQmd4Li0P71ejKY5e3RkV/GH0UV88CD
vIN4b7KnjwReiSV8s3byASIrjT9BWgFH9QvUIQugKyryFLbEt1fHZd5fNvAcXG7K
UcNvUikEperAEjYc9eP5e8f6vn0Gbhi9mxVnubV42rjnv0bspXJMCwykmtdW6+O6
VPhnmGI30Tn9OjFzBNPI5aNDO0HVLe1vREshCHTjt9Ta/qH9Q33lZNu2XIQrXJLy
Ju/GRGjzpBoInD1vfrC6PMzs+SC6SYNjs3Msn3IIzXeuPkek0ULOFE/x1IjAlXhq
KnM5kDHaFv4xbGmMUciMHlJxZJvt9o/wNCJLIHmcgIs=
`protect END_PROTECTED
