`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBOOr4lJNWYXhmQvcGn8ySvsq5G20d7WahbUvMmK2btE0o9yp8RDBGa3WOUpf7Zg
Zzb2AeivCgq9O16kIc6jZS4POvzJKwC5mwIrNRM+ZP9WpuEn6podfk4rcEYfuWaz
H73dYYKHSJ+IhSfbeV94PHAinyhR8e1fc+y8qRbsEFUaZL1owXuh6zw+yh9H2Jzh
/rqQ92S5xrk2yAy39o6IpI22hMC98mkfSzlwDk/M6+3wqPMsC7pBEzTLVdfm3tN6
SR8LX5kgzSiSc0qUE3PUHYM+SgfBgUrlFJ9lTmupAxTdOpriIizf3XC6gXhbmOKP
TznlQrxGo3sb993fJs1fXVh3myUg2TFfkNu73ZI1gw7CchK+xAsRyxTIEMVk3X14
i5UMFiBffmqXJLwLPdkeNyzVoFhgaDCSynPAHir4riJT9ELBrRCLcZSZ4Lydh+TD
Ed6QIh0Wk3avqrJdAtRszr+kR1Ks1mzVo5J6GfDvdTznVSTZqXQfGPKfDmT9JMgW
`protect END_PROTECTED
