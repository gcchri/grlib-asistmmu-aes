`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v/GD4Mbei0lb02M+JYGVq2WPNdQiM7g8O36gjyuJlzWCi+lXyPMf+qJWAnAbmvnx
XioIQJRwGF2ZIuUz6cJBn6t7aDBRqY1EoK4kH8aoHQI/DDZxToOnFR8dm+69IrQy
po9sCteQcZwZgNVk9Cnomk5q1U+JL8vNRQMJG0cHmr8oLmXtn4CiAks0d5MW0Y+m
2wZCKYKor+GlBTrdInCYuJNqB1sQjrVAWL7It7O5cT576SFZc/X6Be/fQPzk7N/0
Nn3dtL4lPlujoMfdtAOubNlRk5jq5ZBXfO7s+S/Ad9zNo0jHPib9rdH+s/frMofw
FT3qIjUah6UqCSdFhqto6uImsvzfOrgLlI/SjPlxc2dYu6Rezh87IlFoyXOe7j4k
GOF80UEnerMx+p7UDpBUFD6QeOGpdx/fE6jFjjAG3r02JtfMy5Z2jhIY1ktVGxzw
DuPyUXBAsn2iFYqvSfv+IQ==
`protect END_PROTECTED
