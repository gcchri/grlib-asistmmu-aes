`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4hl0UiNmZ9WUfo5Wjs/w6sydlXzPUL+xH2Ihs5IXk4BRKMA5ntbzSEsi7C2SIdcZ
c5Fliq54WDpuY0/IoFEslAEOp4T83HEQwQZ7C7DCbGfNafyVxNxGckkiDHz20pPN
Z6iXuFfIGZ/pQ/K3dMe+jxwDNAELpP+wwa9suQ5GJvRgDdFPjzZkCvppUEAwtfhP
J8yDv+gGu4b4UPYHMKY927E5S5l/zNoOESy0EDmwSKSPUPuDEyDOLzjN7A0sOiS8
yuz0IOtGtwUOVYRMq5cHcFSXLUGy4wtgwXGNb7216d9URSR47/5g3JpsWlLEaCx3
QUpkx/STzFFFHBJpEeNqIg==
`protect END_PROTECTED
