`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jq8BH5Yh57Dx+NKL5RdbdFGEaclYcZzqyxI7XGe4u91WQ2FHccz9nxmDearkaMW
0PWncxBnp6/A7+WefXj1kbEvlSU1KRZJ1U/UmO5WO5fNgILOeQ7n5Wj3hOcPeidr
lxwPB6DhBcSLLHMY2nm93n/EwboKPHQtBWjoxvQ2LVmN5h5Gyb7AmL0IKoFs5BIV
g1yWXogiGw1Lgrxfj9I2J95x7TcZAh8NVMDuUDYuWqtCrE7hA/b5m0aVoC6KrpeC
2HtWYKe3PivWucseODDGYNb0lGnGX/moXnuuakB2/IEbN1MROxImdyfHSDGPEuTw
eD5ngpL2rhWxc3HFIQrVWUMyWn0bF7GaSCPlSLYFlh4RR4Ntz2PEu6g83Ss7UlVk
`protect END_PROTECTED
