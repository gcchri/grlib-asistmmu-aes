`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cq+/2Dq+JoxY6dun/7Cn6xsRIMq2pnMVfcq5AC+mP+Kmo9kCb5Z/Z7gkIG/zz9om
cAn1HWHZW+iC4wljiwkfXl4FbTtMNkE5o1estEsMy92AeyQttKRBL09/T4R8d89V
KTS2E2q1NUP+6YIDKeKPa24uDgyPqFmBkFwwzH6OBCJhsuW2GXf8V/Ebt0MiGsoT
exxmav8n8G2ziTU+8pLpLLvcsJu/GVpr7wI/tZ9Yoo4EygBk2Be3s2uGEvFx11Bq
aFtOzNWhIjghB3J4V1BTfQyKAwpRbYk4j7hyQhHtIpq1fr/I8YZHJv8W0AIctefw
0D3dSefcMML65P67wRPe2ynnUG1TdoYFS1qYopSHYMnhNxder1CYOWVfbojKtA99
6SX8Efep6EFCVNXhfS8MV/Ly4t1PPWgsB72d1rR7bFqmVVHpR23vS9F3UnPs0UuX
FQbZ5BwgTy5+vsP8bpZDYUfTEIjCXpv0pMSbTm10v/k=
`protect END_PROTECTED
