`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S82SMHuB9OZqCuK15GohXOUB39dGAeFE5r96t7q4kaCX3erfEuE9ohpsBPnaUuyM
OIHjXSqk+EoYqiPE4/hPuGUYuo7/RCtjhCYU3KUup+iNfPMwadRTQjSFQpw48y7W
G+23Ocj83zgCk8dN26IahCgRmgKomEPmMniVJgDMey7m21Fo8pLjp9quUNumj892
LpUolKrIAN6uEfxkuFRoSvSCIdgD9wrzlXFbXGL+dmY4U30DDD2ZCVh33Kv6hWZy
+vrLu+4N8w/7T+BmgF41ZILjh5Xvb71oOpXWzzm0L2+7/G41vKnRhj43HIfU7znL
t4jp309z2dvrFhQHe5ZUl+oH0WUI7EBTzz7uHSs9mEo7jeWQn8bitBftqVUcb9ko
UH8tp/WbsIETPhz9+XiGlYFe8YyEZERsaEJN9yhSLWa3nUM2CqFezfLq5E+51Tbb
T5hgtUEG/3F8v/PPJglyU//ZMgZilHGVRgIpHAWkDInr9itsWAi+SoAnXs4gbd/D
XJp8LjEqWK8YPqANnkhU2GEsA7J94nEZgURWTKmg1jGRt63zQo6x6OdsR8c21QvW
vCC8ERppgEeEw6aQeY1bvoYtXbZz1kJBNkR8RErhZ76YRh7+1bSw2eCXtf124R1N
pBsc9WUsQsIcKs57uesfZo1YpVsFK+gQTsj0kO7qOpxkuRnXjmgNfnY3q/qDTAcS
5KkXXs3kWD6cJD0pNf2kU2EM1/u9WgMoXw5NgvHtXLXAR3+0R6iM+17jx94DQVPw
n3+awH2sayUzsqcY5Xi4xsTwJJyLPI6HcZb2dzbhZQTO2vxHGkKSmOX3CPuHQpOj
`protect END_PROTECTED
