`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iPsr7ftqcFHrVhLrCvcoSPtrxRtjCcHJhK+Je0IHVdW2RIhCqJNH2EXS+xj2VLi5
LXzZjB9l0UElEQkMVjLKoQS2GDLsg8uObGrH1Ptf4eB+GHSvB8GGdSs4JojWpvMs
kof9t3Ou+iqjaGhVuzXSe5K2ZrNFEd8Vb8FMfjQPY2GlccmDHTf1mtLtnxRlmBXf
+cLVqHyeaRlI2u/AwKvvCI1j58HcMX/9ChHjXzKgun6Pwh1FEAthGJeIdveQLteO
`protect END_PROTECTED
