`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2xtI98EjfugTLsGaDNuCaOSW66gx3Z6GNXVsDNOPdmEw3JKltzND3Nb6Hs7kmBv3
V8u/+eeuHPbS6k7OhLUgyS3CkWZSPHfMHWguf0g4nog+ZJyJSmQBtVyJpztYYcld
jX2VzhMj4mlSGvT+CLeuQP1XDOqcSS6yXfM2Wj0nYkctZD2lnP82jCgqneu28SXB
EhBGSf/vfVRJmkx356BJz0xSUpoIVo7OMReqpRkoGWZonZgSLU4A3tYjJMW9CNmR
I8GkL5GJj6ZJhFf4AtnaqKyJqNrVAHgHBS0TbaTmr3ErMlHUjnrYqve8lds5vxGq
eZjBaIBDV3Hwv0zsk7TnWOudMF+EIEK/jwzI169uQ7wOqdS6XKVhoOR3n1cci9rN
HSWY8U20yXLgFfaegvHqcyovfDWLGPZxf8SYmBWAoNdadxo2Q1sVB0vvGzXKlCtQ
yp9W2tbNaHr/9EWSloa/3+7hhAAr6YMKsRSWyj1X0jooq09aDOHfxeRgysg0FZrX
`protect END_PROTECTED
