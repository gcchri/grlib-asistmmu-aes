`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2yiwq0TvyXFhpiR7MGdWSEScaUCjEXm04TRv5oeJTUOY3ifzVUkH7REfoeIg4thF
nsX9+W7qtjyvZfE9cuiej1PG/RvaG85QuLrAh+wT4eVb4CzHqZ4YVtkWCv7R9s2x
UHBms56311BnckirFwDfNcN7cKiU1AiHRsMecVw/OupYrejKK9ID5dgCNVVNxUZ6
hFkuY1uprmT2jsz5Lsz8BQTUq82oBI4MxnRbOjlycIUw6E6z4hWrdVU0cLRlGNby
xRn4dYraouY2bM/wvvWRqSv7HJHeyAz062418BPYxneniJ9eg72I8fhvLX8ASE7Q
p+2+1Hfrz6r77K9KWNHMgKKcoFRDg+2vvP0iwKAhuANVHpXWCKVouegR8cupi70K
uU+LGIgQmc9AVY84zfgcObMs4gLOiAe0lgQ3vEdr/K0=
`protect END_PROTECTED
