`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Obth+XKDnt3JE//cDX2U5fd3QSiotEuuHkHlJbeM8+31e+04/JjzuJlbE/xUExtU
8WkAwlVljoO4kqLSzGvvAlF47Owp1DT36WKmr2MQZCROcRGN3dUh4g0qWRBIELf+
V0gAdeD5yL4H0DALyU9eb+AS2fVpUIn4GBtBMbw4TE91YjwbdnjnClvh0fu2Bl/f
wTTevi05BEf72dYdw39JvZrNNAoy2T9bCZp6EdiP4mHuG7xTFvjC/4fTvVDnZTYR
7DNE/aypIV+wPa6MaphdNBaxbgHaAORzG7t+PC/L7bTdcj/SPrNrUxfcxNv+vvx3
zzlMwPDK9OCrdXPWoX3sN4JsSHUwM5BAfZDIGUhnGZbQnKPCK7RVeSQxeqTHO2eT
VHxUicpf/8xB01MWC7wDsJD7yG1BlUsh0vyE9ueAtDm94vC5OFBoQoDIfJOeMDMr
`protect END_PROTECTED
