`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NM9h6U9tQl6XzvmPK4upApvuXm3pDGdaFf6CVpCUgWYjvZliWNYHKuCUS4mT5HtU
rmlcPzMD9BINn8MJAsCzH5ez5bpMW8fZpYpBD24n+kYk/T4gnIPvpcxB5xvIC/wz
m65vebpZxSfw5LMijsVQ4ZlVZuGpsX08NF0Svt8XCMscS3hePpn9VFsmOJRU2Bgv
H/eDgKX5W0OMFVaSMdLuONVPvHUNKPBj8dTdGtf6SRJbncJspAQtBSjcNNA1Q/UT
mR3eC/T2Tk0X5HvsOJO5rZc5Q8bpv7hDHt/6WuJuQ+7PxDcG+LdHavq7Xk21wweQ
cs9bwnERNd4VSVC0fTrRFUXE9A+HtvJqyCE68kDB0QYCKy2p2yjMLnSyE/YqnCrx
JHAxndCp2RlYt+AjdylLrsiNCK2BEeq4cL0DtcA7LlmEv15fylw4X/H8M6nWtKDh
qihtVa4tRIbHdLuCvr59jkiFAacDNVHgb8ex5S1yum0=
`protect END_PROTECTED
