`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wkcunndrXO2vX4+LumSXpQn9xGkXA0Do10+0yQFr7Q8MIth9ncdDG7n8tRZVNCI
2qXqfSefMLMHkvcmCr5Iber5tsgs9I1yfvDEerLqxlYkW8yNp2GA/rjVDv0H2NhQ
Ep/mK9tKeIbRYIvx7ECIsXItuB0xNvFpMIwrgsJu73/qXfayNZFVl0MmMqUY9xBB
Xbh5D7Mb1L02PLJPL9mu7GtmOmbEVBzrB6wXFSJ94J/Ux856OZ6JK8tOh4b+AGxH
82WgeNolKt6oiP2Rx7tAaN4H3u7SuyU4yOUM2eepRd0=
`protect END_PROTECTED
