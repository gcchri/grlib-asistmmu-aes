`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2R/sGY6g6WF/KIg0PnbTwYpxGwJN3NcGnS1yhEhhW+fcxjqp3zvk4fVELJHvSCa0
s8NBaElhpbrITXgOYAOTiCt2G7u4NyVUkeCUuVBPB9DipZZ57s18FItKXbmm67rk
cf0la3u7bG66OYfctdX2HuJQ/1vyBnpGsFAp8UGV7no7SwQlKffofKjBa531/aAO
h62/s2alWaZNkvoOlaG2Qwxuyq0CxHfK/SFI/wTznBnAgeFbmuGznLsF4e4hFfqr
4fEkgptk3As5U4ZwWp9uYILbUY3vek6yQIFJKx+Jp9moT20cbX9NXywaFX5q3ReE
JoUSEU3F/IvZYK9JzR1uSitEAkVbhEFiNtxRZ2NrYYBlGZP2BQ1RvUiH7mtgvaCQ
Moys9P6/SLiKiyZ/n0iD7x4tNxe1s1sfh5rHKgDXKPJFAWa29kEGsR4FHOmMm4bi
m2iF4sooKR5fdjVUOAVEwmjdpwPdHQ2CrpRNCgTlwRfM6DoqmBBaMhgHOLVD7IjW
ws5/r4+QEGZ1d3aKRANYXntHP9CUB+gWf4jMBBsbvbW7eyWgOfaWt+UPoF/CXW+B
9zMQWDF7bq/OF+0eaRvU2A==
`protect END_PROTECTED
