`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DEpjf8k+PgeWNm99qxXaeiE6EXXvz/wDaOo/1oiwtAO9L1I0ShKLyTraLAIcE0el
JhAPXolo52e0GNOkFpFRaPADXPXZLWXq1zIFDP6F31tYmcawIHAkVkkCzcVkexLF
k2Waer5Z8ov+1vwWijFwFfm6CzhkY297vMJjbs//wviwR8T3FbmFWFYH3tDUht6G
zgnnD2b9B5tuztDWjm2KtJeLaRsL5mTgfG5i2zfvORjwXHwBhlwDBUoJMgvNBeyb
kXPQAeKWm72n5Nt82urgysVFSVWQWRPP5PeW7laoo8gpyvso8+sh5DuEAvJijtKL
PMFQqEB2YVl1pzoz4fvKsTf0k7YLbcX/7EVstahIt7HgwhY3vgABjavRZF6SIrhc
lZDS0palZEhNgML0S0O0viTrErERb0G0kuT6uCFZiSwno+Cbj+Tc00Ig/VzW0vcN
3g/8tL0Jf072q/Kk0Cb4CezScF3Up0AiP00jUnBgWD4=
`protect END_PROTECTED
