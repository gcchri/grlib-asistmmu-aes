`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i+q8ipYLE+PiUmAMyXlWpB+6HzLf+YOcmNqH+jgfgVFqpxfddVTXqAg+TwLxp3nd
sQHVN+xXSqXahU/B8+fWEvdOFTO+D9PSDHcqnuJ2TvKsHcRsRC5oAPIhFk6i3x/A
oMT5rKQb8CgmaGS9soqslISJDuJlZYkNuETnlr0VHqagdubSuk7FzFZSi67sKJD8
dZ1kTQjZ+lxMHHHmYbqjiGHnLQ4lC8e7ARt+acVVQu7bzrq4kW0123CintNZcjf7
ZBRJJ5x4ClmfgmZ7Bz3N4xeaAiOKC6Eiy3xY+sMbaDpsHcLpIYb42RIHtPMYbrlg
X0oBAhiP7hrEoZbOAyKNpkf0FrtVUEhNT+jUvUuOKt0UnGuqYtFhj/AfRq4mX2q+
BN/2L8wORvsElieE3L2RYox4SQMsc8UFCtTRNb2JuXMhK4ptnQlXi2GNdGZ+YSrh
6FBKkF7v1nsYSZN8y/VLPpwl16oZBUaMrN2GatUoFi+jMWpjgG2jPH5ITKfS1hm5
FCXTL4WvCWU8qOotcpZ1OHzR9vpadLRCC+c1KgGiEyr+FeDW5oGNN74HIO06agHE
v3bbgKCBjXdVDrz0s+/Iq89WCCxoZt1EDCkPDAwLo37fK++En+YJ4uDiKtLQx7+Z
FVi/K7fzH8xnnOZIvNRv63qfuMYDB6559m1bEiW2W4H1zZf7+ovlHwscfUY801jq
WO08sGnCca5fqFWhUf4edvoDN+U7vR3uBE9duD85APH/yVrRK6kOAvFLYjgDE5jG
ittEVfl4bynXJWgtwUuqrNb+7GKSaDcF43DV+ycmmrJNO7gU6gj1glUxWEoR0V3L
hbgbAsrIyDuI4dT8IeS1qPQnqAHwfzD4MCRHeuKZg2Z5RrytpQruqXrqBhXJFWMg
rAez7oDxWm3gku74ltGio1hvhaib9eMw1HFPrpPCJVT2zBK2RIf667rqCVdHhcF9
45+YU0aQGUozHZIgfRorXzjw000qb8SpcxgF7r2QN9v/O0jQYWqGM8xT26//5fq1
6ta5ynjJ55DqA52CqQ/0M9ZT9/EOYAcgtZk6Ub/71cELc45lSdX/hvC85shbACg7
QoqJ9KqSfm5RBQYr6flV8IUn/Cjovo4zDuQqaKq0/zJKJy1uLi8qMZMTcdaKbGN8
no4FOakXqhYx9KDcXme7y5loC98VbmxumGtAjha7mbRPLnT1u5ScBn4+5hQvxAwR
KrDCeA6zxpBD9cHx+X2fxEv3ugldpMEgYc6Z1UvKPuqGM82WmXjF5EEOj5iTUfmh
nsP+hM7extZq7DMZuzTbfpslRa8LGev91r7MWnGP1EVhcjwtxNU0wnUUrc8NbrbM
PMxbk0h8/20u1COll1L0MU1aZNQG+rF00QG5JQpOWJp5d4X5+MGX57TuE16STvmO
DLOEo4uO4eD6YOOJJlDqlEfXZGZhk37vxwwz5sPxuZ0CWoVhe40zmNyaam5sXLdr
GcJQXub2RyWd7n7KVvh3r2ACnVGK18mxXB7ZHDNklORCRCokrhk4dHqyCqHEV5Hm
AeULGXRl60LVGjBnXBFz4SD/tlJzDsPQa/peq2aSizSL+IenAnQXgEg1W+nTGZIQ
lzP4Xllzr4uu8yYDf77i91vsiL0hlZQDrHPjtfXjBDO5APByQPZkNt4fZI3dIhom
N6hy23ADc9SwBKVPNYP76LFFZFh0Y+aKgwbST2MekmNbByQCIVgnvNUpUe/1Z72i
I0PcJQNQQQUEPozmstcEe6x8cJNRL8EWIYe4rYjZ5g/EIlVs8VAwIuuQAU4lEWcM
f/GSnHJYemSy2tjxyTJ4Ddpr5JE2VA3c5eICKiUkPSFbGrtH1oLnJU723iwGlp1Q
opFGanhp6TBjOTdw7gQ0l7s2DuihdN+t1rqTEreza4fz9j7riCMxOMQiPr3yAEAC
4gpx3KEWb9Acg6rBqQOEj9iXkCGHjjCNOc+bJjkIhsmgja1POpzZhPq/eOadzZm8
auhus6vqCxTbFQpmFLTuxb9uBaGnHEdI96rKpoVIJdWxVcG81eMyhu7sy+QhOY5h
UCoEGjEbVLy6N9QJPKY3uC5WYxBZdNPwyDRV130T/z25EIfzeqEwbcukYqsgDw6C
tyVpRBw0oFdLgqVI5T8uZuHgxB+VlkNRZcZFiysjCvHpuhbyGZrXQLYuOI3a6m9Y
Qsq//YlgRJ0n8+JD5AeS3oRT1k3cH0dwMtLmKlrNyX67XyF+W1QEVYA+jbtRK1uB
DyKZAsEC0HFq+D7fuJt+kkfSaO+dLjggVCwooKwGVCH5oUfdd4sV2sFzNJzJBX7I
f2Jo+dxszuWyr4r4DzBSorLPbfNP2xHteAgSzYi3xPIgKltRbMUBSh90PLpa1jqN
BLyz42/UHW2cLYv4qGAC0Pm9pluRqrfXO6RWQUgOoUkImFlv3bKbtb2Z4QzDmzmm
CzBnllu1JTcpsyCp3xlUPdRIbhmHNV1Qyi9eS7mPFTPY/56/w8BtjZDtbQn1WAAK
jBUuwwrdpsLi017T7cXujlKo1fHb551xjMwiSB4Bpl5eiD+25VQxgPUapPpJHSBo
FQtpLSndCCbRUx+FeNF1G6Q6hfzSp6baFVJLUqlGGPX7NPA0hFULmboIEWP1Y4Xm
ArGnD9Qt6SiXwpVW2NiEyc7M5ViDXxV988CwnQJVKgioS9P0Z+4H+fpsUrv0UYjd
YCPaJDt8DhVc7Td+1yltBNBN3guUSs5LtFlem/CNpyQ7rqurZwInGlKyAXqbz8pX
gtF1NXa+YEKu2o1xxHSpT51gX/SYgCNsui4z/FPUIztHb9z3mWdPrQt4xQWAdhrQ
hVUt1GbycUM/KrtZnvAaJzcqmQr9iP1mXXDyeO/U4FtoVjOBSKdIhZemUEZWhlMe
26lO9Rl1ZI5ehvhs6BW95IUN/R+nZZNflPZ1Ef6WAfvNA9JjZwif2PZe2NtCfzaK
IhDd2bcNDO/oISvCs0Kk7ItNtSF6nCT3D4D68alsC+I7eIP6diyp0Yx1IYiAZHe2
r5mJImRGoLAJOacGIz2vntqRL07FXInRwTNO5jpLfXfU/rfIXqCnJ2wfATTHuTrY
UKy1EGo5gMXu6HfS9MWhJl7kwswvqyZr8h0fUepz0v8fkv5kK0iIPh+MQAJ88091
HsFbTNEtJFEOxP5eUwVSkWh8EVYIxN4IH5Gpab4h4qH4W3I0cmfBm7rRomSID+hp
4FAblQJqi4STlPYFoiqjX/hTSB51hp+/GORRXE1KC4RbztZH5W4fY+0Y6myFiMGB
sbWObKaJmqlOkgTiYvH3039j796xfiOuasRskfAtwBE4NnbbI64gW0VHs/80dGjY
KAwA/bWxHNr6Oq98fOpZmg==
`protect END_PROTECTED
