`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9BRp13seZpo9EbMrhuEAKesakzojoLxiTKDLcnD+XnVboAwZXIwe/ajGJtJv87u
HFEhD1cCwt4n1g3yzrmhWda13PqLu0D6Yaisp4g5SASbjn5VIM6HC2i0xEJnLJis
N5dOvtRhZRUsgl2evIZAK2EvoGi09X2yL/11pI4jY3/k1uBc5vScGRtmFtShHvlD
40YOphuqG/J+BH8mTzBDxkKsCNZwg42RDmRka7ybr7RsBljnTWSaQ4M/enKLXY7c
e5N9iGRhajdWd7nI7tXiDhAVfUtPsUL4ajJ1Qdj3pIPyEYnJAR44WIHHGkCSYv9h
GQdU9USkcXNdrnC0UxXIig==
`protect END_PROTECTED
