`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
48jOgxUtV52r/SGWgaqgpwUT3wvKWdtH9KtsV6e5GQKOTjHvwyHj1N4Zmv6dY9vA
NkpUCpOndJU7/oDfjQQyxfkzQ5weMRqzgbF/CTfU+rYbOiiR165jhEkkfQ+A1fTA
83eB1OzDjry2bFC/ZfPcuHPvihwRxmzf8kxvs3jPecIS65jXw0Y9dEmFUbnqWw2j
Qf5897fq2/rEQb32/gqaZen4mFcPyEFdltVnZwu+UsS7g3Pp2mBcHNawBsEsCnsX
dImamxg67zdnffV5gq+LFm0DKGjNV1TP1dQGI3n9eHU7v9ZWL4njdOJRxlhIg8XD
b2hn/3kfYQMmHapiAj1Uf7UaVeGCPjTQf2EJQuw+92HckJvqKL2rSDR9R5QPhBRm
jxknSL3mfxC/GnRmIODojQ==
`protect END_PROTECTED
