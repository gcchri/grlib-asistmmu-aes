`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nzATe0gXJ1I0FwclzOboEaQYBIb4+LjnZF0KMILwE2c9Kwlww0uE0m0HME7tkDIY
79mmg8Iz9f13MQJsi7vh/RIyb8qymPpFHjyg8lxykBwrC2nkSNmWXolqg+WVD6mM
c0bSkfDE4RTTW9oKMFsTkOifMidS0odEmXOp0YTXjjSW8zDH638wFuwiN5FEoMZd
34ZZgmiEvVxqOtbRN5KbMMv6cYSY1C3UJbdpcSQr+znlZwS5z5sNbB7PWoFNoVmK
BgBSt2jIxBYVXhyHuvrfTU2J5i2TKBubn/UsPOUFDeW9CEpzd2kQJY4Kc/QJlR/j
D9D8VivYBwUoOj+83vsFw0flxWkVCv8pbaUj1LsRVilzYd8agXp1fLpfeAO0zdQs
MtTG3r31z1v2mY4WGQ3Iixh1KSWeiCFV3nmKdh4VEsSvRABbwqzm1D7podCPE2dF
25SAGAtXfNMQjcMs3FL/ovJkDhOHfZ2CGTK25etUE1ifyYSC362MUvsXTwuAnSr2
vjgBuo30/kn7KlznTn64hQUIJIGDPlZvXo2epUYhvofPblMcaZ+m8ptZ+ZhlZ/u6
5EQZEUr6razbw+zX8AtZCezSFyHtBdkHFOFrLEWhBvXxBUAiFrcIWh0woegFdY61
n7xHsIx6g8TqGDp2enXs+vKuMnW+DFrGIEkRwfJyBNKXUgJT2ptZU52O/OIyDHQU
cyOzTKclaauFcmtbiEQB9lSg1VyYz9OThHy/b1BHByt7YD/ICwbwAurwsYCKFZwE
sQf41Gd+cg79ixGFe5CS4+Ou1YzKNurmW/d0a056fk5zpwZwn8XbWuTXkU2Ny+qM
KlYNT0le2FHo3P6uV2Hb15RKBIvDoLG6lbQfDbQb2Lgi9qawE4ZVtsIbqeSbGmSY
IlPuOBLkWhKkIs+Jzs3q6fdp2xqG9NfiRbiZJgKhJaeyVRYRRFDastK/rhM8/J+H
QDuOKIkY5EmWGQU0YCOcLHUBmd8ZNWHHHeURHFw/YjyPhHY4dmQbIgs9Sjcc8oPi
`protect END_PROTECTED
