`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vLA0+ZOrfUag6869nC6wXzu4peGvbrNh4jOWbUENBzMGsKDi593Oq4tZGSrULedA
ddNQdKPiiL08MTwmjIC49hbVaVPcdUOyt0WtROCu7C0ZVv451CuPXFD0XZsK3eSA
MgRS/43d500gwfjzIA+wdA7czTPCv6f+ddUq1Z3jUbWA19AhQzlxNsgZpzUi/Wq1
F992l7x4j2etWZV03le8Uw3OjubXIdyEnElU1oFdk6R6Lnp5Wfyk8wnsXtOLbrRY
PleFAjuv/DDU2hyrmjm1eqDiK+NYUW2enkm4Hf2CfQYf25yFonSXjF/zvWffwhtP
A2x+UvI2D2mJ43pehl/BjXuzjd9Jo7sQCo8IUuRraLfV6NzKHcReqWiD0qJMHm9B
PuD/M67tBO0lM4lUYvyabAdZA5oxUHGCxydWulQxCqld1ZmrhskV6sOqXmUoTyim
TDlXyCHb5RGoAnI0ysdIga/QXquIOZWJRiwsoxnk7zLm6txagK+jwe65R6v5fyEo
jHB0iBaz1ykA906N6e/r57s9Sra2rfvRYIFu+HWRmL7dAf0z1lYIoIov4/1pGSNs
`protect END_PROTECTED
