`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rZStp3Eae6y5rnZLGnncp+RgiJuHW6eT8p+sEMTB4Ijn4B/i3TU7nRBVYLfOy71K
StGHoS7jBb91TD8fd8it+DzoGyBtdKlEDwHYmWO6fD6UR8rWKib1MCZsNHfsMRTO
QmMq3ib6atlV1uUv3dG04Ldm1sHnImwk70cKjQE3wNQtRGLpmWquvktjout+VJba
2lxQjMGXMQaxQJUPqh64KsZiNeu82EINGh/gQwAx9BSbKIgPqRHvnnHZYNPFGKlW
q50wyL6vC2HKe9M1ZOaLbQ==
`protect END_PROTECTED
