`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nDhXatk17ddwUfrBJQsRbox2h8urObwaV4yTHHTNBAIdZ3sc7L/eV92xfMyDzihO
CjLSaw+Ze5IlUq3yXQim5SzcNFcMm04oo2hCbq36nVcZz1KU71APhDTBfnQX0xdK
aMfBcnHf3eIMjsM6QZK/TJMVckbXlPqn1j+81i6z/CSCVWmcAIowOBq5Jo6s0axQ
g5A5yE8wgoDjPeOo17KECcervgh9CpfgcZzSW/TB2Qz0Qdr5aP0ezM0hhqqRlIVj
v3udE1HmdZkynkbDuMZGSK/RBeDBUKnKXXDUYAzEtifzpyqNgyjG2BVgSpIaTNv3
vhrf2YCS58Ep6FO/Pm39a0Mp78YMaFg5limFrjVHyTLDIR+tVHAGDcHuVg6R6Gae
XNW4kWGeoYXtfKzI2CkwJv07ZlXyQMLr72AEwrHDzXvRA6RXNmaLQkMN/QvVjrSU
j35jfLUcv6vWE1EvBXlrDySBwVSSoCBJNXnZuEJ3uNVJDk/GLP5TyyKLdymkLiSl
pm+gcFyADc3Ts/MSMX/SnoRS3nHdy1+nqQrxwny9iaq99lWUIIDQ1/Jx2agyXEpw
CFbaUAHeyAAWacNTd2Fh8Vp8CvG+gMD2dQjl+7dYXQgS1lRBd1poNcRAL+nnQEqz
hlAYSR6erIs/cjgh3YwWSgEBo3fNanWh03FsG3wAzXWTpcWyseonmUOesBgA83IU
jAdTyxlXwnYlLv8P3GMau8TyVYdV7MbeoH3BT51I2TOb4y2275R2mbhkOsNaMSrW
1Z6wiVKJTIFi1dzlOay9srtDhu0KUKZKCScan5CzZWCk9oi2R30ioc9mCBJNDwmE
vb6s5slTMkMDr/svaUVgX26+ktQnzDopabG2teAAcJbD3zBtPqIXtt4zR7wNb9XV
ISuOJhtYMhqJyk4uUh+dI6CoIHv6kZQc7J2RLjQWWyb5UPi0yuXQOZcrNMmgWFcT
EGUmFmdA1AS599Ce+yFXzjh7+YyquvCSlAnXoJY0Q2Al0I5QkU0zY8sPle8enCM4
1oCPz3y3CZPtqVgFfF4UqhiMVMxm16oSSk+4nJdF23+yH3i8DlJP1eMPaTYwVl+0
8EtYFoxVF0F7K189HAv+nThjFa9ehHpIqDRRYIivvBoYqN3mmpdn+kCrGfI56eth
WfIEiSq7EhRNwrGipE6kH2VvvUptWhnReD3ATIhQLgRasOV/QHe3FR7R91dYRPh6
U/c9uurez2KTkdwKG1wayv+Tlb9A4o0wHac526bDcaCPRdb4smPVk0NaL+hJMj1u
+1o31XNrvS3BbOzSmYwXOC07mOmQEEoxMLMkNEr6gTtkjtZxSkvJ3+UZeu9c2Aou
JZtOFDoGt95fJWA8luC6FkqS5EHqs07rRHBZEXV4IW4FgY+amId4lpGbIZtOC418
SgtaEQ7YhCDbER46U9mgA8Z2+g95mUEMpBaZgYr1kr9Ij5EVn7YUk46uQPA17iSC
Eicri2QZvfIHj1D5McqxH8ZRcN5yDA5qXGCbnSrw4ygi1EQZp/TOfLim6D9tzA9r
DLd9a5HBYqkFjfpNqIqSVPyZEnfh1fv1baI6IuEMrZRfOQwmwCqApU5qzh+RNVzt
uen863wHkqeHY1VzoxD2bC1MLN4ZDQJR5ZzIcXjFMElnE071lqBn0BjEPTIZqCI8
Mj8FrpCT+SZPYJqfjIFIwwlxqwrCtNr66QXGSbnda7TB61HIUK5TZIT+sQjBexjY
hOhP3WduCxkphplzljCiMM26Oqq2eNVIuOb0wfs1HVs8MIPDZdvwDdYZOxqs77FM
AEceqYqOsfyRFhq5gUoabUk7SB9T4vH3Vji0o8+aNrWtqOxqh0RL5pfMfbHhOVAb
dXyPZY5Ne32Hc+OLKeJKoCQd+FE1C6IWkGQUaVhLHz5Zr+Xlh61J7gpsb8ie1CYZ
nNQz3RVB9zEzlU2gINd4vZCx1tnbVEADlOmDOFd7O+A97F9umkWk5WQOXwXoZjsH
iKywJ2G3XCbOJ/BkiN82cSKAyIPPB+Sg9PY3mP1oWRHP+L4Xb5dcOGrUYt33hdTl
r6GIInI7EmL9tGNitWqSy5+DzpQmIzaEyKFnecCKgE81Sw/6Qh3O6V99dDLpTbht
HS4rjH7PS5he+xU/Bz/bbNoxbQXBE8o8SyMVza7YDLDMkNGi4jxjJzgzaJT51iqy
dgih5xCyNkJ1B7YKvsEX2pF8Lzz+ROvQZM1rQs6YN+j2Eq3sytCnT9ODitZsi3r7
jaMVi4nZAeJRQ9ME+DC2oYwmaBgPhMgwAP5rvFG/8b4kfmshbL1ZoB34BnLqaaY2
51pQdFq0frRZ2Xf6BH1D9OwXWV3O3TfO+JCZJCe7t5VVKFzHxE0lcXq4hM82D+aa
A8z22xDsK9axi1iaqv3VYkGjEvB6yhoMGnGLPcnAKrlJzqJni18fNwZFPYqyDqNl
vl80Ib+rCvMcR1pwC7xlOmGQTvgcpZAi0WoQ9++gUya4JYfvSPdPAaZjXUI6NOGk
/6R1uTM/IJ8B/e+v2ISY86/70yMuVk0VJwWgGwj7IU3GSs0f4EOBU17K1+Ljig7b
Mrcdym3em8nnPVZ0EbeXmGMrU1rNapxOEqinIs1q17gRk1pzVHUATTmbjWFdXqs5
7EJ0KTzjIgA/Y7dK2yjoH52pyGU79jqo3eWCnxejwerqxNYupmDQMcqqSy7nDmNK
S0a+Z14TM2SaHfa7Kjcm2Tw4sE7YOosCqf2ETUqifoe1xc6P7LH6DsUJJnZJDfLz
qVxaw5vzSoLuQGed/yW5oW7ATM1MmnoRo1LKdlRFmSBczDH/r9Wm7Dnx5bEaM33U
VeuZXwz1Bykt1cbKdMFd3xNiwKFgUB8JVRC4cXiOV1lq6zk4Wbq4wVWPmGXog4b3
1A5UBcFyMGk3C/Gt3bSTJyDAuOPMPweTLsBnpimy2ANjnQKAJGsGQQDW6NRgIu2F
dlUwxE6RFJb0zAnE67KUTlA092g6rSzAHc0b2VaL2sftD0ZOBMfEMBPpOeSCTpmz
C+X41AZwMKAVniYEE7oRIPncE5uKGOyk93+4HypX+cfzJz1eClG4Uzh//a/CjIIT
SLLXhJIUIJswkSnap8Yly6A70Y0VJ6p/zYzZDMpzB2J8wACVFxXcCPrWSMHOkdDb
OXWQ6g/jr9MjtR2FKh9kLsciiseLtsrEvjxvCmsp7CHh5y5kY5kdQadHb1tHPt7i
7UeQjq8BJTXh7vU5hOdr86VDehQxr3Qq9SvdxpL7nZ1eTgf1eMMn9bfxfuKmWAb9
odGd7SyRA3OM8S9qZVK5z7uFD0Jqj30R45dREQUQinDdbvCtv4IK5teJ4/jfuxIV
BBzXif1+wIkoEXDknNZlq6z8m8xi4Kkomwhw5Cpv7C8+RR2jE6tU/EFB4aladn56
+JrP79r7t/dqYhn8+yyHaulULdVi09sxx9FzAPW6LTx8Ug6UJKruf1KtHxFPzmJ5
lwlVpk33nsv3e7q9pwKu7pzS/RcGllx68aF1BSjK47sytWid48+xSNAYqQBzwKrz
0rClX/zbRVNGtH+w08/X0YQKam8zMOVFDr6dKfKma+62krkV65qGlPVirTwKFnol
vWbGTX75nWCz0pty61YoKqrUv+tV+n+8Pg/v3+pBa3W7/MP6xF+tKCP9qt3Mycdr
D9pSMkyEcGW6edVjikrzMjiaLITA8kKBVHnDYltZ+ai0rf7xAMC/XwcsYIOjnSir
cvrSvOLQN0aZF5r9a1GEimD3RVqsepO6raJAHV2QmHUSC85VfcZysM1NtcfL+WNJ
NLqWkG1wvDFtwYUIBoicx179DtPxGjkCbuD0X1MDu6rpQhPZuaJt5OfwI63pH66N
wdWGScJZEktVjbeDhSWEvGnp1AUGRK8vhvLU4OV9kZoiiHO5tBm4dxLDiKxXB3VK
D2Q1kEaQOG7+ojO+6izLRMGzJ18XhB9EWoXaDv3UMOLlbZTL59y3zSVBq/75ipww
5iIdd0f0E+J9DiJlWd4MVWHPopR61E1vxp/wZEW9aBsZhw1ntF/3/4UUUuLlC5yl
H+4KWLdnNqZqw8vxf/1wS23p9xXUR24rfVGJ17yzoETcuf9npZ+ZD/qrVktM8Dom
jSsLpmfa5HlnLUMIYbdkYQj3tvUrY2hsw6mYyvwhZMFC1dqKzZmKlUDnkQFatnVa
U4DD7DHy8X/AsXBvdygINFVlAOc5PME2C+Fw2W3HzUTzk7BXrWua3WR7zTs8NGJD
il6YeaYoKR2TbcLqF/PxOunBgHOl/q5gI7UjfQOgewv3NPlBkqexyYz5EJXjHgEw
NEh2s/ZxJUORxv78Cjv6+IrEZacMVTysxRKKUHXOUDMk6hlJ+etA7u42QNeU3vGC
HE3k3qV4e83EIx3PmnOiyaw9Uw0AR5Wtyn+KvQVHNkA+fd0Fx435LoGpiorIn2bS
IU84RzJicXPjMlvAOODe7+m1mW2rl3571NEIZ4NiddZTj7PDzyhtHDupUBh3wAte
0nDY473eEYbgX1lOn4z8YOb5oko/5gOFfgxI8mLczDcf66Rg0jzjhpgwTsK8Hw4v
GmCSlHwofE9dO11X2A0l+IltkW2bcrWVIcfAuUQzakg6ApF+iO5tybzNXuYXhDYa
zqZK9JBAKWMwQknmYXNpsmhchJEkriZ212PoNy+DOhVjYU/CoTCAE0jrKVyUmibY
nwlRQlob5sTQMJqT1954sjAb0KeG0kEfhTLV9yJvPzvtz2Ru5jhuG3E8MhwP6Qbh
iGCG4YIN0Y5Z78t6Kd/1m+IQfXoQzfRuyuoEMQJmQ4+hMuSJkZkpNDsIIomz5P8j
E+6B7wcHdTtxfGxPgtmFilZa70ObTLjLD2RsKAD+ja2w/vr9425vgUcwkUd4LDp9
t2orNhX9TnGGc5G6oHAogjSh1MkiZvXHkSlu8Fd9IPvvpGm76U0cuW7FOesNdTZh
w7GurnyOM8koyDuSq9lYOTOY/sb9gJPbL4atuA3257Bi5HFnayIn4bX+1ZsaImPa
T1D8J57MAWAMZrsKH7ngd9+f/eir+O8zSWeMvdvXAM1wO9hd833yv6XoezcggQbD
djp0wdyQ4XCQON6YbNlzH5/iO2S24RDGj+1VPqXEqQ8DzIgBJFX5Z6p/TjA643Q2
uYHX5Jmq4GqHNoQJSS21oOm3VAbcSn52Uhz6mLLfaSG5A0vPCNgQ17Q3aOybvMMr
s3dJBQePkCg21aDWdAev3GFj7E7r3YNLZtPblwZrck8uOfe76DGZpDSfsthRuZK2
S5dRrO1um1OAH8GvZBbNzFWw+wL0hT/lE+GOm0Xx7EewlfbwOwFk17LQLhr+ane/
yspDOSOk/dJjDWS3wW+6h3cRi5JNLF9eexg8Hsw2W0YV/uS7fgi/X8hNkBi44pTB
nLEMzN5PMmbEOySvm1EmZJl9pY0FELADsiY93LOazNeWPh6MeAoyApi6Q/QS5WzY
5gEYZvqXpI1x3LwGNgaePLHxe/gF7lbh/uLRkl0WbjnmfgPis5dkSBAti6vxWd+k
aUkdJ/SP0waFnxZpUYPb9s47ZScVep+0fw9HM0rVOiXaQ6KW7VIBvXIMx9aGUAQ/
WTwJqOW8vDKd3i1giGqaJnWq35XNog95bMVbAanxWFUx64H/9KUdxpqMdY5XCArt
9PaGtEpNFnMDTb4lI+N+EQMxBVvfQm7l069jFMTnYfcV4/FwX+UKFf0lf15xwBHO
pJa2pOQ3NFoiTZG86jr7Ds+V+mNLp/EvvnV4Lad6nY63dXxA6x+7FLd3oZu5nQaN
hB88gMsE9ZbKGZaOjfjzYWW6uG+6QDkKxo7V74WKMgZsrMtTSMw2mdo2D4TGPGCJ
fZeqHe1ydMmm6AS/pl5EK5dLlnYevBkmzYqTbUIiKJ7wZ/E2f39jg+IA2YbGYXvt
5bSw7/JUhXKvRz5TzBemJOY951YFbU3WpwcBCRcJSJa+P8zLhPMNjd3H7lU2S45h
iYkl5HLObYYQBnaWfvZZ6q7HfAPSh/WM7AMM245E+8w8RT0JkGsVV3RGH5/tvgcg
XTPzgMYx4+hrnt332BF/rGCXWXJQcD36cWiShe5kY0s2hfpPoZHFFiQLpnd32HfV
kY7KTaxfT7dapsGrUsk5SxSXFU38UEqeKKtOpxcfo9CDVhZSPC/AEjqTzA2a0B4W
udrCKaZt/nVXlRltdD24wbhtRV/b1NbC0RHTgE0OVX+IZXuhJTEJMlWlP934TKY2
3ea1VkmHqb7VleN/wzGuVz5cQH346gEWQWOAdnDdvtfPae4N4YFGzgPhn+zNbmWb
LCX2PkRLKdAhL07ECmgbtPeHV7K3lE0+kgDlOGhj6nEe1I6VmttKVvKzc9naTAqo
ZXHyKN2tbFCe91IXEbcXe9M5mwcYKdwRmVdgozBnKR2ZXd+n6wS+CqOELDnuZX9X
cb/naVXXdZb1QRbhtGVfDsKIty3bBQF+a+uXjJ08YkPlXBoWtVG32UrrSSdncTsX
6mD7byKuyB/ccQcgJvDt0YFA7iI1r+DkY6L0QfCwnILq5a7GBBfRywYcyJU48Rny
AxlTCAiB9ay5UgKS31TDpBG/jDuNBE3lzrp07Q+EhhZ7bMOCU+g6y4PQvvj+V73h
Eg0PeZ7gROBfxoiBqOcIhZkRt4Off8oSf6YQYRdgPEpgOAcC2gsn/sNnOgcc1S5f
d73ezIHPn+1XeN8KvTP2ZGy2DS5UUQkB72jTypJDTKoiZGHqAMnV1POF2NZfrY9n
+AeEE1TgsQt6bQkKs6rcmv2S1WTeOhdjrtjAWoxYJApXilGJtYzf2O8hD4Od0zQX
6faFrQD4wy2c+Rv2eVFawJjSlxXLIvBPmRmTWDj1n9uSz1Xtkv+7yoNdHX6gpu98
SrOBii3Y9ysCLtwd2WOVxDAJzghucODv7ldtujTBKQeGKyyLSheBCeqlCVun9mFF
KdYcymvue+Z9d+PqJPpYqrvuMeroRdFdsSJLap8zsdpN47Dy5NzLwgMT6+VYeZtY
RlDdKwNpH5Ul6JZbghrSa4J73IIOH7GH/jNRF9+kQCWF71/AQaTm+kJuX78C2nEB
NJKdDVHz+JSn5qQWnAnlvxEVp88/kEJnWaVljrFNgw9SNIWyJFs3X9l5vLMDV/YV
YkdzfeTIAA1vB3zzhgYqf8vI7EeAJPxrqo/eLBk5Ct8dIweLInvh67LgogZeBBJj
aIPDjBDbps0xChE0W5tElTRaHNHznLPShxkJmUfY8ofm1B3uUwNR2OMOOZSXGOIr
0Oh9bZ4Hsqz9sKYQXdUph0piwTYUFMdPFz8vM9sXsrkan4JxdazqDfry2u3paTnj
Ad6A1jmqMye0tY9K9kJYKt90YP/Fagim8fnQjEFDpgh5PAsjM/9KXnPAfWTQAN68
Rms+fCZOgRsqy2khGXcNrD0ROYBY4ouX3CbzQpUugI3eR5DfLXr2ajSAKSp2ploG
Z4oRo9UKCOBfFXEWvRsBWzK9HppgMLyevfrJjrccKGloqdoskZOuNAeehLxZhHlw
2DSGw2xPqUQkrNt1stOsntwrbwvFKlMLZhntVcAkq2Lk/SRsCglolcMOmkwGbFnT
k4jscynSDXYHHKFkKUBxAbAPdKBRHcOmdr5H0vgmgkFRPuOsinfgxqIelESMlQ8n
1SXKLU9rtPwsDmHkyNwuOlB1U9FlWPwNZC5d4p8uhNIs1F82aLjFz5LLRfYtS+Vs
CSoLM9T61miuDXcy7czOZG4c+9bQu0mTaXWUFTG2wVEKLWTlbaV0QlTpngKgpeiU
biAZRsT/3eOry+mmDSSfIkeBXydu/aStN+I2kb2HWJlAjBEnPwMXkmIkOYZbKz4j
zLJYp01hxM0k92mYAYsUwQS3PMExz+/As6U/SPhISvbSrQyjkW4bmwZKkrnTTOa9
4QnWtk53wArPb2gfxO3zv78B5Qv99t8XQVGj4Nii3pRiNOMXXvfa6pnp7SeRMtc4
PRn/42z/n8mOB9laiWvPBaz6SlrYBTSBcIV4UbgXFD3FwSSIxb8ybC3IGGFk142G
pbxyRWCy/ZobWHQVxuhvKVVD3/VnLfmi7qAxlsWAm1ckUVkrypZapxHqlllxyJxz
klptvqvHGHxneMOBepqKaxbvOhHwNtp5jPR8YypLfccUW7b6MOSS9Fgr2vpQ0ueD
+lONpgGzGOc9RSBMEseKj3Qz8TbJNt1iGqRutUuOHPZ70TQgXELVfrbENOIPVcs3
CRYrYv0pyEX/HSgYaZqfILKOEoSU5DYJ7R9AyRJa+s2NsPMK8WMDtOQeAWkY+VkW
oCn/jc7Wu9hkUvVscl24LchKHLraNjUQI8JaxSndRD9aCqX9M/ken7t4QN3BsB52
4PZo4PKCRcXPlyEQ1MFyn9N6NKw4wRehAiqOI6/JrPbz4vAz3UgS6okRCDsEGHrH
/5s5iQW6q1YwP8zm9ToTtLLvAXrGpcv7Tbr8/BF/ncQYTmlzxfZDbQiGpYqJFtFn
ec6ehJLUvMnLYEM7jppxS4XERB3c07j7vq7sx625Pfn7161RIAfabqmG4UWie2/v
DRFWuJ7hVnidh9QC7HpoGZ44f9FBCa6aAkg3Qhha+8CWmbgG2olVA8nUsYtVIC7J
R4RH0tzIbCFzzWUaz0N6rWNY2EIqxJbbtrGdyYuHhTMpTStYAOtOyPGLetzO0NR6
p1euxvjTc2KqrOmq3XcejjeayPqoHO17hJNDENKZdsyxc1uI1sjwupkHdQ2MpxId
f3nXu3D40ikcGlLU2IS2AZjq7i5OcPQokFw13Y1687BsKwptr4jA3DVZsClxgbz5
23r/tvPyqAgTL5XguGKsN9Nd48qMx108dnUsASb6bUYaODMVm3FCVQ7HaQzFVK0M
5grqTnJ302MRvIjIQX4QyBNg/V3yxpQXEgnOqv4OS7Z8iq+xbql8BZxnG5uyhZNO
26QxLUWJ8XrbhoLKGE3RpytuqzFZd8ByNCWCuOpae556TPoK0FeuKVrAlXQsSk23
z/jJUE6bLz2p32XfqbmaLs7xM/LyOfPrjCE2mQX/eoZox0NvfHkMaRCr3c/5MozQ
Q8Uctw4HKR7bMz7egwSR5p27BC9wMLDfudF+10eNp8oDOAB/rO9IwB/BAfW6jlr1
VK275ITkuZNztUNY6vyWR0Bo6Qj9oT+r/uMqU8z0UXiGSCiOMRxiHb5d3Jb8q+yK
RZNCrk0ESOGYgP6Gr2LXOo7K93djhwkbqSPyKZM5By6ueeYAUv5PuUweNDwAeV27
3eed22mw37zqMx7CVzHjKs110hww8BIHsMo2SyrcNgfVxWjc2L+Tufa1jZVBiZYa
uv2ynu5r/oOyllUTDUl1k6dKxr3wja2kZPQO1oRfcrDtD6EB6vKx6EoqZJZHaLSv
yb+lpY2vdae2Kkzce3SKWzPobLEt0tvxyUNO3JV4+7NeOuVjVIF/jazRHy2pPADd
JKsT0s7AaVipRHU+12CicrKwvt3zJ51i7p2CWEXBwPnKua2m8wcpsWh4gJe8tHZw
kuIUutNqdzVYV01UrmkehNh0vh44kb1CLYQkJ3b5AbTmPtafdZFY3lOUKjc3v2WL
G+vN9ct5lkpWbYpAcKCHEp8Dnvf/ZMYCt+XIrR7QF5vlk1679TQzF78CFssrjQAF
2bnUrncA42sxkcG0QGwruy/yBoc10+H//wBlQqvFNVcWSamwz3oRj7ToKw14MH2r
XvknKLLd7YSb4nssmG3rewZxkJWUGEdxZjH8lBuGgdpDorLa5kJ2aDLaaT96U24M
sJm9qk1w4f9N/fVO+2KRABbg1GSdGmL8+lWchHS4Oc4nCPHij6MDB3IdzkpSkSbE
TkfoaBqZfKP3OOhu7a5kpAmRxuOjSFmIfjsJs2M3tZFs7aL+J4Au5ZClDaTAQerQ
72VjAubenWpQNPht/+y6rN0Zn2F9X/Mf+3yxmsjGc49O+2bycLMqQTc21Eg67bPt
pM9/GXfQOJ/Jm/Crbi9q7dIS7rl5VoU4VNAUcXP5CvpgYtRq377+DFViiy7DoP3S
B+r3p4tIHIIpSuxWHvsk4uwY/u7l7UPdiCG1cPZI3QFvz261ZddQXBjh1R6rF05R
W2ICeQDFiVxccy/+clMWjr84z9lq0A+Iibd7XhlCuqtU1qbcA0OOrmWcmfYJmVIM
2vn2wEiF36lyuejzGv7VQA8gCgX3G4EVEbtOFQcAptfYungM31NC+Rkhp53Lj1qY
IP3UXzjY4jOvUQlQWtT0BZb27C7n35x9p1dluq7xF81196Stk8MhmFouJsYIxgOY
M0OqyZj8hG3DMBYryS6uosD1P1jKRaHqjp0gJdLooTWgrJ2z0yh8FjiKjTBjjvbj
uETJdqOfZ1A2mUP4ud1qqnXVeWEpR6Miz9bhZHp6pMy1+lOAxFLgg5Hx0lSbibUQ
HOmHGX9wJmI4sWv+SYB5GEWLVaGWfW7gmYGRujSBLOkbQKn6BXgpTXjs2AxEY/xC
7urf8Z7UREc/sH2UeBDC9KLx1SiC/YMR/0k3rgB8YACCgzQYgLeQ9MgBfjLrjmSo
qI9GSRpCKm4emndcSCi7kYO4pX3drQFuSkR395Aud3SyYyupMMq0W7QAvnbweWKw
8CCGP1EqRsukqsuEOqJ78Wn4DU4v6GJ7IHIiIC1kDODasd1b4h1UqUvrdEfofIaD
uarJVrH6ZBIIh82XFza6ACO27+t3lrD83Fxv8BKKeZBSa/sLGT/BvnimmZPk6E3H
T6snggL8HrGMzV1d5FCZojtz9bWRjHNDCUpqOt55EImzSY4rs1kERy6to9cVNg9x
y5opuZH9JR7ZnqVLjWlj1GwBVv+umZmWeWH1pYzEwi784UFshKNMhiZ2WAiph9AC
+JLlURLaWu1gLJesVzNfh5rLc+XOmgKw7ndlcfqh8IILbXYLI0CItY68lYo27C34
v/zgvzPaObQ006wN6S4ud8VqYAtMgDJ6i7bgVuPWXN4KWTtSv5V+YVbDxh/QdVJV
dfkgbmR6QAuV2z4nu49Eqj/9bGuKXtzxt6gJJglB30uQFX7Cx8sLymp+S6UHjy0J
fULBH8iF6ttttUlzMh3NSxJcxnU9M4An622dZFyRZasRRpHxdBBZZ4a9CokKJxw9
rXS4uzU/dik+8lvbhi5gHBa2ie/k5jSstw/3DreVG7++bE+7xL5S8W8eIUbV4JpA
BjLOBWowGRjlqrL2jM5gdoHFMNNtSztfG7CGpcs0yLQL/9y4O2TL8LUqQ4qiYSpV
nO5kP7ubI5urP/Wlb/8bch+k4PwwFlz7JdSQmq2LafmnfDSTKHz32btS0f5+3r+R
ovO5of23kpKq63vdLA4jIJIipsnrGpI4JlWr26J53aPmPuAu63LWDrJaid/SXG6d
Wm4ZP3VC92Ojw9rqimQpiPd81uow7fdBVT29kx3r8goJ6a8/oAAbz21GSsKz6nHM
cmZhQNp/rR2q41PScOy2btQnNZyaiIMsSBM6K0yvrVOteZEk8+xnh+kOjuf/Zi1x
d82FyxvhQHfdfMqGKfVxkEH1+2aKB82bK5gDcY8v+Vt0e3nYEB2WW67DkI7pcJN+
y/CGkIZv0IKOe1U7xmOxIdj2g7BMfohIh9KVrwqcfVOc6yEoi3rjE8oqGrNNog5O
myEOASw9Kiqj0rYzTmBrTMf9T7slEIqv1xP4N+Iu672sb3F46z7LagpOzTXA4sJy
cYP85ykHXdjrWRzt1KvV4nYnTurqw5q2lf39BnXkMp/eVnmo8beavK8UToO2Ry9g
ODFCysWgBo3kDNLSpi16J5O3HOw/achjdctFTl09mH1NQViQo55Sl2v/dZCZMN/l
VQkpSz9cM3fJtw2QQbduaUCpS9asqm+dQ+uSYgNL4hdf83kP5Xr30n7aSQ0DbYNr
W/7mCckjlp8wj1FP0cQx+ka+S2f88wRRw8CmoBEs5el0xFpCtvHDWwBBC0TDwOem
bpAt659mMysOBwzB/tVmHHzQbGfvHv2A+CU3zx0GbZrneqtlzmfAhseCCEK2DR7O
aFDabQVeKgbL6uLLbh4ohb3SBxxW5pOeQkXnBj7rIht7bnGaeZkFa1Es6R9ZLQ0H
JKaHuQKfUFWbWnIbADpueWyQhvCZQIlxdOM2cJ1CTG4R0F3REw2V3VyqAntSbzj2
bgP9wxBWaQiWnqOCKfkus9xTMie7r//Df9A65JKxZm5Di2NHJR27bFSJNoIxD74n
f9Dq7+433y4JQCkJlCvOlSsujKu/ItASoB1ago1/SFsSAAM0hdmanF93mXaEjXIP
1gLZQTCINjwv4AFlqTI5M4oM1uCbhHz+nj/nvLszeWlBm0DIkzHsN3RaZPRFvjYZ
cfnW94qiQMxOW1auCaO2wa0VO6iS+sM01WVA071+HCPSXN3PAejnhSdAJ7IpHv3B
7wsx94EF+cd5yNjk6xefvR95FYoGQbyzunGs1gCpbM42byZ838m/mG+gL3Ye+vFa
jdyBa80KCSfoZpXzbSJlTRkY4YT3cQI8IubJi5PNtLGiCWcMmFANKGuZVkwEQjvf
0qb+Jsjy9yAW8J/LbcXmBnECjTXjByseSxzz5Lq1xgz2J5jmdg3jtLY6wkdwHJUs
F58GnEFrv78hemfGuTAJmnPNAw3trZHPm1BGhDIr0vZwcJiYpGZoP3GhBg8p20+F
a4O6aY1o1q16Y6DAN95WaJlFw1wniMe7nf4oRQwIK3Gh53WG9ftcesC4AucTtl/T
YxlqleGKXOaehO1bViZ/7dqL5uaZYKyQ0ta0FI7ib+HblA7/3YPVNzBWsqzOFCtV
XRezqgmcNlEUfPUdCEgKkL63qNRHmH4YYQPFVkLmp+E0R8o3LZx4mYahZQtrYsz/
Geg1eh+EAs0PZbcrB9Zx7l+7hP9b8wzCKFoAThghI9l04TNTZZXybe1F55tZbLis
r49o8VF6Ak7n+XR9k4cUtHivlxElTJcXLhyTmBx3uwM9tYitb65PrXG+NM4kVlmf
NIkLaLozT0Zds7OK3DdKk8HzmQ0cUtZecqFzqk9QNbWoQNbA3oNngLxROnsqWBpt
OaMnM7qSv58N7Q7RtIFLxXihHiGFyYCUQJvZv8zM1faKtYBXIxoxFCJx2rc2BjMP
K2SEVtPNs3KiKf+WgzlAiBEG9XuZyQBUeVGOIzvGch9npJaurg+CgNxtH38fMj7d
2MpXsBcgcrCzxh0Ozn4ZWml+mH1YE3TkjRpGrb+X0do66U6y5mv7rxYAVSJCMDRd
i3WL5zxJj+pzhxOqg1kGBxSSumJI2k+gS0yE/rzDNxAWz8y/GX6INVj286jxnnCr
/MORM2aj0FhllKZlQMN5Z40kf3mwxTOJaUf1c5PZ2vowi1ptrw0Hc6nx/L/8ZOUD
hlif0NK0UV9w29jnkV3xHiMF8sIYbqJ9U1s0wBx1TeRVd1dlj2X6rwysLBDH/LLi
/Xok1jrRiDQcWEz85J7C6kiTEr/FN53WR2RZFk4zawk0d3DgOZ8TVPk2s2JD5JBE
b8vT2fck2Ot3jbHRDnhoxDDb84Un5prsctIwdvFeaFf8VA7QLuwYDhMNLnEAZHgV
ca0mVhC35ivHcbiNquc2Yjy/HWWl0eDVQybfMs/p8fi47tmI/j4g78rJvhnbIEil
nUKqhBd7M2HgiQj2s8b+3uSBa023yee4wVdYaUsiuYyPRWjKfe2TxcvHHtzV8u+I
gnPFF3qd2tRtnMugvA3Cc62+TPbXMqedPdYYbvD7b42bwtfebKeLRpAWVKYLXONr
5ufCaiEMbA4Z2t0dTLaIm2zSKSURM+ZYk2FttDACjW9QrbQU7/j2oRTDp2rNYn7r
TotFXQ3wWDdxyL883oNEB5YHDTnaZzNLXVPX8Do9Cwjb/cInsjbj8bO9zrP61zYC
t1l0PNzid3bgG+xdrZjgndIeLxy+HzCXGkh6AiE+rRiuuE6CsmOZg6g9UhZJZP+n
HheF3OwK9eQhByFdlalB3dq8C1fJ1aLrHZKWBlCIWFVjgwurKkPmd6LP4uzqEl6f
nGith1WDavzEWtEbhLfRZNn77z+Rfl8O9ohzDnGHf+NPu2oM0e9rqTxBOwSpoMkf
Q5Ze0qmr67ktWbmnDeMGmMcsPXew3ZlBq/RW95TMPNjrZKdJ1yB6HDnNLeBFM8Lk
cQeAKnHpX3wOCiUEUIEvXIQSuGWzA/tTdJSBRCGDayk0kjzmDy2w2PZz/9icUXbU
H5oz9jAgVAE57vPdIXkLqfCVWlrLnKpPHvvg2UQpqA7Hp2wKA5TYNiPuvLNzjGtZ
b8mLKvKBYq0gauBWl+qXuqoZ7EQQq4ny/RIy70mPk+3SyVsR9aT8BDj3Lx+v+Gfk
ZCL9tIaVSMTSqTSilvaXAyJjM4zKUaozidYYzSHE+K9hbM7xYL0cABd9kZiPh6RO
yZ0ZfQdyIT7Zagjj0RWz6GzNWUu6kRcR7lEL+AKkB9papBJ9hYHukMZyh0gCk2gu
KoAYyZauJC6gzhTv1Cwus7L59H9Bv/jCj92SJH3leCBH2bgmv4tPhaIByujnzvjS
UnJNozlfybg/tcC0FfywkkgGthOG+apM2jSIKhqd4bs4ivRpJNDWpS5SIrt0XCJu
E4N7VG4umRwCGVel6eqtUR8cIb/d6n0juAOKbv2Zy2Av81JWSYOdLd+Sz6jsIShO
sjJkajFE9ocf1GBH78bNfMo5uDZwVyjUEE1Xkigz/JMxLZ3LaWBNXB22C9Gi+ENz
ZXMSoPnjkuvnkOXAM3CodMSYo+lM7+1x0w+cUwl7vbG7RSg38BxDNFGYMsH9z7n0
BMfQuj4Tz3eSaPPTT2qPigZYbpefLKpJ64XRKbSSVFOUdcHaOWtR533W4y6CIpj0
xFSnz7GX8OkyKjBEGP6D9zSZcT/mSyz2giNsNJhTor/Qa1WZXn236+kUAvLfXLt9
+kKoylM7n5/MybQb7QWgy64UnVyQ90OhJiAU67ZGG/m+JhX6z00amXGj1erYsLXW
+UG0YYeIY8eVAdUaCi/KPQWM1hdQ12diXmPI0wZ0zug24A7+kKvtqXFF+Hi+f/nj
+MSE38JdY5UBkGRBbtoKvzVuafqrppETRhC6zCkyHa6XFqAY0+lfS8XWAiKwNog/
C3ez8Fsl6EaPax2j+sv2F5RzjYQLBNf+OkJx0cFLrHVxjrwPaeXsKWyr31gG6o2h
BmUaMuZY7Y1tfP6Q/w8vonhWzNjBP+lOoBWpt8xY7izQFo++4PaZnnWIdplxre/P
vnRRW0ajIBJgRDgFUtD2zAB9TMVOe3hm1jnw0v0FC5jQ9y04pQ2xFNqtZGnxHrmk
zmbMx5G6A5mzuuYFDUDKEWq6sAT2poQCgl6HESTFkdAKkpxk+wqdubtoQt+r/Vbq
5SDw8lwHb1Dp3N3edEKlXbAzUb/Xqy//EEc1tEuL2qryhO+Vh2I6x0uDbb9hJxdh
LmYiPxUl9XzP+VcvtK3dOmUvviLC6tdXmzwjTGLLXQvwx0+hxuVwQAVkyOYyNJzk
LhMbsYiYrjoBBbk85n6Da9NFFgG+zegd1a/01HSDt9MSaV+BLhbpZYAiBjeA8jDp
qNnqmobAc1eK0W1+27Ub2LYYYjcthBb7u4u0dTwL+YV7CNT/3+OxKaQpb+I5Af/s
ipYG0oafFtsa6r+lrRWnclANpDlLY7TIYoK82MPmdfJEjtbbUqwdMonZDNFB2g3+
dPQEOtuX84rK15OGSmPrGwSLfKNAFHuCO4uWTvQFShrvY1qhqOQz+upcbkqAzjLm
XpMJcpYU5qxYpiLr9kcq+u/hC8qzK62/+jPfD3VbhmnMUts9/J8CwHGcEPJLZIoL
P46Q4+MFbpvG43yon78zof+NawbLRPGddDJnQtfQ3xiYT1y34P5AfJEPVqAeI+rJ
tGb/rd13OB08CnVfmAwGeFNBpH7wGrgb/SvUTo2p7eQxFqoLn/FIM9n6mRakinrN
jsxkuoeIkG3LiJBi9FO6a+sh4UzA3GmIyN2R89pd1/JKzxvhS36zR9muQnvGBw+Q
segjod0lyZfQoh2BKr0CmE1ALHYsQa1UhXicMTWxogv2gPu8PgpuaHKuNHr2G/rp
jQfqKo/1pJgk52f/PmHKjykUEARcHJ2NpeMjR/fP9Cyc+B/pVQtL4WU+cMp7ElCg
GuSuuxd8YHrcsP/tOckPJT6dj0JsIxj08ZG5f60l6zRCEfokxCoq4LE6N56sc3QL
3wkvGMgixEvL+I0CmZ0ZSm6ZmpStn7akSUZ86mYoZ9bQEOZKhaJR1SsQCKWnmITD
hhQ53WDw3u7l9QzC3mxlJ0BNkcRTB0gh0obvYUPkEuad3n2JPC+ePAtkC/i5kujM
5riYjkx4/hAdYKDYMzla4sElApFd2PK6MbBS8cj8zluzhiJeJtNa9OrV+j0gyZuk
pD0XT44qXHS9ENbteJCCsTqRHd25vwgIenCol6OdUTmYFVIPpHJmkH5KmBYc9kbS
GnAt5ZrBxpz/pth/mJ9kkuvD8rsGyGKiNhfIrnTAj0b2FL/EhPQ8aVEAqjqj9RhM
j8QYVmuOeZBERXLE/Xq7tB6RBEHMzu7AKp5I8pZ+2mSG9NFJ/z9FBRro3/ijj1nU
RztM8k1hUNKg/yJTviRcBWQOh9UwdeOvtnZ0ProCS5UA9o9QnOeRLIWH+6nvLOCZ
be1AzsMFqNHZ5lLO7Jc8sJCY13KS3TLlcX0CfYI1sq9TlGZ9EEoz2jgm3DP8pJtI
W72Q1a8VdECUr/iZnQppqQV2XoYlcERyrVjHbQNLrgMTr1nQVxXy2d966G73hAPS
OBkjp7pojDg3Gvz0CTm722QWxA9uZUTaSJRiOoP+CUQlypoZg7yf8+B8JDbbTgFm
mY5pTZMaCvnmgOHuQprUyLxeEIhnwvk0zZlGqFryR2/Cuo0fwEVICImUmhVeWDRg
5EygYgPwjMpBMpertfC8Njw93J4JC4MYUSaZiYZu/kgCchcO+dm+0pMaaxPodSZO
adFBOyS00gKk7ZK/uQ5yYWwJowbliVAwmBsk2U2K6ble1KbcGkFIIgZm2MFcmb9t
vj0NU1choXNSpKQkVMXM9jgKOA30TwzQ6e7WTqp9QQ4=
`protect END_PROTECTED
