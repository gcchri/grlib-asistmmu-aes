`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FGzdw7p2zVg48ay3ZV9axHAn8S383KgkPJJ7TgjOIpHm2FbP8XEJ0Om746+8vM2I
xqWdYlKRmecjoZB/34hsbORPgYW1ruQ3tMaZEPgzmcB6yUZlD27NN8Clc/+pMA1S
aIp0uPy8PZFZiseHJhimMBtjkuxGnL4U4KxD5nfLdKuuT478EVRG7tQHtLKxeoyX
rhx2df3qomyxyHLq9v3QYTpzLPG756W8CutK4aIS+YoSfEqYJBm31yBYxlcGhJaI
LL+41u+8Z4khbHFFCAGFkYEGr4H7hPmFHxWOy2sz68jF6BVENJXBv9UuhGzmKRdJ
YL9O9dzhPhblyxJlKeauXdzvxNwuI/AJItMbW/4E06daIiTYDMrQgbGL+t89wn7/
fj0xqwMbzdukzfWOSdgGWDdJ0p/YZo8L1ELj8FK3jkFHtOFwb8x7zd0pQArip5mA
`protect END_PROTECTED
