`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBLjl5+M9qlZplyWSc2gvQrU6PENS0C6PT+8e/N5GhGy/soPFtXiPWEMyIoI/MX1
XLK8xxPJNRc9u0K0zNI7Suwuy028Xb3Q7GOQIGp/UiRpS/U4EmHzgayIZ22R7q3+
S897KmMprpyZJ8DPJxpRrR0bFhQ8LNrkD9HL6HQ6GgsmiQtram/tdM/bN80kfkjA
MEOr478V9948rz41ms7iisZ5S4YAgG+A1vbkm8vM/BFY45Hv64UPItPdSvg4XiVA
Ku3dNzjN+18+p1JJaw1fWT+BV1gklQsyAqD6CkMxyoJEllm1Wy+dTVNdrpQzEPUu
cIHRaGAd356Bs0vJbjJmNmgWVNqJchw5dlloCyRzRakZrCNZBXOADvVVd9427yfC
bYI3PynkSVWyRAd0bAy0Sr3N0FvhANJeVtxoV2anwxfFn0BfZo1qbdYSgICdgT49
tuhwtPn0SpHSr00BWLTA2b/f+pg0IDBtE2k0zS+LFcDjzkf66s2uY/2QRo7urnBR
mxETOpGY6EUtxf8PZNme39UqgHK85FU/049Z6Fy4HDdpjbRNX5nWCKUspWVCl/s3
0FPVsf+dhR/7rRtFLaP62I6B/ic4VDd4t0l2epJmzBk=
`protect END_PROTECTED
