`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIZyT1kMfCTOaa3To63vUxSEjgwnVjFVpJ9a7ebcXdcl/00fvPXzLtnKSBN1d7Vp
MRxxejr5w9zO48PRcU8FEKd3TQ/f9R0kMy5d+faeeKlJUrBZm2YZsAiWkYGVSMzk
A+mrHhnU8XBz1krfcXxQZ5fLz4whN/UxvQyY3jkMq7Lu6lvD3SgoPpLOAE1tLkty
1OHfc6YUA+dANWXn1PbtRtwHTGJaUrhPcx+y6QMVKGQIQI6HFtQTNGWRD294dJci
vTAuK2uSviD4Xn+5w3slOXi5PjOZ0+aKiZbHLaxRYHzMHuOo62TPsqLwvn3YT0kH
r/KDHxvSLwCz0fcZHnn9nsDZs+4bf1Ggf89kJwMY0R98Hko1cJ/jJeFczn0t1UDK
v3i3mXmc4WJHv8h+TbxaXR6RXjD3f8LxKiypMNZhbQ3yir5USE1/FYrus4xeHaNA
Y8GbQVhAQ/WWkoaWP7I6bA6zu209mRnfLIkLBZSNPwFI5BbGZasvf9crf6S3MJSr
HBCZPF+hmYXKxLnlBLDdrTryD4/JiEC8V5cPf+6LlJvC8NIe+spIuJBrxlvGm3B4
VqqQfhJUB+yrH0LohbaZfdFo6SGsXQyg0rCrsFpMg7ZGiegpOn/pr/x54Z2qsJwv
LmzLcWIFurynnI7/6fawkL7vUYTDJC4zKzulIfV4e2Zb6KSM0RgYgIGNEs0oWJRv
b29H/mN8Asxs+MucWsHpMSGRNTNrNCDUBfWPvB63TH0Z63OJyANbjUdJ5TdIXhCv
PgTJeQI4aP+j3YQL84BhesRNaeotFH08zjDV04KD43GUCPY3UkueKKEaZWOUnukH
fW6Kbra969X1NHTbxCvi18ATZttS8alEpyGTV9lum7KnkIw/EU0uin0fJ40579pP
Z7DjJaM8YAtSz9AimaxFEg==
`protect END_PROTECTED
