`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEz0wS1bA9FcSRjZ7MSpowVBMhv6WACosQ9WkAI4Bv4j2dnooshBPvuoaTkLktKl
XjN/YDvokyFX436ijPF9YHWCC87kanZW94OsT6aS/cWiWW0ZiANoFFWFwueVZHbw
B6eaJB3MEnycqyRsOcyiGJxRcje4yBWTN4dYYIUXim1u1PE2kvhLKaj18+PzvL9T
dzrtSGzHnx5Mm8cJBuWutnF3nNemJkwIb8bATLRY0YGQcFBDtGort74i0cLuboVB
wj9wJnAaGtk5WeikeYczZTxhqAKiX92cwieiVsgkohZDbSLinHGRWr//lhTNloks
i5gI9fZVslIiYv24ksht8RBYv4R45cxgvQTvLD34sUSUSxjX8Me2HXYe0MZu4fVT
RsWRoOhvS6XDsKtv5PheZQQOW0BU01ZIDRxBCle2WS8=
`protect END_PROTECTED
