`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MYyGJC5wF74T+FNU/Ym6/geXIQl0/BFke+j1+WZoffQaQFA5tIaPt7sT7qAfiXb
Umx/EHJxT02GtdICPr4+KddtSzcYoneVBz2OOAI/P19bHBJd/TA74SYhrXZUUE+A
pdxaDrtW6ThysQZHq+zmn1px71pcHcJyQcdqciAjsEmCakM1gqOy11csBBRs6JJB
3L4mVjGvcJvePA42DW3iUO26yJyVVgVg9vZxywaN59RDwyVrhRWGOZb/A8ZVuDBB
kqtMe+mNctWX78PjAYaPhcEf5vEFF9Syq6HYyWnJhPNjfZV1KQYg6hjOOrRw5gQQ
WCbHJQq9uxDM7cC6edmlisPSyr1MtfAWxSRBPX2uKF9b2JWMI/7UF4VS/YQrwi0y
5xryiUoJlBHU1LilWCOdxz00Ba2KA87SsBWaJ2Payy7rdA8hBL7VktroukLYBKhx
p9UplwWIEhwtqnJTZgvYeUlNtBjtIRy9novsqZIZrqyf408iYtt/3KqNl5TMk5yp
zzF18KYzfqRD0ik70rQeWX9E9AuTtAxm+WI22wWA0nc17Hrxpi4Ue8T8GXG1o/6o
8+Gy0kGN51f23aQXEh4x2+Bbvmb5twZTOuV0F7a/dyV45f/reGlaz3wyHmMVPsJb
oSJQ0cgchPCSzYVjMf8VQ+AnvKujrWfw+irBjderulvgOwZoXqLyA2ejEBNg/amJ
hN7BjRIa8LgU+0hpcs7WJWFAOo+8IC+nXxOD9EjWZlBYLjlHhoHu1ki+Mx5uquce
FLS/fuF7Vad1jkfGzLclGiS5MbOINYXhwJ1zvq0U6PEqdiA/+oLxWTDZRnKcwDBU
1XVHAdS0Mz3JpCSNL8cmEaCoHgnAri/O2T1ie6aGrsuxRY1YdYXcBm8XcTaCJPPr
pf9gPx+z3xfHJyAeejRzQHB5mm1wBvxhGcQtlvD0dzByd1Tb26LgcUNwYfcmztCI
`protect END_PROTECTED
