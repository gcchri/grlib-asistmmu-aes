`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uhCqfE+ulu4kdx25ObH3Aub0T8GHkMwTaQUymZ9VYnOQLWELRYPfx0007WyQa6xZ
g0TpcQxYCpBCQubGvrGGW/VifY+o9ZexKG5yac0xzIg7uMc2w670hVsF4Wgb8GTN
U7W5XNP5BUdhJQbGRbXsyBAAxDSZdPt8fot6U8TBM9lLJOrW6jAZ8zCDU7sneSvR
91Go81r4Lek8Te3ux+t5G+R/Lo2VHV7AANcU8WUzsl5OlF0LwsPJKWKT/4NHghm1
YWblInZSik2U3GfBHy67xLZFu/UbwsYKgP//5cOm9Ee7vEmBsxsAw85Gjqne/xeJ
Z3KaP3yzuvxfuDkBanty0+eEmt5zPjTO2SUnAOBatVtYnGjwiZfoVelda0nHKK9x
5H3EUZGPunq+Dup3QBjMzYUX4usYLhzLqYLg9Z3aMGL42EHqRb6vOyeqEuuxLviA
55E2ZMMWpqPUrGHFDArHkExE1PxektdGRPmmyJ75ORs6FX3DgFYFodE9w9+Xspmz
gJOcOsAi03p4OHT7W/0CE8hDlXR8ImKvlLQVumjywZV5zxKypx205sf0p/V6+uVZ
m6OrorUQHQ0f29k+yhEIIQnYTc4Q0FenTACoL+uifiB6r7a9plOk6MFOlndamhIq
KauptKkHCkeXUrODm+CCNauRgw2PnYFVy7fiaDUnxFluurIs/Xxmv0NWSwjWns2P
`protect END_PROTECTED
