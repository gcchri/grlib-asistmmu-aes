`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JFeMBmi/c3ERD+Fj1axGg2D7x94u10kv1+2rVgg6Z0CfRlfIbS1LvRoOaG/z0kkb
9QE3eJyHCK00FodxnNUnUlbuXnneJlH1Hmg4xgZ026lpuzf3lGTQmMmG+ajoucX/
DbziE3v5QtvrT6cG9qcMD5VXmqF0l+obsdtcj31QkeZgA3gF4zRqsI+BMCIJ0OSR
gMHXhcJxHlORu2zr2pc5yeDwJnzj0q96Xc/IP4638QVRcYa0K7UxmOQx5Mop2/x4
j2lybF9Vv7urM6sezWb8r5iQuTPf5OM5lmOiK7AYBE2fbfOR16SMUWXtfIDcsf+p
SFUUuqWxHwsk3gGtQ08Q0GqDi+GXR+fLUOAccGvU6hDJkHD95WA6rYcBgGjHNnF1
Fw0mH0aHfzp96f91p+l1Enar6ruIXGYxO9EE7YilDx6dLr8SznYYkGU4Znx+hSdB
H2SWKwD21jrPZI/UGCmVYP92zDdOsO/YMO2HguhAiQTaoywp/f9WqSWjC0rxTAmw
UloKyM/FfHrqYoLLwvIDB8kbawPL7dfow7Q4WQTGHIC5+UqBwrKterpwvTZ06NbA
Bat8ubcFMOUNZr2cJhWEEyljPiAY79qEMKCpNvWgL11XVsnWSN4cBye0dlPexkQa
2U8+0/IPV/j8xW2B0yoZQgsasdMt8HFG6/t78+xXI58lbeaOSyyT4x96gs4Wryg8
vetD5ATsWJEMlahvdDsRXKQPcXttVTWGSBmm+1KwZ7WKlPSdw4bOvxgUyrU/tWt5
MWRaUA3UlpipYmcNS3RinKQ5FIFJ3mgcfGjFk+Bz+zekvV1ktpERjl2pQEwPVuEZ
Ye2uAeZnNgjQiZOzbgbsJJs5n/6zCPj32kYgv7aepoLiYjYW7xEOARV+De3N4qPS
mHdg4kZVPCUA2E2eZQCGp6SsZiHD3gBDVsytZFX3lxk=
`protect END_PROTECTED
