`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7VYfoc/ZMNYdbE6Qd2TEOv0fjdT1bqvB5mHhkk1OEE+SNTlA17Nw/ldLJ+4FpLT
34qzEATRU+qYavV2h6yWJ1cOEetPD4HTwnnExDno6qqtitu8pK5miJe69f04jpXu
QpgdA005ZV4Uimn7+Li73iv1whTdOya7ODL49J0QigiJhRgbgLfKABAzGtV1wi2s
RS9aJAfUq6pO1B2Q9LquMDBZb6hIWNOE+lVinoxWHzBUTATTcMngj6yh1U97lind
mkVMiwN6VOcxf09weFm6TxcY1n3tkJI4uMEpog4I17Ar3kYztEL0+uZmrURAfU2v
CvqGWKKAkVJdTKMha2/R6Nr1G8N3mrdpY7QfnzNSfLGNQB4JdNZlDPEMRMMdrOaM
ZZ60ALEEwRopueXFLLJxARA6jV2EbzImkOgp9saeRNLZvCMqLHWoji2beodLFVGn
p2AqnzJHvx+HYf1uVTtEqjSGsGALcPR4Z9XLMhjDeMVvoK87Jp2FUkqvUqnpOgcb
oyi42M3ri0fRpB2S8R4jJnfdZAVf1VE6eAXVk8+fn92QPXZ3ggEeSSK/7XsPokTd
0Unc4g6Gw3kZWUziUB5E1KwrEXwR5QbjVrJkqzSzVRU=
`protect END_PROTECTED
