`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRkzObLuKaKS1Ao3KuhOT1F9Z5tn6XhpnUejAJ1wvQ1Lj/KOEHQu/5JQ5FPpHj59
CyH54fY2/91p9wydh3sOMSEMML8FxUAy+2ZGKdjmne+1kD/EeaIppI0erpVTb5Jx
s4bpTpsffiC6d8pf4Y5YfJHThh+m2sjTrtYEbTw9GmmOPCRyralteR4hJCQdNfLT
6sBvEzkZKbMQcMauedJaFaCBMtYjmb07Y98Uz/pCgasyQyV2clGq0wFP/uoVbD1x
44Kp+zCgPA5t6n6B3bF7UqML2xMcpR+5DPbrWI2THAk3e4QSzN1ki0AsCs9G4ABj
WKhxfw7Nl9IgzElDwAvlkRhzHdD46I0jnaFvahPauQQGR/86MWhYl9TRggt2RNO2
YtXYSceCSSG/OQa1Xx6auu4akX6SlyESHTMecNwYgUvL+HjqFXnf3fHIqGFY2KuX
kVTmZqdK1fP2VwM/LROWWH+mXoSHpgNNL1A2L4FP0dmk+darwC04BsX4zDlxkk8+
wldJS4mvYUguR1yIG4wHHNPwuCuQgQpU5KR6eA9RnW70RrqbmysJ2ElE7JQQNOhz
`protect END_PROTECTED
