`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDJedrR7y1epQHaDRWVrwkgH7dz74YX+a60BGamK/t0A8GctKZgYNGWNnGlUHBAE
g3wHOkYHsFcY8fRqXOeetKtIDpjF/Tw4X5tYHFVJsGhJBWOeSsE8qNECMBqduZA+
DvhVfdonu3Ar1W6NVSNt+oMwTxF4YlFaxBQcujV9GlGNdNyuvgIonA54GKYhTMkn
ZHdXUoEmFi9nYI+zVq8r4xd+UFuQDPUPzMMVAXfe9lrna9BxW5arBJWInksmVkiV
yQsOSI33y4ek0QwP2y4aAJuyPmxSIQ6IW/E+zOZBHOccuFBwBxHh4rSLLGxrgMbq
CJIq5LdQseCrGlaUg9JDGZ0lMzIxg5mWgYd5wAXRjlrqQZyz+aJdnFjvSjsW9Mnl
YVzD6veJVlVdtK57pe7b+qLv8MV8bFCkUy47UtUjTTtUPJ7I6DVa7tC9HEfzwShe
YhpDEhh3OKvksFo/s6RowUU9FGR+KxYkjlkgh/bmRzWbRZUP0VFb7sPDLC5l8cb6
B2+75GyPdpAMAHh6joSANyo1+jIGTvkuypJmMzhteXE=
`protect END_PROTECTED
