`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DX69BYu9sKwieX/GdEM0Anfi6PkmKJUaoXDB67uji6Km7Vo13nAOyf7vaqdmw3nA
pyRg7/zghEAmSifz4Jzlomxqm3xlAEOI00b2Z7bBCB7o04WGEKbIAK0rmeRVJSbk
T8FLIlvAFl3ghPoEZr8NSuFXkOqxKZmtMXzz6NDANLcgWQDPSB/LCIGeY/Fr6T8g
0eMlMqbR3tbYjLYos418IzvLLjCd6OqXp7O3D3/FQsXEvnUIVaP3Yl2KApwUqaXd
wuUrzTl5hL5oU99WGwsTHa3Sv9gCy9SZ2w9yib817vscyQE8wv5ocXW2htzfTOjY
8aV9/00MIp9Kt3j/mTzeKvaykpNKm1zBkROCIPMGzzDfuzrKlYi/weRsRT0Fhet8
zk7AzSP1JROSAMDd/XcSDggyWApIycp4MA3QQi2hf5uWGwaDjtJqnC/LNA0k2bUj
M5SYjFS2G+5kP8/orMPh/ANrxn6kr0KPtFbQhZtumT8nkeuEwBcyHLTr5mbs2net
hcfpWgFKRGKB1l6nyrV+9irdpRzdOiTehT4/ls4vi710Ygg+hSPIPmc4XWqTdz6V
5esWQxcrLg2uzacKk9LV3t3aRaENMc1fDSt9eSXm+vhva1j6onoym5hZ3adGb2U9
Df/p7YBoiwTGU2yFe9cvP2lx85C7YZ3yoWSDdkbWBlVP6QDjgwX+p875cBGKYXOl
HAwd/UZ56kNkNBxGaf4Ku3FJEvsgjspiDjaO4Rc19aE6zGHgUWQtilBZm8sjv4g4
JkpdYVPqvhljTuwjmS8mtQtkSKEMCBDLFfgZ21xBQSj7O41l+3L8bonex/dEN3QT
QFvrvasvDzFlHe5gaElWqA==
`protect END_PROTECTED
