`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dETrlZSLQKpqiZ67PYULqOTjEORnkwYod01OgAXuegTQZlOEm338Bn0kaexbprD7
0E/uZF1Q/zw6h74ekx/7n37kM8O+x8WbKNdw09mUePvDGw93x80FCYAUMILJYEPy
roWvdIstvOjlKSlLTSOL4Z9yIlSvQMwpSUWIQA6t3jiaaTy4JhADAodwQDcOwf3t
02tepwALW5K9TnGUTx4dgAmcj5q7Bndt6Kb+AzBXAfB0vHLgfKHwjWIyyU39gOrU
ADvETIuTq/oTa/Xv/+gjb9aVL23iD95MHB36O+Rfbrdqki9A7jjISJllDQng9MRW
C0oGN4IycUCTqtj1M31jPJRDjj5IzYPhT6nD0MkJ7jvenAPv04tX8IWHlG+n7KXL
BO9InwJ3xJgvjCdMy+iVe4S+0B2pHR8o85KBETLDnc+UqJoE7+b6SrjtR3Sy1uGE
ZtjO8nBk4TMdZbLFDSgtzkTwyiDgBEdlGb1a9BtpxPFAzEy6yRLplcFZU6OOraW5
ET1vKptM7uuAGPJKKnu8QJpkZdoHksQbdyVlEOzVQAXXAlbD+QXEMIK0eiF4QBJb
Ay4eX05nfXlw4QEwaKPYKjaHOgn9oC023P4RwZfOQKe8aW9cZns6wbFgHUtxzpdH
`protect END_PROTECTED
