`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wBqZ1GiRdO4lTWzQoXBic2NyatP4wvDbWRXigfB49Ck3Gd7LPuco48VCkH/tA3X9
hxKBlvBUckHkNm7IgqsGIPPLuyicBG8d9sMMM4wojF01wTtyXZtkTsME6meHuJr2
codhxpvMYX5R145+PoUyacx2SMsnAC+ntuVQJKS83vUc3x0WpAMWXkAocXub8YEC
/xvJ93FE9qsZ3fZd/NUoArNhKa+eM6DwIVTOOIg4g01Xx6MVYZKYX6duTMR3A6ri
ICAJAziScfDsHRyrJ7VENv4dDhq77bSlVTa9JsacGmrL65noPU0sA7KqA5tIjP/U
X8PGkWmjuXG0TrMLkKb412Ykrd7NQ9z5mKTWXCEI+WRAtJwNwMPp/8t+tw8i2sgD
lQX8as/7JGLHaVDhLZ6zJor1AFByWMt/QfPouXRPuP4=
`protect END_PROTECTED
