`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6jilJH7s3VtsS5Hg7Vns20iFib1gROSCVY9OcXNXstfN+4iA7YFw8SwOvGTLMvbZ
R/uW72NKtLk2M+jxWLsqeCQU9qPFLTZ5BKLBvUWoIIgrhRWeTxu0CNYcFpsKa70Z
xTQObuwpy6l8hA+F+UIgc7b4AhyZt0WG4FcgL+A+iH1X1Rv6rMv4yA7LCrLluNal
I8knqQ4T87XAY4Tijk2wKCvjYOHYv2WJgWdUNpFhhPuhIMh9QX947sjQvovxqL6f
qlojhsjn8clwQeX+9YFGoEJIxiVYXYUEOEo3QTIGLPXu+uTZkBGZlxgywFhIkQfb
oTmfPMBK0aQjRJrWk8MbefJwK4ILTY+mYlMd87Uw5Znbs8ZXQUGExR9CnnQH2use
FARd6EDayVlLgk6wFUzQPyhZh2kgLmNGEoW3LAg3voeAOH5uJhb0STO6RoL8MYoc
ayoDT1tpHQWYVYeA8yEbB3O0FwTuSNkxof7ADo2SGezuJlUagsNSZNsby7q36yDT
Q2H8yUsqyXCLLxcPp/wQyNlMMLTYUcgtTXIupt5zxIE=
`protect END_PROTECTED
