`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wU9LzKZDVbVvtF9bWDR8VwDKv+/h7IQughImRtGC0GhNxSKrKIhBOheqoowEfqGh
vd8FECH4P0h3GZSF27K/9CBT1f++cR0YHLh2f2AqYF8qpFP8EFdcrxgUiknKB7Rd
VNx5hbdKhNICzN3ua3DwZp15RDP4bVUAOqHOidEEkPkapiP44UQfUOEyfWvwUymd
zyBls7sJ4G+XxiWo/olHHjrkha5m3O8342y+uY7r7W/QVARE3+1sqK6qLR9KQuoI
hRHvKDSYiHDY0i6HL944iHZk3ZUqV4lTKIiWnGvp4wsJOUsaWiYb8nOZr/s4RLep
`protect END_PROTECTED
