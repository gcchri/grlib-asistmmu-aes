`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFy545b7AOXtbSPBjuQD6vA8rufXg0waXofTczkl7R8flwDRfP5WFbB8cOvjtzVh
WaZCnYJKaTY8WEW2ip5FpMIn410GtbdlpcJWTPYW9O/KcaOa3iEUo5je+Y0/y5v6
/HAtVvsQ3D58ryvvOm3dxQgsFuubCaU/1y+Zaoy+1QNQS4iom6ZOyi8Q2cokChMv
4jcrQFzMhIRn9S28cg1tNohtprpKV1aHyZ0bDAgx77xOTgV7Y7mHUG1NYnAnsekj
ubwrmLzf/kpgbkupFk6iVIacPmEu9aLeGVkgF9kixMIeB02UL+3CtMugj6l/M07V
H/pieWnOgprfRM97y+9m1zwlw9HrTit5cGxdAUfvKUhEgX99eeWgaAWD3zu8dZS6
ZFSxAjvgiPq42YB2P7kHnL9C4bwN5wkdldCNlLTqoc0LHV0I8Eume/3K2C8Ch+rW
Z1ZWHnIQdePLDl5xbFgwmwDaJNJZNTSBrqs960HgeNLDIuuui8QwkeF/XTnbO2KC
9xyKyjC6gsuQoK1sAIm2ohxXmNES6ie/HN9jlpPkaqWAehpXANQbXuX/ypWfF/C+
`protect END_PROTECTED
