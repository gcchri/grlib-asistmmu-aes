`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hnwo5OVxivm9WD1Sd9YFm/ZMnmo7zGzZp0+j2FoJuICcVV4dwse0B8GmayXUr/mg
QgPnwJSn2CwK/XGaHzksxSwmcvDQOZRkflwODjEz9FG5hEykYgN89/Se9NyoNlaA
JuV8GlqYrkeCJDu4pEBktTyt+B8i3h3KkZEChkbVF3274O0JFEx1CpA6VPMmqEN7
gE/IivvndPe5JO5CJlV1HnlepxmMLzb3m/LXqzvxg79L+DfXpKiGs4M9Mc2mrPmL
03x+gg8dz7BMFgu8XZTR3wAJdbf6FTNbOeGfb8flDiIEYalx+xsT1v70farJshwV
/E1uU46Va6BgsW68161P5NxfWPo3/M5y7pICCAVTNBrk0uGSVw9SrIjgam9/x82b
30/zGFEZJm3Dez3+d/OMqU5fRtyoexZ53L9dSb8rMBZb9KNnGDpUinjHWKpNdi8H
q6QOntdW123mJGcRlQo7e1yOMEOVB7ISN3iK9Jo0vycamGSuWwa/jeoa2IO3elQa
`protect END_PROTECTED
