`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tICx3gdFlwFeLWmdzjGOfDNknYNH8FpJPkLqGo6/8NneS2fL3j89/lf7jYYFf8mc
3wAOTyNzUxB58gTJ4TcgUaUKSXUZj5FbXt2c2m8kDNSrSM3/fZ5gYM/XA5v49HEn
LwMXEdirt1GXbS/Ot7NONHGLZAzqxxcRirhRgEJ/MsWuKjgZjJsEscHQVzSMlmwe
hnP0RqOP+KHRBiFppCq2wicLPBqeDuwfyzo071nZ19631ReLB+PumG5EbA6O9LGo
ap5b3TFUfih2LEFUbw/hecF6KtODSUDHBaAfO10W8saq11CKbgnefiCHHQNvo4tH
YzMeT+TahIv1wJAo2iBqWjOLiAxa/34EgmWPfA3+dORIYsDFu1uLo+qqZm2wvl4O
B9YMGSllvbHfZh8xvNK+yyN8jg+ECXZ65FLEbTrFJhKDPFhDkTa49yA4GJsmG8nL
NnFXElcTYmgZbBoZsc0JWSp3tVIkyI5sliO0xIDPg/BR7fYsP7Jp2vvBDXtHoTI8
syfqq/HV3SF6NUJEQ6XbVBh4Z7msm59/a24w++4ggWvCK+a03mMZLXxFs8qTDPn/
KTOPs1b5zN6Yi9CWNKUYX2B91Ki1f8Vrutz0D85ZWTFqiLZoAIC1AcnlESWWFxAO
21jdC7djt0OUBsJUDI5Av1xJbArJiE725/TROiUET4isWJQipk91seeAcPVOUrQo
DMTqppiIz+5B7Dms2oC5DzMGzW/BYndSBm0vm2lGOi5Ke3vrY7UvV05TieGpB+Or
YV0HNiGo1Rr8Rp2pJ9SJt+VneDywuQZBiO5hBMX2an8WeTwTUIYcdc8aDp5Q/p+W
v18ZrkwkNIt1Y+QZi429YQ8Dfvm8u0xzibmaA1sE6xi5pTJMNDBXWsVjIXn6HUjZ
t8YeFPffRIFH7J2QzqXo5BSZF/cY0qwmyO4nUvyOlmDQmSo2+HWFKMYBc5gMyy1W
c73V7rJzSCc8YpMmWcmc7ISnicGI8xGHxU8pZ9plO9rpQa7/BmFQBOHyrn4mGyi+
`protect END_PROTECTED
