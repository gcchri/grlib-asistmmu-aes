`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EVT6tqpdYWe0cpgpCy/c6hLvgZRz0vMTtl1xKdR6OifA88J/5cQdYl0zCgLIjgIW
0jfhQzLxYtpNfQup3wFB8KgypqGVUubPFxzmafQsQK0Uuv2zBYsIPdIMKKiyoXmx
sB01YnJMjdoqfYOI5bSW4vYjxQinNnJWbB6y5vTEf8v+xeLdoAJGSUYXcc/DMcEt
x0NhrwDN6edK1v3MhoaT+TeCzI6grr8MkGSm1NUgFzA/wGMpe6onwKIvRTGrfAmk
P5zYgM5mJvKN0RbCWqOcDGOlG9SP0jSnpNw5iArZjvpfoT2fHS9e+o4BJ1hVlY4/
/LkzuKq3dN03vh6Xgpi8GHHQNRSw0pEQVR7ussStYClTyUBbsQrq0STefSZ6hxsl
nDaCCT4QoP5PKSHrjEfptPZ6kEwcl6ZzTTTUlhcFm5F48A9hsJO+eZY657vvg3pF
5zvd5pXLKTEefkTGobXHS0BsZIOx+FsVno3pcvZ8Ew0TC9KY19fQd+M/ByO37fSM
86ESZE++eYNSO3U/5BbWBufTmOtICSiTGnaZl9zObHAXz+C3OxW4jfsrGxFZmOdZ
5tdRwtndMvjs/GgXSo3wPyPFzk+Ot+v5QoyNbU3V38YKa5U/93exQI9kDSAFi/G9
Q8g523fSXacGTHKdMYjrfjcLWPXh7vfn36ltOBHvKQQcF6gYcSXqZht8fZrOq5QQ
F7C+1RTP8FDjbojxaNBj3lK/XAo5vq84UbG81Fy2kXBAhYk2JP+uv2lZqP8K+1OQ
x0a5dsqTBBIGCtTpxbXVGmC6cSFCTfAAjD4+GjoLPeIqHNViwp2BWiLk3NtL+0ZY
fqYthjm9LDaATeuiB+X3WZOSU23U208Wi/Xbq0EZAnVXFncIt8Rmfkmh5yc2X1pH
VHZydh03zq2y7uA1l6GdGtucg8/sWCA7es1qBPM4qTVOL31N27Qu2V5+/84jobaZ
2Xo0STO9VdFC5qozkW98RCkNyZ1OkZ4v3GvmTw9CoQ6+FMpgtL2gHzAWGStqi3VA
K41R370+cSUuJ/IJSMauNVDUZr2VRP6FYTTQvpsi8sZf7GYL/TxodFBkA3NbpSUJ
XJC2Fz/NMfWYFy+KjBd1c44N7il+DyejffqLPtmK9Z0m8Lvr4M6evmgPjHO/NeIo
t7clfKqWO7gWCPnrTKuT+GgTyieNZzY4Lhn67RMmo5tNLMZVH1ZMHb0y09xjSTeM
BuEmEf9IL+54NrPQyCFkPnfLJ8eFtMs0ZglxUFl+QR23OL6ZV5KrGsEYZCUyAS6x
B5ey/T0AFkCOdkADnD1lmjcPv0JKIQIvsCTFKkZTVpRuWSlwkNDr46qCwnTa8VTo
x5RQGhCqxYHDvF+aaaqnGCqIrfnmSkZoEeL0/g8V8YURWGsmbSuri31SZw3DMPbK
ZHezGHxFQJfCHDDVc99QX5erCAEOf/PA+5sgtsbwwVtijzM//d7Zt7HX/kQcwYr7
xUuReJos7PXH4C5uacc1EH5omWp/PDZfAn7hSMdGQOy1coJYvJzLJM5fvRXdPrxu
opfyfHLk65u1YSVQg5MZTwyPaUjf5cyaUw5H671O5vhlSKENZfkE+AJ58JPc8ZrJ
fME58Podg5OTAee9wicDEhA6O2SJtTD8J6cQwqrpXI9gxHc+5ngbReED0mfElA1M
KzQz2HUyATkqrk1dei4cyThkZ/4vXXZmjGjHjrVdtreGjq2Qkd8QZL5N0TRam/qx
8+LpAxgANkpk0zlVAnrE5SIL9LiDE0yc/peWSwpCzaQvpKc0YuzAhZG6CAT7+KaE
YOcgVr92DD6dmir3zz8O7s3lVsKI2qApgPAI9tsEPt2Inj0e9jELeIsc9lQT7hXL
mhx/Bjx8QvMRV86GKRQrXPWVx+30CXGi8jgSo2LCoG4OlCqqyp6eu3+rucGE27bU
cecKsoWjhkNzGTLjkHJj7idbIn5IkzxP+TOonHu/sNfMZ8V6eWH6rY3TrkETc4bi
KkYfycsmbGQHqSSFjp+QXmPRykq/f0Sy+o1PdluQEn4Fdccqo5eJQFfUVhwnILcw
lb1aKlKInOnkfxvAePXDaTss2nv1vZlGCe9FDKOqGCVbJ9sJCQWo8EX+o2Fm9OzY
a4ADkcrFVtolDa76R1jk8P3kTFDD8MBIubsBDvQBynxNWC735CcOAHjpRLPMnOt3
Od32eENwwS2fngfL29q/DgLfJzqe0XwuFYph79VS11RfLbU2YSs+IxswlhpEv1Mg
G4TGPNfC3taDMqUz1nbOEzUQCrvXqdPRf9O380SsRU2y9U9Jjk6778TNwNDyQi5L
kZ9M1hiTME3rXWHkfObsEsu85OzSpyK5DH5L95mYsLUYMN7GaXwenkNlVtCRRvD+
mfUNIM6UDXE5yjV2ZKnvbVv2vU59b5XGDs/jV4PnnAdMJgRQMyz+4hVS25b96nXr
NJqBG+9Il4T1GLePlDuv2ka++JZUgbL2+tkItfw64Y2Iqs7NoxaSjzo1pgkWKhID
3RYSpSD7MuGv6mCrY4Yf/IICeWq+sMAWpvC+4ZV94rRwExMN3dDx5jZAhkYVBdk2
MrKYwFYBTqd8UjERmMk446QnizVzkHA/qUeL8hdt4sH7LqzNBfwReUR7sK8zvJst
ONtDW9yGq78qIPpCtT7+0pFJeK3ewfNRYLdYN766dgrPy0Zw2SwHCu+PS6s/EV9z
8fYh9k3dx6jURPzDy2fmyIvi5GSqH61/73ElIUVW5fS+b2EK0LKcxpkpNXtc5ftd
hmcIou7MG2XkbKq0eKrS0B+09/2RbQmDalB/VDex2iNVpfyiBnN+9yCTQqlvBV7D
sW8yWIrq7y/SY4zAB/haBvJxKLdvw0b/sFVXBAhL/GZGchL9WPF1NOiXdrD4DEfG
TkCyFK8v5aqdjsPP7FbfyGH+FhTfGyKfrs9Z+MOL386/9+959K0BzHGfHxjsuVuH
gMZew/yyzwG4jJorQCZkJwpl/4Oxtaq7bJ2ejKER15/3yLw5P7248BczC2Zs9eI9
hXyZkiznv7CaNUguruhyaUMYusKwJczz+N8ezJFQJME1YdJqrphqyEE6puojW2df
l2L79Rr776I8XX5PIqGuZfARCptHECKpbIomPKmeptpzu2uLIZ2p3cBC9Upuzt7/
MrfKo9LS7qz5rVGvbuNE0y8xZJpv+fkQv+dCrgrRA6KWEHKiqamDvzUsYBmlO4f9
V9d6LQSgL5H7sSrN53qZBZL50w/AxMLNIXz8DCoTnydyTPN62rgqRFgn6niLnb5t
HfUM9NGoI6ZN8uV3RUhDGgWzkVlHI5oGfLvFFir+yfPAjIfpiUD3Lp6+sCc8lBtz
qp4CJx/hccG5ogWqTDndOKzznQb0W91v9C6rAKJkcGs=
`protect END_PROTECTED
