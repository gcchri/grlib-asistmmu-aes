`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sHcOxFYBhrR4mK2quwQKd2XLXq2pNWj5MDV1d5qxZUTJvVptle5XAoog1KeBFbGR
NN7GCkn9otMlyLw+5+hKmErhvhU2nNALINahYmpFGZ1zB6unyMO625+2oAdDlCCL
KV16UZx7C9UaRPn7sK4g4DNLEnLMfvAEb1iLmsNiX0/ChVnuLdIULuP5QCvI0xlN
9XdJjrRH0eCh4KdQzc4pLqmEsYUReUxhEoonMx+XzINqjumXuB5tlQfa5xUfBCRW
v4Y2eMOYqolybT/Te4A0QVC301wuzGaJ2ubLsrjQ4r43rM6WyimHSnx78KnNrF/j
QlFpqwsYioTg0F7yz865DhfvUmPxu1iUYCVxnoZKj+vBGhTNfO88FdilCfap72A2
49uroQr5rEHnDrTK+3fFGKUvXzxhX4dlzPGsfNV11f8=
`protect END_PROTECTED
