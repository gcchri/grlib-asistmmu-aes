`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iHI75SrzkAAxMedlv/nlR2XQydVAYBFpycM0lHri+q0I/fDqSByGRJUJNMtEzsjY
w0W6LHAWxS1iEN6GfrzLRinEtY+Pcm41R0Rd7gUCIl0udg+y/pm3dzH/zjjMKBAS
RFJWCMhQx4wn9UhDWFKn/d6XbqOjk4qCsdz9f155JrY2SSJ5raRAQ4YFPFfC7s7d
npdPZj9b3MQG5c/Rnm7h5U4hEERWezadEdYyuumxHeP43JZSqD+LGU+foFJzhize
WaS1ImpSlIuK/PauKh7weAV4vpBwRC/VTk64Yd2SmXSQ1bxKbdMI/B3Ne38HEjxQ
IH3gZuUcYJ9ksn1v1moSKae4nLxe+GOuSYD9NZrsKMLaaez2ulpqHxTopWlaTV7s
qQom21yv3sv43IOck2SvI+3O8T/g4AAmqPNFILBrFHJQr2BddKZJMomPkyWl2+AM
MNvQ+sH5MXOECZLGebGnx6JVsAtPmEBOtfpv9rNW3L/puBptXBQIuVjGCgcMylyc
Zt0HPBUq6QKy6ia7w3SwyIo6sueq0+J4163eezcUDWP64xVhsCdDPH0XjzCcf9s6
e2gLgMxIPGZz79VqofMSXE1lrRabRebzFeBrtWu6aEuEfDeP6Xsd+xQDxcON7mFA
4/K5IojbET74x3bl2/awAN1MIXcjIqLJ4uJ/vGnVm61ePQCy5q2BZMjnmiDXreD1
ffcyAJR4eUMN1hihHMi2mpoLAwSGpbTtuNr97OqcsYHwgOLCtzUkL0gSuLWwXcNM
XIqtVadDbGewNY3SsmEZ5us8tuz3LRgE4Ma0g/l3a1DPfnsL2X6LSkelBTi29CdJ
yL4PIZPNbjNnTWSV0xanNjboThigoeg8pQpZZO7m/01gePSeKSdmSEcAKMcU9X93
kZKXw8X3QIuD0x50VaDH4yQU8Qt8wMrskC1CjBmCIf3kHU+88sQurtY+YjyrVFkQ
//gn6/dkq5RGNo4gflVCfvUPW1JQMPDpCXImBflIPJxGZ6HiotRpsseyYyeqonk2
4zqpDQHuHgF8G7MOs/3wusK1qAFoAV1wxIfP4MnVXckDwYYxFAC42Ler7W9fEgT4
FyN/JCzCY6GUyuOQsXzzKILDxBkJak5wNFolYxrEX/NZFNTA243VvyQz/P8DcLRw
bOHD6FB/qSsm9MBkXmHSncQlLvJFtWjCMG/kbtbXc2Iq8bNw7Qw1gQBTiKGpEF5d
OIdc7Ayh0bdbW91+AJaGuE/I/V7Mncu0RfEuCP2HQExsPVrsY9FEUYdA+c1IjBA9
6i772LFbFHJt8EWZ9WIia7Apu//eV2SRocI36DcaF6SyB/IzIABuIjFw5hPGJDCA
kxhRK33WTinRVvMBXeO55Nids+71jbCphSNUXFEgVylf5Gr0jEEW9nwPsmsTOTD2
jQgwj7ciwnTpNoMOsuwokO2yLWVO32fr99e9osOfERyaSLbkZYXsbNzwJdZEFOll
wCTAUr6N4yN+CvTrdfTbAY03woq6QdHvDzuvHcrQDzOIFj7WD9D18Ua9QLJjl857
tqlXijDPX3hvldFdArBiISYfurZd3n40VROm7eV5Hv7cQVTDWIPROE3XpdqI99zJ
sg1PhM6fLSa+f93+2pGOwWTHEle3/1wOkvgA7KXWhxBDwzv0EpihedkFUHM0nXQW
ECSlkE7sqDahugMk77QWUGYYBU3zrmJTpITZRZI2Usuq0mwu8y40jZ9aRPCa3Mp7
0LPL1kz16x+ZoFm7cRPrRvOI42mYrbV+33rO9L4XI+3G22MGOZw6we2IbAakkVqS
3ESYQTp09pDJxxDulEcryVXMkgPGteQyOTkzNnUcfQZpDVo81nxserCPF9yqmn64
lIGQRsCfqB+EB3MevThZMRhsv1ZDqyqrvRUzzWD5rOy0gyx+OKPlFOdclh3H+SoF
/NF9GID8DAcG7nvj95SVzBHQVXajNmO+8zphF53MsFx1oScwcEoTe2R2Ta786SYH
xlxWdvytCtNTx0Bw+avKS6Fjp12qhlFwcXZly4qGbVA7O3n6oufdSIy0qtrrXp/I
jOTo61m3YA65Hzz8Bvt/Pn+QhDWvMK7HpmWNhzBRQP8RvBBdnIXgFbEccZQnuruP
HUi7NGjmuFGIuWnXzLb2dAC58AGJsvMqs/Wof8zpmvZ4j0L4KEw2EQWFFJ807Wy9
o6tpcCR4gzAhu4PRF0kESJIFkZmkZJuaFE76kigYbWk/tNvaTqqrZ67bsyLSaYky
lqG+jx94ao1LwJpW9t0U9WVaBxsOl1N0DQq7tU5CrW941nznaCTqpr+28nnzElG0
fuen8oQ3D68IzPTRGBDdOWpGVl591/k8ORMqe0phYr9id4q1vz5N5LYCLhewj/oy
E9rto9Sy+ekGyFoySb21mQBl8CCTOYW0kha6A8fCkhZCCwecOq8rhYcybE2x1ah/
ggu2z/xnNc+tHLAo+zIMpXPr6lV2fAYP2DYpaxL1kUinjhR2Xj/budpmNntCYQYg
NcGxSwsK45OS31wz/enuGGyBzNjO43zOC+H37wSlkxlxzxNXcFAIdh+wAEaf/mto
g9FEGgKJhQpKbqgwoZZeHx1C83Uzz2UVxtP6KgA7pNsx9H4umIYr4MOj043x02Qn
DdWesvmWNkN8CzqeY+EctU2YhytNsqGoqy9rxu7QO3NPkBS4C+b7asQ4Ls4aStK1
QsPc4KQtjzbojksuO/80ua2Zr3KrnbLhDOMPScP5vUtQOWMHZn0v/9UEwipv49A+
trAtzI5+v7JJDxPAt7f9pjKIyUcYZgjFDa1w10y+ll8WDzzA9PnXAAV4k5Mhzom2
wiHWpLc2HVrSRqhC2H8DHtfVdKKk+z9iTA4VcaffsRidOstppNSYLxj0ecE0unSU
71dYbcoCbUUgW4MPzkq5WXdrO2JSbXOHJTmBImv3pGWD0I0o/FLZ116Oc4H7IFTj
CYh+C4KKTD8W30au5+VFtyd0COMrz5C++XZtuo4aFmNskTMMgu0Q6smt5p403Qba
0rkfttHNs242dCIBn6/Grnwu9ILPU4gx2HdunJ/xrgWBnOPay95Ye34wybpY+RBc
EyiXJ3PtcVB/UT6xbu/Bt37+SyEO/NvT8kC//MDEgA+94QfTlIl6ROF/GXTiFAA/
/nI6/+XEK4BhjaqUWcpbUKEA7xOCEIXzIyk++OLZyH4jr0IPvkH3vskRW6nO8rCE
xFuQ3deqa59JPomNI0WGem+gUq7uUxK0AiYUIcnMkdnyLBHvZPXLqgLAPUX0vNyN
`protect END_PROTECTED
