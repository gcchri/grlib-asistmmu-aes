`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8KTiy5rKBgbGM16lNOQFF/ltlUxHDzWJia82WEz0rMCsOdS0N21ktyt5jF2D22I
alNS8t7EOveOLzuR4RzENZHZ1xrwGJXRHMH/ok7/VED26cFNER+p0HKHOiEAP1RI
Ilnb+SnkDoCSAexebugulKjf72dArYnH1ly0c+u01PkC67lajBrJlBXleoKIEjDY
t+2v4HZxS5IBlV+lLLRjYOGjeBQi7pIEhQCeCf3A79Eyw0C3Emx0PldbM/U5BbIX
+jwKgEdl8z2dwH+dvqQoOksF5cQZxvF7hbWAr0o3MYdWB23FZdnQMbdkGVYFFxtZ
73tzase0SXeKMQLh9uSAjNjK/4a3kdlTsJ+ekl3qJlwgmiFsgSWSOXieh6elfNbm
beqkejFTZKcv+lrkRijqOCVsjbXw8M6KjhNQRIFEEwPr9EGg+7pS7d1ZgaMGlfLa
CLpfWq29sA0TUIhighjCpMduqoUp6T/qNLcWD6B6XkHBFmZnT6/9hfJ/a3Y/h2hE
F/73L+VJzK03dOKBiljEbi9nFUznKubMqHJWuqWVZqkKEduVSSzhFvLIK+lVUAqJ
oDAyl7kQOc+4mMasU4QdA+4FsZwhTCwu/dB8sO7Ky2i1WmSULmy1Am5XpvD07zNT
MKW2Ep2VhO2tH6akj8ysf5HBegIebKLc5zWhv+hpOmFSOgjL1P5yxnvZUGVn8gQr
AAsjNlMIxn3v9OEvJXe72s8+n3EmHS2HIxDn2Z0aAyTliTic0fNNIYCMvltJhZSz
Jy5fGqfUnP/KxboTN9XM9A==
`protect END_PROTECTED
