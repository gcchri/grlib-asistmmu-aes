`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTwu6XsmcQKeu5EblBl0GlQSff8OtaBnkJU+HMnofI4o5CUmGKFXeysb++gMbIJn
l/SukMBJblELxrSAFiaKPNx4eeT9pWnjeAt+A6XvDaW/pIaUfxNy79sDPjpjya5W
c6MPe7eTySW6xw6MDe2XkNJuS/gbm53WUu0LoFSrVf1K50NyRNVVk6P4scOMKcUp
VJB22j8FUjPsmdUdrORvusv32Fhg7aM+C71jF1vdv8mx191XeUOS0IgAJKDugK0P
YOj8QiAbj1NF8wat6IcxOTPg05ehzWdKuoYNI91FvVnXiQDo1AK1Q+QmVpuyZQC4
iIqbYMpV8fELsclwVTBNZNSNj5lHjaTImMUDSSAyJVEOG4dymIcI/LKGVaCqs1Mu
IeFeanc43TJld8VxZHhkhV+giKew0MkHp+SJK0WBNThokr1DzRbohHUQ3Raih887
t0uFHtFLapoTzeb4TKb7Htvn9qpJt12QQk3e3+2RBGDwrd2ObFyWNgeTzxGygiIQ
rlQWNHqldhzHVqlEzQhZXSb/NLD721Cfn2qM4GnmwEIjAYjlLsDwtuN29nDZK6uz
2UGvC3q+kN8zzFceRgO7eaEnRLxD+dJQfSzl8VOn+5Y0ClpUrLtsKABTJkQFtUux
OBSCUgk23r5qfEdAyh+trvrmkFyZvIeAFWgd2VDNDsy0V110qVnX+pJpY3FLWaxm
VwOldmB+BLA9A1ymjunHpKM+eb31ycqCZ16EwSvx0qfckzw2UPWcaPD1CvfVXstT
BVa6Oxrsd2M+7lNFKQpQqiUAjNuPgQFdt4g77YpsqIXgwxUMAeO/YoqxwrEdCOTC
RJ5pAoFVvY8cllBwLEvlg9ivpi+mQgPP8EU5vLNmk9ycyIKm3Aush219fu2z8r8D
jZLrfbFTTR5JOmNl3bKNKK1PYYoHiAZHYTYA+mm2w5huehAec0buf2m0bmDHZNFh
snNkr9T5zWs0GhJX/z2ixjUTGfZ8O0FVV0GqXXFQ2ISqCaY3bpJs2JtLqi7Ktawq
QiMllYJFegvGTqG5AiaRRGzF7JNX/D8aEUBoR0aD6GA1jxxCZsn93Qklb+vxM2+L
AozeQj7L1oVC0rnNSKVg21vXd3LmcxCKVEgIQmo/0DEdmIHjPxZuVlugqLGhfeIM
Ov4aKAmCXlUoLsjvRumCRfD0C6F8ZQUcUotc4wcXAZCF7lRrvlmLRuryPQ/L0TTA
QEHxGxdlnVUkbFLwGPEebHyytZHInQ2tQUbflwVC47cJviwNG/4UfckaihLsBxfH
ckCjQ8WSRuPi4o8jCNDtMMDmIZ1DsLDIB66HjHdD+X/cHSN5jO0Msx+0rgODjuQk
rRyQ4CqKneGcFuqo/7W/YFC+vVDO6Qi9Q0ht9R8/VDXVJL00BrSEUq0qt7yCuFhm
K4S/zN11agTh7mfqBcMQN2NTEt6dr2uwfipLD/LGi+8kgYhoArIkszNKmumcaKaY
8NZMHkLzUTh4MwY0dCm1CBcjMk9kJnt90V0H33k+k7Pxhgs7eCjE/n13eXWc/CGv
g/Hpy1olwtIXaE7cZLoTWqiV+W3zH5vcLAIzSFlNV4zTvmTW36wgIy5xvm37TXci
eWAAjBfNJfP4C4wqPDhcEUhe+8dbYBlFIa1X1Wtg9gOlFzrSWJYvzs0dK0rJazS9
sEZTeHM+PqjA/HVOqLqu60P6UurxZckKBtvpb0HPx976Je7CBniZGZelFTM1YdE9
xAFIVUQYzD677uXLWSEAx0q7XxEtEFbBR0urPo9aOL38anMbM0VY6pbYd3O9VL1t
L7TnoM5FFKzG6X0NvtEdZnUT1XYePv+Vg50VI2TlQR4WkdqWGxHoUGuIMyTGoYu2
u5VMjFmTP4hqIOwUhKysb2pU5Tqvv9Sxx3bivvp5KfvY8U/opZq2b0DP3d0C9sDT
kKGvc0HNWfiQhAzr0HAymd0OmvfWk9uVjwSMveThUePzMOGrP7yMW1vH0/16CE09
PaqcyOybspgI3+wremMXMWDksKjRBRMJZhPMzEuBkhkNm27Uxk8kt9dlKhedgSqJ
`protect END_PROTECTED
