`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z7Itvrhr9AA8t05NtN/qiUpvcXzsHB5nIeT9Mwoh7nRWnF4M+jE72WngTuMXCD7Q
6fbx0471dFrThXbGCw2U/BNe1vxJc7ohWv9/XzpKWXNx2jplHjUfrVIOD+wc2M60
eqB0YhVNOUjgmooEpZ65lt0ZNnQvhsa5n9zbqnqcrCfp9DXrJ3FUiXF6iN4CY/Ry
O+FUimV/QbDlfuaaiygpHoE38x8dkcEJmaaba/Bun6z8WGBhG7FleF/5bqDf0b+w
Zf5dZDgNklB4puTOzxTCeKt8oDgG3A1IGdegUP5w35lIdizkUsaSvPYt58sUHCF8
3kS8gGD7xrCFlBooB8Gk550xH6n4dYS+Nl0BacJ98xEB/X3Rtgg+6/22+FeKEQjN
HXKsnB7TCWuskmTbysZginbJy+wM3dRTHzIBL8eGs6n0UW8N1s/pxtQik5RxL28/
h0nvrjhckH1mNW1ucg8XDdI9YvS7ryjAeoMJ0gthF6BiP3jWVRg5OG3LNfZwV5x8
KKTzQ4mIegtSJzEPe3JU5ynWnPNu7Co3wX3MTxYxMWfdHPfG4zdqNBipa7E/kpES
WxpdmFPwPXUpCu/u+susig==
`protect END_PROTECTED
