`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkVl3KIrJCEDYJF7uVknOuOox/wfR6E4y7c34ClJBlrG6tY3ge1PIEg3/ssGe2gA
jvxT43/c6CQaPqM29HU2MVjErXYHLhOUSEnQ+OLhKsmvzQtziPQXEMBcLsSPkVuI
y8Ss9JSusGTZSb6IuPbrCuRM2IjmuXAAl9dKFwQ2iWOIFYgGv0B5GcsLusHkzTH3
w3pHsPVYAhOXiW41rop77+TV+o0Z8RcQSflnzqiUVDnlk/zlLjgSXrPEbzk7Lp1f
g+NTWiQzYa555/DNEOx6m382xHb8PpwWPZb85A+k7ohnR1qKBF6eyVxPwRxZVpIX
OGWERPJoMmnTjFpN8Ifoqf+QodUD1YGuhHUWxzfyob6+4aIYbjlSfNAM2IRKRBJT
OfQ/BzaIvH1ZbcwMLytnR5syKbiC9fr6/jRn1CVgdgZCqZwkZHzQsVVO9+0RvBVO
+aY2khYGY46eXLDo9GALaS/iv9QpBTTU7o1Xhgu1LqIVJHcCPZAhQ2VJ++2p53+D
o/aDjvHVtSbBq9fgoswG8AqW2MSzkMHSaKUZ3lSHv8vVvSMwRcrDgLlj4n1fn1Af
VGkEPmr0Sqf6tH5RHqxbNOhbgt34XFvAIupf8S79zhjDh1/dlotuERVND/nJKtVB
S+noqJZljKLmDS9jwyBXinN27jN0ysGlBsLVhspnZ6l30HR7nFqfNY2l0RdUYy6m
DvaHePLpxcJAm2IVngbk5FPpDCDNot52VZasoDlEHxc+8AKbHCCCZvZgM/iOChIV
dNvCtp752QLIt9UoRKIY4VDcDamZUp4UF+jk39RhIm8g9i17DFKpprDpo9pD8Z30
sOemBPxhAyGft8LZb5mQtKhfPjLfSuLrFOEgaj48IC6CmXMh+hOksE6vjpiDoyy9
MY/TAD9B6TQxkB/qT/fabUiSS9K2UjNUQEtdezqHa8v+UjF9lOSOjWysLBh0v9M0
lIV9i3RRZ1g1XMKInNYjUBZgdCyk++/OD/eNqaA/wbGP98Csgao0VxcPbz3yYfgx
uAAzP1v5aaifdvYZD8onu3TQH+SLCAr0bzpLre+yf2nrQHohDjWdEpcifbkgY2O3
l0L67uUgdIp8KdQ7tPJbwgkY7sV9xQ5jv8dCkT011lQq1jHXKq4SeS2prqA/1M0o
+jqQvR/XFHIjBuyMKDVrXSWhJ1i3HTEw+HtoSeK28TXIOzf4w3UTRV3V0IL7xaVS
OBuHYq8nVtCrkr97nwFPdVjqSp+AyZFAiJI10QvHrX7CQnYScYfpCJ/OrlXw3Bh0
mRrbge9RMYmmC6m4RtdCchSIltTl+O/+AZ5V/d6dcpOTU9k+vZvkO2Qf9C8dyOT4
w0v99ftT3ZCGj60Av92FzPKdOk3yQHknmTv82DEOtx4mwh7ZCTPEm7ESYRbgi8+M
yR5AasPGNWIEt3LPJmhquAqnNiiHLHNUE4152Eh3OwZotbqG0mffIuv79AkAbJw7
wGt/H332e5qndH6Qv6qX12a0qmrWc6uFbUU1Hhv2dpRm0n6K0omejh5XlS2PJKep
a0tscPB4WTp/rMs5MC8x/cncNf1f2jd6PoVvDGDfR/5XX/E1M7+CCk+jWBac+Es8
sItY0gikSjhzFxs9srV1ujcxQazOfDq4p6k3UeJp9B7km3T6Rz5ME6JK5/caQNS/
6US72AUKqQMUPuuWhjAghCuBdlbB7prrsEfvD3E5D9PBuVsmzzZpxChuOmm6flEj
WS3qFD2Ja/FOVIMKET++Y7JO3StTcIbs0C7Pz6YQOqJ2O/lvy7waCG4YfRhc1Do3
MdMOf6/2CHirCLO861PFZoXmKCst5cFFut90qA29Amx7rudISMk0eo9m6ctUVrRC
zAAWY0HNSsM8cnti+t9NJXjIJKYbeUu4wqNH3vZrKQQWChjqOj7ZMt/yrW5Xr1Lt
1p6Jx00DJTkfTcHgJUd9vYGiAO2iN9ZDm3StCk4lysHnPPXAHSGbpm9/xvIJATfg
W6X+r3NqzXa/jvZuox7mdDU+tfIgJBthjan++lQjIDs4951wr11mOpAB3oufaTHx
S3ibSha7ROmnLzlFW0wcf9yydNHLSxvlFQq8it4OIKAn7DHULHFltpEuMX68+qUr
OiQzN5gLOjqAzIrqFN/qYhouX+N25nRez6fqXm/P24jrYU1AGqOdP1lKjj4i7D86
K4YZMNjxd06G2+t7XqZNVtACAHp9ZQn/PzYQDTxO9YGLudJJKF7PWS800haKBwd5
93rp4LBFWdkHIAu87t7jvpfj6I1QI2MHtw93+VmH9KjKlaXjcZ8CZS/wJf8PiH/I
EAlirfdhTS39HqoMg7MyBbTq5+Wy693YDUKvM8LJOBfHzUVSs3IEyKo7HaE8d8+i
pJjO3xLAkUHXxMAxQQdfLVSfcJPdbwbp0OXbEzCAnyvqL9ItdTEa2sjiqfKpJ79g
VpuNF9b5JwtZSkMLh8GaqTcHnfwgruof6re8kwgJxCm452oRSeFY81DkX0F0cipS
ZxgzPZGKmSilpv+q9IciOMRS3q7vSY+zrL7w6ySo/NNOthexg+iwStxoLCvreEK7
MO2recB7ZP3miteNuw024fXhykRpoIoLx+iR+4WKqXo4Kx5u4Z4FSTA+zqsuXtlB
7SKwwuq9FsrON3OSrdZidnAcbhtNl6en36y4CO09blLg9JcUl6ktCMgoG4q7zYPy
vrtN5RhUt/sHIpf26HfnSafpSpmiDvMWAgnSfKVZlWPPqbVu/L30QP2U4PM38ZGo
QK2FIziAvykecyaKeZChuIjg+4YSpcae5FIRbc3eLVWJQpaijfSUG+1KKaJhsPFM
+Wt34zt0MwAaF2yfQJeT/hlQb1yTynm1JosiCymbJyEA3HmWp/SwQnSMB68FBQak
`protect END_PROTECTED
