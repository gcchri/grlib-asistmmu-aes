`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDpG+CdhJBad9iubChNbefJdTYpbnUaKU2hZYkdCtInLFvJ4lg8DgX1SdqVlprX1
iF4Ri7caPtOLa9Et863TrUmE/aonH9ijYpCh/9iEjKkiEQIg1amiKJgbHOcIRSUa
JE8rlrP1wTNOV7A1ROLgY+4XkHsaylkyKg0dSY+jTeo0i8kd0lltzUkRjMMHtKgT
DGKqwBN3CpI+cm52aKRUaAWvkNmDNPehDmzb01+nfBo4EDhrdiHmuFFZLdUJe/TD
E5oxcwqmZW9io+2VYNQngIHeIyb+SQ4qognFps2xy5rcQpRQjhuzxn3iAcQfIw4p
oNMaGmnJ6vvhT/Th+SoXtGmecgH//RVRdtQGVaxe5TCWa3B4MeoHcS3Mz5z8syE0
`protect END_PROTECTED
