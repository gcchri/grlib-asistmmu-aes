`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WiwChcMQCRreGmRv4zwS9/t/xm9wRkBbW3uaRc9M1RUDFWUhH3rcl1KZ3MvWfMqj
RAlYW3Q/dxM2pknY6LUnz+u2Ez2f9gYUhKIp8tp9ILHvv+5YgW8YXth5NMHVpbLb
54IAW/4z8EL7LP2C1PTxZFJ/8++dUY67LBzvLgiqtV/4B28huOUy2rjflFai7H9E
UgK/TmVcLvNcUov1bKcchUZy9evlt+BUp5agwqeYjM/8TaeyLFc+ChejkNGNmIFY
cdFfLAcGmqz4Y8BKjV3xg1BiNfl87oEWg9Vj2DwrYnE7i1TT21lqE6YhDzMjCC4d
`protect END_PROTECTED
