`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9n9rPFxTM0NJwbVPFM/bwIpdWTwZ3zvg0UiVc3wtz+pySFIQAtapqrn1P+7RXh8
qqyJHVFdpPPc1GUysguPe2spcGQDSKEJ0gQtwrZTx/paQbbc7UyX8QbqFB7QyhGa
K1VoESUdHuQHclB0jcqWCW4E9gWTje80OhTpg9mOmVqyGEk4/S72nH/cwnqjvQB2
RQAiEl/LaRZOPKV777tfQp8orRLsnpH7eoyFKM8ymIK7tZ8umMbsK+wbjA6gjjg0
Ba1jY9/ZUgv1Xr3x7Ksk6VBtI/hTVN1gWEsEeHL5UzQTAs/+wfi8DKNZI6w+Cr02
A+7s9vjOXVL1GDnaL2E/oFGJ5BK/y+CIOegaX9boop4NqxEwOULQgjGeDWldyReH
8axODDB1YuHZrlvOuBCXqGFQzMF8yV7eZF9wrUiQ8f376omdVyBHe3h3OFUnIF/Q
oWDIlmiU+jSNr65BJ7t1Bo6wvNhGSwKowpKHfIllMNMbu6zxQ7vXta7UEB2yzo2b
Y1MuWJqCS5tuwZPwD9kriJPXItSdOELI96bO5efouaeVnwgXeYe2yJRpLsS5vevi
C0tsBMHE3/JYaXysNEeZXG6GE9SFA+EArSiDJLvGJm0FbSibHgka0Ied0nLZ1Q+C
S2pGqJjaDNPq6TQzl4fL1mLisYRp8tV3PcMy2qPbfFj1O+ElxxdmjFoWF8JtYTwD
UbsNicTE4OmP9Apv9GjM/38ViNzC0p0WeEam0v8u0WT/XvHe9gu2ojuyo8iOa4NX
KCaDakiB4WZi1yAkAmoCqmhutl7ZGAwIVH5xZ8JAYaNHKatZXo1GxqCqruoQQgSj
GBAUJQwsKUfCauy0nZGDnNG18U9jLB+HEt+ZLO5RsMZDcMR0k32WQjn2Nt1ZDUPa
Z70zYPnVFUjjiFSKcDw18G0x/nvlq8fIRgNiwAO7B8Kp8me8ozHZZ5MypCL7zcsb
YDRz9s2FurrZS2csi9OStJcbpKrTNR95SwiNDGvdBNvVQ8DceQD9rXtZ6QurieqI
F8XlakpnsYms3LCfOKhsGtjm7W+YfjtbrZavHOmj9pAlak9RDoC7ibuXm6k1EmkH
9z/+ZWPER66E5Pn4V2Oa9P1SJneICInKgqEcxi9e9zz5jB2NXUl5TYBj9PsBUdYX
+opLNchi3EP1QLMM0iK0EoRC4P2bBGjI3duu+U8eFh1kwvMpr9CzdoW/73TQ2CZJ
mmpwN5F7Rb4U0Neos2nVew/Si4k6f18chvAS0Z2lAJ/bg64P2KmdoxqrSmFEraGl
BFM2IOCK2HihxtUTb76ypErQyx2AdGCsbjv1dMhWgQaWNqKvGjCnBxrZEP4kjrzF
9OS73ATwpxFuDyJRpo7ZQ3fyaDcAUr+S25vStLt3MMTniMQhd1UhMJL/l49wRsco
A+5fcRBzQYKCXG7kIDhWmeIrQyAvnm1VAGVwKuLDVaUCUfeXwyZ3JfFKp8X2vlyt
3FlCjWwJOW7mKJFbetHVkz8h6xLXjIWPUoCQdFAJcDhHLA25Ou/ALSQJZHN77c6Q
90j3omYCUPU1mH5JRDivd+H+5slMDnDRVmk6SCVdc24V+5/RKt2hCfLLThH4XLzK
+vi9OwmcvN9E3WG3Ue3ERJEbV49KKRAU4ShSg7ff75qZMw+ZROFJCKpgmf+ohqV9
UAcqjF+GjxTNTnRYIIMY24Pay60H5bfZbSiMiAgsPDqr4sZIbCN7EIjJwDc6lelJ
E9NSgWBmRRDEW8QAh9Ub8IjA+VBMF9SNvyD3MqF6e9Y/uK3TReKLJ+OUEHp3fYIk
SfOnbXqaNy/RJKhZQrT3SNO/brMjzwRqwjUIcd5yj6PcaAp3GGT+pD/tWCTPFecx
8XiqchM/gJ2HvLwaR0k5wh85e/Q5rGO4N+qmOZBnzoVRqL0B516eOuMEg0KATM4D
TJ0EE3FmonlCcuDxtg7Zbfv4qS0dOtpfP3G9nqzni01GHYQg6jAMH/CGijoa1JqU
ucLTy13PJ7Ih82C1TN2bFPkk2fTHZeehI2BCOCIsplT9W5dWnWM6q+1GcKIopZrT
AnnLBpurkRYfHAgMLAaV0LYA+R6YxmQvKEuaVBFAatrCf5vN0Z5LtCJkJ1WGU+UQ
o2G/Qd3dYgYFbPXDalvp6Lx/qKnyzWfk5jovNYyw8X7+cRVAK9VwQhzFOp8QYNk8
zfddCBVBvrb3+n/zs2NWR0wxv+h5ufeeDDMDe8x6MaDICmlIbgJIoSFodGge9sLp
IcQfU5Xr1DgzIiDxxDDnFcrm4LdwkmcC/ynAfW0IkxoPHLHOPGqvq4jvVghiiCLC
sDKAI/dPjuECPd0vcS4ifz5kF7vkTuWvqMRA7F6gVY+56KbHG6YcMAGYx8nFT5Tt
rnvkFRJ35CV3a6Ge63ern83f6IrQXeezrUw3k+oKmjKkT/tz57/pdf/ClRdLRPQ4
OjWPFaMHD+Ld9k5KIkuo80/vskPkcVUJl+reOEZpsOPR7LYIMxkwWfwOG9C4mJPM
zhlxtW0BlMy5MHIbhgfpE8s1PVJw1XQaGiRPdWYjdQnJ3RipLQpjg/piIVqmRKsM
UBzhrPR/NI20vnzCuv5r1kkXwByDOWmtWBDcBqbg6qnGHFC9zzkvHuQsbzIWi0Hz
O6vRw7Uh7lcH/sbhKsfiRJO1w95AtGFrcFrZzK1vpa3hlym2d2BRkFDkqBIgaXp3
/EUC/GqbxEDIYLbd0FBv/uedqmXgUpS6XDSZy4s5e09q1SqFCgXZt+K99bNT15K9
DZzQWcO8sQpRNDjHjnBQ42Edxd3PEnhELBY4E6tsmKtdWcb99orTN7KjX36uLJ54
tqUDRN/bg551biOIf0+TUG3jBXfJrL8j/vQpBOvxLMJisxBZzCMy8JImL1mhnL0a
6nCYRKQypDj/Tx3Smh67EH5HOjcrNuf9DMK5xMhx43A4/+hM8uCgm88Vus96dWEz
lfi54FtY8ef7ny3MqzyuN53meo/O/xPpqgMp/RLhWGBqJdded/pfGl5MR2YD2/wv
LVYYbC40p+2kQfsJyLewmKlPFxeqyleBXwWoqRSgDywAPvJEmUZ5KI1dkchd/7oS
lMzGBah621G/gl3w3HvyAOATkaWWykxweGdJDJeQJCbioxHIDb3dCEdl9u25ratk
TSVarSDXfFDYY6WVOat97CLIPvMHeynrz2sqfVCxpR4VF06YT7GF7ZTjIyh4+23f
rLCeCeGI1YYS1Wt7ykafuhTUbHCDiaDs/omA3alOEQ6wuiGFGCI0hM8caZ368e9w
EqW9p0YOJwW0c6dCZurPriX61v96aY4+Rja03f0c4y1lXGYTOmMXF9mPZ8r6oo9k
OiPV/vNP7w0objPLt2zEPGCTDcIso16Zz2p98bMFWSfzrSoRnuqH11W4RaudDBsf
ehk26tkWBtHN6J/nI3N9ny66mO17IsQoHZTI5pPIv0GF70bvEioQ3xx13VwPU2NB
kf6sW8hwNr+CT2ju6CyC0Ci36GEWJCUa0h/D8yKKoV7XcsoXdr1q0SJghKErSlS+
SAZBjB/6tiXpNoCLT5D3aTXDAO3YS8C2B5+7SyPv9VQkC+CTyNTZKA9tIKtwx36v
6vpX50v1xlRgc28l+SR5zIjfU7ZARUi3DtIwo8obBU8x4om99iRvuTo0GkMOVcEJ
RnjO418jO7CWymnP1ZYA80WMefHnDmju8Itqi1f9ys1IasBmFdAqC53fcW0i1OGR
C4WiHB7xlnYcu/n2sFfqG0h81+g4yuE09TAO/VVDKlmi75S5HK8xV1WfzoLtuGGN
Uj4/G52JhGe8IPjqlbwLL7ax/f6E+mvQVuPDFZIBWLRWTK8ZqCjcVxqTpiR9zxGn
Gp+10/P5DQ/MyeBWU01zvFpIHORUxbDo6Y9vvOm25P6LmAijqoa49zl9sMSGqvo4
ygwPUZBG2PP+NGbXMMo2BTVQr7vHM5Wgl8wOzziK/7+l1sC/Q9BhreiZNe49nlpm
7h/ahhXbPJci/RVLoVOXp1E3mo0apZcxwzI2OuZ63+j4/uE5hGqNjzWBHtMDjGpP
5qN4kD1xgzwKuhaWYxTSnzm4skH3qe9bMHqbfyrDOxvAFa7XsX0aQ9prCPHNSvzZ
4WBS30DHm8RPiLXE1DUKso0bCXaonAICaBhjWT8C/v6BjlT5MoVTA85tnK8s51Sh
qMUxSLwOVxOWJq90hK6+YHJXA56rnlL5MAz2ABZYla8acKpJ0BrLrqvuk1NNR3AU
fvhjeN8Hx9aAryv9d2CMpjbmNHJ/8SCIkugJBarHDjB4Jj41lWi6l7A7pl7KAI5P
14fxpWjh5TUu96J4yDCfMABC99r1bAijjRyDhBJOUqDVQkMqT8ldLWTDR64UehUj
7snM9KccXNd6GqmKbM2HmUOuzBvesPj63cCIkO4OMSD6h671k/WW3EuGl7IePARE
Z5VsSFlFebzHlkn0hrtuvltpy4ttQdB7gGcFMnxXusNuRZmjXk33S0VoOKdwF4a8
BlFCMub3/2TXa1Gha5EPMFU6a4aw3fkW+StkYhocxTvHjtB4fO0XDSogeTWaIxzG
0l57VJHgm54HdZXV+RZNoQ+9B8PaiGylwW0Lir5qGe58pSThIDsfB6zpWP3T+EiI
hRxqwsr+xMj/fhdKBE/03UAIP6zSVopmAWTu3xINVYuGL5Q461zmOCMuOX5ZLe7l
gi8rULMXg2N1Za2ZieCyd4AJ+dMMF3ELn7JPlhAA47eYW6UUMzWT6SKYf0r+I9v7
es2M/49hlQfxga7glUvu0e/J6VHA6f/S/ULOlkbBXprLR/SUbBcTmuZd9rU3rLkm
rRUQDt1pklF+djq1capqxzU3v8kpXdPu/70T6e/zIAsHdToo8mDcbO+S0R9qR0Nh
9Hfin4TOdcp5CvbSFVXbNo2rlbHfdJpSZPd6lvcq4773nq6LahG8JdOrN5KE95bW
/YTi0snchi5fu3qVyh5PPonZRXGPW1yu6xpQTiNYi2oHydsxGC7A5sRNNxbKMNVd
ez8ePtTe7nLbRQw1gp/QEgjK3CIDPLsTwjXvp6pRp6md+P/s93kRrgyC9gNWxMBk
cr/NoruiZNhKBHaHy4MqXW/VBsdgbLYnqhVcCCedqaMPv8Z0uD8QOWnAN0z9IM+P
aFd/QztYlKdH8FQS6CI/JfMazrEY2FUDg7l9J794P+y2lppOlXTny+NP9AU5z7bg
TWewU4gBQKT442FKewg6Q1DrGI6DivqecnTqo69WSKuZ9sowLqI/UEzRR9OQj2nz
ZvQ/zYWAYEm5cVtOzNbYvcKqfLmmvaixLS5a8wlVLHuSYclo53jBv44XOWdf2uck
n5NCYlaii54WuQ66H841Af/WhvyO9P9vitJdWCAz9SqD6EPyHfcPbmWc5kEHCY4h
o549tz6PUuemxRYuDdGWIrOzq7ftdiOT1Z7Ac6+9j4z8dl+SLOYcPv+9aaW7SBN9
xINS8biU9WSaxvotlBnOWmn1DYHlmYYNJBvyS6zj4hk=
`protect END_PROTECTED
