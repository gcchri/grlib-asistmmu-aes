`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jDhsRxhZMfuO0cUJeUHSI1AGMLGyFyNRN8bU3GhtWU3O3hsg6pacqKuRqmP9/7GH
e6Q2ibfnKWMhDYuoL5GfvcksE4zhR1W8/lLnmHidFLeD/FtYzia2QQR7wLg9Ci2H
tiwS/7dxPF+aAEhbtrsHsq+6QSdLodTA99nXhysNGUk8t1N/u+SD4zvwn37N8tO8
h3J3eifg0xBt/uGiGtSXWEB7BSjbaHMiSDNeu8KuqA4kggQP+XRe6LFNIDuHG91+
OKnOKnaTsg6Bo1SVeQyAJByzKesMEBA1xFMhD35jlmZMlQ0Erc/v9c4/rYwbw/xw
KAwO6abU+IeDd2jDMrFtAehHe7v2R7dPdsRLDwDcaAqYDBGNfgYwKqIZrTT5+vzr
X1gsH6zSpkv8ygJQHEHimjK9MmwbhjVdwWnchKjmapgc5SUOGimD447ckvuOUDJa
`protect END_PROTECTED
