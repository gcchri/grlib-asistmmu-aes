`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FSVi3WnziSx72GNP6Z5V+amjFViR/yRH0WKXww2WmXh8OQKfQgkdrN6GNyM4iqHH
wxubJ82fp4T7Cx3kD23/Xfccd4Yf/R8gOTtzrYYoVrQRk2k9K0mO9ExzA48nET3u
5u696y1iMNuWRI4qnhqMT7nx8jH77rsBwx7PR/vH3tw7FkRMyoFJQNx5lhvR7StR
jiaaBba1VelrN5clC4n5UtLx8KOO4AXiLI6fg2uFgdyWfGa+GefyfYYK3E1xV3sI
uNE4omT3UJ/IA3TAJeK4TJXr85dAom/ZhVgIHpjChrNQZqyfq426vX2zCZy7Lsyd
bhF8YtMqZZ6K+C3ldKd4MiWv+ZjZa38BO3s8wYAOn/wz3KRQyWFMEDnAfhJyvM3t
PI7C/wvfQrJQRjQPegkpf0ZXxn2q0M1yGTztJD4jsxd7b6q2W9MOq4kXuWMXJbJq
qpj7BxN4OuGt8mCPzyTvufnP69UEtSXA7vkXinux7fWNl6D9iGFJV5yn/0tk9JAh
262UVNAxOyNxihHd6DdQhXN3ASi21qqlCUgGCwoeAZChStBrH1HgzqRFOg3UEc0U
TcQbaiMoc6WlvYNw967TtN98yHvXec6d2g6qZWzNaV0swAnA5IJO7YXvZ6JGfNOb
OgB03QPidCGV9rSQ2aqLzBZ3opMFUucXWhe4ZFRsnj73JgfdBDRwhmBBzrjgU7Ug
lVMrznqSP059agXeuz2+iQW7CFefduT0pQ70c3wLoERpXoNNmiDRkCsOUHT2CA5b
`protect END_PROTECTED
