`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e0z73EltpdhaBCFefMEMRO4L5DGSIlo/ICq/xCX4zIfSZPUjzz1+Fo3dWCxED5Pd
PQU04ylNipDEr+zbc+y+Isn8jqDuD+6CjAzuCdOpqPUB+bXUlEgjru70wkz86kij
RCpYyaZbJv6pb5vDSp9lxts/2NrPtkJpTO7FJu7m622GbOTm76N7e2lNeqZtc3NJ
3bIPbpWK5iaOLstGYOlCsCaSjw4hMJA5CBAzLgiE5CoiOtmJn5C+6Y6Lxw/nwT04
2k1xYTZzYYwBItLA1Jsvr99nO95HBU3rIX0nwxCbShde71jPXzbD9YI2V/0rUpOb
r3WqQOazFAX3eR7r4/+5GE9tMj5zgi+KXkfXre8t8kljHj/iGJlIF8U0IVvmBPL3
3ncHAFLUcA9PJPRi6hHVZ6ye4snJmgLnqqOeG7GUD1rBgwKLcGk5joDXqxiOJnpR
5cQNKQFtQXY/FRGfF5R43CZPQWhJHABYjPHG5IGCOUVIynriDdHb92X01cEnQnQK
1TOnzQEtnJH5FqGQxJG+h7fNxsleQoYbqB1tx67h7C3EEER56qF1hheYwNqqdqRc
v2eR+MYFhj6ZL8IXl5lkiMlwR6c0TT5aQtq1YTSysrQ3bLxo1yRSG620VSrf4l+t
u3mAGB/Ex1PpBxdE/GssxdabZ75Wck7jTiOVAr4nFb0yMImUiay635O6GmPbVGhr
Hs7g3JcmhKngQujqQ9bo0lv7IEvltN1pX5jLzIySqFD8HW62IK7S03TpsybvVrAo
ap05+gQMQ4OV9+uX5s9yYQMa7KrLpiuRQHkSvZPgXcYszMXELriWX+axmrC+692/
SJpKALMld1yGWGVdnDM1vmmlyK6DMi3VdEzQo/+P+M+UCCxDFQomn6NW77Xr0hQA
wdHC7oEY/mjcjiiSeWTIkr1k7/vo+B8qroz2uHqNFpQEOXFg+YB3DKJ/igY76XLp
PUbpJuvB9l/sVdtzYOGB0Y0GEMrcE/EM0YReSVL5T+bJbmA4F31gLM/zW3+IIEuS
EXnD5v9QYnRP+kp3QRrQFf9mYNdxM+3QEG3Y56L2xp5KtxsHV0fki1+fOZoQvgQ+
krMwfgeIDom6/0wPO2CYA0a869IU04mifiL5cp8U8bg=
`protect END_PROTECTED
