`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCHYDNBa7z2rAQh+qVWvwex5vo5tL2ntcyYSuMPSeOelHiFNEuFFPWiJ8Nc7Y7or
6iXQ0G75H8lh+CvcVRGh+uLbdhelDftqAXOj3oXFjju0n2a9B1FkidrhK8I5MbNx
F6CmGpPL94UQvg/gO2w+RSbrwvXpjkt27CX8uujWxZvThl/ZSZGZwtLf/Zt4eHtT
utI3j9rGzJl529fnf4VDqZhxPFpS1xMAwao38SCbpO743yfZuHWq7Pwuzdak0als
FIAzC0lZUdlnV3Y6uT3y+A+U4Syzjj8boVo5HRrcuewN3wKIGrKgLeb+NPgCFPR8
nAs/fbJ0yfX8XzitvT5iuxE/3Utu+XAlWUpY8hBtb4VAscoriVoc/EtQj67o92l3
`protect END_PROTECTED
