`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l5lobMme3PQlFMvKvmhtdAFHCsM47D7KwAawDS7/IPqXLd0si6JJtaOuF45sZuHZ
QWpQ3Z5jo3H4+a6Iehlf9uikwSRsQSW9hnQ2Nw8nfHcxnAmpZ73ub4U45jb097Yq
/mFuZJwWkS9rEZbbehMETTWp/oYU99IicZi+Z1BLUYYh3/4PFoQAhIFlvDINl9vs
aDje9DmPDms9E3ouaYCxA8FgQeHmFa+5FVEklPk2nMGTi2hwCyUNBsOXDGsmesOl
yTesymKts28LluFBBV+iifbhPNKHyRN4UhITqtDNb5w=
`protect END_PROTECTED
