`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9MT+WB8tenAlLWQwwTX0c9zGSS/0R5o+Yl2cFJFyci1Avbno1rP0MFKS5ktOB9P8
4Rltc7BlOk0sOgY3T7KhilC7WaGqJ4pelzDcH1pPKTGY4ezhjLN/ew84rBkPTHjc
ez6P3RsSywUnwND6g1D76x8vLIZvjECjW9eDSgsX7m/ifyHcFTaBWToGUNDcXmbs
RrN7YWvOQ/ooldjZFkfOvJvpJz+mi92sr/W91jiWxBvtg99I2vATZivznTY77y4K
HOzoqXdTDAtw2As2dcWcQQvdZV5pZaALQeWTAY/ip7AmC5YmMb9/R+F/quOWA3Ja
dtWczhan2TwJQc8qgKddEe7G92eIrJV/ERy/5A2ou6Z9w5Bo4XgrpnU8zx+oZ6aR
qCdrgS19LiZZLYt/mghhoin5FEsAUjlmmwRBjbDIchs=
`protect END_PROTECTED
