`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qBubL0FOrhlW9r2hlXKp9UJuaqL2Sicbf2AOjIM4QpJnyIM+4tfo6x4gEbUbvKhi
g6CnTF3q0z25VnlE21qBF3baai4wRFEaxM3E9v9VdWx0LwjcaoiKJXhZQgTFrorG
vHoRyP4kJTv+nOjt8OH0+ZTlI8GGXP5vALYuU8yvNH1XJYimOYoEB+jAVpd+QRwW
GNQTA4YwN4qNPHAodFrZGhdWKc82bOeGrOWlus1JCUaRL5JckCIjSkS/rGiwo131
FnRwvVyW7p8kCTUX/Z1Z1Q==
`protect END_PROTECTED
