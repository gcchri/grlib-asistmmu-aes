`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m8R7wOJnprb2/iDNYM+LCSzaHoduO7yiJ+xg00zfOypuYTJRnZ5bm6UGt0vJTLFG
Lyf0TOY7FIKjkShyWCUwNmaAO6sz4xiL6fkYXoOca/neTh/a3jRoeKtVrZzb7BTP
wgB7sazk/HYrBZ29YKs580CQ2emzGgGsjnWNTZ5d3G8r+9wr9+YS3+FkO/RDIfGo
QGb4hZj3ydKt8PltsaHsZsxjR2XtebBIu2dpX6qoIz39U0KAwK1YQCAIk83UDhdA
qnvTZJNvGkP4+sImqZTsGdiAFnbb1tAW96MYJrt06THDhaq5prmw5IVgeCXsIa3s
VoyQjhldhiBLt5vnSiZgrU+ugWmZ73wGpZy7qpquCoaq5x1FVgVm00cH/mplpoau
toCNqssQh74uvcPbCbLLynZ0fyGjl1s2xFPNC4zv1p9ZEeBfFGB05PaXce9Fz3St
ePxI68kiPc2vCK5NMJ9lpstwfCNs8Dzvwz1ahG4lwhKTHBUXbQPcjhFgTE7DBX/W
x49+cH9e/eal9ua4ZXgEdA==
`protect END_PROTECTED
