`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d26aBvA4pdMxxmsmnxHR22CaRczjC0Ggo/vBgGHcLF8Eq2N2Qp4XhR696Kc922JR
0TtnPs1U5+CYvwEUsTEIo4kqR3iYDUYXTjAOQiIHzwjmBB8hXMrxRGJx/D+3BQ5d
8bliR1rURpccT098UIjMjEE9/4c2lBu+duKr87cyVfnOnPPe/hMBzUXSbWb141Al
3jovyKjHnc+6Bw5frPA4HIWNMcNb5DeF497P0Wj3E119dt+Fu66asrthu4T3BI6g
JNNwOx4FKzEhmFIdPA0Mew==
`protect END_PROTECTED
