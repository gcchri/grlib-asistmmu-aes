`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zCtCbN0Mh1z/y6DjYPzdIF6dTKnb/riUr7YJHhovYAav6knOpzyVRIiGg2tIJGnC
arIJTuutKDf8ftr0l3wMwHB8sPbEQ7UFmLcDstVIaBG7G7piApy7D0/UCN1v2Tjc
Iy9OUvNw5PE72bsbN/5SVnCWij8GKwc2PZlkaJmHOgSD1q2+kkfbHJiCcGvaDyOm
EQ7Y7ct98vU4Lk68HMQaiT3C5sFz6lrHC5WKIqaKCP48TqnYXvnuXCHrwweghMau
RjzHDTS90tJ2e35pRtRPIL9LwbNMmjWed3jPNa5jTM2f9uS+gLQ8CkYQS+5hJy/6
4Op84hCyN/moFzk5/wNEFJobsYclCWT6Hgl3Vx9GI5bIoyAVGV1LY/DTpqKgH/EY
m37uBeLPmyouQa39wpDBNK9md3bxu2oIcehNZSaBFQWG5xBvkN958JBY1G5YzCey
F3QKRED5x/84KwhbxlzkRRpjUdv26e3VAf0ArBSC68Hg+sGCvYbA94nGIiuBMMc+
82cvZ2TAEigbZdZ/di6Vtllj+ISN93XkjhTWwEFFnhoDJCgASBgFm3O7uZ0zN4tX
jzQ71aIbs25SkrUO+kzO4Mh0lciN/Eh6dsRVwsRoIH5QW5XCFgA6+oMTKQBoww4w
y/oS8r4gEutsMN0gAdyqv9BCJnnwgmcVSG998wB75GT9eVwNdEuSsHzQH0Zr6XmN
mwGI2Got/hB7yM51DJm5uGh5sVYdjcY23lBrlTuehcQ=
`protect END_PROTECTED
