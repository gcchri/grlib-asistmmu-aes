`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SlBDFwS7AJRBbqGX5oQOHmzICSovcsiJTDubzg0sO4gaDzwMID6Rxyip0UX+y4jF
RMp5VBNqOyAtzHjC10N/Bqq0KJUWw0rWVZTErOh852yhQK7Ktebz4basyHHbxi+x
FjND84/0WrzVUOTjiDYqldOogZcJ+cyvrzJOnyXMTcGYzJnoP7aLVW5oyM6Uamcq
daw+nUA4vjmlK6pn1XNtQ6bJiXaOPl1kT2pfnuu9iwG5KNUDqNLpRbSTLPvRaSmN
pwWK9Cg7K8hgRFakf3Btef9guD3Qq/RyVgFavLdxlXGfyoY860LemagauNE7GFt1
4209xLFkdnECuBL0I734oougRdBcEIilnhRVf1g5RvenSNrmqw4mEBLwZ/VcKPHY
uGoSK8ebZzYUG4POMUOTaQ==
`protect END_PROTECTED
