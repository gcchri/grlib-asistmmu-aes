`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IX1MFfm1v6qrwPX0GzpsJ3vthAkXrAYkqPu39aWFhheyHfPpR8Jv4b5iRTdQSWt/
fOJ3hR3zXtZAHBQKnmmADiOctHLIn/I57oSbceswnJT713/N1qqT2o3ErIRTPVx2
mDxc0Q5x5/sEXhHfXJqLuvSBwuKOQVWBFwg39vgxFBu4+nA9t1hvtujmOEHFDGe8
fSMjI5QxdVloimnVnbz1BRc9xZAkbwIMKdew8zp4E0qlxhlq3Npcyxbb/qhE0qZ4
7BYgRrTHEOTeDVMSKNdShEft1KkusqW5v4GBvFJVven59iT0VaF2mKde6Avbu+qw
n4IWVY53jGm0Iq+lBLMivlU0wpzgXUBA1CgOygzwji3OxEcmnW9ADTr9uyBSc/f/
QT/8GqSQQAvTJ9aw8DXe/xlK4eyqypQD2i/CZsE8ZCrofAZ1DxZeBFIi1ctxjhxy
lOEaqiM83GMX1sI3RjRLbHdt51LSF1+ctuhWUlCegAkcBtWHA9dSOZhAfFA6wPM+
yvSi7YbXOOIkRR7ZrOwx1dokoSpiap6tfu6VdI8CfXo+zH5g5FVGq08YLy70M9yp
1UxjAn8OETI5Jf02nCQg/zeH7JmjpVnpXEfXOAW8zNxUov5YtV+NMbsjJGlEXsm1
GpOuKRdVltF3OzIf5bDutHhZSKtekzlSc9CiQ5GpYY8jCjGuxpdVpRaYgXMrPAZw
uhG8A77SKcygp9VbdU2w8quKrB3hFbdFLiGrTdncyMoAR92oGjxRt0rhxIo7LhVl
hoR3JbQQWBznHiCd1/Kquc0AnIhlpQ2qXqgas6YkzHlN3wvt/2Vw+K811r7CLrhJ
Fzuy0pC6/IYqIcUiS4X2f6EEG2AuT+7KMuy3A7ESHpnIH1GjcvQxuiyyaxvs3eLF
HzUY1tILorGbfF+x0146h9QfS+v9T6RFZtgKxm63Vz3x/YFC3kiG4XM22qigGmrc
vdjJUqCnk64qW39X11D0ghGiJE4F+Ql8sm1iiNn1uEia0y427TwJ1/Tx7IeXsKmf
`protect END_PROTECTED
