`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBAWQ+b7//H8mpbKyP9qWeJSs6GIY1hG+7IlrHno+GqytRQb0xWNa09jX+Cqio1b
BUkzXVvwtZWbKb6ERwltUXSWT2f1F7v0qEBlsFpt3+LUuXABykSWfEah1ThLGPbj
3kFEI1mwsEYfMgIIJFROmxSqHeBwgb65QUia7iL8maZDZjMsp10iwS4kMKcDWL2b
gmNyrTp7vJgDZD0CF/jc6Cq0XiUM7h5c2ZqTt8S2lnqJadoe0tsaV25M0fRfRcSv
BBRDDaAm+F+HtYE+3oP2FVjUUa/3WVOrLtCSa83xSzC2onjBJImmwnUyVVxLMFfk
10SgiYUSvY8NWExvxJWhnA==
`protect END_PROTECTED
