`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAsLVb76GXWIkY7RUQOO+JKxT9O0CBmfUoxqH7ziC/OTN1eRqobL2ZJjOOhyFpKY
13JnnXrJgWLTIbFZXKEgmjG5/2KugbDJHwCg0ZzyuCLin9vWhQ+gfla+jGLBA7in
MKie76LqSG36QzMFPODH9jd7zH28MluOyYUx05gTGUhSX7kCks/7FrTEtZaKRF2x
WDJDSc9UKXK8cAVs/7aSMbAihUxaB4TFV6Ts9tQR34TVDKCej8wYauM0MxneBYTi
iPfpb5qRz9Zneud3nlzqb4bRJ7XhXtaI2WnZAzURhSuSg+R1j8DvyCk7FD4U5Cl1
OnZgmOqcOClb4Jv23+gYE4ako2Hs1R0xDu6Cs2VEFU8XyRO6u5fO6zpV9kLLZLNH
ezCgeWKlRNeSGB/mVWYkXvemE8UtX7FjGpkbxzKfNE45vvPLRwe73kEsUWTC+IJ5
cnGPJXsfFQ2yKZ4x11PburrZLFJ7t8KG7Q3ZqRs8vzvQcmHHC499LfPqv7LG75eG
CsUOSaR4DkPaGONC77ojOhxFRjzyEBg1am1/spt9IFtVyijuqaQKTc9KVlD+7c7/
HrY54YThjKCDKlhvQSFpka/JGtC5EVH7976przolAnCx8VDItMZot8e9/pDDAOGw
kvsUIQmIuUHvdZ6+K5WHiYxaJxzV4Hh776xVZGiG9Ctm6JeB3OQysvgFUCo90tHT
x03srvsCcPtnBM5QXwClhIfkgVY71OFzUeI8DUCHce8cKeODUlkA8D0rRgZ5/F3t
bpOV8QVY/b1h+wy3IewJ2eliu442SbpzFYAdeGAJMUodmUWkm0s4YMTBF3KngV5F
NovduMFkYME86q57U41NJhSJKWKYp6vcbV0waZKwflmirFY2t5yb/SG7wsdEV79s
462C2UEvEOwH72oqaOIa0e7pKH8MMlF9bYPmna60UZfiXFgifo1tUUv8kbFNRz2Z
`protect END_PROTECTED
