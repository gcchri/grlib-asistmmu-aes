`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ilDEkNMLutRWPWBm7hhpK9V47rgYfWxYf8tUx/Afp9FGidKk5yF13hvHgFa6Iyof
L877u4yqzwT9PkTsr/pU+YcUpq8Tiqrpj2AQtfBv+J/OKd2urlsu6bjEvrd/oBUz
ytrF/lyhXsbnoJfBVrc/m2hBrGXownVgIGr6mIi4TuQBMl9VtgY9mW5xO6vlClBQ
4nA+TkTrDyMWV17RZhPZ0I+SLJAJQGlyBWKxsM8bWWFlD1aNSXcN9Hsrk+36Z7QL
9VJEOLxZu2QYfIGY7lYp+3paf78iOuVFYUa6KkBJCrPQsIxc9u0wEnjLg1hdbkC0
/3OXfYE0elx5y+2S+5DlxzM+29qmcbky9LgKLwty5ozNwbxvcfxx/CuFVRzI9dM0
Salj1Zdz+l3/s6L4/VOlfePsjilEzLaqmt1xCklaa3TyD3bEFetJ0l2OtCrL1QXC
CD+60n3/RDOOJXCHV6XnLlxgUbbVogrXLwLJSf1XyKvnPLQJj/f7CbmmPVtw4UV2
dB/UwzezkHdbwDovsoK/i/gDwPsg1jsftyRfd80mqEQA53/UEHu9Evqf3+6IjSgX
eB6PtkKd63zPWWIqIeWEZ6eySjplboL6gb8I+Kjxe6llkjtFtrN96+HzrT8W6ONi
wHRUnqx0BLBneM9PpX/+eRYh2dWT54kYGjn7jkAj2aHfijlUJTBloGR4lL/eP2u6
ZISgfFQmrtxQaMqnZRagti7l1ZbArDQ+M047EcfjaApJzagvSG+s7HLY89GJ4PRj
y1nVQhF/kw7fo08A87mDbHsG0/akS6oAUzKBcxUt0lkBMVAz6TFqzfGRo/bLyfJi
ZwfAjQgTKKfF5gzyaZgKL/ElF+YDwd1NKhYvvAXTktEwLuqrSx03F4mLf8LGP3nD
0oBwvyRiIcpLnZq7viSMUVtFTqdfWnoRmzlMcTaYvzMvn5wxhy+NLkORlIpRLL0s
YUlCismXtHegdTkO6wX9szwfMyEXVzc/NokgPlA0p2tAKZyUWqmSSUFUBymtCR+I
oiDqXSrj2RvnpDqvood4si06nmdli9Yh+q2UEObCdrb/x3GWWu9MP2so8NEjUDV8
ymNwn14QRsAjFxBUDhZV3p6t8AjHodTOEYrjqOVdjgmHGAIGPlo3flm/KynldJva
yXDwWG5Uz1X/Kr7db5YHy7T1PvbgH6oXe0666zcWH+H/09GNOV0BjLRvTs5ne53q
Jh3kzOLGx2bqCnMGcqqlo98YQok606mPolc0EXwDEO20qoSlwuK99utwb9cxwTTQ
cB385MhozYokcBKSGxJa1dX54M+gIVVsFEVGOC2eeX2jQFzRA5wtrH4fKu+xatGg
sGhyrpItMMLDr7M31T8cDW70iOzMZfuwsCcHnmMBORxE+yrPFnPXTVXN/J1eQNvB
oYP6fEBXX0t5iwaTDaGVXL9T/aP9nVO0FRUbxNO5JlXyI0lGCksG2pGLE+JpXy3A
I8a+ffzNv67crDCOkQZWPI2/Jb/1OcJnin+vjRMR/yQotekWF78elwfl0DaZP90Q
qYD6CJsdpBsu0HURT5gQtEQFuB/reJSxBG1McLgSgmyzkojc9VW/w+YmP1BCVkWk
9ONFXGe2Z81nUMRH/+kN2Tl90YRRiCEh8TxQ1bL2FBjXU7ji6QldDsL+0uobSiNz
dR7p+vS1CoCHOuJLi65x1Q==
`protect END_PROTECTED
