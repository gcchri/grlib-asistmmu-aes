`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/m3nqAaA2xu+o0wVWf8xYB1hUAQxvMKUq+xgrFxw/gaSwwPe+TzWnKOO5v7kQE3Z
prwjsKZb7SF69o6rkAeOJ78Q06lrN8tnmD8HpzJOamVo+xAClAqCnaBgcqBfNHEd
I9D/Mo2Aa52cpDgnmz6ViZ7cNB4Aw+Q6j5l0VpKf0OsRQ9k92KPH1s/O0d3TiO3G
pU0F0zKUKSEnTa5xqFtgePpX7rEr/fTRs901SmeqzyqzCXzu64o23UXgnLoIm4cn
lhOT6zM2876UBiscWLh4GjHbC1JSl3pzhYKze7ZnyDUJUeR360DeC7CMK/F3xoKv
ISHBSo6Qqqj0/G8ZMLp6jQ==
`protect END_PROTECTED
