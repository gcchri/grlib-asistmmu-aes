`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TlNWDIm+UkCNq+y4JYe28OT/7oi6l/31V1FjtnrjV9oy8XDTLpcnyuk42JRyV3hy
3qNP1hYS5vMk0APi+8Tgs+X8tgJDjxZSrfoaP4tVZzniNWRhVsVslhq5ncVnBY//
4am3JCZbwl+fdUbUKnqZYMKcQTXxZcucnCVAAxy76kSsbNsIu+YaUI6jH5yT8VxY
lF6yFUzfN1PDE1tNTDEOHIGMXXPYPNMBcMfpVt8IKV1H9MOOeZcuwO1bCMcLd4Pa
kA1obfgXmwEsJXTpmstwRPOCYDUydcMx4CdCo5NZglOBKzvKI1WvZOEBvoR3RXz2
/nvAxbFaGk4TMnoJDcSP0Q==
`protect END_PROTECTED
