`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
07L1GBsLZEYP/6bdyO+UyeZcjBF/qTPqrKcBPlOdi8pohSD8XD0UCQcOLIbaGaLV
HYzLHsnpb871ELHV2XtpJOCFtOH++87G6wAziq+ytK/3b+YTAUkZo+606CqUCbcc
P6SpDU1YhRq3Pe5/uAamRiy8UdzkS3gcNtAy5yJSe77cZx+HkEWw5WkwSz+E8b7Y
hEp3un6d+Ok/xeb9neHk2KrGuYHpQ8xkQMLzXs7wI7Y3urM+u/TjbafmVtj3kobv
fiHsIDMvx0C6oMY3gh9cX3Npm89X98hzMkvrZkTzqAEFyv7TKbfnWpvqWAzc5Ml7
1fmDlacuf1FfWTOM416gmEB4bivvgEnCu1oR0jgnbDF2SCe5n657iV6HFSiIJxJh
IiIm2c3wd/brosYtRZEDAHObEVfB2uOqNILVVRA2q2mwrAXNRzXaopoLddX/9bZn
7j0vYi9yfVxFIqVN346SJ99HfSG2PBMDFkbh5eYao04V5a8F30acEhSCKEbw22Ul
IxdKBLTY0dmcJhytSXUSPR2WkxDSyEJfLTTMdvJsCzwuuDkvNHuX/xnEYoaMii4X
EXW/23ibhFbeEyNx4GPrZ6zOAcv45wLczHhR9rr8SUcSN4sGbOYNn0s2Hwd+5Lmp
XW2AeDOitLq3Ogsa7dB4lcxmqpkjfZ4DulyMBdyGF1AdWWvBtNUQMHULy1nHtoTS
1Uscu6QVyl40tAjKcazKFvATX11iSxp3Kr6Q7nEKRJzjFiVa6hzCQSvEXjzCLBkZ
4/VdXxGGTJ6PEY5XOPwFFLX/qBYDnXtJHIlM+l50WOihN4hI1MX6+TK+gjI8siEr
7y9Q9/6bWh03eu7CWLmXnz1qIsLwjiGKOloKQIDSuCudHu70McfAfi4nm8tVCTrq
WFkvfA9yqthwbpkNrdyVcmnEV/XZHX+q7eRotJHXmEPwS39gCEFcPSc9v+Cz2zB7
KJh7vIXSDlKgGlaPHaPUTYSyH6F3T/yS9E7WNk+TcwFsUk7BXXGAr8wKt3lNuF0F
aRpiU0c9g+3P318GJvEsktGU+c88OnxVG2yCf3AAUPSlzSA8WDlYtYljxT6saLu9
NrdQCBBrQZCi4XHxcLsh2sxHGJlArTMtn6TppXuzsVk9Ar1EDxkDjfliZfB21V75
dEK9GCMItgnutXYr2Py8+5TpYOrU/6wz4KIlBpm4WcPpmeULwiXkBNfZ+g9q6tvc
yxFuJP8yMTt1id75nwQXlGY9KrUfAbkYouQLO8OnPqzrhIMQqzkhMeioRB61GXnn
O8fvxVplZlGZGQiYMtWEmtPXQUUbEnG9rf+vZG/lr41ylRM0Sto3JNL0U4feCpqQ
XHY1QMtCg2MEsO+2mBri2LiAJBkarsNTInI17jJmcni5o66+oiqlcABfEVVKoWtX
LyK3yqvY61JzIdqLfthsDg30qZWUqO/6M3fA/hwPqTgCA9fLhbPxVY5foeqDS1aE
iFVNzi0Qe1QaMv94iy00+cfVKUFH8HsmFZ7updKVw16XZtBIcQwNJDZ4A8cd0k2A
1NX6TGzl+ULNWPoHWqk/fF6nxWPMdL0Qa/t5r8mJCw/ew9hrrWZ3Ai94uvSsxoRE
uQnmipEAqjx747IVKECZgFJ/4YFce3nmNhh6zvqNXXSt+Rt3b2BhZVzl/ogk0NKS
5qHYds/J8uMAgcB+J4yujNq3FbTxdPeTx64VGase3PoS+mmaGrYixdW6wfC7U6OR
qIZkLbtlUGEX0rLfHrv54ypYgaUJ2XsPAJNi794jTAwiTbwcYxbDhUjPOgSfzO8h
5p6ccdDR9arTjBcwjHIv0sVDK+DDR6rDTOSx4eOf8h2XioPNhaEgXDdMcKuAYnV7
p7OCqDRVM550RiwNYnN/59yG2tpseJxAZmhCVKNKxBoNbKZ/OavzHL0cZXFYo4jJ
yGgkGi3A/8OYPzYgvgrIKmVZjT5HoIlXPIkzqSVPAq2gCSoGizFOawoccMmWcxI2
61EyTi76JlrHGTkOHJsXX05nUdU/A854DWXN0HalVxlUlPtzbrkRQ2EO+t8Nd+Lm
uCW0lZWj40eOHVH3MGvUbYKEu/u9ecRglV46WIZpdBO7Y/VP17qhlP2VIUkiBQnK
K4yfBnepzkprfmXoluG/puqgTSBuUcGYDzqmHzjTu78GG8mi3QeRRWtDqZqC6UgD
+WCBk3ZL4NfVw2QZhix6iFyiSDaUODAzvqNl8088t/mSkEbGCNxN59+JjOIQSMzH
XrGBrPds/vXYmxvDE/lEGGmLCVJ7ZZac4A0QjYPJlOPmNzWMr5qt2WhDa4lpKJ5P
URSm8UfR3JLCRVlcoVFewOP+12yYHYTJIu1wFVhrlIA16wuvuJPQmGy59TBgSTdD
33NG91ouySxp+3ilQvvEBkv5XcTLbQEgK5YQijswJVZDrLLgZMTRPvXqX2502QKJ
5t8hoAVGUiM/V7dvol8G8gP6FKFSD2IlYK5GjgN4NbpIUkBhXiZ666VhXSSGwBp/
6R3XT+u+lp+DxV5SSZIbQh1enpJr8qnzDC89nAD4NzEB9epbM50NI83yB66YwP4n
+F2L+u4KWhz7WjYmMdaQuj+7jdeMPKwVARHslt2lsWxjEFJcecRSjPa/2LW4SSk+
mLFihdsnDi20l1OeKCOfcY+vLKfByc9CWsilPV6PEeuy4N3bChEK+DSRP6q5w9vt
DYv4FLu5byOoVSmM0sTE61cQ3N8DHw8hwYRZNTkzcyk6OoWjQsUN+cJlSSBYWMhc
KuzbLZc6wxO9QYyLhqg+bFIzOsDKNyb0liKa+q9sLE+bQhSWENTYyb6NRZ7kM05C
7jQcB3G953itNdG+jC/umo2d/z0lRdARmKEIVlpGkj/qn1vIUnDkg1j1j8RlvXav
ZLuo2DTcsF9gnCZxowvrONm6y+AlvjGsuMlpBeCCrWGjMG20OflbjESGDooKYwim
h60qjiuee2YAcKdbqMcQ77Qe+ip9g2uvjg0VdLFbbI0KlHzQjzUQ73Xtm9JoY5gr
wYkUUFPm6kBuYoyR7qBh8NDaFCe4C6bHQKKe7+rxlFxBTn3waquuRcTDagjMSYty
0kZr69qiKT2iRwAkEbRmz4Y3RP+5hPi8tgdU3ovxpjbDtVcZKH0Mq6wRdJ1Fa0ga
C8oP6PmeHpVqOAG1UT4CxANLGChkr8Xfqj7FDk+aRTHKy+3X5ZZiZdSIjcJu7xxM
DpZy6qFHwEYJJm7r4G0qZ3A21a87Zgh/p09LGfUS7pfyr89mHTH0rGzQJxjCfDrw
Y0g0tkcWtOjY42W/L5QKo+B/x51TbMNbsvzrAtmag6TzZ1ECAx6gFz3y8OHnYvTR
shisIc6G7NlpU5ehziG7xD7ItdrSL6DUyJ0QrDxumbv4nnklk0rHSR42jUzRIONE
3gdS9MiBYN91FNe18KA1JB93kxHAgK9s2Pf5EMUFmCpijqJFm1U65HPxXiwf0w4i
5LZLxBkJ9KLJSkaXRnxGHaUtYq4RXRxeTSmVs0NFM6cisuE9ixBwf3V9r1qVsyCe
UpIRgdsgQGQytVUJ4KWSQjHVRW4W9fQLYZye2OXaC5PGG2aXuiPcQEj9wF9IsH+t
X1njI4jeV32DASso2ZM9FG9G+cNTubNtk0YZRYLH+QxbTR3RQeaWdb1yf2g4XzSE
tq4SaEzB0d21dmGAaOL83evgFzQPTQqzoORBzst3Lmbvn4kL7+0iQJtnpoe0hqqe
jM9kBMBVo0qK9R5HVF7oTh3yQnL0IXEnoWEPhjJR0C/N/pS2Xy1ci7HH1SidHeqX
BFj52Rgs0gv4EickORh8NWKbYm5YuohBV53t7Yn5TUU0HrYXRN7aBtlNrK/WGkk7
GAOJDXFapJ7pxF9qr/4jSZw23dNQsyeULGDFDXWgBfOS4h05LoNk/iOOZ8gkQQ1i
rmtKmX9CjZwODdLALi1Wp4qC/zvOjxEduad3lV+vaAJAPTgj/wGjzcUJaxs9pTM/
5StL1fh6CAGMEbIUSCAy3Xx2rNqGk6dUO1QUV4nBr5zlY6S/df7yLN4Rgh3WSV1w
kgLZCO9pQNoYR802zZNCrl93FL0AFmkiS75qOGLM0g5KCiX9dbIlJCXsyStIYHNF
KZZrVrf3Uj0Ptz2GyeyiCKAU+StvJIlpEwRO39hlmpC1VMe/ph+rd79GlHpjhfzP
VihyB/yT0cYsDXeF6yTgW2R84rkSksKLHi7HhzmIIOglgfcc4xqAexIPsWogCAwV
u2PSwz/XwaWFsloaz2eCsn7asJbn+48iled7OohKm8pmdbrY3P8gFb2cnEWZUx4e
8J2wRp8KFCoAVAQbpQdCmIosbxhP2MD2MBZOaz3NTUbkMj8UXErU8MgEqJLlWUnr
wcOKaa1nXvmbVx7kspeU2CGwLyb9UB2b0hAbbGL33Lj2zHn+us5IpbyKvPkYlPlT
iYLv6kdk9939w8ZZAQbjQD+u5GS3dbmTzMT1FDnyKoJdtiJ9SvCbUKoWkFmZcMpK
Z327o6JDSvaX/PH/P/hrSi//Mmjjhf4T7+mTeO1TxAfGRmQuOO7i9CCw01+oKG9N
GRi/eoi6PxSKHaP0zX0dxw7qRTiq+viBq0Sy2FJEfQs3GbpYvizAmy0FSJ8i2LyY
cNsnbcrSMAz+MyyHwv+KrRBms1oMlarwAHK/MDOp5xAz/peQ1HHUxi0MAKpxdrZw
BJx195owoTNWAu+MjDX1Jz6xRNd2JCwakY6Chd8A9ol9TrYWL0f4pEkIkRolhlta
skyykmOAspDQOtdwvG6VEtO2qgHX2Uec9guwUsz1HCRvF222lwRG+opdVKRDyqHO
QtjjVNL2poxGZuWvS2vDGXKDZyZDy9gj33n9nUsuckv7n4j+/sxsPqa4PFNzZI7m
qLBKVi5SPkm2QP00JEM8nFfx4PjktsiixU1hEEukrHz4bw0nd1HoJNFf7IC4Drn7
CV8E8Jam7qomv3psYksuHR+rBWthkWv6Eso6YFa4quN5saOTrV5pG19DrV0C3TIo
jGbanimUyNyfWSvgBoNQ1aXFruXGd8vyiECe+xfFIIzPAOVyxlYMx6AlPbfvQ2XX
VH0gqNccMnLbcsQP05gk5eWOq+kL6Ytmy92vjf2hAunnIs08pMuLn4XEdc1oJuPz
qI9E3dC0V6EOEZiAM0jNc5wXWHH9t+R+dASqYfcUkjwwPdERESQqkw/cEzTyRjlB
E8SliNbvz++sLUiJNg0r08gvkBSoXeY2OpT9J/MLrwDFSrAAAlpDCBByJvwsDV92
TNjXqwCvt9NWO+wgresQQ+0oAjjEOTabN6vtrWxvkUkg6RJ1k9WnhQSy1+Pe5Hhs
eOnMH2F82lHduLb0Prgt9aOGE80mZeEcHY6yIFnnkvs0mMcJfvEQV/yrqBP+H2JZ
faC9bPzKJB1DvAlZVpwPzIGNUFxVb/xoV/x9wouSmn7o4Xyj/eKBFjP61UCTwDmS
`protect END_PROTECTED
