`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2eGCFQ1UJ2oRSY2ggUUN1+36lNfh4z41SvI8ksHtjpX18blFsM71c00uRBhuBhai
7x/sQ5WCpRgtqGWtY0wf7f6GvV6Xfn3B992YK6Lrl4vyjDuhv2PUERwQ/eS/Ts+f
7E/cbC6LtqFTJ4/Tg7ve4h7E2H2GnfbHZkfBE/mxSBm761DmSOzTCZMkUo+qgLdW
ImRAnIc6kHVlnMdCaYwIlxREL4D6wx+D8WkruX5fhgkwxgnR4Su6UylU/ELKG45C
+6dhKVAimlLKI5+NXt/JNe7n7JoEiq4+O3EWHvmPSPZykYayOwqCeinAlkO6KPnE
rxwwCZtgR5jwMhLHjXGy6ow8q4HmGkmEvMGx0wVxYmzOKXNSLDbbGEfcooWbgf6d
P5VTpzBVgBEJEKR025xtpaRlLylsdaUzjB+9d4k+e5+ZSFQMIDGyVgaeh1By3Une
sSvceZFwru7OukTjrKI58ObQ9c5tRvR7Mmlx4HhzEAO5pRO6vyMD4ln5E1gE/8VN
kCvuSjgDKuOjSnDQ6iEPStPJzak4Pw6yl+3Md7fdQBpDlhKoKhvdBh30Eq8OA5Iz
3LrN8YVXMIdF/vD6KhLHJhHhFTAv3j65giX1MZoOZ6xkxtS2Roy1Ymh8puA6i3Au
Up8J1cAdxJ6ALuMuKzK4OIw7UYIBdwV2hx4mTrhM362/EcxfjDDiHeOZ/zdLj5Ir
dQI20AyZMFDj71h4AKX2s1JfkTQmX+Wkse/Md/I4BOf+/aVTvxhRiEgNErmXZ4in
4hCU88tXJiJQKMNzEi/XoHVwX5H6iA5Bi+PLL6DHUrRKbRGvwMPJ51+4+rgquKcd
mgayAwfa1qApt2TwqJTOjRB9fGJuQ83Ei2LxmBbAKMw=
`protect END_PROTECTED
