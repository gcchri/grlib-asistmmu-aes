`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WG4/lD6+fQ2Fw7ZI8M4jIaPmWQc9tZ+2iorASFdUUvtQKYW/QmOJxhbmg9Y/uXbv
ygrDtlwzHFjTGrWmtTmS5cRkepCmYmaJakaSf/OqX5HykL1az8o+5Q33GyB1vEAL
RACVMxowLpv90wUT9SPkEXLa72tRYsyKW2NInCqpgVOsQvUI5ugVJscoGwY7wDMg
8zOyEw/YTfqyeMNv2snc1RfP0XbxHsmeG+//RX4/cj11W49qSoiPa5kpV8Mx4uRn
QryalZEEil7mPRReAGN3PxmIwYxp6wPiL0NBpVgblTUyM3LrFI9yizUNjJWD/WWS
86+patBgn1JrVALHm2P8I5sXvtXoOvA328UqHejRI+8K31+rbfBZixKA+7Dentf3
lO+jzvJWxMe3tiGmMO7Gz1Z4c/QfAMgHKV6x3A14uMpBPQyJ8qIBAEdNTidz0Gvm
`protect END_PROTECTED
