`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWo36j4tOSv2yrHMxIU3TH7Z0RlXMa5+3/G2i3FJ48F1/ydJuloDaiuiBaTh7fgV
o6YaCwblVeqRjVN1bSgzqF8quEcj5irLtdAxxOT4CDn43xe8VgcjIQ5rI78zGBx7
KlAIbMfqPiDotUVD7K68kwoD8cGnm20Mitu9DxImW6/j+xezmZPhbR8zdNThLf/B
8VvtnXvAu+w02RkQ8hdG+z2tQqSisgbqmPblLs2BZBIZxeIaNwgdtYJGZ4/hRq84
MzM58IdWtwzUDDLsnjDqZoN/itjQ2yHFJStgPe6de2AHjZi9tq/sbGP73xINcPLv
H88DcFI7Q0geCqjL/DiX877XSmuzLOZ+8LvS3TU/fy6x1kksthp1MIILC4k520oO
9L0b87TLfbos2cQfVRG3pRIK1oP+Xcr3hhIMYSzMoUYAFXmr7T7+4aFNTNFnjskT
mdKUic283HnoHqld5hQzeQsN42LtC6GMBmRU9V5HwqjhqEWZdULpjbuedBSDdDlk
EAFaolv2F1WvYiSrWQYGeFVC0rrdTDUMR3UFNQibh/YJW4GfF///1M+Cy5KF2G2o
FpWekGrnEcnQipYr8LgVdmTaG7rLCbwnf7835ARBXUxdx2M+PA/SN/fsVbT0+CKz
vf59EubxyxOLa6ZjkbCkwnX2YBpxBmc5n4kEz1yTY+rrfYCfNHJJ73X2qOb3N56w
nP4BNu05ELuldQxPc5C48x3xKkeniu7AKFZJyXAHewAHUOkNHvz6QHLh5offfgo/
SGsfuxJTFsv/JyKZBFqeibIqjKbh+xOnqWrwPWsegmzI1J3HOiDlmLLkAA0fxhBh
YtpjG9ch+gol7HVTA9UvDHZEfSe0TdP+I0NpNFzce8c=
`protect END_PROTECTED
