`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cEH0r5+6TM6JElm2T2Zv5YRHwnMf/r+AixXEoYYQLYxMncr1RazG5s53rlow52WE
PTy5FeKB0C2XC6wX1BqJ0cIzCQM06jcpInCwf1layUpJdwhgTtuRo0D4UQeaPYI/
s/NG6hU3PJdgVrp2Vl0QeeeTY4MyRiFGE7VkN2YZWtuDf91xwpI8AlkgD//K7MPb
9scIACp3ydxjm6jCD+tJSudNRlBKx8VLc2WfCZAxm9661WcPNUoSTs9hL89UlVuY
cPz0nUZETHM6Y2cxltYSAtsjUOA58dQGCqKwGOuT41nBpS/UbDaGTEsUYgWyC39C
YbumkJHCB4cbygNlruC+HPwhcEojWRbaXNmLbgFNCl8as+Bz6eoKNBYvQQxehHcL
jAldvFcZP950StDYWuqaP8+3vQOR3JF7A4iLTEL1/Ldrws4fe7ZJsUHJn0OWHk7S
8r+u+TdH8YxNE00zcddGDAfhGfivQ/+Wee+tpjfPRd1MyMX2mX5BDcXdWgyUGflI
TA/PFCDqgvD3wJEeqnz53cZamYbDbdDhUljHMwb7AZIW+gX0jEgTTHQ9qblKoX1Y
yMjQOF5dBURHE7eDUjBCfbFa7VPm1VAcq2QysmO135HkPadJ9zFhtQau7kmvCbPM
`protect END_PROTECTED
