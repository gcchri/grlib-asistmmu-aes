`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oQBxETGsStDHh8px1pMv0lalPsl/HWHzMzvEFkRdKYxEF04Y7QPUZPgqcODNzi2z
KwfR4eOkUo8NnOpuKDJSUi5bPOChrelCed4YZVGhsaPw1gtIJpJv97JJjSir98p2
nI+c3O7nas0cPRhMDVQ415n7NMVfQM0ghxYdvmjKOa0jTUbpN5JdEkY1b7f4C8Vr
efI4Y0h9Pi+usE3VWXNO0pOtkYWwSia3wScPgZ3cAc1o1O9J82k+a3nCLfsGxKEm
9S+ZzPYQo3ZDCsGMCRUWGxeI9Tw/ZJO3wcQRhIn4MpU+Y50mlD/88FDqXEEL5WE8
`protect END_PROTECTED
