`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xdkgRrmds8wB82xzE2+RBFEefAlQWepSkuHkIifBr084x4LyTknxmx/iCNPB9MWe
XKYspTDggRP/vcx7+Flyk2YUVphWP863C7JiVuoe7ODAaNjgYeH1QsOHjAW6xLXB
7HAZpsu/yWtcd3NFfaXSqT/rov+z/JhhZ0GLk5WhaJhVYdJBFq/RLqny0xjbFbnr
Ql2yWdhig2QojjRlB1ezJGfd45YgBTjKt5UiQcsvbbpmlxs6UqX7SLEfJq/EwK6l
t6hQLN2ojOI7ictInkWlbtD1+sm7pwUbjASlLP5+H84USbvjFvfxLCPnSY+WsEGa
YlV4Al/a0NrUY1sU9xEeOiHYkvn7f4lVNFrjYnQJKYOPLz+RKl+UP1DiPVBJlozr
C/DnAEsOKc5VVnLYK6HmZ/A+BUYT3ivxC/It0RSSgv73gRI/SpJwpKNFax8Di4sT
PfFePOXaidraztKv5pRTthtFzxzq08ajyunihDZs4IDQtjSJkzDCTQipQUqyGym5
SeftqwoWuhzEQ3MheF+N4ZR2V2IYrYlmsytauh9TaKBmnUtpdfX14CT9G01by/AC
bepxuNgS/NLUJHZMFlX0SzT2PDSRWXo8VQGlpwQxwZ6tXLCMvFOp+kRKe7pHnDa+
xh00zM+P0CFCWtxIU9qU/Hu8vUNkM9zXCIEAeyme3nm/QnUjNdUgkS2NiqymJ24J
W/7C33GyyzvqZJck+H/xXCMDUr/pAsfuRrVB08rn4J+Dm/M9iKvxcfvnjmFCxZWU
DajCOpXTP6mokI61EcUSPuD+Oo0zwPZd9MW4xA/7+oTaMcg9QFZpOB9wykY4nqWf
ARGVukUGPMd4ea9t+XjyN8bzoW1wPg4KwknDmEkHyYRH/ODqAkhZn1/Vd2LA9zYp
HqADaZzNnVDNeZ/F05+ysIR3Qhkxt6K0j74x6TnlIIZCSN1M56XbcuC+WHHn6dba
BTmm/whyfawg82K5pH/l4uZRmvqeGSBtD4DoWoYAB0flxvqF24zyy0cvXx3sWmKq
VDqoH1wKcB7B8Ms/N1/FkxgNNwtzsWfplBlYq5FjCrUs/EOG1TMaDxLbeLi9b7Eh
NJMbPHe7GCsjmhqARAh6pQ9DmGQUDerHuOra9Gm5WOlUReZkAa8EIWqutPiKmcCY
4ev7v7caytiFKOMJjzW5LzKuj5AGP5+W1ns+RnlDHlV4P+MAJNzc0khCRT4CJf7b
`protect END_PROTECTED
