`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dl9FkQ2ffoDpOHjq8TTeDG3LicDiPtiwpIourIY68yY2cFhObrqJNzk19igpGnnT
WteJBM6hjXvIFPY9fb7xAjK4k3QPcIY5XaMK2HKzZBByzmzdyQKgWubYZIpWk7vY
Jp28a0DL9yYIKE1clvzH8nUCfA9LsDY5uh6V3y9TDiZYhErEMcrvnJYl5tnNnZMA
H9S/1wP+UHf4n447Jz1iMFnc9BpXtyxRcSzV/Rzpe0pnxigIPHUXTCiqQ/spmeVs
6xLqezDi2seujH+rKEYnDT4oKlJPSp7YMyR2zhtE1Gfm/PALYAJXPj08Oq05UfC2
aqhedCRaeGX2i6+SHl2EE0NI9F6xmd6JLPvb53JhNzZcssyIZCWRc1ZdP31/ON7W
+ffvylDqVyNgmTzbBVNqTJfcpqoClDY5YeGDRsgvWMNN3GEFFNw7nRlqzdhTibBx
eZ/fiZ9vjAjS4eFOyGncAu019NVfVdj3N+mxNuLP1/v5ty031Od+uXDyaLobNO73
v+3OyFKLGngPym6VdvtZ+Q1pSn0b8n5j8dNprTesQxCnFtfkVfFfNWGyT/w2Z1V0
+E/dHVzpamgjTBPl61h5y1SZrPh2rNsI5wvSVhmwDiecbPXC0tVTrlPUW0Ow6/2A
YdYFMzLJ3E2zz1A/4uC+mgEkgETc5/DnIpTW5zLwERtCmOmi1Fej9GUPrvOmpUpZ
wc2Kpv6qobbGV3fZbPTm2VQSHyK+cr9VcH/+O0AtzFLeVfwTBOptyV4MbEY6oPk5
T0v2miX9csVWWatPSbM36g==
`protect END_PROTECTED
