`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R3wGCwD3eoZaBeTg4CnbDfsRzR8XzBuyqwxgBY88n1d5XBuWLTS32YMU2DEygCsY
7dG16KHBie1Um5pK4xzoe8TcR/QDzoKP4fpIuDS4FQYkdWjvlfnoLxSDaTNg0nue
FToXYREorwD+KTn1uUNeJMO+Ysy9yFrVu9TeDvaFVMAwNJ+uvL9q9dZDGsaNQaya
/HKRI6Oc/gw0YsIQhNPgsH5KM3AUVkdarmkI5kjBBk0Hly/YwX4ClB3nIo6pykat
gKRW3kMcmUpx3zDp3YCOujzubgJj3KWOb5yrBEqqXt2AZh8XwWqisWNhLRXNR+A8
DOOi561LixrzPei/yENMxpaCryvopaab5yJVLGs4w/s/2IIJ9asf/gJcn9N1a7bz
KIEsGysPvkmWRJEt58E1wX21dJf+V9oPFvqjWfqR+edAnpRnZvZ1y+0iBG1fuxBE
PXwHubak0XZflEzD8J6RW6zf74iJLKifEdQJgzSWjBYhewBqj8D8WaTInbecfeyi
N07SddcyC0Ovj15U5tR+ovEC+6S4AyJ9esHlbLByatNX8Vu1vo4LrpiNrA0Rmv8b
Y6UKsgd5GLAi7UPFUuYYUmjfmD4dFo7FGGHSDIqNz/46hmVmuaK4AFrX0oDek+cI
CoB4ln2zCMScuFueZGx8IulF7tWnxKEEHS5XOSnLAtof4nytpswUI1dx137/pANZ
ZgXCUdVtDrOV+86op5zoKvcKP6c1bJ0D9nVVEfxe1GI+kf9YgKAQZY0eY8zYTv/f
VwAkSNvOQdsbwGWsBqGxIAOOeJ+Vmo/Zf+6VWpDCmfc19B3H4kTVeRM9+GCwp19z
JOvwA+p4NvR6PGPVkObpYTK+pvFu4NzmaNpqF+kejpVXj3PmX7W2Td6+VESVZ+IF
jMBcdD75yWjFxtWLJS4vbQ8fJnlOItai1LFKrz2gtJ/JY3YNYnRVrivO/ztXld9v
A8PACRHUI0RQhmBdjjQA61uZTrxxswXhy0z1fBVo051o07bMuBB2aP6s8AhdmPaW
sHmnLaB257ZD8qfCp1fyW8HcyKZi2bRrw6LVsEq0DnTgpWF3NB0XRvhzcDNuOsNC
JMPPkffCcc/xn+mUY+TlcQ8bG98jHY09FEPV5Hs0YOi+Zq4OqY+LAGjwwKC5Mv35
kuwDhj5UXGzxH8kxUNZgZ2npigI5UBffFa88dYtVvrpoe9zoxhyzfZsXkAdKDT5K
wymTxN5WFhsY3KoIFR86JWKHIZF91ki9t+VJEpz4VsbIP3Q3tDIFJ09WOzvqyXmd
HRhUy5LF9JMQTfk8ssf9TeXwp09s4sBF/aDH8x77B3R2ebCHhCuGrTo6fNtqCizB
xhi0wDx33fAYRyR4WKdM3dTVL9phwn0E5e6RItuI9Q+sDPQXC/5AYwmkfH2NL6Eh
4RMSKUqQJgKFWN+1MPHK3hcUvaeVUbSPiFAtV5hb3XKf6q9WghX18Uih2/8YUWbp
mooscUBlU2eGCi5cEoB8DHlFaR8Y4kZkCuD/FYUtIRSPrVcnjupg2e6xNqFVV4/N
rhuoRXkjQYzKwlGSxzreUkHxb+cwCQpmy2fl6dZU1P3QkuvlLOkp4R1JELGiuuya
m5k7Hx3KfR72IwYY9DxeG4nRkFp2LKzscNgKa7H6JJm2ER5OWl1k2zwa5fNsrFLU
np68+t52DO+R/SyhyjzA6erkpugjbasaxl2RFV/8Hm+XU4LFTzDTo4LvjP89emMn
2u+A1MufzHn+hkgDgTqRnfFVcWFMe1qoY1nygCyL678bhulehX3Vd13QVZbOHadi
diBNS9dzKZaEemzbGIwomExbccWFx5gxt+bSqfYgZb6CRB94bb3NhWedo1+1oAWs
5/bqxC8afHiKIqx+tq/F5a1sdQQjqXz1I3koLG8o1B+I9uzo/SMJ0hpqC108wHcb
uXEu51ZuwD68Sb3SzRFo6FzEyRmjy5O5P5ZYiLgvz0jDYKGHM3ducRJNnfhbdVEw
DaBMO0+/ZSqmVX5OQG/pLo9oUwsF1AtRbqOz4sQVC5skXcJ8KKpg8iyRhFhwZuJp
Fqtg9k9YUB7b/0ZcTD4ZijnEKIokTioLnmFBNhDnEHgp3UZqvi6RckkH/HQDFkbg
OVnbIVVay6wqKfOBowUT5hVX1r3Uf/ym6PEqiikZbb/7uWJUnlYCy2nZswBiJ3Bq
NHxCODM0gErtHSFvn4Ws/98qK4nM5xjvC9SD69wdoAoC8LNEM+6gvRPLPEf99iNU
Q7JpMEaYU0NnI+/XdTMwJ+m5B8oYGo1+jmOYtXFevohClebd2iY96FVsWibmY27h
KLu5smE3j8zwgTMVYFupnrKD9O+jDsnqpMdT93xkRRFO0KjqV0ZnxZcKvIuESChV
U/Yi0IPoYWUNuw5u+TXmBAlinTXOihlPdUc7Xlg8EBQbWjcz8FOdYWjkg/Qx7DYV
7Oxhq5y2vJIjrtz7RWbydhiFJNzrp5YCGkQRI4o+hYTMAGhLEVkkdaJJm85WZK62
mgk/1lFVaHmkdONjRDZA8enMsSp8RbeSHhWg84YyXZJtXkrwkLMQjAT0YEBMlapo
7KoiBjZ/jJcEqLE/BMluzg4ny4tJ8VbzYh9gjjGcxIRbsCzFDICyNzWZ8Wem0trn
cuqPs9K1n9rVZyoAY0lpHrNEA4eEyZmv10B6e5FepsALzf45qIPScklXPIdad0F6
xOfNS25HFuutrZpRWjRFAQX9v+1aWCwY3/rNbA3pzG6ipKjanEyYKEjOigzfLpxz
gA9PeT5XKwQdkuBKFRUUOnYS3oinPe4kHpNwLxWWo6jI31ILMpOnd/srZOlmQMD2
XbtdGo2zEWA/5rlHvB8cwzb+iMkyTe8ThhaZcpjuTNGsuMj9c+wNlmydY7U54O1b
6zmh84o/jRUMI14RupbfHhDgQPm1uASY76Cm8zRdShlT/74Qn4UbOgkF5hlu9Jar
SdLldTYsO7FbSSZCXT3etzWb4HmxjtNjVjJj3HBatFRDr4pAe5Rl/s3WUOGTQeVP
XK1gHBhDVQ1HngIri9cKfUjlzP482/HGlxbSwtzjc21MDyCx9fckb8E3RTG38VPF
P45mUg3AXOv4x9uaUc+d0MSndKp31BiPRQ2cz3D/ErQDLCBFbEIZCUIwRCyxaAR2
/rusx1wI1tGl23QuzPJSXzT5CiBDeIikoMs9+oBPBsrTpe13kzBBlNayJmyWholc
q25ljwicp3UwUmOe1PFlFdvvN80tf0GGys2j8VP6hFqxgs8wy2mj/D3UbBj5nqkr
dF94UZxfRGZqyIvU0pobOqizertHYq6cSjUxq8yb7rM2dp5VB6XhknHO9amNbdPq
CEJAdO9tQELQNy14N0RkCLkYyDrjB3rwfOBIxra/aMghmen1SPOqfviTag9LQEWK
mU+BPEgEUgMM+mH99cs5KQ0JBLEKnJblF7I3YrOLYztauas5vIZqjZ4KgO9lqxOK
Ae6RK9dg4TgNwrTNgqJD6sgt4d/dxyzOzpaANU/RCWY2QgPTS8So1PSg6khFgp6Y
Xs/+z6dBnlgeNNY484sPa7SCF+hCb9iZgNoDspWjfYRwHyUd6QMEvr8gnIfIJitd
Jf3HYAEPSPSoO48ddCOOPVbFgW0f5NOqSCqa00jcTlTLNqs+zWJPfMfX2d4PhepL
DkJzXNdw+xbIRYRgWZunlofigunySExGojBrVh9ho1/d1LblcilAAUaynHpctDyZ
uYxcl8PtFw+s9a6kN1Pl1YrHkTaeiZRHsLYmCBCR3GU1dokk14twc1cuhv+Mc6UD
yICnMFgxv9XZy6ZefeN4j8wjM1U2SNX3BNWsZ6Qk48an4Pt7kV8igWgYTOonlNpG
td/wpAKLC4KQ1l4DMbNWqF6aTWR+gacgOTMXu6G7pHtjlsmfivYo1kvHs2JO5sgY
3gyjgujm3UWO2A6ZWZoSls63BouXKJX0LyQSaYet883LiCaUsy3/kZzuJ0SxrzDi
eVZ2UHZ7oqUnL5eZ0MTkz4133lmtj1bYHfpxwH6gc62u4MRmos1nw0/zGYrmQ9ej
xoj0fvjPkjD0S2AxhjoL2hwXcbjo0PD+bDh75k5Fqq8rVhHSl/zvJZZYwmkUODjt
HTgiNbntSkJaEi33Uiy0eGEfOKo7ay/ePDMau6TEXXD2LyEReHV3z+Q7ZU72z+8w
T/jcQZLn1tTTGeXGx3aPQgycgpucZphwWWyXgzoTs7F4vxml8XGIjahaiW8Sbd8Z
/izvLBUw3THJDtz99bR0wfVvqUBK1VnqFDejVbFY7yg0puksVxWuOH/ExOwAvU3M
A5J4GI1X6KklDNwwipqPuVbBJ/eN3MFFjw+HCS0vSyllQxUAVlnnat3hOQ7BGNxf
SNVhnuZ1arLgoLcojxi95pUxSruZ9FpyMh1xCZ4aIeP2yOherBOYR9G6A9KB2PNZ
JLFdnm4TM1MuVqjXToHl+w37kT5IETuxsUICkUpd+EcGbSY6qPN1fJh5uTK05VQZ
6Po71Ij/N9c9sWRy0nN1VetMbb7ND3YplHcTXMJsIeehonLGG4ftUPrSqEDEgVIv
QRIHil6fyY6Y8ypyH+phIj7VfMxuTI8STl2yOCJwiSCKNs0Aqs2k4RBxWVupgTjL
xFHGvvTOeVm5b1Mj0c7dkRziN3E1lqyXwoXiDUWBf38GC3FhKT1tP6ay/Vqi4HCc
EhRliwxW4xROctxOcG/C6sC3ymJaG0tUQ0ZUtv2ZJsCOLfoDEXdbKtJpHGkngi8C
yhfBkmuDQcFVTkb8+gnsMXyNozzdl8JvJraDpTB79nq5q3nL2a82y4RIKnP822ie
9f1rWiKhe6++C+uERkKQcqkBrT39kSjfeoA2fxWaMPb2bFnSFd1LVy4aZzaefiMi
6LPykCfzbeLxhlNa6cVZny/ENGPWqGX0Q7Jn/Qw5Kbyz6hUni2rpqhtR7vyBpFGt
VzBPE3QJQ0o/77q7Jt/c66T7ZioYi5PyFyb9sFB1w+qtIp+e7jVBKdyHdAYf7GQT
aj6TaWPZ3zOD7ma4VdRsmTwQOhRQ3rFFMGd6Gx04yQJqy3tAskjSAHLrf3T+RvJD
vPfoPpB5s98zShlYTleqgRWaZvF7nn6c3SIwBQXI6PgzBVY1S7LmmGi2BEAkJ6Wy
4Va4XzSH9CEldRfoSnhQyZUSmPfu3Jh8h5TndSxE2crCvnqKFAeKtcacAvhIPwp7
T0KM8BuS2gE5WbiWzQIPKwtIPyl2OHBFxZo7zfcp8P6GiBUr2jpXyBx801qAl2NK
vvzjqcOZf4C2dxqiRShY9Vpyk8EWExr8RInRJl7GXxBCYKKV+dEtw2e/VnSa8Qp+
KvxyiPeyRVgHrqV7vjo0AMLSZOkTKu4q1GWerlj3hrIi5sz8OSxwktgFmIN5C41C
ipDpFmYralnyiDuSlDZhMcgBE+jZDUETk/TKjr6yCy8V0Ywcz68vfh22Bh8Gquzd
HQ7bSR/Cab/DtZOqbJcJSNa86WPKbUjAQKhQu9jRLA0vCbQ0YqNiZS+R6BoL/dd8
/uVqOJ3FtITi2iWgeIx0z7lEXqVXfGjDLAIdu/HLlUOLwyQHBbr8tfnhOztZ6MIz
ImKQR9UxALlzOmds5b+S5opfTr0G+6s8TgF6NHABtHF0ICSEcJ0x3+OWHy7Z5Qv5
53rzcwYeLaLMSzeHqSXOTKGpiTK+kFD5zt+8FEiimTZZJbcvuYvkR3cCM+teUDXx
fMJ3shbOuCnEYtDL3q5W41DISUr33X9F9Z25p5ARnrrSS1OIvqYsAWaTrlQkHIdL
AznBNEbxvEimyD1IDpPtsQN1I3ULPHzEHXEpJLRtfdZmk6rcG0YkTQMpMBpKbMG1
5m1FLoZzoN8qlkIQuX0sPJjS4ggX2iQ4JXXhPXgU3oDoxe6rOgkZyIO36/6dpHmV
gGAnqbFH1gQLQkImzCTAv64CGbnszBvVOG7RyAWXPnwqvz3m19TV3h0TtqY7nPPl
TVOmvCZ3Q0jyGkLLx64ylw==
`protect END_PROTECTED
