`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HoDi2n92xaSGsMc4v7Rh8AnuesJpw6wrm9/jVn7KS4fafM018cj9INr5sCF1gbjq
ReBmM+G2RNANj/2tpaKomuDlLKt5SPE7UB7Z1Kq8qQUi/3hdui5+NIeTPJIF6xuM
4bD5RYNkTqw1TYvCSNm7+La7dqGinNsFPEH3zjFjsEqOAueE5Dash0JHQJvuBFtE
0ADUpOvb2xp9w/dIS4vkinSlBlYSLWcvCm2E2RGYeQdgP1FVYN2puOKoZvcHxllG
tzWK2uWMBQFQ40khE6g760kwlxFli9e+I4otfgoRH83aMTiZfpGkYMkQEeJkMNi+
GR4b6HHGuNEsgdbvS3hpyeDhiqBkxxamtQ4fu5eXzxi1/hxre+9P2XxMr8UNFrjN
66AqWWESnOpQPVvmXBS6CwgGfxeLkBejanjO+NL9IS9cSUsU5mXQCGwtZJ68lYz2
4TIwZUR6s4hRn8YqrHMumfqLIK+Wxp8jT/0GWFV9ot70Q0QlhjtwPDxpdFKVF/rK
hIs6KOCD9BFudvSZgfCxhkmNL0yJj+H6TX1jFcF69k9gFJpFWVJU9p1+vLMKf/XQ
JrBBRIB+J97Zb/Vvj2aV2dUBmbVL1sI1oFzMWyTEORW/u9sIETvNLS6lci6G92h+
PPFkhQMsSJYda5z1hJxccg==
`protect END_PROTECTED
