`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/IGycc0+0lx1RLxLhDGMM+5lZdm+wT+i571uaQNE0S195GBXpTvCDCCxEuBXJrqd
EhDNM3E1z/BeFh2CGjZKpMd6nN/H4mv/45usvDEh6jdFqRhp15VgFrmDYofkXHIc
8Xeo3r/gs5Szx+x10WYUh1S8kiqJDdjHlUMJ8LB2zhh4gJLcXOQSJ7UwbF+KCOnz
9JsDarEFJpogKcmspiS1HuV63gYF+yI56rwI0ypEoLXHGwa2YuUJqHQ/53c4Fh6F
sbfLfBp36GWaQEFd+WRSRx9LB0WQsJo3BjJ/csx2n7Q9oO1Fv5Gtt0hoYtlnceHh
3KZUmVvwVc47n3wdK40G931cTZQoj6uMEqwaJN9KZTz5LUOlwIgYr/N7EiIfCVXi
PZcIird5F3eyBsneNhKTAkVIERfzKp+5UPpmLTsHVmNvt9DXmQb9tuht1IwFK6oa
`protect END_PROTECTED
