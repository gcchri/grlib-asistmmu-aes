`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RHZq9zugsxQxZzrMc0VdcT/SumAnWqsQL87PuyhAqSL1crpu8tWFK6HvxrXMxnmU
c9QawK+xYmj8eqEPK3vN6NiHw1zF0LvepTRaG8Bz8JIHZ6YlGEWY/d0rJbBAIUWF
e4GA/RHw9vh7yMJ1VANVomDJiy+01pEoPHNq6LOSGri/W68KOjPvBjaV7bGWTWht
qu05qcxzCKQ2kF1+H2W6k627OnjNtjhxNHCF1CzElXcZvzx9LKrXVrrF6r8YATFc
djltTxip/+W+JDXlQetacIHlgCYK4FYIU09ZxEIhBKuCmwoH3Urd7IyPIcKBvhBg
X8gpBQEu45GpY+6lukiuK/QcCleGSggCSs00J6uyLdkhPXUEfelb2YUEB1ati2iY
xk/kwv8w45d60WkUtDSZ8HErx/t0ljoTuoOeQzaViy3glp1z3gf6gJRLk7wZGBhD
`protect END_PROTECTED
