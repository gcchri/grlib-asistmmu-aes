`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAhakg1pqJuHtiklJNUCuwWNiI6jP7jcEf341lYp9eucvOBkCyLl4r6BVhdNQA7C
tLuFWBBNOiBfev6TJLK5Xs9El6scNTQy8uwJJc05R/E8+lwRV3wpCFCv5vYYL+X5
BfmO829Z/k2obL3j/Otldb7aPSuXsh2ewZyhFlbTiIIfbO1qJhTiPwoEDD831ZgU
/J4RqxF99FZcwC6rCQEsKLD6lxGgk0ryF/7UMQhXP4/0brcarHPaX3GKLLd8szJf
Aunj41qVkHWV29+zVU4Ie7Oz3WcJNgKHPzMmvKNLcCHhWc0D25NiD0eT25+DUrRF
CfKgZGbB3RvJ8S2NKb58A6cDy1KpTOkgDGBG5Kvs3fGIlHR6TUVrXCghROHOWYkL
7pn2ky/ulweYIQl3lFjLfLrDfq2G/oMLQ7V+8bpSksY52SRc9zm+YL88GtXHj6TX
6b6af8c8Lw3W7fgHsc5Gk/eD0kgwnlKb58dh7p8YRUree40OwL8A45+r+hY5yHmz
`protect END_PROTECTED
