`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qutTkd2S1OiBmZ3RzVxELiS3n30SXO49t590McNYbDcUirHQIiWXJMtgMtZkHcNH
hN6IT1XNCX7uRaMT8/8D45snLH4OK9Z1WDfSsOmZ4Huv3c6GDYdyxoesEEaNVzP7
/u9s51LBQXzKh35VZGXENmup3H/21XATr216KCJCdc/ZhMAlI9r0x6WZK4lQjYYn
i4Ha0UbcX5jBRAv03dm/GTfdgJuQLUz6+JzZfZQlNgkf450brzv65wjee2XJpBdO
Wgvi1gEnSFwMKwqD/vP/jDraCL4Yxt4mSX76b3gFEeyWU5EsYfvt92uhZgIdn76V
nxAOIZQlkAUbhugExazUu3ORC444MFcgwsWovILu5KA8CX9p0emaZiPiLUAg4Okn
L3P/Ug6MaVqXAO6Sg0m2tmJcb37XtPuJL8SW+OPmyYLHFjVqLks2cboxn5G0STMr
CFMIJU41ZpKPvcFT2xTAY+TgnuOblAQUlfi6DdQcL8DL7kr9vLUrgjxPSTm+TXig
8qcKHpbNBUEqexgmrgYwjxWmCUjiKxQzg4hadfGD2RI6rWWStyeW9MY6oSTqtHb1
lnY10OhX4XfpSCIsqONWnciUlui36XwQVkcgBKZO3NcovZSezhR6iTp1ValzpV0n
rh+1Qj6sUngiylzZwlLVdOJtmF0kDQ54pnkG2PNEepjjO0R3kRIXfYHJbBI32EPJ
D7M68i4Yl1mPIkAyrts8EQ==
`protect END_PROTECTED
