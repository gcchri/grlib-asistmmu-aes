`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIv4iUuDR7752MzDFrtFxu+KzDCzbTQIfmkEcQjXhuE20DqpBQfOEWpnLlFBbq4D
g1OuLWzldA3oDzGlkE7eawaT4BF0naCnPlaxunVc+3sEo6eEiAkwVXZgu4GG02bJ
yu56Um7Nv4mNYwr06tA3u5sLx6Z/8tomfRh8fz8cDiLrEkPt3U3qdfD7HZfDStrR
IX0Wh9kLTRJ5TB4r+o6BRVFLwKUxIjllzWRaqHlg8mPtLMpx3LaqgCXEno+THXvp
BseqpHZkStzCB8T+vBUI2NDgNPXjsdfolPP2EL/+fLQza4aormGf4x0GlaKdwrbd
dJXT49Mu4d67/0WkzYdUMEfk+5QtEbNPjgag6EVIvIltyB15b6JzchmiEVjhsIeU
w1+NcVqPxnUVpQKMnU0wkkr3mTvxrgKmp6MOD7lN8Q2RW4eOfLp9yXN5o3cxWT2C
pwBoHR5ePrfvrW0sRWadR7s+RJUS8joc9V2vaZrOBNWocc54feCSdlcfuPeefV2J
D4q8HrxOO0LS9XeK34Vi2lVlkVdc2yxWge7LWRYJP9H2+RdIKbPv9UsnJvfTqPpv
4TkVQG14/KOjvq2WfBADu/HbgmaVvdjmBHIZ/lKG6eF3xpfFFkPYsEvY5ayAkdvd
s0kqK0r9lTFxdL61mbpxx4Kxuk/bu276o8GxysrAQEhCI26A9C1d+d6jYUKSm2tz
r7kt1pUmNSqnMbDFi9To+I6xQj6vIJC0wuiQOLdnmuLVBwINGED1c05jmDysZWbv
TV5Y+Mz+zRCRAq58gI5jYw==
`protect END_PROTECTED
