`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NW0/b6MVmRs9qMFXLHO2iQ1a3T8rgt7/w7fRYhos7Q+8GCstwf8YUxhlZxevNk1k
9oY9O+bJ0TIMcB3GL0s0GAm10F8iHQaZFRB70jiAm4JMrWB50h/CqpUF8t9EuSl1
fWLy0VevaBTJUOvg6x1+z8US88Ar5VILjRPBv6WXHue7KvciOEGF6YjlTguyoubm
GVVXDACtctQVVb1UXo52LQ81FqJKd55TGt5MPp8xhYk38Ae/CF1vtk9LDtiNCW4N
GEeFR75jGCwe7nb1jNVVFHFtRINdKCsZJvfbkNMthP11h+v3kI+WedOwvTjKkHhh
KvZXbsPACd9XL4kfOeWULJBYvIpf9M5rO7kuBWSLO2l2FKe0IUICvPXsGiGRtJG3
Qtm1lyeqYTngwhJcWnVFaW1MiNqPFRzsnJ2s5Hch3HSPgPyxT21aqlRRKe1PGfJY
KQYGkji43QcTI1i7NWFnbt8j+5zssC5WaMlMyftmbqOVdSg0b3cLxNC7AIwbcjuo
9l84tLRq6zhG4iUcvsgnEXM9z9z3j1ZdxK+v8boxEDnGdoOhnqvlPofO3pa0GrYH
oFqftZleKbcCXyMIO0Ha6TPN96lDVB1vc2WGLF2rQcJNdImTE4+Bc4y5dsw4EsOy
txvjPPL0CsGAV2zj+m2cfQvPxjEgIP/XHdkWbJiVISvXhjrILSobyRFTfbdwuZKX
V8bCN6pfKvQfNDdgaHAlzIyrPFSn87A+f7pBZSJD1AjZFycJacegKsaHdryIamds
uHHsBPPCm9oVXzBGYn4e3pM2beoh9HpM62UWR7cJJA02HdPnY/ftB5XpPsEqqEU4
FNTfzPgy0cdN9v5wPI5ygnLmfLMrQzkjtybIFl8JxNSyfdnfOq0bm7ZfefmCWfsY
hMWg1OVbH7ZDhmsG5ImY+bsiZ9VE+AzRvfiFXtijszXfpNb4yEs8OK6CGO708kRs
jHjZQ4wFMweLnjzgVEA41HAeT9rTzn7bBE/5n8TXOZRDvP2iG+Ou/zossXnwSXOc
37VNHikxsWUOaMdvB2O1/t0Ek1qjxMomylNIwvDap5gnPYdRr3LhCy+RG39jT4af
RxCbRV5MIr2qxEkB8yN9o0YThDjs1OOG6BTg4DAx4ICfuOmVc0IBdk7G+cx42HXA
cEkviHPZQezFlVH9relI8meeSDkem2Qs/mCrY4ye9jQXQDQItYvtko5gozb7Xgro
tmywLncxNy/pdbCcTXbipJsxKSqEbVJqaHt6SRc2Pwt6I0zXOwcIHFDdS8/UUO3U
QMWbwAFAFdrO0I9joJq3IVqfIBk6QmXCgmnCUydM7Ay9uslEEQaPzohhy0JmfkA8
SARSGSWSqEKaep1FIRpu4WMJRyjoKNKtbesmCdMozGKNRcBAwsB5EvMUCWcE5ykq
hhAkD5nkngoST2fRRjcy0pI6s+An6uxIG6/bx7L82gGOmmEJWUM2JUfuCgObFk1i
wjfwo2c26lhBn6GcFXtWebHHnKm38RcjQtDUuYKsPleNda8sUuELanNV3F3M1ZXp
uZj1hia8x/24LiFr6HsIL7s7bdeRVyWTIaPpM1OUkH2j9XcrjvJwyBxxSwoBFTAD
4+GRQ89dc1Wx3nOgRnIqAAehpBK+kPnAjxUvL16LCODi900PpnvDZ4MlpUT5j5wN
eERWWVC1552lHci37WntpptiDiOqst7M98Xlj88OmN7J+swd+C3q04Aqws275iS/
HiXbhV4JeIW9xTpgUKWCtl4RyNTds1WnhEVmxd8eXSFHDuy6eULHbh5//Rp4ulQ0
PPG/62EfTt6O2nqSPxZKyb3yvC2CVZB/r0hwJ7mbk5o/RM1uLFGJMkejxvrkt0eh
ASD95NzA47Ll1iimNl/epHvO0HF+V6M8jBoG4X2AkPvv30L4/TUcvvHCX/ycJ5fa
l1ZGTp00cKx0Kwc+6H0n9kVWYu/h65QsLw56ohSh8As85CCGQmVkSJexbWZQqw6w
NgKFevRGmpx3Ggl6tr8tvZKyl8+W10A6KIAezpFEl2r+QpCL6ok8/JIHHyH6y2M8
OsmjpWU0ciH0AbVKoH20W8SLGHRNH7y/icKMtQnm39w4jd3eL/QH2jjI2GWL1Cwx
2Asfw0cixWMUEZyH42Pspj4oaGu20XtmE6kYtcydZUGBZH95HxsV136VMho2UHWJ
OgIe2gXpjR20guBMTychaaDRCyOC38dBQ/TB7WNR40OZ/ES/uSmwz+LtijoiTTqw
y+S8Vzraqszvg8nKgPkaJfuQAMvUfCOLBxFPazOZbUjPmX6LxmaOJzr0ATdYwO7s
cFwIIEOxiTZfxPojLtOtX3cf+CyHkm+ydAV7dnUZAYeqUfERgbEYEtC13XbFCw2O
hFPCy1Ze2Z3Tz+PhiN+iOdAcLfdzScUht4VuAiT/NAy/3snN+FjCvW3fzUKFtHsP
fiRi7Ao11Vmiye92sql1jJAJyA8/wUfN70iM51E+4NagdjdzrudxG5KtJeDQSW8T
Az+8uDZJANXek4PFRw6RiQcUHNDCijg14gHsmZ40U01Huz+G/Fh7IIuOFe9WWrDA
P5Wq6YdJ6OddYvHY5H6uAmE7/LfCgtxMJtWLNtaTWA6Lly+lQVEulhAYkXAYtkAG
fqTEXnQ7c7ldDNx/ngEJN19VSabXhWP69S0ok8wxIs5eA0jeEv22vyDr0sTBYDi4
JklgqgRpbR5Uh/xMQV4pvaU6pGaiypF/KPSKG6Rm4YTFqUIHLhKyuMKFiJzzd6fU
1zDmeu5IIlgjVNNLKQEAdq4IBdmzxglOke2EjX8bhMLFWReKnGSpXkNaMUUUkWTE
nls3SPS/BZnkXS/1ad/GKYQv96mYiX8jRdETulhPdhH2xkS3P148Tms88C35qYzu
cC01NuZk1gU37iOsZKjwEmX3si157M/kh9tPuBTgd/Kvee/G9CBSwXCTBW1rXa1v
RhTOpYquYIagZtr7RtNSrVAFBSCsRt+n7QtgEUx46tzFeppoGecvwQSZIEc/yKKR
dLkGosZ7pGuv0q5cy9Y54ptB3QFoX22hERJ7qCnTxQNHJisKAdghQFqZfZ5uHTkX
SwHxqHG9GAsi01o9e+2AbsEb+OnhSw7KEthq6QqDV6NwQKAt7Q6YFph11wEb9XwR
YYm7I2pHG8b2XyyOZmBgA60nuS2Cwdf4SGWPo1mfhfurMIQsmjyqbsIQ90lFACfS
bbO6MWowSPZw/NAdZEtjpRzeCJEbGO7xESKMHVTfSp+Ftte3RUQcMptaXALNHsuJ
6wQGpQm2VRXXYAxf3v6PtA+SvFsC72xg7Y9OSeGObeP7D28YbCF4gfT/oeCL5naj
L/w+FVZeyHGeYe2CO3wD37P592j2g4SveC+iBGJJFGtxb2pMRMWKtZ69ccbdwHGp
77r95FTzaUmU6+3b3qqxF35+nGqdayp7FY5NLOGZJj4xca3TYEIcBOwjWeH1bZ1k
y5hRV/Rp/E8f20axgBSRbo2P7/kQiTNa1kjs5gj3f4a5/zlBpjOjgtR9DI29OKuK
uygiOFyz4eB3V8sOiBDh4ubeYue9Cd12FsB0M3wwhkcUcoVKHT1gRrQE9J27lZgn
dOJlQxcysF18a/3JD7xbPXkrXhlQUoweIPQxU4L3PROa65U6XsRlN0680nWa4CFb
CYqrw67Qk/2Kw76NLUGymuiRlNOW55idYrtlFWZmH4xYgTM7QkDySeyLWT/VTqoG
IHLI2seQ0mKp6ICL/gZbCA8+ucqsD8J6sj9FOHqp1rC7bU6hqn49O3HfNgCA273P
7wYilJdcsxjzorKA6DtnQT1C1zvYCg7XN63OEaeYqL9SS4xU5RlcxowEvHVIVNcs
6UEIIhKZYAc5nx6Qrt9XzCRTNy59+Iy3zz0bUXM2q+loXBjIWPE8bW364MMK8vAi
qWC5fTfmDxiowp+FpiDbizf/1LGmQ9olLxkNT4+WRyrmBwoJF1GWGFbzUukb3OxX
jTPo3Mu9HXX5vUHgfBarPOEKYbiWCG6yZO//pjVVRHpVgEnQWUljuwUyMrLbGudH
BMW9PyiVLnPKkOAWQ3HBZuDczt9uN69mcxuBeV/pbdyGuAd+YczJE8QIpLuYgERQ
qrMV8iwc5VxMsJYqBkBr6NujFcIYAXRebd6skTFEdo0=
`protect END_PROTECTED
