`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lrKibKxMfq0WGwCRzMEyWN0fd2DeqvNaeTR+org9T7cl2NnaT7LMB/y6WfAs4U8p
udgV+ZWNFYtMmY3KVQhoexoFPY1Fz7uF69wTADboli/rf1D34j+hKARtHznZlYJS
usLvfznls5QRaMjMPCA6zp6Lw3u96j6uj/ibCed97tB2jIzoWdacNxLSaTbN7J83
rXsPJ0n6VgJnDqyrgTllVrYzwRXhncQDuxtBpAMejR0jKPyIutIvgMc4nCgLbb8x
8K3Z+n4ErfEkL2M0PeNswzF3Grv/eMEi4xZu272GDH08AYLdUxmZgP1IRg0xww3T
IarBxMwr251gdVWF4TeFm8NVWto5/1rQspFY/gcx2/gBi2lfNTy7LrxHGMZMljd2
TQTc/qCdeR6StFY6Uw3T7ycHD4c9I3iZaTySFs7/YM5u5nOLhcsBNxprwFYZ18nU
sWf9lccspWsXGi6yuybu6PEVOFRMR8pb077V2BEVM9AH6Ivsk+PpCL+BK7mUfd9f
FBpSZEEinER/8cnv0qIlDXmzFBP3WEhBj8Jcdzq6jaOtTKAYgN6XFvdc4AQNdlnD
rQ2CIhqiVTI/2vzJ+CzJtop0++AFFmncgymvDofaDSV2jUff2JkhwbYbsFss0vov
dDMLGZSr+IwV6Aq/4xzZ4S6bi3kquBRhy2G26mxCgv2rEGccysEKHEQArH13Es0s
`protect END_PROTECTED
