`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35b3y0bKK+IMDnHwBfi/Z+P0CGPGK5JrxE0hrPofjb6+rf9EqGQoSyEKon33A8s5
0jh3DcPznv1L81++DXkCmqCSFjWTaemo8FFU/FArhjKq0dTx2LJfgGn/WPItN+++
uHZ94urmwU1xIW8l1WscWJVM56U1OIlGnlrheSIU7b8Z62nCibYVf/4b+nVthpb7
Y47EaytGplQ+JnJmnhrm1mkEG/Z3/kQTLYPT1gyunX06RY2/SCHUOKo7irzLl8wd
zQpsyLu422lz345DTTFvR5RYaMpu4O7si6G4L3idSEuKeJ57gI5l3isSJGILmHhe
Gf+W44alQk8n+U8kNE3wejDIYvFYcIXoPdeGwleyBWNn+ZurCmlO/z6hg7llvrke
YmeES2ki4GXOU7oRkUy/CyJfgzzpXk10zVIrvRta0b5QGT/O3Pl5+Y56rqNAyUDr
w8RnvTjS5aYxb6WprE0FDyLTcvJsoaQdePohrzrrqS/18U8P6tCLDMFg+Ba+jSyy
H/tKRmXW6CAPhgLmX1aYhDdecOkpBO66vmzNLXxXDfkfQ3jrdq9Ja5sfqVmD6e4r
Nkm5xJVQaK6dRxiqL1IuIx3YUQQ0T66xMCfzRp9v+9hVy2n/iGG+f1mq+z9SlsWs
7E8f5HRNJrbN65Ur9W+L0/JlU5efJSDAGsX7lleyYVPNhniSSLIl/bejKreuqDJg
ULJjLxdXe4ATdBGP/9CwKXJGeM+6Wv/w3dpXsnD5JsOLiCcf3CEDfkuFhWdeC4Bm
M/m2JY6P9yMW8NRpKiwMMf5U8w4qwB1t5GwIKg4W/BH/st+5rEfPBPkk4dB282w/
o34OvzhTiFKrXzEOuVVYDemJepa9sOJUlE/YwuLr5rmRSuuzrBylXN2NAiLspfA7
rf1liFUsIxZfaMZE+Z9SAhAopOmmLf+4of/6BLRDJk1EgSr29G5bwgRc6cwrKcU9
Eke3pdlBe1h/0r2Gc2YmLopU4ENbDNnhvq6SSyCKCxLX3Ny/tCvpsWfMefUOFtsM
Hg8+NimXpKo+jyvF5XZabqH/j+9C9g84+YonBLcX+nF0md7UUsVj1QMZR9HT2GxH
nTRMLzt507UZVOeUVIpa3QI/cGzjIepVNGm7u+ZVNd3nPdWgEiUhE9rUoGN1R+0y
nbhEvC4Fb/FSd/tEJo5E44bvyLeJVuk3ha/HB43e6UkQU5i7misa/a6DoW4R1ypd
nmojadfoZO4Ue7qTsAsX9YrCOd9hObcxmmXYtIDw+UZncs2N2ypmRGA1Blkq4z2e
`protect END_PROTECTED
