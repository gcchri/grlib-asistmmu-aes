`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fMMZZmvCBBJlf3hJuWP1qQoHG8lAgjmeCZRS4YG146i31P69L4Ur8tDixYIclaHK
wcm2FJ+t+1KwdvaGJjL9J0doe/h29tBuiirhWDjFwLIWtZOKqTsoZI+NVP1Xn63C
hZyym9UAF+UQbtu/sNbuDPpnU2rMsn2cnnfQbSQcBzJScQgVOD+Rfh0oJjzJf+hX
M6hv4CFcx21xJmtL3xpNTsy4Q7ABPtVCEH9SUJkLFNL22UXijIIpLXnQsLzNljO3
C9kvrNjCikYFen8sjG2kTxY9qV8raDwNuVtbHrCYv21Ox5jSu6BPsbFo2FHnwCMv
cfVDMogWq0975AhFdT/udSpGj24ZOcYrUexzL8Ixwqbi06ep8SydhMHkyPomsOwJ
qNt+C1MVPzG3LQdvP1imqXOLAbknKjGhKZFamfFJPfCfrVkVrBFN/fw9Ck8+24oA
F5Hc5jtxFl49Lp7AG3N+Rh2ZtZvNApRO0hIZ0CU+PLcnxnWfptvL44u+oB8f8ILa
FDer4SEXgGmqhj5WFggVXfe0qZP6tjmCcNuFako19Su8WvIYfF4HRCr4fP3VhvTP
/X5i1fEslsaHAijTnYyObQw1Ky+lacNGMThrjWLI/8xnT83ZUeKfpmEB7KUO4x3/
IOGdTpLFkfrPQDQAqZul+xjhrbBCGfp3jZoQOBgqXcb0SLxpOtkPNWgdNdQExT+l
3COI77RXlILG905vMljhikf9dFguCx6rfIaXHRcRdHgf/uwhhOHA9Z4K8u//whq6
N8628TnkpMFaXVrYANrQ0Rv5RG879kLdQoyDVOyzS6TXUN+4Pk6qlVczjRXQ1ZMS
lcLPPmHmWeJqLoXY1n7StBaDvIH9wM05eAj778tv1ISYIleScs4aWQsqVJCwOI93
Hx/vLCdnenWy8t06pyCCs39kKjbwAAi3cnzVzMMZXJqdN/5rvnzvgFCj69A9tnQ/
j9mDGlaF05CSseVmzLbbs8wmt3kEVkcpq4YVzBIZnROyvfGp+G0zPXYfhj1CCD//
hlgoDl06cQFYKs43M9wI/y9HOPbSt86fitgsRTjvCugKp2A/d8Yp401c7Vj3AzA3
p6JdNkcnQlZcAfibpqXmdeAsu3QO2uVz+K5J1uFj7B/PXCJnhTxiYxjZda8DjUPt
r1V1+BPRUAaZ2eYOXYsHsQWBSZLwr8uW4xvC7xE77OguLl8yJGrF3VMFqO8R7Zhk
/VPPmsCJ81VT7VO+q9QdOkQEebwraiuKJZ9049W1g/IAOM2W2amQgzN/qX+j4JWo
`protect END_PROTECTED
