`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQ3AxubKC6sVzregRlbwtd6IaiOG3AUKWYhmucQg4z8j/Chi3CGHu+GpFBh1I+Tw
ENTURq64K+M/mbOaXkBfYeShJu/tBFA5AL7kTwMOpEwDwyJ3FBJKroYjIdbTsITu
sfDk/mxB8H0QvYkMBSmqGpGNEq4yjt2Uc19F3IVF7d0AlvlJ8lZqFKTc88lanwi8
DZwRkF0NCWduh2zwZJNZJFdSl2tZi3mAuU1uDyEOqvcbeBiulfNbuvJLNKqM6m9T
VKf1LqCe3DPlwBOVpQvKAqA/xHmyfHeZ+nojQwLMp/Vx022368OHw5GbUwkpPghT
rO0q8JRppLcTwZGGf06oQUk4XBSrtBek+bjvch14lcOrjWEqrtB7RxE+nfv4YXnb
Jc0zSZ8yir/riZiEetoUoDXPvazeqG39xRHpnFlB1Dtm5XiCBSC8FiFiSuOeh02O
BSQtbgBNetLZ/at0Ce6yEiv9sV1RK7u06GMYxh8m8SRywepFUiDVuCbE+Vk2vCjs
`protect END_PROTECTED
