`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CHJYFkqiDrm+9g56gEGK+euOOzy4KzQRVJSpMOoFobkHiGIDRNqxvZenZufUK5Ga
fu4IjZ1Fs067s4wdk7EXkIKdm45LlQxob8EdbdNf9ZfClvo0gCg6yL+cE/4C41Sk
7lS4c53Xqa1BLRq+jPqo+1r86lqBixWhzIkHQPWPUkejqWbl09qY7wo0x4s0DLlO
H94rP8ggc5lIXO9SvOKMBygyXyq939NQrCqLKIkeGbOWEN9DQC8l9XPepA3KB08E
QwYzVR1S8ozVZidWXK2Vtfr73UCqP38oeu0E7+xstXeabHW1XxvwU/rsO65i6/GL
k2vPnL0FKCIUzAtOJJy73PrDico4F2eJitjr/+ASa7grvvXDMiKiPP7tnZ6XwS2f
0acB9I6nSVsaYrilk9w++cAf35OZW+1o7T8N+LlLppAs6v2faTBI3mtebZHw3dmP
t1GgTYnngJOdlfoHe2s0Ubma1kOF3UCtJaptD5RH5rYifSX9t2olymxvKrUqLFqK
GH7A0Hr8kl4SuvQGdshHy2TLEjQh/Y/TRnqWx6R7/aYmJqX/dhW7Jyb7hWH61HyA
3F/nrhM35z1AuwYau/wvhV6paoPcFsva4wBZYIey3QpH9FBXFgCBu1DoJ0/s/zAF
S9klJhNPCqS4epzGwquxVQynl3WI3JyOBZrxNkqcf4vGMGCngcc+0vXspSz4Jnzv
FHfx+PqOjPH+4rufyXh90n9X/FeeyBNOJzud0FasHsuX+I1ClIxgezz+SceOnbxj
RWFRFcsb9gywMUZPlMlgVTdJGvvVCJ4Nm3A0Ai19+d8/TTY1d/9k9GZ9JM72JjgE
5TiRsXz8Ew2TJxU4Bmk+dKPy0Wfxa0/cp0AIVgAu9Phs9+Qx4hyTBm3m7FQwVNVu
ri25Ky+avu6osEfMSKFsj4fn5Ojfww0QDT1gqtkG5xpmvlCJCbvziHP5qVA2xmj6
GZYzkMZezsyk1TcuN6rTGhYInoeWROWb0HCNgyNV5Gyiq4jX88NEMH4ZJO4Eq0NR
LkbxHGzAC6RBjNzu8VsE8kEC8M4MuKAbO9FN+9sms4MMeaDXoq02kP09VlZsCuqm
HDs2nNRGLrPQUmgcrUC8G8RXRxtep6iIy4pYU/nj5uUX+y3Sl8oFaHJAUiM84E6j
llBnpAZ8VDiODBr1sFV//wxytsJoLyHkr1Wuu55ORfjpzUcwK5a4MrWgC51IvuQy
GPCQd9FEDgp9aL+07A57rW7BCyZtEoRBhQEdl/nVgkHPp0kP/0HdqgY/AsUe9L2R
gTw+P1FQbcr3bpWC6ECymXatReKHxec6Zw8qIKt7wVfBjRThaxDunNyUiFJqXWFe
ZiWU7Z7QLaKoOtp6RMS+kjU+t9ibo5eCsY6cxD79r08nUa7OPQasR9/Gv4KZp+ey
CCcXcYqsSslDivMj9pL44s9rGP75/J+Hr0KMAmZzbxFB+6R6GyKLumpCpddu8J5N
N2HbXdkJCKjf70ahDd2A++sBBMBm4yia9l58Awjljf/Hec15mIh2/ylaMLX1zd6I
V9VN3OcvmRqMCmSQsWwX4gZy9rao90YslRJOuBYH6veXJt8NmKjkID7896/adwAI
nKd+WVF9wupEvvYfk8HasJ2Jkx8U10/zNonvMPkhqFndLPG+MKhXCdO8dyiQYAm7
a4qijtw1g31bEIe6YKKOzpbCf7Fre2S/9cHELkNuzbEHRrrL8DK38n60x6MPA8/S
oQ7cgnSA2ZmGM6qx4lPX7n84rGdODwpkdthF4Ywc8fH8YtbGB3L/+NZSRHkqZs17
kwoBAZaF2reMBlmLnKRUUWh9o46TCe1mydQvd4YZ6/qSfWi6kYqsTTyW6RLvyhsR
t0SHMWKMLck2RHMmKGiktw9fZnXngrjFkdQXzSbUq3sFd4yarSPLKueBwuYnHyvf
uMS8E+cTNXN+9jN1sVVvAaqiPg3zlnACASxFxpPUI/AM5aoq4mtZmeL+lc6vBI3s
MqcPJZH05KywXJKUt77crG6uRSqx0lsj6/bZ1hVUoVkuAGV7XKmYwnU3mYTQ5kZ7
amXk/Oo+ouO3cCb7meUsYe8hrskmZNXN6uM9JOyYO4VOWahnmoRSFP2NQb1oIeeT
8vnI0cxlRktYkVcWmHNeIsKyYSq0tIGO2Xu8EkMWm63jsyHcS94iDyKcTravajaA
WY8RyyksJqYXmUDREOY6R7AwIkj+IYw4Q25tkZNp0ZtZI9D9W8ERA/toc7ZcKTG8
1ojWp+FTDrvnY0j2oAQBm+zOYV2Umbg/hxcFUt44z6TZ68UkUCtLTOzyVL4QqRPA
SbRstmZOcvZEHOWPW+yG24KbldF0qsRzmOxAuzJKkVlyqUPG6le68bcsQdAxmRhm
TKzn2cbtSLBIo+Z/QartSC6Hyu7DL6496zpfYItO4zc/zKcmv78WkmvmBZezQrPO
gP8OhqelV7y3TRhFqemEziGIPh3d1BlaRgAWekFm6OCTJM8jNNneQXIBbaYP87iE
iye2xjH6X4bfqxqAaOtKnTBGkKZ12nRs2A8XB3qMknPVGPPvZx7SqS54xjBHcq68
ywfP99iTVqVw4jxrivo8qMj0zaIPRI9Pt/WMO0rbnpD9Ul/U2HgsasTXG72qNh4t
xzDihZlgIqMpG6qhSWGAMV/VYPKc8k3CC+BN3vFVz2RX/QfuyOcFWk3Y7BJW7k2l
SasWn1zF7iSFqf9uVG9cMOLYKLdPVC3Gx8XNvq6FLkr2FeoWcyf76ExIHgd7bbZ2
2HmaQxwd3BEElwshRY2wyTEipZT4vr5Ncs5xBHM1XwIhX/Vu2movbMxfZo5ZGh/p
WikyX3cvGKLy5FfQUjIO6wdUx65u19+wnu2GBLKj4CGRnK9s7REHH60zA3IzsoPc
KHfGAS03UXBMr0BhPO8bCkR05JlNP+tGG0FJSieSjtLp5GnXVasQTCONS7uuKEXL
MGUNLYDb7ChuY33TcgN+QEKs/TWyEeVRauT0j5wuyhI=
`protect END_PROTECTED
