`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0YA7r0QvkeI85kzNSoUk9VpIVb+yduO3UuzTNCatIarKKHeNOd+evRzXe06UUeEN
XlNay1WjOn+omiltAOXVSUKFk8T62KdLjoWFU3AWYz40o4hifQmpk1yt+R0B8/lU
QqHaz/iyROPtQbT2D7zulNxZSaMghEHqseiijC+J6xmMw1NaEVNjKK8HAbivepWF
F9l+0/+JhF2Og862044Bm+Pv8b0uK6V6wiTI5MUn8YO3xKOANW12GNUwQ+0LYCdz
Z/5hLWOIgcLb2BDnMIEptyjupcVy4cIHpsTkeOq5szA/tn4xT5dcbGvTLnq58Tey
AwpvCgQ0XH8z+C3XOux/si94U5kHgaaTTQ+t467BR82hvuaoj4QEp7SkCtl4FgB1
+4K2vtx9OC9Cp5QWLSZfilmFyemAHlqwdRdp7s0c3u5I5WTpvAwU08uqlmha6CQA
`protect END_PROTECTED
