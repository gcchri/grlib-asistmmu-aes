`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p9djE28FUNjnac7JL3iPrIEBDc1AEvFwNZt8guBPQ4QfHwrbLEiLTfZgYtonkLpJ
93Rb0kWV630pskBJMCSKW3tSvJu065iLAtl/2MSZ2ZIkgCP5DPjcS6KYNv/8bx8W
KvAgIta6xRPlZGUZjl3YhWtUKNVvbTZWvdSBapc2/l457yipIurNlRLRPa9EmQJK
YkqBMRY/2x356XaoFgYdGWmwEpq287W9YYzqbhZUUdp3tlxnf1Dnd5CXe7oifoDy
4fAb5Gy1n5OuuVrtZ/EzFMzGAJm1dLm4l3Io+WbqHedn0qPtFEnnUjRcGTf8KC8P
laCOJxOGBCsxSfE/KK5RNdtniNX8mt6+CMJqMhh8zbUeYScdQmspCAyLB0LbWnxc
nGWO5opU4xP7eBNSCq3sFIpqsUN9tYPcC2Ga6+kEU3MDmxLeONPzyjO+ie00V4TD
uq9hvuMbMvPpQUojO/Zu36dDsrQghNv3Sr31r3Rmnpkhxir2BAP3cLHDY0twiyKX
0KyyGwwgbdLPwvk5QlRNMMupyFIva2AwunVsyQdv3qz777hhJt7EB/sXvO1DMB9W
wrNtX1D+wj9XLLx/tEyamr8cfWi6CGXPgjx+oNs8d+5+fZSA8jyywJxnPQQKNpCG
SLFjNb4R9P/kEDwxq9sRTfqia+KuUDTQIOwpZFPZABgQ3cd5Y0RX2JI3RY2xuOCU
OfspT2n+SJooERzguGmgKodU9d142aSUEOmwr7eoB+Htx90434r4yQjE8pNt1dPX
saVpafyQyCRhTUvV5dI8btzt8d7iWELHu6+pdKERzOXjFhCETDtXc8nGV5pYLlSz
+hRN3Kr1IObMZzO2XLUGVdsUfIxAjONrAJfgzjj6x9vvs3fHjejz9Yqd+NUTp2H3
tk5NWII/pts6YnMY82nVmA6u+mNrVkCzQclJk4xrB7hoK+scmqqF4YgtAqhOTFzr
kjLYLfsVwFIbms2XwtP5dHSyDu/x1nO1BGycn3ZCWmsOd+RzvWQnjdqAsVbKqQaQ
GUpqcPuZ2xoSQmTws8dAB9r9kQ38yyD6wqaymTpFVKE2rth6brrLorYgx16YRb4d
7P3WZ7X+cLfSQTMgyeXYLcxqwt47DhcUsoRb+tueG6RweCvHORSOVew5MxWwb26b
xufihSlVRg6GP8KWHr19BfxOimezPgmRs79GP4bpDVYSW5+ZXic7n4a5DoaLh3Wz
Dctsr7tqIcM5YCjCnoKTl0O+KMsmx/dhockP5oHM2sBMhwNo6W29n2KVZij9C/Zr
KuHXPV6rWzjQARXJV8icsXj8ag3WpG+Zks7gH5Jea53oIP22basMEjGxfOOD6XIN
vqU6TaV4TAQw0aEgEVMNUSKXMBanzCvZkYBsiThdgyDyj1U0CIbd40B9eTyJd8Ce
0VH13zEVnux1tsy+6j+tDeP4ol7eLd2TxUiuhW1DtDIa2pgyXBvMtlY6ZtkUHdju
bPOr8IvudOcmE041HlgJp9LDO++JITJbRsx4HLLZjZrbH5LV7NNRztUPDOWRp0Gj
BMat5wUHzM8/VvVy6cYePRRs/9WyFmbNpPSWfp9PMG36C6VYglCrZkBg/jqgPH0O
Urhyx6SdGOZLLmAJGrvfqplEtNiIl2UjDHuV+gdm/bc0e2h1Eh6RH27ItEl8eSVR
Qhm+ulILwI43Z5ykR0dlhjnRjI0QKHT0rDUfUNufWc5gaUFX3fdfQeCdAA6/JLj1
IAVAz7OntNbMKf8PcB8ywJZ7aiuMnY0vI9i3iMRBJN9biA2/p8txGm9t3SKy3yQU
h2y57JI9viyvIdMy0D/LZvhg8hn0EwYtizi7DDp1cbDOillLHTcAMj1OR5kc9yoR
FokvsuK9+HUtGfbycF6v8TkdsOlqwWX/bE3WZV3hnQ0=
`protect END_PROTECTED
