`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fBk2S7TNxGyOcPSadSxNOzpO/O4MrmfvZxRi3sfxDV7PFIosaTOmkSSmASVVBtDr
zP4Z2Hi2r0oa1e+ukMjluNOyEqxqnqkm4/jC109qcE/ijycs0rzAjAAot27TTF7M
yTFwrLpRsR1Lk70Nh3ppdM9CAYKGn/SiHg6Xe5Vx11KIwhLYzt17FfR9t1pj4XGe
cgAQX4txw24gwxkNKJnfigVjPTkKPd2rpk09DVHIYmWDwdlH/6nVxMCkRyGYaCjq
EtnAEeXTlQKVOiTL3vF7Ejet1oE466jIWpNQNv4bBil3sMHAz0dc9Mg2v1mQlwL3
PKzeko/UrD6nA2E4OM2ZxJjx+L6wRtgsbpVuvk+rfvscF5wbon4tP1vKCnlvfI1z
h9KBZOrNy7y3Q52EiiQh/TUf9tYhtHnKi+c7kCUQ8N3Wtiiy4NCZ75gzAR97lXE8
Hlhnxr4SnK0atKBSLEMydfBmV42zxL0PTMyAeo/IV9JsCgA+3YZ2EUFzl/MgNc1o
1XtJexls9vGt6rG4dzz9SRhQtnj/+IfYIiKvFG+CUdyjHk+gzIjtdoIOFo8IxdYR
+GIW4lHTQEBpVvW48qanikJbcwQgu5EhkoITM0RTD6yShLrOF3QmPGi28jC/3fZ5
AJQ65w2lyrjNIrkiOHXtZQ==
`protect END_PROTECTED
