`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAOuYyQXbd1Xv0jznCTfxl09J+oWprHIe190PkAId3BC2Wit21DHRO21xhlf7boM
DtE/VwCzyB057C75ejg6pczKRiZtkZC1rtTSQRNOmOQkdsFs8P25Joceatz0PiwX
COqCWHcgTTd2l9PM97y3wFTiR8MylzMBKoe0vgmHqT1JmmMEDlaZHedTW45eP3y/
a/2nLOMm3HSwEKbSXPAe9pphLifDYfRuyhmNnIf3qQz635e/Eq5iZiQi1XKy1juT
pF/ZUWE00FBefWFCxAbyZFDcWZ7bhvdibF45JMHiDQ+wN34+uMJEmAupOR+WxWdJ
NrtRNeQ5t4AwE9V2e19DlTAWFBk6CC3zNTkKvPSUnv0Y7dVwp496YUURCOF2hR3o
HGZm7p5nAJFKHpStxCOWuozCAxTobigZJvMYKU39NCwq47uicEBu/jP2Lwfpw7n+
TA6alyyr5XL+0jl2BQioIvFnoD8+Rdh08vUvFf5uGgWB5ijAW2mBwo1nZ4gi2uUS
mhX+uhE7F3nZOyucHaJD1fCnHHYMfqf5+3HC1RjgWhfrVcNlCjLCTPnKja7AzDOU
SD2LA/Pb/ssBoLmQeoc6Q49psEqm8rD1xPlPd+4CNI2vBPp0o20q6gqflDu1sK4V
7UYCGyom38vgq4Qk9irVr0P5Z8NlFF52H4gwonEFtr1oA86+7BV2xxzHfgLGxUvV
dOanTJ/pcYfOQ/t+wXqX5fmzvGlfFMUHsBmLFFiPTb1+ZfaGu4p7jfqfbT/Tl+Px
JfDRM5Pf0BhOjrC0rEI1I5NhececmTVyWQ7nuTJ8QrNP1ujMI7VKuwpNOTA0sPXQ
W4y8aFZZhFDPyrHo5/Iz6bFf7yvchBMuWERtHPjbeE31hIhAxBUz1kC8i9y44PIb
NRXbo3JPuPWWnBu0HJXr+4tms6iJWJmb4EKSwxBt6IatZKNdSnikMlhrNnDBva2/
wMZQitl6bGDZEB9e458BYkzy6SBI0eZrMHeAS9oBpSNgR+XY3duF5hR2HzS4hS42
IUWBS7uXN37uVs9+/IrUCxJLzb0J1+uwvepHDIx6p9BxtSSOkGXuxQXPPs9Rzbq1
W+HyyTPb1NfJoUEct74PJ/7M8dK6kBvxZ8iDYYL/CDSH8EuKJkNJiPwsUdUlv2+v
nNjR2sPOjXboiBPbIhdIwItD+yxhGND6XBGx0XUEEn6M0FziCACaaCPGWmpnR/gU
+sKDB1rlt0CCY2XzfBmCBjGuCZpMRR00VsRiygcCl16YsOs8IvcByGGRaXJEn0rb
cRnae5u6yQQsEtPZYmOla1Yaw//IN2iHVm47NkP0N2dDzm5O4WyYDwgL71Zqf9Sl
ctKPQPTZSDeF/7Mlmv3d7nkJ8nTB5qWLvypubUezlu6w0U3khuLPwZsH1GkbZ9Kg
n6gAUWHu9oqFUP1L4n+ZMKQrWKGY5CrimfrUKAnPRx4tuv4oPyaLg1Od1mcFj5Rm
sQ1I9kMpQwsf3tF5pqrXJLdix/YA3b+SujKoeR4SU6Qlv3Q0dVjWCSp1T1f5dHDg
E+kPYVQrHUJ87fRotak1PWGAm9xqh48oXQX7t7MsMG0kQfYr1QicfES7Hk1GSZvj
Ui9jEGdSBXOgSwFqXePrlRG5fKrmGdYkL8ABNbEBHKvAKJf3IHmZKBNIovyoBblX
IxYC556oZ9mrzLT+np0znMiAOscEDtHc/URGI2qhxPUDsYn0SG1y7vmQAyOVUoZJ
q4PIfT4zZ8vThmeZ51HuW1uDo/ZF25RL9o93Prh5g7wiPeHst1QqHFE/qW/OewkT
1eQqim/JbzpPsu+yXU7UqIkDEkOK5ML8fLSttbDgMuOvN+FqVcQYdwOI7x/ukeKf
7+d/mISCsXTRdb9+McAKBu3jpk8TWnmRM/TB9RE93RAm/Arf+g8azVX9rkxGuLdV
HMLmX8f8AM5062pMU2+5HMIWXykIeU48lRHrA2u98mZ19gtFJxMZRX5UESbxSJU4
rMyhbq6tzqmMsm68/AUB4ZF7EyQwvNADtIuGGJnRTxRYz3j8dHQdHrnZrOpGzoov
o6l9cf0t/T7xXf/l0V7bBRs/jMsE94tZ6kY0lXzx7e4tGplwTAdor07Yi5r0vMEz
i5MQckz2l7kIIjFZnsF+0oNphqUYDigKTdAewRMMTfey8vHdJMUZG2kXoqHs77m2
SZNGp+0z/fyIGOCegVSaEnFoa+s2jZArrwfrEG6C1ChxKRXDAPRdAfue7OgIb6bq
DYvBHyXL6kZa6AC7mvc8vnkL7sEgDvWSSea8kxKHIPbM4s7g6nFwqIvY/cpbsfVy
Hu1AQ55qWhwVjihjm72PAFs7ZkUrk5H0DXgC0+ZtBBW/nJg34imx6YUKSt8SSos1
GK7Y7chxkUO5C45W/fxtFOdJkIcaSEV/PJRSBD/FW+j4voO2Ora5jf565RcZmnAD
k6doBdIyJaUdUVgbStU4IRfaQEG7EnSnppbneERQosFS4Yp9KOmsKMNE7sliWLUq
YSQ94jj7CU9/nWszWh3GkNNWgGuWSDsev46xDNA1Zo36GplKHNpCckpUkCS/2rzY
`protect END_PROTECTED
