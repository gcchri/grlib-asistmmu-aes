`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F7Oyg5sq9QCc4d6X0iGcCbm4RPPhcmMFQgkYqQ+3pWTsEt8nMQnZKz7jOYjT7YCd
HZWxx4yotHXNAI+UBccYs7TJAMzcaz19ypc9QtO3cQCt8aztsfbDgiDbkor99vsh
k8VtO5nLuo+2BI7y1j1S6L59TeE3u4N4g1dpuZiV5anIvT5nrQDu194NuUAUNn0s
Brs1Z0NNIbGt0T9nd2SsWhE5kwPB0CwKvFq1NgRp0HzkyiPNwvX/kjL8tVkODnJK
wQgq6w9BBBzhAbTSU5YT9eXMLfwwqOEAOMCVdC4jCAePQldThZKR+b0HEa+ym+tO
uKZstz23z8RRqnOQN40V8hKeCYBe7J6Ms9o/VcI75X2YAbOqfvgBHji1zKEoil+Y
rN9KBguNoBTX6eGO4gKYQHbWgC4dbU3TOI4CukZSEXbG+978T/FW5NmISi46LYJ3
YA9QfXizyrcxe8TL8vQMrEASlKs+IlmyEi2XDq2FX6EpcPq8r//2fFlNT2DhUld4
9I6og9OvrzIM1iyV1dmaxp0aplb/yIDWG0KgVnMpdBv9DBg5WVHx9ptEq3xHAJSb
WhsMR5oR6beUKCuWo+cYBFvUOnqHJ8NFl3cAXikTQ8hflNXczV/0bz4M2dcScuun
EQol9gmzaNyjElAXbxwpdajOEhf36IWWls2+jLrD3az0H4zHSmoZFKY6BgjnSGS2
NHYm8mpc3dEYUVTJY5P7BBSDj/5vcUAm2vnWq9BY8yBuhAvK+9Iqy/pceUx9DS6m
qykm4dBDSGm/obpp40jmpmfjaEPDWiZLnf+u4fKDdwqAFQmnGM7Qv5QuL+0sDwNO
zK2GqD95mwTT/qDxldS2BQ==
`protect END_PROTECTED
