`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WfaNpR9zIxB0xFzMh84fvjPzrOey0d9zdhFWGdfEjw81Ayz4YFGmiDjnf/MNFM/0
JcMCTCAtt1SqLWdaPDVlahCfmeAQOD72Nv63mQIeqrAtoVTZ/rtUPbbDaTnkqneb
ZsonPyy9t4vt6OvanTlRE4T4zHkiNYkSfgGoeZtsTBeko68z6Uy5Yb2+mun3/yuY
jM3PHbtEnTBGZwC7zks/3alDDSGnYhmBq837MdoYi/fp9XRIOso4E4yh4GGbAwQu
LFHY8ZzqMKKatVPG+gyzzq8vEuRkNeXaGHjAvedojX1BX45btWy000H8lasGl3tO
5hsdL5u14KPJUlTa2XaWBTwwa02KMJ97rMsbdyjzMwA=
`protect END_PROTECTED
