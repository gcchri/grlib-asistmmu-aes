`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5670bq20swI5p/eKuhyCPGVW8IpllcJ4xzacodxpzUv7C5X99MflATDvyEARJuC2
0MzLw3w/9lqEMSE0XmlaUCR0YjPJ8vW58LeORTpgB9dOF+Ld8d80JjIAoUJitF6B
eiH4UmR4LyoTxml/euSrCwtXrnfKWx1LUiifHgAiEXj/PWL9cfROr/kMeshEeBcX
+vcqkKmAEiSrz9fkaXK8lZVd+vBcuI0kJnEO4y3sh8l4Jei8aWXFmauEvKqVqgDn
4rhmO76iQPz7YV9CIkXQrFy2SVekQQze6T7EiCrabnyIRIPyWij11DiFy6SbVEYq
WciGhGYHFL6MU0hKaBMC223gBbjA1dA3SLj4drqT7APzRLRiKvnO2p9AnBj5ogEw
yT4j+Epk7KVfpuF6S8dUP/da1maIT0w3TlNpkArom5qb07MzVxTS7j/4KYv1eF9e
/rT0H/Pjc1gVCsvpfsZsiJa2716jTH4Ugh9xFLoYlINc3ja97tY33C8WN1rzT5Z+
1rLK9vFG3ZBWDGH8xr/HxiddcGaJ4aiQvbn9cS2kNe4wS4pFodKb+SwxlFZ+SkVl
v59/s2Ml1Y1OnrsfE4wxgM48m3lg2Q5O8Dp51YQ1zbXjZU7bA5UWf7ryw0DFYkmL
KH8g7gNSGj2AJ8Zt1hGAkJ8SoyIu6N9JoC7V5dA0l0tEAFyo0JNwGndWjqSSKdTP
8T64W9CN0BSIq37mgMKJJlx097Mm6QXe5wmycE+5XY6rBpF6Jx+nOxQas/bgky01
zfSRIumTYlPCLDAm/qHCNiMs1rrLRb7XxHKpqVrlwpQoIqdrJV3AF75/PZHY9CWe
7CArOe9xMCcbqBho7j77SI/1qu4I+NytTbO4sC8QChto/ZIhF5ZyIv0SqW6zvYYh
YIYhMryhJGxxC0xb7pfbAEgQrXXz5RCxuTTMPauHcHzQrgiKrUKhuB6MiF5lR7m2
WDsn6iQj+PESkvUEKK/L55nkEgeZPUmcj9C4nZ80m4YgWxiJuVLa3MoM6PKgRVlK
41v6wahMyAfsCd44wCu+kGmeU0FnbZ9Z/8eO15KlRBtwTYVnPJLE+Z2IiEwPwcEK
XBQDhnWujNifsWW9GvluH0QuHfZsGb7xgEjdeKlRv5YnnMGdwlBAResdhQVeVupy
oLdKGA0/WT8ItraLWVBRGvv5y7hBe9sBHSg8k21wghDBy5DKaB0aewv7We5q7dPX
6dAKEggForFy3+Tny9h4PEGUYrUXX1S4y/yqZBZz5fJuKK5lo2dIWb1yuhHx1z3a
e0rrAhc3z7bKjSZUmnCkE2lAugvTtdKCkAPCJC/nLZa7LTRkKDEeKdTF6Ir4rPTx
ZHZKr4XeXwAgmJkYFwuco2627AijQ0BdC17Sl7HkELl5oZ/gvQITmO/E80Q2bmro
poU1GzO9H9HGQQWlp2bKR0d2A5Oddtzc25zkuV1kN18Ibg5r8uZUN020cxfbuTES
LemAKHo6mJwvo2Kwqkckb0VMQobrgSkkWWBXFzXQd2ABAcVJisbUDw6K4+vt8WLY
toI4fF0fc0ucKFVMPR2cWUcL71KyNVDQwE938BUKdxvei47aBqK52ylBhjPZP+fg
wLzOfWtj8b4RKs/YweQ6i+4fnKFCQJt5TUwNU27MwjQIsdAskR6ArCqAylgDzCvq
hCDLmz9DtAorOfTGPHbGWWQUTizhOegYG8/95Jers9aEx66vjUYpe968qtZ4d103
scQwDAtrhFReJ5Xzl7RBEugqUw+OLp+x38dJcVC0nVDL02Pl4R0QKlmYHpKw4RAV
GwXjXqpzTdNsQbD0LeAItIbaxyp7PU/gKej1H/TL38q4kpiQIlm3aIp7d8JaYYqG
T6m9nwoXrvXO3NXTe30CAW8Qf08UXyHkyvVRLwNvNoDe5bNt5X16DeuK0fLZNMOy
ouiAit5by85ZAm8NoVtgaLD4iW/GAw6ZRSSe67kisPe31XBzPsamNBo+pZNx6w0b
kuFbuyfkr4hYw6TSnYyXypirpxtTZNBo5UxWTA+iLENErpDvBZ6InbGm53RmAesM
87V3jRgoO07BS2i4UzVAHwfamLT/Wo/CF3u61oNtgx2JzRVBWIVz0Vpm0g9Narvp
LBCVgbWzxvYW8I4A6Sl4r+FqOLWsncmlVQwNz6iQJoXygBHcd6vgxed34vlM1D4t
1TXt5e7j6AoEJnVuAqcaFkeeXbelR4vjNnc1PcBf3sCiQbOl9en2C2Gei/n1MXes
c6IpgLLcVXurR3P8qxM9wyQ5yk5/5irFUCuMnri/qGZDuM7HXeiHOZ9haYVXm+23
rl+95KRdwRuIJkRqDLx+rn6OaB1FXQzQncHemOitWQuz/G1rRWxbFQRGSJMiA8CJ
Qa2SY5uX7U0syFfy4yIwnfts79rGfG+VmsD/zgRXplY3LPyrkhhZg7jjAJX0Zdk7
NQh8/Mary7/X2V/V9+PcHOqiCK2QhZYlBI+/pQS12yDkMltP58DqKI7vXe8u3dIf
Zx044vNjNLSTLBKaeydMszLG0RQB95R+BRxtZSOd2gjUMQUPqMolNzyYLrlium42
2eBdfPPZNgg2+ayhWX40+wjbi7MLS2pTlzanpYWpHLHr93qmIyQorpQtoux0v7J4
WjSwwZSBmFhK2yULawpqXbntvc5J/WWbu2w60Hav9jlgo4NUCcSlhqagOR/eIU9U
gGGTjPDqkuR7auNhPU0XiAFubeFggh8AYCV0nk0tb80G6x/+sJ+FR7z9Cur4XZlW
w0fcCI7aoHdeJ1RLhflwmdY3Aq+yDX0a9f/r23my83mnvZsk6/5h1w4o2XGVFjVN
3midRdYabOyp3sgvjGjtzQfJBSR3lWqIFCjrj77JqIQS9zEO4UiFg7/uNtkdjEVO
SS1cQ4F4W5E596R5FbBmIU803yt1G5PVyrepEnK4Fubx7vuuBEqTGYLs7PJAGyod
fWOeHJVpum/Q7LU9FxSSie7dgfQxWIG1vFpZGmCfwciJXsGMR728v1QwkjpSUusz
vHwybN9lh5a5GBM1pRhOpRqjbhVKpSvtAEwDYG+WAzfG6usBb7R61puxbyEeqvPz
kNKw79JQOhKZkMdtbNm5VucywEKLGojASPq/r20GMWpJURUoe7Ij8SQ1q33jnHI+
csK4xDg+U8ECoo5wKV0/lx/gsa4IMI+6Tr9GMYQpzV/2TT/J0+STSdLjN+Vrdoes
xmPakp99YBq7ZWX/p/wCMO36lMc4EOk2Cf3uc/IpoIZdIuZR+unaeMZRDeo5QJH1
rew+r4/O6CoxlOZtdHy02rzrXDknL1rFTke+0iFfJMmVZ1rQtY+4IbW3Uyhm/4LS
iMjT5Nbbs0fTpr36uHq9m/CtujWokWFUXdAFedaQaxbBW2pDeCldPYYewiqJCm3R
pcJC/ihLuwhHqWvrxGRsMEYUk5X0Too5AfHk5Vw5gt+1L3q/XVvmVCHEj/vDhKqo
FGdgU+4vy7kSRqwLAOm4ZLLFYLM+U8UI4vQ5i+zb5lGEfWkR/C1XQlnT2oh+Olcw
fgPG1deOaeDbtixhlT2QQU3MZZFMMmtG9NDNj23YXWwR79BOovGoFefaMZOKA2/I
y1uLJ2hOygLy/Rv4gZyhtypYdfa3H3TSwVGPCOa88+bnCf8896VDLsBBoTTTKTj6
ma7dsdB4KToNuP35zLRO+hGTNpF+FltV+Z5JNs8pCJx7RCIyC8W1hDQycOtdR2xv
n9Yp3/khZiDiwkhxtE8K55bpIHYHJmCq1E7hq0NLSaiiJ59lOEoejUrzSPsjpNol
URxzpw/xrSqY1JIfi8UZXH8sLYLJUw0pfdpwbLIBMu7fJrZcqTOXk9Q4wJM37Pwe
GKnOXi2kg4sla+sqMXSedGsfYRSZgWiTezjYAGkhmGxELmVomNmItbuC5N3eoZ/F
mqgWN4avbZjFUEqKBZO0VIXySpIQvoR/uUo2CU+VmOrd3wVWRREgFe+zcNul/DyO
pUxilJ3UzVFP94OITJqdsr30IhdqUVv/ohT1BDOx3A61mc4QNy3KNYpGtndXzCBC
doqKMz7r3/pwKztbnpVt55CcDlR5TCg79obZgUjx1ImwLstXjGsrja3X9rZmZcwY
wUTL5eJ7mGquClb9K2qt9hrLSpi4ZihX0+N525ehD/+pDJoMPE/Bx05QNh5qIO2j
dXeZ++r3lpOyNgLNCAG8VRjhWfaVWyvTnXlnNRrCorLlSHPakSl5XTChXLLBa4yw
xEJSotKUKYoJKMdoE3HuSHaB0JDF0ayYNMzZa5H1UwA/ror2VDcUOq/us5Gs+S/r
1i+3gV9avQ/9xb6QwnKXwll8etKXk2XcsDO+Ozrp2I8zyPLplpl14owwJqORIPk6
SgUONV3Kttih0OvtBLdDfZlI1Buy9kXxbTK4U4GCPx1xsgxKvthC+2JWTmyDAK10
5//aBKaBeW5sFMEHAFd2fBwGTm/+QWpzMTK5GWYVFAfLlqWjoT5k8UhNvxdb++Wb
zqvNc7sMfCykwNlNfSeVe3hNpfmcgXpBsmZ4ktrFFijpyDJb8XwswwUX09yEubqR
ZBAWmvepJSvM+QIxeOplUhgrZu2iajFhkBzjc9CeUcOcUKUzl1KXZJ1SyohLZ0jU
NrNFMpWwz9H+ovcamXi8JRrCtVRzUUr2toqTq2+ng7WSh7LSAKwY0BeS23kynwKo
ePA06GE1ipfX/9qdPPojbzRaNGq9djZ+71qsWL4pkr2gE/PLyT2XWnmVhytyKzNi
9HYNzuq/cbP7uX/21tx8ncnGLIxNgzd2k7s9slHXW/y4+A46t0MKGjx76G4tCHgF
TqxIdCoxDJWeBMsZSNoRxu6yiMPTXdR9cgrpQ/Ttjnls+qzIQPJG9xi5E5O6ZpAa
W5bTOd6Vdgalt3Ph/wTqa8IjrM6GoaNUwrKcjsnQhFRcCsKur/Vlo6vCwz119AwT
IOWXuUAh4x8OJbJz5GSK3WyCWbgvyOqazYDx0vCzUdqEbrQGfaGaVVeRrSy0X6b1
ajDdHckWeT6zKkkBNeL7+iFNDU3j0TNYpUPPRwjQfyumCNcRCb3Eup6wAqJIYcyN
r7sn1vhFbBsxuXejukiDeX1kHLXsYmWi8Bcqt9rdodnYFSfsgwmPyPwztB2NG6pP
FUQ+nOGEho0cJYOaSG0vftv6D71THuh07Zx94nv5BZbgWRh9YykyZPXPDSfsl7Y4
/Rs0biidCc8kYy7CZrwzi+Eu9mDg4s8ekMS/NusodEXmPCV3hRAaRk+KOYulz/z/
8y5yX8zfbAFqBQYmJGeIscTD1MGT0UFN/FdHPbWsAZ14jyKqe7xHHLtKFh1X+Qr2
lvQrSjxuTTCkkYU5X/8WG8ed7idheOz9xWSV+hJT4KpVTJ7hatqKlrMMVIsyjQ61
6FFjBI0Ksk4+QPooyDrJnZ67+ePAoNPbWinxG2FwZk+L3xgVWxKGkM7HYKjrHd8b
Zh0slvpvgKMG8xFXiKi44NjBJ0ExnE23VD9Um6XCxEqiLxX1UMcLf69rMFw2xsyS
qNePydDHsQsqJG++hZRGBre7VjCUPOwLt98TjtuZOBfKE+3uwLJGbjrczkTMxDUP
USJOW4wOGLTwd1lz3UhINec1A1gwoCCRXPIGWr5aKU01wDmTZ0VE+1eS07401+sf
JrVQD6eQiOHOiG8e+jud/zjShJFaULmyPMcyQTJeHuLX8sgRisEfTWCDRq1j34lq
oJv8E3ZqRbPrsXClPYnLaGT0OKPdNQNd1bm8KeX7xUx+eVGU6zPGMTAeYpgIx0GG
NCLXRiQY3xQ5X+LZftHOUgowNgM9eBt7TAE9Gc6gs2ssrnrexkru/saQIu3fOTWT
p2PXoquS5JAc/LJ8Km6hEYNHBHoV9A7Q1j3+g6fmK7rW1ssNVZogaZpepjkLXlrg
4xPyNo9GR+aCevpG56KVVTtYFA+r0ahvEqFGxn3lUBGz0Ujz0MKYic38S/ZuivhG
AwbEdDu+bIRrnAH7VCG5T6MdthAMu/k7uWnDVYKHuDqwheMRDl6NNqefKVSYOSWl
Nxr42AD2n5kFOFxeAsgt4kypfFJJryLGmSREStAPsojqyhU+Nsfavcjw+pNJcAcR
reryAF3cjWX9fmohuW7fOMJd9LvlvT76uq8C7Kfm89bURFsA+AryeIoTMSWyc6Ex
YRR7doCwQHsPYfubXRJOJIMXsWuUKwYLrp30ejXsS0Ju0ojxXsx0Kk66H75MfGs1
y4HX9oStE4Q/nD3xeXAZx64XZZSaD7sNwDjIU9x/XZabHIVG2R7w93J+8qElnb/z
gPNQNOFogZ+j+P1RvQRZj99ELt2aOgHq9wAGJ6QTxRSIU/QqBFiH61qXaQbDjTbh
Px9UXX5uw5+idIusbwYYnaj39I0h4p6NtLqd2MAOIWfgNyBZo4ZZTJnOzhSBeuJh
RPIpzWk539rU+taYp9N135KBZOteDFjrUtlu1HhtHLkmgI92S+gU4MB57acM5Uo0
Stf654pbkHa/LL1WqJnsffLY30jaHfbJSm+4aMaDe6GFtuP9OD+Zz9IlptU8pplk
q+nZUvxK7XtdttSMCmHHLQ==
`protect END_PROTECTED
