`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1JYBTSVeByK/S3ywyIx/cKBWnFc5eaNR1Q7wn+0K6HPWj9z+U2FpsTD5EIo2U7Jj
V5v1M6ACLK9bp565tDgHV+LpqHwz2/II0aJwgiLsve1lc4d605c6kcMnArGkFF05
0shdwBotKG14Z5hbtraiMhOUP01wwg7vcNyb50xFQcyWGwq9hmvR5OCjOq4PQUBD
LqqeWGUKDPq32/kLO2pWNaPT1y1U+HKg+J5Jpw/eBpxI/+GaRFxv0+A5E1ErBsGY
p0+IqUFyUC1ZqXLZBMxSGMpqxLmHRignu4SJM+aRwJWKGSWBh+v3lnD0Fq8gEoj+
c3vkSsUn+7KU8GsmZem2+oY3yv5zvy+f3IGwVGk81P/E76X12puG8g4uy/z6PvuY
`protect END_PROTECTED
