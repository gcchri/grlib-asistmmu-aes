`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F1MsAk5XPFvAA/DonTGrNAOBBAvuWi4yZDbwpRPuOvdpF+eEenUamm3uZcfwWcbe
ShJ5Z+Yc79+pO6nizfPi2A8jaQq9L6W0wRGqDGeeJ14J6reZYbbLwMb3M8lvM5Tw
p24p/Sn/QCbouPLGqfHPLNZHIlLEh/cM2q1WOPWKJmP6/9gq7zluOo6XudjeY18W
ZhMz/6xLbNknlCMlp0NXbERdKC9hOVMh7ER9zGEADbZy/wrWyX+ryqK37QMRLArs
Qgc5TeRGfinh5mxJQ+76mWcpXUQ/4PWESNvFNWpfDrLp4O9MnK9YdENE2HVruDGt
2Ie2gkeF8IiPzBVxmolcntTyIigJ2fvk2FQoQmQpc8ixKgQWp03GCZF7VO/g4V2W
yHjD/OujEfUpdnSCLcp95L4XmuLS04jpHhxkvHgpDFU=
`protect END_PROTECTED
