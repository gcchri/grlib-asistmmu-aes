`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5fYZuhRPZP5JorXweGGwOuP47Qi1ckzC2Bdxp6UYKUaeD063MKCO/CPbfZeL5db
M4Ru+5OiQ8DHBU8oecl0fVvsgzCy3H/Zudo9D5PLkAFNqjHuRRwv9lRCgECZPRvn
WAcyZqOMgMoJs5wTOmp25q1YC38xEDO6nn40yFiOYlOrDC/yZry1qNoec3qBkEbp
YEF9DiQPavLOy6XwRIbdZRXujQeZTYjsmiQd4HofB0QSBih5xYa1FYf+VjjTU8JQ
YNw8b2KKPoXTIl/27gqN45vCZuEWwSuootypFRn5HlQiEPHwUGAdTk/hsHJ/ijeR
2NGF2wFKXdyMZ0FdHq08Mg==
`protect END_PROTECTED
