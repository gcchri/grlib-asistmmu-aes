`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iUGTweb5QFyASW6NTlsKpsDl1QLVKyX1pLG5Lt/DIgpK7r/Q1Pd43Hi8jtMKT/xR
Pb36Otyq6vgMF/N37LMKdqjaNgTXZB/981s4ps09yAdfEpZakmd/y0AzsXFQYaRG
2547DkCKFQnN1I9BMufj836cO6PttaGzmNzjyukjw+2uunlCwCpVyubICi6Q0U+X
urFuaYow/oL51p/A69IRcJIcPjNL76BjdGR+Dc8yZBk5hRLkRdl7gM9AeSJU/GUB
MASav2xflacgZ/xdRua0eKgI7CajNoyzEMfm26crv8rrt4tSd2hkgDsTx+ymVSe4
xcsxMBjLSYNqJ6rqnButLkXxqKISwpFc7NUUXEPTWUwKS7/ljLQo5f0F6zBeC/uh
XfbBvEJK4mRcjLqxxpnqRG8Qup8qqF1VXoAAVEgBKtuqiNa6yua9mexEX4JVEokO
IqSWl+2fFcARIk1luiE2sqnWyXC+jBZaowjep3XUY+GUFLwLSXQ96z4ansFK/f7t
xbS+guYt/NN4NUjcYc13iQ==
`protect END_PROTECTED
