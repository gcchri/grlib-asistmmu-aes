`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqoQ7NM9N3CuXHLnmVRMzozLyiK3NNbjJ9L0M3o5e8FRDK1Vd49+xWDVgWyHmW6P
+NWL8nKlclvc3VRQBXB32LVt3oZ/+apGfZMSalptByEFGb/4L2D3P0ovAV+VIf83
p8DiSwMXZ5zUIO6viyjaJMNxG4LmbKvlN2l1415G0KoIWdKyXwVtZkPlap9aX8kn
jmdwBe6u0qSCA3Ffj9ORupCtkh4khlCzxEzxhmw5dGhNWz/gugXo7cHn7rmwDtOx
898pEKP1pl+y0S35cnIDxsoPX2mDPP7YVQ8CNAzvi6SpWTJarH9QTYJUAz2ykyd2
hZFKwU/1Fv1u10VZ7hSbDeEOosQSHg48pd/4PROnLK7o/GuF3FFkZU5r3ahV8A2G
s5RFgVoBvrz0gOltzBK6MtlNgPw3LB2CYG5iK7iP+1K7UMRrNXuwevhAk00pDe77
CgZypFpI4MAKQYYNfmw75G3RrNVlbnKT1f627Z4Ojx5xsbwsSmSu2FAR2uWKPKew
`protect END_PROTECTED
