`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ia5hHCXnxsLIakZZU239ywRSFAKlfsH5IPoBuQbHEhxdS3Ajs2cAyr5QlWP9AOkL
cGE8ewzApH/K2or/wK/QBAcZSO8N0fIzpFoNt0LUWrho+GtWw+AHGq8bpa6O7iUe
PxKkEVAJIfUnrSjd6nHbWI5CftDyLCr0QIfvAcgz7mY=
`protect END_PROTECTED
