`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6zpGYyxXXpUHKtWkIyHVxQDS6IFbqSKDAZsWmn9nJeM35ajTIF+BQ1GAo4y5PD/i
8A2jlIoHUlL2f50vudU7NSt3ldTJr9miHch+eXehj7jjzzbgknVnJupSM8lacjt9
GrLbS5Urak/WOLYWfePfoQqTzyRyB3s1EWKalfgLHHFmKHSLp1Wt4Q9zyJeisTzx
pW1vUq4wvOD8Lh0jk0TBeydZ5EOf2PO09tQZYOSJnzvoldKsdvEveGNTlPREK7Sx
2wH5eMp5wOYmZJ7+H7GK1FSD9AjNkx4ryQjjDRSTP+ySmGr1Db7ShRX6fQImcpI4
ljFuOrtnBP3ScsjgTS6d0HDfgHQAffDHR8Rt5n7JevKmFsO6bXug1esNe1UV78KY
EAf0l2MH4lN+FXY0I/wBlmV0+roGfR15BDtxudRpxmDjHcdEsEwOKxsKrl4uf8K/
hgvV4AVwpWBG6I1n63DmRA==
`protect END_PROTECTED
