`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTmGRAY2Kr8JNIUnPd5dj205OBzlJ6fFCSvoNTHw6BtFvQhZF6iGYB//tWyDF/Rm
jYJHDRTM99VlWeJ2rfHoN4BsR4GNzcoL/OGyjm8fZ0o9pcdyeaNb0579wj/dxXgf
whCEGq/K8IKRXQCdncZ/pRonwA4j3TwOJMc1YJNsUHAEKB/dBDpuANGYAEp5nGU5
a+Q9m3mZywEH3IRZmkdpAqmK8WUTlWjfAOVFFz4Nx7P/Tk75EXfl2p/4R76NOVar
oxpiLih5+hbwaMxTYrQlR3m/znV7UzygPgc3IwLdgmuVxcYVEm8LTmg45q0Iiqqp
efV18RzlCYmcA0Iv4dQoMtgawApwJgAHcbtRxYoBdY0=
`protect END_PROTECTED
