`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XL30hpDW2rLFay7DQZl017d7d56Q0FL9RRb2XN/EYp8d5qY7GFcARdcngdolmpWK
AdWBCVqkeDwyDO44/4xsmrlYcUBPGSwWUarqw7VogODiTKnbDc5rPeFZ1J9bZUGs
o4gDLSnMzIoB+7auyMe+el2Y36/EpFlPNGCtApwfKYaGRs2DFv158V2MY8nv1m+H
twW9nBCVEtfUpv9f7ES7FRpR6BE1IzoS3xSl1FV0Oc8DQQaAatfL3tUsGrA+8GvB
h0uDZZ43thX6itbK3PB17iswPOlmVbV8OxwAS8t939K6cqGqdzX5ab75KbyxWrW0
2WRRFhxkSBH3zENj+mbVM1Tr/4TtrEnFQ4T4QpKg+SgDXRyo8C6Yb0323XPq8qrC
bWhinHw/xg4plgPOuse+C0YSYt7qDI5TNjI5/tUs0mvRrjOti8eNusXg2QI3mrAA
uFXrhpA3AEXbdv5d9f4KdOSdN0ACAcqq6YvhjcK4dJ7vx3B6j1ctx0DvhBQHpQBC
iPVfTkf7MFEpMCw2/QrSBB463RgQbUiDRKc2sxGttoSvk0wHvDgkqhNYR0hy6SuJ
crfHKUrWqffr4tIywXVpQOPfoDzKqdhl1V863C17Vt3/dKvEU+evnFaxT+SXwuoF
tPXtAb81aCOpyk0BCrHYgg==
`protect END_PROTECTED
