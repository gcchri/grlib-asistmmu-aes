`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PSwDcWkzp9Q65PRfcYxIxr967G+afMB24MJ81ROozAyi6McTUagcqIh03fjxa2X6
I+ftCedkDAOYzxUw+3TGFMYGpRDNBf3YTfjqPoXarJ5lw5wTSMIBGzcS/+zzjqgA
aZ9aMsMlYKm71edDzGXjYEbx42tZBfb/2BwYapREnlYdbMfKPhxjq2MIWZAcLXnr
USrgP8XJ9xOUZlyYPG/B32QNv5b/QLWE8czhBdqhTvvN0a6niOnh2TcqUXyUmBbQ
wVs31TqIYOK+d5SXZsQywHbNxYxXbsuIX+KOiPgeJn4=
`protect END_PROTECTED
