`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDRIQRAt2vHlWZhZuS9eRmZOILaaxb06vX/2/bOX1dpom2oRsscLmHdGlm4n1Hbs
C7g0CJT1bNs5f3BDChLz0LDLZXmepy6fTvobWSAna2QZ66GNJYhWhXbe8KrJa2VY
TFYRQ6C1IuSVC/CoUZgdaGGyNDM9+tcEnZx5LNBusxmNg26mKDUhVA5uQt98neZw
E8Xx+0lhiWlwWQuKnTNWKXt+8unFdv+Uew8a8Y3BCJtmG1VncMCpD64gPrFGQohW
G71Z7ICBeQcz6t6ieIjQcBGom4ktvfbJZJ6i4YDAR7vbeLSQtrg6QeHbcv4oaKJq
ERkgo1rqYIwnREWiLq2MvyeuK+VnaDkQpCbUeQyckDvznBEFkR0cCAYjns+knQbz
amQLr5i0VFqdmvpDwMrLH5QyolkvSBbLEKbTr3FAAMuJsAKGQ/uh8Q3gYfXORGuv
PRag7G0hRvmnXneFnsvj2RkuYQSfqrdDJ6l/pFczOGQ0nkrQXOlOh8fMyuE8Jc9G
1cBp8XFZRjDwQ9mj1GX2kxZ3nYbfTYNCsz46PKJIEfOLW6S7Q+EA0eqpOkLDLQm0
0MvYN3wMMjkBvturTyPzgGkR8j7nmBzIhliK60nYGhcj63e8PaNzFofjz+7DuyOl
v5wB8EEX8uCAH5Axz++IMHVZM36OOKySba0k1fS5z38WKIaEean/H1LSSB+8Xt8+
/fc3wgvpSchiL0+k5caE5msNqYfRd8eJMXvnpDY/K3lNOM3CgJeAPzjqi2TYwKpU
deZlHv5KzKJRwkfAHdLnUdwm4+H1FSTbWVgvJAvx/EyTlsQcSbBxIl5A97wBsSjd
X8uPKzAmxCVav7LFBqZ4ecL0eOfSis1Y803dBL/B2Bb5gM/c0R9USb34uB4Mrc9a
Fu6Hs1xwNPRH9fwvGwTRWuDq02RnKQLGd+GwhVmMsp7gH0KsPM/GUl6S6caRjfT2
yFUqLG53n+gVyOT3xJwULdev2PdF+7P++dY2DvcMvqDd1l/MRJ1jFWGp84YyO1y2
pBSePLLK4OOmGfKUiZYQNcjSFnwEY8vFUOI4DMJDQ2M1DIcxNv9f69qeNW5q0CYp
1J8Mdbvks60NnoFFSbRSMrHFDLI33V/exDI1SuH9GItmUjBqRDLv1FaDcpTBOhID
Zj0fhvzKE5zydjtlOm7U+Iw53LRP5lIKOYaixj2X2VysFmSR8Jr6AkGRXxj8qAGZ
FxccVNgp0BszenLRe2yiyAYEzgwgkCoK8RrM8YjgsQq33EBWuWCU3qg+KZFVLKS9
dUm1KHvXzcKyxkq6EWRe2Dnc205vovlP0Et8+7PZlvTnhj0De9SrLzJDKYs8EUUg
16vg++Z/ElwpxV/4c4QAZGZRL+8n+FEJrsV0+jgHyqo3nCH4Oar0ZBCrZU1gFgB+
Cw8nq7Ufvuf23fC2CgC7QIbbGbh9AWkub5bJGLNbW8q7yRjs28I4dDxSmU/cUAyR
7GXFJDpGGrqpRpZpXul8Jrj92aAJZqGNRVUz3NKWeI23JCJNVJhKoTDHNe1mtCPs
4KrdjpZQ64qJ0wqwbjREnqsRiqFlvpkGor8EmhVjlcRqAp+i50PUaD59p7nn0hI7
G4jEK3a4F8tooxcSKfX/nUi9Lwceyuh7fzuTNBRVsyGq/ptvoMxxyi1inaKxsNha
t0kaX8P3WKG3dh91DkP6eS6mMBWilXlHXLHdvcBpDD2T2habhD8WqeMCxAfRsnPj
gDjT/uuiOWMe0bNQvO6A3stguQgZx2Ve+480aQr2ioEq2/v160EmDNgpiGAxgU0t
GGSG/aE8UARyrHA9xj57SxLMeYeY3Csc9cKZtSe/SygZ+2TzFP/cxMJv+yOjshVZ
mr/fCdRiEHupLgwULddJHrp5HYPB895mlV+azqRn4CscxG5yYpOWym69wb35ryae
OKSoNXAw4GCfqwMdggKHESRwj6dX7+OLOg5nFW7Qp5J+iGhYxoTWFNT9Vm14moPH
Tk8u0LwtnyTnJg66SD0oCifn6HIKgan9eMzC31MFnu6PUSIRkCxTem+7wwkWbySh
rzXhJd+ikMk+lF47xpjo2CxMhJkoXYrgE7cm5SI/4yrLAkX9/8vdXdMB+7Qa28fu
rILv1Na474P1e8q+Wt+mVclU/u3gFfKuCwDifq58H5IoC9Z9k9jXIBznwsQ/5mVT
NxmmqKH0JJ2d0EjAHWB+Jec8ZZ4nuOOy3fsPc5Bh1KOEFgJjsxMPokEQgIu6VlI8
xPTGEiFbFVlVfctod2KQGMzC+67IsRENhoqD+4BGgiQFRsgm+kh5elNYsfDI9F3d
TWv/ivFR5eXgVujspC95S6pQpi/oEH0VC7QVKouHWftM/33k3M3aq1ABtFy3/NK8
haoazVEcWySR2ZdCqzYRX6NiN91OIk2qSdXt6mRfBhCBJ6cbjt983lim7eldqVUB
kw+Mg4llOpI1PqbWJBYpaFQOdT5sZtNlsgU8Q7A4jFoD8SgsYwB1rjxrisUO8sa9
cSTtHMu8CZt0ql71jICqnyAVtsGkHIc7sXN8Jkl/hVyUj9pWF1CkoK7kl0MWL4yn
SRzQMWdFDa6KNFRdwg0U3UjEnVusaHIyY4AWuin87T8jCz4TJRq17ID+zFMOrTdi
nVl1MqWEjMKB5Qr25NBq+db2d9lvp3jZrusCrr3nefW+1kNUKuaDOGZT/skF+1xT
Bm6t40aPgXB3Qt0jYT0UxogptMvuAhQz41OEs17RFnX0oN1r7hfguBiBoHeGDzxg
2dB2gymNSFOaP5Q8vsNTZwOaTcl+JBcJpEemduN0h96EbqDP/KIT0WmrX0Dm989u
LX/6YNtxDZsmlGs+roWxoaKs3r2pYcuriJUYA9CS5tiij05u5I07XyBa+ho04BmI
9WTOrqlM6Dj8VXEGz7nVqHWlb1g6LlsHWFlSvI4XjSjHu+1cCYEpUgZnuIhx+4OB
u8DcNWLAl1Ewy503BrRZaEFAiYPX21Myk6DIovnHBiaIgr3rukGMoK/+5d5Thdt6
oVsh5HFsCZ4ZQe+6rcjeOd1AnaEzM041gKN9EhliVJken+LoLT9rv/74hLdBGXw5
QDNTJ+1wipKveXcthWFsKAz2dRrjtsjqKn7UxG4mcrxSyfXkJRrawTC1Mn/T9wUd
9RDkLVP1o2gt9t6W62V9OkrpWC3I2lgO+wEgvN7/HKvgU4ibpNDfVqH/WXSnA9pm
6mKLO6d5sVfJF4jDb+eUmq+4t04qDR8AQNPk0/R0nWnVe/tXj/UyLphgd2flieEM
S0LzoItXDkmxa5HqTbhoENDJYeGrcHzO4qcd2w8WKm7rR63XQrdPssuvnkf5IxUZ
ZO0UXYeGy2ekqVpbuW0yKwey8mzjed2g+QU9W0cSU9GbqIZPwlR0k7Qp/QZRqR2S
yIRrm8XcdVbcVcSZ0V5AhRNdii1vnfWxKVguZSKCukvLBWbtT5Zu8cNPjVmMUraz
/X6o+wLwKCmA+PO9oDejtPb1d63tKTG3YsnNzHtRDPuAcSLN8W9dLB1emuqlmRiL
fFYi9MgidxysaEBRrOJJB7jSW3rrEa5IZ2Y5OJM9SaWdEcFlN+xZELuKFO/genNy
okwiSY6M76GIxaiqcJfNQ1y/PJtv4GhKIO4U3PEbQIsqaKnw0qBWh7yq7FG2FaG4
NFsZJZmUbZwKkPWy3xSxddpSSEEsPi32IRjee77dgfWhJ7L6A/O6byuZI1O3cXDs
p3/WC/NgJtgptx14Eb/WJfCga+hYH00rDtgJLhTCXBcgNKUzDCnWlhF4H7EreO0N
`protect END_PROTECTED
