`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTnem6I+bR7WeFrSX7MPa9/R/uCtsVOj7r3OMmwnxNb0w6hz3iA4GLUdiqrj3orR
7v3VJgvTGJKS0s2G5ejOIzOBDQrlIjtMTqDOCpulKpi5aV//2ZMm16bX/66yFHRG
vCDvqXDvDRN23VAsXvFnxPO41K4rG31WIlld5fE8wZ9agZc4Nct/hL0HiLArzI2n
+Z2HdRORMYk6X07O0CUiXfQRKmQQJdMbCNiMM9KQNphkV+ygp965PCGt5NfcbHb0
ZLF8i8Ecx0xx7ABLgl558+RWnrJ+nHHRUiElSAZvDsNL7h9iZRC4Z84nufBUyrc0
iw9vBQUcxU9+3u5C8gATqhm+kp8NGAmAkxMKu5cINyJM2voE1YDVigbtufTrKcq8
EIPw54hO8CStQkn3c/43oPzjs/nwJl2c9Xv+aBP3EKc3stkG8zqTUWdouQu4viQJ
WqwcYpy0we7pN9rvHKUwbVFB2s5zqiz+A7g0X22fW+OYJDA/WosxKEZ88DB5wvYc
`protect END_PROTECTED
