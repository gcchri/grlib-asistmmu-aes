`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+3rCT+QwaXG18KFPjijJnoYQ7nDoYTMAzPhqXbzYz3R919JZYmTMuznQzfMHFKTH
lRkl1Ff+3mTEvhcaFpQB9wGEpAQ7qruHb4i87Nv4eGvh7QtNRctejBbE+6H+S+VA
DQ5m/vPiBO1VYG0OBkF3a9nvMBJ4Yc35ckIaq1XLNPeHPi562AW3QjkcSKS+MBzA
8w/iXTkf6RVPCpRxZ2AuHO5rKFzTryaotXQ8qmOM3m42/2RZ1uk4rYVDb5CKKnSI
+ief1cvoVrNkBL8hVpewjg==
`protect END_PROTECTED
