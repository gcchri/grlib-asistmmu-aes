`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kY1cuk3Dycy0KMcPHEQHjnCJJdB11KGioPClrumxchG8A/ha1dxCnVo5aFwZj7K+
AhOOjktVPSAR54w0iTKhscoxlV/mjrn9VicKurSYHEQK/uDgrZQ1inFb4AxO1Z+2
nxJ4Qcgck+EFWimRs4jDXqDpVmcPFqXvf2u4alz8wLJ4ZYfODME7LVhNMGjomlTP
Jn8IztB1NsMO/lpTt5Gd04hQ9Fd29H+s+5UPvi1s/0T1u75bf2KxSTXpoCHlLYQh
pDPQvkeIRoCQyXTo6QVNgdpbYucdLVZP/K3LVnA0Kw9pDvIVCpidzYFxR/igHH/0
Xj4e131ygefTL/63vmfzrg==
`protect END_PROTECTED
