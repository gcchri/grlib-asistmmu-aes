`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YkUKc+bL28KaS6POzFxjDeY0Oy7TaW6KmR+UT6pNXc56iRxs7yjqJwj3YBGsyE7z
Q0jy8zgRMhF2fjkHBQZ5BPaLqMU5RtKmrCodZSjuitpSGsrkNbCnKab5FL6H0uI2
59AyOSEcdgLSg3mAjuUbetJOP1l+LZN9n9nNNJDrJYpOrb5NbcpKNCGv7nZO4oIp
imtiTs4Yjt5aKZFDFr7Ivln8djK5ObDyizac6QhygLRMVLakbzbl3EX2eug5tHGG
XfKFwmn7/TZIWWdwRkZ3INY2MTdbMFek2nmv9yqhXFAy0OnxInJbuar9H9J0nYBL
OYmyZjwGgiYryALjsuk5L4tspEhUi6LbmnbMDkeeWKKxh/3uLj8KwfIymKDw9KWd
3h1bSPtiAvxQ59PTeUanMlKu8y8yFMPS4Zed20wFwM/Kmyrm5HcdGa4HHhAgd/oU
`protect END_PROTECTED
