`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mj7Y6Hkou1QVbTyFh0ERHLzE5urs5BOPkSI6EJ/7NRYZDgnmY40h4DPU1TWtLxY0
jfBAhyM303ugOK0gDFBMRO91W5S7BSRnvpTlI/xIvupuTka6z2rybVyTEgwyyqgS
CLCd19W+tkwO/NJkKIrSmpbkh2IClfK/P69fxBNL7yn9u0lPHkiRhpP9qP6e/WkP
YHzdBRFy6msja7+4RHJAUMmwP3IodCJiUkja3MR6KH32k86LrdQ1XbRA721BURP2
KyhqwAxreXwX3274hKL+OVIb5l/M2InbIS+rnqpjd/N1rrS8PE6SQPHda7kURUOQ
ksCwNI3JZdHCWZoeQOTBzpvGBHgRajYxKaPv/wWd8L3iTYD1KVMqb9SFPJKAp9so
WtIxQII1Qm0XIQlemq11DzO/YSm8GZ+FTO/e8T46lrPMoI1ObkmysVGNiOX/naPI
MNGR63RhA8eKwIHKeykqrPA8wGB9B77+6ckIdLKiGVVUBsG4xAAV2fS+JrU5Ygx1
FSyYYb274htO0H6Tz0ojNyz2SvCihHTTvo/aeak9/YYc1b41D4m+mzB8+FBSDAqM
y+cpo+rhFIwIIUqWVhnAgQ==
`protect END_PROTECTED
