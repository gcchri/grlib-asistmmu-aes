`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ugYYxE+v7YlcPZ8690z3hhjpvFpC/moMu6RbEu+hVOMPLOKZauDpD4Wn4tgtTmmL
2B+pPaJiFlyOe8lmbzCKhBj+WT6gXj90IR2ikcVIeUvG7wS3rX9CjBGPQt4HKiUa
7pz8h0JX4lDYhKItwxUTDjBWFY2pqF6SHmfn4YJ/rh0BmUAwcfqjQLT8zi6cJ28M
Fh52OyvH3+GAuVexjaYmveSfF5ltq1DaZyOr2zRd5LG8gPv9hp2t6atzDvrZj/T2
teRN6AiF4HXnONDgAAQmO4zLk6FBcNFLdA+CRos+TN8=
`protect END_PROTECTED
