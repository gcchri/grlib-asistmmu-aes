`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8OAmZQd0GT1Bqy+G25kgiGNB33ZfrxfAQx9/Jig3NeZtHoRMjsailH+2UNY2cU7
qyCmGnuuAGGrYlxhz4xwi0jOq8ohb136lbWLJNRmIQHmxSD4aYaTTliFm0zGU7gG
Od4E8/Erra6VETE324+v0Odpi7k2VhckyWBnF3hERfWOZTIuAoIRk80ljT5OsL6F
5k7DUW8A6h1O1Y/wlFnG76AxI47y/zqEhUwIqovkY+dEWsdJ510YTBfQqUrteFRG
UzNmPUo9D/W4QYra31kp6qENo7WjkmodvfTmLebIvNUhjsrwwzuGes1btDOl9iqV
V7yvs9l5VG2U3uX0SzzqsNl67zd+ng6l9e8hYLV04w8CHxmowI2IctFuKz+p9R+g
0Mr4shOAWAfaScf9wlZdeKyLOGWP7SGrmInBnczAg7GkUWUO1HmVaFS2a0Vg5ZJ9
ZWsMH4S8F6SkqjXck/sfBf4xUmA6qaEuq6uPmRQOn9OhZB6Nv7lwhorvgXVDAKGV
U/eWNaK2zFJJP2sfylljWa45I7tFj1uo6CNYMPcdU3nZLzVPCJ+9sOSVk3+1l6Rr
WFqHfBLvSfujpLrh2BfzMw==
`protect END_PROTECTED
