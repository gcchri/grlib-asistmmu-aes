`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JedVj8ARdBnQYJB8N/X0dBRW/QGQ+SWakMqCs+2DLTQgAYNMQGQI2CJHv70wcHe2
7bAdPDw7jr165iwu/rD9wH4x5WZU76JIonLBea6A5PnMOm6Ttl4cMI4uksNJQMlZ
0MoMZsGYDSNGmwHaNa4n8i2Ic2kMVDXmTe19F0iH1tkgEnrNUo7j0SAG5a7GQcIe
w6k5hx4gzRKod7cY0HoxLpWILACYi3N8Da2KENF+sHyrsv5iEX0sEaswjzMZoC08
sh4NMFAT1DmlAozeUzOb/01DtoZrLr1tMOyjMKOpapdrrBYY7+7LDJbxy7/mgJJI
l++zU8TGz8mU1rej5j1MX3fhLvJGqzZ1yVDB8bf4pCT+8B1N8i/CMf9T5fEgQxGf
4N0mzQL6dL/l0+lvJkd/LX+iY4Nu+WuqCNU80CbTb203YxPR+nP07sAAyJuxq3KV
A7r7REiU90/lNccnbtRKun/yV50Of4GIRsnHkaDOkDL47b43tYy7H1RPyTjyUOow
qbghZrmw/uuik8QNJGYS4fhZKMGkIW2SQ3pZoIu4bZ1YmJ0yTUrn9g1uM1BmwUEG
e/3OT+2cAN892163FU6g9T+rpuVjsWgMtdHndo3yBdisK89IkFQw8+W6Rzf1ba+9
vpG8ASwZSxilfhhIFXmCr0XdTQIeYjcqtnj8dI9ZgapXm1Hmt0rQceaYhsJ2GIt1
KhpHe+3w2pgPeyL5POYf2fTbD6wCCMWNqc7MNZOOn+tJOBKF85Nx8TLU4F1rIqc2
6BaQ2to1RM7KK5EUg9e7c7mIEz8SMUW93LnnNTNKZlxOB26PJFES8bwl0WQ2hoVB
wFsX92dZOfTUbBK4UIKL/7WvNGt675iYQntOiNOhGhwiZfzO85EALYF0FKA/cTFY
/G2jjW/GSSF7ADK4TQoMkHLgxGtXH7v5G1RPt+hPOmn1AlLt2a5KU8AeSRXR/p1n
UsQMnh4pHFt9ejZctrEXTdtQTHYz//WvQ4yHZgiLDTv54ySvgac2z/eQYiztU4pg
CIvHlUkt+5mKTZEtFjCwDirLlhqt20IcO/8G8jkIND8GrSeWC2+uSkawH3tZ57yg
LemoQhN6WXaP0BH36Hkf75wMx951CQU0cIXUOJfQX5A3ebg9M49cqfFidOkxiL1I
OvwrZgD1Km1pz1Tn/FJhRpK6dKjEn//7UnH5fTaRfq4kzN8WQ3lPwKMxTbIZ22e5
ex+XAILKLVEjt8OsVt4POV+cBNHJjjVQgZ46CP+eK6IaZF0TOsczrbxA3j76LhcT
e5r3rfWO4xHDfVSv+30Uk2YuPXO90Qij+Bv2EUGpY+jpdaoyqIQ6nlMM05js0ZY7
pWYz0mlKwdRFzcB+Y4xXTqGwiuo64ZWO+awaYumHOIFWhAVmBnAyREO3Qijjk2qf
9yBanuPTIUrje4aKGi/5sK2YupPoiymKuNc9HfnnIR0h5hXxQtJgIsF1su+6++AO
1tGRBCPIbv+jgRAI0/oO7ZgIbNuyYtpo8SW9zF5QGdGD1pF/pqUgUgJ5LGMcKCd4
1w6HcCnMHU4/NJp6FymJSTeXXzpNVzdkIqJ9iAcdB1pWuNwgJjfBDjDfdu4tP64K
juKjkGAQlbnjIXZyQKUE+n5tfIlxs0ep2tKbFz96+ZSppQpP3xs7zbYPKcRMLvn3
r9iX2oVsrRNKFZdRvxBciRitlKdV2ChuerxWB7yJ/xIGJ/HnYwz87pfCwCEGpySt
/w+tDxtSXgU0XEumm/a5QP32sDEiBTHXRgmlOVS/Hwmq5vJke51P99ZjOcc2Mpbz
4I6vyF8p6uZb6UQQ5rkFGqYjqQPrmrwM2g14qgTWKtTfHmS0s9xhXRbV7dA4Em//
+FwxAoOJVtr7O9pf2kN7jrQBva4vPn7e1R+kqHaT06RCf7TS+ycz14yBLm1JJcud
xxLqRQ6KAWp7OzmyN/bLP40T5BC8tzrVgyFtTNN6p1sAJpYvzhixtwdC0pmKaNQy
H7GaHfGAJ+nEULcS7eczt4GrQ/3Ub2C8sX7plrI7ujE32TsH1zx1asvAniuWUSh8
HT8Dd/2XN6QseFI7NQEXKLq3adjmS2Iaj4nWJ9zlnGHI0q/SETPPcLqUCDEz59GN
4dCFYNvTuIRy6URvHQtBbn8uEX8NFgzswq5PbFO8fCYXZoJioFr5VxDlmR09fMoj
Vnxtha67k34UZWJeDoW23sjDQFTmN6wNBmS2otsNkh7ENj70FZsGGP0lJmJINkkP
HzKw5xKz623ufo191RwCWOxLR48EuNx3b1yBr4S7kSfEI2g/9yaPbDmHhnm805pF
TzwVoNZMjT4T6l+zSWHo67u8rytRNHimw4E8UQn9FakK9k7mDhASNmOCQuOljlgB
fQ6ASGVw2ZmeuSHkvuNtEHJjfQ+gY3+J/EjBKmO3GPLPbl4vfrmExdatO3oSQymA
t5/d0URjnWOYC7PWuOiPiSh8Fu4t+zB+d2mPkA5eQDaMehnTSuQ1oft7Sh6CTIT2
HZ+evii8FKFb3y/Dp8jUjeDqCW2d45FCql/P07bGjTrQLeZxkfWdITwpnVcs7wq6
gfKMRAHy/VFHJE4aV8VXhca2o/UHUDvyNXNfunCF53W3yAvAicU4LJPKemc2zFa3
6gHeviTbOSyuv3fVJQneJbaDlxA8S4cTLIh7goWxUYx5nWcleUphxHTkwigs+Sls
NkjcD6htCcWOGnnFODu+gbrFm+2NcwrBNQGtf01tf1O3sihRaTD+eu+rglO2GCr0
+TV1ClujJUeMixKkQXdIYKSY7dJmEvCc+FtavKnUjU6H9QJ+QfzB/ylJQMwWGgFO
GZ6ubLEPOm/r+7ai5oRmWHm08a4N6EDkReDGBxnFHnhwxd3af7oGi2mLhqape/Fj
vsIwwYcmbT5zhtoEWwzK0UbqqGqTF5XFvijF8cOjcMcSpAjJUAwVI5BAzng5ntev
WC5FfKbSM+fLiGYLavbQLLeZtYpqXaBZ4BX10h7PkzWfG2mArwWofRu04jb5yGhy
eNWIdilggV+JinZnWCSEIlIVbzxpQ4Wolp9RKX/UJtExeoaLu0oogSM/iqWsse7L
m3V8m5W4S380YVUkyXwsM1kcut1EwjUtB94hf9Lk6aeh+WiZj5e9zUbH/VhAtp+0
IouKPAJVL8ky8tPqZR8PRQ+FBz7IKaG7L68N1khuR2fiP/pQ8kX/x6hxQC4H5aqP
SPxoV9pnlt+sOMxt5Xa310NugyQQkE0YwzewPjJiud2kzpIaoE3d7xheA7icgk+L
j+d8q5f+HVkrFV15MRCq+V1fBECsaOW+36HmjRIcS8HpzkAeqKkWEe9UXSdf+GrU
Zy/ERKQXfg69d+5PoapLxqfO1Ag9qm/k3Sio3/28kKbVlEMblXTJ/s/AxmSLd3ke
xz3zpelLIlPfJhw9muvxvZHe41jsogt9Fl5Nn5q/pUvVeEfPvZU3OgpXT29PLUAA
bd/fmU3B6rGWEeMfKbj9E2g1jpI6G0fl1Oql6bLwLF+Kxygo3dGf00X2Ozqqe6Nn
gECsZmiYwLjxT80+9EnVobKgdqvAF7P7gd6f0hXmhOxhLKTQzIuMEa50mP9ipRBo
Yb6B0W2wDzAoPG+YLONaSTGhV08vPVQINozxvgoKAuK9UpydrJ7PiG53mKKC36kK
P4pP7xA0hsT2ACf7jDzN+x8ZZ1C732vqXOL45n4dUGFDeG5sYM6LY8tR00yMUVJ6
VTHdjtJWow73YUkRfTxe+sStp/U9Rj7qEwF0K4x52UX+iJN59vrbhtHAV8B+Izqz
WoRvYubo+01IZMa08qUc01+YQbDfaFF1ZaA3LEqXnz+5FNPRIsMpzECMMRMyMZ8a
OYNMwURy8A4S3U1FmadS30GZvi0yJOu6UdvVpm4NipfUlE5wAB93KgPne/eONNeG
AAjFVJsKZop3dY1YClZJ9XbiXs6Nku+9V15ePegr6nPPiniOVsNk6M6vn6KXYFOi
rNwQwxjClVimklEA9NEsyNI6YSDUAO2CLiF1ALSAGEVgJp3VN9dADG95C4d0BV6N
+UYDDOc0pWJrJyMTDhVXxTAXb2+bj7uhjZ+bYcJBfjZ4Q3mcZzDc+6pYzY28vawQ
GtCH6wDxPgEnTNPAcd3AXxrQT2smOjaA3xzbz30+UY7MxiNumAcRNVmQcL/gw3cw
fFw4jUjBe4cVAr1Ek5cMiW64L4x1g0f7QA3dqf9AS2ZUiumfaBhuldT+r0oyjjc9
lCaniI3WqsCH5oqxq3QyxlLcZDvzkziHp2xQL/3fvm0NPaEjXrru8aARdoZ2m8Rp
KJr4+u8lq73iQQIymSfSEgeVp/RRb5DDuzarFqyqpLUFWbjh2KUK2wtZ1id0+YEs
Y5NXz3hLQB80CmcAMqw+zWKiMyHyd+OcrM983xNQqsZliVHrAf5CX7jvZrKXxH4H
la1XMfl+UrZ8ymG7xgFsqvlQWKm3PTJL32bVpFrjH5gEoF8o6rGxou+P3lT4QkFs
J1/LJaHWU2D9x1Ptq+g4CfkC9w9y+Lx4Ak8/90YAys43SOALOoQAJMCJfIFT62bn
Z2Ft1A+MvmMTlEAjBT0rvX82A18nEiUXUsNFv+QQwbedwM2GxRuUXf663dTSMBQg
mnfIe7goOFiiPvY+F/xNQBWHM8OFWt0EGimxrHYrDkhOsu2OHng4GeDgzoF28N0X
yuqNgSegUCZLurPMfmobcI6AVvs+OdmrfA1nmX4gFA276k+7qKCeRTGyDBdICF5Y
4n3+C7Z/THcNsMdAA36H4SkR92RJNYIymDer6N64cGfiwmtaqxOVlrlAApsUfYKO
8MN9UJRPCCaV1DwlKsnORnHXJwzkOG+RHg9pzR+hdY7IYPDOFe7gj7hZ2IBJEifO
n3MJCWPqyze2hovSpxn+UW9Zt390bpXv17J0cIhbc7vmlE0RYp1OiXiahMM5RHbf
10S1lJfqxUkKNHxxHdSSD+HagzXIkf8WrFZKJ2wLkmPv2PdzOhhV3n+JSxQSLtea
d8qyy5WR/ai7lfZQVB1Eqb1rrYvPHaTzOOnCBFSI3PQiBNK3FmFHYoqaIqPc1Ch6
rzD1JKf+pe9JdADSFFjQkjwPOzinSYYXsRUIOqTE2C+GTtiPmjKYJWQQRJbdD9Xd
dhZJqU42bIO+EwnJfhapMa9rJZbTQ9eghFVM4tO+HYdFIQllNOBXZkN712TiYPri
ApcGXaBndspAEoaLROCmHHIv92/tiZlum+emkdhZUA4t+gyx0koVTDZK0RNWBQQI
rqj0T+1rSzOlSKJZrVN2zP5FZWRK2+JoEhNuzM9d6A2trrOQLwrza9w9v+cbCgKg
VIm3CEEsBDNv8iaaDhCVtjotnVfoLCf3yMPy8qC7ngXFGRI/0HP93/sOMgDJDSpP
5PAMg3vwU5IaWElzCsBcYlOnfL6vYOi8Fn8qyL8Z2YWzk29TXTCYjMlIA+9vMCNf
Ol6pTKfcw8Col7opRRqQQ6sklsFVYXnjxt3NqHVPDS9VWG5gCJHzjZmZBQz/F+zg
YaifubafQ4wHrbeA5GyRooLfb7t2IhS7SPZmXgBXhZXBxPy3QJ/TxnpqAS+F+LOD
Jcps2oTE4oMH2LjIlENxJJxjaSPUzoEmMYqI5ZknfohLf1lF2YWqGRXAsqpm3CL7
yveORbi3dPAe7oQAMNTRwYf7eErtHo72E0GJytMUg3rnraDcqpl44WBLoBbzHy9e
JE2jZ/GGE3OV2Det+8Oab1RS7ZC0VhLeDDXLcIdg8WTg3ZKWQ6mxXlexnWgBEvxe
PxsPdFADmHff4wac8EA8vwzOXLUoBjXF4so0PDEBrRRgAMnaf1sAeZdTuQSrgJsP
0SSEPs4nlFEEUB53kcxzvhWfjL5AEh1TetE6zzoIsMa6tp8pSuUwSilON1OnYoRZ
LCCrxkZ85+WJOFRanVh7vO5lPgvwvTg5Xf2nzzny/Sbf8n6D74VzwUPZiYDLeA2s
FuJmncd7FPkslH0p4ywOk9wXpCOWGm3yKpNswEUYuXYnoFcRUuvuUyARz4fzRybc
Xd1TI85KbM0yD/dodYYbw41xdT2MITRgMugBK3GM4C8rvx9yBD5s+hYLpC7SLLzC
W+x7l/eRrkIlE7P1UiyC1+Zdb7dQuloQRQiPv2OKrX6HSK1dd/Y+qyH0F+IiEVhM
5UV5rRaL30OfetZ41S4Z4g/OP0A/MD5ta3ha5i9gEU0sJGLX/HH94LWT8GWdEQ9D
M0CELfOkRxfzHQYqK258iiTG2DoReAQtqeCVBghsKpjp7V/Fc6CZL1t8gLFO+/iP
vVAsgznnw7nO6FKHyqxE84e+cv/21Qm8If97VZKZbTbNSnUMlFcLCRfbDxCH8a12
Q80Mj8sYuRWHaNZOHut9wPSSTNYJCBhcODX6Vwc1xwajWEAdfkz9D/dG1rIFPs7N
ZvmkIpaS+VIjgANfq0kip10FK7KhE17mHJmDMIp8dDHOMPyP3s369ltpIUNEmd8y
cbaw8wPgkqM7oGfzEEMDMJu+xzbSZTZia+H1fPR0E+tq6O+oKp1rEOAFfj0i7C5g
fem/q7bGsALGV8SuzxdUx4CRaTgmi4Z/+rY6Bt8dFtRJkkbCAsfp+lKpMrD0um5D
JW8xZMU+LMg3Jn0PO3yqe9Vk24cvgzhmTq6dIt5r173hiZuleR8ZV4gpjxZM0uPP
HvgcYx2Ik6qxnwZ2Up8wWbfMRwKFvmFZ1mNUgvy2lyREG8AFvpCArLG/pXNAYISO
zhU2VaEDr1egrtydJYNiC89PlwK4omvTS/OifEURWBwQ1ydePijLfYRsqBDuIKLk
s+LMH9eMEB0UMIYTwtwTo1LLd+a9A0nMbmTsvPCQ3Lwrxwwyvj6AiiBBHNkySxT9
gEGfsuiSBMiugKJx+zI1DBBRw9pTzzqAmDfGk6Eqj+NrIgzljilThoou97vCCMak
ZnYk8Iee3br6SlbKue7n7EiwB7T5j8gR/xyHE/ZIKmbC/FE3gOw1Utm5RIAdVKIO
rHFwuaTEGtJsAgzM+4gAwcdRDvmTdn1JrHBQ2K6KZeii8T6xte4vdbdEtOr0jSyB
0Ej1ExOhCdyZtEiKqcULq3kU4OqPhsjv4kK1zi5Ub2fV9tab3RlU/o2jU0UAvJUg
wgytzJrQLePwoc6G/g7A3oRJqTWvbJfJ3gbSnov6sYUDv9TmLvnsULZZhRSa6nDx
6MF0bQBFz7X0YUFGrZIcvT6MlXvmxGv+PPGUeWRJyyOPVKYCn4Oan5r8RVect1u1
XKqr84fQPougagqDqKZTc9Cp8dCgUqoyItsLdLVp4HmZMbQdbwhafHJbYHQSXELe
2/0zJ+SvPOTFSa3BZcVIpYurKMdQafH2NwMw2eZO8Ir68flqgTeBkQx5dk4Ui8Gp
Fs5J/5MGZSf7XBYF0Fp+1H5bkW2wNHMd9m0ePK/jVE64zqvp744c0TM0kKDV/zdR
U+KsVaDKSrm2KOHhBRebAoVL0+hkUdv4MZrQ316Ch9sjI5OqrtCYf/HJWwYtu5c0
sVfxoir4kNTqwhbs2Kjk9EPCtqQ6H0bNNjkIEdjc72FBS270qKOSC1uTNN+h/GHI
AomeGrP2YZpMBu3wTODNhBRIhKTmD/duJsK+AetPAq+XvDaTlO+SZHGImUvxEix5
ETCT3ZWM8X6zf7smb63DvTtrP7hdRsuaCtla5GkLguEOpjB3lkJbAiFA1fqil0qU
WFzpjQSRwbyUC9zSQ99pWVcuNr4ON00dQllpb69rlONTqevdsLjty6Y1jRBsWa/Q
fDYulBacLMCLDP3fDvspDu6iZ39sUkC/qPFpWV0Oskdc38OvfdQIIGTD36VB9015
nrLhLsKHW3EYxtTtFlyLFpb9NKE+lSfah4YWa7zu8c538QVhwe4qoKYv1aiAxPm0
++ADz2pDwdMTYxrLrxZGfRsUN6jsL+Xag7tbSnZAmfcO4dMndOh3PJQw2isIGwX9
kIEbN+Dwkb6YnwU6CIHYkTBu3SxL1PuvPAxQtrJnovSqHreXp8BDTUsMIIcHsEVt
PO5WF0XpJvw9kZSs5FPAg5qaE8a2+dwnj3Qf7NSV5y4bfqs14cHjlW3rkRIUXUtv
NCAnQFab6NVWg79DQlYeXzoRTQuVIcj0opoeQNZjGekCLXcdhlWEctAosTFxrvkX
ec2n+Swj4+VrXJdWhl9Bzc+lYh1shMjFoV3JccprlhOjs6YDEisDUAyS97yZVhp2
asrNHiDxFjXTCFQZ3a8On+6NvAoMwlXE57UuaabcZJdBa7T9cqyaUkf+VyNtKCcT
5I0MZ9mkkI9MUtIQn3fGdMUoBsOmUp7PUtNxSPtiFcW/+wnYAcnf8Sg0SS+5Xq2E
zLFf83zlZzMCXZmITNZrM3gnb1fiPJAB9hBsZ5HTTDGVZ3lWgTHVSGn2xuTR8Edf
48U2rkQpx8NDgKoTTZljWPEB1Hu7vKsz8RyOz6/SLzTjCsAE2YoliPQTMlowKz3L
BxBjUMyaiXeC7mON9Yt1FZS1B1kWQN+AfT7xn90vFlcjrdslEDuavO5v4knaojNR
IQMF1depGcH5pAhtMEefcEvMJCErknHIrKa7YkxY25VGeTdM/ptAIRSpBfnF8aRe
j97C5WdNvZe26Xs1drzPovbTzm94YfvYdZ9UYOtbrWzLudPfQEVDRJSsr7B+jQyM
5DgJShBTlRjlyL1k2W+QVGcU1Trfg//fYA9ICvyh53lROy9k5fAq/oYv0Bu/3/ji
DlHiZEi/Mq4km/5fCBYFp2rqXyqKWtTmp1fCYra2z5tneqPJJf12HcahQZPrttp5
kPsGy97zquTVZ/cT/7aRnMimA7LcOBZ5ReFv6P2sqGqlNZmC7scFnoJO+mv6mCUU
cFASsplaKuUSei7dR8tuRclHz3GVReryVGbvMKfz3PtUbshjaZ60YHNaU7mSRAhl
eDhs6/pWOy5qKcMcMaEc5PUX4kgT0lGqCtYOoK4UqYPd9Hwa+j5wq2pIzCe8LdXt
yVPuB+sotO4tXK+nV6+qt6SDns90IpzXLpEGlRzAiHYLvROA3P9ma+8TN60o0L3+
pS6Xn5tp5DQukDJdAvbPygbW79jbrycQtqG27JMA3zCMffWPhxhpwL0Yx5QYTgFc
9w0LCWn6Tnj+bzmsDsEIP8Tr9/EHzjpBCBYKPpfOgVYY6uLTiAbXpVMbq8VX/Pv3
z8Y/++drfUBD9bUw1kJbg2Qb2LChCQqXXpnQm3k7lDVRyIu6inHv032Aj4YXN0pr
lTUW0qWwepv32923I5qMYMXnNN8tznzO/Dq94dVUUFfsCVGHiZQTcZQtwABfjdmz
yMqkiUbiCtILEuQ/mWp2XKov5gSVk+d5zyEZ9kmh6/UdYmC4SnlCVUIsrhfk8NQU
JpUY5im08+C2bSaOOnEHmq9qb7XFF+CszGg8mF5tzVBYd9yQ0ZHbk5VFikEZQotG
qFL/4YFotpyAPYBBaARw+Uv7E/k8lo8uRTwNyzxSTogLnQz+sdD34WQETbTPme1b
B7L994j5SWSQ2z9KS9V50zpbKDl/jaTYdcni1Ouf/Ntfwu4y/RKnxbG12gpijEL3
ZsX3y0Yg9ZJPUB9j4Lwz91oykOxmKCZlzUXX+aArILTy+tpshFiwtNO+19yGGKZW
N7jLd8vUOURgaSILSEbwSTU8XRDFC72DoFQwM8MmuPs0CpdqvhDijP9779gBNBll
7kDtk6fi8iklYtdvCUEuQFNf3VOmfshoV9mvFFjzOehngj7E9bECkALeu3JQWDmi
pH+VwslNnzhKQo5lYoO9k+jfITUS6rLvnznLhV+zkZXQQEfDACkD0p6Vl28QQxzn
khB8I7iR2hvxo2/iwQeqlCoxkVXF9REV7X6E3NdCAJbwZud+GhuVFZm10JO+j8CX
KGXsUsV2h/PkON4TmxnXckdRuepaWe/Dx59l8HG/Rl4=
`protect END_PROTECTED
