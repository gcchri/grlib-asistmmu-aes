`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJMtbtOfgy3Q6qkapXdbw11UpU/A9cbpb6TihiOThTnMVoqPNUnpSZFHwZJFPICl
CUSFsvgOmvmpE7WaDP9w53Yn94nvDL+rPTTI5f3UlQUdurisOanWSRb6iQdfkSwF
ZMS1AVF6NlDpEK/Xx1sb3zveq46+PnDTqo1zDYe7e8Obfntumxb1cUbs80HM8m7F
HRNFdwb1n5S3xK9w66KnmVFsOJNnaq4m4byBHqTkYu8XyUH/0q4o9jGhZUTVcg07
iJvninrJoDOmJcmUrDcinCdt0mdhW14l+1PcbW06Qfkkc7LMGXnu+VuejcqgJTQN
VA30XCGO/7MXlV8Qs9X83tyPTuHGHayPlmetgkFZj/lKuKI7Fcr9UPTEelHQn7NQ
FQAT9bcJAXeBloQIGmTjlB9rSD5Zm0ugHOOO5bAmbNYh/xe+yEc70FqEbe4k3d2h
+qCZmtwwAxzJf+N3/MmQKq+iRjwCoYxGUEIlq6AczU+dwDRE7fJqhTQAa1Vgt7A1
LYvJScZDPJuI2TXacKr0lg==
`protect END_PROTECTED
