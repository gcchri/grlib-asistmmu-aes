`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DhxU8Zd/Tgsfsiifj8qv6aN6pn5F8n7JIBT8VtdIZTrNhZxsl5gSSHcm0hp8YaQX
CtW9S+quNbFU574zBw3hEGo+3kxmAupgvNhT3zpXq/oVc6deoGl4cptrgfrOoO4m
poC3JBpo+WntbTwCFudemD3BV3FppAh7wtoInN6AImGM8Uke0J5C+9bXrW+pEPsy
DoxYzVJWwwIJU/DXCV51237Baqmc0X6CKdxKE7A9ew9FKslNcsvRPriC/3hsPoFw
a+po/eLnfH40FASeTplBvVem7AOQN9Fv18NXQaRTvm2ogqakBVGysvdG6sNOFmRf
9Gn9Lu1Hgy3wuT9IS99bEs0uffJ6bp9hbgFvTK3eSqlVBf+L5avJh9u7ssRldoKj
mXFm2L/Jo4C8KVpgkhXxEpyIInjl9UhKa/rNlvWGgzJSKTnpmdKY2z/10EVvT/Vk
/sdjXsgYtuQEnV7YhavqrFybPcK9lDRSY2IJnRLJputoJHWTd0Tz0d9y2xpI2B5y
HcqlJurMHj6Te9F9WH/qN7VHh8a1XIs74CPa1EbSH32M0NsqVY/IY42eCHzXF/Ab
j6JkkBp2rxp8yqmGVr4qe+I0R4fq6hH+5MhBFxkEEmD23vehqY3YEWPBqn1eYIDG
SjhGQmlU5D4AGgEgufblpZkgfptarc4vm/azQVWGKE/4kKOzbtXUOXIRN3PkaIFt
jq00WugK9hvlVeuXfglOixJBAwWpK2kEgylwcMfQkH4E/Hn0jlz3oHrp9M205SdM
BExvIz1f8Qg1RWjuBPLX8dye2Kvb8qV6EZe2uxn6voj2fIvSfUz74Q5Zlt/6fVxf
Xo2S6UlXGd/vqBs9N4CgO/dBbD2VqOV0+7sUTMib3rKqC4kxJpEhG2XnHwVerCtZ
zNFdGjjIKCnuJFpi4Z3jprJ32Wlq4bEXCj5XOMvRSf/oc2dXu6+VCt8SvqCmWUse
FtumYci8vd8KdfWGrEIA2+XGAdvou+W/aEmiHgsGGaGnxqb+G+Ru8QS8kB8WeKH7
AX5399uMUfnjFuMruwCrad6m9E7xcHU/PyW2yRrVKY0Io3u/edRsbXQhwyoKmec2
a9pqcLWjLVktKPaNf0M7z7JohM0LY8O0fiK28gPUy0BFgdp2RP2xPYGnLZLgKT6l
UemxcsVlYqWC84QoNnzXsI8CnixEyMwcDeIpCvMC0m/jBX+eW51CFseVVErv725U
fS/U7K9IRxrbAL3jpvNWF8CY7Rg1uhW4CV7IgSbE6EYCgQtMIrndwHaf3XALpgoV
x7uXm95z2f2CLQm5nEC+fguhkmNbV2/JpENVAOb0DYDMDOZQ5QswV5YAcLF3CZtc
2xjmUvkxGcb2/VVjomb4g1XdJs7fW+Fe0T4NV9Q4WX79X4KbFgDvfEC5bZHRQLoZ
9xV3HB5t4oD2xceQQd54Hdbv1IAe3I6QWZmJtCEi9rHfwjO2M8kLMj+JpAH/C6qk
Xj7oJ1HGrwLXKZkIKkZqjKAO1cCMSL78xU8WOeVTXWit8xdlstNBDVIoRlGDCiU2
ZRXKYV9JCyhQCHU600aIiIkoJtqPJ8/zwf3UP0VkR4Bxe/6+DXbTZtg19Oe/SQTO
+yNHIDtorvi+nKVHpFechHqcsEyhipei3qLVfazVDub8kHj4Dt+XFKqjhf56tJxA
VSbdzMmHqT4Asc8NBRuQo77RdAIfcIjQyIzJvEw+2zBMyyRSWyV3mc7vp26GL7Je
3gKL1Up4AN7QnmJkg/Fh41ZI+9yQGB1GjRh3E4Zh687E+AmfC39t6R+CW5U89mUp
vZOlv8XiSK2Ily9Iel/TukZSFYgIuv2uVAan+vlkk3LKQ+zmDcr4EDXdJ9FphUo4
`protect END_PROTECTED
