`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQHniQwc/wTgzbN0RLhS1lXRqQaSME4PW+ltTMEO7KwRATXD9AWpmc2CKT1sSqjj
Pd+chUIb1EZcHa8GIr8iywRsvvWjlKfsjdgIc6BP+ZGFhnW3HGafVJFa/b1Md9cT
gpttKZfqAWBe4/xFJYCx5wSwi+V7g5MRY98xfhmbwusF6PuwDPxq7f9bU+Bo55um
1XL1sTVTJ5gH8P6YuScQHfZdiwD3q1CLcXwyjs6J0Kn+uYFioAAiT2KXf83vcaSY
46rca3ukUv4XTszH3RklCRNCQolWHQHJtex54WS+VvKCTmeBZSrWX0o4oDSvTPmm
7sqrepCHzFAcaUVQB1ZI/HuBh1w3p70nDhb0cqcWiXIZnRMF5A3SeEsUMSBE2vE6
FNpOGQlOg91BFGIoxU077wp6YxJthLa2L23856bLcGeRhy13EdjrKJnv15XeN8FF
eHAaqu571kuECTPs1Cw2FuevMvbIixub3WxgNA5/0S0=
`protect END_PROTECTED
