`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r296zvJkMW/bzIBYdnGZkLqS/qCAl2/TvdUSwdMIp4AtuvpZCh1P5xoUzyT7mEaY
Kp4TKKXTx+gSy/2F8vARiXMJ/z0Fe8aotztckTn3DowCsg656u/SwhxoZ8MVNE4Y
mZG52lkP+CttbgyYoEdMfGWZerSKK08+IMbxwP23HWYOxxKXeN07U96IFDyxXU5n
89H7PoW5V/cnRnZBZv25XjQL7JQqppFXd1whYMOUfrwIBeUvG4Yz5yGTb+mKX+n6
WklUhi8bo7AbOkY+7cRJ3fuvIDHOm9jskYxr3fBd3Iw/U/tzAfs2XxEEURphNicn
E00nkNoCmFOq6NXjxoH5bw==
`protect END_PROTECTED
