`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vYDaJRpYWovVw+NsCNoWG4WCoh+AxdveMwYyZFkKJ0dH7CdO6MsimgdYNfGIosI
+dB6XjysZ9BM65JBEnDIWSvdh/DHEQb9xx7zS8ouk8lDSWx04IhLaCgjwRfaikr1
7dReDHXN8c9rF0GCKEtQaA8gPDPOjykRAwZENjCjhz2hBOvp6w7jdwlIa1yr6y03
CHdbbz1WZOltl0ix/EbYTtkFkFYTB8NZBs18FwvXH10hVLxhIB0W4D27n5elBDkY
x11FyvQhdg9RHoImDmSs0WDo3vTTvYhO5wcoYP8CBO/RajQaZEEIHYO3yRbBtR9V
Guf4IzIk1dLLKTVfWMaUo41pXm7XCXC+grINHkjWds7NankHnJoS785oViqB/hLW
3myLgTLnVKpPRmupou/Nf0G19YJabZE0vLcJxZrxvrO/nmSzywnDU1YBEwy4DRXe
tXAMyDyfpuKnDyzXccdETK5VR3GigboAGY9RNaHMvEzk0bIWSQgyyhyez9sjKnEF
1Z6ULai2CVGfUEOWchzIYjRxt+ws08c9MiPCUgcDGNBblqJZTrnB4YNAv0Of8Mpf
DL+QbnQTIix26Gl2VpmUhMi2ievFzi6osMTBSohWwcwb95dnRTFlBcDyT2wWdraM
/rLENXMnKDgWVRgAnczgN5qxCJR7U6xhBtEeTqtcmDl3/hf7Sn+r7ljA7X42Y/iB
vZfUrRFRcK7ibm43pPG5+O5OKlHazUNm7YOi3C4FuZDuZ7YRwjbWQtatKeGB49C8
KIQ9mTR1NBgc/43xlvKCPQ==
`protect END_PROTECTED
