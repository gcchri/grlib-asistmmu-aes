`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U3IOYSypUzEjLnWevOcpnamrAKRaY5sM7AevK79wcDd/xlTT8KquK8HKKsKx4D5F
sKlRSvJNZa4FftLo0xO2xbxLiYeMBOpLyG9/tDt/5EyVgbYqtkLjbX0EcgNv8mHK
1Q7/J2gKrIqOweOC1H9wih5Sc1U9vxn1R+SMI/o2eAwHuN9PkVmGwkEB6ZeKoEGR
qkjajzCP+djhnKK3s4JgiPPbZNnV6dgFReM231MtQwZERX9Bo4s0A99QAl0WXkOY
lm/01tCfZOde3iww2zJBM43V5pcX2aikiwFWYXnOiKLbNy6yucuoPEbXEneoUKxr
PUqMZiL95hYi0MQrwwhGJfYZubNiS7qRHZ1lVCX///aPEZs97w30KOqyeWGGlj33
bWgEv85BagBpzGfWGYLCym4jeKn7iRdlFE+tbYF8n9lkr9YDxg8zUXrXrEAPwokK
ek0PKSp0QHLpluVt5Yql0TzwWymBpxhBDvN6+DTZXLkK8bIjMtIMpBwKONAguATZ
UTOMuFMEOl+pBpjj2Hu0Pqp8VszXl6v9pcs98IXKxQ1ub7RYw5iUDqjtkooUi3S5
IGgkrME0GpAAUNd1AoFYZfYkJdn3zb9WzfE7NqKssHJdsdqXwcc3Fue37hEKYtK1
coFv3Ax89PF2OMd50PE4SF8hvOhMqhXxvBDJDDcxm+d1BCJxCLbjnsWUv5hN/z7r
aIQ585PGpdyLCDHdP1xJ/MTVhHD2ltZD7JH2QstgJVyHGWon4ZCBj/R6eXL5K0Ex
f6MJt9OhMQFNt5Oea8LdFFmn4HoWOQvVCQrfQ27/PzCMntxLLD1aSO5LVQVzKGyp
Y4xDzcPZ6wQEh6jun+McgKnZziiw62uGp9emq7ilVAGa9ORpIYfI/lyH2WODv1L0
ES/V5ZpjHC65OQc1NqeWl/sJoLfKk8OLo1ymh8cWLJzdUB8WtCcucP80I4VqPY9+
kbCvuSZTj2URHAh26d1pdiORgfiMNw1nLTYwTqulOsrOrT/Xuc9wufPPTS/YMfw1
C0kxQDWzCGaZxa4dsiLmE+DW6U5zFOijXbhmOQHNWVlApDBH63s9r5DR/ENPnlEl
s1+kLrdl2r6/Xwg811oSefWHWo4cc9MaALD7KgqCqHn7LWt7LHpZKB7IcXxT4QRa
p7iARJImwiYHr1ZJpdV764L+X3qclyzvGlANfcaxzPkkh4ENkjOpwMj5Pf/7dcxy
whYZql9Y0qb6u4osmbH6QBmal7j4OgDYapoiENTSkHZPa+5Em/WKdgBcFkEAzEGx
n8J4cJrXyvvQqwAbA2EvOc2nsipTwIod5y8Ewzv6OLlDj7/4v3/3JqerNnIO1Ovi
ae55FbTM1pHQYV4VgpH7/tkNzz7g7sG20/WDe2EQUDPfyMvu3+8Dhl783uWFzPgV
VhdgdA9Un+//znNwvlwmjUz2zybe0ml/NGZTqIW7AMAxx3LUm2e6QOs8N/bfYVJX
7ZqB96cjV0C/cY+rgaa/evGZyTqSaCQ6avAKrgXegJdOSlaosLs+hGTe/l7EefnL
CKipWeAODS9ZUCdF9it1B86xwKeMdSrNHX9nRCQNchbRTRtIAFnvbc/7RrBeWKgF
C2tnD2Kwg8R7akK/50KvOvqBmYKs8obh19B3Jnr3xYdbZHTO/yJeW5DRooo8ujtY
C20jpxAwxYOz6SmSz0ZB4tJiMiFndHb7KlfnLqnby1dULCIdqIbrEv9tkiY2hpLi
un6duYyrwj9UGN/j4rMlrQGF836MWerJLeFUMW7RY4CM0XTqQyHH8H8iVQAfn4tW
fTGwyYOhkmUbla8UDcZt2xbRFGW/yrF27h0k2SYxFyYpYZqiZin47zTD86pZaNjT
mAkbs3NFa3xfsPRsJEC3+TS216Jnc9UODLdOq0K3Rb+MbwehPEOwMdf6wk7O93y/
LVjxF8qQQN5qGFO9ui8ZPEqgxitrQMuN3uG1g/UL2CNpPx0XIOqxizzpsSLcmu9c
IXDcnacvoTEtXVe84+GDuOVbHqU8qoWvWxKS10Eszn0SFjhKVcm6aZ9EBsW1ocOu
bfJtSajAFm9BUjwGE7xjr2mont9tbtX+wnP4jGzy1QvvOc7e5n708mG5PM9hAcDO
MVBhQlUrpZOP6fT6YfErz8VKl7iDZ/AXLRGcJ5DG/bh8lTMzMnpXeWnN1ptj1FhZ
6uP55JvGKIXzUKQjSdkkf8lZrId1PemHDuKsGm+3z+uuPhNip0c3zclc54hyq3RP
JGvN615B9YJhfOBYOQ5lnIUEkClk/0Qti+kuJSF7giCYksvJM1bPPuqThV9lFtn8
q79J5opib8ykX9GxpV3gf5eW/kK1gJSa/aCrBkO0KiNTYowHmDK5NpAkePDIXuAJ
cd4DYT7VZMCgOAFRdOXaoDC4FoYYKbJGmei3Mpa/52ZiJ7+1CcZ7clugM76Czese
XuSnbQOmDT/o2WbvR/XSi3I1Pv7PCjwLNp0mt9MjMbs+SSkGeJdIi2XBhhhbAz+Z
PTWMAU7+6K6tUudoee/gOadnb2VMooxEdN82h7k4mXGasN819F9T3jfsl11dNqiC
KfaHAyEBTBjU6ktAoXrKeZLKAdWvK0gnUkBldUfgkmKWhfO+9IXw8Zx/5UXXjVxJ
topWbcPma/+kFN+OI5zCFiKSqqR43MUNpxIwzm91qcnhi69OSpd8zadJWLJ1D7Kc
CQMfp/sksiZpO57dHZ/ut2dJEHZS8PsSlIRC+fTxmFHwUicvSomszK0KPAy4vXWY
M2tu1t7PhUUMS0sMMZqlt1/4OWzFBjrznZB+iHsQyMIpGj+Y4ja4BUktibNGn6/7
Zzm+DZ45TPcdTbn1VwtPGgvtZXWcsVICq7HO1ye+pDNM9K+A+UHaKMyuWWN97Do9
pNGm/s1M07hpBkYLRdQch8Um/OGkN1xo3gFZKPeS2R5/cfKF+qgLhAAL/RX7T87B
9E8CvcLibnPRxK+2VouMpOsa+mGZ9KfLfllg3gYw/WRYKwfG2h8Wu+cMMUwnIjMc
9o89JNnRIqNvmEKkIEU2S9TlzSIYZgITMeTNgf0yBr43L0vAFmOyDhF8M5h3naUH
IK2jcZif1RxmxM3i3k5LRu6yy8AskSe/s882BuaKbIagKmvEXMTcISyghR3SP5Zk
7SBzKY/Vx9wnNPA7G9SmpaeHYVVpu9r42sEqoDKV5BcOhY5lHfeXffTPgPJty9H/
ov/ov/H2HUu5q6QKvTB3gs4Qgjcu2dJ/JHob2L+hfuvqGWKCjZBP/SUOcL6TJebp
6MjWeaSELp+Ym8Lf+6uUDNQnd1kIytLdhXa5odBMkkh+5+5cYTFx04KBxF6e+o1d
MEkLT36pBH8d0nWdVo0JwKCpNW+nCAt4rRIoovl2QB/aL5uVhDBwwT9bQGRZNrO/
aKHmYUIQqAPL6rWkG8KzB4M8mgHg3bKkvOx1jMRgMuw9PmztPpqiUBSKFc/V7idk
df5YaW5gsI6e1mOL6ptf3a0j2W9VWLG4cXlVI66U+VU6+rWqn0KzcOV9PAnC2qkO
Ux34ka1Gb5o+z13GD3mrzYGmE8TmVMbz0mmCpo7GCBGRXkFXjiY5zeRf4ot3Dk9a
kaW0o4BbccYb31gcuB773EX7hYWwd2u20CimOY3ePd/ac60fq0YufYLK81pnLKdW
QbjfSZkrNCyPIvNqAOQ6HQlA8DG/9gw3LZikyMHNCiyvMGaWcmRLC8oWejqnEQTI
Bvb6ys6lpjZB1WwPz86CWJgnvkD1U2X306Fh2EcCPem92/tKSBoIf4Ash10tOQIg
CqsFfixdlSa0ipK09F7bvWhAYvDjYOfTyYyHR+zhMg7QeIyDPz0T7lhrtX6fv1AN
oDpPCOMwXR9OHSoTTHbaMZ0gQQPh3ORH3ZM7LRVPnAFkBYG6EC8uPa4i5MTxEUlg
5dQFjHK1WzC75zRSJ+k3HNJGaXIyb1NHnKSbQZHNYIqaDLSZrnyU5CtDZkIyKy8p
dEUTa2rd5eSNcB+FEEVGXm7akzpnC0PGhLhTWJvTRRaaHGc9T8ZQAG7UFCN/5DVj
tP7AzdpOW1pb34ij9KXV1euVCiRBVBCmoDrjn3OUAuxYN7SPOZWaWW3940jyXzpM
kQepIxrlGxyYEedBk0DALnH3ZeE8ZePtd1yb7LK8+EqbmMx+9jl81fXLGcZukgVI
N1wGHhtjTZ79r4h6MrGIIYcKk6+CoKpLD9PosYkrEBXao5eVdN4xnGSNxJjT/u1C
xqaWbgJonqI/7hIbZ3p+ozioUHRp+AfZ2GOTBZB205KuNxlD6eiv9lJ2GZd1s1cr
E4O4N2lslD3gD1u7JykAa7v3VWvZiZqBeMv2bczIMnAxT2WcqIZz9Fl+4Mp6Okht
DM0MVU9oLoBUZM0gMCNJ25aVu14dHsxth3O4LZmAVfNAaTEATzQoJxsCjggBfoCI
`protect END_PROTECTED
