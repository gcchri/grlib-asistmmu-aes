`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFSHu2Jb+Dvu9GGc5LFA/7iav/bcxZzJUWEqrwmtniWni7xafFB4CiJFhL/+rU51
4GM4CekjgT1LEJNNKECOcb/7pZMT3sAEkNTkKTaT3UhvWmV/qJIhRYqyXoZZa+Z5
GXht471OVsD7zst1T8nlxs2aV8nmswRs/eAhdfaaLkqpB+Hx3JjuuyIU35CAUr7V
ExZ7Kfs1lefVtZ4gGPAxNmkxGR3Wp26Wc+42TNAKHBgsKnIq/w0PMU8BCBAiwy4+
RSznpAv8CBiTXii+YA+x2g==
`protect END_PROTECTED
