`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eU8QpP9zvvGyH90cdXSMqzrbY+nu3OnZKFiey/BWIodOTvrIrvTY7k6+C3WfPOCp
UJtFcdHaEMn6QK5xg39SzqzxLe6EtTuqeEfFJFfdxAWFqTvk3ZJv08+p1vE8WG1g
/HpAd+Cwjvx3RmZUOr7lq5xhCjKksNgPp1MJkndPuziKY9QL2rE6dXR02sz4XFae
E7vJuYfEcGoxFZmyFNeDZCxgEe8ZAWFWl0Or3JlIwM9xXyIbYlWGCTcVPbmhwfmP
6on9Op0KszI70P35fOPVsdQ7qy8g72RGTBa2xF8aa8k6BsOoAb/RRDyZ8IUcMRzF
KpfShOUMQJw3xrwNIHgXhqzg8/uUsjq8+wPdo9HQFXeMBGDbjr7nqHUD6nn3ReTx
v4DzFSeAW4e+S9ESefmeAGm6dKKMTnxl/LtSaQw5UbFh57gyXZJ1Sp0kHAeyA0bb
2cfwM+YRIiBKFtBgakcEpc6oOFQHFcWlZuBBxXz4bIC3Qs0Vu+hdC/CSM1j5Nmnr
T5jp3mNqIsW8zkQJq//vumwWSuNuEGf84eAy5Y5KUhvOPCekzOFAqGV2gF1beFtL
FbiVpnny9G5LFUN/7vyMSLsYyJYI4xc0Tunui5sIqgAMNGlAwaqtSHC5ezFtQiR0
cyTvKZUiWifeO2e7HKGkr9ApNUOKZZayAcPB31l0s9VA/yeuUu6FmenZjPwZcJjT
i22QRNV7pDzzbF7a2or5y8nNzFTNmG+7KCedfzVVURPCc2ZuffnaBbiHYGHhqZL/
UV8IbFDxWrAmoauUt5eDliOP7ZsLdPUg0sVF3JO579ZS+4KclduGMcVO+rxNd3kJ
If+Zg0Zc9rycl5yJ9wwDhQlr29efcuLeZdXD333ttRlOrjgejKQT4PxQbJr+m0H8
leNlktkUQNOhsI74oUqv7w==
`protect END_PROTECTED
