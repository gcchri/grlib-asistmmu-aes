`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTl/Q3/V8Y7sM4BxDEj2u/KRYcHA9Nn/+oOz6fGWW7gpJ/8rztQ1qHlpsEPm6EC8
10T7a6MYoorUGkYuUF3pS0Ncwh4rMNCBg85rHhh5/CdrA9ak9cy7OUANu17cVahz
Wks4RUWP4hcAKdv3NgFR4zBXcJNAI6Yl6i7yhqh1N9/YTRNZBxXqNCAchY80o/Yl
iUb3twOR40x01YEZibESrSdToSUwiqQLIIQ5AxNFay3SAC6iF1/jK8909IqfzNsO
YKIO+WEvf90Wv3REzEfsjgyCn24Gh9+VMx0p6gAsf7GD/uv4TpN4BwLClQ4NBGB1
NLJmEthyQ9vqvhGWYTCxL0kLPMzXKmtdWgeS6I55/+7GzGlnMZ9FMdtVRtmggvGb
1Ddb/ArIjhIRkLg7jXsPJFg6VsKiQFPLT2OvdQL20LJolJ3mf9O02q3/p8KMwwot
t2FqaS6XYUesT8LFajFx7FYXqQUnVcpem1C9+G/qrKuA27GB+TnIN/0+o/NBX7xN
FTtCm0KLJFfZACVDeIg0HlOhcu2YE8AWcXxq2Eaa+76mmd4AdYkaVoqoplblkveJ
KEiSceajhDs7bWKZxTJ537iypEq3F0zaZT8FX+l/gfach7yUgAYxKz9yai1GHWfb
Yn4bCBaAI2jwQRTsPE/SBAHgIr0FLyH3wm5MlG9p6aZaR763kmMeRCAMlqFmUc2N
ulSWFaFDVHMNrek0hXz6MjsFZLrAqFshtdco1NcJQM4hE842MJXzE+DKTMzIXdRo
dtxluJBNQd5I/RDCJ+lgxTjzppASGpjInKs1unpL2aRFYcBuSXq/WYxfRPCtP4/0
pcREjZ8nN7aUef8Ad39S2Q==
`protect END_PROTECTED
