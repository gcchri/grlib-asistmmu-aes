`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkqCEaiMjfwfSdQx4+vRe1WmI7wM94+YTfMMdABFDWPYTL51cAJX0/ui7cHFe8lH
9bM+j9X57niObbm8Sh59ctCp5co2ZAGiAiwiY09+ebvTkW6Y9w+/SAg4o2gUfQqe
+VZ34ie93+wRms9wNo+D90Cl26d1Rj48X0ivabRS4EllcmwBNHjXWRBDEkjs3w2v
GrUKUGMQVq59Fi87MPfmET0gibSoGMVft6Zudoc5E/+b0vPSNlH4SJ/dOx3KfN05
8tFFKn3kbBhbH6T+OpFmEWub9uByWYQOT6HzKgm+aaT6dE4hZrt2ALbNi+dGD1YT
ggG6ZUC2Ny7rIK8NZuHdsw==
`protect END_PROTECTED
