`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWRWP3eL3XHWNAPSXdu9lEf2BFhaPFoyLBkDODlTYu+RteO09V1auiNuOlpXVLie
YJ8ePDLOWEXu0T1ak2LY3ooZN6705Lsqu28A/mzftD8UoGqm1A/91109IGVXLKB3
HyozSX5Uzfb4sak1KfHZAMOiv6UEk8SdLG67hZwOqXpDMZklCCxyrgQBCDAlhPV/
3rw9BZxdnucwOj+znprhUZ09X8rffvJpLoRuYAED1HAFaxMvaTErqfJrTBhH0CzW
IpqIAzhAXukDEoUk/yTABqSmSeMADzm0obODAX7CL+CRD47N8sul0xNm4B90ShMN
58icgtGPEe/M4hzJCB+YZA==
`protect END_PROTECTED
