`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FLvBG8PTWsG8mNccrMVJm6zSDxBuF3Uey56ge0bMGatSIZhHQHUH7l46gy1a6OQj
iu1xv4zGkieglvorHjpD419dR9hL8s8m1iactZofrZ3v6L/ywuWrZAk9DI/wI9/y
NzN1kwTW45CIWpcL1AFYygd8yjNVQ6RPsVWkc1dsl/L+K3tpYxpSPGaz4KECfz6u
5Nb2krywrgJI+fu5u2k4Cpmc5pLv2Oe3Xl4TY0QR9lWmW+aL/cyq3KnmICy/xXzQ
u6P4t7E/t7qW5slamhHnMw==
`protect END_PROTECTED
