`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FFh/pvSOKFXOcd17F2IU2hg9IhwEvU4cdMkkbMK3fqqZjl5wAd5ysSafSClBvL1E
BOjjVHAO/U3d9uHY8+uIRtDcsKgms6JwGR6R71qcZgA3QacxO5pTyTvZs1KgRfz+
QFXjSCYSe9xo+FKfsuLpQukSVQiGc0vRa0aDxynrHwDJQxgVtjudldGLxaxZXDS7
grf5ytucZFulQhKeRvMkqs29SerdU5DjeXUKSGCZmAMsNpc/hFDH1kaXGyhoL4V0
7hKwLowrI5tGrkrh9oM0vHgp0huNT517nX37mey8PuyqoRuRRN45l3AP2AhDcq3A
yLDXslLIQYyisAUQgIESEW3gwM/ysahzKrGewTOcrByEWK6UvqeuSJ/A2GupPOxJ
OKDUc0nQq1fXxxfmI3z71Pc4qcyKYTJNcq7SgQizoCYKlUmdsGAPT4xe084iaBNo
17pnXVnEhU+6PFWrBw1oicHH8UIjbQs4p8GgXxx1u/7Q4ab7pG1TkuggVFhWkyQR
/iSrLRjeoAp2yoHO0D4aVekMwFlbsn5Zo77eJrlVcxh/kOD3hrtJffPBl58D5HL/
/sr2SnctbRcd84qXNQewSiMaAbyr0HCeLBicMQprQhLNUh0iix/wlzm4RI+6eCgE
/CoH2sp4dca4Dh4ijf2P3LV3BY87RilOJIBHAmMA0mVFQte+U5YXr5BkA0SoBuJc
peflc37TvPEOPj8kLYPtPp8n7BDzlbCtGhFZPdrkMQF7i7z4AttlDxRXV7GgXKqk
`protect END_PROTECTED
