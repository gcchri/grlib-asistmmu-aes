`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uwcyiBm8lS2RfU4t8o/OeciAOw3wCMbbq/lLWM0irlciQDlXMRpdQcnQH4DIvSP
QAqd4EpaDwRNoUOUa6dCs79dnnES+zW2Jo258aThOePAjkYy4Ajf+CZGHBjMKpg1
IuWncN0BPl5x4qId5AOcqhCbYSmSFPu4+ZH+K0MkWtMugMGu4+U607t/KVKgdSb4
GkYJ8fC23HU9rolVngVwTpAS/BeEwmtrUZiKODt2hE5FYQNDgKwWSbIJr5QALBaU
HH+JTcANRVcmARvbIRot6zi+h6wNc/y7271x6NsmPhnxValRJ34WOphDzwsQ3sol
59USCVTRoc0J5rpD9/MjZvCQoP8BGrEM+cwfDDVmzkwiaDgDqDVcy1FsPGcumUfP
kGCrDaig5mU94EvjE39HCPrTjYJpqFdspfqyRh0RnD6bqamQ2Xd55tPVPk57wjq+
mI7h7hzww1mgoHKsm5StZY4cs5dfMSCishLIr9nuvSlycJbW7UitOjNhePogoLIC
q59K7zkClgURXNlWrt3s5jA4Mpk6DOALT5kLqgUgaSssvJUqzYbAQPMB6H5+3S3N
RrbGBA00sCrzobBRFuqqT2fvxzIDnCFgMGZ+pZi5ULycXCnJALqiaHCgJiGiU54r
/Zn3U/loe95qZiBE0wuAIeZWzzrhPvPDsQh2dGkRQTb2U0j4KkdUgMGZMSfA/b+X
nt+ijldXsnvHRxIv+JRKhrpazhAVDWC8PHH+ev6aGABZHKn/dZbeUoopJog1WYkB
lnluwbGg+O2zYlG4+v3rSw==
`protect END_PROTECTED
