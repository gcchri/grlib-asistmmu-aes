`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yllM/xqpzCfenzT/29zlO/fK9HoZlAvPoyXP8S0aJ23j1qkDKc4+k62AFNkr4Chc
byguyRLhE9LT7nasZNNJcSrJDylPEm0xH9j2dg/Q1sMocSM+z+U73kzLhb3qtRrB
h7OTbsgbhqzKUJZawH+TwSN9t03ceOOtzqrgVzPKSsTIumc4H7pLVBxWN7WID8fa
TQIzG3Z9W/RgowOf3gicc/bxpjMMnXV02q/t+ZQcvvx5ORW7SX0GPpR+WfIztW/6
5L0ChDV3EHdrJ21eAPp/s6gedgmYkcIEFSGfBIdQlA1WE0W2Y1Y+er2iFzJfHFpI
/t7cT0FnCSa90wrwDs6hMJHNZvW/A/k74taWLm8RfUtDtURLytY2KLhvgpXbeD26
ro7kGoEPo+7gbBqxPhttCH6gNlvTUx1L0PEegCO+FrHBUabbJhYfJuXkhixXdBMU
8fevNHZfg5I+otG19v/yxWz34vJgyY0/2jylpr11TZl0jBgv8Ht5w2MgbrG+g5jw
`protect END_PROTECTED
