`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rp0UCdjF/c5WIxBUsCErr7gODb9OTpnzbryQ6nj/h3He8bP3acjN2uDsoAWa+yJM
epjzCwOlIEEHnM6My7SE+QlZthgZNfcEt2u0EsOTBvoX4ltEw8Yi8e7ck+15EH9/
a2ZWlRYuqkCS/bjuT5OXc3OHFeyYAGNDCO2G/WHJ7Mdu1M2WUs/nYlqsB8Tv6nT9
DVjzzJc/joOIItC/xupywXCVz8FDoZ6/NlV0mTbymVfKDu1c6GIfmlvsJZ4BRJIa
q5PyqrgCjvirYRENO5h1hbljKsdGrluc0cONBiKsORrPk5znyUWTRpiz6WycOlc7
s+wg3W8rQoYGYXpu4GHEiIVNAeQww3k3uyrhJLHEZjWs6WlzFS5ucziHIsgAS+fe
qeIx7k9BXt1AH3nIzhGgl/Vd88BIV1q+3cnfaULa79aVzN9E3fvB29QvQOX6pzoH
2E3qd4e0j8EbspJmd4TCVDHaJgoyPBtwnRhUqUybm3fOynp0uBU7h1GOI2NQ3gsf
xWK0LQaxx2+Fj90FDbRPpbgkpb9Zd6GYacjsfCGigjkX4DuQOAom3QiHQh1Nhj2a
spB2uFvuZN/nVZ02krpoZlWCdloeJtEEFezJUAe3kjy90rjc6O5+61wI7x4eGtrZ
A+ozG5pRudAnUULDJ79iBzOYbOgKMerQuI1shg/WgtBqg+3S2Q12ByAPdST/338Z
HS29CZ2IjIZVkFH30zakQFHvPSOGJstrATxoh/3Kzo0XK0jSHGel20xe0x7GnxBc
oucpwjiH7Uxf2lcM8KgX7PwhYnUqqTx5jhBlIcR3BXDzn/67IFveiG7Ytai3aXsv
SGt8gLBUnD4H0iGnfHW52xGf/nBf/vtBlbGPg0oXYJgsN7PUcfchWAlr+MFaZlXa
9K0bVYTB1tsAKFOzTdUJ9ggzGnJ9ug1iJeMwxAZZNcyZOzWB29TAQd3jqSD+9Uj3
oH6n0iAIulSaZgAZkqIGDTAtln3qqBt4jtjYLubeX3UUc8wf2Seb9/z6RfdfF9QW
`protect END_PROTECTED
