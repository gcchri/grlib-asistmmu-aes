`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsNYvSfb8utFM7vhL4xdDGqnRuxpH+XIMM9K8E7OLR5bJYNkB7nd86tLNOdC8SRy
/+RAG9UO4d31yHEwunokRgK+3hmCV2Vz04DghcFhXAxVzLJiZS/jIjYATlPLdl1t
64+KK/R4Bba7nlSJMdm/Avdu8vO+B/XVF/u3YFw9hILPm1AGfUOpLEhzKJb4AeyB
97X/VGqLe2DKCKAlNNHj42fBeDaZqmMtlsoaeT8txC2RYl1on29KvBdYRdb1yeeM
XG9G9j7QPpggxlr8YZb46yZtNzd7rvQADX/yZK15BXzz3B2MxdpGjdUEKg4dREwt
TgkKZtu0hjOtp6IP7g6aF9hvmwMnKOdOCqaRUG5NhTEg5ZrQuCgRqbIn3uxJbIY+
smw5y2fKuOryUihZUkVKdM0tdIcqJ58KxSvnRUkkFpHWg08B6vY9fwBEzCm+yy0i
D2zszxKN679xCaLMds4y35DQAddiIjbWAkbh3brqfRIDk0mdFS6/26oKnbxOz/Kc
tNjYmlT5DfcH0Qq40/mCINZKyZilwwWffUlnOH/vxgAAb9g4hwV80T9zi2UL08rS
ADDcnDBIrCOmQqQW+2NeWSI4Ve1Eg/4YTPOdBqxQdoJo73wB860xQwe62/+yt1U2
6+nIQBdcnNrJ3gGMd1Vtjp1owH4SuBuyTB6k5hVU6G1hrROxhk2289j2e316jCSe
eLG3EMdkI9RE8KS5XWi8ccvFkiAtgnh0H7KkmqXPXsHc46y9vK/vmJ0k3ZeW8MtT
ZwpB31S8uor+fWRv6JqPYAVp5CkGblOhCLoT5/59D5QZW4/ZMAhtZnmIC6z9XYkd
KJpG/fc8LfpoqUKQOOM35oytiXfovpKu39GlTAn8H9NKl2Tss4goq4NQ3Fi4qhYs
kaIckK01GcMUfQ7ANnLE6cYbtlzsl6hxhXkRBDE7rlB3mZQuA97ktcKXKjnnAgjm
/ijf47akaWYv5P6to/bcWQR2dBkFT2IIPDr3zAgflLXC0I7g9kGgDiiuflkFVgyy
YWMckEli/wVe9dwKfXjeTEyowYb2CQaLg0fz8TnhaommEIGqlY1lqbeylUlsN13b
fXUqSv2T+wwai3G08ClUG63rBwSUpoGphu8SrHYhIpT1Kcy9gETdkrSOn9yak3AQ
gGI7iOsTVFiTYGNPcLy6DdYgGvX5sucQnhz5Jk4u5Rtoerpf+ATQ6iqRcC+qLaVt
Ov/5kWauNK2HQZB+tumTOQbwjYDmnQ+xu4m5SvcJZGAUNsXwCu+NLD0TQGa0aVdy
IgXf01s44yIzmmsGGyKAMd8TDb5UJTSNei+cqVTks9jrmeyfRIoMwmYU8ZOAdd8/
5yXGSDx9GwPTPDZm0MJTXRL1fH5WcVvjaQrwzJoaD8efEnhuyfrRkQWlB4Hy3Xqj
smjy8Whq0Og61uLvTf2NVw3pT1fGHtT+o7JPy7Y2Om77HHD9YtQLFLkVdajcujir
/XFYQXct6oS/wkIxIDM5hvnm6G6qXSlvr75rZ/Q2ISDOk4PqVrYZ5Tg6woTnLQWU
dN4AwyHe0JcVN1e+UordnpuW7WGAwEMH+nnlMhHJ5Lw0FxaWqGM3k4TLHAWFOSeG
gwtw/KqziPJ0n6rRGPUXvKDkeWXdYxsfPUWIGVnOS9R2GoGIdJQoOYdwEZs0YpH9
namBjvMUkWc5eTwkFMD2QX+a1mz5OUNUlZc1qyCXfC5PyNVJ2v7l0iHe1mgtRl2g
GMe1Dp8HxLuhjJeS7+wv9BQXPRigQciG9r+ZcJywVTNNTFyfilFD4mEPYQH9UCrB
QNFYkpOx1+5G77pLu+CbIai8dzR+aHG7dKutPXSHjynhvsM46g7vR8gRqwqgdL5O
FuPE2XaB+dCaK6hYh/gdFdDQiFlU60ISlgqEXclWfCstdqxSph0bA5VIljesyYM6
2h9ie+Tbr1B/v+Z520dIkHtTC+t1hYjyabGuOG9eggOG5oUY9qAPZPLG0ZjnaR94
eipdEJv7YITDVTlMsBM7EGMzVIZsxzMYFhPswb4nl2xG2S0ESqqD6dheIYgRmd2t
EiNvt1igeQCXquCLN7/4cxbfxUjilPUNx59KUekragBpviJeR4ZVfwGrzyrjsaPO
Ifm0pNPDL76AD3gdH/VGxAOgXoLPKkiY4Jqu2EV5i/4CiwY5S/MxEqj+w6JWKPaj
5wlQ1KvAMyS8qQ4dZiRVFDVuJ4TcyqZsmKewxUS5TnG2larOfVifGQSXYzGVMCgk
advfhNMkQnzMJe3WwAiAJQSzlhFFWJUugb86U4ZZzSjJ67Pw8hQd9oWg0VdBgHsE
FSC79Gkl1uBJx8/QZUksDQLhxN4ySQyHnHu4yXhquKqvXbDxzMyoeR6K9OLj2V2e
fOhzy4ftHDNEPZG+1mBITaa6MlpXPcLss1H0DC8Hl4TeizvDT+kcACYgWYYGrnFv
83j+BfoXarpVUJS26dj86YRw67BpL/7od/YB62ZzGA8f3HsxT6nQiAfVGVx9m+iQ
eooYZaBdLfZjXDNPwo0Iy36u2k3HrmaZ5i5qbMlf4KKn5IjjI9DO1U+Khxx8nEDN
STyK8QkDR15uzW0OOKrvXSYYIPp8wkAMN/CMwiJw8fjuEyc8pbv7szstQMv/cyTS
q2IOrCWLWMusrNTIrVBwJTWFvxSMLymFjI6KP9eJ9BoxmcXvFDG+ZxPA6+ec2JDv
1Hi9SEvQbS4+qKoBzzXYIMKo+vAlRd3kFSR+xh1rfJ5VFBeakhUQpMhUgImlDev/
`protect END_PROTECTED
