`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SnPdOfd+4kuO3Fx8QNFK8L6wckbGNfpRiQ1ZDZas/LqNOfDVsqR0TWOL0CxCXUSX
61wlBNXiVhi3vJPInNqWHoIGWvhOZgEnCHiBEs2EE9RJKN//w04QZiSWNe2kt61/
wvQhjkE+1uNH3MnYg333rNxQCTLj5+boYzwaEcr8PwVapiDRLwzdozo0ypnlITxR
5iwl6esYtNwL5GaoNMy+yc2etIcCZLDBDEFuflA4PVu+4+ZIMRNZdp1YhF0uD2rK
Pg372imTE6ZzBZTPf5+MZAKBC5MNR+e+DndTl1RkLWh4xcVJPyyWpUTPkiyGX/z+
hF1+dyrFPWQ1v1Cxc+CvTA==
`protect END_PROTECTED
