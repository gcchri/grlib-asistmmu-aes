`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R293maHEHl9Q+GHnMl2QSEaQC54JC4P5rhkX+nHqUdyR7FgDq14cyAuNEn/GCVEw
BxAO38MStzrxm1jthMddxxwnXPvmAuSswFvv0hPBwxaW6zgQqIfP2Mm+MGE93RIJ
3HfV+FXbLQZhLZg0z3RAPT4HfKjcLTQgEJgnZecnDQWXjg++0/LNMrJ7v3cKy3b/
9rZ68oB7rMqcYobZSMFB7mtqrHYfEbzB1XkcQrU7I4R+123PfgXx9/lH6H0q+fbb
vQDDYFEXMDanq+sJaLxsegKcjOGSgSinD0HzklNKLXo=
`protect END_PROTECTED
