`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ID/ReBl/5BI740xGe0mhE93X4b6gKZkQg6wo3LuQsRBDRLFNINsuOiCFL449Eo3v
UUnAizNvlQTgjFED3b1ZuHEGMf+7PiVl0xGPxWi1XwmK1UiBlGjTa6CsZtKbrdyU
P+u5LajtNKfqFO9tfA1yxaI+k+9SLB43jf2JwqFuIGq86b5680go1R+llaREVwKa
619TawAazzdBtBkGNkinxftGd15uT1rSR8FuPy5+80cXn72mlVIY/Q7RiT3+1OSP
BJ0c3SPpIY3GDPqHSrUeS7D7O0+uzmyDVoU+rY8p7aV4/7qfIxaRr49+zClYBjvg
1KMvujR44VrF0e4vJfvancTlQ7fPI7psbWQLLHpwKSS7srgwuyarqJhoMiOYlQC2
2KU6AIsZ1w4Hx9VsAbWTzmUG/28/+VgONrzEaauNNpyLXsXzEuAcV1HZERTsJryG
lCmWg5CV9oa5H0CijGvjUyxPDY7qtNKIT+iEB3jEi4NL5Yc/Sxl280LfTSrBAj3T
hE3yW5ellloNCq/uTgjMEAQffHePI4dNW09ObBMU9bXPd8uo9P69zWbfypj6mcQR
OlRZnENMfmpNqscXrc9S2BuHm6zsS7BNro8Lu+3udAGsPZVK1pcElvYo9IkVcxG1
HafkOffTdsU4237rBohFU6eO91TLWoOTP9hrGbYrYM50Ly/8LbYMmT1tCnB6V39t
pYw7Q+mNKoohuYY8Ju+Eazsy1PvGPACauvCmti81yYJqbkci3QOsCdfGS4E5kKyD
eyIPpMWiwmukm7MqVBpLXbpzEIG+ctLX9eWjxVU3y5Ns9xQfTrBn3jkPgoVnzasj
QRqqeGkYFH7T4pr21OmVio0DBXW61CuTiu3guUbQBSl1CAH7PtnuFR2FOgPlL5yT
T8pR1s4j0WOzlnOBZZfGKlACnyz0qpPqtKOty4Y4voM6exNhb5Z7U4aDlwaQKtLb
uGnekle+WTe65eUfvmj4BRE3adH9TkcWmzfINhr2QbNwNJG9AAZlenqXCxFmCb/m
Qx+92+VE1sCtNB19awlMybAPnaPqInpZC8gNmDxft/L2OpDVhIRNcWut9KZB3lF8
ueVQH0vdARFw7GL3F68Kkg8Ld0JGd1U8TNcdufQ8hxiS9xv5E8VJDx1vfaQghTEu
+Y24yXNhfk0lDYbeKhj6O0xwwp6jKr3xiHD3J/plUVBbYatwcXIQ+uwWByc58ILC
0/1Au3U61hiczngsocK8++appRoLVPYSmGDtf67yOaVqJE1VQJz9wnetQLd/BOL1
wh0twhledUKWEgt4obhP7R2PNRSCVVc5yG93IUmS+kzC8E+sSstxjbxRVLkg9EcC
LI+IrBTERGxiiWAibllqEBkqdC91xsMCH/Eh2bSJPzD4pTsvBB1ZJs5FtbNzGqXG
2Cwbw9AdWsQhCfRmLMe9nCWZCmTp00J+I8kmW90MKHEE/MuL5zjq1SDKJWq1Ki1x
InLMOSayLPfYElgIikf5FmbN18LPlNdNIBVykteFgJMvZcTuT/YYOstsBGKI018w
XiWTirFCLcipknh58bQHvM9yjIjkAfWYkSSBEEEpTx2fT6tUUQWzAejtorwL2rCY
mRGtN1dFiHi6utb91O1aj4KqOFvt/R4EiqTLQXZpkbbywGDPFQFl/4Am7DC8zjLT
sdGbCvtQy/F4IAjeIPrmsvXuDAK87jIYmTruFQ20wMgWZe+AhBMs19mIQaiUVP9V
KiwI4GA7A0rIbacgwq8KT0slw7sQ6GOBoqmT9M7QerVma7ofvFxMNsSLfsMjVOBT
9Bk1q69fDOwfGDdd/sW534OibfXTAUNzdLcHmIIYS/GsuQbIeCdGlU4r/PBpBkwD
Oyx4OVafJ8xmN6I4HpIRhINezLZICFacGqSmuyeRXubsEkkIaJOcmYnSbjuo+4Ts
ityt1OSUPifMcfk9rMNuzCbKZZ6MFeR4nokEtW1/WZkUt0VsbQt0dwibT120dP05
Nmst+WMb12pa1GYsyAs87x/vNwCJS3BHOgs5XyTW04bkvWPKENhDU+C5z2q0q+9e
/b4UIFY5gv+Ps6StN7G6PP2wWzS/2jRafjQMBlYAXAGqPi7CRQbjX0vva4muJqVy
XVRTtbujXNmtEBoqi6S4F7MABYDFcxEhQvGOpTxDTzpJbRS3pIx1z1sG5IWDbqO+
KKHdRAt2n4oDmDqdMNgj5MXh7+NBPvrJ3g/HXr+vSdMHlpm3PjgiH8AASGplEnXW
42jQHrO+Z4iatBAXBXLlVyLPjvMYL+0vWDIC5ggfhemvvpl11LAx+P/oHGAGu43D
SU+xmbAO1PJ0FCua0T1Tgp3vlXRzxokEoB8llP3UOp6bDD1kghHk01agTwm3dvA6
IjOxhEuJjnjAVWmyjVPWG4OsP+3dTHLyQ1J4eYA/gcuHOuTT1IzH+RSqbgslnFYR
ENnSTK3LA7LKxdVEKFNOCWXZ1Y8r5zkhHl3ZHlm+bP469T4jUpED9wLAWVZJCtDr
DWVQK0lZvbvqk8U/cFisKGHhNHDgp55dvkuy50g12MPQl7sEjVj0GDdy3yNdGLo5
5I6vBMldN/Qe/XLBs98qVzWp2+tuNO/kK/ldCY/BQaNiTI0HQMmtIm9/rD4TwqU3
Rr2s1I9nOToSnre0zETZNpcfnO82TpSWw+WghIRas0cwP3nf1JhJ9f0rkyNK5cUV
VRbQzPZS0pMKV4YkUyGnIJB+dYLM3IZ7x0st98znuywAAWyvROt24TcdVQ/9lr/H
HcgzJpII0f0sqNuU5ycvyZ2Kks+nhoB8wcqvtZkGZowqMyM6L4hA6JEPzXyJKMJe
hBfYqpBxbw5BGQTDQaKVhKQvxRJGCYXzeNYzSLS8lUNNnfOuKej3sphM0RmmTkek
voBi/lxrVTPwRa5jYsl/b0WS6jAiN2Lyfje6/gh28gioi2JrUFB7gGCqQq7EjVF1
vlhZNG6zhqK3C7D8nP4hHTXK0pk12x7vZkSz2/vMPpuwPOtcoA9F0KMOG4VXgEVh
gK79JiBI5krFvQhK13LrZkcWc0c8Vm18r0Dap7BWK1n7TMpVAIw+ZoM2nr/ETo3v
KvShwRtjl4ya2XeeDomq2/KuHT01m0JLi+wa9/mTs3XzuAN4jegCpcSSSC8uDuS6
LWY6/rXAJkpX3YzvQsldAZS37CPyZa5AbD7FXScNsJ+6PJMEIqZvwBraCHFIWejS
ja6Hp6BgDf6DCkRNEjjBhj2z8Crj0OCkcV//NH4xpX9cfb6GFWTxeIwSnBzX6fxk
EZfvNNkJBHsdgZ37+XFi1hAfkKHdcl7R99yj2obR1p/bFide8Xsbl1ij0tMpIyt/
/eWrtnEz4s+ZCefgfO4Ujz3uD1x8nUDm+/TwjFY4Q2koAikcwFNWDAu9kRnT6Phs
wQRk6/BHICmsDLsKpMTmE4yinB2Bbtykh6FBv4R39E76jWG+2OnGM6WCK4HpfAQf
3yI91yvLQsmqYX+K99DSigcPJph26CecxpYqFLChxHgsAuy0r9T5Mc70Bxq+vjh+
zbuGlNTDbS3AMfhGEER7uKkQ9DPmV1LWwbVPhcIAFZ7thJ8TPwMnUIfNtho9+inN
Yh86VwkFIjCz0QL3CtozO3hqRuO2RD6q0RXiocGrBl2GKcz52lMK/ASUW2ZFRs6C
jMxbNN2wohi68aX1N7jJNKEx6v4JwF1Muty99oyklVCnqesTPh+SJTVYDi9+myJP
Lmde1W1+DXhCRiOoIt2V9FlP7IWB2NTBqOwxKE7t6/sqRO/Itzo84GEyvsF4I8kD
TV1RPstIYjgwy7gogPLu1CeGCdAPDQ39X/oQ1bMzL/i0c9ZYBjdSHMumFdlhxawv
ORPyezWS49TYBHeDMqng24AJQP9Q7XBhhayGHsQ4G6+m10XXIx9XUxwwFV/YbkQL
1dkUlIZqVfLMiOu0pvbo+aKIgwEvEdIdYSf44ZwUwtigp1wn43x8MfZZIlUWrJNm
5egOwfrF83sKMaaGw3YuZRlojO/hXOI4prwQPboR0ArdzuxcCJ23XfvOmNN3vP1K
snloLau6CwsmLmtdN/N1QC/T0argPtCFWADdDHUthPT+xHsWXh2uZyDkFxM/dlRj
a+FtW6vduvgBjxx6NTQ86SsBB6LNnW5o/Wpk6Hpw0WbW8kSTeSfs//R3DLdBRPC8
GsUa3OTQZArAhNoz2PigsY1VFOuKEImTXP8dFXoa31kYMVOyoz8qPhs9ySGfIDzZ
+bhRRXZJsockMLYPf0K3VSgTshK8b8Egz4zHvc1kJNVY1tRVx5Pspxxj3xk+fIV1
tMNjGATg6qZjecIXxzZwjK9xCCG+DITNFJUE20S4ebdnvy0BXg4RMzCdU9CFjISN
c+7abPK1kuJyyJ+bExyTGQoeKUbqWuYoksxGcjlrYBuoWSKLOQyjl6/b6XVAzMkR
An1FVJ3Iw73LZPkjIFdyx2usVLCwO615TZV5PhsMnHz+lF5/l7JV/i+46MvY9nCQ
k89T0gxj7yH7NusW3yGmRjSNmlHP3Cs6+GxBi6NxuwEGrA/MKATPGRd9WwQlDK6G
JUx3RswvHWN99epluBCk8l2EU9bH0VKvVONB7kTOd16djTP3XC+hg8lBTlDHWHZu
rGSy4LHk4Fq9aW/vTDR1LxrBE0hvMueSdXrG5W6cn/o6zohllMDHW5mDPnuFrCln
x3RZxdzxKAgkZ58N9E7itJ6mJ2grePUGdM8o6dNwwCcJNCCjZ1Wdk3OJIdNHG7hg
B00Jsm17Py8VV30uR2etVQwOzvsQ6z/K5Kz1wm0VDsAmKfn8uQ5jqAoEXCizLd1Y
FtmhTYkwDRuR/BcrHa6r8QkYrCrfsIHnoXPV4lC4ShXQU3TybdolNZX+kIsKOY7l
cIrkHNcTSISy3t/iitXP9kyxZFzN1Tc6ydaYMH4iTjK9vStVuv2PTlk65rAcjdS6
rrx3sy5fTL5hhJlhcs/1g0pzulI7KrZ3LGj2FvaJt/X10yTkbou3rWY/Z53bUGUk
jUQ0CBOmsT64bd6/+QkmKQDMNl7amxBMHJGFi2scDj6e3J4sp2ooI9/psIAWu2AZ
D7XxVpXS6ZUwJdVOmuJa5sl1mrKVy5LOWoM+klzRbp7RB6JzxT+jlDIzCv++9ry8
PKVXjDGK44jboSTMtuduDSt3zPgj3nZ86R+rNqTTyb1rjF3BSkfnk7F/d8Xth6/t
Q4Iu22kgbjVnnPhqMwNpMgRDEmQHRBhJaWdkYVx/vHkYgEh/IDnJ3a862M6/ZDFU
q2p0gl9mF98q2o5KqfByTVpEXT2e2LsfI5n5GZhHFgO072R1lmXjZgyzQRkM9DQr
nfmUynZyg1W+QrTNLPB+ChPn12ChAzqMoYNupHEuk5pnOk1RRbxK7W6hD92OfVJS
9abWDGHdLcO846wT+zY4FO+hANnTkr4iX1+4oAkdrV8GlnK3LRktIranlcp3ydsu
ZNAMgCwCzPyhG8/H1NtrV6SAWlU98iqMRtOkR37L3rFzRvScrzWxG0QjxotbllAb
CGJzNy+4OzqEOe60Wqr0+omDFwQ4InIGtSr5JT+rr4qaByxZw8E77XxWX88wyyE2
+IcxQX5DxxVu3ibsMF7DWfY0lK+Brg4XGUo7+BCCxZFSqZ8avqieuEo4RGyKVeY3
HRPbDIjH/aBngy4RxrrXptEy0jVgr/cR/I9DCltj/0YS7TROdMRoA/dMYv3Jz1lG
CqvqIrOQn/jeV9GFdYE+qesgjpZ1YrLoXWTWl9jfMi5gAAoBpij/6YFJg+s3msMc
fAVEePphC/Cj/n394UjF+ut6/VX5MoOMmV3j6RNqP2zWrVy2zgTwBD0LrAMcECwF
vxDNTiB4moxOrqoq8HuEgnZ658gH8p6+/TqRycoelAFl7/XDCgTvw9cErZyVpIPi
2IIlJR5AQT11iUHzNWVdP9mS4nQ0Thv0fWFxfx8e2Vi5LuKh1eLPS0lXCK3uTUCk
Gxx1pzWE5DK54DnIN0zsdCXpBVlhAA07W7UpxcRHpnPv7O+rLOhevGjDBhvW3JLp
iOxgyaWX3K89j2e/N8svEiPbFBfYtXv1d80E1yUzOqC9Qcj/y7iuYAkuJOPtseAm
EvH0hOq4QZ+JtpVAwsUW04w+pbbs5PJj3MQIvjgZXsaZMJjLn6uBB9P/FbhTk3kA
Ops3VjqGz4/AIpMzn5pVgy+j64BgFv2FplRwbjQiTlAcYfxFPbPNGgbABfxWWkZV
GpE8ykF7vQJBW/iiXObZtrX4/YE1xiYmfubjL/ux5rGqJ9HbQLz1nECsN0VKSAqC
wAH0k0eW2NLP2qlFTFplQzzHo+xoumh0SDqKUdhEumyW3MvneW2uqsuULx/J6qcT
U+ArrfmADpnDkPIrhJtpQU8Yx7zy/+rNWwmKiKMDwGRiqEZDonKsXabMv4P51iZh
ETesEonEE4qVwnuONJ7ZutOF/OxzcDlplp3ndPt0O6fHb2ijIU9aDkaaE0r3WhAS
VrabwSEeHkK+eWmkTq6pX5BwFAPhlPX9UZIU4aERE+kAEFnYAAB2ov/KbzWbsAKr
SqBlBTCLJ3ge300j7VFvQCKuOPqedFN7DUILjFCzO4lXk7xOcTSSSzjFCY+ns3nA
txOv1hJvJ/IqeWAI3NCSKiKEhMLKg6cNN1LRXUSUIReQoNr22KDQWefpFSXj2I4R
eTefqqVA7fkTZnhUS8mT888LfjdmjNUeQTAZ8JvWYYhIuQ61oZJLiGGTWsK6DySh
aAKqxomC28ZPRRxFMB2maiqNfZRHuTdUPCwj3YaJ9vUnXes3CKk3sQS9G4WfGRS8
mwrN8eXbEGj1vCJ710mJ4DXgPHI61nLFpm5b6F5vIgb72YBONo69OFq3/Zah7/HC
YGWR8x2RA1vd/V+0m/PImuFkyYSyxNl75GiPkqtSj5Xb8kx+b+WoeOIlTeq+RzI9
hQT60WRs36kptx5uJxLp9Xh+dDqAG65hpoFyFtm8o4rnu130XCDDzY81z2+cbX7t
7zQHrSxjC5V7AEdPbjIGRoNT+WYS2WFzYI1DtAhsruXbHi5cn8Nab+il22Ah9yQr
fHUU7wH49IUGcN32ziwkQtX1Y1MxkYWFpULf1umYokrJHApjKmaTt8TJad+uB6O0
hQ1Ojb0FE758i6m3S5p5g8kt86RHlUVcYEJ+xSM3CdF0KXBf2Swi5ivp9OXR4SUc
FIcn8C6KxN9L0jwy1ZT7GcPILKMCTtiRC0BziO7GXUCZvk0hv0C6OnsUMdXRGh94
x+KaghG6hyWTYU1MREerQavIaEHRds9UzQIsDMIFu3ceNqIKVbSCf3O2Ip0DiqnP
f6oFQQxQxOM7txI3WNA9CSb/chsGv2y7WKrGLfE4HsRx2RmSF8VtXgo4/yIm1lEL
/FZZcDrOI3p3zMNLPs6NzyXPrNlSKlCCy927Ul1msx5ygkR7T08qz3WtC2TALG7C
2JWBdbSojKYyztmGFa/NnP9yJT3hn0cjEkH3r0AM+wjmDzZoFnZ4LorWhrtOVPmW
uYNe0U8dCCFUIDEaND096+tuUHopxIkWts0dL4RPgk6V90sZtxbh7IWuaKBPLfVG
IHD+ysZWz+moLXX9M262IQkjYAaViybd9tHK9FfFSzdiU4Rr84DmqIUDEjWkFGdb
mH/jRgq5w3jzH4VeI6oTqDC/Y8IP9SW1jG9LLFlKy8IRKlps6rlaorOg6Gfto0n9
MHDFYwUqbAcixXlCnH/9HNCGhX9rMON1ZYKfxORD4V5D2oska59EGJVtxZySAZ69
Ib/KSyd1k3999a0gUeG7C2Xp8iC8ogrdiQvUAWm9gIOb7wsLDcTk0tFiaAHOw0Wz
EJ5BTQlSbERXQTcLfIRCtInoqAZnQWVDeMwrauhbB2SgbrbjChEKbZfMtVENEtle
vOZ5LdAugb3mk9H5gy/tReMrx9z5GF4RivIBBn+d4bNZHKVdxFWWI2cC/HEF4LrB
2pVOs9aybN8PW6YHuDrzFxpSgnbiOWpNIjoJLprRshAY0pCT6dHfTq+T6z34Dy7W
YHYvXLv4at4XJ6lkDN3UKT0QxkjMhrXODi+iv00/2372X/Vib8cw7Wby76ys3gX2
s3SkguNTaCTxy+1xeLe75qZ+kCPhDJTLKDzOgVHFEVdVdvU+Fe4gb3jonNBrSXg9
ljkIEMeaMQK3x4yyGkqXtal9F+GvYJzCrdaazXxxsAnaDAsAVmM/bGn0FCNxX8Be
9zXqEwYTUrUB1aZ3y+71Tug4/kH+wn+1cgKuxTK/VFEpZpOB7rUmo8aYLik1LMb+
74Yub6LNAjm4NFFuCBPphHMbPLF0vCs5fQEIBBfuEbugFDgAuZEBjQgaGCA6RANp
CCbkG34yLKFBqX8bus4rNEPRsuubn8FOLsO1chwN/TSj8wTCz1JyEj/fSyD3oXNh
hkDL0tLVU2S7Rjpc98f/mYe7pUpo46RfK3dc/LEXQ2s0RHKt0Z0cknOwGp872JAB
UeykBcrBYuk4i/hawsjG8FWb7SqUnne6vuz4faiUAGw0zitRNqdSgk9KWQFJFikg
6xvgBk211BTX89+yd56E+kD/rnjuz7E9oDxJmyBqVhBTLKuXM+rBUkxz1Hgl1q5M
YUUGPsUzsT6ISBj7cmWmeM3guj923KPPCFcaI8Ef0iIuCeyzc8NZT6yJdHc7F+h0
YhwNtx6IEUYTcImkZ2KMlpKJ+v4Fhmos9473Ou4jRgTHo9g4mIhEN7LFCTnFAT1R
fmxZHd+DQ9EV1EQpQ4P34qYaQch9qjZdsF4QhSscWvpK0uHcDWnixlrtTqo4WN1m
tXfV1SM7e1qGJm8eAf35EYA/7tNd4nUPnx4qd/87krw1zXFq+MH6si1cL9BetW45
lDBwLPKkMqIsAhphX3uNkuYPAl03ZC+Ty1akxjnGbdDxck8u1asDJVk5g1OA5ySH
ZKTSJk6+xj+kzz9ZWS/Qqlv1hYRrw0RA618Pon+1fb3h3gpARC0IILb/a4BrKeqX
2d39bP58lgtVjlgPwKHo55RU9bdo8E+WFJLupaJ4bH5DgPk4KmkBJwESORIZhQ+0
BFexrAz8oSE96UoTZnx8m4Ol98ZIP0SO4hnAmTgpZrrRbPVxx1eMenZBV2PYJ4Gs
l7cQ/2uJt5Pe92WxDvZLutBAP6qjxlP202NCTlH9jKoj90WRuzFw7aKwU7PAMjye
eJtkrYPHo/SdwmnSsqoeAB/eeJN9wT+DJ7no3KqGY/dKGwoEUHYHTCXFpb8j+zP/
IZX3ngCISsH8caf24WzVuqIEoYQj1wcxxOM+GVGqTcG+SPC/Of7vQPwTbLXjatYj
DhTzj4JHjPWMqPS3zAZdnh2ryDSea8O3fTgPqcUQgQr0DZiQPIvUkdAEfDwY7yKb
2zCqIRGpSII5JOO/8jTZn882rkGCNbdh5A6+IIPT5WQLw7YCq9zaGveubjzzAUdF
O3eU9szFunBKxsu7NoVSzhh36RXOQ2p7oBYdaZn+zx/IAOSw6L/pkput8q9c+uc8
p9XtxRmLVPBkfHdF9pp97wcWBXSE1NmAZr83hz8m1fH8lvtpcN4Q1vQsvqgnOPnJ
9FTnhYFhHQMCoARln6uTQwVJSmCrGHNZyU7foP42AxaKhwJfPMeV4tYOppFXw5Y1
4BP5yIT831B5QfIALXqv2FhJ1WFPpV1zZu4pl3GBsto6rJiueZYqVwLsXTzd4m0S
R31Ecg36FgNACSo8MhKFOSfknrm8BcyliM/RiK6Sf8dbbzOTe4MCCRBkegUGDmHJ
hG5OvOPNPnXTa6A4mZKTlX/Kom0U95svo1IZ2GRjX7Khykb8rHq4wrF9aG8lTz7M
hPZ9w5Kr+T3dEigSMWd8PZHd1Y6sob7i/OnrJGJ1Lt5pQvc/J7hFgf/LOgE9Ur3z
e8LoB5gaRAhmccfHzCp3Aqbky/Dh0bZnzbrg3qFTOkthclNObBlb91vqmgRJ23Gc
pLEqW+jDXWRZdjhvpfeXSgVw86WnOLXClWk2gSYDgRp0xEMSLawafUsXVyuqmiTT
mIq6wKWc7EzCabgjjrRdIYmqjE5nQstK+r43REZ7eHypQkHbCIYN86vFAq4O1J1W
rI8YCpSDuB+LwSYgAFd0FnsQ6ZcNvUoJ5k4d7u3YPtruriiJ+Go+ZlDx90KnEqoA
C/b8SNSl9ZL0g+yXLnaNKHadnuGs79ozyVG1KzC9Q7hjk2S8qFbG83mC42EA9+rW
dS0gon08369w++2YgcWy+3YMRTtJvr0BgQKE+f3brIeA6w4EJd5iCTBPDk3gebpn
3Ix5hk1l38OXt8ifS4ScKYArvPZKNbGKX5ECVVihfsDWw0UmuVbGTg4Lzj1X934p
NFpL7R0Zv0lkuYTI8HHjJmDRnHeBKdMO0FuMl/fFzvhOAwMJpqVfzmi4vNvA1ks5
EpG0DCpuPfpnUyY2VKAax+JTR2+cE0i6sEqkOemBxJ0Obw0alwpHiGGdKEPRXFtg
c2UGYAbFCI8qeYLZSW3trd45hKCTQ+wmz0/oB5AA7Os0FLFJxeVUU8VTaLZtbNss
2IaLFtlUYusfSgW4uYDdpgTvQFR6Ko637l39KH9wilOvhIgL7YhTArVuGTjIqeGp
GfMZ0cUEOaKxKFK6CE0ct9S3ew97GwVBHiIijRHWDMrOTjBq9efA77awLaxoamkw
R+vdqqvHMXU+wsJDLbq6z5CikkhK7ihsloNo56nbC95oD3bt0wj1X9ZuVPXW0S4k
W8iYwFYeiuOLInEQNZHEp4RlRVr8yTH5aarh4o/KIy+kup7SYqVzcFxCzWOAFd9j
bRJJKhCwsNfweSD5t+rMIIGbCLko1M1eH9Abeu72/mi5e6IjYyXa9+4NAYZsj/PX
yz60EroHqn0Pn/fhsMzYco64vZDwKNwnkCyrfQvywpDVDyfWuPkNh/PmQhUuWP34
xkvoTd2pbaDT1tsQw8VtI3Nfg98ijBJxNKpD3dNrLkn4/eRfn31NQr3rf1+NvTfm
aC7sWWsw+f75/7Sv/CLMyqczHNVCHJDOarMiGrnzg2sKQIuhws8bsuS/IbQxtF+a
PSpaKTsGBbfD7lLaicoZDZWwb/4nVLFbDl99z0e+lRQRvdSAESLldsMna6oloNZW
oazm7J1UCe4aU9KWc7WjjLbD4+vD78hF/Wzatv0BHzIcGFw1iVb8gut089Mqv4fH
P4I1jUvPzARHvNJ8E5/xLU9+hr2KK0adGnHocOIA0l5yJlDMutpwhfA3Hk5wRL1X
s0Nj/06Gmv5Yx6FUrpUAetdC1kOwnXs+3w5fQn3bepG7Jet26brBPVGGhfh1sC/1
Ni6pxOggmn/+FF4wCv+voR4CbsqGntWV9LkmY/sDfx/Se8f54bQNfJ6peac6KZ7K
+TK4gwVmFg7FJQJ7wW/5IN2rLElPE0qPeAdpSU9zfDt1HibfGMJjMKzERiOC2x9a
IZ2tg/gw8qJjx+EWECosG8FLKOD1tMMUgOpnuUR6EL1yXOUUJPq4NrPHfmxfgcBM
rzUeAqbHLxQNIwQB8CD2aLsHPoCvrhSgD10xmE9wXS7fCkQrqFwS0sUqEtuFXvOg
MX3Qb9IrcsV42+5EoODgr2EZ23x4p5PH9XkheOe6VMmxVNnA7dW7ii2AHLFvxgDS
ZIySfmtdyWuUc78e92a+DyZVqEx8tqj3c8ogvVqR6Mo=
`protect END_PROTECTED
