`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VS+cstJwO6RZCwgyi8wjnFViGNL10M2Vg/ovBfR6h35cAb2U2mmRl/a1oUrgwVYe
+PflGlbJPOdVf49X8QSEIbFm1tltsvu9j3EV5e8IHyFIVKgEJlimFcoSzWyUJcHu
2ForIjxhQ9SuBRUf+R8UPH9yaYeZEuLfqfvC6DthRYK/I8AYd/RYnRnnULCQtGyP
rmGQLBgO+Xg/mWVpSaGOFsIGpDbj+H5DialfZHAWdhwt+u3sfqwIqLLBEaiBBHpL
lG0EQPZI95kOfv6NADdoukNing7cYhhDAX1Vt8qw2ewqvHImyS9eZoPBAMNbSOCU
gEuHXbV6GUg95FYc6DgnFGYMLI+EZp2GwgW61f3z9TyWU5jdNgOgQqk9Q5Qu4U6S
/VY5wpHwmcOWX0zpf56qFpXG3qjaGLIAxSRth3GCXSzDHCzBaS7xdYibk7hIkwuf
cEEGmgpuqYBiycvMGCuT6g8Ti5f0hOAscQ/ngJydRAGs/9SAw41Cvvg9hJS1cIyz
9NjEjSsUvpXNIpjmjm4x3eiSbYBXENdLchgfZ9eD9kwHm8KkVmeiVa/JsQVtorv4
Ggwnoi7UKXZ9su7uxnt5CGXLibFxqviRdTXHRIizQFeSZ1xF7oZJOOhVTO5toCeo
2z4znlWlAyZSDOgopoK5AmdaB0FRVNE/Zwddl2kcNS3Ym10i5xslJcEN/sfEJRsr
hywN3ibjhzSPSQB6BRBhLDEwllvV5yZMj6WXiCHBdH+ABa5x7P92MgdTSy9V/amo
utFJ+CSOw+gezqgZrYXtrehaH+dG9jpPI2JRE3d3mOUvKDU42UKYfzUCwTjMPkxv
m1VT5cG4hZ/N9ZC527f6BJ2b90aesmTu9KiCutemCgh/U+vkr62WfnV+g+aZw/3T
1dQIX8Lq1ddPDT8vWIt3gPVdUDURtW4zS8Rzgv/38B0vssZuNvf7ILRVy2zHR5Uz
nrGy0egshT7UFgv0FxyN89/9N6KU/unIRV3gTxadvApCmb1b12A2BrCOjAQsB4iT
YPCZh4YCdSwfiAa0VQLU5o4T/EO9RJAKWpHk2rCf2M5itBdsJ+jDYIf3v0DflNNu
cDC9jiv0FCfTEwAH4sE1B77hR+nrB/X8ET6FWUkhEle3Fpe4Mz6LYNf8Af5wjvqY
fHuA+/vDFMsArM8Su/u5r5tQpYHX0eVtN/C12BvyxhgjOdT2wGUi2W+Xh1wZgYn/
T13esvI/cVp3eA1g/TbdpYAiXsV+EpXBZ5AAuXQ3YsEiXHS186iniyjAvWb8+H/s
2xvKqAMxSO+apcxczP9fhG4hC3REwWBeWkmStjsrUwy5HJIF29CJuVUda8goXe+a
DuGFh5krV/8Flrp4ppjqGAEq+xJTTfj40kAMdYFtyvyAzzuSaJ+UYLIB5S9PBirG
90vcChu4mbeYZ2+AjwFzFeL0ndfPOjaPOmbi7b2Ht1DUbJNA8iUWBGh+HKhZLexN
6wMZ8qr6aYQ6rcsUzsZx8IYqW14dUv/4VeXcSYDOpqp32DirBBnCWwY41ZjIjTY3
o2duuS2psaniwp3aj3DjJaMdeta/Lc+2Oz3+f4ZcGkc9BlA1rtPL9Au2t3hD5Eqg
H39EPClvMISh5TNuqK5vM6Dg3GCx3FZ9EprTCyNxFCZ3MFEFsn5XrYtxckVJuJrn
wr7YCzf9YXkESG/3XMUEZd3cvIroBIrW9WQvJWAGK201gfM85huBn+8kH8bfiRFK
j3PcB5FVVOZsDXIkGjd/0lcFa9qMcBccIWgNnsv6W0sV9ySFXicNcmZFyOirfZhG
o/LuPBST1YYpUGOVCqsiPljrLIwk6gu7HheBpCqrPoPnw9LNggKyaW+y6Qy3SaNi
ow8eXtsTsUfeVEc2Rs3TC3vlNxyqYQv47EUQqu+4Z4f1wv0jEy2mC+dFNjfjCktO
GXKbpM/8cClCfgaP+/ZwWK1wRoUKHOIqBXm4vtCcXa7Af1YJQ+B5VKiE0IpDJjAF
vRN01w/CH7pamvc+RhDo4pj/rm+JUqIo+7uvDCRsOamTw2FMuNE+5O2xJVmPivha
HY4WwGxmRZxY/Bj6Xy32NoShV5uinYfCrkOAxLxU5x8uKrMIpJrWcPdop+i65a8k
kPbb/xoOoqAOg0G5XplWB221Eg1EMQKL0aJv5SQrvKwlDZVkQD3CfoQgag6b3ISi
6ti9ch5Ja+uSUATs993st4uN4rMLCa7/f+lAsDp6v5+eXEdBifUSUAlR0C3VGddZ
cJJRAQCH1+e8D3fKG0iJc2rVCnlYiAbdnoE7Ubm0kUbP0G5U7GG9yC/FjeYTM4Fi
UYynOWaRH+WGz96rb5mQAfi7oNjtzw6mK+z5WKMPQ1kXmthMgKs0sQ14C0uyYFy9
C2i/WkbPMW4mWuppa9uRuy2PtavJh0nfCmb/iN8stnLgVruMvkV71ymq0wEdCGC+
XtqTt4YONS86viiM7kbzDX6u9BybXpCK+x3qV+1wLNbHnGCpjFgAsLtCgP7mhfpX
EL9Xur/LGNlZcxxgxpk6jYOa3TUuiRA5ZQqOZM+CeN4=
`protect END_PROTECTED
