`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xnury4FYYv35OpIALZPnRp/iAqKeiR7Ah3NbiC9cRRdH1Ej7EFwzFZjoXax7cg9
KB2azFRrNK8XORXvhMJBVydohzOxRNf0oPOAaDcocAEhsgI3wbXEhyEdN9Fpzlw+
wveXtfXSdq/9B6xkRCJP6MEZAUl6m+Q22cSFzsfm7nlf4mfroe+hGgd+OpdbUPZO
DiE/8GAYms6t+1vvp14U9fnyEoLSqZMudXc8RgsYHXFNacjZJ+0DMHgu2Tvlh8yl
uoILul3SG8tLqFlN8AyiuZPD/7mzPVmrJaqXOW0BzToc8+b3yOYfRbmJitHN9SeW
aJ+bIUbrw6f1Z4clB9uibIVK2Sl4XrsNW8MSios6VNT5J3+x1XzcVNsAAW4UoX45
1EEsodHENza+62QdmZdy/mpjKxFEaIg+Ici7iAJicP0=
`protect END_PROTECTED
