`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sho5/8uljgr6RwQhwf/SQvXZ8mH6PTUFXwhjJrf7lfQEgzkGbV144G5cIwmeMqek
OLTAzq3oTAdWhvdsI5xRoVSSmLuCR/QDo973LRAUmGF/7a+KTXx5KD72BDqbilBE
Z0TGbWu6J5X3mQs2JRGcsUiGMEKmcsTq9pJuro8ERiCKUF9UFh7p4DGRMiCDdas/
aM6lunrG+wTZMhwET64kmEELlTH/nv+xmkWAX8qO080Zg8+fPjZ7I876wKrgSgkQ
kwv6V3cfGY+xxYy0MH9DsAm4eBvS3nqPe1Rw807gqqF26BTRq0dPpjeSRWtUehpO
YtTCnUDEeJIPtpAJD2QNRm2PJ+Im4EPpqJV4Dbf7PugFJLcqevmnFOnyeYB2UQ66
/3mmWnZbWA/fVVsJQZLlvMuYukwIDj1zD+hxzbHPi3YoOnthXJ0Top+PYAcQqWXD
oEMk4but0DsIX9vZ/1HQ5sQYBDNitUc7wBD9Ks6GSXAQXg5iGSC9P/TziHz7QN5s
rP6VeOICd9IOgawjNTVcmeL5oVjcR4UVKYSWlJOM8sE61vWQhg5rrNDAEgv/NBSX
JB2OE14MY0LwJh/965NNVg==
`protect END_PROTECTED
