`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFoezUREcPWTKdmK4llRlKLtjUuueJYYetitNGHs95eUUuOafoGo+oHm2HRMva0n
m+JJSWHdxB2gSdDSnASQd+PKoipJvSjwpLCulLP7CHh9QTWNrkiluY+5JWiZKuJF
w5xh4uAJSu/oBxno72bYfK5S7iSKWyHv9RrMzxDmKwORKXuszl4lhOKVapUPER3a
4KxLu+rL4TNdobWBJx0fonGnz+NgusAXhlFi/18dl3c=
`protect END_PROTECTED
