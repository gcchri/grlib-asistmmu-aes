`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RaN5yg/d6BvXyrdskZiUqKTAIxxmgNye1gZG2QnT+UVh4oOWsjartGk8fwOxKeBN
nVz1b/udgP18PIlqOCh2fkGf0J/6K+zaUDsgRsAtaxsIE/4k8+mJnMEbt9kWhR1+
YKpisKLvD9KHrk3JXuxl9nmUkx4jVtTerDk46qAvP/xzaFA4jH9qVSEnBCcnZOwj
LboDB8VqLXKbz+22rbal75mhalsmgvfzDOinzZthEtH1m5BRqVtg3SorJRPa5A2w
QgC2AxEFXNS77GLuNsaIZCAjdDBxkV42oFECVyc8LkA0vBFP+g6fMOfKE+U9RCj3
otxSmR7BjSOhloCesFFaIFsGyeSgG++KRVSNXfTDZG029FV8yfQr83iwVYFmCvfX
WmfAPPci6Omy0oMDmsQcUQ==
`protect END_PROTECTED
