`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U0U3t7fvSzAfkZek7xpFNguVejg/X2F9G6TECDBRT/1JXKlnpqBvZuWf5a/DOPcI
gm03M4LCVWhrnablPFjoMFC2gGF0uiES7L48TwaFCF2HwbOCVXwEG6AqlYT+2jOr
onLpbDPB5JWqXHFnFFpqrKHjBFTrWf4AYbkDYMPL3R7vBVSrAkZiv7i0wfC3t8kT
yLhMQUc0fgrSTlnrhWO4X9vYcFXQqBI6QOHeUX0QCWGK/SBT2x7/0vXMVgsTsSXX
TgufRNR2SsL5IVrZ5G+HNdSaBmJ5jd9AQu05PWIE/n8=
`protect END_PROTECTED
