`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
prF87gysDACOEPQRuMnfB1g9cyxDir0XtewVaS4jVAYBHe+oXPwY4PMJ1sDo+HUt
9iAZmhQeTDUdx7PmzFlSkgJPRGS8oXxmGqAkJEVT1iYtITD2g/zfS66VrAWmlKID
6d9gHpsDKUdzx3LARN+yE2z9NhYReQg3bXaQ0E09TsjKMjdwTDMVGhJZVW1OCzRN
xyAnMAxswajwS7mUNQOO3tNNDodIr/Lwci7dCl7LdK2QA7K6whi/blxbm8hAxM2F
XcXAp9EOWiDRnVhpMz/Om3B5MYqOf52waG6sWk5aoDEFABinDVgtxt36bRI8MBss
0ilAr0d/3+t2bc2k0jzgaLsTi7jZCBMTO2j/hexn6BbDAsOOC7Ct41u23WyfraHG
4we/Rlz14eXw1SjaJ8Xd3Tz7E2t+4zCsm8TUa5KiOplqwN/5fj63hmg56qjVg2hf
K5R3/w8v9OP1QV0mTPeEocIxE5ywyU4KAzDBMfYsK5R0zSN1LEkixDuAcG/t5cKk
Gkxpt2v77gY8EVdGiI7/HZM6pmRTzWRNquH7HD1A2oiKdWuDMKqSWzvSnVor3bOh
KwdUK3zLWVV5UqRxVFeAow==
`protect END_PROTECTED
