`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRgCNoMeTnzoKfa907EElJ3vT/9CzktWbZfKPC0Qm4bhy1CwxXFJn1sMzpQOmwjN
INrDTR3fpB6mEyNyGGh7qQ8Lr/rQmlxrfNvDUq1RBjaYI8yIon5kkr3YTNzKAvFZ
b82vI1mj5HX+tFl6SammgW/ZjWH+sVpEl/2jvT0w2kJ5A+emsjwRgvwY59ELdplp
vHTrg5KWPlRtbiDgBVYHZlR+yMx28LlskKdYom1uZxyeGAHUcR2WFKCaKEzuxbny
1HhXN3B5D8cSrqFhlBUUnf8PTAlFxlHOGS0hWvPtKMIntbbaS6/fNd5YhBdSGuWD
xC/wLdIDj44+KXqZTTjZ7k2p7zQES7cQLTXMtDzgWNHqNnXpX0AmxdleX33zukDK
xrs1EFQkUCLXCiqkQdFKMWANAtNQncbB8UWFMVi0A5TFKB5EL5CH9WGuY4GrTmm1
kuzNbtZbuC1ML+KGef4AkwBUlAmQ+Yd4mZZ2gJ+Ff9Bps8tCNwS+qmyeWL0m1osX
ZuUAy5n0EDi79ZvZ5ZUgbbB1fx/7aR5Qsimlp4CpN59y1AiJnoFt8Z9rYSZyc202
oy63e9OqtmAJdHNPlwqcdQ==
`protect END_PROTECTED
