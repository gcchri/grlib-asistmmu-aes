`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qu0ys6O9aYJH/isKAndOZKV7QU1m+CvUe1o5zSvYgU0I3I80ZppVwajgTT1znZzJ
n/7KoZG0mZvppGj6JcLN2X6Vh6pnXPapCBLVdUqY59+B6wIhoNH4EMqHa4Bf7f4C
OJpi+VseBl85D3jaY9Pb1mfhW4EQqRFkAmCOgYSqEwM+0ynqqJ2C6In1FQw2KuRK
Y3mUrDS5q2TNKQR1qTsrRMrnrvu7ul1RrOc7dfUHRdEudY0yP34FKliPgB8Uq7wN
O8vVYOxmK30vYjBL/pLsGrKFgaOWcsHndgb9PDP4nMG67aBk0VPz0jmlAyhZAGR5
5l3C5SuvL+4Oa+OitXa3bjRH0exxPfVEoAkYxyxYdlE/tvHIWP5Pw0lhBV5wQH15
+sNjgHu26k+SnCUjfy8Kq2T2gSCqXqCFg/bWtE4RpACY1FMKE0st0Uh05uLB1+qo
eVW01k3TjZegL0fjuBHXjHPtdfqDYUTxIDA7iQ+zqC05N9zUZGkqo5fg+6DmlIq/
qF6gnCNfsrF2fMDp5RxVoyhJEcCyoZJuQuw41lPgc2spKwYzkrvkQlsUqqnyT7PG
ry/27Uuo1Jtx+5QCE9aRUD1I0/wCkjm5xKPIas1DMauG5b2c1xU/aBoXfDAnPjug
M59KX6ouxRccu6rfcNFnoIad7nefLQGRcBNda0C5UgxuaS+fGE169NTnmwZdOhaX
`protect END_PROTECTED
