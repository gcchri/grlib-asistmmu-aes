`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZobSLiZj2Em3xfZpDCjh9OP5AOlpwSifcOb/njMCbPVqdjkcxCwxVyzARZxSGLx6
FfYFiitJn20NSGzx+UejrA0dBT93mmkQG8UmSaelHt4x/0NxzGWa1W27Zv86Hmec
YYCXHIjmG1BYQ9bVUpeJ2mDcCGSz/6oGK0IgU/SbLu3YN3zU4XJBkmFJLGLbZx6z
6gGcRy7Z/II0FW4mZiCC/UHajzPdSdmNlBlGjNmZIeqwfquuAwQbZUvsiQ0YheEG
Ok+2XOMF6we3h49vPK5UANImL4bgaRdXkINI02TOsEtC2OewhXYewbgzNjIRpg42
iz6Xruba0KpnPUzQtzM9vE65RR7njw35Xgf013F6doHI1H3Kp52nSiaaXFKmjrR3
OG57EFpuCnuiFC4M5+4aGhP25s+SslZxfPDRMaXVm3bFrPOTHBryIquzxsN/0PzT
AHFHpMTX38w5j6/NjrTQNiypeTg8/u7Xk6PddMRkSd5D0/aeBJTKaKB5njefZa1u
8kMVxglW+fmCeXcEA5h2zidAIGLUOdIbUNZn09vo8xOmHzCKAOqsxivonvRyM6gq
ww5gRqLzVmzaUz7ErPI0DxvtcNq+k+wgNBI+ZqqxCybX6FnycJNemMzr6dgpZiYm
9d2lk1QPVRbT1TrM+Dy5D/O2wktRQKe6dZ2eiqGDrcKN06ML5hWz6gil/b4BR6xo
jF5IWBH8zE3CATm0JA35VcJOB/gAdCeIYkONvA0SbsjmCB35/mNzG9C3QrLnXyb2
fmBu1DF9Zp4D1t5yh+E5//Y6tzQuZPxsBkYCfROtS20dLFPFrTX0t39NIlJkUGez
L403fGx+hH95t/s/N6QZyccId8tvVgCJ3qBCTo8Z9MX7JyhZMPDpaLDt3y5mPkZ6
RK7VhGIY9ppjg2qsK57nHD8MBo3U38xz1yyF+YkgF8n3VasoDMZC9mwj7aMUH0+b
`protect END_PROTECTED
