`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CmLsC9IryQkdaTflNwCVkSoE7ZwVd1V03C/peaufqqEiJ2VVj2wC6JpukLTs+xxA
dK7ri3heSehZjLZReq5PNo+ZjeAPx5YRbapPXj0JQwMOdlJEVZDq+fPuxOgMpesk
VgvZgZeo1waiBkrl3pq4cud7UmPIQw+fNDfqThR4kPoGcLXsl5S1THas4eO1mRZj
DlFnPILlzaiKuUoh5F5IAk5M1uidI0VsWNgDujWVXhg4AKVggzVHPlg9iY5Aptlz
b1eSZmVlMAZAX92ockP20HSKnF6QknWZRyAHq070hVz4sMbnW64N682uFXipueAx
l8PeHGb4r7ozUb3jnXPV9QHeT3cUaf4lakdXktBhSQBC+YhmBPGXbsDX5btPeeOw
XN22VDsZ7WG1P/AAWYXsBWSm9JuXohXYAHeEtKK0Fn6a+s3GBc6npLNxZ/k+VOgC
dtKaDlr68DhaqXf8CMXs8eeB6gsPryQU5QZN8DNOso3iqTj+VmVD7+JuX+iaN7k3
oJgNYDJGIMNy7jVFuak8VpWoG+yqeerCQyfBvM5R9y0GlN+jNTYpjPDiCjpriPo6
3WNkt/itJXf/u5chQp/z3BcHtP/E4AQCCbowuW8Wekp/xmeLra3ge+jFveF/HJtF
KWcbJC9XPwhqGO3g0aybxg==
`protect END_PROTECTED
