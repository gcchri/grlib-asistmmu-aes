`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/g2hVNOSy93xUTW1MzzerI5qLGM6e5K/6BCdxEwg8YFnUf6rQPD2zTzz5NbNUIl
NrlVH7xkRNzeg0lbglS/eKI6NS3s0p3YkIlLzdMdSjADpDwNIOE6sqGMAcYutmLJ
RbVSCY0Xq6ITSLe8sDUk9T8ReyFcMwyvu8IlfiKMntzDvpY1W1eIv8qp7I+rU20e
XJEC1xA1lScZx8axIkwMEBMgYbqAqhZZCSLWLuDz6bH60TnLoZqpsTDpkY3f7Mte
GkY+KNmZ7qv/SjZuyCGR9m403p/kMNtqo1DXmk05cZKAvRFTD/dk3ZnHVaP3TQuX
ULIg9mQ9xnKcjF4OVti3Xg==
`protect END_PROTECTED
