`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8h7lrlf76rYH5w8GdpA67OERaZTANFfruDg4SP2Gnvz8T2aV3o7NNx/NfC12obPK
r/JntA6KRK1WnHjKl7A54iL0ejXIIH9m6EqALdyM8s+pYupoYyKsf8sP4hVIiGKK
RSqHqSbLA4XraNPSutjMJbwgMqcgcvJKnXRo4iQBlq5bA1MSIzEE50EW4fUL6Oez
koXBBrQch/5oBHryr1BYuncghox5fki5RyTAERUg1Ooc2aDwBbpPaxbg5NAgbnUB
D9N3dkIYJExVStLdaQipgsJWyPdk9qaaN6oxSnK7MhJBYTPHpwEJiPp8vjRrSruQ
pvsAme7AOTghajjL5sOiZg==
`protect END_PROTECTED
