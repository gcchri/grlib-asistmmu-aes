`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdpWvxyi7kMelIHRamg29GqSHdcsXgMh4lmNmDezIReMCHtEQCYNtoz5i7t8BCTS
GrKKi9v0T0CrYq+z1uNN8Zv5HRzXadEgZOiMddylzIQrdwTkpr5aXvgyPSoUZDdm
h6ES/LZyfkTzZb2LaOuNDv8AcB+05v0vy9YH6Cbmwp8DoBgISNy1Odh84emXXej+
uC4zAxqnzeFYKjDsi7MdMVkLtoJzH81yM/7xAs0gt9TPyfwMXuRknKsqn97rX0Z/
G07xpUzkIEReQWEOBrNPdPgOMDfqXiawZP1AdYex/zM=
`protect END_PROTECTED
