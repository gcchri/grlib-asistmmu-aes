`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/AK6l405S2L7/G2nU+ss1OEj+rpCmZMgyEFNtgG5gzXJSz75AeWadqVz+Ny911p
mkrdCZ+l+e3MKXDcWDsKgpjzt5XeUJdywZqjzOlgCLVwfLdbgUs1F28p1tr+yDXF
S1JO4/+p9bd3BNYQnl38fw5Sj6OoogYO6NbbKDA0GA1Xz3XFeSTjwBFXE+HxtueZ
H4hMgd8Q6DoXlnBX6Jho76GuTRD44OMEaJLwgTOFIjM+Cv6vnGA6K1RboNAMCExG
49biYjFxD4r+nYVl9qd8j+HEwLX9uUY8FYDrmMUrl+np9rY5yUTkTxOopRxBs9PL
KW9mdqlf7yJf16pT8omF1IDup3fSx2dlarwUXEDNL6zeKXYh/0IRj+XzUKBamB3i
YmdCA5gC0ffAu6w1uxgpM4x51+F8i7p7dsCHhQJSUmoXqYIB9ZXK4ehhW1PTmy/J
gD2kRTa3ALGtPBhIm3NycbPx2+vIwY4aDQCmICYWIuuYjeLjR/dluLIJnSwasIkQ
X0py20l39wc9fzp8wpAQ1AjgOYo1bXoSpsrK8U2xZz6iOUEZV7X+m3PdM4vZb6Gf
Z+I/oBoX0Sju3ytZqL7qkcBtQqrtm1C9TmvfyoBhNAzl5U097eqamRuGdSngiDg7
zBK1xrG5OSvS2fWDzynUmKS6ReNiO39aYHBNgLNXWVl9NbopDG1V8xMZg15ywbhL
M4ode4R2GGoDnGUkrcWXZi89JmATJeOKu85JKN55bmLiIQ63sp04KTZdeFZXQTD2
Jeg4TwkSCBmgj10GYquERDzorN3QmHpXYXM1CJs+Pjll8/AaOb+RbuZEkWwI9SrD
JcTy6hE2ZusC3dBSOrd2hAhhlbR0ZPGwair/S5vCvIJXm+brOlAUuWZXLtXqGXcc
QkDKN8mBzhSvTr4h5cEIuNdbBEpl79nIjeI5FzKGozK0y/ThqjoaCE8e37/lq3NG
D+ol+PwqvOb8vOJG1sUrIcKXV690JSU6FvDMqHpqtgT3zBgYKlF5JbcZKkTH/4Pn
DWaeaPbaKsrDjW/XzXTx2PHC4IbDdK0gGMKahMkQOcazFFz1QZvMB6XD/1itxa88
UAqMEgU8wo+obWilbEKL12D2L1OJe+1KmWd6rrbEVMRgk8M/y4GAgG+1TjW7rPFB
wMM7KyO73BYqnVfQafuDGiDAPIkrrw8Er8QK0AoQUMcXFlBoP7ukMFtUuzU+55/t
rs1Tk8imYXYpqh5L6XMI9DzN4l+IrfDR5a/eT0YeD8EB/AeCWWji/5l6g09fwtey
HWv0Uw5NDmz/hPMybGl87N210eNc5pjcAPH9w0le25gBNMrzkPvGTdBoqR4XeNH3
iJ8WV9nGLbJ07t1nP97RtAf2TITNujhU3iEPNZycmTFPj3cCj1If4F13JvYv6SZk
6MVnE1bipNDGKP1KaTy6KY1MWa3CZpdlxwhpjmlWS+zJoc2UGmIvQZTjtXPQuzcC
Ijhcb8pqo+N94V3eeopsK9cyP8/jaFINx4MOkAV85e8va8xZUx1EPeR6Sl2A0TE3
s1lUr6jW5LpYxW+C4VkhuR7glgfs1DUk8bNlx+JzSIepOIa/ukt8cEHei26t62RQ
IkXKRUDBNpL4UklbdnHKAX8weme4xMql+tjgG9D+aw6JO1QdofFDZoq1orHt5eEn
J6ZxVME3HPImX/NtJZfjtsUeCYqZgxJnJAb7CjabwolXiLU5EoVqtGSUnOJ06zPE
3jRtmfR6pLc5YfX0z6S5JlSZuyixoOrFBS8v9sO3w96LgkMiK2JoLFbb8VlR3Njv
xpProBb6sAsU+JhYxJ0IUxV9ExyCbFjPqptwEDRgbMe345QALAHGtT3d6Y6VWKMe
`protect END_PROTECTED
