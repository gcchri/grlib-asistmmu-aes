`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XL/GK/kwEDkRRaAW1YYAMj2SyUrmiqtp+4Ezqw2w6Bos0WENasATgJs4/W6Q/9ad
XDg+ACcACub8k5r0aRtDXF31NHpUg+4opvA7zVUYQxH93iLv0YzBrL71gnEphyFJ
AHCVt8MAZsPtNtk78TP3+3kz07wZVqXYgQJx/4yXKOxs07SY1uHnKFdS9yWoDCi5
HcUFx6CwaYoQJVugyQurJiiLIW54+XIGpr51SiAlPDIchxaVYHawUP909C7faxIr
ytXWUiH1PlbyNF/Ih+IwCA==
`protect END_PROTECTED
