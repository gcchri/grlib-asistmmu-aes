`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9JR3h8OkAlMCdfDeyTTvesJGvCv9VgoGXLxhJgleAvzph9pajBfwPho3Nd/6Wiq
NdBZVJ2DrmDiR16xQvPb3S3hsxOZcR+PjVCRWC7g1zh/aKOOh8e1M1eIN9SSK4qQ
iDhXfCnzpcotZmFr3180VG9IITu/jJmNbreS8uiHUs9/CN4SnpUB4aE/xdrkyQsl
ThcFUojL4MDjCPlkncENlZuNomASFRIjmqreyPzRBIycfrN1Fievk+auglA/heme
OrcnFOM4WiMpSQbVQltQgUqjU47r82bVeoGKH13oDxO68jK43sle31C6LLpu+L8x
1V1fGq3xsventowkw4yd1BC1JdPOSeiVu7Za61UNyHNexuSgXV6lgImuSQAQED/q
KOL9mQ1kaUWwIa1ikNNULQzva0VN/qBrgmcb7dyQh2zMSzvUlzIEZQx5vcL1t/pX
IA6Vykr/zRhZBwYRTXuATx0swYfuGuw4o8G/pLwb9eE8B3lRLxFcw435yYPnNMs/
TjXV8ZRShEHq2LM3KU3BIq0HX0lKN8RsCHflNBuaJfHIkPyVz+rQrZQokZoBy+aa
TOIhjIXyKZ/+MAkw0IDM/f9CEqqrbbnPqE9WBMk1mHX3D4tTzmNzcyj/1gEtz3KQ
rbtj2T7QViJJB0EVA08t4FOX2UUw6rjY0zzO9f4KPL1tcxvhPTHuXDoQTGC/tOwv
Ctid2eQba9/lhsJntGyS6cq+jbfL/Y/lnEugs2DvqTNeJvSMikkaRqWrGjyN7iic
UNaJFwlTza7pgzr6GzEVRnfZeKzHvhwUvbgtuRhm5NX5dGYWBrZltMfH+Hf/ba14
ugJHhpTurbaIiTAgbzGwcPAPMEv3NMa8hOQYi/5oDI4gFb0YIrunIQTcjGxUiZFn
RTC/Ry1DeTiMWYEXjp65ooeWVjNhkjX0zsMPL/wJxl8g5lBvJZ9MOCGmHsGCzIB0
tWUO8kj+vr9lht1J5/29Tw==
`protect END_PROTECTED
