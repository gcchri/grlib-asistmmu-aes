`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GVGh2W52hNOJWHXcpr77Mz0UgLRJ6S45dayL4UAgDTc3StYDkkvPaN3lmTGMDk9v
7LCuqZ8yRlikmZINltNovYVYH25fd2VlEK5O874u3ysK8nEMGuE1DYAVcX31UZXg
9sCs7t+B7l6Y5c0STz37DU/9M/u4zutqtMu59brk0t3ls4fzNL1/Dd0HwxitGhH+
yJpKRUDf4qEPo5wN7in/rgk4SldKiosh7zSZLDtEabfEmEbTh18dhDnz9fwGPRIj
b0q9vVrVExaL59P7eJISKN5f6zaoGpW+3KEb8XBKQeXwJYG/em4UrRSLs9jSyqea
Pvttn6TZoh/VJFgWBvmU4Js6K/AfVfrJAtiV5d0Nd2i/IuyM9+4V1CYkMfvYDvAB
ttMz51s/S9QEq9joId3FvrriJn4nEJQcm1PzTTbpNuga4OYNlIrmNfzA845XZnQJ
n6xlM23whFm08LV7KaEvdIKPBQAcL42HWXvmbpDX4ms1Gw0phgbT+EnX1Tt+COxx
TWuulJmx5A+SnOOqCv/+zQ==
`protect END_PROTECTED
