`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qzfvJfLnxpVXYlq+A4lzS0LLrus/f/7KQOUsIujP9LG+gIwKaJtMJs1M/v7eS71d
9nSLYq4gX3iY2A4xvyxAJg21pJqiAw1vsssny/pRD/o91VucB9ODFcccE9UL3Knp
ajq8KKNw/t9DVMSslzdRDHttkOhszXSqGeyqT3qpugDaOkqoQtXtjKDYHLHDGP/9
idOgfJ5dmpUDtz6l1nmvMNt9chmbG8dIsqzEQ4MZfwHFue+I6wAHdN5GA3n+1ltN
0KGBzfhYCA6D+hIwx5GZL4nYSTfbym0vKFiGbmlQ+QNrlrT35pn9wvaRJyLNGmhH
PjrMbWfcNnoXcguuSKa2C8wsDiRlyFTWkBsEYT5LxkPp+/Mneb1O25BoQDZSESPB
glok5gr5S1oOk38nH9iKnBpyaorag7armX5DvN8kaNY=
`protect END_PROTECTED
