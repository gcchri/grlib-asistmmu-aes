`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QI7odRG2VpD+m2c0jjmRDBBjJx4bulwLrNH66BD2eLWdRkXYMYgIVYbp8DvZZq7B
meqBI9L9Mh8A8xtngdHlueZ6bOswGgPEKxQn3cAtDYV8Ezkq5jnZk/C/4EAFp9WL
AQ5VKGeTT/B1QuUbppSa74qZ3hYpBU8ARKDq+JNoA3ivANgQqhSzViaJiAXdVyEz
cXnNnvbw2G6ftpdMueJoiJen/6cOJrWTno5AtEe7mNPeek5WuKfUgCthsDFkOm0Z
y1XJ89YaJdJ8+cfVnDklpA==
`protect END_PROTECTED
