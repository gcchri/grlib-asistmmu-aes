`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1PI8O2vdPB/QMcucquUEZfZhbeTQhC1LXkMmVNdzsUSvUdBQUzgjVfbues8nW9/
oFrzrHIbLWoMZYYJUBmgPM2h67LC/zTFkL4fxiqW1tBvJcseCnMKMSprc4iwp8AX
KSXeRKIa//5GHp+zbNbkHuUxKA74odL7J3IVUDmY26Ay66fOb+8rkQCNt1cL/vqr
FOz4vgH/5RtU6/fBay0vP8ib3KyRejFxVsllDpHSGFj42P67igA7urCapmpz92Yk
oi8B0YaNIX+f5geUjSk+ijhDO5rvuq5cebB+pcDrdTm5zfzAiNEiVOoCuH4757yV
BfyLYW/sqGNEh/SK8d5oD6HdOBWRzMn74Gl0jP30iOsWiCQ+XzVslXxvczYxaIE6
jijEAqO9GPe6Er9b4lWtlQ==
`protect END_PROTECTED
