`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wh7PG6J8XmVKF/LSQYdt52BQwH/JDOcz+pDPg5L70//b8tU62TMG04OnnqMDWdwK
VMP2urZo+fmlWbW2PEZeQqIse0puwvSMa/c59E170Q9V+yT/4Qmi499W+zyU7hxC
IKT9+FshyxW3ETgnmKVwuiufmjQPlk6xCJREZz3GtL0iAMvxxq973pmPan35VY6E
HL3OaqSR9w5Udslt8PpfP8doZIUhSw8QSxpS+Du2oFi559yOHZV7bvpzXjMAi2/T
bcGignIYlGfE6JODnCy09MCp5rEl/xXd+SYLZgCdeRHxLzUvtNT2tj61weocU08u
tQT6Z5a+8qU7JzaKLmcq7S2VoyGCWqNWegbU5qSfTGtdHHMY/YQOVjK8ViDoGglj
1gK7dmZm2KANdHgwtoItDW/Dg0cQAAU8qxElwydlVFypyMaUJQ6vBIc2awFiJikP
D/t8rdsr581ur8bA00TGpQ==
`protect END_PROTECTED
