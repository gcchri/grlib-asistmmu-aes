`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C007A0SW8x4dJZNYNX/bumgFTnLqJ742YCaRvZAOPXkyNonPCqberwPPJ3k7FIFI
01HjZaRaXbCbj3KBbKeXNR7YWskAYNyWniLyRbYBL5+R/SnuUt4E42dRQ24ViQic
wfM5dN5Fv6DE4mW4Z+x0Bql753uSdziW9MpCYhZ8h5H/w9oW5vZLNFa24yr/kmux
Pax4zkUMfcglUfOiqAi36jBjxGamXfG2rImxIc0xH1OeYTcrK/SPoapsc0VcaKey
hiUT0/1XWWxQLIKCz3m6LxrrwH6eYndl5dtBCwyJ3fBY7cKOa9Mzins482333JTn
YbSp9JLgCV6VEiiJ38CqhnnPa0BVa2TC8he/dIJOUm79KxCurP3aP2NvTMYOs02K
4y/IltEJt9NwP0mrCSVNnMthARzACHuRbnsTu25k65rRQfR6Zy+4YjhVdC4+sVQ8
i+B8W/kCb9xSKNoenertwBNQzeo8H61vCTapzg8mK3/kSLsdk3S4sEK+m35T30sa
0fs2NMxh47xzmCouULAKQVnJka24a1/kMUZ+q9zfZPhG8+sHJ9HncFFJdlINXRRE
L8mUpA5Bf1Go2tSNnjHjtwQMmHrl/PaS/Cw4IiqeB16ili96r3IyDR4s81Qtev3/
dzoPqMf2E5n+vY4CmpKKOM6u/MbcjwdVZK5f0tdi3MnaV4zRGgFG+afgvVRtj2WC
Xq/5l7N8mvkWVmxP0xBPeTWIGvAoP72ClX3rhqZvr62DdiHp852Iwj3UNMC2h6Ii
ktjKPyaFQcFmJCPZ7isw0u1KyO1Lo9NVCjKleFFkyFMqbE5Wy1VC6DZ2lfYYq3jQ
D9ZZ9it3c/8NLKgC8xQixg==
`protect END_PROTECTED
