`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxjQgdSSnXXuYs/+J7fKxR2W4pf5VtVwliOENo2Kj3jZoopSMA1isypclab+vJ1u
DSPMaj3tdYQNjv60PhaVYTJfZu9jzma/1uKRgp0+T2FFmQvq5rAFrqMRfVyXayGC
cHvdYXx7DSaDLbv+TigP4YRoVAtToacnmj4ez9OV/fkcZ+s+uUHRheRp2qHkL2lH
PlREWru8PatwtnOwaNqMYaLDTA3Zlv96hx5qAtQDJp3LOHJBHeGyZPcYmmk05lTz
MuSpuy8x/n80LnuYhp5eMbdRtAYybp9rQE72OYy+W1Lpb29eo5lgAkrnYyy8cs/F
J7ycxU6XWmooincl2FoXlPlAL/kpCdjkEs6gdjEViAkhVdbWhVv6nCrTLl3GNsv6
tWeuBx7nKBNqKFWfPzA5iVRZtTw6kgQbe02QzXoR8uyJdajNBe9AuuSHnH/DPrn2
3Mk9w83W8sdenyOXSfRC01SemhrehQEaH61Lhmi4PYew6KnSogvUUI20hEzRXQjK
zCV7xWcmFPyxJUh7pt02f9YgVP4VIoXlkl7V3cU/LOV3sXqLo5MhyBy2iaqCRESL
wJ6bnfVAVeHVCbBJ8cE7ypSQcPIidTVJIDFytp051LFAE5B+CHEk/pw42XS7H5dV
ohlHicbpFnEOHTobAjPotUreMh6FURXRcIlvNRyGYcKVwC4HOt9gERsNAeFcLi3Y
OIzjuT193sYUhfmZ059XlxULO2Kyy4Nr1zxI6DXLLBJzTTyEZBZTDRiXEmEj8JqL
NRGARlNHrVN3rgczQwYxQVFx+RZYA7p/YXr0pqNTUY/KmXvkK3pkpZzRAyaHGO+B
kmh5pAr7GKZhUmlafL2BrqDzknwVDzrb/EnwfrogJEIlKm4bNEqNqzaD2fvieBii
4eyuFMKCgz/g/890MdPs8hz7mXtFIQw4owCYKcd33dekcnRJqqFTNxzr2Z/kIpxA
d7ujlgUWV/PasmpygL0gEaKcj5ME4G+cr/6mINtr9swFVuhLqFBVJG1k8jUDu281
zuuyMNVfD0vrRmlyAnz5cK1LpgLZBu77Or9ByecDIbwwfw/ADABmXtEV/txr1v7v
HYZXIdF+Q7i5CYsK/KTrelN8ZFb5sPfxw5ssZC29sUF+r65JCT/eZu9OCRze/UJe
4emR1X7m2d624ibNZxcz7skaoaxtJ74FiP9IIvoQyu1CCOteGG3t0p7nNRW6OL3z
6cE4stacwFJMfpFxwo36MAbpUILgnIAiProYiTP50ICMMEiqLv5hblhaf0P4kyMi
xisg9+eq/PpppHc3xRitiDeoVaQ14j7NwbPpOfei/CCkqVW/4qTRmb0JZUQ78WSb
67jn8tUqgQsvLaHwBnEFT4gjZFcuSGVoFHG/OvF/cELogsXVnsYxgvF/Ja5XQzvo
vo3rPsXjdhhtt/neO0xaLu9kDjYVN/DxtzA7yzGNDoYpGQmQf1Bwu2Jt+sDrmSIZ
L3MGj0/AT8gLOMGQhLFhzlfeS9Wf7s3cfbOq1VyeMMXeTEAmeXBkyKb6JEIJWMxs
ql6WhPVE6VeMXqifVeSwx1Y/euFyrSfx1GU1p4g7thMx82Ck6yl801uDi604+5AQ
uGqeocMkxks/6/mQk7tSdVW2WkZJRA7IXtvN5aWZv0yV0nkbe6TJ4FF5SP5Ty9oH
mMoVkd5sDZ35PYJJBCMHYaO1DjrdiVqyYJ+z6BXQ12w8MKoOA78T7agcDiwlIQYL
s0hQJweZD11U0en+c+LpN/HLqc8Z6TgF/HgpqNz9TLwkxSlHKS8LstL1ciOBINb4
6v7v4Fzm41Si1NkK4aKwKiJd5lTMyqEax3PpuSR1V0vbRjdzca6QiBMebqd7YOfv
c0wY7obeeMK672oFk9CADDnRh6QspGjRYUasqecJs/KQoGxVPSP+/53fTQjJPNXB
`protect END_PROTECTED
