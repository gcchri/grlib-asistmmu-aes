`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k4RtUPs8h91B69I+W86JoeFK7PtVI2mgQYoyoGGmh2qgMiFsItjqqIfXbXpowm7s
eLHv0Ube8+T4qEzYnLfEh4ZZSfwH9nuPahjVf/9QgQHXTyxV92Jor3s9r/45RbB/
c/JioTgvK+ws3I57OHeBuk6ap5BKxWh/J4IqgodFbe/ND4551du1Dmv162ENbujp
LD/+pUSYcPC85ZEsYFIX4BaPwkAIh+Py1SV/t5Y18pDHie81zcl7IDF+3bXAsEIH
iNYawAopWfZ+JrGhbru6BcP+UhnRbnjZyHAtsM8MhZWbMFr19LcvCwEddx1FMukz
TWl4//DUuwbJQHcKijxVXey8g7qE357IRICD4y1/49oATy7mGFCiqTjx53MfN8R5
M51D/FZMufONdbzexIl0iPTdTGcBbC0q8TsmaEvFny53//wZB0kkn9+0aU4LZqx6
nsvjQpKzDfdZFAHNuc4wRJP8o5Oi+lfhw3Q78L7Mb8XeC2XR4PbGLP0BkC88PVoS
7g34SEQ5yzt2oYOZaIG5tNaYZ4C34O3W/TceMcS7KTElXQGXMB4p8M4QJ2RzxT8v
W7rLiMkDTOels18uo2PAQAMpXfm5wgtWC3M5D+mnc5VgGoshJ3evSBXSHwSHml4R
9Pi4YDDBdj42oWmLzu7CTQ==
`protect END_PROTECTED
