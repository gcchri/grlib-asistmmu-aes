`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEl1RefCSyMR9IaIEYgNJNUet1DbhANiFWCSiZintuQq8RdU/3hAOXS3z74GT2WK
DIZT1n4Y9gXI3/YJK4Nxv3AFotBH/c1jqIaSMUbaR+uHR/f6wm4XaN+xJcqSthei
TJsBVG2eHS9K85yh/gqrF99Ub5hCB0GV2My1+Mh++X1ghq8O7W+qFtCZcldweTvA
9G+SPNjbvjYh1iNnyZ8SRdc8mLVvwAXbbSLXJfuVdf9gUiK7E4HmybRI/xnsrBGK
hfclC8N+qT/Sm4loA6Jo6VYfupjm91qnovyH+qfAv+hu8DollUSRfa6/fvUpBK1M
2aBLc2e4OcqUUeWrg8jdv61Cbi7/GGmFBUn3GqffhSCT87scXBnWNrAL5bpS4+2f
qn8MMEdVDQg2ApeE+I4bW80OhKT6sPNE7VmYeQUcdeLD6GtOxMrBTdM+SnCZrveP
qz50DzLAA1+wCXTUHpqVrCF8jd75zoZiZmhkgkDp/oU0GT3xzCpBOKqDrDLnKbvU
aETuuE+1zxsp6PPkbBbHBP8l4rw7p4L6i4ncSLE6h1RqLgtRsiD0sJerVoKltZrj
QAx7kd2fY39jiLwT4WYQjQ==
`protect END_PROTECTED
