`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gANirETThmxJArZbBr5pm1dj5tLg52Vf5Ibl+W+pb4YsRjTTelmdHpP01S7vkF/
z49AdDoX6l1H7k5/x031aRV7WvJkRR/NmRdR3KloZKWVd/+FoEiAcg1YfJPUDI+1
4I8AVqYU5JgvzsJabzO03v58olGYjK0LDGAjfXT3nQuH0HxXzPQWQ7G5qFt5EUX4
i1vnZVw3NwlLXiVbBecPqsL+Uaocsa6mvH6WYst9/alG5qevyKi2HeksY8nkFojL
EzaM/Z61boxGxw8Dw9Yf5cSWhgGfn39/5048tnkKGMWdboh2elu0aeqD+5ZphGeY
zl1sjB7x3vSBOn32a3HJ1YHI9owgTztTMrmvnpFe3oiZOR+16hAGCusYeT8MwoXt
SVedW6MUshnHp03FqG/LCVx/DDx+9X//V15HcicswwEQnSUQSJOmIbkUN4/ICHXK
nAdmRi+jzLG0HnCdjT45dOh6Rk1au2iOdxm6CtKOXriGOVQrDFawg1FIZGDngkzv
zoB2ofRQtY90xKs7R6wn6Vz4ychRb18gBiuefqExh9cfOM+wFLJ26e8aD8pTykVP
TUoXkODtq5mcGEBxNuDGuQ==
`protect END_PROTECTED
