`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
agpzfLC//HzT3uSHLPPTTvykM9+7+O2vk8fiHiEEFSw7RSW3Q35nzI4NIvC8ZLRp
FDNqabrr3con/K7fBBtQ26Kqtc2UADpdbmYlJrqjSr7C8ayyOYgNLhm23HSe6RWV
zA+TyRxcZJBfgcAdmIxgIuo6+liu+Jn8tEk3Xr++Vc9977C/kLF9ICYdLhsn38kS
cxX7zC+nxCZzs2xs7F7ndlr85rsygZjOnCVhY3nO53Q7pRdwAv5RTQsMy3c7P31A
QN5bdf79rObRmqo14IvNO2u4DHzWdA/T0dgDl/mCu071lOa5UMnUBu9BGw2EbAeo
Rk0xWgdwabokVUDCKryHD3jY7YiZ8WqOUupQWEU6dDb4Yxo9AtiCWkTfFAE9YzFc
Xbr0tXK7LL+XPu/GFjn0dRJwwjUaEbHz0WW1QMNEgHAAkK3K0h5js7Xs28qHlY/a
bk57mh/iSzfHxhKdekmyFqo+wz6SxU9DtxSGRDhrUzgKFP9tV8tcbbyTXePCJJGE
IFod2wl+5IpPJkdthq09AlOFDwo7iMxMfhFEIo47iR8H4Q2GK4G/LLEUBEGsv5A+
N3rnis0wGGOgmGA3ld3q4BvuqzbhfaXRCkASUDu24y/isrAs4pmN4aQjlcg0ciZL
6N4Lkt3KB7WcAHBHADUvywmK/6VxMkoL2QcXLmgqHLw95p1WIa48CIvQeVBBcBh7
wnr/f5yFk3WauTMzxPoI5ZvY9+NENgARvyYfLVduLmAXV3G7jZq1pwRq56M7DOMz
yhGyVece0KA0wZlc+BP9+N4CBAn9Yt8/8t6i9jw0CentrYVsga0G/9FAzJvpIyHi
nMrnZwIlg2Bnm+eDg5HzWD57/VMPgun77N+bDUrpO1k0AYJRt+s74KS97Yea1S/h
Bu1Dv5t6eGKNB68B1o0lrnkLa810Y57tMC1aHlS0rXkKbr2I3fuAACq+1hNtGuSU
vFk80A6JnprRE5JVjAYse/Ztre0kFFGVUFbfVlMlSx6OXetxiR1Vbfj5HBLD8RRv
rsQc96hpOKtXyFkDwFMbZFqzmuc0VL+q+Cqbc2ET8WWJNhiQPKDndCcyNfKyV+Js
joZ7XGdegt3qgpZkuIlX2p6SOq2cJ9X0Z7mMvm4x0+AmV8zLgy93cduTuhepWH6a
C7R7vLbj8z4xrZYD8M6c5EUa+OsHWJzKqc3eqUjc5eEByQ0GNjNSYsmf+Pik9YTo
zFrFo0o011ExctHA9dr5Qzf7y1zZoX7gvC/0jb4REMWvAmxTLkkTgWX1WUFRdIIj
W62Uh/4g9V3gIBdq+F7y/uoKG5QBuM/jovREMAVBwfAhYfEA9MFv34FWmSt9JB6p
U2ORnBPIbtKefR4u4Ua35AtyRQ8e3Pf6exirNrWppIR4cggG0qwbUWSAEQNil5TM
Lw+1CERWku09djE2DoYBixznXNVuJZH1Hp13vSQ7xrWSi84S7KRG14TY7+RehQLe
WnCa4/L7MQRb+82ri35ceGE4mimXIU6HTSlGz3bsGbQ9D6sKDuDwVGHn8k0XO+Mc
00OYU3GVdxAWMq5whCNF+kfWw4RGFypbA1tMEbEPF2dctQYz+n/i0rjM8XGF7xdO
CcWToBhzfDcEtE1Dbv6nuAKjhfHUTg7+UIoiRkhscVq1Ed0geA7E0csVcybJLAlv
JF14VYc3XMh/6GZsyY7LVoqs3qaKlmDoldHlmS/did7qH8YHoBgAiCe4uhZpVO9c
u9Tx0HnQ9IvKIEbz1/r2EhxOWxan5KY7Tb/UTVgzM8rWMw58M4tJn7YjUCVLeFvy
zvY4eRqbNBRwR1zViTQsusZJxV0ShnPxb3b4N1m10a1e0whDtInB33O+qkUTn4a0
GI91hTZOBbOTSYfdRpfIBv7Gh4/HoeDvjA/U8d/jTFZ7lO08i9j7HZd/hM1JEhkU
YMuB0uMNvZiF0GA3TRbOZHzqNPdqrwIZiOQFiGKtpPBWFW001sC/yw3G08HtiNx4
d03K0nmCpAK8jQn6CqWl662pGJl6ZqJK0NYI8R+94Jz6ut0Xemu2nk2QE3/+WZ2A
jHDvKiDguMRNexqWoWJNopdvZogvNUplRzS4wu7g/3W6hnuDn1Hunm0qgc5WFbwr
d8awnPaLdgRZInnnF7wxIr9XJnqHE5zW25YZ+zkHfn5pcZ0qbLpt1SKFV/p3MeeL
q8pIg875EYhoMTGiaVDRRFJoot8kkJXhxHumR6emnxxy4nY5875XJEIzeOsaAZHs
j5LrHbcDT/TFoWROH2ML5GCPs29OGu5TfD/zVcSUI1YftQ+naNZWAmFgmZ1mZdO/
WjavAj6iuhHUBT1zdtUoGEX81QFmSkfiTX4I5jm6DbLHmga7hKOPFNZeI3u81tYD
ZufJtlROSHGa87mUF/4lWnO9Hj8awM+/D4NxKHHAaEsuTVtDptwXmzJksliJMi66
/KNqsiK8HCNhDNV488QEIYnx79EwRn6BS8u7X5Gr6m+fTddnXib7uSR+mLbNxnWq
VMPrSU4gOxK9VzMKm83vJJAxODUPtaKwkgNmUxuN2G19nCqLtuEk8bXkTKYUmcAT
GQcl6v9GQ0u8v0Ie1y3N+MYpLKfAbB85uGRQcNSd86QoHYge48Mj8Pn8cK4sowrX
KKwJWhPArJy/XR9151pse0qLmZQvfFcHL3a+vDayoiIixMzKw/0KqRqPX2BZB3pZ
jfFHgwnPxI+MLxTCkdD9dsfBVOXiChaiha4AGDpeubdjcH+JZ2DO2defnPIPLDJf
kD3xKwl9SBLYAJcLYPpVSQkeLQVW9pazBh9zmygsy8qxl0Eo7bZxBHXUiFXaPcwJ
nJAcaRFIujaF8O2ytjkjmIoXsFhehFYqDDoLMQDFUkRMUS2aWoH5+Ukp9eSwfGH/
xV72aAZV7lUJjno+sPdQM1Nc+2lI/45+jnakHq1mCkBbsqyHEF5Z0qFM8FFOOz/d
Qn2USepVT3fOksrA4YoYW3mmThmGz51ia5S2gW1EXdnatqxHKSMATCigAFOs/edC
Yk4RJL2nzA8oNpHvo8anR74FpmN5L8E+rtp1KkyCOjuTLskAVLX/i58lsPyCPu0Q
dN8sVKyOJlv4+QgyvgQZgofQFITdbLDrniN0FX4hK8dDYbPK2BCl1161OlLIVbzI
6Z5Tkh9071U9uCVHSwQpDYWW3bodSpOg/t8Z0WHdmVhDEq+WuBmQtU8unB4t6t8V
+tx3jfuV6AsmDRv5npRUGOJXz7g2Er5C6K2xjgfi7SVxqo2RBDuKjn0wU4rysBVl
423tYLjQzh3hkzY5Tc43Dl8NMirHijDrjAAuhYUneNxPcLaaYFmXXlrUAVGZwPpN
ESHZ6ECxA5hxSlGT/miIs/RKLa4cOgBoVhY523/BrRHeG+qbjZc0rHQuqzMsVFGH
c06rBPFp2imk2w5QI0NTJvfDwtDqOBlEiLoJwHBla9GvWMbaEXfNySoCT8ZcoUSY
5AoF4WgwDu1ePk+MWMYue5t+aKgKNuyHdqvje3etKRYcaAb64eb3j3mdcGjzKy50
o/NM7GxXX5Jt6rlLHnHEVAF1iBIEuUuRWcnMxntTRDw6Gn+GtPSyRNoK+oMmcFUC
BOHNp5ihHwwNx6TOXjDGPOHJ+3pIbqlY60D8XvB4KafNESjhp+4a3blA2UVUCvhw
BeSVZYDORjXhQOvivXUVVfKj0CcfOBjfcOjp2cQFwrETVTXFYMWwRwJ+nTxDRtvE
c40ip0WeCEsnms9GFWXao4qxtQtcTYaTQoI7Zg9iUPUwZLdOaNx23UraAt5E5G/b
ALM3zhTZZCeqTLPOQUGRQ9hzB7og3sEHPOdkfdVPFg9SVzv6+AFB4AT5+7I+vY5O
+1mI0bwOvHKHk/dWC4QeepYLZzydMs5F7qeWB/oI9skZlNYwX0ZDQKEm2iJ20Dnb
rJI3eizeJKCyKIF13gBklXIUXI3Uz65YR7IKNqyUGWX1gwpD60o+ViV6eNYDPjxI
V0BliD26rwHNhyQnHOTIfQwdKoRQ6MabILIH0wiROwjGLSyaf/BbowmnM0NwAHj4
WhZWVrD77DP3B/hXQutaHupYM+HJE43YW5fIV4tzOPFvH+zyVNPeTQrm+rtVour8
bU+Og5CZimQs7rJizgETM4m3xMGpZRgTiJHFKcX6jQfDDU/J+Yw0eymay+I7udQD
ptFMpNdluA3Kmfu6g6CwzQFP6oNdTBstCPLr/BhgsixBqaQveA9lqYTRMhu09KEh
KPekmttXsSlPWcLr37L0zWTcoMxporHKPHfTQwsLZsiMBHE+Je7DmbO9cwonwzhS
NN52xwQZigfLhWdeUTqFkQHPJMv8b0/4fjlBHCIRcTTup4kiZ95tDkTtHba8kW48
TS9IrsceoDGseqrBzRAi8o21Jc3jBn0PahEyMVfKGQVrUD5OIwDBQgNjRE0KPscr
0Yqro4dlpmUD2jwxb5cTjQSL21+nVmoEIIDFMOhr8C4NFgjuhzOF+0ZVCyFlZUYF
osd8+BZB3yN9ytKWc8+So2Rz07bMcUhIK0fgz363F/3HtftdH8ve/R+TI9e3vOD9
q5O71mHI7BUhQXTJ12UUp5CMwx0r/tUl05tAWvglWEz+fPpstTm94qTLAU4FXk8X
dCxeMqaVcUzRazGA3s/6KEYV31ukNj+FbKfzjdkb59Maad9LWBcu6TQXSrqszVoi
LE2LHHxtTLNoqGW9N41ijVDRCUTeA4hWEYjSDf0bMveKuqSaq3jqCxyqaJ0FPgDi
dv83vYd8kQJnHhbS//dTnHN51N+rwYtOp0KV5ZyCMQG/FSxVW0lIY7ds5vDpKT6P
bDxZUs5X8fbGqaiR1MoBikY19li2BXMVp6Yt3aOq97Go8vy4OcQw81H2/H4nTz06
gHIit2bs3xVnyTVtYsoadPsJ2Vn5hFsGzWngKkzScU3j0CDB6SnxtHSmbl4RIQHI
k3ToF1/6RPEOgcD6dya+vdEeD7ZMhs0XAI9MDjhaZYZjJloyRDCwqW7n2T8fMj9o
MP/cbECk6c8JZGLMcoOu/q8NwThqfSphV2WDt60M9k94APX/UU6deKAdRuovPJCh
HeVMK45hTuizlr3ycdbcw/IUFtMsxZdKyPMvsRAGC8WbtCsIDuK4kiHNrHfTwGcg
gmcslaVXZGsStY/WtUdrJpYCSIjqUQKoW6BWwvTO+UbNxMzIoTvANCRcNOwzJZ5Z
mv3o//ZxtnVxI8cFuAzVp4AH+144NkcUtTrCQ+M4kJxoZaOMAHL1KYDm2Ov1Y6Wl
0F60KIdreZYG7ImmrMF0EpuCFmlk5nSpXKIFJJyYL+RedObYqODycuhKWxqX20O6
gkpR1DutSLPjVTCfPToIWEhebAoz0ZX2wlgYT+w+YAfWE0bJBLlNsIYgvmg+KcqG
ucQKzLKZZ1gTLStHy4cul7gdKcXA0b//1DJZjWM0UaglIOVP0OtkDVHeySdoAdkf
pdFaTRj4st3PyyIhxTdrR2KaYcAlbPQndXTF0V/seJi3RtwToZyjmeYffQCkUTBd
MN0wRffpdGLXg+xGiqVNuOEVkjkmT9PRpCaao8gFMK2ciQ6ZXMQAteVlmfFjV/+u
pML1NJTAu+0FXJSrMiJCbCU4rp+tsUOWhuPgQSX5IaMtyjPnKKf9qRVAzD6nap+8
EOcE70TO5DHPryM3Y67+cD5BtWvgaigxzBXiA6ig+6Je+DADYm99K4p7veQwZ2D3
YV7dnuS4Qv8eYRFpgVNXHMq6cLog+2895PbSIT9nHYJQQg8XDPXDvP4Lj+bqW6BD
pgGRJXPo5is0hrBFt6+5B9GDOn3zC3avbirAmu3b2J0dDIN17I2yAB6IXvYRiZzl
QgZ+BG9Br74nnVjuM7Lz3tHVX0WMQIigZmT2TFS6NP3ohkgAw6uCecI6Sh1Dii2t
yvhtEwxrkvRyEg6Wmb6p9f8ZA2JBJHaGIYslPcHVsDzw0Gc89Vz/4P8woyavsnK4
JbSwKB2pJnPJPA/vLq6XAwzAGlmBxT5wqgC6GR7bEHfrjPv1lO97OjAandJm7vw9
CbfXeT9QLZDdEzBJ1dGlXxkLPU7r4NvO4AkR9BkR98Et1fGupk9+Ox3u2cX8L+lx
axQ9IVUYrUxiQM8YciBMjFQ0zsyJdwC4B8LHY4T5h0jKrN+efSGV3Jk9xGOD7CbK
yQTUbe0RYw6FtTFMxZVT+8JHXfFJpy0VrfFJMJZj06WcDnbYgZ2RfClMPRDn/Vz/
grzP7UAnLcqnPaSxg3gcstkRjvrFYD1cSVlwBJriUBqUTjb4tm9inF0rLLkqu00f
F43XvqSrED1hv5xUK2/VfD6BgU6WcVDzavPP3/eG+TvuoI9/uSQknBrLftZj9ru6
oPdhYQu40ASoivh3z7rHIA0APA+TIHlXV+/VzzirOH90o6Cm1Rd5XCJinux3z3Di
4O/zFDsvp56VIybbJAEXa+kkLwsM1awKYcnkh0LVFEjJwSkSRv9Cp9n8l4DJkuJL
IbZ3GRRUZE0/yrl/0Lsqr4dohoOFulUY8Y++ZMyLzkIsZM+vur3WBw4mjwmNskmJ
2gJZgXthTNbUfYsRkPkEanmdl5ghwC9HrVPtZ2jNMm3QM01NprhTIWNVpvR55DFs
KhMKHYWE5x/I5rsSQ2O59OUf8F6WwaOqe9ikq7429J0vrtpT59RlzRGbgxHj3aWb
/AEiQfbcM9QAiz8i9aToS9gfHOOoFYXM3b/nQIzzqp//s3GNBB3RHeTp5V7GuGul
rlB6zRxq8UT+wyWXMZn8Vn6lJbBFIUdHKVIhaNlwVJdaTWnwJT237RSoyXCOw6mu
5Fyn5zqM4zMKuYh9xMJq2/nAVGEyxlBeXVkktGdquKpdPpD90Nuv3j99prtIeCm6
4wDreLPW5xRihtgYIZhqHDwZ1CJRtbCLBgAGrDSJzH7rLrzEZVX/dRlwnxiUQqSY
MsJ2L35pIp/SoSD1S8PH/UAYCnkhbhBl7RVRmyz2DScvrNKx19i9SXIEnKVFBYPW
kio4WXZG9vXDYzrm9+ChHSfeJ9LCU1mE2lvQDJNZA2I2JSEaGJOXWqP0dz0/apPe
1PGPsVxjgTb0YnyryagQ1v1wro6qVJxgbOfhCTET9U5hS/RzbM3VpZ2JFK4Yzuns
msRrMUFlsqsDPSkjnEALPSn2Ox234SGo3yKUerplA58LspLhHRuGSOiEHn9DStuE
a7EXa7onM5b0UC+ljFixMUJLEOqsR3DrIDcHKjgBumGawbxpbwoSogryWGUvEMtp
0Qjl/j6rbW87XwIbsSTEtO/JxwQMWkUelwzPczZWnL/UGKMkkBoB+n2WDZBL9b7D
9rb2dJC5fuKgdw2qsRTvNdpjqYKAy1+Lq1haIf/M3Fw2CY2OAtubxMQ54A0y/av0
rUPws0jeJCrDtNXq2w2xfCWLLOejVyjNJ2ltu3SF3m74mFDSRY6e6wijGbRSfus8
BJXU6Rze0kJsutCf8IM/Erh+tzPKlwDeYkZ95JTrFOgWzcPtQGDHvxZXZs2Gtz9c
UHE7fpd5cpgTgqiKcumkhhrfgns6j0jQ3qAH/UNYnmwHI1FNmQzwRpaUXbGbfkv0
jV4nS/nB+aTm1VYpS3EgBv4XyAmjj2YUMkwHEaoDxn9OChYXgdhSrReyLlV+zPoN
0qgRwQGXqMp0qw6xtnfgH38y6O9Igmyg5PKUc4+x7xZNDbNQltgbt8PXbI8jADGT
Lx+QLLiu4CJlf3D7uYGf2u6rmZD0mcSnswxlF+mzVcVH4TRxzmV7vkLrkWeLc7KM
8vOpu01V7VLxFEJHQcKzUSK2VePZN0vxPW7cML3AKOg1Fs1NLTWDXfIzHiO0x5Iy
8StSRcsV7k4BXyr7nvXV3cAn7jFg8aeOTkEP8KrxbGyQvl1FHTIIQFssRA6ppRWa
JKlRzRd6nU2RmLNJ6VuBVUOAyRloyv/mkUDtjj+FM8J+FJX3v2bNqKMdkHyAsBKw
IEx7nuYXySw7wYYAxRMTEDS8Mn43IFOMpd7TV8Nb4AXQA9JrUNwBBUr7t1kEfeGw
iG+T2tGNHyKzoJkem0cNa/tGfw+7QuWYTDgPtOnPbiHPzbQfzwMhbpvYEdE0DXEk
SRxejBLuRpU7+3ON08H2Lq5CQkFqr+/b3JQK2f6aB7tAICXjVYWCZWzok3rtcjlz
ji38Al9GFKRzMKtmPBmMdSS1Q/LbcfBzbdHkcwqHu5rvNB+bd/rX5DTPltctrsZR
Xp0i5zGXpcT76sOlqqZVo88YWljUMBxh48muWtHA9HQx/Ip6yupf3ajqXVHIqDtc
cOWqV1deZDReShl0rwtkfwbztR9uOV1c1QEX7M/IqaSpdxTCQmLMpqhg9+mHWRFw
ilc2n9WYVz4r8Z0O//wITc0rNCP4E6L/YwJ3E+SOtZ/ownpbNsMgCf6RHdiIZGFK
2Q67YhxETGVYRSz2CclejnaItsO/37dtsDjjC3bMo3TeFjoHdIt1G3tSwDampmSR
GwW+r4jmmMWCmVQz47Mt62jt7hxM9NrESFarkE8BWhSPu8ertOc2F4jaYWY7KeJp
hc+Q23MnsO+APF2Qd041gbmUDK+GiYQ0LQYrXGNs6WIj1t5uQb3rpAKtDO54OUwR
NmSN7JWCvwie5+KKa8JFDWkVUvCVFrp1A9rAXulu/aTz3GD6Pg+I4hWZRLlfEgtr
aljIoCMNReIceP6T0oT+oZFFk2Pc2mkHVBrEP4DQVQOe50MujyoVtuywd5dJMIiN
CWP5mEVq4JNe7UirPakYJOlZm0Lz26lVjZZP0wY5BiuPrTREFpVvH4zjHCggV/GM
OZe1ZOsuFZaqpHmC38akIJrnvnpuOkbI7VBBLduT2QIOl8UIl1WZfVbX6Xj8lp6e
3nhzHahCkB5jk0zWxNL8tF5McfKmkDiytjb91+zO1SFh5Vcdz8PeMRxqip9HG2yp
U2blWHlKlby7Ojk44yURk8MqnuUHvxcEFAcXUfEoUN+rozWgrFkMvEqwaN+ivYdd
Li+EhkizuKKZEXDtFVivb+use2IExOOs83Tl9cj0Eu84gJeOTkJFXEB4gEHajSdw
WpcJmbhN51tmzJS+sg+7wCnUOBq3wd7oSMxgslNaimF54rJQ2auIAHoiTOLumyU8
P6w2YKtHGRL4gjShyclRROaXo0VBTltuGsXl3CdXw45yFyLV1S+NY2LLOzOv1oX8
BXgxpfWSSAjQzdq2ULqZWIZwQgEnxccca8BVzb05TpaL+2c+fPOdJIf2wpYiPgIc
JgJxJEWD6dN2t8WYXzLSbVChy7YZvA8HHPskSM4mGsc1QCynIoKSwTA55/7XHXEN
9lMLE9MpPLWwigk2yoQ72+Mj7Kq9ZW0KwQqYZc/iXZDFWUKAhi/Czug1FkzffCNl
Yodty2TK5TD7KTfoZlcvEwilh6povIt+xTJEKn7zOiraaKkpJL4113f89B1cwynv
A8BMBSwl2QPHZc2Lh6vQAxPJSycMLQW8DTEXdruzCZ678f0kB7EsY8Mb06Db84hV
L+acWtShbuU+0Sln1S6k5dmgcfYIqotVCicVTRZgLUPvKnGvcr3z1QL6D3pjTPhU
/+VUQksMqEZCOFobk384JTmLFBu0ao2CdndLrGC0y+utBvP5bbadVtYrE/wATCIF
NjQgJH4IgzQPR12fC719ziIfWqKvCs9/uch9yvVmF8VrRVsqyGtkiJvydX/Yh5rT
zWgq2jll+MaF+njtbDEcvlr1P9MfjQOWZb10XtfOVzqnQGxOGTVtMgWrHbkgxT12
nKRuiqf+wHsonpXDaQtIwJp2X0P8yU6iHMKj8yervF2e7oa2z7mJFYdQ4tkpZXDd
jfVho2htC6hf//tCQchI4rXDdc/XP8oRb44wuFjawhx+pJa3/8b3+hp2hiCS371C
EOBoyFRoDI4mRgzO9afZRuO0ZfOFRyDlRgJs/r4lDLIqOE7IfFw2VdLcKqehHkHW
0jK0VnzpFWPv6ee7IGqS2rlJq4BM62UN46eNdGuOEhLF5Vti5dVq1JbqVXf62Ask
xPM1iwV8h/VJvASafDvFeTG6+0E990B1UF5klde3P4lnhcvBv1PlbjL6l7PUzNiI
JY12BqDq218EXY9pXiChL7b8us2aN74IkGSM5niM/fBMkAVzFrNTvPuppbWQoD4m
vBjZAfKG/4TVddfyBhvCx/J3tx5OVrK/PQ1FG2KW3eG94HnhrbIh/462fC7og6Ox
iHiQXATH38yjWZ3qKWRTWv3wAtC78LTizvLV+xyXLtOR1OBQLNdPE3oSMNknTUmu
Digv6PiLFwcrdFFWgv2pMmR2hShNu8ik1Y8fbtdiwVXjom2m9qS9hslwBuugyFax
dQEX2VZtEGwCyG5P0yuv1RjLarP5WlTgC9FnnZB3KHebZRJcpmP3cLxrIdFBsIJr
copDik6hEIG7CpEhGubjyPYkzJ3AMxwLN4IS76K+380ItEslcM2pX4ibYgKFidCb
Q28Jlt2KhHgY/ZGx5WMmxWD5zaykBLIP3Esscfvkzzn14fMSRLegPX8+bmd7Otkd
9B43ym+zHKNrb8/96AgWxTAIycDRQHs9xIDuCjaMXrUGWjluKZin975J2hruN9M6
hW4cSBLC3NXOc5qI6QpkaPU3bC/QJGvasUEbnSdzmwb5OF2K5DFj0dQ58hUSrJBE
vRNycZt2CX6QFNrOu1R20RLpqzmhnzPVdCzmJ8bWVRuIMms4YBwNbxV6yPj3m9NO
r/n8gBn/y9eH3oDaVC7PU4AO6drzXGOCjnm2o/zzy3goblMv94uXcwKbkwfaIdtH
M1jJw02NZPBGOqCHvT/yED4YG/H63TOOIOo9Et6/MQ7M/j3+rpR576oWLadOO0B1
pHW587o9QYhZH0GSqKlI6XdHevQsNs9XXQBGV02oYqKFqebVSWxlmP2ntx2zx+Ab
/V7KwY4Y2jyAArLmVGUfO/zvr9VFEO1f88499zE5DpHTwRudSUCS9UzEQ7wpiEWU
xfYaCzXUSNh/dnLB8SuzUL6sh6sA12cxsQ8FRgrYgjxw4kOXp+B5qSdZ0sfa0CT5
2z+Df871mBG0TGMAkCvFa24KNkmJaF0OcpiJRAsZ1p7ICd6B9b9eXpXNXtWUuIKd
kD7CNhxkFNDhiza1RoaFf/Lu5X4/oCqdOeZNRmA+HrgElMqeXq6lHTdufZcz3m7t
Fot2AIse7X84OdRt8i7Rn6qjceJHTn/jCozLyg6JEhrcey5viUptzBnQfDbC7QPe
N81Cf38JwhowffqUTbju0i7/xKQRGv0gnDwdj2LQcgh/gk0zsuOR6P4vwo8QCZPj
FEqk+qaJF+nEtGxj5InjtPX1GgRrUq7aI7ZmSkqvOSX43OuVCQCShPWthl+/YZ7x
6bX1neFcxJD1WuIri6aQFAnjpaIWQeUu9LLNH4Pl7HvCIuxyE1J9hQ2xnZJijois
YQtNrSFjdpxUfZo40WSsc+06De1GrSFmnbxuvZL7oQRXJx+MQZdyOhzn2ghsnbSJ
KXv4ojJAOtIFcCzeiX8768jzyD9FbwhvHACrDMVSPX6Jr4jjzkuUzBKGl2ts17UU
FYSdlG+pxtXpFE+5SUfWS1s4SLc2ed7O3kg5pKlWMKunZooXZNS8IY1Ev+2sPJwK
m3UunbF0+VZBqnQgUT95metdKeE3/8kjrVljZmmGZ9s7pTUA64TdSbMJSx32Rpa7
AhUb8MI3vAGbGsNZdsS7YFx2CxuXIXfOKB/XB2GA/7ZHm0jPJjaY2EzzyqZxzSd2
bKm2IJ1Ujq/iWPTCcNWMJ//jx7J3+2gRDUDYAQoI7S5imPEnA3JCc+IpWRcnvu1B
ZCEmXmBb1cQEHx1uiiK/IqWCOFy8k38tj09S/WlcsoVRnqAteJ1j00GL+cPfc/Jx
V5ej4IPCrllKPtdXencMM7S3MSgLTrXCxQvtCodb0UyVJiR3coCDGhQta5H+MlBK
P3ZjqnK8Ea0uUkGnxZTWCrtWn/bj6a/s7fQ/7qVD1GkA7bJQQHtVMQB62a8t3LZ3
AIy3fpkLuKwkiQ5etupbzuoO1s2kGk73Ma0TkhDeorSxrsTELIEiEzSKMQVWsqDN
HXQFYO5i2B7FLZJYSDOZ+VRfCxJ/oaLEZtnA0/tjX1Kzkls6OeE7jEdV0fW+v5ZZ
BLHrnwr+Y6BAoc0Yhi5B5HLeQxk3b/NmMzAevtZbvHgrbJQegboDmDyKSB8vTc6F
4vLYxsPaQjzMdoByKGLQmwC4TAGb593WAk4sr988ovEEg6aNiAu00CaisbxN67Ov
g1Z0hZp1jwmP7s28CJr58HDSMiMuvUd3gFTtTMk0mepUNeV5mBnCFdTp2ABdDF/W
KQciaCNjdlicSbRwtTYLnihjKcY1aV2NFxyu6fJj1CTd+FVke8LNuCYiG3t0nFi9
N2hfQHqteCZ6SMe/RNLayQXxdTpOdZoIjjUanLP1QQ4aysR5UYjBA989OHGj4OMI
k4ukr5KdcZ2Ce0iYVxQbdef4CIWXRst4ySS5rRMulnzmIovcctwXxLPvuPa7vdRH
20TwRShd/35CwdHMuYez2J/PA3MwtJ+30ZEVhGWKPtUtJWqqIRo3HThiGz+58r8i
3mTmUP2A6UO2El/58/SGMu5vwAG5y7HPh/togMRAm9xt2HbNcr2DGHCKG1SvyDXA
3vk3GDm1TTgdl+w7dATO+a7OfexLuxFwJVg8TzWRBST+KDWANpXWKeYtjDQx+h1e
GrmhLi+HbDfSN2RDWGrSbJvoZp0G0/ErHER6knYdQeW4CKWm+KGnUPX8jI+QYWC1
fSkwJQ9Mpj5uQcinWoaxxvM1HesGF08urf6v2EB0i9nZXWPGpPMi0XjpAJyKdNXN
YeB16TN/60E2lMxmTh0TtHZrXAzKhcbRywmTmudMqo0QMhDSlwEu1y3Bq5IK7alm
yp4XeswzO7RS4p95/sWFvxT0g0a2RViJnZjudjxoP1cX/k6r2LQE5JoNDcmn+2+f
YBMyWnWRcrnvHeo8+ePibHOd5az9ziH1434Z4e2aWOjMyb7gifZEfxJu63iVw72h
FXPyr9uy9sFpypelgK4+ro3TkFawCoyzrmp1t6l1HUXTX8FtJMP7woFnxNPHjTbw
c9cUXHCJtfPP5cvomjZEqh/XRw2HUofBXuPgPUr4WmvcpgoEmUkAXd5Xl6xWweWm
r0ZlFxFBsFF9SZPtvM0RpAARGo7ZRtTTSzK1fO43w5HpumXOm2UrmGN4dS6PB9F6
6BAuJHpb3DFRlWFFasHrcnTRUY/c5YSIlwvGtff8IhAEXVxRYYCY3aLENGjDRAZH
OqYB+53l5lJEQFjr0dgUSGx/ZLM+3MJLFWHbZ1LqXUKp2ORzwIvQW03ZN3Sw5AuE
WVh/lcw9S4pQnRkDnG5eCEyNBH6GyfiDSe4OueRGedYjHClp+xWbMDhcxlqhOG63
d8fFEjXTDc97hC6QxK5Fv69ugBLzY3q0lPDhV+5acgyiGQD4Eho4cKz8CkGupkCa
kKtBc1zrnfz/EBtRpmxOV23lkR5DNzLMyanTyWu4pe82HKD22S3NLU5z/frvtDjN
nv51vSFiI/ngzO6Q2geeMGfv+DgrnGIr7EWjqnxMxb2uDBn3klgftoTgis+iJR+Q
ZXcTBa0knfzF3jrvOrEdOInIx+atafDJwRSwRUZECx8Bo9RY3Gq+HpVIWJ17WTav
ockNDWjk6Va4lBnTx8ZihJTfOFWjy0ot0L2FzQD8xaO25Fy7xanm2dKT+/Q9MR4v
x0/c1jPFo26c3b5dAEC9FNjKgMJLWOf4yL1fBd57l40NLL14BeYHpnan/U3S93YJ
JUvnDbPPWL6adI4UVYfEgQP8Tcd17ELj/DqzIgtHHOfdfd5L2CFAMS6DiiRrqMZH
/Qho+pt01L3XsNiH2gZO8jju8crZAee0+Ri3++sZLvTYdFNT2+Sp5xyXZ5sLSksH
8A1HDcHfXVRcJSZdSIkDOC3uUKWZn+VGTqXPWNxsUfXVc+VZFnu4MmgbeJ999mMg
aCxeuxowVaAGe8oF6Ua/h0TeAQaDQsPaf26RWeoMUDRhOqnF8f1e0uNiS0y3l0jP
XibnAHWKcZaQIubof5un5CrHJ13lyH3wvIFs/4ec6RrP1uBixAIcqmsDS9OknwMM
80PcyK8OdZcis9PP9TLgvFXj8/DcCEIVNkPJgEyjtzxyKR21ErezY2ZEAY5J6Tus
oNFFMHGoq1aqMscSCkED86nHLiKwJmTPkKMM1G/nouClNZOo33cyxKkcABpMIU4S
zg/r7pIJd0jSs/9Go6oj6AbTOML/pmOJ8YTimlwzEXHEjvZrV/plQ1eD3raydP3j
cqvb0lcTsBP4yc4DeckGXSs2pS+s6fV0zT3vJvKFdVgFaN3NaKrQCzp9HFUoPctO
D0KJER4uMP5KgnzSCB5tKaQ3rv9LyCiJdk+14v/n2a+HrI0T/gZe43WLK0pYQIgy
eoX3h6Uds7216HQ2cp7tnB/XDDrHAUw42QmYotHKJR2xoaG6bm0N1fsK95V8ElpT
dL+lFSdy/MgfjoI4oTOdAEhCho6cP6old7gwm5S9B9CBA22J45WG5pZxSsgwWZls
ejsVmCiRbO2m196ZJD2E0kHDcsyi64BmKTFM2paVXCdbJlDxjUL6oGbOaUnPWY81
8Iy3+klrQb9ZNqgbNwgXIP2nI7clDm+uWJ5fmYUXqMN0cJ90zxqGZ56mPgBng7PS
PsrYtHNUJsR0BmUOcdZ3RLMPAS7/CneCxygzsJy5h0mCBaCN2+Af4iY1soklSa6D
KHbwCjrt3Jcbk5iDYIrQgCoXITwspHbqcWUPqjYh6p/upcoes2Vrhct7xDqWutqd
rKH3s/LCxrHUe3miq+mh29q2c6GcRDtlUX/1J/ai426gXnq0aUx5iGNB0wube6z9
9/YN857HWBCurxYIujxJmW6d06mRZjy0pXC88+DBM/OufXW6r30YnnTnJXbk6Jf2
kS6PvssHyymCIADlOzsPWaJdKjHP42LPPEiTEnDkQhxyTYhCCbkgdFGldgMbqnDa
ZnITlDSNOM+dsiViMRg3MRuwa8+/5fHw2uEOtR4qWnAm/Rjanf44q7wIr+LLprMw
XAy3zvSWJd1f7Q8DG200xwfhVgpPkXeQ79xLrHTpqXsgegw771mKGCF+wb/51g37
JzSD0rGTGZMtWtexLGu80ewc4cCHYHGQKgGrukjSDTuMlBunEeJ4vH/uJ1PPdWPV
cXEIMunTy892KP2qDJJuDYFp05LUrjBKiOgWgIQ6O84bbycsgpD+6xtAiHUCJYoJ
hm64yCAI4y3x/gwnGSEmmj0ZITh7FDGls8QRNRG7yvIxr5kzZv0JO/mjrfvJIIR5
BMPKRWBH4W9eGmmajMxcX+EeQ9H4UGD1gUYP5nSOdCsiglqfOZmTVJ8udHNK2sC2
kpzeh/+PV+LwIIieM6XrLcrVrP9PYfQT5RpW89/2UvZfEfHOodh9/guCebNw6/Mz
Z5uvLOWVCWYyIl2v1n6L2UteXmle3oG+MW1QOvfgeAV0/WMeHzNDrhFxBX4YDJ/H
bfHlH9KUSbp1r5+4NsoKY3kQPbHHVB0LEakrlHatbzOscKzR9tTw0HffcxRIdm+g
ouwuqSyZSWUs9C5LQEGmlBOFPg6Plhl+Uj8Ht4+w3UCZAFMjWiM7I6JWjGXnAQ1H
o/jgr4sS+ucooIe6MyWTD81pNZv6mza/ocT8NCpn1eB3xUAV0LoFg+RCf0mAWo2l
16o1X8vXX62inqIsvW0fz0jcneJJ4WNGt/I5M4zcerjBMTGTOgc5kUGU85RNur13
EraPGiaAh5E2ls5fsk9KNU06uXW1pJvyQUJTL/BpUF4n4cCm5KLPvxiOjC6eOb9d
K6rkw/GFYLZkEh/opMYvWzEpeDh0mW3rxdAUR1rKOqp6OGxPyT8N0OikFfyPwJAq
bYU6qMD6bg/agQOcd3IeSuB+gGVbEr6GFo2yMoF2TS4MhUnaADXX8symL1KncgYl
nOel5y709yvT4jz6LKy1I8Zvwgmzws5pIJI62XyOC7lwbBjZZXrj+iDUNi4qcINE
O+Rn/Wa7wYEOwP+FnpkA36+/th1qt5x1EpwuGJvt1k5IPF2HSk7W7FQQIE8bSgwT
DpEaYQTILhVlNXhVSKFGdbed2ywkCqb+7EsJid2VSDiNc4ycfXSHdrF2dj4/OklC
YjJeguSpoHpXwvd+omkKUt1FhpwGmGQHB3/czFRBQZGUqhHKfP+yf90XcX2Z5ywu
aObfaXoREX2bbBm2Uppf56hofwc4E1Nzp6gP+2CCUO2JxtdevkITGjSQjXYhI0Dk
AXNMMmiT2ccZz7NcZ5cdijyuxVqKSd/C906Gm0x8rH8HtrZT09EmIRptW1RFbW0I
IOwWnOeCReU08hePKHKK9jNvp9vxH8/3ruDdAYVjaWje4CzUrImoA3Vk4x36WOvZ
nZeSYNI5U7UQ9kkYT9ihLEM6J0mor/Tt3CDz1ZSv+i4yClWCdZaNY1rpxl3DmGfD
HdScJquqkT2CDrG8nsXjR5OGKj961v6H8+YCm/HfvcKoJeWCsWe2q+8sgMbYtyi2
3lM0Xc/sWsJkp+VwiH364EMyM1LfeAiZcUSNxtwQmG+2gb+iLkcW7KWMUMkggczs
o1O0Q8vPPn1/wzwmERzcPL+myPZyYEZKkzKHC7UMnFdO0oKCGLmQqub5AfhXfZyZ
+WuOhAg/+PAV9vPgsbpO8Y9j33T4DLzGFaW5lP6Iz9UmI7VlFXreR1DjLNxyJTCv
4KvqTDAfpABJepH/Z0k0UkmQEti8vMdiCjtROwslF6lX+TuP7+BQsEsvC9GzoCNq
fvLFEPzXuOvL2JnCc71ZDSSVwhJyqO19sarXTKYOuyRcifFkfcZRNEVwY38umyDz
4Bw3vRSbd8EEca8LRagoUFP2qXtn1BNhMPs2JgSdpCpxtlvCNwaPtMg/c4jCvgsK
LyzrUYzoD0b4UPzghHJ1wUV0gefU+RmLn4l6ujl1pF1D7hS57g24N9ShLr6MbBRw
6J11kowZi9kBKG15jdFIOzEzLfBrNCPjJIATIJI6SRVVveVFdzziP/R7kOwYOKql
XMLsOiGBV3tKf43fl+Rht0GI/H48Ak3qKDC0DzKiv71OKYt9ONLmLKzGJWKCnS6D
foKknLPsCAdUUo+YIeMLcyxm1gEPfTuEeH15w+DbzefJy/Rtgft0qHEjDW3wO4w1
OvY7GYFB2v4/aUZZsKQYh/hS//q4t3ITwT26ovJFfPn21CgA3Ze+D6tGI6x+bDuz
+hnqeHrlzXoAIb437QIoHir2+y3DbeD20aJs8qMkH0LRyiUvAGNEIxN46l4sPDqS
U+lAXCTcMEDLfyTkiKgLl6cA7y1zFMEnib/GhtWMsJRg/vzbiD54NJ657u797CHP
fBJjC3x4tkOGb68+79U1EvTIJBZzGgYU1N9FTeMVBanLOsrn/UNoqAGDANTGwQTl
M3cAB0AL1L/1iQrRxcP4jt07r6RjndpSX3In+p/lfUAGG1m9g9Cciu/8xAeUH4vv
rEMHG5ljqFMBAeqBg1NlF2iogXuLzVQjCr0/gQpcsg38P1AdM9qEn723g4tVkK7c
cf/BC3WdRjYtydi+y4LRqSLsGhMsQt2OQxXi0Sh99dvpJ3v+u6QtwJEmgz3qsyWI
X/l0rkuJlJRJGMSykpNvVV68NpFG2QjIO39mc2oR1ddsKuN7M2qQ9/0GKHAoIrEI
9yslz3QbehDenjr9PWS/quRER3ql+WYxx3nCLmvHq11BjA1RaKjAz5wqCNukSnRW
wDox5asQaN9FXGjlamzdD2ShtvCXW77w9/NCFj1Q+V5B02lFMon22SFPYwYNWgHT
pkNC/iZ1GF/pbjcqbdPyfZ945CwrDg2dd+UXYnV9J/TGGI3kkkV6Vu5ylQBxHyCs
q7qCSgf8JaRgcLFSKvMkM9m6o/UynGewfR4NwuEt0MkNQ9vItZD2ZRInyJRKTe6z
UTaLgkVHQdWsYKuT0+iIfuFjHs/Z7OyVoz7Y/JjRvv9iH0uExLOCL5bjI1t31U4j
NEctgXQ4fPZL3S7/pmP66RFcHTAZLvDh0NXrrTc7BXL5CwgFbUUgJLBnwz7IHFib
9tm2W2Mbj6e3QoqV9zm8vrW7buhY1Qd/3rOkr9zN0P2GnTBrb/TihmMok69EaN98
z262Ha19RmupgjBfFAHxdiOBz7vjBEIK8ePH5nQxUdiTeA/EpWsVB9NpYARJUEYw
K/Rwp6IY1t7qsEiCZreJ7FKd56qjU0UmR9+IEaPz3F29p35/GOgHR5BxQ+cwAzGQ
KSXE7Wd/RK0Ou2WJ9bzj8ttF273vR57mWaG6J4mUpndnJiL56LvZoNRW3wmoNvN8
/yyXFZ12LjPNBuvQxLtll2/qnrbD90Sr4XjXQ2/vuzy0yxK3vS4xJUIlQTJRsmjF
2kqh4j8yy+0FGE4LGQvEjBdoeWll/XHt1XyCoaR0W9Sc5QLRgeW+6CmnG230rqoN
WQX41/WIRaPMXZAkQCFGh2A+aF0BLsmvHMn4HxX5tp8cuKBtl91Tqu5ZGajR/NCX
GxfI1a4C1bdHT7RnGcI55qNNrX0uFtlyF5emHc3558YCRJc3VYwqJGfsZSYv3Xs7
MyoB6vtY/ygrrwbLZRuUkVDnm77upaEGG18OnfQ1P5NSxleF9s+WWw2JqnOBf8xe
TPPDZZLPUzY7gmfcguopsFx8pY4SIkjDSd5q7V2/xz1vf6ZzHJ4SECpMEXF0Et4e
ryxhnEj30Sw96w3o9rmuAbmJGqcvz13Emaki26tSG6XRy3nVMPM9N3rJ4xQoTpFl
s5ROSSCWkUxjlDBfnkBXBpDBepxqfvxRwNk1SYBcrtc/OyiyuuL3Xx1/ZaU+FLQH
Qnb1Ie1RUYAPX+LJlr/nF0G+xmxxSlOdsIjd+ePZxS1n01P6ss+rKc9KBFn/DbDf
JVP4YZQWyHZbCzUjoiFMkP9ldsuc1YT7LcqAMyYxGdi2+nkaiTqV7r9aY6ElIoQ3
nuFz71ekuFzrK8o1hnO2iMt10KhOmx3UUBjt1u0WH5pjXfrSnJ0i/uP/Hj6/pXhb
eoi/GwNHVNbniGgxLvH24/TXWh2QbyatyWn0znsICVg5BhvIcZCm2hCIRuSEkeEh
YEGmHV/CK09FarS666agJ7GWuGpRYNEafT9ZUt5OqKNCuuSx6L8G0/g8v+ZyJb4x
Rz860tVeDExXCF+vHzFpHqa1TLz87HDfnNdls7LvbfbhDVDcuqN8/tOa1MQwXTnw
4ZU1wdirVmd+IutqLFjKVpNsfAQHYj/AG2UAUwJMXFM4TL17sFrPgklzZQgQoH8O
jiuP5tKMjIL3enZ/FOQHKLMr2Fihka5pGzZgCQv4vcZY1bHEr9N0TLaxHZpXPf6d
AfDc92QP+o2s82YjjaLT4/5KNIIV5V1T32d0JGl1TEq9EvnL23+4MPbV/uBgOJjy
476W7bmTEz2/dnNhPH1pr9ZWhRGeqrIYWCAJJ10GOaGOgyfEuHsT1CSjzRLch7mw
jT4Ntl+ODbt/oi+GC8Vq7Cpgu0yZkooxxorbnmnE4wx/VvqRtphXVpG9wMs+rodi
F0Z85rAARbOlGl1dBpXF35rdWKkeGSNUcUcDq/FJsd3eURfdiZX4KdPXX5ZOeeBH
aiq8C1Lg+mOAA8KNshVeuIws1ogDuMjmF7kXVF1KLWNyBS4M0YaSDpQddZSJfPpf
k7LP6wAHIqkPDKWAElV8oWWq7zyA8QUtFMXlct8piskWPzhUABm9F64joiaoskuP
LrRFkC1KzRQ8jV2goteh0IRgvG0+l3NCMgD82dHYKkhHDlmSFS5nsD3mSnmJ5qgB
dVrlXBV+DMc5RrJJ2yjVgjS8e6oTQiITG1STJHOhRQVVlSc/WthhPRheNwq8TqW2
G/p6kjSBJJQPO0NPtRkL5msjNVfu89wz2QuiejjN8HPYUe5jTXZ1fB0k5RiTuF4m
1pZS3toa56pebV7jBK1gp0eScoxwKe2rPZJL2CP16qyZ29vmanx930Vsc8FjWviM
6bE+vEjCk+uQDuyPwvHTNPvCfQqkKMRBp6eGy3mNKMSJe7w6Op9pY0q1ilqRHsL6
SAGHb7NHCiG3NK8ZIiJNmbN34lb08D6yfY4Rk846Ke+eT2N27ar1/4vtcIl/W//V
TbYnQPBv0TpLRIlYFTuESNPJ/ZXpOAYedC7Wy2zK/aFSoRW16gBzf67OlpE3dFk3
tseGzlMbwFOddFF6iRLAX5TusNk4mSeepDEv5/a21ho4kRrbk3IKd1edNxvhYHGp
CzgVKwuVXoEPgFKQFu5x/nglnUhKHtvDoENDlRvpDLyvprSIluwHojCM6h3qPQWo
f5+ysPO0gDhKVF5SZ/RHbwjCKTGJdNzv62GJDxw4jcFKRRvseT1DKJblOpBJ86Vi
vN0zITDw7vYJ5kP1snFnZalS78BPt4MD70jMYmwRm7geGp69TPfWYi2LsJqcbwEQ
tReX4a0x3QZUb37Qf0+R9awofTV9lM/NcxbNOMSNpR17e8JgHwxj7rHlPjiQcWrz
rp1A/qaobSwF5ZtAoxE0uFbtPpM4dylHhen4+CdZO9880H1rXHS0gCfCbFGKahcC
gioVu7SX7czq1u8cL3bVDTRJ59KUxKA5wxnAeyzcK1xDfy6kDTX78Tdi+dyAMTbJ
/cydgq8APszpD1bIxIZenhZ706X57egtAdjaX5nwZqH25kr/xuM4DA0hofb04TUl
JF62RrgyXeqyh2hQnaDkrC0U1G5Eeh5vzXdOW0e6FzbqYAwgzNGrR9ZO466Bn7Ao
xixH3DNeMmihiOYLVmV9olWjswLTAKbMgJsPou0U4h9uOzaMxRD0S3QrG7Q5Vn3q
pMpSk4D8JJ07k/29qptkLvZd4Is+iBHUjT7kRaUp68CMwUuy0NMim9G5DSES4I0V
4DVAXwDCqHyYTUO0FkEW/gunH/o2GWGMFJaKVpQs2jPFVy5XpkbKhklrTkXCUhzx
XIkUgcMutRjAdJ5pbH6JBb+qfLlLp61lxXXQgjP2gkkMowfhpmTmh7tzSulmQJoJ
bJA7+UagXOLmkU3paEj4LJk0e781JDnpJzUTKMAMNve+uMkYZlkLWM6QkvRu5qMn
P2LIOsfx9DyjToRDLtIU7M8DaGBKQ0AmHi2HLqWhUheZRTBahOm6Ss03UrVPubI5
JP8du1iMZDZNjzwLUSu6fGDMEieKbT8sNpM924tVmNQ6I0zCYszP4W08BrPEaryg
c5h21v+AsSYENqRMvG2ZmfvCbaPi9s7imUy5SJ8HHSVeTwwisVhk47GGJWpfcBRl
wfejEWt+tugblef+ivBBL8umk/hz0KCjCSKgrPZ+FREb2H7ImCQpb7Vfe15k1eZF
qeJfIVQbjo3OUOZVUuQiM6ZJLOh7W3WQ9Olq7hsAXUnJnd3tzm/+aDq7x1UtaTmt
GFgSFuAi0HXnjJ86U2zQ8p/WJbqx1+J0CrbJN0Kl8C+f5qf1kvw9fbZHzBo/zuKw
Thc/z0yz1sV5QUat3jPK9Fef1DdOA7lXZ+bOVQujb7yAfsFylBD6hetKkW3RRKJg
M4EqDChl27Rw0SfQPCDMPMOIxf8+L4JnYJQ5W71pXJ5vF/+PjgFYWMQsOXDuMm1z
CFvgg9OT4J0T1I/iGG7PQGiVUAV1rkgEGIcVzdOXHjY2BDBcV+AVdKe5UhorCP+/
U5gJOqAC/M0jtXXji04M0I3yHjv7ctOS+Jnp8aVnyUce811lEhJZVbtr1xOOKyKK
5DODMessHZ5eGnyn14hOfHX4+wdnbJH7ACJsrtzAYxKnajzJiGmEo+Hl6gFQAinS
UiN5JWLQTGfiXYwRQavrjkSvTLHYdy+lV7x05XOug5SK299xxfOQ1gM4IhcW6qf1
XXU9d3mET2G/8o4YEWBWitfn2muUpQO8SzGXHABbK8FF5tDcV7S0+XA9vJO61bD2
hzmCHKzD6vRaQ2AJ5aKPtD6ulqflsJcK4SmE6jcnoLoUvKYTZ2OzjXbshK3jLIx4
5GHI7mhCLpcJzNGsHhwuK14QzmLH+1tsTBRRRO/Fuzz2NTCZF6fXZ+DDxW6tne8A
AQBYdfVT/zusaBluzPYoPgBqBUJt3mCqC42VuWiKMV9IY9bnt6PzXXC6NjDmAmZD
ftYG13MXZyND9HYqBoIkDEG6eDcSgnRqd92lSCRAI5YNqJBjfoaCucZwB0SXAKhU
kzFt8Lk/36yvBW+lLz91EAy39oFCcF2l1h2lpTWtswmU/GloinK0wxlgmS6f9/e4
59XksKVGod9cbdLkvcKAI//iTHsED5b4IPreSPxE4sKEsxcNK0dBVlMAkg22bPt5
55zpv7emi/mutPwhJXuWy0egQ43TTrT9AvRBFx8KPkurr4mCjf9CwtbfjHYsK6N3
+sh4J3f80KE08ElVJn8RA/OPMzu0hGs9QAXIY4jLI4x+qObs4ulKhcwHm4pcrraZ
/GK64PNww7XRB3rdyYP4jenIG3Iz2BPRZELUT/1mhsHqQToc1t8HDdG43Sc/4wPp
VMtg4dEMg2Jn5Qywrzb9i4v5VyPZOKblD7Q2Z3jzAcezciYQIkdlzPfGXIfHk5ar
l6QMusziBO5aLSMnsewiYgwwhCmars+HnWurdEHcTC91uPejaGACN0HNpnVSskqj
y8+DKdc4rIbY4gvfFKYArNjPoaROIkPUegJL9KjlYqMpUDUD0Jy/koxJ3GlNmD2d
0l6rQFGlGIOPIQkfVTjOJvufDZp9KY4fKyzWFE17ZT/sP7bDbVbv13a0BrU0jf3Q
hjjZUrOXrdKFGAAUrIAvlBFP3i6ADZQRdMkWGw7h5FYTTVD2KCsBZW/M6buys7ef
ggHIll8VMPn2yR/tD0fcwwUTJClAWCFGw+u1erWmZrH7Aewz8nIjHREk05ZbscjD
oP7Npqzf29NPyrCftSA0HHUOCw7FTMJrDGj9IGbxaiFFRQT1dawYy5Jl+RcQLU+S
whokEYl1BwWJfx7cPd/IdsURI72CVvSYwFtxn+cpHywzZjJhDbgm9bQqUPgJYrAd
ZQNjyluxU1BLT0xoNefiffqrXcN/Z6V32URZUKuYZDFCNOn3TXf+ZURQgUEi2Ni5
r8PRenkQtHbgPFg1G2g2Q7SCxFPcRAGOdUS4FJtE53jhDX5MC8dFFG/DjRopQQJP
Nd8u9E3mt1qIMNU/n2jBznYXDBc0NJ4jZR3BeWmjlRTSgn5zywjAVcGbcv/rJNuv
23V4Ri99/PtN88fykgIumRmPJ5Z5bfJeo+v9L5bACW4GiBZt+FFj40P43eEMZa1e
z1V64vBq5aeXHpiI8okHMIe+H/DIclsasg3r1ZAf8WXuor+dcaS6R2Rzr714YBoc
pChE+hYSidiSfk3ji8Lajuu28b/X6ylSJp+8rj9GTCWteqUv49T+s99ZMj8jiuEc
FzWX9G5C3Fb7LAwZ/Rz6fp6DV/iBeLzSdxswlqxVohpCNePeVDJ37e88ijoxjutK
kTrXOtMoqFUbthQpZpCegZCvtDLLp3UgDxnvLl39r4eNPt4WSGlkopI0WQp01qd5
5agk+RKEn4HldsD1y1cWP7A9Vi5dOG84hzS959Zi2EkcoewF5omvpch/aKT9XTr9
SMtiukkgrS9vWluUcRz8NDJThIYXejbwa+tGR5+9iK7SN/G9SkzDTxpuPbueymDs
Es9miDgX/sYaxEzPy+uL7N5Vg9DruPT63XDVO09KQKjcGEIcsZ7V28opW4XQuV2h
evMa5dBHFUxoJR61SuuPGH5mRgXSpn8dB9yXcPQ/5qV27u7wknxwQcTFxTwTqgW8
7avAgj87t2/KFjhIt4ZFkqtW74y48cj7nkdb+5yuCD3IXByeplBavwAExvoHU+Ai
7DU26NppMk3IzxIsal2NRzOxNNAc+hehUCUw/5XiFPEdU5+RU1Z2t8xZDdCyXiPT
20r0hD2c+V7X20MwS0UKnn5y5Vg8m20PchjHApbY5BW7xDsWdt1xm+C7C/63/gF7
VQMyw7V8Sz+neia/izo7LXyoj5NWwTRnL/A3yoKCemwGRrXDH2OtL5KqG4x9JAZ9
7Cv9JKNuoD5ecM2S1pDyJhIdT9rbB1uLtyArMLjGdvD18f6r9sjZv5T7TO0QQo1q
6UybXSX0z2wtNDnvuSOHGlcFLC7ou0E+QbkJrOmEtz/A7lzJiOxVv551SpnRfYcH
m/6ICED44OHdnj6Vi1RF1UGW7oj23i6pfQOKTkre033QMPv+a99sQO4a8+FUytnO
G8VC0NiTR02OV+8a6tmoK8YCeYkfgFTtHz0kZnGA2qw8pRo1cRngr7ckL0UGQqaO
l/88e+RgzIqb+ncQOZAI+3HBY6DiwAuYUe0Jh3TkYbTxquWSmohX6CTMtvG7KKht
qyueMs5DwkjwV2UmixiC8oSfee736JMOI7/8mgECyD95vAlufOBC3fH0wfnNvajs
+n9ozlaDFDJcLPYtDEzp7sjZR7wJxev+FqGz0PHSa6HSGh3RjrZ2Th+EshlLbyAg
BxAdfUmqRQMD/UwrL2cpkQuY4xRVf0BrhbvGRPqjpNf5rrXK0JSK559NYd3g5lEG
a4SqemRjv4gjCvqOQVvQa1qTvfZBQExCLTcwjZGirhUH43Dn52w3iPWREbKVrKVo
OT7lt8GUA01WLiGKGMI6NTeImwxj8tYLlU7m1BkkfJ62jHH+LDKRXqL4sgAzT8+N
KQs8F3O9R1CDwKn6Ynzt0oTh7+s3kW0PzbWbDM/qLIQp3C5tqvA01f7RyYjoyiaJ
1Q1jUCtyVlTrN/gF/JC33L1NE3qydkw4jbq1nansOXuoU1Dg0rxNW4oG1kkLXdu6
cJwW//2PCgIUavSPR5QcxzeToW442ELyJ06ycY1XVoC//nihoGEb2IMsH9mHjc14
VUM85Dzq5dI67a4nev0qV+KnaVgTbGmWmBueqet7m0mo9rZm2G+a0qWy8sFSRLUZ
ODygWu21ZPSL3u/CJ0LdQ/TREEoz0y4ZKKC2emfzataWxTOkdUd9NWrFRV8X7hyS
I/4GIk02lDNzYQgvJWvGl9DWVZ07zoggfZSyjzg6i8KiKapcYQSBOjz5HvxPB2wj
bC9nz0Ru3ltKDeJhCMyrGx4SBW0I+p4gCi4MpKBLRIBVtvmgApVrMsXrRdWorreF
hA58Tv4RF/Ng9pGxLqFDcYrUj6lpuPFpWIB4A/5xu7Tuu8zctot2rWSEYRSo9NUV
IT47lT5MUtte3UE/p10NmAYG0cuC8elNwg3I1II4OT2DcAf4y3jOFTpTCOIsdSK0
+DAqOzkLw4lYhqF1hfAa4RJfgdJArA4FcSK/UyRhE7VptssbbWo1kbS/SPcLa6UT
XWalkldBeasL3bTuBT8LjhGdNqLv/uYOxJpzU4ga8HwB4aP9MDRMC4KwSEFFOv03
4xkuBgCnklTSzxtpvpZmdqBffivjHLjrn3RK3NxUdR8xSjnvdbUeB06rPEhUQwa+
km24ktHtc65S+VtoONduDqCGtIgWiqdCGwwPTYJGbAxlXUSfZ9Tp4wleBfZKbWUt
CNkeJPOs+MqhNBik56zjxRk89lme1Bb1fZ/KfGsgHsgRsmT304Wtv2Gy9OT2GTgC
hH2QjAx1BZ1DmE5T690DhMNqIr1NmnOoFO3+DAMheYnXppbswOjUaqSFvozSJQBB
RYLfkcvfAJFKSHwdLu1sW1D7lSZbAyvK4o5F7A4GZE+gJYR/Lu/vzgVP7UJo6m7x
g2/Stj+DPR5BcHWaB5zQmCw4BpG4dXZJKB3MWWzlSHuK5ifPC3aBvNNzwi/1Pdcx
SJpHm4l2WlADzo0LaNm6R491WobfzGsFoLm6KTSM4YdjIo+lDKtujUK5mvWch2a/
S9Pk1ja5mKGxGU8x7vGOoIyA4ZVFORRB9e6b8ylHcjnqQh29PGtbP8/Rl9F/U6Nr
tc5aXNsCdETgiUZ0eT187Igyj2qR72adPxdKSWIb+A4CESxRSnyWuewcuVDx+mOE
lbakdWtJmbqzMfE2BwHxncDHurB/rtCeO7WgU8Z5Ale+VlV9KMboYiKNm3SznWg2
DeSrO/WqFltRhRZEKw1n+aSOe9tb/Q+nau7ru2nw0Iwn6l15mJnusKsZZXXH0cp/
2iqMh+1VPnObT3q3JOA06hdcvzEDKA1xg+zSSiOlxCT1IhsgktrmbM+5+8uMIJRr
p1FBzBiiERLJPDgpuMSwIfA36IvthJmLZFS2QGfxSg2GxiCCKVKfUTqvkO1DCaAt
Jn7ZnCSW/EDU6JM60+CsqWS80QbmEhQ7n2mC9zQ23ZRhf0JnsLn6jtXFfBhHmjl+
AgPD7PDP0aWCF2rn1SUUwxKbGhFS3Hvrn9nyJbyqiIKSjYPR4Q78XCGb6RPakagw
ZQExBajZCrnZXgLBjlSX7/q/Cgp0TBG6LSft2+vQIHAlQppzUxVtJjyEQE89enq8
eCP1Zrn6jrSpT2mqfwR2Qx8QVfbdAAoKa6TbEM5BVqU/w9YpwY60qVwILO4M0ybh
BC1SDPd3YuipJMPHZw2RF/rC+6xVrDSuhSfW1aJDYiBizT3MuGBqHGFrz0UM7Nu5
fatixj5qYO6XpvsQcSGzQbzCVO1DBleOStWjwXlGBSfMbDS7Ebv87lQFM4kO3GwP
2oCDzurAr/jZ5o/yyA6Bc+1k7QwaVE23GZhwAY28nlIO1gDTgAu5AV7XaTxdxVbK
`protect END_PROTECTED
