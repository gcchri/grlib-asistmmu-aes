`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LfV4hoyIGt2wjy9DeE6YrxAhQGcBq97Zf4aeZ1QO4KBnISoTm1RowY/Jiwpf99su
CVZAouDDT7GCZIFpg6eKJaX57R4EbZ2aH5pfMg0rQuLlZBAN01+p8fi4xW3Ptx8n
mI04GubfLjA37t5bqXGO/ADVLi8pSZkvKJs3ZRnozZs0ru+fYQt0nlPIEE2kiJhj
+uiUZu0ho8iMgRHDbqNa8i0w0zrZCroiN31/dCkG/O95TG0XnAU/RZz1259zk9mP
9qdrKVAL7Se6Pmf1Euzcp0VVWeM3Bg/rIMxh7yfjS+PHohR80K8+x7kc8n5XHdYR
gG7Zt48eclhhFGipftr+VcvOETlc3ZdEPaQGEcqjHPFmf64cmQsxUF+RqyhV59U1
/EaUvjIMFTzFsg5QPI6u8s2flqvxzsyPyCLL0F8SFd2fwIYvVyvyIJ+hAvl2vP9r
mSS2psGPE3pBwxCokiGo9RZRmmFBXUmOIdkK10+tQsatulm8FBcAf3PDSQ3EjHq+
BoltxLKe73fyCQxbChfSzpVt0ODB4FsjEEOktJPT3WGsK0MfJa5kc5Unsf4MNQcJ
xaEvFKDiEN3m53cR3WApq0cpfbNdqOKPhu1gKhLSYVWqXR3HZnAo0T4uwazHBrTl
7pwuo9L8sIyhOFETdI3QeH5FYhOKdCK5FWw80GiRvIUU5IaZIQhTE9F2ulj4KEIP
5ga5BCj75H9gOQe2MCJ0yGl9Bn1tLNiQZt5cMf37mhykt014b4X/7YWDloYvp2vP
WirBi4y63PqWYC/+cZYbEwzPBdfgW5emfHApRrXNuBOW1NcG9J1gl1+y95vArKd+
leMV+aeob0/p7uh02ZJhO2CMYKtYY0NPGN16Kaq3aY3ekfQ+HCsoa8l+b8Vm9LLZ
`protect END_PROTECTED
