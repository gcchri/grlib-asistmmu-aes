`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
byYiQRxN9ANdQbP8s+HuH3dhxtTktcmNgu1IO0dJtm8zsO2pnNbzQf6Uo9Z7F0h6
h4b6n7b0omu4UysDfikQeDoM0OTbEIBHdHplQRbGO/pgqKg/Ao3gmT7c8nC9gUaa
KW++IcXrEeVDIAGtGNWnOcsllA5YUh9F1UyUeWjxgzezz0/exCc5sScrAsGPRamI
jmqF+rojE16YWFe2Oj6iV3z2NM+/PNfiiZmjKurscaTfJAgnsKG3GaB76Ff3qzR4
6sUPAxBBuZxVQjdnW9++BPd45I16ZrTndobqLdcgSl45cDgyPq9aN8dn9i309/6Y
xG/fcI+42Rp6/Q/GY+1CjDi4GQ5oS4ByuzJ3R2Q0GNW24pdsl3bVlRgZB2gQ/eKI
1FmjJxdHW2pk2e7nS2pd0aHTcHzyRsL3Au9jPqukEyhrnavra/PO0TNJD57tvvAZ
2XDyZ1QNkrJ7nkNVgnV29urSEDlQha8inL0wl1rM4Z1va88VamTbbSn3QabzQFM4
p7KGH+EDhJ6zkIzG4tWEmtJVFH7kFzhqllc8r+rYWkQ2PkcHrNHWPwDGRZUqZg2L
phNwmHIUwgqbJL7qGk68yDykMkUNR9rJXqgnw8Q1xD8A0QOMDcsk5EcaD3mbQ9DV
AP3gSZzJB5znfuQJCF8ewayuQJu/1ObGsj0yJ9k3U45WjDuRC/Nk9bJ6nX/j/hi8
`protect END_PROTECTED
