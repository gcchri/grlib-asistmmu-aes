`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HWxoWOlcolR5vgh2gVVOLwq3hWm8B8EvhMEOPi49GBKYBZARh2XNJjeVc4g4b3IT
wptItaAygV5f2tMdnGNysP5SfZCIVCt2lDxvEqTwRwPW67fV7yqwvhSOcA0WEEib
/8FuW/NNbSKWgGRInZWX84VZFCqIjWKH7s3xUg/RynebwTnTKhMff4mePdAhZGGP
smTpH49vmYtm4VXBlA7HlE+cVi7AIfKSp+0artKj+keMQhP4qZCJM5I7QZZVt16Q
s2Jy/L9QcZ7mDoQF/HKU83Vi0wZ824LHsRX4Gu1Q2zPIyczx6xVL996zuhkltMsw
BBHeRjOaxSM8e1shVvwO9nE4Ko1YCsg2ZF5G+mGjWtW4E3a29sb9LdOi3x1bZLNo
FcCjoHwd4chdpUrA5s5ZfTk16qpMG6uo8cTQmfFkLTUvDxqpvkLh7QWvRXG0ZqGZ
rxBO8n3K1ZVRD24EhUqn1J5eWJqGlGwFe5wn3ytg6Iy0mIHdwg3ZcLLctV547swf
Gs406g6XPhTcAe63TA+02pniEYaX1RxJK8o2e0JDTDnbQVgih8+GgTMAy5PQagPd
`protect END_PROTECTED
