`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMviLoNzt8GGYt27ePRxccqs5AX/ccBZZw1L9gwSbVLt13lf6N6Hsj+ZlmF86AuZ
2ee2nJmR/osmKVcQETkNdOGxREa9VnCFRYzd1ePRjF5IQpz5pkIE31FqWN5xX6mb
Q0mw/B5XDJXWKpRHEWACk8qiROgLiBhL8no0rKSIC1s19laPsHo7yTjQvZaEJLSK
RxsHUcd3xrET7Jezo86O64zq2b1MH7r6QrTpqvj0et559FDpLimgcY3o5iOigGsh
tPo+X2WVs64i4uzDvivdJuL6SngmumdAyG+fvQuGiD5Fwg/M50l6jBi8U23jyK2b
kB1nbIaxoqiYcZYnccMzpMNcNRsklYfiZYh0Ia6rNYte5v7GakeQPPaHID7p6a+l
EeZzBCdDjj21D4IRnyJxaDWhEqBDoWUA1FkAE0Nz/fR5frb/o6vEwTWTrx6+8X4s
`protect END_PROTECTED
