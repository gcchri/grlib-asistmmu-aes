`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hQixBieBs10P3QT4L6hW5AgRPUEgvEqId5jqlBdex9twvi64JCxhwNVmLigf6+vG
OokxRg53l6OvpJ9vGuB0TFedxbY7g7GLy2zynmEAdbofE4mADp1Mmc/3YEU6ZvfD
5pRKlohs8oHnP45LWfI4fPMEMZ351swOZXuo1bAukY60RMwEuwtAJph0uXFKZN8h
trSVicnNAqAJtew0pabEXiZrUUkdl+jsKNSbMngh+QsRhtAG81TwSSznFduGpFzO
sTpwWryq8+JtWto1OfjAvNkJofx+HuI74zViKiVkdISEf/oBHBJ3hDSWoDeWHZ+A
2rUZHFbD6G8l6yPAwQ648Szly7O6jt1JT/+JZz6vTfbYrH+RKEDDCi2SGs4IaIOR
6GByXeFZRGEqEKROPYmQh/eXyazK9grQZUxGKOWtP8KY1aDmXAOpAvxZEOIR5Len
Cj8LVIHT4YXWUt3lTPI8Dx8PgFHiaR2tc21zj/sninsF0s0l2/uce9XK3Vvyv7+D
kTt1KupoDTVTtW84pM6r+6FKN8RlAh9j0IrZj95etmpVWkbZ3Ae3Algj5B/LgqxD
YCmgYyQ/bgmzlvAIQSQM0k3HBc6eIIrc+r0d5A4T8B+7kkqXYsFr9XDdYRnl5mra
KFUDjZcNe4ix0RzYiR6EPDnmGlVggJZ48uq3xhitQnnrFxzYtEnMn2kpP7Wd+m8d
0GtzozL/yPwkAblibCv+9OrvFKn988Aew2kjZsRz2InqT0iHX140KI27go2LKSm5
W/3zXMq9FW8oYrcwdCWVINLlWaK+YI9WhLFDSRcZ7jpd6dK9ULvOXs1jdOj39gip
tfISmK8dve8m1nUow8om6D9ZVTlryLyWs8rCFCk18JrrtE9htPVu1JVe9rigPpIF
W57DJKJc6dE7Qzhg6BBdJZWXjy1a2RZu4DJOSLrJn/jMvDaoyQR4Bp6HwYnbye0E
D2he1cZXGMm74p1OVqp9RZ+xeeQr9ethX6pLSkn0gHJP5hVZkz8vGzYdP98S5vNG
FNIgTpdtZgIdY/50Y4WxPA==
`protect END_PROTECTED
