`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pz0teTN3hWF2IkUfmICvQspzTVnfZMsf2qLC1XmllK2yx+2tccNHS3WKixF8AFVE
sbL+Q4MyRo/4XkHP8aciokTY2T7hNVHJgVdQFFk6nSwUE0OrueQ0dlzANDPWMEJq
2uuB/4IjSY2jVfcv4DLsjp8Ou5hlNLwSrMN+25jn4TJm3Ww3xwD8y7QSW0mCiE+r
KuSOIGLZO4mkni7jy4kDH2/D1eyYce0qv/m1vvh66Ll5wHn/8RDybFti8WK/6s+1
TYR8mXpKHdAsbluVGn7wAANfjdd7+Q9pZZg8Zy+kitHILQT3THVoSfs8Pzv/h3uP
7Je1ZCup8WVGRxwNGNlv5AiTxus3EsmLKJi653yokHl6cHhbu/sI+dJ2HAiz20aQ
vhaphJwyo2Df6P57rlfSn/JrGOKnK6S5M1h0xP3fAkI=
`protect END_PROTECTED
