`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXulnBOt8znCiiaxwlclt8VsZOjr6cvBA4O9frsYSiKGcbGvxNyeiy5EAsJpHtjE
feDuAKsglha4coLK3+A5+aKiZTf0kAODytFcIVBYy7ubsIBmWHFhxpvO5Z09JORM
AgHLALF1deO9ArtJzzOnDGgtJKn1a1+wlC9+XOe1NB7W2f9OpEksudkdeTsnWzHt
4/KI2VFZQMVAKIS4upCainfmrljV+gxTgrNLEe7KpwHJM7P6NIUl8UhOgswebktq
ULiAjQZF8oUmjp6xI2wRkDy1G7n3mvYlQubVlm6/bG1itmTKmeMVNW3LmrhdI2FE
ttWUuTxBFZPGTKeMxI5I5pvSENPdMmg73g8ZAu5Vt9JXUsYZtELQHHmboL9SZrpO
v+ZXjkVNgpymFGYWcTlj1QW9f393Ja6nq4WCFMQ2632wbzaui8vnICOLNTccaMBw
9hVdUIM9azG3VFwXCnPY7Im3RWq0JN6LjggoUOOlPqxjnf2vxDL/LfJEpA/YCQrJ
w3FNrBWlJpGvUGMHque640UEGjM+8v95/uXrFGlmtIuDwfuzow/jLw59T9uS24+t
E1q+wrmbme4WLPVhcEFRSEvDHSMg5q4kVIDGtF5MMnk=
`protect END_PROTECTED
