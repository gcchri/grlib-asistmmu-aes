`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ziey2NUYKpI6hJ8sbywuoHe0+1hSv21OQdsPvaxgKz/zITZ7qL+jJRLOgoECJPDP
BVdqSczqaAtVWCVZrXsNtyK/qilqy0Sq0qwKhXKtDS6NjAB0u9a69vNBtHS3B4u6
BRlfg8WNr7rtgiNYDdl0NRi5be7eeHd5d+zL09Op39WlMqa2R18wtWphgEPq9sXy
Bd3ABgk//U+gzWdtwv1lusAWiHA3KID3ebd1zy3KxOk5hjToWzpB4c5kgLygTcHZ
OZuRk3msGspKLIsWm6L1WjgerW5xY7m+2joz7hyofy3uoNTE/oW0udb4KhrYCwWB
RGwz/uyojzDcZckq5POb8HRKoWtTALHbpITRxC4d7Sh+GmL6hsPhxUDdPhCGPiAi
ktgn6vjC6l3KJJSuAdAQ7vA7xWBmfA8RYXKAQZrJbEkBCV1YaIlkCVhzEhtB6h24
d9GCDOOADgqgvj06vq3Qlg==
`protect END_PROTECTED
