`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0GKfWTWYT0BgzFtlCGvJP93bjhcwoh0mnLfzdvsqLPBd2gALXW1NUexxz6HKVC18
inidrvBLA9t11NmKNYXpmS+O+8JlOw00jQ0Mj5W5wELIecZf7zLQYcjtZDMSkVqq
jbPNhHUL+TpO4/a7xfAC7YR9j32Qn4WRKlZMqoNIGQdj1Sri0215sqAafTzntVoV
iACgh1TLyNGhs1uQntFcojsmHmXqg1LO8j2jAiluAmddP37zrD1BNRXM7+qrCUjI
n/LK3S4vCqcFRdy7g+o6r7YXPCUTxe5cev0Ag9HseoM9jjhcl3oKYG80kTsRnz3y
MkNFo0Dfdb2s2XHuKbUecg==
`protect END_PROTECTED
