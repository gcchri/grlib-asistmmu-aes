`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CU3mGcSHyh+41GB2IDqJREo/qkjYjCbZStWYqf+fRhpTu54LIf7DIAjB9poboMuE
r52cWGWO+WEufGQ59pYlZ/03drRmPDT75Zhe/wKY15UTqfetkfeWy+bY545exZEk
/bdr+vS0vWrsj8eeXWeYNy0XMC2v7TuZ3qn4pABONqgAisJqkYO3G+CLOp2JOTa6
XiLKpUUkjhsEXtj1e5tYHcPGN+uKT5HOrifklqMPUnwmnSrtFFSJrnpkH44KPKq+
8MOkLCHibYAaQ90kTal+KqTHSBGU2bxq2zwp9nkOGTd8Fzjd3EFm4b+jJBpJFLVo
9BwiXbMSH3rIbuKmLmePW27HZDTMOlcKyHCjTSqXd2NsoAAaQawJBNuUgmt3nKCy
Ax8B/WBST4ccrvqrPAMZTZqelrmZIC4md442b//3tw4ShKho2bB8Vx+sOHtd7Pej
i6jtW1SMviUfdFu/S8tXkXAcx3nAOrdg7nZK9IZXH5+Beq+2nAJbSk/88m9Pz1gZ
MEOS2kb2wBfazqd/TW1zZVKS2ulKL7KKQopVPk6Cg/1tR5eumThUDrNjUbbXjAA5
s/bgDYyzKSKk+AtLTcUXfGcLu1hCB7yg4rk55AATuaTu5T6uubyZNsJ05bYKYVQo
43eXmC0/qj/OchiiDSurk4AU+npnRm2VM9vdEppNBAup826xTxTAyZm1ujaoXngy
xtHyrWtxiQ67YXXptUOYA8uA2jPCV/OfieCWjhxsnDlrEV1QWIececWf11PSNact
a9UVtObInS1srLvIVmUZnb1aRB+wFyuBfLquzwSc5S6Yr+PkdDQ97u4Q3fQOi/TN
ci/S8hoorlMv0UEukfXagw==
`protect END_PROTECTED
