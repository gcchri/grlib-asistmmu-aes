`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWKjvM9iIFrkypcUiWauT1w39yb+Yc/DE6/DDMUaEsYjEYOl+mJ4JwGHqX5VlIZf
ec9GmQDoj4TnXK7y9EdfWHN/FcQJKohqH/V9CDaQ25VNp/ADtVO3QM4piMVF1x9+
RzZX2/MIX6u+Q1L7TwOakYF5fd4w/NLhCv2wbsAV0oIYGJnHbCkFXNsIpHlWzu06
RNWryfHiDxdmASf8cnanVoHb3t03JfsMfMYK3azgFW8yphTE4DevLv4wpFD7CSan
c7cx9muF7ODnK8f0Q8lX1DUlGmApQr9Sw9EJ2CdCO8M4JGJUZQJ5P6ck34cpaxh5
QJQaHDFngYYsF8pT9xKRKwvIrNUkMvjyEkrMFg3AHtc=
`protect END_PROTECTED
