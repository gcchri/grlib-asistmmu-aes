`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sKlBR1xvgJfXYfdr6TpOL6zjsaZ2ANElu1rl2mmuGKd20H5JRwbgZlcYDNCr0Cry
xIOQs/1bM0C2/tyHu8Pj9m15xpvcq0qqOiiOmXUXDz8QjXrdcoUHlXoqGEbJZ7hM
o8bPLt74hMJBQV2sDIqPSJYL2iGffKJ9HZyomuvhss9J3mRH7iSebF0cpNO9CepG
wYAkQr+JZoFdEBEkktyw372EJ+I20jtpuirUWdBfxc2/D8SV9W+VTg8hjKqe1S3l
uttphsO9XW5r/1rhrl4hSKerSjguFFqB7sV84MAB62ZiZxYYIBJzAhByyOCB6PYa
QmZddkknJI1iyPzmPT0q/fCiG0j0IRK9Dy4fM73f2n9VrdXICMI8f00uf/GMH/RQ
Z1kWRrrO3tXNuTwcD08KrLkDhnoHVr5CZlrwxPIPDYozEgCn9kIctK79zoJ5NwU6
iBtzuGeTTJ6hJl25xRYeDy10zWLXpCNOqyPjm3dnyinYhw0NOSWBwO7D7Tcy+8aN
xxqbRo3pmFp7auvZZg0HlL1JKYKuLORJqtET5tMFOgR37JO8SF1rkVMua1kJxM7u
jrd9+zHpUdPOyFpDaiC8A8+/x42o9CN7FXtACoutn92hwHT+3QFxtggQsW+CLHic
A7ou860H173NTm0pavNktqHkTUKW3+nG+QG04QmcP21e1BfZhHSClByiU/GMv8iS
8lqmTn7jiQ6825XUHUvQAiPC2w4cgCAf3mxgYUfH8DQGRPpW9Li3LG2W46xbeVOV
4FJXz+dmOWS2BeDOTpAMgUlYhLwGKct4WhT6MVwcBgqc38criC5ka/1aCDXVIU+/
IXIGkIKegPGlKNZHFwtZIxgT/YLwTmtZaeJc/xGkHTHIQtaC0Vwfn6GkEN3ezgYw
oijufO90N1hHdW7SF3D2kYwKdmfQEuVnTENO/ysqG4WCYIkhRG4akh6xRWLgcAZY
gUEUUi8VtK34/7Vs/6RWh3IIt0slzd2pP17N9DdIhWLzHjB+URcLldb+wbT94Mj6
QCVI5fz45jFbc+9m7fMMGSK47ExK/oQRR1d9SaEYgqt+4XCtI26IBdbFptFPEV9F
jpyKWPIQuGqRIsiCGN2t/f3jHkkUUeyMOgJlvvXD9mCaJ0Td/TsTH0B6pDQwvLTz
dyMB/cfzs+DsdCbE26apqRuaPU0eOzausqvTQrPSYe0ojUzFVM04hpCJHlf5167K
ggoRt0UjTQyV+cZymEbmcUbpa+vnpUElPQseAont29F3UBzGMNEkcdnsEd8iS+kr
ZeLw0AGW0cLgTAI1Gx5QctA+STtk2ySg7SGcAG1LYEGofCRheaLkcH+oxUq72lIp
DjlqrsuCKTAm6kkIXp6FimGwWKoLrtyxSWeCirif/hUYApt96DitfvynOv/ym2hh
Y8FiIelaH+JTbOLkfLsHGhXuLHPKsHdUhF06HBYlLYrTBXM9SkEZ6o6NKFDMmqtY
CrcCmknXohaHHU0RvMguBG1MoSLWcj8fSvGhJo+a7faFqXmthd0Pzyj60NRcTFKz
j3tRKskNXlSO2gy14b/cINyBCi6VMAKjGzd7WQxfDl0tdupVIYysXDiwkbuFEPFE
1S1V7D2JrkGOMiETe4vQuL9x5/SnkPI9wdkVR7PvJuvvhLPEYnKU27cyIUrGgwtG
/ZH4RqZMQ6p3v9LVAx5lXtkfysqCx4P/sm2IkjGWfK5I74IEqdeaWvtmdVhxibVj
nvDuQ/BYhI4eeX3H71xTSZL2TQSm0ClGswKBMfXUyCx6FBccfPcDNRLTJbbE1Yoe
/6dF2x+4A+gAG4jUAKe1kWxCcJIK/iSSlATMXsNwsuJ55yD46/r1e6Z7CompEDy5
oeso6zxDfhHvNbxmIIq/VS0mt4Xn7YejLkumuQyATrqWyfCsNfdUxOK2/mt7R/XM
cVRqXPAkjux7gefbH5jHoNjaDjfugZvHz1A4qQ+3AIS7uOpg1Pw9axb1iQwsWNwn
SbzY1yv8LI8nzLXQKyE7JI5/TGQWSNhZ470PyLigAgarlieLps0wktsliGXKUKDS
PSCKesAviIJD3jSLQkTQWQFLugur/ExX9iZTs5ZraIze5E8pTpbE5z7OgI9NOi9T
G/Z21zmofrMhm2hGm949g93Jw9VVwAbfn/jSbx/W0C5hr/nQVkpfCw7uVp9uSU/C
q1Zt3/b+Jk7oiFOt5Zn2NCZ1137/iqtBPnYn8LD7uFiiAclv98kulm3vQXoDGlHK
GSRwn4Fd5rdGQrCCs7wHAtB/Cpwb7c8i0XIj/rip5qNuNZQoPJnr2ThwnIvBIXmW
lY2l1M661hOS3663rbluqYhkNbTkx9BtIhRjE5xrpI4bcyr65Si36vmD0H9iOKKT
0hl8Vun/dkLWTGzO+3OwXiVjzzz0M3nKy6mYSw/ySe6Nu/2B5n9wA1P0gZ+vRnax
hNQfRSg5UOkf8gp1MWpXUoPj91U7fiLqGptY4lKJCJW98U+qz9kes0sDpk0rU+d0
7fL7JARrd2mgYWdvfgXqIREGVmN9qDY3dANSqX6rcnzhi0uaZUA786BN6PzDGF2Y
JqTQG3qZXxBKQ+XyFD+klY8QA7xjO9+lFCdBUfUVbjUA1eUeDvsjtTZR1GO07nhu
kdtbV/3L7qbzsdJGh3btNmCXoiDTwGh3KVqQmKxknIcgALV33aX/BpLRPV4qLHnD
gZy10YIomnxY6ibonAkj/o51sRcntuUL5qoPvWvyHEMu0ej14+zdJmkMZY/f6PM7
ZvLUm3dbvtSJaJAhfKqKzrFm5Bi736mWkNfAQUqGDLqHmY4zXKsGBYdlBtHpqiwi
ph14IPaR96+bzFVfmU2rOvKn0AXWliIwOUXseD1FUsExVOAaFQ0c7ZEKix0VffeO
uVtu2Q2Aru7VlMxnL+IixMQA1aXDNOG9SpPZpHhJcGt/+5r1pHQoMAnF2UBOtixL
fCI/VFD51kGf/LIcVyP83Hru9kU9lyTSghf2zb3oEynsFXJPZartbdOWJMcjzl4J
CTr/sErWsaclbcmm+Ha7ZIfELl/SeF3UQKiQA/X3d6netxoTe7KHcGnh3YhQ/0en
Ms48Mzw3rb7a78LOxx/hI3QRjpMI9uSAAO7xFyXvR9ZOgzuADu/letjCIZCSs3lc
uDQ4445YBByfmwJVKZiEuynhCpVABP4ON83bquGMQNYOuvggY2XHUQlXerfb6btc
ALEnoyJSPUsRdBNFd/0U0gaItrieD5Kw/WQuT6SMYxCDLyw0TVcLT+H984ph+BSo
CYBb1L2Ml9njCYQ+C9tLrTLpceVLdeHDrFibj0dprKjHbIGjuzZgDXT9xmZdYgTe
WlsGLD5DoEpiyPGU09CTqScjxmGrQKZdRsgDmdNmP0ia2V2WC4/Mk1+qyPQwEif+
3hHCF+sa+L1KjtprSJqi7xt52s6Bc8td62IT1l6mpX7HBK+YfH0MU6yWVM31aLJg
rGuXrciHoMCAmNUKuFbwU8PlkCmSy9auwsSGcPROBwahyoKDjLv1a1wugMT/ptW6
pPEerbX9Yqnai30ziWqfzweDPJetQAtpZDuXYJNa4OhV9XVfLyZpOgjSrRqioocw
4bYE/16SVqOn+FV6EP9gmuV7KGn5QqO6vll5zOKnv0ZM5vZzBSMd6ImwdO7a7fQ9
E1b9RHFlWYQs+QcQj5idt03tle1CvxNunuLVRuXGinFwAg08sOCDMQSIjHUFXicB
yodLlMqbGohWlk6GCaVjTQeAfMsnhD+Ktnrvxrl4kkE0sHz0K1WX6pEc7k0xikVS
MuFsX+o7WQJd21ltGprmLHc+jYmGVxjTNph0v9Kjs+VHpLk/ThMeH5kISgulIqKD
0hGvuThPwmqgsCYIxt0ZsT4FApV7HYgmIZGL1+41/g4=
`protect END_PROTECTED
