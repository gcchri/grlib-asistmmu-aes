`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZWzPzgI9b2VdjDE+uKkZnt21AAB8fojuReDyD89jJJOVTPVuLZFcK6Qv4sG13sE
M669gXFfKUN3QlK/T9DKVGdi6LK1e7Bh+g1P5BVa+TVUGrVXRrQzwtyM1LhsRHhy
YwHqqdE3BplazTCEpZ1dEfzwPg/jouhqV6NeJgliLU8E95xmEtJfyZ/UlkbsbJpt
wekgBQSyI64ewyDYWobL6Vf97vi5Ubs8SqCUrHoP4fuodNU1QXUNpVpp0jFYKYzs
s85xQGkLIy0jxVUuk2mbmRfH1JgYkM2DibSDJG1XrnusuN/20y9agrh7P7WEZMwi
OcjR3hv5LFk/2FtDBk1zXQ==
`protect END_PROTECTED
