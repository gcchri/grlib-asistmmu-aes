`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iez5BcLf6XIjwKITDbOEmsxsIzYDCWSQC7ykfP4gA7gEx5FJFuwnjrit75AZOwih
Tq/sUaw9h08eLnQXcY7vLHFJKnKAy2AHWjTwuFKL3N6HxW471x/ynAMMzxNmvnGI
GTq14NlkdROqDbivonxP736QU8eOndmNpPtDJuWPyb3TRcAocWtCkJrt95EnoaMa
o19TeEjaItU4TKEocbeQA9DstjDMXrabf6w60rci+X3W5i487LyjcK2zTIYP3zck
QfhXIDpguNfHUZS+TxbK8gcCBscmBVBxq+zmKk7ry4e3TKKU1bYs522qfaEjv3xQ
WccfuNMBnCchsGlBmHw5gQ==
`protect END_PROTECTED
