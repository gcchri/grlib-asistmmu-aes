`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vKspaCXIim/MsMXwl+BBF3/DSVXs6Z5XRO0RKemlPr7bkAfo6/lsUxxZM/q1Bqr
GIj0MOtwAIxT0GFPA8JGyuwtiRG0lrq2iPJAHsbxMNmMjLfDiJSClln+Ev95A4ZD
0q70LJE1sVEp82ZzkpyY9gPUQpMcYAZXCzvykQrBKIBQrpoGNcweMDrxE0a0FRhr
06w4VE2VGofT1iBsOzM7Z/zFepR1wtpouQVoSdqMBi0WVbkaGq76K2Dij3kVK6bA
VG+Ay8xcP7Kp01c3XUsREN84i3FcvK4Q7lol2ZcDU/g3q1N3G3JjulvTVq315Vhk
eLrdVVJ9pzhnquK/DdMnh9MIGnOQ5rL+nbbccEecYhmNwTVLhc/pKQtImsd315cV
AW43Zx/R10jJ2GiBsscl7i7TtiaIZYrjKkXjOwW6tz5jLsBrUAbtlBIWAxQLafJl
msONhZomrPV7pP2zfxdn3XDOjhOY2Ev4WmuS4hx9kPDOwUIn59OTtMmmDtyzib95
mgk6DPfBj2mH0mfh364xfNm0Nuhlctle+1F/SfeMeUvtF/vuomIOWQuE8WAVWZsw
Q8IN53uhKOF+Y3HL3d+iegAiAAhKqkhyuYGcVyB+aEqm6FzcgaFosyzZxCBOrRqB
KXVh/W6Wi1gwZb7njz6llD+hF94Y4uFd0t4pNbDocUh9UL5QaquNhoHsQKE59jY7
3yrvgu19t6+lGQKd6oZNV1mknUE0BAqaxoKwewFf6Ev9lIlp35qeqI4WKHr+Wg4s
OhekbKrg5D+h9RzPV6DBdTfDXMpu03bNAaY5op1AsN1x2FMphNQdjsUaGwuWC5j/
e4iH7733bLvclE+nnl/R6aBvT1W1nTCFJED1CC+kuAMFKFL+I1ekKBZXRYT3xykA
taPFNlbCTtc1LUBTJ/tKXNgtdHECKbLOqhxMbx3bPXjcU8zrVOeaL8NV61kwmbUh
z7kT933mInMQLucKSw4susyVOO10b/7ja74mbHyV6AKEuo6oak9zVAtQHFN57BUD
/idUHklKDFGEumnXlbJuUX19vZG1QiSNftauxcsJR/8b7Tivz7lIIWNRHY9ggosI
wjXZsmV+xKcaONYcOcISbAnla9/mcKm+xAKlyf0lSSOwqXhsrumGK3QWttDiXY/0
nSpkP6OZGt87wQADnsCb8piF9xLQ386lR/viX/iK+2PMq3CqdyjMp0jDn9j3Axp3
ynI/0BSc9SoViEHc6uyb71vm2Nr+EOTYGqJt83suD+reRLDbyz9MBBxn1rNqTyn5
stdnZ0iXGNi7tU6Z0MEBSxfUd6QZTWvWwCk0kJzuUpUvNanqzj6MfUD5bJ/iLXJm
pE7GUcuTyBTMzkBkS3rlcNzxjBCvTEtjtj4NCTC/9TAKFuJlyvbbKyUui5UZ4087
XcVx23NRzAMcIXfBMgDLyzb1THqlhUnM11WQUC0MOmRPeBbL4dTx78SB9rUZK2eG
RDowt2vkRo3H4feVSdcuq0PKLujhCamNtb5vdcp4wJYwz6kM37FiCrGGxhRy12DB
ZZSrJi5lLVnPUXAoCFp8pBB3p9qPP+oIZPZyIAiXwgFJv1epq2mYA6xY38jF0YrE
g/cYgJMm/C5DUBt97oubTlGspREFZt5J/GYKZtQMweqoAfc6gPZny+buqwCl9u7D
kox0vUj43db+9HuzHCq+bYdeZYhIfqwRu8pBdr3r/XlTMjb9BgG0H4A2OGCuU92O
a1VapQxad7bPqTGQbmWUw5ZpwVAOXxzQ60PPo9goAKrGktfRv2rntyntbksuB9EP
u/2lLQANgHnh3oGI8p9jgQ==
`protect END_PROTECTED
