`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzadL3LHuvt+RB2wOv2oQaMtTyiPnOUmgyaLXaSkZjpUi2cAbOksMjVkSy2jZGTu
+/+0tiP0TmmMXSm1XGUjjlbTzuoe3ez9Q2arDQF6K5ReKeC37bbjD+DgXgpsPyu3
Jkk1cTJif2LIORn7Qh3VbF40yODcBetSEFWEnyTUni4QuQoB1UIq+st4JcrrPE1e
SomVTtl2TkLmdv4gqkHml5J+WEcBU2a5jOSexmJ15B5DwkgcOtx71nsJ6hsiEOP0
Rrt0ZHHud/6ROD/GZ7HbITRPJra87i4ymhBdXZ0dfhUmshYcAs3bOIXPA7duUCwV
5QVtbvO8n5ZErM+CAAyziYEORM4Gzp6RlBZLKzT90v3sYUt6Gi/HX3WRQLUNx7pv
Ckb8cJW5M3ieV09kp++vbw==
`protect END_PROTECTED
