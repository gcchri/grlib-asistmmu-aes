`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YN28H3yxz9WP5jvfN3iQTYa7hZ2J5gjYwsfbtCNgAqeHeB6/Yxyqzan+Wx5WAApE
FvWu8UGmA0A6V8/weg+hvIQuwNcVfcPjS03AdkuaaTwMxBvwoOB0TpViqohIw3Id
Ek3h9Ir9k0BkFuz55zEv98WGokB0YHWKF5lhyN+eOnuYAuRpM3Ytp/eK68bDso4p
2ZnFFlUYu++3JG4RHPKusduIKuPW8int78leH0uXTCDGGrDjoL+qWaXtsX34tr+V
oOA/HUE4pUKA0lup8Qg5RA==
`protect END_PROTECTED
