`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rjl+GimJpeRauwDC8JjFTdxeu3fxVF992eu3JAQwejWMGyAfhT+6MKFL9tN9D/Mt
MmFDcdrc+SqgrBIXrwNKeopVr1bYQLnNZxDFgfsA6JSH11pjjW+1cL3DPo6vGIsa
ZYeBXFsP7xHH+nhqImEKbTzsbsuHeXkbKW9XW8E2C12rMTXhZpXDIaftv7PUyyTv
mXKvPmLOJtCmv6fY0MJasaC7lyBZuHXD3lmcA3af3mFkuNTvc/74JWe9uyFweapN
6VgWqUwVq8b5C/f2K8Px++MT+Hq+01sakLBfBuTwWXg=
`protect END_PROTECTED
