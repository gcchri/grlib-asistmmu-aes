`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aya+PyYVkf4q9UzulQ1FWArMDOSG+VKcK1zdPedPNw5Jt10lgmlZrNur17aCNeuC
Jr9PJkjw7igerXMBXABk2it5xBQeIT8D2u1AMM9qxuy2CDgBI3LV2+Pmkoih+JOJ
6lEd/qA7fh24/iSQEu/Cj3joa8/QEjZmMK9LGb3q4FEFZjOAIqlF9Bj1S7cWXN/d
/iVzTaa8XFMnfQfU+2nlUMOR+E0ITl3eMkoGh7/qwKVrYVFxIw8rMOM2cE+oEbGF
BSRPIIzET8OiqYF8y5j1wuAxNEUnGzNOXdX8cB94J7oqAfnMBxKVy5tDZnBVur2k
`protect END_PROTECTED
