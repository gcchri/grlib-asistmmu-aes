`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFtcrJQBHZh3DAr1v53Q/yQLSgvijU09AdMFNTuAlA60MzWsgnRSusakuIo1KilE
NZ9r1tHbLUvMllXuGUByozDlEXObQNOgbNM6HdvIjfBJKfj3n3GaErI0leiM1vDj
5YCzhlDqJ/ehz6+6z52WuNsbY1pukRvshUEaXIWS0kU9gJvdpjyrRjZD6K7cqDNk
FK1I/LeqfWCcK3IHl0lrlhDoYuaAJnSypOsOB8BQ219MNJtDvklWjwBa/Rs90BhT
ZmWosFX6SqSF2G3EaBHFzQwuerUp/01j4PKYPibsz3ShjjDR0h3FkV5RyzssNeyu
Q7fSUlM2bdquWZbD4Z3Pg/wpg0/Gsw5nAHHIbVtm+Uavzhuk6PU7XlU1Hs4pjznZ
sMqyzTevR9M/K0S9zRI8a7zL0VQA0shWU6EccKG/RjQLFFaFMmoyAliSJ4JQQxKC
9SUSZol8PEVW5pdIYs7oDCmghrlMlQqS6P90H+rhGXAxLX/7BbV38n7Wo4UTcY05
17aZJ5iB4wCR7xXFTkNEWizPlXQunlITtkXRnmbh2O+6zDyiHStk55NugDKxv+nk
nEAL1uV8mmLTeqwTaxDqZA==
`protect END_PROTECTED
