`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tjDXfqQ4jzDDphtRwdyk9Y3y4pGaFiJhkcMSmQDHAUZtpXxTV5ADHuLxg/qVu8fa
4Am9P5OuoTvJr8xnTgh0+msE5kvvXHiWuFG/TMYU0yT9k5tZBpGRJ0kGmok46zXn
EqEJFQv4NZ96Tg6ymFEQ45ZEWr23HxxbNnOuHLxFRjZIyI9oiZydVl+M6NNbVpJH
KxL61DcXFtdvCtbrHQaWgPNz7BxPnEsgSKNVlmzIqiopbgjGdHk0ktKTeE/lTXuH
R92c+Xax2X3zlryOpV9fsd7omr03QWFdp1rVOQA7AdbB10hhKTjUavdr/Tx/4n6y
rNANQE8GB/y1LNk/c5IhUTEhRKYgo+gQx6N/us3srI15lztZjQSdXqDYiyhdglcI
5bpnHFU2oCTcdlwN26KWlhwsNzcw8pK9Kc8moz8vZp8m72eEvyOipEQZeN6SyKan
lF9DA7qudQGmELYBbJDK9UnmCziL1M4u/ZPolWCANo0=
`protect END_PROTECTED
