`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UInT363ZBSEzeZi85xURdXZwcnwP8OCo31BW6oBPCWsYB9QK8SPStwU6q+C4p1po
bDpTQBnUPN5ekRE/OizPf77DsbkeVBAA7PRWVpL3owNgkdJf7Po+eJJPsxfpb/4d
KejN8Sz1kHRmKwDsw4cQL8AzTqUC2ifBSL14ScYHZaEmCEESavxLI99ozlhO6pxE
IGlhsTO1JMKmv6Y1jPGFbCd/krFHjmQZo0jCD1VbAJr30wkPz6/SaXi2JIE42Aqv
+97WLY2c0eBSgiknJMoyjWH+hS9YouZMtWlFljz1pCX5T2DRo7LjV2nRWmdUyLu3
N+I8E0DAGeoPSM38Yy0BUDqmJYVpf316gKh/9TG4D6iTOPIBdU67nWVI0ehEQI+R
3Zzn/trjsFv+LXx4uqY3RsEaJKVWFvcbXh/7jSnuFFcmVw8VrQLb7DwjiBAU1Iv5
awEsH/1m4kkkDE4d4n3GjbhhyZDcWm4Tu0tiEKTQR9U7c2nGq71QGXGMNVK7oRh0
RVQziZBev6eUWSNvoRFa1g==
`protect END_PROTECTED
