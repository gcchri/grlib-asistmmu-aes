`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XwSk2nBj/rIM/u+dfnpPNSXgaANtSuyqBOJ9IUBkldy8FdvhTj8UYbQzjYUITn9/
9H9v79iwmPCdvH2EPURXOL/hwO35yqhELuS55jYdOwYqCAdMD8aosCbAi3YKcJ9S
Toyrq/1cS629mSXSGTn0qBuQRzqc4pvue8KpSQ6JA+AyFpBh+4m8Ec0GZQpn+F7g
RQl2RY9O+AYIoeaVI17yOJOmuPXJAy3g8MDUVMMrBFnIwHW4LB/6U8jeoP83P+8T
Y5dJeB9UmBnUtFG15j51JVTCaMGl0MYo86trRW9UYgs1XvrEpo2+qu98p6cQWncX
ZrnW9GU1fzh/RzxzxP3BZTEjtOuAzypK9tnFXod5jOmeJPNzOR0CIvwCwg/p0/dz
w7vf4yic2PjszNrmiUtnGlR/g3D0fV+0w8JUIhS/WZdwLVBFNISRfXOEqu8JstMS
Fi2dMC34dgazA05NMo0+iD0iTpSV0bcncGmNvLbQJJG1FPLXsaT19J1aHrcM9DGI
HYer8mCYmMLhWFo8oiXe7cSS0KdREDOONa8o9kc+8fAWLydfafz/BBoRwFeIPOTl
`protect END_PROTECTED
