`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thtPjnTQpV+e9io688cdeaW0l+EF1Wwv4y2ohljRtDjrbSGhIRQqhnDpaS5bg/ia
Z4tziC3hQm2eD+COuxcxQ1OD/JgvdqhMGKPK0sf/YqRRpJAAp6dd95C9CDCM+Wvl
3rr4j6rKomvvfJAR+hj4OJj1AhrvyworV6fHKL4WAkLvNqNJgLkc+tkwCcXflNOX
6Q9dMdjYz/W//iCLfwPXzjW81gUx+fX4theFvm6ijJpGmY1hCQ2HKxn2cS/RNz9O
8sG3ouRR7z3lhVv7jyDKBQ==
`protect END_PROTECTED
