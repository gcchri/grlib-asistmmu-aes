`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C80/1u4G79lVBty12aNsgXlQUEXIZ8O6zwDKTlx9MiE1k7QiVHTkWodMTNPOmWtC
j2T1E2Zb88O0MJEuVMKz5LN6SucbTDh9qpnw62VsaE6426XBv12meeLIFQS7ijIY
fcsD6vN9jE+wTi8vH8UIaJ+Dl1eswjDKdcv3ZwB5VXFjjQTvYAwVRnRs5biUF2p0
oPWlOblOXPgIBIbP1Z2l347LrnqnGCWZw6GBDc5vIb26kxHgknr/WU9dW5QWBxQG
dm96p81geSZM9ugE0j+dDS3RS75ljg1rELGFfQdCfco=
`protect END_PROTECTED
