`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mxMsMf9YunNVRbMiegraAp+xJT3dj5jjfKkvlPrOR3bNpSLj0MvJoD4K2z9/1b7w
TLJLUYia2DsJY65t79nwYPhDDwnT1dsqtkl9EHhrae1fHaweVK3E0VrV3jxVYFrF
mFU0J2F+SFtN8F2pf/Y2dcggp/E3LymgnIbM4SJieqQpKI6yRpzHqpUX55x/95fA
iRvqwnnLj9bdAYLo58WDD9iRo5xjg7qNLSv4z52+NdMG/uoJGpLh93K3EQf6rchs
RGFncdAxIVavMGIE5zhIu15p97wrqbIOsYq5McHO9eauvMJlO4hOkF5aOzUPdKqW
4Kdg5zHkRyRh7ytT83h/M+UYtwFvXnzqe6bFUK427kz8DgBAgnk+Bs09kYMqUcQa
341jKq9g0tZNg8jpVDYyLHO8GtOVaPQIzQR5J0k79j42EwfMD7gIedPV27p9J7h4
SkYTFBsmIf3NvCg+lRt8PFuS83Hm3uecQZWCqibOC3DfddhDnC49qS1AdPzAg3nf
+9D/Lj7ZJKjYO+bReEfrRPhYl25KqSEQruDoSU2d0/hUo77CSPS+XWKYOs7K2t2Z
nrLRcmNfuAp9+BKxsFfjZy1XkXMJFiT8GY0Qu+8t3W6C0vZKsNuPzXsJ59aSs0Dn
3zjvOrBis7FXTbHqDoItpw==
`protect END_PROTECTED
