`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZxZ0rzDuhSCLnGA54gMjz2JzOtrEz3BYns4T27ElEym2Hk3ImM8WCud8+VgidNwM
1IqD5XJ6cYAmVjtS7B0c+OOFx8KfO9F8+MZ+mG13ERkgRIYTRvtMOYFx+FXyF/mN
nt2V+W9LZn3dn1zW74MJg1vpMB/hLZbLPWjANmZ9Q/fXFfjSjPWawzu+Rn3WDQvV
+7DO/mKR86OxjNMRdXmBk7BookTccpFf542JEQgvSQRgJtCMRdG5VlP36T6Eg9fp
OawldEfRo0Z1nD/MQo0+wgqJywvHZNUlxtF1gRC1r5w=
`protect END_PROTECTED
