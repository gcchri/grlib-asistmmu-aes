`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Dco3N5r7OHi4fQXGIuurU17f72xK60Ac1tu0PqqMZ3GoXeKa/AZbyLDTYPKNAcC
kJ71KTfEUc9Js+RxkBi+6oZD77rZVhSpz+SpXRsIDhlbFUFcyu1CWzEFF+kHNDDt
Cc8+oQvQ+wOVw5WvbYb6hSHw2f2v9m/BAEpawfjCQO2xsZtWXCOeRpvXWAO4SySr
R68z7fQp2snKLzFGXm6nXcCkyVK64uzo3/IPxsAi4yE9RYjbdsLris1dyut6GNBp
RMUhv6J3ievA3dBMEZYHQyNh2htoAwKwZams1PCcBBK1+3cXj3NNr/kZc3wsBb2u
xTBMwjsvY7YatDBU/q8kM06q7TbgSrvnC/AvtHnnw19ykzC7hscNHkwo94EicH0u
4RoZKBhsergp94tBP8Q7g4Y8DSC67FdvESbn7PvQRSs=
`protect END_PROTECTED
