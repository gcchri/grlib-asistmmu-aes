`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5xxyyDUGq4XevvPqWVS1JDWKXWX2BfbGFCgMgFqcvDpZ8l8+yERl2/yvFB4ehu4T
eQQinK0vBMvrVvnloizBOhZEb6MV28F3ijNseFDfqRAOGdDdGlNeFHZfHp+sO7uD
dkxwHUTRhIY+eXOAXYho1x+4g4lZmUGfdmEM/+TM0hGnrx1BXsmkQ5y/7trrGtWc
C9+0JnXNLlU+01skSZKlJHFV5PNqR5AQ7G8l15WLdT4x+4zKPVldklqrhK/8xXXg
pDl9bS/QPFyvbXYS0cs+W9D6R8XulcQevNjA8nFlD0jRMhXNNV1zMFfPHRwCR+Ls
jDWIRSldYtHddYMpVaau61AiebuXMS4cMjgcyUIjLfxgObqaQabPJ4tGBwawwaPx
s15oJSnQ1Hg7LCQ5p+AmdD+5rAnV7wZjrsy9tIyXSVKVvEitewTI1JplBO2Ex43D
1NJnIVvUnZ7M9YfBRO4TaMUYwUKEbTN8IGZwXoWtqLPtNHwme/gN/SD1LjVkkH9u
pjUKtjA2tLsNpLBzfY1IVF2OjT3uRsha4aRfJTwPyUgSskV6Lx2jB0eCIik4a8dB
E9Z1aYZXnPf9wLVTTsaG2YqIpvPrth0VflQH2Wgrr38wQo7JsIrcAWI1s5F1DHQt
EuAmEji5x+LL5Uhn1qHZPg==
`protect END_PROTECTED
