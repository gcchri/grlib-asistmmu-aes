`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hKa3QcxJ7fDesRbMxqdmK11qL3QpUYKxT/i26SpbWMV+PNovu7HAM7cwe3d4DlsN
wt/KI+VPLLQKPw2jxCjIr5dwGGdhdpY5tPuxdVzhibu9qIzcxqcUZyqFO0a5mrA+
hOv8J71FTE4buGVSRrmLCz5qjA3PMrY1LKBK2aW048fZfe5GY5MC82uTrJxUcsM0
TRF5vA86IXsycKS2+Zva+YCe6f2tSMTe1friSLYonvT/svqI2gZcOMNBAXuKsnzO
cjEX9MCA0xT6z/xI1uDBHlwWEFMp1ofFb4wppQDV4HU0m7m0k510f2uS+NHfKrid
qq1j5IGZQM/E4DedUWjNm/1/VLZRWixaZluK8mJAAOYX3tOh3aQXWgRywz96jEs9
`protect END_PROTECTED
