`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GqWLSQ01Ck0GgmaSyx1WVU5PL1oRjNPTh+psY/XX5l/6rPcuAjlgproC2mYBX09
vleJc4l7hUFG7jmf0rS/1gtFlvRL0TqUX78mpLJoR1IuDKMpDwr1qDXy528ltCiZ
wKjZGYjeNbeSz16jnTRA7XO7Hz5qOkPcs+4C/kBmBy+M47KpeIDRZflpxFmS/dMS
oxEEUMLF3KJT+ReQeSL9bw+O9E0Ia8nJQno+qkEN3Xetxk4PiXySbgInyZOF5Asn
zSUxBtGwjaP90JVgy3YRhzw/fSYrilLyWdMWNTsrjpF5keIguBPaUdVbZ2/4hHV/
uJRxYJXcm/s+Jt6+p/RWXQ==
`protect END_PROTECTED
