`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DyGU0ta58UrIxVOTi4OATgRChKWXZomMxsTkfO8TlvO7wL6XJXjPoP29V+9dMaiG
0Wx0LH2l0GmNJr8V6zoEp/dLRVz2rm9twoMicbd7olsTWVCySPGrPQKHfp5TQOei
4nFttHoCJ1vxDeocPo+fM+cfCDfxOu1BjLiZu8M40Dcrn19cKBNOWNtkmazc3UnT
wa3TAuJxJZcgjZutkaAewn+teUTZDEEgTPAExpMkBmPIQr9CV57LudGsUfAjWG/Q
9hB5XGE3U5JOdDg6vcQRxFl2tRqJKjFKlaqP8doAQbgXZjXATS1oFVyCVbzVUCig
2fn9yqhCGG75cBQP5cr+eSDgbsWuD79OOkKHvZw2ZXbN3L8uH1fzJH70lazB29QB
1gCxGRrN6c8DIKVj1bz/26ec7dQN398q/6XOz3TjqsaDjbCFXmP58sWbrfD2g03m
7iADQufCu+fiFv7lYZjNDWz+TKm8ryhUV0v+paSWcxETGi7BSjJkJWTFqQzFYBHN
7UBh+ybfzlbo02+Q/GZ7YGdt3abfTCe+XxxCjNY1RqkwOTxUFURDwybzBtqFJE5p
Ez8I9XnEhM+0gHW2OKqnGRdL5JAozDAx9XaJNyMDwYhsP9yRdMrzXm2wtdSAf3ZO
yD6pTiHjM50sWZSFB9+c+Q==
`protect END_PROTECTED
