`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
riojUoNTcPKPzb/4AZi3ratywH511L0hWQdenOcFGaaCn2wWzCNeCd12XV0bN8Mt
pui+8JwGcXUETTvjL3m+nHoRwTcYutdGQbu3UimTKA+Ac2jToHxMCvU4KoThIlZM
ScH17Z2VEhIOcg/fL5zywgKealr1Gvd2FWuNRltkAet6uxSZDa/D52owmQ//j0UG
hnuEIWEWkUesPZZaXvFLxpxCOMOGkvicqqQINOdkvkAuMJ0dLZ9HaaHZuymUlg9L
8tGytqntiV4CSVBZ8NUq2kQ4H37gxb/6agmksJ+e552/+A9+WNZtB/bibDpXtlxB
XwozKp3eVCLzsWybjdZEJklJVQKTvZsEESOhz3GCGhUB7xJziKgrU9Nx498YWdVP
PTAsLC0vBGDZCZ3noXLKXF1YFUcDK0HNdmpHRtrLQKsk7EHdiMucSV5DF2ePaHtI
xrq7r1S4h8zDc5AjQHAw0MEnpSTVffttQ8aesAN9NA5C2w0KJHh9l6wwpbvgQtiU
uI//gWWtDoAX7XWJ+ajv6Er65TEXVi0B1JyRaIxJ2wptD/syStBFRPrL54ip18bP
2p89ptejiOhfcZJP0F881W+nTES6AkVW3sPc8z3AsSYGyv2liJ7jmniagSY7sAG9
dY8fmvOchxL/x4jfAfpJOCcaX3fqtElur4GSUayWk/A=
`protect END_PROTECTED
