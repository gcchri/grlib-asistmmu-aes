`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHjcEehuvgubLZ/6/nCM/4L2gSxhjR5naDYjeN1KEX2FY1ujDcqZebKjqW5u4cpd
bT6xLHeqcTct5JWjRpOdOUeGLtZoK4HQNJO3LT98Zob0LhtFTx1bGtAotNMUKE7I
KgE16EL7TPFTGM7xjCCs8EGKIs93WPENSQtGAGLwfp6S3hNgNx+HNVCflCirGuzV
6nl0dW5WekalS0sD21cTA74ed1kNQYiPslwpLFq08bjr38sHLsYyH9ZjFOgWvJvY
6NVG1rjjZoJO8Xr5XRUiIBP0OjSUYgzHZntKUMKmGDQ+gI3oJssLUzrZn7fnTyIr
E/BqZ72UwjL3Sk5Lv2m06K8xkW1C5fCbgkaRVKgiklp+TOKHX9YNkFh+5pQnzAfR
q3qGy5RQv04oT8EMgQwAkYkb+Mqinxc6m5ydl4GsDMTUsHnQ5bVTXMyY1umePpBX
KF0xXZDUpjH78P6mN3JU5014MymFZcRfRYX9hsoC8nU2QddGkmhBAIJ6EMwAX0ed
IinPq+KZrMHGN3gK2LE9yGpkKD8Ni/Bhq7A5D4hWKBWWcwN1ldDVQtw4Xmtu8OjM
t/coNifbp+q/yIR/tmuCBFStFDwM3O1Vg16FJ1izLIuCO25PuBNcu6/i/WMzamOi
ukabownzQxvQUfXNuR31W1fgiCYnCCiOm21yzyqb5a0ovMXQJFaEbs7u24I8XNt+
/+TUhhnXgJcDQUTDKMrSa1hX4sXJDYNNlZSyenRo8gRHUfpJ/2Hl6VcFDxY3v8Or
PxSltIY+GNkS5/oI7vAEwB9BkmhJR6VLP+KmkZRkGq3j0v+BEuSWt4EuFO5mPtFz
bFZVcDrzvs6/cXbdSZg4P6My4tegYzUEBg3v024wA74MNJ8EZ89ZWnEXQ3As+HpZ
aLcxhR7Tsm7uraXY65ERTLVPPkybd/a1ePtzOvt/lBM3B6RjvWGNAB2nBDY7mfEV
0ocGv5YzZxXZuJ4Oxk2lEbPcPyHgH6jvExZp+Wn4pT6s9ob68AsQN7fwtiDV24CV
ds21jOmABxX6bq3bUio2S3ugMrOMyICLoJA/M3zhFZ5o3Xr8mLQ5W2Yh5Mnv1HWO
FnAERxB/gDnu0OEzemYRzXhcM0bBOMLsimEL0cUknv8InxTxNnstqY96RCPhucU0
RJiv7/kH5jTrSOVJ03KLRk6n7Nym8ISJtE1vvBnLjd31iQA+5Ooihn2/u2lYhBWq
RorHch4aggeCG9XiCKg9xTu+wQYcKzOFXzPeMfA1qZSePMYSFwjh2oxJnd1Co0EF
Bz/WtJmJr2DqcefhW1AnXzSvNGPPHnJjVQOzAcRbLEk4WeCWDEcvlDubMQ5pr6TS
eCCcLYQSBnxj2ksKnkuztjWXOvd7BTpFrW8wX4smMUNG6w/MrroQUIIM266gbG0j
YM2ZMZseRYT0/+fQ0wScL6DM8Nvj+Tn+/G0ZngYfK0nV0nY14fOcpmDvXviu9L4b
vgYfw9EP2gOrg/K3hJRW1tU54I/VK1CkW5grWqUDfNsRMpacPvUj97SZp5Lp2ytW
V4FRyFkULtoG+IkuBPvkeVjfk+Hxv8Gf/a7s5ze4fmMSf1zkuPq94OW7A1EBUp7z
oL+PFx3jEGDB1iCwTMwYykiruscXONjJgG1tP31y3gDNGEywUXEkYGvMIGOGTPNV
wX5Mw0qbNZW/0rl9TTM7n/H023fvbQhH6es6xwlFesQCV6n/rqcsie0FGkfEvB+r
NVuESeIGMmHYXAc9pkEA/tdx97VV/93RgpX5Oi/XnfPwLxmoTJq/lCCenepsy4yI
kIsqmQhxlfhfvt8XFkRn0BuWFMatjrd7/gwa5vrq/PfSuBevWHo2iTNt4qwo73xN
sN08wb86qs+jBwWErPk4PdysyJCpGU/nTV/o5zPVNrClk6YFminayBzJrdI6zUBZ
u6PCqR+eVuxk4mHw9kP21TLrpjTTfBNjfHR8iJi8peDniTZJS3UlOgN9gZv7gKQc
5X7C7KjGKm5gl17LOOEvL0M/ijvjV8cT6OR2zWBI196LVKb+qlKAI0P5LSAkNX6w
phiLHzaIhU7RFFxok+/CqhyHwJB/7Z0maCUWVsA0CQXftCgz6uN7Lg1oOo5YhB7a
4KI9pLbiEIV8g5QGJLdXwQLYTEh8EVaL9wDHiF0q9q5dmx2G/DLTgU21Dc/ySq3D
sz1vyvRVdegztGcvz5pLDlt+0TfoYihed7GEuDNBiKld9PIdd7in/xGzGG0fkirg
pg7NO814MwlL4Z+FndCt3Ktm3E/oAbUp1ByqZgV1m+lior2nhCpcC4/rE5/7EdSy
2yxeVY57LVMLro6t9V99sSoM760diYm+XCpcu3FQA8pTXjOA8xuF5BvYK3cBZCJC
+BSTdXJhP2/Hs8ptP2x4Qpef1uh1U9myG5zApFn+A9EkN47/T+YSecpk62gKIW6g
ARSUgnAzXL2l5ywltVCaF54YyotiT4gSDYMOY3y76tOKgaRpeyb6gz9LdU8bXrsF
11xuAgOZKKIlKI+f6PXijUGnuXfqAdeeUv2R5y6w0Vgo+0uV3ZzyR5FVU65tKliW
ja2ay0DdTrZZ0fxG4RvG/XKqXc4zrfhYuNc+UDDJC1GZCizszCW38EWs8CXedm9O
HWBtdMBSpzEc46KJ0h+A/pqHDiphxvGS/gAwX6bF8jjbQLnvdL62C3jyz30DZOok
zu0qLh/P0hSfp6dtkrm6zz8//69bMjB7jaTUGLkCXPpr7g+uVrS8nT/cBgy4LWPr
ceOs5M7Nn4yNqW7WNNcUO0cKBSeTK1tulmVjvu6u3JjmaDcNxPn5A/FyjqFC8zd7
BQfOE1xICWtnkWPIUItJG3IdzL8e3lLE9ocV3uHh/xHomtHxPJoc1xbka/fiq+A4
Prw3LAtJ3BP7OQ7t95NgByuWMmTK4SBzrL2Avef4JvW7NH1mqddRlO9aH7vA4UxL
uhg9E98yHCEj5Vy/DSRu3sS/TXsTMDTyr1UQotlweXABLFuFJWl2odg9jC37xlvw
FidCcXp5/GS3r/Ys01O1gXWgZP9Q3jlqxf/Yr2fifQM4ocjBzoNpgMTbi59RlAkW
ULkTUZ7SaOAL/GranT+Fr8Hz1w3sdwQ9yEEH5fCMYCE5xxIY9wIYj4L5DmtLxI9f
Q3Xo943MwGpfNEYh/StroacW1IJyqru7OPv05RCTSPCY2z6v+cGMwF8ag9Pv6kZp
/Of328IFNlbrNLRfNsHqNOxYsyetApKXfD1PZyFI2RMXbuEfQX6VbWg+XwgI1ZQQ
0gHU6XzgHBwXBWrJIWgtp5JEu0naYOSYVR2mylg46Fy8EQX614gmSlIq7z5e5W2A
jaAZ9KjOVTSSENH6I/7PmEFSNTWyfOT+2YnvXTKuFdpGpA0DyVq8D1Uznmq5e/jZ
KE6LkpJoJZH7H0oYO1wi1FyaDufnEWciwG1H5NYKl3BBdL+mxi0q2mCTIg+El2oh
JR2S6c1BJx1Dg8BafDy3zkxWqoDIY8m8xn+NRGLkyB52IS5DNwDqnFchCktkHf44
ottpRzOKnh4SrFGP7mGXS0TUwH4tiZQoT9rRvoxuQwmCN0wjxhlCFxZxbmvjic8Q
K0V8R17sR1hTCiGHVhPLvoVEYj8yiBpSXnGVp7Z4avnpViFL2Fb9a2SLn2HyujFv
p5UbHpA6sJCjlETDCb1WSI5Hi+5Lqmhx1rBc7+NlwOTetwNMG1o6WomUZkNMff1r
Q0FZDT/T/UmtwnFWKtg48BjzES9J4Rmv1qqA8vZrwLttFKIq+BqRieg+ys+1fMMr
1veRaC9QBDip8qAxQ97qgzsIHKTBPC/KA9ZBeE2LvpqQKNMmcVhq8SBMoSS+kntW
S6laKFAC7Kjbodpg5vEWjcnex/aH4xxV3D6ukEj0hpfSbxaNfJTQmb/NwFh3PxHf
LHq0r2UmOYBq/R2g8dq/N0p4gPk0aE4MHmD2SEgOPgi6AzH2MPONmlj/C/VkeQ1w
/GynfpXFpVAeESX7xiARzu+3wOwbsjSffuKGI6x4bYjIL2EILcpw5gZTQh8HUFeX
vTe74k6TvdAgxf7ldnwj1/1GQ9UkmkB2R3+hRq3RQDfizdlid+m6A86lzPermDRX
3y5D/u+D10zt5qEtUWSwmtZnuwn9ri0nDgqBpt6uAPwbw7hr0yml1y6MbcHyt+AX
0T0XOkNuqXqkQd3713XkbzAh0R8G5/vlX9uy1Mnik8x1wJnvCZ00CSTBDoMU3sOu
KeuqjNAhCLtxKmAXu07ScZgkDJ/gwnsYAOmyNL67dg84qlizInJ7kMkyeOIjOpn5
si2obzvgDKrGkPUSx/sSB5JWmI8atauiFACOK8luTX4B2VMCKvTbzouISYP4Z1HM
HSSy2zZ6RVE3chaR2gj1+QBccgiDOlZ4ilLcyFoAhc3XJLX2IZFfXuj67iLsXXZl
u6ScZE2y+mF505pIQpL/fJGQoMWCyf8wS2HXShyWMMgW9ZhktJd3oDPSlFWYgKiR
ala5WyJCwbXzPIglRYpKt+oWgXQXTy1QJy6lSgfPsZ2pDkTFRULIdreuwG9aiwIB
`protect END_PROTECTED
