`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j5v/RLGQ4zDB0j2ZhdbFTUVOAs2kCag1rrZE45S1iOlX7DxA4Qa7v+d3SsFUN0I3
xv+YunJZsI02EdehMIX5QMpdI1HvRgEfDGkB1MbjqGJwp3HtQWrTnl/zw0wbbMlE
JzSMe6oMjutXJBRTykAopu1ztQ0MXsSwoZN3Niego0YrYHFTmTnE9niWe1YA+0Pr
0793E3MaRhuIwXwNWYWupvhyom1kjgKk7AAQdJuN98KM+zl78GnRW6jaHsP21wPe
AGw/rWsV54KGMNvR7CHf7VNyBCgzYogmMSjSGEYw0/P07FLMMdCPSkSGnJqHWhfS
haLjvq8pAtg2XGwjfWA9lPzD4pZjzLZ01mKv/PZQqrNHLTSYuhDPZilJtgxpYm5C
/NT2tohJAZRJMl1VJxABybGfTihrC0S+XLjCR1OjtnZqTKwsrJ8kA/bmug0OtweD
bk96+99Jckt/ZYTYJ8kY56X0mcWGasW/MY8c9XAJPdjWffktRd9u6vPj2uufddIz
BkApdIkeEYXr9UsdLzq/LWIAWaQigTP78SKU7IDnql5e83Ki8DpaXb2Kcptujtrn
256yW3MCWHOpzHi28zQPq0hUPdmXalAMMcPccvMvDegWtTWW7w33nOcEGuVGetKN
nV1U0peAHXlTztZh8ExwYGDt9D1YI/zahGsHzSkiO4QMvVRfp8JtQFH/isYnoqlh
`protect END_PROTECTED
