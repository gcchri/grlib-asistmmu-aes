`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxRwsm+YBlDGCQHwuDcE63C/JyN51d85AtWCPorab05aZo91ReDgPTt/UHca8z4n
pYYD+2qNOW+G0hxjN88jMOsAc3cC4j5ppZ53Ij4LkOnDOEom2DUkX+Tmhmtp7rxA
IYK/kyOpkkMHsUtQY/va+xTr9ZAee7jkHjNNcK2964yQsOPSmFDoCK+jpvMJodhJ
/vl1CvJ0b9TXjY+jb+8uNYoGi0iNGur6LvCWLiWI9nDzkq4X1HwAxqoNgYEWhkDw
b7ft3ukrgVedT2Ajs8etpXIP0qrcwfz5lc/gBKQAM9B6dbvzkRjnJnCDk0YpKXHt
i+98yYzGKnBOGrjfn6QSbC7wP34ZrP/Fm+1aslDFePgmhB2+0GQfJ+goP6PwR2NU
YWP6VVxJZIg+PpMFW9yV12qj5a0xkmyEyJL+ehSQpL5a/fEEY5lv/7ghvqtzcY/Q
PMqCzchNiw+Zl2ptKY5zoXdA/GLO9fBz5KkS9OdM30XBl0XcEdGGkHkoMj3SMcVD
5e2RnuH4kKxrdVEOKQC8xtzhapjDDiGCyDJaPZmaZ1rg9NuvgoEZ3KrNe5gJBFxZ
AvNOEQeMn/Uu5KYNkpDMRi1mF9iXrcTuFdVyJE6yKIUQHIcex7CbV1sdHjlKyNgi
3OKkYU3DM5KUEJFxKck1z5Lf/Ot4VrkVtsICMZ8u8CTzMM6/g8+ETi6YEM8CBoB2
h1/4VBxvcN/Zoo38B7LnKw==
`protect END_PROTECTED
