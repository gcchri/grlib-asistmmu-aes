`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNiWFtEoRh/3BjgMHOadWNzklenA7olMpfZdxN11ZqP2NE8teCNziI80HXVWUvax
G0ofPIq+kpLKBVq7qb8fBdF9xbelygXlSQbQYcMR2H6+Nud2H3TBdgIcyw3+YXer
n/gPh6uhcoGov4smx1nm/ei50jcrnhyPx1yJjyoBZh23w74BIRjyGbfmz29984XV
ANnrC6G/r7vUFOfHuONJby3DWsghXKSMStC1Wr8Ifx9N+fn3euEnIckb3dcTXYzr
wywSXQO2ubVl618ur2yWUh6gJNLXxTDD17RY6L6wq2Yi0VsrAtLUBHsb9Oo+emfS
Bpn8o5ILvimeYj1gTARlA97Nak0nzlB3Zp6jpWnLo33hcsbBW0m0LNqx1Hl/6LYf
xH5BM7UN7ea+Tw5eB+HUDh7dwZe445Om44O/NrTgOaFYuXT46n1JQ8TKn3v5t6Vp
YXvIQcfx97bCjf7T30uSqrX+eYpB1gM9+ug/1XsajhIhSbnU96vfrVg1jJLNO0WD
ybn81eJhc3hTIZ/6FxnogCVF9vG6XywngUMjGLr2NwIA49Zwpk5utViMGzqr71rM
E+dJPV3tzNtFXZCheyi4K5jRGFb+CfFK7bm/oauWoAw7ljkPyluY2I6FM+fD15V3
JBB81gPyvKL+KjhlG19KL/rKdm5TKhwtfzeZ6yp7HAFk8Bz+Zo+vym1jQZoPpn85
VvlXtjOs+rLXjNO+cJJZuIPhvGP3X5CXO4RvBQPwEPhVlgM10SVoS4E4hNHMuG45
rVoMCir7Com1+8/LtMooWRYYGoyM3CPMEMq8qmiaFNxS9ZWzucgz7qrlmqodwhA7
Zs/0oVGd7gh0VhbgecmOp7Zn4D5aBeyWrYEtzNt/wbLujvtfxD2uGtcXkD609pJn
LgZXqrG1IuEI20xKRt91TGNSlm8WttZdNmk7p6Ib8apP4tPpm4s2zw1+/IGWSHRY
L6UccbHnaU65r2/xGwGa0BJw8JxD3Tb32u/vdFXy361vsRsa+wsSoo3HQCyhVnFr
vBgRjXnW8AxUHnFiv4BHEeHq/86brzhSgRhuZlKBnbETbO5RroE/uF4FXDvfYndW
u7CFW/ztCWpUewuVhTHwBu/0Sro05zp+mh2VMyTvObw6FIkIuAQzrbS9jCnPshSf
+XwMFDoWynsZPhrgQU0kK6Zr+s0UPblZODLlybEC0hvV01p9cl0dFTzknCwVDt/P
ggsjy1DZyJ0H7aCUSsM03j/230pnItYn0MPSiesCJzuiyhNB5ZcdpgT39P3z1wBw
V3R3buuAy77d0eB81Ami57k6im7w1lMqiSaE0lmXEM5j/8M+MO5f/WsC81Huet/s
DqqrivEk4UQbASfqEP6eb+J4bUAstCiWqxdlikO2AmX1YKPCw8VRQlV2enR4fRm9
NNe3W7jBHqi5i83mCERQguiL30kHRH1li9u32hKrnWQjQXBaSMSFm4aw3Le5fq5s
PMY9r82CTKGDtBNUx0teEVv4VSvoZfQvyARQB4qK2LHXNKz6JL72xXIyOT8vQGLY
27n2j+p3/efFq9KM1Nn4cGkuU4sV4AyKX3orySqCrrg6oS2AQpr85HvKsU2XWwCQ
l4C6ex9geTdKUvpp3q6LEKe8F3VeCoR6mGMc/WE76g4+LbWW3dygPh5VwKL9c0nd
/r+l3JYg5mbHNURL+l6mZB1kuY5DqgH7+/7x1MWRlv17TSGUhy2U1OvYOLkLsTDb
ZRZ3Ne6jYy5o7JaPQZhKLDa4mjYKGn5Rfh2uk6vfpEfxr3m6ojvewA1wXr+/XrH5
qYXIdJpDHe84sPh80ULwGymL/lpuQqvan+OFo3bd/yAqDDmUOiaGDuaqS+5bdBjA
dEpBJgt+vFQr8oRNoQ6l4vB1q7eP86MRQ+MFYyPPasHpD2GSeez6EhcEIRmFT27J
6mlLq7JZdS9wfVkBek0tM9Urb5VSyihwX6UCJUYnb8B0Aw0SkBlqtkobbc+4FfY7
z7KNK45iCobiEEasPWNkjzbGb9hC9SAvEmGRDkRXgaMlNXZQU/mcd81KDG0cr7k7
ES+/wkqPajsZ2b7+e6uVulodJLIIKGcRyMFVbVGsoVnuHgHPzzvsUzez78nVs9Tf
DuLDZfif47WO60tA3SdbI7m+gwrjaYI2IsSaJvr9e1hktBMSHBfKxoKaTDcmv0EM
fjvkE9zZuXdYldkIfOSa6ArOaOB3nEQAquXtTTiV8qJCeRslx1C5YM1nWUi6ljQi
DwGZ3mgpRDbYuE2TNrF/RTkvBTvvs+zZoR+9azJ3HGOYRY3vHPsMmDgm203cv3Co
2ymL6qxCgylAFbd6qqVdzFV8sRnv4JHcxspNIivXH9FLGcjKgXNsQNwHXuoFHQ6e
iB3VeckRQXOByTBNEw4gCj7B/WjPsKia/CiyIGbljYJ7lZGIgVkyMtwXkS/fieRL
hOKVDz/XTsH5F+w6eus+H+92wzkTW87FurG7asL850REGNPr/olDfBc1XmT8cIgs
cI3u5XUCN1sD/3Qwmh23kSxsUPzc5AmAEz7mDOCLXQFY8p6exa2kaR6p+bVV+oiU
Drui57DEwJTw+vbba1Wdjo2IABrfyJ6K6oqaiSVZUVUxLQvOkHPNkqb/9QHPv36Q
qVKqhXPaqEb2OLLEQYoWBqBuw0x/mV5ZaCwZ1QdADZnh/F9w4hrzXOjIhfm93ZYj
ubceeij4sfJH/iofAVig6g4iiBWBiXN9Vx//jLmk6cz1LY0GwrJYPFGAm1LCM9bm
PHGEC/L115lHEjfGSVmMxNHVo2LS3KsDGe8fe16X5Rkci8fJjV5CnP8kpJQ/VR8O
xJuNZGJZbyER3nGiL3LzYcd5MCBGd6+jUxDH8DqXVaOScLUoy6UvlLNzl4XELyk6
3OtZDSulCVxb/1Xpph59uOh2aVz6xaUZ904xzNaoor4QEo0XqBIU24lJkpfZY15W
OltI8hvkOiK4ZGCsh/ow2Z59PWIV1G1Q4NyQrkmhUcnR+NUKow4o6W+4Xev6GimB
pQGjH3EGi2bMXo65WFzgzQuGxJTz68biHB6sQime32tXPFbr+Vu0QYojmzby5gk2
+hpO9kFqscr24HOZSu7ggPrFijZvGuGobSBiK0hoju8RS02Kl86n/kaas7dLGOk4
D0TgivBsa1xyXO0kv+milXOSpkV01akBW6fgH0EUs1Q06eVt2026TlDXufngz+YH
/1QMprgVCjLkqxEArCi9HCz6Hiu6eBeDPTK/GQnSVyotzFdl/BQjNvjWzFA1IV+e
DhsLZpdJMWhBAFcRW6pi589iz0S/JU4KncAOCUtIv7WhJw4DeCC3kyQ/WnZkTxJd
UKMml67pXms846i21oIfpxeji3D8rok99kiC6UYB1EGHbj0dWirk/YaesaQBmHEx
lWdHXEATtFWWHfs3Cv4AaPo+ZrZZcLDxxppC39m+6NLVgCRW4AVfyeSUjirxWN+Y
AlQLRPCNc72pQZ5SgB8+sgXL3F1ZqfRU3LoJdxrM61Z+BrHPRDNvppB5JRtJxdYQ
ic7qrt/zmIbQyOtQ7OD3DTm1GgGEma6BS/Jx4yWqj2AIbaB9szOyYbDySwjNKw6s
ZOgITH66kF0twSn5DgiqcRantxmL5Sy4xvtRXNCQcdlRalsRb67rbNPL4OT/Kx5T
ZrDFuvdmJAt4CwHc7ei/hTWCuYbzISnhYmw+hx/GMPecLcm+pVj4ERxsvgwpZS5O
zuWbQ6afNw+M3djeipYMvtaKG2FxwBo0gal8FsQJclhJfjiUdbD1mmN0T7LTkPhB
hAvy3F08tXSy4ioqxToM4Lpd+CyxagEt1Val9pJsbwHmcrSfnYSwkMvWVDAI33D4
G/5eDf2cNY19py9Tdp/d99cRrglFXkiUG/XbyzdjT3LpILoVzwI4sTjuK6Jzp/lr
m5kKXizOBybGDpz+qXWVMITzRHc2oOBdjpYb9GRj0xTG/Z4CKeqyCzPjByEF/arO
zDD+I4g6QQTNUboHnEHbq8CZomJtcFMOAk715mHlgTHSS0TQVyLCi/jIGgnU/Qy5
8NKBhuSAN+s6cKGV5HOYu1x0e2P7vh87w27RiPoXC35vuTNBhJlXevV60BZWtwWJ
VR+lCE7wf4YEA2Z4LwYpn103/+adOLrAaXQfF8tWLcGb+ZmF6TV8GZ7HyZCusZfv
n2fg1B46NGO+qSRxXB7ppBOBAdrbHF0wi82xhQKXCwLwPqwVScBYjHkLCOkNGC39
FKJKJNVJjaYWfui3LLl+mu4gz1etrIXD0DLu94VPhNSq99gHQ2XwsYLFvX3PWHSs
ZDpUWEmiPuyHvhU7c1LhdKiHDMhhYLNjaAioa+fFUvEPVe+I0kwSdFVriJ640S/v
vfZZsixW1XkmIAHNfFT6tyvmExta+BryUdwa3BMU4+x4wNMIfRbvLwcXfppuT/rG
7L93+Etypr2WiYp/rZ2tMZbC4nT1Ge5hrweYEoqbwdrEMvuxtYKu46jt7IAedm3P
HJj8SaTWmU/ugzS1OS4N15msTgGKVFYEVJ2jMRB4nhLNLbOm42hzT3ONpimi/NSi
K6BCp3z29jXyDy49swBx/6AGlptM4u3jGR67TwYJkZZVMXWg7OLJ3L2ZdACyE5O+
cP9Zk76d5RYysaZJJBmTNV0UtZB23ZXRQawu8zM9D0VmH7sgE3v7Iyl6clOmQE/5
kLYj0CWYH4kBhpSCMLQdqTVSNZqwMvgF5EK75QssiT/96ljPTRjhYU0jyp+F58eL
zFicBEQ+HRtB8zcrOv0LJ/yFDhGf91uY0VZNGGI64sjeVKHv1fwNr3iuNUNAb/UU
uSseE9PwyTW16Wos8qKfy61UMkBkcpgnNIk5dmtu9TBxdYuoOlpU6QlLGYzwEzvY
Iu54Fvk9RLC1A2Q5hGCTW0D4NsvaLsZvUWoE+bdjkgH92TweTvd47MueWoLyr/4M
DCMp+nJ+XNygAvM5T4cYhZHDzpVV9g5nVE3laBBcwh6nwvVfISOvI9IuUzDwMy05
tM9nS2Rj/Slx6rkpzWAFlo9anQ5hbTlDhYlqO8+B6WslYpTt9tPdyE0CnUQ26Xpf
2Ml/C6rTIFtUo3/FbEM76cSVOxWlE00wssNJ5fCRf73HqIZWTylLjaLv78vEsFmj
kXHEUpJOaqS/caj5cr4zZ9XD1KiVwjG7k8TMwx9Qdgd0YYl8f3uLRwpnxRCEjvH5
Hf2pL9hqBWj8OX6QlXxlcTp1/Ym411D9FhNydugjdzOvqN6isIRhHAEs904NiTQx
vZiughlKfO2/gsD/pvXftNY6GgMdayZFW+6TG/Rs/Z4EqSCSTXGbvnZ/bGnu+pVm
fe2sQoYuJUkxWIiiuhcWJI+MUZtRwgAnVdoc3qDikUxwr32vXwGZ3S8Px6mH0/PU
rXDLM6+gCKPwjgr6QdHRvZ3cClf37UWDky+AjZbAP7We3JXNNFY7txuc3PL7h8FK
zPmBaJ3ZV6QvSbTwPoKKjTDvDUL/SEao+O5lAWnFFT9jmFCbT0LXDbKkqiWfPm7b
2uAPpIrkqubDF8fXmZWmqIipgtLeZrvLJajov9yGDbeA+TCZCohmTOpob3T8p6/o
ysh1zt5ryWp7ly7OWf/myyLKL7GlAyU5xJvosRPqH6/Gq7t2Da/u0Q0jIxqvM8mg
lndQ9Bj01q5ZrrCqG3GckWaDBItN9DW5zXs/cJP1zqP+ziznQZnRonBQqDnXk8Cg
sCT8pV1m8qU9zenJtRJwFOL+t+PPo4TY2d8bxkB1/gCRO6j+0HSN/Ov432uGDg+/
/6iSyXQB1VFLQAg2XwkZrVH/qToGUT2kLAqlxT0RCWoUzyn+dzapz9vIYp53HRpd
YEtuLqo8AdbLa8heeWb8MYpQu1/Zi31bv429ugfsLQtykxjz7+QJpROn7gSrzRth
VtwS7GypC/N7TuvU1uS9u/6ZztFLqsroOAbBJbLhhwJxR4jndh6hhEjx3WvSMga+
9rODhmuNyXaDn5d195I+2MF3/+yC/n7y5b9ERbuh1wilJvD1AZsMtBF5csS5gHHc
rG2NfRR7cekk5R9zU+zIdW3QqNs2DREVfGv6zXpYCBzAXQnH3E5Rsfj+CuPYU5Hy
VdNnVqapPCEEkPutzhwWukzpUhPVjxgBrAX/vmrn8g18Sk1ruiLqn5dgksVUzB5V
EDCK6JTwt4GgVbUjxfS3jaIACJLsHIUqlgenlL4OqLM7NwJh/otfOrmmBkMAapFO
vm/Hv/2lXr9mmFI0Ct9vL8v7pQKZ/rPB+p1s8iwgBXlP907drUbrgJyocR3VidlC
mRkWZ0VYoGEjVo1SLtHvsU6hwdmBm4r2l3AzM38j/lr2wzNpX+zm6fEawuyN9gPv
PnX6bOHdk+A1YzZrseebyYzarxGYKeQX1SeA02/J1cJbpYssvbcXSj5gogOJDPMm
ruhFiHWX6Qk3O0Ol5QxCSElhjB1mtdJtIY1tvNtw1Vmrngi0mhB/8HAkH93UTYVV
B18wzEk10UxqnxZjAyK+YEFf3gwd1Ned8DhnkgdZQFWE0TVo2yvSbfa6Ex54XTl6
JlQPeclcbRP1pfC91NBWZuVxVX/RmbT9DhjgawUWT8yOXBiRAicZ7A6MN3ngWw4c
liX7yVUDMH2VwNRS3Kp7Y8o53S/vuP/bY7C4Fb+kfcZ3FeWpyl6QRE1SsgWQSsGv
M3jn8opLRJqToeGDdsHuBaZqEgRcuVQNtECuXrvueu4bFdPhtL58KPm8adWy1guU
GOGdbIUcDHbnRbZR/CIdtE1qgwTa7gY3IpIHAQZuzGivIl7ass58+NFB3KfMV6mb
fTBsSdZ3gZuFEt0c6L5rM7GhnEIKvqSRf5J8J/lmznW6T5dySe5ndKf005YUE0rU
e5Dtqda7LCnRdKarWXNuvmgXnwl0LoIzGLSta+Z7A/vnG94yew26s9uncEiGCnzw
Tt72KMePbn/0mH40K1hgpDUe+6uU3KFv+hCNZ/GQn+uuf+4MLqL2NfsvRbp5q9s6
AJZmshc3Pb9ELFGMxIS+0zOREC+Ymi+DPXJB7Pm+6TbxQrY5SW1G2eageVak7wuA
gfRmXw53qmHszJ5sDOoQ/vLyefWG6g8IWR6dMUFkDTEmLodiVI+hOOWMB/1H8EsB
A/uieIhD108tHb4AFLxUloEDxA3f9aY1IeRwBTriFOpcaV7Q06ozxlI8fobkl38g
Lx2hPMkHQtRQEdLMWIzfJfUOP2gUiA5P2CSEBODm03IMsfO28TnrTZzZPMleK0AN
sOKmjS5LRg3xiAHo0RfyAIGnJz+e6AVKPk1kh7w/4IhhCbUw3vz+qqZhT53QdvPA
LohgtunCMnfxKK8mPuA1l/YObXmkflkV/G8Hcc2bdCwMfWx6bLlV/kwBeJqpiFJR
4+yNBMGyRhG8gWtxXSOBndXX3CU5QHWfODF8Ghrlm1Or5nip65IYwBa6RThW8mYJ
/lLapGAqfxBfhNYJIgobiEhqiA40xbkscZ3Qf26RHNpxcI+dn3kZZbHqdTISGYit
KKuuzha9bpl5AsRr+ILZDmbAZO9peQRa87BLsBDmTBDovX21NoZquFatki1QJMhZ
Yj0B3bwrowXQ/GfCcAs0CEInuKcmrpX6jNApYIr70fSw36rUcTaE84VNShgz11uj
UAxzaeTz6a+/8w2XtQRwxgB98/tzQf6oTeFhvliujyat2JaubsR+kBdRqKAw8ruw
M82539TCw7O0jtpoVKHMtV8+lGKgC/AbC2mpdNmfx3tf3Ahj6LNkbBaP6/ZkA0I9
TjC4cUy8TqlkQK1MfRBHKOyDUq1OrT1q3z5yWMiR2ywku+W6827qAh6pltpyDtad
SUclLM+HAFUQzIjnDZ9JMyYzMCM6qtL4Pyo1eNmENfXpCS9NmlaXuLPeSWCPuTl5
xSJRj08jfE/bCQkUERledOJqAk9aGBxJvBODG36KFhAO4yR3SabnpBNaqQs5RMTW
dMUetRljoG+wyE61MwYcm14MiVlgtey5gUjsT645neNLsEG9XIr0RkNmRECQjkzy
anhlQShsxLFLLSUQZMThAuD4TDYwfdxWrWU+tU6sVC1i8LBFSahOJVNKSszJflIB
S9AwdIM0zYK56pQscR5pKrX8D3ekhZUtUcnfivAX/rbgwsWQd1Hp31lg9nPpZHuK
xJ5f3Y7O3CDz0zpcq9boP01QMli2i370lxm9rsXFDESumsUiCBafDz9G26aUXs0q
cKOYeq+pMLiPQxqoZYm6OfeObbxS34zh6YPVQIo4g3DtgCLi+OuvVlXp/F0h0zut
03KdzE3BP9+fvXlvAJOcxqY30X4LW6Hx0bK5vPEYCNPQbMoIf3K6B0arpskpmXyo
vtG3bZOUiRcRoTLpbG+M+kA/90ORY/ObO8C5cxpj4NU29WcOuMiFn401j5RhhHBV
mDvMA8P2dymp3J3asZDci0K2Ip2O4CCiAFqUmGceQ4OattjKUfBwJ4nhEH0O+piU
DwZgeiWTgqO8jwQJ200a0Y4SBifkHwShCivDsGhavAGBAZQqiwqfMzXjCR2BWk7P
jcXBCWvF4S94C+1JWIxbhsdjJpyBVABeDQ9r+ITXBJCwYDcJBiiqtbu9YJAdheU1
Qdn3clU2osL7TCbNRfprbqV+kmoseVyolbcYCM7st9wajccTJxCo5yRqeW+73TDG
/fuX4ZvpR6MI8bAby6oy16/0GAOGgseu5BytM9LPwHSZ4qf+BH3U3L9XDuNODyNI
GDWXZMzxAbg6mKJ+Knc5CNYS52lwwZi5mmRPM3ZIXXxKnBx/jv3wPvkr5aqrBDnb
wGZYEwAqfFW8CqbXpCvl+zz7ENQEazraUsnrEtzQhmA6j5OdVrFZLwQeEUGD7DIT
cGXqOuCZHtbwXHPj5Z8Ar2Q+oXdpwTh5mk4x7Osj28GGNrXHFEUBd46+FZnNxEHB
GSdfV9yMnJFyp/cQdWgPDHZ+YVqDPvrvH51CcPB7znP25QapIeAjWfhE8FhZIe0y
TJhXlCiVCFjw9k/i4vHGsMjCk+tP9tU3tLk5zUpSn3UQpDndbouIFqioHLGyPSmL
oBzQpcnbB7Gcf1VRNQmaJ8dvdpRG7D908wUNrGIWsnX2o7Vgrg6tNGVU84c1teuz
QgYV3aflFlc6PiYmBQ41FvZuHaFE2z8FWOuG0MaLTp+jjKeXs+c+DWWsqNyZ8Hlu
+A2NeZ6JCXA0QjZVaTS6XGKENGbINfrFZQUbp/7dxWXPUzTgcpB76WNridY6LfXL
rcDmr1mC6KgFgg68nvFkj/KHv8B51/mLkPdu+ZCTfD6Jh3v6Ro9Rtlj3ubQTsMhk
DOex199KidA1qi1WNt0DGmwb+Nw87G4T/OrXJvcA5IrFaPNS8g0Czv4XFmYeBa/j
DdxvMqgCVRItBMojPnbOi0kiEK55Y04X0Dd6bvawhJzqjcN7JDrcvhVWFqgXLSc7
jHU+XYrNVEAmcKmpLgw2TSEZStecUp7BktIxQtGHmwxyvQxS54GOoa4vtxec22nL
4BW40Np/fx158dyXY2JXNV5gq/+e4rlxRizgkPDAJTdrWnz5eNoQWi040DqEg1J5
6X3u9OmTxWPawme8SUpOCPWCDI4MH3YCjcW0vdnI3f0vjRmymgiy5k9qoMblOK8L
nsBwbvLttzdeS1hpAif8sSsupkFkZ1tiveiMUWtr0wxh0E0M9ybwvE5JJYYK8jDT
iN5pqkv1vm1KUty6uMkxlLvyhOgA7LP1FZdDdx7X3yiQIfTYykGVGWvPPfiovpyH
gGW4OVBEILyxMlr3iEzJRZsil1yNGwRghCQ/18SijGRQsGEfKeLPNDkbQuRQhMiL
Yl+kovDXBl6UaclgnVo3PPhBSDXbg8nv2eTesmbWHs6cH/m1YiPXichnUQ/lgaLc
5dm3z/zGv+Ows5SMoq+yG+BziRjGZjP0mOoTO86wJh8EE5hwjr9h76z6WKG/637E
AgSJ7B+RrjIZ8fSK8PiywWaDHRGL2maAuleBpP9rer//RQ/uuaEG6KrIC24GZT7W
hnApYNw7YWQVIyTDY3zraM5zl6GUNyUCn46HHncJhw7UU+bFjF8WvZZ2Lp0WF18M
+pZARQykaDvz2pUaIJXcm5ODN+hb5fx1tAiDexzelEEazQQV6jfaQtRRVF9wzmCR
OD5PQ1sQQbdRZ3WYv4sp4NXIIIpmAEwVqBdNL/9lG+AbZEHDLNmuKcM0WNX87AsR
afQEZP7YZTZanQBSPvoWsy7NLt8UBBw0dq2Q02Iqxdbp5+Eulvv4fe3MS96Ik8k6
luxS5KNvzpKeJFW8+86R/gVYFEcEjOlY4qfmQu9fwHGa+0FwYY4HamWCQKtNhQ0W
P37Wm8nktq0subrK2SvJ+gmkoiVhru3lNf1aWD5y6YFPUoWFaPQfyD6KoOTafp/+
oUin4fjyS+WnGjb0IdfFjxCc/35a1q3JeANMS4v6eqLy4pimQDIweEQ/YnpEyOW4
frBEq3rOVR8lNkqU0Lbf/tiplB+T3mspW94FFPufl03sUICm+IrmnzVBz709PVpT
eSeGQ6GY8Q4VLlaWn61kdqaGdgGFZLuH7BS/DtdXkDCXqn5A+zsxvOxaoFRmV57U
0uByu/fNojQllZRJ0/W/q0PfM/WOEL6jDFk3HsLp8BRZdAPUD0d9XNqp7Gy7V7+o
I8HSyicJtTdWsE4FGoCfzJbgXXM2dsg7jTXyAOpvbcCb0nflWtYbB18kW4xBZ2xr
bRGDhB9trLiou/q7tOPzAfzVEtpblYCcBODnhujasDtJHTji5I5yW+9qjscUCXOF
PfRU6dLlxxVUGgJtOd7FwbxY/b7yE0ZjH4itzGDJ4hmZ4HFEUfDZFAExdjqNbLPZ
I2Iq/fSEY4QQVKMt9TvPlscQ29alPOGP23Sqt4VMR+MvK90vxbjC48A7gaqu3uqK
Aak1/PQVXpElKGigoszMsvLdvPDgpocPXwLfxZCkx21x1AdLYWQshll0Nyonc7Sm
2Fsl5DYW7VQyDA9EnC7MVPTHAJIQLxMlwORVf8hCv+IbwqPDdzxaVDQAU5UPnx8M
C35AEk7SmZpYOuO4ABke6oJcOMnlwUZcoUh7NFb322vHRCoriQByepe7hgUfi+e8
9VJhijJCyDEc01b2ywG9ewFpTNx44HibxYFyJ7S7leU59NOWX/onmvFpgPqQUxPx
ZB7+/mpmzAppZ1uGdubdPS1fEiKQah4Q45aD+lgmODa3zQjGJqL+IHyCzT6BE+8y
+rspb1M3bni2FGOQf5cBP34e1iGpW9SVbXJq9TcunOiGwVLHOjCccCx1mYl2nMbP
ydSw1JE91Z18iQOkUAFDFf0Wy8mgrb6FSUuzGp+AItdsty4iYPhQaCD88O2xg+Tr
nBOAIPN+lAcinKVzqWpMdOvGesKtb4a6IO/6XBjuhyV0hJ4PmGdPt5o+HEUxo5E3
gSigZi9lQjtk96wmyuyA8b+1Op5Y7/3VhDNKoDCBdXilXeY5WDRuuFkFosGPIwcS
QJMtBpd1OFwGgrLZcwB0uEBaY+w/16qJctmZu+UXKlCXFXc4LvxLa/pKpEuVT7rC
MOngl5/+G0jb73pB1x/BY7OKQCysbEr7BzRz+I6M5uIZ0x4EO//8eiBWy66k5b32
qGeBcQD0ZjMS9amAEKdpMSk0yt5YmJp3Dd1vcrOjHkwavj0Ui/f+m7CGQBE7yF+1
nUJQtfWxM7CvloWvJce1c0uIFz6bL1a0G+5COewQom57foKmx8mImIKzfBHWMYQM
mAdKm509TDjUn6obOHz0H0OyJ/UuuvCv5P2MyL8U+UvjDOd9sX/GhyiVK4nVHQTI
WVJFCabVRf2iZpLZWRLiUn0P+s01zx2TUeYDH2oRWsPLubgxU8m7WQmowV2Q0jR9
9Oudbh9VCuWdnGhQG9uJvfLoGXphhBJP+dPwvgH70CeQ9DEM9NFFGEuqXtXfWE5X
RRbtsPfMVbS/Z/lG4tFUkEIClMGHumaqsy+V2l2wj4paAxEVa994PQsMrb+ARWcJ
VFO84dlrIFH93uvpvSNACRO72d/5vZzSejck1EBgMv25bWBBFXvcNwFVUzc21bKb
8G1wiiIrafzptbYi1jzRGeim3oP9obUF+gN1R/HE85lOLwkptWKaKy7D/9Sl4XFR
Xl7A/HqeHJn5z57Yew5AVRCkuxQ7m6Va9QJk/8pnHdqcmlr4yB/Mek8rg3MN0/g2
hcugTdNF27w0e8F0bm4ZzpYgFStkcBTXKNzFlsLYhrFF8KE50P3wZjtru9A2mzOm
d7ODTabiXZOgl4MwF4C6YBzmRfIWbn0LDFalvHk95+C9Rpx8kxOPBRFDlbnkDflc
SDJIJGoiRTr16EAk9QxyJ9+Q+kpclI/MXSUP4rAiYtpj3AZnc6nwP+xpXUrUmYLN
K9KbYx/NS40QZBCE7nTnD+s2V7mQaZp5Ksot+oW0Iz2jVxbTS5uoDjIelxPJEmcd
C32m5fmPpUdWuVRsfSFitF7iR5qkyK53yWZe79ySjFvxxz1NZEo2s7clOOD0bXgz
fcDH5ibtP+ARKAjZm+ygNss50cEFVrHIkC5/UuRng5rS+k52Ou/YJolQ+wQojmLE
BH2moxhOJVzzoXdNdd05w6CjlUNSRUWONfNBMl9ziQCvXtzJ0wdddmBzYFOFsszN
rUOUqDFJ8BeboON8mjDdQywncANigyboefcBQcFJNaKa0OCSgoOCUy787aukd2ri
tzsfCb3aupOUUzdTwdE22/6cj3S8fQUd0MUbqOD8niu2DuaKDwmsQ3DorPLlSn53
JmqZA/7s2a0YzS3gFVRd4xJs3RB6KYmZz5uAt/dfKtaAuUU2fDRwPFcwXALg5WrI
1e5BaIa5SnrU0+bbEMPc3U1oWImP78r2Xun4KtyPawRzMTbLmiMNnjU7lBRB76Mb
qMiECfdNG45XH/pc7oCca1z+P+XU4n4Bgu+QVfTexfS6VFUgxZIivaDJSyNt9DzF
SjMZ5BLJPirj3qPmxeQGnqE0hm8OlWtbKvHqnvxB57oHSrpA4eEphbfCpTGSz6hZ
kLeAxACd0TJAw4ClazGxpEgYWb0VIFpfngcxk+AcOQzj/rsSZTJLt2OoLTTjeAnf
iTjJJ3DoyknYAeccTuIiL2agfwSSZRHZKsbASmfmdIZZLmy0e4/6UbNuGjkqED8U
eMpqQLjyyPEkWsozExH1qyjnl9HSM8oMxXggMe5x220lFuS4Cg6wHBiCMWx8ciU4
zIXKqv2++YniV+j1+AXp/g59lCXE5sxBgQAxrIObbT3Pa3p42wl2QSykdJCfiR2F
bEeS3g3sPu9VE7cCJGzVr/glcnXfSDNIMWF+rq+XhsuV+dF0FtJNHZC6GKwbycQ5
FUhWQxxD5Ui63xMh6vr1WYtlxLXxT2iiUgdkkndQEHQ9nYsgyLZCpc1deZjymL6c
5jAFR58O7oKd78KDm8Nysn/LLhpx00aUL9RsRPvtxeziQnQNVgKaH9IQx3xhU3eO
WhOaU4IZqyogEMptEQuvcLjoJjLSsKsOmahxxYXVQxMYT7fmWYvnsDMjSDJthZ8y
qkviDHe3L7B5L2xyPsYAkHZEURY0qvFovyEFkHq2ijHkn0uy4L4WUgVShitviSEO
j2MIawkBh5aFVo7l/2yU4vR+9ufZjgoa4e9RJL320XxYjHJXCSL/wrUYAGXUyGPf
q9SslP8swyvLIpI1eHuHoXuMyAt7xHOYcxGUV/bPQ1o6ka+G5Df7/7uaj/yIQfaI
1jV6nPEUOx361X0PrNRbLnh8pn5Hu6MKRIyS5bpBdcrRQXMPGezqrSPW3qRoxztg
b/4gmgNm/wuG3EP2S+FRZF65KVaFathyEofPacMhLNF21OwHtUMa2lUEnb6Wvi95
xOa7JugkBizuUJ4UjF1Oow412rFRw/nRmlQLEjYQx5SZgYADOYerGMdGfbPMX48Z
zQY4gWhJaD0maOP8SCtNte6ue4Vn2hkODtdYM+XQ1EpMD8jKRDx8RGXEY0v1cBi8
4E/FIaHViGW5FftQFl2+WupBlebHTtyW+hg3YK9uwtlyr1nInyOMmwh1TwPi/Vc2
2Z5Ck/PCMmZcPV1Y863R4/G6rdnAh5fyBsbDD1yJz+O2hkNwl2GiJA0OOnkUjs4n
F2RugKR8gq0QJpo5btZT10g2n7uwHDFDQGoyLZSxnrlqo387nE3vyD+kVtMSkB3/
GDLicFG3PTw4wdJYYW4DM/7zkURlU2tA8gzkVXvZOcLFaEAH2j7+tBVxiRT/wxs8
JzPrsRmDea/92QTWeQkhLzI1+eN26zZf9mv1fUjySi3fGtVz1eAqsPDhgfyO7P9o
mz18kV3n+AcqVrwZ+c29p7k+F8GGnygvDa10LlcXytlpWQ+SlgVpe7E9Jf4wnGTA
I89VoRV/QMISjpFvTgi5CELxRWr8us9NHLOvzT2YQ2YrNDk0Ac3vyeTzYpEZnmmf
VQNOYe5NRnYRByYgx2vdLiYMc6n+gXJjlH/1Ps4OXd66dacKVQVKxIJM8Y5xjv6a
0ieqqxHoli8d4P01Niw1yEuKdtaaQn1XBJbl9408PFJQIMyzxyf7z5i6DIsbSx5f
KU3dZUiaN7RweeZpb5yYHQiBYrIsqqg64f7yRN/HZIydE/+p4A4y8MFFKUt7e2tx
hUsBFhK4l2JtulTg39Ey9KNB6WLFHVumKHlNqdVwRRpj29HD7uOgS73ChW0ptuUH
xWXvhhQ09kKIlLaULWAmXL7ZWta48qsUMQ7TxmTaBWQUljQos+i08m2EZM2Op8sI
gSY36E/TNHLhVUWTHoO8Xk8LRIaz5BvB3wnrlrntQsUsLuTgYjr9TRacmP43OWSa
8PwgHvNibnhSYrDhNCzaD4MQ+sr4ans8Nxoy0Yhje6CD8a+GyyajP2YnrSpkoQvt
SHmrhAgACG6PzCfxbDobZbSXPjWROAm+v9zh+V4xcmLQ1u1Q4FgVLGjrWAgd/TFf
BUx+s+FWitv6vUrSh+38o1ZfPVh5DqXrevf0/hRYicsdz0o6yLg8z1ObM1cRTxXb
PWfIYmYx5QhRO+kwCVGcLg16/lcLzgDOeZtGzUPZWhKrxZWw6W3PLRNJTdShte5d
q3UbqzuGJx+uy9qLS2L4yZDXjNlAK4Z+gCAwL8ANcCuQExZDjGx33HIl+NyjQHLz
bcbyJSIV2yBxiqVxJWJa4HgFMnQiv5p47mYhzvTS1+qigyRZkS7BQu16lfmfa0v2
kCPTUkP7rg9dTwKa9pjqj/ms5Ybl+wWXIK3jr1tSANavWfpfECVzXs/WSff9ig9a
znEWVGOguOgJpiqwTCIKz3MbgY90qSDx2vGBPsEFgr7H8VO9Sb2Cy+Cs5lb0XzqW
+sWmcyDzZjNNTyYxQd2cfGtU47U0ZuqslCHrDHCWOkP1AH882xkIefz2Ud7TsEXi
T/QHcMfVIuOPpdD9DDTh418OACa8yo7U02qYDL4EraZ3HNTzDqTIZ/TPDMxdL6fc
nbowuYRKyzZKauIJ4NJwLOXQeQp/3bcypEwl+wqizzZ8up33WXeTa7VITmRpVAyN
iGP/936JcMPD2aPd6ays+gdMBetnbtaNCAOVETo0He8ZwuTd2cvZDBEHSRduW1a2
6Cd4sKNzDmtOeAJ/EYbiTKc6bw+hGviWa7NWxzsPYH2M9fzE22mxM2JpFm/DR3zU
As62SLOHy8aq1/H3562q50yKNDhjpFqo32LfYFue7Pwyf0JRVHN2LNqafdEZGZxY
TOStmr6EY0+B7VO/JeWd0G0kyMwmOxeTsjosVXLs4ETso0SeWGJCOX0KChkqMAEd
SQjDeZQucUgrSa+9R3/siH7R6UE7ohRaikKX69+5f2ELAqPhuUKsLSi4HErcvI5D
rI+WtBImVXna1UyikyR9FtsEjhFyVPVy3aKP+MK5OeS6UBJ5NTRxCoCy6/eVqi4U
zvhey2dnzzAiG1V5NRbnYnvIYHDg2m4HOvBF0l5FdDEQQegMoUtJJcJZ+Djvk9Iw
CCwi9noVitIm83tWtGqijYl2Gh6cmjLa6RHL/EVe3ch1pruEEvYUYA3NhJmKWltH
RJMIyiwQdd2aKriPutPlBGdwJSAdw/Q32eLREMNMcgqy0FIe0CfHdIa3r6pQ8ijw
QkOQB8Khe0MV4a4kuU3M4D92l/Xw7cas+36nVHnH3vMVq2a9NHiCgIauymQXinnq
zmMi9noaKW8GlVg122R6Zm0nYsbnvjI1bTvj1Rw4TbtNvurISET6EfShfr2O3wf9
BF77Xy7U9apeTET4P6ubo0pohplkmaiZW893KSsY1Jq+yWqo6P0ILAbXh1rnIW2G
iXuvaMgdt8LLPauDVCMHvmf/6MOvWb2AFbxZ/bLY+XqILy7YvPK2XfSVA9IcExls
CkJpospVLbpkx8LskRkSy9OfaNZCutoaStfHEFzkxuIHDPzpQG7zfNLF98cYh2EI
2I6RtEIuhpXVq0Q0XQA/IWXfWlrIQBG+Xe8wMmZ+QnMnG1q+nY+NikOev49F9AH2
4yqOMFydAC4uvS2VF7UvH9VYWHaEgj4VU53WPcus6gPCOoXW4biDfW2jsBS+/i1k
WW08sOMIGnvQsZiwofyDUpD5lZgr4VX6eoxdJfuNEZM9c5LC7nZdsaKadGIXKj7P
5qrOrnFIQTka54yDIIHg0oZjXuHUl4Kd8zs8iMcCPuPmol9YmBJtd5MFAmFtU/uk
E2gMVIro6RJwEDteTUX5emi97g3DOnV/A8DFxIobLzUpnXiPQWofcl0GWdUSGW6w
TXZTddkib2A/adcMujakpmZbRmPGN+QZHaUDAPCMpXA93Rm5hdIhWOUti3HNg99b
9JI3hFri7sTGqHffg8KjRq1o9S2zjKoQvGN8lOuh3fUopNmB8bQUihZDiSXxHzBt
WZbpTZflV0jEtxkIzNoTFDJP+pPTCS3uCUOTSSG43z5zk9ip4AR7DjXOFhQLzKjg
Hb8vjaknpw/L/lkGfgdYnr1L3LG5BWCH4Y9y+EWrB55duYe+YGcD0Dj0Ks3jtvcm
Tit172/kApeZGlBA/3VMy+g18mGP1vjSsguZc00TTlM6boebRUkNuDRLxwc1V/gy
yUAjFYwelO4+trhsFAHWqksM2aICnfiFKFCTvfP0VepSPiyd6vjLM3v6lIlmsnOJ
0kEYlfxvEUBMoMHD0scpnbk0rgbdw9CAnc3yQ6jE9L7t4pYXF1kCZV6tVPapN539
dgUp4pP8eczOx2VOAdUBYqLXY3xDXZIen7+qM3hozkRipK/jUwEoCHTJ6Eh3AUWl
sVcidTr49oc6uW2kwMSnpmny/QD/V7RcI8kz4F3ZIRwa85gn6W5nwRh/SnO4G2ad
h5ew485ul/hFUhjCKsp9MoC1tYnmeyY/pVA5LbwY0eVv6akY9sEHCSiSRNnhyGn6
PrOLL2hSXg3rmo5hKK68Nio5+AqG6zsRW8JVnIhKgO4qL36xqySJx0oj6b5gfLVw
ECrHg9Jes9f43y0n2QKVTUOxySxms+JBURvR+wcEklzamTkysMxDlPUs29uzwcsl
yQ7ihWf0rZxyz1vikUo53cGQQ+fIOUKAQOyun6Jg7NfQZdoMYF+8fER9zH8EhNsK
KBXEblX8TmHACDUnqkerIIcZBSYNoKBBVGCqrVcDSM6aBPVmCK76AWDr1pxVi2yn
9pN76B2O80qg8KF5KkKeds6TnqoJLlVuldHsK5lw/zuM0+cN24D1J9dEhMIzGEHw
HNsh7VdPQ+rph+WDPR2ParEHqCHnkQx17GMR0xsA3cPyuKJgWlgoLYTiMX3/BmJT
2DD09di11TAncYComhhmwMIh1Eg4Q51Mh3TmyqBWiHrSsUkRqx1pQYgQ00U1YEtj
falCd501evEVZLJSQH8lqwfME0VbcLe+jsGEhDW24IO7kWQVbvqWnFV8Cn6HvweM
A9rfKu0s4lrYvEQfxrh8iyQ3/eJsNl5/Ue/v1blbjsm8YJ2OTUp4WOtqoQFvZw9P
o8RSUeMlp25Ws4QburfJIg2YIL8Zx/3Mf9Ux/sfcPLfxyG5gRt7X6F+lQI/DzLN9
fF/XIcJcBIz57yfa1W9YOLf0vlenLCtQJihead+zfeR4P7FCuomQ/CN0Ef9PmpxE
huMIOWBN4OYdjOIuDp6jye3TYHBAhccUG6vlOxXuNEzU6eFZ4YttSKWOJBS4rytn
Jh8FAfhkoA/9by/60nWM7yK8VAr6mG0Xdk2MpH0gfTe5igvmSlPm1NYVNEFWU+DI
Vfgud+iNhqzlh46Pv8HtAK9Jm+IaQW8v6GKu5rDtwAFEVHT8wwSbVHFZ1XGuTuzx
HccJSKWAKZot3lfBwjaU/8D0gBF/ERHBAQ37XQbGZZ/XSTFUEcC5UNeUboka4sJP
4ui//lXzbH1RI9A3AViD+HhZi/z5XzIbtB+XHs8qWJQ=
`protect END_PROTECTED
