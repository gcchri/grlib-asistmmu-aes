`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hF+FjmVsZ0R8qLRPx4K5AKJK1u26wXGhz78DHjWH1AXoh7XDRquy/1TfEmniItAE
dX293CFwbicvYX0RW3vYrTvbHQTLzloGQ1cFCvK/gqfZWkQdGDf6t29CKSa5JvRY
BQW3M06eL8M49Emr6kwhszKy+O0VXaYK7UboyD7ofPyBAOtpBAylS/UrDSlThMVZ
njw/VXFqlCzwX0xHKlZlQSUwp87S4bF/oWBsrkHUSdqwToYO8FYw4/wp6b6aLWQA
/7GdnmCKPXHrD4Nef5+2pAAKEsP4Z8bYeL+P+zonA0XBaMaaQI//2ucUmoI0KGyf
b/A3zGIzTPnDyWpfTLn7SS2B+rKMseLVHsHsrNBh4v5irngOOo8H+LFDcpsh7LzX
bN6C8aRtfP9KCondV/td0VPPnIC9zkY1tRxgvjah98T6hveIjClgxlaHG7hdPns/
`protect END_PROTECTED
