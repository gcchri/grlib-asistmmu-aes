`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SIEwL29TqA1FdLnE6kdGqfBImkghEZk4X9LuIxB8feTYlM0jDV0rY0g51LT/XVKe
hxFoWLR4FcB8UItEwl74MFvmap671SDsfCJyJ/Hns29ocOBEGqtLChe1Jbmp6wol
F7afxBdEpQqjhHU5owv5jHaPe8w8dUL+/2QGbcjxDrOtL6G3m3/S7wKE8C1Zjzux
3p3kLm6GGNRRk/J0At8ugvNB01t9GPQrJapfRA/eyKPFCDgnFz4+q7YSiCyc2V3r
uQPsJgPgLUXW0YAN8tIHhvv3DdxkgzuULe0wMDQSEKXRiMvlDkQc1EJrkLgWl2AY
0uRP38XHZZuOzjU2DOk3amhzZqbNx+7Eefm0Z8WO8OVVy7gxTDUnEjEh1kjjXWmu
VNaZTLkBUe119w2RnBNeEM4wB4zsjw+ahjhkR8r038Hgf9pWozwpGnlFhZHRGVgP
DwHlTGG8D7bOTsiOadSmlkse+LqFdAspPrnlWgMtLTA=
`protect END_PROTECTED
