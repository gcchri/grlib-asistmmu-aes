`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BmJfaxVDTkuB/VC00p6EYI8hB8V4iANcEso8XwIu20r01J2+Jy84g2yPRIczgyqv
WWdzLJ7AHdl4fwWbBFXGcGRLZR82qvfTPXLxSEXfI8yJlTAcsTNqPB/9ZPZv/KOX
s7H5xF7Ns+QJYnbJmUYn+WnTFtNoWlw7ttFBWDL9PsUKGBeoi/FOjPbZ1Tfww0SL
hg+ipRyBIRJVw1aGZYEyqHZH5K8n92CXk8tTVQAhmftoNXxlrpp4Oklqm5P/W0QH
Nj10RQ68B/zovx6+M3Us0OkfCHBMgs1C3fEqpN5fX8BWLWUhMefTbdFFdcfuOuXC
kam7WB4jJyK/xbBglSXG/avZX6wv5hiHUygp/Lpvn3lsCK22DB8509gxfEJow5rQ
su6UEZc5/YzPqqkCzA0cIpJMdoQdTSOCwt/+epDtZvt3sugVGa64rXVWb+yhnVb6
NIN9hd7xZrRa0h2/9Zv6pRg9Ww2nbCiA4bscJxDzoW5inVGJsA6glJl7dMwscSYx
T/ndqwxxRm83Rgm1jR1v0e9NO3mSdX7+/6YR9KbYmhXv6iCyHKkdJcIh4LuAfgD/
o2fXuA0zXoA1QIiQGuek2A==
`protect END_PROTECTED
