`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQCS7pZ42T9vkEFk2VApdgv7XnjubM1QVaMuzRmmfQmXOQLCweINHICexVgRMDdU
ipO7Lsvac277xAqTiDgpaVEyaHQW8zAcoES0YgcbXaLmV4dgxTKP+YQKEDEgdWfU
ELI9W9eAyRxQZ6LDfURqveXhy9gerxxcmmsWNvx3Hocr4fUlpvUHHchSXbNVIaFO
6zXJfY6JwI/XHkp2CcvZVgiLK7Lh0oPPNY5F1Z8BOuueLrBoPq+T2Jjw4ZNLtvCA
YBh8wIMcVfqme1JGesIqkHHSs9LU9xYfkUaZ6aSEel0X8Y4XSFYVarYzHtFbclLC
1VzOmIqGK+X8x0+kFR9It+yaiAFLlLD8TZxED6k+pZNZsNQYGf8Pmow17VryLLS9
wcLr52LA89HTy7YfQc95KDk3OTpH11LlSQPBcrKAaz9qybK3UCzzxMMVNtb+kHg/
h3CCgghxpP0WljcZvqqENA+b6E/qbCpfMYw64Dw5UzROvy4Nw5/rVWhHa0XAqS/z
YGuUvW5T9OeDz0EXh1NUHyIC7vBTfVRxhXBslfn7bHc=
`protect END_PROTECTED
