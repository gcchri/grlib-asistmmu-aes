`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+err24hcAtlqtSUZu5r/2RYr3ZRRb7K2a8gsZn6I/7pNrv8kc/Kr2kgEY5773AN8
sFmEaD/I44tT8rqdeRvfVwu1fXdoQNiLa/Q0lv7REkZ7Od8VMCY7mULS8zgaeHuX
KwwR4aQVBqELnNw5nhElfDO1VwAHLYDHbhj3F0eW/6M8b2pxRLOwDBtPH7Fk2lEA
dA9E5WgotpFTeIn9ZK6noeu5gi4HeEWUrbS9TcFKF8uXaq5Gfz+USz3gaw5nKIBZ
t/b04FBZSNGcGfBlEl1vqsD18+tVsd5K/k24zTVV7Fj+5xWT8YgsmNb1ESkem63M
E5phAUSlrnvd+FDI6c4L0nQsjh3H7KOnBc6/ZeEDJEN/EIqn4jsR1zQziCyNbeiE
665eqBNjSAo3PcUsjVbsDfm97IeVRBT8gZCTbt+y/Na63VNfXU9sYXFUVzm3DkU9
OnW/YZUhNxh4LrTH5bK63jslVvQbuhB2rPJh0rvDY++TDn14BcYL3fUjM1qWLfNf
7tflxOPGI2JebjKzN7ozbc1RnuAAtZkuyvdMPemF0P+FOQTLOENEgpCLrzMYMLhr
O47L1kgv6uOCkR1Y/kkmENVkgElF7rVEJ6u6fXT5VI2Oee5qZbyJ2lfwGmd0p6XO
8LpxXFsWV1fFVgiaHVc9Esx0cQFDPRffv+jeRtTwQr5AUJYsRFlQ3Gl2Izv6YsYX
bUrayvLzVMzxepkDBdxXjGJj4GdAygysy+B9RLyhh8O3Ed0/Q8jbNC3wF5viqfT8
XcEWbdmJUyXO4w2g3LZle1YAtlbQFs8NtXrZ275ofbM2ac4AzUfW6U2BmUGY9cZd
kwr5Kn41jCDrDoeax8Zs4IPCzlmf69/xFulPfaENNjLXcGiJ2aAXQD/x7wMi+PwQ
f3R4zIu5EqsOOK8rZrnNI4NkZ60d74RvWsEa7B16fmvGmdjtT2kPEwBvoHMK1gjC
pqqmd8XdkvBPv0eNRbZsD6OF71AWFt85I1tF5qYXjKrHWx/3mRmjjwSMV64JcUK0
FwuRv78kBS8z+s8rR+Yg93vBwN1yRR0LOsoO77dQIkmIodGLxCoiYyg0ZR/kN080
YTV4jRsd+RbvZR4jkWhuMZBrwmdw/PxdueAZvvUKeDWmvvo8LDBw09GOdLncoaqo
DA/cXOT4jXOfzJwtj1Jj99pOyM2csTI9oIgQbJR13IzcYqX9X6dfa0KIdDoqP6R5
DKe4z3+RD+CIxkyPsShjnnN5enGjKu3v5bFkHzl4ixWmrKNEfI/xv14tvzgBJ8Wg
k+f9WteYNKGj4THGEqqoNLUAaWIr3crW+eR1MOa/nzlYyv4UQA2MbK6Jt9cMfhe2
FjD5aRFs74G3dYV50xmb/foQo3KlNeX6ZZ5Ca/pH11mX4hGOgaDAMmpjybb8HaoF
+VpQc093na7DkYLhevJLlCk/AsvfZJXWjUA6ZCqJ4/kijirwYlTNl01dO/3INEzq
eQ3qSovmumqgihO36BZeVkwrCAJ7W4KXk0mm4Foo0YN6hhswirjc7VVWrAiDOC7J
XOei+vVVMpdGrpejk1WxJ/cJ1kUGsfDeMVCccTCr3lqq/PKekZ6MqaXD2tfRJaWv
ryzCee4coxRarWeiyE6EQFdjPXNPvxOT1Qf+oHwTeqdHisbqyKiUSEmR4+xxAYWO
NzczIU3rZ3A/svNCFCMXbeD6Egk1Mzk+tiLuozUXUxbkvrV6kAJ1sOZ83EuNBzwD
9gz6DFSk0TOha4GA2c8HJzlGXp8SoGfVeuu1e3iPq4bOqx6RysAKx6WiI4UHxs64
ROblbc9ojmgmozZn2IdUWABFaZQSIis6mnjK5rv9ZZsY5ELo8oAWN0N4fIpjIfxq
W65eEedgvwI8CKlMFMoQ+tkzTQvpGpOsr0J0A2KEyjBsuNFwDmosz+Sis7j9KNsk
70/DZb4k77S5wEJVUk7sI88ALfQ/+8WqFiuBvgc8Drgenb+D9NQ4WwpVLuafe6SK
hRsUBwO+py/6ogwIuCEzrvh3cHP6G8Y6nk51jtGUeyurnU/kVwDGy8acqMz4EKwd
fiCcgDAcsWA6zbwC7Liu5TBeGcHcx+taB+057L+pJnuh4ewsOM2iuBIwBXJIHM9B
p0cJNpBJswKpvnx6aPseu034R0BwOz13NsTs1onJ4SVhpN1ZKk70DXbXFX4Ruj38
hmV5brxLt8jSud9Jlms0aP3pdK9bVggUtFWsT145vDfKv3BGa3koWSHZbf9alyH6
YXEpa11MAOniDGfb9dGXxma8d815FQ+rfuLGTsAP3IXklim2DHtCtwifL5fu5BMj
DorFbbbfWPM4Tuj/CDXc+ZcjFAKfrDoQhq7fRMuAk1iezlACZTPBhk2RN4Cdwx7Q
7RXFtzmcsnpUVrX3d2QCAw8/n81Xz+DQf/hBk5SyLhLnpRAPnQaZcAkOagDuDmtp
c/RKKk2HUfmzcczj6vGo8omqDVW/nm9uZ4TAMiUIhGWY3NfmFIv3RlZhAV3YUXgh
5M7Srhwcuf+qA3RixCkjrboIAgXFlybWFz45Bas0WcATCGyZ1F/paGz+dPo7lVNn
LfFOhJ26HmMSsyvkANK5tz+Bc2ZPi0H7Vw5jf4xquWYnEaJt/xzLgMVdv2zLW5eT
a8ehf1D6bLIu+cTxUbTPg4kfHdHoxrYnOpahNoxn6Jwt5B4tfyAShaTeS+7k4ec4
HrYQkWq9WLxqdtoGotZFjnoaCdej9pszmrXiHUeD08YWeDTayGf++UiYCDJv7FxF
ETqcOM3vJjFbMqmRVeYsBgwuikGunKY5+3RkNVZ3LUi1L856yY/Yb1CKmibu2k9Z
a8sEpabaxoIPOJ+n3ApHtegTyZUpFan7XMANCcDLUIpcA2E+/SqSIu/kXsCwW95U
B6R+A3P7nklFLWlE3jQkiBmreSOx8DrJ+gAxaThWeXBC5HQOFAhOTPlZTfI/cc8v
yPvGT3MO74oMJqXtHHmGEWPpPHsH+lLssPaxiM15onCL2lItIb5iuzB4aYEaxOEu
pUYMLDxzq8Ie7t+eNFEqCcbnc+EbE4bI9meVT7Qx+zp795SvVtsI33PfOWYFKFel
GZs9R0tJh5FzI+UIwhMcTA+Z9SQnhwQkLDDZsmI3E/6cok2uqqJiGVtMO9uHESYY
daN6S2l2bQr+Y6NTUyP3XLJhkVIcHaxWK0dv5679dolqfmtsPjQTkR49ZGdSGgEJ
WT33knWl0t83aK8NrgdIPituTb/W8CbJT9gl8XWUDlchv4KbELFcZlq9qHg/kCy1
IiWE8xECaXtociKyQLsgLlf8NC3HG0WKwd80Qov6s+6Foj5mPWuXTXmBXOW4CguZ
lGoLNdMgqDSApxT3brlsIfuZIiG3h1eLN4UIXkmlMLfTYP0AItUDLnm6mjNA6tdh
FAt5KjD7192/VJ9c5bGhSjsEiJsb4A+N4J/P99NpHm/mR89B0NA2msg/5AyhBAfP
35hgwXPDYR5BEjM/Tn8UfDM1xmRiQQpSlCtbKnzv8hPGm/0x38U4sneVcRhWLSAk
mBSr0Lx1+Teyq84r2JUsNhLZA3yNZNEbDJDvq+sstFtdkkqSHstX9MKCOywMFFI6
7Wq/h3gXqLXRwzdNWknHDlF5tNvnwUBxYXil0p6jcpcDPdaj4t4SMeaOBuZlkSe5
dDtNSHEO1DNatkT9/r0MK3J12BhnYqQ065yb3T6q3R6DF9t1aZ0/SzX1pEJeutvU
qMgnh27qq6DUZ8njwIv7AAUOekN8FcpwOSjl5/9B5Sy0efWeHbqaQFPtOMoPY5x8
c6pwwIWc7NPIaLsNDqrIiOwJ0gGJVUVfCadVm/QPrWMXStU7IlWZHbG8rfOT3ApB
8+jZlBAYNMryypva1t9GUoNL3wTXm+dXNxN4ZVwq4kzVeEG3fdmxqKC2vKoxKxua
4uwm1SjgBS/lOnhdBDs4iMpXI20LqhNkN4wzBw+1ERJBzj5TVNXxVCzB1GtHK5Es
7gQ6UITfOFEUAZ9wqewqFKNkjm5I1YQzog6wDoWLrPfPGgBxOzpdYqKnjRor/mAz
Y/hoVHJgTNxJbQhAr8P1aHdINjWMI94bsnRGV0ckG2ONuFHvdzMn+Gc3SJ0VTdSx
+8MD0f44GRL6lJOANU1e1UKz6xBslafi+JKEAQpWrGFGgcEuzNM4hEhA1rsscFnx
ldCgmOShDanjD9F7BuXng4i5/3c8/Ml7Qkdx5zMPvFaiVwnNrzaRy0YyZsdOQSLe
WwYInwqZWRUJoGrUVaMNizsXdtyf5ytLNaZfe0t6M0OFfIy8tZZdIvH+z8ubvTlT
WfXNEr8k8CkCDBsJJN3mbLlNwbqzsMqnOxzPpw1iFeLs5dCJovmRr6/IC2TK79WJ
I8PYWaRsBTV8iyhy87Xse6HLJ77TS5q52Dfw8MG4MHEe/+AnR8ueRiunxLN4w6T/
OMckyLQzCoRBdeKqNhfMPHRjlpfMnbbZ7LhYR5Q7NtM9i+VZSQfvE5JXKA/9OtjY
otc87ewnSm04LoJioMPK7m3ROYOcpcHZj4UBf2udA27cAnW+Twc9DG2vrAEbPFmW
lj9CG/4KmkqTWf9+aHL3QPdXr7addqEFPqkoxi6qHIQQpg+OhvvOkjZP5ClE8KJh
c991sKjT1CC+PsrmEKQssZyECtjpSfOYT2veczW/u5Y6qLJh/KQWo6ODU2bgFEyx
puMo58upbYPn/2Sfn5FD5KXH9eXaDCPGxx4Zqkz7UOf67Bphgf3E1mxE7KbiNXU1
Yc/i1BPlb2bH7pz3Yr5/auF7/9uPV6gb4mHYUiVRz8XbGlECWAAgQLz3vJXKMfHn
BmiL3G89YG/G+mLYkQM1N2i0N84+kHi0t4IPT5G/XtD/vehPP3zV52ByEKTE9q2y
PksD4mGp9MP4vVsstSP0T3PVlzyWod6VIN1kPl4KdEbbB6NqN0bqZY2AfJdMFdLF
z+xIsU3MLxSMA9bT1Bto/HwO6TiGFl6fL50H4lvoCgHFGGcyJrvpib3RQeMUumSh
0MITAtBOwOI8Adk19LCYJjQCH0j9c9HwGVsS0sYXWxwXSF0R+4H4J+dRQ2Bjonvm
3rixCR4IZGUWW0xZgu4RhpEHZVXEf5TayFC4EFleK5O6U2ExKhucNby04jkA4b93
FqjpffetogzKm53u6hEYfKPhpOhyQdvfIcHtAgzfoXpra3KOBpaeNQDGpGj4+cTg
+Y+nndcbsGSZu6gG8XJINz0jictrhdKQK1UwMn9Cgzi/5JhZ7DlVyjsoc7T/n4qo
mF/ts/fNuixbBVGyxwDn7BSF7tf0v+eqNDJssD3lb/4RdUUjlox2FeU6yBFqzqGM
uDYYkDe50FkBAg/jSNNPXTqEkF+Uh1biLggrKf0fBZKbB8QBAq84yxoEmDKRgIzC
9nltz4GLx+NgwthYlAooVyD5MUAnV5bZzi76pbpQdOIa6yK8pWoNDxuvG81tFJps
lab6cG6E22RAOp4ocmHgfdbR/ArwAaSPuLgVE3zKYpT/8cnNJ+emSplHFLHHUHNz
OxT3/J8/YRrDWUQI2q0FAQjOj2kQ6NbZZEOKARZQ3zQ8JuZLy6PAtq/VD6FwPw4g
NJdI8JU5YQGmMgxvKVWGIXEWVUE8cxedfAbf8v63woni3znuZY6P2xDoe8a/q9w7
Dc7GELaYY+wvwnp7qUedfzcYDA/Eh4quxrIVsw/cuDI4HpVb1cRxnVKvCWKBO9Kv
XYMCjsAEo+SrdZ8dtAHT8/3tnShcktNx/ash/JEPF/mlU9YtkQkmWt+MDqMvlrWN
VzNRRO+ttXM4qs01bNpqQgXkABOql4+0RWYiFb6vTA0swF6EIcw/iJcqATYTyBok
ISpe0isY6Fj8UVLCDg8mZN1W1qM+LE0GdHwEH9nUAAfxyrrbn2vUS9gumq5F0wpb
9SHZeeCZ3Gmzgy+t76j7i/0RbwZtJgwONLrD22EQAfuy/ngWHyCyJ7zQHnuFNMD0
ArkucJ2gr/gQjoYmCuCoRSd4SUB8Kyk/EsnrcwNZVbfBssQYI/Clrcb04nZsiOBA
0S9nZ28HahkvIAk8SH/yvHk5fNeVvzwbtts3ZcL4GBdM381fqiI6YvgwE/m4z5NJ
iALmVPw7RWxs875lEXT02Od7Y+uMgTC1qP8zfRVoycOY+iHx6D3Zd9Wr3ZKC/DWZ
19yaafnZ2XlSqtZtxM7gHmZx45mCQxNZc7ELvd6Ad5+BZS/V9oa2zv5i7JAohhO3
ncxwtSZh+6ADGKaKxL7Qyq1qg/mzAQL6n2c0bQvDdkmjMXS/uqqujOsZ/OW9XaHW
bSPHfKH8Cgki48iUg9GjTQqsBYKjtcM/Ybq1eHIxlnxeq/96GFJn5z71oj4Yh/GE
/r3RtEScJHXnapCcAHbzUiQZTOncAChilJ+ysnrY5Kh0k83uH63mqp/bxitRdtpQ
OPAHP9oqdy2dfkkIAWZivnTUz+RmZz2p1+VGsd381Pp5/wlJnHDshQ9owM8oXZ96
BO3ZmnElfRx5C9x9mI53MlHWhY8op1dhaY4aG9X0j71buLrqAB2/ld86NlHNdgLI
DuS0OQTGw0G6KKRwPglya6pJH7BrHJBmXGc68N8Ft1hEvKrKa1wsBaUs2LFcl1sY
M2HCARMApuJIhILdJerR8tBq9NGVYPP3LDtRPR4qlJFiDCE3dp0wbctAQqtFNsP6
Grg50MU/zkFgj53TkzXgJ6WofdRjBT186fvrBQMe1gojna6yob+cBa7o9b5FnEhG
XVeabQWH+Pc78mEYbla/ONbF43/bD+PrgbsWvv6jNN4MrAHFyw6e+Eir8F2ZaJbL
waUoHNV+QdHSgOsHSGdF3EDYIXvteikrs7+nVwD+j5N71xuvSjpLRA//A8Vnmu3H
8bFpjFq/Yf49q/uWCkDsayz3+XcCj2WrMwxRmmNn3s/yN5+yl5tiwAac9pjfqMat
ubHQvsSflZwZbAI1h+gnHH04nCp6IbGQW63hQhxifl/W9v9XfZIVvlTGJQ/GAkHl
jdRkajyyhNzQsQHqv/m0hWQosbgAZTLONHkI6O1OKFl9TSeEN/QZNwOIuE+gNZFk
9wuHJKY4swA6GTaD8T8ME6iLirmN2Sw9GlExgYGE1FRZR80P0eDrX5eav+JoTqSE
JB1sLKvNchpcqKKbI05zltNLki6VB3MMfuZpmJba76vdaxg/5FBA4SJLkoRxysRE
gmltHVbeUaMFotwcEbw2+hO6OaImN3x6j186/sVIS0ZimvazyRss3TRwZ+uMVw1S
JqgISNionUXaM3CGRc04moFHxlwfvWBNVQ81gHoE2Uclw/rFjSsz0OIMd+rhZ1su
jR0Of7fBGzearaiOLvLIQmz69bkiso0FoxS5y7Ui0EfxLzf/Bsv6T6j/6RF6qwY2
6JDFJwSlIK8noBt/bdOsTUie6FL0grKA2v7VWTZt+oqPGJxR77vxyRQMuXa+UrV5
xKZYy2ExjNnql/9eZqr4+gXZlebCFpZv5oZ28xl4FKQm9H+1PLknvW1uzpZ+uRhn
7TAsOMDeJ1aBG7+T2FK+mPmlWn+hQhxTvyjU/Zp6WgmdYsScjtYtcNGGUmvLATAk
Z/lfYuqiNUPFUx2pFEfrTPXrjzFWOjWonL0xubjq01YxHkR66apX+8GN3Wv2nrJT
jY4fm/dD8CaCWSZeC5oA31htGHHhauAgZugvkPj3mBluYaRkgvCwKTyuihSaOh8+
e6jdKEnwpaYeNkHO1+BgP4NHVlveD0hQOewFWK4hAY1DmEj7biFhGmySnAJpkrYV
EYv+KJ01i1j2vqwJAUcOthLHfv11BSRBd0K6jKswDMHeV7B6sNAqzRVrQirW/0xT
7NE6trpKGjgxLXbH5jKpzdzDodg0qdO2iPDXRHuR8soUxO3w/IFUtXpPg9IC/F+G
Ap2o2BWilOsYxfWdk9FJc/NoSQdFu6V34qHWmkWyK2WyRjhIgqViOuIsKoM4RSAC
cmsgmS1A4v7FivVANr1+1a1ozi4WG82TvwEGnFiae5pGU5iXiCERsrEYpR53JxYP
krJymofJK65sQgBYT4u0ue7P8YZ+VynlAcJua260jTVGa6UGqBkIJjTpY/csNkAy
FoRKYTNKe8uz40E06VAYxZ98D4jG1NhyP27yQnkFkJR5WfAM5A2nV1kaJ4u4ntHp
EZCQhlbGzoW6ZRsgsbvI64heEnLpPNA425zZ6ca174e2ihdGco7ZTzgFWk89s86q
e4AA7v+6KvcXelofpH3ZOikipDObztwmQ88U5UaDeBCm8rmYcqeBVwuRYW5Yzsbs
BrfLmxpN1sU6zwUdZb56W3A7uUoICRMSW2eoTSX4CcSEYeEwOdeACS5NV29I9q2x
6qbwKy+nFaQsQWb6bdO0Xe42HAxxV1MvcgyPuU1TE+MYadIrcMvviCC2N4DNH8zV
JXmKp5z+ZmVg2ipOgJZKV9OFKRTb+wtBNRfwDk5kvDeCf4RHp5mJkPf+Fn9G3XtB
DWHeBEJeU3ucGDbL2LHjVOfVXt9Ic45Lu7Hn13z6i/7r3vnCvZFI+HUpabco0Zyk
PnX5sXCoVuozpcpqBPfU5TEChwSrWtAgfC+leavbRiLbWS/V2X5gUTtt/EvzdFwT
x2j7O/0lM82j8RdSXvRJAlngOS/eN22NCSXK7zGMGvOAs7TurBcUOS3Yqzqvx0k+
4YH9brDxHVZ35gQc63y6nVuGTaCnicQaSf/IBSuRW+F3VHM5voFczNiFkVq1tefV
Oy1XqwcuBtusKH6OjuCHNrH3nuuVF0sdT2kJx4wPSRP6J2hFIocF/rVga48R2QKj
2Mwh4kZ+pJRARkjOovERRVfj+qGJzNZas2Ug1GGzzN0Y/Pqb3GhKX7S7GxzYFsx3
p0tj/s8Oj2c1lgVV+xPWwEn+Vplz+u81YAthBQvQyXiwT7Um6qwh0A5Z8k6svwt8
Zu+5WNez+7EgK6i88VrJwDWngDBYtft34w6kRXBZF8dFKy9ywHGmN8MRaiMIZumV
rEt7Lo1jiP/nElZUopYzSF5N4fq2FrziuaPFs9+f6X6i3GUhBlrKJNgMC24zoMrI
EnY5ALQzJRo5djSzZzA6viAqj9E3htyJronOfqPzPO41/J+zKDG/p5Np5GUz8B7+
140uyDULrgiTFEXL2t1knYLsZ8fbWvn15sqeXN5NNo9sNyLAlZ4GZmSodE8nxM+i
/iBB//tRUuwN4K5MsUsaZBpAo2WKNqot2I+zU7+iRAqmUdLqfuOQ6lt24/bxoZS7
ji4WiMblZMXx3ttC/Myo7L5eNATCvZ+/4IuGW37U+xr8mj1r1ISBPxlhoIVCQTjQ
uBPRxDWZA2cYlJeYlDrP0lClZ5h3O95R7oI6KvIbEfR749CBEBG2Lh6K9CfEiJtE
ZpXsisl8gcoSUjhkJDhKdb6KGDnFjvOziMX5vWTsZxMAANJH6KpOm50IaSbMZmjO
pncmWP362rbRZ+Rp43veGYpnGPWs1VM58TSB0rqnGb3La1ex/mm+Fw5ThHnK5ZVL
t7DjHE1SHVKwoIP7lVJRMr/R8Nrk379rU0PZivV+yzjt+KRE9EJStVAwO+uxDNZU
3eSPS1UQd0fUxVU0L1sdvlUq3kLzf3tWz+hVbp4DOPs8jh4nNDrwdqBSTVx77CRy
bjTYr6eVVfg0vYNMjLi5+58Mxdl6TXe9w+wr5OWkrf0FwICkS/fGWF+z0SpzW3x2
++8dQyX5JEtXOtYF6N4nutZ9guCUfGpjY0IEUdZS/qaloWvycaRzGqokIQyIIkdY
79yC4ECjO5GH9KAcnArsOu61lPoR4BRWmo4xVuqb+9ehoYL8pRB1w4b9Pgfq5w4v
khToM8HB7EEMngjYQnHBjuOEawb4SBBfYhgjoGMZM2QlImir56nKqFbgvVtwKsv1
GfqJfaIeNxbR612bJb4/wMwRCYH1NSuIDvWBfKLdb/13PM+20AYUyUiyIB5AM8mD
7q/1EofN3yO8U5eWgeFxZUcrnOR7eKqEaBm0bRmn4j/YvRfcdDTeVkUQaypqmEEm
bgaKVk1tCuVCrmV2nYII8YINiiqkyuTh7AU8AOCG7P8Og1X68+d/21pIsjTvozn2
DQ7qJXnA1JK0fuRlnkjjusJ9G+C5hCOgv9XGLbUzIr8p8anSuNGribxbasHgnvVZ
ZZfw8s0qY6+/EeiV3H2MVPfAOvNGqJvsOoP6oO5XqrRXW4PiedkatuWLjiiQTfx0
cubq4407RmfXAxbyfUjfNXoTjN9ci0MdC+sSPW/YLYrzMCqtdKsC5Ll0fXdLD5Lb
ZvW+nJ71ZBNTuDaqZat/uRCwcfU71RwFoFz6YvetoitcC7TwO8jPGmWddfh/EKWn
wANWxyfuILDt/qird1NE8mGfE4DC3JxIF+CIS2d9IbrqCGfNf1XljnRB77LulpyJ
pR4QNJhkb8EXuawIVNhxQzYcW0HM30SJ9ART5w5JH53X5n0gMy1RLa9PMwSFDDbn
ftKtlGiIY4rnBNOi8u+TtkqITNhf6lIvjVVAMrfPksMB5vcTfmcT24+K7P3W6q7D
hba9FXPAli1rH62Cn60X3XUNe9E3Z2xZTjXk/Cxi4B6tJEeQDRqsfDCpdLVJJ1SJ
B9n3WyOyma7xhGRf2j8mxxE86AIWX9k9oyvt/tAu8h5glQfDBekcJ1/MruMfIRvU
7U5LmJi8ZmwIHlOC0snzrPZlmr694E566rBhoPXIxF3hZEOnG0L41UhiTvAmWJYu
t6pn+P/Br0kJXZbcXS2U8Y86BmbVtKCqI8Kvljna2/hLTxZE3EPnaPhzwTicnJR9
lLHs/VGLXLYuSBPyQAlL2eMzcIlGwfwGBZA6n65TMhsrjJm6uXxCDdv1ZvkygpRl
IJHq5qdJfq9uUVyYp9T7ioVk3O/QCABVlpXLURVcxCelHXP82xSNa068R5veMwUU
q/BbGYSUE9gd9GIYaoDDOfNZGkP60RyfSs4c+PnbEZ7QLyhtXiZ3x9/fr7maS++g
R2W90MRaXYUjX+X8Je7eHxGZyDLMk+stcm6Jb6vYCWT3t/uEzmqJyeHwC0VxN+WQ
a2CRAMilUWEM90HsyuKrK6JQYga0wBkW5Dv1Kr5RQ+K0ncPC1AZoVZVb6JudTdYy
cuLZhCDehr7LWZ0Op2weg0Khi4dq4Ab/fDTskYcHKevcdg1bWA2QTmorFykBzOYq
mVaqQco22K8ugLSwsbAO+3hkog8y3IgqWsEIZm0YskGq7CJLNobKAZIbo+VpE25s
FziWPb19MzRrp5RdGxSD3QAFTZOe+EA7k9kHE9RE4aD0gimdPTgo6JS6UrHWPinY
N14jm+1nvemb7oCXuLPPq0ofPPsUIU4N5XjQUjhoWie29y7nevZqlWcghOygyAGt
u3UNz36Ksa8NjgFH0A2k2/Z8sWT4G56TW9Fz6RrBl87yMQlxzsJi/qJuGVIaDyCa
dCuojUz3cEOi8V44lQSkUk/7/7aAtvZPVDZZgeFFLuVwGVtbN7yLOo3mTcgSZ83r
47ItbrJji1qSM2jP4x36PsbM+D/AjoqsZIcfHXw0uBdjAVXdjLpxmdk2CfoT3gMG
oAnFxY2EfLLjXRy6lBrmprk/5mmUSn09rIpVD8boxHvw/gmdJ23rhgc53Y/swnc/
MkzoJVtMgYL+hGfbgQFBRh1Wc1w2u0e+2fi8tklqW8RIvx7Felmbzo3ag+yXxKia
4Vg0Qjxd/q1I3LVOMdUgSRhgWS2rXnE4jtFCw5I6tvcQoW+ArYDuhxI7e/gLcm5g
X2F2ep/RGchER/z5Ivhncu/DsVqiYTByS3XYejyu/tCEQ/TRbppMSgf4WLw5N0rO
wsVbDnCc+pTM0aMSyUzxmFMb+4gxzTXBGi3JOEGnW1qTVFyf3V+dtLDifYafymlL
K8gdZbYGvk+KZSpxTAXa247J0rNKyjdZy7urAhD3b4s0d+/q+qTB3VIL2v2iHkPJ
f9WdtP8y5u55IppmpZUhxpaLbXZZtdbXClHddjrdeE9RGMill556HAsWt+pBZb2M
nKjt1i4cO03/bc+Haf6M/f7d9hwC4fuCKTEwsIvQlEAQBBUDTlZpPzMusdKFhrDI
tSVTKPz0OwFXbfYHYUxQ9EHyydJomFvqz/u7QM5/IWurh5UjSD2E8e/AnFxNZBt3
LYqjB28ARRfQFIBJ6w7XQX+TxqrK+pAeriKWKk0EL9SCS1jSj8hpYjy/2hbtt0vY
oDVVFk+Sm/7GNUH1vFLtdcw64b6XkbrO7S7kkx9H0sokI9QUnCJN7b++HSUQk+9R
nvp8QjHOkrXBxIzt/Rf1F1sXvBwCGos7fhV8qoCsKwLUhqfdBcyqyWEkzebAcN15
graAJ18MX4AGF+VK7vjvOa6z9QfzA4R+Tvp3BRnXVTXp0waYyW3ar5Q7ek/CilA3
lDzawSMCre+ywEx2NiwDqjTWGtQSdkeYEwPi5GD8or0PSCJmjFBKoN6WdBctMgi+
Bzn6ZJ9nMDW3sWQNwcMVjXtwghEV80btjFrwNj4A1oHppgSOGm/Bj8Z/26A8wuP/
Ubz5PladeL59VnqCiH5H+CGkTClzWUqkqQkDWdhVyE3bOdXSt3az+gmSztgSGwHq
wcFyLG4UBkYEVYj5WgdqVL2QiaVTkvu6tp6C7BZ+abPDvyl0QT2UC/QUwh/bpRjX
gxjd5TCB8hPfpD1TbF3yIbzU5aHZ6yjzEk9nl/h5BB4OR1PZy4YZeuznxNMNjPw0
zjPgzuQRQin3YdsArvGXra4cXvb1PHnRyzCSsKCwO6wlDUsKPvutNBgB7il8tPqp
YfOTNAH19EqLmze6LlF9qC+J5CJNJwckiUOioPLed+Y9JYJj0g0kLnvYnYBXwKfb
zV5rnB2XCMnIqC40MgNufka1vOa3tbZ9VwxPWM+PX+W5o+2RQwgdN0Fy+wIbiITx
5nTkQtkJixJgKz4seVbW1NjjMmxwhi5YLZsHnX+rf/bDXOL+nEilj9DjpsFyj7ZT
yIxp/D5Dx6tfr1MU3qW49Rtt9w5SkUpGD8znkwxeAuJ7O/ouHRG/Q7O09fv14E7/
yjxE8AWQHmEGRrDRBnb5cN5Q7cg1wU1iQ8n8uNuk25id25jQCYM9xRyaPyzi5CAH
BTOa9LDdM65uRANVnPaC7PqAqKZEmB2GV+p0JjOlBYovH9sfWiMZoMJGEz2JsuDK
bzr0xsBs1e3fDepyf8nJBmuM/m+nUoTAL5dY7kddyoxoCwtH5hcuzj3d+hACny3I
`protect END_PROTECTED
