`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j1EWp4GOapVAEIkF1gGUzkZJg0H7FELEAMUdhShC45udu1nBbtTpJsNRFfIpwkyd
H0toGSGI392f3DLcU3TfvU8mq/mAuXmPyrz6vticuCdQYhtpGVTTu0JRKkYUioQ+
hgLXD49bsTYEpDtJR3RctuGrpJbxugDW6CCIeyWGa+uvZBByxSbnz4gZSgnUrnJD
3J39lNjNzpup+aC0yD5zlpXAJ16nizrvnKyqRgl0KLh7pEy3bnDOKbq8wmqaCkuv
le0QeqjeJHW37M2j8kSxcNh/0lQ6gXXgnnPRlRM0Xy1PuSeORtLMcBqRX3S/fdxa
xmVYHQe5VVZp+UibOLmZWfM2G3hd8bJJoH9kTG89ddlEjIEA3tJbQ94YJH82AjaT
31uWs6dSgTIYA/1HJJWtu6Kyrl5PRe1QCPRjZIhKaPxo4+zts3fLWQVQSGutZprM
DCq9dltqp181t9y7H1aQQP4453Xm2UKRPWCiG/WpnkC10ryj+Pk+lcSOMkm1v2JD
jPTEpiU6BBGbWNSk/Vuh6mfLtmagsqDJKtkfO6mjmyP+VZmH9PtyIaUgZ4JknIeo
`protect END_PROTECTED
