`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rs1emQ+m/MPukfb60IH/8Fp0HeH5YMP2vTNwpiJrvjvvfVSOLnsxB8W6ts7vWHZR
VT6pKwuP1R6f/fmjsmXeSyDLH3HuImYsAXlBhNFLyk6nHpOf7KNRFVJ0hhwfczkE
CLWmcdES4+d8F9pZ7D52w3b3FQ/Kr/LU9Z/aQLQO1e8KHw84PuPmImJWbsmUHyOA
47/zsAH5hOZyS0iweQ/du5g9LvTfUVT14tUdtIGsI6Kb9lCq4UtD9vk+kTvRyBpd
wKB6Nc8gRodMTWlLk52+daiQR6pQf8gWu/rQaE1G4RNT6s43E6de+PTS6r6go+hB
vC52H4UBLn1x52Q1ZyGFH9StE4cJbyBcFyInJpT6eATqpz30UWw6dDCm3/B3zf4m
`protect END_PROTECTED
