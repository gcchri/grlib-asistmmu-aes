`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DS6eHhuesa3R7t6k37XmzMfm4VvpWxjII1qaoBaXQrOotcgQW+ZnYdw8Zkjc4XwM
kDmny0PAhfepyjD0K/NGOiyI4yJkhNjgQ3TgnYDXtSOvFKIsRpID/62GdryzyBO/
UORZWOSozZtuxxNPavqFogNuEiqci46eR5rt5a23XHRNDIBCGEN/gBMyeKdMlwrv
4Rjmlbo/4f+hPfV1fsx+G7FCgO/T8BHS7kvgDtkaT25VhaPRjDpyuyi12QH5RUNZ
oHKpSM2o86wyWaVty9rePEtyr/byVn/AjoG272fWjvXzaesTAy1oANjLmrD4+yVj
DBcJVYy2BdQ2xdmybR+UBxkBPjarTeCSiqwpuYbGtn0l+7JfBuSlbsRrebQouHCy
fJQB0n9pvahrYkC3rWqekzOGXwLNIpcTra5YQgOyfocXM5MTZSvLjkjJGyp/bMaP
X76pUgN3qnwSFLF+xUTYiey5aY10yUaZHRSy0LFdbi11dJobvIjlTCv/R8khRqrE
`protect END_PROTECTED
