`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YutZln37RAmo89JHCw1iVRB70Y7I8UM32pwXFUV1QgJUMHYeBjEB/f/gCUvpefNr
HZbpP1krXuqRvRIgRSONUD06tocx5rsVHnilX8EB285sK9YrixgSWg9TisVodvH8
35BgwroFiTca+3u27Wk5JkNFJg5G351hxzQ5RoC3ENF1+5ef0MlEsfg3/EHyGJNz
bxi9jptw5wdQTEp4Ff6f7oJX+XTQRLstoH/JENWCyIEnzvCJuY38FRUFKLKmTbvg
e9dmKTflNykIchIXsOImG9m6jnUHplICRCbDktmSd3ESmj9X/uAZTH8dI1wHsTLm
62lXfb7RALDXAn9aftG/8VHfkIaiAYM1UPVHcVtHM3OKeicLOHlUi/ZnGNRrfvD6
2isxxxWlEZddYAvdtfunKQmWX5Z1hFii8SHkurq50hYvqD+Y7nhBDHLbBPbZ8IEn
ufL5Zk6CFs9fkKkdhTUeX/lUSx9v1GQyrytpTp+DtYwCO6gcUhBA3c7FQCT+GPBh
`protect END_PROTECTED
