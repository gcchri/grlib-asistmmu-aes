`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfMNL8Yc9l7glEI8XOymLRtoBCtQYFHHbabTlIrh93iY1Gz40lZo+YJtPfjxQLIw
FJEBJ2vFDAMxcbJqwZiMpDcTUrwN8YBFY0BMseLWkZfhGjn0FNd9T/VMZgo6uKzT
S5xvx8+jRyoOTolqESG3L3Dh3ZDwf9+o3EHTbKGTVTOrmA/EofSc6xF7Qkp93cNZ
9LjsZ0Q3W/SksK1fVNmcHT91ku78HpJjp6EGF7ttkee/rwAEwsoM0KADD9WZPpCS
tFi9KJtJP4APbViCv068P7+hU27YoFzzpHqdLmQage+ztZ6G/zNdGVtHB9cORI0a
AMej50QgyPIfNAOleT2AdCGxfslxeX7a09Nqate2rPrvPzEGdoqy2Bgdo3BG507h
z/Oav8gMIF6/ipvX5LSnSA==
`protect END_PROTECTED
