`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ge8mSBFZbgriaTvC6W+n2QfYX5BQWhzTCruDAFgREvogD3iQCOvz21t2yLrcbcEK
NoY5RQdrPZLuarOl/uMp20/CMLTotwV40PMZGB4Ed4TP6QtUI8LaqAcoTL575rkY
Nn7FPqKz7BBFhRfdGRgps8xBxks9fv566EuMXeQHCn/DsWj8zadw8v4hOqF/0yzz
/hHA3rgAz172hSODBWsfKwBFWRQ6j5WgUceBtrSZCt5+ptBAw5KUJmWeqUvGoNHd
ZUI7rOKDNBN8kt5YqrfhH12K5SdP3zGyU+vTgF950oa/VbS8W+nwR5M3sU3CF9tI
IRfNbubX42Pn5gdMI9zS+8bN3lY5uj/TnJXhf8Zcv47Sqbw7AeEsw3lrDaNCxeaS
g2ECQFS+VSbk8BwA69kDYqIz8fUH523A9P1ipJyhy40gQoOGPBiW6cbCBoaZmrH2
mevr7tLwc4hj/BYgzLkqDI26OS5tUp/Pmp0aPQGLMvyDFLjUiq5VaFve2cfa8jAP
FPF5cUM3NylsemiiD1ITeEybLWR5k2k5HaCUb3tH03gqD/J/Cx5atPmjF9RQuJhK
azpRpUZFzu7NUOOWnFchdBGsDu1vJtNJIl8qUJVhlArObKhILtetDDdmsbRteBRc
uT/rNeB5RAiNKQlHnrxDWy5/XNPyFpjBJXlyFIHm+nW+1HoQHjwg20mzQo3/3uDG
HDsMp8EqQ5RjVmTHrNGfHpZZ6MmtWmbmQQjBSo+RD9j1k+YiKLHBjv0afC6GIFIi
21+OgPrUD1rhNcTf3f2B369IrZhe+2sYs3KODIG3QawAs65+leQWfNnT3PaZ7dLn
pwIgZVerG8Ckk0bG05CnkdlkN2yVjiYb+MsmuxtF5pvvOCvETXr8tL1vNfU0J8kJ
9LQih1FGODatCnmoiX2cQSSHVTndyytnidpQxqZMDFpQxrud1BZ63u7e2AsjueRj
rRqG7/aVtZYNTCviEdKok1/sV4ojiRDm8vA0P7o4zUQjins29y8ar3yo6+owSuIh
wfDSkzZ06A4aSYpD416ifSkVq6Ih3gdP8HlXW7RV1EqxyjsS5omXEc8K2CNPRr+m
0N5grat2FkmPGhppE1f9fMjkmZxfRGXYfTo3oeHodab8FDOXLLST9ocFHF997WFh
8Z0anMgnWr4nMTClIOkB3Y/0Iw+dcYNKy+xVr0PYWW2WNr/YRZFXxdtL0Vm1ENSq
vk+lJaQL+DK84qbbPopyqsL1NPNq+w/zk/cJQAy1Nt8s/50kOwViYQwXqVJF+o6q
Zsj9jeHhIAMnuGjh7fE4YHV5gXPM9C638gnWZvDHkYRQ+no9/LPU+jYvT3nyRqFf
BQgCqJwzIWdCUxXULGyo4I3mqLuyL1zHbSThe1xDMIluH64fMwUbsaBOpvaC8KS5
e0DzVLUAcV4uiQIcOXzk4O75HgHl4qjccoEfUgQ8nA9ycItYVv0FDS7py4BbZyeI
3RFnQTHm07Np+MnyFIG2bpHC/jz944DKKAABm8pgncJUK8mmZ6JkTjcs1t/eoytg
RkGKQ1IGWBDs9FbF4Ctcwe/Crn/CyW3P4skLCfAHC4fkHZ65gk+repxNLW932eXo
vvoCWJ3HARdA2hjv24+0R1h+M8iLfn/ohBnlBA2HFo/GuubiAgEu3V2dP8m0B6/q
IEkbr2ejOMQWGfD8IKoX7A9wUWJTHpHSFWD2p+ji8SkjzQIeW3gKoS01/XFYkYeG
K7dkSdi2taNyPXuhdtsHe41W9hMeth3Q/9y59/vnV24aTMCVHFxW8Od8HuZhozn0
jSCnrztS2QGtJg9rjeuoQ4CP04A/2zL24qucPXZGPH+Vn/V9B4DQU8nwZ/jpem+z
pG4ttwctTzJsWkIDznhX8JycjStB0N6ixxk1O5Sx/WTGyo506hg/myB596q7j6p7
IXr/IgSs5kYr3gYN42j+2DobCkrBhn21V/aNT1gL5OPr9U+zcxmfwaHuWQCQP242
l3EIRybYNVDaavj3R0uEOCgAEQF5OqbryHFt7bVy/+7jre7F0w8AO2KQNJhhycKN
REaFu1cxvgwRDBWvKIwM+KbxiJf6M+oj6/V/k/frQGv1owCVxzOP6K+VyhJgSEUr
ETXc28BpwIkk1cRuW8VEnz2Pb7kgmJZPG2CRL3kVelNbv/p8VxA6R6T5lr1nEa+2
E2b8vtPCS+HxRJZEUAFmUWWlx6n5S9neWymyiG2+T1V1MB4LXI+yFX7MkicboKMR
I1verklBtXywWPv1DlHJEk/XQkuyMgaGSTlopLOHho3fF63yKmHO+1eI1YMM0vCE
fPVb9+ZPUUFnomb08e2cAeK0G8INeEG+Dz/Mn9yaYHq6oMyfTtp8p6xTUpzNpWGK
jhZg8sqxhDbfFkpP6Feb10R8L8LNyx1ylSAR5r1eopze4j3261joopEk66lRdxLY
3XfzjBWeFfkCPuH3cbYMLPYjN+gxvHhZ07MR8ZkghFsNht9YW/Kj4DKHfqsJsXuA
`protect END_PROTECTED
