`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k/zKdw8LlaxukuBEY+JWuO4ZUZc890+oEG8OB5CUY9A2QCFCzz8jVl/6WE/f7n9C
DDL1FKSfLXujRCUpcDNNRjVvphR9Z3N4XQygXTZsOYx4HQ5gn6El93ATT3dorn4j
a6srgTmlIszevRP0P3kJBudHkWKnfcZHzlDWFHOsLx69ucNhfu75sebKRRWRnhRd
CxPtVD0GJlCToAxvF7KaiWGp477Zuy2g9/KyK+Q8PuD1XKbvT2Bjha7sVeBRR3eL
F1a0GO9+EnlY36V0R7NtmForvfQXqLCDCCd8AZmoHErFbdV4u3AA5WGSKoR2KV43
hJZCoWtsnmS6jwg9mcrd93FqY2dqE8bSMtqdCTgR3BtX8CcWhVw74rU7lnCwxQXD
`protect END_PROTECTED
