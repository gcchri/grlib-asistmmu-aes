`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QqTxAuGuP80YOnfVhEV8lxmDvF4uY/eU/0qeJW68maD2Oa0uRva8HjxPhEmssSku
uvEmvcP2qDxVjG2bAKsUKcxVnukl/Veh7PiKGVXSbkYh40yupx0nUgekPoZFqrX5
La21Hmo4NMwzKDeE8zaYXmUklgY3Th0qUIal48K5v0UC3fvSD3fk8LexmBEnM8Pu
Jp9UzXQOusmsuFExG4gAYIFnlYxUX4Bzsicxq6jhpW1dLVwwlH32VDgrO26OabXv
Xot3bWdlBPtN9X78BytR9uLWhDofpMdDQRE9BfWmnNXlEFxLHp8MnIxXvqRmIgFM
xIKiDTYZFxc8I5FseQ4mUCABJXWg5Dt3wRjDSoDWfgnhZ3DGZVJmYZDKhRRTFxsS
aTzlcf7jvUxKH1ysKcBH6tDCV4uMpJunb7qy+GUdQoyxItHYE2CzwQmL+OI8TuTw
p5uvC7BRtIOvU/i6gmcfr+d6znb/e1MC6mo8DHTRKYtsUvP+okTXsWpKpS00VqKo
55W6wHj6oIl0ydHureIQMd/ElFeJBPnUxkphhFnKd7OjR4GixJda3RJn1cXTQZ9g
bssvr8g63bR8ycmpvXhANlGCZBc7ZIUT05uLiNnmH1/B7AGEtkYub/XeveH4jTQL
k9v89kC5ug7Ovi5YAcGCz9VhX9g63BT7JvsIz9zFCwJzXrDy557/2PRs4GqRgCUc
6bgkldQrak6+iZ7kaAqqZpgS0DawEFVwVO0B+KMgwE1IL7F3Smz5azhqXHKqbIaS
Elc/3QpLXaJ15kyL8K9N89IyrQ/nJOHpK+mSKEz7Ch/af0EMgIWX8mnesRfQnBQa
N3SWZAwNxfS7qS3yUh3xB77+zcuIpV6dPg3dRTws8/RBln0jDZyBZa36+RYu2fNW
lZSXTE+0id5766D3e9Q/0CNH9kIWa+I/XYcChPLWerDxWngHZ2EBYb6SfjNJQNaW
aPD7JH8OSvX1ts6MbeF5OECWWAExRNlXMsQY/WtR2ncBXJC/s4lkq3kD/VdpccJv
nXo1tRMLjmMxRVoRliUbiw==
`protect END_PROTECTED
