`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgelN7FS29tZ6+lhcc2w6T81RqlKo5j5JlgdI1JlfUcThI5iySMU3mVpXJvv2+dF
om9T4ifxZW+W0mse0UfHVsa6ZPVsxGeDEqNlzjR3TZdAdmZfSN4JdkDaZE16ynKF
ZVbYSK3Q5/8K1zfDL1JbS5U01o1vNIQ44qqVGji/ZIIyO6/N5i5m/XOMI6JpdF5i
DEUX4GoFUwjqvbYfk8QCvK4Kox00UgJDRvH7ka7DWsR6YqdOBvTpH8v7gNmY98s+
dK0khquVC/rkbDJpufxCjO4hnrQmZkeaI+DmFHjs9Kz8+MJeajqDmRYqkay949Wi
NJW6RbhivLQI3pDgdOoWe5erJJaeYdD7sWMSi15z0m50GlbnHnbKgco4+1vlUfIW
QNpqnxXvfxHKSlB1NaxpnjkwOxarTzPbD8hJijp1EhcXFGXbBCADNs3tOLRKMj+x
I03pwW6n7nU7ZNonTupp4ZYj1Y/477wFrOp/1Zqj1L6cqsmsNYfnUIVbFG6gdJH/
LBnn4TpqcLNDgaz+TAOixmxLLHxc4C0hqJ0bOTWfJUV1cEW6VfA8M01Vo0R9p7sX
9XAB8AOCrgTTL7xMborzENC7EQk1Y4T0NrUyEZG/9HSny7GA1We4I+z0FPBmiCyx
ythmsOucdAtS/TMWT3ThirJKkozgH7JP6UUqqqKhtxlB/d6E3gdg2u5XRmZ2WiG4
K4N5HO4mCZQJ7vV7kDTXFgRpmOn32gwJK05DH2/vNA1Expci2gtS0vSbctUonv/7
xhOn6bH23e2Frzcklsa9uMDGIzUKEE5FYeRY2iUyH94bkbPP8CxCfp+dE2YSJgYh
FBXpuw8IoFBdNMpq+7svSw9DvGO6cInfhgC+PL1+evuZXHj76Xxd/lMK4cFpSeOX
HauFkn+JcRSaQSi7SLb94F69OngvRlPnxHUE1/vQeHEsajSaxiv+xdFWghD1HFLH
Z+biZy33Jt4FtcbFthYBKCTme/dW1P2z9RHve76vtBJgHkaFnJegpq4QdnO/b9ly
jA4nKoDCbqK2r1lfdlQkkx22bRbBVSsJfwSpKRONb+RVD0JLhIosei93tLigHDuT
+i2s24CK0h05UJuV/ZDDVfkv2/6ERt6wHC2hQcwvoQ8ep3wKyqyk/RVXMLskaTZ7
CcY34+1gMusdV3yyX5sH73yCM1jCwi1fPLgNgTwVHqpJUMN6s02Vfloopvyl8I6q
nJ6OgS9OC6QzWQE+UkAT4k9nE2NacREsr4Es6sMkEG1V8XuwFNMCt4TVFBhEn+i+
nCtNP6YQqW0u4gpudyaPkZKWx4pqHm1gVMw4Uwx4l/6doIruP/nhLXBADTiiU7h5
3HICDfbakWm32iKFFj+HisetQD9uBtfs4QF2Ym5O/tE2CWhV0jpyiztn0V4tCWfA
kneqlIwWF0Z4PU0Zf1vLS0tyt6duSkrmy27wr6Dca9bqh3WCos+vTnjgcsNtqUNe
PCG3pWtJyUWQSMhj8zXJP2oZnV2Y1JbiDdOx6nEwF77yh4Hfs4ekjqrl//uH+uBy
O1d/HAYFlWEB2OKpQ/HGSTJJewa4FeuLbEmL1tCSpwScVP2xd4FqlyWgcjaeIMsX
LgA53nFLRqBaO9TzrdFRglLC+u/m8bonGRyTC39B9mWdBMf9QqBQ0djn+KA76Z9v
eTku+7gPBc4XQZioEIa10lQ0zzFKQe7UTlXLRYuVgEWBRU4P2SqOT8RT2TQyQ/sB
ndcVnMV2ZObLol1ZJhbtDXHL3tPr4xpwmJjaDDqQZc+BoojGyDH3DY71+i/CqrZB
6rEiihZhfhkEobe3WsuI3ZlDiDk7KsspeELwwwRc+GPxtbsmP8jNQ4wT04HORR5K
j6Mat0rTvulWlOejbzTEAiTqGDOQ89KB1WNKyB+0aJLaxGlV2h4JaqL03xG6mpms
SQ0g6p4rrf5agrguxlajUafuTEJCjgBW0uHVuboMTW23BcpUqxtmhghbnCusb4oN
oobsrxw4meZp6bfwe6Nkc0uUGredVeqdhD7Snv4Eht3/Z7wRQdrd9dbi94QdJgKW
OxXOWXlS9kaUsNPXyY+E1N5EO0rw3aIL7Q8yodB8bJu+55RvChxjLxyJh23eo1L5
wv+zaSAO0tfXDNtKMEQwFCB9TSox7hRpJmrBMrnNZLbI8R4aQeswG73klUPLJ+Kr
VJmxc6iSdNtnR0JNUJ2XDHEpebdbxey0QVWzje6H7foKDeu+eMXGLfZ/JKsSLLr9
dJbMZBMcy3PILMTdUsM936Ff0BKBitFgHbhGOVLulprMSCx3kpbuDrmGCR7sX4BD
xftf8dIwoJJF9kSaTcoDW+253jZ2mIpZIsGt3dYoh3M3MP8agBm6Ltdp+o9crSBL
hED2dbFwMvxoFqxwgjAYtWtsh/mmxdYj4ADtksagjiz0+SbZZ859c2NV1BbPJO9B
9bAvfvfD6/dWC2V/KhbAtJmaKwrbeaQfVq2aJxW6oKKF4G+5tfHtKkBCueMLXHdM
WmzzJRZTo5rxf3+kxPv3V5WgNLGpMV74mSwXkDy0Mo51OWY3htsyCmbX7BeACq1F
sKbH98mMXCtaxuSpGC7fNFGFALVQvg2t+9wvbRxmVJ+RDk3TF2PME1R4gIv0vfWL
b7W8aWRQdW00fqula+FZcYHTcT8omYL6BpOm/oknTUaBsVBj2WjlUhapdlxiiY2/
K28aT1Zgeco2X7ISeg+u8TM2V+eXSAOU5Dwy5+95bAdbmTSF43OzM1+AXkSfsCoZ
/T/yI+fDBN9ICsNcxk2K1d6WcYuRqsOx/VoDz+qFtJbFAxwOEXdx8A2NKOKq7xRH
FDNFyAinxuaAtnronn1IXO8DeO1w+SVP0uCMxmfQ8wSzHs8er5Yl73f2XldR3ITz
rSAPlLx+aj1unxNgpm86a2mvnHhK011NwBWfYzjO/cbq9RN+lDYYJ/Ysz+17s5iA
tTNadoDo/t7xWTttHh+ZikwBSJ5RTtFKBfMWIDGBXzVR7US5yt7f8QL9XvnSc15o
LldkoSvwsXpTgPsHISzocXTMJlbPS9nDNofmO/t9r6/ttllMePirpILmGuhSebQw
Xo82nlnxpqWcqF2/5R2J73AslRCbkH0yQJYNQZtqt/JIxHKqlpPYRM/R23LI82oG
3u7c0nImq3o9xIV8QQlv7Gw46tv9ydRNvRr4ZTHgrPy02DBLtARel7Han/Wr9tYz
tZZHIlmBroevPUqq9hEYCQ==
`protect END_PROTECTED
