`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a5gLBuZQbFJtfJDXgzwm1BEhvUIDQ17Yb8JqHU/19ZBWMQvfu3BOwRRgaiHqqqZd
JtjWFe2UkzAGO6WrXJfHYr995PsKy5uBeZ4vJHVOHXYyDHTg866OJWXZ30yIcScU
7DXNKxdwRhparzOR1sJz6yQHonxr5VVtU0D4gipqti4PnKbVP0SzcJfuz8UObHR5
9d8Fz7CGIJxaHMBe5HQ6wf+ZWacWLcrtcAgXc5JJR/wJKIB/uzJQVHXhMy7WLfch
P25dL20sOnwut+EBlZA7aDgsDjhrS24sx/MuUW7fpnKMojMQCCawRly9JrDByp/N
Nacl7a2aSMXaXrIkh/ZHrVtVOZ/Y+iph/5Ozy9POks657ar9rB7Ns7UuC6sPtZDA
F3iIp9CdLfBCIBnRFzeQgAkXq4/XwGmkVyAC/k0XDLGB1rKlCirSJmHaim6GVn8T
+xdCXZgFJB4rh5myQR2HrfMvpDt/K3PwVJEJbohU1vqIGuTocLJuooNLZnekltnU
dQev+xIrpuR7LAuR1h2J+UL7DHx8BnUGBYXYKvh/6uo3RgJETCUIZGL1BcBXblF9
JIONNQ3CD8vLSPGs/7zULk9ylDJMDoV66+fd87DDUF+jIPeMQZR+Xte3PQNkBtvE
i+gplQstzqEuJQJamyHH+kVgfkFCEuxxFKOJLdfC+ulV3Ycv8s9gileSrbLR8SYA
FVTGsvZXAgq+H8CqUZ21z1WNoMnMkRUNZ+5RiDZNQITn1ajlYu9Z0QSzUnwoBslY
6liHP27T+NE/BHWrvdyh1YOdoBAD+hye/2ierKCYNeotx/V6IETi7fmM2+9j5JaD
Da3nr8ToRs/ssGngYCkZF7M4BqoRDF5oRw4ST7/SwJ8=
`protect END_PROTECTED
