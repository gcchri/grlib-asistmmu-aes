`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNxFeMRhrHojuI/JASDYrPs4aGQ0WN93lVfcDdfh3c+dY00oZqwU2YioAoIVOeNT
1sgCkSa1+pxtTPi0uS+5NF9s7HoXcuzswMjwvT/EhSq+9T5jc+YkzUYh4RpN07Qp
D/+po+EOWyt65oGNQ9cKtSb60fOm5L3quJB9M9JE8+um8OitT7RpflvDkoDaKpDI
Ie6x8fuKNyD4X5yy/l6medrDTa36+k42uho1U0yIwr6/J/bszkVA5XDNvDfbSxcr
pG4eOBl2uIdVML18Zn5rhS3NeISmwXgC0tU97ChvHKxaRpD6cIU+yB8vu93FfqZs
bS/dUyPlWxJf4qQzeXymgd0yimyKIDV6JWZQkt+td6/iaIpkzSPe4uzybZ3gNcU2
oRhj13mlKrVnlgR1b32SZBev5908RfFZBl+CEZCTKc1McswDTF7MotPAnfCEKZrK
m3QREhMah40x9iPBbA8Vb6cm44eJCXr7KL5lktzX4vUMmC+wx6JgiwpfgnNDqOih
qI8gH274EHK5ISyz0KanBU+XAOpSm95h4D3G9GqyoAAAVOoc7HSxPUL5YiYfWHPR
TOQ1RTKEogHtjZkU5YWHwZjwNWqy9ByZejm7vgk4NSIcyuZyvNpXvPvjYI7e3npi
C+2MP7V79lOKCNletxkXAKuYlRvJ+xnvW7QrQrtu6CeHqlK0KhQdMTxLEyS+5VrP
lVTMs/lxqzEliv3suIFEV//9dW8O2j6mLG2JZqY0H+b0qG8M7XPU4qYqI10k8ftQ
ryH0xjxsCUS+yuJuUUxDjyARiyKa1Sxad9617mIxGDIAy1rVJMjnilH+akL/ZkBd
6tCexNas6NXRWaQlJpL8FKLxYosuh0drJQhET7//tEutpfgZGBPWB56dYf+Do20P
p7UOKYMviD+tvl3JsoWpxaNth0hbzYtKJvAuF/Hh4EmRrYlNWijredPHV9lI8hho
IZMt9w6lxudjPvsWKHzU292aB9IY5jlKdhUBM5XPw03vjnIpVujpr3k/xEgGqw2S
`protect END_PROTECTED
