`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8VjT3PWsv0DgIKiwmSHEy712cWd6s1Rr06RhesJWd0zrrSA0Z/+RuR4FnJd8XZJ
F46+GVBWyeZK7w6CYevOuiymXsUi75SRcS3W5lPdeoscYoPv7flC2XqE+frK446Z
+e4DUDLAK7IwVx8HtkLpYoabyvDjS2CQQZK2FKHboRvRSubbBzyez3gk6e9Rtn3T
2E//VJlkTVWjuDyOh1KEXN36VLYyLYPYoOaIKE5UzC1vrJovKMFIOJtv9WZsi6ab
vYecDtiXESlZnJi9eVg/xw==
`protect END_PROTECTED
