`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVd/xs4wxrVnnb/2uWMTetN6vnNGgyx8KRsMdLgNJV6q4VAIpfWm4tqMshb3aPvW
1HrLV5JChAe2QoHyUY1w+6oqiFUtAw3+e+mjiXD7Ho0HdFvYcQuZbiRWf0FTt3kb
tNXf8KCMVGJhssu1KmWj1Dv0dN8INZ6HVgfvQByDe/vT+9wMMd3CtLE6p3Pw365R
K7g5/siUGXIu8xQZ9/F6BunTRtlIhJog9ZFasICqFFA03gHAkSvp0xpBkidz/0pq
ZgW993tNlgxyQZzgc0ieD/GdHh00p1SomTJ9niKNSlV+gdGMOJtFmVM3nhtCnvCF
BevFGoj5S6nOkmUgvpQbABRXZmQ0Ez4HAWsQXefRQMEQNboCyBrTuZzLGtDsWOdB
oA/fSt2xGmq8rbDaUvymWKKDAd51fq+nZGjHBdRhgbpvHsE3TXUhii1zEBlZ99te
63lOZJ9iGNSpMnEfFHJG33NuBgYNezpJ2oPT1wAsHgaJwwOd9F1gaDwusGzM6SzW
BbNX/zbrcEu4A/AUvo9vFg==
`protect END_PROTECTED
