`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vja0WsAVXTRfPK3GxX7BOqHHoXx3g01qied+F6nM5DqiRISJiNVU+jTCQCydQ5l9
YY8Z2fp4rq6Dk+QmjHLMwSJsz+TfK48rbJzWhFPXnS7f6IOUQFdTlcxcW6v39Jou
G0H58mAkEHpNh3WcaBu6+/IM/jUR0xkHSPhkUQPV0C/kat2W0c/x1wTC0pa/tUWz
ybaSQOjpeVP/o9t+zNKyE/Y1kqSXpRlTvfuwZD/gRr3QRZR4DieHSBsfRZ2qdpQs
WDHZCwPyuU4/sC7hde0Z4raGNd9cmWZq4/DLcaUggXdlGUVe23r/8jCuAXPvP4/Z
iVIY7dtLQ1F6WC2FEZay9R1v5f0eDJPS/NNlliANxOAHPGxnfKsiQFC8OdYOhbiU
0P6BpQs2ToxsR7GdY7dQwShoTTMJROA+w2G+2lAn3B8jOyczMWRCTy6hsbTJjA+A
duVa346B6EyLUwHniQRsjRtfq0B73aHAZaXw527zsIpFMGyfXcrAERKFxlTK5rRv
CRMqwWGk5/yKBcfqkHH45VOzOj89Q+QzRihBdfKFOlwUeul9boLtOcLAoJFmP9jo
TI1Bcd1VFrTzVtPtunnqLMkYRRy0gGWEJPu2ek49VvpsGzvuWBNmbcYDvw718PRe
fGP2fZvXSkPIfuR8OCGrg5x7ltlX5oth+rsKdRGFMZezAGFYOnnYRvNprCGzumAR
TuEM5N5/m1fp5wa6SJPRjio8Lb7gwYn7OweKP/XaXaPPY/rIpdzPxyI1Dkqs5I+Z
GVV4EXWManw7kzCkCRRUFv8E7negUzLUx4Bp8fk+6Lq1ZhWBjz5aQAi8Ds8aYgaL
S/vHwP0EJCKu8j7/W3wfjuj2+EaOeXlw25clbjl6e158OhSDuGZ0Q0LWfx3GoNEi
Nkr27gdojwk5iYGJ1+N+xKREStbcXRiVBCI50cueivfZFJTKXHWX5w4Pz4C2mgdb
DoSZGiy3A8OfCDdcwOM1L9bKqgzXyGMp+9qx99DSH0BivZ0mbJ+O1gHWD6krzUf5
EC8hPkWvvET5YBP/NH2Irayf1QaTPz0Pp+BHr1vnnJhm3AHtfXZqievCCQl3M8rL
/SKnULTdGhL2BxgJEhpkDw==
`protect END_PROTECTED
