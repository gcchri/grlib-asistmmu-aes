`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sj7IxtAyqg/srbeRZ6mmWSTGOjm/7hnHF+EVQ/Vw8kXFYUD3oRti1b9IHjh6Meh1
xIBUEkDwq14B4whX3ul71eT1srQ9JEbz7OtAwliRrwkWfrxGEfjxc4tBsyLPawEa
ok2mVe541CZ4cMHtM+93pyl7Cv2mel9XbB3IOAcP4iVLD9/0oShaMOaJt9nY787F
2SDGi6vAJi4ttOYAH5E6JeaU9tXzIPXCGLwQ19oznX7jA8pgqnaTcPN+fl8PxUKh
MqtvSN/czf5rLGJdcRv3P75mfXCZ6FAN2yW5QnTmo0c+fCpFB0h2isZZ8c2tS2hv
KbzMZ8nciCQinrWhdtjv6LTwIOX1zcFK/4yCARQ4+zqcqFmhg5R4t9oZSazWtE9s
fnUmVnZsd2EMplnFgmU1GIuW2C/efogAJsK50wG2iU+0ZRbaWayLi1Y472/QeE57
k4Yk04F2kRNEY+tpu26rKoSPX90BSXSUJOU4qY90QwNkJ25Akwje6ef5qlLFo5a3
YEaStI8TSUu7wmUrfnueebG6yr+BU69KcE3t3MxEsxgcSV0guSvlzXbSRROQqROd
pNVLtDjynd6raKYfVkN5Zp1VOi4sO8SWth8y8lAcNef3BDcJyFwnOB/AikrLjSf/
NX85V4dT9Gpv715UpTlz5BT5Fv9a6pgP9lgcSIDWeQY=
`protect END_PROTECTED
