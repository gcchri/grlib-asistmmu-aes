`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrsU0bhlUO9Fx4d/IOzhgGgKGUoJ2iXThinRTCg0sKFq88/LTuztGVtv2JrNi2TA
dsV+gxcZEYuqDUFgffZhkENj+4gKmi4aGRuWl8mkIuMTmigjhaqHcJpOnAc/eBzf
Nbx2oU3t1cpwlsbvNVEw5BKdDGm5rLDPSoBdNt79xaIaxsNC4HjTNI4T9oJuj2TS
QN0+M8IMSvTLQCVT/raa6z68srkSfT7N84YBxquUE3JoEi9JLkLd8pWvRgga6eeC
zt6eT35TufQg+oclwYiezSt54m2SYhnfGAlYClK5760CBvgE5cyGo9a1SGc1MQnb
ROUqNFyY3ge+hkBiLp3LvBvOJljNajDNyW3w84OLzrFvelMc8GmQKXKgezKyAsh6
wUYbJWKiTNSdhGOhoQzNDaM0vDw+XssPhfP248N7eUg=
`protect END_PROTECTED
