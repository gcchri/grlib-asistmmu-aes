`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjzvTNaRPd6C7BOshVEnhd01EVlajQPjwtIh0PCm4F00/dRhbh0Fz20TanFrCS7D
kiGCn80lrjyK1Dz/TqlJ0uZdpHQ20oOuuL2Zh1V5QLGB9TvGodJ/sy+b+oQGCNp8
F8KkF0aUusjexd1QGKmE5xm4RTFZ96hiWEsffRCPe43z2ERFDvHeeu/G9U3RXf7w
QxVKetbeXgTLIUrW2XUuWu/4OK0wQGSd8kWctnnK0YNsyC/nf1orX8eagnKTpLVU
kk4L63Xnpj6Ct7UlHGh5iS5teA0bkotvniYB3ZkvqFzNb63XYDt/Bg/1U4W1jOPc
pJV5yCFlA3kTCX9dnFh8mN1nLYixP0qGJt0CSYFD7NsS7fsZzTqtnO3eqmQ3YV1B
E2VJMHhZXfZj77guW3q0rKA8RVfXc22qMBKKML8nPZ//KAftezh5itQcmR1MTAgZ
`protect END_PROTECTED
