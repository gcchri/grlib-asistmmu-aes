`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Led4tFgT0At1EMDhA217uJEjr5kjmDr6fofiAUzdMi/XJYRYScBdyEB9KByeS8Z3
S9/a1RODDgXnSQm7Qh/vvuIu9uQsR3PbEo4ubPxNzI0wzNh6RgMugvQhF1h2/jLf
ox7EWuOE7hMGq7aHVQJg/DvZdQoByYs27d6eEbLjwnwsSXdc/099kdYhJF2VWnDK
0wc+QDSLtV/nj+V0u7fS/TxEzIJeRC0DMqBO9U0lmBALL8RpNKoacygKp+WaRq7U
l5VLrIvaULwHADwEpVcA6Q56J91GE251sE8FSkxWU59R2lG2FTDMIEq/8IYy8nnF
kQIbCNZp6X4rjF67WWJ5q4url5wlpk+0x+LBgo574qhylQI4lXtH7UtTOa81PG20
9vtaSaGcLwPAx2e4GHWXKdTlTOKfMfMOHFVhtzRxVzk=
`protect END_PROTECTED
