`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VS3Nw3zww7SQ+0n6ReQZGbg0+nDOa76At5bJG4QLKNY703R4uGmR55HiiO/WYB/q
yNKN4naJQ7+oATULYagcjoFzL4hh4HKDwMP5QLryAvV7mKOwSb7ZrRRu6Pj461Yk
XJa+zmrz5LYJ4bMjfQHDY1KhYJsRAc0h/wtdHy4hX6zwaFA9fYmpmFvLCQTjTduB
h2o154oAsew4UmVNKKOgaaCb1XEyaNrdo2eAK1/egoBdsVeaDb3BzPfMn94OMkO9
xYQNqxQIJBdCGiOZFfx0JOtFbQRXFsk/9gdOldnkHdfyt+lye9iRCf87cSvVN0y8
neUPe/bZavF0CPCeka1PVMM0x8Wwyv6pxxaC/jcHuVFnhSY7Ur9hxK+xxLUvX431
yb/J/fr2G7U/P8P6sGNoiVIhTF0U4bhHEYOijipnNKZ53uSXtWgwxVCKoD95Gq7U
PbUiJZp4G99D5fPQDAo4inMuy525JwAOxQz5/BOsv9dGsansZVGReJyMXAaUARSy
cVV6SULUUbcgHkShJ5AiGHNyGKE8t6rzmkfEMo29RFooAExVhwkHnjBq14xPKUM0
nQ+h3f8Q7TYFgDrR5fvJkZqp/wwFlUsnGCGe1gkps70hdtwrwWClQNUu8WfB5fez
cJcFaOPq18f2Zyvc9TUD3hI/4hfpYZp+n1g57CfA6MM=
`protect END_PROTECTED
