`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iVsi7ZUu7EWDfnDjCLzyiR+y9I4kBBRPIG79+BnaV9nBqbEfrUNpqxM2howGdwoP
WVs1rjkFzxSMS6tw86L7CDOouvAeBDeqpxJje7B2CPAlm08w8jpzxNs9HYIixH7g
EKpPbLVivp+MiU0f+dJgVgxKOIaBx11aMhgfU7xH7UO2+bybb5IkdjMwEL0qaJp4
JyZm8edGppZq5VxyJlo8NlajKjurlb708DW9N9gFGg0epsXc/5qoiOtvc7kwU8w2
kUED2aPbwArsBqQ9WRyjw8g/icyCai2vI6SkUMVMSFfFgkNf695hMVOfrYJV0z8O
CNKkJr8dTV1769B/IRILelBish0obQbkGkWoJAdTqzU8ltXdrfqfacpQIDIskMfb
krnHpF5XuBwIgUhSYPK9jDUFwJuRvDwjUt8ZO5QGddod6+l8UxZLXKWnMTQA4Oye
oye6cwJAA2UmsQWqWFgl2RGGTJhcNKbZiWXV2dtXILEbcFa2CjA3DNVVPXQ2RyO/
o3KuFFx1PDSZBR15LBceOCfNlPY+XMd3Ry2wnp703K1xd4e851nKtji6bHAF2HOQ
oTEIVHk0H7gjSdGhuxkfMcjiHLAeSxfejlEeJOi82Udl7OxSBrKGJJGbnB+L3yKf
T/heJVK2wPugnLW0Ckgj7uQVT72IyW21KDYMUKQ1SY01lPWWxPcoNU2f2kLsEvQQ
/vsWlehnTwoFWuIcn9Vfn5EDDbQRcOcvIpYX2+ZNygYqeluyb8w+XvOrz28z5p85
w/im4bm1NBf+/Jq/Ct9pP5rVm81vipo8jV2vHRsftPY9JW6bqEJLh6zpZccjAH4Y
lpzOT8k8fQnBNrvyQ3+4C/6jSESoXEZ966G9EodCbSuI3C9NyWDMloYPMfLlaauL
U6NFb8+VOco5WUJ77ju+aDr/QkacZyk05vp/HgMz3YOlmTBr8eoe1+dsW3J/gJDo
N10bTZNRBv4PxB3XogKMKBnHAs/gqLXkiMzPGrIpq4ah121nxb3bFT0m5/3hAf7p
FXkDkp5Xh7Pjt9dqd6X8BUxrYiMefh731JxgjmOStHy/1VAaDPXTFLzKoL/615OC
Rh5WPWC3UNV2GBcZYl055q6T0MkEs4bJtpUA6SUbyayW3LN1Vcf7PNtAYaMGOTyB
AO1+w5i3/NJuLQ6g7jBJ69B+ftreOuVb6KS41sW/otwAMsmuOpAlLLNZ7LQmV4J8
PqYQWvYaFgV4lMrSlQvUQBTQzfSIVfD2wfuF7X/qC+1ILyykQMATKVuRRaoG65Sa
Exc+33QZ6wyQAbotkmwQSOWg9x41x58of51mqnK3/0D0Wq91Y9xj3ugKnjJ01W9X
toZf1qjC5nJGRmMqvPAw4WMi0nburSQqvl7KQU92w5lxhl63WHVmP9MlvRdzyO7Z
4ulJxW8OrSiqE+edz0DdA39GUXhTfIW8w7Vh+uDg/4Cbki1lvweN2RIahhiUQEjK
pY9N9vtnn+/jJY/g+TuoWwqwyNRJqndAHWQkPtXldmxOqHv/WYEL5nqHYLjUisK0
5SCAdI1V/TCj+4iUvocSDEMwui/rKU49E84Xd/2un9wyK6sfIUGZ7nE1yykHiYuw
4Qg8EtoW9FmOSesOQOH95c9RFZTGpSEk/H9cUo/S9NZRl2IQxhbuAIk6EX8iA3Pm
lpPzo21v+SIgoEeQdPxyJThUIfPx+k4qLC0JGW/UbsfX5m67A/digHGNCMCIbEoA
GW/TsyBeE8oY3FtPiSrFLEpoNAq0oWvUPC9MTn2CcYdQZ7q1l8kDQ0YnCHfjeXZ+
aaz6aICwoLQOaZ0TAnzEHkxZd1wh79ROBqqzp0kxV94EpgVx5QYkHdOfJJNEGKDc
GtTAArwo+YISV4LJbP8VJejMuEBMd/ehIU/dFP+lQ1JjwYUDgTvdxzukomn+Teio
+3Y+Gd85wEDzORr0wP43g/c2aZvwqJ0dNd4bLZpyreGYynC+CbgkjuuUpfwu09fL
WRQQ5D+Z4Lj3Kt+XzyjtGA78wRsDw7xXxBKxTm/30PZjzCjMCwoB4LD3cpOfWdw3
a8qFgYEMDAYWh8Sxn6k8BPC3ZeBfQWQaCaLLfErUZnxYQp/EKwcOlUjb0HNy+y+x
L9kPhtJs95/jHkE/+EQVBLFAU3W+twN+d1rBy8hqNkwm81Y+abWC22y09SmZOfSs
DpA0dDY/BTy9pc8q8nmJIBp7UTP/SKI/4YrBmVme0X38uc5fRBtl8zw/G1Ygtr1z
g6Dw7qakEycxS/RvP2em4U8hafySfyXoKhpxa2wr0DwSOzMCjkzOO+0SaXe6zArp
OaPs1nXPcP5Ud8KKa1aU9oE+72V+PJaWqGUWk3CG5RxV9K0UfwkYgHsS0l9lItzN
EvRlnea0UlYr8Hijlp8Beda3HigC90EBCH/nkxFyoMtLXC11Q1Q7It/Dk57YtQop
SvcEmS+iu/kBjj62UFl6nGYejOzllM0Upanh/Y1LDWDQWPWTB+7O5hhqLqQwlz3Q
HlW8hidXh90jk+74LiRWgpIjqRoUdqtOid5G6Z31bZlJ/8qdDijFtVBYvSwkx61c
244+hqRsfpFcRKzJ7PRx0QrYwk7OiR+4iIfQGx2ZW0tZv+RSmXt2pvNkjMDqx/5+
DC4HTyLvcKBOy9aHorAdpmKjUo3y+xPKadv0dpWKxSzm14iSsG+eUWp8oewNJDIQ
udTbPnmFBsd/G8DQSORZgDqASHTMjDAHv5pfAJubMaWuA3Q+Ii7XkyyKGAWUwvvy
ZOusjJHW3G0xw7IDIY4FE0sE8cML1ilyTFHlqf19XPsw4Qa6ZtElYeNidpwMbrDN
4H5I+hBFwUvTikJVCinOUAa52bGcsaXMBzLSIeTem2nKvJLWZjNva74snBtw2ZrR
V8zoikYOcKiy77rkLzWwcdIE60dkSq6AwtWlZSzRtXfwcOO3aIfUYaeelcZ8Vk8y
mUlr84DMNQko+u/W28PKB7AyJTYP9ak3a+IcqyzimXFrUi2WkZczreMct3KehtLp
a2pxZw43FqLbXQqktm4JnOk6UobUfBYfJX3n8NP/8/bbnqYCLlNFIW99zu/j05rP
9hO/obhl+VOJvY43HRNBwiEV3Ftb/DJH9uimQGwuAw5drVfAYwG/PSX1hrnYkBLi
ru0ZLbzkjm34eGfwcBcWLMGA45QCT7aIW9icA/ct546DbsHpvI21gFVLCZHtXPHJ
fcRaUVmicGxhDBoVI02ZtNb7Qqii7096Ts1gRUiKZz74OYiw4ItSC14MrYDUYUEg
fFz5TlR4fW/2trfTv1UmFFO7ZAm6lj/2KeEvlEmI/eBWmrJGnVlXSzQlb1KLl5AH
98QgQpnndmj5bfkmlPQmB1OpXU2jBpBpTG2OC7HjPb316Vr+WvUAjh/qynVf2KQ/
mHa2n6qed9o95VcdfqBQE/jQE8VBJArZ7ZussMAwW8FRhXYUpDkZ7o3SYLNe5uWp
ZGOfvCdqQnm3P3qr98VlWV/e8wKeAinKrJOqvZXVaCKo2vaQ8mPkU0PKc9uXOA0q
KSc5xzEftLI06XtgLBuZpv8BU4xz2ORycfPpK6cI/sVDfkQsBla1V779nLs/fo/J
Mtf6PpNjFcHckSfWzQYlQLqEgy6OqCPI//9HRfmiJIyG9pzeU3vwsYoC93oE7be+
kNPn6yXGUXQRlN/G3/c/cpmOeX0ZtKdsjhOJ9dehwdRe7bO+D6Yeo5D34ZWonLDh
R+OFphjzmm1AJAUPqnv/KDgOH31Ld6lUHb3vRICT788fZuzn6KAgFHrgc7ThWUkl
8F+jbZ8jBCcc0LnL3gXaQxXxNJuGq5lW/9f6K8QRAzTCWQad9VqHZCoskOuKgWSd
XMFd3OTwRpj8wbHWGzhU55VAMkZWQzvLFP5hDh4Cfkvd5bIn8vc1y64eOom35brE
VxhJnRnLFbczm0TXxQ7ld2ccoAEgT8SoSJ9MXlYUuVchBbggKhyhJorJHRIX+VwQ
NWOi4wvgm3vt4FLwDBDABqqlgH4f7Q3wf5Mo6DaZncueLsxHeLVbNvjhrWa1tUwP
s71y8DTMOruTaW8/TWAOnWfbWrAbrraddb1FWi3fHCZHxYwIagepazKfRZi8R84H
3s9ErF6qloIq1rJ5AwpYebuuoO+xWbg000GIbeFFjr3YmKZvz+Ud+8mngYqVVmIJ
HgOBEywm29eZmwhmMnhbzBh1kNfso0pcMMaJJK7dKgGEQshPoaFkftmAulCHdaNM
r74NjFkBpD4U+E9DlmwznUORXILv3QeW7Fy6iwaa6Yc=
`protect END_PROTECTED
