`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y0/kVVGYp0AjXXEWBMjTv6Ff/sNT7iVvQW5ON2iRAeryaN+AB/eQ6PQTFn0YzVvq
J8zt77j3tESAXkXgy0yfzVVk4EHtN67cO/3uZciyTQMidK3dH83ad6nzBRAO0iqW
hPscK8+zAsA8XOydlpbFXilbfQ7nfr9nHTEOSj5WWO578F533wFljGukOPQFyYSD
9MkSZKLsZo9XfylOBwydSDf935CGXGHbQ1NlxdWcwf+xwCqvFI1LOg+rSFvt6Dun
ZLLMu+rXjajfzgym3Z336tJ3gx2WcpmKBlJsEan0L82nR4x5CLfDd1aI7XitpZ2a
v6Z98HyBJMtAQx3xjt8um3IA00+jNSDW5TMTnDboOrGLSx/J0zTYIfebz1Kzw8ut
tbtUTWExWhiDGFVytIWeQQ==
`protect END_PROTECTED
