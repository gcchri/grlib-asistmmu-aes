`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7EkCcOHVX1+ujXWhglWqj2Bv3mkJpPvbLe2iV/0GxM1ppR/r+kqa25kPTUZUNgV/
vbLAvgzdLCo890DrPYX6BnpFDUZgOwAyB5zm1ostfYoIoFK+CmHL7IfRLl4k3omb
nKu8twTeeg2VrFIt/x2xVUyaH1N/FBMakDrHqJHR2YtBNf9u6xurLYcBwNM/t1z3
wuUAKPZ2syZPScCvnrojn4OF/isaMD3CxVPc9bAbWIIP6Mw/yjXEhjGhYxIyZXHL
3OIgOQ/i5D/h9lkA55GYba34Vnutj5BWwfDLInOJvTB9lyG6ZA1gB7WQk7dMYZQ+
0tAeTjJ4o6+A75oB8JjY9JlcW38RzurmItCPyC2+T/rLH+mfhr0ZSiUgRigGdZLB
KupX581xQCHdUeOPd8F8TtmxuhCPnd88esI5KwZgG/BaiJLBg7HpJ502L0Xvzwap
lqsw2+Wr6AdnqgfnyEw5B5rL2o+5eOlQiYpOGMBD5T9RxPATdYExuG4z4gsCSFrM
PKYNmTdZek6l8uQT2oPCkbYcyJ5fJfqdcDGb/fGodjSJNMoMmi+SjZEvkh6Pp8o9
1JkEEaSI2lPA5O6IDKxO0YUBSwVOj4ZFR2vdYG58ck5J1STi77EIoPK2RSweMHRl
`protect END_PROTECTED
