`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJW+FSXAJUxmVM8XIn0lTMg/ApnAGkhCCrRzayyFdq8y4tmaA6dZriMRhkNeVnb1
nw4Pa3TLNnK3Lw1b94/mYLB48YAO1XQtCiyIAOHUdhw1z6AK6STdMDKnX/xQDvVo
9i6Ph6Xz4G41QcA4UoRtDKhQs9LSE/scyiZ3pl4+2Bx/JomgozLXYtdSwjk6PN0v
qDTAkkY4UQtIDVK4DgjY1ndRe4jTD1MH3cRdx+Ut+dH1MT1Scfutom5Oo/tHBIA6
yRfqLt8satiRgHmtpCHWHZnk10BMgbs9NaCZcw6w59nt9USQFLkH4gaa27DkEPJv
Cy8DDaNSPyBzB/Iq5WURVIxOQobP/f1BA9Cxcglg6VwhCjBZD8e5hhoyj1sERdGp
Gcw2NAFLcDIjcUItuGzR3geltD6mxLu3nBcadJ+sTO639dLLiXSH9+WReT/C+jjt
DSs5bvTdDtGqGcnSN3BiKFVtVrtIU2TVUBLPWMrOmtxUFfUVvJqgs3AX8eiScEla
QhUOtIk+i1DksONcayPh8mEkUndTs9DrwNJ7+0nZtVR0GKqlRXh+2zxhsFgGCRK7
tRXmWrwhkvBDBeTMV+jIBaEv2MZHX6tu76Tko9WSBZwRnogVYUA1uF44r0n7hJw+
h9sxncgfnGmSENttv7lSdGnZCBgxsnImyc0J8868Rvgt9mnpsOheu9Uawz4GXvmn
OYqAT6IwnjmAIZPx8P7X/r6Y3c0pOD3ol6rbUnyF50dj2AOyLe3E4MpmDS1P15Kd
k1IrC3n5tcyniM61QzmWXEfnC5HDKX80QuCRh/y2tH8J9Hlu3R3raEc/WD57Bt7t
lxvl7fFFASMaWArSdkf/XwditqbdlW4vMXBqpdi2y8SOm6ABvlU3YEs0LdDCzhx6
QmJrcxd457D7nsDW3NG3Wz2B8qKrQUs46fk3zbCUSVE3RNVyjIgCHt7WMce1RtJd
`protect END_PROTECTED
