`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGLBg677M1D9XoVNA9h9X1iIieHI+9pqsv7yny/mYnxvjvUujctIpNLzo5kUZ5iq
4FrgkLKSdT7YHIMCJMZCJxV1dox9UK/a9/PRw7htkJE7sGO5pxWxiL5qJZlkrdlB
52nyaFiMryzR/mJwN4Qc1fKHmEWKY7n4YympywPZKyUKMPfT6iepo2k8PuO7j5Zg
12t4XyvnOtRyIGGyAbhzMBgl30nVK+OdfwAV7BhBsAgw1+BOrErkC4jbnZScanGm
FQVf1f1HknyZ+oEzrh14YCmbBdKimzIYYLpThyf1pevSE0dBJ5y9IDoT/lwIvbmT
Yp0us1gl3jnyQ7f2CH0jmq/6raaZoavuYBsMwXJ4pjK4WtB8tOi9lKvHZfWI4D7E
/PolBSsFFwZApJ78J17I1aCNIVjlaSVvnEx9QFYXcszthg0JZC7jk8fXpJbmMxMA
`protect END_PROTECTED
