`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZzWmZXr9AbCKzdRMXRw3ntODJkDGhnxkNh2bLtShE6PENjeAmU41iNSYBIc20BAN
UJSEAWmTFa5+HYaiLdl1XFFoNBxFe9KztCu469kWig/OwcgTGnNOMGTANOUDOgPu
r4A0Ee8srsY+O4NnRd7/Q5SPM7WyZFeW3J8OSoJWdi1EUKAGdodwJANcZav59sTq
2UuZ4d/jAgkKDWDPJk9ezScjNQDUMCi5nhD1mBVMHv5F5aK6iDE0zeZ+bfb0Wzt/
6q+XsIxFIpZy71EI0xAKLel5eezQ6VNSCBvXy5pHFhrjokUBBIPFOilKaXDOqqYH
SVS5MWTprhABKhsz11IO1PGQ+TE7WSqQAvSW8Fz7lBmgbtwl7m4CYl/dZqp7dcIG
DEYduv6Rn6s1cTqfJQci56w7PZRDQ80eLsotfhIkbRTWWr6B4gPqRYYG6y1ODRsZ
Av67gPaVcwkWY16UAmM5D9lDk8bk//0CCG5vWnwxoVQQZTmpnUboTV0YP6oiwaUV
sjHxhdYgjtC9zIy7jeKaO4b2p28CqaTioPuTFt8iQ5ibdjEAdxll66ebxOqfdRGa
yHKYPdhMxRDhy8UX4cuNYxLXM1eLIsRzyMB6buHkxKAi8ytcwOQIK1kvRaNJCDz6
srKqJkwLh+v/5iQwqMsaf7BkrTfxSpYDT8JW/l8oI9HEW3vhzASohtZn73EHpGOd
VxwQlVl+FUzWLI4w/lhtXGXI1Ejq+m0ch3UFRpT5n4qq9k0j+cCVWGcqZHiNJ/cr
NUS4rdkxoB/932uxKfRDO+Tg+qRzQau3Q3t9635PbY18aWpG3Yz7tm/GUUHoJrax
/vcE7uyf4TxY8tsBYCLjhrUBdvzWUANnhaV98dsMZN2Rt1HlVjmN/JsDu6mJTjuK
yl0XpUs/N1NRXeGe70U6S8Fvh7BhLByl6nkUbfvFpMtpaGHXxOLgfc3wqXuCl0KJ
x6x8UaVd5i2ze2Qn7o/r7AjI3HqOHSSOp0K2ZiRyJgmG3QghtcszgjYCPqwIGECo
GJ0s4UvLY0qq7hn5EBcJar81SpZG37pUBSmeW/eplpangctNlgL8+klw3rv6rqNf
B7bw9TcGrxrAgz3rw8vzIw1LZRTpMzUn2xmfO7glHr6Cj+o09D0DYZp17dosupIC
ayRsTWSMJAu0uBZecBZezhfGouwoacxkUZEi4PMBK95gSvJNLn40UB4cgRxjDALh
rUPhXFdk87LtXdavq2NWgyAR9JHjFluR3/Voo80JdioXJLaISbSglzmvPMtLB4PT
8m6AGnHdEXO5xOmAPy6A26v+O5GTpkckuK1s5C1iKMmbOQGhbI0EuwmF748BITll
YFEBLo58/C9VVVz/uwLDuwlWvmI3ZGFUyIsgYOS0SRNzxr88vVwdDcI4WxX6BMbJ
d5Os9qRMqUuli81ox2KEPXe8rIgqJOsCahQTj2CfA5t3kXBFHsXszZsE/IKJdmBy
ddkk9ioO5+CunkNonmrZbX4bHlSefJnNdIMbvP8iDAuC4v93fzB/xa+RRX9Nb/XM
wVaImLnHzKvAaNYJE2cmqGknJ3D8OU4e8hbMag5ZiPZn83sB/lwLq1Kx/Ho0i/D2
JUjt7PXyLzfeYzqXAyN9ihnMX55DQBkBWzDn+DzClseMTQUywsuKL3VqdNdloHq9
Kp4hNgTUJqZP90bcdeXWfAX4F0eYi+PNYHHJZyHVRnrGGwHIY6A9H/M2TOxZ5g/A
JaKHTqEUCMmCf8QUGbeXNSJGB3FfznnHiBevfOyDdyfOnuLnVorVZa/XunQb6ZGZ
195vDiHW3ARRpSGgaomwjJCXc3dKYDIe1Rgo3FxZHTsi8hZs/fwKsWDgzyM9Tzk8
ud1fYotu70khrHCICr4071+NqL/u0Da598ugwa4o4iA8RyRxF0cIoEECw6U5+tuY
VkmVGiZgLIiATVmL45pEDO8AjmW4nwy0fOfQRp4UZpYr5QwUU/kJuaN4lrqXZWrx
8Twl1JUYRDx1mOI2msJYOqUBHxFYXOiZT48hHErbHz4LPqacKMzhczqV2CLcniUO
WJz34SCxHj1m6DwU/KoycdapUP2Mxa8iz9QbQiyw72yZdVhlmMbiGSag30NpZGlI
kK2fNnQhZhI/kcZ6CzWTWk+P59NSCgvARzp0AZAivC0whvvM52+AXNfqIjKQrS8Q
efkfsvtKeo0tPPu2Nq/DRjAgSbKf9h/nQqGFf9cTsT5fk8o7AsWSSDlTVTJJjhFd
l4APj1WvvHUTy6HYI9PxiT1MbWScvBAyoFXqlLKeX8OJmKZ+pZU70cGX0wBgFKZj
Ap5ENSbLfvkPzRxN4PJw+WnjGhE5RqVNt3SKqTS7WAz3ryyvYKrX4RP5alpD/6pS
4gQXolD0kPqGHpMRokDawzODCBNuVea+nmxryf+ESkVm3suL3lXRBjrZDlRrwIFB
96p0hr6HttqGbRd2pr8CoOrY4S37DyWfJuxuXd5Qb/7k731csgLKNOWA1WPsRU+I
iTCbjT9u5GarwfTmOPmXNQZhnhpiefyJDeDogGFEvm+bBR87YrFiQ1q0b5yZKWtj
rBJecaeYishL52s2blaVjFn7vlnhtymerVDoIqlfX2ac7QOXD8BANB5rYtVsiROT
XAm163PwJviyqcKDVHTfYAmq8dSDR5yws9jTiyIfAHrdAQOFA5tnMKfiujLuon2P
OoAcndsVInN+SKl4LAS9zkgWyOyTGbanQtoQMtRC4Gu8t5aOMPwbZfwJBDLSvDfb
K3QsH+n/gzPG3Y/JR4MgX3TkA1PU3fQDxe1trTd/rT2jzymdyvSPNqSJ7ieDmYuK
rnGhW5Y8FLS0HJK25xOu28MnLrw0g81MmHQ3g8UsyPw5NYJOBjvXvJO0txX/9cey
cdRRm0o8adV60sami4Noou8o03cwkA6XoVRRqD2oCRn7GdoI3lO0ew/Gi1YUcCpI
20713bmpogEmyUvvS2dx3qvJKARzMfusNXSV+mDWmAn+hlILz4KPJS2c8/7BNJDe
unxssHB/VW2E792644PYhHymxDYZnE9EsUSl7bwJ0Tqy7BZjmM2ztJ7AGp68shH6
Pn48/LnhZNcD14R6fCGAVMkAUBPejMK9X6DZsEdhGe+iL8RDefIt7rYpyVA/UkGI
P1cRuB3Nh2IacpVtt2FWCBG4fZBk5KoAzXXvAGImmijwgZjuXN9pePg18diVK1El
eP3lxMyvtUJ+z3UjfmiZt2slxmgHrDZHncgiVS5E5y7CDe0dOfbQus+uR7LHPt22
mHwbmheDbvanpNEGpm5DUno41nbY+oxaL4fzwRs/umMohN7HGbiC837nKDeeas5t
KLXEfGOj03RNj/z+PP1hwTgaQsQemRxs0vS3vJvE6mJBRVBF5v+TpZcbj2qi2h/V
F35FllI2Sw9pRwoJCUFHpoI8HDUiNnvhNjjaqz6w5rE4o+5cYZfmIfIL+Tv1Wiir
llrEogMTadwCcOc2muTwXTZ1vMoOflC2a+ToKP/MaLbkk2TWjNP0LaV+9C1rcMPx
POLWM0OBoalAjHEdEnx5VNrr8Dvm0VhnIwKq008CBMnqaBK6yFnzUy/C1MdVeX9P
Dw9MvV04//kW+nONK49jhDVOGsG6cxuKWsYi7pEBx+E+7yvMMabC06tHX6Tx6h0H
MNDGagI9byffmDWFPA30eeDJOJ0w9hvo77fyHlaYwuzSes0ZA8UxiUQOPmyUsNII
gHIrn9AA3LQRbhA2zbHw7hZpvXYYEGMvBwKVvKyHz8Xi1l9CRxGqQFF3tGvOF63u
1nptF/hI+G0etiPteTss0rRlPWGS84zPfRDJD7e35BpCiiS05uN1qhcWNhjZBWVh
a/VYWD+u+B2xBPKqafT4EX+LXSNN6t4RieQB+LkWlgiqpTfjPquhDT9NAprU0yrH
ttvnZwtUR1muKHpyhuYtJGq8RoZb8JjShXe53JapJnYfb9vF/CA/8jzJi9bf+rwN
+OktHxN0n1XjLt9mYAtlCN8+vmm7JYVPrVUEzb8jlBMTUl7PCSgB0nEEks+F3oZ3
jrpqiJHgkIKZHr7wzaXqc1APuKmTmOKtqHCFqdClybT6QWinRaihCWuoUfe191O7
pXzJu7KF7y+dJ5HId3fZdzwJTXT4y7HEunVQ8+zDj4zPlmE/5PIb7pAtp0EBH2uf
ue6+zzf5i8VWFLa5eFHqhdG+kH9RUZv4ftMkx8reNgdRtwc22oa/n+Rk60H8il4j
upehPRioXCxa56rTwud1TmlLzzgO/Kju8Mvo8emeRDdg6aeYPGZaFaGMUE5cg+f8
B8Amywty+1MxkdlUdYQ8GKMMIAljd1XSQUq0Qj2hcZXzXWIV5npMfwDjXPpOn0Tm
RbppQ/gVyLRZxXU2JVzLRnibnoyfpj5Jl1FIqwWLdPvwOb6D70hOGUWDoaoH2nQO
B7qscCga56ByOz7CeD9ubovkRqJEv2E3IgyjNqHQSuY9lpenX3ecvhhjk+1Pjy1T
/TNrxR9SOmpwxyQdZT2H+k0KJZ1WPcoNUftaBpGybB/A1CVerdhiKu4rG3utE5gd
SvdptMEUXqSiprNJ3tlcguCqxYKHWXznEhYvC5cnqZit+o66R2v+zKfkTtNx+txX
SxdEYmMa/U98JKLwxhRpRTpxohBaVznVxWfR4kxhDDpdo4ciVZDlKUSeAtzjDELR
TVgxf6ZcanznI8VhsDmveVFKHx1CTLfvTZX9lzRta2tdyl2QzXhjriUH+mL+WvKR
v+QKDx87uNmRvJGBoHLhU1nu/QBtJC5kpBfxXs+0at72Rhj+ACcd/AkTgHPtRSvP
lrL07smlYdO+y4Ymimvn1gQ0SQx3/q35e6QFJExB3mvcaaYYc/ArS072w1BxSXfN
b+lxV9SXXz3NgG1VSNSBrawG5w6v+xZub6GEw/xLxB9f1oW/zhOkDxPoRCyNnRCH
GDKNZ/Osoun87hL0gnxVmbRoHqtXrHubiJmAT6YBDqQfiUg5IvRYGkhZpcZqwsg8
Nm7d2pIf9lI1eI5ioqJU5V4aI0KUi0dAHjeZelGlK/Dsnm+gfibtenOlfVGWzPI3
b8Fx8BECj/s2V0AsGEbej7K0ZygyRAOhxdH1Qd4gYQAgYz8sYjX6oqk16K6nQkOs
A4VUoZhmaKTbsaEABaBOmXXYL+xix/xgX1cuLtYDw3pi2pa7/rNnTQWsVWPYRGrV
kiBA79SbjEcJ87maPWuXupKcPAREKbkoJfudJNHfq9MxIVsW73TCsJtEkQCPlIDO
CiZfKV3uJXE0PendUxzxzG4P16aei7UoTmXX4GrYzUX0LKF7b46N6VJo9/vHu129
+tb2djDCIYzuuc/UYoP/WBwmgAMxuxX5fHDmdfFA3fvlBY8gRtrCPKXO5PjqxEU7
pFRyyHhBN59hXaFLa7zr6hVrm95SlJQzt0YKFwWg6gIvTzumHLyKGMNLFMJ3asKL
a1vILlDmJDACzHhczbGc93f7m+D+lXwEP3LDGDJg03TLqyTK1kdn6JN6X6JASdZq
k/DQrusQEjYGflUqdJnN9d1fOyDiEbV5aI9H+mS+Oh7t8xMISHL/Z9Rr1RBimmNn
opg5dzrasJbenGxvH3iOBqc6UpLiuGou03Kv8TlRLGGjat4oHeny5vFUbG9MzI2n
7l3sOVI/NjcrzeyLHjHgzak3zM4vuuXGLxhIINICUszLNj22kQnD9MMw+R2zHW/v
21WFKXK0vpAn71ppGS5O1L//oM2ukvCV2y0Cc0B5dL/QEf7IRMMzvEo1fseFI8bk
jGscsYLvMTD89/TtyAgR4LngPFxAEWhVE+Q4+FYzfFRJ47jChDlQv3vvLwqEQX3+
diebSgCMligwCTgPSLeJ8w==
`protect END_PROTECTED
