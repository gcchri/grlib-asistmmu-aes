`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/CHdhbyEUcs95O8FBYL9H3wkgX2vqv8aCdVlRDfdb/l3CcqprTChl2eQGH/EhFb3
R63HadliTSEIoR48hGe2lZEkOxR2HWslNL0al3gIX/57kXEW+UUWdljMUeQjfZT+
iKvidIGGxJ+YaSEFwD9Z9LL5V9sd3r9U7YRUxemHW0G3vYAkGAaU4UwVD/lz4Vzj
6TtrsqQC7yqDDxdKLHp6lUR1i4V/402SZltrlO//ml7asLOPlhzwksjlcOv1WvWd
OjWIeKVBnaoabkHxR48n94kA5eqwMNAW7nLq4j6DDCK2BIRYpsTf96lNUZ17q4w8
d8Rk7b6UAMwG/cMtoRRjnjq0bGtpCHky5BGnnCXO75kSaFLZDhZxxPspiS+LzmsR
E+Qz/VBIKy4PXM7egoXiGOoe9UCnyw1FFYJuJErNa7DtoOs8HYrwxwby3NgDA+jc
hb8D6HYshal2giwhDKPQzthjwO4ktx8QVPGPbkVTPXseDxG0QmsZcsl5XZWuO/0x
SmMeTUWf1QrJ1WlW2SxzXJbcLKurx0oQ3DVzmoRCNaUcJRS1Vde/B5lL7WcZ7BtU
N5jiRqngAgD80CNzeX+CcMye/tn0ldw6sA6fSCbfMc8SBqtXFKJ6RBkQvPi8dRZd
mUVSe/3mnfyj1qe36s4VIDe0DX/XtNazq6+cVjRlqsLlR+PgMk7ylMLv+qYT7L40
44ilLdAPv1o19Y5WTLVm6eSEj4DUL84PCVunHQu59Mo54iQ4eIsfxPgSawJBqmCU
85+HvMbqqWuNPLfk5b8CosIhVHdjVGxBktTlQThNfMovdWVaRL1EFLLSHuujn71Z
PvQXyD1ZNUnvJucpWTBAJ3VEAoJnKWxfCuqvFDCRbzqppreqMlEklEpPEeaSBTVm
SeSCa3PmKCErCnxWspu4Hd+NRnBySq1pJ0K6l7pCpLyuH/+C65L91RIPOpcVldaH
hp8iF9qwNSIzKeGfxv1vRZ9q4mJUZ08rbO7uJl6lM421HFbTwKLtN4G2xFG+bZpi
mPxTOhGcLosYZ2iZZrC5NmQQ/GnDMdjq0vN3xa3+mlbd1At8fAfojsqXPPUu9s5x
LiwlUWOz+Z5IEt9sO6qU2+x0L/3vu6VJu6Mu5N+8N8aCnfBm9dhDWoCDuStfTcEI
DBYHwWg0vl+ms2ZtV8ahLtIRsK6IbyttkKrJ7XIVwFltFiIwKXYelCdcPXCQhGPI
mUoUVjBJ8YwPeZ9+SoE8axgmHTCS77O6LbISIySy/THE6EXaT3hdOELYk8nrdQr2
egmc4DZPi9QsWErmxy93hqXIVcYW+ZQ3r0/4ErlyF7oaW4LGazcWlZdbfrfraOs7
BUVdcATm+AmcLFVBc7Rpo2xtu0V/P6VJf9voMqP15pzCCDINAPk9A76n5sM0PiBL
5zq/8nvPHI/ZQsQXDm5b9OX2H1Maxg0H3LkhB/fI29aZb8XbtVNHf2GoIgXjl7vz
IKy9PV+yM2s7Lv9d5ZaMct6wKVO26oS/H89QNtD03quX3vAtePNCQrgCGp8nqPSd
twmibffglqh0iiVjnZbbVC5jcuM2hka44FG/jaFPyQ5pfsjwSfcZKC35XBGPdQHT
iSid5yJUVXIbl+ISF1CRsJybZIP1I7sER855tHHT9GcaE1EOTL/YK7miXeCUa3YA
CzhTo44yh8XX9dEcyFOUl3a17CPaXR8xQRsAcfaPv+CkzKbO2OsScnP24cleTHqE
qs3forVqXOazMX7UHafLKNAcrq511nTogXksn8rDbC+ui4DiH2ICpnO5T0IVpW6d
`protect END_PROTECTED
