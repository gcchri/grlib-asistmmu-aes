`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pkoaaQHkksaRKyQRTnvvEzRp7+03hMsVcYayKJgP1EWoc46ycRkp3czm6snYnMma
U/FISUIqH8x43fn2+Z7IDH1TJjtn8V3a9oeuyiuMKLY0RpVgz4onpgdnud7oneAj
lkJg9sQBtEJX2YaLnLxYfkBWdf1LdPfooFGRKjDynhZkcGv1YtsrrKFYcEEOXw5e
ahrLHd4hXOTwLJbYQ0w+pQYOrkMoLRBM+Hwwy1WXg/sn87PCZ4fPcNmDNT0Sm9J8
KhQsrMSszSonJEb9cLtY/6PVe6z91wIKunaTZzQk0T+2iBdyqbfq74FO6hLWS8Xk
DoDQBYcCx4Hu/DQ2I+VSpx+maOwKt4uVLvhOK2JALi3vfAKqQ8n9u2iN/W+ashLn
6hkbvJ/JJzbM2nVjDe6INw==
`protect END_PROTECTED
