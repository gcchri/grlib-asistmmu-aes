`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ymuvV+n3vPXgJkuZz1fFKFkLvNFVmPPzkEYuLavH15We8nO4Tqr6DZvuetrZif98
QF9B9Y6Dn9XajznVcUpJNjVxD8maB7gr47Eg283GvfUr/95yyvdoVFMLvNDNyoE3
37UsvGxqMB7S1nWtYfBm3+ajqcYF7bHQvnN7eyvgC73Il8OyqY+Z1sLr7BC1J4gP
Z4lHylweuIlLp177Rw5Nmbr8GDzd3qZU67DKpLL8b/i7vthcdfMG8ukEWJrrwHNT
Kwd4m2KePPxFd7/fX5qBEvQaf4+hasLR2cYUvSGlyltBTBYoetpFDKh61tQttHG7
a/RAQmt57sHFxpBHvBMp9oOaAhCXIM7psQXvrYqBMFQqJOVnD+JpAWDhO37EtKr0
GRekrS0Ye6g7nDu8o8oEaoLjECCb7RtEimA4FeF5rm0WZIW8d+I/R6EYVulu0DKl
qvgJ4hrQhVPxLLnbu8paIMPEPVMJl32v0o15Rv3/TISivO1YlF0wzMtrvYrsmrxJ
7Vv6x5lJLRWBi67qdI1tQImzrtlB8nn27m6mPnFNNMVgq1hY3lIi+PjI9lz9Uo9O
onsrzCXvBXE5vMQCpjqo4nfdJ11W8S/K6au/cKiangkj8zj3zxHKqJKsnY7p555o
eDEn5wcvHd/oJuJmQ3R16NVcLq5tVzc0fvU23kLWD0KwtzfgRkhXN/soTIf2cIf7
yfyhUN58UpOBICjH1ZU4Uz4Ogrs9zQXshdkzM04/ZBq8woPRN3H+RF3ii8SG7jLy
/80rIlefAIcYvCn65bqDgVCEh7XGhuCOOfYaZKGcg/A1RKVlCG+ORlF9ClBVxfVm
Ptm08H4ceWfzdGAlPk8A20UhxwGqN1gGIuh5r4XYeyvR06jtVMOwaaA309ZALjLo
4HUKnBct+MRQet29p0zCyQNFODNi3ZFt1z5098h4yiv0hBtdBJLr7sQXEseIRixe
e96jKHLQGE2e0kD/9HzhhoM28oZOnLSjKeYs/rBsTQU=
`protect END_PROTECTED
