`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUx6uXho/0lcA/QvfjS9ta2s4uK56hHCi4cgTMvdZF7Ab7GH3EEm8yzgjNurULKn
o7IsioIxHERLxm3kDldLT1vZ+7ataSkuzhdN5COMSB/7P8mH+5+d+J8A+ahTcpVa
bxh8lgZErwW1KyxMQ3I0sDUiQuoHUXwRdhqe2ru5zgULOjBUOyALthrwdyi3nBJl
X2mS9zQV/2LC46MpTH1sL8yr8ZwsBKWWJusoRQ0ZkxSNJjUWO4YbLelXqROcceil
DJsMkmrEhXGmIEeYz1OaVYwplwGeRmylGulsR4/bqPc=
`protect END_PROTECTED
