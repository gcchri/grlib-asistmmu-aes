`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
001S8CI5NrxjGCm8fMPh6sWDFBTvlAVrPGNj9aY49XWqd6yOnC+1P3yuqssOudB3
IBQB8xJDiGfh/BCLQm56HB7nGTl+9tDA6B8YP3XKVYpcJbQVOOSdYMBJqVK+XjAl
Oke1O+HIX9/4e6o6qqUzM6GxkFSCdRPclvtVMxR06YBAPtGyrdnaT2SHFOlHdGAF
ahjZJKUF7SJXiHE2TU38+9zWE2eUZi+OaXGpmZC07KkSDor1eXL8uswDpVEvDjVe
YjQ/xDAj22mkYTzmvao/UvqQdHYSI4lJirXl125l9vEkXZSfRLl2Sgqe31v0URU0
pfxrV4+TljjqVwPL32Lezg==
`protect END_PROTECTED
