`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eaFBsUCulY2oPWOPQO3XPZfrryIvnI4kwZyuKafdGsoLZx2DizMgYb+VA5rlrKwF
zeOiFnD9nJN7Mm4PUBkOs9lRGSRvDaYq2Vvubl22bxqLrTE4Jz6B49df6yI0OvRp
9sy+Q7iXpvCawLVPOvduqee73UVRaI0iH4qFgQFMxZ/nPhFShjzYZ0FjyFi22azg
MEZBGNteKyx9mzGdUkbIZ6DVRtSXVhrpWqTNBosmzTs8mlNsmHs2VGMaPvRbVSqQ
duZm2rSZTzV+CqMiMzC3AXFJ9+9RbhT0xlFnZXoI/OIcELeIiGkjV8cbwCr+T8+c
qjUv4O22flDBohUP+9c5SdYLPLU9O79a4moruW9LcqijNdWqiUomsG5SptCuXrOF
enYKUVPj9HBxXd5kyGZE+TMI99s8ElgPQqA4Vba6kruS8HdMgxs7tjMIfHF+A0kf
dZT+171z2Zrw7NVC/keMGpMw557vSzhfFiFdW/FqYw1iXXOVnHQo8p3AjGj8oczP
VhLZTIVEMn6nVP5ujMiNZKyi/97s2fgauN/GpSw1nRLiyweG2+XaaWbVq+naFjD4
MmLvm2BVAPPUNquB7u4qvg==
`protect END_PROTECTED
