`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DzoTt4nu8T1WtRp5b5vfl8C5W6Ci8vJECWoqM8MmOlF0A5HcmbU7NBVt23JbWiSX
n4gTH8dPizQQXLIx+xeycNt/WxAUhPQ/b2dd7ABrmsB4L5VYbPlsiNZsUxpC73BY
Ace9c1UU6NUEjJFM7eA5ROi9T+Iv46xdLIp4u6tMVns2M7pkpnurFR/SE1zdum8Y
D8fMiHNNJ50cEVUhfNgewifHLbktNWjLKXfe5Kqr1u7BF0Soqp0sjNNTswPZX4z7
ugNiMYYk0Cc2dPrvx1FyoXytxiO6yj3hJq2L0YRJHedzKoAswC1kIEmKJsQNG17C
JiBzsFVJGPRaLKXQzwHF/b1sT3cwnx3xap6UV3A+EKD1g3OjOB2i39Q0H5ynElXC
C6UmYw381PCFFjn+x+YPtQ4AWDEUE7OQiIajlK4x4no8AJxgpBkq6obsXofunsNn
wCRqv2jobNk1u0yXn54lVbVko6fGh2pwe0D8Z8pd68VJyGDoQnOb+9CrVtiTVWLU
Pryb1PxpI3HC9lcQ2RXPbyuPHrcRyxl+8picmvhQcY6zBTLfXrmlKOEEwI8sNbS8
E0YczVhsBwrG/zi/wEfkPRZ8gkKekiV7kJ51wxYliMwU+a3vT5ElYZ+NpyCBOFVU
BN+s5oVKeEwpNBa9jtwpOjnOG74gXAd0OwpN/Cy4V2FsEbzR9TwcndJYFCRfwJsA
7iyww+HEEf1pi0zXyEpywAU6IlOL1OCLU/9YA2NPsAMiWbLd+9YePJRwJbIFM2tC
/aVPWGP01+pqD+J9H36QYMOxB1RQ9Pd/oE6dtyIyzSI4mHXJ38TiaiLP2Cqi9i+q
HZdnpCxgG5APQHUMZ1WFSJNzk3sUQ3svtqkIXbievmF/br57aXCAN6TMGTFauWV8
xab3x/bfx+HtRpwpPMyxquEMHkFHTEPqMxMTenF/hEo=
`protect END_PROTECTED
