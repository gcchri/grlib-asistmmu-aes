`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ySehFuNZS6DMbXFnMbLDt7HkuD0Fe11EKge7M4cRhlHzZ4lAxhaD84chk3K9Y/oH
UzEoi4cYmicHfkPq6uZ0Pn1mS8HFIP3PFDgQApiOnmAbJTw1WlkHArMiu/tkRNzP
8OVBN7wQ6aakEEC8ryEZxZZYkVJ4jp1adUpb8K/KSSCW72e9M4f2FA7erAMilLWh
xcMlS8SF1nAzVYOdWOy3S5fo1YpZGY2KqJoIVKEnysnLyhHIGgPoKxTh/XxbrtjW
bSbkTMGDoLefkFViq5hLfePDCria12KWPCuW+EEKoCstTArq8Lqz5JHGR0cg/GRO
A/sH2SNJdPyVO2aojYBiEEYD2Yv3xwHSJ97B7bv5V04TRJYImqbGB+Y0oTCmrMEC
2ULZgNqBQ45xgO8QQfOPkKfQKqXzgDpy/O/kwVTO2JscrQg2090M5Jl/BClssQNP
polM1WumTRVYc5Rlim5me/tt71dTcOay016I+3oAUFwUM3NfRM9VM9eaGfE/cUjA
8EE2IS5yNn8MDp/76QVn41XruDQAfzqKuq5bPeJuKZHOY3G1OPrFP3KDVHABKPZd
`protect END_PROTECTED
