`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/llOrpmeDcT7Gv96GIFn5QK2cd3q159lqato+UU7qCPoKBxKRB25JzBDoj6DWKFG
9W/k2TYTEIsumeZl1A6Gn17qqF2yhWrSVy8Q/DABSQTT76j1zi3uXMgNk4BiIfX1
zgU9HQ3z94MriFmAlXTRiJUlVpuSHrw/tGjaY+do3pJk5TEpvi0pZ3SFl3QKkTke
aSP7x9Wajoqq7uV8B056BT66pIOghOF7fKHDc716jRpE1KWs9TbHbmtx1u4nDmD8
sW15VSnvIeuOL41Mh1CdEo1yL9LTiIkrWsJnQOwSB5EzNOIUN146rClPtp0T7NFU
953z5D5zh5dTdsgL7HkME6HI9pUThrM39h0CZW7dIVYjHtu8w3y2XEaI85d1tu2g
nzuGSQ2tX0O47LNhiV8puhDWRSVq3XrJMrh++SBxwebjtMKoQzQAyccoQrS9Sr4t
tECx/52kjbp2NooLQ1YDPbwrKB0MSutwW5T8Z614dgQ=
`protect END_PROTECTED
