`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZUPzIIwhHpd0wJ8dKRi5attVG9wWiVIGj7s1o1ZvPdUp0It0qELWyH7cIZAJUCLP
tlvyJb5hdsg4e6z5bvCj4xRVjjVWE6WvwSzfun/BYKcT9YbhgcpgROH+ruOQOAGO
JUwyHC2zvBYsI/5iNppx6jyjVcC3FgoNfxqWxFnMLHtjXa31QO9VyxTDZGnnoFAW
fMo2v8h/2iaDSA9HAP71SlTCU9ljwx4ErbPqZOL67a22VOtAmBy7XF6lQ+NipWPk
jbGxlIyFlBVlvhPRWSWH4sJdRWLYxRAjaNN6i8C5gNUNXfWvXFkEiqzrINqaGUXv
wMrk1mIJyRu6UXkCXgYpGY39Hn/JcOrGIWOsCkdLU/mNO0iYB46INytmAU08sDas
aSRLRU8Bl8FNM0OwGJA6ROaK9d9SLc8pPapogWfS/RLDmF/sYnNf3XSQtEqITnPX
`protect END_PROTECTED
