`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mNeU3liMEhzienw56HHm9y3DhKlmlfeb1z+FAETMT5cFycKAfNALFDd3x7SOphTP
9dv+aoS7M8n0p5Zt+LEi3WLfPWZdAnakuepTQsPnyfGWLoH5xjtiFW7+FsHrrJno
u3ko/AJqMcLfH3EhBzeXpoxhaNKjriLTbTp7cohTDfJFsePGTHaxMV+BeGmuFv51
F+xKvHNYOspao8YG8QNahf3vja3SmY1WQe6hqzsNFs0fz0YpICLLcsgxLa1AMT/c
KsSlLwUQVBfYKjTxwVCaEA==
`protect END_PROTECTED
