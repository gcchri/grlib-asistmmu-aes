`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CzuCPiczwqvXfanoaZcoGLvPcZQp+mgB2kSPkIVQqMp+aVU+SKG0q7RsWZ26FB6c
CxrgtgHINVRIjSoZLHnr8tcChK19WzpZ0TARJNcOSHKDCZgbRxpkNqyYAeuGMZV2
+FliluhHNTxJlQvo8yveyBWzsaefJhV+WdtUfOoE+1neRDs5B9gUTsbelFjer2qd
4st9VgL5CSsHvw2ojep3XBwbPhCAMJ/6NfdqyX40n682GrTs8zNoUIHl9OC9123g
89F4nhi/cHc06vpLAqVEKCNnwWj0kwZEh6c4q9bI+fZT5vvBo62Ek1SSJqNb5LsS
IY8yeGOsCuDdAqT3FVAp360xZvO23GQ4IoA8nf22GOO1rjQeqn9qwH6r+hwts/RB
SJoxZLqiz9XFInZ63KlErmL88G4KLmxb2gm9Am63wHEokI5x4g/7ViPbTbpfGph+
jI/g9cUGMQGwZ+ZHOlBZ+L9ueEAk7Egsv+td93c5b2MKvKvXH+lk7J9274gpmvo/
2rM9QFcOqSFzzIvKga6jrfB/gmErjSLKnnKvxocVEumhXZyWJztcHzc9yp1vqBZZ
OaVkHp6UgrlTTBV3WBUVUNGtR6U75QjQVNuGGdg4qm3ZZlmYoBpXxvqEQNNe3sb9
+ROFU2Yv/IHN0SVxb9x5ZLz0Z1cxokIdRRbAL3OxrP+8XF7I6JxRxG5VWF+diwSx
x0Q8nJ8TrpE69rVBuaT9RB04PB5s6NfVD54vgVPLa3VKfwGTXqFW3Y9CkdtQbBmI
Unfx7U9H7S+xDFOLpDG0Jnt5rp9P+RPX4MvJBbJekInbXciWOcKlqu8SyIKsQsx4
WhI9yQJFhSrSImuHDRXYDi4AYKC15CNstsNvZRU88qk=
`protect END_PROTECTED
