`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZP+MfsdjJ5Y8IqUoYUPB0JL/fRPQOWSf89mVnb8q8cI8UyieXIMynORZsunnc9Sa
TwVvlCbXBH2s8KohoaNc4KrgHtQUHpdq6yfMIrbkzEkwcfAWRKTc/c/wgcUkFGeq
nBBI5kmnlFZ/EV7iiAuSSqtevx2SOOK0fp+PE4jccngdohtEFVIcIYKgApTgLRkN
59aVU7GMamr1Co2/tjHIbtdb3PU/3X2/DIFJeWJCabkMqsKWASjPBrvDqiJt9gd+
Q+EC+U7EQP143CTmQvA1KJMaq/prXhaBcVOt6SdIP6hmHk3vNRqVxHzjQmchKel+
mOD28Mv3ibpY61KCy/d3VzdD7cyDkghMEZ35FoLPbWM=
`protect END_PROTECTED
