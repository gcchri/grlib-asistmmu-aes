`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BqKNSUWM4jF7/f2kiz8NA8THXekS/MYOjaeFS69J5NRhbCNJKqayQ/I2udRLWtpv
uoXITxv7M+FDUKk+KBTdXUnQ36UdBNu+EjYhrCcGlXeoYvA8uQMoh+74p4m8ZQWw
KTjvUcTM9JaouC7RLHNBMS+3QqK5Bcz7xw5QJ+4zbqMbmNs07yMX28sPn4qrf39U
eVdvvtYrCTRlG/Vw/8dLBqLDDVXs3zBmDAX3YMWz7fRAzaFsUTheVpPa4AyaTJkD
BoQQIEe0B+TUxeaH9C/+EYgB3sLH9J+H82f8pVGnSG44CLCWuHAN95xySLkNNvLq
F2RQUiBxP9hJwz2LPZN+e4IHeBOZcAwMrIaeBUjHX3px0IZPvnEO/14R6oSKtM4E
XVlXiI88O48Rrzyl/Dwl15MNAufAtzj897K2pzdMkt/riW1W1oXtV3VvZztt2mdn
WyFyjLQIaz9XSz5GWPHd4vEkx5IjqrL/zC22xM4YisoCT1UbUGLREBMejd8mGhn1
9PH4t8LwuQ+/Zseo3wr2eIDrVGBS9nm2s44/n57lqLg=
`protect END_PROTECTED
