`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WW0vJCvRHjvOFEQi7GSF04G7WslhOPXhGCQAvI0/6F6MuOs9Dvm+6QP75fgKgpQ5
b148qhZm5FunpCm9XluaHZSfjFJkKpjjPouri8tw954LAEWXcBd4DsSWRJQwGnl5
MmAhyZs8htbZlsFNGRMVKp7LWQvMo9zEJWt+itwPms6GgAAkNCnpYOVAz8o0onH1
yF2dw6M3qxEZpMyP9uZw9nL/aNGisLsfVnx0r6JCbzgmb9sR65zPi0HOrWHAtip7
lowImhhfj94QQPdHcXZ+twZAtXRDqJCuicT6Sfw19zd0pwyQV9JgTX1HsF2Bvuca
N+yKKbNt2h3mZotYSkWsLWgs2ZMjVuptwD+ZRKcVGcpqeIJCwTW4DFX6eTVTpIhX
wzuNwwJfoUeePq+Py4HJlam3vrXp8jcibkYrkDLYboVuX2HKOEhMfqfZgya28BZl
si04NqtMPJtut4PWUaq48kVCVmEVfagwzt97hZEJcq2fbn/jRVVjg5IyUkrEw+hK
y7wSXnt2ilS5l7klyH+OTdNLse1tSbKFVo6zu8JavRjAxyx715HoNTj36DeWSDKF
5VFOlH4l7kc5Sza4j1eJojIKn5z+Md6lH8IpVCMTSl3whLrASLb9ZDVWAZFyL1NF
+FpeGDj8pU8SfDhDOwXDuvMscvaE4tQByk9MhfTLqvn4TTMLEBs696Ed/CwurSJd
`protect END_PROTECTED
