`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QOFBiAWV7usKnx2LbrPLUHqAlDtl+0LqQ7oZ5Bkp1igz+irL+sNapLXfWhxtAh95
dhxzk9KKNyNYXtyrb9d//C43oJPMiYDsTvO9E5lCxxOVJMzHvAHmSSB3uCScVeIF
f17aj5AyRx8eX+csK0+VGJnktWBuv2QnqMxnOTPb1Fc5Ps4hgbdD9mCddh8O23jX
jvvdwQASTZhngxZ+Up4dcYSqw0tvdSXEncGTSUxbxCfFXOEAaGU6SIjj22S7BE96
trllvPSbFJaXYnenB7bKJOOS0haH7F5tNYdfroSkPlTxAzaAMUgQytDK+L4UDYqM
cmYzh093CM0zxEhWtwTlqx/iRV1UD8xn7zAfLOwYtDhwWgwOI2PhDt2J0VkD4+FJ
xTDZ370wiuhMgnqxXyJ2YAl3t0OYt39x4hR5ohCCIZj++SAWRQFVgmX1yo9+oqER
k/XMneIdgFGC2Kw0Qgc9+ul5vukr39NsS1ziMrbQbvosQPhdja3ZSrLDYZLJh1qr
2ErYISNG6ROBltimdJl04xu+J7lRsx3RcpiTyQEWomKiVe8LOgqf7L/AiMlzaMzk
YdQ1w8gkdaRNQummhUJAYrBZqbJlQXOvnmnenBCgV/jPe6IgwshRJZGdY4f8O9g+
1FJswwzCsuGCabA4Pnuv9eggO85fQ3P702AeR3f9NwlOYmOUX5YXsRuKp+pm5B6A
AO977zsT5yg1kgMIaXMOTezgTm03lYhGN1ghIUTUFOMXcfeQQIEgVeAEFlAoPQ6E
onFlm9BG1dQ8q5K6nS+UbmFRL9zdvGIcRqHlRzgeJgGPc+wYXn7yVbl+Ywi9h5MU
`protect END_PROTECTED
