`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aAZWSvjGTNRLBPCwzHFpcqZxaMKa6yeAycyutXusf9WV8VDv9vZAPZYOvDfENczP
ImwrMGPmbE3T5jULZqpDj53L+9IVJk8UATEOP7/c4a1J4OPKJ+075yS522F1xkBd
/RZLrAstKQx2Tjwadtm6p81T2xO3OcObqWSyKOi3VSiHzJ0DB1KxFoF/NpLdMZXn
I6Z4nH6flCVmXNwl61i48Fz9dHL9GUwj0OcbZTBUiMza1YSvsypgDGb5o4ymAuTo
M8ssS+82d++0mUooOap+oRRsX1aWhncZzdURVF/5WTOiT67O56sXo7A7OWQ5kbJt
l7f5PrKLB0XSTBmLEqMeI4N3B56WgUTOJWmHSEZ61OpiWX6bJSZ8MGT+2a2uDM2T
FCckYL8VA1BQ+UMJYykH5VYr80pFwvDOP5dK5MwX2XXMxBf7OBnKdrf1IA4Ch07j
oo+cWlL+VC5Isoqnir6Y6k6w9BrXc2nFksXEn3gNfG31dajyol/tAaXuXFc+2iIw
tg8el/0h64VKc7PhPLeeCS74Y3eN6uQtx2TfjCslSWXK38Bqlh5IaUyrJvRhPGxr
B7eHYwSLAdTBa459R/jX+PFuoeZyvJhkIVn4jqc+mIywx0b7ImJISlv3QhHZ8vVY
dsjNfmjkIzMHgHl4jW1u16pXoaSMOtHKNBouYiSJtL7zuzoLNH8n1qF/B5pJwvVu
S3BB47n5xF7ZLOhWpt6vflpqPj5voBakNF362DR8tE7j+VmAl5h4yqUbd3uR47CH
T4AgxiyJwtRlPiytkqpLnA==
`protect END_PROTECTED
