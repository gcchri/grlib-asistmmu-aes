`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w80jF+riaTRWEryq/OVL6vgARFWkwtH6N4JRFMdL/jRZCyKwqKTpUL/fbmhWrHy/
8WZk4IbqCZqTP1XqnsTRYjOOggft+hmJcfTQELFlc72a8+Zs6UfO9/d0/MFk1CR2
CW1YxBH/sRJzSx1m5vT7SSq7aNpoLERuVIL88yLYIUzS5LzGLN7PkneYS5ix9MUW
Gnz7QtBevAPlUcrEB/H2bw/yLyCIoP+TiAnzJml9yMd9TE7RHm9v7T5RQZcT9OpF
p+Og0tAMUpL9e/ZmXeAjaGAB+L6JiR0vBABM/pR0IWRe6rRi5G5mrz4Vne53myHf
EIXgncM33L+w1QMHEfRIQK5l3d7jt9cp5+SVwnh+waV69JT7B8ba6mzYwWEw6Y06
elcZhilZ8WOIieYKwUqRRsCl+iEjvQEoZmPtk4aSMSYDMeOUPC5IeQh3w7eF19UE
RbW2wZBWMAYlAEE/EdpRV1AifUyMY2Nozr27mDu9Z6AnQlVVyq3xQkKQ0n2mEGQB
eCawSEjYAEkY8Nvfnp14RoYuF+FpgCtgPvXAct+cdPKqlEieEi+SDgPcUZIz9Pxk
GVNDLo0poHOUwSbBGAn8zzIORUC2bWLxODAp7Wtc2JFqVwffTBO8Y82HzfrWP1sx
l5l6ElACH024BIbuAZ0ynVxO1dVwwuxTIZ/vYN7gtpzHisahK/982PR1Dv7xazZc
fVW2Itw09cDU0SyZ/m6y8piL5b6uXfb7UVcKwX70/lrwSj21NtqmuCo0UT/ceI4c
4pMnOP48D9Zs3pu+rph7b6jH4NX4vAY1wohw3ixZedQGZIn5G+qG6aAX+DmSIx89
0gPKmP47ac233nKlqROk7GfuA9pfSTQQ87l2wGm2c5EfeFJhb0S1TEaIDOhBPTt2
8erGhBQBYZOk+sW2+mU7MFAv+fuV1arfVOVDyS+g1FwSmCThU2uGKM/bear/wPRw
Nif2QgzR8BY8g+cA+DNnNAcpkQBfeuGeT1nvFfsb51D8GXDbSCdrCY07vNlF3kM2
kSjFLryNg8GDwgKTRBlKXL5YLgotKgAvd9XsC1EN/OMjWlGIhI5zjU5a0kgwNnD4
0fRnde/qGatlj4b+6U5VN4xkri81guZxLfIXVpkPpcn/jAj9GLfZvaCrC92Rw6oF
efSCK6mBqevn/prdAKXE2ox0NDteF7tWySQpKZfkYe9srtRr5QGGUWRsOPS/e5Tp
6dJFNgy5H5VMNOHwxS7lzS9fgZ0EfBLEDepX9xG+PowZosf0nUtSKbH4AtLMMxo5
4wmyHRjhjvCrWvNLu7pXEX0HtppS8DvCBE2oZFWL4opW3rHq4GStNHAL+MxsY+aR
0LL24eV/2C7EBoTP/wCoeJPUN6S/tAzumezhPoO/BWsN+g7oeYeM41wLdB1DZ6mY
owI7JrnirU4UMW9HD/5gk7SN40LPrRcnOugJ/F3nEJyXB1ejd4UfQ6o3nSagRc6K
OgiDS9xNr7asryVilWJQV9mVKlZxctcWx4KbXlTxauPZMgt4ifsAmhzrR9d+h896
G38/Fj0g2n0+X2wbCqLrDm3kLKOiFG8XM6k6XDhq1Vaw5heVuv/56nCC2CBLTn8b
pK9f+CyYYS308T+O8ruY+oHxuJoi2nlACeJU5PN4lMGGrp6PozVnrzVu2J6/4hW4
UxfGwigcYpZuW51NyBB7uj5nWV1CLFAwWNYqVqcnmUYok+eg53rah2V2IQngRMwb
mZg7OeAmH0M1+zb8XW0qfT8JAdlcE64zRJuPleLkkIo8HIID2c6jHjMjZm2KOBBh
ZClNAnU/nGf9F0yLTK5UDv2O3Gj1e2kLgSFxGbgij5YNWCS25CJL+qy5tyL9gV2g
hoUFoLsGLCdk7z9JmHMefakBWJInWlV0Uj6XzeP2VuDZlXxTIlXJ5v5O3bdHwT2U
WyVjQfGakudjMcYW2F40bPQrdUB/xYMb+txUTIk29mED6jfyGZDjZQeKOvxKZfbA
qxhUgw8nb4LOdIc9MEMzDQC0vrn4rEdJfBe4qmLPK/LgwXsClh/FVnO6xtXjQuNa
O2ZJiZ9aSdALsb+fXXOFmOzUlh3AXUD31tD1O43PK9GKFOq+Ubkk4ptb2IfFbgqC
6Dv19GIFWQTyrroUZ3DhlgkPO8TuCpa/3ebXH8vQ7fl2Dot3fSaUt7+BdZoYIiL5
V38GVr+A56ijZMH9u/hdF3jeKIqTjHYRhLDLsDDlrhn4tTA/KENZJDev2czJOwJH
28K8Hbe8BBgzeOJAKVIL2oTPbvJTlRSuYMDQWI1/mXUItFCSiFgczivhSWQScyR2
pw3axbpqVuhi3cRF5PEjg3NWaRL/bBoz2uwhq271TeFEo39do8xx/MRBHHLS4fLn
GnpbReTuyOM5a3yTCN+Q46py2D3uwBbZqUsNFaNyvyYbNzkZ2JHhkmNU18TW7mjd
dBkhjgNVZOoY/ZjdWWfzmQcxYELVBcszBmoPbXo1IGSPHFY1H44RoyreCkHX/qcR
9uk6LnfYV4j7spaRpG0QxKiAvGCGlDDVPQ3CQftZxjusRPX6NTsIK9XAVV2DH7AJ
KBkirw+dajyH0476FfhVP/AofUpSggo202Sliu7aL7DWvGxwWjfPDQDYslPMBaLQ
nL/TQkmf0tyiMRcp3x87PG1K/dTP+iRe0DLUAFwc3f4Aw8ULOQk8QlOwlueqzEo2
o/lfYTRKtBeg3GjZiX5MEv4+mwpzigT+ReSrbagkdLn5udIJn6Vdj5SZZ3ZMNbge
TgnnPUxYF9NEOGAvJ2Kii247oioL1S7iH9jfIQMjxIzvuFtWBErxzH88EAAM5bBb
LpZP16UevG/aDV0zdO13NR24AWWVBTV83fXnXL41jTFkJ2CYxvH24sTeLnAYmD6K
ZxiAkC6RGvZKo2RLoVmJ3Qa6qS0kzRW8hM/NhrIE7I/OrqoWlVfLfam+qS1BN4Xl
htAjnEJGRzzZ3raO+xk7IzfEggzsl1cMKNsPywY2/hJq+vjcOCLN7Ntv87wPt5UK
jdFJjAo1U+dgm+zS/l4Aro9ui9mbKgtkmz/9It5TIx22ja64Sab6Khg+s3gFYUjI
5fRMbT8G+rPihC5p4Zm6k1gLZxHR3C/djaChhvu2p+72E+nS1EW0XqdofF13d5Hn
QyQJiLBbJfFzronXJZyjIKTk3iP50X+cMw6WYV/Xvs6rIIFBFXJ5ae4wTJPOk+lI
LUGMSXo/+BYjONTdhKKlOjMWLaO5HGGvaXiVgxKuQNZiGlrHlEIGFETOWMX4whz7
ZkvcFa6breNZjLxNUOnjqZ4wnvqUZOP2JFHQjvftnwjsEr3kQp2t8P8R1Gtqnf+X
ywpiTA8hQTa3GhSyePQcuLB11IVI194cd8CK5ycb5xn0hmj1H5MagyCH6CaQHTmZ
XsA/4xhJvLazmxd8CbMZIElBOy8jwgPkL34IPklIc9bhK8Y32xH24D7r44qQ0qC7
SzHuCK6bW3L2l1v4Ep3tspJqCdWl7GpUoMAJHqqoNbFxc9/7FO1Dhipt/dh7CVfL
AUFJ9HC0GM4JF8Gv3w0Oq4W2MTHrzoQYEKNGfsO4vcDjwW78xqTxsx0h2FELbhkD
Wh+l1X6YsRVLaUob/yHznKiDDGtZgy4QPmg9A3bbu4Dbzq1k8+GIPpdscGsUDzP/
tYh9LJKfuSNZXxtU1aLBgL5UVmWyP+Toho4OanKU/p6sqi6f5QjQ6R54eK3F/7uf
NYJgOY8uuEe5tqbEmFii6lQFjn7t7lC2z8k6oF5HxWgZqhx1mSKd30/9Ywgg/tdc
J/Bf/h4QX5IsVPUa+9QXZobyeTHEFYf7f4cUJO2+2S0wDljjynIOJkJoEjt5Tg5x
TOzLX6W+Qxq1CdGt2bC8bqHLXU1//1T7lUb58N5Q1QJf18N0LnpryhA1fUqkeLxd
/8SPMLZiIMSeN3GrtmwO7pGOQf/wbC+7Z81DD8K/+RtiFjfCCtOjcVutFzRH4VOP
9YxWqopIYpf2F5SPgDzxT6sPn7gkeyvc6jTHD5QCppvC64zwWQ815nM/VnU5pA1c
XfMH/hPI03fpVIJY9ua+v2zdrgIvj8lGFIoK2BBS3RSjisVOFriVigZWN/xlpRvx
7jiKmEgMG6eprm9EX5og3HLFCztSE28txmxBZZ3qaeOkD0Pcx3/lOi3mqSkx2oT5
`protect END_PROTECTED
