`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mDNsDPNhrk6Rf+MbEzRTHZQNfCCcvcPFM7TGpQ22yw7CCRhP8NzlgpvYMSZGUgK/
KIgqbUVECljARZ4j/z/ICoWtjvd+eIs6EW913gLQ5Z4oAtD5XsTtqi3nvr/nLKeX
p3zmCakGU1Ww1GhuSmkYaduDLP0hSLNXaGHCHGfEY956T/5TPfY1cRVK0qnHCZic
FNl/r9M2jCKQ9SpGNOF1qQIvMePEd6BM8VdS+OzihteSvCyur7f5pm2KemjwiFWC
b8eBVDq8uLv+nMG43A4YRpPtpX5jcMUUoTihVOY1nih/o92JSWefkjaEeHAhZfBz
c6K8oAWC4M8d0LxwGmech1/DqfO7xDNV6iBjTeRoBxQ5si29b2SxDMYovFv/ol8J
S3x8ehpWtoHKsHM5nNXhMoBYMLs7/CurbVpHD7qO9dI=
`protect END_PROTECTED
