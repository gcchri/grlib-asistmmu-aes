`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O4kF2kKKBsuyoyP/R7JKigi6OEhKwOWNG8J5JwFAX0HoeSkVqyYdvlS8OkuUUx9b
qTOxXNlI3lfgeyNkFoiyOjttXmeOmVOcBM4NHDHcnWscKqgCPqiLNOwnGA90ucuq
pssNddF4EY0JkkRscDf78Y+n+ZAWSVz4e2uvTMyf+kzya7rNHO6b7i+rMleNn2oo
yTkhu/t5lttqIhbXECzMyCvvTUV3lo/qeyMaxZUohO6Nl6TfM5nmXeebKOLAcLg6
G7exqMqhvOQH9B+fPJl1BGZRND7VBBzz+s1Qs1JoGFhoxncFX0++mELkhdMEZA1T
QBDqpJgj4X8qFmLAH4Ap8WSl5I6nqnNN350uYdAIL4+JIsYHruZns3MfYSobMZEZ
HIBQyCjhhCzb5e8xW+neDSoZLZZxELU2FwgUAxNeNtAfLs1dRV3gr90ahbz1m7qH
N5MBurjFnN2y2RQa+FT4rQqDhCNMp46JCf+1DQ9gwnZhig7cOnyLKVfXF3R361tJ
UYxKhdhVKv4tXEF9lR3XibFHowpVRZDF803oKRVqXoo/p2rOTfHuNipPiR2QKWaY
qEokIalZKzP6rztyFOA2JRKONq0QasDNforp8iwxwxX90mwdXAvaizCgvPE59bDB
mmGkavgMjdTJv4de9FAKLiRjbRgaAjeckl5tFZYglCJ7t2JPGQFT0kHKylAYVGJl
sQ0W1Gb4gQARfz4/I9xY+qwaIYqPCJvq58k8Fj4d5LHFo3VYLmbYynV5IR/UvtUL
rzyDnbwvfksypd1VgmHR8BRMPsuBeONxD4T3AoNTHoXY/wCPrp50mWHWlETJJVPm
yBKAqdPcRyXMCp0P3ZbkOUh7+Kc+k8CGfX9QiMiJ8IMMnVWfMWjbu/SLlb67zXGP
tOzH4AEaKjrJTH7XJnwD5lXyYrgvJIW3jWVnHeR5PgXM2TMarHtrHNAslHHblqcK
KFfrVhuO7o4dXmBEmwzU0c+Mv0qUynlWkn6UBAlJ3IqJi50IIg8wHpeTRxEK72hf
F9WakhRpvzbYTdcQEkTMGh5NJRBKv3Nal52ZtqTBv/bU+PiZU/glKeP4NfSUUNb/
oaJR76ddeMRZ89FHcDMOXr0Ksz2ZUfOwUTgikaP37fa3k9VzH2cEap6j84i+JQIy
c20t+v7f33Y01SGa1r2GJwvFz9PudiXMKL/ciiGoRzaT4QitjhM6jxHnOsBsF2z3
WSIz9zkFfMKfvXTuc6JXCw==
`protect END_PROTECTED
