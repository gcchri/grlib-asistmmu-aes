`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/kMcx5BDxb1iygiia2FcD87YhV7IZeJIdD26VTusSxQ0MNxyRN7FYseScV1WSvc
UauLFco9QIj/DvYRvt58B18cx6f2rtjuGs36W7Mz5vQcmx8S6gLFCHq1WcrjFRGb
hVBH8wrseAxJ+c3F+bKrL2LtmMq1xdNMSatbh1xFwKfmqvBcnC2El5vVM2XOiiF+
3tQhgAPrYOhmzoAAIXGRB8l/fU7DiK8nHjH68CXKGHC7gxHt6NgXrAW2uY0Kpp6Y
NSbRYCIzFtw0cmXD5d5eimBWG0WbiL6y5VTidRcqvAmmwbm+9TLokMgWpA3metRW
3foPIVWqcScG5fSLk5IMCdtZlGAnr5xMih/S1CHu+wcSTvSadpVv3KHb6brMOGpz
l1KGptBV58AHF/3Djs2J61n+5gng93SVaXp718GwrHtF0K7Ny4EWz026Dayeo8Ih
`protect END_PROTECTED
