`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PI6yKj4/v4Tzd+yVcN/NNxOxUWcxu+LrI7clNApQ0tsSnl6eNulnZmf2+6MJpPvH
hw5firKCHrFtaHfyLT0sQFJv7EfbOR1bUk7lZV2INqJKePsmR50tolN65PHn9WNh
2lvEBSsi9yeLrmVVaRFTfPoe6nYtQZPYYh1Z6kxejj/G3o4ouzsxWEzYP9khLF/s
QUwtcD1hAaWIDBi3zzMXQBTSm4sLalkWWMQsZIfZGAct148HKKb9E2XU1KMhCU5P
lrqaFy65SxswzLNnKhL7shGf7S9wVayngHeD610Csv6X233kvPkF79QgKWtmcP3l
2l0ZDb2cUT6vMWyJIWTfZL9zZmEW2m/m8/6GKYENzRk=
`protect END_PROTECTED
