`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWr1lINgsMI67UEmGUyD/91N7H2+jTKDGRyfjI9hJJgK0xS59m6hGqIjJSuEgIdx
QNuTNeUbfWo5jFOmK8ze8EIPsoemLkvPnkn/HMYn8UoqgGxzjXH6R5bsdSMrRxH+
FQ9PRHLKvnO1vMeFFhe7NSpY72Mi6xASaDj4xLixn2GpPNwV+mnORt4/uOu1/Wb6
VtrePEX2AscRU4KZeIlK63cgBHHbk7ebPDynU/zuT3v4uA3D4LAB8TXPRSvF9vpt
tXvgqXf0/Y5nhRDKvX0x4LZPtHmOQ5j7Z5Zm3GVWipu7VuwsRytKYF+5swZSxxa5
viXTA95fblLjwufPIW9XGh5fHW6oi/4E77u6f8kknzFrKVlxqt/wj4id2Y5xDfJ+
FQZgBHH1OD2Fh80e0K0aDBYBknUDeBbKJAG1BU9LFPuAdo6THDqRVuxtKedYmvps
Y4AbUUr776AZyQCW5cG1Bjm/zb4aD72HAkzaFL6Vpyva7NE8DG5QBIIY+INCkbqQ
DcxKb8JMj+RzKa1uukhutQTUNG4+AXIYxc8QV9G6eWcM5udr0LqFPD86hzmH0es5
SL1u/3jnqlU0fNXU/pS8HMnP4oqjI8rvqityuQbnj0fsX3YZ//jnUKRNaPVkdnMj
tvT1t/0rpbLV2HWLm1APthQ0M5CyYaP18yc9kWSGL72KRjDW4v7v2DDjQJ6oB9GN
Yskk927tEit6YmN12Xm/3UGz4SOOSRHL98iSsJS/ZrVYLv5LGqPM2+GYmkjowrv8
59lcSlaHiqjS8DfqhFmjuIgEilA1KWaniPvTpSPeT/FBKWusuTxGSGSCeAy1h152
p1S1lsOOrcJ9n9BFeCBCm7Msr2eCL/aCcc9AAk9uRi07iwXyvDv2LRW6jZ0/80zr
SG2/Hwv829HVRM/vBQWeQrmDm7agoHbpHnvY1sdOm5qwXlviEpZzfZoat+dWfp+a
VQHmIYzffN3M6jZyl9XMf9vih9HCtvvwn8kaJIXmweGNaoLgIUG54rK6SZ3M7/aS
O9z87cbnPkd6FMEtE3pmZp9wNQ9hsC/Sq3J3bwvQFK9A+q/a3qwhsPOoRgRPT2g2
el6QkCsmxvoxVlrMHxFgD1OOg8yE7q3vpajK7CZ7Tpsepd/lQEeMwxq2CYxkGBXi
G/MDkwSN5XZEzqO6Bi0Yu/8x1QiDDPYO8ZLNOlQyYb8qm3ouydHPGVloORvXz+Cr
VrfajJp6OnEexrop5I63MtaWL64Wtk3rYcRNNTDocxPJuOKxiMm8cQ9Nhp6yzr4c
`protect END_PROTECTED
