`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ghWxeAXGAGCmWCdIVfjbL+W7WfZtfQUDhv5b++roi6THFWplW9pQKz8LYoFYZKE
NidzHif9TpFkxPEGAGMstyVgrx45il98MEmVBlrnEDBVpQZn99sfeTNGzqAI3dEo
KI286/JlPknrvDzRzo53z9lyxaxdoM3bv1Qotu64tDeKksg6CHa0doMpOPN26Sko
zTb7HhLkfTBU6EagwgLi3Rq361P0YVExSw3b7PRb6UK0fRtxbW8pHcwKVmZOitFJ
lGUHcK5C9gdCAH1q0JOhzrgGk2FHSDKWw/UH5DqqGcr+nkgwSfvkXHbkhIvOlA6r
K1tGN6dgRZKjq53z/I+YhYM4k054SZGUqAd2AkRb9AxpR2nkSb6Xms+6Qv3Goxl6
`protect END_PROTECTED
