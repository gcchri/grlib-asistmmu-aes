`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLl5qNMm+vQf7IhY8O6yjrw5qIxEIhGFRG8uknRcBQmdEzFQRwB+1r1pd0teqRws
OK5epaOc2744bHQzq6ZMaVKnk5wRW2LqGui9vc68eDXIp/XjzsS5aGpmMaImLvWt
SLjXrDFEIWJYfvzsDnAlMZ10QNobBR9hL1olj8zDIG56GUPtuwE+1RUgKDDzK0sc
7XtYdHqoTnb8NSJQvpQVkmmZ108q9WgC8ZnqTLIsT3NB/o/K82TmuMae0sgGc8n0
B10pMlXEDuIAvegxZWtFEi/yNYbSglhrQK2hRbqao5cFyMiom89E0TDH4Ai06DGW
IrvqNq1b7ZHbpeJaveNCyMDfT+baveizbosdA7zAE2N0+OtL3P/62pFRAsvhohMX
ChrScQPRlXLep+VZh1F9y8Vy8XZ21jQr1dJlcv+Y96yNmkvTQ7f7DaDDv2/dDAAc
G/0OWokUwwojv9FRvCVisnfVAjvqVtuG2WYLPlxZPBXtZyow6ahZSxtuBjywvBZQ
7HZIlnKX12hOpbNbF1NbCZzlOpXubvd/BAkTG7FXM/CaELgdcMt+FuEM7E2MqTk2
oG3OTB0r7Mh0j3B0D4fD4AUNO8FQVg1vh/275oZFpwBUJ1mqONca4pGTuwSzIbxU
s2VDiQpGThctETj2rMp2sk8wULBddDYxEvyMwCNTMWbi/+lK93yF/6xJw2GNTvi4
MXYtXaaGc3Xh1/Q9ncWVFBeziM88H7DzdFfLXRFFxN0eeuIUKE3oFKone9Sow98m
nAYfVL/z0OqZuXmB6Yih2fe5Iisf4W7SmYwHzcGjPmjdrb+vbJ6AmAA9te9H5e/s
Lae3/fszRtlJkZzOT7/U7A==
`protect END_PROTECTED
