`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PThKUJL4E1nfQsp29iq9Sxhm7QSj/w3Fsb1kOH05QH3AGNCVFrICzNQ0Ls/jN1Tt
gJGbS1rhGvur6N+p/VLVdoEkNL7GEUartn37jUerBc1fapkUIi3arrauUkgVpm2A
vP2GUrl7QxNq1DKybGINcilTC7FMe/28rzmCgJDLv3rrZ+XzMR9hlB84QXXISDxp
xOS5+DRwUEATr/sWe4Gh02zmdzpz2pPhz9EWaleDBBSJ7fxT172Gkpt6/J1DhdPv
/q2IjtEPimXpQ7zdNVyGFtro7Ie3N2jTYc1O5cBTIBUGLdtELlnLKI2PelNlVDyv
9dU7qtXoeXHPdtYh1Zz4xeHkWHD77/7F4IZkwXJCRX+kIrPv8RNhohr6yzWvb7mT
uKyfJC84oF7jhcXLgRYhqQ==
`protect END_PROTECTED
