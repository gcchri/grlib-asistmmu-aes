`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wbmULX5r5g0FReEFxLX/A/CqPkmslo8Rx5NiowXAjWS2jLEpxRU9FcMQ3LqJyGS
qHQwOFM2KKY9jEZq75oNQylhhkcYtpq7fov17B4DGNjHzQD+HdrRKJcpzvm4A6GW
u9Lpn55iZgOHrr26nhkUp6qqwoWntuE+Xb+yXhejpAVzqvJtu5WcL1TAnKB9dkYe
qPbJzyjxGDnpQZGsgp93xOvCQnpOA0SyubZ945Ory3FIYqsXUPwK6M3oko+aoZHG
sFEPCX5l0Z12xASPgIiYnpcgbrRnoftmUBGm+/X1IrlRz55IMmM1x9U/RybRQWfJ
wpGRRnpee4faXwO+ooXf05ediJr5J5EEauJCqn1x2Ti+jf842KzAnDo3OjD4t16B
PbhII6q1alwax9FALIpL7lJa+VtF6GOjoCpg40qwdR+v/CJpgEt+wxq3c0kLY6ip
LuDN8nHYTyZJcT0p192xcw==
`protect END_PROTECTED
