`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWIrH4G84BqmfpNS86gKqeZPxbP1ubI5UvdWuJAOF9t7I0O3nQifDGreYwxbOHFq
u8oM7Mt7DnrV+17BC/FLvxeStuhXTjs+PBHKqLMcJLmZQYxtTjhYpMCzmij6CgbZ
+xrwQV7C/owHACPitNgAZ5KrGLhZ+J5Fc6CATpHVi5nilG5J/WldYvh6DTHP/uBb
GFP5SsqBuThGV7Uqol/2Su9+HFOtHwHutnaGmVx7JscNvQOtiGdIjXhAvloTi+nP
0hp74lmge4nokmXOKdDUs/eS2lMcGeJAd3wBizBDMzfC1Fsv0uaDBbngpCHLlVca
EPBGzc5V6K8IJmGzH7QK6ADLzLCKBZoSLHTgxp/jnK/Y0nk+h0uEEJxuYX7wuIgB
Rxts+5auQgbzC/qqPmLnrW37kTnny6MOog1dM0ovLnaLk7nMfg758BsDW77Bxkmh
lINmSTw9eUUXldp5vJ5dT+2/PRppY9ys8Mso0w+MmiVMiv4c/6FRZ9gPPcOjKlcC
5O2UqPGxZ0smoxZ5fHNIdYsPAH0CFWJMyGEcFtYI+/AafMhuGLzFYU8n/ahOjy4f
VMCwf83R9PTaNZATwpmXWK9K1EiebKGYYVq9ekqe2V8HbKUt70ZKldEk4UM8GFDd
3w3GHKEmUtqYVHH56tu0D+o4DHbSy/LS4XqFSNOUKwuL278N1UQwaJYNmXPEtWsg
pkrPwVGG8hliUHCc6NTzWrTqETGlHYGzMvMCCpjjiG6Jje6lUma18spqo0GFThx8
ei4GJSHI5/8aLykOPTIu7hvlw3v9eD0Ef2/9Ubt6PjtFyp/DFQIabqE372g3uilK
ZlgX0xlgC1WfpMow/0z88aOopsLL88toTEQSsFXKizxwAI3QoYPRMb2QGiDUd8Bh
TigC36A1Udt58R2yMZCGXu4vpKijWQHfyUCM7xpRi+k+PeaaS+ETEESlRlnvpXS/
N8+qaa/yLNagR3Srng7HvezplfO4yYYw6w6AQMmdgglavU4iFE6uc35exW7aOxjY
MjyT21rUlhFDDB8VNFmsFonQHaVHGZwN606oUfunvz07cFzmMFHzYvzj2tG0FWve
r2dgIxDVG4JzdPb8T7fU+GZpnrkgbUwn5AsvcFE54uRqX+JqmJBluSAe85BpEYS/
`protect END_PROTECTED
