`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
as8X5RkU00hEvcc51vASBDb/bEqf+V84v8E3sjPupzwtWih/ABAAGs4fD10EFyKT
3S594AZ8ceYGm2KvR4UNK4VEfswoUoamBy7v6klzy0JbEIqHSBhQdAEh1OdfcTv/
iBHy1w58cTxzVi3WedcO3NAXhZHm7dWqhCW653XtH+YwqisruHeYH9uLyVjkVYXy
vJUEnkcpifiAIZ6fCrrmc90yMOYFnLpBPZ8xOLoXELgbzScz8UFR+UjwKlrsDRxw
iuRw8Zxp1ooF5QkjvHtDL8PIjvoY0HkdMfFtDyaQofE2Fa/4wuqjWeWmvdfrHOl3
MblDmY2xzTNr/WllUJWL6HYOoulgXv2B5bQlaKDvaW60FkTAjLhJYT4szY8fiqhL
bsG1+2dfv5pTTaIybvMngs4vS5024oIYbYE/3RSOS83Q434umKFxK8VFZZ6P7Vxo
XabfKhBriRCdjrtlQwaif4woVlGuyV+OtVWf0diSXDEaQVgXdBe3ugbyh9D5a4ZJ
BtF7o3V5J1tJ2vkk1P1rwJvUeeLzR1+fmrPqOw8eAF2/1v+T0lDLU0CseGnw3YWg
RAAxIw9R5X17Jj0MQpCaP/o2Xh0FEOQCr86Ie+tOFjrBcWTQWmUSrinrDZpG1fgN
8N5BZfbZZKTjE0Fd2Vy1DY+F5EhgVpt8nuCL9+UTs+VH3hRPipnHJ3lITpDZVW+P
VKzBRikPfCZEwIuFfSxWQvw7SAfKrK9kXzSgUrvnpmBg4kpQgwDxanwJTHQaG7Ky
6+NbSW0vnlnEBqqCgvrPAkBV6obD2nHfasNcZNI64VCAQ4xpeAsO9AYvJ6KASm2k
wihdJWul+MqExCFILQVYC6ykqnLP0jt9C1kUAUDGwkdaBOjkyI8y7X2qiHCDNvXz
2TTM1GlAjroRycIRPdfM7bTwH4F+ajs2Jd3Gg8YBYYkws97wtk0KEyAhQRKLg/4w
ZdUiuQX8NMVWQfwP0N0DGCEzKFa+0PCdc2h2ftG/lzk6bFcIQDEMNwCUoStF1vSN
kyRWhWCkxWr27jOCGMAw9b7mhDVp9WDowxjSykhqXhwat2lanX2oGTnA/hg3iokE
zHURoXvu7suAtAPqiDCydfa7V1gUl35gGiTiYkLQ1PQLv499ttNMHv2x7Zf8Hl1u
owUanceTRxVMrJj8QJFXss1ZJqwbIxv8V6QdFAwYIcsJYKZwQj9BoaTROqpMi4tp
qOEREH05k39eV4lJYWUP4cAiRJuXFwHHUK682xgu1LGljsZ8iIvtDBaR3tWmDGFB
LQ4xxkYX7+Zht4XnMnC9g5B0qsEmEHSXrFBjdtDqdgfaQOvUvelhCk07lG5U/znX
rMgDu0gjIlHuDp49tuPzF1jH8Fcp7nDIJVF7S4Wb5KBRlG5wWRSOY3jVPuxbuaXQ
`protect END_PROTECTED
