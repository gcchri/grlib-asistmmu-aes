`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xSZT5XpKy44zT84ueCZUIpljeKo9Wd3OFfOmK6aN5MEjK8oJ9pt4sig+Evs302Is
enLIffl3+/aBwq2ve75rtQjrk8kSxFVBUalg7DPeDOEtZo9zN5ljBUzKfZeD2eEH
PzpU8SP0XzvCTYVl5GHoAhlVf9CIMHtZiz7V6RFZVPGM+GkCyeme0LjWL18z7RPn
KoKWAtcFO91oB2flAJ0cayX01Un3fhiy78bFEWSP2WKHQ0zBndSBkEOC5dzOPY7Y
Zh9B2yKaFgkBiUnKMO3XhG/cUH4CeAVBx1aoPXFncNcBHD/NjFxf3uOIEulkFGF3
wunVgex/Tncng4sA917XNyvmdJLEWD49+cgQNPGQZXsXPee3Df/2UtgFOfhqFDhp
FPrUlSBxHfoCmVs4E7AkjPeK+ZG0w3NxjIXg0O+Nkt0lgW6j4x3bjANwjpnsLa7x
xZvoRGASLFCrHdcTYixUqf/qE+j72cgEJQindA91nsmjXNgDuOphvpADh4rBIT7O
jOp4tw93iD+twrfeZB8ek0ZO0O9+ARq5Bhp2zc/vH8Y9m372l/AMn4FWiHiiymVm
02gY3oMd1QJhLMrZMmsbX9+6fanHkrAjwFKWU4nKusixYLw6VAtPfJb2kMmlem/U
S7BuPSVf0wNvkWJA1bDVkvj/LtmytvsKczdAcOCZHg9m5QouxcychDqUTQBZV4tM
Fv0hN5fnoIdpen4AO2vh2DPFOyXk3KqBvs56UPVPeLMz52GrKlQA62NPYhU/1x8o
wwyv8r7W7hvEk+V91muUaw==
`protect END_PROTECTED
