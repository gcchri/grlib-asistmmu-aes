`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2EXdD+uBmB4GqgipdPbQ1mJQOjiUxf5UMywI74IukDFbMLS/w/WOpRlOiAqa0tq
c++Guh1I+IxvwAgwLp3oWszsrPlvG3Z07zF4Kn0WMcz3lZsc7ZSVTr0FszEV1SPu
D+HJJbZ9acqI/pFD6FokcynpxwB5NMu8IKRAnXGHiuaZu5VoBaP9eZ8vVgbAHKpT
g+UpAVkB1qmNHcr8FMnfIsK2h1I5q3dwdLoFvNI9tq76M7IGQ303RQZxG5DwTSoD
A3ato3/pWmlwUPvSPNPinXluwiakYtu0DkIu5NnBsfEGtZErqc4A6lEHNQFGpG+r
fGyD8QKOouWNZQfKJuOU2ZGo+kPZslrrJdPEipvV35IZuWZhen9OdnlspqlWgMjB
vsq+HDSPEzEmuT02ZnmX6g==
`protect END_PROTECTED
