`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kRAQ/UEw1B40+9C7WFUdpEBlrrL7NzUu+/BS3tJZoeWXJ1ZuknAPj/iY8bE39OEr
d0mdrvm9C8mxy4mB/AIKQP6LOAFIjWqR1DQbGDTf5gceItlBFjoG0fvJufzLGFI0
6jffcMMRr2yNkv1Ls6W99De6jd0cORALXPhKavhknzW4+OCYQ3qy65rP88K0Cs3X
Tt/iGyepzoSeFG5iwOouTPwAUGCB48YnkUjhCmixLptvKszY1nENNVZtCBzpm/Ag
SN3Eav7qP555t6/A9KqvAG4obC4O/p4WHTWimiuEUmOJ9Nlp70RBgkzJLcm90SDF
1qvgvcQ+9yLiD2/6JWR6M9EPBhtb+0fF2b3a33Is+08oa+Dcm48DqBvLf1QU5q80
`protect END_PROTECTED
