`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rw/AmeSQLdhTTboLsBTWuMmyMPEtSl/Y/39hrdYj2AxvcS6mw1XsJMmxeQUxHzfO
TwIrUu5F+DdjAqaZ4el0Xjye45dPpdKJgxj557S0lT9WP9IsIV6ZDGcql64FGoj+
bys0iXnJmZ8uxZu1HORvuTMIzuRKnJ8KhUspRSrjz2mRTpODiJCm2HqKbLyFbVzi
h6XRHE34DgoS+CBKOieJrkx56/ZjeJ8yJqMvPx1Ppg9/jWyfMRPfafXSvlfWw2HM
xcURT+bhSWGYkUWRPX0lJrcys9oDsF5piWSaxFHboz0XGNVQ94sNc7UYIKz7GxUl
raSBzZPwbe6F9pYAf05peE6VjtJ5iiQ+HmHT+mpl8qY7dYrV9jc6gJfJOIgcMx0w
jM3lYRtCy9ObAUAMtz87oo81D57lgwwk++D6OpTF+45SMbOYdTGctJ+/hQyCbaiY
Yzgv0ueTheWTWsq0snFyt68Z0J9za7bqwNVyMkSvcOSXCp5VP3leU5IXVT/fUEHA
`protect END_PROTECTED
