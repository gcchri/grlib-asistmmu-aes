`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YIEFbOR+C40TKCRGf5fe9DEHE6YMMSnUmfBifpjgl3JT3/Ocaw2m8R0OODnv0k0j
edsk4hL1OFoSMS2ESP26DmTmr/M2nNgs+KFP4WjAQgGmooyYruEZYV8b1i2PtZT0
+YNj5LEgZopHdtftcVumxaDhp3pV7lFvJy/VlDUVUi/t/TQwgRVIkiHoLnWAUwaR
oWyMgwteyB3WqmaI6VxcafyW2Y9lLBK6vEXhSEkyASEvc4j35i4PLXykQU1Q4s/a
uKlSGOyuC3ahOUuCXw5YRPNc2Xf/k1Xq6dDJ+ldyNf08ZOuUNpFZ9RwQsz8/WLEV
IX4gIXPAcyZ4g2IM+uM8taoTVxfKS6z1ed3zmg03iBYTYmv4bGXiC8Qh4zN/GdTX
82A3IF8qK+9mJO7vOlts9icaDOvaYhfhytRe0hsfw7GtG3gsBODLNbu/TVqAhuLu
ggXum3NAY+nZW3kFgsqu/Dpa7M3QFwUivaHp3KMeS2dmdZSs9DwhoJve1BMBxIDq
6+di0jTTp20Yy+5HZWdGhg==
`protect END_PROTECTED
