`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EE8NFNwIGty7rx+rPHeRqqkHkMOJe9Qn6hIs3xxSGZfS4HDfmdqB7AS20zGHjub1
4FLsPJstEgHcMsU4rYLFJ0hWIBGKn39sNNuF+j4LgdHOXiqkyFxXTyBDpVZpgCHp
HeAEjdJRHqLDPid/f2Rj919vVGJsACzKHey8Lf2B3vafGAyfSti1YGNnlOVTMM1C
c1jaaj16Bn7DmPrVjz/wVdCmM68aFm45+vxDXgMIFGsF8J145P7A3FLJ+J3XcQKb
KasazbyfMy2kxyg9JTEdC+MXtJHykWxDSE/6EBw7nrdUANElrXssSpb4o31sXc5k
RI7oUazbwb7F3L88uMoBXNREjd0hEXH3izTWIQNvDh28giB3yQqlup+IofEumwFC
KFkmQasoDm4XGeNu/67TtYuSH/V/K033sD113MBpCjWnXEEW7gVH5zL6YRiPdMln
pU0g/EmXJW7mS9Dx17bZGnSV392VAMScm2QXFg+5LnyAfUQeGETGMYhB08KSET79
auNvcMlEwDrQ7fEsAieBtTIWym6ntK4KiV9PTz+WGPMtDbR3q8YiCSB441Ve/L/m
EL08LCVRaVtUqA5Pw6fWu9CIhpOk6qF1g5z0UvIFwBHYcmCd9idjy1nrGSCoa/lb
CljzWZlkMPGYroaBeY8uJY30UAMLNurZGpz2tKL0xaZ47nvtQ66feZpEySomgdGe
R1vKHYHl42RlANjRJ0Rz2XtnU8k3rI3FVH5iqvVBMdK+2m+KYUEhMJR6brrq5x3P
YbN5hFWhC0iCOqxnTLt+My2BzwXHok9K3ueDl/iCvYkhY7MMDU1UBMBKlV6o1n1T
svsoFppNUejaJqJHX7XE8d7JE0R8ZVuUGklHBEbqWBLegNumm/3clouTkr13xesl
++ixSx/xJil8SIebfqeYV+utFrusEhsZyZB2BXuvNFw7yIsoENgIFmsr9/GoGsBh
zi8UNsucJw8AC6c0KzAWH/WzDBaywxpgXSx3NRryHdi/zpeVWZDTLP8HkzwiIjbY
NCr1WfzTf5Fhc3ocFhikO4BcVDJFs+JNL0+djd0QtbkBFMSCdYKTHjpFIKN9ctiy
NK1f2Z3UimC81CKs1fqkqAnR4NT87SGJFAAAnT1izUU216Gy/Dm/Vx8uUbv/mHfI
aFMKck/wLXF3So7y7sc7qWi74/Bmei1+Qtf3DOdSy9w+CUXSupkmgnvyUYwSX/sv
Wh2vAjc3NfrI5zRHl2sXgjkd8sW1aZqsVvX0lw/TLfNorBDyknQ7abwn7mr+Nkx6
1o6qeNv9eFGkoAoGPcxZ+r7SMsKOs1Oj0hO16SK/e57LgeDC3tvIuZ0gRo8FpwEY
/duZ7LCOgqlkE2JagIFVX1w/hesNgtmn1MCBs3qFXaRfA6oX66BifvZQD80hwKLG
KFVBHc+U9amzO/qaSpDHEPpvaJI6hlEITlMNO1anMqF2/U3FQXQgdw8dhoI5kT4E
VTCQGr8/EMnWNlXEYD4JnTF1o3AkzNueRgyEaeo0kxZkASFFXBAjcYJ3QOpWrIbD
avu0vGQ/0YNrPo3o7uOdVQ1ugvh0dCOJ2rDYFSqa+eeS51oN+b5ZqN7BptaYGYug
puDlFt7d/EaqbHAxtWbY35nlDfo0KwhWrPhYz96L8ABDgdvGepFihlIaQ2sl8NoM
rOUpuzdTudOOq/KWvkM6/eq3bG3kygdnYIvDe3Uz3HJ8/fZb68RrC/hPZAV5AWaV
h+FcEClCVYstNkO5kI5T9hMdEgjp098Hw/IqyxpSRL85t3wgmsq6/ibKPuzMFZST
8A0Kv3Bdj4qWKxglU4xE0aR3vn20kPHhsde3VqraJY1vkxUPV6bXF7Og9iYJAREz
/dmQpYE/XJWoMk8IOQoEfMd9CWXvQ0LUqKfOWUc7eBeP0YU06rYhl+4+kh/cX6n0
CJ+oCe9gCoHLIbUg8DH2R2SY/vxpCyOWtS8xV4A+ATVpJ2hkPs28bJEiOHuv2Cva
h98Il1rGnmj5Og2l/Fn0JEVvrvfml7DGDwv8DygbGFtBS5ebI5I4vBTkLgVJ16Fl
oXLgGjKYw3/1LVhakthlK4OxYObosze/9arUqtshlVs6Fi1zgkMMTo9XP013NBCx
AHqjYE4CDFrvWHTZadwCiLFAckldgrl4QuR62YeBWWyit2OsYzDdn0uCJNrecbL8
+ASxbGnzMJ4bdeHGez9W3ka6Y8jEu7b4+Ck3XXh3Y+UWo96Hwsllrz9tH6Bl50PV
zId02qiv6ghOid1sdopGTY1Bc0ENyS8kXV6jkP4BTTEnxi62IijnnLdJsRTViqXP
lwWGL/9kFuvyXJK/0jNRHY/XLY7HXgu7mQ71ucvUI7B9OsP1yFA1r+D6LU54hp/V
0HdxG3rH6Z2Ja6jjU27S7RyKrrrWRD4Hf6eHkCfMCazr0+jD5pGhPrTQPgxQBA1H
`protect END_PROTECTED
