`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTBwkz1ci/oa3UzfPAtW/65kWi8CWHOSSR9WrelV8i7PgCcFI+qz+yS42QE+8IyA
qj9v/tJktKT8w+EBDBuIFqaovHmI1UvTgArWQUfaAco6YksAbq/5h/7HzZiNABnC
DrvSnWRW7uNdTqky7eNN2nq1L39aAjL0ecIi77KcMM7m0/PmYYbE13u+uDWvYuVW
H4UE+VbZuk8y+21AQctaLn4wmYNjSbRzFAHlEKl+ew+apJFwwvyNRxITy8qkEL+V
xluyT7k8LBEgd3sbkQkFLQSrZL7OoFUt8PNyrMAF4xDQjW9KaBsKBSsZI0ihOf4T
tgCpHJ2RwFGejkFXh/3uPsYvXy1cuD/nT0/Sgoq+kCHZmODa06CmAuctIm+tkv46
5ZhEFAIX0haxnO83RndUiPgw4Vx0m2ZYWdpqAO8FCyvKNw9bbQ7zWM1C2es40m/y
1zoOBx1HuI/JN7U24K/IxFroVPxmYRuUnPKJJc/ftRY=
`protect END_PROTECTED
