`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZacOP/YRX+O80/3dha4QHGsZYNDyredBBSib9zPZVwy+1rmzw/MDnKtWl+9iCFBc
+wrt17fFD35ApVmWWODtcRtN2+d5ShfTlG+JlnWtFvKdR/0vR/+qHc3BRU48DAop
T8s3lC5w2FWSs3HT5g7LthGL9rZBIC63UrR1N7srAX9Ij9tgZnIPeRkam8wEq+w3
quD450aXmTPh6Yj3ouywKlhTzq1hQqHRlcXSboQXsCl8tLkCPxT1eij1/ztnRgt2
I4IA42sYhwOepzMLSzFsgEBmBaQBw8e84zlzHs0I+Ec=
`protect END_PROTECTED
