`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CUyU6xIYpdeDWJ3ies5znD/mYhRz90hK97VCtU93Gz36t8oEA4sd8KE5WSn8jzxd
rjfn3n6H/rYWmE0zCmnnQXT+1Ls28bYtBTbyS949tJ2Qs6hWXI0kJK3ikY0rvVEW
o6etqct9RPsNw4KjRnhZgUVWrpvLoxYYMGGuiA3ziXb5z5fJ7cgM2hRjKgNJURYi
i0oHmZZz4I7GjLiXFO39SeZYc4WFg3hZS9vMwkI/uu+rDtQsAkqBz7IFCoyViLDH
r3NEzVYGNkQpNJQ3Aqb0RAMVQn17dPuaFSqJvtrr2GWz9riv0uRfuVnIHXEFkCPs
oFxCJuPKpDabDUj1WL8Va1s7EvAfqEhm9KoPRX6gQnf2fTJaGHt5tJ0Q2sSkVBG1
04atelB/7RtlobWvAh8+QQ6kK3Yfoqxc/KnmXDD+wp8A/swkPmfHnjJWCgnjiBW4
rufzmBI9lQyTcApI/S9DdtBvVAyXdKtICersSmjLPMrxaOmqPMkew0s3rcgKh8q0
V4lJrynoOnIvMRAbQgt601Fxn5rtR3MIHDmxrJ+xwtBGmoJ9hM2er+1tN37vroGa
JB4dYnCk+hKW04WmLqTgmUErmdb98Era9iBkQONRMIayvBKIkw3tWuJX3Xqp21aR
9QH2ZdvMb6gPJcR3GLObIMRg23jXQHz+8MLE9mnLTMLx5IdgG6bxs+WCrPYDY2yf
`protect END_PROTECTED
