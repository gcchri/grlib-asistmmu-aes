`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLVISgtqI1aqPjDZ4EtacjVPDvES9UpO5KA3vZhLcyx4HhStvNAMf683nmQ80nUt
FSC97klSxI3jrDQ2lAKt6h2fx3QTpbV1v7vviPp7vVkN0RcR8BADEMT/jBl88zYp
xbnD9KRDNvXJ4s7MYUAQvzeEDw/1ms12eljSdoRAZ4pus3ImBAMQ06XzC1pcmmkI
wziziRsWsfgybFCFH16BNpCkrFwuzOZuhf2shutEaUGr4VzfCn4Z/ite8ICRIv3J
iIdXYHYWXf39qV/jwF4YKBGao9f84qzBoq81CA66wi/UlWZjQJ1VijVmCNXwaBUU
4vUqxE1BaAb2mD3TB1yJZ8X0gP4u1RJHh2DuXjja27nd1baNsddfjIPRhtkxdpGP
PBPcYhKnKDq5EFjatMREwuWE3iRPWBnsxB4itT+SEUqxv84Rb3Ru/RQUD2xdjhPn
uZdgEoQ8bNsUfFJX9MSkfWTgjAGIbGy7EjiF9Up70996QZxia32ub8BefSXB+zlH
`protect END_PROTECTED
