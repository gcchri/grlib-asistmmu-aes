`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HDjfsSa4U+fMaMU+eT8VDM0IsYv4KmO33Jda7B+2cT5jbpd8rFASiFpYKGLCBZ+Y
eEz3NcEWkZU/7iAeZHx4KxBpqIvgq9JCC4VsGOpcEGWMCCs3NBX9j5ir2GxDmSTP
KbrfeOY3YCYr44FrhREkGQzbq2fWe5eWiM2WY4M7Fo4jrSlAwhPwqp8X+N+aYIfw
cZrj97/QvsgWMXK5Te7UZBmsfhRkY7beytyspeD29IttuPBM8B4umHS8KZtyMOZO
TDF6k+PzP+3pXw9AU1OI0fD+ewBSfHeQIJv/juPBlZAOMjS4ehOVwUPVhUsoR18F
unpGUbPNvWWJgLAwa3RbU+JdfM94aCaE0x2TCKLkOkJowKnV21/oyTnuEXIetPb8
Dy8b7RrovVthBs0nwzvN3oVX6Yzi+sD5bMBZ3IvSodAcUiXpk9ajt3W+AgrWxA6c
/Rlr2OTYh93h7ksfK4xkjKmPndG8wkzjTXsQOYXhjhoxrAz4dMEeSdwb70BNa278
WG1LbgVe6d0zygT7BZJYhoXl1v2q36yXhjiah+qvt4ITTBRYJ4TWooW1JxKM85nQ
4sdG2GfoDdvCK516fvOcTsT7DhY+WRb27UKqOhNlpqM=
`protect END_PROTECTED
