`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0n8QWX8lzySv6jUqbQtPF5NzioQ3EoqlRHwGx57lW4XteaoLkMV9WBhQLdtw2WYK
BnUU3kiVnWZhfglqxvlHXy8Xyu8aKlqZX6dyoCyQqJuxO1dxUlDSoBCM1Siisc/e
kgXHfrlchdD2a/ZMd36AAinraXq3s6YxvKkuIuCJRNLq3ZxV4IWZr9VVzmGQleeO
FbdIqxeM7aqat8Z2t/fzzln3XbmvWsf0euloXOE7raD7/AqpvxG0ExoYgTi+5INh
jhTCIBg3k0ZTZ6t6chmxMn+uA0EqZKHAh0ZYM0Y+xDEH3O/+OqiOKkNDjKrNX5pw
zdcvLg3MB90+BMxn+H3yAZJTeKuMXe45FncwreLtUjzQTH1NDfwQqnO1RC6mGMkk
BuXVSSdqWtitgCE3A5SROOf9zFBjKxRQhEXTE5Sr6yZXk9kr6O4kTg+rTWS+5RXw
PcX0AX5SIyHyuCxHunJ4dh4TEXcdAMwTKaxN9bxT8Mh4Pge0sOFKPYgPlKufN71A
qHjQsyrZWfd+B3pcxw/H2A==
`protect END_PROTECTED
