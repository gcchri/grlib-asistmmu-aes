`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6ylasaEMJCOh9P3r3aLfi8f0r3IQy7g6fXpRR518jRoEjG2Vkj2d/RC13AuAObJ
y05hgGaX8PxUx3BvLw2AsguRlFigN9CJm5tr7fecnHVHQcJKCvaahwVF9fGnBQs0
0xSSaNIYivKjDr3oW5b62OvEc1zAFZV4Z0IhYYEfgYhUsLxZ57cdHgxjdHm0BH0R
HfxyfL2DKD1v4JZVsBcGJwwA1mpOKtzddzCczArn4IcxoHUXQLQLMAWm7JFuucsF
g2F+m6+tl6Pc5mQKGS3T5Xq9+BzKbnJiN1VL99QbB6oxsugbt7Ucq1cn1ifTD5x8
`protect END_PROTECTED
