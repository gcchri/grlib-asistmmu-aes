`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjzIJxq8W9MQ3xYuEvY5wV/gtT/U7fyob5sFl7OxrNGYCmx9mJQXkVS4YlJXoD9r
uKsaJHDAHyGkuAUrkUuPRJMhhCC8sfHZiZxGAgIBl0ls7ssFK0a91T7+InjywZdc
Ge6ZhqeasAqjpG1ALzj3EFxPd7G1sOr2VOTubeUOhkeChWhONLABzKKSRJzFJuJ1
1cJXICzn6At2Vrt+5ECFezxAkxXgHX+cyPfyFN1eNnav/PsnkgHi3prIvF3aPCUD
oQLnyxzfCBeiB+Ugg1fuDN46z1OF4GqSscr559ZQw4yBonBaL7ttrB6TQpRrCKv2
d5V8IYEWzU3JUYUw12koT7qy/9YlmuobWug8QHbPDBuj1QKnqXAUK5Ekbx1XyU08
Kc6NaBNLLKmF5gNaTXOYlQ==
`protect END_PROTECTED
