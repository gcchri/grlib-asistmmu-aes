`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Va1ICBu0vU+zIDQ0e2GS+1iTX+6dmNI6DMIxBgIlb4K/o0QFaY1r3Vs7+bx+SFXP
L64pucebfymmaewEJVc+yq2xp8i3O+Bq1whE2PRlATWXYWguiYF6fVC3yt4Gw5GP
4DFam70s+5IPrKoLtTYxHQaPFLkE1N3kV4S/jmoKjHDsuKeEk8aAEHh/bXXli+vi
S4EdQE1RivD6SxbwFMct6uG9Se5+4w5WxztEdfKVPHzmK9DVnabjtnljz/lk8bgu
R1zZV6X6PmvzURYRhb5e24hqJAah9mLVK+k50sKF5XY=
`protect END_PROTECTED
