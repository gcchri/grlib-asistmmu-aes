`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JmMGPwwFDbkwNqrXBrO0O/DE17ClZ7DGxmkWl3fjWYIpZYRST+pqMvIb39UD8tDm
5SNlzk3fin4appDHkYWEa4LCJnDnPROosZFnHrPYqVXLgIcOBDqhfzOR9gOVOmO1
U+NfzzX83CBccL8N7u1kZ7j25IPgh1RcNXeUd7Mi/R42evgendD3e2C+9CeVAewV
CpcxPPSfpZOSuyDhSZ+1QDra3KjOIOlZ1TNDPZ1/gYPMGwZ5m+E3BkoRH3lIkeny
GE4DxkDIKzh6z60AK+r0B1f/C3hM6btQANnUj2yMjFBDBRj6OZKGrU+mkrO27VTo
o72VlHLl+Y3pNwdVlPVj6XAzKLAP4QLfWEIuGuYm2NXPrnbA8kJLk2bnoLZaAymF
tc8bu0xoHaPgHAUkpKhPE0MBAHvHhgUCtBi3xe9vjKxI4cdIRJD19tR2jYpmtyFd
xNERWyX4rVlim3z6Y0Sf++FsdbAHhdyJQQ/hnvrGt7g9M3+8kRkh6iWWPtSRZukh
`protect END_PROTECTED
