`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2WhG9AJ+Ynwe2QmE4LWfjt0DnoFLKtwtDoIJr9ZQ6Af4yPrcaDPVbzjj0E84Ltj
JqmEZ1EmPJ9YA5yc1wdKnSK5EfsaufYV0rbLnK+ApPKaTw94zH0021O2O+5jCAHW
l7oyikkehdUYal0tJl3JXgxoisByYS9XRMCxfA0Wy9yso5xCc2qM4UEJ0US0dCV+
9+7bqJIn11Hp93D2woIcsph4J9UKevhhWURPkwEglU5QBswzgqfUDdhRTxqVBjZH
Sci2qXtaE7aUsZt3gzOdrl5rFmisguoB1ACNnAnl5wisVODHPtYcBeBIfvCmMXS+
l3XfpyJboigDaVi0i+yB8xhdYP3uw+4XoGleryytFaYN75vjmBUXmt1lTL5ma3gF
9aFj33481s8wB3XfkSkzJ++MzF/L1qCIVFT8X3z71d/6W6vtwouGKXY/T+39kuz5
2kO3Wo2+mOLGB02cfya9sRRpStmlmNBx7cc4q7Wqx/7hkIE98gMa5yvL72/MzVY0
Tk1IyfFw86rNAH99vuZwK7foFQ7xE9hEzwAdrFfMsHyX38I1YYDrE7QB6Ckg/4YM
3NkbS2ISFjLO2MTuNMXz0i0HbuGZLnzF7W/EvhOMJTIby+h9xigq1APUBKGLDI9M
T4Cq1VFb5RMZmpN5vCFYNVhBh7cxO7NwG7KuL1/rc+BvAbwxlsCo3omPFoSmApkV
Z5nx/vgCdGalvoyV9j7MdTYVkWc6BRSGOad7vOkEmqKWunw8I0FJD1fkyuDfHqk/
O7DpGLfvhGmaELtmXloOKCK4AErdMOMzYsHZqF2+dbkoTKj3HoXBE2jDwcqe8BQj
Cl/USKmuTHMabl8mdYseMRTGvy7Bt7Do+QNSrMppe5M=
`protect END_PROTECTED
