`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cySp6qtQAYFJzSpWZV9o8MuJxuUrR7GDI76aR83Ku39BD2gAbjsgztJ5H2z5YZ13
nzArSA7yOkkxLVuu6pKucR78KN/t5p0BdT+S885Pxnpp7ROt5/tdraq5RToiMgH1
yau4UT7vBLysupvZ/1GT3wUtsd687XOZ1ZyY+/uCNapQdhFdMH+mOSwOVyubqzlz
UH2mjxg3L/Pe/sk1sLQImaBfcOMoYAqCrRapHhj0bs3DnSDglFW1171dHK1B+oj5
Xg7iSrpudg6P4wdTgUTQu7Ah61lDrA8ao8s6ZROdXQKR3+BwAwk9bwJLcbzd1IFO
LtFaIvwXYGxhT0PGQgGKEf9by1Iiu9/bJagoq8UTbW7ZuDWh4EpU2+lWdb5YWnRd
9ks1ID1LdlFnKYEd205PVlgq/FdizEv7Wdcq8KksnGZ/ltj6eHyRe++aj0FZ3EuP
BhS9E1A2SBYma36Bik3hQkH9KCTtKap+JWarVRgg+bctuN8dwaLAR3WxIeb1enJV
37EKcOBndM/iTRYwJ+kE97qlHgA6N6SZ2xwwEM0fKpxR2PxsMpDOCpV99SYs9ANb
HWub1ANQPl9mFxJu18N5itnt6tXBkIRC/DpNbUtqeiY=
`protect END_PROTECTED
