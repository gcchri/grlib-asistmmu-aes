`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ugShSrC21s2K82CpZ4ihSJRaXwvB79DSArqA226iW56TLpFw1uGFfgLUK2cUCi+A
ZGRtY8uup6ErozgMG3nnfkzQV/15YiXHSBTKZYNhEME4jXqwOaEs83Fzs4vQip5f
9YHrP8KkaqzQfvuMBnZodQ1qalNHxBonemzHULM7lpE2uGXZj9Oker+ogKewuUM6
Os12lM3iG7Skk7pOcei9rlFbSrKEkxr8F/EpBAnG2VwinkFKPwMMZWZrpmeKcTSt
e6yeXcqnlZ2+h4u4bsHK6Dh8JSWDkdocClrb+MQ1u39IEwz13pJGexE4o7TIT2gB
TdQyhVbn/LY9CLGVXkFhYlTriKsjdp/D/nKuMFX+Tc0nn8cBXMJZMNCZEZVE/6oq
ZQXipRmIs+3v/xVyNgcsoZSusJ8CjIoqMqiQqG0yHsrT8JUQyywabxE3oPWexvvr
umn92MLstrI/cBsIMWHRd3SjGbkP4FrnEDTiaZmtf+6GQkr5N7oZBQSSIoQVgbD+
`protect END_PROTECTED
