`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yYvFvaP7OPlUXyCPOtxwI47xhW+nc94f6muhXNMFlifnaJNNEoqXk/ix2JJvT86E
x5mosJfkOnVGxucVxsASBQFcBQSuI0mPWAyGomklMdANLGa+rNein5fgPwy5/v4v
bBwe8BjC1zaSu2xl83Fg4ruxdum171H6HNTqW8xtPHfT6wsA0XLAmYDpBH0/w98W
B+gmSON4BiLk9BsKysQtRsm1LyJhOkZJWOX8Z3FGg2w9/XgTwTmepc/kksHwQprw
8n4oiHwFszQd7X5FexafToMJ4IF9F1T0/0uVPC3rUj/lb2CnGap4ugXtvGk6Etg7
EI3QIdbLZwG/liuOF5EPXZ423Sto4sVTmjAs0a3qoQrvLaGyB/sV+2YvLsFMEjjC
NOOvegAn82CQnaZhIFjAA9QIgHLzQ342DACIMvlCkcl+hQPmfsuT9TxYaskl3z1j
I7DOXp5M3MmsRy8Hiu7V/BABoboH9SwAW6GnjI8TSfit99YVmClorumCYYdNXTRw
MnHHZ1kFvz43wU0SlsEeFqsZPTcQU52x8dsH2buZLI+bJ3fd9Wp824CkR0FhJ/+k
1je3o/qDgysk+MQCaRCZH+coutS/nZD40jHXDLbhDefHX3+iMDFXSpNQlOAvWfGA
mUDQP7MHKhXy9JvBnieFJYcHyrs+AokZmfRygyugywH38KKq4hM+mana6NNKqrB0
IHDvDa91lxCC7zM/WD6F5Rq2prh/NVtfOG4Vb/UvRtkXE4gf/H9swKvYzdSAX9EZ
spaM7Iq90GtzvjI7hCp+R0X6KM3arQsZTT7rPo4M1JrJs6JrsXEtQNmIwYyvUMP/
gi2oSlzAwQjJHfNw/ArkkcKLacev/sdGHirhnmGxPbR7A0j5cekxGT2fyyvVEUzW
0YvkxAPA2wezwkMK8KqGWGpHmzLuKdiH3c6RqRXOOoYUMk1Fb4OneqQiRNIINras
ayjBKa1ydUcmTciVLeLGt4gRrt+LYQU/RV11ohDX2ebDP38DftMLr4Wkep0OJoJw
A3rnFaNr2kdOarZxGoCntNvrW+6/GloRM/eYqp8ZAT7v1WZ7a4IouAWy3tbBgQrt
`protect END_PROTECTED
