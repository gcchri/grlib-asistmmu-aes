`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sPnk0bBWEpqV6lWHonyQkiDRtvjb7zZjOyElIFywCfkws79ItlBsBSnjGY6gCBZ
5X6yrNMy9TPh76Ae+K84oFjjFlPVCUKgc1FvBICsM3Mv4JcVrnZL5VpoXL5kvlSi
RTB5s46E02NR51LnVMyozOOa5yPjCBGZH3vrA//Lrw9CxOlqmmWvLkL415U/L2Rd
nBLrZyqh5J7/QuSmZi37Tzk9Bkb8guTXc4KIbZAUss9CnKzrSck2qmGACEDrOS9e
UuKV8NOEkr/mjeMxO73PGMAMMrzwQ9Pbp9+CF8Z6u7Lka2Eu9AH8qCr5rFkLpiKu
DNLXj78kKM6989KVhDsJd4AWbFBaj5kgq8JpxH3AUm8XoWYUBZEcEOr5own6iME/
2boPd3yNdiO3CNkEAzHLLfaxB+5BpZ43U9h8kCma2Uxrm8L6ZtCgRIt68uFCESn3
U6uQaTOE/xPogIxXFv5Kx0nHnYZ/gnIaRzdYSFY7Apb8Pf1XaZRc7AlerIYB7AKe
vyoHQEBXBj23WMiP9Gys0Se1xT+p1WfWRsOObM3vq4TNnJqeLioo1mN9VTJRYUsI
+J7wlqMqj7fPXmS0dwtzlK3r6pag32GTXwvhSER2LeTjEkwZ8Xkuf0uzfs/2uiHn
bMXLa4vYNvcDHy3GXXo3NXyy2e1X+0zDhU8lgSEAuvYHuVqncH3t/NIsIb0ns7lz
yuy0ORDJQRv35IVBxSzawfUDqkWSAssyl3pcRKR2Bh4JOITzygu9BCPQ/uxrdBMU
1DPYwZHO6Trx5C421mjZ7vFiUfwFu2bY++4h4zbtBqrIl+h30LC3Ijn3rhKQ7vMh
3wbj9V/A0o+JS3GX2OCGeck2Ihswpa6uW15L9gmd21GGSVT4X6n1cVD1lLFtMI6p
MxGcD94t4u39jPJlWtqQckl9xI88jsPlmJuq9eqrNiXa/G7x25buE+phnWwyia20
`protect END_PROTECTED
