`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6NVI+k8YE9oKPFy9dqW9kgQ0tLjpcTHkzbDxiRk9JvuIb25v2eVzwpHt+2xvwQF
QJa3g10GjsRAHRbcZNuaPMHo9y6YFDMXIQhia+avuZkZPJsdQn+wFxSywMjeDEho
vL1RHndjzNB16x33WErfmxtFEeEc5F3htnkLJOjSTfZ0k+dyAFdulKAr9k5O0Jtz
1kewMSAeHEK4fB2zUEenPitGi2pQ5lPTiHDLq42b1skYM3KpTDqC2OsXFvndBU2P
RnXmOOkYsP+APJuu9XAuhHgsVK/2IrA0p/4eyFSMWq+Uek9oap2x2NJTrClq3TBV
0UHS9guREo9mdCk9Wq+V1/3lQx+VeVsXeJSoUyGIi1NOOYlaBEZmMYGf5aGg/s+v
JCjeRfoYQ1lS9ZWGxdiqQYcvEGJQBydQ7Y4/+C1uMH4xbUvLLDJ1h3s7BRxVphUh
jqIMozT1DrgyDh1WYmFBbcYL49mU1vyd/PqL+1ppKUB1kOGDRt7e/GGsxVXTR349
pW4V1Q089yqQtSlg7rYcDu/dLiEL1vpUhwgl28tFhAc5ccaBLJ476i9n2joz6lZp
SV9AAYNihmBgs6gt9Fx/MNqoXpfeFvvqAyJ+0zMSn2kZ8mOTt4Bu08ogT6SzKHXG
6WcICG6H+zK6WhekwspS/N8z6SFJKCEJr2Fh07Djcwx5ur4TBXepfTm7dt8h5YPG
c5IaMXupiUIBN1qOeSj+WBWkCjbR2+OJkBcVURifnI/5m8gjrV/aW0jJkaLe/7Xd
gADvejM3U3JI+p2kZB9mfvKuDav9ksvzu/wthg1cgedQvg12lye/1dnElK/MAPPN
LwHYXSUFxy4v8x80LcHrdHga9qtZVRR72UxR34v1AXCDiB0xZEkVYZ4XKsXrO8KZ
qb536bDDG8Dbd8MuKHEUi4TpUG478Dz3+5SKDRf+3kJoyrmuEdAi9SJ35hzW4UrR
+XrK34QdI2c44p03AM4bJb0BUA8AoVx/qK4G0itGM1idpmpxpZoKTCRKWKcUN/xJ
cvtC9HXuKYDORBO9Tl8/SPoGuLPC2UZquU/ZDKvLoTu7teQtnY2J+Jz5AqOdihkR
vtuq16Qr64b9Ext0kSBZkH3Twck6JU2Fh8fcOQzp37y2UC6SKVdDgwM+w0XIvVQg
dag2vF9Izj5N+ZX5rKPby5mY4bIG9Y0txLzTe6dNtaGHblL/p4/0b7daxx3Lptu4
p5btNQTIaG5MGx9OByw+FqU7UWpuqahMZgB2ThHCERsmd4JQpZCaDQ3YSa5PEnR8
3aCe0iL705+eDRGpvMb+EV6EswztW6Q4FtxM2lScvXfT9bxhpfXbq7rAH/td0KsX
oeq5njVUHcEERgdwKAxac2paJF2Zldx9ESgNttqh+KXb7Yn5tcH7lMb72ELIidNa
iXBdr+yS5KtcEnsvUI1CNeQod40rzENP/yYoxi2t8Bvq7XMyu+s0zsNM+bhHAyrs
mK/jq78ZlIBJp8fC/CkhKVgg7XBPYHn1Cuq7eH98aLr7gsA0DvXy04INviyQzEyn
4ZAMcKjWOrGPR1fHLvTQibHa1iFWC5gd3aP69ogiQoed13rciYVIXsZZAK1SFIfP
KGN/0wWyAx7No3cGGQfh0HI5VYIbvSxKVABYvKhmQgz4NzTAtEVOmCt1vq9C1Kgn
fEslWLyDKVnFWgRx8Hz89r/e332I2VV1xaYWICToPBzK4yeu9iBezBPhIoQo70gw
Pyy6svuhdWIPv56itwUl75avHgFh30KBJOEfxx/nBJWEWEX/x2VtCfAcD45Hr0UV
jXyDJjugqZirtaMZOICkoywAyve9m6uXfwLkFJhIgFNYuu8Zq3p4ZsupJuO06vv0
YW3wKCbR1NEBDLVXEVGu4EudNbaWbDXTbRULGHcdqEn1JyLyN4olwpvL3YOgD+iJ
sD7sBQM9h3NcaaULxhGsknTHX/idDFcPpbuPtj50+tR/8KI5C/DBi5138PCnF2pe
snvh1i+U21Rc2hxoPuONOGY5J8sddCfVY5si7FGQeELhrLUDJb7iUsAWZyC6UHP2
+m5ji8KIwOU5yk2JRwhoFTaMLO/x7GmeOW6zozTsCAtH418g3exuMBWR1uq+h2SM
+/BNPHGYyZHMMI+JWLBYsflmpSUFS3IPb0f0oD9WFHEY3cniZp9+nmjDcs2xySMv
MSH1OFvpLT8SuDiZOBnFEWstYilajnJc7xvlfsfg7PVn4NzMW2jV/MRAwYE1lSZj
xhlF0OC6VqbZO3evMQjBJHrMASleauYXsJ27FpHzZwDR/SzKuACnWQBQ9+btxmjF
K+p69iQmSGmNdUyw+THYlW4R4/FXrY2vCC/rI7kv+iiHRDOHJKyw7B2dmOex1Jc+
Bm2B3kAZaZmHGYUNO2HvdB0AZ88+NV9T6KqZLSLu8xavly5NvjipAPHQKirjDd8g
GeNsM3m8nEz1dcuqXqdWfKf27oIdpkpF2WFhQKvJJ63f5IdGVnT4HFKAePRuVGzs
d65gsM+qtwcznlM/v0XLAgEwhwGIQiFo1O+wp/6qkbQVbSw8hn3eh9px06ITRMHz
+Y+HbvUzlQSTvQkOHKx/b3t3aLz5tf25tNsYcXx9khXiXqnfL5icvMSoja3iKk/Z
VlStvXYSjQwIRcV+KPymIueOuHr5R2QdD8QDO7qYEGW1/W4LYslsmutmbn7PveoC
JH9WGiHOKCm4Sog3aIdo9B7XsUknXKmxgXprU/eQpG+rVmXj+7dBlNXsmvPa16gZ
B9vkotKI72eun8sQW85quqN61WREBqlknkG5fvrcZH0JDhnYyR6hxY11PSZII+sV
wdWLHgcv1hH8APd3f2TRN6dEun1e8QtKjQVPoyiTOC4rdRfm0/rlKcrALujRjTyQ
Uj7zZNHFhIrljBaYfKSb+Nn85wmTAVPVXAxgStOvHr+fSQtspKwSo0K3RaXT2nmE
HcxLiGfZgRzZI34tMsOtzzlq60hfXIE3ZClkA9q9Z0PnmibVO90i8bRJwNgMXAKM
99v3jRp+B7bvVOUwjbNdthCgfmY1h/BVRoyLwfIF01S54c/QS5rP7VwV+qqDop4L
9faUoDsuG5XFcFxPlrcK+A526ZJkIYts50V9XTbS3w+3eCrGkPNWXqAzoHkCYgbT
WXczAQLqCaQeDlJ4o8P/XR2gLyO4BJB1CZX1iIZGAMQBMg70bPTWGyvp+a6e9Hpa
7jSnxkcjpu77ZXy4he9xY5QvWt4En2gs2k4zS+N/wn9murjZNSo5w/y3A0LANsm2
IUwZmMc/81rdJ6WYAO5mMLjwOB1Ys02iXZquGbq2iQ/11fJFzC1cz6HzfPDrc5Zx
k/MGnh5Yd8GteVBlls6uoxMTi1elft7PXmpGmwhrgDMSY+b8672lZIRKRgBB65XY
GVJHNDdlzRoOKqlDtIiok9mYMUDIPaPIPOAJ0O5WATgfSrs76kXQPyYLr1S9LFtw
72BMssrwhroFJTXnd99P6RqAp6QyxBt6asUmcNy0FyZdrAE0qWwHBuU0jRYDiUbF
Ij8iFNAdrR/XuqvVh7vpkNcRyPYT54EJEIBBn5oaOOM4p2EQxndEvODP6fn991+V
r2TKqH6lTkt0fH5OjqfqcnkVyAfJ6VVyJhbBWFCPvp7EqVUPi/+c/1qoYF83L2pB
7JoseHYMFlabw0lN4yxGg8jctLU4n7ehvi72SbqXUTsVfQJLoo2KbPWhB/vvWIDu
rbTDEl0K9hKfAOi8eSECt3BdzDU8Y/ywp+6eoeBMn437xdu+rfx81Ogb9FlQGOsp
EMg5wafifVPuBXYy4eRsMSsl5L3EyMN8a1Ldm8tUozRhjSN8KVhw5p83jCG8LKHP
Y1m2/YxSHJwawkf6D2kUEa4gVhnUBPIe4HCGAPtwtj0sHEyPVgxd+Zw4kJyUw9+L
UMebXbDkb6x1FBjbFfZu53H3zTh+alIK+fTNPYtMHF+erTF6CygF+WgrBcY+KZ17
UXXm+swvUFhP0MggpTd3o86ZleXne8QziNgAjI4TJgBgiEYPS5ppjRxFEEajfYjU
EF37i6DEJqBVBErLGc5yQdhoguTEOBT1o3gJ7l2h6coBr/WNrUATyxQBtrm7Q6TM
pmcjXM8Eh+LH3b7Mj9R1kdpwwJGShuPknWr6iAq4CZbMCnlDOgVo4EE67LnXsvbl
e+/iXoNPGnQgLo+ziMVX9y52fF6LXEvoCP3rV9thgt9qIjvPkdI3LND6Qv//IUIB
F0qQk+7wZsuRNgc044vT2LdL9vT/qmxTa3pWRKyoiDS0HAybsSqRb6q7GSXT+jlZ
Z2Mp5+HsP42dnuPPgWDxPdGH9F9r94BEYpbEAHscezAksuKbJzvAFQ4wRXfWwk0s
23ZwWyrGi73vrsgme4Vhp+wQfHzTpAHHSEpSLP18Cqfq1OXCldfaY7XnWPaH4ICd
MlgXp6cFuR+HS2cYGk4EPubVeMXHWfr1rMuFmWD0ZF/JLqauwGomu6tGRtmRxATM
CjQssIEjYBtxbmQTtHe2TLG5BRBpO3XLjiBS3ZjaPmcKEqc8lWY0ZkFP2RYf/I7g
zUhF6in7YRb7RtVFXhMUWEKp9DW2otoy7Ff94G6A+URhlfVxvqrUDgMHt/6CZ2Tz
1X0/5Z3N7Hbn+subvLVVWR3r4vhhGGDGCvKx5/Gyje1v5IEeE7mH5LrKjbBWgk5R
6GGqhGo8Q0AXzVxfAEIW2rjsMQazwUVd5Bnm1dZbsttp/rgjI7uAju3mROY9oaRi
9BeH1eU7ri/0dAv+RacRp2eep/meNL7STy7ip6UptX0bu1EKopU3Lxeh0GeSf/9k
WigZk6j379sLElT/VLK6h88mhZIv1JGX7owD3d7NNEnYGBOyhfcE6PFRsrxBfEFX
wzfsvPZ/ltjaRp9cbwZZg4rklcqX3MroOz24DclBsUvm8LhqC5dGAsJg2/t7Gx6A
Gplic8I2mOTmoRYYW8tFAWszh26BTaNaj/Yz9J5u/OJLmNCNZd6tPUuguhZwYbNC
DU5ub8zEa41rYURTdz6PPwiWKjZcNJBGlnLmwjUTx2S8WYOvpB/VnhtQJwlvWe9p
pB7NPz1UigCWcKdzioOiBP0/6k8PlGxtSWC1qLmSsRRWSt5HAPGLZdtpHwWHdqHs
EpO7Guqlz4ExAVev64OGuKS/bnkyM/ZtmNMlq8cSVHnao7I8DMaxkPuZI7+SD1C5
Lf8k+eO3HNvqRhsuDUsEgNHluhfp1rwjPHUy4C9M8hm3Py/5IN0gUKEALeE3Ik7P
ryASomEH6nIqhVyYv2VK6c3nTrE6M+n0Y4fzOfIie7uUHnUbp+/ouxkcFT5eTPib
KJz6PVdYPbon5OAxiQ8sfu4cx22nU8TGAdNEguOBwxllLgcXWiD0+ObIxAM7JtP7
+WulmAxZdsVH6LdtWiQFpAgmYBrxuG7iMOoFt7tl9xnuGLefqFTEEWGKWttMjHeX
E+mmx2RtZroWqyUOJeO3jxg0Gd01gzwLjDPg+F3OWr6yvbDwNlqFKWzwp8bLMqZz
psXQXShZA39fOytg3EsgMKu4hJejir6LL0QV36kHvFla0Tc8Dp5baX98QMAU2RFZ
9Z1pJbrqLK8+a32vrLcUySe8SODc4aYFNqHwz9EpeL1MXVIqM1jO6aYbE8CgGkEa
U0uClUN7JQvl6iB7fN5wmJEjq42VPwGGlSHZ8N4JgQTqNYejMV+I5Of2HNae0uYq
1OHBiyXNPOOS7OD49Ix8PcMKUknbc9KTCiN7qxOTyZN0DP/xLKpeS4xvhRgSRp+y
l5P/SOKpwV05W/ue/MqAaUHt1F6i7i7HPunjEYQ57F3tui3ormdmNmWWv43AlBuM
J6/jhSfgoBN7wJkBkAG8gtTB70E/P3JaI3+8loFKU792Dyw1SIWp0sxgsgVWRMLA
oKYqHmgXe9my9LE5rUtUZGKr2sr72BXfc4oN9IdZJFvG8jrdIupaJF8G0H0DWoxu
1DO6e8AentdmqrquwpwrOe0BwIz8jUpTw9e4J+frAdhUFJxbtI3490HfNsrStX2M
Gd06e980kdTOEQRSx3QdUl1zkbqU+Rm8d9w0yIUDg6Ero+8r3YnJI7XC49LqokKy
EC4ZH2z9ptLrFIWUj+bzWVmeklQOZojBNCAguJKs31QvyFClL/aJV7CCa1/W7mG1
1S6NvJI15aOari+KgDha9U8f2Do1/Qb4hZ7Kniafe0ddofJe8z4B1hChH9rudH0K
gxvMdaPz4sRmTpqbXsUXaBEVnZGQKU+Ajc9UFh3Z4siGw3aGmp33e7D0/7yBJjm8
Ju7xR+pBnqWkwwunq+6I3R10Dk63nvTDANFSlsn1XFCHhe/Y0uT0uZfFY2920z0O
622EKj4ShSKsMXCJ5zz1qLjuQJ1PfnuV+CkG26YxLJquk+JDm1Saxh6rUL1Gaofk
M8qF4DyYkN1AsiZjJLG/LmNYdUO2QWLXe+no+WJaD01tq+d2++F7G6pzItnCeOzg
vkTm607S1neDIaXrsF/sl0x2uD9/3SYFw+Isa3TWpEzQvyqGUsAfOcMTu1gtWL//
ue/ucdAUiWRj606uDgiC2VfnWDSl1sgtM6TFNDc3fu0OLGwYy1ScPyQ4InG91B7I
3BqSDdlavyX7P5HkDJBqov5ornGgJ2beXK6BHSfqbBJ0kUsq4k3l3moX3ESKYnlg
KsnzIfiQDgBf1IVwMg9SaWtNamdnfEyKvnsceVJg91SEmtrdMC2k/iXi+adzxPXh
MQuqRBW0uM0eAW9axoYZesi8+jM73oFyGqhAjv/+X/xsYsnCZ3uMF6BqwNIflWrq
I/vMyyPw9Y8QzOxdcl/63RcQzpu0qKOvUJRZfRuNHv1eipDZfi/6sVfz0QlpzLfT
H4OFDkym9SiAYD9IW3XwdfzsK1+YvUwGQMdv3aEH6Mx5pfOH+ilLXXXkRP1cn4HX
WWjzZRKCXxr7ybOLGXVRwT4OtgPkzjHfw1Mdz/A3y8ujaFB/qLJFw+5aG/uE8Xwl
i2HRllDy5UYChGBmVXDYW+21q14+0EkqpBrMQVZTH/087mRxWghzXTSw3jMeZ5k9
dRyR2rh66EiA70shom7ONF94iknyLKfVrmWC81QrLoD4qstQsq4oRZTY14TmYje6
M+jhaOTaeeZrDJ65JPrWtA1KBCCDdY2dZDljohPtRW9EMLl+PiPfP9r1YOCySASe
HUje7EKDUmx7DRn4xr6Tu5Imo0HbTv6TSoEG5HjoNJ5VSfaZ469WtHglfpplZv5E
BzXJE1MnT9GfNk/2gjNz+STscW5pI7EpfKEW9ZqzP4g23pmqOcV5GB+/2JDrtQxQ
x83XNrD3sHHwx76IVza7DobLBdGC9zkER9jBwDVnHo/8WoruyjjlWcmIStnvR7HC
ulkACjvG71WGC6D2qMJ/4P7dRwBmEWoiXrV4GO1AdBQQJTE9n1VKH4Oymnw/Vww8
6Gl/xsntc90SSY/wrX6sRl1FKbdyNtgcbBBVvt3ETzOIUf2vJx7ph9Mj2+mLfYiS
EWDFByB/MhYTpdLDqPCGQdP0JmC5R7Z+0gnLdOev4tni0vxm2b94r+29BAaWqlsd
q/KN7PrcCpfxLdLtvIewKNBO7mDQDMNJ4BcpX422VFI8Lu64+YrediY/00ClGRyI
IPXB0jn149ZrbkRz+U/6gDHoiv4pDheGIsuVLX8ZKVhWRC6i5iw1cyS6sjFJOnAE
nlYueHLmsb+MDf6NoF44diJTcIFBzoM6ThN2+Bkh4mMWgou6cm/Sx/BDaYAr8HAL
yrGtH9Q90HWApGQ5bzYuFBuav4qfF68h2fwIKYS1rsXs7kkfwp+8f4n8coWS1dyp
Y5K87DLW+BEvotGF9XCc+esvY3f/gN1X12ITaAOKggjxTyTfiXGoqTc4LYWVXGFI
Mbrw25qAJgV93uNJfDR2jGvtS3sod3qY5t3DFs404kIOjZfTWiK8exTenZ9bwjGD
6UyvN4iv7/NUf/F8qj1rTrrYs92Y+3x/wXPjzAk2hb91XzBubP4DsUuYYnq7k/Yh
4rj7Io4hrgFyyBvbkx/JqaaY+vzMnlfG48WG2jEmZSHMah6aBmNYQcCKLr9wMlHA
xRNj132DDmNWncD2/eDKCguklVS/bMJ+IpcHfIW8FRM41ImO/kqPV+sowd/1P333
NsRzgsU/S2KZE/NJN4XDhF8rYhJOk0gCvVt1+0KaT4LpMZ6FX6IMRmblcQrfqZeM
UHGFPOlZajPblrczOuqs9ilAIwiz9c0CMTEpjfnhLwtofjyxB220Dp5YOztr5SOy
9Y0oD0sZqzEcpg+2G4QJYgmS0gbSH52aEw2uirsc9TtWyZB26oXVx6d2Mlp8+QTS
9/4+/+I93ZCyOAJpbmoLhlm83pJMiSpauFfGWwq0IbsmibYZuK7Tgh5UVEMI8CYJ
mW9d9wG5uMLbBF1jmWMaCcir/l3sqqqGzaAZ0zqzUiToqYEejay8HrTKBWDyzXdi
0DpZAtZE2dNf/SZRZJzhb2zSiI7NkNkdmkJHzl0yNrxd9cKKyJ0VqnkYG0yORMyA
Q8UMX0swvpiusBToaDY2tp0dPFx4VJKj5DZXBS/Yk46Igp5jzC9LGGV5dyCQx0in
dLgLeqIk6HpgaDY7RgI8FVjInkR3PVBF3xpJ4FljETul6oGI/bO1ZhNDOxAdD5vC
GyNUj9z6VHoHxp78ZUOdFSWpfDOwd7Y3VzkqaKgfF62v+8a8Vv4ADRVGILQakWbt
gahlfLc2uoSd22uFTfpkJOiUtkzkmhKCjmKCJKwlNSwY9e6/fcipIH7S7w9jefpZ
ONRZBwYINV2QOugAwSWFMc97kK9RsCSGGBhz3PnHRVx2hvrAWAS+Fa6YQ5lvMd2c
qWdeY9XRcqL9/f20jH6VelJBvwDSbyNlyvq3MWGuQAarqQ/M2T+HfdrBa8VzPzqD
iDc59UPgUPRfcwMBzQ0Hgwc4fcalhAvPZR95gwBDMwV96LejICoK+2A+7Z32pGfw
yip8smlrEqhL33Gi4UbzzGJcsNIVDZDQ5yZ34b1zQ+S637myn3Qx3SW6PxlUwCQo
QIXz8fxNYJYyQmwsED4CHGskC55mMfReymqeaWgHgqrMgk24UsqvUdRBQpePCfvU
6IfXqjOUc2HZCtTz1yZWaRyb9f1LirEfZ2sBaZc0GI8W+YacfWN2MJPOd8V1sAJq
X83CdOpudFiPFhu4M6dGHXNSSRPDrn3ROx0gvDKuuVJ2uwbKHlwKqMehSchy9NKZ
271wbRiPyX0JUMfIbWn5PSF8XEmXw8gD5pJ8kjSeRAJVXb4UliQ/7zNaOi0cpxLG
quBOVp0BiUDqJJLgdyz2QajfdpeIA7gH6sL2wh1EWKUMlUIKWggizLxEinFfgWFw
s67C4+sDWQLisDkrl338g0U+L5m/ZAy/H4p5u3j4SuSH/LGnvvhxbVgNINyIl2LX
cJkRMhAAHZ1Lk9LlpGl+lQ+ADKsp/yNSMiBFVOqjL/y9+v7u91yMo7E6txQK4uHE
7nOkV3qOnsMgWHi4CxRSRCKMAnK1d/u5QaSLNJKKbqkyWdQ34vrMQtiCQoJxYbI9
sM0VR3dvO4PAuJqU2KoGL+U8NqM00RXvQY1eEcHohRnW1KAtRaKWUnanOTixymJI
QIUvrbWgNBHYUbVfPIKAVTjFz1qjFx3HeQhySJ9ey5+3wz5KVN17k8HGPW0ACCF6
D2+4Vb37MPMuJXTOdjnUPTLNyTU17f7LsNdiaktYNoaib6lENYfsBT9lblYW+V2y
RKbWOaElo9Q+0jNbkZyqmdE1tR979rlYMZuwUWIsVGaXyOQe1/8/AQ+B5xwulXck
/9CPbO8pRd+lX4bP9cZKkGk+xyz3G/hingxPSu5P4ENiTOlJBAD6tcjlflRzsFE6
ibsFG2K/Gh1MwKdrV8KGMUnDbLiRQbIPe5iGbQTKMrNWvAaQf6K6w/XlA/iorKRB
YZ9Eqk163LSB3TgPzWyWnBJnoSHQsQQrwOMN9smW261OBHcP6I4KoJvmWjX5T7S2
sftSyCSCiuYbbQr5TxTfwK8eQbg9YgOZtTAXRsszjFxO4JaJ5z/Wkavw/C+xWkys
a64Qsuw+pepE/26UOx6mnz0n0BxYAnSkZ2xyJeb04kRTNiQt+P+sZ8FqQTv+e+ox
k4uXalVJSPOZTfh8Knsr9F7OGGNwh1z+6EX4aO1vnDTB3cQXtOwi0SD9U1HzWTKb
GthFkLsd2v4rUQ2KwkBE2ZTOq2iet//OIEzL3aTe0Y06iwWttM4qmLDAsgoSpSUJ
Pzbukv72QrZzcMB/sKPMRkE9vcqU2zXf4KY/e5Kqvi7KrlNH/wEEQo9GzWFH2xcg
7csIIcMVnjCk9G4nSjdTyjAdEmcLS4x0dFBKhyC7dJVK1kcFLfas+RQWVAoHgd7N
uSRhqiDK43l6BqE4pcS5oqpBsn/DIeV08mQU9LKprHH5HYXmzBkZUeOhJP8lYQrI
nm7mRYf86wQy/hamijsoZDbtytzGzqV7pD0E3ndU/NnO++6CqmbzQOGXeCeD+Cjw
tDf6FAGujUn5XxSaWkZlatUkRML70qZIdNLjUSGNY8cv0zUyk4j+AzCw+6VrOV31
SSF8KNVU3DQRE/hAx3GBa1DVTeehUcbBlfRrvoAYa3Jp/4wiaNMJ6grBnOu04Iom
XKx+rq/BAsPhMFqKCBFDgcO7KIJ3syhwTt3rWR7mkiQ7mxB+nH2jRswqNXTyi9zT
V9XuGxK5IkbHCDoaOM+XC4uznCnFzBUwL5+yGJnOM1yL/a7wOd630NhjOfvENyJD
KiZ4BaHitGxyHNrSj2qBw+OkxI8e8yubG5nOSYar4zkDzd5hO14H1E4seeB3gRVZ
qBqXm5Ap8jSbTjsFONNPfbgCARY2ci0cMPOoR/S9LGgfgmX52IwTh6lnwqchE2hO
+EL81tVpgMXmcYzerq1saAq/TaGS1iOMNuB9+HNM3dpwGqEyAa63Lt+UNK6ASWSA
oghUaIgQlktLf6wBD3DGEJxL4ZuuU8rLC22rm1XdPJDvPnm4oBu9MZFtEiC/uRcQ
0Exp9NlTfz9+hoBRVZ21L82Yzf/7UGZ6cMn8XwcN8e18AqC6erud/jeAQ8E58bkl
rfTuXxwD5nfQsT8dop5QgPZoApErlwt+lgxKCPvHcYCBTj7fr7gTs3S5QbLIvOfr
3U+WkgyaajPQO7MVXYtWpmIrdgugktVnOzx/nc4yepIrwslZGqzLCOFHtoJBzSxz
D4IoIyRK8FVs82Bv4bvzMptclrrgdqVz+VQ/uj9vIYEyPfgV7L0dpFJ07gresKT8
6gI/yP/aVTkvVVyyX6WI5GOZU+07zpRAc8bVthYCjAzRx1QhG88bph9Rc1qVgIbG
ezzTZHXHZ4ei7ghlQy1O3DJUM/bStAZHUXWqiFrTzkVIet0T8PRbSOo3AM/CWn+i
djzzC7K2DWumzF0P1IwL0WY5EfdaUY7yr3u088iztcRXzKHJFLEX/cz9UmoJXae4
cUlapUPgd3zlRdwTFf6JaAy464e820/ti1Na0xwLUjhEfp1TyvdhsbVwcLVVeSqJ
IVjkGvPfY1S/aP/w8DVqc50+HB4TyvQRa6XHu34zC+/pAGE1mm0dEsFGUnUYBLx3
cx9d/jOI50lukcBUepwzyvWqZSYcFl7yz2nhvkLqykoK1qVJn97jQWCWZ8NjIoya
RJjabZK5m04qmNVlb5gFJplRaiDTgZ8t3h/p5awBN1c8Q87EMF3kWlL6KVID99F5
hBITFyhG3vbuWVDhwzcdfrUKxc28DryRdgkNGzJFulTzn/4VD9m+TjTB90N5PBYR
OGAmGTSPbBAkziyLerKBgHh1AkkFnv+rn85m77GO7rs65XsQrVEzqeRaE3NWLjL7
O2Mtt/ujCoHTZvlaC++CRM2W7IV6ioAB7FlLyoMQbhhEidqj7SMYTnom9VBLHpWn
HYf068goQfF1zHOL2wnE6iJlgXteyp3oBoHiQnMU3X6T2FWGhlY6CA2e4PQO5kSJ
P3CV6+BY3hnayuTKhUgwOEfDnI9pQz3s9CwP+JCUQ2F/hSRugTLV9YiChwQ20cmO
tBFu+MABxB4yM1BKX6aDnB6ZBe2Xk5dJeLJiCsirdlvTd/g0VH+vUg8qEhXFzVFc
cPDeVe+CO/7IdEk7Ef6+3P1wm/UOA3Mjf5zHj2Uc4rzuxJfK76K9CQPmR9/wQbpb
i/RuHTtnPwE86s2XI50NXCW0JYl6PDQPCWsFYT/xuSaZeprE1VF/G4F3WW6AagQz
IQ3yT01NcKxDAp2cW1oMwM+dCKnKKvCbDvBa+9VBLjPbl5Qbu9qlu8HqkUnPcESn
FngukEZyYLA/Gpr1OXz3PR4XPkAZX3C7Qatstqjoq5ROLxsaINQ52aZIwDy+aqgh
SK9537qpQyQ/UixwZmJUjy+4fqMqXo1D1CnKlkbXtY7awDlLP32biR756fG6Leh5
R9EOD85H6B+RCopgOQgNSflL/dBBPetQRYGK54E2hxaH6GVMrQASGEDAQHaMxpoL
iHXJx1zVdRGKd2zLieJ/61O1KEliK66pBXToUpOsnI7B71C4zLH6Yivv057N+n4q
iZIkhuuVQ5r/ta24c7IL24Xe+gIG9BETm0yhb93CLnekhP33db3sOz+FL1H5NXEU
M+Tv5SGH0DKgR7Gcm6mR9/21bjb4x3npVLmZy9/V5j3vfZyRDIKgQyzi5ZUXlRVi
28uD7uOPfRn8m6jW2Pz2QgoJJGbSZFn2tO8XirahNfOFLnN7W7e7VemzVsRK55zH
ACsQuD7Egh69Kg21j0C7IMGEvnfruOvUdlI8qvfGIKWmirSHkUwIelqiVcYTqqI7
Sjsb6B/Y3PNRVfPhsvtzJOYapuZlGv5BzsF7wDe4HbTjkju/qy4TTyUEQD80K7U3
vh49eq1PnY3CRtXhlryrVZmdJmDdQOfxP9Vd45fAY4R/4xcHczorPiTk4MYnvazV
W3MA9OqdBItbPm+OzfawqranOFbtavJ+WWJQlMMiMyioUt9zQVjsJWFjFKu6FXb7
AbIH8FXCmnXTznU3gRYicRS+0A/ugixAC/lx0iPy+QnGiRdu7LfeUKol0KVLLc1N
S4gWW5WZNhzgckthVpNKqW2DxZ016ObFsoCszMU9YHTzpHlBr99Iw/KoXz1mrNPD
Onyj9KsqtNFYNzTdSHvz4qOw4VEIzvkt5tEBQ6hOfVs0i+z0jtTdfsvmNy9SaHbG
UZy3O4bZIAlaSPT0u/mYFani3R33e0/aqBQFteBGCiQEABrecUbxJ8AnCg08VnCC
caN+MDeX59SkZkZjTSOA00wF19qqwPjXlAykN/DDekdY5CUWNLsr/WGIiKpl7Lpm
QnO+MLU6dAZLzLfLM1yIchijYIt6TgDIsuQFy24Az1mOgPz1Vmb10A2sh7TkjY0F
pzFzHHnSXOmvhVulqyoziR2OBcqjd1JaMy5dl80fV0v8LV+xdVsXt71H8eZy6DfR
dZgceCMCRhqXEZwUkzE14aSFTslCdp/5hXjeLBPAEIWoJvytVV4Yesqntz6yJJe5
zvya+weWDl5AUp6uZp1XniTD4lx14JIE7aQG7++U2HyzcXX/ymeSMf7spl6s1Oo/
SEf+75yrhWtG6wy8ySowvbDNlfOTK/u/Zpv73VZetnKYpKbRgP40rm1Y5yQ3IVGP
CqODQmqbFG9EN1Pvj2Mq5KJ73ld2GyAmcTxx/xDiVp98YG+zq99OlQONecx1KKCs
M8KulXulUMVuHBQRGuuFkxEC2idsc0I5Z2nDk52akAhZlY2CygluGgc1XXfUhpjq
P3Mg1F9jga/3/9vFyOuBiMolSnwMxk6bZ/mlddY6OrZNdgmHYgiqk52b+Jn80PSH
gyTp2J9YiJ6ynKVwqHj1/0pDF6ykT4Ig3xbhD6G6w+cX/P4TpKZEV7ylCLst/tdr
KcX5mUvfATdHIUJicuXZp/2I7R8ao41B/JDARVS6pWR5avZW2t+/JFUYEMD/tylJ
huUQqpXupbWXAMP2CXAzXfVndY4ZkL2DGe/QJSbLUW3Vhn6GC0kk5YeVnxmOja6i
C3ZCq162/ZOif6/qhF2D9WUmxpcnoc4XU9AihO4UHu5XIrd+QCoNrrlngqqkCA0Y
3lPAEuPyZX58nPiT5g9VLhigTkoW7pEuns3rD2Dn7HfcnOrsqrA6YY6RTc/R7Fcs
x3ychUF1wE+RjSs+lJUCOUujhSPyCd1KK7pz8s8oRyMOQtWDBHk9un+aNEf9Aedz
xaUe9ivgZetdH55NbZWXdC1c6dRNhw95C4zz+fy362Q0t+KKKaSllmb2mLGS96lx
I4iI4q2qff+FVJxWwSoo2RDBZ3X397TeA7iJS+q3XzRbFw9QHcGde1Qa0Coa3bu0
69tkTmgslh3vHEu9dAEIbrNSErPL3EFWJpHpccsZgixcPUwl6ljSAvM32sh0V9X2
e2nAEd1z1YyQZ76JXqbE6N6SwutdLVSZkxuic3QGjCrk9Oce/g+dTJ1CtRYxwHdN
i8Aw2SkU4Ood1j2y6F/U1mFF7cpNA1Dx8NYOa+sSq5T8oF4KqrC1H1dHVcnPu2Qs
4vvyiuqGC668rzCFXM4ZB9HhqFEnyoemEu3kReG7QTo14Un650j8rO4WYgrE35HJ
yrJtZCB+RpsiQbAt/l9lHVpGKPq76QtCr9PSoRBObFuwGr35kRHek/rsJQ5pcFR9
bE6LUM45kTEFR70jfJ+IxgjGO0Cw89sHixIVhlyazirXhGC1KxKNdkqTHGH1629Y
QI26oE89DsB/SCPvKjMNvb6AzYMhiuxRASGvSNrxnTuBDpij1uM3YrKdhBOgD2uv
8cdqZAxy4plSGbk9aoD+R3eLp/MV85ohg4iSbptjH5dVaEkyV5305Zx4Sha9+qLJ
eAXLvXOnBYDflRO7z70ouDmWp602lEvF4kxcyAIU5lWFCI7x2PAcpNg/IKaRHrkG
x7YraTlFaicxFQKL50nHFP+7CB5c3mTR4zi+Rwub2fGxRgdDAnn4G0fGebRd2MCG
mjAlGkX57AaoNdPwpWQgu96VMkKhthKY/6EigUbs5ZklO84jdcEcjyJeBSXOUN5O
7iaz9cHsjs0YrDWPCwQyDJ7Znre592r9Cs600AqW27bkDYXaqDhLn1dfD7Diafhs
bpPnvmCJjQCkKEiw+ScBKABfFW0SEp6GlEgQyDZELXTrHFewTwp+hKHk4bGzVyUy
HJ0hwRK2POdkNw2MNZhijNTwRsYuFJR4Ay6ehSDDvEpoJSgqgwFwBjxrwIdEvEy0
B4nBHN3x1SCWgbRxxQDtN+Sd92EyfPF3z1W+Te+nCcX5UFOZ8KNwPCGNFhIC4A/m
rK8DUNNunkxKY70VQnOagfywXchwI7w+Mx8xMgBtVXnwZZSRjHOsUy2MdjONoTSV
L35WHwDQdBG5STBZXLLbE7sZ8pfaPCUvd/6wPVnR5U14xKCPRx6SjAl9KvD8wFgT
BMUsVA1VupWYLZ4hHR9dMqQ2ifKTIqqK+bWeIl5o6tOrzwockTuPXMZO3IPeQ4bQ
J+XnRniPBZ9LVKyCxuOW2LJQEKqHwRAzwrKtjlqN3aPgSAZqMB9biEjAKu1ZHJxL
QzyVjgixM/cOXqXjixaErL9BOKQgdkyIs+tdlzZHHCGdVjBJEuyf7y03WkDqVB/+
7mf9m/9fNRaPf9l9pz+BNBLF+/b9q1QLMA85zzQ23zuMhAbwQ2CZ713acEHO4jtM
SIA0fncf8ckV8Lqgwlob6X8WflppQ63eQBTSSzuQCoJiUwYryMgE1tQMn6ohf+fo
XI0yI65AdnO8X9vHqJiLomXAdpmbEDh7EeBAGcngpk+JseYN+XONQfFD+adsV36a
IhaV6kpNgqrC0l87IfX0pkLLJHLLiSeeT4RAXVwOvqTGsdIQ5QK8SIfUek165oka
YO6i0Mxr1w1LTdXxANtakbgXR/0Y6aZ7pUv/GLUuGNYS5yeQx1YjraZsR07/D2Nh
clW1cOaLM9lm3Gi8bx1iT2Z7GTDu+klYh6medGgpl/Wk8woZH3UnDPy2siVOlb6N
L/6XQFXeEa+2fa4wNvi+EBa+XaAekaeWthHcTR2+jFoWphdr/Vwy6VTlpyr+YqKB
E+P7X1d3uBGdLeBmNCVNpD8DzFz9pjgC16iqf5Qq9mez9BUx+OMES81OnpaE4vFA
X3/mhaylaVLh71LF1/39QOZkubNM/0TpR5XhvOyBFa3gDmIkQjaE+wlh9e/e41lW
LPC2vqC7ZqvSY82rszz9QkXgimBeyKGKVC6pcQDkg8FqZS1TE6dsdpq8/JlZAM8w
Z+2VCDNt4PSknYA9cr5SiagWAOyBsvHPVoJXCFClhDDWK6U3nXE2I+CrUm2q6HQ0
z9lRUWWC41AH8JRebLztkLDgZA5S+ZoLo7JZ+OQ659qsUtjDDsFT0QeiqMhHYdwu
2qcdhwJPfKh7CmMJfw2qKK00PUuLWSwxOqisAyCZprAss64pWDoO9vYB0vQQ7Hph
WUMca9WyF2XKegPVR9KvH1VW47urpgOt8U8K7iAp+gTG/sECCFxsclv+sux2mrYp
AV0pAASrE4ct7lgCbgqoofAb1JGO5q/L2WgPJrO7cNiNCOklH9w3ZUlSQs+vuHKm
Z935xyZi187lEYteKIL5OmEN2PRuUZCcTAtnx4dn8CDma/iteNnLFumv2j/wn+eE
8hqgt8i+iGDn3i+TrSJ+7CllcAs9wz59vRV0u0t4Vvx8hB50ObOHEaxGkfAGFkpU
aOSPJl+XGFwgeSj5xxnNrMruBuOyovXpws6mwqdKSNy+JEvw/fDKJDVEesPLtt4m
FTHcTUQl4hynKlQnGtuEBKW6slq0yqcYgjsazHTYQi9/j6LfTnWSAeFARNdcgjf+
4jl0Sp3Shnwo4RSoOfbq4znE2RvJLwJTJ9p2WSK+cVzstvxSDJl0EilFbc+iQUtA
6Qry9m4MdS8k5pmdEjwPt2JoKhRag9tPJQZ7AnH0E4w7ySN1x3HDOcKcXojBqBg+
XkbbbMDjVLk/rw295Y82AzXok4XuryIEZfpCgbpKRyfWbsS6NestlhBNSsZrnUgP
CjHGCk+4mGbEffnnXcROhPR1jG6FYb33YS17mIv6LN6jPACBdfPbJhLy5tCjKAmW
9Cdurklo5J1LtBbBVaWFiz3GzI87dUSJGyaIrPUotGnQvGlCsYH9f5iK+b/zl1xb
TGh0R4edIOoAsnG/6/2KhCO9pAum1gjUMU22riBfkn+UzbKvfFXfGNu9qJsN+hdk
dcVI8Fh6VuDz9yZ+5ZwMXN9HVh6w7/8TCcjPTC/pATzQXmo1IajtIhACG+3CQM0Q
LWRuOtAH1CMJBeOf53HcXtAOgPR61yxGa4xXUhvTPeY1FYDiPLi4CPSfRboxABiI
JXrOfilildiJE9u+n8joEb+HNurEWlHPfl64JTG3HHkqwoMhZlI2IQO0Q33PYfPt
//RfQ4+NZ0ic1ePIKQnv6QamaUIei8Z1nSnZotfldb9OCbksrdYgSl36a+1KTQHn
ZMSH91UMdCx/igozMq5q86L6hqWa1Jog5foUsHjqKq/FkItVtB4wW1BY3cVNfAbF
cZgNKCuV5vDARY39L14mF06LtpA8md7wJ7ixLH7+98oQ+0BxTlI5jkTz1X7yguvb
ro6kXjn8IB3LESJElcP/2J9cDvOZz4Y3WamTP6ki8K4TqgyLWDTTtoRG1fFbhc0S
1F8g5ErgsVHHULjBIwsLsMLj2Iab6wyl9kVrjUuqU2yZv4gP3DQ7VdRGh4u4y4XL
Yn3X6nrCln6K64/aBjR+r7EndqOyqaYX1ryqF01jipu7AhdBMH6fo5hm1H6pwsV3
UHO+vLUOSwrOB76aHam2sODZ6Q5+3888E3Te5OiqxANWROJQ5CQUwLZoTlvj20iu
eL5ZycrFeKcnqA03usC5tEIES6KTfUAvVmYoCvekysZbXRi6QLj/AKMMhEk4TEfX
H/k9fIsRt/K90QSfcV5hgafD93op/pl0GN4yp+kJUnoXPZP3XUNe2Pi/m0kwdben
4dPgOFljFWSUlp34fmuWy1jg9BrI/b8t0OSpOEkgmj/fTuA5wwf2NcWh/hFbEQr2
DLxkShNj2Y9MrLAJA7L4+lXeN5VPVMnaxVqtAIqqeadXgxCHfsRpwr6KSh0EPAJ3
PIpNbQGMw5bCAc5Z8YunggSZ1Vvo9Pvpnlz2LtwE5fPQkabR7cxEXwAfcwsvGNn5
m/QbhYKUNMlvjRE4T5/hPZbk8scOtNKEt2OUP1+6Mx8fLf6K7xAgBGt6VWMrtgMh
FPo1Zyd2AD4hejQv/SBD+CbLaLUC64yhLiw37EqzS74513rz4baClQNDySlOn79s
OTmxwsTP7+Cj3mDawhgOxGUJIXlrdgVMY7pz2c8yoQLqY4qSxyMkfEpPWBagxRSM
jnMRXSI82+GlvTq6J8GOEaGYy5vE9kR0eWnwzqRjVc8owU3t3iIIDS64guPnuBk9
sNkehSkibPj7dT/iopSdbEqe/YXh8tfIQkGrsjUB4x/ZoGZFtFnHOBJt7nF/H/xy
76LZTgIGYIUQdvw4Dr1ibx3Myf/Avp2+Wmedhq/o23ikETNZIhOW2oVJ715nC/z+
kjoRdTem2sQ3fycqLRHC8zr1O9jOIp+OZrowwnsRX6HrH7LPbrWsB8KrqTJWCGpl
vDk4kqXEoCizX4+bOXNGQj+dQ2y62ubdXnkX+6wwuYDs9UTxyWHwAwTvf38z3LYG
oqbMJm9HSEGONRzKAK07hP2oiEfLPdd++eC+4JjGvea17GKnfVCwKb+5NUXoeLFI
4xGsReQgeDOSOj7a/lPzK8whC8i5tltjVDDEsPkACYJmQVskcwKMid4gMtQf8+CD
RDkOKSOX3w7oHpwyHAtZ3koJ0ngMdz/s1wxUR28HiNEStMS9CNz25v2Uhqb2hJce
5T7HD53E26zBE7KfQi1pEJ6uvvjPvma54tHbc8R7W4NWLP+ueTPjD4jaFz/1EB2C
I7PWdD4iWehwdEbzIMmsypVQmMpW4wVVZ/Im5K+iPBTWwTNA36Um5+NjjlGM2A2D
f9OEycIEp2RIibQZ04/f6WvOqv5wxMAIlL5Y5Liw4RGw7iN/2ZnrcsJw2HOJzIPJ
uoV77ZQlPmCImr6RQTU9x/Qf6WzUPSXAvC6u8yx19gBlnRw19G0UDJlsi+5YX57a
Cc8Q2ehIf9CaHcIxV3yHUzV2Qmvmk4hjH7LRDV9yoHvCRHFJX2Zs+5AdGc48lgza
fyPqmj3PXyoeBoFK4R+dPpEy0DOq15/Bcjf/plIqAaHsSf1vqWc5z7zRgeXnmrLt
MbpHNXqFIg7eOa3vd2kbvevX9AVrb5pm1Uh03eTjwSIDVmXdzs2Sry34OXf1zVXm
i4canlZ3N1WYqmsTgjn5Jj1VvHSic6fRYn1xlWrtoaUeIDQy59cfogYy4y+/k57H
aMdXHr0cnYz6H5c4zdx1i6mD4Pk3ZT+mqxYCscNkb83GRfREpgaFsL5FNXgDS5Tm
DrY4mD56bthJM1J553KbiAIlVNhmSBnLh87i1oJVPpEWOWUbFRyqTyF1DssahoGN
y3Dyyj9Dj9aVsy8MF5iO8gNkt5t/bQxnTWF5vUKR/flFgxT7SaYBnUXEk592cf1U
k1GurDWd+vgBsb3MlVpcrs9en1EFj9eRQdRK1y2vuLqKLw96Ux18dXjxmLZ5v1pi
VfCFPhVJEVGTI3zo+RBpc2TQ3ti2G0B1am2pKxyLxgk50daB3j+6lC3Dk1hoEP+j
cZsFwV4oG0F1XDpkjUtyZ6AhK/L1xy19R0zbq3Dq2aqOr8LvPuS9HqhE3ZiFYDIX
8xadxvZ2Yh6/AeobaKPRK3a77cj96814ih4CaphjUCxHeqjw86MDt12SnBwktt9j
yyXTWqsyDO8NFwfj93RcU2909JGs2sgTC6Phc7twWIUqQUDrFH48JSIQvEw+S004
YTrVcwzS5rNS+N1FY78fdezMkKIhWs3aTCzX20kjhPSgrT6v6pQQ88xXdlTyQN1T
O9ZUbDCqE4lh6d50sLr+6mEuDxG3f6u7ooFyJVKeVZBTS4qHWZuTupgFgzBqwD6J
unrDBDAqI0LvU+us5GkzsLspQOqq+/IVmgSFrufBksLOJOShx/mfTmTjmoUfDuO7
hp6PR+GNmDJ/bFnb1kLv0V/L/1ro0dQs3+7GHqi2J5wEqbStHvCQpejaNeHjyBZm
cZiHW87/vG/2+UQGG5NCxaiUk+/ouXh3d8F2T1JI9Y89fXmAneuZ+TkzY5QPpBVw
d/kLRs1wWCHN9qC2TP64/hlg6rp9lpz7f8Q64SJ1/yJ3f5gnpFHwSUxF52EC/24l
r6xv/KxNh8TWBxcJrFWj154JIDZPwg8ZRVsHKH0iacBx9g7dZ8WDh3om9/YQPPe5
TIQP7Djz61X9gLL7YWNmbUhV0g8E/c2pOOHjr1JQxZtaFIhdOum8c9fqCGGddktC
x08KRbG2VkLJNeAYCaRKeyWjDu+2IPfsg82oiEcrJ2/ATEwti6ePR4EH/Fyz3yLH
18umlKhoNBulXqQB9bjNKxM96gj9x1dHaMw1IdmdBVsKC4/Dw9Bk1606YDfnSLaB
9LXTSwOSzFqVbSYNGDMYMolx+ER7gn5cu8twzuR/rwrpJEnLiAvh+PdgZw2eKPtV
8rxztwWh54JSuJHvfM8XBLfq8g68NffEiCqcNFyQFXVPr9dtWwSyP6VU100mV93/
GLjekiWtkOhJx8rUyAmphI7IYUl3U1xO2a6gzeLnmki261GqXXIMZW6wqTFJH40u
RSPTuqQgvcyoJ6laBHNLDGZBJrQN6njtp76rEa96JomM2g6So3pIsywionBhmOWE
Dbr85KNVtjSMHYAzxc+GpNdVMXvnkejljHPtJxZQ0KYwnJDFMT6l+bxENgjkDFYU
Ey0cZKDEd44LJxHkYFuYlYzPLfhIYyQf0kKydBMy0zdxQlK9l1WBdDZHWxw/jF4o
YocOJU/mMsW2s6Ph4zKt+KFqX/aeN/gyw0tWlysO+pJWUtOwD94MZ02OoopirMlz
rv1vYJ3EySOxcSafczTr9FvM/GJFiYaGDDUpwwVlkLEWqcI44ESlzQhfjOUdHyZ2
CIF5Ruakoay01soGrpYdDeohdBE6ZXXYI0jpMgIScG0I7Eh0TuldAbNbWfsuU1sq
Q2DhHOc2LAF71+IHBMiqRktlz16KySEcq2xdjvQXrJqt/HtHPkIw+BUnGmcZ4/99
HLRXufN8ENWzxQThqBd/e59zkR0pSdFnEIr4bTmUmAVOvFubBmiTEXky6D4mURAt
UK7jIyKZGLFOosIcfKRkax5KSdt1ECvPJaRGkefGFiUiFJQE6FpIBM5VrLXUwa+z
Xa4XTJVnQCOH6v1MjFj6oWGiS3duHoMMwymlt8ToOAYuOm/rcTYzScTQWlW4pOQK
fwWa1pXpUSUEmjJmrTDZ7XCgNb/suWQMTfcKBEtl6Ufgsb7GOO7qkF9jSeheECCE
XfhdFy2tkMXH3i2bJSb5CEwVIA8U4yEaTAvlVbbOOfmzXfznGD46XRMNXc+/yZ3U
ywH2uL/LAaIUxeDYQIA98olLkW4J0p5fvK0TiE5Qc5z9/lYjAG9cpU2kSPDLCjjT
1fSDrpvKSP2k28TCCX60LYoLfEZYyzcWJTBg7hwEWBilcJFfHouzBz4wcP5Bqor+
IuhCrMEZJbtDgfGFU5mRHw3b07OmR5UuDmmgpttg3WQ/bPIb7qT3d7bnUSG+IQBY
deTRH+HSl4yCLbeGCgRT4yTBVgHnS0qfkklb43m7gTrAPR7f9l7LMsik35YMriQ2
Q4QRN0PxbcMidAK5xp/PSSHi2WK9xOLR0NZwiBBE5kqGKBl6j64Y8M/pOchJ8x95
F9JqnZetuJoryFlhmiH3OIDj5xt0jSwd6YPq4Kk+AQJ78REsOaj/WQkiFhu0mKpk
tnFZjS3jOTsSCOPmoEtAhGzeSscEDT8PQUknl8fXMjWBMy6BG4JgBdiam2Jzi4Vp
IgBkvH6FdqqMxayEM2Qii7HcHABCPQflcdWXCLF9S5diDtlJ0P9ROKxVfHRYlCvy
PWqRDs4Wi3PUCgdsr0X2gL/QBfXA9X6vpHy1TXqrGRdDGoQnivkL2exh9ZiR0JYj
Xng5sATbLNf1Fpr2yF7uf3PNQExJ9Hdt4syUiev++P2LCwBPQI/FHTTwSl7kBsJS
R4QLpmF33mdMW7U0X0wk05HgIcOb4SVyw3yQZn5gGNjFCqaO8BYZETDCmA61ByEO
GzGCzZ5Z2Kw4cEA4+ajZszConTYKdNK00XJib08Vuv0eyp5bJKNv58QsGuh2jVEv
69cCOQcqNib4F/HWq7slMy1ygEXn4QkFBhGNI//pYX34TX4MOSzj8xRlG/TFCf7u
LW4kHbKLLm4PogDiJM1TY9mhF7yTiexqYnXq37kAAE8asEnHHfRSwfkFkB4QH9Pk
hK28xNskrQIffyOsPeA3ziwugD8ZxC/YXfvZGPCNoNCGuucaxvFyIBp1Xfn7DCrX
g1QNdDiDcpXxuzrugVDHq49eMB8YeL7KbgComNxVMxwn6Xf4P+EWDutg1XCTk7ZA
q/kJEZpERi9A98bLiewnV6Idnr4E7kTmMNJ7R3guuxSULYwDWg2vNwolNJE4KGmR
rwaHSLUhs1X9qnFNr/8VsTWHVbe/WUr0AeCvJx/KjQmQvq2f3BwN00fyWEN6KQdP
Fffl7Dm7BP2D87gXH6enk0UGh6xckE/DfqqYEBk8NanJVx08eWxuT6s40O6UEmFE
qI/8mMUyPrsvgw4jWQeRKPg6Lkzcmlf6NJclmzl0LWEv9+Zdx8pHf5DCdKZ4la6U
IVNKGp5kz9hPkqeodo+aPsYj6M82IYfAGo5xZte3koaigaM2jAIQW/C8OuOWfphm
hL8cqNpXsk6tlqgZyZOACPSw4Q4eeNnRv+kgQyHKT+zUWc0hqdkEAkgqZcK42FZj
OTSXccz0F5mla23ftRixCkmaYV6Xo4GyzKddkOicheDJHA4KJ8FbxG8gGhf+DiLe
cD/tny3uG1RvTREu3CGD+zYEgO1ouypmnf7XNy9zPuCE9m/+Tdys4ETIQPRJaWmG
xU4Gr4Kn9vobUsholok96BXgkNGRgEVeKVQYo3ENwbN0pXZAoEH9kUbm53oenVwO
neFV4dtR/nQk+ljKUVsaEPLoq3tb3uGuAhVZi0XjeFEoXMdFXETZcurq7SIgojpT
KGlYJr+LtSbjx4cz843dDDx9xx7ahiFIny9EeAIBi1KMiq2XycZIr0RzqUZQIbcZ
GoZMf8ULrrArrCSEn2MNcS0gOP/FrB7PskRyHEGugeyjusBjYQxMtER77rQR3juC
DAM7G25I2NRnj7NMVZTZq+1mYIjrZWAIRaPnrvY2dCag/1BEmfJEk/Y7WFBGKN8Q
oXFLfVGf5+c7j+XmKe+r83RZni0VogYGdVe9R+mxe/NHHbcH9vlPIyar+NsXCvpx
9GtNwmyVO9v0OJzSkPoQ32svuYjwpN//5LJpjwrcZ8+Rk6KSKmjxbEgDHBSGRGP0
tcZYiui8uFbTv2DrfXF+vgb94qdu929L7dYVgB0Q9U5TVp1V7w38z4FmCIFcjcpg
mtMwUnhlCyAdYKs0WCQeoTEeomu4saMsFxg9aykMg1d8b4rtnI3k+Dcn+YpZFmp9
Vr+onTYhdEWT8jxMG/VdE4FRbBMfoILHBrBicNKfjNQ7uyCe7O5/vcs7a/vjdjNN
Q52MgisacKdc00N7TGWR0EHrkawXQAnu5VaeU9ty9BH2Q+rkNpzzEAIGw8rNeot9
R/B7gWoXVbwx4s503Ukddvc9I5BmtAeKQLG0jhXbeTIqOe19f4UKaZpTa6gi+7Ta
jpQZpxJAuaXpj2Pa170f2XL1W0r3ce6R9/ajCBJddi9X+nSd+CyspLznlzANfD7O
lUZ4ND22tKmzvzoQu+fzCCMz/5NoR+YrnXlgtIzEXeBEvbnKeXc2E7L6Hqndxycu
swcZ9k+YqhewUU67HCYz0ly1U0Msn6cqbaxQUzLefUObhch47qKgO2TgIWQwgMJr
HwEO9390AYRxFnFZQoBxwUNYJ3ywDXYkVEQ3b4z7bdIo3stLAi0yOnd0Ra2neAnh
j7lTVJR16R1eFAPxsb3SRzij1+j02y6SIw+mTfpQvMRL36sd5aMN1tt4Y/bBrIVR
Y82HWPuDIW5N7M4/peyX2njBj/AYAH9rPGRmKEAxgklgCFp6PzPjA2jMhyeF46aw
lB4TGJ/HfbWKB9wdM02npCWvXA4Zqt2e+k0a0lh4CJbI7shWzGp0iVHeZ+nlUyPF
1DEQSn9+VoLfRh0N2krDP6Fc5Tc/EesRt4yiGoZeMEt6hZDo2v8nKpTXokJgBodH
Vphs5Gjtt4Gfr3dmuvaTw4N80iL4S3DJ410cCS/GDyRgkkRYukxNdIiGpZrMAR1Z
oEzfg0NsQnths4sK12xU4XNMKfEDfWTkHp+yD1LNXBJhM8Uo+fHEceRvDf5hF/88
iDuoJ8MWMUk7fqy6sGgzLLwTJUriwSrp+nq7LiT0xgr7Hf3EmzIchF6ygGFJkg4m
jzX/wbJK1eq7aAheeD9Kw9e++rWT6ZuFuD5UzbXU86MoI1g2bLqhbRIO/tM2h6PH
o0iwY/9StEv9GXMlGg5M0TRbFsx70wE0wk5q5ttcGo9po8WXulwVgbhN3GRmZhp8
qWH/CxbwB9J8TJa8A19EL2eIh6rMmXKi57vqDyBww75dAmWdE4mTNt4YgTjMCtfS
yvEWgmpdRcyPNaTpddbbRKzehcD3ut/feJzmlvK7KpPQaQf1LFPUvnOIn9FZP/WC
kI5ZjPB7IKlWrkTcYFeFV2fZEXcUKMIkYsnihpVjFEwTbKV8lKR7U6cXytH4uOrL
Ck9n53SzbzTEj3yt7wT44YbbjVuYZ4tpBjHd0WRt0o52MT+PZ5r+OEExCV97TdjQ
LLS3I6YRM++bUZEeXoz/RWt++5kmPISSoD7YPcuRTvfaDsowB7V8ThCjH2ouFsW1
K4592qDyW4CV4X8YMuEYaDSH4+Dduh17fb2mIdO+qy7mP/ARmsNQv4RT3C6MZ2bE
G+fjkTr8In8xfgjBcfkhrDTDiFkaQ719X3p/rZqTpol+smQQwAxGV8xKKVpTlTJr
x6kYWlgyR0M5pE/GzYDFEAV5dv1fbwvtvC6+zGG8pKPORApKQaMyURz+nwYd3XCY
c9uzYGg7Q9vxv8Jh8j4jwa2clPNfYsQtrNbUy+abJkrhNiIH8BBTDE2PG2ZBe+yk
KcNrTNc38mNlgJEJU3toqHnPAlQj4yxBU0F5T8fR0wmxhPpB8xPiwSNDUIohB3r/
VYeHU7AXqdBxlcxI9r5x4QbVA7nwUreQFOV6tE29gbNoTWrKOpkn3kddcj/rkYo3
CVDnX/An6YxS7a+srBVFcJByugbi6i6U7qiEtQnW9lOCkbKJ+Mg8rVrKzYZdoT3Z
d5pmOHD2Nnhy9IDQjLZ64c3ZeJvtIrZrmuVQt6vByxNx605Zm1GMY+4Jqdw420M7
9OEaFYMvPBXOsjt/VpEGWDB2O7SURJvdlfZleJMByDA7Z6tidm/Kgyam51lUbzR2
k8Se/yUmv8FONvH4GNtAfau7Zx42aH0vSSBpcmIH5KhUEohkpFEWcEcsELiqJInT
kWQEMHKRoJ/ISVOZM42vk2vofEbqHPBnNe9asP4jBb0trteZBPqJeeXwq8fYi9as
zSbyHTu7/nDUqQaJbjtwIFKqZperR3rbmy3naPjB4cDvx+yfcX9iHeiHvtp3wEhV
Lhm/P5Kwgr/cE4SgfXkt4TVttUytHdp5rhhIreN0N9lO7HApHjQjbLzZSbRqXHi7
LQq57xm3DFoZKz9l8T+yJT1mrQalen2nswyKlxll3Mk7Qeh5OgzpqNH/ymSFYmsw
r/jlTWcwmA1F4hhhMYbWGaFwkF5GdfTgtXcrey/lhOXvrZOY/njnhjtVsd7eFelw
vrAzf2LE0vp2pXztMzFDMTGLUwzchKi2d+vxjBkdNIrB+gwTKAGyaOEBSzKwhTra
LKjPLnRU7IgCliBZlG73d4sx7v+GCDMi158LNbS1GQoX6nTSZ31hADal/8Gv3Oor
7oveIB9GNQ35/D+1oIhLCpD75Jj7fBwoNjVprn03VxX+dcF4e1uSg0jcgKo/UGp3
x+9Jt6jgWpjZGNydnkeyKaCpnmT3clduXN6fIcd+gUiiBfQ5AEJjJyXP9j4av6je
CDCbn5iMGbYJbebfbXkCZ+lnb+sbgGhvtSmtQzaU/XUIPYoau/FMXNccqEzifMjE
T2XMugZX0fKQ34zUxWOaapExAREpVJQRFrr5vFWfhLFl5ZPkY7s7PJpY+5hJ7egj
n2GuKYD7tE6lGbpyAMr1rJdfaKO2AM1+Mm0Y05wX0CZ/rXhhQ3trSM5TWwU0f2n9
7ciksMCYqA8ZM6VzhW+6fGv6ZVxysZCaGBm3fwPpHDk4ugV+qV/BZY9i4omhfIkM
HZhzOdsrWpt57MbZv/lifQITIyfa23lSYFRfAHMJNazQ0LzMLea8+FQiYO4eZZqc
PqXT5WRR0ii5ONK9vfdvKh/BlDuIdPHcmJaxHR3FEDaP4NqpzVvmDHeVLP5ypBIt
jy9F61D/mw8SCindIBq5XiykwPECCgWiZEprQnyMpDbbZPkDCpjQVzzmCyjuyg4J
hBqUAksTh3EKgm6QnHiUc5HGEDkG9B2SsIMa6QJ2M8MaXHYU99iIRG5R31jGJyKs
SkSmqNoAkp2A+9Yvnlhh8Ff7T2Dw2MXGfpa/TKTRdss0HaB+zFeyxZt5uR8YoDsq
ozMNF2fJDWlaVm8Dw4vHaoCdyC3RwFyU6FA5fxLm0wnyVq5Uj8CqzUOwo4k0SS1f
oY5szCYn8uJSYQS+iTv4U02QmZ6DY1OxO6Ab3r2eZ9uaii2C6YuUK2E1jhHe6/9q
jIw5fVSDSVxEZighFHhtRvnSUh64TpvzszH2biUuuwaQ1P1TjQ0BkrAY58BQsoxP
QNy9UEvRgXWR66u99MCEeno87JfNHMjm3sqWXbLqGCDMxPH8jU6IamDdg5kF5RJs
ocaZKpoRd7/DAqRgbhICVfF4nSYzTw0yrGcz5j+zJ+N/So3vCsKJ1srFu2Em4SAm
OjNkRt74qPK1ddQpH3uJSnrwV5dNs7bYirxhw28q+uZAybKVmzmriTSCwdOPOZQy
lYz6Iy0DcZ6F6ch6gSdc6Q==
`protect END_PROTECTED
