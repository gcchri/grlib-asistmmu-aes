`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YxFDB2GB5fygEOgbmz2gkh+mfjpVfzD0ABuV0Qod+atP14VDjnH1dTuq7JhKptHA
ogK9km6Sqz7vpkCF6LPua6qeEIKu1wkVH8+k39jtWeJ/GqWPErX39wJuXaO60saL
Af7AZ5N5vCqJhOPH4Dikg4G3/Utu/2gibk2Yfeh1nHrjM4MGQNfVrQDhoOII3SLa
MOHY8klCR/i28pbruP74RHUNv3FkYoAhBpacwMVsYpM=
`protect END_PROTECTED
