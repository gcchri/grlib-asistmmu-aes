`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCTYFjOBiQ1gfNqXHfdXYrkM+ixClrazki+cJvB+W21J+TyDplTWcSdGWdKx3h8Q
v/CIFnLROI1DibVN64ZxkfSMoB3CouGqeVv27p4C7ogi5Ae2R9ug8V7JTvdU18Dc
Id6C64M1NFx95mrlKsQa6igz3y0MdNMc8/M9leH/LWKgkLTwABTdE2AoHAtxBAXx
qetlTm7alp0uj4a2eEp0NsbZ/3S0etB+ABT7d9kbiFOkKI3bphwugp+gjvgFtGnb
yyLELxK+bneXqB+Qcctj5Mu7M7yI2yoiRq5aC9Zvr/fZVJ0spTqssC3qoG2I8LjI
JUBxpgWxTJwizO5QYmQ760sctUE1DwSJ2xE0xRoW01lpKzjuyZ/nZvdiDq9G48xQ
i2UhqkJRQ7iaaOkx6d7DjybQxAFunXkBsIfxPtNVGcVZCbrnKWWqkiFcPTiGvBsK
6H2gCb6+iDw3HNp8e2SnAmwddBBP4Gu/SugC0nD3bOk+SD83dGKMBmFwdEJY7BDE
bqG6bnKYtUGy+YiWo0oArnGAQq+2p/xDQh6Vue9qahfJiczlsGMU50mJdPpz5Tv0
F3YJtxLWLISJpvVuOHjuKSl544FC2FAMdQnpiCHMQhEWNIIQ91vXhBu8CfwNtwty
OeBtZKw/x8jkVJRG+A97U5F7p9LYolL/xs5hbSAUvjEjCM/8Gu38gJPM8OVnCUMM
zQmo0jgcz77RGlVr5mFzSdHMnTu7FUf5t+L3Bt6aZ7lOZrcvgNraI7ueMAYxONCM
yBv5i7+jLxrsiHdHfbFlA+X6LvQImyGveqMK10XOTrVeKs8J9WQEdrvmf2jeJ9dm
lIwmoVpqJBFZ2R+jZIRMm6xXdRNKcCTZCT6FF6PfFJYpQ2u3qmQO/f/ao7EuAOT2
cvVsnGxUl3ONalvM7oAWTlJclw8yKS7b1ywiiFDzeeSQZSW2qa+3DCs1HIfc9/mz
3rOhRxB13ePFonk660QfvdC0NVVlrp5nyB9Ogyw1n/RWB9ALrext15WrWq4IFnn+
HEe+/Q5cZVacCzBeQggEHYSNriKUha6e9SuQk/8TBYDc4yunJX4vQ12tuoQyrcPh
D1FaQlhkjswt14lIgof7LoAdOPOCHOkh6MiCfEgEFHvvZNgszH0TMIgrTTZoMmX+
`protect END_PROTECTED
