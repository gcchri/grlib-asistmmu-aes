`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1alxM8UN3l1bN6BNbUyoROMCyvUwd4b0PxPbC4YYY2wjrTi+x514pTQGecjUG52
zwGg3uRwvHjY5m+k9WyBHEvOqCHibNWw12cN2eUPR112MaZ/pgzVCQ1xlNCjFyd7
DMqEv5yS3F5oOkYk/JptpDQZ7AweDY5qM9hRgpPCgp4FMR2TbP9FJHe6x6/Ra5YF
/lMxmHiWVaBPtJAiJWoyJ2tLzeJgKeFNFUC4pFHLtxTf6ibXUt0otT5Fn6BYjawd
20z8K9MSqIukuPVFIEDkQHKW8cQPx3hLWOAaw3gkJlSovkeXLDWyb2oOG11fiULg
LyM4l1Tg/5fInKTbNI5TL4oq1ozdwLm62Sbtglcegz+azFNeO0yoblkF+3OOw0WS
jPH9MDBYSLA8UPcUlod9Euwcxm1bqzoyIv47mt/DL70x5DTDk+R+e/TMG8g0ienz
5TooEs6W6E2skiM8sy68E5kUHf9NKsmPwrvBq+dAwvKjZl6PCaKnNXccshf/jr/k
kfO5P8aaPrLgUSkafq1qFHQ3PO/iYi8UkS+PYxoGBE7Hc3uoZXNwAGvoMb3rfx8S
1ueLOcBGgMQKvcw1KX9bgjN9fLuq8PO6btRe4cZ3QQ9W+nBlXhtKTuoQ0jSGaSyJ
CiSyLjYTVMfvNsBkSdUd0ZsZ9vZfWgQIihBtml0HXdpWC05lpM0O6LTsH4pk+XNx
/SnhGZmS3SBCEpfupVSilXmuDxGOzj2iB8ZKHAeFHp/qZlFjZHyKJI76a8KiKnwv
LyiCj1PShBdb4+ZQxh6i9sFoDE3HRY02F+776mVIodSmqjRf+L13ZvTJ5qHBj85K
5fvGaV6uU1rI7fSdprhLrnOpiU6nsB055HknsSVBQdIAednpzk2I4wRgBzph9TXv
ShxJFyZITR54CA9PdF+FYwPRjzb028K06h1JdcxnSDSBSVH6MMeXOdEf3fVHUNb5
tMA03IAutnFCCAQDbXBjeHk1Gwc8vHfbPI7Oa6oLxaGp39K9VnB58N6v9qZL1AOv
Yg8GS1ZbIex5ZklcKA/vF6CEc4wzxIpiPMNTNm2SBMG5TFtjoFR+EuaQdul9w1We
aQjfJQi2q+XIEoDox+LxVDoBeK7nqZpQJG48pwRQ6aTtuzalr52xejjLlp27nIGS
QBo5D6uN+ZnvOlREKXcB7Fp65DK7QXTrYJS97EvXN4cETFZsQclE7IlJ0/bxXorS
Jj5oxQ9EeObjpszxmid10tmmkjUxFd8nuiZM1Zb6fbCpx8tFAghTqTJWgztflipo
C7X42f0MUiJw2ny748nOei85d2txTHRhigD3djcyJAOG/y61oXzuj9Lk4AHzBITf
SLKFfFQvDgJrfrvjycOu6VQOd/3sDszHtVYvax9614bHzM954G3AANd6elHWeR8u
G6Fd5WTvq1fTkMquzLhvbZ3tlAhEhcOkS8p7Aba/hg/opmzKUdcas20bCjM6cAyJ
kItW+wFPJgAG/Dwt7HdCywwCQvD047fAtgf9xPaQdDg65vrRcyWGAGVnUokq8piH
RirrRwTVnGdPKEXjqJS0PKeOYTkMgmH32pWDB6VsjdQMvXP8GqBHZGpDyfE8+a4z
2dQcXPLQLeFougAxufLjdjC3VZJK2hiXpVJC8bx/PVUfUSoiKvb0LLq6w5fDmWJD
3WB9wS7myrB4zZ078zFAWQiSfKSJcI6uLKR/01l4Fx0Mf/hzxrZnIehOm/sM9XRc
J9/sB5SMZQHjPECQ5Spy4+LXikuwls4cQBTLoAb1BptsoRWURB6oUEqyeDNPD1fN
u7RMlDtYs9ukk6mSQZLCM0Lx5Qc9wChB+twt6BxugEPbmPmM91AxtharaDQy6bmo
pgQZKtUIDXaAaa1tQmA41D9VdG43Bbokk1PbPNxSajjz5X8LCajllrcEbNdt3nrI
wL9KJ8EFTpRmQQPnmQTCDC6VSYrAEZidJH6oI/CuQXh3PZY9us33hs70XccX1IwZ
wbb/zxwzs8NpUE5kVpsNI5PbNksbNki6zSa7UHGGxJGoi50E51yy1oxkmysc7Mdz
MUj7yINVlSWsn5/D6z6pPyd09OjI7I9hwtiM3tdEeDSf/15g6uY2mqzUjLYenAGR
5+yKdcNg9S7dZZyI9l6rL1c6MuR22j6ukbGB7CmjNNFOVNl8ZcVW0iDVk2I5LJof
FMA4b5oPJZk+4MatopFJvFMRCND5GMh8ht3YCeiP6MQbLZAfqYbZTGw35a0cr6i+
+I1SjWsLHJLzsAuebJhsJDNWu/zLAGdoWqZ6APMwKndVFFMOlWDTPmsU2YTEYdpq
xXRmcgf7/uyb5H2hzWPom+ljTfpKWyLH0J8xLPDgr+Q=
`protect END_PROTECTED
