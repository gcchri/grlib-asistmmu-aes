`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sALUztX0ENopSULKmnqRdOCudWrJZdeIRHN5Cp38wiPKKWrIEe2korHpmEo+Grks
UPDls6wKqTN0WLPuntTXN+2P/3m1X9jL8ABZdvM5DfwZwjo6x5sn6JBdtKv7SVl6
N9Cv/H7yr1k+v6ddOopvmnqvwE5UJrreovf6Y7lOBELzYQ9HyoDhhh/gyJMYMvnI
WNwjZ+5K1jbZ2IQnqumFpdJTC5wN2dzvfGXfxyzDAyVN7aRG7TZxPQVG/lR9STbc
H84BkvsAzDeME7wblMPOq4yryRSrd4ZrtBNMayNBcKJXkf//0TIxX6/01Brc/qFt
qRoWtxITweJ8EbEBZ1UzzLvhWdT/NyfrnECbFCTgJmbRr3eZ/NHtlyy/CTAjGAGy
s4V9wzTXf52/EVUs/VhZwyGtanB1AcACK3xmTWeslX216rKHT8GBWdItfofxwI48
RSLHcqNuH1fSNKcINzqeErONjVAriU73LDWk3rpKZ92wD541nRWuj9YDH+vqjDT3
a0Pc0ehgHB5uCdl+doZGpO2DBKE5DsoOIBYQ5ZlvdDLlHBB3Ga5YdlvoatZejaxp
b4DfvBDRLbhYLCAvcXUliLIc3UKAXyXYEPmfMkhhUXvmGJW2EiBVkWfDCSbFQPzR
225avSdZFZy9L3kKGAR3oihmAGDC49F50XrgELKykrCYv3oA4IuFOtTTlR8ACVxj
l/Iv2G9Fd1444TiTc7QdsNNx8q9P83QFPZCFdiNa4SeHA7V1k6ArsUM4cf7qfbq+
LPYkQL6sBEkZVkfaBI11OtVRZoMq7wOBcazoKZLjAkxYGx4bZvKWgS2lRotV60IJ
FjX1+tlKIHs0Gq/+6QxL3xWV/KrJOnuT7Pk8+JJLcKZZtCK+Gq1qBsgOwxM6+J8i
brrZhfCs4Gzc6o3qd1j7KMtpEwyfmjMokVIo39ZSf9c=
`protect END_PROTECTED
