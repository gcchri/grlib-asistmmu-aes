`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vxo1RVKS+I7AyBrjuqG0IDD97WGlf7xGF8CaACPXaCQQxCWybsYVz1LKGap1fpDr
ounyfbZipx1NDUdSJr8N+ARdKwVVTwJh2jK8UPP9/cRLPpM/KY+DJYytQofT3SA5
oHBYucSpItkFPdOM05v4V30Pm4qLpDjpUqjvcjVAYvuakb1lTaoAxbHbJ7SwXbuR
2lzGSnY5l+KE9xILGzHN2oIMoZmapRg/btUBFVyvSMhKYbVGJoI7UT4S0qVY32CY
adVpnN5MXIjJ+lu4NQdsFj/aCbieFYxGnp6KpsPpQYA4lOI5jMDOsZBfPGYPhRgD
uzl6SxG9YcH2VcI50hs7eNni8f1iYQNr2l1syqoQ/QzYvYZxQIiN2sgHEUgAaGR/
uaJHHVZWsAh5SFz3BTZBE6c3opk9MZajG+EtNio1Y2Hq9dCCl+xRzwBJ4INLQx+u
BVx2VE79t/Dl5fJD/c1RGGKhDqVGMCmOZ7miwcX4yWi9aNCpcq+6TYkwj7nF2uwH
8Jm0GaK66YECxlzSxpgVb5DzF0NE3h3RZ58AIKwuk8y5DCtl5xyG1ivdVMQKBakW
BvrF4ePRdZgRtKgDBW26+baA72kcVi1Wp8kS35mCfEamUMgB0Rdk2bQZ7NKJS0NC
u6E7o3/5hE2tPlZVJHgrPjqEOSw70j2d83JrARM/WP81dViVJsgbvTCOu5YN79QJ
V5M1EQA1aWaoBkkIQq2iC9N5FAGuWMJ5ZmTktEEK9Fk7kvU830F7fBR2SqP9NE8W
jXNKuQRScUAE4jzdARmwOucA8PT8ol+OxeZ4qX0MU0UEbxp+dRwM4fw9jCEYX6Vm
f/nyfjc1Lwmux9sfmfS9gDNv9yCJLc806kwNTPAEqkOfSVibVFPGuj2ZPGpgB1ac
41jkWQW4NJLhNi9+ToI+ohQPjOaCKBVJboUoFcVDUidrLtp75iQ7OoUaZsqh5xn1
c88n/qzvpPPVAubGAowDqT6f5FiF+9z9z+b6x3MNY2lctggSovSnIczF2o4VHG3d
BS61gPdgO+tK+QDwcuHY/uDVihzJemNK7qEWlaLDA8EAA6pmM7smYL1cZ+bVHf2V
FxEU9kQB0yXNKYDhfxWBWu9HwIYoxiD0vw22Q17LAfyJFlR6O90KFyb3NkzUkKfZ
hVxpZJRJBicllNfXOXIOPWCIhEkqzonk/pGZKGAQGg3GrDtrNozR1OwgTUXrq/sG
BOPQ1hPLIA32yL+QOhkbDiHZ6S3RMI9XF3Ifq+VX680qBpadtvsi7iOlFZ7yza39
/Popasb0WaqIUV/OBBADZ6KcodTH3bGhHHHWsH84DbTSTopFkzD7ST7JoK1n+q76
9AzyNDgA6BgbXsRUPUt3RIQjfFgxMZ2iGBCG9QXIc41INldNHustIh7Ldes7CeIO
d01p/xUw6aYygCvGBsFajrrGg7VGMZzQU+UvekDgZjBWOUixRWt9D3jfsFYukzX2
56s1dP78PXZHZ7gFkPNu5IWmtsVu0VV1jtNTdGbP1oXfX3aZ7lmxv13nDA8wWkju
2cb3enC6SjQZDa6ZrxFwj+mw/BlTWK1K9NzM1AdzdP7IsAzL0YIx0HhW/HvxxcNd
ae96ElIlK2FywC9Gf/lF5UazUOrZ+HhrUXPY5/RGOxiEg+tXEGF4W/LzWH64YC+R
NXh4jXWvX/ZDqx6CPwe2NQUPERaMQbpsVfPodRT4Lm9YcAW0uNykEW4ivFIsH8oj
XQE+4vt+LtWMc+lcXoVIVyAUZfVNk/MRIoJ5E6YOR+b7T6jXNx3QrFsqhqhx/rQJ
rVdhfKX9OYhmIn4oHArnC4p2QQ3sr1AAFBie3kUP4W4FMnDzctU3S0kO2/68GynB
2DVU0thYBgPoEwiver0FVqh3J8xfg6T4lAUozaY60Va8oxtxDVuRy1JWetOnxLPD
0pnq7V42q4vjfGvSaPzPR34W/GewHlqCFd/+kqg+Yr4MWG5TRGdeZ1oWSiXbd7wy
z/iqa/yRGwiA1JjE5XXaALuNRLHcvQn4u0p5OjCwydFAKyDLuVS7m9P/T/3Wd7WK
L9Xgwr9H5FVnW99piFb22kCCZVWzo7VUBDOEnn19gLeDmyS5uPRVklEOn9TAIsK2
Si6U3s6FaBNfpMNboNBZKkPkcLXi7vYKvVKC/h91v/g6XQuFke1aZlmiMyQo24Br
q1Mzaubkhp4Zm4VSI72/WLlmPKhcOotCXgq+hR1xcylNqqzqKenqgac33dXHrlLR
7OreWsbIfhwPwBE45dwZ35vYb5QC/QmOZpGOwZgXvO6VOUaIwbGj4Xfa6eAQ9yvL
uqviCtcVMKhGo7cnIzqJdTxIXZEucPqa0CiGlYlnbm1s4c2+s3THdVRtJopE7Uld
RcyY0FFhpGArZTx5+B5h5sn0K1zUkAdHLow+MKvUxW8AHToOd9P758CpoS3XGyzc
C+u/QhqyPwzLlO8mDj1WkU4cKojatATB8Di9eUkFadFmFvWb6LOgHLKEJq+sypHH
Lr28VVf2OwClba++hjuEIwmuCNHPxQPnA9YGw1Fe6FmjuiB+vhFWjy8XXs78G7ob
qo+qpdss0yfdbpPQFNOk7ccOtqnBOn8qwEoYycKcsODmGWLilvPZUJttWy1DTY4E
DOtWGdgzjp1wA7vTDIx9V4QRQ9y4IWNVy047qEpUZzso+KTE9Rf5D+QPm874aC2n
C2x/o+uXpsd858CfZJQIQi4QSZYpLZpVx7HIZ2wuJaN0YEjVk+QO0AEoSD6UdrPM
bVYc7SMVX82cKmU1GwFj8JIWjIZYnHluTdRoNXzT15r2KZGgFbMVWzd42UJIx2oy
aIjmVqBTVZ8ZEIGCuQWxP7YRLIWA3Vh9xVwmX2iEcQIToNpFQwKlp/balfahcvp8
ED4+Jb7sol63+W7FFb0VBgIDdlOj7vmc2JaBpfHAXJ2n/SxVHEUaGpA0o8/5cYmJ
+8Q8Q1TFa/XSLU2vI6Q5fT9mxJSDwxnjrN9fHJbWKADw3TGaR48dpfXRj+SkTB7E
JHqf1rzjToxhmci3v/6Qdh1PusVZv6HGOTloZPMcl6gvwTmwzNK7J6aCsoVXDWie
leUOSBrnexUWQZMwdUeqqp/0DV4fvBI3Dgzcvif95yJSrjdIrwe8jlUvHLSskZr9
KEu/H1F3OK4iuOKSNKeRA2jmE0dxZZCxLohmCUnWih7xvxMaTvv4k6GfgG1ah8YV
CasCFuiBDRZ54cC8IemoHw21QzipHn+GcWgqxJ+tGmMR4H1gRbxV61jxEr38o+vu
C1hWPvO4tDifUp9LonWc8Qe0WyUarCNoaArAKoNA1GF+AcexmBrWkm4dTmCkWtZD
8FqCISKos5VH5hWEVj1eFZoCSG1X1+u7q+jDBgwCnversjR4VSaCx/9mJ3NlSmWf
fC5mErYFHWIkyijg+TnKF9FuXngFBYusUmupl488RFYOH1ebpnOcu+GVXEpD0k1x
z/dZZZXHDeLgHWCgEWMBMlWUI4RXxXEonjRjO575WSDdDhtk9XhlZtEocRNYTHYf
Q9xCVakFPHDmrot2uulOjdTyFXBHsVrAg+MqUdMhowRpOs7IiEhI7YpIFPyGZJUB
XByqJNHCcjsNIUihz6UJ+e37oub+V9fIpc2biM/kYPdwdTl6Wi9857WDaeOco7qj
NAZf2U9aoFu+i+DtxUQJszn247hHpeo+ryziaGCI9W507KJbC7UelxK0RS640XnW
tVmssgNELx0Ek/1AZkrS+KnHImM/1TNpygex1XSrOXWRW2QUcJ8R51yn48NcA3SH
Cw93DM3Fz5WMucWXIDm8NTcB9517or2vm7Ux0zeG48tj1H4tB9Zv63rLtWCDTE4I
o9p/tAkFCADfDBXVf+RXS3QUpq1IiJe113MJCsWCwJH9rF2fRNNEuNS6ycqH/pNZ
iLU4HWrCpFnEWOEXDGwG5Rb1flEMY82zspXFyO8x0OFSxVQ7+gmpXs9o1gqna9FD
3EOnt9auSR4oiONvVAt/ZGbqAMtZQzbSDGny5sZKhpe+am2fMaWkt0JwbXR+DZM/
BUfR3kc2kTnIqOGiRgunULPjPWClT9tqKXzZkLTPcCNg2WCeJogW+znvnvl8gX96
BBT2WK/4BtFRhOMBP3aNx1NZmEcxra5mh2dHm4mpXOgktxTdW0U0onL5gChEn4qO
qNOtvZawNRy9iTzvdAJKkVJM9M/OBNcgvdg+CC7e6Uhxr76Fjzj7C9JXswio4n2w
lgVSAvpyb3CmYesxe0alvg/JE7dTo423o/1U0GeLw8Yf2/RCqlXWOICs2nHypnpy
I0723mlfH0rdLYTV67t5KM1o0UcedJWXiqsIvKe3pSpbgXCNaJR9CZsT5sTa7XPP
wBWTSwgRS3LAd27RH4D+d8vFwcMgEe36SyBeH+zfJrlwVbIoYavSVLPwdwpT25iO
8QRiLg1qHEjM9LVHLm0AFV4wh2OcspOY/6gBluNzqVazAT4sBqfzLICBVPN5NJtx
2TfOPepWwEkGefrLltmSC29ILJTjgerxgetp8TY7pEQetmVQ2Hu7r8IYWwtEOnz1
fkJsh98fIEeVZO0Hy6eAPejWNVwj+sR8vTNhSDpbUIuKANDNs+AQrU4OMpBjg1me
7DzehpzvrxlcH/kUwUYAhTJRHBQ2FRnCgk+5JVJ/f924rQGUTD9X35/nYW5/dZ27
WQpeo87alFbQQ0KPCgqT8piTNVED99eiGQdeCNerG2EOa9JbfU933R8JpcP+OWWC
6b6mOFMXPTU8CyCU6bXtmmGFGtANS7dsbO2vQIftHlDQdCjBLkH0D3AnpXdldgGB
yf4ynIZ7cBFOGeCTJFmDhE+WoeDUJtmgfGnJyhBZHIcjqmbwzEWAGZucDI3j4cVC
afxOQyi2+FBX1Dj0DdAMJG8cQSWdebkSTjZtWO+dqFGpNyxDcZBzWwGvK3ffgA8G
KJXak6y7k8OIvR+EHSrBC1WRb4fD+v4rs7eefiUZBIBUpt+WOW5Y00Ui7xGvA7he
th+DbR5Dxc3h+s4oJuTaRAbRG4fDDDq1982k6NCU9bN3bS+4dCv9JkXn+F++zWq/
jPlIuRs6y9DNIvlV4fNz2JuxOQqQWzb/eKwVBc0T4BFnQmPOUBazs4D8krxXPCqp
D5JDTN5QGX6jkLMAWvEtY/SVetaUgDsgoT8w4kmj7tD5LtSOCeljmts09r2+78b5
wTUKDur3znG3WpXPbb7/Fz3ZQh1gJA5siBiA6yDDhYg5kj3h2XPEmrcKixGfE1Vq
ygt23KmpOTZw4QaP22fVEviMpWHQFZWqqYZr0mh8A8z+tK9ql8drEXL38ny72EKV
eOuJgXOHl0hKOHqgZCacU+2yTnOOPDU/dO6NG+d3D1lGlKuKfX6dTlACzhd32DZz
lRSAYXr2PT0GNuZDHW+6aTt7+JOT5oY2FeG5n/BOvhK2SQ2qYoAgQZoPVvkQvrU1
DwymX+zWbkR1Jgv2j/aaBXvKiSq+Vusx/LjJ4e4MJOPULJdYtMaKtJkBV2K73Bp0
qQFF2oECR5lZ2dCBKO6SJ2sJIk+caokx1L25CI7I40xKjRMu/Mnpth6lbmaufocX
ApqFFdyZkxW7dsYBLql3LKbR+WSrb/TqJTc/ldMAPkNRHpUr2672a8p36LhY+tRa
iQTYOe9VD/WzuApP5P3bmIRtTT8Q9NRvED2gTvhQes/gdxIqOlPQN31oraweoyX4
QqaZ/RCYiGsgcBszkrMXd6+6WiAksMeD4pU17R3h+bFwjPvMEdcPW/4hOoHz+7sg
XoqZA0O0zgltEb2ZnlVet3fwvIt8SKSIc5mF7QKYbcpfcxDR2qoXOXTgrSjKddaA
C32ZLUZkD/D694YhjH7JpTRwgaC1JTvh6dvzVSERuTmZ7t3hVJv603Ssw48EGdGI
aowh8AleMN+3SX05EyURQvQ4Ef8DKuiA00PZurYUX+7jUNIoT9LVFBswG55BlKIq
4TT7qC4CkQBQidKMxTeGNXC/V4pwiOlO8sjk0WXk7YlywDOKJrLLi31fdQ8T1b+y
/GvhMqsC0xNe1W7S+CUPuP3k+aJ0DJZbP7qzWEOn3G50wzYNABpLZCoP63Hrerin
mQYcYEMDrH18t5nf5d1eSXy+WoK3Vu6IA+/2K0k5eZiUo6CYAa8K4rI/oigKCsHb
b7fhLcBCmls0SukrwoFAnn2uo//ojbwx3nFRW4MaL2KKS7qH/VrH/VE4iIMOmchv
f8PH9SYDNwHvMFMAPyzgM1wjuJqbby1JMr0rzA7bElMTB+XLfRi38V9N3vWYRTub
JCTDiZRqWpTuH0/Ukjk/zkX6E1PDUvHLTNsb3kvlDx5nVX+fPLo3xIvuSgYa81al
PjXiJ+d2OYD5Eo92QeHpDPDliIxAepoDBo11bR1KM1NoSX+0DkpzpQdzlt3M8tdH
UzaNXlIPsjuQdLu1Mc95wC5vkQo3Q8k2NTBSwTvY2xCOS3m2M8uwRZEb1RvgusE8
u+O/u2UH/LhtOVk3TPFxi0kMBujL45KC2KAGteiA5Nh325Tyv/8Q7vm7+N6KvoPd
XtEe+by065OBOshVmDSlKQ2OxlB5eYx5dVCFH7C31cvOXQ0BKiDuG/TQutvmo7hF
HT/TeCeL42c9fpud8uLrGV7ZDsLptjwy9av1AGff2AlXMgVMpeebHRdn8yk+nn+E
k1B2lkWucPOgbWjG6ihxxTrlCXfuVMmMJVUDTym/vn1J/HOKhHA5jIGnRNOtroYN
mbNW5zEo+dfy97PTMWQs8oldOmQhCQXUAvRzVbL1ZQ90Mh/gaQzrhExfXE2T+XoF
AcquVJb3XKsO0gE7Z3QyE8uZJxdKBLkSbI/lBhw6/O455Gb5uxmqdrB45V3gVUR2
vi6RLhmyX1AJTncRpiwjkupkugNEWL5SXOkOw07zGm/x4uLMSwvPmJn84cGOI9+H
CKLX3NFZ0l6vH3S7l1PjluwHx7Z37h1OBmkab0UdTbFuAb0ysTnP7l+az3kgeAZ9
B5lSE3TaLTpo2Hruccp864a8xU0TEGiOB262jjg9A8+qBmNWG6dcjQrMCqa8DgiI
3SeieijjLAMqjshN1UmRSnxp6Yi/Ap44eUHhrSiKoTjtp6qwyvWOvcntHxTRFr0t
zy6BfhG4N3xqJkVdR/mezcMFr+ZBUjAJ9zqfnCZQXlGuSh0gcKrcmA9Wqjcc68qW
wYON1IdqlE2KIjWt8aSocGzCQ+bsDEe3EOTv77QNpy3r3mCePS3r20COqmi2ba3N
XaYxyan9NCZcbsjM9qkya6p/o6VHgwG3/vzXwjFVKGWx+MnXML6QX0cYRHyWGb8c
eoy4cW2LHq6fuDJnHOoHa6r4VsLiyxYNZxGAuPoC0u8ORmT39hggmNTEonZSqbsg
MUxno3EAg5CFENcZn8HISYXaGpwZmJF8y0gB5wzMSX0hQ52l8FuEoiMGd0/uq6Tn
x/YmIxzlhXdZMzxrd//hFuuoMnRYlKrXqvbF32jiJwfEFHs1YGVtGNpY7RtTXtEm
G0y62kPy6tRY8YdQlnE9BPVmVqwlSXaEpqopSI/nf9JitjmaucBWO5yupHsjo8G1
GmUCW7NEeKxdignYQRUgA/UPjds98NZFd3dmeKnUQmvrVWkO9KYSXvL1FosHs7Wc
E31ezi3OCU/eTILNtqVQqGEnK6vtcFVd0pIupIGVFk/JRmMPZpb8NIErso8ofdKi
begMLe3ZQ/XwXK2pBngwlF6PmA7bsRllMr1Nguu0yHvvSvLRlAVRNUjmawfx3B2s
1VEpNjwGCNNlHfU3A3CA3YMa/xcA8wubXIT6tdPcfuPqrxoay8JJ9ZOYtIfd04W+
g4wSql1G8ay5o15rc2XJtsH6L5jJDA42wDyJQyOd41zI2KEdmH6GiMi33Cln533L
8yAWE5luXovUb31+7cGKzXBcM54sF9ZKPpCmuVhT5MTSaM0FsiAY1aawRbQiMSza
iqBGKB2H3i75QIxPLZe5GlivlX/Cds59HtSZCf5QunJuQK9mW85Lm9BXPtz1905+
PzkyqRVn3ajBSHi8ctWKGpJ0qeFPRttwm1ccayj9ixLMnLs4pTa1/BUPHylc0lXi
Hz6U1aSy0pqbYoh/PvJJNneidWiyLKpYNd4rAPn+jqoOLBBY3+w8wBXiP7mpCbDu
yrQH0Ipto0aLR0MgM4KBM6Rz2jPZOVcVnikR/IgE4Ij9VKNajqoi3xpBt80a2Np/
hHY0wIXGMz/yYdHaL15kPbTd0pOqNM7JobUhSiy2FNZlDvrX5RQnyo5kWBXp85DX
26PFl4oo1vWFKQxTNTg6BODFBjm6aPARQP2Q1YawWt/wIgVlsvqeNaPf8oq5LKCL
YDS/S+GhTM+juEgjs+jiTPLC2ZIU+FmX5ga4GKhLhTTMs1fjVc2D1MYjGfQDNE6o
6ReTnrgHhetA24ifyw7AmT1G12DLRYqfOKtSJ6oTlJb+3cmPbxHl8Uk51s2jsr9A
OLRzUqbstTqOhMjRgPFYyBeaGKrWqHV/oOEPhh0+5PM1T5KsIELuW8Hr3W8KdGaw
3b49x6yUAGDiV6ecqVVZRwNKVIjpEE88t6xv4fgVeWshu+L4mVRLhAUiXNkOek8S
mZvmeVCozGJsi1CJzDjSXXLcJA8OY3HVRtsZOzVAV8/QNqE8qwqvt97IdxpbSVeB
VPyjFr4rbJMFiHclgFoJcaAZLECz2TdKN3pof2YOBbrzKm9NcmNTkJFx7zri8hu2
kkrRQPNWaw5nc8iHt/otwE8ljo2X0LCbBvEvnT9m8moYVRZO97i1Gz7FtVDPksZp
cjyVcvqkJvf/BzchwEnACtVcz1EW9ODLIhmOAIWbjruIg49qNBETYlBUbJ+D/lYS
gXqy+zap0JowhmzDtjTkp85x/+kDtL7mx5nXWq3QsA1JSkfZMDA9o7sFl/DUEYgN
inUEcUjN5L553ab5QsBiBT7hcHWgtfnjiU1vi4f3JVOIhm7iWO8pnrAPbm/08I9R
tV+iPMfNWvK3Wvrqe5g3FYdC7+qoy06U5oe2caD0SVq6vnPu9gIOAzpVX+BU/Pc+
glHyCRsDXZNLvNMNQOzpkhwLe+934y79/JLjyEIVnnfW0tIXrwmHO5dq4NWvS+QJ
V576zgGlNAQWfyvm9+H9txRX4c3RklmVon+5wvApBQ86rpWEXcCg8bTbG5jiSn4h
OG21PDuTQ5XvZtc7DPR2lisMUo9AOOsuvFkfGOBN+8H/XFU9uVrWSOXuk8JPq3+m
1ulUqeV8cH/1za647ffBQr2DzasuasumQNJcr2DIsikv8+XB9Do1AylEnqPY0fEz
qcu+9KGDsFWhMZI/GcJCXMBAf9Lc0/TNeclcEmH++MhvYyeJ9mNF0tmIt2xeDExZ
1l3tz/Ml7T7SA5EWz6xGegrC0p76VLlje25RipYN+uYM4NT/XRyYDAr1PXNoxDeO
Q5JqzeTOIDzUj8STRYDdKAaU5AH0w7IWS/pWX2BiPaf/r2IOvu7lfbCN6m9fPdJt
QboAKIDfAPbdiSRQ1mDYYIrd/jimo6tqOstW+Pv5K4S/YK4STX60lQDU9DSox3OL
N0khmh/sl4+TLsa7/JJhcibWSHQ0DJgjZp0BtemTjSLbVjFMHnEhBE0FaPBpkzPB
b8mWki7YzmfNUk/YMNsCZIAPv0qNESZa8I8GyCKV48QUvJ4vCv4YA3/lnUFOVBOz
FgmGE3csfYCMT/haXn9PKefZ0kaPxtxFd6WEBa+BwiXMI/l1DbGMFW3MEzW5UWl4
48TIkFRSu2iKLwSp4u2nAsFDt++zrA5te2+0yvfTw5tk87QsZnAQRNyrOgzfO8tw
x/LqnwLB2o8XZkSaEUStru24cgrJkbwjpAJS15nPsUyWNB0vHIdwF0+tEdesUJmf
d8fDyoJbFxnc2ZDwpznRY9kTfDfLWl+3BuxTaYTiBeaZ2elXntTiDy3FOVyJZ/S7
3qpxH31Opr4bLxiUK/xI5nIG3GjgTE+Yz1/Xxc9TFdZhILoGozaI7mwj2qPBbtvd
wNQOfnzijMhOD1aLc4HZCaOJB8OwIVFpH09UsuN196FkMmEkcmLYcuLycWlCPeGa
M4TnqEQscfwQBOqQniKpcEwG+pKURqeFHWOmLZAsBMIVaJxj2+lgAR0WIj1RXWVY
Rlm9x++letL/54qG+gxq7uKLbNRwkj9mHWusmjJjq1jIWG3MD13dTo4gda6tdWrz
iAXD2QKd1w5LP3d19GqPwzLZp6aPsHyjmQ9SFZgLT3LQqR8OX2d01c71PzySIQeq
lZpjAuVsIgA5jK6bOfdfNtgPLuwvTf9gGixtKoMThDlk4Bwvo3q4HSiiyASNSGh/
g52nOVwiKiHo5KAiCRiE58sN40MjPAEaKP/yYjvjwxYAac8iFf2V3ttVQ4X9LLk/
pv95ib8Zr46B3izlfCq60jg8Mq/3urI2q5ZlBwGmg82LpdoIYn0rLaNSnZo2XXRP
dR7laIDIWTbkF4f3/Xpg6FKaqAWyPCS8WvMN2CofCJxm3dCWABJy/ltwAPdBxM5e
avYnmDehoZ8qG8n/bgQ9jtoJegx+18/zqt++xVsA2mt7CFfHwYlBvVREtZ1vQVoc
YA4+aP5b1gCFvGJ7KoZDzhnlHrvWABPWHFwELdSRKcCplQCYfdbwA7dY/dAT+IUR
TBC55cfykABgSgcJe5ZQ9tg8C5MsCSVLQ3kbY8TCLbR1Rh6NmkkD5PHCKGDE/Vk7
bQbrQOZypyuBwlFewbh4yi+MNPX0KEos4L7XfNrJj5+myZeT3/95H5hf+oL863Eh
8IHMEYMqY1tPMXN72Lgzl/VXzlY3gkBo5DmcEyqF94g+zxlLstIIisJA/HmiQ1mV
QG48xUgwqbIh0dTQzS0DxrFNLy7kcVj7KGQTKcLVs9IJAHQ4sP4ZCt0wk8ZtVp1h
YuhV03hxdD0GZIIufOxDJDvbhpdUzZPOAeyFwnj+ePecnIGaknVMq8a0zNb4U/8L
s84jkFxCfu/UCrx33IlQmylpkQuWuklMsBpr1O1v+SyjxC3HaJdi2qTyEwmEj8rh
Ce7q2eAw+6l8wc1Zu8mglro1a6BBHKOoXWolZzzXRwB3+a5Xj6yUhnYzkTLiKfch
nxIsi3Cr6VGjVJm+JfYpemQ1maEIVss4ppBfaNehbW3ANUvq8f9bouXT+ZBIDFLa
q8ZF1zdgblvn1LRtKm1vuDOHmFTQWmFaeDxaKT5Q+gZ3TKw1WNZHggsJYTrbGNRA
7R1ET42wo38TbUD6mIus24ze3KFT2IbW2xVmrWpa43jyC34tN2GhQAY6wEmm+Bsc
zkaRFpaMlTjQn58X9pMP+7fj/mx00g5bgkBDV7ALCUnU0qR3ihhn+3o1EkQ+788h
/M5z7pClNkYB14Y0NSt6MBH9vQ766184dkTixApB4xbYHfWE4adzVC1qJ+R8AWDy
ut/yIjeKsSlRjqJnrDGM8uPIzg6QKEO3b4/5EZqhy0c3CtQrMg97ohE7etIk1QCP
XpHryv+TVg4dno75Nvii2OL1knnVs3MP0Vdf0jh9+SH3+MGozbTkTVyEdYgMjSwz
s5UKxlPG3HrjkJNSS5Gdo3Q90HSiJKDr2ornkYBIC8K/aZVOvU8cN3hI2MBX9ZMx
9CWHMVxcp/se1eed/5sTWrOewzGSigrPApO+7Y6Q0byANPuOsOJffaaAxee0gGhD
dS4HUXsfmwHqS9GA5DbVJaJNBEGgIerAiun1qcF46ce2I82m3+qNld9R8AIg+eGf
tk6wTqGvUjE9GVWZ7Thkc61RogtUFqdtg0IH47f/qyyHlw5yM3FJ8ZVTf7Xx5Uym
E+DXYcHDfX6MeNC2zOvkFVWtS942J0VTbVw7A/DXB9kstAd0cR9vAF8Vw0/9etmy
Imxm8lJoRIx0Z3oihvCgZ/EHxyYSrpZFW/ajG1yujOJPOw2A+Zo5Z/WpzH2WzV/C
wK7AL6fZ8L+NdNPoB7SRR9Lkgm3oDoT+UbLVyFm1UJQzlXGi6Nv8rIYtoBcHNkYw
rqNmAezQxyEzvQAnMT6AThZ1IWE1eBganwljelU3XCHo4uoXXpZCh17U+toAKo77
5OADMDHghsEvQxkac1wOGKyg59fLy7sT9PqbngVERY1zwSxd9IJ9GQy3iiQOrAAE
w9Kfd5SdwWmv5roY2VNZfeEbQ2fFYsPP+uj5esXAPIortMliaJysL4gNORgZOMxC
/vHuoWO+XafrQHHjUq8KVBQKJlJIQdA6gTkLyIFeYhBVReJHNNUlwn/xzgA3Q3uA
ngL/AYexuo1K4w29P1laBNyAu5KXocYZqTJCo6vAg2vgS21Lu361xcK1J8WTXcmu
pI32Zi1hv6/WufoOIbmXSeIM7Fb5RW2ybYU0VnDCQ74k8fkSjzDcjcvFGUdmZCRt
lTc+iT0doogD7RyfpKEyn4kOFMrFo+7hnGUBszBkoQ0kNvQ9UJZL6zxY/XbYOV5w
g5svsJUVz5HWZzgjWi8a1Ct+1JjpeQXMaTsoDzEFVbXXN62D5IWpodpiOPONOs/8
uVDZEsDjp61fT/lGTWyKNS4D0wnaO5gWE/L399TI/501S2yh6BcjQG/4XeeUawzD
KPEOe+8UbVyY2WoZ6vpv6AtGAf77EvqbGP9fnW5lTXEnelnJK24vnyF7XqPb4s5O
xmU8W3iui+Xapyx+Puy7DtrsMeL/O9w1U2e07AwYHHDhySPqb7ZR0pLwDz6Isv55
EL7piW5yte7U1IIrBerHQBnKANaSiFYkTiZD61pFzSvXiYrEf1ZY/3P1vIPQGzks
v3ajGb7W4CrIadIIdI8Zq42KR2/vlOM3iA6Jgq5RjFqZyplEdHer/LxgNGwL4c2N
vIJfSueT4gFSJg05p/OoqSALM9z6WlqPxJqFVfWkwJm0St+uClzirVgLfg0ctNi5
I6mFytKGdxR4sQysnDZg9xTvFa2SdYd2/eAr1Tf4cl2Izis5LMJn7pg0PzOSyRzm
QNdNUGe4wXmILlk74a6V1gCX1az0oVXC2qto+TsMkYaAX6MuLAI5LWg/vAHLE2Lb
h63IyfczKXs1IJ3C9VOjTfoxcpoyHAZEg36TDsl6PcW5vQLpRQetKbyY0vKi7mdV
67Gx36AJEdZoGT7R87UszmwbZjDgUvdJ6w3iksCcQ193QzuHbmWuhw6kPvnCakZU
F4xCR3yolgDRWCm6SIfVVf3Nit1GzOPjJB1M2Bd7ZygNoZPqA6X+hwzWSJmeV3uJ
/c1g6gWK1NGEPtQ3sJaU1cAE8LKCp1+Br7fxQ3zwnRxgUefck1DBq0ZwPy4H2JmP
XNJtxkpe8jk5XMQyQDJhSeT7Mpm1gmMpBAtkiEbPAkdtWkzdzH8wERbsOF5m6CZw
KgpHRO/f398zlMjAqTWKy30MPFpnwQDtva+oQ9HaO6mGvjPuZWnMajEsWMjYgHB2
IVXZvFgOn8U9QXXISqjl2LLgW2NOEaKYeYK5TXKbvXMs9iEQq+vufkaP9zAnrsp7
erdmjrUWbvaqgU6FzzFjV76jgGkSVRdj3Svg/QX7irXuc2Mcb8TkM3LhAL66zxsM
zpPiPszeOueUCjJGfU66Gp0O2GFgey+Y60AoJw84EHxVO6AGQl3KOmjZqkm7/3Wj
bZGn3kCwBzrBWLZEOpjFzLWeaQrJCtHKi5xsN2t703/yNPjb3uMrYyGEkD35GSE7
8HO1I64oGqoS7MWalF6LHDLOBy5/sL1xqNwBXXeQcOz5kytOhr0ZLMRxa3vZviOT
Gyy/A9shamjpdgD0q/TjO+ok+MM6+ZCxCTEm1LAEmnIVYsGUnLXM8xgyLNGO1EvT
hQ0GXvRYbxgyks5pRUCby1/ymix1Vjom+rBzj/Xdr6FkJ8KL0aNYqCA7CLtriaxh
9gMMVA+JEoyX1fRgelBC3/gkuCvV5BUj6YwtwilFshnYy0+5Z+owNwddWZB/hO/t
pEKtG4IqzLIcWZlvpc3tqY07St8+EG8t3MNGgNkV6REZWTwDwxL1JIwKD4BIs4Ab
ROKYVke55A1kIsKRQvQbhp1ZzevAcAhXKvk6ER0rwIhyIL1aRmWp0fmjUEhwcpjA
pjDo8GfGk4B6ham17yyBeXB90aRohf1qCf5Y8aYmQFer156E48tRng1h2F40ZvHV
qG/1w4RiWHSqK4hW9874Mmuef+zJUPaAZ6bZ+9HGYa1k9LjP0mzkwQMTTbbkS3ce
wPIaz18HQNEhOZqWyFhGtQwtLk5xRXKFGqHMgBx6aF6irBxjwJ1R4LqE486XkDoe
nu7oiLvpj9IIsVqOTw6w+1WBZDLUC1elWoTDqoX32XxRqY2FA2JcN0RHdmm42im0
1VShyY8N3F5+HNuwY2L94h7k47Qrge0NTob9xn6sTDAJZik9G7inyb7IVe589Qlu
tr/8beFPIZlCj56/4jcBh4szN7kS4tiW8D3TKZlgA2WFJqtAfyzu+WTn7Emdhj4I
z0GC4+uL+wpAs1LLeMvp//CB2YYXdiF/SmZz9HC92ueWS8qhxTogVVXmindnubRi
I30IDazijhPxdpNZHAK9PKdVqL9Q//FVKs2lH3vpDXU0GLE44oUVv6B8a+wne/w1
BQ8JyrKWwSN/cXI1DZ/HLvUMM9PGycUk1KCFBLD9LWt6KqqX9I1fQF9id0ZVpbXc
LD3Lyd0iuc/24rXhnQ9+XI5sXitnbqZyRe/l+dp4p1OLKTlI4AjhdoDcAekAhbtp
jg7RRfmRVjM4fpF+GQPnkbTFkx73bC0gXxsBNBVlRzs8slIXfY5ELIi1P3eOZtMO
lIPzxb2A5r5NudBS0EqekMunHBc366nB/qUL4YEfSlO10MmEeTi5Zh8bFnNTRxKJ
3/vDj2QXfqAws56nmU+k6osFXrzsxDCNXFsoJ6AmzE58I2XOl6L4I93v/C/Sn0hG
MDkAlc5Nim7qS4E2+r3wsfn862/iu+NecXOkaQ4vJom96lNFEJHEgnpucjJ3v20A
ZcFeDcWyg4rglohgyrVMZIWBB+rrynHg+CrrP+F0NiEnjpKn5CdEzE5690ePLeqa
1RE2kREJV1peXQdz14KvJKlIopvyjNuGkWkvM7RPvUnqBl6H9V7JKuda+t+X27+/
UiFbVszicW7RcDTT15Dhx2w+QW7kkagItMyeJNKEAF9YnjidgT+2guH56SWC0UZs
alABuL3i10Fm+/s4tvnY0uf4WdIxOKrG9NmB/zvUh9mOlZQ6j66K0FVDdoFbPtmY
C/xKLRfIVk7Mnn1spfb78q6FkLYfZeIuI870hBaVefw/P3CYA5GYdaxe00MgCQiZ
PekG1Y79FlewKgUVzI1Ug42aGdYWmKhyrdZJ7vkg+93gMYKbx6n7Q8qTsEU7I0kg
rx6QBCwuPQCyFHsNKzFsZHPNABvMre/03UzZUcoI9dv6Q1gzgCvW1CYj3RLXD36a
/MxgUlFgYwvx0InbhJK/tALGNhjgrRsCsPHgN9vPPO78+56j+MopELpavIpznGP7
qRTTIicW6bPJt9NEC8FUq057LTTwiELAbZ0M2djrcxioJXl5YsALxJsa7z9hXIFl
HnGVEyrvCf/m/7xQWe+PDVxaHS7umpY8eBNYd4JitartBWBReqCFLAjXgLjFZiTC
7Kqz2F95Q+wjUEPzLepTETiJIibpFH19Rlk93zvAM2B5+QpDWlc/ltEORqhb/znE
A7OmNqn1l8HXPAEu41NLR9bdO2EM6uOVRosLgokAoEYuHdeq6MiCHXQD1Z5x+vyS
XnQtfp+bpXryARzPdLE/Cj+hnpvbqwuhvamuMSNLsw5F4XZNuBBk8Uovqfs14DL+
RoJtBMv+37ZpsXhlNpici2/UCdA3aNT5Vid6bSWdxUeuArlE90j4HlOjxMxbPJTr
Cgwgk8y8tmzR+fuuymftw58RIzAg/VLdhJI0zWSP84DRgEgByRI+LPzElrapi/EQ
/UH3PpyzVC2wKmL5dpp8FCHfw3nCK6X2P0qV5LD2mczTWKPzz1VQd50ZgBWNRI9N
K7QnzW7h3HoGE7drmE89sDM80sR2EfdcK+JWCZktqxdoAPoMsJDdcK9kgKSfRr9u
5veq4s0arwFGMH5/pB5XpeMP2mPmcOshrNufU8i9H08hJu4q0eWGVzbMXpclY/Wf
AGdIg/RyA+mJRwG3WdlidYDoKJgFRPTd0S/TLnOqyAjFZYgIqfPYU9MdmjpvGAAr
j8aYxkZ4FaG9JXoj4D1fjN7MUapdKhUFRjUwxi6kALTXTV9sIh804aF1jj59enP5
X5NK/5JvaK1ylNPg5hLCw8tG0uL4nVA4wFUSQvr7NeY9ieHjfv0fCFve2ABcTgnF
lNTiB5Z6VUiZWLO+q/Fxbd/CF7bQaQPg/ksdKpGpSLYPqkEOXJyLKMVrE9abo+9s
leyFPP5Zoj7Te51Z71dexSjaREpNh+sKPzJa9JraL4b62Q1zLUt32ruo10E5Tglb
SdmH3LIvdGzzbSIMVSX0+8/PcCAIepqB1sR/fEC0hdHVuLLWZSdExe9G/IzgIUlJ
VP4domuTesynCrkrR1od/4zyuYjZOACsdBp93McV/mxmGAS5ZWfUJC/C2x+IG1Zx
Esmt05JOycvgPatAAyLbbrwMI1aPJG/+32PXZUzsWmuhnQxit/Ra3FZd9ZrjubIY
ZziVa0JHgft8DeWGCesFHfJzd/Tn/V4XZw3VDPWRGiNq4bIXsht7grQiw75vCMYq
IbJBpPdDRhjEhnIxq+3/P5YZfTieUtAgllDi09tDzn2d5WLSAiMTlLDqUuTiRfUy
ufwU4njhaE/TAvjE1Mutzs3PQBnWh7UmEmmazrsfVpYb5GxVEGJ2Z5TlPoKtagFI
cfMJW7CAqf0RgtfztOdL4x5Obs2ppQkaiJYhLGr2vVIGE8y2gPrQEbystPX2l/He
68qr1ktPQ/fkRpb3mSDxHcc3ds+X9M24OTNSuhyPeDUWRtAmMeNirTTr/pMxPejx
oXFvfwQyoEV8R91/IKZO4odW+UcRyyEDi6UsFPb2c6xE+vJMa//Fn2HGu/B+Ec+b
xR0IoT1dnSzujDDiXXGj4fNgT6EQ+R8Fp5T0JbU/203IjdW34k4oM6qIn5RG7qPT
6ZYJDe4nuPSRYd7ChI6h5BmOx28ucncMkokGB64hpYZaK/iFfbaH3BHN++jXZOfu
1Ri55s+mh1ylPzyBkFJOSIYd1o/oBIYIy0yoTO3e7XBFwKgVmaoc4EPzGMEEV0Pf
nARAj5U24e01nuGWSKdXBkVQCyc0hh2KhjFxi7MyF0opnpXBgKCl/slQ16PkH/a7
BAdEsv8oDfL4l3qPnZ9gWCe+klF+TWxrzO6QIgWXVcCHfjYxBzPG3ky/Qme3/Ggf
aGUroudUbflhaXYth6ULXtGoZD5HR8ZslRUE5aGK+98mKUC+o0DtHmXjwo42k7/T
+VVJV4Pe262wRHOS/rcsYtLbPm62wgraovjVWw4c/4ybDvwZaiOe+Fw7LiIbsXVK
QZ8zNpXRgyMeKIjAq945rYznvcoFyoqjIa3rDCeyk9WsH6RielHky5fbz6G/tJ8y
65fEAA6o2KDnzKj4JN0iPcpAddqLTwzznCnTTlqwIKrs6EQyHlwOMxuefscJAdbM
KBZ5gCOlUAouZdWnaP1KUfdh33BaOWN4YNiVmvhB2/eFQSHkUedMFhMfMOVAZGO5
gZDKZor4W5+IGlUkSGXzh7TmL7d06CeFN7iK0b+qLL5LLeQ0gh8d8ONCL3NiIIXo
EDD9HVX7umyB7yrKZo729MVtGUgqYh1JT3+l46Z+EWwMCImQ7vSvH3ohYeBQvaF7
K0cHpIF7lOBjy22UeOFg5F1oVHfYfH3Y13awA4gBadKfWZuccR1FMjdNTLPU4L9l
KsFvJWiUGC98HMYkK7IlPuf1ydaazWEbjwAT3T/p5Zd1N2N20ibfvy21ZIGB5FbF
lJEHUVcOhmDb1TUY9lySWJq4cnURZZhmpyVvJ8LRKXnMh+b1uIkrpAdqWAMy4FEu
u5vljyPYZ35/a4dV5v8lMN98G8jYgwnaPx2/HPPgUIVdX3W45iHSaZDubRvcZA9f
P8qtebPj0cDrhEwvuboooYdUyBacPiQsPTTLUofjM9qh3FBX8RnAJI4OXVuDtKEB
CE1FPKGuHdXsyRX4eHg5QVsiOmb4R1MR09crwulQF1+uZzhf7larsNFQN8OutgS1
tgrvjoItHqSxndYHtTro54YjrdtWkx3dRN3zgQTXis/HzzwxmmpWOvo72rbrpvuz
UkwuI+oVETOKgVUWQlN0PCRrYhhx4f18M2aY6lVp+1c0qRvWofU96My7kT/L5qZb
AmZAP96dhQZsFwEdHpUeSv1ku3UfPAI8kDqiyWXgmhHD8VPEqPxspFGJOPL8A8cW
nh6f+dVJCrLougRwLNWQ3Tf7xYNjOGDm9MwjgbVyneSlzR2g742g3zl6JEEi6ePY
R74BclKTT3EKjfuTb5KNF8tIZe1y0FAHmG3dT8ftaRPpZ7hxCGk19dBDYlWkvwfb
EYEWMtIoLFYWWb7F6FomvWO+tkCRsaC91K7S9iA7XX/zrFUo/cyUJV2YS4sLcCpa
p4hPSiOD2Yhc65BnofupJe/R1Uwxbqcjw9VLbjW9iulM1wuB/UZlhQ3ATMfSkrfY
G/Ax3plYs+/KJl7NS87EKL2LxAraiLcc9276XpQFupZySLg8z9bgeidMDnCaybxw
sdMCwodG18wKpCF2ofkCygXyAZVhgarLrvpenVVacKXflwzLRHdzhvQboU10GoAT
EsoGSjCiquF0JrLNpRB/s+X3dfdAAA2NXx4iEdUNmQkFFpL49qC4/LLxHFzQhY21
W8QvRKtNqqHzrr6ZWSGO1Jfp4H9riLqoW1MFM5QBobCFJzAWOfX2sSBHjfBCUC7F
+PctJEHtNHuUMWI780a/H2FSkzZIovkwuNkr7xTbl5pZ872Hr6dDReffaDL8jqL7
yse+WBfml10L6WffPSE/sqZWPa1atA9pw4+BgQxtS4TbYc+uKqyEQ9s0QVIXTXo9
0OLgwX042iiD7xK4C0FEvecjO2TZdqrJddbSAUeUkAQvZHoG9ii7LH4SWMAs1K8R
rc3Qn4rKQrcuygtEVtbpfFFJkIPc5PASgyKaRs6Fv+Ziy6OnpXbEsFaQxj66MaFK
du+FyGyDRXn1yRvhCqQbxPATRpQJEqDZCcGJvSFPZrH7FcQvfdJkfGoF9JAiEDF0
DzNfVscLYOUVnZxQ/97iS5nZk3ypvpGuaifu8iroOaDilQp1ZT3i73vpH6eOpmO0
+fAldC5+k/wu/X/5JxbCOGxaBS0jy6cNSDJUQayKgY/nvBaa4CmyyzmmqmGCXJLr
9sNNL/n+tWUfb/ss2piSz+dSX+Cqsvmw30GboFNw9haQKwRxvz2USUVkFTYNb5BM
uXlV3UdluMs3VJh2Uyf1+FSbhqvR5ampTkNY+R1RxlTADRj9Or1pWnVwQ6ADs4aD
t2lc5spcRF36eFQscqLQtlC2u5IJ5PezOTsiisNdXUZZpUrof5pxAmrxL0RNNEEI
EMt6lq4GJX+gZK3HjxYa/BKpSX6V5kIU5TKoc3rZxXnCJRxqksbQPBhonFMb1TX8
1EECthg6DXjhEEHNGvhnRpyq0rq0FhJblGoYjCbGyfDuDutT54eJXZiESODu+k49
IIaeu/MGFdYH9EbNNBDYR6wJ+lNy4D2KgNg4ZDwDyfiay4vfYqWUoRnkc1N2lu6b
p+LLJVMx4d9oWtvGG3K00eu+2hRuVEgPzX0PoXgg8Fdyo/N4ZYR6fHDSaOjk5VNa
aLW28L1J2zvDXUzv/6YckHKiDWZNj/oNjhXvl4BSTMBdgz2YXcTEBzK2TNabkexb
HTCwVDV7m0/3urfyINsUx4T74OfrEAyrxZA1UEKYz6ksJP/SdwxGRyAXcaGV1R5t
TIaaiQ5fyxee1/bCzbrGXQ7rH4HQcTMTClWmKwOPrSdVSSuZTHBEIqOhgpca0Vl2
1L4roRobSQCygl75rOGEzsgYpWOK+rjtycMLbFNqmr1wzTzkQWlH7jrRyWotNvOu
vF4GLp9wZ5cg0W5AEVJyoF3wTiWkj29yKBqppXrvbtBJNcVw8zalDj0RGhalpDv9
GXOd7clYhEKuVIwBCGvDXFvm+MMMgidMMfsCfuQ4Jbyb9GedgylsXsbUNtZPuc6h
IYf27lFqd8w6lo5qM1LARIfhFIC5qNozxmp/K4N+M7rKHVR/RNEcnNMBN3EeCND0
tAzmOe4k1hQRdgCdCrNr7sNwNzPdixWz7QQcH5cV1EIGZDBOSz3qFgsNC9nPjNSc
3Wex6qbmJ+trCBITGdQnYIieltBPbs418YxNNmk/tYRerRRV1HZBQ2XdBgYN6LTO
MQnnHO8+KYFT8wh1MJ4NvjpC24tVS0El1CMRmxDt3Zs8B4NPGucbPLhrOYYW7OzP
jH342dSO+zNzlRnE5++u9qtc8u08wToJ8H7B9mikWWd/pcL6rq7VBO64a60obpgW
GpLuUDs1GqGHL3Cx+3HcXG8yMx7gIqVeYb0Add6/7Yjqa3qG0uSnniruvnQ8aFbJ
jCwsn3QaaUN8MGnpdCAefzOuf9lXELx1UrmSulbkXHZoXSP7L76YDpYkIg8xncCt
liqzaoT9xYpWH0OUcrANqYAVL9sCCt3vi7o0WDSXTGcgkAmzu2wPRao6xRrUcAfQ
G+T5zrNm8Te8mdE44Lmfe9heVmgv2LTPxYyf2HYPS0v9R95djfifyEKsyXY8g7aW
6cvZLXMJ5CIkMPkWZ7MfgrS3IaX0K+wZk9bXqdB9mYS0oLWUTjv/GflYk/DNPL5Y
rteLOkyChcasMWYCm3WKb+DKQSxFoYEFeCNgSv4y9riLuhMgtEzKEQ04u6Q6egCJ
KZfun2Ub5TfqdBG66bB+A/uk6cjcvvhxI9O+BdmTF9zd4DqENQbsqix+NDnFBzbs
DuuJH+KbJ8+DeBaA4ElMVBczUv8t9MB0MjMBJ/8Z6EQ1sUOt7gTBCKgT4/SqzBTD
0sAIr1TK+8SPeMEJrIsXbnI7PPLvJF7qOssuI+sE+xJhmqbenYeZGVZVkN4Vmn1F
oq8OGQgv6WNBxLJ8zOxucdWatW4XwNbnO3Q+/ulMeBtL0KIA9FYWq0swurUWWqkh
f+gBJnfb07gh4QvSrag8LfJVOpZsBdEfdpTiviabbvQbdfGW3EzYo7a9qisa5p2Q
DNp7uZV8f8Le2ItEKK3BGmKLN7h596lX9FxUpYTYaVTIZeE9Xa1/Z1qyIgncwMHb
mWE4Pb5KdKAkOriVX8RIANF4xUN7iS1kIpZUItu0fWIh2YxndY2guc8aOsP7b1T5
pVQXd4d7QC4ZFNSIiI7dWDt7fQxBdOWak3SzFpCm8DXX6oyOeg6+7qWIZ/wtntNj
SPnXLeukIVSzdbJzgutcoYXnWBShbU2ZBnrSNfqEiCadQPT95ME8d5RNmnPszQFm
woINpDGZZ/KQI7D3DJQGmUnPKcmRlJs0ObFDktD/mvhgbXJ5wJURFx6DtWe0xMle
Y+j+28HfdT7nE7uJ8vmM8hyXFb40f1bPT7mqZLPVWjrF8UScDjqYwg135yV3tzpZ
8yvFTL6IKiz6z0NSXafsOYDqz9gVaP0qXFfhOSVPFvYOSiey8Au9Z7upzfewaBlW
SZx1SVuUVxXmecYWMOZsGiiMnRNKtlNYxy9vrdddVHrR2l14MKt8hsb7ckqCFhR4
uVPU8tAV3FbBlHyNyosN5FsWwGWIKeuIWteogBufy44mJu2Xx2OWYfn82WYfALWw
MccLfSZTXUu8teOz8a08d8jBAGP56t3gto4kPYZFw/kiDayJwTnwBmmpnyM06nS2
JWCXmqeocHI5wen9S+JIQyWlFB+e2NaOzkNuuwskqP7yE4BI3quT4bV6Na2Ze452
K25JzVPsyq6mXWOcuz3nw3zsfiUsZEF+mgCK4SkYhY1nmewhtOQVMVpPCl6bBulC
XUX8QmAWGgKl+TBTXaxXWlTFdvbtKLLlmBBZSrPbMMXwB++cXx8o3pjjlcBiTMvE
5xj17mPoyV2CcrYmg2Jc4OgTdH5KOoYxOAyacTdJHMpOZAuXXGyKGN4HuzzGjeIF
87VfnMjoEmcrpNuyFE/TWKMqbypPobPEriBPkr1VoOEzY4u8mxc3abhdLblSlozV
s7A19YzS6u1A0o9jEXOV4nW7LQCL/AAuZWi+nVW7pMCHK4A6nnyMkgRKV27CjwBG
B3VyaUb5REycr3/Il0kh9ilm8N1AgI8gOWk03T+X6eVloICQII2zKcjFPf3UWxU8
SZ6MX2og7CGEzALuSKhNHvhz35/jDXOEpdYrW2Nq7HJjPlkcuOAaBe6EWNtFDZ4s
UimWqsCG3C5bEv0oADliqbYfp6BieJcKQyAtl0iPZdsE0hZc8Tm2F2jRhuiW7AlZ
+8CJR06fzsdSuYHWBgQdzMthxxTFoyBQwELmyVHPFt9ribCqWIjbTWPhKEUj4LR4
hVF87M28tLCoDcdGIt7yiiFadRiH+ymYRri+avEzvIAqSXKzWEX6yPM8Hlw5KKLG
h4baJQlQojpNrsYm4UvIT3saSZwYvYRelR3MhNEeWN+JtEiWxLxSmYvHEdBeJk/X
UMnn1chQRukMMa3RAurbdUv1Vb2jVqxwvP22IVFYTvpzfESXIWK8Jvo47ox9KbW4
O1c3mF70rJxAiMLRZqNA6QGypNWT6RGj2++6UYMuKrUQgZu0MzSd2SIqKrv8jIs1
pcN6c6ZbMUVDi+Uf+dnGsg/mZap5vgxT4DRUg2v58TEPpVIdEkkARVj+iXtKhoX1
D3WbegXw3A7hwPxCLoZwCtGdhMseNWJ9swvrxBqrY2hadFh1GqIZVWoJu7JXNz7y
ssG0+YFxH5iG0IoDKXenRrNWcCISCvnOYLBjQDUW6xZLvsWcimLqpxdnZQNG4KXs
3bG7c9pZJed0xs8f6q/8Ft5p7lZgzYWfJJNo95r/xpL+Kldv9GXqRJDW4JW3rk+v
WpCBatYO1oKnBGc/gMHtl/a8fBfIU/MWBSsdgLGLgtljq06uKoHjJijTMFmYmcbZ
mrKGewk5jGZ4lnbFoswp4CI2IgAKfaSPGy59wwawssY64+WjGO4ZXbfn+Ew8LmhY
MbYhAhuukMBwZS24Wq4zmhuk+/pM45jk2BiVOaefdj8sy14ZIsi04H1gqxN/nTAZ
odETgknSDdBZrqK1/XoUu5BEm5YdgUaa1JvmkiPRZR1lhs3kEtKfqnJ6preCG4SD
Sl1rTukTJ0JJXUJcpVi6wrbKCpDHTGSDIp6KiskEWSkOeO2TEHFeCZ1qxpk80v1J
FoHjcWD3D6mzLuIruTRLKDl/7JnOZy4BnjgjdY14D2AAneXgdG1VARbLhewpjT40
A2Xo0lpDK4OSNg+y2Ixt0reDiPAe6ifhWU5SaKAXBLplQwy5eHU1Bmdpv+icyOY2
I5JZVei/nPQatm0XtQvY/Tx6QqouHsMEwvafBL55kjhmHXxmTkgBx2ZB6MKhIhAq
qqiOStNXucxqeIs5uZHkLZvuq4N5gC2hVbtKQJpDKOW4Vby2uy/6T29lVclk9oMB
T6w8LhcFuPUrEoAit1RbAW/a5ntikVdrb9eug48NUL5+gGJqT6H6RFNiP77rbHYc
Xe44TiXxPsg2XoOpN+D99zJ24/DkbFbfjra2puwXYMOGd4JYtDyMh/kbOsfVOjNZ
UlCNnjPPe9e454vejHMU8sfMta8G1U9G7ZfSrmzt0zrShbcQABVYLAbuxhweKq9c
w/MzgfRTVage6Nk1Xtjk0VfEK4WejjCmUGMMWdMf568YhBv+Am3iCiBsw7ojdAAN
Uj4eH/D6EKqzDS6PxNBTT7whM8VjRZh6y22ckOgbMD6M7fDdLhO4ltfjMhL3Ya15
2ljOCozVT42NqV12ImqLiKL24d6kSEg+ewtIy4JIejVtUHTzGkfOV6XOYKYKO2uL
5xT++K2SCFuem9TD/vRm/bccmdWuoW1V1ZUvrlLKKTnJqY8b6q2H9IXne6OsO76U
MfEAq6ftNYVfGKyciKzSBeyC/snxouL6Xhvlf4ay2an7DmVO+jR9i31EofDYGbio
hLMEOPwo5oRiJL7vqTw/iRHqKUQyxSEbBCfj24OPcsTKemwQ3j8g77w4vTRjMjhI
+vC3/TXubK3ijkVqGiJ9rmmnzzpMoPT0veVn0iXFh5UpOAiwoH8+EndeDxX0EjzO
Oa66GX970Tzk0lDs5PFewJb96tVvE6bDdBNT1TF1+XqUswBvU53ih3pH+3TWCoG7
slyuYJ7j0Njnm9RRmfdWZskNXTcSspgUSk5HNofDaeNDneI/yleb/0eB6jpBPKLe
ugCvJDJAEFGUeyKNpg+PKg+oul8R/ZDHuLQoxjXKevQ5wOAyNqinQNViG1OyQ03M
JT1+p0mMZve+HvOyXovXLY6MIUwHTNLVxe585LGsbmBIQczuhVmGDJYmL7zYKpw6
eCS/OTWT3EAfPO5X+XWEnHGYOCmzDDans+7R3407MQLveO6W97aiA3c0ax/Ep3M+
LEDT1LiKSrOI3VUjUU+DJn21HLcSuIz64c6Rhpq7WpjLNI1qDuciFrOlsr3/0oW9
n8KShlr82eJ9VkpQvcc3ArAWR1jPmkDVa3WO4qw+4WKUS2TSfYel65yOVFFTcDUv
Z2yxCwk67iei041QaIfzuGETu24bN6KVTzveGvirFMn9dRWctEaT6TTZIFU3XAc3
EaoN01ZjCZYUwGGsoj2266lroFEK+KdSoJqQnuAiYW1J0BEHhT6njhphK2lPlpMr
Fu70cmyBsWqtWT1+VI1Tbo2chpE5W8Z094mIPgd78vJTb7BK0ZnZN0Ib3XI7oocn
pq5ylOrsHgxgLwGXU16knL7UMRAtCVEay3JyLkPmFbFjwmwOvTgCn1HDyZODVhSu
qUcVoTgSXYTHDUQ9CDV0FxwgcpOTnicZQZiInwX616VV2usUgZoaMH4nxWp9RnuR
ZZYnaOqwBgkiNFxTK8RwGnXx+pt9zo7bgY2tnjXU4mjqvIVziXSLh46PRR4up7bA
QsRB+yVTy/IrGn9XmJ71ctXKDSi20Q8doRp4h5TE1MiLgCxUDT96gY6hPIFuZw+/
LpxiZ3X1nK0y1Gv95hOwxG60gPDV5rmSdbU+PtZTucdMlHx3EOLxSbXaZINHz/EO
QYGrRue63So7nzrs90YpDTtnZ4G7oX0UFMKCClcw0xxWmJBNK3WTNFHljP0DcKOI
sS/aiCDx1+RyuMdXj9OhOWaWneONSz6kilhMg5KkpG11uYNIqjFBpmZ1iIc4iKR+
r0VkVA9LZ5eTpm+bQsk6WIj2s9WOqiCyaUZIr6tDjmksEloZotG0ZQaexcn0v5kd
gPKFr8qUDqWt6XaZ7XuCLs8E42hiPN268N7VmIM+fNFAzEwsj5g15qz9/Wqs6g+P
h69E2AJnu05cykTExBLX872sAYPVrwTT4S3K3d0fFdn98zAJir2fZKxoMCquQ1zo
7rYc/LNo52rrg21TVK+Mq+pQqRtcFX9kch1R4ZAsYP5V/KDaYQI7ecK+pMB5zxao
JQyaXwO2w/9m9D6QOgXUcLXNAli0sPsWgdoBIz1HOENmsqMtO0CWdfL3gHBwst+4
ylP+v+I7UDhBfUFzKsIPbMkX+RpChJiY0nSV7nuYlp25nJJ48f78fl0Ac0N+pSu7
4DqpAzxZgxnMD+KjTQPj3c8GrVFdHITHwtlHuT54Fc2J9NYbyMjv53+y+ueZQzEM
vBXOEnVPG7C1mw05UIlQRhjpiDYhIX+gopKYZIAMqUyxB/7ZYv5Ao5AWLvFFnEeK
3VlgMIZlOBan10NMOF/DTI0XXNqUsffLGV5qN5UQqRUHGD2xeS/h6nlIPc5+4i8i
h44oh3H6QzjMramUN5+zZfRF348CP3DMWWjnhg0rlXVsBzLeWk28HweoJvxCnN7+
zFSFljj/Z0YXEh1I7FpqwG/GsP2JIZio3oWdtBv499kZO/gqoHYPgKzGjRTDXfCy
ocd7ZEjPOiMKmB3Z+IG2bvsOsYBzUPGBfj9smTVZZJdywKknngiIfQHNQ3kmgXjR
+Rtihf1XSFW+cCj3EgP3IkcAWaoK8SYiSq6jTFa+tctJc2wl9staPyIgY3RmaoTp
gx9ffoJ5QdmTgfRHQJ2Abw14zw8ceEe++u1Imi6gwkh3hlwyKuU3ElZXDuAfTlqJ
ApAWNU1uyrPIlhfhiR7RYeBRVmEG8SjDstXoCvFQhENnXaW78cqgXaAW89O8hCW4
mlyg7tjllJytm+5ZGbHNPCOGD8HryP6MICKNAtkvF+s4E/tiAtnLwkyzoSy8kWOw
AEi8DobMc6sbJjS/g4d0One/JNCbXatqRG3ZXUQ9rulcc0ix3eWZIfGUpI8uZJv/
7DYBOaIWz9j3yIU2sB2A6prX3i9VbdujIVzY9Mudg/nTS8w0yNGxLRWUs8BfPsQ5
aY1R39khZ5cZ0XpKrUmN0/FWOzZs5fGmMFckFH+NFlJ0jROnHBj/ze6WREoUmf7Y
lI8BjbCRkvZiqGDs4gE3kYASGYPdin8gpaplh4OwqlRrYzfeq1jncUtQq7sCLYPI
gg1JG0+8SBWVVQJjbSHfuToY41qss1SsxFHsW61VaFpBL1q8cwKjOilcDCq6SW6o
+5fnZ+eRo8mPsF7Ito+2ZhOJy5m7JoPFVCkz+jEgNPl0Cm0es/TRphfj7VYSaxct
qIi4lNOlhxInB+8Od02if3zKepQV4ShJSyHRIjBei6I/YxMrYHsD+uaAm8jqmC39
8mYEQwW4vt8F+1XkQ/dU/hZGzm8Uivl2JrXj1T+eFTsSmON4SrZnZtapA8uMw6Kz
jFhDec1VOjh0xFdN8wFGGce8ofqRK3AAhD3texFQjx9dsbAZrdQU6n4VD/HLfflH
qmGo4c5WCgQNODzktatB4CXsHoXqR/DXVxIFz0cBMc5K7bUWV0yLxfpEn0fQjC8l
AVLJ+4ArbbEZiXpt/okkbbmnIdUiGJQvXuMqU+npQU7HVCvwAs6TQumU1MhnF8zp
kbLtfOHpT3MU80O+ezGP5uqjOqBkz9J1tVVIe7+zxj5mxJkQKnLKU7hWr0hXpn1d
BAntcuInnuqWeRPfutxx2Ue3pBJ0pu/xOz/6e3GOYs5fXxXy6zz7qfvH5t1PC+JH
eXeRxxevbJjO8wk0avkQXsZdhm1EoaqzAnqxv5VgVrE0VY09k453wHOaJV3JuN81
vRSNWwpORvHcdNeFk6QdJ+cZZC1xXeCKWz05A4ZQnbspka8ctzmDDKLcBWVqpMdK
Lf0raKYs0GuPv59XYa3uscGDpBiwFSUIMYjKOiLOiIP1gPcCEYSTcG7jVGR2TrLt
25LIlJpnhqtDkO2aP7ZqS/WzuWEq/7Wjt0LEvjL8odNH72HFVR7dxDtSFHiI77Cl
Ropsh0J96Rb/evF1Dp3XJ2F0b16Yv60/7PuOIoKq9RRXjMq40xrkTiv8NNub3I4N
sAD6Jm5TtAkm0BMSKVJ/07YjWlYbNj2DwBFfy6qS2eXjCVvoHPZDMFyN3QhS9i+D
MOzuzywzllEm43Go/ppKpqkCKtb3q8TasiP8XUy0+xj+zo8bLsC0JRMEdvs1ptV7
lYv/1CG16kAqUFxABjEaDNOYDT+dATqmYk9zlh8JDH+3uysDUIojoL3G1ylRf2CO
DT0LSRKQXF56UvDPrBJmZf/hMBxSOEG0zek+a4nuU8IGiUMvFAftyfKhBk5/TEy5
BPABF24UriZP1KENdCEAnjh7iGvmCD1i09iTh8buSVkdytyxyHHf2hIiL7YucUEy
4ol7Wa0M1iIztvFdL6nwMLJ1Ke6WqkrbhozdG2OPXpWP/GzwWEWZqfUx1vyBVZTi
3w5h/pgRO0SutLwtyjXUymdF8XMpZn1vczWAck3scccgv7DXMyOMKFBQWK6ZD38T
hz3J9KCRNShxGXqPH4D5GJ2JojkWvm215J1ttd1r8sF1efD1vszFxz0YMwzt7HjQ
F3SiqYZNrovpPpjcR3mrWWhHgRt11IdDuvnDDkj8VpHWGZfMn7DS6hY/mYmgQ2Eo
qslxfBi0I0Ten+x4HCrV3l6IA6R38+2wSJMbALsfHlBOqaZ226WMtX72pv5yEKEG
vDKis7KsmjKw2jn8wCdHJsp9m1fngklpG35GZHorFszRfSA+vdEOs/385PbPy6yV
VkhJxOezw/7SJASiBRtswn7wZM2YDqSBjQ3f9RXikSxgOPWuus9irF9A8jof7MUr
2Ds5+Fn4XWyxL5raEW9RLAoRGqqnIz/wI4d4jZA9auA2ycYh42deFRZTw1NiuJ7X
YjZeA/x7iywOzfHsl18v2iioAJQf/pJvOsFsIeJf8erV6F9jJ4zrGeNKiEccpcD/
RY4i3owRJb3yHeC8t9k0zyo8U1q+hHzkLX3dpwzntzc=
`protect END_PROTECTED
