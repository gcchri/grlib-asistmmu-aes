`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJR4gllsxkCren2IrsFGhjZcCU9uRmLeBrIxMySMGDTL5waSw20dnRpfa7npt+1L
3sjajTWdFgrV/OlKO3xCIdlzVAKsx2sUAX66gmMQ0uSbNVSsfXyVErYAzo9+MWVj
oM7Sp6LsTvAzBq9Re/ZVPd2LjA7pu14AJFkr5IMIZqNjFf/9FEiKSX9qGJit/vEb
cMPqvKEZbPaZDYKgzWEgtjjPOdq37aHRPjPzJIKdeyUQcSOzUrPO1S7wT8exiK4w
bKMlueoD2RLn9+RBAlt5SgaDIRC2VbWAk0vmV3LIaKNT6morxDJEKj30muLvULY2
9a8FMCLkD1AgTm1rZ7u4Kp5IqBWs3tu+Bz47zFf8sjp2a9Isq6r5a3Xz0REpTA8d
`protect END_PROTECTED
