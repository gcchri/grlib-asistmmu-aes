`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rXhnHt5gixDvKGCXW6uZzgvfg/Xf0Bn7krr06MRJWuOPmCBKbFsATdwnwkYXHQSJ
0U0xRkWZkYEYEWZUIa8Jki0QfSr7CCS4YkU+dourvQGdvg7YWSk3GFtkNlJLUuXU
TqOgwGHhgT7WeF81U+QLDpnpbPWcn21PTctaTBP5o1CldZMTBOWBnj8V6gJ05Ylw
7b8G5O62jC21rcOyo8TP9XQiQTwaEUM5gvxftUAIbSEbgxq1yUvXZ/A1S3U30Sk6
GtDFEE2G9CMFVN5OKDOmO7n8vfDp6nt38Ec4Op6jy5rpyBY3c1UHpV22P4hzwMyh
5nZYJVh/wGafpNXeQEYyfBYv+b63/5n/rEU7a9bDntdmha4A/WEhQbryLDaqw7ab
2UGSbP9yk91YYi/12eIgW5zplZgOzgOeIpQJcMNsSjBuwHzvene4oNpiFEkZW6/h
m43ul+2CYtvECgPCIB+eC/Hus+dDfnBrOpgoacAkoGLJTbFO6AhGZO1Tl8GwXu6h
Bi5E+YaWHj/Iqjyd6X1f4/Gnw0EtqbcKpk0qKBWCB7eDg5xahdxeHwhR9cxmxDFC
XyMDh50aCfRJlnafE5WoOhQqHKzHRxxiPaKFCAEYqma44UmPM64/uY8GtbP4HxSD
mU0B8uHEKX3W5KyndpZmycCMcjMIcdO0aHKy5eEqaUKvjN/DTRfR0Hv00+VYLHg3
t+aYzXrzYvKUj+zvpvXGqhUKE6BIRBs+O5jXNw2RX8/FvLv8G6OtLbVmXP0DYKEm
hYULT0B47VWC3fl/X2Nd0/S5UqMaHK9sBqPIA/a8j3kpmmZdTa088ZtY0E88GsDO
Na4v4uvfLkwjLaERVhAz/IWZG/I9UwWN+b1eqj5kkWVAhPPLhPgpujfzjN8Fa/bY
mclhbaPmEPnMxu75+MPntBSmqOqqdoS5d3fGbHS47C9X1jCdZqFntTTakmondfvi
bo5W43oXWyMjsHUcbu3J/W8eYhrBpAip8m0WdhrzkvikmvF1nc/MYMGoSj0xardg
REfc2D+DZOWvYZVhF1wtXZIJBI1TR4lHhYSmG6DgSrpFeOPPjc6nzbrkx36Wy5mD
19FgKgPn7vMLRj2x5S4oQiW238B+myquGFJTT2sX9SLOC69G10+JBqId0SUiz2L1
eebp0w0De80p41gUoQb5/KU7lSVMMkPhYZHgI994Tlj2NXpNK8aqPvgpTq+3QAom
qkZzddq3Q6FGU1Tb6LI0t+FMfOaAXX18aD+ZK6sDv1CQcozuQxJfsm1Yj0L8Z6zH
Ywe7ZzrVJ1pY0cXiSB3pM6dF5dBW+Yzh0sitlrUdv7BVFBYkV0bbVSOXpxPAiArE
tAbv9KwvKdja72BHJVPsFO+VL/ba4QplATdsuCuGw4lM77sLZS6qnjQFl8uRYLPc
4Jcf31YYZWtXUy8QVRz1RnQYh5c1wpL3LUtZFWr5Rhg4UVnSVuGcmCXNbbV34Gd0
O6lSYCPZzWDwV9HLOj8pJipAgYXLtkrtLTl392CI4qdkjhNwHSXoFC+Ul6GAZ+yk
aCmc1QQ0Yye5oi+mgrjU5yc/KYWP/IpMonM119yI58S6ThFG24b/+V9IDzgTnufH
rzfRPqjY57A+sJgoYIVxJnUdHtWFuDw9ZW8NoiP15e2OpNLlRoNhO7GNgF1SKzCU
3HUYBpzjlneOZ0f4WPWiHJniL8TGJX4sLQqazQzUwuY4KbY2YXgbJEeawo8LRLM4
RQNRaU7FsMi25lE71XEDtcfMHnXxVc/hivcNBBRGrMh3TNHSVnX+gJN6wdRnS+pT
jSZBamjOubrfaA8lPnEX9RFLUODYsjoHnB3wBLwosNOtGptV0B6KJ5hNxtwSeU7Z
zJWEEbD8ontb3U/rdaOh5Hle3yawBcUhAgxCXNPgFthpay310gZjANNNO37QodYh
1GJtWXBie6RvCI8Yc2WGvEZHov1vGsC9SHUnS5lANd2jmQuTg99fpunT6xM39dWs
09PfGHgbggjx+vHJ9IyuTuiWLCANaUPL1KXJJ7Mg931/ObC7rlhgmzx21Ci5kviQ
AOmYV0a8REHHTszWcgBS2LfR9C/pQnjdg0oRJ04DVGZ29b02zYQCr6hXb8Vr89u1
pEBiudGS9y9ne1C5zaBDZxlXZKVEpr4uf1YZRkLzpn9V7YlNREkFqkR60YH/uQpi
VK1cAAoo84tw+basMFmZN5KxEoKxnPkB/5C+r4MZQyQfsfKvPDO9YxacLitr5c+t
HQXJWLGexOiJjj5nf0DpL6FZZCMlh/2SK9IdLkEE4eZzALm2fa7BN4grFimHeHyZ
PGPTIaMM3IvZ4Bsp65m7SaxL6ER3riQyyLmi5Slkf2yhEpCOKRLpLd9yJrnlewvQ
9L1IZcgO2jrQLkyekZpO0UHBINb1xfnljXU7bsNRPXdadXlI+PocepMKPBObgYwH
mFr08+MJQU32q9AD4kl0Vq3kOO1rz/NJD8UoOWgkRN58QFrbLH39l5bkwFremT1w
CvOcQ+Wp+/pB7WHPeBQHKxjmIXfqy2G5HYSa+4IL9DGlEGp7NUplI9AdoPwvQVYy
2x2uThJi65Ye52PVwhM9v9xh9FcNfKfCE4b4gUiJWMai9HMvmMG3Nxhp/+7olj2D
WONFIarFt2dAMdnjoNJG3PuwGCk469y4bBeirwGEhkKlL7yUNnVRdnXxlqjSNjY2
YHOQqOg9NuevZw22Sr834UXtIS64z/Tx/mnWxO+46uxm1MQxGvuofHEXKi7/D8qg
1DVIo+r/LSCrbimSfSPReyWPOw0TFU2qLXW8HT4Z9NGSROsg7aS0N9SfO+luCEpd
DqdJdkvIaqQVu81ARvbMWx7UPquSMxpY5FFwxpQGnXrzTjzLSD4lTVrBk35k8dsY
cqz5lkyr77sl9fBI1WUnS3y9WSoH6z/Sr02VXdc6MI5sB6eEpvr2BscT4yCvf5iG
YcqxmNdxqHVloo4jGQN0PakoWK8hkB13lt98WH41qpybSrASY1nZgGnixhUg7X9e
XuBq9HPziZOW+/wn0lqqWfTe5Az7BI1GUBPfJoXnqOCttIM6rYnUNlXHv3/uWdTu
X6A+nRUyruq01j/XTNdLvBB/W5QIFTm/8A0FtV3BYTYs7el3xSTEO0mAhGPxTqOB
mFcC1+qYtmXnimaW5DYxTmIxIYubyWfqkDN7FhV/mXfcPS9W9DOwUDlR99xCyFte
u/XPa3DUFjlTb5C8Q42JBeDEhXpbgU6VT6l+wH73SO4AsK5AdyZKHNa6iuDyFUNe
PNO2XoqLAVPEx7b7qv2h4RCXl+jNNyxeu99igd02E2o/IRabfwGONZSWQrICbF8N
86MgC3wt+IBW+nYix+obQ6DpJ3Ff19aH5W2mEBioKfCYZ9GaJrgN5IBdZG/pAPVH
xqfdWbOGoo7RxJmFDVzXw7R0aGwys8/YG0t/D6VLoye5BatL4SjUqwVI7QnokBb4
rY4NTdZNxxK3xyv2Ni2qpwar9kWg/b6llho9id8fLrqS0hhXO2X7N12aNH1gWOHk
fSXmPkpBNUfKlxQZIEyXAcFpbEGf0v95zyrzONn+ucdZYpVbOvWeoLKFNLnGxlfP
eh4fhG/TFle1u7jMkzehCUXEjmaORoTSDmh398zLxP+qdlJXIJC3pSTOI/duMVG8
8sy4rk/jg+EjDBMYXfhxnCjgtKnP2ZJVT6xZlP5q5mTkR4dmVRX937vIg5Y1fI3Q
J5tkKj5We0U7KqozIHL0cH7lBo4m+LtIUJ3zuASmCV22sPyV7DG6TTfgPy9fRtE9
L88f0InpxTkTl8ZIc9Wq7n2ZwBY59uVhr1uVe6wYZIQVR5joVI9WpNQIUs+3NoLO
nkWpbIYeL2r75/wImcoCy6dDITd85zutkjI7iYI9tW31g0QZvUqGlNn5BmQuCxdU
FqLzLstdD46OdPrqeHF894eST26bmZv0V7CMdBrkwnu2j6KJFlgU2Z3ZO7JpM7Xz
ddaBEVkT8/6IikjyQTsNNu5ZcEUY1bWWuKnqJRfEu5isMmnFd/AZysT9CK1yhwCv
Rov0MPONfCZjC+B7/sCIxgMIy3sNt8FShWDO/0TdsU7NwbG6MP/DUnFQWYE22gU0
AriIlXSJ2bLudexS4I4yXXcsJXadUjuRam1nSEWO6T+eiUhZZw3hkggBqZ+fUuUF
+Zk9zre5LtVRnwp7bvF/wU+R1rZ6waGP9qqrQxy0JSTd9I0y3BjLbW7wzEfFC7gn
EWzmnGDrHtbRRcrb4DzrhpmNh0xssy3v7N9WMCFzgZ6go/F6U83ja41V0hl7E3uY
iVpTEWXNRxilMwIq+8Xmz+oIbPt5EXtVSknX8RBNhw343iCyMmvtDVE7dAt9D7/N
7IQPgT571Z2MB5bGZSVnO898twOwqUooOcs03Fmegw2c2JabUhI5CT8azmfLAcTJ
xInl/CRPXh6QRgjfJTZMS5IswmkGV79TDmhf+GGZIoZb2Y3TZxfcKH/Rgk9D6Bly
zRQldV0rVpRDcwxmh0kDFGjSGWWZ+fDfGBqfihHx5CWCkQBE2+OGEBTHAi6PPxR5
pKAWRNeDkSbfuFFuM8f/qkz5xNnx36hzAiIU47pLGAF03sfvOEbIc6Wqx9X5ndeJ
Bz4kY0sJoIRqZ7NgI5+d0aEdYbhizYGnsyzxN/Bj5EgGy0TL+QNc7VrkbcOdagev
oF6iMU1RKfYEvOHsQxONTkerf+wBNfw7LXfhIByUQjd7tEJ2695To+WC/ZmYmj1Q
HExdKI0IPvxX+CDrxWp9+p50imZgN8FNufn/t7G6vdvOaTFjM4Kdley5fXkInMEH
wJV19WgQkoYiM2ytSGqlmGP6fVGKRG2M02bY4hgZLqnTyBhQQJ9omu41++XANBhm
OCpTOa4g1JLwE6zedWlJRqJ5/rzzNqrRi46qL2HIwLOuTzdRK/uwKgIT3aXPzegq
mjhb5F/Bp0nCUt1SnmRr6bnNYHuO+CyPm2z9MV/00gJObcpqAURwayFHMbdjcAgd
lxisMJs9KTJMaVCcciovPVArhYcO7dwpM0eKW/4hS78aLKY+tXbuXw40vDLyeUtp
iP9fk7D9bX7AaLA3swXsWrKFEsdNFm2OxPLoOpwTwu7JAS5OZLym1ny8ibTmMdBa
/p61+2GIz3XddsVbJavt8KN7f3/ibaJmiR8x7IDc17CLDZ5HwN/R84SyfqwBNSaj
wsazUBuTdNv6tYErhk40jW9hR5XqFOJqorS7yzsGTw1tNPWSDjYz1xbPpC5yflar
Q3QBMTp6jpgaYyoaYHgXfTQuhLf4CdUK77NO4hvf83OD2M5ctFR5GmohHS9/MJq5
3Rldwml4Hwarx42ZO30ECYAZAtXEm8LlPCVs0b28jksPracq2NIZErfy6auk2IWA
BzcBk+8I1YyTYxpxkqfayKRrSmb9xQ6hGXV0dGKDbSCueh954eo3Y1hTU4AqKEtg
HzcAw4aDYwstdc43EicrtPhcr3jKO/k7S79LRgG4KIG1q8IGSCRzghPtEm4Tve9x
kBl2vvAstazb3tXLj8WGEi5o2Oq2pT3A35uMf8xwqAkZVQLutE/AUJh+AIz48P+S
Pq+zSLXM2LRxebnQRaKdB61xOKmgYbBxFKYNbyh/aOgROIYS5iPOTfrogwFDMnHZ
RFK9zPJF0bzvgdbxLvr3o31fRK4c7qClgrwMMGcvIP82OtOY1vWb5FMs0TqzUkIw
sGmRZHmxMPKCQA+9sG56goEy8NrC2DtrN64TMMse85wR6V+WzUvqsLEeh13ItHEN
tsks1oro4E3zHDcUsCJNfZetmRaXafUNd8jAhHB0EX+L4THCeZ7naHwxW5GHcQ1x
YiZ7MWacQB8p2iR1ckPH37Nv7OS5zZ4flwMIC1Cr4O0cZBMe6v5qWj7wUBY03U9h
B4yIzWWMn55nGoHftk1jK3yxGctd90Sj64PeJdLtnA1IClWjqs3eL/52SXFu/zLh
9Dxy04crJJIHRLKdww1z5y66fzeH4b2i2kfeco0fqmM8GOzTPY9RgE+1Le2NIeRc
diK5kAvpIXUpDi8A7g58lkT9801STHi3iS9sNPaQVESN5ymd+2L3xZ4Rnu7w5tyX
V726yGj6QUUMHSdK1gNJnTyc9degpl2iJOeFfxM278V8Zp+fsgOSDNINGWW39rya
/EyV5FVp97nC/TE3SMJIk8ixVidjddg+k/L1Zgw+RjaVTVtU4dj4NfQB+FAnqjbB
p/gWFaTsHA9TQ8dS8K+U3In1UllLa+4SaU5SF9/BEFP3KAYXerW0Z3+gE4x+/jJq
zqPt5j4wMPxhiXcnrc35Z9mqr5CF0WgA0H6uwvzOf27HvWmhp0jKACQ2NvIMdyM9
wNsIjLbW9EQDr7IJzsvXf915bqkDKY475AwfYn+Z185iIXj9OipXuK/Zw8S4eGCE
+5hCNgEWwf0aPBnc3QL1G6Iqubz+m9DQyVfa2dHxnOD8VIvPl9GDQo7QpWXLY4zI
h+GKjymKmhA2YwI7DG5AWsZwYuWTyYXAVQQw1BEoh2XZhu9dH2k7g2lN7upDo5b4
u1UbM/mC2XuhRYXtR8HNH34euaAjzBNGHMA6ZTr64XERn/LfZKhR7NTZqU4G0O6f
+RbkeTtZXMeO/m7Rjl6TRV1M+t1v85NdRDx3w0aCsBilYVqosIQVFJUyeCFEvlr1
yybMhtYks1R8RDK+4FYvrqvMySqu+eoSvKVQVN+hq1GsHmBkCU5YsnRC/6rW8CeJ
IRhL8IuOBKxIwwnj7rfmuoo6zFIDY0yObW0+AutdVnu5+WfJrvu5pfMvx0K8OJes
gFuX1SN+Gb0Ik7rELh6ZSKK4TSdlrFGQBSsU3PlKzmZfUTKlZgfa4gZcxB6PZgTx
A0uP8poGsCPDluJMyGMD7ZW0yVwOWeodhP8ifnENnA+mGH4Saj92eSamfoSeRN3G
jN9ka6D6r7gZn7NE/EaA2TQD8H/ygcmMdWB3pbEHXhlxNqj1E/bS58hDrraNpkAm
g9VSPAG7apwCK4Ljv47qFUxt1/sJhpXwBE7E+xK9ZaODQ4ANYs8nHx6bFQH4vOaq
ETdOpJ4+DFC2RSGRu7TOnvanAcYoU/kVrod6E2/mv1YZK4p3D4IztkrtfdzEFh7S
9thVd85ApX256NroG53JPqqpXHyGUuAG2lO0lYDLHTwcsRNeAkBL+vaR1XwobjAn
l5cGg+3mgb2R+/zDaCcdPDuE04FVlezO+utUpHHBVkZT1rVmH6UQj1ZEUlMbvbR8
LRgqH/GWS64p51/faVl6CpnoKZbQ7AtkR5m+fiCS/wLq1lDv7zoTU/k4HB4MraMv
Si2fr2/ybLcRfLMARS7tEf5fHbScfZabQEbm64kCsmrc2Xgba4Qkc033oGgZ0aSV
EkvcqDr5xeOGSpm65RW7WWG4ZfFCBKHKnlzAn45SqUJKpbK/Lj0QE5M+zqbbngOY
MebraDZjUiss0T7e8UX62zRTHqOZS2cIUjLAWz9/85Mo6ou/ow99mbfUex1AETJG
tA3wtpZaXzJ9/XrzpOpn0a8Hj/fzt7EYTZJEWSweXaCfP9BWcUqUwwsZ2YDKhP8j
jJBYkjquhJr2ip4h6JpqKupTnyqSHUbwSmiJIP7WQlnWU7/PQKz2vGk/9j6+7kEl
woDU1tNPDgAIGY4mmmp6i5AfilD1qwW4hnkLW/aeROUo3L4MuUcAgi2znfMxQ8K4
Rayf8TdJnw2z9jqiHu/POvKF9gRaM2xNlFIicPyr5TgzHNuDqiy4VaZmi0PclZcL
iG713e9AbEzWTBEzX7I5q/lIqaV3IRvJqPCu0RV5DzmdkWm0WqHoey3teM0ULG28
Al2mO7xJkbZUChgBdnce/a61/j9CQXkf3fP4qvISCntHZu5t8A31NdBLzcGBWMve
RbIQPxuwSIHrd/yvKxmWnkkQLFGIrjx3SNyUe9jLHxYGvpv/vW40/TKf6hD/bVde
lW1Xofl9EhFISG0Brfa20NXVnfqBtu61LJer54TIg5UNSSaTPOw2K/hqGXqCgCwH
ilMpMdQ5dk2t8+5BfEgDbDPDkZ/2sQUdVMCHtqK2Khku5YHt3R2uqXld7avND5KD
at8WUZN8ca2T6m9RWU43T3IlyI47cKWfMycd4YkYjSGpz6hx7rmZ44Hd5jNAWjF6
TK10peCW5mQlXqHhWzFo2YyeLv/YSEBudYaU5VzJ5ara1xCM2VUn0uev1XjChhxc
XsSJJ9HP4SwkyKZnW8g3P3hF/3fYs0l+NjjXSHtFCCWSzSuN/thHpLa+46NAzDmR
sOPlbA+1wIaUmMoiwnn3aRlxw/ntHQ6znAXBt6DL6Ocia8ED4TRP0xtM7QFpxgCa
LDGNi3KRlaGz74WbrkPjkoYn9vNqqrkgbWMkv5w2YHe21bj7sDz0VBsY72ZpzmZo
ibDacrxRmSwz8uH/hUZAtX4NVpLQGIWqZ8ZGr0bv04fdBxt33MY35fIaF7G6GuzV
v/cqpa9Gr7i1z4W+ffvbsGiMJudn+auZR9oganQvbpoHfG3sCkqAbad13mLhCkwq
PB+oFNN4dRQhBLywDcs3rnaOo6HtDuSS5eU4eEp1nG9YfS3qoc8UNh7gXNPE3JBk
GESqiow++n3bSH6xn1a2E0mAIQnZfmhNfnNvtFifRCKChjjiMpZ4sjEe90LbnxJC
TGZ8WBB+Sfx4LFTqUwqd7Supdd66s/VjT9QP0Czm5Ka5t4zyzl3opId6v3ZDnVPB
6aUVIEUI5W8NVOvh8E98fw==
`protect END_PROTECTED
