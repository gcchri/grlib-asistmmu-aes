`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7YOoO1lkyYzyAKMXlklbnjpx+e/uXe5x4Kd7moH+0A5panCuEtqbCqnyqXAXqUND
YNLVk/lKb6/CrO9g6BmJiOZHTxlduB0VT/QEfsVikPSLi9/B9r/uia0NT8y+LxvS
onG1K6zitcD1NV/ao9BbhmVBYxg1Z/hl82GoCR9w/RbiO5aWVouPBiXmr+5Ejpp5
PXH9IqxH3h4w14R90LKvuqscbqglnilBNCHVBKLdnYKQIiDzeh5XwA2bomOI1Nti
8io0XqgHvO/Gg8sYeROe+aaAiXN58GZBQ9bMksayluwZEjmN85TgHpA54oBUek5z
bhn4/2HMkJfiahZP0KwsZMkSDO1+XLKWF9FS1g6NFzyqONVD3kXctjfELEokTYnT
hVj6Vh5nB2Z+tEqlA08hIt2kKHB3ZzCaejlly0enobsozwaK5vPq28skpS723Tqi
KMoZFARckY32KS9vMb8chdwVYi3Cr+arB/vePpOKKhKH8zu3qd7Iue+ZMofv1ZpR
`protect END_PROTECTED
