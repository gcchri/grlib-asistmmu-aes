`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLOiZLfwwnDFyq4m0EPRWrJ6fgjAeqsJxM0iBRFjD+2Or5g4BvCs2mAMp/MDV+YT
PDaiKHml+Yr5OGTvyvb49D42aYiLeUqL3UbACHt9zOzVRhYitpqOouG0oqAcKQQp
UqDryVhR/9m8VzEYt8edUsEcHrTyK6E3cCxyGXMywv9ucmUZ/E9OwLPkDRrRWnRu
ynVinihMMXAzhrrs2Pd5/MQuWSTnaFE9w6e/EkMFeoOFKCmIpyWrkI6ki3NER85A
fzXUXr3Mo21uZwopj+puH5JkJ7IQImr2FzZg/hEvNVo=
`protect END_PROTECTED
