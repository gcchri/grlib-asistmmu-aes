`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
poYQeUqi0FZguhv24veeukxt5JRIG2F2ahmFeOiRsTtgT03rV3xmLiZ94XOJgTNE
hJM+HnrHEdUlFCQDCLbjeX41Fi9GbEI0OU4elVn9/1+tBfd9SZbmQTzhydBaip6A
i0NenDHVCMcHaj6h8dRS8Mh6PJEox3QPv0BtIerdJOxuXbX0DpRpPvrELch41csb
nl2rYf9RUZ21E6i7maJ5C2sS6ZrW6wyLW7FkvIYPEh2AHN7DZtaVOGY9YE3ln/6H
AmzwQIqG0980U00rNCUJ0vuZl450ueoW1Io6c1c49vac8qstwv8rPmsZhswm6VAg
qVtCiv112dX5tzjJ/FU4AxgOjlj5D2QAbzLOmBoRhHDbZ+iKH7gQ7gIytnG2FWEQ
4SWidC/C135N/AFJhgdZKBV1CL+X86JVXPNxf4MjKMbJgTq0t977k7SfsG/Pw56m
FGBdsUYGSXQHfWji6WUqKB5q6Cc8OE03K0Y36LNb42V+ndBso6iNjHybBbSDZ0sN
Q5rc9975gJfDRItlgYKLLMSp/L+fLpXtFxseMqa9eM6iNgRjZas1ItPWw1VcUlFm
zF9gV0pHhCC8lq3xgUrMI3C9OwtuzTW8EI5d0BLYlK6C2mclRRRsPqoKXG/mQ1+Y
ymhxla04comOFaLWixbXuvcRDEiQ58IPv33Te8LEKpAzD8eA7a/ehWIVYcn9u9oG
2AjVabQirSOknqw3X5ukSpKHyeyQpYRWNElsT+dJadsqIa2JMIG3Q2vyVxnqOloa
/KDW/PXPdj7hnXRdM3uaE5kVHWl+vgWm4qb+qaIeWiA=
`protect END_PROTECTED
