`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tL6f2WxF2f8HBo3iKSF8fabNf/sLcFSUOtLS2mQ9GkwCCVUKkt3NJ0PBpSq3oCI3
ymP0qxl6ateuZ/mSMicuq5EfPnltHtxNUDBb13QoEL2NgBS+f04inA6Y1v1mosdd
H2rGv2ZyN9RHGsaPhy/FVOCTNg7ZFKaAIgscxqC6ZXDwUicIdrb6csMAJUXkgpyo
gBZfQnpM2W/S33LqcM5ymoCOc1NrBwijN9Q1ZPYChcuePo0CX7cpqMj7ds6u60y+
iX43uM86ZBoz9CoX36pUd/URfpuJoOILYSyMr+RFzeid01G5boiFlomfaYhy/Zq9
HQQup3DVvQaMlvXG0/o+aBgYNrcTc2F8Y+PiMnKdcPv2XBfyCrmIM4X1knbuy5YP
7Z/soeIVRXzqKLVHv4JSY+wryqeuOlB8EI+dbAze59cyOKXeF4qBFyyhW5QRpVYG
RkLBedM2JsWkGymupTCTOIHSdWmDJOWXQmOof4ZbOogsktkI+cB8fMHCswRIBwg9
u36F5vo+pBqWdv9OzBxe5qAoT3TZKHFF/xxEWbIsKovQvzSFIuISnDymDkMoV4Ra
usO7LSqjX1gNI0HXjqdHkffH4/IqBSLj2Zt6k0y9w2VlW8rxZKTUaSNB+30bQ3l4
6Gw71NnprcTXqx/iMJdD4IUUp4SAVuEjMYFut/hmU5yLZp3Rz147ig6lRWa//YdE
AdkZ0t0HI9NzRSBH5UVtGuoUMJUVTmfSCaVUp4mPodcvcTLwZ1/uowC9zCtOpgbJ
evmwg+Hah3DcdHa0bDTDvg02yVQIWuEdh9BnjBRp/zUxYWVqXlEZjjtgnGyqLFmH
OagdMgzB4HITjW1KIAsH6yo85oPF/1T/GzJul8r5a0h+CcXVP52ax0LZs8jq2+rs
jEzQZWN1PenhlViEhuQviugHypN0jJ3gXbS2hqzEGFrr0AwSzs9TGhpj8uFOP6BM
wcABYM/mqxMGRGOyygRlFgFHguV1XoWd3gK7GZGvSpI9HilryJlZlMsxtgnRTWsm
22ghDIUaxYFOC9V44ITe6ktkWc0hR8ZUr/QX6Q0ZZwpxx34LjWXeCsXQv29j96ft
F4vk1fbxVvJq9wXeN20z0HkPCZZRuj5QtxVjfXC6vnkhEbek5K2IEu+R9kK+H7Ve
`protect END_PROTECTED
