`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZlKomGhyBhRAJDNlo1qNhVlcScm1P0ASSkNRp6NeGmMzqbikYJkQwHSFf3P1uRL
jJpuZxaA2paz0WtdtU18pvckj3ATCQml/GXmpFo4YXrJ9mtFGSR0xTO1DWgFQYEd
Seu2ePMDHxW5l5oz8D2lpgrn7ogNOjTWJEwgejYZAYPEkGpY6lzNpvcLq6sLXeBy
8XashoTEOapuiA7kz8NjlYYQHhv8tC4dX6YXw78TCwwg52Nt6glM3iSKNLrY4jlK
87a6Qt9c3S9FYe/AqprdPMycDL1XS3HOYbZT2ufLkbMNUH2OjMk5q9Wis7sIOpde
DXOa593BeiMwGXqH7F42iZQpSddouBleJbkvoB7ym28ImazTlgKJkMOJYT68klle
VXGSshyGqZ6wQKFWpFAVPQ==
`protect END_PROTECTED
