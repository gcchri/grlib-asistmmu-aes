`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yyw3OLFR0OeO13PZ/NWoJ3WbbEpd9xc6HqfW/nJEyqZJsPy9Qr62b2Wqa0IdLrrj
9AvEXZLunibHjyfX2LXHEkF3LEK38GwpcZcDd0vyfchhAfVlDqjAI9LcerIc5kQP
Zf3gyKmRbfKWWx4lmaCCuG/h1g1OCMbwuOFPmzCtlazvDj8kMUsXL9V/xHqdm4/e
pPBs6vOzOlYCt5rUhUqwMNoNHUV1TQQMoGXgN4HBXGTw3CEKkDBqsQUY7r7zWHYZ
X00F0zUGHCYQsZQxFi5lqw==
`protect END_PROTECTED
