`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLmeJ+FaavV2/L3acJGg8KsHu73mqS98kRBlN6CL38TUxSO9XjreVZVDJ2P+yUq3
cFpa+VLUqF5JT9wvmQMZTNWLgUAtxlMvwPmOs/QEGfUBsFCz9CFeSlr2lKF4neeL
FuAFgcXRL+ZUfpq/uL0Q5EVmvNM9KOjxUBIXPQMJNcn9wcWh4pVOBQRNRaSimWUE
xtt5/osS5dinHr5QmTz3bOfj5hkojS+AK0WH8ppov3psIrpVALXyGbjgfHB3rT06
ymwNzY7eThRLcweYg5MftHIe9QZrH6Tzmyb1LlwwJCA=
`protect END_PROTECTED
