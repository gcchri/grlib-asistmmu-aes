`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7q0/EXmYAEDVAzDX2b66HoR1he2KEtccoZxDjMzPIpKL3MluFyTHKpboav+r8VN
HUCDHpnjKu2ATSfPo1AsRGy61CkSbTTUo2JpCaLZkcGxlRf1Ih5F4lE57a8kJ0cv
fRPEOuN/dvjYZQQvAj0F7WZgXlJdoLpZhMrdlgmmSvHMu5mECF4KGQLuRTbIXivx
YOJhwT0ZTbxdZ/P5Qf17q2agrhbauKH0wIDuw5kM6HWNrCNoqD/fIbuzl/uhN32k
tRfgY2OdW8oRKo2wHjzuiYyArGf83xbyzcxDYpBpGrHPHweURKO7vCTErTIt5md4
V7aikSu17Sekx9ey6PatHoPeJ/Dg6OIEvUFKcWiyeviOOy8dqPV2/HQG2Yd/rDls
VNs1SH1ohSs5nOioruIQu5ZBOv+X0tU/Zo13pL+H8RpREOFOkNZiSGLFLFMTVDL5
HJc5GLFHAFr2qeXkfqEhYXZcd+TMgTioj5AwpKK2n+xQgSeLIh1mcXHX1oZPtSSV
qYkh9hH70hMHA3tUkIrQN/jBH3HnJrXuU+Qu6M1tw3PCVAvdWKA3lxZDglzGu0OH
XiaMBB/ai0X3i7RZHwE9aaTmUMsdelfVBWzqEEW7B7dmEqbdq90Wdqq/315DjYkp
tS00mEckZBEedRe37C0k1YgZtpmFts87L+PWBp8Un09J6V/SdrP2ksEjrvq7hvvQ
59SCHdm6PjkJWAbNPDsQ59PoLGFohtXS4OQhshod8HapcCLeKJRqYw9VUBuoVxs0
5Nzc4vay47j2JjozZa158NbhxyCQWtaJ+7Fa5mqag5nlgnvibfMfoJ9qBg/6Mup3
aRMn7rnQW44Hpl0VO4geXkyn4YWS6dvXceZAjbdjadSlIZVaJy9Z2blNF15St0F/
WRhAywFe0wqamOHcSi026Iwxgq5+4wRqe6Wvdd8oFlWEuUukSPCowUNlHtbHQAO4
TvgWiV15UvY1x4JS11ojPRVsECx39WFX2nNFu5VOki+YciuV4DgV672G9xvtg4M+
qpgCAdN/mIpBeMuFl+kaVmuXbNjfsp44ttqRlEZrg3T9goRz5TDJUcsvhMdpEqD3
N3rI3MPm07G1/pDUvsejPwqwz/hfO1hTRYLPcTBtL7sK6qXBMHNgyaArCtSTdfRO
f3N2ZrRrMFnXTcUUBibDtl8HrA7ygFN56eIjjUwIC1XFLFqS15GaVFunuA3oyeZx
9GKzCwJXI8Clyu4JcFYLHATN3HdxzvDL4vBj78bzW+H4Tu/PnohZxjK7NjmJZMwu
ipIGXGs8XA3VPp1t1/82lK4yGUPADsD2KB85rCXPb0jLc7/uMXfcnNHXWy72e8Wt
EgcPD6TwrlpgK8by+koQ6sVPB+LlPYiNVMQY251LEnNadkVEpWoQf4ePLLOB4Np0
TBH1YyyGA592KEU902lDEzQSzl5JEZzjCdguBgo+PzOMeju0YMgHEj1/NOHnrUwS
YxM7GQMzK6tuICml5kvNO1tC4igvhe9ctkOyH83UJmg9mnX8FulukyMCqjY7QMXr
/PlBQAnr8huBWMWUmFSOOu1CE22opoCnR/pbheY4ANN3IRm08/nxO8GyEDhwXcJq
ersapERgD49jirprj8I4NubaxLidk3c+exTGC8VyQRmNNfRhJGJBEXmF8AS3Gpma
j8ujjL87Z55+5cC9D1YzI4UssWsuUBRMHzegFtiR9HB4zcHCtdOw/zWJz0VUwGfC
V3YW53M47/rAz4EC+LoPJUrLEFWKCBiTaLP9eHu5wLSnOmZOmC3i9dgoinJ5Im8H
bawJUKLT+AaXcTamN6ywEWjebiR/QpP6zBUdUxTXnVuOPA2x7MP6hOZAPoYur5TQ
Sp9jujg7uZKKnHafrzZcxiQ2bCrfAio3klzzbi36qrLGhaCXASgRxsgOBm9AurUB
uF2WHHFzz2byOo0WBoySSxjjNAhQC45/0VSpF9I22UYfJpftRyaWOMEk4Mn9EKCc
SIf+U0jtELlv6y+1DXRPua7TS59et/V3L1amizuGL9jgkyeEPnIkB+LHw6IZD6al
96UUd9I9Twjj8EdNrgnlXKjhP6I4qDaGxlc7Ff6dKGvFbruNuvEV2dxX2rcWcPdS
srRZf3tx4EqjVkg0pXXwii8eUqy1S1a9fdpBZwR23iEYFgh2ARWl4RF4jMAA0rEG
SAmiJtm2ZzG5BDJCH9zRBLNGufZxYW5XB9HOxIYzSWVTDIWYKUoC53H6mZ6SwRZd
zZJ0/fSQB4hMb5xERzSmQBlQDA5g8LbWpLOcDtA9ovmJnG5cNVqYaENgrsDsTFmI
hor5xayRflsIgBgP9qY+LCSO85Ura5Rm77zisTsyL6X6LlxiqHMMxTPj9cyAEdgR
+VphymOhYJIQbtYkFEzf2H1KSpuLUfTVooC0ijeYk2OZiy+QuixnVjYlIoz89Rej
qFbNlenPirmWfQDptG9maDa7KTQEKBav4saYOyOqTHPuBfzN1IlmKFvTpd0+v9H3
jkgQBDCMcGu/rt2x9NgYEFD2Aut0W2cYdbe3w0VJcBQftX84tJRnztXp12631TIK
7Cx9yKrsyZ9NdPqFNx9wm8YxF9AJw5d9Ptd1btpywdlnnwN26tC9yYg2VnZVFUDw
+yN/cSrRsh+g/eCWBNN8QcYQ1ebUfVAYadoKOJd0kFVuBsZqwsk+rKPv9/Vi8kp1
Qo+/PLKsmyU17sXdsSUNs5LkPXZnW55+VYiHVFLMTrwSjEVdO/Ncpini3FiXVuDS
V4TRdEskxJQtIqGKaZ/9tr4FPnAM54tjuBH7d5bCAH/RbsDNI83KUnFwWFPR5/oJ
CcyrrZDqNszWRonq+d8cLP0mJZk6YB8kFGCpObGMbOEfo20o23g0oZK56sPqYptg
iDu5Yx2Ak5UdMjAAA+hd+75PsOV7zSmrjfrkuwHF3OL+ksLwYBIRfQ+Wm1Evd74+
gahi7XnaoXq+161D3n6J1LatMkMbNLlJcuUiJQ6QIPg/aV73TY/DxWmM4Yk9qCPR
BpZIROc6tQ/pB4AImsi3ULXOWkKWOD2PeqnjeDK6zwDNdTeFBF/Xli2koJnnGpYO
pKVhQVOfmicRtkPTUlIv8mxwAHSh7giNQjHbgzHjt4eCjrOT/1CF0sixsBL4A78R
4BW+V7DQUq/Fxb1m8fYTvd8IigFh1PscixuIKsge0x7NA6sTxVZepX4+tZ4NvJjw
bgOxeXZPL5k4kSACsNtdKi8PmHqeA57bSi7rgOFdIZj9chiwl88DA2ALeVm+pb4k
158/9wUpJrr2gzvs7T4aXp4/ACmCDu7H4Kn/H3OeJwj/vcF4q/LPWNVKov4sAKBP
5upwSwat3vZHIqNw2+m5t2nlzS55Dra2c6igZrZo76GnMTMLNL/kb311s5jvDoTv
uGFyGQCFy5rWB1pQE1QAM/JQmf2FTQKWrKsKylTrvzgVtpNLP4o7+pt+adx2rIri
DL/60qzKmCpcr1tjBtjSHrHY+lWskI2h1ZyzH1IWAD/rmUwlUSuGgjSHArOv+Pjq
dh/ncqMtLjJ1R/XB8kTZu608lpk4D23u6hZWTBgzascp3XHmHSnl2WIiVzwBdCj6
xCClVc6OpCixxZlSluyY3WEfmV+HSXhf9QyoSumJ+IFqB56cWPGklQK49mIbGvfy
n1hHZB8GvEUinLi/8eCjLAPDR2y6WwjzBLXVwAWYSvPkoelTk3qTrADf8XXbR99U
FzwJVdVdfQK7lKyra38Z4MMSuPfJ2+0fzvl9d80f1TosPU5yUPw0gdk3rMWJgjhb
blFWGaBDzDoXs6WllPZsdR8vDDOkQ+erxXnALLkEU7JvGkDFWfL0WIA+YyMq06d3
kyIPz0qNAHHvQSyLwdwpPNOEvtbOSkD3mdzH3qErGabLXG12x+DaB4an7nn2ZKBX
zeIEJa2plIW+YsnHv+ajFkf+1zs0uX4oWibfmpfAz7WcYnC8cpWGw4WXBQhOFFyn
r3oPOJSKaXq9uoYwnBpiKalkYIiK41tTOdp5CS5BQ0Q3JaSwEdGLZhELKxauTVS7
GAiSAjaIM8N26AURzSsWt7s7HOj+YR56US1+AyM5MQePWu8xcX9q0eJn5WcK8wNP
cYvyJ4glXM4B3yrfQAZ0QsfKRTcVi+4wdyI/Ax5WRkAR+jitCp4G2D0WT3fUV4y5
7VPc9jC7BIVOIxKcJ1fFZA/8HWh810DxbZ+eRevLCXSoB6kDslQAgeKRUqkb6Mfz
WY4h2MXHPoQUEsv6D+NZudMAR+B01FI7BA+kDYbR7GXyF1rB05QbvHKVd3f8RWIQ
4rZfO9qMovChZOaVMh5pWAOE0kMHC/DT0LoXK8hsRkfH7gGyMNF3+rNwRP6iJAQ1
wOnpIGrbMFkR0zsrfUcUgf6pPUEg7VFfArG+Cp7LH872hu3pF7yc/W6bq1Sbd8y5
FT2JahdNuZhq7c9OVfXXsSWp6hPv1bjq1iSxY1Gp/dwp6JCGS9ir4AG6qIAyynEO
wIx1+kArSGow63ppgytsg5FYFAJ2xohygePY06rBqF53xLkUbqcDWB01/2FJ9KUP
VJ/zeOXzufhFtKDbfGgANp23HK/NLRHTbD8YieHjrJunyDwX/JPoD+wVdbxZVtuS
nzE9oy0Ta459Ot36vebkja/ceH7+toVs3ODUOZOd4ByDYMcAFpzIK7PT5/OLYcOW
1tdx3xiNV56O/a5nzPGnQ8orrUJQ49JmmSabxv0stxODvQXOljY3UltB6S5CjAJE
1c47p72FZdm9AcEKUA3LUVO8q6AeWsJFuGPenXDPoKSsqYpgHxgf9WLqs2+q6E9/
HYcRom2tXnUmIP+g0gb0AGofN/jXoT/FFTEeV5rKJt2gqIVObpCotM9lkMRyTdoV
ATiUjct9+Q020/vzBjMC8FPEM39KReSz0+pWQqqH2UolVfeWQb9ZEINb9K/qVD5p
1VoF9SfQRNi3mImN4ls8leRsRM1Ych6EuqKAT9HotUsg302tUTq9ziQBbS9zayJD
xky9QoVTYv5xqrMZR3FrO56snQMgtWzpOLWSxtR0dq6lToa1TVr9x36iBaO1KVTg
QWySFc18V3wQIOO4dkaTue77/JLIYdrjqjLAmj2eHabsN1MelmXosbkxoMDJn0+F
HT5Xqort6PxQvRzZnqbngH07poM2SrwqXmpFlbORLIjOCBlSABtS3TOk0XgjMKXU
u5z4wkQwsAZ8/Luh4jOjIQn9M84MtCUnao4EiMGn8KLCd6v6leh55rAk18j1E0WB
oWfWFt8YapIdrVOrvxSckyrPLmty36OgCYgBOgVb/7dpQZu1boFxKbsaOPOk7961
iesMSgMBklh/FLbl0j/duZl8XeHjrtID6+gTqlqPPUNUhcE0e/BPaPneBBI0Mbzr
0Nu/KBIOugRkbnET0ocT+SCbSn5e7HaPT77UgIS2u4VUO5teGD6lhsgL/Ash6MaX
fJk6KjU6c9dyReEhsRcVzHYQsGfOnYAtkkqxdIld9rwGYGY1NjfBLr7Y/A0hZjcA
o7/+evAXuizXTeYHd2kWEMDxvL7u0t86tm0fsVE1W6SF39uAzm1cRCN/26aDksSH
pAgorCfqw3oSd4vRwxIWHq57TZ3ShvUuLme9d55VWv0VZuSSeIwlYUsrvES2gMGs
LvI2M2pSgwWxgAxDsThreqnFsktxm6CJNLxbAmeaYjA9EgkdpamL5HDpJZVwyqV+
oeKErlERJUQ95XWJ0ba76o1kpBT5XOdG+zXcVB09qU4Q9Xt4e2QPElvv7IKa7yO0
EAEg54izYIKx3GSFuNWf/qXctjKl2JTV0cGyDOS6oTeOSVe2Qmsze59R6ZJnAGku
RVvrhTvhkCMdAnF/L5wevzn+KffMnKl3TcEn8fAN9aPVSJCVPtxWZx0ktQ0HTRMn
BgHvMCjsbBkOeYVVx+W3E5CZ0DZ9oQcFDSnqdz1R2ga6XlVyzaAnrg4/GsU9NRxz
2b9Hox3J1GqDBYz2tN9PLQwM+/N0t94PLZ+wtgL/iv+lago07yFFd8aFNC61N1dx
E3is1tsuNNrvvYpcGg8z6QOPD05mdfViFeD9e3GsxPh977x13fqb2AzA+dY5doUC
1bjKma3uBl1OuchZYfiJQAUzPOZNeTGQdYYf8BrPCWBjqq2XRjl/L0J4tgtOu6Gq
flh2SKnbADckTiNuVRmBXE2MsRhc7m4BUuo9U24eKBJCfEUfqfZeuRAWppWlF8FD
M/8k9vplu6zrynZpg+oFO8uszlpM+oPi14RuSbwEiBqty8DqOxpy8ozv4cDY752J
Pmi1VOD4IEJ3tSjjSKYw3QGmNUamm6LWkcdtLwlc/tMFnFGCOIYRMNQYKFGVySbN
WFLgCyBBkLeq3RqcOQgz4QhjWZM1+zFjTFoM1w8P9eW/leegNHV7J+T4oJh7GOnK
GVwSee+uZNgWAsS1d431dHZJguRH74HUYKalfSXnzHHE2gGfBdmrgwPIN4QfDsWF
HRzmbwHLUoR8m23EueOeP1vbtrPU3xvK2xnFYYZZaVpki1a2JdyrdJt7d/7sU4A/
vhhCZKEcCtwqidSDAx2HIHFOhqhhpYzW2eGO9VEpqDzreeBWawHUO9TgpgQs2rSi
AIPmSyBVqPAhLkl9S3OGpHxpEYndukwiBgHJLgr5lPMWq+Up3Eh4gUFTanqr97Me
c+dt60qyrE7jj8YcEoWhgvHwhvzwlkJzV33RmnbnGonRJYFVYSIZGcD4wRroo3LN
g1UcYxk/YQQks61vxSQ8hhko190D5f0q1u1jgBWAGNo+b47bPyAp40+BA6Okux2M
WZdsH4bi4c/UJhqVJYpwyvdA5yB2QM2DDAbfR6+U9FC4mHLPHMfsWw/rxwja3lPa
R9/t8XzFP3iZosp0CrOXM6gtvMdvKvHeogme/Xksfz/GSzQ4h4TrVhl7S8wkZ7C5
BwpuMBJke4vFZ3wvg9wMdaVTdfkO3FJkxpPecL4jShxxwYrcviyLFb2ZW622ZRu/
0WCTvn9nGH3px5YDdFDtm04GMOP+bEmiziE+hGWPKDaoBt+sbFjCSKv9QaWcgwHk
mEi9nxzy/5xJ/yAUfceX007Ch37TZJjC+Jga+aIJ6ZHbvuku4fEXTdpJ531ceHmg
3uKoYzS3uN+zN8Kno805yDfeIa+CpJumX28YuyUgqv5uwgdj+UtrUSJLBm0/WNpf
SuCYcDBTucPIN9NVrloKD+70S+NDJYJ+5aJyAMkGOjszW62y0B2fZilc3ftA1WPo
sTIN3K9Jmfr8qRohMOoYhjZRULmXHEMR6jH4FfY54GjsfQBVi26eZ/1JCMRt9ktw
8rpBRhAtEeRxKgs+E0svvtdGog9x+5/bZo7C1udSaSNON8bYg5YIrl/gtOvf+aH2
RnNz0YrS7j0gbhiLwVsH+J7scwOMl6pvcthHfbd9kVK5buOJaGmV2wB2oSg/KJIZ
gaoiUysvAwW8I2UQT1+FL93dkPIZe+g9+Ujyr1as9PVyW/t9Hms+G+reet6vq4hP
uWM1xoX8+QMTMrsdgqnemcKI/tkPGpqWSZ0ciCX4k5e+K0kjnYfoVDaQctyL9e4o
gALvzKdfNKzP8U+d09S+LfwXKY7j/0wtANSI+PkSz3HrkwSxS6cAK/MceQvs9DH5
LjRPnu1W0B5TGYjXeEHO6j06xIz0VQWgFskQ620Myo12b+7YxrJFlmNI/xoKIONn
nBQx+duHpC1/PvI2fEqcua8CclgBr6cs1Epr06nePZwACrmKGVplHVHepPjlBYDQ
Jbc4xtU9ODleWVW1SwqLGjyPuQEgrq30GyP5dVmoZtmjgxmEO/wREagxm4dDtd/E
/6l05VrnuUbE9eZvKAYFhtU+bLN+wq3YFr2NUZfcA+BD401o1Nf+qRea5grG7YXj
HHJ7w86OQKwQU3FQXqQ1PmJXnEqXOm5oeiBvko/Zo/tSyASUT7gxQ/iVirhjicWh
2092m2NbqlJSvX+NYMzphV5f4wiH+HodVF49KLhEUtPna0IpSULymMcebUiqX5Yu
EkbIw1SgTRzkwUjSD0DgQPTfkTbVF8w0MSDMlKyWTaID6nw8DBqu2BSBDtc/E6Sm
utxknx0m6EyvMByxdgoreXAzfLxKnoGIYitwX+rlrywx06vlUJOiUyS6IGrYJ6yw
TnasKtWyQ2V+xLrdt+hZmEOgiOCPP1Ddr/f4/rBzCnjNBP8uixrBAyzsZCaqXwk0
oMgmJsjaEbxS+pdfxYmUwwKZ071TAqLO6Vc/c29/ov3mbnPvnT/AlwsR63MIJ5dN
ZaEDvR9/tbxZRNPYZI3L5kFdhZLvQ138sUNBb/hl+CMI3b1luvt3GSsn14JBari1
RKc5eqYS0hm7ATaJ3MkVtwjzPSkP69Kfq/w40qByF07eggcQ4De4Ixz8XtulktEs
IqUYAsFmS1l5a5rMX64z4TKxQobw9NUBh+VR0C36y+mpkcn1tivUvHYKHrvms48M
IrGfKfWwrII9HlUwME6jZ2yCOkZUU5b5KXiPsXgbhl8gMIGuQWQOTlanTcZaQtj9
H0CWnWmBo7vWo53tLhekcfUEZ3389QtzLq4zBRVTJJplPgWIxNuZKsW7xDOzuXwn
ZzAAxg3AGUc2umvfcpNhfK8biLGacBGcmbm3cPywMPVuXy8t6DGy0imWRb0w4pQf
wQ7ZRFlqb4U55z+JenlosenUhHi0za5Z9Syd2teGuAhGlZtuWExh6UbCipx8djR3
qiEytHR5bq/7QwfmdJGEfuuDO9nOHj4JSgdX/jA8UVwlzvyASAKt4Jbb0OeM5gvD
Qoak2obRWpLR9hh51hu6TVxTJhi8FdYyMUVJI6SFcmlmGPv6BBIqBjSfwCnhRuRM
lK3pQdFq73HBKzqOGYxiaR057Z8K7HWqOPjLoojs2IOapTfmYf1ffYHvst1xm1NA
Oz52cTWLNF4pL08M4UojSI8VszJDx67AeWA5/wxpE95sYRcMbCkSsVE7ZPj5qw+c
31hur24F3ts3ECpqElUMlAH8VeJFVs+HU4B+ldxtQ13fpsHlxHg5hMvyI5GMTMOz
EAl7IX6CIl9oOoq0xkPDB9iXv3/4FnukP3+8VMgBEoPRlbNR7zJTzNQAMsS2xFL6
w1LBKEraOl5HbM4+yrG22v0m3KtA97WGhCGg1X36ZqG0Riw4DQ/b/8S/zDH+uLWQ
oJwk9Qb8H8kOxjiJI7IoeTvCXAefHLPSoPeaJtiCcMEcCfa6q38SM4J6kOIgdFI+
pGGKBlq1IFM5cuHAUT7F0CQXRzsIxu5XUvEgbJ9r8rM4Wbl4qI53nmA0pdqk96e7
Vc3GTO1z7WgTozKIT9OjW0Qx4178M8QTMQ4rxvQpoH27VmkYlX+U4W6UOA86kQX+
zc9ePifsPYDeQS+15O4+n0RWkmEMhqMO3Sdz2ub1BpjSchXhm07pP9AwEHLLMDtx
BMvaplxaWO5yZWyLVioEl7j/xozQbmMEdbNupjzMT08++ZgNknwCgn7U9p/Tav9+
paJt+uaSBzmUpN28LOtE//tetPj9veWDIBjUyGfDc2842JhlDSakGgYYKwpBi+zy
sAU6zfPsqOhnBVuOm0SEV7kg7RdPe6NLUjgA48JXV0zlzsEzvHqYSAzx1bd4xOC0
wdvJO+aes2qy2Q2NFd/bFpIVuPdu+UpR9dhkf2HBqr1w0x7t5DkksaYI9ku+jlyF
ZcwqjOhaaJ0TtgiK0EbKuSYUqzGIq51sV+zb/YvPH/WG/wZfXxTG5+RiQ175+oP3
qsbxwzCIvlSCpoZcP3G5U4kRiby7SoBNImXRzryccpJqIHiRQaaxawPC72N0XAcY
dua2mWmPXiWD9FB4CKkEwG9BBudtj3TIrm6bXWGFF9c53+wHC3CTipWOU/4ywzd0
zycOe6H+Wf1w/7wCHlULN9QrxR+BlMvEJ7fUTgXCrh5IBaac23ZQu3nKEDcCfXHe
TaHM1UUFqEfIZ+Pbc2omvIVjrIP6bi6i9s/JwuIBaVUH94TInHqOeoB5EkDjM90d
zAC0C4ZZzZbSJlqrbcuEyiDu49kQ12RK2h02TGieEaJ9R3tw2xAoKzCe4dc3UhUP
VvIENroMIbtIgC8DVK3wTWuDUAfnFknDizpJVgJVaKSmgmryts1SwvdO/pG1566Q
SyGta9XimgUZUPoOk3JUpstNRIUUUSj7ztIj/HVzIg5RIq/Q3a3WEu+gVJHLgJ7p
k1m4UE8yLXdoV7E2zQSxsQmLlUfv6AlH5m0SBoFKz8HlY60vWwARL5orFCylv6jd
VNoAwu7TzrOkx1+SVUbpdAC3suzgrmbgWr6GGtvhizoqiM6IghByLqTwQTv4WNWJ
CdzDJdw0sto8fow/1ReNlc0TMgII1JubltZwaNNPgAq2fV0Y41B7qNR9QCHpBgfc
cR1rSOd5L9bO/c697hjWaOEnvf6JM1jWB58WjxAFeaFuykVRsKOcxqjmJ9WBnh+2
DTpqvgF8tIsTzdJwC+zrs9H8teD9HmAz+ExRp4SVOLjT2vs+GOlKkMxBXExJ7Tsv
EBDYQ5gK1u1hGILy2XQ6gl9vQQ2p7GoY9FsVv8sfnMzNT7eaKzInKzE+/2/TeFDb
HNNDeJucBvfXmjT4Juw8zdTiW6bvb0DDQQykkXV+2mVMrbYJ9hibaZLoutpmpJG1
ljCFaGq09mKP3pVf0EWjn8OzBjg2S8TiIsuZzbk0+D1AyvKi1Ek30cBCW7zPFHX4
IKkWA/SXVntej7XOWSiQ4LJ6Vh0Q270g5xA6ygMVax7HLE5RJ9XyU+HTGWIwBHFe
l1MK/boqke5J6sTLG+lq4x2UeW1FIo3BBzje6W125wkZFfeRDfenMnXrlKF4ANyI
C6dFcyUXEgsg7M0B0CNNBdKnoI6/ENEPpjwMqNFODjMNERgs3x4ZZBz+/GhK5oYS
ff8CuAedDMhHLrVpMGq0Llu+2UDb/xf00J9aiT5bWwVaPwmpeYZAgWARoJjEz4dU
ymhP8b2KCQc5Kr3aKsofbuSAXxIqIJmLzHSuSM60GY5oGtJpJ6gZWIdrtoWn20fZ
MkNDjtJh0y3kEk/HC7eeOZFhdp2fDKjMetAQiyWfPR0Hv5Msp30uG4JqwVxCNsxx
QfSF3k+ft20JNgGMHLjHhCF0KhRIve8WwHdggVx2KvtyktoN33ZYlAfFvQb+f0Ld
XZTPiOUwp8UNS33+dFWn/hvRw/fn4U3xjAOBFr28n89osGZm6TCICoiCGx/1Hit9
9TgXjPhMDGlOP93dazMfuvVYbo0Lmu5exRuk8xu8I3jXBHQZGk+c/eirJ8zDCaOB
/lbpxSZ8IvDpMRK0cBIgCEPmOYhOeduhahoFns2Uk9Q/1QzOCHbXD4iMk0VFLofM
1pO3Z8plAkw2YNzqRwGBLeoFghUHXwzOn51IdlA+KEGt3MABWS5EXcnM3RoCXiYj
EtJgCuwPrMSSmP25AQiLZDxxhc3h5PEMm+P+8h0OxKRmM24QxRM3k7RBZ82TtP3Z
bcw3hxHofGwitAZtZ32EC0uzmxod785S8jKqIQpGZA09Lbdo5PgATM1OlDa29Phe
0nZT9+qYnrHSi/1a/mb15Vrxo5liaRWhDVomQemLfY0g/JvGf37hDCgZyMM3jWX/
5fmRT88fIjMEEVJfH/3CFVDK0ov+ILmJT2NEsiVMkCwN5yPHHWD1yvdupps57NNP
UWPq/foRU//dQ1H8+ss07ZXHw0+/cvjsGmQCVRtA0I5bW4WWkA2sUBuqGgKyDqse
2oW8NPeW7dYPP4AYZA20TsvAkkM1b74jomBEO2p93JDULYePpOeuJZV85hHwT3jf
Po+iYYZB45xocb8dOACSKQUSWE7g7tkJd9BKfrifx+/i+N9GsRRb36abmglSra43
qckSxf0ZOjkXXCZ8+T4UcGw9ajCdenyZQ47yz0pMzusjgluNE/nT27fhzg0QiTBH
HmOsixdC8HrU6zs/hqYKOVsC9WQYb30bnCc1ugufrwFXqhniIdXt1S4w7HKS/B3N
2en3Er8A1o//WPWvLkDqUjIbtvl+Nq/kiIEfumVyJTBJJhgJ3nvB7kh1PxIM8gS8
F/3+PO0xBKlkYZ0TAj64nNXcLqTBVG1p52quyleznLe6rShXSopxFhTweJ0Ow/oj
H5KDrLtitOdiDx66taZGA9N6bY3Fr9cfOczjqn7eMCSQEC2UwjZjZQyxZvGtWZ+d
aIEdO35FrPUqDYE9qxgkHFdpwqV5hpjklBLV/Ll8FZM/R+RvTLxDx3AEl6goJkiP
ygwMNpCLbtY/ukbtU9CbscoHpnRovtBt2gqCSyxTCleOMV84AdAWaG+flQZKESbT
M8ZGqDArmELOUDFKnyZrjQVO36+4CNswFWmhlU4HQFLMCSyHYXU6ZMAZIMXj8Kz8
KN8O/W7wjQKhcMHDYSnxWL2ql+L8f3qvSQvwZVt1xIPp8SlX3nhjz70K0N2UWO4x
CNXdUbanz6sKd5dWKcKWXZxI9BlTISbybR82ckCmd7NUhURYrEEgWuPLpyYZgmP/
iIXlxWN+YhF3c5ao6AjjcF8jnF6ubU64HDsd4lcGpgMKnSWrQwn9DHq5dPIm4GSC
sb3+wrvrnEIJ16KQVJXoTUyl1uUnezbLpq1K3uePIA6fAhAm+nQ/ORs7UsWnd5fT
I5iiHbtB6m2t1c5BOxBGN8kSmqiISNLgIRjgdj2MixCc0i0Qj968xCIbQXXi0m2g
9WXhIv7oNbB8ybCHjhRCCT/MPN7DbY0URc5FfXUm/GnSIhrp8C6Udl72OW+mCRVD
uIwVvK/HCg7+RCYb0lJ4O92DW3aZ0uMPDJCmejxguQ+lAfjKaAcfDJjEU/rbFlRe
kCi7nDS/8mpbrPdp8EK2ByZnmD6Mc/5hyZ9msCko/ZLWPq5xC5hiMgSCs8wLkiW4
wRBuAj+IlzQrLPN8EDjb/B5E1VxPfE4dLLke1vtLqcCMY8XtlOIUxGSDVMGZovCq
rIxq2ruq92YkVCuKIPItCMoOQIS0dUcDcaWSdgZwi8Mam3+hrigxh3I2rRw/qlL+
zHvePS7zTH85SHJI5gvwJy59gM6l6spYsY5KNputZQtlqXoGhv5BGqzDGIWDDzmf
s9bf4W3KcMiRuUxL4xPreAi8H+bdD4zKVKlqTJzLTPUy72Cy2cxgUJKgXsmZR/4O
MraxoeYXn57q1ywk5BeslMy1MPp5D+GqJvfCT4a2c2ERu9ZrLj8UTgCMQ+4PpQFp
GBhe30uOSrvYTabFAS3MdK0Ibt3ttqGtYVKMoWhNA2/Vja4jLN8bllFeG6tBXoVo
JfRATC0ayIlncpq02ctYGtKGwATZuJ9M6iyxSVFwG7Z4UT9sjlfHb4oSFnNn3TUa
tdnREdLacBvTOpkugy6P9AJfKwunoScb38FRzQPGMfi17WBTmPaBkIdEyUgLjyca
93QcVXTn29YBQQXkNIGQ96c961L+4oEtRlcYw7OAxqhOWx6DgbEgLh/sAw7VpQRQ
Iv7RF3VK1PVUzEQNX9x4uNjRuBGsWYmeETXwlJ1bHWvzN2xJvqWyICyqfV6I+CiT
VdoR9AKZpAkWVJERSJGTst9JrNQ+wOqF36PRyhglR2JrDpm4LPZW/+nlAsNT9LgP
HTdxQmj2IFJ92gsB/VqQUhXimWY9XZQc0jdmte7F5tZ91hPr14ItikFiZozrb9XC
m6t8q5GRo/V5fvmcadAD/VeVcmBuDLwVDzWR1+dcM+4YurnYxj72dLFNoZj73Xmc
xGnGdasR3p+ncrFSC2W40EaAwl9GMfrVmOHUO6r0SsVInfSWi1laxvEJ8Oz95GpS
v4flJk+gqMgiCpR5c4MYsEXzfca586e9+TW1/zdBI1klRFjGE9WUcQ7EEQIlx0G1
VTpZ357YGfqweR3+oNOm7LJwVJbgezPCWCwyuxr/MBWHd5IjaBlXKMb+1irbwcW7
FEOXbvc0/qMSIzZL0a5pxBKZl9Z0Ewek1G1v32tW2j1rbuAsJDnWZYrJPS1dcvSO
zqNtKw6svGjstEf9kzgdG+vfYoe/FwiLyyF1b0LrId/rYpgpFC2mwD16FaHyM/LS
ZqBbXW/YddNGRnh2HxIhOapcliwAlqwB6p2HoHB+SPashRBW/o72g9wHenE92+yP
M4/m3X+KTTPhvZt9wFtV6FYHZKbZnHLHfC7q5pE3/SCWrdc9i0883S5zktvDjOeL
CEnN9JzV11WTm8f0/nhO+ttVlMgKRzujY/NWXAf00idFdlmhUFvwaKuxCZqoUBIj
jdApuR9P1ipeERSizgqBg7Mmr6O18UxCXEh9/OOCF5tAHXvuz2dpTYPY8J7EoiYt
/7zOvoZ+1stFgJmfJSBjidMa3CdhTUnicRG405nOg7TrZKmp+wsAQ7WD8r3dSpsn
StF7rL55wioXROnsQ+Dqe4/UsmbVs/4sgNTfBaRZkOODfgFs15MMU0cFWZ3mS+ib
lGTjJAu8P6LXWUQ9d3ifNcvDNgyT9WUN0DWnYwnVjz5At6wEHlOH730pENe/l9KS
11i1k50apwBoV1Kj/3YJJ/8OJqQweYZCrragYqzdrp3s6ybEFdqMgKXflkTXOtPj
gDRx6nmMmysUCCojWRUp1Mlq/sSaHk+F6bjGuNuqLa5zr25IJIyZ1N+d9pvDzVhb
YM51GRRN/MO9XfSLySTMBR8SjXMm1HV4NBuvSf5V/2Y5Pr2i4GiM4s9badiJ6Vto
7Lvlv406qgOrxd7JjtWgZL4aGc3/E0x9l3ndFhKm54slmLJnT7vYqks1/hsgGai2
qrZO6mECMnqHt/xAFrMtzVhLY7m3/iUq3098hitlIfdWGIIcye2zkqgwAd+0TD9Y
sTv7KsY0p1CCHslQJB8pWQSKr1R012M4NfIHcxptUBWwu+fvu0j7WRPyngUK6jZB
ioJTHrcvurgVSqZaXtS3VOSu5SOdiNSppJsUHs7yPfjcDwSJ6DEstKkubd/t3UFv
ztQFuZ6IvWy84tvMSOkR2uN9hFn9nThQWBGBflm+YOo288k83IaXR5yHpSi59WDi
xKuIsi/JhvAzO39QKrvLj4AopwbMxWvNXOnsTWI8kRRh6eFJhLqV/5UMcuz1gZXX
DT3vThbbklFdA5AgFa6o84oC+0p1T4RXK+TZeBtaZ8AmqqzGWEZnb5N9ii8Pmjfg
zhA664xxj5e4os0aqKGTLNMRilxYx37nzhYqwcWv/JQZIvUf2aFQya3WKkq3jX7P
WbPvM81bPyFx5XfkCqPEFM+VvSrvaZD0JpANmmjULT8FoHrre1wdRsrIh+h2s312
+7fL+WHF5sVpaztjcz0jfLE9e3BESuxRkqMPBARb+lDxPd1JmwPiQoMwfk/r8nS6
mAB6aT07nVSfD5eklZyY3BylPCaBytfPlFS6vAyOovJ5wnVu3hbOefaeCy2NmvSW
LWG/olsHi4hKMXVRmRc0aSuHYQlKMt5YVajN4umfmqjYKpbDSOTWmQ6Z3M8OPERf
ouskh3mnd9ArehBZXl3qLaSPqEv39Mtp96tcZsC5G3Y1DCQNYBttlguV49QG9/aV
DI4xGeuEDR759xlHPJQ6mPu8fQBadRyxSiwQgQlg17u1/IlB0RHKWLWwHH38bDKb
YjClHPgbhd054cl65B4X8v48xrMSuS5dtBZKeDLN+viBhDmqKc/0C24RGJPfEC4Q
Jo9HRGQrvx58chv9F6uDsBvo/kI6ETB0iAmvbAfr/5sryDzBxsIXQ1mfdHO3is/Z
8b+jkF9+U6Xh4Ilxavfc0vWbaph4iFp5qguiowBg3KSou8OKO6AGa//TQTXTnwOR
PyOoSBdbxGsKR8Sinh2N8/IWd3dYbrsnUHskVJ1Vpw4d40YXR3FNg9yaEnr37/wB
Pv94dyU2hw3ypkGh9uC+RKAumqcWhuMRVukUfg300rQ7hRC+Dcv+E0YxoTx6cRBn
9J+xBJJTYNa3qGb55twvYb7+HOmLcyywoHSOwR6WdhM3iAC7tWSZrYnXhmPyUxHV
4jAR20f3+9QP6n3+YlPLG9pK2oDK1jdrlBTSdgE6lDS5rgtHDDKhEdMRq4AZULyO
IxAux0D3v1+BMaLtGr9ra3w8MkGXY9PLRtqtqlG2AZj1LkaJEacaHfB//omwkPw0
pgn0D01l9xvaBQ8BqyLv2c1rKliuzKNWb6ObynYTY+SfEROkUG9nWHoF9gpvPDit
XGD4W86tdaYi/xQavwjCcgPA+COUtm6XPtz7vU9rxZWYivnKdtmeYaQ+s1Rb47ji
cvoaKvelNqphWDLXsR/zkXJdewlddv1hJLNeuib1+7pep1hDky3JXuNDDdb6PqIN
pmuE84m8DKOupnV+r9OUZjYTp2ulc7vHj4uAGeRr17aVTqSqRaDZcqeGbt+zowYN
w8A5jqGkyZ8otdwrwu6kgZrBqZDa0gbXcv/FkbO4rOmuzUSxxUkD4DGks77NyWwP
lF/KqA3LiO1LdK083RDGWsPEH64Xln+lF5Q8lOkA+hY5dZj6pGYneT2GvVQsEgHx
IChXz3PRe5DPyurN99lfRHVRWPhZICkmCBWiFwga++hUWM0H2H6DfnqO4PuAFro/
LEJDwc4C4kr7N5JaAH3wd2stg8kfWdepIHw8ryCcemNvGaTUt3oqNnKmeDwTMYOh
Qsl8fNg0/siQ0yLtYSjYDRFbVkP/0iZSkF+r7ARW2HPexvtDRa0xf0Nnao3UZJr7
+zS6KxkVMtXylMJ9goLdyoZa73ZdVYs8DfKjt7G/gcVHY01l9dsXrCV1K/PlR5yG
5a2nOhlwqsb7dRXF9Iw7JhCGKpdkjuJJ7X3kSXasdxQ15WnNSK1JpL5j/clk9nnI
dxmSxffD3hodaW20K/OAYmSlUliUt4tsr0B0cXEYg+XOwLmLIlwqdks3GeUBPKST
nJ3Ya1D50UVf0XPgF0I+dkvYrbtHJvJc8R092gZjYcbgn4HZayE9+qX3abNk6R3x
8n2fInH+4+MFA6qF1RpsZNNuFT2ddShQcjC6U9hC/9+gz7peSWWn4AfkgZ1bEiQ7
TqXK8mFakg6yhEDCEtKa3Aihuxen25nH5BAtqCq5MwnqZI1/1xQsLs6uO/3SE2sk
IPC5eim7rfRt1sdsyPD0v2mxR5qKCAmz2SppAnmir/qCEPbe3FSFV4NRNeOwjw9T
ocI/yHJ6kMQkL//qlll6D1tQTxbazgwCfWw4EBvYTLIWVZOfufgXk0UFZyrvTMIM
wQyqqrrLmzr6ZRElDXBWy39S8wcSGRfEb34LhYG0kGXNJ5uMzlCVVu48UFcEN9Bk
mzGMc36+xxmDE0UKu2ml2dKY2NI9JAb65SonzhwVzoEDCR/VSVa3iHQevPcNdwm6
5ODYHzA9Z9XXbV2BgYPHZcIysiEdbgCAhWtzW6X41zU55il16riyBFPHm3VNiklx
iupUA3Q4K3KSbV3xwcKQ5Y8mv6OV3r/WoK95Fmxy95h99dL8U7Ro101aHyB1EGkG
xeh4KWzIemGWutV/rbjJ2yLeULt7OGzHVY2JbyYmDKa11Rmw94gOP82e1j+7v0Gy
o4k3Fv81cEaS+u9x+kRaF8GHj4cRuwwZEK0o/hjV8LJKyVBslqFCZChcIQcYPK8z
liiRZMw+FzwO9wrq4t4SivIYEpKlCpZXJv07yRjch5cYNwOwN3cRmTvFX9IxccEA
eGw389JKjcLQUOaQDvp57pgfdSXhB4y7mu7dSzpgLy2DrMiXOIHPfcYLx8HFDCDZ
sl/PkuGIIX/Ob/dTdlDk0UYAyckREaEUE7kmqHqgEofNM2srflb2+6NqPWJnKgQF
Ji5GkRwWOGp3vEi8yQquv9Tt+UkXAKWxYdj95HU33anxOi3y0Eb7NmASeSEDV4n/
YzP2Ng2/jQRr7kqgj+yZrz+nga1CVL1qzWuw9ElouqMp02sNL7jP/vfoxfdFpVpZ
Nl0ffD481Kif0SxtW0hx5hgFiKtLDXELWbg50wjVVGg0G6n3Yt1C5ch3S4iHPczq
MV3A68O6jneViicr2VDWdzFF1UOCoi+0jNWOiQCat+V7bvzt4st6LacYKSVgpFa5
W+2myYUu+PWYvKufZfpE747r7yt+VwgGTFcX89/JwmWRtW4ywyGXVu/h0hZpkkPj
iOWE1QZyVFRq9o2xBA0Sx3z/6RGIXuPuy6mQnQq3zTX+nOjnax2BgqlbOnaRgSe1
wmVBTN0y3oxMOOesbrWDkUkdyzTttOWL7Sq3oXLFej0l8gy4qWmgYOvsSWtuupkT
YnACP7B+27EgDPmcG4+de1cmXnC1UaVFF5Sa3sVgbckwJZYjamWrL5UbvckY5cbX
iDMCf9PG8OyE3g+e172tAvwLlb/tfMFl7o2e/w3/0ga4nRWqky5y9EKmpl9+bj9k
eA+xYwUp2RVfwonyQ9fI0unyxeNvWysePEOzbELA4L4qJ9+tceLDBc/eKzfrvtQL
T9e3CkocyKIACLqkP6GwxvNjb2uBCG9GTjc8bLu4H0L0hUN11P0I5GINWghu0Z9k
rxIldJJBZc22EoxACEOVtlweDVaKWdpoVYpJ77lnZWx/6BM9JrLuc+V0Cg4tKvMX
GjMHt+5zWcm1eSkM3nsS4DILiqizarP4hC2GxK9HeNPcVLLi8rEhSES7qqb5sL9i
D9gfc4rT1AGOnRPr6Ouf42KOyxcBZ1bcOksRd/Y7Ha1ohywlnTB8g8OOXsGInP2g
9ogcx+t56xTrjO4Q2OPLW+aMzFHI7XdqkZ9+v5qbE11uce70p2sOjf7gw678M4JC
uDN7ZeDNiJX40eI7CRtvHSMbRdRuYiTc4gnaYcjfMXfJihMbxrTjmyT4qvhSXmrS
AVuFNYtLSCPN+d91sQCEM+CJMDxClSgT5IjDYNxEqHnsl7En66l+2axW8shh/NLJ
HclfX5xGceJnsHKxBvRdFbQ2w3GU+TEOQkNEKDC/iZe2CEXexpihyWZ4uEHf4R2Y
1LzFwRJc8AbqcxDV+q94UqdTG9WhHGVrHnArU7NdSidIR8fKs9XRS2H8/z09YLHv
am79owDIVnjEHFEdV2wMWadxWotZ+LN29mrDeiAd5z8iumAIsxBfnKhiBOwnUjuA
g74ev3HJ30pySvAqVAm1kAXhnPSvn4pnHHKmbWqtKBUsv4sUOaEej3SlzSeAdkIE
AeUFjNsn3KZI3fLwATXS2AAM1Ic2tzyI+ArxMXqMwXm6xI8C6WpluT6a++F0Sbud
VNLYLIOJ3qwEYR0OenzBYeO1QsCrPG3BygLNtAnHiT3UTPz4t/sz8DGCpIlMTsWi
Yclfn51IowGRxv3ZQCAwkgAt1SCAAf0mDPqEbj5UBbYkgUAamEMNYAaWGrt82uRt
WWICn9V89K/yFzx0VBWRCaiVOHQqpNG7QQSzGmZrZ3qQsoJIEZpEglyyIWfrMA3b
YmsYpxO1QZCFE9rP3ksN1KM07bZQa6eL7PNVv/NdyNdbTN/dTssGXptKWeF6oEwP
HgcixXS2RZwtcD1keFV+y7ch18R0FF4Rcqlyp83jTv/uN0mgwuZs5dzLeLJnW6Px
v8Iay+XOPa1N9qpxSjdT61OkMwTmgzYvXuwwOOWPVqjh1ZgaqpxwoHXwRHJ8TDrq
J+cd+G8ST2NTeNNB0KdRrZMyjseVGiE/Iw1HAlhU3GIG+zLPf1jxRbfyyUflKNnu
7CuhCBdm9PcDBgWhz9nlnGFNbRszqyo7oHSmTbcQkkwVRCz5vauE8Lmd658yLEbz
YStjweP2GKhbdmGM2GtMRbKZWhIo8C52u6hcr3IFsy6vp9TfHR8ddwgyymYbXkjt
wGQhxBUPwOBf/XikEEtvZWZnDbTl0GOJ48lThu+Kj2K7rbMFNx1ZpgmWmrPsV/x2
wk5NbsaH/BfcbdASC/H/WIQwyWUUm6teNqkXoC2YsaH8YlNrBRcJnFs2siWQIpAi
Ze4kzXUD3A++kcaSZh0y5Zu59ath6cjxriME5BndPityKnOkrMyBCetweKQD/wOZ
QR0f+7kghDUI/eqa8Ggq09BFxdit+pY4FVbMamIFJc0G9lcEQEkzncqtpeoyPgti
o+fDMC5RbGYFshM9+rkcLlkGyOy45r745MUpu9kYEUyIlG7eRRUAatGUWomQIDn2
5xjztPxgfd7Cvldfuv6duHyGM0RkRnGF4+MuNeSSB1sq8AV+TXHQ4R6xC1cN1I1Q
fMJhCC7n5IA+tWE5u6Aby7D2ixucuDAuVxsgHJlRLDfqzGjbOYsEK0BSlZaG91PU
xOOhcnIcIQ6sonb3egOoxnXv9H8nJ56XooWPR1x1OxPAM4dtyN/zLhlgZvV0CzVe
C/G5vpEYH7ATSoZIWqvMHkBALQQLTC3HckzILaui6F6u/Dsm4uKj9C98mYvuBfjF
HBdyD9Ds9MAPop02KdBEE+SSpwCIz5Wp8FcIBcn8504PHpGDP1P1rlGHbqGyBLV7
ZTFxGhHrut7d89BVS+j3LZ15U/GDQp9HC086wko15GyEmsY64OAjbcWqHQ6gsABv
38kA52tRJRjifSDz5259vrq1bTEJyDZ2/sjGU2+yMgIbH0R0l1oTU8D45d1O9men
naSdIMKKrlwE8uvkAk8/D1APnFRdC+Izdyi6bfLKVWFgH2gOVCzVZutXmhfNRkZa
nuthBcI0zlxTMuBZF4/OKjfSH5moVfDXSydw8UGRaeSnOmYIMFLIjUnsL04gf7YH
ms4D/UTu/TpXbRG7/xccNjsdH3wiO1mboe09mAO8yNEMXKBu/GI4ZYtTIxWZm3JT
/EVFuS529a/f4kDYv84OTneIrJf4vNSAOeMt8Ic+i4X4oBu9gx7tC7WhnDCeTdee
OS1g/DrV3BCqCSkX9y/L4PJHKhz8obQqzXKUkP7XO/P4SmeWDrRBieClr3kAwcqq
6A6uy7IVSYWne0bMBk7vOMNQZwPJvkGEidbnpfTiJR7ztHs7AQBSelgA4KkJHrhA
ETInu3hMowIMTbl57+gU/vkjAOl/F46oaAXbTgtaQ6/ZovOMNfAOIPfZl7Pq8MsG
uBeLtiMZ0bYB+NCcqWpBBX9b2DWaZ6sf5q+swYwSS84nGm2AHxvKrd0S3ceWd9Ju
wCGkZ74UJkzLbmSigHbofVpV0RSN1+FJYbbIbFq+QZYYTrW/eQte8a6TXXTA937b
pIxspXdKcbUDHDImJu2qBp1kcGyaIFMii+mBaDqzPJt6qFd/w+awqDsKR9d0q+s0
4/eBFnm20VLEXvL+sUZS4WCL2EhiuAWemWclOm238VmokkDYxjTehrQDL6vFOWCA
3Z41N6zIBium/3SosZjBDaggmi4brzEfklmyQUOZEOG/WmSCnwESZfOpIzVGPmTR
KhbykajHS1fER+1S+OJzrDOEFEwAbYoESOPItjOahYlIv0M26fyW9UNTYjDAwyT3
1oKy9XfE3nmlEhsZimgrFbwsl9gsgy0OnKWzv9iKIPGXLzZZcvEedWnQXgKPlnsU
q121y0TOOuMMIUKh0ABCZkmaDDyE5zfEkaNjRUrdkBICzyzkwOkUY7+PYGyZOIzy
S5l27MxSFNhYpCO2kJP3rvylBHisq19wDVrZzy8a5xmWRSmkvLqCZ2lL2mBGUSvX
mNbO47VcuPwafrF8leuak8ikoKXy3wx85U9ceejvggAHb2GW67DcEkqNBLp6RdDu
P5gMdORr1lyss8btMhR7qw1iSHos1TQKeh9lsqpzqS1QazQjnYlIFO5hnRD6c02j
xdZDs0hYPkJ1+GxR4IuHDgUNLx4le6eQBGEfJ3h3sznSQkXC7oyHNWoz1JXLBu90
hgB7Ui/v+JauWSJCiVdvbp16p3Sbww9K4ym7t9/j+7Y1oeobInC8Trp6FhjomoeK
b7CIlLz0cavAAm43DaqDxOCqpdCQIuTif5KW/68qXasH49qqAtcJSDYPXIqe7o9S
6QlAIw1VIM/abm2PkA1LqKEJM42AF/6wyITYvgoIR9DN9f2D5RcF5iOgP0w3PWMT
WXujL/9LWVBmwLbBxFi2TmRgXvcfWZxsvmEhz2ODqdNbPGdA4Kzb6FomXTXrx2e5
+JV8ivyUoSiadobJYy7Yz2yXO/FTkF5mhlxQPdkPxfbDyHuxDSXvokuJYOETNmPA
No6iK4KNOKxmCvmjctv5AL5i/67khexcbEU/B5VIgQ7zr3akFHc19bsyoT5rydO2
7u4PJPwsS09var0oHuKo1H8SsldEsRDrhQ0GoSCbUynzE1KWDDqCN4oHlocykRR5
VDtjcwxVQRXUT8RtAIUH5+ix0CRXOyJ/G8FY3yU8BXHMRoKRNkZMYYJJuyIIgBC1
6HHpo/xM7XtWWuntNLhVzvDSlwbwzeHLSZUitUh0g+Fi8E01ryJtZkoOjDg44h0K
7eEdMygwA3JAvVl6i6yYOWOsfOudu/As5KclWVL8sR0lEcjTWExlUbmVmlU2tyYL
hNPORMod0SIHl0Sfvq81ojJdFrf1pOn63410QtJgQugBNnP+a29r/3BXmShaW8D1
oxJeQj3SoToXZvaWcpKICPvaGnho8JRQmMhna0o3H+g/XIxNRrWKUqr2xtr16g/8
IsZeAKowQK9C8DBOj0UfyoOXg62sfku6ARaffX4NFPTywGRwBjUH+CfU/C6MJeZP
gd8e8z4ClU7/PkJLUi33l5U2udEtzPHP56hIJimXlDH9DYKKRhFqzadMRFlJp1el
lHgYiUuzV8BhGemo5XYxFvjZbOEdbPPWKn6pzxjYji8NlF9egQ6FND2pOXXLtU7l
n5nTovrRXnrR3wi15U8+ZstuAYVNHsqCNW8tKIOmrgj24beEzFRQje9X/pfaXGea
2nK6py/MDYb/E5zTOrJJeOP0Ravj21Abc5WwbgmV1CFJLSoPgC9ZMiZbyLujDFTw
QW7F0kM7h/Vr+RrF8GbMucZX7mh2glwPJ2RMGPf8BFhu1JjEwiCWJsriz0pSZRCp
9j478Hk4J+36RoL3D2XmtUTMUhMcGLAsyZxS3Tp4x6K0LSoTqRih4Re/IjH9aspf
xo/eUGWc9/9s4Uh6NIr4+1SWkLKTp5UKRzhjm7kWsl4Wzh4SddhD5bwI1CrmfdZJ
qoM0ROQbMOcp3UNUAZIkqvO8O3LoZd4k5jFb0NtP6WbglRRdSojepslSKGtlz4xV
D6KIh6mWrvGRU0wS9+BGfQ1P2coZdKB94g3BrxxVvw20lqm2ZGt4FXJSWY5kCFzP
+CmHOCaUatoyZLzhPjDAcXs3VYJDHzOdHNasOXNfwDmHkGDX75XCXlwOuvcEk5SO
fwKSZqwsvr6g3rjFcK/foenZGIfyBSLDgnWNqmkPCuoBjhQfAF8y8NqajGdFSm3N
sfIzB8+tT23EZgtNxaqYmuKn0pKZyZygsRnjxTXtvW/2cO4Ecv6YxbOde03tvt3z
jZ1XbIkz7lwxVFdpGKirslgrJtwzphFPEY4+MLo2ouKRKeajeD6uv8EatZPWczVj
JceVRkMjNcI+0V6mQN7xBjAWdrulToj2YB+nG6fiMk4UG321N3eg0C/c47tazeO1
U6YcIeM+jjnACAKWlppSxBH4zpp+cGCutmt3/hS5bqiD9fUvJiyTJ3A9MbVI17RV
iczRXceHhKA5ivFkif5eRckWxnICl57JppwLvurUZAwgFScMBGuID4BV6r3JK1Q/
388IAjMPRcYVaqUF/J+aOjRS+Cg4h/mZ7IFA9P9CymSfvbK4FdJnhx86MuTCTgj4
xykboMdZeJQ4kcro26CHxMp7uQjsQqOtwwwkxOojLdpmZ7z4/4KHIMPoTI+3gXj5
7UcNrtSBoOoWjIfhi+d22znIG8oCVMsQkyFbhLbWPEum8cNO5BBgubwwd7J+gV4u
3bBhZjcN58W4sK8iJDF+jw+xHQZeFsNTXqYmXWESploZAvm+zBPzco3wQaHwell6
y7OQw4rNZJqzkUwI01EeRyLAEHm25CNk2nB0y/mkVnZRNDsj81IHBxsTBdmvyaJp
HO4ih3ISJbdW1K0Sd3gMJau02yL497RXAL6cf3cCuiP33nKudr/jrOfFDmFbXjH4
8T3IWh5mfrCEE/oDT25sBETqEBtZgQUqQ/gFGARLQ7EenvvwOdPbSoNPU92nJSi/
JEm/JROFjmsmo6Jy9jDCTtOv2JU8rcnHrxXGDkStXJiB3tz1Srl7FEqNeHLzQX3O
FQhYKGZ5KhfPCvjTt8Sce/uS/UQH5eH1P5cpmmnaE1QtXF2KyMsQLC6ttqzcXSGS
AsTIEgF5H9eyhDdYaWbSEK668fKo7hKAVwLSBdlzRbnxaNrZ9pYRRmpvBfeACLJl
xhjyYTzWSVhiCGut4lx22mJey4TNXt5T9JB8xpO9DNxQHavKTetpKivULFKx3UjO
koqVEKENP2lTlRuCYHIFOOYlYZH+TPWVrK0snm9gNrPwM62b+WrYlV33xYPafXlZ
4o88gWHK89Niori3jb4TIjk/kdw4Yo6M9BH7iOI+YBIT4EnuuIo8iJn96Rx8bjI8
sR9ASUHKin+zdItefZDBxU6pRytMNaXRf9FOZSH6gQKrKLSpgR2TEGcW6H6rocOC
/Q4UgHeCFR+RPSqanHbbgSLp+A3D3oguEi4aZZ5gk2ZE/9pGgrF7yxOJX18QsKav
y8RXv/cpJaWLI047KyCwpdIwQyYIKvfkbr5+5rJriaBT5DE2q0IwDVEJQoGSjn2k
8s9Tg/xXCi01Qg7A94QRoG+nYabmyPkKC3Ag+gD+WWQ7sgM9uqi4tf+ja8BKeDiS
LWwCmyWRseyrZFfRoJuHgfC3kR+srA9LpqDR+MvMW0QuhQmyT22D2prqq/t39sjW
ydl3HnwzPwjISKx7tzp3yYEhD1HlqJRjk/PZ4Zxx9+MDpeCij69E2+K2ih1v1lqh
w99dEUuge+ZmUuwDIvRrEdf0H5kofEdGsuwjl4/hGeWh4O2AQWSXGePlXZBigTHo
kQviueItKIdhYXWt8tFsWIFL28Gfny4hBAJzYcVlPZ0KnPoKukBZuTR2KZ9Wv8vd
55vV14+El6ap5xpatbGDedf0EhBjVm7CuuypIc3Rndl96vL8U4GV6yxWrBe2PqRk
tf0zFTGK4fU233O4hvSoNWEUN6I1vqOz0A54a9Ed0OEVufnRfnsY/GYYQPERWEx+
Kp4OSnT0qNo4Y0vN5PrVBXUGF3tVXlHggSbib72dJbSHGsOjdM3Kz05BV/AXd5Jq
OqccPWZUVFzzNQVcBIcwxO1beDOboI+Wi3LnMf5Q7DnZvOlOpg1mNiZHASOu4QBd
KrkioFNg2dU+6RlKST0+K12Nqf1niWZu/LC2dN06X2XCc4bV+n25Atg6mCFRL2Vr
k8wyzkzt4jqLZChDMGvFmUL/W/DRMJvc2323vs4WkHKG0QvmocbuiljSzMCIe/XE
V58PykTiVRDz+AmPGIFrAElon8qYTVwIH6HpGUT/dDih6LUT0iqXhisU2Ne/zsuk
fZZ56HHIhC8sqNlshcX7VqWufph5oJHp/ZCRHAWFwIGMAw/E7Aan0r/OmJ6XM5KR
i1SsKj+8CH/bu/J5Zo+WmzpFMSWytIwyw3kzfjOAGGtQeg34vj8Dgr2Fvyqv3VPH
Qd6SxjHmy2hMavNbA0cSlvYIkeBCksXYQee34qIXxU5cuVZRe10eBwqooiCh3Y/k
yhBctmUNQzehhVbkHuN+wLgD6gf0Bz4CzX92iX1VHDmGa6VgTzRnZBoyQnRLi94N
1eVJi/swwpD2oHYaGvOVlCzvUOWMzC5EcdP1yx7o/rdvrRMlMfHoicYKlA6Yi01k
yJ4dU0Pjh5cXS+dfCW0BBIYpezJcXRmDXTrsEeLRNrJqH1IK8wGJkwO+KxkoOBOC
Tb4sBEEOYweeQ0LrQRMjgmNpSEFkEpUhPVsmPhB1eqYdEbv2yVkra3ZB3Nq3dI+9
U0+Ygz/ERVTr00lJTPNtgR41Y4LC3zPzQ7SYdAJh1+j7odDrabNsY4PoVgg2oYVZ
FE9tLEgKNLYrjGU9t68FDSOf7Y+x9T96b5zZXyuG8M6Tb8OANh8yvCJgA8Sqb34D
YwBMPY4krHUMkLErxq3F08tZ/6ZlDODuqSk2GpVGWUkuDIqD/r4RPtRhx3vqQEfN
qLTHKWq+zLqowm0RsnIW3ALoWRGb1CgdBhvfDcbLxko2sgzHhpQ3GUTv7NgERkVT
o+BS0rmZY5baTGpCLK29RhUOyejjsH3ExO+REGDTGr+BcUwzZzENTHSKD+laVvBa
peCn5ZKXlPimPe65YbrIG6Sdeqw7huIOQIts9x+co+dE66bDhBYZbnIDWLCos8yb
+HTi5bI3sMxhQ9A/v5Iltd8S4EiBZ4aIN+6y3S3XPpA/KNZH3+xDPtyICVjj3Puz
Khor2ZrqmFagTF7AbHw76S29g3bT+4aRHiorU6wHzrYcOaqOJTjVh7aCef7XM/L8
jkLQUcedJuPOCgvLlDICZo5vvQ3YZXkZxxMGjPVHEmFFCUdDCCLQfnSYCzs6bJB/
0rAiAuLX2hED8lKokbq7d6Y299ytcJLH8aUIGvv7ryCoU7GF2vm//E11GiakDNnT
HkDD8yU7Sfq8hUZa4JPSmmzbeOCGW5uagSE90kFJNVNtMTiNlBYM5M1ApXRxtxTm
cBRJ6u5nxjM92N1TQ+yBtD0FTEo8OnU6jnnWVJtRY5+y0EeP0rUQpvUJN+19rtQ+
t/5eevapPgTgLi1XlB6b+2iFx1Gl+QuPGp8tdTaCV4jDGZrFAhAAYpR12gLqg5+W
JlipyBpEZ7sJSB+jfLngTp27tjU+Q3ooRdvOlOuyKLAdBUWj7cZBE2jr/vO7Ga95
pWJNxkPn1hf9jrdV2RcoOSwEMA55VYQBGIzJlqI2i8gtyzV/n0dgUNOl8JJPxQyl
OvNvl792YFtHd8xSA2xSEp0tHy2AEcJKYKhA9v9CbPEEfPLnxa9dJpJI1q2fDwBG
nqmca9g2JkD4C91n1omEWIXodeXhnek5XTe2Ki4g/exEAhQPnCukTt9DQTSPEEeh
EHDH2NCrp6fral9Zsw1/l8pWO/cqg940uwIwPyVRWYGv3c0nVBOqq1E41F7EFE6T
xZbZPaVTvRbzN9EAbiUFjO6+/OcAmAa6QIVuv5R7eLVmgfYkqs50MD/GgMUNezZi
KKPcfi/F1+F89tIw1fxCfJoG8cX9cxW6Fs98fXql+A1revqO/nvRVtRbJd1zCDhN
7QTRU82ownd/E2HSetl0FKZZ8KS3mbPpKtLlSIhz9citNYnOtgZLb/RidGE+ULKm
8Lb4u1e87yqZ4yQmhNwOjKIERxxcWCLwZ+SonpqoqTONR8CAa6Ca+aJokX6tzeW9
Qd3VhHkn82pdi1pXM3eg2yRoN0R+6K2MNbOKDlSeVI7pH9ZVCADVN3TSSnarlJQb
GQ+ndL9KhqB30FxHRhdM5f+kzFOfQCEq83KC344gavU/FZD83mdcJYHZoH1FoTJx
IexAxPgotNfpYQ++7+mjQwcMQHQr/Z9rohe6dO16rRDTpYspcILMsUZkKOS4onRk
`protect END_PROTECTED
