`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ce7eOOhy02j/Q3ZvAyex3Pog794UhjQXcEj92UNMqcEOdPfmKndovGdOe6fDvDRl
Erxkb5+8QKRJe3/G0JNt8FGtXNTLJYo7E2VrkOGzf5XijhHmlzKcK8oyNGKgODf5
1f96g8BgIJt7nQU05do0jVg4bKHZHjLkVyOUTVfK+6FJ5jq2Np1J/3d/lws6AdMf
yDHVOcaya06Cb3l0BmBB2QPcW8ivTzTukNqm4wdJ2vdkSeZWPHXz5z4wUvIbY9Af
op1CqDwKG9v7sQsEHR+dAULBJ38thi8VRXgjA7VC/ZD+hQvgZkeDYG/8Iu8wE00e
aaSOmuHfhEfY7t3HzdhJTt3oXZgqXHe9o7v4BnhOiu1UGmAMd1/l/TZguwEno8yJ
aBhlD9jdux0nf5wCUwcyG56LdpKJyYNu9gLYJ1Y42/Xx4VHiPOm6xC2K8TTXVTE/
7JlcCjoN67uQ1Kd3ZJFqCB3p2YdgS03tReFJGEhf3E5k2iDYLuG0VdcZqUq8Xj6e
E07aaY9Vbs2vjAxTXdyaqKU9CybBK+24ZcdiV92F0a76qBzMpaMeUI6EGsLQ+Dz2
GkrAHIjtLGUxfMQ6JPzH2NaCyFaRtS5Gu1nr9F0X4mFsb1NW+uaOm36+UubJiFGc
ClCVo813ZW8JyWpZTA/t3w==
`protect END_PROTECTED
