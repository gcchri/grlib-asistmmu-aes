`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Yjjg449y+kpO93vbxJ7mUq2zzrXNXsRyCUxRrBSJhnotvZKC/D+wEyG+Lrd5+6B
UhaX+aCbSyeyJ86DH/+MPfD/7y/HyemcWmAQb0vC8yQvH9/L44lNNAIPC+vdeWAY
OfF4H41DtRidUg0j99HckvYDAdXozRbZkUXIOew9mRf7K4tXelB7HS8stfSk4C9U
PyNQLpUpVq1zuI02SiVevxeqwrJ0gXMqdnzbGbf2GL9C2CMezWKPlRhCi5iNa5bM
yfDnfdX6QcgTLcz3XV3cwiWxRirJfszzhHSQ72bJnoxiIDwllzvj1Wht8cgfcrhp
TAG3K/+vW6j6zOi6NOzgvYJgsJr4gs3ZjU/6qXmGxQNQ7mDZHANPGODI+M1DZ4QW
hSTxf04uTbz6Dkhi97uN0j1aEHAy+leu88h5Cym4h1dj/Zhs9rBGxCmtV23HSPNk
q03kEXT8Rzsr3/89ZuKDbVgxIHsggvRHU9RW4v3CreWeBYT/9iYJBL58S3c57xSK
gJtYfN07tJ+5hYQ2U7/iePEqKsM9sNdSoYIvXeLui2n0y/ylmWqkOI5QBy8VdZwJ
3deiNq3b4Yk+UEkrk1wr8fSZxQ8xCGWKwisPWJRSDwaQx7eKCHcR/rfqh3it/LkL
GIowI9X9O+gpGcWfMReqSULjXNzLqkXwqMypwy/ILwtwAYyrodrIaZNDYoBJ7g7Z
R+6DcmvKudWHrJmiX8zNiNL4pVHt46UC12DwEfIR6OAHi94NYfDI17Qq5Av7ovKA
A8ScxuXutUib/MGTS12OvAXrIhDbC105pusLXQw9Zyu7XPYad0yY16+ON3mE3xlb
NtbOtAQwI1GPHhoyDsdJlQ==
`protect END_PROTECTED
