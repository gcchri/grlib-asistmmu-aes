`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
inuuhTY75ChA8/kSgK/o4USfnbiLjAoHHlzArlTx+TZidYjDsPUjFPWO2anSqbkY
4MqGVs6gJUUXuFEc9lqV2P1+tVbWFF6Nb43JaR3plruanCCxBgZ7xE//+qBQWgLz
kvb7lKaN7JQz++61i2M5jLj8br6/DSW0lHCHrBnE+IkjhO5OmuhvTMGMpw59MT3E
giKIVMGhqiJjvGWzt3gTNLPijEwT1QXdsflEvh/4uaWnD1HQi0fnIKeHX5SYFGy/
dLWJc7/DF4WcWNTSovCo19gX6UlWl49TYu5uGuRSSbU/WkMLtcu1TVuBy2upXIB9
`protect END_PROTECTED
