`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4MqrBjBdY4c2XHvbGiSkfbv9+d266njcYZiGZxXNE5XEqLHF4AO6lO+P+avi5JLN
oI7qqHCQfvFAqL+eD3qWQTV4KgxvcntwBP/LUYrVDaDLy3W5tbDCrZfl40DMrxtF
jrFFD+bu3LuANi1tn/Tarx+Iui3JxksPkp2CL3iAy4NWwBydu7rgqVFaySk5abxI
bYlojFuRqPlxEig1gGDY7EcK5expnHnz5q7XaBthfTRxrHNg+A1mfHsjyv7oFBRg
4YTwIIxgO939819YaVzfFB+JHRPcgW8qSqTLK/5ACAaNQC94/j0/g3sHKEIFVK9V
fXTwtcoi8Zhs2EM0nJ5zxk3ABfw9rVsz7FeQm369utfxwrJeJtxUWX5ZnWf1YznP
Fcu1XKEzX1IC9Hx7d6kG1CS9rD6vnHVv5rNY/1NHXAbwUS08+1g7DicNYpf/UGpL
Zi8gsBvhWksStOmAABNwiz0n03T59TRdwaYSN9EKLKwwPNv+DmfOH2zlOFEz/O71
jcXxa7vcFxdPRB6ceIlyj41foVePw1pgiEaPWw9uSZgH16J1frum7J8jtVUOh+8a
zNij2Lp0YV4YHSPzRv5pucmHvJXwv15I4TZCRSlxX7o=
`protect END_PROTECTED
