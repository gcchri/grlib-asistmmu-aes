`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9nmNY2YAVHtO6KLKDtnvmwPMePITnGgnWfnWkV6djmlaYpajxdaEAKEct77ry1Op
vHVKCeyRPblqt3/7lCqoGpGb4lOfVKwIAU8IQUwOaUT6qg6goCwWq7N1kofFKZeG
KrLhcsGF2oTdd6R+FnNHTl/T6Nuq74rqGoTmFjNr0KMajBiKW8Fo33JPRs2sd0WU
8aHWpq7dKK0Gg/7HHk+x5ZrMku4E6t/Zp+6w1fMk4EEI3Guc2hmvPcTQvSwKWZPH
9a4FQHMxco4wW7Wr5BoL04Hl3JA5smykBprzkn4goORUoLLeUYPw0OPmyf9Eg1UJ
gbqXeQ3VT2HRag89LyPGRnR/cU+JkDXfO2aRc6LOXOF4s2ui+NYhIF8ogSbGHNJo
hBbvKLeTqeGSO8RzMXKC8NLOCSmIDZv6nDZNac1NAivzOO+SeYUOVYAt5+2sa1h4
Ok6ibxM09vHxGCxaITT0exGAXFXJZ6XWLel7kSarnVg=
`protect END_PROTECTED
