`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBWyAFutl53EBAA3nw9lqo/H+THV4f91MsJepcPiUsAiVoLXUIXdL7otyG5RHJ4f
LLOSsMn/9XMYB1z2o1LI4oW2zZWmISyadD7x4APXuTBkBo3eN+1t8yxWb0fomH2z
Ee+N+vRcgmG8d1fafnEqR32rPI/Tf0H2ev0LlZPmDW5xLzyWV50ePuEIC0kWKoa2
oQzn7Y8C/FhrDHa+JHpsK97uN+dJVJB6Qu1eEz3kLz/48UQeA6G3UIaLeXW5+Hg/
pgyTTyS9j1fXW2YMtglTpYU6P5cX6hDsZOHw1k7zzwj4PMZOp+eexzJLOu2YJ3AT
qQfJm4WhecP25DxXli4EBrqMylfwdpRHmd7cVQWIw3pRrb8Oqt9BaVCru/+lsRHk
JgggaMZjzpKoGOSjnpfG/4yNeNcxTsh9dE6GSagsH6iwxEzlc/LX2mhaDLE2+EbR
LmVXVpKnocSqxV8SLHyeOf6MhiNSlDIdh+XVUD1naHvuZfECaB9nFb96jD8tBZPh
uKz7VFg5DYdf+g1RkxHMbSvZxhELUVVJBb0kIfd40z5Q5LWcv298H69qaCR7kpqi
mwfPbO54thW4sIXmKN1TVQwAFIQ5S/qdm8A6TVaEapj1LPA+eDnNFF4R7hqFEyhu
7VB7jrOonX37egoYMMvxJMxJefSD+jqkje9dMOvFwkCS0vW+nOvDAAdGtdo+fywx
PRZfqsFt9YwoT7zhxe57XH4io4WPcPQpQ0jeoWA2WulkYrLXqUS4Hdf2MWFY9Taf
Qv9wudaCjPOZibfFylzTCpdQsdDYthawrfm/3R+akF77Pnn56ZY75ARebbrKMKfk
QaxNRs4Lfv1eRFKpa+QdROVPdc9P21WnH7GMHzzkULpzDZKhosMJhtGFYjUKd0S9
O2GNMNWvdy9/inPQbaND6JXLVsbLVqtt3yGjGCS90hoDqK4/PQBaxlv52CCBwtqR
aqAWcZ6cI//yfdE7gZQRubOm4BEBxJG2pqAk9juFtmsmbfUhOOPYosWnRjMhisJu
LUgvvuAKqxSdFbDXonKRFgBun3RDYfDeymdrDAUNLDs4wd+GrNj6J1XCE53MuY2b
SNYAUfDMHbIUIDgLpP6kgW9mkSuaIo8M8OmExSQGft5dqBvZvxgnRIuiWgiL6B4u
oELf8kppGgJTLCrU/h5/y5T5uqUv29ntaQvQfUk/G66mpYqgx2KRgDPSxEmc64F7
q43pAp8tNGTvQW2T0p7t9tDa+MJ6rUBvA9Ln5Wtc0xp+MQL2DZzXjAEo/rAgmVMu
5dySLf58vdVGCwy0tnQuCCTOShQQUTeKZGp82HWWYFX1h0UfBcvuVc0VM4AvCjTb
NQpVfE2s5ASsQbddo90+aqgvkn8Y+F106NCUauBFaPdgIrGASees9pEGOKFSzubE
U4X1/HXFOTJPQi4Siz59/z8XwOGIdgD7LaaDCDZ7A6pkatPOl0/iLe/UKJGNsalK
zacIhTITpLiBxL9LJYNZ3D5QoE6RKpMCZ9WUYf718RrwtoEwmJk2yuTqI58MymJU
3A+SN59nmtVTFrc54bNo/mPjp0aSPbI95jjLnJoha4wdoQxnJhE/bea3i9ZshfYc
wtIUeAVimaQb72WM/H7OuQXh+eod6Rx5JCs8tDyBha4RXmuoclLaRmzGoLvzJRf+
DTF0NcnoChBh4UAJPb02DAb1SxVMTgVrFwmC6XHSMG3Hpwch8/a3q8x7WmHfTAv2
RBJ36FYnL4YsiBlHWxmgOWQVC6z4KuG0IN05QBddbj7MxNewHPR63w4piBegYK5E
7G6lKAw3RhdVl5Wkr9BdjO87njoSw91I9BQvHPB/llva74hQFEGgyxmRsSjXMFZk
`protect END_PROTECTED
