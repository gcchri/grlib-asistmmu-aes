`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7bWmklZbZ9MtkIGDc+ux+yP81pP7JKSc/kk7AgOK5qErJfkH/sIkwsbO8iZkuwAN
DAPeVeBT4Qqna/5Kyx0PvOhQo/Dl5NHBEeqxwyH+7Jkd19q74LyuH/IxLzp57ugP
En1orvWdByjNmalEDxW/XaiQNoZdDS8BUhG/ZhntEiAzVHqdQ36zWHB6pGG44q6H
514uEPfjdw5dOIjA9v1WH/4ylh8nQmfMxGVP7f16P2kT/tJnM0vxu5s8stT10PM4
sgRSYIuq6IeSOjFcCch/Q8ErAG/I5CjOwQhX1lv3W1rzII9SdtuGHQzXrndwyCa0
6TJgejCOf47G8zVDTxmMYvx87Qztv15n9xKkgLjqjtpmvUaf9jRp1mKt8wIlVEQp
z1jv9QTMoHIQh9F83UF2z5TzoXSgqm/ACo5BkfAKHq90Lc3yhne+2Es9XGyhzV7d
V4MOPxSfAnut61rKE/KEFHg2Tmucm7ktX/EKrwA5Rh5nMbuR4kMp3DPsSZYK6ykm
fT+0DZs08aWb5ZNFDF/KU9EEDbAxaIlGqfUQk//QSgKJ2YftqdgdRpDCJ0BKI2d2
NkwApYV3k/apG7AG4OjUW5wCk1MJ1VnG0tZ+qtv2PS2ELECqAlgXIIWI/dBCID34
pZE/JiZ4qSWG3Yq1T4OF93W3fbDHBDCXYLxcP4A2GPBT4+ZQC9krDbyUzLk1pRVX
U+kzOompLfzkxhegRin+TGiEZgFO+dIbRdpKm5u/SybjjBZcXKf9Cs09WCddjcij
nnsld33LmY/pIgFVht1VLBPj/oUZgH1O5NMr2QPe1GnHoFuC/ugERUxnhGBkilLw
RLpth6BmEoavqfBed81nGS841xYCVsVmNN+MqzF3F5LW2tz8HxxgQoEIo/AS8CX5
IK98aaOE06t9JdgvnaMbIS/YX6fsVnEidUTXM4IoGOmtmSZwZji1kTjR0XZgf8l0
+Zb6hKVunp5yiMPw/yQoqAlbS3NMTxMv+WxNiulLWPq2z3R4lFsB6r46/J1sOHvX
pPNiqSWrGzutt4y+RVfXVBabk9D8aHHo4Je/AuHYC7TVKsA6IgHgN7pc65rr/1bY
l/9eNr6GmItXYVLenOzew18paYDt9qrnF1LIg/+v7pAo+55EQLPTbzfJmf5FBm8l
uXWUXSTxd7025x0R0IzFinsL7uaQYNwmdWqAbB43EmqqCnoqGjNmiJlhiezgIPi0
AtAtzgoT+U/nA6dPmN+hETg8cHy9/0eG9b/tKdxV2uxeReuvT3lLyJ+Rhiu4fDNZ
ScGogYEmav1LqKdQr3ORTDndfE4yXzqYAtWCNHdLm6bsGmq8sNoZXv3aIQ4+1fVh
qnSGYytRfQcRKCnvvnge6seKB1NlcJMYFKIpaverPuOfo2t85FPiVPajdNVuTuYt
ctcRPlrIUIvQcRIQbfyDF+b6oVw2wmKuTN/+k/OapMigH7OpGnqe6dhssQG2xOXk
PIEjoAaMTNp/WetWaP58vCG+DWqNPmPVJDrKw8PVC2RHUAVeCb49CETqtrd62ncp
J9r/S5Satkqqn+LoAtfDqajZUqmxFSZkIus2zbQa0c3N4Ij4m+qHWYjDUDUlkFHL
GtLnuPOZx/4gqzfR0DCBo3aG9UQU7qR2qMgPfPFVi56xYrtOCArog07+ejk4ymdU
ZmYndXxEklGnLLw3+zKMthj7rS9PwqhArKOX0Dp9qHlh9assJnd+eUf9ZclaKlxU
6FFz9y00UdeTr4/Dl8aOgn5ABhtdDblRvm2J5nJ0ULxEpqCu1GKX566HtAmEdINW
WhBzS/znHDwKYCYVgCzx2zpzV+PmW1JCnpgsTW9r6lzgJGsA+Rd+cwUOKBknHMXs
0K6XUx3Ntmd3uzaPQ3Z7lg==
`protect END_PROTECTED
