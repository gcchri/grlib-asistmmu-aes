`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mBzjX1ksKNd6rLnJZgH9kYuM2toZqom8KIiY+ZIq0g0c96xSQXVdO0odyNMOS3VL
LDK8hILo1o70vZ5DLL6o9heoFV9+xlMW71eZJJqHztejIlN/vLLTthp8ectYDFj5
EVjswHC0W8mGzlbBFzPGjWUhEHkKnIdu64N+fpaErBO4D5Kr+v98AfyiCZuOpQe9
r/RQVzZ472LD7wrgHkprxzpudH5ISlD9M6VnzV6iU1BAISafeupcWow+AvMqxOe+
d9fjqFBJjR0Y+GKe5L4bhNQV/w+Z5NxRENVPk7zAHuGTfx/92VY0jIK5vLoCX1ob
ZjbPCLVQjojlD89OzUkjhBqBkW8Uf+/OCksp9j+hM8KkuR2Nq8M8yVhEdKFiTBM4
ZRwnE69RLNC070vieOuO7CA6I0KJ6ZHZXL7AYbtvM6e+Ra/F9Cdfk9jtDFE9DFJ9
czV1FG/7ixfbGoaOARGQxmbRu2kgSVWhF9j1VbYCW3TNHHkoYXRyFfNz9sjtL40k
swtl59YvkDddzY0gtA/sqBH294ku+tgJiCfdA4o85GamvOKp8M2tWqsEuZQA7qLX
OAqVjiPMI50snFgRZV9aEW9t0DmOLvP71WZoxxQuu2A3PThD0daxl/6GiiuiEL+m
XQNQw8H/HIEjYUm8gcbGPh2iQwq+b1TIr4dLP7wNWOUhYmD4nXgKtdjYJUqa+yq0
fpbEvvh5VRrHEmeB6GNRAgr0XWnBRIkNEe82GGz27aOjGjnE9niw/Aa23qcpMJ1d
WPjVAOeu1romlbWf8EpBItL0XwzCewxWd6YHHdGTQyFZJWlHK6HfuxplZNvAgV8G
RTZJ+jzOn5bwEGchON+JAFMmwYE6DU+enntb2HrSnN4VRt3Vjg/mm4LTU3n4kJnU
e8Gz0x0c086qxusxbe9PAs320krw1fgCh3HRoW+4d8RB7lCJ5LxVJVC+oQkkcjJp
rNz+KzFQZnQTKJ1JlAIayq/WSziTEGU5vGtZ9KB4wtsln5ywo5sjg1Xs3nBX0V27
UG1ww0Id10vMha3UYYMV8DRsVJPiDhwIrRYFKMAPzbYgIMBf3avw22aSybpyanpQ
qk+NsH4VM82628TUraPxU9W/IrLIZDTRTdGlewG/T3XIY1uTfbWbA+libZbNHQyP
tooBt1Ov4KBZri+MZpLzrMxJ9IJeVm3ZKvG72bZBNls9B/N/sPU6FLzVUY+kOxBh
GVE/ZR16ujyN75+TLzNUL/ScaXHMAsncH639klKUlqz4IqptxF2YZLOwikDCCITy
gGosW24IcU1SX7MijbMoEuh5r9MdMRCdBU4aJMLz2DAV+j1KbkjRn5xVTrMYWW7/
XxorFfwFxPCDhufAnjlIarM1lyJtUPO1VBvC01S4x0I5bzhyKGBwirKXnuozvclg
9cXMEF+xdDKF+4nQC2mEKpcFOFQEOklUI4LbF3sNS9IlJYq0KyKRyhBb08V+zQam
SBon5F2n531mM0ktgM3ukilXhK85pyUSrhFIU+vu3E/ktl9jSSgG8oFbWmJPN48c
9Qg9561/uxcUrbRZ++DIpIfZMnEn9QSEym6kPqJPmZbjEEPKpOHWD36vf/zSoWWC
kRj5X/xqbKpSp8pV8caeMeyM8LfyEVTPOT9N461ywD+y/4x3uFUsWNNABz4xfJbB
slN7/nRNF0BtyrhxlEITLM0ueapJD8OzmivrLkmF1s6cv7ca1GFyQmOLPcJnO3A/
HwPv1cotY7/Xv005CCimu7t21FHPcGMphdB8uHoyC2wWBDpPvf/mF2iG44lOUQ9o
PO1gBvhpLFRlDdhPkNI8JXDFgADvsrQisgVUAnY+V/rH2US++KT4WWhxPGzSV5lx
+Utc3/9kVyVHzDhm5FjQj18vn0I4Qn6ymALt5ffnzy8vD8AJ8SYUfkD2632X6uzT
Ev7wdteXz4DWi8g+Fgg3esk4GX/BZqsCUQsHdh9W3KeGyiucxJstfY9mbwv/xY7k
BzQd3X5xA5y/bF3meUUe/sVau48IV4AAE9F1QoBT+w3Zz08TcDeKDHXB2WNu7g28
m+JkppmKVaxhrr2pIXzD9Oa8issQVUsom8HGKUdFMk1K4lqQD4inkOBZ6GEgE6Nn
rFDJW3zIa95iWZOkn9QGJ+OW4ro8/IVOrqF91XrB4YncH5QLBP/ECmnTa+VcQomk
Tplw46+fk9SO1ct0yH7LZxymGGF6lJkUuknpqzNboWFIja4MuHbxxNZWV2c7GsVO
IrEUTf6XT14Z0HxPWRpyMfGayMrPj2+qWfpFXi8xAE1yoORVHT7ZcRU85e/OXa1l
s/7Ybs8D8hDLvFezYgpNy9yq73msEXDWGNG5QwjERARG0x9Ik+kWO72ktwvEOOjt
nydcXVRvRDdLu4/be5QxFcZklPOho68hiKUMq6pfM+U6x76mc/gSSujlbF+qtS8Q
luH64QLtyxnKLdJDo+B7iNJdTJH7FdOA+5y3/2WycHdLl3FsUniU/wQkvO/0BWj5
qsb7KztlLvbu7ildUNlbz0Lrrf+i1yqVCb7kE97aLfPJIUI0fJkjjrU8O7u5udxN
tfc+o9PRXBt4KvtJH89VArgvb5PPCcQ3hmwCoYDlCdfDKjMLZ6eU3eauhXYzhBAr
A3C6LFReFp51Bi+UHk29PZaUZzcQtKmhSn8SA6CNvZ2Z0SnRNS3k7LWqe6bykHnR
l47rITXW9LMAtgNv57IbKP4M3JovH9e5NGJ1NtVuAoLfoYihbEua6QqN+wBf7bxl
47fInFtxSzXkPSFnnlrBiLpnPohaFaSCJOIA+Uv2XCiBPxfJxv6FQiyGpX4nWBzB
sC2o8sDkjQCICwgsb0kr3e9tUZdNRmP9fnKnE3q4jNbs+D21dnM24qbV+JoI1X9f
mQ8qTV7L+HYSLS0vjf3Id7cn8EE0D2HacniUfnu/AVYoVWshLbzjA4O5G3au4keO
fjscomIwKR4BfLmAA/Xh2BHw+lbZ8k4M9H1hI4qDJUxMSi2FRWuAAuHSsQF7Q0tp
P6+zJQAVewfps8gTV76XoqepAds0cXCfJo5ACFD/vUH8Py9NhKxkGrmf9EO7zp5d
nu3aakzbjlIZxlFdGCnG+RDvUaPiMBZQxehLhSwtfWukHlqlBnPZsqhJBKaMDRhd
esybzdo+5LvxtKFpFOQRZl3JLLaYByoMRrprxmcaqQ90lV4BF+di3el64kQxdlxn
+rCWXhPqB3YUgg7WLmgXULJKMLmgbct7zOz3zFS2Qfi9t0stIU5krMeUTuVb3NPF
gBQtLVSzwbxU2ekjie86vtowtJRpHYBUZyZm0ddFUxWRwKiBl4vhdY9AoUDY8KSg
qC5mryLqrQ3ygGbStoU13ql+7tKgPg9YE0nSB0YIBMaO43UHAQUeffgtKSuncobu
po3+MzG02fVGM2PwUKSmuH/qZgCaFWzfHzcvTLlpnfhGzKvwV9RXnhc8uWoARHu9
scfVYZNmg3Cct6a3PSEiPtvwn+SvvW4i6zqBoGNDDc0oFTsyBhxaB9SQLelKfgLB
MS1lRe6Rs5NYLLh4BCaiNsorzCmkyVGTUUpoMe6fSh8gyV2YQfelIgZ4DgOIsnr6
KVdaqHr8PGXfhS0fhqegUcFR9078laKZJrVwqnOPF9VJFCeVWmgN/TOuPbZ/i3+x
iE0KPjuNbDRrshnxW0E/k25dqS2HOr18bncv+0qgbCs36urM1i5koEgh5eXmfulm
xVBX59xCi7+OllngnhmJEHcNMx54ZxtF9g8UomjyT21yfF1ZsPNW3h7CwTzMauWZ
/a6ghzaexepp2+hilFyqseiwQRj70xxFP/kvE2gWdWD6yJHgv6YO4UYYdPYQordJ
27jiwIKpACgs5m/mAN4TVYV+O1hQF+IgSWe7gbM9/hqApqL9/1qAP/Ac2Ff1gz9Z
sa6xIBAP5rQ0XFY0enIUg10Lo/LqKiO8LdmIyn3lr2G2ISdiYM9+8lFwcgnFRu9i
Lft6T+/eZ4h+Sj9V7kHenOsKeYU6Eml/6trP8EjNW1cO/xoP8dHpxwwWX/4mcPUP
r9KFelgNGcqdxrvdlGmfhsAQ7LPksQl3N1qQYWeWXIcMv9iEbQ4V8Yxco7Ez3X9h
GlURjem6AsFAN4TqQFvt7dxFEC78tRVfnS0aDjqpYfCQAGzGDT5H50ZDashRnApX
bFdZbtAQ38ujv8w8noLGHeZPLW/WOmeTaBLFCEBh05jtndCBMxdZG+bU8w1Az7Hi
nF7T9hXODtWCzpe69xIFdtngZFNdseFkImSbMAmRfURnPkVQQ/lTPsg2EOZGFm0v
L2R1hD8AOnHecnUoYwKc+W5wiNsfi8/fm33As9qrfDBEal9c8oe84bFhKAtQ9w42
e/nzcCm1zAiUlHHHfHiiBH9zpjny75/5s1+OGEnAcEOxlJiEuKFK31eLNh6BLwAe
gg6so2kpduOh+k9Xf2s61Q42886jvoI59QClWx1nvbB9s3WWScvOWaBrowChIi0H
S66afyG0Asn+ILAI3NUjsRCnwdzGT1YtME/5rp7J1N2T+mGcOmJtRnWS4uSvXW9E
sFwLU+x+7PLQP1Ew2xA6/baF+f8ZEphFR4DlhztEmK7NGoF8/rL4RE2m5zUiDe3f
/W+h8V5AWrJhuieRwJMo4kgTPkCCvwXnejd5ZXW2NhLNU0/zzmH96beZ89NbehU8
FSjFAD/07mdRb+pe77b4QPpERufL25EbSPUqXjpHiDG/Iw7+4GNQXJh2S0VFal9e
4VJE5OHXV1npk6qmZmaZaXFPmVS+gotEav24a3okaEjA8a6AGWK/ZuahfeMbb8Dp
LBwGQ1jNIyy6bxEXTrylzb/q/VFKHaNS7Kpl7L0bcueORg8u6PbGxT2QNH8Zcn83
+TlQq2eptRj6PwVblRh4W84ragT6SU6eQUXN1bZJIIu6HUTaD7Mc8JAAAGKWaYZs
Fp2t6Pp86DssGHm7z7Vs6CwCphkJM9/fhbK9a1P42yyM5SED9mcReUgmaOsejzBz
JAJhxJ5xSAWqvu6tzm7rHFaovoqcWx90nHzR9xrreErMWhGjpDV9I2ARTwEwBDte
Wnj+uc7fKY9IQD+ueXuNiKXqONRDE8c/LVDpp/Y6LqtDiINNiaX+i+ajQvvwA690
vDwEdnshRshFL+eAgtmZJcUPFGFf0Ur596lmCpsnemfrEPqYDNkPTPsC4o68Drjp
oN5AI9fiBGb0qiURatuTin2v6djVH1aHGQwjeJOoj8qFOax3axBmHBBkhbTI4PSB
fTrcrv30fcPgLgFtN+7KJCmebwn931157eOLZpw8bcTOqO/6jWbJlTQeog4OHSiX
jkAFM8uHmD0qoPRz70CH3PaN3Oj5I1VdHF/4uaxbNEVOmpfkNRIAD3JjuIonQk8P
WqTDG3ht9Q6cf9/ci7K44Si3wbpzth2RNAacqsoZOfUytTTBdL4Oe3lGRWfqcWi2
rRprkgB8baIqhGSzi9tzpD+KJc+bYG4QG6lqPBDjKASx5I6rLESA9Z9BhkFCqMkl
V+oWti8tY07EB5+0SP4ExHkuCmX9QEgr/l9OD1O/uah5k/SV6nHtaI0Sudd0UKFl
/f41rKx1c9xhxY8xVomOqDOnFN9EJV5C5Eg8pdFQz7I8AXD3nXhbqWqRdy2e28Nd
VGctMRSWo895SvcOuthQ79D1NOuWkuTS+c6cZFUfJeMAANT8ZiR/MxzaZF6npFih
NePF0rc0q0t19B0rXMBr1Mt2ZyXUrL9fNNDWYYkUSCqJzuER3Vc93VMeYV8joIn2
aDGnJ/FVox/tOoriV084QdGkMzu+Ijx09h9Oj4zIJzG/vyUiCjW9nFgPfNnz0SWH
4JwCjkAhYXzUCvZ46iCBWbREPPHDx53bfsVp9LDJLCDYJrccvt4VmF3IyPTcgBcA
eoVER+lsUoxc8TaA6E+BW1wjSggzPljxLfgxlMczjMMLtLJH/8yQTvBrrY9EFiwM
+sdGChd1DL0aPDZzbEtu9V5EjREmCNflbzmoLavh/oEjTEEoxUO3nUThhsnodcxz
ZRertTuvCRyVR5xksOyPKaV+RJqTaaBlkFLsOZLAw+NogwBiz8yjy+aGeodUyq4d
bYZp8BbRHg29dOsvxosfuUptXXuWZWlYHKhCNVTF+eNQ6nCtPKtcLOCjh+WOCimb
2r0WYZocXlsOSf0OB+43bZZ1frPEgrtirTE7Qa7+HonCxlHmt1Vv/KDgbmAt2De1
YNpPBID/9LC6tYZozTm07mXo2YbzxBIsgXYkFb1Gq8JhntSINoNHC64J8hCCWhir
JgVa3Qm6pXKGObb76W+SCTyvioQGKrGdyNvPmJlRsofgfSsYvGUIkzmorNT9Lq08
4ycA2GJqJtjkI4qCuYlm39Ae46j/yOXUR8M4UajvCvS4Pm7QMxhkC3UxBOZL8Txx
wiYVCMK+RnSfmjZcKfgqixkv+4s2eNOPxbrJZYhwNhSWBI3QpP+l4GXRih8bAUFT
9ufmOt+ejDd8wR906QHvPdoi2CF8OqW5Mthg0tirV3tENZOzIcNe7PJKj7o1huSR
I9t49A5/1GoIfbhB34P3yUk3+g6JJ7UxE8onoJgp8pvpXh3XS+gp4+JizQfxXVsZ
9b+Q9MzAWgj+EpTjursjV3Jp27ZvX9gA4X3ysDys8Pt0/rxASuJ201ntX719JX7H
FB2Z6oDX/EiB0aprSVzTRbFdwo5Sy5xCHW62yphPragYanLJVRCXnpSluoH4tB0V
U0U45/J62UR1Mq9ThqKvwd8vBmJwOa1l/GocPBAyPntQgPfle39qzyJTGrmI0MWf
WHNHXaWYO6hYvwXAvbqJobUa8vGVutgXtcjsHg5kSo7IzDK4Bm6Kptlp0sEgN6zp
diFPAKdRcuuLR97LmWwN+1pEGmDqwwEo5vRhw1v7axB8R3zgNAluwV7PxkKscK4h
fVIT1OVwzQhvD4U3LxggPr9p9QVdtHTL19dmBEf7p9luM1+mXgpSQUW6YcAJeyUy
Bi0z15gCh+K9sAGhD6snGl2Z2+bXv0I72qGUTvtrJWDR2hfyp4JnvAGFTS00hTvk
I4tGISDA0Ob8VVphXkwPml+YVWzZQhfOwtCGWxCegoPib77WTg5hX4eg0EERHEi4
0VTm7OG6XLtNGi4QyapV8fDg8ImZC+j0OARBm2jDekRXpdUqlkV4R19lF3UgJ9bM
28+Zsdhvhcg4ttNAAQzFLUuIrwND0RL3C7AlpA4EuAAFa+KWJxXmqoO/HtfuIAfD
gqdt4/YRlt5frb6e7gJX0io4RpUDp2MyE72d7aZpjHbFJ4gtOJLcO50vr5yihFPA
NvK9fbmsF5A01lJPx9A8T6QE0A97cwd1D5kGs580ho1W39cBdhfGUQxezHbo+d6h
0yt+AhJA7Slpx7Xnb24J/2NCvcYGXbD3mLoXnjVId5+gkIf3Dr9kd8X3sOEgx5EV
hiyxDQxV6VPW65lq4tfjdwIPrP4VtXTkHy161pMp3Km0ParOmajFt8EKV0pES51J
`protect END_PROTECTED
