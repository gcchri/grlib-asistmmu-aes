`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BS7G2g3Xhkeo0Culxw9HURaS1dGwuvuPnqX3Plgxd5080aPaxwbqhCipgQewjjIi
0Dzn2o8+EyD/c0waBlvESTD9S2w3VUPjNBKyTA3o0lqAwvp+V+4qG0khOIw8qAk0
b0Dcdbs4CXRuVclvgzN36vikNHV+d73bc196RsRZ6Lve1PBsG+2LTLqVv1VWmcpX
5MTHYHLLzuIGKuGSGwkbfOUcy8SRloZBjoWXXFlgkwJNLPmhfGk3M7XA/PMWPHp6
btOwk8xKR4fpHuFEEgxnnaUBzRBApfx0p696fwABP+nyMNFQSeHPcaXMJreApS0j
z1+0LEJThQnrY7ZeutIakQgoKqfRPv4FZjWexB/b1R/emzlrctxMmFdXxWcFk4ok
Dom4kWPyRloHf+vt7D8LbBi/dKE3hVqQFbxIMqm4eIxajTd0rZY8lTWFgtSZ6w+1
9DbUoH5arCcEYZtF6tymrg==
`protect END_PROTECTED
