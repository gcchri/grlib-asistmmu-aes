`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/FGCGVOCf7F+KsVe+VVuhv37gLd8DrHtG7nRfVkr+U6krs+tZtaWiWJa5x/mI3j
d3VolZVg6dhKcSJjmz9oYPEE4xqSYdWXQW6bTvkdLKlHiVX3VMkCwEtmYZ5ZWO2x
10D+7Uuw7zZWuN9xuHRa1EVp3KWm4NcxAqTGP8b9v5rPWu+AEnG4swlAcCxTFSMe
BiKi7X5yRz3hXGx8u/QsyWPFzTdZNCxayaRCrIC2gXCRgYGRJzsLTlVYTg2W/K1S
iuHvD+NLn8UBKw0niV0LwRmI8G+8r/uP6SuxdJ9xV45ShnrcwBaHhNlfyfIQKkfL
pqS1zH5V1ql/EnvLdOLot55cpPd59vhiwC4sMtCiDBu17dDxoNuDtQpvU8T04dJj
B0fWowDCLKxHraRiL4MZu/LBfcJ9MQds2u92zvaXLu5VYxY+YM+lc8KCoOTYOA2N
R2XpEN9LjMKCTHoTYDqhV1N0QnblWbfwFOmUJhRfG8tUa5/YLl1ykVtInFFOcikl
b5u+EN9aXqh6/tpqk7Dh4vV+q2jM8MJdM+RPBTMSZB6qvUZAdBuP88GbEzXcKUP5
AI76z+lCzeBJnDoe3UqQ96FwbRUp2xtgZ6TkehgpNGvw4VxhOFvOyE2ozeuvWGoR
pGZbrvz+m3Fn3mt6Y3hsdFOKScEWquKCHtnkWjc0zUFFqMJh0jDv5VN+dLw8Dacz
SCbtllNpS+cCi6dbBBu2Y7cx5KFsl6VlXw6NmdTXSfWYsz12Sk48OXP1Yy67lgnN
o6qT2j/2njVMvt/gVQYZeQ==
`protect END_PROTECTED
