`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZDb2DAgw9VVdpp18JaP1s+siT188IToIFdSR7yxgxNevrd6j1j34jGSGQSkd7O0O
zGyQ3WFykAil8tG1Ha0o0YA3gQnhD3i50Jzs5ONiZYyTmIkYw8FC+cPHi6oiJZIX
3rJtBy8kJ2exJCuywXzmQ4MSVFD5GoogVs4iD0UBAYgAWBVJDW5Sb20USNREdb+l
T7t7yP83eO8y25gg+g0+Jo8qrnbbgFfkqGW6F6qHpgzFb72WPsjlRwAO0ND+BLAm
2GT1NnRocYMJzdi7//rwk1V9XMx8y6ClXGAupi/AuaROF/aXrDMsbb3ucfTstEGB
A0InSa9fCxdQVrnBtQeRfsuI6AzB6rO5UsTDnrUXGUJ7R8tSiSzy0AZl+h65SQ6i
QW0L/vv3jAC6cylWn/lBh8eVsWjMdofI/MuIcQsIi3OE7PFMSQrTrhDnWIiMDl0g
T+EUpr8qXgfPQKkJCeXqgjMda1Hf8N7Gh7hzKVSEZLKQtR9yNJurfKLJ69U/CNKW
`protect END_PROTECTED
