`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rM4UR2qt7hS09L8K7cvLlTMnOmmnfDdPpYxN58wWuiqFY3+kjVIDbjACRlIuDMPl
3dr0+QGQ1zmyS8jOfLErhoL9EKFxJi7mZltMELjFUQVeO6vVAeAP5TuD+PX7gYlL
uM9GSPPJUz/aV+Qbmgi3fYC69YrgY6kSuuwDskQZMpghLkUs2X14bFpqD4wZlaZK
+PFLj8zYI20kbSTpHzDlehnc2B5EkE0wi13j/VGjYUXmIqbmvF/UH9F3SuIzpwTd
D77pCUzLwx61rPG8aQo5Krj6Rx4ZOkiXrXGjsqk+dts48alQ86szBt58qfDrZvl6
wkC8aIKYNgR0tNyYBz0GRcb94RAU80eEcxez1g/tYxokDHBn1iab9B5rUt0GACob
bHZdAx0QiPaCgukVnCfVWSCJfHcM4xj092UB4jdLhgcrCy70MX8LuprR3w0ixAq/
7XIi1ayH9NK82mjFGoBzVjCtbMoHapLRe+FZJ+or5BU8MaC2T0cqLd5jWhZh1r4M
8vjdnBdNQZQqbJO67XrQ90Uic9yiQiJTOrslbQlYB0nqXQjjG8wQOSE5NIdLIeUt
0r28elYCMj2scZdm13sHxxMpstXqktQnYXPW+zSczqo=
`protect END_PROTECTED
