`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BIHmYSIWsxZio/TEUmiHlbsLL1WwiD7CcN79Wcqh2bCOi3SEXBTnUjclI8ZXEZ3x
VPDShiwz52gEokGkSB0akiBfhM4wytAccg70fGot5u3FCEV8McIHWuRBJ3aC/oMb
q98miMXQ9v2e/Br8eeX004PR6xBE+lXO4jGqbmKBlHCH/1qcOh5c1W+3e+DZqUSO
mdZ7wSTZU0LYfIsAhE/9qF4GrV69Lskhw3KYbzCD59Y+pIi+XsXcH/3SYruhM8dW
m0tOWO0HBnR6hc4knna27AlP3W725GAmnPcK9FSh0LZ/QfJdEZI5oEJcG1Sl8qqt
PMANWtT/ndMlUVW2dqJuCCqQ4qB8dU3EvPpRjBa+5HjRJz7p/lMVItCXbL7U1YIq
Te+TKhypE2SFg0Le5PBhoQ==
`protect END_PROTECTED
