`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+BkP/E5eUtaOAvLJsrtnOLLLPm63mY6z/LgxLKR9IBsvq5/z3Lc4xlPOQY912Ed
wYjDpjovWbKKDQHhyB+arrppIvO4OO/4BRHpC6qwFeKn900M9kQD/+2+Vhzej5l9
0X0BlE3soeWI7wgHan61UXySi+d0TiXi23eSVTOZMzWL0zkRzOcng7RSAERoISLQ
0za5es+gu7WM1bbvtQ/Di0aULFLrqlZhlMy5KQeVQuGFQdFYElJNoE5e4DzNJVfe
WULiFHxaLf4X2EPL1avC9FZvPtil8/FjtMWrzy0cvPdocjQOhQ6769kzOnwbM3Rx
NsRIq5QcHBAWUxZAxu86smlfZ7bS0JS3Dd+mPRKmvdE=
`protect END_PROTECTED
