`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0kfOEjfjUQoUzMoJtbNKHveeTPCcu7Xr79DRa7WGed5e9sE4TM7iaTEf+WTA5k5i
M9pvGN4wnOBEpxuMnZqQ7nCUV+AjxPXzk8PWefFEHYoAuGkuOn3/DxK3nhfh4QIC
VcAxWVD4yDz1+acz9jVK4PuZpekUkcNgk4t6h9/m5esF24KG7VE6nVShF3KFntwW
8THV/bgjuwB4ohM/iCba5AIFAMVvlscKQtlgVo/i3T8+cAC1HyK+15kmQlUaMiaT
772nghe9anncY73+H0th7NqzJOv/fK7E5Uju66W9LYetrz4Ta07g/Hb94duBu6wk
obKklnHfaYXE34DeX2TMkQ==
`protect END_PROTECTED
