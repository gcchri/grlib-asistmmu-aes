`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iIvdpJwlGiV7y3QR/QX8qp9G58jr5SqGKx/qcOl64Bg66lDSZTIsRVANk0HwlUZs
Q2bnMuiyO+n3/rHeSxYtdpYr8k28slUm2qM8GjOiM66PHZG9+b5FOIDgIKQJb2np
G64MNoENxl/00n47XwXtEo0GZ4R0FzuLDOh5Ug2KcnfpdR2wW0k+muCgS0LuhzkH
F5ObQTsaxRJG3CXlVa1aa1ENOW6Dwr3vYA5hyCFV49JPr4DDE5H11RfPvHd5pY2i
MfDQhZzfvRRaT5PbijmkwkQNxkKNJy6A67vnoqVop6ZKu+zc2F1wp75upbLK4ice
Z6QzpNog3AWblB5oYEW7oA==
`protect END_PROTECTED
