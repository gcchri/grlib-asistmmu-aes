`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5VCA8fTb5qmmnplltYNv+QIldTG021c2jZtYO4hGniTO/Je3lRQQfpwiGw/dl4e
D2b7gRNzDYGyLkQ3H0X0KTE4xCQlzvR7K94RKBr/1wzRqZtgBp6YwWwGEILbSsOt
kM1B7XFdDmdXCxWuSc+VryDa+eDSTSKkyWN/DO0gdaYSL6FtY4HxaHHAC1ezDEO+
Zl9ryGp75/QwJPY2Xv8dqdfYPYtDukLg5lKB509RtIBTvwOU8it9lyP7W9GNMA+1
scI8z6SmFB5OXt8SXHVuGWn+RHUKws3aUIVPe3UyE88VzeFMWFOIVAe3RrkQ94AN
CFtKLBpxG54yuXqcsoD9k701uPAFjeAw/pDJ1vxK/O9to+kccftgrLcIUseZ3g10
GitYtqq1wyB7jlOQmZV/8A==
`protect END_PROTECTED
