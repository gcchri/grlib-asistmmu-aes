`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OvLl0cRIs5FFNon7bi5LxikujVPK8aoA4eH5OOKiv6qnLaZXeKduBxYeXaS+qcYo
nYAJ5iHH1/cpDqIt4sK6OO9faIRBGwLnsJZ++E4bYnLoBOTcHXKsjZpYi6p7mANi
wN1AG4u5ScZZZGo8NwZwj6FCSqRztoHZYduixAFToCPXcJPSitZ4mPrZ9r2/93Ex
9L6BuSveGOisERqAfFIz4v/QN9NS796UkE2+4zxplrYd5OasDH4oRoz2tH25tv31
ceM/B4DbHPl3uq9EURIaOof8SiBBYIqX6BI2sG6NYDKuB7QD7kP9dpJH4SvKeDaL
uljl+H/1GJHUGmxs/xGTqQ==
`protect END_PROTECTED
