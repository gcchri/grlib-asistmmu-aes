`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xoCwHU3OlgQzzOU75C0Nvx0UVL1DuAkf9bg5cmLkudBoVBNqu6wnE26A1iMug3Pm
qSa3ll7N1fvjGBaStF/1Tw4PPssBHtwFxr1yBmr0CdVoKD5aOUTRpC1DOjMcQtuU
M8XXTUBKKmZ9dU+SZm5ofJuwd2jXeGhaU1rznHl2Wz7BP85XYGGnPc2ffXtVF/05
GyY0sdviILZHPqrsqGj64FrKqvSWSKeTR6CwEuJJtv0kN6uZeMKHkCATLDeGMGEn
mdfxWSbes8B36UxvsqiHtxzZqi2tC8PU+UPCqV3OXse9NMM8hn833FECYn86VvIw
wMGiogurtZe09tvfXKuDRw==
`protect END_PROTECTED
