`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nh7xby5RpvW+kf+jgJfLaBNZWSELhX2cab6QEWdZWTGBI/TEjzxLFa0D/srHub6g
sXNBmnVarr0rBJF8awu3iCVIoyBiVt/OZ48cgmmbSdqA1TAeLpbT25AP3/8u1iWx
KnUF7mrERi0pa7KTZ2sZOPAl+bizLCAoOO/XSa3Ozjrx5fIGeCvSw8lm4JqngiVT
U/pqExVKZYFohpazK4GkPFrAbEWesqhNGt/4yB1oN0gVpdlFHurH4C5jNuqaSDuZ
eDs2we/3GkSkwaNDr7pvhbN0BT3EeroZeHvnVnXgoPi9g9nETtv4oQox6sGdlCty
qzABVnea6I54lgg3hq9qyeQST7+xxxQtRuJxMnynrqRUZUASNGTcd7kkp064Ms3U
/Pjp+wPEuTshQZ9JmxNplMY/vD5hFXYrveTHyvGborJ7xqL+ylqiFj1IF7ttqgUt
KrVJpzqGily2FnXLsjuf6C3REq6O/AWQMTM+/Umke/f9ZfDMI7GhdKmgktA0a0P0
+DDtiyAMVZMam95/xiifXEy3LLGbOO9XN3V9czFX0c5/6ChE8gb7MASyKXFyK8lM
9370HzC+YuDAxKqXGcBHaxhuRNqOpmOa/XiV4Vv2e0JqYPS2HV677waK2YDHPJeN
7ULd1Rd6Byld1IZOb5dtE5l7WZhPs2T52uFMZN+ONpxm0HS304UNzKkMWI7oXMgo
/Vlo/GsgcvWfiC61xe6Jv0GFBDcNXjh5N3c/hxemGKb5n0VManWgGxF8D2yEFCfY
SmWDQhTlFHOgpMldt6/8I2dMEI7He0JA3DcePXcPJHkveULHE6CLpFKGd1pyuMS/
lTR/sCA7No/Zr7ByAtnGcr1EcNVGVjifI19fowi+JXu93E0oQEl4HsqlGIlui5MO
KTFNgWJBPKHnOV6rUp+/CXONLEyG4L2AhcRMuXOmObY=
`protect END_PROTECTED
