`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEYX8GfoemJpqKNvHH+RqH8jFK9jCcIfm0tjYaLlYCl5IeP6T5sxi1w/ZRSah2oA
4Xb/b/pgxTKTnxxrx33LTHN9gOAj3Tn2Va+IRYZZHbQ3IAgfaO3e1K4rng2NLqJk
Tb+2PvTQ/XoF4HlCEB2gADyLykSvkbGzallVPzF+wGdaRc1yZ6xQFOnGxk4Kobtf
Df+r/SUTBlqjqrKLuHEHXHnFyQ/Nj38zJldQUf1WM5BwiXBmq4X2W6BWxrrv957i
xv/snoSVxd8QCrmRmRtkhh2g0DSLpp/goqRf2XVdURulK2Ua566jc4nLEbT8VD5G
3dM0+rUk8SWmiSVDMejDJA==
`protect END_PROTECTED
