`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Osk9BQZCrOmoLpV1miV7Q2GbGMUlmUPRMiK+1vpXXyn5ZOH/eIVHhxf8KNRNUl0
z6mi6Tk17QLtIejtt0pOZMuUsElQOweCLJpbSjkVADoabqofhj1UBKUD5r7GsHlh
Y2V/r9iVxfX68BBg8ZR1rfDZ6fSJ4r5n6ptow/4FSaekcCZLxdgQzmqeFGB4ml31
qK/JWUoNmISJCvJ4WN1P/S4jvkzWGn4AdwEWz0ILjVuJP940/ZPF0Mq261bXzkRu
xkIBTBU4xnfN/r1lM1W5CxUj4xAOYY9QRlTekBj4Umf+U+TDcqi31yD0HrMmTLdE
s24oeQIfo2Vry1hEIuj7HIXgYNmvSBE5dVwlKs4Pd/4G6WAu4IDTbMW51nkGYU3E
rzML7h4GNUyCi/fKWjdZw8BwI2feqE8OqTWQUTl8lHWcqB9HMD8WN6QninjtMOC7
dskfi2lumW4rgd0Tt+6WZQfnHevdMt+Hlmnn+Hrl+Fm+402BUZS3eH0MYt0HrDx6
yYzfIdI60sfNFfHXY5kX7+oKfmnJqJ+1ReDdJC7GwDnGISHVPU2n4rcblLpTeUO0
NDShNmDDcadcud2h2dYz0w==
`protect END_PROTECTED
