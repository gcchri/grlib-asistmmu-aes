`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iBD94pqBa/LB1gAONuXvZ6hFs1mJxZbzUl0NunAi4/1xCcRq6+yw7L0MhlS4ELs6
V38ysJm5PgUFftO43cdJ+WUMYX3+6qhmo1ENVvJru5+K4QxoxHB7m5awka9dTubl
c1JKY+LvwO7rNqTWXgF3ooDVw+J3XBeIYPBl4aF8NqQuPWieeBhymtW4pZlr6pSR
3Wtb8o9HVdi41uqVfvQh4DfhUPPQfzWCC8eBuF8IHF9v7qU2ggPTtv2CU+Hyaip6
awLcL4pyRwdpW9m4HNDVf6ui6JXHTNudsq5AeLpVp+2BB8RMsrXRmEZBA3KGYi+K
NF8UOmHVfzha9yEQ3uHsYQL0TvZOP7TrWeqwulfsmQPYJosp0RZ6l4QCc1wbe+CF
82FvBlQc3zuXcEt0JXenT1FjXPQ4rUvcLI4qbqZmocyhFdq/scyDX1glw6P4rYpT
EZEOmOSr4xp0Q6ChPuq8AW2/qazg26Y653q6cGqi7pqOCO7BEy/evAwTKFt8PPyt
bzeK1j41hhu2VtVbHxoeZbjirq4OAgIIGmAVv5jmz5kymYOj+K7T+ktoh1/7z7kK
IjwquiT8htlsST3MucR/mA==
`protect END_PROTECTED
