`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWUTvq7bG/0h4oDRicKz/rY1WDmhMdBE4Wdb5+p8MVW0Jcmgm96fO41ZrqSBxRfV
rOTM0aCxLXk69RGrBcXglCy/VU16E5etR+sE7ZZbqPS6ze0zoUPhi1pyOnCTYPij
DZVp4KLLcs3nGqJVklr51hKC6OsX6zaspFhvE+CB5nSWWYwgv9LTXiDoQgVMD20F
p+sv9+AY+RmG6D4nMAxu/oe7zCyHVgCaGtiy+0P0HLMb+p2be6gWG1whmQEDn9Ws
acuBNzsTdZLpzKyfauicCKYsAVsLJXSSw5O811nMc3sxRZV2Oup0pmDMFZQHOV4R
WfJNciJm7uiekZ5NRIZZSpUYkZ+8IXA+bSupc/Gzy4rKTfWECKEar/7A3tETXoIB
XTif/h2usHA9ZraJyNWfB6pR9k6LBTmtmulUu2REEh8=
`protect END_PROTECTED
