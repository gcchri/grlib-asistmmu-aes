`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPZkOTduVws6CeVNfk+k9cd95RRyNck74DKUVcMM7tu7WplFhhhbHQwxkIGNy+xj
2cHoO1Sg/3rjEcdonL1P8C1fZPHK+CyewpXIKt6bTEFYzJTbrmdO7yvDNjv4csAG
s0QsN4Ujdtnrx5BoF/asWl3KAZd9J7NDvumlquKhiCSHyS2gddCavQ405aJiueK5
7DnVzdFNQija2+ss4NHOvSycFsaMZDfFZkX9AXJadLEjYFkxgtB1OnQAqPyHQLSl
oLTtbcLjkNSWQSvGYNPPkq/JK95lDKuSR9hc0LznBAlw6DPOb1ZouYMcavBwYyF5
en4f5A475dBaGBq05xn8rXGGFBNS8pFJibJR1sR07hFa3H73KTwcLqCBK/QH4f2Y
rm7+Evm7hSE/zwg7wtcDqggXthue6u5mfOr0G6EHj3BUvxUwh8R6HlQzkvrpKc6K
+0vqxXtp0zTrLDPNYZA/rkfRt1w6chKulCqvuPWLM3dOXFm1NHv8VKEhGPqhKp9z
NKLYaZlrYlNszwH/cgXXw+qk3HdnOURm74yYNXhrJ7ir/jhyEtw2/RaIVfrI7/1+
1goBArab4HrhccvuEp+C5MrmelEQ+j6UXBtsHv7pmwX+wszgi7hfzXdT6ThYTtzs
`protect END_PROTECTED
