`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JzOQzJgUI/2inyXoHYQSaP7hodvjCkcUFA0LFByAXuQ2hZ+9SpG/vEJ96Bsi+FVf
Nc2lbdc4HY9Mtu1s0EV1QaHDsQUH7SC2rIlCLalGo1KtC9fY5b28VteFD4eOFUsg
UXceuNA1yI00k6h7OVBc9OE7UnhFCZALDUnsniO3M61f6aeJu5XNhdmDi1RMgxD4
jEn+DrKKPr3mrISGIACmFvz93/dmh9SVyBaRKGsI//KPq6g+sKvoWvMDFVcf/EDx
JSb0Qn9bBpXAQPUoldtcC7N3NqHOJIWidSvZGeatifSDJ/HrVvwazIg2fKKNQ6TB
`protect END_PROTECTED
