`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2LZffTJgLPf9sJ/fTtYej2nGRxKsbsoKELlvUDZabHOPTE3LcK82Ls7KAEOtrug
AD4CppMIzZczTFOPTYdSoauqyLojrtDuivjMeBbbW9SzPE4fvhpun1d0gu/vQm2c
py4xecuB6J2dgtYJs+qeLUJYK+sBwzpv6WkEJSE47GA+D8KgaRUEslJoDcy16gte
tFxwAnsUCk+1ChKfQSZPDK/PtsW8yfrB5L0cCcft5TqtKyrqfh6DePwHhF1SiXe/
D0HL1XbQkg48cfTDdc9qhEHwNvn5ZPZFUlwxUMQSVfYCvdYKkN4ku2lPvREYF0xP
0kQF7URnd2HTDBKbQ6oON1waMnLr/9XHans/18tp9gv4wUjtZPB4t6OWFyxp78OS
5C5FOSKf3+QzYq22I7vQ9LJ5Ci7fZLrc5Gx2xqNUxY/CNdac9qB7eDzrofYAo18U
iBoWrzBMr2soyj4jVTiLP3Dbhkao2Zd8+YH9q/ZGb00GOgt4mKj0KFUV9Arf0CPb
vya2MpPoW/c9/Ne48xOWwZInxCIQR40hkeUwmQWMdgWAezz6HIp/otqT5L/FJbXX
vVFn+QY71kwbJJ15zhzwFxm8kZeRBNgJ1NwAJZImbosDXA3GoGElAtHyYSLuFCZT
/BFzgtPDPfwob5Yi+TuKgTpSwNY5KvpsHygzCRSdOfhwMDlyfFmoNQMaoXL9Duch
qYUvMvDVDXTOu22zTLD/PsxKmKBtNWkEG9D/X0CnFFn895+VUZ5DUYZ8qXAmGV3d
Z2FI4Ss1Fa7VNAd7y0hbGCST4FyV/Nr0TXhtw3RJfrw0ttj3+Vkbe1m25tsKGYfF
PH7SiLq1hnQ/sbwLKsHJ7zS7eWfRdREAGsbC1CCgoRq/YiIs7CBtF4ksU6LIBDCn
DLnUhnA86rB7pZkEcnzmVQjgJe9PPs7hS+Ez/PKHM0De4nNpyOBgRZ140ZJfXHXN
/nfokC4VWpOYL0vm4DTRLFINoSYG3CYhEluD8eIWNCtBT2lDTmsjEMudww5PWc31
PZWac6RfFxhRxnzpWeaEjPEbil4oaRTWRLcFNn8DJUQpBVKurQHoXqXp8WbFXWWF
T3qjKbxVf2QQY9nrwe183Ali06ay6qjU6uA1D9eYCPJPZv/PMru/hYdg+TJe3ySw
p2W99HQs8YsWRhbMqhlVDhygxP1jEgLn4A6m0bt3EKnyAP+lFMOIFyqWpDRX5ZC7
dWTo5tbtcTdu1FS4gsymtjPLoGApkqQmS3H4qXNvFZBHMs82pR2qhOcIit1qJ4xK
QxdQCPqY7k+XX/53yKxWx+4pK/9nn/jv/QXDVs31uPnM4nxLNqltE7+BoyMSkruM
Z/cw/+IcqbcK8T/GlQD+PU7FI/JSrU5FA4SVwjAQPvCPgsbqAVAa2n8yKz9G81no
uSvDK+BgOPwY0ryBA+794qZle54FJU6J4tZO7RYlsPL2hivFQX6/hAxQmPXs1nNr
f4JJj4mrxv9YBV9kWgFb91YbkM6Yx20PJaR2BWBdgNtCG5z/rbOZfy71On0lSSNr
PJN6A1yJzVesLOmOzXTfEgclKjprvWPmuUfBZgyM7poelgk02WYpcKidgCyQUu/k
Um02Fa1HfeN5HygMFvYAPW/+HaS3GojrQVxAVR0Kzu79XvQHktqAZDT32YZXSQHa
hFmOg9jEz4cC6PKIZc8FtQWUWNIeXSIZcCQ2Oy+LxVTct2HJe6flK4C3Le4OJRBB
tNY31VbLlugEnlRyf9Y64KKKaInsP7/Erwa6Ar25FNMOVtFrLtGX1Iqk1fMBBJnx
rM6axAIgb4rYE6f+hEU0xwyrbZaYY1Ti9uRuEKkdrlQiMh0s2srNEJ1kHeU6UvoJ
dtqX8nN3fDSbjlA87pad+nIObrBd/iZ4aEmVBMHfgBAG5UYwuEK8WxdoYPi3PPJw
JAw6gFre276vUcoBU0QI+8RY55m5n1cmh5lcPUuKQaeV8cpqhOBswhZ/km/STQWi
0AFgJgSExEIQnF8LhwNhCx0rjeIQPVRlKtcaRBeNcnvpqBC5wzr5afpQEjCXwdOx
fEdVJtyUNfdGrkyvSExXHRVA6tL8R0unhivYJab5bra/TWqeZuVSe9mQnn+0Q9ns
hKTSJL9E6wj7st+Av1JIRfMOOUQZlIXQUqGw0kHGQKs0YNbW3znY2ExptJnU34w7
bXj7Tn1Z1USvIaQrGQaH1AgEsIOA7oEYSVuRtR8S3SS6BxTVj2jMV0W128r0c1x5
NBg6SM+W1oA6LF1nbo8spW/tb1iMV7DzeZACdYoiLj9PNKiV73dJQu5mbvuKecRH
HpRlCGuhnUY1s2ODoAJe7l+Z6b9i6IxhTc3eQ61ReeG6wS20aoJWRH3WsfhP4UwI
Zy6Iw1ZWfy5YpBLoJ1wXuuSIukjN2OgrDy+r2j0to1xKgQV+pH1tOUKWQq0ul9cP
d+fQ9Cqka5XIe6tHjw29nmpuQzRspeCgxVUcZDr06irxGw+fbjoJpOxH8Us5Lj9C
qAifcn7rCiMPXXJqzeRv0IHLs+DgLv0crJOvfjjD88A5qw6w6OnMjiuj3H67BLQl
T85JItlx62tL8gDx0zhZlnl0+P8It7XE0/EwFy2RERNaimkp6lnhsmIHHF7HdhT3
WK3+PX6iGHnoqoZohly95wrWGO4hLXNyHB2/u+rUVvUEcLqLQlJBxcfLxmiQUauT
81JDjQv9K0P5kTI2kfQI77f7l7vE6K+5LxuqTXB7tMiRI3F16FGAPy1wUvkIsJZb
KuUEBSWBm0mKN74oGOvhket8E9Wv9qSSucG+8tmF2gk2GEDyVbpjWHkMcbcstH1M
`protect END_PROTECTED
