`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RL7NbEo/n8TEvLhX2Uttx92R0H5V4BtdEaDnKNKZDchixjVhiMWTY4r3V/YAiqij
AchA8GhHLxIRvtJKaoKSjHLNWPkefA+iE95drIRd0HnSYb7YOFgdbQXiguvD1ZTM
oe7f9wBACS+2gyWEmyFGqEoHKXcoNKJua2YQIXC4z1rADzmZTiVEYHt5K2ZZTuIG
3ReimnlctFADd6XjfhRE7ojC0BgQ9GRVT8PQFu1nF5oy/IxyASvEdC05Zq3Ebt+b
k5GO3WOqINBrQgOzC8RwWagr/8g5ao2sQtsfYUK/OJLizHZZd+n1SeC49zBByX4b
2b8RjoPmnTAz4gsjOb6Eb1CytoqViyX0Ensbv204B3p7TOb0bpXDb7FODZ5+n0Xp
1bwz7YQmQKpHHYrXL+T/+bXGsHfOjMqG1MlCKNFTRHmDlYu+bx70FWsUjZMbjewb
zgw2av/8n3sUYAH+EN8aaGPA6w76Ktq04m5NOBnIt+EGqj0paCcSq2jI0KyE1AjF
jvnuTP2CFZxGSYSSnr0wZmnd0oUGf8zI5OVcxUpy+61K+pK+S+yARlxNskiCoMn7
/B+dnYGI2s8AhifTZeIbfgGbl5+gbv1kgBXVtIeY6IiJNiiLnjfjJxseq8kvIqB0
HIRzJ9eoA56SwJyoV/Fifav2U+6FRF5PidItR/4FMc4=
`protect END_PROTECTED
