`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C+GmndbQxFtwC5MxmTFlKfsQccNv60JwbXOdY2ZHvkenPSQC78/gTC6OujVceZrg
ePsD0XH3+d12JbRbk8NVy2nP/ETJnjpLpIMkGqrq86b99amtIBgzvOqhDqPoGv7G
mtqrBzkIg6r+nLwrw0fpbjZ0NsKZqdKK18AnNTo5SE4AOw/aSuSBRRniPxk9nNFB
p5NvxDC4nS/LPRJCgakyTsy31o4wrgDaz6yqoIAP4UGYflJ2nLPXsJlrysoOXxwa
rXbnzNQSwEGFQ9SqUbnL8BZkRr5q1xvcguL8qc7shJgM1wzA7RnagLUliPBkc9gY
+0kvX5ceG7saW0oo7YK7vSQwb0rfwYpt2t+20z1L5oCFx0yvrOM3J29CRHpr5y4E
AEPkBBXWkk35MpDsJf2cnv+FWeMYC/L62Lrm5cocfVvi159iHSIKTAwWmJQCU13C
`protect END_PROTECTED
