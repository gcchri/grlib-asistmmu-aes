`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8PDjWhLlwApyx76Ah1S+ap3QXY85FkIYGP0vHqYp87SK4mu94QAFB1lMz9twXYZI
s1Moi9vEQXquwhchvskAEsHxw1MRftCpoCPs8O7huF5ERMammotGMRq0bWAhprmY
IXYtN9RHBv8LA8uOoqeceSjCaxRvMN4Q+Y6OgGGJuVGuTdM4h7PguOJNx53ky3Hr
idaNlNCEt6pc59WrrFREn7PDKUf540pP3X+LaRtv0+JdZSxz94rhOZiRAicrDSrg
boWJwFOFZqSaHIiaHNf3fBMawt0rbkgU7EvHG+XJFxnQOdB1hz2DBCuGxAYjL2ov
2/asDNkqZTlVOX4Es0QCpt/iZtFrrcVP68NrGZSSCo6SU/YuoPElEUWQNMTxLzqR
K9vpirg7lX39XZ64LSrV/g6EXEyKy9pKUEvtu6vHAaG2L5W+Id3y/rXZYrxN3sWF
aR9gaPL3Qnzb9K6pAnm6uLzJ171YxF7o+mMTbw+Wojn/kF+PtUiBq4IkrLKXzd+T
nYcsrEsWF8vEBpbybY1z+yCXlFe0r/3jTEZ9xQkIsp8rGwlVzP3zX8SL/P2TkQK6
TwvXxxFkhaj4p5LlrcugBe+IKKDKp3ChUNG3AqgBfhbrSA397cLkqLSDllYxuVtF
6l5bR69ao4aQcM9wwNnKfNfiNt/bkpZhPq898WbIpLXTdkv5SnMk9/aPIzNaD6Zo
itOkFTZkNn2H8twYklaZuRHAL7u+XlQIQs/t0w/XwBxrBM67XZpoGT1KJkbz3t+m
`protect END_PROTECTED
