`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0ZXx8wPVP3tc7X7jS/WzC9s5bJbnPCNYw+WgnzEDVAn1d/E8z2E50MYH1+BKGHc
c6Id5Q4+bLr7m8waazhrdpxrSMiFV9vfg81OTIAjHlkGXRCSQHC2naWo0FS4COsM
VlD2MJGniBOXSkzrQfJSeyAZRB18/ynb8M0XqHIsrC1yf0LrCCSNZ26vHhYuTj9X
OjkfFBuIvTidqvtIiMTA7RJiNyv9rp1/4+Zti7XWXPC6LrqHfExTMaAZSugLvapn
07XCd9db23WPshx5lpKElhF0pnwmHVF30BXA3+Wb150XvfAKMwiYOSo8foo0CBC1
HIOYQYqmJ1Q7+Je0vTBqUJORzqydOFfFEGmRGxGTYBGGuYsmKNmjEWTrz+YPYUyc
K8+fpzXJfFrii2eX9qPPzd/XVbGGhPHfQQdlceDyZC9zn/mJSntvLGXdecyHV3Pe
XMySOzWZoCbJGSfxcLl/JUpZU8IulkpcyWESxVfXQ3yO1mka0f7qn7Vm47/AgJQf
7IkTLudcTjJw5qaD8yQrZVD++4jPOD4YKFLQ1Hx1O9EMlZ6IHc1CWTRea5KQJ1Fo
Xm1dlJ0yMKbqncJaWO9wYud/Q+ZBVXWg1VLyyApI3QXEGmwBy325sV4r9pWSJtrs
d3Zf3bifSsIbU4BnuA2GGkrSiDTFf+Kimyg0q83h2KRmZ2YcB6A/aMpnkV24G3OP
KEXc4uPUsHbIZeVmgEfQDPWH6N58DKHk2/LfpOx0wocOnWcYcpqkt5R8hN5XuJo2
aTFSK/ZYrz/mH8E5bopao3G/0gFQdk+fcf3MG0E89+s3b7S4rmex6vBoI96iboR2
tYCj/JSC8oNvUZsIOEk/h9AYdEHwbkeJ57kh0Dxt5QVLtEf7PHu3YcMxeITLoVry
/qSMf6WZzgCSYJSeSHqcXOgDagZO/GNqxS5kUapsVx3P7nYm2EIlePdfkad2KVDe
GqPgyqdar9p+ujUAn2wFqT3o6daW3zvfgfXkphfzsH5hQceHHhglbiT17FOOUhnE
0y+8nLvp+WP46BQcU9ZflvQD0ZacQhM7biZ7+Jpsev5RJ5lWkjyuEHO/iMuY9vAp
6cD1YSTHL9q5OhC2j7SkcXAuz/W/COLtNhsTaus2JncdBTlLz+s0FwKe9awfu0e2
PXQD/ZBwXCnxLL4v8h9+OR8GGyOCegBSRD0mP8KxACUy5C5sjfKavL6r+J8Ue6jW
7VkLooJZBpCVRdv1BT4yRkfW3Pfv4LB3G69YXIpH6M8OSROuZy8zIOE9W1A/OF4U
evihnk6izAykyq6IbtVX7+2Mj2ont6WxxrFwnzPIn7gg1+qv5WuvccZRZcNcJvRv
rIZxVWgHLD0oNj5cx1R0XDfw5E6QLyLYFE8bHRO4tNHGFPOCmwduQgfPRMDfsAn7
+Xz31S7wdsMQRgYZp4U13Q4s9FBUNRviiUHELEgOzNtAmxAOdI3MzSzxgDm59Tas
0swlXBUqWpdHg1BS6JzGB/3qRCZT9YgGvbvmqTuAovM=
`protect END_PROTECTED
