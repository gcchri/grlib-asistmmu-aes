`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2PGyKtB/7tE5uMhkwLUHu1z3SIgOrrePPfhKCUUktFkCZYK+pJyGE/buAD1EUGnF
q/3XSyOc858jKg4U191nUplA18LaqoQRPpV5A09dBab1p0jZS/Z/67IuyXI2k3cR
ZnpbSbVsGSTT48ZewvQsDtSwRxLHiy+ZWimRc3Y2bPMPHoRNiSbZYTjDTgol8zLl
9zZ4jOig8IWcwfScsZYEsumkxldszzkq6MzhzzKmZ2N3iUc7l5zveWqELOKRtx2O
dJn5B76GKjrRPYN9ousP2iSkbY1wsiNJnDmHu0HajG8ItsBaKy5BPzmr9rDWWQ9/
NYx6WxqZH5ta0dijlm2TH3xqFlJdgNU0ZQujCXS420XKYFaBrOUKn8e3H5H0W2WI
GSnSKVFgxm4NkoVDW3YyUQ==
`protect END_PROTECTED
