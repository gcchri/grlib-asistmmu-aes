`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiaF4xtPfLK2FYKI4HFdmcsimP1MdvYtApUQEJvgFAbnlNjufByAIfhhRszToMKw
FL6TGjoDNXo1RaU5m0brn7UB6KYzOcUecKPztNW8XJyNKyzLipA4jkKQ8uNCi5mO
ECPDiDCm80L9fxUNsQMqV/f9Y7RS44y6ifAzuy/x0T7W5/VNL1N7BFkyG+SrwsRL
YPriStnr7RgYjp7c2eB9Pk/Ze8oSuuF+x4/sD/ken4Mqk5hy6a8L6SMsWK/zMja6
T+h1X1VJ3OiB8RyLOmk23XBpJQkv8urIR3ki9vXMvxhyEwTWIcVDVum2YkYx5h/N
w+tqGp5BNnVuwyX2mWoWgu2DxqLiURsdlarDTkypw32rvbB1n2STRD6RHAK6n3/m
NH83cY7dqhC0uwQqU+yjfENHP4okzthgX5GN6sDv5XL9GbUBE/w+9qhQ3agRhozo
RfTSnKpMi61gnEHsP4DHqwoOq0akAC+qEisAJGsfZA1TUgAEixlRqsnm5KzkISFy
b160sjQ6oTVoBW5y+jmx/7rbQpAsrvdapKjXtCKqglnQta9i5B7OCs9Me3Blb2J7
`protect END_PROTECTED
