`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OiGxKci1Qzu31Ga9DAglRNtNhsuOO5zbayXeIRrbBaFMK4SR1ESfPiAOtWM2bv4E
sqOt28U5s4PVvH91cZojmiccT06d9Y6lFvKBwseCOk93ctvV3CGBYa0xcR75UL3G
l5ZVULhwVApA0/lxANMx0p2TXbKx47peApAbwq6DSWy0XpEiY4v3DYLdmbvu5eRH
2SdTB+GZzrsm88fVF6yvyZ7EfLq+pJmkUwOF8A0R2SEsH7/+WQUOXI27jDLFVnMP
Dj/Hv5aVqo5PcrfCFYxqyc3/BbRVxe7KWM97hw5uU7CV2/2MV5B/tNFI+jEcIGrp
Uba9g6Riy62NrAeCIejzDvVBQQKE7qzwOy/Cy6DXSa9tT0St943Cgr9SRd66vPGF
EvheFgOOWcUwQrSr3KTD55NHqvbnRFbv6dX0jWgAOiTY+Ic3KReEI+uATLYSNu2K
G8zhpYKAW0ltqYRm2gLDkJpAvOVqpvV4EjbUq1d/rWuYqQbXzkPI0X0+dXkXT4LD
eKeQ7qr7XK3Ur7KVvirZG7eYymiM70dituN9UuigKJ+GV365uVRVeK+RIk6ANH1D
`protect END_PROTECTED
