`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSs72D79UocHqEeXQo7e3GrYw/cTsREABEg8MKmg3/N2DXpq1Srd7vPw8jXR1J6V
TL+TeqWEBQnRtCgFzNGSH6oPFzU7S9vMC0cpavfDPiLMT9beRSFNBMkGv4huWB/n
qQ4jU+fApaUDQTdSYpfJ0FGARzeP/xv/rbdc8CEFINdlMd99hiNufU/DmoK+Fnjq
frqEpOe8P5I52x3IaKGCD9FwLqnfl7iGGoa12J3FFbkZdg8pnJlbDBIcWXyjNbz4
wR4wo5QgQ5v0cwDOwju+c3YI0a1BkZ5MA4Wo76oCMCSzEsOAgrX/Gu6q82pVoS2U
RVnUvB3Q86j84bRoZRaNOuR3OpucI3aULeR4aSocwHP3hVLNZAI+Lh8HmyVyu1kj
JSr1a7TmoN/BrtP8U1SsutEYVjD9JoQShykwJWGT/BKxOlgv16Y337rTLZterqB7
Bbs4H8Ts0rXXASNwtXi+qg6UWuHfTpjMwZNeJDmxF3KoSLDgbFD8Ibu3oFGXj6ZN
b32eN0MlEeLiiyFINjzf9UN1BUT9sRtxcppVFtSE0ToBUhVqyyf+LnYO7ogcxV37
qo82nkLnkVhP4+kIjEg0elSReA8BY5+g7SSMcW34x5sSs2jseKP07/qfEY2U6bt1
Mj2t9rT9jnrMu63fUIMFywfDY7CXe6zMEC1UxhzQaN35u0/oihcCETfEd+O/wqoy
KUFdKnAWx2Zkp0NfBtz3Q5k7aShAc8chL3BAaJg9e7jUBGy3GVaHlYqWiWu82bmL
lBeCLYukhMytv6hLGdcuDGFvnSbdPwgmB/Bc89trKPWK6mk6NicTYQQFs2VDob0h
l6R2kfUt4oUwj5lz5GftdJ1dNC/3Fsa68B1DI4fqcdoawt3lCt6VCSne2PG5CiC+
lSQMwxKSf0j0HVTTW6jvNbOOU/pWRZIzROu5pQeUFRxoERzkkM9uB57UjKlYu3qn
xbMOq7Eeonk3OuWvZZh26lrG74SY3jpBIkt63kj4ntL8aZLZPNAKqoNbgZiFw+ES
CX7xNlhqmeZgU0qEtJyCy+gXkWz2GI/9JIc1XfprzrH2HOaaLYF6W37RHmeWmfU9
VCooJSGmHb308+Z+TToPpbSF4AbGxKusOLirXUdLtUu3m1/ER3TLpjeRQHLHiFGV
zrmGG7fO1RPAmQ57EvhMoAALAJpbucxAy8FtqC1MmWTGxlH8uX735/LZqTw/GwlS
x0Qv6W7nCvlPk89HWYX7OoCzn0C2DbDul7DLYRii0/MwlKCeoTi/6AjSAa+ijjWs
9NixlJagITINvPNp+jFwrPfaXDv7TnqgrGJEQLu+9dOQw2wdqMaL+NAKlWashqr1
Rh6tZxLLhyBlr9zCv4edqidM2RQ2UJoykuUv76OI5D1+DocqaRo8nSj/BIEy2FlY
vVJF3X3RdBekoqToTEbqT68z3ycEQcMMPaVY+hsXUCYbskeyZsxpIVrRMbUxUwgK
XJbf84r27tFNX+J1hREr9+3iA599WuIP8wGguqaB28opG9oIGY5XI/MlEie1Xijt
4030CBuuWBDDBg8/3FRFjQECxqMKl1fuGGeyiZrH3IlNOeVH/3chCzkjEUePGNyR
1ME4r3JllBqX90AruTgbP11yiRFUdo9QtefU8gvbcNJx1HJYQZVSUn+pfORv83rd
P2zGkJT7aXrmqhatuEcTrOsfUk0fx0W7zHFS2qNxIW6P80aw4kR5x78HhBp5w/Ym
Q7Myw14jq/JI2nM2YreWtTQHSCKf6MJA0WY39gITUOtWsqY0+0TXZArCB5rQMGPX
SJaDKEwKxPQBU66+hvtiypFPONmWDw69W3O9ChxTpZzuh6mOcuRpniFHB0xQISuX
T161EFjSu6T2/M37e9eMGmpCZ3QprD0LLEipzxNh24Q/zrHrfuY+m4NIe1o/TJZ+
EKRlTTmILwvyMTkBNIgmQyhAmtfvLcGUjS7SUHKhWxeWv6z77YFh0dXRdH2KtJ6K
0TiDd83dL88O3gyLHNWnhemH2tYtsnItKIfHDLlKbntdCavfk0f7BNpbuyfZxIY0
/fTchzyxI6tQRsxy5yek7Ostwr3XE/s1YDrqawUDrvM7G+kb6ikEOzrjlpCphXQs
IoRIlwsjeGQ7UaSC6+fUKOlNCcvS/LMUYJhhX/5bfoyEI9Fj5tmvgTNzbiVDxonp
s3OBRdpfPMDhlRf8EdGxKTRQ0INvc0utaLnIJTAZdFUcUcAftMzGt1QFXjDspu24
nONI1SaTaJShLDZGbdox7Fv87YkdQOW7xJ/7mQoEQ0NN4d/5ydo1K4IbruTWVX6R
XsGnBb93AssWlLe3B8rjg4bbPJ5jyJC4G276RjjsRt80gCgLMlsdJEfps7joUm5e
IBcNNvC52tvssk4f1AIOgWa+vac9LZxEXuf/YnRwQgizk74fenMhYf28NofNMHVJ
NcZQ1V+qATbRuyZESLFtfMlrxGaYgiCYo/fNr+uTi1Xm+aqY+WciD9WUX8H2wxim
jkzeksOHrCarczK9bV2t76sPB6NMpDEPDNldkcJPf+B8VDOmfZvjh0Wf8RwKSPXH
jNvytDmP0PlKK9+Za40Ah1+caQjgHtRa/wvG84OkSnB+mReA/jvLYx/UXNVPVlcs
J1ybMDuShpoxCxfKlKyAY/6NXJusAPdGrYMfG2R0jEfak8jMtkw9B+tSp4PShYzS
GgiX5rHwOTKVSEbhbwSh5pTmcS+hAPUGazCelGmDWd2cEkmT/AKJYjwDqqfbvBZa
aAba7DzqdJiqeQk+oqzX2fSTZ0auuW/rR4o0vOeISCssKg3yr3Pttap9qL/YIphy
29E8Hl//w0pvpiSR8jHWSXCHkZtJMJKUS2mXkrPOSvtzqXSV3bWpOeUkRB6yZolQ
w+9mkDFag+goRaK7EhlvqUTtKri6V8bj9yvqOZsvwz7UT+lIgqpMwbf71QIIXzZ8
nnslk3iT/N89mEWrISId8s0RN28eEI8kp/ApJcsEJFRWYDy+sdQdakUjnjnT4bvE
/xHvvL+4ILdpX3sgdqNQYHkns4eCF/wTLhuRihdaXVVYHvNedWMFgndT6kdS9ADs
ZmK9SN1bui8U5XrpPUno7nh8Nl2ZMBzRhO4tNUAmNYtkooU1jojptm7dXGeGJZHC
wouI53tUY2/PWdwOpb7VJHYzotfrQEHGmqJVBWlb8WEAniWQBV0iWIrjvwwQj/j3
WrpriFTlF/rfnpko68/uBUHs3kc96QZKYUZncIV6b1jZ3amoxBM4uFHxG7BTJqiY
2jzkx/57ktVEGN4iBEZjcbMd0/ivN3Qr2IjHTyuGxKrP8sVGXLQIhbNKen1Kamdc
NJhfEaHMIBqzY/XwfF19Yh3eRePDup0LXSIXjiBgyM5MwR974+mzzwwWdPYb2L3z
LhfyqOA3smsJl8Jrcev/8VjwVromclt8VFsFbT7nkoQUi1YfnIz7tqvyoOIPFBCe
iBjESlieP50p+dLDc/wK02qzZ8e2Vkdvt9b2qtzZQ8HebV9Vfhohp84j9P5F4uOp
oLUXgz8Yq9xJiDtE5g4xDfVth6r3CmHYjP0ccqO4D0VdOPi0zQJ+mnsRId0flXIY
jOPw2PNAILg/7T+yTV8IXzm0oWK/zSkCEj5mv2hCrDcjax0I5Hwrnkgo2kcdE23T
jCROvH1Y3YkSMuTcZjsdkZ61V5b2d9rZ/GBx3risxIORW28oicfSIwbsvR6TK24H
v6oYAeAkAnaNpn6Pz0muV1O4JWQLqxO+PB71NtjzpTLRAvvshLq631qX4mcYoOfN
TIqUm1avA/rXmO/v734NMlwTQDroykyoevmfZanq/n0eJf7Vl7S9piR3SIQRp3tu
UQbiZTcmBhMNeQt3/TuzUuYIogg07K0VATPbHTI+BQh70bw7fKGs/lSbHcxuQpA5
YHk+hSb+au7zcyi8x3gFCw==
`protect END_PROTECTED
