`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sUjXaPPN2BQj8EeI7mrUpLAEp5WFVtNiZGXYhnIfNkC8CMTsIO6AwbDpRBuj4hmh
nsrjdHnmMLqTaV9J1A0YWMTnweAZ/nuCANUBgXXuudOlr/JUI2eRH29gyyX2DudJ
GufSMdbcgs3xOR/cEG+CqV1AvrOKlldyEhILVI3vsE9rgu8pv5r966O7IGZmdC7M
AhAX+4rHKFSFItC0Dk0kh+6hKvtqHCS0WLRiGQOoP01XWq9663qd7wqtqTQi89t1
dtFAMtK/F4jRavAE6kNRPNrzRBDFOx0aSQi1oWfDJJXVvYBkE8XHk0CwcJzaA9xN
h+vMzTbXaOU9tbf1Mesi2FKWO7ZJ+7Gv5Pmp9Ykj4VBJdS+fGIsSABohlclqYCKP
AF1laxjLdJe98p6XB1hMN3OFQ/gq6ScjPpzBP97X9MQweAOQgde8WvPJ5pm4xlX4
hr/fdXmdBc7ZP8HMcKzij6MTiIhYOa639tT8GBrzRUcPmk3Zocr5ORaplxWUEEHq
rnU9IzUkW8T+CB+cBP0eys5VSOjGmuixVgs9GiK000y8HSzKH+K6XhPv4Dy69e02
zsJ14lsPafg8wm0G2AjISTtGXeDidSF9bgZRMteD9iHCinI2rcox2iUxa1niX7Fg
FMJjKQ2TFdkdyAgggGiseA3jR1wB04j+XPXKHnPuJnL1fC6oLgHmctfwtgPToK3R
zgqx/uiyEUKhRwLyHe+tR0GrurtNay4XFTcWUESRGvAEMDkTYETp+oKiLEvPJEf8
IjfHsD9RTAIv27W+D2NPvGt2fGRaTBWHZ37l5fHK778tkdv+8HYVI+pC3M+o56Tq
rtAGtJf/H/s0vnCjocwosw==
`protect END_PROTECTED
