`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oaCI1xY1FdSo4B8Rmrax3keww88qe0w2wsnT7bHotdSLY0u6rSsWQUZog3xJV3vo
/L5PpO06kv27r2X8It+FxsPuM7dfbUdl37+QGbyqlPFUHJ51pscCH5NRPx5zb9Ri
T00YXaEV7erTuh9NuPEc2sKPTdPZPEi2IMYK4zHbkfzIqPm4i9l3zpgVEZKlDxre
Oo5E3/xZq9j3xMYFNIXWyhBwacdJ60k6nVx3qBmyZFNSy0zxy5VpU/McuWbbp+1i
xqgyegAgOUk8f1ukyf+/hQJsrAu1aKzjHdcNNu+tXDvxkfBuoalg8uEmpcImLo69
KGSEAPv1ckbPJBdFr15BZRgd2QWBfXMJ5wBUOrH1vZAaF11fibda34Uj+R9rA00p
LPrLoRDJ2/KegVNNDInA29MITCtU2h+kJnCajx+CZjdFaMmT3WgEY9VlkwUZCHP6
tZzMO+1JnhtSV0WIIFW02NgN6xNMH4+EyPAT0aQsjI6jKlWRwz7JyoFQCsd71DqQ
We0HvoKgse3LU7cFabWWtdLW6buFgkB9SANXOeTFCnpX2hBsKtqcCFZqpR48b/vD
nzjTDJjkdqHi/+mBemHl9MNI1c2/d0krw0HEbWwjp7QUsx2fQXFpnIoZERIrQJID
dss9UQ3cPZmFPv6/tLNUSL5lwTrJJy0/bN/rhgP92cPQucUIHRMIbqc8fgl1MikB
zRcMPCOwXoLdAtu+lZkaSMoSHurSYjdE9gQS6ef8LGdHScRI09GUdJVQGszllI1r
94WWgCX71StcyW7RqR8LOrD0Enylr0RsMEvrQSpJxl+zoH+k1fkUhnSQxADwK4vn
eLt2U9ii+ZtvBitbGCCpoaPvGBAcMWnmsS8xfxWT3O3OCeWGQBm1DvqLUtJDwuJ5
VFmHtVLdgM8hgyJAqxjSJI7Wq8sZaW5mdk+0l/8jiu5WvyzNlO7dWGRDnIm1S7M1
frQTtVElflEaqw6HQcMNMuOkrvWWv7Ywg/wJP90rNEcj9t89DlXrK4reFg9NlG37
Rn9WrBx4vmIos77s8S1+c+y8A24WzhxE8Cmr0RNkKoggF2tXMRYrq2E/TYAC8Nvr
1F9BcydmmVsRejxWXKRi/y/8c8u45UfaWQR/vdRgLdXUGMBZvnogrdIFysdaJS4Y
a5ZjqhEqf4VK1ddURqRTBNRmGOpZoZ6ietmaliHMoi+TKorTdnKpxqs4Jl55TAPT
CATadsog402PzDwe8lnF7iMh7PQUhcmDgIf0HOSwKa3pXE7IYyB10YF+oXhOyZT0
5eDAAvLvOD4Aicdd8j5A5rndxHeSX5FSywZXP9GP8Aw9+GXd2sCJKZYb4AT+LO05
l1Gi4vy8J2TiTlO6/Z6jZZVoOrUBdwQwsFopX0fNYtnhXhIX2jpyIGdqxxNl0Clq
L1XVhoFICyfYz6anghm85oFeZaWpgl4aNGELbJMkfCvWiOEvyyWTfIsXHLkhd2pA
B4ROwxJ6v+WsvEUEhQXPfx1tu+tL57DN7Sumkcdrz1f/kMrMdAMaGsV8CMmzll0l
hb3jTO0Zba5/q3lbpJA/ShF/EQPHRMv4U9uWpXUG4/Pc2gR/ZdaiAzn9Zc99g8Wc
4teRPASD966hGQ95KH0gyUAdwYDTKvOKNYl1phMWkxGssZwZ5T8Bx3Y3n8RK+Kiy
qxd8+K5VLq4ID0ci27psJcAjEPY/CAgzp5VzCRWg4YE1Y5j4cWdfctnE1+zDhwpx
22twDcggklchGtRNQtZkThySaRoOE5qbk2UqZro0uLxVDcScFcYTKqWXKzLAUThD
gDCZ1lJGPv4EV3X4lThFOZuxTlQwnU6HSgawvh/dBZzPDsUCeVWYH5KZ5F5agSiI
ff1qkAMVKL8+ChrhSRHDEL9LjjTwd5JnsbAnxIMWzL8=
`protect END_PROTECTED
