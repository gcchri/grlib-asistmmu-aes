`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N83g55ajzPa4TdjY6LK5h9RcJD2I0uIAdjYyvfjOht+s7uIJqqKpIw+c7O42/05f
h+bR1jmMieX2MRP8UONgYgsXEeabvEz66eo9eNbSDeX8DY1/BOq3/0jMTcOrcjVD
87otOQrA3p9nwqrGeZMf7XGXL/9e28QxovpjKuf+RJ/yKotUNCdO6g6C1mP/WUuI
wnu24522nFHW4p0vMFMl4EQ6g7fY/0Tn/aQjMJaHVVChEUyo7I62Dyxem0Xag8Al
1oUqQhEQWjF/8CQuJm0b8Zo0sU8NVdSQqw12+eqcl/Dq0zn8QNgLLEsYKGnW98/0
2Qt3uJ5AR8/oC/SOUpBUA0/g0UDINd7ZmaP3irBSX1e3z8pYgP0ihqQEyn1W7wNc
/JcTvjb81rp4otR3LWl4UMTYGwCvBJt5yQZOEeCOLMA5Cc7TkS4wetBC0sFf7tvV
kJukxy3C8qJ0g7uud+xYtrifITDVbyaC3OoPl+IfYxxSVXOKnjdZF/MKmJx967ZB
FqwLCBHatPTTGb3KzsddLtg3LHIvPzVX5IijVWNc1RJHH+c4DSQOLNRvsmt7NFx9
TxZyKYYZ3Q1wpQi9cv2rOU+yqmGjikbUIGAvydktqG7Z96U1zbOIBXAVJURXOkKC
cEa9wuDWy0phKxjF3P3BK5zWk1OOVv+b7BC2KRjQXec4cBzWy+qSepa+9V9iOOmR
w7+4WKEdHr6obyJlDdpcihrMh0aB61U+/SlGcVjJEYvAsah/XmN4brzJ26uGIaV1
UFDYDivARwozW1uEoGw2c9sV2d8gslPSX2ut9I3lOKZLMrs5rp80UZkj2ndnSNSy
/bCK/T+hYpZQ6bvZqj5ieJ+/Zh0+zhXsxaUim8G+5W/zOm3ULj2eEmeR9EcJc28e
O4QjWLZowfRPnO8esdOE9c9uCmM9PXfUDkKG/9LxCRw=
`protect END_PROTECTED
