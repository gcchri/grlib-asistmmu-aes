`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MpK14obM6lcjYWiDjPi5t3R2XBU4Jvpee24Gx+At4LCqvnO4B1u4NNicWhs0L0Dv
KmTT+9YPCx3d1mRj+x7Ckj2lnFo4/ZyW6yqEnIbc3jVBaNH6M5yblYqNJnUu43k5
6R7DzB69fLiGqXrfUH3T5eQ5p79lA+3/Dh6BDGc8HD3aM9RH7i++XOn+91TKmhAT
HbRv0wt51r0XaYfN3EceqomxkfGHTsYafCggE8naL035/5FJSypRCs0SEE3TTIFF
rwusLQvcYanNyPESO+8Hvh4gym0NzxAnos2Fod63pBwcpbef+R/JLBIEBK1HirUx
sOhZR4SrsGh9Pe1OxEG4Ex6YrFSQ/feSbmIqIqNrFlDjYCWv0F2ONRy6V5CP2jeL
HS8G0/EhAVjzCAwaOBCrVLDDAqD+iJ+CrvvtMKpIbhJG951Lmh3wwYjBaYDW3Uxw
+DcxumJAMmr/J016efyId1tm6/GYjJcTznYP+MoS6CwF6w+TdRGYT/6lNVHqWba+
1V+ZnFAsXlycE7FjhCjTXXh5BcvulCi9yxO+wKK+4AqT7qqMwtWB9L7WANT6A/rf
HnN17kgUQIKkDmSx8YJSQYYgSTKHGrD9weWYBz+HKshcR6EZ2z6peezf4n/ZX6/4
p2gW3YPd9IFpZBprxSVPnJfN4ICyiG5Cq5Ep4mcYz/1H6kSbRyoj92vA/PBfROwP
dwCHqtqoBU0cGpd+wfcD6jX+raryEB+xHxLcLu3W5QyVne1D/Mjx+EY9g1+G8kVa
/2vIkLwX7gyw67QZ+Ow/KppDLRciP+I1gSznohvVtgy7kZwU3J7MvstmEJtpYnpP
tu2OdZuYZDbokFjpJjbpg1Hzs6ryn9RVEQqBvvG72kHJZ44t3VQc1DVb0T0ZPCqK
`protect END_PROTECTED
