`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ikl1oKKFesEpCRF/grUJpvU1WRdE8tKZ4Nf9yv0iyvW6V9PA4myiu+KjonuzrshE
dJ55dp3fd+YMxiIwflwvDssidrJp6TQzU1NKrdjcC/rMkoU3XYzkZ5dHmohVFGYj
txfGER8y9pqEKr98aKJQJxUDudmE0NO0MCJYk/3ZuBKL3Ialaw+SznfHnaZO+U/b
aTPdt8LS5sfp62n/IWQm4+oz56D8dabEg/IG036w/01AnvNfDNKGgaqBm3IZg14P
8sJRmhJQm9gvobhPGX9JlZ6JURxahOH7prZtse7yaxl6z8zhpMkchpDOn/6ucmyh
dP7O4pSb2D48N+HzJaO7p9InaPEHq3kVjLKFmooc86Pb6UoQ4htlPOPzDj53jGkh
K+XfQdXuh/Z4vpPYNJWiH9v98WrhDR8s/9oDjpuxgsE=
`protect END_PROTECTED
