`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bU1L5/E1JXYm7CEyFBm22QWLxKRrK36RJ+dxGU654ASZLCGF14HWWoBUPsy5EQIi
bUbmPhJJhCVl1xzmaD6KZje8uH0tTJPpUtN+xiXThf+J463+G3tVI4qILGRlxvcL
u9kzngFcr+jlnHqMo+nkQcxdZ4+NKbv2st4dlIjvlFR80aWnRs6EaBCZS6OBfivN
EhnyNdYjFvq3qQNdWXhKpmonhwZkYi+qV9t4pHxPsoN/n48JHj+v2CKNIfYwhNXU
`protect END_PROTECTED
