`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7FyMLIHeTPyrj4hOmCL3mmlO1YvyIaEf6hO7Mub4kzZb0xzL5QZ27/pxe+rWO89
twHQWIVfPXzuCy1KGzmTvdeZncvXJMReMHFvcNktdzPgDSBlumT0tO/68WNg1Izo
bzryBxwBLNjEjxwnKJK/d0SZiqnmD1j0g/QwO44Z8Vf1euWhV56RBsXVK6Tk2I3+
MDGefrbwHys0YBOL5LntNXZq+3TUKDSzRZ8vW6W7JCvCORmqVPQM6ljxBqUpPukk
EfOs88cxqpdELhwA5MyZfcEmpUHleJvkqf5zz6cJuIH+QHms/IRTFSHKHNZ+QXMa
Kbg2/Is8GBSGx/zTmneuptRvJfkajZgoleix8concuxo62ryzko0ETVDmWH2Lwjp
Rp67msRNmL5B1yOJPSWl9ysRX9HrYnoVKpuQJBXhfeov/WwymRgnqkxCCu3YjYSk
Sao1RZvFjVm+aXGUYc+uUox9/QZ2tloz1BuD9Ee5Xdj9PsQ9AdS+vf8STN+qczhZ
+zgkNgkZCi1+nXnmjgrHPYlDWsbC+qztiKb6na6SH6yWJtVhbjMfbPo2yRkG1Z3+
h1HgRotGYtut82r07ywC7JR7tivBFKJtFz642ISdMNY=
`protect END_PROTECTED
