`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hyl8L9mt3rA7RcncWKOFQwedpsf0NXulazsYYxW/C276VhwNfBbW/1vwdXDjlikq
sJ5XtmKrZQ3HqE/nSZG/fB49W4jtlNUYZOlnGD97ZY5aGmf773eZKXkvb8I1EnnP
O6z6h/WhVc0NccEcRaH0C1m8HOvzFp8v5Dxoy0XSQCcw9eW6ZQdTlD7sQ5A2cq7w
BBeS4R+He/OTsV95yFg82yzSdgjqwteAWBuvlMJfMH8mSOJd+5GA5TzvDYEn7q4a
DQXSwL6CRJDg8MD+Drx3CrLMv9aZtjlxrr17uFN5RJq5LJV9lHubLrj27XAhD6Mo
e6TE4GZBR2u4eywavFT2Zlh3fXk4wKZGuNlkjIF6JV+fWL6XdbwX6e8dC/rm5UrY
O9XBLBQo0K43tTSfeook6ul3Uh9H8+eIPnJ1/LW9jc3vqyDwNiZppvM2eSMGED69
TnDYQkYF2lIzliCbWyFfqwYfvcuMmTPrTsPWnzTg8BU5WRnIkWnwDoTVzobu4Yoh
wZ9XrKplaPUZCwjtaiceB7lOrtaaYPZT90ZEa2PDN/xdxftAaqnBhYJUK2QZFqYg
2oqdmtnYCiuQ93Pg8f2WLdYv5r1bvCQcKMOS5Q2m47+/cAzV14Lop1LR02IWOFf9
jPXiUZa+N7nDaLY2e8z4rlP9Uux5bn8UgUfDH1fVBp8VXBtZh1K9J34qzoGCWXLw
yiT33J+uObREPWfXkJg/XA782s22GZ8PniUQID02GimyRaQUqHhtFJY+YcrlTFf7
lLnhG4KfkNXM+fyMRyrUXzO+OfP6Rlk1S/d7eg10kqoaMKs4w5OcPzNw3YyP6Fz1
AOtfIAsymsHxsjUwxQvJ+RARfoY39MNT7FoQeAMZ5OkVqYvPliVsFXVNUt0A80IX
sBdsqQxQEIf8/tgMI2XJBGvQ/7528q9N+/iwcz30x0A=
`protect END_PROTECTED
