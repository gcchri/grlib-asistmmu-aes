`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxoIzXFOrPwGQF9peXQg3MZq4+LK41AACPWWX1VPleTJ8OcnEhX8jEgm9OPLHJOZ
DmhaJ8bQTS3jObhY4o+qSQd8Bz+GJzugxPIsV/aC2mAZXSoNpfO3yyktLiX662Cj
grl/V5mgOvo1T9bPGa4IIEWDHXSjYRwpdRFg1IJUPHCI6VGFkZA+0CM4kffxyMq5
/D+c/wej/0XWUb61q58oJk1aYii4/lqR3nk22AaXZhe6lbrsd5GwHJAa70dEE65F
lPFf22s53JJCVdqu6zbNwKs1A33GqgW3dNGS9HhGqixI/+bOFOUpmiuxqC5L8c5m
zQzyCh7lnICeWlqQ9e9sE7aNnQLGWLm9FtLRDYnxhXL8VRS4V2aYH9O60AnnfzoQ
8YbS6sZGMeYFtfN5QXaW0d+LJn23hdU084TFHPSm2ljiP1VZ226c15/w95UmrF5p
RXcPy8HhYLnomtH+Ec5skw==
`protect END_PROTECTED
