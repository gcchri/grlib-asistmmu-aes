`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M1jjyfCy8fQYXUkWJVcbNxB7xHSEWRxPof3QHcWK6TJLP1TwQPHXXkZjSW/QniEA
TxOsJsdFN3Sc7PDikcgP2PVpeumx/8RGGYCLWNbLnu1qpnZRTPH2N1jcT1lw8Rfk
rEpPBsICO458utfl5uFsddYFLuFCta2BJUj3RzDHOge5lyCspwDJeJziGhOb17ai
TPcaQqRFgt4TzyFdIRYEOpp1ypfCVMopkt8TUylGLHWw5uhDuB+Rbqr2xILXdbaR
Se3JZnccotLsYBDf9SzTOtW0rJ9uL1e7zqI5ZkBZwAojkGGUZkWVkC6x+gkSGTFj
PzXwtKEe0EqSPR5ZTKxIOOxyDPpUJMZgPrAq96t+1DelTCwfUduenx3dDXK0WLTR
2m9CjVnuRMzLJA/c3NmqzVAybcIloOk6OAZqac7jHzl6duaKuGHMtiFe0m3Y5r6L
skXQxDVbl3au37DbM/G2O6Kdz+OudWe3zmkjAdZOan0=
`protect END_PROTECTED
