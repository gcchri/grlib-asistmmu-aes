`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Guy+W3oUAHJsK5eypPaEAlRf+FxEYeXBBlig2qjEDHXJwjc72UkZAaRZIymXg+cy
ppTPKli7pzhJnxhfOjIdm4vrd+M9iKZTItvV3+u+w+g/VVuf4eJCGHH7mnAZ7g5x
ytZmlv5BcmSnt2EmcSYSqPkwyugKLpffDUdLdFpWPPYniznUwHy7i3kcgkL+6iNF
sIoqdG7ne/vLZf6wePwU6SmI4ExBNcJgriIyTDNFR3APTbobFzGjZ3mjwPg4fRIB
SkoL5n8vPEPP4p6xuxhEylg/d9C5fldxcZK/QR9+wpZeTp4NGtPxh1U71ZZJIi0p
`protect END_PROTECTED
