`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nINKxPqzq0RF39osKAw41cpu8+SIH1LgM1P46IYjywGGQmPVNf/DqHJ5GqjXMlJ4
mVLNS3rSgWWoBkT6rYnlojfLBIAPJ9OAX8DvyaDJSKIC72u2drP2NY1gBfzziCQT
1cZ4JZwT4kKVqKn0JUSGBxP7cIYvM5EyHfT9faM4Lue4627gCn3a4GpPylYeeQAw
KbUGz5aMbYxnSlhW7dlpoBa5KeDRisjoIk1jMjIPLvs9o2mJ8I0azRBRmSkVbLnr
yGZFHIFCu8rLAisdCPEYb7mEOibsxSqm7jEt68aVF1eqgTBmMwd0ldaMUYf/VFah
g+IlNMIy3myYNXVMN2xUwSzWs/un8AEdabwnpJed++hbWtk/UuT0xXXGCDUj4ccr
BLsviA5MmqOAJIyDiOOAAGGUCpHHt15YsrPtQxJrp6+v7xMTy4RgzUxvGop5fy+D
HwVKOm3vQUYAJI+ivd9bQQoC+k9+jYW6KikJt7uRESWG3OiGqUVvpsxp0UFIfx0r
QoZjVzbN8FLjYwH1wBWa3T+DjiJtaSQ7m3NRXnISPAQ/EyOscKKUx2kK6CVYb8nC
cy8XvWddx+ECL+2enshp+mn7XoIiIr0fcAYsY4aqculX8SJYWGPWbaITfFpo/R/m
RDcomB399kIGu2kdwDIwqtCFeYNXOcUDhnIkc1E5wPKzxG4jTYZDhmVgd4Hgew+b
Lg7wQ1EBjI80HTGnn3wygIyaYb0iT4D0+EZtm5yOTpvD91dbfqgOV/QMZecdR2WL
/hgtoJjAprqYcSKFNJzjSxFjS3lEr8i77Igi9vrNam4mh0PfhSNtnuwQPVKRvPNb
t+E8SLsBNmU/6YRgcJhvO38028Hwkx8n06lebiK3WDkhuVwo8nG54Tjnls5jklz+
X3vFUleM+RuHxhvXk7HLVrluxP5A++QR2uDAeCCu+JulrhVoarpcXC7fub8kwLvb
TGQ5NWP45d9ejMDHA/VUQArV4Yn+lv0n3rbVd9/EkEyX5B5KU/tjuaPa6lBbI6tD
KIBdr2pmj9GZbPJAtXFEg7/wWjVgwaOcqRNlmEfDrd3NsbiulcBKdwvPkA2enZ4J
4WqLbZMEsbqEjgx5Nt6guEdswAQG0Ulxe30BqcB8sVpN5LyFNEcyNF8QLAVsR6Ek
rDFoFs+bmxOf2kfHrvsv1iuAliORFZFMoelk+mSzNvVP6nacGWtur6tXo+W+rPuO
2rgS0G13miKL0rCRYRG7TW2WDtqoASA7C6XOAsdowQKRkYZPutVD6g6JGQaof77L
rQUHnBAsPQVw0pbHzdHTvP6sO3BEmlqFX5qSKhvsmRMzlfrkv/49bGLR4cF4H0pl
kgQtq/3GzPgx2ioAAxTHRJ0lv3hjzfOYHw5/CZXnPEpUS5BDIxGwg97rlZSSFS8a
JOgMteUij1MBgC2XaZOEKw0qvZ55eB2WgBQqprDmUSn3H13lPRF6bJqMeThkEdo4
R4rnl7GBJXAPDOC+BZPOYiOytwMcqzf9ThJt6kleHUBmOUwdC7OlNDtGRoB6TOB+
DY3J2xjPVgR8gjgVnLEGhCwL7KgtKlZhe6u5/N6m6OPfweywFmkEt4ir8REqzvDj
FUo8Rde3406BX+1ZsPP4oU+XdHSofzdzX9jhYkkabNv30iWxOv8V+YZqo7/GsLBA
WhIMBOxZhjesSsSlx54TlwfvqgohDOKoGlOJ0nPYGukSe09acPr4A1uUoHhtMFiY
xOYOAP62sld1NvS/jYOwbG9kO3IQksiid+t7vUSV1pttfq2ljX3jAtswlfFmA1zK
BeRXl7NVMBv7dB+dyupOIbSq0AWSng9Ev0dY2MDCfBivzqe+up3dB7DW81V+fyW6
vx/vSwRz2/yTvKE3iv+UdIlJdSHr31m9/o5kfwCzZgHx3jL70gEbGxDZzLt9IS/b
h2iuuxSPu7T2C2yBOjo5C3NxnwqEVvX4heH6RUCmZxvio2+OUbpfSZEYfoLQR58v
qq6d7cjQ8ifWZi7+Trn0jy8nK6nFnsnNU3CUvY75xzSVXgMHwprpCinlpFWVyaOe
uMti2fM5YMHRgzpS+grxfGv14GVBGNK3cNUBEhYskKvgqymP7Cr+RY8s9N4mlXFV
7kAb4KK7LyiZF6Osj6JKSCTyjYANqTrdal9f/7wVK1UuZEo5sCjcDDahFoX3pB3I
VSjkZnQoorCgWYysWNXE/aeL5Xfo70a9f4QM4LQb0JeyRyiXFnAPRiLXIykc1Bzt
0awMy7ezyCiKTsJPHidTRj3qgUOgrC1yiJfdxeRwjZOKM1HSfg5wttfTS8IMr5ug
PuuTseY7qWNDLfHYwwl/wRHg89CyNrb+t9o/a0zQI5ARdRRbaQ6N9ZrCBct4hQCY
0VAhonnTomC7U28XZijE8TuVBuGaJybfxlGV/LxQ41q+9ib28kfYT7UyiJl7hiTP
l/UsZv5Ek9cVKjc9gn9JdhZg2HUh0weCjv8tY2tlVvklfEMSSuoa4ikV/J9pevyN
w4hL6rqSgTq/hJfnvlZYQ1AjqnbsUdWbto7keIz6SGGMFLjPsF9aPThaOpl6yBRa
TJgvkWXa0sZoZVwpJdB9+v9VFBkUMe560i/iAcgRGwTdmmqCALUYiA34zcmcvpsL
sra61J2R6tB1/HOb1HhP1djzoZOvQsRLBq42rdTQBJ671Fom8et8qn4e+wbft59m
Pz0h14Hvr/ZqjorDdIxJjZl+atKUuzixOptkskCp0uYeOGzJZMSMrIs7k5xcGmQX
ipqzVriWORZtrHnbEHjraQRvWX+tNo56L/JVZ2OcxlvOxTwINTZyZfXegoL2fDLB
uf2Ywe2Gr8Q+K86yAvlonNK39B7vlOuh7ICo20IcfwwOV8QvvF9RO6e7kxBNfl0B
7THVbAngC46VE6zQbOhaDKOy3wJygJZx2/QnDIaYtticeNCFRBN8XOweUIozK2PD
A27+6KCMmQFYq7O2goPJzq5kmm4IV4U1BdEskwsCRBBamLGL1UDnFaLbm8fVGH3S
oMO48neTe+UGryDzB0AlMthpgeJk5AIVmH3S0q4DCoQN5mHUeZgUfjYycbR6zkI8
QxQ15WDRHVp2YC/rf/8dXqSQEtMakDD4cyfMkzYBvy+wP/9bWtqOs2J0u0ohHFXH
AheKPohfI8EY0g9tm4fVF76yqb+glziD+wgy1cx7XivGxMpNT/QHC9AKiuKYXSJ5
s859AL5S5Qxd+Uh3Xpu4o8thlAkZMdxJlOXERxtTTtjIGMK1ZlGdbdzwU7kFyMpV
xtbmHbuwnxSivlKQ/vrifYlMraYLSj32mVJWY1A0sUJUe/XL3dfy8Q9nWhadCG2M
1h3Lbvu2w6Lx8ycewMrrAThH/E6O+f2JGV8zrQvuRDHg3MZhUe5hgQqnZbpVM8Xu
fx6BmdT72N+LR3PBdDDGc4KFhvkcE0A9fKEHnm02WBbxGcimSSbmG9t/o/RXPhVy
ovDwYPquGoed5EOdJtBBeZTSHsUeFs49K7hAoO980bYPY7xer5z+Cz70C6WeHH1C
rlXNcB9AhAPAgMxtuCxWTKXwcFtMaS8FWAhIlpAAJI2RCpCZrxyygZhiyYFe38oZ
8oG5OG+yy2bOjNuTHWR7rTleP2HRQnnidzbI76DsZTj3n9in15HM0l7yVHkvcwJZ
qcoxXUwMDHqX/mILiownUyzUQ63twPkCWexmhBOedpf8xxh/mAx54OVI7N5YnRlE
FhMERMXVhkLlfGYs+mkFsr9jHS8PMBIyMigKw66Uy8cbfyU3Liz36qi33dRMsmwu
wv09JFPi8XiyvicTOcKEvQ6BcxLRQjqrCsGtJppaZnnj892IjXeVUl6Q8OTv6Atq
5Lns0a8Mlc2EBghmQK5ct5GQ6AXtHbNzIuWxXc4rmEoZSgHzyLJcrco+wPH5SeU2
Y3k6HdEGt4J9trc+DJGIOChoU/BWj73zL1KCKSBEkejB3bh44Ty6V0xyJtBE0VGO
Pxka2JHp1UCHqNGh5I1tgaWkvCb2kqXiWdDIzFxBIBapgzwjRZ1b3STUmdX6G+2e
NMtg4cHm+DJNbLA1noJ9jRX6GUSQPasv0rKysZX47iLTsAdEguKQhWDSKqDTVgG9
WPhnSAnlX9pJ6RGDv3HbTqh10K9pYwTtY1LCiszfM5qBEpfojbd7YGfyumErOsPH
MLh+4FwEJDLoZvAYEZZb1NF6tNjcNTWlZydbKqbuIF1GTRFCSCvtne3ZiUr1EFcX
xDLxYwmXJV/fY9aOgLxRnkoIii0zkXrET+fiUmCCoTvs0fZa4/ZbHPk1V8Uo9JQY
MhnMa3d5/4QrM5TBIFYDxw==
`protect END_PROTECTED
