`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kw+4S5yYRwek5RgN+Nvtg8uQBH6kI7CbRe9Fgq/UPy8UClbJPz8MK5unk2Tz5A/K
DrO1oQkZTTRjvVXXgzjSnCdNkk6L/HzDP9Riakh2WALO8bXqO+SRpQlT17ovKgQy
wwhAFoDS+7CmIrusMy0P8kQzvUyYknoXrwUufS9n1fNQZCLaLquKCiZxdSmJp3Od
Imk4+c0FjlX+bG3/iWKY/FZefYDXkgtB4w3iwm5PoKHyDirOg54sygcofRiiXR3e
qFa9pgvJe2aMLXPHAGF+sJKzw7W/qpyfGVdoEMO7k20eKS17HCBlB9HPM47dVs/8
zJQnD9He26ZYvpdagSb48pJojbDSCOHnU1HIe+Q2K/SB8DGAXyoKM6w6et46qu7e
+ST5abKcw0t9p5p8KTPcIqEKTzTy9PCfJ54ZtU8IMYo=
`protect END_PROTECTED
