`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XizxOqiXQ0efj3WgiVw2gTdKwBz15CEB0ZkhNKYjPgOOY5XuLTr5Oz5OfdGBmVqA
RfQsq9MhweCWwpyhEErz52la3gAh9TMGa4zGCC0E8fRhI2Jb2yV+Y5Cjoldd6qxh
OyYByzzI0BCOGHb3lncGt06VG2rKwdYkyrsbzO/x9mtOHz023G552vNots1thCNA
atsXpH333649QSYW0DkQT/LRF3xWKFdDK03lK/nnx5aFRDZEx7ANej8g1ntA5DVz
P1YVxuxkulnQd8wQzXrGO2ZPxREJhRWQLjflg8v/o/FqKDIrJK0b6u5RpttwpBTE
348oG61whqiEzj5nPti0Qa21S2Yh0wSO1nqhOBkpVlmaK+EWwhKzfIq9LFFekgXA
`protect END_PROTECTED
