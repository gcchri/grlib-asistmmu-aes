`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HaCQGZYdW5a5JgJYGS6c5ilWhg27gC9Xc8/WNJW1BulGr1qUDj/lpFybzrRCW/RX
BfbfdUmta5NZ0QRAmLYeA9h/IvjWiDeoh6GdycMgur5viubpt7LQOB2+r47B2its
VIba5dCkA7rNcSghFsf3dhIPmJAMlfV2pZCGUU+xF6te4Bixb6qHO2qCmXwxBA6/
D/beAR87c9U7IoMkHeuJDSbgcIm0B5JVNaPPgPlu+OuX50r1nni5kYxTRYa6dvt6
GqsBprwBR9lNrSgtjL6xWeuEXHDyoh6LIVpkWK9vMvDmq2G2X4XBF1xlz1ZFi4uW
liICMq+AYjtDHACmsPiV5J5/O6Z+J6IOshsSRhOtUAQSvSe16oeykSyDfAnFqQFE
wI7ucuUDurg72EIri6jMN/byYCXSvTmM0RrVRzU+7OqsIy8bI2tBit7LWu21Hx27
dsMOnh/2eYIsXlmy7HFKFA==
`protect END_PROTECTED
