`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xE9349673g793iQbKm4sd3eISBPq6dRJZtsdrZoN0em/AjR2LZBXfq4kZgIQjXOp
2P2+dQIURQr1+LKUFi4LizDjvBwEqjKBRLwIYChpwMhiV083IDXtwQUzZfAA/Ifv
bufwhZQK+eGWuD6CE8vktBhONo9aTtf14+rM9aECVZibwKg4NbhhnHzZfZ4m0+rz
lraq62Sap43wRQyp/RuFPom0gZS6GAXIVcZ1v6ysPxWryPkuP/XLXuWDM6SI//CS
+iGh93m0mXk8bruxnp2wNJkLORN+yc6lXBOE0b0UJk7zcWP6cx5ukKwbFPMwG9gO
Wq6qaH7+Ap+uOiZFx8BJcZtGOZqi9Vq6/QlNVQNnXkR8H4fh1edFERTrehw734RI
9SrOCV8dMx9FnWEPiseMKR2bp1bd22o5JInwUOG7+dhEY7+Azr5L9xdln1aZ9x+3
TQZf1BPo7lGwMmrcc0SeTTbfSgUxwGiAoRCo4eDsr7wNprewJiB2SmJ8CRf/meWt
`protect END_PROTECTED
