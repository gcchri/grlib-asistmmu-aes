`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MKy73Tbknpx959RCgRiXG6XTxs3rDIvNZUnBsmtJfh7ZqWrpJtYJ1e2dipV4dPI
lO71hs3dSlIfW/meLvTFsZdLUwtcHhhXbY9S08VxhhdZN7w9/o+nIjVDv1mW/DGy
wFMlL20SrcbdawJV1y5te6c6EFbkDrKIBXZxU0U6XpqqKOldYL0BaK6Ck8Ir/H2t
eN1W/NE06FA+R1WJk1F4ATg3bgxh2h3ZF6HVWIFWkYA6Xp3aSwDnPqYBO0X1bajp
vcMqI26KaJfc3tQmwEP9ccO+lvI4QS19rxwtZxBZB0Cs5ms+vslx/7qYeQXqxH4n
gK2RGc5biwk7U2CVXcwGbcYIb7/b6LZNBzp52CcYo8s+INQI+O6f8W9W0BQgWIBq
cgjN+Gp5jwr7hJET1NoAV4FkvHR763DlMhZ31EwLXpMOkqdNbzSJXvJenpkPMPO5
9XCWScWvWRI6HnuBcXkLLxaKDgc57KPtupOHe/Bc0rM+3l7vZ9TlBpzyeplkdn/w
KQYmcVXYHA+YpdtUx9WWHVWGWWaaawn/aFat/txi28M/nvpbFgLoe+WTcrxID1vF
`protect END_PROTECTED
