`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjBccOBolWL4JPLky//WXI+spVO3AcVLoQ4BopL90i3B50seQJHPHa64/OQkdALn
U7tuhhIk9MazLVf5oEQMk0fOeVHTNgyjsekYs/x/87A2phIdKNLEaM18ulnP/tu2
C5yDgCTcnHmCngzpoppn7lalOjeajg915Wnz1DhDlByyGF3xyFyNaKm+j+rPT+mR
+LZxpgJGKvuEr9NumDfY5H/r1DLZQVp3BY+4+b4f6EwWjk0OrzQ8yqtj8P7Z2Axb
f5N0sZSycmzkqRkcBSG/iCWFhGnGUpjmhjYgGNfFmss=
`protect END_PROTECTED
