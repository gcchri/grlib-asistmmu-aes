`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1FWlNBdL86k57UNP11FkpHZOGFzdGti30qFHc5ntPta6kYfORFxUksPJcfqe2gcM
ARDb/0q3ZvI1JhzlXZipFr0kQ7+1vt/4p3yVa8fUBt7rQfXaI7qFYQU7PNKvdvTV
8Th0xLxxUX70kvE6ZNauxTldxX51Yco/nEKx4Age6LOTw8wYAPhbZFtA4vCRmPle
wJKrLBQPXkGEECawDFTLmHaKx2voCuCfFqSA0K91MY+GODmNPLjHiDwnb0cJothj
4xG3j7ShJLUnKWpDAk0/HTX/tSuI6dTu3dV+WXekkuSFvgk6EPwsey0PUcRgPZuv
JH3QCU92HIWQ5nOMcM9FtiqBhmjOOmwJG7MiVxdWYemyjYDnPhtS9V8qmuq5DgFF
vZkuOirtKoBdzBvnnCuidluSGpaVdgp8T2BX845jnZoSiHOXesi5qFUCGpU9CF8x
aQumfDDWlr3BJZsfWowaCSe4m+U95kG/xeJ2JAT9YNIFtdLMFGcrpD2lPwJnFdAW
QjhnESBu0IT7LyB/Sxe1ZRWYFWN/Ar1GsmBGvK5Yx2ju73oxrScwuwA2UcV+D4Xz
FnYUUzCQd01WLgI8Yw3dhOEBJJBuSBO4+PAPZDmFzFSk7XCLqhLJKnpdFp+7mHXD
OCgJ5/Ag5A/dsSf8I2xE7zds/V03BXVBZc68cswljYoRHXSrrnSf748a/pntGlNj
83/0/CNGbiK+rHgNMwcXCkuh1cWeAlGEWFTA56Gqvyj7l6oebFchycgxwQvQIjwh
CgbV/YBjwjY2ernN7/Vyu8NYW7QUKrC9sAnGYM6Sn3fG4wNf5ScixRBGR8GGw4H+
sNwxu6SZ96LefEnb+sbfdw==
`protect END_PROTECTED
