`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ROJTYYiIm3mVz79dYvrVTYYIxPkWrm2cP+hTgUwaVQ02N5//eonF6QdzGihiZ9D
3moShFalSLH68SqQFREoQ5eEQA+ctYHkKrWEnML0W/5EoScO/YtbtM+d6BFSoFMH
YO+fwXfkV7k8NExR4bDXF/mAiHBHi/H/N4eWz5MA8fkIIE9Yq8ROYN49229jD77D
OM4ziNBFx1aZlL5uzZtrW8tG57WV5BNJGDrohYniwl2LdLtqOMrRjmiKvdrD9Qx2
aQ4z5iF+BwT65KXyWyKXKkCHe/5+XXreuizSV1PYZWmjYH35/2amFU46Y7BrAyWS
RTTy3UEQUK6my13skHetlmLcw9oWBebwG2BLzpPEU+PnncOyM0WPdp1wudqaj+Bb
pMOCFmr7DUU8KFX4lydCFbwYwa02kn8jHZ9tNWPDCxQ=
`protect END_PROTECTED
