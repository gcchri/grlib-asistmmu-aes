`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdHRZgQZWtIos+cnBWsqWXiklaICy3e5qCdIarzQ+tHxCsau/8PL5IS21WiYJKbr
uWlefy3rL5+08ZamQU1O04btFhJTDrSA9PRtZkO64cAThfNn5atsr7+d4SAvSyA/
eNukW6VSi1SKUmILqMLsO0YjZ0NcEs7UN/f8V4bW7qvpommAGC5Y6cvT8/E7yZrl
Y3IjnvW88gA1Em+hNXqHFyyZ5vfkST7vKSMbWkcc5opOw9WUh+/gjmP7ZvWfbhW2
I1hLrmzmNx95gO67xq0zHTTUjrKNWrtzONKEOFKKhicDr3Boqw9qLHOw+rXUM0OY
z0riB7bHG5AtlF7qQ6Pl2qHxtYgenCYaqjB4rhLHHUgnDHPSerYN8zvawy/7r45e
xTlC2K+G2d7se8yO6m1syb2u0YdWR/uvzV2k6qf7URPx29y0GallrhVzDPtdARho
81zI2hJSCotux1DG1FgnSgDDuZhi1jNjrJyH7mkz/mannQoOPX70uVxVV0LHLDKF
fqW8zvlR8vPO1UFafTpxrg==
`protect END_PROTECTED
