`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o2z84aFzjXRXoEmbnvT8uxWUTLOuU8f2p9fklp9SG26EpMxaGrtO8XSRrFH7MRrM
2z0QhYTBPP/p1Q4dXHO/Z8D4xGJ8BcX2wXzwhaCKE9fgNGvnnbtNBJUFdjUHeoTK
Q+amMGa2O2ahyMfo33ZglUXN6ud0LoJ3uTRT8GUD4kK9DbduLeeku4RZ5kstnrfC
N5+KKqiVB6Oycii91A5EoAAgKH9eX434NYxMBTi5D9Nn5/1K71K1iHZk9sfOw5g2
VfL1FlJhFlyyli2SKAXj89HNp4qa+qvyifcl7bLdQQVhsi712FQYbr9kte0lYA5p
HEjmbTLcK8FNneEDYhyKvWgWxDV+PxrWusVWv6wHhySWQeKIK+vc2qyJ25GrWZ9D
a6qicneE8NEIr3fZX/QuvClx5z6OxQDqh/O57lMpEouoq7YybQ6cjpA6oA7m0g8J
t/kDYoFjwXY6VLGMYjw12Lo11ktWUN1ANZjwBicstUVzxnTdQJvBHBoyfkoWxU5t
q4ZdBKXMH2hYl8Ty3ToO86M9fFuQ6ZLoK3oTXLweHnRNszgF8bF0xKo00fXv6rba
lOfNhSBULLIOHEim4G18aiLjGyTBJwetzdig901HVRqoxI74UBtmy+7Oxl0Y+jQ6
ZuBD0pc0fFs1lb92CCz2Lf2T9bKm7sZ1m3BC0J0ZApg/6qDWCtfhKPOJVSDxF0j9
`protect END_PROTECTED
