`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FoC+dwbJ5J55J2vUJFmFbzw3a8raXsleo1mo2KLaCUjZRa2Npb63fNX7zCoyFngI
9/Xw1xsHPK3NJSFsNpbALapAHTh61H1hU5byr4TlIAClPyjEjEfX69tGfxU9UYkA
sonlWKE3MtMx03TVDOJhzRMUHpHT80gwZS/TMELyJqkwe10D97Ken34iKiOSThr3
1BIgVTzNFPgciVUWIT1NvUp1JGyGSTOBv9JtPA9iEjlAiaF7esIjVqZgNDYMC21k
xZd9yY/UyL+SgcEK5uuwL4O51YTQ9rTGG2Xc2cH72QYynTdwIT62MgM7hTjfiY2y
5rU1bpw4j5SxHYidJsIpPzvitZ5jziCF5g9AObuwDGVZ9XObpBoYauzoNpJBPrx0
RPW8fDv/6qgzQKE+36Yhq1kvVC0SUNYpeZTF44cPOuOuMeHo8nzRn1kkySouqLUn
OmzNteNPzkc0C/IPWCCwlobxI3LIyJRJL0uKL1NQ4dG5iYXvdDmZ/yCmp7nDu1Hd
qInzo2o1pME1GJ6O5potWhBu+yyM6jZFrJgqSnHbgupOkVnTDriAl0G1frTRciaR
ltMvRqxgst77GkzjKIliMkZFX3UQFAR8Htfqwm6rkGInFnPOqPmCW2ArOG1KsRzC
jMlABhFZ7TEhekl7epKpzwH+mHl81lfYXryj4a0QO/ohNu77e7BPlthzi72r8XNV
CCEgHg5lQedPbbn3+Uswz2Ud0Seyess11o10djc/6tURqNJwCmQNehZm6A4FnuqI
vqfWladUuvhPfX/2mI4K+dkSy8aflN8+np5C6x8QqyCKgWZkdygSB5j2UUJFCVFC
lx2vZT8jkdDFqrv7iB9/Vzyj89CGixZ5Bf41Z7oypCiAU2aq7SR6zy9Qy39tyJF/
ooaW7E2T7JH/4g540DJ8HD75mK/n9OrHOHKljCgd0pKt2R23Mda8lWPluj+NIVSV
hSFkkAG37qHW0vDKXVfFvfiiNXfPObOBna7/3vYXSuWlz5tS+bma32tqjMc2J0IO
vLuhpKFEvJcI8Bkq6+oWeYkwA9NwtU+PaCa723jxH0WFJf/axTrm2upykdhbllSZ
Vh3ZqJsc+Ua0H2gGdxwZTfZ4R7rBaVrzB3sWGWQAvovfc6wNKuRNtxrBNAMYv4bl
o7m8vRcU37SxObnFbxu6E+pVpYrqw6rjTFYoJKBW41FVMdFMhsfAABUcr4fA5yMn
M0wLOkmp+FiVSRiQLZ831xwaJj5bMlrLn+tnn2mSqasuX5ClK5++vg8vaZ9olIXG
5oDpNnJLYmX0KtsHjRKaodJcibiXUYjPZlV8pW9T6kOaCXjt6KU7HH6iDUyEZ7VK
xl7vvNgTP6BGHVkb+h303JNr4rISjQ0cSezShASgtHUg4DYEt3OWp5dV8bA28LvM
+CvTmq3Wlaw81j3+QL5J+kI5cy2vLRIdg8ME1eaLFX2HX3TCAFzzgIxGZx/FUk3R
GkwCWiiwB8kmZbM9vWxTsRcXgtNWAMVaF9tEWLn4h0U+8+FPkIx/ga3qRcqZnNg6
9WJ6/JPMrdRY/Koc4Z0egpWMaacYaJ8BsucITi4iceUwgfFiOyJq5SsGD+xQD7rR
Tfw+NnYCHWYLaMCU0EB6aVyJhX9VaalK4IxTH0Dn54bdovaaSRwG/llLv57W0UUQ
OmrcxWA2qx27940Hl3vTgMAUBOLuzzhL6dmZyE+8Ny4jCYq9KhDVN3kkc2J/OcE5
F+O1JvP8+u/2kc+5cPw0V53TaiCIUp/QHJtClHw3oAgDQeCzclC/ZVbXPtAQHPfy
4OjpfaKq1zLnJr3Dt0NISexn18fY6bC4lbdmOF2ELwGChUCowrc68VnO+NqxtP8Y
JZO6xuanWJSwyU7eKSm4lFOZWjG691ft1+QmunJXFq4ESRCKqnAEF80lFMscFOG8
TUSidODEcRYYh2BrHvh8O/WQNBVo1olJLutZWYanAhaP/4NOIXZ1c0yRx68bzKhz
HjCyhpot4TIshJzG8OJrKNVu2tLryxoYuaoUtcj5WeeKVmKEv7872pSOrBFX0iPX
cOUM1XUzm5KVdO9AZie9GlLGDMrWwF4PaZnRAbJiW7Z1qeknDrYv4wHoThvmuwFG
Xcqjh8OZJ/9EPuSpsEYms7dJEJfoSPL01flnTAnVsBJvZPallmP4u7ch05uIvoSC
02LiYnnLO4FJUgTbaV8cGAJM16GcbytS/o8tcjqgToNNXiLIENkOfi7s4khaHGiK
YY1JLVsjOqvMfx2gvBeRF2UFWNqBYSotcrP8FwI8whzD3JgfgjjXGgSEAr5ZJIIC
1Noeoc0wzJ/zSGHZD+QbIPunIPBxEFSA4DYApgTQDvN0RPDCrRGcG666KOAI+eLZ
CkZa9osvldPTn2rexgX9nQXlQktRIEON0aqAfsb3kw/X9GdMzcleOqpiOrGfn9Pa
xcAErEO646rVvYCf0U6DuPbVlJVC9Uwfl5Li6VLhJ+IYeDzJxgEaIWqb3dixN+l/
1DBh/i+DiEZUQYTgYwGRXMNhXWkXNgAOgP70+IqAe8lI3czJzr+ExdRtwsKm6DRu
etwFTjFsZSJjPNPWN0z5a+O/2aHyv7W2xIANF+PpgOpeL2DetEElP3g56qHOzqvf
E3lX+iCNMkvIyZbJcxTCPoj7osfWcQPPwf3gNJ+WqtZObpv/ZaIsQWrmxCbeiFKw
uVxqERCpQmVGfuAT9pJjDxDrI3dIi07acJea9Ou5P/pfTHiNRagc3t31XEWCZm7O
kkjBWafIW3+5IKpE2Dc9FpjXBwqVpwNT9Mjg0rkiEgLbVbhWaAYaC3la61v4ChLm
5N9pogwsz/Ktgaz1ojekH35n7eT+jcTlzgEiltF6bY16NbqyxCQgYneALr36SkDb
m96D86FAlEVjx4iAMK5dA3N13hMkfjaq5t2n5EQYro3qCEszpsDVEOW4yF5Mkqu/
XnqjWhRW4tGHsDKIfeK3FVhxQ3Ex1SsFfUj+32LLlbUy4ex3fXqEh3iTAb+BazyY
833JPGiPe2lMV+xO+abd6tRGh6bqeMEd7Q+EsXP/MtcYpS/OHRQu7s0I/3SPG7D+
Bsm2698mUM0Mr9Bse1y0gztfL7ej2CTBPbIlbt/smIGdqhqwNfG3h6BNXxN1QE/H
KPCTurBy7riZD7bCq7adpaqqq1tdzPxSrUJvVcKEI7KyF770U5+uzFyMPplVc0Q0
5WqulpRwRZO7wjKm562/DTY8HDuweMpr3nHqhRAOk5lKZixa4sTDcl+pwkfCLdgQ
QfQLlY2lqAH75d1LBz903WWXOKEOxG80JrnSHuyqL57Ytd0iQLZOn0QtGqRpYl9S
GOS2R3Dr69OqDr9mgslSDB7J3xMJAl3SNb1ppdAf8DXZQIytgMzNuwQeVOL4c6tj
WR0IS3xe9ypntCyEI6sPp7GAGuRjCTre3gldmhWM5zxM1VVs+qtliXB3h4zME1ug
ydSRK2GlyWK9SMU+GfAZTVeciUbUJ5lcStpxFzhytQM0pD+L9m2taOAPnoYu38lB
32DcW81zZaXmuryazLJIkCDnNVO1LWQdH+N51I5DD12rjzhP890C7swN7ywvEJTV
H4BmMtDqQvvOjPBLRPv2hSb1VYUdRq0z3yuJqlBV7ibWXucqfqmexAFyOoBNbPAM
REXDOTq9x/IVr71hzPqjR/dr0K5f39Jzh82j3Vc0vGtKiLLWg29EaWupSl9Hdg84
GSl6R1jbWFd1S/+AbcpmaJbP+lIreJOikyLWvsfOob7uXggcTqMUVVHx6KLf5ryX
rjpt05CErRHsWtRNgLm8/G9DBB7YHTd7H3eiCFHug3/sXolpk4WMwpZXfvMMt/Tb
OqorfvNsM1prG0T4zR/WBgpwkrbkhHUH+k7x5IkB6djSx5/C0shnxy+NdESa6Fyz
J+Di1B/oJGzY7nzkkNr1tUfuzsVIJz8qHpgNNkd6AXZf6KHsREuuDlRNjTd1HWlL
Dfl+jyrWG+HKF3t4kMwj3IrBDDDDItb/N5YPUXxrXXHl3Yp+/W/ih2aCemrfuxMG
ENKaF+QPE8asjv2kRTGD37zDzkhA3jDlACFm/GGS3DABzOtWviTQ4RHJfLnbKpGC
tIC6WUCK4IGhvQYh3EzXX+yeF69XKHRSgSe48lMK39gGAxPmmjYov+yU6puS7NG4
S1dzuDGH0IMhE8ok5mCISkNLjv9Hh702jaSQ1lq6TBlI+LyNjYMCqUxToIBZgAbQ
YbebwUE552AQz7YiqDMiHg4ThM/jvQHYymXIbHMUfRYVMiQlTkDq8e+70VBuT4Pt
7P3GD8D1slH28CpDMxLLcArVbEO49GmQSALcvVo/npZgt+DHqZMU4Fnr/2fv7gk2
YGfN9RxxZQYiTXjsWzvzagKzZL17j175HfoKF9CuXYlfh86job+DuJT7oMb4Yp8Y
YFh0VG01TpVzLRUunOYRzAzPtarazVqxmdcZAgVulBcFgbHVbtCkoWIVOcZC91GS
RYwNU4G5IevXp/AxAPqfB2PLu2hN+w6Qjkk5o7LqHSrGGqhDhT4NOgDFtR6WiPJY
TvZ7VIebb6OpvZy7Jwy6FCBi1PFRU+swCdKzfX4SBYCNq/xijIWyQkPKjemltwcD
L3W8V+8VS7LkF5JT+XEPkxOpQ96YL/oeyYpxJkTYSbFlL2xtJ9CN7BLu4mbBr5qn
kZiMwdqISDSrm/85F9sbLz4nDKhAvXYmBJ/T/+BmllE3xQPalj8HtwZ1ECNq7H2E
pehTBflN5ZH4Fqei0tmFKYpM4ZaxP+0Vw5LkP0KHSm0tGzXnKopn/5lQoZLGMcI7
d7VSPCvtoxJt/l1Cs/tjU/LdYUCrxWUnY4v5J1pGPL7M3GtU6jhrVijx/GjdfX9w
n4Pftm0KjXuHBhwQoCOgn1dYem/F2VDwFylAX3vPDKY4HvyPszpJB2HMaqYjcC6l
Jgetz+ya+Zb3u35ImOoHHyEe2ShbaHV0HOboj8gP4USV0bWBfAKhE9Swxezqptis
PUOGZ0ZwTPAKwQw6QVzdI5PoL6yWG7Qffv0VFdvo0DoAfeNum8DQyVKgpH2us+Hd
dUk/ObXKPwaqI6oDNeddLx09dDyE/PCD4hRImwr6z0LYlkDR0h3t1XVpkwjlcFpL
Sv7yN9A7ztUTKum8RjpbafyWOC9fHGP/6dhfttDJLKSx3fAA0eSHzz4SWBFAqEQ/
ScYoX+QLxAn+W/zsXiBGrj0nQDk46yXUeAHoVtrGML3TGAorU7OwMHd1DUJxVvU/
C2g2RjTK8LZxWn1PiiXzrleumDH9Hr+jCZkGlSLP/eRb2XiBKLG/BSESiyv8w/au
ux2Cn8rjJu2/pSYum1Ty90uhJRudiXdpTBJnRnDkma13/daGhYpOK0Nlwi7J1r2l
gFLQZ6nlHaagD1JL6f83INAOKPM33wxSYrwjZFkVGqWyhfifssyShWbIl2Gt08EE
jnkYi3X2zqi1Nwq+09GaTaIJDNFQ2V0laDd/fNaUf7DpYYMLK0cCl3hh+xQ/Zy3T
G6fw1ybBu/Ho3EnKWJ9wZWNt4JBkUzJdcJn3MLEEENSqYQj6KhaTg7f7BZ5j026P
UmMrmhtUsIj5AEdF99rIk6+R+07odrGwqAlmZtecdCkK/4nmg0abIYK2qur3cv8Y
KJwXPhlVFxIR7Kd0bpls9EdjvZIpqgQCZZ89cXrBxI/5vyJ1WDQIgfirSTPccP8m
3RI6AO2CjXqAnOu0SRkzFxv53thqFPpajEGCFYt+aUOdrseIia/clbcerJu1Aw0S
w/jsKaKP41Rr89biqfYCrWMvONS8cEw/y4IZ8u8iqamln0MSt5R6MOWSLilZHIMs
dtyvjpVxUaHnusqpLdmdfn3dEXv5TDcXAIouomQZ9t9j15CKm13HY9RHvLLhVqeI
/nQJYp5v3LtAm+EEoF8hZI8nuToTY7UCW8gUYrSiMy05vpswWLNLZeXZpfQf764k
zHI7yZnpm0iZKMGYJkt97sxQEwN+ww6gm+Lh2Wngx04mYT4UULNI35ux53NvqE/c
SkLroLU1OKjVaj3oPMUPB5qBnxPcBlpehNd03JR9oVO3z/MdutRqMXecZalModcq
BJke4XIyvinXzcujFf136bH7U49P0miWnwslUFLH6FO5Hcqwg922sBINM7QGPb9Z
4BxN5j4Z17RYBACnKCX+9i6aMJ/i8TiAx9CZUXbGFRNEOqZyn6lwkjc+DYWN8wY4
caCUgCYqD1B6mY+OC5aaGl+f4Wyi6sQXtK/Jl+ReHzblOyGF+tlNxW0vKUR6fNB0
cZDO38YcKAOg3cngCy1gjVG0G0WfOKypJcbhZ3xIqMHmwL5+flunX4bnqHExl/Wx
CsMQs3iGCsdJDZBsA62S7Aufm6wiY3KY2WMJKkMx7eTEyBAImDmXla/76ZLrqo1g
YfqcPOkvXQdsgXWPbHs+uUO1prhC0rnxlNUUFqOZdAkgnlSPoUIOnpTZcIgjGsOn
lhMKLZUVN4hMYSkj5VXXv9NAPNA4vxFW0H4i35Cnt/WrnUzPWtkCfkc92u5ZJSL8
lgn947N5zMl7IFyVrh/MlzwUoS4f5PQivcS0VhGaFVpJCiBgaVNFabd2XS8Mvg36
6T0+l1hftc85MbJMUeN9CmBMLVuAW++Z/G6CAB07FyocJGatdo/LmLmf6O01mYJe
2BOqlgqsy0zBaj025Jwjq23qR6JcOcgn5dOtDZG/pxNmu1t0rxzCEQ6pMR4rm0I0
BjUnH/2vojLeuraqtAWlE93aS6lwjDh7UdpgGVk6ln6STjZUAozyRBdFKoS3SCiY
qHdWt+BqTV/qNUlWRAqB1Lj6X03f782Tzfo6j5D8yoXPlfV03mQ+YX5Q52rJvsBC
o5pnwP+WaoA35gvJdKtlGNWWnDG9PTH6AsJvwP8ktBBCM9Kvmxoou3aDo36mnbc5
wsdPRcYQCAQoi5ZvAejBcqdwM3OsvHyDJsj1Cr5t0E4sxyzTXPNZq5nnESU602w8
jcIeD4y8HGH2LzTNGMnIVm4lk2ba6le8F5yQnwH7Or5sA2wkG7Ase+JrGnV+e7/b
lL2VOhtAnVuFMzahC86r9uCo4bY6U9J8308Hm7q8hxyx5H31oEEq1bGOL9sNmC/3
Q8cmS/H2o/w4f3jVf3zlxl9a4KkjttHU00n9Ke4MwyKdx3mF6IqNSv8yiebdrGnY
T1qeuxHa/vVoQCRznKsUstlj7zoytYVK+pdpglc7NR1pk3nt/WyT4dmOJud8a3+S
ww8OiI67B7dtGbYYA6gLUGy+ShRHbvyQ7KnqiiCDkYYjk4BhBWaCnwAegfGOpuTH
70QPHws/Z+u9iT99Xr7iI4k0AWvG2eCCDqjFJ3VHem7Cy44/EHkoVER3EB6lefFE
RZzbUJXFEDKI1BD+4Ir5J2/6+Bu5r02GVy2QNXBBCjSMrTLLbIv9/+sshEZ7XhUx
plSpOkzVVEnN0GLsApKkdI8vOjzNpwtjr7WN+V+bMJgvLFha7L1LLLTE3ZRFhUQT
ePFf6iA30ejyj13PTSDyXQaQn16Is6uHQjZ8+rNnxovoI5EzmNXZbX6rngAjYBUe
Z8H61aGrpGcZ3rZomCWxCQPjshRcBdOe1E7GTULbT4UbTJD6P2BxtVafoYFoX8Ga
MPgmNRAS3HuEbQC+e8N9mdGIzufds9CHKwRRwnQLcrzkyUSdD/ruwxQS/sBZvhJX
j2WbmTIOpC4+Z6n/V/qXHWxiOTK9hQxWySP/my+YFnZM9U9tPvaYmQRR25Fs0uBl
29GmqGChQrifH52I5Buu+AR11AHQde4pl2vrwuR+dts+LmoYhz/tOGrXMQZY7nZ/
OwXSsQHHFf36VMjSH2cAlTB01jhdovSkRD8umRmCdhlAa9QG1L0ZhiBjmn14iCGR
keD+/H+M7JIVz7skXw2iaZdWRgQC6VnWot95KtsX0pGBV08WxBZIrE6ISmTZWg0o
SdxggOoGIU+3kQFmAyEwusQc7SVxGoYp6RbHQ+9dD1cR7g9d52ax6GfXCTcQr5mr
mCe/R73A8O/HImDJrwtnJsvRqp87zbY7qNzEox6vUkgekiASrs/P3CI9zSDZuoIL
+UAL3mKs3ypAYclbLA7X2clUXale5eDUFAgcC1CsKUGaltmUALAoO0c5UUu7luqf
U//vvBXRqaBxFEq4vJTrTJRbhIgA0TEvLlLHh3gnVofGQ5XMato/hS1aQ6/bcjy6
vesqhKE/l/xvFFHwOMgXFdXalXTIAFvPKpTbEGvtFMfZDJrFkiOFPSRAgMikSVjT
8hDtRG4ciw6iiQiEsBL8j5OcwhStViD9hN99Pm+ufOoF0DXJ5poIqEVaTaN0guUB
nto/407Ut/yvp1+RwwMp9ArI/B5nwybvfF0+d258aMKmWiBc4hEql17ir4xTHqnr
fGLRpfFyvGKTAUAk62H2yUpFZvrfMaPWi/WhzDRdNWmqBpPjncyikH6VHGOY9uDg
wH9vP06Ex1AFOm7S8m2PBfX5DSUm52hNw62AEREqijkezss2ukyQv3crPB+SWAn6
HEEQLvr6ZuUeNGG3vz6YXvsRxmveYaj2mfkOqmH/MHuE7Fea2T3PimNU5KFbo1TU
CHC7V6jebfcyA32zwGPOBDsOlbTPx0MG/t6HLgqLk2MY3YyYKjRJxDTl9A9xHhan
9UyubuJhXN1aTGnO5/xnwHhQ5ficd8/PJD8F92z61mdGvxxFxOqbtQyerBdMz0iO
xs3t6riTYmLn8D1hur6DTayvcnN2RQyW1J5WS2zN+JMpZ7aCjMaZEm7J72evZN4i
65crGFWch4bL3GvsyedBhAaM8YnCz95L/A6EHHUt/HTbV37ihv3D4ttlQ1KLxrrD
/S/3BhJrazfWR0ZEAuAAoKa02o7kH06QoWUcS2xAl+sBC5JMP0jCHGMtwLPkD9/C
m3WoeuSXH8f2WAr74xzJWtF2HVAATAT6s8hu7J537auey2XNFQ68fU3MlR3ujyvf
ILZovmuxK7G3tRY1gFc7mo9Dwl/T0GlVAESKhvT0yXkguTUZBW54a01R+vbIugmq
FjHjOTqXUcdPNNxBZZlMVtcLgONWYkH9GORPME1WZ2GAPC2l+379tU//vpztsuCe
KCs6L4D2mcCVwaVAP2Lbqe2KSxAcpE/12UM6wmTFidLWzZHzDCOomf6WqI+ALep0
nNATW3GfGlQY/jb7/vGC6PnpP6Be1RXrE52dASG+0jQ+Ln0dnaqcBwi81qPAkr9d
AQ78UgwIYbORX1LNfCJOjMDyiqyiSILFvJ+QtVVoOMQuE1VTpysrhSNTc61ujUb8
Jhz3pC88eERNjVTlT+UwjTAtMer94YYfYyFuiv2by4bK0MdKJhuK7hTbB2MQzJkq
MmIxRRkStMzs0fYhqUuW2W86WGZzFPCe67ts3KXud4gYi2Q6sLeM/MsY17cocR6a
oGjRrmqQXSTmaGFaxp4m9tI1gSRLm6WbUteBIDlBlf9qHgfsk8CYysZ/z82T8Sd7
TkfeQUc3RHS84Oa5oy+8JHSkpMgiWVmYyaD/lenRXkowPeUHYJuWraWs7rKAtibH
7ZVfX9HipinpnIxOj5nxTxyN1KESb81is+6+8Zb/fBYxs5lMK1+1i/qfSnkghRCn
tTdni6+H09NU2C/8c2KQQw8jpqTerN53es5WVxj6kJTKvk/LitxwVbq4fIxtbO96
mYHRYzm0Q/cdI/2PmWKJohicQ1dPdsyBpgUhm6EfhZm/PSrpYRitBtbtn6AkJMjL
q5EmWEchikTLrIOdc8TOm4JZblCHY+aaYIfB+c+TwtUrqNeZ0y2A+cJOrrHDNBDi
4dcjRnLXZ7mc0DLeXmATLyKnqkAim5dj2y4w1mZfM+wiqg2H7u3QUbkI9IXvCRxM
zNveEGN8y0XesWlRgd+7ZNTQjGFaKH/kkNX1wTYMW76kODrLfd4qpGd8SJnUaBOi
datfC2KsTakv+gOWOYfoZldLpUbLP6sI1LPrOL+7zEU21r8JXyBIs/B3u4huV32v
9bGyS0R88bGc62zYc6dVACp3ohiUAavDXhmZJs2eqLfVyul73pza4Yp7iYP+9IFo
pYk7b9PintpK8qOrMnTtbQpd8JSbSGWCRWhIIp7LbDdbEiX2Z5pUOFn/La8B7h/X
VyZVqVCg8AiwLkdKJAiVgIJo4DBvYX+IpbSE+wZQmvoODtIYv4XLOrkxTVtGJKq3
lkiGxIW4P99eQihgDlw1ce50d9CIMFKalk67W78mnfhy/R0lNAp+Md1Ks7t3JERN
6gQv0JD5mOhs2isl3Pp7z/9aSyddKhHjwv93t4yLUueuelkhydL/KtODeq6yYxZS
2z2scLfJD+t/j1qVPnLuDbcWDjHk02hPWBZsm8n+HhXT0UcScP4nBMUQ7gMS2DYl
T0PYAdTKo7qRpiA7Ej+DMO9KbSTEefygXhQ2iG1ie1asyhnUHQDty8Ren4riFXeQ
d81z0VEe+3DEXek0K7Su5kbgGcCUZzYg7ZWUGlMFceum08Sf0goKCIcu+1vn8fQU
LPRR9mQdO1bGoN+sdbIKHaJFtsJcK761CYbsYO7snwWiRshOQHieOHPYvCudPYHI
8ofSbyzROGLmnkSysUD0KyB0yKMpqSZoh5CS8l84bDD/Vs6gAnlRFGNNonqfMDJp
4zOhG3gLMPtVrbTeGw3v6D1hPyOzXGgVJ278LtIHH/7Bitjew3IR23M4Uufb1cTC
GafXUQiIWp+3gPBJdUcAeo582/hhQhLkDINdeyTgQ9sllqQJhuZIWO2szdKvsz9l
Bv0d0RNdD89pXWYdWDmn8iI5Gh4perhqeQX8VTIswQmYYkSOui1L73VkPQgEeBf7
gWh33Teesr+GS4y420I7fNWJ6AWOTFugX0vcApD2eQefqPR5GAz0zWHQvjhvhcUY
YEpF1tmN3auAlYYVInUB1CpWhnFo/zXi5d0pKB1OFF6a3a2aa34Kil6KSDGv2K5o
bVGGs5B4qFhkZ7Y+uIF9kPUOiOc4oy9voidtjyBmUUCOcsnRWpXu456zz/AXH8eL
IYmCHo4nSUlPFMH461RoymkSrz7N+7/WpGs1u2C5UPRdSO/w3LhPLrCFfW+tnlED
WVkU1cxqwuTZ9zdios/VXoxfxM+qhAKWteLmq8hTpswd9RY4Q20ergcK+33JDUEO
nAkPKM2gLjxctlGAK0yA8TNc1dkAWNDxEhJ+BgDmAtvSalZLAfuUzYYOsmQ9kUG+
rX/jvwGtfV2XPi+4Fvq9t9gse2PArvZgw+SQ1bj9BwjWW7h/DgpdE93U9C/Q3oOl
IFopa+LX81exVnlC9TAbUs/Au64+JGfnYE6afCsJ9GLxirU0tYIGm87BHM1NdSbp
prNCdLqdr7FPlZy6+58ItxVOQGNzoU1Gf0QczYDXob2qEXby9y6BFT3qKPt78PW8
onnpynNositqSRJwJV36taAGXpudbmXLUMZdwSYG7C7GyRUKqtkNOzcsu31uhs7K
IMK2j5cGYqPAUgXXiRkFBwCzXNFsFtiAOC5BCyaWMR1fK/eIaRm328xJLW35wycc
rTcg+OC6x3LjXajt/iyhoLVzUeSfRHWAq9gmQUVzMJ4P2X33H4k8hX2sFvq0M9/o
S9mwqORckcb3vfp+DaBQugMpERmKZhDwbUhTmHPkaN23ex0oJogQkVRWoKAV8m1P
2F1YxAlcbPlWQE6YgGe5rGFajI/q6n+pZuzQ8z6CaB3zlvX8VRmWv1P5ePxvrjYV
6KGc0d8ZTTx6NfyjmXR24hBG9NWpICnh0igdJsige3U6COcKN5VWmMXqFQfdZj1m
2ZsKWSXBTMEkjAubIFolFvKPFo5Oy6b5n3skhHMtVD9/Uj0NOQCcBbhWuEe8M1t+
ZWgcx9/kaOynaPdlwdreQjDKiFxVqbItkHWfA0fg3eQWxjBVvjFOIK3jR7IaHeeL
sCNrnCCBTkYTnTgT3JGovBaaf7zLScI4MrtZfdp2jhn+n0rZHu3+ccf53X8GPpLg
UJDB7FKwq0RblG/9iJHZbj86Gf2NYomeh1ID+RvkqRbTDEWEgd1AyGjSYqdV0QlE
CP/vee7M+wYwgfh6Aq5eh3AIxAQfouKt515fp0zYh7aS2j4c/H3gIy/WY/50Wh+m
+FAxFAksa3G9HOfDkMupsqAkanPT2CjK6bHscGkOVG2xC/TApZA4lQX+o1ZJ594a
4v3BLGqk4W4+JtVEQemLnrqdARF4Vbc6gEcYJOJ1Bfu7mN0uGGjqEklB4DXqYnH9
XYntmczZXsFTH4lBSSADvgTv5laQ74lulvpaOBJ+5mgiUKwR0g/0o3qX5cEJvSfW
psRns2jxfD0xxwp3DAxu7uYcjsQuDsUij/mJdfGc9OPysAVZKOJVho383fVbmAMr
hTFIcnq+6EViRfJ5jGeVTLDrL4U6kGIroXkW/bToAMyKcuohW5nnT2p9161DyRbq
+28EM2YXHLNyJtpiDsyYX+KLspTh5DFXooQ/pYMKqDguZLGydR3aFSzV+JxQbG2H
l4cveynKwc71rnjFFzlGR0bb1RwmoGpX258OiiIaUlHTy4IkdNzZhQbffBmZuaS8
Iny/CFvBjrVkNsFC/xXBe+1LBbn538isIRK+kbTJ5oJndFnY2/N6OIWfHmBPF4NV
2lHUFtEtdiotZHs9Dfs4BfnmUbOmGokZOI3yi0EBdzg0OyvDuVjpDS97r896BTqx
B+YTr1ezKZbDdL3u3nubX+gVHBQ3q/XTHA3TQjqeTfYARlM03JZ2B05CdG6rYNpl
P+jwOeLJ7viZsV9IbRvYm8Dta4SJQKzhdNDjUDGZRbiU+8tI9QVxmYLj+Znivbeu
k5WMSYtSbfYMhNOumLKl0tIvIutPAukPxi4t51fDV/oLOGMtpHnsAe8nekaFBFfb
n4KJWI0HA4+wJ8AkX4Iw4dgMM/XyjbXmBoux/3EnU2UfqWsmN/c2PwXPjwgpz5kz
qoVZZiKNWZ0z5VQ5J/vLke3IxoYmnxK+QZUNugdx8rGr2JKZLlhQWFDY8sz3NE5l
SUNvt5Fj3MV0e+U1xcH6FmYADoc2W1y3bT8//o7K0PmXmYx/DMFlHLfRLy/6dUrV
ay3zU+XfvdsE4Xv40x1d/h/V0S6uHA9dP3uculgwk3GUyfmdHbpQezPgNOPnt5pr
mmv4Bz0XJ4bQ2MDOt7jaB8pS6C3fgPb8am7mfIh9C7l/gBF0cp0IYw7vOeyUYDdF
l8XbJNXn+IgaGUFPhZ42aJNTcSraA31Am1waI+XQZrYQwdomDsE1shltGX2W4bdX
4DDinVDonlLvpCpTrT7Vaz7cbllml6okiFXNdm4CHdxdvCBOVSfTSny7pDoNsxyM
5Cvux6XJxKTZASbtc5rkCUBnnwrj3WZaWpyUzfTCIKL1MEkwex6N4AHPtlw8eDto
wW4XqHlpN2iWNrphKaKs0/6YslDceKRqdurHYGTP+eNdkN2fjQQR/7t8HTk6W+CQ
tneIrnM9NFYDWjvFkCwERTtFvPu4bwcKhGQh9jvkpyMno9tXi4DTPdpM/E81hX0j
0Y+ndFcjbESigxxRSYD9oLtKhKtiUezpPn+pzuf5Kv2sgM7oYD46ZUQpZZd2Gt4a
B5DevMvFYMxsmUMYA/PQ89GWAzBGEOyeqICkvi7tod/jWQkPnsx5Yaj51OpycpSf
5sDER28MMqROYQG4leMGE/13dfnNA8CFtMMfU/+BTmoln2oUZMjkZmhbGU0B8Fae
lH6y5yNCpFDlFMPu9gMhiFBA3WcwTrkVawnqhuDw1bmFaMBKRDKwffbasDZGlI/I
Vh1Lvdjs1lUQ10m7HS4+4l/P1TA9eKCslKWEIGGAlL/Aq2RkeNr2f8WPuyfX9UZl
5K0KS2bA7stAH8dNhSJmzP2U7p7pf+nMGedaw248fUnqX7FZghNOPCnZkBm32Nhf
qATg429RX8+cIu4LgBchp1hLHL//qxXGLFpASN7n79QKfDeGUhV8DDbYhC2/GMOi
G++hnS1xVTvYI6NjpKtexVA9jyckgdostctoOaQrML+rkTVA3lf8pY9C1nF7T/Xf
e9nqESWmF8tHbPSrMldVAexbNYk+Q9grkW4NhI94bOqGo5cKFqgB5BmtMRHLTrX4
TADNLqv7xJUFb4XaDauk1kha4sZrCmXM3GciHQsuxzi4Hv1o/VtnOZB8SNEZo4aE
iq0hmqC+H73sXiGBS4ZkV6911EljYvyCXZXun3uYE4SoyII/RKgv/Z8hBFUV9FzT
asxVq13I9YEmp4+4iDQfyRTFCeJG3hoHYlMcppQmjCBhJS0PmOzbJ4zMMT0HZ3Xt
P2CUB6eqzVBscJejE8oT1ZSgFOG9G1eJP1/97nHdCOQGfJzeQnG+nkVYDuXngah+
9gaXwYP07MmxRoZippYWcvP2NEl75aICWrLydsbdyS7P5u9Gu0fI8jBhvtpdmcT9
ftio6Xm7FryPUjYAcJJG67UTB53gehlN55RotVUV+Kp1GrqyUmyuPEtJ7iuC1K5h
J3gSG062U2Il55CAEGv3RuQoNNsOf1IipRusnvie0Dy0G3X6rmUDQ0HMNO4XAnQT
OUhRU1mSeSdwYpfI8p+p9eJ9XTv1UER5Y7yDthLx2PaB1yd7hQkoNv+CZiGKY4Vt
lF8QnjxeMuo7uaJORMKvdcRptsJY/FSJvcevBL1e7UzcCjGmn4lroaypn4hH6mHn
o1RWTgyFezamPaFnDbTO0VJlfli0IwZbEo1RTJTei9vkai0M7gwzWQHIyn1U1ret
9EbLGAvoeEfJNbWMYx3rQga1RmKLtpntbP+bLiBxTmqGFGThr50GHy8/s05Xcqtv
H3e4lo8j3n/kjBubKarYtGLH1wT/VgqAxhwQpchtjwFNXko+TZoPfuYnkoqPjSzg
dcHnQH6SQmIuPehR6BK6CYv3JvVeS8Aqe0dLBOLtIlKidYA4yTErjyBdBjxSsmqp
FQbi0Er5pDN8uwNs1ZRzI+eVgK1Ggm6S5kwnYQmbA61/aVLUfbn4HhbnCWc4roAg
q2CqsvEJeefQlI36yfVy6uSRhOfKSg4GN5DN9VvbnSesIjR96PquWTd12cRRAjK3
wnNGb6DQ0lmtWi6tiFc3DuH20Xz/kCi86L2YrS+TL3SKjSZZs/0XoC+zHdIYrhJz
4QTH9tb3KevASLUYOhFjtWkMwcFTIL87B+9Kd2yQjeQPlJmGFBKGqntFCeAzTOGO
v0SmsfkSKJeP0MaW9BwZipkoJ0RMp1TUimiPl0i0i8LaN1kXSPDO3HT89PC+p33r
cwJzPypSqZND7J2MAmrli3UOMvMpvfF2Iyeo/kaQAJ5qyccsnaoc/xXT/nYIsGxT
DVX7MIHHNkNmUD5A5HwHUXs3cT13BjHgeCFyMgE5eh/0D9ZKyeXji+Woi+T/UBji
NSMzaX83Zoj5lCFzNxcvls1YqGoJvTnA+x4lIweaheEjg8S5dWaSQgJagmWF8UMw
EeJ99KwzjR7rVb668IxlptN3tHl4TDgi08KltzagXUny4ZNWY3uaeU+5SUnf0Mna
8tTu4cdazlz0atWPpTYlPWa+QKnbrMOp8Bbjqo+2VbPrlY2uL2kRPhUKhhcgvntG
XD5RHUOY/uYJ11ROvIM8xT/zGrYX53Mo5fGhPAitN9PY5hkVMK1LlzqHyRennpyU
cucUsvBaFdGocDoUTkcgwmn+vocdcswMxEzyh3taCr0CSi82vGKsKgDtTpPi+sa8
9M++wjvwPPPJso6e+mlQ2ZRByk4mdSBLPRSs4RGNhdaD5Qa2L4dj0L5tWw985ug7
7q2IOh2L4MRRTMZzTaeM4hvlOQOu+lermJpR22gD6U+7aLfcU/HPogqw9lgZd9yW
xI1K7fyTRkHAbQtCz2pi5Pwlz9lVeGlbVOcknQsaV1y26GufWTUAVGN590vaGTYk
qgYmP8K+f7f3Z0Bljtu5ARLWfP6LSp57Sl5MBsPTzN37QCK1TpGexWkcboX5niSz
hesC1Nc1H9QREMyDOFhepRBtAzCNYpYIYFUsjL+XwUcLNrs7pPsqdvFVkQTPhXpc
btele61Bq91tQOLLgbChrruIAoeCVYwAQvtZ0M24SyGiK5iiwNQokpjlc9pbOMR6
jPG1IlFM+vF0hgObrM8LzVjMwlk3V33uKUDfeSNQB8o0iLsv64xyfElix7/PMip5
Gs+keYZUswNM1ajPs+YjkfEKTNv4Ttyzb6ssTROgBdLQeKflCTIvlTS6DvRB65Ud
qZpvtLTggNI9ZWm4sfQBvdWIYoC52JXNMcB9p4p4S4b/7/0Pme7r55P+XLCGdMaV
pj1s4Hk8fhcs75sHVqxDPY+/cGoZiOzwdmcnNqWe6ntoChjmA8vfwcATGVlm8QZH
EPLrDg7B2zNO7gBq7ph4DIS4FTKaz2EQ6hwpOc8nxoaNjKk4qBrgzb+babdY7J2Z
T/2kMuQMj8fpVCdUeWS1vi1g/yGnXjVCJmYUhZTkidZDxLknDjHMIpfu6xwtvlnT
/sC84V7J9I+5nSoocivlBjWBPCU05N0jnOnTGlGpbNOi9YrYsaKDQ109jxEryLkc
fDX810sNpoy3T1aJwNQv0SrQlPvTQ+ikqxuvpyOJhS+yApcV1qFYqu/gQKOS1hzk
92k0IhsBgw8BBnAWUp2e2IHqFVf5IwCG2zEz/4MOVBj8wSqNDNnXTQxfFWiuJx5x
OdGEpwJ3wHAy5xrH4RRrcu1l4rb4x9ypBN6DwE4jVQgoSIVtx4IU8C/qEdDnbq20
OsL1gbBqilqaVcIsC06F6fROkU/y/O9hRYcGA+u/GPw4F3w981t7qvi+Lof0Ssge
kovin2+KaFL+itv8B+BDBIYABIByMXaK4bpvVp9ktMchxFMOwzvpf/ylr+D1gE5u
dsVXFQZOHsIhlE1iRw+PWZZNR4vYoz8xmLW6XN9IDWSTQn5/7udwhY3ui76ogRWs
NEDsq6qKtqCOwFi7rHVSMVb0oBi7/6Kg4qaL8f42z3RasHP77Srp3HBGiHZTNmuJ
K1SOItRZhFQPBuyIxClXA8ucX9RBPs8RDQzM25GedRl96hfs4/N7Suexb6hmrrAK
DkdXwxaegIjWBamB5wbiGB8hjpslJsPvW0BLgy/8N1SgGqv+Mpqf3wNgN385Dhim
lqdPMmTAWjIvVzj4YH8oSp1m31lKV2I0Yyb9rg21btpGG4MjFsUtGHeAtJRly55Z
mewCINMw7s2fr+iZdbjOQdKB3/XqOeqBjCDR/YXOJux7PwLh/9RQ37RdYbCRnbs6
CKsNcKOG5qj0JhUWE/wx6yZt1VXlxsqLZe82ehB1OHGYf7iiSuDCDkxbImfH9LvF
7x8SOeqXF5VFWCsnDbt6AnM8jrIrKIqAQT/P4ESykTqEF5vGvkhIDoOGVNidDk+T
eoflh1cWQr3C99Ho4WlCnG46OmKYnG9Y9he0IOaN7rF14RfA8fojugzzRH4OKEIl
EyMzLQYjDbiLu+XCmuEeYTE/ci66+nQCGpcnrQwnh23mFntXzswR2RqTEVmatGF6
MxlP1AhvC98tKpafkBrUcv/qONg51YuxdPyaectyLEE23yVXADWi8TkYnF7k9t0l
xkv1bgacdfHRyDst0YXqNchde52byl0GxrPPTxtzwVIpA/y+oot7wwNcA0HIov3T
as8rf8Rb1/f8E4NazNTEqtiAUtsBDuLgGM4zigfuOPYatx3AVe3AyKIoBQFqiDyh
2Z07xQiyIKBPUofPaPTJt4rtxi58a1hZOjSZjFtE1I1b6Qlfc/7nDz2LLCfXfsAz
BDJfSasIzFW1VxLm+CqJzok0G+Mie6yy/JA56aWIJ0oNftidpmUBwNCca5uSQXpX
mdR+QcbgDm38d2j7zYWB5LZhxohcJHz1VfjW8IVvXmGCdS1tDw7zjtkQODpM6SO3
500dLQIzZqFJZfwCeTS9lY7mcwDBNXXmsLnheQZ/a63ybp9cmRjd7SWcMeLYTD1i
WwHqfr9zewn8KXqQgHQeRFrSNBIDaEaqJzmwZNlX0e08aGeGO3V9QV/A8JF6hnEl
w40BRTz5BzF0/4eqisqHwCRdFqxx3JlABFCY8QWEmhTACefZlRPmY73o48bCaPKO
vt19Ug07yosrZ3C1A40gGv96ArLFpnNwRPlPs73kH0Wmql23QttpFyBiat9a/gE6
X3xW7kqvQXjruJfT9I+j6O74EWc692NAvzUb8Pf90YoNgpsduCC8WhDE1/98D/Np
TId8wZ2kRYWphdvn4xz8lzhwau6cAAR9iyRJUr6WAk/awLtlojCgW4rQRJq1xrfK
EZ90qBkgcHlzUA99A9D1IN0gNZN/5ukziTqy6EhQeqoFK0s375A1hLENMIMb15P+
EXZoRwNG/9LP9jyT1cH6ZXk324s/PzgSSNDwB3uteI6+ZvtP1GECUDB91uIuloN2
o4s5UajYe9+jY5VIWFEreRj29jupgMrlBubgDlYx1iSZIeNazNu5dhzLgUuy3hIn
cqSr9RFwK5AlnRn7l+k8nAYyzIQ4B9w88yLswvYyQ7OEy67m1WEf1anovey9JLM7
LIGb1Kflf1sI7RRC3oxtnYEL7l9LngNP1+T0oA9GfO+gT5VwtStQlrJ73sLQmnDV
4mEhpyIBcFk1RbsY1G11PCAILL8NNl/7Hh2i1cnjDmgRL3Kfussyk6z1Ohqt+x0M
qItEbmCIpIcXaUb68jBBJ32hUB4QbBRHT5zTsZDOL5HDIKfBnnte10W2ges6m8Vq
K84+SZC09lxonDZ2YphkMfTMiAz57JytY/l/gGQ1QDrYQDW5Aeyj4kTVuR98u5R8
KyEx3MZpcv7q57Vc5WsQmmlDIKZEy2O/uJvbClqsLjuJQFhZxa1I1nU2963lJpvV
QMvSZScuGiBqbxP7EnFe8PPtsd2PgeiWN7GSNvtPUfNCUk4vDsDNa1cmlrsctRVI
8tRBglg0wL2itLUrwgEOOD4bwFBC01mTR3eBnHhpUovKmKTdhetg4g0YWGMyPbEc
ErvTfkeSu7hO+NUUdXD7rkyTRRsJcILy6SwwPDSzQ+E3et0KAiXF8VPqvYCcGFap
`protect END_PROTECTED
