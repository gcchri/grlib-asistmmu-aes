`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dczdt0BLCYr6C1NuBVWWZrd0Ohe3Ov0Lo7NZvlEhrdlp7uXneFOzJSWTPQaP2S7o
dPZPFeA9Zxzu4fz52YFBjjiGC6dPhsTamVemDnbCVF3HjHQEvAH1HE4oBSZZMlTJ
AYWk7yiUW2HX6pt/XEk0LbQ/w+t2fu+0s6giMzqUlmiIFS2Gi2zgfJgmJOPIOI68
5rO/0TCwgUak7ITBPlaJm10TDm7t9Pp0bf6x23y5+LsPCCAVS0nwG7/64SUi8qi7
JsvbizoWAEmmpKScgvby1hHZw/D7vF5QIJH9HSzjZrZ8jHcrqY/QeJj9o+4NKvvA
OK4NpOhXUY4PHMzy4/SDXGFEL6DvV3Ot/CFLtxgqyJ98FawnqeDJQWGl9Age4/v6
RFFhlwl1pYgtTYZLipOjBMvuEWsKUXIpu7DnZM8CE+n/HVJqR5JeG4RtzeywaYYp
jdaEIeu6CxhvS1ooaMEhAUXpK5LT8Fgsrw4i+BZvRi/a6zghDasY45+aY2LveIjU
MNsvqfqWSgwFWC9ViJ75Im2yzzGb9q8XwjuzFq0XKcopnFSVQU6CLwwGVu6MAxI0
73lYK0jPjT9UPFQkciOFN9Pk9wRexCKJl8fOgWlsuAJaYGIcu+7U65v73EciHdIP
xpESCTtkADLDCYPxFMPS1pKI3se+XSPpgbmtxSJrIwFhtE1FWnGPTp2x12jOE4Jb
1+1f9rIbi87kDvQv0BAaziQ8RjO2EKMfYEN9CIL0iQEMg/g/MKNDy0KMz68OMWqY
vWmY9kS7u7cnIUju/9syaYwB40f1sA1oRGnnACMroDBweafmy8j7DueqlyAEPxgx
mk/NN/i25tUB6FWYIQF5CPT0mADJKyrgPexiRe+2Vm904xj/ooLLh/Auqb7ScSpR
+D8wdnXX2F0Rcd9RY5XlEYh+n83ScTgJMvYsfYM9kx+gmxpzjez3U2DaKIjXvUQv
kA6AySuwyJRMOBj+XS94xCpJnaIoi++/InC/mFDNV38N9uhBpInSiESKLQDwlak6
lwSbjosyF2IAhkPhNxfgG8VHmFVoNAWiZMK+QToGE5qYeRlLMZRc/wpmGfwp+wJr
NRFa0oEyPiC4OrRh/nPu2+hyaRudiCd/NwHVxFYSKKKqqWvRv7HO1cQy/8/0IC6P
oYDHh2o3x31/elUaHhS+EJDLwGIcldSoaGC3ltYpD4tCrEbeVxq6wYupLCl05yMt
TWz+wiwN3ddpCS+2o+OPAz2ZyE5t57DApaa8/HYRKAzw59wS64dMRcFOFKx1SrCm
Qw4ox38fDuxGPH+hIU/1L6L9NhwEDj80kBk8grVJNCVYIZUCtzQbdrHpgjQ2C7FE
gDosuqtJDoftAWdTlRQetdEg1yuihLgyH6rpwyLr0cyxpbugkBULpVovwjcgEKsc
w/a8C9I/TaFkewPCgtp3aAmGpLZr7oWo73uyZ73+sXEq0gNfFviAWpY8Re8QxeIU
S5VouGbY6r2IEaDvsTB1eWyRymKwJSnH7dwaaTA7e4lLKzGla9O2rr+LdLU2vapz
`protect END_PROTECTED
