`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ouch8mz1Yo4cE5oH+qJK8UE+JIu68YbqsMhWFhTFVKpf68BCoYAhll9FPW4RMzNI
6W2etjIaySQQE3pRSPebjj1ZYO6liyWwt9Ei2Cm1R2iRqWv4rS04Mez9t3AuR6F+
s/eqxoh5UPiXfcHcE1VMylvwRDwfEU3RSgsLwwg8FT3mfLaez7ecZhZFYfVC9JM+
luCLcEmvcPzfBkUu56wReOMoL343oAWwQwsiC7xUI8q26VruFMx239IPRjAMXm2v
nZVUYIRC3a60lvnpHrnHwg==
`protect END_PROTECTED
