`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9p11bI6Fz5Daq8rQQWJPGoScuGn6xVZa/1TpLhz85M6yZVOVasvVsPbxAAh80bD
mtaKHIRNo5fpz07ZydFD1/+z3kcYg2g/APA+2sXzDynCptndnlywqRhvOrkQNzB3
g+IkaAE1cnG7H3Tow9Wigt8HLNBQIeP1bT9I3ppZVOcty4tzoifofJ8h/0vLTiQ/
QSB6YQrRtCBea+Off36euhI5q5WNZHMdR1A7sccTstY3PU+EtIR8pSByYpc8cT85
PcaU2H7AEVm4SV7GoeAqe5oN+vjcMJ1ZroM1Zxn301fjU+Evp7CvdinJRkv81mK4
nKY7NiCow4MeNTcm8FHSbVecZPKMF38C32NSwGDnuTS2JhR6m3jgq2DwsT9VTDeO
E9BAh7PuwKFtHI9y594DkCEgZCbKUaXqGj+tnobz6g/ShJeQlbXk+voiR0CMqItx
0iPSgFzXZQzOWRWhAcUiWzim75e68f40CUqVqomxSwX4eIwHXtTfgqXLFbclyQox
d82jM4VDlAW1Qk9TgqIu8GiERmuej5+wObzYmCWtXPRAjT/kLz7sYSZZzDBncHwg
IponmEvHjvCn09OHFcxNpXbq2QIMG2kiKbkPXWiRF0eJG0gUoN+foG4JAqXPR/Ws
dcoVz9vlzGhopNuQPVlmDQ==
`protect END_PROTECTED
