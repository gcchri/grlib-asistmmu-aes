`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhMJb6RuzkRQXdTr10Yp9taqNIu8c4D3fjFysGED7fdUbzcLoAovN8cFPNrsfiH6
uFqE554y85L6oo5P7Hp9ApF3cUarxC30ligDVIh6NjHvlD7xCnAF0fxljWH1byYF
opvATmkoeavwNnrwePKuTqcmmDI6JoeD3JCIxA5lPcGN4rO0DItbeGhlC8WFkE47
sJMFbTQHBM/dQIdGJ8LR7X7MIPxoWXXiDOqsUtI51L/1jVKcN3kpIlPxS33FzVYI
myIHBWgG6K/OeElYw5sORw==
`protect END_PROTECTED
