`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QLOr2GhBTm81PUaNt12UlmsHXc78pP55K7k5ISbFfPOq51tId71Xywjx2mSWbqL
Ou4uqpckR4doRD0S6sk1GfOR8x3qaLhSHP3360mRWC99AATc2dMYE3j8vevOcfJ4
fdpIspUtKY+JA9TQYt+2lsMT1AKEqql9EOjycgcBbHNFbTR+SoQQyw9n7xtv65h6
UtvGk8P91HJp2/gVjYi5I2ZvT0TJV2v8vqOMD+NOhEhkTtkznkiQfv+5e+mScFD9
LsoNY+Zp2TZH7WBNT1ZPazHzNCB5ONYdiRmD4zztEF1cwvZvOTyxF/enXuCZnKq8
IK4v/zFfJO+iHMmCS0d6YqW/j6GcY3sP5uIBi1LZMQExtRxklMA+hEFk6wrWwqAi
wOAye5ckBrtAPjOLMqnbDPj3vRCmkfv/goAS8oxOVIQk7tGag3StltQWuTZ6znrr
Kp9O4szLmdERDiYlPi7GnpjHFGkNJcKEqyfqUj6INhY=
`protect END_PROTECTED
