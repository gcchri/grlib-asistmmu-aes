`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B6rCtQAm0vnxp9Xu1jQIAZNRsDaY31s7dysMakjM+XIfA0vXbv4vDiFtOhbo5vFT
KXZm95Jj0x6M1JxAEZYCcKI9/CPlBUTcuUUUJHnA66biBxL3n1SmK28Aia1fVc/i
fu0bgi603xeXDpjz4/FNr9ihOwjAocizwr53OvUYAj06RqkcYLA1Ji8Eu8G8cfUg
No1Z7gXBeyEoSy4H7essRKbRMrGZ3VF6P1vg0i+c377FdKeLwYgYuS7HETxrca1k
6s/AGIVqAlhKtl0IpNiy4Q==
`protect END_PROTECTED
