`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KH5Znjsq59k1OAF95Va/PuBenpGjtzBRfqkq4cO43ncO22oni5azP1UbUM9LSc/U
LXtpuYkanej/jm8kBnd+H2o+vYemGHQw+P/79Aq9Mu7nkKpMDmyF5L5cTg5w1iba
lminDid19vrLUD0z/hbMEg04oSZtKG2dqF4Ai1s+B7vVnPz25C5pwGWywx89YMgK
KKJTkf5P1AmLYBNitSrogcyF5OjOSlu1iDXIonRvA7Qmbg09dyzUP6FYnjVcRkBK
sNOfBCgau0Jz0qrixiagyup/a8DOGe69GW4nKxSRW2CXkSoRTYa/lqj6kwS0KVqL
dH3hSsLwSo4LBaowhTLiPklRpRFQR9BaMiHLiHp512R0pN+YMpFF0sVJTMRppoKe
vfhcbXbmewPLbP8rD1lVkyduWclQU/AKo6m9OliPWtc=
`protect END_PROTECTED
