`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a2ZF3J+KUC4+lrSTxQiRlh9vJMkDD4xMLG0212qSdqQZ7o6tyVQXNQZaMdphuHvP
kbZkBZadcxi4MraXoJlOVQU6oXntt6jFTYg8RO4xw8h9R9ABaHgJAt1wzHlstEg+
BDl5lnVhGbMu4DRxajYzxJNFwqUyeI2RRjEVca5trbeIlsvlYpz5O9zFRYn84ZpO
3dSusup0UQSccpVorh1aHh38JbUI9L99YxQZImiV5uSeW4awqKuarQH3aRG9Cr+v
CY8oyjSMs3l43FvMjCv4G3Ic9dCPQqe1SMq2ab3AFH1KaJS3JS+TQUlg6yS3XEZN
PFiDlD6KLU4WP6zunjH5VfWxDBjQnWLGGL3kpLgH/lQykqKRMmIYcI63V5p4O79b
HJBE5EPGGSvNF0AmA537vOk29rXE4evYfJ5EbdbzSmA=
`protect END_PROTECTED
