`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Etl1Ps1vjep7eCcA1GTxETLXORILEPn1KbUQm112Ay7v8spzQVkDz0bLQM4GnKtu
xwm0h2bCrzSIxI/zSKqytLwud7FpNCCf0mHurOUqu5PQLqdKRSE1qQhM6YLLITGA
1toH818p8xmZ4/NYBjcnCQxSOvYqD7Fela+QyVz9+UXP3CyLgF/+gA+UPyEPdstL
YIT4ZdeNJUj/ehMVKLysTz4o5x55GgMvVTDSrRG2zngFeOy2xR/torjoBNi60IVY
7AgC3hZDv6aAKkdbPqoAFEPxGVL9rgz37+f5Mz48gto8rdP7cc8OfkKHiluqxIW8
cEDZ0OkKKhSrDantPRXj51le+ECM/Wtn+XBVJZImGgoVRFeOLHLCJRuh6Cb7K82Z
9TTd0kKQGL9wgd33hsM7nqyDpscoCtrZpP3RN0n/OlZDl4OEuKj/DTg7Qynof+AD
dbxizkVFuvnf3QuQBD1LLU5auy55sDqzh4PxJTbgNSlnNTl37Fo2vXIgycAwX6bO
7wbw3hK6mUjjcE1q4jjP5tnw3DqGk3At/NiiDlhU9zoADRKJkgnYazumy7UFA6np
MMKRWLRQnlzRHgX2k8mMgAvo9iKePG3SM+ZkYeoBQWu7YAHFwTFCr2IcdHnSJO7K
b0zB+F6holkJz0hvF/KMvDs3x3ciPAeIFpV0n0Qe0CLs5SH1vJ/z6fVX94MwD6DC
yzbsgZi5CVa6fqpn2f2Mq+ldTRVv0Cq3WDuMODp7tut6Io108r+NTpy2tdnlLXyy
rVFJh79svWMXXdSjwoHYhEHBeRkUYpYJb0uKvo03k22oU4vheaaV/dl0IsIAzM1s
ktYSenAHVh1N0PoVS6Wqrz0bisp8R71XT/NkhxXUkPUMH+svihIU68PX6PobE719
ccCHRraN+NGPJBleG5PPYzV9SnE1NrmlKGOhb7f6LQDH0AWqk3usMUzJncpN6bRu
IDnabVsml1b/GtVGPq0QvF3VnKWNK08FOsf93B+USwMwS6qOX6IOXtJ3BRMHqBLL
m/ofzt+bhVkuJepmUE8MYPxvUp+peOLd0PlPiFUx4nuZeaOj3ivKGy0SwEIZpt0m
ny94521kE8RJpET16hnbSfFf6bA0GuyGm4PO0GigineotIflF0yk130Q3Udbg13P
lY+eRibwjgBeHgMm3mljjYH4S80uYl4Xoi8IKUVoLjWLGsxWhOVbnNFnSAercLvm
h6/m9kltpXvW3VpBzq4VZofR1ZODOC/CI/CtNyDwrVUrZLVv+HiYlyHJkQlk3E9M
ec6lg4hshsUI7mhNXaLYV6XWJ2CsA4tSga/CkZbGh4P2ZH+fXTzD7KPYl283UJu0
aZTjcyeKhV38zBg33QlnhaJutnJ/sezBUZHZOGxdUUWXIzkmfeoaSzAeFeDRZxSp
dXjQXUnz0eaSpev1q6VuvhZQnyf/SnqoJM37mzGQTcPamyyWzBRTRWTpqHoHTAYj
eOCZSMBj+7zXflzMAV5gblIt6dDGnhoJNG3ZgAmZOeQ44Ib8ka1QXohUSkBdIkIj
/yH9tfich7Hx++MTQLagu+tNQCRExFoOrc8GWraEyOeRuh9vQyjF/ljazO9hsZzB
sfysHCPu0NKy/QZ6BkcgjF300fIpPFNR1qXQjcJVi4EFL4W8KWux/eyJJZmxqE3Z
+x+KqcVQ0n289G45zrOhnKpjH6bKNHX0qyeTPvbfEG2QxdcrsEaNfJzIRm9VShtN
DnKWYUiPXjS5jcxt7+Nxs0fA6upNgp620IoRAKoi+8ADaIEDbms+6Bxl0GicKsxP
AhDt9nhyIjLiVo613ODZdVg/NjvXjUnfgFHBFfG0ulGhn5NDJ2bz2UNG2V8b6wcJ
uZOOjci5Icf9E1CsUJifZegtlbJQ/JUFdb4MeUp6t9abvVLn5elOuAcS6fslQ+Ag
bSEdPZlVMLPx7kEjnJP/JxtvxcKb5iuR5E2jkSAQQppUQdXb5SLRHkLV1vqTQlRx
t+bWd4cx96PUf71elOu8fMhZl8V/Hnt/lm+7rnibu01VPX1wgAkF6oQeskE1WXwb
mDpESuBCO14aB5iopZV2NLRr4OUq2xbwmCnOdI0dbzvbOmP9IzHBUjHR8jXtPgK4
xpu3xEBTefrrKHORW7IoE+Z6gHetsEc4mHF3DHjGIrkYlXTZGVhrhBe0qXo/tD0D
rXndYAXEZETl/ZH5FQ0aP3gz+pviKRj5pXEnczq0otmqohrEfsZPNc0pGCWGwC3Y
sO7kPDQ4ejwWdya8BAIHmWgHwpr6///JKGhWeZZ9Xt3H36ARkm4lAnA+eiKdsvmU
UJLRXcWUNm4+I5W6zxODqMEDOZbe2I9uIkFSNc8jQYKB3G95PvPkURLrH2rUPOVp
H8TPJGyCK9IThgrFvRlSvYvzLPuOWMwiE3DvnNaWX/1zWbNp632azC6M5dEcXavo
cxKbc2ptSWD4RoIA1bUdU9v51zdUFdKdKiJZq1YrIyPP8kP16V4vtIXoZYUpdBtF
3MzqszJ/47UPz4P90R2GCzyFYmiNoD+m/Nx1TMJBEMQHML23hTfRPqr/pV9XOGXt
`protect END_PROTECTED
