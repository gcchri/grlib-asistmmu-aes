`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9WA9uLpYaCwaTaqVQZVbKT6QKROkEq5ReajcevYN28XgaMvBVdEGSn5yAkMHSC1
kugT7fHHddNEeZZz3QezH02M36qceaMRCblzYqNptf7QbGiV+kskM77K4iA43tgB
LFMvtikMPWYG7wN0LcweJDaJCI7Hm/9H290e3mNcZ24Q3x4r0HLtId8XzbEvIjal
NiOSyT9LmBqUx1rErhUb06LTEpURWnuSe6NBERbsZowB9rQRUdSLWOSJ775Hxfmb
8Bbz3nTqYxtDJcrenADMsX/9DxSQQf5u2/G1uvqNVr4yCPtLoaxuFGGHK2DF9ggE
4+ywbDE/2+Gla67SbNmNzdaanoLsixuIfv17Jw3cRBNMO1Gq/zm5liGQgMCy8SgR
K2Iro+2xsR5OHOhh21ijfpM17GspVM4rDzN5EuIxUh4=
`protect END_PROTECTED
