`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUE+f0Rnb9IirModgSL/TCj8TKPYCZ15k4jxBE85CZ6o98JR9KnKiLykuMGyBnp8
JGDANnYz4QbuWHLYW5EsC0W7z5D6t72BCfnxU+/d4TrYVzHS7c46UdAWWPLjQ9aV
lvgNPFz0qW8kdx+Qp9Eso6NJCyn1b1iKVQFZ5oL7TW9lLCZw9P5f82nryHTzZcxb
QLYLvtnyISM6Fuj676Zf+07+Tj2ketqPCTlehReE5S+l+FvgyiroQPTZzRoVWcEa
adTPrkQNG23gt7CeoLLt9+cmt8TmD2kjS3jQg/hh/L/6bKu8fLmy+s82oj+j7snX
/B952K7V5yxtExLtKeyEwIimReEx0hB7KD/NpIbUFJ0MGrNeOqQX6Djkm7z6kfUJ
Z92cl/eW/HA9o67Mcgr9wA==
`protect END_PROTECTED
