`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Nb9b04I5DNMJWIc0jsMiGXUeddDlV30gu+CM0RgbvffvIKPkhPN8ghQR0NmupJ8
XgI913kt9d1w8I9ra1akj7FzCGLLq6RvbloYAw2HT+GTFoOixsY9Lq7GNh6IBXIN
gGdXkyuKVU26RXexFFsTrq47y4RmkKD0OSPweSaUVclu+d4fivGzCvXakeIjSanq
CU5RHPJSb/jTWZqkGTVANnTLHuU4qwaTwc38ipTMxNrVWNy/NZ0FhRRU+6ll8CBV
kqInGLmbw9ukE8BmU5bcQuR4zdz7xQkrKw7W+HjNHOLcPpPIn01s/xUXhvCcHGA2
a11IsFcYbDi6PXYC6pSqvCVFEFznpQN1qfwgX6wIEwwJdPQbxGAF6jFOkt5pVLLT
wCyFbnMAS6ipHgc20fQv0uEbkUMTUAU5QL65M6zM3lBEteM3WckugH7ePnpQbjr4
5zPtqKKxa+WgjSLeUjrvAl5uUE5cld8eE3vsllixXMuWbUxhL0pA5Fqe5YROtNTl
8beW1KopQpNdXvg9Ww4OwqgNEQRbkRqQ94i8Nk6e3FsxLlr/mM0TawBiGEmTeW44
0KmD8gv9uZpToka0UALoO8eJJr5OguXPofxnAXiy3T471xTnIO17eHVMYubC/Ody
UP5A2kLQHCrnUhsBPOZEBdKCpajigp3dgyGLZHzoDxkJBOhF6Xk/R631hxeLcLH7
ehKvgX6dtH9sKw9c4jVF6W0oN1WR0HYhVHWJYXL5tehGSi5lATt+55+0gPgJ4hi3
HF3kI2yti8iD5hy5QWG21C5bawiYTxN+Go//dHVjtz4i8bxVlmq8aoapEm9F2QfL
8N5rEfNbuodJ4jk3FYjTDazrUnqER88c+tJC7vog3Hmts08oQFeEID1XIJRIPElu
+/Dj2s+xWTniQ3VEGMK236bkv9+0sSm3RyvjeO9UYxc3AwXTT2KM16mcbB8xE0g4
h20z5CqX0iyzM+bPHym2jTO7FMmFefIUzEHY2dMkesCmC+DhzQZMftjkqJOF+ElK
uIZHcNJDxTT0OKimryYwdJDYOeXd0FuSZL/DGG9NGsZXgIpXh8YkeT21O7IEnQeF
0QA2RS/ZmtEUAK8ith/Uplb6HShfx7+M3zKUoM2oryZAeeYlcBHRIZHi/nq3h8rD
+PLzUSe5qzB3X+FpfzHtGlCnhACikXyGSnYwG4+3ECTG8/0sE9UeNtaBMGSRJp5I
xGLD9Ru2x49XwgshBeBwqvf4mcR3d94TJqEjC4wid2epePZJ5L/5pAfibgHUQSFu
wXWmvbHByc9bF4jiSfLuKEloee9CULkjnsrTcAYUe/joaNA1RL1xqY7GOTk8cf2L
UQtMR5ocfZiJ6vbdnmicKOOMJg/qrWHqZ1RknmaCCoK5IQxDVJ4g8rFTD7QamZyc
kVNawfVEzcJuy0sjmrvDH/hr3xwBGPmEtGNZqWiRcKhbEL4saF1JGrE+dzB9vkPK
cu2KpDnt1BM6rUfS11MOclMAHWu9+Bjucx3CkyovGAA8t9fnHHc/0U2mT4liZe98
F8UngxlXvTsLYQUjXrj6ol16GtQFcx/P46aLdntff29C3ew1Zu7J2UBbB/pzMegN
exs6OsazH/m3fmWMCbBWgBHGWoOqyr2t4Ccv14HKIDL7kRO6MPrR1J52Hnzredaa
A3NXVVatW/qGlSMikQFvCA==
`protect END_PROTECTED
