`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pR61pQOry/zLgf8Mu6WbLY1yzuvidLdiDZU/LQcWvEau3tSqH/CKMnkg6cCOeHw6
sNGjZyQD1BB9dHWvluLqHVwelqq6hU3qtgvilhlBYRZ27VYyEME8GqmJU3st0p3G
MgsVcYFoqBvOdT6uSH3fmC91kBcAUNE1//M6n0FgKV9hunNxIrF7uNsrOVhcMGuJ
NdVXj4sRIIdFEuB05m29s22QGOqNexvLs3SYZS5D5gC0VvHQB95mptM3qAm79ft6
JQ5eIcoUIdROxMPMU+K4H4mJcJLat+2jSB4rYyZo7u0CP7FuHF2KVVSug2heNVDv
7fVJSqXpKyTfzMOD8pkfCdrCuG7LCV10iE/pC8qt7dyp7gp+n4gXAin2Fd1PTmxr
9E6YP/BZTHtPgLOZKZnDNRFZg5L8FyCqWVkZHns5k/Ftv9iqAoyjvqqT/4N61GRf
cPeVO3wMo4oMpywLQxcYAPrnhrkJvqeysVQ2NqOxVrDl4EMRDyRSpClDSqCs+eCQ
rkFYVVTWjDCsw/xEDuM6hGbi5jrPgCoUv5goTXo18YEvQvbzCnVW6Nxij1uxaXDN
MNsx4+xsmGinYF6qngyrldfWIO+ks2yox+4aA6STdUdY6LQ2XxNfoamvq5p318yS
HK96ODLap67XhXEXvhFgOkhJpjTvu4wmbbm/Pp6ogfRUCVPAcrNLLZanRGOEjeEO
b/4x1Pyojl5b5plwUc1hE7CYPzxu9F2fUoxMeuUHpN6Wr5srDpuuJuRAS88aXywO
AVN5eSnhs9//DKHZNxAGWehm7bKx6GKB4U3RNnnR6bTqoZFnEO1KzCoIAJvRiPnj
Y7E3HtyCBHr86B+0MtrzHs/Uwe9cF1bbkmKSzDdRki34i8i9sj6Gj/roArbH/4A6
6eeA7NwdhEmfYu+QNKPJROVK1ksVxRsAh6QpFW3AzzkSS6vQcgFAGbMxr6OrJgrq
tJmZSTJPfZ/+qlQwHkbhEahOKq4wD7uaz1m8khWsI3x2RgH2tnzRLpAWQHteDruC
kqc1hu3rPNpGMCnzVfQxre3ViJnrAbpH7nfcOxwwzP1p391dsP+tYg5N42kpEKSL
RCucrTVjfCdDD2Gz+CMi/k2+8vnjqmgEUuSwJ+CsVSCF0jP2GMoPdt8FrTuGaDdK
u0cjUaQJYc6ylTD6lMio+mJNLXJhJBxjbruoVGRC79y1lmlWM62QihDamXnl3odX
ZFLgnDkA4Gd2zrH8Wg/94bxFSxQM0yP1JEYCZ/3lk/d2AWjdSKSR6FnJYIayllJO
2LtMgBwSs1Pe62RMzutvHVQwipUw8cEodDx7yFLDcH5Kbmw/XeRmSCJXZe2KPkHf
56QItifOay1FkHJu6hwfdYH7ZEPGYFKwTSBvbGROGDwlVYX2wXxD1PLZ/xPLZYQf
GW+phoiBp+v68RPpuvSjDXn4p2xgbRiezL4f0aU4Mv1wcraSBi2oNp2+f3Rjq1Aj
ajiQoRt+igW34lkib0yhBfadvAPVW6ArGF6f7cL8K6nKrMq0Pa6bc/BxImg1Vv+q
7IJz4xNbCa/Xw7ReNCdYGB5o475f23p29rQ4DG11ZdFs0+0PMOKBeO9x92ddK0hl
odAiiFJQ8hLlDNOI8tX/CKhu8XAsVwcSdqCsvqkSFwch7K6FllYN2S6IeJcj5m3J
BBNYCr2hiZKpdYagcplr5JzGGyGhuWBSgYdkzbCtYmitf14aY/u+Pf3CUqvB0el0
9BNS/3qDtGpJXtTjgeTla9XbdlKkMlnruEOYX2TVHBsqhazfM2wmwc+E3J3GkNS1
RyWZKKBQ9b56jIuB8DK+Qm4MQ1YMfcos3xEWTOySJPNZonuVnd/qpUAjhP6gnsbX
tcsc2SxDKhf2nwtGBl/3aOdLELytldAco9Vgy6BD4KqL59czy/2b7W7WjLjsjkRN
2GV7HeKnz2oMOS0iMFBzMzQS4TC92UQ+j2nKVI8ft10hTQHnMJCU3z1Vdvjm4aOw
+OevqItmig7hlU209p1i4zgNZSp2PjHnuC3tkZIsdn39YckuJHsPYQKLghaFh6JW
efEKOOcmmO6eMEk0IDG/N7HIWiF98/49vluV9fcSFYPSN8byGgQqhjNEza6MDB6f
naVvyLhP/F1cxUnVDdtJsA==
`protect END_PROTECTED
