`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wWRFwsMERzCLF9xnm0DMMIdh2VZPPb0JYEtXJJapBJHy/DwX50RsLTpZafsPyb4k
Nsl6cAE90N6pjPSGUrmuJhz9pvi0LYs8Js+8IUcqIn2XeyDlFH6VgSl+KjOo+NZ+
fv/DCcAMNGoJ6can39NDg09Sgcak/1L+hn1ZIACQ1SJN1m2CZbaYzAj/AtcjKzZG
zS9xlJ5kvciED3enrPZgQvEoTaZz6sedimMUNym5iZQtGaycvs3JSVnFtUIkL0Ig
TB/1TuRKY/w5GZbv0NnoDHbC94dDilXJV94Zo5sKh1uQ/+mHe3H+dZOXAkQzuPFS
dnerDycQH4xLFKUflYz2AA==
`protect END_PROTECTED
