`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n58YwWuwgi8I2HavAaO5oTtF67ypCSZrO2M5IOZZjCAU2tGtUKM3HxuLKEogafEa
DGjS2Mjtmq0ElewvBF00tvfgpLE9dWwyQek9+RlKyeODOEgxElWwjX9wFeJdVFk2
qBVCyF++8cvWmClKKegFiXBcM9+rC/yskXcL5+Y+P3JQva8E/iU/+9s1y7+gOu5L
IRUGO3aS1s0g91MIq3XD+4AvqORsyr5OKbQQCuc1y3uoP2vuFXq3wEarLUVZtRAe
95NwCzcU4t8jCKdkmtKOQ8TwOPqgZztUO71PrN6o9tv/qkkCn4JFL0TgCzPz6BXV
y6XI0LNmH6RS08tFIFbYZhk43RXCmUL+ubsJrZUWnzQ2lxqtC4uZKYFvR+qM0hfF
2imIuIvS4ioNig7bpXgVwMvqWR0LBTe6qcKPyJ/XniAHk6my9RwG1UMcB8TYx/Zp
EAI52ldwFOIlys4Lpm69xJ4WTF5HvRQUNKI0umKDJ2NPM18mUNTu7T1mzPcs1WqQ
SBzb2Gdmq/kSYBwMY76YULvNRdlpAZyDN5rVAyT7Itx/kEnm+lZVr/9lY0kFbY4G
O8T7Zs7WzXjVjbbZ3nFWn0R7A17cDXgK55/98VUT2Xw=
`protect END_PROTECTED
