`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZTUA01pI9a+NwsmtWNrE89pD9gpC6d+cEVVZc3KgJ34nHqrXW1pAQBgEMNDe0Rn
8XHcyALYR92s7mdFaRMN3Qgl+n4t/MTrEW3PHoddADnaa8SwT/RWWNFgbxQPL0w1
xCyiq7Y2XPuqnwBwWA8tl6IhiTUL1eCLn8tMUboZXoeQik3PyztXz4Cx7hcXXBRJ
/OU/thM23mopE9BFRcKh5S2Fs4Cva4ctmRVyyb0BIjh75tymRYUIz5obZQzGH+9i
06hzNpkQmPBVe9lmYvot+oMWuNp3FfQaGDGzHCV4KU0iXkwf2aJYsxNV2yoJVGFH
w4DFExgGp7U/YMhG9PD/5bmrR8biQhf4tvn4jfmZs+ouQ9J1uidt5hO2lGVtCJuK
tEsENCBdEWSGqR3v06TS6I28AvQk1ie/yvBjUKXN2bGtBBsxWIZcHtSd9O3hs/wj
PZQ8q89VzXSNu87SH545TmS10MfLdeQMolXoDfIUm8rT+ciIJXrTmcVsM1W3wVm+
ZlqatGdS2YoNUTMRLhoEXCZw/SMRqJhJrrsRaYvgHchLe3d9cGOzdz618+XBNSLu
rtyXfkocfiX02liVVdSEFBFztw5NYi8P6bosta7wFt9HJBFIhlHLCpi/4FDzTEzV
KUpdIR9dgyWRz+ZB4Rk2991A4UIS90yBZEQ2BuW0TQWZCR3+oNFW3GanjMmn/6xP
dj3C6L+JOgDjZl0Ml4sApxPhQVxuZbdF7Bi9/keEaE/c2SgY1fIB0rwR3cNdtLAO
w623xpGVxW3jl2Ta/DsHFk3DedsWzL/OC+sfqSmD/GDSZuaSu6/J+i2brcVl0JK+
ZTKwsnavBH3mnFRGtEEac9kKKtdI0UeMEbM/p4fF61ot8b2CvWdYYX7QyRX05dDF
eanl4CctEvOrbE+yJMH6DDNm9zUvYR8uStzPtgBTpExDMvbKHCKKiiZ2en7RrAv8
zbdzzPhnwy/md0LsVFMEzVEtVZifOrwSm+BbrvBfa23KV9VA3XY96IcJHAmGUEI0
LeDKY/C1utb/dx49A1UsKkmRBcWnnrLFK7RlqVi2pkrLoyL7tdUrX9wKDNp8z3DZ
K2fb4f45gXHCGrFLzFSszHR3ulvGJb1xiLr9+R+KmJO/oWwCBmiTRB++8KB6Te7q
3BPZ5+1a9BOeJZWl9qxu/wK1aFRD4BLUhu93pn+A7uYtzHHf/M3bsZsjcvykqhSD
P+TRAceWuAXcQFc4zeIyD/sHw3Cjddp5E720NUt9GSLKLSjV3fXAFUOhazWemUkx
ct4oR1wYdrn0Uo1QMA1NPC3ctQcGBo63ybxTYsyr1vFnzg6QB/fEQApu2H8fWtTK
k9whzDp6JinqDt/nL5+fDwcfcSZ4TWIT2EYGkL9wOsXcNa8jRYSrBtn74F58fGxH
RnH586yKZOvNRWbgF0e/yCj52GNClJ2D6fnFwL8mER2kzBhwL7lC2lTTql/N+45o
rNsI8OJ0mr/7kPLwsCgrTgfNRVDqdawGtguMPQTnpNg4ZmGg593w7IocFvkCBRLC
JjwXz3zFYlyyczm/bwXL+IGQ+hShe0l5zXCyxHNGLYcaMz8643ESXh/uD9ANSfdT
Fh0IvD9s6wPnp670Z5k/DoCNBKAiPZdYYePIMXndQyV8oWdh5GTpxlyONCrolUbK
VMkaHy1j/Y8EZ4MxjWDLtU7YGGeRhXI9UucgGCeLvuUcM7BGVzUu+kaGBxJ2/Zu6
iMMi4b6fa63m46jKSbuBw+3svPd8zKR3fQKjbJLe93H/x+SKjdAsaBUxT6LfsdXC
0091RZJUjTrri9RksD3S8w/skgYUNA4d9c7jDIIos2DSc5BuXeGQCI6qTwYZEjGJ
Fjyk2lKVdVy1GbeZRhjUpsPUvrmD9t3am1BOwX0zrYs6s4nWxnkY/yLzmVrfUujj
wKEYpARDeSv9vhzXigNvGVIH8fYlgZFXyzQy2W6p6of8eeLCz9fPRuy9UAr6LVth
vNjLesMNrAKromr1wgVv3Sr7feUh6pQJiazj0NSt1eHZExY8fVyXccaRLkLHfZ/7
GzeIVyD9/qi12OYArSHCotORGQMVesq6PZVHbhmOoyebyUPj0Gd9Hzo5lBTu9xFg
LJ964e5bUDEERAtkTfwRFAvJdeR32/qtVrM5Cw6XrqtBebhCDpsiSp+mcTFgqrwj
SUjlpyKj31D+4KrsiANm3hkDvaEtd9RoU9bVpulUX68AvpMSy1jRkQyx1INgxiWu
Ry891OXAxcSGthHLLiUdmw==
`protect END_PROTECTED
