`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TEGACFA+2l8zAYZKIMh5Q5BT8vofHUKnWal7bqz6DdyPrK25W1xqrE6Tf6SN3l1E
9WfVwQGZdq+dPi/oMrEO7V0r8AC/c5Sn65+Y+HUL4SEWOM73VUw9bUQQhQawkkQa
xZgzZ/TW6Gh3Dtnb5dVv1pgt9SSUwYO1TQySzv2tNijtBMZNoI3nFFTWpjaul5o1
gLIRWiJjipfPnJSsRM0niVAkcYxSNmRZzGIDTBnh+s5P7oKP9nIf1EQkvvkUj4+F
Pd/zxGYo31nt/LAWG40FEPG2l/f+J49ax8GCYig6v9fPvejNTdkj4aUlxNU38ZK0
fmw+ooPFH1x1rpd/C8Qwma2ulVSB3JA7ahvjmh2En8vuj2aRKL7c2ixnOJu4jiRa
SU25b+8FjQijzUqwSrLnqWeI7S7nj7JsYPUs0Q5VzdpfiiQLNttcq8Y5ZD0dqnK8
WOslZ0hs6Dmz8VAZZiHLNA8tX1Nt2VW+1XATnd5v6J8LKOpE7xtqEAA0sqmY3EGW
WZRRB7VkHbiNeKwXig+dqTVeDdhEN8h+YGQgKAs5ubHsos4G2TV9fa9rinVVjb43
YzfkmJJDk1JkQzWt+SsxXpYX4fzOURiZBDkF6QpILWbvoPC62Q9wefpBzqYf05V7
bpviBGtqrTm/R86x07Dh5q+puIPXzEfX8o0NWkDAdH4AhFyzD075hX4TvxaBXTb+
6TD8Wd5DBNl07RHfXHinKM5tiTktlfCxddFzR8kwg7NXc5bLLEvsRHKvPIEQ2+k7
AR1FUJ7U9VaTaL7Me/UwYsmW6JYVI0jEnsfx/ckbb0NtBJHJRc/Gg2+xOIP0bhV3
94pkKPiQ3n/AB4JMT9n+VU0VBfV/73+pKKj+Ps+0dSvsDPRqPkkdci1Lwwn7PAe+
4B21wryulzhIzgW6s6LGNg==
`protect END_PROTECTED
