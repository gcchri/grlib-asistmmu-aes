`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7rmz4vioR2o12rJmwfkFHL358SWslot2K1FHj24gMyDQzSiAQaEM0Yp2VGWUSpjy
Xu5O/BCP8m68sjasW9FNMyd2q9vltp1iEfwePDwSR11XQ7bSKAx4JUxwP0tCg2/d
h3eGaoTBr13HDS+2Sshtljwft7jUFi+Vdj2s+aUDHU4BGi2L3XN1DvgYFbYCjkyH
1BZY9e8/ClPPEdmo8UhLxp3PATohSij6bu3XVDB6MRhjpX/gf71rsEVMX6VNh+m6
/WklkAxtnyxOkgjz0LRUDk9KhM08Ns8q9hkeidpMGfVAg86SDoh9iVi+pcsMGOer
yehsgc/dnJpB6Dzu8j9qnZ0hFShRhECF6jbg04ZJGUkyZfDgM9PCmur9uklB3PE4
r6triTZ8/q0PLAyVg5X6aYoziohrXMjG9JuY/z3j751y9WRV5Aicq4CSTc1gbeAF
Q5waU+LnjoV3+WtXKPwbZOQ+4KsBqTan0t6hMS9X/jqCZ3NLxTSgKfWzXg+PgfPu
`protect END_PROTECTED
