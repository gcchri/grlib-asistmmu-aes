`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YEvphlz8BKmDqB7xqQs23updFEq1sxmGr46Bzsdn61+PLiBNgfbTp8PDUVYHuZZu
V0FGOtDdTHi8kWOVG1Kfq+SldwOEnSSb6pQsltskoGUhbbPU/RkEmCRtZdfV1w7m
Fm5GNVnVxu/jKhlDn/1jx5GvcaL97rnz9zxA1vkFMLx512YIXZpZ9YjHSMUdhkKB
ykSXfqMpGZOybHUPnUaPME8Qb2FB94hCUVBQ0mCAyKY5f5Y7u0HLzT4huA+MizOL
/0AQkcWr55HdFkYa12bUVPM4JOlI/SvAxUksFKZqEUD4tMawrsk+Z+w63JBeVx8p
Mj0IWpvj1cEr3mG3UwTtQkGJS7nRyUnTqimipBDk4OEfh8BxKouBBgsH8PFNQAQv
6KEWI4JWrZGSaJsvQjMzyNE/9TTiWAKNfTRCbHlba0ctXL+vzPhb0hP2CLQwJncj
k/HVkK1EnElsWPMcfzC0K7Y5qjUX62ZJeyXCrys1NqoEYaf/iU8C9p+rUwSyOt+X
Z3NXddTA8hgKg3llUDqwO59pAfv7pHeq3+YcJgffkGRzKC1+dtaSYPmI5gtq2dYG
o3vYBARdHkoG4pGq0x2rcWkoXr3TacqWxH/9JHzY8QH7thH5k1uMXKNB8TpS2K3L
FExCiwKYfXUgmk4kN3lCgjezvacE/gU5yVTiloEo2GvrjlTBB4sERhQNbtfxjEMR
nSczfORN+UDyZerz6vR2HNmji9u4SyFu6bjXB04BQbtq5rPgRD/jSOri4IWM4rA5
sK39fpoLj3fa7J+SVcOBtfwosZ7wZnhvJ5Lb0WUXTzD0TkVkVPDT/AW3pz9Ixusp
CYOHLUMRcXzAosh8EMDXnA+FSVA1KbdaYPVVJGmSw2s7VxYFg7qfqSl3rzVtl8uB
O+iDyxdXquCpjZX4EGSp8sYov3kV7LZj7B3vQgh1xnU4Mio07i2sbVoIokaqFg6l
6xn2538j4nMWV1cxd7IB43HicaJN1RBRPsgF0CTAGAL+LNUjaA09NVkdM3Yq2Xh2
IOAj2LjVQ4G49mpPr7uLVy63y5eNg4YlRuEDe2hjgyH34MIyz7fz1Hc9O6qjz3iW
1uYuVU/boOV/FpMcXtJev19CA0LUFa/ZQTB7qh/mMP9O/zA9aYSKZtwohzFPCa3d
`protect END_PROTECTED
