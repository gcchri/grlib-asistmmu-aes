`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCdVT942EL21X5hLlqQt/7nI68s9GgwQtwyVIyqnU9zt/J7rpQqnfb2ByAOXtANM
hVb3leemYUPNOWNlNIaZePEh66e13QFZNDd4luSL/8cYt9YQppgfyVEkhE5VrHgr
fcYS4+4XQnAFtzQ0Qer16NGsRy+mayGcL06NyYfONGEiUgHAKg9n5JjZNOuWh/07
nw9ufsQFZjciHahul2ec/c2N0N1Dp8qHykV21ibrr52T1Zmj6sAMpOSe6wsDGavX
alovpb+aMKeC4YaZuxSsQ4AmWYEigg17VayaNmrGk39IEv+vwx9c2U7pMIQUF+pu
ErvtImGCr0PijeNZl9kAdm6N/XGALbdDSwzqHj3yCKeEWHEI+2CDBinbT3l8XT27
sKlkC2i6XrzbgLJwaH2DkRWJrhCgBfzRadlJaHyjpBaYTy8/RZfmMlktvW5V7kvB
/hAUsPOVkBZRUBUJxysxYVfDYK/Ou9iDyC7Wy7MfHGAvnlg2y7ur1/pFGaw/nG7U
aRFnE0o/5OI/bKZudQeLlOLSiDhXg/XvGRwoaSAzzE+ziaG8KrDdLtWwgjs0z7xt
CGE0Bt6rxEQAutRQVbylHg8uyP0XGIt2SK2n066H1JKZWFXQSls9gNwIrEgIvazq
Zw7qGTiogKItgVSVLo5koVCsSRaMt9dy3JVfIPMfTQ1WeT7w+pEu1rKsJd9UaZF0
Ee46aArL995g3sj7y9D5RFcyQt5KU9X/PH40A4Bton/P5hD+DnxodZKm4eh4YNYm
iENhecX2QihFZ6mT507NitfWDeZp3/ZVG3fx9tHHJyOQ6CEazoBKNDRNi+hwVNER
7qJEIEeMGQkvs8qybC8NXKw89k8VQnzmCxWbYlcmspY7rImCG1NkiRU0MwUmoiL0
WiAjIUnz1+VOdvdcEqXnyy4Z4scgzOu8TCxPof884K6hSm5x5ZVWWyzo1W4q+c87
d832DLRg6k08gmOw0cwg7/xLJuWvaoAGcBdwnBdDXj1G3AsjtQ/L4prPXk4OYdes
`protect END_PROTECTED
