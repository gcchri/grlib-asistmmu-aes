`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGU/eYTmfQjpiFFrE/rvw1rxPyXvOo81bGUoVTn7XnTgn6Vf2indnYL4fap0MShT
47WlUksnhUYZS5WV8u6J+KpeZFUOA8TrYb0bFtr63BPZu7Fww6bDiCSh6B7shTm3
oAi/Mca4Tr2/Bxachlstmu009OFD38rmsW4yGiL4QaQgawddtBmhH8dZ1dAd5AYK
ybcQTOWu2zioyPQRMPJWJBT8NEoTSa+xDhN0DlfWKwOinf1rEVS7TRmG2tn5oGT4
TWuW4IarP6WSCZrpZl5wIIieuV5xyiQQZhH5FQ7+PSOds+vcEDxV6AX0MUFI3awn
A7wfZg+TEEf3AadhMlLeEoXZkJqziagvmHWeQrrDVUObs1kfhuoMIFToFn0iOAw5
wSLMjw7QHEhVFJH6tYtCf7UWfQwKe5xcj+3PIfw4sBcGSsnpv8G9epCVtEfj17Yn
u+zpMJE29rydFgjvXqXX4qCgXXwuvXwJm8Yb1aFBBEsoSmhLFQ8NmlCKfEFsLwNC
+K2Iy48tSRIrG4NIQdmo6xSJ3DTNuIv+z/8Jy42mttFXCf7RIDkcPBD9x5UFlwLp
ZCFFTWZ6Ewof1sU0BU65RPlLer/udK9dTU5txpXhvcWAfX9iRtAg87lBLMM733B2
gyGQhulf6IOUu3iGfjCjVupMQgbS/3EnBq4pM31fvasxNbxlqurdAhdPR6+kPcFy
iNBRS9b5Yc6B7LM9DLTUqSKgIkjgIBfhA5qRMseqemfiMeWzDK9uSOrijLuqmIQl
ylFZhw1ERCVeOEl5ayBaiLCG/u+3MoRXFiH1yxhc0duK7YqA1iVKLYzEKF+ZVos7
OTf0IqSyqbA7q6X5coxWxzQ0+2q18dBd3cYi2v1ZVTe6clwIzRmQm5t8A6CoISSS
cDup/9u1eH4uDOaDWDWOBivkjDqknstXi/UkMHc8ou4nTQjk0G3qlcbVKnK/voN9
FTviyEPwVLqR4jZxR7SvOTjRiy5kQHGHClKs0YpxYbw=
`protect END_PROTECTED
