`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfSDIlw7HKxvqVBt3a7mp2SsCT/3a5OOVPXVJp6AL4d2mMaJcOmbBIwjt3FutNjX
BiOdSRqjyDwQfb5Vw/678BqMdakG7ZSg4MY+SmWbfcIosYiaaIbfrcx2QG7rTFIb
8VUz6jPP2bisedW6ShlCFj/UWlxIV8OyP+Pd0CFppn43ngJ6uTgzwt8WSoGuwi9U
/obzQ8mRTb2ZMcCWn4t5BlXf0zSyD2AzrPJW29Nq5KPfiUYrcoKct/NgeTgT0zMr
ideVGHRFWUEL2RQeI/qJw45ZtDehP/Rk/x18I7DQaYEcnsfgzZEdtJ8iuV2dz/Wf
3ex2xHe0lq1xYSETmkURbVb5TMR1sFuOkE465qGn0Do86S36o8mSdBaRf3t1fHVw
mAkyt4SjgOHAMgqOxiWZNU6+NueEygKE9SKxNfCpmJo=
`protect END_PROTECTED
