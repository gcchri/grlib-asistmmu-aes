`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pM1aQENApAohUwOkq0X+e2ATyqgEEU/V4BVPK++Pl1BZ8MSlNzg0036v+SBNcSmN
/82Jq/CHliIoDV2LzKxu+V5ghMKM4L0kG774zjHcT8m2zr5EEzzT7Uy+3lb3VQeu
7aMUhl8Mpic/NZy+upjEjZslpWSnHbLLdcSJN8j66VG6QUD7pJXRtUVJ7oIqqF4l
qo3hANSfY1u/Zr1hQVDci9ce/GsZ5/wPmBiAbpuo51AYhRR35Nuc63pKvRgRWT0o
yhHnNCk03Fp0hdP+icmPaO+6syYMUFWDjj4qXl/FeQ5ze84L5tpQ1S3vWoXnKMHQ
dfBwrwC+slQ/5CTS4TFuO0inpPVapOQgsqxciBW/VUnbzQ7O9quyLjmdkYDTQ3G8
wemA2CQ42FShYYb5zU0lcUV1t6S2fj1GJbbM6wPyHeH3+Dttb1SVTLTLA21F0Khl
XlfQjwG28ApH+npew8wN2HIR9xsNVfp9jApVCGcdWkH4O+sAIb/XZq8vHpdlMHn5
2G1oOMzrmZoQeOi58ersHZHFhy7sOTyuxngEJnWyXG2lBZDSlxuTdtm7Ypp5sS9c
J9NY4Wlc92GLZW/SD2kn7jC9xS91qwQ/HTjNiHcYWjuwrpN7IeQVLwbCIZJDZSQk
zal+6fnuZIuj2Qb/nzk1h//BG8nFEKgQkeSl1PLi709Ul//zqh/3CNHX3ek8jwwM
AjlsSmjGQmkTegYz48Zzk250E9Kfy1Fai7K7PXaZ2fA=
`protect END_PROTECTED
