`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BcypR0HSqWUyfLNs9p3rxfKg+VchMsp0Njq//5BmxHdzq7tFqmAJjPEnZMHJZHEE
vXRsn67rQMlPHuabgUFM1G+/C8L9GHjKbGUIqH5QZuRzGsXBRwW3vUALSaN6pVaw
X2fpPBJn8FVGBTGaiv36wKnqeMl/HpJ5G2lqDE0ABP40Wn73sB1mqJhbVeDus788
I++S+bhU651p6zEIFcXHdwlSBSalTXzWr35EjDJmgQ7FxkKyJbH9sRjj+RL5Vgxt
LtekMUw1E5w/JgysOEq+0QatDSlzUwrbFP9u+/Z+cvFCB3eSCYX8tiIKQj9WWzYh
46Yc7xWgwAn9pRedC0tGFV76ceZpdp6MYpHAhx22ebpdUp6SwAwPRB75I7gGjnQP
EIRlswdbmM/FA5hIGQntx6X6axHlW9wEiaE55O1KrpydkMsKBdKG+Y/GIq1HA8fH
wKNByoFyAlQQ3S/cGJ2koLhR/RIu0XYCAAewYBcF3pW5H1DH7OUpj5HhTYTq+VVw
Y/r05n6X+MF4VyqGKkAsfe8Zn8z4HfdU1m5CjMjDEQs3T+WWPeGh+gzOEQ9X5OHa
+NeCR1L7nkupEP5lDPRba2yo1xxCEPAFKcGNYQX4w7gFXw3UHLx/ZHeSc7cYfOek
0zCyb7gcdAEMOV6JzAkKp0nKw9E8duSYfegBwyU/RBjwP0lG//sIVoG2k/x79NUp
2u+bT1fMj3ftl9mMPxt3nA==
`protect END_PROTECTED
