`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gxwl9+5jfn9sNV2RPjNlcyCs0YcVOv64TyaEnn16+wEbHFPnImdfcE0aT0FC5TgC
a/SL7N3cmc/5EkdP3e0Fw3Uih/k6w8ZO7v5+IAUASnxKGOv9UsUhlYzT7pcCtudt
Z1cEg799f65Bksq7nqSgWKJ1dp1njEa3OV/vglB1zPefX7fTvccco5AcuE6EdGCx
qCLJRyelAlOYpH3rC/YJg33lrpyGTkxJT3i0Vn1GbT6CJVEvIR1ztAZ0woLOEJh8
dRqywvpqiBSsHDL68q0e2zvsvrpV7bIGRNclrN1qKctGSP3JaJ0ZcAqL17bNectR
ET4AWgU6ILtMPQqCRSZ6WVdaGohF3IFRALG9HCzz7s6k2o3NT5jQDiEUclnt/Rrt
wUiGfM8Qz1Ge92mbKWA1kqax+QLuDOjPkqJB95HoowbUCKVU6aenP4xwAk5rHQQU
RIqyEzazwH25z+sbF70OzIcCVkdpzb1PLRjK/aK5+KwP4QG9Yh6XBOsj6OBmV1zy
2AojoPt3+LoEP7hVJWpBZ58RDtJ6jQcMFeBviT72ZqytBqx3iCI5bXu43W3hDF7T
U8U4h56KqMAsFCvilD2gihRaNOYG/FzFlHmZGMy2RbuYtZCVChYCZXK5GxZAOoQP
Ks7fdeycjKwDNilDOKgC+8HVu+AMiZseF44dMtUlOpObFdVvbzNmLdgo3wak4T/y
os2EkWep36wiheYKK68X8HTQa9DhixhWOj3ZjluxQNW3V4zx/KboDdBSYNsoKsJy
hNegf/y6V2lH+4rd/AkXQPpDmY4HCJ4FrN7lXMg8L2KQFCVsjMcuzKfcn8X9Lyr/
OZI6NO19MiYg1eeV8U/TQh0KpRqLRhb5AXkDjn6wT3xKrYw9LKoq63sD6NwvHgkg
hxEwkzvnKwe2nVLBza6NL3mgjlJk3uIuQ/oGXEiVUNX7Ci4bZz+g09scny3189R9
fu85BczZ83+Xk68fjzNnEhiWvlXhRiB16OjHbNIf81aJR6HrHVAtP0tkM030UTAM
HPREZgfSI0krbutJQIy0ObxXdRh9GtQ4o20teivkyW69+0wPMScYJLJw4YRqtlAJ
HRN9OgbtS4xjy4YaqfQ+opfFx27Uq05XwaE3bqiuKkSp8EE8ZWyIRRfgnBpVE44c
RTptVUdMSGmdDkleWG/5WYBu8jUzUXLBmn5UX04jG+Wwaq7wCSlg7y5aUWnqbPdS
/cNXa25FDHmoazZNNsBK2xZ7+gqJmibhnkUG7SHfkD9rXGiACsWf3E3VD4jgRpgZ
7Ec5V18JSlsF2O33PddachDo2KOY/1eAF8Z/XUI8/NBmM6tVDAZjYyZX8EPEqFEI
0gt9Km6BB3csB335zNCLTeI9ll8zOXnmnvlLKqNre7Qle23+SIwa6tYFXlRo7zc+
JNk4tAC57rlXZUiC2//wohKNzfQH5Vw2bP/PhE7NJzF7Fp5Rb3YqGZdC5Uv+AASv
YusVniFEVdBYjy0BaTRmNEABRTlpFVukRsgquyL37TJO/sS7bu407uTuHbefwpLb
`protect END_PROTECTED
