`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i87qpdl3qjl2q7Zwsf3p3o3IS310YRB74dDGeRfakaR7OcrQwcrJP8mAyjIN0+Up
4+KKrxrcbxaTeA1zjDiHRYpMniq4d3Zd3iPWhV1H2xwa5mjQj+iZAXqOqwdYouiQ
8xBviTj+hMB/PAM9R3qkHolYuP5G0FU8/SROT1Fis+z0kLUKrkSFhhNCHcv89gdJ
jxftlFkuBZHdzwZ1TgQEkO18Phk0K5t1WF+6gSZTb1TfCKFRHE9GE4rCO2ZHyTab
K2NhucMMRwABRxZtkY0Iu0StG/ynDRmk8Wcl8XiNmtb+rI3Iz0nW/DfSMTMMT7Bu
11UZImcFuhO6RKnidSRhl/gZdf1xEMPNPXzHsvSukeuQEKq09ZPjChAppRIpTMje
FHlqkWUJh7VwtKHasEqn70zfTMl8lB/4M2+GbnHY0K4=
`protect END_PROTECTED
