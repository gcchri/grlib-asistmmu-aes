`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dfh7P1uo18LHZHK+RM+WQnfHNr31Gn8GL6SeOdyCpllMYcaNovgzsWMK5Qr1b6JA
jPbWcKig9do6oqDqbDwwseSpu9cp/zsolaNHEB1Dy0nX6b/ZDLFsF0BlKdSm5B3j
FHVVx4wBmum7ND+aqKHa6S9YfLmtKGq7OTyRCNC09sliMTKF7G/V5XNFeesa/s+t
PYlmm2eThFIzhqr4SfeiAdUzfcoGXpsOWS10wB9fc/UK5TxU6GgKLfAmXi39cNwj
gteEs53PIi5x3kBT8lo8kAgfxe3sy490I37njTcGxKZ9CEDHVWrtyZl8ZUVksmjc
gbI+LgIIANTMf9M/21Taz6vmh61+2KnLAooRqbDpRQowFIa3wxphR1DMRlwzXiE+
WS8xCBdQuC7tkXb/xJKNOYeTJ1o5q43ZTQ7fnNNLlJni+qHMPAxu/VwnqCLFHVwa
/sOWhA/67S6u6acc1x0jH5jTfrVCmy6uu52i7zEkN5c4604S/kLw4ZP8hrWNQDR8
R6KpyU71wWNDw54LAJdwsgsXyVUMQqk+sz8FwMmhl0q2DA6Kc6dCPQkmnJ/vKtij
vp4/0HubJa+Li+wNjumNnGcJAa+8dTl0seCGAzpavC93pGPS7yslN+ptp6vXa2KF
jYE4SrTx0vn4b0Lf7FCzB47A5Hyttkyy9lEf+21rFN8AzD3UTq9nrO9V09XuNg1F
q6r5Uy8bMFIqhQCBgW/N6c5ixKo2yvnKFJ4s8dTk2Bty1pNlbDTu0IEQbfVvg6vI
oKlrNYgOhCj7Q4Br1Ssu5bFrXe3ItsnOEvKPo0KFMN8K+ktxxlj/pGFHzzr4yVFp
TfDBiAAHog7JLnrIFjIwjewFOZN16/npXhVdxd9a96+WE8aLozsZO02Di3mjfu4d
NGCwe1q0LTczWAYfUUtz6+QmU4mkDarZVOI1zI4PVuEjgtTz4xQYhsspKnYrEtOs
uQ4j2a0URXWkrD5cuStOyM37suiXuRqFTNf8AORRRDxzrvc1XjCN/58w5sSn8sEi
JJ1BlyG8IK97VZUpdUdCYZeToHpxcT2I69DfJlS+bus=
`protect END_PROTECTED
