`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hf+ZqoVA2zNhySNDEuh8gw8B6LVUbiIlqHSAlwul3PmcpXLDruWZ8OosRgC6MKBr
OtYsr1n6I3KlCWQMAEA5IGvA2V+FPO64ra+KCnm5FOHU25ykJzYLpjmgcDAdEVEj
n5T/AzWGqgzCh822io6kHTzhKlmQwjjlBJTFhrazd/JUHHnSNtmAF/5u2yjmtLdG
Jzr6yv8h/64+lLgvCRpVuNxD+S4KpAniQSLIyLrtxAyCnT2RsVo8DAXf1/+RgWVT
5Uk5GpqRb0CCXRwb2WVZY8VqblXhXb/GSFaelU171PCIWAcrjk0dzpkbgiwR0dB8
a9xXDvpxwN8WEgzDQb90spQq4y0qhRAWU0UZrsYhH2Babu95AiKGf7DlWQcWg6CX
A2yhhx3y41q3GLwYsbL3a488b62oOXsAFUhGPVSnXCnFoWYHPSVVtzS2YrBvAmYA
Vz5C67nA/UZhcFZzPg9Ci+3MJdBpJZhwPHxlUUw5hmk=
`protect END_PROTECTED
