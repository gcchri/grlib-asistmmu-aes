`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hsT1ci4ZCHbEcCKajtTgHvewaw3iIBnGKarNCNUzAGxcNnQy6FXLHmsyWMnYleI
Ga4FVf4XUuzSp0+w/fFBfLgAH3T4K5VLchbsos8jfE33+RFxCmr1X9I8doYfq0ji
ZUMD8nDeAZg8LK1YXDU5bselGhuWQQv45X80Ba5xu35sIh83a52yj2JI8X9U/bra
JSNkxPr4R8sqXc2Jc7XdhxYe7kEsnmWHjAMp7BRrDFsKGFnvGpol4uVwV/kzNtR5
sRd6rD7rsKPnESYm/l4QyTucAh+04t5bS9D5K2jkzcXt9Tqxu0rEEQLajeRfKW15
+d7IelT95XCE6MQqzd1QEA/EfB52+tJRcW8/tmfiWZ7KZs9Pcxt9zPipxo9CAfg/
DdxIcr0hwRoUdPMaVilV/juBQvc1yjo3mWcAjFZCTiS6WnguuNWaCEFkNkSz+tRx
5oXMKfu5K7YqkeZFEARF8rqaebM/Z+VVJU5XNhDMACwJ2KZtrDq/2vhcKhZKTDZj
iziSlKIVSfxxFmLYAi2TWWI2wWH3GJ6FrlmB/7g/m5h4pZ0dyweTC2hkzBtcc6O1
La/Wa7s62WurPLhfkJJG5UOteBPU3Q4xVih8zeNCEwnGeBT7BClPtsad9h63gVvY
WojOH6pMwHBIodgI6dFqbrNDMnMbbOrWnMuJEoPyp6sYHVr6nSNzVgTaExJ5xTlm
iSq+xrMbXzUfAvOrD72CqLctSWEx8heqxBw6hyd1vNSxonJX1k9L5fBNsMoZbt7V
aAlUmnP2gO0oWbTh/5CI04teoWclVbbh+Oa8NdzK9+njQ4f1zwyKuASowUJZRZig
7NI+RS+POAkBE8n+h0WsOOUyUmm+BdOmVVROhkBfQiLgDz9TQxj6g5m+LF+/2eEP
ahBNOV/heSsKSgalhXUxY0LHDPYL8mvPuaud5OIFU66dXbUBNXfO4dmsWNmYceUW
XVepwFKN77LsU7GbWEt1HfwYCS0go+2wiQE8Dz710CSX0JQ94YaHjFeziKIHN6zc
5XPZXx4p6neLFAOTHcHA+V/fMDj+k+ot172W/S5PhQiVc1zmi7uB17Gd8gFkqaKz
nYRBgIiY3cJMCHH8sVi35ny+n8X6NvTWxai3oyDKhZ4jI1asl1NvbDS3eRWs6DMu
fk9qYyCO/ecFx6Bec6yIldJYWlBlLGtiUAQcgQPn5QOS4V1O7U+UAbwyJ9y1SkHY
DBGnwE8QP+bGcSGJ3iI6OFDUN10935yf9T75KNc4rz+tING3PIhIUnm3XZ4SiUMc
0E3FeximHfh+Yx7LYxievpHsfUCFRQO0Bf4vo+iYgQtndfHbmlikOMJLzxcdW48s
BZ+zp/9e/FACyRryBa9per2Wu9oZ33hY3EeklSuT4X6cm/gm9Xh8LlHbwJQQjXd9
DbEBJrxlQROOtQMxBx/ZMEXUwytfbEn30L3OBIPUm5NX9J4pJH10/cMDe6HlPYbs
3Ue2OfqH3ldfwdS9RUTIkPDUEigflTWAHwPE4Titjb7Z2QzeYnZlcgZY+7Gt9a2g
hytl7WE4UT5qNkSPXcf4wEJz7cHV4MpjG6pLjsDKlUUfCApS00wZLuyob7Zbp/q2
sXR4YK71T4FAyo8tnLwB4CMPu9kMtXPeAunqZGf3p/pg5DrRL17HT5leHJCklD2T
YYGZeJE7LlTgp3SOV3tvIFZJMiGqBZ0xO/MLqP54Kgjw+MJhO/lWSFlnqCtEyryh
3bOncZhM80wPhOhJW8DaAywEhIqUqHpdSXcWawYhC6evWZIFZMurDejdczlWGHp+
g07bpbwVrMuy212V4wPHsO0vHy4xonVrqSgZZHlGmoKusLz7/wQMSjcbX0kRA6on
Dbpnvvs7u1Id1c7TfG1nX3PFCcsPgr0C4NS6/SA04dsK7PPV4w9Q8enp3qI0cIN/
oOczRxGKtZihrXqun4EODtxk1GWeemlpOcBUfA5kuBguIPMDUOE/dzVVGL/U/xdc
rvAOcSsDpx8CLTSUOz6rEw584j4ND3TcF1xYPz4B4r8yS3iyAtqywU3/q4PYzK6h
GuToQMrqithhBUli07/w9BvP+SrfChjou0/XTzG8tuCgoj7FNG2RVxGFThVdpHD7
7aMcFHFbuLpylbqr/aCvyjMfigX0c+KN1lSRE5h2K7AQaAXgSznPBMJ00jRwpw7N
Sti5RO3G9FC7weZXy2WfpvLYrn5AzKdU2bmC1gPk/2SDVN1KYjTRIZ7BLWeSeQMP
9kwu/DEPHVJugbGIKwgpyA7lE+IpHcWfonkz55GT4DeGWRiSoNC2jTfw66PsA7+X
nZcC3w+QAp7CzpBLhEHav6oWRP+JgXXVR7vfnpmu++u0Hj34fr1hXeve0spaWrep
8a5W2Jns+wBGKXzlda3t9kiGfo9t79SYQQ5Nnyz0bpn7A+Q/n4mZjcZnaDLm5wQF
RUcYIV9PtSg6ZMdPo4kP9Iz4ekgigVrWVUpD/aDeqTY9nIpxpPOJuEouQh1IXWe3
n2MvJQC8/OMIyhcQOI8GmAKNQbc8WpEbm9Tx69QfpaQQZ++FqnHDLLFTvufjehXc
FlgugYWGlf0YwcBCU3ELDH8u70y004FEfGIzWcIRnbX5VzfWxuKAMc1SgdieTuJs
YCLt7+qjKgXKj5C1CDezXCLr6HM71Q/0sFK2wvFXTbQuYsgWpM8hy/ArzkHuFwn0
/5THtit2DpNd1CXPgQiwLp78eW9x1Y13hC33ZoololdNiI2tl0DE37d1FAHOw5g7
97zwP0bomKwE5w7auYYtMhdDy14Itca4sQEP2nZDhV9CXzsEiF+3EQLqZfNSs17w
aDqw/e8sjwkmM0O6yULnw9Uuxiwx+dxx0rs75IIWwzX98CVKPM2Lne0kNGLHaIsz
2HKSaPuqsAuAECnXUK7HSTtUUJxlcQXMIwAYxa0CbsvXHVBYvMZ10l+NaLld3NIh
rGhkaBVqJ03QU3nm3xxwWjuqvvuOlWn/TOHriEXns/nNEfTKmCka60n6PHofsb+K
RIGFXP5ZZDKZJXm86t3rY6dwwUvy7CLIMEJKOpLgvJVo5atLVwPdoIAJlke03PVl
srpzPY+38djYxAYdmfGkITVzM2jyAwe243SBA2AORP+aMR5xGQ+i1d+fWBpfuDPU
8azEhBOsHuWZKIsX+3oeRCm/PZOFkxYMJfbKVtLK6/kLpEPOCuDr2o+2Gr3XoUJn
y6SglI5TiwHG3zqanFkiuXyjMuHGOwKEwaIpfd2rrdi0BEjFEyCitmJi1+uOcLIi
PQR+4XujxkM91rvgu6XFl8mduWe10v5YjlekY8G5h5DZ0WLgZ5Ly3k5Mnng4qSzu
zYASolqe5cOXLuF3SXWPSCUsvaymAZ6TIWHmcl2d+9u6Md7CQtib0gui7MM8b51p
xzaVl4YTYYxOz9vf7IcSRUVu2txwx+dDWnfUv1ELVu6yBQ7Sx6D+srQZMSZ0Zr/j
swxzCt4bgun9GWsoQBxI0bMzOyeBmNjVwqKTfShrszYiWj7IRxJVKo/OGh3pP+uN
IqH7fQIP3ToS0VwQRlfRoGJCjXhB2ffonan4bqxiAbx0C1cCITo5L3xid7OVAHsi
YTYkmjhTPf853w2ranEfsRtF0UDpOW8gQauHjJYK1olHgFDLNr4veKfwlBKMsuHM
IHpmu6tSgzrBFzwrAeQaOiLTGXv8VDjshMphN0NAnQ5ZgFslcDr5FPOFSffWmSel
Gq8mZUmTfEqOS3PBMTtRB3RovFgB8x++VAekZR/y5MQjS/wppiL03g2IXQyEumH0
ZnUxiYjEN3P99kWyFx6QPtSs8Te9SK4cHZbjJ9092TIlEROn2L/AmGcWp6DyxFpo
55Ahu3YiX63Ij74pF2S1VXv4HKsDLBi+k8Eioy/plh1yk0BhB3YZ3pHX1O33ZtoG
7h9jhUBZvEngQD4nEceov5uaxjU81f2Xy9zVpD+r1ZNTPJUMpZTGASPO7/JB+HHz
gCP+NY3ujKZ2FiIGlwmtz6Qx1uFig1tFhpSFNZSVPdfztmhvuyz5sfOvWXpCX4aj
Z8tdXvRDYCZ4VuyCMwgzzwa7lDKAxwr9invxrimQsecyfdOCsqth3TQ6qT54Gd9x
wwixat5/uKO6zwiQTFTF2oPa9849tk5KuUDAGFf3rK48tB4hMALyCgm99hgP2Pp6
ukdXP0Wjj5STGM6EbdMqoNSpM/7EuUhM/Pt991sFO0Z+r9I2GiV0opWRudwXY/OB
AJ78lgy5hkcCafXKZC484IeuHhFou5vLYcJaXOfniiGeRPluLEeLXIBAdTyWFabm
K5n1vbZdNASRkrlgBwff9ZNEWbjsarFHaJsE0iKSlXPUM81261byAWgxHC3OrQm0
j+QL0KHTQmrC3GQ8zodATTaG3iYGOvbyz0oEwnHENOtm4EGYFzFdiZE+MxBvyaNe
H7b54VUqAzAmC/z8wSWYl8IYBLY4bBn+rn6BF0I1gYgCc/KAJJSDc6wp11yofGf+
fWszz5HCOZXf91JN/eUqKdgdBGbKaKUGhv7zvGhCEP9lNJVA3Pl3rLODayTz6uf6
z8zE8fx/hq0jseLQGiG1kt2aB/6LUroY/GcaJLq+pMN/SMMLc2qIe4f9tB4ajyE/
3bKDPUlW2dlXddt7UCFbBgzD7Ls00mvisq2LNE896drCDDycpj1ltuB722yOxE1r
0Y+R/57in6UIG8zBJZAZTDYKjP/uIrcm+e4MEwmvPDVHpQ/QjytykpNlMYBzV9Rp
qV7t4VH1VWoCOL1EX/psmTOPY4ZvW+N5M2e1BuTYzx3MYiqTAyvNrszhhFg4zDki
cXWCV/8BmGomormZKljHgd+vo3Bk3IT8frCozr4I7y8XZ9Dr+7MiFRwVcG16WiwK
SKrLaURM+6cyRv7awcM6PfkFdsFyFduJoGj2FEbuxNx7yzkiOLMYenYFw7RoaYL1
KbaedmLCtZg92cJiHKxk8P7ES3Q3Ua0ijJzIHGkyAukmVZGhlpy/qeEnXhKqNhLx
O2eEqfabHydTThUQoCInhiEtlrAzjmhWjIlCw0BgIP/PCAqhw+v456VkAjbqkicn
q/MMmvpOamoLX0hH/1djLO9D9iE5yX+zJpdIgfNVC9J3qkLHS9URHRAC5OqIeaRW
g4lenXKCt59tZcT/jiXOAAGs0nhSx0Lrjt1UhwfQzVhBWZZaE6n0HFcb4hyr9faN
nXu9f5weDD6UXzTcRNH/hPA7LPzhAQCvot+95+3mXyPhRA6G5SJ/PkjBV77Gs01P
/QifH9ohJSoouQpDkzTZf1+KnZdbNqV8ADYtCvWiovobHAkON985RmavR0/nGLxe
ocahDAwYAKeVRrOrTvU/Tbw04KO9AC3FPpHb6lY6+4ae3EdYb79IUe9LKuDCHb9m
f0IztqlMSiYl4R8wRq7dPKhZ5r/hdDOKnwn2ImD8SdsMZBs6WslJmlfQLQgmt0Mg
lgu0OppEimPffemxWKtIkXVcez3i5HD7zcjJ0j9Trh/ngBE8SwnWvxJ3jgc2unop
zZs6sC7D9uhligvuHlIMhYQDk4Y/z5EzkhdnM54ayE1xZovVwjQ9qqxWtwkYIGsI
CVSIDpVZE65ZlORGU24KPkXHpEr4c5GkHUXKUep+NgjvRGAFgUcrTA1TKzqQV2bq
LOF68qmqod+XmKyhpKWcaEDAtM6lv8xqsD/KDyem6q8CGu4pdFnIr9ATOq8SMj3r
7xbmHAdSyvreG2F63ZZb/qW2M+AIZDrc4QZopm+bWNHe8puzz0QPsp6pf0A3GU3+
hCUfr6pctzgj+xqYEF5NdOOkefppN7u7+mv5Lvpr7nzravT3t+Ta0ehGf/n0G25T
kwGowZkv1QkX14ztOPS7pUr0/0lE5GVq14elA79jHuF2n4FOn+yOiBRE1G9sDASZ
+NneEu3zUvUCk5hrA39XyOE1VOS4lp/3cfnwVKEyiMuoA0RHIxDWDqWri1k8O/Ai
hS+J5zfShJNgklO7faftvL9iqyj1ug1/mnIQlpYsbzk2v/OKFsy0IGd56dIsusDk
BUH3zbaDzgS7CCDeOdPBqFJ/vIMJ1/r4KhzFcusHeesL/6fju6wPdcD9k5sZ9ujn
4yOpnkC50CwRfYngpOfaCSpUJgR1+qgACnBV5/xqVBASZIl5PsfMDVF94B7YBfoa
G6ET9EJu7DAAGbWdB5iFnx2UhQuSzMD2W4WGdeqqc04Q4sELSNNM8jihqR5x0qob
FrMpWNrXoEtRAtaNtkAX22zZIkb3Dx+iTpJS3o0IJx3HrB7PKLDObe4fL6FcR1Q9
RZLdzA4mbcQh0Vv0/80F32M0FLVAL+/bK/dkiELxZ+w89dOi/N1L1QKc/DHQUi79
GsETDqRLqCAEIzuYIoCRofijuy3f92h6n+i6C6/gSgcG6u4KrQUlWxLvTf8A0eQ6
L80fOOQ+6g3elYloCH+vy9BLAc6DK9g+oKycaNwxJpwgk5A83ByAZ/NRFkdim8mT
VwKW8XE9WUN+KZfZYQ8VpXHrYzoyHiK1Qoib4lmGcug1AstBfinq9z+U49be7XCo
npbH0bIARe8HAOZLshilSAvUKK0+hqD+GSlK7MpYv4ShiJWmEIJOUsvSZOVCj9/r
meD1YM6Jh3CN5iYJKvGy/z0rmt9yLBTXOKVtgf8NLA3e435fPcxjjwTHUl81zuhe
hyM5EifcK1GvEU4wmFaV4nWXBotph8yVMxBaGV1F9Jq3lLj0I2MTsuURdnxUaJTw
/hFCEMoAfhxqg+Eu7ann9o07Ns7uwczqM/k8tUcKgZgXs5kUa4P0o1waYO2zXJ8u
l3aSUQkgsLsKisNNHpzWG/Av53rB1GDtttH7Bw/FNZS1xXevTnHwHq1GoARmTQ4K
nxmKuenyqtJXs2DocRad7uqq2hWGvWfq8FNm7zhM1Mu9SqtiBh4F7FwolMU+JCpr
1JPc3tQXcACI8fp7FPTMHHiCOwQje3ECff+XrCvE97IhAcv6lV4yb1uFlqya1+2P
ne1TD1ZabuaLe2u7pGrQPJqLVUGwqzx7UZc1IneNzaovVgkMQmXZ1ovRCC4x1dsM
U8DdKGEFXsOMbFSmtQwOFom5+UrKu5vNW8g4zxCL3xbpm8qkNU4wurmBephoWLH8
T1qZGjrwBj46udpxBm88EMdJZJJ0iHl4tWvnCuoI09CQirN7O3ZFCp3eei5Pq3+4
YvRd7VW2lQNlquN6ZmQurgOM/mKhdsiPpN/4xvu5EfiuOfZu7zl3i7ShPCDH1TjR
h1gVJi+MSsUvnSMDvprd1WUHa0ykzB72OKWetEHF21gnDlMzY8IMeEWMV3Z9/AbA
aCNJwFvxbbw1+nH2gRCyFz4QnSMd9XP8oX8t9HAqlM8NMMunDEODGkYArU9X99DV
FIP5evchyYENf/KioI3sbSkh4OA44eMnKPZk0LsN+kdwNXURC+OIUmVeU74zo9xt
pliABp47A6VKXotP68FwHJ8rxr/XD+xzfBsUieP3Vr7A8tHpUPbkSz7GWonh7gdZ
k2b6Gqbv4GyPuDfCDVJS3hbiZXRxYLp36G49Q6U/A8dLW/BR6+aJ82UV9Mr3nhRA
ullc4aop+pTZa4C7DwZf85d37d4L586aoYlzaLh9wlJJie4udyx9Mrh5SCAG1a7g
n2+4P1StAqyR1wTzIJUUa6E7PXhMwPC9AU1FMBXf0XyOQ90kGrgs+lgxm6U91Bym
iYmoZi+/K+pUetEeVJ5zHSzbvAzDv2ROaD/NXCBhSr7oDCCXlbDGvUzrMkzsxKn7
nonuNdYa3gOMpki+TLxk/DTtQHdfG8uts3IZg2Ewh2qtBO2/Ort20LGF9Tng8LwF
lyJyq6cMe7eM7Gg/7CGY8MP9fDGTWV4ae9W2DbRlx5ei8OFgclldoNsSb65XvzkX
DTKDNLphh6DCSqkD7uMjz8ixVLV2cXxH756VD+batym4fYlogxI3sRMyjc8gjMAJ
9PVUYiGYiKJS6McHwK+2wrMKiNnYMsH3M5GkitABSKnKdti2NPhkZs/SYubLki5N
7Y80Yc6vYBw3DtQC9vZZEftu3pdCO8/ue+Ntb1im2rTXFL31behVO8Z93oMS0OTv
+hYbQg5jbhzVM18BshlswkbHRnNrtFr0gqOjUAbZNRpUWI7+KLBCFULi1vXv7xeL
K/zS4MsDjBJnGIdJdKnQT26EomjqduwXPo2tQDrsoBigQvfRbiU5NYnhmgV1bkuU
cYWdF3g2qbepP7fWEfPt9uWellv7hHzp1KZl6HcjfuOFVOvvd+eJYBkBbxL6Tixg
sD0sQyXITrX9sMFpvmLM4e/eWmq8i92GmZPQNfWoVwDsGg0pBYPa4qOZPPnrdPoC
qHPEq2dwZm1Jl+ca5UdmqAucbeEBBXumnOtqkLXWlfyzLPSDRi2DAWLL7dY4IIh1
k3jYlzDOgXwTfzUG1jb2f6Bed21tjlTk0uDXTm5yJQYnT64cTtFcrN79GDGRYZSo
x4fm3MQIlQSmEGr1oklzGtn75nyDfeM7Go9Jjs+yi9L2YQg5V+4l2RX4Ti5BTTaJ
wJqnU/KNvpyHakgvMaVpGyrKu9ON6SbbfFZkig69y983+Afgy0/j29DBzccAtfei
hlA/TAehrsVc2ZYS4EiMB3wBKCaSxzdehjdPyz5VbeRlIpkCS7hbCRewWwgLooQE
/EGjBvqsMXFyHf7f4jgQ5OTLiNWM4QNzoJ5KpfMdodQkhJUSR1c9DDY16PU8hd6B
VVNY8w/LllbIC1VmZaFmp4OMKKOWleJ0JMkD7LyQIVaBLR1R0xGENxCgkX2AjkfH
o3YEuCTbUBDsZpGXCc2xA5BC+REqCkfFXpOo0LuP4TNho/GFbXgK0Qx5qoWvlBSf
Td6eHd6EbFApqQIsYb4SFR2RT3w9M3/rYT3Egg5T7VlF1Gq0qhEpjUPpFpB1Xk4S
n3kPS3rM9FtS40Fy2LdO9aoOmRNff2T5eGkeQ2c4Op1y4jyvPXoDDs+GCGqlDTpv
a8uIOxg5Q/JQZhfZvvvUzQdObFPzJTJIAsoWaRXvp3NBA9gUjbZQZsYv2D2wP0JZ
ZWG4Eil4Rj0BVk9cqkKsymgtVvTzlw03jGINX54qCAgahw0N3bPlDfq2Y2bT9c9w
c90BDrj3Eft60uXpZvZlXzKtJWzPc646jgtc7pV43sJNz+UbTImFXMNYMkKHeydQ
xjntLOulxzHejRpkXcGJC1h09SUPQLPwQFjy4AXWRjBEc1E5YmL2ma++J4xL4bED
jlntpWqBMGh15GnkNemfVc3xab3wGsdMQ45yYNNsZUBYiWHPUV6gbbsj7KUFY3zt
6tQ1K66Bq8ohWMENuttbsCWmifUpiv6UVTFvFwseLMRUX7L8pZviS/oyrdufki8x
cDHwOZTCI/GwYnVLA9gOnv679kTNAs6Rc+FwcQOuTPVZYvT0GGJWLcB+XrBUZhPH
S/8/sP4NVLX32tvNWRds9Bk/wBUaIX3am7pwIL8J77rs6oTYk3Gio0s7+GIlNgIR
A2ebGGsxL99OxAAq2ZRaGIKAPz0ZqR1XEzPmiTL5YWwqGAdDWHBSq6H3AuLRew+m
e1FsAOm0xm7kmOcPp8p52Hwc9YBvPeLaB64bVPqm7sjgCGwkfemsfOVu6hMkFkva
gHyrVMvmNT5s8VQgInnvB8eI+3wAew1DgvDO7z8Nu5mI3ebuG3+xNrS50MC6+dzc
EW+FvPOGoR0T2oW2RByYCOjTerPrJ+qMHf8GTAPKT+rsjPWVegS6ozTnzExYscnT
UYE0NRFvb3hntLD45oMEwMvEC9wt8VyV+sVFhA/+eRh1t/ObAoyZPo2xHrzTBuVc
3OK8OxKUEamJzNpbprqmHvkN8mkOtJbYAuMdAiZyZED5GfgyrGFozONru2HTv1QW
n4QheBvB7ly43wWyGObE0nKnTw1wMIZvNTF4rjRlD9YYlXiWBdilaBXxt2dtUVOL
Hzvk9CAOtG6/4qjIEAUytKaHIOjv58dxRCEQgK9WGj1UveyYjkh0KlDeD/JIQBBB
w6B5YzGL1RjwYRNI+tBN2dh3s3kB/77JW0TnvVQSQ4xuXtFB602rc5D+OcRlTHqb
c9bUyoFBEAihuGQ9MuabaS3vxvFWhJuplzAMP8hTFkchgFRaK33PRN4x2JXVbJOd
r6yeIHmvBrUfFDuVm/lpMUizggZRLimdXKbKoil09z1Z+mXsdgpclRWl0DyuYQ0X
VRBxgAYd2vVw+UbYJFgCKT31eBgmGOTUyewfhHjCAn6c+6B/UTZiRxqzwGe3Jmca
61aYrUY9Fj0uFPefwkJe9ewrCo/6gp6wbuT0X9aHlVpv74u0H4W05QXxWR+NvMNp
XK59CFVbzsWrvt6jvKzr9vOFZW8dEAQQrccX68Q3C7HhW0Ap+7AdgXi0ieaNbnAN
KZYcyYJLcwHdWzgD7A9chJA4OyMlusT2Q6OOWd/32cIkl8cVdpvUAJKONOPnTXjB
e4IcjVJMc2tpEPpKnqCdNSCRtARw4c7A+m95PRzlvcHGQec3mZSrMkOyilfVrBG4
Uwe+jWUCxmEckDv+ZWgW07Slwm4f4019zKiPtEX17ttlPF+XcwgS+gNKZdQBJrxk
BBvrqRDsCfZIUgzWN0bPDeCKjnCAozrCTxdD1x75d9ml21+FytsbVBAKEcSE/h30
NO2nuYe7tGS01TytjFIaTtLp7vsngYxgFcVgcvCngi02vEoQZocwwGQdg4APjWWe
vGJ4t8XhrpeWiqFBtlBq6xdDLc7LHppzsAR3NXeXcNoKyVB3gGhIltqhJoW+sAID
6KT7zxwRvLjN2pM4qao8ZS0svN8QiS9Y9Lk5B2qOa7nD9MlRgm/FJL8hfT1NXDkT
t4+mGDzQ0mDJgqdiuejkLxmrJ7RUXK7QoErc8xOCd+19wTAaEwRMGjb8BVqCCWPV
8XUR5beAsSZFzFWDI0PSxL6Xg8dbY/H9tFKLH8u2NU3VLOePA/aYhmk4l/59Qjnd
gjxtpLx3K2h5pDMdykOrScNVI4WyMh/QomfEbjN3u0GdL3AIOsh1oKqwyC5a/PG6
tMrdpMjMte2l4OlnvGpLBG/OD23oHY2LpejohS+YkWEZv1DVM2U72kGgl/amyQ7g
7lUwyOwxXXhkH7GydkcjrsrzqimT+qlvWytb2PhF/RZHvKu4+dX3zFFWzhgQ1+pA
+98Zlawk2hWz3iSfcFMgRPtv5ab31v7cptLkK6ZySA0v/VipEtOd855Gu5ViKm8W
wZzmEyb0YUxgbHFoMEwT8InkFMQkVI7wobox+9f89KIc2okudtWgZK/8ZSlgAEWg
RF8NMCAnmOzAzquoUQzR8JrZ2dfOzw+htcJWPRfnCJLEaR7gBLABIfAjR+uLQmnm
OE/bo9r9FNLH7n7kxszNkqaflOkFXpQjs8A5KilyD2YAGnTAE3M1sWSuNcVVTbtx
6YRbhb1aTBO+7SAq8BUDvrpqjkoee1DDGzQ+t1hywcQ/6hlxL1TeZEzIligr/K93
SahRcxrtoMux4a4RP2Fr5KNQQwc1fkAv7CHY/LKDxyKgthi/5ylKoxfRMLUz/p1F
3n36q8nXW9huwms1atiFxD1AS9aHiCz4a897wKeopUVvBeQ5jjuaNI3sKnECrIHb
N12tMYAFzm8Cd4qRDkROpQ+gEIkH6kB+DLEqEe0vFXpcPNXZprL0AqalL9oZucFJ
cwYYfAAiW3eBc2531Ob2YCRJItUCnbIhGgJcDWTZn106YB5E8s+ozX1pVbjIOKnE
iymCUz1hoLca7UYpTy8a14a2Dp/8G4dIGFIH0iljw4KCnpZlgYkgGlKlf1EjFWGc
rEbZQFiH9fVorF7Jjm1YVm/467PxSabfGoHKhr1s9yur0UYpdCSxfjoRvcmQ+pQV
FV4Vg5+iwfI8i1nl59D/2EQL/RCaIvbhrH19/bMiWRKTVMwQ3yWGOqUygSIfnDgz
psMaFZVMg98Dfh6P0IKkKf4c5lZSUbVqz7Ac3nVlsd8JO8JKp7A++JiKC3VgpKxF
C5oI0h+CZy49ARwQMe5oQlaQ60fCnB/S1DLAakiMvOBO/W9CCXTpqeq+AJH4oCG1
yWVqnniJxEQmRISs+TEtV4u6xvZf+btTtfnCz8aQ6mYzPPiXlaKL0xMtV5oWUPWb
UpR69r0gsLaqxUKCfwQv7/aVzG6dVBr1MeRp7hMXiOHIefxwSrZnUIkzpBARcNtF
Me8nvBpTwvP0FxCdm68K2498HoUzwInwB8CrtpbtBX4teo1xCb6bDzksssUuSmnB
6QUzXFKrl7aAqbGkQ/0Km8uwpLZgdaRrkHZ8wA8TpU/U8xJYZBhdkzXysJeGsrNn
WLys8CvThrABzvFmiIBnnjSn/n5BYQMDJy7fTvikkPOGuzuooRxDFFYXzS7CBMZP
LUgF0+txL/uynV+aTJhid3hPw0HMos2mScQw6pjwo0tQYN7gbfvld/qVFgNC5lB8
K5l/EtOEpQs/pKQmWZEqqR7pAF14EmcRj1gxbLGXQvCibbNjpZ8EUj4Lo1ItJOCB
/58mGM65DHJKJaTn3yHFvBKv2tOgvHOxihNH29zUiNonQooDo99htiYzuunHz8H3
vZpUqntOGrn3dA7i/P4RvfJcx8O8ETtnuct3BSEb7NmaHUhhsaSVtWctua9PRcz6
AKEwNHWA6rS4FWQIAr6Eb1h3DE0K+LOaO8AnZc9PIUeg4uj5ykMzRQKG8LFHQBfg
ecObxqWYc34dcqWViyXS2Acl7IcjjH4M6xRCRxGwz3OH9LnU3cEfBfIYEdyg98YG
wdoVFWN18HDQP2LvDjwquiS4cuaQTGFZHnAJzdK9Dck24mtdxMJYJQsYZj+DPIwb
vxj+kFlkHHZjKOFUYm7HutVKLkpH4P+fxgoz+ZbtzOg8MATk5QM+FoTJbZBnnnI9
VTvaWACj5ZIhyjLy83K8C6XkUZ/BO4DTMpcq+Aj19YrqAdWwwJ9SgjdzkkHUM8uV
/JHT0dTHJvc/is42mIiY+LhDoeKQOtzyMEqqDbx8dD88vLy41VXY4nAarAVebyeg
wgcqgzHcnorVflk0MZfgeRulx5o+uJMS5qZLI7EihA3k9DPX7FO3DjY1H71Wersd
JkivhPCxIoyJ9npNee5OOwNkAKyxD/2devW8ozruXLrUAVrNHxO5RMObS1aM/5q0
LOfZn6FJDM7En+9N9fvP3gZniG2m3qCOlUad7/wHxQ+g7+S6hMe17NGB3Kd2gEne
bK/p54EWZzz2+2bVdHUf5h8y13BQ0rT+xbcU2v7ztPFcxZp/i205zSrMrCtYFSJt
SDFnls0s19+ko/oVKsLw9V8Zhgx2k+zqEXTP1EIkXk+spMIPBD6YFL5c14F1pgya
nuj5r/Eme+nvkYLP9xIRQkWTEiHCJT2xNj1F2sLRQyVk9SdyaQWsKU2v5yPBVzT2
WuTcIbU/ag/ENQn7D6pwlJNQb5aTqoSxPBiQpp2FZAsI2fpVs3dn22bQQR5jgbwd
0ncvtI5+7YWGyb4maQA3LmvSlG9qhNHmCuOQUQEbbOEaCtgO/SeprVqyxq4T+RiK
VC1w3WjIdQAAKeSFVTUbhGHDOoY0Kz1C4/EwFH4ozR8NhqZpF3/ZHCYw9ewgWWxv
0tqje4ob1VmAsmLLcVqxNNOua+ZK821/hi5iKf03ZkRkcvVCeTw12m8Ul9Anavgb
3WIWv21mxehCCoJvhEcNeUF16zi2dPeOKyRLnNqES79WThc79CWC+w9YOeUg7cwn
BmGF6N7WI0X8Qua+8Gqqfk0yHjUp6VrtACwykctrJz6H/KJsYS4cSi7RKSaSGb9f
0P0uhslkYAx380UoulQdrVVeTOvqIm2v4wXsZY4WMSGq+Tz7Q80IWi23g4e+1wmS
yUVu2K7Du2NNwMK20dDyx+Z9vYDYPhSiuBJrxamXwfzc+Kn7sFF+RsbkpTMnu1W1
GoLyOmkHGRyHOVKzCjrZ7cAfGgkHELntvant6csJFFdux5dD5gf+gB5dJ1ugNHD1
wnoOQeLwguWTPe3nDL27/1RQ+Ta3kQX4hMHEHVMj+8mv0m5bZuvrKzqFNXOorObG
HAYhMrXsR7dT+Sy5fHRlUYva9CKpEGWObSqZvLpv504Y+8Te5XfLsappOD5csDJT
aM/Jt5qW0Ok5kDIEa43hDeDTFtMCGb5MMLmpvvsjLKCZhJ0CuAshdwtFprp8+Jir
9t0e+kiJpzmBGcZ+DktFVGQEINbvfj/XOopiqO+MIS8AlfC2JqIju39K3WNMqxZi
gIEv6pObvf6MWLpQUSnbp6/KYNCLeQKWl6HKzvPTg3zRC965GwYZiyANNyCCssp3
fhT+FkCG8wIKRfzvwbXQXD/Q4tBa+LLYzTgD6lDTIMKxj1FKPx4RYQsiRpbUskj9
HgzzcID/b1Jh4HadHTQiCReri0403tHTD3nBkWuvcV/KtC+qapiNrdc52Q9jiiui
tEg8eXgmi4IhruAk/nTMZFX0epbFoMy/6aF7RdKr/lao49Xa4QdvkN1yEMgQ1T+D
UBtWTzIQKXzsy6bAa4rCl4Yx0Yt4Uky3zQkuH0S48Im84vBpoIhXjEPU8QSeO99+
hq+I5jCCtJAOc5nbeHsstJLHF0s+DPea2rSKTkwcs1WBOTAq+HHYNuswel0/2eyj
GNj+Pko6M4lkwd2JHUwlWQ3Pc0eQRPG/AXsTrhB7hPxuikrAlyyBdCzQjEMNrFXH
TH1TcWjVyCGbRlHk8A/aMiBxDDZQi3YYKak5OBzcyQiiS1nDO4THs4EFbk3oLDzC
asJiNZGtQB5IM4PbJW0ELs4X9yBJC5QCqDiOIQz5jLBDVuChDhMDu21plZOMuYvs
MHaH2fDLhNTkM6rqSNVI/n7eBcK/qlPiGtPlkgZRodQ9h5egDpiJ0zs9/PfXfTUx
8qNpRl/Vmk6bTVf++0LHHz4tjIKg3/mEr8U8EfR6r8oC0cTOIFUUNkqYmJJwUeMB
/NC6AMLqUz1aiYFMzgy5H1n/IXbYR1M1OIwOCOZwzQm3O3f41BreDhwFFneS49O2
HggpVABBJ3lyFR9q5z9qdTQzzYa1njfBa8rXABDd5c3kV1rvcittcvzaQAk0Nhyb
fmTT7An2UsAkERYG3hrwUdy7XvuQ/dZQ6RJXqhJ6ZR5iQVSxr/m0vVhK43NbZI2r
lO87JKsUNsRpM/dRksi3Zpa9PEebtzPFCLq/drULys4E9YlcghCvJ4SpQtM0Q8fX
MCOtFEldSsAJspiKP6tohiGqF/SVGP0AiJCSJIs13UW2csOUUDTGlERy5fFQzeOA
HWOEw3GgATa82DHTbYXil2UrM9Lgi9GxkSXWRRFIJLTup+XQ5WLfe6B82rRVHAsx
wYDKcdxRUFJhKYU0TCRao+m+FrWBkJKjoaJH+Y42rhLhNpO5s6HD/S5E/l/EFS2Q
L9rQqd97pKlBceBuxgdjz0SfyDTa+zGKKMO1017YvH2tf7aYcwl2TMyKxO4YriGa
xWA8fQerl31DPOTwwlKkUz0ngtIm6lNzdNBS+N9sO8e7TwnpBwMa+PJ1BY8pgMKQ
jafg2QjthysP2psNDV8nIECrjS9t/nJQRswpnMnrYH1p64y11RXZ6w/DConsUupC
VTJnZDEcZdmQEjMk5xGKoNGOtN/ol761wRBQf5Z2UQpPlFCjlwAbZuXF06YjyN6r
Kqm4iPKHEkUoGaA/uecaz+86+GG7nbBFGsVW/EO58MaEHhTApfq0mEvarTJisy2S
oSn/lmOXH9ylsLpJgXdaXcDgvIBOG9haOr9lRqKA+4xaU8Nla9hZYeN2Q1I6+Yhr
Ci+kmYGfkrKxB+DYUDmXIiZc1bplXtGgFEvt3dXKRry12NIiwijZMFrqLv6wridS
5OWRrKi13EHtVS0+zAAidHi+E60jF9IwYlPlzvB6RKLUT3V0wgbCaBzf6u5brF/w
3fOxxoGnVGDnq6TwKgqtwvhND0TIHAWoMM8t7BvjlLfUdznMYwgEQ7eL8kNAlNhc
wd7mKm23Zq3Q8jSZVZhT04YKeMOD1HpC8EESwp9hSpT8C7KZs/kKUTmoQVPGEwGG
b6lZ4gp1GZxH3n8RKT+zRQ26zm/y6WoWZofKlVJt9YpZ8JX4XbzAXb0NErfzhSD3
Gjxfj1j7kJDpInEfBRleaXypLXzEHm6/GNt+r8UVWO8Ze+w65u4OEVOMQ7kK5bG8
f+al3NejUFaN9313etRkZ7D1v5q+oTMQZuWu5L8HG5vu/pVUgnG8o01rdYDc/DYL
aRL9JsVGX03R0eFcw3p6ZPQhuuJ5kxg9GmM84/dzbQI3CS0yHKrRKbHybn6Z85VH
lEMu8teJRRJluktF+mI5K5k0gvYSB7RX9vijt3lmXgbTpAIrl7Fcx6KJh/rWHOsN
svLRi+PkGunERNMH1iyfO/xhwF8+QirMnZam/jxhOUPFD9/JFQN6iHT9ubrGCo5k
fEWKnCN8qaM7kS0tMtEW3Dq39PJ2yHJlqIy2I5Qj9KuHfPj/V0txIPgvflu7ChHP
jWqW6ScSgGmCNeIjiUI3Ia6D5JpMJZwc+r8ol7tJ8vw18hRv1U+y40EqEl39WCO/
4jCwJG0Q4ktbp4g22Xri18oFfl0D6rpJDByb4kG6sR23+ACx8tA1zAzJiS6OgKuw
MW4UDgdIxXcOrLOppB7byPVBeSfHjgM1AoMBql0kbkCC2XVqLQLrQSEEe7npc10c
e9ZXgj8UikPReqrTFnvUmaFa7NmKub+0lQgg2jiEGlhaO9RHTtstm9DoelS4oYDs
9lj5QsYwUj12OhQOKL/xJzu3sBe9CQXtIkPki+4vQoODtgvMkR3MhfKYK3AffrAE
NFHjkNmkFv00wDst+sj9mbH9om7tzvPRHKZmmvuBZ+oMI0o79/lOJf3uaRZrVlrY
jz0/H9+pXGGQN9JzGX0ozZuJlgwhkY8fhkqxHorMP+MXrMjyGr+4317bbKUaDAzc
isSb+zUmUmd0A2F0pOLtDnxrE+gV9yz1LfZY7ViVK2TJWa3thM5gRSPdXjXLV5gx
wPtuXU9D/egrplj+Zlot7xUbm/LSsHb6qjiaBTCyf1BOFT2OL84Rcx7rkqzfFrks
wHVkCWZlWtxtAF9kQay7zvX5cNSCSfJ9hVSO2WeVz6+J9D+bnHFyAVjCejs1jckv
RJWONLr62Yf1B5QStoq/8s7MUuuCBRrjpNTfKkzuChGhGTQHrR9vSiC9jej2diF7
2DcRXjRcJuOCvmff1Wosn+9OOPglGhlKIY8oZOfXhMHuyNCl0m3h4WyKqe2jlFrA
6V3ocSovyKO/QelGK7X/+M4REfUywHbZ0luV6mQ1Red6qqp8jl5yVCTxcZd9Y/F5
iaimyuF3+DyG7wvTze/WEobIQbpVYsjucpk+TiYcpxWrTS4mtsSZKsxba5hpkICQ
BNdZoKPRYD03Hv+HcAcEhs7frhIkQ3lyJl6KW9wM/DosE7Ra4w/7809EDg5yagnq
t2ScpHofawI6+iiJhSg/QQd6Y6horUZi8gpaGcx49tdBthM5Kurs9MHBstmwmYc5
VKJA1WvSJoSApnHun07ZiS5p7uRymLcbC09yYpMjB91aN55GMvwOO6eLyxzhN8+J
fMmqgzzp+X2RcnBBUbExQvge7DNEE1ovGUSJoBuhp5tcW7WN4G3/hf/l1FlMORSd
/NCNi8YLfyIot21rh+FoKIGCbB/ltiYiHFr28SCfpSXxEC3pvi3byBbwmv8NIiHC
9OtNgvzSDUrofYMBdQEAJ8R9KS1fzSvemPeTD3JT/LAJ7aFjSuHemiOfimIRXMzN
o1HQ8mz0b76NHd6AuKgRh7Fuoxa9joCUmVcOra47EOu6YgkQVrGDPQnyayGhEsbk
K7SR5eJsPsp/OjzbQBpGgluAZ9bRccmgda6yq1Nl+mBtfWH7vxTtyRvfwP8DD5Np
mqdTc0E2rycyTE155AFZfAa3LlXWUMrNOjKA8bkT7M+jOg5gMq7ighONqbYd0P8H
cqq8pNezMkENJ1RK/6LcVjoo99KfBXGpjQORhxfXCaZZX3KxM/+TOBIA5vN7k8r1
8kE4xQLyV5ppahkN6Y2EY4XZwvMW/tr+FNrf/RfZEF5QR7qM1MkOPeaLcJsfhQRi
lBLOnkecVw1KZaBFtwleneJ/ZHVcjhyL/RNyFkOlzV0FMk4m93dcEnWEbCLcYk8Q
Ms5jcN6KBbb6PIi2yFnn6dIngTPyZQdcpDgJg3yDxLpWBiFOAeM7RxD2WShzZxfA
jLndeueRAYFRr+vmmXxQpokitpk38+IgMm1Qw+k5x5Z7PR2oSWxy2RxhdDHZN8Lb
w3O8GGLLaOf2v5SUkZvctK304ibHG9CeLhQp4jRrC1u+YJMm3MUsy+o8gvbIlcdb
GuwOKYAbdm0V2siXaX8m2RR+0bMF8bwA+QyttFmYyh63OuOTsplb0+22aUEqtmJg
lb+iV9K+R8elx2LC9e/FtekrYx49H21a54QnV5BXh+RYlo9vOwYNAAI+0Kn13A6G
9PZt+Q3PyS9G81rUuMI13FFZEhXY1hfdRm5TBfYY/MIdsiesQl0Tdnf+UGwFnN/I
NnzeXenwAecllcp/wlF6A2LvZM9KZKRVbx2gcwh+qb+VJGfwzNhEaJlrKQqjSbmZ
jm1P+djg8ZSaEjK1aUXF/6HRccejpul6fUzhmmliuHdz8ImXZ+kFsWBOWGX9P8iu
L5Ebp2sOHzmZ2CfOaVsiTZJzIkW9bhXf6owPvyIv9nfCE15mcFYbVj+Rlomvb2sh
KqdQnk2VQdHmd1s6WQbsOVzFuyQctGakYTdLDYvSfcRKh4X6sxKtVjgRHZhTniSX
Ar3vtJoAJzwJh94aPOWzVSeeWz5s7UfTLJ355swP3BhttTY0ZPmmYfkYsgiNJ9k4
YVgbbIy6IwY0qHtfj6LQYzbQM4S7ixP1Z6xBXN+tWhLgX2kYo5VdcYhM685vTmw5
W9TmNUqZ2kn8ntcXh4rDYx1gJtIvf8n1FtP3oQ1FDeJZnEU1lZgpFGkVD6XRKk0h
19mnpGFJktnic5d3HlK10L9IVjbJCryxDAhES/QuWCFPwRZLVtv4Ga/mOYmLQX4q
hAd+xe0cmqU6xQIELC53AdplmDqzaNGoqyLRxQJPAkSI3+as5Oib3h4MxHjmz81z
JP4RmTwCxqiDOGiZE9FLnZ5Kk61E8wLHvZBYLXhFalG/ZrX/xQT8lxvx+NtD0eW0
UWS61O34CFvfLuRUld0Qg4k6ns6yOauX1moegeF4ecMPrSK9FYWnOtbnVxCO5Zs0
dDbt8jOKmxtpXnZdkNZkVbLWo8X6Z7cO5TaHYXztZzW9VWDTXfzzMq1SoWma56A6
y7vNV4JkqoVVYdJB9K64ZUrQffTeJRk+sxwqV+1wD+nQEz7clr8LcUUha8+kkzWk
qwqUr1veSL+YEfNrURIubFgZGTpNZMZCSH/szEwXVxloCOWarOF3aMIagVUAfHFK
/sAbKjU4qtKl5RSGxOTBnFgrduyEWEd1b/5anWHjXjfJev8MhDwSGgM2Tjv0HmxE
wZ+ax0qVWCCErSjX+k3qFmfQIbb8M8iHLFa4zcwwfP/oH+9Ejk/FTZkfhQElh262
3Iw4xu0yEzYEw/U26jqsefbIEoaZGl0cWYsYTMd2E3ge/mkGtSL76KaiP5yJtkhS
E1rzMDdX4hGdnb8EwKF7K9ue8QWpRgyZnKmVo6yB1Oa02avlAI4X24sbfJlUqVEx
Boaspuw7haXRm+5k4FCacHEsZRYCewI5G204gRK0ALbXPFMbEVYb5s8lrOuvgRqO
NbbvkfufBSimpngQxfsRVw/zEdS7q7va1nVj2B+YQZUOFPVwMAEnT0oOYWcZVZB2
T8D6hxPmovUuY38/Cm1ItcxqbV8mxH4m1J24Uwmb9NUz1OuqIcjXRPqWueHpdfjL
JWacTu7LrAQUNRA5KQCF+o8mChoMp7N6TnKQbFccDsbib7/UpU/j9esNntYPyMjm
OeU142oekeSq8Xa1BnNxU0J/NYARKr9oDlAAn743iTdCgMJO/SsawtPBEPWGBNL1
4WCxzdJi5RKlYyZxEDTatopD6y9nGSBfa6hOpnCX50XayZrhH+0uwagDoizUEEfw
VJLzhyxJTBzRPWLlPvfum3plGXSKrjcejZj7QD+sJj1qv2M998cdAIQPNxh/Jvsg
aaRg5PHyfkNSCQv1O2RCSN2Q240BjK4JENDStXN7SqVbE4CXIZo6P/AaINllQEgi
OnFPhzQpIKm+JpniReAbDB7zNAcBDql17FL16ddbZm1HPccUMI9CN+1GTjLXcMe4
XvZQqT5jY63IpjLNIznJEXnL8lhdfbcKOamG08OYITnV6iMOqIW5sRjhXLCYr5zi
qdzUe+AYxW324V3l4N16rV8Jj3tXTP/B6FpCc4ygKjo4vhgSs3p3BoIeszosypYW
q28PLYLcDXeXqaF6Tqjw3uvtxGs1NHL/Szzv0phb03rUOaq8pQsjwlEcDnSVGtWk
wJYASpXJyKDBgeNlxdjPxor9E2yU2hcYepnfc+4PDulPAdgDmDY1PQlnvsPoXepU
s7ftaX5u01KPzsipfbNlfrGMZrQLj6yf4F7Hgqcqa6ZMOejwx2/v7FuERk/tlXs2
w291oK60bz36ZCpuION6Ww7sjmJVHg34/BRi1mYSudlabEYyCwc/q3eVTmXIPP27
sVp4v1Fv11WeeTrHe3Lh0CJzhK9srDZcRXnFIzK4hUO7f/f35XacN1fIDo48HoIv
AyMgsxzIfPjZHSkUSHYbapo/Y5mWWn2btlEJ782NyCWQYkoBrE4i4TwzErrHwTxg
0eJS8mlpsjnWewpgmlNwJ/SO3FkNgiDtWpvKzvhA/jiN5iwt6cqhq8RAuY3J8gZD
vbpKMeHHnJo5um85XQpkhdwhQ+fnIJdW3a9nYzkhWtnSc6diIp8j9IH5tOB3Lqfz
3FH4Mi/c0LHYpJ7eQF0bCLB9mTelQ4P9aQfpwdb1CAgZZOZ8y9CAVvyn49krEDDK
BcyFFNwnbReAEiLaIhLNVBOB4Hk/JVaRK1m5E5LMV5O7A797ZT//eBlsQVWnl/3h
z9+3imSD7t4n8YttXcORnAFO+hEu8NKWZLNijKcvJiuCCuB41NRv8h318WO2vcrV
9n+497kY7vmqldvu/aq0ZSYobRsSGHypOq0RhyIp4bFFiVHvOIhN8tCsxwIf0mS1
s2kWGS9T2zniDRUzz6O9rUVv9leSD1X0O1suwYRDgSwgoPPvUVpJh/eMHrZR3+5R
FzFWPud1wQP0loeZzT+HgvtcXqWPLSZz7QG+WJ6TnzB8fI4cGhQqv8QN5CI3XOOV
4fJQxn0Lv08QMMze+1UP7qsLq9fQz48zMJjQz/D4/PpMoexjzmskm8IEotkXt8ur
+CYrEJw870Gb1sSDVcWvMW83lbUau2CE0tlzudDZYWfRPcOK9EcLayvQSprUQk5n
1WowZFLMQdxZFGk9CoSLKl/xHNIJjFo3bzJKZtINiAJhiDJD/s1P7+ybjTEj8Be9
qNbZx7qzWpV3pSGKTdBa0KV7sBoJhsPqikR8ccJ31hOgD3muyc9qUwfo16j3dElq
501e5qkbxL4R1qwLDsF84vlbPLssHlbrEXCXyi3PYvZRFb9BCiVm24AnJCFBO9Fl
lpBX30vX+ofjuOZnYPwCfQvrQNeV2RBoh7nXjedEyL/CrM8dqTeZjTSzqfs5nza2
pil6BiuOW2vtzKrbvGTgAt3MSDDQV0OwmC8obcj75J8QRC4WhHEZH1ggw/qoboKD
Ua8TKIFTvPHtiiuM1L5kEpFiALWabZEr5PLcJj3zKnHgOGkBpp2jl2Tb/ShYTDCE
RGaNjkchy+qKjCKtfv64j7zZcBT3Q2Kucmkx5GUVgGdfyk3LRzXnVKGuiNAoLL5+
B3Tjm6tvMRi9SCMCCe9As63VlLglGcXgZcI0uQHQv38yg06nr0ErYLmD2htdy+f3
USBG8ZjdUVClOp7UhrcB7nvDRuoBtio+PSKy68reSFAJEEH2Z5SPcI2GEohFfRXt
Uh9ev/SAUy65Blo0lu7mnTev7cEr4r+yHKieXgwCqhenRhSlAYkbBT77qNAxCdSd
zDzPkemi2AMHT+s7f4FngtZ+VKo41BxpfEhzSLZw56CrurTXMtRIRiJ7gcbMLdK6
xbPqhl62FRApPWho2Qv8MbLLY7TdlYQyAxG2syi1eLu7Pf3sbxKLXJ5k48u7qAqS
Ca4Qnh3TnrJJ5+eZoy21IbvS3E7+8rxHxfrehT5JxUEnPnJOEwJo1d6Ix7hNKCzS
mgnzm0eWm5iY3YC+wHcIdxtcfaqMm4uJ/uY3RBmSqBkIiY7YYhCGATCM2KJkVrbu
pnYhXDM759A7tdFF/yL+8WSFokmCNk/49FevvY5c79QfWZsBl1Prgjkgj4i0ok/f
sk//JAZpM6QO88ekc2BMZQnmd8GCN40nkuCLinU5ZVmdtgPym5pDxPbJv4vGsFpe
nmi9Kt4RlGHwKFuVHgEDl1nrkHHBWfhXR/MYTnAsBlhnVJgYYzYJFD6RxohC5x4t
LBwCdzIUHtVPt0sPPkFOYeanWId7C/NWLq/fNtCLcSGdX9V5NM8Mqycopcdc/kf4
WyLOO3VtRRGIjXXnWqyIB/VSg3A4CegyvYkD1CQiml2ptwH1NICAnSBi0qNVL3at
MJ72ELshCu9Ze6Sv6O0nrN06Fo4IfLYrPxfCpF/noSb5fRmMKwB2Y2MQ+pdLmEYR
grrtj5ZfDvxOLN/VuvBffonNTznwBwm4wh1j2MyvkWtCGOhczd5ff28ztruuWHlw
xi4tpAPWzTlMs9+Cfar4CR4rFqDwMcr4qjPckd22QrZbua/BwqK5X6yf+ZF1VRzl
/4A3HjBZLSf5sqTK5tA9vGrU39tortxtRnlDOqQgwT4hR4r+8DtlIFbsrx4UA7cT
+OsJIfWh2K8Oqic6hNwgamQFIGVTgmmXnw/P9YVRbllbwkaad1opUxzc8nM5Zoyh
yE3EpTwQby+vfazM8Mr8JqPOepqKpjvHAzuA9MncYbw1LbEw5vV9YwI2Z1l7aH/m
98a55hIxTW2uVwfFFA2ZlnLZenYWYH9NNvC5D/V4Mei2d54GFPnTqTr8OLLnYVBp
8fezqGDbjHvKguGNHVuP3QonK5igHX/rFTXzNj63NaBQag1Og/yClF+QinmaPlKq
kvVceEQ3vG+UgPV1l4YqO4KVx+O4wT8/o99laiVU2Qna+VUINiaK27fgTxLmZ1sq
Xh+49pPrfkFf8E2+fd6kk/AQ1CgrrVStx60w0fj64mqUIxSMeRW5eOQNHBE6SieZ
g8ABDz4pRz790hjqamylpFoZYcYS/oyZh4aApz+AFeNISK1Xx7ZVp4/z7E+OkNGB
ZtMJcRCCkmZVNcAbDB/x6lJwbYzXJXXVsSeIInCmOVNJux+/pyhg0q9qpktAV459
1u/PfIYgleWTKbZ115NVSIvsM+Aj5sPXYTiVdkfbzAccSBCnA6a4UItwrj/7l0Aq
MIfd9AH3/84biJt43mZgdJDom4VNezgweqEk2KX5TY17th1r2CqJIc6CXz6ZZ/AG
zkEhYhgytau6chELyMdEpkPztCcJFh4oLpqJqZccN/X9UcQ+R+WcmAqMpgxTlX4J
VgIE5fyPu2snbg5kXy8i/Gjb8IALbe+ipkf6Tye6//t+Idu3252yrTAusSgPoX1V
9uy7/KQ6p75vgICG1JJ2VceAlpgwqMLguGEvcaSfJpJaG5kKB+AcBARio43ylc8S
w9UdTm4FDAF9DfqxQC33NmCjKE6iWpb2EpZY/BewWBLnmn1hGo8avNrujo7ZmXYD
XsPaizF4aJJjUtA6EF+j3SVkdZRwkTns2qPqHAKSSP0YuOjvYKBZJNFjrlTADwet
WE8ORYYUgiz9ScLQM/0uKwXI1nRtid/1KrivrY3LlFCDInEAV/KC/UAD/A/POTzI
bjNVBASL8BFIgp9PAN2Si+pygNmgsLOgsrlhRFCbJrfHr8gHtbfykr8nPWuk+YZC
+xlH9iu2Oh5ooWCywE4MZ1ul6KmY3LZOMswF5wAjH4Ruk/K7WdsgsMic3aERFam1
FILDCjc2qQ+q6DZlA7vtb+1ZhlqeYaL+MJdaNjSqnbBoSouLEpE51v2+lscW1gCb
iVHAgosZyw3KwgHqucJO2D09aywSmsOWzu7mM15paR2NR67c+bAr6FRHdkBhDGB2
WV9mZ0Q0SsYEKvsJuCq+kgAqb65NvcTxV8F+ArpUN+9OKLpVxH8baipXxADWB884
hY7MF0vmnVcE9oGzJKrtweGNSFcSBnvlL/COimwxfAg4T6/GkaCkwxYPbfizr2DP
oHCMfbLL/NF6isqgBb3Saq3T/2wRknPt8N3VxrLMyo4gaEvhdXVj6m46TtwAn1xm
hqAReVuAFEIwuXkQpuA6wMcgUfesm/uMPN6qgC2ojvvsG4XDbmU76QIyhxLlLAvV
6qasynr3gaT7RIJdo0IVj7JZMzbAyFhUScUKIK1nm1FVZ6h/Jq76LdMHNxzxzC5Y
bvoXhsnHCdBYOSXH7JXue54KqmtG9BXoULKDFI1mRg1NhzdEwQn5pN0MKPBBQlOC
eMLgGmiVrlKx5hlCVe3W8IG0aIU1/4e2QYjJ8OnxqH3te9sFRJYwpJZSQ+fqFGkM
H5jjz7jAPJV+L7vm9IHC5Vz1lmi1peXRpUbqHj0oB/NqY+g7LSW2TrhnZe96af1L
mwgJM2A/KuC3fY/1NWqtt8wTlS1vVl3NsuhZI9flBo65zISvJ4osOZiqlkt3g0ad
Us5SDGYTlXpcP8kncrtUpqpvL3H7hcbLicpiPUklmvWfCcN3k04q6LSNF9NoSi0W
NB4AvcU+AX3weZJM8eRD+ctgALUcZUgx8L70ySumAq8XThLG9aDgvQYMGWqEycHO
ugynjEzZU3tpuVXC+/zQAHJkBth2Ez6Y3nOWRVUpYXzNwbqbjO6GTpYEpX9/XL0d
YwTB7sjnBwYo79h/hzfmMzFiOPTnbA1BwQCZ/O6j8x8DECX16C6bhjid5WwIwmZl
wmTFUk/Mk7FGWtp+TnTyNMm4TnW6iPIPKTluNmhCiWlCN3682HomOLHKQ2Y/Yf1l
YRgR6vURwBTbMhxm0xaFo91gZ23XMXwQv555XelBEg5LQBbJZC9qtTthMZ7ARrH1
b7lFZasHHnDei+P8GGyeaaAcj+GrK5H7w+As/lgFV2QnCm8YGG2A1JqZY8VuaI4N
SZy9IatCdhbcVYD+bqHxMAFsNk5aGHjpHzearbNdY7izvboEhoyTCz0XLfgPRtoD
Q1oHuXAsjQQ0awNVO62NEcBuf88Ia+r29eXEqr0nk3S5tjvht61++Zdtqo1+351S
UMNbUnO86wO5FM9eLqwIxXTrhmYIhPkxbTgJVE+cY9u2ApLM2My0hPBTAxVkzdRq
1eNIwLjC/Icy3A01m0rB+QocHGLaIo4nFeuR3ffnilIzqDfSjZjGgbQ6eyq3IIlj
w9rJ0Gxy9jVf28TQZywqW/HubeoGPup9JOWB3ErBZ7SFYPTWf//9Yd4LRHcoRsQv
P0RFTzT4xiXZN+5D5+THh2Clxn/wW7JwF107d4mMzEGwP7+aGhys1CWi9YnkH1JD
zDY8L/srjTkgbV8tfaBhmvS/l0ncLkKqireySTxg1tpghYZrBa4KWjW0QqmiI0Su
JbnovhcLazUfKmq0f/4eM3nR+5XZdiyBQa/YdhNVTXGhJtDmTQtDmcIcanijfM9D
LoTQo+HTot6ChCKLrvGa5HXYbtZeqPYx36ASJlCOHvHjsPcJjxWntOcEMNx2WzEY
9CnjVhOiabAbJUsOeogX/Kx4q4DGU2yGCR0LBpUBdwUvvy5X3vERJvdeE8/dycaJ
+fKVlTWwyMvpCrDYYg+HQ+cb6vPdSw8NqTi5XB6eNNgR4U6FrNzvpZ37BaQhbf1J
Kz/Tt9ZEPj0RA2/jxKzdYyfKq+8Ldr3InL2ay8fvqkwLI9TswjH9wMl+x314mybC
Mhe8agH7qbFFoiUPLAtr+44O4+HPCx66WmxvDc0EI+Lt+POi5Rro9taVFfycMUe+
wfXp2P/e1cL/mWL44yfnKnH/XFTHG6w04Xae1Sfq2UKUgO/FckgmRcAf5A8G+ttA
gP+zfP0T7DKNPQaFK0fCeEARqpR2zd0fOgcLzhcKAMYpkB3boiNFkwB3fTq38efC
PdlzIpL1/LK07rOt3utxcJsp1VVNLpN6ZNjmtVAkEm1CG2xJRVcTTTiNrFKbOxVQ
dEHwDCD2rkSv0Wp3/ZC6D2RLdWASeE3vfU6AyGqEF3bLYPEnRokT1DBR9UYX/cN9
pdrqx5WyfBgQBSglDAyzOC3W8Zs+zTAc1H1TWpOJMTlKRZZ2PHFAXQLkp2zO4Tl/
2psmMDC3A/84OMUag8Q1RNZlcOkA8gDnprmcHGVHhNnK4gqqY1rVJDKlMHGpl+gj
Ov+p2C2pMGhAHhduIjREsU8cfkOjIPgilt8rInxD6JabFm/FV8nXJz3VbL4+yy0V
9+3jy3bVM3SL5E1r6QWpG599j0Ux/5XEEO6DMknAFMaeczhb2KSGfwW4eY24sIUT
fBVnor4+ugdlNCyOQBglNxckBAwlMDW6jwEEmKfITfshjZoJYM17tqBis2UP3Ow6
D9kiPrPLo4VhS4REop2+oPzjmaywE5NQfjlxYPCwVjFxQKJK7vFjqwyLkGH65LDt
cdfAf/iifP/MtINeaf96i/HBmT+KykSVQhHhYZTlstbZY/lA0Avo2hAwIwcQObrs
f4uL0kph+55bA7LsTkESk7S6th17TMxHKgC+nOxpSb5+071id4EzPUacKJJGNy+7
meg8jAdfdcc1zYmf85eC59eAj6Yqk36U70pWttIirpPv3hw1Eh+U1TOGPJoVb6/e
mU0q5ckCOy1HcTnwBbvaMM6wwE4jV2poYOFpj1lwVm+XJ9VKS+8f/f+QNg7b69HC
1R/rLZfQyxBlQQ09vIpmB4cUEYV7WtpMiuvsQeUnrvCJITBwLuIcOFzuY7G16Bdo
0mFCyI4XpJSYIpPXa2btik9mzAOAJhsZf+LL0u+RGamGU8xSFQe5HkspsHOjF27L
bESu1NZFMQmiJXsYUfTDDOb8PGHrltTArMXY9PmSeBDHBoJvcjnRufvWlZy5ge1Y
NGGpxbVkapNONz6ibebj2JWh8vrvr1WNsmqinCnMOHACuzRojcQFU4g+1OWqs8SM
KlLPgt+KwpKft82npZfyIJD2UkvswEh0u5bW0k9hgVYJ+i1+qcNMfeyCKapSVe5X
Kc4WiMmv0wPmVYkwuVMPMk53yJjZU1/SYdVF8e3DFsH1j3QSLCyNR6Z7g7uuoonb
W0j0YRw3RrWjZmx8FuLIdnoKSPGo6qhrOZ1EmfTAC8R8CuiFuJhzkfr15YVBoxQ0
g6H/YcKakDvAlgAW0lGMNU8jUzekKshcbxJAKmLy8Rz/5w12E2En2VBTLspbJ1sX
11lVIB4TNEGAei/nq2aVdyg08ey61+iAGR9gr1OKJdN7J/VHonFBj1etM80nzdnn
LnHX23+0ipAU4HsOuXeYMqY1YhnHFO3gpasyQrZtGmLXHXCPC5Drt25b32seMDTl
NdwzJ/90bvHR+x+5NGj4uwSTbR0VKLS5IekV+FlJxB5ujR4tCzVLR4fUO9nWP+40
OrHRS7S2JgjJcU38puhBB7YQ2N0QG6YVMtvEymOjV6DYK7C327vKoHhyJWaYXX3v
ygzYyCbg8nKC6x3tw1JGriB0tIAmkR3KVN2dHob+spzKtRSd0JojsVO47XMlE6nu
cVI7d2LSMjMe5Jy8bMN/CR4nioWOI1xREkUz+rVFixFphk3maawF0ccNpFGXk7PE
yOVgMUdY1AvGlmv9RXiVpFy6wacngPc1Iay6PHHY1Jist6j9TPpQTk7G4puV7DMp
+EQFoPa1vhNNsrjCjUUv4Ivn+ApnXMGkLEp4Fn1pRWgs8ZtDRLEnbT3FA0hqxVnr
dkA5j0KG+llWJu0xBmfbrDz94ImOxw/plghtBOKFFyHgwYX/cn/J9AOqGl3awb1I
MNJQB9zlVwn3V/VFsBmD6Ads7+8VK1LEJaHfR4I5SVuizFGn0sUaSXc0nlQA7u6Z
4bbFBuanI6gkg+X8cABDJZGAdkZqVz28VDNFX85OKfX5p5Q69DNAR6mYDf2ecobb
f+tCurJs1A74aTCZ4H994QXcBkj8m02YHr1OALoOUFUOqocFV9TG5hGxChrHAaXZ
jNZqa0tLyBKWfp/ctRJj5/3YUW0qETVJQSVn267mMW/FkVnOrLJj6PZ9H3f84n7B
+3s17VrUKLpOBAHFRBzF6C73sjdmUyX+GGdiavBZ4oyod78pq7zaknjRseFvm2+k
mLkH9UjKRUg9aL55x8NuHNri0ngyKTDsloXdWoYKTHOvTNrnm9XXfXeQtBvMhkUe
5hlI0l+0QOtvqayIbXC6h9pPnCzgqcUz0ZKP0Rxv8ogR6aQJJN9FcwuymMdnaE3P
Nuang1kOeA8wVvZW/o57gtNPjzKrVJL73r2SDrtp/mgLkWDYnvAZeI6lrF8r8JaB
EPprf6quQPaSEjxwYqEJ8HaYldv4TlEcF85lsC3C5CPS9WBppouhZd2e8RyGNfYK
ki7+8jOGmCqEV+SNWd5M8/w872gkrt7a60rXSS8jr5RYrUQR/Hw+2j1TGNl39OvW
S7bYz38rck4vu6EZ7cg2W5Nb3L3sWh8/8dW7ZNDuhwRkzZqfv48sUbeydhJocAVL
wNir8e867gr7TQ5HjqlzKgHgNLmS3bZAg6qnaFLa54ydCPHmG6YZ8CSFUlL+dtbv
636CHPVCQcBlU+BN3USobhiL/WRGUF35oLVRB29WttBSRJS+uFQz4ARv7cvmsuak
FBNr+UcsCe7Fc1MvrqTfdQLRd9alZy5lfHvi6un6RdbuBkKiRvTCdN/xf8LYZMsG
2C0Ss/GXOdeG0Z/SblbdTx9ZKmAHztannACFCvCWrmwfxxEhqMJ4jDu6ATZhFWQF
m7qyVf7ynVudJOqDlNQVPIYmLEQxnjEskCerHAr/zATvYxQm9AC1NA6gDxqMH+2g
6osLzhyhDHNl+ZU2ha7N8IDf+4vVyPFRAefnNr0vUmK7h2Lj4YxFokQmW9k1OLxr
q3mcWxO3D5d6ZmbD16O4QdiEKYrk8QutbNsgMsyOnlo+WZSZOmE3gpsb/Nvfkpy3
Gs00HxeQLOlJJqaGJzPZK3R/ceL0VAe983FXg+89XTFzqaEhk0AfskW4pMGKvcqH
F7nsbR18bojGgZsiDs0G9NAe7m7FcwXLZRvgryFqWIHjxAH0sGCpuZfGi6IzNvXy
/NA2PLXjgo8r4Y2bRK21ttIuImxxLBilRJSsXHKP6M2WDc7lTtYBVIbpejhiqPxa
nTZhQm+p64q3X7Q5KuyjBPOJBjLuhFrjhybeE4uDtGC+eDGUh1qTUoTOzjPiL4S6
BVq01VuXYdv8mjx7qHCeoxx5XCiJKGRH/kzfj4s9ZFSKmRfAi63lCGI9tNceuz31
eK9WpKyHVu37Knvt+3xWGAZZmz8S8jkTcsUFi6GSPaBYlmpVUJ4l6hyTMWjw+X28
jKxxFtJtbBw2WLuB9+oYzBCvu7OgBzsMI0xoDquLFLBedcfftT65j6Pesw9x6Nwl
km2RREK2wSVIBcNF13qT8Kf22ulYmJlbXTx7VZ1DFzcisXlYYgyi45JEX7PqIb6Z
PUzGxMzszx+xnXDtbuK65PGbaajWc3UEcsbEObI3xyOBZ4uQVuPF8gquamK5s2dq
OtJTXkvOUkWcziCfmJTDMhe7t0qfcUaKmP676iXDg70PNhebBgtM/9V9f8ABwhVy
PIo9JeViP6HcLVbICHNrJf+Bwuz931HT+94DTAy77dCm+Aj3bTLSVV5qFCS2RUR5
0XVY04EojjfLSSctFzjOaC8NyRMmujoE8meHTKOigQ19CaBlDnXIixl69bBhh5UZ
Spm5r+fcSipROP14d4wUZdt3TVVz64dfCnTgrAla9KQG+NlIECTsaRbXEZyOqbzd
2ZMwy2pnpFYqOdbGgJudXh87Su2MeVverODxm9k8jZIqmysY1POb5VJcHhFCpTbT
ggRNWyIKG0lLa0nCgOKheN/WyHIxJMhA8BVGR+7c7MYrnwR4/oKZcsQm7hKnGcGh
jGB2FhxZRhkvjabtDYCo8bsQ0aL6vhAOSfLVJdz/hy2NKegyddMg9KoMsyegE6RH
99dxObB2m8UOYhvSYrq5Szma5MTZkEKCdJHwXd4Lcd8EvoSgnhKQm1DWcD7cObMj
3dgQj21HeH3XTmoug2pOVeJxHf3p4Q5UfGS0BUWjxmhZzb9UuOpEGeGJO2i7Pgfp
YGL3k6fTlSdCQxpK5zls+rxoJOwdspwpbHuFar5YfRNfeCQ5M17M9c9UDWE1I0I4
pL1j0YxpC1to+ZDus6scUM6a+RBEsJY9R4ZnZORttYPsKUb1kanxNcaLfLE89eGK
TwmZcbV+yfA8PJBiUfk3zwdjQSL1MDLWRUfiFrJ/D3mf4uMXokGmHm8U3bKLt1w3
gezSYAOZnCPd739YWUQucH7G1XdUJDPslSrfAYmGdAhYs5FxrbxSwHwOKx1EWbNc
7Qgm52wN0QjINDe4C+RryoFoplKUIDkIPeaAokpK/ZaXMWyPLgDPuSRssxeP/poh
QFjgqreqrxYA6UBEOoTRwhXHS9uHg6lFKZpFYJ2MrrlLclF3fxx1qIg8MpuPmN3B
kMiMLjkvqLYdbYlOwcUdZSuAQOd/gp2W2mT7SXtbfzucuOsW+RSABdBdWKaHyuQc
XnH1DkLENLrL+HT5OTo6N3nsY/jEfBXUp8Az74FeDEPPFzu4B/8t752yPryBn3vt
j3AvtVgtEm/HIrgYoFLzqTFUyMESyvF0btlx6GCi/7+u1wBaKPp5MhohhO0/+UoI
NmdnQPhdAFkVQb3uTReCMmlak2INcOxWQVST1rarMn5mLTPrRf03KSOu6U5Pi6cd
RHDNf+DzaPY3EVvfR/Jf4Rmx20q+GpuZb5Y1TtV+6O8tmKkvdwufi1cVSQbpeDuZ
bHXH1GhILWLk+xmQ2gHv08s0I3LND0rbLTS5a2ZkqpGUDrTS0yQlgZtVAIjMRO//
1ynubymAW+aonaGv6UHKpcrJNq+nZgDTrZCrcVHuVfr1f6xWdFntEVjkd2pI38Lq
OvsbBDd1Neconrn6Gd+A/sl6ytNuUpBhGT9HPsf6Fd/OLm8cRTTNjIkkiqS8Moyx
XXjrkcNqSocJIRgXgUWh9qTQpMaOZXse/N6lSXmzLo4iAHQsbOCFBxhkgPaISVLn
pntXUB8W3AbowRPCCO8WFVWgbQ5Y7ixmbYap77FyFEAv3HUkvp774D8sWSBA6csY
VONxD5udbGplV0SXwTcP4Bv/gC43oPDDrX7pfcnbeC908P4lNDKT0K06xRboO3gO
VtUQKlfZSp9/Q6hQlarYjM12QOI09YsCh9X3S997rlvy+zoYhMTB707CTlHrivy1
FLx9cJWDratKx69eb/90LzO73s8pBCwgwHce5poX9Sr89Ml6b8mLIpWdBx3kBlx2
cqKjcly6a4mtxxXHNbaGWwWcagyFd058wmsOcZNll0GwLd/xrc75SfsXhhx0e4Yc
PO80bo29RsAg1UBdY1qBz4yd8HgGUf2UNOVVvLQbngDXel16AzFw/A3ZbB+qQHwF
RFgGxD5FFZmEf/X0QEpwrOWJsMGZwZUeh4dco1RUugR/4ff8iqAE8opRqdm4xqSQ
6JRC3SwA1IAGk9vLm1Y2i4XxC7xzzTJDI21V/eCKzq6KbWqnUyAQHnF6BibCa4Mt
i9xA3ZF7p7/INk1U4B0oQ2+LAK+sodaRqn50CbdspKR1WsSLxjUQtc21e4Fn2n3g
cqStK9Ap5BfWSYg0iwXk/CZANYUr4i75dpSG4BOTJOdBdI9AL3dhHJIhbx/Uyl8j
267nxN9Ly1MfIfT4r9maEifdhmLc98ZMrPwNEgvXQwS4AeK+risUNcUrlmW3Q9b5
m2ad+pVwNRwX9PY/w7RJM5rmEz2I/MGxIAXTJHZarzKiq78KoLWzpXtWQTwq/yMN
/9CpaKi2UsHVbC5C6loAfhaxnpFbRMGpJPisdVreRYN3GU2qIz72CbdNHP192pQ0
vhxu84NKRtoydXIwPBExnB+f1GN0HxGxIG22vP+e6PC1JfE8St4PgUdgOLyAu9Md
Om3MM8sohw+lpjVLDw3EBM+r1DwXYsdw4I4L2axzHFFzwxaNw5GyfD0l2pfKlaoW
ntQvSr582VwY4oNjakfxlJ8PB7dZbmoSpqHb4kxGRgLCNAyO8WpCSWzLtRtkZEk5
0VseFHw908AfeYST3wqnKBkWPukvVYDQprfeddpm968w0wiY0IbVEBeVwKKTOB+c
wfUo9vPaIH77C3HNTTY9EAlyZAf5aeJldYAhqOhYapCzYZjvFPKVT6DfbxGcgqT6
XLY/+L2kPU7Qospw/OjSOGTS8siaaNmleRmbxg4zmQTxl6HU9HpghQLzsYI7TZjq
Bfh7wWf1+px5sNjLWmz7KzUDsINLuFtV5+VF3SnSPYdCKQq/gx7Ujp0ayTuyTthe
qzLaKCHQ4VEhIfBnZIvp3IOwRIiLyd0asiSJGf8ElX6CfWTuePgTGodvrG7Sgvtz
R7xG+7fuEYlQBu1Xxa7Swc2Lb2jkFsKI/y57hOA//iP6wwww+zc52vHupLG3eFEW
KaqXPBfia5O/lx9Tf2T7/WsK8aVkl+kogUZWYm7QpauVwY8EP3q3OPExpPUxYneV
k7jGXLH5CF9FhvRL2TR6vCKI1uPJv7Lt58IAaNukXIPK0G/cC2E+2Vo0CfMppvSP
EHkf0wqNoaGbqK527mM5udiesl8x/aTSY8TXJ156esVXpAX97Jmaf/4BWJ+UXh/T
/s5dXRqtckSHwwpz8zaH03jSqwSkd/8eV8ZYUFAVWO8kcH+ofA/ejPEN9vVpc/o0
WxxAXGXLce3GTkjat3+YezqXqrmAh75LaJmhkntihXx3zswh+bqw7VcsUtMGHrAP
vJvGVI3sddq+HEL9IqYNQLael3jZ689MJ/VkqgybXyktvUEeeBOUmBvG0PxVZhy0
zfWhoDCyOvQJQOvEggbbxkL0lUg35/bAt5rPO63bhljviGMlyZ2y0SUcZLAHox6k
qHS3jP44mgjTUKng1NuPVgYMbqpQF5d9NB482wBWlx4ulHjd9n9GEjP/7oJ/FcEG
9AN/PJT71T3N0eUSVXPLaaxlNif1maBs3MtthV4PVuSJPPj5OtZTbGFi+KPVAPpn
fLtU4zTrqaT9zTVccV/iDts0uDxbq9SEp0fV7h8t3SDhyxcLV4vbRhHKmfmzTXql
aP/5KbwJS56rnM4ZTfoQFWWklFapXZu7kR64a7TXa7apn6ffunR3Y6EXRFbQh3bp
/jrmglrRLHbHQn0mLBVv42xtvjH4mBhnbaAj78Y8ZW7H5yDnX/l3jwztWKiys+aE
v5jH6zQ8tBAOVLP9YGyEUuqLAHw59Gaa8uVKsduy7m7FIRp0P8DtvYHI1OMIvY+c
37ix6HN+JVRgpt9hPlMfkN4bc4I/2bhhdDQ7xyZ1nKELc4WxhNzEKZV0nyL+GNLN
VLaH5CNFChItJtVhEhHSu/lVQ6tFGGQ616+xRPDK4TyiYXD/+dX1CBx3d+N9IGZI
jbB/QMgMLRK/d9jynpd3obQlQTynDiYtyUiuMJTRy9kNj+W5xJpMRawIrGFGy+9k
XFSnpDlKf2pwi9aL98gZj3mWmaX97Z4Zqn+ybV4UEgaaIhEEQ+3Brd2JejXhMn2g
+qjsLi3cVuAl2LUMDxYfa1M233+9qgP1tKEAaXMU0flcWnxcUTBL2C4hMRzNNHWx
YYADsf/40qsB6Mar7LDVY2PHxUMZL5+p8ZcfHoiA1d7GMkb4/6LGC/kpMH+kXdWv
NVZwPbCEVEffRr/kvMEXfl+sk9vdTUdBX1i7YQB79J88bnQWGLv4lUoU/rIwyhc/
ypXe0qMiPXKoAiip7Ii7lNz2LmijIb3fDnuOKwfmDD3BDhtxHKvgmDBiGvw1Zgj1
0nXJK4unE3wNIq5z+E5dVLMyY1839pYPxVTa00PyI9TyJ0M2Ucte3cck46RA5eDz
dmkmRMHiJRS17Nx8Oyh6nXE5GfvqxJ+j6L7ko15WnBfUeZnq3U25mywnTkPBpyfw
GAkPMqpEUCqL8eyCIQizWb/bvv3aZ7lETd3gaRKin8/VJFWHAPfooBvcoArvyCBb
k36EqBvNOFOw7kzFJcKJZC69DivumTfqJtZ0cOT0JbhQ1jIwJCGoYAtnbiNjGwCl
5qpXjbWraGhk87IvRH6jjZmbKJP54w47TqP2jRhrA3TfTetGrsE8A1qn1Hv8BXZ1
w5Jx7XCodXeEb2xZyWPABoJ2vKZMwr5NnIBbUgSwhASXKsz90wCvWQAMS7iE4GCN
9/61EuwUR3TwiObwR81T8QvaehVxPuUcBaIqrXVzUbAbKu5QWcnJZC/jsfmfWynp
jfRvwiQGCfOCtqnb1Wspw+w7U696ixlbpkPZhxl81M0AA+TBmdgeyDpj7NvL5CaR
JBNNqhudKwElYgQ2Aa/mLud7XIbYKPvQx+TL5KJWPS5ISAzXn3DjZUM/MTW4ECoj
yo/+p2+h9h6Vjhug9Xmb85YJG3u6saNj3NF2FnGAEKb45MFRThqF6QKWglrl1Jkh
BShDNipBSLZqxUc+01Roia4oNk8yHpKlrMP27brjj28xKpyEw+kgbSMPcuyqSPH3
YmYZhUSo/qcMtvQZeqpQbRw7yOpQV/nzYMsgyEGY0lmTYLNEeUHOrcLb/cHhA9yc
v0CUSs3ND2RBs8k89KP2B0EDMsQ2QKk5WFvO0gJrlP1i0db4zsZEtgvWTRqUxldA
ZjjWurLGYyl8s0neYMXywoUHu8GgN7aPuF3YEWQj2p1dNANqauyj7Qs+3WFK37ws
a1jN48RfPYdFngv31c+gu3E/13HPMtjluUx1a6webBjm87BB3fxWHl69AzrNcpP4
/CIRyC4SFCyO4c7Liwr/CpKandu8dgJYiBtoarH0LRHAcQyxlNtDDuyDXj5XZaSp
ef5J4Ou0kdq8PSiplwhg4TwHiHpb8jGtA8RESg1TteEMM3oeNATfI3sFEBWLhiQe
td1vxwkJGlxXai/DYqZzcyFcx+JBCX55K3EqU+8nAUX0SNRLWu/ZWx2sEVh5Geov
TszzF5E5bax48gY+Es108aX7qZnF1sIKLHxyXXPIStivlOsGMcdG9CRbhC8Z9a15
6PI/vEg0fhb3gDUqfFcqkxIjwtVU4w/8DQtL01dpuoUzTcogBFs27e9Ax22GCe5m
bmcYMTTIefDI0x6bbBRbAH2uh3W+fm01+ELNVsKaRVnLttJCpV1MRObfmnumtWVy
k+5Q59g/V44u2AtQLV6cD6w2kfjBK+bRcUiZli2GIyTz5rVJL7loCA09VXh7YUl7
9giyd9LRis609BVeR0GoShBLYeWfCobxo6poi3qekSzmT2FBRbhn7PmcnogK0kU2
PGmNfu4M4XRTRq8NjgIVHf1f3kYBdmbsgKDdvVULy5zzYCH9Z5kXXtCV+dybdFE7
uNhpN+/B/NBpp358H7BsRo49r7wyAYe8QmEEikfiIijexW393NcXaoqe5RbMbiW1
AObFjBljd7c/6Aqn2TCTviXIGa+NoRwC24S3coltK1E+lQ5MTHch0IOKEcPlDmrC
QfizctfGl+CmQT5YUTL4nx7fcvd1oRMp69o3Z8fkrnyamAjAkocQYV5JWnp+NtCw
4t/KQym4IeM8l30P81hlEFd+Np+42wL53dRK+U8QJvgELOPDvfVmBqytF/h3oCMW
oOxYKLTYPaLUWDOepBHDfLU1vUFoC7BocuyKVWDnycznTsAKO9yaUKlfKioyf8AU
OG/TLi2976VyjwTZsd8XCYJsLuNE1RYdCJojIroH100U5nTGcpUqe2aCiaYLRq42
vU/mMZD5OMy2fIy8T0/EXBXkGlV4M+68/EylwyBIK21FYMG6RTZXVnztAJZ0if91
6p9KZK4VvCRFQGujK/aFkhDbT1rq1bYSzNWZyOEwi/5w+26vsn51xknsywnxP8/K
efUGXc2nN2MDaskLnIp5jgtEVF7/CAgGWmedxg4Gs60GrpQMSPY7ljVJz/742PVY
li06fZXU9/h9L2EbALMmJJtX+e8prbZIhyduhmY9qMttbzC9q7sxGlBtAQFzUA3C
+dDqfoVfwh9PASbd5bTt64vH3Xv3w3CRf/L4/knFqEyM/wbxDCzVOHb8GLr5H5Zc
hO8Av4Ydt8TPYCZuPYhDZNbkNYwbNte7x4jJXmk7AduNVw3Vwu+aZvM230x20m0f
Rkrpa7eV4AOupXXkBC3xtEMPjQoIerstlm28kbe0UM1BM3VugJkUWdzenyhao/iU
CrOPHcXgpFpsJUQ/xrFPePzLcNBu5O2NIEayuTQQhCu9EElE3rcEOhNpy8DMtHO6
c24pzl1ugm6kBjq7r6ORWM4YJCE7M73U06mSjtArLyKIEMD/GbwYXYRiCtkFduWM
wLeLGatEjsQr3OJNoUZQqD1sJGO1Ji9esMGmG5gVX27fZ7h0ehnA1YzpWRSDrj5E
`protect END_PROTECTED
