`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gfRuuxM9flUUTBIPwVEW5Iy7/MEU0Ps712naHXsf3WMQDi6VBWNco14TR4wybH/t
KRsSyUv7iTNgrCSYQfrAfQOXxRQ1lZ/dL53P2bA6cMh+v1SRrhNmQcMgr5fPuZrZ
Dl3K5JyDp2A428AcpCfmWW7vJDk4duahtVJTgnIvpKiZ4Tuht65LQUAcXSSuQaTk
j8dZRm5KEcN6FMp2Utgpo2HOaPFZcV4TRB8goWVkY9VIFmE2Zqz0/qInTQqhVS53
+0/zEyBF44yqD2cw1VMmvYBVTj4huKTAzp0uda9ifh6KRUNUOyIxiQaUdvKzEws1
0wAJCsmCOCWmClGGtJYXqktsvTV/j0evLLRoGssFs/8W6CStqGHbKHMS9oOTeEpr
0LvBvl+E87JK9wUE1xR5i3PwQcRkiwt8ravuSKUxKnEc6wTwUNSkzorp3yxLl1X0
WB2o4Hc+hZv/GaWnQhb/MNcTWEl0Xdr1ifjbRMhltisL2ivaot2J+6eH0T0YsCG4
Gwwg6aiR3ARknKktg01Dc6u4efxEbwwYqor/0KRrjJu+WCtJJyfw5L2B79+GQGUI
wa2kVELlZsD/W3xN7DQJPhQ+xkAvxCvMPq1Bl/O2XRkc/VBdFmWtGkGJi2vqoDiT
L33UvrKKns392UttdUAiYlE4LkCoCapXBttknOOvvKb0Eqk22xq2ez3ip39VtT/J
`protect END_PROTECTED
