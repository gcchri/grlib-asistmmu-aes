`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Am+3bx4n1vER1QqBXPXdxm5f6jBY5HebxOUvWW2s9pbl/cRR9Fn9D8PW9+TdNCSo
dHe+UTXCvKKHMQpdLdBpSz2DsZUhl23njXI/LILfC2v5nEt3RtCTN0G7PIGOlYht
reP9ZCSLe8AEZRb84HVtvW10coZTzP/ZROH7C4StBe57UtEpchtUjAaRwGnYHbZ1
oZT2yZisa2OOVt7cSIpE37i2efLQ3+5gd+CDhn+y5dA2mILJeDuZ19VJHZj16XuL
h2GSZghpfcSTlqdt0aJFjTbwdXpJvV7yAeRlCkjiwHJl9krAS84/1P7FBH6aLRrv
733sWPFsaBnfAzYNE5WGdCqXvs8Ji3EFl4F3PMncvGPrzbUToLwRyfuDiUqXqqFs
jOsXcbwb0fguZCWaopVTyUCp8bfsdHAdxlH+OD7vzuF+G/JCZ4PWbUTgg6Rx2zVN
13hfH1Ke3pVuvYgOOGYwnm85rn9Ol0Var519IcLtpb1RLcplYmGktjxUTFwEojqY
UeoRa7oOhhSIm1N19g+ZOgFj5ZKQk29II6Ku8bx5wLrzH4JjgSjRE3QpO1TZIVLk
Eqrnjc7EJDIFZchLVmOjxqLLXVfmgMTAeYV+nFbLy4tYSoGG5VPYJU4tg8GWm58R
ZrYZRPl3nbh2kVvuu7L7lC9SkYkOIbLtgq4zKBYvOl4tmyDK6VeIBuGhwdd64JoG
Tpw9EPO3pdNbXzBGA/8xpVtY/SzTq+ENucDNzKe1TpIh6mI7wac8UwfdJMPv1sX1
11YBHxToGFJhq7nio8TsvkcBPC7zIqjov4evHbzt0slz5cur3+ZKz2vnO9hH3tP3
9QaaslFqR3j7hRpANG5iV510jnD4/i3pCf4o3j08bu13HbMTZRDU5zCTlCLR0+BT
ViJFOx3ByBC8JBABs6xE7nuqZzIZ9xRUWRjX9N4yIKJNUGUAlyoC1bMJL+atdmMD
7Fwkma4VGwbget4Vi1MHCg8azDbANO/wA1X4EGacIVpVoqsnsLoMzJ2tokRIxZRU
LHLgsgedZm3GW11+lLpzBkMfcgW1AAn/atdNrdRujbrBJ+5juIwJ7a9BwqIlSSmK
uWPpDFGM7flj1A5OwqwERB1JLVEqFGgw5WGqBL8YsXe0U5NIEX8erX6yaHAm41W3
KsFVKTdfEEx5RaZK03+tAFJP+cd8kEbUlTMhUEmZxsR1CS9yHvn2fOM8BGgt33Bp
wtQxW33M2kMXc8V5+FxnCQIuVYjxC/GJR3th3oRWvj5ZRxgtQGnV0QGpra8Be5iE
R8iHv7EpnpO+UOWF21gVflQT+kqKO149fCHpwObrse0gwG9xm3Of0huPiXgcYySP
WZO3QXcYtXy8KCE+d0NLEfvuscD9aSQu7ee+77KP7OMCDpXk1X8SBiqhIBN7yCOH
F0W9IAvCLV6C8DDANOcuaVSNW5KmeeB1vdYBH/cbIgHXIbX/Glb0uR6nb/QBVIQr
Zpve0AcYc4dWLNfvyR0+/w4Dx5YSZA3fE/T7Mk1VIvjx+bYZlBHHwV3fI9FBYGiX
MckEwLlM8+s4qn9JSt0p2n0SDufrSXI1Ygmi7qYHugAegv6GZO1iMfL+s1CKk/S0
7XJD6dl5jxzNDaSpLKygxLcDKR9wn9jBaONkXLX6yzJsqzYuIn7GihYIwdgh2mlL
2JGkXTFseQeLaijhKFtJMM/wiXhfEGeAKslJ8WPVdJpCHqZXn5UtYKFYEw1rWGLH
VD2zcP3dHKsEQjfKz4ASptYabJVy7EyM7L2hc30kSqYTKl9lD2bHcRS9LTK1PHFq
CYO1pqT9rowCYSqr0PQ6V1yv5BoydewFpy8zXl6vb1alc3tjIK9gSbv+MeCvVU+E
nmugrVTJ0FsAlR15WzLjon3KKqgSdCgg+UkDDokoB6hw5n3bD7r2VrBTnwf8u12O
qRZMCoct5bx8N7qS1gjksaJIUQyRFNIPDPJuha9DRodtdYeRT5sSNdT5Ya5uXq9k
IPw+n9R/NZBP5OXFHw1xfmMpFNjDoFTngHi7XvBLY1OLkL4kPhd4Ammf7K8dFOfW
1HBkglbwYEnoruvMZ9oyr01oSE9mbU7so22H4qWVvfg84QFlrIj5IxUuHL+TX8qw
hCwQSVcbNOrbbgR9/ZV2i7PClgXM1I8/qw8d5NbUAtdC3IjF4S+UI3sYSZHWLZlY
IG4NO9nwS8KRP+N0/lsj75Wd776kYxzIgipcTnrC66diCDeApSO08Z1KrZB84l9H
o05ZgZyn37PvzAUcYe1aFVTlDSGsrksd2DPVR9NVBnyWdai0P9nxp3jvFvb79T2T
61mhvT5UhEn0eFH6uAthta0fZG3+TdWmNsYqST2Q6Tk9vsBe4ryDHQppe1meIYOY
hZJM4mlSTYneEE8AkKqbKtjKBpqPk2bkwNMCmJEjZgpGZrnONSVExEmFJFQ166Fs
qlO0aX+aFiFjvW6itIZGYUyJn1vTCwaaA7gmSkcotkFzmWkdyx2eKceDbSgR2qhB
IziWww08Jkc+oqLJ4/lG1V4DW5WwgD8Lj4rIZdWv8/6vjE5pm7yGYX8Z+U2mrT8q
uL4p9zub4GgQlYi8r0WAjZTYJiXoqAy7AUuRqafy9ne/eBRAeVHpc6zCKlRqq6a+
wFaQeYr6tRA/lW6i2k/yDvwKXActVJQiuqqoBGjSh8G796IYJTI73EZ5+2PXg3FB
YRSId1QimF2zh5ZeJZsJzWO+yf3qnGppwX+8+INc5EE5z8w0gDoUkGjFeQtKT1wI
L0qNCwM00UHsBOpmFYwwDgML7M47/HO1z4xO5bT8S5ramertM/d3pdGTczE0ZFBQ
FcPv/8/bPxT8+64+cRkNCfrJzGEi7AsFfcO6KxykRTdmH4oyVl1d4GZQVKr776os
cmB89gosN/l1vzfuHEu4iwR1Wl0sog4WWcpfxDjdYkG2AvlO5KOK6mWcncYChgt9
UhqsWKV/pXentjIvv8ODTg67JXXWPD5Rrx/WHYi7zodKpYnpBa+8oE+BKFubs96+
o3i8OsjHh+B91fie1eYSx8i0pVKAEgvTISfzK2V5w8B0eeCzv5pAW4rR9YeJFDd3
b6DE4rkWbiefdwKsHQY8indM/sx1A/5b6GXsfgxLFxRsFcIQA7/gmrPiyEQU3D2W
8ooS/ggPmag4PZiA/qruncZcBdXiKBonHgZyQbBc0BT+2ys5p8aSdGopoA6ooGKa
9RV/f8Vj3hRZJvOhyRCEXwR60aSHQSfl52FKb4AyonrAI5jDxpAg06287YwiSxqJ
WkJNa95E4/DsSq0uPddeCmU9RhQebOyWDjyrHaQSZEEUI8PkXKNO1xfhQ1+l2/WV
fFQEfQLTgn8osniWqvWxtz8d5vrIJ75UQSZ2Dzhe1jibunrds/w+gIir31dTUpKs
jlbJ8R59nky6nli6DQUgmkgwA88U51PLYtY7J/gmhPnGnb7/V+l5JQs826bbJY+i
zG7+M+fk9Au6UsQypcFXaXEAyqeAix+na42Zp7GsAeqqNcZ2ubgermyCSu4FQEKT
zYtI9kwFnWGXmbPT9Y4iDT0SuTwcu3TpQ1a7tgMDebaOjiIfPvmFLjsnz40ZZEER
eDzCftgi7typIZbBoJ+et2JeeA/R/WAHc8qgRBC7lIxfPnIwnDXSj3bvQ51MEeLJ
Rg2WNdWZDCyXFSBtDyWRXdJWMxuatImc6BK7aOPuoSUPHII1nr6nGkPUASpAtzX4
D3/n90fXDWvqFYRiTTLcz2DBun6rXkTqczUJG+om38WMmSSImXi0bA0XNpowU06A
ILxSLmVmcj6IoDQ5Vxbluu/vVcuUeCyVt4jKBMgZ2c6mhyvnE7BXQke2ZnOWhV4H
5i3cP+/TzCrW0LZ1A7HTKJbUsGOJddHXfiYRfMbSe5IvNRanlmu+/MVpH1bFs5tt
QWew2vw1HpYNTIexgrk5bydrwxHKbUDupHfMRhCZRyl8C+Bs31noQy+4KEvY56lg
qMfVDUI26VtR7zpV+kRDEtTBTumyo8ZXafwr5jQ7Hf1l1ifENKcHAGC8F3clvIyt
qYeQByehKU8ENVGS5SGSRfiIwwqDI0G8sMEURBPEfKQNz0p1XmYSTJ8QlAmr01EI
ZIuCvrFqZHEYcyE7tWgntuz/ahjIrWACzsIHoatfGIFVNaB3H87wSmowbIy7PcHt
+T/Vbw7zuwkkM5nMvPpdT1YBSy3Lq6Ih0vBcJuW0tU/iBNSn8YyN/mw2LX+lpqdU
aMqZssLvGe3GdDgz4CE7Iaf8J1OEz3lRN9lKEQwuQVxgahe10h8C3o3gpKhTQhYV
B61uzEwoPHyG7XcssoqtCUasySaZrThcPK3khxoRoCDtxaKHBd4nJky+iASlhZ/p
4rWKE9jPS/+aq4uZGruqVUthkADD0BOONffgSqiw2hBrf4CJKu9D1mt3Vh3Sp6Yj
zJ8Rux0QfGofslOj0k4AZj+2MY8+h+2oITtqGuw/KqdqsuD7ZbxDRmKiqEhIDg43
LWwxiu8iP2P1iepp9qJrQSglBjN244j5nuvisqzLwkRJrKwW0TB/ZhRCgDQcftER
msYxHSfQ/XyAU9QvjfTFQFSqmWHOG1abvs9SwoZM4U56sB/dUpOAd2faczRBxoSq
kymSxSdPUODpVpEj/3wguqVL/VQHGo20Oz5/YqfOg/jYWybal5K4SoNqA7vlCJco
aB7F8kyw0T0kpj3xjWVpEiYiNBIN6ezn/PC58wYm1NA3eQTiyhEDpcYBrwxiXQVk
YOVXchjhKdy+3DdYaAAz+aoeoRbATN/r9U3qsXhYPHSjmU9K7cLSSeOCpdZhM1W4
nYlEyiMyXUcnQgL4LlpRsSzRfSrBHHYCobwAcBhTmr5QvOLZZ80D0q8szZxnUmYT
Bf/AAnEsLDwiK0ADQpAaOR5H3kvSDVLJQ/z8xv508DpSLZlhCalhqjFggHUksxMu
78uZth/ss1skw6ptLLPou3fB74rI9Xy51vbJHWM/OnHOanyIlmNE/folZLK8kHyj
smRwv6QlBSM8ng5g0JKbUoilpXQ8TxCdOxsxK3XUHk6/BkZv0j6M5mOLWYg3/8rD
uZ3e46Lj4x2O0BvY23dZQyh2dYkJM1HwP0SK5NtrVVJi/unS5PyvfpF9odLwF9Kr
k1SsPa6CW2k/6nhwSyHamtc3rZz1k90QzA6MTyFlZqzHwpo7MrM+h8OnVPB4H3/z
WXl4oZdGcOjyFKMdZt/gxneVfZya7aM+puz5XJXW/hnfliwWQwBMMCHJxkc3mUNb
nknX0ugfNyRaGY/ezAKi1p+E5jxamQ0+/qUv+8IMbcliqZcQCKJZlSjgK+FX2YQx
OnIYXF7Ht9uJVenRP36T/tIXUBoT8wo8etYVNDP9xlQsbobsn0kgae5XbkeOugST
NYVNbIdSAaIi9jP0CVzhje/sb464vIVri1Jq3eX42YSqnePT2hU2v+Ejez8Z08UE
1jbaI9+lWRh2G6eLywpG+nnd9bk6DA59Y5wWktH5tY4W6TgTcthUo2Qp84o11XRt
AKEewg+ZxMsOv+6CTZ5lvSbfFrw+hjN4UDSYcXFBoHFtsfxyAa6Yi1ePtRu8qWWF
qJaeZdgDO/BHgpnMS4dWpSC81D9VwBx4gtDOdMn61rNPJn1JojAxeXpIZuS2NdXX
TlgdXuzR0jbMsnIFkIus+GePWF7xV+e//vKEUvsAIHG25dHZ6ja7N0ryXLlZwoCL
2I5MRKv5tTB/LfWiwVX/aub+hL9LQstQ7v0gRUozVYdDyV1O5QbBjr+AeZukn4M/
cj0WMYxjNCdE8pDLUfV5WOncP2jNLlPcH8mqHopaIVKD5CDdgKJYUsIdq6V1etdc
NPHvuqSRNyzRAJ7xCb983/7sDqKgJyLFIWxK65GX9vP4vXtxVNYl4Kgywg+7yIw0
hm9KNyKrCynK0D2pv/yBHn/IOcKFQwaxQw3rpoKnwlW41xaAUMGcj4ceoAdoI4O1
wpPYSzNH+ePdMzpDo2DNVgXv3vAKzSKkwKkRm0NUoZo2TpbcQI5gLP3CwOhHtV53
td3H/AItC7XdNbEXU5SS2YQ7y+PXw1mh30AFUsHn7TY6B1N/L1I8S84EZk4w2GmV
PuLb7pEsh0r26uExhLLUDeWrodC+AoosI73fuItZWVri5+kqKQdA8KQgXaP1Ao56
nxl7tS8riRkAIh+OfJEl4wmA8YxDFRqHGmDiiiVg1K1lQTZJe71fNfh5iXir8wJb
fK5PJs2FOmbB336MKXlrL+Jr9zrNjWVUbHndfbOap1Xgj1VY/zxQ/nAoFqlk0IEh
gAfKVSxZcmRIYn424E7k00jgbAfh04BLSofzIjX8xFUDv3TahPsNl/YPYpR3BdQ/
GDticSU1rtq4RaM0tYfF+jvZ97hfIi5W7s1C3kdkHG/CI0eMsEo/96ctBd63vUV3
UcGeHoGg79sj5np0dvyrjbEvYVGLYZHUC8Mo/opKqWNwgJNdCJhb1M1yww6tC+N/
1eDN+EqKp9sjNgfZLWKnxPkVnVJGb+yrAPOtZbaNHN6sHa6dBvJf3yCcPtCcZOcR
PRHcWBXMubzzjQu5j+sEQN0wuMPvvYzQaNZpgraGI9NH8vbEWvYsJyDnsUSHE9KO
kcD/+bEB6wXtOEFEtpq0LXIYYF6BBNxDyOS52gW7fSdqF1ElTEvHxW0eruHSQHwK
dkTz9MmnyYIiZ8OCiGzk7ZTvn+RxhOPgHbgKc0mR4Q6SZ+htmWyednhDm08tstum
YXzXG+T8B9lhAnr3MVkCh1epIHZx6ZwSE0sYJ0cCHFQtU6BvyUKPFEv3LkqhhTqu
eFOgNUcRf9+NEj6rLU94vyjOit0JAmftbzbTGMCy4TNiD5ar0wuNF85S5AiWSj22
ZldsZLNbHFrhogeTDrcoNdlCNeYKkpVb918fHbDk64ZJUNbBRNW2mxNhui2oQWm4
hjeMzZ0Be1SoX478mx3WA2tOtJlVqFouiVd71Wv1xmoqP9GAZJOplmSQYn+kJBsN
XHCh2hjHT30q7NDp+M9MVQSFFujcNpY28RqZr3+9fnh77xN5sQsa5fbvs7WZ50Mo
PJHEBbLHGTm3cM+66XAQZd7geFy0YwPkorfqFBGR7P/mwxg4xV/5tN043plYtZIo
qFz0Bdp4gCk3PTJ6eTSj/DdzPWiEWDnFB6Ej6Et7stXvCXz9/JEhXUlNmbsoep6N
J1YudZ0OrHmd2r0+dTis40KoUPHPjXKnhgdCPhmQdVwAY7wRiRn6tAQS7YfjHCKJ
ytJZLmTCGHqAL049Ve+zMrAlCqbd0YcAeVQeo2vOT99j18UqhwlQ2ETiVKuUsFvv
CDWhKTaByhLcf5+K50xGTDdsWKso39joWEnfPek0xYpNjo9SYYMA79CuubjG/nKD
iWG9riPIMBYDIWBk1c4ptHOwJt0NPG9OtG5V/Iafwn4I2tQWP4auhw4eDtb5UE4R
OXCTuOKtPmbNaJbY/XMLLP/mgzDdhsrq3k1GMKlWcoTys6XLaxCcRh3/w9VW+vbx
Z9pCIqEc0ON4q/KP9Te5G/lwckh5igZ6diVmcYpbNKqFK6Lyx6K6KA3PTYP+Pm3k
cVbg4+SzRES23lxFfo97GyeA0bpUJ66cTBEIvV82L5+Qu+B6NxYUApkApCxRi4GH
p3TJP5nODgGoDPfBkb0saZ5zDqRLZib5VOAw05LiVaSabnwUlaNA4XQ7q7xVLbpL
Kw2hbO7XGYgXJi4vZm8ao68EfxkTz9mH3Cx1uB8+gNYFYMnqvJyOfMj8FbkxHpbJ
TrUkP8Qyjluy2Na4J0fJyKBKq/wcbqF25O2ikB84YWHEzRYqo11gDe6LhWRuStf5
EaXwtcVWqRlbmXNKJZ78MVr7uuuxblPW9eVltI8SOeBwUucYe1xTOya+dIKpOYF+
Tb0JOAHIWsGh26EWB9lMzxBcYqOwlrFaJRo3W0L1rwsaEUm+SYK+Z6DQFUV0sKJT
bzAKcSkLihSapeML82mXQG3dEtaqiMNr2tX/Z3ttXyv3/Wp7tCUeMD29pIuMEv+g
kBcg1bLccSqB/Tnwby2tuUHrwBycFGoFTOZHvEPznLHjTeuED+mWYJxFwFM2qZLW
VYjnfbYFjEzOoFf/iHw7Gn1rsKfOEz+hY8pxFlXYNttO0bdALfzh0IDIHqlpsfBG
du0pa+gHXNqHY20PURDRk7pwbA4tWO02CYd8vTvlwuVjMAI25wHAibLEU7f6LMyd
W0o7OG5ecE8k0xAhUtJA6rlHz34hbhCC+2ltqUEo8fg6qy04AJUry7i4jiNAYJ28
zYgjT6j7QoPFvfMvjgXRroKQOith7z2wPtIadIjILIhSmyGac91rQrowMEsj+oRg
ifmegFW8U2vsV+2yLL0lCzS4dIvYq1nRX5flp9uO+K+YEJoAKv84lb9bp1Dt39tE
DJXDy9cWctHAAvVxVDorQYNXw3k1JIt8PYDLckfHBuSQU379OIR/xmYlwOFTWybe
xr1x0WUF3h6HzG381ghr5xSMQLPRwqXM6vMlTYCci34WEvRX5DMxK+DkgJACoKRe
azt3aTLcwEaHWxe0X8wAG3HoxwNv1y5lYiwZ/CCXzXgKVQICr5PrcmYaxwoN5ApF
aXzAJI99tX0FU70tYjyqLbNSpAFNhr0g0RagmO9Qwgomge1xWUdKbEN2pDOUGMnp
Aizs/0+hPIHcAoO8/7yzwkJpayAzMniLR7rwoqVOrN/65cqJM0EvCsmGBaN49MGm
aA9RvK/3kh8nfBN6TXDQbDnlyYm0xBuppapWGW8lL1EQhyBUjsWsahaBO6i8jfKd
ArCHNJTfuts0+qyqm9qdHGS/NKR+snso4cU4igmT7ee/HxcSkG7G19qjneYI5xte
mDHUSNsnKSCLOt8MOK3XvDaUTCSPEWB8U2OgdqzLx16nR2J6rcGUse7lB1XWF4v8
lBcyc2qI1DBfIQtk9zPwNHpi8xX87fmk3QyxBse5HDUo5hr95BF1Ybi1t2b7Vuzb
bwA4yJS9HSULtF6AsKWvGL6cQQu4U3erY3RMZ1azVTGDKtENzHDbcw6n2b3gnwp5
hSGoq6PnccfTuRdPMHmOTkFLmkKW+Ae9TgpQyzbpKlPJz9rWi37aIIo741hSBy5h
ZKgeBhGGcJws9mJZ4CEPnAIxzdwIIa5tUbmvL62Ge7IrmR/ajKTE4nz7pYqyeLRY
YJYPF8S2ECvNC2CR8nI4nCQ1iozl3hwLiwPlMIWsB5sWdlQ7C3bJImqhUwflgPfd
+rzxw+RMFQ5z8qXsA8XuhHATeFYm7w8rPabPzwn1VZPUVEr7jW7RE7bqfWsRBWeZ
fd2dL3BuqWSC5mRBpPAvRqt6yA493SlgfYux+g3b9aVI3zjNbUC/onZa6wLS2wL4
mBEq0JrQ+TuPO3qsot4BjHbyWn2JqIt3emaj4c8m+LyvPUrMYSF4h5ga7X7ibmxK
H7ahsaumSqSaUVYJY5BHn1cbFrj0FuzlopzyGrWsC98XyZX/HWnwJjMitUXBt7lu
i8vOmh62EpVDCIPUEKuXbbNoEFzAuBchTcl1Sm1NsL4o1nyK2gRywd4SxdazLrsf
51cDYYVEsrp3Zo5BIrbcViDCMJvd7FPkwcqE7AVNeQ02/rcT5feO5l9Ht7owpQnV
vGJaNEY5VZiA/ifr5FF4cLs8DyD9x3dNoBTCU6PqbP4xUpD2yD2gQJJqz1BZfCrl
Tvd8fGZgTbIvVnu+zCvC5vSyFcppU4xupGUag4M7Utksp5Hd2XDR7uCj+GwY41S0
jPS9vkm9JUVnl/t2e5FLxPs5jNjTVGwVUx1qMu0zi36ipnuHo91NVjSCQyu3+iaI
GvIOYzaH915O5ef9m7Lk2SNEjp9jxnhDPxfeN55dBqtgboMNQwUI7mK+vUgQcT0X
nchZWuo5G5CppgKZ6gpvMwUmbZuedK9pmXwrN74JYbl0yjKWOrhbXr5ohIuqVJWM
RTIAa0dCkIMAsgQdjtGAxNSiZh8T4GSuu42VC9HdyMiRq7ccdpLrmkmtJINtOsSw
R3BgQE5Lm3VvUXbTH5ISkmadZkhkxnVllF/2R1cO4sKU6TB9lC7bA9o0dJ0TrTIx
RwKX8FHWVrPvoDQ/RnIptXuc5dDn/taxoW8jJcIu/UJ49HdmJLW8vncCEYllpHMn
39tNGNvjZn2uBf/FDGqz1BEINL8z8XVsGzhOSOsFPv9KhyPoJF7doRRrT36LPMjG
zC5jgR2JUdrTZjqj9OutwHmP22y1U6rpkEoh31lsPU/CwoUg+G5bUk8hqHwc7DHN
fDfJ3bTSreq0iZNmK7FoBWmVJ8pB9KEKfYojIEzSsWw/OF6pzMGwwW4aNhjlDRvP
kk9WRFgvVW+KBmyZdba+UlHauKq9GmfAhzf0FTJtH1SgrJ8xqAkg39oZO2v8fjJh
2aIhWWLwWR/kL6serIxd5XHPJLo6MPUyzDaYiZ1lob+Ecw3sVdP88AMhN1r4gDF5
KpBm/BxXD73rmDQrbS8kl4lLf+SFTrp0qsKARJuyIAILQDPbZYAPYfAXr65iE+dJ
DVwXlqL/xCrm+/IkqwW8Df51eBC0yPdaG425o6whmZZRx38k3xMQC8DofJdxgc7r
RyPiF6gFHJl3N/5LaQlQYWYPj9hfl25wFRlSTP0X+FdgGBEqNjc4QAnG1XxLPIpQ
NfVqsS42zND9picvc8q1SpFRPsWyaDWfgKiuQ838QCZDFmJ3I+rYSEQTr3d4m5wQ
WMv47Lf+zb0BfJ2WUXmMUOoQ/yxHSp9zdWNbSJnaULNzoqcwukkm8tiqAvc3Hrjr
HjnLJgFkMeTeHMXZU0JtnUOP26jcJJtu5cN24xHDq0P8FEari0sZOwB5HYAcgpZJ
rYXV+xeoTugaYaMExwEctkGXajKjnY/dykgpAsnsDnt+fFUH08B0bl3vpBdacEj0
pUvrY7tOt6X7a77XMLH0kdfsPeTOjSQ7VuoJsRUPd0lrV2SzaAPQM6v9PFlGDYd9
1fQd3ZzR2w+jb7aLEJZ32PIPAAjxIbgExKofGimgpt8jdXufZLnEGDLcNr47ok10
lff68MebgPCee3DKybYo9fH+6a1jc0/eRhNwGlnEzjOgO6khZf00Z3N6HdhdMAFB
GY2TRrKv+G3lodot9HqA/ogumDRvP/DGM5A/nrCRuf1uYEkfDWVhPXfC9lqeauCL
43SBMWFJgMclYk8cFkrOMSQc/oNjYsdQWiuENyDNEdePEyuybT3xIdApFJXHKz7y
fj9mtnZ7AdEddUAmGqGEZK1rFzrDTVc8W8GklTHDpkv9V5ni8bZP3nSr1O7m3a5b
b2BL1tUuWvvrqJfNOlY+mIoE/oTygkB6ZcxSOwKHZEPaS+8kUM1C57sjYiJXGZGn
O5O7gQUuFSeoxygzbtqbaoqS1p9wSR2Sik/Y7+tCVqAMl1az+3dqhoitN97DFba9
bQ7wluw+E0sXAMROpqt+9j7IBaMi4SvQF2qIx/kyRkNd2tGMtmaGD7LzkWxTwfWr
gPUP0GiVtfrOE+TugnT9Sk//H6zXT7qBYGTIyvzFgJX6728AGwsX3DeBfxVywJj0
GL6RraYc8e58/J2WFNvYWeRd/eZpfxQDcLn6P/oMtjb3gPkUFGTmHsVHNHCJKwKg
i49B1d9PXxkoMgA98rPaJvonfKkAZMUddIZ/cWiFyTdxOLx87AczwRoFZKCQ4fWR
/pNpvEL0CQDy5k5aT6PvqbrSXP16mXATcDu32czpUK1ctXO+1FEBWd7m2+eI8g3V
X2/Ixyrqzt/5YViGDseIeXmiyf6JCm5PIwnD44AzbWBnNupnVL4MBXrOgZFuhIxl
Ersjp2GcWVnUk2qk4eBE3Kip/UK4in3KkX36yqYmsmT0jLNH999ik3ROp+Cu71yb
GgqXFafwPqhcyYqldZvyNPu4MbUKH2FZryjhDMGWI/z2ET5NZ4e1xNS76e2/htfd
Tz+xs/HTprwtR48+TsRnxqGpuHGzgzSszJNH2TpNC7NUfBFjpIxJe4Tw8R4GNnpp
3vObw9NMVaiwLF6rFZ7gq9JI7C4+gklqMvTPsEsA6oTXuBiyS7tfsxVDyPuAIK90
B4KmjlszjEiROmujuT+9KLnv5fRWLvC6Xl92l/9yfLxqTvFJaVRJU0NcU+iBBs0C
gwmEqU/z169z7hGK0T2PL4DBgRcov/PKEv0/TnbwYrGNQWh0YRJvDlPwmcqtRRvr
SBHX0q5JoTWn1e0kwQhCmogar87VSPKcypQS0khTeWm8ReSDIcFGUIQMV7rU8vT1
m5wiOpgjq3jMJsyxHRiWaJvPlQ6Yu4WciJr6gvlkc5avXNDBYNohsBFlWrTQ6+WT
1HS4RI7HNWR53MqWx+QA3UeiNBAIsKNTaiKXfea611c3a+5bEDiafWVfMNAyJVBn
EQdWjHF7eb6Sf4QBhkGsQCvd+Ow+gJMc8v+SjBx/9+6CndDqB25zlMP9gQarQ0Cg
iWTzYJwq8tZDEx5Yw9DPq8GcB7O+SyPlltJ1pfnFkqg0UW76GFIAdqevHH5A9Pmo
w5n8s00sMAO+frPr5r3sSRxdvBLyKsXed1wUSK9n0CZr5z55dzDlqdVrksl/IJla
RM/fiNSy7/OwPw1IliX6Si8e8QSke1R4PPmqNd3AvlqcWpCYM2uCL6eiK28VugVH
tiK/V+Tsv30dgp3cgbwxldy2VZ+T0C0ElPjmgzQkZ6E2TYDKtTlK3Hqmz1+JU6k0
5mD+2sfSB7sNLT7Fu0XmQQAHNrjlhMPfpCeIiA0VmI43hFhJd9r6P+K7Y4/6ELq+
wI8A1+4hTyQ1RPtkB6l+G5vvPKIZ4tw1bRQdSirfktUwpSbD4tqZyEu0kixb0Vg7
sxdlH3sBFvDz9i9pA6LNPRCnKWK+KF0AO1Hq7TXRJ1wJO4cVFVpSOX1/rD871c0h
zKzLII6cyyA3OplcpUPB/OOhfvtcun6ILY/rHk6dEvYeR6waKSujb/+G8J/ruDx5
TRYhqrP0Yf4S6DqrnconX5fhCWuKc9ONNPVxbzzQdCNWg1NvnbXrBNpaD8Dbuafl
tAOaqJZWkmpe2pkMUw55KqxF1cdFcjM2xlfTGgQf6UXLu8GepAMaBEauJHTAYM98
s2s/zbR9WFDVgp+m+qAOvwPDwWSqJrGw05pm1yJGfAbXZOKA9JmTlaDsFBs2yqeP
6MtTJWG4qfDCasbU8/aRI0ORUInJ1WxXoAikwNcJSZuR/k5TSMjfqGo/AFj3tlwJ
cNhJq99WjM+R7jrl8PQB+J+CphQXQ8S+tzT+GG3ItMBPQ0dezR6osvvQX57OUoxQ
FlDY6IEZZZE5zmA2eA/hkgiyQYvrAO545vy3SwEhTPx2E366Sbun5RBlJsWVLGrB
wZEy3lTbhaJKeEvNxgF48WkRBJ2VAYhm4YRnovdI+fh6RS5YIpIf3vkX3Xf75RmR
8JcF7q85EOhWxgcE+O8NCj0hFK/uCYDBx9BEsuMzqMXkfs4af5Z3rJGQscRN59vh
cY73F3Ps3c0XYEgQxebPoaZB45gl2xY+rXFcp0M/3CT6O+g1Yw3G88Fbc2vCqaF8
mvocFS7bYS4ACc4/PVeHwRIUI7smZQBnJLkEBs7S9M21OM84JKYcrqfGmKlfQR6s
34YrsftmIhfb8ed1zuPo6xWmEEjQVvQI2H+ObUE2M4VvQKzm29xXT47AWeecOI78
ybbYlbMWdTTKOwOdPii+SPotGfo0oWCi9cjCpgyXwRHudw3eWfd8pxtE5/QjL48Q
gUzcuf/Hbbgh+zprzvEC1BRYMrRRPnCdMamLy4u7psDiHp1HMAnN5gug5H1xzes9
B743zDEbemHUP3tS2oAdLucIsTxdhT09Yg9HcruVj2Bq6KsafBlNY6L9B88iFtXS
ACcnEY1Gr4F/VqOeVhjffp4QOj+wdTGk4SoIqkgqJ3L7Z/5aas/6OS5NV+wMocnk
IWFZVCdZBMqLq0sRbAYdKUDY0GO4Z40th9dIRIs8Ozt0brRuGWQJ6RCRoismjVdl
zlznHHFH2QbSwthGslmcel7b7pU5ZkHngQadgtWMz5XzI01UYpESPejHqyRtus0V
pPG5L9FISo4L5MxBtsjgilBQAzxGdcMhuCcoW+giQkzH8mTgAS4XDT2nL+uIxTeM
Y6A547huBLyIlUv7ircXNAe2yFcRdR8NhbbAJ4713c/znVBeVMSsm3ipqrEYT22E
tSlBW2ZDNH6Vp7nY5nb2Glx75aWkllsUJHi6+3u+IaH5lIwiwgLRflB/D7JEvPLs
fqF96MMIcqZvDKeWrjyBPlr5KMx3r1nMh57JVk88T1Y4EA3eYOCk5nF75OwMF1HA
oIzPs2UTlPTCmJxRSbAqi0izDOfv2xptn3W9Psid+nnB/HgOsGB5G4UpuNBO5jAb
Akyjh8qR39OqqkhuGugKoeOtS+jiZvtX4J+PVo0A4zFqN1PJEpIiIOsRRF4JocIC
5i/pft62beAOHln/FPZNJWffLUb4oa/PlIYbtojSHS0T10pw+Ab0/yoDKi7V9oEY
oQ2MK6Db6Wy8vNTCWmESx+lq/X2/aljAwFgApbfvsA4XZAQee7SNFtAz8KVR2HrZ
jKR1j/OyCpeponm7540qfFUFSQLVBPNSBt9ZLmZAjSbSbS1j731WzmNvFl5E0ulP
NZcv9a5QoMv1A7GBropaDFmYN+V7z8w2hKRIeQhofEb3t4kr/6slQmBdqfmYzES5
AD32ozehZNHTQ/m0OnlCtZa09x/h17xn/IdxjWjaGnt32+mvPl9vZn+8aX0+Dk3t
Kc4WHTI7Q+h64Q3044wWvdb8tsfBanLFp8Cpjh75VqtnIz5MECq4i37SjkaTaebe
BxWx0W1hhFRsuKX+eam1U70ZHQYZMzEvNVyEEWlkqnLj2kC9TMsOtce2MuSm8Fqk
R1cMZbKhZMkx99CMJwN4qS/++nFgnH1dtlKUOXEdSq2OaNIFFuWIIxXn2REf+CmZ
dsLWMrzMjsHgjeyRKnuHSKQZnB/WPwGEDGqk/nBDQOn8lZ1prx+uM71skB4WK/Dj
oj931lHN6czjDLj/SgejBYhwPPrrDCxX0zXiDDXDKFK+gbwOwTtOtSImduGeN89E
wWPAFSU94vrFSDuzLlyI/XcZNdGgDoYjWrVU7aWb2ao8CdL/+LSqRgLJtdw9kCtx
V8vqzEYxxDNNsUIzZ2AJqRKofubCeqQDzLuCXrCeO+zuUbHEgMPgqulqiSquoyHW
Sd1qyGfr8EnGjvIDkJrZcQwsRvmS+AFZZj1hEOHYOnQc8WpBfwsh/h/tGowLV2XB
EfEg37GGxqvObF8Eflc4mPS7zUk8yZBzaDrzaclKk+ITwphm0YYS45nGmcjgQA93
/uWJmFq91ucluCxy53v8u83V/Mfbpuh/4lLo/Y6eP9WREgNNilYnLByl+ePLWaTi
eDiyVaQKxSm0e1WxUWkPOpzk5tTGTSBaarL+12m0mo5jnGG/EMtOLnW+6snLoQf+
G5I3BImjQzeW7xZJe8KhwrzhnjJdaeYAqViG4hpXdx0uhY07xxmRZU5owRLx0GHv
F+QdvPEvW92Ndhb15uuE5uMXFClM9MdHg/m5Gjz4/21gi1jOcmHPU/0XlrqXZ8yU
3yIOWfrkfRhKwWAAXgMzgIPf7+ouCHPWcWNNxHxyEWgOr1YPbBjFkZu4VdQOVff+
x+LAvff2olM/Ear1Hn7XSbDz2NEtQ0ZioZCZZix2SHKlxpLst5If4C43TvQLq2u0
Rkq8WsN8IgwAYST8XEQvKenWq7FPK9zQVhVeywkLWoA5ZcT5DwCweSv8ejXneFBM
7dq1VxeyJY5ktsdoIk23UIFBWgPQLIma5H4nxIWpfzc3HMDRlzUWULMnA2UVmwi9
KM2ubctgrwHfXRELRXeWPj8F4Oeh43T4AaWSPpEMUcPB+ugoS+4lPchuazdBTRx+
eqm2eXsKMZ03Hh9CVRjvmEg8f2/Jg7P5F0itrx8vQlkgDBd73JLnnJE74Ata/K19
ym7cyazyVRDt5R9F/r5eJ3yhM+t6sE3NFeH+mBagWWk1xkinUbeBKR+4+So792fj
B8b55eRmMj5og2N0wja9JSkX56o5HNjPXaVA5NI6XONSdsiM4bWC+GRfKBOPWHe6
/lWjwP69sPSXRxghxon3xP0KCOXlYhDbDhr8pEuxHOExKE78xTGwMlXy3Te++NaY
a7VPA9oT3kX1DBkkL5h+u+EO6j7Jy1tLlaRf2/993OzODeyM4iRoyqUZXf8JSkWd
rz4Gl5Njd9YCDfQiX9mv4ME8qupGTykMvIGLylBMsDvg/kqA4CZdc4sEBzG5QgmB
rfY4BsadMcDwAE2kB7aX1RinVzVPiAtOobNmyj4zjzTErX94K+b4wzpcC4lwvnPS
Gu9ZMRwlq2h05kBfczydZmjAdGSpZkPCT6Jkrlfw/dHXzbtIC0zkUN58FtNZjEcd
bOLWDAEXYdZsMQKBLPpabF+kwZuA3Ta0j4eBQXsIfkw+lTkNvKCdkds8e/bGjN/i
ZTLe5hwm58idP4GvWxrRVTYH+tdgr9cIHO1KD50pbF9SrgeAOoMkIob5oeM7yi7b
OnPgMbytXlNp21eh3YsdPp/sROFQbFfMFJsYe4aMVBQfQ9NtdDtwQt6Uph370M8+
jSpbSJLK1P281OLOqNZg7zuCAk1vQrkz+muea/gzKoR+kltu5esnLq1MscBTMZaS
n+BAZ+k5Ynl9o+9EDjNBz+pioepAmxqsX6Ya+3v9DrSprh58Oj8UDMWC5A/IoH3u
8sABkPwOjCBBzRt5QaBPw5I7hgETu+QXJT6cPNd0kLbSTeq33AHoWnOuqhZDGG/d
RG+650p4p90bQi8N51XBryGXMjreEYPmH72KyqQ7iz27HsdKP+a1vp+8EO27Cn/y
HUiejacC5AjMXbr3tisgVm/SeahjruXScOWt0H9Z/oyg4xIMRPKax5+opbhterZ8
/WKy95uo5IddkRgYxXJ0WAOKb1Rs011+UpgxHQ4cm0YzYPcXp39kx/3rBBOEoBwN
V5DqnNfJSaFiYcjSBmi7YKNLNxpKIdwLT+Df9RmxPv5cMUw+sPV8x6miPCqP4wp7
OPaVy15UzHkTbEaLMM55wTEv5B1ojZGnelSZcwpc5lCkDAT4MwRH8p8aeOK9S4nK
/fhXfn7PXMEOephBfPSnuD87FsKypdOI+/xgJthpQhgOxGU0DyVOMkz3bQHLTM7W
/HlAsYysCC8jkdtAxqRACVzOb5T8n0k0jVGzbrQOxBMAujmd+X/ZwLymFn/t+yFA
PPqOlynbeFwpJuCZ6ofnNqsdjJ4x39SD2MaFLFuLOwoIzNFzft29HqjfLRqhBot8
j/e7oclPvYmT7Z9imXp664UT+kcyD7186ZAoZhaMYDc4VnieurmYBoOCWI3X35eN
sSRvnnUw35LlUlBU6yDcK4fpdUATA5PPXgr5lOD7RPwu23MZfBZgSfHPg4pakLrH
QL9ePeppdV5dc3qFt4ZhuPoiqU3ULv0f7BTJJfK/dmCsNdkCrOn46+yGeTZGBiWA
rAP7EoJzLWIEwTxwNfmJDrk4C8/NzOq87ycP9nRV8EWPLSw9HdeMmXZFFsh60fC5
wELWBj8BnO/8G/m+pywFjBd1TvOoCMDDBodqITsrK1Txb3DOu/GgKiXZCCfp/CUN
W4lGyxhbrhhRvDsNtiMfE5Xpv1QzuB8EoID1uQzGmzDZ6EfHJy328Rexq1DSMqRU
vYMkcLZKDlbjoiuEI12DCBXYwVt/YoOXLHrtvgJPm1cXMdNGIUJBW+BPXPdvPYZS
L4mmIkbx4+qrTOzJNJXngpE2jf9aEcYbH+e7C4MU81aslZWrjtcTDyhgxNwFdaBF
YkswPRicIMqfV/IAdsdemrdFOGtLzyUwOePQkKrGVLF2Iw5EHGZLZFtlW2FFroh8
WeKJI2icmjqPNNAPCSEzeLgdzflAAIaS1IZOLV0EJGHUmcPi91XnWhhuDwy0hou6
C6iopKTGS2ofmweZHdFsuYOIyRFIfuVNcdxKbi9tcBcaRnxvy/eYxqJb9DVmCu+c
OZhNxvUjKtt0zbdjeaFh/WCqbZlu5I/CVxcNMGC9bXpBgEONVlRWnPwKT7xIjhy/
6pEbLAktiVTDjwqR9kiojhINnP0VkCNxxUkz9lSsN6QPgwtP5nuAgJJUrE2uPxs3
U4m/J5iSnmLAYzjINWS1qpsuw1q4c5JlARtuSYB50H9GpIsE3VmZtQB+sivK0dt/
+XSLOzpjioQyPkd1FTZM1a4etvTbvy/JrRMS5RRmxMOV3O9PzW9RMu5EY6g3rXsY
HHagpepK7olfavBOvC6BUgjfyql+k8CuPUfXOSKkO7IFoi5nfVZTQKMXZfaC+JhU
KRPFZrVKwhSWooLV7eaJhyvldXBAdW/UYqjr4+RYzJlXK1gD9PRam7zXbcT9b0gb
XoETpN4889K6sk2L4KvtKY0fZ8WlWEs13crCmnvqHq69GD0qytv3JpyeJsFajYOM
6LZchar6FOz1vCUwxs4G1WmFt4+F4lVARXrQaW8NDAix3ddPWwV/hXYs+9ZVJvQz
vy7cHn8jczMYWh21w/t/00IS/Ea5UhUY59A7tf8v4T2zpc8o+fnpy0d1czkg7AMZ
3DJx4nXNLGe6aQWU4uyDKtzj8LSKr4GUU8s4wpkumu58AOle9IIYBiBtYD+PeU7E
9z4JBEBN4CiHXOUZKF8cHbnYWtEnsRqOe9minEoLwYT6VxGClG0U68m5h0N/Id2L
vsqxQszZ0QNaBilYekiPyEEbVPmlpZQSbYOKEzjXVP3Zb0PzXvSs0neRDRlxIQT7
KBemv1KKzKEgBBwNJ6AUtZn6gnTNgHAltN8jyfOH6JNFLADa62O1s5dyKoAuWQxA
VG2rYywWKgkaq1SMwm8ggzGDIk6AgtWZN+tMVGzDHZUtTDRZ5NcMb2/UTqRLvO8s
S4l3rfz7hj+gj5SpR2jBjXrswpX3BYHSp6HBsNel4Y/HxET815JpTQONfmGJyjSD
7zWpfcwnJ9XDnCYrQX9FDbY6PtQrVS0Hgsa6GankZ9oOoOLPEh5AI+0zQ14fCd7y
gewb9FPP0qoB+PbW0T7QhepP3sDFx8UC841DSd7TQFWQhsplhidwDmaSFEMhjZWo
1MMI3Th4HUBv/DnAxD/lpcfXfeNsOKkruLkjc1YpOBKfF58pgklkrChcnqg87vFj
q11ZjTTrC53dql6cRsplAtw3DecBUpVJVj6AirQAeNZdGmxtHXwq90BwxYzKYE0T
udkH6OD2pfv7q9wDLRQ+WU9TEoposWPT701F9mkXCP7x4exek7mvJbiMshsiCMPH
wzEiVuWEFNCSrl+gOXJyrvYfAVuOje+YoGb2/2HcBkttFerQL4nUe147bb903uPx
s6KKB3VKqddc/HhbM8Aq5TLkLD/AaJCHFraYLlOFkEHX5fv9fyslfSU23GnWuhTr
jOsML9iE/kWXacuFMThc3TiPLepuRYHiIm7QMOWf5SE8wwGhOLIHwGF5RJgezBzz
qqPx1m19wOzPzR003KUV4+Vm49m/bf1kP3lMUAn95ZjKBjY/UvE18L9Nqn34Dbde
tyYaayEdl8bl1ETHiraTOufM7bsxCmAUGOghQGvevuBXnou3+630sAetpG+mmbSR
rTmy3B2EyIf32Y+x2falvGi11wEy4mUs/aFy+H42e1Z+AqciEP5XykntSC6/m66Y
aIWqtmiI1WgiX2PbHZiTxbtIK92pDwUHwor5yhO6M4CwjnVxJnhNddeRInnHOuX6
TMh5DEkfizpX8kWTYnHcFJGdqX1LiIWMboD2Fr2OAhKdLXZF7ClZWHDB32hZJdEp
88A/1263mJFCICrhCI2SZpCpI2nUUhqJyEYYUyOTLS7UfZyICm1ZSF/C1rcDx2s+
Z2Tc+2RzPiTJXiAU5mYflj+HrlhieMFqBVoilfLzL5y21ne9cVaVd9BZ09h+K3tS
JrgpeJamC779pkuGuZXKvs/fQ1YvUoJy/0+d88YQC1QJOcaedOiXHrtpdkI9WLMd
9hCrfmAKoFdSLBRFYrhZaH/1T2fKAuO+hxZlGqTTNWBxfvJFvn+dbVVzK85C5b5e
joslVrM2/7koWOeIkV3QKnwa9S0plv5QpQY4GYcpX9ylfuuqFh1eb2QiYe116G/h
7iVeCW3wIWbuczuRFXzDAtox91MFmAlU0a9LZBVJUXxzqrgQHugsOTCHVTvk962c
j4lpcqmQ6ormz8x1J7U57fYMZHr5DKv5Gf1Gasgnh84unozDxbQYq1Q4nwXOEUP5
30Br9PIWbg65cKDsAVX6OeX4wn+cCJr6hJOMkDOiMp08jo/3MdYO9q5uZeKK+Hv2
zlZ/zP6l0qg3bMktSbaBTqMHWgtGdteRDGIp/8VrkRIcsChBpIPzYn+amCbDFznd
rNnjtgVKK2vPcp3UrprEHS8tAdqCfr3qscXKzhyTvfVDsLTAjmfBUkmlfeFwXz3F
chkCQiT1vWctyA8B3DdCm8fz01iSuycVUm41DZ62T88/ChHPfO78XC4/QZk+/ND0
ictEg8a+ANOiWfCAiaioZSjVGy3WP7ne5eVWLXbSoDiGzDOYvy+Bnddg6yX8tCXg
WXJAzdn4cYCMDYWqO9JUE2PYZmyqJEKY+L6+aa36b9CxCzTOYE5IRRexOjz5cCYK
GW69rvneTZy9xIwEqykEpezLsYWkBX3T2Li8TQ9mXKBH19le5jTlytpudXyoTWW6
XyRv7Xqag6G+cp/H5J1uHaqnKtZ1nwsq+DN30uruKiiVRtH//fbxI7iD1KKFJUmz
S1NaSCD8gNTm1pI+7X2er6Q15bY/xSZF1y2KSNgJKbO55S82D7rvCZZxSYMeAqJz
x8ehW8yLMaB/aOgIdbTfrBmE+dwLT+M53vHLC+uvf5UaXf63IrELORM3148DROz1
anjQGfhw1dt4+ood5BfDGnrCr3Z6ReNzreounkaBqujMlCEHfQf/zrz2+1mIxoQd
KE5nlZaZmr7IS/Gf0Oe+1Lc+gqzIC20dotW2FSYKpJ6U4RdQYwBWeWw7JB1THb2j
MVVvf8vOKti8BAinZ6X4k4j8INPMiYTpE0n7GgHUxMsHaCi5VErgTeKhX5rGy4V5
81et1ZMqOzlXw1dtl1sVBdA8XqM8QWOgDnnzl+wvU4bSCGucLq7cRiX7FZ58qIZS
DJU3cvew9tL7wCT14Ndbj4eRIPN2kRuCBR5vopXnSzx1lqh4IqelQFePKiYKFEBS
y2svH14bT9gbObAWhT2JrFD3qAM3yHvV1pGoZloK5mV4J2o76Oiul5G1PW4CgEbI
ImJEd5+PCbf786wPLVm+V59NbIc3dIAc3MjnCCRpnMU6j7Ohr0zG8mDD1eCVZA6N
jO7gb+Gci+U+HEY6kXFPPqxVC1RUomEJQV2jXResi+zgLMO5H0pIJUlWuA/6Xs6c
XTIpYaIJYm9CK/e06SimzD2zVq75jdwp/wqCaM6Rm2uDRYgccNR+pZZeHiybmPU7
DH0+r2MwkJipNyrF3zlQkbTixD81wwD6itC65pu8K/ytJN6sVDj64xgvTwLMi4mX
Hq+ON5M8xEO+bXCLPLPEkhxu5Ze/OAx63eqcEMupO9wlh/R2Q9/PWcQ9zDzgL1Bu
eHoBSjKsUJqdvwfjG9oiUuHakzuh7WFaZ5vrvwIkemYqEEgU+wXagooSiX11A6eN
2m4cFBFogkauC+PeREl0f7Sj+D39wYylD8riSRY0uY2Fv7+urqqihafhLXTkqgJo
03yo2cRhtKs/PkqpTVYyn0ToyJmEDRlQ6w5euGonitAoCzc1007uaSuQZJF14Qip
23oIP1jbjlSlfUVTNvPjDSl9BZxa3XTHg/YcM4bB6nc0eKbhxHKETX7YrxjNOLMj
Q29Sl/c/4oyV+vUkeGCg6ZcjrBa4/Z+2yC3s25/IO2q8uK+cp5mBDvXyQFMB4/wm
9CWMMhqJzVZiua0cZjLZRLP6LKwl4hj2Jp1khtRV8uhk0n9cB+BmcCkUkEDoXQEy
rsMcnTcuFfsOXCi6ufbh2UtbA9kh5UUxU0z9iidR9CYFxEiCMl+IE+OrLn+fcRLS
zjjX957vgne+oXr2kdok5x0SBNnusVFObVudg3ep+5XnJokxxwgUuZ0IqI2uxDdx
Trm6jaxXBqldFfHjkeO4Lsi9EEpIytrG4rvp0DOGC3p3KgTHnuQptyjY+U/F62Ix
1TG2V5iXXPyMM9g++XRbIxn39aFiv2AO2TZkgZyuS2LpTq9K1xRXYKI6XVJibKhi
QCV7QdrK17VqvW8l1vuweyh8PGz17qIuneowT2/TONXvOJ4yL5gpZ1Qtq75ynnoG
a4mF45FoMK/AnPiGSrwdyI7LEuIeAyI0SR8XWVXQgogtKujTbso+JkrM+SxGJHLC
/khx+EH800JPCQi6+I8O73dnRfLOfOWQ6xedvdWW0N8IOIQ4CYuM6eD2psb0E2Yd
JHYgzRlfOlfJ+KyLkAKwS7cK1N9PpwigynVy+EaZ7VxsRW+lOymhpVgDBa/ZyY0E
S+39faXlsdpRYfpkLCYUrrZVh6Kv5nuzDBDfSB7g7PJRat1++M+zypXBRgJVAbui
OxjZINguWYttsMxjQt9+GLALzrQZHfGz1YRjEtnzw4e5MQOlJG088wxBld3ox6Y5
zZhOH1vzJWqRRyp6BOh9carF9eaUpK++5bwfSJvRHYucGr3RUBkmZhZM70r31/QU
6NpsmgTN9oTkNluytPVVxVtvj66emw/JL1TXCWGfLQDORr1XhAtl8bwgeLOGELLf
JP6ipXiEXzyF5UMqLRWMrmNz2A233IvgBBu5LglraY2p0Pukymlj3QV9G8a1c0W+
bU30Tpxki4vDQzmLQEt5WeNtKQg74XKDMUB13uS0vW9KC04LOr78mUYhdbWM3vSB
Zo1B6YFJwmbQvXDHxQeinyv22StpJ4nV9zE7vy3IAxLroKSqrwrp1P58AX9fKArU
tFsXVRAILHhEHcraCPdlwrXRmdlpsDRlhmHReul9ju7BA1WKb4u5kvdxWPpNA49P
nzewJuD9z/X3j4mJTFzboOzUHIHYWDRlPkGb1hvfelnYbsgecEctW0aPXoozu/9F
fC0GiWu9MAEAFpVUDxbS/BBslIuQPBkrg5kGNSmz5j5yhhojAPJE2GlodjpPi9+h
jP3993swf/sYri5KIHbKN/Nuh8m6Bz0v4nDTYTfON6Wuws10is/u7V7iQ2yfL3CA
cFVJZxXjsfgM8CxsbRNxPk8+jsFXtRZ5mhS2CjnbcHBGxsJy9cTVwApSwoZ1msfr
6yUsEwVNMs3bZ4Wevsd7JecbfxPmADPpUggUrkjZ0ulRLYOUwInIpohVBr8vW2SU
oqPUpYhJj1RIT+e6x3gR+7ZUzx2REDcPjdcfS03ZB2/HQ565RuLXQKEmwRS9SD/y
/07DUaajg6QBKg4W794fhyI0wpni+IU0KBo65oxCFeze/gMs/NzjNa1xeScrOu8b
iOj1TAAFxxqoUKmu3osRonSWgEngInoFk94RZa2nxJPzwPvTxX6Uv61O1TjhXD12
UI8Jai9LFryxcDI3O2TbGPAtppVbpHR2LudUFRaWK5epEMOmeGS5mHT3lY00rTNX
uyMpx+Tw/JAiVx83OVKhwQwGC7x3Oc459P5s6uUX4PLpowR3yrJIeKiLId/vxA8m
i9E/E+ciys7yBGGdDmUT7I9Mk/RSl0VwhbVlw7BBR/qLNaYjs6PTQ3z5lrbXU6Va
UCYVFtzWb8UwoU8mYjsdtF11Ksy11au8jjjd23KdeAVfr3lUBwf1AUR7zLGXRCdA
gUsi3gJSMtUBn5XCii65eWWz851yTrS2MxjDOsereLgeLFAShk7X3pf47EgAiM+J
Oy5IBkBZ/tgnV3UfD14A6pRYxc/TeliQ/9mswIsMlDNbxvLJeeb1iePLq5sJgDBS
QJ9Kg+YRDMHXbaPV13NZ7htegnOBe310GG1Z2CFOxtFA/GZsEe6rI3X3LkCQ3mv1
YqDsbzlrDANIJO5c+ma7ly0FRFrFs+PMzlXbCVUYvovPKN6i0HOwQ4HpJthYnomA
3MrPx78lIwGv0uUpDlNy4Xi4VBLWlGKTpqN3+aV/hZiQur3ZI60jlUOT6EHWbFxP
loXhbuVa+oP4l5E8NRbGX5ov8XzNkpkRtADrQe8SL0+de5n/V+r3r8pnP2rs4xz2
VkWTywKgJBzhZsr3GcdYHxT64Sm3iv/+4NCOM91+gdAnrZYGRNuTxqkmQwt4pWms
hDgSCNw6YSfZawLaEgXR7c14sGf9w25VnbaTacGSEqeluLDy/URjQWB45XDKji0k
3pK7/MAAjlCYl5Y+HOnGeUJ7lVkBP7fIr1Kx5q5q1Ej4pDT39MHzBxV+CtlRgOyE
eECo6C4AscNmvF/3OvOovl/VHVMXnVwIErj6sXcrqiWDX1T8X1qesoCohzQJhF/1
YOWTv3K0XHdfaD/qLIaREKbNLICZwXmNRSYUSz2GiilhRNkXebjBd/su6hF9tk56
vJDx6A5Gi2L4/47iK/oeT/CcZd9Mxoj77kjAXONZcrvns7UT1boBem+z2gwEKjcZ
ApEya1VZ80gqtkDei8SVeCoMjYSfcfF3gQVLDhrThLG0NprejDrUf6kqf26PVQ1o
EWRnsgs4ri/L8EgFG7+1cl5wvLiDwOecXR2tII837ESu8NsVJGgdI55DQ5EvPQrh
ZQ9SaemmyAL1nMtzOy7hydtFYE4vcWttKXOdTebFb5xmILkp5v1zG+5dJhbFNlYX
D+teekW+6haaOkBYWUyvT1tifVxu5SSdmyYvroQdg97LQMPdS1yBCRUjDFWRO5Ir
BpCmVtPRjZjclzGlZZpTRHVV+CRty4Yp8RFmzIRJkrkfXQZMEigcuG4s4bBfeph3
0qkDtlXbmPDaeVcNQJQR7Qp3/PoyeMW2GRsfI9KTpCSHHnDS9uQOZbs/dr3hRNOI
KX3yvxyZ0b2iaCyX+l8AWoEZylQJPapClp6bKfAmW+0EoyGn/5/4gIOqWNWUghTP
RVczoEDovfREnT4dGBERNf8uZXQ7WYbK86oAwZd1o46rbVOoYfdMlPTA8B8F2qXr
bWncbSlpAedABJ3ToJcNSXI2AM6VFBCCwqJY7Ffv9ACm7rtfESiFx20Ytc/xxJnM
Z6CY/MmQYF4tFI17EZar48AVokJFdc4TefbbL3Fi3xByaPa3Boc8IxjSYIItJbZJ
GhFvNlb0iQGkJImB9Lsd1GHqM0Xscwb0Hl/4BuHgF4h8JOlmqGuOr+KE12W0lomN
u27IQJxoCtFMcNLv39Fwv9f+iu9Sw/Kq9RKsS++pHw4FmIrucS5BBwIBmj5jdzhu
ny6zN4zytk0N17J1eI2wEGXmvZiOIg95R5xyZ8d4WW6NAGyPB+PAlIuER28lXIRz
Lrj+An6ZW+dUmIz1lr9ClMvOTGneJFFtw0X/vH+abKIDRCAMh6N+61C2k9Lm0aYO
9KII1LzJr4wpK8LlMSLzeocpzkTneXO/x2eMxONQBlccbWuvWVaml2wm8zyNtTEl
Oi+0T7fFJeC67D9ab2FyGDuhXTccLjopGuYs33G57a0yId8s5DhEz6apGbJwGGZQ
jPXlpS0mvt8BzMWcG+cE1IwaVxaGOKiFY2F/nd/M6XFmcQRV7U35cFhjv8VSONVT
MNv2VJiZHt/D1e6kgouwMkl1QP4homGx07Gdo6ACBrzVF+gx+GSiPCYPwBPNYwsQ
YZKUHTqJdrFmi0SUJ18APulBP4fenCPh50prDym8NvYEghLYIf00Gebpz5lgALyc
Vxsmbf4V03jyMARAcg5lbYpKnpMhQln3NeEop+IkxsKgMUVgQVfKwVwVx0VxAElQ
0Ul7/++4T216q/BvdNKHIh9FYe1qIGJXcmmKXIUekHEzIacm85ettiL7JfzVBO7s
4v4HhyM06boLsS4Oy98CGo+Q0v/cULCUNih+IeeocxFNpEgpbHMRa6KvBCQA99ey
Vhrt6hF4hV0Kx5/Kfdn9cRCNUHXv2aKM/WWYtNxxtJNLLfqByCO8MNMYctkz8Jvb
K8bJMwMJ+hqFlj2TgjvbbbrpZYWC+VM1XORegg5BxAORXwXKSpEDJaKZDTp7avFO
otAjalya8pEy636ITzKYDOqWpAJL+LpelbPxjHpOhANK/pqEw00RAa/mqtwifMpd
nxQk1RM3Zso3NhfTIqJKsR8UokQ1lU8Z0AEAjyefnjIde2gMhAVWY9om3p1b3lRo
2e9+FyCp4o/GDaiSyXKCGkscVMjLfeFWxR+xLi+fb4/CQx3w6tbaWAWy7kk0jWyY
Q0ASxmSmHUFbJnWOvD+s/dumVx7xE3V4j6kv2xn/H0fI+85Gwtpsd2H65PE8U5ci
tKQlOVWvB70esyWZR/RZ0xjTGv8RqlveulioA7hZ1rKk9F5nTrHFpcsLtAeP5owK
FxCZlc35TyhCPVf9vxfWlluR1xU7EkQmqD8vdnav2m3XaveGzt9Yr9lbcF/TnPzh
1SL8/XQUJR2hEFmKQyKMGyzTzuP68mOmfnYrHPdUTzPfSEYqce1ZMfyL7db+p6st
j3EclvN3VllP5xTGtKC3awZ6yLMpo6LdCWRZS2vnLQi3sJVhcs6aC9faEPnfYLJZ
4VILbFJ5sFk35Mv17BO/o62hmTnNjNAaJpfKrQ+xJmEOQN3D3aFWrZyjfEfZXqzb
z1TqlOZK6ldSEx0mzhoBPSp40UBe8RhKH+8ymE/b2jn8oIxJla2qJ3DSyii72RXh
L9Yl8JpAk2k+7kl2iwZsrMEvw8913crPprm6icICgeES5kavqX0GeKow035u9xY8
DJzXbTbEe+irdLaVa5oiRT3M2bBIcQWXgBCKYnEx8bfV9GF7UXS0q4PVlo4XAY66
Rid2YMcxLc76kqFfFrq6oHVIaR8qbdTClsGN4YCaTN6+CVIlIpfuAekIpOZ0DEOS
6gyt6SObrqqY36XGH8cysWQIbUnBcpRdApJGmIlSc2Z07vsKDY6UQPUnIh4qzP3/
lFgKPtzq6VwuYgI9M9SDzRlp29J1rMz3tYmDGcWNp5v+4nJYdKu8tlSOE/KvrgxR
S4tO87FNYfbPnyfpP2rUD72h+C1rJGQQKqKkZfPjiWC8A8hkvhiE1UCuF5EDP7Pz
JhYpbGpHsbWe7+XFhAE6LzElMJOJL7ggcx7fNzONHEY1H0inSGR2Hn9ymTIU/oJ5
MXLm/G8Ubip2Da7644dlmMq9O0DZGH4wFeVBilHEpu7RhNbGLiyReq2R5rFViuTf
imREOQk3qacy4+U1/g2moNZY5XFK5kfGLI79WAcmxQ3fhPhoJOwKgAYTqumSLaxZ
QP3jp01LUyPvejNF1EgqujLz9xRzVfO0KF/xSljbtTZAD+cEnCsm9TGC8X0I9Cf4
+yIHYamCTufwTlpd5WnA9K2d07NVMDMrmRQeHlram+X1lHZKMrYY1wh4pxNQQvKF
SfUsuINLC9QEzRuVwflx8Hpb+Li7V7ux03AuMnPTL6o8/DQpAdmb4IBLvS+g17rV
hR0C36Em6qm5u9njZ70LM0Z2MjAitdkadfXmokI+MYNtxyy4es5wqjiXKu/dbCGl
MmCHxE7ztxZp1visZSu8jl/qEmCRMSfBeMvj+sPPjQYHWTYA9YIzKMt5yFd8VUFV
3MV9dxGpUSaRst1+y7BX0r7OKpxGXC0Sdi3KCTIZIKeoO7xOCpNoXJZdUY9jNGxM
Nz2BRmLxMQn/nfxbf+WDcbI7ewmsWt3kybZ+r2Z0J1A6PCMG3dpjlOlEHN4+zL5O
rarT1wLxKaj25cRjYTcUMygNTtKZJqAY1nEOp4/iPT5LnEkgcyKZp2fmvdD/uhqx
oy5qQn9cAi9HMO1PsqdWWaL+UylvdeQhptJX7OhkxKWmnLp5JmD1Y+3w9EbII3T7
0csphb9odEKPdHw9fJS3FYlUukWkgZU04zppyHmTZ6fpVMzzXBdWtIU/wLYRqfl4
yhHULBiu+VHOBqeOpI5Ha1ug2zQiwje7EnS5n4CkvTt3P5bOuMpFAGh9FIpvcR8I
SFiB7C4ALd5QwufygF3q3nEU56O97F6Y3Lap0hRd1QupbH+xNI2zimuoyc/VmlNe
0tn8Zl09VZzolNWRXybT9G13Piz/i8jDtHfn3xITYKzX8yZPMfNosJE4zJ77al7G
aIlK9BzlxN/3Zy/L690RM5pySO0PoxQB0HWepwtDoSit44dwBqCPgQhulatwsh8n
HMMvezuJuGI2kj6yVCSlMBpCzLO2cPzN9a95lLodIlgXC8W1oe+5r+RmUH9gGgo5
`protect END_PROTECTED
