`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CuzYbwKTf97exioWyOaZc24s1hrm1pCoXc0agKfwukpuKtUcbqcvuElslD2adIhU
pZztCztD5MYKRvcxSGTFefmwn5xOyTT+UR0qKd4rk/I9cMhkftGYNnxVgeny/QDI
3kzJWjmaVei8dngc8n5avRUOcPzQ1nPicDvWGsNzRA3DlX9gP5KPsYb1HOIyOfUI
HxtPJcdJR2H6MuRfXfXmq8BZLduEDP66KZOJ0XWhHnGKOdvtHcpAXZ9dO0G5013s
fDktcMXn5KhJIMJO9k1dWc9Q+NhzfpfezxXrWeiEEHYqxVnYTKkjiLHLYKDtB8Xy
nzEMd955YDDJK4elWF0rC8ZnMQ+LA2RbtIbAmYocoVxUTlsVdXr3FokzmhQhD8yF
QzBP+KbD4j/rAtwKuBuJz9VxAJLwEacmX9NHp8AO00X4CG56ENfIeDL3ZTnWQfx7
jwAzktKm1jrqjqQD7tRWbxZDOBLkU2qwYUzEpYPVcHM9Of6JqfmAoPR20d+a9GGq
XVwrwbgp5Jz9zMBr0dVuRtPukDKZkXFlPjfD5G4zyuA=
`protect END_PROTECTED
