`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CyLNmYqW414EL6NzFp3nKUs0V9IlamvzPkaBKzCqsMDOlT7n0B38KkM7AX44KfuL
QYnITixIFJR9C1HzQdUMcno79taUkVmqjT/xmjdPphJ0uL03f8ttbkJZLa0VcB8c
5I1/9BpCeeFRzczYApGQUBOjxmA7CrrUCMRfEj2wnaraXuesCQbI4iNHZ1Xh7cX9
6NaXz6WrUGIcdN3PrW7KAsmTkM+2V7yFC9DZJtdcP64yia2VnZOcbYC3BtydBrIo
+C5A5O+LWgyHcA4vhVRSKbi/1gkjkcXjm1fx8F7kSlf07UFkvVEZn1nhy+0Hjszu
l+HYzuuvGw2v27wqcL89Z3ksbd5rEEQKs9SQXuVKfX8r5F+0vdpvvEO5BaPhSwEr
KJn2qO/5QozCKZHgmeMNuA==
`protect END_PROTECTED
