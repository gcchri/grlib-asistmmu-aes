`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3DUzoNm6FucMIHSE4DnAV0sJwDiwEA6HFvsyyufXtj9aGNbYwx2ay7rfkfLKLn3l
ML2uHYhEVp0KLiV0yKBFojD8WUUIGuy2VxmJrJxAOlXhEHydTDpPfnJkrQqxfZaL
vS9PbfgPkFztinIbNDZw5T+xS+xo5OtdR2RYggGJaaw9etlQJIWNA1M52MuQ9dwB
95WwgiXHKIwR2XsMt8CRBJQy/qtIBGKDfI0p0XBUA3cZA40OlfkARzti1xRbkiab
9q17TEUxN9wGJ0uRNYKuMZFx7cYvaLBKNSQRFuQABgnQuM+YmJgJlZsWvuCHuN9T
neMnIUWAu1ybJH3P478DKPl/tLQZiqTGDh8Ree+6/ZBJ0N6pTI767F8YxJSgHZkM
8iOmLPaym7w6+3r46WmUt6b6CNsBkEGwzML5Th6IiOkWgUVnJSEYJAmXcbhFSAgf
qm6tBYFqgCFexeIUVxBQc56jatOVFBwi7yahf1oYl+/VqJyE9CIpYpjTkrfRD8CO
IeDO65zUMFE63bbpNjB4LNX3thQpbCdRmS2gZSP0US2MZ3kFzFBHKAlrv5F34/Fa
7IoM6qelBAmsR15OA6amgH4PKjUGgavzEujRe5Fp0/1zmckH9dlmDx32EP41Ndz7
RiSiC7iC2/N6mMpQ4HtelVv3BqJykUJH0KMt+QYOFio=
`protect END_PROTECTED
