`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
clIHoZe1Oq1MfSPIf04pr0nmqfWlq1FZEKeB1ZRklJD3vR3kuUFlMEXHZiOWSKA4
QPD0WQOLong12t0fy2ooPHF+IYDWyZyNrrWmldhEhvjgUZOiYIifR4+CF6PMFnhq
hUrmkbMVN7iLUbKXSp9Pk+BVF/h6dWnH2yCAjrTQm0kvKLrpvgEwchhj6sBQhvTQ
Y5KLVFRndsR9wUCDRUJ9+padpAg8yMajSmfuz6ABtVDrLhZ07yjA5XEY5Erufpsi
XiqDei8uumVXqtmCVL5vgA==
`protect END_PROTECTED
