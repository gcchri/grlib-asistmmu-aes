`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CtHTvTWF7o/4RU5QfLDTbn39xed8szwlj2zHGOwyQFCFup/zIOkPMdexidKoCSKE
6Zcvo7KJ80owjOfJzFPtxBcQaQvd+I/5rvVl0iu9QCjiClZEC4pCkMxRczh4WAZn
8Kg6dXab+M9E2/sweSUJjsWHgB9xwx8W3RgVo9VPJY4kX94++X5LDG1MHtjoZKf2
HLQYu0ic9NDVrv9PGpvNzFhf2YMuIrFclvJm/xNtkt4aUNqVD3GKFexxDHm5RgSK
Rle1lWfGw7uztT0Axdj8FelQt+SWM+Zd+LIJtZK+dnK/Zb9pltezYNMPekb6D4hB
`protect END_PROTECTED
