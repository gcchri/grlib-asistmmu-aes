`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dt1sXu7NRh44R29JMqNq3wEsGCYWDyKFEFVJfKjt6oU4w9SX7zuTofxgKx9e6YTx
SvvwQb53FtgCSX5pH+6iXs5d+thE6X8gGXym8rjtO4rpVQhD/5jZFNNuWtvJDIeu
bwv9gEcUny5ZTBudvo3DrydoSt0RmLvw2qUDCOmLkE+Gtjbkf5u08HqIW09EDFS6
39vz9TqDGGhVzgWboXec4DxseUZj1Gv5R1Cd/B70arU39iEuavq64VqgCOdtJxV3
T76s8IHStkuWR1XDlIpcXg==
`protect END_PROTECTED
