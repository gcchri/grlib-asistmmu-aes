`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKeLpkEG3cQ/VG4r8i2lau1r3h/qSqxPz0hJJIP6hBAEyLtQD0ttmjKsqmPdrN/s
as+PmrVc8VbgSd4Dtc/tU3Gs+2YEVpagFv8cQBz+TSOVtPZFxR5trSdXMH8cV5y9
ZH70Kq2SzR5f6ibEox6xV0b9BZNbvP11H9grMZtheQkb34qXx1kgvV+7iAcxs/Un
JPorUuLJOkFTbIPeE64eER4dWQ73+RRK20KOkBKisPanmUbIpPkBCb6APICrs3+b
Ccybdwk7AY4BCnJBkIF2/6Pk1sUR/R6fl/RzhdvBDp3YdwOKsMButAcjiTXHpy9M
NDN+ZpECPZq+1KwH9Qr9vXsATszQ7ik+ik1GvItdWMm6/XpBn3sQ0qQLlLYJk1fP
6U185TzbExLiSHDGbjNRQiyF5gYmPgF+h4QqWMq0+CZuG7odDj/oBaNEAEFKrtva
OS2W3K05YlnBBHmmWaQUEw1xaZjELNViV0sBsi+S93KGB7fCJ/X7RGRezNWYSc1E
o0AaLi3JBcn1Xnes7FbcyVIQwB02KMfZEaqhCsIjfQdlhsf+zBbe+KrWB6mAEJ9O
zoKdikuugBtXcZIyQTb2Zg32ZJDEBeu2VmSWcDNUzh+HJC2t0yZS2NPC0EKsmowQ
pzRcc7zXNQK6RpMg5qkjrNYvkz66AzreJRPexyIpk33BwZxkPFwEF6gNU6Xa1Nfl
sE1NOBLKVPCPih35qFzzQgTQFFKjLhj8gFNfp2kvGI7svnzL7UgocRErD6psI9jy
937y/BSBgYRJCg916F5PyM2RzslVZXHor5UHAPAaJ9OYPrHyXObBAqoK5WP0vlZ2
Gc+F68iBq/IIBovQOf7FgqICQjy5ZVi3hVv8XcHR4KHsHSXKDGyNt2ahSgpXLHrJ
ROIW+OGNfXH6rdGPZrvxwFbStXj28S6WeMeWX+6GvmzG90+ZiB5hkkwg0Wt67QMa
GdKz7z5wv+8HcWPqNvzmXV9zPciq0X4odOINjw7zsMIddGHGBY2jltgcg0d7xQSQ
JwgpLeYmDEQZN3SmSU1KLC21NmllD+HVmQDze59VCQsLwJdyt/FYpecwvlVJGJhd
pYEqw9MauA0WHFSSPilVRcqxrNbM3AxpS+QJsjriBWB0FifQiHnTz08MeuchMoO2
JxqXbDgXQJItN8nPqeUgtoPArsLLmqqyNJg260h83AKX1XFyE7d3eYk57iCNcs2H
c/94f4q1dvOk/s47y1k/MoabY3XPIyA6fyK8Ucr28NunM3a5tQMRxl+gvb6edxHc
oS+4Dz7moMBk5AZGYSBLTSSAZssRMrXKrD75r8M/lSSoGAdNZrtFZ9W0nnaYumhH
/QqstVsLD5ufWFmp+Dege/XUM3zcakldAOIjIwHCReGXvwAEqa6y+DHzZwdCtiXW
H/n4VqZ4F8i/rWecK7+NGJlu9Hm5iOfjYOegag3DcPzth8gQDTxXAQUlstQ2yddY
SsL1WdYuZGfTQdcCTZkwvoLDj68/2FNlysAGtByqUVkgPOp/01zaRVHVizWwtBXV
BMSX3hWdNFVnlxR5rq99YqNrJLNMyBhiMTQnGZIuv5yw/VTKW3bntUfw+HmbWjGr
Z7kq2Pl0VNHWK13Pw2h+frg4dzXyoHm7pe0PQVPrfkzFewS49q/77bgR2UWw76Ad
arObjzf+SPlWLycSwZjmy/woK3PO3PkJOiuRX6taVNfED+rABvmvK9uLxrzbfrlJ
xat6Day9BQlT1Y9xti8SxF2QP/6geULNDRtHnUcwTgdCUBHMiwFqa3h+t4icE+VF
xA5uCTFgEnN99TwGzOFaPg6h1bi0u3z+alLNFd156X1d0MuLXr5+nfz6B0SqnSFm
1XY7o6lho6RR0OXp3c6+Hh33WkR9dZZzk5EB0a+rqv06MeD2ZtcZb852G/vjK3ZH
/+OI3l6VlVpuvwDTDRr3aEuCJ0BBRya7pMZBSdl7WExFAZzGrzCTKGEUIRaJxniA
5yPBxbJp7IcLTlQNIuaaLrJRsw9PFUaevAw51VQjfw/S+gj0IKEauFfBWlqQ0g6x
hqnNhOfwdnaALVjzDKavfIu4QDkeepdYASeAOTMbgO8LXegGwhdRJMxIii2SZ3Ux
2nzu1+YyTC3FdHbYgqXEoTZkKAU48fRfbfPxq4yHRqVvvMZxt6qfgnvxM2VuKqUW
MRjzdkV3d7jlst1ybmSBlR6mwdY0DDdHmZ0tpQi5o3CR7MPPJTa+Vdbbx1DGZuWX
v97++WIyFGul/+AqHXZxH2MGv/DkZUVHGZNQSQkaD240k/tB4S+/xseCGBaTMr5D
xcSOiz7zZUqb4s0XCGlMMcMCFhUVa1ixi7jnvnYE+b3q1QYMDMR6rZGSeJ8KoikV
oOg3VMPmiIy2cBdcGOF2wVHrBpKJ3mqvfrvyVwHvekoQugPu1R05KpimL9gwTx9L
QYE1cUh5FiX9j1uPMWSLjLGGzMvxgLfpXHAmCIyPaR0BJyk5uO2zS0BfMd/p9ee9
rG0emyYHKItx35zy+O/JY+Q5i1gPvJf+ZvXjhD+kLqJiPTgJBngAJlFmxaYmKFuW
aLIlPO3cYyMOPyA35l1XIqr2AOmPB/JNwYDn8B0y6Xx3WTswaOiVuiaMsABaebkS
mTqPVeilmiDEiKLffjmyLIbmhQLdyG+DbuUQLTKjDWdtVTP4pqHz77/WbJn9BvpF
y37OEfMp2sDwJ6YI9Ue4DZr7COeFk4p6Ck5i9ab3iPlFeaiZvjSv++VV7FgP5+dC
dK9CG1YI2pN1nDf9ha0nIGU7xOYG58YPTJvR1xV3RZfeygHUS6Plz12s3wN3ddn7
kGVjftR61NKV/JzLQuD2qRvjvslM8bHoqYFsppMoyMv0qTn1KGi0XpfdRZi/fXoq
uhe5n9VeKmzXrsDnG/xwwYXGMPDgetuPiD2TzZDdbMmSlyPCSmzulAO96oTEy05x
ub2o9qpch8dMd0u8hVuRVhtUyC3oy2NChqU0vfnoUx2MtMDMQq7gHXfvx9a62S/H
DCuFuXKL0Cl/Dt0tEs6oqwR+9DlDvuJOAWggYgcincYgH7WTOfPHZvHSaIsIFVIQ
0+4GKALFZSXZzks3v/CkfbvRffzRP/45IUv9dHi+4Dqafy9gtxVEyim2YfQqUYeS
kTaCLiB8i6dhl1agEKlS+ziQUVMJqsnEnbE99Ps6R7o6qO93pYuxSDvUmnPbvSMY
GDDVRYuFTKm2xzDGcLBSGxD8X//4nbIkQi+MzNCnUrpXnOn12M0UYlu+SJWsdm1d
Bj2ITbkN3Zk7TWp3k9njbswuooVqFug0L921Dq4XaymDHo6GTBQmH1CUWrAprtAn
`protect END_PROTECTED
