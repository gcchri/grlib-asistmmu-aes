`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLR/r+Oc3Et9EIi0L25MEqxYk+BogHUJ/t1lt3GOEVPl4IouGDdvI63NerRq9lfC
d68N2u5Zpglj/LkmSKavZZAXK619jrlD/1oKCTkPsKXsTyqegOwW0tHl5zq7vlNH
N3W328s2MJpZAhqLLiVbFUIdoupPIV+mmbKtwXD/eOE3shWZDKuKzPosUA9rL/+c
6fmwkkBU+LJuGA2dD3i2LtgdgYM1yzZim09zhHDHenFJKUB+2If3rI+KgmOXQNnN
5nrOWeQPVSwpCm0QCMWx6edtSa8AyOQPWU/Ny8P9uRcqToP2iuMy9gL9CaSYGqHp
cfNSrN07EJZtK6jFJYbXFOJI7PwmO9lNFBwrjEHRepoz8n+d4WvVThqZ0gCJQ2Fs
Tw4/OwjhV3dyCnKis9DagJubWa5I11MzItpQBqsXz7mxk7AYgE1NwqgaCwAKMfS3
`protect END_PROTECTED
