`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXq9zS7ttqAF3OhrOfIx7fd0RmSWdaxIe+yQmoIi2Ie82Pr0YPsUpz37Z66nKWVV
24P2jttBCeIwmvfOaezMZC2Ic5cPqbqr0HQICYZFGvcrxKsFw/++8bhnd2Tv8m1z
roX8ZyXEQXWHMXU0KiQssAe2mQEiWLwItMHrNECgAFJUk7ygh6xMtQjtAcO+nFMC
ZbiXx05Kz0NvEitO1TDl15XZo/VOsjBFu4VuVn20EhwguCHOdtCnGaD2vF4qBboK
NFzon+gmsHqMPd1KruIIafNoDnSoqMN3rNRYb2GS1/bbP9hoRv5Ls6S2zAMV8cYw
y0Sl1EbfUlfOcXK9cIqdt2ImMkzlbdDLHoylu/HJqO8eik69w5EgVPbbkR+SdwzQ
cRYuIUesyh5iYJ+DNclYeLWqrdLsS5EC9WJpWQXMt+z94A3L8/mADFhs3fjA2Hvz
2D0AMf/LEuKt4kkvSWbSMkXyvHrIwslbUddUIRJzFmydDNNbtAtaY9skuIZaAxUF
u71RCEVCJV6auH0xXMci9gx5JtlrQzfjiG7lrJanQqUAPdMhy/t8WQJ+cnO/MeAH
EWLaTPCWnhBvzWZV1Fp5C1tlWYeHKD6GGBjzLSciZ7uc4VdJC16g6x9Y6EfoktVb
mJvNirFuVXg0TXx1fqYDBxP785dTAxXU1cf+XUHcfv0LHiyeBzgS8EmvMC92NdKP
uXwGC/qgYYTf4+YSiozOdEmmz53e6D8LFDdWUlQceCt9qx/X7fJh/EIGnnYkvDqK
go46c6M0wYs9N/fpFN+FJR0JZkM+5/FhxXCi5/p7MOe3Q+qvdtMQgxt3+i4AsHAc
v/cVHthM9N/cG6BTNrlBzzwjyodXsp8EDMHR8BpMlTQkJ4glmfH7bG1mNdwn8BbZ
0YcCSejnnoc7A9bUD6p1wx+5VEAf8JzqQcvAoRdLuIGuWsoIqvwNb1aPbIURZo2T
FbKNM4i6wN2CSzXm1k8R8Le0tlrlvqvYUONvGchHllV1D/q1MIUdwLnvfRPkNkJn
w35QhGO8q9RikdgLstnaAJgqUxcT9Z1x61+3Fyp1sMTz2SFSJ8d8vV00QQ6rUJ8j
gSWBv8j1l4dIwVteE+LVIC/VjDlzV/0XodVFjfyOERgUO9Gg6HqhtgEo+Uo/oWxO
mUjz5/ysPq5n518799FAtI0MnBcGvVMlPSPbpy5hAK4YvSmRok0yhRvVf+aaazP9
`protect END_PROTECTED
