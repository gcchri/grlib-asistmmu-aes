`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6v2Cf75IsI9zyTc2KLS2ECyBNWe4A/kMQrovF0W46Hbyy5SHsPEGtVt7+k9gkpB
5jxn3kw6zHiZq2pUP1XJFdy0GQ8cP4o+JwBwZnk4Tk5bXsg7yPRIHofm1/R7bVPL
W6lRQPsaQqZhPtbSRFRego81OJpuJRYMXblU/R2gzznvUnSYQ5FqcZvlpw4Yk0oA
/6v+aNbhiZ9i0kBsLGVpXPE48yzQKWJMji5t0QmPPhfmZRFxNpB1uRZzFk4BY5sd
CKPDgF8rOtStES3vf1c94CfQLnKbg4KkMAzcFek57QHhW2xrg2GJI1fYQsFtNQvm
tjRXxvM0ZYPieARIIBRaxeBqVNLA/BDB2qu+hjuLk0NhOfj58zKpe4RwV2zn6UmH
i3BL7hmHJXCLCThBf/NMHJKMBffC4A0PQ7JDGpuk4Oa78obsck9HdoMpz0qoXqre
2mFuhGgGwgBU5tqa4eF6l4aIsJuqSYehkEKtNGmZFqPEZvwx4FSW6bdWH+mO9ntV
mhYhiU1yCe6DW6lpael94W7C1PyUP9aVfMxtqdjOKWfGAsivwYc9atbIP1PAAiSp
axOxSXjksqVApfqJ2h2HuG1PmtSf40t6EIfeQcOR8k5fZmUbf3nvgWyEKGiBYsj1
ot6pzFC3NwFnagAKIJ1s/EehbJF9lFyBdLUJ6hASGkZVTqHeCQwl8g4ZaHI3lkyO
DjQ/E4+EdmzHN5AXJySuvu6uLzZUciT1cOxZVbT0WRWeEfvCnhw1VldnnT4Z/hmB
OfORmdMwYa7VDzZYYDqth8BoLGCl6NWmw+4WTaAbaQQaGxK1Pifn6KSMcoN3OM12
/lbcsFgz0SNL0VJBW8b051jhdp5ZPt2MYCI0r8lCautTjMCol0Ira2XXqe085y5C
7nq/QiVPUOFnDYWv9EujGsSAdiJD70OwtEtf29hhF1/c7eAwJs3VfH+wlv7tJK2p
KDqQX2n1P+1uZq9Y8Af+UXVgOdhmsAomIogO4hwQpVC9zPujyZMTb7ACwGYWOlkl
wKxu9Kh6r7Ud+VcmeHuQE4X/cQtaVSc4voEmzRFxCcReaLm1+WDPr4y+7+paPiEg
aWbvNQNO+n636UncLhyvhGGfAC2pFLQyHr/z5RLd67YyXvTNkyOYK9Y7W3UEglvN
a5GghJ3W5+R8HTpw984lyHAscBNmpfEyN1gjzwbvgfs0niv5psT4IybKyRHuwLfJ
V+Tc2Ko7OTax+71iDwJMq9IFwbprQpNCW36jI6Tb6BSbKo4/81WnmkKXnHC1O1Ue
6I+bUSNhhBudTGqzfPX0DNkQIaZ5E0i20KuMg/Ej/WPtuCrAw/BsCWh0nVKo8705
yLsvU4c7kQCXFL04D33sovWFUylg+vUkAJpvC02qu3MgjjI8if83P2j9BxF2Um+H
tp91S+IETWtTq1WVVhkr+tKhum4ut+YWfxReCmL2kpsgRA0Cs2W7/ehkvPLgJhNv
t84gqcFsZP3FurGXL3tPstXrmf/KFRlxgbho98AdzOf6dx+9qOdU35o/cvfobQrH
k7o3DhV3iULOOsB0IG1LVJYsDfRrfZyTrIzs9mk2EK8=
`protect END_PROTECTED
