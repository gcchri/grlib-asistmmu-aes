`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCSTSA32KFCh2HxH2ov/yK4LVb1qQa75UqKlz8icnldx2ffXWXhyaGMdiMpR+LWY
ZpdUdVAdC+52YPxSX93Jrx22ph0qv6aS4phsB3K2qwzHbTwp3L9g9MfvSyWXyGae
Jf5HQMwPsK6deROpGsj0PApCtLrDk7CbRp9H0ttJXHiTH3p9rTZffmzlc9sKOlte
/yeJlu1OtnslAxlW1H2HeGzcW2E04xJdroBeikh1zRwDwn60oI3rLB3O7beog6iL
Gx33WbFeURDFtSRHpCbBs2l997G7qUw54qAv87T1uNg=
`protect END_PROTECTED
