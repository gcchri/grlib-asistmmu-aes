`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJGFET4/EXLXn30fZBqjg22htfeOqpPI17CNBY3yb7a0Pb1LgBfMThV0cCne8JiY
PWYtDriIz0ovZ8XVyJ6fsSTeKsJcKKjyCb1zs9xo4cvWxS0tDR7OqKq1qwybFcWr
xd8qL1CGmiVtLg5wJr6PnalosErcCMlK5v5Crsw5Q84drfIIKg3qMealXoKf+Ey/
ISkU3TC4lt2lHHqEYlv3702AMXNF2sAbbu2w70u1JMKHbdcBBdR6o68ervRTMQxh
3gX6nTMwaZSjbFVGTeSYYw==
`protect END_PROTECTED
