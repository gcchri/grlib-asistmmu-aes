`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yFxQP7KKYjQa5oINCn/5eSOmpImKKCxnavWRMc952WzTHNLJhB3xg78bywTN6YXs
QFpVVqyTSBQ9cBWCAbJFeN7x6phY7EwA3njeHwpKWL60bEOJWirmwCojZK2TERt5
HkiNTsq3LJt3LRfkHI2GCQQUKMrYbT/zJULepKGI1NA3vuuf1ComwKQi6hrLdZp5
lEeckKK+ikBKT73YqXtNF5HbD+LmEZwUsDcmbIBvQ2FEJAudrWzk48xoqWrDalrS
VbOg+nDiVjU/sz6cktfPhz/xgGPm527asJU8grEQpfZNFA9TAZ4qK3OX2WeXnKAi
ZExWFevKvPcuBeD09Vlb8bbaLf81GjUwdV9U70/z6gXzhl8jLdKBwM2/7gayo5DO
`protect END_PROTECTED
