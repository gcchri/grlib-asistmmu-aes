`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iSV2n0oAibNE3DD8lex4XT85vOy60Udzp5Hw+KJ8L1lKjyvDl1XnDURpSqNIixq+
1nQbN4O7F4ozfYKh2fFm0jdI1gPRZFULPbZ7He9LPA3Lcvm4c3jcmJFQ/f451mAR
HyjD+viisCoX5JV3Tlb0ci2YeadrIDRGgfVY5supZJZ1Ui/b5OZ051OupKKEXKwJ
PhEFYSF8B5cTzGr44JQu3cpRTLciubCoTYz3OtHirSCzlMYQ1vHsJ2KjaGFvQvEN
6BghuRm72ZJmBpHT7iU8xngBcDElIUhDibWngmbtCeE4zebZ1hKCh0z2LaMbcbVW
0hpQ5KqG52oeGh79GnJ+CU1W+tQSkv5zS9zYFC9XIWfLMbHAzmX4FdC8zcwJbSyr
uthYY/0K+jwnfb2YifJdRg==
`protect END_PROTECTED
