`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3s4/tA3SRIXNmCu1m3ccWf0mtSFDCFMAmkX/Dve6xfdNv80QicOTxfiuD8d6LmBI
kOOK8VlMD/QW8EJCuBWlI9Y2nBLktBzreiMqFEKW4bzmogb0v46Wy0jXQDSxpx6B
d3cHzZFBGVBF33KlMEnPGvyZ3+LbSMsx2DifiFVSPJWMoCn/579yIXpJ8MyaKMzl
WYMzmUqRwcZLNxeI54upa1LBUaaXaynckBQnmKzyZN8+8kYlZ9IPRGUKhnA0ZZfz
AvGyNJtiZ0cAeiMJNDzR41VmHboMC2wN0our+KCejFWNC/Rq4fjBfsf2CR8574oa
EywDJd8d0m1WTV1ccnrG7BvjDWESBQlpw8SI64fL9vsz0Tjt+27RdeCMWkXV39D7
WfdHbyNQFUjJW+ADjIUtL4m6XIIrlYsZTI/o4HqNDOMEbsg/qrrzOe//KUVYYwtq
cRg8E3kjYLM7oMvbzD2ROFJiiEGjdERY2mW1mAV85Ym4qvzG+ep0+g5kZGE0XYT8
Zni/KdXW0baMPbkG0H905yMiOfvW+ZYHCU4tckfwsx27Dk2OeZsMeBzJy4AZ0/39
`protect END_PROTECTED
