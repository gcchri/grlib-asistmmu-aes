`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rk7j3w1Yx+RQo85F+2Nb/cSY4pm0azDjAwD61h0xggzkvKAkjIrhYSkrhtQj8J9l
QoSgdKXzdwD5wftsdr1G+iUy1KcgUEUaGiaxzfMam3tBqJQmeFjKOD/3LiCWNr0+
9SDhC7CXXJ3xPW2KQiUslksFE6UIxgSopM2yvTsRkDw/9zuqR8OIrAtLhIzLIDiD
Tz/2rtiXDeY8JQ9W8/onMJRCfAnTJEliVPsKiXd9Q127+GPtDjfU/KXjxu3ixpQ3
FvhJFjHMLkMF2jd/dgQzFKLO+ep2mqRG6m7zqBMvB+4oCvUcft6qO0/YlrCG/1rY
piZ82WVsAJu3CW87J0uYtyLrGS7r7J0Qtio0il9elY2hJ+ISU4sf1rknmUkivzjH
qrvIbx0wXondSQHNMhx8ucG5QoFvm8eC5j0CdSrVSR2nOe00pPdpLbHYabMctu04
8qpidhjW+P3DOXTEh898giSVBbGNDOBGhiNVAarDhjsXarzeazIVXDMLPRo3dgZH
pGzu92jo/9aEaH9OQr+stnZZ883flLv9xklMBqDnKcy7WgU2J/JZq8VYorSHHLzG
1tPxm5nHYaUtbqKv868aVCI640NCaH9kFAuFzij2SWlgwMddF4YdnwkwOsK/p3pa
5fbIEVvykVC4KKIcq3J0LGIsd3vz25bp/2vmjs0e6d/BPgy1d9+OTDE/sJ0FcKo3
CC+iSnPY4JpA1pnho/PFbwjFVL/M++xXIrYQIR2xIP/9T9TUI2nE19cu0/IdpP59
DggvFkws1sSwZrXtUQdzUPtfODthVLDKGBbnxGCXdYzMjGQEcJr34NN8NdlxeWMQ
Bcufg9dC9+HrRPGuxM4+CN8XqqUTJAkBJQzP/Wv/K4KzwwCJNDwI4pZxgX5mbPMo
H7qb4PDrxiOaHDdKArWjM+IYuSSACR6f+7SUUKbG/Ba6GgGLjJI6nM4YPYkyERZY
`protect END_PROTECTED
