`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naFBbhVML5gMpTrr2eB5cUH4MepXmW4ZacCzM4aksLSGpkSdOH35xR3AMdInNsV7
9plUy5+Z73jcHdm9ssqwvtLGW/j5vV6AIidDIH3ISz4H7Zyl28JgqODFd6hWPVGi
kjrr8xTDucXhhXki0sR8QZHzWcGoBlzWsMiox8OHouk982T0uyBriN99mMpHDmpi
+Sz2+iFuFqJbIb8q9jQEbDMXB1TeGhdg9FlrDEeh3prcEwhLmTDcnfES4jZR8Ab7
QwfGIk8a1MQEdB9Or0HkfQ==
`protect END_PROTECTED
