`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YaFOS0xillk653RhpVjLlg8pLLniCDkyfxQgMnl6RZLyY3/SOVgj89OL7bh7FSoh
A/WwvG7q7g14AbStSNtSlFyI9QNccqYquAFc/NkYlgIUy4B/KqNhILKhfvU9Kg3w
ysg5zUtRZKf4ssQmZPpi7zgcXJph2kda2+62PPenub5kSZuZKqKICxtiYFrQvVNM
/hWiYgixkIl4kurq0COsqInv9+Tk3HqcwDAQCHV1vKfvh3n/XsJugm4E6DngK70R
CXiX5jeOtIqHkJ91uVOh8k3JyAXqD9SNrSPU2oLnsATGCxCfmN/pcDjFUbvXmlFM
O4ad6bumjiq16/azaXA/Lv5wOV+2BVfqMBTmFQdCad3yNtZxSXwm5A/RCcBzErmU
5mgNIEpUSoEvST+qhooHAPB2Di5jwPe3HDTwQpymcPLtlJB0TvfeAU2c9Ww/CeDN
`protect END_PROTECTED
