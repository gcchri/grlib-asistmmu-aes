`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4w1eLQf8n/waI5MPVmpieFVm+apqqvDjUzCswXF4s9kjZ7nZAlZYDUlCt73hVm9i
NN+QQl2itvTW38Pi+8pvp9KuoQzmdgm98fVy95jhIw61x4JlZg9lFSKwiytXWdVZ
KGTHveUsC60NQarnNosmmFcXRILtTzQLPjOdouvnx9DDgomAekMidsoB0AtWE21J
n6TRrAttAYIFnQYYXNeq8bVXD+Xn3amOu4NiDZEaEh6ls1iLHK51K2V/rRQr518n
uPqO6z95bG0Gw6jSBX33TVhPEP3LkB2S8ipkTO4cAb25MbD1oUXSR23fkRYC+sk3
4F4gCoyufe79MmftFzzVgkX3IDx0U7ZqCexcQN/eJwuTxpCNRNGgkPqf/HMIUM4g
8Y1i6032PdDltAtNSke0InWZ1U3X2MhaZwlYPaLNPOdr9C/M5bvT/LtnZBRtsXAh
woasEE1v6i6yjEI6CJEYuA43iIQSSii0JeUuJ3KL0U5e5F1qE8bQBVHhzQd5gXQu
YIlGAbBmxMUg7ascz/qnq0eMrAZ4FXyrUJCqvnqS6R3DCBWNmpLJ/zEkYmDBOpCf
XADZtQwRFvUf0MGsIf8zWA==
`protect END_PROTECTED
