`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vvo5ahNq900+SZpjLJmi3tkMRFaNrtN4JJgem/MatkgXapkkgGUKIdaYrLRMZADH
vzVTJ7zTIKJjc03i3amhZVOxbjRgJisyM3MZOCCM2RT+f5vIsxJejL8d/Gq//1/i
lJHMxLAKm+TNLui2aLD9aUiwMpKEWqFWVYYxGjBeTUw5KE/7kH+HsHBfL6bhbx9U
9hgtozKBxwLqcCH0dC3WiMIXL/1y6td5XGdIOjdjZpcUFVcYwY4L/hChWJJnH/tM
1jD+gdDLPJfOg8lhxvEytcwS25Kv8ZQu9jYeeKbaHEh3nyBU+mbU338voGjkw34E
HvXsvznQ4Xwlcso06Xm5ib/9M2/ndl+cGDflQpMjA8WlJMoLKVupLX1RoI7GEC6f
ZBCOGcZjIVPKwvRn31MPlxPnZ86Z4DYQAp5dSSWpLMI=
`protect END_PROTECTED
