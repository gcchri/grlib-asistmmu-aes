`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z7O8vk5ktpRJyNQEXmkWYGVIGYoMW3dmvVebr6Qi3Q4fo36mZK44nJvQd1L7zqVa
Ws2sqU+hrqsQa4rMfgVmSQQi31mVIsD2CQB7kipxCi1OpOLY8sQk6eYRPRi1oYsn
Vm7Tc5yux/9obdKVdMS/LAKXtI3EnxLr2O93hG69jZoKla5qww557osw94LCpGkH
JbZ3ML39rSZ0jy57IJI/xLyVq0F1wWBqeP9shY3ClYBvZCphAEMyINoER72yHfo8
gnj7IhIywcBj2BMs8OdVz31kzLmIt8255NBvcn97Ml50iop6CQrIO+D2Rfz2GpuK
z9857MG6gbnsvDk4a8e1ve2iwtVP8UelX8K7+AEXQWSMiCvt6dV3S3Xm/2S/9uQx
K2mQgOD2ysWyVyx0fsVfTikYFA7+uaZCAHhdrzL7ePO6qqUp6BM0dN/yj0MVs/8r
g/L8g0g9eBJ2EyxX3gn7L9ptErGNowrM6x56L3XuyP3/8fB+VAxWw9sEl8C4DqtP
U3dhgG5fZWgmp0A9UoI4t7u5tn9I/YbBIbdquUHc2pg6Ma2YZXDZH/t2z4h4Z/OG
Hg8j7reMbK89PAdphKR1O3pCp4qbExNBC/6Tqae2HAZ37oIDpLMUnq+bGR0LMieC
8Oxiu/v7SbwAb/mEdTHtoEKX8nlkGeUhIsvke6axfWgtCnfg06tESi5Ns16P5LuQ
305rr+U1XQsfrF+9H4EVpGWPb3kIXuXeDen4Tn9FV66sugHZb+KllXAtEuw9pSbJ
diIJb5qcl5ELuqHtDw7f/iJEV4WMn/rjAyhPi1xX+vhsnmHBpJi4qqf82ixMZP/t
JpogFxZsNvaPZVrXnbYjx7DYthL0n9WuHzl8OcMXoway9JqQTsMxj8HLme9EEhUs
WOQOAcPya9+/rOSKjc5YNcJhwgfWWpEEuO489Sz6WC09r2mUJILyLh3fN+VaED7a
`protect END_PROTECTED
