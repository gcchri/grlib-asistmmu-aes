`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SWr2HUFZ+gsCE/msCTDPhBH/r84Dqi1CJ5nH/a+4P7cpFNs+DRwiO0H/gYyx/jlM
s36PxAFkU0A1K5qz0kOzuiMTl5eBJxCN0Duyl3xJJ84sNWcLlk5Z3LM3+MAvm3d0
NZPiM0dU5WmqWw5P69hIT911dNtZktSwM2aXOCsrMjfHmktjlCRPWjtXm0tTb4pb
jyUmzVIa/uVuYv6JFxGXpb50JWtlQXrsgAtxVXt3b47ijrW2cA8mdGFkv3iHlene
/DIKABWP01e26vFDAaTYkiWEGmNNGxxLCvxKw20TW7TfVlhH01Zg/o/2p+ftKltd
JJmCc4IYWLCfPTy42zDTb1vith+GuPe6vYj90+8BVAsKdY/hm6zKIID7hw32jQFE
WIPUF5sn1SH4gU4kWHo0v4CQ1sd7ZyuADadAYGPQYbHU0vtstapYfrTwZdz92esh
S2IX0r+r0c9r2bjpdDcOu2D0159DFjvwfANzxmgbQoplCxo3dKoCmOooVV/OV6Nr
iEGzSh3DDM1jZrQ2PjmY0TjRT/r1RCtFW95bJ2P1n3v8RxDnV9OOUBFoDD+mqZp5
n+XdlUpqSXkHSF4YFWyu2KS1Z+Q12XVDAoHKbJ3MSzUJ4cYPNGxfLmJhmA4q6/tV
AjLjzEkUZkY6JQIYlvJhEdEp9hepQWGpgZYo75b9sBT99VdwSaG4n0qDT1nLt8ha
`protect END_PROTECTED
