`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/PmZ55DXKfaHwMLIZsjc2H9Xlik5GZ4D1xYzQwlm44hJT5Ry2NXFBO2H9NO/Z8hJ
6c8u9mVa3T5UuUteHSaDMe5Jy527SLreXlYCGaJf3wUgoMY8lssgF+jUgAaiT5og
O7j19/JZbOYXQRMCS/lRaatwuosz0cYS/d3JhZRJhlwz40ctWUfBwmfecEqc233m
TwwomZHYey/+kSlP3890lLvdOsdWyLaXCFWDM56Frg60D0ZtD3/w8J86/TAlWNIy
zK0IRGUVGSt+E2SBaFX3nUcqwCkqn4j9c1z2aCNCZSxAbKgWtUj5qlypZOFx+ja0
jbZNSU15vKlbgvZ2wLgZESWIqUMrOQMjazv+WlUNMAOnImksM7C6Kro2MKoNuTue
ceCe5FUlx4hRXpMrVEOmOA==
`protect END_PROTECTED
