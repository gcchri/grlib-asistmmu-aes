`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXc1QotqD7eGRx27uelL0JzENCFLhEU5uDmn0WYxK7ejKOkSGZQ0vAQ4HjwEUTej
pTRPWfN1PY0qxM8mZUHZfmVQWClz4/QmKBVGdsGaxEkA9ulBql4aephl4avLBj3a
GZeKoKYLZVaBGKn6R3hsUXijMdjwBRm/sE15/MXxfGmECjt1Q4fLau6Nn9vLEKXq
/UpUpRT35WOyBaPsifKIT8u/f1h1kE26lS7eWLeoG5sLc6Q4lX9C4v/9uZ6y7gzR
Aw5ZDsiTh1C+XPFuZc3wNcwY1nEtG72ibQAzGLnr6zNs3UMkhUJZVfnQlMcPB13I
sANYCmZp5AK9xPoWsri7uKgZQpJGD418BH78/0lAbb4SgDLmUPlFA5YMwKE2ewvs
Hwogr97zZABz8ejtb+Chx9h3Rbt82ZI3nb0isN8WwtPzbhNuo3pNac3koEoirtkp
RmTOrdLG2rck9jQhRT5tTVHiZDnkZW/IRxxb8BBn999reSgKBQlSB2wVwwzAdmqT
2UgGEhfpHJRb6xaVUxRThHq9+EAsg4+jpt6VVU55aBGitKpUpe5t49LjB5g/OCBW
5+JSWYgtEAcDIrS1aPK7D2n1EDr5UQe8cVtk4fqUW/PqMUlvhjWJHYDtXyoDCApG
CXKPpzVm3zo50nKBQUadT3XwnnW0ZrGPNS2m0UkT2zIwswqr1jic0qxajv5PDX4q
bJIS/kyv5wkkqXgMR2Q+ArXp+u9WMGkJ8ZDS1F7YTy6E7b2uN2d8UDg/nFxxzJlZ
I3K5ZTCz3B+r7adQplZ6qgIQXHlOFm2hrAfvfFszDIKbpPjh7ZDMabXcDeUTs1cz
b72Nrz5lxbhQ282GedJ4j/z67InceEi2SpUG9ItNeeMycwxDqm9ga1c5qIxaZr3C
nSCk5jv6OIQUreG5XkYIQgMpGzVwTLl4kdGkmtibSGgT4Mo79pMs85osYyjcqvP8
`protect END_PROTECTED
