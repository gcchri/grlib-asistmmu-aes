`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WvuPq+Mc1GEo/jbj3pKBOOv1AnoE/5pV2y/a8b+Ef/iggOp4fZtfJoIj5+I3YNZy
M2ITT3dvggKx9XaH+2vJ+VZV3tagmqR8P4HqoSU3vdu51p+4CfqTF0+xdYmBfzEw
kXpTq1XjBvsoO1zGtbsHhXZxn3cG3AmBmH+tPcHA9jhQ3ko2StFlr1wFmtSk7DSX
Zpmqn3ouj+lD0HT0xSGYMBMIQuSZO4kRIdJ1Fy4NJWQSZk6pzt28nz+3hKebS+Vn
A7I7Nx9wZ1DeESJmzoKxGRSFg8JQpOe7sj8SEqJ/asX+ZJI6nOLNo7lRIFD+A9Ub
GkErAZ/uDP1Caedld+9yKie1HTZsmHkz2iDd4YdTXpHcUy4rWM6m+WNFlr/A3a11
KepaqyEom3RL+fxoBKZ8yfR7bc2/6aYrNxKn7BbQZQw=
`protect END_PROTECTED
