`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zuaw2Ux0A4wiA+HqTK48BTJ0Bqqv6OOyXfKIzHZexNgKF1eCcur7qeTGfH6w78V
sTEZ4Cuk/RMN9AM4DBeudgPzdjU6pT/DutdBB2Ht5T59/ZbKLRT/hDkkiFhBeAwH
c0U3792mH4MFmYGojvnmFgWu6HcQRgAXnTxIAWQT5N+pHpbdYwpm16Y07eWc4Ml0
wGZgRoaywyyrX01ORSHw6SThKosN5odORuAVWCdCA+cwXOruRiuHORUrm4G2VoVx
PX6TZPjFEBiHpDLwayeS3nAwyqqyBgkSsyTd8ffUVEBNbXlWCoV5oRXrqNqKq/O+
YSLViC3liypM3fEroaRzna/bfdnpAHPtS24fXHfoSIka2kFf5js6/5zzcG5j5b+j
dNNB9uzxNI3LPZhwJY0yXqgzEV3hOENx0E0mnWgbysTGroweEax9is029K4yA1MH
C9NQVLxCVmGVg4V3/XkWPFeKgAIHHWtuou/zi8fcvabyJbU0O4CRvtn5LoeNvAgU
tMS2jqJ6Ik1YG3sEsU0pLOpOO+YfiDpbyS0JTyDSsTBu6wRXHS6eC3Z3d/eFF9N/
+Qfly4MerfCB2X3Ws/Qd/7eoAO+++iBBp4t4ObdHa30GRqxfHJ1Ab2B/+4HpFeX+
DOC/q7ZXM98mLZHUpdB9CEjoAJfIw34CPfTHE0C7VnD537yqTG4QN/VHrma56IUD
RhZSRWL6nVL/PFxfSRPXWc29MAxnXddawIjBFFUn9m6V/v42dTqx/hTHwNwFXpT1
KGFflYLEX9KBnrEeqvMC75xsQg25TWvsmW+Nt0fvtz8Nh0P3yMtbatAhsIVSIUOe
bov82HteawSt+nSObyuGeQnITvDJgTw4RKYkfHGqbqpE734HZuakvRetDeG6wg02
NXrk/wWMXpjOlox8QkgbPogZCKoa38Cmu8RLD1nLGq88MNlU0bLhoHGIvyaKBR8U
ujDRsksy6NkTJCBmN/16U8K6MaZxKw+z6WIyly0QCYgxjycWK7L24/LNE2VzI3mY
RDnzkey6vqf12YBDP+uaSO4zqhgLsFHXTT9+BUioQxqqYtrT/TZjq4QtTQbHQkA7
GBtBX6fOih8P1chGUMNWMEPfFyCRp47uOBRcyXrW+6gOaxcUXWiSxc9HBGVjjS+V
aAmRjWTfditNRTFK8rNUV/a4c8odRyKDu+i+b5dLGJnnV8K2moelp7UBY2ElDRL9
ezyKHB3oMmoniowSp7h4HKAkmOx3EnyrlV73Sp0Yz/dOZlN4gL8H5Qw8J3g+QQT3
lKPC4BmSmAvy9h1KPdhVH0Yjl8SrqEP2QiRGGclRo4QUcvzJp0nwYI1szoahO0Vn
HAJynJ3R5CshBsDHQhIcPQaCXDAccLqLfA6nx4GYEkWWUcW6Xw3HrdMKZirAUjfS
MPpH026zK6KdWHxgagzns/FJ9xo62CMBrfHV7eYUQShb+1+vmr3kP4dgC2aJrnb9
AWxftHnkNPluR5/V1D0G8yr50+xMXSQu1/FPQM94F4LubCaHkVIuDG0G62fxwiSs
VV1uh4Oik9dfS03+GTq3VBrlfpvqNBScNbU89+XUKXTEi0/FWz4V/Cp4DbSdvoAx
jPUb4aSFivGPnijqFUolw7qav1pbNYq7orfRz6nOQoyy32nigN+8Q2edAM1Q6e1t
UN0vwg+i9fE9BEIptXTh2WeiHb2CciHoMpf0NWx0PPL1xrMxjofZGjlYXrdakhrs
mLOpZUOz7MlaFAolRh0EGJAr+iYhC84KDUqod4J6MsYlu61TmcIlfigMBjxK5Ken
St+TSsYQ4tc9YQjZfij5GhtZSotBzy5W3oaoUHUP6J/edF50jzA5o/5BhJC0D4Vn
vU+FCTTyrqLDb5kr5x8haxTlWQ7bZn9Agrua6D86c4oSyCSm44JHuu0XAXxMCnyB
hUypldnS6RNrVEYhDLkWPTxu70epQi1y3UYjecppJ6URzMnFdtqUA7ynHKizj9s0
t7Q5va1X5CH7zaV9i0kHuuLOWHiAbAjCpSm4WV95+Xk7BKBQYXHiUVSbLRKGjpgr
ealWoZ1nF7EOXUPcS7smbVYhqpJARr/TjXbD6lbrQKsksOuHdgG23BHmXBG3v+Ue
gFDCxiU+S3TTWxQemxhPh7I/l+fZce24qVJwa4/uS4wGvcC5VZ6XmpN6C5UQunur
TnH3KHqQJfeoYkTr7MeJ4HMNP1H5P/jfPw6zuX5qps/6oTaUBAoTZw6nBQ6tndjr
6oHC8C89EUAKtTYtx3PPvbJaZEZOJl5I0nFld55+Bx+SEJWrkW17qhQr3aK880Ez
REXSBq3QaTi6t60PboBzWUoRe9e0Q+YieipUNGp/Bz3oO39Evz6hbhkYI+cwj/2G
KnS1d2UnLmdY8rsRExzGWL5I0mmljXyH0YFoos4hgX8HMX9RSYXzNDRD9aFN1SBo
yQ4PiYxjfnBklQ4vB6wAjv0mP0an3nf7VydrnJ7h5H8VNsZdt29uuDICOVOPIdWF
1QBdmOypstbP17HEu99lfzaai1471mRQKx82VVnqf54xYb7TbJfg3PgCCpFg6Vt4
LEc7mMciQuMtCHLqGah+uXx1+KeG4IHex7JN/AohqxgKe4wxJwyEcQ8d6iYcxHBi
xcEUGyEEHBsXSg4HcPWwkgorddW+6v+nBWJda8AwPM6rCEoKxD076DgFCMUpSZwn
eYpkTjclXeInsK6wBD1Teeee+KbNcdPm40w3JNfpOP1FeW9iphQbnhvWT1RAMRXH
exaN6h+EeGzzSu/Tfgk8UV6+2JlQ2upsRHpg6m5qSACW4N03iTBOGD0mLmwMQqGI
8McacYFPL/Gl4Q4tTo0eERietMb4+CIKnqGy947oX7R+zLUaBtGrQGZyU1tvQnBo
XnEra3DGlQKeyk1u6PcAHGRK0dD/PcfLtd6qTtGdmpnMXVR4CnI2DoZCZ/i9WhMt
nkR8Lasl/ALGJRU+Y6/vGnfxoArOGx3ePzI8oz4/TDGSjT8BYKiGLFEddhPIwZqA
xREhLfzxE+WUwXeOCPWV2SKA0H9NOjNQ8s+Iu4TYRF6zHxSmpRGDkALu8cI67zjQ
w6D5IoJxg51OzqOk7oFzT2cfnfq+wJvZUCICmRgXtbpHjbMNA66ED0G5blGaeeEC
2HMHLwSAS+212Wcvf1RTgfwONul1wwekIUrZZhXFwXoXtjxvjsBQU70bIweWefMC
jwSUqg5lDx13Juq2sqDjFVFHX7Ff87FeE/P5eAaXY7A7zp62sFfrGnOOUsOC3q6U
YPoOk7xkO3qa7qQCxRHHbOkgj0gVuqHBvN0GpliLWeuunoNCTW2DdCoxWr71Uazg
x+sn0mnSopTnhJcY3cDD8o4NNyN9zsQuhS+x42pmfu2nUHU/l8UKtRcPrN+dMqeX
SWHyGQ+TnORzpOw1lDW4xu+6IghKzyV6Q8Neo5Bi4LkEXde22zDZ4olMflY6x0fQ
MvXFDbsnVArhojHnAbg0XVSKdL3iq/sLw9B5sT61kKsXew8gv9VcQrLGvLvgBxhS
li7dxcgfHE112ap7I+pYUqh9tXmxg2H/l1eGtPLXQAaANFzpHgqy3SipKBu0N9GS
R5C4IXtomQRtN/4S++FK/6LCBFOzDr/bQxH90exSiAWYearMXDKYfR6VldHt1Ce7
zafBeAGx7eVR2v+VetBDDwQCbITSArTh/OtOuoHRoLuNy4tblzi8dR3TCAI6J04Q
YV56lKYQ7aQ6uyd55o/yaUd0HAvhK/zUlD8vOBGT5uYGlFRB+xW7UxXwi4fzAfDh
9bkTDsRLkJx95Pp3VUW5grWaSdkm5y5e0g1u87qMtsKqELSAVCcNWeDlOzti446J
2CPCcG8TFc81B5u1A5cP5GafRRzhI9d9NAOfdtB46lIh054Gms0mPiHUmTFdhMk+
DQJJ3SvL7ofe5s/6FuatdbuL2r4W1WCv9NkJI3v7Oezwng4MBw9xLNzjVZ3OIY0N
IdELl9H4U6VV5WTOIVRM9QasnFAplg38w7fvggq3a/8pbnv4MR1jevJicDq4RIxX
/EvUD+ZNCz0xDrVxGAbDoVUZrNJfMT7KkmGs1vox0gGEkA6UqyxxgYNLGBMSN5p8
/b3uGC5o4QY8sZFPjd/u04qiO4rzSJwvdxV1uWkKnmjbK0XRx8ndgacEXd1xkJXC
nVOIfEhenHmyvWvWNymaqELHl8BIjFvVj+aD58Cxi8CNIkSARJjc4y5+2AnFYoK4
yzNsr3y9TQBVFZBkwHbos61iYfFa6fGNMiYLPAUkvRz6tAnoavFh0fJ98Fn/LQww
wCLflBoRpPBjDSfyXGS6X/eRQibNgzxMXn1lHghCzux8vvgOL2nnavaUzUXMidEE
BE1oR0vrsn7HZk4NBeWf1sEwpADfbDD+qAYeh6gmNcvUDtLRA4EiwM7G6o1/6B2I
z+BvIP4Si14Nog8rM4BBosng81b8/6ywv3luSXHg1v2DLdJxr/AIRTv91xhON6Nw
lUlxyBKWq2MfMWy/d7jXO1DtEatY7mXLBt9hbmVs7vgocnZg9yhyuOGPh8ADshOz
s7FGCHQ7BVwJUhDNSZ+7v0r2yQoV6YV4yoreROyoowFsYBKtYMEs9B9K/xRty5wZ
GYPy0H7cA5HOewXcZKODo2PTvculULyU8kjA2pXLA5Vv1Y/pw7FidJYUG6p6I55t
BuxX4JZySRS80sp0CjL50XkZO+QTHEVYZoXb40HkC4jTAzAo0RbWm2eAEpBjSp4H
OUJezh2W7sx0+vLQx778bOCAcb3ZU7w+ySPjBf1ZgRh4S5QWQrIfu6F2RHZkk4O0
PH5dH2TuZpEn0VdcCx4UH8ptFexhUdWN4z3nXYgN9MItflvTk+VgAm9DbM+nQe3J
VeM6l0K/D1RGw1x/Xx5t/anC4OP9d3oBlQWzFqu65Ui3mkpSn8e1lbiG7KzgVRXu
r/1Y7ydxkA2Ne6sJcn9k6l5PiMBY0wvJvq5WDw+qv4/lzWYqUlAoLN9TB7uuEOl5
BH6K3GHFjmcRetGFvSkL5odUc1ujyYxoCT2PTztY26Ps7YdUFqLod6YUQGNyQjkB
QfZ7xc9wgsfJLcZj3TifAw6oo1+qHUlLxfcz8pR90JDLQCnWMpxS3ivWWNbXgr5+
QcqeqXN47GRoYa2JIxr7TRWRyf1zG6NhbVW5uEXB97eUZDVYRTLd3uHVlGiio6+2
LV/yZkmCzjH0q3nncSb0IRV4uLWkMMXjoqi5dSTBWSwoiOG8XlyJZECcuDbz9hdA
J2OqBKhGDEnE81MxFZnq8HnmOHh7ajBbjIfJIryRHMpIU2gD4l/IRaZ4SwxCGNWA
pVlWw+KRzsRXQ/vXQxAkzVnhLz0OwzZolZngJZNy6bzF8lWF06ErOvxLT0kMynPd
sW5DI2txXUIe9xHK2DavBx4/7aoIdwoVnYtUB1OveFYFQbE/lVRQ9fIFlaFgDBZk
4UBKPHWdE/Hv9j/1OmdqLt0lZqKY0VgTz08HMYt5xTxk4I7Ndmnf0eVAVk4qN4fs
i5nx1gY1WwG9OT236iJTtu+QybGk8m7ZSNAQzcegAD2YFUaETRfkHTWPY9fNoQjA
wuY3EGdS+LxOjDqsT0fXFmr8neBVCsmGRPoryRqniiVb+m+qzPuHmk4kGPI+Li0/
LB/huiKB8JkW8gO/qiHxC1O9hoygPrHqKzshbLQoJJ9AG6imdqzp4T/e7JBAy4G7
Z/vDH8u6MprgFmcGvGhjtZimvGDuIr0Cy+RactAW20x3lCH9njM8nt1+L9Zok2aF
1dsMT71wktTmV5UpHYd98m4b6q5LMPqOgiA84yVGOVM89ECzrEKVOFck0Wa0Lbwl
QBGi7XOHwz1EXo2SrSUR3J5xjuhI3q3Q5IfytwqCu4VFw7YujfV1+xDFwpM0+zbj
LAvvZjwGnyMbOXVU7laL0S58XsBiCCXWscSTNw0oBxuIBWK1QtmDvTegXpoOsBNk
g5ZvUNS56XOdWHlHXCyjKbMtDkZ2EMJ9bKSL7WMnIcjeewlN4gTz4aYfDsTIopdJ
lQCmt4Gg2XABbNOVXJlOK3DjLsocffbgH/woBA2hUqfJZVLh7wcCMPLKbzkQQf7v
irSvBjtrB3pNoDtX0rjWHDhQklUE2oCU4y2w/mjJeK9aHydbINTBPrSYoLZC+4CX
Dt8Ue5pE/VEbPrAz19nobfoV1rbLLpUT2LTO3DyvJFY5BNXqTNKe3V6ts44hZrY1
XS74y1obAaZhMcJgXG67AqPpoDUahIwTsnI4sTHLAJmaZsbRdHRpsn4JGPBh7+rs
N8oQS0soH+8l6L6I3Lz5G2wIUf6o+5JkmBwwDwWveuAf2jpvD1WkEL9w/y2hrCQK
eIBtykU3+8c8UYpiEbxb/HUx0BI4rEHrcLxkUFbXSIQ76gH4iQApUR8FWgXaI/9p
SPN9TOjX50FLznw0as4e9WGWq5hTxhj9AH5AMH8UfliCxPmATq7ABIdfPgcl51Lk
8BWjJaSYcb3lh4LWZ4iJwyan994FkZba6ty54lKTLqycWBNlp4FkBVglNdJDCeld
L/lnLUQLiciu/KA6WzHBZWMqktrgW5vL8ff4ISfy7AMmnR98nNCQK0wNGBtDLnc/
IyW+BiJocb7Njt3+KhkMA/iWVs0+zmQ6utkqu3Q5KlbGOC59Q1I2fAZWSDlnYPlG
D35xeusHqCSnPP0wvXcMQ5tZf0h8stHB7+qr3AQhJ2NtmzsoyPoz0AOmj+0Y1Gp1
Umn6PoDuez3uaA+GkI/vPC6d6fg+EmZBR1RIR4jXJqQFMixvtTzKH0M6In6qx5CN
jWf5lC4IPN7MU7W3VPhm92rgFEIQ/Nxt2DS0vCzRbCAv6y8nfHRerOl+TxN9gxiF
KNUUqGMzVSO+yBH+SFnQue6MqfDhMk/M6mIagqMZaA1b8TDbTBICHMuIP6JgTs36
ItmCpGJraQtPUYjEuYpJC3yio637CyoFxXU0ztrIc2hA3HAjlDN1gn10I+zjGpsv
xGry7/La9AjUAu2NCxHaJccTTXTsDDtRF2xleOD05uN3CEr6QVBg7Ciu4AUwc94i
k37JCJVzf+PiYoDMI3ZZZVVuXncxTEdqE98LzE23YrHRYCt/sXonj+V4vrCr7Nh/
P01k/oXYYiptbnZNqW3Kg+FZvzOKFRnw1YHjPL21se5Mw03DlL6u2OoriUyrng8k
fwweyoc5+KHWI7uOFhgu418QjwBIV444oz6seSoGzj1QYlXAzcK0xSku8pUEovno
MjA05rW3nrEGnpBo2fK9WYRSnB8cz/9y2RCd0TJnHdunMuSM7ZAd5MV3ix6Qaw2U
0ToDfM98vFGZEZzHTB4o3KJuXQn/a7NjtB/0t4jmI1XaTvJfd7iYPoODGgV8OXxA
9hdKZ8FvMQzwPaXuUGI5rX62LvvwJ1B8rkqO3rUyNwoPcORdXKwVURkghYk6XEqp
n8eksSGt7yq2kU54r/p00AxATsw+LbnIYrJq735m41HU9y25Y7fvWquDzf/WVCBi
sqf0pY2GEV4v8eXUR5hQWCyC09hc29saqOlL8XIsKIB84Mld3LZJ3W31tyy1UKey
HLhWTFXL4dqTMKHI9BFKkcBexbvqSmlI/I0MHdFl8YsYLB+oqz9zpInWw/nCX4p5
dilziajP08S+U9rnyxE/AUJcMpLjuKU+aFg40wtqp0XzCIMZ58N0rBPG/FugOEPL
BLKMMO5xrE7wl1OHhTujBu6FLt8lCwI4MZ1Op+Hr38D72Cmg7mOG929FtI5cnNvj
VeEEhOANg5URJTmwxk2JxRsmRXuy6qaFadUUSM0audeWqFSEO3ah/LLlFlAUsyGq
Z8FEbF4lKHOE2RVWCTIAhCOSfUKvutwzColNJM67j8rLahX3PUvXEOdQXHyIKI1i
PXJSMEFmVsrhgYWm9X2EbNt6/tq8eoai4kLpCtBfJKh5YjvITRp+rewGnXNEFxM6
wWcwzAGSPHSO0u9lDDgolUxP3lW8mR19Tyg/IusGgGJTd5dCxOQHgqLpDgrO6NDW
NeKZcQUTbW2k4TBpe3O1E/gPMOL4kMsVZWIDgZHcld/sbOJsDpFwS3MJbhDyLI/D
5xvDZ0RS+iITSBsIHzhaa/ZM23Y18spVDBchYhvwwTKvZjbZ+UPEiVg1lTOj23i1
W7E+GR1M6BiQQsO6AtH4BAyioA5NES5AVMtOaIprOlcAx5Bac5U6ikaT0+0TFrvM
+fAag72gqAlW26v2H/GRzqbP7ZPA9dbzt+NBuLeh2Y6HDVOdnIsCEabTCd4R5fMN
u/x8nDQgIe4xex5T8rs+UYr+rXCkBNBe5q6+Eu8HsEJjryFfHyLapY1Kg5gNZPpB
9ip24cHAatM2CuUBsT/fwmGfzuP1sSgESPnpNKCsJljSJwEkPqEAmBj078NczAbq
UTGRdxzG/j1UE8BgnYPYtouXwE9xroXPuJjgbkiKYuwOD5ClGETEjuqJUPJjgTZL
442wUU6iHRC53dNvbwQnaBMqlWKDcQjjbSoLKjxEcpqAkHmh1MonkkiXep03shxc
nK0oEv9H3Cqb6Jfhr+gu9aSwR2/19y7BX1bwnBxbc/bf0c/SlKF8iP2uTTP8wFcX
Fh+hmVmBMY3rsI6VmzdGsjxhQxkx3kv6rF5An9H8goFksasq9tkOoAYznkWHBOir
FmHJTNmi7dV6gqqY10Q5Gg03rkObREK4lUWA6nF82NYv94ovxsSQDjOWymIuFH5d
jrce5U3iJB/RVbBRm4dK8Ntgn1CV68dWYsCURRSHLr349p2m22rgAAK6rmM03d6x
aLrPxPAkzkE+2lc9FnFqxZZlIX7U2rwvEdfwbNzmDojHRF8rQZ+vyoUdjgyml37G
dxgrXEPdasQLba7T0SQQKpeJYD/EF0eHok05KiP1ViBj/brt3fD8hPVnWYFfVf7A
uGR0d7n2zouXxM+JfovSCPurVVmIIDlPoRrhptBmN/OrG96I0QRErYmIZ+Yg1O3q
wHtlcgJQw4LwyyZvZBT6I6sn8uY4BUf1X5QbBznN4cMDid1VRzklP2lX6RLx564h
M8xyUTs9TjFlxIBnIlHhvF52hUmcPFiyLrbIg2Ss+4eVQ03IpSoVgdFbaU/gWJXa
+k/fIE8XywQ4yMbzciG9urwhRGW7z9i3CF+ypNUgiRnLV8vQJl1PSrGjJKeJcYVa
1rH9NgdyvwWBnXQxFa/kvuqkluiME+Xjbi1uz8Huu43rjDvsTK8lNO8LCFUW8qQS
N4sqio+GihKCqr0m4on+Ne/hHSn+TB6XOxdiMnaJNlDkIXIFehCDekx+0EKCae9R
KgWT5SXtXdnJSk+OMmdmYWlEUqB/EoKeSiZSOQmDoVJAgs+T5W5EbCyw4+awyCwv
tiLw/t7yIOeYP++osYEtmA==
`protect END_PROTECTED
