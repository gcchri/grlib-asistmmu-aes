`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jU3aYZKGGhAoyjKrFmUbQ8UlStPDHiCTzJXOMFYbuzeGbsIr8hUAi76DIHitSCNi
l+15Z4ghDK3g9vJIxE3mgcNfL/lQVAZDBbW6qozSMe3u/ycqyjSNYNmAfSTN5ji/
j58trHoIkrXB1JmZnaNqgrGCKoL4ef2ytabMfRnk3VE+3GFaGCpaKGiLtSXUOAEU
6bXT5xHS1ge2z5nCAkDS8ZklmTSQgw2330vvDVV4oyXvwVtCkZyyjDwD2Kz1l7EA
kCv+vyCTlCsyCJ9YzTPEEYkWwiYSyMJFcZw735WEmebzYXD6sl8vPqswKN05dSUu
TGqsjuKR1+chz90yyE6UpkL4zp5MMUvigUIi3563qZyoWm/SFjADl0fetI7dFB/7
qTFiqOnSz0Vag56uUPwhF08Oo1wGWKXEuOlwxSrKaRg=
`protect END_PROTECTED
