`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rA1almkzi8KHx0IiCfknBU9s4v8VQkY8ieBpomxzE2mfR15CyWidcbX0Gunlyctc
kA9TXMG0nWkAQM48QfE8xKH7Kt+OwiObw6pVXrucAODxoEDBLnZjm3iFFEQgYFvB
oI0iscwyZe4Hk04XUCO2OownKJ40jy1gvtsEF291INsvYEshj7hnmJSNLmuYxzsm
Ofpn2NlmYZsuIFPAqzbDne8LLUOWGkqwPXZa1tCAtjb42YfusTpdA+d6KLJUhlMc
8MjgcFt7VdrmhjrBsfCqv20gkXQGYalWBT69783FJEyVzRNbVCcYWzDiEOjvYfJh
Zr56F0vuvS954m4gBicQB+Xv6cZijsUEotbqsTfsBtuGYY+1ODDd9NU+z1SLFUHF
oiYZDvYaysTyyMMNYprIfsezlWE2mT/e5PdcVBB9UKwFq4iPVA/reXO0yFoqNz0w
2msT9ULfreEzFGUQGAoR6rNBo5AQYNTgP/LrzCQpQVvMJNQHzvdJGK7UpP0Q31aP
dxPzZHb6hQhwCZKQkxxm4GbHEi1/97WJuYHii8YzAFstyxuITRzpzmPR6grKHj0K
OUkyHxn7ycFHP2+yFmZuJF1TpLbeElmMXvjHf8jsK1ET7nuag9ZBp9btsw374XJP
bQBGgyEpL9J648O/A1Gxb+xoN2JGIkdusAfsuWvLqvKyUjMtndxoNSCJZkBj7HoD
w0eynWV+glwiuqq+xyefteiTAD6mIr0bIojNsLKDk50cZ2axCYyxl/0S0l5ARHaY
vWbEFO4qjnkGEGarkVxZB1yFQDYrHjJt01NlFYmbC0fkecrhNVwnshlropV2a9gO
K05ysne6YFYkFtH2Fr8He19fEhBBvJ7qV0J9f1c9Vn8s/1OmD/VA0Sdi/xl5H+63
vIn6ltotaAQfqMAxijYksA4R+WE3KQdWgoQhHGzPzRm7G+yedOYvWf0S17eWBYtL
Q116/e5LKSQyzV0bz0+DgYmUCEKdlGh1dWKsQ7tExqRUyY1lpXN0bxV/pXb1q6OP
q9LjcLXsHIgLWjDWsrcJdOUgrTJxJVfQ9a+/xpWjDXLB0hMSiL6p7vbhqf4a86ID
xTKFca4/AfHc4FZ41x4uvfd2zEr3+dblU4cUi/otEeQy2JKnTRJczoyErK3iRNI8
NOkya4EsCMub84RGUBFSGXZs6FRU246mNsA5fUQaMzKnMsZLN6XZzJK8msHdWyqh
4DwP/IIFiT9W+pvjwEI5q8IxMRWeZMF3t6iEHorAbMa07D3ZnmJv8AoHAR+S8Dr4
E3RWQ7dPOaHRXsCp6A7kewNct3Wn0DibQV6JIJYxpo36raLmapd+LhxOQDm77K6V
B84sosxUl0DINrCTrBPVjoR1OY6nlzQEBk0VgHw1ioRhuTZl0+xTzdBnL76KRzA2
hscJMqc7Bd2rUgoAY4/I4WC2JTMMMrRx5OO+dT8iQtzi7hJHu1rOjFFQTFmvpgVn
v3p19ab9A7oHcyOHkGjPlqz+21Fah0uOqxNDPvyq2HAGdslcPIpAsntbpHIRSWpE
tkBcGxPg/3OiUHkneSTqAKUVlOQnjo7HG6V29Txj2/K6yjYRbYjCDvnqf6dvHfTe
`protect END_PROTECTED
