`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1XMlxEJC8VlWyk4Y6tZKjnU6tL0sTjAVLqXg4HhApcDKKd/9oSIrCJzK/qQuC9a
lFsVzBnGdiWi11ma7b9K5yhnHX0ZaFndWw5gtKI7+me++X7hMw4cooVYXdANBHXL
z1QyQkjLM1Rh2dj/Zazjs5VeBnGcFvgN7wAbPLwApoGBK9CewoQA9eGPP/Xp9Na4
A5y/7izkrtouqGhrhYoCXWkwHGLNAKQ5OLBCtIYCzKB+/lDCS7kqj1sNxPw+mUVi
eoeu9IkUS0aEAji2UEUenImc08W3wjigxM7SP5ifucUaz2br+DN3uqbC3davCGUW
xbeKIN+hBeG1Q7/Od35FVOCb1acDwtHovi+Ynno2qwMei/9U4uvL0bKyuO0xeO4D
XGqGL+8MIw4Urgop9uLjWa1V3V9FYyxAKE2GVXoI/QPXcz5l5vSon8RWIYUAgEbB
BER8YjiF6aMUDbouSmAUgquDlJeWIAA4vzCa1W0i+yXc1kpk18euU+tS5NH7gx4k
O7kRTiOZr+527sRbgrcdvxz2fbZvpH7+kfgNFMzNr+NslHwoLGzfDIQH8OtG3/1k
OXSr5yUckZYZhfX/d/RsyvcyvR6yjjCPLqSrv3GeQRk=
`protect END_PROTECTED
