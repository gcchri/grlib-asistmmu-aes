`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jCskmuW76VOt10kw2Dk9Ctz1rMjzpz9rCB0hVQ8YpOmO1FvVqZwU+RgL9sN2XjKF
VHtEcYqCxVlHOtkfTDrHokbgoHu0KZM258w+Yq5dKQE37viDEOuDCGb3oMR2eTK4
17Jf+xuBAC1nce4tB7JvBLCaS77uKRVyFAzN8DoUsQimNAhR+0hVDyHoZ+4VEbYA
dkZjOMMu247StVDb4P5V6PjhQN16/CdDQN5ltAW27NWcdZkyzmbI5VazYQLGxcka
EholKHfAqe9H93jKhs1CdVM+Qb6h5FzMzkTR8wkORvTcApuxR+No3sAn85RFw781
BIGWFhqQUyKB+BJSKKKdSpDQI44nBzI+Oqgye+/30GPBWDNWF9/NT2Ibs224x2tI
zdygozqBLymvQh7L4T/kQuIPoQnL3PCugAy4t5m3qRPkgiKVI2w6RyEOBry1riQh
`protect END_PROTECTED
