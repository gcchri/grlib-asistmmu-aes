`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fp2PSRtcVnWrVpV/Zd+UKx89XHEZSoMYOeIGkAyFK9cNz3Il7OU1ADEDuqVIxXZJ
N13lIuRHIDIb7Oe0aSWTVw6E1C55GiyFopLJYvZqmC1U+2HaQhGXIi0j6OElLEp0
gkuBXhEQ1+MTxdRW4jr/iPf4nqTOzEwQrO57tX0IN4k+9F8g6EBUat5J2cCVLR/e
ge6Ll7h1TsZyT8a72ltwWgqF465DDFixMBqh3u+ncNJypZ5f1LJ0pd6VB+izBVyD
LNllmdG00DLynyar5CVYs+gZjThYvLFXizs8fySqczreX75x29+tTSJUvk6Fmso2
HN63cVoKIy656yoIbHrqm/oPnU4e+k5192f1K8red6OSu/7fWSYzl+jSyDYCShod
8qtklS/oXaqsfp1CyTH6d7GyOYf5atJLrVAqCvWsksYMNcMUe2qTahR/wfpOPaC2
y70kPxRFY/y8Y2ZADBohPAq03OiGCQ4K1RwasM4RMbVdS9CODNlDT/hM7SRYMX2J
z1d1kgll+Lp1EX7Og8xYhKzM9vflQr4h5tTaeZxhyG2dMqYPe6GnaKn6nKA7uZjf
sCFCDN0xZoCrJJpZMjawRlBVe29LI5anjgJiz0tDPKf+5x3yPdo7imF9A9nS+vKE
VGFXfc7RS7gYB/VHW2aIQA==
`protect END_PROTECTED
