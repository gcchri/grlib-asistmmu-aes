`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y7FxTcOnLkkO6qGIoAP7ooGknjJOH3vG2kwhkMtZMFxvn592KvMVxz8cSNLKkpU5
+KiDCCmN/eeWj3v/wYxvJIKZ89P12wpo8dB9hX7frBT0XBdH9a6I1H+MVGVc0J9F
ZnGyIBQmlN2fLKaJ7ZsFs8L8ElikhJlbP82j8uG33IeQYhQ/PZ+Xpk3ripm/vgYT
Gv8h4TDoOTNdEN9SQs8BuBorA2g1qKrxhE68BRcCeQpjZzG1XjJI3cZwHbybdoJ7
hrZrbVoPYeFZPgx6HuV/FfSkG+vIoV25VpSF0+im9B8+9zm/eFrRhxG2sOsht2M0
w53r0ttYDnYuoKD0VOeLB4HGds4Y7OFWvzPG/lqP54O562unCiKOdLNnwgYrp2/r
/3rNo1kTa2bvdqaIPN2MkpM10dn0SMRlolK6ucvTESQHT3HjsWqZlWlpsd2ZBtqW
x7KPgCYhXu1d7rcUihbsoX3AcuowZru1606wZSej+mP9340ECG7UEFXGsojLKP7g
4rcSwMc1wBn9CSGmYSLIuVYqI0KgPJz9KXvxU6yEzU3qwCG0h87Pd66N91lJpXsB
nbPUuXMuz8UioRvDtg8sj7IqGosEgUoigIqRlsKeJ/uXyHyKOz2rCgUT+NXY8cnO
pYWbr+WjZPPd5JXisiwK2XdvSpKu/5DnprSByufiaKxm3952uNQPuzwXu2QF6F3p
WOn97UAxaZ8E09uI/tBlcERkeI43DzlmDvS+xWSWQ4tjq3KHv6yf7cyn/GkwKB+E
qWxyYOJxihp5YkmnOjVqq/LKlTExig6iedH2C8pimW2UpfkvFAEimIAACutZhFIF
5FkcXIbokclydazRazSn9Q9j4ZfWzTtaCrmZvepQq65leTfTiZ/JEk587qpUZWam
hv6WfGDIspfy/oJpLiCHofc8DaeN53PyetJGJ6IQ/CYt44rAmMXcIN7Wq7My94lP
`protect END_PROTECTED
