`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sLL/J04lEFSs9s4qaqYqkIN3JwJMYJb6BxvVIom+/utP0acsRLlANqzKjRDdvaps
SK6VgiqfSRVvfI/8Gk83QAdxvsY3d0Tv4uXzG3tej4ppFZBycX5oNuCligaXVI1M
uPZAZko3YeuOY4jxfkDbvq1YY2xGD0NXSXWJCmU4DWwhth9sJgKeqkI3CTDZpRbS
ZJpLakiPeQ2dA3qKmivU83M6cqvyfOVv/nbY8NdwuKTb3Wyqrr+OAbOAEo+h08S+
Nvh1/iRrqZGjYfoUehAVFvZIRITFtf8C0Tn3gt5XOqY=
`protect END_PROTECTED
