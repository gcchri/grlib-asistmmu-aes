`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9i3zjSGpgBo/1uN0lcBtCjmm7F6M8pKVLif2QfL+KyAMZE8jM11OS4R3K3zOqw+
jmseEK8NA4qr6w7krh4j1oSqlDr796hWPjRFUoZm+I1CSihs801OosFBc+ALs4Eh
Mv8Z0RYxjv5818ztsOgluHkHubsPwjXpQlozOyjhk9AeytbSDZ4ucF+mn4qzQ0Zo
Um/ccTSVNO+20wY4y0d8YNhWFsqzrU1k8wPQYzX2MYDTTvDYtHlP1UzLVYmxuWEU
bQQhqTzakOWmV71cgrukO0n0oIHLVzo9fd9XR5c2Fz0jz9zz215LgxOW4q8jXndd
LCIUIroiLFvpkkxEM1Z6v/Jlsxlhqa9Bavob+NmUS4skLQNOTN+4tzmebh5Q4t/H
6TiAixptSxtPhEvxep8KRHs/RXiNFCrdV7o7acjPNvE=
`protect END_PROTECTED
