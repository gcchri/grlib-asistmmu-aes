`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BJbmpp1gMvr5bxQubK583luRsW7XPh/YRNyeBH9NER9G6pTsLX/YQ2KcKDNQY1OB
5jOrJ6/fCFoqCzAO0YeyIaUv9LzvZ0Xx+ThNGULjPkWQHJVeH8ApWIubX+KQLuPA
1iL9dUZBQwusOloDgIkLD8P99+Y7KBex1EkAXpAooZ298jDJIJ2HYURgCdaBtf3U
BXdnxwRtdoF7etldIVuxeQd53BM9JvgDHO+W1YwjLIdJjzlh3flWCM0TV3ZvDg7K
NV9z++nQrYmFD8bEiNSd9q7pDybQovgrppvczBot6OGLHwDKgpnyiXQ7m5UccOUQ
pEUeI0dxgW2FJg9kMQdFoiTeE/GraQCTb3+uICzLPkCr4u/szEwIN38XkPnFcNmo
pSVMZfbnmd3qSXiMGi9ZLXV1GEnOitbBjZEuckOqtnAdt2F7mIqrCloR7JV0m9o4
DxJUOyEyO3OOedIHNzF3bFVfMph/oz9T09/GxQfwYDYk86MbR0fcrXdiktSMMCz9
knAH67p2e6bAxU4TXCKRRFxOGE6fIkcmIsrjMGuODwfHA5hw1p2BIaw1fngB391M
FsrvlbJ3GQC+QVczcZYjI5XG707dI/0zi9gMVXzxDwBfARJAYslZplDs2pufjaM+
sKeNuaO0yjJQLLuHt7PdK0tFjwRGdv7PdgbDYySqVB/wxKIVo3H4fVjoBRfI8abk
+pXr3wqtDOM1MMWbwZQiMRtSj3fxk63bfVuq9wLa/xmZJQikif5ob9mbxKkyPRmu
M2D7pPkJiBpV5QtGd14pxenHUZhc58WmOZGmZQ6NXOlImwKUfBX2vr5XOd1vjqQm
WBk4YGigLrrbVrkK8N3b9BHrdp1COD7VY4PdaC03gHhSmlm/OcHbaMyiX94NnWSH
B2t/x57hGpw3wVDS/uQ8vsJA9AfbGJscssQvS7fLIS0l6x7FocT8HUEy8i71CY/N
42LbxtfN1/B/QfZC4jbeRkeGptpD5IIlYO3L9R4i3NxSXMUr5D+LhqVPf9+1WRvz
/Y97/3ivWn1KqE91CFPUArhunfLdsqRYWkj7VTeXZxo5Kh9fcyBng3JY02m2I7WF
GxHoynk5a5zsOMK91YKJURhlrhe+vOV20cGkjwh2a05lGQRGEIpYNpsP11Usp0Vu
f99Ccxo/asn5ObOJSquzbTkJHj2VI763M4Ss3aIaIKLSkbr41N8MnHJcR2A+p2n5
LsYdjjO+53gssHWS3450+tdpwFod/hgCjCzqLMhlp35cJT5xBwvKtWKv1j3KgesL
jTiSbz1zvkoqGrGJuX5/23CahojMiUF2M4swqfFv6KvLsMsc7kVzn82knent8x+m
3gqSRqL0XAJgS39ohaCo3PObO4zvJ0/6stKufKhxXzKmn0rTtuD2yFo+PEm8Cb5r
OLlpwjWzr6f4YoTmeMxW5iTfHq+zW0xNqoGkEbu4rynmERyGD+DjHol3uYzU6BpX
QPsF5Y7AAxMH7CPmQBx2G3CZn4vuXOQTErOtEJ1TiUn2D/YoB6vEa8xDd/Adpzbz
ULLfCkevAonU3RDz4eBU7+bt5hMuou1GnH+2UAG9FBpktujzJxets+2IyFJ+WXnl
CG2apLuyMW4oCNVxclyzq1S+xmF8wXuXu1bomNrVsUU2fQx033yhnZpJD8j4Zfyd
7zyjI5novg+Rs/CMegpuTPhdt670q94P9tqwhpb2BVWvmRv95DF/CA9MgUFPxV/o
mq/GqR1kqtn0uEalkEjVNARDe89meajPwxGTF3MqzW72Z8FjzLZYibBddeG+X2jg
XOlUiGF4uDR2I/qMGOP4AEgUtiWPLiW9u6oU1rZZhJfBvQDhZ1awHUDp+codPUqK
YvJjeDPyaKvX+5FuCEKTBNM7yhZKszhqdXGqgC7ttVQhZ2ioaYwH4VmSdeCNXaTX
4lf+7CLpOzHXyletx9mXTIjMFAVhr5FLCh057+vbErYNP1aUczohqOHQlwJ9KOQC
ygdcd0T3QGFW3VQn97RRDIIwir/hPhOJ2JLpV6tTorGvgDHPlpW9dEO7Ud54fLPm
R8fEtO9XrODphbuyRGYMSCdDwuvtXc86P5IDM8/QtRqpYK3L3U3rzakBbSNa1lMy
DFTGJ4o883+ri8jR9WdVcWAMBkDwzVuUVtXpe8oiWD2+oeDyCXXfURGsjvd500yI
3s2q1h6IhyI4bKuzPavz2w4nvO0gD9+5YF75tApf9vtUJ/N658+zsCfyQL17N6nb
HlBeO5r2drLnfCpFGFv7qUqGy+Rn0l0zeaAfjjyJNOVc4Hb/z5iCKDyjuL7YlJkc
9tLDCaTVSa2DrbsmHpKAqLOQDOrCct0QhFgWOOGOUy234tyr43OdUG9XI4vrMrXA
xa62wq68Je0S3ZUfVfxNdDUm4WBU2IWM2bIp9OvpT5nDqupjstyyseEMYd7CS3LY
bbIhgMlCSpZtaIeEjyKGeje0oRXtZiHNrYBKNl16bGwHF/1i4vQjLFB8nOFJ2MYr
x4n0PhtN+4/9kzu/hFiQLcT+Rt5qEBmo7IznN+cY6p8JLjsEJLy55w5O0JcBJ5uY
kJcn05wKb1tOxOmHxYBATM0WMmJ/HeD96wgCIP7QaX7W2/6J20MwyZMsktYkOrcT
/I+GmP2CYZAH2OJ6N2w8GDVC4befxy5x68s3vU1N/uln+vtZo+6M97xFm66LgSEZ
1a4irZNO8kEq1hn4Lcppv+Q5HU+ZxavZMYjSBmoLvlPgCeKDY0UVNtglSt0Ys8Ic
Da0lIw4bqBscwasNOu4ccZrt91YsxnH7l+Sm3pLlGVK490YXy7uh1R/ZupRTT4BW
zLGGqSHnJlMHlg2KbVap66QcYqtX7aEvGKJ0HDUtFI+y2cM4swOzOMJzcty1t3Bg
juQOg0prDoo1GWhzyV310SD12MDQZyJs5vZMzym4ugCBbpX5MvTERpBeOepM3bnu
m0XM+zP25wvThIr68pxJAxMS12B974zTyOZ199OCfFL9Gv2OzSxRUvCjI2j9+amr
P25pc3Rzy0YjHvk2fuB64AoaZFsKdGuH+zH3Sd9KJi1XBsMN/MZbtG1K0d2oZXB/
4i8paUICwMBL3bSNr4YnrUREyC1OCq7kQ9AeFTZOy9RMbuHEKKZEQpLfbVuSNHBb
0ityR6bVETOIX4g60lsVQpPwcnyn6nnEfdI5IJQ1t/4PxpNprl/HqzDJ2FiBpFXy
r1zXjxVgw5jl95/WGfwFzBLr2BEQ8eITP5n6yR+esak8U2aIbPpL3nDuwGUx/Dun
ZnkmB+GEcPH1F4oFPDBK3fDpHTl13ae0hpCv5e4HotDUXlggc80ZI1/LPXwhnXcS
ej6xj4GbEr3IX7moNYrOORnEx439+UcLR8IsSQ5Ob3RPLJtBsDHmJM/MDQnARHtS
uZ3zSeeGYra7vAh9SsT71idStdw4/hTYdGT7YmWAKkr6j38gW4DZfEYPy+k0SApk
gZwocJuMZmTP+9qfBm2CbfQqmbjfJb44Bfav/U1OahH7WVriiFDUJ0CtnOU0iGqO
3DTq9eWaj7rQvNzH5vXiMoeaVqVXlQ8N5pU1BbCyv8jmkKASBquj6kRVDZY3LFSI
ot9hprFLh0zPq1qd5K1pFld+G5JRIr+1SrGaxlc/0a4Jcp1tsPk14/VnNnlGklKX
BXPmRFmg1IvbkTFQ5kmPTKRGXHAUOh50umhy4bpm5JIU4OS1Li5967Abu5oiqK/r
4LLZd5ala+CHNuyOFHTLBWjDLJ+eqo3sA7uaUgm+bhoIJJNRT/jatn4N1Lp1VPYR
d8z8x30tEdhlu7bH0XJf6H6fYfz+ozIy8nTPQpq/t437J6ip1/TP1gX1awJZdpwV
CDUQCgRQgx+rk29fJ6or4RprvbMevpFoEPkiU1M4A3h1HMz1paF3cmeiqZr/NETd
GFSwhVLPlCy15sixBZeZZxU4fRBfIuVNWDLUMrkw+1pbnHhpUJIERpL41RRSxha7
6Zu4nEbxdYo0jBW4RvUiuSJ+zS/J8AA0LYf3os2AX5zyWDi+GktU5jP0/iqVPhLI
QE+P2wImhPUymT6xPaXsla0AJwmCrD3FH0akUtuKCnebaLXxIntEjbK4mRTB8WhY
iWVGRDmpQAPuRozGzRSHyeHMSPDtJoLPj9DuPFHmdTZvsBGUbrKIq7epLY42PDxa
jyMnCZzphUTyV48wIVtY9lFMuOSqsBmwp9VlL+ZZQUnJQnzJganf6hUMokTwH0xv
vlPp4EuHCIa8GsB16Y4jqQlqz49tpI8u9fU9RpStRQH1BCWikTphdgUFszBuRoC0
46E92q6xPKclhI6iUiV+I/lMVGNWtqJdZN2Q2dVCedIpviH+YtI3wDeIq+e/sU+Z
NybM6Ytb69jJKGVqappyjigUwfhLYzfaualz9Oz1xmxrnm82t3o9MrwbmQczNmDy
99RI9U86O7rb5J+YKGkqGWmfKf2FF3xCdmyxBGGmz7hi3q21VmDVtzcSx8yW1o/N
UfFIiGkgZhIDYkJBzdT8I+0prWWZJm96rUuWn58xBQiK3sWJGcpmpVYVAIisSNow
ma0VWlosq1UpPOoBjn6U1RIt/15E+XJS/MODaiUfVwSa3yNiAm7QR1mhrChYSCHU
vOavOm12xWpcFS3UqBNTWTybWsqftuGEUXnMWW8QCzYQnwB0yIT6z+4qtZI4eFWv
E7wAw1psuYokj4KyzoYSP8IDMm4HldBaOCj1/UQO3MGDIiuKulmBODsVw1FyMdKn
VIsj+Neuk4/I7uMzktAAC0vu6uxtoGGI+whgihuph4yYUv4YV+YY/ScLqMcSCD+z
GlfOfsvIx/AZN2tkkblw4DCGCoLQqEI7nzXYbc+wo2pmvg9qVAmiw22hWoMEH1Us
wAj15+Mxl5Vv8aJ+O/wXl1XBYvKWIUOcNI7G6RrKJkGhECH/iCAa6khy7u5y2L14
AUVkjf2lD2P1fiEtanU0RVYQpKXLwMveOhDxsfIvg5MZn1frRjXnMYEW7oXC5QZq
aytSoxig293j0sTahmPXkjGiDCm+9dJ78BxzdNZgc78hK90vPfObh0nkVb8d1SoS
6gxipWiZYiUS2fEWh2ud3Geywnf89DM8PLAitZHzB7u5nCumZCM87Kk15ZPlGJD4
7pZ3QMMV3nfmNZt9HdyipOxHt3hrKQjcfuO8XkzCfwSZWxKYbDzRo4xRuDbM1jKQ
x+Lo/6JjxiRjNXihTft7SWWsTafJa3mphdFqUY19f7r0NWmUk8I1ZDSdKywgk+ct
Al0ZB0Zl1v4afChp3Ent3y3JZvrxXSptyARraUz4j//tX00d6w9rb6DiW6UBT03Y
K5zidzVGVnsg7jhNNfre32chKP8ktIBPdpLQhZZP6rgBz2J5IFnJMz2yGyM9sqWo
+UjMIckeCQH2rJMeNgYwFaTLjKk3u2h25VMvIPm4zVs/z/uad862daVoYuw+Enqv
`protect END_PROTECTED
