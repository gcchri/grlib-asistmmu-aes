`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
odYYq6IswQABNzTdNbQlgccfrPWyLH8S5Sx5hp4nmWyj+ap2vYnLRl8EIJcklZGz
cOTPabI2bLVRKkZ0zmJ0ef5fqZ1WdHYsVcs5HRI+ZCwXBl4sDg15GsrTujpiW0Z4
dOlXTjI8cF6hKeDphOOdOS7efsQuTN1AKEqKfrbVcuDQXMm1ShoqCQp7ctQyKjs4
LQvjrf19TIuO7I4pAM88Cg==
`protect END_PROTECTED
