`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+jJgJzCwiFD10mPi47L00WEMeeQLOz3nyCm38dyzBiaVr9gTwoQ7xHTOGZnkqYY
F/cUb2hIf+s2GmSTc8xTeEeHCB3amjLJqktyr22PJbl9MTwxlycwRxIZepaiStkM
dKWcQYnLncw8saBoEdWGog20O3ap9tFrim2/PCxzK2ZVaRLodFZeZN9dHLPrUGsN
LtWw1PkUYcmvrXYSfym/pW+kQ2M8DBz4OnuIQbhsZu+FrVPXjYj1TCE0NSu/t7y8
ex8ep2buGse4OZcdLcRyiWpEfiPH4LsmWtfKKvP9j1J8dIq2NMfT1UDVoKopFRN8
NpS1rjyfJfQlTfJg7zZt6Kh3JHXQ3gLzu9U0GSekYkoLYthg3vp8eGHGQ5p6iEqQ
2egz6Q5h5h9L09AbFqyQWXjODuaRfZ/5JX3XPPPcNyTewTCTXSoE/9HD8LyC0Vjd
I3bTNnFhAYuGEbnR9PR1R9fW5Gy4FGXg2SCHRn64MGLdsGvrMAKM/Qndaim6LH5c
`protect END_PROTECTED
