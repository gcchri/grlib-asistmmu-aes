`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulwN71RrFuhgrPQSruTgIuD9hGW6ZjKlK+TeR5IvMv77Vf4JUR2ZlnMdKkdQEhNo
Z3QqEck4UDS6JEV6VMa47Dkgdo+FGWsGtfkMo44A71HQQs/jmMR+KH5MRBojVpcy
qvq4p+4GuzgAJgLnwLq4p3Tkr/ixvmOaugYmyPY2bcvwPWqjzr8UcAoqNJAy9ZN5
O9ikTE0N3V9rCKmSGAO0w9SKhW133eJWLehQZHo+QyhOmAVpWMFCOSMiHf2Ubp1E
x4B9YmSiN2VDde7tOeg/zsar8STCulJofq+Pqb3ay27ShrcUkTOoXr01nXSXdYuW
PCwVxTcVwhdo5XIbqZTCdydROptG900x9x/2bARXx+8FiJe8IxotvCWOBfhSKeRr
nIliDKYKyjAEfBEl4RvE0EO1PDHkK81DIHeuLxibHxeRI4P4e4Oeugfg7tA5uL9T
Q4vt/FRuMaomnElVF+JsuSe0h1fWHWgB6lGUOaZO75YTND57MlB1LecnjDfFitJo
e3SieeCPNty2FhCa2xFbZgAOP6s8dwl9LITwWZyUjRknFsYJWToT1SUV54n0Tzh8
86JCnflI30Beak4tRF5PB04xmV8LbIH0/EXsN23yp4wPYUAj30V17fX8QYSmqD1+
27DrpRhkaVCzpF3J82Wx5HQBvHvV5mX4q2qkxJf6Qrh6Jtv97YjQuBqs9wIEy4VD
1CyVfuElizO7nX3dcxPUFchiA9IMmUOWNYXMVSulsEYM+I2/dqLsgDlPC8mCMd0l
`protect END_PROTECTED
