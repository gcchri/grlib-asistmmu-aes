`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ADfur7yXC469W7E/pnOfu69meKQac1QwR4KfJbnxELyJF13Qnal53si+3ZjHXYUR
zkQATuE74PxLmaBIqTycK+2gixr2MTYKw4/TpQuMXwpuVVkIGpDaSqNpH9AB1OcV
1Z+epO4nrnrMS/IrnH8aEBFPAO1neF+C/sE5cOpUO12qb/IZbS0K0QGRnP+19Ajz
CT07RWZYFIq2W70ms3EU/XRro6daAqs8VADct3uW8RAYZPaRa1u7n3Yjh9yWzUtd
t7i6t85qZkjvvm96HxgCmZt/3WoFilyjn0BrQyGmUbuA5pPAiKCj2/XRnfDjaM9G
H5fhAjn8Ka/zLUr2nVpYqavscPG6Tupuajo4QvhhJhEY2EERg1v7Ll3YDB9YCwyf
rsEC793ZVoBprbwF9GLpkWDekTfFjbt9trvlvFtn4mnDANdhjqFQLgji0sbIkuo6
N3utsv0NJbOKs6bwR65I/N1XnHJlLdnSfPbuljhz+Zg=
`protect END_PROTECTED
