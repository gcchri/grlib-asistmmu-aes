`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFH28ZDMVnx8jbNhPCK1TO++bdD31ygsttL5x5j9yx/T2w/OniuG6DUk9T7NIedy
bzJl0ZQcvvEx1CIPyDAJMdV0tLK27P3y/McdX3KSIP2MPOSWk42GzESckWaxzZj8
y+7odBYcVqRqqErqkNj9DGgz1gfAfLeAJfl5vm0YAm/DM1dHaD9zk0QQUJwQcN6F
CW0LXwedOLq0rhjN8eDru8QB8ZpWIdVbxs5J5goDiRH8aS32n+ftJe0FsNkqeNM7
AUwy8+x/VAWjcJJaZMLZzl0PO8l0/qQ4prNwmP1erjFW/e2Sr5odsV2wCkHUgjuf
Bt0kKnsTkrjyupPEPbWS07Tm/QSV8tZqe2a4qbAgoQJOgrd3IWYX2oTJF1W1rLmb
BFDDRa3KSaKfx0WVRog/tfKUBIo7fcVdD7wjAFfVM0Y6Q+Tv4MdkoVjkk5rJ+wQx
Q3XsQhUD21qckwaDqAhNgFDus819X5vDKQ1t6SSv1oh4RRPleteV6YOecCvBjCV+
`protect END_PROTECTED
