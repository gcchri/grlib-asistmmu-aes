`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvQHeZqhkMd0oC9TNm62XdiwFO0Zb25V87J2q68e8BEZE1ZJudr86A/1pMgwcoZi
wHSlWyG95yi2D57nIL7qEkjPuwOaT9N7WzfbtXrCla41O3hpU/MzuVfPJRBFJs/x
vBUvDKWDxjOnrSmg7AdlmPUni+ixrpmn89K3RF7u6b5oTktfXDcqeCm5A1HhBDSs
PNSuJNf8YIX4gvapx30lVE3iuYCm0AbEt3CQG63JWWY/Onk6sz96P/R1rKhKIV8K
8X/upeJJEYlli4Q1M9tXk7CWclc+vgGiWLjX6WQ7dleFSGegd6yk3H2bh9ZMTFPN
wZ3tgAMG/8zsqt/qFvWyRCEXh0q89NTvpRe6MZOE+OSMzQ4woanGLGVqDdTVTQmt
saqDh3HuJh008p8Pkwf59P3rpBfBeLxuqkwdnf2iXZU=
`protect END_PROTECTED
