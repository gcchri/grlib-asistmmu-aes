`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UM8tQKi4l6u8Rc7P4uUpDx+YWBtzSBptUVgbboZWuXIqJkz52wLfEyuwDKVI9mph
fhoZK5wYRxBx4NNKC5qOPHbVAlk/E7LgiWGY1IKkMd2zshrySe39a9+b7VpFWu7w
B3i0GTG8F0OC2hJPoHIW2yZ7j3TL2yDqwj6HB5E3nunzQ8remq+2ntBnDk/70L8u
8jg4QsOvwkZeWSS6QHfPcYXF4wt3FzTY61MrzJL6VNpEBlPqdweJqa8WBuoKblRA
`protect END_PROTECTED
