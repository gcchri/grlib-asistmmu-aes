`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LHEryxbh4sTNipm3+N3NeNLXn6t4stlbM/3KSSau3vwfHo6cA+ZJYUSP8bumi/3+
FncVWUWkQM392+bSZ421hZZZl998Dwdoa9bnYZ5kIRC2LM38OVrUd3Q6RjpwMoBb
tI9iuJ41pK3Z9MgK9S390YUmeuSa0wNgxciDm/5o2GPUdSrf1JpxeAjveTcMbUR4
fbgqvoU06f+NaKywN977UpA5dacVSeYh+YMFv3U8m+/Ocrai3UejcvLZCT5JC8Av
RH6nPU6neA2fUduMAI1xZNst0G9uTv6PsN2iTiNm3AFcQMv8x3L1wVv+R2/HD0ZQ
bVK8IXjIcaQGkp7K7dWstrw37y4KQeo8y7jm7YbTz45q161aZqzc760JHBDKkLSS
b1BaP69hhzjNhgRS8Eb6f9DICg8I5+8PxwlyGePr60ndtK/6Q1yhZRNN3+NIH9ga
4hH+Bb9wn6F2dZRJKevp+0FEeUviaoxcGAjZ2JZx0BIV9daocTL1JGhrXXtSfH14
upwoYl6QuPGpBtpC9VDfbCTs0KOUg8o7XdZ5IEypyj4oIardQsKCT+Zjc9e5jjb4
igev3davxq5HUfwAPacPoR+wL+M5bCmyxf9konrWWFk=
`protect END_PROTECTED
