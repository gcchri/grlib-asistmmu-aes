`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Of8YKl3kezfmreFx9oqiWq+BCHhKSWjfyei7+O4RiC2l6ZR1+izD2L+okMJMj1J4
oi05DNLODsXtLaZ7ck/pD1OPx1NUM5BIUzlJqrYrr3v2PdDXViZBdnddBYHSIYj1
3VauL6R9H5kB8t8qqZcphHzVUfQgS8jv9cvpWgCaGHCEOXg8ct/5kcuVkUZQxgxP
4p6kZmVWeb4Oj+/xW/TMb/cKotZsiIjqFRcN6O+RVgxJt7PBY0qYjzusT8qp709C
PXX97vMiWp+tuvfnu3Dp2kD/NEQxJnziX2VCToouWxIIOtiAOlnRxZbKMbhk4+Ic
gVZxYgp0Fa8LtjEKK8G0pmd3H8gYrsJ3vQW+hBUb4gmgiH6dBOgWlkZoeCYCGZB5
UQ5q3zkCpog/tvqbI6ZBPA==
`protect END_PROTECTED
