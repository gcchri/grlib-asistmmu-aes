`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S6AsxUNX8ffIhgLEDCeUvLggZUJjlP9g9oteaxtbyLCBR6kASiU65bltbBDntqGw
UyidVl1VeKdPsr2pbp2Hwuf8678eDKNzjEDe3SmMr0Nh1P5miuX+epzRL166IpfP
TH6lTG45tYQCszv6ct0xBVq5roavTxxZ5S2JO4KC/7n9uO6SaL7KiHg3hV9gIAFk
Dn8i3GX8SKodilSWbWkqrjm8uFcIYJVLAOX2H1hoLtJf0isew/ErVv+uHRkesJgy
KbN0q0bx+bwZKxjsF5XNXosQt5uKTAqzwB1S29ZbCozqf2fO7ZX8Popgh+xrkZw4
wKs16eOOoTxeC/FdIGS8IdIGMOrQkC9cgIfDRvfFqh8PTvwyI/t96V1Bnu5Lqzqw
ARqY8wcncpvvSpJF56OLcWfnheH2UWXH2rfN/WMY2gklpS6hRCwcZTiFb0AZwj9v
ylCZ09VHzmwhCNTH6LL0hOLnO/GLIqClb62ppey+tAGCC47lByeEY2Aya0/rJ36K
fVokgx9v8kzT+f2VlzImeY9uQk8IUcAmTIh3kQMxU0tT20ZgvK+kggGmeD6MhQha
mzLWcvdC2yeg9khh6Ith8cNqUdBz+d8oFbMlkgkcWSwX4Ez4zW6/1sAodyF6KPOj
`protect END_PROTECTED
