`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJ8quLY/EwJxL77CjGg/OALKMj/MaAH2ar5zcxRppmXy4XjcnuOkvUGmhaGvMIDM
6BOJS2PyvcQWIo/5LXHmdf9PYf88T8pfjNcTS4OIEU0XK1pDyqOR3OjP/lS4uiq+
rah4g4levTzaBuAsQcs9WVsZzrUrbMlPZHsccLQj7chsN+zxJ6gSfUka1Ny2tyeD
M87IQS1IHrVIS3eqq6X9ncrUyfc1amkLNXeual0mE0DZNkvv0JUF6YZ2rEsrkfF4
m85OaIdf79YQnW0vOwECQWo5p1YQf86vyM9RpDZFmFo2QPD4QPCqm6ilKADXcZ4u
nQrMjd1/A6r/ie4U2uW35r57ujanTe1W/BHDxn0htG43zs5i/xxYpy001j6cT+VS
jHi7OKTruYDsVjzbcknsaw==
`protect END_PROTECTED
