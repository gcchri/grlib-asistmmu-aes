`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZY7dwu5YGREsSfndhp1767GoscciU7d4wMrBJ1FkMe86/xzi7O43K0VxBu3cRnX
UOEbXpuaY7fP6Q5qhZbeDAXTbCFwJxzo44H0hCZvSsiLURAKDs3bghaeN2lz2GbX
6SAUT9DiOVWHF+7/f2ASJ2Q6Pfh03v4hmcIq4ewfSVdbLNrca90iRAU6+6JB/bxS
aT+s6hSMDsBjuwg8dBrdc6LvfeNxV1swyyqmbW2CCNCzQMaU2rHz8X+dqwKF3fe4
NL5/07Ic2VS0OU7Vo0M3g1bJVSNCUbAphwTTASvAP24Pkc/s3gLOO6vtTWCumPX2
k5LQ7mmKw7pIhzcTSNhaL03n+GGclUuGhsT4ifCYkIw/7VcWx6A/YiFzeISZNSbI
Z9PY6V0uWfeWMNOQRDoLIMDI3kLtvU9I1BTlKagOwZjsnISTZbUpcTn4DyaRu4cR
dr5fn2QVcq+z3iy8T8AvsseG81HRygFAhTfs1ovegMmUQ+paLjZS+EHLQKrIqkhN
rbuMn1/drUeQTwICvhl3/FEWyjPaOs5fYiphFNPEo7/ADZ74UiQbOq5QbGXIfHqq
iqlSz1F7VlI4jubRSWB0kWfGGI8WKuBLMIEZoLeQrUVMW79u0cyNJv3cZQIOToRJ
hP0rGu4bVfnBsow92DPBRXPQSWVbYKqwQleP0b9Liy70jrU4iVj8oQrCq/kf8zGv
SHiKzPvKDeXxRJVUWZeay67/5FOo4Rq9qgA5iveWd/friotqzuLp38YY17WyvKn1
lZY5q4kDlt0/J6JJMtYLWw1IFVsKdJYGPRUZNFgD5iNj5LHYzvcBBoBH9yIiX5uM
k1PyLPNdfa1VE96iHaesP8gGMq+E7kEuHMmvdfd4u5TSpJoL4C+M8JX4QTx6IJ7q
AJJM85ajsjsSit0znpJvvF+AnwXqDjRJd/NEi6U+bmc4c1ciJfbfM3w0Xzh2VExM
am3ipGnvlxjnbAukoy2UQIoGqna+Qy29Mb5Z9lGVra+NZIrioC0l2cyXv8OdD3NM
JynBd2pqRqSO0C/nJjnnstl7BFBLkIXMLf4SP9ooNRPBBAi1aLuUnTXJH9+GwnpV
dGCLaJ7TV2nIMvBtp4xCB5C43wya5mGFaSI+vtMKy2LoZ8e2kculRmuvQlYwuf0D
MyCqfjHARCh7a4ayZBQhTnCOPMP4hehh07Qgzjr9NNJxA0nJVCcKrYkxEQXccbrG
bLhn+RjdD5aYaZMGP2PQwVmIBv3j2kfxBVkq2aecOrY=
`protect END_PROTECTED
