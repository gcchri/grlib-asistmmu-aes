`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6pZRc4Md23BCk9WLd31qWYFrXnB3JYIu8r4AyMP4TZCcVuXcfDSnZ7XcMwX3bRl
wodwD/7v3DQ1FX7ojpA2lyLiALgwfBHVJXVklVeGtBFACEyrXKioND+XwvBUKM0O
G1s9ZoI/XOY7UrxziKVE0CR+qrEbcNbeRCoGhwbPMDf64OgA2qGkjdddH8kOEXA0
IXtkNu78/CSbPL31/QN8Orx3HWcNUeLAA6imNVehi1gPYHrr7A96rnzhI/5LOuB5
xplkkxb9y/kWJYiVigEacS4pxOTBKsBsBTPI1aYFGCyRaIyuuXQLnmxrncn8gOZ/
K9lWrbioIjpAOaFS8+61gD7yM0GFDNP0dpIgKOucJw037zn8hWPArU0X1XuSoTD3
j3TGB4SkRjcFl93CmfCqCrNIiZNCh6Qprpxn1cgFdKFQ5Rj221cQqYu7lLAAeIkJ
f+4Z51zCY5GqoSuADQAl2co/mx1oBlSyfrCI30aVp4igdhv2rfAD65M61mzwerdE
`protect END_PROTECTED
