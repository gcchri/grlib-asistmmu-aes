`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bDLkSNPonrTDutrK0UH5M5DyMc27cL+4HDopm7p9ijCr3nkE9M3SmFgCPka8xs1Y
LpQ5jrUe5FIm+ihcwGWlvPukDn2Cglu4p28YMpFaWwrCpAv6RSMQveL4f3g3rT7F
bzkYhuOFhDrpt6puWjl4xf278iYJNHyzOc0TsxN/suQsqPgyvMF4i+woPRiEppjT
RVsiDpJFmLU0ptRfSXszyPh98wq+mEaGjAumtFdbgUwZBXYWbHa2OJyM8lqD7bkp
9n703+rbdqEeW53bjOti2p0+bpexn4/T9d9ied+AlaEKyh8otb7b71vAR9nAxPPp
i/H2/OBPHmtC3So0idz/SEZxykmc5evORVnKGeA+ZOh9qGCGv/av0X7pGv03G0dl
3l1lumYzH18M2rfsW/7em6yQqfJqqvur+wazCNCtq4wC6eqY9M8rBzXTZeDeJovx
jaEEzFsN1yYg3gRA9cG595lHLUNEMq8E6hIbp/6wyJWPKJ80JuLysOczja0Lqaqg
xMV2RL1rDWckXlBn4Z5N6w==
`protect END_PROTECTED
