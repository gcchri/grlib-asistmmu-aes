`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDX7C93QzUL6ti/sIla6kdNLerYz1ND+oDie+8EBQ3srAH1IRNOEXZ3wl9j4nHxJ
DMKAc6+w0Wjkw0VxKTXNARTrcWeGmwmC1OK4f9tmZHMARbha0/UP952Wgk9whHen
+giQ19Z0qwjLNkwoZgwGgMHMS6ANUNXkEjwOAicWB2aRtfZWmJVobGVKWUIL8J/A
+AbZaVtAK8bsNgUIAIC3f5gJb2pHtxrnd4TM5X/TqtQk2EEVYtVktQP7kXaPL9aG
dVzRSbBSjMntVFT1WYzNqVwKX+XHOfoJ/ZZHcXn9A1zPNv6RRnM/yv0NdWhuFvUH
kfJDMthxgxIu4Cek+mfJHpfXNS7245PgiZMB07R+yoymbtc/Virlz4tneoK6qIRH
rJcNmdLsLXugS6qFe8BWh2XoCsYI8vFgYbJcDt7fyv/hVAy5YUCGOrxMv+B7eI97
LweaE6LmVycRiqwE9MwVN/JtCte8tG2zZRRJUeF3xb7uxx52u/EE/EQg/M8ebTCt
zc5orGAQPAmPCeHlp55M1d9bTZwu2pf5EVHL+qAieeqwB7CJzo5ouNXVlm03J3OU
6Obvy19oTa5Np1oWDMERjw==
`protect END_PROTECTED
