`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
br1xiv3cnxaoTN/hb1jYGqGCrVRAShCMK4l2i2fkbugaz1dQps6lb3xqZGVXmx47
TlXD0HZ4/hUPp02WWLcxajcj/fldpY7BY3VCJZg1E5UCD40YpZVnKxZ0zTHImatN
2bRbgB1AuTJrCqxM1Z6yx3K+UoPVsZfzixpqiME4R+gapQKEFltwRsbXE68g3Y6c
d0JFDCrNKg91Qv5WGMINnscbJEJ4+LfuorOUTBNAVA2JudzIE3/57gnfhONIJ5Cj
`protect END_PROTECTED
