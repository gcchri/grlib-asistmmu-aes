`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvYUiNYexj8rwQXf4VShabThU0nFL1Ylfb2Uel3GH/tigIJn371+ZEKnbW6Zc6Iy
juiBQ7qVoO2Xd4heZ6wSiql8xUf7aMEgs1q8QdlylJg/dMvDnTVWYSvf/fiFQMkw
pvjh0M6YoUz41ABkr4QO6KeiSQAb88CCgcqNvqleMhu8nf+77SrGXxMWeF+4nKcJ
yAcQ9U1tJOW1HyoOK1sBAG03axSEyPfOwLuuoGPfljZkNV0/GkYaW0GmXQZbZHAI
4yzxEEYKgiEYaSg10aCEAJIEcJfkIQNoCxjksUtVLIzntBF8KhOVrbO/GKWFawev
WUSgMi9p8kvA46OwmOW45wN2cpuHEzDrOtx9QcgwX7RAM1PuPgQxlGXMSpECYIJl
Yq7w3iYcJ6eYT06P8m/8SJI/tkEG/3FV4MZz2KPvoALEfHVZ6xEBnACwsLik+98X
X/yJPHeRSJEDOqLyT7OROXJRzUWhqlidkpyQzoiQ6sRUTZ7Npw0X9kVj5qRhFDWd
3hCzOq8exCNBTaasSe9iBsjcU193yMdXLEYbkwGHyAh3TdTzpjeCt/7rOHzkKllK
R5dmOLyaNyq+f800f7LRTwuVJ3CGvJ7RFqn5iqwwFWrKMlvM46gX1KVYEbKmY3Of
jEQ15NQdvAv0LnTl7/gQC8LnuWZlJ3CUmqmhoCrAFBo=
`protect END_PROTECTED
