`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTMXHtZR6A1Sbmd0jXxAgaEmrlsPHr4kHlC2uGoc85kAK2I5LijTSiaV5/SrUSKH
TIOk2DZPOg9NUBoi6u3mbznxrz/mL1V3NQ+4dlP4mmPjuB7VXbHOPLw+/M3ABV1f
yyLycvTF3+SErta3fWIsmNmpZuxztnuIgDVo1xFzChdYNRomz5MX8V4FG0yICYdo
1m2U/kxcFhBXK/eBpx3TZnOQVBIe+rzSdsQ9ya+CY/Nmq4L8fsrN4Xp4664tXY5O
RBsNYml1Q89AjIPeI3aX40ff+U+emienBg2pel1VkggDU395+AwfLUGgoyFPGO4b
qq4IUeUyAsjpkeEbdWzAzOLHD+RyeyAmO2aPYL/J/R1YpDZTPbniiIS0Y83SBwRr
nsnNCU2ciAWCvYoYsDYEPXFozTYQdsIOuPd0uBZDvNn+JQYMnr57/pZn2GhoBbYg
`protect END_PROTECTED
