`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PG672YkYHoUqoFHDYuCzYz4P5Aj9Qd/gceju0d6ZQ87a+QQ15DKK6Nj9QDBWr3v
lSyyQujT7ptKgYcS7D9vtLXhJke7W3veo1bgTEWEdQAj7NS8gIbLNEippRbqmQ7b
8SaCLztCgcGNlsiIz0xvtT23COHrCIv0WpiTkTMf0N9fT2mRWhHKKBFVVHleZFcX
BLb2QoaPfTUqXmMJ6w5NajblbaLF5O7UZ7WJWcbEIApM5vEa1KVVyrfD+9WCq3Qq
UIbhelG6RDZIRhet03lOhtDtF01q5wflei3WHicxco8zlAWLAnTwVS9VRHgAPmwR
/SzfcpKyLNcDBw4W+QsIj0jpv6gY72CbFCd4GqeIvqS4itKP0AT84DQYHNC/gqlH
oIVs/BehDOzsVUR9Picg41/W4uC3xBQlREyKXMnYYaHzBDWLRDszpiG89gqpGjww
HtNFk5IB/wUIrYAzN2kceIt1yR1YUdTyvCgsI0GTgVpkuvJNs55vYsrO8Gb96Ild
yCecIwf+9xRFCHNyPjHdW8KOzQ5M6ciqESoy8XlvVAvmIn1z6Ix7cKSSkVe4bQXR
BNovq3YniU+ylKrUb42iImnP9jNsJc7LgNRTDwQDeHa1ys4iJ2SWtzae0EWcGfB/
6be6OVvbGF7BusFTIRXVoxKs7qPpe7BrPm3duAr5KoqI/BddgwmifQe1QxoYsK0T
vWGvUIR83ihmX/BpxlgAyyKS1oxZAsuIkeLzJ9cAz3e2Yo/F5b4KrChxXeAloSrz
6/c1wxlBq+IVoT9nq3OT9Z+96qqc1kQaa1UtCnhC6MIZbommHBaZ/lIbC43aZuTO
Z3q2G0uKkF1ZXEMak7mbAWu1uHA0l3SDygP/jjPCGnvfrgItMJ+V3e1x2/NrxROD
j6+9RxmwnihwurHxkUNBkaySIsYtR+i9QXOhphGCrZYaib9hHfnFVooGniacwZBR
+gyrEowt6kA4LUMRnuTNQDKuvq5hb69H5vIRDh89RM7FF7AqeM+XLWOBxQt29vt0
4nRUK5l0+awKefZJbQmOs/EhXGDVpvJDwAKcr/jUe4QMEe/w9ApMqb6S07aPO5vU
CC8s3KyAgXLgRt/QJJBmjH4b3ssYImk670c2zms1lDIcBAgJed9mvjoDIi/LqwPT
HGo7IM5OlPnvGP/J8niewqR+8p0Gvlk9/4n+YvMCsG7LNZkgM0jyTxfXpuCUfizG
KV1S4rMJGvIzv4n8aTEEXQwI70fkF0fiH7xmLIORsvInkoKONxEhqMe/F9qlKGkJ
dOrkQub8exugab5NTXr50BTiklhpdnwViAe1hf7fsQIWmfjraJ/40alGgJdUbtlF
+ZnQP3SgNIJtRq9DVw+nU1FH9dU9QY+9VwphBcE+7ryKjI6ux4SXvWZ77oI/ExNI
1t9EmTNi4YiqLVdUApwq1vozvvQV56r5j/Mj3HJ9JF3BEaRsKCeDkg/DGXQLvgwC
kWSob0s+qSI7K/4JsgoslFXV0J5kzWdlEaI3Lx943Fk4BbhgSBXInpjNimYKzB1K
rKhXRrIhomDXMsZd/QoOF9OFnpnksVuLNADlPWiG9bESrae9x1aYNOjcOj1pP3/V
1p76salO4KFEEShKzQ5S7Jp5BW44184OiYZu3w9F5poOIaONoGDVCtTOhtnbzc7F
oAEhvs/2Olz8EuLpi7OA9AwsQC3WnGgRhOeqd3lLS1Q/08ufuzn8A8zlaonjQ8+3
ihK7GekDvatSIIjIB2PmJ0TzLXflgGeptsFTJxQVEvIJKMTJwOW8c4ru7CyDRTiU
2s2Pfrfcw2TLc8P63dS3bqQpmVG92Hn2WXmEsoN7Ra+OZvAJ9ZgwbVU4j5cnFt1U
ttA5GC1T6P7ZYfFc2n1KGmWhGJOkfFU2/lU1LCVRAqoOdHNPff0gxeHM59nUP51J
fFRmwLN/9hR7rn2azpkK6XnX3ZTdNURVKvyLNOc5FNElePnxMc4BsgOButnRhBjx
jg1J5JNQwvhDaE95huoHh/ASPpQo8apFPdI3JHdSrCMDo2CdSngjWHc1FUGIyW6D
83sC9DUvHf7bItZPx4D54GREMFC5m16Hb5BN1qdqJBrHN1l7GTaOcXRbuXLnIb/H
VEBapwrUnfHI3d1+mkCdBf8GHSlKnoEQzSiaFtq0nx2reLbdkoBWlaPNRsgQX8Oy
r3aLTGIkLVOlSqpUTgKpPWyH7Xthi3cBJ0/aMpkrDQYOtctOtPUeBG+HwTZKki2n
YOVFSDbgvthLHsPP47mpqNzzUTh73hWFMv1LE2Erbzim/663N1QxfGvu5mI25wyh
NrLjckLMgzm5R+NeDOwqmrV/z6L+i6LwLF+CAu0Gqk9BH58gCeOzietGoTvx8m8l
bcT3j6aQyIVOM2OT9Zy9TjOtqGBlugWH3TiGvclhvzRMWck07X4/+3rzwEiAzFAr
B9I05inPkvrNkkgPrNReBWq3CjsWkzJNeSS+aSZdvn1BkAz9Qd7XA9aSNsqiQCRT
vl59ceocwDQqxjE+BLPMYE916aJVIdv5ilVM1iWsDa3MCSH+yDSGnTi0scdgJO+5
JwzTWQPB2KK/vUTwR3Wn9yj9HLPvFhUzl2zBTC4ygfi0HclrkmSLxlvYfLwfCLBb
OKi956amtjnq892MODEmutNouRPYNy1Rt4Weg4IfKqrCE/j//K2w+EMCgg30/wWu
ZfhQCEISuitDiQlkNbgMhtDaxutwfd+/pQ8O+nwSPUacuRUYBRI7S9DyLrREUSIb
S1HimL3+YzA65aBQ4RaOWDR+n2V8aju3VHEThPzCapJ/kxTN1+kfhMtnjMmgQxTT
kO0QDji0h5D3UDnYs7SLeO1XNwg393BKxUerDZhAYy1pukuekiunr85u9/Fs58Im
oMrDTNxH/dVlApABc/Hcxu5WWJhE5mR/mS9sxdbuPzLC1rTNXZLphfLsb/Jz6KlB
x0xy870GoJub0hWuVG7PWByx1q/7y2pThub5vwGtv8sktlmV7plrpSW5BVBVgYF3
1LgZGmgdc+0sNwOdKTqsJeJlJCkfk0dVx06+xaRCj7QdPi73MXCOgu0NP2j6agpM
aVp3Jrrk5GxnRaZQNCJnOOB6y5xOfSSDWIN7f2JHYRdzCp1Q0XPraYQYG919yIon
+v7tgZ+DInFwv9jWvAMH4Mfi6GUuVFLS6yws+HJMcYvi/G5AgKoFyVbCgJmp9+kJ
mRgpbU8xdxM29lV860+UZrHQQ5Zd/n2Fxxcz1mGfLgtGH33GYWT8Y2RGKKOWUBBk
+G0enBphSpAxkeYcfe5jcvnS71XQAm3Os354hKiayuR92PRr7584u95LqdIHT6UD
QGn0hkGAwEF9/qrM1Dt1ZKugySprgUfBT5S+4mN/PbySOveAOsHh+3XOfmDxh29t
Ujz+ZNAbbxyrquH0YTus4ushnMI9N9n/+nnuj03Paf5nZSSh+Y2gEC13qSmege1J
JRCypH/jgJHEDnpdXYXX0n88UpLzU48jROoXOnKV3Lw0ARWBnDVBRhMeb5BshArk
MfkD6gqd7gpi6jPZ2m0WrWaK19GFXthKa18D36mnxllqbPzOvvbTQBGyV/rHFlTt
OS+dSt7wvb9sr8z5QwlEWPlF+RxK9giLA0iD3tlsLUDo7IsBDEj2NzK5Lj7SO6Ik
v8kHrVAjUvVbKcyuRQGpFmniBkjSBGcKxm6nFXZy90MKEBHONRj8BXnU2/SjzXws
kv7ECJS2ZkYDnBEMFFSKnff95sKTltbsBaiDMX/4LHQm7j5WUXM4Rqs+Aip5DtuT
eG+QPTe00LFzcH5qOchoofJSpGuTNc8CJFONRgDLsjrqUyhY8MeJ9pS48XdpBa+m
+0RbV2rLZfOmRLKthXu3NMxHTPSE+42+9BGxndLATajuQ+B0dKnKg3D0n1ZO4bMC
lRifgaAIa/AFi3FJ9KMxp6aJ6/C6utke5K6wSfq2LCbr+qsFza0NDTxgWi901/Ld
i3Rf1iinqKUScpmFejipuZI4bMcYP9u2m1zTuF4aXwGWsLbiFr2cNuBl5ILFUszH
6mLJyAW7osrQPgW98pCs4yrdgxMcnPR54LKsrseJxImAE2GUFgAXSDFAm3sF7i0S
skLgIMm78Cmsm4taRe8/nDraIQ6YyoHfBuyxUUKGL43QnFIYMLXoRTLR+1vG+kGb
nBrQlytzezsOt71SfpRjTKLdk8DQdRqUmwsWZ7komrbXKh0hbl9sebyvwx16xGVP
myA9iGT6uqVDfvw23sZfMQrJjggKr2xZ3vNb7FsmpNbxofeo1wdGl9OUTr6RH6tc
9pQ47jTIM2enB5RPfU9ga5LXJzFlI6ehEM19J2zolxDUH/lRkL+942GNNsaWnGW9
Lf6LVFDN9qef1fY12owcKirtrlETJf/3bvlVHzBjoYPZJYB0I7XFMq1mKl8lrmUQ
cxE3N6MHfX6tV+fQFkI0Nx2SIuI53hjiftz5md4Pm3CZB7R6me3WKMW3dVROb4nR
xhsy0lLR17TiMTbDZrYX09XPSxlbNY2d3A1oNRWYidkFDhIny+TgQBRGCQMtPU/+
Q8pWKJRdmFQb/f6ItHSkL28baEyhB/adK/irYGMm0I3LQit7aH5d29UgQ0riqcZy
g63B143luc5GpPG66YUtlZqJNtrITQ4nnwUaYbZiZhfx/+zKLsHUf+8zRzxp0qmJ
cO916kcIipOEJPue6DNqMwlLkfsJo/AUAaj1JB29Q4B3jA71oTgStRvcy131XT+c
Nz7+1IVjZ7zmN41Kkk8be3KHHA7CwfEAhtEHNU4fPgLUxtXlqCj9stjGxJVkbbXk
YqMCNjJXSN5QHdF6JFJuA9UyxsprCVtcII7cysuxJs9iiGuT5wuXhOJTsDoKGhFN
FN0rEd7y07Pr+ShKthDXmqE+yY3A7kU9cUiM64dATEtT7TfJIVorS/XVAncTLooe
ds5q9hOmn8CHFJ5Qf35yYwshsyokvgAaGKGGLDXIHAE4bBQjuelwgdSA1cj1mwtr
Q60bYR2kNtVCLDtd8ZCjJEnxWP+lfuxiefMrDrB9HLtTmRC8jiuxHfUIw+AM8IYh
zT+m9H4jQhZ0PV5twdKTOW5gr7AXwfZGsgVdrDTz/HBYf/vMpbp5dUe8z8C9mcrC
HUhjMI0hGsKCxi3VIM+eD8cOSgIf5S8gO5B+004ANlBJAyG7wLUdSAeRhR10qaH0
S3GUTqbAiqHHk2+tpP8akQ==
`protect END_PROTECTED
