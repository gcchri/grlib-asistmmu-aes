`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CptzQDwd48FV+TF5Kg0pEzEqFoSwOUvOxHzB7WcVoDKPzXoULmomq8yv8qzX+IFo
fiNCIObctC0VHcaxo/0djfg4rX3JG7MJiuX6FaFMCO7TQSAUww2vD1Vr+Wl5m0EM
AiQlcRYZv35rdkhIzob1/w/GJHQ2MQYzz/ZkbF8jPlMtaL18g7szwI+sMIceW8eo
aysbeebAdqZ0/Cd3Z80xc2pWzn895nvaeNCbvvY42igUr+VNn9bFkkeu7jxJCHcD
H9U6N4AGF/GQhRQP+kdi8g3HaW1anqK7uFAxISU3xKLM1XSr7a3fbUAjAa33myPg
KxDtizc1tw6Hucw+ljql9XOoVlnNjcsrRj/ppvs25sEAjs9/tfL+/99Z/SeUBd66
EsVCRyHq+TgQ/U3VJxFG/w==
`protect END_PROTECTED
