`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NmzPgb0JLz1cSOfvrCwtgOKz0dGuy7rq7qidLbZr1E691JAEVilB0sn7vp84y7PJ
V0dvKeohpP2Jt73W0HDn/ls4C0neQyo52TDbSKrvWTn7vQtfdjGOeHDSWwmGoTQ5
SQYoddF7ytParw2/8mDtzfhXNjrPcajBR3ghiRMgezBKrk73ZLtMVicvqqyPX+Xq
ljhNgWLeVxNHik1Bt/OmwSUhbK0dstUkCwF75Rp5NC9V4GIjK2tzh4ef2tNPk7Sf
o97F/vK06+/ZkM1NfWVatY1iEoKFExFJlda+ni6a7utarwbdHsaW5UMOwWmzGwsi
tiXF2AeV2CEKIMHEnSMxwznhpSRZwt7OwgGlGYqshRUJ+FsUY19QpWIxe2Lbp6zl
yX0qWU5IEEsotUEi5eW71A==
`protect END_PROTECTED
