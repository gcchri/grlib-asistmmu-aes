`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wMZDzU98NyHV/ysB/dWbmlZ02yzzqQMstGJB9lAhWEwrQxrWB0P1UeHl5rN3cTn0
GdOiH/W/sQDqqFzFXJWk2j4pPz4sqJEIJH10DZBA6s9vixGn8PxaV6ykUGReN0UZ
T02pK5CPJPU8oYgqvjVuLoURyQN77Mb5t5ZktdrWF4ZeiWTj9ohQTC+34MLZRntH
q8RKD27CDAVKFdfLjluR+08bgJdp0Tw9Q1j6WWBqA3zLCSzjSVSiGKsh+lPfb2mL
PVLmdEpL2xq0+qO1rxFgwzSTClWHycCA7cLD6mm/drdmzt8W/FsH2GJFX/c98EZB
A6nmPdknDvmfb7eE73L559qQZAGyjgQQED0Qzje5CTKewsgsfCknREMFY+oXoimH
OT2e0ViDdtZBEGFuoIdrBcZfSXnCF/DFY+Wzxr4oDpDP/Q269IDeRBy+UjrzW+wq
8iqBKLVTRQBx/Cz4MjlfUP+iGfnoEUitlJGGerh39meY8N2C8GVg60uHBlnq8uYj
uzirgtRv6qE4XByjVXfK8PJt1Vei9GaV4+zAyu3BEVOqfXqm9WyZmYtE+j4eQAHr
U9eAKw1fy8naNJmy480W/VY/vctx98a/YEbIadFZ535v0+mKw4U8kccvzJ7ETnoq
bAtypwZakZY37fOWAiW7rnXTNV2tU9cpvdtvZGFcqm3RoWi1ClcYV4UE4ALo01FK
YDAWo6R2gTCYklCy0G3yRvAr/HK20pEghPIZwG+cvIc2RtPLY58EJFKDb1yxrV8o
ZzMZfP8it8vjTXr5bn8quQSSLPI/tLvKT7KFl+N6uBAqFZYm336DG7b7VtO3HOxW
xkyCFTJL4rIrIvZeYLHhUpYd3pAAB3fb/i96NZr2Y3OUaXbC7FJ+MAG5qSPphun5
3gk37pWOLCFloSKI//6FU9Lv35wVpeYXItfoufv8+15kCzqg0lPExpDMcuseyZ06
FIii8yoovtG21fYJ3WllebGCTs9Bx0plV6qpC7Fh3tVrltk0/GBRxqiZwJ/weRay
gY55yrBR4W5GqyaRjGYDzAzDuv1XDjrDN6KYbpUJyix1GR5Qn8GAgywGGo1gnU15
41d1FNGmx7cXZALvscDhDBs0Gy7zEysZn5H1tn3wrlZtS4TVmotIrIQRlWQs3SYf
ad4G9QAayxOY78kdt14mM5IcVhWdhUKPi/u533BqQSASeBdfF2z9t7l8QkDnuu7S
hy8/cjUbgFWxOWDUp8PaUQWtFp5uYC8Wn7RvuuDcIoyzo+iBXiM3JSXm5PJJLDnj
kjMDwDuEKwNXzIzneVZOMWdRLu1y10ejcv19bpz+irJlCs63n6RAKWbxlN8eXjL/
l1TPKHMlAtaOou2NRayp2ZA2QNL4his8HKlbZnFixEo0dqr7dMFik1LPykFYglT4
o/4SxCwbgd0x+l59S0RI0AFJsmzAF/tgs2MbDPoC51PSSn4Rv1cucIaq/q1KjIwV
8/l/8ix+zW22n1xBjMh87xRxoYcVZS9KGCOY+8I027mIfH2yKL1VzH0puR2CDdzy
GBHUrxMWhYJSxAbd64MSqddV/+MdpBdNa6wt11BAHJphzrOzFhNesVpEQqhyMHwc
nZcLMLV6z+yiwwaMPaHnyKUdGIRWM6GSVmgEGFZ0ZWlSA/Qk6Gfbia7aKXBVjVq2
bdbmH0fVz9smjs42OiAM8MruotRe7Tu59nWgIk0eGf9KLzGFYzBj3TVxKTU+ILEv
FO3E/lGfroJ2+pBwT4yD4i1Wr3x9UmF+WJLGadH/DONTdoYF7jKSHis7w+Basp2e
Aha+Y8c8Vl/4WvKshdyyYSwk3ZC4p1UwYfiLdCk0WgM7su6L9q9p67mHEtr8bNdK
bHhvNGRwKUGVvDoiCVZrvxXbTZ3epEiojyGNZNF3v7wb1gisyV76azPU5PI5cHZZ
gqxOzjRdprhoTriLiXjCVZfgFxqTHsJtxp29WzbgQFc6dgdIluMMrfzwz0xbSFgN
XmK45BYIL2Ueni7Ad3FfmxAbHwKLerJDfF8wXwZJCdV1qu/ImiOpW8ibxGhYkEBk
AiYdUWB9NU3zy5hPSAyImv8tYUECPAcSY3PvoaFXTfuYUPh2fC/lBy0Qxf/DwaMP
bvn0CkouBxc+UdC500hWl22ZHO/IdhIdUEJBXyKvfUIDbiEelIfd7ySrNgYxboEp
KIDThJTWS4oq46B6NsVBukIMVbuin0L9mcuCviJe5u/USqtmcJDoZJ65EJWq5PbH
F2+eQAaismDYVSg+qinNqTEh9TzaE7k/kmHiLdkLLq197Wmu9pTUeNoM6r0TpcSD
3UAQV7y5rWgig5RKdi5hG2j0a2jXFBPORkow0yoSK2jebSlgPUEx9oZ1GsL/lxRd
MUWuHxMkQFUDdOFYsU9GUScMdmH6g1MkjR3INznt5nSRpFyrzozpzRYc3PXTWqQR
+NFqxYjBRVbD7rNlZthoeMlZ/14BqlXxA9MSbQZiakpJxbDBmE/kpXEQclBsLgBj
cCtyZG5l11aJqVBLDBEdkyG6Cmo6LmZg91qrllRVA+7GEa97UENHA4XCtR6Lbz4C
RIbn18LvGpkhPCIq1LMcfsiOU1qAW9bzZ0P4pMOGIO831Jn2V0V132ILjcBZVq7g
u0ppCmxDVoC75XjhOKKT3UmuGM2AfiaZtzAhb9PszPQzZ/ld8hjI7iag3ekGnzh5
dj9FZM7IJrt1OxylQLhU3M7u5b1MANw5a4RJkM6ogD/KknkWDRk2qRRZfjGjwc2b
H1oBUQBOIwfUhkmjKeDBieNq5o17j5I8B1Qu8mjtE14eDy0YCBUx0UdxoxZN/kiK
A6KNQm6uWCItCs0AQzW3ewzCwFgttzfFh1CsCzDIfhlPNAb12JWDlBbIgS67CGQf
ZNLNkTMjdoudFPiSb9HcixLdvXmdYy1D4DWAr+F3qTSqcafp2i7Sf7R8odjQyKMb
qbXew4tF3dkNiTRSAPAsuHqcPQXl983Nr4UsWh/kYjR/pt/1xbNHiOR1eHaAVwCN
UuDvtLzPYNGZyo9KprDwNDzG9UmKuQ/WHS8VFwtoJv2BSd8Yhm40RfHJxVK3KjPE
qKkparGVDiS4emU6GZH9BwcjVYj5/p6rd/5DtGebkbYnT9wvrktgoHMKObAKB/nL
INKm8q8YXO8sroFbptThD6Lxn31AMWRErdyIThdnj6gL65Pn7xjK7nWKQjEQZf4E
1nyMYFvRBRL54aMbBxvZrt04w1T/hzgUXh0Ir6T1YAB2gOtr6xmtsSwnelDtYL1F
Kmjx9gIDYaI+oWYFgd2fs005xSRjpJWG2+h3+nyQRMCD3vo+MuB7DrBa9mUtMHkr
SEC2QONE1V5dL2kySGdqS2KuLxLJTvcRofkw6iuRcewm/Uz0/trMrAuPLkVzGD6d
d3l7zZ3jTILUKgOFyf2DFAeY3PKNkRLmUfY88qSj3wFgj2qHRSskag2p7f37CYJ3
wEtKPuUadatuuZ2jvsS0hqHNOfY42plIYd3g+B3oSRf5nTaDuGQ83EjxLiilRQ7E
Ja7B+GFfG8QVrAwjVcwKgNaqpEGP8fnHkDTCdNmr33r/x1l/QGFl44FHuE6VKw0C
4rcjjYseL1UVRzvh47YTtOQSkvk31JOStjt75lYxsoFp930Za4gfMbPRHvgFn3ea
HR+FPobtnRbbJlAtpe52ArUrzkIBjllSPTeYSCvfwb3apMTEBRrevlzXt+kUcYWa
q4lHu/iXuBK5gHbo8gQ47vJAT44DUr3cBnm9mIJTiuUmIMpLbEvu1JIvqHxS4El6
CBa6Kkk2avO3G88RYiI9p4RnY2xp+Olzgv33wPi0WABxN6prDkFsbHDgIQdH+/OS
voADfbqscjTOYRYtRy0HvnWyhXI+3R0Ygy5rAupUMq3yCvYqkD18x1NBN+L2+NNW
5NAFGVzFCjlyJIn564j6UFAtnOKzi8z/5jwMfLVezqeLV4ZtmoDSE1mNgFvfMClu
5z/gPH61ptYrn0HGn5QU3UWwe3vHBinkK3crg5xM66237wRP86ZnFlBn96ckVaA7
j19VoYxUEMxcwDHdp0WFL2fm8UveGYWx09/OYQYcJusj8T2Kp4I0x6fMcApnjkYz
mckDOlp8kET9hlrz+WTxJpfAuMzYOhgp6MMpgJCa3UOfaehfr/KdCIilobLO7Z20
jnkSq3ClGHnmjcCrAXsRyvipydgYQMkYrqkqy03y7YurPtzj8rhaLYqurkX1ognK
AVgJFJxCb/Vb6vQUtwckZ+oIQ2DhupqB0bfmcG+nFHqzZKfxuAYEMSPK188Kohc0
lISbyoquV7S3I/jzhqp67ZQQX3pvqKlJ3zNuA7787KTGLbQeeHuo3EvtoZj92UrF
RlKzU1Q20mL1HzQcSepWST44aMaOEslulfj1muzUHIQXifmar3gDXkG90OEWc9gB
/6RjqcROucd7k1vWlZg+eL5kc9MYrHJubCGP4CXrZC5n5M/tr8ylcY7Aj4v933XL
4rZGSuHgUkvLwkg8W37L1Apm7IpBvff+Z+ys1eqYSMgmCC9XAXSLpOsBIHuyS4cI
4W23frbs30JJzty9+hHAnpsHD4j5KUBbILYHzrdVuj+qci/DtI8AsB3sapGmVXg5
2M9SSz2ySH50Di14L1C5ZvUUubgLtqyx5KU474bseeJqS3aML1KEAUGGSlpyQXqJ
cO43RiDvIoyUQvRFZxuv/ofY7xCcdwyEeC2JcM941UWlolU7FUP7WwzYfuMcmX3N
fKZuPhbhIlVCHSrctksRTE+PURauSps4ESHx0lLoNOJyOiM7nWFx+ugjG7s/LDxJ
rb1k68d2Zi+PtTcU5WQeQbEhdpgud9pwjFk+wgjwWIfDcHYmpiXBu1QUQPhGdKpC
smioN8oX6V1NtMUVueE448gB1cm2T+5ZVDDVCN7itlae+PZqgGIWTih7P0NlQKw7
cJk+tGlDd60nzH42h66JbU9/6WL4OvihdPrjlMxdRgcE87IPDLr2r2wR9YapTVjF
QoH4SmiC7WRm8XUN5nXFi1GjxbGplkG5YIYhsoH+qaBcG1hBRoTOmTiq4s/nZiqN
p8G4ydZwSegeHAJixMhegzPSQIKO5dmMuwfQjioasjJoj8urYskw9BIWP69528sX
Nnl/jVBLHgQ2Pynp4UXDW2PFPReLycTNpbL70TMm7VCydZhz4TL8QNUPdxmF9spv
i5CD5VDkqko/Q2Xv91Ppg5b8dO9eZj+sbqUYNAWNzi3tV472bzgfg6hZVDfhpctg
DWXSEbyIhMQVYkgYgbX34tWGX2CcoBGUKD/VXgyqGYtNK6ygkNPiOUQkoyunA31G
MdRTXsC+iLgwBRmJQ39SNM4jtIbfZBD3F0cVtC0u0xbc78uKSQMLJ77TYycrXNYj
R6dsvmPLmzEzwV3bCASvi9/R0E3RYSMmP2ytHdVXnI5WeSiPToUUQkURvRPdVGHg
hpWY0Xe3xZVhMhhVZg6IYnD57q+3am6O30aOhC9wzvttiX9xVoGAr6qmtCmroZH8
3QPK1Eh2i58csXKMyQUqEqfTP8ZhE0pOMwnoKLDegXb7T11y13L1HO+baySvqOdz
zpkGd1dJenKwuHVW0Nj6hO12UjYZR0t6454Db7Azhkf80EkbxAfRZDoNsBjsFeU+
zXwdPcPH+eLtTGj5TgyGoSXwWNEt5sxqA5yKfY8Fsg38PG4MTyyixCOEPDzJRfkh
`protect END_PROTECTED
