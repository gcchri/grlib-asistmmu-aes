`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BDHha3iJw0oZIVQHwvFvUKBpLn0/rCSFtE9BzTxgKFUOIN7qqc/oXRGHTn9JwPbw
0ITh1vLraPuYGLo4zTDEOqkchqM1qbTLy++whXQv5irn2F0VHAHJmpYSZyrAfr3y
he1LTTid0w4T5gSsZw6+UNNOEs5BrXDblApdeNcuJjjf6wcPkFw2cNFgNnEFN3Eq
Wp6qRu1vKQIu53+nnYg0rzl5l4hxb6Wrg8d7bkKzaf9KW3Xnr/ptYlj5FJbAKlU7
HeQ4kE645wxKoIYRtgsG2lGCmipUGXVnKyTn+ZLarliv/rhOz/Ll34deU77JGxe4
MdKV2l2AnIIxwFj0bW10CA==
`protect END_PROTECTED
