`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ro4jK85Yc1hlnfR9MaMH7KVpUsJK1NBovlDL6MBKUAXAPjqjW/tOt1K1Zvt53MQG
Bp8odpYlz/srNKg/aKfGg2nAiRcprKBOzPe7Iwx1P7l4PwscfpOKcXfxi93DZr7e
0/DYh2ew8I6OhbiHUB+UlEs4ARNoVGR4/w3Z/5tSITW/ea/pxLCJZUMynmyLYhwO
d8QLdz+u4czY82nPFGP52MlRIFCbg0b9mZKWBS1M/3bbjq2Adzoeqv3qhMEvF+WB
A7Sjw0/saJ7WP7nBYXUBIu9XxsTBxO44fIR/gv6pmnQ2HDtASC9C1jtcQQJAmQWm
jTzLX8OjNtMt3IDDURBm5b0+hZ7oDv2bCJQIergoAQ3jWo3VwnhnR+likfwg3m+f
7qByRpI2oCsrD4rumNnOAmHPe30WNu1MjjBQaDcgNZxFV9FuXVKtcZnOXoqqbVbb
MDi0GbssPIqeUoqv7HfQ2UyDAZZ8Vap88btVOXtjb0BVLR85M8j2BvhqRBFTH45U
`protect END_PROTECTED
