`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aa3jODAdglQuoVqyIhXBXZ+4DQolq7U0x0B9dkFcBtmg/sTj+AV+VVK2DhF9UwT2
8rgdMW5FfGtNACaEVXeJJKU+QYq13uXk/FU9AdMcITMZ6uFMPPCLuOpnublReV0h
wn7xbGa1pjupTLeHvEDv25q4kPckia6sY0++508BVUETnjCOltf513Lg2kF4KnAY
aF7wCKl2kun0yjiYUgq3ll/FdzH4It/S1kI1rWVKMGXlP+YsikfXzV8RiK9SxsdE
PvXXQYY4tV/7qtIpGN/wlCN+4+eOIkyWO4Ebeuw9R4Dwbu6yiz+zJBlnMcDTTyxB
rqXvg/tElUZC4HBKciXb+L0Y84tj/zOqEEpCeDdze6bvpQjBwTWOog365gEZRLtg
`protect END_PROTECTED
