`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDyqjPPJ3hkfV2TniJQATOffjA6WmuJBD86gZvcl9HtS1cQRHkHq550+usjBN6un
jPYBoUTMXOPuCrIBT2E3SpfqXFaeaKezJxs5csLFjJP+TKkKTEZ0EDrfRZ1lClAm
iR3cAfibKVKt67E+PzxbSdwAy5r06JIgnfXgpKaF4xxpf4TO3lMKBANSJIN2mQSR
KHx7L30J+MmXmSRxlj89w3EhgwR8NWS+uJ+FRLu58tPLTPYgvkgpLokwROofpN7l
UlC4tPCHHgn13lUyZbV6PzN3pNq4udr8pvK7xheJ8wB2VuyBwoLltQONbuQcANBI
1acNk8NgDLQ3iOq4M/61+q7DtS44FEeIUR2fX26YSlPewfXu4dTBNe4iSvribqjz
iC4lAHRNiWI1qlt24FSH/0uX9FtRptEgFPiTnSkt9Dq7k8C/WPbgKyOyIi4JWjTP
9Jib9W1nSBH0LnTW0SL3nyVjIG/FpTn2OV5dTY01aClkWp5iSsI7ih6ZLjHBWRD9
pTm8MYcXG9Ve0J+3mkqYO6Xfg4ukNcxz5FOeVwf6STRXNAfMAUmiL7lvH2G3UihH
0PSyb9002hKvPldRc6HeDb/Vgvy4uxgCG0NlnbMDEH5cml2VbYt9JXP+CAvsw7s/
yvwMae5IQLFAjyB4Ggz0xnRaJkQzZLnZN3poUFAPNgbfvsJV3Z7yPaGu1M7R52tB
`protect END_PROTECTED
