`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
96AZyrIbtK5dVh3vTebh8jy/49vCPxrx/7nm8hYnGqhq7dsBwEpy878DRLwOAsS1
8yu7Hgnb6Hh2rZfeBWF6vwkkEa7oxtHSidrrFz3QGTcv4sAj4xB40yEQS+cUODUV
+PNv5XZfD0iLtKXOEKxtUsUvOUuthqWMZ8c65lC5xXcTVXDlMwHQhfGtbb3gEJPe
UxX+fCqGbh20VjgbxJe5CBy1G717l3oOzhlDJaZcyhb0mgg4pJLiO6PSjQotob0s
KcDJ3EqwUhv99JIQRfmebLW7kqovPMRx4gejIAct4Kwz90YBU/2ZKO0T/GpOdHju
/UqJduqADpLb+sWtGlLQcA==
`protect END_PROTECTED
