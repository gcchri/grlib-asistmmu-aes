`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XE6UE7AbwID75RKkt3xIk0yGBEzD9HA6puPRfW1NLVcviXA34DvWJ/byiVoHaN1F
PbtDGJbrM4kwtoilI3C5ecrfPoaF2NN2GOj9uCiU0TOJBzkic3Cl481CohMFTTfr
KKQZMLMubuLURbZWx9erwoqzeugq/RC3+JgdDdhX/Gd1FjhJ9U0jFOoqV6aZUGjp
DfkeJ3Kik7Yf7RFIHJAuyM6XIttjQKY/RbPwnsOj9JHILutba5QCUzquGNCggLjt
Wv1vscIYhfqa3dt3LAkGCEUXZiCuEWKocIDmNiypusHIdq4NapItVY2owQfy69FQ
TFy123mN2+2c6H/Lt8rbpl6eOLuQJX4CPfu7KdD/FqvxBpwd6y6ChCv6aGj3brkW
lb0udhpyl26l+dRPW4IqnOylCKutoLnV8iX7mvne6uHeFTddLjG6Wb9FNJxZJqRO
hyWu0L4xl3hLkHkNJ8yStb1JneIm8KH0AbIaccb73pViOCJjc6aqvC16DV+GxOzT
2uuAgxfwmBfFBqSdfUP4qpWvzdZAbwoa4iI8QS1ggFYTiEya5EKBbW0uP7Y59NQA
MWsnD4MPd19NYsjPQ0X60tVC6C6C5eTyFtorVU09Db2sSOQyZa+aXPeVC1EgNl1+
LxHXSCplVEG6V+BLMIlLioTCQ4jPshBGb9CSCbRD6RFsiGVudcHbfswaD/VpHfQL
GqvwVuB1/Ar5tbNf/EFLNWACf+HVbZvHdMYRiyVn4YIb0uKY8a9Td86VAsdsWwPQ
PqAhQyomY0+oDmkZe2IoWDmOQ3kdVeEtKrGKlGbOGjhmqv66CEPnm9kNQPnFapoc
StkG5K5dUaoKKPC7a8X8wp0dmkCmBFVsQwnwgh3RE2lS4MyY7IzsgL87BJ1JlJJ6
+aNiyaWbWZ4Mio9MB01iLbHUSHjmJd+SkRt6OMADoEeUs08Zb1i4B/3c8dBi6YKn
0eEsP8mcu36fF+2PmSQ59gaRmsuwZuLK2IkJa/JCDAD5MCkgl1R7Rag6t6KGYcnc
6zQMijDdgEpN8DySjmkiDszx7DLmtqiIMHn8LBsuEEr8leb9w8Dg2E5wgJxTKXRO
XJuwYfbu6Cu1Kx2+agdREX9wC0m1HT6ZGrIbnuW8u1tvC+0wNP9RXaRdNL/4GpB9
SPeTgVGfGs7SAcBVhYrPuRTchC/KWSySfVSIIYppJUy7A/9vjN/eFbsccPu6i7Vg
NxK7ZHc5m+a1rrYjZLUz5/GlcMBSAW0pv5CJqT6chzAPE7Y0DhQ3AVq/dXfrVva2
qwe2IEfo8h+7HvzoeJhZc+q9zvtxoTctOChpRCtdW1dfEptutbo4ZAk9MfWYQ6JZ
j/BXu6fMkYPPdbHvqMebPc3NK1efcngST2QLVLZim4M9rnYohN35F0cvSMvLAVMZ
Ckknu93TfT3BHq3PIV+UpRa9ce83xCa3gLw/nZscnRasLon2CPFEAnWUsVGZYYki
UJJEG/d7jrezVH3KVoZ3Wv45eLGocNHv/NuH+KEMK4XIB+B47WJw8aPxq7j3uraD
qRqG3xTnmBDB4TYR2UvaJs7wF6a7ApFS/TLlWsVrVBnK+R7Ou89XB6rkBzRlLng2
nzd976y0PN7LAQRu53z6rEhx/RkyzZ8p4g3erRk7OMcW+9oxq07OSFz7Zcs3FgO0
UJGT9H5mYjQFc9TcGrkzcHIQvHqwCx9jAtUE/LYp7v2BvGI7bsq4NwqbQmUONEPF
teXfPo6rNkaw29nX0ZR/UFgTNsQxOZc9MMbD6zyBY9GTla+jBNx7cfSxjK+/h8fv
Gjqwl2PjdGC/Jes0ARl2T5P3oDsFVcuq3VXvBOsTqefDsgbKudF5iIALOPakN8Lv
DU6H8+ply6UEB1k44s6pJvLgm66ntULsECWD1p96gxV8sWmIN3fwpLgS1uYYeJvC
8og0eH86HexOc/g8Fixg7jI3p0WruYV21bmz6XFIegNmAT272/LDvOgShQJzpLHR
/T+TTdQqoFHWtAGph26ZSg/3OHHQK190S1Obc9QrYumbyDc3GzBbHVUTbBKJO3Bv
Zd6l/xALaQJrIjcR21wpGoflDO5od/RpXCbw+v1k0PpC4e9iOKhFNM20Yomv1bnc
lcHwbWf8WwXIOW8Xm9kl2IHfCjJuDClY172c8GZPW0l3soEVuMnH787txeJEYtvy
`protect END_PROTECTED
