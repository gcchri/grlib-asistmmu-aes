`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYAmBi6arYQU5aVJ5aT5dKoJO6aRkeL8uAZPGQyRzTTIZl9CxCiEGTiYByoeG39w
ET7/bEEWEQHdFmh4OgX0vkqKKlihM50xSWE93cdjeKtsomRvx09/xKgC0rm+1Z7A
fR0RaetMyyFVmz6t+UY3sGv7WM37lraQR0vlKoMWknnzUPaICJanRYRY1JQQKOA1
8zfxfxo+cENOPcEtTOEz7c4Gg5JIaUpwu4lffuQlP3vUTjjZJ6IrbrBOhVrNcOqR
RZKWk583AZZ/2aVFS2ZiR6Z+Ib55m7M8NqDau4rZthMKUOSCyXXjEmqVRSjNDiWt
qP2e0V7VeLgGkLJzCQrvhBp/JpLa7mlsOj5JZuFwljFyPW7osMJIPVgFjj+VV+Px
7kqEyBCXLL8eRNUa1VxwyVceRPo0HxepRYeZIf+O+Ob+iQubsEMD4bwo4CQ1+0TF
MXvqJWSdWwiGLfeVPWGmxnf18F9IMYpssBKRQKwTbXtx1Y7NU5szjiOnOgQTNG57
RFhfEzgrJQZ4hJyFoYSZcUtnEwqsi0AjG7vn3f9Msuz1HK8DioNaLh26UJPzB8Ly
xT4F37/bBE8gVVKJflyXH+u/aOTnSlDswtkOZjehOrofEYAc+kmaB6yGH9S+B6g3
WbD0g8UcPAdVtLtaG1BU1/mWC2k6kbUrpR0u9OESFA+fz/K+7DMAQ5zwlSjAt1Fj
`protect END_PROTECTED
