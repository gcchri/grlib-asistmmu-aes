`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxjZMqQrOGsxIXUcD523D7E2vluIOeoe57LA6bJN1CnrJq9ia2fQ0yL33Ypy63uF
DoBRok+K34FRrgG/W123BWtYcr12jwCRwnEIWCC0/l2P/xE9dq63xxfP8CTDCWoD
bvQrM2ggHuoKVKGdX5Sf9aNTaMDp8JMvCGrdzroHOn2rURVWqSuXn3YyKCcRcwZ/
zV7rVYIzTK9B3d+p3H3+Tz41Egw1jBGLLhXBPHs6plrx9qZ6dU000hI9I4DaLJwR
g0K2sd8DR4LKIj1LoUdbPi6KN+wZyuA5yKE9dlG1n5LoxZYj3qylXOIm5BZYCn2B
al+owASMa8rwEDUUdVvvfWULS/IZV4khwhB6JZAWNQlzGBq2daZWXLOPqlXpETPp
f2+BuYewPBKvhTkDsh0D3RNeIGEC/tChi70zhiuPr5qt5yF7iixJXdukeB23Kzbf
J7QZbp2t1wbY634HwKj3465ovs3BFYqsekyGyBpxPg8RQi4fc6WrjBJzJhz8rfhY
`protect END_PROTECTED
