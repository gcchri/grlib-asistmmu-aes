`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHUaiQKQUNIz5X/+FXJq2S8udSiLMLGbbKWoK2+ZncFs+oDYop1fOMzawfo9jZXW
S/84d3X2kr77TBhQzVMlsoIPqZoLYL+J8k/awAI13nQwZ6O7Eydy2YXO90oRRbuf
FmLCQOZmlokIIspY9s9G37dcDyf2YADNhd6MON2eq8mkTKUD8swjgYWugbAWpQgl
V3+KfKk2sNdsxgc4ZuSaQ77yDUhoyt10XpJB/wnoLhVz+yYZIpEpB+uKRMPHJO8/
sZ3xFsq18848c4T3+5hlpgG46wFj2WWHmBrs8f8kOm5hnBWxo1B8s/ZPACLlSy48
8yCy/x6cOoZXEkemUxuSBMgPm8JCP1wu9ObC87X0YvcSOrDigVn5IfHCczODB8b7
ooKCvtpe8qeeMmS0fCbzCG8W6VNErX2K1gwXqv415y0=
`protect END_PROTECTED
