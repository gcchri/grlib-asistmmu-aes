`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rnGcRKRzWj2mqQnqFb+SOKOZOAAKxmekgWUDepOY6X6yBX2zjJALi+1jfX+LaPMx
ihbmACOAxkO1K8ynPgv6OjDgh7eJKCVXx6oGnp1wzVDeZZFPdQ6fudpU9YF5ymZO
XH6UEO0XE3UOBk3RAjv1Ce6wnBVugJXYWX7Q05JqRn4E/3k931aeNQU6jextkUDT
V7mx2XksqtVvRV1tSKmaTMLUQiWp7B41yFV3JW/rETfXWdnEC7Gx9fi5P/3Io/hJ
kLRKGHZBOZQY5b5rv1kLmvnBkJyyvmAWfgE5OfpAASGmAYhMYm1+i7SPE3dQTFcq
vfqpRlb7kH9igVpe+CX7p98JQiKmBpg0l3mOlqDBOzaav4B5AIO0im585g5OEkk6
OggKwQoFfib++FUX6W5zLNKN8Zd1ICkWOY7ZGg8FowxMJDt47mbpWuqfRYyz7VdU
zjmTXZIgQhLbhbXtCFeh/EY8InWQnkHmPf/31s+aVahzHwtiyyujqPKPTGLrfXQa
jEoC8F26i/Jv5MYQebuupxrROiNBLao+S4UJW4Q03hmmWCnqugIy1CSnEK+sVqGC
hMy/L2J/ml12VgbCp0nsKVD/XkysTZUpEQObIl5pbjRZWCEyflL2a45NRT5nowJi
tt4n4rlL76W49zxRGIr20w==
`protect END_PROTECTED
