`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eC/w0vOFuYCTdvr6zVmGT+y1c22squd9Zhghaim1BEZqFewLdm494y6URlbzOZn2
fIgaw5Q2INiMivLE8b9krnd2giuLgHiGqi0cdZNydb63IHJg0T04iPoSpG8uJVVx
OIy9xqXvRPjx23qO/bXQv0YFbk7+jYgJBiBaZdhlNkX85F0FNv+PzoWm+Wj4EqtM
JIlrXI5vhaRMv7HyCtFIQVvqJenRWJc6Wv1nbM/5hm364Gyw84Ds7pHC+061pa+7
F5VRBYHOt0EqiBxb/2LVV0JFJ9+XdIPa+pOeyYMlcm0T1YVyBmHePq4bHJZ3/SIX
WObJChmaG9bVllwSgrk4WCKCeBfX3miKjUnYcN4i8rpuEa1pxADBV3+f2AVk23cx
A7sg4aSqRTqNUP8xEMFZHZEi+TxcY4AYUHI+KvRcQKh5oI//1Tqg7wLD0BRkAobO
u7N6hfv/gguGDahszRcnwAMkuYk2jS2y2rW2A0oVSOZekAusY9Hm00ICRxrgaV2q
28RvPYwtEC4ZC6coex6Du4WbgdmBNOXN6o5EKxSe/vOHlc2Y5/dqWU4rM2jw0FxW
B/57oNJvOhBJTOS3ZQxAHKxb3sDN+Zc40F6HgpT4JbDLOK4Bac1UOeSdAG3SzInu
Dbqu0nYmJkDIEfuup0CaBaKEP3raHoBJc++MTcBUVM/wiKylTC7hX0nfKEfxTVaW
anF0UvHwy4z3z9ap2Kf7q81URlayMSCIIJlTJMSZJ4e/sV3MV6+CZWJf0XvzLJb9
4I8C+s9xYm4fl8f2NIyLLknvBBsxhuNvnV1IpKMUsv6NKT1CaPcF6uDi/ihM7koi
1MjY0XkNSRNH8P/7kuAK2LOUH1NR6hKK1vm8lioh/2HLvUUg9NsbDGvripBs5o4h
w88oVVxQAuD7ObL7xd1kHCuAc8cpI+rLlQ689GkZwKp69IkRuZajqIlZQKPBwMSn
WrILnSnA+BQz4KE4JJ6Jmoz7oOWrcenGQ2hWRaNHmeYx7Uu+f4pg6xulqyeROglS
n0hhaUqjtAPutCuq4oKS5g7ydrzlnTWSBpTDVyg8br7DEVuSROwtp5LGrWSzdXor
Wtr01WRV1ze6hsr4t5vxMC8Kx87Ebt99a4Zek5VyccVHXKhQRpaFKNUR5QyWDFdi
cLs9ya+/a+310sHzbPZj4or+k8+PSPCjBShMHXd0jcqUkM0FWxYg4uiyEtRTd5pJ
139oagWq5kE0hwRyXHXxaEjtTJ6Mk1etq8wWv3bMzo7JFjvZNBDzKM2yB5SBabjm
x8oduG1Aj1BFCXJbsPiPr+cVh4skPQZhXq6cKzfpmLXCYygwtH8pigMCbif5DyR+
yGnaJeXo6KYmqRMAK1YWBIsfjxzv5WQBLqIbCxJ1Cy99LBQ3sHqzSDzt3Nw591tr
uydGf94RWYveqsv7B589hMMkSYqMrK6YWWY0jY8+QlT5jho1Naa8y6qCDyhk0lWZ
knVEMLM6J9loYNsLy0on93TkaQIVzaZlJ0VKp1UAzsE3nqZ96s6SD+qt3LPPLEAW
0Sr6fKvX2cXraFsXtL2croqePN3GHq54dlobR0L3C1NwQ69ROZQMiFvlDg/57Zqb
2QJVyIp90SoPYTrKOMFFr8lsqgew6xPJ+EHD+R02YSvMU/O8KRTfiH7wP1rx9lnX
L+mOPlomA5akRoV0wxaOf4fXLiOP07h9/0HI5CQMkVN71z+1YOHTS5IwgW+6lwWR
hu8HSeR5Hgmbn4gFItJS+Q+4+x4MR2DduDuziKQENK2WoPbJRcxlg8RY7+MDdfJp
6utq9rh+BM3WTLLopx9N1nAMF+wk2gdSlZtOpT0bHGDNb+Gd5dIPFAlmrdrI+n6a
MdK1esgPJWyevS5SRqox97/kGgVrOhDTaVHmE6IGpPoeZC+dCYLOyy3xmLWnO3Lp
3j4atYQIB46HnkNJl0TRZ2FdiHUD/OBWitvMZFII0Qp8bvexy3oV5Ds38Bfr1Nrv
lAdjnZPQk1kQKcutAuyr0CBdlH3mdxiw3X4xoy4nlavSvZBkn6B0nh46KLP5g6ep
ItP9M0+fkLUWf6Ktqgde11yeZdil5wg5une2kyntZAt4MMxmXyDQs7IFotA8gZRn
fQBlhbUpBYMJ0L/xjjtX8nOXuTYSQuMi7na2zyZyqifA5NEd5McX/oTpHKnt6SRs
T3wKRJicF0av+zeAuCVw1IqbC61QDRBFA9oSbsxyISm7GuuY5LEn92GpW//4JLYO
BQTt8qPze/s/JpV/ibz9X8ZOft7Qqp+BMKdyl23SQjQWu80T2cZM8xtr4ynCS50v
7U0D+6d2gNT9dIZGH8YfrQZkR4awNudjbbzQDKs9QucZgB0lSqV69imffAACtRsI
XPpE9pLAZHdpQx4sAaiLPv/JuNKJhGRxs0dPO8VYEe7YzHcgU5Aa9rIiIS3LnOfe
6hleMQZDsoL/xbyIyufIDtQs+sFF06IpCm42zj3PkSDHuaKahdiQghn9ZBdw0Cw/
1VapqqeG3V5sNZEJVEAa1o5mrMYJQG9v1/L/UBbu+Da6C54eS4lVA9M8HRPPPhO5
TV+2XAJb7bPPIMqwDiwxGHLaScaNvzIHoLS96tjWZGgjqE1VV+ZeqAweZhALavnv
aJmQtWqOhiZQg9U6pYKFjxo4iYkc9D5jXfNwAg527hkPy3JqsEdhq/q1Wv9iGB8S
Pi65byfNHx9Y0+nBuYP8tE3E6Cm+fRrgingSpnrsfPWQk6JA6nbetLzRdK6j8nHw
pNkRXf2MESlxPYTNWdfkczDh9OrFxCzzh4tvwigeAoCI1y+25cgN78dRWglsjuBU
EPJOWDI2az7NYRFyz4X4ug==
`protect END_PROTECTED
