`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJzcjdqsvzmvq6xEHjGBoN1B33A/M9HCXoHutvcqvLs+Vr8wxFS0TVliLiaiWaUJ
LVnVXWmJ2aNi0GLJ3WqdchZC2+Pj5zwn5bMCackTX5Hd4Hp4K81XLGMLN0zfhlFG
Qz+5heI1pVF2dNT3sXpgRkXZT2IP0GBunnOGH/KThEaeKGmu+1hCSWi+0WLz+q11
VanDbzrXHoEQNK2Gn7ckI4KjopGgVZAYbf4XqtnCbbJgEw21sD8SBcJGD4sqJ8tF
QMRW0Am3WL10EjmGu5sR4jGPFKPd7t3lx66X8p+6xtRg6C9g7edK6Ud6D1yIFc2i
ctge5Bmlf0JHkXOTZo8R30eXsIIt7QM4M/WtMNYWN2YqdnLIEph8QzMHfNlnPuSs
gb+60EepfAn5B6JlJ2ZLTQ==
`protect END_PROTECTED
