`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TgbW2qQDO01/MyE45mW+2bEZLlvJiNlnzUj7Cw+KQN3so6J2O64uI/WdFpHNb4ay
7MrCKI9Mlw48hBSJ25vUhUVTPvuH7p5m9Ca367CLTzutVBOuUHPIAG+yenoWYqnY
WdGvNkFXZ15osar6CF8Mz+0F5DxIdcQqyD5aQKH8X06Njxmp4qypke4aSE/dFHFF
cGOVnyGyLtHG2vs1rWuLpHLNEwAuQg4LDjB6RqNTFL/jhlH3CCHYIDwwG7IN4O4c
NNzHGDuS8/vosNac4YH+WNm6wCFyO4HRGtXw7AayvOGRGKNbG4TfLgS2+7lF4bsg
pdIhPiNCxYwXQbplZ5Zh1Ihg8nr8IUKm9JzmoV0+qAQ/wm0+pt1Dv7MYULoaKFaI
R9s8z/7Qcj8p2jVPrI4sWrYP5E19P5AszhSBW0KvDfaV2KvFJ4fo/EHu9yQ5BQeU
dIk+4s+9FadYy5gSDPpzL/G50LUogVmR+BWALk0ZXOEVkK6aeDSz9Pa1JxOYmt8p
zIibdWNJUWGGpHqYVopKmb/KyFm+tFTE4jrahaqKz06+E9DGfYURtp74bC+QchxW
NklSG1XC7vCAPTrNiy9s8oW0fuDVgS9NUKLtbuw7+GczCkIRCdNd7pbHEUILgkm+
22nofnRmiOhdwE9wd/9xKl/qS3WUskz3uhXjzSmhHK4Dc8qZywobM5Qz39zyO77L
IejjdWy1+VSUDwCWomvflBm0YYITqBv3+U6pzrpqr1ZhjK+1MC8LmvZWZtwyVy8P
3m6/UF324GCkrQKLPU+PQ6I0Z4cTD0a0Pgn439vLodtDfbC4SNTqjXCvtykMuEC0
iK7Y3zycq8Cbx6pH/5SdHFxhqQY4wK9bKlhHYuh2+619RudZGri9dti2C1UB1sWE
DVlop1GevRUH+uhmYHAcZ1Id3gGomV3zbDQIrvZTozX6BQwu2iRAtG0r/2dOAyQX
kUGxxlHnd5Rjqo039xPsaRuXICPmId1MSwKtffDv43xDpH8qWOHHLqgSFwCFBSTE
NcHaK96EKsGnSyMatfqbuwq5Guo00DxO3UGD5tywLlJywpMlOUjVVD8Iho06q74b
uAnWwSQ9W92/E2UHrdkhzSBCZJflEemOzpP5iqABofxw9+p5mjFqv8+lZgWLkKoS
fNvc9oz/mss954B2JmxdCZuxQv730bsUFyWHDC0G44yqWwu1KYOrv4BSqeq3PwAm
qOb2yKKh+5CcJfPAHpq/8dTG8/uKhXESvaUb50h1tgPFhAt6xVCxjgSejzwfieZI
8nLXNIkFQC1xJDR7nd/Igs72uEqmfvll8qnfYVeguVlrVfooFNwHmSV6RNeUbLew
1nhcM4ImOrQpwtyYqCiOGYjnPz6RV8DsYr4XYl6mKDWQaHRxUoUjC2CL51A8ianF
BuDSiBFXczHNxNiiHSdHIgMx6shi4r5rxNpu41N/TnI=
`protect END_PROTECTED
