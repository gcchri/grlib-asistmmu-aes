`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpFfKPxwg0/iKGT9tOvujMgqj2yKKCxWCQEku8x5Q5aBRy86B+36vbHJKTvpOyJ1
3mS7RvehJ3u1bYzUAhsXkeqP5H9tL3mpjU1C7wlqfLgEyoMGeLRBtdZPifArRQGH
73xhk8mzjYWikAN4QFwLEkloEtb/b9C3Vu9+JAF9fmzkKxY0QKCmt+UrjROtF3WY
GypWdOl+GdkqVI7qoBzm1znl8QA5uTVlosb8TzsduFrIdIfyE9vHdj3k1C4WkHLr
uR22iM6xTPCqxRFhw5UxLN4uTUNm9351HOJMzWHykkqbK+9E891r1o8IVmM4IXxl
QVXq+b0a22xSgH17qKWBPU9KdZRd3cepJuooatd+n9WMqyM5sNUP5F3yn6wdOt1I
f0wMQdMzHRjI2gGNQ9eFlp//ZbDpfw/fffnhVuTnhefCM7BuxoctLk7TXcXErfoB
FMP63ZzBGJrhpSHU3gyF2fI1e68tt8Tg/WZ58R0+Q+1nfDrnSUyhr8s2iNE0lmmF
0f4+GIWvgI1OBichWXncUd5tsTxrCm4lPqlvoLaqOU0LO5xf8fvHepE9GENy2txd
L7ODwCM6HckQq+fAgZ6W0q/NSjW0MRnyKScGSRS6+X8=
`protect END_PROTECTED
