`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+yomUnisSKNIuYYUvADuATUKFRZZl14FicI+HShWEKkWacDAI7V2wzgs6ESavs1H
nWOW1kcTTUu0rZ0AM3IeLdVhiK8EmnLv15V7PHjEvF9aVO0uEW6Z9UeIRKjE5K0+
roo3KosfdEOdwUlUZNSqZaehIeRi7LhP7p1DwQLFRQ/luBwWTUeIku0RgPekJvj1
eX8zZF6qwzeYvE24M5qlCbQ8wwuvHudSijsk37bLv046cIX/y7Hj6b8QArTTjT5g
jM5Do6dUzefdLAZRE+Qcr1TA723D/S7KF2RFoxdB+mJMIZ4WX6EMQCu8tnhBLSCl
djUFm8qTNR4E26jsTnbLK9oYNhgQjnU5p9ftI/CNtFLLUNk1KnABUQawrJYIQBOX
XPCooWztCIB9KEGOPq2Sxw==
`protect END_PROTECTED
