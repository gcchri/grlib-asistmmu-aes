`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RTPOLPcNEoBje08HxuPh1tJK/utwfI7hGH4emgs6b9s8jC8LN+BHCYzPZxu9doLP
1qnF9HFkuUZLmZgG4KfiQMtG3fInyOFnvrjzuph653GEEXC3lMpvStVEChfNrDA5
1CS+Rl/eKfa1ugiWX9dKWpkJ6azVWcqWX9Li1laeWt22mdU9PHPtXc4tG5875dG7
dcJWEIkvNPrUA8YLKpaLaP6vg8h9zC0myFCnSgrFkj/NIhzgp8dqpryPJ82bISIQ
1DsnhsZUVoCcaKG7aWxWQGyYXYrEtpZz6xecN7yT8Bu6tP5ZBANM/ic+8QxL0Yb4
AXGmScrumf+uM5DclGITKfyU0a4QAE1SYMgtBHzYZPKuhDc0xe8Bzyga9yRDqlET
Fgz/7GVMR4zfBRcsDB805S2SCKceqPnZ0BU609kLccc966YlIT/KgGxnj1iz2nLF
kf2FlfCu+JrmKvhNOtcF99PheZECc+ES+Xcjvgb2xQ4=
`protect END_PROTECTED
