`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYTKsWBfqLcBuVrWeZaXYC2W8a4zgeG0nvDhXttnCk5wikT5LvjHw7TEnoQP0yl+
ynaxffSHFfpZuv0+QY67j9o2sCpErK92u2SipYG8LIvERtpYRjzVoBx/LdwiFwMs
ln1DYZgBC4+Yk/V7fYJTsAsUFNzfms/mBksPvXzBlAaSor/mvJiO5W4y/CvVgaWk
scXUUf7twjLLntsJCBQONJZC3mvQnz9jSNCSdh9TOuTQDzb4meXEHYYuWtmogEdc
h1Q3iTuvf0rmNTx2llmNZc8H14bv8bamJXlomkDbqjOEcZFhfmOZknwEtqfhaJ/I
zoG2y+AD7EhCofqyfU3JgnUkGBHlKni7COiNN48ZKctXRcenTSVs281fcA/48l2f
Zssa7pmlzKnTacR1hyjdiYo11Yhy46Y2hvH/koWVdSyRWi1ZizbZueQNNlYDn6cy
GAPQcZ07Ys9ldFz9owWCLsAtrYaPLyH/bESMXvKl5031gJb4gASNOV7pSO5OHoTt
ZuC3qinXR+uR0mI31VncoH4EEwFxeNglu+rKuZAa9ozDOVEOMiH1azDwPYvPHkBJ
aK9duPdXUpM/Su8KOKExWNDGSHxc40P73sItieCU0No=
`protect END_PROTECTED
