`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdR0pvyY+9HE/Hpqtsx5TeOKKWbt1Zc/t4477c+RuAutopzk4vasEKLm9/llQ2Vx
qhJqaTcgTwk6be/Xkit76MhG2zw05oTQ58EgEFJgyc0fjK0gMUK4b8nepD6I2+nX
Zq0x3c6/8ynh+4J8RH2rKkoGTi2HPc044l9oXJtydjsDtDeHQkIZqdnVw4OYwqqd
G8jMCnv5Xxbhq2OlhvOfBVi13CyNZ1tZ8AY5SxiC7ceKf0i6/vrkyUj/urcb0wPJ
4AGS4TBPd2ba7qvtfPfjOFDrBgIeHX11wgMuEwaBw5tyyA7TpuICSdAelIngxTa8
czRRuXPeBf/3EMLJHsx3jONt83x1sv0i883d8A1kP2BZYZir3rMwMl49AQbJcY1F
`protect END_PROTECTED
