`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MVW1RcmhJUbUdiZHoqvoEctFvnVb1GbDOy5LadaL3OAqHfuLi34qFirCpFGZi2T7
NXFgCQHnd8QDhlTZng7tAI51JVFOipprtON686JWZfEnJQELCUZ5JsbDcFuX8ejm
ojW93GdMPRvfvunOAOt2smSH+7p2NPyxlkQGjMUCNMNcyYVftpqnNKcRsC75s+Js
5XXO5zslhs3ii8ksCnckTDC+GJ4YrEy2UcgqK2EGwvuYPgNDByHhbS7/G/OeluH0
E/6ejuvW6yjpeT9oo1DOBemWiHUqB+2Y4nR75NAydus=
`protect END_PROTECTED
