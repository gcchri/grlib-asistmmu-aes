`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+sLMHkL25MfIkdCDUs9srTbE3dfJLTG/4KcSLqR3Zq66acdpvoqAdTsLX6XwwKm6
ABOKFLHvMrvTXk5PFdEjJtupIefEqjHefuKde5ipvrU6fksodbNIWD1xRoex7Rrn
AzNyirqrpwuFpxdQJPLIl76hdSE2tGi5bpL+n0J3up5CA/hgWY3FQ5EnAAE1q8Qs
4/CXc7AVQf8ZvJA0a+P/IfhzrLpvZawc5xg20z0KnLbPb9cLU5KkaxfIbBZSaYlW
dwFz1HzOtmRWE+yTbEahJu6JSwVXKuOeFGtDSkxzfpz5bUDmuersRc6eEH/wjqRs
6/L6ns1xFDidAKmL83c4l1KXe4YQ9PNn1WlMM6Y28tXm97myoy0n8z0une6uVK6D
MXre+qkIXL3XeBj5gMLPBZlGw0JcVYPecwBXm/il1+gwdS9oz3EuYRhUhL1X4MZD
xr8T+vTLNwwdn0wQFIqXB0f/blbL2hndsI02lYn5z69xpquJbAIyn6GO/IjansDZ
VRioYUDTW7UnsV/Q04ULcG2TrXca8kRY5JGbYWMpbxBG6lk1bnr9mExeRd2XuzKb
a3MRgqEVpIQrHGbvajc4CayiJfSMyjU1GPaFtmExQRKL6Xp1//oHB6PUYJQfXnH0
hqC92E0B/mgVIk3tmOAk2377yY7syYJKbXlqkjv/c24y8SwAge1BRHhPWHFyiTnt
U5dG3B7mC65TuFlv8DA/A7bij11lgG5fs212gCkf9UZUAYOxYYpPLGipaf7yUINN
X8p3zBKO6kz728wc5bMpK8alOSau80uneB67Al1AlboeuaVWTN09GhybYlwej1oV
q/tYyKl4UbRkqHxJFM5DyGNWp4Tw1H5nMtZZmFXkfFx7G1hlUeDSlnrt8jrqcHaj
JpIQlPT7q+q5cn+lf4qs180+BnsUmXYSsPBp2sC/+As27OeRa6mok6D4yA1YZXUa
edF4FVM/mg3wnbQseEHp0g==
`protect END_PROTECTED
