`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61W/hlI8FLwRqG25OzI2FRcyCkyT7O60BVi9nrxsDzbflgT+5iop+ndB3cMgn04C
rBfb4liPruZZ8W47bESukpdcLYrOnro6x+J6OEjEtWDowXWYOisEAqVjRn0a+Jkn
wjyB4dABZS1fNCSVQYK7yTZjuymBndM+ly2ZJAFS9DvN07jeABWUHBn5pJUHegFs
X/aZVtNE7EMpJZe0nBqpzGoWVmahqKKmgqXxEMsFK47IiY5qRtAg2RiZCprUfOks
ksSb6npvb+g7uxHyj2ka7U+UBFlAhP4HXB/McK1w/LC40es+gXkx0r8rHEfsEFSS
jvJHtOGE5lyxNoIzamgs7VSUlkqNpT3JBqGlg167k+UC7UG/ZuUVzK7EgPhny0X5
Ik9q+TzwVoa+UP7qNMCwirrech4bNO47waP147jYQ+9jDo9uSz+P1n/amKSkvn1T
s6F9mUmTMIROkQEzLKGakUUS6gViH8e7Rcgy3tdU+GjUmRY4YCZTHFSb8hG+ZQEy
iYsvVOp1HRHD5P9hkzVijT80RHlOCyDLa/jowBGWKZiZ5glflM9Geufqpv0wf74y
y+04z2fuxMJOVsTvCONmeZR5lZUvKtDOclw+GpTU4Edaw0fg/ABGrtnjcZhmaoxM
5/phf8q4Hp47LtlcWTbuYswDIZMHiQpifvaMg1SWtlnnmDfcTb05r2jhy+ZAcdyc
AD9/gixqs/w4PybFoigAoGN1WIxAJSuAMvRci/CxMw8gE61aBwe5RZ/el/MR+Zsk
5ZjH65icPhAHPNMnxM9N5rs8J6F2HZIOpbQx5MCXYA+yEobGhyVyFttx8hPO8JBz
KIQMaqTZGUbejb1C4lOmYjZnFm7snfOVuK1PFzgSYDzpc8IgvbtkTONJC6P5J4cA
nI4CdWT3SSj7g6OQJC5EwwQw5r9IY5+UxgNiO8OJjnIrUcSOwWh8erQeWqzFukO1
BtuSvdEab09Qc9SHuHBC8bqnpD8KascfjXGBMxgQK75M9MN0xve3gj0asWvQSwpc
fUPbguiiDdPu9EZhUpQubrB+BNrEHV2t8FXZefIqIQXYJeGxY7r6dhpAMrvTsbEc
BT5HcdTo1b0FsRD6s9edKF8Z0Q8w48kA+JhRI5aMsGoM2Ju1BizmsuWP3/xTd8mD
sad0L/ea8tSyCyulOBOZtiBRF6OyaAWAGNjlqJ/Vhl4ZvYogRf3CekcrUaRufQNU
quTlxZ7ZoPuVCxY251ltW7qrxUOjnhz+sPJv6XEsdA9WPD+H4rEd4YXdg0hozBKA
XA0mUz+MP9KCloWrV9DzYS4ODn2rKjAh23aNDsbUqtNiEm2QMWdGVwi64buGg9Gi
U+CEBOwj9opEhakpAXbFOxaJHqG10Lla2VGRG3xEJOqIsycRRCUIF+9nJNZX2vEj
09YN7V+2xK7Il1VrzV3jNYpwsAhJSYkvenKlgpZv2tooFCVz1SiRXG+kiUI5XZ2K
CLF/1X+Vdv36Z5uZLGF7LR+cs2p6AvqXp+xOFgRPxLXxXvq0YSeb4uRr+hnKg/Cd
4X415CnhLvOSZhtu5eM8jxU5CUpkn7dgmrTPV2K6LnZhuHS6Grk8S7RLQRpiezDq
OH/zKCc+Vp1DVHUorKYOfQYD4VkxupCtKFmHbCrQ60YWyxOQZBUqIkmjCnCkhMPP
EF5/9Gl96IxHiAIIf63cLNFfg8ik3o/ihlMe2f0im9ncZGF48M/2ChOrBCxg/4Rk
2KTyDVECqABdBLZjMMFugCY6cZ5BZZBrvvT3XYLaaF0rlUupmXz7O3H82/0BCK3H
oxscGOe2SBmAXwJ0K93/MDcK+ZBddLwB6E+hX7Iaxlw2VL9tlLqZgVcS5hqr08/h
SMDDaeILzYAenBh55WiecNIMMdqjRldWCAaAjMhlwilK06uD3diEJqt8cAV2kKQC
`protect END_PROTECTED
