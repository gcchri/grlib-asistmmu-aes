`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkWlKXV+AQ1o8OpPzPpJcZAsoAeuezsSelNEesaY3j75D/pNDXzxhf78nxFYJFpw
OPCpxP8hqroXFqgXOx5mUC20kF0sk4b6miiHCy8lJqGOXCAg/WU6mAN2SbbLWBHt
PprMDbhSuk013YIcRKwhdWbHCECTjtl7xov7rpvotlWeuhiaxdWfireLYFNP90WU
5bvohCZdVfDxclIoeoV/Bl6ow+mjOcHT0mtYQSWYHM9dlOYuwWOxDbQQycLHof89
IZSNKZ+FvFvzKwXbCVTHmEBDyjJFU4oPKhZohBZ9FwUT+cQ9sbNE4oLIEvEM9ZTG
y62PBsGmLnk5FSLdzsCkVtP7UYXbFGdoa565Y0YQLjw8UOH/23/et/lpAtOoz/TG
KDyhzmqXhTnYgMh0ofrplASoX7jktRRdR0J2MNNEhi2AFKgobsIcjkPIwNONqjuX
QUj2YPsZ6QGNcVf/U/9EQ3ePkUF9rVVNQcJwCiOdVCNHRupZ+4XQtQJ1h7rogmfw
m/KLWqm8gQVvdYF0m9PArc0ucN2fDoD3oTmIoSoiu66BsNP7sM/OW7Qa2RxoaYMQ
`protect END_PROTECTED
