`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1gyNbZPHz5yYSCIHRtV5iRH2HFFnxq4bfMiTL8lVC1s4FNpIzY8Xn4ToOic+d8Cn
lvrV0Wu1G4yo2W9fbUSu59KvSJyUJhQMZ+jt1Suxa5wyX0E5w29Ewr4vl60q8Y4G
x6VgKYiBG3B33JABsnBsy9qz8W/O9h6Ys1rr92fg0WOUHWrwNrSD7DMxY1PHeqC5
H00GDH9iB0A9bcJv6LZayx+JuoIWcMllgoPr2db9N90ve3P6WpE9orb5AZXQ1MOv
c6eL8TBusRxTj7xR+Nj4D6b1z5D+QutIFfXXguzukmxwJ90ZtwiEgyhB+ZznsDIW
t0kpSIq8Mi84XSPU5234atgYSgWCWT1zJBu+50QixbAx4+xj8GbrWrSIPZscpuef
`protect END_PROTECTED
