`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
weBBoHKzdV1iMnb8/WQzX5OKkQHu0pnOnUpH8WCaTFn57ygXecNjapsaVBvOrMP9
kB5vWmghbV7sI84DEYdcQcLuJMYiwYQWof6oNrLbNXbdiGs3OhE/LiRu0FFKHJjP
Gq/dbPoEYFoUHdJQjXE66qmSXLmLfd2LxWWinAXde8MEdI1bIe57H7dAbcVSlPlj
E83gNJc41z+JFzTTn2WJTQco3fzm0KMHpDbBphUvohiAFXoPOMPTxZcCxQ20U6qT
2DfmXIrjjH/sdLaO63zftW6l6jf0//6FlZus1l+vu+/Xw9TKFNcRKRXeZaEJacMK
T1PHvCyXKnkkj+c3U4au9d9vMSDNY3/EapXtOKrJugFv5g8EoCcsKpe28s34ZPfR
7/IVaWcCvcgaSN1nnDw+dgeZpX1jbkfDw1vd1la0fQabToskQvX4nCJR3wMXyLgX
B5iMlUUgTKkbBakmpJUja+WnwCE42Va1U73uW9pvl6DE9nyGtwKs+yqcw9wk8XGH
Di9sZF0tQLgIiR48r7qsappM5qDliKeg28RMLyT/urOCJSzx30YpEgvnpX4FxCMA
XhbTGgyTkTWBcJ3jGELnEO575zQHoXuUlIYYwRt1ms54Cn4PEUu/U7WA39FtV3Bw
2FWRMxJId4rlZkBOeLbFHA==
`protect END_PROTECTED
