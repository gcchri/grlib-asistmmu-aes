`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sp2lCEKa+/VAhrUp12Tuv6r2AAVfbhHYXpSfE4ZuDqnD3yT6xLxI9A7LnU+E7Pue
DvZTgo4rRbAm8MFIFu8W4spivdeXLy6PTlyRgQterFl4sK3n1B+6lhrO0KVXPVKt
eKLAfkPYjpMMsu5BdgJ4Qo9FTAd21atG7d3FdmztvxD7iFnhr6i387rOsYK3CpdY
6XGtWGhcWxLxXJoq/6iDrMEoy6hUoDw6qP5CAds8OPBShULPy29sph6HzlQz7RLM
VH/0Bww5RX9UIlcAkbZ297ch29nCIjpbZDGjGkgqhng=
`protect END_PROTECTED
