`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqx6l23V8H3UR1oqJo+A82tsiblPjolin3p3C1xpA1cOzxO8pN4zJ7lctROvso8m
fNJeDNNB2E8O8bmHjzQPJy3aNFXYxNH+pyR+CilQduNgBK/A45e1zfOOR6RKN+ay
fiSfxWDZ+SulrXvEEXI5a2af/TnVW/vAKI8JyyoKXBz9StTLmU4K9aTQffUTJJCO
sDDBptMlJGJwtY09d7BQl4iXuM4AfAMFCi9FieS5yA5raNi7DXjsCawoEw4KQLNx
EX0Ksd0GO+k/nwL9G7oY9DhAQJvj0WLWkAL8DbK/F0YBi284qQIBJe3x/l21Nvzm
2Y09p50Y9Bb+aqdpK3VtZeA7QVHnfAHvuZrlY+nrlOFNo3WiII8TvjALb5gSDjLr
7e5gHSqsxkir7BD7f7njbC/VX+fyRMw0hvgyGFkqWfO7x2sGFtwIIfZ7TvyegM13
4JVICukwCmiA3+Fu8pgxpfEbItpxMu5QI93+atY0GqN+caatOJM0tq8L8viocyen
1s725YXjJyLEZFmm8YAV1CPmiUIKZx7NKBPow7v2D5RwDARA6KgeS67lCYrDOWDF
UMrx/C+QVfuVgUeqEzB3sD3iduhbe7N3c8qT6dpRb4VkJMK03tVNHqSB7IDeNrNe
t5n34r6uckqUR9WvY5hWxWgJH6g4Yqos9KUPco1Hs6BPFE2ThfCdrDH6i3sf+UVZ
gsPkOuM9Cjp2MudC8oGYQ3n0RFR//8D6oQVjH37bICG+EWvKzNsyvlEmAU0QD+PD
JGLixnk2S+EPjs9swRFC1Xk3A5od42B5YDTjzLdq4j7wY8fPpSzdBuQt+EdRsRUv
tDvrhCrpvg5rGF+t0R5/dMrf4ikB32ElVGIsLdIhpDQmZv+8RX+kYXkNS1nyZilm
/nslGjBxcfry6Gl7S7WafpWZ/om3orZr6TbwBg2PTRD9ekY7MorxTNofK2Sv3hu0
JeMbiwSWQSz56XNbgTIcugz4YXGMzvLnNb8W9lE5ZOCqaDwaGF4tGAPl7r49CbRQ
uBTheMLlka42u11bDJkScjlrW5zgI9LkTWkVaJjUJD6gIEL+RreecAMpOzyx6E1a
k3+3qwE9PXx4ZTBg9dNfYojDWf2XhuJwRdvVtnwoE6hoIWwEh445LlofzH8nAQ5u
VOVElW/Qhn5gZHoljYPa2/CKkG+8rZYUPsnd5VQ18+H4LLrHLz0UC269TbjQtolR
4O5msQLV/Fj1zvzfwqnGMP+qjY3y4OSbw4ikuP0g+hKaiaCAtrIrrI0mkR+QoU/f
qxq950ER7uWUQjLEOYa9g8Mo7iOWEymt7cER04SR8jpkqqJ3zy/vVJQ3n6i0/KOU
XDp6u2AZIibFRBK/FWldUDT8ndO71qKQgfxPToyjih1MrdNLKryAQgB/WK95+hgG
QLP2XBbLkP4jXQB69dgSU1U8MCcbl70huXnq0Ec5sMdZZFIW2m8amm5tI5j9QI1n
QvEjPtk+NcGCB/hjp4pI6g==
`protect END_PROTECTED
