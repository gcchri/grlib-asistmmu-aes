`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1G4Q0WbnaeKPGv4tQK9dZyl9wdbpz7ukmQDMB93pSoQsvJkNcdpTHK7tYA/Z3H9U
uiIvyeYUb4v/u9PuQ06f8LhDdPlJLZCRqYUdpYdZEUB6I1O1zyWL366ve673UnR0
eBahNg8QKMKbxBK4XyMaEGuqgn+gb3fOHenZhYBh6IxknSrWkXc6SjHh7GOnrrTE
Loak0cBWrh9F1hzHqpKILsoJLz5UzpHIjFl98hcjZ06H7aFvPDc17e8Gy+ciXqv3
nfYT9dV0sJNHT/82ydEiw6giZzUrI7MGAXtoZn0TGS3DbIsj/L23RvjP44nJH1qL
n2b7+67MWUqduCoMahGnqXhv93E19F/nnDylqkOmuRxexE+g/uJinDW0u0UvEh6c
`protect END_PROTECTED
