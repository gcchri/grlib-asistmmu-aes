`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWcyBl+PCiFiEvfTLRumEdkoZ91Hp57v9AVAnSYuMuXIX6DKjIfDejPNCSZubiVU
h1Smz19Yi93uc/Uzw6j6P6bthHnnGi0NhZkrUleyOw79EVoAcNhewXnwTY/Uyoel
5c9YZ8KzrfKCj4KjQ075zzsT+oV+SbyEntXEFnOzZMViue2TXtldTlBJVnLp7mCP
RiVdg86kjM/CDeu12Hn4hwBWCQLtvoCDDGG5RyvCop9r6/yr7n8LhAdb1WDfEXIm
fKWTmp+iSF0w8yS4x2ascgQghI4ZUihUyRgfUcwmeXYqtayqBgqXl/JG9l8N3zTn
Vgb5BuvqKPryL01aufG+1MVHLNIoi4X+/r4YeTgE4SleykIScA5rwnh0wMDr350i
O3G0hdvP0sXj0QH/ywYi0V5Xy0QEM1h+3nG5pDb2WjspXv4qpBKiH5i6IoOKYjjo
DsPqVzy3iX7bhyqtS02E2UF4lwRliKa/MB5YlVCZWELSiGTshq+Zv14jBtEMXRSJ
`protect END_PROTECTED
