`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ff2RGjA0TZJMOQAQLk+c4L7lgf5Q4qE1gm3vKtOGnSgBBqAwue1Yfoe8MOt550Gt
OCazlqMjUIL4LhETz7URT/Vx5Ds0hcqLtFTUsQ7jBUqJ3OxEZPNUAC4LzMGSZpXS
w1LOjTz5V/n1z++ho5M/nm7ekFpfoZjIEXUPa67e0yf6qFne55qi9iqfRU/gAEL1
/Wig1bo9fSkhcdswjxKW7VKgUhAwv+OTVnMjcDiZ8UZ3ywXt9aMr3Nt3EQpciTOL
Ra+hE9w/ii446P2rOfJWy0cC1jAZeH34f8g0yRua83ipdQsD5WRZIJZ51eTQ3rij
AhOMiDyEKR30pRsFwzhEtElKbz5WcOF0UN1Q+PY/RxsYO5Lnhjq3igtMlRbvFVYh
HwdKba48O6fN/H0pAVdKe9ZKrUgnIQOBUZ1BDRQOp1sx8E+eRDpypVNchq0icIvF
7GEmz0vRf5evkBN8rfR1Sl3zLUNPOyZYh99Xw5ZUMkYshilHAdx1vKe6bJPU3F+5
`protect END_PROTECTED
