`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpWtshUww5H0PTEuINQ8brnN3gqDopzFfNFTQRtERAsx2Or5NMa3lL7lKl9eiHi2
nsrA8Qu+fUGcGIearXDt6vO2GgqeWpAzO1UTPBt000D32+ArIsyEu5ClyEcMT+Yb
xyOSjk8OVLYp5MR37ofCblaglmSgNytaFWtK2HC7n4IBW4KaL1XXdT2EGZIcdaZm
2UjLKXzYvf3xmA2y74FkhdDOsU2AwyfWN3TeDLEoOfs1oRRs8HfduhFYYTkOmzkV
k9lG2ANZXdHv5bKAFUvzT0h1gZYl9zkPdlpkbOcs/7cN3HkzkB8MFqA28KKV4xdn
pkTl3tpC1BHwCNJtmSEzvRbK2tml++/kqSgBZMUoFwNQ6q+TqovzwuvnMNIJLLrR
75GHUJqZG3WIJC52ylC1+PjFL1jfvWtZcP/WM8X0Wxd7E2FtBo9wqGjmcHNLkgaZ
HS7YSGWw3NMgL/trqX2f9PWLTBOjzfDOreEFlfDH7m30zIL3EvODPRtWdzzSt7NZ
t/sMAPDOhg9MHSF938rpr5T7DpK5mPJE6AO/7Fdk8dwEMSm5C4+8DQjdUPUu97xj
ykc/YwhfxKmVYZXSRIKdqlePqJnq7Oak71S91rkEU+Uozh6IuzliEJXMDW44kVbv
dwiu63gSvkhfQC7D2+4sUg==
`protect END_PROTECTED
