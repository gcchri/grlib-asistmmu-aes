`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VIg9CRALhzkDMDM+NDTpKWHNckmhQIInrNbvIP2Zv8/endRaBkPC3siJcgMfjQGq
ioOk6N10nkW1BIlfBOKUVG93pomqypu5viMgN1IT/WzA1iQp/oX07k6zjBDG+Tl9
1cuHOTaRDIHjUJWZQyyhZDbB5WvQZlR+pNO6suLNW9h/322F4bq+sDDvDN3+Aa2p
H2W9TbMDFOikwwjRn28P0G2/x0vRVuXKMAZIk74DltYW6qs+Rwchm5BFl3OpimJn
CTBSd5R4olzZDHyQSp+N1gK7X1PS28dgBYk33B5TfHoG/UPjmRmGrX0KvVOuzADA
a+/+F/tAMS5i+iK9HaEdc0TMGFcZQ6bk82qgZk/iqdC6tAa/cpmNslVzc5MgIEaK
nxuHektocF1F4jrSamQQvw==
`protect END_PROTECTED
