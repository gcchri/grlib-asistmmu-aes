`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uaBdY0aws7JLx9YdrfhHISFHDFh74Cicu6tajif2fNFMpDN2WQFjWJUMi+pVHBU9
ABuBbSm2ehcs2n+obcKHmne4N/uNeNXzv1ixvNkfLNPl6oD6ZFjrVt/XRv925oN+
PjSP/PnSjxkYqvToNAlKKGElb+IXAkp0SsH9MUQElMfGbtkdsvn/RWad70YU3C1K
BtodmXQRDr4wCH3071Dd6kfk40sDJp2dkrWaihx11+CHyu2QMgvglwfSk6jeByUc
4DM2smsH6js3gQArMXyUPTh4eWfX6Q0MHEmVyvaHYRXURRgkUxdzwFXBFt99G206
e/Ra9fizo1JsH2gUqbmAMOjfH2o/NFhWeMHhZxj4G9i0tgeY0q/7YK0xrm6QRvaK
draVFhhjTRMZ449Idds4KayHDlzXsZinRjPuX3MKZlARZLktvEtVJ5tcBmln5teW
8BknsYoBY8jVYF/3ics7nysxNtvlqIavkE266lO9joYNCKzCizorqflwPxr6WwjH
tT3mk0QSGhYu5oVbdDsnJyyDI1B3Ht+/VphDhas860T4DjZpxOxWOQ8c3plRJF1L
/B9Ln+HOL4359v1TE0kR02d1h2a4/djDGe2AuImo2F+ACFtocJ/iUuX3ya3SQONU
lfjn0I+/Y7wv1K76B2ItGZrbq8agdETn5Ye1InuQUwU=
`protect END_PROTECTED
