`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qy7oqXlPEzJaYtkxQS5C7boE1swoDeq89VSw2Zg8f7210psITb5qJCk6IK4Y6ZN0
PpjUjqmkXHFJeOWiUI1j/9F65yQaubMyBMKZmcclAlCruT9esK/x26fiLK2yMQ+R
J5izuLj9yG1HEvTTq2bkiMQi0SxUdzWkquN9asiWuobpdH0X35n0iUcw77gTEHhO
IGZ4+VQJMlg9QDUcE9b9+QqZ/QcQ6kSVjOic1gY5g5iMOok7vOEu0zrGZz8R3TZn
MBHdAxkpzasSt1KJLQd3o2ttmmA5t2Sk1Wv3Tid+2Ld5NCKtJJe5mMiyuduNHYp1
KHpHlB9WopqqrFo9+pikbBb0Gy8A2gIC3SSviG9sjaGr0TljYW27MAFIdDT3X1WM
YQZadolEBcH+Tg6S9Cmy2so2CCWefFp3oZ67d8wFvDiiKUvSC6GcYF23OOjEhF2G
sf6iNCDjskAcAjjsePguJSLcez8jMZ91RoeA5rbpuMhY+qp9GJjjhjAGbRUsC7So
D5gGOYsIY3mcMmVIN/vVCsPFobYv1ujxauVfyy/zrn86AaQdycc7+PNPhNqEwzHS
GjmvJ4haDlrdno5gK/RsUf5o0mdInpqTJrw29YcfpARnPWLNjaH9lqNJmEK52nYk
bN7DJ35MVYXWg5R9vm2KW9zp18W4mtK4E/xtEv/OcQ7jFfNU8CX1NTQF1bHY4YP7
nM0e+Gagt96vwXidA7C+vD2pXa7YSVF/v69b9zA7TLT7qcK2ByG4bGaPj56ERql/
c74wrMdj02baNcD51ZfwN/OqsjHSwCu0ZFpCZFDp5nwhqodcGk+7OoQnwly0vYER
2OA1ZquOLrfWvPCAYtt1igA5Bd62ITqArVCweWvL4gbHZmPVdHRGwpKSIgztAa56
C7PAYCnVGcJ5qfm8ODaPvikMqI8NJ/Y+0m/Sr7k+gZRvtLB6LhiODpR911e699c8
Xxcj5tyDL3kRXaBVJtdUcp8C54DWPu0O4NjU85f90q55mlhNDnQcgv8tY2j8uKpV
s3Zsfy14W6RMkKeG9VcmMxVQTKbFOIL9jMZvMHisFh8bly89nGG3jr0ISevLeZpJ
Gb90lNHvwhLo8W5h+LvFPPiPUrkRKJVYC+BwjcPtoXNoTqNugP+9+S25IsNbDmWF
WwyIBRje8wYP28GQ8KmNYFAbW7fa4eUIfNrbOnuc733jegMtyo57In10dQSlFhhR
hi57Tn3Qn7Z6gePP6D7ZhcFZzMLrD4O0bR+dr7KTP1lc/wQMDEHPBZl3eP3YtUT0
Nj8GM6LKhE2dQa/jwRl7LewwvMSkeUPmZGiaDtab+Snz6F/+Mlbdp+dfGZI/T37P
Z5tUWupQ7zSF95J+69PLAD3/QAhpji5GGAJfABFeud++ZkslVs+l4nCrqXzydhxW
NYdA/FGqUcHFTGySf7todSF2LNNfvNvb4nLOJacASKN2xkLhQzCuDd7OoTu198LC
Zx+jD0pv2HgQwkyPnkv4sm/ibLGinBT2iYmjd5EoK6+sChAHWc2WW5jIbeIbRmwv
8/dLp4Tl57xei97d7op0trLSImVGG2DawOqBvJWMOON85jtlLhULdkMlhGz6cRuh
PV9UKP7uy3mUlUSveN8vtq0IgQAdcVCODoYuobdkR+y9NhOjXGDMVGgvskC/QzpF
SfHbY38t//6/77MnRR6zjW81/ljtMVbA2cx9f0A0U+zMAlNIUZPh1IlsuQ/qr9Oi
P7nKPBNbcy4rcM50ZRnTioExt3cvt/m7+3YvdKM3G7u+wjRd1BZ5Ma/pqxcbZfOD
lQ0ACfIHxC29hSk164mR07WmZSfsiYBNiiauQxyFuR4=
`protect END_PROTECTED
