`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iy67ptq8xRkmgWSaeqlzb9A4vQkgOgrdK5+kXyOZjzA1ablnmR/kR54HEZ9wWgLw
1tA6KLeKB+2boIwLqogOnpesidgcZdhaax0WWv22HpDBTvLLILctFTksHDNqFTo3
gNokgkdoWvjg2XcwPDWx2/5uuceWiG6UZpDlfMFN8npt0AwLEnaLMbE7Et0ESdUu
ImC9muzMc7+AxoR9tVBmYSn4edRXtri0b7eKvoLBkR/7FcOCDQHLMQlKdMYJudwR
oAMefTD7Hfm05zBGrDjoQcUPRdZGf3ra+6idYLDoUJu7T9dwl5jTFXzsEUWOsUq/
Ku56zOvbSs16VDOyplKEcW6uJrDv/MAIPz3sw3atwO6R+gWDxPveNepurG1TCVxD
sTOCPK9qsBVWChAv3XAfMPFdbXmsTUjXMhWVpQIEvzvYD+kAzWSPo81lVukuffyD
osLcKCDiXC3GzVMSijT8l6OXmQc5u/KNkvKR9lFP22A=
`protect END_PROTECTED
