`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQe/ZrSO7rxkwnuYYnGPf4vHpJ0cYd9E/bwvKzAxTNBo6/t/XuDWBFjruso/0gPE
FhSvmTZ3tvvwQ/aZdlq/+03EhIwLLRnE5jhJzr0WTg54DHPMdLe0oFlechrrO6Ho
lD2epaYVzhCBko3L5EnCVuzhzLyXJUynlV/kPMcKwyWCskc432LZhXgyTLY6W5CL
kLDgSe5EW6ogby/oEahaG4mRDrwI3jGQVY5ScSQcLUQ+PWCUOqedzWXf3JdufuTZ
Mhk4LoJZOeONjhCW5VAf7SAfbkMtAp+Rdxheya/RkGlDAHTaichvDrCBiClzx/QP
bg2+R1lSgYKV0fQw+kWjTrEuSWmJtrba2Tqm1HYc9TCJ6jl7pTN/6Pwfuwle0YzU
6G3NeO+pGRq4OFGJtl0pDFB/R9WBQJ7HX84BSkViX9PuHbn4reV0XPqxtN7dbkYa
FJzj/i5pajNC3YjbjnTQC6nVeLpEdJ+A77OLMJuxfgjX4dsWUAUb3UvfX343LKzH
2y1dEQluFEscAUBTdP1zkGtl240HnBH0Gds/rQ6M7/mDtHgmwUX0QhFgsz8b3a78
w+HsVT/cDU/gUFnFCzcA9B6Pdv/Xm8etLQVYcjvFMuaE57I3BDNYdDFs5BqNtkrG
pgl0NqzMHVxGqH0NWaa1cM3DQZJMUdktNnjD0fx5my6KS3Mw+9cvYSFFaV9Mlqoe
c7gKzRFtShrlEXtM3H3mOSO8lFNCV71cCiTG91oCUIUh8mk4NcZ+oQ+QlYLdtSaM
n9fDUzupORg0e6/So6tgTQ==
`protect END_PROTECTED
