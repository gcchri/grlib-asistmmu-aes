`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCLddk1wcCwma8+H6h2HmEvbUOI91wcv9bkY1dxQzU1fMHa/wOO49MLJSazwrAuI
0PbSAzAFKr6HONgGlMHt4KUcepQvThD5/ic7uQQvkhkz9CpF7akMa7Fasc3DnC8y
H+ovPwEyoBRF4U2t+hvlwEsLI0wtUCx3xS+wcmC/DbdlOqNTQf8TtAmQUsIB3nqC
ZoVD/2rd8YqiR2PsS9DsST2KvWyklWJtzYo70hWReb6nKpz9q2ixIzGAOF+lKaTt
89If3i9Eqs3uW29fgXceoJw2egnJql1vDDbYZuSv0APqZi83sGkRl94fINjgnpcF
tTYsBy9tcYM3dKghN+iFsDYPz93FOivC45SII2XxJYNL0DQTpRG4nv6i2D5zKX7l
/MJ6wavqUKr4Xu4UVY2Fr9A/e/+waykK3O4hl9NVWq002eN4XoarckWH8P+XjBBc
lyNjyFKYv5PHiXV14dgEkw==
`protect END_PROTECTED
