`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yIV++Wyg4AM6YfxVuhRMmD+1j4RsoIUxNJxIHqbL4n88ezCcemAD7Tj7uuMMblzO
5IRGnued7lzsLhKkJzxuD14d/aE+ZpvLaDsmgYh1Etsjz8axPyqovbDYU3k3CnHX
ZoOpvieisX3YZLjUq3yibUiJhh0vV47h+f37HZJ0gM8GYpp+IJOTtJvp833VZZhg
JpgdpXnOf9mBYImAmPyKb2BMhGwjF13TWhRuvQLODg0RBKqS7v0aKLeILbLLLqKZ
/bfXkrSL/AJ9N1FDu4J8We4RRbRroS/Lng/sJ1QBerizrRaNb8mzaQJqj+8D8rDd
0Hon97pbYzsfie7vt8uANGOCqfHNnPdILXEmFRlOY6oaxz4FLmZbaZ329JjODADd
G5TxxmFKQfDcMLkxWg2+DpKsGIr9VQkAOak8VaVtAelscDZW6mUyVxRPGi9mQHss
KHGdXxFIHF5zDAQRBQdJD5LTcmKZqz9z8uawdkiQbzeb8zAyWk/Vuhj6LXS0o9Im
Fy0pT8M9ZZB9xUcf/uyhLbCgKRx+SogtcPmVKLxMUJ5fQ3tLAUlpnu2dIO26fmAB
T97bmkpKl0XCUvKwVorzkiN9DngfgvhlKQCkxAACM6F4Ek+J9Tw+baDyvUwbM+y8
5kz4SJGfV20LxyQkf72SOSeIGEAb89oq9M/tlW7dMYDYPnX+9+dalItQM3q6fv4N
+VceZ76HPRPX0oq0TCWWnQo7G2eTRST+ROvAMA89AKdpxrc1xco7aBOeScfHFIiC
UZYO3HBpAcYq5z0sZYyX2hs2VghdxwMfQNTMvsqyfJZ8w6OdMPCmNWy5zZR50ae+
6pbJnGPOXlVBlUhWEHvOEX8/3sFUS/i6vG5Re7kUcSo2QPdqzeKfE5NvwTC/8hPc
1O/PvoN124f145Hyr7yIiddm7GvlWCiY77icYamNxJU34JI+5Ka7d7OQtqfhrjlU
FsD75w0K7mCTbpVvPQgeneO4HWoSBPAOX6tc/IUIHlbsk+oYvAr1oWyI4X6rVSqs
teA1fjwSgRpj8+wrKXpCdp1+Zm8LvIC6yG2Sx6FJxQ/qrKMa139LXpbBW05BDCVf
l+Smq9rZ/mUE3OIn6swcvSewzMXaEyi7ZKwvokKTlVQtoenPY/YEmR0ZTmp50dVE
7f9ccWuD01WxUonPVSkuD/xWuWpxxJnoewZg82e0ebTE77THSLcgq4NBM9Y6MRS6
G2ve2AIYupNSREhGRWG0Z4lKhC7aon5N24zsMMfd9vPQifFWwg69uirPRcQMbJ8+
`protect END_PROTECTED
