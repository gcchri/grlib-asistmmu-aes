`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tPMpyCq1Nv6Mzucho0275Paarf5AyKup14uRVzfFpv3tOHu1eo8W9w/Kgrcil5S
iB4zOKyXRiN6ivAIawuuufjatnchW3yqZRCkcpUFpSVhe8Uo/xKUCf3AOVPrs1BK
n8QRt7YSagxdTlhXUgbnPCrlCUQwtASf2dXkBtYqCQm6FzXZdZUR6q09wPDNH4Pt
9EkcbBUMbLO8PCnsmT9GpiDuhF+bU2F2N4Oz69T7RIaB33LObAJZ//00K1Cwfrqe
lVSMWHQnuIdgOWNOwNyXzRbpPKPFAuaq26zWUWA8n0kXbxKIdtH13Jofh3E/dODs
U/vQbnIOVeDLjAz6p9XR8eCS/FXY3ekOCuqUv2ct+2FUJkCNZ19SfigXaJ2JdG9v
eBx/MWkJ0WmMTsgdksv1iJpTC+2kHRiWdno8n2gWib5WYH1y8DFlzaMDu7rGllS1
EsugdjiiWyJCkLuIQ3bXMH5oKQfp5zldW2zYu8Ya9uAuHUPMjWSR/4WW0hG6b6AW
dhOg2xsn/uxUsWE3E2RpaacuHrE8YO/YrMPExXFpOtDf6CG/L68odDU3JKcGjpTD
/3DO9ndu2l50JCdfjDnXGnhSlSZhKv1MFWliHwfLmX5+bRsuqAYbFECmzqui0xnR
sXp2YQh+QAPloniVZxM5G0Lm5S2RF0M6TtG3Kf5oUFuRjr5fr0CxLFgNGUCGJV+X
JO+wJPxImTYl3572RwQp6kYyH7ivEVKgOYrilClo3S8UBXSpNYrynz+bPDc7+SQW
`protect END_PROTECTED
