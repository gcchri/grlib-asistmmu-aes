`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JcEedGGCo8bVxt7LqmtB6KPs+tDClLIwfC95LzMnlvqpXgjayfQD6CzuVuqlFS5p
6eUIOO+O6RJRbM95Olahmnw3+Q1yzyn7yfZuhCa7OSZ3AV2IqLgU+p3RFgKynKWc
UKPLv9up3O7Q38ivGiTosF4IyhjlVdm9y4hX7swJSZEIFGl0e2dPdskJjaqMduPo
P9G2z1U7dTytVUHawAPUxjvBg59ieDt+Ibcz9ufG/R5Q05RXoBZQGLFnqpqnvSHA
IMYM9SivgAaxVOBDdoL+J/8iMb2NxNmfLeMXZ2ZxxZolCAl52W56l3B45u78HGO4
augF/ebh3KrFZwG8ZCWr/yVqIxQv1aB3iUmwe6qOwGmoV8gd3+WxETUf/P5hraLj
`protect END_PROTECTED
