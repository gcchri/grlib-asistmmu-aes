`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GxMqsoy90ubOfPN7qrrJLtIDxiu28fJ7hr4MkK2ocT4o9HNcniQT6lmbJO42wzWs
j5mmeMGtbh9jHAIgytIRmHJOu6wKr6FVcHS9MjXHm6F272L27Lv+tcLfNvQ4hZzI
cJYcYSlL8bH2kxFFEfkyFxgqn7DfZb0f5rSuX/f19aMJhH4Nen09GZKMyNIyOAY1
r+kLwKcrUV93i9wpF0jQsdC91c/RQJrYMZHkTZYn31apI8hHgiisJ/X73ZtV7LDf
DENZAtu4dX0fUHxhs0yCobu8QzngCalT6QwFMWKrRgA4Z99WrgfTlrAuM2RhAQZM
rIETTfooxazYGP+2+Vv5nVoeSn19MDFfq3Gqy94vn5q0FlQ1Z7usfLJBZXuFjiwD
Vr2VeGj0QUzvLD9SUiEe8rtb8wmFsSdDM9mYagiCLKVFImrwSQLxGwzX+Wt+nw1f
t3CaajlwL8A232BZyJWuRsSvBBut4IVrQquZdqOj1Pw=
`protect END_PROTECTED
