`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZ8hL+tUkVUi9L1bLa9gcaRJkh1Mzqanro/+3N7EcVw68LrPEcaHt9exB3x0Ofky
QLWTRcJls0hO/xh7YQ/SbcTDZ25PLLSBBgKV3jVd8m73yDZ3xGM93yPVyhw91tMJ
4hipfavMqpEwwlZT60D986FeXP+l3mvTTSO0huAN0O7IkrIokK7w/f727wBnKwjC
2pRuFaI+VLsZm2x5H8E8UZBsu9+uNxvd8XrMX3lmfMcQz83+LKrh9c/JGphCI4GY
Vbi0+HwVbHxZxH9rFUtswf/E45+BGWbTkMJOS4s8L0kZmsCk7RggW/AGITf1gYLP
PHPjxNWOTCEJ/LPyWOslN8iWJx15KW2nQEPuvKTg0YyjyxzGwfk0J8KGEn5atMl/
9evaUQcW8JCGafBZ+GQjHoYc4PvaXtlJLvUJ59WtxdI=
`protect END_PROTECTED
