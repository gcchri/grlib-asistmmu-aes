`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8y0IW3+fuCkhbl3Zif4f3XYaixFu9YUFXm6LOzt/7YIJzFei7HlxxTcN8XRAFR6O
bcmCIqtsYzR/KJPW3ewr28NUrhyHqrCNd5/lop4HdXy61nnrO9kFUpmt9Krhklm0
v1NhMo1AzHxbB5CQoOlfmOMfNbfj8nZCB6TvPEUhLS6bEEX8tVarZKxfQDOx+5Sj
Y3q6D0P6tMHGV8PC0FPiVHA/tsvepS0s6IYTMl4bKVl1n012wjDvfHvGavtnZoiT
LwcJsX3AJBtVO/efap6vHw==
`protect END_PROTECTED
