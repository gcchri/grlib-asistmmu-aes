`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10cw/9sj1jeW25iwWKkjqTRIe0uXQ0ibrUZ01Ou2OU5eJBSQHoUZHA3uM0JE4P3F
nvjBmziqnh89L5Nlnqs9hRcsbSSG6iYpvMnPF33Fyiw1jrCiChFZER4Dcg0TycCT
pmZc01136yKF4e6wVKCZh+54+13p6LAUkzqUKhYudJ1zdbZoDUiUnj9HY2z4F3y7
ODdLRRRVzx4gzmg0/cOcZl7309dsu668stikS7o6tWB7XntusFc9xZz4O+9GTest
lQO3MPFcr1bteThH0QHjo95EjHAUi62pceQb5v3C0M4thGPMdfFNxOKCxqtWcFnc
RbZE4yTI1F1PRoU3F+dWGzIB/mitQIssaLaob2YJAMjM8CROPWZXDC+k0ZSukvpH
ySt4WUE/a3pLZphu+hn5v4d0jHlXQHXEOcxEdV3FmyvV0M1ZAsPv3RpP0xoypwTO
4zl2VTmZLlg1Uaf9V1BB5Q==
`protect END_PROTECTED
