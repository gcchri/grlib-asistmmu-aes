`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jsC4alehu6VNjAL2SNW5XIaQawZcnzv+OQ0dSvVEW1UTx0gHnfWNhRrYtMGSbzg5
XCknXQqR4Uxpa4qELSwc4kXDcDNsXz6x/oQVF7CoZDr5dgkUiz47opQfjb9w4y01
1b+NzTvV6VWKsivNKzCw1bKzk/XqH37seEXXTc4JWVJTbUglPo3R5gLwzJQ1Mdcc
tjWQH7VifdFLG3Nc8TDByo2OcPjKXznFzI/1lt1la7me2El02Mmgd0ra3BPSiTII
fqVa66cm5/QJCsfUEazTNDDZre6l265rDojqeRYO/ThGgdc/6VunfHVy5Rm4vQsk
I/Be9givATMcOgTM/04XQwvSzakDwga5xBS2o9hzXrP1zLtauVRQcT4+v9mVTtum
DdroVMaT6KniZUt1dD0FfpWuhmREPniUIJcDV3DFwX7y90+zcs1rBLtC4Ldix6m3
n0i2wNBiYR+UjACxcUcWr7e44EH6etlze3HC1YbyrLzH/crZc8hu7KWZseinNyBO
pRQRix943oobH4dQhDcDtx2bKbRw7XLOscdKjZq62/P6I/XyWsM8mriXvYVCE25/
mFlrCkuIE0AA9LUhew+vWEnwV2MpAjK3+2Iw7SM+yorFW1P2EitS+dBM1IHSY5dj
s//bWju88UP6ApENio7QrfhA1k0RAXaCIUdHWXKjZgha4pgoyRx9j4BBJrsrGVdN
ehDVAmUBCxIBiynpCrqpIgCTsj9eRJfSV+HmWVobG5wUjrNA91z2+6IQr54JLY+g
ULnYpZsUxN0OWj4JScMusrAIPqpOs4Bzn3F5UzeWRNeP2EWZdFc31bvbM3x2tcQk
kpyIoTuyz5e5H/SicU1omg==
`protect END_PROTECTED
