`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BIPlzBtw+iC5XtPFYUznDian5Zn1HGb6AjOBPLrYoqk2XvQl2atGeYRt/hV6CTi+
noN37P9ipo5ei1be6DjgjP8C//TPMtSiQUMg9Bcvd9gDW3cSLxXPf4DBu/eKXz9k
hhhspt4kQvMk1JgRS+KpJfeIvP+s3PDru32bK3aSCxlKO/KCAnxpNck3IPeF7TVm
67kFrwrbZAXy/dNsm6sqfFiYmO9ElGdA+V5oQmVAXjDE1C5pemBdCIYfWfciBXxd
4kw36uBU40RaIkHlNdtdTt7l1AiaVMxcNEW5h9GPOMTGNLv711AO9ihmRbAy2bHi
qzzfH/yQbhq8Wbqrv6TExBJ25+sn7LfYiXloNCVRX8vIzrZHqeCCuJVtStyQYaig
La2SD5AQqMzExkxLXFioXvV9oneXNR4pSTguRpumKUmo4AFxl0tSK7c94vEAGpes
14m9eJ0nxISS0kEkJrh7OaaI/GZ+12jNQ2MFaei0AG2HBSWxDnYStCc71+In6pbm
RPdJY3rXU97Q0cE5Hk2hgwpb+30USRAYNb38KZBLqArrlZ/Vc8OObvJal7zkzAzQ
UAkjTWZ1oXVawiI6GbjC79i18Z7Ng+wRfHhgKaEaA9O+GhJj9nhCdziNHsTGhXc7
QfZC75doU+8qcR1RlskHyQ==
`protect END_PROTECTED
