`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5RmDITjsYkhuT5CcSj4gTpw+lvD4O9v5Q0cCkdmIqhfRkSouIWk1QRea+DNJbSp3
PdLy98yGdD4hdnUdWBwstEf0c1Jv/i/enR0n6KR9oYGM9k7q12QOLntlVGVpNdba
TS1DnEZ0BOhQSNxPJb87MvifvWG4kxSvidmSSFICEtuTbvSTHF3+/UQkcmW8o69P
MRowMt+h1rP/s+hEVhE+SsgIukzehc2JXqpZOx8zpOQAXwFyL3nAmRtuEw6xOU0R
UiSPVOvUiTiJ+E+sQdd6RcDmSwDadN0vyLxjq0cOAKvg/O6PL3sjjeecU57YQ5Pz
pR0Z+AQLSTKVy+ImQgAGIHERPmbhhJHMPFEabcKeWo4SHu4OOdv9z4nOpwJXqZQV
SWM0UQSi8RUQ0vHnb+cVJNyiJBieHNMBSbRUHeqYQJ+SCIyZaElI63m29aFkU/yG
NLwFCEGm3LsLnTK7Z/Bqpw==
`protect END_PROTECTED
