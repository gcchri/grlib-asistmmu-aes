`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y3bl6FuBK+ye+YXYxIwUDa3SRWVNpVQou/wRSBEAKnLvERcSXoJ6l3/+yxQ4+/ar
OzVq68rPpTRhRzDSci4zQyvshPaIRGL9tcF3b5DOD6pLUA2LuT5k8QGCE3SkSlr5
+HvGdHXH7UushUZRrIK/E2QCO/J9RFJRVl017oAH13P8KIoIhJ26JFuztr7RTgK5
JSDEBLoOaqZ5fFEDZNPJb5/Pdv7hTVlufBh3UUMJG61yMQDmagyxqGZgBdGtZpAh
opdC0DUN6MCAgCLZfqQpbo9dgRbGgNGU4y3eXmQuS1Xa7X9bnW6mCitcbwGmCjk9
S49HWGkpjpk/Ixc3Ov0B6uB020do2LPgoyqEK52tfva7iCyvw95j6l1OKNbQ9BdG
QDb/cCwRQVgTsz//Y+D9En/LI+JaharIC0Ccbp8Zcdjka1LlgyJpAC6CgR7V/d8V
eefuJEQaweZX8FnuhgR5agKgH2/t8ba82EgFsL1jR4aM6HAwAAXg9XprfoY8h2MT
ipW2JCuk6hpLpZsqHEYkgF0nR+sAYoaJxsVgaGO5e7R5D1CrSJj6ICrny/pccyDa
8YCt+uxWYj7xHYVBy26gP/NrgTe14fjS5lp6K1SLtd2CIVtZ/ThGC45Sh9j3YAa0
8ALp/+l5Z4CM/ZDStr70fdJtGHA3svCVqY0Vbe6tZObsy+NCbkRpv5964B/fbaWD
smnaZRY8W4tCd2zdGTn7x3PiJU6gjJgp21BWYqsc3Xma6T5fr6+DppUTki88C+kb
8EdxIqASi8x0ECLFiUHGIEKfsGuP5GpkAGDCjtFwAY3rMq+BnJIJWL9FVcAy7RDV
RproO4OaYurjs/SNS0YE5xoWwUE9yFH6F2bxwm+3a96yqAYa5uZCWEkzlpp6RKVF
EnIYqp4uZ8/hvXT6k92KLyVZ2LDRSy4BFdYnjkyP5GUR2egE51DLFatMTL1iZ5IP
IjVNi9mjvFJdyCFy/JxNhJLMOPjr3KETXnHaQAp/Gf02PRduBNSStR4LVHsL6NoI
jXY5Ea1qDpDgvZ98kLtSCMOznKAGXO7W1gK21/hszXIE26+kKVZPoXZU//WHVtgE
RbTEBUDhDsTjJkFMIEG7FLOgZ8HdQkOnMJvounfgB3q2KPWW5r3gO5MK0lDTmMRG
9GS54hA7KrzQntoZxNP4BQtfohzGsApaH+nNrPQvBjYQn+PBDog9HeRH6zFc/01R
QtOcW0hgBR+G98J/+2PWA0nr0ecfFmN8TZb/X7GlC+VKb+YmpPRcGZFehyExVZpM
HUsIQTFrxrb5eZbIoI96J5xjbrClFioa+BdLXPg8PRKHnSCS7PTlyE6T+OjDGzbo
DWroTqbT83vGXSrOZBNTylQv4brqrGCVIeiME6GOOWMSHfeZ/sRtE3G2lVx8t7At
vXgeZzEFzHUoZMrxuzaC0jFPJWirHuGc7NmK1BuaSdsmhJKubuVaOl7EiYE8zTUa
UAKu/8XbpHalFIpVGQec7Vfd2agANhNV2K4K1HEdX5GfGTL1XPBH7d3TdrhKfGoG
fI6PolyYUwQuq5yrRhOnDVU0S/QBC0VS0s6kGFgORWYZYkK9b327Irl98S25IABM
0i61dEqPWryxIcVVoUkLmGVp9Mk8mQGAzVNMeBxKMhoI/Qcg7bHW1PNc3cAZdIo1
UT+Gea8H0bp9BFL3xsHaftoBXEsGKF+qy63aF3MiEH+l6sWuoi3s4w0x1NY6Ozj3
Afcy0IfmT5VAt/somcIpHu72MR5AbaNtYUriXj1HvXRCeZGrRzytwgXsQuqYPGew
O9d6jeroQNSbwMV2QAfkoQVjTwqmu6sKVWjHlDJwVw1KhoQ6xw4utAATYQXH9viC
ebDux9qZFitw2v8E4q7qLDcSk+/CZQZQEOTBsUbchOsKNGqTDus2wm2RwuxzyNW3
P8VbMcfC+SP2Ee0UznHheeQQNk03JRXzzRcb7EWJPM5qYtH7AxRKrJdsjn0Tf01n
D98/vLZWupIgmnG876ubjnIpkz/UMhwxg3yeV8GBl2hCkLtSpdnFdRAhsh3Cq8Zp
PJaucEY4+D0A3toWbIxu07fh9f/szq0PqZqYb6q661DS8B5MBgF43nZa9qipencF
7/0+gtiBFuQtHwC7qvBsKmnW52YfY855pCNaAUMgZd28ADouRw937gjQ2k91HQXG
P2PW6bJT+IGm1pRoYLIXTR1pVRIjA1HbibVWbBoGjDHDsZrRI+ApwQMBsvVVFzL2
jCCrEh/bymLV5b1iZ7pP4b7WsXRSznd1VzJe48s7tzrdZbJDzSMI0Zl+lNnkJg9j
ZsNniuYpPWmUgMn0oltOiQWlbWc5F25V78vcCHTMpyl8estUeR5ZjESX9mEcF7/v
huBEpvpaQqoUQrikc1we5ukefMhpkDGFCNYcaeaX5Os7GWKgUBIwQLgroPrIBsok
MBwoHe9KwyW07Mm6Q6uY0C4eV5w8eNegvkir3DhZaeuEz0Yvn3KMeaX8jtywJ3VN
BTOYADd0oDgJiVzf82FRdF5WAA/Lts87PkNqNAleGNh7d7XTV9DkZygKcf/uM2xd
VsqSO7eYwlkYHjGra5p15QQPUGCh0Mr8ri0GDlWhzYuvml/M7dELmlMTEY32xK0x
7VK2OclCpA+7pwFfU3gN5JLxgoBEoJajSYVv4SmiEPq5ERY6AGM2p3a660XPKgGD
bXPKGqUKCFeAuWEeIWCtOA5dRY4vDZ7zOucsH99LSHrrFOnY+FgJ2BQQRcrGWqxK
`protect END_PROTECTED
