`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTf4B5RKRyC1rKQAx+fFl1F0W0i5018mRQdUBYrdH2HWRovqV2VCL6F1xeBR8yRI
XKWYTlnJ8Sq0mYC/2TopFsbJS/Mbw2uJpJ6LBblghe/KMSe28RuvKHlAipgGWHrB
g+b6jcC9OuF3G91dL3w5dboR6zpKzG7RuovX18+FBhQk8dAplHX4s8z15rViBSDI
VVbSiQ+G7ZhVwmTYHPqBGlCK+P9d/uOtAkYyvTk1slKGf1Pkr8tf9ssVU9LZ2PcQ
65hwJOaoBYRx7YqZ6YUMr9ymJPu12zozW38W9ZIRcsFZAs1d43WXWU1yNTjsO21Y
/GRBKta4X5TWejUG7t87Tpl3gJZI95xdJQyQQ0rveVsHepvZ+ugxPbd2X4RocwEt
lVdgK6OJsN8jhNqFEOuFIHTvbHxRsEUkjsN95BJl1V8ff7YweHwvjkYyn5OrSk7P
nPv2zNf2CRXtbT4QBfBXpdMOmczQC4qsGLUSqvJiBdZR4YwSyIH2TtTv8OI0eGF5
y35P3NFqB9dKLG2+LEuM4mpCvuUF4GkBlcdswwYgOWqHYM4Vvn39K6yq218VS5qG
Ze/gTpZBIFJumlBRQF+Hg5TOEtcmyJDaZ34kdGbtSbmki6oFv2SlPdXYkIO+EySM
gyO5nKamj6n8Jfvsr/7bGUE4r4TMYnPSi2byAvYNSQiN0KKHGqMVWsyEuF4/xMo8
v9Ohy5Becejy4iYVd83tfBNnZC1Z6ubGj6m5Vt+giyF5SiH8Y8wwyjHYwfmJKQVg
hK/OQRRu2sE8Zo2qialuybB40hHOjSwh20FcEzLKzYob+5tYanl/PBo66mTt1MMT
ABPcXnCljrLxqpYNhPp+PkAzt2ZvC4vFGGlNOVbWf6ZtxmWL/WygONjAD+GzIaFf
ZY64e+55YAq9IeZXyYAlHfsFSsy80SPn+kmA18kDCkuQt7xL86NH/pJPH3x8MGik
K7Hxy4a56am0U6s5c/bx6cJEcPnnvylot9CL/ijmV3Le5J9RlaLDIgl3wzA7BWY2
RAYcPdo7icm1U/z5zE263cre2ArAviG+P3XHD1B/tQ1L89w983LMinpmKidT5P9W
5sThawN+iwshgdT6eBeRWOQwpLACIm3YuJgXuudsGwnPIK381IK28yzrQQVYQ80E
e0PAnUMdO+kWgR+YN/jn+c6u8McS4QVrMVYhcFIu9UifKjIHWrVCbRu9UZLphpBu
0gmZHe5QUoS+DcVWbIzILPJyAy+qiDD6DpNT8C2kLQqIW37hK07rfJ29QR6P/EsA
Sqy59bCo4uyV6z1Ad8dtGn5G5+Kzrj5TjjqfUH1nChNh62+J/PoCpZbk6hQVT7jI
nKz/HMCWDme8aa5+Jexera7Kela818KV0/K58d7I0Jfa81ROp2VwJxDU2pOgpUkv
WUJQ0Ww2KTNOxrM0HVtEALzgu96y8LRD0eSBcKvvHnewgme3lXtY0olKRKb7+SgM
shvRjEQX54KHdVL8tiP73uIlCzCgLGAgnGyRllVBFX4xgpLijEo1vEMLZWNmGW4w
/2K82UnpnSgLKCu29+lXkmSpsARwkr/vJrKOBv5rR55snZTun/fCGNErIOn2Z4Xo
ZbgE7Sl1Vy/gqwUaEZONWMzH8c2gXSMzOUCvUMEI8r3aIRaR51J21zR7+SZK5Nhb
Rge3OrC7B9/njHor7rbVHyJ9fOVhwh17/VcfgbFYcaSSicTiIi7fDsop/OEyLbib
o8XyXgeq2RFyI5W6fWRWhMj1gfa1nsM3RZ6ED13G5J9Y4Kl5pJ7BTpAK1+FuzXZw
4B0OcMftDHGJ740YRcCmS0m941VM9fl/lxqalqm1zmzR3trBw/1RFxzSdrcczXuK
Iu0X1zl81w+bBjUiWWmQYt8K3hbXqTc66Hh7bVctPzsUjGbYPn5OsI+cW/qa5Q+e
50Ux+hFSzYFeoV7/uBMBROmDkQ7Mx9DOV6HH34uBsw+5ZY1tTUWi6HyJdMSPF0C0
YveZYsMupN7trD7pS2rOmvtgb4vU1d7Htl88PmiqH9V821cnCCByU0znsChpW0bB
e0/5ajlqRVTHvv3uxGWn9FF2wejjtMlp2rJ9ttXKMm2lMKsN+3TMjvfb88iyvEyh
vnbJGe5TvYq6+GYLW/kJusZOxCYDasWqZ/0irPdUWWVufJuLZuxMQcO7DKK0j47E
TiLA5I9z690HRIepXS/PRVjgJU/d78lgykp0L6gTDFLWMFDEEO8KkY1CYBz/ZPvF
gYt1RHen4TectcshzNLMLJApFhVOEZbRXAFuFb16EJXLAieCoXCpabZS6xbaunQ3
42Czhg3TgZcmsw1OghxWUeHusUfH9dsEUCOi9lCfu5FsyFIX1jMkOiCZPw6xawtK
A5y00HUxp8aU5GAFxfm0fcZPbJsD0vGt49KXqfu7zC34u0aNFRCTmqKr3KwLE8AC
/E5TQquJ1dKVoWr3XtVH1ZC3L+x8Kc+6WdINlNRIh3InfENn8y7LOeHLfyiV8gXo
iD63PKRxuEENGN7JpvGSfg==
`protect END_PROTECTED
