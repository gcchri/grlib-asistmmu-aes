`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6ywr/eN1OAeoDYxu1rxvBUqrmiCMW26i7HsL5PSxiX8a64E72R7BB04Zabu1LNm
sTzb67EswUuPveVuKy8XPs7lzZqO0RY6LLQNPtd8Ei4H/Lw1B5TrZlN34FjESdKA
TTQcSz3ov8ahTLL0YxGyhNPb5gPyIxVlCLEYN8yv4Bu5mz/+e+TVYQTwatk4GGdX
LOVhRECi7JJsnu3Gvp5xIvsHRYq/uNZskhx80Sr9D6zobCGXv/aXloR5IUDFPe9C
DXVs3r0tIdtLWCH4nvWZdUZUTtJcUonZRNLY/NtEWGMcx1blzS6xPbseSP6nUC7H
RoGEV0FaYO6lu6XWdhl4zuk9ChImVBY6bL53nl6EjENVVbNnkNU4gqPsfChGfeH8
vlIQo0VeJL0L7QuY5hz0DKyD4QqjjhBFS8Ztvn2bgxMy0151gw7l6mn/UKjcTqjn
U/tD0LOpjfDNyHPnmmc1kRqwvVE2d7bXHw8z5sb5A1PUoKghB+ffs1vANoCr0C/G
IQjtMc6VGLKrUFjsL5y65uYEDcM39ljIqGmJna9qC1KQuSU+f/OYqfKJQ+ztLDS4
ZbcbgwJsXLnsoURcQSTXKxTN3xy9Lbfb4jqMxU85fCNfVWdMl0KAuZl3V1f6Xk4C
ot0sWfWDRGg1Rw4zHg0TWYVduNygRlrjq1qUC/UNfvB0RaPgShqCzL5BRBYOy9uE
FK/dvwfTy0QbItdZnyaJF0PFz7abXrfsKoU4ctADi9HUd0ZD+XOM9j5dNxD5+jkF
gHSmPBF5NPIIv+oosp1lCGMIAOf1kcvw+a5/y0HDav9ygxAulONEcbK0HCy/HFZv
Wf2cg3amjXBQo1lwG7Zjjky3myrNoeWJ7G2Hwvq5FmBIsHMF0YhSdsmxq+A3/RZG
wkCZTMhpHINAVah3/WfbUiOAHLvPdy8K88XZyzGIaapr9fVreFj1drbHreP3CTL5
0uNAxCopl0IcWzGv9RWHdTeSPoO920lnJEXIyv6nfk5hreQ7MNb4PSu7WBJylvoK
qaD+SyA0kDbQ0PpCi5a2D+wDodbjsnRwbxV2auiCrehJrgb6lwGzueSftwjLhRnw
wdCWOJRWELGRwfu3n/Q0Je9AODJBP18Xon2p3BXA72+mpDitSDC+9rSl739bldxV
k615aa2BAuLH6Bq+sPp8uQZhjGaVg1K5RYdhGdBCHqwtjHXzWSQWfYOMqzmt4hjZ
MA2B8JDrkIlfMgA1+HAupCjs8McnYFwRtGSFn0c8yV1tdx7Qb7SO8z0EPTgb9sSn
mkMbbiCZQU7dt/d3sn7FyEKJhfOcoGmH8fk4SrVs61uhDBMnnrlLNAQtAKiYM4GB
fr9RnLFczTuC035dyLTUoN6lpSj2qlVmUMKb/poz8iByV/36ljMgvYMIvbIoChSM
SvycvoRv/hHc6noMDNmd1f3ANHETyHuB+Y+13igKUUUmmCIk1u/qya/H2Feh97uY
VOk/gVsyQhr1aYOK1QZNiF7JGurVuz5cZPGzncPnF7xWH1hPCbH9iClcmBfOlOp8
sK3PXllrWr92QE9yx6v8UKPig6bzyj15awDpdPv0N61kKjkfLJnJ2FOIFRcPqPwb
yMg/0tZmWWOPZ58KOh7cfe6IsPo+EW33rW1rP9B6quTuvXTN6DzVByfZ8o2T9JxC
aN1hMkbc9IGeaEtXlcl94JFu8TNtHkHD+AvN1VT79fwBs3ze0MY9qQg5E8iL8GN8
wF2m6fVcniHea5o96kCTt3GHRtoAh4oAn0heqA8fgOHaCLlTYsffulZnY0fi+2cH
8UWFSlpw4fsRNXUgZ7XeoRykW7dk3jTmeTd8Ild+2lEUFb/iMYB/EqYqrZ/GvYgw
g9Gb7/nnIj/yDuYOv5qUPrTGbZcvhPM61F9ZwX6FN+NPLHMoQ7l3y5jg0WWJ4Rhe
P04xy/iVz0iyymBnu6a5YFWr9YQMFHGa4Fqyy0iXebWBGBgi3Q4HDAEuoP0b0u5X
Reht2G3jV/KC7o0U+rwZ/HhDPAnBfZ7EtO/cS7RzxYUQVtJSSwAQN9mvlnJNExZ1
fAEZBx03I4iYjEuTiePGVUaO6FI5n+Zwbp60SZsZPdnuctg8NG/ZFCC3w6dsS8cw
o95TlPElJE+U0dp2fbhJyXhQ3UPhhVLnK2oeVUZeQyy+PYOZ/Z5LsBWexluut1mV
9ScZcKfU7tfRxHFBaZ5LnK6SfE9itmBPIdgz0IpxFpw5S0QSXGTFjrXdddbwaOuD
o+uUBTbm9wzw1mNp2vRtrN5uqiDqSs6X5sQp9WSB0W/C6d3OOc6o7yy2Ne/Pjp5H
Rtnt4V95uUFMbwjFo/St8S9NR1s9z4ZVL6dMOOAVJaMb/S22GDSCT2R/9Pm64ILO
QxsXE5TPhXhsCXDkZz7PqE2s/f5jUn2qdJwjFj2IoYuHeHicYGBDm11RS8fFp5x9
tvz975CRi1Z2FGmWB4EJ9U39wK6N2dNkA5u+El/xVFPI6u9jRYwxL0b6VzXY5uD+
RIQaiWZOHMeXpSmBENDDCb81wU2zSGTErOpbeH51iVBDqpOyxiBq6UN3NaRdr0Q7
uZ3YSn8erqLTI5M21F6DC6ra3Q9xulAiPgArzkkETAVY18at6bZpE8sQynYt7s5p
A61/0BDSuyGSxGt2FURL3v/Cm3MEcH/n171Oup4I75cNe1pqfuJdzpwiBINa7IGn
nj98lupdnduUMkNCR1xAzpLID+JvucE62uzTdELuKEC06zgeXck0z7JsaFFS9gZy
vxbRFPOvnt/hmudBpCqatVKEucoNh9/1GAnYacmkNlcl6fEs6EVLoqZOkBszXw2T
ziGFRny3uLVT4aHNd0igAaoQ0XzSSO+zlYIgYYb38CTyXuQsdGO4km39sF5kUz/g
5rsfNczoxuFk2+J3A2sx3zBl5v0FY2FColBFTzU/Ok98KqVfOAJ3ffj0WDXr8+PI
UVq7lAjITE8SeqT5fnUH895S5eJ4EcNiwfwmpd928DKlxUob2SGztPHk21nCLv86
SmoY2C88h73++s+kiimf3M4dy988YsRdyQwI2t5qP+guiJQ8c6JTeX+t+xoGnLdF
Rk5Q2hDpCe35Z5YPO7Q3NOaiyQZKpxPxsVw7ltF+yztL1mXHI+aX2X5uCsVlb7na
9uDluaaiwT3SD5eq1zf4IRpo4FN0VMc0c8DAhohHXvkGOTklzNnEGgcVg35uw4OX
h427gP1S3U1JzIEYgyebtX/2DvK8VxRsofiwvpE8cxVqxXVbIdtL+R3+yM0L8AH+
/VXmtG1im0nVGFDoiEdkfApWGYmTK7p6oSwTwKgtfHwt0dswRb54dVl4r4r5VOmK
Qvm8M20q3lyFhnwe6dFoDnKrMmtTJaycsfsVGq3a7+i/+zqGdY+gpdk9aZJpucvM
10gEMWH7gJIKpiOJwjx36k8Cx0SXj6p8GEThHgSBOmaYn4ge4o70Cca1vR3wviOH
+h9gWB0n8zzvR94lTU3RAn8EnQmm98RzBFwldbH0RZs3LjNn2go4+G7qAn1Jc6rf
c03uPAOeXuNHExJAmbmMOYep1SSzYXuahORGrgROr9VAt8qtE3kzO6ev+pcfXh/a
Q2TXsc56n9RGQDtSnpT/pURyKIzop6wc2k9of0BPM5li9rB0qF4NbnDXWWCCojdH
`protect END_PROTECTED
