`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3LoUEkgejcw3pRRQSRqFCrnZ6fvZknZzc2A+bJHsVIOpJtbhA5TlcR04YsfItDx4
8bo97rpyAZKUrD/6x3VA7NyW9/I2Szzc6tnrMUIFKK7RoM3UE1EFw7cWIq8e7dQA
KKhJn83a6gpJzgT49Hszn+v3ecLpxij9rZlLtq73aA2JFIQLs9099Xs9gBwvx04m
BxGEAQ3cu7HYEwapMHN+5tyIRUt4tSdzSnVUg5a9mqNxOOVP4we5EpR3EVJD03wp
BTKPVySn3JnCQ0YLmXckHgFdzhzrYfmmfz+6kReFGifY/ROMaD0HpQGNQm0fLB4k
+I4oDFovWqArGFh275/M39URvMTQKEkIysyTYBkA6hOV+lnypRKWsVHH/viyC2tQ
6bzeFy9VyGc7NbzeL5jSxhXDbk97dhH536zugDFbLFw=
`protect END_PROTECTED
