`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HNBP+2F0+F8leZqKBdlXpubKdIBpRNDu9H/s5H1rfIwTduHfsyH9SSgwHb539gd
joxgzEkHsFwNiVyOa5isaAAwu0m7eJBWC3XfLP0NLm8WK11V/hGtn9BZt6ZOs+8a
4lktTqw59feGHsOghwTU22FYG77rM3bi45nmgBdXHCFKD8pJoC7s4Rob6AwmAmsx
q/AJ/uwiUoTJCG69sXJ083QceppeEhgWmCb+MAxz1DZuYm+xDpeIHxwXruJfrEXm
r1O+k6qMaYmx+hdtMU39jxftSbVm0omQpONZLB+PESE+yZ+ecbQIDq4XaEqM57TY
uyCUEAVGscsA4rT5fViqTw==
`protect END_PROTECTED
