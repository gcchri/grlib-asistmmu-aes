`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f0s7eQQ2RC63xjm8dLw48tTo6NJm56y5Obw6v0/VCOFJ5Q+g0Krnyw5jiC9COd09
+8Lu9FO6YRrQNY73tvBmBzDj5bSus0883Z65VgQshM/QlOfeDI1clxmeXW7q79Xv
d6nghLBCF9Q6b2OsEFz451jVdKRyGT6VUuO1FiejoTgXkZOsnL8tC36JkeNr6TX6
cI8BQ1Q6QP0DRoExG2JTTCo9GaAL67WtPOLD4ec8iJxhLGrA0AVFDpQYWPgH5agG
EZWEgOc9oTS4L30FX8pFxCr/DooS/B3OCOpN6HTHQ6tOoNa59t57NY7lRXIaG02O
/tOe9NKJwmd0Za4tRuHa6KAAuK+boxW1iyuV1zZFDKr/gPRGv6Pg5xyr2C0Hskkd
BQbAmNJkaprxZUh24vo1mBRd81voHCS1cMMLGRjikNFYVCyLw+aDY04gUfzIxBuX
8uPWQDNnqQX321NNtiK5qPP+fPKZDSsuvtVd1nhWR+j5SIWbXAwZcrqcfpaM1s9v
eLgs7oL/GEQjgh0CunH8l/+eAqY7LLkaJmCRszI6qE4zXqT9o+TgsF/km+9YIFx2
RPfkFYVq0pNnLcTgbxjaocPe5Zj7hPXQzd3hfA2t1WiGuz/GukcCz4TfWpQc+MZs
8duwRQxPDMM8EMArtLLD84BknFhGBEAmipGLeRT/9e5hYczfergeP0b6sdVKz0W7
zpPeMFENb/zpKXjy5gpROWnjYGbdGbMszaKQzC9lYjGt0n0BYS3J76SNdNhxoxj+
0sNkl8vd1P/Cqc6bz6UGfw==
`protect END_PROTECTED
