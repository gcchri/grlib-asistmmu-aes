`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nj/lT3ZPLhsmlM0AK9oHQ7lrNCMBdOPQgK12Pu/L0ztT0ACMFkpOrE95QWNRlfQx
VTRZfSd9gZxPbNSw4D/NiVBRzQNwXMjkl0hORVQXoXJtyb06v7foPVlaTPS4mKtP
9LmEFg8iKR/+x9lj64yOkYp8FiXQVzzIGDkQ1jf4s4uT+D276yX79wZCWPz/WMNn
be8iL/uktNwIvh0oxk/nu+ywezIl6dJ7OkLsB2VIFgP8n5wI3k5iS5zZmlrvmju4
qIUTRGHc2sClZdrI390kGM5/OmnD0LuR4aAGO2AiC8qGMJkjrr5Rh3EqqODQzCbD
qg9Kln7ccrcIP0OirReKQw0LGy+81F69Y2S51+vO6Pvtg0E9zJ5uQ5lx1k+BcUQY
uksT5TXjdBqedveUvCiLA7/VpUtmEgvIT/N9gBxzsTGn+niD9/gnyA9WBTeIqSx6
`protect END_PROTECTED
