`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bv0T5HgsX6W76PAWM7h5rG7t1eXPxvcLVT8AJw7UaeXkmdgJx/3zQpALJKsCSFYM
oKHV0sbWRTkZSnYFHGinNRnnSM+JBq8eIDgceTcUkOym9RnLQcGsNMCihnubJ9TE
u3rmxLVlfo+rG5yukalnR1Hloa5Ea6SfB4wsundy9D2e8RwejJHr27LqSuSFIxTv
rqY97Zqd9fGl251XrmOMOAoSwhMpvvm//qDXncJphmx6Bp9iqteHCgComsjOlF3H
ncQA36ih+rqcxki5A3ytsrKZPEeDaLqyjU1ysI789dK9KnvW1619jnMZZx1RdFGX
LJnWsbCRw8c6yCmiMeSYuVeq9QNeBuDnoPQLoIJrF0g6Cgzm3ZDxJ0+27nP/QlDw
DU0O4EoVw3VBFBii2NsmTbpGjflaHezw5/xZqZA+N+DXQeuxfcSXbFSiVS+YSbcN
P1EzFX9thPiP2001zzgGxGjqJX8p12vYsyXvwgs2EWXEKxYBbHmdOW5R4hjms+PA
GWISri0IRtrro9e47GAnqGjxky9S0mg0ZhLx3pzYuYhIeqMAyuhiHiKGTrAwCfe6
4zUIo9gfBE+L2M9SRauL4fMtN3olTOlqsO9Jfp0yBNu9WYA39ow3mTZKK+zPN00X
vYznQjsC84GXuxxQDRrXLw==
`protect END_PROTECTED
