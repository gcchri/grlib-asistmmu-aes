`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f3AGGcFTMzjrvLhfZ9xbOh5+JDMjq0wKDcZ1D3edXlkj9u4IHFObpQy8DqLS9sF3
OQZ9msD1C+mGOs/IpbfqyZnpr01kOJI6UmM2j08R//WnTJh9+HEbGEcBrc6pVAzj
yrONMLZpkgdRV9eY6LfGWU8uUeQ9V0ZKW0X72Fs8bwFbesx4bdkELvkOt+rAb/Un
vSqxlX0wRowXyUi63gCiwp7JXr8aAC4gEkCYGiolk6JqU5QZzXJ9dLL7sndNeRET
urvwDvKEU0ixGi91C2qU177cA1OoTYfT1mBDrEZKpeHf5Byrfq7NSYjAMPNSG1ou
wEpBMhA71UqtWfd7cpv1GSRcfHucm3NES2seXNfRv0yRXJAzGPI6q7KstXLSntg8
oRkufftcklDKLbWdou3JQeWO3O/1EX4euB3jIF1YTI1X9XoWjoqxdnmOhPZczRGz
yYGP8Kf3p6OgcJX23GP7E7+GgKaWlcDigxoF/m511D/3nvpVNPsZ4yLtDGAsaV/T
0Euc+GwvqUns7rUcfz+2y6oPySy//X9jEvTG5pVCmzvc6y9vK6AFQATClcFjEM5i
WbIQM2hxR5V7vzXjvztpceXewaRg7IxcAfxsK/lsNBst1LS0qv+3lsUMHqusHN7I
3P9IUCZz4X0+l1HoWMh2GnV/LNCVIJI2CsBrUYNq/S19fhm70oU7CrMGw66dMCyq
1oFnUP5KTm/NauchdDLAvmVEzQEqt5rv9ccW9+tcHTf88V8h7Msy3cuNIJRkp5K8
/+kF2DEBnvcOWs4bwRzyRsNnxNbMM8sUY04t3btn/Jt5l0ZNNJAA1cq2FMqkEMRR
0gGu6q9mAcS+c3l8h07dAaHfsQEkCR2XZLmqABSI1OAqi55bEUkLfxGr4Sl3uYd8
LUozGNCNFYtDt9SCiIQYujwzPTDKj7JoQ7rtcJBS7YUI1C3xX0LIdc+9RMXNinjr
r3UMYiQQDtdgYKKmNwh7sA==
`protect END_PROTECTED
