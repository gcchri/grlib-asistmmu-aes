`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6DXheyzTLfHZ9N0emfGJOmpTl/2l+/uc3UkmcUbw0gVddtkL2zNUz3ZkSt5Z8zjQ
H2C7JTPIUBvlTdL+KuHNIHXB+g1rFAayE9x3zDnEsFZOW/Xuimd7EvwMiLB7mKKv
+xzxUyM7ywZdDnOgtVAzmvUSVZPDtKjanW0bjWRwYQcdSwuUx4FcS5CUAqZI8jnS
duidGyblTnozt34cBWcd3YmFV8mw/V4qseOmUL8NWbtVVxsh/iHvOdC+WFte1y91
ZSy1OgnQwF209/YI8q5JUm1bfu0x/n71KZbaMmzG5elZPdHZzhvS8Ct1kQ9g/IRO
xqHfWDaf9OLjkCoTh3eA8xBCSXImgzJv6zhz9/ToAk4pEsGUm8BTdJauS6XD3LYr
RH061FCrvqeyiNIRNbW36uhcUA765oD9en70DXPydFJ5OOj4OdlGydNma89N2Zsq
jHMyOK/gpHMau5z3GR9yGNYFimf+wHWsUQCCYUE2hUvvVPTD44lEHbemglkRCwts
7y9HCtS5V6VNa6xjN4Z5bCwaHI7kEuq9/+mAbgcCobNRKp6mV8oWh0rR+3ssYGrj
6Je1BXuDEWYkoyU9VxGQoMnFgTy44RxhzcfSL+efqygGm/Se7MrZk88BkKAS/7mG
ZtN2zUj5QyED/bVDMGsu3SH5l07QI9/APTK/ET9Uit7l0BAdChi8ooriNFAbbc2D
PraAl0rSG0SJe/6/AiO2Mz+9hYOAfF9rvDSzst0ddYH98on4+lc5z/WULTwAcIVH
cv6mmihoICe1UslIdmUaf0++tz1xTX7Qkxok8hWFznOR+26Eg2vW1+UHEp5L74nT
O5bQLt0IlTrLxKzj6NNHIEcUD7ZsGe++SqiHrud550Knay8z2Yd0J0XgIo7f/txr
7b1Oeei2C4aZ54UeT6Ys8xE82VUOWcdu1cwiRUFlivpdCkOM9el354Au1zD97ozF
5G2EQ2syUIfvu1uziipcgS2pOiJg90LLRXKTzhFtS2uddZxtnsKVLR0C+rMRyQo7
VkAJtZwZaPO/0+XRzpZ2XeJzCPv3w1bEPop8IlMBY1sMkZvDHCgRsPqusc7U2OD9
LtDBWnihfRpKMo7Mp6o+RfubUaSDQ2QlSg4lbst7HhacH5bu9+F44j63Se1CgC9k
ZvOR6NIhDyE3RYQIExcOaphAPPc1xRN+pW+kpJQqBkTdEf6QEZj+GjR6+WExgGW4
S4NRVmGsGbYwUqrwpjh/TA==
`protect END_PROTECTED
