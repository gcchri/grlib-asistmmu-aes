`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BzaDqFgmx+LFdct1xH/viqOmg9XTXYijHJ3YUBwroRMypyFN/5QyDwXBfUcKsGm9
+9nUGtMQLu7tYk24U9sed1wWWR5RMP4byXDka3EMMdSLma0Ku7njMn0QW0wsLBxt
R4RB+1TUj4krJQ1bHd9vTig14hRuVhZ6+i7oz/K9WutW899LoORfCZ/9THU3GHxs
iUwZpEzxsTS6hoEbRNK6XFseWmCYzamDv9ztVuTrRAAfsFtYpYAQTiw2u1moygaz
VQ3uFDs+EsZNpSG8/Yjm8D9dSzD+8Dl7IyvxNtFz3gwxQ3ByzJuZvT6dVwOR95G6
6cYf5AFCWI4ZPG79umZNyX3SKAqmpKhhoBIUYwPnENVpz+TX616E6PC2K2EIfJ7g
eqZo3a2Sin707NrkSzsKXR4dywO6AJ3oN8ruocmMMFpiGsJb3XgmKwgc4wgS+NLI
UNQCNztLs5T2N3VqEr2lBL3r8HpLbPk6YgW10icWFPE8vI5Ty0FN8cjaus0bwpm/
x00YdoIGkzuOisECeeRyA9bphuvCS+7MN70ZmfkrQezeohvdXuvdzJ7LA+V5Nlfq
MUq9UsY/ueiDO6qz4p5babj7rcxQUI5nUASxk732p1E+INbDcSA2nlfXoUozaJMb
weOVtCjXRHHPLmIc5kRPeN18Euq3UARKxswbLeMfW5BcBMGHfQ8Lx4ixXVs6s6Sx
hely9nVb/l2W2SNglCtGVouS58cx2WL19PYorjkKpBVOuvugJ6NgG/ZM+DhQUjAL
HlXFMUIbNUMUsEu+wub2Z35+UKLE0aGQ4g8z0mM1Gj2uhRLMWatpf/ZvuzS4Ph24
oMNNOyikBoE++x8+D/Vwgp7zN05ISa0pzjhjm0u7SUEk4cn4XeRRLSLXwGZLsnEr
cz4LAoMpFwvCzrt2RxDiEy0az2khz+tHmqrOEirbyHU9qMnQKFBYdgswEhMNPCAi
o3uD/Mnd6n4SPkbSJB+zAgVNFV5hO7BXhpvEEVrP8F0=
`protect END_PROTECTED
