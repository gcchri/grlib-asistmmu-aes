`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FkXOB57dQR/5ecEVBpTdY/YQi2CaypAccXeatd35o3kURvmVw5SAAStpv1onYSh/
5s+NioWjKPtwph3gj2yw7D7M5lQhoc4AiqnCjcsCvsJd+7V2hBuXcAsYfiT5GbX2
E34zNJVSPzl6bOkwvCEGp91sCp0dR5L1cPwuzKoIgkF1v7eAygvXi24pQRGw/hoo
9hvhpCon/sS+YqjM7f2XQzBfDWQiixm7YiBqcsWKetpFfRCU7mu/u4ig477KRdDz
QXsjfFL4USoXlu+IMmXULSuCtqHFwp1woy01pNgMQRGbJXWPBWuIgh+x7q7EcU9i
ZWhL4DgrbLIdxP2TU9+L1JkrNWX+c71ECSyF1pPIcN+bb4O2jUvKdehts/lcmejg
RVdeuSnu0AS28HPvaBvvvXp/A30ulY515Sx9HcW1Cfe80p9WFP3D2HKVLYfb74VY
+oxtGylhl5UoCqh+MQMoPGCxzpuseMuzKOIB6qs6yOGsbMY54i9fvXoea00hGlMN
YIGZnXUqsQ7NrFBbaFVCGo4M+YwnS3YQG5hBfwCAZnd0GRrLjNT0fa4yCECkYYrC
t3jU18kvtr3Ctw8BfVqgMVx6agrYsDyMiYEO5U7zd5/KO1Mj6Dsh5xb4Tzyq4JKv
4XhslPqEFgITAYAJ4u4ocA==
`protect END_PROTECTED
