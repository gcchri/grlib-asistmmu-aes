`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVSkqtLViPZ1RicugVY0dF5eUYoHpgrid/D+rkLtnwykLoQwq51XVrocwQBmVwVZ
KexhBDQpTUW2OmgVyD15qDM8g0+S2AR8EvrJzxJjQogylAvMMxcXi7T8JXSMD4qd
kyjalWjKp9RrFQ5VNCYrXzQ1Mv+7cbm65onfTCqZAwGm32TR637CsZEAavxOhYN8
rs3B+5PSCaPVgCPNqMetojxub0bMB3RqBIbt94HJxmLVNWpdw+TzICkO+GtZ0dCd
vYLrWL1ybWph1LhRGyC5GgK0cCiQQfx3GHARtRTQ7CzCNXewHEXbn+YEev0+oPib
H1birxMyub3CMA4RcD2T45VJ0FTrCug1torbAhxnz0un74ENOCIQlrU3W7f1qO4C
Ta+pQswEazP6+ZEwX51f1fhqP31hCaVFmUFiKliE4pZYIceCp3TlUFvEEcuLK2Eu
3djLv/pt2zwFyIpwpEjaWKIZNKQe2ydm5QNPFssjmYrvIZtXwhmoZLiLe2wNei8G
Ie/XjbQ+/PAOLTF7rWzg03RIlef94HpgZ/flUvuoOttEKSOdY5VT3O1k9SfUePLn
XpyhI/UAFsxIWRTcrc06Cq6vkisD5r6WiixY4k9ArxuKNll0K5AqqZL+QgmHUlby
/CC2qjYEOvm6I+/5WtHHKaIoUyz1fCgPu7gjllXpkug3EqwwSS2h43o8nIadVfr9
jtDq8HTD9YIlajZi8+OsXW0baJAHRUU7Qaf/SWHewVRjFGWzCW4ozvichpngGSzV
sNU+FOrnt3zoLPon2OKI+zUAUcieJ4TWppNjbmHhIqhvOc4dag6Xuhg3ZI0cZ6Qb
BpLblUMhRHjanZikpnEkYSHWtGo+02vL+p4tePTwqF7l/DMq/Awo281tO27xJIK3
Cp2KjQJW2ILjiXBH0sDKSxwXY4zXsVADBB6+R26saTXWUiTJLcWwFVkFyaMi57vX
bnlHIUR8vc7qBTxSyZZjk9FdToOtBNMXa/haGLuBmXECDNgcOmJswnesCuFyXVdA
vv6YudDR2iqZZIipApeGUygD5CDKJFIEkx4OuZbjxjPczSBO0HlBt0Qa74XzfwZL
D2JGZhsLpBQBATsGvowhqLfcLJIFmWle7ajL92+iOS/M46yENlFviQ8EExOhukki
3+1cjcxB0m//CIEhzACxrmIwEUii33ZEPUu3ANzeqGX6fAAG2z5hZ40ezqKIGhuN
N64CbxY0zz4t3ZtTk0zYAzuueUgNXBTUFf27GUs6Ki/OJ3IMPY1VrNB+kfh2QeYe
a5mp8D2T5iaBuX6N7FF4C2MJmOcG09iSLM2r6Kf66dy0fI3/8B2m8CusKZRXfrTO
C2iVanJpTeqbK4MwFgELsqmmv4nBI92YTQGoRskg5GQVPKRHs0wl15onPcMZ6QU5
OrH3FtA41BEYaDbhOoakJTluZ3gRcrznTNDICs8dnN7yYnHjm57l9rUsyogOj1OA
ro2uMFEiz/uwne+0p1ycSEGfJIteIcnzOEUymiIiZbm82Z4GF32RRHrS8UCXZBq0
XEgVF8UatHkQhvD9uw0ckCH9hF7q2aVcbq4yKPQ6i7Mbwgj1sJYnl31yVI9D4NI+
WNMv3y65XDH6Be8ZvfLZR4SHfbjCAmo8F3hwDz9h70+7a82yCO7xDqFq4SKCdHrS
je3t6VvsQXqqjGbW8JIAYg0E/RZmlq8Jehw5ekoEPVxgBgL8/AnZNZBbzLPj9nYC
WsUENO/9qM8HAX6f32Kk7QI3yNu+v8ss62WNILDerm2x+3C8CIagQ70HdCqnRaBj
PGbAMIdQtWA19iqHsEmQ6D7FyhTGvL+3mVj10kvYmP4PAegdeMrYBnxHsLNK90nB
dI8nPR/0g+mZbD8rfj1eAGwK2dBgTrwkEjbhRICGNo3O15xhsmc4uy0Chc3BITHN
kKnJBXJFa+U7+R36uJY0Y1jATvDwEFpF8nqFyALgMILKJGq7xtqlOy36nmxY+swM
mOoscsdr4ty5TdGJfSaxlvbaSQK3dV+HuK24q3ljzxnvUoQl17qYW47Ws7zFHiUc
vT2pqZoCBbvVt2AWE+OGR5hV2iPjQaHBPsGwmwgc3SPsNCVz2eX/RZiFW6ix6sk4
hsMNyqmHLYtdHl2uJ+2C7APZMDFitDVVW5rNVC4o2bwpvwUlu1g8r7tgAaqdfjLY
DiRYpKf5ThOK3yy9vYbd6qgfLo//FS/vhlh8A9V1hEOgkhe+nTyuJrlon5zix8v8
dD+RyWgss7dq5/hz4E7lypXn2wG+lSgNb741WKHoTGVg505nO1IfzjzQa3Ey0+yn
k3qdFVDeKg0FUx/5Z/KGdTVqVRA4Q+oRP9ViszCd0y5bfgzQjoPMHe+fdNz8AErU
ePEpdPoJEu4NgeZvj4eW5MtxgsxLHUlRT6xj6cEdWSQx20JHz2J8yfk9RetoCrn/
bdH7br21dbDe56hbZVXoXMI15oKD85t7qtbHSNZr9RvsiybZgrY0cNBlAGY7J+8E
B2F7DhT/4OnPoCJipLW82+8tlTUALQFOQn845llrX2ju3OzMCqUIaaEBW3VLfBWb
WtXAgx6ObEq4srsq4HD0rzZCvWoM9NXGhOCW+xukjOgj5IjJ9tToJ5JlkozKCyWJ
TxCD4ssHmtvl/NL1la7/Wiz75algtyLdvaPoQdQPFzsPd9ZOf1nPSY6KMSS0oYBe
1jo1vJpmjEFAcGYUPCP76RsOihqYXs3z/xwVHKh7qlXMaA+LvUWp3IGeTk18vNS+
AENjAxvJAp2Ch/6uIz1Grq9ie8PCqqXqF13MePiFYMElJvvDO8JQv5Slkfl+LaaI
NecRYlc7s1MankMPZB6Q+RZCfrCkgFdGstuMZHFCa8Th3JSX3+lwwi9Hd77TpNpj
Rm9ftV3BipNshYqPyjVI4FffGVEG9nuVKm3mLbmEnRlXQEksf8a/QhwVbee61m8d
OJB6aIF4U1uamfyHf+f+/7wkALzqRxTrH6yuHjSszb68UwLplr+jFfJmSZaWEMn2
PQjppYftozhMJFYUWa0C904PUomXLAXJUiQFFOYKt/Q7Sp1cqBKn7spBw3l+X5lR
v2YlkVFGLzU86lf29yF6zyNZ2KYuiHxwF8VJm6SvBZY40jNtxjp8Z/9w20xMH3c5
54X4GXdyqeSVDE9WMGHRHnSbiU0zE+PjS+Nnb3l7Ti4Xa0+c18J757PUptx+80uR
K4xKbL/eckYzl/DJZJMXwOpAJlwGpMY5NmcVu/gEvXZp7b76/3ygmBhobff50Xqz
k54kdKgDSSkaUp79Knz8QNIn3efRIozGOkOezeHsohPWgu77Dx5ih707P62egioW
EHu69etolDsUskzsw+by2RqQzKvKJt+t745Q723Oaxf6ws5fkRb3kO/YfD1D5wYx
obydizQIQhU78DSfwK/ZIhylarxOePbetrIgW51SXE6ciH468s8od1iZvFv2cjX1
Dyvy/sEHjuWlLimOKG2gHgGFuTempZsv125yiKRgND+J6Ea1dE2J3x36wWvsP8ta
XKvNA0cge1MbDmuovzSfxJceIHUWkegmPrA6GRZFFgCCRH3QYfADc/ECzITtiBSn
fQj4wrBiq/VCltuOruABazJ9moRdLTFcywZc023FyXzER/xYLMF9tRR2oPk02smP
PlI+PUsaP+TVpj9KMbBYkynQf2S4O3iF1Hq/MHHaiS47XFN3DSHgpXX/Cq2Gnp6K
0KQQ/RiZIOwg4nrCJQzq1k9G4JegK47wG2aOX0cJWjpvCNFUbjC0v9NQdcQDZkFy
sR+GFUCRX3fRs56Kil1Ix1pwQHAHnP13HsFAlrgc8xvUwepufqFSVdO3E/P+iLao
3taEP3RRR4JjNJQ19/Cf70oiewukDPFGJVcScQOdztZxOQFAJoJhFKqKGCeLcWrJ
DigNRDiDbnV7ONhpHITbWgDHh0kIUvFggYGpaTW4phh6SO8qD7GS9V/+ojMUjtfW
9H430dySlzB3qFZXxqNDZk+fIZlfyCwz1eUQ7VFjl9OWi+oD443Fl3Fin0XcQNdU
bSwgrL9irtFPMI5NuNmg1pseAFjs9cdhM3FwcLg0n4ZYN+wdkBUrmqx3hXsZoDeo
Vt8xMj5wbzOB4eDJxgKNvjnDrcqEuCvlEjfsAl1E4GJwXsjC2cSUEAS9CwF22MBw
OqtovNQgjrqb+tBqLQOZRn2aHjTIKRi5BtH/xzbp3J16tc8J48qroUdPyC97Ivyo
zd97AEDw1NQU/Zd0EPbTliTAUDBB/l1epmGKg/tq3Jo4d2TF2B7oCePkf6u2yvIB
3GP97xqzh4GPTwgIADdOIQEE9N84Ct0kphr2f22IMcDOIWZM3s2ZEq4HTfnQf01s
UFRiKTo2vAlsCVUFZYWoCGN9WVRDLhSiuiNG1qvlxJXDHjogDFGdlJ5dIiepjwOl
y8lGqi3aomvd7pOKQA1aTlP0+TDxQ+dZcqJdQJ0vYicBl2ZJSFb8vLsQhiPoygGQ
KiL8S7woleSspISF/ObXOd3MsOPabI/XJ2nwcRs7oaQeCl2M3g4lKqwKwwkbP5u7
0uUzsT56Ih2g+Y+YH9z0jvJ72/KGyJhoQIj1b7xGZuDgoxunj8BVZGEaFgirsB9d
rSoaV5o2VMlavQbbXQuQZmvCwGZ3yQFryMPj4iXUD6irlJrxQAcUYbbDJRLIr0Jw
RX+6LvRj4jVXj33oPibmNm27CNRpAggBMQXvbJXbK2nvpn2x9xp5CRr+WLLzjraA
HIpDUB2tdcVSWSgXrZv4uMoGJsFjciI/k36FibEW+kCuheAaplDFcNe5Ma5jajp/
yNJgS8YrC2f+n3VUBQg1TWpGLQ244jgUiimCWamLXGbVJaHXhA/9HBo1rlA7C1/6
r26qAsbF6MJCgt+LSINQ2Yyz73y1sPtCj0tbn6Q6oFgNlM2Z+3B34u+GZ6A+i57H
yAEyC9NjGXyGpwfVVfowNheHkVp3Ugv1dBoRYdhlwgL4fWVBPXp9eX1LCeHaCdPs
f9aZFxXykGvKIs4sDiwb7CDsC5cZZcb0HBkLrYevp0U3AKIr8nVY/NFh6BSaxyt2
Qtm1XDv7RLZADoyqz2xRjWBhfM7j6i5zDsDzTnJjYmde/muXmijIbZQmNFJl0bt6
1DX8cX3MFsIT9SuyyFhNpABImaGREY6iByP42FlJcKVHlDz06c7RPiBn8rqjg7sZ
hc/7r+cRDTlugEKOzyoKlggInLkFG+AY9g1n4h953iYQ4sl9UpS805WNhlM/1Ib0
l0vgr29NeAG5jinz9jiY+1MpEA9yKDYpcJo9m9XH6DuvHB22K4xEmKMQ7gXlfWwJ
f21DMLijVC1hPubicb4e1hdBX3ALVBcBg86IZMq9EwoDCFgWsPPYPfQnYu3r7xr3
lxTJ+kphHTTmIMygWQt9Tyj6MQKNNfQ0FFe3s5TxtEo1C9WfRNkDX1PqF9lXm4Dy
rNkFTuMRKbM+jOyWGVyl6Nmm+nTnjUsmAjyQS1aIy3mt9+YfeAi4U8GqHlOxtdHH
igM7VOrAvsSocuCcxMQHf9cEvo/7dJ8KG76bI9/F3sU71kqH04ucebu0b27nLRfB
fC7YLRMTfBX30W3sOl4NwChu4ckMNSBc+wZk1toCWPyM/ZTdAzatZx36JFfHodPG
Vsz7PS2BwBxF0l0VAzP2XEsv55URyo6BFTaiDmf4oc5GtqrMfngsH5NLCTsjAE2V
9ZxiVbhhRNcybJ24e7eTCRrcOUQL44wpRJWWBQx7EbSqncsgEHQ1VNueeIOz5nSy
CxW5Pxz333H8Ps8l4Xe1+FFVQxO8PXW9F9bhdlnch/VJBwwrZqVMvNTlzr95OJHe
pL2m0KXoGmTO3w7wAW3G/2CdlIyF4jmf1RIO4vyln85bt8iuTc9uS6C/Fk/lJv+X
ZGAedFwOLc52IwXOVBhxT3aQVtchehPgpe5uq2f2cJrKA67kHctFDQcat2eNY7r+
+gFVTZ7HPIKQuueROJ7eQyug01ha2W0MAlsTF0RX3DLcoby/m2SjHO7rPfE+wRGD
OZIOwVinuTr5UkwqUykIHDyFjeDqcN7T9wsKmUI5982HE/OSI3b/2SwNmuZkMStt
5S+wIsn3m2LG2g/lEhl8OFI2qWho0UozK9hbro72EXTM+9vDK3o3hKDvI4kGzbn1
a1kHgQgml5alMw+H+bSitmYd8/yqL8jE0o1MbpxRpF4wgCcxuh2I3RI5Lt11p8nP
KFHDM+SvrcxRtai1H0686PgBoWfELE3wu6+XiQAFFurnDAmC2BXHwEjL0EfLLIkA
bPu64Af1mgPU2/NdFkkU7M+Vj63w4ejDXd7KUBTrq70VVsSMF1VV2uIrWLsm2NnK
GErkhECy3YlUOAF282lSP3AdSeOJybsbaT26C8QIBF6oI2napRIIUr4VwGm3441m
1eejyZig5IrfiFXq4Xu6M+73P5u5bPTwepL/wiaTt3/NLzHJ+3RPLs6s8ijjr6Md
ONOEohtcViEKjufWTfEvlr8mutY2R3Udb0WzDJyHcr82hNn4TEn7QDMxzMSS1dZk
EV1X9KCuZ1iQNID5vqrveXD633gB3VfRRl2r2VP+Z14GfumLKdFwbDVh8GKAcH9L
lrgNugY57gf2W4Ryvd1K+nsKICbPSm0hgq2oUEzF4cYHV+0iW+GJbMUT/L2dHlFS
JAyDcXepf+dblG9TmzZ/6+V0uw10w/JtLAgpqPF4PsWEv656KZWZEkw5p8oS1mKo
iPHXcL8i77KwzGG/eRQ0O1bN7iHCyJgz3hsU+UcDSNI5jbgEBH2WPUqncrWpd9S8
r1QLYMy2jQPuEPkINkhgwy9DpnkZivguPYUuZn0ADgdQi1toX5Y83LmNLJfe5Rwr
rRmgVh9cJogRQQCfHQQNh7MNmruPZEe6oRjmpdtlkAMLHgRQBcM6gy53gmisqrfe
uCZA3yPM+OH4DMmTyn72RJGt2S7+WIkoZ3RLrn1Jjq9OJOyyrcsotYhX4wEXuzrt
NsRvBT/BhB2rKZDVFMAQ0cY+dOWYak5hiF+bSl8pHzGWWdH2s9IldZ1YTrmeXU80
AfNY1JXxkY03fRbktGm6mbPp267cOZl5j5+d35ZTyFBxBpSew2Bd9xu989EJIPHT
TYyygjRJAD28jSt/dxxo5hpBAGp6f+lgK/ebBinkGUlosiSfr1or9fXIqlmAxCRX
pDL2gCZ1MCAn3DM+BQ3TJGTSFY0DyODFU/4R91peoudQjA5jr71KASARGbC7DxRe
/TFr8eGdtr0mDMAdMbcECo8NsQPCBWG78KldiA3pZIKjX89O9ogk5ITBu1lEFvip
k8Gn9PvzGYGZq8VY6xg/TeSMp+RuEOCpiHKU46a8ylDN85wgO9/zpdRjUWluqtsg
ISHTzLm2fpfsypgptZsUmCHLp7PwWrqhCIkae2YEBhd2oCHBdjYHug5fGXZ1dp8x
BzWlV7Zz7NebGG1Fu61nfTn8NAfYVZ8ddQsBiEnmWXZP2LBGdmQsSJ7OG8h70aAs
Gp90U4BPSGfnKrYk3BdM8NnAQhbQ7h6Ccg+jj2cvW/QGAk9psdHibaCqNnUJxoqH
YO9HktDTGoZm3Kntl3mcE53hMTnGRDQzMpX4ZHPwNoA1mxLriDBzohdwQuVvs5m9
BYSp2fn76CVrNxzPruNTt3JjaNz5wXdmx9UYW/rzUPuINH5zznm6FvpPAFH65bpl
p/9dTDstklhcBoxO1oOPMsWQwXVzcjT4d99XyeA2Ulro0zO78gldghx5GxiZvrGM
Z8lC3J60O0A88Vvj4jE+GV6Q2vgLnqLUjIU5giEYYWoancSlRYKUdpk5GgrED0PX
QJNEcbM4GBhzf0bi5O+vGdqb+rB7aURsAE6P2ldLLaudfZvFdZAwp1rECGW8hE5o
d577RWVP/cmh0wwvIqme3ilpkgg9I3YU59Po/RMwJfEy5dJJs86Y2fGDfeqEcpok
fGEJFFZvuKprXQvw2Xq7BZZoBQCR4GuZO4mb1qWej6wJCG+9DCJJQIJvrl1WElk0
rjUoGbo1PjLrojgL0MvNg8ttmDwzFmTyNQdW99cLNnIfHXsWqdgknTCysPzcXi2R
OBrhKZ8QZU7gORfYdX2FtIWUJiY3QTZ4hP3gZnvx2Pr7GLl0REDk9VbFyOv20e9C
Aqceia8k6VX8QRYWa7eXEMmUoFefjh8ObfnmOfez9sNLyfzy++cx8VC/+lebdcB9
kTR6uvlEmS0EkqFyXtM2UmIvyiKW/MId3O+vfUjVTy8r3V0Uymgdeqc9pSE9/psx
KjIws/JF8j2LyAg1VvbFHZSWWWVzbJLjGxbCcqOT4WCC2hSGLtY+W0obWQQ8ZjTE
QEDM4NM55hbhmueKnbfTmMmTh6lfasMeSv5ZXGYKf2Q65tP1NeB5J7+ki+lkOhSV
yrLc6HStVopURndyNlyfB0IszaZ0cw4H2H71DhLqsbjadaDGH1CD92y7bpYwm7m8
GD2LcMHgt4N8MqAexNhn78jQNh5WvVKzCKl7PRVfPEWjJcFg9JxM5NY2PzQqdHrt
II8laM/gjjkDuC5oWZ/lAsJgblsup+c2rkYSy0mQX5QRLNHw76iCggMI0bLIS8xd
URiVIAxeLqn78SbLZPP+GqCfbIr492YG539mlfojCK6vtQwqxalKA9XOuz4n+EgD
KITT4xEMQBFPCdO+jR5ot1Wb154ynAEduepsbfdbIQ0WDTPu76Ktyss+wZnwR13u
KSaESYDaazimeSF7/9CEAf7AkzXQ6SGXta/SefpSzrVpHDuwxxlBpG+IPhS9k7pV
UrsNYk2OgS8ntnPHASSFra1ViXkZi1bDizJn2YOQDu0RXOCe3q0uYPKOYxftr3eE
`protect END_PROTECTED
