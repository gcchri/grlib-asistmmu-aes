`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qfu8fTx8t1uAZYWO4Oz56GQ1OBXsn/2+X3fJxTWCCFy8EdC+PwbWq+2axcuk2ld
T7AtGDeHndBXajFZ32/7JzTIVsYVMnG4FRlq3XD1oNvc+kVXjbYIUWKKnylJkh65
wY6I3WGO2xbq84neYylejwpV+a/SUJHpU8ASje/cp6nX8R8M0CMGlMqqbpZm8dkc
pzUdmegoMV1VuYauRCX4X2u0khOMGpk2dXQLZfBuJVDWd8+PRPTT25L5xf4+gpR5
yUOmFBQ/3CwTY79gohy+lcSnj+e1b3Z9xV3CQIE8T3Sf9GboMPoCuN1u8xzuQVUF
nOurxnGnff8iugsHldw1E3fNrhb79ktZgpRVwfFWSdgFcWUcOBTP9n1uzBaTm24Q
M3Hb1SrP/4DuNa9zFVieJbSN/RCyjwwbFYaQ1bc+c5Mmfu0y97esnuhd0SmACEpB
CZ68h/rcMATRUUIkM4QE1i3kXMmoGjf9D3wXFzLaTfWM41Xfs60BemRjeCRK1DA5
cq5BeJrKblvQ8oSd7sH6Lozhdtz6v5RbDfovwlzH3vMhDXdP7PBEIR3h9eu/PdaU
qj4TN8vcwXX6G5+IpRqetKYqP8s/hFkr+lA/cbUMSagKboEs3/Bf9zxBbKZu7BI1
ZmtgLQkUHG4PkeI/CNwti9/YNll+beN6wZGhEF6EcpiBE2aZV/sof5gPeFdhDzA0
uxPZF6D6WKClSQKo79wJaUeAfpoZDK0Coi/iFYGY18WSovinen3OYCMwRcANH7dt
a9LM2B5r+rH/V2huR5cyHoW378k5T6nJVHU5OUe3lYw+RtR5xEdV8dsaji71z64G
Lp/Ca+4XYDijL4Jl9RVB/pKhrPPm2h7OtuBBK7pEhgS835rp/PiH8Pu8AJyyK5jh
ny/YC5LROARrtYvbCmd94YfsXr0hMjYMazSavEqvVqC8X2jnRx07HIy8bmqgFMje
opIvph32kzHQdrM+NNbMKPElJ/ytySGPwnfmUTArHEct8+ppp1/Hm2R1emfTO23G
qzFSAyXPidO1HcXQ3phLcy0OZA031SKtSQ4dq+Fgj+ebQXYteb7jZ2bWbfEEiBDr
sAq3dS4Tqka+P9/3lAUtmOncomOJWSNC+nRCKUSGSXPXgHTRwUoqsn+GHvxymDZE
6zmXTai6h7DKT4cCLTlOCDyMDISpJIEIvHLY3T8jaQypvxk3jrAMr5CBBBYhjb+e
koG1N9g5E7NKRn3ymo/z6HxKh01X4zJwBK3rDBwMuI2t/QziZeohy8wK/bF1faSB
DdeBGaCoQVXQDgXCA2vK06cUQ1vKcbYVNod2dLufjawOMd7X6HJrzcCl7y8U8P+K
lZ1I7zoymw8DKDPyJGNd2qhYHKYArulcJT0N3+q/FILcEISVCZVptZU9xdWtBfDu
vaB2JAgp1rFbHQ/VxXAhFgeemBMBLEcyQc9j4sgptL4jl7hyHX/1YnuUOGUw4j+o
2bJFvAk+5dchQXpAQip/Pv4KOjBQHzJ9UghG7di7x2mdT69WbjLTD22itZn3CJS3
m0dmPnggvUYRq3/FM95hC7I+N6/TBuUoemZDygZlp8kEbxVVc3qE+MJXaK0xOQ/q
K3jlWNjc+Kt89+mHce3kVIy3QPtkB3xe1TSM57zH/cZ3xJAk5uFr9pVPPCsRlmUE
/L4cGZqoMMpSe7v3/0hzW/469Di1UPbPFxyPXu/+ysUAwfl2VEop95DCGfBZyhWe
PHe3LA0JeqyaQhHkCmmx/9ZiplC4uVRWqz0yIDL394Qg4E7+Pd6Y4Co0NGdAMR+c
UAWIUZFzL6CjbZ3kaCO42OVo5MzDjwRoNGNkWG64DjamtI4+/ZJN0uS/+5XRNPZX
BN2nmdvTmuolfQykmGdt3s9RN871uaCDw+DbAvgHAWwr/zRVzIfyGk4+DU//Ajcw
v+rtHynnuddCufBBrUb8Fpr/g+1RN1O5uJub0sCmb4hYLsccf/8R4TNoFqIYKJFj
05eMsvRg8bw6ObsMEtGBBCLmFtTFaitX1H+RfKRmybrbz8/QLJQe344ee2ZOfql3
3jwCih3SOCBO3IO0NGoD+sPgFwmb95wf80k7g+5adSR910tcdm6glU0NI8c9hg6a
QnO7I+QJgcYVeTzf0PG6Cgmyx4M/tjk01PJeJH7LjoigISvgzqY43FID06+OIz6f
GKDuM615Ktzh9JlPV6T1WideIbUbQWhLMKcx/dbpoaj8xUumOKN4xC1hLWSz6MMW
iEvzmRW0q/P0rUnCkG5E+6qh8cUPmiAm/ypM3mdNZX6HT1AOOcI98T0x+Vz/O4Fi
eRj9YVtiW64pYropECfCE7+KcKogqCEOHD0Ul4iS8bj1qVzoBBaVFN6A2vTGRPoI
kIXNXONyrIGKbtKCcrRBFXGD4ChP5pt6n9Y043lWB78RZUxvr0bvqVQIhecewMZr
8OuANr5yb3M0GsOzfNmDn+sxWZQHJ8d7/vVG1EHna72ulGP3NQpaPZkXbTqUsSLp
poCuf03X6QBrJxrg9Z/o2qzpHq8/3BGX7N6gI8/c/8BpCANkPElfvdvo/n6PU6Ka
ARX1Ev2bhZIf+WUYWHHhlxDPjINqkdQxkNGeD16qXpet41eLO3qcCwmyy+vq3v3N
xLK4TqL4Pj1My6jkVxv/tJCphh1SPdQGVqndmlzuvA1uu/Pf4pOhZw84/2QFeaKQ
m1OrhHrdJcgPblomW52EjWhHouAJ9WDX1q+6x3vyeVWnN+TdA1yittbq16H0EA0g
CG3YwUoHRbyD20zoMiPNKA6ns5XqlBzDgUN6WBAcYkc3BJcTxvxrsatDl702zWJC
JnDKHC4Aic+3qVfQ6PAaNnYOftQnjPOnDVqjBuPzWf5rNdBx/HH12DKQpo6iNHjg
z1mAbk6ymVa/U6BSU3TtzaDB0RsAdXmTbYl6z53jfZahDlMrseV2Q71Cthn5yHoI
syfb9mMi/erRr7VgzocdHwdbJmxuXgzvAob4ed7oTs30inOcUlIWMJrWdTq00IMu
iLgV71nQC7GgZyvFEHIPAetMPA2oWeEo5K3eZ2lMdCZDu71hJT/aaThqsV+EHfUJ
c+iPV+KuUt5DGKfa4XHeD09iWdbCCK/Xo2P/IguwZT03qYooP5iygJHIB7m49Caw
H0hbLVtu2KTAQT+kPEWPVMGkktufwaJXxGs5hqAcbRjOVRnBo2Wi//1Rc/mSzJUw
hQGVVlxroLMcY27UlTfRD+uT2Qu9kfoVakzYO1iyxKAZK5iWedhpKfjfAQQetuCq
EbCCwxO+Z5Hvdj8qGhTnHr2192rvZMw6kVAOL33H+uejlOt5ngyX7x3dZgzO9zZM
okV/h5ZQGIyRaGHCWkdRUU6anbNwnE2AV527WA7DcH74GnWbOrVe8to/8wzdHQBa
F+YFyn5Gg2IVksyGIxvx9f1e7175x7BUds6i7A8NnaqRnkFzwtVuMu2RqkMSjbLA
3aaRo/r8taPIhuH6vJfuqZjWR4/qrU6OovPjgCu7zrmu27BJ2wT2sZaS0VKQ7XdK
6m8pn5hllqefVYSN7TakMr8Dfg6RxtqbmtB3HtPE3n1I6rBTA6WElVJd0dQeV2Xh
J5gLt5UPpfNlnibVEBikmj189fLvCeA6KNjC12LXRnQ6WI1c2zyREoPXXs+Q+Aul
UtYelX27FdxNpDicJzNfCH+UkMjildAxCvm0xfnMwSWZpqVsxZRA6ljXS3Z+QrlV
8A9cYNEVQsqcGvCmxMWIzsjM/FfqnzBD14Q7V0bKeyNCwAIBcDLOqRFOjZu2v9zz
NUK0QekjY2haFKtZcJtMzKo/TFZT377OLiycWdbkMqj0EAkm1NuoUlt1BmDr8E3A
5cDV4TWYEdBdsX/5TwnT0VY2bHORKDHdZ60op9n4/ox6CUFbMvgJUQWhAatXi8Td
ETotMs/nIp3NetRhQPrTiayyrRA0W6eAT0MNvlQnG3FtIzb1SIDNN5NWAIUM39YT
A6ckdM4XjjXRZyXFkeQ2uyJ2Xa4rhlIRviSGXYRPssc=
`protect END_PROTECTED
