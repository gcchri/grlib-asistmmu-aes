`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vwNjclLcqbscyPwO+N0p8I4TAqrLn+XAXlUtka3DJqXeyD9fYsl+TqIv9pLrNCtS
zXwYw1cnFSZ+7FxeByAqCKWabEfR/kJ6BVXhK5lPyHefyO9aKK/0DUmF0d7zjKcn
QPUQwe/laIM59zGefTxkS1zHHYHB9CMZ2i947yUwLet7g62HSOfjlKQkQB3FCNzZ
ROgJllPu5HU4TGJanm9nNvo5smCxhOhpS6obsYWEHuLXKnFl2934RFF8HCzr3dpr
aUozW2NCw9AoiMIn07t0qyRX1M1vlGP0bs5h4sanZyi8pIylaxkhncqwmNVZZ5Wk
aA1TLl2pvTuJgwfjJm4As77Rp0EPtu2jhY4oKHhgdAClfywgNeNkJl2C/iEDOLPR
3telltstFn1y7pFj/B5YLSWijHzwleyW59yLiCG8LUjX+A0luettwtRYnX5niNlj
6tpBZIe0Uil0V95G/A8yJ7qBG/gZ2Ut6+4KXPVSdlscvTZJvFy34B6xPvZEv0CKN
GYkaf6mTwbgpxR52c50Q5qRLU6uSb+R37ZQPfKPkm8CNh+domxMqkr8kQG4rXzPT
CnacGSRR2ITrbUxQN0lrSXwiYhTPWeMT5oqZxuAwviqgUQlMt8sEt+eRe+PY2i8W
wsrj0K6p5GeoIUgvyCi/DLFyKAAboH7uzOY4UBiM7Kafs0m45+HFf+Ik/Yad1ug8
EvFGdBxrQp3jTMZr4mNhTlJrQ5L32aF3qBL+92vH2PL8vqHf4QeQmhcbBPZ0dBoW
E2jbW7X46SJZJsJma4a6nTuxGC++jyqzstX/UzRXSC6HWlY85LtDWP/JSbrNltJf
pB20Zjuh/1QKtrSnWV6fcOYcExxYRkKU0To4b+320sqH7kr21WOFM2Cld+YkCkEY
IjPmw7Sod2lTOnHt0tHBsUPFoXJhYHoiCCNiVBRxockrwMqw+X2Itk+gM2/Hwl/Q
LG7HG7aXOT0NXFdwZheDqbVZSWiFMfYt3Hh1MeU7+MlLLC0wyKh5PmX8lXEHg1Vk
G0NwHXTwVwk0a1JDdjmmvXkPaQ8L0Tb3mGWIMKK+8NjJf5kN3406KKTl4nlMGZvX
zrG9RYFnwq96MHKtjQx9rFxuy0PTztRjp2UH1F7NQ1oXq/fgAVCnF1ZmxbdzIoG3
SzRYgD7O+QijqXaBrpf8GkanHQuB7yeS0itw41cGrOadwDtvWAd3EBQWMi1r/KeL
BwRq0lvi8c5mqOfAcdfoqlmwt6QUHnGRMt7TlS2mwJnt7L3iKz5M6i0MT+sIc+ja
`protect END_PROTECTED
