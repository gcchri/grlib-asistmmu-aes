`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnmqmR4t0352lbCu/vYbFVAJJXLz5/0GbSckB2RziFk1Gf3GS2yVU2aC068tBkR5
CnpZib7LAxy3N0/c3u66uXQEn3GUP5eseLQ3O0cz4ToM3dcQxZQEwYKgXon3R4t2
VNWOXzg3bF5uBdb2bw4T0otKFZvQLR7Y/rmsR2c2yfRA780x0cluXRJbTbf+6lO8
YAGuHMsPh8d6BYYJjgXbjwNJqwLcsuAPd2LwJyucdtwUnr+CfuR5vb304nePpL5n
dIfsXAP15S7A7aOFvZeh634/5PfIrxg7YVmfRKiPAOAJxFRt1zMIVe4hOO8KxbU7
PkC3we2+ayMhquvTPvw4SP31DoIVYfiOJLzzABcl8gyVhUXZd/Pd5qh4MyCn535Y
9pSFABEq3OnCoytHgjA5n+S2uFpOsRDP5Grt321gyZDcCojwuRZt1YuFUu2Urhlb
DC3J+vSLV3A0eAVGPv5yJBqzxgGsesBOL42dVeZhJjIqgAN5XRTlLNumr7mXpWCc
XA1tg74y/PRlRfbMSI+Wu33AEle7OVgpOWcX9kroUIzpDi/3Ftg/OGjElwdOrK3C
fR85lQsweSxQRjPILyErBcnfWb2Z/1H4VDeFCO5t84kHkWfVkPjhFqVGJ1eD4UFR
vQy1lXkWQwJMefsG7FPsSmNd4M3822niYSaCoSp+cxqkYX2uCeEsOqu1oIIOlp3p
uPVwNSOZdA904dUAKBNVJmGWMH7JQE4WTBtMdIHEUYS0na2vzgIWPg4Ghp1qKFOM
SiPOfqCsmWBUh9agCTAvfl3oradXiAeh62Yc2419oyOVo+iIi7JZZr+RuMqsIxNP
zPI+X3qUSgMpffpH47dinpgMeRVpEvlv/C+uwoWNe2t67fo0KLnk1rQ8byVMP2Aq
Dz5wlGmrnCwBQLglErg/TuWl32t65Y94V/0HoyGjCqoelOVTNzJo9MHqqNZUv2r8
raDu1h2iqyq08UdiLTL0pIjmK3s32EcR9FlU+EM2ZH6AvjjO8T5I1ASNO6cgK8pG
W7YnSgcNHo4pRMLbF2cl54eOaUU7Y+mokZc/iz0tBhOQeVr+/J/NlOHSeWU1+mqk
A0C2HJjVZ7bqeoN+x36oVCdsfUtu786gijxqsQCO2JIOklyuNdLIcRQA/jbAk0hi
5wU7aMTBaEPLeSuaorZjB0rRkqaBd6cI1fzwW6TCQc+EX3FdTFkMzS/s895LmDBV
s14fXrPWoYeZZ8FEHB/hnpMFtjSIcqCMrLH6r3w/Xj+5i795cveGUzDgwQPnd+8o
FKwt9PUgX7i/0hq3IL/KQVOVtQa8xUl1xpfxVRjmHmvQNnDn+QFmwudflJiZ698L
IvgQACmX0Vp3AI51pEel4dhYh4bzMO8dmQa6y9Fz4WjRQFOde6z0LSAQKWITdI17
fvKmtfYqj7FpuFuaNfHOXXNV0h1+tSep8Rjf8nl3jH0uqN0ytQbJWhe+LY5H0rD1
fUBFh3EXOJl1pcCrFVVbIzW+Mxl7mv2AZgcV6GSLyaCWBc+JkQ2WTqtQ7pKpNqk1
y8dquiXxjz2B6Die3HFOh9ij0vi+Dl8lqEp7qbAPBKb6RbKK/vJfhmCXsNa2FjTX
abi++aPwRwr9saCyaMq0QCUiyij8rV9K6TvIpEWZ3uwGT5q5NkNptMR1shSmcrvV
mMy08EmYBORI8Z0zYgH0ept6C2+b9CplvZdmeCXFyTz6W9H3R3wSQ1T7SJL6zKqM
QjiI9GYrR2Ds+zoJKHrnKx0ePtxnwSK0Q+cgg/rq85WnxnTn0QgIbUxy0CAwt5ds
X5OwD2mxRCfatDEI4PzUL42ZHVRC7th8Tp6+LYh7R2tqW7woo7VTiMIQ2Dhz7SYC
ixDlBqRA9ahoNXY+JXtqGegmeeenHfDiXYCkDV5QntD1ZbUqAqrkHSP5URB2jMr8
WJOzc3Y6t/LIEvoRwV5FLyJvxo2NOU/eZiAEjdupy5nLNTKsYtOgEdXtIzDWB/Mf
/e68GyTvfZpDXNl7wSY8YiUXDEX+9ZdtiTMRNGqxoMgMuyxyCwhmptboRLr9fnyz
p/5hyZHPPsoXUE7GmkRIT7ZzSVSTL+PCV9ewr6j1et6EYMYctI2K/KYlQqBEJZwl
5zNbVf9p9GXHpPnB0+c5/oCEweI8GuI0+/hztz0s3mad0FmCQCqPyOTsuOWFxN0w
MAoorJ3SNL+W4WidjbGLntWVd6ostjdVabXfY6w0wDPP4h0161hqUT8PMTX8rMFM
7eVinW5N+cauygZssa4fMjIWiW6OnHlnu3H+r9qCaUJ6rLIIbPRBtacjzvjv+oDU
GVzZ+n0zYDlRShK62irwGSMdZmh7cYZ5CP4Kn77ViLK0lvlVzED9LWO/ozFarisB
dlbMrb+YlsOLPxPOj99oVaXnYxIIZaGU0X5pjLmvGY3t8KNeq7HCc4emUsCO9aE8
3BxdSwpwNu57RpB3l+nBes5+9711vyfrY8lXjYjF4prz8DFlP73L2bD1k61u24aF
38L1T0ZqQ0ag4+BNw6YcjiO0Nij1R27Kf8MBE2DY/92VJZP7kclipnLz/Hw/0bEj
OXS11hAjeTX58EXQ5vQrDjwDxW9DBlhSnfsiERv21Rxhbj93nISEzaJO0xhUoPdU
VRlTLJW5QgjctYX/s0Ekpfs1OFPoxS3ClWOM2H8bIiLriIr9il434RmoJbg1S0RO
5e2Lv+lwBorf4npEHXpReVpDJYZblsbNmtM5xk4apM0VVT8yMmZ4SVITuGLK6QLL
TXq6tSE9boxbEzIdIVtYGElCO70Mw7rVS1JNvKbyoDS8DoHAzsVUNcDpJDmlT5cr
4zjL/mj0IZlkX301FHGSntRgqFe6qG9r1yKDcTZpI539SmSTiF61j3SKvtdjYg6H
Jif+150hctPEtvMSB/RpOg/1xYS25ahiqG/ObZyLh74M6J3ZB81G6fMBjEiDu+M7
8xkUHmbcXbd+xXpiKTYzwAXezYPIcwbtFUQ4i1GOMzY=
`protect END_PROTECTED
