`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y/SJBFLM/LYwXwXL6DAFQT3cvCrWsZxP8OEMTyBsBX8Hzg7srnJK+APpQPIA//Ki
XIdqRN4lUklMBfNruTOC59mgro534ZkNAerJDgd/kHyi8vX63TZhqwJeANq8c3wU
pkNAeJwGuAk/IF03msErejYfHfbC4P6cEJDowUtG4Xz5SM0JnNMXFbTIJrfxiuir
7j/UaJAqjAlIV77lip6bZ1r/LCiKRpuL4laWqEVim7sTM6nXnsAcEX1DdX/4geL2
Vowd9s9tXhpOdTOs7/fICRDndCNiHlUsQ5n90KG4Ofn49Q1sL70ZsF000OzJYCOv
wI1EEzvRXgh56UDTtjiKCQBJB+aU2ocrUflyTUIlBTgV+VpG1X/mbtjYWbfPNlyZ
3akzrz5usBv9FJn5fOVprBta4be3UsXhK32lFJnE5KXt71ggp/+SHL+LbuHwOZKO
8wrqq4VGWdGKwdC5sRRLnYNRUbMBdEIb+no8yc7MO8bvPUVNJulPbkzo0pGiiMgM
lngdhflynLMR0oidMkcO33YU0hvZnCrxIDXJmuTRGY/uDD1rVGOZGdBF4FjcY+uz
impobKja6C7ITYzmnx4Vn7EhR2Am2mytLhXPthcrFpOZC7fJOUM4QPh5HqevXYfl
aoJCOnHym5iO97stYFkYr5zeKWcKmSHxWVEodVFnSEo=
`protect END_PROTECTED
