`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r0MDj0nsCh2eeFU99d3WcDF3fq76Ca+nEHUjJmqdLsWCucVvUkozhRNdOq5bllxA
GtQlwbugi4aCizMYInbrWc3Ovlcry+X65rjC9uq8udY/Xa6odnB4kqcbRTnhjr+x
P8/EaFazmGqZOC4bvc9EU09nejB7eETQqhMQf/65woTABXXVYCNz/YFuu/fSmUAq
uzZTd1n+g/NceJ+1r5J6EcowifomsjqeybcGigd8ZaCm8ywQFphJNfzouLVCQtQp
+qafe/5fF0DuzXfNV08Y4JTzgjvORaCLMUysOMLbQ+s=
`protect END_PROTECTED
