`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+ts8NgHZI9s7shNHFruc/Axnx7RmrsAm5aUBrxLos4ScLJkxJ/6GhJiGVICetxx
QP0J6/EaMZ1PcFDih4R4v2nsxssaOIHpZuV3pz9XrcqEgfQRPHzdGonQes83H7h4
TYBHGZNfO0VRWOfEoCMQOYXxPfbgcipRVieNO8NRP3lIuQYLCDyimRauddrVsGwJ
bQrVk0VGvtP1uIu3UIf5X/PeuCxEx7AUs13tj/DmlXUGIjB1c8mMACylKvKZt2+9
1irF2mFQubRb6aEM6RtDpXh1GcDy1cqmmujRsuJPWO/lLn027jd3NJrjkqiNOS0J
J1yELQ41tJW2ZnY39kCrvhnhoBCF7dTZdQayhrD34oHZX8u5aKf/hual8wzKFgR7
H6L2bpucAsRJ8pjIwDPtG8wECUO6MmtXYZ3xYifQKfW0pgCR+cRixBmDm4h4Q5wU
dvKWKFxg5CjmuMfsD+lkXExPepvhhjB75EjricAoJHjdvZX2JJqEDMG81G7/sa+6
IfguZCv/qPyzWhqVkLtxj3G7OT75rnPOppRnQMU4n8YtN0z2vOQs5TA7XAF7RGoI
SLFvivwBnQMMwa2I86Js7h1ZfsPD4+mu3+RjwKV0oL9kGLHr4/wgW7kMdfvsKYPc
vwpy+o0kMsBP2ukfocNEc3twTirv1aLxWWt4IpS1f4CowzaQC3tOZJSrckwYPlsn
n+j7eP6DEdV+6jNhObq0Y3HeDMMOEnjtJBsEnFadFixRkDklTPEoPzq2pnvvYEpb
79DruPEp23Tnde/2xIF+6OsBntxCpc8BwYzvYhl5PhS8BLyCREVn005hxJQxXIeC
znWRvUxPmYwuIGgV9pfXMNskQfRVavB4TZdPi78+NBIaQqYe3wOc5EF3elI92Un5
ZoRm0K2jdi2SvCmEux88YXM1nU4f3B9cyRLEGYiX+0DGeZZYwyNTgyRgRD8mw8Ak
Ytjk5omOLnGLK3Q17LQLKh3FlTLjGp2yzlLspwDrIfUg1DjU+Uu3rgilOBlhe3Ua
XngGWYaMHRF5rjn9Xu8z/L9cAY7cLslkV6RzHcgYfF7oAzqwlHsk0azYy/tNQ0z+
UAHi3OcrsEdUSV1JK39uRA==
`protect END_PROTECTED
