`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
od4dG86//JwRHooEpoXw+VE+LpGdPcj7nFMLhdcvb+WbGyThCtKzGKVNoSVlWEGl
DJVMr4k8uDSFC0YmALuxPCIhIq0yUNjdC8uDLFsNU017MOd4dDZV6GUeu2JswA/u
ZwYFDOcly92+dDU6vSzcbw01IBjHr8PRLz2cNooaBeI3uuR325UwW/Pr8Yk5ijt8
QxEJKzFP4kMHCemCTR1x9SqBB5nfTxis92fxvt5aXz6Tf5p3LdTea5xFFeNhxCQN
gMNkFTrfZ9d2VxpeYO2q7MWmDG3We01e8XxBjdDd/CZJ/95qwWrehJKpdrBaO0+k
4LD6ymPxuVxIp6fC1tKdJD8fLu2UtxfzdKdFlwp693I4ei5zlCMyk22O2EMRako1
Vam/i2+ypFFUCghFtLMcTOUChfdC925N6PHqEuP7jCHYcptueQeNMFs18QrHPNSO
hGw77jFShYkTYgiL/nS2oW5QXzsZLpALTzQPsgYarQz5x5ChNvZ5XhjP+IGLTJae
8jWVaVrM3CLt4FDWFb03/YaIIdmPBedcrGi76P87Mg5mgVnWOGdfuHLVmSk6DV51
+IGGkteFdg4nF8/Ikgku/X+xbusdL45HZtWmgY1okzL58NA7715rzwfybqHXtp1R
HxJBxWZqAkgsijGxypiS++/QWMlL5kGQEKGFcyxu/MkNVl5/Ci0YpNXL8aOgthS5
LLb60atnJ7YonS+ZsMI/RFaRNezTJpKQAKYrUWbVp3ygHLZPRxmsWGhSkhwcdyYW
CWvIOnMDsumopTKF29jX8v1rKtwQMfd9L6CUQqbLeVa1tZdM+qUimZHaIaLUhUnY
dW2IemDI5S6cIrOHc9GYKdxB3N3D7NfFuKOvJKZK+h1r9/zjUwb4o+3WC20Klkzt
XeLdw5msX/+KAm7c2sfUAO3wCBrY+bPWSLCDOEIWXF0gHMic72u/Co6ShN5oyut8
dEioQGb54B0XbjQI57KFSHBZjgA2H6YbhIIHv77W+24gPnZ8MpXo8viUYBBVivWd
XIKuz5gHmjKp9bj+DnM5DhzMxbnWbQ45l23BMlHyjf9ReyUpf1Iv9pka5M8shzR8
3mFhFbqh1lwBqojiZ/AzuWPdSrRAxQ3Elw8Iq4gTO5+0s/7kJQhmvn8vZ2i8cfvr
IA0v1tob7bEZ+1QgYmF7CRhx4OvbEOgOX7BPCXuSdawh95BaVGlwuAONyE8h8kJr
u3FFz0ZEDHF9w8Te4kzcYJL0FhHZSWVS425h87mVTiqvud3WFXuVGGnLmUvBhYSA
0vjDpjrq8e4m7qqyqfAQXCLDSGCx3xhkVrB9pj7VrPElOuwEqQEJsqLMMMb5/kdP
12ykfj5XurPeO+bUVZJG2N2Ild5ZRCWdtj0KCtOox1q1EZ9KgdZzDvgAMm/T5tJB
Tj3gW+Gn7WeoBt30NpJ6Pidfd8KrRzHD1XLkmAGlYcd7TYiUA8Sx+1aGzdU8usTA
fyasahaW9KP3EKC5kfc1EpM6nYD8ozjg6rAjv34br3G8v5n8uMXWYaAfY/ba9koC
XOGSeECh2bk14e6INBxHJfD4ms8Z0VI/tDF24i3Abkd8X2EU4Gpo83/27rhD99YG
SSCCYbYi9cBe2R3tMJ1D2dBywPmcxK4ohxhrzmP7O4jwR/1zJGxzfsT9t7To++Os
iu0zEdFsqPJCouRbcGeJJmog7E8HvQO1t5N2l8xuGIFQ3RzapVbKJSiInhnA8cwM
UfJpxY4Xex43J1+q/gqTf8IQSpR0CI7ZtLzsxq5qd8hmTopESPqF5cDql/RFaxvV
LuHyhTjzuPqMzfy6IE+TLGrae3kkMhUHITtfjXGbwELE771BKCKV3tfsdFjMIA7o
XCHyJcJNmTUXHtV1cHAjJFiZ7EACVZH5oDVRy3icLbV1u1QSC44sQKsrcVwzQPXA
RghZ5iGOZ9XFBwo0Xi2Y58l+NiwTZWhCd8m3gu1ke6brnnT8s2bYhQxTKFwebFJE
cmjePU+Pn8vHln7aoZI2atvaO4ph6TxVOzckl7DJUbn/Ul+3aQSq1sSXVGboV14j
cTYMJfIwpim2jyjO81o8GpJOqHL1m4w6N4C9nslMhFNizarmifVDSxirEXOopbMP
PHev/tlll06J3/4kaK0T9rOEI70eegUTp10lfKTccyo5OpTXA7Tuxfr7omoioXPw
9TCBbF/zqlsE1oU8cqjnx9Uo8tkNxAuzY+tvcoELjqvDLXv8LOv1RtHgTBrN+Ffd
K+BANznxxiTOo96WJrvyqEn8CCdhq+W08n0RjehnNu+pU5dF4fudQH7tlu3FkRKB
SNkiRlkIk0o/m1yx5PH8cbREaxq9ugcGPB5fc6BJ1xgNBCFE6x9mjXnsPqjnWrjC
C9OyxHbawuT8AF/zqpb3I1pBz6uDqxT3cfvWMVF+56eqUmx6wiM3VsvHWTsvAv08
gX7TrnB7wW9YfwWgcffszy/0L9iTqZtEHvTbRqFhBWC4zQrIa6V0AnfRNP/wwlBc
F11mYRA65++wcklxbHcarugxTlZJHZiWl19IyYgJvtcc/LdOxMzVwScmbT/kPlAi
V7Fa1+DX4PGBZP1mhXjkaVtwQVewf6on6vAJby6mR3qOoCs89v+5rTS3dS2wt7dJ
GY9jh2FtsXIISKc59yWs/3VqnqGom07W56MEcw7FDXkKO1sAiquAvJ4tjvZBTEFL
qUP5q5E9PRbdIzxESuH3L2ifupMzdzP9kI474aGDEOsiARHc+a1waiHAGXij3X3T
1DU7adrKFOgdWxkbAAnAFqswjdXtJsiI9PUSzs4NpFKZm7K+S3Fu2WPvgseGfeHu
t+jmF0r9u/p+8JeCPzFAWsfuEX+Ybc/9YgjilhHolJFQmAhG0r5fpjytzrtpq8m3
W+JEPKideO8XukNOGN5LPpeL7ZtC1NpTiVO09dde3u/Ylhfzmueq/m0wSjyxGnn1
rB2cZEEvEUKE+p6K5vhOIdpgaAvVX3FBR4pKFGeTi1c=
`protect END_PROTECTED
