`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DowyHB4++dkq7Z9/YcPugbLOe3xQ3BPuuvRSy8NM5eqFt9zXnVapMhi0fOnibNIT
MJOtyM7K//oYzKQPByJzpFtli5ytTv5s4cvRyREVbD3artR2bdTKvVRIZlZQF7NP
pSLyPUNDkMC6bA4tApn9S23kXwNengp8YBECb4ykAn/2dq+2FUXN6qAt90TgIjNF
hRu52eKDGZevmCVrUdoEfQJWXfkRX8KGlBy+dwHPS1YSwGvOBA+ByI/tp7VmlDFx
WiUIOu0wr29sp1aOa6sC6XC36I8HlBs2e4f+TgXiyRFSw5QJzV4IM5ie3pETGWM2
FjTdK4HJat2rJlXIe7vkaikai6W7qOJN6rF7z0YB6s4+TGT3htzWCiS7I22eTyE0
cixPDoIvBlwXK0pr4OZVJCgA+3LZo0YaNcAa16TJpbvOSVt0qCo+tJdDCLDPcI8n
PaaytKxkUouzA8PzpsNDHM5qdDczVcNoh8QD47IVQcSr5usHy+4I94+Y1qkoMq3L
AgSFoyir7jZhLbeDGoYTfszDXgxn0ye6QZvAsh30VwtDINLvSQdgiH+hEQH2LDF3
/Xq5mlJsB4F08FZgsyDLgDN4WU9gdJgrE/io/w/mJoZAiufKn1rntxPxGlE+hRvi
rKMSBnhBXwo1cVTuKLPC9uTeT9o0DxNZIxHUWYl0pqHdBVg8xzssJfASwPXhj2Xa
JGrriTBaagJJsFuOuJNJ4ZHyDC4k9Lgu+8Q43zAe4elarLe2xKFYY7bqEulwePqb
8yCy8CaHbeO+hD/oE4eQelvwmBdsB4vHQUtAnhLy4Ap1sCsf66WNUZRiyF1MDnzg
TixnlgaaMtW/Br/FV6uMDbeHqIjOys2SRRvgzJqmvMyKqNasJn/tyFv0KnHFJBAP
KamMKztxaEZok8+deE5nHYyOqU3WN1ECWx7JU1kLRm07iL7DfDynKPibVaNL0D25
njlJxSa6SvPzyKL7oT2t++9lnjrahin6MpGkhv5WXNgfnOxF1FSXxfIOmBDYxel7
8yfPZJKLDheHGrdN5DJgBUIi10AFBrASmqL1EgRNvi/ylJU6tQK2J+hyg6Q3UUHz
ORW28INRPa3Wff33M4Ss0cNsPWT7/vL+zYhg/bQ7MBPeam140E80/f9YTP7DsqVN
Edd2Ydd4YjJIJPe8aTN/dMwWXkTwz9JUtsD65qD93LnlLAoSLiZqQCyi0rhbagev
45eS3Nontv3mCxT+DgT4bsnw9FPsz6Wp9BSmWm6edQsT+fLTqbzafLhN3RGE7aJ6
tPoeuehSwoNiXNJrUJuNjOJdGi5l6YydwnYWoJnAgqQoDPYe37JLZ1s9Nw5XJBcR
yDz8BU/rvnm2PVXYhk1PkDCvd4L/sRSvEc3Y946WqcYf2EtHD6xopMAbY3PYEx2s
FkcR34EcNiG4xaruBJ4Jpc9KrQKLXGxLkK3e9r14dUYXOpJD/Qm/bugJT9O3G7KM
WvKkoeUACLAxIKGURrWkeCxYApIsfMpJZuvhmjpsMecgvfNdXdHY5+WAHtOaNLyf
XfTwZhBmTFMWe5lp1QyMAgvR65THjdO4+kb4KS2pYz4hiVem939C6UDS/G/STQ1N
ssy4XMSbtFxD91BGAURPXdKEUqNuHHV6kYlG1k6Bb/JSI1gRwz1bOSqenLMjRb/L
b/VTj1rGp5icHvs7eZ+mnps2oxW+ypZb00+boNMB4xSDBxFMmkK4BWLP/ewQfMNu
26PpNRzwtF2kbffiW3FDiv4eUGyN5ZsKamB5lkYuVaDB6LJp4L8OIhRU2RktOK3N
4naj15H7Up9Hz6Vsd2JqPbM3IwWfrQLI0eE0G398KQqtEB2cjAMNlvrr0KSfTeEj
8cRvn59cTOIWztQzWg301ynMcHtWX+FFO2rXb8p2vLHGXNUXJLmK1vaBO/nrE8oL
KFmYwzin6PNjDawnOlpGbg==
`protect END_PROTECTED
