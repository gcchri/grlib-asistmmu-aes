`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OhV/x8fot4C/YN6kx8+VKDOxJHWMebW21SlRwZRI+gWx14xxyhUygEp5/bAHffS8
s9UpaKyEiMH3DpO6KNO7+jPYfZ7pSBGlMXj6P36FRbxorLTAq58mzUp2xoNKKBd5
jRRNkbKGbzuBBno86J84gVQf/U0CvEUSmSO0nhBJTtRqaTlWqlG2wk4eCEnU7MdI
vtvzkEmcSaycNJf4/xALEzxv+2UFreJB/xGTRpcKIOxQRkjzAir6kQ+9MpCqdhXT
d63Ww+jsJtt0d/lWiVd5xZiVINteuDZgbCQkTD3tBtJpFWNaz8zNacNIft7Wgo2w
RV/0ANxW15akl4MQefBFNlMhNrHNTyowFq/BCSW5RPMIYkbaGZ7As3okvWLBdfXg
`protect END_PROTECTED
