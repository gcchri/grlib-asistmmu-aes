`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kbc7MWb2V0ra6zG1MR7AeBOx6nkNj8dlDoMscsRRIHfZShBXUpS55oOK1cXzqRS3
Jk0WLrlQq1R/wEe0eukZYu9+crM9E/9x255H89ot75n6G+RR4aTsoOXBB3+ZaCPw
wBQmRNbpBhKDWjONVE/L9Hlg5vP3h4g13zsD97/tymvQPizyaC8LOpt3b3Ovvd1q
y2UwtfWpBtTze+b+bbjADpqnwP58HhAsjK6570jjGgFZSBPYHN2aU1hqqljZ1Z6G
U4EICDWa1S7v0+q1mzjlyQR2gGkIfPm04mPpGg1fMKpRKAqAnCGhpD4WfDCoozPA
sasNoIfAhqe8CYhrS4AXCu4A3PxAJEJWLGdPE/wbwVpCjhnqU1qQwyi1LSbg/5rQ
ZjGIjBHWjucD84Ah/h1ZoK/2jqlZTvkEOFIIUXJKQUFP9Dod+s3ea4uxPTNAWrrc
6zx6TmGkgsiNXE/JXikclCc7StVYzro+uOJFqMcsWTk=
`protect END_PROTECTED
