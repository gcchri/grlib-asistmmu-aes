`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1vaMsdSthYQRDM9N0vHLYN0lXj3+xYEhELbaYeS3rMwB7xRwFjiXn7cWiEzoCtn6
ZEvOEpJ1frNFGH+8yUjkRz+KClo2GROdtldtCGrbVmO8h/S/sqOMsM0eYEEdAv5g
5gW+1mtEKFVpzLE3DWD7ppjNLM80pB8BGX304BAMUwioYjXzwM8H0Gs6YcwjN1xg
Ae5pSda/x5/VC21LnkXYHVtE29SrXhmhDtpDnNSHFESbszI8W25oZKHP/6mxtGhp
b2PdR+wsoIGXIuTKLDGM1uoqJFcbR+JXZ8siimdYNYChJJ6snmVt/kKXeJRDI1jR
9Q19eBewsmsak0NgO3Vg1QVEFXYnLDxpXpC3Mi4+pej4jr86dDovsBNPUH5D1GP7
nzSbgkxF02jLJLDNu7NIrCwC5s0MZAbc8/JeT/15u5J2ZB8g6T6uH8+e7wNaNpx8
Og5XXHM0WxOSGCQm2MvdPCAgGq5c47CoTh5fzH1BgUQ=
`protect END_PROTECTED
