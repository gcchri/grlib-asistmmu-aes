`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bluY2wXzL10J7Omtf9DY0rqg+4QiDM5L29wGTlQjXw/2ADJlANjXaHwGKsp/SI4W
wwK0Jzz2GhTFij0YlMsX33TtIZ8Ah9ern889dNxFA1vH1MIbccA8D+wIzar9k9o2
d1Lt+jOk8ISnEWaQf9Z2TYLH/Zdr6KUDVsWsD/EMJyeopRvvFbrikiHo3kYTpqcA
+TInDtqQhnf5wTVO5D+3X1xI4Lg4sfT6t5rp4O2l+WCdBPlE9dvCYUdB+AztKR71
dn81CHIz5cmKOJPbIy3dxbSio1z1+hw+0rtk6eUpUSm2M/lh0ea3ZGU03CmYTX9F
SwA54RCEE2NYSNLAeSPnTjk9pTmICVkcfeXkxPzDHZyrhTxKPza7mt5QNL8tnGap
6SYuFYJUtNpZd9VdpD4tWXeg6d0p1OuwaMso1K5BeQKdzzNLyV8Br2gXrqE2xtUZ
rHSk/oU9qyNKP+fd74n4Su+cIA3GdaKAXl1CkcQRIQb/9AYwCG7koEqrBexqoz9a
QWwu40N1A/ur673S0PEfticALbKia7BKtEMe8gym8ST1LxULoEfUe5kczTgHe8Gp
7osdOo3TVXBnzAIOcorC+DRVAJQ7G+3rp7Qp/ncSEmF8jKUt47VLgkUfyzmNemAO
kQz5xVx5KxNJXJfob/l2H/HMXapyQfTFuOfZF98+u6kOorlK8bOaFkBCSS69jFk1
C8v5H+Duoh92/PxZZZz25TqcsFYANFvg6OEj4U9N4BolsV0bmq14XCkycPD+KZbr
lOdh9UNZxZ2wKzat/kykfh1bYoL5KJCcDHp772ZB5sckX4n5Cu3wTq1MnlvXTdyz
+C2vunyPAnNR89j9la8biuzgoKDhlGPhLUyfanrGcVwBgVCJH8UX5bEcMAwHBeLC
81afKjsLYl1HNULj6hGFl9SJuQuTtQe7+Xh0A8NMtjPpKxiAFGre/Ape7xjlH4Jj
AmG7688X+rk0JeooPJ3Llc/8ZK2/mTN8rp92seldxYkxRYH8NfIJ5XUq3M4IO6pj
JgoAaUUZdQM2DeBW0szZx4gqRAYCpJp81esxiMI7aDHl0aIPvGGwhZaXrS6flawB
eWp5bWvnKZl5jTTJGzTMiiWfFibCGvJDoVBSJbYTKvhIsfaVEMng0R7aZq1xY51r
AN8j+8fgCbJGG2a/I4fnwVa1rJdzs3V+b0fsMRsvDm7cW3pavpWDq8QByF6TOVlA
7O9ukpNKsv0VXkAKczD5V/kfmuItFXlwFaORTCbJqxKE1cU3P6cX8ZclqvVvjsvv
X9/cBXOK1zCEyhda7Ze8mueqFF7wmisRlExwpDPJFXWmKVCnSTScD70kOMo3OFwe
d/H15aGxffSm1TAyV68V7e7ItwsMwm9akZrMsw+J+eK/IhH9vxuIuwUxQUYpQ4PR
Jed1dJ8VELthE76+wuWqPuH8OWufiy9hySBGB9NpQ/qO1kCIsrFfrOtOEUTpkIhH
0+VvriZ8v2uSPUv/yZo2trbO2XUF2ec4zCNSQZO6DvLTsl3EBEf5Yuln6RC5hqsW
ByvWg7ccBRq11tfp+gmI1vzotX6bZadAdh/uhxCjp3KG6X2GfG+lvFDa9ASLPxfX
uU5Q1FCbVaHY2/VSZK8ErzF8fsdpGZPm+MEHIahynVet8pqTOuKjHlpzj+OurIMA
q7EzoYPWZNSe6p0vEee6Wqmj+OXaKBKiBQ2ZESn7kjYZeZ3OwQExhwhOm5JI9pax
Dtnr09yqABh01V27LiuR/x2VUBK9o9S0WnwrEQMr2BroTzjgv7a2EZTZXlBVyG+y
Zg9Vy/f2dFlhIec2HEBQ8ZV3vRIjc2xe6slhUEV2nTyjXSBXoMHOgXiaFMepUcKS
MYrmNMgJh46oK/EReiz9teexrz6Wdt6Hu01Pp7UGCh1RIiaz9guP2HzJFDPGn/0a
xIKw3dEV0bWsCesM9Be4U7Afw7YWZICkpQGMmqfcXK75kKtlUf0xPAdKVg0V39qw
nSgpaGdspW4g5+ulY0b5hSX5AJ7+5pvqTofd0F7Th3QEakWgWGrhhxdi6UIwNmeN
DQteKQSqGY0msYECHTExg62/F7u+JcrKTwWjom4Qe5r+ItZHu7zNZWgYidSb73qF
57PmzOdiNpyv4MmssgQ7AN6YC+Dj2+9ac3EsxfozQALZsh8JVDv1/o2DaEsBHodj
mkIJdvlpoqZ3bEF7ev8djjo/ZIiEpBC1vFP5MgXhs3R0526NKKmUTvcMAlPUItMb
8uiwjxvRHHoi1mIYh82JU3TdhJsJzZ4838ZkKqJ02N5HUaUxMRq+0SWXaAfndBOV
Q46R1MmipMGtLRCPh/BfAbPIpCi5chaoxqQ9qhfLabbyHTroSqZnFv1Xv85QSDia
57XuC4yM4bLt4qPTz6uzp3YnhDmOH0TdlnwczeWm8M1nrvMym4+bQPxEJWioLRqc
uZ/YpWgip3lBP8YjzfiRio65XBWRNxV3hr2Nw6Q4lsMYSTQ6Pd9BHrQEzgdn2ZFd
Zv6bbvVYfTUHbffPk3PcvCr7pGloKQ/mc3dWYZ2GPyntdnCiAa7CH2jHvQiVtrUx
lKG+l7mpljOA8d6XpVD2m2yE4KBdlDIiHi9xQgWSKmUtk6mOBtBe2KtovDFKCYcV
eLTL6fs14M4SZE3T2zWum5Q9DYIAaEZLumVGbj0Jx1eonk4OTU/LNz7ZfMLDbwiQ
1zBh99j4q5hJbu99Tyhsz2e5++ASlZpZ9IT7jFLJYamvQkpZiOiIuYDFBcdtIZuP
b82gFWd+287qtUbHqR74kc/ItbtfJ4b4DsFnI9SBv26qHp2NpWP7+/7UmxC/gxXm
gUDA7zGwV5uQvHSUrhmOkAKNOiSC4ETgMYFd9RfEsLbOpfZLXR5fR+WfIat8iEMd
+GNFTZ8pwsxB0kMWqqRLhmDA5Cw3M4rarrQOOuFmW0tPbV6SebxnIonlBtCCmUPh
MmMCZz4R2Rg4/lgMl3G6Wc/QbSi9a7sgRfvII7V04z15ShoPjeTDdaTpc0WR9Q4P
YGGrdbpTiXrrMLSAk0pFYIrRt1DEc6C+1kpxCszcUHMeibdVOx4pfAJCj2FX/zUj
w8VAnMaOeSwZeEXsMMQ4/RzOKc/1mvX9FwXgj3I3nIfMv7PokVfvj79479QSpcyA
QaKGU0mq6f9ExWzFdTgFpI3PtnAYjTNvUneaSni9Ivshaj4ph9fHdjhrlDO40w5d
ml+ntITQoinSwN9/351r2ZMRdyMtXJYQ2GR8Ek8jIqNqv+Seer17R/eyceGfTEGu
mF24plm0/GwC+PGaPLkizPAbWhLf7UMLtLHiWBojd2Lok9SH9OoVrX3dDiQOyqPM
uYa5vmmFjB7+YULsmH+yL1ticTXUpfAjc/RDIILJV9sRL9GgtO5ed8KyW5fMhvcn
ABlfR0DtL5lWu8Hq56SWlsNR/Gbh0HRRNdNV8XT/l6JGjO9V8HeAbUMcqivlp2y9
DQriimWXFg7Yl1i32+Sw/jHHn0q1ZwV4J5xnBz9/NtoB2qRaRt2/d1mrg4hfCCHR
bvD4wAiaP7hguXRcp7MGcrRDAw6m93ikTuZ0AQAZJw/bKqthCESwSSODrt2tjjd/
GsolbcpKHozvVinSEfDC2Rw8cSbuJBn4TVGV3xZnvQF7N3aLewB71/HWMCPsJ1o6
l02d4wbeSHHG6Z6HL1vMVtZmfZy1NxPKvGJc3KJmbeZykrURDf1hu+6BGcC6Efet
Kr6s2SnpNRJaQ0NSwPLQ0m2d1ienRap+a4ip0lPN5LxkLAG7Alj0hgJc/bAUeQwT
BXH+Y0mHqADGZqV7XYuN3t2zr2FAP/pbR55KiLj8FRtNNKJyDBeamfArKo1xw1fE
Md9BdGNNuR4i9HdMcuvVk+XyNiGu0CjHqDO25l1kmFRPNHOC5XBezAyfytDPrq2Q
dUJys0fzN3WPaO4pfhbqMADVTIVvJhx3b2aIr0/eGXKxvP8it44WSalCOkcXTLZq
NZyHhglwOo9cS0A+yQpSMDvP+hhndVm5ONyufNU31aLEF7f5TXSdhljSQ5yzEnM0
1RSAWSFUsQGLI8UxaPMVl973BVES4wS5CXwPejcbWyXZ9DVWCmG+Ee9y88CnuHlg
c5Ht0w83Cyk2g7Rt3tyDsiBfb2sR6lE/lLFexjzikN0O/eKnzWYRpFnPIuHXzFLw
9T2XIzO35gv+Rjo//CyDl8LUwJ6tYlGF4xTq/4MJ+26pXmRnqJyuVExkCqB2SNGX
yo244Q4rHrjLpiabguMdc+pg1yeDwOIChUzcVHIDo1U5R8VgWRpo6HkIyJrwz280
o52I7zHbq4bwFCciK42TLJzIAlpQRBtPxS4Wxk+RLyBwJRpMUeeNGgT7+n+jS+fb
+CnmFYs/b5nRwqwfWEtMM3Z/ruAw8JiE8CG5vVXe3JnvVUtG2rb+Fap7gieZPe64
W5GfZgQwYhRtr8w9VmrLVsq5swmnln2fiZBqqco82EIKiRfRtDXUehGRsOm+Gg7c
ufA5A45ZQ3rpRlwGtLtkQ/XR22AHfFZ5tYiYv6270qar0POPY3+lxvDbL8kecCYL
akL+pk0FMnY4V3BYXE84lNT5AFjkXTH0hOXOpFWeTTcAPUwhUSf9Mxw/IESd8jYU
Ahv4D1kq9rr+S1b1bhZtY24lJC5gsBhZfBywHGol+0kkNNcagy7z3ERuPiUHXrAt
9gFSbx/cWFACStCI6yLoMESfz+HHQHfk/glBAfPCrIUPABqugxbNatztvvMjgtUl
UVr93WSR3cHiVPMvhf74MANxdIeLQIPA8QQ4YZtrUVqUCapkZdQ2Z5UZ9/NJqvW4
e9zH1NcIH5EEBGw4nXh4F6FDmJTZiNNp4uxxCfncw1YiqRp/dl3nGMbDdmQVQfTD
si8NNcspmL4nsn2FiKWcqL/PT5EFnyMuQzbxaBGphPBM3Trovg7WamyOqdD8CMD9
KLF4A0sboGqLzMWvuNX4NfZWsPJgU8ihXYx1EZ1RAz7BwF5o+WtqCCpHVp3LRMc1
vaVUAy5L2sPRUGTMrvI1p9c5J5oSL6cxPRskdnxPwdw5Fn4NV1yuAXSqRTe/eVRk
LoNEYdaYjcVHMq1vOL95XVNzUf8iGZBMy0EBlkH25jBcfRQMfnIGqYSY4LS3KQad
dzNMxItKM4YpjDV08AvOhFOAFV/L3unhgzppzV3XzvaVGjS0/lZ6OxQHEzslQJoW
UbTyg5vNPO2HWLp6NS8uobMx6LiHBhU4w1uY5PMvfUhZkLSXjCqnr7I/MqkUp6on
Rz1FrdSO2Q25oKO5FMwMxxkONhywrGjxLI23vH3q3dWeUhwjLJs4KBPoUrDTT+Ho
+m5ViV9Ax7rc029NHJHIXpVhTgnM8K9MGtyOyMkwX224MTeB2sOP23IacWhoTtow
6yuy6EMtYg4WIQPkJzN3LLu2fqfxmNBPpG9/UaOxhT0Cq3RVk2Bqb+sqXceS1PJ3
Elj9lyXxR9sbF+1k9glZaUy6LSlvGO+p66oiwR1HQxY4AxwBhFqlVRLhdMQ+wYx6
2s7QtrgYdVcwc2vcn16BU6E9kyddfE9rivtbreIMCU8DZ5iK4fX1R6HANyeYjM14
3ElktjinQjS2XiPig0CCOXJfnIorHzDDyEhECQMCTlh5OjWDKqmXUw2W1OWb06cI
cigOTLR2aJpZJXoEoYPJtxiic3nlj1hU5RstAfoVaGOSXh7ZLlD9qFLzrMxfqEJP
aYOIgzhndgMUOy2T2pmuW5s8inFjO+ntOVFIbogAAso2ukVxIZE0zKCrd6JwapaD
TGFzY9PakhMpPpIjbNqnqnXFTYMya3WWIdty8LV57jE1szqYwjc36QW9Ha2s5E1g
MRGspD704hMgdpDC6s7WF0iNPmLjKtvnFszQUvk1uGC6WoGDRjt+3fHkm2I/ps5v
WWggYnBMppkSOS2MB+vfYZ8tRHeuMW7p+t7fd855+Zd+MnZHkoVADXPomO+/SH/0
1tdUTygkALP/F6U5Gjlq1b/OMF8EL24TjHj+cFpvmMaNPEF1t8RzqWXQh2iZQ20C
oRPKU2W3WfHX571+VyeCYYD2+pSkAGdVYo8uQio0pPK9KS+wiJSWy1RcSb0mj9Aa
oSVeTOXpbGIX2F+JWOJIbrGSrTfeCUNuuFiUG72Hchhz60dd5XsoKxVw9+EVgVcT
nMJfFKM4cXO3qjRJtvePXtGuDOOjyBPLC6tyUkl9C6I5Y9GLhfN6g+BpTUke63eS
9qHrMpFWD0K/gfXJO9wT1QzC/2LK5v4pOaOXY1ISX3wpS/pjFp/t2Z2hpTz6HiR/
K7haMgp1IIB/w/3QZLuUhplbZpoI3hb7Vam62ZBv7Ef0evsjzxshWWziu/5CDFlB
FIqOUPfqk+yF56JvHi3UulerZvCFMMYip57NlUUaX+hUEy30onkmcW+JHYowjuKS
sdfYVIuX21C0cSItCkpmHtrIlVZCP3o07iTLtL4hEjCAQY3Jw5SwnzCA4kTnPQIg
1+2ydkF8VzpeiChLUgZV+DA/w3yQyxPM5K293N5+W2mk0ocgrxcJ3lL82J4bIU0r
SLUv19LUAuXXnelb2vC8QQEYE9v1kizFQvRx8BUYZbdB/GDn4dPTykG2vzVYZqRz
BGarw9mC/4NuP0TpekV0LYde4tQHhCiZae8aic2gdiFp/r5MGAaE4KFzntZU4K2X
7WlWvR9C3IJGDcvGwJHU/Qmisgojg2l+cS1AqWf95AjwWrU+0hN0R2LEMfngfXBD
j7RHOwVBdAbOLJohOEDR2BvAmBkrgw4duMh3o8U+KC/34TceqgoTwunXOXXCR+Ti
Qs0cwyDHP/TZLeoUhJnoYoUu2Im06j9Xcop2jEyJP790YtqQ/f9YS984skyDbDrv
dlGGaDm4HyU3m1AIuZ9sZkdHJq0q6CO14LTV/6deOnec7C0DePs3QS7Ft3LXPgx4
9XGCCOWk7QUFjQODHIfjS/VgU8g1BjWxjeNR8qYPx/+gHbAfMKRdne8fB9Wo6Vx3
NAERA0k1xT2K/hOWza3hyfMUy/Ckdxj0kslM2xIvfhkMdJE839+fkeyB2FGAW0Dd
2+oBybAI546zl9DKjWRAa7jMiRHrJH8cqxCH6lOulqMmU65BR1Sf+83BwtcQX2B0
+DV9F2JIRt1rrwu80h3+X9DWlynDVHToYBMKPmode+0oFX7xJ0/OFMNOSixheafX
jTzmsnHmKfFbr0PjyLlafeEQuFqmlWndy/IPo2orZGa9eXPDo5q1qJnXXXsw5i4p
vudQIUnY7lAAhzWgztZbn3kvmrxliyyYot3XNLrKUkbR/r+lkpAKaMROfwI4MBFg
EeE7UKssdGMv55Sp5TIgIV5hQ6klEWqv+gEroryoVJvJXwbSmolhCFZq98Zq9uPJ
hkOJIJJipgYQA5TBU3yFaHLP5rFxEM4KBETeJQRCE2Nk7oPG0pRuik3Xn3QEzH13
7ec+7BwP/lerb87zYP3NMZhgIGFUoYvlWNfQeWeQXy+Dr1Cqgyz3rxVol3eCCtPU
9g6/UT1HA5ecSXRtt+NMI43sI5XbHjorSKXFfZKPPbZnL3b6VmeERAdINjOGvcxs
MZ+y+OSmXVOUY6bQmt4aq1RO+GrfMK3ducKJvVURyaVghxuiQZjB5JNzTdkVqoEC
02PPu3ukBmjJwHg1vMVw/4mRsWF8wTqLEYMpMKZR1iEkal++RtDkOZGEo6Zn036R
7tEmQ4dlMXZHZ+cj1x0Ac1HdyApXORCzjge6lGLK5yZ1cb18EAE/OZFFascQC39g
dfEPNZvCk68yICiqGwzclvY97SivE6dwZeROPoA6huczFRbGfKIRuvh2/KgzUECQ
blvqPdvvCPGam2ThvzFk3f+eFncaCBp96WNz6j/2c+qUMA1bkFHi5GgoZTyHYiyh
sPgAR0RXS6FXYGHVqecaO+XtL4qO4GHmUl9YUAs3nwUpjOnJAvBv9IouRrpCxevE
mL7eQ2ZS50cV5fs7XLw6nqMNbE8ADVyB+WA3+fmavprSBopU8VVazE4sOg+fBxxh
++WMqMCdeq9ZoASNbM5Qc8UGzADnDGkE6pe3RpcyGT/elk8gYLS+A5mzYu0vbvDa
ASAqaOLp2rSqGYz5/yHNo+ei6zT7EywgdsBuXPI6Nlkjgr+FUWNb3Z/3j4pm/WL7
LQRFbT3jOBHBVduPetifY+5JPQw1emrd+Yub945WBTHr+rjZRig6ceCcGx2vQTKC
eQRKpglDPYOOK4QhiRTgLErYoMmy1IMYAGgRTr71I1stojNTO+yv8EqKV6ytjVUr
7J5kIzrWztrRrHrrjSjeSsU1oZvJ3fa/YzkluDEBcf9lLTJj7KEPpMNrPmtTEYb+
XgAWsemO7zT0KGW8H1TCCVmy/TWd1UlRMR4c6J05RgHkLypgdcNYt0VP17pzCsjy
Bn55NJwUrZOyB3vwxO0juPC1pzbpa0DgDjnxOR2P5s+hg4/cgXmNnRFq6TCXlI9H
IZHrlzcIHULCn0ZG+Gpy2/t6ABJmMKD1VKDehQAq0JACZlK6U9VeA0kNxhqbvOL4
lfNKuBW/6KhzZVA8uOBvk5IT592mKTMYQPZFpADfsGd90FUkki3ospFKoTgZAPWz
Zu++zhPigt6Q9or0iPy/6gzsEJfUNfA2Cy1dSdy2oXxXHsvWdIN+IIRAmu2+B9ul
Ypj27sjmyvRXIzwrF8VUkATh8DPvERp3IW2U5u5poPoqXhi4xgiSwYyXdnbAfnui
ltG7+0F/UCESrcU5nPNHH2eLwNBHVydmDKYX6WIUOxeDvGC+wRSg9Vv+eRGGU9Nd
daK5YTYRi6Dvg1VILqrYHOT7J7fxqGCL/VslvnQl+zX7O21q+WIJ4rpz2grcoKUw
bDTjNoEUdbExJBwSP0eWZFpIQMGIhB1tywgMpv4ETAPGE0c66nuXjevg3ErcqAv8
d9i9qAcIQOS6wfkUytRA8BfzEbQj/2W68C/tuI3AJabM7b0MdVqSJ4ZVxSv/DemE
cOi3H5kcLrDU58Ku2qJ/IA3ExFkCSO0T8Y/zsoZMC3hod1j50TcN0XCBuQx2a8o8
PQMghduYLeTChs6BJDUJiMiQeuDLK7Oal8lbRngrwYZCYMzEgi2gIGAT7vmvNA+q
7s9Meb5yIhj0qlJts4fN1uoUJ1sFDTLEsSEm3C7q8vahr/KcNno+LEV7jadOTNPD
o1rR5V51RLOEt+KazpwGpqUCslz/V9i92Kruj0SpnYKqcMi5cCRrg4bEgayri/RJ
J5GIfnpY5+SBOKdjd8KS7RsY2c96ONmV3Q6Mg9jtkF/oWQ+HBzQ9a+rsV57YIdqv
Q7K/CB5ArgZCAFoW0QatWsYMs6VUo92zfSNja5jQJs0DNokkamfXjSRacjpgOGrK
s7X4jiVFTsKAAxbSAKRjwNRj4VeHc4sGVWNr7qTW/mnS17xjiMAPuXENdxNhS5C+
bae3JFUNWASmqxFOgFGGDYwA7BvUi3RLFiide2/pT0qCeGY8AKnyFwjr4OmZvPVN
Pnovcb/UkxYgtX21V4vKboMWC7V3idGhykb5xoiY7Mw171EohkFMLBfmkHbd41Fy
deVhDrbVtzkDlEXkQaD6BwZidzjl4ij30QmH5O/MGOlbsAFaF56Tp3ZtvuJUgZ2e
5WKMjWAIe1hU4zewo8xUuzBC1i2Nr/08qEdYHvdfc81NaFvlbVk6/r6Cu9u9dPVj
MWNSLid8jHK+VvoX06+H/iMKEtlvlwgHW6hYGGdyRvCLSnXLnWrMbSD7eOdjUucY
+yjIlWvMek+PUtSqu/IqbqEfYJStIS1yHzAh8GmnzoSBlaVvCPWyRrPGGbmMsUw3
qoJhtk0TN0zszwXjXRP8KBzfw8XsQlJxdynRzWaIJ+OUFeRrzvJpFygaLyC0kHel
b/5cIMsI1lS9DvwgxYtfA66GICslqrVdor3H1kAu+8K8W0LUWwBejvVAsvYJTAxn
hOdydXmtDg6LffSam8YU4rqpe3PN7+pN5XJ3YkS0HlD+zf41CfbBihpGoRHuZ+me
3GB0BN+UsbqDnUP2haFFuKzEgzCNdVrnh0R6YMim1Q27XGpexfQL7wCIsbcarrmO
r5dxpJvhJcuZ1S5t3GFKQYBirMBEh19WCoBUgcbsZDq1pn04WbPzJKRwEuBPsCe6
YfnfpJYGtLV+aVnlXiFovt37NT3h4Kt7XeEfuIsoRu2XpBEp7Slwb/+m4rfmofjN
5Vvtdbo1mJdU498CA5cGn0krNPl6YfyBQbglXDt1zo+8ydaRmEcKq2flDSxQz+gT
gkbKZyJ5naJ8EC70fMxQ7NSks4BhwP2a/GOMIzLJmI/B2zlHyB9r097GPMpBF0da
vJME0VPHkwlKjjAWE2rXwgsVkdIuTXGSG4P/zP2Yyc1F77FoYBj33wfnj6Bd40nb
44v8ikqCv+eNkxtRsHRN+WgT8UT5HehtCA3l5jMb41i5E2ixh+iDrYAaXuIwacYa
fPyf6fkLJD6tuCadgcT6hpP14SqIq91+CBGDxJnM6j3fvaXwLucrafDgk5N44S4P
d36gsfF6d9vZIzi0BPLRjBJag0vWE1W5DzPl8MkWz636UmZ7Uz606PE+8mXur+2g
vhYCwSBcawUtppIMzy09XEg6CZQH7QuhWb/KVDSujoOscfG15YwAZ4BQ6vpysesQ
y2ToqBb2rJPvPcVkVNo7QuGJHMHjr3ji3WjzEHJp6RCXv6pP/Q5nddJh7BOpKQtk
opQTL/LvHNhIJi0QMgS8KOZ3Z6HV6TaaDb/tidYN6GgDluMqiyrMpVyXrXxph+so
W1v0zo/Ey0fdmcGbkHq04gprH4Js1UfvVTxq2C4CBG5JjadNf8XO9j7qj1v7xhJP
te03wMVFmUsm0kZ+Ikc9KuWi0iQ88GswFo03IhIIEygOYoFsYWKp6TV/1J0ldRma
S6JSm7AYrZCPj0Zm7VVU43HNL/eCW4gZo0ZwP7TydNjqG10OYrj/BLJMy76UppWT
Dn9eiwkweH5AuF54DT8HvBmx3Uky/4M0ePLwxDM4r69KVNgc4DmJJEBVm17pXEOy
HbqEM8yOfK673/dFp9RccyLTGlG7dlo570dFV776Gk7SvCMzrVcznF3TNVGSo0Jd
qUbqPb1DFI9pq/05LaTBCgZIaoP+itxM4oM7ByLLztf29kaSy2F/awYDQYSUE5ZB
4dyhrvAhFDovFU2uxXkszgId9CQ+Q/ihN6EUpxLQsFmpoNZeUao+nlgJxIq581Bx
awpqsxmM24t52q4ilhXzsulDo0MEoLvTjegy96gqKNUpf4syEx9UjeXlFgD9WceW
7Zz8ohTcD8GUbRdVTuiRTtUcXLj/aygvJyTUZGYUry3oXVN6gQ0SCWw6/t9iM28Q
i/oVl6dXEtquYraZBaTCLqqEcn2pr/egHOyWFhJ1kTwZF8wSlnDEv63q5xDJOjQB
hhqB2xr5+7y/19S5fFaj/G5R51N0XhU+c3Bhk+9Q4Y7kJG2KwkLYo0MckaI1+Jea
wFAt//3UAzHQfNRF00DyGFk3dWVnae9+GTQ4bAQHCcYQJCUjU6cms9IraZmn1O+B
YgQhBd5DuSQhPS/5lIaQjM/MQu2NlgiDLBnGfx6FD6cpkNG1RdApMK/Jpr273Hnb
11ehK8AXbe5qeVqSCJulCnjqWrjGqMzm820YipU8//qduCHwJ0CNIwB9ZUYacNUX
zuUVj0XdliDJCVni9MAw+nUqBxA7us/xPSIBW9BKdkzO4eb5b7ILd0B0Tm81yv27
skPYtNwdrbU7RQ6uYnmxLz1LPy2xaut1WN+V2FMaWO+bB/x0k4cICQcgWiAinXR6
h6Mx+OuBYPKFBfalwGYXdUK25bs3PHa5EtrhQ0gn18tu7xu0700OucK8EkCy3+Ws
TlT3Wqt6vaC/GKKExOkP2+Mrp1o6bfySclRSSZgXMvgRY67Tx1LefFDkfJo2j86A
+pqQUdR3kLgaKi9S58x/RKgEc7dNLvz0qlvu8WXhIQdqZck/FPFgGAfwBGfVRRfr
CDj+SFY02m0Klim5cJujN7et0LAyh3HOfkon7U6AMnFwdhZEtgRxE0Fb0Xeu/BT4
wK1Kmiw+vHWkDt2NdN3XGEFxzHOgA6QuC1XUQasr5Y3ntoDVnsU4+j7OsEy364Ei
8fEfy6Ne9/sq5qI0LEnL6pO81hW17XdYmTO61QSSq4RsyYxN4WbTbNfX2qWNGWPG
HwzHbbV14ZpNuEg9O/T4F2MB/FlXkpTThRWYBc4MSxI//zCo7HKYDfxvq3Py7X0c
ZUv5VzZH3vumYO8lW+vhBKMH/FU7Jp9vQ/o+o92AmFz+ZszQjqZ5lbkH938oXUZc
dj7KcU0C8KtBz/oh6DiiRkeQcF6mZSe9w5FIw615mpCBUicDXphr2BPLWpgWjGf/
X/jaDbrh1KBLaHyvzzC0pevH9/ElflXK9nmBIdRWrPS3VEO3OTq3lS98lhgeBuoS
8pCkA08KmduykmJ75kwy31xAMXn0F3OQojN3lFucACY0hZp9vdSL1sNdTmWrElsU
tHNtR3Mp7m3/XMkiahMSHGdGLVvAUkASEWXTcJTnH/RMZV177ov9o5kwfNzf1gNE
cQxEDhhME44vpeagJoI99zqQoBxvviamzeKcuBKQ34M2jHBxPgrMD72qrM04xCU4
9r8boTzU7FwHo2+hJSY3T7bzCU1RboDs8EcCixs8Y29rybn1QbmigGOPV1aDOeyl
LAbrYnFfmkLj37fis9BuPAeHSddiFXtHzHWv2pFI4T+X795JxoUr2ItAm6EaXESg
e273CEZDuzRHumrigAmiYqiiKVeMlM1bsMLBq8jDDqPCa8F+pWe7+sGhTT2sgk29
tF1w53smbMBisclgDq5G9vuVOgrUiMo/2LrtcrdXZ3CiqoVpAJHiC6zJgTFLXUNf
nKl7s2ntrdaaDt2JiD66wESqhzdIzRqQwTCgZRVrM4vz4gBQE042LkzdKPwNPpN2
rIZV88oIpuYRytqhxwDj1ty06RQ9m5r2PiSfAahFjDFk7f+GgcOyyBZZyv3cGytV
sWZ4f5zZ1qOR7si/vVBukwaTq905XPwr+hoX3YJJMqTimGVMUpy4+bhEXB8rgbmu
20viB5ZnMZZoGM903d70K3bJgk1h5Uio8NzVdkp+w85Bzc0N2mcQcejwrKZ/snNX
wv5Nf77vaAM+f3k/c2XQKaeN6uRZL7aOH6/vnWGOwPdKqS+kBzRHy2qbwKsKQMpb
uQgYccTwHEdtqv1JIU+Kr4HhSm4/hhkm0KMUxsnHWNhyCIrSJcIGxmjqDXR9iuCY
phOAzWSsT/3qDZySgooplfpCfFUcJxCceOTWL8HVk0gYnQm25q/XXkdWcwca2rBl
7bPRlBaLRwazjOsbFPxBlllLswZdon1NRfVHAT2FNJb9ukFVRhahXSP2tOtMUsQn
AMhYp2u2GWA4/seBStZdO7z1/i/2mn81cVcILm8eC5wSJo4LRYfN71vgtrMXasvg
jWSlAIZ/UbZk4idwE8VMRm/P+3cO+lE3y9wJrLXlnTZ0eFavUx7b+wWBxLLC2loN
DaBlBOE0k2M+VBRziwKGVbpy8KdVFoBRr4tX26AFZHpInkh1msBWVDKbrw4ts4+V
W27ObtdUnH7oNdJ6fUAD/Ot4PRjFkSRZfiE9pejIry9xhmVu9suDQlJuWXosl55b
UztTf8Nj14zwi0ANiSf/IWVRAkN0N0IIunE5lWE5TkTS7WtTrXGbtmjpp8t6SPvN
WYDWsmm5qZ2rudAm2EBAYUA62EG6McfU+PQK6WP6WIwpY4LQqFc5uWtutIbVIzRV
yCEU5G15C/+ipIL5Y+KbtTtfz22pxLBLmOn94cIbKeWqAzBj0/CQnxhgZ++lpxCA
lddUZsg3tnP09DgFHSTXdMkswmnBeh3ZdCCTwE7zhNokLfFnjkvBEWw7Ym6UwT7s
+SMF6q/ORY0laXUuc7qwE4KfOHskvhkomIQobPoG4auZ34/3DZ2IBGSHm2WJNEHC
CChIHOvM0cHK6wq9H51Qv02SbjjUyHbR29JUeMTlTTWsucwUB12f2nYkMglGrAir
fWMeUFMLdqop7KKfxA2SsNdekrznj3NeRXL6Tp4st2WgdEmVBKrAH3Olx+TD8Plt
6iHpjCKo44oR9zUkFBO41Lrg8YJcXBZ0+IdTUuZ+6qNUTLrsPYXTF4xphJDlj1Fu
L8Fq4BQh/kdwiq04P3mAW8/IlROWUYJ9qolaKX5dPOXtQfTfENMJNSnN7rIMtFMC
KA9rNQL5ju92F55ryeIkFIOaVSFC0w53mszqwmcORDT4PVY01V6MOnbS6UyqunCj
uKMr2uVGCUiAnOr0viEwnrr3aJQyK6Zpkc/Kt/pZms/DkTHsrASEhIl4r8zG9+Ul
GNaGEQKpzURZT+VtxYnEmvum3XddW72I0CByuE5kOYzvTdmOb3Bdo8IDMUjPHATb
YCdGbKns2KAwHELXl1a60WGdr0kQDbrWrTosokSIFI+Lar0f8e7Ikr9T9VYtTfWj
TfCEHYN+g4pRJJ597BrPy/hVfJUOyLn1qmJbdaFHjK++3u8M9VJ7P6t8PnbUHhbm
kF1NuS7ewK8guAwVKfYrX4kxTXTtpsCdrI4yXdw1J1lRplG+dYGy/ea1IvjTw954
SeBZsROZfj0Wi/WhnfywHcRv1nC15SOw6w3gaTu/R5k7mRJV93mQ+JGmpE5a4EaN
yCpndCQoeNxZieAqBZAFZdJ3Fx8efPUFmGqBLytlkwWi7iYotHQ2MLp5PnJGnEKE
wozj6VEiAO1I9INCHbVqYNIlAnssxcMmzRvbvRbZzmHXhhxA0N+AsJJzQSoz0XpX
Oj4o5pcYJq1x3a9YpKynvSSSlGGJEvEYHyoTUa1JNOFCdXppjh8+cIcQMAgweeyG
o0MmI/rm7+m7KbACBjMumGBX5/OUZUrZ7MamLp+WZOHTQV0yZtQ7F8nSwWDJrEG3
EQZbDw2FeH+xEhsPWqxwLFinuqZE9fO3IjLmjPRxISKNKzflWiMjCIZe/MNQr/Eh
XsblFQfLFKDK7MB0ehcMC1Rv1KmwN6lkep3gGJ9BeaThEVQFLc+3FqmXN5Wb+jiX
umox21IblEQHs31MS1pLniEit6cLC+1yXyfFIUoXWs0nhTnMWpt0kG8JsI0SuzYC
wMeBD7RoGP/51K1uSJjtjwOEJL9E+Mc281QKo5RDYgLAXDyMgMVSx92chlUnW5q1
8LZ8xYTZhVyu1hBhYASRrs5yYX9ChFHef8W51gysYo03VWz4qigpt5Bo7yHTXlJ2
4/71AMBSuj/Qae+J29fZEQd9HpZ0pmuhoB/6X//DhoKYP2nIx7JtEdkD4v+1wFLR
A1q6FASlhykW2x77moAgSSsCQFm4O/U//FgoBvbhcXS1pb+CipuNCMTbD8Id6IRh
5gd9lYSRH4YGZJEencqR+OJzf8Blwn+rQvL3H/iB+VvnIdI9REHp4z4mV1knq1rg
T3VuZSiTZlzwSkjpenbwRNrWX12GugzP0y9lYAz0GkeS36JaefD8+8RcuPrcuB2i
gq2uDKTseq4LiwqDytgr/JD65Xe1xA5Ehvs/LCrkt43g8DXuuW0QQ73yj2AKfYhd
/akgSg5khTgQ0KcBWSnw6jm+HnCmY3CuTGkjVg+hrv3xNr29xn8ac981Ek8cjiEs
+B+B+/gb551fRE0o7KNLNXJ+lc5YTGLeupq4nFkb7bCZ2eXH4T1fZ02BSFtMbgcv
nyDiEYpx2N5WXD5FCL6g4h8pkrsZFK1qS0VqfNQZq5+YqXgYZVBh23YJKYzoDE7e
usbTAtRAukdqA82SIf33D/MCUOj2/DFYZ1EwDIEXu35QwktfG1td8l/yEEFS1X6V
MdtP03Wi159v28SWhh5C44fleExvxeuMBAKqicMY8iVJSEd7HUcwZy8pbLXwfIfD
BH/jZhEGNz536QOLYu/c/hyVw1vydxnrASfl5BlXH8Egmcd5J/8UonWb+7Ut1BE9
Tq6KZxP2agNvEvYGVytd3pXutNQQWqHzZJHOHMFTAUbDPCNszTBrLp3uxQSF6YAl
Q1t69N7w3oBF+IDpWjCywCNLeYJs+3yW0zF7YGW2L0owv7uI0Ydz3aai+icBE1D4
chhSPkhgoFeC0D3gQqDw10AbggLe9xfl+uLkacwEyYOQMq6UtnQdLnhYx2C4TNLK
c+2K7JKctO8uVfYwpo74/1qZxLUr2qOLNy0UsKRuok/mvQ4sYcVWd+8nAFwl5W8n
9HQL06OqYztcvRqLqWfdaQF2IMxSE5TfD2sjQYG7+WoabOeyd15mtBkkyqmqSaSa
pt0zI/4IJffVQOonVXwHd1QDr4DHAp326+fkjLx868swPILPdPawxgZ3GUztG1aQ
77Kc2ybH565oSg7rDKtqv3EzNcgpGZA2KM5mNamPQBneZOZwaPuARi9R5ScOgVlm
gsVsKlXwlBVcEEDFUmo2iTDcdwure5nfzZy8wMAFlqTQFV3qVs5zMNn0dHegkGbO
20kW3iis86swuI9uxmsOMUu2nhqhDcD2h1969aJBAhhxDjrbDp13oyihVdcxuOpO
z3tk7ogdNqcfWYwkDlBgyv51TVb1k5l/QNN1SM0D7Bu4MwQ91msDy+/VcV6VHac3
3ERhIP3kptZk7OjNMA/AQ0ski125y2eCgRD4V3b+xQxhTpMHPxhHz+dpVURGuScP
yC+4WQrv+7axSkQVR5NVwVh70UtCFGwXKZsS0Jj1bggVcnPz0lgIWrSUXLAYhl/V
QorsWz2+LiBf4I/PkgV3Zh7POzeAsj+vXi3mIfOFS994QRzGbVYkBmeV2pr3aJCG
a+C/cZRsgkexzmrTxBa483n0tigSEUlHhhZ42vhUANdu74twlpSJG1Pg+MbOxFct
wP1Q+1c1/yBBYtw/LAAjDuYYHcbb+TaDzfqIxh41k5YAezQma6vRb8AAX5IWzx8m
u6K7lWUIiSFp/uwq9oC9goo7/W7ktkGE6x4M+M/xMMrDdEDbaD9F2R1iVDn+Xl1t
6BT2JS3S/6Mm7Dg/Kt7c5oGqgieXFgpNhzhIkBsh8ZkKDKKhf2z3fzTLOoPpvMG6
SOhkrEFHpXNmOqNG8cYy46M+I/uQNW2DJJOhkskVsQUvgExJF4KuAsvKNU/hId5L
iDC05Ado5MFJ6jSZ9fyuyVNVIc49iMuHOb0F7RBmPy9meHg/YHFtxsMrno+NOzD6
KJoTqtqJGLC7pugZdPWRNRGF4qI0qGK9+qv9x+/q8r5fs6Y2gEFLIIFlOxIKY5Y1
ZhR4k+etNLhsU3tbM+CRGbEb4UzZmL24JUbRqyM3lbicBavSanV3Gn4JZUe0flFH
Gw9te1W/OP0++xEvj76ZO9MdLwpTZUd00FBaTuNjn0PCn596FUB9iLX7UsOgLBhG
n4+9AkA2OJnaHJUOd8xjrm/WsuMA4eIHrytDN4OWIem96CiwuAq8GnaR6GvREXbv
FTktDdDqw/6UogA5r6oUFXbraEtyxQdfd4W2xuV1Jjm6GSHQfJzAbHGqNPmFNv9F
1RMtwfEKDpWfvIlw1bke2GfjtAouNuNA6FmzT7wmvYqb3A/3B7m34qA1qsorejqp
OGQmemQv8tqm66skKTBI8oh+wTp2WByEQIxq0KJqAFH2/VcpaOqRru1I3fR/6g+0
QetRRJ26vRlf5Pb4ThG4nExmtBQr+ljrAar+m61S2wFuGQYrCbuAWtceIlp6mFa7
6WQ2jNNKnLJzOkI+MwE9ITusWq04mEs6rW1pvm/lnXOY6IrGtHbYHHG9ThUACtri
FbewZdXneSmovKr8fO4Yqv+A+wNuysm8bZIzWcyty2CMWaCUSgM6hHwWeZsDjl8L
NvIcc2RBc2o1kQhUdPHDlIKfqh9ShmsPwhHWNFkF4P2XDL1UuJ4QiZ+7sT5J1++T
q+9F57AMmPLW1BgUz2nspQXfn80M22ZcKBYpt6bbhNeJYwKv04+JpYWYsx+ZMgty
29fQq15bF58/0qYXa/kRf42Y8Nbj1hdMw9ALgwR67kk/s48raz2P1ifgxasN1i03
A35dnyvfO3a7BdU8ipvSXEetbqKq/xzep/YXyMLFCM+i8ln7YxU6IwSTpDEDi+gl
QWkA2nesMybW4d1M8IaRH5MXJtnTs72V2pf9GPm74ZtGfRWgkIdC0QZjLWOiR/Gi
qX54BFx1GJjyvWLQcFLDR8a8nr5KFIlQi1xvf/SsDn02vCJg1YBlHp18Jya55tQu
aOLhbE8+GicUL9zFLGmDIXBI98V8K+/L7vEHX+QXlm4RQ05ZFiWaxNS5JlPSay8S
7j+nHwWKyzU/ZrbXwcr27D2kmt6hbFUPrCWm+ARYXN5P57ql7vQyw8n6JdLGB6Pr
86uueV/BbZHnLLl5XIhfSFhctUeeaF6GC7zzkEz568jtLJcXpRJNHWUcLFXKoXN1
FLVSPbKlWbExHT08qCokp9rNL2A9OMNmCkGOY4mNIycNVqvXsGWLPGraOt97YL7P
2qmaOQpHUgsS5KHQRUfnxu5l7cnmzBibGyXyeCSlI6ZhSzzR3w1fzOZeNLltr422
c/tI4M7UD6pC6io5PBKMxYyloC1BMm9XGLx+1gyZmMtJjYMrcnUofAbOyyowmmOD
f4R8JaHaxfmDp4UJw9IjJ+bAtElMuv27E8nXINDSdbrVl5Fp/aIr1271DB2Zesxd
okr6UhOJQMCOSK3R2dPyzVjaj0M5nmMucKlIHIvXC5XIp5wsAakMQggyylFeAErA
I2JqNgBiKTcHAe0Hyd+BZGtJYLlICKune99g5iXyUdeEtNTgtYeHcpoU8RLBd1zc
SHx4q52YZGR4H8Zz2EZ16P7vjTLqA+CU7+u31ji+gLUqJN07wBlKK382K+pxKyd4
DvZzCQWIzqBYNTlkN4itvaKW4Rlh08oQN5+8iv+tVKkPDjl/00j9loPYQEHkwWo2
UX0I7YKWTEUgXw+v8y/749qBumkgKlFZj/ohW9JQtIuHNA6WdsM8Mzn3Y73C02+r
EXNm5ESILpwTa+YDd7y9ssb83kT8Lr/QPNedHlihLz6oMl/BKLkWmD28uP5RA0dR
8pk6i/mn5vZBR5nnb9NxLV6figOMPE0bqJ8B86lqJfUwPr3JFhYUoYwrHdjZbCY8
yws+UiWMSEKVj84TcbUzS+xpcZlKFYhPJbDw4x8kupFZuvQgg4qeXX+1pYG2VWux
39tmOxmD+/UTUUmiV94mGdRlrLrrEW5k6Rdn2G4TyrCx+JFhFxH9f1h7EF972JgZ
Xks2aeGcX1wf4An45Kd6VS6APRBNn4z7gPEyH07HyJ6j0ghWLMyEdJwO4J3KlsZN
O4+EWzPdA+JCOaJD1rUK1YajD2c1DmtpMKS7h0WChzVYvB9LR/teigpGnFzWp4q1
ELBZKEaxlP+a1VNDIxWjrV6NY2V3cAYi7nzHRK5Kc12B68k6S/rgw4ky14ZzdVg8
6WPxZ3qeHk4O5qsWKNUTE0WKmKAU6crNcY3cjvU8P/W6R/XzG7ijGoPhdftIHAKD
IztqMm2JPfnoa2JBV+nlyd2kCxMoQ7GSLGzR/S3dfAhi6JlxvTcfN27iFA3+4rW+
yy6fa1eotWi3xIdrLvXiH7aRhQGXzmerrL242HXbK9CJ3o0vB2vkRlOGBKrQEUyQ
1VABKe0cWsU4Wp17jHWBhEPrl9dvMzZ8fEUGZA91w+2Z1sOjxUdXrQOHn7MqJRc8
ni842gwzgjJgkiWoVRorKph9hqg1pEppLwHa163VpBE3GyTdM77/uRtyMP97Yj9T
aull7OMIxZ+Bg5ZT37NZ8vgl0Zcv6Ukj8Yan4nVV1V6e0HWiWyfe3orALjmqKyV1
4ABccg0T/+c5LpulsepCezw3+erE+kEdVUofwnVWopifUG5XZNd+z0ksiBuQXudy
QP0W/cf39ZhT7KHAtckCfBv2c6GxM1hd8wBZ7Z48t/3xzRV9+5kIKKIQWThP0kDE
w3EcobeDpIRN4EYlppA4jKyFe2hsYZn2avY7J38ChNpl5lBbaymg6Z2fxa5wgh2d
dFaP01VM7utb1fh4PGdlahZc1Mz1zik0YrJYGeu4RoGOc6CdAqFRdLZ4CrXQ3cr7
aGsbw7bS/nzuw9WZRtk824laKQ/9v4KuN7R7B6KAOdoDPiB+B7NyJP7oWEsqcqei
C8pVDTOQSrDt4a89Y3xdaUNa7EIIwxHQOMhiBVwyND8hXSANJGd/W4aAIr8tr/Mh
xHuhxqfE1WsHw9XT7TZEbl+2Dd/90uJGYiyvdg9O+4ZNv7EPmVIKlnYojW8syCCD
q93Nox92nbyALGx4HTioCzZXmS0hFeZjwn2D24Kl7AGbSSEf983ARsuS4eZSaw4k
dZ1xx1p9BIj09B6Gxegz6w72VlCi5QXjmi5HqgCnoM0YPiEO0T8H+UGv0YhLk9jN
mzckbufH8leBQ8Z5Kct3uLw7RoLSf/upbduDaZMHeEln4ovanaJo7GruDR0hfaZl
ksZMmbvgS8yw1QGzh7wCI2pLGBC5HQTSVi9+4d/XZO3mBKfRIak21eK52048K1/K
H9jcgbifY6Ki+TjHlEnOL2KkfZPb9x+U+1uuch5DwaAzEBD/OBfWC4S2wmOIQ5OL
lJOG0CtLg8spksS2sMpfDC7kksTCGB2p9uwQRGiUBG8enKFUgB9HpZpaQoNkm8VT
T0nyYRutJtQTukd+BMOmwbPQ9i0+9R+0nllb+0ymf+75aIn74yUzfB76W5d8fag7
tTqKphOVfgt6Abh+UtpphGHCQMkSNxS25Nrfu7Hltl+4H5C8bJojwJyWNiHHU4/x
ynlcTCJqKRUy/rUGasJi/ByZgxMqE2No43wp/pm375LnAGb6KRFEsQe5JKq+O8Xb
OOpL1wi5sCm12m0wOZXJOSVX2cq4XnQAbGdv/hvE0i3+bgtfYCpUTcGHoj6oxEBg
T4akYxpwttXNR57+1ZgTaze9afQASWhp6alvMGu4pSwIRwfUwSuh9x3yb9TtqF1+
MDo1s04D66wufMe2Y0ud34/im6hWFFhBITQf5G0Uep52ofcBRcE86GL72qk9yg7z
Y+lM4OedZqsULp9n2dGf3PrzcVJIqNJLapza/y4GZMsweeUUTf91jug/K+CsMa7W
fByBXZgXY68udn4ZZyQSuCvkZz+BVOLaQmz1J/YxfFEST4th15oaC6089o2BTRQ/
phOpoUdNoa2oU1+7KhmET8x0o6o0qjwWRLuYQxN2gDfru8/3SJ/f22nQAtH0yVAW
TECOrzJUZzN8QtaeRdyohJEvi5SBTHdi0fEY/htf4d56D8XnEiVrShltwz4sVwwh
Xo/Iwld5w70d+0+7l1KxzczgZuvSSz4ybnd9hbfzlOG+ChalphJtXhQxsQ50iR+8
UHoo4xG/Oywlgpq/kalqsNtf1UXwqdY4dXl4Qnx+bzi/hd99GOyE+ydfyRZb0O9N
9lWr23MWB6V7WxZztx8iBu7DUFmyQa9LWZUEdRJ4T4T67A5tH4Tp5h5U+2IHJ09N
iHvOspTqCh76QFrHAkV9PkF0LW0meyo1vq4R0InJ1Oef94gEVKhQ8OWSwZA2tnyI
Wyc1Jk58MLBQB6YtS2dI3yy+ELpatZLsCUDq8ArirOmjyy3dQx3X+iXMRhzr/VVw
znoLpwZ5uqUlgml6EnFmUdr1iQ9RWTpH9nGszBp3HzwGz+sFdk+co2cA6iYt8mi4
QQD6IbpfTSvA9Y5l4KNREmwcu1eZDZPW9uKcsRbPFy5f68+Y77kvUivo0XaZXZ4C
jlvDtCKhknSm3uE51gdtn4+uyaHeICokGFn8KGnV8sm+aX5H/Iz097rOEKfaBwAP
aT6zkXSymv3OWDh9now7Ye0duzzmG6opWIKzV3Gy5SWS7h3h28Wv8jsVjVBtvXrd
K7PDawISKluf9M6qkqdDWzr5Sv+ow97C/vZeFAffeiu/9XrElld8YNAztQLgTWp7
mWVTd1xBL1M6Iu4L6Z1toXbkAOzyWqApxPi7NhoUYBZdlaT7Zre9dRBqXUVW3+2O
n0xD/9q8EsQzwJrlFT1+OTtleo3aO39jqoPcK2Sm/+n2fsgEIcwHqfGO0V/WTX7w
zMLbukPADLTq05+kNX1eSbkLHWNUe5UUD+ROK3ARhgNI0RU2IkOMucDoE/G80JLI
S+USD4YwFtpzNDkl1MHYggEdNjx+75G+l8wLmQPM3IUAV8aixsTAe9ZD4WYsol3s
xyZAGUiN4QWcyZxBWtNlVOdfaoXTasJy8Hdc2STVGqd/9ZQuGIF1lEX1eiiGeKMR
vBjM34X8B4hcAI6s0awWFJezB3SMC1PwUzQKC9z2oGgOgpR2KWa0WvvhbQnj9ACn
QUTud+HnDfEvHkAJdITVONCt+HKhJj5OLyamjH861C6dnsvPbTM6ZMy8vQXnnI0s
KjJ+ClG7amip5IRpJfRMG2yPg+BsyOxPRzK743/f5eaK0mCmyPvAFUh3+VIP3obk
ntaD8QrGGJezsnSLUA0dMYDwtnuDExAcw1MZF6g1R5Uu9xuh762nNi4R4Ji9LM/0
Za48iLU9H6iZw6OK3rfm58pyCGDWwt3Ks1LNetvDSVTG0dCYxgVna510qTv7jl8K
2IjTYqwHP+5U63K1kPvMToz+gfhOCmKKBEwVT2EDOWacarmEGsO8HcNdlxUNIjPH
1BZkWLXYyq56z4Nm6di+NbM/GyXpkEtCtoeaMDZNfTjSblQXS21CqueEILxklxAK
DrES8oiv4WW/vS9XzQyiBnjakmTr5nIhMOhuWc9MZr8aKhiCSqK4+sE9xhYyiXrh
9bdPYqvdswHTv4Facg6j6tFnsKvEItUbTGdofHNTglaaapec4ZaBrL+mvJasKtZl
ZiVqO1rkHCQJPvGHDEohPtvm7Dx+rztrQhsnm4rSHwS21vBPB5MqRTDG58ljq/go
8J0ff015yYKYPM8HPZ9L4+XdFDxinL9ZZLbba8pBmUVLO7mMZthBHHla8EY0TiZE
Gp4UgXVvrlPXdoRFnwSbE+7+5naxWHF/m9lGYNR5Lju4vaizQ8kPVTVLnLVJIJ2A
MgMh1UuB6F9SCczj4cPl75tRiwz2JFjjtSpojY2gd7BLIcYI9EFkah99ASN0mi+n
rOdlBos2L3rCu2JsbmrKbDxVvuleWU2ZweaoWXsctHnnWwYZDs2Jd0ubxvAYgyir
s0sI9mmPG40UwuKiAgDRYr0gm3EY0v+ITuN3VfD1tnD1L7J4Rg/ukBQvxtWsIoHN
RfbS5/0BOOFF4oUHzy+C9vi0pOECsMEEuFoutN/OaCAXqE6gus2og0yISnNbT0YY
sQYnglxWUHdpgAr3nn0NF3V1tGZfGtZDPlerMIsYJLORbWuIeAISakCmdHLdP5y0
BwKHnCFg8YBoCnofdwJW5sZGfVJ/ipoQCDXI5prR+A13HreN+Gh6LEGimiKbECav
KrVjVkdujzy8dZoDygzIIJF1aN2aEkJYDMOHN+/NXRUEcd6h5+7KmjxF90K4gbLn
zKNS2lvdXII/gzNdS67OhUo0urVz9wUNiEZ+3H4IM6Aeau4o6wv1GMLD+6j85SaH
jhord8g/rM4/95jHPRz/O5MXJIhbBMI2UGNEdKu6AuMr7yYPvTS+06PKTV1mxm8i
VO0WU/JTP+YsN0m0Lpiwn6cUxF55CRu/8wLhrxsKz2wXqKgjWKit6Se4/fvIp4+g
IFfcquHmgnYHYmdp+03RrMui5axlToDSEzMCclrzf8vBFiKrCQZ5vVH6u2MjW9rc
2pHeglqHKfOFAT8QRvRDrz9q+C3JRXykcP+JYx7VnIUN9hlDkwbotA3PgdkMpP8a
hmt4ZbDt5t7P03dSAM1gvEwud/tsM4aLOHrw95Li6KLJk1vsnXkUPGUdCtY7xYox
+TGLvBHt67bhPPgKcMqlLCjpopYobIjIA/JTq20ewdHr4IdJQdV9j/8s+tGuOrSU
s3cbDT3osltkjDBk5E743mEaQEkokv8qHjkk7ahGuNgoucZcAuTiah2LzMNA9DX1
xGqIR5IM+oFEXVSde1arViMMn62Ga+vxO/O+bjUcW1rDOkdfCIJF1Cr0c9de/n46
agpGLXJfJTnm3dxicObIqv4oPvuevQ3YTrvHcHUi04oFf4V1uWvqPNnPW8dO+jIg
Qg4iWJORzuLrXQ9n/SXTxXvyByHmQWqfRVqGzms9HNEMghuJvnKtA+WGLAnb0RxR
09Zvmdkdfu5LPg6xnP49aOa/GAROpEcOjyJH5TD123ykLQKlkOC5789gJJ25/Hga
ZReK0kszr+C8mFRprRddkYTtMegosqo2ok5N+o6nypZtQC7SYQs7+evnryG10uGk
QssLf9VWegQykTaEvwEKs22+Q97YBMSbvajQxzyO9VD6sPnRqbQGqn/1MbxkHiSs
3AhaiOu45uMPpF1IlQfdDEYIintRZfJEgAIDOz9wZMEKjJ0kCHgb+VW5P4vMxjcm
6+gbtjB2BIDlpW4a7Icq+7QsDwywiJEO9sHgiO03E/WS3lxhkC8pwfo26O982G3j
aQNofcZ1WaHVmyZzKqYDCa9sCpo40AJDja3S2UqmjpfUG414Wbr6T+cl0OecbW4x
C8iykO/SBuzalPmZVBtxOyzvPj+8aR066LMOHURfjjbaTGNOoVQgmX1RA4giLbO3
ALhBKfS4J9ibBj5YIl8WRvlzdD9HHqMuLtAlVnENCnfg9XN6eGkxaD9ATOsgFVMF
VZQXCvPK24A6kjRoVN/RJNCpp0eimiMBjFxO+oCKIw+Xe7TuYjVrLlBVZdFoPkRV
G+cIOZqstZKDNy1WJ8OmtZxlU3vTZygA64aAkuimfvtn+Ze8XBW7zMeNvehMu5lD
zHcnY6fZoEZWg5MPILHJxGCgES3nWCKniac7Jvp1X7WqW9xvK0Lwas0YkYl57ivI
HiBFfAiTLwKozQD+m2mSbNFk/AAqMemNpJnutuIyKnktF7YvU08F74YbjVK0T2vP
14fBVDXxPEMnrNWQzfOxnMAW1xv5X7X0ma1jeXTY0aDeuqwEJPCqIXMEbTc84rS0
Jn2ugiGgk5fqll8HWNFDFgCvkEq6XPOC16VePZZpfwr5mBxycqxua2ucpr3ffX/Z
4MYfEdVNiLhS2begdURfNo9/ZlyGXvh81YLo59fqDDFAb2DtR5bZ5L3oysxeX8vk
AaM0EpIpHHGNc4hQ/YZE4PllBdkP1lX7IIX6KmiHUNpQHLcbg9C1WDTnfX+3x39z
CYqu58hO39mqGeR1skSDbmt8fgh2Ku3rLuj9AacRwYwZFyyO1G27lkpEGG4YAmLe
1MPcEGew0QBNAzQuPUJusy1OJNsN6rh8gcjxpgEI5sQIn/jcRdgn7e+cpr/fIg68
5+wXpyouiHLLvJXjlrLYrYJPfXe48QmMq3kaEL0kHeZKFRjjCgZhU6foYb+u5izX
ZaucWbfeF6t85enln5LzEn00nX8Doj2+jnUmZV7j/z8d9ObOVtqtF0zNwS4fJd8e
eNg5HyC7NmQy7eV6INWEeCrEwtXYSOJTDCGyva54uBsxU81tSnFXAbW5DnwRPtuT
BBhMpfRkLuKGa6UCLLx4iwt50VeglWM3Yf8L1FS7TnAHDUnkTRQGOG5qvDI1VB1e
yN88i0T02XNXswxo7a6B5/M47wL1P5yFq85iW7RXEB5t7ohqtFPtSqm1oB9Li8aS
TEnhHvJep/AgIIvPg/gH/Jmf4XrPYYTOVCb0D9F37grk33mzasAopayIHnSnA/fg
Kx2mng+UYBeqL/e9GpawyKKQY0Qi24mp0XIZXU/8bNoTbj6X1EnW9c27k+xq0Jtd
qbP5ombKQ89YhGwZL0qkPwlPPy+CYDf1UH2Vfzb1xPrs1Xxcs906clvjYZqFcV5b
at3WAld49oWq9XQwX8juf23iLYgEkbsIJhfuqf5yvQnYuHZpxwYapFOjuFM2LGlt
fP+S3ki3nZSiZzBR7JOTJ7BC998CLx9SM3IoLdnIQ00Zs+G1pxvvl03DEJkZx2ff
R9B33Okpa7ghbj3wmKwYzs7gOwYLxSytpS1/cLWlTK+ZaE3qh1nZB4ndpVqAMmGw
yzcaqUN23TAyPqU42F8Y2aiU87CH7MbhC8jRNmeb5jhoCfLON7NJlj2Cv3bsMeHU
pdx59V6bhWjSUWa0Wg7r1BDx17ndQZcfIZnPOtw0Ekw2KyWNZMrJp7Z94Y6TP18g
r0HV9jKCAkggx9zN7WAY5z07z8LFleAciAiIjxJvmt/mTCAXqO5ow/G7+wZT0dR0
pGbcY2YCMK+nFvVH3MqAMhAGwXZziXpUmIA/8g043shryBdzFssfT4Q0YQGGIb/E
EluxXx/iUq13kvA1VYLM3G9SKZDT2YMZCOENxaXH70RiPpzMeGNsKR+9xVRG+QDc
h72nLMUNeyJrxz+h9S8UC61b9wORnTRC2PqHr7YoPXUn4D3z5wvR3hIkFsJICSpD
360+UE+rkem2UytwrmNkR+9iDohYZhwdJs8U8gPQEe1VCeULzY35UknDDfldVPb8
uChBUKtj5FjZVhYF7ZY5fW8AJVRE/u5R1L4vN0nFQRuVeGtfedcbIIcTOu2NVyNe
1R4smgF6mtP/VJO8pj+SL7JT58sDtXDql0hXm0FVB0w/Jv05CVhnvNy2qmHqIQdS
30ARssAvU2tej2FggNj3QbGgLhhbyYvX9Nq2AfU9fxOY1RGyV5q4yBTTHGZOkhV6
WWbmYINEPjJ3CrquauCNOuDUtcNYLiT7OP23ki3aOhKZ9B7+RMlDiq+jUNDiAS39
3oUs4eZHm3RSlPXibnFFl9rfBXSkqqvpXZj4Ci61icVL/L3BVd1oGZNemOhgGuma
9aq6EHaE/Xgv+4AP+5F6r7K2vXPBNunQkkVaZF9FWLgSPD7AkeQCaS/RsV+E1bWF
o46/LNukdJb9qMerRA26zEZNZOVrZouFPhQKLh2hmS/zqGBafe86e3sTEcOnVFBj
h8nNgs87y/N4cOsmkeZTHNqFkFHIyh4Qe3fp74HXrcNKacYdi6lMHBe0LwHycGQ0
/D0Vkoi6uTQbjckR0nIqXdlVLNd19184HzX0UdyT1ydIBjWV0wdapLnCNJ2bU1iQ
FLN15r3Bj80ebZDJHfv2Ov6qldkqNO9XJx2EBb40ylHtdwSh9Lvot/+spPhLpi81
awDW31xJ3s1O7Z+4yMkrNtd+CVdAE9QQsDNubivde/R1f6y+gtyPLPazf1s+UYTM
uAjKnvxP/BjSday35FiPT/bVZSxes86ehe/9SQMeQiK0VUNDI87TlYJAjAlkLcHL
ckHlUHJVh8TwaZSB9U5U5yrRNHfwN4YyWKVyWVpEZddW/wPZ8C9BpPhnDEbNHWop
gmY+WWpjG8+nds7G4iWtFZUTSIpvWWHERVNKUuUWM1nFVmBwA+4y9QIwqm4QyvpW
SQG8tcJo12E2idPu+qxtg+vl6B/VMrMp+oqNocTHoR5/byU9/bz8u3G/Yd/LhTOH
+LKcDYQ0iNwk3NrbooiM6w9C560DQYTGRIoSt/MC10fmfdmBs+jQicpJua2NtzVy
l8zb6eGnCR4U3Ll4pe9X4LWBHHfeoU1kaowZa/stUgp9QopXSjY7CpwpPNpRbNpQ
qWCc5w7yd+xZks8hL6BsfN2ULj9k89KJfZkt4FGFKCQiEyqXFbgQmT5BHA8VOMl2
oSBpbCc2eAPcAlJbh9ejZB6dBY5Mwfh+rCg7Q2mfU1ojCkE86kKTK8Az1Avnykpw
/OCrfdBPT1lt9pYBwUmLf56G9QmNFPIqG8H8pIUsf06RdSIGxLnhzaai6DJnnAFu
On5q37ex+4SBscbqVEp20bm0p0IVB5OrZl0eKVgM5nYNKwf4mzot8Gxx06ls61aH
pw2sWImYAmD50IyZbF4WcNHDQHhMAEW2e2hSAAYVKcE9JvKyucjPeAGD7/DYYkZv
dMxIJ8eEoOYEsdH6A5OC9PIcWhmUc9nrSBhQAg3FhzpWUoK6As/43bftFmRmXap2
LaXB+lPNuRIe/JLaUy76qUCfEgEmKj3AqTHwUtVkKJeht1YXC4MsnbtPkrzuQoXU
mobjHFnbC2yhEhHAcocaF3glMpSMDXPr3cBoxZ6uH2b75B6AGCNzKlKZn5E1cuJY
Py9jyP90z5hLS+VnaH5My7wFVf6jh3UrFTE5oSyRTtRTyyDN+y+oRQx11et9+c3Y
uflGphxQDIk3Rs+RoUBEzkz/gqKdxc++PF9vQpJ2gIazF6kaHJbw/ghoJs96EerM
2Cq0KdEO8CAqmtoO1Z2NODMQ5FV/B+mTrpV4OZsNndGhGqZexYM+QcYMOgdDlvOt
YuGKs7iFc2sRdv82wCl2UDZrsnJ8WOMwmMumCbB/sY8ld0Tv2v81Dq1IJrOJJ0fh
jt4ioGt3bIs91BzDok98fxB7fFJpfQYFVQ6PkS9cqbTFMctA20uR12IexNdUAcMo
kxHESpyl00QfuxMXEt2V8yGT48K3S6IRn9dKsboaxqLBD1MOd7YJcB/cq+3gSLxy
wsw35CPx8eA4n8tK4YT0x3bywchNx8uX9+7K1LHjNgb6xr9fcE8koQId8BoKW54/
yqK0LPqGBi+YMxPh3PHNncSNvOMnxs9qtHQIYqViwdAavqXC4Ds0K6dFxO3p/UAa
0ybEX0W1SSl1P9DDfeFX8w8qim+yDQsSSeASIfYQNf+3plKtur/Te5eAJlIEgEuE
BhLQzS4yK3gGabTj03AOAiMSYmpOz8qhCuypPHYjxed1mgn2zK2NgqLIx4xTAEb9
J/DW2UUkXlNcYd1ifEwhUAWe3NyYhvwnoIoRp9THxb+5/BjbCcBTe6u7+Cv0AJH3
bEXziyYGbCVg1v6mGNAJHoGCgHay8j1qLUyGeISTj6DgXsqCqu7h7NpMQs6Xtgym
SOZ/+aauxWUYLHNUYeUSCwrfiL2lxs21dxiT9/LhnBXRH8uEJvDE+DgjiUIMGTii
qR/9zEOzwuc5QNEyhaiZIJdbFsixmv92opV8JZXEFZ890D4r/8DrjbDJ0ipbyuve
CIMnNy2f3L4Acf3PpahqbMXwIATArPfG9z0lQNQplvJYllL8k3mioxiXfMaWHf46
E+Ses2MwMi5rpMdxirfHA1t8R85NDVwR+PxS1Vwz2ozlwk/bwbxC1JZDgaU1Kox7
rt/v8eIhia6LZUAC6ue8h2KPPJPuhGy3i/v2TJfXZ7syrw/QcgtN66AsgfFDd+P/
MHfftHyyJ1fAYc/z4Z5RoEt4L7qbGksOZAiKQEZCOM9QTaFaq1h5CPInGMHk01Y0
3Gu3xau5ep43cEyzZwvAi9jAa884bez10VP3bXk4iNuRV5+kgfViKsjfCKnYBnJZ
M3JAGWvwWGQ4ratf7/zPIK4EupygUG9E6bSPCLq4UpPQL4btTFBRMO7D+zFbslb0
4zdXJFu3zl6FE2pIJErVDcISQc+zZmQF6sjhgONHNCNq6sJoSrImHssixZR+0j2z
3TvdJGxiSIrWSMxftzzwiBCH6N4cGPBcnnvhqi0srdQQMG+l8lmFZ3f8Zr6ebTdZ
FIo97ODl4R0iOBzxKhxa1yI+nDSZ8MyfF5o9mUYGsrMUFHEmAxj5gdvvOTqtUQTM
ihjLJ0+qBRUQPMhzUhr5ZJErM/7nm7K/r65j7DzD3YKbRIdqCfqSk7nHOuk/plrs
r45cSKXF0dGwCNikaRtqyis7uLKgCxPAQtfueazjzDOJEE6OGzbIqc6n7PYj/KGY
NY83goLgymjn3eVlxW0hW4I98GUKxlqswl7PNikYPbAW+2TU+rEP75StG47+JQtD
p8koIIa+cy3nr7QXyFI6t2DxXxahqLefdXuEZ5Aszse/Fr3/XXlc1OUjyP6E/3JW
kQlHZitYhu2FRY2LD09NhuVkp5VB7ubkR+o84WT7gSWQYthzOfQPvSUvPyrrbzGo
asr3gCwFufZ4ZMgJmK2VSzYL0svCJqUPuZwy+d5LK8EtnOIPoQfvKt09iVcQkkn4
PJMm6qGAwmFsdA3fhwh60sKn4fIQeQ71RJGoEttPLelKwmN3FIYdOKi+6utzVkbP
dXqfOKujrZP5h5DDU+dnYoJHyPWmXSBgLudDKoJqdSHNLKenOaot08lwOPu5tzP3
ydmnNVXSjF12RtBoexpdXAeeMULl469Xw7H8UQYEJCWIkpc5aKmD46TfQZUDeHMS
un4XYD2yHEoXBrtm/zAqA4hlxN2acoLKWTqI2H0wPRfYXsV4th6FHC35wkWTOq89
RyXh9pjMZ0/j7b052/Us/6jjlK5y2/iHxbjCLESNueaKdI3NB5nbb85oaIAJq3lb
0gEfTAKW9h+ou6z609Hp8k6lykQmw9oNTt7oObwSTs9aFD01dOYEFv3qrzqSVGby
FdRrcyWPsdWORRI9KuYgTHKKbFybGeSJek232ykpyjCFhkRAulKDhn25lcs4QKe1
g4ZH2A97VybE2XApuxx9W8dDZULjw2eLHBjZVG4BmK9mtF2o1GuTADPoFpVOipHy
I51+RYqthEKw7bDh/kj62vOCoiv/b5rRmWhnrqMESS8pt315bpGafUul6Y8eRrDN
iULl2ammEiqpE9WeFd7g7epnxHZkZ80hNWFg952ng2SmjDy2lO74fkL2KYb0xhFY
/ESOYWgp8GeSjjep0bUFvkqBcGBT07ExPt1F/JNH8o0WqHnjqG2CvIXOmoNIPV8K
0HTStjcs6S91FEVCfVe/GBz7vkqrQuausNhLHbrlznnxMXvoJkZSdV0BIkwteX6M
3yhtaRgIGXaxPHgq2UXB+40Uywpeuy1s+NrSgOFSL6cUr0EBrY26xraPD8SJ/ULI
RnW8VWp2quc6W4lLH5iNpp5c+GpvILTmMTr0/kuZKb9iCUH/mRjXvywkbxvNOkS+
9LbxjJMCXtnwlP3Db316mjC1xN+oQFPhGeefNzr/PsZdG6qDnZLTLacIMd/Lu3Vq
z8TmREO6t83sEBEmXEC8uuWg+///l/AwY17WxO86GbXYYw0UH8Ym/zMtGkCWdZc0
Uvbay6i8bpfbeQ7DxuTAPpgML+b6haJ0HYO4fQuQwm8w8Z8st8GDmFQVhWp7/6cS
JiaphiZ0ZDOrZjsK0aZB8sHMBwJ6++bd1cUkHfBQL35PeDBVNJ904QIy9UwRB7hy
YExLVbKVmxBVPvhigMHOG2l7qup5WyE3OqBdtZxNBkqn3N9690E0DKK/9zfWShmi
Na0Dc1+TMkCOBxsSgXZN5vnmIScrznV8kGwG3du35y1gLmEYYx21L7jgFyNApLCa
H9fkpyzDMXn7gYsUz3DQSDfTZ6xRPZrsKsWoItfxXVYVTEKtBfSLAJk0gIR6YPNt
iCZu4C1YYCi6f60NtJHKy3ArmDJKIENF4HFrisD97e6qBalY8FUzEQVsrqDYimIP
KMgh4DTGgWi25WRZy3au8CRcgRBspHsnXZX2HYn5Ws+0Mfirxy4cRL0FlxTF8/sP
RuOrB5DKpVQi+Pk98TgqwqNM7rqf/Gd9heSwKPlgQN1YucDGyQptYoHlGAlrGk0D
6ont8Xf6sj1LZ+PwtyLRKLMygrW7vBkz4czTigvpgUQgKidHb+uNxObBHTcrR8Us
k2nTW39gD5MgT4k/+CIrHQSd8syVwcHb2f3bKBSJPBI4msPWGWtM9yhj9Zb9A07A
3EH7LqwfA+yjC0bKnq1zxH8Kmu4h490EbpMrIUozUqCeImsj32ft1ga6ngRFzBoK
M6pVImOLrh8PxziTUfB/EpIUOSp5cw740CbilZlapCgyM8Oe3BIRRnNcz227d8Qi
jZwgFD7SW7L88ES7hEO/ccUjnugYP2u0VvjxqZj4BcOHMwcTQQfh2sr5QZOPaVjA
KxpDbXClIZQQ8SxOEPRZxvkvRGUd+MyUtTgp0hCFdTkzTGirDlK9Rc6VOln4ec+C
58nSb9DNZcX3wyApdS4HqWAOCJjgBUXsZCAnY0wiaO9fVg5Nh40hH+JWnkB9s7lW
tgyGCwRAAtT+efWU1Adc4JS7YvdAabSljwtYPhu+X5LpJBKi0x3ikZkepgHsgOOh
rZGEWoJ6VSQeKqV3gcNGNFvNzQPxBU95lEW9wimXlcOqhQMpztep9VY9Lk6Q9/r2
tfZislgmNDdEcBrRzqkVw/5KaaPniRBAGlOHKH1Z+/dzsiu1g27f9g4jhPkJpk6J
hE3T90OQ4TlPSmoJFWtJvMtQFID3PwAEH/gR8nDfTCCoDthyapZW/zxPshk8WW54
4RnJ3wzFhGe8xgTuYfCcAEj+0lc1kEy+b5RxYQ/beARaHriGSNbhKlwmfBfJv3vD
5C+pP3ZG/3kVu5Rv9nMs9bfysfngRjQrLBW97RXBsgXYXaQZ3rzkJJuRveL5itiD
C8ImvMbCoieEtQDQFG70KpfhjoX86T8ih917p/9ufLji1KPBxU0DnLHdULB3fngL
iJLblnrRkC/h74nzGFLQJqX1MbR+Tn+tiHa0PuRKH7F5lX7kAKIapsR3N5vYgTMo
pdtdVf4de4IGvX21D0FoWl5npMgkz0I+cMS66pTEtckN7GTRFTAri5uIavkbyXk3
M3VXhujrWCbLPaDZ3E9OZe9W3SsNVpSfR2cEju1Has5XElRhIzQl9TDI8BhzXJP0
revH451wAeh12ZffTDiv6bjHWNSFSBebl4ega4PZ63VpYPVtWgspnflMMa+YnM5z
eUhsxxXAZU96B5y4I39KMaMqd8NzWM2ebUH6X4CmbhJe73doDLeWCbO8uJSfMZFR
u/Vx1EPcpJ19Fjz0jICnanaXWshjEvZG0JDtz+lx2g4NI1na6GCCvzn0tAdA5478
dsdJsjZ29pzsfFk56baC3OHTL/xrYoGKptWIwMhibhT3Hb0r/mugt5YGeJ1lylZX
GBJouXiS9KBpSiMlrk1XX9Qv916kz4l3JbZJAuAgcUmbRBbVdRoPR06rWR7SITK1
fqX7ehPlC6CiWRDyu1b8AIbxhwuTf2o1+C7xbP8uT+1AMsV6rSQmBc51XkP5hXlF
nlHIXkkCCjHrcimsE/1v9KvmEgIZPb8rDCCEut+qlzSc5OVeARClDekV/gfAMpdI
aBJgj2EI29wyl5YumiHoPkrYKjJBYuif4Ns4dMxFez/EJ5unIITQj6i78nTT1Ogn
e/XPzWloFgZI5TGnluQyWIpI0kc7ldGkffvm8hbR6iuGuHv6WDO3qKCchWxc6f+u
XLhvWPtjQegxrTmneY+j0HWDzfjpAMiRIsMI215WjK29XBJdk0GqIqo5lS1mYHPn
JSWHgqU1gRG2vQxh1X1luq9OQUbwcrKrljeW1PeGIgJWIkBdh4nm6+sqrVrBjfAq
gn9/N9qhSAXq7uMqlKAlcewFFRL/pgCoz0c8HoNIfxRxgYHpWSD6XlOQAzUI40+X
y0iU4Ms8Pj//UPTuPxTry7+9f4B6TRki651JjMhIC3FnSkj0qqY8xF373WrvlrGy
lhbJFvGat//JOZCHTlw7kFpl7nIFFjbL9LAG8iWHjfk08M+0cGyMnhUwtFz+Lya3
BukzLRbjd7e60dvuqFULxTgd2B1fKF4xQtTL6Q/hWuwIf6L7OlzcqgzZgqz8NsZb
KC+mto5jAU+Tp3jyNeVXBf3K/DLbJttx7kUTo0DkP91U0BLGJEHeUWPLjMp4O6Ak
KsaVBdoJdsjU+F3sv45/qQ2zDFSdH+a6UxeThF8Rys1kHFEZ+YUD9d9ASrBw7oMk
Vm0XyXwZu8vFRNCFTnceE3PgXs0tS+jKp9IhFnyaprQIyRV/cMlvqOWwYSIHj4gQ
NCt+UP8Ly/6tkIwt3bxMjQLDZMNANHR+P9aLEPlSK3DzRtzT1j9jk30ksfhswEu3
jqTcmXACXwjtdYquRx7ASzhsa1LHZHpHzMQZsDDlaWVfHNyCnfKzzOPTR6H8cBbS
AM7fXHeNuUTeUUwfEHc3m/kBTIH6kXCOYti27zxJNeNt6pcbALi+ghPfjluKssIS
FAzCG9ZIu645rc7PlB8gSH5asZuk5zevmAw6KYq/WWGP9fOAZiQZz8MkHtGwwgJJ
/Wu0+E8MGFOfx8cY6y9DERgZbTtsAX1kpj1AUYlMVaW9ZBTOntxAxGknpCVoPQXi
uKH13LUjvmrf9gS245hrXHDE5fB7ZmEplCjyMO0KJO9gSKSM6iyqAhNzoviBFQlW
XPj53LGTnWacqunUOI9OLb+ZFdZS1BgTZkPUq0OnPXz5SAmTKru8twL2SbO0FSf+
p1woEFQgswd2P6qlA49uRU0LXoRZrWKbIbRsr1A1Y1Yvrw2iHXM6yAxSXb5TBc49
4ulxaOpz4ayMHn/ego+C2vL0nawNu4rk3Zw68GpTyWVMUwLsHkJlT4pGJzQCCfwD
FNIo+MBZgHKsJO9LI1wydhz7qDmIa/+dHoYdyKG0XP9rqdY6T+z8R1F0kGGMrDRN
f9ggSryLqaVScbmixJ2C0iv68Gw1z9CxVpOGI6qONt9qPd2n3WiGps+l0XTw/sNd
Gd0V+vJMxHlx+6SNoHqngfSgMxoXDZBDsg7vm85KJz4zb0VfvoCqwhtrYN0ah3rq
Oez0rtRPPMy1Gk0p797vi1FhYWMzoFBIxK4Pn4XhxMJjn9O5d5fpXZ+PdiU8kMGE
r/1AFnn4uvcCtDR/BVY4DPGrb38bdsYZL+6taGRl1npmjYzEsLiwc2+Uv6OOyyyn
rKE5XASiEFcB/SfSB9Omsn0ddidJWlA4JHnN0xkJd4dsz5JSgBiVBhfWRmMm3mNh
qG1Wm1cbCJW+4sbScS84msaBRKtFOA11JD2NTNZKwa5oAYo/eqqbsHF3jYhBgRPQ
xIBQaGPVJq3pskda+p04Tqb4fHIfa+ML3GczwZmAXRXHuWjPrlmTZ7LTMUIMEUYy
QVfkNGBiNbQZvy86620h44qHcDvweBj369WUqdsfqpaHolrtCbgMsVMDd+7411WL
j8p1j//YIckkLyko/6tkoxMU0UwRxhY96XsXpdqlK33WRCDaZZmTSK99KLCOwIEb
Ld4+ZxGTw7hqHdVDp/taC3VQX/gdzwmtBB1LB1GQZHKTt7WwJ6V2hJHs0uoC8eMg
8wFDLY518juxOxpFs2dqnb4YZHNCGhunNbQDCSV3gdM0JOrIuKWawEY3suiFCMNv
VP54pMda2Q/+A/kF3qCZNNzz4Gd0ef0Gp60R9n25mhr3Lf1i1BuyyUOY4TNSe/HY
1ed3qoqsb6f+izDYa6GtgUkIusrbW67xaNzgt9DdtDZUcE3GkapePLmNIa29o0xR
YpIdI2xOj+Na3qC9uSbQKPNqPOlyYIyOdvZ8sxN6Ujyl33QxO+WcLrmNVuc9Sy5b
MMPm0LRpa2ZwoY7WrrERaUX5UXwsb7EfsG7/+9KBbUdg7BuwwPQxzdyr27CCL4Zs
Ka90RKlVwvcYZFgIEeHe5YM4Er+D19JLm9nBlhsEI3F08BZKkpQjrIl+rAhuDHhZ
U9pbKndsmWrrywIomQiv7YyKVKmtWqU5zHM7THBYZ1YRD871LSoMAkshaPz5eX8X
G+NZA+I2hqcuT67KOGs/L5ocN6w/E25I1+7kTLfH96PwmVKAjBBX+G0r77nzlyUM
wB36l1FtVV0sdiLzJDWTuYmvD4PLpQNnXY0519qlqqNHPn3wZSeT6exYyAeELekA
0oLtYCXsw81fc4XVMYB+mtLbAzSHcWuozdf3m6imNIZotiJlt2nkvoV5RicypmG3
BpD7sdus8oM52JFALvXy2v5QqlFNBThjOl71GGOgeu8JOtSsyrYQh/BizPhJMDzk
pYPCFuSxkRoiKDJQ4mujbzu4eYs2msL2Gxg+sMFYNK+y0dapkzwl7euq/sqZgLxT
JD/Csxmwy16ZgsYkt2wbbMu88Qz6LvlRTSjNjy4tVwOsK2RxQlLJ1EGI/espVBEq
zudvqobOYJ3wwZQOnPcVjE5J6NmR9dwUF8yDenMwpUFQSw3P3UkjtmLcrs4d0u6S
qwTMc+KHOKvcciET0HlqWZNTgC2clcXltLm7LnZVX7nCBHjMCIg7ryaikIIcVuma
jjWS3perhEhedIlnjRVt14KyjeYAJ7JgD14THih/dkhdlKWH0hP2awseRh/IQzt5
JaTBxQE4LhYgqJz2HI3l1b+D+QsVH0JNGUPVeeIlTVsb7wpjjqBCUzXEz9ZICi2b
nsZ5nr8WSsEaaqawG73Meuo406nWW3tG3WQSdEc996UGbnz5xjGgtgwGRi3hDIQz
VFFUf8Fwzq8ZUBYDz45gDn7X61eOScVu2NnfhoLPIQI4/WeQhQnxo9hUoChVxohX
bxPyWeNDnlFN2bObFjr90r8134+WA9gheBUj8BROf3SXMLFBeIfwsgxcZmIpdwOM
GWiCIbq3WhOYmeK7NNn5PCwdkgdRoE6avoZjatPg+3Qr9l9fiBaSeX6JG2VPo5JM
a7zUhhwFCAe75U1VL1J7YiOyG5N+pCKmIyM/Pdf9xK8Qv5qaXOvkD5yE5lZcltwU
//JKsppPdVqkVRvJVdCOj6Y3HhMZxRqdZZ50MUJ7Ya8DntSQ/5GHYThklot4BGW/
FqUklvngvszlg/Q8AoVcaQ7DXSP4vvh7WKtcEq+27A6oTRK945NWe7UiKSvJ4k/G
P2RfG11VroEa9YoiIQ6+NReWsvCD4dVfHtrQdLzeqxQE6UebbjJCWDhltvwVNxUF
zH6I0HPghG49w2TUEPcHvE0O3IPSNKmio5Z2U/Hyfooc/rFSCiW/2s5dJ/GsrO98
fIvY4bh8tKpZFNLIZFrWEg8bnyhjPHkxz5dQmYIPWmk1qX82ZaXDP69Uy8ez8c/P
rnYchX7Xx2CtIozpYA5+Hb8bIshVZo1HgrMFsePR5+SSxbYGYKAP1hXEzLcjxM3b
QQNeb1GMZV1vDJqIjaqwe+Mp1I6dLESM2S9ISVk5y4fKkooroJQ6lagsPamwtmL9
MDzMzRdBQGgTOYvXCU2izudSjKdiv7SlS91Iu9rJNsGPi80anIHji+X9GqzZpQwS
vduW92h1GM4R9xHjGAQrtf9iRhYCyhgV3qmrufXcUTSVYTit+n/7v8wQIvvADH5c
O+ruD48AW2hHjUt/2XrOlvECnd5J4kqiWrE0ujT1R1GcrMdOZv9Z0nJcqErQ4XHb
zbFdW7f6VWMY/j+FCiZ2U4zbD/UNzPlvSNFkE8KJ6P8NX4A2lrOjQeWhMg1ak8O3
0GrvYAx0szGjjOKpTxa3TtOztCUzDDOXws/pgC9KSid8iafQwaSuYVzm1RBGbP7P
FiNMQbuS1jBaLWM/olr/YGvF6UbL5S141O2ltlbpd4JKs+KRTnmhVxo5w8n7oyRO
8ddGwIYlL5wRILYEdws5La2yaxWXNAf+YGf8+c0lcSQsWZK+Kq2yR3Z1XvG2pl5l
2Z4httcMNSBww6k32mC2j7vKHo90Lnt6SleSh2iUM3fXg4tWm51nLjYCCl5HTfS0
xlNOkoV5se007axGmxd3t1HjJOG/6FifBrQhLylAEQUVOh4zAMAHP4xN+prJPRr/
l0CrJPCfmwPAB1NX/fZBd/V9siLmWsXbMKEPZzb5bRKfIHf1cph7QIxDKnjJ+d/M
/FEZxlN2e990BFW8xvx9253epHMWiGcjYQVnYaJe7ibMIvUKXRBrFG5s2MxdYxpf
3yTEk2RpsqTB7qXusiOSYpwrw4wrdj+vhxHm0q8vaCQ18LCyKfozD68f0nkY2Oa/
nMy840JP77eShT2KB2oRnf22MWzaTY2et9qzt2EWzB14WHeWRIMeLyNKSMjefnqF
0G1Id+B8xuYa/phicaMbyhlYjYcSqGeDtf/ihzIIVy/OyT/Nm6fqVXQWeJeJz8NC
U7Q9wPlBS1PsML20SAseLVIjemlCUzZl7ER5vaJr4BQLyy7cF32iq99a6uJxj9Vc
i5vOrLC8e7By9Zb9EGR4EjLdwSAnpKAmery/vezmj6AKKelV3kDTgBY1BPjM2DWF
Ri0Vn8N8oqAnVPw2yk5V2mX/cYlf3UYI3OtjQxjqAjWyR/xEXL3ZNh6nKdkpPrMp
3bQP3IhJWX8keDDDRi7hbc7cu1UK+pcPbdpgP6bFTlyEnbTY7CTg59JbTtA29cY0
m+5GTByVV+91Nl3CN+lfxCcVpj2aYZjOt0SLM2ycqJC7zQaGDRuQDEsSZxpYkBq/
Rbc0tc3v+igNdH/GUWcUinWD0vZKgbZ3Dd1+511bNhQxO5fQgPgQDBmrnUbIsilO
0wHMLkAuemMtlC00aVAcGcOC5K/QakIIcjbJwoaPCOcsCVrOKAXEd9WLt2CRz6LR
5WIqKGXUocnSmjf7fcOmXUIWRNPOkZYUYIICHEJnghyOJEzdrryiKvKbw5cpgkZW
CF1LBi6DbkV6/7fzHydoU6tv78O4nS96OXmCSLNqDUdwOVa3taBLxk0CXJSD6Dk1
kbLhPec1wTdYlro7HFZROkYlXdVSJHUBnpLIETOS1g/FQOtaxAlefzxqsgF7f0WZ
QiFsUIYpcBdnOga9quZPZRGE/kyY9oSdhOxKgakoYDfUlN6cQrkbLHrBZwGpQEGM
/t4KiFspX2r0sZEYIw1sUp0T1YAWd9DXDwvPUHz3wbTKEaEECVwdyxcILpuvn4R2
ej21JeeGSBC3XaiRSHSpg/GHm6XW6ZfW//3IXTkXhGGokn8uNaiAw2eEa9jutK02
mMEa9V8hWXZswsHu731mXJumd23o9YrU8zE0bRkpMMJO4Eh836qRyk9uM0hkeWjG
nBEQ1UCxcRkt8bkBJuprV0djHq8PdxZgK/uRAxSrMPrbVJ0QgtShlXzXC2XQ7Ilz
mg95B8F+KZSSGOPrsD0U/hHZVgE800DsuRMQJM1qYCmYP2dWUN/UDjV7Cw5vQnzf
W5ullN/15gSsSgTDrobNxl1aNAbyx5EqBYTESLN9HuqqtjPzB5qAUFAE0QxqnF8W
yHufxcQQqEbNy5L7PsbpB4CUTr88Wo4h1+kLpZLM0NXh4HxjCXHkP3SRaaGBbe/x
4BwDJ83asnxuGuoFoFLn9bHhvCIprnlDwAWufWTmzfzcHjRVnhbBeZNh5nKteZOa
Trl5pS4uGFaDiNqLE+eZsqK7HhrJy+QFbAais9Yah5ZIh64Ud1dV5VADODzPLRH4
KuawThRh7k+FVKlbTQYBA+OgjgQomXW33N2E2A16ptNTMDr/CojW0rfbyDi17oxy
6vkAZjfEO5hSVt7x0tEv6llQ3NYxp+BZ1HV6iiKPgRyZk2+1RLXp1XzMlWmyE9/p
PFdf4VlIk6zDcoveTLjLrSbQdyI1JhAOTKp6q5JDt1SpL3+ALo4IjLRFfoWlpX/K
+V200rgdYza/JBcY6qfWGamJ2NIJY+IvWYaOU2VhtsoxofnkI9+lBUdsZlYVJSvY
w+B/hU5jW/JuJyeSQ33QvUawt6AhKDecvunSTbdHfmzV7uMqoLguJdnMfMtKV6EV
VBpjk19o9nFWX+qJKWM6LiJtexzTV5fWT+rrLyYpRf6M/9E/13DxbfGd2nVf2d5+
/vr16U5Np2vsg+wSCn2xEkLEdvmlgyZoesVaibS5durCO8s2mTI7LqJK+FMMOC01
50yWC4NgO1tk+32f68apDEzZxciXMJTy6j6k/TvEI0HxBjboLo6PCixeZdEhcrcX
W7jSfDbTIpq7iO4dHJwMPgNhhaiKtSIcVkfLj4Un1//+/XsH65tLaeo6Odxt8S6j
czyRFOxQonu5pHqMLOa2kz+T4HRJklsT2mPfa06T6ag0i4Lrca7/86SxvFu2cl+3
F6677d3s4LdPI91E6Erdj6cUfB0NQcep6Zr1GbpCK+JHIDR9OSXP/cMQBuQdYnhI
LCMN9Jk4G8fvO9xopXp9EtJuHY+Q81iWYON40/hHNGI7fo27e1r6UWo1vLMl0Ngd
S9tjSYFYX1i1h+mtSIeNCXrUN3gqPLtOf7K8qjFk96NTqz5zIuVjOawpzMdqtPl0
1au5x2BrKCWtsWc0VTo/+VDgOciB4lMERx30Kbh8U9Kg7WoqvMzo57ge/dkd/lIe
bBALeYxbPm5JsDWQ2ScgC5Eg1kB2MMZH2E8WufU6psizv9EhC/uTmvDC5L72ghCH
92RyEa9oO3WxTuJlMDUTrNn1mzf1FGXEGiAdd6ey70Suxm1iGYXBHKuCmNphAhjF
AbB0R/ffQpWMbgJu43SzP7C2mWYq3seuhgOil0HvzldbB+upW57VIB4YHkrP1cvI
qOrkVlysB0uTkbMbjeI5u0Bc6EyRqalFfEStWQxpU89nzy+KYp3QrT6h8m1+XXtA
K0EehxFfsS79inhyIJVjfEwAGH30c7ztuoTgLQDp/fQW/bP3l+glAD87Ihav6n9L
BNvjfPy2KMUSRshKOI8P4vmK7BJ7Z4m+8bFqAEENi36KWgPz7+PawC5eD9lh2F/r
q8UkG55sBKD6qQesq1U4K5upLeeMsr6AsvT6618DIyRW7mANTs59wfMRA919g64V
skJyTcmSxnVbozQhPZXL/BtstUeP/Wc7ghOFedjh6wFSuLOuW+JOeJCePIldxbML
6aorb6zqx2wek9Yl0K9+iWugAryrTZgd/EBiJxJoau1O7ZXQRbd3mFNAsn5Tul0a
C1TZaBoxIHnI8kfwUeS4A7rPcrWYiWkUUJvrW7LJHxMlF1IqaxFdfmh9U+x4ujT9
C56AO4qOAgouheTb07US+TFn59597P38ZAi9kl14H1VQO5bV4XVHxS+MR6USaeO1
VSGve0ELzswWohQv/r4Ri+4ZwvzCTTnTHXco4OTKnzfXgudYlopsF7N50K+1yEya
st7JZnb+pgeUeYgXQbskICWRdMUNUxsH6Mm5GSvDH2whU6wWr0X0XvrqZzdbof3a
dWRfQHOhocl5DbVQjBFkLmwCSHhV+6iPZM4/XaX7wmb3mV6L1TUiaJJf7UmLX5ol
Vdbcbd06O79lFhFghQA6f1lBdpy6Q2R+Q/6ZogxpqQcrRZCLlIH5xf5HGYywX8YH
Rz+hx90YYB0T4FB11Jb97MDy3KArgZ2vF9k0VenY0fweCqxlbR7xe6AMjTF9mZdB
IgkearVa5FxnA5jnDWuikzQGaszQLxL2wZB/uE30Glw/6PJgI+NMwQfjMRozYRzW
GpDky6nMFvMSdy41KlhdP0jNw9rNLtllYyejzOAT6qUdHcKDeaAV7Lsfr2sCzkYC
kSVUFXPUj//1sUNJB9xb5L3GqigD0L/aw7zVCjK/q9BvWLPDCLvmopz7U0gNfX44
WcRRil6IEWDOuc+JXDxm08sSIr2dQb4V3WFXOYqwurBCKEKgjb8wVCEnmY+q61+F
u/IptmmtUb4l6WqdYEh6d5R7WsT2fbm1ZKYARf/ArwH7GaYQPZ18sf2xAcmGbgXJ
PZfuJfcom5Y2VMmtzWehLFh8c/TXr8nNFsr7B+dYsfMGggXYq/uTEfLoTITOxC7b
v0Z1LC16N6iDttlRovWIhzatOrApDYJYxS/j/zb59B712QhOkuVSnzwrKfcBHZtW
rFYIuNKDJzo34N+n1WJstbcWgnUMS4VNXbaQQfe43s6qLDoBEC3s2YSXBjBpQ0Or
gpoYQZuIAA7eJEzIM7TZxc32Lx5EwAE4ScidcoJ984ADpbwpejbyiRrivY7GqOBq
Ir0KJLcpNQhSZWQxr+s9tPxtPuPg8Qrba7FXtf73E69Qtaver4xV1n0knldn5+Vp
NBOs1xe9MBg5bwKHGCkh+VkVICuS+IOM6GDxMbXE532iAF4mhfrH9ajt/XMQtiGc
3UQPdwlGtbqxAoLiGvQ8Oy5usvpkcKCwn/k09eF4ugyRfX3EhMd+jtPYB6IaGiAX
HDcgEKscOX1vml1uiXbW+xINn+/6De00VrnDUUr0zyaJYMf/j3mFuFzbB6rFvdbY
Edm3Djd6Fbvv/kR1euFgzearqV6nDGFJbuUAWxNfmfzjR0/Mmlac9fZgquQdBXYw
VlMzt/7cbpjo/tZE/GRr63SHbWwYgIvyfUNAGaAsJosjQvIDlJZ0V0x0dXjn2xpS
Ps+igtbliJdvqvv9sRwZmFYpY1QJOZfxMtFIXl/+yZxd/F7BQ1dQ0z4l2D0i9oJF
19fH8Dz1uJLh4xECeqStse5e40Q8JknVR+mvOwOu+7CSITgqv6vBqfpvK7IOGuFb
u6WV8EXXA8lI+WaiJ22zU3AkkD4vISKTPNaEjl+oAlfeDZgxcDdK09zgek/yAv4n
JGV+USM7mQauyl6aP2hisr6ogsJgqIJo5ipbv9sZ1EmXpdrX+XJCXvEQRKp5gePv
WPPln1AKiDgcb/KnFotoB1l0s9iHk9YY2dMP92rCqx8FHzzVPQHcA3V0VgXA7CsW
izcWyFRed4KOf823CitTZCTcMDmm8JJnh+WWSrNXET7T2Fgj5e7Y5N+nnxAt1G+t
8IO4V3KBIGI5JjUZ6Wmra2a1EE4A3rETg60rI4fY1pVwVJGE+KKzBp2IFuvZ96O5
qSWYVTXlkSblEGN/mplvSMbkTIHjnEH/PsE1vOZMuNV+LnSA0oxk4tNfTuU6CjJ6
weoxV/tDXwQoDWoV8ZrZ53uyB/yrLYCLuqzWiuWJw+0tNwJ7h83mGYfqLzig73Pv
Jgv6BwkI4ToZ7LGG0OnDDaMuvwZzi8NUFzNsLOio80s0E5jq0kOTBT2NFsu51tLf
p9JyVc/xYAoNc+GCNNcpYZxv/oM72oASP0V34oPme+mesc97eQwarHfyhP7ZEoVy
dIjnMVH4o14bTIE7JZPoGjaiFfo+erneS926sdHJV9TK+9YDRHUe84EgljwJIpq3
fiMItb4KZIywIOxytR8LnpJPpX6AoOc4YcCAMujCPo4bxjkAjw2oC8lDTGxKYTWY
kaV07Uo/6UQGlL+Ta7JCEq+WXu2fsVBhOOUeq7BtX5wbByu0cSFoGNOCxm+eTiBF
C4CtmbHl7tZRZO3lfkmvCH7Hvda+P+wSkCds/ZmAPgSkS9VkQOAv7SUBaZ+e8OK0
hc93VCFClT4Z8VHp+vaDFNvYyvy+eFKWVAzzSF736QLZVXGIsbybcEjNxuLWarqe
KZPPx4byRTiKhgowUMyysq41C4Q9g+KT1oB4ioZc4wNfPCvTPKL0lO+UuSJtiius
Ut+f5+7ajKcv+sPWgbAsxAaDQ784msrRLoahFN/WMFP5PvWzpoOlziGtEI6ibNkD
RFVOnNw/c1MfgcfTu7mxkwOa0a4Kadvm7Os+WgiNIv+8Wt1DQTDSKvjBDqoqCl2Z
9k7ex9FLHNnT6HLa+xQHfYHjq5oN88N2UlhlJJclmyRiOjE7jXd1EciGqS0axooj
uhDUaY0GbTMzhB6CDZpzB3lcj+WYyJ5NyimtgjXwdVTjNPiUhf/KNXPOsxkhFdAa
hgaV9EaQLhM0f6+LfabNcWDFg5wpvNPqeqn7fCs3oEJpIlei9aH8LJS+3vJJMqg9
13q2B3bmMKKBPnoBbngeLf0FafcLuKx1IkfPFaFyi6IJEvCDXHk1jnu4ABy2ITfT
X7mALJIKZeUdsa6Q5Dmp4W8t3IRTklzh5CzkhUdFr4th+c/+6DuVYKxixRpEpLfc
LDG4UiFNfxWBdIQmg8wbdVML4+ekwxCcU9CtZc97xvFimMn+NKHzia8OZGfIsiKN
vd8gy3azjsgU/ldOzZnEGxqafW/Ee7KwQZlTLvl+hNnOUznej+misDyyZiM3Xpxq
IydYZdBgOvZ87pX+T5eOHHENfTbQCicedpqFffaGkZDQU7AhGuvqJRNwCVQX3Xr6
4K8KYvrUHtRBbSo6cTD+LYSJtOLb2bz18Kc1GqKk9U2Z4NPIxnlKAvDKN28YLumX
ysLP5CyBPYR1+wUoBpHu/2S8F6W4an3iWeVq8VLUm7Kh3/T5f7/fimMis60YF+c8
6a73niSaruJL5/9PfbwMJfyIIvzBMD8S/5xxXVccsxz7ZmeP87pfaRfZxImC1MnB
LdFaeiS3s0AvhamyH6DJCXJ34thX7SYKUj2a/GUUvYhhDp0vI5pa4In+E+gDVJww
/CDy7fcvqAd+jCyJ0qe86JWE+OecM3NcnWiiprunrj5c5rMwRK8wpM2pwiKxIMgN
6RDbFT3cvCZj8ltIrtBk+vMUUaqDWHh9XCaS24si7/MVJmvZah9DPVhA5jvYFK2V
06qW0/E6Ys4AWOca34VZv8P+ulSSSNXlAyOSyLPsF73JoebxIkWvDnUvFe9Ybo6y
iE8SCstlf4QTXHosb+l8vQ==
`protect END_PROTECTED
