`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDQUhATeoMLJf51rJS/D5/yFq+SS1qizHL3UQrKD3GE2wqanxXGbrNxM6UHO7JmT
EK4ObxHk4E3F5gYfQe7GikXN8bzm5vhsoY6jRR0KbpRYwfs1vQRPInr/6tH+Iwg1
Mm/OoCA6wAXGMJ32j4rCaRX55VBT4MUjNfv2cg69NJLdbB0d4oYE/mb2Ac1Zj+iN
Y12v6caowx8DvRmpFcy+rQiRl1z4iPRF0UaW8RpvYX6UvrJBhpv55IQy+0wpa4Ry
Ih7yP+POLk1aBBGse73Zxx0dyaAi66P+YfAj93od9HHsIcVMU6ut/r7XSppuG/ge
DDZcWTktKp31FwZZp3Rju9eKjMKtsq8ktGarwXZtfkitOneRkGkwcbKmt49wK0qo
`protect END_PROTECTED
