`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VBQicGIek4xNc18YAxoabJtQzlevT5QMBepOFFVRcIJ8mnQ4EMiV/XnQO/8Z8tjN
l8E+jPNB3i7XeuMk6YN40tAVwvkuXSofbhWTQQlH/OH8Qk5yQ9Y4d+PSYvfy+aCr
BDqA9S3igGj0GPO+CsIn132PmAhOAiIRWUsj6IudFH1A7Z56zudA/u2LTFOdHIRE
wJR/d/5Lyhs1jQbE7MnJ63TMF17HaSmFVm79fUr9Wz91zn+3FlGAuul9RmLzPoRl
unopLNRwQ/gf6xBWT2nT3oLYWh+r6ngJgmkemRHteoeBlAVZzgx85fvM64ASoN/Y
KQDWLCJbl/rHbxdH27BP0JvWoQH0enouEV9LJ1NFwz7pHPks/VCK5pN75O43w0sm
sqS2iq12m65d0w1A171wH7TuKA3Ic8ZMEmghsToMBEQ=
`protect END_PROTECTED
