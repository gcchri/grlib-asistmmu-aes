`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXiLQVmBHEimkutSDPjNwjtz2w9lUc+dVVjmen/Gc6qGUap9OGhbrz9mnIzm0pJt
tOzUZfpg5j5ZB3rgeJKWbKr1Rf9wS5ZGprtcPorKsUnW3lVvEgtKNDfaKd1yk/Vo
mbIhgiOb1tsAYZiw//fHtBGSawQGIpu88ISyPyLzB6wnJ9JtW50hfEyU7S9Fcw5A
ISFAQcLKMW4tdDPAIhPYlAI+/yJIQiuqKItPQmKxXnSnhD5cEx69wqJVxr7ra+Oo
gZ/a4PJ2h95WfBvXJZfDXsujpgZkLxoXZCVLXt2es9UxM/yqtSToELCh5A9+Yqyb
X3oOMSIG+OAdB4Tyi7lIU+VaCR8Z/Eua/FE93CglPEQRO3BCoB1+jVcaMupz80B4
okeS6QFFAJe4cRtTLqgnPoZ3ipfwHd9UoayfSwLDW6u/NMkGcyjCJcolOrm4WSYv
+C9mO3ufF7NJAlS82bWR3Ohh1CeVB+l9su2TaLcbp3bgqTBvLvz8cyfKl1Nr9Kmj
T5lAIvbh9Bn0O1zCeHn/cV7gQYdQ+H2fLjSLwSJgrrMQJv2F5nSBQLf5k/bpHq2J
lU8G57qQOnH4d1KVqncsuLNfwprzcZD4WJxu9fIQl0k=
`protect END_PROTECTED
