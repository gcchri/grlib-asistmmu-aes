`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LnM2T9w23qF9qy60bJ7WazUM6hOwR/Hnl3ZYAd7E+ja/yGRnNDUTVzcSEM3DHHcp
EcFy224Re8/jx0pp/F+Ym6haRMmF8ryimDI3p0O95/R4VQn9PDP2wfn1mc+uoSgl
hrrow2KdhIrdWkwUkYzNSBdauo5nOtfF8MRe4hv20V3rFclS+E6jBMDl5ItDITyj
p3b1+28LoxDS8wwPB6aGbXtm0V9sWbEprsEvq/lJId0idxXyByBZu6kU+PxfgAmT
Doqu1qhmWabrCoJn9uh9M7mp1GpVZizvqh/U1aXy/fbDOSpvpWtSq9L0/insUq6a
H/XrurQwN7xufOQdTEJsj+Njn1/MCdJeDf8b6KlVH0VLTjkFVIV00I9mLwsJtk0p
dC52ECkMohLOGy1oE1eVuRs78nwdI+/Sp+gKaIhfbEzbtTbESgYMerRKgNUZDxOK
RW5Sg2CwMyrh8/BBIE9HYSZQBcqPIEMei3Hk90HmefUR0w8lJGPcptV4C9KRq4+/
4VgIS0mF90JtWGxl+/RZhelNJrUqSDunmGpQHYVNWjrpopu8SfTE5vs453Q4EHx4
`protect END_PROTECTED
