`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gLtrJzINDdMPmSBy6EWUCBoD/RXKE+EKR98ytAT9cbmrjiy8iGxfj7KKSvI4o/6B
eMYTgH+JYv6uJeEYw4GnJRYNK6JVG9UtPnswMCdVSWDA+VEDN17WLAZioslQdfSA
Z3oGG0aZcZWF7T2J2RzVi1UvHX/sxPyLFtowwn2+KHl9HdGSayDuJduzEYTqmZSs
qwBB1rdC8bVNzSHdJAkicAoxPAIIAiNkcDAF2ISX9dF835QIrTkRORTPbE3/vPsS
N2Vo9MXZkuy5+g2Ow6PHvf3jb/humCGXftzmZIlze41q7NfL+o6enY3Ilo+KAG98
qyiZOTGDbRhOjHxQN26ZO4YIacQbnnhD6ZCaCiEDnenq1pTDS1LKxuvYXpnkJD3r
IbhotC4ujA+Ev4A4LjsU95eoSK1ySbpTCUnDKqnvwH8=
`protect END_PROTECTED
