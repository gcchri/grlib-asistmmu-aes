`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RVQvM0ZBJHWywcs049MiNLH/MRkC6TNmGgz38Y2KCa2BHUxt4L/V8Qwu5VwarZzU
VKpoj9FFxDVx5PbnWrTshwnYQuuaWqcLD7UzSAe92o8V9uQeQmMvtSl/d0ghgG2V
LkysyLc4Tk6OI3pNciSfwSP/D+YPJjAnEVLMtd7vJmfSaxPbXhfLsLvx/sYCs3yx
ioYBmrIwJYPe4Rh3BBH1DxU9sCcvskKmaSqb8LWEQgS6h+0EJ8vef1jpxhcAsLLW
Uv/vtbnkMXy3S+kdVe1rnN2IVwlZRAsCICiH7KmkzKCjDonPWNZIQ2edWZUYlmvg
jUtUoKIwShcPweadqESWn56lN+k9aSBnigCM0yhlINRE7eQlmRYVWkhDibQf9WYE
9ILUvbFdQB02P3PDCs0qDWYEYjYwG1ODCVvH1k/amccOzEs7Map7GizZFYDUDgZy
k3MKOKBi1+NfYp3Fo6fl1FS/fPI++n4sCzb//C7rJWb/bxuU4Lz+kejxRiG/Afm+
wwYnRaukEJbUaW+RsvmS/cVFoOUsDtxgexA5n2sr7EsN3Cixj9138gtUwv5Ybmyl
RuphBBKXUlw2HGlxnqA7MQ6a1dMNPVLeuOZD72/rCve72jaX31Yw8Zgjl12DZbdL
ZaYTOIn9ujG/u29W3cQtQq2bZThSN3lRpweDby1R8uBGoMOy4QMTMIsmhz0grP1S
MnL8MLKLOxfmNVFWN98nFe9nBeAaejkf8+wJMM0Qw5/6YUBAFCawh/hdo7/F6/sj
rLXAKMvEi1bIMHgToWzoYo7AzWYOfte5IQQqOaTMXdxtPa+NM6BRRRsSGSUgQ7OM
iGW/ZJvTsqodTj773G3uSES4qhk+ux9td6DkLNcb3Z8z3I4vWW5H+OjSLgJ9kdXl
pI3a+BXM4GQGydJ7BkGd9vUiCNHkFd7nGETaWc40tGbPqSXRNaAfcHHxoNYsFGkX
9WZn12ukWo3nwBpdb/9eQr4h2Qf+ES9RUW9v7oddW0ELmu4cq/4SflRfSw9y0s58
GYuCNwbZVq8LH5GrDYQ/dj8RKIj8ota4qt3Kj0Fe8fRPGpd0V1ltwnYC2Jqu+Rr9
U49nlQA4X6X+kJYUTLWsYpY9HiIZG+gmwFTjsviIJVUV0zGz2+Q2PdHZp8h7CQAy
sOWpUhI6T2TR/Ko2y9skekNR4p/yX4w+MPRnDgFTzh5NLHDjSJJz8tZq30jW/Q4u
X2Jea7ZQ2uM4o3zDBUgZi8rLu4cPG+Ek+j69HEfTgRJTI5vE6r3+7t9HCGhC3iYR
/2OmcJcNzcmirWKnRI0d9FWak4EowFmKUwIJQKzvpAROlX2UNNhzOkrl4rWbr6Ai
PCvUQd5NQacouZj3cN2yuz/97shc9Jty8G+1Bg5AHBVrDujGIWeAZSsygAJVbm7Q
cdw8EfU+e03rcpNnJsqj6rImFjLQRDSswy1lQNgLl+kpoCJZIdenTgpfvawDE747
Ak1dtNneqkkAWaor5YYDtCacYnr5eZVKbPBMzm2Y07m+mBAIesh781etf171uyKC
BGlTZPbuAdM3tSIX3833eiR3J1eLPOmo0MljowaD+vuG+ZVymdFXWJ6zIBB1eDjQ
tcC4ckBaM/5N4/9/y0GVrvjjcGfV/bIL6shofyJRkUKtZMWTMsAQrkiNCKfN9omM
0ZaTBWwOcrYvuIjAGM2TWXefu2uELWDw0KDpTB1eY4yWw7g/QG0Zbxj/h9bGytCL
B9TyQfpZ39dU/m5bKvGLY0z11wcp+mQtoDbisadEMe67ym6dJym6T51vJzXz9iHJ
cYTTL3FB5QhU7gW3y7S347Yd61fkfiv5549jCb+jefO82ZbTD440mX7JmrxLMZxa
aPvsyAfB6YWEEQjXoTnVCh2DvaQRF3CwNkRrBnXjowc+/v/hPTsa/KL3wUmU5RIL
ZNler87VDsWeigh9RhrZI4D2EwcoNPe83e1YcuwqaNnRjwnWNOSoOIkVHHvZknvq
AQWX59kXT+vbdH4p90Jo5E5WXMrfT4f0psWXdKsgsjEsrV2RREYb8RvdDuwkvRrx
jwGFvfRQwIwaptCYwye2BSTlvcF5qNA5Ej+J1uSAnDcOJkZS2jSex5axJ4bTyecv
9gmYCAE/Oq8iURn0wpQ51jt3tTnxpdnSlnzdX0pH0VOddTYOMctO1pbtZ5mNWXYd
95YbrCWcF+1j5uBOCBCM4i/KjJmqn3bakpm17DMzYLihHh3ZGh0wYpMBGXj8RvCv
Wj26n2TCiNY3azxSYdwLLJxsugclE3dI7ITyxJjfnMpVs3oXaka/gl3XXrwwLy7C
pKFSdQw9tvE+hCrzngrPhQOzCz97ncG21LClzXUofB1cWfAbJ23YVqX4snEDErf9
xPP6w9JpSxfN2ECb9x9M6E/AZcpvwV6xnNVHq7mfQabU//PRQyAwhq2xSTeg4HLg
KOmfbHrHUypUgu7VStw/Pq47B2bDVs+MtNnftNfq2XJ761iF7JcmG1DfD6zRFO1+
/mEatsU/R+EzANkd5W5UhYSOcQtYfN92sKJdwD048c9EzJY7m7MMb8TJsJ5v5SRS
sIAKsiqz+zcZYIXdvq8BJFehnJKnJjWEPI9OI4E6rWa7T+RbGYRDZhsr/u+mxu2y
s8nANEn0QTrkvT2Jqf1AtCYy5bRTou78BjJjwkQHq8fGb9Ov2hIaItlaGxC2aASF
mfjbGSA6V+6bREuQQnh10Wr6UQTYjPfNMeh/YLfOhF6XIjdUnMSRLsUOZIN6LOM5
fpLMFgDPo/cVwCEBeomkKPkwbPtUaEVtmY5DYWzn348CPu1ovYej+zsETIcjWrlt
Lp+cHokXImwFyJK2wRATgSECnSaMrlse7Kl4qg2LxdKlnoNpZDfGoFG1uEy+Lsb5
Snr+33OdPW++mzRnQcRyVD4DP7/FeSw2JophD3pt5pcS2ALts9ckdbmaP7I3TK/r
YPeLfTx+eRDB/v59Yb5jWfGxIzFmP+8lE7/OsdfyfRrZm53Ywj12CYPpFEF7/OVv
PVMskVsjDLnVHLvatlexh5YL3yVBqokEbm23yOSQuf8rS80LktDJMCgxPrb+BXzg
4bqnVAO0EFidIvWZNywoNutj788QldxAj6p5kOHTlAinmDoIv/GzQkqpT75C3oku
V012uNFVQHCqFB9iEXsDqTqo0LvJQGskZ3d/DA8ZhaZPCvDl4MUHmH2DV22N0WSo
mJrQ8HTyVx/cmaTIHHVSBBEwyUwaP9eNOyCn2NOQsMbS/Iiag7jzSwU7iZgccI2f
r7VGF7LqdO24GZWdf5I1TRl6wp/w766sJFSPlah/4C2B/61RqMxt+kKAsvdX+fTa
CuWC6j1VRyrhXmQ5e/gNavvO9Mbems4S6AoJ9uU/1Ek5eQnWy8EU34oc1BjPw+ET
gjrPJQarc1HkoPYiTqEyR/nHm2Vf27buarTrEdep1FATpEm1sHOf6elhi9H8KFDy
J4jsRMDhT3EoybF5/BLYty0CPmP1MXu/nwvZruLOD8LN8Wm+zKBKSU1JZLQlYJ+8
NdKLBeumXsC1fhx8K9I6Hr6oxqnKND1XCilI3YswYpjsPUIwVdeinyEyLYEWgWn5
LIXwb7JHibLOJk3eVUeH7txVSBrlkMbr8WxJYdKi0oYJPCWIrGk1UW/UbkCfmdKa
gsFa4Yz6ldbpfuo9zQdZJwU04x+QJYjXSo8gzexGQjWpXdlqgKlGojxwjljP+sYD
6LvkSAxe7GHFQqyUAizzfpJHjJnMlVuwOKs9erpiPZqreXLoPGhcU2kKvWBtVYOc
6JnXUcg65X2tImyjGnRPz+lKzr9pkAcyASWY66szZ6UMRFMW04MHluCLY4zmacLB
rdA8Uk0tosmi9LpOugBm7NsTCUMWxPLFgkzAQWeD6+iCZ/hYMrxYrjJRrUdJVa/X
yQaXOZE1j00Ldy4/w6uHL52aVD5B4ZeTSzJZHO4A3UedsF+Qufx59WAR6LyBoZrg
W2nthiWyxJirZk0PyE7C0E3Z9hg2LM6hW9jcy0E1dUXx9XA5B5F5Rn0t+oLxKr5R
SquDFXK4ecIdTOm3OOEnHO0CkFmT5czkNLt+fU2GX3JFC0rv5TViFpBJyS8nGdIH
/74Mv4yTCQqXkJA2AvDKVAtBp7t8cCCiaNy/okZT3b2PTaTL1PcVDys2w4K9j4re
plQlphbe6pb0pBJcEdWtJpOWa38WYVq1a8BBqQIjsHjNNlzwlQwXaYgV8WdHRPrO
UkhaFbPozUgRDIBbjvczoxir5taHVyrKBGlXL1XCVNpJvjiAl6AQCIA+X5+6PskK
QeRMhzHz6XfDXJ/n8l+Qvhd2ykomwuPiPsxXWhYT5hZp8YJadgZDTvuhH3qwEQLj
Rj2i4iKAFVKmRgiLjK2Sqif91z4AhJRLhTdZTu/B3u7dv/6+8oeLgSuZz7K52kFs
NvWKCu51fCwqhdgGKP+Iur5oiwxc+b6cQ9XBJf6OD06r2O+FDG8W3ccSKz79Nxw7
r4ouq/pVZB2dypmbeYPOYY0C9EswXfcyZ2YhcGh5FUpLv86zGtlG5gGlaUBJXw32
bRpF+PCydUSqPVkbr4guKqipfg36/wrC4ity3vnkZNiYQIfdQZ7BSBnXBA4p7r1h
4IJuoaIW2G7Dc8ADo7fMmjMU1Kt+215JtYS73picAbTU5kHPKTA1eoePEQ64EVTo
ChbhUdY+wKnJR4NboAgXjcVlz3fCWrqMyiZ5255L5bNhhozo5oe3bXxLr1eQl+HM
WaadILusinM+Ae+bECDbT/Eqj7+PeHCm6NZDrRJMse/TJENUbos9tzxheUZfe6gH
hrwsY/YjDgqP+BkQaOHYylgilIJMrjtKgMlJkAh4fKJcbpRtieYbawIUEr8C3knc
OPAvK7HTHNeiq7H9d93ChtLLqwnJaF/8J4NTwdAn6iZQLg0A76HVmon1UJtBAo2k
416cHUSXtqPK2hux5rgCpmM5VK3OfdwDRdgXpj8ucqADLBQ4FFWO5XakrOaJEgOV
j9kD6QIjcERCmac3Fb9pOLgnWf+iDSJrf/oGeWFwQu1HWpaXfZvv7NLDUzt9bU82
vIp5vs61cXqdTy5k/64Ca9mAC3sBxa3clS5HVEhZyjz4QV4uwbFNACtwnAvvHQWb
z/g+6M7oS74znS2Wuixhn/Vsg3ZLtswmQrs8tSF3chqonLMqFBXzoCgEGd5gcCPb
ParfCGtsPnXSc4XvnFQLL1W9R6TyoXiCbwF+wFO6bx53n4BakIuYzqWoS6QJWc5c
0eFDz5xcTy/HX4Pa0X0O1VuoGXYviZ45fmzWYjRu83RDKXuOAQ4lDwLSMTxAAJQr
VBl0U02EEM+/gJeqroaJR8kimjFMUt6ggbjfL2TgPwBmwtLzYjsqTMVrXHBsEhfH
q2ikxkiaU0cPBos4udAYZz45N7VdcLkiDHa9iqEWBhwKV8EEjgO0cj2uGqdRY8So
Jx1N4kIukpF2VGV6cIVMqm5UjlsPujKhY0gj+rALr3pm/vxvCkqu06p2RLp8a6pf
5eN0PhCgaZghVyE9EmvkYg3uhZf1l0Vfb4996+7XIjOBI92yO9+u8cpcZup1kBY2
Zz5qRXyiO4VvZUyNAo/LEyuvvELynaeXmp0yche5SUvyq0uLHM/7nXKGtOr3x3Y8
ZScxKNyVIsUMKOVZ1QN/p+OugakaGcN7STd2uUva+f24fO/pLVZ+UvMQmwzZpbAL
7cbh/Sm7RnCTXazPujWKpcvz3FmMZPW6GI4GF4gGX0wEn/2Tq0/k5eQb+oUqi3KQ
S6DtPFdTMxQIQgC3b271ZevLmhTebbss22wwhEFSVjh+inJBMHdJZmcNLN9Zckyn
omHpFxzcdWv8sc9j1HLrvyG9OCpCrY0ImutpuFrNu8uhvqf7b0cwAjoEJWoAleQJ
/9w3y66v1gM6xu1AgO/XK/hqqD7RjuiosCQLwbOo6o4BWUbc3WWmntrHoeU1A0UJ
l83teA4uD9f0uv1WIjQue1Tl+NNeoVTX1yHKUfSzW1aZUN2CHm2ZurvLP6Lv1UvW
NCx+wXb48MZ7RQKbTbl4apK8e7b/ke9JphjJpbOlFhP8DDjAsmS75+rw4ShRbHfS
x3HR40OXAmOUFYvNoALg3hHJOkTAY6qWhfLQOFm49URgES/wd8fdJ0XlE3taosoh
WUBMKHi6ShOUXoeqsKG46khig6aXEYsLDzbpSewP+iqEW7V6V6wJOxHhLaOhAqFM
yqRD9uq05VKgKS4/btXjUn4VluQfNWvk2nmuCunBNaJrL+0nAqvlBEtZGxUs4srM
ofQ/eo91ud71GcGXBRheYADG8cUBJCBnrx+cPdbWXv5NqcXJ8TBjczNzJ69jQLI4
3JAg09EIrMS6z35T6kY0X0+DMPSPKSxPPJz4r9nggu1QVFre1WttaAsFQIlvlkfY
DyjPBAjZqcM7zLK5QLQbCpHiK7NszB8bBkIyy5czFqCbx4ZaZgcoHHaww/f0yBXl
WZyNZ8nNwoJ84ThvKawkJpgCqtcCgIE7EO2yakL/cjdYGHsnMffZdL+9DaA5KPVy
Dan6MeFPNviafv4llInN+WzxK3BzdKMk4N6U9uPOORVT7DBuuJOOpT6IeW2LC/nt
he6UGuugk8wxvbn/z4pQrtBjt65WxSc5I8eHif9LuDFhUY5+3V2iXrG4ktCeirlY
SkHdO4scdipSdCo1lt4ew4YTx3iZGPOs7ve6pPYQBBxDLyiubNUIQMdL1dIEaCt8
W+hyS/48sIc8bBQ5+gmB655fK6ct5J3mgklfisyQRi+U1Uyg5+6H2tiz7ET8arOq
h5LdGRWnDpJNL2IHZTWXUq7Hra5nFlsHqe2ik4gk9O6FE9HtelnX+PnWl9o1umDM
J1dVolNGuP+9pHb4AOUtUWZ9nWahkm3IVlR60+T6UWVZihtBwrgy+ypc7ViJ7eUR
xceC6cmLgJ5KmfBlOtUIM+GQDorz1RJjfU7TFO5PPni0XQ18ykt1v/e4FO3A5ZP7
ZN/yjsdS2cknkkkq6Vm0JrDHf38fyjCT0zNXfk+/22hoK3sNj7FU4GtZ7cv2tprU
5QB3wJRPoKfGBcrmyzem1Sm1nydRsOSUB/RvpkYQiDJ8SHtN7pK+TOTtW5QvIREC
29yO6PnO1KXuHpNUbYiuYtX42kMs4XyQTNjL8yw5C/QVv+AzSlwGXWNRPfdL5ycK
1E0mAIPxoKbOoYvCLRWwlJ9IllJeZchFMlOpIy2lCyA1UWmnm/335xEZ/W5og2gh
JAlbq4WppyqrgKxPvw69EXjzvXAQ0iCc7gR3zTS2B9tfg7aNb511u1vR8xe9WFaW
NENpX9JWipkCfpaNndI1Kliajv62e4JuR5buOZSroYG2VJ6279PBs3qCxLDD6gTg
PvFiKC2R9O0rWcNj48rIk1kEbNoVxZAnA74DseUlnhQf1bDh7iHXI3nAlymK+AkS
WO0cvv65IO2sXA6fYUL5G40aeOyyiZM4cfKGvfr8nBmubadLi3Y6nubRN83in8Yr
N9rD7qkxy1nVDCy1Z+9TrILOgeCEkbNxGG0QVcy2iBjTotJP0pplm8Bd4zOzFypT
jLCgTpFQtdBluLxrvjQBxG5e1U1bdpKeH59hPNbpK5Z3fY9SUqrtOBHIPYVGfykN
mvR9bRV5XYUR86rl1+OqVd1rRYMFUvaxloa0Ya6yzO4UkNcR1QJW1TxXMy7HwF/o
POEIElFdbt5suaeK/CFKi2jpDmI3bh4YuHykiEVO4TNnIscXk5PQsj/D77qppj0F
Tn64NmzW5zkCd/nTmtHaRqQ+d0hq0GL6NVrcoV0UrwACbRmMuiSg7wCKzPUH6F5H
zKSPHnNb+xVRUpVF1/hnw6ef/nfxaP55xYI1ZSFZa0HQ3vgSOZSmu6LtmELiSQ5K
/p1ua7WwY+G/SpMoYCQ//JsIjTdZiBavrBuGenk2WJKVfCCABmXxxwlvRXDsY6QG
qZS8z1y3X8BIdzsTx3aM2iLTde6BaF1SSbsChFNmUQMfXCDzsmeY2Q4F9iGimSTl
b2mb7R3ikEjYrL0hi1p/BBdPuh6+Y/7nPWWpq8jBVlsfr8nxkbWPEEZAcwvnEyIp
B2uc+jkMkgmUwdUCyb8MTAf5iUZCAcYx7Vo7QPiPMn/h0K2OsHohF2GFajGpsF0H
UgZ6BlMncr6vLnoZFwr+Fi5DjbZxkoZ7umDJs5YsfVo0TMC9zVaKllW+hmX2IA0m
Gu5lbp3Y+93b/eutEoND4+x1j+GGDJmj4CK91jFpFuNMax6ncSjzkGMtzrY76Tnw
UpcEey1RSmtvzg3rSWsdbiddPSurgAKBXMFE6DirVc2L32bXqPlLUjQzPWlrJQbc
FhxDMZH27dw7CFJdKmAtuibUKzRU+8YOCZxt2J/Qt7rKQJP19ZAf7QAHM0jvYOKR
AIMzemRzpp+Q6wKxMdIU/WsKKNAH3qwqMO0g+UOILIspdEEYEsMWathBj+TPYuNB
pBNusbKCvbR46cJc0t1O2C+cRDjOg2BKzIbuG2wQ1NNg2WRKhPeCPFbHdglN23B+
3bQ9637IUPfG9mVlujeHey6dO67dZ7cmkHl7+wvoFo8EDEdj5uluvDLcbt3NQP6J
iXcocVRtgq+6RBpIkKKsOPfpUiyLw2aBJhTfLbRPmGSYcyz1ioYZrkJPd4c/ECGG
mE6LiJMT6azItsCIoY4By2O2fa+gxmRc9snJ1IrSUPxD1lajYJErA02hzCvbHWhY
CeeDMsu1ncgXtZiZwFaUlYeHT2bumw7GGP7t+yM57JdHkxVh4uQFJhQXNHphFNTg
opS35Y77EFVl+7G0OAeIa2x01W8NU4U1FraUz42U3C1nKGOkr6QvIQTK9ioCjOSh
HRY4DjHOXkXYJNusKO6L271AWhJNpIUogfqAmMKLy4AUsN9RyIISnKAoBMTpJfTX
fSYAC8apwe2oKQpyEsNl+298BaFzFndrGihuAV/Dn+/GUppsDYvusfMLfRgow/fr
vp/Yh6VmKg0BX1ECnXWVCvB25T3Bv5UkjZFqq5nEGvhMI/JGkY4WywV+pCmpqWdF
hJ0KnXZ4UAaBmpggE8CXJavZd2YpW+A6JNxuZVCYSkbdkDlvjRdlKn3n5pZidohP
AafUbz52w7+x6TRGJYPvCkqjpN/bssYtukepgRQ789iTLdoVq5Ya4/V+zgNwT6Bk
Z8SQFS5MFeuZMKWfmcUHhAcuGhMrpfXUpFgxIKXzZdOnvZshwx/f5ZZEluZL7fCZ
bZyiQygqxA5Sy3UDHIHC0565UHI4AuPTSl/IQ1aUDmiZEtyVJtiRbjd9c+E6lf3L
3K96VK27kmCFM5mfWSXmo61gdqnxJniOE6FvuNPt0N6MKI8IumONTsG6ncXCjzE1
3ME9GES1mRM9VecBdLqD5Gghl9QDPaNabn9cjKvBsmFDwE55AR/8fz2ry6kSz3Y2
IOfKBolC4zhPhxTyIQ6H85VUagepRsWwtp6hCrYL0meC3BKuSvCMi5JDfW8hDl5G
Kdrf3gSr6uqXLDdESvYMBHTlgF9zG5rcqHC+gjIqsRK+NwSw4BM1ed8P3f5XrzXt
U0mzHIamv8a0w3YWqYS9CtxTkpUAMTWzyPorPSqCA5rjzmSC3O33jgj1Gz36+LLF
ZffI6NzEmKDzXihhpAmoMVE8G5ipUZBFUNGAh4zJsjPR451HQoU3WI0P6FjoprT2
38iKZwW4UpbtjAahvU3+/JfRI0m3innhDNsvqFRZxFbH9dChHZAVxGTEfM+ieuPm
fynHVnijLk/jhpv5HvaIMmu2TYtX4n3BNcdquazVUEpGmroKSJPSqqxyOWr3o3VU
MgEQ6GqqJhZ3c+B1Yo5yXWOWnZW0qcKKf+TzplSE705bYPZKXotwIXVywXe+3qQ6
duzrNjGWKmH98i/OO6lV6RMV06qAjgvGjW+sNgQAgfj41JJ+LE1drez/yAdeG4Gr
XjprF0001hR0sorJPFnvLJGUxWnq4/2hBvF9/EeIRlS9TPFsFqlcrMzMQj9PxG2L
BqdyMtluzXNR6j5icDijaSYVv5ZhMuFUHiT2OkSLxyvcXq4Vapkf+v/4dtyFoiYW
GI1iLo+fPVQem4daG++qyIOa68HwxRqg1FnvILWdD+vyE/xDB5Kdo6LdJ+DlooUe
EYCgEo7ZGLhsv7t1uUoSxLxP0WW9wWHjuS0m52KP5FuVfNtFdf5qPyeruoEdf3Jc
C06F9KeRmh8lpmu0QNZhFHWGJSwrzV6fstip8FhkZfiTR5EcUjWOKoIirOqIN8zp
5ip+hEwBOnWW9WsMJC6xyTITYdtXAfb+KW776uLJVBphrrk0FvKwzTBOC400xAZd
IvO+h9xoijvsGFBGLBKbHOu8SAEAe/9k9r1rYTjavqtq6SnG+sIFKNpmZSGkjcOU
trm2aJ4yzdR6notQNsGfvONQlXetHoAf8PBfZB/sivmjTJvw8cRgE9bTATmlZJmf
Y6KBfxuX+NrcxYr10Z3v4b8EBAf1kTknJTmnL7X4R8JNfk2CekdxuYZtrYeAi+PC
OgB3w9asXIzrpaYHZdeKF6GFFGkaszLCEM7VJI6gITa/hvnE9qS0bxx1lCVAzUzy
llPDKYQSxbOOhAZdL5+c4IKMGxxIv67ceOIFY5WDuDFbabVNy1hs9BjAtyL4tgcy
qfjJPoPPJvfgBJVI4P0Yt6LHS2w1aNMtchmHZagaNLrqm2FfdYLIqp+/nBpYCkiQ
604jVkm/vSZPiozNd+nJGZjOvvnTnrAfG/ut/+JNfHWerJCdzChhbmkCrEddfijV
7P/7z+h9JMOnE/4fpQ4UpzjqzWd2DHal3mOqCBXfZ1W5H/D9KQNJaHzNUc8o74bH
AONLjem6BrZH3fPpqeTcScIBEcT8bIk+eDg1etZNgF5WGJROEBTFPfVzWbkjiBBd
fLpBOI3r7LEYPP+fvdBVn4XUNAAS0LcDJA671vsOIBpjJ8jnPy2Zr0FnOVVI9e1S
Uz+BeQYua5O/RN5JpeQyFf9dxqVawtan5bf3vcjJasiEMCbFTZlvgruFo7dt+nrC
mAGDiegurYilbGBnvEN3OPSfOZX26lJkSy4R7EN/qvh4OPS6WM+8pF6Erq4aG9i6
Pff9ORCH0xQLkbx43iZ9i7DmyHTCkVxhMkVggm63LdGqiWxKjT5S9z7/zSz1XheA
ERTrvxrYj1z7eKHgwObEmimCaiyNaheqKMDBjsQA/ogyK9XBkg1UkHh3fk9VTyDP
l002Wl33uDq6E6qMIKg1rCGZE8EBvJbH4Rn7029r6s62nyviQQqu+0xn/RWQ8PdQ
HjIOos8I7zyeguFdK+XZxbOOLKOz5lKn0huE+RtC0ENn00kp/WEyPa+pY0SEgozD
hC5Aew3KAFJvZLKxhMPhqo2GVvHEnfj8Y0BjcECM/OCE0S4ob7RfUnJMDmkBNxWx
QfmdeVo0qrlnnYJNxX/sFEHCeOwGllPLPLTwASY/zXfllifJr1//c5u3EotJZ389
CTgaQYjV6UxF+A9lxf+5WbQx+zM0iO6Kl2QBidv9B0dfXYN7pyAq2dTamAf/TZMO
qancK6V8OT2gUQuSkKk0lOtc7D9iwhnPaQJc9mafloEKjMsmJr7gyLy/bgMk751u
IR1xVAqgumTIjiaIE4wnt1noebBDBWdjpiExK5YbpWbCMZpSc9lZN/98sTfOPBrf
Ckj/IBWwNaqNGb7z/ZDkhCRPE0VmYeHPcJVWRgYAyqx9AXG102Fh//XQjEuvMyeT
gQJRqaiJmD4POdW70RnMpWNf5A4c4lfp6Pv/2Oh9m0VfO+Xvy87erNkm9PczAM6G
SsW5WuITHJbEJGQ1xrUUJamJxGoDFjugGKZ6MSgp+wApplfgzCV/5gkWth0rJYBO
EMoEQ2DP8OICOO3OeDc7MmH0lNBgUnRPVQubLJrv9hkiQ1zajz2ImcwE4qaa7Gnl
LTDaWDlH0Yg2X0TX94I5aRAyIvvdHlzQeOZtg9xidbPYRnNMz+LdSUEsXerNrY07
ROvRaSGFwMSAjlARhdkIx+HCqxe0WwWztR8JrEANEU/CIjWH6DhmNga0qRkHM6jH
5W8x7p8+fS9jkE7p0SGt/w/xhLg9/xQqnkV16a3CC+kAsTNwLF7ykr6f8SqGyfZn
EQWBmyg+8kATWqqCYWGgiLgRlkgcI+le/XNaYT9rijuWujAoQNchasuTuMg0Xp87
0FtMmadDG5E8W2VP3jWR2jJIuc2UA9TJfCGvLwhwcDd9rxQEWs/LyuOU8GDlD2Lq
+sQ0B4nKreZj7RQ+iXWjaQ1yOkUuttYZIWrVaO5+oHDUyAaimdc+7UQ3DnuQGfww
YyhYEz6duHZSmgm01lS7eT5eCVTdwZKAkG/eCvRuUpgqAx5H86z107g3UOjKLf36
yRr3YZF1I1rILt5Z5WcrPK0Mwt7qabM26Gd7VHiII95jjxrf5x2zM8Y+/5gevbNh
qjLdpRcg/6g6BkGFqMlK0IQ/kvqovaKfP9XrpGkh20CZyQ24/owXCh9pFqUxWcR4
PaTg0d6nH1elMtAupNeu0aBvMEn8sHXbZFCqYuT+43ZXJH7LpvR9jC6Zji2YRN1r
WNqyvDLlF74Hw7eFtXy2sm+EgaWnC2nSgrV//k83JHxY2IusDO36JoG2WaoI24Pd
++3j8Xu0jaqUWxgDTXnxyAJoD5f/3GDedlht6dBAmDW1tWn/E0k9RIwsXRHIDNgM
PSnL3yApIgpjnD2sHQUF7e0qOse03k4ruc9ghH/kHN+zNYxiK+O1l0UrxZJDYWRo
Z76skYxbUUj03ciU++S7P8hVCo8TddmeUT3+Bsb7baL8qvNM5vRGgFVdLvLrvowG
iXn4pq+minjRbUJUqWS2S5yHYlXiJQu63VswlhzTFXdWOga4RItnTQVT48aTPrEA
sgowV9JctIXjXh2uvVAesDVC1DyDavxxN1tacjYJT66kaf7Z5o8PpCwJL17tgr9x
9ihgmULRXWO7mOxb3rzsuHKXKiTQ89Rh1PYRxTiJeI3nmYt6feHMC6Qz5oU8I17G
90NLWyBAR3/mzxH8Ytk22tMLaY8m+IZP2dYi73Voc+lNtiBNkdOpJvDhk1lh5XzA
H4G0XSHPD/Jq9wnkhvP1iDIicEzDuXPcKIWW/fwv6Cs1bfBPC7vxTDzE8Yaa9wia
IHiZm5+ZdiWxTb8zYHpM4kP5pBsFWu9WrytfZTlFwoN9W2pAkdQ3x66bR/qb3R3R
IITOBjRbK4admnBgRxgr3ibVIQycCd34Z3HjjyD1qSoLC0eRVvlHl6o1h7kHPEI4
TOShICPMyMFOw8utqyszGISUK9HfbbMhK0Y7zD1vSXx/GlGspfAGK4ub6EzNHrFm
wfHKwfL/fkEHhhd3Ca08r26SrtuPDvF7dq6TKV/mo476YKjLKvp/wB+bo5TtUwGG
vqxiN8fqqNZsx6vUnchfnXKJJ7eJ7OA18GJoVXJjfn8POoDt9CW9InUN+amGwGab
ejzpZSY5ipxU+IUETr967XR4LfaVFp9outZSNkLizBXk5VFPc4d8zkAy43AlyuF3
tBubeO+11cUTfzU2Z3MHmLgoIKckTpX60p0Wua1D3umkHYH33VP3dlQ1fMsxZsHf
7KW2AVScwoMDM1ARc7iGB6c2eiR4tEgPu39F95LTLFnrjiKSH0Rf4S0ztw2jKKPR
9OBUDqiPkNS+0s9/y9mF3CuK2DozGIldyV3CO5jajd7Ap5MZuNRNcJSSzBmtjjJK
3R6qpNpHdQGH3ROKHc2k/AOJOJoXJQiL1ya5Y7+br8oHn2xkeiTQDqkNPYxJVwNn
91kTrdK6CVY/LahM1IgfNLV+0Belne6nRL9p8odoasi4JF703vnVVogdtqVpSOgC
2wuWXn3KurMy/u1EXuRCBcEKxPqiGUSDnC7WCwv8LIjT7H5JxoH+AVu2ecuCoGDJ
Q8aCLOk0ExAxBH/8WXwJ6bhOT0josbdAzdDB5sOf987nCYaikU/yp5tw6FeXc0Zm
C0sKcy2/xgfqGnJ8wr6DuDHCbUmivWeGc3Bd8Nkb7y/wLCsoRO0s/PIAWgDl7Eix
W+4IrAmd33UoDYcxVoWp/J5TlvMBXQcitgsFUm2liyPQb7c4y/2K2vWKhhB1zjb2
D48aZS2oKQjDgNdeZZaHJRcoJo6J4N6OHLtt4jJfWfEjLD6XltuYmd1eYD7FfBmD
WMXh2c0VucgL7waA6UY+WuvYx7cjBTONwIYIX7523+gT4dsh8YnIukjezyVw0UWT
O0mVITKPZS/tbi6nStteQm2ObwMFFOBePz0u9SNOWVWPS70Fr23/YVxa/ehigcuz
8DkotyLd1uEqctluDg8UZowNHvl9aPQTtU5OXwagsY65o/bqe0zEMH9AGbmIzT6l
b/mkS/amyH78OejRpoXm9PV+fh2IF3dvT46u4XLdO6kkt5wvk2A0kGe6MROoTN7u
RFqt6gFUy9q49MR1Ugybi8UQUnsU6Nz/4epjsEKOLaJNHVAlB2Ya/owGStnKgER9
xC7B+QP5cYOawTH2NsYkVSvqdNQdyl4uCUqHZjieUYUZxJHse168jkrS8/vF3CMN
kBR8rIacXx0oy3562OH+0qaWM+FdcLYcW9PCWYAlFMNP5Rd/VZNSfhoNJZiMYV/Y
mkDmbw7Rmat8sdUpqv2OhA2/buIm5YfBTjwpXidUANYXyuV6hIPAXtJjxhQwVUvW
o6IVPoDh7q/DZBN8xbbA16xC9vVquTJ39ZIiyuu3HwDeeeN1sx3EEX3Fy8g7Gknc
FXOZpvDKcN2igc+NohvLFi14cbS8CChXgfwyNTkwiYUS/M0KFgYLWtJ0i+Ll6Upq
GtolkZ+DZAuLtzNHk4dlsI9iAa6LiG1v6pqiVa4ChkvUx68IIgfN8SQYcx+gxHdT
cgwEefGcPIfWFz9C3h9bZNURShvLyWTUaQd841atmoi+HPCjRxU7I84RbqXcvnN3
L4uxUoPEdg0+xCvbXGhH1s+Zrzso6vcVHAuKowoTQxKeWTxMV+r3SRCT8W+Bbesb
nIgP2Z6gZ6wZuODA8ehJ24e9nLviNb/NRkPRcMocFCjDlJtGt3v2bpK9ZpAbqjmM
OMQuXKU0Uh/HM86JUdow8bZfabE8vmq2ipI1OfL2/d4A1OXrtbl3yCm1jFXxQL2t
wZ1FPFShRWFA3PbtXJ0WdJ8wVyS+fErS+7C9d8z7ZiqUASmN2e8AUhvIFzZW5Oso
Vj95/H/MuZyAzSnPuM1pK7iitQAg0tqXjT55Ov/OCBtOiV9BvILyTwTUMvBmGTsF
jLj10/yC0ZvmUqpYuwg7sLerx5s4v6IbhuCLVnUoZxMkozqsvsQzKeIkCZwQnpTX
rdtcsn4JsPW9D9FRvKusZegCf+8lq3IlgbN6bbK9V8KTgzaVs/P65DHbuQ2cMNjB
gngUUf3IJXf+pySWsQSPCc2cmXbqSUJhZtE+HiFdzTSreRd2aqLjHTwsTpJAAfn3
th335cBB/OSBgko3M/Nv2W7SkFnIz8UdZW3XCMg7eECf4XKo1I0aArYhGFt1qHsA
dbwLNxwslVjgqypHyScgbrQlfwkhSOZnK4VNI/1hFJyciH4bRAL4tCCdMkFwegqO
Uy3luXzOfWkjJWsMiCwV3D2c+T6FX1dZ85LOYSIX0OdiXPyv4oOy0i1x4dDrvKLx
hyr0dZUgn+zLMX4Hqb/AMm3jf8VtRdZrTkIQzFS6VbehUZCQuVYeYRt4EzBdPdGs
J2l2RpvBg08XLSaCGVXZ5Ku6T+u8J59xt2dmBbSpX9ZQVoPSGD+UeRbfG2je2zuE
OxTUiu1xFbqGJyII6ICisQ8cS0PPFe6cOZTWjGSz6g6arF7ENjJYhacYaOlYSLhh
jMVP5X/v+9E2XKkePzXeFstztpRMnwt9pO5KcgSslsGpB2yMGEd4S9n9+ZsvXWYE
3lHNMmyIvwt9gq9vKgNeJAG9GkR+ZKVNskVrbHN+dTaatJpj9NFzzmjm6e8tdEGz
1y8HbpBB2/SArMy5KEFWBh6y4aS8IKY9oZ1Tgb9oi7a6l3imenA8cGA89Z2pK/vH
PGz22IuHtKj8p3VE2xc+sR03/cOZG0ZnEwMhukAjleunuFAsBqGz8NORvcS4h/2C
YGzPIF6Bt0xjkJztNCxuZMy6or52nOXDQ+qDSIRdDyCW9eHMF84SLrkKXLlMmX3A
DrTcH1NDPvknw3Rozhypeaxwl0wCi4b8RZSQY1NkNt+v56cgGfjrizjUZzr2k/ZZ
s8eLOfVXsjyUm6jFCaYl+6O0TAYXyH4Wn+Z9O/i3RN2zbLmP7Lymq9ag+vU83lrg
3q0d01pJaplQuCOtjldlS765TiHyHC7V/M82umFiV4XFWBjzs0IEnQwAx3XxczGy
3Lu589FKHlf1pSakUDXAHi5+Y25YTaO17t+2zYTzBL8DcWw1nUnUvi/LCCuFZ5QM
5oDlT5QeLqyuq3mx3H+wCq9dMIV8LX76Zc6Lv2rz432t+nJKGqoU1KPL55jMVUio
q4AzJ8dH7/s9HIKFICoFEKIk6gAX0uXH/xzyz1rtMwo+J58eakjYOVKVqFnw2n/B
CekHcpicQpUuWcLVFxoNJPZyjG3CqUhNTOzAgAQTxe70ZBz8fsYQIuAEk9HVNdvm
VLi6Noov793zp1blGzuugFnZOVawG+HTqCLtKTcngyCwF+leqAS/WOvAnY2yWFWR
ytBT7sUZojVinHBO42OtZyQBZ+YWKPHxYUJmF4M6R4Vq4nlRAW8pwvSznSXlg5g1
KRr2migRgXTkyj2fW/pdDRoCvk8Jw+aYY23U23UQktr07v/EnaHB6Qmhf8NPelC7
HcrD8PPZdp94NTXWY2UxdJ8y8rMnAO5Bb/nSRnxAtiO/UvwEHbKeMiM7J8/kg06r
4VydaEolAxydpIvTMG8iawxSC3iDsOqqJrT3tqbutPqDlJg3b5ZB5EgH2xrMqMFR
weZhJtHaeC5ED1L+pMF92ewxiIG+WsTUigEG8EJn0cFxNd5CCWexwct7LJfxmaqe
uDEykFOaKvBMJyi7bgxR58frISm0VVGRkYE8qASfoTVY3n9/ni/zG/vWmfMoYSz9
j8gX/cvFMH4h1x68Xf2qDqy5Cohot6+TcU13eABub8a52Zn3KjfrocbJ+vU7M/en
L/5dJkZ8XX9rXDEks75gVcZ/SjfNlfWDXsqpo5NEapVsqt5VAhPGVlwe3Oy8IoCu
kNVTKoMRng+x3srZYOnFPN/pHoqkXHSoSpmAZd1QS0gxQyPbYENAVgTYjFLVcL54
Yl4mWBG13l3JfpWfUBHFahUUo7w40uFy4K08hYvXJFcB1ihGmkiVToTKw6d6WPQ5
KgN55sqYebC3nIaeyOgzmsMItE8gz3gCMVPtYtZ+X/ZoX11GQnBq2O3HPsCtl9Ex
SNITkgSO99WJnr2+DghliYhQaIrpKNNVYldoDqGOIvdeDZb+dnMlHV1HFzl5P4V8
p7MKzDMt+bxU1neJCOonK4KkExsQYqomDDgNT9fhczybnp0Ya7WKMMaIQl2uhfTy
NHK/sN2kwv8h8etKdR7+vnKJCDk5otMaIfLi6ZYDQLDs1ie8bGz3cP7HLNhPPivp
An7S2umTQY2LvMy5WpN/lREkug+7s2BSo1vc0gGWFYARP+khetpas0y+Rjkax2LU
ZGjAd7pUT9EAWWsBIYLhgKEWNumFDYViia0zbaJ6EzSvk1YPaLpOvVJUDs0LYw/u
VkCVvyNPeeMcHfP0sI/DldeBAk1RwrmPwX2nPoUGF5g6XWwek4BJnKcwCPg6hfkq
VBfIGkoKn4n2PnErf+sG7X6rCov+LwgLHCWg3QMMabg7dlhqe5SmC8j2Jt8NnC83
ebj47YTjaCbbN5TFcQ+XTbDnU36ACjS+lALNjEVT1Ga6oCU8dVmNw8jWbZ526WvH
J61Fc+xj4uGahIcIdS+JXAAA+/rNX76zYap1G/DgC6MbavhvqIYoQogHrXSPFfKz
ufNoz9RURlhHc77TeQwHKXTPxSZaS1Mv7m+xfMn43Vt2h3WbXlDuek/h2AQOmF4V
nsJrc2uCxtSiLNhxMVvlzT387PLBC7FVMoNc5mY5kZiZVkiKi6+7ixDszPdyrJSN
HKNGlqJ258RsH7IxZSVMbPtQXIGM/q4QO8rTA6/pX+cEI6UncNRRobLuDEmXrOaz
ONbHwqi7ATtfKhfFEok6WUkc1ndA8cSqB4cpR3P6mi3EYbYbq2Km5ugF2aZpNrd/
mZUgSiTQYuuKcfY4lJCnFRHji2E9rjLnCrwdcNION55ikm58KoKT/WeH0v/zLPWv
u+kcFHuglQd+RxkhLyLB8jZmwHtGu6S3mGe6va+jkPc/KSZwrBELXQjS5UaiC+kM
r7ZMgycirSz6lEDAKd1/yJZ+yHQ91PpTzZaKUijdV+d8KwBVDU7JRAZKAMMzh57W
UpriDckq/ELITfq4GTPH24Cv2j+1AUNxRt+Y0SnYNTtWNlUSmAD0yUqyKsI/qJUd
c3/vDwlDXqbsehmHSj9XvgVSOSD5JWKRZ44/A71y8VtM+sIL3xIJyMuDA9js0sf5
JHwhefp0YQ0enqm4DfniGuIoWQTDoA3ccr2eiYHOM20iW8a751qh6x3MGf+MC31x
jBzrv0+BIXxoaJpTxXgaNd/lU0oyn0pwWwVwl1H/dA4htbejrqnz5+m0Le7L7IiD
nD5lJKgw5TjSR/Lz3dtFOlVfpolqr2ld9raaEcbIp3gbtK0rQb0Cj2UY6VRfPN15
KwYB/8nYt4REwwD0GpvRM+qajQTS9mtsUipmrD9TSIfe1BgQWL52+aJLRWRwo0J5
23NDtlnYoctbXGkR58tWunKFn4CU/3wq80i/ytdxAWAbheou98QxjX5H32VoBZaO
rRvts98CYh9V/O6+IcEZ1iarMatZac5EvzuR2zw0EEXpCey8UdlIkGKPwbEemi6W
6NJlI7obw20eW+Fd6ngV4ALW6CaKs0GmSPPfD5Tno394PPKzJlCyO//Sa9pMJ8yJ
TMhk1VtcD1Ob5JP0motGEIL6meqQ2LeBVKYGtGN5uKdeE2yrQfbxFsP3foly2ws4
ncRpK+ZngTQbQosrudJxAaYPNYeVDxXeswqP04tAjsGyi1dQaB0wlafYK9bYxrv1
TtIimohTe9IzZdMPq6Na2WwpWTTTluFuDu6z1kYP3ZHNa8IqZvZ8yy3PdPgrZgy7
I9a72uw2Q61mg6lZF4Hsghxj2fek+xoW7vlF4AwMaDXOvdfzL7K36oi8sPMo5aJh
66auWrdk9m7v3cOWKyWs2oKVEGkTvMXR4UR/tl8hSBsdKZd0p3OhURCxDLHrDHxP
69U6iIN9swRMt3tew4UgErfyQVZko0L+rw5NA9SOukaxNBJnWqn4Zq0g05LLMFgT
HJGNzzK9J2W1Hs5CklNasc+Sx3oCKX+oKQYcsttAwZZLK/UjrBKJNi6bFRCbP8V5
2TqhrX/kGrmSAYGEB2B4ydXPfTV8o8i6aKj13g2fm6F7SAARqK+OjA2IRsLN9xtC
u7gMLeqXd5SXAMpkUowrDyhP6BqMz24PdKXJymbrHeUZKeuK9ltB7tNGLxRgPvdq
mPhktuwRHGEiVUn/T60pjF0ssaUHgXFab5HSp6/OTs4QK6XWA8XV0NvPTWvJWDkW
67Ihw4ANJJ3ZI4DHkrDPhlYrL9LxndTeR+KhiCtyFSVyMC5D4BMg1iz9QiIZDkWb
qL5M31+hOwMoWJaieARwmYQIcRXXW+BVNxkDaOb9Vc9i/c4JCRvSjLOIoZ3HB7Ei
ZvQdOxyFmx0+iSKnUz0CrfYbKtM9rkM0SU9j5Li8gEQ8MvQ/iRq29cAbtKTGhARJ
CMW9Q54GtPN163RwdAHFqNVm5eCq3RzNiUgvzwtZD5tLBD7Uk3pG3XNp10sEiuo/
rCr78iM9IUFFtb+t6NG6H60s76IOE90mjoU8+8TIhMsbk2IWDdp7o+p3BKNrjsqL
sHrJlFgME8ykNJ4SKp+1lCFRo3ug2YGtV68YBfdV5KUX72bR+6RsJ2lP8yV8WIC9
pyWCTcsd4REWHXMkvrR/jmFFvt1kTJ/rc8RmPD7Si0/GaQ4FFPJ0geOqVlm/BIkI
w2XjUAR0g88HgTADP4WIAkrVfsS8DrBHH6DV9GEjqvPBmqPGvQiOyhwWrZPA+LoD
/C6DoQh7Hgqu6arBhH6jLg4jb3DsDyZy/lSsl2m9GHgWqnsCPrbVxkobP6U3crBT
4BylJUlrL/NIW754/uPsEB2kS/jHZ6GSbE637lRVrm0MWJhS9HABHsFXGbgzBohH
hTP6cOsF37nRM9CYqgKJ8IN7NVJV6l77EP8D/7OdcHtgLkEHDsslqPp5gQZW72sn
yJoaSEVxskuEXeVuU6TcTJvkceMzdbr/Iu1CH5/nx5aTlE6jfgsNBAVA01/j4TTy
lHK+2UitiKLkAl/JDAkcMteJ/IzxY3oCwImqggSwKz5sCHVBVP2qV3tQoVcOEqt8
8DZBdQ1I8EUnBxlz8gXfw7QUdZRgpd6ck2zPHIWyJpGJLeECeuO9qyc7c3mdjmnQ
nKc42Jg/RzIxWJtqHc5mr8UPB/XkaU7XVL+CNNF+Hx0eyHjasT2AgBqyDTGKzpey
Pkk3W77GZxvFBC6tY++NnxKbbglMF/+7e+Cz3/1CIPI6Hqk4pqASMhe2bXuYHlfO
/apdvc8hlfiw81DJGJ/vNfHsRxXnw2BW4JlnSP6z3HFvTuLZMhVo5rSdu9HWFHR6
ahx5d0BsGf9FvdixHE4qXWoiWMvqSIRSPUg7+/XAQrl+GtmSX/KQX+k0Jhx5yAyh
ylUiDDUnxmlc6gWbfa64tgRTDqyzjGj6d3zjA0+KS54B8a1alwTgXk9+xu8fcoAd
83HYZsffexR2Dyy1xf5gMc2K5UnaxxFKI5BsXP0VMiDDVHYfJNhFySG3s7+KSIt3
PSgCpYW1aR1E0tQhdE2D4Ul+GGUzzKM6OHg2PpG2HtdCYPykJF6oeQEDPMIMMpbC
Bdg3r8/77xf6IraDVVNR9vvqtxD/ic8dRsMCL1OeDTLt4zcquN5NTxQtt+qgNWSJ
/luEBDzj9IXiV2qZIIa4oEEL4d/THQTEgjWm3eMHdo/hyynRYmnifbxY44VVtYnJ
6DKrAB9VRJbdR3jD3yvXhwcn479YX7qwTtz9a8TYv/D7rL6TqfQNCwvhiMmsHJ4Y
baXS0sDdsg1ACRSnkZvgFZsAqOWC6YSqdm6aXPOsLjD57UkUONHk84ZNgUPxaKDP
q27SO0ZZTLMmOs5Xl4FiJYgKzTD/M3yi87fMs7gDjEmJU8ZAKlZoqXpcnD4ZdDrI
8EqIENcmz3Gn0hxj/BqX1H5TH9VhdmMI/KjCtO0ELmCP+BCTQSeZeeKd4CfobBKs
891hgt/8g0ARYF+WRSeQj87Owqj5XNK1uZ7Gh6I1I5Jrr0+iQ3OhuylYbO87hGlH
asZCFGOO/4/5Rif4MJi8LFPFQAejVuRYGwa9Eq6ISIGpDUUeOZbQhEIJagp+MyGp
oCjq/khYNxi7rHTRc8XZN8m5NrePDQvjwbYuzuFf20Xumhnbv3Ckcf4ya/VwaERq
LIbml7ItHIOWbdBIs2m/d6b2u89j7iY95oStkqFnYqDe5EpQ1cmSacEYEtqn9YpT
wQIbFrBIg4c5PMqLu5zYC2fMX/CzJmONABB++xsjuzB7OCVjibMhhol1OjKKF5b5
EfJRHnQP7VhnIMEOt5oPfL2hla/d8u/dj+cKxRo8U0PL2HHMshmk7Wyna0JjDNwD
ZCX/nTYcx/5QMJoY10oUY4Rsoe7SK4uyBIdQaWzViUcXpmmrDfPn8ZkcIvh12spA
axw16tBlm96RPPrhiaD9MMX2TXNseXt52sf/DAhODBRskzFX1YX5gYtocryWFNT5
j1JRsOo/De+18l8iHQGC8ElkDLLAVd0mpV1nE2JzXyUOSXXZyxNYaKZRDYZSqZ3T
jUFN+0u6pPI9LO+WRiLp0aVHJJ5a071m4tbVB6UmzqN/i38k5Bdg9NAlVyYqp3VY
w8pRQFZYrWJzV5+HDU/20ix6UopTkS1FL5kdf82sg414A92c/ddN+uCv9ddp5pi2
nXgjADbx5x/8HnmGYnpOC8tVik4/uxOYh9fR3C+xIc1heo/Hlh4+QpaEcZyQa13K
5E5GxV576Hl6izrm4RlMClugtOKxFQksPP7kzjPKl2N4NPw4Gqd0q/kk2wtwsnby
NdufytdgGXPfPVr9mnZ9KVXr+xhMB7UY8NHvrbWnN8j9exBfQeCzTit+zxRH3ZxG
+BjOxaf+z7dBeNrsDebiWAILhxkd7SZkJrxazBDlhWR4EKWnd39q3ZJVVCHp0TMN
ewAukpuSDuri9NOM8ef7cO9OmEln0YiY1eMPhc87wShTWyeEvtUEb02zLjhFlnKR
ReTEnDstn2uZUPUkv+wRKsAHppGCRq4mC4pdH2bP8mVoeS4VWGL23ufc7vHg1J/B
k60uX/u9+62K0jAv2sGQxC7bnjQsvn1BNzqQq2MTbMfNHW1v+00WR819gH29akv4
kfvfG0SfdHrzJeEJSRxitzp5QaNRGidRnjedmfLkm1BiLpIcVKN4Oy0VezftDvUA
d5Tpz4AnBVTDXE0SDxupyNws7yaasisR0b2zJv+9dyxgVvewCRzxDCl6QGMSU2iU
Y0ySezzTbkaVRkJaErzEotUP9r6fKX693agatwN3P70jgqPK0rG53SOwzSvyFBD0
Q4MkQpsInv/DdKTDSRZ5/FO+PlCWqCfxwUxeX15eRv7Jx2t95n1nl8oaFUk+ty+E
1xtUujSmpvM5fuFyQJZyPXf2PEs6TRflKi7QGOCCHgdYhR44rCfDcmygZnuZ8fgX
3XVizNEtNshrKp+QxhJkdcptH3J5yWUZmWuqRWkdPwKPI1DOazTyfCiX0T+00TPi
6ymconOiWSiSDnIIkRhEMUdftiZscGMf+7YJPIJIAa3W4bxx8cigmB3gMoybLRYo
wkUVeL6W+Lh5hSKIYcjdCus0TPvUpw9I4WLwTfZ10l8UTljj8oOCoW3Zqe5JPD2W
EYEbDbF+AFrHp77YAP52Tg+ufpZkLdoIIGBRsB6AMKpxiQZ4i4jdqAdBLZcmVTHh
Dch+boQeF6Ys1roXt31ai3qsj4AIUl984TEOCUUgzJqgVyjFxqB70yQXfYrRHE/E
pbY2wgkRGrFOGhNCLyRM4QPfuHDELWbavqeXhPv+GurgwCPt+2RliIyh2KbvCo1L
+dQ6Z+XzXpBZxBqPOUGJogXpSwVpeX8k/zMTswBxGjd/g/oAG89i6a7ZloVNPHPa
YjTh1XdJfQ/QIGW7qT6ZbEtCMtLl7Tu35BhoRfTlgjKSMSTNfPlA9V2rDbEAeEnY
8qPuQjq1QHedr0K8mfHLFdvAF1SDVUgV/F702iPSaU6Go0wJB+s12A0lgUAgV95d
WWMIyK8WnYLP9dt2jzoz7N+58HgIEmj8HUNvy6gMFFiPIxECaIZ0mziGYEzi7mbf
gbEzErmtsvU6f24r8gO28KRb8JkVlfhUS1K2k0WmPLTe3rIMF7hyvnYG+4QPg1HQ
Y1yiA0vkL53rV1qmHuSJvrjvLk+jPn7Krfm8Il0QZxq3QcTJTfRY7UpQFL2tixul
5aOUgdTjzaraO6VqH6FGuQfbp+weyiQf7VXkjopIwtW6eNhBisYZP7ny3Vns4C+J
Zoyb56LcE1c5aS6VG+vHpm5uoXm3Lx51r5yz25damIslx5TjNFBvW77TDN7jiQbg
v/iQYaZzzsNcUHQx48WS+yPf4RYlZy5dOR+TEcZQIAOF0I8kumSC8VU8GKSITAFQ
+03x364WzVJwpdlQJ3HU3yaHdcSxpvGP5KEotybHF34jmeTxA5xieDD4ba13B29L
LhTIM7fFC+KcuU1XQF8dQ+MzqvQqdpkmWTZhUJhvCILTf1+F5SEb3PhoF03o8TRU
cEPOyP/VMACfGLIWuG8Pyv/dtZjI60oU4MhzPCapeLVM81nUeps2zmxvWTZZmXhZ
urnbRUk1BxUUZRYgNYM9WXeSp8tW/kvyod1tHbnFlm8rvDShc7rE11JjidxYP5lm
cJs3yCmPutCP2GKjjBlDp501FzSrbfEFFgPDpgGo76Z+la4z7kHGbHr+bElZ6jHm
RFkQ1Oonf4IT7Lc8cPY/HbUy/HoXnqLXa8rVhWofBUqXFlrCpYotWM8gWX8h++2Z
rhVd2vZ/Qv/NplRAqK42GWBIhpWe0nzj1gXQRwQht2NPrh4F2/v1mcLitwKAaied
fHklJ5PFMfwTe0Ywy/yKHrnNxgGI3Nf8ZBqva6eH7LvOPSg3kbs0iGtx5gm2pOEq
1qX/nuAhJPJFhyxHObReF9kjRxLVDCYFkOcykqn7yznSLEKw0TXQZvciArxxpZay
dVrTNAvVTTE468bgOV8m9truoUvP8n52ETxARp8jKhFbN/3DX29lnoIifkd2wZ7F
iMiRJnV9UrbtTY9CdU0ppC10q2bjNgeVktF9N8QML1QXhvCs039I6rkqFmnecFyG
QyP8mHPMoish+WKSNJYVK13kVWcbUvwcqP3Cn4Hq2MI67DBak1MfpecT0GYt0HyV
HgHNmlyNEEcoYSPEatdFnuO5Wq0W/zXQE5H0nOROgB9mHvJa9uWmEEzC7t/+m8gJ
IxHohOTyrMHXeKag+/YRr1QIBRiMr9Zw+1HVKnUHGbgToWTyLzbZuTo3lu+MEZgX
OULel+hB8nWRs5zk6AiyTBN7wdokf1LWoFS5xFP4/NvZM2rry6FM7JkLJa/eOI3u
LOoYmz0VFn9q9ypcf7Ixe6Ug7B4mQPwpC1Yrgmarfz64SH32CtF6REQKRg3yTUaA
xD8/dsg2MVNPVEEfkIsWx61ZQLHDtH63OTDiGE9YrUmeEIlf9zB137YEGUpYGRFj
PbOY8kUe5HsOSxzP+DeUwYMynivLQ+BKjOz0t50+VAQ0H2eDXZz/mCcwiU1R6JCM
VBhFT2NGIYefXBvUtl1UM3zmh/4wWV09l04gBPa09TJN1fM4bS/YHMI+u0lw+fD+
vwF3Q1+0sw7Q10xwi4muF1Nj/s00CkXIuaavxw0XekNONkTCp1nouKgwMe2O+a9Z
za4IUQPVbE3bNiua+KVaJ64OAe0CZUyMCTkne/p7heRnO2nfP5WyfnyhwJO86tfd
qqKBBeiyQRdiTWNQy+w4z4YwSrTdB62C9GL1mih0Scqy43VgOVSIgWRaoJAwwIYI
eVUNULhRoRxGXczJozSuCJfagSJ0b9chpCgVKYTowAxSW9wWrVJswhs+Dj6ZvGAJ
pCssVTEUIaTd3X5ekNC7DlH+A0EpPD7ncJ3OlHhguNjeezI1ATFCcAaLY2FYwNN5
SK0/P1ytPWIRBCbS+PYKKJovdfheV47fFaYMXR6prI6/Q9zWnE9t86CKcoAxV1dC
Pt8stqrgHnxkCwXOq38vbyA7KtIOOJisobKs/Z3S/u8OyE9Nk7PAeJ7HCmSaMoAz
yyRdGEnLVoKJk8NIvuVV85e616q1ZBszm6RZOrWOtd+RAkoqTZ4z0FUwXnjCLv3M
uiN1k0dFRFkhQGGQTN2n/drTpvJLyKqLBj9ILDQ5XU8uaFgnx/DEq1YYi+N3O87S
sT65zk4L9tw/rb7ja05YYRrK118owG+SdCokzxtvEMiZu6w3c444sqCtrcKWpmYm
flYzmgW+Mt9BkNdbpghNXD4FcTk+QUFO8cemOMCrGZIO8xxQpBdGhjaEvIAOrre6
IO7MuomS4n7kwDqJRSEOSJEptZgI3yt8MUfTqeFvMraH40Ieb1KDpKKKRaBCjeAv
aSIcfPFBwqkV+hOWtvTHyWYo5wPUOjk8PPL76oIp+euA+CgtV/o8GrH0ogxWWckA
AR0XdvUEG0riSqVeRvYnv+x4ieVFirBQHCRcwJUZKtgQuAyTJG5lXSNF3z2r4YWW
OLcQelNvCZdmG9yz6RRNpVrslJNQ2mlJFhVopMbmjPoPMXxCoqR9uOakJpsV5h1Z
zdmnd6aLwq2YaCd9vZh5GwvVGeghJbD11iadfJG2BUeBHH8YdcXJi6SFFX/E5bC+
E2WF/FdDSkqJRV75zvazS2qiaOE9Xt8RlGwywNvE+PWJyJOiIVb4ADVaD1if0HLM
zSHo1x4yW97Yf/iyYje+lvXcT8lSrP3JY2fOsi5BJabjfS7YMoShHPdfk5+2ejcV
Un7pfKJXzFVMeSju4pToulddBTDO03gGenDn+Yplewv9iqhAgTmARzSDfl/nS73h
LIhr7/UbSyd8gbUPAhTbiJBgb6om+hy3gDcsTewdmJw++wRrax9pKp1PyJg8jdHk
sHjKsNxvmgXfsRvxUbdQNb70E3rkkedfXU/pwVbeVOp6iyYub4V3odWp4MSv5z5l
0jwJpCIjEEJ/QOldQWrv2YjU4tXOEseyw1b7HO+IKYznTYWTBWyYEvyob6kFCnUT
xzXbVwUq6aXoENkFyYQaFVB/Tyn1qFubIqUW31gp01fU/H30iKl/c6k4tr/sfwQY
mAaWH8setvmv4+v9AZFs3l5dl8lbMTj9EhuY0MOg6gIEqmf4vA1/shtcOwuOnnus
usVEZn4CROZ8GBtEqqaEqxQ1r71rOM4vsyu4E4jAz1+6Ehwgao5i20GsTl4JpyxG
ox4jJUo6ihxB+0+KFbm4b05BFRaxNdwH4N1mTuc/h1FOMxI2N/oYOzEuvWzXlKo2
1ETK7NgwLYJyKQk5JtpppNjr/iqKyyXYQJ7pKkAnGHqquhuWchh9Hj3aqO5JT162
Sbg+sHm5/ZTnjGUqQtZWOrbVE6t/h4i5YNJMLqiYsHiXgNh4i2et2wrjeGl7bOUE
F0Jbc5/FHTUpHUwt4rMk16TJeVo5ZzJ1373lFM/tfFU4GRnwxMvpHNXHNkNQLlp/
skwfn9ZsqmthnRpvp20/VUUvLFLvapIQL47hK3xTRXqE9GTYK4Sl3Da5cngby9mS
Omj6dSeNj2dGFhNsyq3CJBAhz4t8Q4qVvzz07SSQqJf0MKPp1pWEoDpid6HRcm7f
0iuCHk9PKhLdKDtYNZiZ3YtfmC8XHD1fWudlMNF5TZ9YoKaZFId0hBzrYGj25A6z
R0T5ykivx+D6ZF+DRNglKW48br6uwObOQ+0U8LZ3hR7Vp4W8PKyTxwKaVo85DqIv
gFzUhZTdEiXgFnfKb04G1IW8xGtRL5pe/3MwHtfp3HqEO7k6F96lNuim34cmc/nE
g1pyT68vTR/X0KmdFRKIqs+qjqoJ5YcqxD/46lUKH0ulLaA7zGqWH4QlovMZG+uM
eg1xC1aKEDALenhBH/QDawptfRvv33Tw+p/IulhbmfWO9rp1pWJi5mL8MwpchGyf
hLcKDBNzIWQ4vq0jsh6hzpbKmGgnwIkqekfBP/qw9KuArby/JK9uOUao0WrZ1qU+
bgo9xH387FzoX5pbwLvo6kwlST8lHCJjuHeOPSELscl78aBiNqhspE7U4/KzR7+l
KbSwk1zQZoblL6cO1EWHaI+3tcuiIFc2Psovtnjd7QkDOt1Aw0XZOcxfPLGe6Nq6
ZyPlFKU4ZahfhWvZz2Wy0P23gLIkJK1NXPbxgu5yuTx66am+SBU4o8JkamiZGYGR
Gw52jfv+ICKBzeqQAavBSA5rMug1+0AvTSfplQPzOCvyVVZC9djeKDNOGqJxT4ad
b6uK764534dt6jL4yPToI0J7k7P+xX61Ji8FheKs6ZiPK6ywkp6ErmLh90ahLgcF
Ovsnf40eEbXW+c59YWIqr3tJZxhbMMSCV8xlppCclMcH43RyF7gDQkilObVpRaG5
Yk5ZpJ90BVNHn9GLdTFdAbgNYii1roZirkIuMp5NliYzDoBr7760f1IrQljhD2eS
yC4dC4GsivqG6VxLwTvWxGeKGsxHAGfIEMTW24cWMqBAfKEyV1Llo/7RcgCcO3Zs
AQeN4ptI1h/2U2Ihv1Bo2geLL+yXenMO1Tf+7fPB/GNIhBWp1QkNcY/UrxkBvZLT
EcK9ySL1m/fmfnLkwdRGEjDWAXf0daRl4gGRUdsaQf2yaCWHJQQfu6Rk51knEh6E
cgUd79lZElspwJUs/xOVnvTWjMDatD5JKcWIdQUZ9gbMFcsYUBcS2VO5QxuyoFTq
uuCi7ExgEm8aDEDNEsPPOSDlM7Wg8AbXI8ydj/eQbhikHw3OnLCrX1fptA4X0OS5
ZbM16+Is3roxioawMDuuL2URQmrPHYQIiUFyNgwBdExnOAVgjhDBdgP4jDHOabkb
m32UWCJvuagbUN7tOB4dXuZ0142dqtM9r95LtKh7bKvpj+70zvaPeytoYzMqtZ/e
61U0aY1kCAAp9bBf73jsyjdOQ6Ep3ijAwETYW6047ENVgq2lKA1+4t6ypYspbeUL
q+qy1XeM9HUPlngPnAeKsWUREEGf7L3sJ+CkuDGso7+aS+CWVUQG819RoVyzlR+D
pbNeEVhvfNf44T2i+Cd6AmL16nHpg2yxJIIjNNDfy7NH3JX9hN9pTyrFyAXMurrQ
//gwgEaSDf3o8K8kl48nqhb+6gGmSVfR3OKYFaGnKwbAzgMchVqOHy4cgBEgIER7
uzOnEBhvFseG0FuyV6xEJcNaXIh41gvY9aF1w+BifiemTM6Bf5MzSIMPfAAG/9bf
JDnTAONDuaURt63/rJt97cZavBq1espA7R9V8w9kYCWWoWiGireZ5kxYyhaYY8QW
FIeWXpjkeOxQt5cbRR/LYE6EnJqjotLst/vji3yO8TtTB52vShcTte0N2NA5lSIF
W8yFOO09AeTuOan9jz4bO/8dp+Yj+3eUbGIGOH2M1XXLkOJC2MwMLKquid1zTUhJ
cvvkk7j4OJSUz4VjrfL+g+GvvQ4+QkOyIDHTE32/O9VogrZzxdGW+M+UKkkg7961
nAynRB38asCcRuk0za+U4PAMiwStHlDM2hBkoePiJkiqcisQ4ls0PwJf+1hBV1h3
QpynIwBuf4JaPCobqhPAHxqA1bNPiHSjrQgKGQx6ivdizQ13F4/GH4d+7NgKoQn4
ntQ2V9ofnKtLvR5+vYKUzSnVx8iG0SYM4Pd9oPRCh6svLjzSiI84XdRGe7oypS4p
32HAHz6Tb95XBgt+MnpXdXO/aCd6/3D7eIR/NtY3spEaoLv2cAfVdaMEXK5bOHUd
af/qM+hfy2yV0QNhZeNDLhWgjZgKm/scA+y7T0CLJkNFERdOceyWcNfii0G/wbjJ
Ot/3tiesreUHDjha8/UKVKEQJ19DXPphTVCAd3tD9t1zap7TxTLz3+jn7UZY+HLg
dvNeNbnN66KwYTZnrMjrEIBKcJuBYn2zgmDeH9TIcmU/vTFFLT28DqSy9IyfkrsC
CpTniChFharLC2fiTKuy6few7jZ79q8GCphELedJJHvMRkRNjtuN68T9qg+FnDYp
nIfrzBzmkc7ButtNxXfLfw2wTd7J+pVXxpjL92fvL6cdRs8s9sttlRsNXjTJMgMs
jVnUvFCwXIoeQ+OzQxxsvyJDx7+t+4+O6w4E8G3IjtmjDiVDi3Brg3ns7W8Qu1IA
67ne/FI0JhBaFSfOwlWsG8EI3kkBglnhrwiE0K7xU+OzUHRxTp08S0WQgKqlBC1x
2Wwzg4fvXpPly32xzh4N418b7TjIOVIiqZucYQL4u6pOg2VqQRT0vwy7AFi/mlVK
O7kybsdtE99J3d++o4qYY/tQ+rlZ3nV6yKNAVRvgmdAHF2BW84iSJNNl1EvWyFbr
+Ey0MVdht+NRUTX6zyjgBbecmOyudWJvoV/HQpsqUuLirCGNS6JDqMWtXhtie8Wy
UWDmou78JpQBiJTXlNMmTq19f6PKLjxtoLK8VBtwZWNa86gRNKVP2arRM0OD+b0X
kfifM9koMXDWu0FLYB1sYg1flaEuTwJ8UTHALBpnhYlz4AcO5FVwuIHtuqO4hCni
FjYNpe8ptbG/xrrITWN07FXxHvRvPVjBeCdJdGzzoBtCANPbdmHwSUPUBwMybIHK
qRSJ09ChwjPWLeGP3RSfybciH23MA3vDUfWUk18lT2+/iS2hp8EugsYd0ftJRjki
bAz/yOXgoIag3k9bxcwga6k8W2SF4+DF11WnASlaTl/2nOu3iRsk1JfK/+qZbDLQ
meEOsm0VTY3UF1RgYfk1/QL+2wo1djmA1rTL9GwKH+NYf1Ddtak4jOtHJvhz3xMh
VHW3tDQ9vQe2rtLZTg5VKk7VEgrVf5ECpII93N5nUi8rJkXGrGgr/aFYW0Ab8mCO
Ff9V2hx34gDomyi2YMz/s9lejeOmm4xvIOYU3J6adMH0g+F8rbwFAXp+1TU7Dvw7
C+x5L20Isj9MetXRGp8ovglwMyOInEyaAfRLF4E+nZNWHEFif8a56Pwv2EnEX+tr
OGthABOjYVzla+aC+AQqWedV0J17krQ9sr3O2rpvRVItrm1LuRatPLYQuuMi9DJI
b/9aN+xN/zMwK96XLrRrOwiTEVDnk0y8A/JfZj08aIGp3+hTmqDUnLdilB1q/Sp+
GA4WCRfePSCjZxJQ85u5eRCSHTMY7PuXniwsPRqmvvIge1Z2d6EjIkkpFnfKtLfB
Z4pRYYxzhnv63Uv/Tk5pXKH6KB4/89ErKkAnO4JW5ZINzMLBi+NBYhODteKGVqe9
Sl9klB14bwWngQTR33CfuvWE1Q+XQ0tgYkL8uzuraP1b4vtpI7sHeu22MMsXwi7N
YxM8q+/V6bVXVWwH1KUzdl+4CaonpUEwGcMGQc8vnK2gi3+VPWt854x+OOQ09/r3
wVfFDEjKOq4mha4t3WR9sdx8bKcMzJBmCfY6TaqHONiXk288SnitGkCnvY/b3TyQ
BRsyUta/pCzSwDG2sNCAYLVXJrWcrFtNbY3FhODXU30uap5PzlFYKlaqwQ0fFL8w
TtSS06O0MoadfT1iN8qxxd31vJ7/OGdGuVch9/WN6+mRtkb0/TV7LNZzyrncxBnb
NRPq+JguoVWfKihvrkbb8shK4tTO6spgsBHPxMCE4jnM7915vtEFS3LNknZChMHt
OLQnEl3uBd0cZYndWe788cKazbkEmwV4PpG2K39JrbfW88mXiBZLAL1UVT/WO8HO
Q1KEkiL1olPtC+uenRsMc+oXEA2OuXXbqNt78bbySnyPb4lQ0U90arDqwzPa6yk7
YDg+eWlygXat02oSmKiBEMwWQMujlRZ57F5SIFVUtyvvMvIlQvWGDVFap85VE3yE
x6V7OgeRBqGdVAmK4hyps/boyJIovvZ81QLCjbBc/hsRHiOxcxc4EfW325SldFvt
ibs1j4uNZ+QCuNC33haBF8TVolEjcfv+jLal9YyIE3AmU2T+uyUfeSinQ+4iB6Cl
APY7FsaUXhi69SwdIrWtW9EG9xM3IbF1h4ZZ6SSjO26ORPcsiohXXw87hGGDKpK7
wZvCf9IUc8SGkGKomTnQh35E3uWubJErlvRov9arOiCc/KSKunzMI5ssxQtGF2sk
HhgE+lTL6JKQrEkYbsIOvhO4FzQnEDIAk5QcM/6AL4aZYM3DRpHWgJwa9HBdLpjo
sGZ0F1OzB2B58vIcAsxjWhsgGw8OBL6uihsWCMsTd9yKF59FYjKZJ3dnrdyOsFgo
EINp88z3VvAzQFpCtHE9NN+YAhrID1ZQGFwt5+PS4yQJkHW9CAWmSaKyGIWJipc9
UeMjw+eqbDzzY3TAOsJDcDBYO+Wvsx2Cucvz1gHibgaKhBovhsTlKyKdwjeH6kc8
UcjvMhYGU2nideskHsGGrx9mwyQlE6L2gsgb6hgqQYJtX4WghRp4aequeSdoCmUK
9LfNJdebeWkbMgT7j/5dv63qWKD7cNpu0x2iqCEViIs0jT6L6H0VEqEobrqaETLI
DF9LRObE4i+Z8fEskVq5RmmSoykg2u2UocpL00X5bRWBJoOFtJya2GnlDQ9akRUi
TrbnBVD+0AtfLJq0lLBiNMoZ4yukqns2wK79UXK6c1AmsHypNXetjiB/hKKMv7zo
KGk5vl1fVqwDFIruzvxDU2rNT7wIzXiqyB60Ea1i7j9zXh7hJVjkrcFqyWgfnkbT
fTsPyfmnxJ3+9VeKia3fL/oJxkt/6QU96ml+N+zZJMtYPuLrbifJOQu4l76n+rH0
36NmCgznmxndMb+hoJXr8vntGC0hGYCnm/QGFRpHBfKJBgJ1KrW3WBzCgoOwnsgk
7m9e26V8CgQv9G6VCHANCEMvyxUfTtuMN4tudMfMvgmo57o83K7za/QOHbPrnJs3
cutGUDjcB6lG3PSoTxXzkBLzQd5F8znS+5tfMzw62zr37y0N7wMFPC1bg+4/5CoD
LAIdrhgKSqymcil3UE0TjqGlUoTVu4vhvHXZyGFh5YShW+dIWHYMtP+Fo/RnV4ub
ULMklnSaO+Cl/uUJFJSJGcXJS1a8qQ1XJAqeQgIwqdHEPPiTMHnOVl9Av7Dvral2
o74IbtfMnwtjfOuNAufY0V5MsntEocN4/1GopHrkjTQBkat8YRn0XV9J1HD4GvpS
TRZ8pPC6NhR+gLKB1aB69kftvtiZUMfyfwaQdrksBcPIwPKjPrG1d/rwXmvotmZY
J7j50NQjZi3/KuK7X7Ulo1cmwerHjnaTWJn049N/6ds3jbtz/h/fmnelJ654f88D
2JcQjg7/AXZMvgeibRsPBYUU8EYjcGySkNdwZvvR9ZZJ6hReFBMuf2BY6EwncZL4
26bPlKs4SPaLZ9XMFWPvrYpbneFCbaWRrZ8mZBOO1yAREWcyyqVb9c1+s8G+DpCE
JfrsJ7rPnEIY0BR0MgxYXbeYXmkyNjKJVElwlbIvS8QfzXiDl/B+eE9mjBRbyr5F
TtI7J289sRSt1NVkjbpuxL0grLtiSj/SxPjvhgTfChW308F8faxUk/acQgcYU6Xm
s8WvgYUCt7c33fy6cAs7DEpFiI42Ol0MIpQzZPgitAnxRWN32b5lrzYepg2NRqCf
36t2JrfjweQeWABwt2hkifMHdanshb/8eR977ogX868DYAIvakkKmE2QZKfexxcJ
6T5Qb+FQUvOssNXUOvQgYdQf5XszQWNSth7/oygO2cPTIET5csZcPHaxm/rona3N
N/2xJ1v4pVjmMlwmZYnzTRk0E0m3PBY/ON06iDuy2P3ba2AtAFr9L/XHlW0MU3cH
/e2PapG3vMH4/coMlvWdfe5HNhMCJcHms915r7DJr3+SWcaUZu2a3io+Oxih7PaU
zX+/o0PNd7S/avBOYgiusQ7a0oV5BvdNaWnPjM6Vwsk/G5g1ORCpMWpsImO8LCO5
oCtAUFtMFdWu7cHrLwac+AZW+WO3yYKU0ASb550kang8IvSutx6ZOo/qCg2w+6KO
I7EkCh16YY3DQncwXWk2xeXfJ1zVOX8WrbL54rvjEgOJRphjw9o1Htu5o/9mevJZ
g7V4nSCnKCc3srD0hpYhrgcAeZnC+6xiEV0GZ1TxIKadeWCtr/LkZWGTWmZXCta8
va4EXyKFCAMDG6nuI4M/nRTpyJtRbG/EjB1t+ZGNevGkYqadrDdIy/irJhijG9ep
h9i3XHdSb86vBddXtV330aOKn/eDP/mQg7Q3c+XiR1UqlhO5ipfVgP3bXH36JiKD
rP1tHlgaZ+uzgZ0Ro80Mf4SeR+NptPahRzZmDC3JkV4zGdlHAYDQWcjkCF04kwmq
+71/uDShZP69bGDfpkSJDusfIVPViUUzrlgebjtEEcpsNraulkWr489f7Y5/rEe+
OG6QgcDd+iiuAi3JXpUfkerwltrm8aAdT+DTniyFr3S5qG6WFqD/gbEp12rxuG0F
a+iJSAp7W4DD7G73K+BaETsLMesrbXgUrn2t5GJILuvstkn1YhddEj/YpwIqNtNR
3tBR9nfbpxTpzRGzd/wSXJqBlO7UHqWKokGYaz/S4VdBFIbCh2a1Mjl/D1H48ny9
jO8mTxGMsN9HsYjwbl5Gb8RVX1TIJY7Ewf3qzcDUU+vPqUu0QqJSVA5LZsNfS9i2
Y/tbYl6b00PeEGESN8I18OJ6E+ahrJaIg1Iz+cGq+GhkD9io2ZengyXP4X7I1wR0
xN1b3k5NAut6vjhyVMC4UZ2W6gHbaOMTgMCuGw0cHAguBBNdNxtYqc5zbaQ1OTRh
tPCQ8ARxNTWPVrQQOOlq4+eFIDYB9aqRK3hU0zQMRbmoyf97AxU2MjvzPawKxZTY
OBXOvE/rkIPwvcSJ8evPOAjiTC9ZOUv7aS5W8mtTm8YaawGpnK+UyBjDwasX+shY
cLKwctcNN7OEu/3lz1g41J4lHF7Eo5vTU7ht8H3/Om6+CUB6jhegYsBK3uMtGYKn
LceE+ry5Y9EZaG9em4aG2LsGbIgWaXKXuiOxjR6lE7dgHDSEwUAbmtpCDtjzQxMa
Z3TYcIS4te/kB+StiHzOWttOfGKREJvAUPeUDAXjT7rJTcddAIie7SUndWXFeqvM
j589ZlJe2ONp7x5IiShrsz8gyj5SBi8wNgtUuh/F94ENjJB5aAvWxHPkiea8PYAB
3a9fk2WhF4m0FSYCY12qDzscJB+9jeSniqufAvVuLB7+nPjJvVT1FwrJt0mFjUWE
GaebOovKwvetz18Bd3qyPiq9D44Yp6iVHs5F0vaIKCGaleC9ofCj8KDaDsKpMSza
AfhEuKI20ucFM19sIzJho2NfH4Z1ms+d/zpnTD5kyxzQ926M0A+dSyjTKklRtx9y
83uxwrk9qtGUInwqStyAZ/XY2bNS9LQdYhbMlc+rCdoAZz2/bopGudOlNhNuL+BJ
zcDzspNeZIymwBt/F09ZIxzq8pQat5X/F2BJ4IGB9bBz82U3NVtZC4OP4L7M7Ew3
7AZktE2hRcIzF4aVdo+31zaF5CFApqnZ7xyIDml8eey6c4YEwLPnZvufC0ZdFW7A
yMmxca6OhAycaZuBzLRCAuI6x6SUK14YzWuCV1HUZE7MlAdNt0PmFob5apin8pzr
b5BdmBrgyZLRiEOQS2cCwQ5ygvZLTdmWml54oEb3y+OEGmmdj8dPvdzzGeX2Fpiv
zbF+mnU5JlyXLDe81uCSzhHDQ8ikfiecspFAdDB+S6AkkZlQ4ASzIUTqzE+TsRMB
wgErnm2kYcSXFAOltwB8Qqo/4ZtvfZUijpeOp4h9AfrTjo3DtpWayPrBtgOJu36d
Av27C86SeF35LLwd/EBECuOt+ckzB0HnB8O/TM+ZcKWlghFlqOldPbVrQqaCWj1t
CrROYoR0Yi1OQCpAkXDh0nGAWzOb6m/CxHvrKQ2+jwtGT/S1+JRAWvYrah7yCqfz
rrcpnkQpLIhJEzRpgOfD8dXPobswXpD4y2lshsAEK5s3e+ksNqHTYuNqjsRqRsmN
9u/3ItMzUwdxpCLtm0VFSMWNDjbFAM4cw9P+zyC9z632u2n/twoofSFubdbmhVty
5CbC2S65MiTR/Flo7818adWUZbnyuwPD9TY0knqY7nDrpPmDYtlLbQEQUfu9x1l1
6+cA6fGlxNL3wARcqh88Q5JUVxeuKI7GqOxlW2RizWsrDvBdhk60s/GDqLnhe9N2
E5pb9wsBWoaw8aHduuz64/RbGHiI179YH9hmsjqBmgqO4Jdx8JZjJtKvqB0DHO3v
qQRzgbuSnlWN+AlVTBIQv+oUbScLwDbo/lkJfug86R1Asty//kTccGzGpE/KBcyC
LujvTmGfAMqRjj+DRHBtb65A/WN2WTKmQN/iRw1P1ltnSBtxzlpuMxz8LO6yE2dS
hiVptKlwAI+YdC44PSiONNgkxd6MFhtE1/arJn/M4Jcg5rm2FpLjmuPb79/3mcNC
CAFdGgIaH9XTds4iJoOUBODYC3Paglelg9nFI+DGf4HpdiqMrYvbSYkt5Ne9E2Kk
FIhxgMT48fnaQbJCQDOmuVXjwtkEquQcsP2cU5LcI+cXDF6u3gWJaD0HEV2FL8dr
EZ2ZuvQgcpKs/PfFSo5yYudpf0sJ+9gjdPHxv8mxtWeJvEJrbyXuZgza0eaXP4ur
gmNKLHd8JM4KmRE91uOEQ4bxX9MgfioR0hshZXFogeDRh29+hk75tPq0MRRXZYVI
QW6YvakA44k+rJKTWknpdVot0L8HcDPLzfIaXzbnNR1WCsaOz1E5cuPO2wgr0dJU
l7vU9Tmjt7MLGElWmnPAh0Dcv872ivKVXMXrG3Ttd8so6Mc12PPyblDTSlSgv1VQ
R4o6I4Gs5qNJ2s5hxyKPri0IdYGOki+VmiI6ex5P1ppDgWNkPYG7xwPDrQbWoUra
S95ShcCS50Y2XVcox7GO391EY+69SUbNwAbashDR5RvNPNL7CUVB6UhFDxftnPUb
m0sL5cVOae5vv7jcuO75BtWBFVCJ3So8SWcw5WBVfyGMlJlMkymEjf4sd0tsZcwm
860mf5NRQZffe2SLA5jcw7/BjyQ/X0KVOkzP+bfR0pe2tBlb0zldMX15r0npxlaB
Qcz+lb9CZO3qp8sC3viskfxkLZDQ5w7lUKkbxyVa8x13zMQRXOkGUafRVJ9MaN5a
y0fcTXpq1Q4BStJFjy2ZyDQCd6y6Se4cUNcgFyVvMUog9VZMFn9ryZlarmXXVU3A
h5sPVK3JWZlU2yE5tZjw7EIbQkeXY9BauFBwrNZQ5MY7vFnlpy8zu1zv0EDaNnBj
CIuofoObsgnULTdJzcipqXH7fl+LOCThqg/B55YNqc+wqwgTIb5VX5UixtG8osF1
X+f8cBb+Wx7CBifuX7r3uXaifdmgELAYSXwPG3mp4lKn+uPvMz2UR43EcbRjGJDE
PAMDJtAywiEsatJ3y+v6krsd9zqkT+HTuHpMev3yDGVbLkQ1Rv85VStCce/0ySnS
kly5HTOEueuDbgp3PM1QkCTIEqtXKfiL7PGHtx5HKJbM9qTXweC1mF4sga0yANm6
2nVNjsvLU7Pxn8fU9o+8qPuih8Y/HIBKIU+9vNcaiks0Hi46kJVZg5GzleP24QuT
92/BI931HtSGx5oHX1guVSMT16kno0slC5uclv5X833XFKsnS9MaXx8VYpRZ+VnU
9GSIWhjixf4F46Ps0a6A/kzwTwHjairwo6iIEM1MY890wWduNukLTHcM07pLHEFy
nXzFb/CEk4/cZGOc14zYrDl9+8Wf5x9qHpvvOjb6V5eCaMatqWWyDqU+goAQqKUg
OaRMrOfgJdT07v8G7sfCwGkwjJQhpiw/BoYBqC+ggvfi65vvvVh0alPi0Y+6hgSw
0slljNFPT5dE5N0RUO4M4XSZL0NXWBzZAEUyRlROc2lt4ZDvEmY/V76qlDmUVRWc
FRFvy9cidBjUdrUM6Quhg50Us07GZ9xXUKZ4lh2s6XV5+IqLdgiwHws47vNF1wC3
G3kzcVfDZ0M7NYNltY3yg4wLVQJoJDvgkxIvlEeyEtD646ouZQq6mMqAN3Y/iz3W
8vzo7x6TNe4/MWBoNNoxVzVv6l9yjwFPAMwN1ego88Pu72B+BZ00ceCmpyXJQXfv
RglxbFhw9UkC7i8qErj6blJjlGjGe077FN2CzNBApXDC72cZFVpGDnVtXjRQMo9H
ITXH8USxH+uG992Q7KVs8dOEEeieFm4AC/KkTEefFdn7JrOe36USOsvnhVyZWfdV
mIWgzBs2bahFkLncw0jtIbWhsb5u9VOv10+qpTk0bnPW+cdWJLz4pT6xcYJ01Rpf
tew6GAwAbARmHqelTtmDfN7B18ed89dvXNXLUJtxyIrYph1JGOR6oVwcghsnStCA
FomyNQrxk0/xb6iR/GXSzCQ0gStjPvxE3io9RxEGXs9PvrgaEv5LHdMXO6Wolbnk
nMLrENR8QO7mV8Td0k2GrOYifC8IJ4vTj2loZVJ6BLmAJhkFA9faewrbhrRNIgLp
Lay9X3kFySLLBaE17rPCrj8X8MinGmgihmSNh9eeKPlH/dAybQWRz8oFC1utzE27
YpU+JZ5xgFDQpJYm2lk8/OUhUd7Sfare952y0VFEV5a9Q7ePJ9y8D8QuwTP/OWqJ
jbC9Ndlerg3MrCyje0fJEJ4rEnW0za9Qq+H6gt5GKcVCwIJuxaoXhMq3RoEF0HQD
A237hM5PEXPCkfFptQaByRibh/JST/UHqW6FnW241XTpaUoXDjOZ5i03uGQrZjSP
mDq0ghqajmRskcNu7/HCyb49sFCrcrxPaCzTjU8Jp4u+SBwShZRLMe87KbXirxbt
kfbulOmE/2zBluf1C1J1/p5hUuTrRZTZni2I15YWQUlO6nASjPpd72xInYNALOmW
LwUgeSZwqevzq6cCFbbxm4gu9X/iAUFol5t8rc6JfAog5Wg+BNXhcpvpebdockJx
FEaEqlugQ6u31ONvM6cN8uKin+4jKiTcMbXh0oEnN7aHPHHtn+YckB8JV/xOXEJ0
K4hNbtdNaACZuRlR5i9fr1HIA+3yU2pQWwxPnSG82NxsCczJ91jUoNq1rgBNhHdi
XcAxJvl1s6OK39QBormkKYdUDU/zwu8yxIYk81hV/sWDocpTHqJH8LzV2q94t+VD
is1aup5wBJPqnQcVmctMy+ZbFuDCclsCPhg4UMP9CY1MLPs1DZtLpd7Mjob8H6PZ
TZsyg3U4ql+e3K7eEW/31atnHzbWUSiro66Fh9iwA6Oq4t+jn3fpgLfqRS5KA4IU
QvYeFkrPZSXQKhLzqcQVqDZRxFv8Wk829POw5LdX/xofQq6DaRgFlHCpXS/zbcUl
KK74uK1u13qfsqNa3jkvDkBkT/Byo9VSqu6xtTJaTHBx4PGm7SJtT5BS7Da3iUwy
O55XOMvpiEwl01pwvmPy/jXS/29bDThLuzu/qWmrrWCf30tn8QuNE1BK7I+1585N
4T6Nod/DBklxU7wS0TWhOsY0V5bwYf2D/ZCLVzeZI7wMRZYLTskdMtAROZ/iZFrA
+0DP0OTB6+EvWYL0ysrzoNEFtBLWywG288QaUsYjleW1+EmTcHEacVb9kSJZ+OY5
urD1abn5UsuQR9Dy0Avjw6dn5DPpLO+a9OAyam9F5h367ItQaLrNANxeVZIpBMSb
BoZhO8moF3Y1FRgUX6Nx24RNrHwr36qS/fPccBawVjNg2OG2wZG7/MLT8aGrRYXE
j++ExuipU1ioJNUx5dAlRtp/akLmNbmBWgZikoa1RCK0TpdXZfMaCcKb2+o+P+ju
0pT39avab7xO5L2LSyBB9bYlnufaXRtx9my7v+S3/FOAmkcSUZlkXAuovP/2xjP8
VhSe1hCjmdy85AKV/HZWLRf947zYFqDptrv92C8bru3Dp7TlzDxRhHNo5/tZ+1UR
19R2LqUoPXomJplnTpdrBJ+4BoyJLzJ9cOvB9uZit90zbHh2/wO6Q70keTwotlPJ
VGgal49vxJGaBp4BfsEuyp26aMcWagtKPslQrSBgxYA4RTKdvZBgZagclXdscVSp
j89kaeSm+HZZU5h3l7vO7Elj195TvnLKk7NkKxJta3UjWDc9IZKX1GlK7XTOxUvx
gkWzXtO162yrXbl8GRqSyQkgYWNgJ/Vj+6ZTi4g+F7CJY24jn65EyNAOnTjm47pJ
2Eb/ebsC2Uph97V/XPX3jRty5KsbNhMILD98KAaFaWsquqKbVR9161clJY+pK0Tv
7wsNxooWTjvp/33xQ3WTKHyCLC1Z0S0VjXEkX441rNIKA4FRAnfzzUBNNBNAnZdm
waiF+at0CH44Bv38fCYLvUQTdIFXC7w2OAHdgvQYEAxKz0ZheYXY2Hoo4f64r16h
8+roIZwn58ZcHViy7caHNxR/mlXnS+suCUsx+OKA3AjpcGg/5GHzRczz0h5SCJOw
0i4S0THomh/S74X1ZwT8Qbw/S7PO5yGtIQnOi1YlkZan4EP8mEFT6ZBXDAxa61QS
dwbC0/R+Oz/ok45y7wzigyom/vZlHnV8zOc4nZW9wcFOS1qF9+5wHC+N3ByZu33o
7+kXJprQXevoyBqChm1pjrHI4xOaO4cKBjP+JrepDoHA3x9GYhgf6HbOyE1g3OwM
/OjpkF5GMjy63N9vo//jWjjIkd4TP+/Aovj+qpnc37/yMfqTAmgzj/8lQjK/UrqP
d5clMTutOXKLilM9tj0LYZCsyld3WzRnHcUmVXtnzxsfaTurO9jqWGmLD1Yk/np0
91E6dGvUhxQSbIxODbY9L4BZ9TlHaDvMEVAjh4x7XgMXmjsRZXjdEOugMCc/I4VV
/+0vT/BkzMTcx4Wraa7Kk4WQ0llVr48Nv9plNWABzTCarIGrfsrPWQNAdjHITTit
xx9ErvJrOd+APDeRQaB8twLZTqwlRbvDoaSnWu/+C0xDZWU4Tk1O9eBzbzMxPXpW
ZitHnJlRcx375xBKmt8o3V7Jj91yIviSvVNYRntfjA4BxjkO1woj8LGFZXZHB7fn
068cukFum2hm+KPwXVHFZj5l4vx8cMIMpfzuEkaUV2bKp5egDEFxnkGxFH53k2Om
/ovytF3Wz7/t+WXuVDD+CWRXUieAL8ZtYHkDwBDNwIsyDNTDvOBUqV8XwH11uifc
gso1ARbehuAZqkSkKUwt+BJcN1WBXWpBEMVE6mWHla0EL1IXih7b9SgMVSJZ4eCV
FyDt6I92roNT4DMLhsGa5k7KtSYlfBoRaabGUjCnJ+h9nvqtuXG1Ru1V17G/GuGR
fZsKgoZDVj9SOt2PK+IJSdlYYnofnxJo5wXwcCatM1ogj8XQg8fekm2rToTGVxKT
I6YJcVS5rGcNEvmQiuLo5DdB2FNyvSrxQbwa/m8klgBUOYvB2cylGqm5qxn+pdfy
LjXsWhElEo1+LvBhda8ucLNiQBgUHNM1F2JHUee5KBJcNr2nc4IjWTiGQQJE0bbl
sjpx6QIwwkbxJFCkhPchoZXI5IF34IglMMuFldnh7me3lGysBTR+pVEj1OyxNVbo
A+DR8KxNk/01cAnrg4A/kn27ozwQ/sE3iM5UtzD6txYxbcJk2VKxvzv8nwUBpu4W
9uYSTzj2WR1Sa8YXNc8LuUbsu8VoQbJ0Si/mmNy/00sHA5rHbg/KCDqkpKOqnk3/
L5ECffoDmJEiMKv3/2XsWA+tmNndBXCXF6jSapsoVlFV9jTDWeN51ag1nxisbvR9
dGfC4+g8+ID/yIe67bQL9g2egtn7VYiIXAIIrOxFf7bQUEFbCvKyYDjgogcfUvx1
ITVMFjESJgByaHWAoUtpVElOwEEqexWRya8awZQ1or2enf/qAM5xSK4phanhc3Ae
KgZVDcDDnj11ZM/hA0uVJ6WjKTX+haUwYroljMoczcjcwd32K8Fg9RBy1mphncrp
OHjSFqzsHl/7ch/ww9frQW5dQaQeo2Cyzk5j1LS234EPfS8bGIbvOyxp17QObH1Z
KC33u0HN2avuoS5f3+u4nb/6gGg/T9GNuTo0ZvTYTktLmXYi9k+NY2ny6LbMbnqC
GiK37hcQ7jyTHtEUMA+t6lT2iuVmj0Vnv5drH4NM0gnehUPePWpFEu4TlqUgbXey
fdAgNEAJsrQmoeQw4VZ167+nnH6ncHzuPRZs9DGiCM18VW9jc5V/jWwggVlMy+oo
Z6gyG0QLmvTClFwf2fuIrJ235RIGa1PyVrdb+A+7NMDRy1fMRYa9W0e0W/Fuf5Ri
+mF3ZhefL0HSwtwcIZZO6IBLHW/piNno6xc8H/AVi8bwUU6GgwKiIMkII0NGGxwe
WeWBwurO5phVFjwjJqI/bLf9ScWa1HIhsA9wWJVPeojD6k/HMGFW1N2wSb9CSqTY
X2XU99ARRwxR8kweYPIDAYalLa+P0rO0vtVKk781+hnweaKKwpM7zv+5pCFjmi9g
jQnCeupasvq/EvRoWy+wzsZ4DDXVuX6zgbQc4HLswr1o2t0cHv/tbGJYQi+PpGLv
nb+GFc9YVjlFKHJgtQOHicK6p2dH7PqC2kztrNvClYqFPSWGkslSrpWGAkHP6srL
obv9RXcxBoYrR5NY1VY/GbtYVqTSaBQtZT+zlewjuvaUqnq08firBed8luZzJ24w
c1zNkPzo9P4WcQ9NZgb6dJAcLd8A7mnXOS+VsSvT9hNLynhaIJPH/sK/J4YZKbG/
WSVaf2yun78afoiIte3CkwlaQlVB/2xYQ8TsTS++6+Po5+9SbKqN4WWiqL6YjeJ3
mPnhBer1DRbdcj3yu1pT6AHQlmYE9H0jQ1wzsuWxm0yKVDe7ZUI6+Ioo3pqAWLO0
JYUGQZVrBVTfnBZ7aSO8AEoHWwxv/kMX1QSDMvKVagM3GWR2P/EZ9KnoyGZarqKZ
Sv8z5B/9pNH+FZdahC/nE1R/xjxtDIO3Nzb7iWCO5/tiHAKpOsk0tFehKQjKFYx5
+18pVXl1iHQIeBZjCXGKlO/b0uo3oItFcgUMy70CNcNbc4vE2P7sIvQKjFiGyhwL
cOOHQGxVGA3V83JXA342/avPLKqFx+O8iV7OvblLsXWwHk2UTC7Xc3fHAZ6p+77E
ETScmpY2H2Vyny9d3vjUrIaOQJmOVsLMO/Q+uBVvHk9mRQGNWkAO9SpwoJCRXtNr
rwrlQ6ceiE5fwcmRIhflOCsbkvG0PCcWhZNDAV1UgSg9FLvxQd1745Ef05qoapW1
6ySXMhxyxe3KSkzt6EcxtlrevU+Z2V3utHf8EsM30C2Rl8OJItrOYhHtf3apI5Mo
8vAjvAwOFJDJyCg16cRvhJpRNGAFnr8Jd51kBy5pBPC1DF0Gi3BPUdXhiFJdwtE4
LwarzzE5PC4RP1xEwMFI1b/FeXsx62Q13Z1pA/Z1sOZlsmqFliMjJH+c/XsU8bPo
Eu8IIVKXUeqJQOYU1AWYWsSxurmeYIX8EhDYQi1GIk3JTKRcRGdvnnOjng2AGnhn
927uocZhyf7VImfxYzb86K5DTAib5Don4No0KYFc7FTLLLFU0YgJOZD9523zFLXM
o7WVDNQ+EiqgpdBxM3dX9EruNr4Y0fxbEbGTnTXuB5GfSK5t11ztmOYzuoX2IXi5
/8o392vp7ng0bol0T/H1VcXzQwCugi4X5Y4JvqlZ3g7aZLnda8sf0cwd60t5sE/l
HHscKIvDTgj89ZBN67U2GDMwgU6+KoI7iGk2ymL5Zo5PAWQAiOzirZu9TJ5YVpBU
vsNdqf1yYJG6bb61wRWeCe+GAB2Rdf5OaFLdN1CankdX/6g0He8SNX0aI89/CHSN
IsS8J62+Q8y4kq2QTbzh6FqwnqQFz93QRu1DxLcL6YvrrDVeUDtFH5mv4giflMYp
v+hNuiHh3fGK1Rr6eQjYTcqWh5kqpOBR9cmoGPaZdcbqe9DH0Wvl7IJPuW7S77cO
5A166FTIJL6z/+XlOU/q03UHjze2jXWanrKcXclF3Cwa0wExNhNBUU/HsJhSWR0K
z2L0kKbJADc5F1KuUi6nerbYG/31uQa2w8rMyu7ME6Ol2qHo7KisVEN7LY1rjKwp
k4XsEiei8YmxZil5qzf3qRzWbAjIx+OnWLX0u8KWE7uE73ZoomATFWbMZ6vKSRsQ
B979t0HvO2R1CLWQ87sWHK+a9zE+ednZgzkTZNKlNK8jlw7dNHQDN1BfCUyrqK35
obYNmTQ9IJ50y1fUPKNKkfIFvQ18CoQivCGAzZKvRjBYxxwBMFDyw5B1g3dXhiXp
7mqAaEfHTl90qQ/XpqM7nlPXhQ+MdoJyaWiMQq8HJoar2idWmkJiNPNIQ7T9/62o
twBUxYmnw85hPvd6CDjKTlifdgwXd9L6GEKl3uZuZtOxmflAhK432T9RqEHbKPUp
FeysR1cs2FgE7rwKOKqUvGXyTf0Ogv16gJVBz8m+33LC2T/SJvYsTc2klP0wl/O2
hwz8WZ3y7qHkxYRKk8lB1pF+LRpfrxc6jkPEjAJAuIASnRzmgmTyaJ6FWwBmSG9j
IPLzqwR4Y643ZwQR7OZ1BJ6mE0JYHnbNUjpY9c2qMNtFUCYtFNowIeTAVUBZuLN7
zDOwn4QPjCHVu9QAdQApBqoMo/lW7JXCZDUMMZJlLK2mJi9s5I4zsEjmxjGU+oPk
uKrfMZlDA6fBr/jyfk3Sk8MEgaCagP/Fgc03nZODYKd3AqSGLeiRULiZ9Nk2iE7L
p7cVAOGXs1nrUwWGJVMdZUiElFIQtaCasAlp/ESq7Pw27PbPNigZpx1qKdk4oimv
G0AMhBqHkxzOC0NtQMV2bG4fa1MLIVeQKCBhGp72n8wGvG/cGe2YSkq/HrWgYFXt
/ebPGiGUTjLKoI9eXh02K+KsJ7hz2KFgniEy3uFeUaV+nGcqjtJnqYzfIUgB5WT5
J4n8rKxh9XxTQGn3H/2YiY5lajYQNje3Vy6VR6WtAltc7gIUcr7znGLx7PiCHjEQ
QL+vL9ggmhhjlPA2aCqeScTO7KJj0KpcxwcXkdvoHMIw+7ZwNy7J7sSmoKBgzmaq
iCxmO6TFgb8ykue2y5qAPv08/RsfiokCYNnJaoC1jpa9rPbpMWbXf8q4vxEXHa/H
bVMSC3EPTM/Txi0BuTBleQu7dLAWLcRMZVbCuN0zufpk2wFCbJI7thZo+jrHOg72
onA3hPBgA+qI9vE/Yyl/4K46JS04bWhe+Who3BzGb4CJJzN9ZhRfsmvu+CL5Q681
r5DhL1wfHXvLsdZFUJ69raghm3nXrM7piVc9G68k5p+r4Dy2QO5CKJrsQ5w+Nmil
jMd+6yX6kMV1tJpBvfKutUs21TMRRdV4QKrWtclWLkXvH/RRF4SMPMqd04AUOeRs
Hrk1zcEKtWW3X09+1505Xbxr/emFX7OqWaQYQeDEyP+vkiCC58Rmo4bqMv07Xpov
Gtnq8ogC3Hsh3HmLUinJz6lPODAphEVqtuF0agXT2zFtcUdj63yZAqodl5ZGhDMT
ITFFJCtE4GGwJT0DiGha22SdKRpd2KSSTbRvVLO13ME2CIzpZwaoBj4hhy3WMMDN
BDfLBeMbWrrL9Yx5xtlBdYncZUP0g7JYCZelODCMSzoGZY4wtHx+JdLtb1jiVoz3
ZLxY4yQWYgsfa9zpJiT0CrV+E7Dcj3Sxs13YzW0RhVqk8r5zZrf80g+ENW7DfMAA
UyLzz+eISWYNMA7wswSKjif5tsycKq657Ud0wp6dQA6IKvG0RNu/2AGh69s8JlBB
ufENuN9Y7cruBx2Xkb3zPGxD7PVWo8syb6gASoqy2qoNbvmq+QgaCGzpDEtg6e+t
aidInt1KubIgIatCB5OP0YLD4bfNXi06xzpI8pz58te8yywosyT6Heh5g5On7PDh
NZ0Svyi5oiU8EYImfb4pXplp6uDrsOX/9Cu4XcN9nSA8AKrhPsnG19NIgB2rYXZT
PXkB9O0dVy6qBY4qDTrZrDR+wXqkSST/jzbBK8o89COsotDJcrrvaWFdg8DNeN5E
vbFJkz/O7mlprVMwMBfTCbpO/0PxNEx4egWVwTEqLPFTD/C/JmqPmV57rIejtIxl
2+fl7TK45PmN89namq1qC3FOeTfmWScAUnOCc2IB4su0E1++EQ1EPtdsHF7tiiv9
/56834WaqTA8qqZWlOosgdY8fYVDib2E3Bq/dL8aZQ35vZQ+osBpzwXgog1qQXA5
lyu1e11tApj7sobDgm803uIdBZtMh282Sz57QkcdMzUzTA3EAfP1F1GnbRRpWBZM
33BKVuI83Sc7Wsl/BHeKa49nkyq9fgalNcSAUPrXNdKfkD+3UnP7/LOPfxHVy6Cn
GpnW4W/99orcxqXbj37PQwddcnToOz8H7rHryiGxbwuNOlJtZRRAQ/ITEl8r6o1T
Lmha3oXBlRkv99UePGEdRVXsnsIC1H76Qtiq54Ur7eq2FgENnwyjJRfcyzzpntp+
NUkehW7o9TVe4ukgITbN3uPyW2X0tQrA4FIt8WuBsOfF7oVrk4pZkmgTN6QUTKcL
Zh4eHYezeHDCpcYBOnpkLlLxnA1SFvOI87896OEXXidEP9N4smAvxcGUenv7IA5e
9mcwri3+7ARkAUN1EltcYGFKDm1Z1qCmpkeW+7167k/Fg9cJ/H0Mt0dAakFZZ7/w
HGlcW47/MGQc7rFaxqFJbMOiHxH7QPDlujI8BwaA7wzYGMV2rnbWPHJM504Q0lju
6aniq8DpEiBN4BmbJU6+6stldAxLnV1iSUFWTy0ytQ38Bb2cLWh8wJFed+ftTmjx
nBdVBIG8NfQ3597GFMFUwNksbJB/iMUH6QjjskO6DhLgJS2tZbpZvY8Mz8W5AX0y
yw8QEZ+7QX4XP/NQRH0E+LHEfBTE2cvXvzIce9pL8istkPSji5zBdeR6EI6n/4Fm
ect8S7I/j9OD/sxZfQNlMacjpdZVv1pC3f8odL81GnlJ66KtRv3G6JVL4O2OUKAl
eRziUszhUcnGL8hhcBpcGgh6e/WcNKQUZMdQSByRY7FRzze501tND0lWfR+Q3spY
kk3xvwvn48GDyj9ewQ02APAqR21eYEVSwRD+pViB3HUVobsoKhJSJl+TnTah6NK4
CXvLfnvD+4dcQ1by+E3PR8VJ/h6a1Sk9qS/1+rEIUu7zaPNKLN5W1rFu6bDjB27n
5qDb/yxdnLD5rjQ7Bq+GZNGCxvfhl9vR9Q8tVqPsF7BdAjIcI+PX+1z8h8dGeuyX
zVi2fp+wP2kK2E2cpvIPU87LP3ESboC+A9C9kPxshzI1fqBGyhW4ZNe1aJkDUtOp
hlqXMA3ECP7/qYhV80aRrTPwLqd2C55O6i5aA1qcMkZRahPE3WBFR5Kf69cd8H+P
ixz+R6aiRzHgx6lgbMF7Xqe7Qlhah8CJcpE+jCkpn2Kh90xtXn5pfSL4eN24C68T
1f5dnT+fJ3U4NZJnoS+w4oog4Xr26k7zCIkNE1ak0OBBr3WckC64xE2aN/kfPR/D
e3XCl3jz/0VxYn4BMvXY7hS1hsJcSFVYBVIY+udlk8k3eBnOd5dszyNHq3qdr/jk
jWE9MVrccdwvn1Cj0Oae8B/68XierEhEWIbo6B618SffqJZASfOGprN9pDOxwPzk
MTwT+9bjwtzVyUcqWjmILfBGKp9Jg4ugG4dFQtBvch4RhE4/SOerMJRSOJE9yFlb
2+gthuZW6/M8zO3IRUqP3oeDQKcTn904aHFGBKj5AvNjFBmc83d1fmE0qVGL6jRF
iH7EBtjD1CdgzHdkiVFfnF5zh/nhf4GUN+NPnGh0sDJJhsIWINSRGG0/ZumiCUYr
wbYqmw6INpUjAM32de4Tg9UerrP3ywnb5ERpaxK6eCYyUD3DDVYJXWp1Kk4plh4R
dbVfm83CKtl1dyH+9xxVpRuybYLRGZB7mxhOikvgJPsxyi/W2ma0XhXqCxD6Lq4O
Bh32bgr8bpfWoxSPJSjzFhyqxzCU9hghQmibJDKyLzyaeEyrq5c+dCmfwP7scOr7
F2W+ly5hZns2rhmNKiZxcoI+TVldeZNyp5gXcVqfhN8T8H6wBqAQNhvaPMAZvtC/
RWzatRjhpM71jukNVarXdaBN8Oqc2ThGkmUzp5VgH1TzLfOXMWjmRVUAUX2DoUdE
Z1WUSVBByd3A8uRJTraUjMluRrAi8qhozON4TRnTVD75uLjQYLci2C6uAvlcMUZE
q8whvnOgL4G/7FQE6xfVpYDbz9hwXHrC4RPFeXG1M4k/UOlUMoKr6y+sa5tRUovi
4Q9P8HcnsXuHRzB/y5IJn2bRLooOOMC+M+V4+JGZ0jpcdsoGxxahPEZfjekM51HH
IMOsQQAjVKj0f45f2aEX12dywNgOszGcPg+9pxsSkYP7G4wNO7eLa8ryrML4c4/T
6v9+CsqlKY55r9oqAJRs/poWigrBTJINkg6SKbD3AuBYtvfx3FJAMgQWZIo6BLbI
q+PjjmMFQqPoRKbQbEnmIacs18zIWyLJshbCaZNXUhE9zp4BqbrLz30/+zJBLeXl
Z6t220/lNxsvhv8F3b/oi64Jj+7O7MtSF+l6zJDTy2WmM37QXbVQDGJeBHwTHmSX
xR4HrgZDJlH62unPjI3Z4rQT/4NhVfzsRqYcYhG4zp5HSy7d+lfqBs6P/VoBBZbR
F8FilnhDFo9HaNLOLQ8sECLxa9oShuotl8haanMcDNFeDsGXD1ZabYDy6fVV1e13
qATNj7zDx4mMBcbGiZcnHbu5GH1BI2AJ27EnLHskT0A9GbsYRJw089JkzpDGRqJS
B9av1o7nQmbb6AgJE679m70y/wLqI1nXAMPwFq0UbOkb2cPy0T4x8LLs/OPMpJH6
SpNEWYifa39VgcR10gB6EHndTPaCEt2YdiQZG93tZ1tVkRh85ElWFdBJIJbUrb4k
`protect END_PROTECTED
