`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OF46LB4heOwk5JGFKxfmg1oYHHikS29F6bsJEox5+zTnP7InZmtKm+97Scnh6rMX
zmnvDVS9gpSceC2gh9cSni+I6FhBlfKO2LcD0Z9qTv3QN24PH17vg38rWzI5qyJn
aFoNY/RuOo5N9deQ0W+IDFsP/+exEAYGGwQi/+aCenaYEcev67nsickrRYryETAa
JKBJSswhysfu/wXCVbghqCmx80rCWOU8i3+1kp6/3lQBcndievze0PxGOYYJITaZ
YpA57omxAKjV+vIW+oals+BIyA91vlLUgogBBnrzP1yQRR1tI43oLRliazD683y6
ZZOUCYjbOfnwfasXM5EGrclvIGp8tNGWiZFy66WIH5dmmcDiVknq3ExUyNSIDgWe
ODRJDJg86Pz9qTVJVpSbdDVCxPlo70UtGcjGa/753E1Z9qds3OBrd8eWS9gcQuAF
FRgpS18IjQDMbE9Bw4rPFBlGQr7A5QUUmWdTq48Jy+3sJ+qy77xBEFjd7DuYER88
P5G+luBCvz8NM33yLK/mAqNDmZMtBflw4JS9dIyQlM+USKdXeR24OfVz/NV6GxdZ
Asx/C43RxFYZwSBiOB8PCOZ9rFnq80/Xr4+bCvEnCqNogMv5RcvVo2If6y1SZTmR
y7h3beG55gw2+H42fkMVlMiG20FB12H8Qgr8Oqunzonq6z3CpZ3WF2P8yntIpotU
C7sUQGnLAS5oeDQwTOcNoXxR7YOpiC4HnJvmWZaDpeUkY26mqQ2ldK/t8JTca7J/
e6lQtNABO2YS4vaJlTv5IPdxJEZq0NFdlQzK/eU1iAK5Nz16h+Vkkl7WzH11Xn0o
cn0e1gIkUpOePdedQL0nnc7HgifOygQn9IErGGOFJY70mXhsD2U7bTRkytO6CwbP
xeS2isINWpBsyPJaUp7vFDDZ5nMgZjjsx1mQhCPN9qqir51TeqM9pCJ2vxCnZgYc
4QYzF7b1DG8kM7bBf/pyt6Nl1iFf/wyxKbP/rr4nWkQvRQmumMp2iFRyzfA7OttN
+EHJvtNYel3tyw4909Gm960Hd2XJgVU4rM4o3JtaTIhvxudEnZWTb9LBekRp6Seg
sIXqfNF7tPLkZ4chEJBrpjvtb4lT4rtrJ/NR6ERXcboEQg96dbi3SGwSpO8hEnG7
thbRgggmRY6u23QrRrWkwD/WhHvVVq7QcMkv82/4VEKrC6s3oV28SSNdQLqboDHJ
BlNnIr+ZNtnWcI9X6rx/e58/dAmgsvVWmLNQCoRM4oL+Q29bTLPNhzdHYPxJPkDA
iwdP3Sn/sSXK01aTw1X1n5S++OePkYsJ40ET1GtQlQzJwPubpC2sYG727l08rDLX
1wEDSkNpCa+XUKXvXPxFwAzdR2WjFMahJ3aBHvNhEeBRIagk+ISSFm+AfObkEOiW
qBYTyG44+Q+C3HNu/I90tAyTOeobcNFj7OWfQW2PW/yBt1y4UfQBe4AEDQBa7u2D
sccXsbIV9/mz7bupE81pNi0M0JFwBi0/qQeLtFrXiSfJpCeG3B8LPs3FHeVW3V1i
DWBksotuIhGnsTdDSoohtrQQeZx7VFnGX7WiTJt2lQoZ1dITQ7He4toIxqXx3Jfy
`protect END_PROTECTED
