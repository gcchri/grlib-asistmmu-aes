`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mT7fYdYkKh0Ud7+HxZL7ovc12KOBE24+AHfgKbPFUhYF7bH7/8pMIuUiIopEs2F9
ZGLwfjjVFPf0C6Ta+vNOtKugPNKlxWEgcgpKMv5QxRbsiB46P2vIGZwFiMF3cr7s
tl33d7Zw8sZVKTH2Z0YpIJITw479+OeBdhccR9k+FyjPUkhmI/KPvvgzh9uDun99
KSaUKLoxed0Iq90SGlINEPjBY4h5XGbho6ZIGp4KhYnwBGHki9JtxlLYWPM1RIHF
cPFvxsWH36pGhXebmzr31JSXdHsB7+wi17EVBTNiG/Y8BdcM6HqL+zsMP47naUfz
Fkjj07fBrpiJiGHcTh6HpUIaCgaGR/axCini2LvCv4ETBdoXyCmwZUSKO+T1Lafe
bhM+41PrPycnf8fc80bqT4dXzcEDfKDRyupghqeDNOkPDcHpc9oGiH9IXDLLMIHZ
fHlqbwBLAlX50UhAScrFwR4P/zqjogu7LovDnD1JMN86y9A3tFlOZII3kzDYkPcE
o+sjsol09U50nM/TjG+GPu47tIjMf4ULQwV9VJknk97agYDOjaYBu2NVY+5MpCY9
h7V51mTBDD2iYouO08INeA==
`protect END_PROTECTED
