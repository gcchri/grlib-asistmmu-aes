`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QISDavXpM3UcFMI6xUODEmKs3nIAM5A6mdWX9sqlaaSlDbETTYlj96UFtUhj8y4F
VQGw0vt7nMCEjz4c8LOFg2nRFfucBm2OrGbUbU0BXsU4HCxVImta4+dkE/NOsbxS
xCdWS3wXa9jgRS19vT+WTu7/mankaZV8LgV8aujIHHKYz79hBcFfzvRGq1UfPaFJ
E//70IadhBgYG1ykwC6Aj3ufrgPFMi77iEx5E0SMdJiaPzxBuzs9F9L8HbEcXZky
LZCZU6sBsxWuKJ965L+/TkE+QXmsmYk61Q9E/gFHoPe/kwcFNlp1RmDN3KD/4B7J
Cstn+iG3IIdM7g+35xEH73vk3cw2YWTqMMWsq3yZ4/pjQOkgaDiZW7JC28J2YDLI
nxeRP5mAtj4MUk+6I9HQsA==
`protect END_PROTECTED
