`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MWaeHb2fv6MKW0QuOekPGwlWcycu3Jx72rfP9jak7jwM1A2f328c0Y/ujMVCHvKf
slyl2RGD8YXLt/xODWq3OPZ8UvFD3UJVDGveg1RJSlyzrnwcRqWjl9J8xettPzK/
R37VETInPWXkiRXkzAKsCK5hW6wSSy9OWUQhDaJFt8CLys2LDdaz7foDNk9NPqA1
DpwRSh9q2tXXaN9qktpv5TWPKj/cvhKRYWYfC+RxiG+/dCv4eiM8W/zhE7zSydxA
CifInEgthvBSZqUDPtiZH+WwCGlABK/VoQKxivnWYyHpVsdSwqy1cXiUrj/W9PU3
v/9qTRzzcWZJ1v8tryzCfurVbdLofOyYtp41Be/mKjVJq1x6dFXy17NiNlb5YIzl
vLNd/tIXHOQ2l8XneNsYpG31eAztZ/qXBuH/1lj2z9hCPZQI41/TbK4e7cVb3sbk
dg/SXg/HxpAsE4+e8J1X+tPth6CkVjMCuiZb/URpBUbV2wZa1v8d9++sLvFI6eF2
20BPpIkR+cbD4Ai9XceWc+oDdnHcxDqeivWhNo5hz55zvjJ+WVk1Rg1B1zLZSBPZ
9jA9VaLwT5JdTiyGdmYAq53ruPqVdKlzaXkyFDIZCMawnTTC/U/rahzpqhCI2k9+
syY8BIyvGxlbcA5u2FgAaKKaW9f5/ZahFfBtrl1TU6Bvvm3Rc4BjekeLysC5gYbP
hwNY5d9ZCx2WlzZx29S6Vi2hgLvnAQQ6VoLFUnKBcxy7P+8qvQTiTa0q70yUb57W
PObcys1urc9mlRorAYNspofUfmFSz2hcKqo9uy9akjjHJAqgsURbYajo8UKJytzA
FHEI6eYsthf0YyHab/s2/2Okc0C7Re1TffKiHYmXEdmRnfENpnMZ5t3qA78vugJp
zuN8mqaHEC3+zbVyA8BQ8gcEizsdRW78pqFYVdeWl1F4cDDm461G9ulYIRyRsxdO
94GyO8fSiVS6bOjC8rqiMmRJY6dCS2vm6zS5OZ5TXzMtVZpgcDFAi8oxwXD4kXgb
+q+4Qv0FhpiGjNkuKBRly6a0l7UGoW5LRJIi1EbPn339Hw7j11REQl3oydUMc6iX
uP+NZL7eO7ElY7s4KQzE6/0uZIxXDwVFmpMQ6Y19AZH6C4U91nnLcgQJdZeQtEUm
igy6K6dFdVTG7DyIZAlWAoReG9UexbGxm/QhvM+X5L07CzWmNhi7j6u5SPWTXQ63
uASgJkplcvO6cvrpATD3zSvPiv9MjADKiiohf1Rr9oFETe2aa9nwBhDzzrgFl5+N
7diosdpD4GOaBfYF1K0ncaw9a+7J6vJV9acyc2Rhwz5TdJWTVaWEGkrmGR7QN2eq
aMvK5ZhW/iGR2JeAikIcf4oB6jvLLJbPIj0COCQnYgj9Ki1FcRC5ds3dvso7/IZB
DXsG8m0sXcgG+c0la38XezkBJN5xDO7ubuOcX6KSF1AbThxDbR1hlN/w+uGR40UP
+++z1EVLiltTZWDMs4v8atzw1ZyPEP8PlhpbV/Hh8Dt2IWdqlxTb2hcCPox2WRlB
qtgbXjQ4gJxIxfw/jaaarFsv/o0j3yE2cbWHKmvM80/HOGefOawO+FvtiSp8S/p0
J0klOYRqkmf4DNa7mWbmOQQgeJjrofgudwhOvO4E7LtbkLB40ws8CCERA3hoWjd4
u92afJ6tLxRaHSsK/VXG9pYAW+pa5bXx4f0zdw8GJwkyC6aS9CzUruzTVudwOC1R
xtyQz7anCriYoSi9+3AG2kJ/ASAJGXIgeg9coT7Ef4/tGV6tli16CuqMC5PHlf5c
ry+po35QESoVyKo0uch0vvt5cjaYFv7nTEhH6HMpiguF/S8s/vqaYQWEGFCzttWG
2JH6iJ6lwLqRUleZEc+a14Hfnb3iXX0zYzeGFEs3i64khZeO0fvEM338l/kLttIr
IgU5GxapXIYe4jnxb+YFfhydpdPzmVMrzs4mx8kp2Z31oc4BqJ43BxGRX0HBzevm
BpND6LQoYM4HoYZY+iMDwqDcZVgnMzaTyCv+bULruF4hV9xWlg2bpLgT8vKdeJD8
7ZyK9+VPeNqei3RjeBkIzGj+4+WzpiJcp2424zrwj4M0ZeECdAjfFKowdgQA2wWA
diOnsJMfJHnZ6FrQ2oAqJYGg+KZwtWPlbnHxZxNL+6WlFLQ110EFvjg1g6bg4yon
wlyuH3HYVPMz1wWFYZ0QNsOTcNwxNiA8jwaLmc3PyqpAaQqcSlLcc10O7zFoA8q+
eKXk92enaszrXRT44V8cI11pXgHTCxbOQrCcvNuRBUYWtP8vwMHJCzS7/xG2NUNt
yyRHChDjfSGgD3xl4QxBlbXHdluJvNvF3Yz637NNFxtOhOsvnf9dZ57SxxRMrOih
UH7/Fv0qxkvVwXWvY5BJLPjmvI3dhpZj/G+/AW38O/9VAB2Jm1CS5+kIQHtCT60h
arpIIGF/XAbUo1pq0PNEDNbwAlFDqD391pbDplxSNT9ELkZiu7tjYepmwmeEF6SD
xIwRTp6GbE8qjumdzSFJiQEFlKd/BPxgQxeYedihxIx4ezzJUlVMff90ZrXwNkTF
7SLvl5+mMNphCu5exOPkUMAmWUFbHM0vImiynYZvzgZ4Pz2QqwQTfxr5Amr11gHr
U053k33lcqQwqFon9NQIYSUyIpEeX4/7AbsjrobQGbV5QLThoaEuEqkQGyB5Pc2i
g6Cc0b37JGwu5r5N+RzylEhiw96xd7c2C94Suv9DSXk=
`protect END_PROTECTED
