`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z8d+cHQZYQXCsJ5hoOGGQPi4DhlpP8XIX7p1hkHY8yGe4VZcLI3g+Um9BwxzRHD7
lghm95oFaBS/5Edf4yYV2cPYfELpYyJq/0+6xAglbIuD28puWzdFYAny1JiTK3YC
CXyPbziAX6r72qe+1LgGqmMTL+oMVEOWOPTCGAQ2WKjz5MklZcWaBaCx4k8b5sUA
ZF/FFnVxP+KB+nPQD9EAm6AdbktnT6FEbzNrO2AFDi134Zphd2KZ1I/EIWhVqvsb
lTIDOXH/EXRz/5hxrbdOODRzsnkcbRnuK2ra5MV3/t2WPx40kOezrT9PRC/bFHjy
W4Eh7Gf8P2bzUoxJxhpe5vIzdLgt/kQOEWHJ4hA2Sux3oKg0gTw6VWNUtIb2UMrB
`protect END_PROTECTED
