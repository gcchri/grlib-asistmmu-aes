`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/9YZS9YmiX0LYx3uJUdQjTTaulNRQQ+c7f8P97f8KSEZA1qh/TabGpNmrYf5zWiQ
XnX0xb0SI8vq7N8YYJLjponZUBubwn2TO91oDGSRDksIOB3jZ8WloCixlg6qxI9z
M2ER3cTt2j7/Ycl6AFO9NjVvpoMsM8KtGURPF54esjoqqVAxiNJzsLRWys1wcGBv
FpumctgNbsddNR+qSpGBSANw12EpMoH7VEekRAgHfUK2+TRDifRgbS8jOTBnCEpL
vxxoTQ6DDbjwBowmO0UNQlfzKJOap8YE+yjpHPuiwYgNl9bl6b4zpJGyDL5S18pn
LaEK8ubxF9PVU+BmAco854hsGVjzVWGh2/70O5vSzbuGlFEKa7bh2oZ5S+Tsw32w
Z9t5rForxvYwYlPg1GWHWUDiLELmZ+6/UwSw358gcs41HdTub6rcumyLgftzVUov
Gt4zhwkBwEw1Q1PCAPWfC1woNmX65QXqMU2yGULvzUUYURQuhO5P+PbovdqFuqjV
haFqiqB6KTvCbZVXfnCW5ADJB0GrmflYQE63HC0R+I4fuD/k5//ejseNom+g2TwY
POybg7RaKm9eBIeqGEV5IC5FLiDFtKRkmChDNIneWUSs+70LSr9/Pgl/aEdkwdvk
uIz5u6pAJl0+A1j7jHtgGEeAATOeEpXEgBbm5J3tXS2nyzyFcB/NFruXHMMrkj69
prkiCgaPfYOvGvMQXeoXD9zKP7cN80Cf95r0leFWF5PtSVOO9Xv8PXpWC7d92+vK
ZR/FsJAKEQ5ulcNcdeQShkDSFYW24VMV6HygGwbRZDtj9Bh8aXNNu6EwCWH8WiFL
dYyS7ik2TEOCdKeDvf7D7JtBa5mmOZCTGAjnDmk0mC4St3Uycd46QYy8QyUEX9cb
nlx8ztzEBJRe/+aIhqg3qAL9hzMQLPoY7FiaMaqlkSW9oDvzhXO4+fUiAgiXoIgh
Dz1dDc5oe0qy4czqMtmjLU/uEq8f3bJWvI2LVKSmSTTfmcb0T+XTfzp7VPEelv2u
t6s3wVZlUHxvPsfT9DubwMzzdECsZi6a2WwpMZQgfMZS0ChVi5Jwrw9nQLW+hFM8
U0d+qG/c38gLM7mTvI5J1wqmE69MHFdVagozszzSNgBNFjisxwsUxZ8EsFxseDWK
vU8IAGj9MJDRcaF7muWqI+EkH5k1Hsn8o1akV5YSdg+08AUKYCsYbD45kjg6DEWh
9zHuqTR9AWKeWBLmrUnhsA5oT2lkHpo/dKnf/sgL0UfTAvr3ZyKyjUZMtrsX4gm4
4y82hpdglilapGMKtGH4QUX447dTVZjzTL9TXeZHs9h2bIs/DwLe3hyX6HYdJNUZ
Ks7cp9wVZ6MEDSE/0TiLkQ6mivaTQ5SJ4F8BY0xeEDEl1UOSZlssuOz1yEqH/YX5
6xI4e35L3Q8q7ut+zX26x1ZvqbfkSH4EF7qA1oKg8gkAsiBYVFtC6urNW5gX1WQN
0TezFArL+gTzmstPUDLgm0jJUplGxORXEpj0w7LBW3jt32/aTvt8IbG8gMKDV6Vq
vR78/AUS9/9k4H8MmNArgVg2HGT2kWjAL8Ci3THRNtodEJRj88RsvHqmqKeT4vzB
vi4ezOKp4R3jZ6zkq6XB4ltFlBptwd2l+7wCT5Jj4YKDV1RuOPzYuK90CCOg3xyc
DXSP8gJyScFAaEr6g7mfIB1mPDvMe7JZVn0jSjAsI7F3OBG7lAecZjNtH7jQnv4H
ze/yO/ALMEUzz9VlU8v9kTsrS7/p3nDVNLhQTQxO6HMcfp0bkcbD2Eo9Rxzt0vxj
6iETPsNoYcpm0sBCgO7w00DsjzuBxYF3Hy1HYu2BBSUx5Orj7vmnTwnfAdCE3faR
vjLHO/c59ktn0w37VzOaTZYhdubj4IpEMJ75UPqFgSjnY8SAMw94zoVPjkKn4LX6
fxqr2XRZnHi88U895b3nsCdActduP5Ljn6uXhMGSbUKWJSF7GvQIjtuQGweEFat3
zPOXrUBrLPXFfPEwQ/uXAu/yCKiG7wwCmhx7RJ9wilyc5sIJoqrsEo5oGUctqzLg
PQUq0C7oiXwQenXY67a+oiJKvJWToOOwxZSH9tUHy14MdB5RAxtRCBpKlCjV7AHH
H7UrNfyzPsY8FuspOzx7+2SNlNxYAay9kHm5ePrXABktw1eDYWKPdw1wA0gBaMla
`protect END_PROTECTED
