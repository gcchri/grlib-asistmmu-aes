`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jh7EJrgQPdi2LqGvzsz57tGM2zcEYhj9vO+KBngpELctTe43UsL/YJbiu9PUhw48
3j8XAr5ZRUMSmZoZOw6tHY7oe8ZGIp6+ukbsbgCCvoEYUaUWaqgRiQkPqZ0CubDu
s0jb0E9WcZTtSABlp1RS6qpaIrbOc9/D99V2IH91d8jdE9GhWP0G7oLoJA8XZd4t
sKFNneT4xdnFbFWRul+3+Bddivb5xp/K7HciJW5eD3K6K52aRV9/VTCj3KuYjAqw
`protect END_PROTECTED
