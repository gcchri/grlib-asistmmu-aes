`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BFtxMuQn+fEAwDLmkajXTWjAubBVYbiP5cc4zoQV+ROplF+4Tk9z2aig9JkTN2Fu
+Xz5MOajjmDhpAQprMNZmoEWFGFA1gQruSV2SFwMFhHoebcQzKhPhJbNUtaiqcXp
TvSOrygqKZMPHKaklHCO9epYnFlKS9+PTfqtOSpQ01Vwfqb9XHaC1LGEyQzF5BkE
wFF4fnQZULbxaF9Op1FELtA8hDV4LbNOh6Migqz7jSwFQge91Gln6O+P19q03v3P
ujRnctmkp3oZB19A0Foc8ChnxNxCCyaRqVwLHqNmm6cZUd/wp70C8v44RK9zk8ut
Q3nA/HFpfGaMPTnWHu668NZj/z+JieXTaA7ZtDwSEB6k3QWAVvvMQRxNNB6QZR8c
SIqv21aibula0x67K8ru97WK1mehPvn0WMR9Twvpvrlc8d7YmVuVSIMmkS3KaoSW
zgQsf2Q6DH7AWalq7XAB3BvJFn8u/7Qu+ex31oUgY/6SVa6kiPqf1k/4Yy0qfjxE
oPuBd6wRBTE97EUt76bW27sxM3bTcMmMZRilqpE9dFjIZXkiuaKgk4J7+EXcAmt0
mslBV07Wvv07Cn56Cz6faOr6Am8LnlmvzghXVJEyrAWU7376/KQHpKvwNMeaxa4j
j4A+XDvZcfQwZPz9ieF8u9lWkwpfsT04aogLsH6HCSzACs2zDDfa+nkPWlUcVVS8
evmAEacz6m7rKW1kVfG6HyZeWutu8ZGfUAoSEMWYnsvCt7GasyYpoDcYCEQRkKhv
s33VklWZv1xuW2g3PH5W8dCHDqj9B9roQ70emCNIAeGBgsmrSGw4bImIAGO0Fy6x
I6y/6P1u5Rz7OrXct9KGCQ==
`protect END_PROTECTED
