`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CRyhNC/ny28alWOQzkTEzTdnMMjQo7yhCkzGM6rXXexFWbYqToek66TfG5ROev9B
9wo6xBFRQCshEapoqHQ3eqfhOWRDWRvbf8z9oS88gqJjQE0x9pcuGFBqUW7zneC7
A215O382aMrXGY1YDHD6ka5v5k4T/W42CWqh/5C/lwHMuZmZ4fN7ayt9oZN3Jkce
Cr391Zr0BNTSDHtB2hunGgFfjIX2/tgLFf9DyjocZ2OV8ZfoaYo4raoHPODcBjeH
It023bTwV2XWNwgJtKOVvNKmhm/5Q0ZXrys/fQr4FfRwcPXN83hAnTX6j/IcwmXf
6/dmiO0AcfCtVfiSae00Mx8JF4A8u+B29Q9XxJhmmhV4KSdEd1f76nzvMpqpWFE5
tsSW9Dq8SL5mLE1Y7qKD2sG3UR5HrK0M6fP2tUi9g60bGuIw7dQW8XAsyiJFGOkK
zkKkOM54DsGo4bNY1xhZInhEZGGL0ns2qH3LfKtdhB6gBXuaTUbPk8nGEP7t5SxP
fhGTpVF/acMTjtNZJyEvxPGZ0W1M8z9XaJF64cGVAhb+JuThBVKJ6ycn17xvODAB
MeWzKUO8yGTKrM0tz9wUIYsQDW96nrrugEAWYUJ+ektAlzODhowK55+XuUa58Rdb
ffrk+xkVv6ZiYsN0uNW1UPcx57HTZcwOu+wmInQMvuT1P4F7XSywzopVt0YImcIE
tlNs714ouDfbL8j1psicalmQYWnjayxeTFm8IErEe+Q=
`protect END_PROTECTED
