`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3ajSc+ZIL+iL4mtoi/zkYMk/GtIrr2dxui+yo0md3qSktoCC7KnovSaBlTtkzuV
pmyg7HNSxBVeOBoxxmHP0RG8fB63Wf7bHjMhdb9005RJDRkS5Rlv8p4dbcL0NJro
VpJgQm18bDMRTwqQau0vTDCZ3jGQAA+i7DV4NI1llaQXSO5VbrOP+Aanl8PtwyxJ
H79/TIUF/mHQF6JsNK6WbbMQ+bfRb+i8KpMsdXcaNwiIAyRnBGpFn959iVG/2/IE
05Sq3+5hpGVoOEOpzQTIpvcxG5SeouzXSIpqGQZk11D34wnby6CrWYL1lgiyw+yT
/29+pG1pmJ5T3sF45bDKsT+GyEzqGxQxK2+FuHNXfNh0nJaHMcG6Uktn4k2G6pun
p7tL56vh4XLcfnXarDBGYM9PVGHPYooL/ahU7ti2uDidEIzc0bEbKglfpGsjr/M+
o+0hg+1OBhye0/Vo6a487BszZ1n9hJ6mcg7NO6GgxgcSHj/txF7TI1QMyr7PcOu6
EdQA1KU681xQ7P0WhZCJ6fEzwRZXMsWypeu7DctxWv8N/Bhr99zMJj041QXa9/gn
DTwPZKX+OufFTuoYiVPyXTEE30OBLTpO+OSnospD4OBBJccB7KJRiyncVMNpFrv7
v0775KD9sQuNvtD7fWQ3/7P5t3WImhHwjc20oeyIOVxi72qxezOU3S+zJn2viRXe
QP+2jVZQnr2EsIPDlb2yrXwHY9MGO2uCfuwcY8+VbXFvmHiEyzqldcdmNCqyWba4
770CRLOSShUNLaiTpv3wKw6WNmBS/nmY72spE9FZ8NwHf6SPxr+6gW4H2YsueTT/
D8ENuhk09QSSRxxkp/XcTWFXwH55nvkC04uWBkckboEMGB9sokYWEtkQhoMP025f
WA42IACxLc16Q+t/y6TMwDQ79kJ6/bIfG0UkjGF1sjymoMeoLYigtNOzKrMiTuu8
MB9BUWJwQv3z0v0sjX7gltnsc8v+gWaarmQn/jQ26WamLOUr/uhuUWjkryF8BxbI
tlCyUxXI3vkEqyg8qzhYRknl3JGA1FVM6sEf6ZpZHSBEuQmIj79FEamfCPa0/HcC
HM8SvB5GtrID8rN18LYpk1FgAl2ZI3CKLNNLC5fTqcNn1MYoAqcRkhTJjYrEcD+j
YptUrd478Bg8wle55wPJ2xJGtZN6wb69bVe2G4EHesCyl0tIjZQJfw/GAb+QoeXr
T/i48wDC0pnAG4R31lde6gNLVXQbfMYn4Gy5+Ff6NHcTPmBSY4w1s97zzShNMCCo
Q/z5FLRxGQUTiGXsO+BYYH58WWXVMTVC8y5DucTkSpHsJgFF1LwX1aNu3YWjGxuz
+H71bjZDLgt4IBSvqiSjhJ3Uc3GHWAL/g1RN5M4YiHCgsfPvYMiopstl/UFgVzw5
w0/FGpVNEG4Zu9jhLxwMUfbLg9qxtsqIpjvFlB159mHKeAjuL8bBE55qqLPkbD7P
7Gj106GZ5PcrypcNVw1q6znCPikItP5VnPs3EgQ00W6lD4CFiW5vjjj6sWAV+Ekz
WSCzbVIlJmxEWXFlz3BNxwrC+YONDFCBMol5JLui42fdUYSgUO072qBkYdyo3TCl
GaHuuUsotcPDASgxh+rxxQ++u7feHKxd1cZEWm4k+l9WOm9YBBS1BwFJ/8Zfjoow
pfjvnUZF0wdoXQxgjeF21ZOZdSCofa0xHLjqvPJGn7l7ap1YhmqqaH3OWHrOQb4F
MLieNOcjoBJg3Gan76Duu9dvzZBHZ3UKaWyokIQU4B3UQpKFBLQ84A0cig73tsK0
wgAh8a84hd0zlX64+r4R6ez4Zb4QJFSO2Hzd4PNhXxLgJWDQuYsez0MbrrhMQN0O
SvG+bh9D04D8Z0//3OokFEY2SWkgX73KNmUCUFAzVph5Z2b/bpWYUUzIo64mj7u3
Y8Yo1PPKZ3A90RAcOj7wddAS3cQ/JUyPeecQMYeDQ2UHlP35NDI3UbAkQxf6Y2h7
GPuudoJs3jNsLN8vxziOf4FDWQzDkq8C6ctk2xL/nqYIOaC5hHkxPEAB881rGwB+
CqsilfGtNTr1JGkvYd3SW12Vq8+1uGJRnIlJSanHGoL/n8z7SGx7/WIGFv6IXJ5E
QBQrVQquxNtdiV+bpSjQr1xI6nGuS8yDL7qKuMiff9rZE+fo9YNaX92BHaexRefl
fbqYYJcaClzBtN9PSiY/KbVw328C4JJWJCEdWJF9WvHrEkgsSCVAxSS4sDzuChxW
t1+fydVTzG6lEyPkaiMNNaqOT0q8fq7/Xf9PGRRJjboixoKC101lu0sOVSuA18GP
yjZaDEZMNk2j1gLP0jNeFs9Jcsoizqy2mmzVN2OkpjvSkT2QXzaATmJiUoBcFLdn
sFAd5jgkVz+H9yTTzAX+n2eMeUTwYr03mmD+2yHMOw4jCTAvJHQ36KTFc3OeeDHg
XlWTDUWtFqATEiZI31hHc/WyKHJlFV3yWAPVkbwDcW99/qkON250HcdfUrVOq8uM
lHjrcvAPm1uJjZ+E3xKVhzqeU51dVsgIFz1NpyYlNZOjIDX+B+kowio7Cm5/OIFv
7bI30ltVxaZzLCrLiLYmFMBrQry+1R6DYFSQps+uHhEFgVu1Gectm9pC1bHmbjwD
lqrXEykLc7ihNQ7o87yR0XuiE/6tZeN5BGTIZgJ4btMqke5Fpj0rFigPoUJr/f9A
ZWO/GekD05rKmZd7ofr1Muy9EeXpSS2ZFbKV9FhmD7OTinFTPIu23riegfcdvEjU
MYnIX7dKWsDLUWzirOfJdoPnNWz07CA9aC+QtUWCaSkJFs9OLlON8HHwDci+nAbP
Y+gn6SGZeVnOkAc3iedUKTLD7Nbxi1qRlejAiTCByS84uZH5vWXZMSfBf9D+nyM7
Qm5BarrKZrV9ZxCsP+ucCcLrJytEREEhAglCtZIvHiLo10NAK48oH7BSzxRCmB4O
YQIGOwGvJE+T9WtYAP/2w96R4qLMWHC0vxQbuh06AD3SgEvLLd8aim16d5GY4q70
sWIJtoqpFR2pn/lmpRIOjJywiK3tdanf02JfubV22Z5CXWYna8T4b4zteVimsQwH
Ebu6Q+7/tN+j2+LBNH0S0301gAhwzhv4DKcXYyxkVVVcYIiu8dl5W/VvErS40cwm
ReK2NrlWV7FY3Gqsq7YCz/OUQdwy27BIh5bElbZFLPf3t5aARM0ht1Dg7Mxg42Vd
Gl8yqlSSANW3IG2WxIrba5rtce4S0lO/TcOuxwp0Adl1IHZuthxXwjipsVxfNeGz
YKvxI0VARW8i+kmpOa6kpkrMTXh33LWt5t217INQOtRSZgJ9DkktKfxhC+SiJyHQ
HeBTSMEmL/vaLsRL78pfb8VuFLrVgwmeZsn/hTkhkBeUtiY13oTuEBjkuH7E6IHY
BYJ+rLpOpPIuhBdlyhP6ipIIHPcKRpeK3Px7nmZkytSdVLA4WFZ2c0ihncK/6vkT
mpF+hkfkH+YyyDoRFm0+d14j0Cf6YudxdOuNfCR32UhBCQtG8I8dDNlcSpTbMsgs
9bGabAaq2tsVvtaC0iXHLQTr/phUt8oiBt3FifIngE7Mj1vNQuGP3eqbpubi/4Sm
x3Fen1X/iYja64zg2T5JBAldurhEbbBpRZgTRTyMf9HCurNlkZMRSYjwyyJ/+Kmb
JNP1aYwj10vdfjT/O0aXMfbkLn5BZ3UNxdeH74qfF5Xf9QQW/8eGU8WL0Tq6Rpd0
K/R6mr5Y9NrLb2MNEWuChDvtX0Z6L/c5JOvsH5cCcWJdvznbWr6cxQ/Yj/H9+UPP
9wcPawHkgLJytrx+emenVgWLMVoz7v0wRcqPo4oA3l5dJxdbHrD0ZuSGPdJy0HXz
J5CApkAzs5rFauu08lmAN+Rsdxz/r+dF1MJ/Cs9z9r5y1NPR3BfAka/iEczt2ckk
TQIllk5K931NNirIyxhKvz0m6G8+DDOdXyXgRbjEzl8mvocCoXTe5R3jpG4pbU4g
9PFd0D1N2MEJuJXouAsB352NrFapYyWPI+tOXfnMq8pE2ur2LWzR6d7tTYiNKbjw
ARAjaYwaWfkRm5tMQlyeVNPZFOEsGEd7K8cw6rpPFv5TxJsNt+3kHEa0npZYsvmY
8YaDxg+QwDDq1BDTppCgeCr6jXc9VDalBlp3eahtH9XQEf12qkqCurN3ZMR+90MP
nVg5ssM21AQI5dkgU3hjn+dxF1Ip3twHLg5Yo/sDMGHEDlDV1ub//j6AZvE5PV/R
bhemEmtSsieZ7NBzAGxrbq09bWvQxAlNPRa1ZpS59MnMHb5BHt3Z/lER8SLbAgOi
CNyMKnWu2RW8ypMo2hJw15T1Su3AOuns++Sj/SXqtymUgWg7FZBOlO0lpva+JeDN
/rxAoc5AaIoQk2uAsSsx5xuGfNbB0RMpLkgwWM9mawgPM2CaMdHzNUCye83yLpa0
vNqaOcmje5ITe1dfEIwLWn1pg7fo+XAwV3PYyDfmXxg3p6zhD5HgP8rapttvik2d
ADb6aRi4Xrcnadf0TWacne3VVgzyF8SiO2L1BLBj37g=
`protect END_PROTECTED
