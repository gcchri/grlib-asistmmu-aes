`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQ0y4UJboV/F7EyejmvYRfMjZs5Lq62YCppqCcuTdZtzG9GJcDBL6YxC5Wy+mdWv
1HTaoKhZvl/V+p90Qm9M56BIMy4nyhajbqQ2I+1+40F0ABasGv6gInmg9PfaBtgT
TFL/NvGJMXMWb8J4o/QpIl88vKDdVWZiVwnZmfjwNObi30Nw27C8HKyQkBqhmAH6
4NBr/4j+Xu+wOZbdYavP+el0VQ5d4+oguGDHT5lk6BBk6/JYj9npa78QQu04Zjuz
1zVHlOeUBwnR+EbuJV1wnSy09T20jDr/KwbKiKGWE4nHicci2BDhmsMquV+xM1TE
NN4NiKnEzUDGyPyXewgmdFyF8tLNw7+S2sgrPC/SHFdoVf3G4vWxJBrFMCpwJEEa
i9c/D7J+kpJkju20MpmV0FssSUkIZL9PT2BoMIHNWQkgR3di5ma1JOq9J4i1U9J/
+ZQCitguRtT5MZFSeT3jbZ0KodvSPoMKspiSa93niUL6eK1ac0eS7RfkATkpeNgD
01D6k+OoScnhP7oRsb3kQQ==
`protect END_PROTECTED
