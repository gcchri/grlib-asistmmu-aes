`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vwyJw8MRDdVRuZUT7ZUgoMiznrmLQIcK4Qgxm132COCUPxN7tR2WO/Jw+uDiOxKg
DV45IoPZRPdqmxw4u+KxsI3E7zSTf/fJ5qBU6C1JpsMYk8ZykPCRk3hJJ+eK6+F+
yHV4az+eem6q97Eg2a5/iblK3j++1qBTMJZoLOucq0ZvEmG5i0KrE7Arjh669+jj
AlOc6PfDFt/govmSbAA14zk0b4hJvwom5I+dq3bfZeEC+jsGH1vf1o4HM8YbhVSJ
6kDQmZb0f2nef/Y2FZWWy3qCatAocNg0aUoUE83HGqetuRndqZSQ/J7wQLD6ghFv
QSANNUNwj/+5ylpa+Q9B+Ry7RFbb1G4ZXj+SpdcHA8Zvu0obZB/Kwk4NeeKMDXrm
SRSMYyWk+Hj9yJ59J19iomLR4MsKQ5r1NGOdIov0DaUp8xFLZravSe9VOTWtPHKN
9UWO/X8MfGl9HZGLcoX5rKDniHqIiTqkxKjOcAS0+Edx9ng6E4f8jhuzToos9Aym
KSgwJqPy1B3hQTGNmUjE/J8M8h32kbDZUVoMmnZArfejy1cABdvsirDCdbKDILaC
fgbXdF6T+GGNVHbWRzRCndcRQbnmlp+2O4giZyNiHgVl0levTDm28i5LKNs760l9
Ds2tf7IRQH1RlwlNy5QHobpuLSbzgZNZ1JZ1FsMkIcUUZmzbAZH2lD+DQbaLcGrl
`protect END_PROTECTED
