`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jvXmFH4pEzxebjwVR5tIIinlXAoPayqKrMdmhqU/NDv6dfLnLrcASv9JwdJNQIqc
ZlI2CEuj/3lmvkc/fxiW9ysq0HoEkZK3OoT/yFm3y8mcrH452FBM4S3/SC7bpHDD
q1v3JP5CxmaHExuTMTMcF9NZUAcq8t7NNrEu0u8849SUM+FToAwp6YF3jl0kOgmc
AISlvnCnk2wI1zBJGrpoMqoUzOL7o9DW5U7LtVyiNJDCrFtK98nx5P+7cYVhEUuO
oqmm952bXMJolmzsU+TDHUxUwhkDAizxb0ZkrQFfiD5dTrrT3jEHeW8ZL+hhhRy6
1ZLXkx7bH4BmgZZRdp/OTXUSmNyj1MwzjGG+PvWwr2OqaEwFIqyFeQil3xrefA2o
vUsSOXe/607busEsgVWqhpfTm7OfDaT/103lU1lzAjLw8hRGN/2vI3XjEkknspUB
2QmNp4aPZ2N7OmXF/xRL7Q21nSbksb7GmyBfCwK6wdQo6PUjOJskR5iB7fh1TBC+
1LfXPaO1xsRBw02I20H2wDp1dn5Ai2HJRIFxwXdbGCZUf1DLSNYAK7L1+p1tqc6n
KiztlM1bjQvwLt1L9woQYGkvbjHkdM+4jCNwHGDQH58bzqU9NwTP1wBTaMQyM/m5
aXt7w2CTYD1LEkL3cgVbUqcXq/xdTvcxIfzfa+Nb52XPnGHjyMeUAm+WKXThxtFV
Sum+EQVKMfXzw54F2q5AWKXiB3H7mn57dM4JwAARpQNM5+IdFJBXjBSQS6r18+nz
Flg94WX/Zl4TmNxjzQ++5g==
`protect END_PROTECTED
