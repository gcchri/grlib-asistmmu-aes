`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xp/kPI6+3P7Ns3T4LNnrT+9dvmtBBwnBgum4lg9NDcUHkhPF82Yt0MXRo567tRZb
sFJqPo7sQBbcPXYh49tr7gBluLoMiNMnmHNaqFR75gUw+RszrbQe2daTtAecJQWD
Zra1ubOxqRC2zTwj0TcuvBXgiZT0xhNc7/LrDnPUjAe4e19r9RQqaafy2nOs4GFM
z+SH5GH/MrugZXJK0TiM5aVzhT710r9FjLWOuqA3Q79UEkcvx6Yd7WKj8ixuMFB0
C+goz/B3fYlZHSziilTY4fuv/V2vqTU5iolZ5yadjDnn5mC24fDv/j78HxyaqYPZ
B/cSrOmt2CzQhN1o6wNaqd6MuM7T/ksFECFQehGkmMqopg9UNhQLvLyRj81kKW4z
XVyT2WUVfhuy2HXqvv2pnkc2uF7u0nW/sOpc/ijjpy+8Olmdl9n0nmmg/pGQ0o2O
RysS+inWeCP+0bZjUVe1AI7lNGUCqL5nG4rAOhRrcKslU137JazZVDxXEDAFMaz2
Xj7lf6jCWkO10ydCUN3GwOD5cGOrP1gbHhb8AMW+1/NkV8nZ9qJ7Jec+NUOpaeEX
wg9tmm5EAXxxUlImMuzW1i0AgVVg0JebG7l0ZDUI0ZzAHl/lQ6iHde22bf1+AWQE
MLW/51tddEFlZbLCsAVFp5cxFIk9I/E3W1nIFSS52I0sEw4qFzqYz+A+/osjHoII
A8VmH7EKWBOtjFtFa5dyON5IKEUlsxUKgEIOSoJ3vUwPE79BGZZQAoRjymH7JOB7
Afp9mhOBddGbaVWo0Hn9TeNeRNslpy3Z64J0bQmgVHY8vBKHQRLvfcqZagMhquBC
2leMUDMwTAD+X1s2jwH//aOuh8LrB/6qkvRO6RI/VLBDgm7wkOAZQmBP+OthOh7j
Adjx6+qrLgyHcHu/RrsPk2e96g8s/oTZxNYqUO9sZgo8rq7+0Dg4THpvFAL9Yvim
fHaGbPSlZS9WBL2zaRkR5ty24hgZTUrLsFjmhm8rPsc=
`protect END_PROTECTED
