`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Mh92cXX+SY7BSVG1qkdT/pOXyabsMmLB+3MMSuc4iOTRMPTGht/PZi6DKzi7eER
P6K16/PJtH2yi7o6oTycLrb+mjLLlkwhDie0tnnHChesZLmso3/XCbx1dmLBubXP
p4+3XjVblD7YNNE4KRtnqGlhPZ1GPIJJEiEBOv4HLqCb6+D+fDZI0oIWec0Ph4+T
tbMzkobjU7uER2B5/e7qWk4QBN4qLQ33/ROYatTJNikrZbOK8rPo8DYq9IFBm6ux
YsSOEnSK0wowuIJSfUKNgfeEApNKj7/XAlTeAMcpuorzNqCd4jfWYY+fb1aT0cAj
tDoYMVvV1bQCay2/C5WaG4b4NaCFoO1PLWWtFWNr8sXeJPlxnBtlzwnWyxjkQHb/
OuNlakbRH8+7QT83CkeU/VkCScjpNRWWN+B2S1xgWGPb3BX4BXaZ5bN8zc1fMhjL
xdvMeKKcbpCIMCQ3aV6R3rAie0j1HcFFIAaStIs/va2Cgjc1U/LcCrkJWA4Ms7Uh
TaNa6q5zvTL3wZz6PGFMdoUybn+DauNoHPLnoZ2e4g+1sGxhmjeEoW/Ad5x0NRsB
FbtL9o8K4+eqZoOLNVNETBHbCzJmGJBaSLzekaGn52hXN1WTpugUGLqPJ/n+MQME
O2ENho0B61qOA5oVd6r8Kg==
`protect END_PROTECTED
