`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z0XB6my4OEoVQHmSaf+H2r1oLE1ReprFUxepjqo2RkjZwmmPosQCfT06tRr1yaAp
983eGNjAicD7EZKRxubnouoTZO3HbFtsWcpqPCsdgD2EQ9DdubBQa2TI9QaEFO1p
RBDjmOUKKmo0ZMRUEIohLgfahmllCl0MVLypEksygjsxGxsQrGShIcw/mFlfTFWh
94ksCgpxq1jpP5i+Btrp2Trt1VX6IoGyUoXWogVuAVSUFK8fATHb3FFd7zFOLTem
1PygM3G9F9VO4I3r0JiUhdtqrm7dKR/DWOjOM3qxaE1STtc6OuIPp5bc1O0gzO2g
72m669dTP5UajQ8Ec3Ro/FQUL/pgODLeTVNUk762M1Q=
`protect END_PROTECTED
