`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qiMiMJ5Sfy1pQtVrcuPGMnTAuX6hxfOsWm1lQcsuYwbEsUQb9GMSEMKWby641Oyz
ZAbtUR84RRv5WsuMAMO4cff71L5TThUexpho63R87RrLjfUn3UExdwcUXR9QJrNK
3rFqDCiNuXugGng1AzCOCoChcUvKVC2PnB62v/lnGgp8vQbDtFice5Gf0hzT6vHA
4Ay/YaOsocP5Lu8DdldisT+LEfBvzJbxekdEkw/eN7ksixqOsN6OtpK9OarLT0Zf
lbq0PDBcmfrgJxzQ3zfxMq3UziIjrYQm3sqgsNPEu0OLKyOSfsiPMNFNRBSacvXs
af9O3ZQt4E9YEYu2RpQaJqiBLyNQxiOImUKx4mQ8OPjtNMnd8phYF81Jca5r7vpp
aJ+8HHL/6cNZtOp/zKMlOb/xH5VTCjUpzT0tT4wyqEcfypRKAk+vZIuyTZx1FMXD
V/ajBWcyYXHDwnwvNORdPG1mOYS9AOpHLYdWH903kb34cM3ITbOQR7c6oxTxhy2o
JcW/ONvseqyR1sRTlCHijlT10+XsueJfwoo3lkXEkx8GNEIkeT5YhdHn+CFHP67C
z3xbWFouSLXdqv9Ry4IZpfNsqaSdd1S5EG+RSY5N955OEz65NvRUEk/CvVKMRneY
nCsh7kWYh9aVGC7qAplyHcogh+VpFnTY8KzwvaD58bI=
`protect END_PROTECTED
