`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yFCLvfMhwk1newNa3HBD7RQ5KDC4iHi2tDexnYzfWTUWrJxb2ahE1Me1i8DTzxxt
iZhGusE9ZuTSTOfg7QabasPIVfzjJTYj0Pn+1v5t2IGF5r1UVr4KaXm9oDo0tc/s
FnYNrURS80p3TaDEtOdD3RwILnWAXNh0WrLLjIPDeNxQsU3eFEKPxU5ccrUA8nnw
F9tvxduNVIP/BQ9nX5rFEbJsYex5MvQVA0PJOI5wqobFeGn/qr5K3WJCboWu+KQY
4GdNfUB/Ek0VpiuCP90G2g==
`protect END_PROTECTED
