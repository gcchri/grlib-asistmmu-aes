`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
okMNlzfoUsEvVj7W40JYETHEGO7hcM23u2co/paPmdYV6xbzNy2PCxBoCUDgd4vv
MzA4kz/SFwzadn3MwBkeCcUGVrLavwVeF/QZILcScN2VatUbUMB57WUAimmpprGT
1I6uY+kxWp8fC32Fpz+8AE5eLYMtg+FovGA0tKN21Ii/25mnF2DBXenj9ngOZtSq
SynUiAIpGICELGm7RsyK9fjEPD4BfdOfDjXjICyf81K0ej2EFAh+YXlmYm2+/hgx
HqaObT0um/QYQjJWghPk2M3253Ppgy5U7JTFBrdVDxSixR1k8DqTj8qbflWFnMM9
d2Z/dek/XBqMeuFOzV3vXIsHeUkoW0DbR005tawfyhKjpo2N8TOqIHUGWL26feTF
F3PQz7py/qvhdBEzP2vKo9HWh1PWTz2A4IK1UrPVt4c=
`protect END_PROTECTED
