`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMViNI7P7eg331S8abBr11Ar8Nhxw7LWvKNiJ/NFFu/i2s+mzuoWsVbitoYM5BbL
E2ka87IaUxN3RGNgJjzFYYwGRcEbbN/W0v4rJ4CjsYMesOmRjP8ucWawNtOV3RWI
p7PFUkTFYWBGzF7+yrdyvanp3iRDCRiffwvz9jcCLLsNdDe8FvpNsK9fvBkadH5/
5x8e9ULvEgcMaFiZLdbX5XDqe96kFyeccnW4pfL7zsHYyOK9UyWA+4JKDeS4yThg
McSxaOxPXfEYygPz14DFgSYqSte8J0hjCU0QcAd/9A9WH7arAkuMcYnsJVvEckpW
OHnaviv8tXbOj3l/oU2ywM6/m+XMFpu5lgmZwiR2E7zyi6rnLmz7PqRSf3JMlNEm
ZBJ3xRASBttWgjNfPQd2bskkZAjVnMcy5yKsPKdkN0UBTZpVwXTAT6XNIMQBn88S
UUrBB0cc68XzNfBw7WeEECAKm4+zGPN4ZrzdfbUFS5m437N9YHVB2jVCyURvPdNO
Igbrki8x/++PvhItFrs44Tau2tSeK8J7B9989tefy6ihaeDgR/EslWIKC9onbxmt
`protect END_PROTECTED
