`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXcgfdf5Q/Rs6/uYK8Mr6SPXHgC8WMQtgLoCDLB/Yfef08cphjHjYS/5xtT3A3ow
8AmDCdX8GP99ZNjb+1OtfGpE/f/z/OuvRZErmY5sniJ4tWKhIs/FlSeAkE9dGFYK
erXx/R4o5LpePe+fyPaxLJnNMwHAmQpkKVvE7mdRQ6Z74MfbjRjsDvhFDZW38iu+
kmkLPzch9o913xdde4/Eji/mQ6SEtTetN8xhKXtsbEEdHgqT2p6dyi4LDdh6X4Ue
p5GbcyCJ2AzXswCCnPvUvRehyLJ+b3Z62ygB+UCQZXhVskHWdJ0jZZTu6h2EtCio
/9Uz4QYIPQaQAednHwYA8bOXxgWtdI+NOjnNEvrO9nzKoWaYlJrg3mak/1vBo9uw
ARL9hGoku+dnFOeiM2eMNrm2Zku+jL/CLJKmUfvSnJ96Af1V1oCr8Ne/+1etbXLU
2SmRMRIvr/mAIuXTbviG+3gLDF6h0WGrKqTIr6ODyuXh5jTOGRuDFyY/UWhrwfj0
cquyj2JE1xSSiEQp+xR0ukWIIx0AvRq+0r0vBi7gHMkFSOPua6xN89b6rxzP39Z9
gAv7bHn1XRsgnmHzJyWQ/Ks4B61gKTgydEWYtb1SMZtR3qK2bvoDKUos3ixwvPZW
mwFZYWdZOqO5YJTen71BhQd/R9aQZ+QW3CU47ueG2ab7dyHHWLj5/fKACV6+/lrS
2D0iFpZ/Y/+FModTM+k/p1KdArrM6w9MP+ioi3Jr67/z4oGw3IeKOTDDd4AsICww
K9xS7dT3Fu7oAjtNHCH1zrtTgRBv6NDi4LQNHLf1DpzL8x3RU+o/wvYXnd3gcpt9
eph769QNI080fsQ0yS6Z8+4UqVbiai6PW4Kt09/qJ2fNJYpPb8aB4/P7kNcs7+pO
+fyZxq6L2KUr3vtT7z0iybEgg7674gT3FzTEV7EKOXfT+4Xq/3xlUcEbm+7jBSSb
8rEpPYG7TZVfiUCagGFznp070E3gEP31D5SM3J7zmlTtR0KbwpxMp0zh2nMkqD5S
5Jvl/N9a08Mu+LuTI+W43nvXJywQ+zDC7Gt+Y7Sh5L6OBi1DtXfmpZ+0cM1GT9L6
zoh910sDEW8GMKst3aco2c2DEZaYlnWobVruTAVCKNe+5mP1RMegXZ8yvrFZra7J
JQNenX4por1V+vs5cfi3F3mb/SSHe9ReqB4j36SShDZCH6eoo6NpGoW4BavYdp7b
NcShO7kr4+bxv2UMXaTiYbBDsg3BrA0Yo17qfjJJTSDLxFCD2oCBkZ7nn4BTlbbS
LtXZ/SYUUf2niYwrGMDb29PLGeeVjK0n9vJwX26HIcZgj1f3CDKdjnpE1igCuLjN
gfcivLXp1G77tA7bXM7epA==
`protect END_PROTECTED
