`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AOFHGwWDYrnRYcsMFReuVozGssIXHRPms+yPPp33Cn/xsyavAtuwEm2FV3Rf55Z+
PM1eq2725LaWFuiwB4+5IPtiQ02eF+r/cADRyiVc42E1EAKAyHFs77ghB0zsJbIP
4RFeL8w4sdQHFJ+RhUo3I5aZh2i34VbS3A7+ZEJ8uUFdOlT7FATAQRLnL5HbD5K7
AsFR80g8aHFkHYOF0OfU80JNhxQRAshturd9DMN9ju7vUcur0SqIBeYkWKZ70vXz
gYkFo0McmtaxhBkNiHfYSr//HiEaiDOhEwI55tztTWxwqQ7dE+vyNMJzuVHRimMX
F0DjrtbTJFM8TxhW3UsHpn6BCAueKx4tkR01YhKw8C/VeLXaohmAqSvWhVACpBel
5PnKHJkqepjO8RzBjoGDiAfolesrWQ5nad2L4ZyDn3P6xQ2OuidmNZDU9zvBO9TK
L7nvOsNzEOxWwx+Cp09pKR1XjxL2rWayrJaWRuqgx39lo6c8ykIUu2iF7aAtB5u2
cdK9NdBNGl+N79E6ToCeoU7ydjnaJYiw/75qTP5Z5feLn/NscgvU09arp0LItaCF
`protect END_PROTECTED
