`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJb0DVH1LOwNXYrRlrFqoI0+1tHXB/K2cu+Bsfp4I0VU7iqSxNzlTWyYBQ6EoDnn
kaqJ3S0m3JfqgR9hxCcIduXkd16FR2iT+Xlpfse9EVDQPBg9YRgEk0Kvj+gP2X+e
iKzAFiVkMQTnJkrlAcF1uy2Jq7nIGHuPfu+MUFbdPRaPUrFlkCr4WRPmrwDzEIhX
ugUMnjjkyLZYK0c87ZA9/k75KIGZ9e7zj3gYK/Ac/3xXIZd5wLUWQ379NocOFszJ
gL8XQzpKR6o3qkYVgn4iz6lPeoLBd3YapxVDPsimKZrMeLZw2MYqzTV0XfEp2s2I
GYhypAEi2B37+aCztsuxxWYvFMv/p4SUsq9I+AFb5AQ7WWboP8QJId5/r27ZWJbd
xsXJwxIE9HTVmQzoEt1DtA==
`protect END_PROTECTED
