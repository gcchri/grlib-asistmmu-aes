`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjrZ1WMfzweiPTNPkcOvh5gyULAkLv/j+HxKhTSX2D/5IMxNUnZW0io4hutOEqv3
8TQgi1EqOp0nmltuPkD5BxbtYo0ELDqlPPvmzBqix2SBRzuOkSE9soErYxveo4DZ
a8vzAFjL8mIibngTDy8q5IhAJkVykzu1oT9pZLxTs2hXQ21RwaDdk/ipnShHaR7R
YYoYqIOSuhSZKWaWHMKBY+rrfmKmaBSkdqjUzJb+PdD64T7sVSKPi4hOFU/WejTD
pLFe3HwCArxxhTLAffyxrlKfmiPe/joFKB4d/ZyQK9ZvhZhpLcxo+l+/pZOXPSnE
352CKdueAj1xFuFtvKqZMRy4u7RPoj7j6B79uW284IbV/qA9r+s4ZaBB72sovnq/
YF1K3Kfuzeq3xALVcycYgOfux18/aAc8EjPW2XOfgE8Bd76z5kYWzm6YUWqqzK2P
X40IowAzMG82YkXYZnqvdrYTGLSWO7pyC0eU0Tn35S4GKTh4e6ao05zcCwJBHf1P
a/+9Scb/IQgo9n2YKcci9EUVmQVdKxLTKVPJe091Vv/U22bCkd++UZy9od9mSgxl
o1R0d+Nl5qqrSWuczBivvqT5tlL9dw4mv78k+7L7H7PyxaiLpD+wOgMLVosdVPD3
N7PWTt4F7zs2SNaKkrFTicMVLZbnt2YRccYT8AbbXADwF5RRqN/rvaW2NhjjX6z0
4JEfLmG6SOFcgzRpNpJfFjL6l5FFi7/B4iqYi2KxUDYneBS8mhkeWWcaDqsJp/xc
Ri4B7PLbcyyn7PpC8L6LF13FK3xiR3h6vjhprgZIooyUbBzbdR8laYpAq8MxlzIE
5dVWDQOlgPFIYy+HqzG4XVDJtg7WZWgB8tS/vNps8bgJzOQZDvaYm76DUGNUdSEW
I7xMo9TRM97U6RrFk6ECO00u6PSXbTFyLwFgNVhdPCl7ntRTERqgIvftYoPmEPGf
qco5PBJN6KNDQwUemayvWQ3vV+bjy61FHKkYMQbAlyDXSFQrnk9guO+4MZQzwp9A
c/nQjp9Obqoa5QKvWSFuu4kB7GsxEFeDwEAaz+pgLC2SSBPXma7/sc3saSujt7Y/
mdgBBbFekIzhOKpXTGIHT2MLbVMB7GU9pM/B/uFlzESVDrKdSw1TJBWpyfKEdByY
QxoU4q5VlPQ2yIxLsGXCzGl3nDW9bT8/0frYi7iWCiQ25tK2TlKPmhuaE+T4pTht
1LGl2tRL9dLRt2s3qaVFR4a20N3tlcQcSoittkh+a2AWnyBfVsa/sPBLZ6wGamqX
4+BhSx/l+FrtzAsksk3lV50Z7BxIjxDjLMO2oQnY8koc3lASbvgN1wN1hcpwFo+J
DQyRR8eaG3EM/1LRiAAZVSr2BRtEq03Ifdcz8uY3fR4/lPqOJhz78tFBu+bpGueG
MhGRccmHBjsQ8t0e7ZO2h9EsInrlDWBdaOdle3JzYPxR9FtU642WU5flA1qcReqZ
aSGX0rQY0wlTYwnMPdhFdHZtcS6QK6tCvdbtqoGrFL+PdT74HjFWcIYggHKak+cS
SKnXQZqqSZiGTwjjAKrfgEBXixYlv9ZdY7IQn2EaL3Bh4vhpOj6TtEqXcmbAMhaw
ctZgrluq6DcY/Dc0fxV1w6OMl32SSbI0gWTZnQkHtGOfsW2DjU9wkPEK5WJooEKe
hkkgFOs2TyvO50cf+LnoesqIGKniRzI5WlFx1it+A6dK20TKvi5/57szME90KIAR
Gf30IqJzLAtTWEBI+uIdwYwNlG1OuV/UUVdsHGjFX7Splvs9Wki5YPfsqwIJznQE
IMIgY8c4Xku7WIOPVa5MVXTP5hNrUnmp6Hu7tTt0ACqTXVAjEL/UQuVrDPGHKkGY
Vgr4UwrLe5TFXFPtoGFULVzqBBRB8LwOO3+AtdZcuMCkUEfvU+vJNOL33loZt1hQ
boSVTnhz3LOmmueeunIwQPBTCjKke+NEcUNJcR2SyQu8NdXmHdFnh3qYe+Q+PzHh
s8fxq7Cos9VvM4qxymqrZNViVtvpY6xchLNmwA9GL77AMiHJOhgWmuDV30ZhLeYO
9tNhXNzPf8qkaOQBCrnSE4nCzN20Pq1EO3btYZS6QxyvmhxQRFQuPrYriUQn6pA0
`protect END_PROTECTED
