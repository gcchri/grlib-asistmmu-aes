`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2BI9us5YtyYiEzKMxneYnhig4CQCqIAiuTJZAK/dHekkDR7WYzNTdLY5hi+hBE73
4ebHTZX9LbshZwTZ6dY3gj6+8bK8nyI5KpqcQW+4YlyrN1mQCrY+YxAQ0ffExEF4
CIWpWyVogKNHo+Xf28rTFKJn+kVx0GRS7OG5hvEldCJYU5WHMoz0xSuxapGCmW9n
NCuXkRSSGjUQ7zufI4aZMoG4fY5vpMefAfTw8Quxzw+DFBa19NjIslBNU/qQuYaP
Dc5u9XlrBdizwj9q2qyHzEd4+U8azJ8gJawz2qFZxhCndLeGjT4XSIyLWcX/HTzl
LZbgE64ZlZ6jMeLVW4C1y4UgfYvj2Zj8QiTlhUmScMUc5lfevxWmcdpQewHmUhgG
80tMpSWwmf8ikBYdw0dYUA8nhDNR7CNjkBuO0eLWCTF5llK+w9c3Pn0n68R6C7g+
i0FRebX3Gdegabmd4Ay8cBpd+pw/VJyr+7YzQ2A/ATz12XkFSI9XQAlRZmwj4DhU
d9RCjqljR7S9jywKqsCGQghVenQykCcbyYcHeF6DdNASrevRlTqgUpor+i7Y62Iw
UMCVqqYkMnU1e6k9OeLKswWoH/GP2mSttFnz37ICu4ypXJ6GWyLU9ncwx2ti7ThC
bVdtvzzGdYsf8OT6rPPEh98eWqannO44qhRlqKzQMCuHjdKGVVn59ZrIqBtVPFV5
0oYg9X5xdx7p8E3atwLqr3w+sjeIszZ0IixeiyG/6wY8yBvnFBxGdjnES4M+JuKz
z2aFHWGof568Bxrrfxz75l14slMTCPqqngpXnrjW8nOMsfPXqIC3kn7nrJpeo4tY
D4bKdLMCsjcsunNCWYCu1jrELbPg5BWgExTBsTjcTlo=
`protect END_PROTECTED
