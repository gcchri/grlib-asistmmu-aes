`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQSydXFv7/qdwKr7B/8ODs/Wz9iPJxGTj6p+lA5TII+adJEoMwOfuSXDzjBt8SYn
kFnkE+0jEvl58sshgeLhO6JCJ5j63MKrqGCd6F8aVyzemvgQAWNY7Cv3qpQtwfVr
6o6ndDkj+8E6/zb3V0mUW8wJPMtuTQpCy7oQDSIZjgnNCt58qRQWAzedrvwlGQ6Z
SaVRNJ9BeTfzJPtmgzY/wb9D15Oa2pe5Sy8atNmYKnIiwMOApwPyYmbCT/fzbdNA
OHUhgiudCBX1M8De2mDuhwDSPgQbBmu2RoOHPxscZiEMaRvnHTQ0LAfdJ7qoG6w2
4dOol1dbjyyvePWDoBLn6Q==
`protect END_PROTECTED
