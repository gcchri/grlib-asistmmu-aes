`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xMP1Rvv2omymkkYVntfWecSigw0KxTkEjhHhgQzF2dGWqF2Ansn6UI7/O1RG42WF
Hh31g0oMgFoZ5xWx5vXrywyet/FApthTbPfWdqCi7l+0iADgrqcmJ5GF73Kgghvu
XUdIL2GveKRmp8uRzjxUabMRZhmClzIctdsr5UguBHsQelkezbNuGUhzgd/t8GuF
M5Co7BKM/8jRX2cDTmsUrBxPr/x8JCOqcjTSoQ4x1mSBpdOy8insB9+o3iWokBhu
3OFF9r2az5Phm9p+bIkn3Pn3bKhY83YzSB1H9wC0Ndh+hyQ1BfqPtspnjbRaXHZH
hHl13WbeCzoMhwfYbqJ2ninHvp1quS1idaxljfy29jLDbnkZ9rXkHHagQuQGJXz3
MmEmh76eqSoxhH3XaVaXvg==
`protect END_PROTECTED
