`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KsTFT4N0jDqPvqQO64INyW/1OMD44nNFxrCxODl8XibbLlJl1vHS7/8StPJ0357h
NOUIvth0wWA8vdFv4YUcENbjV2MO+ZH0NTYwcXERzARAJkDelJY8FaSgEU5fsvje
M39Wq3EzGFYAeiXoHTiBWb8wdy3AvIwSofPkrXRG+V6rXjeayoIXskHs1RMxtug6
JNLZcPn4TOfhm3gdUbaIJMYrI8wZczE63FoZERy9hofN+OrHFI+QzciZq4lJMn2D
B8uBUtLmXjdw5D4fXIu/Cbzix3drtSrlMRKMy/Xn2ppz03Bah8pkCvYRW9Q1sAcV
Qzkp7RMrnvkSNyXfSlsbPWgC9u4LHzyb4cCWiNuy01V7ReRKkTlZq2gvsVn/eJQA
Ke0M4lnrgt1kZZiBnJccksSXfsQL8oT2mgTDf6eBdG6XgsTkTM+Vu2ejIUFqXWKC
G/nLK839OkIWJC+i7txMvLkP0vrDJtIe94iZ7Ee95uvG2ydRur/sILqPVoEx7UDg
I/okkfTt8cVLxeBmqye3V30w51P4jB+hnF6cREqOM4WbmiN29x+lv/QBYl1b5pIo
cYcicxwnYVufzkFGmau07H/ij7JHcs0t4wxecuvBaoEKCSTEyAE1m84TidsNhtwq
f2sEAxiScmZNyk+GqmMXbSSWXrLDTY9Xlyd0+3gAZ9mTwpVojH0/xFdTbFe4PRj2
imXGEfvxCnlS2kW+hhWGE+44hmLCNSWzQrjzuSDj95674Rwxq4OJ9hXJGpVJB84Q
Ws44sdwRVge0IJFwu1gHncp4Md63oFh8Xb9ULH21zouFjYwTKczjfM1JhlfFChz+
Q4gYCRt8Mo+zAQYPFB52HJhYUoaKo4mnUI50C4N9REWWOLTfsK3zLYLLDdG6xow5
p4ZpMFvSo39aPeDz5+2OU3bbI4xEsz7Zo6AWxmYVuFosV0xjNhdQWbJnM5uBRcdB
IhdeY1gKl2wxChRzwTKu9pHo+uHowcREjFAsoXrn/Uo=
`protect END_PROTECTED
