`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WK890ponvoSgL7Zm9YRBg/kui9WYfsMNBu4XGfsMGSAmPbFokLccdDrmyPrL3gT4
HJWPYrWR98CtPO6z2ptOzTBtYTmkAImddWoSHlARiTdxpck/G8qTJuKS8bGw57oK
qiQjCWLilW8xKCFmf9EQNdmSYxp4dLHkl8N00TGRJZnWOp8rpMNEUZ/LSK4FiBiu
CTUEJnnvKsnIiBIkjCXEVW1S2LZGays54RTG3uAIL4iQMgARCbvHFCd13REfTyNe
M7ZuSUePr3s2sSQxu8wc5HUO8oZO0+RByjH8K2bgJGcu5D5Hh73DM0gAA3iMTZhY
7KX7yMfzzEGg4XKBIpd5RsA5bzb1Eibx4SRAFhipMLn3muDbD4nhdTw2sGlPVoj1
uuwHajhvMs3iJljz+rSrXxn2zAcj+ZQG1uHcJf1+SY1kif6mSsFVdtS2qOhowFKP
xkeqiK3OGuZEwg7YnCe8kE33kTNx5EZyUJI7KIJoY6pHR/ymahSF7J5cqf0L707J
lsE9qZNHRvIpjudV0r40NeZ5YIhVSDtSdmjoyLK85f4k617pv6W3G5l1Vdy8n/P/
DP+AqRS/V7kYPMIUatqM1bSPZHS7P/m1j0cxBuT/cT3x41HGlE4YUFoUPgt3udTu
pUUUCR4WSAu2nom9lOZnVFg7xN2Kkt52tt7DdewvByBJmrQKLPtRKRyz3zC5aPYn
SNWbfqfOSwxU18MrUlcR6iQvA/AofZLeyi4QsAX0p246ba0uiroI29LT/NLDfyby
st50xs5RmODa9EuJUAaahFPkDfufbAB1Clx0sNiaGKRrYSQlUxlMONTThyk0Ggsg
QDrOxJi6OYkqgtbKHpB8dSEHYz/W5weOrWnm0WgugUC5faCdM0hVi09CFgqzcZA1
7D8eqOK3pX3R2MyK+NlHnNPWh7Klq2lPYax/G50g7UspZHsKww459fgJvQ+SAVFS
QZT2Kiik9McorJ4oA7oNblEkXkyJCSGsrwTse2DZCmmxiorJY1vgPdc9UxMRsBAZ
1U+ysj8zzV1HKrJ9OnkqNc0A3exO/ngDqYAXjJCfue8tCGgPsr03c+J04V4cAJ5X
4kgy0I+lA/iQsPv/NiljRARFt0eLRuIQdbSIZ5ETnA4Z7WOlV6qJCgTuHn9b2vIP
H77Qqx8EAWpoPwuhI0zJ1qT+LFGZzvmTM7gMwS+Usj3Jd/Wo+BjhQsglPoSkVuZ5
MSbL96zzeH8pCxcQvJs+2FOE/pQq8w441ED/hkEVtPfDkGSadHzN+4CpWC4tQw4P
eWynv1f2iUA1yl40WEllilyR/u4OjcCc4Hd++WQ6rrKqdPxOiWZXUgmbMAwX0gJY
Qcj1NpYw4HyU+8wIGz+A7wAxUW7LaJ4TeyoITZtHM1YcebG+EhY5SHCNNqNOeVt5
wOdTYFAw2eAsjHYfADKA2xM7BOSMIWhAO5CLTVZYwnllT5L/yv/hPgSlmUKxN7vq
tfXAYNdxXsKOnELHM4OXIG1+GNvGIh+NE/eUH5AMTTEeA2wETgrXGrRLh+RPK9fL
LaYBA95Cf61yLB+46HQXOcGKryB65TcZ5bLjvLQdqjZfR1czCwfGUk7Lx3qtwx1f
ohWIoWcTCTQi+RjQdDbOrq/8os2iiNtRTwHH7TXzfH/1sOw4FZ8KrP0aUx52Q7XE
L4xFGcJhh6grRT1H91z0IGwrwJckLmDCQ45KpENSqmvq15eBacf6Ef2GNF4k7/GA
v52kZ06GjG5T7ZAHJgIoyL+p/dXMCeiIKtUu3WW3NYmzKTWG5DIe62ae8b4ENeFs
S+9vq1HsvCXq7eBJa2kFJfjkmmX8C6AXJlz/SuhseTDLouZGzqpKqd8C+qxtXlrb
IB+WUml5icmuNxekU/ETj0ftoQ8c4nJT3UzpST1kiSwOWZkc1L7oxVp0qfRhqyZt
V3I6kfGVLYo2ED6yVxbY5jodAmZ2/5N1YFjdrJkC3/OhLt/5S4EwH2zgXfJi4IJo
Pjctr8OVQyLAh/izg7LMVay2uFauUzFNh4D+3b4oLcC6UGNG+LJRFM38B2LriVVN
bi542JJxo6CH4RonYQu6BY6Goadvmr2scc3BVgPsgvoN6gYI7mdKHeqWByfeeoCP
FWlLCPUIMD8F+NREkO4W/EsXxt+DHazDjJaXdqJxC9z8W2bSEq1LcVnRQKLoetY8
3wkWZ/SyyMswO2u/qZi+xLCKbFVRHWtdaOO0PW6C6uNvwEAG12X5xIj+rh5CzAt0
DoB3YGESksnovX3qwtrE245Z6kL6XIy6k4Trlhkki+KkxUzXkTa9hhXDx6YMmxap
OeH2EE6bwrkWlwyEjH3f64QR3HCP9FvXPUjOop3csmyfZomz3YCU95VIE3b/DlS2
lYJhFQOdk5SSU24wzGwTwu/GAyUtWZiDJfiWefbTL9z2OS5YjDpVrZ/saVrW5zas
WHVajmgdxapia3wOWY7jRRqFpI7/Z12IY2okvJpvEqJHDtj/VXIkwMh1puImCo3x
lHGjJjdwjpbfPlqXHPHX1tjCYEjuNjqv/t2pDJMeQFoJX+JrmGHbjM/Tx8KbIZwo
EH89ukOY6kXE9WZvxOjI/hKHjmUQh75gLexRaHO32YxhLpWo6DyOOF0sDQzkS2qt
bPgupAWIV5lvckTIX3bNPCIY+Emy+WKe1Py3rQWunlLcmHa+EdKIFBN2XtxE7EJ/
vWbc5DJy4RnhJvzAkmULvspExrvNa8Lukj71cCbYQoX0EFk9fqQ4BB2yJ1Wo7a5b
oczWoy7YPuZQntSdN9oUM9Y7qxOFgLgVGf+KnxHv7GGmV8SI4Rs3cTKMWkrE9hM5
V0lnxKfFt/fltVoPOzZyhlFQGx1TSCtwg24Lhq+KJXlQSyyh9uBE8Ha3/1pNomBX
cKxdRitjPQLSLWSvcUjwO0Bco5ObJ6A7FLzoJMsenFU0d5eE/jW6dbCeAxzvvbhZ
iwRPANR2XN6qelEi+Gxf4XxMfPTK1WOiOhxMZjjNSG1UPBlYUEaHLJTNB5hb2f5M
/hd8bDsp+3jkLGFKAradm9MG6PRbDVlJRFW0Fc0c79gMj0njZX7uQowUO1KciUIM
v3M+pZfkAUB8n/9j/F/rvS2FphYRrvameBUs0tPADxB/R8EgHz1YumIvGuJXbJ+7
hE7aKGK+C7oS3zGJ4ziXATJGXXA6wI6ou2ADdJ5LUltbPl98Rxb18l2zDac/Ho/G
EC1D613MCq3Td/6t6SGsVrGGH7UXyo5PHOUBg5cRoE/tBYmyRyzk/p+YHW2yBppu
Uezoq5jxH4A1rG/++kpl6GG0+6XPk0jsZ0gUqAlYfQeWWya+s/aVXpjFw0WDlwmQ
UOTbIPirI+vu9SdTdTeR0258yq5EWEUuEo3rGybDv5V2GvkvPCJsxd5+/c8quByS
0pSoDtLNGOJZhgMCgpumHT4Y00Q6pzBjKqQ+u+bz4j309C8Pc9oP85iojVQ35j1T
lGT/jiMPvHU8XvOQivKrw9FEqkjyDdPmX3VcVBd/J/I5vN51qXIVTQ3bmUPYdM2m
zLDVuYHDc9c21ZULnC0PvZdR69afMWcitO6K7DTVjY1lOu4t4sCXm1M43QLiW4BS
w+mcBlgs5yWt5B51RNoOjY25E/9ReMH7WteOSBQt9FTwUPhkRRFtqmDfs3MoHTqG
H8OKN0v69TzMOuLiNIeYiH7egwpX1bw7Lpkkd6JwHhYASu33LKLffwnNPaXu+Ukr
eUfB1jOgGKKsIFWCtoPlrBgV7mQi4h0Uy2Q4sN+tBH1RVOb0zVURbym4kEFHDSMI
/DhUPARVeyKn7mgAGVro0fa9HxO9ffmSkiBIABg6oJLOepd30ySM4uOWhNMT/JmE
KMWrL9NaC/q3DlYkvLPRdA7LZYwWpntfuSkHZ0hEWMg1pFNVneM5BUBaAAjRkdUQ
3zsc7gsKKli1CjtuALMPK5ckKOBQIz8vygF+dFCIDvTvZQ1LKSyjfqDvqDPcVamg
1Cc1/AEAqcG+RcGLpksdJUNrJR4ITKb2naJHDEWROeguhShazqewnZBZN8pNmRP6
6BJ5fslxZBEarEUMdBqO0fgrBPur8NJATq9llMqLmC/AvWGfhFIxSq7grKOV6NCn
PWquVVy2BvJYNGYY6dh5kdrJjZT90GDk2063SDgPOnqMmaB1soPv9xPFkAz1DTPM
MLMBHh3sLku7lyRONXRzsm48Zf7JuHUWFGIlGFRoY43WdQ6rl92nOkh1Ja3i8mjl
G8uNMqiKaYBk0vp6ZTgCiXeNdfNXvHjYI8icNfk3moLvWihkTsm1vIoU6tBbLPr/
Tmb3EXLgcOlMpMywPT04zjiVIJNQHjDWlKOxhSIXh3txoDgwSb450lxaRnABozqE
JsbowOh0YRUvBtPgAYOR3IKsWH+9NY1wzvO/fEY9w2YTXCFs2hrf4SuYWDQabwu1
8o8xzw0w5QNTSl8rVTsdakFX7IF/Qi0/YNsLV0vv5ZMmSyRJSp4N2M3wIlsUOsCd
3k9qWGxaiQAr2c5Tp5dQV0xOzq+Ah4nV6Mujp4wKk5f4+UWwqqa1oQyxTcbm4BRw
s+f8dydFp+lrwO6+hlUXhgb7NHRqd+6ieX/yVJK8Hn1Xk+0s3H7fbPyfUTRI48cT
nnBWtjAuYwGp5kOaVk2duLi5kqP7E+MYPYem4qZnMFEp5JUtvkhL8DBgJuVMfolq
DgQ3WDsaSkaF83tLUtx2W/MyYzZThVCzV5dbWJf7SvcBZ4c7z7wVLCuic0bAqi23
dUPP3Nfv4mHjNxPx/tG3LjmfDTBWuzwn/2PEHoG7aGnpIFS1xWPyl2g2XNRNhGWu
4xsVDkzm1HJpVnhtd5rKpts8OvAB/sgEF8TLfX1YI4Lf2JyOu/Q3g6xvTsD+kE1y
GnoXKq5r3Xxit78Iw47o9nxtMTLzFjmH4sP12ouKbjTQCI/CJtayBFlRSsrbe26K
CozZEVPUgRDDTJlU0LFKjOPzaEMK2LPHF4oK9Jvvz8KxYXEtFhTZTYlx2GSp7P8s
chhnaywYo/tZANHuuBsTy5sOZnDP6KvHcOn4jrmgtYzeDwbovyXYcLCBF4gBMfpT
Azhemxkx2OBZwd/eIj2PISwdDeVEFB5do77aH9SYHaFNKe8XAuu6vFd0mbNh+brq
A/rNdN9BnSl6gC9p3mQ46J1FazNq/m7WSI5AZ6UmohN3BZyEs9zPXo7JQs3EEZ/Z
fpWvwn1hsYi6LRpOsgV7LifHOgkeLDFpSNA/eWuu8TGHEdColWOPmikOG6fRN4zb
lGNswdCZLvd3b7XMf6uaObzP2tF+QwfTk2mGNGIim1g5pm5l4NeyiphBMSB+j/Wd
5fYsaqWkcmYmCc03UZY32qct7aS4J/Z2+acnH6ApDa2cTCC5UTpCQ/Kpf2EXPuwD
zGKXyoXbhWsCciCRdqIZxDss7rewxP9eA3uKb/Q2stj7ravcdvW3avjrxL2JXNCR
qhdR7VbSl+ZgrgA4MiDE8RNg+4sybBGJ5ZUtNmSWlpkrqZPHRtw+yFD/QXvS7TgJ
Hihfr+j3A1Fdnn2cDWhtLcS+fMbSf7hMmiWsRC0bBxRnq8p4a0j60kPRqfxc3xDx
uh7oarLgJl+LpFf4H2px0QbyCKSM9YGENDQUd2AW590YH5IOKnml/qmLX5/LX0W1
X9sR9V+fGoyaJsRpdLpRYRx0pkeS7SNZoSOhHq9g1hem5Aww2Psq7pxIuuA/MX9T
WBg5t4HMk7RJdtEUr2jsBAT5yZC1j5WNExOVZ780o99H8YXg/Wc1k3HW/XDvQ8Fs
8rgee1YGSocjLoWF+Iu6EeqPYCpaAecZIOq5VJkCMw8Rv4jtNdiP3fsQN74MRT7x
IWsrcamz+hz80A3huVA/DCQFmi/kYjE0scU0EcRi4Z+dRbOc8uHDuIhlr0UjxZxv
8rhvcFoZear+oQckc68ziSoBBS34xsv/LlZ6OUiZgMVWZGo1cyp6Qe1jzBr/VK+L
N/OUpvfl8BLQz2qeH1HF+LeqXeXdBKOWf8LxukwGjsiyLDXzYsLjk/Uheo3VWHDF
wFTO+B3NeYBb+DXcVJN1aJOAuQVZvR1oSStTqoTrrxRa+GKtwmC4aDW0GxPGSP33
nW3DiOnPSBGxM8oOSKVnwNCmDZfXh7ZXz3DWITsuWpciU52agQtXb29rlcZW+kUW
soxa5KAZ8WXMBYIH5Jr3Uj7mbindx2VLoUsnjlchvBreSCnnXPFwkxzyXMVYazeO
wX5l/U2cA0K5Q8sNEstVHtQSwouCV/DgofMsc8JPR5xcvITA6nD9O0UIysJb2paa
IWgw5HL7Rwy9pZIWz4BM/Wrdu9OPDao8HmgG4N2pL5LkpItZtCkeh27XFltsFPHy
/neaCh6dtR1VZ79jyMG5IzQGHVnCi6RlnysPIJGLqdD+GFiz6V0Eo6S60KlJFN1g
1xejP1YmhUiNjf5bFao3ww/hJPu2Phv8ORMa3v+/AH4lERMRpknAg41eClxtEDHn
87QYDbbpNvUHpjsAHKlwCva2qTgjQ0R+rXhMBlkUxqp+MTmfwm9RFQKZG38zgv8U
wYZf8gHf2tufzaXNionhdGjBpiiHAcR66okPwG/CG3Q=
`protect END_PROTECTED
