`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWTpCFF/JK1DF+xeTSXatTNXAHihzBJU87eex3NO3GuIO85bkIN79kmuNTISfbax
3XDjgtUFQSD0ZdII+acOlbnWzJaWWGC0Eh/dD0wVWXqW9xOV7r/wBlmbjdbvZwBO
qofk9Jo07c+KHtWHBYV54GzQul/uK2IGrefZVylraC9v8NjwhhtwduWnut1VR8nS
c//dagA0YLeifgj6RCB4Vpi4Ie7A9+NEqRKMQUqdHmDSDwyJmcOK8e7LIrfUisF+
xPVbAShuC6dJ8gjfhkl4lYYxBfu2DDMVMiubv7kCewpD5mvtAO4UsZHS/KGsNocp
Uk6PBDA360lfv9YtTP0d7V6SknYvJVf1WQuovEi2o1OuQoeTSxQiLnG5JlvlPhdT
jZdwXXJ4UIHn83tr75UC1K/wZwX6GSWt3jkm3V7ig7foreAVtXH/G36ahZWiuewA
EjueG7F9/yEb5LWlFEHXoqhFLGNfboVp/QX0dQpKDUmhovjBSvO9ev9UQk4RmDwf
5U5eKB/gKDtPn3c92t+FDVU5/LIjA0hLw12j1bewmCnrg098KrSwDbND/mTZh06A
lx+Q8PBDTPckeBcF/3LRJFLmTCq17rlvY1jym4g1erxW4uImXklROhlwW6c1ZuYw
icv3VVLC5YTwhuSgFQUcUWZmWmCOKH09osg3H/rOtlpo1n8wXD+EUxxn5Gb+dFld
mSJTsybMwbpM0isKajWCqQ==
`protect END_PROTECTED
