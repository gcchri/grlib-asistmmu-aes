`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xS/XDK8X7UoxAZ756cQB+9XncDGJFqYYXkyd1iU6cQ9H5qGcxlS3Td3Zmd+iSGEl
0G4x2IP/PdLP7qutjiyV+hsykKOUEGVgB/A9N8rr2lnJGy8G1p5F/+pPnKu3kvAs
mB8FZidjkdTNVWHciCDTfgbA41qqJk/8ryGCd7JmYgxqB3JIxT+CLqkHSgdaArlY
X4MOlSU3O2EZ60th7ghXw2dp8cQ3Emfb4XaI+HVJ3QlLgTwHhffj4mSpekqilcv0
cDkAyvtS30wO4qWSpObEiJXSPkBGU36KxldcCsHkWnwK0apoq7wMRCH1qCLzug/Z
nTtFbquFYIioxZv1W6yUTPPtenQ9GC2Fc+kGiUIjBrFFRrpblusXZhWC4WHlWwqe
`protect END_PROTECTED
