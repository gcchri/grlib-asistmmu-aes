`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IFyUjvdTx1yEHSe6D9GfmqqSR8MKJsR4f4xC6i4gmhVdXLhMIWbq/AcuJF8LaBYr
QTxblpehmH59XwGWuZDv7M9EbmAi25CpI658T6sYdxz8GeXP/BxnUXfCdUAxZFzH
1K57G/lqPrrGPG/qn2wkkWBONjF1CYr3ZKRrHD23E6skZ+Gq5iIVaFECzxv6kilb
aOLNxmCDKNCaDKicIuenPgInG/PuMVdjz/4Db5dXqdI4UyaZaH5bqyIbqRlMiUPZ
xX5Snnd8gGSrZdbY05G4Yf9BgE3pNkSh+FmXZY0mjuwfM2gcdweElaIR5YwBuLQK
UgSLqyjsjkY1rON8iz3me2sdYz++IwPleU+xTfxkSFnDBA+niJ61Vh72wznmEFgy
2CxXFocIYR+Zb3crRT6prdMAe99ZVQ1cWDDHVm2dEOTXA+82dV9iW4hKXukQjZYL
`protect END_PROTECTED
