`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5cTydziN0/Rlc1z+6gvEXO8BktznZsoKkeOFCEVZW8jlwJDGv5SVhz6mGJ+xBjNY
gjTbSqRsnqimU7Sl7D0XKJSQ2PSY2hVq44nN58VII3FwkTTp+Y649L03Mtqqw9WH
HuKiDEOGbXZnLZT0j0QEe5E66TX1eh+mTJYA3l3VaYHe9E7JUpBn+vBNCXe4uOd4
v3yKySUIPA1QvQUREk+4zMDLOQwc86xHm4iR0IhXmLysK4mXXewGLkEkd7SZkBEP
NS5BksMDqzZskIY834Hm5fEUVDMpc7ynd/cKyMDPTYW+oyMmzMSzqQhpVpN+xFpl
SSquuGEusgG6Uwc5RwAVdEea6lM3PqpQ7YWw3EkSD5K/KnK8M1RR60ojgDhPTSIE
AIqlAh5yhOzoGDRCPUia93Dpre6+Vzwk9EZ7C35ywuCDaGHQLjARGMR1Qo2PtC+u
U+8IAlgJTSY6zHuhUao/mrnZfkAyGdzKJ3L5XULrxrMsOuB5O5e4XDHmrG6Z2nVb
J3LwDi9awC5VGI/v1coQ4VGBWSQHwGNBPVlKbfx0TUm8WpyxE7LjnpZv6dabMjit
RZoX7atPZipBWFyPcUbpgysik9DS0tOhqSujmYzfMZNW/Fbt20IYicMbqxjsANhV
8vxoFhWoX6dFTej/0CSYDLsU7TdIQhCCHPW3iigVjEAdYQ6VgKX+bPJHOucMtmot
ddcBRtTNj7borJ+WQYYnZq8I2pxWrdRMzPYGjVVG1Kz2f3Efwl6C6BD7/Uq6QH7e
g/npjCPlIAPZb4p811PtBhokuYKhmfD9ENQYGXISn6f33PLyuPVFpKRZhNEqWEL8
MO04g6WpkiM6daOcg8x6ZUfJQKrmSX9nVYl8+amO0y+PkqIELn181onvXK5Phws0
2V46veKxCPH24/eJgf4kewcFqUY8th6I8mn+vAVWgbRl0DBFuIyWFa2VAG8vrhrt
znvIBH94g9MRDS6Fg7HrAYcVBXOXhcHx9Otz11ewjtJAIRbMAi1jlDMS/Zoy1YP7
McDLkV3LHPQoxAffH3nUOS52r82VAckB0FWEYq9xyoj+AEpwl8NUMDZ0XOxcURov
TXs0zmueBGMqsYaR6YxgIX498ut04JCxWF2JPwEpvQdDE2Zl4AkyVyxNjD00d6oD
sdxGKDbGizYLcxxlZ8d8zwHr1IXgv3/B/vFOVuve8cNUklDKe1WlQwkKhh5LgEzr
rQ3Kz4e14anfqsblB+CPwKvZojccAWfIq56Tb7g3jqNFIyDNTS5kgNOUTH7Cbp6W
zjcsvx2qTmIr02y+iEQgCMTcUYdn8Prnv4iHMyE4CFtVmrVy/gsmCczUyczXTWZZ
LK8Dyk2lizLkrymVoVyiOHThuScLBnXes1Gi+8KHSK4oWmCa31MnaXZYZ4Ef7WvN
tqzYY9zdwocxiPqwWqrPyxmMXfW0d8YLXVu1wyd4XQcNv9mutE7WvoEvBwuNhU6I
qCRm0wbN7hY5Gu1qAE1D/gaR8vMGBYZ18HlxfPPYddOHjTu5QnQyb+OhumdtP+Sz
4D4cn0rnQNG1G/XUa70rEMcOzhQBVpCzxsqbPk/ff6Cwch2tuISvq4YTLpuytqvS
VSh78xMvL/M0UdxbkrFl9x7MP0+QOFNqC47vwCGQxxmxNgZnkDDX3ejy5LnmSPHS
ctwV69e7+MUyGZIuqDUf7aULbchDfV+YyM0x99ngfQfyXPEwuC6jc7SJ5RmENJzH
klYMVo5Mm+AzjgKpTgF5lvGbVyIRYN9uRaCeF7gR0JiF5UlSOMCDAFyd6kwbfk26
Qmu/b9QlAeAj9d10tg5mauDJjIflfIOjSxMnKdZq4u4wdFuuWBDJPQ7YzTdw+OFs
l3LRqJwgXYGY/moihYv60aHmTWiLVaktNd1gFopNWtl5wXiF52YlUdhxu4QFnmdy
tH6de0bPFgYd/mb2xXZAEsUEoNyWl/9pHySqny9fvmcA5CtqpNlpIomUgJ9JNgPS
plrnw2bIEvLyuIOTBk13EZj5MHtb+/JnMvRH7nESGZj17Vto65zeR6fLoQcw8DdG
iRVJv7uMGrEjoxqVGN33/tmqFbEsKzEykLpbf0Gpewp1VzHri3BP6Lobr4tawHaQ
FuF+GOrl5hv+15sUPIxvoW2vx0pHj9ExVCF98lzeN932x32RpRLI9m7lEk5/HpBX
MaBXBegPuY4/VBJXUe//6IBSSACJKzD/HYBrvPwvp5/P4aO6+Lk1KJzmxJbVFTUe
C/EyyVQpdLvaV9ETlwhK4E+rrNumcHGX2UEtTbAsxrJavSRSEVM3511e62B9gwMO
ho4FN/mB1t873uem+HS+/3cR0yOZU1HCyUUKu0FgDUX5Pdlip4ovQPFlvR415iwB
APZwOzL51dspQp0bzyz8aETgb4CcuBkId1XIe/XN+q1NC1ZaZitFyqUY7IysEzvb
SxWf2fnIpUwAYguxx/UiKCCBe6B3aYEHhOhGoCO8mcBWCHsdeLoK5KFOHz86aCVf
nDOBgcV4hRopI2Yc3r1Tfq/ir8RA84xGezl8kCANSn6sGhRKS1AZDyCnwa1Aaeqf
7v5NptdfNfmTyfABVKX3+b8egGOVmoDHyYT/XXUicV8YBcXrC8xkb/AT2qOVWfzO
8rhDKj6snT/RAxueibT7Uhx25zlOaDVnavQl1wa7nBbThl7tuQ1Y65ghPm6ia3cw
FwFrw+Y75povNoJ4GTGljWqhWtUkHBYucAdFADP7ziHMzKMqHH29CWNZzPqMSqLb
mhBoncZeD1qjZ0P8wFj9+rqzmfAGkKMQFp5t5ou2Ce9dBvKaOdBVkNTiRylq2tqZ
RpDRoNT1fttvrALfwSqd2acBLCIsV1Qas8KOo6IYLIIPMacfmGxD/QgzUezqN/C+
n3xSpYVvfrF0iDHWFnZEW9FDT7Bh6aTEfbKA1r8bbNWM64ZRElAszlQso6NcBhOk
vVBVGgKaQD/bTwyWdR7lOlNa5MZIO8pBtq73ZPnFRP3xPk9PdT0zqxMQO0fCj42l
j2Ka85k+/ccEnbzMhpigONF6uwxilIBPhGNqDXe1U78=
`protect END_PROTECTED
