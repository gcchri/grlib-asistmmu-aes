`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcEU4vvEhp5PTW+KpENSF8TRg7rYc69i+DV4XnrUDG/+hcmm1F0abKCrxX7b9bC9
RdPKe40UWbKv009+P/gAfPn2dSC0qKy2G1iF/BWubK0J2Gd/QZgUD563M8jeFWhH
z72VY0uHvM538QJeX7A1v/72drBOMEYZpFK/Pj+xvsUabEBkjKC2IDXbwg8MYWZl
GyN1gZfuZuXzbM2lzIW7xJX6v+hYfw4xHsqrYT8RWehwS0cArntFE/mFx1lJ+IH2
lEWXSjs1CPFb1+t9VW63R5TuFdlqWyUHaqxPqtk6Bqt86MYgtx/IYsz9LWqxE4Jf
s5ebaijTRD9K/yr2ALe30fbqTX6lsmN5GW524wusXu4w87YVpmG+AQf+tYFEorUs
CGWwtfEf3E/BYkhpKmmx9UOX2u202tPgTKqMFFz9gg3vCueVMJtKOxBCJw0LGp2C
7QHp8U4B1ItIxanx/HF+/y23DzIyJm6dAib2hsSSiLwv29bcosYx5JGvywhIDPbo
6bbp85m3fBexZ62UJ7L7DRDpbENiIo5lF130mm/mB6h2RzYzKh6JSL4b88gEHs48
bQ03xgUDJ8P10dz22lCQPCe9Ho47dv0VMZ+Ke7qnpng=
`protect END_PROTECTED
