`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGau//GlfKHIwU6c2LgqGSq6PG9qm9aerK4FwRhlW/InqFk4bzWk6DI/bgvpYZHc
jewULIzc2wnU975mum9mvVtw7ZFz10bmVJozXSdZUdgEfq6qOgLx+PmhhKfuwxAR
S9mNQl/x6rkEzAlR0zrWmJeNfYPbYZH76ebFPIy+HIzIP2cGjxlU8wabWBvr+3zs
q/f6rMW2nkG71LxQ2qZdpVoHJCKwC0I29ACeWF//Yv2eERyfPohy6lHiCLBFF2oW
RYgk9fvIEd0a7cpk1+rwgZqDEw3mjeqOnnvVwbYls6z0sq6jZQxp2qwRwrj2BHH2
M2IgkKAs6EpGoMX6ukslkKw0WdJC6s3jZyqbwYnUJFBx/SzdW4C701ndJrUiE1+G
XugxhpLN6CyT5r0nOKXxuOm5oAej5MqGH4oBT4CMSf0=
`protect END_PROTECTED
