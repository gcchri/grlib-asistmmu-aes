`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eTH6K1bqgY/n3C59AG4BTwqsvFz7/vcQZrv95wCSHQlz89xqbavQdT1Tg0UAkNvh
jzCieyPOtcf8GOtR+uck9gC/D0u4wfPgr6/d/F59qiSqOMTw6OL01UaJs62Ps2cy
Ta538QKVRNMnlwT5Bx4kVt4BMTF932ZD03HWfvT6qWyeyImmY2C/2ZUJXFiL0p1p
KJhszBzU23lm5tPfO8vRc4svvXZTv7H8jxCndXcmTbL5zTEQ++79WCqE8HORGwTZ
qHJbJOgd5FU9KWcucwY/sy9YzedLMdXtGsFDSWoxNNy6A2WlIAdGj6bVXabxNg9j
ruHSvUfRH8K6HM7HAtV1rbRA4Yul12SerpTTH7Vrzm9jcEToHALwqdKPBxo8mZ7t
8LPKQUDb0ew/vzgCvmF5rg==
`protect END_PROTECTED
