`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6GTpJadwtUh19b3tKfEOOPxFDnQdQi1UGS51c1IjqEX8YuXomFYvGyWdAdVcLch
p0qezJcjSqdzfPgS1W8Tj+rEyfY0cGyQ5diEnIsqnq5pLuT0U7xz8poHTqyh0aID
nJUXf923G9SKmw5Sg/1PCKxz7w6dA/N5Md+C7pX8gxbQO6Mk9/u0jNFTjzj0kvpA
dkkHCTBodVKl95yp64/JnhBTGko/OY2auu4erqTQyoJa3kfvtuJ7LbKFPna0Uff0
KjyjFnzGw9cnc1Tp0g9psyUh2WolNSES83g2G2C99SLPxHgf+CAyByw/6gD8wvYO
E7Ud+Avh1c3TeycCcKLmP/D7LOk6a7RjjD0sBlsgf2c6noqqJ5tQcJTcx7SyJSAL
YEIndbGSxTN6jRzkWgpGgVZQJuAvx8sTpPC6efwXcuvdnIIngrAIJ62nls8AYUEs
`protect END_PROTECTED
