`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YX/I3fsdQYAUeLlTX3Upq4oPthuoLeYy+Yoqrz3eG/+KAJ0buxp/hhrUpY+t0lLn
Q04b8VKx68OzWkkNksFWRb2c9ifIi9Bvg+pTVVQwVAvQN7abWXS5Sq0pJekqWTSw
J2BOE3TnPe/3K8O++Hkq/EbbCFtb6bM0yVn3sfNlXLm+zD73tJCnW1Em53VfSeNo
bcolPo2fD7ZolJgd40sZS1VZNgpu7rvM3Gs4DDYLGkjRkdJFdKdjWzB+8dy+MgjV
k7LBfAZy7XUOaHxOiOCYEg==
`protect END_PROTECTED
