`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FuF8yaPrV1kcdrUaygFja8CNZpVlkMrar3/xgdiuL0hdNIDyVA47WOBcgjDKPkvx
GU6KG03kcP7C8PejFGdMuYMc0atN4PY+Th0ekbWCOZtoa16NqaDF8jacGqXpwHbf
6MYVylO3TV7wJCj9mikHKfKiR0ZUzrrS2E3EMBVBvoEu/ScdSghJLnt6WrSd1StS
zOhpskWj6VvIOY8ik2NHhyxixIVFTLWngYQtsCAeo31U1VBKQXmt7YogarEYJ9V2
0KrCAtZZ8WHpVV8ltL83OkxqElRwsXDvqK3YkZZxkmBxH+1H5j/A2jMBqgos494Q
7UOVk/9l2UTXdaGMGOzmabY2/UPvLAl1NTKlbSpskxTqR+ck0SbG7q8Weyru8XSR
ldXXqTMeHUtpsS7ZzmG+tRR+eNTIY87Pw217mplTv1NpeZlU005gNoebytKlZFnh
cni6IrGqca1/IkFUDkZj5ox6g2MGQydGxNvSAkDK051RGPVwXwoGudwnRZPu8kfi
A0b/WYPoW0hwsMhFJZbjNLsr95D1x9hezQKVChm2VCo=
`protect END_PROTECTED
