`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPQPRCAHRwc2xa2coWEO4UiETMmb6hWQgDwLG+PKPG0vxB/0UsOf2C1CRjlT9GYJ
epBhb1tK2jxBCXtHLpHEcAf7JJc3NKIQdeZi6O3QWSeSaRgibtc2f87vGxyx87vo
32V8ykeKj3Djf8UjmdJp7Uwa7v2tpp7A/MsIIJO6Doelxg8YliZtdPvGBMsXaC0i
kx+xXPP+YJcPrb59SeXZuIj02b0+b5K/nvml0USQMLxGCpKSyNOgDmHGZ/sarm5k
GPXw8yUk3lbVVNLBFOaxpbAsWTOgCukgd94BR2AYT7N+eGfxYa0MK1yIOUrvB2lb
fMNO85Hi/wrlghDnQUmNv803ZW5jkrB77YA1UnGOqysFf8h+uYU2XJ6YYAn4TCYv
nBc2XH8SD4cftdnyboWAt6O0WMHuM2yqT5hYEiHUoKysKrShjslCx/Hb+6gah0oM
RaxfHiNU959qYBAs75XPm7ft+8j/Zz4SDFBoNjqW0mUiLs5w1a8gYFrBYb72ACVM
H04Ejnz5qdzZ/vSKokRvTkg4H0IVPLFvamI5AHFdoMmoyp8vxUcivonKgEO2qOSy
HMPU9z4Q1T16g5jnGV5nToS4f0nUWidiNkvMYBBRszUajpP/rS6WOmaYZ4GVCRfo
DyM9yK54yKVUYgk39ABE+c8Xyz30JQ61cC0AdePHG88=
`protect END_PROTECTED
