`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+SAJWn3RQKqu0pw18oTHW6Ald53cfbiljVOD/JRzkxf05uWBFJ0GFJg1TIOOdMD
ZF2boJOzbHTX5fADljpItxtQqU6XKlK4NzUPJmUsco8NwCJJqUptvor0hiFsFAN2
kcnkokO647etj/oWxXVAQ4hlx6vYy6dkXaFCBUyHW9539WSo6p8NQPNILVam5stl
R9k6U3VZAld0B99p5ZQTyJLg8G1JDcX2NFqGTntRJQkumXk5zEmhd6984SexL1a0
INBV+ITV/MrqoOgdaHtVHp7fHR4pRTkhRiNL3itpT0HWZXByiKO2pRWHfbP3u+Zk
ndfU9v+gLtS6nyJMLDiwevRanyCnZ5nFPCDpGIOIa1qHCXneMvriA6jzub6+A7rC
KRxp44zrc2NZGxXfTSRGICWIVzzECQbR4ZIqX+W9Nne1aYA1MaBgM6/QiYHK6DCi
`protect END_PROTECTED
