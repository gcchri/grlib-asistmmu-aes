`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZcyfMM7VwcDI9jPaepM0auZbMUtjbloL4mYVrovvKWn4D5ObIAKI4PyUN+cR+eu
EZ16wEabMTNMJyNFwLJn25bVtltEIsAJgypNJ//WRNPpV1LsAHDiHA2GcayWs08k
zPPl0RJIsvhve6UZqsZTom+PVXALf3bGbVuz+jDSbYSRCrwTBoS19iGkaMwOq4gO
b5VbkEEezReZwOx9uq5qrjyFC5bJpFvVvM2uKBt65XEoABM35BN11xpKieuEWAEL
ViwoW9omC3aZVd54QBGx+BbgnqpSRYIDW5sC5yuFuN4bqoIeEWeZ28R2/xOCWDUR
SA1Tqf6FaENakHozsOQs69eGdhL+F+f1IccdYlK+O223N50p2tPQdpjnzFPkPLpG
Q5sw4Jk6upmwqGUj7eCmxQ==
`protect END_PROTECTED
