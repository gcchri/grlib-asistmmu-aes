`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UsSj50N6nptjPuGSPqvByZsmVWluQhVy9QmFa9BQfVektnBFadI3DhcbKZ664zdz
BBgRhRXObRfKet71pJXIwoiETPrV8mSZiui0l3oZjrhxcFDoVNBU6BM621QyriwV
BQroLuVP6gK4k+U6f4RE+cXyws+DRGrXKroYly6CG4qqge3r/RyzIsL+fTdjqByJ
gDLDmgmzNpS6iq9VtOdbSI7NqeXHzOzUnN7ypgdstlsxFyi90jPvtlaDcX29eQ3M
VW54j1LpjtEgf3LzYFMrGBDpNpgMBkrbX9k5zaGmMKIWxGKXiCWvs/Iq7r3xN2aA
eiW7jglp/aB5vECw6zR8OHKkDyIOO5KFelW3Y/y4gHU+z2qhP+8uFGs8ljUMrfpz
+CMv/rqrDgDkIEnqY6ZXkeKgM7UmGZNKrhW9o+TRBGdSQ6JQiZi7K1kv+MmQFKlf
ZQQH9Z8ySo53WabjC3CBChi1zYWxk2g7Lk13ALze8ByWqBc0EnRsFW96/XW1Vid7
oyiXUJ6deBsh3JNP9e/RI47oum4xsgvdFVHrkb+QhIjixgBUIP7WQEvdxMaDkRJ+
tK1+8I5RX6JjsZVQ3sPknwuQRqbC/H6KdRtoi8FnlhnvXO4xvraGgJclgfWLhqsp
d6L/l3ZOhR6NYNxUCWdnWukufT1/8UTbBIOhU6eKsfHiBwIr+JoswqwlWApZPLgn
lmRA4xXgQ5/3dXHX68acy/mJRbrWYv3Mt53L1dk0fr+a+9ie3MZI4G0zRew9fbbL
iSH9I86fWWwoFu5TSh1XXT3AUj1eEv0BoX5oJGq59vP2FTt3HfiORvmTUZpRkEJa
YtmdvGUuSYVfHN2txABS/5q/f+K9EwOH84GlhooAHTHOQ1XZx8hzp5fLXMsfl2Zk
UuHqs1g2il4hw7o2PP7y7SaZy+q9OnxSn7A8q0T1CFBTEbAWobGe1+xYghP5D7Iz
wh8HrL7cfjq5iaBclRPLowVGkW1yKR/zEYqZUJiU8K0HeGmxixY5K8gr02KibGOm
XT9byy8OhvYCS/rBAGQC4fvCakVJalPKDmaxki2AsNNVtDn0Te+VgU/v562e0698
6nA98NX3Vpel329Q+SqlyOG9UlQDC8FDG6YfqETBbvqGv17m9IhEXCSpcOn+vkuA
+o2xXjD/9V6ZtposjCdYgX/4CFXwHAlEM9K6+B00VEUXI8FMIkUPiR5+z0Jx/rQk
ijs4nxcQzdchS/krPnvlWAWyvIMJpjRilCj+7tF50Ubngjmpcfcf149FqyKdoleO
3njfhEk1WYtTBO0NU3KCDOmYMgTxUrtAHU2DcEEHz4J0eIVs09NC7i6/cFAg6klE
iz6n6IJTrWvGUu7BPfAl7dPAwv+vDsK+uaZN0WHWfnoTj++lKX2cMi9MwFiPKLD/
0wj0vC1ILLCNAdLdKlbBzy+6jcl3auGZp4Onim+vO5LMkFIkpRmkW0pBDd7RzHci
IdjSZK48759jvCo1rXBm3ktnidb8P8kyeq5AphcQTkYpz/IIIu3B8HVJgj05kacK
+l60u+wjjzFsg/nrD8JnAyVOJmPvblZSpAcWAksLpgxaP135+u37PBmCwiyTJcIF
/6RScWoqF3as9M8TB42dd78aTmW/xejNp4hwVmS8pbWNNF9cOuAD7aYR/DpefBj9
9Lg0OQldFiJmMLkYFCGRgMxX8CakLLD9LLKUYBmPzMPOAFIgPjlcZhl9hb03fg3y
VIBF79w9iY4ZnUYE56vDlPTTrMEHv8qvmtu8kOxOCf5tIoSOpntBDdzdSHTEs5f/
YMO6thqJ2A3ck4C5ohDyvTIyN5BeIr49yoxLlT3mhTVDqCtg1dPQbiQJMnWhO+yh
XhzEQbhkXVlIMQFPut+FI4//qknKZp3i7umnoKy4WmiNDy/xH5JchLHAscNQKjMN
JakJGwpDwkvyMsCZ2Yssi9v+BC57NkKUg48iGFlTNNxk3aHbBwECYA41dQz9QpJJ
v8zcjz4X0l9lIrUjt8GlHpzQzopIZcsUYV8mWMASJLpcQphhPNXAYdtROrRWwze8
3nYqEVjueJ4wJ/9p4M7adaWMenRHSlwcrSedxuowN1sRmh2JihoPDyvzMWJ4//0K
9MXzw+Udpa10s9K5w/YOVRt7wkQGbeelcF6a4NrEd2aI5zhqiH1ZvUFz1/bfW+eI
pBJP/iGxVd8LH+YK4sYbwmAaBpWoRA/vPpqZ3Q8Q8EkExWW+n1A2qUe03s9Xs5MO
FgDjhGAdu1r+Yr63KSZA+CLtYqR3j3P7iJVLS5ClqCy0SmVk/lVWLjLEp8alpLWN
wRrFpCRhTE5vo8dr5QBRQQtP0Y7xxBF3EM4qTL7WIawhU//QmstNRYIRJ6+O9uLD
GW4qQUn7TPZxWlmRGTZB5r9IKC3pYmOxxLYSDA9vzQBRFSnC6zGH8LhsXaJAvLU7
S1wIZ4IoTBtTtE9WfWqegm0YaZnWymiEZ5zvy/P8laRguxkBtPzVCUcZKaWypRVL
j2Apyp6EE+w+N+EvNBazfRFRaEkcPcKc8z/7FnTJpbV5QeyML+VyO9jXq3KSOG25
mNJSZoq7FdMXk6SXU+n71oKxuzPebF9gVaxR1IEGI9BLCQ9CWcICtEIVic6luTR2
UD6AOQxouiUzoEd4Yh1nFboGH8HfPUhYwoNlW2kIMMhOcSdQ2pyI+V20fPkWcxSa
WZ2T0g+0U5EM1X5ms1svV1eISjuylVIMxCvObfaPIgvFGEpi9gXCbGP8od7LYTm+
UkNdpYip/B6O6FX6Gg52OQ4XeZHvByxLsojcPni7ag2hdVxsqZEswm702mfs0zsS
dtzLopU5cVggghLunG5Q4v5W/ib+w3qK5sKyoMr+jQ/w10wT1HkIB4Po71WIhKPt
2tXjqYJ/S8eKcbw7Qq3ReFBDcG1HoCFNjv4aPSHxUFLZZ8KivNjx00qybInVEb/P
2fX3JSEWIk4r3JzbqwpWULJuCgnCIIw+OWkV1Z4+cmGTlB/MkoyFu6ijyltbv2n9
Sj1Lt/yWS9f3z56rDY5ocY2KH31T3Nooq8toEVekgCU+H/WsO0jaeBYRLted5exj
/u3pAYk278/rz3bQFnKCFprytBb66t5RjBq+eOkzrh2KaT12WMozau7Md5KeCuTf
PSW7o25D5YXXwbMgz2f/nMKYTXXx+rFCIf0A1j1nkaFmdeX/TsfhQzAypYuTqUN0
h4QtWDT1A0igjG+459XuspkTANegYnhn+zPt5KQ4QTkm4sjd4+/ujPKKMWzx9GpT
GM2Zb6k91zLLAQESMm9A1nD/WirZtMjoSQSGoNbmnpOPS99A8iiLF5KIPwoMQKgw
o606AgpiKnMSvx25emXxUQmOmD2dlaaDAy5YvhoEKMfM38KjtCm67bNFZrrbJ9tp
2CL3QRCbxBxBOIU35xXXlVdcWK8ZnNtQe2Dina4B1X3g5CSPNDsoGJtNrlKAtL/V
mIkjnYCluJNt9lsIOk/UsZizVpKyWjTWlEVjbOroxNjcrxqZXEE4xBsQej7OlxIg
rLCcaE1SCdZwYKj4NZSW7Gerz7DcUNwdEZPv0Mz5VdtjjAyMpAQOzU48mncSwlSa
LQELkf8Weo6+aruuQwISpnohgakZvzEq4SWS5vc2LEn7nMrzSyfEQ/zeFb2PEDfc
V7BN312JRC0V+VVklDZInVrOYIJ5C2I0nhsgn2m8HLD1taStQNNo/ERJqgydhXpz
9uVC39JYKXRNFD4mtU13OQMfMBlufqaVt6RFyV79fbqcgoro9qSuO9y8e2Lr+AWv
4k5x2c46MjLEUNDALUKZiTCA7uUGQLqgHf0YZhZ1iCWv/XS2xCVTakh1381koLnA
`protect END_PROTECTED
