`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OOsDW6/xG6j8nrcoxJ+wzcUjo2aOdRs7ZN+bsT2tg+/KnLOHCxtT7F9Tqv/Nx1cS
tBHbqAO8ZIMHd1qa4Wm+3BhNiLQK6SeU4CP6xEctLAa6MycODJ9cRcHeDlMNhaT8
c1zXn/glvfigehuR8uhwwYcFAY5U3gTDlUXI6RAGAimlN7UGcpe0gLW3SB4aJGBJ
aDSxSt6Pqj+RuYA9E+9LBs8h1EY3K98bAD7t5FFwLIinBHHe9vCxYRyZEMrvK6BZ
tKangRhCVK1JT/RNs8D38y3O0azx2RbE1LAj78PxzPdfYmvwv9RL6fKjHEXNk/9z
Qf/gmwDRyd42cLPZzIC8QQXY4YKyKlSaCvmhX+Qf6c0KUqgxMQh554THYJ25pTbD
688vYMZ/RHU0BEvgXfAx3Yky9Rh3BbsypGcRFO5L28BhFnjvLPPlwmPm9KRArsyi
lidLf2W769N4cyIre/bYuEXI5NDXjnHjOOnpS9jLnpdQDJN5dszesNmDW2uCzW/u
L0Eb4iPtQa07H2ln74wDkO3PME97TLhPelBZlJgnl/PQXnCEDIxmH1hIA7zNo5JV
SUJM2qsVXivLtyxjdL0/l3m9vi8q5vt5VeCkhWYbl1Tv5GcDb4L8ZkPQ00Asf+7h
15PDVU1iUe8xRMTr6iB1pD92LWhLiMkqfR00GLoqVYpKXBMUnqPT1xoAfgq/hvVK
`protect END_PROTECTED
