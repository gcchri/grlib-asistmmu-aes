`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UQHea6PybMj4/1ccdjM21kcnwieR6ruftifrQAdtxmUmeQIrkg78Uxgcl9wDL1KN
bgXJxmsNfT6PltR7fCsEquabAtnLH6btI8DkW/8TJxI9DM/baIkCnbDAZZaT5o8a
VIG7WO7w95oU67jPRRjdpGLuAuYsVydVOGymL0lWwnr/O/ruzMHt5zymlIWbG6Ts
15e4bLpXDLmZkdOuViGGaUcpsd3+CtZdHM8BlrwRQC7ujcTsjiCBpeyXQRsoc8KR
NS6SA61vQdcCzN5TBr+xWxcTGRd3e47IDPALfBd2appDZ9H2LOuO80JlV92vHNhl
gDSTdqwrt+U+k+cTczoaPm7UUvnnGoFrBmt1yKgTRycvWCVb3LG9zRByhF7ZxgqI
3a29kTkN3oyy3no3oDqWz1of5R+nnRDANg8tZNa62XUck02J5q+eiOObmQLEmpG+
trMofXdi7VvZ+dWVhMcNApkTCRGDax27iJq9Z2WG+dVDkoMkXqD0hgLQq1AVyoiM
TV+NHfMV7UxJWjN4nMAQE31lBZhicSGQf5j/XNoBOXY=
`protect END_PROTECTED
