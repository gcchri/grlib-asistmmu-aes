`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNLBUsPHUgCA9AgjfQote0bblQxsoJlQGFS4WDufuthQzHAg5teFj0RABeX5EjX7
N1vhG0Z2Nj1GbmzfSkK8Zqd1nBuAF1leItSNLcQE7iHJJorw8KqMyOGF/qczyHS6
/cMi0Jp3H2ZWWf+Ug1mUmkxZMINxqGA3V/ADDYQuEntWLrQEANThe1jvzckYbSrE
zOAeEX/Wpp0hNW3NrUZsFLlEgjld7ZnsQTvSnjgG8EzdzPsu6ldTQKVxbbQoaq6E
l/LzlKXPOFlET01R6crLA2F1J2H98V24jK9jEYu6S7aY4cSes8PP8QglqeuzQCLa
UDxfkwEI8XffCXXQ6SYyXHLPGFu03bT5hUBTD0if9dZUdsX84ZSQ4BSMmmoHiTSh
1KA2kUMiRH2pYikC8sido2QxhTbAV8alfbX+3Zo+MuE/Ke5rKrGis3M0GUcIyX4A
unQ0KCwbhUxryT0QfhWM4xnWsEz8FWEwpBaidhx9HcQTbqYRuRFiT57RyzsVOp8J
MdYJ/4rHtr8OFmYMg//8fv+DrvU5ItBDs6YE2OBER1kZ4Uvq90zvrugpLtivE52W
XLIysUwW6oHnszMhl7tMNg/F41i8EbVLX8xmq/OYgcOJ7Na3iEfesTko+S7//f0c
InDaiI9Sv/Py5SBMEvDfC7AV5vx75OgGuedqM57LRGuc2XApwLmNr2GqLzRn6n9i
Qo32DuuUjyQSHqWgcYepnRkKzHZIQwincaiPi424wNdVobHgfGCrEjGMkna5ZLj8
DQt4oNcNUocNfOdQnCcUDMzT8mtD9w6UF71Cg6SdIQIMo0y+xDc5RMA4dEbbvlDJ
vmBgV03k0KhJ55YNIVElNkP57ADGEOuZD/jUqcIwaNGI1LlD+MT+4BzYZs5Q3/Sr
o54ekXfCPp9vnzZrxeRtKMygSBgWtMduLL8Kxss1RA3RcCfgWLPbuMueQgMmVCxP
3AZlWoasTUTlsNv8QRt/9faQ23PVFo1RCnx2FFgKSqRtaKYOjD1hSNxaWc+lAMvi
xBRyZIPGyp8ePFyEGfVd4w==
`protect END_PROTECTED
