`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3fMFqj+C4EJ0VtNqx4X9K+z8ZIv3l4ZGE96SqqGAU6ajg8FlyA5fGlugZQ3obrT
vSJrbbTucgatetMt+WaPBzUoL9BiUVlyzXl3fhOVzVgafUh+3Yr2zgnhiK8zBL0C
l7KHVkyZSPvAwViRKiNWBjpYaGf40MD0uPyrx0c3uDd/MBzToD5jbBzguSovtgi7
qf4axuppJzoo6wNPr6qsvzpAfAVd6YUKJy8wZds28T6HK65nvRzqtVCQgIPiK7mf
6+wEcJQJwVVYCw90YqhsUH8SG0bjdhMFJKi7uo86w5dSVu0WibxpovAli/CRyK78
BnE6fbA31twGblUbXm8xqlDMle5xSTvJBXpCgBmAd3/kKkjATuWrXT88kE5DULzA
oHZr2ljrFRAQdZKi5EU3VM2cD0PtrtFz9D0Sp9W0FDAeoH2sxQZfg5Y1qErxq+a5
6yNWdmymyJBC0jDOHHWa5peKXwfsAcosbbnYckKpulkHUMzA0BjP/PCUXMBnbHUu
81j2GJ8lPr2PuFFLLXFKR5MDvSfoTzOgJtYdSYVSfJzpfSbjNUEge1mJocCx008N
4LWLNOEr57dF7c1sdxUZ/f1pm8M67AdNZ6neveyO5LHr4h4yNZC513F2vibynZf7
`protect END_PROTECTED
