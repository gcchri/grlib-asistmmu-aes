`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fngifoR8/gGtLgYkwrQ+qNVWr3JxzcjLMzh0SMBN8fgSL3QibPm+pdLrmLwQP1Dm
eP9Jm1n3WlE4POtXRuAI4h7T+QUU/RujVXQGh4beFgHZzYQwFcqmB/lxV6fXPTt9
y2wKkRKJ6cc7mmxXqiyvsOuSzf3VaRmklAZBk1c9D6NiXvZgHHw2Trsv3sJWYOn5
1A8IIvVfsUOB99YDqFXJChqgEPxDeNjomU8lCnkWTd2IEARa8ld5bRbDX00fjvAH
htoeVMUXHbvC7s8r5pozmDCZw4oh+owffC1wjKPtjLEH9vLHJaeHkZtTsBek+FR/
ZJFBzqv47Lv8+GmK6d896Mtnegnqea0TiAPzyxotGj90p5I2nnbfHOeE74sAnX0u
+jhts1WAAQqt1IADvs0MLORdOdJYFRy6FGqsJMpPQv/xv/ThC5BtTabUG575GWp+
`protect END_PROTECTED
