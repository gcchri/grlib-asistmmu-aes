`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aNxubnquWaT1ZqhpNpmZmZCW2OHywewnJiWWDUgMud6lxt8ffswShNzPRPsWzOj2
zFi9ug+mPsbkbBMQckbBEOJQbDNmG1w+bpRXJumrywcli9LO1/qUXcfl1E+iEuN3
mvTMpTQSMb1Iclf/5nNfZOwC9BRoYx5pquLkpjPr/ZVE5M42Jr4D4eNZfrpeaLTb
aI1koCea+oQLsg7UErvZv8FiWcPSG0Au3k4NSqALlLSZI1eCgD5TTEHixOBUZEGY
JMWdy7YgqsX+bLmh7P5bYQ==
`protect END_PROTECTED
