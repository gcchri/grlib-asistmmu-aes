`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEFVKH5/8i0AXxJZ4a+z7sAZkhwPbFG/W41c0Urn/Pzl4ldDlCohGGYIrIZ64Bao
u51ySwCBU/FcYg91+Xpe6RMsuQGzfierfV2JcaMxCxa2fMd5N8HtNhOPRfGc+k9J
csuCGyPY+vkpHY7BCVh67Aag+xwtfH0sU4DCEu16DZO7FjUalgSM81yNDP53JkiA
ODxCbhOi6zIqTVM1azD67pHQzpCu7+2NBJn/Sn0eBhFgrwGyFcumMVKhQ1q+WrwG
q+6Pxgn0DnuRm9mQ0riOilZY3/1oBkKeASWi81aDaVAYLjTbxUG9HIW/CjdbJ6pF
YhUDFxduqx6D2O6sZLDBdOkBFqBAc/YRFHB6VLbyKiWYHNNtS5f1riD7Uj6Ufhn7
+63UyIBDMxBo8+mYMldpyDuYtE/98+yO1CDbQDuhCaPBMT1Ba5aI5OiIP4FjKnLv
lHL715XJq5OW5b6H5GlFjBUrDksx2+FSXZyBqn/6/LSSfnZmaU0jx2Y3Z/rp0Bnx
jSGcK7WC//Zn4B+W7ektcxrU7I1o5GdmXGWiafh8kINBSgjSau+se5EDhXsp2uiQ
HHEfVpNKK6lIBA+fVlQu1BMA+IsNpEYLEMQS7XK6yt+ecpYACM/f6Gzyy0GyC+LT
7ve+0kfJ9RhMyNEiHQPTgHuxuHd2WXgd6s52PoxjF0bOtxKWC67zFqqDYkJ11J6P
8XQAb0pOX314azhzw4tpfQJr5EAXK5nl4906qz7nYtzdvliB/kP4UugdkG6sPm/N
YfxgJhsQprphAe4J/IG7IV8Q/wnBh9R+QjxC/6pZ4WxeavqRAJR/hjOY26ZYrkO3
7OUIvw08uDZ/G0LorUe/rt58Zwwtv3BwnG32vyjNEroz8URdI0Km/mc9DlSYpZNf
McYYMwGSmxmXxY/YZ1T52FtKl8VmOj+eE2YxJJdFR4BsRV1n3MTD6Zg30qlXj6RC
xDSI/OxDyRU+CnX/lq84NGYnyZiLpcXgOTQTsrWTD+lzIky0+7JP2LRIBY2Oh9V7
u8KPaPMJy7Yt+T/p3IiNTTA3vVB5+POJ3e3WiWbtfqzSaO8RRVtiYCXFFCDp0oEI
JLFL0yCWdRfNxDjnpEasUa/tZODalX3O3N75e5XABbDT6CJHumllzBWuE7bOcmV8
sP4SUQB8nd5SlWmbcT6DLBLYptj3+F/jJcWY6KxKBgWLzWvRPtVEPNei+/ISqIBB
v7WQ581cTwkU8x+EGC0dlxXRhlI2pHs7oU1x9y9R37WZ699kSqJoXaCLvv+LqUuM
h3pAAR58dXBU79gzF/+wZNvDeMShapu/inyXcSaFgOlnOWCWI0XfDZgBkiN0wy3a
bNFJIBBiuxF9pxaNmwJixSoIRERptEXA+jFKKyTqk3AgtVKqxsgCWuBE+V+s/hOa
sF9pJdZRP1Wf26DcUacNX21oul83T0jMLv4rl7CEweYZgR5zcLHfqDwMygg8DO1h
w3Cist6+04ka3zbIIIoFbuRXWh0Kfja/p6Q9vjOfc9ipJdXZimnU9/7cZPqcBDsv
V15SD/h+S3PdGZAXF2btujfKor6Nzjqrpbe8MoRnczy1UFNQVfYmZEWRvKFK++jk
QR3RwJb48ck37kBSrEYT7Pet+toSJ2ptk2l7IbW9Cvt3RaCIG5FNxJ5fMKRzg7Wj
`protect END_PROTECTED
