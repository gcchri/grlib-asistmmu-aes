`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TM8s58Pnw2/4ztWwDfBWxRaC3TmsXAtMyY2rm9lARXgy9rKkBTcptU3701KMSFJZ
43blY7qRtrhytPcHNiP9pTs4q0TYG01a+scfeRHh+lGVk/zs9JwwG+aF0mKmMVi6
DxTaCP7T/gHD394MN2a8d9/8Ifax5b0C6elKKut/EAy39dLjoMN6s27T78UNI8hf
2lJeaQqYFOPMvSHlteO2tYbSR83pTmSsIn8XZPRFbolL97yPF8F6ffGN4z62pIAX
jlCUEpbDbWrchXX0m/HD8gnnzxun2otbjTm7smtsNlkzgoNKY2aDCujIHUIZpOiF
P2voKOTZuzGNWxLcZoeX1A==
`protect END_PROTECTED
