`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5a0odX+3CVYefmS/zdUA2CZ/vUB10CnxaH6Y83DrfZ9/+LKKZ/qGi1QF+73va1+s
R1aegtF53d8DU9asICpbE8ryr0G+n3Tu8J9Kqz/Se0B2Y4q7sIJwDGQe2IpX3LOl
cR8Rne178/217a/M+YvmYbJfLkWLkreHJQ8cRi0lWHm9bfICMAFlfUYzDMrAk5WX
E4+m0ucj4kwb6pPfM5Ia8xhMmWOnCzewT8cab+ECpsGolTKI4U1gT4yw8PTD0aWB
KUridADrFNsBjGp65o1EyN0bO4rDerWV+a58/EAk+7548LoW8jWyx9xFBbRifxj5
El50U8usaljWQPcJvGZOeQ==
`protect END_PROTECTED
