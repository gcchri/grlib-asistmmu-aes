`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1pvAWsC28AG73MkHT5G/Lmba8hKMPvdEVrnE3AVszx2WrVMm9SAt/KVnjgkTfgA
moFu2L6Hu8ZCFMWuuAbQDypFzDk/GNXWNfCAqivUZpqgIZ7/m4s+Y6mzXyrFRziK
R5UheBbkQTAAyj5lKHUSUIWzwioR6N2Y18ctMrqfNy1/qKRrVcxce9Sl6h1pcTYm
ffeOX5PqebeidV4CDCY9DolnLPFiBqQfJxgZUNCEEKiH1RAjAUzDPh3kshJcZyEP
jMpM7b2tRh6xBa0q/GMfLX3OnkQdqBUwVFlMhfbJbuB3ns/QYADM0UC6feOHsO9K
oN455bcdJaaUxkhqch4Pu3RYB9K4MQ098XJtZAPrAvVJG6WAcjpoQzNhs2MJmhYJ
O9TL5fuow3OmhcfqVJnoHZmo8lH3JY7voySW0JTW3nw=
`protect END_PROTECTED
