`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuhbG5EBoWN8u8vFZzmhKKFFGbNRfBdXU6xhEZm0a319ag2RX/GnjaaC87qyL3wj
NTaveMD9Tz/LKpN+oqNHBy/ncx0us7G0VLKasDCHffi/i541bcgKtfxQBO67Q1Du
V4V+slnfjHu+llcOKJyNfWOtylTTn3WvKDDoIE7t0J8Qz2mXgxQi9JymEWkCcmLv
rW1ZtTKwG7wIGjuGlGcOQ55GzLWrSr43VPGz+PIBOgQ7WZFQ5XPCV+3eKRDMumk9
zVk2+ZwtGS/upcCtWUi5tZScoL2XQTe3YvN7cYuuUjWue+l6tJ7yT0wlYu7NOrBv
eAWtgQXDVUh7jU9gdVTibQ==
`protect END_PROTECTED
