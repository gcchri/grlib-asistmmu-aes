`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVNZr0p4V/NnqrXDOeUtgkIoHULxuhIT6lBME7M+HF4p6hXYmKMN18NvGgeMeR6r
uzZLVv0iC7WCz8Z9W1pA9VqdVP1jcPqPc65Hc6XPi3xGXZQUGWR3EWgQOriy9StY
jPVJFAyzuykyBrhPxKMPpV6L0yWOi61/Ml9DpEKJzfR3dLPhq4OMHPOZ+TM9oLrE
6zbMyt565R3PvP5utPlPaNC19IdScD70goyPvHd8S9mWhaq0vIomy4POhyP72UOn
1MK06Dg2pvZOhEYRypCLew2P4/fbQAf8+Gr5BQg5/ANiQaW+gHhXJvhRGak1A1kI
n5VPrGtFKASBus6ckEp1qQ==
`protect END_PROTECTED
