`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjyHqvMkR1umn566kSA/SOp+RyvyosPfiDus6Crsdb8ZjvzuqeV6TIo+J+reLnir
2Py4r1tFOiYzueZaHYbg7SV6bYoIj+tjOLGOIzODveuvK+pt6OZU41IEdtKvq/rp
26Tn70el6aw0zfWAXc14DyjJl+DH4BAN3hDiCKwtdN74NOsivmaNZnnGRSkRIJ54
PIlT0V5OsMJsp+1t5TpgJk19fR9LoowDAnwOpqIivgg73z+CDqXLIEjcmT7D2dQ8
Er66cLdNpLk6ltQ8YVaop0yvzZ3ksq6vbN8g8XmMglJ92h52fnafXx5pWb67dp7b
OcsNfGFVNNS6+Xq/inXI3skPQjbS3kTLNXBHjvkHguUhZqicfBUaMjh2lnpDupN9
tai+ez5BBKDUXyz8PfZYqgIBJDzj9ygmWIU63Ypy7hRiZgIKEc/v+rGyOqT8xTtU
tK3+N3Ri66/bFV8nf4i4Zpr73v8CYj28m4DAyFqomyIfE8u5RkSQyRkNwiA9N+5i
rzboFqGQIUEmf5KwN3jZfY3jLysDgzMOJXkCFk+p9FF/q3vHd4yaXWbRsqDu0J/G
ZsABUtKLpQEJdnGvcddgzg36fzhtH78UTkyKmtJRAFkDBORsg04kfp4Q5vM4a2mQ
b/wVwvXB3L0bv2iS4BWkTBsAiwPINO/g+2UrIbqjVjs=
`protect END_PROTECTED
