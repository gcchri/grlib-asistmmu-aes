`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nAI/Sm481EIqJv2nGSULNLQk22Ye62ws9jYiifAsnVzY5qu++PZpOkxLkUPIeP9
WnXz3G03xNX0MxEr3DA1F5YjdqWimUHuHu0WUGqjtlooNuQKND0a/1YIopvTXymY
dWBglQ8mReV8171xGiDe4NLsIB6OAOBtf/JyKOATVLigiOz2/YPdadXiBh3Qc/BX
CaIlPiqkB59QNgG9uP9UtiUOWovy9f6Rf85+GCrEWAknKksLPRXzYBdFed/2BsuC
ICmti9Fa+eUbMUwMUU/nsPGutIGV33imXxB3XnlGA549Z7rB+rMqQEHQP/Zln52x
CfKdV0fxNDYufmUaIEKWvw==
`protect END_PROTECTED
