`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
++m7udjmej34TnXj6hUCiTYvwsjzvTQ1D8AGpZMOZFmvUhCPAjIdX+YsaQfxLxPA
YXWbDyMmLiuML2/FsfW1qTrJMpZNVmqWHKrl0LYrODNk+g+YCxnM+v7EcMMa6v0A
2h+Nq/AjnVgufdygMNCrWd14i7n3bNPgqPtmwtpTk4CT5xCmkxzoeak6o1B0uvll
OtlubebBlyB7GeroiDa2ouhBZIZYer/MGy0V0jD1MSysUqdx2Ysdg9m2R1i/To4Z
JWGfM6d2gO2mZrhk8H3kci6Nc7qkAdo3ZKemuQyP0pZPNQn0bTaRf4YeuWoPRwa9
vaEN91huFWA3kQn8rWPzTPFm6hbWeB8628XENpCQI0d45H+U7YEaoynhvHH+6w5b
X84rd+pxjZ9yYAoxV1wHaOEEPL3+Wjx3B7DlNiUWRX73KBKezaP5RXyUxAp74fkz
Rr9AwhKplzzdAEXcU9kJvSe89Xa4Zb8q5cKa31Uiejg5QSGoElzvcOQrT8ujFvW0
aj/TjaCI1suhSJJOAJ8RV1jG3taxFHbN6ViKwmAi3iNoQZNagMsFS93yLXU1X9Pp
piz6yweevNcB4Jk9lt8LkR9EB0q5SX1spZr28fPgoDK7pvxKfpX6qVjLQRz7uSew
YgvbQf6W6CmWzUgWGAZnYSzz6x6yCmNz/UxsTfEX+D9ZXRwehgeqJoveDom7JVii
VfN7CeZBi2qxNdfb/rEhqjJnLT5qMC2La5PdJo9W6LDZSLSNoOP+8qlvaK5hEkBb
`protect END_PROTECTED
