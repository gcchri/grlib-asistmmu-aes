`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
04AktvO7Z7pWNXknAr1tC/nETBDZzOoauPM4abfZZOtl5TyV46Wmsh945MiL92+U
yHunEP3GA/Gb5loXHh9x6hTuV21ZP9EgAmBdW7p9roklxoEffJoRKXByHWvCMMf+
SQrhOLXT1p34n99LPZCcIegEeYZD6p5UxAvh8yUNjYID5rcrYztD+MujbPr7PruP
EbZb7QM0LAFezZ9e2j3Ev4Em4nJJLcQXVHy1r4Yb/3vY5yGvWZLlpgGb2sQjnowu
Cz88jM9JyOXuKnPftAFnr/chu90SUeoOUBC0M2Kdwcw1UbaF/2aGktm/h0Nh3cJn
zg6Y9iAMmCgsx2OVywbaDZLJa6n4n4H60vc5hPcOxh7lSK7ZCwvYnCRVlIvAt4gd
fUKHmnOAJevmuyS3ac86IV9ylbCpiOnIrB9BrZzBZ95QWBuYWz0lyDNMStu4ag/L
ORKZUbAFU7M/SmvKyDqZd14rGdXu0VnrbHXujGzvktwFUwr9xLG5coo5pbTO5YLA
d/MY6pBLawABGAju9bDuWTrFOJS6x1mptnkH4EEPwDWCyRYXH13fvtSLSio4LyR9
1WJDrlUftXmZdhmVRBmOUo3Qpf6XcxY071m1/uSsraLE3bj1oW9Afdz8wHIUDXWT
dgRfAvRkWlpEedSpg/JOTOGpFAZyVzANC+fDWPcNBXtUveFpShCZsrbboE3llCuZ
C1aS+N8wa/ylUTuZtHs7LTIf2bvOOjOtc2ZbWzzxTRp/3mRLWUiUSX6iP9IpyNre
wMkjDgTZnU2IaGHqydu44PDxVjLlO2ptnZBYGcul3il7QF5Mw2WcU2xS+Cl8dGwl
2AfbwYooJA+6s/HjpSfkkdWxSJaDs8hktr+EVlVH2fk26PRQad09P0gq+kIRsJMu
74+7Jj+iYcbJrbRJYF4ObjoIuzlEG2KA1Ma148IrJRieceZD+XBLimRpT3D9vJKO
24AyxOr2OKa5EoUA5iX0kA==
`protect END_PROTECTED
