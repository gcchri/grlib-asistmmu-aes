`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mmjg6Vs7ebnwcAGhRMiG/83KC6uLyMjeWOPv9ktiZEhdISqmyNqX6WoyscvAVf2R
89WC9icwHna0Yqw2xAOV3QFqmn/OSE31ihQ48uUrJ02qWB21w4KPrQWfK2ct9N/j
H4HzovVpONZ3zYOku5B/WkvHDtN1Ju+zC8oJB/P/EPB7AkPHU0t4P6W8r7Hk7P9O
23ES818zuLSJ13KuRIFeIhf8NRPBX39hjVpbTQhFu+6k919myZUAMVttClSq3z+Y
T05Z5C4aLE5jYOzVwyx6ZzWdc6Ncg1EvgOv9NcpcmYThhVsV6dnuTl+mIWenDtxI
Uu8H/zJsVEJEai+QJSaduLFTlcH5iJy7ZrkJnI4iOvzR739EwCMubzFAa4sZamZo
12VJrGYHgnvSRCPdBRHbYXZMPfXwTLWjqFa0LbEbIG6Uc8fT6f6qxgSagGDGc4NZ
yLVvfzjDopNJZyiEvB6inw==
`protect END_PROTECTED
