`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzyWyqieFHXw3XByAOrboeFLCtNftjuACvTQfhp22ds3pLbxdFeRSN0rJjD0yrYi
mGIYmMLgaLV9D1xLpW2hDtgqC3wYmS4Z47Cc0ZpLM3/CXxxHwPR3q06L7jvClcAb
tfhEv275O4oWWt73QCQIaH7OjqvrWcLNyhPP8awuFeKh9z/IwmVMxUN+2Wpk34ok
1u4w7TmT2OaqrS3IMEi4W3SGvbHbtnFgpmkgELQNN3ET0pfMkHm/OggzSW9vZWkI
ZWkz+tSjqlZiRHb59DjGMvDv23/IUd00iWvi4nkFVrMJMLLBQ7Y9IszgvGM/1Rg4
/On/MGd1ZpTfkzVCqWku/fMKuHS8sfkX9VrogFpx+XqR1YcT7uDi+O8s8SbOIprE
Voaelip6Gxu9/5ZcTxGJgOMurTszG5TYxlHSdK9qk6EgkKdpnDI1evLjPod1J09d
`protect END_PROTECTED
