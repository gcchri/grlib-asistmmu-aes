`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hQYQyemx63ywHUrdT/c9B42vP+Vz1BAV2RoN4UpDegTTV3F90IjySY8zMvZ8V1zV
AMVenx4OftTe257RUaAhrdbsqPqFPzyh6eBhA6z3HK93BQfcmZeduKteL0ismBjb
iVFe7nEmLi0Ndk6/HRNnnF1IeMi/luYzKX3IjzfbnRN+OUneBbhaRPzeUZUwGs/R
42ffl1MjMgGaTCXpw6BnBjj8dI9xhDCjIzlO3Xs3CHTJz1W2GVQGUrz+SJ+PPES0
zsGEtkQzcC0f3KR703YApXvysbkB2LeGIki9x/L0IWIq3ik0EvipXngl5LxQIrc8
B0mqeA0xAohHNW62/R3kfNRAlciJveyE3N7oNS3lO+I7YQoEXqFfJdna009nL3z6
zsBMbrulb/zPuVXgjR2Sz2CdmdZL4b4HFxAaPvNcY40ASEUvx2ZYEMT2I8VyUHsL
amg9NLRefgk8ylAE3F2nL+oLFEdwoHxXU8ewHPbsKqM6a82I5Tp8rhWlLiMpuPOX
55VGemkV56B4pMnlfsgJtQWoTpypDL128MILgXXz3KEO+2Nn+gboYKlneyr78Zx1
OZddaAth9+RWya2yopjq4QRqTFmWZd2jmYXVU0BlVKnV8T2IjYqywBkFxVEdKXsk
tptet9gwr5CI3Sd07E+NfTsyF/K5RS1hRbkgIUnjGcjiUPpxX2FpxnsH9C/9OLN/
/3E/HHcVQE5uPxHSER4NQkS6lvZMcZrCfUw9DDr1eDoRLxgNWotU4SM4Gsk67SZU
sMQsVCl9YpqBVso2sQk3OiUtRxy6W55C8OEq5p202cK1h1Ogpg2yvKHXCnPlthPL
pTn3oEdgw9xS0nmjVspHSqweINyC9nUUM+OdYXU+P/Vav8eko/FIHjSq1AlG7v1e
dbiCOeBmIBebwPQmk7YI1Adw14QWuJBLmSv+/pb/WlkgxRH9YYeeT/kPP+qbUZJK
I/GNNKPYpEPyIN3zm8n+zDXwyD2/7d6j33u9bZLaDPhSFsGvMFoNCpx0fpltrlHM
M44hTw82gwCAmOCigDx0pBTo7FydPQtJLepaOipNzI0=
`protect END_PROTECTED
