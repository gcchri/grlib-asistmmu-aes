`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFdW5JwcL4zZE/+fDp1TKTuS7S+iDrYTPcc1Wl76JKDlkzmB+iYqEQY/epxt9p6S
nt/hK/3p07ccjiHTBaQorTMT6YU5nQ5zZXkYj3CjexcxDfGeQrOqgzB55HSCgPM7
g8XtlcnoScDmzgBshU4qn0R5Br7ZBplSL61yQVcsEoOm2VWdmDvd8FYRsP9Jpxwg
4kpOprRmocNPhfqWn58ihtEx0hwKhjhpei8ULkofFtaV7udkyP89scykJodQsOU4
OUqn8b83G5KDK2AaJgw1OAJPFmpf0Kik69G2MvXK3930KXG/jAkPQ8LgqsKNv2Vq
xEleugFp1y3tnh0fGZAAuptM7pIrtxr5rsHSFMEbcHH76gRSd0SyaGltVyG7HDIb
WpdSgwamXFe0TVoh3cDiyJGpkx0VzJ7ocFbMV4Utby/0yJwFMdxGfsCY4hEjs+Fo
AXPQviovQFQkPqpBYzPScOK9ib99H6CPmx46hyx2wr4XwHOrxMxAye6AaekW5yMU
kSEdK53etuTYEyqPvSBaQN4+rVucwuK7u7PP56STUdoasgorNFuHs/5/+DTtYvsz
Is0TX5JdR1aWkoLvjqc+G+Toojk14OtHPrfpCE+5rZm3a8jydP+ahdiF/stVozgn
HsA8rrpaoZ9bux+neEROhI1dUjjdQBtUvy4h6X96z8K2480Rdr4nbdIRErG6WQ8R
b7K80NDEHiVX0//FJvm82QZbSFy+KAzvnsevjsvJ5h6bnqOLx4Mna3FmYuOw3A7z
s+ZTO9v8uzPxakAYeKAKNh+hfIBmWNS6DUlP12PlNhZNoGnRXKY93DS5UbP27piq
52xUXyXz3H/q7mWN0kaIkpFRdtRBZ53M/SAzggGzYTbxJS7iqzXocy+owDh9CGWw
Ilt6s0fL+ZtnLGuvoKZNk0o5snRfeZopK/ogsqs+WWFCShSm/MM6+Xp0pkCpFDQm
4i9VK3PA8QEFCdmOLUNAJ1WPuILrrlKSu/wpEG1U5MqmKe75h7Z1fwc2qU1CPgpy
DDvXhDtUR9mPMdimwYnLPerKV9G4ZaEL8EiQ5hh4DgYAVxj0gQ0tyKtllJCOeRJE
v+NZ6ODLXfuY7MclJQRjRWK1cbAT+eFOZbubIWJnTZyYUrLlQJ61nykyZ/VvFzkT
0k+f290LebrMjUCexs7IiJOsZE0kBVS/wWwic5otWJko3wxkpOV28gLSQ6AEnWjH
AaBoiMSEKE0ms7zlpNHTnQh7lGXNI95VSX1G3v0Kk1Kii4QUt51KFlnznv6eTUs1
dKS5TzkrpVKyHYIwoMMHZG1nuDtGwxrOg27VNo3TcbvFEiPwhrGXyAVjptk1ZOK4
p/pE56CFGMnNju8w7gDq1qoUXoYlAJGBgADBiu9HfLxa3mXsQfYXBM8kd/2pCZjS
WMNuLpcOQoUAY6GjCOyA9PcgZxrrnfAGy5k3PYGZzU3MAmwYOsu/kvD2ZVXajRkr
9BJ7pjy5SiZa0p+5uaKjrTxQwc0cg62S74rgVdzkc8SMBMZlWl+oUiBnR4LrLUef
Bdg9/yySJHbDMqOLAXHzgAoAMIJLbzNXo34Va1senPYjeKBkz8EZegcsO5rhiRLZ
79yei+uqn145SWpqEvtmum7k4rpmxOf29dpDeJlO3DMTDLQyH/yrLOqec4aadwFI
fHw/LCWL3Pfi6VRrc0CUa5rfaLqFm9XQ3/Ny1Ze3auEn4acmub1unnn7uis5kM07
12Ca4PiUMgEBbV95hZJUik/To0/41ExL+VjEZs6bf7RtzFW8iE1KdYDcCCKXm3qf
o8/2lMWv2YzJqTiwpldFF7VLM23MzDtlwDKrunwxOBNOuZRJ8z1YcP8/nNHh4Iny
NOnNcYlWckZbNIpU2L8VuEOvU0d6DnhkRQalY1rB3J+/ac+MCPK0lb5L79uQ4NBh
gPMf1hscHWpKdbnyim6G1rAKcqDGn7+Xkf0l7zpnLGujBHJw52DmW0FnzDhPzYaS
XUXVLUlCcuwR0dHamkMhYp4ezDSgewlOK0Lg6A1U+80ugAh6GrP3e3sdEiBWVKNK
EEyJJrdrVVkDkldV8tb+CgAge7CrJIBBAW/wO+EMNKyam/BlUZ+TGfbHHq1hm3WE
cPePluSlM4hXpOq18iHe/S4UUQpLpmqHO92f2vmRSR7AuT2ymJBDDEQQxxoR44pV
WW7uiYaPwU+Ucd3x0mUaggDBDtucozMmhYmL/4vq310Pkwmb9blc9ctcut0E1AQW
0/mukGOifa0rsIfjp7jm8jIj0tu4QncVdxtK3SisyYlf6782RCzmJ5UvvdjDXEEW
JfWjb0orkZOEWaW4SukIs+0E/VpBQqXM/xqViIKvXAfY9vSDb35UH2BZY31Q7qPv
n1WFcs4g3IlT/y8lQ89PpuAwDG1bIwJKe54fkbq631pUrYNXFQ3ivQ3wm5pD1KCd
zJ73vccEJQ3D028X6WZDRaNiCnZRQWBeQlHg64/jpeH4i4m+QlGeBBfr06NLgf/n
QfDe3YGXAj9iCTwcELmy55qz6TmtOaiXEe43KtxgXwuJ0VUUsMOTJ1g6jshqVoUa
NxAqqHxTMMDgAPEt53cOxB+9m7aulAmvlJCEy6GqRaQiEq9DlrC3D6EXES2si2eS
j0liaiYeDEmE3FJ3Lm6HVdUHe/JXSjLqSWlLCcykIFyYnU+S6+vbLwOiWTcx4wum
NPCKOLcG6TINGkuulFeiYnMSMr97og+FHk4z90HBmXinpcMmZTDOunOM9zZJSKD7
yccgbKiVeD0vAwtZW5DfTrBUW5gzL4qQoTOZVhXuBuSYaWed6Gu8zy0b5AsIvz40
EW58yMx7l9mSuilv0HOO/7WVZSgOoQn8sRr3Jg/FXYIrJv8MNVy9qMBv1SPpFpDF
hGUFxlawCpF37BiB0smE+Xxf9M4+1S2Bl/uhmzS/34u1BkF0hpWl9kjMFc0Pur2Q
MRp7Tqht7c5GqkwZMcdMyR4BztKOxYTje/0CyKyJmowBfCVWnZX3JhKdEzXY44Nq
f02wNnXsmJSy0wnPF3Swz8E4WTgpD3POkkgGNz/xRNUT84kaYbbDz+RpurtgrR2/
DCqx5jwOk9U8+GGgeGoiQ95ERqsTyQZSMOw0ugq1zGF+TyelMp/JPnDBpw/QIC/v
suMngrECdzHDrZWH9ql5LXMk/Rumzzcl7GY/kDJZQtHXW4w4hWZAxvJh1x68kygA
0AbYmPi5RA+xsrcuidC0VCEDLrv3WWm/LJ2VHLJHM2i70PuhHxDRUA57Uj1DJLSs
xg5uorWDzTmhuEJWV8jKMDkqBNK6pwCAfJOvEWUOaGK1UBHLi5pGK59WDAjTSFch
NKat6JuXIXoM48dzgbBcJmvycfL+9jBURzrVesKqCMKNIKVPkvRQhBAfs9/S5Teg
msGlVvZZqFIfBoKzXmFCkfUiS2abNodV+qeRzRvKWCCqyAiH9Rfdy7T0fdF/GynC
VEjCXTCn8FmVYPP4j/71roilq868AgQEqK4UQbS+/EMuWgzw4uKVcbK1LLhrH/77
S7mRsftldTIA1TWyTK2Xo5uGAE2jmPjFe8Ip8IgNlrpvvteHGO0mQvnE/cCcF9zn
/ZO16dH+882iYHFb+CLWjF9X3HV4D1Es+aX5FZr29U7HEoEplTxMgrzC45xG/r4t
+FjAdknN9+2UUaImDBTcEWRdRgA9LkGhuuTets1+dZordaEdTXF1j51R/zv3Yje7
3IRWmJdWQR/gEw8Ofzb6N7gXdJjSVl+PMs+s3D6Li8neFNY2/0f08c59XWN2amgJ
UCcJGxa3xmhO1uA2exRK8CRZk4WMm+d9c3tm3hRk1vwkRTnNkBWWxkPjw84wIgMm
nQo6N4+yEmXN7a2BerGxKeqZ3DjttBS5RiNFqcJD2Q/D23gtJEbNFJmIYy4HFKev
RWo38DWGXR5F+2NyruZ/+ErE0wwUv9l2s90i5ctJanrVSSRYgQAPxDy/xe4KfdAw
OjQYiBGVcFvUk/44UQdoLtcCk6f8TU4njEXDoHuIJsLzgT0cqLjt/KVtpXItw+cB
1+TVknLMjoETDiXv3t1qqkHlrQ8dS1pbfA3tEOYBCzegZKoSt37vWuzOfxLpwWC8
IEhqAIbAsVkERgehHYQW9Zra9unCo/aRNh552Ue9Zhr6WCP2adJRT+VeJdDuqOP8
dq1pItKt45UM9V69u/LMr0EoTdm+5EbFrEFUfKn3rRadfLOxjM+DPQMLK/5dKoo0
jlio7S3SFEgeqDYakELkmP6ASEW+rjTP5Zm9DXbu+kB1O8FYAPoskIbuvYceLGPA
2sKBC+RYuM4rCAXYSdr8JV0HT56G6wjRnpxbNEe29g3UsiwyL8Tqyd8cdYymd0gh
KbefenqswEYDQvuNUv0uskj/ZjsUyYAR5CXKix00+sga6/NPDtkpZaeSiN4TL0dt
Vrx2YSUrowhTtrwdtPlm33ReCq/l6ob9RlR2LwM/HSWhBWCqCYaKtbnCIXQzA2Tz
Wuh7fHuKcqfsCcXrxImByUeGSw82P203Wuq4kcrTkO/LmJMUS1ipz422o2APaLau
MmG/fzS9gLPHgzMsUh0pbsIULRbEYIJBrvN6mbaNRie+XaWL3pqgeZhL1CBB0uv3
6OS/MBAkBEQ9mXpdrX/x3DN6huOdGFaTfe4K8488fsGZGJY8c+xg2LdnH37QoUxp
bBMScRdLtuPTXmiRQ/WBuZWhyczPcjgaoM/ebsxvxu8Dg2f8+Ef0UZfrctsOJsb0
q8ycAAnv9ZJmFbO7+xj44KE7nd9Tzzx2MOrbKjqwEiYg928uB4xVU+dPWIjilZkY
DKXxdn+MbuixSR+lXcV4tB+HZ3qslfvLDLIXJu+j0xNsYorpgpvBmLQUaJ2jJBwl
0vh1Ltb3/NBKljIUeDxTqXqmevbu8vf9TmYbV2xTXfKwENevzLrGar9Np1jxlHe1
1BDc5UoCX7xA/yzUBq4d6POk7Ko1FL0jKzsDz2ikPMcoSWND6gX7F26lem6PWCPt
6dyfxBUPFzWNcdrhiInbw3HcAzbVCALbYn1EQ7vd7DA3MEC/QZYIBcRDfL6+jiAU
8t34sFxkfpH28idwSpK1PRHwzaIKdItPcAPO2p16bO6l+ns7CB4ifKzvZx6w5p/X
dh+FMBSbSqdeUcJZdl2FbdIIhawc2vm35BfFTrTbhjlEzmhUct+gAd428/lFUvQu
3UuLSclWFzKXLmhNZ653XhSlBMAVO1uu+rfp9tTtH6PCJn2DSBbffiS79IWqKTrB
m+YSosut50Ma/e6FFhOMAcsE+ypCpbmRZptpMcMyjtn50ktR86bRtzB33+0WPZT4
I/rPmSbhHqkUxysPeOv1qKMskltCorAjSyfrkrxtexzvVHLJqv2r21r24CZR1tAc
64csBwb5wea80E8EtUspTDsH4MGBBbxz3z/+uUYYDCnWoPH4jkPCb9SXm2odNABq
is/GZDPCrMoynfK34U4EzA6gFZEGgzkbjW5tSsN4Q6YKNRz4elffscVi0C/3hOQX
ipRBCuOXVjgJpDKqxy7z1uIy4MPaW4fZiEMdhWTJ0BzGR5NTyXr2pTXnTF00Osyz
qaSfDsVivqBJlEEvWh9aaf0D9JG2Pu/SCIhTV7EcKDwRYOUQa08QHNcM9zeSByc0
8/QWLiBQLYdXObY+mXcBSJX3Qo167owTfu8NN2gP4iuT3R9y1LrjkB0J3OCAImkc
qlkufnSjyoF4iG+FVCrW/RPjXM9qybcI3z6TX9k/SNmhgAf638v5sxjzKHSBwUU5
p49kwHoqn6D8FNZ23ibRlW5ta2gT3w2Ep3kpg/IUIUmOgs/0g/oHgTe91JX8z4qC
nYA3d1Leq/UKh75YIxhLLDuCFv2eVGxA9EQa6aPkqZtreqV8jk71dEqZBGg7riG7
FxNGKieXKg+UM5gyTF9sQYOSxYr3PPH2yJgtOeh+HQIV21qQ5+Uzt/A8MiwwwPbC
f6JRK3RnKlLqNgiOHuDha6PxAoInf5y/3P9FLiK67uJGnsU3D01M2HwHtIuYAPX0
kL3e4HXc2+bFKVVcL+5H5L/H80SkNS2LCAj4H9nUPk5CznDSjspDr9f/zvLA3qVG
nYZZJAFuS2uf9tbUpaQkA9q9rOXVx6xTvjcgAlUT3zgo1zvnqOck5eJBZRSiUid3
ah/8fzo2RhSL9hfvWk7sj6feITumny57Anh1XEYA2RWHTwbaTBsmR0Z6+IsNEZ2G
jilcWwNQsW7V6LoFxYc321LzGfWth9BOhq9a21kw5hpFDvtcFMbaLkKNxXB0jXfj
ncKDx4l3SlEvYihQ+U3pqUmPXU7yQSz+vXFqw7vDyL8nLzrRqKxCPy3ohRy9/lJT
gxy23v3zHMzoFdl2VhC5uyL5QuSD2XR+DDI0K7JqfnozeZ3TUSwOAgK5wjQS9fy0
wU35qPeIvtehyofCmiE5KLSru6cYgY+q6sOIAGePW+HBAVeIRvCqhu/wIWciAdZr
FEGSzscccoE3ks0IadxNnniQtqAxdME+Hm86flZa8563Qor49PrlXehSkoX5SJWB
ZZSDGop9torXhN3Ar1A5ZxkqLR9m2K/qSMkXLprHebjNNB0Pep6onMhEd3PMU/jd
Sp0qFHT62xv2SP72IXkuJEiP6WZTU1CoIxzCt0ziyJ0aW+ztUo02MD8eDpjIbk8q
JX9WcAFMlOvv/doSwa0s6lYj9hywR7yXHX1A+9MQG4+Qm5fTv5TiIxnaeRkrc3Dw
LAmwWIXFK/aREsjba+WPOwb6ZZEJ3r/F28p+eCHawK5eKjF3WWOo+OKpf/0JujQd
ffiRdZJm7MLQzVVJMZ9BuJ8NZwwhteFbNGLjVd3KGyiSsWv1vYaE9VwmI80Mr8Va
QVtfLWrHmtIkZnYt7sOVr2YEgWs5oXOW4ts81vkKbxHYwnt4J0c26PorKNu6lahw
qIouEXzuufJAfbModOHBcVmg7R77mCAlfc6MYdjQout9qMR0bOGdnP9UMb/Bj0RM
6EnxGPPFJcIVAkdjSAwUuM8q0ZwspxnIdy4asMfQQTzAdG4U0x7rIYUdyN4RUyIp
++4RifAAEcugXZA81Fb9SOqGkvlJIu302vYF809WMq762ero3UgJ6vFvLh5MeGCC
gr9RtabUvqtLUKYKMho/eeePPSB60owg3xym5cj0YT7obDBgvV91SuRm7sy2ZFK5
I646ob5bB/u3jbc4BLZHmNAkP5BjzSPF6jogwPutJUzv+xys2jWsGCtMuW6MihJU
EDhpjSB2scLr0IOUgs/mwHtIEvFAI85/UnSAMC3WL5DDwnB8690AxLUbkhpZE4xS
ZvpobByab924ECqNt62Ef/s2njfdfsfF+bo8XCvh/rN94vKIBfRt4bewGnNF67+I
FZpjW6SAWgcwIO5jJTZK7El28owwiJk6cI4FUZ4obHjpRSD0BmXHASMsHzInXAUV
/gQ8ZE8mUq2stZAqXBZIRUso+t9RtrTQkvAnbbn8EJf11rqGB2oadTDiFAMmDcTt
hlGuV+XzyLgiAxDt9lOTAtjWPANsPLECGMbhv3KEB2wMkNo6P6tcOMfptqickNTU
zmQe7JvqOU8ygwG1TofhcldaDWLF3ZyQ8XupH7BWUII6C7o+tX6DkR+5f0uS9ODd
ma381JUP9L+dZu0OIXTe3uySYVNe0urXT6dQ0nkgEtkNafLO38JkUcXy2rKN1wYo
I8WKPAE9RgT1qLiBqOVCMuqcNG4krjlFPNFNgGxN2h5g/fYkx+My/haRGZxLRK/D
SrCXLQMGVkjhl2lg3JHq6jSJPC3LueE0E7B1IsxcUOYtMMrrc5uLggCjaRYAN9am
SJdu8Kvju2l3To17+1kEr9/48vtgDqjUoEUJjPQxmy66xGWIkkK1G9cXDjXtEi7Q
LAAKL6WmBl8VeviIllSYYVis2iz2SYe79mZ7MUplwca8rUwGN4oDzff83vKsw2bf
eBm6th8wcKfcIAI4kzt0q9XgrMuqaNEbAIoRCrSAA73/xqeyM7THxRuc+SuHPk9s
NdEuTpZDvKDHYXomz/7BNqfLJzuafJcuhmrYG3BIW/SD89YtYhtTEIkXD9GTvCZT
hRZcAmhzCIMaweZzjjBPsQcg46SizW49zygWQZS82x8rlb0RZkJJEk568jyxg6Dq
gaBx5So5I9U4gMJIJZRmkLAzuTihQiKOShk/rKrVwMgT2LXQKfqBmoV0/e4Pwe0V
vvSO+g4+ZfDdqGXDC4ZSEzIx7sFUswh5Rg6XaWhFEgfS0/sTZSCOZh1LAGh7jECU
z4LetMje+vz5crpC+kRqXBvyccSIIP2GxvJQITI2Yt5wdzc/xxRmJlOYEnoPe2Iu
ITFiU1QeQBMxvh9rRxAKzVFnhE2tyKggf9ehc6yVEve/VrcGoJurWp3ydoaq2vPe
vitO0TMLWjDe5B6f6hW2uivW/N33lgBAM01Gz/NMcY7j0i/r2GM4XNHF2ujDmhvu
ZYNEjS4N9I1aVFjjie9Ft3uIPIEreQEQgdknaUXDMq2qvBh1Y8xcyzG0oLBbuKN3
O+UBGvCNR7YB68kSxd4F2Rc4Xj8IcFoIbAFdzaBrCMUPPzq+JRjGJDcYUw83OE2S
WGdoeJ5zTxnM4kU9M+xcoqu0waVK1sitUkvT+wew0VPAOD/FdRUw6PoY3Gsuqgpd
9+kCPDLrBjYpRMfF52eaVNK0X0DuAUz+jR3A/fjRPqMzLNuWHlCKOl2Gf5LLtZAY
g4amuz2oAxkpNlFCCJudJeY9nFha6KqjJQy/+V3WjOl5KIBxybYZUmi9jw2l64TW
zgSjPPI03N2i2AtyywLjShkIs9Y8nSnf7H5gpu+hQDZi+2Bgf3O+RPRCVbnJoeuf
8Ue14Sbe/KvtO+sQ5ij0c3ejediC64WRBro8cegQnQYGQQbcu4NwVhXqwCsaQSKs
sevVnNNDnQxyULrFbP3QD31qtnzLc1pZbAaH5TIP+AFLK7grvqKD7MXBf6RKr+J8
aFSYwcEXNMbrGEJ+WwAELTiTEpjZatufzBKqBvmqhXhnBxlIiUjjOoNCubc2ry1Y
i0Kw9AXymMLWmy/0ek/NeypAvw8/QXCSEdF3i3SSMcx7ESzhTquZ0R0OHwFnX8Mk
xRrTq5hP0Jss7UVOBGErQVJMhjtNj1B18R5Xt6EVQo8dNju7q0gCgkCkEmJM5WQV
aGZYe1sbLp5rMyzWH4uEpuUmsxHLnKTtN4+iE+LtFiV1UPfA8YLvjXoqIjZdgsRe
qyF/S0zIUuk8MivesPXB9e0ZzRNTCEO1vgqTzytsWTK7a5Rn7K0JBgiZGIHg6c3Y
MVQYbUV9aTkTfJ7ClgbsardKmEgdva5XXCSyjMI0yQtDZUiKBuMb5+oRfdoKQZpd
DbBl7sWkp1SvsymgUyHqbaZxsnv4zuzKbY6TIlMSyxlBEPOqPUDvFPPondCNixwC
yHYHQPV0LPc2olFVN1gLY8zp+VmFiERD/CxgJfOY1RwhC8HOJ7DgS7DRJpUZGc36
qXpvIVaSHEC9p1hVjkXboLAQNdvbRy4SrS3SNahbqtgPwRvUTUJKuyiGBeNcGA4y
qlNxgovvGbFqHp6ps8GnRRSsL51aKULzFCOU0an4jQhqZkzwdWqHGNAOjTNwc2PC
lRcfc7atG5KeDzHcAKxrZVA/0DCOndAZhLWZttzA8cjs1oXhK0YCXVRn4/8VFs0z
IsFTSJDRughVurphu0yQjXThL4rXctwAHiISkNRkPbo1BV7nmP8b4sEabXiBjdnD
2nLdExKme37Y3KkeYpVXEnhwT2gYDjT0byFOnNo2gPLFQqbd53Jk3a9oaqco67y1
llpXRyjPwvJv92wQZFQhT2KQqAziVqcsJQg1E4lfsSxNEYZ8F7qbHWKe0ihSdRYl
Hael4CYv03KvmS4LlA5vErwIEHSaC+0ihMC38CIdhkFSvPBREWktP8SgCnqOoQ6S
5WeThbMGiwohFwiGJHfb/CsIZSGOUyUi8pGn7/t3onoYLqdwPR+xol0Vzd3uwSJR
BzLACy7kxK3k+U62PPu2LkMP0fSPS1PwOMJtZd9aCBVkK5YLGFY7hyfkoH1Rcego
xDncWwys0WqRXYIZUZ1EF5oHxQdfo7g0BD45kYpbpI2gZ6dHKDkpE4NVSuOeuMaw
gyIQOoJ8oBC+JgPAmg2ibz7/SZUnDF2Ncnl4LW2lGdBX6oTrJivuz585R3TVwgZe
Om6On/ogxTmVfgpoe7h9W5RqmMwjRg7uF9julWfiVkfudyUeWNf7nPoEcRUwelYm
YTD+VZBx2nLGOQaoI1C1I1AtiYCw3X+NHrsC9GtyyW0XW4VEy3qa/IQbo30NX+9a
Nd1Cqa5hl7vYa2NiprMly3tbAreTN3i04Ku4+uTZPgl/dU1bL8SkF1OOERj6m1Bo
3S03L0ihVo+wiRYWeA4Px7iQ3ZyEw5goulwLbC4+mbOlI3XZLT5vKLHdKdkpXze9
3dbIicovcf6fZW+1iF6eCWZCgrcmDs7Xuky2VqVNoDD4cn0qzVtG9U5Nt0bbDu1+
AaClDjUwICd60ARbTC0AIQHUOERSf9moxHglS1kihQyEnVo+GStRk7QRmNxPkv0r
goRyXlJrS9K8IEDcLmSysbHbHV79QDmfWW23SJOz5q9Mm4uxC9ZBa6KzWG+K+eej
xffMedrYFFOmM57bRUc+jtxLr9lGnHeTmauRtzcmtvmzodabae7CAqCDOas5kxzk
yTPH8mZTFembaJF6Wbnc03o7KIvpBoJZu9ouCbnIyd8t0TiQbLMW/ojxahFnsnPb
IPKHHLEDwImcVmHhfrQC/GoRBm5w+CuzDbAYYJDMkJUGP1nrlN2vUHaXoncAAYUJ
FtS7jYMef3kvlqoN9kpwcHhm1E0chIjLcAzDxVAZ7XbQopVSS5e5ecEdGq97Bjrt
N0RC7yWWjMTAJQLUj6G4EAYalUp6IqLNVZRAhwgmHvDH2MVnW03HIk00bFLg9GF4
3s8xeyn73JRcHQFWq6IJhJCMoFwXOUqPAsn/IEP2LBUo7NO0ukBcz79nltaVhmBF
l2iQFkQCsp/Wkshh90fF7rMSCwqSWBGZDPnNZ31zfL5YLJGm4EfES0yxfs9aliaK
ac/qswyGIXQsDbCXZcK6SgonDr6++0Hb2Z/sIAdcmk7GHatZ7m1YDIdfalhQkXLZ
iZiELq23WweU09PqTjVUOVIeueuEQdy4+5HV+VS4K0q3lp5gJF+ETS5MzaTCn/hr
qK/UQByttboo9fSswTFIzGEt+LMOdVQFX46BdzyjOCjLSKCR15MrdVxqUHSTz0o6
+ZqZ2xfIo2JucHVjl/ZVdbhGdgEK5ZPuegnx7p40w9xQFi6eC7+LUO1wgbQ5M5Yf
pYFiXYpDD8HPMDgN+3LRqJlU8/y3G4TrV895lagbKpadtjZAV/fcZKHlC08PrZbn
W1m8SBvgOD4x1EqZPPOAygot2PdDrBv2yMcRN1bW6nzFNSEuMHFjeSXQHvFF5OpG
ZhEMFP5PS4UtKIlYnvurS1T6XDAlneWpcTWKiEOSwciRfFtkMm0xnRIBagxvXaAW
OVW1s2H/Z631Bg31BqVGitYkSDIy5dWXt4H3JuQ9YwkaHdI1OpCHRNNtPqrGrKCK
AN79wXQPoUSfAMY1vgK3u2efRQV/znTxr8q1aH8CJYTk+zDBQ3oBl9GmwgchU9Zb
/B8M0IF9Kzr6W8ktGxMqna3mpuM6sdHHXdspCk5ZxUTWiP26Ppw2Z2ITFckpB3gk
UdGfP8kRB6mzDP32doxg2Uym1a0oCGgdVaJgrZAso9LhHA8D5+a1st9EymloF8MH
QFVr9+VZPdpZKI7Q90rI7r+q/Me8KCdzmWm1nPnQs+FcQ9ueLSZ2IQ8UzPd6g4i/
UYcLhIBR68Oae5VYz5ix/rJ7ByPRkTyebDcxj/hfVjhANgy+uEkuhB9CPerMxYhA
upkFhUI05zOHCDfn3wIF3zMMBhQBkr4jH/GGTEaKMrFYwvAvz8xcKr9QeRayV6Ze
qYtDUZujAHyzYrECOlXg2vEUEKcF4l0i0DCPY5TTqWd0+aKaFwB8btk30Q8cHTYT
3wK2V8PvZQK6oEuOf8R4THm18b5UgDE2LtunJej+SfZvdHf7vdh0oZ/h8I3GBcUp
KrcS3RyjBId1zPfS8gVVPSPyFw+W+OEn0omshQ0VeI4w/J8M36a0p4vOuT4/1wOh
ArS/h06SSNmgqpqEojUmmebOq/jpLskfQXC1N4RI2NWqYsRQnBFzVk/8PHDm3pPq
CNDXyt+08wUdEXzAOe2zIuA8VXSCX06qilFAVkXkISJy5cDm5OJCDT12ImQBH8da
P+mdp+byxhuwyZo7KaEeFC9lMW6MOsAhXBux8lkUKANAuJ6AwaG7yckQ9S7H7WvK
3nelhnEnVbACezZJpB3td+m87j/i9PmjUKE/uL+foJZiBYRw7+7JkKKO4VjfktEt
bd/8dbGoIYRlhFx7d3wqSKxHc/FPyqIih+Hyow5u/28KdHqWOaT8f1z+OrvKXOIo
2/I4pv72cfaI8eR/dRQzVkH1hHrBU6SblsEQ2tFLafZoRPtWkaewoe5QlUQCYBLl
BX9E9DSQlZkftbSw1Zvtizyofzz/tl4J20RW8QgaY1KT4g89nEpNS4egLmREAAxD
fRFbEe1JLz04s45Kcz13dm0d3Wow28vMNznrm47fj0qEHXumazlyONfoinDihI/r
OdTZ3KB/JaiN2TeHh4tk8SzQJ4z1oM2I73aKH2X6IRnNYnayYGqvl0Bfw2mrH9ui
EFmCZU1mgx1d6YFUk8IwDJn4imNH0BSDQ/dOD/30PrtIOzDE+S77nf2q9K2zXjYR
fYXOWtZXjoDHskzKhezgck6oPmqRKTNQOlXtzYM2Unnq4wyvBcbmVlDie/R+S7E4
qURyvDSE1GY+CkPbI0cPyDgmxleFVVrde26SR/QnxAdyI0PXE2nXf9jh/jP7BEW6
hAgZqxBFU1nC9mOcdtOwL4Rxh0pxgWKg3LCPoXD/gJSQenJzx+jNENnNarT2SoKw
AVJsEUeapPNJc/ODNSVfEauzUaUkS2lDdA/spJgJfbvDjDSdNSZWJo3Wo+OKzZxp
CoOuI0+kO+9LkH85TD2JnfkVlxUvdzNNdhuuFXs4KHmaiAM2BziiS4+f4NUSFCDx
w0Ciw2D38Ds+GfK0lHmzH7g8ph7ljsSP1iQQyS27JOtYY0hXG9M++4vj0TFuOatr
DNP1ZtRlVSsCO3ZK8e9Ldb/bHgPkbX8T1LNSIvSSBQObrIzashFWq7zEn3Xiv8DB
kHdU1COwcCENmQ3u6V3E7dlqp1o9u8S9HB9ZabuD79/bIkk2nsJ7F8h8tLKz9e1Y
5RUyculnv1liCOp7VQxA2bUCamRbytsOUaI95ZM0shb7df4HVilWynmeIQu4L9OP
wDnQOg2Rq+Md/606GriksPHgc0GMY125RCgnP8gQ92nPz5xb4/+Lc1RDkLFRfWpb
G/25dWm/mKJXhiBMbDTFrmtFrdQQd+6dPQ6M3Z8sCLCNIl+zBroTNBw8s9THjrnG
OrN+MXQSr5bVMC2UcZ8p3jCEj/dRXEmkpHCWolu9zZrx2foH18juxkh1q67RCEcT
I1mAW5bXDqKMqf4weGD51qN032Re9DeAJAw3tIJoBelfHi4S1QYt6ZPk8qVofScM
TzO/UVMqVeyv7J+lYFhnir9PmcJ/D3FpXpamgjKpJglUmZC8wI7ICXvGG6VyW9ba
PTqMfKGuCdXJmFis7a1eR5Y1ld0puzwZURBjANraiGRDA5XPKSiczcUYNwYHBO4b
gSxUa60o1A1K6CcZyEznNjfFirYsBjQobs2hIufKn36CgUjC/Vv4z2Ec6rcJyVWV
KgkQ5K2MF7xXKMG8S3Yqp2rx4Pbc3Gu2slIofxiT8eUUsr4VWFOFqZwQDinr7nE3
ov0QAssnq14/HHgqfXGmfSSfQDvJNTAxnbuPyIwNFxa+wGf0LZdQm6qRbkL1nM57
IXczTPA+6SLL996MsmUztr55lqytfdiuX7+SaeLxK9iK99mXvdDFt85VHSlymL66
apjROEyDUnrqmkLbXzh+VlWNOEWdk+rg31BiXfG+orcpNf+4TC6ob1X14kRmqd4/
GBfeV1mWqW24HWL2LaSr4gAU+6j+7ISW0Q/CVPnuLkU+Id4GQ29kc3rg+YAZeYuQ
r1I76f0IO/z/QaF/u9PZo+KsPAq3VvUObn8O4lwGyGVVZNjRiuv1vZj1b/dWmTUb
ASdlFsQnVp0mal5TJHGCHcnk4CQdC56Pz7KlUUioz0EmiN6/R9TlAAcryjacemgv
zrW8lSIpwmQ589uo5HEsothKgV5Hv6BUKER3CIWhP1QZl3kWv9d84FQxCVvL3wyu
Ax+sE1B1MHtTzIwR8tMS6Cw9Ew4jz0ZCo5es1V7ktoFUhkTU559JXRQmeTDZv48p
2XLweJAaF3t1TDpvOHB8SVncUMbuWbNJTu9WCWFDeYfnqRAwY7deXcUuFw1QEivb
+0Ezl6waYfhVKvHPjhdE4JB3rkkQiHG51ArJ8HFBIH7YBuUo9qkpnoo0pVbdV6o7
hx+ii/GurEt1hCCH3aR9ebhc219xN03LK1lUwGQ6pmd/7fS8VrmtsIe6xV4X+AKV
OK2il15QA5FeVMHOKp66U7afUkgeGREBiQyTBr28cjV4RSkZ8gcg3hGB6wO6+03G
0g/Pa0gGgZCut8mY1Jv/H8ZExEbNjPMhXgKU3xZldNsOCsJflMZ2ERU5e/wWfOkZ
OfNC76NT/ZsaH64LChW1PgnWN5wy9loACiGBcJ9PasENycQd+e70+qzLl7tGTtyP
fZ7KhO62PB4Abx1WZpW3pMv1jw2HOtabkHHjm8hnre8ETuDISW084qdpFsP1iGqd
ZtanaX4tvEN4S6yHOcVUZAvAO3U1YhfhfsZoBZt1u4LcqSW4zcDGvSriMWpVRz08
Xed7swBasCdfdoX+c3uhQms41w+YmgLN3DWmd05dGojKyf9eKpXBPrdqahM2hh7s
rFFIJVMe3f+3YanzTAYG5x+v1We0TvVO2xf8h5Nhy+b96uWRZmsX2zxrtmHSnDwM
MDUsWitXQqzc3L4CoZyLOaA2i0ra7bk6xEHCVQaNz8o5NUFkg3CpgcGWI+E9lkJv
E3fARmCiUiOAYb2iQl5Udap04ZEwGrxy2CCfDV+u/OlcYVyrLzIBAdDMaF88FvQn
+MrwLrV/8tuYlLQ5GDacxCNyi5ngf1hGRBIw1Dq2Wi89ra0wHFFurL/0cWR4N2gm
RqjvtJqQbxR0vTcg7mv0W4nM7pU8v0fliWN5ekdk0f/MBQ9ViPAqqcOaS/Kju7LI
FmDcvzoAKt6Yy872NQ6lpp9/mt/yRC8FIXBt84af86I/Ros2Ou1XNoBnvHSIb27v
V3xBT/KB3YWrHfTsKCc8ESt74CCBRQ6++0R4C+GSo82mWMLJwsse8QzfWpJAsBGf
56d/xi2TAiEP6ANP89hQ5RXuVQsiurALXarqtI6ibTRLzJavCEdP8yNoHUK/2Szc
16kgJUKfkbunQsfrcZHRWiEdQ7E14K4Euy46M7NquIX1kQmREmeDBBScA4LXz7At
wZwvZfEx6dR9u+sEjM62Lz45qTeXhGrYQmhLECo+LEBjoruLWYkHtSQQXcOoIJLS
IMLG74GPZ2SDX9TG2bF27fpUrC7AbrHW/wOPDxtAYhny4EGBENFQuZP7S1RMOzja
voI6rxQk/1nV+eJEVVw1dqe5t/vTkmmZgLognbynj1K5/bfT/F31uPnE5ncec2Qb
L0ubdkeJ4d9jCmHAW/ekSXiGmNc9I/soHPzKX29CcFEW7UJzyqBcfHeAmVJ35yFY
3h634VZL5BAqp/MpDM+uEClNYZdZZDttz09l27SUT8SDuL8P0atfbtbE2UNGaY/N
IGZ+eu55/QYE7VxgJk89bquLFSgY1p+XGZxwiVGU97+BJykOo+PwOeR0oitPg59b
C26sygBU1FC9DITAyAwaSHtLRH1WCnie3Vs2nRHDRSNgEq4zDEDRg1xo10INcYHo
7+CiqtuSZUujEy0ZEDKdPqYlOB+W0se6eJV5EEcsJnOMfrreEDLszAOU2R33nIAT
A7/ShqD0dy/BqarZV6oCrEAt/dBZFcPeNhbaM5ixvBz1pNDlsOsjHtxaxdO2vsCc
7vbTL3JOGhocuczyLKVusyXeUDA1Wh0W7MxzCQlNNbMfL2/+2j1pyA7Dl0/FnyEO
QrijHH0Sn1zKlO6DTfclwMvj3za8mtILlxSBlyy+/fYBc836zgCXnfthc3pOsz8l
kfVcaTi5yObJ6nmIXOqsooIGybV+Ndm8tzC1dgoxGIHsaJdMEgSdBUXhzQV3CuOw
MD+dkJIhzj3xn5aBpPB2BytieNZaJyH+yOxhZ0dbuE686ZeGL/ppuMxAYq3XRCoJ
XXlNsV8eWlUfJD/wQSJp4JF34HtitGHGNlGN/HJ6G5p1oRD/S7HkrFOPsxzLFDQ4
h2S9uMYjrmqfj5t0l9+zDNU9rF/xk/jsEY53BfAoh99ztPjj+vpltxuOCjKbDhAR
PIeJOYm0hqAULu6s/u78L7UzDjyP4z5FPzMqeXrOLQo4W3yqNyPHcNdEdmt/9kXG
+u2Zmn0rlgz+fMrIJGaJtVNQ1hFyErERtak7jbWEAGPEVo7891dVwnqrBNHGRwPu
8MMGMHohKV3dYFmFk3XTN56wdgRd2K8Lgq1ctF0Fsq3emsechbqcFzRPhjZMBXUl
U588zZd87D+geO0KuReBgKNTwdZXoSbFqyrORG1amXTFKtIa2PCv4ZuGla12iKY1
+uDaJgWXnHNbEsvFsYx6tT+jfnRRhxJtZPwMVJJI8ujvqZVZY/j2+VYvdTQb6k8S
3HnrX0qpsHg6Tyumd/DWT9DTz5sPlRE/D7Gs3nvS9O3K7NYOFvSta7IRiisVAmzA
15hQYbwPsPwOfEFhxJlct7dt2EpOaCX4GhxWoWU93JAQeA11v/K0+bb/kELYPVxQ
S2YlkZ7ewHcxRDDxUue1JhxlH4ZOvuKoLWbLOaaAfseqDoYM8Hvyfu++8A82XDpn
jYRCdFi4sErcb7Zn4Jfyo9wOeRgYmS/E6ibsk3QSuG1oW4eO6vYCboFDfI4wfF8K
f44HCZAAfS23nX/OPqQ3aIZVHbenG6qVMVNZbr8DqPrjl7oolYK5bz4TiTBJApAN
pXtc20D5vbY1vlTG6z9MpNOuzFBCW1uupcRzoHwsvPgPj4cN6FeJsgWRsrY/Firo
tTk724ExkYfYWYwqyY/42rh4lFxV5NgWWMQ7Sf1twUSJbxKVrtf0Lg74TObgJ0U6
yh6s+erdWJ35VkmU09PuKAsOXTBjd32ffOIPOcrUYA7BUUcrDj9ZFmdNr0eobTKG
s/4WGPl4vDhhQ5uV8yaVTh08J4plDgwFKop7OIAX2Lu8opEMRVxkJ/BTBC47ZSSR
9UsSG4J3RvzhYteD+3bDUeeuOLDT95zE3reyDoO4nA6cWp/gXWhuGvo+JgVV1amI
yqeDF2ZMM7g8i4wM2QPxBODECa2jJUhnNmdbfFUf/tk1LOzkiIwoXz/rGHjPryOh
YWwibOzg4VSN69pMoDJPewKca4GpAAvP+YyPpRvqP1pXIAO20aXwDvWMVelhbYeq
Y4mtEHNEQfRG3ip0cro4qcCmgQNeiDZ0K5tlwKoLKlWgxY+gfMOxr60Ne8gYRcH4
Ofa18vCfzxbAu+8TuSQx3huEbM/WSTXzlHBuKuzrg0zp/VUj+wGgkxI0a1QFEAGQ
lCVXzvl0cppOIc37LYFNO7dVNqf5s2RKlCefO7O1KUw51+ZHmXIGsdwG0hk1P27n
OGO91NCmTqeBxkryKbmTITRSVJ8xYubDVereuKxkTece/hW40MPHO+DOD1uEyTiH
fAUdKyl631ya/Zy2/UbuAVkawekactZRpJXqcBK4pCt09yodOfnLrcnRimyHJ9r8
6uQlhbbWjbrDZxN1OO7bVASexl1LoB1lQlWATCCH2LuukueMIDKi5NJ6BBVJKoTW
nMiLLnic2Ujt/kL7BIA61CuTfzwST5h2RW5649ilvTiE0RRozrSjJ9F0eQZHwiKE
ky8ER5OL+u7zC2Vjlh27rb4UiMWppvd5z18CczI1tZEAdkUvVcw/SF0KK7gwtsaI
pzie9VzzkHr4hkZ/S9ZZp7j3VsYbGXWDu32zOWFb3IQeObUMlJut5LhULEcGTgbY
/BMKTXBWpTI63CaFW4cz9snsW2Oqhv2fcpTmJ8dEf/ssqJsqdxFohGQKTmdsnwlj
UCyBQJ1wTVHYtNG4tsuw5CfFAW9uarEaXjAXge3J16PPyw07z2dQirCFMYpUtHJp
Y+d6e3oKQJ3LpufjwMOFl58mkFFQseoub4q2fmMQl7KKYky7Zp8yrdw3J+fg5jTH
Xe1KBewYcJuwjXKXJQy1ZoXOJninj8NVUUa5utKBu8rwuO22bJkiVqGIMJ7Ph/3s
rO81KFnhxEWffdoQlMG7BEMrdtehzBcMm4ICX8Lj3OGXdmWX8hWkPOUBkaf+HL+Z
qzXzmKWdwu6a+hIsz1ry0L46iXiw7YAh/r0lEH74ZulhQU2tBgZxRB/Mai9jeSAj
C3TadaZ5lEjUu7qlYSuc89pIjvERz+waIJOvQmclWp4fFG9e1jXpZYT4Q094KBOU
8TqBP4SZ6whASHjQhjM+g0n/4GKs8oXP4qKVEcLexiM0u+GoTqkJzfzlP6CF1jDf
uVS3+vGBQv5rJcy9E5D5/Norj3mTyOdquzWp3DLU6aQSstby4xa/nnbPLpiNwSYi
3Ht+DYBe5h0VtDJMLOxSOex0nuugTP2mjPepLFKlybxck4uv36KoT2V9aGW92ViC
NfZXOdF/mkk9Fa7yLh12ilaL806nbaePi0ctz8ou7+FthfSmaReJP7V6hyyfPZM4
5uLJKqfi38mwrJVbfaCCr5OPJYBh6vMv9l4S6bDkQsslTgCNZWO/mP1u0ZAtbtLl
Hgjawcc5eABiXFMx96wNBpISDlnuLqg87QIR3nSBK/keGiTL2EXs4ocNUaY6DUm2
yuHxkOS60V8fUZ8KyFaondNHbIl2u3wQ0wRoxT5Cn6zIlN2FERFtbbZeryUTnGd3
+vL1GdbG9dO8mLLGeRcK9TzaO7U7YyJPt/3eHH87LUV8ClgMCDZc4tOrO04JGm1A
PxeteNZJCRtE1WeEvySWJgkdddsnvR3YIt9Y/AH4+swbNVjPpe0qQBojaLrozl1w
RO803q/yEQH3wOS4oZD39g5zhX+SWqkoaAWJAF3Ic3A1Z44bOJVfxVtuQZaQdziT
Q4xOD+9VlMUcEpA3gnokpUKg3Jnv3FhFAH44irV+7DpEmw6LXoe8fVoF8ITKEAul
Vl16F81n6D65XFP04+xSiLPV+nsIbBxtHAI1pzZtsS6j72CwSbbaa5BCBlDdPu/T
ddvVz1JZUL3VgdZR3jJYjpFuz3R9slWahoXCudsLNIwdfOfx7EzTjhCy1vcNjMAY
i7fIbZr6zxj9y1JJZ/PbGaH4X+j9Lft5RiAgI/blcr6ywYUoizy4K2s0VTLBU0g1
w9fXkNjmUsGAMsksqaimwst60IPHDIPXEHO7OaiVxGr9tNHLfPG+oK+7pQBQYBYJ
KOUIyr1wD0lBOiDdCKjRq3NLD3XqGWAcnN8DLsuPoRaGseYAeOa40+AK752/UbwV
yy431Ag2Gmp616YWhsCBQOjkmt+BpafjJMJ9FcqXbndOFqMu41wKO7PE/5oyKcLk
BzNGSrqwqDgEtnk9ABoH5qMoB2izRnyjdVF28EXx9C52sLhFBkv25BFv3VIlhnB4
jeC07TgwPnJC6dibN7e/6EE9G6WMerHGoh6/5/LhhEORKStbcjs0rNWeh93DbyiJ
MuIyCgtLCPiEN6Vfw2sjrxVrqSoC2PdQer1VuMb8J+zxMa7iIZyD3ibCQkaEJzsw
hVK3Aev7TZXwufzYD8ktRXjv2hNgthMF0hLGnVyBwVYfT4qntdm3g1dclaHYA9BW
QRAZ8nY34r7nbnBnUpJorfwAFbmtNFN8AalLVDd+akXRxKSzZXZvSdXUc09HEBTS
u5vVstokyhNODVyyY7VJo5YRHFPnHssGxDQIS4QXgbX5045JQ/Cs3bhs4zkMhyGc
2isD06DlhjHS1+/deTq+NCvXf6jhPFSUZzE1P96aJltDP3JTeLmhV+2PEhgNJEe3
420+4xwrIIb8taDxb0Vr46cIyswjJ6Cvda2pBQgXX0qBQYpM58cqLgB2Y4I73pTf
Um6z+ybJ2xjenpAi2sius4Uyqf65lrQg+WwTrpPFxmB2u9NgL5pmUx7AphE+3ckS
aJht2o6DJZmppVA4fxv848KnfBlumaOkwVg0aM8RREGmVQQceF5kt5b/lM9PZlYc
aaUGIgQeoOOm7WRHOpZywwSOB2HkG6MwUHo35zDg/sw26h7q+PH0fju9mX3ztt/l
pIcZLg3bGene6EVLJuE21kuXaYOn7n066AFSE+RX3r9LOzVACAqROcKoidAmrIHz
fI6dZNIlqsLdMEEmU07PGCovm+MHCDfbweBGOnjDUKjtjxDqCQFyjkt505RAqzcv
qxuBuedUbNe2xQHDuLCu1JyDorY/LmvtyLC78qU0VrKI3jsqpsi9By7Ulq7C8HPy
xX2odYQYgSzBQcQiypGmy51VUapOosPB38A4m1i03KsZcChc/BO/uC0VQ+c7PwhH
v7ysJ5AkbpZFOJO2O4lC8jQNZcZtnFWWIORo/sY54C9yfLa/+Oos5z1WTHm4/AnC
CzET5BMUIjefNdITnuDJ+bpJq8UOLe238KoCcovZxEZvkTT5ejMs4xXCHsWMZ+8i
S17DCfitUd3X+2HD5zVMBOy9XmjHC6bY37d19cwJuIkMjW2PpnbwWxBvhCmEDN07
zIf1OV3XI0JsJeS2poctnlyl7aopjKG+K2YBm1DnQ28+SU1y5N6pmbX7wm1YYUBE
R5Sp6HDvdx61xfS5iieKMhVP3cqolerkS7XY7tL5fQELKAWdUQo/f5s8T8s1cNgx
gnZzugUlKQpEpiLsGlLM97Ynj1Q6+o8H27uRuZxcpmtArAnVmihlwHya6oVAITci
ON1Dl7iS/Ct2Dadp+CHGyDyXU8RD8PgDaFneO9ZJ3/cOAbZ75dXiWFJo0paM+LlZ
f5ecpU1nQxGmMNSi2+uJrH2hnopTfH9uddBglpqhuJdtDVRdJmT761gkE6y6uYX/
zMQ+qAtqdu2/8KLvEDU5/ASN5zKZPs4cdHjaGtXvbhtIL6EKzuU6Nl6IxUM7jCdx
nP2WlHwP1SnvC2Tx53xWwzhK2z1tsT2l1f2fuTjf5qxmk1cS5X3mSsHDi9StVVf7
QvDQMRs3NebhkfKWIhgvHVCKgJsuBoRnGnsMdwuUobBImaPgzxeC+/XHU7bKx9zM
q7I7nrrbLJ1N5ng3eGZCQdgnvwk5Qx+qIwWEK9O1C9rw5j3XjS75nXzy80axTGis
U6BbXe+1jsBaqzWLDBSmXNClaqw+YRIZVpVzGM968a4SjfJ3t9yAwwZlSkGgfh4Y
O+XDmVnghpZTlkBo3HOGmb5NVfW3peshzWM/FQlkYke6DlZLyguEH4Pg/7oHORfB
kTsK51P0fYimfsua1binI0JhXLRXwqE/anJwmmnJAcOS5HILA/BZH0giH41r1Tao
zRPRdFrNqDeUI9kGYuKzyZXrAtXDzFFuIIYreTsEhYo/0q4kZkr05AhAgCZv05bx
H4DjB2SqexKzdR5qLTzS+a+lqmZQw8kmY0iR0U4xKFIOH02tbxG4X6+ZDRLn8pjP
PzfBxwCBnvcirNa/wGFAfvEON04IGOBgn5LBKHPe+RddHhVHn+RhClbZLsGFUTwd
R2C1wmxswFB/MXXi93e7euyan1ftnegE5eBJDbA4Nx/3xp5gNY2BnJ0UPYKX8H31
OPGUsnlKHIsOVlVYwquau0a/QrVb+7kVSin44iUpFCfEE0SPRjqDm+y+9/IHTmVE
yLKv91PTT1uNcwLHhRQEU4QwAvJblMyeosWDuUwrmwIMJK9rgLW91HAH5biivood
YzhH2avEZQukw/R9qpORXsZd2UdxYo9SpQ34gXizV0m2ecSNe3uaoa+3lkO1aahy
VRp9hMPrrvwUFf+VPfq0DK3Ov94bq5hEi3O4ss4GnS56vpyXXox2nLNGoX1wEddv
t8KvoMdLRKmb8jZWWv3v+yCV3hJbgmfXnZM4HBSOUj+PhI904JkSWlITWQ5Ilo+K
W6ybGggxq2MSdsFVHDbB2E+ahayI2eY7D26z7bfA07o8jDyt2ZmpDHdTCCjt3Nnm
x+9eJr011HBdghXdL6vSkRiBHsWxtHhD6CNPSibozgqru9hyGVXqB3HpCIwOUXKG
iAkAAk+Ka0k1Aii+6tqd2UGUxQaBrdvMG9Tim/mv/DgsYyH4WhwBO0Kn+z9oP0jj
kfZMM0xemFZZyySisuML8Hu/24RRyUho5uagQeT+hWWDJJOZYnKAjpZLKtM88tpn
/YNWeZj5OOWJ+uJ0DreFbCUy3B17BEX4kAVE88rTa4zzqqIBZVE6naDP4iYXV7Ze
AdJtymHowqtfo4Qpibk1WCAyEqH9nn4rMlQOkocUAbVfON+T4qoweMV1sdMISIML
h1lrvvceT/HJz7bQxSeo+dS9MFsHOY2k5Qq+Qsb1+U7QckB6oiFASVAFRtLUCdpw
JD2yvkw8HtKe38svQYkk1Rr2whlVNXy5C+pTIg3H15nMUh7DR/9GohBAIjuR4w0M
zdEmMeDRzFnNEgcPsogYBMmUgDK2zodC3oE+3wVR4vvFkM4toDGTbuKRfwWuGZBa
P83WQ5LxQ2GYCBiScGjwc6oNZGzPpaLzc+kPHjfe2h6nMv28D4e/sCkfiK43k59d
7mfDiKCMZFMLaNqj1dBxnIQSKX22W2g0sCnTYA2478mTW8NxdQp+s+onVxhkxdfc
wvuYklxtpOeDNz5IwWZXDZEixXUgbkDCCWtxraWmxq4jdOaAGGg3/PI2cr0rMPiv
hxdFAtIKmuV5z4IXGA5vd9QYpsGhG1CARVZ3R7Hrny6J0SacvWDTVqroXSWZ1gBv
g9tdlrH7lkQ28MYacCacuAM42k4Vb54I8FDsYUFGyrQWrYkemGNFKnvnmSEmEWOE
tqNB7LXfApxe5NThIbz1/A+GYlXwM42fG/QJEC5M0WLyGjYB5rgji8zZ4IlOyZEY
zE7vpFuvfAkk10WNSMbOYz58PBjk8pViNVOHO5L2lM0vQnrNhoYsus/qbI6yQN9x
0SVYOo5dasI/L6WaW7IugfKIm2/Rn/L/gFbKB4AXKp/rjwnwEFTKSOEh01QEvmzX
7lFSpBxXyx5X8Ec2QJ9x+qlNE6mFEGoptLtWpfXGF9w0EduYFYrA4LziM6dgiYTy
CsKrDyRwR+89Dc9+Yq3s2MA3d7+n4msGpTCRnOFmPWXGw6dqbcuJMV+tcBDaQZFy
DrGZ8uTRJl+1nI4hD6TQBgcXaIYRKJVxdSQiCXAyLIIMFBdGoevXyEPHDk5BK6dA
lmlvX1AmjLLiDmOZQSostAAyuSzw/SjWI0EfdP0B9M6eljiu2X4FBZsF0m6NNZhG
DK02F+dogU5jxb+zbgKAb685jIJXriMRwMyhoD0mDI0OampDJQoWks6Gbd4aHUfw
5hXNNuqg5OYTOFkrooLfsk1xltRB61l2iGCA23bcqHQnbGJE/zF70Kowm3MOW4+5
+dhTSO/IsAGKjrSe94obO7y4xotzc0hVDxvr+H/wY9gZDHjPVkjfeBPX/cpwj6SW
7nylEnUPgBPanPM3WMXG7fFUIgsDC6uRduwC6T/rtzBCURqQvCZd7sh+ddsP/ur+
T2Ni8M7aM9teibA1LBQVqKjAepMb91YWP1nCxFdfQJY58+wuBYH1pea+n+6V033N
TZJl4f+p2Nk/dOvQRIHdndfTEy5hiJ/DNc5s3LYF7WVJKvSMQH56phKsjaWDC2tS
TcP3lPgMK+P5grIPcZoNZrSUCjTJdm9XIxl/5AHNNnVoSuAcsUYlsn7fX2epdLFv
zYVcxqQ37da3HNHADptk3I1Y6z4hvoF4F495Bu81PBxrpMgM8Sc3sYDEkHZqYEO+
s4fNmwHd/BuDyVNKBY0bnpS9JYEAc6J3mpCFw9b/QWOIWySVSmPHXiPT0I1W0ADa
33sY8mPyL6YI3i/gJFhgpIER+0nov52lo2009BDxSHqypxBD0nQ1966qriqEiUkk
rAWQAspAJXaQcWGp0JcQazMHu24wfyk1aIZtHsZTa8YPAlsNXFB4oH70Kkb6K+sC
AFwxNTVlWcta7oGPwOxphxjcvDWY2gND14qtlbcTfgGAyQl+6xRb93S2qtTy2Ro9
2QpmRfJGDYXxiaHgjiVa7rVC6ZALHzGYeVvU8+GWl/ufH/q1xAdcSVjqmBiXBlKq
h/hHrAufcTuz3640nzQQekiu85lxKdpQ81XJd4fHC5w7ywjDp9Xi/68LWlwaL35q
pvp4tOSZZMgK8KISBKcctZ9g2H8aKrm8vc1n0hjxEMOBxIIFnuNbyCRh4AI6CC+7
d7aSMeYwSadPyfbHhupph/R4Y8Euty4hAgNfy6TA2rNJaBdA7gLq1O3OcEf44mY2
lNM2vA5aoWYbB0CJ3ymcPL5Dc1xGSyt/PTplZItBB3zdH87mC+olmXswtI/NPlZ1
+mlJN1IzW3vtXoSWDwShrEQQViuaqLCp0Mnz19sJDns45qmn9ZiZbT62pxpPAf5N
6H3ZFHjEvQtUqcvOHaXj5RgzmjqwV142ZbcFDMWPSEreeuL57pADDC/freUymV3Z
eauiZkyUX83+ocFLQlKYUsvTXAUpW2D+jGeG1IzCzP64kL/HO8RRGzCNaS433SWR
uo77D8dOjJPMgjRFe4q2lBizfBbxuwbMAcec6QklWG9Lobshd6mO0Zcg5Cn3bc7c
UGegj/KbE1qZFJyeZhBUsffWKbcn4UZsh75zhKx+Q6DE+KwxfOmClfKr+26+AELE
L0DKxInjF8RAkbl8T+8AxPEXCZZ1Twcdkc1Enolbn1Ps+LS/j3prUPdrUjOVTLSM
w3h7F91xhGbXbaljaYpuiL25DeBHfqcoeMTl9TuPg+OrQ/VdiiGJodqOGUNh2t7V
UjdA5CF4zfCQv4FlgBFkDSoJqw1F2F4oAQCMnTL3v8pLvLBK1pPYg0SY/6pTo9dV
ze4XUwdivDPZgpIZBmhsjAoYuNPJue6QnCZcVtntZAEpQMRiW/u2fxiF9QLnYWbN
0yyyOxdNBJQpgXZV4vs2xfp/GJUAPOKPDPHVLOL0T3unIhCCRhdFkGtR7HXJ2Po+
c55sgmD6wNwo4BCvyJ21oYBPJ94or6Ie0Lgb+U/d5SFIaFHWu9mpAfJ6DCyllvTd
p4/5ukJ4ROoOOVQdu+N5WjXVhyOu/4zpIYVwshpa7R0Gs3MQwk5xyDtmui2nizQ7
/sTbqt/sTBUt+24deh+Rv02I25lIyv0YS+o+mLt41DeJTzQrWT7TfOOIBeJCCYZN
6NzByFstNsRhyPvFg+rhPiWQF3PRanLn6MX/tfHdHc1a1rS1Y1QtoANgRotXDEDG
SNXux7jjUvm557f+2DiYHWZUJfZy0vkL4WCzl04d9Jhsnu4Mduym26AsIWMky2DO
jG7sFafnKPm7Ta6zjQYsvZhmHbig4X+NLEueq5/I4znN9pANNDbSNXP5hQO7RlhY
lkmBxuPtoIVzs6VxVPalk1TuHrEscDWUwRsNIKN8i4Q/t3tD+Q9cNzA4e6I/L7ZP
AXJGth4bsuglvtPWETcE1TXhWqfK6cxfdyoi7xnc2GbjTzvpGngmlNuRF+jyyWrD
LawuScbFNVyBTF/W+pwAfGK489HmW60PQoiNfZf0pIbbRcug67Fd6L4q51hbnxbc
CnGfMlDMGF/chRqBFdPAbjh5e/5wEZ8eqlB6luvz/dWMPDHSUJk8Q0YY9CTsXPKU
2Xk3VlNFOv0Wa50AruphFE+TBDha4VQwkYvVrMNo98ky5dSRZKxcywDYdJPwGMI/
6k6nMfj6vS0tr/yr9PSNi/lO8gU1NlxdKZOfzTGusUt6PUENO5WdfanuGHGG74Ve
taISbmSNymByGYAmBvHC7aOLmtqND6UaPQzJEQ4csXGP8w2RsIsg83IESVxmjVE/
/aKkpzD1g9j90KNC8oFmPqR6qq3RItbE0auYuPlrwVDcSNTYMmi3NjSR8WpvzBAg
+6Cr+YmWToidEjAb64Fw3QlTzdOCvvmufM4N+TuM9kuBm+UV5+xIQEidlQuRwl38
83SzUGg5k2tdsRDknGSZwXSmFH2WuDpSoaAsCuHseVYD3VCsBelYE6+MkZQh16A4
fBmR4RqHnKRhYP0hHnuROH9KKoygFcA6MpRm7rgNg2QGsM4CnILeW2xt4vsU7DhV
fwDLr/fg1CtKkJClxDmaw0KhzNmhZUCnRfPEmrshkFaQU6RSMlveaPtAs2MkH+uU
wpEneiM7UXx908u82LW9sVthF8jaQ3Ioj7QmO2K2jxOYaRQ0mt3AlCN0CzcuoDRO
pX7vmej9zvWzfueKCX9ArTUpgxnw80X40TDVTW6sZsoRmUTqrc2xoBkBgXIqE4Xg
SHdh/ck/x0i/qGrIbqQrzIq0bGmFPUrZW1c6TXz7fIx/ho0FOu8MfjIDFaq+u7oK
5xri7YeMbYG6Lwdk217ihBAtps8pdyVHlYIEI3OuZYA7+R1XiZTDSX4as9FRa8iM
/6tKQKOtk6fJpbMf13E3v+fVdPuyfd9rTWS9c0ydV+NIm90oKafeu4QDvYgKfAdp
7ujyb9k/9nVH1E2PR69v3PxwBD+VCbepGr17XEpivBYp4HSCtQtpKuauSsGdqnND
rC0yq1S+gRjia6II4CZ9IMSmHrRR6IdEKD58cvG1ynv08PmBzS44smGM83vuDLGV
/nMNlRTmF8eKR2+mFDIvUrSLZ4pugZapI5srNUpcm9tb/2utft3c5Z4RhVCtCejm
43HXY9WLcOcWcFmdAjK7m6/HzciFBFMCoRX518QUrqzF+t8+9iJoNOTH/NjfUJOQ
vTJdxb9pJ/5y8yhy1l94lya2dnK4j+j5QGfSW3XsWIXAK+znfUXJS0Rg0LsUu/8c
jp7EzPObzMf151AY9bkds9nl/H36Z2ITRLBlJBSIaVKQV4Gd7KAfIwYExVzq5VDq
kNeK+bId1D01WBDYSmdO+vge5cRCR7l0xcsSJFhvwu7EZ9+BdLsgGQNi8JtsG03b
cHZ7/BaDPjV7b1Xtfs0v5Gtx4Zi3bZjlDRCCiPZZOv+ekB82ZlhO+6n8WeahpkdB
qDMpgb7RGDPeVZpGAt0YjgncnMUBdYi7kqbFoaqXMt1kDbq++jyrrFg2nQb77sHr
zpH0yf1BzWCVsjXgoa2TpkenK3q1ko8xVIexpUXh0nryKri74nxN+3u3YHEEAYSv
KUQk2dOgY7lwdkoLbcJwQq8YkQOPYpOKo5n3gT+VZDvZmxq/AwDI0jG3cQY2SiO8
7uaKMO0qcaqZ4pWgZpWVWjCgznNMFqKFN3cBUs8AstE8YvJmW9r0upBbT3iESMnn
yrEOpnwgIWFngHPqxx9b9J9AOGporOVV7OXTgy+Vpr167w+iEaCDdeWKjHceHhJm
bHLl8Xb4Vn2pcw5Mci4oHe6Fkibi05bZrKzU+AuVjbYuS5FkduP2gxS3f19iivdr
srv45+8Vjsw2c36GgqKeGr4XnDiTQiXBF/nWQpbjQibMP0OIysPAvCHRImZ5U3HX
BPgxBj1Xm+gd+Rosgr9hL9tw7qc7bkYiQVXTG9V3daxwRUFXFayv4pSH3yi8tDfz
WmNc0iMwJU36WMgSXFtD5EsSFL565SKA+fRBbWdqVu6LQ3nMtIwSJgEQFzh2ufqa
YVVHXDIz9jOjKA4IXFasVAOk7ShFC2a21u7vdJMWuYBB6bSElyZPzxfGt++YGb8w
dSKToAa7i1y5hgFev6L+WRdfiXoh/smU3rL8zQrK3WFx8KfR6zNpzKd6SppGxzfg
GwH5AfEu7brZeG/PgbJ4QvZSPCcGVyBvJ/0IQLXeLAOkL3w+YsO+kGFido9ikLOV
TbMZpEy1QGO/Oj4sMuRu/oc+FqpnpsbylKVLDkMExW8YTpHpGauKrG9/q79rga/n
0tN14SE0x/PpDVZgkr6czk9zejddMEqYKxWF7AeisnWf9J9plaHhgq4gy2HcsEdU
3ltv6MxmTkXOD8OeFLN01QPxIrB6KXimybqkp3M+J5jrAJ/IB5uobw60GIaDWJ+Y
Yl4zc8RCasKh1WBFNRSXN33k0+oBEwsOPIDtiI2y0OGal4CRRJjeti4xxreWiUgK
WxdlxNJd63pl65nWN27ZO6/H/VVvdy48XrCMdJ3rK9wrtwfAGFe0+ofrttYmLdPo
S9W8Z1/aDkKoCtTe+RUIj9bfRa99pDDUh5Wsk0mI1me2hThacaBm5eZdLYTND4af
RcmQ0PIUGAWGxdUlDRvh1+QZjiTRmbdWvPBNlanJCNwEW+UFvDGGap5i7tAxLTh3
NxCjZOi7e6BpD2a9gBVM1M0pduv8SpbggJd09XNGstL4Kan8h9qTPan/fhbbCEPs
C2lICSyE2Sk2PY4Kp4bKwDBa7qriFqN61Iyw3kTeD8voMtNo/1isfAYSJTMT0Rix
hhzU2at4EmMmmqX8EgFw419zlI19UrOymlocgJy52mGfz31aO0m5F12qZyd1hB2L
d4HYDSiVRgm1fzNDNVRWLkamvfKIrdFozuf4N58PYSWabA5E5thbiffwNTFc1UFD
Pu7hiTXKoLb815Cvrx11K9n4gerarbo3tiSBMS6GQnwjDamKRoo6NG5x4Qk9fxQU
vyUF+ftP0e9VoyxTStp363qeMs93PVtrWSn99N7jjNYsHHrxB3idb16n+ckXDeRD
poyAtT61NsH1LWS1X/3LnCXqtGXJBhmZjkeix/RkHY7aYD3jrF8yjoiEL01Br2h9
0/VFNF5O4DykXqZ0PhbfXqCSdCtsfYft08EEggMFk6/HxpTIL6sG6GJO7rAFy09D
ZqLOeDZ3w9IJEtmls9zP+EV1d8PW8jm1XV9DctNXbB1dil+Huqi0o4r2C8GBqsfS
C5YXXCCadlkQHxZIubhAUp9ldoa8ZVFgerxl9YuZzJ2Xwsg4DSA7Lys0jERJ4cXL
j2Ut7MWGzGC2smPXZpVM0u9WkkOIh7N8/UgN2xc79Ho0CeuedFhfUymr1/N/KW3M
uVH6+LjGpXCIOSYS4XATwAwXesyQo+7svAFMCWLbfFEcEYFPUXBYfFeLkLLwrVhE
m/v5soqcD/s0aj5IEX6b07g+3ESSL3+oHvsl81fuAAMb85zRE5wRYk/RSIswCgFX
LlScBkj+7hY1gye+1gQdBRHnlJKMZ9vjYuLxRhsZIgimY275n4SJK9dIcncfXlKe
MuvHijL0idieuqDWj2N00RKjWnSMIY1iwmS72665NMmDwlWcPf4ZUxSJ2mHxtGdf
tINpRCXf3sBK3pLW6IstOWOflZKrIxWsjOQsDSymWIn86Ul/undoQIBFdmspV0Tb
uaXjwZveqdhVk1oFsPx5N/ZDUCTv0P+X75cjNHlPwf8mbCSldj3i7+xPhbcZUDUT
4LS3BsejjrwgilNjdlGU14bXY+KEq9Bh+1kaxA7cll6yMwA2JbRlbCOA7KvqOAwo
mCnc2+m1zoKZlttmM9kscvJtYyVMA3+wpSYb5Lzj9p+ONNvDClEsRy1V0fLpSqRb
KnMXHqoYmx4SeqU+wlFmy51HfztsWuxMK9SHatUzd68RZ4oIEX/gdc69PfyyXeEq
hl+9RCqQUhD3DqAndrUGWZSoEoj6/4UWDCxvy+U/XxlD2VKjQ4jvt3zd33ZklDxK
cCiRfr2JL/94RYahlR2maBHPsw9l4/UbgoFdZtNllQyPUJBodRCe0yGUxfnC/tm/
U/n0GeXb1wN5d68C1qTM3VDg+xsyyoAz5a2QC44reAipBRu9LctvjItdYM705WKS
fioKoBBK7YGYNGbj2F9bSyCS1rBabq8A93TKA7D8lGoLd5A+kWF7bGjBKuPCq2lK
uZS7w7Xv/FK4H5eDU6yGeBSF0o0+tKGaRpmyKOAjz8U0EICBIO3PAEjXXtxGeI2m
XiDjX/DShOb09IjVcl8BfrhveXbVXKZ8Bx5CTkbQUqg9uJ81m3n3BqGPmRR4Pimy
aofjfFypx8al+wsv8j+wzs6/1F0/Ljuhhjpo5Vjo1RyIMckLebXNUBKpXwGLXoeF
X0pTwc4m+wp+nMxg8Bv3AYeC2vuAyf39Tr4l2+1yIuFpHSTJq42yT3f8/GTOfK/R
i6SWpNFGpLpXs7Sy0a1GnQHc+Z4JrfUclJrcJRIMyHLzLZJJBcdROaQGVdwz6orC
dxRgGzf4laRiWAPE706eVttgvCo6FXVjyZ7+VXeDpliXUi4Q3rmzVijTT9PmQTIn
Wqh/1hRIEFAxeSlUsJchYSDX4pr+yoVI5HyWb0wyZgLh9h0YqB0WdG71zBdDr3bB
BJGeRfTEzUujRr58mNg+0ZnmPkCDKnufSn6lLRwx0SP0tRKZIsDk4/9Eu6b+g6RP
SmBMPIWAc03EZvpqVdNVjg/FM9OW1Z4IDFmKqu5LdMFc7+o7uYvaPhFnbD61nSNY
xyaJ6znkgrM5uuUU3/IkM5PwxgrL87iy8oNBYftsFoa4KagrMEkKLj1mAXpR5tGc
CZIG0CFwmoBVOknJnE91nDHnuM+kcryIS9avFbmIfxcrsRipaHqRznoHVsUwYqgy
gSETevTtRmStHCWuCEV/pQsyMoiXBYA1PRZ0EFpqcRi005dZjL5zt65uRs8vhFza
LvzpLXTfr3L5tfCCaS//YACt7YuP+SxIZT6t2Kv2PtHVLm14124yomEKFCfYUh9p
VQa5I0vti5F7/XgHXE5vSA77Bsbn0r09bPAH0RiK3GKGUe3M8BFNtOtzGNWF8/+q
c0lrxPnS8P+yT2AZdroyGgR9coj8Pk3W3Qpig7JiaCbIXUx1Z2HVmQCmAusMhJg5
yh2ykdj/zF9GUYmanZX0Oa6OVewuZFdOm37TwC1ea4R6JsT5HrjgfxH3xL7hBEVO
R23+SyGRZWYtMHfET0ApI6X4brhVh99zOzOmuordV1IGul79MKkXZ2MtPiPq7vY2
4iGB3hz9lYuMA6JH/69gBYaw3hXOW1sqzGcTLfvh/1b0npSUz+w83Jt7FWUXWfPD
9BK8BzRn4rQ3g4mTT3ieN9uCFy6KxFn17xh0Uc8Ts3n2hwlqzyLMNQMG+2dHDqOr
kELMKzCyHTUmSyVBKLKM4+naTKkiLYMMU/O3bL/bJlOIJqVAGvrQvX7PVSHzG5Ok
7Ziw6NiRQQmoFpEuLqgxKAAuwH47W+HtEZWpaIk+sAQRwQMDTUFQCwDMh+bNI2Jt
KITsKFgTjFIZNwhkgXn9p+c5XGHKTq+Y5ycXx/0QDknUOJM0ZLGlSZYf+8Pd7WJY
qcVns73PeMuHWd0KQC5qclFUnivAu17o529UqAaVTN1Ezu/PkNgkqoQ/LnJCHxsz
1KmkU7R1GbOicOs4WzKtSuwE/08FjTNdX0orQYknoDiPFA7MrIA9c81K65n99hJT
8sSeCkrGs9VSixDnj/OfE37H7iigQHFauigrt2WwHwfT2gP5H0CjSmYumsnzskD+
z+xU9G6G4LCGJsEgJ8omsOZwG9MF324cWYGnFAinqjV56/CdkUd8U97n02TM0cbl
xQXHmUrTzQ/KoKSQdjGjMGMyOjRR8uW0Kp1iaA0TxdoBWpjSucNQS/sMQ7iqcziO
cElMbr7uLIJdFmrWAFO6HXcxvPopR6JTXBCdr8nDt7bX77L1Ni9nbI4iGpSdFtxP
5gaN488RMLVJawJP3EoNiJzP57skCdTpbYEiqdk2/t9qf7TzUX6xfsEgIiK01LOc
NxytyeDOub9sLVou5mdZat3HSNQJWnfEgLxVGS8Hujr5q054jyjMMd/mbTvoutFX
lfIE1RPW/+Y2IefFSZnMZpWEOZEbAQ76EIebLVDwS41GkEFITxynhr1//l+Q3Oro
NmPI+XHRh5de2OmdixyM2dQKOxP1pCgVELc7Lm9ttpV/jlI7ppHGAJY7ttECG2gD
nxnSNjgnXb+xDxp8i8Xf1BZqquifypJO+I+ni7HXYVdpuN+MIJ9sOG8rwkd+WGFq
Rw2u+C42AMhy8WTYyTtITfr9E987fFCDJadFWvdcOcwzLXiH/FFsl5NCWx5DaljQ
nQ8cC4M97ZW76cozRHBo5UArc4ZhAYP6mRa1xeqhJaLaD+vp8Fr2wazl3ajsE6n2
Op3u8A4zN1m+fAtCoLOzRYiTSxeUw4nztxKZbWBkT+DuaxyffRoUm+yWCnuloWyS
G8pe/ACV3ztSWYo0H8Yi6Lk2P/rVkYFy0gJQ/Ds5yEi45+ieEonPBoB83KMSYBuQ
oBOHg3YmXwKrv0mp4nZHGzYa8sllAo7/dmlmxdkPXcBA0UO3Q6DyA5HYkIVdpKwz
WaXu4UcUpQJWuNoz3she7q7wN/xJOs57G7b2897JqKPJ1RNy/MUU9Vku0ay88MZJ
i+FTaDGnjr25cl7jEUWh80Dvs+eDGOGYx6jEP4gLUBsxh8n8C2NbnFBnHcj+x9Mc
mhBu7bm8sGi1xT4DhL+mlTxV5p2MXYksPu17P5HlIGL6ZpwUx3JfMCLqa313NIS5
xiBPrUK49rXVWncYWuLBdq5z+ZtH0X1y7HfAVQqGGydis2nrEksTrxlvZosYddyQ
mXlu1Ii0MCrjrkZjl874nMm9Miq0n5m66JV3VdF8Pl+sOoH/0zXB4e1HUk5WIhUC
su3nKWEUcaezfP/H+GvTMsQBMln/CoFIyUPfu17L5um4cyo9YPzUHQZ0cRFvEiGz
g0ICvnhPEwwINFj8w2dFrQA7mnk8dsYJXWe5Hponj+0zEEN31mdhOPhizgYXAJAU
9uP/koH5AjmR8zJICMuJ78LuunY1/CL0b1waTcaAaw5Vdlmlk8goJMNCxD6wdRe1
l2AwnpaEEG4QRbNq/qSi8mvaNGVNqmynvGcVnmuw7RJNTU/Gdb/uDxNRU6svrAB9
AlRCfLdgZ2J3mYUR2xOsQ5NN6vO4EiaMkB1JzFeBBwHH/IBuLS1ezlFh11puDUwO
4Dq/zqj+Xm/Q/cG+uGM5Dk1Jb3p1i1+khLbJugha87qafziiHbnOF4yJGDopPV3o
b0gC2YoHiFRHqtD3L18SPAcoVkfHzGkZkuTXZYLJyJl1aFk47XydrcBBCPoLas7L
Za8Nt9YAgg5iws8bIj+qCWp4eD5C0/bDNJKZRpV/zoa6dkyNjoXP7K6fVclr71M9
RyBYiEsYiu8GhX2FlxCEbiWIqhFS1nOFlcQwbg9V4Rw1l7MQ/DmQcZk2tkzTYD0q
AoCCFIxGQxeig5hORVS/5sU5R4nP07RQ5gKHNlgZFTktbSAhlhMY/TQX2y2NIFlF
nSd6dwfRHFSLrT3ywSu/EuAIW6Wp0x9XTBK9sabd1NF/uUAqFUbeJcBjg33CYdbx
uk7NgLNa016SgLFpqPeVxCW8FAUnyrBn3RkldyZFamu0GFl8mSugbTT6lkkq3+l7
7OQjLKU7HoSWr6v+cXc7dnpvlo5uc00jJPAJIkW0Qtw3ENTExwLw9PHXxkAFJuHo
2FTDfZFqDZizzTs98tGjJsLyz9ebcSeEkZYC9LxkFXb26ZqLGC+ttBbhu/O1DRkq
8PnDLJcthqtECwf/K6OSVMZvo8CZx8mWzdz0+9UGBwueiYiFNw//gQGbiGSvFfar
W1Cmvv2o0JTOThvO33ogpBur1b7E+70c1gJvdyP/xXe5pTPDcoWGbA9+sUgm9NAe
ee9KF6SFtP+5jj/XRZDznPetSMcM3aI+prjQePQX2VDK7CalMpGqUqMQzgRqf1fe
kWSR9hK0WHoXF2v6rVzCvacxrLSSKbHfj+cPPdFOJclGj7r3SrkMSbvM4E/rPZ53
/lyzYay0zAXbCLaXKK9HjCDCsDGYtLpZENWNjZAfUXTAt0D8hHLg1rN2y0y/SF7K
yc2bOBsGbvxe+uiqp0ZuHRBPAwNRWLBr51qXE1/AlAap8yQF4BH8A/ocH9Q+N8+C
IZKlBskljabGpCvlgCLEqCWYBIExTn9znpkzRE2+ANRPKT2gFPW3LlfwvJgqbcBZ
z7EW2dUUckrSiLzg8+8rB1yDl8zLtHiB5S6C+rS4VL72oA9Y4nHuwv2VdShu3fl1
a14UTHjAsIlIvSh0v6Zk3hTfqjlxkqSeBE+SXAYDL1/Bz0/NRm1FnUiMrEMbdh/r
4xeXKMHmwUZ4mktmqf7FzOmtCVmiCO7YxGv0xro/xLuaV7D/A5YYDXNYQMCHNg9Q
qM2KMYwD2LgtXK54iNezGF7g03irB52QFYVvIf8wwQINbhOZRFUwSDSOivK8EPNY
+fWC6y9AXTUx0iRzJmHFWDzj9ZMSCmnXbNEXFwVCADaklRnOtGE/Vu87vAZnAvbs
TA8Rd4hVheDsMEFE93imBMmxt9QywGUhSsDHK9yG/XzLn4rmEUnc0GpxjyO/0TFV
4fELRX0jrKGkMmbKZV25Wth46006jSsi4tUyW+yrdphe72el/zUT6q4kMfEuTsoI
VJEsGzlFZatplVZLa1uURFpM3kBVp4F2IVAbw1JtkR0ApaFf0eVIj/wiTakyqF7A
5ShwZw0F7ENOqC2ni6xYcKkNQuVwndMDgKMureM0e1Vdt77rVv5WtVB1GLrTs9ea
vQYndBVbxel87z+FvnM8MrAOitPDDTFYwzCuxqMld6Wi3M8Felue69ifcQW8RL99
c1qLoqm6q2+b4k3Qf+tEnMFrwsuuouZTjU6FUZu0s+2yctnbT8HJImL03V3wLVdX
h8L2+h0nxgagsVavd3sljfe8FQDeHZ+ewBlDnMpPEJ0LACeKoVhXFxbUGScBXi8i
eiTq6BsXFfPafv+Qdmxh/y5EBtFqwC1r/YMbd9hO5PwL7zprBiGKoJ9kgtxq2G1D
DQPSL+vsiLDGGYqwF4zh0g09/Cj6UIYCGr3i2jU4vuozDtC/oHL8XCyWZlxoMbW3
t8ZjZWkrQEWSG8p1cJyA+2BbP6qmpnpP0jv5EJuW87y8NyvH19ROjIkkJVsPH/8F
+avZp5BDsOt2MH8A02nlwSlseYZaUuLiDoH+GO/+wmMVHtOwEaokZc1ATfSNEvqa
bHlRuolRrQBHTP2pcbj5jMBemIndgBvR0wIks5/AmPU66QVwczRx9y9u7fR6iII9
jeKY7z61/Vq0upT47V1bLB8M3fL5eKV0/mGPxT4aF20JySojY97IVRtJSZiflJHa
Plhv2rz6rjlSW7rv/K/C8ul3VqZulDKkT1gaJHryD9YOwg19f3Kl+ZA8srUyJ95S
0c0Wd07ZRzLn6Uxl+JdP6hEGd6b2E8LWrndhD6uDQZHgkCvGYgIKQQ1dUsZ7V2iW
roiWxCEMhldEmJgBfQOz04fAJeDrx8AdVaeq/rhTZCRJTvd/f7I+N0GbdDkM1CS9
19buvLav1rXsFJjkJ0Z/n0LutvBSspEJv/MqbfDSfXvtnu+AOUjDgOc7j6CRHjoy
yytn3KlnY/RbAPxZg1OYTShTj25LBrIVEapInoToFaxkTkaRCmdZbP4OEMbthKLF
pieYvoI2OxKiDA+K30u3T/sKwuesKer9fcdgs+9/YhQG0g/Cycrbd2EBLKXSjHvU
3x/HfykqNe4G6mWKkGVcKevP6gbCwMX7uC3et/brNil2EGl6e4/c7ixRB674j545
Y2kYUX9iZEtCC5xaS9zuqDWtdvWAC+iAquY3ZsjuIxZxciGUP0smm42H7ec1gdnd
IjG/ZGNUGkcH6Ytmuhe7ECdK7TsS8AJe2xI3DTYruvQ23mB+CDZtYITmida/+BSr
JcRQUf3savJgo2WX4VtqFCHobLrKaEdZ14SPVMSrrX/RwiHmcJMwxmlivY7UXnjY
fCnv/3DR0pFyajgYEWwyMefONq/6wkFJ7aGQTuXqUvQdb6kWg9aBgNWJ5IyZ6bvE
nnpnLK5o78TnO2gdBpmfZojIG6al7x6Pbeo+qn5AZ+f/vE91itrT3+YXbF5jme7k
t0qbYdc81Egf5EdkGuQ2YS4Lp6uKCptFumAd1y53fz3NuBwTHdrCZJTS03kcYSDp
L3whiqCXQ7Ik/wsAnAvZPaZfp47dN5hIrIaZ630DFyymjmhYVSr/vGj1QuF4Qn51
MKebHVjZresbELLMxRNjk/XXBVykyMUHFTWnwzMRDuYQkT4gFpSEr4G7yaORHLQT
1cGB/YEloERU6pAtrKQ7QOMqcicg6PUpz6d/JiKz//R//5nHOv7QcbEvu7uJgi5E
H9HFUI5ryn086d2+E4lrM/UXpHVqNXKTrZwjO0vKkylQ8/+8AGYdd7hTScheOt5u
UsonOCGaNmOeZ0AfF9OqURVfaAImZl5TMaf5+H7N36CMIpaFrscevSwrxlM5K9UY
aMnP9VC+p8APmjGp0m4f9O21x3kK7eSbgnVnPDCef2gbJxLrgDcIG848I+O+NMdw
MpPe8t0YBckSsRGEz5ByyA9VAoM82s3ub3RPu4lLtiOTYF4bRJi7CgQRAAVdH5F+
AxtMvU1+XUSDkdnZqCsrWBnhbuxcyI768N7Sn1LR+9CJvxqxWTE79vst55HelSHB
08wZRYyHg7xmYn1vp+7F55j+sjPqg1LQXPOe89ZcDWQVVme6AQGCOSJsqjrriFki
Fkorcz3RdhjOu/DEn5lNyrH0BN9ewHXcCqEx5bYC9iBA6jHP9A577abNaXq31e+y
qOHKdbuq2J6PWv0RhGXODhTwJtDDaFAx5NkVOx+9W9dN7hLbXR+PZNH2zSckFixH
81ogEftQQP1mpEsgnX8sSyFE/O+cibPJ8j9yuZAn37s5tTjLN1ogFbnELflhb5CN
orvIuRGDE4wKlTakC88yr9cRy60LPFIsSifWzmWQDw+7Rp9A1tU4Binuctc5ch0+
YzWYareFpqD2E3lmSYQGH1fEKawo9dgjS4oq8jzrXQ5Q2IaaVsjywNeFPak7XlbC
m52A2ApB+QsVPJiyyrsLEWjR+MCl4mJc/0EzOvaholxKbPFqOwGPwVvJakztLYMH
jthpozi9S+uDGUv7UXp1KvTrfseuFchm4GjxSl0+FrUE5szJTfsO20a2CZvsFHPS
JEvX7MjMrYuonFAgqKv2OyIRWnWCTJgDv4nLN7MABl8SiCo64+N1JntaKZvKuvAw
79aovLKVebWkaVxky/yEqFjAteCF3gRLoqmn+JDfkS22aAJhuG0rmCcpiyP+FNB6
0RHjvHLMfJKJ7AKfrQab+iBTu6fTK6vr3acrgJg5AMlzj9DtVOwrMBjGzMTFMVgr
KlExokWDt3LLc6xBN1VgHE7RYpEMjl2oqw0miOiHjFN6t7E0av1kYhISTuBAKWz1
DTQP4t3LcNYoWfQJjMlNjAV28DgQa1Oubr7xgo/AF2p1K1avb7Icc+l/IGgSBYGE
FJEQI1XM80LINvKktpkg6aVMKMZcaSwqJVFiF2YZzm5gKCqVCZCFCo+9Idy4Oj9b
v/mpt0C12/wYXETakrTUwAANaLJbfXfOjqUmUqZJKGNwTBkIP2jOCnCqUXCRoPMo
TH5oAVIsV5PZs2OWvxqNksIo7N5ggoI6zBG7HgOFVEZDOVcRDwRNhjyh9akoy6AW
AjOS4XxwUVk8lBbBna0MIYo2gFky6Np3SBqDuqOYYKzUQsJjVvSX/3WDadPQ0bw+
odw3ObOtA3UaVlPED22veRYb0UKyHraSHDpo/ocX//GJgKZbfchEt09OqhtBzbVM
tINYCzsQlDBXo1u/PmqSvEHtfH6aiDElCTz9SOdi7wFVjxD9WPzii60B5alFIr78
O47ctIOFTskk7G3xNfXgaEZBFj7cwrbj6Cq0paNCaDV5OOHz7V6ecI1bRaw4xZwL
7UXEo3Gz4v+FrhF842PHhEFDpY/22wNZfOeUHhSYL7MUVL2sf3y9fExuqf0Hlt5q
6oipeTgnA+RlXoHWWKz0l6cttJxnyUxuI/+pwZslyNfJ3Agah4zxVK4riRNBAF4S
3KYD66cfaoMV2/drzEAyx9HqHORRGVWjp65j/BfR2c/S3Dqk7l4pk4mWmw2Cp1l+
mmycMl1UxZ28gAHGv6UxnbAsKvhQ+ypY32wgAI4lHhgm1Ce+Znww2B/r1of3MUda
kHHSV8aEIx4ZssRJ3fiiOALutilqhHZVbx97ILiEQRaodmKHhlTcaHyWLWO/GBq6
eNG2/9A3Xd6yX94pnCLbBXZOw8AKAtNW3zE2deYO+GJVBJ9dDKqxfYPZBMxVwKmV
zlKOQLUnhhgO731DBauErmVrWBArp72/k48zxWb0zIvf+pQL08wSc2byl2WauTUZ
p9eQne55X6ffVbJvHmPIskDanlTfrX1JADa+l95+K/XVjsmPFCIWS4GCKMUJb65/
yrdiiXo0O1RjO/TXyjaXYzeU85u2tUP21azp3hXwryEWZLNQSBF276DzW8aU3tHL
COrKlqwBWUBLexBi+N+fVF3iOFpAfY2LfFcfPsqrN4wlITif+aJ/emoQdu7+bND+
A++j5Dtm5A1JgFtkGJkSEuRYHFzqtjNRT6qB/toTHfJdjTlq3jxaYIaWGMEjxJpP
6vZYI1X/byMTBW4jlcvpdMpF6sg/oIoKfyQOOMVtTYMuUapW/fn4KhmjPlls9a4l
MmMkPyZMr5ZWAWHpbq+R5uPH58H7mWYdmBexUQ3dw9D+EPCt3hsDTwecROhir8sV
9NCQnQ72b3+d1qcteXyJNNQw3g4Ob1CkGnHj1So8Lue0W3W0toPYs3zNbjIHvG/g
iWbESDSj7dKgdJ4uOnrcbkDIBUQNpzE7RWLnZFCxXOyDN6nhwMeiXW4x4SmnooOz
dEHbxDEKQh1A66hFLEAYnCpC3UDs96zppyjfShnM8Fo5KyBVwLV+9kWbchF1erar
nUoRIYbMtYyjscZDP89D5S7RpvYX/TXdLNHzOG9kiTqNdZxtOXvERjbzzCm1+hyi
Dr1cA/ygLod13smzbLwvsLt8ZrbZhalKRJoinH6YopMdCTHtAuojGzMxJdaXfGD3
LtJUcIhhT48UgHAnWn6NDhrKtQclkR0Jkl0uHjgeU+9b19yk+EzlKPDKnq45aPc6
RUwlwS4n0zuS3ndTR3EPW2AaWNhoh1EJ6ojP+DcvwLride7seacbNKS4kXep4QcK
+raremncPYDe9eElUlfE23Dgh8lkQ405BXhAfMeWBqkJKglUOxC7ZYahUuDLc1r3
ZBuGoPnB+BQfcM6r8xg8ZZ8JgnxiQD/XSWrpvloZg+jabsM4fS1X2cQlIWOaUHtE
lQb+nWF4PchaGgsX7U+x5yku+9VQXadOVt7cPRZUgai+4sgqK/sRqXZo2srFIBtL
i7QEw4V9hMT2F8BkYTxIeHD2t+Oj8hKcldtNSy1Qdh4PbFYNQJrHNk9i321kYuqQ
b7nwZ6QqzEcUOwRF2yc+EY4SJkiMAUax0Shj8eojyrFtTrwaZwx6cApW5BGbxP1N
JWTM+XLKN8AvoELxV7q/kxAzIZwoD+m/MZ2R5wu0hHaEGyLNin4adzIKmvH/frJE
8pT6edBTeS71XzNOrBKoI8e7OzTUIL1qcMumPgTA827gxrnuA9HWE9RcX07IoJch
ZoHJdtn2Kux6H8hf+7ytsn9bqEJIAFNoH3KJe/yvjyJ+mo1N4bpFEYx7Cy70p6lh
DG7btneMwQkIQS71g3YBMKPGAqHpAU0b+99wCHbc+1Pk7wBZCSf+vylQQy9/2oez
QmOrTuSqezCnTwRaadTOQqh+HaEa0pU5Jz3yRVRr6TY5BSw24dFE/+04rVNJw2cj
oxdSL+tpx26kBaDHJ5IG7biQbaSCwSVDA7tjX1gAq+9RwRaFfvUIeOdYNDeqQ/qY
/8iEL0wyj0L+EB2/vUHseHkbLaF2JZP3CKLNUhlzgV1m0Ji427J/ZdxQvVZ3DlVq
Iwcm44Df50tgu7DoLKASAmcN2J3D6wegw6cpbFNaXK7pb1GiY0BMe3gVtAjk3/wJ
bNdZxU+Pw75Swy6OuQnyEKTBXBnhZSosLbOTL9BgdmNoJrxIwv2Si4SLiMHuSp9n
quT+YgPeLkY1ZjA67aFuch+uuSsMX0YNL+Hhs0+54wJGWfjfa0go0cB7gCY63MJe
bQiWeJ1+niptnVvI/+0kjziQ7zLn9BaAIywibDpUcKYR+laHW/zQaRmZ3c880XJX
7kdNomoSuo8QkfNszNTsINMy0pHfZc1P517teglcFOU3AqV+PngxfTZjW/VXZRCV
YDV8KQzp5yVFSoGsBuN0RZULdhAURKd97tE1RPxAySUuZ2wCsqzFg0Bkgl5msKIl
dSXM9KHy+mnb1UZhq/EyK0fYw84eX8DAXDQ5XP0p1hlMMYxbLMTzSQfZ88s/sZ92
pq0mzXhRJUu/xCXbbA59d8R5f69CGUEG24JxS7v5K48PAsqQH0diSlOt5lZiD0Mi
NxXEmoURUMiUUazSclTG2sGpyrbrcLBJTw9E6mhZql2AMlnYNHJ5mmkOCl+TqGWG
fl8G1jqgfYlzfCRFJZnQ4l/QKUnHWcD9Gyaa9LC6q7cQ+EYWRLB4G+w/fYHdsNdt
A9WyU4A6omHDVr/WOrwVwjuX4rKCm1K+zs0XLpCSERRvTJS1nNSzHTx8nGfBzjvr
tN9BHalTvgNR2PMi0AdfNDNlSBNltnRIbD2UXnFUkDKqD7OWz9uphvKVlGwu84Nc
5qvs9ZWYpiu/k9ouz88OwONZGRRK6XTxcJp9BN6pR7HD2RoAsf3Gbgw57rAklUtE
8gPFoJQCmulo2O9bWPgqbkfVUQi24oZexhWphVZn1YH52D+ZKFL9nSWsJ2giRnVA
yMOx5z+c1EP5q0o1PaW8n2/4MPQFM7oF7HtlOuf/hejlKrFZ0qG+GLtAVl6rOf0K
sm281pRPa931pAz11ujHs8sMrrf3G0e6rQydCX2vfXbcj014XAlC6ap0FHTHqSQ+
eYpJoOu0XAPvV4btMHvkBcHJQ0bs9EP3VPRa0YwqEObVnbs2ytlNXyOIYOEgcR3i
y467auxjd26kmuGxes7BWlXrH2gfA9JH4d31Ch8XJ+CWwF8WKANoGna6daMkptX5
EfMUH3Nb0UWmhokXO685wJAYwujFTYX7OMj0Mm9wTsqY4u50L/xDlbkDr4GUZGF2
8sX5yMiyYCMP6sbtx8GEutVcsxSekru+GwJeFhAANIAnZ6rkq2+tf4rRzAVIrOgG
1AcEufXJssiHguM7KQnSeHfdFI9VKL5yJV5nTIvIcigJDTqVHu+FBXTKpSLhx0o1
DWv0jRYot4RtqMChp5TivIq186mkrRtUTdnZ1gPzNIPkqpDSNMOk/wftK15qoCB6
Vyz5XIxL/C97VHI2SOqtldY4Tw1CbiQCsGO8qxkWAFYkblFBA2ArswnX+JvVP1I1
Nxfsa0AUqj+VaYgFWZd3idbQhptfOPwGXUg3CMPHLZr0XrGPz2PGIRtkiHYBypmQ
Haukkr/2q64D9Qwh9JJnT2yYpGqHMYKigYn4F2CRdFv58KlCTlpFQ1hM0qOeVYzn
eY995bDM0Cd03sTQdHWr+FXMO/Vz87k5ddXXH64IP6dLncc77uN+sgpneI3qBsi3
I/VKn13+zBmLFE+7dJUDNkBlQ6qV84Uxc7IqKbQmZCaDQJ6gLbNZ0wEBqVvv+3cf
Afijx0d7NZh7jY8BJtguSYtdoXMv4tHRY3mtVDnsS/IeB5kQUJdKabhCI8jIpwju
jagvmHnKAAXlsb3Uw/4JdjKZHajHcDPLPqVw0fX1DJDCLjiBAaNson7XGd1RHU10
v/wF+TD8iBaBhGuZEZDVMEkA+z0fDv1CSGwabbR4kefJRebg/W5emlJTedw44ehH
zOruCYoqcLFH0KKulZ9/YnA3pISMEJz2UgCsi5Ds6K6ANf8Kn1uy7Ipm6vVTxSev
a+eiSXV44Ieph8Lc6DFurF3uocism6tgT7ESHiHrNwwKVlKmoLN+Fiqb2tbYhbqr
N7qMirG5nmVKrmVcDkeL/7OdnWxANwjjfFlUe0Fd/vvgFC0ScIGToIxAXZ5n6Qh+
em251MZIuNkhcFyrkn6XI8NpsEH9uxOzhp/9XWTzK6CkF3wTHh2T5I8/xTxP5hX3
p/0a5IHaGL4kqF62dw1V0iuxLCAN+9xfqqnvLwZLI9/DJau/Nt1e39cvqAWn2kCU
kguxwiKM1LSyXOiLcWNPWuD3RL4rm1/sCiGT+q/vw5BPnWenr7zZGpqsqA2S1Ao6
SMK24CG/4lLf8u7lcyqPaTdt1BU3FVS7hQQabSxrTfdUSrJadfFlmxKlFnuwlJeg
JBK9xFLDPXyS/D6eT63eJChIx8STLvXs7s19BDZWLUrOxgjGaDxa//PH9fLcGRR1
QhBykw4MIG9cZXEh5C1J63nd7cLEpW42nGpPDGQM+aWrj7cXVMk7+nDrYtmyQJWr
LFhbtHf19woftbZSi4yhhQ8x4QOYFC+eHDp9fW+XpEIlJ8d/GsAD2YI0UgOy0MQ/
1QnrWewSHf4C1f7JgZE70YoyZmsWDIM5fofzt+VA0yWyOOr6IL9Bxggmko5ZpsqN
hZT0LOHO3SxVMmRdU/8GT5q14M6oTKKSYbjmNdqkQrROz5T2brU/dWDXvh6TJUr7
CftSuB330ZTcbNQBOYMVYtxYoxbx28eeFxZeXc0QhZTVl5yNQ2xwhYZnJ7JLuYar
XnHWyN8NPBr6aZzhr9uUvUZ3htWKBJXT0GDFNYj2CgylNff/0OY23sPDhmgpfujO
jBzdS2hiuKMbYVNYdQ4sYFzNxqVs+bQRIBvtaVDTU3wYbXBxK2Dc4U55hLzouAH1
aCkdPX2xW31XSjpW1J7e7qSWgWV5XhRQXutJoLpwngTwECpGcyZt85eeJVq0Spus
5mWItQEo4g9wXmtxECNp5EZ91nXRS41romnK9HqIGBSQjGjVDKh+qL0HkPS/tzMw
Ll+BwzbmjGs0J05vvg1+L7jKfrPsl579/CC/hwRxtYDCv43V+GIqve6gdscOkUnm
kHpv5T80DXxHp/48jIWRUGWdWG044PHgAelOPsaEoOss7EuxMh/KNtD3rcdvYZWs
atxqBVM+DwDeXuWg62fUlmJj3fx/RKr5C9BjVXUE4Iz6HXfq9vQATJdXw7a5PaJ3
cWdUuVWmvl9LjYME7InNZkmgEPG59mvswt1Zl59jT+CySYzfv3tzytFp//LdzO+a
F5EUyZzeUVcwgvCO/lMaTOa9OKUYJdCnbjFTOqGFmC8Q2ULVAl8EgMhN3P+i9AEh
ufcT0aI5VRPdJmZhnHKQsf0ceUnmYearBWvqNqhe7UWrZn/GMowtGyaAWEkynhfC
ZNng2IjT9epdSokHgSiK8g6zde21fuQQP2c+swT+bzAwBwEavJhG44sAQT3qrfLG
3FAIj6ZFZUq5kEOUeXPUSb+O7MtBNRB146IRDLPTwqC7Uw4y7wd7AIKlXJVgKgkR
0DO2Kt4RAXBqx+kNzzJC62zVzBFPusuTL1km6yllcFZf8F31tWvqwZ8ClVYgXb8G
gG2KZwVtPd7+icn/7YyBCOJSMpA/9ZGK3yRdpREZRxGweSsbfTrVawT70FNdhNwJ
x5u7H1CBvvnJ1MHzcEOOZ1XTBEFOPF4q89DG10mJEOfbAVizos9Bqvt62GHbe3sw
ozzVz26MUzkMWlZKU7yfQEabwfEr6932M1hwkOnQAcZPsqfNTZCaZkfsVyVzhmEQ
87F8DF5y7hmII3kAUcHeY+rDmqrdCiCAzLs9ocjHiAG08ITD3VKoYd6QHEu208ew
pUg3TAPFVoYQtBHQD6YXGGgvabkC1uM1d8Re8E08WJvTqb2DgV5QC4dBrAmx67gJ
5TFlKxnQGPskG/hE8NQRmxEvUUCL+yUbCeT42KCLAMV/FEI13GX+xTyEhiM/Zhh3
/oJcKGI2aTSEzP5p5z13SIi+w+3iWne+dMjz8I3kkNRtDExyGjCGD4fFOc1kSvVQ
4n5JhnsLpl7Ag9i/qAB2qAxnpsp+uXshK3xJqBMpDsbiptgMOrX+71XLTS/ucif+
K7Oleg5a+00gJUdoD6xKvJD/wq1jKP04N6jc7tdZX0P1Z9didp6GS6Gkqzjaooqy
98RCqnhCyeI5cUL/7GUL5OIiYEhQwtTlsPrPaR6bhPeF1FrkZrnm8k7NxhE3SscM
T3Fa+z431bgq8pGUC4L0YIlJK0dzsaVnRFT0/BItRpasnz5cEXGYuqsVaWGk+lV+
gQe6Pzz2tBiiZQN0fukpWhXBIMGSqZo2i+DMIa5L4HV2hDdo1iuuqBvr5ADXy5ha
hjHffXrFDnWuzCAZIx2bx46e6rUtqETZLWEgbGg+OcM0KDp1TkaGCFOxJuOuqk1v
QTBqEfTtnX0oUg19VD6pJQ/NO+zJ7/cCKBShWuP1GuCQDdIhFtVT2iWSDfrKgkNg
Z/o0oieMtdD6hAfAXUGmrkrleafcDBuVhA9VlZN3Sevl6pZZRg8lvaVS5CgPcSNS
KViyt6ZYg+OIZG2jzDtzvahiz5yB6Q6ePxGgfsR78B5ICW4Ra4M8XKXsGlgV1in7
oJzUGQAWD+ltGA2q/ilN4UdqfIe165n7kCXSvIhz2pE7FWu5uLf1TYtfwjj/gdfa
48pbgG/jGikHTMWRkIn453lqR4lZQQW2MCO+6IBH0pRkfaVzMSvm827/emM053MU
FgJfap7BHrSeY2oUlMzYs6DbP06Sq8ZUqnUHJbTiM8L3f1650UoLF+dBuSCVVlEv
7m6pagPzb2CJWIo5QTXoymJJ4ytEXS34d8Am26IORvQMMdc47eDvY8MJW4RDvt//
1cMBMwzKXagk+wD/xXNSog2hnhKsYaCClDzF7oeR4uzF1f7R/sI7YnAT0ngI4x8W
wQMam7xmj89wo53kY5dPphZTTBDryyYDIRy5uRGIAuelYDuI4QJh+BHAH6A5U41Y
fW5Zq1GXrsYi0WZwt8Iup2wXWGOdU2j6O5d/szpoEOKAUMKkQh+Ul6GI/fRftPWV
beP8KVsGoc9QnBUQQkeHpp7NBEGCqwKsIoAG6mJCRK24viLnVQwx49cuVFXp/IP5
ygUF1y6fPXSBy/FLVreNn7KROChdHR8gQrOQZEwHvHxbBTytO59Q4EfEhNLz2P4h
V8xPDj5ODLQFruDMd34Cv2rq0wcRWtnOucH6KHNt/PJ1/dRvFlsjSZ+0E/OLOgfw
yzi9mtuW24f9zH2M0txhjS3sNR4KylcURzroW9IMmNzlxP2RGr9UcxlfdyraeYbJ
U1LvTAOd0+mHDTKXgXBt7DuelEfqynNeW/iE8c2zUr5uT5uuN3Aw3skjHZ0Mabmo
Z7DVFZuMvn4ZoXp0k19qX4VOgKI26DhVD6NfqEJlgRnxHYC9rA3sJ+vqBcsFWLd3
L4CusOBojTx2RwqbO9yDK9lqImx7XrLIzSVYZnt1P0lDZnhGyeMPACmZBgD0/Yjm
OzUa/ME3p8f7LLHMcpnJn6KFQvXfyGlYu8COHuQtGi2Rtg7IImByoiRrxV7t0f9x
lvJ4V46gjQywg5vULfo0QoRIQevXh5txbqtFIWlxyypTHtsZ6Ji2epDa/SVKQr1a
ZooZao0MLqjBJ+MbjVuo5QssRxI6HXwqmeoJdmFnoiTr7FsDK6Qspc7GObrf6Rjx
7rBpJMlc+J1x+re+tN/ixKWjT2z2kG4lu2bfJ0eq8bRQaAtfpMgiCQ7LsrVZZHRc
Mj6domhn1tcUgGRxqToE54Ms4Wxwt1xE+QZBuyNgDtNCaWQd/FdxVdd5Grrh/Yoa
dB+iNqxOgbRL7hlUVMyCx/+tDyNsqDK0LeB7eMTVKppI4T7jiFG8CXig+4gnAKGI
FCWOTlV+fhemmFPZNLv71SW0tbskdcL1FNx5c4F3MKIKgt5NvEYeY/m9MbKrGDUC
RwBodGOK00zxiYpiwpB8vvGz+ncp1THqEWvtRgYoy3bzcDXtOC68kLlssuuMSeMl
YBWtFHfePYpF5wU9uQgssespAZwC+25OIdUZeStIBm7YX0WJbnJ+UFeRrs3yD+QZ
SgCr6AmDL9PHgwMSEDlY6uh6f7lN0qp7oV3jrRZmp8N2QDE6POy3isxR0zc7lARI
yqBM0L6/3eKV2TBEd4YG6yQLZOijd8r8mNCvnGwC4KXWMYk+lDPqCSf3I2Y3Llca
dXbEmutqBGVUZAIEjJXn/hqh4UmSUMFMK2mlBnYvMfI4rmqxbdaJfWqaynrp25FP
mg2+lWbQ/QhGAwtoFKRkaxpZPHzs68R6zbDPlIK2y9GE/ieHVavmWCqcZ1UGSLyA
icWTjwv1ki2asdoP5SCOej1LjIScOVIxy/oVtUCzgN7UQPdlRpydoSt20iHIjJ2Y
E8gT5R+THw6ZiTZG+1hrYe+KxAlm+0jQUDla0ZdEffZR4Dvwj9/aTIMoFLJEAofr
iza7GjsagehmIkiRfZrI4LOs006Nla05DKeJT8Qd+agli5fESs0e2i6EvBDdPTjj
35hUTJMRXlE/R92FxYi7byh8Wu6eLSLeyHuHb6g9WRrITM+7Y6p9Jr2iQly2SeDg
ruLmRihiXExUTbVNkHVA09QcOHzauhH0Xc9zlSb6q9oipox0ulCucq0WyF/m8VWx
FJBxIZgFqTJ/U+jkAUbGjcgqbaTLl7kr0gbGHSinoaWm/GVi8m6PEyxEw2/jwHxQ
lUO/X/iq77vtdwfENMZRLUo0owpwOKYcerLWSH+7mMMDOPxEf+e7bazPZ5j0vs3Z
aocTlXx5/TGxeGU71yunxE5sj6ufdbvr0Iqxh4sf67txJLGmBwenN8An6UrfluRZ
cUuMdEqtV2Z24Xe65cHZD9Wgp9/ISn/cT9VWHw3XWOhBESL5lUQrmLrF2BqMIsQZ
o77Wxp2ITxXQlrT2m9N4mumWgKuR/TT5xIat5cujL8svURCnUcFa986ZtLguZjhN
VBbNkMAJ3xef5CWGCi+4REoTiFURFbIQbhOEHAL4NuZqF45PXJpf2IAiTgJAJZaP
OW8Z+QxxthBxJx8bV/IBanl7evy4RitYa8vB84agLFXmo86aEdLRNs8/ycag5nUK
Uxfh5pbtrN9Vq+cZpclTVbhmqDjRt3wZ/G+JyFS3DQ9tV3whax4ZV/iuUT0CZCCU
v55hIR7dgQ3KcozXt5ou5xblZqkCwZIB9JFD8E44/819BQiHgRNWanfDlQi9yoX3
naLhVMiOBAq6y8e3bpsEX/taHWxf1cO2wGDOVG8ZGPD8Ny86rKAGiRiU8FQBfgjS
d1pKdIlpVmxjDVhclXlbCIHf8m3SYaUCAy9y2U5JBN809BEdQjCLP/KPnI8NfFC+
MZXfymT6trGgW85F3nI9h0Eq0yvOMQ+2umbQ2EE5+urkYGMYir8mzB9nAtHyud36
DGVrxs9W/3PRgxmysgu4R2En4brnF8+ZBZ2yYTTS3ZOS8heEOYKcOc0hozOh6JGJ
Pi2pECGA29m6GmDyIxe90UExlJI1WgfCc9hVsZLUlQtjzxtKe9UF3iQzwO6dWLcy
KuNZA80QTpFEg5t8Yp1e+edU4u58Kvzez852La8zzGf/oxfhQcF81xGP/aKaywje
hoU9fQK0zIj+k1WwceRzKTJZrzDghoyUTiQ+u5zfA9gCgTJucHpaW1Zp1/xRfM7i
NyepTU4FtsiV40s5LTw3edWJ0gl5sdq67KrewSG8vCf1f1NvKzPfpmdpJaXGGR/4
9bG/z03uazemtZV2cstDQTu5JAhDpm/sCPjOREb+ZD4Fnm4Vj+A4JyBTyGHbjtlf
MmCtPfXQ26OUgEUSZtDrxk2Mgk7XcqBgXzcb/dTnUuPctMdPe7EW4fEpxoaJg9Or
oPZJ/34lshemLOyb+K523qW8m23hAvu8F3FpBzS1xaxuVSX7vc5R0GIHxvNSAr6r
A/ZdN+7pB2ik/h8W2MrPifd5OlnIEbSyf0UoMqeZ3DC5rRK2hJ/uyINzff22WFs0
rn5VSXqfzVdTIJFfisiL1vxgyV+HE1xeisdzDSNm/COPdW2fRkfmMNNdX/BYJOCU
RXHedI4lTj3hsL2IEJNnoiUSgwkz7ERKtPWq2eFzQK5rUoy7WrvyIfnsSycDA9rU
EuQUrC8ZbSzKf3V8I96sVypWGT+cPxS8xeKDq0tw/7cwZPO6q7fHG/vgaNp8PZXW
Gh4N/ORjS0B2PjngBanlvs+w44kR3pE99ydEpKOGsAYp0TalpwzONpROliV/XjQ3
Ya8iCiPbur+o/tanQy1AkQu0SUaPsM+OVY3Y6o/GK7LCKfBDcoyS9SM57Gmg8Yrs
ZYwmQclBIFpYoUyb/j8wSVPhk6W1NccTq08aNpTBxa+p2MWwMotjzbcLUEwAIt3D
kUS6BLPJNkshWjz3txdXdXX4k37/rtKduQKxb5wA0VzkeHniN6/ARZJPw18oQmy8
04bD+LyBOM+vzzj8r99eG4Itr/C6FtCohA0Zz4/C2W8JNObzVHF1Mo3T2MvmlYJq
6oJyqawURko1tYSpM3FNFiPNRX560PfJI9cCQNb6JFpM6cBMT2HAT7hkSn0URjiR
EDIPoSUF7fo9EpRHnhr+TC4Q1QFoffvKfdTBR1LA8gMCIhxpAyrqqzJDnLMN1cjP
uSbgPF727k/ipiCVRAUwgb5PwrFgCzDePN0+PIPa69r+D1oR9R6GgLeF4ypCQTRZ
VQYCkqw8E4L8TJU3rHSuMXP59xlr3ro3K/pydXbHYIw1xz461QGyrn1ZFO7bdErd
8ygBOJyW6Y/29NeoQqZAJNxz13wlYfoio+b5ce7/h1TK58XZq8EAiLtQ5apaKH8O
a0iqiRJfGGCCpwtTGyoywpTDFpSXtNpzqHdIEXd5mphp262hskTXVp4LrGhkh1oR
A+JK4/a9ofAQA5nx9uSSK3HaOh0FgtN2GZHheBBjUByIY6ZwaM3/PH9u7k2bzwOR
inI6W9BV+5Mp6vbnDkojVr+VQ43mxRq+cs7Upne+OgiIn3nc7xz1iHjR2CZx4OMa
nExy7+U28vcu+j5193Qfq1l5BdCl9k5HDPevluRGDtei2OIUysiTCUoqnAfenZ/M
SqQM4wvQT+mZfvCzCkL8SrGfSm9uJWQK1s30cPM5Yt0UECsI+Kx/84bXTH+Napos
wrIZXm+VyDwukIe8bHLq0aMuujNebT6zR0KpRCtILaZCuxUPU6qIcL/AWnyzgwEh
09rj0DIvdaMLTuWQdNJuN4nqS+cd88Y7nrvE9++fJwVtA5bClt/lxrt3UUVhz2LH
tsLien7B2atyfbmrpZKxYWfMuftocaL9Rtix6XcRYsdEbGqTf1CiqO2nPOh0cu0j
1g+AKDMb0SZArYPhHBubrOE5XRVkycRmDjhynz4eto7Y0N7mUjAo+g7VIxqtaV7/
JYeIe7Y9DV5YdN4MH0GhnI/p2U9YYYnZxZ72QqzeQ1ttIVxmQp3YZrMQ6k5+39HQ
6+FJxxs0AvzN2Nz1uDE87BPLlCkV5YqPUMifB2dHi+Om+viBYG207oSY5hjaj9lv
MstlkoAGCePe5UQYMPWC/yKwDrkmhTg7Z5T+XQ8PLIjMDiP7+X+stuwE9OGqqMXz
W89j01S6tlSccsh7HO+cBnBduEfqUzPWrd6U+hOFGEeOd9QlWzhqYygzJJVbAdo6
92Qikpd/O4rOe5SAkz5Bd5Cqrel9AqmgwlXIM1Jy2UVmKWhqQe2Ta1LRRlaeamwl
zA0cuAID6wARLOVyj6MocoLI/rTP+8icRS+QVhDranRgDje8OUcAt5Yr0lz4riR7
2SNFM3JAFwjSC/QdrbooH7liZvf9jSMxPTDL1Z8oso3ZUjBp98U779RvtnqAJM0C
HdAj/K+FJJy+aGaeurs3Z5kyoXjhJhxOre5XJ6jqlburSpqrE/luxYaIhVHQEDjg
e4wF+9HpwVblxuNHZz+02pPXbl11bhTXCAaUNDxi0bD3gvZMJkIpNLMTREXkttfU
U+0hok58Gh8fkfirEm2EhX6io8ZsPR8vrJB1EEvj4vpHJc9cMAUyRf5kQV05p6iF
rQAsniVmY4BthW/ha0r0w4+rXluakT1n+9UQGEeMYyEoCiDaqLQS3Uy0v9Eln/8Q
tNKwRFHeTFAM63dFDVzJoMZmRhi9uQIkSKKrf8J5KPxYjQpGW3L3ea3EDWcpaHIq
WFtJIL9auh1Bm8XrI5MwvHU1wdeTsAWgT0OHDRMJD6CwBg0tlz0cXcXR6yFYyCRx
kKPXytZQVI3pv0/kmTSELdMZnwBZyx/F61N+mIZHP84JqwK03BIOWpwhXxzES0Vu
3Xa9qesecKPb09H2uDftDYn8Xx9c8EbEKxxkNZKmPKJrhDZLEtQKkg+zIsEeUGNc
AAdLy54hRvFBbqX6v0lWp9wByRnKjCeq5edC9zOEC0B/UGi0LojyM91Ic3pokw+7
xlLQ5eqiWi57BIDjEC8I3LSylPsR5TFh0ZlBW3h8nZcNE74qXks5iGYC4KdNdvU3
1byThy+CQsolQnbc1mMh6FnVzYYIVVUdi2OTPV8pEkwUpXqaDDVSh51glWwmrC3P
v0hK8OK7qnbB0WfDwpsCwffjxWEkf1y6WQsyVczNluKLqUwURsy/sk794oq10xiO
D5EZNsGX3Bz9UJ1Af9YNx0FqX26Q8POju3gcnuwgNN6wgEEzpsBr8ADO6EciM2RV
DnNxQPUVvixStsDnbrWXqwsJiWGQ50S8eaD/TLIAXT5D3MxCG9vU7kgICDvAQt83
b/Tp8uVcYHQ/xGLpCurn68i9SzfSXZi4/gqNYFwHqKDpsqXzK+oA31GGMg1ZY46F
vXyls8HaQG5pskST5XTUALJHcK6uQIH5f6foWPrf6fBvzwyJcfnTCZnjo4hyUikZ
NYe6+6K1Md3oPwPgiZhYpZvgSeYExbO7DXv8kf/4SUb1w5zuc9wIFlqv9zky/bH7
/6Ig2L/bhBMzC1JKMn6NS+FsFiieB3z1QRjwkUYvm97fr5QfzxZ4O5SOvBkhi++C
osP6kHafVfsmiSD47vN86Q1jDmQfuvZ5loQiaFJSB6CCuuG8ydRuO2lSF/FqC+Di
R1bYfOjJsCVmyTa7L133KQd/JkVvhVTxYTTESlY6R9dKUx2yvnYct1KidTSXBtEI
LG0zUBmpsARc6oIrsM5lbsK10qXniqxCx75ASqkXv7+O5hD/+DQJPFuWTPtJ8yYd
cbobjOY5E/wgCjBSzohCstiYZL2TUHTCghgK8finQOBFblNWAWWoX+BRv2P18UJs
Yzryr4adEU0Dv36UGzZcf/xtYBancgulGQjWT3Gu5IVRIpfc3WOfDFlRA0Si64FT
4D4LeW9XZZThcCXq5tIuKwbULml/HvKT2G57Dy6Fd1e2lOiOIbKzNwViaVSzcFx/
0jAB8plr0aZ1LQwxNMpAwp6QQc66y4Fhk+Mx0IzL+fM/tgDUXR/7ZyiarBOSK6Ru
OK56XUSiDIjbR5oqDmZmw74ZgRG7ws1zMUGVtY0RmsweSAtmVObPVgdsBEWS99yE
R3NmICeLNO/XhOFkgSqfGavkEM+3qPG4SCqSjRINLCTIZ6BNs2BoW/j4TFuAqRkJ
kWvIKqH+93A1A9JEFxQMvfduJ6gvTDDoEEv/RVi6d2r/61JP+HHRJcxH9ZW1bXkM
E68B3/jeGTc1Nvk8jRxpRbYmDhXEmaMBdZaJQouOfgocI1XGTPO/8u5+YY5OOI5f
c3fxmL0FqubwaglR6Kp5PYoQfm2q+2X6GnJXE8M8wkTipWF9d1nqHWl3ABEylPgj
Lm9RSR+/gtAfxbKbJumtlPOlc1Jr52SilzyeqA+akdIwAaejJgJTTagUxyrAM/jo
aRDCvmN0Ve4KLDI+kbi6/xe0MxW+oHE/4x/wBN8sMVDNp89Ogy+Iso7vy8EgNuRC
pkP8ebScttfYuLNn6ojk10TXyTdc5/AymErfCfeJ8hjqYARmS05KNWsmTK4JAJLQ
LjWoC8csqsH+U3xecxB5XCmmCQpBc9lyyHj1TWkCB4Fd2v/9i5Tx/9Z3kWsL/UPu
D5WnzPEOuwhyPJhsVGImwKdZ26rTtq5JWPRt+BlGwTATr2leODu+yQx17WduT6Nr
6BfbUxDo7mal7THf9pIjoD7z8izdMvjX6eYH9c5qEjt1eFpUd/t/FUpteVM0PQ+S
EvrVTDr8clVSScUxraScI6iOM5HxpojL5woUcMmt7KSxJdsUOu+mTz79TXKePpMc
iPi+KMQqTQGqdr/aFutarpEBBi/4HGngIN3gcTteS5O3oWmdzJse4yTn7iD5mi6x
feQzFSskRSwa4ykf5eOWaq4vVOzDybY/USgxk0V8DjYGnsKiVvZtoBo0HWLtPNf5
h+i32W7p78/YKNTp8iPzA3+0QLfkVcXOE/ES3V5kY6bKCK+eojUspmWrhTMkKsoF
1VOfwmpF3nkN5Bp3LueqClLce0KrQ5jbsSV7prmuybc+N1Oa0CRH1/QTluPOZ/0t
sDB1XKYHZy70Jh1VFA1WlE5uXEP+04Jmshx98j9nr7o7gDQLGN9k1BYuhjbRUX6F
zdVeATAsfIF/Y006ggrga9Ahb2xpGyoY5KLXa7IKmh/PxX8WhFGgGaT6cPJbYJS5
K0Xbyb/ywaEuHIEr3CHN2AS2+I9zSsQ7wFFJ1JWz/UnRb4Gwbhgd7+BfOq8+nAIO
4VyY+gM8tE5Wu9r8HUAhAtVvsmK8wBRqQC9ab5IXc/PpKOdAjw5+rSnUtZgZxSph
bVPmh9OcbXy15LJlnw/FKCyGt+8PEceQyh+7JTI9mw+L/JWsVTz+npImaPKSeCh3
uWCm8Bp6ctxnEpQUMAdLmj95MEkGLs9fhQICiuyWK/wX25J1kjoXR7kzjjpHUmGC
KqgJrfI3dQbo/eW9NunxAxH85z8QPPEn3uB95RSoOue77w4ECB8oe0+FBD38SfoY
iveQGkznXZaT/IorKsk64+PvDi9FyiGOZGObTGy9b6wL4GxOKPD/yILFuTLH1q4R
6s48JAtGpo9iE02HZFjag18H+5BTbWOjbco3iNX4DuGBpXataM4eRcil7TXgKNsP
lVhQaCcG7X782qho8vZjDnfRk35FjjBNP3BK0G/OAyyYoLONambIur7D/1QbBr3X
YxnUmgUu19J0gFF1YNk38dySP1An6e6zHRAdBmbvNxXWxKMXHMg9k2MOS+RhpNqr
YpzG4SaVfjCeAh0cX0Y9ZDnbK/0X8tP5EkxOdBU2ZTgG/uV2mfd3TPNAQk0gnHFr
i0995rYLty0g+SvpaMO1mnIgf1sV+fvavin9VHt7NWfVEtuTyMa3U3aFZtS1Yk+9
X55MIgk0tYCx7vYO4QzSC38vy2UxVjFtlbf9C7/l5P6aL+2JRCFu49QSb/HRwEDF
Y/oz1oLfDFzEMbXlOHqxGjzrlN00d2iRdD5z/o7DftDxErNOUGkZuBJI5Ev/Z3Nh
9zMStcmggt6STKRFH8eoGWs+CQVPsTC6C5YaFEtyA6j/Xcfiz08zQSyxQe2psU8A
eYzLk+XNDQsykprlgamQWn4RasZAEj7WG+P7vr+W4UyW17ZWPYTd3d3duloouNan
tts+os10y+eugFcrKqTA/uLC/MPtyQfIgxjTJw3qc4LwtSieZKZFCcKPecxvgzyK
RL7ESUKfwpk7c8hQ241b9WLaV+SNuThQ3A2www8F0JkaBBxHaoBnaSOESw3YnioX
8vYaSztG8TSwUBWWZ7Fza390VV3mtkgrXZnIV2Ec/cxSI1dClEiSdE44iG3v5qc8
WpKd+mr8GxAtbS/lF+LLdEfvQTwv4i0OQXs5XjQQgRYosMOPFaZh+HuX0yRc4MW7
OnZPnaJOUFRMTyFciWpYwhUVEMAgIzFLwu6OJ2qqOfNyZcjgJ5Z8vDrjMlR1u+1P
EdSSmuu8JzB1sj+xNFFNc5mvW8PUlxJop3HygM1Ui0x7SA1Fu0WiF+SJrdoJuvag
fz7PsdMQge4umH/M5ohAxaM/WyOkBlfQcJlagKHA2wfeakZMaPSpaRI3I3Q+1t9N
Z/rW9DgLWa1+G9kHpEysj0HvteGwB5sBZtEU1UMxHdscdSZ24bRG6jhmMpGFHbK9
jLzirzSmBcoofVymp8bFpYRxgWJ8Gbg095oGtepTKpaQs8f3+fVWJseVrEsc6lhf
LjX9G0nZqLEdAIncL17z/VSQRT4XEU28is6SLoK1h+nrUcM3gB+HGZHgSvRpZarK
/9q8IH7BEcQztP4m5vRLWd4L+tlHCBDnUnbUgUV2kOlszxXcMEwZ1QPF8Jyrie+j
ngfoyFkjc2ibzCC7JMyJLTzuUE6oWbelFmUXquJS9LJ8ufQzUR3X0tnGgl+BIvve
wnV0A3lNKsT/q3gftRsIqgSU5yS4KpiNYfvWXULgbBld8xjLNedJhgU2tH+yR3YW
QyG3rlM48QMZFk+U00/IPaThXETYqqbJ5BgNcNhbrSZ/iyBMTO6uceGRPKWjxEy8
eGvWOUUvWlqlfQW37HdClSltdOXxY0Um/72YFt1DOq/hgwHsaRMMSKRC8IJOJMUU
/Z5IHiXRsBzu7B3rQ7d3Khre8UCRK9Q4L/KUCWeh3kjN547DEESyCu77M7jIOxRg
aVyLgH27hbwfTGKpdIzB1nSu3nzc4DUPzVtI1FoM/QqI+jO6OjjnYkL1dgY7C9Xt
wZMyse4K85y3/PJS6vsccrZh4E1Ti93MmyHoPYQRr/mxaGPgA32HGAWxSkgJsPQi
dI46rMAIo6yZXJa5fogbWEtKjX2+YXWKLZ83yLXd4cOr6ku8mAUmN28auEK48cp/
V7EUpsof5ekgrnF6S8UOw6dZYdVzZFEni7E3dy8sj4M8vERlWxyi6pXTPdrbZWOP
e+vEXrSQ048ELYMkZ+Znz4A1cqIkERbpMCjaWxOdzewMvwSs3pKL2PNyQN2WWiRN
rXHGz974EMbafcXF9UbNKvodfbkUOr0DgZDBj35rmJagyKvV87g2+xHMVx1Ss8r4
JKcgJ01u+W9eAmHPwsC/DczsAVS/5f9KNpTOMxhImx8/FsgOV19ja17WuvO50XbS
nWpgQqQFWCwI9JuLxlt031wFS4cAoTBmHzxhsBdnIQOFwdTjYsFkBIL2iF8EAUzF
hJ/xu3aI7fwcD4KR2NNVFpljP07To6o5P93Jl/nCScOAHM1hYNYh8m2Kcl9PlfFr
IJXxMoa6/uq9+apvzQHXnGQFeHDUnsNZm3LJxYvlK1ELhj8SHD3qxKxj3xLg00EE
JuiQGBHLuF8yC3Mks2TI4saLyHZ0aV5/jDTSsmB0RDVWYD/uC6VauBembvBaXg7s
wFtNDqMLWxtXKCy5FAjA67H10LOYtw63Qdq/1rRXpH+HIE4lzL3hiCVMlaaz0dy/
TcuYpKgloqMQVvZF+xZ8llnZQ/94e8RkdYu+JBZo2U3Mk9NU5++vxL/z/JGjX5FB
ArOGLAV0x7eHf5yO2QlkybONHaly8FlbX4T5EzRZO2frksxGAnUgjxN87oL5pccp
BbIcVfXfloajx2b4JG/KaYh5ZefSSvsUZ0824nDyu3rqgdrdFKf/DoaqwYFF4SH3
tlLSjL3UL47VlqfV13wm7ej7tLcSuhjCg8QMwSD2E2GINNAgHdRQmOSoBAvGfUQK
Wjt21fFGfgTGHFeQq28zATbZB6kOwbZ10aR+jYOvIBc8ZNvRmAeyLHZutTEAj2Ps
I8EtwPhjppAAcqWtug+/fKRYVyoBZYLINIKmtUv+d0PN4A9P9YrHlERaQYRPYhch
C+DWj/eYbCCkqKW91pqSZHgvya4DQpUxJPDRetOgD2ForoTWnrzazlCV5YSIInGW
SA7pfcLEoPmm5HrFvr0gSGAoU4bTnLydO0y8UizSiH39wYXxKwwg0goDZMgXY4v3
GV8m3JB2Y4NAnTuGgRaqIo33F9bsoBBQpVFdRD/tjgZppQMHqlV4f+m9RXa2PW+k
nhT0nUqOv4LPfqdXIE/HqclJcCy7bZGJ2yVUArgXq+261n6Kclvx3ZMc9ACB+tF4
kza7SuI6Kaycyuy/WFAYOyE0uuXfUOht2vOBLESZObnCJGmADhVTP5n9NNl1ogRH
HJTD6TlF0LzurIjUx396iV0/J4vl1FqgQuJNakWc62ujd/vSfwFL85nHd7jLWRDi
dItRLKYBdax48NZSnpBcHBPL4eThsT44S+u8TKrE9e0m7cDSvPq61WjUKebzHOeX
MpLY6bybJ67N3ACeYHw1gSSUJQVirrlHQ53EgO3OsB+t3HGZZ/cQz4MftyyatC2Y
ZKdsUnSSfpfqvqagAlN6y+qbqad0hK0el0iR/77jNNWpAJJBSOckm6UJL39/UwPB
rbxmBD9ARvxP39FORndn6ADuQgEzM4xOQMeJtWg51NzYyVOhbAkmib7lXRsHHwaV
lfTlQLZK9R9zuQfJm5w3ijul4D4EAL7uzVkonkEtX+J+9mfKr5BaHGuFpm/2NmUf
xr7+b9ga0K46F1SsxUIQZwOfC/Hcodltxo/N9bwyUq6dg++vTNUnyMjtQ4BSXoI+
PFzXL+7H2Igo4hZOJTrbMlEJ6ZJtNF2kWxhaNFXtlyQ1oTlU0ld+Hvpd5KKB4KsF
e37viRrwq4lc+PpfcGt4POo9EagLegLwlijXrXBylgcCUJpUFf7tktfx+H8YN60f
PvIxdJ6Od0OLFdaJbE6TsBQqZ0DiGqDVdZJX7IdcFP2GPWshr1D50P3XMtuopfLt
jwgVf8L2IFsBHG0OQe/0ZGdeUvmrpKcCMiyEQMICw0nS+Ib+X6fT5U4SuB4KTKdc
WyFOaV6uYlrVSnkBQwLdbbNh+/PJfT1Her49baTeRVZIicRwk0vIU3SX65QO923d
A4kuIM7y91q0DEL5LkMT9Qw9puniEPvCIUCe2u9mfxCzvop+YDEbeAOuASfkjNtw
gmx98bfTNate8GFynXHhasbDn9Atzw5Ms0NPH87gEkhSYWieIeeyvRrnUMIj1wub
QQVdsGVZU4RqQ6nfwP7yDgTMZsHoFRILolU+YYOBbgbiKfQXNBBK3VEN6MqMbPXP
tKF6mGqCE8+12h0lTOi8IONHhHfts8eUpAtbI4joyAku9evh9wa35ZZKdnaYcBgL
5ToGMNMtuASRXCdy6sv8F44TG7V8tXJLIVKejI8dlTyuOJfYj68AfQ7m4D/a+joa
pS45ijimAjjERvvvBQOJYHzjbfB38sU8pX1EqSNEtgCCk+vO1RVrEurlQxCKaSgO
zEZqMpbF8IUUKAAfjWz3V9avMPwOfGilIvqDuhZeA7WQrQc9rR1LZpPScKznjdxZ
B7HKxEWhX944WJDtT2BX3P8QJB0wqjLZA1eytCVp0gqxYOV8nO4v7PGHHAe6qi9u
DT2sjtT7MnFjnC1v/wCYZOUTw75TEPe4c7xXKUX7rdvSd3HI03O4QoWTb8px2cC6
QJfFSEJ/FqdAnQRW7El3SmzbnnCwCjlFP6ojbNE9VUqE2AnPyJ09rUOjN+WuSdUX
9EpFemX520sIW0XhM5J1176iJaayaWCjhO2XnM6NQpVrpf5J+BQlBU9eomMn1Uwa
4Eh+HAWaJqfpFliAgId1jP3cYBXL6Oc8aj25w20B39JrbB/7BDrUiSCnmhS31pvS
7jEnizxh0HbYXeMyvYbPBhOuauQIaZ+qNhhoOHiRxxcKfc6WoE33WlEZLczTjA4g
S6JPxV9E7+M576L9S9gXjzrXxBn7ldbYuRim4cjtjKGmLUcDNI4bKi7gulWDhw/l
oOvs/hgePcNy7HPjRY6cgZQBG/qGHzc5zdtB3EYCkp4CVM700EOmWu+p1aOih5K6
dI90ija3WIj7kkn01xWwUuzOvcSAbil4HRm8qsjXpW8UFJ2BtGGhRxQrpTSgAybs
t9s2tn87aPu296M/jiMrBZx9XpEXTuvmHvxyoSIyJzsY4Cz6SlASraisLtd9ZHAZ
fHHwHXUnEOhNr1ZzoFMg2j+4Ymn2AwWbwwEunbsvvfzLB+F9DwueoI2NRXEh0x8m
hxqrXmIzM3BOnEPr2tiADjVvxgkGYdhLZ4DaJnkVl5UUKZIu9C4Wt4/IaW+1jE8N
St2nHp49wclkGBu16ysaQiLvo1mwCYfrRISbrBgs2kqJIiYwUtSr+ZQX+qk26EL5
DnRcyV52Ag1tMpQ/iaY+1ueQMvyOI1EwwXkrJPmwJS+Q3JWSFnCuD7ZZMRYbJi/8
CkFl48//FJLTxMahb1SJq0+fWr1nwyZc9QbIv8n5KtPrZ9dlwutDKqDHOiXYSIDs
9moQe3JeroGfuzLQRBG3HCsTvTVcxw5ynTSblhMPeQf5WY7iOGd6iN2i9CbE3g7W
elPxax/bl38JerrR9CrXghMnr5TcZkZ13l9AZjjUyoOflCiseR/f7qmXnHaCgF3p
QwpNjqpeL8oWKxh3wdAgVOF6Tdl4P/MYroUYRxFi++9sTSwy6ZPP420v3w0kaWKS
3TrZ2W0deew/16VXrrjhPjvs7Plk32THFg6CP0E48VJUQEJNkcub4ETPJy5Cl7un
LAGY2F0yovMiARvgOENLQ6TY+S9UoSiSYAZGKmO31CcIUZiGTqHMbwHnuxfVQF1i
Tbw9JrvgAuoNsMtELDLZDXAsIoBfxNv7UGQanvOyzEvCgNZ/Oxc2ZhVg9LkM/RCF
H8J5Uc3SvtS9zJcFnEGYt/q8fyg680cB+u+NeRjK89jpemlcOdAe9eQD5iRMwoZp
whivyyHmLAfVKa+yCHACUcn92sB/NF8t/5Awcq9wnxmeTvWVFWX4B8C3A5GOqnW4
0KacxYsRNxsbZuTEyhpZ+FAJgsFvgCCcr6BVniqpm7jpJMaTSUayOcFcjElZR4k3
bj5jMC5hm2MlDOtS9lj65jTkpWSOkh4hyKAGt5fGk95DlplznWz5MzqNEdXaw718
mPqDzvfkbU8LCc4gqz7wZVhP9jpr2DwgI/G2QA36GeCbxnRxpC8+PVjxgUpG801z
SUuIqC2Gyou8Up8v2QsSvO1ojTGAhFVel/83dRslp6qzoF/xzKZeSGa7r3mP2tUM
m7WNc4FyvFejbSvWWVftb6yKdXnxLOwXda7ERGBmze+b01m3mG9qoQQreJ14AIva
k7un2Kj77p2TzrdhcaC0G8XXs3R/yA7eAnL++pT3VI+hW1scGNPG1hkbbpjE+62v
gpSiZtrk1CsIUZgWfAzEfuz+MK9f5oTSOuv0S3mX/s701iq103vzhLnLtUsuuBkO
Rl+W5FBv1vdWTbrcTufS6qA7im2oABwq/f9MtBvfX+vyKGp+V0ELI4zSpyMpcwZn
rdMJOgf5MMqH3f4v+0ntWtO6v6FvKLCyQSPXW0tdnJycWoeOI4VsCExeiLwhU33I
AhjKsKU62NC+jBf6aC10gacWixbN3FP41QlQL/Y4HxJo5Ig0gAzDI4vGVdpUYTCe
YXhavxRTzrNi8iNun00pq2xHhfDc3cdXOzLS+ZVRkxN4YJYTMnPLYpOQjQuVd4Ej
D5np9ZM++sgIEGslZoxbryZAofoma+n6AaqLxj+D8ba05lhLIUpoWKBMAlyzYiUm
px9J5KDgkrpALm2KgutwCBco7RUItTrnIWR9Zb0uwhyeeyC5H8tdU++f2FneRL9x
pmDiubrhZjLS5iBJQHxNKvfcvqzOHumRvpgmKElrBHkCkIEJEaalWdTd4ruo0Wam
a7JBmCz0jEUlBh68nH6alfFhu9Qk027Hh6UiqLUsqJ0Uhi3C6b2lsdGw4mVdc4AY
rzyob79hC814oDWhXS7rbV8t0ECt6U7mX/E6vVOXI38ReOX5ozGD/6ukZ+oodFF4
udwnzzaSyYXANHLr7fi4G2KgPhSjcLtEd/CZ8y3S6voOr3Pb3I+bIOy2rbN0A154
I8zs7kMM9ZB1DQidgUA93MPJLGuA22w8B+XOBdg9pzYuOPZ1YvuiIEpbmS425VDD
dXgVkixa/P8CHCtSK5C8a8wc7sXV8I3cnddsp5oArl2HGzJKq623/8AFv0Il4e/5
L6ARGgAuAglcUG3HP3ZFgPz6M2gO1fmXFHlU+/ye3k0AKVUTHoFdBMWQ9182p4j7
5mRz+hWlSMHWQoZv6wzb5N7p7+cD7plrhrnQbVqIIUBvSsqB1/rFFnR08ixUZFky
hXsUjYPvvvoA6lgjjtuiKIF2qXG9SlneVL2kVFkE5zYXlJpLoJzfRpir+UIg9eV5
Ct0jnPk4DMvyAavgoqnq/D4CnUo5Meh0ZKd+eEJYpbNJk+vPlJ3qF4SSrn1N5TKs
IIHCZyRs4v0V/ZplRvCzfgX0tmbhT7+l7D4Ys9pTbdvpb7OTT3C2iDio2sk0vlHQ
a2Bs+DuddtAmvzJzZxaCEiU8FiW6GIGhpGrwS9hc1qyghkCg4PATuS/PkFzA6IBz
bz6FyldODhnvThThF2PsJFDu1e5hCAgycvOkpDyM7UEfb05n7LgNYcPRNP6Zw+E1
pdnJEiwQCR4JeHHNsbHoonAPFOYbf3zHuScKNNQME5J7s7TyNywb7k4f8WkOXTaf
yhhJ2SugolgM0x+e9LKkcV/5X6BvafZljtw5AL0+5Cdyd9qafhYIbOSe+tbCo8B9
9ldEfp/oJEqOl4h91cp2IipRwSqhppRTBQioFiCgjyXBolI+4Gpywe86cjA5GlBf
VRK7lq/3TZJ6hzEth2VghEP+JxCRG2HluxHK8Tj6kdkiYok4+p5/POJy48h7rj4s
M/XMGA2XslOJKJTIlyoAV0rAzGRsSG8JKD5AF83MoprEqeZDeDFPTyS/4Uf2T2q5
XK0wzDPGa9eWO6p0aIHFG8bDYUwLcoOB7EwD3IBqn7Uh1/1pIzUxzewbpu/rYus2
BjEZQuioOJwtP/+j42S4Y+GFJ9W9p9RtmEa2jlK/B3OA8j36+L0KDtq4gdNBIzhK
t2v9UByn+u8V+tyc1wJw52eP873BoB1w5n7gjATDYwLn/9gLAiUrNahDOSnfwtK0
uqimpCPmtoKX3Aa/D8OeBKNUvqh24quE/M0MfjE25zsAOSO9kmvtaN1FxEpqXBCP
QLKNwt3j+kkZRPD02wTX9AbQ0JncNm9ENwBXVn9zKeL51xJcsW+2wEW7y/4neb6s
K5iUQrItRY41Q1N6k1wR5sjY+55vkKPty+t66nMSSI6iTgOdwemuYGzDH5hmm3nH
hchFGN7VFRVZ78W3nyALq/CHIpaDK0pLwDtxtLweX/7HJWbH+y4K1boL/um/dBoN
3rskPLxug4cZ8ybKbaZsV33AE4wt8thKc8+uLhpl/Z71VqEWdAorKoxliPyqowia
EibDjD5hKAqqnfbS5B42GXEjOvGaZWri9+9nDtcegO9BgJpPGHEUEd3CWH4M29sG
wPtZZzCuWcEqxQYyR98+Vgp32QgRijuMxnrLTAbZSXANQslFR/J0UioqPaSOvqFi
dIlKvaus5LbAKvdZ/W6dF8Nu3IXXNKDb7Zek7FghNkaIy9zPEijNoQtX2sl10pq+
xXyQtHi4fo5Zo69qWhX3Dl86mUhyPKg10uIcvYXLpGJ350NiKncJjXRC7yGR6MGQ
75JL0OrFaK0uKbbIv1uoEDkOjSAalbsKZpVooUF1eYhzgI9kYWir4VLl0dGfIMtN
mq+yx/C9EkNnWPH+wkEEFL0uYccR2cGOjzUke0J0j0MSPwoGzzrznQ9Rn07TfPMd
3n9Vpya//WLP8/eEl3ooWHE0HAVYjnMaD1S4/BYw+Lb3RfaG69RR6LeYLW9VfnL/
E91GCkOwnHLPn645twEuWasDkwwotEiSaiZKrDbw+qTZO5yEQYZG//spW4wB097g
U2ZrIXKIPJ242EYktCwN15LO44nnYfpdK8R/qdbH8tyqkO2QjR2iJfKjXf2ZrStP
j8KZNpHaPj92R02ji36maI57wTZ+kDu2SEetm7ByRb6+3Xk2PA0Y+LH9IpbiXZ3x
81ZcsWpolSBwF9Q12dAl+J/UpxGkN1gTOem4ILmmmHWnf2+fY9deotw+HqJ/er0j
tc4h4inxliK7BCY98QleGThy2jnbn9PJjSqpgeHiTj90ds0Ms6V+BAuluwMtsQwl
iCEfFPw5zQIM9Z0vbZWzXL5kFoQye0vrsh8LuPgDUh4NZbtQ5palNpLhDy1t6RS+
oXLPCgM9q6IC51DISBhcg91NfZ0tI7mjug5NVYT2fZva7CXjFVi8gPXt2jYyYBei
XCI0JyBcSzAL5xLQEK5YLBmAo5JGLW7nsGSp1sPvaInIQCJWkY6Ibo5nlMiDNHCb
alpuAszSSu/hQtXFdGEI2Y871QfRUzT70wqC/i5O1un9h55duEttWL/oB5YYphg6
z2mC+tcMJA83cBfADcdzuD1Sc7nbHCrwmmnrGoerasnCExVaAGaH+Ya9iLOACnrX
+VJfI2ABa/gqmeXAehykqRwY6uqpoykZyH9cjC14YKJ/dcXqF5s/PTbh6IGNLAqF
Xj6Y+35dcjvXqDxkSw5qtFkjtB+LUJ1jmdeJ8oqhxPHJM2i+sdR/u7YPRNh2Ir5y
3dvKRupaAX8u8BKsjX/UBF4SX5T3BFRMQsn0Hp9W8BC8SsaRcF5rxa/lDWhIyJYh
yGmN/TZefj6FZ1TiTGP6aQPtySDBvoEaNh/ZymnzTu1c40+MVCN5hfhrujpXkSel
6A2zU4eIOq0hZEBeapF52Td/gCPHXMEPcfXQFIjn9HGvcgIFP/FwTmsyoyHruKoC
tcQlOe419cv1zfKYjiFPRpVSXbUxVZ+3gQit7W9fLrO+AcsZxbjyWHtTlacDnedv
RiAMELn5LYT7gT2uQtUnrbgF+UZu/LrIWUgUiYPvA5VvG1hGLejGtw0/a2myaj8e
6KFgseSrjH/LgXYJFOAgP9QqegwnevgJjqo1ZtzKNUVw3cxZLU38VOno02jM/SH+
QQVOmfP/qyWU7acIDtsXAo+ScIDzJqvJyJW9gdyJh7C/AXd1/XMglXNgtCqCwYh6
yX/MezcXvWy4BRO3ib8dcr66utUIb1rez0osArwBUxaf2ton5lvPuDYfVG3wjMV8
zzAfZL/28wI1Z1QHLBEvaGywoIewnnE/i8JxQ3FDuhDwJQ4q3o591BlHpfNtUcG7
LjNqUzgXHQsJjH4iVhSqhgFwXg9CudlzcUnHoOgExyvvD47mYKu9Q0/H1hh0l1Xb
jZT86UVJaYF5KXpkA2Ygjke9wHn61JOk4d9IhNJey+8EM9cDPm9taFbp4Z/Sc5K/
4n1WKS3BBFrrzpCXPiCWqxEBwgqHzC/N4QOMMqpoN3WSdvNIsZhP8U+QISYrLKGy
S6aZYRLd8RQBbNx6vMh8U0/9m/06tKM8sFp6j3ilS9zTOZy9TbYdwqk/Bwog/PrD
B6DX0pUeTWUa5QWLo+3hZyY04U3lLgPIuR0Fk418FjflXDCZZxaqbtxQ9RZ5kSib
Y3a4AaGmU8b8At4C/Yfn4AkW4YsHflW7dEjFOBhJZ8JPSIDndg+3UUwdliJsqKdH
tpTAf9cjt5FHsKR2XNcDoCImqT8oshWECR+NHaKNqjQHf1qtVeHtNbMjqu8QE0G+
+RMZeOstCwPTHVyDL7JTbY9AAPY/AiM6wf3IA7U5uz4N+MQIl4o7T+52qxB761xB
DEomj9u/0v0sHE+l1q6nnSG2V7SoeZmAZRXTRyQh1cUlFBs86qHA0bZJ6QharDYH
Wc6VACULTFr+NGpXjnbAyvgT9akNl0rbvDmHiqvxoF8F1FwHmQI+58Fn8je0UBfh
2xQE8S5CN3Ju/QNemH9h3nmcW3i5SDSil1q7sDDuQ2UNiw6Dev2jww/hyD0RinAk
uawzioPuQJeUzRtXvowTEp8+745mVsrF6j76Cl2wrRH36gTNY2KCpNQC18HOAD+y
PSSWE1jIwpyu5Bh08eOglZtIpGtRmmoCFP4/lsr0CR2ECxkaXO+CEzCDoEKwvcTn
rW5Vy9gSuvjsAY7yeILe1tAo0MBJ53JP1ATovP+DZYe1S/NYNbDUPjChABQoTn1q
HLPTVqWe78MnVTEzSsSq4Lyj4aOusAJ/Nyc7afWcS8XBBOElMSC4t0Yo1z3As2M6
u9GOdOx9qRZbQGSlRRTbmbyCO8/9dLSvzhADh2YzgHlUVJWAVALw/bJURTZAQL6x
qKPbKdtNtNE0YROlPshyODi1vbIfiZKE5EoH6fnEsUmWj2e+kHJLd1N4Ba7EmzuD
0ZhILKIGtTp5dKwDa+lLF9zfW8qCDKqfH7/ZESuxwS33FGX0LHSCDCM4emmtR1pb
ROuJamol/QKaivyHj4yD1095q/PJZAbvC175BHBcbJhI62oRFgIMBUKTfuC3TuGx
F6NXUdNmq4uhoNrC5Om8xUk0FuvMO8YYjHAcOCCVT6o1FxY8aIs8+AKbVFz+pxal
okx7xowy1mJnoFPUwKSFU93shNvpMMsB5vR1I7sRDc4kK4tOv0DnabZPNvZ2JqpO
1HLzJQY5dAzsu7qBc8uXOV5sGss5S8mZ6fB9iRftqeq2pQkGEd/M4RPKm9mDBmIB
OXVWHr4eyCNhsnh9W1KM/b2xYC9yeBk2IhrDsV/O4ZrS3XisFRRGnaEbTLQCGaiv
IJPXVXNPtOBndgHKS8CBek2dvvb1xiZi9B2eMB2DjUJUVMXdSTHk6IrgRyFJQdeg
jC7t1zPhJWAYMp2gSUCnwwNUYzBzG5w4hfk3i+MTNgBFHJQF1vj7I6hSaJr6o845
nCdoPLBFQ2RkUbssNQgu4eeJ0RdghP3Hee7dUYxZb8LLwDzmiUDDvJqpk0p88cbF
W/k0YIsbTjepebeeQwSndXqohMYHyFoahcs6O6AErZpidAEh4jWyJLMv6qYTqVYQ
OWyBGn+XhBG5jkCYWbcgzthlNqQ8FSD507WV98UhX/jxcWqju7hsXOQjt07K5k44
RlAzDxCVrW4+WPkN4sZmEAdGH2nTggwmKwV+W+QCG930W8sK1dUzWiDNa9A//w8/
UWSih+OOn4l6B4S1BhaIIucl3YbW8TDtZfolq8RAt9qvPMxcofRuuoAoWGmowV27
FT762xLXz/PPZbJ4hd64gM+ETGCxtqw2nAxR2MO+qUEQMhjlejth0S/MyS6rXIJG
C1R3kf1E5PT6whSxq/CBwIIZWYnYDojiqwFBxQC9Dcxxred1fSlPzjsPkbeyJXpb
BPlgAU3QtPPQW2UZiMjxds8szUK3OOfT5YztW4T4WrH+waKiB3lTdbLHjfnCQEvy
5ulnuHA62WHsxfFL3CjI7065q+Fvyhb6OPw64HFzyZu+X28CA0gBPN9laMxvT3nk
uR8fM/IPQzZMYgRoz+Aj22hSX/9GbC9g77tikz8pMUBgTYLoiAuOuf1kmAFgd+pe
xNgRGs8LjaiE47vg1DcVScTkwITur2dDLIHmFc80uj5X00InrRno63Sz5etgQYYd
oDzKd4uJDQlr1FEhaZvSVb2ffX8OCUc7fCSdynvP+SJdSofLS5lqqYF0dz6kzD7O
4K6lxi9gInEc2J7pmKFknEEnUI8UN5UUlOJFJu2mfpjejY3Yyqyc3rptNsV99dW/
LttLt7cWfDWvQPUawjFgTbgv30H9hAlPZ9X4eeZjUFaachhTbygMPMiCbUtQFry8
ZtIoQo2fJpfFXx9CGrspOs5AsS0JYhQHzcvLmkNxUXW/nmrptJEs7AcvO6WBdhXB
ygpqLHdksF6WWOjGkOC032P8vGq9WZNlWB+NWXaA0u+zZIiLQyKgAlERI11/Ge5c
KSd1EEpkORDlrKYOsYPgzHX2QzcFGWbCScVOSrQV538wH8Q8r53QcCPsmw1JCWEp
XUfeIR6IfQrNNGN5XjbZSQFYKjr5ticdE4AAe4xifjqGTX+tU/UeLBZdts5hzItc
sWRFUxztn0XUgvtALsgOFTdGebPkyVYeM0snPF5IXMyGGqToAvqfP1uCGwKjLJLa
oXYUP8LhW2oYPNdPDOxbrv7gnqpj7WaMYopVvWrafhf/VeHGAlUwpxcVphQDDE/c
r41BeS4/VVQW3t/thspabvbNEjcPJ4vdauhF8lqZtMAj+nyPWfeypvJJPZk/UTp5
drG91pOp3VJDAUcM7i/5FHwiHh0PMiWnTjFidla09hye2BUk5PIFLgDhxgkaOfrl
kudl4seeM6IRaP00lFwTNGgWABuDDlCDTTcBV1WAOM1B42+Z0HI/FD0Nc9Jaobf1
hmiA1yZBTKLcu1I5xpcxwNmQBcn4TD67lvNBLLP8aOXUhsTvqhpvycbBGmIAU5up
zVEcEHp+/pWMELYd+K+AKNl3eAuhFXp7wErKOe9acM1PLkBwv4oOMwstmxLQ9Ed8
iZru09fnevn5UVCrzMjPCJib/vNKYEd8wOD/tnNbzUQatbEIju9GzJT4xSJHVKdr
E6lQlyTYjKVb56MgekUQkBeVMdmZtkpIAkgGQyCZ2asNNwbGXfPTrsP04Ep3bIq4
b5lL+KhOSoJgAgJs+GmYtdWdwf5ZSgAN7qEwunqKOzT2Yw0tPUdaxowgJ6d+HX/0
2sUqucBeLP5vDZdgfliVSwSgiqlT6EWVi51/q4tAsN7r5y3tn1QaJXSyMeKelMtG
Qd/vEKJqO7O0NoGQyaEHJV6WZVepxGMK+tSAOFQGPrDKx/VizNM6oZQQc3Q/5N95
WtqWkU0XTrKjy+/8msmEkRGJSN/xhadTWDd96Yw6kNmkurU99bPbSYrmP3voMyF7
KoSBhsXWpQuJLTI72Gp4TZsLwd4Bk6Ktysnew/6lj5uAA5Nn2vl94KUwAQ0q9C4C
yod6ueCDq9hwnby2pYIs1+KgvCkh8DoHRGr1FscWM0n5FQU46rv0WCUqeVgv50Oj
X5w8pFLL7eFHsCDM9fCK7XBo+zpDXgRPJtvdPX1NaxtP9rWHKjdrOEzXWa7YtdE/
egqv+gMNahi0IsU7nOGTFf9GDwzaJNgRiIYauz0qpZR5lIPpGs9NcT5rjdc52qax
jCrPow3uFo4srrVkm3Xd1d072Kcn195eDSUmoplmTSI82g+gQUwds6OPZ12IdHaU
madYHezpA5unS47AqlR7qwhz7lK+wowCvH9fNKfjrokrsOlQH5BVjX65wYggeK8l
ThTcVCv5yDkca1NmEeEBS93L/r31AqW4It4yiRsXJP7FJghmu6uGQlGVrTFVAR7a
NDI0bP4uQsBbf6ei8/HbSebHEgcPHNXNf6dolai0jlgjXOdUt85z7zNGFFd6KqRu
5IUnNVv9bLinPkNAMEO7cNarm4MU5Rr4CB5YIrT9ZmuAbs0tFPRPLOUgWZuRNKTl
IfMvrmHbBUQ0HzRnbYqwnhvOfvZVOyElH9VeBvewxMJr6sJ6zi/I124htx6uIJpN
NaGRyeWrjI4LXeGsz73CHs7Pz4DyA1fETs4/EGNYNH79vZT1n5HRwWseytxBjL6W
7X4xuwSZMd2WtGgNHPluPqOFcOt1P7dryncOrNyLtcXwjhIaBMHuYcWA5EBAeEIQ
7vrwMIQNMxNwLGWwGWaN+GgVoK5TafQ59+hbl/SR9iXreuMztQn1GJEX5qOUpAhN
zNN03I5Gy3eXDcrBfpu2jPyI+snjjrCSNcFbSxxC6cegdRzAeG1iTskfghFHWUd7
sB6LA57oMnUryqqEaLRukxCNMy/VcH9MITZnp8UcJTG0cYJ2svRwYXgDctdB0Gkd
3d22kyVvsRZkobOPQKEFj6XMrRmtmmSv09KT+1Ddj9uSaXa3bDwAOX3VEPBrTfyy
i7PmgoUy+BycS5ApXQE0ex3GaKd/Safuobxt3IKqHN/YeJo5nIXX+IdJxOsxzkBd
gF7/6Ir0skVuVXlwisX0w1IGimTeFupWItn+uNWy3ZlqcumZk/y8F7Q/AM5gKs+l
wfIW+YRo4jLW5Hfj+UkH8GAX+3JVfBxMa+baYELCy3f6Wkezj97dH2YSa0vLr4cV
SsNnxWIyeMstXneKiWl62c2birYXRmZI/E5qMHBGWUeTgPsjaoQaRDZyO5VUw0uP
8VomtZbDbVBhxKD15PXNYfTsusYcVbHCh+knR4Vv2f+qfJ23cMmZZ2jf3mpLVRvI
YvIUuigLbm5kJBNsJ6odK2GpuBJsNAm+O/p82KFzAVw2HBzQlX3Zs1+o5cB13at5
a6W4Tf1fk3ptimomvwhMv9wMBTmNoRYUQPIYm1qoIByB0VHMGI9IMcmyxrq46CVl
WPhzzCPhzXCdkorem+VZndfXEVK8EaINRzyZ1Y4fCSU+vEspKQr/vWmfThhU/0lv
hBIDLL+vPhFLISpWkL1RSxmPp+E6kNY4Dt2gJcIVKK/4U1vMr/7n9hOi/6gFQRUD
A5DGZUooHFDaVowowSqbXDSnHBuk/zBEKmIvNYGHgbzS8JNXbV728Z71Vd+furpu
AdQOeoqor2MzZdjA6QGr4gTMIPef/HZM8EpEakyWz4IdHD49At/7sA/k7JPcUibX
VkO4a6Y1fPNWpYBMuPdmuq8e3/v5gtBgIy4YNkp9WPacfZzzjl0hccYJfuXBe68o
y5yLQb1R1965mU+eWZNrrfXWUJqdyiNPgtKNRQ8HneYiqS+1aUN6kXf0uRz3X1tM
9s1NUBpKxXbg9TZCdcsBdbaDF2UaR3bApYdXmyxz7p0MpZKLFDVXXwwA/nSWekoz
e4yt4iWderOCJ5zPvp4jxvNAnjIYtGUfxPePJlj5XicUuNz6HtreAm4JzFVZiFJR
2QY43HfMNiqT6DviOmNxU758JlZG/C4lj/e94it8bZdSerykntJQ++GUmJCjq+nX
WyyGECkf+AkF1IG4DHxqROk75dWTEMZf4ezdkZ3enafb9wUI3fjdqM6W+yI6X0lr
77ulK6XUtnHYqMZUyFrIkIUlfRdU6UHRMBHB8HmcT9wk24Aibf4OcfWTx5mdoTN6
0Y6caod5F94HUbT4MJP/3ITUpy+yDPL5ISDLPXgkmWrpDh3hWBhVSHQp4RczTAzg
QVZ6WYrWzEYMddHzYt7lDkFD/g/rV6ITylZK4EBuCGs/LiH55VobOdxvl5XxEUpg
gL1IDPTtOxIYH9Qlu4eKDX1n1DDguvLTctThqUh33Y1A3gkM1ATUrHHycqhNyg3u
2RUGyFnV/b0hNrOOMb8xcuag4XVfDSjNKjBbQeGgrQcSkRMiY/XEZB2AM7djHsMw
Ay7h926Z2f2uDZl8whOoFil0sXd+h5r9qZVD46jfUZg/dFjRe0Fe0+fzGu0+ugH4
c97rK5HyTFTYQccZuLIAsYxR587UXULHjZIoe+4u1qlzmUbQUJGTw5Erb4Lra3U2
8irIdX1wNRldstrV2N8WF6WFNvlNk18qUAUU+xDR5FJ1xLSHNEjHFgUudKFGQdVK
EDI84B+WHQRXZd6z1v+7fccvDIbjYyOs3AU4aYz40UJaoeh+dPGNiQGDumu6lzvX
H5MOJxQQLr7Ey1lVxB3vhRj3QaSLZTVoH4T3uCZV/fIL7Zztj66oQ9tPUzm3PoxX
lFnP6RifeQlG0UnYsAtR1buhF13cwGEdtUFNXISc1x2BSimk4lj0hLRVor9ML4RK
eQmZRM0zkcju3/TZIeSxbB7yhjymn3vfD3JQWmpsKdsXkgBBK/WZJAvCrlTNewUq
AeAWHxECNZ8chFWXgMExa41WumdPuMeejj1gT2xhiRKi2dQV20cXleZFrBY3/dBH
Faj/g0EBEZquOSlx16Cqhz5eZgkapGjqtnADByzFu5jgzgoL5KnohaZ/DC6enjXp
kQ35XLzL7fQOIyxt9uIkqYnJ0DS8vN85NMdand2X6BOexQo5dHqS2TuPsc4Un/QF
PySh6HPCVXHp/5gFHqaUecm71PMeE5KUFP/XFrZ5073hZUDD/0s2oL7Dt4nCVaDd
0wnHeq4DfAHUxZqNlkmTahaWIuSl4ikQFlWDVNgcxv3vTuPr0AO0cBhMfjTeSrF8
s6xMIK4b76N3R74K/VtiOAOYabUES+fEce+TLgd8LqUwAVoVlrqgUq8GVWzEqujx
0xR57v2o3w3VoimAuqigj8HZdUt7AYldYztCrG6e0S+obSduE8/gHm7zd49KHmCx
5x1ATl4pMTdvzSrsB5glOhAf1NjBXiItn9cKk2p6PWBNPMfxS/JduzBFOCzrjlhg
THu0fhVvmx/4tVp8EMfKR7cOVvn7VMSE+uDzotXHqNoy4XiylXS3zY2o2DLRJ01m
I+aLsUE3XBHrMBN0NwAcIPYiL+nU0LHMDsx7OpkNihLbxyHrHxy+bydJscI19c+n
XxLTMVJaJL8RyZCHPKrzdqv6Fb38SFGFf9HypwPTRjZ+sA24in6p/RGbRpdYMYXW
i0+Tyv9gVLe+oItY1BK2TMTgsLugUlcwLkU0czFcFswDFuAUAIaehULGqtoaW8Fp
cGr636wfB1SlrFlwblB2MBRTbMGUx1tQM9outf/6vlcFNZv6z3YFMX+AgwQKkZih
sb0IgG95bc7B9+K2RqYK3/JCAZrDWszkn1Xg2W2k6UQSCS+BGX317hP66VeWrUYS
a5SDqwL0x+ebk+Es2Y0J+FGJT5gDLreoxcrEXvEWpPgxLI9BF16wFCUJgcrrQ2ew
rGrAT0VpDEnacXPzBNlKh/7I8zd4C4W3e48hqu7nK4ARJPUhCg0akEYYJbYmeytH
7cC26oqAXb8Jwe0+p+M4giDsi20BlSHhIrda94IUpGnK9eAwsd82Lw4d+bALR9pJ
amn2dUCVjXkI6+tcOLVyG/fLgL0DoRKaPWTmtgCOmiSi7rA6RgMjlPO0jQtNqOaE
HgZ0uIQVCWKz/hMhhTmixL1Q8G2FvXod5k7JQXAt3V20G+zkHThlnfwFHCXsi7h4
7AFnxofkMvd3eXClq2Lm369sJWQEMSgz4ZBhQUouxE8nPchRa8l+cdKOiWA9hQwh
Gx+SMBPcy8p2vYf4Y+hUlgtMliC0jDVFl0vhWUX4OBpBY91e0ZHLyFqbvp8pPiEW
ZZOKpUfuNR9a2ViWBou8GiN92qyzYMqr4ZXOfSmPYaceu7LlrpiFBSdh44EGiult
Z8dJX6rb9VUsw+58puQzjuEAl9Vn3KP7JedUNAv+BS3Hqbsfql3EUiRHfryCLAxu
cd8PDAeEvyZvywj+piZDIwrbVa/n5xNgq8He3vgFMKRttNbxDX0UEZX9tVDfhqJ/
57Gt3MaTdrtIXkrzfQO19ppnl+L7J+CgRouf7pvEmfMPR/V8wCs7FP4q5l0X6sze
U+cmWMT8sjH4W/bcH15GGIMe0YKFKIhNJ7dCvl3K5ISoMj/X7Y7q1qDIFEKRjNrA
XteeJ+L6DpT5nlKovc/jYDeEWL6f1NypXPR0LZ98UiR3W+n4z1NIjl9xTgBENVZB
NYA1bKteHsoTRgSALW6qfvzjywYZYiCmnFPxFBC7Mo+mnHZdjO1coySfRKOdpI6b
GWFXWvxhlJ0pnau3+/SqfQddbxsdw3mEFqwe9ERzTsCv9+mVLq69jbrtzJuLpow8
UDCIckRnWAQybEwhstEQGvxKgyIPoqfGq3vcAzjrNpYeJi1Xe1W5nZhyguQ90GTT
cP63rOyy0jf03++6to7lKV1NyEchGmTEeSnS1Yz6wmWJocXS+0eJ7v/GCmvTHKlw
kwqsOlVrcMmGfk6cPvnUvJStvEHQcYExdsRSWNNjFzrqtQXonIf0PeNA1ursoCcP
nDJumv2pJFQZ13BTN0EfKeAqoGhT7bjgiIl7Bi6vdLLALjQ1jF4ETcFiPU5iKGMk
STahTX8j4vCXPrxJRVKZkMq7RXzvE09dc+cUMGQ1SW7744At/LCwEX6ukogb+VAr
LeDaBGUJ9+IHQQQcmIkhkN/oZwadfpK4t2WlUX0dfMSAuVwVHMwQKpovmdzs8qqt
F9EhV7UzIHXH+AHTHzWNGbmpGwPK5HjU0K5E0AHa2WTLKgLiuwhDTZkdRECJ5wKE
gUpRH0060VlxpAZr412ktsz+RJm9cVtq8C86JXBRICtj5AU72nUIHk6z5BqfvmIk
kTlA+W8yFaqpvmM1q94sdJC6bi3PZgY2yaLRL8sgp1U2tUw79GQU/BsLxnI41KOB
pbXs1gpJuIq7V20QHGO/68ucbStNfMUDkqizevmxzTGOwni/R49OrmUJa+W7zE3u
OgFGhNH2dyF71YWv1+essC0XAQHdWSjLIPmr5VF9ZNgGsfCTFfemj7Ze5PenO1GQ
uY3bO0Yj2/FCGElSJuVqmVxVNl0fr4UsHE0ufXPSzOlRhlXFYPVPIMaUM0/m/zau
h6T9ZDZEqDy4WtBZ9BPyN9c2awFFxRDpZtnuC0u0cStM7sT0j3S6ExbfxEzy+S9T
JU3CTGBfXZ699b7JatStJ9aJqdyBwaFt+yTRRyQ3kn5ZrcTnFfuxVaEfI/KLg29f
hyZQx8xw8iRZ3kzdsT1H7sCPeedC1r4fz4TuiFY6zfSYA7zSQwLcXxqBXaeQeV/i
Mtl+PMZKuORN2Nws0fo03RfJnwqpfKwd730zP1e1xAYubi13ueZeMXtkIMypF18M
YT4hgpNb16s2lZzxmI8d7gzixeZBWARtwaZ0teFtW/qmkYS64evtaz60L4lK0mij
xkkUWip3dHr6YohrcozYYkq7ScGrACPk7Kvpl0NmzyqXRNEQD9sqpHBQPsq2u+y/
FjGSPbFI/kJZh76qA+6qO6ADYX5VUunUVzD0hV3ONxT5/T8n6IfCJ8IQE4ZMmHiq
h2F0KY/0mTE2TStGUTScG27Yl/nnbTTj97YuLHd7LLBUpmsiDtKY2TXBKQ4ijm/8
gfwwt5vNEcbQMHkIihLuioYGlSDZdVG20Q8IB6ugi3qlYjo0sRp4K+iFfyaUvdiE
K6fODh9NX79ROVqxb+xrkhj4zxVSxQ8N+40khqMPpr6eDISrFJxBMXVYowM3UXOo
4NJE6+sNoZNhmTz9d6rhtrwPPX8J0ER099J+zYccCRVQGhptz/K+qzqKnmfQvges
PZfjqgGuUefLTSdXKNMBTne+4q+k8mcl4C/wvP8qxV2PeCJBdF58eqJhGMW7qkUo
4zAyaaGmabosWajKppUkR6wtjNHIib3P/nw0OOwJ3vsmVbFF97H8I+KMqnWKHD5h
qiTuJKHWnPt297JsCuTD/u9GKnmtEuc1rvL3mi4eANnstsc4l7P/FtVbjP34fJ9X
dIZmh8K2a+HD2SDfIp3NU7GFnqzsFnOq4f/W5y+/mXulFZYhW/Mxy/+iKxUkcFJg
BbjmIXnxVqETdc1/2BxDr6szYrRoHRsnBTtpJDHUuxT2Mtpqss3IfWAJa2SWRQ2J
oObmDaKzaLKU9KAtFvO6fBg+kUFHtGqihPYs+0HbXTEGUvCNRwq+APpdbjOfWpMZ
TDrUBMoMoXVeIdnv25sKJlqaaLzCZL88wcFFGzqJOrEs0IyomMV2FyKhMoZD1Sdi
Lzosr08sPIF98edpjyyYD1jZUqTGjMvpIQRftCi2ItxsszhbBC9cfe08L3qoHmZi
AoThrqq6YrwsEuPzfRKFONpt1AdqmRTWozJVdCgY05l4eRB5ZiEo9A+HUNctALry
jXEdrpGNAlrW1wcM3Dc41Gdq9pQSDRihjceIWXhk7MKh3DP8iXwngZ3lN8CjCS/K
3N8dTtYhftrxwn3bkkxHHIIH/qCsarP2nlwbdLp+BIZ1NkhdncsBj6xE9zfwqXDM
6zhs/e1un/Y7CHDJE33nmOvHi7cF95IO54/utH6niOMA8rzfeIrK50XCaoyP7ID1
kekh8mkAce+gXQdIw0sXDd4C13hN4z6YqqooknhvLEacwniG4yuRH+NRqcPvTYBI
qPLD6m/d49bXwwsgr5ZlkMqsF1mUYrbKWzuUXJENGp7QzAugTLS3hSNah4qtIbus
1tvdGUE+/q9NWhfE3q9Aai7OuKdliytAMrlSAhJuccmx1GDakuyeIyNdQo+UZKy8
f+uNsFhGNLhoZ5D+doU/Ot2i/ZqKBpvC116jjEM71G3fDD1xLZK0uVBQTlduXjeq
42HHjE4yPKHRs8AzjJTIIkYFyd98VpylcTb7CwEr07XZY9Z8XzqFjrXmjySDz3vn
TyaxQJLokI8oq4swa+sKKzhgqIwyvam1vSdhpaQBvRNrYFHXXWFKyZbOxZ9ssLyC
mbNk0Q93OXOXe5lj7kLF2Lgzln4QaIEovOtIum9w+4eHm4Fu/qLhUl/Jse5z2XPe
koXDOXitp/PJFKHeTA+OJtwO8hGRoVUv/CEnns39wNXG9rT4i65aGiVueU0A68+A
F1uftU0+5SAGqS5pOA2u8MFHWl066IVTgGTiA63txKAVfXvX+Y0Frsq858MMHxgN
6OpxMsa0zBEWVe44sfxi10XLlErFpRpvjDeV/zy6LSINdkJtIIYhww7kOi6NlyHh
Qml9pGplXL4bQ7XRuMdh3srG2EEFv5lRzolH+6YJuSxv1Do5DgUB4VCr4cpux8aL
UyXJhZYLIHSUxFCow/GUZlmeLRwxiEAxUmLbHgFhT3W/lkzmgmYSawGDmK74F2rl
p28m9ehM1TDPz9xQeLa3vzk4obHeYXLcXuehAV3wTMaPRUJ6VgHbtBFQSAB+5Zg6
Gob6SbKGq8BTO8l1d26vdeRKROiVJbb0rue24SxZ8zRD8l6vFC3uuWso144h5Dlp
UTvwQttMgnD/ux50rIhSoiDJisT4sLwC2UEb0gk1UsBwCJBmSOA5Bof85j9FW8f5
WOExV2F96AMJuuyUhVGpSxzCLK6JnP5yYvN0fextkskBWotJ6d/Ot9fUB5ems0W6
ctHs6c87y9w7xG/HA4E5RBmoHEo3grQUwms7Dtd0bpJk5Sklk65hEhSrZU7yVBDg
JUqQiF0OCXRzcpu43drEZ9FyGEG1NpGFfJAAIDdH476hrJ/1PmIya28anryrFkA6
eOfjnWbgsU0UdQJ2EsA0UN8ec7/eo8lO3f9I73wlNwJlROu2v9O7RexxbGz1rN/4
KZtBndonCYEgV5AVlLcRN1gnl6kA6pKbrjJNlqFLNl0nHXSBeLv9FNQOLt803J5D
muP56ioqtuhbIu94CwpRwfbWC44keLE/CKXTxXiqeYe2I6cpvtMDMTT/oa4SEvdN
o1ksGzjQI0CU79iMUnvDYWfY5zkwCqgk7lw7tAad57ki51nhw5TX0luviU6WscnP
cvhM6g+B/Yy/md44H/QGyV7ygw1aDdZEAFO/GKRZctf92rRlsXFUdSqIK6Fu19I1
dM3U+u+XvR2LDwwtBRnmFVPEY+b+FqMatOI8LwsSeE2TWeDamzmpVPWVcHgLeX0X
nrdZiPJ8htCynCvhySZY0q9Jdl+9DVmph6k950IfB91Sr2bhjKV+jJ7wZNyTIBFe
PpupXO2aZrBiHKg4SeVPx/JTp8yszZCZTU9XsNeiHLK+IR7UEbkTio7kXQHl9afO
vZmwjKPYglVnhDF1nSzj5YmiovVuLJ54o8dlQoF1TjuI/R9A3iswuNnLNV1l8XUs
IsJFzO+AX0J95uC7yFL6jYyTuap7kAXvw4cQ4cqzN0LxbnviuuPB3FzbEUXX9yLE
+PB7w5q21ag2uU7bHsyAI7xGtJbvNIHkYXAFURs/AUKZ6t6Jw8iM/A3YuNo7zsCm
tNnobynNvOSksjBZTzaW3kowoD2UX9dIvF1IpyV1hwSxZbDcsvBqLfEvQ2vqr5hk
Tuf2NFw8RgQyFOmh5X+lPClceEelYqu0tM3QGdMAzTkEDOmpyTmtqSL7ypQk+zK7
CbR8TmcOODuLz90+S5GLKaaGnwMsUHUKz18BeelfCbBcOklDveqFHGI1srscvsBw
VwZx8fN7b9JAiGea0hd8U07YfKqFRpT8Y2HPZx4K484U/kHZQQWEgHPnJhVoOpQ3
9ccji2Zk4pkIR9rrvMZW0GRz0OnCPSptL1L+H3LBJD+uB4LZAuToLBhPrsAGQrvA
lC8F/JDEWeXXBkhavk+PacP4p3IpJuptu35i11Ebwa1lZSbZxBcCcwh/52GQGxQn
3Qf/LxTEacs0XB1te/eNWFKc4wbf+yPyoCllPCpnIi8xH240GW5lgtLTnIZr2zbr
TyeGe7aD7V5qX+1nNS3PZzLbIfHoe5No9j9ndmhXxxEwuEyISMbghYzNnAc/zfPS
+LVKpvw3Msld/Vsc3DxHCyOdN/2QfTqdGqtQuQx6Vd4URaZOzPlaYCxSFuVGk9Yy
87rvcHS8ih4THuWnFlLSa9Tc9oR/Xsoh2vDNZfZOJDXvFu/HxwZcRcQgLm24MOgr
2oYR8eD8BYtkX32JSIcth0WzOjVPdpQ+a1vg5Xl2lqjqLugGeDAIV5Iejj+ObLHa
PHtYpw2oFvMZ4eMI7eWA/2ehBR2rSAT+Whk2zN9Qh/wkGbl8Wz3SfhD2Yax6cg/V
AX0iW750eXie7H9ukRt8/f14A5UVJeGqQcV3x3CuFDmUphRU0JDwcv5u8XuLrWwH
iNskYBsWATa/7wmaXTdy5BOcVgjXjPuSMolzvZuQxtpLkUcUoZGbTVrWAxn9nFcS
TRbJaWYVi1hcakW9VYTIPLbRjZtGKGvGDNbpk/pWzX0m8/pnXo3WmCqVFRyDe6go
445Fa1tlpgVBRJi6Nbg48suqI35BDCcl543UEXMg4u9GYsyxH82tkTni69D43I8K
CekHUQIHIjtRvJjRk5kAvhhXJb/Qh/khlOH0QO1tDP1bXTbOlbB55hwWrFL/VwWX
NZ7DUvuZVtyraDMYKgTIc6JHYDDwGeSWIMVmQLmnBI2T4SM0p9uW3IyrSs5RdW+a
JvGUiptiHbCQoIfJ3h72VHvmw61GgUJApDoagJDKeCMS9AlCwLGlFXgmZi43UpHR
bjXIriFBQ1FQNvJa7jAZg4WKDgsr/3PdlqrM4Va1vWYxk1i0Jo166WOJvKyUqfNq
VLqhCxLPzRovCtuBvBPkBJ7XnUSaXOfvMuCpSu+qrPPbilHsS0zFCRTkrRhb+STQ
WfBAQgqhhsl2TW2inG+U1i7EFeEfXHE9isSdYOf3l+TJdMuKXnJA02sSvcHGkiFa
KXqNeFLEyHgcQeJj4EJTbo2ALHaU8wyj/zbXLk/6th/H7+0bIeKZdaJsTw6aoWzy
W6yRlawURizO4bcne8DsKi4d06bI7eT0zZ4834wjsGPgcy3VOKl2gYcIPdooXJm6
lP6zwF1de5NTnMbBb+8X9XYWkNFdYI9L8ZbSTQ+Qmk9XfSyoHwtvrIPPcMS6SHRy
bmHo+5DJBIt4L8WY2WTKaxq4ABa5W/EqfGrg+ITiMW2c3Ru/8m4j4r9VGbqK7lYo
gBfAQTKv3t875496WM/8kUFj+Gr7FGBidU9Xvmi8f81xBaPsEuYkoaU2DHSK0x+9
hOEa8qAhL9M444gsUUCb1pl76TweRSuqhevTf7cwJqvrysHzhioTZ6WOKZbOKEjY
mlPZAuuLRTv1Jd8J9j/XPwKLOb8dHLhwfCwD6KT3qKveGjBU0+LEH7EmJqijaSX9
YgmaiqFe+B9q/BmqOediPeWuKlklrilZiGB25D5KEoBADQD90+Qoz8SKsA+AJdUx
1Pg1QxFr2RglAXzdBhhje+9EwU2JdpzzNuh1pHtDDjrQaOQnIVTBUhniQEte401j
xqpTFqyLCc7iCDMYqlhQPrDMydEOGSiktnhsRy2RJ4VLR+6jUE0RFQfyh/NmRHaP
duJwAbvBTbVJS4XtTlC8weRZWlOpuEXh6gfe1Sim5G2NnQ2EWco/STf3uzzRe4Wy
v28Ji5XYmHqX6c5gm3F6HHpxZHoAygGYfLfvnMNQw2w+zmC+nlqLBcRz/1ft699z
WHzaiHaAx2HKXKvJt6jjvjf5m50azHEbxQnWPlEAcn7oDhdldYdZyHCyzst7mkZI
TLT1uWStJF8iSgjVi+3CjmfiRjZ69sHzAGI4fxok/+AygMth2MOhlYV9QdzXqGf5
fwurjRijDT+rsAPfTOqYztw8w+bj/S8P4iJdnSn6zWDfzMmN7zU0FUJ9oJo+QE+T
2ds021rCvl/zwTiiYjIHfF/eWuG4edLc8CNtXPHf4OtsfrHHMElQeD2/cSAeGqkC
8jqvevhs1A2JxjxwygJ/oJzCPm2tALOyYc6KwS1k4lURuyUVftAbzXWWVlrrNPVQ
bLTO1QSViHlpqIfkK4kT2u2Zp3IKbJyyJvaNV+F5URyPH8+bDTDISRjYqUq/pO5j
dx4PC1CHtusQ8NWs54jJkhePVToXdf7FZFNpch+q2ZNv353wcJW75P4NsfOcjoaq
j2ngNo6jP4q9qXPyfHHIEkdMugbEJoq+uCcVdsam6ZlzQ/tS+e/r0BXfwrrf+DVv
I4IXE1rp/xHxzNXU45alWfwvOc35Ji+P647jRUBBbysuYy5cyzsPnTlgECgUMrDf
zkKVqdy5KLt5Dc9a6VW+ujP1OgFZK2ApYlfBZDy5UDKU3/Tfa5aJrUoSFEhyPRJ/
RmzDGKXpa+OgPsVNMAdTakP5Z9TfFZ+R+5WZ+CyhWpZWboDcCELWYV/L4mE2xjeP
dOoFhXc0ToahwuXDdec2tabsbiXpWt3euKnM7MP4RLeNlxVvr85Y52rRmk0dVNzm
588hAhV9Wf8DioCByCe2RK2DlSc8XAi3lmWVHj5bZ2FOK6bLYo3Zz9shK93M3R87
LfhpKvhIqNLxrLj0TP+wxhQohnlj2kqdGLubcDgWXxM8yx5I3WADjSDlmf7C7vDM
P3P7+8aW3ZnAEq0I3sIuGqKI5kZk2s/MHt0IEBEiFVmOaacnpf2tPA2gNDtIOWdx
qurxiGaC0bJ8xYoImn/d3USQCFZv5+16KQ3OcS51R+2+wZ0aZAzNxKd+4XbvRJCo
HbkEo3Ajv7MpW5F6sDbzes/NoYx8v1xpD37W2OGpA7017K5EMVWR9tHcF/rNwXWJ
5valmbOWSXt3yg6VhNl2tcrPFt9pBDHFoenzFgM3l8rjiQXReEZDDpTHI0EFVk1d
sXi6W2zhanE24bUn6BC+X/l4uK/elqKiUUd8o1WsiASHH+yXCBLc7kdkomTpi2uN
Wv66okJDtgR24XF56LdShRiUfX6ZOjgp5Gui0usLoQrxW8heRLlrKbVM0daCKWuL
TygN5z0syy8mndDKcFX1TeEwgj0ivzytWwuGz6hGrnMxsYUYMLRJ6yGt0TYD6hun
I+f4Z6D9vSKZOdTBbDMPD/DCxBqV4nXKBQYxzjxu81qJFqHDhgm0sgZUqfrbVmLn
iQaOmitngLAlpwSQAL6uBSkWUn6fJ5u1ddy1Z4385ZEQ11g9s/elZenUrrJNN3Kj
xP3TV+yByHKgiZRMlA9RiWfKuyH5lKCuPjMDIXPm3g/pHx2DSyORPirFsMpVI93b
O/CXDoQXD6FQMjBv2pCZiO5n6hinGDT2Gy6sAzEDCJSdvnMVxaqQN/lXc+qjakNY
+cTL49EQ59BSnd6brU9Mi1NgMOEMSEZWxnUhOkqRtwKkVG5Os/uiTjLMI6mcA3a1
cEuUV5h4+wjAfqRj3/yPDhWZ6f9QJYnt0smNvDhWLrxQqVZZH9QeAeFrS0siqWqD
NWAz/OOdd+MrwXo1ZptGso8Xb5zDvhvya+d+08olYZtp2fDcFQD2LgfiDNwrs2lc
oXj4kXjJojZSxFLVMhiFecKcbYFKlBRiLfMbcjnDscJax+ZH0zKNKU9h/TUwM5eU
QljH3SXW+dqHX8HfFt6acuCiH0MQyP5i69ziTJI4uhsqNnxqD9UJtmicXpff7eXC
kJrHTOMMB0yx7kOOMAokEnK2ejUF/iSyqlXBfuNEJMapG4hupKp+ClwntpKKRFsQ
knzwSPjgZLthXjA7ggUmKxUJ4LCFTFSU5nPBNqmG2mqSixEspHq+n/QpKKoRb0Ng
pV2rZWV5RxqBdSx/OvezatnY8hy20lJ//eSjNOUENyQQJHFUN+3bG7TwzpmboGpb
iJaeOew5kVKfs1mYsNgurSXYb6NuQi8FD+uOHbIJAzGDHhNFYHxy6fgBntSV8/+q
HH0h0ybmMuM4vayQTtkWaOt/wt1oHeXLb2n/MwgbolcQ/KLXdVMdblXR3hY3uxmk
iU3+YQbp4vpw4ZIAmu3yxNpdZRBAPRCl2tWe9G4nsL3RKEdk+lMWlta0Sv1QUvGj
MrI3pCnDtpnN4QwUoj2+oQnTt2WRb9RVoE5bHkKtOYB35DK12P8Wb97A0WuG+SP9
JioIEeT6NgBG5MeGp0cgUI0RahfkdcOv66UaSfCVpHoSK4HlTOJyUj8bo2JWRAqe
wPDGt5+GwSgwSnkdZnR+jYBEUoGMC/V7zYtrbD9ipJ7DQ+zQ3t9i1CjQZwOmoCqb
XV24l4yLhkO2nesVnjfP1TMxTrUI45UcG5OhOwrD90vq0kOCT0S8MthpHeHMvLMk
wMGNgbmgh2/DMpSKWhZoQN6B26oy8GC6tnpB2hKRnnSnUcuKUnPUnyg6KPJ3XxFu
9IY4/WXYQxcbp7Hfob6YNtbkRvSzxBQc4TUMU5k8wiNJVYCcxQnaHRNoA/gQLngV
BaV2Notd/DnOVDu2ynrpm1ZXUL/hOdszEQ/D3CmkzbcS/AgDvRJHS1mTl03qCpdN
CnmKWzxtNm5YQsMoFpxaOMPOg2EW4yt1/CsEj6SqtQU69AROuWd6rZjUuQyouoa8
x5mu39QgBBf9CgiRpIqhzo7822rHObZXImrfxAvi0be2i073IK4DGgXusHYiiDMz
hVFRX9i9+SKpiVXxasCrTv6U4jms1gA5jjbmOFI9U+ZEz2ZwJwcpCi5P7dxyPtBq
ZNbpdvyET7PwqCsXNv8rGjn5AyTnR8WLJolSzEOSuE5uj+Spma47OBnVCKFuDezX
FHkV0Mwmpj7hru+APyNRLS9vUDnglHB9uVcG+E1GEJ+Hpmu2nC1D5QB/e7tTe6BP
C3oqPb0R+h49yGUR7R08cDaXzPPfBj0CdJHNPjcYGB8Dnr97tpiACfkynm72rB9x
4fLrsdvD9VBiWOdvFi+PtrNYfG4lEyFN6cK5GZshYoE1xWetJsAYJV5gtBtPehKF
0zWCnZQzkRIIz6phEICGUdgntXYi2RUwAf6Md9b7yR0G/yPPcwn4PPZoZFc+rqlD
ZBwxcI8dry0r1hFKpnUaTzGQbhSijg1LRCzg7Mlru6HO4K8C5zGu3sFkyq1hPoxB
0hGidym+REaupVJzUd8RKLloscoRlZE9bJFXYvz1KrqaCW204x8+OkJvTSeaSr2E
06YYxA9w5U748eNnKhames88c7KoJXdPJoFp3CmN+NyO9akH8nxolsFlgWAUL3Gu
p6TZgQjL6jlQ6Rw77je9B1B/K59VFzCgxQLfY3nJVagacZ2iyDvFbyC92r5IOBJw
Dx0lAFs09Cw/MoN3Cy9662wFNoz1jG3XdqYxOaLO9hXWz301vQt3e1fQedkGGXam
maGCTW8LBaogFWO0VnHQpBOKNQr2P84tFjoxJH5oyDklLEW0OH1QughsUp8REAel
Kzcgh9RsyVrVt3o2Kd8X6l1tKNP4hgCRQw6lD+mPbwOj6F4rIsLJev7LwUfO1lXO
1pZDEP7DeHlwWYaKDTt0Wk55nq64ruuFJ06KF8UyY9z041WKpQADqwCXORnWhZBJ
Ki/V8X8qHig3QZvtRnQhMx4w9L1znDDXV+2Nbfehwti0sQ8DOaLMoFdIpc0fLUiQ
UkcIkMbWFnZKXiq/nYFMUD7Jl3eHywzEZHJNfmrKFHPGcqqGOXolZKYvFXeKZivu
AFqhSzM5+ZxLTm0cVIXeOYzUQ9Jk+lAKfALUFsH39hkZD5CI5XtQaVSc3fbHILeU
3VD9u1m6iTSeT8h2n3TU9YHxGWg/+w+OmgpO7+hXnOYr21svkMq7Pn5kOTp/EPgp
Mc1tVmpsQLLDyfMgTrPLYnAJybbrmxVKH6LV/+JxY6aFUzKvw57JruL6wIVS6saU
6iQrubh/ghhXCd2YhzNhctQURyh/3+8OLKcACfaN/LytMD3qfcdT1EjjOfiVXQO3
nDUwnRJArHCrILj8yp4/cYVSWiQNoSIjzwfe5WD9ciAF65Mkh9sjx+ahf1rQEnKP
s+bOK/f/4T92a6xoTUsc6oFH2Cg3bNdXdZ+jZUvMUvQmu5ULm9gBSw5Xa9MeP6Xx
Eoo8xG6wjuOuLzBcwDl1VLX6ZBDusH+CH9d1SBuJg8Weg87fejTEWlCPzM1J5298
aUr3CmUOcRBqfa80oNyoSW2jVDuTS96hJXZShIZ+iJIDsuwoOjjrzYwheQo2fpyZ
tcLmvUkuY0pIPjp0jZFZ0hBvhN9hoDckAGFjnLI3G6KhUQTHzoeSXRFOSsEvxite
hV9qO7YR06528f6306534oqSi/UZoARKMigR7mF9xf1SuKdUrocQAMfUvdCOHabF
s+jlzYF60SUeY9JVql3JGOmgtpOGFV1tliqpEmWezz2jQPx0gJTFOc4bxyjPm265
kFXfGjvkkYVAYsRN13WyxOrnqMTjbXhwdZSwKKMmyLJyqi/ztT/fsaFjYZmcXBtA
p3x3/BOXjhNjADLvZomNoIArW6XMRzuIEQpdEFAmy3PrspBKtpPYSInqbNZ04lbC
lguASdTt2AdSSFsVT2ucZ5Rkd16OKvXT1d65aj/Bjb+OFkE/tIGyeZgQNwqvwI+f
YUCfKPZ8/fuJePkVTVrfhBwGYJ4rBG95hrpKfJRluHVy+LsqRYKIx1d0mkVZGpLO
iKb3u+u50MbKpspmUj1A9G5nO56Ble8aMV/GCQU0k2fytoK5Oyh3nzfJm/Rh7Nzj
EDJObdyPKfJH6zdPI/njqqFekjv3FBZ0bvhN8iP41drSrOJb1QwWpwHiM/w8GOW8
ovhv8iZWsDRh1yyMcjHo8VvK5zbfRZi+zoN7JxSN1/U3c9llEyiMw0vAQU5g4xoD
kbDlw9fC5R/k2u8od8gM+7/5fBbuNKxHgv7k/iu9vttfdnyl0NTGbP8Nw/eQxVF3
CNrG1G8d3dQbCUhpJJ3ZCARWzu5p9YWgrirkuerpRy+9s2yqIJLGzUE0ApdH1j2V
KlyPVD+WWh7w+HyQJW7KS0Rol6BG+0ceU5raSKgPPvRgx6ASNo+stfsnjA55W+aV
hl5YD3yhda9lOFXkIzMdrm9Qj616XISqiZ2T6DcbrQzVvsr4Xq06pG2Xa6AB5+PC
D+qyUMUKHxY/arF3ETqwRnFZ4bvCXux+ll27EeiLfpVb0XRnAXtHl4pEoAMdDiee
IwRxtJ/9MrCwhNbgW8RslaqaDQkCWzdHyHwtJTCuACXC9BCN2kkosCY0dXbEJc8u
venGa5fjavAiCUIcOj82GPYTb5vnsVEmSn2USwIsr5LjCCm6XoRkwLRM5a39vRT3
ILa1ixJuygYOUkgN9t5uH4I4NQl4p2O/4i5ch+b0W6tDNeBjbjXeulFk0Ym3iwUC
ZhFqHI5ytgcJLPuzrw9BdwkTBliQYtaR5KDNpOUHwOTfzsX9QUVPGGp7i9nFR+X5
Hn01g0qbzIvqXmYNfIno+JqYraZgWtXn0NLB3BeIKA6MINr8tEwXBNKw978SlPdE
GaqQzdjCc4AmEi8b8X9LCbsEE8isgtTktgXOtMFoaecEb88preEUXmGFQzid5FhB
5nYmho3rhUaaBc7cI6WyAA2IH9vsy5O9U+YvM4/S00UjXiOmYV3eLn8BQNjgsn78
3fJPOkqwV++cLOXiSm0sD3mlXM9QGjAtnTCZafoBCOb0mtl6dnbkWPty22ZOoURe
PwINUSqcgp6S1Q/VQYN05afCn+GYPyhN5nRzTe8MNUPQ5AkxiDwteowvDjOXtYBv
pTVmSvSmUgXHLddsgql6Z6n5DpZLnjU7CG419S+jnH80ucMUXwiEl2cY2VlQXbCC
wids1VazpuiTuumTva5O2i1+xFYrFoS2NOkK5MBiobEwBjdNlDMoLkHRDY+8iHhU
4yNrie1sUYkshaMc4muBbob7iItPZWhj1BM0kC7r4NtL5B09RVKxtQs+Rx+A3U8d
ZwNgvyqctL1iZVg407o5HeaFsMKaAyq5TszRH7lMQnkVH4HgqWaqVoZNXrWHUuXf
scfjq2m1U3Gb+fJux0e5Lsd867IKaskqrxgB91PmfaOM/CZcireIk6u7qgb+K9bi
Y1cId9CUB7PqsgaHDdDnC2jJJQ/yk+1ZiWAA9oiSHIG3fbwJ736S/7d19MT1TGnC
FdgOHGYtirHpYm4PkgdqlYme/jU9PHl3q2fOXooalPbRh6bDpVT0USK/2F33HVGd
kLlXBloawF0YsLUvIlQ/eCtxs7keGhoDc2DE0A8fNknFNFXyNSA4q/Pkx5W+nvfF
xBFFa7vW5P/kNqg3zIocY2OjRhzYZ9+ZmreT5+7siWeSxwfw28S7UjKIahch0I+p
e0tA+237H1Ny2u5uaeBe0TUQWADcRe/BV1aG/33bhB2iQJhwvq2SFaoNZcLf9LC6
7e4xlLWBiecMyKIgWx3FYQlr3mvHwdHVjRCuabBsfyfG8uzrm8GY9gObz7EmUjzg
IA1TOsFo2FMLPEd9T7KO2NqfqqF0s23SxnWemUzDILg5Aioj9vxYhIiEyoSMFzBg
X1nArgvQug6bR9/KxKgXaZHg/8m8ZqFdsbRSyKyhtnutUhUCSCKoxBAuqYxewQXb
MggGNIP+hH/A4WYc4YX9uk18CTRimmBpOy/2ObEdqoK4uT2xez//FPzqsSqo1OQ/
jBhKPN1bBr483qqVlJmxK9ChPwAMjIenxvtBKA7lTiknrLsvghaDfK0g0jKcPiLO
RPkR9YW8hxaiEhGwRCHsxxiNe75i9DjQx3j24RfnEGX74FePuL8crVFPmO4L6XlH
3HHHzY6/9ow8CMnI5t26ByX0sY+h4L853XzHiNIs5VRz6bxtWFwUYweRoJD3faAX
aMXDp0+YDAsC83MMowo1PTLEiCVvYv2APaOrmlcP1aC0Ho7bhOv+GON/kFz+CjOx
MgJd4dYjNfRGqPLNrUQZffJzcX1UpqyvXInUfaushHSliyKe516du6n//kONqHYt
2tmSq4SbdDoajBj4fIk1KroGZJ/YeEoKFjfheR/QMbc286aqhUvwkGRcmrjiw2zG
EwDkgE7UB444bsrJOARP8x2nxu28oAk7tW/h5AR5V//xvBGZx2FcPSTs3GWAoASK
baWMsm4iOeU4Zc92NEJ0/Me9jLqJRujlyca+CGDAP9lmKXPsAA6apV56Gs7/bO/P
33y2jB3Kfye6s9MMFc1S/PH8nbTlOoLCb0dPOtx8nh+9qpoyVt60ZYYPGikSDBLd
pvO1FRQ+rWACyKSeKA1lFz8YC16yuqgbzP7FmpVjfyeoBXvaSlfAxrFnE9mkm9ZR
RkFS63ELFJAYoW6wSuWZcznspZCyFbEy8y1EfpwJkIHN++okwY1OLlXYFzbHzENn
FWV7uEkFzCvX040jFWJYvF7GPm9EzGOpS8yucNXty1VWnu8hV1hiA8AhJmlxVSoY
8LKsweGvHUONDo6XZsen1oEjlaYiqOSdbBGJyGu1c8GacyP24vhjG9lOQ/mAq+81
go8+mdWMnkEalL+mwjuY8I5jO+zhNbjfRJCuD63gjZHymYETV5dwHX3ZVi9qih2n
jYHSzVaOO4FCo2wKMijT7IGOzHm20r+rWT5niVEYVriG1kiaYQS8nxk3X/1rW1t8
MevcpjKZWYIPpPH7ASZPNdkfwMUSXLhakDRKce/30dSouxSApOwTRkKTqM564vae
tTr7VkcaQ/F0bh1LgQ0UbfWfukzcXHPXAEGc2gVFzoeNunOUMnPDfx00lKyNJ3zH
wab6iiRQuqMumZy33AJI5dzSzeQoNbCrc2liKCOAP4rvkYEsR14mFPdYPgX3GGnN
QzHuTBEX4in1pnJQLQcdB7nm7+euWFk2fyZDoXHFbQcckE6umhUW4n626bu21hEh
/1HpQ59nMrP1aqBmF3p5npt+EJHXIjG8XkpldH/VVGikLB66+s5NhuLl03KbHuaX
JyjsL+Z+YPeDW61I9lidzpc4siXz50glLtWzF3I+Lqj9TXB/PPEzw2R44Cg8+aBU
T/T1ZvoWWULF/AwyKD/NXYvcjtcCjnX5Bl2a4nuv9jivH3deQiO6RcIi4Y3RYzYG
XosufV+t9nf2ngBWTyGQwjwAif/AXlVaG/qiuoIGQcnht6c4gVQ/lnJ07/BXc9sN
MOyooZHIgRjXkpI4+vYVLGqvGSjAFLe9r4zYXP32IqH1m2MP/HixH2/k47q54B8f
AhfL/6X/mc37z2drtZBjSlhdCCu/z6doijcmcYmjEe2RNHag8rWDXqi26K0xWFMj
6MfMnieXZD5+PdfiDthtyr4PtD9nzsxwBk00eliRaf8lJdXOKabpno/hn7vUXgX3
M6HlTx29LFqxotrv6oUxnMKi31DmC6YVOeFGycxXQGmVVw9ULGsP7GpV2tdcK4Px
HbH/EMYw4mlfiMyzBhy/8oS4PtrcxA6hAT0IkNTWKQJvb28106Ci+aKyvZkiocY/
fVmW5C6mjVX4F1pNOxzQFay/V1W6I30Y6MetFzn4qsHZR1HQdiIl5nnBNXy0A3g7
c8Qp0IEee/3rJply8LgJ3Ie/h2UFgI5IxQ36obA11+KJb4FqdWA6yZj46uIC2AFx
HJzczb4P2dh72xmch4aE+vtriymULKZ1yrXAKuhoAJSHK9fvmAz4F1OfsBk0o6GM
KUnQ+eyyWTKzRQqCT/jDzrQWgDy7x2/emP6IYY+hjUXS6LHj4zWSLEQP25o0L8NG
pWTK3/5pdYrcFAJGKFqFI20OMAnXYXhgmVo6PCNM9rykNp036aYgo54p4heHF20l
NcVEiSYrsZgR/k/8YrDuLjn2ytCQJR4baU2Obmvt7dNLEqTImWmP/8mtvIjRgGqD
+F/I0T9CD9PHeLSAFpBuxMd5No9+2baYgXCuyLDxAXrewhB/ZO7v+wwOZ0RXnzn8
mzlbMLirnrKp4HhmClkAoHL6LPKcsziH0Qjgog7ZCJ5ivBwuuuqmo/b+DevP6bdZ
41B9T+nJpEZWmk83HTzSghGukCTjYSTTQDvY7vD7fT6J3BJI922jiqfCT+NZXbKb
v3fdfUerLVLD1vJgog8c6mOI0i0e2ee8etqesuOj0ojslHR3ys20wG53Jcten+1w
chZWorPvp7Ou5Gn4oq+7p59k3kBdl+ZsXMXWA0TPo5G2Xx9a3Odj98Ryo7tDHvW/
el6dANWFd6E3VWFG+VqJCuVVElP20dlmlJmj3+kfqGX9FaY1+phqpKe26tOz8iOH
b+APy9wUbLryMVVJ55K6vGcevkTutp66hnNwNI/avpCzlEaB3rJlH6wU8iNKLrWF
HaRj8hJJvVuLMvze3hH+4lx1xe6BI1AColCPsZT+c4vmZzGwnXHID8zjxnUzoMQm
AahyPdzn+jqIyFjHbpKxaphI+lkOdfkw1RBPPjzSRUjo4TpN8rf3eRffXDdzOjrf
INT3DeqNe8NmUTo4f/5vjzR8wlyPVztLiryWSufkJLQh2Z0RZduwr+YSZDkJlpeq
an7+NeUbik0Iv8bgtijIOEXpPy3jV+B3oTP7YNoBQhhysgqe0o0Sy5CRzKRYB76i
NVD4pnANYRohNgjoCSjxtydStOPIXwiM09xinXwEGoAh6V/QWv0Ju6XyMavgRZsn
/CbEe+QjCjhMSWlDLnnA+1OhIwaHhbFPgaWxL8PQ8O1qLFPCzhe+6+Ndatp+UVII
YDj5pDs1SWnKKULcRGNiYDDcA8TFepbOQdeBIG4ffvrvFBKiJ9of6lAB0DXGoua2
a4A/I/u6ORHoTrgB5hQisOuC4r+SI9/Hq5mFV2q7wL0//uYBxplnC7fuyKns5+Mx
P1rIs81Cg9uxL9ev3xpxt2fkY8/9yg1IPKR1A80NWUpCQwRMOhjJFUbdWig29F4Z
RV0s0JIxyZGOgKwTgf5KpSvXrFmOJrk0GB83MpxXkKfguSNZr+PH9mAlfpVOj5pH
jtElpsDIrqZYPsBfgnEUj0QSVFXZnpM+7Y6NU4PBq0FfwcJ2qxuGQis9CDWkxY5v
YcoUtWebEWQ2vWPuhrBeXL3cv9sDWNlnF1z9TdvzfHjKTixtyLWpDeqFuWAe0SGA
sSENTm0FmY5RZ6brYJV9katihpp3iiukJal6abpbyE2OwlG9xskl0oNH3kKbj7zx
eurlVPsgtfCR8apOlJUvUqoj9/sKogsIdK1xCoh6MY83JDy84WMM0b7qtQexVD/F
Wfn1fO1G4r3lF+aoSsaHXFPhFJ9bqclbwGqqvEqWtspO3mudAzFyIfSigmwyMBKu
DdJIqPaeoaI/WkaKBJYHSecnpYkHdieh+2j1ItDINZAjVL4OnCg5PCuhseO3XpIu
o+po2I4AFevAAxHW7aiC39IgHG71vEofcOBL7I9jNU0VGK4KKHC5Wm92zxvtMX77
65b2gI9WDQ8U6P7n/yBl34kOdxwg7GrFNFQwC+tFgPOOev2hrH49v0sr/WyKM3Hb
Ur3UOegIKprQQyKXz9cvErLfJNZUil2pWTET7ElcACo9K09Di2rzF3yfBCzmu7RW
JD+Td465fsCtG4U4FNFdonJ7OvYHpWobqleBQJSJkhJAVFFaa8trqJQWOTn+VrWn
RmgHQhwpW49h7UJdjHEwIu8mooeZX/dLEoRY02K93ulW3azwS10exAF2UAB3ZkDz
8qwHNtnjwKCB5riRcmPbS7xd4H1N82js0moCoKedZsMoSUsbaf3jhB3cKYfYKeR5
qhExTFAzdpgDHCgv0BKjjyTnbTdTCZANTAhYQHC7eWsNwXNs6HHqpehpVTzPPbiM
RHMiZU1oDW9ZQG/n2NI+gRsyrOq7TP/oq4Yt1b+RmXfFd4cRj/1wc9VWhwGGbkFD
W1IIL/6rbgTsqt//O/u7Gk8cpYvlGOTIz1OuyWm8f4ebp2rcR4K4rgxl4wTb1DQK
RCCfNqvrm9CY29aH2UimzT6GH75MN/qej3CqI3j8NDUfSZ5hhqH11A7uO7VdiIxp
rBEuwho4DCX1+d81KLglWTHXV2V9wL7i2DPf9bCZWjzOhb4lgNU4go5xZK8QAYzm
uWczbou3pXyTloi4/oPwtN+G9WMSA4T43xBQVl+1Xqtna1bPC+dK31Ml48EDx38y
paVC1uzjKw0z/8G64TQXu+2cyaeNxkffGMfG0dP/XInWNxW4HD5bJ7jdxyGOKW1i
8QR/B78FsKmrlKG7x6nAMrq1b+skwqGzS2XS1NyUC4mrhNqoUGLUNQY4ShhV8M11
r7CNFDb4Zjon+hf8Z4Jxo+wZLBk07Xg04/S7F4cLxlNKHkGG6+WAasF9Y03CYjcL
0PUyAZk7U3XC3zNjGcT+nZ7npf3T+idJ7DaYXwUPs57Thz8uoe6hLSa7ILliYEM6
8+udbImeaGSVEm1kZEg9qsQlGX4LgSdtJ13eG+bOFLdK9aqzqCA0Es6tgYcH7Czf
Khiswfdbh3gOVNoYV1u3vkUHqhyZOhCfG9BNeeeYRZbCNjOJewaS0qFRqvXLGpHI
VUiip3JQVLQJ5FuRVq+2aAZ9x7HX4/l4iI4zDdpfATVjPnH6rDMOew6xRrwYZbv3
pZLDgHslQM93Au0bo9icKb1NmUAb0ISTna0HyU7NsM10WWNBORzfr4BoZ53k6LI+
SoPgSpMXft3RoJNhRzktyWMzEtifVMAuIe1FEyT0CdrGtX1lgFu5A2KVGA8KSjWf
LPfLhHx6GO4+94OCi93b/HVOrHuP3GpY4CpGKYpR0ibkJgSiYxWvUvVCB/aWVFhA
BV5xSLhhyTm2/bCtkFfRHkiLD3MuTJBTx8PUdwU9bR4AjvPJ7AQvZ5epLV9jD9jq
wIVFmlMBk/sUi6z6p6kqPjf/eOWxvDS+QRwsJJoZRz1cikQALxQ7bVVK4wPPHUrP
GO0tyLBf+GU1qtP05WVJu3fHC1Gr9u85P9mZmQvBV+iof8jX976MjDVxiiGZJKps
hXYy/ZyC64dqyLkbRz/IzglffWjTPHHRkn2DW34XjJ1rnIMiZYjKS9LSlHAmP0ZC
GzdD4CJmYUKrIj3IddEyyr5UO/GINqgG124zrwDZ4zNfoJ9mRHH6zrDVtqZXLhIF
mY/FQGPZXExSH2GnGOTXRlFgh6pxQmFLFWGLwOPe+01RVxFz9DETP98QyME0iLEF
5+SXq1rOu2OVPj1z1+gnP1V37dlfuqnMGPabpu8DrH/jji0hoW7UfcI23JM0Bfxa
9eT16bJAnWZwUZQsP+N+hfwQcyQtD3mvtFdbjOOaFWRmayUgBgdUpsPYZE6LCQYs
fSTQ0qmcYd/b/J/yiwo5BqdUVoPzj3jNJlC44JeSzDbd/YPK7e2CSzjZvYicVG4K
CaV/TZLHf/x+4VoqUv+1xV6atXUgCiYHcxFmC0o9tr7dRXfN+8BLsrAAfJhxBq4d
SUfV2hkpB+WVzbTw51qwXMK6SVPkwbQO7U1y5FEydV3yn0w16WYoAK25K4DK5rxs
sAgVEwa0ZiRGEK1/EyBcrgxonZpdQmkov6PDxnqUk/mB9lkqUVoChZBnEzWJBCoL
xhh2888d0xTYvfMOQktoWvUNJnJ/RsCR+Ekjv4ZZ2i24SHK4nQ4qqm6l/MIX9Z46
LNIftKGm1xyAzY5pcSFvePZGlVIeTH7beD9+3FoWICEIhF/SkCNpqTAbrTPZgGaH
C8Qd8gYWvAlQ51CIPgR/lm5jUUTFmAqBE+WJXw/P1lWFJ76nsz2yeo/NirbXK2EU
LKd6oYW4LS/bS9IoYwAlml9Vc0q72mOb69MrnC0OTy6RIBoki+jiCy10WSp5h0s5
L5a7ovtz1Yy6sSZ4TzPcegjCYXXKwNoTYumFU8Ps/7vtSoIs2i0lTTTyyScFQJno
OmZA0pGdmgOG2OVJxuyePx2SYDJGPDD/YpGEfK2rQjWtlQ6U1jPEaK5c0hXpDzHD
lVab/2L+6PqAYP7ecS6F+gYln9v1XvIiWJWJakT4jboW5LQziMwVy1W+m1ExQiwR
YftfeMtuxr0SdeeRex0Epl6DdSWYekd590eM0jm+wr2uyLiVPnSC3af1H8ZjKCvu
f81MXxtZK9/bi9vfmIB8YevMYrZkGdn0cMnheVK36EHJ1EGzkdZah1XKICqmxFLr
5Z2Z933p8/iFSUPbEBLdQPuAIxQeAMCJBurrb2nESrYcsEvBUuCT5CbIzmpV16qu
JyHcWUZSzkajFodbd2nBFykGSps19KgLbS+cVFy9+5oOWhy25yrFsb4R0u3ipLF9
NZb82dmCcjMDpfEUul28AJ9Cx7udIYOZ8akgpLEC9ZZApYcBWUF/C4GDvSTbKxKk
ByphTKnjmkh0Xven++EK8qaiBVlq5XT5W1Hwz2jm/X6tk9JwTEyMTOoCiUvDi32S
UDwwDppHeg+ZjwWBDg5gfsjPlUu6eteF5iborHrCbU5pfPCPdAbu+G+Yu4bWvJpT
zwYK3gHO8iAogF9+etQRIzBxlVL54c5odkKXnZRMVyfujfj/aSlVsj6Fhs2ptfgK
N/MWkJ1dFQRpxx1QgAk2mhupS3wOwyNpVp7CDcsdb1enD57Kxo1BsNL5bUYGij6i
1C8SxIImmPDUcO8st9RRTKwYCMYkN1SSpiTajXgod6VYBdtrJ3i4qWfvtfPSRMqA
frWF0ywAC1rrwK6wBivoH7RCwjq54hxY2SBPpklki8mv+vd1T4uUOzgG06TWlu5c
9twpI9voXu+TTCUcNjBAOxhHaQybNCfHAaQiQVmBKFO4/DE4HKkEcykx1Ny/sc1N
vAFc43UaX1BPTYLzPoa8Vd5pBgtCnKSXUwfTD8l81qdRT5TiO1B0ROoRKVvuWnLU
j2yKJPzaTyO33x8A4uCSiSYtUTaTJGqigbAYe2lj/djj7kRKIAB2z4GOSwZvW6rW
XVsRFDHTi+4Vvv77lmzHs0BQAbWjrmN7LHH3dYRZIhd9ach1YI4CEWKyv+ocH4iJ
dc6Eu3muYsC/sYIwQdbiCYJLMNfnN0PhoW2il3tjoNsKqv4jDdq1sbUHh2sXG6HQ
QjQHE27tlNMUJGnboXwXAuGUfCxQ4WMP4H+pOHpsNkn+sh0lZgcs++D6RkELwKat
kvJ09IkGoQJtUIHmWhAHY8jQqgVaFLyszMP/n2M7nglie4r9QWecoXnUMziC6FEN
EkU+H7S5c2D+unkPovt+c5hHxW5dsBJgsOpXJyZf7SY4Cbo4HM9MTPglCsY0JkmQ
Vcx0Tt1298eN1RCqtXmyEGHvra8E1yzkEUazioASrjOt/aG/EqgwPtiCphlDk8xh
eZN59XkncXRENjFzUGf5zBI+Q5+c22ARyYzUwe3f+AiG8MzKhgsk+Y8k8YsrKaPs
taWqDf8eLYaPxGIRg0eaxi6T9sIyts3se7FPY8qVilh/8cieTftbFegnux65EgwF
2mdSlyKLnJcu1eFU/iK1706J+ka2cHnIk/mfNdDVcshOtqF9oDGyezkEYnQ3Lrwo
jKAc36Yjl15b6V8EtaFGD1Bx9bH8oHuzgJVthDFqeqSyLYezy+RWhwPfAXMUZ0PJ
OvrTzHNBYftyw2hhwl7R+3XaB+3mwy5djpvJAulG9Sb6opa4+7rd82ocja9yG0mA
mnjbuqjLaKSoD0H3PKH+n3Z0zSlDGe9AciW+09ESZgLOIApRmkDhTs02huWwennq
T6FDGLugCnrV5KRcSP1b1wx2U/Nrp9JtnWNvMSbxAr5CrFSLbnfmf1lvWXaU9WB9
Oz8CxtPA66uxO9au+qtcGaNfnJNkY+fDgVXXdcbVkz07KQ2n79odM3M+zRdVi8rT
k7mptD7qjD1QZeUdBEYwN7+G3hOv4pvQQenszAAAgt2UEwJPrJPvk5ft0w3ToChD
UQfjwAqZIFakFoxrDcwPMgAT9Z7FyKxd0wTC+p2Wok39L5ttNmfYWEVlA6luAHEG
+pfiCq/4C85KAqUwYEVG9ryVv8KHG2hn8UgJYr0+b3R9Q3v0yc+Atw2+TLhxi4eO
KIoZWg/XC4alMfZr1MBLGCoBsVtZWFpxUGSD4jdGc8UypP3vQCzdPyE0xVC4+oAu
RNKwGz2xguj0OltozsIwqvy91kMweVYyUfXBTa8hwhzJTxXDcYJD6LhG/qJiyYqi
3s7KAHORoikbv1Y9LuAjDhAGSO18ZBWHxk4MLEbDxjAizs++qeckiLKnHvHyBCiV
Hph1OH8XIAfmvs0p4VO8aQEFyUR1LW/vIJFr6ixjhvTTke3DkiEXw9W8oS/Qi6gP
xeCrRe1e9Dopqs4fF2eC0H0Vs2rKXJ29EjgicsWImMMPzDTP0jeZZn7VpdCfcKeg
J8Dd/etGqkgtzLooUCInbv9vNusgE8BwLQOzG2dquQfFiIGLfqZADtcHRGsXAF7p
XFCDAjBPvVcP1x/oSF1lBHwjeJRZaEE1FVj6SRWu02NJpOqFErnfAmRjnYKQKqFz
IZwfgbqajb4f279Crm/iI8bHZ/luJB7STuMapq6H1peFIyP/gP6h0VGlZTMoucaw
E2nZljbK1X+2zT+LP65rt2SXZzigXY0bnoUiwV9UrDnWDIm22hmjFszg1hmwYjbF
OpTlQcdGWx0mhY2KZKaJSlndP89mpW2FDkQKSbBjcIoW9Zrv3M0Ynn7nXsQlx/3o
W3M3JhU6arEuUg7KO0POMuexmr/MOTNr1RfQ9F1//OyI4IadhKq3Pok5zajm+H8a
EaKXxYGyRx48YC6Va6T37vVhYIyICqKjXJ8AYAfk1wypOGjDmksxLU2hSbE3VP2V
ats++F0A2wPRRw/+CrUYVqMNvDXVTRr568kfxaQmulTGh3eE9JJdLmo2wzsaVIgS
VL5S3m7zCnxKlO5+7IZ4rVekUHOKhxQ0bkD2owh/2x+8PhPlD8eU9BisBaf1LGyX
c9bNhcLXJgTX3efoXj8aUuVR5cbUrlu1zurru/Zi/MmKurR+oARAxQ7G5zehLq6Q
eem7kYb197S/4Z/gnEI9++StFW8y51fNSKR4st1hLfStTTTaVhhTHCjsL5SdWL+7
BeH4qXntr+Q6pv5sd4DCVI3zrTtHDmgscVqFapP5k2KPGvFpBFe0PYsghBIM2b82
rTMag+GCeoMT8qyyOAe2qSQ+95uMNREQe4PWs3cruktzN8C2cr2CeKU1UAIOETYa
qQj3YC+Wmd46klbkOHDHsngGsqbu0n2YOKHF7sHnG4CPo7433plmxNkRPRSRA+AU
JtC7CZYp36XmTivPXSyB90hfs2P4m4O2hVCK7YjeaGeJZa+y2MgbOPerZNjMC+zw
n3KeXKaVPVgwzPIlcLeIYrHGUc7iBcwGmXEmKwdO6s3nzH4TGRJbdnZo1sdRD08H
pjcxqOdJYEzYrNN1mOR0mrcTpvD02q4+px0yDWhO6PH5t+kI/pghNL5kbQCC9yrK
m1UdZzk5HX5V0o7dpbJYwjHGF2kghd9PRN50Zwv5WDpPWVLOntYO/HVUZ850r6eO
jbdQAkXq6Kbp7V5zyp6kNOtV7g32y2jTOrFSg26jc29pmUzW3KvpBJ6BL0/8eTE4
8sr4ddFmHOTa4wWwIh9YRMfO5FkI4CTcAiAMJyiqsNPd+6v1sS1Vj9okl4/Q806a
CzcP7kbaf5EQwtsnhLmygHf97XVUUoQ8Hl7LOoE9dqEtah4TFRO8EdK+dWCNyCm2
icgzUxzQsteHmEq/xDk77P+j9y23o32SX7iW5pOCtF4/ueVmDPc5z3/ZPWCqhkSQ
ZbmV0UjPqhCLzDzrqu39WKMiXm4JHiDoV8QWA16hTz1gY83TiF3e1qDMUIjhNVcx
sVp5/8MBfmIzD+errYXy6j44pN5PHOAkw7Wal56w7MDvdT2A9kPy5qY4QfM+QLJx
iOCyEKJpXMOyG9vOPtBC0i67mPWxjyoAe0plja7C5MinYvT+IeOf3x9tIaFAu5uM
ZhhgJwCqFoV1QRcw7uQwEGF/ACM7AtjWyoWH/XmbnmXzNR7+BKtUYe3Z6z7nmmMR
pDT1Rn+SHopoSjKAFRiYukOKGh6AawlFm7AM+x3jgzvnJI8NxIJIm61xX++i1DDf
Qu23vTHHNRF8xKsdYsKKepSQL7OuEqSyzHnvprzW+3Qq/GJ+IFxwc1ExsJEdiexq
UWIc11u9zkWWRkPmuZF3pE6pJU1AS4bgDYL5JXDSnILZkYL9pknNcCUzUhTMywMr
IH5YCJBrcp0mWrtn1lr4/QNBMhq5n4t/TV2YtUp7q8iqIjqDBuXY7FpMzF4kaXY5
jzJPi4/pbySMMKvl+cKUZhB1JtngHqRvd/fGFv7MHQl7W+SSDwXy6Nk4fYD+5yMt
QI55nuIrVlESGJQes9iyPyCX4tvnfpSzkFxzgK8VWrT7mwY0MD2L/nop3vyhjaLu
O6F0P9iD/3K1JFyjd51iJybZquF9UcyFmmCtVuM+7c9WpWesorSQY8mi3Fc3kVkg
KU5Ya9CbeiSqZaNVsgmMLulIDk+jSDPeZoYOIJq5nGdzQ3ghfG04ldYiAD99uizr
499/n2oc6NDxXk9LlmPG0v42juOGs9PyjA265AVLBYOfvxtXjevVVGggiUzjSKwX
b7aSwkP8G1shhy68b2RAwBcDZI47s0V32Pnw/jYKp0z/Dtu3Z70Gxv6fsCxEivZz
g8WPyAFEBK+ipw1NvySOLj79zKKxOSwpzfwplWgyk4hrHxYwlfPi/6uwZ1Q9EdNP
LJ5VseDEVLoMaZxBSDVEigXn1Q/gmR7so7JsoNwbjEo3vxfr+KZQBa/zo2bQ1SHC
/YWgxZNU3VXsU1A2TsSz9x0V9GB3o2bdPrUNb6UwHGjYpFm6iy/743PFdPIDGKLD
pKChvrdIe8kdkaougjpKRB1/xqCe8zq0zPq5cQ57M/qgLzhDA+pjMapdzwSLntCk
BmM8tViplFnD+HNrDBcFvkD6t3efarAa5MkV06FmbINgaIlT09hDSM6QXJhN8nur
KdKgxqSZk/Acr/0AnPlpGp6PlYL6YQWSSppXcBR3C2TPOnEOiS7i7V8mJmb81RtG
lftaK2kKSCgCd/AvF0b1+UWxykyOatAM3nRlS9mem5izNg1WMMFD3CAI9x7DBfoZ
TV9FyW3pP8HEjl6IHhsXmjuj6SJ6u28KSiHlRFuZo7xWc2KAnFiWeq8CECgP/uOW
Zn/JyLk6v+uMV2K1JI98iV28RfakxJ7zrYr+mHIbhMtPH9GguML0o7lFjXqzq4CX
WfX586TzDQmbJHeSL9iOx3NhPCHbSD0ByGNO1cusMFXMWnydAS6Un/U7+qcmOe00
4x7cJ7XOptu/Ca0RIQ9knRc88/O3ywXbigu8+o/QqHtriSJCpZZlswBYEjS3uOMn
2biz+8mlU6BcM0vrlz7uM1kZ3yE2/wLOivxL6kJ2Wawb2GjZ0xLXmamtwJJBNAV1
PZ0c0adkSzqwXs1TxRcqaMWocBZGlHyzzjvFFXhBNmp5WPO09zSJMf0gi555ZRWJ
Msy83Lo1fr1rvgUwb1GZAOMaHrybpXTDql4XQWlaEO/shc17+WwyDqm2/tntkS8x
OkJANkmJVigkIG5u/PXvSs8uZOiq90aM2GHG4Ja+6/iHvXnxN/DmbGe8gxmtVWGK
bDoytkEc0LQgOpSvQQns6Xr+Mlq5QfYVCZakV85tQu3UeK79i+geu6w1QgYPWfCz
9zHk6xlqFSO8vwRzstVwF5az19T+H6cIjHEP7a6hPx9e6YMT31qW56bnEZN4V/f0
0Qx4bUmbjTwEFqAFCpkBIFpi/0+mbyFPn4MxREolofmJ+WHsg6RFDaZk9XKEdTb3
n9nCiBfeTaEF9rL2zxJtMmD1hYmh578iRqpPqlzaOxrnkmhQn/I5g71b8acKRXOH
GEx+gETOjTM0WKzVSbd4/2WnKKW2a0faPcOITQiatDbG+ng5ImfoCoBYXvJkvHlE
kXnmFFP8BaCbKQpJvuGXtw606BF9+40GTLZSLiBH7pK08MVwxYxc+2ekugNnkxZI
Bt/IRBgQlU2CTaS4c86+tWgJ7EPcXoAIaM0kWRA1/6t9PsUcDthnmUtqeOoqSvbF
jTyFem3VPla+486FDXqJqSCFY9NZ2HU9nXGl0xDbZchrhgKZulD0Kufmrs4iuHC0
J16H1ey7ne2BvDdcRHRLKnT33uEfUjFGCMC6WnEBc/jGaisSivty9BvKqezfxWYe
ceMExDyGrW64asTwVREqs49mMWrN79oZI+SGFA0TDFHg0uXwV+/sKOmNIHUwiA03
sYSeShZwkGNwHDIcx7HrTtQVooxv8BjJq/3wbHupSqlAYhv8z0TPBIeG/AS8FINR
4ORKVK3YjVdEnlCn8tNi6XxAg9p4EafyhAlNNQD426BLtsYjsenPoc+9Mou9KsAe
5U+dQ1MBW1wX2gZwzaViVvrKYiAFxtfJiDqlk6xPTwJS3KmnMV1U/A3BObaF/Q1Y
K8t1I3NUnO9Akq2/H//7LmCLLtB9QJQRTpza+dFiI9WoWmon9uTK3FawAnXcM8R5
y36y/fhNidna5RNQL6MNB7wmxJZIWByukTaPiOVoVYy9j7eRo6/YhN1Z5JCm7lxm
OYlsrOc22RaDW5chVh121rhfF59Q4XoXh64L2p4bRT15uEJv/Orx/CnV4ChOaU+r
diEXvLXvEMVbV4DZRJY1uX2FNQs22yW1uOWquy6N7ztzDBPVIaDqOFtHWbySj+E3
wutsbxK2OgVLCzQ5mydUvlK1FujdCJjrDaAiLRFeuYdUUYZ0KDaDYGwY0U08uFgC
Vxr8OkAWD8ZEPnJ+U/RCYeJ8H2o66KyyCq1BuYlqRQHqAQqoQxU3Aemz0nVORlNz
yIQ10HJJQUbi2kXMt21AnCbSuIhvu9Ks4Ljt87b1CT31KU0FcUfiALboHmPyc/UV
g6c4qWv8lyCQ0ZnMXQlbxSyf/xk/58mUlLxMhPyPhsjw49767Ls0Bta9Dj6dnOaE
g8/hfktBAdsP5E96tJAnMrCDH9P5NvK7wxfUlag9inqvf2bUnwx6D/EEKJIuZBoo
DXE9vlpTQH3gBVU+uDFPE04Q3ak/QNHPNnk9CnEHB6Bad12w3B9UcGW+ivLrGNVx
Kdf5clKv9KtViENxzi14rZXhZl3Lacjbv9DKYcRg9VPh+96cfvULIA+eNea3PMda
Bn7HSRtPgXz4IV6tPxB8h0AymtL9SRQHxRXhzdRML6H81XHML6JPrm9Pd6Zict2f
oQRovjzz1K8e4pp96cepxWaa5w0UJtSN73332xG4uwrT59UKSh3LzpwdwRvRLS2c
DS7SO9JTjYkjM0jn3lSN7DiwUdqNvnx+VwV5QjuN+pRsINsd8Q2efElCw6C29qU8
smiAYWRDDkeIIvWP5d2gDdcsir9+f4L12dd3FB6uk3knYYObwU24cYIXadcdHisF
m1x6e4kZ6Y6JvrcawF51CnSzPPBHgEoIYEZ3Cr3wPI4m01vg4OXt8uJn1q7Fnj8V
Jhg5PcB5K/s+Ra1fvI95oe+gk3esfWEAHJ3MGwKg2polzgnpR50L2PNQzMfHYlz7
1QJhmS1vCL+v6tYE8mlmSBH9jZmJzBVyHki7MIgJl9fXVsAoTwzbi1F+q2yeEYZG
jCmuttFJzUqAa6cjAh4nr0wM8i9G4iA1k/EOYKl6UROgxBH7Sq7j7c/rOtxLyn6J
RRdIuRxmVaSMM+aea648nX0jZTFRLqRgUqwF6+Fw4vWN0hpNK4jiH0rmwoAu7hov
p4tn81EW4ykoeBnLG6E5YNCxIKdv9AHuWltXaut+5o7zqycjXaVNTm5d3uyn/tiS
usUUOXYX5DUm0COvE7xMAmGBbfk3314KzohtUq/VZeK7P/LbN6dDBKHzeIq7mi5f
IeAts85rIN51UC36YtxbPRG+8lMpMrvTu+zRwbOXLYl2V/7okoTPOV/GUCKoozyZ
XpbcB9YFoblh7BqPlBHEf14vA9WWLTA6A9YMp5HMCL02X1hl0KKJYoHLqvskNETd
uaK+lE/HcAndQDRt5s7LWVpIvV2Zu+VmAgzn7Rs0y+s0mtef+tKU37WqWb+sg8Fm
cOD50NkFhqE2WsNo6KEb4A/TF8Ke5pXgdi2h8nTtHheqTpasWD1FhN4mAb0w2K7I
g9QDzT4Ha/Jdab9F+3aJ9D0KMu2QnC4mmyJtXSTNTm1C/znuhQ+J5i7fI+AfUp7m
9bH/pLYt+bJlKBodXvDleVjxHO8xiLKZTRKe0JLExu4ss9xpEkL7GQSCKwgTAFk4
2U7w9EbPTLeP2Xn2O1fZRDDPpIMMCjwDK/1J5VeOTBuPD27Fv8jvKeS/35GXtGjz
bkhkNCk6QmGmrf4Jhv+aTN0bwAVjZxOxpycCaxuS+aqfHdYc0OwtPXUnAFLELrlx
vFQ2a43/hQK7UskXqc52FUtwPsiWT4U7F25h20sU+pETC5WfLy7GE3MVuemKqPA9
n1m+EPTba1u1RV3xO49/9mLjwNXidPOCxycZPlJtmkDqh2y03ajMGg02Cq8+zH3l
H3HYSe8f00032s6VogrbITtS8wnTM01haDVZnZcfwGaSXxZMVuP4zqbMShI5Xrjs
Quz/gvxtB3oZ7iv1Y8mYCiBwm7wFGspsb9A5vqxr3VIxSAcVyfoq+FzMtms/0eS0
j/kJhxt+8348zYN0YoxWxlWzOdg9y8I15ULB3AyTcx2WSAlktYuNsXXdfZZIf5cp
poz1gL5fblhMyBTAueRUcZPoigtApj4gXOTlGRITOkfYU07znRM05XeAabxoagrg
K9fSyWQ/kgsbAjqiwooYHt600/L6N2AEg8fK3dCzZtkfDoPd1GA9kACJEciK/i8c
Du38UoSuZJFqm2jyR/H1Qbmbk2Y+vdEeKI4ghOD/UsWKiFw3dnD60WI0Bl1qgSkn
VWdArsDJoHUUK7m5rFU0qsyuPLrKHVQlDERSbFy53MHK2SlMH29zNV1IJT27Jv0J
iwt5G/5aCUXPpd2NW6RrEgM/n8usygCMy/q4CHauemp2F1K+CZa8dmQRqS+vSU7U
O97AKuffsmZTZiRD1ME/aYfmfb5reiD4c5ALOz0QM1LPnzfIpIUCOaK6IiIHCZLS
ZCmVlC4ZdJ9OGilz+4Nmx8GIt6XUNwtyXtvrBrQsJwy9sUyS5qg9yRNZzhS8JDtS
LpmfdrZlArRbBLg4hk/qaHrLqYlb/K+iSLMumO6kpv7Cjjdacfa+Y6XS/snWmLXk
DdeKVGy9SYTijUs/ILc8O+bSDQmYCY9TPsDrm+kJpJDSPbhy5EBkkRQ/hlKS8R5y
A/7GxtrSdnM+fXiPtXBkNvi5CRHcBaRw47cW5fL4OKYqvWxBI0Q835/CaKV3Qayo
5iMsgS+JBirwMvia4AhRF/0ZaeTSFzfmQua6i7Oq+269im4mK83aqS1Pk4305/Cp
IF6TMbL0CQBCw63x1WtigzsPy4yfmvkzMKTgmUmykuMSENx9ug10JftqkHZD3AA6
9lCRQJ/+smIiUZABJRP8zbpkBtk+PZHzQVwRwhsfd7CaCNicC8kBdd4S6+TV9VEd
8aNeUvdBgvAOtp+AcUM0T9BN6jmrQjlygjO5n587slWMak1XWsNdB7ue/TIXa9fE
x+TYxyC0JW21kKuk1HIqCG+BGu5IDK4tirTAPaS//6usrD3I9ZwNGRB5GQbgR+uZ
RHLPU9sTxjdCnnjT6TAhnpYTTdZqXFPynk4zxUDeGvfXs1Mnh4tVGYMEcIhp3eDt
4qh1lrqgpPcGslMvRJuMaIToDZ7n2RqEWiiCdrZJUFO1Mn2GhARz9WL1hjUAfV9P
mOZ7waQp9qGudCEAjZre5Ugb9gsGNggd3WjYSFlKreW7DMQDG8DJzIBGKrUtNxL1
Vra+Jyx+9OB3bSNDL1lnimfhr97/zuyej6hFcs7GMIWVtL9LNoLw82DC/JJBxNH9
7sgV0hPbUgZ8lTVyWAbTHLWIm93PYGJPkQeKQtRaoWSAMw7lxikBsLzIDpYybXaB
MNQDjNtjbVonCA8QT2xuTKuUH32tUlqe7cQ+W/upZY/UtJstNB0Hz4GAMkIQ4zx1
ICv9+FAfiKWudOhPZoWNOa9h7cRXcOQNvMzKnsD5MkDsZw2OJRUq8Ef61B/vdRsT
dVWDvx/OEq7Da1v9+Qdj8nGQfh9lpuC7oxG3WTErYdALpz37O5JYO/r3t3WZ5W7y
efFgYYtDYnZBEAcR0ILk6p1mMYqZf56Qeqz0ImpQqMnkIeFu0R6fEiDzkWyLeuDn
24OdVkuW5LnambmpPSijNuJtGMIwdGyy+Fd0sH9aAk5fxBQ3GyJB8P7fSTP+ZC4L
66NQOsl8xSiZwLrkIVzxdpNw2wrC0h/4SaA/x+e0QfM5wiJjjHL1QMSAqljBFCz6
X+5mwL/vHTY0/jW6j5LVbHjEKjsmCSRFNjvdjbR+xn36k01fPII2bYF0lv8ZV1WK
KIezZ4GEpbRlvDt9nevC+KaUG93mm7tfonsz5mHtYKy6vExDqOxi/jWLcgY8T21e
Xp9tI/ACMQVbypPu+eNARwOs75sVK9NBHYnMwRybf7ocHgMiwIiu1zOPw8+cPPYN
HohTO9vNEaob1nPUZYTrEMPdqF7PAKn9e7V6DEl1crDFBzhi2XzGs/YDN+4eEIWe
vLWc9aGZJOQ4rdaMhEgIL2fCuGpo6clRhOkY4obhQhg/C2mVi3f1U+hqpAyDM/6Y
N/T/ZAxKrZoO5OM9UK15DeYJWuCpOKX480jWGXTmxDIGk6C2MgIigeOR5F154eb4
fU02h9k3+/iNRb4f7mgmnb6/5TQRXMDb7EDTSalhjaPJ2E6C4bJbwhgcJ5uLIqBb
iqnvcOBfUJPZtB2edYfupJSHKT/9HScxkWqeQANt95AOVe78ByKQX2J3YDOHClws
plf2EGjQFMZ9Yccz3CJQd1zZwcuRia1sb/VrGotV9aPq3GVF+G4qLHZ043vinTqC
v9tPXiXxl0gTkr5MT77jkiIhHLJg2HsJUTawGioMlhmsp69rUabhQEWZYrgY8jzm
qSS+iOmEF9ZvhF4h/kL1tEBXWdcKjwtc3icYZ/lICUMxgwkX+fX+PIm97VMm0uei
/FpDP+HaoAVsE05eL1hYNl4DhXyUManMkGt5+lPtrweiWAssuVMORdfaNVCE+g2+
QJplur2zeolRocciVpLliJfadV61JxGKoxHaJ7QJy/IM+3sa/pF4XWN/6/Etx1ct
RwIQj2/13Zi6afwn40q0VR0KmdHNSr60lyJxRbvijFZwfqD+Lml5JoAG8MicNm4V
XOVSHB3prStfX9eLrZkjk/L3fVEe0U1Hqvyo4jU9rI30Z77iWo+NF9n44cRzx8Az
5BPvL/2AeyEtVWDcT77XP1Z4d7Hx86d//PiYk7lUT6pWrrd185xLrjHpgRiBIgFg
Ly/kQCJSSPC0Ao2rvEHQI6beCW+ANUyXXdWNw4rpTH5VQwe6eHgPSbLha0cT9oBV
+GK7OBqH1zrHzbtMAv4jOs4ROAQg2PQfZ119dB8VnGoXMQCHSGsEpTO5wvu5pHOa
r779XJFHOazwxY8tx+CsV7thhbPH/FML2WFzSVTBFx4bCgThX42r9rCBdq/y7SFn
QsAzMc+9SeYDtO9d5hAv1kyHePHDI1e3Msn5jEaUGZWeg8fY31VUh0hgraWK1S2/
hsQfOXUKdRtRlEkyt2MriTRWmsui2pMJKqpspBYrKx0ArtGazu2JkjeDrmO6FRZi
3UcDOv9mtZpCgrSQYLhXa/gtqCOfd/ybVpDwL3Yu/AgF/bexXpQalx/ISbg+FBUz
ykNeLBTYj39kpBA8rbtnoxyw6cgNgoBKvgAd3wwo+wasVMlIdm1AuWvI5d+KGeZK
fPXNgVxoSoysXnCtK56NQmvrwRpAZOnCxnVqXYKLDOqmXU1m09NAYKSvX+Q1DGg7
mGf5BUJEkHt1ctqNbCkgd8vlk4vfMcbPg9GBtsUrUDuvfExarYLiDnGU/aCO+eq7
fr+KSndQkprxgnfyYnu15dmPusvuVcVQL0EtdQWquKYFRApM+DyP/FVX8Qroj5Cb
Worjq9JMje4DdkPnIIgSJj7swTXiRbzPe3FheboWde7harrCfXJxuo/RSV3PvT58
rSwdZs3F6mrYFhdIcjGNyeiB2Ddetvuy/vDe1f8jAGQnYA0ccqrIp04NThWd+oj0
6ttPAuEpMupMkqi3S7OQR0KGNv46o7Hn/rIoq+EjttCFIvtb1EizkRY6UVOqNp+m
1ec4AWVQRSRD0jaW6YXI6HS09p/jjFbntLIrfX6tWdAkJsx200JNlpop+STUn3vv
QhylVFFtSVdDosxK+cTy0sjrIGWW2DV4KSLLy+qEW6UmND/TnZt0h+NJRtv1FcIz
XKCQsJgNHEBNYlBIpnH2RFCWK54LJ+n8DjGGdTo05hQAWYI6XFhJc5A2SiVI4xOO
DxXAmCaHr4tUxbCimreXPMsUqP4oMgXVk8O479kfRCIUh1H00xWoG2uB9LQSfPe2
safJzLR/z25Eiu+E3xKuIh+goX2We+iQuGRajOrGosPzwd2P18FEGzD43YZYL6W0
lmJ2gBRoEWupaIKe+UFwQer8cyMnWXn4GQeZLo4VNavoArOGKXOsjvkwhhLQj241
rp/ISczMk1ZQm4HplWU2y5o/wQNl6Jzrmt21A76mN6r5E3VMpPvIoNJYZDbmdfhM
r4clrziuAm+9HjhZ9V7Bd8dpKDnFzwgQTq7AiwDe9HxW/3zLoYvz1svvOTV6DLN2
062n2uKgXYf44nKmyiqgLTz3TUkCWlOI12WKqbPWrBm0BXfqAmztwKsrUYF48c19
kMTCTXtbWT4cROQlDGDwT+PCg/RiozzgttSTRXAbT2c5RFb0b4bBMMJbr5GM00Wu
zs6zBhnimxJSXYqHbHyWRbA0qx3f4c++Jbqepd5iN46r7W6I+7QRh6gzyE8ANZQu
F5q5/UkqVUjKCM7PuEse1sPoUbkaY2WjDuJqiOiSUlOK4OSAf+CqzIsNV3tJQxiB
GL8mnjgkMAdYDad6ELg4Sxa/2zorPr41zQFgycf1stbBqwG5rWAl9bsT1pOO+ObT
Au3OUa45uwsokEb12XxDCXoDm7eBSAh/V6/PEnr7irpExz3P6Od8E6K4R8JuNq0e
VN+tSYm1SRTg3DTQYVYWf3xnmdXt4PUIg0c5j3RAcva35zFocFAiTcw7ukhJrnwd
m1UlJMmhO4qUotdX9UbNEEusRz7CuBQkxvhNonAk/X9i7pKxI5i6kcYr99yO3ZG5
AUfgjtdWs6c7Spa4cnzVM7ZMemD8y0MnZ4NylZ7p+Y4L6vvzGqEses7Beq/5BDQJ
zpQbbS1YZD76/PHQbkcpZRNndp0SP1lqsYy25iuAxtX8BmjL0OG1NfMNFCQNYt7b
1CPt9Z5YCNulmxAjOTH4UcPnZWE9OqRuAU+Na3VS8RDIfPUBg8XXz9jOSK4KUP98
lrbmxo6dcsFwRi1sVnOhi/nsXNzf9Gg2UDnqGHze23gPU/yFtrkT4AN60UGi6HwG
Wcl7BrO3DNjX9lCEu3iEx+w2UBV0a1Uu/P2tbXS6vsyMOCvSIZoeAOebyOQD/cuv
IuH3XC4Dd0oDB+pcebTvcbWkrz5aWqeL6LTtc6gsV7Ga/wDfGRN0GIbr9l15zL1k
c8S/FSZyWzDBzSIWnIqA6mf5dXpUr26x2UfvicI8sszBIpcTNlSIPyBuse4yJmU0
PfrWUEcdqEsipt2REsglFl1oI5hfSZGrdtGmzk23aIDM/tMOM6chdDsnHMBRK3FO
sSaQbfh2nLqr5BMXTR5b7miaI038gJKHWQnGhYuONscMcDfS3+H8Q3CG6M1NkCZN
EVJOBrBdVVohfby5kkFcWUm4ESZEQ/EjFYxIO0/unAvTM9p6cxEnc5NEzi8IqaYa
soy2ebxsQ1VqWFRz9UPispBS2Xo4OZmflRbxwtJOy5/FZKqhfc/WZY4NQqANaMfE
yVvCH9b7RKWcM+kR8VTHy7pVlq9HLAgkElv/o6d9Y/6RO3Gs/JLkfKh3ABCFYMYS
84MFFKBnyyDkfI+mxAcZwhUU5kS9Q365oZJlrpQ84NIA6JeCr0KTIpZYweMfUCzH
sS3DzDeYtd5mxUWuZKWPBhiRLmPvcwWkodKkFTN5xon35TIAW6vQmcCcopxEcCFp
lvyqiSV2i0T+KpIABDKzgJsCK6GGHDZfzVsaZj8k4apwCAwAEsfwUzWwwzWJ14bh
C/RitoP7JItk9IpNmi6TiS2n80jRnLLZSpCFodzoC+RTHAc76pLe6mDk2ABYEBmD
KfbKCeKN10N+I9Kkj3oiPPDMFYG/euaJ2CBkBvPDnHUPajZ9lb+W2UrHVEajoJNb
9T1Yi06xwKtzf8cIxCSgZETxt+4Hdk8w8iq82LPpVxygS17Zy+PFG9e01Vfz2uwC
Wxce4zLF0LGWp13pdtnKbdq3L+d/hQynno0C9M0goOX5C293kirLkFriXyWxK5Gc
9bsGH/UrfaMGPd6G4QOneoxOknRQORIyUo9iNcx1271VzPPFxnC1RjJy5Vv4jpC1
RfKf7oQfhsuurCp3tiEyaN8ParaIXjJjtvxU6/9aGIXfakvysbwb9sNsbu9eEbCe
+99eXHJ5bxLBRMZKSiacNIfw6C22hQUpOfJq7SvZiVOl4Yf96LG1DoipkzFwXUIT
T+X2uOJVzyrins3yH4aQjaT19izXlS7nd2Ne4ZTOweKLjQzEvm5mlh5xn7eIn2S1
VAEqEmCGAs5nbENNlKeJ5g8yjFaWlQizguzWpbeGdmIMLcFx+A6WcmZy0GRzZbpx
npXrmXl6dKes1qUpmpLU29lOTKqw7KKOxZPKdzruB2eUY+h47FHCPp+ZaV46Fyet
gdAix3mVO2p+prq8uIZ/H7sUBp3bARMmsOpjx7tC82Wiox8QSPnim9vIkyv6JOtB
v+rJU1n0dsJVjaV5CmcubTNrFIC2qpGrL6ANK484JZCYGJhK7eiWT+meptNq1a6q
5kxe8uAKOzJnwFbRTLD6bqSJlvJIzDHCUCWtqFDSDDoW+QKJoOlIFVhQCzUEKGHs
X6d5087NtIqzvLh5E0Z8bio+HKrHVxnqfwjGa/hX4rR4GZvGNAlzOBYNNHhpax4O
nXk5DIPoKI234dXnuLuFk9AZ8M8KgVax9NTKwehapdF/CwdHT5B9yBVWCx+wH/27
CGVN5vjRxO4pA1i3vWtHjsjz26v6VtT0jMf220vxRf9W2UGf/2Z1u05eKXmqC6nI
cFhhkIeqrzAMIPArAmriRFM/NLGn6tBAoX/4uz5u6lR4iRN36cf774ivLN7Ahe7S
TaQiWuiP2czj1AHsW6sTBjGwQZjXL3K0kRuUwjHC9FMcgWNW6lcfVo/J2hDdKfc0
3T8LPhjwD7vLs7sdXowMJA+lAyDsL6/7BKJyIvCjHYqyhHKCuVCwD/byphSxxGvc
rh/OuwhOAufe0HDgt3sFmEeL8TlfeHepbo8plRnupc4tWsix1+HNHd1iShADvgN2
PinEdT9glGdcezmScpcNtpakoHEetagI5ruSbGD6sclpzxbcZy3UoXxZC05qOROq
tKrTj5VYoCa7EsD3cxbzrj6mE/N9a8vdDB84LSYoooWP6GvktlKvXp9kvYgyWJbi
pDOaPWjDxIhFH5WTSmZSkAhvwuxZDYRP3MlP0XAnqHxZ6q5nXbFH/Qa0q+BncrOM
3RL6scpzPonpgXRI35998LlcBHGnpZraWuwFabFGFbEIvzbHUi4pzyv7p0O/6MHQ
bT6RryAlNMUkvqb+E9SK4bPA906A8fHzRghj2SM1ydLHHbc6t9S8J1lWB0kdkvSO
LT8+e51mcp2Tekm/HmgJM1bu75tfAHGWFIb6EwwU562c7hBYMz1/NFFBXuVk+kD8
qNoSJ10b2DHiTXZHaQ4u7we22RUv14usBtfCJXi7dg3I4KvET+DDi8DFBCokBloK
sPQkBhqiv8U557TRRROtDkXuWep+QMt7iKUkoBOZeCrE2k3p2EL15WUQnlPNpo13
223jMrJRJ4fVkXDm9zNpLP+NqAmoG1gWEqFBLf9QD8sQf+lR+wT6vpG/7gDJAhQV
l2O6pAKme4vBDhpzzKB68UHcrfPQcVvb3JHKlx9FQTtgAGMrTHSkhzGJVf9xtsxI
3+cu+ro+xVuJNg7jGWwWPN6DBd8rdyKIdZB9qWSQKW+o2LfHltfmSFFrfkCw9og5
sMC7pMXwZJGDccz007M1qufydYw/1czTl00aAIvq+8qhODxTV9qk3JJO+i9LiAMO
FXLxiP2jdtfJKSQNoVEczGcn2W05m+FKv/wb6amvUiVZp6rUi1Z+awKIyMHZuYli
/7Bb+8ddPwE/hsuwgVvf/XG0NR/RUCNc5v3jOerBSiT8HUqAEilmcHZElPdZSP+S
eGtsySDLSnNoDEK7xtcqbCibmBtn42FZbwmdPfKzwyiuZEyy3/YHy9ZZTmDVxBgJ
zoe271qkKM6vPndwCFhBBqjs8/itnWF8aCnC8wZU8HxS5UgW68/EqknoeATgpEW7
euM6NLp7jU80xbhGL6he0g2Oq7gXupOWVH535KKC583IISmTOkOcm/uAHsAIiuaF
w9cxlwfKLZHcbBxWdNPt2R/MTM7DzhmwXCRePTmhS7yOKW9v1HCxBq86XZj2Pwkn
KlJWMJKoNdRngZzUO5elKteSVQFxtzopG1MbhyEtWnTgQXHyzPzBQsPh6D4ReGnI
ietcDV5+l5a4lw9NgJiad1yLHDTEx/8AGqk9VTaoLNSSUZ8Eq6tnWe79lk/3Hin9
sqf9B4eKR12nXZKlSwDiz66vRCkGr6BZgzKCZZYcjkv1zVZHm8B1ymJP3VhoMOeT
wAhw3pXnJXYdbtNomqgvlOhuZWT9/Y2jsuBfshqJaCq8+NJd6sF0Gg1jeFX2SPL+
MkMWKnBxt0/9iRkF2nA9VrpCl1qKNTTL5YPj4CpH8DyTmJZBmRu2klvghjwrFxSN
toqv64xS7aw6QpkM1y3bbelqsAN5BDEw/17dj+eCMoKKxX2dWn2iQ8cNaZd7zk9W
nT/wsUsJuRWGZTecz/rgQ7JKqXQ7iGZxFABpxRTeu77aRa2xZ5q5dSgnlCesj+uj
m2EjjBmUUZaOlQoVX8gQFaGkPHVEuB48a8uNJZvcfa2wO1u59CMdiIbWyo0RHqmz
kWJdTrJ4rw15wTsyPnL4jFRhFGvbE4iafGvHQTFGZwtb4hhGCBEyMIdFPvQ7CBPo
QxzyPjmtlFog8pHtAcSFm8WrmASUb24J0e4Smfz2A+gSaHId7bOTdLJrfAYfMciU
EhZmjvMDXPgME4SVGlufQpL2Vx3MrBGCkMzA1hNpJGnbLags4wUcZb2ZN4RCyWvB
edXUC5jChH/+Yh9DU7keOj+5eQ2s0cx8jwXUKU/Q+ZTh+JHc9dnnlkdqzPPNrpJH
aWjJm3rnSWW8M9pMzKQIC0FL6UuBaxQ+Yw00Fu1yvMFsZ1TDFWyz+b515poe2NBr
2BUU8dTjI/2teG7s25Mnj8KABb4bJeesvmus8lYv1bMj5964EcsPiRsEsvXZ14nk
Sd5vUAJKlSL/5ps27lcLxCV3Tz1IYHygk93s0MEBZ4wVf4s+B3+uQ2o4JdJ9u4Pz
gS8R8dbtnBux6DpsR5w4e2RriKaKG5Nyyt32UR5HLmYAYDZk9hoyeiHjA51Wy7XL
byjLiJat8XinDLbSUAAETDT/WkWE45x+VpQazWkkpVZDiaChgtXhljYNIvYxu5gb
70JMgdSK7iALiVB9wcm02PrECsyYKcIUslNx5Con/29rz63BY8WZ0oO0urozpFWZ
GY/r6kCoCEch8onDIT4fadzGNzNUJ9U1o8sXOPzZqxvGy0WAvRDcO4N0w9l9CgTs
u9sYUHGW5cJiujaRU95fC3T34QNerKwCSv9D5zNKSc3oUhRNZspZsOKY3+lqZDr3
lzYdcpTVUnWvNV8Q4EaE7ibFvVG3B4yKGrO5sR1+7KY32P8gWe6UX4qsN1qTFaMZ
uuri5BfE3HGV55c+xDTkKHe/vs174SaOlcYQx0OuznhtAVV5qAGVP0VvPYzKOGV5
Lr7cAnD3Th7SJF77ehOToOOftXd66GQpE1RylB89sHhR8xrRlASwrJ1SCK4IWonV
nT3LMADxRosNqPBZEv5CVrSrr9WFomeu0S9K6VvH3dbyeQ8WKMlST8gQ7ekPk/+b
eSBOW0rOcuaQ5c16XrA7BLvE5rPMq4Es9cSbfDPAbkmVPhM3Jmd7u5aAoiOcdi8l
/pULOQI/Y0ep9A2nq5XdjFyHOuMjA2gjdYEqzqkahz54PYPU1NY1P90U9ss+swGi
eCV9GT907rumwHmMkyQL1d2Yo3u9lQsIcZMFsuyoQrZq86Qy0I774XUzB/Z4Kxgx
jDDYI7kJr576ZfSHTqLejtt+dD9nZl03RplGt4z0fHk6pN3G6KANeYpY+DNHGNwF
5rnLjbZW/FfcWy9RBcFaAKTCWF/deT3Kqg4ERCAGkWdcMWoBwWcds25bFXcWczje
LWbhZcI5G1X4Hk/L6jOY5dQfgthirO0p3HOL+5IHDZSEKpb5IgDzJMINd8YIboGJ
OMxpAT4uhOoYdHgXRvKtgPMxJ7tczErD7dePaYNYpWj+sKL89NwJV9NWaDF3uKV4
msDZJvSScuSfLZthwvX2vIWpqTSta0TR+PMkyxokaA0aFQKT43zE8w6XbI1i/7DQ
Ppd0ZBQ2ZdBvykOWrhwiEwCkwee7hFaWLHw7/a090oGxB6uLBXfTApQ+cuogI69s
zcTTWo3rmbAY2PaI1/RA4R7v1fiJC51s+TE7XZ8bQSGoeLqNTC0S5M0dVil/GZH4
Q0Jg/1M1GV+QLZ1oZp1EkoE++UQPP4K/90eNI65G6QgiulverVhwdUuPdr3Cixx7
Ti8yc1IFky5UTewJ9mkeAfehm9tyoF35QV0NDA5FlD21VtgHdG1ATYIKZEOx0b0i
ez69DLhNX2FomOTvsf6VaCbNxCGVLVO4+9tsaHs2+kpZPyfuEpE7hd/TFHByaLiJ
WowTtGLQEQifvgR0/F39Hdbxo3C3Oz9nYNXl4EywAR8FbIZVkRqrfABTDyer6oHF
/l6bj8JXEyBv7cYUbjDlketit6uly0pU4s9gXX3ZyqWf2Ge4+Hp+z6AnCeJlplgw
98femL4zUwaGq17y1SLqmX6EkzeqDRoyRgIqoaAw+bzaLzX1OaPQt5x0EkQGwtqJ
L7Td3YtAKEe4+IYJginPi/DZ7q1reBDhbJnhVSsRSP2+OR650xo3AG0pQQakBvxO
cIR564+WZtYrUNCFC/kgIK+T9JneP1IduZPDIyQFrO6DNiYMN75jOKIRnUWdSuM4
Vb4m2xveOYPKcHBku4g1miOPsCvnczCE/YWjJrnlvyG1Eyc3JVQI00lFkGFu5zOb
qT3kzpKllWOgJdhaZbQtEIcbpwo02nmthRga3q9SUiwluXmCx41GIZNLZAbWmF1J
WBPVzQC6XfADfvaxjAf3zGdIvfxsUC47WRc4xuwxQauTcN2IQol+rgDfwFY5p9Yg
G0JBlYtr4o5tQ5tbJrRRNgTA/1ix9Dgj9mqS+nVWX+h8AA9vBdXd/kAGkmiWiUu2
uuhE7fsXJzXlMbUz5gCQx6F8bfm4U6ei8teUqvevVXyaftxQF3gPBPUESX3e15eg
5S/kq3Op2rNnS2pEXDllg2cmhjtZsPw+n+iII/mkAiFOtSgIC3w5tRdIK/cw4SVR
Grx/4kpD3zlUp+nlQrv3k3v4DgJgrgm9xJbtRlfy4UtTTTe1/+qRlaDzyLn7Q1BZ
9T+JVRvnHx0/z2txFAqa7wagqJQ3cx33T4JW2kUmLsZKLOweuQ1PcGQcm7fGV6eL
eDgufauaUW7SkgIYhsZyNLlT0Muc/HuyE1n4qCtTKUPKhwI8Loxm8OdNIceat2zr
H0OCE5tEvYTCpgVZe1ESTww+SwhI7nDVRUvWxH//+xoK5+5uTVqbXFiUb0u4zr5x
/NwN2UXf8n4LaWetoQj4IuUr7RCiF0wUkIvw6SNIViJEblxzei58uVqw0+Du8B2+
B6qJhKSTnjevycWXgwQJjg7T3WZqqCnuG/TecsRZkpjBzC8px5Y5MlWZA4x8CnRt
R6ev6DUv1B1xO5vkfZqiBd78VtayVplfqQORisvqAPxEAWCgQYzHL34bEcKGlD4E
dix6tuinM3XFPJBwizb9q0dMSBQJFhigFhR9l5/S7jPxs/IK2rHamXC2OC5m8+k+
g+cXU3QFdiKscviPR492zaKi26+AoTzDyfICWzeszTs3F3czq/aul7rCwHdYvsxd
HW35qPi9J9FuEI+E/hZhDiJqilPSmpRfbiz8MQ5fB/jytEUiFUBgORLjjknfDhtP
zLVwcrp10dmr52lSdSslqhO9N9QKvJ8qQsxrlubZSKVqH4acV02160z4PRs4rAmm
YJdae4bD3kfwkLcaSya+0sOkUXBL4d7RuCsZ08NfDzcB5n5+cR301aTfXCm5vwyb
pJ5IxtLOuh6iSeDGeQ/08q0jGinriWpNUyJ9JEKhRhoPj4otdBj0NPSKCxgEbKSx
o4qZH+LALqh9TgX23xUpTF0iclLSLtprnnFw0oh7Tj+REpw82kkfr5ef19gG4IOq
/xGKdB5BZhIbTy6x++VimqPGN9fvmDLZal9+e9qXinviO0JRGwdBdt+nkRyXqjte
GRCbFJmpitYPn7EvZki2H0hgYTkwkR+NCkSwMQVcIjR1w8AOnnLhE21T65aWyiu4
c/fZqOM86zlX9I+PRW7j10G3cBNKsQxU6oOQSEAIAU0CHlyimc2sSm7vLlQ6/Vw6
rPoDplxvS5BoOylA/cUEPtWxVM7vYUt6jv2rD92XwYMb7nLvWfu9YgVKkwtnYoNq
osItOzjtN6SCKqU8r5BImB7YXdmOeq+WApKG/7JYmhNyD7cbXjNFhzN5OrPq0W7Z
glJu7TTluHdLdnj5berdhz3QWsRHMBSlzcsHtknL5W5kYqG673Bl/KnVO9lxBoD/
ZVOUG9Iwerk2wxVeghiYWcyvjfMyQeN7pJt9LRKtW8gnG6D+VnPKPrncLWHSph/m
tUcu7rvNOSRBZAR+KIih48RpP8uE/brQq2eP39tnf4CEcj95SA2n6SxOX+34kpWi
UfNbskLU1uUA2M2SyWiv7St4Eig8zmoGypUNCtRkyQTjYegi9mjqG6731hf0vyUD
DgFO2f8iQQz7C6lBiN2jcszmEPyenn3j4Td17vtKJIkEMciOCPmqh5opz4ORf+ZW
0n6gt9HgQo5TVhaF8O2GW8lHty2EoEADwkZwpsi/OttGPMiAYyaqxI2lCDOr3IA6
IxN5T9sL5gqDEAhtfau+I1Lr7fkrtTLYsBgpbHTJvVUiIOem2+HcISwElB/kmfJi
dKVXxHf6hJWjYRIJReKyglydXk3eMAdaaPMy9HDmKXUsa/xEZwArSdU+HbhejdFO
Vrb5XN1BbtZgS/alh4PRbUar1803fIbpb4MMJHk2rX4C+sRJ20lDzerUmrFievan
f2yZs6HNPnXzeTuzgoXu5WcIXf5xfdg2e0EQbu/oTlSNGXgXIUGOaU9S8IeqTCtX
JInySU+vpv5oOik8rhKYHI3l0gPk3jTPppNMVn6BsYMN7oSE6vQ86HEuuBX/yXcu
fQfnhc7zBWzzOvAfS8AjqMMxsbpTj3WKk32NN//BNzmPKw3z3FHNw2KlA3afZ+lv
UMFsZQS9xseU+5zwSZlxe6p2sGmq0QthaDgcnjaJabNQQRCr0eSJhKUQeAEidEp8
MPiDL2V7OEDlA3XDnQJShWdNTjSWitElR6wuuWHWlTw/G5gaRBLBIMg+f86HtVuk
5vCeO4nFn37Dw2SHZcLuEttallTKIIDtMi1I22E0Zyp35xOfDrT4fJ43elkx7mqK
iWKLWwpb+KaeE3eLnYyZI4J9bRGSj7X+Zf9+DIMpJTNVCRBFaph8SFSbni+IFISZ
pn4ugXEUdizcReZ0DGgIh6Z41n21cp9k87HR3Y7VVBnPT3+3oFAvS4Us3WL4UCO7
F+TWmN68Lkp2ZMsZkHixpJ7QgEyapbLKWYNC/PkoMHqRPZtGpJXZ3yKXzg3yVXyw
Awyf0uaAm8Gv410TUAEmAX9I2GY1yBpvODpT2LIwOixwLu2T5JHfhWb14/1qBkNG
1HLP7Vo+Ilu11GQW3kiSAmr+n+rTtlE6vQPjWGQI6L2r82ChcZnOblEWzwTvLzsy
VEahCsLaqHlPYCv19DlEyudVbQ/6ukCrzescxT4GGKko9sh1gx25B6FRB8KrleoF
uW/ynZMrysYDxUG9VBlib0UiOktJNKrqmTOaZMm821vW34aRzjxny1DGjj4BW/MP
19RkRaclyAXVNp3g0h4gmBoVdAjPFth6gVXcYU0RDTqFEes8T5zhIfvGTvF5qBJU
Z7ck9wnVY5OfZmvctaXCKrBTKACOGqKTxg5hgItsNXpxkmYX1huA+nMYB8lOaKbi
hUCVM1z54bAMk3OmSKhan+RxxoJ4UMy0wdGad5B1TrJ8+k0Qp1/idnl7iEzi7lGe
pXUwd2idbsaylAyuZ2AkFjY22rrLJoam0kjHTLwDSnod0sXzd4JOz1iq/t3jwy6m
TRz4JybBuglDjryK50dvSn4y/HMOs/XnRBL0W8AkV8I+cMIXwEN6CaFREZHUoMpR
xvnppHroA3yhe2eVZUGyEGBbVrlw5j8nNgQvtQHQOhtiralkKjvegYFzfqGbX0Ax
qV1sFUJ3ueQtMM6F5k7Zt2sYYh6G61OxIInrCsY5snw990Q5dU6tsJr5RgOw9E16
ZUUeJiPfppMFvZs2Di40UN2PyujbqXPimt14xZ+c38zfpHfShhHSQ3RL6eP5cPrB
/u7Oi4QTmfZ/13Nk2u3yGlafjoqADj7IbRWUvOYpgwJdjdvvSuDonOJIXHFlAS+a
h3p75IgjqKHurgbhT4DCUGXEpIhxUW7oNhEzaQpyQHUXvYcVIS5TDgm0NoS4DDKV
j6GetSUPnUOM35keBcqJM+vbF2BdklIo8fqxmeSI8QoR/FsEwetOc/yRr++Za4Vq
VSIS3NTxqSeVJV+Ifj6ss0f5vZXcvPZGAyfozJYb+rj61umkPKqlc7OwX8yLdL4r
dQY8UyH3zt0M2wtDBVPD3tUkz0x24Gn9URyM3DSgyy8WOSN4TB6s2gw33ruHZjnT
KglFnqp+SmQuBxrZj3BbD5GuFQXcHzXxFb6/U8+mPYsqkW61m44nXoMB4srGaJQ+
EUMIrMXeWjb8v4AghhWPVrnwkSTElTTZ1nVJxFNYtzHcvzMfF4aEWkB39LJxi+JT
csHvL4L8FAC40crUpA/eA34ogiYL4zWeEn9M2/BJ8GigHL5db0Rw6v8+VOaT8Yqf
flHVtQPNFfsb5w5/HQaaAOQYZ1oAjBq2ZWwsMRD/dUd5b/Vom8rBh09f7A5FF9vv
UWycDG3ZMhUkz7kjsFPFFVg3lTliJPuVVuWP9ipbzsIX8AdBc11kSUh+ynTqkv7D
ny7A+vavYM4CAE5QYM+dK5JOFheOWEUOMox/DxYXawUoq5JTplh4PCI4ElTzGQFb
N5TFB5m+bkK8Ht/JhzrQGKl4dq0PjuA6LyzkbXzZ+eoyR/lIKCe7w9L6elV+KsXD
U9p/MCoJzeEKiIQm1WQ26A/+944I/iXLdTP2GRqmG23+h4Y4GtNCr75ebfagR1rb
sn4l6GTrwOSNfYupaIOLNktJ4EiReeMdDaXyFdlOurpWqBDGKmvo/fMWnkD4csKw
TG9WwVoJ+0Xtpl2lIWSNXI8JdcAW20w685wh9AZN2lDZ6ttbakX0Ve9tQ8lMXKtT
R985xWms8pg2M51NzQQRn38A0pLVDel/stQ02KNDz83MDljQ/Od7DF4vu2rppT6W
Vps+w4L9nbcpJvA7lItJz8nM7kDHpazbQ8H97MACWpBzEVjebUX6l9h2GBr2A0Jd
ROP7nGbjqhurfmMWl7LjOLkEqshlHzn4DWP2xkbVs8Jec2tz8QgOEf8My+KN01h0
PguDnWECSAhQ/qS6i59ikcxcZquIw7NAFQvRyL7MSNPTDBiblZqyBziu+14AdrqP
1CeS7GSisnXQZVUcQ8dxigP7P9HdC5H+dYkPB9WP/5Lty6yeSFCBX4hXnBoU8Ko6
UDlJnOeb5/Gpx5QE0gLmF5BT9MqJzQz0sOV0lg22zct4iw3mbeWOimeQAWDDEqyM
bzvnnIONIws7wG6iR/RSvaPKXQQPnukklkiRKcss3A1FaAU8iVK4yOsMM7OO1loY
9RIt6le/YUU9eXVanb/xHo4xNxXz7mTdIG8vZrxmFgjebQ/1e4Q4zGyukJmoKt0g
MM0KVX2xLsVXQgKhj/WIhx/wEowtNS3dVcUvmSpZB2pWCU7dRdtOSjH/htg6iIcc
qOYQK69jhkFbDuamIIB3CekfFpU/UT/+a3kmK7coKdwJohks0Hcgo1hlKXLsWnnO
SBIxsONsdsoCFFXIMkhgdrbt8Vd+JgXWdQgemqQP96hGGF4vGi1HSk9RwTlQ4MF/
5EFASXesvtPN/K5eb1iJQ3lsPnHNA/HdBizaxdRrf4iWQi/3paGlqiYJHdE0eEAu
C/3+0ssipakgZhWbtAxGJsLWRs9PrLZ+0aqZT9miTJQMfsvO/s+Gk8/ijE2G5pis
KqsEzxYjAEZIXWcfpEaYLGlP2QBncPMQNA0UnRnCGT7ZVcGeMv9VqKi3OWroKvCg
MEirELmdRj0MxcDQg52ONKuGhA3kFSEmCbN+USqfsDuB2Zgvm6sRLsJSW3A1lm5n
EaK6VLmGP92fvnM6DV9PN9XaiLWi5/fpmA7tyszDYYzB/xZ9XeBqCvottx66REin
FA4/GsUM79Fb37Xxdz6ZJLR/ZV7M/6iKPdlQyUS0YxqhoQgdbhNSnrda/pNIs7Aq
hxL+/g6YA6mHv7bou/x8wB9x8STeT/eMZH/xd7BUD9D4DpkiV5yqOOnKW44YFl1I
hhTcUpp8MIgFiu0oKT+aL7Iftm2NyOgsGz9X8+w1JPJnsRoN4pdKUfhUUHXVqG5U
ZPdsZk5lu6e5QMM4CUJmOPRUtTQ9qqFeBDOPLOxlJSNgtG6Rm5lGQZDL1EgyzQ9/
N+Obvy6jc6g+AA+TdUXCb9g+0ffHSlkgVIcVdwGfy+ryolnx0m1CX0SSouUamOg0
wXUSYMjU/cBZvPxVw+nuB4z8+f+3L5bbRKKnXiLlZ5071wla0++k2JTob1KgSiPb
QKB0IY+O8d7qEKVXmBSucUeUanw+81Dv6mcL0JlEzyPrgJzXBbaJmH9q0zQnXtHQ
bJacFFZHekjZxj53Zkpk4yE1fhG/GOhLfR0IJFFEXenXzHnJobg9+hIGE0xMOObK
FEEZGEYONERVahgeeMqjf6+fTdIo7Z9gIuolmOlfX29TdSWCOwA8EBfZiuLHos9Z
xMh/GuDYsU4PNc7CiPZswQoQ2ueBVpVf/LPsIjnFqdHgu2de/CcrD34Ujeh0VOoi
DgRqL0vwwm6BZ/bS3/A0ITRKwDO9MCacNDxfVFaeUXyLydQQu6HFXehw54qkvjTQ
0muGrzlWN2JZ+UmNUzUR5zuu7q91yo3YbKKdM/f2Z7GxzY2qZbBidplTfABOaecA
ux0oCUsWIX36dnsDTniLCIEAYKXclfPNhmclAREbxozxEoZk5sgWhINrfBjr2UML
APFhPm4eeAcZFvk63wVcKEJRvM0EyvXyO5rXBRybw5apMbIaoGK8s1ciQricUoOZ
/pgiZIEqjYWxavg+Br81LGnm0AKKxDTmQ02THo+moOSt9pnuM0oE5orQFKwwG8UF
Rn9n39Ia+cCzIOOowNz4cloKbOgONWDbgN/hECfxU7ay1wKA814VJm9in9LBypNk
edXboLr1BkDMmJX0NffInG/VCwemu9kLZcYrmA2eOAgYay51nhHfwtiHMXwzP8qw
cih2JP89rYlup4uZD27ItvBrz4V5wWKMWrcVbd8C3DYtNZOh9xBqYaciQlD3UHrU
e9uXMT6bP2MomANigXT/QS5GvpfAXPs80Pt8oYydQmglNvK2D8f5jM/YbqDTrq5D
xLVwdd6xdU4K4pwx2C8yBL7cmI2y6C7hnMppJVWD05w83o6iTPop3filzb4qdkgf
D2/UQmYDGiUJRx9Uj3/gbMzswPdgUSMAyp55byHsgBwx4NSZqn2tonSJvXk+f+jd
66yIV0XvCm1LSVvvyQmpArfuISGEVpuzfIaw7wcopJKZSdfKCIbhBWP7qChvXa4Q
IuLH9Lu3KvlmbTFkIEhDuno47qIV0YUSGcZrUT1mU1MbtCV2rif2TSo81Jm0eM5L
1EBmhRTo0jGewdyZ7czIbZQXNELdZ+1HgnGFWjrt6BoddcA77iNERVxABSgjyvnS
OhpgfO6hNDOIpdgStlAxo6DiKIi5AJf8AcBz+PjEgjiMGm8DeB+ywEkd63CoKuZj
y9YU2j3d7mSELsYhK97AgSXlIYb5Ev+5bFXGKAIGDoGo/e6DvYWwKF/BafaFlYby
4V+pTqnjQtk99Fmf42xhlsxbnTZ8XHe3jawPCC3G0naYvDrxoW+SRECP2vkNrcSN
m573lnIwDXYQJWONVCi0lSUcVdodeFe66yW3cheFDNWxRd27yBmNOnkBSmuJvzF0
R+gp7uxNDHghPUQCUONb4zPPikWfKlqbZ2JuRqFO5NUHSo6DPHsWpAzijdJ4WRHm
P0bTbktPy/KMOzeevXWFQ+H8fLsqmxBLTsG/ocYEdpM5BAHMiuJvjoL3NSNW1XoX
Zb3D9SAbexcB440TAX/QuB4+C5wdQ9iGMkBW7hOZtZMVLmybj98NaittCUHBcvCF
FkCc10poEtCMcFaSaeuPjPI0/bARyE3+HO+WIADvJFWca3qtR73p27JNLDDs/bGh
osUBPowo314FlHUTl0ThhS9F6xvd2uaV0ycGbJ1YXOG7IHh9BPticCMxZT5ZdtfS
Jr1l54f0NRkk8+G1G5H1sHqJ+wqpkqaCfE3kO+BxtCAV1Rc09ZWxrLtxL3dAf351
Ljm13NK9QIl/QpPhUpjD91B4qMvy6bvI5/RpANsYNBvvjPxgcU2hlsb6VtJkzv3z
AL8thdkIcWCJqyd5JA7ZuANai0iituXOr+D5asqZgSF1a1wwEGl52ncvVGKjyLfX
Xr0btmEHiKBabL35h2kqsvXjpKai+tamWrvaqbu9IeQ0bcaCFI1PQ8JG9Iv+El/7
LoRky5ofTFYLeoGSyjtFg5Jj1yxUNu4TjwiLSQ3ua65rGFWTicutIs6OsdHxnBA9
g7PnNoah2vZw0PyhAf+x74+gCc7c+mDrH7mZmOWoxJZROBn4l5A7TrBkdXNoyRQj
wK8kKiLURMujD0WdP3Hhj39KoijiXqwwKJx53JRHLJA2CFPugqvG3HQj4prAOdA8
KvwA71a/udA+7G+3wB0SFPH/BgV1kdpuz6jwzgpT1neZZooMP27xYnowmIXEjN8+
E747oMXxPwE2fIuvdAA2IadK1ppu8weSDZFz1AlZLpRCqD+HaQ3zDEitZDw5tRya
MiMqWqAM/TU0xXqxWt+yejK9FLPipqedFWwn+x02bEHQ9YhzPBbxSL48T7GZNmjN
C+FDAkEpkQd9CK0aeReoWVtthvMN7B0+tmZDStu+NPRhZ8VrtHMzjXb80uY4pVZx
CVpajnQS8a59HygKSrQQ1n5yQeN3FB1wfgOVeG2nD6Rgc3RZqduytykUNA8k9SKD
1v5kkCZ4xrnu1ISsmEqNQCQjPXr08HTFTd1rILeAMPjxWACtNNxocz6ULAXVBXnP
kMWuDsN/doo9707bFp5+SNylZdRE25/+3pM/jzIeULKdeAUmvY/Lr6VCv/xAOr65
mG6/+KhNdEtZ2XOU5Kh1Rnv4LI9pqv87PIlMUI6WvgwOkWCmC+L/PdmtG1hL4qnn
zIdWa6WgARQ9+luvxpOf+BGhaY/74AsG49ZhQ9zM6GqVnb248FFr95ct+kJmgMTY
wTj1LaAVY7eq7M97WV4GeORnoHhJzgx2Hm3fHWhZR4E/9bKduaF96ZfBU5csbcot
UOILEqHo+b5y48Riy8DIEgh1DFPvWJwidw1LYqtjO1oZVxOVR8vDDVvHn78STvSW
jpNM2hOJVldV0nSQ6ZrmOCaH+p2ii0DcA79dPOrIjDRFD1PHSFFP2BwnE5rW4SK/
fi5YeVRIBERwB4Mol9g78YSgmBE9PsojTov6OOzA65hcPGZq02CcffG3J/mLPfAV
2bNlNxxVcJJ/tjzbNhwkBsiIuUMNqfzhTyxryTwLB/CUSNa/8PcPbPIPzDcCHKEv
BvAoS9cAbGNMph+ynhmdsahvHKmUJU8ZlkEfQD1MECaGvsubKpPMQ9QTiizBhKE0
gK8IdhowzKmmw7lpPIyrfri/OVDObICl5Eg+IrlYwhdX2OCEPi0GJs1a/l6twfcu
bw+s9B5wGXTbT9Z9a3+6Um83O3AevnUSPQS82YZ+IHtUVevPca+sECNhGNafFlv+
1trqOUQofv/3uFDQKrTCEgvLcn4hDGG8Y5ePSrolDIdZv+fqBLmrbM/VlPJQMEiE
OVhfAdB3VYbsHIZSABZh7JGzLv3X0UX5p9HM7vRJpe3uf3CcfdYjmoScJCZz8DTX
DKOUTOQYQ3ud6T2rnq6VQ4rxdcWpdh67kCm+VCIMYb4f4IezJevYbor5iGANrmXU
apk+Dy9/nkctW7HESieRofoLKMaJYv6VVIR9rR/mFuSKX9OTd086CZf8irw5AkDL
OYkftODsGd9iSjZA8uTTmhydj59ISPix7U3EMAjnV3FrSNK5lX36OBZtuRqXqHQs
qvfqUBs8UGozVaf2NQc4K4d8/9BGbyK45WcKbIUSSBXGzFOp2oNU6vbzelp8L+VU
It0FB+M/iWDnCmOOHyb8pE0bPAYGeTbRZaSNU2gJ8gGQSdARml9uhPCgfrNWbaNH
/wtZJLr1xARnYGvhl9zrrQ8Gjje5UWLpPPpMbXwvkNAmuw6khrbE/tYHMUwaCvJE
kvtiy2L6xjzOydhuIK0wvJz3Ylaw5is6nMf+OrKK4vmeAfzqSJP14G/PUNo3GJcj
EgaYM90bYakZHN1rCjty+AeBJnAHqOnig63oBWSfEfubpJG9bZjLbiVxI2gbhHTo
blxM8rGXSJh68kaXKjuyyBUTc8ZzEEvlDOoFkQjB4BwwKk/+zwT9859miNumusk1
4Cq8GFn2gpfio4ZziA96YjhvCGPGwEAY5TnnJh69zAEJ35A0FRPmzAKK6REyeLLN
dKXZU6Gzt9DedwUf/kFbDrLxOmePBmqHeCvIFl3RyfLf97tGkRNk1DhG9b+OJm+P
9x1KofyY7TWQ4yRJIyJlwis5ANjqKAoBcsPYzxZ85J1VQHc1YhexabxkKPQZKVB1
e2HcNM3MSQkGbOr5H0+e7fcWBtk4grx3I8Sr0FzZDEmdXYAQqWrvKW3w4hRw0G6D
5y2Lvwjtnz4PP4L4PJhP7A+nhuowSrWeZVKMeDTL1jVK1IlG7uOdC9A4JB3QOX1n
7muBvAXgh5SjQuQtnkFScFAm9NjW2N445thfwRnP/7yDEFiMmgjoySywc8Gqgg+7
RM43+oND44Jk98xoohtf+2jHcoxmcXVnQo7/XWSxF8p88JvoHCu97X4JEcaAF1Yl
K+K77NNZaG+PyyAPpkp+EvNWO0ECkBT4Nr8qd9DO2kkHfMi/7Q9fz1VCsdbvQi9p
9mo3wXhlKdpPBANWaCGLPpYVgyqZ/6/USLK3Bbt44hyaIL0crcbY7zDX5feiuj4B
1U1TAnztHZ1f8KfW5W9bok1STxy/mPvDD/T3PB2a8qgVJWtdF/kYnocJw1WRGXJc
uTr6bN7Diclt6IJlX3lqiIBxjRJ2Gm9SYX9gsFJxbI3+RvntfFZYaxdtvROMLsUo
P19F/wsGwe2SvCR0iy00rUHuz4ugEaYEQUuj5hlEYsRpohINNdRxQLJ/+7GPzv+R
4RCOgXZ6uSk4c50QWuI+qNv+TZmAk52lxlDBDw5pcct8d2SAI3x5fxw7R6cmkKQu
idKtjAjPI8vgrQmMU3WfgTkBfi3hLF14yv2lnjPFBsACsojrRJqAsrkAbrlDTPcQ
+KDKEkS6SaorFXb1Lk/wHoErb8uJeRevH71MU0lLMoHCPYtI34wY6bES9tYtPSrL
SNzLJVLgl6hjZfU81YkbYzzwoF3R6uHBkq7yN64FsDgYIE5t3ilDs8Z3n8T7hrt+
VLy+lH8otjr2Y2y+Wse6MtelXpmObCEUJia47PRvxtKoPBMtNHQ4Suki0txQjcsI
3hLtVZUOV4NtNnKkEog1t9MF4lTDPQPTu2pTei4AcdHXw73DM7XJrDX+dpwmL/4g
2x7xhk4TTN5J/x9sPYqn4UN0gFFZWRwKY92+NfX2YKBKCmbnJ3b53rUG0OnIuc4K
jpfhAa0ma9jfAVcA5nH9MJ2sy9EIEzDjMX6QQ2fmz1xYGu3qJJPCmXtHKKptHQ9/
MnB/sRZL1yMbTUccgs1qjSCnwIDKSecwnFkJTw1rBPg2Qgujhj4QxmdwW4prTv7c
kpIhpg/K6sWFzS/URGWFWGPir+H3SsXqZNTbt67mDYKcL60ZoKwsK+edzZkCRvUS
fplfAYcA6ND1PaUCN6duNX2cQ5TqicVHOyhphUukFVOxNdb/4sWVmJG2k0BCKcAK
q18peBTmKBDULD9m/tXpzmQyhI/IcxFSzvafehn8lmAHARKDPP4DcqKqEx1HENMR
EMBRCQ1mZ0B4RNJIJOfowxvn3N+ezs5gUGo2C/iUJhsHwMQ4oPNV63oF9GmXB9C5
qls0y0Ugv7Eo0WfloYJCCtoDxrpYTYp7Gsr7nuL76JnDInJk0RP8cKCdg7k4BfSO
Tr29eEoVuqinw9/XLH3ZLeo8CC2MOn18Si2mfDkBwU1DCZj0C1fCnK5GV9bIroay
FbxogEWzJXnejLsLJnrkpw/3kcREK6vkyn6zftzNgBCHpFWoBfFRPOuosVZd49A7
Pzgmxy6LTrHLRX/sCAk1zz7KefTgzAvQTEncf3c2hOHGds3f5xum+dWVptUjkMx/
VEHPZIzYJYmBbylKrCwWzxqTAkLFmw/TiU27MsaYKG65avuC4vzAS7vXHCD8KjrL
nGhPC2JVbbPAdh/j9rkcuPizyQpyTV5kODHEEEL7oKrogy4IzZQR0miSOENweBUm
TAtq6woPaMRO8nfTtl80eBbAQ8vSXGqIkK6P/al4ghH4yVrCQV3BLL788tsflXUR
D1Q4TdcuGKatb6xaccP4oc83f+E0ndJkqCyOZhX2JyEAwYSSrguH3tB2kK7PAOFG
enQXrjGmjTQDqgJdjX671NuSDH1mC2iLSAxaczJRZIG/w+Joe0DfnvOiTrWVIqzT
RABBjq07VpAGW43BzLi+GExWG5od0a2V7mjo/uIOFNZ5LxAXCYNQOjJMu2S4VBQd
rpsaKCmUym19sXpzgfgiy5Qi4nLXKw/3EHUT0O9fNHaeH2//1JQQh3X+jJve011B
I+gSAaCADJ7RD41B4sp61jesXLmYIsCKkrWapQhalVT3LyOUsGvSb5vszxXbnoCU
QBRf2dkuV1WS8KAdOfscQiYSu3MEhJZ9InKu7YID3F2SYGaeJBMtU0sDhWdCbwQU
5diiDalCjnxtcNp7B/122aqi9/M+vgZmNnqLR21FRmQi/Qrfh41dxJgltWI+ke/p
eD5SCJ3NkMDTAN6GFVib5uQORSLrwSO8Cimd/Jvj7JojzCEYP1gYlRX95VKO0Uvs
GPWjtomLiONpkG9/z5bhzkj8f3Z2vsi/rSH8VPOVzdKDi2HrrvZYyOeXWmCIgN0u
La8cSOfmZPKlqavlGYWZWSmvgvmQuZs8Nor0UCPMBDX33JdA96BdF+DxThKgIa38
Xq2PcoPAZ/LyuBATHp/Xp/YTQ0IdRN4Aqrgh3gtyDB/caqNy/e2qpvsqsZSf8EkW
x4Tkm4T9tY9wCqV03KzdybSkxxUiMAtZmDLHGDCmn54iPMRHdfJ3WHXfR//Wx6/F
4eIiDDQ2ahVLDK7wxqnC6nJy5d1FH6hlARk5tmuPai9CT/5Ng+aDvxCTtITKPVnJ
fYGosWEdjt1slPB+jBdAbTQHuTdkVnQBFEuyByw6ITM7EcY1WY5g476+xx68fB5n
63d6e+dtsqcbtfU7Ny0ev5b7+IDDwJlIEq/wx04aUfFqvmxshANu/AqgJ9N15M6D
pO9r/lVe7wGTcqkEWccf2l3I+Gsj6Fw8dtOESGLH70UnegNhRst6Ji2eaIA+pQQb
Szs5RBJSYEvviTWhvcik8lV4vTnFxWWE9AFDMuWm21Bd3VAMNZUqzks/r3BlcOg9
+RsDbw4hXaB5eGS1w+aajFtiH7AjRCAn6/ziqKU6VVlyKucZdsyjxmuUrsUBGWUZ
xWkrmLDH2NDHJLAndI9cvXKcXxTfay1q9GjKoDD1oXvNjxvmj/mOcUElHQLFHItP
fHyPOxcOAXpMKSZveMHdZHxkkbUP/HW8WH4UtepadfUUwyG3mBMfMaSzRWIfTwA0
5yL4DRuPkkEzgkC92wsamtqIX9OoQ2fk7N2u8W84d/hwypM9TUfbFBYgXwNlm0tY
MRtB3zcuckQLVadSCeGU6hMYVfIdj3GPhSUQv1k2cYdQ7YjbP2d+iA1904FmB491
3j1ZS40bQu1TpsH/RTkYHOCmm9B9NfwoZKcheLiCR16hy3aQo9WH9o+4ynDAR1rk
yJDbdfyjBdxNPNybgAbyaLTnBkRNj9GobGYukw8Rk+5sz89koATInKeduexN1n6+
rxHbCM+1O0jGgY/mr4ZFwlE3N8XrNNXGmG/xeM0HhvAX/WV0ZKWlBu0MypjaO+OJ
EBCSNHotCGNH2Judt0gxDmZsj/35PteSZsRhzWVk5d4hRlqYiapSTPTyCyKnTmQK
rcsLhONwgKOQfeiDvAkLk5CjmqEDkEduwqz6bx4lxxb3VENVMJJ6VY2F4cog/4lI
TpnLZPds8piBVR67JqnchEmTrkZYdhkewU2fkeUxsk+qfVLjZ9epKSyztyS/VBA7
aCRhCjMHicOQldsuDBBwYXWMKP6m4b8Ore+1YYnZ5ahG84zFh3zZisll+5ZuqyID
kJRDaQ5YpxBjxRdUV9NE5u6pumKYcqTODuw92jV8L7R7qPXJKltUmtUK2SFKyRPB
8GDCA2/MwnxdYsZwUM3rIPmKOzr2KZbY3so4ki6m4zg/INfkhZcjWqutpEWxJQMh
aMG6MLWRlSLIzhWmES5+KrCGln6jeRy1ojCtnERX7NMSw65ZHWq34aqyuCUMCuiy
Zsas6NYMzPLMgoClEy03hMUFXlZnhZSBu93fUj4N07Am3xYMjyPcRVeMWWrZ1N/x
rW8xIjB5I0ydbBuA6/lP2s09xxeWHXiQnZvT3W/fC8rmadTVNyfiWjagr22ms4uK
rneNNl+JAkX515xNKFYypxYiU/BsPB1XBBKaeOZvDmMC5gz59qdVkWDn5tlq/C+y
0L/zq7wqZvBslP90Egbd4zb8dLThNLSWZlTj3FvlQtXmoGS5sCUbBoDbuvFh8Txt
C4qGNF2hJBgNy4BGXAHg7q0oXC99m4sbZV+gbIDNKJC8vGG7ybjD0GDdBMNXBFUL
eDyZR0C6ALgCvHclwzzF92gspJOeSQ/TcbbSiRszPatEo9KdI4cdG5i++PEveXGq
y99gJwf7cs3A3wFtAjs2Il/Mi37iN5OWNvhvh1+vbwdrdqA94w2seLvJL4ZbyQXj
ieB1Y7YtK6ihTpVAoKSRVlPlTW+sNcZfd8nvhqQlcXvott1YhvJ5F3iEYwJQgjcd
7B45WI2f/Xp6+OA7SDuGxVskvkPxjOX4H0zEvas0ERpiPQnprAf7QgODRD9rmp2m
A19/D9iYfGJyZ2NC9P9NsrGeNAp+yCycV8iwJpA8TWkFs0EoTsiaqWw9YvQTYoY2
ZlAtYEyDvMyWpc6pgJPk/c2yPvbYN4myMpow3gCuLBtSAgmnVDuYD0F/IXi2sznk
F5ioXgaaR9qRwjYOL9D1UhEkUbQUZxLsPK7RoYMcUctZd6dCX00aH2ghq/dBb9zM
FYuMhVmifJMP7Paj5cqm7BIt+yeNbQP+qMAFGKah9GUjLGF1FFRq+6O0NqYpgA0h
beMB8gCnc+e1BhWr6LKhvfcMA4sKvWSSbfQGKnC0v6eG6l9YPDMF3OIQ0hhZUkZW
wOEnJaM6iu5x+C80UQZj4IRT7rXXaBnI5ZlxDPWOZeLHVcSY7ztKu5pHTSRLY0Cs
8awvj6/xfvUMUiH8ceejgimKNlDef+PfkigQSfknPCguCeed2PLea/XRyGTYNJai
/+gDdyJqhHnagjdoxXCh8wUmpXAKpnJrbG3WX9DuJOrZzOKM66q1cXNdWzvg3H4y
BnSTlukObWcKW8ALp7weWuVjDvIBXV5JYTpyoxEq0ABZfXtjyP7XHxFc71oqs5rA
fn6cUfC5wuQ81tf7lvnqPSzRh8qVcBt7DOoV00EMDdjImMu05cOtexvZ9g9fjkER
aavphd0kOBO6y7jhM9hRcSG0vKjW/faqMHERJvNv69ACeqh5QhXo3P7wgvABlyp5
qqkMdLL1ZtHtpaJquOwp8vg+VL+8RzxdfweS9iUrfTBMffzjUx5SuAQn6YtfnJtM
eDrPM51CKHT7b3JEGDIVliUWGe7OR/YOb5tC1CDTVebxhv9VE1yegBbJvvbvDl5g
QzWb2rvIlvXMJy8/FtGQ1fd2DBHYpzuMGN6DWXK90nw6fDqZDf8zYDlTb4yuKCE8
D0iOTTHafsfS4eXjd/dJX6ak+gRxxrQs71zyKWfRXy+9ol714tGsJ2MbkjG8Zvrw
7sX3d+vFetCCP24xT1hSpDZrwNGk8rl7lOZeArLrLiyttXnuIRs2XPta6Aj0UL+P
KoxDI3p57xQVP+hnYRSvx7DQXrdSmFoErUPwh3hnuZO+EzDWlr8lpiYSbELXuPhm
rIoTaEMMBraO4HiAwKMpsM2F9rbc+BfUdsbw50f5l4OGfPA9ZS8BgCGVDWdxqjnR
ZcrrTy7Sjv2w8eqc1QqPPlyrhXPqwqdbxoB10qT/2kgv+EjHqm973SZuNlnKGTFj
Gq7HwZterebAOqR2LrBVxXgm+r1ctbXSikym+SpiuC3pJ93KK95/rWJHBvxpu+mW
W5Lew5oizgvUrw7DIS2TBhnJUXJgMKZCHnd0do5VuaRi/rUmcf88qnKvAHm16lU1
hpoHliLnNdiUIaQHVEW1slFgaiu0p9VXVkErcsNUUumves0B6zxiMTE5UjLgAvAS
qwaUWnNW+QxYa6BZgL1iUijNvMxhjhog5Zci8EMW82HJPUyLwjl8EkK3WtPz/YzQ
sfldxTEdrIblss98No4Je+0gx/C/Is1N4kpiowWTcJQ8lpuEAWQimwrMQKt6l9sP
0/HDBcyi2RSUIDKWg19mnSba4ejrSVPD+bM3AOyi80xHep513ZJGaNlcieNQTG8+
ZNYVXFdy7OlU7Kf1MaYJE+0caf/KRMIYdqwSxVfAExAxwHAmHw0gZqToUSZIutQh
Mf/85nAVYbkuicS+bUFaYZ9f2dFGoP5JZ+G6driHJSUfFBICJBnYJSwzwP18Quku
/xCBv6oS0rp/KriflObkL+ePwLKJa/J0DRlpfbukCk3V9oASyCT7H6uesNhrfsEF
g6pnDr3lkh/ti1oXP3Cb8LfhbFplI+tYmgG+Cg/XgmfaOUB+dvzHezwNB1I+phXi
g6mkymzBdmFAQEFGRiv5Cn0wxG9++ZHUjAli+i/oyZ7ICPwzgqT7bFsjtEiEOSc4
1rr4pA+azp2yjU7MvEfOZ+GosX6OcpkOCCPDqfBgv6efg5pFZyy8D5a90HGtnmYh
Jd7gYg+4CWH9Td107BrTIRQV8zaHX0d4qFVFhpZFEDAESV/xFUL2F0QttQjwmyti
uY8FSIduwnEXOOqStVPKJ735CzqDx8LgSOXETMg0ejVBTVvDej/tmWjN4hERT+XT
zBCswbA2vf0hGEIt2ltNJ51npOAM1uBW05gKLcyh6PDi/cpXKovzCt+2rTnRYjeI
wfn/gCf5/87BDCF0YEkv9U2rnUQ02Wlhzj+8qFpFSafqgsrKQNrDzGd71GmZS6d1
EnzVVg/cu/8S6IF9SOCpBHJINhF8sXd2kaGKdTuumNDZCozYeh7IULC4dDu19oN1
X4a6/MG1O2EZ0grUikrnCOPAp2+ypVhCiK30HgJadtOE8/pXGQHUxg6ry/pJ9WRz
tYMZYIvO5Eipyhgx1+o/cG5qi1OqcfTXcz9PxbWL/FrjxlF23t5G/V9rrH/OIE/x
wWTirSJ3u8UDuGm4FGGEnOXrbiBBZNTnJtxL3AhfMOyTUg/Yag//ZFdouEufzdRk
/sW50SOdAxJ0DoaVdZ56ffkXwgBSxaHHUnGq8bhy+awgSwfAYAOh7dC2NVEobhQ9
sAMFhIOLpQeewvunUBPa4D8b207ZhZpluFgz3l9g31gCHQXOOymk8Jl+eWd0I9ny
be1xxUiFZ0PApN6vqCXmO61lMFVFeDDFOAZ8Lfn+8RBm0uI60Y/t6o3NWfmDUhbO
FZUT7Afo8NGaYSJoabH727gh2OYn1glbNW/f10CioBa2j/atjWDIzKk+9vrWo1W0
r8GNXkeJHt5VhsFgP2X/j1jvxHBTlrDhn/D0zmQ7tYdILZR/dLBkxuZfk2g3WcVe
tSNnF1bm7OKKa86x3frJgEcbnrtxpund9t/PkSxYi/bOEzG6WeZM6JeLvLip7hTj
ryxTDfctlfN7642mPU0ep1tT7trfoq+3qj3BcwfL/wyb9Z2ibnpwgIRDMQl1vXdy
uqNI5FQOUz3Ue4C2a3DqafRyH4cYfq7zvg+vaTIYkW5s3NzghemKGC7z5Vu5WrlO
X1ZVmzRUiP2hb49kNNRshAtQgfQSXXtjmN61BNlmpnmpECvTXzs1q3lXAvvQuJCr
AQCkSd7GcPap/lLgPfQQvDer5XLq//IAtzfnhIEjkEsMfNDSgP37DiWvUS4qPie4
oKNH11E8EtzJgeW1UMqdlokquKbzwn2MaUoivQvrDEIESwuJcrRZYbJRAb3ZkVMi
R/G4pZDL36AXRTKbUKZBvA2uSzlhtAKpWqA6Oi3XSDmkU1QqLkjR1xlL9VF/E6h+
UajEuH0ZhHPBI3L5uuzED6voZk/ZPa00WuU48h/tD+BjimiR05OlhGb2WTShb1sk
z9qsEuxne/dpDGeuuw9aTikwLXfs72anQGKfQBjpbSjjTEwSWctAPggWRUo2D6iY
26NsWa/NP/YTgUDwc9PmDhJ2uOldrMEQB1TKLq0HSzkRp1tzx6aPTDqdYu4usgMk
eJLuE+Me5V7dkPDCJvK6KhZ9tIq/lfmmOR8KRFrKovHNZ2WEh+w76zwnAt2EFrFS
CQ/PHiGyPi1RrogK+Njsuj2zjnoMys1NWnXivTKG5lbzODK1pbnTsU1PW4Pusmk4
aaLh0SZyASBq39hbyNnCm3oouRgxgOm0IxyUgVpqMFGDyKVvhVW04GMO1BRnEQLs
bv95zC39dlP5CNxnJtS3Rh1Vsn+nqtP+UAYILsc0bZWyJDziHVF1r/ZWpix0UFLV
Bj9TAmpdraYq5i7GwcaPHuXY89dIsfltxObHZSAdejpi0h4QY95XOu/Fvs79TqYT
ZtnzDrE7siOILyckkCLtD9AHb88H8JnaqeEBgsNUK9dB2tYnQYYFg4GdNcqcMh+T
dwfa11QSWtkAnPfA9hJ0w1/04Ma4V7dYCmZkLCEm82ddxD/ABIqn1iNxmakTpeJp
gBqNu0QtP2C2dD8c6FD2BOiVDPgoQYCwJZpKzO6CSoDYnoZjIQRMWswOliQfb1PS
KakGTqgQIDoxdnGlT5IADqC5ggnBMTCppkne7NM/tj3NtCnJTYSobrkvJM7AtPoL
R9GcqRJq4L+MkQVO9fiffobE4nsffACigzXZYP9ArqxhsMHqraE3j6nJ+sv62pQs
EW9bykBgvUYAs2B/cScpEHzFY76fmsZcTBGxmOvKZ2FDnByj868qxEU1JiG3D4Wm
D5XrSfRo3tk4tL2OSa7TWmfdenFz4iAtQDcGJlv/cCTL5TI9mwLHUko7WDrk+IdI
tMsj2onCfpKEBcg0XFvUAVA1DUayUP//3g9WjnmPidbilhFzvalRLnpWXK1MymoJ
FxV9fy4U294bCss9ZEQCAuzRkRgk3Loyj8rIOeZ26eTPOq8qGuZOMWhxINpyKqSg
jA3HSCOhuWnWX/Enk2ComdlfMVIS+7rHodMne8HnEiyUj/ctcN7z0aazfi/RQsOe
RPM1Lo77R/8ETeFKW+nOG00luWnJXZc4NRqUt61DRjydLWIRwvo73EAwy5ry48hS
ttifKaks43Shb6aPN3ANxN67azET2RlAvGfG4cIyM02tAbXzJoCtvgnxB7/GWfVY
fbStEe9hQCqgg/X4FVa9M2lYmfmOVQmY9HogvYTJ7sRSrn3l8VBMj+f+FnHHQGs+
VILK+TVm5io8EzJihpf/JU39K2IP1kCTcvX93g6wDuh9fBSk9aGAGLkCZEMjxSY2
tNXB9bcQGi13dO4uhxo+0DT4iL6JLgtI7a3x1Xn5CZRHjf20TI2E53ZxXOWOO+Hq
umEuZAHyt5JOgkpF4zfPnJ6e0+I082U1W53T9DZ6t+l+bo5Yannf1SUM91xRfQWs
V6axMB2lwfztqGuPLhNGHv9Pgib9Rq45SzhajXp6l1vLKi9ndMPQX7SvV6CTS14+
kOnX94GSzRpsRGS6clIxoa094Rlqo48KDPWnXaKHM8h3S9qVnyJB5pT+xDw0PA2t
1aqLpIaQ5n2OjWCuPlCIiNBCABiy8Uwr4bxVrdvCNdB64g5XQzW5NI+rZ62uTEWr
2zDO6sTmXB+Ct4iGsmoYhpDUdhth7/Y5Ui5O4Fu+VkKPX6vcn5CxPzlz9JWQM+gG
1DokUY73tlFLs2dwaQVPDJYoEFp28MT2ATEjKRg+JlTge3U8ELSKue9FUBVQ5tim
JLJVya6JxsT7WfeoPhZDlPocSYYmc979gmfbP82RGn/+//DkF/JCqPw3l85vBkdj
JDkYfPBXpJeXn3rEO+SOtsTcFeiYOTAFVFAXzcoqFhYoqIPYiW+F/3OaV6l4boQ7
X9SgRL++W0ayAY7o4QgaT1oHSYfJj3w7/Sbuu5XGX3Yk6QZsnIlOlu1xKbND25EM
XVUrSVGaKNVRa7TpJtQCJ6+fx3cuhwEKY7vWAvt94W/ud3uUZTwmxkXsmDmjuQD8
/iaQZIoymtYbB7Hd2nOnYPHhsaZsUnYAKFq1qXnstvtgJ/6vT5neptIhme5DgRKE
JYWUn+2up7GQGoIiW/oFFXLUm8QY3saDf8oexpq/LtBoRZhCQHsK7uPNF4xdayP8
mZzzu2n7RVpdoTIveQaXzb/wTBsD68xeDgd2N48tEM7FQj9AAxxfNEFfB7qOQ8GP
1dGcSVlE2eLrQejTmHVocmeZG8e77TL3y4tnxRtM35EAoMbdRVoPiU0jWx/FomhL
Oz7VpkSrnEFEg0EpNTA1CS7zwodnDQj7hujhLYAL2hfkM4n0XKpZIYYSajRE6GNg
ABTDXwenPu4lzb+TXocEa+OQSfj1MlX/VPWe6PtN0jTThK6japIH/YvFRlqWBK+1
z7CkKnH8VYcdiAFyFpEeviJf0r9YiUIDi23XX3kAus3pPPfx0IhcnasmSSjXWcQo
gPEAhXDD4PBG80Oi4yn55q9wmn9VIiouqY9brtw6LPxal06f6bNZpPwmQaMLm5tv
cvIHzTjxLSGAxEINO5OkiEazu8E9V1a8V+9UWGnKA440Mopum2123QPIzrUMdmXA
EXgjUhVvwJkJmtmHb8bt5xeZgZREONVx6SxsaNu2kWNq7UfV1JhW0bnimSxOHx34
YKzTpE1t/ITA5tNwO1nJxSs3GrvVxlwIg0fKuDJGha0CNfgib/cT/J/Z1XZd3o5l
l6/as3slE5qd/31l2CEOF5NVoHPi7N94qK5zll5qlzrUhyub8RoHU4b9fhJyPnUq
zNGPZYgG8b7FEXOkohM54zC656pyDmh96nDvRQiGXJCzjQIgdOmx6SWwOjDXKbwU
+mS9ue/n9znJnlnoL2QW2DfABsSJ5VKOj89Vx9zzTjfB6U3tkFrRQueXVkbgXck5
DE9g7ftVgnh7KwNa/lGKeuxvG87qpRiMs03t/RYU6grJRj7ZLVWbGyPhv0f/YlhZ
XG4zgPYkWy9pG0S/biQ2D6Qsyep2LefkOoYEYrofw2YNqLJZFNDrifJrn7Wbx8i3
bdKU7V03g/wDK8jQ6/I3rMnDr9P0ylktFwqqVhpFaQ7jY9OS/jQRxvxUiRWAHlch
I4U/CgQuu3xxG49/8hoPjSgxWAJ7J3yao5MWim+FzS71Bs8atASDSg4BW1IcO3fc
I4+97O1qxNAtf8BnORaM7+UeVeWrwANd8DBGxErNPvLH+X2LcqgH7XViuKNPhECe
BWh+ysgZnCGmzQA6HYRR0p+y34w4w4R0r27D0YGSxigbOeZEtxRCxd3v7xkhw8Tj
aL4l/2cNbnVP60igP05gVaxamtLgsLqjCCW3fQSw0xd6etsZBMpq6kwpZzyLoQTk
+2VJeQGsJJnPrLszD7xjgcrcZRZtydZ0bSM+FogC9mjc1G1RBAQHWgg19seF4H/0
G8lRm8IcS17yqklWU6YqG/QGKXEbZZArCne8XDaov8LN6kPAna7tn8jYrjAHYNz/
esnVzkFDFptWIUpS8Nw1TdX8TRAbACK8bEPu+t6J/9vuSCcYHUoTrla++BMzNKSi
VhW6321e+ycVWdVUXCiSI6mOyT4jH7N8NAPH1RhP8CClnzggrd4Q2rrQrd/dIWCB
XWa5T5WXXtayoHL3IrnOI8xWwA/BJ4dYgnGlvMNH1A+PB56SgEabSSv+qiRWmlSN
jl7Q+/j+r3tWcnMJAfQ56nzf8my4ikRezmb7G48Lq6AO2c/iHcc4N3CoP8COZpn+
sMHTC0s3dKwE2W924eEA8O4ogaoN167/hxUK9qBiUHEmLJkYW/4vnh3ZlSO7bpUB
I6esCtwxVtCPxRpb9k4YRWBAroNdWoFRRqAuzIAhTa3/On5012O58IYuJo6wSQWv
8C344RKhGUdeYyo/Aj7xzVxEAl9RcYylzZoHQ/7UDawFv/SVgLmqRBI3up+F1dY7
CyCduUjZ4MvTB9TEsbYiXpCrD1FvmEZCcf8yZhKDNh/HmQItC/HdfMO8Y+2emUNm
wDkkGCLIulpt5NClWSbIWFGgdVTfaBAQtAFynCvqdYgplxbbiyGUChYYUkLZDub6
uERjVWXVukI02MHwdIr0CqzAKH/7B1FiRQdFQ+Zgtgdf5NipzQMOC0XsAls+cgor
IS3ceVPy6HuQc2+EqwWUKOP95x5v2OEzU0ovygpu8Vs8v8JCx8R8zPap61RNyjwy
thxsBoAv9xv1fFSQUsAg5BSA8f9D8zmu0JU0qTCK8nsJIfvDSklYOJZJ99+JOcE7
1+qnZmU1W1OcjJoTHNDE7sFUqP053HQf+pH4BUJaHkIXEs3BoOVDlGInBrSLPuJo
4UFk+u6lUYvjllhi8EY1UaQy5+vgWRjWgwRaNu11ZXRf4AaRiDvsG/Xo36DfzBIw
BORnkCRr5OsHpG6i0s5LWNYvZLoQzb/Sv4+gdmsjwBWOfrOOUodsFQTlZANB+lWU
UxAiV9Rf6aF5d3z/rWcB0x4u+hS641nHgME4TK8TcMZkAt/56AjuhYCktwmhrzbA
1yPqazRp1jhgaZsIgamA+M3LjSAED4i7Cv1HY3nL5q/MGB4NA6E99D07uExR7PxR
qhTsoXSTGfyzlshgA5R46ClZTbGKm8bqG+qCoKfiMd36iRIYE9DFZJrGWEAGSbVP
R6m7N6vyTUW3hXkl7YMuPEs+1x7fNyEBxUSfTUDHVtU/J68gy/Ks4ghPPcoSCqbO
ztY0hYhPwMQ/aiGiZxPab/53G+wzhse/4ayyhUp8WRAeQV6EkMgkzejIOdGY7VIN
DZYFEf/oPtFSSjEQQV3MX26KqSlXO+5naB8174yPrlP3iDImbbIda30DtgsPw0rv
zC9N1kGC/ya4ARK6pKQbiai3OlxXAwuFzrwwNi5y6pyIAPjoK3gu7m03pAVsM4Yx
xzbBvdKl4NcBzSUJufPvhhqFuU9lkaS0aHmAfnT5ghnKMh2KizBbulafe+m+tDFS
Bi1Emxi2sywDiEqI2O6uMTCAjlnP9lOO+spruodyrsGtfOZIrZNIqDq5fAOBYblu
YFYPWFyeqOBiHUMAcFxHXMxl34A+vKt/7X9dzhyVsxXQfZGH0Ezy/lfNCeB0Xvyl
1LxlvCWR4E148OX/j0PKtcI+RD7rEknwz2i5iq9oMyuLeAC0tU72kgF4M/h3iZH/
N8IOxG90fwUsy6Wg94hmbS98wL/UHX0chTj3MhiV2gvrC3ZCzNyr+fo8/ZJznEW5
HVc6sShfZAx4joO2a5RzY+GbrXnQ0xFNpjXYlhTlnEBO3q7zKGJTvOynkESxJyk2
U2c0IUjLeJBI15VTX7tfp1il4kMM9RO9fmRhAS3KBGsByWu3J9UJqK8U5V2eo3Fu
oqi8No5oms9rV+fIokt7wJ/H1aD+ThTF+LcEUTNKSeV+0aZUZBb5TBmlF82ot2Hk
QmK4Kqn6Ek0mNB5cqXNls3TUl9W5+QnwL/KKooOv8XGw9fagHdgBOuMr/y8Vt99o
ujbF1h0BChLoefdNZnY4DZt4eIkl2dhhMxTl31D6CaWt+87ZFkK5JGzxD5Ckhpr4
mxIk7Yv+KNmtt0ZYF/JGTfENlrk3Y8NB27iztOq3202GwDaW2U3s6XI6JbsdULgp
fcVMlPayI/8SDcXDbekUzNGe8aYNdIRFTGVmeNqiAWc2ncU9mGZkA7gMOQNKyqXq
dSvhSbUbOtpRn9zZMQWtiEPF5o9y2MxghO0blBjms+hp8THZhrHs6SjAbGBtA01g
hvdeRmnGFDYWj3g5J0olFS51CU3K5jH+PBWKoBiFMHBYf20UIKNxjGOMWjE2/Quo
qK8zfLcT92ULRePJfGV9aXbJ+tbJUXlb3jFGvNZgQC0smnVYR4i1t3DLiw/mxfJ9
bYYV+zLhh68Tn9MCG4/9KalYHD9zXgU2OWJ71qE4gJyIsTmlPQejq8dQC+DfMPD8
f2rYLBHjHHd0Gd6RCRTdT7nWsllGLlz07ddnJ63CiJPE92M1Ae3re0cz7MAUFhzV
MdwFbR9Wge/YKxgVsLhLuSmpAY4H1LxtcopdmwS6ITUk5WIN/T11OAkG8m+oVsw9
wIX8ua816HCwJGxFzpzw2r04gtuXyYt2r0PPtFfegHoysq3smcVYuj7oUi+EIFQk
2fs3Od6rMnLKzpgEk04DPJNT6gyprTe56iFPjWvaEx+woD2Jw6DUWto8zsKgGPyb
CjJFl3WBrj2xKYPhlryJCtDg/GBkPF32D+Y612sCaIT7BXT0oWvzW/J9siCVQhtC
eTm8PNiIE2czE/rc2+83ELugaAqHe88eh7T4URXANU4MjzgczWUwJRVJRuYqRx3t
qNtR6050YQ5S3JDsPi1DrYKttPT8r5HJj3K5gfiXbOrw1kpsmW4HB84cIkPkq53s
e6lW4sx35y0rptMJxAVVrrB4XN8Xpf/j4F4rn7FL8ktfqXKvdonXJa/WRBivLcOG
81xQu8MvOzq63m2vd8DF/m7heCWELGGjv2ablj/1f38SHdJndT/fPExuiv/G54Jn
JVu9Saamf+tU4cEgajzXH4uZvLhqtfZpr0rx0PD3rorxuFH9FJdRxB86uEnybgPW
V6U0VBaGyBzdAQnwaks8DhjqdKXSyuOxD1XntSZi7QvMsZlTSljMYEh+KSNsUiZX
mUn89xY7Pii3j1z3rIf6JR6TqDzQx9+WAqDC8c6C2FFMYBwtjjS9Her1zAL1BiMF
nAS8JJcST+DbHwFFfUNbwAtx1GUyf6zkv7cuTF64tujDyRIPlMN6ywFo5To4HNa9
nw8kFFdN+IixDUllphUDj6rBOawN7i7n4jMt9vJH4jVQ+OiakrUHtOmtn8mWoGhG
Jfps7+L7GwUCCf5/x1g5Ck8vnfdmBLp/PG9i20LB3IAv2ma4SUqPP5hz+1//d9xB
w8sevqBpr88YPOFKuQg6evgnHEvgVEDAvLZitcpLCFIfctKauV1GPWF5OEtLA1iW
VGvZDrqjCud92ePIV4/dB2zlcRtqYR3T6EI16A09YGWrkjsO4+cgxojj+V05V2L/
yyoABjutPo7o6TA5gfmmaoXS70HY2ZnHh9iArZjcGNtOWnmuCoqJRlG6IcbylVdm
wiQS4lvzd4IsZ/U4ZolXvrc/guq9S6F9KrI+azVrgLT01EZKUs6AgfHZbE4O6A6R
kepwuGjUcpvyblgTdHYZqDdhQaAI5XtJyNhEWQDU1Rqh1ZI8P7w5wVjDyuzfvcqn
561kDmX537WomgbzADWbBjOih70EeK29+V/BMOuHZAC56uWXsJsjcvbFufIvVUA+
UxS8qofPip+aHWbUp4idKSJisFhYyW5o4tT2anRgcRgt+Oji06/cNgZsPDWU3u+W
S1Q3W69OM54E3YQ7UY9FjzN16MNNtW7BNzkOvpZrNNKGsMCinDxM4b2NyR2vyZNR
QFme4M6WFm0XqFEq6yYoH8Y6/XJevEOJg6I2haYYasCqVN/Qzd1eFUBa1BiAcOz/
JniPgUApyHVESlEp2ac2Uyg/Wlff4DTMeWltO8h7zY3ADGADE4bQ/qlom50SGs3H
+BHritHE5nwxRP8EcDU3QUt4FRR1Kl8twf5EGLDyUTWkBYDZoE7tPYtYeLyxOR+U
g5LUT+mUl+ZkJgf5Z5m9e7D6nGXoEHIH495eH3Yl2pQgWy2TCgSugMLOQbvVXoYi
qVYI3sjZ/cA5LrXrO3YLoph+hSJknxF3C5rnPxV7jl7z5Ho8Zt0te2voAzApRfQV
B1ph+XFWIxg6PmrjUn3K12Q6mEpWizajiszWy+VM79ElrQG4vjVumiTHO6OORN7H
BE25p901jLqGtIQH4EW+u7M5tvKPMinCfUlYJGB4RoN/o4Y+lQSMqOXm84T9fH/t
S6ltprrVxyUGJ6pk44AzD0gbn3/SQl/Vs3ZCzqU2515ZCwf8yYTRdEPD2QwQHo81
NSJMS4oRPqHWA0ylfsbDA2L9rLBgehVQ/vaqIs1A9S+lijRJryGlgRcWRiECgmEv
VMx78U/O6GmsLTZamYI35qsKVCeaKOsh1EnKgWF49liwYGuuOHj89GUbR5+SGzTy
BTEq59pB+jjobHpC724Bn429OkM/OfYRHOsbRLR8sxbVAopcoklWHD1ENy/5glvN
Bzc9iU5vYCiKa4kArcmO5IgHj3/tkb1MAVfG53sBeZTpF1cm/yDakyo461ZgR6fq
0IpduNCeci+bdY8/7+W2k5luYRlFHOUpQhcFhdcr6+Rtilg4NCNZmUHPnETOyHAU
U6ZyUw1hg+hDM7ZdXY4PFbetpUeI2s0EarFT/QY+Ax6xbWkdww0KXofMudxWlBg0
VXb9zxQSfhtmKSgLeLRim9uNGZeS7Tr9QrUh/TPt127NfIFTDjm0Yoqm+7PXTpw+
4U6LYlEb1vgA7KjVmc7FrvnHlHl+StHaZwDUTcWTFwacbELBHPxyjXwRhJc3tln1
yCGYGeThMPH567mWR/1tzRQTTsEfksBVkrIxP4UXvIODf3B0zSzZUqTzTq1sm5he
FHMbki0ajgA5UfISZjtdZSOype6Wn8vavHFU3fGSmvvz3JNUJZYb1/4CIZdBh41B
K8le1xmNAQRsMUa4kKGaiGFt7W0HxjMgSIXajzZACCTvaH49eMx2w40Ura/N5Wyz
hTqit0nqw8d9tjFawt2xV4ct06xSfPLc8UtSqkE/o0GeKIsoVqhduDHZpisf3D5R
0JE99l/8nesWSkk4DUo4rdJ4niF0I5zE91+8mQ4Fgra+ZRjLu3BZZLalU5MTeghJ
RNwxBtufKCQ++ck0sCSrKj7E41GFw9RjyFZUikm3zO6QpjeNrKVsNI7XEmiagvYs
EsEJjhP9Rq6FV/mQBVWh5J4zS25LcdKGo/o+LtzWd1O2sk5AD7pta50HLvcM9XYn
Hsfg16HfveniChZyrJbDX5LzwS4avuWhH+tDtg/grA2PVHpGs72yEqsAF9eT843s
7OWX9V2DSMpulkwV4km6juxfqkXlx6944/2X4Ir0orX76vGHVzWQ6H9PZynJze1P
+stUiU4QxVP1C3LOmHtsHm1B419MWZKpDPDLJHoE5D6QO254M4hA54SMHvg05gsj
Av/kFwCcexnp+FB8/FLmuy2yb+fyQ5xLEn8eQa4OLyYYTwTQTfjTIKqBGM8/MyD5
Kc1/ylxrn8DawzjLejLREtGFG1PjePpRIQLHSjlqioVx2HnG3diBqWeeSSdDwjl/
2esKSmJgGL7/6VtYgkxmb3fWoubizSZUyXKSdJAUSHyqxk/yhfL21XYDRLclqCFb
jqQA3SQRlTSS+lKQU9TaXyoVgGIb5m9cKDDvpMWq5TChvz+mXsmXtZIPhR3MLjhV
BcrGcBYgZ3UWMyDZvQXFWvDKLua9OvXVrYn5IbUalact3gnm+76keI8n2FMKB4tP
ng8sUugGTF3z7Ec8bxe+G+rTydUNCIt56g0yKLcdxsJ1SF8XbYOu+tx8aGA5KFGo
tB4JVR2xU69y8U1P49v22H8iZmMj/ZNj2SauJTjK3UHEwkN8sV4BN13HKfvPN8PR
/TNxr6iels3/3MuufnEoGtqCzQcv5AiT0uKokJrCYHlJXXwcaRqOIcAIqzNCj0vu
HZn6NZY3+PEIZCx/rJ9kkYwZeZDFS6NGrVojfHmunOXbds7UyxnYTszPZJSXdtn/
dTpS8IbofqG1odHv56uZ7kK5jxZ5ppLQVNMj78DWDOda55ynQoNC8T3D2aS+VLiI
5akkHnMcq7xTbsnB/XgZgaoh+yDeJ3ZLQGh4E6xfA2rCZyOjT4PAAe5gJ55o2B6+
m4rTtn20xRvFzZRF6lJRR45ffmnqf6LCKB+ly0g2pIiUglEy0lN5Iu2Ygyh9kWqZ
ac1nwHDRiu6a7zeiDcFNol3ZKlVFoNcQzS6pBvWDvtBBF73Q+NuogUBL0naG3RzK
P3p4BitWiZCaIkHwh2eKMuvi8upEqd8oEF2+q5cjOt58nY1zBts3X4fagbrAY6Gt
20+seDChVGm6d5pjR+C1Dsfz7SYa6rjAAeVzoJ+jxShaE+KSsp9h09RylSX//pGb
tcTZDFfuE5bx6RaQtonyVkpCmPFwQOXpylIbgrjJ8XXu8cS9YdT5ET0v8XliO06a
nMWkwUBWn9E+mf+SH9vSGzMjaqXgTOVD8LpKoXTNvLLS2qKJ3C0Z+qH84w8VsoyE
k5sEY+A/Qzh1vir/3k9d8BMmNvVCJLije2zyJtDwX8twFqCTthFqo8U4j20h7RlD
q699Kbi+hZ0NvHw68b04pix2D2Mc4fketXaigl/YFv+PizsjUL3PCuufs/QkTmny
y+hG25dIcQXgZOneKWZqMpVMOHrbcvxPfolIY7HP4MKs7K6VBrixPa341IP7yMQs
bsv7xJ57l0EQHi2ErSDCTDMdlE5Uaz2GjXAKHmWaieHjsm5BM6oZEHHsqve7iBYi
Le+/p486esFylX7PUquXhwNuWP1s0IEGpFdFUIcLCA/jzvqrmw0itKDwTWnvpgWf
L1zwli/EgFMjOWYAyf/fv2HznP5XQi1+TEXT58LvNgH4X1+GQxOAGrIVNfhaA8ey
Kcw0cbMTkEbvjLph/krU80vN9t1FLiztac0t9VHHCdAzxP1joOvvZJ8nESF+J72h
gLxEzNH14TSYfacXCUhE1FPUQFtnPdObo0x3sO3mreLwHqZ+SadMohVflm6JtBHj
6YgijjA1PakB0KIAcoD1tOyxmMNs04YrgSzgD/PwB6xC/ZYhCtFE+FqofFQ4mQwj
nACFuCEApfSnI5j+GA7H/N71L8RbUdG4s4Hd2wBQkeNlePEGDjhS0zHRZyw+hrBn
nxE2BrLgH5DNRmzBqNq0pah+iKrpX5nbY4CSVQNNmvlmvWjoh2qlOJaV7BbO4XRi
zoAwOdZUDee25vJccJ5pmxFE2QVUxOmgoFgZLZ68ekp/oLoogvuuxmDPIlpufEZY
AQjiLGjnehWdyvPX+Qgrihkk+c/QSfPlw0ZcYEY2KPhK/nRg4zITMHVZI2km68bB
Hca51cG1Nb3qJQopfiIY+hZT6ziWW1gLmFq6cXTF7fQof4EG+AedkJd1/SUvFJQ+
QgWqdDOZYnP5hJNPtPCVimLO1gv+xyIHWi9gVtStvgm2E9ppVeuuOqUeCJgmj9nw
XPczddqAsApX+2EAede90huVcYbG6oPczKIVxnpwXy2RllQEiHZUvNw32i5jwLCU
OscuVdF76yGB4+vZgmMCgs6AcAMnbuDR+qXsdWaZ8GgCNdLQQjw/OfXcD2M656p2
e9IDu3e8oO5k31vPzCMosi1zKNS2NRBpn7gkeZRtvVQq6MHIN3QFF2o5e6yzWFOr
al7S1BwWgStWLXxVfm1Yg434LOlFqfcEOtVG1zTfNr1rlEMNHq6E2uL5a4XdWqsr
nHvJwchOPh4HrB1/ecPLUXtNYFnKEMETi1RxPO4c9WTx+Co74REIGMsxAh0Mnp4Q
tjInk9ylAnTjOletfdrlZNnUDTLVBrxziIjsmP57gnjqPiFR09rPh0+1jbpDth/A
XkS8SJ8AFc/GjwBVF6X/9naa1JI8Daz4wKbx15EBArQyj9N7sjf+gEoSaPfDl/w+
1Pk4G2rujnqjxXTE1jsNKv9atd8OgJEDOTFf4ynFXoPG7PlBU8PNs9QhEY6WQKa9
0ctgekUiJX4HXGxb0+6lMHYF9h+YajpYOfBFgHIio7TDjoiCWdTLXLulhmpq5whz
uXkKhcssVQqKube+a642T4uL+yhxK62DDI3ZtWTYqg3DVuEA/B877Ki+qswSr9H5
qI86gL73Xl0/ef9abjfUf0bOuAwdoCdDNXWZGE/7GgDn7YSgEajrnPoctzziQ5Lt
QMKOoWAndq9FKqefjG6SW9TsBEuxBTGzEOaZS6Zpe6CWU6pm0GrltY0g4DGIAuUM
Y5a1W//Yq4/2oXEhZyFzmSOKii2n4ZC22M+PJalsKg38Ly3h9l56SwwBELdNHmr+
uVOJ7N7AuCgjNIDD/1Pc6YGCl7QutvCwB/7UbUfj3vRZIRZ28zKlbint6u9RuTCK
THPUjmVq72S1YUg0/v24km5mWvuPsKp7FLMjpRVq9eBHgjtO2aaH3J/vdlOO8tRV
DgM4QtFQBI+NC7EFAD+GTokjFwY9pzAiBgd1u8Jo60ldyDJGgycSxUybn3xFwKXD
pZ4eNlRwcrfjSWVYMnvKQFcrMVUb1nySqHBsTYuLWordic5juAcY/SahINBe39J6
j7Uh/4gS/nQSmLD1sy6vhhhTbJaIcfJoLNgyfiPzC1zoauM5Jn/kXO+pbbH8JsCC
nIzwVwO7W0y0s8mKnBEOd/OU9YJMHpsAv95eUr5T12FlDuwNxuwHn+febTiYoQsl
yRMknYKeUQ+ozL3b4MiJIaR3+6Gg1TbM9xFb+y/RPtltUWba5LtqYKRH+VqTNojm
F1XK+Qzj8VJWxeD4KQhVxnAE8pqdmLQ42b2zpi7iL0IDXiXNXQHo7GZ4hysuuYqr
6Ya/ningFbHh4hap+T3A79LTw4ekAImJuFOOLuTM24Y0Pfo/yOLpvDRa3NTSM1Nf
N1kPDdv8AME2E3KnKOIS0rC+3dI7JoBCy04MsHfnPBjTHNBxIRiEG4gl1Hvxgy5P
KfkpWalLuxb7+zDtQBvsbw+eh7a+4y8dYzXmymGwk+HXcJguGdvMstqEJswvzjy/
o1+bRYHjEC+qDlzzzVt234crfTjjDJHjNyVntssGZjCtMNtBmWEre/TVy+Q31BwF
bSWCj5ICMX3mojqkg3nlSaxjIholfqXxZt8Yvz0Fap1R99hmyoe5qsGEr7Ij9oJ7
/8TanpJ4F/piJk1Hy64qk60I4xZmqV9+E75UOMlHEjUrJaVjli1+VDwWfGJLFe+w
Pc8F5o34jM4i3Jt9kSJFnaFcw79WJ/SL2DINYJfuIqL5INeFijlea98OTXt73chU
6/OIEmyiBT8T7fNHaP1LWNr9lG+aZPQqC7trrzqxAd/wGz26mLlP+QMXmroa0ge2
kBSpWRaBningoPs9tlR6gQRUOMxF4YC+p/BrZkHJuNnSk5addcL/EfLnxM6U+bw6
rqP9TtwV0veB3eIdS7HV/n2LPLapeOOo5jiMgUrA0x+Bvz/LHXKoxNeolf6mp+gS
KdH4AYqTEiX8I0v2Csw9QlxDmvZovXNt4E5EFyTHrEoLa0B8G7Hk3gd/F1G7dhNV
3LmTWaB8p+9vdHkbTvXIMrbHLgyP1hzFYdywnD0ovm9R/svaEDRQbeIVyETezrI6
EEnafEshTefnMpIyFoJa1N7PGlJreu0/7zGKRMO3TWTWhH5zDeyZbJuOe5T/AdTg
4h5LVxDqllrbqhK3yNEki0Ph95itwxXlhBic2KKlvCP9t4W4D9dVnLfwa3ieXc42
SXnUQhe9i5IspdGEPvGH97Z6E1vipSUsvsrYZNZ1plaZkUIKXus6vcRqV+Lg8ISV
PfS+ER1GN4z4fy08E6gAwwXsPaFrMRDUWFgMtr2psdb84jzz6Nmn+nVf0xBvkWYU
LPKIW25FZABn4sZEvI2Gjm7efwR6tZaetOuUImwrFShGfQub8fZ6ivR7ljoxilGl
GCSV5MsqhFl7QB0QqMqeIZ+zu7PbGmmFiTOEJCaLdMSWnU1783cXuSFKM0PDo/Zl
iXvyw5Zg69jrBOH9KRoKfIy/wQ28L2Gu5XZX7jbI9TnpTlsaxwCyMTuCIpgvUWwr
Qx7SQsL6SJx2uDnU6vdHSdrhYjU8juf2V6tf3/0CJUhzj5UE9gG6A3f3JfsxAHie
A5H+zgRAQf7R+5H+G/ONSipI28CMkxrUiVZG6TSrSoO9CzPBuEWpLAcNy4VpwA/J
Ico3grjp4+MqFdv6sXPgE5Pze+DIG787XL6ma+f0wwmnRxWberhMCI0VTTIMOrod
oXr5IBqOCYwhRRG3n3qDYFcY8cL6XQPCXr8YySMuC1mfvTC6K1lOtKl6jiRZcO+Y
c/PoYtJYBkevreXuF6khVOECz/IZAZAZ+wCk2STakW9Pm7qYCYxs8XTjYok0w/RN
4ePyWhB2Wv8Lj3XUZcWUiEA+MahstifZLUxQpDuyRpysTOx3bXzAsC6fPW9NKDBi
8jyxDf0F74A/w+zvNHppmaMpIvaiERT6qmls6CAKgw3UzBnYpeFp8xhG5tWYep/6
rg4tebaPaTV4Ed+Y2yVjOLKo9QxodoMhj3Me5kwi9ID0H4YEULvzop2l49BC4LpI
mOD/v9dWnwOIwIEHkPBeG0qsFy6t7h1ekHN+GIn13pwrRbIMy3wtTMbDO7Q3DWmg
aXu0vOWVy/CbWqSEeVJT6WgveLG/MTo9xtvAcZvFxDuciR2BMSBxnHjvK704zeHY
t1iTrWDxkgz3bRy0lupOy4KqSgZ5/SdNhZBw4xv9eV2VHE0VuIzWVknlX+nxcauV
X1M2veR4YRlWPpR7T+V+7lT6I5JKoEb0FpJf96Xj/zBgWXDMW4bHIAtC2djpiFHw
202w1Q8b7kq/fpQHGo2RTi8IILhSvlwqBFsIhsL0eHBAAYXFPc4gXRzrPhM/QrHU
VcuW41jeHnsD7JaYoDK6cHU+vfLrRAJgFKTjIr5UGiX/5VtWUAYeYgZfQ5H+09ki
/AUJgjWYSnqtkW8UTx7YPVGiddALKJNRukOBwzDD+uzpslYsCWOYOZklBfICWmHH
9MiuADLrNLctqd71KsTet3+81BAmI0GCR6p2rD7HRxCR65qTc6Pc7bO2fg6fqUR5
sMjywJzocEudbrdGUWtO5Wq3PFLsjnGpKBYRcwT+n//ZvOHpDXVW+QHa+uCh4XUq
u63b6P2h1MLKNNPyWOsGfxlwU5f1/TENbqKlVM9XoldSC1kvZvLdKSbIVmFX8XuD
qcbL4CeRp0AjuXBGkU5Y15GzoLYksiVM/AmPe4wmo4jkP+Q+plVcayAwE2R2utkY
+zn1woJqS/OJjVvlcoXasjFYj8DhwXbhFuOlLD75mQfXzo8xNxAepVwFO217vzqF
2OGypTdz313DxJvb79NDaX3WmpKFtly2JaN530z4ziEPmkginN8m8JAGSD/+cxyf
HQkuaePdsT2DyTxj28F9hqV6dEr0N1j64k8VCOzLnpXMtaFbrF6q90g/pjjmJEqw
OjUfGdI60wrijiN2ovoX7XffSFUw+CQslJtDfYyhonbftyas+PTUGgVniFXlFWLa
HaUa5JaqY6/RdwOmMHlx/EUcza9pvucgyVRPzrIVpytbDKXR/a3nO4QuqNb5GxP8
/hqRJ98/ETclzEaO/qsdNN0YCQws0o6VRUESOjzPahQmDMuHd4hqEPdP25TLba0T
mLgtLTQrg5fy/QeSUnG5sxEhan+4NLQpwpbAHVeTZl00nUryKPiPA0DiWlvW3+S5
+4ZVYB8eeyPJ8m4hBkN+PC7AuoNCgNTYVCMlUraaQIjGLHwBioO4Iv/FRdQQAk94
E33EDz/10Jh4jpVFEBHzWi9OFHPs8YHI84D0nLVy1oXOxmay7/edGXPGu8ofgXAW
qscYJoD2jqur0Qwd/fAAt2J/XlgbfpIH+MJ4HtxeNmLMwm2m4tEmQWfkYBtcqgPZ
WI8iYCKz4FemGJGRNFFJvEETbQ8ScT53HZioaUBP5RSwFnmq5o0NGvznPbrOtyfn
h94AbRJwe1A12oKAtUhQNZ+IsOiIvoAPHBmHycIEKw3SobzuP5FsogMvObOtxc4K
Z4x1bUQ7oRthkBxNzT4rUZ6OWprwQOYJCacJZt3aMuDsp2Jpz4Z8zQndGZ2ENq2X
LI5r/pfvO0ihK227WvSgB7EcQOXc+TG+2zGJTctgxRo7dP+Fu4BTgIn2FrPvjvaK
c1222oT/9KD1QqDEZ0OCv4bgM95N+3xTsq14aqtxzdtZjIv8ATBXjeqJ3rF71UTO
hrYiqtGX5IbvyMATHYqNTe5KgCY/3Wznodvs0UUicOTwOWg/AlrAEyXfR7PBxhnY
EcaZ+xNMgdizoUkClc+rmICf38E2BL34CpJIpHLrStDqgnPbisIHwDOOdm3cRD/v
m1lGC6XrSkrIrP2nJM773iKi4aPgKZnNfCu4vUtn+WQavW2SvmkqUuVzob7XrQrc
Qsm8XWczhTAaMdFe5wH/QXI2Nj3N9sFRv/vz1N4oENz460YAHTMaVyAB8xNjttNz
UxpFm76bqm2OMXF4X5QCBHX9VHqOVrW/ws6yv7BLhDyTa1Ftx+euzfwqpJ2ZOV+V
SigOsSX+2wIhvGuwpZWSg6U8uC5C2RhNRlIvqihogaCzM70WFWvIV5oL2o1Bnoue
McMeJIn4bYDF1LyzxAEyf2DGB+iMy0GTL6iG6Smavjzk2JcyrCTtQwzxEbVqFcmF
gAgXO720erlDgXGUfsYRqGCoQeAOpFvEKwO/043Y0zp9Z1a8Beom83ooFjNiZvLT
DmaJzDDpkgT5wQbPzFNIfd9ao9JOVsfWvCQWNMudQEzsnidOAHyArgnJ+2l2/XeV
1nKlOA+WPq9OTcLF3JUgq2xtz1newKdg21tY4jhlz4VU22HdvdxGlDiIR9BeY+OM
yJMTBcOcl1o/gr7zFPqvcu33GsYCvm8KlJcuzBHXpKCgGKHaW+ZWeHHfdS4R3x62
IMN9QJfN6OaWDMMk7jM9DoJT1mZdUJ7NCySwQHW/CSrczts8z0Gg1A73zh4O8vOp
K2d2+3eVTL8KAJr1PlTiA+ROug6UEHCrnKoINBIMBkndcwmowgbq9gv5caEVEp31
Y1f7W+iEqJTwhny6+qAltjZvnWxSMhYUFzyZ/jGYIlN0X7OUctlIEyPDWS9X+WMb
puRGoZrF5WMy3FCfQknSdeQ6DSD16KVPRbpTdYXQucFqLdrPufMBfNfyG7S5IeSl
CY4NynDh5jjUW6VDJjOKCusxb73FjxzkvjrcGxrAcYAaJ8c/czgM06oDPX9tFOMu
hfOV5Wv0eiOxR1gj0KaUyo6Fv3gGQcKjZPHrr1kUnvdEYonstiUU1Opn6NWRimh9
ybqRBrd1oYiD5V3QJI5lJO7df5eeogRHNRrmkazqJM0NT2DN0HMXs0V8y+zp5EX3
u2xN4+WCUtANc5bPILgP+uNfeuGODdTABC7W/7dgmplMH1z/c/T+tT5xeg5K3o0T
lWw+zmN7wrb4tkJfmtEHSZSUmsjzhPxj9p3tbLNezLjCWtGUeHy9tPzMvTTaUeqv
AQaJKou+ICtll69jI5vhNuj3LRbARjuLz/s2/vlIT1xTviRXdJrHkiXgtPYKlpuO
9GUyc/gO6OIQ2COIENmKUC/NshAFz1ExfX/TDMolE1EDxkK19urtSkTR07ROEVkH
7i71qBdG835NMv98yfC667hsUyXTHHiayfEwO5z81vFYDvEjHISdfG8uWt8F8pWi
jsY44wjJZOLfLU8AydFNJbWKxhulImaHR275bwq3mc7GE04M8MF8FjtedtW3KU71
qGmCvEz34y+pwV7NGLYBheuvw8o4KYjGHwu+eJIPgbTET1oIH5n9DZys/JhyETb8
yHbVANxPvrk+hjD+13JbhGDTu4lai86lvo2dlG5eRhzY96WuvXN6Ej1nEGizu3bu
Czy3aWdkL+YGRWFAvf/7hmpr43RFOAMeTjJERlIcJqT15pQ+9XEyUETwAtZa2rjF
qCgkiZi4Q/1FrNKpJoJsBZ+b1IFAUHgE1sOz2T5Z8HprlKkAeCusKfcACQVI9wDm
R0UP2lOHNy1Ixh7eiSF1Fl6+Heq0jAw1MEi2QZP9PgqaIvulfpOn0wK9YFrjdHoK
B/g9sWVLN1SlluBtB9V93NFvLW0q9AG8CCYUiJBtVfTO51bMA0B0LOhZNbmh0G20
f5FmJRJIlRVD4ah3jDArFC6vDzu9T/sTvlFhFYj3vgixNnkOFXdyWZtRIx39kLZ8
67S6h/iw7ZtOKIk84kMmrdJMf/Vps7S1vKrzY6YBPvitBGNkynvew8yU2xMlxUun
ejSr7KaDMIR3yvOTblQ1EEnQTd3gUt6F9q5ygrKRjBmOOP8iexSgZeKoXDbzIWaq
/UV64v+ukApr7ox+sjF+BbJZPRva1ycaYT0uOiwL73GQo9NjC6g+2Uk7OsbJX+pM
qhxkajsVUJ9Zl7fwMuRQON77VxFDuqAq8qOQEw+KW9RC9RmfLK0ciPVGDCsnszk4
hjIA2kSfBBHXLbyzggikBBrmKSvRr/sbDVWTKP7ghv1CU/MHsPvo4iAGfIQUVRrz
qdH0qLWhNfD5gagLQK0JC0FLzXa8HBboHWwjp/saBHZPJ6+r9CqNprtuhWqatVJ5
FKLUQLOjTWQ0OtT8cuHA1RNQHTYSuO7MK2olJ1fZmBqpEOWUspZq6yuX3/yQnelU
ZKxND4roZrl8b5HbOagIPprDlVap+vBCZKs221hdj7dzTIYyS1/RlrZcNeZTcqAL
HRyfr4LdK0+s8QzISB2sq9j/SuzvE3pruEnTyp1azLRy2iSm5yRGFtG1V66sSvBL
Pzr/7SxCHrM3NCVY71fb7hILtuu6XZ7qniYyG8afxClfMWoMgsjgPJmekKIw869E
5ycERMjjOHH5qSKdUfOwWsAQyH01qbEXSv9cLUXTGdHy4Bvif6bK0vvmUuwHM0nW
inqnKOIOeee8z0NQA3q0wAzeoJNvdh4OJRk3lGMfi/oVFz3UdpzVqEoZHmmfQFv4
MnU8ya0zZ003nHNoo9921NJpldwhCroZ6Aq+c1SuMG3/4BA9Ydx6q0MrUP2U/ybV
z0h0QypYqTMueZlMaC4prliWlaO0S1NKWJO9M7AYRtx/rZ3WnfinT3IlSR5nWmZV
7KWUbCKASTSFhpRDmfKfjOOKbQhg1U34oT2UjPl3ehPPqC5wEGcu9PhHrSsGZ6Ti
14creL/GDzumPdCBzJ8IncZS6M52zqr6a+0cRIMFxiCG5IOTedB1WkUhKuECVykp
ZqUC/KqMaFPETV8zaKZxSr3z2vkcG3mjzMwLbzyxaV8fCn97O4zxoNMCB/R81zSs
7pAJbONEQUaghHpPDEyJ/MapomugFsad4QJWHiYFmj7TvmXErtSxeUn1if4uqI67
T/W8/mYqEs7OOIEEOB4YCmEUqsOfGnFLQeWvK5Bx6eOIW4q86bN/64GIZdSvdVno
EjK7faW4iZSO/ZIQSWM7XO4TY9cKm1ETH/o5GvK28EAwPKSGmbf/SuVciWps+eWt
ekJyki/qVCT9hylgadqnpfKpaXWgIHXJ6ZuRiqzTcZqmE9xZS0SuD0vij77ZsE2G
Sun+Ehfq44toSvxoWWV5W2NxVRIReJUSd5PKqdcz4hFVPX8X71jF5/zcf/ukqbxb
MjDFDfNt4WV4ayDQ298T/mqQDCz+GogMFFYc8WRvzR2ACl0DuBgFOU4GBQoQLJ+L
JrwKqqZdhp3VteW2R2f7VJuJDwUBJSRjOhYWN+Hq5WqphmzY8hy8veFH5hlQBo/P
oBCuz1mLijkfqrBLKTIqAXwY2Q5NRWtG2YhuBHDMf0hRZMSxEbxgWHjvLnhf6YTQ
MlpauFjtcstTZibVYAII44PZLK0SKcY0gmpLWX9LRrrZsedWO0/0pdm3kOtV2Dp6
yzBH6GL6Irtfiqz2ispD9ebpcAk0Qxd05ngLKUjeSEQfL8zcXOqiN2DHE+2gTV0d
mlqGXlhjnf8g96+othbx8uZ5QkUQ4eJUdosamZwimVyvF7xKhnTZAelneS+Vaeao
BXPAME8Jj1yEvdrjoZiP4TaXQp0sjqL/+qZWFN1TKUFT9WrvL12hARK9y+TMCbzO
qWQLYknOpV4bqfMoAPXdVkx3hAOKSDBqUOcCQzNm/7kNLmgFtmjYc21mNN79pWJP
Lh+hbLXMpGkM+ArzvQuXllHdPCbzrMrCZFTrtzPFv2cThMvsXLnc2xj0W2IfnuMc
dJkEiEosfBgsE0j3J/sZauJJqkE7dUWKwa5RwD1sHDqGB0uPCbTP8/gHEchbx70f
vBjM7vMikSqVrb9J5dyBCppmZkWUFpBsf2u/OznLr7cPtlH3/oSXJftKE9qAMpmx
KEdt2m8rjs3OWRSFgiCyZSr2dOVa62N7vLvZazZkfnnZVkKIw4xAWFCW1+KPsrUH
iBOH+9b/aYG+/5kD8a3eqLvIicAJ88oYYZL8MywSwObkbAeKtaz85oRHjRJYWdPA
zfc7xnjcziUHyW/Zh8raoJgCFhEI1D+ClEBK+rCXIniEp0tNx8MEKtUtxtE5XvPF
+d2qVJCSjZ17I2/KhPUzB36JW6bNsL/1YP8pUYcdkT3Wgdbc3NO+FRZMKJfY1j3s
WDSJkCZfy7P4GqJ4kcl/kOk0gZkx4Agi1b23fCb+kIRC01O43ZwQ8GoHYSjzj9Pp
C6WQ1q600UtvsLWFSrG+U4buo/dyoDHrK6M/kpFjEnTlcIUM4vcQh/vTpYxDPOO/
mLuaY4T9rEXAxAyqeMwUSZnfD/GXT/BUH10m1oxsmr9mLIw9xfHhUEFLPbv5Bdlj
reat6P27BUd58p49Tu77xn3VlybBdwHyJiPjpRd0hJBS7uCIANn5dhTlMsSI0ECO
sp0CBpVwP9gQbjJA/Ec8RLBfT2O6kFDBrhlGi3KGjevjHghrKuVNpfxvBjnGGwM0
TiJ/8LCfcL9setFryGYZmHlRp4Rr2ugJ/JX1DnWaN+SnCDVSR54jiZjJ2GwTN/5h
CIUKDmsaDYAAGUqug3m5JWEGWAa78Yk6biDS+7ZA7UllwU4nocq/rnjWKhXQxx4q
KgSBT1pxGCyRchJI3ZLx2L3wdYXj7Vq8O/u9dAkLxaeUWLm0oBZtmRzasjlqFufX
pJdKY2yv5fvChXo5WZ3rGo7zhqYrelDXhF9HQXrM+HYuT0r8aUyeQsuIG5M32R7o
q98IWXJDShg/yUbKdqcQ5IcI/QAyPbzNFcvEJrw/fByuSqK7etxqr2fIs3YR7FcL
OI2iSaCezYJSJczOFQSVO8ipEq5Z9BnRXoCO4SITJjqRvTIbdzB4lAY/h8SQzlrr
HK+fvfJZuNOICQbyE2IFTekBqc0gX5VECXrYoqSjmjYe8iJ5FNXrA6rRLSrJK6pf
Zz2XUL6ZbZFErn/ec5bHSk/eNjPEe74NdTi3+Uhf8yy3A+oFDzxqwOktx2uPdzE8
UnqBLsn7CtVb0CO1JsqifYivdLopHFo5UkccJ2P9Od+0oDhyXCfu5T+Vi5gnDn3H
TR6o0yib7ZGSw3umn9LDXr8UOxhOx+usUxDjeARwvBX7Vcfwek87/NHr8afgOR07
M501oHBz9iZeNBvlYltLeSeQmA2XLVHgrjVxcC/pf7AAdjdqu+EgvlPXiqKSoyFN
mAfYNu0WibqXvNGdo5aoAKXqPtcoeJUuNLQ/nwpHeNn1ng0tpaCttIiDOH6nKPbc
hAS2e8BHLg91Crg0InBL4ss3p+nR2gD8QQngBYtMwqPfVVKh+S146rinPf4IcbSu
6lOH186FFzL4BWHXGhmXt1Na1zN8l8UVXuzZtZO8oNmdrqNJpSez6mlFkmaMsJRI
C3AIW8M4ByWg3PPKRSg8kY/2YXRVBLifi+b6yySUxrGbq2zV9Q+3S4q2tXrj9ENL
2GAyXD1Y+duM3fDVkg6w6i2wdE5ONBDsSNBCdPxkdyfqxS0qtp97px0tmSTnZSP/
qUBoBjQtVCQCPu2vlCp4iafw3IMrGqEZbzLQMkQtQMn0JXM8ypSLbM2MatuMEHom
gIDya5GQJoxepYAFx+ZHvDWA6D0gjxcxFKVggZ6+o1w3i8jeYe8CN0j9ekooBQjg
Sk0EgVf3pdHAnYkwnbXI80fc/g+i05FVh3JZUUgUqvPF3HcgOPb6KVDCv939ITBN
CU+6SkHkeyIR1P9RPB7XblzrIiXe7aAfji4FZbOscAngM0WeAWKYFOhph+EpouIB
vbwmondmOwZIpbZjbFhcpyz6Jb5b2BDDnJKR5Ded1NZYVJ3ds3KGwQmqoIjhaX3A
Hz/l7PyboKISKC0OY/C6a5am1U0xzGBgntZMbCxrMzmUEdUNri9aCAVJO7tWcmko
JVbZREEnf4IQ2ju7MpXgQFNdjWvLOE9KrvHgkz/tR05gbmqAm7ffu7i/52IV3/Cv
emsTRfFqJ6zM578z+CK6sfI5ZwchP6SvSV3+DQMaEWHupuNvZj1l1gciQLHpw69+
kt4AoE9x7svTHll+2BPveymPD8vkF2nIToqs2PBjh7nNuS+QXuG/CB+oXILMqe/u
qPXRMUTHCA4LqL+5CA4MKO/vMtxWTpISl2ulUi/WdDNhEeYJ9KLEFQDnJXmb3qrl
9n0dtBMCsLX3AvQNOh34zMsHGQaeqqYQJgkv9Rb1hxdAfKxziaSIBtmj7WmKm9sx
bOkvq7SnBmDRoHuSaO+hH/0iUk2uelnF7oNX4KEEjwvZc4G85Fne6XRXDqm2sNTt
Il7z00hkGvrWuMld8GvQUNeq4YC3Dro8rxa9jiwoXAtSJ/J6AQiF2HNxUq8A8fTj
LCeIswcW8o5q9BY6yX6Uq7Gre6nT4i52G+DUA87mxcjuLfLDIt7W1+GMQStCy1Am
y9r172ynKAIMJJSat/lJ5TNPjpXDhzQhmbZv/jDQAx4EhlBuZNzr7oggtK6QK51o
e4vlKZn1jqsFb0FsWoNZcnHUY74co/imIr5XhRs9wm8rwosu9vDHzXYOYh1po3Fe
nQF2swE09JRAvnT+mR4WdgFmRAraXrXaUGNAat0SDCJa/+L6QZxZODZfUzYyjWov
ostF05RIznKs/Zof9Ik1Zjfv14qRTNCFrSHzat0z2B1Vlqku+Z2bVu0y68rKI++M
NtomLJCeQtONUNmhEb7AwNk2bPmdqN7wwF66YHkPWpqhBkWWID53EVsWS8mcs3oh
v1wKIfhSCUTbHzAn3TG/BPTvmeVo44UoBAheuSpL+BbBJrexiNZUGW70CYw+ecu0
qNqbebnAoq2fkLnVnbqyZv2f0UMN6GA7jmHxMRD+r+pvDqvhFRD7/IHSnkf66K0v
jb09JrKkTf5bAyObIUuoXbEfk6Jx7yek9vfdQlH0Wq7cOTSaVwArivuyFlV5BK3w
VCXMs/jhVIEnmhLIC8FJcOfBR3Pq2Lt9poJCDL7MPVFiybmHwaCvyY1WBeNfRIKt
3k5hpVP87T1c/2qjOFCPaEbWbZWIWImZu3bG8ZEQdp7u2xHyOkkwyi5nYzxGWYhJ
V4gbqyVLg2qK9gN4cvJZAaQk6LCjQB1g9HbTD5DDmBdl4HMBlOSI66MPG13XOEv8
xcOyxtKc03Z65Dbjgiba4L0nZjbrjglvmtLXqsrOmFjmpKG8Lzc7MQ7ifqo5N4vV
yqConZnNr6HbaLD4Lcl30TBgRMcAX6+7oCsFEWrocdCpB+IaU/fhrXtri2gL0wll
GKjij95rJe05LP8xnebIb7V/b9GlZg375ItvxRogB3WSUkq9wmaRPwM7ZzQ4qlH1
KAHvQoP0zx99FORGMXg0uvaBNUgKS1SBR/81nwiBxtdwPvRcikFgVJkW79ZHspsY
4mzR18t3Lx9RqM7Okd0Lol61Zyr9ed3aX6DqEZqCfLDo5NR+yG7DtCKWInBQ+GiZ
QcBx3KsFsOYxXztWIQtExs2HlTGJ4eDCIudgSeWH2JjfiAP1X3SM5CiMmY+MORN4
rqwKOETelt7BaHSgbkub9Uc0zzteUfw1G5o4bu3KBFOJtb4a7GBQSLh6cBi5qhNA
WBJVt5ZuSq54zau0CtKnQRAqHYu0ogTw/piAc06fJdknJAaZzE0rXfztJq81wafZ
oN065RMGC3rW9Tj5q0a9LBsD6lxxLAd3vFQ9WYdcPpOWfhcEiketYcyb0iSR5pr/
8BTFi8duEBZJqo0ZHbKEmRB0lGsuk1iw882kX1Ey34GoLR+U81m6QOMfbMCmVs/G
cnOYtIjxNLDfeDLTdMDVHSazVU01YZipneO/Lt6e0NO4tS37H31lXu2ZeiXbxi9U
sGHAsGwOzQAEhykJOyMUT5SY2JwzqgP6nNAMVYhTb9TCcTiXjGAw3jSrWW4le63m
nRVkopfYw7+pF4/vowGLRLGrCCl94rhJkQzKYsnx6BQbtKbBMz3ikxuhKHTTFoz3
tbs4/naEa83e8v88CaBYUlVVJ8lI1h4n6HcbW3dFGCYpXlTNGWFZS/iXxor5ebOX
8bf5bPVTC+ZphZ0iLSBMEmiQGs0iUc1Lz0SpT61L3NTAg/7fmn5DJ0iQy7YE5/Sh
bmuUozkq1XiWkXm7WD3sWiQrHXI4iDBWytyMw7gI57BjiejhSetamgN5iIVcw3Q0
aZfF5qVjX+USufv94yBFwXIELrRKnZbL8rfcAkNz0MmE6NMcj7gMiSeD/oqEtHvL
hA+rOLyYnp16snxepSO0wamVOYScdwtJKEQHgU2jjypPgLt+pWbvAnXTt8/j/i2F
f6y1MbPKy27GYg7M6/lu793ZXWSIB/aVjDwXnJqSOO8tIq8X7wRtkhNRpBj1WcpU
vaZ+8QDBWQaXJFU1B1kM2KBfBd27/enCvJGFdAGGnD5sKiyPd+v08MIXWPIG1hbv
VK/spWESeu6d0JL9InVCP/ZwLpk1vO60yg9RT0iwbmr86LPRKlnjIIQG9B9uU2vP
RQ28bvKLRpoyHwU9OOwiUb1YdIM67sRXwnldr7oRg+tc/xsNLl4PA89I5A0CKeJ3
D1HCoqe1TpP/Lin/TEyQMYYry/roj1PZZq2yep4m+bNtAvRk/j+Bypz/zn1FH5/3
SQZ6uh94PjA6OM11EbmshbG7QJC2hwaxh0Yi4nf6ID4NHbCJFcF4Jgc0PKm6U+wk
U7g+BSJnagRn87QSAQVL2P9AxuuGa8Na2PgzLLomz6M6p/2Dtb6n2CgrMAkqlnI1
bgHkMIq3rqXdgjuVnp1xfyFbkIa6IV4w0/zdtoTbDVAfNpLrWHuDfyT10YCAQSxb
yrnMFfmNmwYOMKql8D7SiVhF+8CQYjohoji+180/94OWCquKTzG3RbgXuoAjxV7V
0DAJrqoOxr2bGFdNrzhDgY0k6a59JCAHc5iF7lh/uitr60ZudjoP4XNl/jG7A98b
kDzHl67H7qh32ue01Km0Ny0rmXMMkN58+G77RMaN4OxTXTfnz0DTjJUljAy0jsvf
6eILuyMDEAyx8/WVJu+dgpMiMBqqJI/8dZx3yFulSVumD1KyiE3HvoozgLAexdqH
Wpa3k6QWDziIb7nMOfRbkrrK4OVFGiaEeUL6KRdznzlVyXLxClfbyjQjJFwGUVys
fbMPe2zN6pcemsZwjf3+O+yUcU0BhHIga/Lct7jr2igtx9g7tgdNwPH4xKrvNQVJ
k9UW5pSNqs7FhAMX7AcF+JxO+mEN9Wy05C16iO2JhWmk0XtFzTEvK4HbcgVbiWnd
NDtRKh6hqTQO4KZmBwk2K2I3KuaqLJoMhuv9KK6DmONOHBXn2BdPzeq51Uin1Kcy
dzvY7RT3EB4wpevUrXaEpDbMR4hjucR62+iHGZsX6G+xCLNCpF7K2LQ4L97RREM8
vuSPCKF7rEH8rPfcpMpVyEl03K38j1FPGzAj1k9Dj2njkD4Y6HwDtZtpgo7OYnLX
Gk8A7s0mnuesxHTEX0lQxgSU1VmDngz0Um9XgSZvFQagIDWzvVzA3qmej4/XzQ6k
iKYrAjY2DB5v6CZHQ6jvHkPtExLj8Rlu+z3Lf2UVJIyvIbr/DJxO9m2HZM15dV7W
aODKJJ6eoWDUaKgeq1l25u/wwt52T9jrjqESL6MvFFFLTOc8esTMbVFHh/rSgKy4
fOOS8rtRTW7PrrbFSYed85WheQLiJDTOnlfKaeLCSAv6U72cFWLvw945UMo1SQ/t
lCmS1KEioe5hoY3OhViNZI9GKWuhN5CVTRRzyyT3JnpnmRa101uTSkqKGzTBMX3N
Ey1suXsXk6KAz1xgUAdVDBdQ+9d8/nrkBId5MmlQfJMloakMPq7gunTCQnksxPZo
+IsUKJjT8gVZR7qZnmPy1+HcMEX73h39wydeBw4d8LmgQwDLu3UkklC/2h3IhIlz
RNjFk3eq/FBUPjgDlIPxooY5aO91V2rAT2OTSX2HE7c0pGgjxJxCiPx0W8idzFoq
7dM7ISaOHc3Tilnxy7y9owgOIR0O/aFp2ct596II7tOKppGbstgT53l+YgK3GE27
1uLjPmNiEL47pBBMY+R+M5JLsqNBt33rs6lUe8TsOCmbRM2bpdA3mLAR9yMZc2HP
xIS6hiL/eZfwROaFuW7ZOI65+X0hxsRDWOhxIPtwS0NCAHuUE1pQwNIHKs3z/qYc
DGiQDTF58ifT06IwK1J190dif7xqPYLQ5CTa32o5psKpxH2quAncs/dou/Z/Lbqd
o/dpmXtQSF8PDbMHmYzP8R3oc3Ovg+GKvw64PCI2Ydyxs9C644ymqYM1PLFFAIYZ
T7fXqz/VpaF/Tgc/yyhEVWS6ROShqVjIuQK8tUAY3MP54S0SZLVEYQF285J/0q3w
teV+1yAFb2j0ujhTUYZMdcVcf28k36XNZUhSFgFvCMvTDC0myfoGReebeD/NLj9h
y5MWlk4M8DKbFbAtRsa2V68k0g5maiFZlIO68I01Futo15M3yF2oAR7OOYG2Z7VA
vs1tqC1sNN/vz26pAcPV829/RZKn83QnIhy9TPVVKSQaCrYe0GA30SdKrPqU7aX4
yffQBWh8v01Er2U0QKIp7iAiBPkICXiQgzEGdF72nnnkXQwMhcG2DFqJnTCHRVGy
y7VrzmS43vxvzkfnEbotUQfxniP8mDtsCIjQUZbj469H9yMgjA6OnI/WJqZPIMFB
PjKcsHKN4vjMucCxDr2r3A0jJ17EidLjbjQ97Vb6BHc/wNLOKKBrgKFlL9jTxfpd
iCll6LLci/FUQGEjvj67wTIwCe57xtkDo74d37W/G5NlLXbqMIvzz5KNIJzVYiD0
RFRt/nobNwLvqr00z41lbPD4t8+U8gcRSqNQK6ZIbH+SjhM/pHpxkjwC0zwS/RrS
PHhK9nE1BJMXulazYNrQ1YzPN4RBubfl+/RJiCGYnKwIYoPe2LvCvGTnso2oHAnH
YOWeGNnTOlGBsP5YV3tA5B73fWTNMbKdiPQmbNH12+IIAEc/DbXRot9e1ecUZ56m
a0LEYH+efu7WOBXSgG6oWT9S26FlcoWuzWcXmClpa+24kF5qM3KD/qYmDXsyavHs
JOg+G+KFl0AVzZrShGIX8/HxDEmqL9UihTxOD/eZonneCsFAiuPkIvJeviuQ5/EH
c8wqeWnyF/5jyw/CYTKGVUElRzloB29qb/xGZIOlOAeUw4AN8eJFXljtcVVQlmRV
Wlj6VMxsfFX34BzzqQ4f1FCYk7kgSxbHy4lTxjALwhJafxqCRqOkren/wsbrh75E
SkWCZyGV1vBNUDXNmHrnzypEfQn4PLlaWD3bTY7pifKdXs3JSxh5sk/lAx5cbdjt
8/14O9cRZiPlw30TPyTzvN8vkfpLR7yayy+24kNnaIfcOTthxSCpTFZsxqT7xGbu
f10kDv0SP20yo1x7ZU2tJkPUReOCjEk4vS6uEaqddfZAjmxDlGf6Dhk507YJHuKm
lTnQmFimi92bDUSXuOr+HItnGVJe0I5uPijAoP4EkPw0WXGFlYAT7oXK5kC+EkAZ
AOFrvQ6WJUHT34wAtphriGwWSOzGBgCKj4mVC8KqK5/1nbZZxZYm0q4KN01Aqppj
3Ryk0iv+x3oVOJiV6ZRdecW00OHaegdFSEPMnurog2GuE9YR7zjDa0D6hUekIe4s
fBTDPqyUayjWjR8dLQu2DjXe10OcLelFlJdauXwT3ZDE0jzC7KzHs1BKWm0mfQnq
/ZfAJBk67TI9LVhJbI7/wA08V2hsDvi8hT45BmG8dwA9USs+hur+FTH/9kxuuP/j
FuQLgt4lmWWc8Kb50ElyjhLzRosR3WwhODqJ1ZOu3vqbEHF+97QKviEeTDtaXYAf
YCvDOAg7i0rcZiAgkufUCLjgIpDbEEPB/1CJNAR6LFcH+8chTfjT66vbMl+gliHQ
ALXhLZZ1WlgH9plpVNiHWYzVERcOhYiHjKphOwXz7jEg312EDJ4xjORrDHJf0KWG
Vof5mO2gsz1YDZe7Ilh5hd7UM3Dl/Y1Ul42tSuEFjaOkykBGEGq5BHugzB83vGpe
I8BpDNLuXI/UxqqHLgd74wDqY9ouTOUGg2N3+QosfKLoQfBCm3U3Npv+KvOpP2DX
zFy9PNCRQL5D/GDeh9W9U0x0USegDQsOtTsinWId/F3LVKftq4Rp+ikTsblSCTOT
4c8pBGpxvs38c0c70mxnZEof2Wl/ahkwEp8Rs89CUgJ/PYvjVTy7dDPsDkYTBMhI
41dLP+XuDA+qrDw1omZiKkAFK9j4cnyE6CUoF9K5r3mCUGmbGV05kPU40ckv14DK
ti+Z7pr4WTnUPdMwf3V60JiCrvA/171oAtz5cknWKPC7t01R9awJCw2XdXDyH51l
NRIrkhiVYEebcPqKG6kXBr8NXlnum4d3TllSZKAXGy794bO5YFhBAGpToBm/eBjq
pNkIsY+PC8q7isVh4QByikuJd/T8d9Zd6UmkAa4Afi3Y3pjf1x6aYbmtN1Dmknon
2d7t9ZdD7YPxDe7Def5dma51t650APdqQw6C7LMHdSQT9BO1HO7ZStmsOfRMsUg+
cTQL8sEmHYDHiOyXvixR5Lq96bxi0CKSupFpxjgWKbHO7Ws3yyn88TEsO+yYzD1F
ToQI8f5HsdfqgCWKHJny0vrP5E5Co98eNz7ytP32+wUiXuKhzuSW0zFMWTUwTajx
qplWByR8Zc0uZe8+kkR3uaekvCC2IrFf9Kjawmk1fJzKa4h0r+LR7jdsozP0xQJf
2N4gWOwlnh1V1EGdDLfxScV9xJyUOZKsqamp/jpyEgY8RbqNTxHTB2Lk72istKxZ
xRBVeNTWLeZhlgsfgWueMXbjVrrPBtRpWwO298Opj6AMMDhpMNwiEMhUNK7rKtLK
py2peG+FyK2eh6PpP4h89FWY8nVzGBUt69MAqpOmdQ4lBlKfzIogW8Ej0UljHWyk
1QTaZLCryHnUB/abwXygwlebKxdlES+jZ4XSlH/c64f6xjKcW0UAOaEAawTeazuh
1r9pQq2wmFfEO87hzXEtiVCKKHTP0PG8mhcI5lxbE6h+1/ewBdCRBIJH1khS2EHh
rHwsRY1qoCMMnaNAOFFytq0Ng0upGhqJGkPDiX8whNynEXyeR5AOtCKelyeUdUjm
G2JRygThuZNmd/83IbJdxO9zU0ULK5WkIDjdfSFVoFPKKVGD/7e3zWkQXv4jAIVZ
TvEFiJe1oBX9H2SBdFzm4ESJ2+HJ4Nv6tWTMGfWBPuSgZ2oYhGcn6oOoV6buylKH
OJwoUqV+cTmIghkDsPEr2xfzCAc2vwxJpNo8mLWFxjLAq2eovPv4u5L0VT1S9K2u
fsZExCOE8RwebUYwgxtPa3t+dw02LKFS828Wt/lU/JDpfm0KckNW/c3xcaq3AaLB
b/0+q6/VHLtEHlcqT6xtq+0dNQQh03scFynuEHzVbapvERX3s0gbyHBlTqudonv3
DehiP5eXEKUN2KZuIiXEwUNudY4wSXskSC0DxTu9qYuDn2dclzsFXEfVtdY1pmnK
JQQdwdAHYpDqjWk3j1t3X41cCN5HGkqipn1uH7tw1mxWjsMzh5ZO5vpufUx+WeoD
nw9fNGi+bl4mGZMT/e5FIzyXYr4BNDvjHprlfRv5ngRv/mjS4VocTL9f5itkdS/s
HMRfaLkmUikv23OazXlLQwVfLYZAdSkq4gKN+UmszBuvplDNliGmXCg5CNhL6G7x
6gYxl41jcL1wZKAemvDr/uuruVI1PrX1wCguddbXPiLKL8FzQ492x6C6o6JgnjjF
+TKbxvTSYTyDOXa/FJmkZ3JlVOF8qHaK3qdJgpMiVCahQwAZh4KkOeF/R9lAOB0l
TT+RlLRbW8C0UD+Sp8h7rzR4zR+2iSOS+m9aV66MjAWXX1bW0YF+oE3FWBJ2xFIN
ISngXQ8qIFbXTHSEmLu2NM/335tg/CKCCrYeyQtlYDPN+LwzkK2JqYU1K2Xh6C7s
TYd80oTXP/ZV+jpFUmoK9DB2bcKBfp3yX3oP/aHQ8l8DmxQECb2e1jM40vmMzwMF
CmW9+JmCGiLavqsfRRnK40oqP5ZCI0Xuu7XGEqq9q/N8LgdVQTOrp48QVwpKf1FG
IkBI0/OhVzsgLWcd0b//YsScPHde4Hqe4CTnGbj5DvPndM+BFYRUgC+2wTqKK7Rm
BwUmsxvJ14TkLp9yIEN8J9S2cxiGcY7RqmaVmrtZLBGcmGfn2q4amGJhEpzGqT+2
Z4FomxfnJGkKtWFWIYERyyR10zy53blP7J0pCkUmyqo9r9RPTcDhwErh+bHF91lG
DR83L8m5URodCILtuu9R6wPzycP4cQPU9vjXgttybqHcyi43G+hby+SnVTPatrBN
kUtXLZqHGUu56iEJBfEsP/sf8TNRfKaWmp+28CzzWyJOiWrGoqDvsJSrPHz6GwS3
ecQR5k1FLhU73tlFOrcURDAyH6SME4P878AbieDObfx5uJYAEfCDM0vPStTBbITn
390kUIBJERWl2Auo2yEDXXBs5deUEJoj4Qkqm3zVFo5kPxuTUiPs9ftjKikujyA/
5jwHylFIweELGZmC+MIy7otbc2yVb+zxys/o0Q8ob63ZDRCswteIjNQ0C9206x/d
thYgt7pCtTr/2yeoLFf037xLthMB5rWxgfEBHlJOqvrNJDt4IYWggxsoP0Thk04h
FdYV4xm1j/JUs84fV9EuyRf+KfYreVfG3kn3sNE8HB/iAZXlUXB14NW506o9s6mQ
ux2YN8ddSZFALHq8S8k3EGQHyeYxEMJuvge4uDxhMMPbOm5qR3wvsEU+uSHZkZF0
YrQwuQp5v9zBfr6yAWasuDK+EfhYR6XoCMqulRZOczhkafBO8CcpcDR9bw0QJLZw
fLyDsWbShBDkRfvRl61LThEoCoMlPFS8EHseGM1aRF72IHaJHMSs44T4ToQBfKqz
yoov6qbdFBvnZET7usxXmBENnIi7UdC5sDPj88V8/DjeTHBOWK5Yjbb/z4Y49D7o
pjJwFL2YSQn9SABiXY3/MTVR6mcs2EsTkmMmXFOPdIdI8sFPzVzEsXyfhGs9e+gJ
JQNXvTytMObd9cKotavpgtkG+W2PSybtt/Y0zJK5vx4Sfpuece/EZW3G9SA6gklJ
UpPVxh0T0THooIqnCDKpjaPOyEv3z62IoBFjGGtyQGVOyeEzrxSy8XoFfM+/t912
sHe23tCEZvtIsuTm/3H6Flw5AInqClMmmlut3l8ddX8QSBZd8L7laq0g/IgCiE2r
V7Kt9dsqbYgIn5jAMCmrrqyzMrtISe/bhkyS9QvLWybgI5e9tUKyOFyhx3GbHYep
KtLQsJw7XlWnepUQPysFz2vHc86nB06F7D+U0e1LBESoP+OmdKLXEsnZejR8koy5
A4/MFc31h3cEGvmAteBTsIth9LJVXd98S2M2X6d+8fZOTDP1cGk3sUItIL8nxZJK
nqphW9rPrTeNCUt12TPKmADLCn75RRHWPTt03LG+11NjVlovvtuezqXgZSM3oRVQ
qT8GRThFG9JfKGHv+rolZcvSnPGguKl22/57CX9fkIoFRtAJWt3gJ+x/4DKJztYQ
IjBJXascwD7pIy9rMwNAVrsKdRKpnaGww80ivOW0+to24irxAaMypI4fpxB8zLNn
avddaqjli2IqZkYh+NEa52+syxp3wh7oXspwHczQ00eiaWsp4zUw9EJ4oXS/WAso
McYVTk2Lqp7Bulfw/EOoGK+7w6WqHRLEMPh9+zhHsY9chImuBkImSiiFdB/cdWB3
zKF+QigmHEmNNyZQVYmKvw8wSMejqPSliLAoMyBq+RJxNVv0zmmtE9v3w7w8sHKV
bBQA9o7qVbhvdWc+in4pewwTOFDqSihMcpKZkPof2iitvEkQEdE21w60qJuP8gC8
JDOHFzrFFFnxU0ksKid9LpMQMZ7KdA8NByaXUa7EeR/ASS1zZomxZfzIQ8TpxFKw
lCS/ZvYRoowUCIX3ZzXtpIVwJStlEIFSbnkfRRt1OKhTWC8KMKn3t4Uf7qe8faMV
SYNcD9YJ2Kcope7UiJEHyIUWxW0Ji7rXjKmp/sSOogv/3P8yE2Gd/uKVli30tsJu
/KEw+rF4+SOu2HzLwqPEcYxwtQI/hyHDSOUMYF9lhbqzg3gs5e17xSgak46tXEyA
kmna3Lw/UiGVYGFdqqGpigx/HSA3WTfWfirVVtlT37VTrZWarQxq0fLfjNNWq2Do
UtYpxVgM4p8ZvSugJ8Zn9rDfQgur/r5yZsqYp797EbO/z4V3ODv/lhjXctOlzeGf
mu4G3WrFx0TDCfJqhJ5zexg13TNPZBSLQ/VLhknOC5ODjyuZNTGiLsqJfEQGJAOs
rugz2X1/hkm0QBNX0H6sfJ8GyBwQgOUoZqbckCFqXsRB053ndY46eqG9XGIk9DT7
DDbUK7dkAfFV9iGWG6uB6RHIhxrSgjnHfh+aWDSlT9rtEP/EkLtk+2t20t36YN5g
q2v0XPY0PGw4/Sb4S0PGC+BiQryN2APe3ze2lvPiy7ynav3aTbSGKrIfdCS2rB0U
qFu8NEWDpIhFqwF8giiSin/x90bLoDYqY1hQN98jnXkqeBnWoxCvEKqxrYEAvub9
c9wVxnekOlyZDaC7VloCA7WAfzHgiwV7sbmHwbCKG3JOXBZeMaFuciH3ZVVNlnRn
PfwrhDqbyA7fqRIBBw/2aM3to47NO4Ct6pTmz9fykLlzxz4CPgn8Ho6NDEsQjeiA
LmVB7lKWKFmg3YgPmDnzpo+GG3xbQqhlYYM3AcwPtFVDRv84hKyduxr97ogPDuBl
w0ztMGhNt0x2PbfDGcmOflY3toHqZkvQXcMG1srScuqqm9k5A0OYJZi/Uwt/fFoc
olR2RqX/fYyBXxqoS5m87+TdR/lshELjn0OLUcpJqhz6TOw8JSG0d2525im7r9R5
TRP9NNP+2208q6qFhQeH2/yBlxxHSVcIUTt7c5B5le7DkZhRD1KbA1W0RI4TwF+r
zIR2zSqCfFIgLR0afB6HcFZ2yPOdM25vxJr1gBfsn1DzzHnM1qwvEH+tMjeAWYkq
fnqVqDBxKJXIH9qCASPT5+tz5gbJsSpS3I5gCEeBOlhkihi2YddSWVdWRsQPFGg3
VdHTKjMNAtV9T2k5dp6UTASvEbtvuMI7xQiwgtvSnrm+zCYpEviAPafXqp3QwGRE
bpyohDF0911PwzBdaY3Og8dzasBg52VLF0gFIWAWQ/5s1gMAxZl8sT4pGZMeeuWV
E7DlhdtJmfmMVwO73Zs0NE+xGsfcZX12qiHa5ylDn6XDDZtEjfuWrXpDOtqcHMC5
LMYVPgSV9ttGeTb4jjrKm1rRPIcfcfJhhwwztbZO3bvJC79k2uqYrjtrRJU0Cq8Z
XbHV6eRIJDQpAQ/UegIN17YnDriBB3/3aD5/DbTIcEQ+k+Lvx341Niip/6+w9Lw0
Nccnfp3ruAhdi04alPgUOM1YWycBGRE/hLyQaaf/DR/BYXtCRIeWs6Z5A9pjjFBV
XulZ6Cr894hqYJg2Sh+TE2qhKieZWy11pJ9eekSUTuS75wH0mhTrZ48qoR5jpXLS
JT51XXD2Ftnb7Jow8Eg01BiJUa4zpfF5RxQMpiG4q6iuLMBBCkUjjzLNIM7nhLfj
sVgiiH9IuaNFuoXpT8P224vxKccx931aQ/oYI8u926xvh3IB6ILU5HTJUFIRNRzb
LqHROoYt3hgLYwvICT0wc1QDRAPJV87VvUIEfwa0H48mGk3tiYIRG62nwCFcBL3n
loJAVbNT9lsX29QwhCkR77NdViRhLnN/omTWskGoPbpukMUCv/bDUwnvuIcajMWt
GUe4MhpUePnn0MW6mWyFD0yCy5C+ig39nqlV2QayYB1KEAB9m3SwRxFltkzMCaE/
KA1wP1DNQJFgd2E5o1ah7P/y/Yq+Kd729Ed23S4+SuNER1qUMylAAofHBJNVBaBS
3zAbIOTUdnZIh6BWMNsF8aQeIn3hrpGAhPYfKyunuNwMvTgMviasxWcCJFxliLs2
e6LQ4db+VPOI5wUrYaDxGSSwRtWeneZV9sHuu/wpF0nJ+XSwXQmHbzTDf48YlVuX
+J+ZM6aG+ubXKw5WkND9AdWTL0vbcXeXlTMC3bcl3zhyc9ORSfmFTlQeKCAwIIkV
rMnMgMDsm/SRmCvxuHerhDHAlabIl7ClPRt6D03Z6Z/e676TiZwn0pd41D2x0xXW
mQoKI1TD5tSolejRh9pJnodBk06JQAwaOO09drCI5338O1HVQNRs9BBoJfpCUfHy
Vr0Kkfs4Lp2Al2T017Th55NAR9FlV4T4EHlEiVbyxABRXWH+VPGkbF2tyNGwBvDO
ox7L6a/iEjHhTgUCwa2yAqv7YBINt0Ki3cPettWB8LlJXXi8W3os48rEYaNHA7ia
Qzik5y/7cEz2ReW3owCRNUWC02NU5j9+wluvLoHzaoduYvMiIQyFUxg+i+J1Nxr0
bYjeCCmhW3zgXSVU2p7VHa5b/M6o/nAY2O3nNery8R/OXPefZRmDfM4SuEhIVLEb
+KtgzQUY/WMYOfCG7mG08VVmGoDgrkf8r4WMmV38LWW/AYBUPNeiG+oMxOUbL3ks
udnCAETITLAWhIqQ9IRC2OWZ8NJQuVgR3aH6JLSuI1TlzUi7UJUvQEAbJ2EO0qBv
IzzEpFxeUGgPL0RcZ2cD1U4BojVBGi1odeCZpk+RLRJjkqIDwsm4r8B7oNPCk62q
s6WqiLDIEGRHt5XKXD1Z/M/8YngXxin7VHveA9vyXh2CCQEZAKtaPt495cSEeHc5
mtvUgm/Ey8a56vCP4b6ZxzHHSYWizTf2e0AToWBR97vvVxLS7gHiBLcdsb7pgp2J
Dcg+5yTgDn5/C06NaFf0xveOvGsKnf8RAJplsQ6Rl6pzPCFijUJbOATmGDpfAoqE
2+qBflDH4qEqhuhZiGrziIGy1uDeYVO+6tbZcpZP6DtV9UQBXnBJRUpeOgKh1oPy
5nMKnhxa5cgucNAieVXmJiFmuHOFXUnBRrlJo6BxB5WQHnwDco5AgeQIAyRhVQSa
EKCbHgfrJWte6+lUx5gz0j0VO/5oEp5LxY46ZUBBqkAuyT8Xu3+c6MccS5rF6RkU
8+gul1ghi7l/c6NFtZ27c8duZIlovyXT+TTs8V/p/wrR8Qk/petTfdwwXngUQqpg
wwS7HFk9IJH2LEufbVEGuhhqk8htQwuerElH1uosvwmPBmVVO4A1jmkOt2OrvTdd
37p5eoMu2xtb5HKKsT0c7NpF0Qhck5+3pyUO4FdzNbk6qpaKsgOjLIUj2BN5vNRk
yfJ6xKV9LBqtpfoh65cHq0UM+uZISUx4YVJSwcrz67cKWbsPd+pxfd9ABdO+3Coy
ugk8TKLOW0oRLssc/xh0uy0A0AALtdfqg6aFQGlWMegSQnio9doY+UipErEmeIjD
bJJZ0zWe66HKMiqVVqesN3+8zBR0Q1/61DjjrKaAuYTt4VVOW6wotYHPFQUsxSoq
HP60R9UUEQEJpwNXptqLp7WJ+CGzmlOXlt/r11xeNUuFyWI6QgTdBd08qmYe+Qfr
MISkmnaaudh3VkzeZrZj3HsvrP1fSQaaZoywRfZeYPqC2g00WVWBFPSC4OZ6qvR9
wcxXmA0fmS1BWZHmVP24L8RUpRIJI4Y2mpDvLLc92VWZumO1FK9CFLf5xXWQRQRm
vhQDPT6WmGj+q41NAcw1HtNUEnI/5H0y4whyinBd4sBuLgOZE1yootZdMnn3qr1O
Ho948B/IkB4lut9VypAHuyUyCbF9mkB3JgIAGIRF3Wxtav25dqv1bJExKtrWmIJX
3EnMXW7o3u5XFMxxQkeHQwe0FZ5bAEeEKYqFp0APLcD39KWS+UNGGuT5ZWEenjtS
4R4tEUMjL4B8l/fwv5rcIBFUKWBvowHZch78eGUBQufqj3R745lnVZZ2BE3MZDUN
+dpMF9DXNOvLWJhdsEcVRaq8qTvbJFnjro6b/Z82W1vU5alTXoUgVnEpJoffuX8Q
aNhfNikh1MT/xP+oHfOjvSArmELkFehGRPrKO3SwsoeleHjOhyskrvM9xIiuffBj
SHIgxBNjjq9xxGiiLmx/wDBfj2d4piNEvthJlg2YaK+zc73LaxjiKuGZ1aHUV44p
R6EBgee7Bp/cQeMJkxzdPLZQUaTM9eTOJE7kFunPvND3Oy/aVGteMRw+fhKpp+f9
jll/lH54Euhri4vh+Zt587X7Ag9Pi7BBdERv5hMRTFrpfxdeiajbweHdxASU6sRW
4nwTmgVqEykGtcKzHZXDQecXpO9d29NdI3jwnlDW4KvCgX1B8+Gvbtg+DupEtWMC
RNYxPzgnG5I6lusQtc7MX37TxjcGRGfWPC12WDUConxgLifDfnb/7lpaRb0Iwtbl
QN40YDDEECTvEGTuS+y9WNmXyIWlwgYYv5nGGeCODYaqZErvDruT2+OZS2MhQyJ8
WJ/cYfef9AYColDFyMh+H9I805vUbgSnyTqGGgaocAdgf7wtbXLnFT1jbB57UhvR
8ilHxP1eG4M12lYTHw20Z0cWb00svMUCToaUJQanW1q61OEPkZmGVgvAn0qRByeb
GVYS9NmTFnbgAOzImYVJtqHGAwPHCMCyKDKIiG9hMV0z47WzRIW6a+GEd49Xf9Xz
EldPgpZKv54jwewNFuBWNL/EMz7Caicixs7oSgSy1QbmDxeZfEmINnmf3VUl/nTo
KZ/XBsDH7IcD15iHVBshHpy/cuc/GlJALcDiAektKRnO0xLd/FHIkcMO9tSI02O6
trYIuRlPcLjtBd1IHpvAbLdRmkBOaeOPbEDPJTgZO8B6U9dN3JLnnHHuo4ff8D3E
OmsKADNf8iFGH8E/yKXmHELCxI1nUClyQzAZi3AbwVTYaQ6vLzqNuCM1KTNCxQs6
rtQdAFu8d7fVoARhp381r2M4klkNGcZiqU1dxHE54b4O1H+9aVIlEVZbuXszB3Cw
LPZxXQa1nGRZAyWTQbH54p+n9BN0ykox+CfGxYZaLniGnJxvLfOVJQpBKJmPDDBK
M5rr2Y2QV/czIw+vEn7OmY0Hf+hD29XBdUyyju2FHVfwv1sXbqycx24JCnzcIjiu
XEI6k00X+4jbF9A8aUVwCnSi3Rd844G5rZOh8ZesEENgN+jHfBGd1gZWLfMI330x
mxQbYQbF62I/wt2s+AQh/kv7mNM68/GDXXy2n2U2qz/ZYJ8HJW9ocQ+IUN0dAUch
Xak0GAIqFN7AYaqpkp+W1GibhhwH/GUp8/iAk9sl7r858iEKC4hwfJ37eKethhzB
HLPFtZN92glpmtV290kp2/PW1Y5IBhfAwdaVcsoF7bBhuLCvGqJLRIqaQd5BhKcN
/8FXFkfrUD4wW+TlybPHoisNpfFcKhHvJK2ggsvPGsMou0N1s6NCEf94pcyKHdve
2DiUbiVlt/um91I+VZpDutsnhLu2M2yHblBHFGWvqA15bMksNK3S9F6sjinRLC7J
BixBr0AWkhyEAOrL43yse287q4wrMoDa+YcSqR+wbedstLAMwjdXSip2DOzOQDIo
iFAeOuF6f2fITcXBzU+Q9flR0twqmnchJcBjmZVZWm6DbODg+J3w2zRvbISlecpS
ydhGYjSnxxZ/rrEIan5DVwKrJ4YOC98f4fRhYJDfsfXLRrErrBq54wEuPSjcNnoB
3tcU1Xnvid+UvqTEhoMHJ/zEmpGvYMyLBkfssNSD1xT1WoGm/LhtNr6rHG8wG8Jd
qbHzwknl21OgYx1tr2QJTw5F0J1Uq41Bb+FNZ01CbM0hBLmXPgxg4IN18F5qYDV2
wjaMe8DPKFVIWME0giVvTZ3Y8d5bf7NKCEbXZnk9MgcWavRCBTL3x0wgcSTt4Pa0
uMRzPEvH6bbMkwSnOnC9VPwDn6VfIjS9hrlLxxLS6M0oxV3r0ynri+VAmyfi6en8
7bEuOqntYg04Dg90EQwZu4wxipxk/BYUCCSzXLwGeCFXsNRmk54Z+SKI4VzrT9Yr
mhpScvbjyxgFf9RdvyrYQDVwwWPYeZR/p4jbvdCZqd7cPzfzkyBLVxZQknukfaNb
LYv4FMo5gbwKC/D0sh9e7ACAnE6IWhOW9xf9CKsVRz/P5GgJFus8rci3dpTRU5fb
qO/CAl2ReKjDPDubrcCAQCIDu7x6QXu9vKqz+Q/XNf4Tqv3PP0uuhDDXRPrASb1r
svDZmUOiPVP9XJQMIAfBQAYhaiMDS0kSeH4q8N+v+RYwS2Dc5hsvbhsl9Yim1HlG
2Ax2LDE9yZF3x4+UGd7dhSQvG5uMNy1YjTIiRYdzpKfXL2JmFkt3sPi+YIepor5+
Tb/+5IJKwyFUJrZll4GzY626KxYt2JqbyHwBrbQ2dNp4uwWE51HqIlDSIGcyJ1Rv
9u/L57YnvExYse34o3zQSZkgMWBNzz2syCNzY1mJlhbJLp/XIGW0b0HNEQBAhGOH
lgsHweSwe9q6uuQHVILNElJEpkQw9KuQA+eSl5a/gTOYQvUmHZQSSJAk9LRrHRqI
vZWezQIQlERkHFGLfZK9llJmBGZGxfRmXrvY7WXagep4+t+4uJLfyhk6s+1fcG8f
WWOdvfXlYDRDwXd3U24ZXZzsBBPlFj9GguPj8VCNF5/o5GjSqHqcn+CIc0UF2Ko/
mls0qbKWpUB0WqEDdfDW2VId400W7HqAqPXcMk771+V5hHkZYPKeQC6pu45xx+Xx
EwJvoAX5NfZZXQ1vkl8P05NGwecSGNCI40qnYKru4+ItU4wqbTz1LpmmA2BHjEDg
KAtvMNe6rmWvS8/HxXihFLtsg0EWgvukY4cuLcFtJ3mBdKWDafuhqtdBTTHUUFxA
WSyP/8lxK8+KqvVaZx26jyFXfF5F3pJsMJMtRnvBnuNroj4Vi2SFGvnaf1zKZx7c
vuu15eqBbCCUVw8mv6WzRgc/oQygszgTR0isWmjEUSbQR1Wjnp4CdN4BhlskBi72
qUz99X9Hebl7uDZO88uqGKopPNUuIE9ewNmAoGQjXMpw+x8KQG0T8wsV96wGV/W1
YhYfzr7rnh+gAhwOoFWYRi8ioQRzlMpf2mB9nYo2XO5SVfNktHXftZSgKKV3mLnK
JkScI6vYXcQ64h+jS7hnPJ/tlG2l13a5lWFv9C9EVJ2fBhxXMEhhXHdg3iH8Ltjn
IfR7blAS0h/jqeVXVzool3XsWqVg5finlDeB7uAY+Tty++IJuJH8+WzYrTsx9pfn
iHyueddfRgOVynCGJJ1vySEo0a6v/epAyV6iXlls3n+0aOIW7soeZbI/TkE2jfp7
tQazpQxzhMvr5sbRSrn9GfWrA9NW4dX8gvNBXCI1q98GbHGrQZ6T1/yCpHFGm4Id
fp2lWGw42pKg2sNvJa4gdKojtheFuuG7VUNiiu8cK6ljieZo8MebUD4XcQzvTL0y
CPFtNk0z46/QlmfAZSucLNda1ar/J0uUMJ0tcoBJ1hsy6LocCs+YcFoFgFZKuK1t
ZoTkMuO1D71JTBRfS3vJ7OeGWiKZOcQTAJH7xMi4xTrwi1asSB5GO1430lk0W2Oh
t+2LKnAKTuCscNVgS36eTfcnYMo/0fLrvchx5oSlBQFJMTZNzix9y/rByyg/L1sc
3neX/2MB0uwEm8Dle+wP7XlAJgI82UGpRp4Q8h6B3cMhnv7/BzqQNLJcDko633Es
HkGHY6Zh4lWIyZCDrDeT2ulFQRzkd71NuAp/iS+K2+XPgsgSI/EoiAesWBeYZFhC
Ytz5GGzlIS4iNuX7NioOL/pkhk6xyfXbOPVKjLxoIVFCeuJuaFoKGALnJd5bx1A6
NdlFElDSNvR+t9FqgzFLR26+a4L5onKYNSelyuhS6wgFFhnKWKonNJOaxa1LZVwF
R9fMQvwYC7453cQZ4QtteAPF2K1e9cd3VzidkTtMdBwE46LfMaN1YMkr/n960M+d
utV6GBV4z2NwDQhs0dJIt+5MBSmTXDW2Ed3VwmQjsi66KU3tZAiLyUlDPX9VdMKO
pAtCLudxMa54GDV8K6Sh2uq762duM7bRZ858uhIDAtztNBrbe6U2Q3gn6u3+kS9h
E8P2pneZzLD03fS0VOAnmCFBMZlHF2pCP90KTYrdF/qkFW5IwTX05WupxtLuB8e2
OkXbICDbSyzLPVLb64S/Pcehl2R01V9911/Mj86xM7TS5QhOx7U2ZYjgkPgPeeHV
+aw5D30e5DOCDrARrpJ1mO2iAmi2ZvMUWLK6v9UXoY0mKg0xdXd3VJ0YNHKPB+id
kSV4rfkJDTAvulBjm/k9Mx0hYowPdrxiACdJW+2qyYN7/71rRSEgZwDzFg2Fh5xm
a16IntlNsDr747DZrz6qs9gWSDPsd1Q9b6aaclFVc34anVf5GAlxv1kuvbtJspUq
4PCMTUlpu+Lprsrn+UPmk3DDUujTr4xZErzCUv4OUEZIMMKouuEDUBDl24YlkOsX
vNfwSWmvWA4WBXZbkZWorKLM/53Hcu9QqaiBMxVAyWp53Rs5HboWQr3CRF/vcqQF
zup5vqMuUwV97Qr0wV5p2agNuIabggPDzheXpH0bTDJBmqQmquYD3tZQZQACn7DC
TVAz7Am7xOFoqWGwEehjBhzPPXKfd/oNN5m52x3I1+PwAU7d5SJZE7xcdg4c3B57
h9K5VQtx4D/QW2RuvlP5wYihYPnmFpKCnMwhvjEWYdt4R7EmJPvmOdC3pAaqpsq0
M8s1BKRrUNYTujWIDgEtZtdFuUhyWo/D7PeT44oSmoL0vF51WPfJr+HrtQDaTs/Z
hjbDEjcPDKpvfHPuuTQmiQsmyWIf432ZwU9gJz8k/4Rg2zKgAAGWpsOmOFDgf1pL
TmO8uB9VChT+nf0iTZAr7H+OoGdB+w+hb0/pOIE5kiJvcHBuOE9m8Fdx0nk3tZGv
A6Kb5ogQ0UiU+vrkH1zxaj7Gi0WmY9YOecGL+ZqagI27LgvY+TZdbwb6DaYanRCy
7jvX6gWtDAI73V5Q0zlDUugMjq0KGXbsqUI0q7PzjaAUeiO0z2WKYT4Jc/fheDc6
pTh9HL/iYKaCjUhZuBWNoSTIUF0lDL6WCW4M7/ATRvPHsu6z49axrm0n4WaTH/N5
6uIOOidJmgnJuR/nI073sEWog+C+d4KGsp8KevNr8TTgEmd79lcniQBAlSeNRsZ7
FPZrVL35ld/4TBKmP5KbG9ES3WdIIESbaYKFcSvoSdP06Lg1Iya9ujxG2k/PAHA6
hwYSEpHNEZbedQAIpPgD8x2GU6tHTtDT5n1i8Rsej1BbiA3XgTR1WFuHUQJ40Jvp
5xdrKeNEAKdxVAeZXoXle15v2QKXYXEIBhX4vVmTfcy10Z6k8od+iqCt1zAlLsly
sLh4SMfc0dIJgm0QEWNifowM7R+i5fZtfrzrobvvMk5FlD1RpGlfC5S3nTDip5kY
zrNgrwgPIndKlv2wBvSpBtWJwZlv2PxdC2KU42elPZlQOxj3ig7o8LETWaZs/lsu
ffpaqZw6pNkwsZHTc0bexkZDI7lxKPILTp8oJNdBiJrMjWxuDB3Nv0qv2OB5QG4c
Qfjp/AdltgSl9fkTH++JBTgNRMKd/tTeo67AfcqWJjbwJAwI/vlk9oN4GLfZzid/
a74Y/rjPLxD1IXWrauteOCzFfwCeaBNhagDRkY+79E68sP7X/9NUvR3VPZvvfC+c
fyLnmpiEnSUMfJSite3DwOy3DRibltLG9fWQpeu9xGDTPFdPdhaGcx70wamSZ+wj
Id2yMRQea+utMsOhr6GBC7RB8rDD2JDYBIz2fQA/5pAgIs/eyVTgPZ4Z7o97TcfC
s6ieNE+97vFY0eglSFtI6Z1yCtsurlxmGnd8pxpFMD/4YZX7WVJY+bsfitlW+LuA
2Xn23dlAf0lbOOUmTVNr5JJoJ81fT0Aa4f8E2bFF7aIPSkNyueyXOCqHaF4Rcc5q
hxehhtESceaLbDEiadKP4ynNWrWrpVKE+59GP5fLhLK90z91+dNfUxwGgS3yVg/B
DmJ8noxDkr7s/lxsL8AM2y7SqgXY0y195TknHGeVqoCQPyTPZgnuHmR20tCv41ox
/e8JjsHq47kWtJ0sjQBkm0K9qGhZCNUlmjMZj4glf9H5PGtRW+/4pQV83OwWjyhs
C+tF9y/f1+YG98VX+X09EdiljRA8PX8ymj3q/yR5LaxKLImUpFhhQ5OZKZ4l/edA
fnGgPNaZuBx1kn0VQi37KczP5RFQwC3aShKzp8UCsLxtvc1xAEvAJM3Yh3KZ0POI
xEAOgOtbJ77Lp9Kbb4a9Phs2eSv9Rf+65w8JVspvcWhGavoJLMypDGqE4ahy2Wmv
f6wrXCiFb3hSyDpY/yeQJWl2fo8i3B4+1rjvsWckEhC5tk3KnSpXJdUfCVP7Hv+Z
dxwXiKuLGq+Sj1qK4lbIVvgSknqnAUlf0BS0qPsupieoW1dkBp69TyxYpBTA0GwJ
2EXrQxln4Wb6JfOBuKzQ65qOw5fqmbv1Gq0lxKefuVeZmCcajQmrpS8F8HIYrWHG
T+XKqPQNFzJ4vjsmQirJ1oVs4k9ColOSCsNw7+Q8c/annchJ7nxnt9M8jBAI0Ace
XqfPpRfshYdKwtGehRoaJ1bcfXoslQH/YgbJ642E20g2Ct1a+Ry+8RI0buKxz/Me
YZtfkvwRPxWvuugz4b+TZkmCn/tP8JrX+fVfSl3gwpTbli0tdGfVFSHlBi+m8fFc
Ik2t5GRBZvqJwbx2w40Ly3d/yCxZCbRVBhreGISHO0jgMIAK4W2Ho0FhheovX0xP
HYiF1S7E/dNjNOYKoCUnvoe1i6CY0SkqjCFG+xfFL67OCYeqxyXKt4qPudEEUYoz
hCDsC5cG0imXark+fYmhJSWZCDczEDrUgHWWm5C1I7P1TpoKS57bZ0Arbk1B/kqk
/at3LjxZ7Y+lZJyMdlhlw4LC+UakvtMD4jGF1aAYl5i01WxUQ0uF0WxvXtwM6j9/
zFc9u3YCWqkuFglL6lPEqJDEVOiu4Vs2RLHmuU4YcrvATCDC6cAEGtmSYXkrb050
OJ32foqM4ms8CKV3/hJNQCV5D4NqhmCU1IwC0G4VilVWfuCY6bPpBsmu1qOG+MAK
vCWodbX2gpQoUziF4vccofnDQVzm6jMFZSmbIu70g4bSyvZ6C9+iuc4Crihy23ah
aVJa2eGv8A6BVGaat91DYx8s32gXEAIZ9JpT2aIZrH+BNZxgg72o09+BfYF9zn45
f3Y6KBhOAdEP4o20Rv199fZ/AKZo2xQjSIpkTRSUpRxQ9q7zdT7taFv5or2rBsJx
zm7uxlmz+J0qnOiUKUacER2ndguIb2pY5PReRFDGZNa6zL104kmORoNL/oX4BDfk
KKyh02BxlPe/1RzSewYoCTvwgHTPERX9PafyoaURtgumwUsRVONlRdNoQcisGs8M
TWZSHSH/KJh/8SUPz/v8VAdxPhWr2ddnflAhcQMNpbWcZNCsswxLv4B80Hewf/cv
xWfL+bXE2BvF5i/amNfC6QGTKFBRfXakXP+olHnkRGaSTxwW4fJTbGk/Y1uFQEMj
6nkfiSahKVk1iikZ/lQmT/gGqwCexJOUWBeCbrkDYPVlyMbzNjMxIWy1/SEBo6Jn
AIku85tSadaNkiP22eTiMi1KhyQD3ZIb0r91xr+hLvbMiJlJnl6R5OXDhf4dkZiX
L6QyDARfjcKYZffFNtmGnSIuUvqWwwqB7jzDecPyEBchtMJYIxTLTLaEqdofLrp1
ncUcVMNQ+36uSSQCDRpsHLnInwuOlAu6esSOUWUN5FR0yEWUy3tHPcsEd9dT5fF0
72ljpT+Squ3EZ3ix8m76ncaE+j51nHSRboL3rbZ8tPct1wMuPTqwarWlMOcDDMJw
X93sxbS8yTUbMm1ZQnw8csKUTiyAH8IOjzfsYE6cy7TJoi6IRMS06VsSrvPPPCGl
+WaYRIpdeRFGmCj+ru4taX6yjQyu3CdSCo89ZP2VKfSlDfoxmyr3YrI/CcwcxSMu
en36eZj1hwxp6yIS/CybP4rBk7xA5BdnLxIzdTBq/ej8rRaMQ2n/nWKBBsViaRBC
rNQHrm4mIluZIOqg6Ts4Dt8WPjBFRdxF+n2t+GORcdFGQLfwzSWmvx9VdHQB4bT+
JsyilkFEnFA7RO95ilwmwSNH6z/WE9W4fV55QS13HNHiK9750kX/xmKbLQKe06Pb
L+cmIWFQXLa511zIqzKeHST/FaHv+NKlclZ2z104G0s8yI76ScEuuefpFTP9mLCu
x5CVe7XHNYeKZ3VEe7Amt+oWghpnCBTBd532GdhEklvrf3wiSKXEh0hks9YOBd/G
qpBVvfYFP8ByhoWlPQvBviqmw04hyXBya0Z42QcOMgnAC8corPNEhbxJyIAsV55C
M0joAUWCIKQDfv8q5slKewXpMKLWy864Wfv/dt52y8AUSJJqi8ajKomqZ80Rrt2k
4zxrtDHYvK3QLrqEK6KHxx2lir8bpgYyjLTLuSNLvpCut5RvNZA+WqHFvsfF5ek6
EzsMD9bGvXDVuBnKDeePaI7JVAycF0+Eq1YancBD6kBqGP9u9YNXVdeE6x0HEWui
Rw5qjrd5sg4xOOwvu6kMaerfob2SxoNljG2bgyYhrjyvTWtoqEz1BZa2TDkxrmDz
iT9T6o29m6BNZmh/HpZ3lpLdVDHi5dgvA4obhiDONzh6JII4Or2tEs/u54it0Ebh
e2P3NAXHmcsD09wILLkX+bZTXHXgTfTWtXOYtI3NudCqKHR1+mQdGo2Gla4CVAen
gXOXuOTxCxfwpy+sQZoyWlAmg4QvNmU8wfwW7WIVOWV/fKMAjd5oKaIKuvuUVB18
20nO8LGWbGCtEvx7BYBFnaxy61CjN81Q5T0ICxCBqwKqQA3RgUWZlSLLT4PEPCVE
ZwNiwgGVPuO3nawlfSih2yFTRK71t8l9hC+R5ciyOS/lBute42XZkryGjdoEqSN8
+QvHxZ9wbQ4VEUFKw2Pe08lkH17Vzz6dVqntuov7N8b2YxQnaiPbwtUWc7dOslMd
9yAAnV11wIILAaEmbN3npUM6h0C2UgqkO6Q01ph/zW6eVeOsF0uLchO1suLweb6t
VCqXaxu6y3sCncgaibYCpibtwZTF5TlmNgd9tgv4hZyL4r2Sy6VQnYXZyqv9XYPG
BeXpEV/dNUEVtocHRATS7/M+ofmv/UurfCF6sjpzpAwSWtp3+RvGSaH7By1o2tWu
BzciM5f3Fx7SIeEK12RAzJ750I9fEi1vUtJuCAZbdROp3J0KfSBYXfWgnKBvSwiP
9L02u6Na0TyivMTq0VdQOituOU95Eh41tb8NOLHX22yHC18pPXDbOrKBx70wpGzE
Kb09zYVMikPF41MVafXSOYRe5pXwUo/FgwcaiJxWzIBc1LlmzIXRbfzlomCxDCF9
+kTWgNkYWggbamCQUvcYXyvSSdTdTclrVP73/PYyOMKkr9uF1dKSiIObzjqunsla
BUdpEBHWmGMYXPfxyOAIKOJRQXNRo3TH67k8Tn3d/FYlizPiLOH9szyibH7iSdTV
G9OnqoiBYPgenldxQ+9r6t4gw80xJlOw7tCaTrvDGGQtItG7gzKlfnHdMTwXStC/
bo4hnlxmC8gbrRubtPaviIbYzjYlbwBACesKZlZNsVPakEBoTlVFLXoLiMJceaCE
P6bwFrUUw0T2y/vfeXCsVnm01D2uWJrAHqSYlxN/j8XUgU8tDZaLH6oqwEuEPxly
xFs3o/hBVwyC8z75a4STo6HCnQe2Y7+tvm8Q9phqGMKQ6TLnfpOo/ixd6Zgz1HkO
fx9ka9F1ocxk0VOZlE/81KPvrnCjg07hpSHkpP5I39qa4EK3RMyvfvNFD26Tv/uy
nSJ1Km8wx2Wt5qx2UqyMJY/dO/R5jFRzCieMtJ7UymKJulyVKIQkgXuuIF9CG0bK
z5SLgfhY6r9nmANqokxzwQFvIHFX6r+/N7seBrWh8uV0yph6YsAWpYQ3e2mmtNge
KtG5rgE+kFWzkw970Nkw9wTmfZsc0b9o+2tHYx2nAkcYf+8LsFjdrHKVQsl+Rr4f
Urx8DkvwG69mQ6wETQAqKamtmOHilZJbZPPRU1K+V1A2riFNlGr5x3tgUPOTCf6s
HDAuc3dXVrw9OWOOVkPbAUsyXy39zIjFJHyA60hjbegMDMMaucZzJEEsRGohdBvK
rpR6ofNp57smU/qBTNC6XEQHMrPCjIvZmG6vnNgcyyz+Eof5pnCQDcMvK3PHP2GU
wzON4RmTBbflJN+p4pCqc5J5ZMiw4G+q9lDRZjifdOFNAU/c4ysSZo433jqDEqGg
AQ2cFzJ1KotNjbXAK/WVspXGAIi6mEXzEKOHPVab43BqTYWkO9vi4SJwnJzJzE8H
hl7+yLTPLb9djt86zKdoZgdbKLCVuC7cN7tts878NCY7wnN6cl1C2Bn4Pw0ng+pf
9uBByDJFO0kCPUwR61M7hksEevzEaZhVHx0ICU3dwTCj8oOT8Y2sVJJve7YkKdAq
7Tx8Q5lBAQz+tSBC3rMWiNU1KKMS872aC0Q6pP1hab2UnyuFwAO5e+oMWGnzJZXV
dk5ri9guxegShJQQFTPkRKMHmMYYrvL/rBV7ewGovB4U9K7ANJWJOGh2cwZiRtNg
jCsX5vkELRDpOXpJf8MGSJWILKxGyHd/SlGyS+ktbU2l9JL1zm8JGKD7eHORekyy
G9Cz+NuzQyQNg7BqE89SI0vnZhsPpg9/GsrYMuD2AAONNObQFhKkiXtO8FGYMXaC
qZB5jlrMp4SN58kJe9fy3OsMDHzpGp85NG2qetwJ0yGAxgC6ymFZdFL+bz5XzmGk
+AC6/FPazCXdoD+QrqUiD6Y5gxxVuyP9hjHlwCDQ+hrzkQ4N3r60SpJMGXZt8MWR
1/udP88R7KSKmsVADsNNqThNu3/e2+UqxcUl1LBj2+Vcs8c49h41BJxM9zXprpBm
Iw36saos8vJ4qp17PC0EUoTOWZotNdhzT7m7PbzQobMg16j7hctyzv76MuvHCDHK
2ZMokaQzhGASaRy3u9x3E0LvhCr2Vpub/02M9VdGZO4qT0UyWoOTwPO5uWLvjImX
94dcx+WmlIUhoKRMu9S37hK/RqH1UFPhRBK4a23ng+aPdGkHn9YcIFV1Rf1yMSZb
PlktsKeujngbJx00+A5R9j/D7NZggwmMjmYD6fy5XdzPNF87+ZEXblUUl2y0ox3q
tyOHnN4ahQbL+mtCF2cVcAMMRYPP9JvM4KjkJa2dLQgfRJBziad2JzGbjHtP+fFI
qmono70eETwdRRPwF5Arvg6Tj5b5T5DjsckUEKJZgdF88gdxUE1o3RB1QMuXHlp1
47eMGIDahqkJbygyYQCzA33suTfI053mYujhsiH/KLEqy3xRRkH3lCcLJwN4kLw1
noop6LhSSu7FEJsMBKSXKo8XeJhKqVXzK8d0QRTklBoW+9+oP3j8qPiVyhd5wKs0
kQH7UkqI1k7eAzQogolWLU+0GFMMOk8wpTKv5Inc4Dqs1zKfl7d67RN0R1F5mNdr
kAeQ1atGSG4kghCd+MUBu9OwzJbQtc6J46QjlMis1bK1WgCWW1s9o0TvG865Wz0T
sCMN43Io6C0bV5wKx3+V2+0rLoYGJYU1aoYvMdZAIsBhFz+Y0TOpYxuNVYCxFyKc
5PTM1IGgLytqm1PLahtz1Edela/jRX+uc8ioZyvMo9qzXWQQ1O+7ot16bQbYF5kj
HT6GRO3fyiNVWF6McIpYX1AlYVWN79YIrZ3/4E8pqVkK5sQQmGEHeFonmk/aBcRV
sdbkBMqb7vn0zTdO3VsyMPpwKdB7NUNObe1ydKtTlFq6itJP9l173JyNKhNHn74/
KI2oQYkz+HskxExHZ4wwuBu2reyO60rcxj8ZIU2cseDbbJMtlEW394bYQ28uan1Z
GIN+rr83tk/r/dm79O2mxthl5MIO5ewVs+aTJHQpOxMFw/FbZ+KnrLWhXH45XhzP
MqxUmbwelSsdcZ6lsGgdra9G3pUsmfzxLOcURoFi+osJTbnn+kxPmPMcz915wjEw
/6RIaBqocZPXt1KMOpVihYiJGbroqrFAA04I/vrXl3utr8gof/51xJR9hQBF4sO/
pwF6mdE8DnTijdoEYusqmP21gxoBAwRAKTnoNCk5tST9jJEmREty2ks078RiawVY
Lm6TUFdnqsWlRtf6RnGAYvmMim6HkZSjXj2TC3tuj/H5fDh+6yPUWTKghN+fofa4
kMPIs/TIVtxuZIPf1SlNrkAGxSl/jjPCKx8xtdTpVdzGABWkFvuBXVTxHdZGiZpH
4oJfpw9omKhpEnct7iLF7o30RA/J2AXo6gYBB5AtyxdzrO9FCFSNLmOTb5JII2QB
voG+0glNvGu8IbKyXDiAZjNfN7Yb2AVeyJ3GtQoCrrn9Ve0KHWg+r0/DwWgWhlh+
hxJo+sQWU0rZW5X9qbGu/47gtW4nfe0hgI/f5J//FhdnC86s1WCQ+RJLP4lYr/Z9
WKHwzUKE4+caf4ploEYSuc+sWdpGSLe/tI6jcTxul8BsEtlWjCdWIJIvTlQDo9XU
bVvBZV/uugAkQC8rb2aAQTQQLcn1WYUvYhd7bBaSmQ1WJ7+ATCETLSxGvpocBvHz
Iwc1H11l2Gg3pEV2KhQRZcl6qjtr2vWtNfi07Jj9Jwx5t7aWsYZPzcFr5sjYBri6
MxkM+FpTxcCtPwF4IYeabCCPXHEsRrLm9UYYOE7+e+MEd1Z1atgz/h9AznQOe/YV
I+95ntWxsvArJxAYWx5F6G/ObVh5i+wan107kUbyu8EM08EXJW4Iiy6JAkyELAQ+
7qeL+DcfvgMu9h22sQoyzoBWhxbDjGWb/SMoIvcjOgJCdyf9HgM5zoGGJzrVc6OX
dV0LBFYYZp99NQZjVNluAghsaPCp8nyemR/r07wgdG4VZyeUK5ZmH6il+9f7Eakc
MOQWqwTB6k4zMlSMHiQd2k4dYqUp3oPHp/PuwbKmfv5UsbmJMI/39YQ8NuItiSi4
LcZf+a094iLN/uV6MkP03IJVFPu/ZfoEvp8YvKnN4Bp8Op3YSZA2QYOy73s6VRA5
2PzsBqEz6M2dKolduRQRWG/I7bjvhTWmMeoHnElgi+TeRPhA7i7GuqgjL79cqJDE
Wu4lsPMgYGr5RPgHcBbIZqtBVbt0r+N3sCovcULd3TjPAD01yPzNvl9diBgzG8gd
W3716QKPZysd7x2ovYh704ykGdCDYmQTOgYY6iFkDyOUQIj83GLExxFghZAIJVGM
73o1qzzsLc6AG+t+ENXoWpjOXV5Vfl+9lbA+u1NlGJG4pX7+3IMgEmWBhVU2ws8V
vEZ1JiS7FlYOo5FaN3wcTDQhsPUia0FwQ13ckFoZc7nz87g76rDRBRiK/pSpIjwL
qVdWpKD58TVRxblXOSZaLLFGdZxeoiyvZTnS7TVBGK+b8xUZetFfPAXUm2dsCq97
Jprz1bHy3/aYJjqD/SjH4GoQPrjfHk4TZFX8bP4l0PjU91bJVG3s/KYIqoFCIBo0
RrEaTlCeqEiUt0dAfIUAygJVXENoxjeBQ2B5aZu/F265NJAYRD6IGJXmj/u8qdYP
/y29b0+79pTGOA5iGkhpTWDfYTizqpK38c+L4sVXh8SIobV+3LwJbzDg/K7nOjIi
dHPCMARzsX+vvN7hK2FmmCMKNZ2pmxRYj8QjfeMJw5P4V5YOVSGg0ryy04dkREI4
rtP8+5S3qdMO/aY4BBx9Veo4mg6B1q0QX+Vmfxcju9AHMszYuDcZ8lsH1sCGsTnW
1tRW3wrE0a3/gY44gej3MNCx4pH8AJU0ZAMU53DyX971fsB+/rQ0OTaylpEvoWWX
NGW8ztKYDs2yiDIpDjs22kC3BKd1IdsxOncW98EwidPLJHg0f1AfDNRo9l4nrW3o
ISinMON6qU/+xm0cYtcWhLT7l4SiEXP8Rbc2PFYe6GiGZhnDTuNlajmbihpvY+IP
+qtbMABy2ZZxa/ecLAhFWERabn9Jk9y+hRiN7PPRTLvdgJB64MlXyqHL79p9Trwj
8uJhtHrlI0njw4m5MVTpN1ZXtGcLRayr32pPydoiCeR3lMzMMnudaR7f/qcefkZN
PdoKO5qPWX64euM/OUItuFoGi/1G06bf81zdtMgdQesFpWpAsJKuOb+VREBbOgaB
CMAGcnlz2suOpPJy9jLEVN5OhXIdp/g/VabZa3Pi+Y2H1iFNvTLHeLgAJwtyCgmv
SpoFM6WHlJSMSuEuTuJCC5M0RS7yGubQ4rM/TVcId8sCYb7B9QIsugKkUPB9SQQS
RKSZvikdW+BxGh/kGYUB82HJFZD6Xz0Ruit3swxobbCUkplY6Oe8WWDFIXogbz28
o2FaT4KvBmVS7mEOCTTdaQvxYZYqQe6EeR9rzXchRK+cj67ZMQ7U5AJUq5DGY1cA
1Dqq2yRC8zkiz1aQW2NsOdXvinhw2RLg+9oJgZunB/1t/xer2xhnJgbBHMjistTt
1E5MUo9xmmswa5niNETY4JJViYTJ89zhpD/+aO85fTlSRHJ8W0ffZEgdkUr91Jle
qAHxpDQbZELGFcPTjiMHewCJCEhsVxkKX4O2physPbtJAok9jlF6ym4ZCiQyaf+W
d2QYsrZZOWRbuwRGaTCV6WGZ1AifNu5LcIWLAzuETu4juzuIjFH9qzOJ6OiNH+6I
/X79X5OXYwr7/XlONcXGZFOOV0a1gCuiRqsmxzgIrQ5c1YIqg7DxQX/GxXGaSqv5
dVkefHQ97qt/7/uJH9m02Xzhk9X8Jh4hqmUVzXk819h3YW4RG+gltDffAiSOjJpX
UEtVJyBJ90hpr+CISptQVTLEnc/C+PwZkUynr5efmJ+uBB6t10WvYigM+/tNXKED
+u1ceFMS7aSFbDRSr2S05QCynWW2E4rx175NheWeS9UHy0teMXWTKyDO8D+64xxS
BA+ozJEbAEmnkzjR9SowxCSWbkKvb0Uczo/s46emGsgOQ38XD+izIXyBwNqGoo2E
8espSW6+aNj3x1CD+3QJv8mpd1AI/dxuPxeLlaVBnGkE154e33LCdfjrjj0Ha66x
ftm8uvi55Bb2GlKzfLii1KgbfG1ZewMObfkktlk48g6sdHjObf6b0Dj5Y/Z7GeyC
ypndu73BpTI3W5FGRTsiXr3qn9cIOxi/EZyoGzSUoaRYIfhbZAJDhESWo9K2/b/o
T2X2wMQ2h0TacHEv/yhlu4aswyXtMvTq7jfbW/1EAFkFjb1aRM9WLLkKWd6DHm0X
z0Rqi+0C1LE+Jm/oXvzAp3m3qN99+LD5NBghsVslTslm/VDRAWTAD0vIDD6Y0z0V
HMC1jt+ozBCod1tWyvmnpoeAoS6Zzbzb0Z+T2pRA2I5xG7kI7N+Z4/dmENCoNOtD
rwNlqt3B3br6VhAn2MdDjXDwxyxpJn81cBq+Ox3XEUI44DvhMjpbo9C7xVLsvDFP
AfKVWfZZHGz+u1eQ5fTOfWJorvAjPbUwgJULFPneAj2UruP5bZcjyjKF6x4lxGR1
m3ggAx8JpyibDPJ3u8f3Rb+4vFkkU76h7Rn1WLnKrq9fCNNVedtRKJjKeUFDIYZb
WL+SOeL5b64v/mhopy7NsN7d5NoNJKb3V/nbqwQisJey9D/JcwX7cxHEOG0jx32Y
u101w9x3hkmHsszgiwocA8gG9t72vmqzzsKTMANxq2KKaLcpiLDEtSWIx8SgcDHR
QHvN56tDYv7Y4W5koL/2osTQ4uUlHJ+ECuTP+dMa93TVJUZRGJL8Xc9PY0B2jOiv
PyhGxcr5yz+LDiIvA5ZV8VQVEvLPowVvf8/83MgwPbEnx3DtnOt9r58tFIYuzjTC
2Hs038UK55PtvOUdF2xTsQuToE1DIa6GYMkR9V9WaVa6BF60oi258zwBS6/gOYq8
ckQl15QEv2AaXGFQXuNF2T3UXVnDubYFKnGCEFcx6s6jpIIVKx7MAT5vCzbgysAo
L5gREpDD3p58tM7wZbe9/Hmm9PjMK7BKqBYlZ5aKQHZxkpj2BL6TJXtXl5s2Wy2b
sTTSHq/qx4cV2wqjs4ZUGobz3TrPKc/YapyWd/NS0Bx9vwQy87oqWAj2T9RZEZAU
k5Jz+g2bD4pGbTDt9m5H7UMn9iyYs45BVbVvmz8ewSyz4p2HhNlC7uYyLuov515t
MvA1HM978zNpInLrDQGpabg1CD3mTBf0HOua3y9apB0hCtogwAW8mvH1yYWZ+Evp
VPjEXr0jn+KeB7SCMxLdK/OyhoPhVJdp7IBZQpYdjxV+Q4Q/5NmiYf5KtYMNcf2T
/WseiSnGTe6oIuACMEjWTGSSYIRehuBMgwyue1sOUFp9t4LvCM5HK25FvuYLtnwd
9aTqpt7mHEzk9aAhpkOsKeS7A71ZdceMdH7JwIqqSggTB3qCq69waHvtk8fFsZHy
bsPFZXk65lFhrAQi17HKuy4RVgKZKoUz2e+i0bspcqyf3l6cJLVNyG3aL6JB8O+/
0JqaQxAHfso2u8iv1/BYpW4Pad7nnDQURGNM1qCVNv+Gkq8VAX2JuAm0rBZcuXMP
/T+9tUbeSPrWQLSz/ooGPG16MJWKxr8Ot4pIfjgDF+Wd5nqAhs2G7eDoZlPmZ3KV
iZ0NF/rEa35JfKnyGAKeGFNyU4a6Kzofg59xeZgGUb18inG62GEiYg2ZJayAdWno
XaTW4L+dSZNNSfX0uWwXB6DSJ23G3V2UKjYIVj8s38CbLJhISW28Lv59YcdyT0mJ
wMUEtNGltcr3WJrM9N8rnid4E+2B3qw4bLwd+DRjNoIv1bMYh1mPDJfXy/I8li8P
trcRyUsxg3RfJFsRTtHQNMIlvmJJ7LymTGQtH6HhsO7saRnwT36rJkciuf8YsqhE
QnV/puVjqLbzoVF+VPWvVUHSsP57ASXUMmg0XZFN8NtDK/MlixpIRD+MN9EkuLHK
G4krQ5SpId8j1grSrb+8m9ncju7fk1oawKEYj66hd9T1vhqOfKEEYUXsdTxMigqo
NK8z39yc4pGPDNP407PDUf4020FJ8/v7Gu6GxATIhxNVwlsIUxaevR4nkY49SN+P
LBjBdccpd/NvAjSr0Itoapg375az19RPJH2kf6sADhJq20tGT03ucKX01cqYPdJI
Dnit27HLLecB/78xCjhsYQ9U5Ofmj2X8bRZ5tqJhBFNdFGt/BE57XoyTM2hsaNJp
KmXnVEeXZIMNX07RuRsgL1C5vgKK1VdK4egW4Gbd1sOuQriCTQ5Sq/QXu0QM3xi3
+i3BlUHL9+4W67HRagCO6XSchkgPm72Qa83IvO0q60azlwOnjRl1humcX1TQiTnY
QcY+vT9aF3lxAxyni7pZgerai+Zfu2dC4/Zu4dSS6fwtHzImtcwWu4ym6IymNtKu
BDG1KDEPVgmvi63XoKc3bKn34eZp/VdPBWKMKddk9j72KA05dsYWA34oH5Z4dU0y
Q3ayqj2ofIDwZIK3xtggIk/T5PyzvARKxVHCZbyKarzJP/OFV6epaCLqaLv7c+4t
PW5D/GdbBmVfP/weCq4udrMrxEJYjVCPhftfLi5LvEp9sNYz5O4oZp8cFSkkj/0j
mSGPJU0pbop07RsxYC+YXFqdw0RjLgAwENxhx1vsHe7XeJ3JMXxT4zhRy1O8DZ3N
PACvcwqFT5rpCU1ekRnrZrE631WmEqO7sxi79DbmqWA1L4IWHkn78EVhDPUj7HZa
br/N3hgn6i1BCj7ZRRDeOSz8R5kJ4WIQCM1yy/rXRFpz5YV9X7oksVuu1IC6+PJs
NK1HMiJKdxVlIF1zjAyB5kWKlsF8heW7JgbwomL4ykeoqH4gAA+kxT1nHRos61DX
ivfRJtZp91w+q8BK7D4FYC26AGoen2qz5TTX+D0DGZITwt1CXv7hpuiIN3TM0330
P0mjq0OVOvEZ7+KzGRy44MAcOUDsQqFvtIGwG5cF0ljYRvRmIq/tphmApwWViAlX
h5lW11mT0PO80Z6jQ/sw5up5cXUJBIMEyma6cLCZR3W0g52NKnH6Pfd40lBp56pt
yQRpEPQgHdPhmUnCXzb6dGXWFCaKvnUM9eJYkbGTc+01wm+UrDLdwMYmNJSPHqFr
mwoptVeSdMf0EfHG+mgQpsGCI9nvZpsHxt5TrWYXkn9KdQOCmN+NV5OlidntaIRR
a2vb4LJNJvjp5jI80lLqtmK+CaDhqwSozLHh1k9Po0KQOacDPtJteh82gHwveNLr
B7tDO91DhKdV8qrJjvSOlcRoPG8iubN8F5Sx9Q10Bfz8cjBcrhOARKAOd2YgD65Z
sVivRks1onTT1Wsi5pCTyJ0I7Ll0Mz+MeR9yFBiW3ccTbrdqu3Y4i9h3d3VUfdik
GLH1s7FGbakzIe8ZF7+4q0lxUr3KO4K1ODKH1HcBsQGZ/u+QBD7lfEAaFKQoVO5I
SKZ5sLdqsgJyABsmtKgFFo5hQhf+ibgexhEgfY4Lfkq0nWMwTh6aZe+om51rYLQ7
vb9KwWG3cfpunioKnT4KU03zcf1eghHmw6+wxutuHD+F5WEHq7U2wSFHb6vvfg1q
TpOSBBXdQUC2/9R2zY7wpkTAaqhe2XynDjf1p4ywXAFIziOmtiHnWKNWXOrWZjV3
Xo/1HGth2nbyd5Eij/xJNlNCcOoNZTPppuoU8EO8TWw0//0No6k9czEd1xMELDui
I0iilRg+rg4MRbwYoFHUwgKy/MWbwRodoz1WmfvMOQYRAUtxOca7eEqZPPPT/jsn
jpuN6cxDGl+fqdWQNCyu348/bJGdHEyv4of3Y4CStbKobo2D7jddzAoXx5ZiPR77
mJHMYnRHg6paoqCJSdVKZR7a25sDn7lsf6YfT6I579EDBbxKE6USHcUWsEs4U4sb
dyfIczZDcOvKuN4z4AwSywReQhp2JE6n5Q4rLr7jHG3xTEcJ4q5wNKoAA8qhBqQu
dJhicE3lv4vA0Q/hz8gnQ72gWAgc+Fkn9ogFhl/F/iOWwVpygkK/oJ+RGnCxtKKP
E5apv7xw5c/+bPWXF3sS7CMmR8fVCEhU88JI/6KFYq9Dx7558TbZvnP1mmSRr9Bl
aOnyPa73X8gLyKUgOypS0eS9kItFC1GCw0ISwhf80CKn/SYcsriM7g08vArk//PJ
wh4o3Gn15CmtxWiAuQkwx1O+fyeKh3XyRL63Dnfy2RCxf/SDwhXF2kYjcrz/YYkH
AH2yK2rB55em2isyxe2DK2b9qkjPqLB64SvzQ+O3u7sLBJCVrBJzpvh+c15d+D5b
FeRXYb6+wejFkIb2j+qAcxeedXueHmIuMgz+Pb4vRlLvZvLbqSKnX2TFS5hmTdqu
qmDwYy/KRc7SkX4XqDGdv9hm59R67z3AyqcGnSN81B9Qa8MKn7cXtRJVJdKJwUE2
58zyf5zM2gyhSNJI+OeRYvilgGjpLY0BiBtxsMnLxs3fYeCnrZ7wprxcZ2/FrFcm
RkkjLqetdomWxrmOoXyLUYQ5srpyK+iuyHIcxP1i0fQU8mi1bXTWx93oviU7ccZP
/Q8mO2HInHcEwLneDH7fWuxYziiAhj/L/NxbTRGKZ42iCHpJxa6eRAubk2Kli0On
gT8GPiGOmWJryijsiYPo+13x2EX7ffhPC2XQ+aIS1ErLgz48bdLm+o6XcX70G1OU
wB1FU0Oe+dbeJZ/EFK7VkdtQpIohC8onOxQJv+nLmcKw4y4uTP8M7xpVQoxaR/6Z
24zLcJlfCEDtm0rv/Hz2FvTKax4wZANEKAphlSmwK3X3UnkYUfIjPh7eKXO46yMB
WC3vWCxsoqR4zFHAVmwQR7BgE1ARIntqq+CUSC7dwZfO1pKvtiwOvlZKFE4WQXxf
tAVGbcMPo4ufus2o26f5agg/33HjRZcWp2giVplNdF22xWfM/22ciQX2mxstR5st
6oC7jds4eYZxwxg+2oGS0EAgBV6r38hmF0aHtxnReGDPS1KOXNhl3yEty1ePV8Ua
NfWFyCurOPMfJh/9iTTzPt0Mj7ONHmU20TpTP0ApQFPAePEk2JUC2sapkzFR5ByM
xBjh1qRMCFyHGcvU6yK8U2ZL1DlDM/5AwwwZQ7Ic2wUg7NH1broppea66zS2z97M
9Ax12XA4clyEa6r9U4MqVudoNPceBBgFuzoEebL7Oma/88M4ey+nFL6zfWhXjeqE
b5Heg5SiQWmHm7eLxj+cCxfI8Hxmt89WW0C4yv8mIX28xxdNsfumVqMCz+bDA3oF
zL8x6Jltvg4OULR0C8szp9JpgHD4C1/z7RDclKzwT59VDxAOp0vvCB2nOTnrjICC
LGoMw1MrLaB6foDhYbeXrPcx9pupUNdTJe5Cqb4Anu5ZwS/IFOAphnHdVNtxTBS/
cfFk/doFHSpgPiCmi9p3xdw0lDzn+JuVWhYzZ7Bzd0CzB3NWu++XTFelj4poceZj
Wd5VhQ+XeG1gjDIkI0qMraeILXQqgcb11Jy61JMMvEqj/XRKq7R+mWOLE4BMq/8p
nKMuTQ7RWrQDEDNoLrEF+gUygHXBCyyX5jPPEnl54SK2VEVPrKL6XMIqwgdPVz+3
kQhjvPIKalxwktYM2oTKjPBL2O6M37Dfcyru97A5SyKWcp9oQW012Eh2DlYEFC/R
Nyk1sqFZv9KqLjQEjDtbZrS1YagjWbHsTzpfNbk8bBW7tbFF9mwMWgtOCHy+hAhj
qoS3bD070hPDJVtqAfcAYejc2jqregmvwcuwyB+YxEikSbMlybFRHSsWScsinMFQ
vWJadz0f3F1p3MjHqlM5cuX+5V6cnJ2gTJTujys/of8iEeXg7B9GokUzywQc6w5Q
HcKL3J96bz5E8W29eSgCqyo1FzAisTCeWuDRxtpU+GohCFPW0VSUX1mGoeUuBC6w
5MzMwLD/r85X56eku79vBQWgm7fQ3yrENZhW/QcrMCZCbzbA5bOSh6ru7hqzif2v
Y1mxBVntWAn+Ko/LWg6619VWszOUTcVIR4vGQmYrl1iqD8wDdS93p1c7V3LXRBdQ
n7Ts/0iXSxMFpooSUjPLQmHB2sQ8SRynd2aWTEVIHZI8HNmWxuwU8ZVBXttQ6K2c
D+QbB3CRx60pbyesrNhXsjIsdsbp9emgGDd4mU0Y3smvAFAbPmfi0V8AhO2OWgel
wGDH7ag7IzzAtLBs1AiZV01WCnWNo2p64sqPx7M5Sqn9I2tCFIe7THQ7QwrOm0Gp
WOrYi2cnNWfl7AXj9Hf1vxyNsPicE1iohQZTyvG6/oRT//gHMk9qA8etpDF+vOt0
yl8b+vT3SEOvzCb5yLbDrqIDbA9P3wA4gcaQqK0KJU/95pKeBfCWRkIsrBIQqitv
oARfU/vb5yvDi1rpX69e/51lhFatQWYqMsdZLiroH+S2IH/aT5pWe7Sie+b6ccbV
kvWaCixxPfwgwtVyDl8oATntunqeqUs+UuvzXUkB8zQDmSXZ+Y7EMg2JhNfW3DGX
Uuqi91wP/YLHVfHjYNcgEA4VMm87isDK6nYWxxsQKJ1Q84xaJ0doNTB8MKqHxiLW
LED9i6ARFH+fEJXSZ4dn7GUwOlYdTqiWdxh7bxF6bSCm32Z3B5ToC/dRKsoqEcIb
BNg0lu4e1TOn9cDmHnM1aq1Cedrjbu32fHMNABPACf8gZqT5LraR00dJsos7z9UW
Q8Q+OmVZ7nCTD/w0WR17bfHXuXj12mnwJxuLHtOudvxe/FVolNS6oZ8sYqNjFRO/
dwzhPhgA98bWl2tQ/ft0R3jOXncqoT3nxPML2XgVGEiF5xGiCiNwgfQx4bDiyAYG
AtERrR0k8udwq+yuO7RF3cgdqvVZQUlOOflrMIv4AFUBRn3oSe9MkECCuNWYIQQX
LbqYIEpcXjLOtgk1Qv/gU82TOvhNR8pNxE3+vwXOlZn8fYGfuXupX76smOHfJzpK
QMYwy7Z0fYA3fHTT7Ao274UjR+swmGs7TcOuk0B3jNRdARx4kjXktYlagKHxTjuv
2oQQ4Cvf3rkv9tMnFSWTqXsKnAIMyQMKHfWe5J3/qJK3vBIXLfy7ALOjLnnhvLco
q53ltjAEFiKqRORYP9mM70rDJmknZuM1QAErmM8Wg+88SGvKx0X26sMV05QnghSe
xArP7QD3F2Y3YfjUYb/eVo+9JH6vqPv04W4D9nZbdt+UX3vFeQ567j8Td+V210VR
+kSFmDW7WCpE+pcj4hbLhhAWO/6QNEXuRGfNWd5Ovg2lPvWhjQRXwmH3+3DyS+rd
6t0cXy4A0a6hkpumW87AhZz/sEIJDluy22V1LK/MVoYrTwp0PEuwlXTti1R18gEp
qxyMvSFFFJYIIKcUnWkfcim4r2WRQQtVImNGKrvAOanKM8OtkAX8i0yjJ8jMSb/w
Qe62thLjy9MTKFvZzFab6Cgopk//pJZIvXsFwrXGrmud3T8BfwRtMWXWUAHwR7KV
2ET/Ke6nYpTbr0tjXKPUo/+ASPnznC9l7A0xLi6pr8vFQAj83sKUaa7RcgBcpNLf
BfAD1wWkVLqfyKW3P8XUcMRHjzbR3fbzsJ2yO+35Ft4jbN+yEoH95QFe1wXLOwC3
OvuLhJyV6dVK5QEHK5JbJyCJ3O1M16oXevb09u/aYTUOe/qjILBvZXt/6FVTe+T+
I9VIwvKR2XGNT14U0miG6rsqtVL4H09Y66y8r4+0rjjGPi+v/pxlgPH9aCpzBMDj
h1XtqHChQM0bcC4NWHSD5P/sRqdLxPxC+vr3tXEovVTRWmYeHoLVe8sa444QcIF9
HH6kLzhwg6+TbRIYMzDVdguB5vMFxkRrmfGSkFVMyS6dAzIgsoPcJKFFHdxDFBbl
GCs/FQpCuBz/JsuJTZgIFtnpWfatwCFQzIHa/FA8AbVzg1CCYOBMFo0qDremzLlV
UMaThx3rU27Hn0vBerDWOGpzOvKOquAvziBUWwh/Uj+gcrrmfcyWw4EuGrgqNNDs
0x6Gao1qclyt4vyvmyAbDfuCE2cGsi0Ey0g/e2J2FGMswe016sdr67KnfMKc7Roe
0crCEa9sGbHesWHtVVPxepMx5JSxXmUw29cp4eJ+DOKb60CG26NjyL31fKgMs7Uf
YBLcEnwPGzC+En3gwPLRirObZPz383sWQWvXmzsbpOSBYBIazbnFLiyxiLN7rZ01
PxxqArpxypxM0ZxYV/K1/BC660i+v5YsO1PECR/C0QdarqPcxPe41NPy+ZIjy8Lp
ixFPhjp46DhxQ/N3lEBWKK5ma0pu4L+DmfJZpNEP/SY4fkvdUBVaoJetgsdf38h6
QbULH6pbnBlhISmL1HsdZoYNQYt/XU65pkcJFqK6IT6af8QkgUtDxYyxoxymOnbx
FsLo5PlQNLuxI0UpTN3HJ/j3YiaFzd6XwKWAMH7V8ZMXa9Hl5PvKw0x8c0hChiW4
nHUKRxnJ2qFK3QEVsTRIbO/lbTTuBO11OdrRAyDBAQ1NSuuaZiZA5OIhXiTByWtI
BK8QsYtgsA27IV42BotD7PoITGddUWENZtx+YkxCcbZitkO7cIljBe5XqWa3g7YV
ucz38JrXJmYzHbPKc2MfwAzrvh5sqwK9W6BPd7HJMzuUb3iDryBIIfjhsDwEtGeK
JQLU3lMl0EQXvFzDR12Pi6esSDcxFtAfyCnvsj1GJuDtmePQ9LYIiFdncCUOYaUn
nBFKtGAbcyZZ7MQoVrw8eg52lOQvC7VcWkgCGnWL4FgB5IbeNDdOyg68UikCbYX5
T7rmPUKtVxKoNr2hfnrkIUIMmstO8gSU6ZIJYJ9kl5fxQZQ9EgZqS/sYBQfs+Tjt
roUWQQydPbrz9GuXfNGSsIa5EtMmPvKv6QLy2VC3utPYto5oe3EKnhzImFqMp45c
oFxrOnTZnaAinSp4RfxyEUcve2CUCvMrFOvkpmQ9td2BjgrAVMMili6HbR/jhNlG
obgTgs97K8nEDJBNCp/mtod4j2xgQ4WdKtjoFcaEN9PC7NrciK0QWz8o4vQ79GYj
Suh1KJID7AKaeKQ57U0FF1aStamzAx84+G4SgIrcu58Jw4ycYguOT2w0dz3smAtu
FPmAMpZorcPJ68qsFlJlUB+bJ/5E2FdzdOtS+RGQqPY62OvYAMH2z3O80aQQTw5h
e6EohzfcMIFvpYnVwvyxUYFirIc6JPVSlt8D7yIVgIV+EmWONnm6kz7Jh80EtS6m
ZEpmYDIKOJya2/no4jDTygeA0hIdk61Kn2C18tuXaQVireSubtFg5WYoKPmv+gma
mRNNJoGB1/xDyJR5ljp09oiQGJ71CFnYiPh1c2ayHBWqKG6XVfDQzMDCMomUBlBk
dRD+SVTuE3WQgC5D2tmDxP2Yb3kOG537rZ1i3LGWi93l5wKvxiOvWFAT7B2qESsu
9PZobHz35vkqIxnV4i1nLhLjmCkZJ/eoBo/miwsJ6Oaes0oIGpGYnB9D8LO63c08
SCfXh6QPzeV5z1dKr9aMJqAU7UzxfveMI4Rqhi9VKHt7rqtJdyhEHKJDKl8pWAy1
nm0SZQZ+H5RAYFn+SYd3bg5r3tnLS4L0BJj30Fn1zTLgzdFp83YW66dBvqqThKaQ
DMd2sGE0DZNLBiUaOpoZiSgtG4gyeafbCDj9oP6mL/83gFGFhxzA1i23nhE395bh
neRXeZ7yp7alHXcs5yovfg5dhYSDuJL0ikAAhbItLlfXOiQf1/U9l8KuAqxaQIyo
/bUWZvHtHq4cg2N6jXyIcU2d/KWWqEx0o8LPRIln0EJICjQMZi+72fZV1VY26dkK
j0Hp/GirYcMZII6zsfW7YVL6Do0JZx/agpMNtSfHWy+J2c8G1nf5ymfYsqwnVfzN
IviRnXgNhHpaJmJphCbevZs7V8gCsxf5R5smstweWLvx5GzKgy1uLCdQ/55a603e
uKrH9X2pOtzAVeJtlnvxu2HdUBFKLwbHnAxyv9rmUJ9hmTrxBuZCDERn0utYDIDK
Wivb4/b6GZPEXdKOV8QWmigxaD6PK60RFqB8uPaegiid9lulyMQbUAkAoFVOTRy+
ZOj2U27ezUiMWJ3hBY7++PXTwkL3PQpb6xOrXCiQTDHQbI00JARfGCudaicXuf8b
1P3lbo+uBiOVIt1xTwFei+7rp9VGvOiNRxrtNfg57RVX7gSgLV3PqXIIVDP5wBb7
eDF1DVwm6E5//jhsdmjTJM7gdCVYYGVdTKkgDYYNS0wDPPz7JCwBV9qmLEbHq48N
Z2FuAhW1wlPYELQUec49Sbxv6C9nwpxIwM3ZM4n7nv9JDrALAHBNfiQ2aEY95rp7
LfGHJwHZh2X8uBLF3cymC3gMXCQqv/JZ2BCyygqSUeyck9NeKx3F9RhEDwjvMymh
876FgueFqUa9eoCsaJXYuj7zaNYsl/PyyZkBv2b9zMa3ZKj/UM5rST9X0Q91tso2
LbJYs82vmJWaIa2e9GGueBFjaz7sZTKWq/N+LHP/9yVQ2gHgFOZ9DTM0lta43/ps
cXHmnp2neRJqmFlE1bzEeZTIueJegxZeV2IblnWuFX4EDs9fLexJ0Mp2iSs4oI3P
ltLqm4Es0J+5YtWaMcpJDdAa3i7qUtdO9m8CevrGXAYSG6ComFJsmMyPzKKnrDV5
u+BZWfhTWd1JiAm1wISNDGyxDAkcY+j3zqatRoHQwbOIcrGp3aI/xRK9r+yJboMs
N8S70oUyYGQsmibrD61WbtaxekcjLiUJoQezaDEsjMwkmA7SGozxd8UDHodEt8pH
qqw0B0D3D+1xN7urqcBlHgbJVpMqttcgmREr9aEnYDdtAftHIlMzXmB7zN4wPmgo
ZUuTZnGEaHY9p1yv+G1Yf7sMlvvlzeo2nnxTtaAtj+5OikTrc2jemnm9cHTevPYY
h0a0rXF02sJneZay9QR/3HbKYkusPpUpaOJdwCizMSGZS9KCWIQoi7Lt/LusXig4
mxzx+pWggKVXLq3vKshqwolT4s7M6QYbmxQWA9bx+PnpHheMDTsqmgajkjRQNm47
l65eWrv6OT3WdIuAI3jtqZGm59gJYCuUuCM3pfzURWbEDIy9pkGR/XAaAI2+mmw5
LTYCwr9xqZRd/yQHhFr6hWLxjo2UW+Szn1/czkCnJj6Tm8sjcwqWTE0+FvihViOQ
tiJ67OSSmUrTaBwT7ocoHnqcZRmKxM2lgHK6QMzZVn9xZbZW81nAzFJpn/nVWDmQ
1/e2VD9wmlLvM3nCZVkwCvApvu3mXGie5q7scWhKVhL9oPHP+CHAxKIPkA23FDqp
FVLZtDUiMtmfW37+Dx8LiAlK5R6TltfDmuWJLfkTNJyEEfZEIm3tZ9rDmsMSx2OM
j1mavVwXPErI2Ykl1e/chRYjskXIo521ANWTX0fNuOOnQjrLrWeA6R8IiXxJScCA
IR2HqMDXaBaOzAA0XMCSCbX37P+TAojMQlnRjP1Q+D3KaIq+isjQgfuDhE8fdRdZ
ix2ZsVJf4XkoECxHnzuofOeHG0duZvfhBEGyjlP0EJ1CVqtKj++GeWG+HkNQKJNz
jPEcgqEZafzuJojz7QKsWam3fedcKqpb1w/fP9SrC+VjDGFr942zaUTOp8Q2cpfN
uW42hzwkyEJgKssici9I0T0PNaQSWWqOC+H7xD+ruvgh1FPFDVZNvPylnBpxeIh2
/gvBA1SZREowsyOk37glFoqiNmQB3lHuaOEcsz7P0rBIbUo0vBdH2Abx0eexbr3e
LBmxn6/ccTi/xdS+qJX3/SesYWQpFfYigwciFOlxnMQDSvvcldc5F/dHsN4u8655
TA2aYP8EiuX3AJC1Pgiuyb9aFg35+gXR4SaKQoLy4BBbIgf0XUkUpAwbp+7paGLQ
W1pt9+WAfGX9/8j8DpFIImLX0agxdgKreIW/vMBf70L6Bn6ddQKrn/wcX7JITpT7
uB3BNh9Ou2GbF77Wd/LYdrLC3yp5p+htyzyHvhL6qbpf20BGG1CxNlM9sqdxcOkI
VXZyhQBJMC9CsJXcGNDMcnMQ2hbGYZEeyl8dujPw0etXGCy9r4pD1qaQn4NF/mr+
l61WGZ8eA+dYkbhOECV303NKpLkplfDyHBjLXi4SQE8LPsPLvOtH/kr/ydoPtMoe
6z4vVwzsElh59BMkK1Q+DMnpS2t7NV7GOJ6Cf2y1gdxRZwh3SK7BVxOnHU/3RnIT
QpDvLHzm5XXjs6+yjGGeT2TZgOFd9f9uu6x5RmtjxaFX+dx/rUYtBcd9GdFAh+Sk
s0/Pfu8yNS2plG0HGfr4AhleRe2MKudDxVxUCXwXmCL9di0KUOzKAVSyX1nXugZg
eqMpOQxcc7iKy8Urot0D44DBFZq7astN1nLTar2d5Ra9fDsPtxolnv7AsCUroKMf
zKPBdaiBhT3HwDjz1nFHCBVwT9BxZY62LgmJoN5/sO5ZMQKORswxtuIyzAIB0667
NmShHMsPg5KgYLaE/ax/RZZSHuHZ87OsISV4Z6UKswm3IL1dUyn6EJQwVBpxVGuG
R3brwnwga7L4DhFR28OyXXCNmk30HbuHhFM/u16UkFvMXN5CIxkMv3WGCZOUV717
QlIHfMZwRvyF5UFUvDIXttX5SRftst6ZRaursRsLVp3EzWZt+5x6oOBp8OL3AHKW
5t+ddJKi1caCRGduJ//iY/WKtzZ3MixEf+Dug97lbUg5gAEXCpm3NtMQqMODujgB
++rHYoaFRrIbk5sqr8cij/omPCvfYKyEBLAZ3D17AwFWeKj7tUpvYzkXHCd2sGDs
2Hs9TPl8QvrHeY9Hm97OAyx60nEkpsGJiPRXrr74Twtnr5mn5vRcFQgmp3KOFlu6
EZLuHZDJs9BKNGTcLrbzNWbqLgYAyvj6QUa2jPIKkOsZAKXHe3+umxESBHBCaXgk
/8285U0HnQCGVV/n5EHoShCbbvmupQixu4KDlllj1exq4P5SnrWznQwzK5ObgZCJ
Hb0B5eNnhNgBTCCJHlkefI46rtZzxXiwKQoLU3QGGkiL5AZZmRRhoOhepgI2wxhh
S1yQLuGXc9TSlqrNaektnDF0Nnm06YK5T0FJupS/z4eKMUZgjZLvRYghUglGhHqm
UoXEYnGxwpyO+w9xOt2rsZQB4aV9zAjxxPj97T23c4mr+cr7cMWIXdjo+jViQiXF
uyygzF2hylk/sk5l+s3CFzgxOW0h9GNVJCuPnTPZF+BgazBdon1r9qw2rK3fDlhm
n4pzN6n8YXWq+ZrimfDQcuXl/M43hpFLXNNWgr683/iEGETm3FMV7ak6S7rviNBL
rS4wt8oHs0IdldW6JpuzLM2asz3baf1rhycoJIhLc5ikqiGHzFSMzjK67dtYUL4X
Vz9tN/lfIDs4zn/xZfVMtJWUV7t8Ja4WldaBnDT6oYceW0IcnDG1pyLASZnl5U8Z
4pDM5auCoBgZW/J6mvlg7UIN1n2/4HtKw5hGcRLXVwQ2BZfxCMXxsFpf+N1R4Gvn
KQh3sFfwkBmpAZ0G9h1aCjJggQODpHvJ5iAbpbbsarPT7M1p0SI2rjgBCByNswUW
iiqQeBaGKdmE546q05pe+0eush0zljM/yCLfwHgyTyGSHCZdch8uNFWN0qLltMVK
W5DJ1vmm83o8RO8RwQLoMXwIPEGUURnAuIiz2UZmmypmyYV9zAZAiX7Hz10mIACu
yhmEcd2CazYGwwP9E9pRL5CNCLijYXNPbTRfv2mg2Le2T9JLlIl5u6GAsbf2UaEu
zqF5oK4DLXqzAcAK/RCftOgq91U8w1HMs3YawDFclW/U9dvdMn8jSULyTtBgEQGU
ftET5zA+cv5V8lb7mDcZGlHL5I9tGE/ez2o3FiZPKB40TiLYp3ZLFrFiN1ey+sPP
6oBmfmP9ruDDCV5mWFwv9dFBaYdo8VDCAbq7TuImj1orRoVC70gPtrb3ILDwX1TU
cNSNUoGPBVQZooqH9/Blikm0De3SQKpBJLArUfQ3h1Ho0jdj8fEw71731e4hLbNG
SNr/ClMJqar6+QrtLkLGU9CfWQY/omdDGz+Qjn9oPLWfjBvL/l2JhZT64iyfTcN1
YOmdzhuKq0o9C1gyH2fZBd/czT3ayZe3TdhWrBM/Fdz7bQ92LdWJkB9tBcL8+MHY
S8SvSj0X7p1wUgqsGfvvEd/7LEZpKmyxbOpbNWVldKJ0fA+dfThzn4kVqXbPD7Ts
TjP37BS72GOdlZukd/KNsKpirG2KrKSi6ksXaFoeQHekwI2DvFisdTUKrmdIVoDr
6P8dCTsgbgwIYH95MbfvJDdIXW39jvfj6/SANyfMwU/BHEFLgiblOH9pP8dWytbP
gkpscGThPblRc/gCP2fh0R1wf5Bw/+TWxPtUNY1FEmECZGiy8A/KRRY7z9TYIsRd
2C0ml3RnBwsPuE97sguLuOIKfWBUa/ONWV921PRIX7+0iNu38VNQAtR60yL2C0pr
yUL9Znfq5vN8eM7bO0zyluWTZ8KLWZUyS0BdymzzK6F/dH6nemWACgCSmCUQ2xxG
LHn9GZJ5D0rma6AJwZp/7NEn+q8w+43v4iMuqObRDRVP+qswi7U3ye2PRG9BqHm3
+KkG/YeAct67wHCELTn3Vt3Nklddas2ASaIJRIrjP1VL2hu83t+EYfr/Iad9T+wZ
k6HFs18nyD+jOwuqgyXjQzqGgzcpYsAOiMu6+n+u5X5ASfMXFqY2J2y7Dy158H95
PDxLOfsuOYkZSr3xMI2zb4+UqY2aojxh8QwzGQEb5uk62si2YbBJQ58NINlE4oty
0g4qcN7dhIKgJZ+wWbWrqnfDUfu2cm8fr114VqOSDb7eTAPhTqqxrctWvYwCPwy8
fYlZEdChJFzD6kcjQGMET+zTTcmdx6R4NLJGFPOBBFOr1U4vmIBeXtM3x6rLieRi
EIeDRxR8YWq1r18IjM2KEV2LtIW6C8N4IwCefJI7urFXHODqW2sxYb/013/g2sDG
YfTv70GCQxGs8Y1em/I8qxSuRX4SHluZwUG2pu1k+tS0Q/QvoHQ6oq0xVIGATaa1
mXlOMNHtOLuU0PzUsX+InoUZc1SY4Wm15u5pUA10M8cnZVav0NdipsVhRzOa13WB
bHQOWKXSSj2lXiWKbV09gpChqIwdeBIshzuYoDY8rdpJkP7GJLmXBrU8nDNekduv
9D2gqUYD4CU4ABVWT4y2JtTqepehjhQ7KTCjJXyNUGvlDbGxRbmF9B3Jd71Osft/
MLZYsAGZ9mpgXWNJ6kjGAV8z4n80GdNshz4+LZ9hl2ERqvAiA2ROdeALzJgFjMuX
w/0JAkyk3fusD5wKx66540GmqXTZcOdvDao5wPuMGp8dMofbCIXnMdrNsygAgWKm
ly2MxyFbDxmXbUxeCYF7tTrRBsaEBC579m43vFAzkQvMnroeKdCIWNd0PGIxQGUR
bYjbUVwGPJx2iGxEpgIZFBADq05kOUglIl9DRx4LPLd47Ts/y1SWFsabYs6SSWQY
Q7DRNXbw/M91Vo9cTKjoXuITk08DmlNPI9tVggY2vCpnPtn37ANxuVMumW3IgXSE
m7SDAK6Ud/FWaj7WA3W26bwlgA2n45nyI1EAzLnqbxgLMjgnaWTi9ip8B4tB6pmm
uWM57obGjJJCmLq8QLiUsVvfwwP+Jb2S7vxg7h+H7n6aB0wOR+PWcVkwZpU1Ve+6
40RcgefqyBSES0bwgktzApyD6JBtGi0vHJybxN4E7Oy4lFC1Tjo+V3cm20W/xAJE
PTTDpKfe3cY1Vz2OmvEJ8WkXfeFlkCgYS5V1RpxXpojr2ZqkTynZj45I9FvFU90Z
gClHN3Y02O13enuk/pe6VoUY29nuXaeNq2vpNz/SNsmbEF/D5fpRzHqqrTUX6vy6
InmJYcQsoGtOIOj8gyzNjdIH6L4QRuKWWL6NIU+oTjdmzmqpQntn+y/16ch+R4ya
U1ucd8KU7dGncSIdiIA8cogGm8C72Uq/TvAYxNLJWJdU8vCl7V5R7iGo7XA4NDE2
CBCCyx0zvYxnOybQ1xsK/t/vbPmUzMSMggBRGPwwlsWZe02z2yzzRP7tGN4Wggb7
xtbeWWTQ4kpnvI4CTCL76zoyZQxiJFFZrOsUPK6rredYOCJSdir4AX3BRSMcbi87
7TJGiVxDkTObI6dIGc18zXVh3PPiWlg49fQD8FShD2F8XF5YIZTRcCCwNBQRs6Fz
VpoqXpYfGu29wv2MfnQArXSGeqUb5+k6zY+DoDHUssQAjwny4ZcnYePvmdnMS7be
yLeq+Vvbu5QZuiXVWqXuBvysCiC5ZID2MPnmeXFTmq4bdRwNzD6qQcI82RgveizJ
tGyykTULD6wD96midc8dQ1Hlw0q3U7HQBy5KPSxbsott65E7HLkDEj4wqFCXfl58
SHe5H0bCck/MEA3DRQj+iph42xHwKeypvjHsdeWMr2gbQjTMbOgGuOR0vSGbuWRK
ghL1cofhjWimR4lv4l94bcsW471hC184+K5o6QzRwZpBGQCcYOdWSVxwbMs1icYj
LyeYiegVI37AzwUCfhw35f4n1tDP2CTITCTPg5ZZKfeLovPlB5MkzeFdwT4Abk9d
Er84SDn/ttOpezvRhsQ1E9IUxJJUWZutmB1WTeu+g/yg8rXaakAl+8dzdi6FWwqi
AWGgNRAOz0UWPTIRv0NEmtG+P9bkzAlM7kZIBQBRuLQWy7PK8bXhL2cqJ10EP6pr
UXKrqhOd3p17smPpNcWHgoztPG+opd+0JMxw3GCjhByRDyptyChPoE8I02ZZ9taW
2YGwiM9oIJa4XPfO7vrAHH53S4LYUKF7UsJoa/rHXAxwF055mPqO3u+8EGkuVHAr
XJAgpf9a+H+WLFqa1YxSk+B+xwYcxMpeIMlB88IuP/RpWlPkrU2/kucouihxpSMH
321JdSzvdN0VnIRIcVa+ri3xFj1zwcLo8DrWnS5KXC2cpoFdDD+TceovM6Q+2AKz
+u/nXgoY/0VXxYUwvanaOSb+26Bw+zitETWLBYrV8vMaMFicxHoN7AeVbgORZeq1
ayWvnaeA3/Yw8wkQipCj+Wud/NwTqCgqKJ7QTRHasTyYJbzNAXb35znz3q7kLzK5
6ndxqb0wKuVSIJKUbeEhDNtn4xjr4Q2XE0gZ2DLYaKVbO5xjxHb5D3BpwJLHVfN5
p8HTAb/JnuvEPRM6lbfgVNshSpza7rYhY8W0repQDnL9b4c+Nb01f0mQcNRS/Q4F
ceCrg1pmXaS/JRySFAlFspLc9UyR4Jw15l5kadvzMl1srT1tVeT/45FXrcizIdzH
LsJFBNuU5jgwZS4XiNP7odwacGdTt9HyNAK2A+CANprLfKtCUThFXnodKyIMri6b
OeYDjvwUkbiZImpF6UYnx+Jtq73LQEs79f6ksyMAhs6fk+eJ8HiYT8xFBDLryCUz
JEijiTqWUMuUJj7qmryG6Ef48Zn206l7mhL9fcX0W1V5/X0ocmAxo1M09+4g4poo
MdSS7EZds2GUHK5gu2CaDmXmi4WCieYLPat6xa3rmIvEuYbi+wrxm68kAgCEOhdL
gVqy2AGuwaE6D+j21ui+jj2PKU1b85mIkI0ZlNdpYG6m88zifTTHy4M2BfU45Hso
P13uoDVlHiecTh03pnaTq9m78uQlyEB6L9VgKiOGzsZACDXwP9w3uprL0mdgDN9A
clK55Rms9Qm3PKoOewXsnH1+WNSKD51v4+lZgFLhbFgiVW4E59GOOWWpdEuxpUdH
63Yp2Cr2+NAkBZbrCN66659Z8iHwNRpUMfnXj0G1Y0VRm023bBg9QFvz94iiibVX
8spkd8xnwiiMf1EH/t1GsQ74RcMwUpKgg4GD6+gSKcmHi6SnKDmParnNOc1gYwhM
OGisK1d9sM/Xg4wX+cCl8OrSpgx9wXQ5H+WnfyO8dWhkx8tLg0Vd6BXxjGZoflXy
5QGPZ6MMsD4w/jxl+ne5jYZar2AEQYx2aph0w5bUy7IgMm3zaD6W33LndIFzuJ/x
mpw5JTqN2VIKR4t/nWCh6h/MBbuWeLeMDxUATjkCSxsYnO9Mc8016+s4xGjAUsxC
gxT6Phz+2uQbGmFds3k5CSWDVbivhwn/3k4go6Lgnbtrv1f8rQwujVZq2pTsUmWw
YEvumrawtDZIX9+QfopXip5xh3NxlGILP00MVuaDoFHGjiSk6gX9uTRD86Fymk5L
bHRcYO6qipA9B3jUYHCfdjTu4WSjmQLloFW4wZ3oamT/TnPzy5TspUZk+jLmrFir
QqfOMjXtwG9X6qKDfzX2CSFWwMrPZ9zWAlQ0o0yEaJILwrnxysYtA2a5JNyXo1XR
Y634iLLBUAWcnXYL/mihP9iqmZILbYRHpRr3qQ9a0d4Erj3/RUOz9dwdVzYjuXIx
GxglenSAeRaoMmxA5kbEobEzUuU6/Is9us+/wWhT/kEzfRzYW/6lLxiHF4c5BhtL
sPeIELvLOeulevM0SCXUJwZMyrtdVXQmlflCSpPqSLZupptJVoNIhZWPAColC5sG
TEE5L5Sbqzj1u/R9GLwMSr9sCVrPjlvmGFb0N5OLXARSsAWZWfRQ8uG48IHS22OV
01qK/bk5h2BqS3sAS+dWP6J4ROd9xbaNU0QwNbTvgeFIbkc8d0Kud37ucdgApYD9
/AJsWyUxoPHBdfSusILAKi2ALeP67IjICsbaDa4U44TuXNkvw0vuVTuz76advzJ1
HYUt1bYdJOGiUvH5SNQ17x8Md/3/eIkPAk+KLYnZG2vfFfiPrEETYIfDdUUA9F8e
gdEIzOySY2rISOi9mnO5kH/lavgPxCygtEJPrV9oGPL6oMHet8Sihjp8Fs4QkyGQ
fBzf1XKUEdsoJ9LV6SwRCAQh0fWwo0LmlTFS5/46JB+CIHPTQX9MWT/yY657T/2d
wDCBqr+3IT/BSJgHUCZFMgn6UFBeUQL31owzhzQS0qXot3jONBfB1oBPzfKIH4Nb
pyKxHX934IiXOzugf7xjIyMqZqJV50bFsWyFhTnI7OO7V9UvAIGfRLdtO6gDFzji
fRvLOg80ui0ItX7eEVZgqQ7I6kJoeUrzOqiAFu+AM1JZTnb/ChuJY1BDOtViaITr
Xidy5SM61xMbocaKMztoL2gqHccWPf0VNN5p+ek5NdQ0+9OIJU/Ij6M1zA6plK7T
vXzcy6sSDSJnB3wQDnd+FKkgmxerMl670qhG8f61w8K1qAk4Uw6ME1y4D3nEne/+
l6bz7kqLfrCeoQ6VKBRjZBk+nbdST3vUkREF9hLEhYCU1Xql4CMi5W/hw56ezrIN
7ywQG4yxPrbBN01Al1NpdAP6lwVOuzkTGcdOgpprCDa76AEGZhNvkiRlBwVod+nB
EbUM/uEKm/xp3JfToKvGw4RhYLx3lACzs8WZHJWbWSGxLkQiFYf1BiRjG4YugC3Q
GuzAiUvJ59FKt8IER/Hlr0GNwmIEldcORNAucBD4AHZwBwnU2isnPprRXNsSpUO5
rvLaZEWk2otjuPrHTh3H959F01mSgloXhbOSGkzoDEvzsX3sVuOPczFTQnq3uFbD
wggpD+Ezi29xnogK8C85Lcdb4TeHmHLdOAPkntuQQV71rKM1J+ZrNGF8Eq73CJJG
dLlGMP9bquUBzC9OspQ+1/8ptFzyRIR3eerMUU2PYe1rBJ95hpehWiAHyjIWKO3Z
l7TE55CSHvFECREWBk1C/dhXzYNlSRfSkiI20e0m5fYuO6+mSyRqXLaxrA0vOu/6
HN5L5IQ3DA6lw+kTX+fRNtOJNt0m2njKweA5N1c6UXsP9Yv7/qEGqE3vOs17IBG+
6z2wFpus6k2acO075e0a9WN3WYzXxJsbiFQAIDQPuEDhQzNuckp97tAQFdGT8U5l
oitYLmADKRZJkpjdl4EIh33/bTTdDfyNb3QkUAjZSEcU4w6bm6tuQzskj+q5ffjq
19Cu+exLnsVul5Rw1vlOb1epsVJmemr7vbsn20nZ7qB7j5dI8HB2W5VvRGhYhUo5
S14St2YERmNQIVYOITorkriA9IN+J7/Wd7fDOsEAcu4BsviEOrz0QvR3GUaje9Cd
9HbfhUjrv549kjbe0w7i4aILKXInJ2osJU5BrC0hxDag1WF4+zCfKpitApEnsIhu
lYfJ9h+iqIc0fsdPf9duVCN1jcwZCww6jH3qiCOytnO1+ivGa+EdU2yz7Ptv1UsP
jbMWttM5gUaIwQnjSEMIf8xar7GbaWhPqMHNRMJUlmbhecI11xw1v4NWC0YkIk9s
9xCIQUY5FrWupVegVXwT0YKNiQWuEmA17XEvokFMC8HyrlUJRw4YGNghMy7QHIbb
NiHZlMadse922xpN7SaqrVo7jl7cRDPqZUqNyTVWm9G28SY7DsO/RzbSJ+7G21eX
nn0OMM0/+z0w4cBFWu/hnNMM753/QnEGThetF/mgGGhjcDoz33RE8MN/4WSy7oNn
XS6XLWTWQl9nVykHR+t9fvd62NQj0zJvO1fnGZhjV8FXbuBp6iAJ+Jf94kwsVpPO
g7nYNi4LsT3LWeVk6ZbZGXHH9x6+HJ7l/fwiKi6Lje77kd0zikOyWRkAoCpxh1R1
DGiUSJGBw4G8HVzoPj4JBr34VN5DztGay6vurf3VC+px9TmAp7RSuIxFtYMXzmpH
mvqFPFjH6oWWAisE7IHExSQj2+6QWmwc7kF3/Wro3F/NJfoRtluyQhGzZ2qDxPM4
SZGSPhmXDI1x3xNny3ytWBsL4G/SewMrZOyU7NPaa4rsN3GAX9oRAiPLUHvBni5K
E+b6tDTjCHlz+BP/szkDsJ/iyYCTdY3SRSVSTEY3J7EmYGZsFge76sywizcrMvyQ
b1G17Y7+hzmzWeSuU3fYznbnvFbxH2z2FktSo3hyb6U6M2J37xNzl/7m4erJMveB
bQf2lrgYuBlDsyYy5BFMnJgH3S14cUgPZAL7olNwBSv4AqcVqA/RcICjEDAHIu4A
rGUv4pWMKBLhdpwWvdvgPOrWao2fVJmmEc5/HxRRBmqBWCTkk+LyD4/nL4SHAHaz
IAt0Tf2ANlPlRUWvo3nHBg0rj8bemLU4W2ziPddTgb8JFa+qMTwSxlvNebambS3v
Rgs/YHqRS4XVBhM9Q6HHKhvzPyhVxMcH8srUGhBDAKevwQdYBoorKXycF8T7iMLG
fDAzCeOWTfmubmpVFGp5f6v454q1+fq6thNolPLrIAC0pXIoSZSW1grJxR9+8yis
TU14nHSfNdQWBcsx6l1E7cc/mr7NUVdAqwlHqVLOWvK91TTr/UMTswwveaOS+xvN
Wl39c+8CkwfV5Y1dlUKioSS1guELuTY8NP8V8OzhHp2mdOK0MATvkJKm+daVZ8sI
rOeyN00v/OvWSycp2BZOHhOKDOE2bcyc/ff4CETm3JR4DlSH4CB5zMwtwCbt9z2j
LJiQsY6zYO26vvARRGqqtBcVglbixH12l4mZSWHLqc2hD8cXzp2d9V6pMFhvQWWU
5kceIWtZxcMNvI3XbmArV3bBafCl6eCB6+wW7Nmip+L2MxxmgnMWBL+v/hAwt/Cg
F4bM6r+ESYy/nkBOF97CeBEusdbuqGGsgYuwR/jz3VY3tkjhiSntbY2zZX2/pCTS
MfBJec4vGANBrOQ1nCxcfwy0NUWtCGLHVxs06F5BQWoXp7J8bBW92fmIpdLtkBVx
kBFBv8AvPwH5CEsy1hIdQrrZ6AL67g9hbQUJcVNilVpcPcQhvyEDy44hjy5/aOWu
O78lxlMuCHlOlM1wTbXIrFYj4ylyQN1uES7munA3zvUeZxHSkqzNSnY8753jI7X3
HwUORUqOGnafVyy7L6RVwl+jxrbJcewVRDLPMGCIXl9ehE/elcR/4pEz9IY164DW
VfZhrb4Qjtk7x0rB3FlELyR8fG3WnFexehvRVJyIFQaCmi/VTwqEBOz7zHqSRwNl
O3Ix38epdvUKDYQ3MchfChEwI3gUY2f6bCj8aE/sbSB1JIfTwVycvkIuDG78MeIU
DnNo/7LyyBxp+DrRSMetFmQVpT3+b8W6Akhmqc/IyHvdBTX3vWiVpWhxqLdK/Z9+
bt/D8WIY/lN/TujzQiUQGgNqFDQyZNxn7MisHWILLTRDc/r7k+1+cJKd/xHTR0ZP
HndKx29/W7cencL3P7sOuPbFzHBqIj5wcoWECy17DRra1BlqUrXfuz+gnIClLlRh
uw0xzjBhmgSGu3e322vvWzBezjQAz1nejuas/ITxoTc3zEDa0Oeex4jO1V/ubjs/
hHFTlYr42TKYuj4kk5EIq7Qu2ap6XaUzBBWVN2UujZdQbmltWoU4LAsVpn/z4Br2
Oktt1i0mUwwhow1GGRIWRoLldaFU4NVayoBOHvdqgUS4rzER6pEvhvtUo2zrsgUm
2pnwIgsfOS0XhY/ZmxiFuh08l6OYzLgmzc9IWjMwYuJV3w5XYkZaoWkyy4d6RxsR
lxeIOz2UQGCRMmFMZmbb+go1GPLVUsDJsEPrXIAFF7nMA51krx3yAjtQSmmLfgTZ
J5G9tZ+wpW6DvlMy6APBUp+gRJ0aZ8LrDw8Do0Y3qt/IyMRfthwpHhtPRweKbUrh
BmG2X2f5N9CKhokuNhs0W5xYt3SUBtp/8PxPX2IRkal02238pCyuP6QY3R914QEf
RcbGyOYrDeunhhbbPwzh5ar0WauWnSyVgmG874QxEyIXJBkY+mD1RwRBCZBNcwAm
I+WXIYAWQifWcMaYnkif/jugSS7uAli+bEGtBYGKM8baJvtZAVf4bKbBTfucAWSg
4wYxWaU8a8VcylYlVog7ls92x99aLETxqXx143u/vkd4EUPJYPiK9f5qhCsP2uAE
AlCskIDy+GcM0EqPxWIy+DbPV/kdEh5Og3WLoxIMMgyXXGMUFWbZr2XsVXi0CS/8
p/Tr/m4OHhnCAGZjozAER+0f5iQlNeRvZhE5Pdljh1ka7FmBcva8qk/VbnQY9m/M
MtxjVXVTLk8qrRFCKLdYnJBDqXjuWgyu/sotSe+UfPzXDBBhiZi6KKpLwfyvulp0
levCAYLefU0FQIUSVw9kdROr7A4GiazPQPWzOH73GvKOSDOYY1/K2JUWyGDuxzY5
oRYH1qdRorkPR3PcXykLWdMnoYbnQGUtWTG2E2798iMFFiRus4oTHpTUUT4yTKR0
QBES/tud6LLXmLiHmTjqBQ+3cH1my1M9Z94SQdxlHwbdN5iUHQqGSnROGo/ewy2W
jwWgBtQOl4CFX5iASmD3SNH/2NYG26CUePVvfjWj4CJ+fNc5mXkCPOLZWQcWfhuG
yiUiufUCjrdiL2XyTBVZXzrIDCUHnA1LA4gdLqWwP+x01oPZn+7FcPH4T+ABbs3Y
/NttJw86aTOQQ7IPtZX1PQT2MYGSx47E53roEDx7yrjjGAQHMvb35IorAypR7Vrs
fQg1+r850suXlquH2BmL50SO1ZAR3fJU8DYXWICHBobqvpMi1K8Yve2SnOuFv/2Y
Pp7oMgYqbABS5ARbnP0OR65dSRxygIoOYJF5si4JP5yCTFPFV+pbSelSPwqgCD9C
RbrsmBQkpHR+vCy+2WhwVbXAKKF+ptBJgMd/AJ2oME2NsLUclxZaZ3A9fOYUV+mv
wYtX37YwvZwZsX3eAqNNFhGBEun1qSZoSvNSFJnzPLK3iOdrH22FsKZRZnli4vDO
ps/RnkrtEd9xWzqOCkcJXZmY8ThZbAKpQ+AK8GIwVy5PW6vOijBmOZxnaq5893ZW
VH1D7ZbQPZ8FujD/jtDhGCV66HTPN3UKIp9QNnupCd0J6lvezwppuVd77uU7TYA1
ov0F5Un7b3OdKsHUqShEyhPC2GZL/LETtvw8b11M68Zuf/FfTmWD3zQJ3St/38dm
hD8IzH1I8bgb9rxozWAHe4O1gUEG/YI6NnwZZWsyFVBG1nZZzfJyRSENA1yJTkco
c78Jx9taHnUFFva7AxnM5DTLWJ4CqlCbPLvibcLzEm3E4MnqaBV63wpmm9/kBIoW
Mac0ZcGimE4rlmkRKlw603FyeTufokMJAeAY29NXOp2NofJsyaTn8Lq6QEkoZusi
UGftMcYSY2rHD26w3dMYLU/XTPTpmDcPNo5X/v3bjGmzDinmpV6btRlqWgKxwLgd
5fhfQw6pMyeDAbiECpGvxbPEmf1LSAEpy9mybNDdwVCCxZ6Yl2jIFtUZCQrPTLux
+Cx+sFQerFFiG5JY5F2ztBQLeL/RC0w60eQJDO2ItVNVHEcHAJL1aTHeXalww8Hy
Dq9Sg/G4u/Woz0M+AgDZnFvH97yLsjo1l0LFW56Xy1kaurv0fSMQl78RWjXUKSNW
FmrSHuQa5nRBGLHxubnETeFO4mPsNZhASGlSdvfwm36SGrAi9w6oSuSuX0/sir4H
gkEXWMhBwefk0H/d6j9eEGyOqBWX93nhv0ZG7aYsgrs0vf8rDYksAqUvl/1T4lZQ
yKNtuLLTjxZSkH7lGxfR+dRw2OO3ha1Jlsci1dZj1bf40dcOZck1/CwYKG43Gwth
w6/KeXJj5Ht0xs3LuE7+m63JwxVqzKZr3k+t5muNh1ZuB4EDI8Kw5J1SM8sSQZCg
mfcJPiRUtClPuXgPB/NdNRzZ/YiEU8crQmX+iJNueNf2dVZ4vroHe5QJoYMZIca9
hcDBdkzF4aRlGGry+h+YjYs1YpMDJoGqjo6OODPqNUrE1/e823fSy3tX0QQO684/
PkvrmxhDhYjh+ho479qxJtWqb98eDJVKSnWHDVdsa+l3pA1yoi+VNSKs0jR/Xi+u
tGw3BNXGnSuUwWNgsbdMBn3qeRNPqqqjFQLJZaCvBgCXQtl9JYNSArvXZXg5CmWH
3MJedIm1vygfZAfanMfihIKSNMy1YOBtoKz+Q4TntcDo/KU1OhgaZxTo18Wvd7Dl
hswixynUh1e2ULixXAX68WjnIEJKxCoZc2VBi4h5v95fJE4nivXUeAsIpPAmj3Q8
siZsbJNnUc+g+uNiGyRxdXDajJKdNb3iC188AUWyeSlpqq1J9TClGJwpQ0MShoGI
PnMDHrW+RSluWgmeOgGOQQZCXCvu1wACCMIXh8bHmmsRJcFMCvbhegyiqlZHl2GP
QkWXtHOAz2+GBi0Rxh9pUoYBQ+H2mheokVICvtl5KtVaZApMAVFQuENkoID9Us4l
UBKV3UHheuHHGFDFg1mywzvm861SUlFpmR8mGoNeDb+ZGimEedK9i5JZDF0/A9/p
ZNd3wnjpbfwSYXBZx/46sXs+asaxSXoypvK64QbiuUYFGu2/LdYaf6ToNK9qWK9y
Tl8rCMYfsWvhDZmjvbMJQNTfHQ/s/bf+eHIeqF2mKMuAMVOhSY45GYWVAA6/vQpy
MSe5/yIY+VEygF5rklFtz6cSF5lbw81uy8fJxyujbj9B9l2+PMSL6Czma+hwYbDo
AabC4nGSA3OBHeVICPdgUPk9wF0kIGCLgP0WfaWQBRxi72i3z38WETvMUmFWmMPb
Tj4W29wGOsugCtRO5qYKNHuNvgj/nIY69jBXR8wYAdt4YEBp2fA+MSYmy8WeqVS0
M67ct+s876sVlvUnrytLjK398VVTfpIx47rE6r0raB8gr20tg1YMWnOiPvG+2c2s
WUlEnFL/MPvaHJQRn1K16dm16nhxyOTJu/uyUXyEI2KlpEts7xekhJojcF7OZqA2
Ppk8jXbgYJEONKJArKY/77CP84jkASuTq3PY9D1d6dB5h/A7cuAV7y2CI3BBw24r
3F0mYR8RZ7kQm/9Mq9kF3rHcCLxqzVN97QO5BJlz4Z/j34wLL1bjszSyQf8ADF4h
7TJT+Uc+mKBZQkeY4IyckAnLv1Srh6q4GaHaOldMRmk5e0hqIzyTF3ZLk+P2ppsm
nuathKBCl+Ewsg3sNNvhSS2cfiY7ZGFu9t5QYZiIMtPGwWklDRAKHgZ6XkS+8Fq/
rEjbia/t5rizqpdKXRUxWlogzGWGAeR8V+oa4X957pVkl8/RrIs0oLCfH4VG9CsS
h8b6a4qtJxB2vmXJVDb1JsGcIPU2FQriXznLVXAGpGqTBFNTS/0oMwJrjJkFh0dV
1l3N9kqDyX4sIH77zz+bQUFa2jrAE8FJTnTXT/o3naYAAPUfK7S4CMJCRyvw1PIl
N+yzHZvIEBAmzeMqiQRscAnCbp6z64BlaTNOEN3ZlhGHBOOIBu3OJDQ3+fzfPSAo
sHY2Rcnrj7jYxkf3X1dFAI9GJwEYvNRTvsghqzGJXT4yAXtQ0mwI7543YVYsvW7J
8XzAWmcM9K2KrLdKsMGpuUzCzKs7XaXFgODm13IFQ+0qz4YKzbEMoDL+sD081Pje
wa1bNOHcsBXBd0dAOdZVaH0ojC//d6+klC9y1wGVREGpYDul04ujFOGJkOOUACKc
d1MylN9sHNR1IepIR7ibfr2Jju9XDFJYH0hKThjpXKpfF9Xeb0542OoB5AoBVTZd
vucGGpwaPJ6VeBuVoIcnCwq+rbuKqn0Wvj/NXu36F1FQJ4tLYw7OKPT86nL78QNc
2xOYK6wrH9uUeTednjvQH4NMwZXFTIKpf3j/jBdWdh5CO8k4pHHzv3Gzs50tXyTD
KT8NdWOvbkAf8GNng95HbqkDbh5pMQxf/zexK0BcPGq7dXrnu185Wn7nTiVktXKI
z7yanuR1FmE6kQuavDm2NU2ajRRBdEQfiIXpa8WrO3lIIscgSTLXYEx6ltNJetkK
VPCWfvfE5I9Wo8HcmfPhJIktWI6+Cjpe3ba8+PTN/pYrw14kIc+jf8GvJxKdmbsh
VsP6QTxGyR3Zv/cb1+S88sbzjn8+C6RjE/cP6cKUBmrm3AP6/9dDkeRo/0nGiGlj
4bp3Xlr7CWHNx7cmr5xP7PiWEz2i7QSfEaNgyb1IF43R7abJVJZYhdbwT+1RpTFl
zdFNe5y65MG5x8bRe9BMmyZo/mTRCsKWZzegmaih61O1iNctEkrEJ3+itI9to5+H
mcs375nlZ5GiEClGb1sUL9/IMRzfAaivsJZA1UBv4JGxaS/S4qj8CyCIZ3LiF9/p
1iWTg0cUtn7Pc89GO+bATnR+pm9Wt6VfEhao5fYruvtTESYiGWwQC5logQ2acNsQ
Fj6AMjE6/+snKpDvcH+78lDrvUHxqa1lBkIyAAVPCvPRO0zFe5V0A3jTClGsPOoQ
V9PWI6FwIVI3GCcNSCxLNuCwpZeSmonGpVgoQb0OFevomkjO+6/XNATrXqtjgums
ghOkOC01NQzVOpSgjBh+TSwJi8/5+CmxrQR10BKbti5Qf16j09BxbYBsR5ec/Ho/
N5GPXu3ANk8fb6kLy6ERlG6t5huWMTvJGgQ7+Q5ClYMN4JBc41rKcwn9yHsS5zYE
Qe1fWikUgP4THXyybYUaBtftSm0d7KuFHiS8jf0ZQWaUCls2UWcKLSdz2ThOvi93
z6faJGcwQgDD7h0rltdVfMFu/2FXzt/hpfNPmTV4aNBU7SqrD+4oV4i9F/stsnwk
nJalfqdJH2naO7l+E1ODyfhB5CLUwZUnuqwUGyl7nckZOFVQ7nI+gOofBsgtjq5R
5M6LWjOWsH/F5bUP77dOJJRMg89yhHpaNMnIAAOKcLkx+U0jsQ8c8XnlH2RzPqTb
IvUAP09wtg4rQIto3albGD6Q+3B7Y808CbGfc11W50G2zCqJA7VP0Gcj/jDnIngP
FpJK+ErU92TmNcxdLGJgWYjt3PRl85OY1D7nBmXnYwQH2I5YHVXtFztNVxSaIb1e
uxfh4Wro+mXsYx7ss3fgkonTMgH0rDM8RKRoMSBx5MMKISVhBePGa5867lrRSORw
JQPYQnuvb0KF1MaSAvhb569pN0TExICoRzJ66r51PZdm5KxufdXCuNKyXEpCMxRh
8gXSVzN+7c4iwzZ/WFnoPLCprcRuZdtzoMNZttjMiH33//khI/J1uzeq1n5WCOKh
YqPhiZZtX/X+A1+e4X+euUz29tSdgx6GYmXBvmDO3jdubzI3VhahkCpNsy/1GKp+
UP46HcvWcy+oTJ9HFM5G8WDF/lKQKFI6vkxS3mzrP7pBsYSVQmBIk6OzGyl846I7
ovYmzkwPbNDIEU6vntDTq2HhH3g/EP3c1TaS2NhdrPnC1T9xqV9sC00FesL0SZ+C
RmxVB78WRBD0SFhpUdSC8tqVbQ8jnRRj6kdPkU4RME0wJCm4DMB091xxQ4GAWA7t
raqT86UOCiN0dQ6wPrr4X8+Maq3EQmB5dNIXV9p+pKaYrKuSwTv7XwTDxKmTBcEh
s47o5DJHDGe7x+VLhLR64mVod88wY2lg/ZCmAeUXzsttesF3Gx8e7ePlnEWzXgzW
hWSV/qNU4lI9LnHE8Y571WDM1WUrJhg4MbiTHYK00KcY8eQGNoXr2+rcFuCDfhaX
zHagITTqHDn72J30nSQAiMNg723cmk4pB76R2we4Of9fF89wEM/aObkfFFxHhHMf
097gjeCmwWtmz1JHjGKqrPV7WRp6uyGDKI3K1N5SZgQzty2fnXqSPEmcxvBdv1or
cIAc2tB4hZFaFrxl5h4LSlQXdZ+S6KTrbDTdvhd+WoAxjZqkkAoiF3NnTZiyrJqG
DxaUV3GNn+eSFNzAtFAu0QHqw+d2f8YnH6s8L9avNte73mMNxQ4mwCjxh6MyJxCT
ZYv/9HkxZdMcoeYGsgymFUJMHH6UFnxJsejA2bB0xybvM5MbACg7IU3maJwdEqOe
mTz2UQDRVmDuBM4Wdceg3rnadKX0fuEaeb9sQFT9hFR0PpLdRsB1g5Y9tJ/UICbF
dT1E9I3r3kjat0qHCA0wwwfzqgSJTi/noJt6U7eaO9B4SIxolPt4zjNcp0PpVdXR
DAA2BQiPIWyV53LxtTj6k0hqNqa4NurCBsFR96nQUJRuiDL7CatAE+lxGtNIyU//
IWRoNaE/FQpKRBbJCYZbORGCtXYbv3fWbcVwleimEkpI55cAw1HBR3hWwD706pCH
ncrP7iurNMTf5oI2J3y7RAYd0567fLKJsQyFviLRiRFTGHh/ef4HTYTN4J6xOPkM
yfR66X0Xsu0qvpgKFyrK32nuFStaX6EZzU6JIbVGD+r1TsAAzvoFA4vMd9AvAKh5
P75sF6TwTw01XVpyEZgf6w4R70Fvwa33UN7mGuvPEsLDYWqQEF4Aiz+59NNXGJ29
8AZAQAVxVQ6BBPndEkurkwiNEz9AvUp27Q8YMGR6wI4DqMj5tkZrx7DeAZhIqrC7
qRr+I7xzylT+afZ07ZskQd9/V9scWgCGFBSK7duBsdw/pQxwx5R8tgmrQirCn+qg
WB+BrW4BM+PvYY+ptDFsBMNGfiHhd+SAVcoJTkBcLRXB6exHlshncMYpbSVgNK0b
9vEq7aBByGVYkovN2uySbL1s9MdAt+mqad56wGKHDPmBlAzvmPirHKGW+OXkBuc6
KnDOym3OPASllWgQeXvCwHB/EL93PS0zpvavLTtpYQqLcjgu9tTks3VCrWuk07uR
KpEsc/NBlpldL7x60lTchywmvFIuOSMUmC7BuMgCJmSfCN8HjHj/VcbgubYtK9zP
QkTx/5DLsvBSdQetNlpGUWUuomwOj4vY/WJecB9CzUDeb+xIO0uAr0jQI7vvcJ8e
dawmXz035FauAUz7FaLpDTP1iL3Fmlxc44yD9yJ0/7dWK1eGyHkvInFZB4VStRDi
c7ild2PtgCwZZMhaTDXPz+JSOttbJ2yWs1EK7UKPof+eGN6ELkDOjDYPJC9nAKyT
YitB/QD2F5YyGG6Zf6Xnejo0vyBtW2W1vyijjG3VXfIfp+W1GY/ol55swWQ1IG8l
r76BVeTQC22jIsQefWRIjxBk/fUfdNXH7UVfxH6vi5TgGMMi6DQegwBiyh6g7Ixv
thXfLC3rk17h4g9fE1gz0vd2hZyBP7XmbFQPAUDQUpAdt9tmcTpRYyHuIh2+SaKJ
/wP2Cl29LBtw3vxr93yxuNgf3QGmAf4tW1PcSKKHqdbnympjA1+soHlPToKx9+CW
4rrAgSIld9xrp7aERixbtA3MggnXeMP7ov+tdfXWMNAMtlufSW8q0nu50iRXuO5e
t6R2seBQ6FWqLjwpHapDefXt3hkoE9ddZtzPGFf5PMGwywDK09qbqX5yAakbqdXZ
n/uXy+3PsawuA6wELP5c615clGBQpbbRN7UPFCzQNaRS+P1A2bLk+ouRSnxYw0rs
67M2nd/qDMPzDIiF36z+Kt0/tytkKWrOGVA5N6Z3wb4xOd0tPrje9VXg4M51bEwW
gPAo1/zKr7OG9SzloLCvIjfKJ6D9lon2wn4O3ilfK7i/R+cbxK8r0LpMZmk16IYd
0fBbqCLsNuppNCKu9PsKOJyz1+P68qKRr/Q5JtueS9jhi+gJiOG9z7naM6yfeb7Y
30nP99dgXtxKtlhS8MmGT2FDpcUBSnAl+1s9pX/R1jzIr40hdjo91PMzVmRGYKSA
SMaCYYJ2pmUe8sS1oeDOodtsnHNqOEJutQto8YxamHM8Pl8uLc+ZuLKr+m2bQkdN
zOL9viH6hHbPG51NyFfCut2APlgSlXtcmQiSzsCuxlp6PLJ8RTfXA0U3bMjQnR+d
GW4VXunQ0ucpciwaD47fgdNReZTdkxyP8sBEXEJIbCrK/8G0HBTJrpdD3s2zVXVm
lwFGnIis+cpVEVddiB7IIJq+dNfqksDss4Vnpo2hoQjxPs2j38Q6gmppxpL/Lv+a
uePjFFdgF1HIqyIs/hDL8glXuUMm1PgsdIgayQgmy1YvHIi3lsxalEQdhw3MmdK/
VPmLAYr5cuon9zRLxYEUpe+SXXvr0nLOp5hACoM89AdIGXg7jiDaBXGg6vPH1gLt
588lTTSVYstefSOZNr5VjYRVEPgIdLi3juLBiRo/T2A4OLrxX4bO3uqoJu1R/RiJ
cHj8vVp1/eecNIpEacDx9HA9btIaMFLih1rB88ZIhB7FzLaIOZ/rpajT3Jl6fGpG
Dge63vDiSvCVuNt0uc0Uet8Lf6iCt3QdnnX+346R9gvjGQ2MSG7HbgcPz/fqS7x4
Z8iS+crKEwppV77F9HFsRAjGR/GgkH/i5vOTKNgvmgaRNsPVPO3dkKVkZsGorHkx
dDaWJwPasZJu5ZLsDlIBL+ktVJ97Qgqpop7hRAMoIkjC8xrfEfCs8cd4r1MY2/zx
al5mt0m9THhKd9NVEPAql6ad/Y1Pv7+9mYS1S9XWiB94B3yewL3/NUAQdAOaKT7H
GaD0fa7nAJoi8Fe2b4bdJXEO6u6GeUjNQiDaVyTTBsBg4pogXBoreOwTwb1X6liJ
qcpu8XY0sHx36IarWwK1BhILaerelm/Ee9BJo1dQTOIVe9Qph3Qo5QtCiPdIvIyU
2DVw+e0yGZjSQlp6etAt3FHoDasYXCkNptsf1aRxCqGiDGx/kxZRP5FmwLOqnjLT
yP5N+V1VG9jlFWF1F78GhMkatUyOYlxAtK+t9oo700jZf4Y8l7cgNgqv+an0v/I2
qnRh/V2AMYx61V7qSjo4mLvpKsOI05o5sA31Y10lPlG5yVdx5mVr93Rpoj68TwE4
sfS76Bv179yqG7LCgC5unwdJjXGVUA3NuzjlXr3tKZS7WmHcYnbD2bGpRtEZ+jaM
mQ5hfFhUBVSrkscKxzLir6J0OGPDL9jmurXhitwc12iFaULEYhHL19dlhX3uIPuB
aR7a+p97011F7he5pqqpxNOxb1KMvWatNgmwiCSMhe6TjAPPxhCwIv2UKKeetAD4
BWhNCwlkV1BtPcgkMbrHmWTKBJtNUFPQ1nG1shh0AVGtpEB9y/d1flTHcRq/K0oT
3mkmXzxfkBuEMJ7UY804urj4S/GHxNBCX2keO1B+WLRyFa+/D7N1ZzY/94zzG3YY
WLMbHJoWT8GY5CeNlKAFqFpbBbPFKRfgcLgPWZy17qzr2aS0TdSFIIBR5AY9Lzkh
1+fWh5ZE3C0XdEEfsDg7+K2FKaWrH6nuf9fXiDoDk+e9aaoZS8Zhslemk+xgIyMZ
ivkhuqGsmh8mvUksZO8P0njpkee1G6mS1vsgQOH8mg/+In0DtRuCRtXK75hERhWo
0f1d0mcJ2s6yGKEwpEI9PKx5n1Idd+IB9uZB3lBigCtEdLVfovbHOFkFdYLB+SOW
OY12SIj7BXOy93LgesHYf5yWpXQ6etMpgvi8+2GIB3cgjqLx7meXHd4UzSnp4vph
SZzhvR1tuxQgxQOYxj5qGLimILwbL9lfEtrwFkdux4mIw644yDUeaUDL/lWyK3hx
QMBhT4Kx7SKorVGGeCToPrCgk/K+M1b930eHPGOiPQ1oewSKxWC1N00U6exfBDGT
3S5KIh0ankKrTQqvuEPkINp1VTC7vgWidJp0JDrWeHblI9bBmzE0maEnHb9lYmvA
X8mmyosTs+K6Gj0aLwC8UivA9GPUyeXtRQZLxrRs8f8HRyJHA1tmF/Sq24WQ3rHl
zD4HoUXfo4P7TFUw2C6he5a3wPkSlJHArnHalDAKNwVPTg395hItaPo5907GXbRh
EHXO+8M1/Z6lM+dVOaZmAHW+Kbu7dBeA5tIKDj2jKco35QrzmCFpm+teFo1bdWpH
cygjixDWQ41+BqwawVtBqwD/pxVWEZRB1Z89FE5DMfDxxXmkdWbFKwgFE2BPBg8j
eS69l7IPbyVmu94bMTTc4PMydRMVCB53soeXFCjQUNM9djqwl9fjbtePTgPJxrap
Ux2CaNTa9fQlyI3ddZoxuO45J9fBSVquEVM+bt67rexvwdi5XDVdLSk8kZGcluGv
21wmkNPYm54gB2wFFq2Iuaysd3pcTrF81IeTmysFAe1NBxicXBc9DDmiHwyFLQlK
IMcWL1VHClDiNlLamY/GhXHievOpCsKCDZVLkdd3/CCf34NmjrytzwSPDrztgyQx
pOfvS9SQX5uWuQUm3ZJACntc7Z64Xytnt1qgmzmY7qZQx6GJWTIC3Y1iO7JBAc0g
4MMj0SRqRAXfaBdwtlNp8ZAN5xA7e7gYFS/rMTJQ/mwYnpCvxs5aD/93oXX6/nby
OqCwsENtpXIdg2MpIJGNrylwoLSwaEx3u+m3GUfu9IzKxpXYPd0C88t+NQUntezn
GDN+m4bLsRjHwpVyM9HXkRxBorHxKJ1iSPZUVctba2LiNDw9iQH5IR05bzhmQSfq
CuorKFqKGs+x8SyGzLsUfqiZ7dy5N5axvShlp1SaN5bnFT2ObSDn9TiNQrKp/C87
u0E86afE6VAFRm0+8jTs0DTm2UyPiyZRqEYIviEJiA4Q5UC16kW5uF5qr6WdBcx1
N+o0604CISrPr9AqLtBL7ckhUYC1ANYckX9j8tdxBJFtpztEne7tDJ+g1gPzLppe
M4nFoXK1CIIjGxb4efZimN4ywvJQHHDE+NfvxfhixuYb5jSKFQseJiJ09PguwNOw
GFpSDwNmn9IInBJMgikHMTKVPrWUoT/kzO24C9M0ggmVCE8GQ4UMnwsYq7NCsNnW
/JTsep+zrDnpV7O8Gk/Rks+nCcmDFD1i3Ww/1mME1CE0cZuwHgF50jxfJEZF4hbw
mDxNdsE0SNYH/x27u/d2MvtC+5wd8FVp3XJA/nHel3+CKVnl20F3IUb6vnYcucKN
/THFafADkGd8IxfmYqsirrqXWcjhg5ozZywq/0SLBB7n8dI+qiwKUT07OdmnlyRa
bUfZmLKGnC0U/KMGxLtFhbQL5KluGfDKBgwNAMux5QI77JOCYoTde3zQ2/kG0PFq
kQcKsjaY1wh7p50WgjgEno9lTNrkZjavoOqjRT2j25Km1MQfbZyHEDtc2aKQAFst
VhySbldMiLR30B7Vr3WpFc8hQ/YDpiHdmDaMYYc3ej2huik8nY8crM6u7fc7eDz2
hmU9lddp7ihg4nstgYdhsOjS2VR5rIh4wh/8Vy+n3soxZF4FXcHBZs/fG2Xsqnq2
0IPtuQ0TOYnw8FpaYBVPwHv5kaOygdG0JrNLA0pwq3KWzbPJf61s/zkmG782KDXy
a0VpOSKn5w1WPk0vRjifiHXkDcxFGE7I8Tc+HfOYX8dvPIdbm5oN1V1/Izb59ETO
J5FPdwmU+NpMgFKXDkqwwB4VoQ4i/mWTTEDcmCnvEw/MKJJ889sWqPeJJLwr5zIM
kMUJtuHzLZV3l9KK/T4mKgVcdIqs7wxYjJqKroxxiLpaZJcM46/ImcXkQ6glkp4l
BGyxvDYGXe+Mu5ognC3pBy+EvHouA9dwH62pmtJzRyKh/JQ4yv93McGHcJtu4mIf
e1BraBAi009KqgQiF5U1K+jKFAq7h2+79T3lo/oGYVP09j02H9BKWsbYUiE/p3nb
PvjNZDcBCzfKpDtNMbBL/V2Nk42FUBZtumX6li26iWTUHP3GU4Cc7xAbjb1b2foO
CxJY+D+c7FuBFHZoLKbc/1mDS5PyJlyF+vhnM3RRxZ5ORGZe76AiR7I3SjY0qnbN
HF0nIHRsP5ir//YMaId+iAE5lWdpqUUsvp4PJtdJVBMmpN8zh4yN3YvYJik27SNL
ODQy3QtlqDiPJDqsIvsF8fsTcG6ndsMKAv8rv/oEZvOOlA7eaZPiNaL0X/irxjO3
YB7ddKv7tqOqcdNZOUXS02dvuq/v88BQDqGHXA85vT70hauRVh9MSIHeS1lFYFSp
nIzvMK7by2NJ3cDtl8QPYpxH/yQdziHm41cyUtmtDtBqFaKkS4qxk/Od7M3Bb06y
+nkNI8tRfLWIJh4gz89iSBKsV4GV4ZktblM83qpaGiHx9KmXY8lm2QfJs/q65zKe
nx3jfP6ZjHa4GUGsCc39YvICybliZbSYjn/vG/923KViPSlHc/z18jpQFEzZ9fl4
bqjwXU6Bk9I0B2h0XMDjSgob+DzztHm71NmbHlty/xUJYP8qU4TkcOnoWDRCaPIe
L9SxxkKH69SHu35EBEwtooW/s9VLZzIRl2Z2nRJ3uHsEHvlVZ8z31gjtXMUGRvmq
6NnGGEWlXrYLZa6U+zY88rxWWFxTkvAZB6LfC58FqKtea3dbGkTBY4amXKypTJ1c
dTnzqo/ISnR6GxisZJVXGQqMc26UH0AFhszzXZG2VRuZQz62liFqla+uk2gVTto6
dXVQ0d+e7qpcqgmDFdV93M/ZPeGZwiaMxgjsh+Ayj9+BPNWWCDIrCmlvmFuW1mUm
dXE+Q6Aqq0oYFhYL2zvnjxBAYMRTHWpc6yhThmqb66jYpCVwyuL9c7txdA+OSuq8
7MfIk0iGQlHPPXg2h9Lz8D8niyMJBYd3GGla1Hp612u/z0fIklxMpdgXht4zYB70
xms4Cp5Zzq96W0gsgR6mb+4eX/yuey7I3Lr9tUI+3SlqIEL2A+AT4/zgNsJzwFZc
8IXUXGVHQt4oxcLpyI/dPPyAkmudV5DYRye2ESYxbp/xKCBgs8wgZG8eCsVWnDZW
F998p+jX65ZsEPf2kaUE6daCla6OnwUxUypPB46WPcUOkPS16nXrmuwcNNCPRdED
jgF2sbI3OfNbI0aTUvhLPVQ+hjxcFMWu8IBvqsGnn7WxOMZFrXI1wyIH9oMgqSRz
WY0XgUFsk42xKR8/pwg0RzPZOkJQp7V1Nm2QRaTyqPZKManmfu1XFLYxvx3m6Ep7
VtMODGkRDKKzoU/svqCDtU+xxNepqIohzyn3p9+wEd9xiBPnNWiAxC5sBugpWeax
A81tVldlnq/qPGZ8qPUsDvkiAG+xhWQk3nNkusKY7jt3wAWG4x4cLz1O+63jPkjv
hgoy2TFoWqv2nH6IP+aKO3IKuyrBtPD6RTha8fCFEs4ug92YOtjuLl2FjfZPYd6Y
p3kdtwKtX6adR/emM449VnR+NC3VLcsKQ3knlIt+oWNHPiaJzAxwXjI0kHPWsg7/
gfHdS3UAPt/El028eiUs6IVhb7nTfIUmOpHXxqbH6njkdo8WipwsVSd2IW0oHniC
4cVrYgbcAQipavznY3/oTnmOggEzznQ0pVNqCVPTATZaXuMhPfgBRA2WU7FhRibs
Z3NhWEyFamILmsLEModjEdpnIrugpRXwn4NGnmzBSzATTLHstMDASsDX1P4EXS8X
/YahLqjJoA814xi6vHzvGT+ywVjs+81ROBCxf4o4yHUdaUSGxwkiVO+rcPgXAV6x
K9o+aovyVxQZ1gastBFXlGf6hPs1yHXXoeVkNgYvu+CPavPCvVmrHOriufdvAfne
GmU38LT+u+CGAo6UT6EWm6EOEC2rxKOsGzsU8iA11d8PN8TIyB/gaSMz6LhSn2wO
IjaBKvWTaxDoxzp4s1q9+nkllyC2ZxfPO6P0LWj665h1+PYViKKyboUrUkXoh6ec
75PJr+4PjDJ+ZAblWYcmkNjPRl8456VrZ9miUvbYgZK6M0V1AZcjX9yrV+q63qRn
IzQHJITGrOMh7idToB2ibYKwqUSiGe0ORMxTeAv8JLClTNYuAebAVrp9f/xFDEKd
wmCN65Bk5BHchDA2BC2IC4eFYn2gecFhrb3blT7npCXPDS5plW2bMeSzXV962+1X
g7oitDuNjzBDbYBsrXW3sNHjKKAZXJP5KpyK8pzhfeE7Hl0yD7eInfRZ5fhQ5Glo
wsrtSTbagn3vjBS28c2S904QbNn2jBMi4+P2xjwE9BOP+yPRTGjvua/07LsOdIKg
s8BhWakTlv0wyh2YeZXLcdnM2ZYGUs8uXz5DynVHFCPZS1ODLLDUmtpmYYffSn0V
2UCHxZYq0OL4KI9B5+3O+mSNbYZf0U905pFbcqpuzGUOWK/cvlHYbFMKx6SyQH12
Q7IAA5yRXIsliQyBfbGXo9Sslobn7I6i2uh9sPm1oHLD6EPTuP0Y3iIlZ6xz0SSk
442n94PlRO3eLhPFCVe46AmDka0MBlQ2WMUff/I/3Mx4XZfLwJiwXEnNyQVcd6m+
CB9rqUw+e2lIUpxv1lZ4I7qKrTW9z9n/r2CsJwFsEo9UHcpGi4btKufsDeQegOaX
/1JjFcMNscXmqXOGYhY0VJZu2ltcCNIpKW4AldGUD0eQOBjLjDI2jL8bSGU8xxFk
8pOiiFSaS4uodQzSDPSC5hZcWFpJHcNPZbFp3jaL89jh6L0yZzr4IBtksJzuEhW+
n4TQvpWDvE/4kRr7xN6ncjwqlrxLbjROVafxOKWSfxc4pb5Zp7rKNmlB99xkFePe
mFKDhurNpVAZF+9ozA2eDaxNJYRarpw/vfPZ6TQ3/LLbdXKYWZcklrmJtd5/lQLe
XBW+IDl56oMDSfo8+370pAYv69j/y4dsyYNJkiAHxnBv3FhssoXZOf028pgREq1m
o9axzVJDEzvCVczrV+JK88SuZGmKQnOzdf06PiVNciQ3d0QO8IkVUTKQjg5798AO
KZC+W6es3FvD60PEN/eoFy99mZQgQ7yjwtMJA93M25lHsTSDJBGNzpbTYkGxSssE
IYl6mdgOCdBWHTcDuhT/eXkgQz5mIXTvzXuGbcFb2Cfd8cAoWQTNK8wBlqh/joqn
WeqzqPZ1Hq1b6dCbfEzE1LgVIVcE0J3T/LkPDrCq7laOOM1QyGnPfM5yUlOBu0IT
Bq/etc3uukBJ6fI+nfKT7MAcyUsmzblluOVmjJTCMhaupKh5naOINySJpPEKBoBt
knTqXoLnm1S58JM7vJbjveI1FU2EQ+2hu1im5UGtji/Z9r3e94Z8ZfE3PAEz55bp
TmDZzkLZzyUI6G4XBy2nJfLvXHmGWrtBLgews8PYYx//9UcB5vbCk4wsdNDqY6hJ
p/nh1CMwmmrOCK+fUoOBnGropJ1uEHbSzOCbx708DSeE3VU8A9uPbn44BPHdZ1YD
kc9WKSfUqTYw7Ps61b47oySTFK4xA3MP9RK0nzFBuqv83Z5pqajFy5SGXE8JdeHd
qKpSnn4/fHYAXq1RpFIZO/LGL8sBcImbvNiVwvFNspDuP4TQYHpZt4oFwwhUy1X7
LxaXendrCEQS7bMku0yp0NzNVpxN+DbksX7yRpDzpnDB8/vAYxiN+gJ3hNgr3WNu
S1SVdcWLUaQbc61LXQP/4WIahGCUFvBfbOmaOansaCdbKHz1mthmwNEv7jOATztA
3PCiyIWkLKDSrNslr0xkkwrv/siD+ig2lHh+926syyouN3bPe5O0pLU3/wYJ0KMB
hGEJf/PupbYC0/84UFTpozxDvS789eNJ8lRo2bn7otlFGj5T4yJNSaHU7ggVTDiW
wvuQXf+93KE7absjXaaFCgwIeALoxrm3ndTzBIvTbul5PM2AoA3gS9dEWv6By240
N5+2D9SIxLNueBHrRwabUKR4pDW6of7vyD/VbA7r6HMU99covUzVplGdlPTA/yvc
uHpK3CLQCP5rii/nwv71PcJ9gWykWXxgbQJRene0y9W5al+hf5qRknwIDtKHJsVz
+OsgnBfqLGyttatLFOYQbYm+DZVjG3Chy+srasGZY81eKmbHgb2N8c96hZkFcBLQ
FbRPooyWK+AvBVe8/W/+A/oqk9nfi7tUN2LqGBbF64fpbUSHoOERvFQzIvKUu3Iv
XxhoQlaxnyk0bwy+rYaZOEGxlp/WNrZYbAz1yuUsrMfUzwdxu+F5NrMvOuZbnXoH
XVPz0OJjv2vnMNs9nootunL9L3mcCHwyDly/D3cckgwpc2I59yU5E9ZExqQ5TGlN
tnHbKYn6XKrcE8qwtSoIiAmwKR5r67BJTzhA+LPDQuVyJPwcQVf6rVQFE/HwVsZw
F/rp6/QJyhe6Fz89JW5EhT2lBNTTPY1EdF7U1KwkPu734yQTbiB/Wm2WuUHs0JGQ
lDyMYXttfZcg/TDTZ4QZ0mDvkFcwj+Puj6OQOA7dPmW3BNmZak3x7j5JRFMQawaC
B3dRe8a+cyhVTPkIgbRT6UGzkKLuUUeDlLmEleE783Cr1Gb7TeIjhlv2l4Vsv3JC
iJ2ufZmIbKC39lDXsj3n/oDp2d38xRdBsOcI65ZdcoVfI2JL2W12GneRuvmt81wk
zzMQ97eBzxbh9zawJDTs+UVuEhq+sk8Ui5e0YCLofUEGCIp3UUWfyY5j52oiDhGE
FjzZF0vD7/YmRIMBwLylhGlovutp5XhMWI+ieSfBoOAWbH4E4xR0/bYYsWfpAs3B
sLyCep3WVm3eWIHORyck49IpPDZZ13PjslsTQgh3CIlqsjj2yGQjaDou1hHymbZX
GGXDPbpHuKbJUnqljb/FMdluFrIUtXxPM7881yhD7/t0RGsB00qkV+M6+qR6rEJg
u/ByI6ysXpK4lNIqGJfdzM9oXVa1JfECWidtwy+KpvcBK2GamIa/UUNZCF3Vvxx8
n5N9gv3q6en5lwtsrsGVgLaEwVImQRYy9jUXjAfd3p93GqHLF2OcHIzZzuF0X7FL
mApkpNEm/xx8FVAAeYDfCORp5vcUsQmSIxbi6/vEZcB6NFOmFMImyvHwon7E+M18
SVF8koUW9dB+iKA6CxqSsIfwYdHn3Cuf+iFg7kNedvqJsO/CVGVML5kYA/wIpRVE
fxKEB1YXBk2PH6YqsA5/gWdn7SYq/5tgtCNxSImWpduEck5t6yIfv0InaJAfTmYk
oop+QWGeKgNJ9jO19UjZ55Y108B7i3E/xQI5ktwOgWdS2a24x7ktmXssGysSP323
NJeBVddraWe2smyGT9ylN5Aiq5pe3ozE9Kku/l7y6jge+k8UX6Ov7I3wmmb2NNve
4m6rfCpXM2P4RIQgTgs8i4Dc0l5LpV60Me1y2uN00X3WUu8NHzECBVOIaCtJzj/g
+6iwncJ4zqVG8fOPj+zzaM8wC1cfEtz5yoaOr5XwP6eoRozWEO97/ExqATq3rYZg
/PchuA+eH6XJJS3nfQUyLVyd9SECdAFZv7F6OYbmP9ugZ32t1jPvvHhqwjy7vqRj
Kjo/Cg1CuhMvDx4DRRWcdGjl24XPoMeb9VeuPBvkNy2YjGKLWepJEKYjFSWggf4G
n60rhKQx90sk0Hs4N9dIUoPeq0m7GruHo9hLbyn5tkWmWsF9qUxVokdKXsE7k6Tl
0r3JF9LIgW9dIX/bgSs/aIM4Hif9B7raCe83cT9e++hhPgVcc2jiK2qTYtxuz4VA
iE8fO96wAYBWzX8gFkr/kTE3czcJlRN4gJv2VEaprjjTh7lkgDgagK/6phjzHxZO
n2iDEzhFsBeMK1xfx6jwvyQ/nmYn7ue99592K/QzvK7z8fyC6MDygBZsMCOq9fyF
ZBXmHBsU+xQFxj+g1lw6SVEIPJDy41wXViJ3+9RRoV/vBWuLFX600pbKrrOhR2H7
xA0iWk9U9I2pAt2R8Qhq2BdPI/Vzk783BMxmS+OngCiEwC4xcFK5Oy2gomLaWokA
6VAV9CAeSKNqpi4ntleoS0MNCQ1enIQhvz7GB5F4B9D1tm0SA2+QSxq5HIduSJZc
9fk6TwNAaQvWmRNM7Yo8YvRzszUfx+EXtqrD4qwj9Iu6DrBc/0getJV86nmsQmHu
rooARLDSILxEo6xzXIfdL/kbcuOjYaiuhvMOuLwemKAzxIYvbMpmLT5A+YeTTp9I
3xX4CXhZkkGl7+dsgmbYPh6tRaCzFw9p+3PM6YHpEca8bmIB3xDB0QF/shdjalbr
wo7saRhh5LACUpCNVZHy8OR9aj0zV1pyEOb9ooMHU/KtEkYqT/OPAVkWLAL0Dm1X
Mz3g98L++Qfd3nwUmKv9VPiaU5PWcJPui0ULO+GlPEnAkCzh7MaBkmPqMHXV4POF
kREudtTErn0wxOnaM0uYAocIJIiT5rReKVdyWgZdd6slBedC7jWJuh0lFYx6FCD2
UcXGd6EoYji3M3x968bwvHGPg+ICEyHS9ksJPWkbbf01LYwR11OlLfu2nQjUDfz3
kBlFBoCB4wdtH3sjOfw5vJ0mEfEz8fuYRu2dzgf2gT/VZOMvhrDkxFtMxNUiUQpg
dBmispBNbW1RYIJFxc8OCUZkcD7VQqsMl071YpuzE8SjBRByfKFvTiL3LUmQdHyQ
gz8yPqr0X6JBEv/XWw7Mq8XrRR4FEOVVNu/yuH+ub6CCvBf7mYD7MGrJCYLZfSKS
XX6iQys3ZoqypoZZtksTwfmPPEn5xEsTK85+j1fKpR71BenrJBOo/P1dGdJugDmR
kd8zA1sa1sBT9ZksFE2sA8Lqu1RGcPS+hg2J45TyonqZsPn2LL8vp9ix4zZrz8ch
Uo3mNxdyN2EcWCsBO03UWDnLjbpl1wy6bd5Ra4zDcA5lv0Ddi8+4UeWaW3Y2Zslw
sPfc85X5KVvDXy5hoLzJzVUf7UK7dcoqeuC7wa5rz3gM2Gt7aUx/lUdnUMHoyGG8
plaH4xr4fsoBGJGQSxatw0wzYDit0WaXtJC+wBQIBJpHMVHpFMeqMpYPV1xdZwSe
uCBp0ijoPfDONOnWafyy6aIsTSi0UZbU2woNw5jHe8/iceXCWZiR9gjVyajMoBFF
/XSpUU3V6YONOMGmxntPlwUG5VFpzmTo/ITMuiE+NY8e/PHj4AJlEKs0Zdcjsblm
y938F28v9eYSB6SO/vNWsf0L5UuyFZRnsZXSevgW13+EJMNHRFRBTEdJr7RZ50fN
pVnDV0TPfslGdtqAktd+3Z57ZBu5hEf3/+JXS36MW32E1Sh1LB0qf2AiR1BbwVGI
6ApKkYpjDNFYAKA9KzjHdp68ZI+LKcxVhyX8vnS8h0Ez/5BAY9NiRX0i8sQZvbdM
89Hbberw1MOL201gQuhsQgB3C6dvd2uj9dNJ9kEJFiGUn6c9EmaztnW+fQT0yMaq
caq8wOlWzFiEceD8OQJ8yld1FgdSnICVplAEVHT6KN8ynQkyiDpEYoA3vdIgqwmi
t5BApDWmgMHoUBbfIRqYbstGbKmjwnWtZkX4IGeYnGthZWxz1D9dLqqTzLnzYIMV
cehfD3lqVKhMS92/EHXriSvUFrvVvXbz7TMZsyVAlm4iWJK8MQjI8G2kQDUL8YaI
8//cga+rK6CtvW7Ngm/8bqdWQTT61Njk/FMbXLi9Regn6Q8q2Jtl5KVufSbvG3h9
AoZhMkLURDr8fD9+2kOdiiLvRbhzijcqjln8UGFVlduB16gq/Nt8L4GFB8N5hPE/
95hTTAfIAVU9LVRhGrfk3AfudL7CfKnImnrcmg+BqvdlslkFCSScTmy+UnAQF3x2
N/36nfIz4zhrigz2WK7+wLzFWEnyDE9TgybvnbdIomDHHtRj4TQ/me6+gbeycGC1
DJv0ZL8W466d3bVKc6w8poiG/zzI+RQ6K56w6bTbC2cO06UgVLUaniuQP1cgPGQ8
HEBQJLtG/F/TczkXwY1fFWWSVNLD/QIjP68+t9AmCvN09JAT7SbYT2mHIqpoCE9d
WaDdvJj6GWE9cT3rA6V80PpTqrXUqWHuCRYnxt4OtMDkyGbNVMWTevlVOoWstq5c
d73/dn2wit9r9KbOeYxAeJ96AnO9+P91aPLNc8C720vZpO4MY6/7pgmNjwlGADhH
xHENaLRFGG/9eOe2Un85LQZIQLV3sUemvxVBu6n1RXJzASoaazsBG9W06ixbXK5E
LVyznNswFI/GmuZDk4fMxieCkP+5al6mrWfS527WRQn632o1FHQxJBGfZIHKwTQr
kDhJMVC1aw8qHDO1GbTeXdi/M53PuJdMVSdq8KaN/clMz3Fo2LNGPaKM2/f/kG99
EcfkYoDCT4r0mk6c+X29ssfHykd8qWgzyJ0kWShHu6wcztg6baGyqr4noRSnInVc
pt7T4EF8ttMpFbJHykP1s8VbRnmWsur3hudIYZKeHa6XdEelGZtFEi87HAyv3NOS
nok4kH6f/x6UN0vaL4Fzhewi4sp9HgZPBBcMTy3DfTFbHWJ6ol17+W/N4c7+nNTS
h/1XLljcASf+P1K7QhJaP6XlRoaCciuYj+/xnPIklkzHmgAJYZy+4e0hYyxLu+69
64KOFUYUcyxMJL52AeOS0yIJnD76bhv8FxmSBiDccVaF/3YfiVyIoWWgkkpghOm9
qrG4Wu6eR9KP5BXXwbiEEYsMkC/Qp864O/lB04q/Ljuve+gXIDfBQ/QeWvoyeSLq
kiNVUR5PLMOmzbkqMLz3hiihl46nbTgNQVtr0StGTFCxBAXRRoW+NW7z5xmDUiw6
vVZjjO+JPEeCbH5/6gLC80cXgl9tPjJ1/KpZIgB39LLwgjElRNE/RHydUs4k/M8M
EVxNgmVxnom80L5b4yWN025Vpohzk7oFtyNOS3bP/MUZU06eQpkcyEN3IikNxLFK
aO0GUIkunsxp7R3NKeuySTpAlgMG5w3EP34kUzT0ArwvfqgZtGhmrWTwV9ZX11f0
b+XUbsNoBJxmz8Vl4dNuRwOw9aueWIVlb6P6KCMEnJFKyVAvVug7JBLHKIqUrHEJ
gqm0iG3cqDObhEFQmutd1TnXg0nkDj86dRh2xJXxgA/G9FOkX9lm95w0ynau5PuA
9pKItZuhwbhtpJ5U8Pk1Y3a1EUTEvLf4jN7y9cHTA96wNasucPl0+qcqQPtXCzdz
+gWO79xw+wRKOMABGclxfXIRattCsggTkwlMOdW5UZVaZ00f9PC4IqvBf2AtHvgz
9Hq9r0r1N4CgF+ieP1ebeTCK+wAKUk7Cf+pEKc6YKCLWBMWzE+LrT6621OjUw+CQ
JjC/PJQ1Bsx7+tLVWrKGkgsOJ6E3r9oObWX7Ur5ZzhjNnYHSCHIbbrzRDrySBpSe
q/RneJA316CF3AtCvCI9gQDE3xMRAJ9Ckc4GCOiFjqrDN+jIVUzIkNIc1B7gu5S/
+TgUCQprcLVetCSBx/JosLsWyV3OtBdl2/EbdWjo89js+bxp8QnRRG1Vp4xT1lD1
uuAxFDbzVMQU6xRCi73IGtIInJh4I9GsMLWOmN006AtWL4FRk6j0z87wt790wYf8
uOgk9TGKxui/3Pvp3xM0NoohSfbxnt9JSJKYo/OawIwm7v53AaLaory9ugWXEZx6
pcizGbixJqO5/qefnQamaYYDAjDrr/Axj+nmVzVYS+l280GOcDl0Y/r3AOGSs1mC
ozvm7V+JN3tDZYd7QuTr4SRXD8Vlj5ICtI3BhQYiN3t8uprg+tcUQWrJkZED8E1F
BtKzsqjYFkKUapflcVgnJXS7Xdh0b1JZawGijkS58plDqCImJjKWg+x5cIESToxS
WBQzC9PosbkCu3pwzdWCDH5EdHmrQ5bxcI9/vhOyK4O8hQkI92PfLM1Gc8aN3IJp
1YuWKlW+D9pMNRQ8MLyCHZDZNhxX7q4iT/wLc9OU3W4gWvW0+p5Ef2T+3nkQA4/5
QD566cou4kE26UJtpsFuQTIcrHHEXsyoucavesVWMG75dr//bCugQToerNblg4qC
niqGUVmlKerQLvVCpnyg8n9pLBRBeKYgMCdLbfN+BP71uUJye7eBKHKgUyltMKzP
yXdVjufJzBRNFoObSAKDfyK2EjU6ZoIJQcfNIOCmIPjTOLupy7eFF2ktHuXtsAkP
jbRFt+qXQ65Ok5A3WopE2LKbU5qBYOOGemP9OASlhwpQXkcOtVUDLiojafAxD2WQ
/saZr63tffL4DWouh8sK+yR1cjMskEgK5to8d2wT1uXFKzvVnYBbT8NCRN9Pm+v3
0AEMjmkdTbwjDLHCmS3Q3CBCE7/o3snpAtkfh6ITD0RNPxE7Nwhhikl6XbZyoKmj
EkJbZ9ES4yiwB+yRxTRbzD3GVBAiMlRhNN6W/IU3Z9i14mfqdFSOf381KLdAB9Zu
UVy2yycHxhGjLfCPmYcmWeGQhRLpe1S8PMpTCcI6v67AoZsX0aWQk9vf7yjqLN79
Ueae3ebp4AXusUqworVHqwGQI0pjBJ0XJoS05sGoXS1/4WFaRwOZC8RYuH6RlGTr
DxzOYpkxoHIy5bm7CqqKJbdb7BarF6rLqMC6PbPsiyPTOod631m56WrCdcB9llsR
NFfPQXzgrvuTMWFd4Ar8rLAbUg8fXcIdMA/Wcugldi1lG/j/j1ocXO4zW+8ICOY8
ztmaaZ3kf0oBKnWf4ox5iHT1mIuFDgltjmnAfRu+IlTLRi0DXS0cK/5JR9mJ7ML/
RjXIJ2x4LVIIfZBOOXZISBDADTclbCg6x1C0YmEHUH8UQk+nQx4DeG8GW83ezSXo
WyOwY3zeYRINkslfSIz92QxxKAVyFRHRHA4VPFYBZS+Zs7ViuFEjiVJXgi+AhKzu
LBEfIyXaNSOfyipbkaPwgVO7R2gpOCFG4kQM1VFJxIxA8x+CTfHZIqSQewvQ8bQH
vDNY+IRAs+K49DAo6iix1Rl2h9jrIrEnCeRtcFTgC8i8ljSH59DNyArj/ZVQmlI3
GxJMe+unG1LNe1brGDo36JgI6p9levCvMc9Y3Woz70tdKqFT+nlqRznrYxqhPhqd
QRkFOQg1Zi7KylwdNtR2njw3C9rgNydYzsF0GyasmCEKDDEw2put9rRi8p/LRU6D
R6/vfBFhLgBZ83YPVbteXAx3mzR3chpPBGH/4gpDWa3Pe/u1izAWspXQFW6v9CSo
6dfuBIZRyCVeSHWyWjA6HhyWC3XfwCuBXMf4/xfn+DCsn+CC4Aj0xIoR5boV7BRt
W5S8NceE9b5xF5Iv6UXTe4dXK+7fjtLf6+r4dYPvL/FkZjp10HMhMUtlZ3GztgKn
BaYsmyuOLEiXoSkDh09YCEQYdSat7vsiUuitLdIbqQr3Eg9jB7fcR9/5LJz1uclv
tDPq4u6uIjSqUslGVQHd+jj4C9Xr1ts0AOqP0E3UBWytE5S/jPG2bGF5n9HhtvLT
42hnyHsC0D+cMfzC28zkFiDUPsTzWuSP0pNBTm0R3x1oHT+SXCH8NofUp+cK7Hfj
xoMKwVhQT9JsoHsJT2p3tZbyOsRHnE9ibp5Y05oNEhw98nsAlskqTlM8Kknwz6dT
tuQYLoo6amAjWm2y3YaiK3HpiNYt0wXCeQuXEiNE51lRQkHoETUmAk1+XHzbzLQd
1D7xkLg+PWrbKz7BeqKBOnklJ2xvzhpDl4Nydq5tP/BBcwtxUJw4Q1qwWncjj1FZ
325hq4r1tGJg+fSApfGoxEGTpob2wjFEEfk4Brim4JDbOPeHEZcIZxKBWn98SNjD
IuAQ5rX8ynheZcaiQ1Me3qyWINaxYYyx7LsKFtX7jhsfFH3A8Rl1d0lQXiaLQ818
RCVNXkGaOUC7R0Xdb2oyFHyX0J/ecJuz8FVHhWHhuP8xQZj+YSInEyZjxU6NVI8e
1M5W25OLsLZiP+MFVv0Eydf9tYVs5MOidHzP2yanQccrY9cwJcc4WfQNXBQ34UHz
9JkAgdpI38DW7HksfnbUcFpo/tXRb6WwKJBydTQFwpKh3cEDTykwzH+LIHJRO0AW
QjOnA7FQpewqs6j0uypH/HCuZBSo+/TUodzeVzhA6fQfnLN8h35jk07d9iklnO2T
/azMqPlcEVsKoENXPcMjolFnzUAFx5DhGkc8yx+Wj5n6bf4VDso59jZEP1REvimg
RzlkL9mQze8lyvzzjU6aedt7msZPRFT+h+030kf15y79/SXSVr/VhTUv8gqrELYp
T5GdYYIIDkN7WS66Ortbld91OV4ChMzouEkqY1hL6EPiv44jtJlslcnJWpLx1O8n
IP51EbvttzoqGi54EJfdAH4hfW3XoHsmmaNvFQf/WMX6nkpluWatNC+nDSH9v49n
IygpQJOJGYhJquGkBKNApSutDd7UBzemBRQRVbYCva8ufRoEuo8Ykf4VqkzcqFC1
GwkFARdyI0Ug1KDrj7cKRyzG+KZN06CZjwwmzvz7jj5DD5zwygcq4BJ34FIoQy79
UOdUVAM8p7RPwu/L4Hu9SlrpnmbcMjmOsQFu6tB9cuT+QLthAT2lFG4VyePvrqi1
Bcg9AoXsgZUB0aPZKhtdckzFWhUR3YzleILKyTKI8XKC8PGivsQHh0ttaXufvY9H
oBGbd6EQcSWCZVSfWvvr6HQx94Hs3YQjoHC6gQu+kMxFDu1w8Nv6Tp63kTS5Qqfy
O8fiKvKRO/O6RF4R3UohfltzENjUkg7vLjtlhCj8aYdA/BuuS3HSR5rvzFA6TmHE
kNVS9dwXJ3ThffEPujpDY/R/jtBLNglZdBHdbfC1BxcKjWGXi5z1KqQYkuL/w21Q
GxUT2ZKLM90FUMxgvLlP8QaWaVGmrWsCOpVHjiXMtHbPk8N35MBJvCbEwZqPRJXk
zFJNoQ4upl9IQTwMD12T101jPYryzOWGPugCX4eDAeGcsKXbt69shu8SvGimJTBa
7nqdBrO0zs0mPPLDz9PMkpwYiybQHTPIPRedm2uTPPSZFmxF9Bzb8OSl25EOEugu
pcBw0g+WhtDlbwPW5OThe5XwRE6V8kyWVlPuINt81aRhfpvl9ER8AD+1DLwpM0e2
fVBZeEz1wpGQaic5WAleAPngJG4v9CYocG7+FrDTtA5cvU3otXNcfQAbQSXjfoTY
QqJRGTs2k7rLlyX088Rp/RnlYRgVTw9HI7A6B+/kQQZJwngOUhpnI6ENgI1ZEoLn
fB92LpPJtIqlDOCtJZRdk5BZeoirneJ1cL4A7Hkgj7ivk713hIaaqZWnwOjGAolc
Ao0c585NiIQmLmNrwyfznkzahs4sDkLYjPXBY/bnkQR9U/bMqfbdlEaa1GZGzykA
BzXN6GOdUZQEqjpwtDDGup02vKr3eTai9c+WkUubio6UpQZGD69L6wWSQ2C2aJnK
zF4BhwbILkYsp3lampw9YzZnTNWp+XUqp9L8PDpIbMSE+9zMEfZJyEBDZVENPbkw
6ONogETOrRqUECQjUQ7dfvDzrl8Y0J0O59OQ7UfYd7pjAvQnQer2PU3+I8PPUZqF
Ubvt/ixECC26A6KTdNgplLxJLEDTqmVAnimGBmSGgcIuU29RYpAlN1wDzUWsQy37
DWAiO3BoQmcO6hrheqxCc0SPdJMXLTsTBYP0FG7YEfXZFHfZ+Ws20NlRuGUDVlc5
PBbUxijWVGXEKiXgXOdZdKRL4JpwQFbpLqpw+qi8+QcCU8Wwgx4w9ZMzPDRFp+5v
PZf13S5ydQMYGn2RsJOltUfJoSvcyX6slEaD14jtwQwJ4es1vKB/3CJreEu+rIyW
FtOHhQ+6e2ZkbpyqExBFnhw+k8BJMiEp2vlQcwAE4YyMZSHpw7zVQnHJmit0XIqu
SuTJSmZ++XMpryjMZpmdrlIwbRAspp26O8O6nM6UGCTljF6bDr3aP3ugNwePi+dl
NM4xkfM8ErJv0Gsl6jENrAV8Xd8O9nl+c1Y1oEgQ4BnRofz6LbiFyuY5eUwKsZWf
pFHdU2Btnxew3ytebDA3P8pid9iyoCIh9vDPp3hiuZJmGgF1T52b5As/cHd+G6WI
HpgA7nOHYL6yVsHIjGxglMDMYN1qqqDFzM9lZzTgQUMfkrmmDF4i/hFoXQ/OYgDA
GXv2yeCEaFtFSs59Dj/o74AmTu9Cmo5lG3helR119y0Cx8u+nENbIisHQJ+rlAc8
iqcBV9fUs8y7j4TTOn0gkfHFMPfOXnhzwl/4LLvfEAYvBMiOBivyv9qu8V+xrPCK
sq9ziINxAuZI7LFnZX8XhWo3vWVADcomVaiqSKJLW3u4Q1gMMpAaoX967mIxq1Zj
VosjOIfdENW1SzPPNrTpBUsVshUsmbrWZXqNwQNS8JYULPHIHl3pPbfk2ujKh5ao
/hARMtEbXmTOLjnLzSAORH9RiGsSA5Tohwp5w/7zFquXR67dhHqgVEyPsavU7jQF
pM1bn4DFQDnG5XlCfSb0Nr+66f7wTVRCckGhKUQ3YgEf0jS7t/GycGIU8zGdYI4B
M+8kj49PllFV3joNhQzPZ4xWOAX42CtEY2Ocmp8Ox4kFadWeWHoZkc8b9bBbQ+X4
DFTJUiqyu5Rk6/w2gSAupxcDNBUW+ur04j99O55algzjvdFF4aIG/HU56VCZ4yrN
+2Eh7b3UwsW28bQC7Q80OtHIpvZ0jT5B3p6QddrPvG3S+P/J6B6mxVwL5n/oDZvU
qFZeEN+fpYg+IPyg2Z64P4/WJ9/DrQMpCjBx5SWMC5swoExya2M980P63+uGHUVA
w4CgK7ey5vwHJn/EfK28r8Xrvj1XjHrCMTtEpRn/diSOuOCMy6mUNQ4ds1r08XmK
K0L7vFt8TLeS9MfXCdl2Qqe36kbuTsEcs8DBZLfZLxAKkfkvcWK36vBn8jcJlegs
DfhTKWiEWOhXdellTV12VLOGp99uC30wW7Qtvcmu2jxW0fxxlhaB+9DDp0/VSPQU
5fWOyr8E1bCIC0rw1pt+EWSGFnYVsRNRv28zukICppE+wdrHu0Lz52Kt7/1PxjYs
kAm48jx7DuyW2Oc7DqanZ/Q3OoOTyTaXHRF0LY50ybKycyucv23KjuOTSKadfIAC
wJotCSP7tU6OH03tIAi9jCI2yULtnzoTBu18TARhIdMNrfIS8gEYIiAprGPceKWu
wrU1hE5Z+xWDGNjrgxLlAzcE1DQ8yVpROiV0DnCLbYa16U6xZZbfypCwFw7uYnBa
ifXLHINUzXCoHXtsstUeguSb3e/XrbYaovxdOeSDZUVRimDHXi7yX8k9ps5Iq0gz
nOHaH5sIqXH0wDvqJzSvHaf2UAKupiCl7TWTfopfmdTK1bv7IkHjtA/+2ritIw90
3iAcrEoVFQgy16oiUit4Zl19xnS+hyrTYXR6W4rQTSECZnj60xV9GCq4CUgZrJX6
tXH0VmF8LeaqomdEevWiw72LHndVfMt3+XoDUgkmoEZlEpcBpngLzD2t36SRwRH0
Ga31q5iXJnp7gMsh+LuXF5wcZ6P/09rnMF9q89wLjOD9QtKzETOuSPI0eGgKgSv0
cnhMaiDb5+RhIGNt9o3urA8yHXj109QYQGJ5OCeEQBuyUvD5fz78YJou/sr5IeId
YMbd0gBbjQa4b3LReCIt/TDQO/2y8+fJw6JdVk4p5oSw1CTv67/fJcBkDTLKrKdw
WBOvHlFPBlkpdX0+taW6kOFgF2sHam1FIVz2NkaksRf3mI8IWge6ATNIsX+/67AB
0TKEhGIfsFlwejdooEOZ03uh5a/ZpeFemExnww60EdX9WZCw4RkOpyYqqMRwP4HT
V42LqOUH6lAAsWgLvOS6jg9+vZrk39tLTgajaFZxVo0WhZcVPJ4lD+4M+LMX/emK
t0k5CEhBeCcTDqNC6XAOYg6sXPdTYqqCU4TSjIiddJLWvlhnNJtk1JmoDiWse4wQ
m9THqf4OoClF30jSnJYzlOmLa3HovTAtBomIJ6dtnyJWJQpQ0pV8LI9YBNPykgu2
wUbRbieFjGlFBEOmujU20gmqCfy+AcW0KvfmBaCQFU43PdKnE0dVEiOehpA7o+ky
VkT+6gefq6bQ3ZDTw+RcGnvL/mbPnrJoeh5ZVF2n4hNYyuKCNIB2D9eq61M5l0Nh
KMf8jbIbuGBO2lQlFsegS0kFEblxyJO6HYFosqaLovIS5t3gnqubq3NC3VmxlWSk
TTWdnnIqdR+dywK4J/mvbIlu93GvJ+RENUz7PgRLgTVUZGkAxMZXWu+XYIA35mgz
G+2FMV9z67abZmTPWvELJ6A3Q/lEcRWQ2ejPRlQ8MYZ9mkUYfviJkksilGZAm6Rf
IiwbVEXoTjaVXc+UGPF7A57LnzPVM2NPlp3BdfOYRb/QjQXFgXxvHr6ucUJz04a4
rpZTfRS/wTyPqU6FYt/z6fZDwaiWEVhJ866VurX3RrvIXgZ0bJbZPihjXq9lptHV
gAcEcoTDtXymPKHRJ2Mt6FTFlt4Aq5MAj752W6k9NM9IJjouNO9LorldL7eZXj3H
ghMGDuKLUg7KLkW7I9CEdoAG06OX50hPtNGkPEBCY9al8oNyU59gz6HjpFU/7mo3
TlTXABO3LGp3XOY+fmiA9w7U/+AO+aAvuNWJOLxPgDVz09OZoWMP5N3dJgCiM8o6
g+dHgKssEphqEasFHJHRm3SGhCb8HSxYb6lbtRZFsCXgvOdSCGUAOe9J9QtpETo3
DFEi+SgTyxqrhwwMeVPZFJ864FoRrYhEubGsBaWKBS5Gkuo3H0UyShB91+RUp66D
6bC0zkSYPF2izxQC27wmqYEhLBSAgG7QgJvW5XyMEOEnkoo2rYrktfuMsxczFxhQ
io0/RdtnmU1+kaBvxezpfDAn4fvWZT6f3/S0yDU86vpMqUsQ2RWQ9my6PXgxnbIv
7Q/3N+Ofh5A1Fdg5YAe3wVsAdYh17ZbpeO9d3W/gHiGDhtSWNGkY232h4W+f3qX9
/+DiWQehkftlwy1Y9DteoyX7kSqPT/ya+gd+0M+afXKiJCKQ+Pv4TjO/ylk+TPSg
eHz3ikaTmWlohk1fi9atF/GEtUdUcDs1tkyP0n133c1Tpe0AC7C3feRQkKgE9Mpz
nnW94EtnRiNNlvi17+t/afM1455JN1LTFL8Px+PI2ceb3ZXICw4wTmv7cEFSiwiG
qzDcDy/LwWMLgrxAF7C5cf54ivkalCJ698VfKfsfo5+j+zo3I3UezAZbXkwM3En6
Wn0dvBUxbBZS4RfVHlyI1BGCQfJ1beeE/SYRIiADX8NDLEn2k6h+jMhu7Lhm3BsI
x21ZNUDYZVaBCTyf1/EVpyT6reZcWbJtAtvMhlUFyRSGdUpyx9oM+TBA7DmE4pN3
GfGTRujnxi6eb3wAXGnTEB04yXHpq9WdSrH8w4NOqhBbpYX6Vp4mYM8IIwUJi/W9
5sT5wRBUaROQg4ySZUD45HcYvPp3QBSEQQ6jZgSyEzzJM/eyAIPSfBJm3v4kiwgO
m5cFBK1ZSTs8Vj0Ggf12Cy1vqGxMYERPinT55dHGsv4SecTkCBZsKj59u86KC9Gu
7pxroFxo89iTmKXZZjcTHReVNXivLZbuKiqxoomFeKzNTxGV7MkEqt+58guUR/GX
Vks3C89WekcSJz6G+Bt6eUXz77mTaJNd4F2peIZRg5xe6EXnYYJthUAb9izim6uk
xkHYOBF/W+VQFFdNGEsGEFUJlS0PjgC8HZAlPwRsAOEWQ5MzuxsgxUZ3EI4/P7vg
Y4XXxTDyJfXjg48gdxGoeqyExxxvcRposmjNM+iFq5S1USpmrEWLX0ZOGWaEObS7
0+6QIsDzYLnFyF70xrq8OTUk/rBpDdPDh0bdIiSt0GuUnKxz/ui+2DbNGojSxOK4
IN1DhhcShmy3ajWNzWPB/H/JYR4O2JrAtCuIeM7Xqdmebmgqb7dikqirEXaeTKs6
tLzm+mHV4NSIQYb4L3kzMB5FnPDuss9DP3BEruiI3CL0SwIeB5fgeo4YUl7S9NVb
Vt8cVGV4KLAzs1xZbKwaujkKJmiOVjaKpM+JIAuOJQrQ7NpVlwjOzDwqhU8Em7b5
ooWZMzSObT8x1tzoiPGDrNyAx/ETWdaS95k+wcB8ENCKD/OphTN9+ndPCGMMGpNn
FSvidtrqZgeKxPwF3dEnbVBPuwbOl4Nl3MfM2RNyjKLDy8VFcrA3guI6M3BRyokx
/axlVnCrkxieNecN1ZT3wRuCE5NBd8l8P0QBTEMVJQwZejkOvQHkMx2/1KiVeoyw
fbfYHRZd3ADkLE/Outu5MsyaXqYg3VvBQH8n9FconWENUYCTK0Oex5FTqiIBd032
J9CY5dTmkJnKVZJW3V29gsfyYmLV1GEaT66s9ujXmjHuo4tKxrFjJuwQs1/Qnaqr
AVGpPRklsJWOFDiOuRXE3fPVgUV4iKfQsNsYVwGdFWNSfKYZdDq8OOPn/74S20lS
cf21Z78Nn2BJeA60t1TQkYQJdUzt86DOZ20vIiXzo5wgiJaTkyPRqbLmt9SJM3oL
APbUftpVZaM+YUG4KiVQzFPds/vKlZH5jA0I41wgA8V8NQm3T6HEmlPmJB55MbMy
oEXDRsD0aSLGuX5tmMXxD34Uo907sfSmwpzb+Pou3SJXvIFvfJYrnHb6bDcRixXl
6KDUzWQavWa4JaYoNHMIs1tqdQKhqginumwTzozB/vcSuNfCj+bUwPYOTQjdtK97
kLMpXGl++N/K/6C2FBukLPqCvx6Yf3BlqLWPfkoC2iI4eCPouNWLPWwu7eK8DLeb
wTOYzZwcw7g2P38T8gc20Lv5w3z3SWAODKTXDNRN6CU8Fn2RC0EyInDoxwoaPBJp
2qh0IWYQrICwFWWMCZNZdecmEdhqLauygqD85RhXq/a22kWhvblKbRbiP41hlEu1
miRCbbbPfsx7vlv7eChVw32ZRaoJvQonObjzrP65/DMK3+W3m4bT+VFH3tG2qM8r
CAI5QJYwKdGxDL1hqb6K7Pq0bGKRPYSgwbL76KJXe2Qfb+4vf2L3YPyHZWm98EYl
QczMgCN1VDpMafaDkIKRHZZAFjYMEFk6fGHvtL4SwI1oCYDcmr+1h8fkdc31UQpj
EMIyxPl9u8A3K3M2MwxO8oxkO/B1WdcFA+1upqaPRA1dpI0TULhkC2JGAladihEp
t2nquG5YbqrdBxND0hjOp2TOb9lr01fk+Rdl+jysGOSe8B+waOxd6k7wWkCD61El
5pBgchAko0ZdK9PdTI+PnFpffLvq9Hm1Jo8DHhlYkAnWjQUVt1GrSfMlCXFJwja5
8TlRtPXNbhSi4CFW/o/34DIwis3dDtIafL8YiJNVvG+lRQQgbbqc1/jPpn4UGplD
4sf6Z7s7sg7amo23RUX3G5vCNr53iP1C0oxKyiHEoFKBPPezbiJN31y+vxg6QFI1
xfmPRhMG26VjL3t1KWHLgRTplnFxYoHXrwar5B09JehEauhkxdjnclxD9cKkyR6J
FqTmCML+wOS7wMnx7jYhojdi7Zsm4Ba61iQLWCuY9gPGjvaApaqbl7t+LUNAZ1k6
OTCrXgmxRBEZpnO5IYVvmQFyh5gO4mqQE9hI8w6RD0BLz8Hwng50J3nmeikGXaIp
tRmGkG4VF9a8AXY1gpkcLjFZLRygK0924PKaQrbtYmjxiNliRuS9Y18OqeLvspG6
UqmHjQL7ahNzG8Wot48A6TLlKJwZMbZVtDxVk350P7plQcVqCu+XnUYyWNMPuOdT
KcWNAr+HD7OBu561kzoz0mX97GW+AyWxHxuE6vFAB8f7vD03iclEJj1sA6KSJY7c
bxKrvU0XNPNnPrgyieGFkmS13kmQbAgPLIBypgkE8riwHOLicGCO0XAikpspvEDB
Wuig62Ub/eLuDXjHnhcgcbLkX2+FD6T5mSHFZyxvmkNHNi51gKAZJrTsvunLOxIm
XimyP7oTXxFPvovSACnxGuztZY8hJH63kJcmcGOoaOaGM78Vf4o6ITppM6nr7SwE
05QkqgGMPcLsswutKFNoXl1I5GG2vq9ty8Q92YncNd4M5JYN4C7E7W/1157V88/G
qfjlN5ChKAIYJWziaOA+Fm7gt3F7CzTfj1I2pCMHutkK2aWXOtWmiq+YIYFOEKcb
4CeGH4u3RvPNPHgPhfi6QiHnFAvoeZg3fLhKmZGMa1teudiGGG9Sq59Te/RQBWv7
QNNByRjsMlRB9Hi/DQJZZjaxNB1T38uBpmZ9v53R7cDOJlHh9TfDpjwxbUhkVL54
UbeTtiYqMufn5Cya0lCYQGwYkwOxK/1VofMlsXOf+Y/d7GQ9lL7nOwWJXI/30/HQ
LSfsdDMFNDvGawiqfVjrYosAXiB2Z57UNTLqiDSkaWltfixJVSZDDm5TJS1tT83d
ybIOcdhm4rfw/SKTYP1tJOp54i/HqdWTlyWQXAIRwwBoz5z6YxPT01rG3WkR4nCw
kqmHTlpmv5rfhH4lkAQc+mudHCk2olFXTIVM8vqFM2/0c4HPAC8To+AlGcBr2SRH
CeOSA6s5/0UeupRqhcymuMtNJq88Km/ZiC58obEMQRXVK26C3g9ySU8IPIzmaaL3
fT0Sx0S+XYdttomX0aPhwi5CrBNQfbWZiftZ/9Sdb5i4FL7pSkFyTC3thnDYM5iq
2cLqFAmwQwwfQDsybeRbM6V85mOy6UY6MF6BSH9reAFidhAmXVJMF5Gj/unwvOuk
NwRPkJP4gMIoWZEXqqIR5QufYDsCB3kmjttXDPxfzGccv4/wgHwdJQA9obNUd3tZ
PpfLXVHKI0ZJ5un/8eNScoae7PMxBz5Y9fcy5qr32ByrPU8uQyZ/EwkY/2dVU5lz
szcPMd5oVJvwQpeK4NSgOudfqp6K/fZ3heZzsVNAAcE2/lgyZIx5Jpl1Pxy7ldfi
BV7hLTU8FzSzhimRZRIJJJSEmjoHufMbuPulGzx4/j/uxcw4rzEKSL2zR/6YkfIl
ZDuWE6wM6UXrzruyKs1xhpxzgQxSGdyQuOfG9pJTO3zyu96idtYsJrCquVrjsF72
ejuTw60fHrVvhQgjrs9+jUP+2xa51tmgVyS/Ei+gALiBIeImZk4uqkM2O6P73/Qa
Bkx1+/scHgG4YF69Yxapdmy7Yxjk4qq6sBvHAytyrV8yAxQ7bbGIOhxn3eqZCB6F
R3jR+TTiD8dRGhKnEMR3vNbDxZcmRh/QFPhjbh0f5ssqiEUJDwllhvVavVGQYJFF
rL19u+L7S5IxRvDcjXTcEusnq2XYa2A+8MppkefgjiIYHBTew69h3HOyjRVafMzc
ike+psVQ0PnioAyfDI22XjWDnomPljk+ANKTnq7j6WhLsc0jr3aGH+NSiLSwQ7QA
Vg6xvOp3ndQ83AwAPSv3NglsFIZLsLYbzyhQdMAmi2Bkci6urSj7pP6AMGTrkiAM
iVx01f7ddNwxr5IGKMNc0AChFTSmq3T3HbmYZAMDQH96Uy1eokwKFiboW+FDlI1/
y2w4Vd6kEWCmxnNtEozqNPTI4mUDaRSwMQgWtLA8TOSMDhMoQshTHAtl916a3sq+
XZViVmWswqlH+zpELPJcGRJapLxRkrsPFkt8/18YX1o5uteptW0GSTEIx0zipoZk
a2WjEMzlm82GO8NXVSpuAJFnWmZVv/NVIXGebXdSgNadpr+gEhjyde5d8geWRl0B
KFiH4g8DJ3uHVXGavZJuB7B+pC1WAC4y/XCpaSQ2Hg2k4SQD7wMhSo7DxWE61HIc
8Qz8TMNPQ+8GsmXD4hBukBklDdDtsrB1sGgTTA+8XMZ5Ol3QvTjU6DRQpzCx6kUl
s1i+XHO/k6LNjEC1BI1YLgGMT+ZkdPKgb7F7Hx56QdH3m4G6+SIY3P5K318F671S
wdRE/nfXjI5Yz8Jsu0463zsHwb1hxnZA86qeWTpgRCdUz1vvjxgEI4SpfMxEu227
zPtSJmlMQPUKGlL2A2Wvnt81PTfaUvQt/PmWtgVKNzekr+ukNl3m+IRWGIKF/ZrQ
N60TFu+tcCiM4b5kGc8lGVT8oxAehP329W9T9r8WJrUu9vXGP5U1VZunkDfzOHUG
KsGNiFuSfTvZh6TswHEgbQcCvDK92voCh9eyAQQG5CVdtzDZ+oDYixq/Pru2TYS5
wtHBdaxfhNRIZOY8iK3njPpQYrLK2l/oVvywL3/KBFvn6G7QTMwrimYZTYiaJYmd
fX1ouebDqyDukL0BGiY6XccCygiDMCKF3Erj10SlHksny4pe0MldPh+MX4DevklG
7s2H+SKr9vrRwHRGN961jPTpV1x71XfRg5ywszc2s6GBP7G3pKJAjY0k4FuS6P/0
2A5kkfDx3C1o0ZFswhvLzxXx4S7INaq6iebP+WMjAA+2TVmmR9gLH4RJYUCHzAdn
hrRjUBjMlmP9GqxZ5+F2EWqFK9aTehinkVD0YNxadV/SifHSJJ6x46Mik40QUjre
LG1qvcd6N37WTFZZIib6F5HUJygznneQ0BhRm042jTzqnCHBkOc9nzZmI5nOgM7r
d80NMjVxhUnUg9s69v7Q+vpb8rFYAqX+IwbG6L3FZgbRwxyo8AWcf3BG5Qfsem4M
UwEcmN/Ixusz04Nd7IKkZPDO8aubVwbhhRQXql9egfgyoKb1GwDHdyuEaFBpybbU
A2dk9VRotMmZuWKvH9yf/rLJIcIZli0nICQAwtw5Mku1pqtvexaliLnztFFq2vwI
+n5ESJxf7AsBXutda13i2/xffEE9TBXPwm/quX2d4Ta8FHJFjb062Wha6orhlcwf
Q/+41dmQzNO3+UAnKA2g2Go2O1QM1DNl6FPcTGM/kaDcbhV7K53WJtH3mOwlgAIj
MMd9gWO7D1xnnCrInlMiQ08kzAPJtDNjjQyDsE2xw2iVvRPKzJk+kO1OZdTH//ry
NoSyVTuVAq4Ab8yrR82nH9vOqLmK6hDxN7BAejcQGa2G34wQWb+QnVhPWywauyLj
aXwMiMi0o5gfFt8pl6O3ukwq2i66S4N74pH41iWAw8s89DBXcHjGJh1tiO+qaxYw
rHPSVp81CpJll1IIqMj09BziW9xC/IsO5kzl96sF2NBDYj1Qn9u2SfQGrL+Oppou
bG7jDj8J6cxfwa6cIOOuAqC03yw6ThaHHXRL9tm231BPF0ZYRtItcg9mfMrsukT1
7WzqzSxzPGq13t9y+NFENtNDsTR79ZWcQVQ8nfeobu1oaJnVDbjD5fQJEzZz8DHn
zFONYFin+3xBXqZ/5MG7/tM7q8h1c84T7vF85QzRZIY7u1nt/Mgb0jdCmtzfqOBm
kEMSoHwk4Eq8U7v10cDHsAIhPL+dG1J67EPt8vQqImBhMwv0MiC5UfYl4ljQF9I8
YzebKt+sO1uSzBCRK5ReczpVA8gciA181RL+P5s9+jjRdUUpwpQhuYL4h8PoqXwF
PP04f4NRegpR8O/IhS1RammjPVn8lmiOvLk03virdIxNNLgdGUaHrluoMAuvWo4T
whC7ysbld6YeZOpBNoC599zGO6aA5sHB4RZgHzkXyUsVslnBFsQPaNQ/m+ASa5Pp
FKmMyZKhUGNV5TQLnVmHclMK/RtHannHN24Et+cKgb7I6RfkQprplzDB2VZYJ4mJ
nob63k3izNlCtB9fWLHSRbRGdq9C2H3B38H1aSPkpQbMbdjelPyaPJvFY1e0j26g
tYdQiuVFCNaPhkj2+67xXbpZanKYj43HZXCbnip1FTtyUY3YA9/aP/OIt4K3Kdzz
uFMBVMv1OTALu4N/gez+bWBp69anfTDR+RcBOg1XFCSYpoNOR2mdJT/cjY5seNOT
OhsQOqjKCNQKm2DV4vSG/vSUWS0k/1KLS//oaBTXzDaqMpNt71vLM7Rl9+9m4xKE
dBoplZrB8pvoEw24PFD6Jw2K8UZG7pqvXYhwyP0Sn9nbDHue9R8Rbzvwk5jQu8x+
+SJGYpfD6iGdLoMvqwVe7WBJr0pYbiTFYVkBubsE+dMdAEzkffWRVRi8B+FWdsW6
82OFUzzo5aOm0p+IrZdfD9o5iTG21vJVAuWxh0Ai7AD/+ZnM6yOtJeQFhp+cd4s3
u8VhfyB4CcXYU9C7SydbuiY/XqcaXHYemwVA5oUrUmrnIkRkkdkQy9Z0bSPUDsUX
uXOSrtBeWITgQ93SuytVc2csC0u5GCXDfw4tCNzN9rHN/3rG4JcejjWl6PLFKP++
0wh68seD4woNbba26cQ3tJVhCcVbEBMvXsV7B+er/fCZWzUI8T4zLci2GA+iGonG
rL8JK4PJu9Y5icx3hULXFWMnnW5deEhdNfeGoMnUEk747ClymYZ1+bbBnMmP1obH
5vDkT3jghiLcLARJUydhNYYNCtSdhKYdL0ZV99k/fZwCCOJikcAZoQz5uPn6TSqD
EbHXzA8vLmhnoBvPXba7LiSG4mk7YR2QUW8X6TG5DFzllW2jAbilPd63V5eIiyDh
Sx+uFxuw2rEy1hWdouNAGeSPAYfli167ZX2r/ERYYZswLVxEgYZkgx460HIaVMYH
9Q6NXy26A9FlEwFZd0bWUoiQBQ3mNMvpS1QRt4qOv7x2ZWWYnQu83rBBWavdLsmX
9kjR8TDliAvyaJW0/xu+D8jTgcX5BzyZD68QE8k1fPLi0Pe2zZem2pv0H6GwLWX7
/kJu0I9EqWLAzfoW5PBwA5Qp2WhR/Drk1gb5WuJH8A4qD4EF08Q4urMb2JQNRz2P
DoWbM5wldl2lQKfMjZm8diGN1T7a4rD3bNlBic/mrSRqpeyn8ctJlF7RBbu78s9+
NQI/lQzFNpBwlGy1gNF16iVaLcuhQm1MQAg/bbuVFE0lseXv4kWntUkiK1Hq9dat
F6xWnRnTpsGfx0Gz8cZKKhgRVCJTbpZpnHHQMQ+6F7BYtRBWOlVXlIXNmIbKZP62
Ygsh9VK+fph0TbB9IT7e5M3dHVwk9LV+1wxMLyfzu0MYwsVAjX/c/0IabuulzE13
W8nb5yORTIHsXLldOUX3dbHj0aXx9d8q+bhItObNXdaupvxuUc3ut/ycEJqWedfL
gxnrsVb0TAF1A33/fRL3BqmRBkZl+GPMVRjp1Iu+1jhZUHGYta6tdLfId5H100JZ
0D/B9jv4DjVesqda6F3+mK0h1iTtErsYlHkzUXVFZ18kOJdkd6BuW8byneYPBdf0
N2AYt3YS6zDjXwBihRzZv9ivC05nWIp3kfOgGI5q0Sj74+aTPZb8ZYAvuOJ2BRBn
F/CjFY/cyMLDcfPoo2osnD1aN0+uuy5qyO+Jnat4bWkDVKj2SPNZ8viijAqWzVc1
nfzj0QBbftD4gqavH/jV4aHRtV61R0VYkP+Dhtm9kPovMBivYG441xomt3IrSBCm
REh4VvqceJ9eqbGqzRM25CGiu8s36zDfZFR45bpcbLW81Nwiijwnph53kbowkR5G
N/heQzXXat4438/V0tdmMvxQH2gYKlUFDN9EpuCQ4EoLV71xQ3fr+QXqMXz6sGIV
wueJ/UtVnsCzKHBcnUths9MwZkrl+4m50yU6UhlVsLeyRE6nu91fFZRiNEt1ItZ1
di3GYhkh9hU6hi4qLhb2VBfWGjopDM/rVv7P2pgpZOoi8cNPsrB29ihn+/4wjyY6
RfjiXA30VrP5LnAlZ+y16gYkAtLrdi142zEeEm5q23JqqbGi4kpILjYy7+eyd/UL
xhrils46WLy3g3jd4PIOjqT2xu/vOdCkpJbeQYWotDUi+w9SRMolqRPrl3v4Mpi4
snVSUT93X/Cx2jekNrZsSWbrWjGbQUI9FiP5ku6eCRkpl6Qk4f7mNPwqSVnQ0vZb
yE6NZj6GK70i/8gt+Vz7bJdAqcT5Xj0L6HpqPw8xnNU27/yZahtyNJzZoGVAgFLN
ZN8fCksrCp7URE6P6Q+cD9x2tjvtDYT4MUYShIg2jhPi6DlQT/mtoTktq0phi3Vh
wGAChAMlfVDTF3c+ZOLCYZszdNXDSiK0nw+2tcFOh6VlL4BxUfES7vPY+aDhNOJg
4ZTeel2QsoOh9GQJISbT1UhkxwAoApsndp8N31H8D06nOBMJ+49LlDww0SgfXgkc
bOJZDAv2KTIBRS2ILtN+MF//5akdUXAzdOkINyCrqg3G7XU+NW4bprdSz1R8QNRt
vqPdGBfS5QgiNSHrUJd24HOsPdoK0m0qrThwRKv3K2r8ONzErhoqSOpzcJnsWvsM
avH68Y9OJKuH6ozMDZAxfiJ+TNZhdvkj1taUCVhTDwRVy8+pGX9LVXd1u1rzH4AO
yzVSBiNb0P1ntIhDBZXpCmP518ZJS07aXrRy9lQP0HE1bag4Wvf76GGQlqC7AX6j
Rw9CV9G905I7b8T92Oz41mbsDhDxt0xOxwaxr19j01aeJmCizwdnHvAGV0cqNPq9
MdG8Ru4AYRszXnBGCibsQpQ0LX83Mku1VmnLEyCCLZp0AzySIZp2Tt9kgc53IDuQ
FO4xjcMr2l5vxEHFrH2wzwQdsHY3z1PGEAJXSk0xGV4m7+y/4C7KDfV5xFxTu2h2
0qrs32s9VS2dtxqLDBcmGpHHZoBThMK5tPXtmR5E5IYAGftXkHHNruzlYaQOnfYM
nVGS/+q+jSqIg8dPco9aIQ4tgjZvpwNpXhaHvppTc6JH3Nay+zqSdtmJVqyMDb2W
P87KFRvuUdpMxRp764p02PwDsaMtmW6Y6NIvEG4ucQ5mRxQ/dgpy5DOCncD7kh/b
ieR555CIdW8cAKkdqv/lGeasMhP9bAUvem5rt0me+BtcDxY9mo96rA8ZvhHeOml+
fp2zlWqh9p0SL+m3sPD9Rs/euF7/0JJ+M9cSRCDNdoK5QtsY/wg4cGCux6gKkC/5
VH8l3bSBtXUvkWoGzKoU/EB36Zzgz59ncR1Hsi1t4lryrkIIQxG9fkXbeIrQ+mTd
d2im2G+T5QtfLH8ozu2lfP0uNp2/X2S9E5wMWx+o1jCJ9PuqFp9Nj2q1NXCbE8R0
BAx1TdTM1mZd1mtCAkdZFnUrIvNq3MQbo62F9NkAOIfLOWn8tf62u/BxhqJ+vCxw
9JFDYg4bgEPcCS2dLircU5FXSap6pzBj/vHBUEnilMe6kOOLrZyQVI+hQvTVfjqZ
uCIXke2k6BLdTmO2abj0EWH7ZTN6PN8Q4wdE29S+wclpjXiRfv4R6V4rv4jdF53C
VoqGa8I9BgoDQNFekAd4EnM7/KG2FmdF9VXKIXdWbrI2QyzHVcVr40zo84pDsFEa
FFKlWM6hB7piaDnSzwxJs2XDfwutSfxtHdBAM7lGPzxIU4zctyFfASgCk6T0gcwk
8oaig23IHbBJ+PgHgmSygJjDXrehuxOefwis9qqxAjR4/HTM4uPGNg3PR/LuDJJi
K3cPsjj4XKCiwau5C9HdksglmF7OXweE/399poqi5ZZl7MBq7EgVil4SYTN+nw9W
kRIms5ntoID1vHWMJugITliZYRABXZZ598jje+/xi+WkI1DHP3dhyYQY7bRI/udD
y2GQkosl0TQvBdyUIBjNz1IMeK7UyAf0tZmqe6w3lV5zL7srX8iWcPLnp4Pqo+O8
9xzDN281jtq8O7N5nSTqcoTBG6igszFWqSWRm4dWplxiMKeU4IUm6aAj2/x4vHbv
PdOE6rRXbRIhlp7XYF7FM2um7um+J6dgVJf1guSmJrkYLkoatFpw52diSCh/7MD4
V0dzkkmNimRjz6u4Cj2cjuJZOFbWkTldx99ZV26BO8WWltoaIN3HBbqGP+g3MemK
Qy4iy8gunVj6I0JNXpezCa8/N1V4pOY0RoTghcx5biEab+dAUqxrvwZX86GpV2r/
RFOFEApm1qdaJxu7UjsZlJih4+W8eNZDjLWTcZ7CiiBPAHViylXenzOtKPLmfz39
w6SzCFePZth3ODO2QU6M2a2k9k/bsTMwoFlhRub3M7RV7PBnH92m7OXFM46abfIx
HEVkJyiSJWQeepKSpOou25Uf9bKNy9c7f7O0DXMkj7y2lxXE2EnJm+2/gyk5gmlh
QS3Z7TvD0/Mx+Dk+8/Z/5UbE9ttBzv2nTchbcPCWZsfZXu2hFQWVbBJ1qMxWUuPh
R1Cn/x2Wj5lIS+KoCRzrkNnBl1vgFdCzvogbAsYYMseLdeWqpG6fMlVFwY3SFGlL
S0ddN/15S0c0DpOcrUVzjIbNe3qWX8atzDpkRSK2jOKrlFlKaZRWgxpTIL4agitU
8uae/2nYs/SUE/aXyRWPSyo9vGFI8cv+WI0bg44aKSPkd4HxB7O2nsiMy8lZjV9x
2lOc3kM6WltfDY0nXUu9O8TQBnsE4zrth+CEsNfv2vPPyzQGDcrqj7+Bu4nuUij8
G5VXe1Z5vL6dMsNPqDIcbI7ucCbWCweDn4ldQY7hwqOPmDFaCDQvT22/xTqYbc6C
L32R4kOb2yO9f3ENvk4T32OTXT8aCq6ah6Dl6NNl2ahBBW7GvI9Z3Ktf2lo+2wBw
ZyUR+wvvYfyz5Mnk/hDXbWyGhITDZF1SMNWUMPahJLWUfVDJazOqIH0VxJyDxaTK
BiwZDjaNS+vv5Omgpen6fpyuygNQQg+5o9Y/GCqGFH1sjPouihJnS4lhFL2JZ41j
k5urtdmAF1/sjQic4LADEXdtt+7A7HXO2MwhzRUyERFRlhPoUSbxwYT/L9Xhhjb9
k5XtY6WyzAEgJI3xwfkkcyYpuxxh9CjKMuudV+yzAhyEFYw4rLvjMBykJyozXwjL
R+FBBoX62w0ZNFXDbgdARKqkgHXtAdjXczMywq77k6c/WVIksw6Cq9N5eR+SAlqF
XgdPBT93+AD1MJcjDrJ34WO2ZwXzvFHaQprfDRtGc9kVFrHU+IbQE/xjN8TvIq6I
JHVtLOklKMN82oxNhmOVgyXKNCSMN/dQirJKYlYPtqq/Yk2jbiSCCxLZ3MNAEDO6
M1S1le2vMdSpYio8o8eh952kuvnsPAzfGdvmQqwoyhEBnb2Xk5qdrcGxpLC0Wz7m
sW4NZrAs7+lsmhJ2RTiX5Ms9enyBp92s+2vyZdw1MsOXqpPPkHrXveQWYNAMiEzK
1GiwBGHlZg67FknXgo9GHr0t7sXj0nB54+uB3amGrme2+GqkBiuSzSDB/aWB6u4p
Qvkg2n7MG6qEOTk7T4b9CQbBR2bXJXXcORhVKo2DOstxXCXvcCTBsGhV20FUCyky
odITf06l7nXmfPTBYFTVrrRErL2B7rdUaGVd8jSiDLzmQRaPawlfKRGOXLQk+3C3
xviX9UCQ/2/cNi3X/agUoAKBgMBb95Sl5DnLB/+TOzW+dK5ctYyjD/Lz7LArqAqA
vJBvpfGudnYZ4roXWLThKQZhpQQencBu4tNLLSmoWOGjkUHWmRsWq9/c09lubmfP
gYg4rTj9whkrVCOtxamXjqPUx9Y9VmfpB4eUwW65LEMeT3DUr4bjeb11m3eShF8R
t8oYWPetkzKo0DMbgg3s/xCVmW+nTNLji+uB9/YW3FItCmpQra+HhLF/PcLgWKvf
XjzhJWNqSL9CQkjzBEMBc8lfhEEovZs0na1uOTtoS2uVZ+DU/VPOP82DjBBoEUh9
riim/lWSmpmyGsDY7dMhiEIm+W041mYpRAw73jsLSLqH/qHMyzakQq7qfBY4trpP
3P5A1LqsYzHHje+2TlaXnWu/4NQM3v5MFOBAaIZcSHC+ntJRmECJvWOPX2WMNvxW
SzAI6C+z+S7Y56ye+TJdDEWzE9s59Xi/tXpsBecR8+LK040jDbTNSfpRLMb7OuRZ
n9XFhTZPxeeW/BFvHvZj/QlfVL0W7s9UppK2uOmnWhSqUwHJzQWA5lNvCOKKdtCk
LBlnO80hmSRSA/rMxforGJBH0VY98KlBmPpUXQ2PJT0ERSiOml9oXPFAZeLa82mx
mWY6xhdD/scl4QwhuFSJp2GFp4oJeywk1IBNdwRnCdgUUbSfHip+SCTPTQAkqhEz
Z6VTL0jtmBVNeK3wBKj5ArQluIhCaxIyipzR3z0LYZ8oFv3XdqkOiemB7NT1dOxX
lv2swlvEXhrxTOZ2vI2elO3U5sGms5nkDb4GjajPJCcC22mjUR+6B6GJU8sHVTq2
tSRSOzmPVz/SXZXIb+Sm/hohxvazI13jIStGgy4yBpVBlru8i024mksW/x/bC6Ob
63o7aouQ958q3aseYk9VDricH+qVyOPoIKcWkpsH1gUwmM0p23LleG/ky0/I6Pnd
b4XUCuY5gL78X/AI0vLa0iTsgdMSwWo8IvLIirdp8t1ITMv4wWDgfqdT70XCsi0d
HJWNrWF6k8Yn2WYnISvqp2jtXHwAXEzd5fs/HL1GYQdnEv9Cq3D/d8sIScBLqkOh
edyPwc6ViEcd/UrYXL0FFdpmEJ/fQiyRyz0Guve/8fRfOZoslr88YJ5CaugES32c
TcM3PRsXoi1p9kcBoKjp4V0sSCs8H8MDWTkAru93AU+cSONj7Gb/zX7J5FIjTEMs
uhHZ4DGsoKpidXYkCmWmNtsDmP/9ZWs1g3pkihTUvKs4txbWb0T0dW66ZEufBERY
vy29H2KfE4kTb5wpOVJ1Xnc2b6YKoy866QxkRL/RQW9vnlcTcSry/JFMbAQJRBfx
KEkhU3AVA10mSqDVqB+/0XzrpNmEFXVcLBjCT8sFYgh05F09ZTB7w0vozolmkXa1
a4NWsepMD6qPAuS7fxTRIof96dEyCI2wU6pZEhhp35e1RwpjhtqwYfqovpd7FuQL
zX8KvZwYg5SzwrLHY7zQ8KkCwjplCnvKmrK+BrrxKd1qt43PIGTSI7BWr3fNBNfq
7kLfwSb+ecJpG2hAPt5hBA5kJPB7yWfv1AFg1IxRLSVd/WOvl3VFRRc+u7eeGkIQ
AgTnrBLP2sowukq8PhHfOf+IA//gtaJYWD1KAY+5C4Kfxn5r1HLRKO0IMHYDHV9I
W8SE+HQEOnRfhcqWX+U126tmHRRA530A0IVmM/Rd8J1vFcXXe96/sDzfd+5obTwv
ckf8JbJ+LkGVUCoAg6fBYHgNbQr/6a/hzsaWsIXiPwiEhwbaNdlXuIDZgs9mU3lj
pEYlJbPaGoIV9ER+WU5KFABDxt4UxFiDh+o1hyIlPVuYoLf+fTjmVmWjpLmnphpi
+ybfhxtS8VV/97Du2pUCUKYfCcV8bBuOZBTwgUfYxhY12WqGkvE0Rigb4JE2qwO/
RhnB5Soc2ckNo9U/xGgFQ4S8vtRCgM9D/ylXtFdVmMOOYK9K3lFXeZtuFLg8aOi6
KPd6Qbys1fua99hW9qZOrPdovaRpWcXAcMbpCuPk4Ejvemxfd1iVrNtoSLBHJ71i
4xPj3yuGYxKWemLtAHCxC9haNUF4XIShFlZdtznBF1N9G4QMQDsnEG4Yw6vXmjPe
TXpdjDKQ4p0mTNNEhtSYP9oLdCB7JgZfC7MHbIYQATk/ByI0j+9sJPFrinvqDnKW
cvfqohmSK+KQQU2q7hIGAbil84LUnIkh0dspdtH8vByglJp4uFpk5hdONXPXuFCT
3omKjNKaT3LKU7mOIedmQ3Dby4za/9QXOuflZiirMNmnoInSfpifu/eOGejGih4z
wDNWu+87cgDMs5cEY4msqAZnQXju6Ty3wrbt+qEfKszLpFxhNEm0qISTzvYEPriI
ZqqyhWKWQ4FmPIOTcsBBkVXn6tj7poMYAGb15HgJMSBjTgJ5k1phxUohgVJ7TUzQ
FpyY8HyobdA3NIXmxCKf2sx4JCyPuZkLMY07tEt5OlSL8VRZAC8iK8U4oy3PY0T/
2b5mL5Rw0IIwVvOzSPgGQSUfwMM8jsnAsmaGkABNYezi7jWhN6wkND0skfZdXNSC
0AjcdjHzIx49JUe7UnsQl1Nzz5lsIRsIWZ1tyUodjTUdP8xv99qS8vXuVwAGB1sD
J8EWO1+0N4Hfabjp6B4IfRPOn+ugoXiF3NgmMkQxc1U4rJuBrgWRrSmgDNIHlvIf
AOp4fCRBovTvsuGCWb1MQwhVH3tqQDnuyORfbjbuIq/ITZeDzF/bJ7sVprPgquYq
M5lkG8iUJ9a5+HlQubtAJYkpePiYs7bn/cQcGMcuQFX/Ti1YzJ3zzhr2jY/exShj
Tk2a4ig7B/3gk5eKGAIzP0ZC03HiwAGXCZGx9K5qotEvg7AsBOKfMlNBWytxu9Dm
12Kw8vwDiV64w8t8CVwjp4MEDfnhFUJf31ERFxNffA6Gp7oI8wGSj+YQdlBg4D5n
qLutzx1Uvssa5XUWeMMQsIsg1L2jzEFTtTK+LpbAyjW9yZSQ7gWRK6DYzpn10u7W
9AhflpGSrLZ7MVYR7hH13hSaLlQFK0Sns3+h9dvEJas+DXGg4J9MIHOueHKSPWlK
3c6Fs8rLshV8cWhiLmepvCocjSJYvU3HT+YGCU/lCqZHDuKPSpmgUJdSyG0/FiB0
L1mFKKZsIqVbhb3n0YThpkI7d619reeD2uzpTLlqXYjc7heh7KtHkGgXB7naFf8l
miP3rfAOUhQC13AY7AqRy2iYZahiVza7UcV/BHRMqT+bwKoDCiTaMVeTko4tg3I4
UFY0lloAy1pSQLOvi1OjNMvw3BxeiEVdjP+IJzPikN/LICH/DtS2GEcCZ7p/zUjJ
VC/phWWx3tfZ8kgMrW+RfbGuXzDofmJ+/tEEWy1e/ZQN/2zt3X6rvgKDx+tRAhuG
51MwF+WThPNpkFOtV0D3PwIZ1Uh3fiMKh3eodp8a87hxaf31o2NW2gpERJSQ6nEH
QZcgahkZy4MJ/0rVwZJWzdrugCOwHLxkix+5xFGnHG1s/Om5FtBNCiYuJfF0QoOL
UrUl8TCIakFjU4IK6pKk8XXWN3JWqb3vd6yPJqh/ub0prVyFzgLi9HTiBfZWI42O
61HZWZ5RhX1vfbXISs/yoWA/jFscyQTQuj7//ODJqu9aKJatbkowjuaJrxp2AO1U
bEtqUAf9zLK/64+dBJG5Kr/vy3UlbYXraXuR9TV3UDV4NU0DwTsdLNihuVKLx5RH
3Y//p6VaD3l9FM7zmGN7FmF+WLmCt+UWUBn6YCyaPgweh3zvAqZdxKO10EMFAoNK
M+Ob8c0RfTi2xt1peT5hel+0A2WGDoNAXGxJFn/x+QAaiheSQ+J1JLxpLIlNf6Rg
0VywU4+7R8XZa09JvVpD9hlKU2Q3NOs3MCPULA2jUzzmySyWACwaCsbk1WGlIV7+
6PCFWtF7HTC1T7THwDpHSIfuDV7yczpyPjE8YKgYrW5FDq/pi3kM+XuM4tu4nOjf
Z7QuVaHtBMf3lKWmeIJ7RLrFMi5TkL5CmTUr5dlOAuQSnpV6JHZafh8fMt/XnK7n
b57D0pXaOKTPHG0cg5T9dTRrgt4KKrlX3EsJKOwwmLcOf2t3GDrQSs0QJ3zvj8qI
rakGkpCKwAVovX7VgiXp/Qo0j7Wvdh/1fpq9Lk+9I9OHUnkd0tb8swaSRqxzni31
9hUGA3BySku2b8PVK5FCni/ek0KXfQ2SQClJ/wQD8/tir/3if21TCpbwrwubcvyU
ey4+mdrTtvustNPjsE8183AgF1xH4h14Dr8p6nwIihkBIaGa19btmYC5V/3qVMnE
SE4dt654Y0qQuztXvaXW0c2jflmfdqTkYgWvBAO6bmkkv3zu368szs9ud+d2PtMl
RxwaPk7O+Gvy7xYXfU44JJbqXndKxPr5oKzJzPK/2ONxGq6CWeYOSlX+3B/5GaHw
0GBdf+lekKNryPu/EDAr/fwG2qcpg5f9NFyaBsbj97/PtyT2kO6/GhPuemyJ4uIi
lCaT6JmBZGY3FI652g1Jib5W7Wal1NT+EeFJY/SHa0YJooG2wgUv3QiqHYwiuz5Q
nmSrLTC+I62B984/JLFN4GQ4GoMYqeFszuF4VMCsac984DXMLJ4gtsb1/pYuf6wi
jVdoUqjqb0WolVKpLb89eNZnwFAVtLzpslyyI/f1lqIyRus9GnXMYXxCxjQBb3ql
pcd/hCPGxa+htho/sq1EAA33PbrluO7rA9QFFTMAX+TrMGYcxxTY5QdaAQByPmBv
ZW+HA/AE3i1gY9Qs91+jhCr0fd/eEruYlDNF7Wd/CK5rJX5+yKe5aNXvREvw6gjh
BWCIj9Y6gNVTAOdB1Q1qbqI0OH5Z7dOVW3ZXpxb+oF8eOTEHTEhEoThbQtoS5Ren
mccVgc9rs4lwwSbc72j/o+P+zeqOEjXAhVM4yhj/svAp6jPIcj1Wa3GkFrHqq9Q6
bdN4bmreVw2ddb95ucIp3McSyIAeAua7+R6+1vLA/g3andxEJK06yAbHh0MDR9Io
6UBD3vfdQCQfB1Q7YOrAq6P3kn4CA8Nk7WhptbQv7L7Ps+GQkKMJrktfVJ8fuMlp
rgcASQocsrfa1NLlRddPwi52Iu+aWVvaK9hkYMsq9WP+dDrFAsq6A1jRa9kIrjQF
KPfQJKxI0ZNKbdsxPhHDxQ7C1r/Qb3gAD9MaKIxt2iu6iDxKlxnr2ARdQV0uLm8x
G4xRZK0D3sdD/3ZhFLNM0jcU0yGK0TRmFQbMoYdKLUFjZUiV5ZPZzGSwj7bslKei
0pQvSQAg0dX9EACI+ry89u1fMlyE253i3oSuAoT/XJu3jXDioovuJnMh6Uqc4P2T
b7w1QNf9n+7xkd954il2XV2nFdK4j+mRTyLKDvsuJMkKFej0LVSNFOaJlj6lO8x+
u7hXGuun48fNrerPfM3RSeEvDfXPCChliJXaKqwDPRiTp9Fte1LxgUBCkU5XNbhZ
Wb4KcenxjSz+23b24vYy/5BkSpzXfDkWr1LvP05hoEhmZSQlP6f6nSpWd15uPrJ8
+sikWkYGWm96k2IR/ERs2csrd4mxTcL/Q42BhqpDQ10kJ3TS2jQPeChe1q+HoYr6
kRhZI8d2AmaKR238XXbDqA0ATCjped1Ei3XSgJExBxx9lUJjhThZNHJLgI3gPxS2
ggncJr62EkSB6fawidJ7djyGPpM5tbDjM61/OAe0WImPLbL5J1wOziurD/+6i1Ee
1T8+n7yrF51R0aGM7MxJAguFodGRqVRLPxiXmku3k3s1g/VAXfyMuHsDCYcNBl+j
EEcnSKu+SjYPJditlWp7/NXEBFwTj3ByfVPJxuGLOuU9QhXX7NroX8vfBc8I/PrF
uF2A3CEip3JHZKZznWWQPncbJ64uDbYOHi+LDwXPHziYvQMFwzybwclz8ROgrc2B
/yCj+7ACj2HXwzxVLHF016jn357Q+OZHCVfzP/v1OVSsZaDpdK3pQpE1O3NsbmNC
P5qkzytu9/JD/Xb1CCIkCqgmzfKqYu3uKpbpclFIS/MXH3ajbOt9eqSMZzC+9wWC
+QRJqvYcuVfQYXr1a90RKkOsH9mYM6xiw9SieLvhgOJu9mMuLpArSeSYbvmFkkZN
z4NwYyy7o35wKzuo9iGSL9a2oD/lQkMNJ+Pq3KNpE7XSmT77ahK4Fymjh7gn9VKy
Im+YswPhRzDflXWW5r1yIdp4lerbgecND+54jTgO/CeH6ptObrlh2CV4EKuhCDEo
N1W5a0aJZ6URvqxsLwHUEr//ILrLSn6uRbGpKhFyLwunnKLjJMLIMxKdhkAGUgaS
nGGi8oORQ9hYVfCUtjKEhrAzw/3WNGHnpmqFYnoq3PwENZvGFnXGqu127axKBfid
6necneeomncBvbgFSMsznu607Mk7kuHT1zUqBN+seL3zFKxqArLazh1HjfER5Oz7
CRQi4Xyc5m5ag0x80ZVZ/EMu7XkGKoJIYszy1D8AHOj6BUEtl7zdXPkiY3wq9dKv
11Opjb3tG2BDltn43K42SVuOqGGygoGRCP1uxPVLBslyxJKoeFpncXo7Jihum1ty
HUuSVRPG1SLJjEQUrHWVztQtGbZgmrnT7FuZuqk/Mbqcqi/h9HkDsfChbibQe5Ef
1t+2b+TRRwAsF+DNqmMXcQc3AAHdbOUiimTneYj3t6u1LquCAUMjdmBSv6N7rPpO
hL58NVCmCMDA13sDNO1nEE563gUw3LloLnE+DkzoyzUQu80+/7okEpHdan+1yUMy
fuYx1fJe+ShAu62NIOb1QJspNCd6YYHwqmjfXlzeP8PnVuMOHK/7mXAfGiknBs95
ajH4DPcvk/jTGw0XHjkZGjLak5pYcNFDQkmWR7lHerBN9s6GvqdcJuBAItD4keEq
6+6NqRsJcUGb0p3Du3Z4StdF7EMl0HabYhzFEtpsO4SL21bnKO0dWHMUD/ajD7RV
px8en6ODiwgglPLKIRqcn9jviNv9mzqSfFSHs9dmvtXQyXaI8yp+JhmKuTpeRinK
T/pamPekw1JB6ohThWNfoOxP2GfcO3I/smV20DcA3B+GMF+BgaiQ8En4sr9NLslL
N2bqSRUOc8Df3C9RUy5jVQO4SCLjpuda9P+brpfWqDkBqlo0fjTmuh56cd+vPJI3
66mKHH9UWAGFYBV3tgojnaX5BS6GUiN+DTvfrcXu19CbtfLnD+q+bZIkxXXGHKKK
6sJmZ8YwbgtgJLswzCAP4DkSwFgaZO1CrdepzBTyZvbHkvNXv97rvG9ENJL+sIIo
2vRawEJ7IqJ2ZDYQdMSiXCvActVPhketpBCid0C0pz5eWg3DxEBhQOrbRCQl0c0H
92bKlEA2NY6TfHAkGxa1156KgkHIaHU+lkDMQ9cCDdbOtnxnMOJ4ZGEOiSz2+Q2D
8EI982rt6TXE0ckH/nCTjiHv2ESM2YUw29qwILSVEKmZi9sltcszRjZWNnYjW7by
+Ev7sOO6clTkYVwgk2IZkBGbMSf3cnncZTjcsOOzW7UxoU+D0YntnQ4wW3taJEKO
8wdJDr24pDll92gSeMiFeCJjnnuVm4aZdrlEIQrZZpDAnULgIgZ7lBvhH2FH62ja
ButB9vcVcCSkE0hkjdOwd38x/2EdhCvsaoJBS0hrL0pnIK3gZMVXwH3Cc2PnOx4o
m//HucOLkj0/cB4Z46W4FtBVkQz1k8k595td14hRxk0tiQAageHWQXf1olvz/oWg
sglVsIbWfZNoHqzDvGWN+jeYc/17jWDDmJVgl1rPgGpZzLMzpRcqj8ZLMxg0GgeI
GDSgWPJ3sniTen+l7hVdBJM2ys8cTZcWxHzCE+o6LiUhZLrom0e+aOCRn0Vt8v+P
SGi3MGF1lG+5U+agVwzk959J5NR9r0ijTRKbpszlyh0PF+5iXr4zJADhlY8EDh0d
QRD08HHYw+/ea92fKFcULIF7ih5LghQyj6/m3S2sv8zFOr0N1/xUQbFnXE0GcNeh
lMzVuZ0l/TXnJkyYJMTVmu9FxWGR5C7fGgvTKFY7eWclDmhcuQRqiTrBcvA3tV0m
RlUEwXyLXOvYHlKZXlvJgUBQGMMonVRyyR/1NF3agoHr033A/iSFlc3g4IkYLlt7
ZrZTWYrPu022PrhlXDdsZ5OEomFmtOSZ8JrsiV6lRShxgLAx3/7QbiscwkA7I4Z3
vvwocMtufR7n/9njUQUxX5qdkHUl9qogEeZbHiBblblPTduiBABMOxznm7VDLatO
dcWxpGELfE7kDiuOZillmYgFHm61kP/qExgFZg//0Xe5vOivK0znr/or59LfeOBT
HkoSQPKYrWH5aRk5/FsCpOMuQVPoyeEZTSZh7Mu0veLr4xgsKnKTUZ+nZy4H/FAb
XO2Nux19akf0e0KgeMjVSVGkxxUrqG22Ie2WF8Qs+v6Sau0NZP809uewAQi68v/Z
9ABoypMSEjhEsLaS/iDwqGZob+JWGABmiZTUjKdt1iCB17XdCn3IqhezcNRPvGxk
WQIAkowMfgYJxoYykr/NJd4PGkZtnbU9kHnVHQIJQbSfVol1nRCcUAVCuL4VF6RN
0WRkYCY7eU4skroX6ql2RGp+fr8oJJXEdPsIxKAIhPmW0ckXas9LlbkoZsfq0nmW
lAFhWATDKalW6kZn+X1kVFZsvVu9aNYl3+ANu6uyh9qOIxy6+Xnt/q6t1UHtxaHy
xfalKb9zNNis1IlraPeIBxkxxQ4ExrM28iTDrsErKVwSyBs39crpbayTkncYxeAY
3rK9bYlWAarxD4TJz/vFdrBoABvj+69RP4LW3JAvLpwz9sUfT9IbtLblS6Yy+43u
EvwsmzPhJCIXvRZoVP60uelyyMIUn18K6bxZXgaZpC2ubNMWjTgXeFq5s2AEOc05
0qrjjCcKqMswaXYUwJkdiqHFbIPneP3nIUfMXxAXyNf9jCLnnQOD/SwxXJfDnLRq
Ee5UZ8Vh6oS3wGQDPj9LD9VBg52PbtAa7moszn5gm/Esm9NHic5Mte7KpZuKRpvJ
UfR0AhFVxJRQSZ5U6x6Xj37K8Iy+CxWOq2AnJxpRvl1YCca8sXYOEj/GBahk0Osw
HF6sSQC+Un2nCIydfBUSUKsP5R0re5/pIXg9NL8/V5526jKeaC3toMw/c5DuSYm1
x1oavXaTohXeT1/3Jmq+eTimXXVJBww2xMOfLaHJ4NI7sbFZlhc4ROVzPznSPGWL
X+m19tF5vXvgzVdvbXkgRoqJJN+YJp0whA03HsNjvEDnsSwCYaiYB8q4zeegOwxE
bKzGEQiXuDki0t4HZ5ZQkjGwpI3hOfZV19WH/1aLmGZtpNETF7sb03oO1n1+I8/e
KBRNXZKlQqPIUhIxM9mRTp3NKpfQPhPU7sIzlNkBas22wXswu4IDZjaTfZ/nV5L2
0rPzj5RI9p+FIZszdm//YWbhmMz9HUNNGJr5HUZOU8XWB7hxDAJBqoh3FsBl7N/E
dJcdsKpKUlSdQV+jhAFhfl3uSCKrY6abOE2Z/KnMtSbxWdo+vD0FsaMmPQ+135E0
Gz1nVN2wTZ23h234rWO07ZeT0cdpwzHoqr09QV71LoqHDm8UI1xufZwbu/e60xzP
ZvJrmCjhylUm6nBdTnohZbstKf7qjztjAH/E0BxV7iT5X8fYjADWRwMAYpvzW6Es
oS2Fn+Wab4NaSjevKK6hELoS+OpeKazaq+7t5SPMuhAisNGkn9pEiK4Xjr4b+51X
f7wqay50fY3/PZPC/TBemNacooEHIe7fFdhvDL/Vw4DmpD9NqKspNYDoQplzfAVc
koVXqnvrO3NH7mgPzft+3+pG1X02MpwhmFH6lhOV5YHYuw2wRZg5S3ejKYG1tjCX
j9HdFI0e2CctUqeQ0i233ehWPsOR8mdt3w5dO8bRVAyEEtsEULsYDS3E6T654jYK
SBfcKNgqeGiCB0KhmSczc/1M29MbUPC3eB9jQQte0OtNDtkivMTeqvu4oaE+4DAi
jeLcn8bTF9XW5UNf9aAaa6/uudbgSt766cZfqsPi4ttxKp2c4binSv5uv/lZNc5B
vS9QKpEeQZzG3Lmr443+bj2ympbjee3QhtXNIKbuZZo8jYocCyjR8USxipE8zcM8
whUJ3Wbwg/d1zjNQXvbRS6F4h1DmY3bwdLqfkivzqaYT8O1U4KKwx03E+RWbr+kl
GmUBPeIPf4enTmgnU1XfAdjTLUxVAZpMs3ERkMya/ooxS0ErC6VvYmpjXypC0HGR
iDR6vFPIRq6Hr6jZOYTGprz2XFGWzW9PT780lwqx82ABKeydmfl5Ygk2p57giZ3e
t0OAzugzdrQrKIKs1AGIilG/HYOGMbYJd6m9At0OfD+0Hk5A1ANB3YjcvRPFkLRC
YEOxcxsuKRHfq/HR1qTc/rdBm5makYQnXRs2IaCks60dO3rXGbqHg9/x6Y03JBIr
eU8XeTC90RjM+MrHFsuvmtAjh9qKf9getvBbOZ1VypDzP+bUs2TedbCbCZuuHGXz
sU8Yo4aaRxQtivI0ax+EQWA/el2toSzZlvfLhFLN8VLsKs/4AtPqEPvWOg1Zobx4
FSyyo6Igdqo5AOCQPj9RdC0THaRH2tUeKPFZgmq2ZewtUOPLDEIw0CyVnSPMVSq7
aDP3U39G4xFL7/l5pVx5ldFv0MyPPRtC5rsyD3gX8WeCiPk6626hGxqWpxC6k7Sg
xEOyWV7FG+P9T6yMDlcF6SWTOk6pyV6ts7Ns6L4T8hw2VTxyZdznimAbbW4lCYDM
cyoFTdi9rSRu3uk5LP7KxgmYEKSwRd2wEgFEeQV5VEptczkY9uJGtBJ6GJWiOkK4
34XhX14D+Vi7s3CM1MZPKZ8oSQ3KQq0wgXcvVGIFZH9DGUHM99881+QHGldyccEW
oU0Zjsh5ShEvpQJbRfvtuZkK1p4LNvVK37Rn1O84XUzwbsDYV4E4naNp2C5yi71b
zh0PkJVtB+V4Rktxv96gN0QVMdpr/1ZpvlyMfyhlGcjwe5pGubt0+RI8uY91fOJw
NM2uMa6/F3kTgJ2AFE77AugaL+Fs6DLg6yZ1r1xt/QIFhPkgukleLFfBFUUgPYJV
2oF631bWNItGRNz8+YEjFDTr45ad/cnLsMfO9+KuwolDWPaz80g0UVI/pHIiXHU6
PQDe82FvuWS/JWAvkkyH4Dsc8a4cQ8TA29Tvs+NhYsV9tVPJFgvIMcE10vpqvA/m
24XctnfJgp+yRD8pOsWysEAstCIJukvBnxqrN6BhmRTyDD3v0uc1voxgIVI6URsF
2yLu74ZjZ1WUhgIPFKmtWdFvxSXvvlOie4SBKwAWxqjMh4T6KKPiPJPvYaGOl64K
E8PJWhI5aB9wiAlQ7t8DN3OVDgQ8eOn5hEM6m6xM/HmcTUU50JgO2YiULc+XB2ii
FsyUoX0d7TJbEBBGTCzMZh8MReQVWRRFlNeH0647tgdGRn+Sbm0e5/aQElYMvfVj
spvxGW2e7T8HnGjWWo4D/oFcYxlGOfOyHfD4eda2mwtM+g67jDUWaSdBenvsRmYW
kCWofDwanWSxuELHczUeDN96kAVnsLZRaKBvmjbP0q44zfDwmNj9k5ytuu7/QvMg
aZloixpzyuANmXBTkNLDvROWUIV/v4Si/720puRecKNrydLG4bp/CphHJLDhigDm
Zh1DZHe2mQO+Kf6YD5R+CetZ6Kd/TxRWMdnvlvghUoeCJsXaW21h1U77Y+gM4JYN
pTV2zGi/2MAXqU6hQ8viROhKON3ofHgiJGxlLpZ/ng6PfXjF+STKsT99+oPqR/VZ
qREoMGW9Xz/APjwT3jlosjjE01QY6s/ID/PcQd7NqLKgERW1vi3yRupqV6ilyZwA
8R51ZP+3nNg2JmHQq7ftmARi49pM6pynMD54Wq5d4rvNheDqXaNwS5RPrj1KBeKz
hAHquFGQJoj22LiQoLlmDYQHQGZuyuHL/tIK+7Xb3hWlk0Ya0ohaqdestKTLsNsV
nfGsaoU37sNf2hor4HQczbPbEa8fGwC4Jnqueit23W+AidK8h9jPkgrgqtq0HtAK
z+78wyeYvzUnm+24qGv7hKGFhefOx2xSUKM9Kv39u80I2/sHBbghxGrAlI1JT3R8
dw0+zG05bSHa0NV9hyDNXtklAr8q1G6EJcrSe3z9UA015E0mwUE0RMUhTkyfpBtf
gPQ5ZF5fUem++Zl8/B5rEYvUJLoaC1X4J+kbyml26WRkhStuBX4Arr4ea2hZDHWm
vuD8SnyCSidF+wBFgwxB3lKgeZGvcJYd8TupcTVvUi3QImjQnQpfPJkdlByRfUVZ
FDJJ8BuKBG1UrDhPYRoBx87q76Fn26nMIXyKKwRMVPqQaxje4jym6PgzM81tcpgM
HIxDBKgxk5IA7jna+ClZZYie7wxeSTzAUoAuhK8RqEIsoy92B8gq4vUBlzq2E8HL
y/zJNcVesapU04pOi4HxoY7qIiDIDTbxH1LlENLhyh93tpsH87ndxH4j5H5NyApF
0BVLmvri6NYDoj9epWiS4S7FTQrKb2a+z79LqsLZvNC8khtqkBBzg+TxQO1UedSh
CLa2LCoMUnbpoR7XufMcMRyaFNw3NrE8FoBVdYWfpkRdXHj6yMxh80sEB4LZOr5w
bWoA8I4YuwMPdOSvm4ld8+4uNTKM/qAv/ktlm7ok+Mb/WjO8piP8l7g6e9eWekOj
ATdcNRvTPCCPOxAZC12upQtuqTZyI7Yy0+pfr3ba/BZwGkjts9xQ5y7aZibimR+2
dP38vLnxrMhg0vzwL23vb2Rbuj64YJd0cfiDGl41ayUn4sybkWm8bdRsdaiICyDR
rzmcKcZbSLE1rtqt2S5PLUxwW3ZiuYM1Mr7T+nfaqabJyGn52/Rr41msce1QrlVB
RndKzX1O2vVjAeJgHOuoZX+pTWOcCOHW4ShV/tcabi0wdGiw+25S5YMJERVEOZ8i
+FkOWkMQ8G/IyNP0uWXF0XECzyzXaHEK4RWGt7xwNHOlqdXNLvJJnFJa7CnApFYd
vB4hKg3ZeNN3lzO1aO7DZiMbIxPXILbP2dpIXz/UQzEm/Ou7eB2ZEAbH6Oozr3wK
kxQdZRtejgjfkdspkJESwu8Vzu6gO54HXC0IEnyOu1dOsPeLloQJ+Yf8ng9y//gt
sKmWa4Jd5WPvMstBvHu8VdmaSH2oAdOtLNuT0Xps/cFS3uK3Tc5YK+NUqgS2eMIc
75yfTkToc4JwPOjuJmANewlA+Yk4SnWiJH5uDC7RKsb7qXBjM4/iynDpuCP8cQJC
YrDebwkUT576ECQC8gBFP5YpFk3HvjH3vnV3OfPJD5quJJO4/3S9en79QDFT8i0v
qQ2M9W25m2s7LgUzjF5UaWXVowad0jIusCVD0ToygS8jwFAFvyioppkn9lHfNuIL
J60F9rsy5xDRjvazB3Mc3lTzCG2rFLc7sinT4ba4nFQ4cdFpHGpwZvoG7aJ7bxVF
yahn7Kdbo+gan2gUovIyN4CwLcTh0wka61S7R42EGaKoc+O3JcNUAZA1WU8nICfL
1znBGadk3dKoLY3W14xiY++Y5U6bTdA/m0Ga96I+bxcKH0bxTwYOim/ymvrIQama
FjCXz+FB3mbXNZjEo2F/Xt2N9GzzYkHczMvT9wieuTH0i3nX95LG0FJ4E40rk5HN
HQVo/rZ51dtJ9pcOaobxZqwrEzY4d7UDJvkD9Ok8IGN0ECU0VBqT5uTXjY8jhN8P
tXJ3E6gfnEll53aVpRaPYgN9+4+nzsrsq28sIKEVjJ/Pno8XNXaK6zDDVFBO+msV
X7pP4Tr3vGwtlLe1zszEj2IM0A1QdKxeIuIutKRjPyuJqDPcGjZ+nVFr3vRJHXpq
jpsvdXBR7suq+KmyjQXmCXq0jSbApIWB8BEPEw4haJxBTA01keGCXAEPp0bTGEx4
9RPxHtLXQq8nr7qhnYakBxpcWe4wzW8UzlQFW5Gf6xYl6yIU15Z9G/kvoCrJ0J9Q
kwjFQ1J7M76U7wK98JfSac8J7aWhkO1DTTgjGMtSN8LhLxgxgejSBMsebAvyid/b
1jwjGaTF0XjgDQZDtmz2TjDfFU/sV4sM+QADYJMCKIHrA4zWNl/BRkFonW2yieh1
KDtRSURcnDhYxuu2J6vRa4QKw7SfPiXl0OWGpDPfWRWZQkwNxfggsdzzNhlkRHnG
6MZY66G2iKO/JG34yrglGFSSqEZlsU7jqz0e3PxHQ4loAASpyasxefteO/6B9wW3
uwnoa+c/lqxqQDxEt5rPzW9UdP3yZF+98lL4X/O0X2x1GNroN9pia6HYCRPQwYNH
m3yZgjGkAc9S0OJoHBq/cXPelZvid+ezILvAGUw1JnFBPfgk2jeSimdehcRATkhc
JUogSWWtZO8PTJNk6/SU8GUSW1loIRBFBAtZerHKhduGHvM+75IBZ1j5DgajlWOc
PP7awOEnky3XxsqsTuBeYPdtA8AROBQAf17GgOPjWwEvlJLHwhUOfYwgtlLL6Ppu
/2FXTjCjU/+ZdVPO7IhyFvlYmnArvqGtgeoHAEckFOWWOykkrtBy9onJTCWaPs/6
mk8rSotpat3ALv8FgV9uziZnf6NY023S1S0vslEpiyijCSAVyu0tqFZ/LS5I31F0
yfhpXoWxgPIV67pUYjdWIKHZp8tNZbYkbwVTRyKXYP83MJV8S/SI18V2b2ocsoA6
VYnnCzklr4fbjHADtk0yX5GWmxFC3AbjTBmpzk7eq2PQzrQi+TBIZjQ3bCIADI+h
J43ErNyCkhanXKSmxxkWvm676D4+HKYcQEwAvzl3Fw5YPYk2lI9zjlZzJPYKML6b
DMQZ0a6sUxLlW1WGGsnGgFFXy0fZ46mT6/s1a6M2+aUeZ436vn1g1eICTqqIDAVL
arYxXZmj0yr8aV5Gwdl4UFGVNkReTsrucb/GDWMoJ76Lrj10oOtCcqExDAT893hJ
sjkvsz2bG/7JCiAFeRjVQeH3PC8FbEs35EmDEIxiyfOVIJ85Tw6aM3Y6H57q+Uf9
+6f3TimNuSwGU1EIY4eGxNisbo7Buj2Jr9M6gb6efqVd4P8un65bcjixZMq5+4Hn
taLBwgkR4c+Kbi/RU8ZoyJdbLFuOiiFiS0pc3EoDSX2gMDomR62FftF7KNsP36+2
nueb099uw2FMYkWW5ZM1FBasVS/bp6PE+BAMkcst7UkAebEtoGawpBjurUFHkOy9
ukoPcp8Po23yUPxEE01DXYeW45fkDvu1cDh03o9sCVDvagKa7w86td3dbNYPeLqO
WK+BvdnEbLPYz+aOMuII2KwQWwUR+FjrHsKFxQTeCbct4N5XuA539RaHiX2TILE3
Pv3co3XpZDNTEnfRzQI1BzmNIjoBUCxxP6Exdz8z69NFoie3b9A3CbqSDaGUbEqk
W8NekTEJIWc7rZFXpvxK1r3d1KWmCa3284UUlN6bV8OHY80o7L8iIasSJqoF2f7M
uWWt8O6PkOoWAow13H2LOo1HQtynhM/SYuAGpBpQz9UoxzsebMH0cLXRc3AxY7rW
okqTBJKAHEonQV10+Fh8BdHXUhtlCahjQN3m7U3XanMdiPH/gb3n60PDYWOYxtlm
/sGDWO9Qs2UwEYleLsZiVY9+Frof8hdNNAlBHsN1E4qljoXK6J88eVacZcfRQbAG
h1UyrTEla+X8wJrlPQfLM29gExpQq6C/ytZYdmAasxRpBaf0VnAtVMaWVwzvt0cx
2jxkMRTIGdM7/u2zB67LXJ/6//paV1NPTNuYwWFj/4Sv09d03db5+EjkT337SaRR
75wQzS2xlTorWedgGCk+vsVsFzOM4WdTjzIrDt1R4ie6zJJhqlrozZqEVzMqfBrL
CIeO3l+8FdMz23osWoErIPgvhz+8/iP9ed5KCq7RfnoWadM8rafGhzul0gSGl4eL
8dzOiX8FiDeRA6XtXQIx0CRRNWVmvEj6tYX8uSsOR9Enl1FmCrNmdz1PIQ101CTu
GpgYGS2OGnsfDr5GjIhG6tij73gl2Uuq1F3TfbrPUANmtOvZbo6PO4CA/R8FDLzJ
iEb056PwDnrll5D77p85hEvzLsHE7WjbbHasUdV7+ZIEHKk63rwh2EvYjqkScgEq
6DNE9PAXMkmLMOO8KRZXkuXOejaj8f5FYgmUB1Pu81BkhcPBbKvGcUNQhRh9jONc
w57fwLJqFqBp8UKNhGA/NEhpD31Tm1pu+x27omZYZqPWG1+xBMXd3PnE9NV+1NEA
Tf0xZ+C/2nmvF+7aytEw7ov/NuQQ0Kpbobl8iUCplIaZoxYrqnEQ1FHY3BtoYNkz
w31rLehWGusbhfAa0ESoD3VEO26xGini2mKEt+OOXCwHIvSkONVUz/gmzuH06Ejz
GwPWkH9eU5/SV/Qg6L/TsPPxqpHoo8Cmt54/Lzw/mPauzf973GddJL2GnUs4dOOn
WMF+tRzJ8A8UTnPuGa3CYEuCjDBcq2PrrGptBOhvO2icis2+VM+yKFT97hbzbyMw
VwKTd8UPE92UcoE7I1NigCUUvplYZDbhW4IQSG+lK0C0UCJn3zeRGMHBFfgtP1y+
umlBahGADBUyeBtppJHqi7G4AkgFlnhb2KIuu2lO1q52UYgKv8zohrR589acxODe
g7EWgVgr17pg+6SUC782Pvcnz2JmJ1SlGAXf6tVjGMnv+cuJSRwQuZ0FwBIv+HND
X4QFRrDDAHKL8RGtSnpqN1ZMdQCGn17yDXCcYZCALE6cgKKWHnNruRtg3pjeNP3N
SvY38CeMmXGWrebu5KLfrjKwsG275M2PNLw2wfLy5xyn2seN1BR0DbYFOnMsWWO7
uUEBp5++A+ZGpS6uIbnVobpfDnTF/BKOksFleJ5DoalRLglkzixd4x++ebYAF9en
BcNblOTrGnECx69zccXACjGhU2qOaUXYqmajszY/CDqjQlnaceFdPi5SmbzxOHXz
sqTzwtkdsgI0BvB9Czs+ZTKbkWbqqw7Kvvkh5rI/iyof4W6UXmuG5jrkIVl47pph
1ZVll1ReRTB4+Vc8FyDpbdkMlwO8CS+KybiYhSAm6H9Eoo8t1bBX8F7QvJPeYRF3
VRCOC8kM3n2TRjCyVkVSdRa+N2gshVKLspPcu91bzO4qG1k3WiQN2U80KJ6ytUJh
bRMDS0fcwfUEsy/fO8HdF8SwOC8nyTtCRwNY4Kv6dUREoZULqFHQClUTPJHwJN/1
Qr5hUJRpSEbNPPF0LE41X6LEvOrY0h8Qg78QIYunwWqFMG5ftoW9Pbqp1AkS4NXs
1KbWQdVzDZHV/aSCHOcbQnkk89rrogpHlUqYkutlr1Kh523jsPGk4PytNkvumk8y
RwyKIOPNwLiC3JChqylHxbwltRz3zeJueF+l7ilzgiDlzry+oi7DM13HAb5oTam7
Db6KCQ6RHILP/M+Hj9ZYOdvgIrUd5ZzBW0qjQY14a08N002oAYqFPLFJ3Qi3ajJE
dhdvL90BKPIsOQ5cnstXiS2geuVQX6ogZq/a/81U7cbzk9B1tZgtNwZ4DrtQJEak
zmJt+Pd3cqGM0LyUrXfCeHFO+mkjCE5YWzsuyfUDXtmzR+7uVT7drFss2bT22E4E
JbGXSHIgeTwOt+D8aRMS86Bx1siW1NNqPFMH3yaZo3VrjXQ4gvR9w8UrVx+0jQY9
aBJQvoEi9qsvAgFWPJ5Ui2ETVW439Vbwg91u1GbKcD2JUyUg8irZrJGL3XMzcsyi
ZX5BG3USaxHdD0hx4tF2y0damZAE6MEjX4ZXLt4AUKwvVx9yN4S4uECY6PdMjb8B
quFJprWSPeNW9K+OmNlXrvtPWY/cNAanjTCP9j7bGI7bflKf/UR2KroiER5g6Mnv
+yuxyPdN6JgQPHmrIaDstIRqiRg3iYBM/xvS4c1jWD9kkEn1pJ9yMuwx0YSqIZer
0uYjAkoF7lKZcCaD8NuRQREoK7sObQ+OWRTAQLJGVWW8WiwLazFr7JtSJyzUbSDp
UwCwPqQTMbN5YMIEDpRWGsjqYP7PMyxLX7bSX/z4RAQ7TMqgnDG2PXlVwJAZnGRz
OCsAuB44TTOu/YLX1sE1/j8Jzm0/hOeT3kRBIg2g8bgrrhM8h99ameIlE2qnp3uw
b7DzSZfcAykkhu6TNFEY+eATmu9vLnY2fDT0FKv8QmzHXeatLnjYvRIz21TkzKwe
W/lImVkN3ApLHUjQo6MEbDBPMNiuBPkTiwoz+03iigxbaRtPXPXxRyEJ4Wik+eM4
WNThRy2+haqtegDqmwpY4pUDzp5j4kf7ernvMGtaE1PxUO2A7eUzXxUz4/F+vjP6
1Y28jvyG6tC9y9HkaeaszFFYHPPjDlT6PufAvK11J5EAogEtOKFYC8QMKcX4Y81e
0BhX1loJO7wD6rk30P5kZwXW/KLXKqQlJ5k/kQv8713aj3vX/C8G/7d2BKHnlD3a
niC5ZBXmTPJheM5L+gnDNCZljEIdYIDApgG0TWHp0q44ee3giwa85UF3dTIc9j7n
eXjg/gffx+Ndp5A9gWD1U8EdYmc9FytsqPItvtvwFXLB+5ZkEPkUS2C0OjQnOunF
wbMAoWX106YPfvl8IZDYwvTFsNeKJcMailEplbnUA3hQb1oTAGP+s/38NBsiKiFt
Va8fCUQ/e4k+Q0sUCbnQSJtMdy4okyAoerY5nj8+zdstPNrbe6sTsq8h33/1G49d
/w0OkABUO2JSWogQdWKreQl4nQjUuY6pqpKUve4GiupHRWUfFhvHGYhJJ7rBWXoq
iJJOjJvHUsbTYzCxhmIx0TpJnMaF/GjwkHj26fWOzLpap7WWKpnBNzntocySy9PV
dDmhfdnn4PQr13/NlJa5iH57cE2S6/SJiaTrlh6f1+nRQkrlS2lg3FQHLzsYTzAZ
kCFVQwfhY9a1ZkUJAZd0wNN03UUJs03Aph+RPMoY9RcYSE5dZU/rid3KZSbcxVq4
zcS4j7pSKMt/JHJ08LdqsnjM1CrkzKGSNunpUZG0GxaAbYl3GXSaYKiS5z492aBJ
k6gSCY81ctmUm61DpOmVBIJsNgWB6eeakUomVn6Y4HPJQQcwNrQCtL5euRtbOIeW
YQQs2EigeYhYzwIGjoqdFIM8ISDOhpvbaxHyQNo636PO3o2vdPjd/AeaLYf6AZJC
Ba82e/6FZc1+pjvPfQKYYGSciDHo/zs2VZ+Ix4eM2OtRxCFtLRmbluGDC82+M4pH
kj63lNPgIKva1tfQR6KjxxRD0mTTVqeONOEKMBUPPigBzX67jPuIY2YEJiKuseSp
l6FvfjlzXAIp9r8vllTa9Zk71N9NBGv6/1xAIZh/BfNg19hDxoADSGDxySH8st1b
ERNLKVexnpZZBcz8rXGDRhnqiD8llpf02YaZwQ0xnx80wiJebmTgUlvq37+6ynO2
mi9Nei0pgHE5yU9zoMvdxWvTD2tg1xHy50oE793QRHDiaN5uc4NfP0kUh369boYQ
5ZKSHvs4vQZtqZUZich8c8+pTe164PU6uOIekCNX2klfe/PQ6NdW6umJdZ3VXqqO
6SpudaMS7DmO12O7xveMgXHZ3SoyQuAxTovutmH2J43ilva61VpvCU3X6unV4aBO
OY3+PXKf0VjUAeE+jIxSNI+AqvtfxsgAEEEcCglf2n6rmHfqlBY1VRWl38Kedsoh
7Q7BZjxMWgMARwMb/qFfEEmDdr3BxCgHNhHx3QJahNneg4MUsjWGt9+rd613XnpR
52Yhhwncz81bHXirZbJyJg12psGSBVNtjU/wWAsIBNjXU9Kp3OjdoGL2J8Ilfbnh
bpKqJDbZhHWLftwPre8FojMaOxah5On9nlagfnOTN1jlUYRiGNK6x1/8nhfRO3+A
747TCbQqqbIE/oI2gXlff/rCfr7fawZ3rdTqId1ec7/lsqcZk1UFqaeuyqZXE8Ho
FXt9ToxnpEu2/hDSRlNELL3nQS0r4SC4ZUZdZ0hzVxW+o4FgPsm7xnujXkJ8zlzk
fL4ul7M4TW9YjWIHQsMMbpmNZlMz1+tibOwVFq+jJ5c5gplBawznCd7vBEmi7GYM
ODBe2OpyR8sf/bHIc+Lb7CiNLL7ltmt9/LaQiFtuzOj+Iz1M7Q6pnmfNr5HUJR1E
3BaTeQ/EYIr2zGQXneyU9dibdvlOVJHwBLr19NaU7dRNeRsUqMczApKt8WJ3mzCR
69S2jqYolGK1VnXKpugcouXMOXmp2f/y1knHVryekTPWUM3zmMwmW1bzUiY5xkMy
1N5ZL0/XOSkl58jQO9728dUIRcAWROvMbZxLpC8LXAncrchRdrvuhZb6D9TvC/4V
Ms4D/kQ2E34hHzqsqnLqDHV/BCF8+mqqC//qTz9hPM/H+vCITpHmz6aepxZLp2lu
poubWJtvnnoK9HBJL0DcXNPpYrd+Qz3i8TQBm4bdaOfnegguvwDSLxkvm9fiPvrR
L5Tj7eR1J5dPE90z7Zw5/6QdKGGSJXyoMQ0W+KcVv+qVqbsqR7/MKXs2Oft2baQg
gzbs1ITeSvCUo1mLk14D5eOgIVQxfQ9DsR/HQLiPBLWHSu4CopX7MOwSFpP0i7Y+
8jDbhaQC0FtZwwRcpi/6ASN6eZivcRS0eRTJWMqmUkB+3kmlAAdkFIWYcT/gkWF6
y0RQsQlo3k4hzklHzi3nI16vXU9dmrFvQksNUfZEsHkuTWgWrHUkD/yHpPkcuJBq
74lhtVUnlvJRySETMMXIO8254rT7jxIPmvOK+ymh0Udo2UcEjAvXg6g8DwX1NE10
2ODMX5GhZXeRHDAjeaLyPIGc6iU/8O+Y4E64BE92erQmUnsZvBz0FwDL74f5AFpf
+j7XzhBVjLcQhWF8qH/dg50jX7OPIE2w4VDaNGV8Ba5BLtiOqk6Ua3woUgIYlCot
o2+S/Y6AezGxQgKO+mj9fuPn1bEeivOWr6/mm1dle/rTCOVRc4/yD0jcSM1wNiM5
ZxYEq2cJNo2dCYMy85EBPyb2Vln/Tj3msiD4kuKeC0ZShVUeX1IogfnZCSUe8YrS
CRW7vYYRqNioBs5KAx2zhbwa4Icxse8BTkzw81akT+54+VI710EbM2zQOCbKg9rC
6ryJGgfYm3Grx/kyav1cmZkindXpBElRLxRoRN2sOgHrP8Qsm6po5TeOeSq1FX3V
iWnwPlOB4+fa25lEi8JXKIHJcC6NDuEKyD7f3OlMaZUBQFpcGBTjAm9cbIrrlgyS
tnCjyNV7XQ3DN/wP32Sdb+ja2eupYQGWgTR35JPmYYvjKhWftPMD8R8ETgZpQ4Yu
zQobxYydHb2I+wfVI6SuJRP3dxDWwF2woBvyOLVdBdu21iRDpBt5+3akrF2Mzq9L
kUwLDQm5i7l2doVYMj7HDMuQZA9UwoO7UfeE2XPB5JaZYj/yx138IOMWOK8yGbgu
j3fXMXzQ1E71HrhFoEktmAnF9GQmtvCmnkpjDz7SvIcwFPX78ZvAFLJo3onS1TbV
B4LDMAJ44Rtjm8w72HKOskNuZ7LDLKT9AM9qN+NQQcI80o4unwuTZUTTifeAXmYs
KWsig7yqq4FMtCcMoB/gNkm34nVbPIyOzDadpnCWYZXfnBxBf8WacBe+oPxKMCEs
cTty1lAY8cA/6u+cY22Er5EMFfFQRFnyPcgysf09RcQhPoCSWjkTbcoGCpHNpQcZ
BTYfEY1N0x3MD0dk1g/gbok2j81YbcqMPCuRc6qKjAuSI5CBoGaY6JHeOGhg+9Kb
k7DDbIRQMxYwTtN/x2J/UvGusBA5SdDHmRpWq4WmfNcGVH97G001yEPnTguMbvaA
mb4JTeusK6Lg6wCqMbosFy+qdZc3nGoQW2brJNIGy2gs/G64YHokeXrSlTWgPKrS
Eo/MhwhtwavhvVcLr3R7wBCPwJbCk+s+2Hjv0O0e8OQCHezCy1Z6F5CVNktLDDrW
3FEQcGbAA8BhNI4GFAf6sJkPSAaIIieQ5zcxt/F4gn2ZiUcQgAiJUiN0EkHuh7Ya
1i+QfjRfJsSWIqq/1MklulemQnRd9VvEDk+zIEO6o1j19KO4dO/J6YkFCjAVuvUl
e8nBscJiLRd+5CjQ0CQsMva1ITX2IZ68/LQ6aUeJZGNzRdOL2zLEbWRda6kuumbV
GZWGRGGIO74DCMZiQBsqNDIrFIAsX0ym+7LKVhhviJj9sPF+NIbkkVAs5N5m85IN
FQUrtZwgN3xTijpwaAbX54RkN3afTDKI8jqEQqTuioL2Jv0aepJh3GpNUgB+O1aX
AT5fjspWpaipDc4d24pJyjnpFhewPhf4D0eKEHgfLFYNpx4Kx+XSroAB3WH1zKMu
UlEyoibg26p2LoYQJW8aaDT/bLqjZbeD3QRqtRW7Zbzh4XwchOKznVSUaJxuhHxp
G0d39mUabMmbtJU2w8tY9z7hFoN7uPzg7e72nQ+iRI8O+TiWGl9N2U3CMN7Tw6L2
1YdHH+KLNh80AqgS7twWa2JaY0EcznKXPj5bDtjLtJO+Y8g8IFwzToxOm3rSUb2P
f48jyRddvBOoPO7VkKS8PKGG1AnNu/BYtsagMm7xeAICQbTW/ePUu37okmOpuxpu
1jUzkM7lfdgs2FDC8McOgqo1yBM28BIZTpIbWFD85h2Xk+EdvTLmX/TMJcpwGvZI
X3zFwovTRqGWOTUtupCw4iS75aN1k7neWRa1iSi3JKLfi2wojjiYuUtp789OQxTf
LeNJ+m9CLy1xLMEo2knoe8klB/w6cpt0B4U9+C2ZTJlygS3thnRoIKXPE8C7RvLs
SqhB712seFoBrwT2XN9Mu2N5q0DgeaA5t6lX6EcuOHoWTuQJ1qumJiJ4RSH6xIUy
yG31mhKNSxdnN+2eFraG1G0/t7su/ilaQh4Yah2Pha1HWQ9gEqGD35zJ82EF0lmE
ddAcdm+m4PW8obJUk0a1zFOKH0vy2wys2iXiuuoFgcddjp4hItC4LVnLf0v0rvwM
xN4rm3TvJU7MFNv54cMuJo9xUt/WCfuQAVKgY4iVbxq99ouw+dWWrHe6VE7ls5Ee
oAWXXyo+ADF27FFArLnMWrkLd6nFcKyOOF5rqDVmFiQlmuj32e42iksMK2Bb+/WP
OCBgT9sHTypmJoRtcWxmJFcVasarK2VW9dqyGls4XznevxvOPrjOcgcbGgz2wsWj
JNApRjp1DTpYqrNoqrClp9rJXNV3jgmyBbE+sp9rjNkPMupZg6LijNtTjGu7gOfp
mFLPI2WitTejqeBNkb2JITzxUCpQyHd+r4lI5Hp9VsC7mQXghOZi2i0Yby9f6Csm
MsNCZGJ7ghui3PaOY4jQ19ruu3Do9dgj7ShFdWtzdzHxnmJnc6s8sel5vW1GE+Qu
SV6sK02E+Ifoq/aWjQwZ58kyE1N7hq9WyfFM9e0mtjg8noP8fvrllTHuaL3bCCvn
4EvbuhZk0bnQH8iioWMNvax2LCg46Wvmnu27pTdZbQljZnSghwGi6V3RAnHuPSNO
pp/vfox/0G72RD93384ZbTVyft6arnrDT1aQIrMJ5O/YToQlgKPpjDvPOzm2OCYL
ma077wopRv+NAG2UoL1TfmWPeGE0jhSSzuXjMSeghbHBok/zwVYRlPPtYlJD1/W2
yEQyIEMUqWyN17n3jkYM+2iFdb2rfVYLnbqrKjn7aNxUfZaLPlrhstPg4BMWHspZ
FFwR/eeAzTsS2ADQdvEyHeRBvmTrALhYPgV01fikwghOMPVWWSmlsFVbCed3TOXe
MehvCo/v04OYtZ+XH0bNoyC/rElHMZQgbK0QspI2RGDa685qKnWmcdAmDK+g1VTl
1ErjEHs3Z3b1mj3o1SVfcPE8TAGRD4WPSSb6oTAwj6bZDj7rAwBWXkAwrh8gw0bv
D1VHe+1fBdNkKVq6pK2ueISf1le7qpXm2BpjCxLxUA6QC10Wuv6HbRowxDHzt/fk
O58DpM+YBR90C3U/8bkEXODQSpLbBbjmWUwVmW0+vzZxFlxc6e9t3BC2xOI8FZHx
FoX9FdD2N6Jomi4Jxx4PeZqg9DcGGWIGGHrHE6GGDo1GitsrbPK98C6P6YmJTVrv
hCGxl8OIRt9KmFJA/7nXH63kMA93r5xGbswlX3xrtD9zs6iem/i/w1w4kdClGRd7
qVTmmv3m9aJvfbZgOmYSspRSVgeXw/u+5Mqwga2aonJmbsPmBaGX9NWHq85r7A0T
LbRVD3OHRo8irLtQMfqKsGOyVqdW4SU8vbq2eXOjzENkyS4H+HEGEvvFa5VFsgG9
JI/5IJAs57p6FI8meHA75VN7BM8b9nweJYzxfsFTW+TZjOYQ2V+zfguWee/d71MV
kLIbe/SvP4L9vB8VOwO9SANYUsKbknITqJkbNsLC17iNHoaoxqoPIvberGP6udRK
0umT3QfX05R/g5kRAhUnHcZ3E0QXRjJV8op1CN7N8QLMmJPkFJNY0uR+yN4YlKIf
+Y3uDht9O9IxprEZGHfPaQi3AjGRc3wZ4LpQz6G8M93qBjhb0o8m+Y3GSp8hvayY
8IzWY7YJVUX/vSGUhJxi3se/OHkhu+CsVNUaux4e4/qAxLCsLCOk1YzLRlowCICG
VgLW6BjO5dvEcmrDXe+HNsLB5jJjyfxiZ6CEIdmfmYjPdbfKusVGiYDgGE4oWAFn
3jwJ28rfv6HFHqiQJDEu7hCtoEmXhZ5GhJ1xiVW6mn42yZqGqOmMm8lwBIa8Y7AJ
duQpXS1S/UA+rd739rDWgkNSaDeMnvGsCS5IKxjrc5Wid/IpelIXLxT+c97IT6AF
Kk1IRoBnVQgk7erke8LsPL0V09l51XuflWVefVquKnrguOkhvxzECl3HHGL2qv2e
dFF785K6lKNHJ1LluMlILdjDOncntWfL4dK3FiwOSxrKqwAuolAuz0E6zejdc/t+
iCEkP5f6frvU0DgniVMd0AUBzsS7sYLEAfJ+JT8F71OBY5B0zXhDwm/dSWlE0LYN
pnPlY8fQk25/CWLaZSZ14/XQq47jdMiWb8JSOLBYMPY+gbSoJuxTEYE5zWHYqkhH
FC3s+XOgyoUh2SG/FjgEnVkeFts8/p8uwHa5EdyNgBF11s+ZmLl+mXHMropKs5+s
v9Ctzlg+iyqyNDPqrFl9E/eI7AkJHDx80+/MFCZjhFn9N6v1e2Vbxnn8DtN0KNuE
XumverJcRcGrs84bZzW7xBOTzEcMspKV9jG/MUCqgDP9w2DDw7uJzaTRrZUuoJiN
MJU8fsQ+VDv4yHBcNRlVg/zqOVl18BkL9mKldi1aoYgTH939FxuRRO39k9wSdxKN
QkuEY833LM/ZPch5qBapP68Pr5BKYBb5KbUkL2rgQUn8ln4yxvdQaSjdD4uEjuzl
U1nCysCSIN87H2jONke7G1pJZGI+e+Eb08TRX5Ab0e8yxzFoSadArUYwSeCRAXo6
Pe/Jv9BjiqPfXhxlKYCq9HD4Dg3s48aJ1OIPP/kzstqUhWaMUizghwD2mwKyxuva
bHRlG1VO3Jjs7tVi94TjIZ/qu+ry5VCOsjbQyPA7fCgx0vZLr09D8hXKNSK0xAsg
p11L9yP6YhF7nBOxCsxyADsmMdJQsi+y9xTmpkNKlZv2S75uTVaOM+cvy1TC4/nQ
CeOiKXPjx0o0d3GYJpQCxQ22wfhu4uSv3ILzNfGQRS9vtJOtWiMpYr/oeUjohCOC
RpzVWXRC8+zDScYC3YE/L8VJjXCRwNhAJolveu6V3UW4IwBRMrdu/51EKsiWiJX/
06vvNjncBW+BTZNws4DrWfwdIXthVRuX/jtBu++X+8Qqt5ta6PxWh6kgfTZoHtVF
kaLhos02qHEtPCY0cm+y1n3HtYut9U7/Dg35uU+QQsOzSbvDxzlMrNBpN9YMJpAF
MnvHgiRcam4hyrRxHIAVBbtW+fv9ya1+ds0FXHjhU3krrAg5RxAggrX/3qk/cmj3
fxQHzN9WZpcjLL7KeWUrOb8IB8o31GdsJLdVIz+hBkn6f3kYk4FZmwLYE8ObpAgs
hfU2zLA6fgrHMyockoyh/7hRah4dH/aqRfo93ZYMxp6qIYduYZfHXzHAtw4M1cvB
pwOkuTQi219NIQsZylZt9AcaYbLDg0Qx7bKfmLwEXWS3tZGL51J79g6APrOlytmL
utAP0xjmD0tPNTsFFtc+CJOf4SHeDzRZztySmHrWAeTpIGgFHo6IFz9Onn7fj7qu
zsq38SX+ZgDBDZLLeiLkqwMPiVgtWQYxAzY/Mq+i0f25Z60SnJ1BqEjiuRdNBEl5
5pDOJtGodeJnJDlSIZexVdNNP1ctRBheR12An+p+I0OeBMPXxlA1IJq+0TTA6kiD
4v0hkQoTQYukFSf9TK4rx7dKxpeFQgwfQaCH/8A8rWO8J6fLHrlaCOmLo8O452Nf
AAMCpsLJBkNDvHvlBSmS60avMdK7UAClqu3pBQl/oCdcpOBSGIeKCFdJXpjbkapS
sXP6E68gqU2BSxd/6HU94pnHUvzIdnnomh28anTMep6TSnU2jEz7KGloYF4WuCZu
Vt5OzKjMtYYK6HVZNI8vc22HtJc7Ie/4goC4Yug5pyl0w5LWYYSeq01V65QDM2k4
eALNT69/9nyUD2WBIDs/PfqraBfjdZsLXtnAY60m/NqNiPGfm/hJulY/braIUBRP
LIQZXYkaxppD69K7Uof0AFwLS/qHCLAJit+1q76omGjYKHBhP081tcI9Bs0sYGMx
sTyRn2yVoA/kaO1pjxGAHQzKXpVHXkYneb1FnZZrC7eMJ8SFmFIP0aV1wTP6oD1l
rqCbNvsGy2YTQvtjMq6LN95rLfwBf1jivxP3t+FfEo6i0OF9f7buO3DYh6kYApKf
GAw+Y89E5wNq1M4SsqcLGTqh0VzaMlw80CnglGFYfH2KexJ9tQf7Zqzviy7hs0tL
Vn1VxwvHYH7YNW66Xv+ziaKRsTKAnCPsx9S4t67gkXARa8ivE8wz+08noVZYdsXG
C8LU/ZhQyjdmECIS8H3nze8TtbBbkCFGGbClRFAp8zHmJTetGv10Qm+tBL+j/xuY
qvjYH8ohYaO/mTEeVc+NyEzEi5JPEcswW5ZAhweG8Rj4NjuicfGUS/i+QotSwhyO
K2Eck6E3IRqI2y56fvt15D3ZVTb8g/ftIouUzApWm8gcXM4gTOX1u9uwUIbkSA97
XZ24jvpK6phhdHLB/e5hBDZHwqA3DykmJH42lVvHMTIc5jStUcbLN1qDnMYX1ng2
pvHKQGK1l0Uftt5noVL7EhBhF5cnr2pBEMa4jnkn4vArbzAKctRXWEHxQII9tUkh
M28BCkPc0Dbw55o70hemp0f88jNP1kOIriuuhh10pshMPIByPC8A88gkXUJ4IXSI
jPt8dD7OvFIISHx2itdDLYrP+UTUqG5/oQZOho1PJkUdhnmuNncVoHVYI8sA+at5
LpLy8s5ZwA9UPSl5fJ3fprTe2QyeQUv6+CiF3ycmmpdluRWejj8RdV/UzDrGjYAG
VBnPvZFKnQOkJ6xt29EYGKqVQ6WGc5vRoyGIE6tYPDgsxIeqraN2UOdq2UtphUH9
JeYc1KLAIcvBos0tR6LawhpFzzyfaIWKexmBasf7P42ysNO4lmAkJsYKlhlQZ++z
bLCQ2Um9MMi6NF4qjjH963pPHEEjB93To9ZVm/4Xe+UFfl+NmASUJy/A6s69ds/K
mfALudUZIlXiHORtbQZp3zJmfbs2jWn2bOr0eCOBLM5PwIH61/7Xx7Pgy+4IAwDo
go/jvuaOzejjwhXYkCplDyqAgcFc+Ba/XkWXlCuYhmHG0oxeGFeQqwd+Y7epPjP9
mJnYO3aFBIsrrpGTsOOaob9r06GiPsQPBRqhUcLI9c26/cOAi2WbZk08z4/lHiv4
ZyXiRQOhUt2kNyyHhYyEthcmCwg5Pu2W+AwfdQ1EFiEFH7ZAU2VbMEfjW8+bU5H3
h+1dD4xKuguOcWfMLxpKoNzvrx2KpDoZmFy4UdrS4bn9xinrsj+vCRIF5d4gz6Dx
HzmpTjQ2fGTSqzW7E6GJQ8siN/G4d9d/wsYO51twFglzqJgcZdX7Cy8mLUByTzhk
tjt+rCFHpztat2wJ4Gi8Mn7wW5F0lgL0l7Z661E+wRJq2kmTaFSBqiNUn+diSL+c
/0EsWuJDaj3uU+A+1iNkRvVp1o7BjfeWhJZ/grpWYR6mey13JpLtRZmP8kDB+3a7
/dcPktVteua9W+HS0Z8/saIWZzSnRHfSS5tGKUtnICMNJXSumTBkxGKocgm0OmXH
djZ2yscrS5SesX5WMY0d4StMbsQk73AbmxQ4pGnouiLwI953/kgKJMoMS6oNPsFW
oFW6hIBXC3SSXy9MO7O+uJ9HmracDwN8hUqm0R31Cvh+FA2uwqOXSdeR91MtJ1PT
MPi2Cz42r+acIQuxP3AyKVyYHSyKiTpkNazbMZ+NlYz+sWhb+bBOBK9Sy6cnm0OP
T5CnbWEryrNPWRppuSL+fjshQrHLNWwGlrkuwgAu66O8/VjKHcpxO2rHfEAF013e
7jerKcUtPhg5f0IevIHydoWOyflsrj/ylc/zOXRKZIoQ4yM5TahzKjflXQtpO265
JOrK0qg6gYUzg+Ajkj+Tj/hlq5DtfpZy12rodOvlQ15zkvq/Jco2HBQ7/WDKyZRt
6qgcnJ16Hu38kdqM88G9dFZEZ0LgZkHAgWM6VoeJBnJCkMeTEbT4NPiLxaG+1sSA
NK/bv3LbUWaZoekrgash14DyHyC+KANHUz4R5InM0MfFL71ws2YZzAd9Xm6MqxU7
vRIqALRSW+pyZgsGsthkFDyNfb5nRGx6OQ2UddU1DLJNMSrR5y/9yAn0yF2mTy50
QUQzhUSL/t7Nx7PxxJoFcSMQXWeDi7+bvIAuS7W10IwKB9qqyX1yFTHPo7oFzJIm
rqXmNZhZzy96iLQ3CjVtaOgVg6UEkFKcM/4jq7jFz91nrX2TSWuWR9WEr+MBUwX0
0y2NdjeMTQJdEyWBZGnUnjGBrgY8N26RkxrRKGt+VuBGNyQ18Vjw9ifio8oEtsFU
jQ/oTNI+IOKW524PQ157HmmkgNXg/tVmgqOUdfMdpH4fqsdglArxhypvwYgf5RKG
NgBgbYDD8i20IrvRwc9qkudFuLuMi38Y/B20Z5fLnnBUO/wXDjESFnWq09mVJNKt
2y3vyqAoiUyKy6MNWH8AG4vQavO9HwNRgv1YLN9E3mjDXuOp03ygWyyDodh3T+mH
3Jtc1jJZq+CUVa6YA8oUPvwG9bfFhfOITQ2vXiIApLqgtKYs5SI4PrDNgY3ZwksN
W+NE4n+VoqaZnFxNTOoZVLW7OzfjU8nSri3J1XCPss3o5j+yokIx2SIfPP0dXMjL
GkkkJ3eyvUf7XBpnCksEwvzEdKmCTXS8wI9zNu8mmvXHrdP/mjx+n3x9iLZgptAg
DQxkNJ7kBFmNI1WA65k9qpUnmucQFWrwAzgo2TFYvJ9MdTQU/7a4DqDILJz878Wn
EvBhYgYLueCAkR0dvBcUi7d9OxwyrWGFRx2KKqT1hoG3K18t7v/E5iHIPM7CSEYg
oMfyBM63L0S1e1z534zXovyX8wOpxGXSTMIV0U8c4DwdqyUrz8QskcxCsQd1aeKH
LjxRCxxuhRKYWuKT56vxY0HLjwvB0ThCpgMXupX577FzV5RVXNPE7U8o/BXjL6sH
byVSdfkowkg9EbvUpqRRCr0sC8bgFnwbA/v3eD3C5U8tOMPPCb++H1uUqORzFVRS
rle8N4xJTuQY/pOcJglMeynHlcLu00XR0F4wDQElss21h74i/aWYRqa3yBMjnsBM
OdMAFWmyZI0rAXwfAAifQQwESnk5YrwQTMxpsAuMdkp75YNAQwXRdYigZ+Qbwzzi
lkJb/jI2ViRhrywxP1ZZ40NlFqgJTx7Wdk/xoPf4kI+SDEdYjpC9GjU/OFeJTkU/
97flLxXJxhor3vYgaqa28CK+gcbzHzPL7z6gMEAoIh6s7j88b1XRECq3PIULuwWg
WkEzrpECJ5Wnh9EHOD9Unzj8vXyVonDSKAr6DkNQklSPl+qiDAiE2ygV6mDhrWj0
e19CNusoK0niEg0rSUVmn0mVi+1OiEvVdPYm9tuExH/SQDZOWnSFhthTAduytD3e
mDhdTbmI7D71AtraEn4gOufF0rGPLb9z/OP1MWjhwIU5a1nmsFjpD7RNIMsAFUPd
esA1vW/EdBFzWVq0MJMsr0egUqNqAVAqeij30H7QtG0f/6+15sqX2kCeVEUekzub
WcIl1L4+8paKuiuZaR2ZEYvG73XBe7sjZB7EcIiSK1VmxlpMhBiMbB0u+yHR3hRy
Hi9h8S1Ca9T5AFwQj63Z8cUIR6VmT0RJcsP4F5wys8VzmT6SlTiNbVy/+6U2LqrP
qZwjeLdHAVQnShXzPuxAUtiJ5nZVYLwjBkDK0W4Pj2iVUzdgJVz6fFu7/l5ylxlC
46u//YSBJvT9cyka2ZdYIWEfC9hOfqrcF4R6byiOx0oGYLSIHHcyt877ZM3kI7/F
aVTbOC6G4nCFKyO/NWEUDoG9HMrwcohbNjBVYUX26KJWdf5UzmV1Aynokl5NBe1a
b25TzBf4GkGH77YGuX+6Ja9RlD+CpPPPOjpbTM0QmesxrC9pV3Tnrai7KjjodS1A
Z6+whfWfyykKadLCtU4NN/fqDHo28NnKXL43/4R7l40VaIjnAogRNtmgOuVRmAQa
Qov8buu8fjfrcvcIK950LNtp322FxpTPr+mNdrn+PcDatsZFHVB61BuNoNvVKYEM
MXpQlq0RSs5W+CZqXbg+EEe3ceF7ltO6dtDhydA0ph4FdasgEI9yk4Q6OdnNSTHZ
v2SPpYoFTXzN8kIZRuOl+2Kag6vibIyttpH+vpMhcZ8dxkGRrqGSxFaOysNkfFHM
+WYl8P3zAztywuZtk2lT7pwC/YgaC+UBSJFQLeZEFM8joy0Aa2+WriLf8MX0O8c+
cb+3PXHnb66L4na7tieIfOKJtDxpVoK9JMjYiGsIIEIcaxgDdtYjeUDWEUFv4J3D
yePS6ZCixqLWvpuubWU/lOOWSs4UuJ4sYWCsIzsR9AUPBG55ows/b/urSbEk+W+Q
YFmLt9bB7NAYpcogaVl0B5O/rItPReJ2unJ/8KalOV1z6XwACHtKfJed/9lOf9Mp
+rnKBP20ukiWmGc7cCPFcGDa9PBM7D01xeKAcLG+DZRMyUycGevmIDSTVy3iQWD3
sFsc6SxdRCqfZISloFt36gX3zQjPVkIddsGdXlVDEiHEjTEoOwf43A4F7GxlBpm6
43t2gDnY96FRw5WOfyTIWr3f6WPUFgI2qu67RI5XOQUhg9VsCC60p9b4K+Usv9uj
JP2y1RGD1tOcgcGq/AiMd+hwHanNCUaSsm7UhFRDE6NbIzLRhmrAjFtFva8/Bydl
Q2jxjzOeNXdozhObk6sKuDw0s6UW36jGvvTIlZWFSrXH5xWGrY/tyXE0ZBRGwzwq
nQkN8pAuNYwyu2JKTwhYYO05h4TctDzqO66IYSQTITo7HqRHiyIylhlxVLJ5H4zq
jdCzbobs0Z8pta2FZGB+K393E7hIzec3EYFb4IsGWTTiBPP5f1f8ofZm5rv0qw2y
SW988rba6u5N7xrKx6x5gz4+GfkU9nTyYy1WCZxQ5gb1af0YjFDUOy9orLbwlRz1
7S7wGlAHSd4p5SaVBwVOoRd8YtggPOebq1KG8gnYhO0mxVuXRgNz24O34ZXHClxq
rOU+YXXtFbIZ3lMct+xXEesKfsiTkAMj5fsFjUlZG9R48mlLM3wsqaLvFEwfW5he
wyNjrkK695Xyc3o4y0obSoUzJpNgO8ySupTn4MWvZC88Hf2R040pd1FpNjSyG4Fz
fxAXz8NaVFZWdBGsHIXa8hKFqfb5fJhsdiKYTeW8W1rYPbPTJnnk5I255NjfmL6N
+J+RIzyLkPWFcsI5YEq4vQm7btWj7ybV6q5FJ6vA72r4SX7FPO2r1Bqu8IGTUD07
yfGF1TghMYLL0GTlKr60GtXeWizixhTvkg+9ArfxS3T+Qv6GUaZqf9OOSdzixrVm
rj5IowiXZeL4QjmJk2qvB6tSIoFInIfN/Ul+hqBQuCcbVi0yMMAzMkLGawru7UVT
KHkpKFyf1zV2a/OeCuFWf3jWcFjYMV/C6LBPzMwXNnCQMdWC5xPv1ir6WzyOmn76
Iq2L/i81u876MwnF8QIvFT737XKmzA07DCThrDnAIu1gDFlFJoh9PjMQagVcdtOr
JUtYgMXIUInvnIFhLHqPzzkHqwvVq+S4uOLWgdbHLxYA0ZVsMfFyb9KUFDfGVvnw
2Vg1UcchUrU/h6JgS2xisuEKCvfH8QvWHKCMMCSLHUeJyKm7jlB43khWbZE1b+2c
O+5SMvmDGQqz+XP9Lh4iIbMCLTe61yWr162ohlCx7Ug4gDSLaW08Qu0YQ3TitnrE
BgA5ijAfu89Q2wLeu8Rzjuh0g3XBdiU92cQtCoOeENdkXemoKIO9povIRlGM2/Dk
8IdZ/EUPpgS8+CxdHKHjHSazkLk51/8P44Dn1cOGwd7jRR4eTdq6MpJXKzSw9fZA
4RZBc17C3m/4NDa+kIimU7//nM9an8IC8c+E1FBW2o7vW9gOKB6o6nM1yZLtKGtR
o7M8QLp/32X23T7aUCemyHnhs3PdJ+gbyQ7uDa+egqqU3MrqsrrFSJbADzpouMU0
WCbqrUnOAMy/ZSvGhfTN0D3aj9k3FDGn1IwlLU6I9D45O9eQmUQozG1XylNu2U0h
tkH3tG7dhVxB4uerM45tz6CAnez7KhCy91olxVRHycnB0TSmkpU0Ky/9ZMC1etgb
zLI9aM147uS0mkltYblUWVNIwghuJQ7MRMU+4ytpyuE+MBNArziXXwGWDDjDCsLg
Tk+GFd8JYABiJERpwomBahWzBYBPNYrKaVMleZN9xv/ymb4rLYYOmkPjP/YboUIr
TePcCMg01r+3ga2tPQGGxmQ5kftiJKUpP+4zaFdTB2yO1TmsAclEaXTAXX+OBkgC
3UBhJVratm42ckeAiTwvD6dFjKh/KsiaSYIBUZ+zYGWxHO0hllNN9AUm6GlRDUiV
wsxpSCpKRymiDK3IgW13IvFnLq6ZgMb3hyjpEkw6OWuHWu19qs7MSmwa/h2HjyQ1
aOSbZKbqhE3dWNOxS6DvdAlEuM0m8FwcDanOkwKxQvCE1UjvTpeZpInQ7eSwCEdL
uUjsfOJSquHqFTMprmctEbIZYH3gzBwYnbj2fV6304cNiAMj9oSHwlIni3FL74HX
9IOuTst6emnTFELWk4FJd5FQ0SmnXkusuGOBKTHYI1e6EVXJhyuvncV62AmjaIS+
ZMpD4dZOC2+lrgEbdMETspHAMwIUQyi83fFjIeF+I1234qbyPPquEQjvHsu+0Xby
QwDDnqDn5ReOz165qt3CoF4GixvmtXQdr6fdTY/0Ey/zqrzsZQoU5cdfj6vISUWo
iquCmkOohYVsbKy4wf3EyZ9DBNv83LoAYe/wtL1DcCKaGHrcvcA7isNybUTzWNbG
8ON/iujaEJC4gjKwSyEL2lnm6Wo933d2iell0Xo9C+kK5VNccZQ2m1oXTZ1FGLUB
odggAZaWXvNr+7oajo4EZBDNxPSYPTRnGEmx/HGzxIrLQdGV1ohMl5Ss51MV/dTx
yAY0q78AiIeKCwsoOHpQldoyJMJJsCZSm4S7SPadSG/wf7vvgMszfvxN+WesGH2O
ox6xSdKFmAhHIKswXSq5Gb5+8gUFwDV57cYaaUTQaVcV4TxoNUksbZwnwMqNRb5b
i8EpX9O1d1sLL89GB59T0wZnKvnJu0GR2NLb8DYrL+Pq0QmiBnlnYW29v32sLNVN
CoaGCo+ZPPianeYuc2DXrg/9Zx1feCNqPKQlqmVrKa8T3XEA1Qz3jnkOSvUaL0vp
2IhaKbL2QAKK9cwp/SRRFrbPwgSO8I2/L7YwlBP4XC8+6N9U7dINPjSgPJP2Putq
bg+tyqZT0ukzXBMTVU0PT4/gRZrPAVLYgAbeP8wHBYIur4TnEaeUbnL8TqbEeZfg
44wUFfv1JBQDxxwybh6N0vRpqgsaFT4BAstm0F6Y3Tdn+CZ5Ni3nF09zhwdeiGoC
IyP2FmUvBs8JmMKbnoMPa4WEKsMHnmTaOc6fEH5QOaJ/EQiDucZVToDQ7O4NXyUA
Hf1BrLGifICILgP0qV10WnfphFOMHjFfLuM4NiZ7S2YTkM+m1LeMcvVMl8vs7Fce
UrEhS9Zv7oCBPjWxX8bT0PHLyQifPZcMgo6YXKW8Dr5AAvB3YAywZ9ypsVXls+e1
GqSFxEBe1b7RTz/iRyxujivXCU36KU2Z3q3QB7u8U/LiGA3UP0ij6cfd7QprDCQ6
vZ/ZY9V633lbhKACri4bbKxeiha/XWPoNT9o1n0Tkh8B+DRwh5Cuxl0RuTDphhZY
BzdHUx7QiAA94qcnzZNIBsaBRwro7EaDkUE2EJVbrFA/hxBOKJOlAiqn4pmDWg80
Tq8SGpCAxtfWFzEbyiayscXFXGCAAJFLo0Nz53q9atEilFE5/R6olwe8f4B9dVL0
nk+LRBLB54fhZm0/N12/C22M8Csrm7qi6nDSJBi3iykS1u5J/njNK7THLpuY4tHu
/KaBvulzAVqnp3zptEiTjqkn79GYWeARJLss1IJVv/ZSmalJeJVsSgT6nlCmfxlE
Z7ItY59Hl08gh8xhzX/sdtMWsyiLmzDahvLWSwWTL4u1/8M6gqAi3eNc6EzbKJDb
zDtAoPdZ1FNX+59yQQquy+PMOJyt/icWtMUUsqLBBHsSqQfl5nbzvUH3QrmHRyXu
POMwNFFujv3R7WKAvgKgWALTNtNgNNOkD9JGBldbMHWkqd1CReH26YfyO6ccUMz5
kuB/iCEfFWREKRVed4euYyqhRrRSNYw8fFB+yMa0ZGT8HKmfhzY6JC6RSoeq0yJ5
fiAVADGqjFNeaYhLM4kInHaEgd9Wk4FusUm0h7uXfpfKcrGC+qA4zaIcSkUIVdlp
I3eziop0FTSOTpPEcnoJn8HmNtLSb9VVxr6tbW3tuqdTU1FeTiCHjNZeBlz2sXj4
pDxXdfg0GQv8dVC1GsHV9raYyGECUxj4DrhUk0/g5hCEbAOEu0tUeGnEeiLTjJ9I
/zlerPD0PUlODm5PyRN52F5i3LlZD/qBRjRCk+nRiZAGSWcWkRYq+AJji3Ye110V
KQ8CVaBIqzRRmNNdDRolbcRYz3G0TAAZiPjz8LeL09RMeWmECCUyWfA6Pw90ZtUb
7gErSQuv7QLJo7CNVgiHvPUeQmBRfHSJx3JFPoHMysvILdpy1FWpoKL8nGQzBLRp
OMF7wap8jN1eLODWfeIYhIQ3W5HJ2tScRI4AcJ14Q2evb4C1qsAzR6q+INIO2wzt
+9P1bAfEceBIqsRxGR/YNu1FtY2jEnwo7i5Vgsg+/KJq7N2OwlajW2tncOAHNqUd
I1r97X90Zs7d7JNAFOtaqsvGeosKeKz1aL3yrLIvIGNOHHyzH3aqF/3O8tudKh0m
rkfEdLNSMN4aArOMiuGz5jU5eBmDtWLHThLfXl2U4AXlN7bOiaPtKQQzoaftF3vS
b0T8JgnItSwyEvAT8bhbLKXW2GsaC4+xBAvP1gAzztlSpb9yIFnUxFG35B3uGOh9
U34LlEW0pfXFDfOGKNo3ubU/gApD6XkyL/RyUWaTaW7uU0tLgYV5GiHPTDzdOoS7
Z2dqN/eLL70JcioTk4uzbDdbnETfK5BOwRkoF6xCRA1udvupeUpCZ9LwltTde+02
pEHQP8Dj4QeWwuwPUsZ9/A7GK+Vh5I6yhduW2kjr/36QmFYTyHilLIG9LPux3e1t
53P5huUmcZpLG0TgCfQkiiA0GSe18jwYJxyszbhYVl91mJJUU2jPwA+9ND7GJeJo
q3ncpPKY6aR+S4qwm5s/x2eB8BJzUdfrVMB3wz5FaviUe5nUyQbDktPBKKgRwV44
R1b71jtxaZOH+oqV3zylvTTkys+r3zM14eubIontlRxEGnmMwHUXiQJcJrPbjF9L
sgaxxMLbH4nTcW9L/36XuPpRVZ9XJb0/BuAcHBmjUzo0+GMuR/hWLGV9mGt0iH32
XCztH8sSanJUEW0VYPlBW7jcH08IZ69i3L7c+jLNSLKgvPP5lfwMmxh8ZCKhJj69
snM/IAXUI/QqXjFQAQ9LqlSbuT0XzpEZA6DT4lk6F4kAOzTyeKQUdmIyAVNn4alN
Usa8pta2u7GHYzZakyXEiAieIXsCxkah+4BYnXqjJ0sY7FGoVRhXrWP5p9h+L7ci
dWiuUGKhfHYiGNYV9sqL3IvSXoNEceYt3QqRoVo7NfTJpkN4yynK9QJ35Qxr2k06
fBijYeUPwSU1TEjodC1dg5hK9cNfqMGu/C+l2NITOKT8v0+s5f7gPCkOGmOC8U31
lJfItCv1jNTF7z1JEpNkyzgnqffW7LsaTL1fcUd4gyeBUM58mM+JRFwnJKt/3AxQ
42nXD6pXJOXOc7fqNg/ZXzMqdxh+oO4Xs5xVZCyenWCC6BBK71bUz07ykrojOGg8
M4NtQER1ygifhH3EztZom9+BbDKWB0x/eXR6NxSaItosiSJzqLCI5xm17TzLgSFn
5AIsK8321I1kXBcaRnKcvB86ieccGGUPhNh3/w0KMjbv9CdjFfNtIEGZn5Nas0A4
ICHW7TGnEGVhOV4T9moEaKX0aCk0RUOVG9esDuwYhsugm220wDqcglJw+IZdXIiX
CiyBjiQ7e5io5pkygTRNfsv4DDLHOmIXNohJB4Ha9qYPyFPUyDMc6JL6H5AzGMZ8
bBWcVP0S7FHAabGTzKv1K2W1vSntZfVY/QLq90AeDYplLsrXTY43jTNuB2+PkQt7
XnbwDRjLwFP9zR2R8xMKweKGNQo8L0RGGvNxP5bQZVERiQ4yl/nR4lXgqFH9cNzm
KcfqUMVS9jo8URwMuKj/TxGCOrPSQYs31N2U3qVCK6txH2A+qMkofxcOmH9ERIw3
A9606QhX/kVCxh8id10Iepr0yOVGDGaLn6AILr8C0FhGCPMMp/PM+6AeP4PZD2W7
rXcsA5tX22swPP9UWoY5qNxamUh3HaW6v7Q8IbD2vYesopVm7LBAyVgs4TN/hUpS
Zdz9rEFDHJRQaU1ZujVbtF5ltI4kW8lRMrFM2R3SxybI6fOIzP4HD0CRB44tY02d
B7AHNxuk+ZJCr8l2L3jz56r7eB0B9zA2A7E1qWsdbb2/7efQ836URC3hNgBPez3W
e1FzJWoXr7A9YBGVT+3ZqutgrVNw2PnO2xWIBBdjaraomQZ3L7EIEzfrNNZswjei
DsD7iTubl/PWZZAWw6Fh/aaKptBGEJJtiaUImmAH1/UIS+SqhwZbwFFC/ajkaZVr
fNNJS78jDGQOVPJbi8ma6MYoGBPyKdj5iChhq1sdx9tgTAjLKIWyWRqZAUY0LFm3
P+9b1avTmga35X1xPHwwT1CQrt35sYZ63LgU1U6SwTBpb2Hp8zVFFGoAMjHbMEZ6
LEL9JnWpK7kIvac8mzTYh8CEy/IXabldvOzS4iqAW+bP9yyHUbrBardockD/d0zn
U4jbRNs4Z8MkfS20jbGVM5HBEywheM+KURNOW5fjuf0NahLW9PD8lJbYz8iy02sZ
r7m+ilslTfzpZtR7LY4UOWgUlYxcTzkqZYlCKUSwV0eo3a/HLhzbVucCFfa+T6xN
2MrT87e8uqThKQ8R7nEcj+tRaDf5f6DlT3E9RSZtFqj4Q0aPJecy69soe/56Il/G
PpMqIFXcMHZZZUClRfo9o+OxhH1f5xd/hryxgkaF9QYNfrWrb9gvIkWjfDHxYAsE
j8WT+b7g4Lv+/yunQMZ8RGkPrgWAwhtkUnaAcwJ1vRV1BsvFso7osMWDXipst1DG
QzK3UljEKP3wG3hgTtl9tm0vu53QwMUZxWLEr5U1TjZlmyhxGZDQWilx1XRUvhR9
sFOnRS2EwfHU3OXtbJ761tz1fwPRAVikeII9QlUg9qRH0vGmGwRWNsyjY/7Hbd2J
hsjeS7OJFGz5vfolPa9faDbOWP/DLhlBLg/82ZIb/lNvE6Z3ucK8ISkoP9kEHjne
+EeZCnL1A5bzFDr52kILs7xGMfBrpFLhtaW4m3TGcxZJvxLOoWWIziPRd0cR4dKi
G3hzCp/n0Mle7AV7WD3pvaWEMqBt1ZSftvClGbKRAhI1st3x7uXPHX+qBsmSHFHV
wkYSbIzYa+JsRcSN0G67czcozLxIs1sAg3TlzeldbPtrWcZgxdv6Fv4HPNSJFyc9
MHWOWO3pu1VOIcj/Cjnx+oUfy6IYhI6WFWFTaJpHH9EBGldd3XTE8OhC4/38aXCZ
VjfXxpCprepo7fe+zk3RWYOoLGhFDeV2hxs6w6p3U5o+c5E0sWprH3Qt0AqSSH7f
VPS8xE8jTl11Zema3/WVJdNG68g8iek7cMCNnKzSH1BrIk8DTZuSquGajZG85iu0
15Jc6UTbebxP/u94lZo6VJ0DlrpV1nFYfSDhsJRPQdC5/HNvF4Bwal3FF0HEaWqI
yq5c1P6qMkCHBD+7lqxufg3Py7HefNvwMtLmhUFasQE5+eQLEPAJetetfu6mbGZm
bI1hnyHoTFi7wuTUseKU51zmEBNrCm/q3nd5uZauf+h6pj/t/S9JSTE+WzDlGbTf
QGJ6BWq13qlqSujwRVbuT1jz3LLOCpFV9keytBQoCQqVwsGO1w4qLbbTdwMdRTVa
kfqKe1X5/hIvzmNzrk78fjPiRDzowZJWKrNqGG8pvdfxf2f0nO/Zb38Aw1Xhqy+V
XNgQPfC+9pX7PVuD4eHSXXuV9h1dtt+g8byOsl57SXy5l2+pvCkwKrDksizrz4il
Q/9eLV1fBaAvITnClRxQLmfRXNYKckPvFkrp9mwA4444TkTb6WNON2AH/ANI5LRk
6rTcuvZjd5NXvAyHNbmFSRwDdS9V8t2H78fqFJPXx8hdcXyhwRoXVw8RlGLqnq5O
D2P0acPnDetXllNmwxnG+KJPjK/REvJPU3JGqNj/fZMMgy1uNvcfXpYgrqeL9z1p
1VlbJ/EOTdAIym+jeX2Yj3O7BpkHVZPmLMULWy6GMRw9vUkOjBhkU5T1SLNn3Fyf
Yy/igNxjvCnzJ+uuJ1iYE8Qpbdg7csWwYZLJWEdZlc3v89TpWn9QfqLsR7GKU2EA
n6LYJJz+NfMR2FMGQEY3NFM1QoaeqpV6DFz8tGKwTCEvSWuYXVYbMQ9Ub0ONMJNv
i08CvwzJDD5ydO5chk5VcwKltGXULeGutW2QLDRjBnx9AXzFJtbAF1xIDwtJHJ1s
/WZB6vISS/WHBYc7ztq0hBJpsYBHB9XHRQTUC3VX0BrdQl3vmxsAN/UlvcfKLbHc
VJEAZNNg6MUu+pvnLDYPbb5fYKs0gc84/oMhdgW5+8CsUG8IFC7xZXnYoqRr+aRM
DgHUMhLrE9jCpkpLAU7f1Ic61vOxHo5LhMODQuPNx5d+UzW3EV+0mdW8a7VmU31O
fr29En9CkoeyfJpHpp9iTZuiIIJYgF7lXN9SCXUXv9b6WJAA9oI1P9ENndf7/SJz
sFQh8H+/NjGdpglf7vmIvPPCdk6fg3u2U4CB9SvmkvPCjjKwEfkdyFfaEcZyHtwm
R5tWsKCls2gNk29TkkUJr/VO0OvZo8ZU0jpC2glQGltM7bQspLKQGTECmj4fjVJh
njZOsMFLay7lCwSIsO94ROy+6dHRc2u71HmOqBkjXEFnZwSIPYqEwmbiZScGACmf
7YE+/qTzDAorVLWnVjJi0YkYXlV9jeqXdyM2aVqXofY6halCWXeRqxWET2S0v3z0
EZaQdDg+z2o24x+jwx//Q5fKT8NbEyXc7i/PzkHJHo2932BtoNawx1PqcsZZkb+E
lqJWbsLVaqkYrH0eoV0KbRB7rCaBZwvuSUJKr35xnFYe6tFwr6bfPWCsmXVc4lK4
goRRg5+GpI8RmKSJGIMLta/FToPezpkuq1leYwY2rJ9pBrPPd/uJ5KO3Mq+oM/nF
qXeketNZdvo+1bKWHZzA+QZ14U2Mp/jIN4G0IIQiA0Q299dslB68YHcFI8OOuPsU
xS8WUrJgNNevAHg/Mb/m0Ift5qid5MFOAS4dihK6NGWk8TkQpIeFkDJDmfrV5BgW
s2uSf5Z2YQzjYA7wytdXObDoX791neo49tMYAqWpKiKNEYX4OYqBHh2o8P3kVJ0k
Dz6SXbGTVlF5MDwnI0sHADxXuc2E8rCd+XnIjGWeRE/RHJbp3EUqltEgOgnNEqRz
PDRdwOL+E1nPK7+IS2jiQ6UHXJlhoUaYiNiy0X5eLpamyPHv9WdDmpNHg1rQLBza
7uBSaZRgPu8OmCVDW+mDZ20cXHVsCUJMtTw2u9ahd6RrKAw9evinSPFRLNArLDOC
PGQ9J5br2bQFhC9bqRnl4FtUIJF5EbUmrkmuxzFZk4A1Z+kEeNtuEOtwPRuPsKOx
zOi7/unE0ZH98Rk6ihQgjVU4qBvgksRImyzQahUdwnFHflxe3GDUIih/X1j/BfQA
Kf/q78SfBaLHpjBd3ZpGjogi9QckHcM0y2CftBwZsarsTac17zoSH4BR+mi88/2J
ismaRavapx58H2BijpM3A9EVFczOxHpJ8BgPvq8ErcRpC4texPuOgdVecp9TrKip
v75ffKipNiIkmD4vcHFSTSZDQaz8L10MrOn8oBMfqnt7sJiBWn72VHk6oIPPurGK
r4b9LKAzzE2sFJ4bXrhH8KOl2h/cSzdUw3SbhNmplMp6NFWqdyyOagoG/bVY/0yV
kg/5lgvJ/BzCiREfU9wbqGgsVn4H0/hM9vEXp1d2j/2g5Scwwgj2odqhMaOGc9BR
zz1ALTohB0LLt+VMQx4nzEGUqa1eeEOl1xUpi4CdvYRPmCm+rGFZ9pvB0icNwIki
GqMsfcQ1GrVz7WYgthUA8f1FFocrxE9Ej7SBNqd8arPLVgXZd4xIlG7sAkyezYm7
BVgTo/tc804E9LzeOzChZg/eSMpxYiYxiS8+WJ/jCZrOz8QRmNJyQf0yE/b4cnqn
fRYDalE74xcSHMykbBpbTow2Dxwd/jduQCtjoQMHfOAYS7m7MP+0zqXQG7+ahOm4
6/Xv6Wsjqw7M1tQClbaU6ZMV9bXik8UqEkNOOAT07353lkwSnWxgTpNERk6kXQEG
0n6HGI4DdlxAFwoqKEzkCF5Z9QOu/ccFCnXaPMdZULY0QRXspwSUkJanjHgGEVgA
sTuxThuYLrGFGH3+sUOcs2n8DudjPBUhgzgz9ySJ1K0zWsP2LVILTqx3HwdoGRho
1b688Oy6WROou/3uxAxlvff12m5Jhp9Av+b4nEsqCwLO2q4ibQboUKg2o5MNrsNi
KJhn4aFqQgP6NmGfXYx3sl2BSSEdaTzz2wsieYkkJN1bLvrHyI7niKvwyV0g/ZeO
XgdFIoxGrRcPE8PiRftj2ScOE2mwvvw+1bn0Tt7OdMT9v57SGu59USoBZFc1DQtp
/GbQSrOGtwa5M+dB9WLU6J/PRwaPuj1YduMI2UCsweO6/X1n0aj/mF08mrjQAOvJ
Bs/6p4ps7TKoN2u2g29uXHUov/9g5kSKrJeKaO/o4qQCmpWszG24b+twCIKtY/br
NNdBVjjnawc9xpmIc1ps6Vm3YPQCP+l2aNZZK9uD66uIWmh6CktX80pg+kp6b0+w
wfXyxREltcScrw8I0bQbzIq0HeG0vHmPF7i1dQhTVxBtSaTZ3HrIjxN1QcvgEk3M
CHm4+YNWtsuD2x75D44QyDjE9dYr4k+0MP6Kr0K6jvyHgFpkLHqm4pn8wjWDHtX+
lnylRojwf2yXdMK6c+hvAljTvy36g8hLVqAoqBghurYvZxfDbjmx77Pk0T3FLL/A
eE+QqMtFAryJw9fWfLQJIaYR0tNnyN1vTIucFLZ+ogocZdvR1sQiWKaJA5IsAYH9
Hr14vcQuCvJFqzkH4ejqUBcifGp73logCftw/C8TmCkPWjNfYOelcz2PWu63G5dS
4veZuANOMfF5Wl3sQrmeqgsoUJ/asnwtjtw2ADoJ9/DANhgqAttztuLnmxsWv6VS
EiyECx/azf4T5V31Vizfi3H4ob8+7p2qsBNsjtBxDMckZ/rA2MXIcmgQr0B+1bso
nz9rbrnVsUA4ta6rHozxWktj9X5WeBPuDz68inRgWslkKCu8ox0jEqou51LHBKyd
jerdxMHBtv3qw54TTUwXqk06UBGvz/s2KaE/U0o0zsMO3v0t7t+9m02rubB5mNQt
SSkXoAYnnhzEPwwAGwX4wDRhp1OaFGhbI3TKlYQ1Iw66hY7yci2QLz4094JXDKxQ
pw2CPVPzLHVjcwit0VqJG9qp5lXmF9T1DAasOOlmesWwTOTyejWF4QwBS+oC4Pb+
nUoHMfZjVq8KmZ7L7eePtcXTKmKnJGw20UXCbsFV2Hf/mIEEB5f0J6GO/yaCb6Kx
iC36/lmNLniL3vQtrvMI8hsp6Q6UaIYe3jBCJB62ZmitM1aoXMdP+7uo4kwOXR2I
m9H302hFV153UUG1yZHZ36jDi8BZP+F/eIdcD4fTtXcEOoQQu6pAbDiY4plf+s2f
aEdegpF47lT6JnzTtO5Df5HJdgh2TTgNCAyj/2DsmwM0rIqUSUpcB9Rppg0FowSS
nIBNGB/BexUAsjynRURHWNKcJJlikcN0WISu8/lKO7OYpIo/8mUDqqA3zfKSZLEu
ul5gh/M2D6T+bDaAXOF4esx3KVgxl0mfqmO0YtCed7QZbD6yxKCl6l0ZvJ1bbFWP
BJoip+aZmQRE6ZsER5HBBy7UBd7oq6J+rMnZyXMWat3IKtdXr6WCF/okpNdY2I02
8U7zOcivlUJittRA6cJv1Mcdr34aqRULwLwhNNGGokeh1wROv034/t30LB5lrI2m
a7/Bb4S5iD00D87JTI3Wpvcohr9iqbh/CzUFOs/WW48zP2urgnNPr9eWFk+pEcKs
vG7zQ1VoCCmaopc3nhIu64YfnIJeFi1PKd6eluTfODil5lFb8AprtQk4MVlTgdNi
NaGi4g+APC5EPB8BcmPt7xUB6H2DnxzhoehzSb2Hmmx8bPCatsn8nM6Dv3eK4RK0
EnT3mFC6kg42BwjP8+RKPelYhxXqoILWBAdo0amhMRzGmlKmD73FpUm27wEM2Wzy
Mwp/vOzPf7Rfw5XbE4TXOzOnuxZxzAT49aBf5jRfVa2IJwwh8t4DNt4n3giMPk6R
1l6iUEMKh077ypffRmiunWGuSufkltCj5pjqMnafsnlab0NrrAdM1K2nGNhQMmjn
ohIuxim6nL0MKImR64ZjdGc2PgTTF6YU0SnuvrBYsyoRIoQ30cvyJtEUNEfRl8u9
A0QGjUVd4Gz4a4hpthcoV78XK3yg+Zq5zXPzL8ylodPcKsJ4jOhWMw1rDA9Ndtip
rMS8IbAqChpt/Tzoq1SxLidysYJX5KReVF4Z6yGpMuBRm576eY5OHt7hGFFSetez
g9B3SnhyCESDCpUBQzqH6mNBsas7QOf7+3EAJaQB1FP95M44643BH6aPBkr579Mv
pvjzkvas/ikBR5DvEsDn6uenupBQW122XTHrBsBKe61vsp0vnb26C6UtPD+5YwSm
SISXFtplc3tPW5GSQNlhvUnHSH/9ySnozVACbkLmaLRhKMh1c4wlP8LkV0XKiwu+
lB0KUCZ+mB/0iOGJjLCha7Wbs7dYrRq+baWAE6cWfEYfOZKoMzrxqtEK6j82WedJ
7oVn0RGHGzhq/5Q+ljhAAwDUnX+MmvBaJaZRpTQeswe4EaP7HcF1GBCWFoeHGShx
DuNco/yjzyyYph9pOL4hOch0gVvj9CtGcVkMbEQvf8ST0m26KRfLiMdGXXvF5P0/
6MRiuYTUdfK/DQdxQn3Lb4UlbVQjVQHnuUUUssVdzzgDp+Dg4VX4dYZpEbMJSQjM
wonPUiw9KEZ05AinoYOhDb/0gqxahFU80W00lAWXpdvHp42/RYHRNvk0SngPkZTg
CC9qAMwRYpzhr2mEohbickwqDZl0Y0OOSi3l7HZQDJot6PmKedM7ccL5hLX8VExz
VRO75C3N9/54dgmZTXmP0q2PRPJcoHB/vLMdd845Pp2NyTUvxLK2JMHEU5TJHnRz
PV4Ye8kCMTseXX7/AwlhghhUlcl4vGZuLFudM6zCgEkEUIFNwJxt0uzvZA/WRNG4
ehI7wyvBuZf8kf9rAn/W1ODnCMiqQxy7lFn2lPcLHqohfyvj74lHTO4Y3oYu2BGq
iY8ewBrfNItkfS4LH5YQze/OzutKXrHquUqx7XbKaNij2NpRNBe1drir1DbVD8mq
rY1kvkAbW+b8u104UDnYYw3H5mD7AwdXpb5JH+V4eskmDgAQVR5UaQ/1FJbP7JT3
9OnRb20VcaJ5yYGaPt84E6bW72RiRZZV00foLd0OxXwOWKdosqRLBwWNdl//uJXB
9PeyzxOf2FBGBZKgfZgm+avz5DqGd1F9/hTJslZpHPkVd6/fmGFMNT4xTzx7Z1xL
PUxZgkYbzjr1X2K9HmXbxvAFETTVzTAiH5evcZyrvML/OB6MopfMpeVEYptyWeVr
o1YYrR6y8ubx5tNpUerkRp9+2xVcjOFj09nkssxJhSJdXOAxSNHwUedeb413NiiN
NTaP0jsSYPFd1Y+M6TK3Po7MgyiapMH8yC20SHt432rR+u171yN+mdvYV3OzWgVA
hyUfugO11rHtpa/9QosHZP5fnzi84fbw2DWzW8ZaOi7CyUuF4g6/1LhKgWlQcJke
bb+whimdJoiUQxtnPiH+sUsOhgozgSNpB9jXq0f+NReL+i2D5ubVYGn86IzJDalk
8AaRrgs4xU3MrOk/mko7K28hbCA5xQsU+C5mWWc+uv3jddgVM9IJ6RLV4u2p9w9i
JcwNvVYLYC2/q7kIOQOi/oPJmpM4aRTguKQi4JuoUj+uf0QhguoXV9ggpvmlWIRk
Lrl3R4npMyGFUwTc4uMpzBUUClXq+n+pLsZ8CMFPS79JwGV34hB65ECrqgRecN7s
yZpkhHvTij5VCFkgVj0wa+XnDMsMTTu8k7lujYJfW2CdAZ1MZ+neiPLq6JOIQ0hd
6+gUDXh5kQckxQvtGPxN5/YX2K7GU1/p/AJ2EPPHytF95F4dS0tona8F9K95ZWFl
jHqkyvWa7BavRHmxDONx9SWp/W6EEq6ukUUmg6Fihoai4MJ1hxQ5JpPnhfMbunHB
bBWGMmk05y+qeNv48X94qkcUzhIVea98h11/3MFOr3Hfgbw1LDGXJkW+Y3tZGzml
eBMA36a0BfzwoDRmrQAL9Etu3avGeKA78xl0cciilj1D9byqsX+9sS8bgm6LF/n4
wjVaGQTAfRFWJ61euHJnWScMmbS0ZAX9ocGMgwPoW4LYV7icLrtphU/EpBqWagXq
tTO+0m1JmWCrlrTuPN4PkiT+Lkux1DUZ9b73kIK7p9Y62JVVtavMKHVM9sY3UO4i
r6qs5M2iA6U6CnqatKx/8T06WnBXv1yKG7+TPjFSegSsC3vsabkmukeXacTSwkhb
d+F3llzTsrVfiioYxrChVJpmY2O/EDOeDyN9fHPPN4ZvXOQnp4EoGjHGTRAsJ+sq
4IH4bwMIrL+5UmBmXvsliPoY8h/IrdaCDWfvgdpHHUTglrlWeQCK4+DjCpd9LOrf
ooYtDW7Yg5FVGi3EWx1KmOrCHn+GVvXZwqK60Z9/PTdm1CM4NO0Cv+/l7VocvQln
VZFnnC5woInUso+MG36h0b8waktf3WtjBB9+Wsk2CZoyU0dmfjm9tRT3HPYR7o+C
IIzU/mUgqVRta0mpx2MNNWniKftrtJ0uyOr8drfFfvgZzTX+dxlsJcojXlpfFxld
gahfGPK0+xu2BtnIhccg0gBfd0m0qklSN0hEQjWsA+knO9Du31ekTFggjRwzv945
aFYH92lcMbMf8f80CGBkLXU1INVgiNe0XpWTSvq3v2JPgbFAanCuVC9FV/c/vpQX
5AkygKrxU3mia0ayJGq1Q2fn74c5xsW9I9d7OoV4NhMz1Xj6BFwTPUuXiceda+rt
HDWv1ZBpBl8Ts371QveVtDgyrmBl6lXyIgiQdXW0LPynmoyL6yZqUnL8UkRonhbd
JW/S60QaPUOXmaqVwc7NKf6WbqqzIXYYr/Kv4HBjqWL3qX38hQePBtHyvEZZ0uQD
aE6LYvnsLvgOgM8kj+LRGNRoLvYdU2NVpzrW3PJAsfQR/OVPCx8UCEdcI2JC6mas
tnEbLIHczgutbLKWqac5AvpKeWAocBPnAzQv8ooqR+x3X3ECT9BJx0X/6oamCWl2
ZoPjaIQXH20LWmEgGNIsEw0hLJvul0dxWK5YB/UuErgJSGoYVxFpZh/fewHPauQh
H/la1a4gJBt7HpgXXTeTkt5YAhNaGwEDzaV2lKoZvrS1u2f16NMHWO7+RPGoLYW7
F7SlLLx88vPLPG0SwpWKGHAMCfOgPPTHoHNE7bByhglqIVD/p6I4eNH5iB33xcpP
ZzBo1Z51oXAY64KvUVWHEAKFfDwloQP+B0yI4xLeyd5dEQAR2ZO18TCf4rMP0GNK
+XMBQuPyjjbs/F3/1QwOqGIZD8eQQAev3khHhnP5rWUsswXU4evPHL2hkXdnHe+A
cwsJ83PIIvWDvz0s4IRybZ/nJDOhkHpkICYTCyUZf6kIJ37htGiuVWbFME+e+Agm
QLLjP5efx/7z9g2lpSlpHEteJ63+srBsrUN1nHYtYgGWpWpQErQtIiLOyJh9wh3A
i7x+Kq1AZkWXK1F41+/Fc0Ir8+HWVEqC6AvRdMljEI0iqjMOfZBqJjwXEGMBtK97
FtKdh6SZ8rQLU72V1GbegifY2551ef3UxmSHaMdOMVnb+gS2Q0mDWbRVSh0VZU+R
QNdSxmlz14ueE13+6PPmuEQFe8EJxYM92qziJtvmVpAdeR5UcipEHg7R8HCHyMZn
/2ABGU6gtz71VZvKVfRP6AuPsD50wXxRn5lfNyAr/m784I7YiRZfJmPW5ht6GtMP
/6heWrDyoi8vhU1oxkqsbXxbl0HbWJo11uNcPlE09r6SfGdrHp4fiYKnCPfw8r1O
1IiYIXCgw8BpbBjXN/Nq8LI1DAwwZrBbe/0sgieKAAtekTyTux55QZKfn17uRSei
5uHlmBhxJFGFJtfAh83OgNJyqVphXNvrc1mDuYOZgpGe4LCWiNdlQ+rubFq9ICZF
z5mlE/IUXh3jy5I6N5Unbz0h5Df0wOeeSC7hRW+ojJLtaUA1GxSl9LPt7Mwq1hxT
l5UEV46R9Cv8OLABfgkwXVIlzJUz5lrTIiQz6rvoX62UAtnIjvUIXJAJaaqKQdsj
LnpfwCuz607qx7CXQjLujZvqTvVJOrwGNEJaCs40jIfw9wQYO3Brk6lRIS+hea6k
8/wK7dyqp27DLiYk2EM+uCeh7nJzTqiPOm1vOkkqVtIO/l2jsavksh7XJZBzq0h+
651DtnK/cu1iZe/PlU+1WGW1XaviW5+6zBfDnYRktxxqHT8euJ3vXnYsxywFFXpm
0D7MfoikPjO86J9Bbk/+A1Yc7wWu2S3H9cNE6r8M9UGHynUaNDUqgmGSTa/53lDu
Sgi20lwGrtXLZyKgc+Ej4a8w9/sRdlAcLchEI3y8PsVXrrSEl3XFLFmlRuReR80d
lQP4ySn3hjXOCXZjsRkOnhO6n8ynYC19/OWKwdVdI5rcJasHGwScaS/drrTjUoPP
d6t+rKyP8G/+UrEjSxlMwFI7EmTI+kO+/4F8DizxPa5d0nSi8bYnewM6zl/+zS2z
bSV0RjSConh0nBKqqkoEU0mZH+K7IDvcX1nlyRltabDfOPuvhkI56mKzPCnKKR2j
nEglRjyVdJINW2AuC9kdFRShlscIzv5aE7Pz6nLa7n9pbPltOQRXXQYx4cvxNYdN
p+wWHCJOnYdH0dD2vMWs60vrBfFjJFvgYxwFwkAYOU0JyfDrsC8nvJo5cG0vKQIH
v0TYMUuGjjx2MPsZvvNInqNftNOhMEFCVn+he9iCDHuvg2a1k8DzlrIS/+UZed45
FsROFsEpwI9PiTONIFWOOn4mVf7kJEz3bZdDDR8kkPVi3vsvqDWXcaWJXuLOHJmp
+svL3/AhRY0RgCk3vu+NAeWgkcpEal+Dp5XjZOfeNsojUa98gTxsr+8LMObcrpWR
b0e/15C803WEfYgMJC6VGVapFO7TfriDZbf9AbH9wslz8qhh9y92yM9iTB6gEsY8
N3F6pJjuiKBxYPH3PCuZsgEpnWdOaZ2KneA2J9rYhINc6LclksXmtfnwVUlq+kVG
EnYqwfPB9Z0jDRGooMSUrzT64hUfZeKS1hept2t9xqW/i/kaI2Sy/aCLv6FPjZ1Z
9UnckozR9Cgt6A0R+uSrKcZSVrcmXK4if4i33rSgqRTtPKbsqmTzr4hDz4Zl7+1h
pUOqgT9WCoDFX0p8UCyYi78Nn8dznVFfEmaxPyRbMkbBgm5miGSILBorAzNWb2kO
TyhuPhrLHZWaqckcg/KTktoz9/C/+igr/b15ebIp4yfu/gYVcNQ5zOa+5zsy5swa
s7zqTxM7MMErLrHKWQ6cIU4+hBLGsLXDKcgHbO5kiyxAf0wT3GC+cbJsL3Wikkoy
OQnO+0hRL522HLOnnlZqrQiEf3lMC+cXmWG8FV2SE1ohCJe1IUf2cT37f8ogMmBD
KVYhgbHpg2SRWhj4+pGgxxXYnxuP/xavangFY/Bid9NGcQ2Y2Ns0joGUcbebtVlZ
W8PwgVr8lT27971hQKrQ8uhApzeBy7klqBJBiPvJt+ACIef0E39gOH3e5VU4wFPi
6A6R37nhdXqrYXR6mJjaxg2Z05Km922+MS++ZOHrNMyFFqyo646W9+sFme3TW/qo
/a8MSvnhv1usNn7MbME0fMqSiqcnWOxV4rKIJDniK0T0+1/aUIDFIpj/fjai2wkl
Tk8ulLMaNkPHZBf65VBwYq2Cigd1gGscO+9JLirWGYvP2wDepqhEQhupth4BMSI6
IBGo51yUeZ9J8L0n3eGsLDIlo6L1DgwMFmVSRiAcMoX4QFQMLFKrGPsL5Zo4ezRP
lIYbzgrrUvS7TRbQ/iOFb5IC83miD8HwiFbYTkQ3r+GGGFF2bqK3Lx+Nt3zYuTvx
H7CnUuWzGip5Yn7w1anxeySGQBYzOc6/vmWX6sBFZ0JLAGvgzfItJnjeUU+o9eNE
0OOeTx6bA2VTj4BwS3QwfXgIfDNNzsw+ckUs9PNDaMSlU0S5566HgGb/G9qI3aaD
RBqHXB3gn7H6zHkmfFbKuZdoLdsg6vb+XcmZol8hGy7CfEC9kTRQAoPy9epa0dkw
+8vmyXVAOpDkO3n/xBY9BmTVf24PPVpaxA2fyvJMmxOFOCoz+Dg8QizytY2FERg7
bEEV0iNGgtz2KazK5FOg9pjTBfX9DlLVZ6jVqyXTp/zfcacoNGfAcb3Seq/hLe0q
2NdVGg6f/7Ezw7u6o+8JzBq+4uAWvIOAETIuWuF14794n8EFbLTiVQ6xTmtNzmHQ
ZxzdEP5CKGYC6+Eq2g2ZUCsVbAVi+qiPqk1QhT4hZpfk0IW/YCR9+zjHWGJKRCrL
GKTkkL0t1yE9IHGUCqRYWDEoog1eNaLLooj7a/skynzvjNwIwfLXdg/hmfaNk+c8
V+zHhttuXFttnjyitLQk/b41YDNXmudgOdVMD2IerwRTP1q2unfl77abyfAyTQdF
2DjRefg0WBC4PD/3vcYRklKUNkeRWgWA9qAb0WJ8WSlogkY60LGzZe6G1VQkSO3m
eisSG+J11A8MyKpV3coLnScA4eRGdvbtZMBQMaG2qy3/l0vDsADGdeL20ZfElc4w
pYv77UdVFLKPfKgJg1PKBdOdQqRsBszTsUJ7bdL4aBX2U3XPg2EG/ap894Y1Ty/X
t9J1fneebZPwcFg6l6nB+d2YIVUHTjh0MqyEGOmqzrxuSCaGXXnmvMIt5U0FqWQ2
TxBIvgWwkUY+lNmj9/ZTduSrtGkz4t0/CojuRtN5dPJtsv5STpRCWrbDXytj8Ttx
YgpPytPzDr34qvaZhyYVb8hCVTcWvlYc4osZO5jZaDXvsnclEG03RBJKvpArGNBX
HphFBoChGDePCwY8vxjiMSTHpNkpx1NSa3ghqbHzH6Dw63dRLcs3Q1/6tzZ0UUWO
I/CH0+y1rlOSchYOjkNHFHNOSPdAhx36ql20kCDznoE7AFn9l5qPZODkIpU2AwSW
QigJKQ0uWCmrSUOEdOCg5vgE8HRaUcUK6aQUHH0z+mpwpTDB931M7Tw6RVvY2SoW
VJ9c6AgzAO/e3Sa/AsEAJc220aRukhJ5lpW7jyUx5EBwuZAYPBY2wwzORMKMNAkF
FweVL7Z2ZrwsDmYtsF6wMGr/C5LU6ACManu1dgdv93zyps/QykvwtXIUCcZAfq2Y
CGRekzcWflH4lHmqjVStha1edr2Y8V51AzvwaQAyEUpxJ5j2y/Y5ys2Vtka0rlIR
Jv7EQf6lL36oFbtzHGo9GvpnKbJ2QhPL4WyP1FEdDboe+pw0hQi2me3p7HoM5rQV
9GYhKH09Z4ZMySkwW4hEy0rdbyNmefc2n1cWytCrj/Rr3iAgJ81hpYs7DPHyK2Hb
nRxNi/fRKGbaoGOYZtAvpa7KMXsBVtGPlzt4K24umD52Z+8RWw09etDrL4VktvKt
0rUM2s/XIKxL3egPUmDMo8VraaGkRJsBcGirVxid1XmHbEFzUHy7Uxk8MYqIA1fu
Qz9wyIWsN7iUxA8FkWLkHewg5Xuj/P52AOm7x6vthsp8dbfxWS+8ihFkCFffhQgF
quz450reqC1r4DygiWfN04MUClyYfQByWfqnTCxKlCRR4AElS5hmllHiS2WQVzpp
uJdgIhZrU/tkevk2/KejK3krqckdSySB02FzHG/iEr6sSSeTxH1JMlm8QciYW/yp
4ZfYrjTRYfy/anq2MrToCtZwyBxdPVFKqupWMIZfSobqKA66GvVpZxpVX4EDIZoF
M2jPn1Ol8AHkB1uC5iK6T4ymvpy7jSo1WzSAL1GoWyhu6c8yS86SoT1UjEVDXQz0
1QQ8/HTwTYcED/F50OLo/egw7oHKGKzsTSodqauXqMX6AU+Ou2ywWDSXOLtwkDsH
SlDim1Rb0VDWqutoJC5sbQCkdezFzzXNpNsqQEmTkerbi3JAiSpCcysRvfqCnagy
haco6SIxOJARQ6Bl8Izp4nUc7Q3z+CGer30VIezB3E8yhV5P5ncJj55ZM/FNVyzm
Kk/u2saClXg9au+rMZXuSH0YBC/Z7T/40++QI7A2rsEfa7+wK2yG279q2IXhjbyV
vDVItd6jh6NsYTfzpMR60z9SHwyaZii+g3XfhDDWUJRu58a44vLwzNzzWeulBpcM
wouVZhFyl+E8oPXGaiRkPbi5DAg+rYk/EraxHyVjZGWQxKNH1C033uaAx+UpZEdB
dAdpoPZnNtZWwmaG3zl9AJlspEpeQ1mQsG3/Xei3CV/JrHv5r3bJ7z1P+7faD/28
fRR/HnPiwbjR5KUhnpnoONCOM5NbdrMP1hUlHF2CEjDo86T9UZE7+pyKjVTpTlkM
F23CtUtZSY0nVKYs0dKnAh/z0/xQGWj8D339Z1Hkks9YEVEj5WohpBiQkUEK95a7
LbFzkuv8mo8xYrC+Ji3dRNtzYqK9ZttHf4vi8BOHoK714ALOfUrvMFM3z+ZzmE0K
9/i8ABucd6bnzqQtxF0ajeLjWG1F/Lr3xgUMLmxSDk4PZsGWiGkRvcXuVhmWuhjL
AU45+R3t1X1Y/bytH0akNVDFuhi+/ODByDObbE4JlyYkpBnDWVcF13k34DYXWTjR
gIiUavDPwA5btpuAIkKGExkrCjJLQnndT//v6Bg0g4nFXFLs7ADswC+32TUYfkzP
HGJnMGM3h9xUGEK/agTAbOJEbxgP3Gqv4uuKYjIrP7ES3QVkKNTG6QD7l2bdfqsR
6ksDxbMc+QNnxolzfWPCr61XoZPCvohCgLPYkEU/iVoxWMwVg2eA7NUNcH9r955+
OHIhVHQh1WOfM8jM/HIt0MNoNeDeZHUWB51gdp3iYnnoVPhFo+/GYKffXqYf85DW
b0P5It0h1Z56vCzs5oyhFN8pC1M+QucwL3hCELdoeH8t/ceniDUwHQtzNdi5UFeC
0LU/qayhN7RV1b0al9EPhEplA93C6UTjO2K54LaaTpauoje3XijfzMfncEgimxr/
Cfjls0kV9OPBZNQkoTyxba1W36DVTTAnwrWlKgnmzHeqHqnYvNt4t5V07RFcXRVe
bFfrrEIUU1wf9zibkRBrx8OOB/Srm78Zu+crnmSvXP4qlPDKI/Z42ur2xAiS0gG9
r+Go7Q2c0yrJbCbVIuOEtXa+BA0E94IoyxRDgwu4Fk9aMOC3+gH5KwUA9kV1ObmE
XxZi5fe1dgULZjEg6rcpl/aN2Ci1KABH+t4DQ2F4I+PDAt1N+B7KC8UzsY0TopHv
y7sqegfypRFQYHYyLqIs5lN4BmIiJeqH3N/1kncJBZd7I/k71Id8QSegaQaTCvPl
s0HIIO6NCPmikhhS+C3AwXWqtwWzy9oTa9WE2fRrdankJJTgSYqEhwdCvSxjnDOZ
ihDb9aG7IEph6OuCd5feNL2rKpg/q0ZQw9gp2j+g0q16Q27kbHVQmSH+hoypf0AJ
SE1oFW0OYAXE7Rt3FqSpNPwL74y8cvARLOtJL5CEmcbZwXiAsww2vLTBQyKQ2war
ddvqioZUnChIT445IDkLED1SB1+C7rZcXPxoHDP4aUqitB/mQvFqH+BcDhtXq2XR
uIBc3cPFvp3+TqRzPtO77cdCCmK2r8ttF60lllPwEL9v1aiIMDHjvlZm9oz5cMmC
KrxZPZUTQsc8uPY6OYF6EGIpMtuRPnedvWomqp5oJSS8FsA9oJT5zf/K6px8MuB8
IO8jkJ9ESSyUtkX5Yzz09kZo2dJ+tNikVrESIwn4/Xd81fioFvT8wScLvLepZKsI
eM83n7wWQ5MVD+Y3f4icTkaU/y5aXIWJs2wa2wtZfn4VjJ1Tcg5IwGoV3ttNxbEO
63UURmo/roSh7sphzHHgSBKvJOfWCdKoT4tfDaQwyzaULsLsEcMtREMdRzC37Ru4
KGT463FZNrFVIGdRp3TV353NzzTyEh4Vl7qU71EnTChUiI+tejhQZ++PfYRX5jnL
2x3jFYUJN3C9EZOHdVoP29UZBzN2u54mFBf0yqTflrW+NOHVl1VR4m1nDjMCO6i/
h3QC/3fkSzAvLv5hFVi4iVb8ylwe/seOsi3zeES+y9zPkDLnUWXTBityFqsF4XRG
5cuEMhdL8H68l0LBzXaYFoI50VcYoNPJMy+ap6ET5WVOAQjjQecs97ACWpJIJHFi
TAhkhisphHsWZXBw8o7CjGvEsHczA1oM1VTMmHpQShPnTTh6lflQRpprKrNlPE/n
dBXRmAXxQNTBE0/xjqSBYS3BsvsTWsk/g4FW3Dt9NBbb4ecCrggghacu6Yv6zSCW
6/9JtcZ9Kk3KzWqw8JB7cly2UxvNXlha8fvYRERP812SrDYy5aHSD6+chQXm7P6h
1KYDsyIudRqexrxZGc3HvWTgKwxxq8BUILtb8XIXqNkyaAQktapkuOua+Y5XMSTZ
25UVxXWeCZ2/q307UhOcgK0Q8c1w6aPlq97KUIIzFPs2IKqkcqjvzJnwzjA1vgB1
IKVgI1cjGW77Qkfwu2McV090seB91mnHNuYVfBpkk+mZTKUpC2yWW+teXJ3+W4nM
WQvaB3YkRiprC2cpLDQ97vhc2MZAvMVA3is/YxmJpdJsMollG8++aAoXcy23LbgV
Tuu35kR1m9rX1XMPQQispsflUkhqlceaBDRZephAbbsfE500Iv+9x5KlIDyIqoe3
OEr5CO31Wd+AFesPickU/w7xVNHkIMJYjVAdRo+uIDofH49hfxZNHUl/Xba1Co1p
k+V+q8rNzsEMTnpGOM/cybQhuxiDZr4LCrldDVVre7CtXDbM250E/tIIQPJz5Mj6
njx8iHNnlVgOgFUDCwztyWu8TczCjS2wwt4CQEFvBRlNt2FFnDYrPYpQ8zyCUX1C
xBaVE0bg4WITs8+YuPCN313R2ruPnlNu5mWZer11z/RcNzFLiRRA3oQT3+i8J1RX
0yLBtVB1ebDMXTCwZRhCw1tYrCJdenYZWh8PNXjSMBEQqe2KaMgcOXIqxBC8pCjE
MXs2YbaBywkek7W3yiRJelRgg85cGrIjodi2arzmGw0bqRmaGHIV+uxOYi/PuHgk
L6JBz9N9eZcTBAXkllb0ZaQvqUYs2Lw4Gmhyqq0Y2PJOplgvLgGd463B5oNkpXkI
VR0SnCuIAqsoqc9ZFzBMh6fgUscK2k09b67oqoeKniGUXNXtmKLMSBWRFCc0Zv7L
EBFShP4Pu3EBr9MNOczyUErQRVk9C/IeViwp5txy3ppCakZZOAmW9/Nl5Lhu4zjF
ckj0hhKLHUwhEMuRhDDcfrHHMKQuceAmHRy9mexyGGLTidLZI7EGr0OPR1907EL9
Ps/SJYqn+nXy6ZmwuvfI9pMfvjPtC5eubkGrTefWZVFU+6V5tVOGv8UKkcT0eTms
3BAlL9pNcgPC9l0HDI1/fxwaZQkySs4qsEqWokVAEPXMlRxOIDoUqeUYraVu/Ewx
Ot7Q81N7of9M5Z3k6yhwMM/FrP/xwlPq3252/6YbBXR/J2cyEOfp890/m2f6/ANG
gDQHArkBiXGx0ZVhfglJlT6te/wHsRzwXsBZbo9ypM+krHXchXlkbfQcozhSc1e/
AJ/8NKWsK8rNjrutJ6LqIZ9zWd9sLmB+kvr60PFyAPltsD1t0oTyyeSWaKTZuzD5
IdiEGIU6fyjzP0suQc5VqJdr/QYeEqjyD3kjFKSCoWgS34DwnYNllCeI/w2uOfTO
94c0kpRg9wrsHoewO7V0A18kk6wg04nDj5j0UTfCqAgBnSKF3xfseQPLwNg8kb4P
Y+q77mjEkPMoLq8ijGWiwcCeBCQgU6Sji0e2a6/EDVmrhBbleV6xEbyTj/d1EQfI
qUKWqlrhNoRhKP/IGYER3vlFLXKHcNcf2yJvTEdvsSAkt7Oc0nOKiEBRvtQWteBS
3vAjNA433xPmTF33+8gPQUpugIlrh4BkGyurOYTkWFhfN/tzeOynxFKpSboQjTuz
5TQT7XFeUnvPvwIntUnvpr7Qsfwnuqs3GM4xBOsk3FQoGAr1TM8BS1tFZLlEBwNA
8gdh8C/ebkKUMkx+RFHscFSKBa/HkZZCg9Lt93PmrqJbRbqZuHiDfKG560wt5fBe
sqSHbUdKZdtsxd9q5PuGQV9GGbz/T8yTl+QtfskDPUFuU/+YPSZI4yiqnbLRb3CB
AWGcAqb8IPpK6P9gZxALbddLZb03t7r8vivueoNxbJtyfAcYf+ds3ejeEULnOmrs
8hV8DYIwn8cYZHfaoxYut7ea7E03HpfRLNMK9IXu3BeQw3hD03xJ2MZ8ELeQsHJQ
1K+AJC4cvBDNKtxKSNqaQK5vZLlqRHkXDQTARoAtEm40unPIOeYfTQbSeZfnlzhz
ilef0JxaP9ioAp0aVG8yVI/QkWJzBXpVisamZW0zVhOMS0lOC7ImXdSkMnwE4Uj5
Tgz11+ERJlo0/IgO3kioHwGHAMkvQ8D7eZel3Eb/0TjEjGcqmFQmAiAdd3nH4bbP
siwLDqI5EWmMYsJCeqEd2ORsEDhluYhowY6FV46jL8qrActkJFoUyYxLcsxrBLyH
0HynpEt2xFSjS0AICcDUSy9rpo356UyH84J86OLJULAWs8J1XXZd5UBa0vggUUoO
gHP6F5SJFYBuzHqxq+nVzh9MqiPOifqD6npwskpH+BGUaj7w83hDOTY663MThbMD
DaqiLI3/pg2wdC4NUbvgyjtns9lwgYI5ErjKEZ+kOZVevM2WxF0Wx6ZH2eZUK8ry
07w3ytcUvrh8P7dtam7dknypFpZWVDrDJoMDv8jJsqDgSqv80coDRVh22LE5F/Hl
qyGGfE2JCv4MYsauQaKoRVF84yLcF7jOEXk8n/rFrCCFh0wIZ6gvltdm58S0Kg51
Cj90PR3WrnHe+qQc7jwii/W6tvEpWph46XxoMT6yn9uvmxmiL8N8bP2I0q43xgjc
xyqNVS3J1HWvU//YoE8HPB9vXol50eacTaa4F1q+mAT7dc4HWjRXTaq/qlUAw0QH
lNqqFx4AUdV7ythH6aixiwMS+vitAgMOH3uPAxSmFEC2+C2L3Tsn7ui/2CiXcXE2
ftSghjyiorMPOdT2iGw3+XaqeQLYVYUfamV0AMyCFmsMio4S9LfI2zodf7dVKFwt
ox04aPn9B61jwi1AWMnLZ/BPRL+XqqoNsLIEIVyNjUY0GCRC4ZAcLfkAtPwjJlI+
rLieTxbbR5C229jxUthzgEpZcd8+NhG8RJSQZnGWsswuZpaZRXyLh40mPfFM0Bqr
bJJM24F5IlKiABEvJ9PR+jdV7P3+npZZrKSYl4fRFbA66qYblch6qPAuj6Av1tbQ
dWnqnyYIpITpAKMvUcP5RWOpvdX8yRWy629Db0kiIn7PKLQ5RnN8Z4tmrHImo3ok
KkrAR/5kw52/1MOIVuZQqDf/SGu8xpUa6ALBi6dIaHKkMjy6IRtoU+7hKhUEekvI
zNtph31JWV6ou4PSNrIwbeSjGfkPSp/TtJ0E4y6fVTd8BroT60+uXpfC5K1LEDE9
nzmX+qLRRs3i1/hqyz+Ur1z2JLHUTUL/IfbaJG49jUdbGNaJ/q14mqJid9zFZpam
iqf08p8S2cd9WkFfblYecmtnt8eABjbcaTcu8/MSIFNT6q6UKAnnni2LDZ0PKZrj
n0NMnK392b7/yWMUyg5m9a8dt8J71ai72LAJ43s1k3ai01JqVDo4iBdASOr52/q6
48zVXfJ3K7FfbuLXF/uJ9jVIVkeMNRRmyfOFoQQTTpb23a3fXWzHyfpXLcKvjIw4
CpN26oYI0wuJoJKDwJQMIpgxxhRVnKj9aVEDMbkqx9id3S5NqSxFE5DwbpU7tMCL
62JPOgAAXkulssKb+Yf/JR7cbIU0VzqZaB4XcHuTG3eYNGQHzLe/tkWzOxg7sJ9T
H2Lgc1beaPO2ZMGV1cWeE1jDWRFxQrGnrEpcZo8A6CofoKPpiQ8nMhYu6vkAXKFM
7KrsDpThiUQexL7VF/7Q+uTfOswlh7o+30tK61l9XVbv7sOK5NjYstCA1ROIayL5
W/DohNmhvt78MdscfzYz6ZHmFZKO2btM397pzyXZ9BCCot/g3h0CgPvZF2NEcQ2e
96qm8Ps+X8rOIhzhkZnq+zOOswqOP1RskmBK1AzEuqUuaCciqZtR6l0POcC9kWkR
uPFr4JgK+JLcNlPrY1F/E82nhDJ0yugskc2pijmA9fUZj5sapy3SSkIILKIV4zK1
I7iBpRXBk0ka/zbrfPygN5ZWNzDgu4cOh6cSjjHXTV7SN2mwQlApL6D3t6RxB8UV
1yb42F2rMiH/pNQ8f0jwoHlMx5YP+aSlQ5VuJQwTR3ucULI0hXIIdgFIkT9Gj32j
H0eocoVfe6nOgtbxgUqmcAJ8wxuGWSUv9/DOJlUCBg1WVV5VrGpntqWYpdEgBRos
NO/GD3R78U3JMraMR2PQ7QEA0M64gJDjgIL0K7ZVXzPWZkmWBmCH7fdreG4SPdrB
skTyjLLiEWyRXGFJBEYcBfn3cs5fSTj3wxGkNBsZtWBiVLxT/kykcQrxRoFbRM4J
QGNIhCY7CtdndQzCDdO755xplMfk+w5fEQS774bTe4Y5e5E4a9JxuwhlO9Nz7PU4
1u3SZvgybDusIyYRREOF9jvQYNm/VNjBptSL2LtAi47eeXuMhb2WxRB11r+AOgss
vAZi3nrbTNYJQSGE+Kg4u0sCgqitszq7Ojl1NBsXwzqFqSSq9o5z5mA8T8jZflJa
HOh7S6dH1HcHUYKOaRoRCzMHqkLjM87SmAILwkfIAmmVi85hutRL6mZE2boMFBZq
JAY71IgWzlLCMSN9HyZrOpVrrMGCVhOKM/PG4zrT732ieKxxJXR+xjce/sRh7Rr5
e8Um5M0A6coqO+qvspFEK71mxAPwGqFKgA4OaiCQZq1CcJBdIgafYbjIoLvdqQsF
+0UFXPM9s/Kd7u7hwwA++c2GthN2sLvtVQJ3U6x6bREh3s712kvauidqDOKgRW2y
isEqRl6EmLEuXUr4jw4v5I41pJqnsNMve4v+gxjTHLQEogLm3MCAlGLlkIMV7IYS
XvY5eePnAjeqD/Y2Rj22+iIqf00keGZAVopqGNj7XXGLyyB6bsjoWLCHEMgyXaja
eoCcugt7XEQs3TgBe8qYQRXzqFodNB96E5umGTSVyAazs2fQ2iSP0+pNUfhwOhPa
YjKhGSefSR6ZBXJHR/Ql1Ax1AAKJCDaEIS6CeNSAp0KZK9+SbRf7FgFzcX0PwId/
HUExntLlNQIP94fI2hHy+UAiGgT9bxsuhm2ZT9Dia+hUEvV/vXCdFehBsqnuwqcQ
EuU6mH/WJxDKZQ94SpXgp+iBXPYzpJDHDVpKjMAW+UDY5cVqc0rgvN/z3z3a961e
6N3F8WY4kzKvye+OCd3ueRIkXLZw3v0fVmMkQxIgoCfSUnx378BdP3JanOgr8Sy5
1nSdh7gnBI5eOOQvupZSUK4LlILV1ZPn97W+L4DkVvhpWksfo1MdTw3v4OXOW4oW
wJNXBolCNxfxxtRX6nukW35c6f2okhEmHcG8uMvusFrF9dHNWDNid3Wc8YGaJ90z
oqjeuqgdCuo/4iZhUarpxBav3grMwRVi1YACl7ybWGShU4/1wQ9zRHgYUg4Dy6m2
ZyNhtfb+L5dv5q9U9eodVAd6ieCTK+Vutn3tzaeqcwTZpb7o5sigUvsa3nqqhXsk
4l6K0w82B3ReEgSQz5WKrx95bwdgcDmDRuWmF0rVL6h6jBAgsc0LO1cbW9sLGcnJ
yutExkXRRSE2M0iyUF4xfaahEMJ72cu1GVEZ4Ml1PEjBsANRpywIxY+618WzUVwY
GawC9mpOo1CO8WjsYAgs8tzJfomkN3IerqT1Fal2lcWGOurygAzPvs0paN0c1wGM
y3lht6uz+XQM3ISwCpo4zOyKc5Ss18wu3kpE+vIHXCGUK9CaUFXNkhWlPO1f1aES
pN20uCvqF93ZbpndLaRAu5OZOyY8pztv+LwL3tTJsyY5TzsyxYCT5J/uYxIrWnye
hB34GcjEw3znWNub8zZtV8YOikkHLH9iFwyHnIqItQJXc8erMl3G1cKhrnCfADcK
iL6GsI2nad6po2LBEG4Bm2fRhsKDue/ulM3RUOZuB5RZIW2RhyHbALRrUyMYBFlB
c5TAOsa2yHXVFPd8zN6qYS0eoX83rl+THG88cRGGvZEd5GrHvUJbIefbBvZYPkOi
k54Zn4i5RWwZCjJwDOj21pCd+GP07OyJD//61FmYur61JAFo7dhHAxpeAjzFxDBx
l3UZhSi1fOZ4oyoAc/PkNivuuVqBtPhiasI3zBL4o1DGCsbDHNraWmxTKYWfztJG
24AQeJ2APSm9qbYnlaJmxEwBsppMLmbmYA6rIeU8Je7r3329k5Ys6cYwgD5AWHFv
XGz+fLzwzfZs2zB/Ulvz22V2uvYg/1jCukWr+/O5xLXKGwpzbzzOenXr/fsJrbY2
YOFvRi+rJuZkHI3jNG0v4QjHM4Ujh4fJDoC//O8Offej2vWw/dfcPF4r/122PwOT
eX1TLDXLTbI+Oi0T7Ryp+qt52TmYjvR1oaS3t4yxLIPgqw/w6QLdwV9vCmGvoR6Z
NrMy6K9+m/JPCn+RJ3MIhgSsbL3Bgr7NFaVNxm23WT39hU7o9S70louqAvOcniYC
1bMgB8cPP4sV5Dut1chYUo/y9FFVXfGHXLm85bQdTh9FleXKBBnLz1vL1VJtej7p
fOniCSE8Cbstv5MTmhEkfwk4EVi5PzUehR4DcfCGft5Mk3GKqPMW3ZNoWbtmPCZm
yYvuUPJUjU/6WgWSrwBkPV8Ur5oKFeiAqypo5xMGaMD7pC0bwwJgfkabBgRFkUp/
ciBtTbuknSfStrZKHcC//q5sju9BKWyM/wN/rmPNvvmHGPvsPx/F/Va3idwkTLBn
Y2olIeVJAEn++0tvhyb9eIYlNaguzCOnH318YNsxN0nFtB1BVFOBFcXUaLXV9CYA
uLnSJDPEyzZi0Q0iwIGKo/x/1hwNb34ApsDn5D2rvYOT1QnTSenPC1wswpegDv6w
2yUPWff4lvU/TeDSjrBvAA+W8gU6bEAjA7Qit6UW8aVE+hPzkMotq4xbrw5flwVi
TYBiTvgleedCmyjo4a/5MztaBHXzecaSUmE2RO6PMCJDCkBIFEpQXXnP//4rVFZ8
kozVJQDMKT525WVWRR0PPPydAq5ktyLG7vTWPH3mno0TcI3F8Ovr1LpZKzureL0c
efqw/xIVbXz9/W2RslFFPs2pEwbmTwEs4tTVT5QUNUQZseLPGpLfbJ88Cuu2/QT1
78bTpCffsbOGOsAS+lxtM63I/HCJuGVPqYMD7z/yKB8LwidrcXS3yhAWbrv4siCg
xicz2LUvj5w3IPc65SatTbIHEsAlTwXaoOEReEyeh8EpRAb7YB96WUzokBqbL9VI
2+YMC+4hDc8hw1Y1aep5u0dMEyTrmBrIWPJn1j7vclDBIInr8GA9RIjkOzuGvGX1
UJdH3GDio/T1vUByJt/gtjx6xZxISF+dGOZM+8dzZTyvVrhTtPbYzfUpfEE4WlQY
IY3TDqLTFPMDDaMe9O30M9R21n/0khFOVFu0ovJM3t4kV+wcbyxvM+EYJb6anq0/
C2hFCmCPYzdjoOkSxA9oc79E16ACSjXOktxmfxXs7aFsk3zZM+K11EZGknsjYvhj
5ViajR6F+3YlCBUCCtjCZAuAAdjaJSX3zuxwtiUpiCzli7mStzmUtGTTzI8Rv6+V
bb+jDTmCiMRRjtVySe9vt/YIaTg+5tpx2Xilr2WWsa/EutbzixzfGfye/x4VdotN
ZfHbkkIeuiIHHY/X75vuwj8s5HgKAUCz/pM0/Sdg4/OAifi+aaMQ921LNfSsQfyX
3iXNyE6L+EyqQy2U92al92yfv1PCZwxB+59MNgDhfFUEQsapbhwX/yHelBHNvfNf
R4D6v2fabJrvlFVIUqZfShxjvVZ1B49SkH3ZtJg/cWInM3HBfNxjkz/XORHB2Fug
WLjWqcF+RlVeepHENDSjSa6BZB+Fj1HKA8PqDPbgS3yEWMVeniDSagf1Dd37BPm3
3sZYVCGJsXUuz3mhifzkpqWJe6s0sLn7GQyejsMX8BaHqj0DZuKaFLNN1ag4Sfs3
8Y/5ADFpTiKBHMKkDnBwOPEFY1poSS4mfmN4aUApDEuOErLYlOlpBL1I4GdKR+GQ
EaQFT0n/W7e67P1suOtRMs85IDfmWrZpeEJ/2RLMW5oa+kuWF671pCS1oP/zIJIu
zXmQcHRvViTa6dirCBU0Ppb1b7vSReAaw0xoMa4dpvp/Jtzcmv1xs9qiJPDpIRip
coS9F4Ojm/2rU7dfFldDoQcL12nXrGm+UTPmi5188Aosx0PqZ7aFjrOS544zUUo9
Z+nXF4DkVWsTQ8ddCFzLDblad9d9YB7EGiLH2EtLmNX0CAxT5kbyIsm9oWWeOXBO
tix8mxb3RAdB/uOkFaEutU0R0s+NNR5qr1G+epX14N7H/y/yYJhqcLrC1mWbBRUT
ZNST/e26UOjIfbAX9IrMS8SUJOYNUfPkDRlLs6hcapBQAREsX9yXA6PXJ591Heja
i6SCxtveNyfKHi6Ug5dcUkgtAnrWGSLN34f0hNKG9xcyGQvYYX+ZCFIzbvLJU+qI
ubY6rUOhdCeGGYF5ePsTyBWqa7e4ES0Khg3MDddE6qxRaY3A/Ul3qar8N4gU9Ses
JMInYW9NeK9gzhq6YlmNCpftawjz1UjHB5EBqsQspUHcBAK8nSQ9IIww73HdUrXG
krDyBj4Qk7YSMo2YFSsKagTsnEuhEbG1Zxe4t/B5g/dOGYlZ/ZPA/qieKAIPGesh
ULGuJ7AagWUznL26xDKYGw9ZwMuYyC/nAJ9YSte8MCNbsoF8zzisSY3WKOlCtleY
QLCzaXMznxGIw+BRS70/lOrcZqmsfRZv9ZUJVgBInUNvXXyJjtHNzGIS3Q8bmGjT
WEfGWhRdIddvQDwbNCxHpZ8bp6tmYFW3/c4doM9lQcJXrKQbmKrFliwltw/7fies
NvBh6+pQxhQldA0fj/xhWZq24LgpqJII0uyKA4vGpT+zmilwj7kuSMpEwbF2ahAo
wnaHypXHsgg93ZZUlg4PQcJRQGxnbmh/6Nelm3rokcM4HwIiJna3/+o/oSnACuxO
D2bReYU2pIkXTjS0R5XCqjSYJUJe/uhIAzpAhE+ilae9/tMJOQful0eoaABPUJk3
61lkwz47TcY+6hVb4/VqqCYjYn9ro8dAQ5UrOphEGi1j48rGsoVN/eUeNNd3LU1M
vJGhfZyPkmPs3ck3vxHjEkmEyAp+qcqd5T3D+x/Wv3/cQqOT7gSeMpM1DMUflzqU
azjJ2MiyRwBNtkmDpZdYL0485gQ1Lx+T0ey45aYvQptZUotjFqoT2thXrYqFIRFQ
Q8VceIrNDwHFUcDtEZqTHdfYGnWNLkIMjuwN3lJZTCWWyUujvhI21JEUq49WGoIe
umJfxXuvvrbkbriaxgfj6v33nAulgkOIycsdivzN/TjSEt/U5/MqIx4Yd3OhC1lV
zRwDDHO9icf4xxpGHicoZtHcWOmhmZaXai/vfa3j7B0kTdpxys+cdPTQs/QlbDew
E1Rz+ZPSg+XhdqNj/l1QVNg/PxbGfoHFXnwNCKkKNPf8wDTuwuxaiBLOGWaDCCkN
nzY624t8gy6XDx7jrMUPSXPKEWLRB2Xx6gpNCtvY+S0iXQUnPdBsMSarEPPWCOwn
f58vxfqVf5QPieTJYOaGmQVKNitR+KLWO/9fP/SC2b1ujei9wYR9lHDmuqUG9w+Q
LUhYegcWWlacgxgivWMRysxGH+CUUW6P0/Yg9Uyvf4nFvWXalHIBC9Y4wuFbwo2T
uiGrl6zWkiYYtufcZG8qtdX3Nhy3IP8MYxaisYvU9DtM6xCqbmlkcaQTm55LRyqg
cJHaarrdKGhNeMsX65YXAFaMQ/KlCWK5E1Ed4t9CEiP+X8+6W9FCJNu7FJ45m1X1
wDuF604v6vbZNgVAep39emFLUpHwI2AKj70JwAjUWq8bDZDffJC0ol+T05HAiaqM
cYCx03Z9ie2R/ONDAABxDpKhSrmVLpjX+p6BVdG9BE4FtOy1YbyP25jpaVAQTcxG
fnAlD3uk7xaymvBSdubpR6slr2xOvNDz3xt38OL8GIJG3vTWZcBOrMP4G1DoRYNS
4HvG8Ug9VdL/h3KDilGeFWDuHBegLYRyiYxRbtht9gcuJ/JGqLoUY+lWJeQKTrVy
WT+Zb+bvQjfITst0FDUG7LTQL6NYYFPf49cBXalKgB2CKZizgdVT/Dzap0SeUvmO
xQ9xQyI0pZvoylV746ZsmroscJn0AcuKO4Hs6mx3J9bytpYlRiQcChez0VsJRAAM
i1qZsvSNYgb7dznUK9Plm9zPbn6FJTkH7fAoQZCi2r2z9K63joC24gMzrEFKez9b
92NZpnx2MRzRJiEUKwn01RAWa+s8nEZairhfUKdtpmXiIzFevgX2Gj9FgqwyxQd6
vign8tSDNVvTVisH6QgUobqQmSIUrwh1HHdXSLNr9MSp3rjkHs+xWmUy2rRCayav
b/0fq5Ds3DrKANw6WbLnVD0E4MBJOHXOlXBtnxRPV/OPI3x6loPxX0Z6TU4Fy7g6
iVIJUyUeIg90KaaHuve7/Mp18u6y21+8Qp9fDxxUzJou1FK55cvrw8voSpjXdomv
FHzOw4yKiL3Y7w1eGdwfN41xXAUgpeuBXtdd2uSGQgWAii3nXWzbPm7c2D4XxIql
OjmSddAN/tievORCVUdWYWYBs9rkLJQ34x0Z3sUcGfcSlINIgtOrbQZYQ0taBdAN
5hSmrhMSgG7TqeIMo+wBSBtZpH3PSweLdPg3PNU0i50uRRYnPv6gvgkUGlA0NXGx
WpsH7boP69+UGUICTaBUb6b2QpVxGIjYOEvR3Xd1wXl7lEriAGHb+gMnQytyWuOj
fmNnbHu07wFkTbzimNw3o5Bl58cX9Kqrp5ZzzsaGWVP8kP9w+zuPEu/E4gjk8qae
wwpNTT4/i4B2YLudmEBjPmw91buAGLjHeC7HHc962MCgBuBxpe0QWIpZ/7Y9cAKS
qDiC6ncnsNgPGk5nPrZl3mX1ASKt0o0/Pz1IePfHaengferXKOOADbcdiW5n/EV7
eMr+F48IOgbcO3FZ1Zh9+xpqfZULhkXxSNraaYHwbziFURG+qCJlZ72F1jCtNv+Z
cpt/DvOXdh3zB7I7jFdxRh3mok+KtBWJ4Apik3/BTkE8p9Ng2I4lXYyWZtOZJcWV
WEFhT5fY7ium4NDvqewybzCfdqlcxlRfs+IDOSpsZv37KqgpgZ2ZfCA2h2w04Lv2
tyZT02V0BxXwjjVegOh4Lbg41o3Thrgk5XBS5clMIMiTgP3O6HPRMZIAbwSsNTmf
PofqO7sqSNbhafBNzTT6iTF1I6/XgS+vrFBf7z0dmHqIekrfRX0ctRGqLL8VQgwG
9mk+bjnFkW5KLGO92JHY/AY+LejSJdgKq3izwoB83KBRvucrsEXfRE7vQmXD3wuY
pIx3/wfKVWHOq3ne97PjfaaJsVTemwl8wJRvYfj+kiwKqjF9Wt4uF7e0tR3p1Znw
jMl0vcKuJjL8G4BSyFmHScPxWXy5VlSthatJo02+hMRXt+0DK7pnb/+WYO+UdFJ4
KJCb3bUfyJbTQTxtl+cX1ofQnGHDUkcVtLyhUfImBozKg6yGEDb55SZWiPwjoWyi
DYyMxeX902THUkP84Lbp5DxH6jErJz7YWiOtBtjmWPf4W4BdwMyBqcocNo7bC9va
60giOUHNapjvbVA3dULOk45bE7aOLbsE5RVwT51IEz/VR1H0hoQEROOPUWDxEGlz
/1/ua3uGyQD2OiIrZCSv4lkYXjMDT301L3UdK+kUNZn/+ddmcfZUU/R+r0gqput1
kWQAVmFkqIAQmvXM1t2ua6+lCkm+uhJmD4Ep99GRXx8QWRvgnyL/Me/FbuZb7EJ/
GZWSw/ESqQKo2Q/JwmEUgfahcfR7SGJL7uBkbMV/eDxZ/0o8kZxRIHlLUHlDeQeh
nYGfwL0TEX72ATNj7sk+rBpTLMY+WuoKwEFMgkORzuWNsJEBIE650bObO+iosWbl
zyQMzL+q7PiD71kG8nqdW1eMT8nhXCjncHyFlSVvDbscXgL2zQ46SDtA/h7krl5S
HDpYy59o8413/h11HFgVfQSzB9nWtuSpHnvIXKdMq5XlLF3T1n2NmPVFsHJdd6vt
uOx/C/7lqzML6Y8awTxSMgVQrJ1KLTUH29ersiNyjos8GFeJ4OG6pkNE0joGrdVu
AqwFFToPdw3bHd4AIs0AYie/JcjMN9KLfwk61pRdonMO6aRFLr/3Eu6AiPR62dRt
07CEQyd2M5tQ5cGFPNenqnFRUBiQWLPS9T1CW+BRWVsOKCFAW1eNHR1I1AawxIvt
ZNtAEOBE8gQ2OTXt5BXbg5aZp+RvRvek/Ou6O2h4gVWCxzZ8JuOkRBMv7zuojXWO
6WUp+G4xZy5YDnFaeB4muk5o8lh5Kq2QzmEGPPGYoJwMlADenbyvP54gEiGOY6bS
fpEeiXutE/NadsD8Chq1tOl87Nc6TYDY3hpsc/3t4+g3yIAT5wqsIxksVyMIzBrA
RDj32MfXxXjug4PC5iFnvmP4N2OuixnkdlenxPi/NzM7bAGu6LwjoVCfXYdRaOrh
B+r+FtdK7fGih7UxD77TjmTjHDhBX3kRhKobSAMVzNsqCBPDAAcVECEhPZdf4pCN
a+IriC740Rwir8yBtNXmY2UO1hSex1qdaa/PpelHqDvLH+YcQ3rnvoTAlN69kSlW
wAn9L1vFxm9n+jXGZwbjr/NK3DIZ2qMZCtdAx5YAhfZeZJ0LDl2VN32IN/wpmd28
4wVgr3tIQ8Z76DqfM4vJomppc9SS1frPhLX623Pgx2T3ehMnRx73c19q5ZERJ88l
NB7q5khmyqgSiEbMPYwlMfGMGtF36wL17VFsQf4qpZ65i01/Z5UY2yirJxvAZhR0
X0xfT1wBVio6UuxvnM97RJQ3Fy8dNEqTK3uPNIzbfcbqrTGCxkvX38Zn7silrIel
zMrMn1+7zgHzWnMGhY07ArQsYSmUVf6Yr1EXe5MzfN1K5Pvq6YATyynwHSONkuGl
0VKnJz+Vqkzh80X57hXNx5lXcu7dW/zE2jgz2kvLBhLWKTL4uhUc25ZHzoxA35dT
D2cqIalZgKyBw4aCb36pGQnE0CAsN6XLPWy8t7Dfn+wlUTX15Q1Ia3mgXJGY3csU
rwMa/y6PHtMRAsyPH434ASEQrVO37d8HKTSbvIDhnH70W1OrcYhUzwkj2pL0EZXI
mq1pZreipnd41JvgaV37unWn08+r0xfHMQ7+tz9qk5mHyGUFhE/NX0c9bRoSrXx8
EYkiXnia8opoMum6Mt1BsRr7WoD4JcNZO9+Vm7A2TELtD8qGBusGgakX1EeNxi64
k5N23f138NV8FqL5jqYwxV+wq/Ngge6hICkIXxUDFUgbQiOpATTeJSa4dcYk4QtB
JGME4nZzs0K2y6eGolaQg45SVx1t47BhThKwSyYd30KEPiUpwe4lpYIM5xwEzNNJ
S4WXKLOqx7+eXPDvY2dInAmOEJdxR9tRQB4RIjCEVQSfwWJbzdMqw/VLTp8kR1Pg
s6cmbsWDdCl/hgQwKmVDvxpxhznf0c+PqhM+KocNStQp9H9952joyy2d27r8BMHA
Xm7dfIgmkM0rzUH7Qz7f9l6jloQl2msB2Ib4Itr0IZSNdTlCfHzCoyIQNlwfTYia
DJCNmV8BkS2TAdUg0z1XC5gtxlQI8Y+0OC6J0ZbmXRFbNNjlGeNHR5CdeHOfwRnc
fIUg/Bqv1qsmoGrwMdH3bOvX+qhGHBWwIBbmQqpN6k3d1CMmo5mKe7rPRTHWrexb
KTwFLLAxnXCcchvSPtGqB0kIYD5382ujU+JaiqPdzNQLq1pXfHsE9R7iexFZ1SgZ
cYKEIejuETZbHeuYxsXQp2sU5l3eUsmzLTxWPmEVAJKOE02tJ0AX1Z6lF9pzZkzi
+sqGQV+n/7NeSPplATgvZ4t11/imeYC0s3F0+TC/p8FejNrKsQPYmiS+CW26Yygd
SW8C0H+D2AI/2QzwdwgDJQtPGHC+ewLPI5CfFc79P0ut6oTzYDdXS+ZLST1/5WTq
Cjv0V5GuVuU67Pb/oeakcHK2GO3MP+4IgKA8NXEO1AKJfg9zPwuhaSDeR8yCLEy/
Ew9xgxDmFgWZRJ3dq2kiUQYP0oQ5iIWE6KdV3dGZvme3+iCQiAlU++Bh0KL2adxN
uUsceoKO2ha9/bh/CcFswuZBT5J9plkMWGtzZijnQcvbstA6VH6s5Ru7Kflggk3u
ArdwO87GdAZw0hfxfymUC5HFhz1sJrqoLnwNsBKKP76fhoURrHaVY4Ymyk9T6QG+
9UPaJg1jV7BHILvRRYXzRnlH2Z/J0ZPcpzyFYuvJ+Cm8hfMBI7vMlsLH3EyLo9jA
VNa6Kejn3YKJfHZ6gJzylx4ERyxJh5CGTt3qK8Jm5j44nkkas5GpMo5N8wlAM79f
8D95R6rFUAUPBPxxeT9bdeQU8+lU5ltGqGweTH0bk6pfglhDQmpFPtBBPFvc/uN9
/vwOjnrORHU5xqDztGE122KG+epvdGmbe7MyrR57Vi7u5zkVQ/ir4wkvTqEXmvFD
jv59/xUc1+/WlXr35kKsSXEOoSWnbCIygHSckIhwxwYG+JqcIytGig57lH1BZkVR
2Th39iB8ujpO04GaDybXE9FCxYKW5T6onJ0pmSnNN0RtzEk3fa+S0b80P2FJ2Re8
J8UeOGr4tCQQ+Gze5fq4oOgtXr8760IDKnpYG4Ps65QrsQbPJGH8OrcSYNjOkPF3
1XHTK00NOQOp8zi0GOW8/86W+a/lvHUviuI0i3zDaa6aimtdB8E/TEgV2kqiXp+0
ujAJgwlAkAdVj1GJ0HREfCgeP2W4tyVqaVjGoVXzXEWfTNOYmT1hUUdth9Gch17r
AXyG2Cg8qc3U1MzCgA/DETy078INfLdOFz0VTzsvTna5afwJT1LF+5/CfmjOKLl0
PEOANiCC5OJa98Sik3Tgz+hC5aq0ch585NR8V6njx1GadLS2kINPgbkvTkcP+rBi
og5Mniu03N0hOlL2WDthB3VEwf2nv1YzQm9D5sTXp+p+PRSjOjor4GIaw778U179
udTrxn98SK34Q5++Yn34EkXuMHhAgV54QZeZKRoLr6N/HwH1ezGZU96aybjKzudL
68nT/N3m/7uMMDItR1byqb7+0JM3HqDBAbdnKpwVLj2OYCTAYuuA2K9G66B9llAF
00eE28F3fkMR3zR7fnbBUUSzWoE44MyV6lXnyi3rs3YycveldkTWyHDjyoVHXJp/
12H/JQWbP4DEExvaJDP9YibaT78x4WA9qCRYT/huPBcwhrJ/7I4RgGxof5qlK7Nu
tk/u65oEZtNM/e5ymDc7Irz2Z428dlOSinkeg5y3p5nvk4jpXdQqBDxCQ0AZxZrN
vGt/5Ui/LkiSMUfjWrqk3Ad34DDtEhu4VqZoVb8CUHr71CT8dU9aOeS7CP2XaQnW
drjdjRs2kx5+kXYHZDa18fRN/dCvX4iK0JWlT6Bo/LOWohrb5mqgiGmiA5piU2dO
v+577fMYDolsHZTV7HCNNFW6tVKquyFoS6BIkSHlx6ZGLoF2AMSwf7R1ngFX4Oww
Ll8v9ChAHCKRlDhgtAGURdpvIMtWofXUfcPr1kVI54Q1gqXf5QT85b23TLaPX+7p
DxGfxdf9Hrg3awjI5nKR0mw/0U9ZPZX2NAQTPrjYNiU0YEIL1yUWg2jiaFkHHI3J
0b/eMFNq4/fXE6t5r/KmlS3J86XmIH0b29idmHI5eCUltMalVCBTRw5kg5nRrV8S
1pobeFVgPIeEworJOXl/8V81tpg7hDze6hnnI9I4gjHMl0Su2D2TUDwd62HOClAS
cbjZRhNioKEsnjDMgljMSB1+SOd8HQQWsebfo9TwsaJsnxbb4ft556H9sJktZ+la
kTsHT6+0m2Y97V8nmZ2ZYJjjiQua5SpbyIqFeEeYXtdWEHZ+gPl4TpT8p6fQIiXc
ltuSqfj6vyAzzfmK4AZojCLKjoUx7VhdDjfCDmgJFy4kYEWqrqP71Ks3xmQtPfWa
Qs4wwZZT/0BaaDnSu6kXQzoK075D7+XtU7T7n5hULKG09IgO4+RCmf2apyfOSx9T
ADHF7/3M7jw9dLiSPJxnUcnXPJ/hP9dKvnYRHSzqGwbysBHzS1pB2VYNDXiANAWl
gO6vYG2/Rq8cKS+GPEC1JeLTgYmphOykcnBZQ+taJ/pl+eoBDryFfRLFeIQvDb9j
d0xuzfUbM0kFGfIPKHRJQl8rkR+Q8Z32Fh9Qql0/haoST34eu62JDKVei40NqcQs
ulL2+LBsU0owM2vUtXJC7JicOYWxXNTMZ0eXKqOSsaEK7+1iRxBF4uEMxHZdiYjD
cvj6Qc9hlmuveJlIwe4EApnl2s9Sw3SczRY++84iL8cXKSWCtR7B4Bd0rsgy40uH
QfbtsJL12lD9QzQElE8gIGT8c7L23nUgRLiEa0h6n2K5YMO1v6Mnu/okWYOb7+xc
cLbGALyFQTqw9PrFZ2V3f/aFmpzT136lfBivOVBbQ3hHqKG/Arbbk5B+1RUh/j/f
5E/kFMbQEXI7xshQfYxuiPDzwRnQKithmsa1Vwq8LsysPRfYwzvB561pt3Cy2c7H
lV2XT0JIh/lm4pJ4tJPc+PQLZGTFDDoY8WwJ9me5qcii8pqGLryBlV8RcQhpQvae
/FAdEn6z5xTiYlS/c58JjI0BdbTsMvy6F0zELlw5XKg9SHwHXPp4ioxN+rFVgtKP
NRYVX/BeSpX7PCmLl0kJaViaYHeIcg2JOuBZlgWL0XURPTOGClK1Q8kDIVhtAEc2
q0df82i8gOok00j7d40w25MSpRNOARH65dhIQcBiuUNdbGdvUToT9RbmQzaOIq2D
qJWGYvmj1JS9O2AClqeMimpnu0qoolxAh0u3eIP2Cu4tjL3kaMakknSdrnV3dID+
c5HEkOfz8CqVb2uN2h9poAC0n3jnX2+xzHK39SXc0Wv1rNPNVoI8vGHYwHmBgBX8
2TpXd4A+xlYYB1z6Yv29NuIxKy58eXDW1y2bl3R/abvVaaAScohm4mk1NvTHw02b
EX1OxrJfpw2fxSGLIIYCU1QFWygWJTfKASpAwB5GQLJWc1aSkV82GX7WpXsFzDuI
CpUWu0BGInK3flfxi0KmY1wai7LZrz1Po2f2p9V5k92HKGH0gI16Mc+OHiWjr/bJ
kFYQDXMOUbC1D7MyAnlvwqiG/v1AufUTBQv0sS/jEzK8gU3LG24kH8La4PUGxZR5
shbJkkoivx0YyrOADYF2bHu3qv5tNdQ0M6EDuH1/igryFP1RN8TUxw2YKnLSUp7n
bOmE1k40TlEY0qxpgtq+SoXrIXCS8zedR54BO1ySRNsVLIKjLBe+5EIHpf6WJwYF
PQ/kQEa14DIeXGimg7FNiBDDyu4L6NtkQ7mVKOQkPIVRk4zqWk+LL8BYeQW4ahHs
iu6pZVqBGikuKQZtOZjJ7Elo68qNPwZ+w5jiPBYWFDiBwTn2Cmrp/GRANyIAGFfO
MgU5L49UrWD7/U7G1c2ewWxde0IFd5pbwzfBPC5q90rHdnRcMZO+pNUswWYqM0EL
1xa/Cm21Q0ONS7C0ZmK/XZ5zEPt2+nZEKI5S3fpVpNyuQrgXISZavjOhvFy2f/zs
JgtBO+Kp8msHPiYqZAXUNTMdherRNFumW6OLMiB/7J0BO6RaCRu7C67m/k1kbyED
IiWr7i9ju1K18p+yBAqffd6xsiZxPC1x1lGi8ql/TFwbE85IQ3+5BYz7y/O+AAJN
AjCwS6AWR2HInUgdB0a80CIqbrO1q7+TlJUhdQA3Z24dSjwOKC0gQavDHJO1djd+
qBnWmlYgsMPApZx02ppFM7iJFMxbMvZPfYg/KzD+FmmqEg0XotPHgU0M2RklkNyS
9dcFoJmgcZb3jD+Bn+ov1FYAcMHicabpYVh8FvlUs+urQD2HQ0+Yfo03dEiyWLIZ
e1kSsai6PpaDYR5HRJplhCTqGP9tLF1bJpsT5z0O2UOPtq/7WIficUHpEp/0JG7b
Q/qAsUs9iEix+VgzIVDUTvfkBVFXt058tWMNI7dpO4rDF9mViGV2EOrfs0L77X7b
F2eBZzVobpNP5dLscpFqYbEQgCkx6glMM/VIsXhG3w1XRxzl63ZaWxg2BR/nc9Bg
St1CNFt8wym6MKsa++MTFmWXg+bba+Np6JPSPH8D6hxF5BbcbAOzv1VXPrRdJJ8r
WYJV0GKI9gpToYyX3srEs7yqB1EYHww76d55XRUGHIPhyZm3NmI4qbRQ4UHfrcGC
xOKyWhed3wkB7qitGB284z3xfKEfV1jDbvl0f3KGRf1cdy+TpUIjmNy5tevTcxhn
U4szc61egsGIlmL82SznxvJPPMgbgT/XcgujuezGhXZzy2Ts+69+ChWiTUByWkAL
xklVY34Au/LXwn+addOJMj0IMSNbgvDYZc1Plik5aZ30GUHlXpNfWqtOBoGvYJ9h
OsV9ykVIrTL7yH7F6qqRBg94sHFqm/HIlhYTxtr/ZSR2YwyTpKIbbQf37IlP1sIk
OMPJUnhtXFMd8Uk5d869mZhuPUASUdb7U6YHm56p5rby+g8Sppvdmjnna5ba6Dcf
DGF03kGF3jWLE9M4wIdvVmI51b7N8gABgduP0SHrx3np5jQ3C/z39rzyJpEC5MBn
3qn3a3aq3UjybDMHqkWCSTDdqjCc1guIadx4ubVpDqRsSADy0z6Q2HIGwk2YSW7S
fF5BL2yo7ahFW6ecowbKkRq/gDkc4FurE36mIAVQCo26j5Pe1uvkXx2A/LkK3UJK
2WNWacIEB2/tPt6hcKf/xu3v2RSeheNi3RaZ9icki3PLnWLu64g548mjTF4IIAPu
bngfIFEg4aBWg2m69ypuf232jkAzQEBaN4oyIZJOVjzMfR03FbSolBrUfJf1QKRH
z0eAcP4gc8AGq2A6msz2Oqghf4piA/ELqGiylSGozq1/GMaHj+ix/DQ0Bb7cf77v
iFTS66Vh0i1XXb5ATlHbRhVv8+VWzWK70cCkwYmh7+QM5YUUz03UlEc/Ek55OumV
zHeGPcjmE5MU3KSTKm8Qrmx313F6E+7g00yzRguX3NugsGl9bBbsdPOOaibWXrT+
Vtje79mKStbrZSUeE2bYyZcJMQKvq6XM/L07J1t+LLkR30gz89QR/sZvGVCpLjm1
EiGgUmSfeqGyfdzwfsSHOlkIX6s9IJqD7gbHU73ZTI0eBJSe5fkQJvrj5oL68MDr
XlAW5RYkzbZqKf7qx+IO6/aqIrNXMOD6bduogrtZM9xt2zTjyuDV/BFyPkEgp3TU
eJCncdP5JHcYPqSFJofHt9BdRAc+HBqTaSHOcaZ323lHMLY1CsZRjfSk/XtBUA68
T+6y9x2+OTRTdpL2Fh1b2PsSTvdVPnkt9BY0NB8/psjV3cUtt1yBjQLCUQaHI6bR
u7trBcfzcaSOSVLQgU3Br6VPFAFmiMHJosHho+Hw81AHO+hFxKkCZII/4eAbbaVZ
oAu2PgKyuTfDxDmKPtQg70ehCrM18loBeoCYiIh4LC5ozfJWOMVawOJVbsp5NAn1
ymQstNcf/DlrdBZJKZ2yQ0mZPhzQoRCCKePYlsvUjxO2Hi8txucQjwwy66wht9ss
tOcrKuz9eTSqxSbPL91qNfUhjjV/S2Lh3g1z2gt5GMpROcKiyZxIkyaWaL7MD8vb
P1Jtt1U7rfvY7OavFI7IJy0uQJGtYxWMHkgyJMXeRFsEjmNDnaLkeFTay3Ge9YMV
6Z94gKMpw6aQO6caAt/7IenU5G7MD4Cwjjt5D54xz1F6tQ5nT78hrW+ckxQaTCtc
iqxs2NPnBs6+ka28izlB20Pf3hwt7odId57mHu7JyxWtYl8ghx8g2Omi/Eq5zcLg
jHuyXFiQ1ESoiB1AjP7Ezywl7krjaC3PD/JEmoWRcIkkxb8YE9cUWj5tehW5ksiw
1wZmDA3cevHfoqFXQDZKVPvsSfcyViadW+g7n6lb9U83EuCI2szxlZMzy+VBMNtP
FeRy1TA5KqINP84kSEmF2FgniGQhByXSWMgVxh5wUMom53FhI+WpDEdvwtat1wWD
qhYp0ws4bo2kBlH3skljz/HmYlIwtMEqKYoenp6SaO+iyltrrtGA9R7HwhQLvurg
69hF3OBw1oantezoiAcZg35eN9q8BR/0n2yUxgEO+1DdG0WXMZ5gSMV16kGFqSV0
IeWWGn6x+UMTFpFNKTTCIo3dKHaJel/siqLtiEzu+SWni5hWK8cOYJet9W5C3wHs
bKJi6rXwwQ9Oy/KbcoSHxrkUP3HgaT6SSMwKz+TK0rz+6VDQPmWRNQEGuw3f3NqE
JZ1HHPo4x7shW/dJasnT0d9EgigsR6bnc6CbSlKZ8qHpDiH+hs+3d9QeAC/MR5Bf
0J4fR/MAkny25Kqvj8gbMJFY1+1jA/q3cE4mt3UtDfF5al2/LQKmq1LHWzNycPid
FLfj/QX+WtCaL/qpqRcerabFe57Q3sTCiG08G5jDPzkixBToBctjoycpo4AmD/at
8iwqUCwnqq1PW9uXkyreh54hdT8EAbT4ZNxkI69IUPXwPyfrXCUVsQXHRd6mP63R
AjoWPXuNxosKG+ED9DlTS3GNny/t24Od5mDCYj+ggiSMtg+3YvMIrdvTFxGqTjHZ
v0LADVMIUrAiVY3DniT/s6TZ9v+O9HjAkWQBDcx+YS0y2DOkbgNFnr2liGgVtgg4
fp/nKvuCvBUkHJ7o9ufaoD0xK7/azjitcp6qK+TyPdlwKhFquIMZAmrImiLUujwP
8P51XfTjbimw4L48WnPE5LeZ9iaXzOBvUpyZHKf4FMnbvkDXvfNQvqRKJbIx1xkb
96lsGvLhZZGGTXYVpDqZ830Usw9ik7W7W+maABu7QQYqme7VaKiITXJ7kUI0DXi/
SaZQySWkA0WurCE7ukSStxm1DYQ1p/+HIfjmVcK0iiQKkhG/ND0/bxGzRRD4FAWH
RhyvgpgJrIvt+9PPeXHsJwtCp2mXY3CmX+omrJJfVWr0fUP7K6YEPCId/fq1l6o4
DwiHq8d1gRyoo5old6caoFBpSHRrRjb/MUCHzhbUcLF7TAXKb4DVlp2lGMwsT5Tj
grsv372rpG4uenw6XuNr4q7+A8ZxMvy03NKkTMLJr1dwvaFFcQU9qnNQeMPNjRCU
cOJMV4//PAKbogUEdGG2V0t9p82FGv98TEm5XKUFIkdcTU7H8S6cr6MVvVZx8ofb
oK1m1kUbMYRkk8n2+IWOLe0JP0Pdk7hxlBm4TFWZUj3GpY8PKUvwc4fSXVbytrxB
4v5yMd5CgFg1A/TyaqlDGkCnliJ5aG/psDqhpTGG/jT9hl+s2VsEqnnS9IqODDjK
quplkPFbBhYzAUg3xh6t0YgsqBepvWZlzAFhENIs3qWu/hg4d2anu9S6EE0DSor2
0mr8duSWHnJOYqSzkzYRsQH9vYfkIj6EKKohX9M25BdO9keogLQrba3A7492ABWw
ilwsgOkFNiAlUvSerGFCKJr1v8JRRqCvVbkfKphb64C4G7to4nvIib38K+arXh8Z
lYISxbOPcihEhU9WBXkaPNlQLbo12XCfFxW8SyxZdXW1eyJMxOkIvPt6Z8D/FRak
w3oxruVHG2jC2zIv1e6cDsiu3vCAE/S+lvc7dtakgROlMLZDNaifi3IIdhvf7p45
m9RcG1HCk9oO89is3U/T8I47rvLqrWc0Ly+USFro/ETpYDH1+kEbUADIItclh8Ir
mDj5VL/WsK87SPthTDUdzL1ffFeREIOqqGIA/1lRbZVrea4uPW0oTqe7L7amIjNe
iTJmfM2kBenhDKdd1oPD4vHCzCgesGK5ggv/eQlPdAPPeMKA1q8FWYIDZA+7rdfJ
tUUfT5L+UuIiYU90ryWS0Ugpp2cqVIGQkFIEYaCDlzuwZ6AmP97kcpJU6cvw7hCt
qMTI4/PSQllzWq1RmBDDDwmYksjyQgWyonyKvexRaNz6wuxO45JEjMGy/kUgVPP8
BFY0nk6fjQJqebEI/XwZbYXQx4H2HRA84MSY6RuE2xDv5iGSNFRO472DN88swtUF
hQNC8f/m4Eq0bGQ+FIm10SLVJhpWkI2wzy12W5Gzv6CT1VJJUvojicoLLy8B8OTj
odcoXMFX6zMYhNKAsKI+wY42rROkDhEsahTIuBbFw9hSV6DrJde+s9Sm0hDOHxHe
wtoU5oyutrasVIdtQM5G57ZrEQyE5Y/8ihcjN4d2L9RHe1ir6MX6xQGAQG9WygM5
ZuMtb/aFVQnZmAniJYxF+/ZUIXC/4xy7mJJgmZRTnZ2EspVZnhPuWZoLcc9OxQDe
o9S8vFDp+cj8KR2BjnH336akKZP20eDJirMNGbJBmqiqVEuKRKQmOCDfs6osZccK
88yG+14j8xB/vPce+T7WzkukDyVBCqhfIX0+B/9htLYWw1kja/jZQzHtFC/UHzYK
BgNlWvS2vSg2WLveNb+bjRk0B8u1CXS+OuHk5Ki0NVvndC9fqkk0QfM+OPTlwD18
XNPqw7vb+2s/yA/d7m2Jc9g0o+npFXqR7bnzsJFzGgmuZ48Prf2CMQSMG3uZjm0n
ijlg1f3mgiIFPyZYwFW3HxO3mUYqGbb+yTFDH4oDvmKMXQW1W+zSzGCrwNk8MBjB
XBCgUzIKsIvRdwqTZo1QlrQaffRicPz6MzbrVmeKed/Vwf6+jy1mncVv3021MSx+
VhrhEarZWOd7y03Wn3gaWMynEuSk1rSqI1mauWC1cGRrME0VwRSoTktws/BjvWfq
cmaxTFAOSBc/FfVKWF8J4mDeUQNGQNk9n6K5PaPSzfXG31XNjN8KMezzFblwyYkz
YZ2LnMNFtxyEEkeWXYdGc/4wy+yOhG3ZCmOboGYZuDtReR+b6WozwQU5xUfk6paW
RvzFQVsXW3V/haQ9xAjNGDPceblV5Nm49tMa1+MeK9xXlKM3odjzzYownxjPRLJu
xn6c/QMXfgVb638QK7IdHbTFxltDZV3r/xOg+Ln5CEceVBYpZ2RjSdswdURbyBkd
2d1UqMy7pJ4weg6n+aAwMuBQYhh81oDyO4M2xbE0QULqY7Fm/0GERgvDtLwg1tuW
8Ojv4WTwjMIM1kACVa039AP8GuCBiU9aAkE+c7HcPiKU15hGyNjeay9eivGTDdlZ
lVoInuk0vUcJmUhbJwYVh3cbKJLSn5WUQmzV5wgCB46QMRZs+zV/MHs/jlSEwHvZ
iJrfNbx8BoYcS+KL4mqp/fTK+ezmnE70ZPNqcqA3+mQX4F26XhyfIm85towKmZl2
gKgFcsBtNO+kxWghrciigxgujwEKD//EGnA7WhRoOH1E9MjkG5ULkknqLsXwqzGO
Y125RVYlpge06S6WMivfhUwXKY4jYYLfxJHoToySrMRtovG5NK157SzXE5/ZqhRm
52E4Ze6motJ3xtLvdgdbktZZE/8jA0mghx7FPatuu2nj+iou1DOReBpK3KGGHsHg
IMpnyCAWlKjCIYSMACawOWrRvKHkaVHd1vj2wIAy5zC5MaNcd5zvWHqqlXjCdM1C
t2ejRLvE2xlSxsvQk6r2/wEmTxpSgIfUDDoigf3N7CA4Q/6gAXkl7VoDYpu133b6
j67IGZT8ZgIptb15+YzokUeCdxGXM2/BGzPvJYvqOs7oXzx1dPHzFszElYDFqRSk
tl2JHuAth2QBpRDbD3hOkIkne16uWvvdzPTHlYzHUWUqEc/yKzqGjVaODmrbwHfI
WabdjQuIex9WI8pGZxl3AwjEhwfJ9z4Gfcz1rI5FGsAYJhy8hYIVuZ0ZRgmTVWaz
/rKsnlur8uDZSmZhbSqC8TIP+kwHOH59mUo9wGtf5pQCS4uEe60KZbBkv2x3JJ8r
2ctqjQ+rv1pujUXJBF0wu9sOoTmtLRTJfbcR3p0Nth3xPfuh70VPRZoqkImi68hE
ScIR95K0s+Ao2CRWUzb18j7CoMEPIH/L6y1fnSp8gyB/XR2I//qVHvnY/yQxqHfX
G1WOgMnfBpdMXK+KzgzjFF4avmuj+DYfkYkBJj8knG38My7VSpI0tXqtxSpf9KCB
M6aPJykE0zXxwIqgjZYzLBvLAnhvbhybDeltOoekdAka4+mTaSX9LA040c+zvhB/
0QUS5g1vfLEcbK/5KGp2fq7+K+vrPEnEI1HtJxs9aaihKxmQdwOdgrUYxZbYQCTk
PiGV/lzgVcgONQ8oXgQn6NlR40RT0A6pJ4Wo2oRjSP5brr9tmQKEcZU5W7VJ4Cyi
U/id7c2B63RCeWpnFhghJa3GaIYmcqexDorO0YS2jg2y6aCiIX9r+xripYuzmHI6
64j2ttilhq9TpsRNegbiq9E4+7Ct0YtFs3PLX3O+KJn++2ZSnSz46EXcuDDxH1S7
aLHgFfVRd/nnIEbZCMRcWRkcqZ4+0inpm3AYU5Se3ENmZ2rNZFWd7bPjjc0llADW
cXQHJ5vPRRKowKm9Wu261km5DCEVw2lBwkPo4amuPqtGJhDEG586qsFb7y2aHsHH
PlYOS+khmNxL/7L6xXsUi45/wzLPt2d8XdL1dni4niq61omPuN7waBLTno/tqCUx
lro/2GWXaY3panBuY0x1og2GJr+jXZFAQyiS5cjn6kMFucECfBbEGbkZzWTHkOy3
98gt2OS4Q6vSFhB1T9Hh+/WPZBHIAzzZQ+HnIaO3L0pJOvZkD4GMH+sWroszLpdy
mBO3z2k+ZDe0Qu4N2ZNTN97LUPi6zRl2AfuiPrXmjq/1ief6yA28jgMrHNePTAdr
+4bBHg/YlHEJskWg9o2+BhQUwk4yZgE2CDig4kxIEdd2KQf0ZnOJawNzeBGSnExJ
4zB1Azckagqx66kl0Mdz78TR1C8xRyuU9899eilpFNtf+mbiXTaxkZD4dBIlpRYD
elZoqPcTLyT12I39+6Cxb2s6sDD19F3LHyOosCIEP3eIdt71T9C9ALMp5K/Oy/9v
XsqntLl2WBcoue2+tzc+mx9PeMVt+U6DZvnKr3HqUK/aQVZXTkuZRuGWmfz7CWnE
yWgk5bkvqpqqhNQo6wkz8Ml4u5dr79+NyDkF7nbho48DMRPaz1fYvGgPiABnEVYK
Qkayy4rA8JFEMHVjXPvZgU7YFRQUavFqsdYMYXG/5+57US4ZCkDnAnuYRhSB26gH
E/6YaeMjpeFu7bweivRJ5PID917hEAjE6OFXp/lR+453UH00Sz+0t0VBENLbDGjZ
NdFVROR66HsrHIPV80BYRqa2kcihfEM9APkdGHN69HmkddHeJYItibKzs87wZp2R
IvMc2huxpdAsBxnQKtYCBEPLMksdc2NQpPKyPGh6QbL2JV+fv2JG/H+nGGeYv9Jn
BZrKxhrrnU/xZGuB+bMddc+vNdW2gLMK/D4gIILTOEWI/miZVSCIcBKMjd60HWDl
FDzjtF96IKDk3D1hoaN8QIH9PbnHzk55eiJz5RXlYROvsG5NVreSXA/ZZpe4HwoB
pLfmHptGVG2jvOippZB5s6aXch1LRhU5PtaWn5K/rVyZJXzxAR2JDMMwgQbr7Kuv
/jclmVNEtIE10U72mqeKKqrwf4rZa0XBLy8YoCnuiP/n2gGNOnfc3K70Emh6p8HK
6ykULMFtxxm3muHPBuByz0C9D5AKVQtn5t8bhkCVjPbpwGC2QD003YPpwahpdHw0
Hkxd0om/Hs0tVAnukRONmuoXwy1cNUg3YnDLcmwzt3s1GGcJZnUmeCRGBhd8m5Io
LxIEGTTHDI5GyNrzQ8hXs+BcZlcQbFLlB51uSm08EZbQBdWfc7YETSjZ/ebHJ2ww
DIvXqm3PN9ix7thKvIt7/FM1jhmYbASXgd0rngFLFeVlZmpxtWqj1/Il6oCOFBxA
RGQPMrCJa9l6uJIk84ndXdYssFKAAII2utXCGt0Wqj5jPRfdKGQnxVleWeFYNGgn
+WgZqZg0NZAn3owqwOUClS8kyOFfyz3qVaYFG78Ehw/N/V7lu/WfhqDbz5McSjUJ
ZPHS4oyu8cEQtE5/ZXV99Ehrso8xiqy1a9mnrfaFHNP3OglEilEZKL8K9s3cW+fg
uywc6TIdPBNFi8mpmueBHhszgD3XzfEFIfEBPUeKqj7LxKAVDXN1GESryzpKdviW
m9DBbXs/mYVQCG0ea+yE4oqlSad24lTuxZIXpar5NU2nlQcMN4+xNCEukKKtISMO
npQarfGk04g2y9/Wqe8Mbzf45f+EL0/+cdL9/OE1NcQH5tu719Q5wL+AWWTpIAL7
216n1pkznA/P344WKabikgWIpEycCrtkhMwi8ZwIJ7+WtEtI1IwFleW1kbQa5moc
fpwC8HaY2EiNIqY6DMxoVZqlf3f7enR1z7bRxmlH0Eno3wbwSXLQlwf9hmKIl59N
IBZMWnxdIMYgcJuN1S4c2vWMbZm6QbG/XWZ2wRc1XAzh19w2GPOeHYNMqT4bCSat
uCTacfAMaNOCBxxm+Qffhz/boABhO/Vq06MhSC/lbkz45YSHZx7BWIUEwzF+8QoI
JqPbiUTdyDUcaLYAcBJ27uIlVL+O4pZcKn2oDjDdJHtmZW1wQrdeIX/pDPOhIlt5
Bmwdh4WdbDFOx10myP34YUgn7eFQ7f5IfhUD4srVHwe5ju5TJbR62zPj8j/hyYu6
6VAFcniItTJQLCu0OST+2h32gVJ8YIihKA+lvDtcqrfD+np25n1DoQ07VjiP14Yr
xVMJIN3Zh7ZyAaODZ+n9pATi0xY6rHLznhRdfl4HlXubBu4yS6M3E3NmXHfmKPNx
5Tb5liccFrgi7PEOdJcg0z0rOP3VsJodkLHWkyYtglv7ykAGZD07ZwOXW/QxKtte
Jwztbljgdi31BXa3eYk7+S22f9Ku+hJo1GRSMSBVq6cq33Aw+wNfw1OTuL63HmWk
LKT+LdhuQfcZmHL+v/eX+HTn27ZSBiDdWLRuAAZIgS8zfY1J8hU+HmLP1uRy1pej
OHLUk6dIWigli4fDcUAx6G6fn7UqKsRxKBXo4+l/M5XxIqDkJitByPSE6pOBLZzB
RYajhsAUz3psy5f3Pj9r2j/rm2VZipiDP4QQiEy4hZXLqr0HIZRqpAor7skzbs7f
8gJvmeH94pdumE6cdX8SwForzci4oJZXt5Bcjq/8L5d1EDySYoFgQBax3NmmUzsb
ulQwM81sXUjTEVnKJ7tN7np8DLg6mMOHV4yGumAvCQkw93wHxdTtE6hZaXCynl5R
nQ+dhNgCWq3AxH0HcrZ9mk1t75X47PIMx1qe4iLTFin/52bXkCFMQe6NAdNQ8n72
JNCjXaS18ISdDqrm+7VGkzVxFLNrqaEUT5XY7BtJCVS9MHk7uHtwYgVtFOygxdkh
21ORJXzocoFqy6lIgMy05QzYABAiaINbxEB1Tmm31YI11wRb+jp5bCBT/Zzw+NJR
K/oogvJbpPmBSYqN/U/r28yH2m7s0yCYRh9cVehAJdBq4TKzjVogFeYExPOg0qLG
1QUbBIC/XA19isSlb1oIJQV1u0FgclXrFLxkVi0njMPnmN0hL1aO4oJ2JknLV6hM
b9ANDakNC+a5VuLGF000gCvKEdDRcG75UXwVOslP+03u8b+i5aqkCO/ZBltXUGaU
jKxYs1ClT4oC/I8S6uGtfC1tzvBIYrPOxes2knwJ5cAssMJHVaLgg9aD3G1BH32t
mlddyJ1CwXk6KY/kGcf9jGYqTZCP8v+sUvwRV4acEeva2+nSAZ4Gxqq7LYt5aW38
2X1PnE+6GlSXausIMYExGbkpF4LdKbTHxo4xgo0fZ+ck6t8CZtAPPG2hmpxcoTUl
33Cqrv0OjOWvdOtett2lFCGhwoMMbCb7lAtAoecIep9dSBwQlem+9yKrw6oRTcMo
MpU6yX7v68Kxolz/R+0k1EEB0A+pVc2Ax8h/LQaU1O0CLFGCVgnNs30a/KlL3O8l
JumlL5IsbSGIAXUxYB24TyT2W3ldsV7eoZUxaFPMIOnorVNsqoeWwm7/N/1zppCk
wuqpbnC8+17b4AL28ZtKDzx+i1UMZN61Oxn5gt5TYh1i9KsHaAp+WTALMzzUXdc1
yfwRI7cXToS2xXnD+dPTUi6U7bOa5dEI44ljTIyRdjsX2hixOuuG0KUNMtdn5Kyk
hcRhGqtj+hF+knx5ALtg91AsWSgchrj2D9ycvnp9TX+Y16Qiuo1TMfWEPjLhr0wZ
SdRudaMkcsUx7PbhBEp8HAUn30y9ND/ogfw8AXKK7KCFMt8T7VMPys6sbP9/VRgl
1RVrBVxmgCWeERsniYwmkFsJNkJIOvyGhejhS1cQz804pCvjad6bro0nUzVtDmcZ
MjjlNtOGOO6vu3fzqRZd6GjmDHr4EICUFOFtXLDxY284ue+Z0qyETzRHFj3Ojbei
1/+Dop4ldq1tZ7Ct2AO0pxJ/mnRVXivs8J26dzsKFUQg3ztRCmq8hYTNZH8TeWir
bI5ivocC23HpxsZP4sCzZWCRzDVLm/RkrNpjBqixqoUtQL70g56a+ooFLsyPgMJD
+rEmjoBCCLdoUi4Fx+0ZlStcRl+FMMHocm1MsHJGVI6+kVIf0YbuPOhvefFDCTUK
f0XKBRZAxf2INpQ1pZYg2za/rXEWKhZX4bsV5k/+kHn+gOhsJWiFMxuA0mSe0EXJ
ziuzZY+28VXaxlTBQGUriyfPt2xXn0tPVkal6DUFk8tslazk2Txyy9kmHG25sKI+
5+RaOVjIFUmgXv61g3Ap4OK395K0ftLzq30e94HsyvPUt+JtiF+ziYFnkLHU8swj
rP7TFrgmHJso2K6odWICtyQjWcaY5ouSc8/5wvkEmP0LEdzqI4jyzcIMt6hgVQTZ
n0HVxy+l+65Bv+W8NU2d1oHb2u2+gx3tGqqh18JUvqOrxmgbvMR2ijhKDZ+O82G8
G7ZdkLyemX9nzGE/pEi5TF7I51mzs+1lJRT4FkoK28daM4/84wLSGSyz1qqG6IjH
WWZ4vqPuVPbvDqV9csWtpepOHlEp8JtrpKK039IxWj5z14zDIQyvSumq3JKRWa93
sd3TqXiLJGE62fWWutrMDhv1SwLd7lo0o3fMQV5sN1pHEebdw8LtALVB/3z+k4sl
2WDKrKD/qsVyQarZt6DwNetydM8pQSSfaokiNYXbp9p9VbzgWgoJSXVTombHrXfY
Si2/iEpj6lafP/TRO0QkdvIBy3KSDJ7in0XflTeJAvke23liKammgQDKGLkI5/n/
HiPI7ydrNqCa3aAkYyJVBmfQs/fG0jZMuDotJiJVxbd4XqIzKYeWsShBFWAYzKfx
evEksCqkSv9/4c/d13j2K//u1hQQMKNlGvJxWBuedPmZw73/TP2yYyxwsaksiv4P
zxu020rv8iU+oD0qOkKY5vSsh6rDFXQi7uY4pFvcXJJqGL5d2Hb7jm5X57sg+4y3
AaG8X73MIcn+w7EO0q3dbuE3IFRTltqaOxQ++JSSKDHd+xMonXw2B6d85yGin1OQ
1pX8/AsZP2sTWOaZEy8Z1DP2qnDmxc+ro47qY3p76iUxH35CG8Pxq0z0jKLmuSHr
D57KvMLAbNnRnNrXf2fwEMm2+CO8iwoPbs4vQ7Q8GS3ahdz1NC7lI7CdJp9m1NFK
/tbXa+f3poNg//Uy/mi9JQB8RY5cSv76BeL9Ij9978i3mA+roRRZMu+Fdf/OKy6u
F/tNrL8O/wyWw0UowZsUCQqhxuGonrUdF1qbbaSPosXKEmO4+Wgg5lQrlMgdKgAI
AuxjDOMOvCdOkS+rMIk7GzD2B5OC47J7IsGiYtmOAmMBWq7mtsR7HI4zCWAJqm4w
P+zNQOqPzxVTQDn2gj6d0n31ei7pg9GmwgEntiy2WeMttNyOgLhrTehBaieZaeV0
PHgV8O+PuLhZAJtD7N8k7LXQtXeTi+aE3o2TAgAJS8LshSepsOIhDLhmsvDktn9y
AAD5hU5kicZgnc4wqbEcDZODjJT0uUgTidwKG4l48IAadt2grXA55WzrZsmnODV2
RPxAckqe+SYgALAADUE0FNwZVKCC++Rnjzrtp3EsnpXfCKBySVDiQMvL7DCH1XoH
3dpu5aj5ya4Hp6MyynHVM6d48a+0K7lcYjiTfKF5geeedecvBF+LOpeVytTIsEKI
ls3kyjCESfwOZa6hGutOAN4T0XBLr8B1dWhA61SPHyQI9WV0azbjWCUI6MU7iMBF
sHcNq+9PGKqKEaNBPdEgHBarzH0FkyxXL3E+IuOveLxMToX+pZMF+wmTV94p3e37
G5m9qneWyYYc0mmWkIAy92NzjtPgKTFXPyyS70g5hrSwZ248wM4DwjPGgdTx5DjM
4J7A2DWEt2JUYTIinehFtdAVBZqHuyNtlLIPnmUUUa1DtaZipnJgnQuepThkYOtm
peahC5/JZAYaEhfqiwMBD45v+RGa4vt/QKRZuYfjVwkAkejxC5cDfGK4A9+3BDWX
sSTOdvDJpCbSw0WSdunrvtvC40NaH9LsVWZxyDr4Y8kHQO0FZhfaK9c5PcJUNWqn
+sCHVep2NHt4hps/phouT66OQ6MTacu9IKb58oQ8w56WEhjf1fVf3AsZooLNXOuM
RUk/m7p/bDC7ul9djYOER+iPW8Dk/XzluK+2eEN0r9NIw9o5MKmyR4Ihu/H6cnnG
4NErCAwJI4w5GwfC7LKXDeSfrRWmJdZYbaNPFNMp8BZ7smO8kbTjraWdLplC2hbr
Oxtq3qYHhkTMYeWb8if24/9FF27ijfR0LyoM+Wolkxe1Mq2HUg5jldMBRF7szP+b
ZPFDkJpBDVLKP8XoU1DqEWx4Q91SnxetHQ6TUiL2Kldy51WyY1VSk7DWewTF0cEu
CywhvsNVPkEVMVAP/BoVoywp18gEt8GXiCXnopnifo3SmW4xMLQnFXKc84piT9tX
ARpU7gBRsSgZJ+VNlwct+edB3nFjeAzy2OD/zjZeEgz7CROobnPBoaw7bPAdANTF
y+Hvl157jmjUIAMilgNH1mEVPwySAs3jWzsCn2D34scZLPnHWz0d874/lHFQigg8
HnnXWENqP3MzY+HYCwvh8Vy6NCQCdP4EV6iLVaBHlzM/Se6By35nQVpxE/+PKfN/
p43j9s5150uKp6NftGrL1E/KUVXEFsengDEz18UPSLzqsGrttngb4v63w/HQFm6X
4zby/0+0ZxBj+NLNgpSu9JhtZ7k+nDiFRw3rI9OtoKBbeXjHvQskZ8FBAYc2rGp4
KZbAFWrE3FvXmcFYC8IHyYCbFCLiWVxZCATNSUlXENZpi5bsKNNAdGoktedxuO8M
z6wkMHJsM+KCgytEMGCULiE+s10R13nTBN4PWyJwO+M/cAze4ODAtiiWym33f2Rz
jXjLvK/d8l/AFRtBqgzaOPWRPxLCtYdJo5+BsfX4pnJRFEo8C2OyLNs7IFFu32kC
A6qe70SXC/dYCDPvtYF3vx+5nQy5ycl0+qJDmyaQoQ8MqF0YzS7jwPyD86gO8n3b
EUJLt3ZbG9x6YZUKYpm/O+Cz5e0s/vZOvQaSXjrfVD7qxlmbdWb9LvpO4OsGs+f6
WhF+grGW2a6wmQMdeHiP7Cu6YDySRx+NF7eT6NM0YePZNZ1n7KbXVY2mVUQQLTNe
Im3ORBFlgjhAYiwxfMGfGaFp45WIZaEkW25GhwufaodDT8z3Hff+hYQMXL1dUmqV
W3GPcn22YgU1Knf/kmeQ7L2GlKs9RNjC7v2si/pAZ1JoE7futeB9K2OIelUzrQTl
VxX6xiotDMtFS80PBwc5TjA/ax0loflvd+MZOsNKMcHnG3WeD49hawPmXyzSS5DG
KE21XShRK/JcwgaDvSuiR0fRbHELsiSewVqZDnwtUTH4/6u4AYnBAOE2JuUDdVlj
Cc1mez51VO9BnqXwdav4S9MZop1FXog2NoOxUENiDNpnSI8MEbRfK8EcLhQ23pYF
lqNsoxq8X8N7od5mlEHA3xeA8LgiGIrYX4LyqAcRIKeNZsHkF2Pa+uupl9QzIW3m
EdaoSVCT3UT3nUsr4adewCFaLAs/tG3FWaVNbTdjXLPCuoB+pYTh9/LxZMUY6o9u
yBD6flkNT2L2eSDW5zh0QSpftIY/2xAhjOf+NfsHUhJNZjOpS01JVfyXT1TuJt+T
4AtI0z/BqFVaQqipUFTo1JZtSCnzMpyLdILtS/uj0unY815Kbqd4AeMWzmaHs48k
PiolSuTtmzFWUuadU/RH/DVQFNtwesaZIaShW5tZf96Lt2m4fpUCj/d3xCmk8En6
P1DN68MPrH9Mbmo+VtnYGPmNCWHpAhRLiCdFsh0V+iAJq7K5r1iloDsR+y2wIX8f
aGrlbNfcVGOj7cfhYnV4huOndUqhl0NpXMmD1VBChl2YsivLC3/zD2oISIlRvmEH
ncG/FQxIotLKkTFCZvLdGjqrdyYGmsuNSm9cLAT551RMBazSHXUEyBXbRT7yN5Ew
Jo4J4X2yds9J15Wl3vOkyoDUWiFMltYl38boLd6iYtWqvwzhqUL6p1z8N0Gx9JBU
gq2/ftrVb3jr7EZlLio0WBBZ6MvrPsw3gCPm17FZhSanPgfmWz+OC5qSQpRZcp2l
igrhZUcS03Gv4Af8ggY335RFLh5lXTVVMfSyFD0S4YXaQCxrxXaTdM0fsHtgHB/X
3zctOgy+YHp3sy42lcRnIDMwyof+kLffzNg5LUpdMc6H4+0KF9xZL6lQFW7QT43v
EBnPyHhZAjQpChM0EBWAieX5LkB8/7m2LGBA8s0CbqUbeiFdrbIJhUkCvHzOpaP9
qnKwh1+GXqdF7hA/kULleHjEN5J1k/rnGR6uxMRLRoyqeNIOA0A4FhLuDxsYLyzo
Bu1Qsp+pdQ0VAa8o8TbRETNRT9LaqNnswD7BLnrEyXgDJM7DSInd3XR291qJjB5e
curFuzTnyUwszFFJhcNxgKZXPxyny01R9licJhvRGtUMmlfe9PC6wPBtAz2VzhUw
1Nm9rj5EsW0yVTSf84a43+34IgOzM2Z1ngB424phoD1OOVte65UxpmWUufuu+l5j
GMmHf9tUEgQVi2aWgagdv04okmk9mKI5fch9sTKF9+NOitftyN5b7jLHzZDjNn3Y
2ZhIuNAnv7kUXJWIQjsX9o2PYhF5CjT3CAt1kUXpXTCGBUUNLN4WRfBBw86auyZ8
E1WsB23BANquEdaKRsv61bTfHF3QnhFwBOIZsukECTpzp5zx9GLr3kndHuHhTZtI
AudGRszwW4muKOcx+CW8ENUITNCI/54yTwkBv33Qj3zS4WZxDUAgEPbSrAT5PtPb
GET15hbD/WdTENtT0JPH9If9HquzbCWWiSk8RkKoPot9DBcMK2HVpUJ6u4wd1cXk
WWumRQQEIdS52RFz1XMcVNgHrTlz5H7UWplPLa6zQ5FXD8t1BgprsdA988/SSutV
YUKh5B3CNquFG9qHZrbhwuwvyrF0sccd4m6S79IlvEUUORmQVLGvWdCOslhz5B3v
pVZsWUij0+coB7NjUS2fEaar9+zhIVbQamHkGNCZId6v07DcJNWqeYK3XnjEe9Qy
NHEJpJqPTnhc72g95g4nsgTAf1PCdimF+15Fj02G6aV4rUotHq71R30g6ype3eg1
93LQQyS+sOKam6Mn79t0uGVhBrLv7gV3o3z8ZbUdlfoet5bdIYBV1E1sJwYZbtiv
KoIsWN8HEEry845j06K/HzILT1zku/qaQahIaWkNcKUZCQN9UMHTQf7TJKi0g2bP
3Zv+my2yFCF6NXYMqwa9XNUarlNdaRbasBd83mmxxL6XG4Ygyb/sgG8lM6I0HB/z
FEBOayhOeXO5BOWEvSS0a+KoEcakeyAhRQjGq0YZzy/y/qA5j2XkDZ8iC9pQk124
nPctlZrm1WGTcae0B+Ag3LDq8ZkiamcKns0p4WLKnN/kzZojzNJip+oSk50iZf/j
KzJ9UafsyvFyKUEij/3QaBRl34kOFIHFHgBZGTK3RD52frLDHo8SY9JaRMPqXXGz
ZcRHZaX6CshRlnZAZpZYIldiE6j65bK+RcvBPIwxEv7jaGCGJ55Kz4T6B3En4IiW
/5m8v8zsQdbYOvP8baEChiEidJjeu2YAAinrJo7ZLxLbBB63xPw3p+0iy/aPZVu5
6RuNb4Uj4HUJlVR/1k0ZTelZYcNU8nRkSmbzzqCvoYBKJ2M79uCk41za/wkeScsk
N3wpow73aV3dv2WETPzY1Nr98ws9x6s9OYkD40ljCxEbmhRUu0N4vvTlEP5HfPFj
Yx7RsLPOlIvcFO1z0bNZepMSJbRDAHVLV6sQGGzc8TLSCcY1DN1gi8WknAX71Kf9
oNfxbsrAk8swHYnnPEBdiJ3YlXWIdtFQ3Z+QjuZU+iBrhECHorvN6zh+fR+rC6KB
7+T3Z5NPzGgvUPYn9dLL78e2URQm9AQC1HHkaO2Vm9Q0TakhrHSThRCQWUcvBJTI
nOTrbqAPpzR6KBNPaSctqYIhZ6PQL/dPZA1+Ru7KVC/Y2g+xVpzw9lCaqWvbg9bx
N7Nx1bRRPa6ZD2hgA6q3uvSR/PvgmN5EGaycHFboWc1DdJBMOevfwGhUlcx8iE+J
8QZdaao0RALKef1iMQF1Hp4nA2AsAJjLYLRfxwo9W9v0wrYmEDAFtmK+anW1fO1f
FZ1+Xkglr9gNKRtGL9lH7iP8vqx148CszMroKAyNeTdDcrs8gBby7pBM9VJVt7qu
zRQskiGOOcu8WhFvHnHDBkfF1vkSDk8ro8T2Ckwt18XIOZoZBeJ/t+TilYONcbss
B8XmBYfbM8IA69hLeFJk3x/MZxLqC1QvdIBVFn3TDV/AHF1wm2iV0rUpruFqqrcz
pQlZWNcARy6dFIhqLatseGfX3oWKS2RxnOqN1Nh8F9zL0zZ6m5ZhlyUIukiWG1Qm
Ilr4MhI4owCZL+sFsXHm9WOy8xdxZlXSy93GFRmJOU6hJzz3uJQzpTPAz6aSxLF0
RDrAaX0xJC23v8HVAhWwyyA42QbEeK4g/B5s/drnHga8YoyiKNkse1VE1sJLR7kV
ExHdA/l2uUszKtG3/XzMr/iyCVaEBEa+xITjF+zkGRvDW6R68Olg42KlQ7M932qv
Ozw1tugqldFKLPwa+//Zp6t2uiegAavh8LmPLCS5wsH0Fo04eyEms9DO27WRfMwZ
LfqNzgE4sBWNbo32ieT0DDUI0dRFFIaoiAS0ZrnRbZWak1wT1nerknhga4FOENxT
G1L59X1bln0KMQlZhb36f0bQFCoKNE92Q4fC+1WgGvBzwUI9g03OpXmjbHIFPjdN
RWCFsslmNd755wCe1G+o9V+W4A8QgCM74J+GXRvlkXNJ4o6t6h9deRJKlq+RPmRt
F2xAschN2Jgcb/kYexKGWsRs8UxrdCwcqdaqq7W4B8SFJzE45LAK9/zBoY98Ddae
FRFGVf06Tho5MCe522slA0DXM5pcvs4UUFlLh3i6LQKnM9h2xVUAE/Idk8NLVfc2
FjRPX+0HjDQm8v5vDb9RCy8Qo4jIZz2/C9YbIs3QEdKQKqnxJm61yBzfysEeEPc2
xvwd53czwb4LLRzA8JwGYZYaLjt30FWsn6BmUVQ+OHCURx9fAgcBeXxNTp+QPO9M
cc9aUop/+6L1yXigAsGMnWeoI1LRsYDEpUNP9YP7Bytr8IJEFFk2+xr730RTrjhX
C1jVP8gCDts2v3pLngFiwUx9g+wnO1wFHaYIssOTJSTPXWc1X+FdWpYtowVjT0al
rIrvI3D38md/mIUhvvYBJEDy/jj8dz4Is8kmI36nY7XbTNKlTt14oJWVgfFRNBMz
tAjO7FmgE31iiryS0rPULJXHmnxcVagTTbNwtJVJTga85xPOb8WUig5kNWaM2tqK
G9mu9Sx7UNY8PqJe6pEVOD6JAM2mteE8DTBVBDnmxQ7C/KiLERdMOV4nr6jUTEKg
Y0lk+jOOcv4jq6YGXLCsM5EJMthGOXn8bDTUs3R6lUytXghyLhQ6u/Jas4k66jgZ
bcBqTFiWjOPD8J0BYy2e6WBZPP/SlPOrvJUNlmch5z/4ulSXP96W0VlVZGjy09b+
M9TgtuHV7KmbdXSZ8p9/tvE7H0bZrV4+Rfjj2fdEFyR6zmA2i0YoP/W/mV7IG3Ea
QYaVB5+8FpspYi/hIbTi/up7gxP214IxPAR7jEBLL8tTOuuSYu4WBLw1jwHt+0Zz
UfHJuhvrp77C0/iIv5URtsZnETqnBrOAxZ4720JXnmGqC3/5uCMRtF/VZIX/aWF5
2/tss87AH0qjpWGfxoScjDd5l/jwyjMEQLPRbEha7PR6I0dCSUDIIPXj88VHG7y6
OgcKzleCfaewJJF6irrRpsjvrUsjxt8QoboN+FAwjYbx+CmmgWYPXOS+gaNdfZfa
DR11J6F3kBQ2Ts5fznqxcjn8CqkLmDiyIIVo9JzMfWhhi1qX4bH1XxTHMQVZCybs
vdjPt8SHoSYddzl5yNr+v5Gg7bOkxT2CJ5Htkdeql1Jq4moguPoBJyP09y6MhtRe
F3OrJLnc/R1Koj80gjYTKow58x2pnSxcS8fWfLsSl9YpjWtXrhrjuafu07YX+rDc
legRjUHw8Z3NpV66raTsFLGcoTX1BF5fc14MNYhVFsimMQzhtChEU6BcuQo7IH76
jYe9Ulk5KBgG0bKW6SXOLn4Czu3tC5bDNsqd8w6n5vHYicHPkMdWQxxwGqzsIcXG
wtmtrTl/sCSn+ogte2fyd8XcY/4kBKy1a/QsKqiWv4gSYhLAyEiz4ypiQiavWK5X
uK7vn/FKmTfIZ6EuWi/4iPezyS4bVxcgFccQzVHbw80lppoKWyglUNOQSdStkq7z
txsJNssUw0prvTz6dQxukB7Bf74nWva3FsnP8Muczwsj697aW0QQW1QjRlQzjaW/
BHETSnCyhnP4k6CXx2LUyQ6G1gGDjE7Fp84xbtdQ/YeX/H/43NUcNQTR39DmogL4
GH1kQqzy9F2+A/jU6rSrcBUJX7DJvi47RYvlUPoaGufOwA49kchhCRe6ZIG6pC1J
5G2IDaF/6p03oOvf2A/NTMuXqovDnCzhYQcjD2069b0xQwDQKgXYDvj4U8zwAxMw
MS8sEkQ5Oagjaek/aMzmL1i324BitG/2oGHAaib/25JioLb1kCE+LnFlToh6Fegh
+E/CWqbkfqN4yD0eNaAi8DKZ4iKAvp6DQCIyWBFjHKnQvxqoFRageBlRXPoH7Ipp
pJrYlEynncXPS99dQifGMZroGKe8bLDQxCMpnwuVGLbMiQTrRthNqVYjlf4uGh76
hQNjuQPRaNCBBr8nXS22MoVKTGP0Xu0Gye89i2JIxFJh2lkvtA96K1cEYhmR079g
ODa85cOAoZhYzNAuVsLnciy0yWWJFniYYlXUbQJup8fzh0kLGdM6mKYlXUC+cuGo
Sj03DMYbVIZLYJL9jLxEOyIzFMGEI8uDtCc6vgf1QFbn1a1eYDMz3qY7tu+L+2xT
2WDcbVuYDkHrqISn9tSBOvz9M5p75ZGnZALhHEmVXPPmKlFyCsS1FITOGnI2uN+j
fJ0S2YRasaSfWC/fKChrNT5PxZWsDAxj24WhT/bJqBPUvvtMlr6AjZKPRXuaspIU
zeub3HBGq8Uv94toelmIm86Q9eXawR9WsJyo3xqXU5foeOa27v/360IvlwOxby+m
9Wtb4DoUnQwiwzJze4Zuh0cULFVyLmcI0T8/ldg/p81bJlX4Q4gIq6gwkzIDlWGS
wC0S+dvWI+j5k8USqg4YwUELUfA+STvbJhqcT+AdX1MmM3VNmGCxTKzZxpSHBQej
sJ/Foq+yR5p6HO8o+T88miyXvKCPCNYesD2oQ4TsSXqR3o6Qq50341zw+M61vzI2
BacXXKDABO3K3ythuLgqPrVAYDc3641RhpD8LiO0bjX1zFYwCojW7Szk9XaRr05a
wvjtKhsqrgMGvdppOHd+qehXMHaoSl2EpIEeYk7UkSn/8bPkjYU/6NtiZtyuU/6F
pyXak0eY8feJVnmtUs7JVlClDr1xhamXPN+Sv5Ka2Wov+4lvL1Zerovsy7rif9Au
B6a8XhP79DS7A2pAOOnQlsoFu0o0BSg73TDbBLEFlLOs9qIjcyQsK1oj54zcKolx
IsotnPDBq6z0+C1vpPmJjyaCaQ1QdUzVd1f1x8AEefZjzRqtBTe5n9i5C1LFa502
lw8TekzpwmIUBp7Ya+LPIHshJGL7hhMnjmI89eWHpiF14N7SwxqloMkeDGdNK092
0fIt6QE9LXMgydJm+7s4CNS9biaXAJ3PUQvvfvRGsGeuLvszhrnKqfYRHRa5qRHO
6kuLzXbT32cCzASdZYoqfzJuNaPVsw9z3mwd4OwjjjPImtJ6HnnXT5VnFQMXU70x
AL/asybl4pHgy32twnjLVFJpVOVL064flb4CigN5+Mk9iJcpsRkJNAXCyy1TZJjk
ALSM5smtXUDuTPJWFi4UMjHY7TjCimGbRPL6f4U4034SUE9FXy0+Z0U5UFXOpSIZ
Rs9FAWIvQG52EjnQHrUkOfGlob+uu0DgEQ6ECZy5dYCsY1mfEeLbEYAQxmF0sREe
8a1xJTN9eg8Q8PLzasVG/EcdNfmaw8OwjmG6UZIzZwsRu8xqm2QvtVoaI+YEfEut
Dkn7QmKihF83yfnhGYtGoj3b2t8lQGdIPoWQHksxHzKVjYC0Q4fMz4/6zKvEkgLg
2RNp+KDFmoa+5oe6Ohzr4S3hCiSDTeSIYYauQlP30+ohAv9TAqVOmOdwjFbmXg+X
QLTKFeaXsf7gf57bDqGb9gqTN0Rmah/IAQptAZ+MreXlbOmCEMLmpo5/HkGdbgSg
2RS9JQmYnilTJcIuWI8XufEM5G3id/1L62SEwEglA4FuBRH7aP8VOUfVT1AdymFI
z1/2csOSTDESCuS0d7srFjqfH45MyYEKrn63FJFllBeul4yOJBYGGx8h409xzxgQ
SPkLZabdySqng9AXA2B5ZLUljsNyrblqwefkbtiJnUM6fjPY1RQFBFhgFEqbHorL
xt0eGnTlKO7AXs0T++av9W4KOGEYrHBpp97IRR/aveD9/TxKENXmGS+6YHpUZnAf
nQgvJB7tejR2YR4DZ5MvD6iPwDvxAfInu2NnW9FOxD4B5hdE2PBc8YdQ//fDLths
2PHcT1/jZKq9cdszNR7E/IDje+9mgf2YOurcxQPMnEscjx646z/ngarzJXdLALyv
iG2vVg9Mgz8j4mQa+FluumiMbTZW5lslZr8z3FRsC0ZJB+w5nGncaDJXUioFRtwB
hqiHhxcvVqSS8jntiookLPlVCyUxNqPtrhQsR+p7ErUr5FLmtAHI5afrYtixe6hO
wGGR3tj/JRP0IBCOQVVMlonFhys/qBwk8EAEhVnXXWg4LYlWgiAkFw688jKwgTPG
m7ZFgSlesmpe4GZnEo7Sm5Yu4wY8ReQmM6s7Cy+6A7T2YQ22H7iNpB8He1lB357K
1cXTkrMHWVMDrKdmkHrDB40jTvEAuXXnJ85FctCJB/CotlSE8xMaw+yE2jcpla4c
2TPu39trvx7IOBNOMyHzop1y+cJ3HXiMddaEK18S/bND3CekR/qma5nv7w25IWkF
MvC1yYXLijaKnxqoRDQmLCrXdrhsJJum5ZIsK6LFqo9dsaTk3UHha3r2j35x03Vk
eROjZVUA/a6UdpW5lZWxa0IVMFwjLwVUYE38ejGaEpeaKENHINaKFi9jRWKWbCCJ
NCIxS0i1wvUm7X3lDYQBuUUSuA7VQg2ThyrzUmeRQdplvTMld0Ety/urfaSR1xKz
UveZaGSw8HuG5nW+j4o5KxvfZrK9rGXylui3jjnPL0PQJamw4BB2bbKup2GJGp+3
a1A5ZyAAoXCF5mAEoTN0WpCEmW8SahuZr3ZzwIxMrNmhTpmIlAgui+C5bAKrWm62
Rz4aM0nbVjl+VEGa4N0RbElOwtQQDfA4Nad8RWwtqnVa3SZxgAA77kRS9HOyED4l
iNeyLh7xAgfpqHPlgBsPMUNcnA7N7EIsl+3f4f59DKzgu+AbhA1Ha1ECBYk6sV/I
VB/lyOTh/bEMu7YAWhD5njuY3+Ua00lm2EAbhdeHJp38IWT8BAOnOmwMqmUh0ORZ
5u28+z613Fhjgbj4juC6zX/TVE6gSCPw3nZfeDergXUppNbHUob27ooYDMeGse2Z
2ChqE2l7pxN7HnD5WGUuzf2xOQiPsFrNxSRkJnRybVHlLj5duPfQ4XLhy6/xXB84
CnRzpu6Zkglh5cIuUP63Qhlp2++6IYszmvJzPyF+V0Lnkkbt5FjWsk1fcBsrJgHC
EmZcdpMQkfvD6RTzfThSmMfq+7ZDY+NvVVXNaSt8ek2C2N4Xw9znS8mlSIVdx9Ny
z/WsWQY5HhOhKVFkWiuEXxy+qlG7wmz0GhVFhcz1jyieaELj3yuRQgGktbjACyZn
1O1mV3qN99hMUs2BrXjMQ9xZwKkkDn/Uc+ffAD8Crq90EK/JEX7wyelk5763skBz
fHQcXhaCdzPtRaU7hxMEDCFxl930PL4F8rt1y+ZKqc6jBljShwNavG/qVKuX3K4X
lgtQ+ep9jOukdG/Ub+zIvnPYgPMwDjXmakM2EfUBm4c+8Vh/yJJ0tvyelBlS6El7
aec+XhmKueq20AAgETwA0WIbfgJ2/tbwSK1viznrlnbbt2AEojd7YZpAzb4zluqw
GQnJTKqGpXitdDTFOPkjQK09TQ1JEd5bf2mrRWnOvkfzQw35cxivgMgoIP8TwZaR
U9xxC10zwtwnVZKyMnRoUdbsiwn+7j7q3/YSw+an7+dZNrknFaUlhC3+gJQ+wLHC
SY8R/l6oeixLu+3IRPa7gUsfg86ryphnHmFOiZmdhgYhL2F+DNVZ/JBJKq/q8p5k
CML1EWHLyA3ddxCcWQ38toRhba/9qHxW5npKfod3RE+xF4CLpzHkO2tuVxNVycHn
3DnoyP6raf7XKYFUPbdMYCxKeBwka0RMriGwQ7cwe56r4ssceP0I6DvRjnpvzVKV
+lm+pQTPWBeaXUJDGsxeRDGl1iwjTTaTw6XUXo5vneEFt/GhyNAabgZwG0lm6KRu
PRO1ZP3GZmsQYBj2/1sHaPV42+a/kwofA2aP4oYavLHqcQzyO2p1iPIkprytbKLO
/E43YIxusk183MXHoRW77jlee7GaPtu03bUmA6CWE18/wqBVwkk6LKHbrb4bQdOw
kC03CQ9oIddJJz40bPLvyzmhHgsAyivS3mevIPYwbxPwQVQJTKk1I1hav4UtPf+M
EUQoG23s2HsCpHB680crv2lM6eUQLAPsQohvSk0sJmRGQYq3w2ixqGge3CJrg6pm
MNjLaG5V4zjRxRl8XYzDs1PPEjSXCKwMuPTlcC6o8OEUzTNvSz0j9Chcqm+DgzRe
plBaX7nb10+sMP8FJByQ1mhzxq/aaeeq4Sx9nHr3/iYOC0njZtlNTrl4d+15nRqw
W8JWsdp2uyizd716B36DOwITiZWDpH+lAmgIN+rpH71By6dB4smc6cEA+RstqGXI
eObscL/GyFm+f5wusB/ngpF1nkQjDqbiSpoZIueartcTXVFYVO3T1E8g1JFiKrIF
YN8KR/d+J1LGV3DaT44Dp1Gc/HaINvSQPpdHa4cc3wHjeur4iXuP6DmH35fijwJ5
Q5o+ApliZl+S/U7KSVUFp/+Je31r5iT7eSBeul2PtCQzwSUIhrl4ID6hU8T+zJB3
BUNUYZzZDIGA+tckDLT5OKlnyfKMuBlEADhoB0BjzYNP1U+W/RyxWNt52T1IqNZp
yX71J2V7nMqj86qcdA/p470/lKzCiXZvJY289QGUgQAgwUXWrBNDDflqIHUrqW7a
QD9WRjDf9tKlTF850QSEZbFl3YwhXIunnBPsL3h6KVtgokdtz20Zv1EyzVH49EdK
t9v0iTl5PQlTZo5GETVVhSUnj2Sjrjyhsqf+C82Yn7jwB6f2EN9QlukM4peSMKsK
iuaXzLk7jGGb4/4MRq197GeH80sqnJHoF1v3811jhpMiR6wGHfW1C6Fbcxhu2c5P
+EIVH3xFF2NIysOHUHlLkt7BJn1OMiBFfae0EeHjlmC4LgG+4gvBJG283PeE5lnw
hZXw9wRDP1iFv78mbPMb3pvoKGM68b9tw1EPt8efK5kWcuGttJ1Iq0/nAcQPYPFs
qEoaPahYZyULXPw9D/ZGZRwpLQT5Xxy8+rOaIRBmNZlBKQ+aSugDs9ZecjxdJGrY
WNF/S+tcf0pXYd6Ci/VuZBQLj8+i3DxEEJujHgBPdSD4sVk4oTRdavy+DKs51aaR
RwKdR+CdJgFwBqKzXdCs+30mpmR5XCLarTnFdGyL9kRKXeHBt3N7Aaet16LLX/HK
XnzsGZ+yPhml2EjDU96olNu+hRAm9RKcFtTQN2eZ9uiaAeEztXwLBnmHTZONf67j
H7vewLxJU5lk+gTBEjC532ZKzu2AX/Tl+RZKBCBY07tPZ9gMuIdsqzks/ubA4LqL
oRtZdrBxZ4GHzyZz+HjTYfip3wKtNtviE+45Oj+X2XpQwCnZYyrQcq5cn+3a1aza
9QDMAPNkVbPukI9FkFCd61Z3mx3vjbfPDjWiWJEcH5LfHQ6cjkGqDPQQv7GqpKdm
4emcLyOiZGyNENflH+W+rKFJC7Cx6JBXsTGPNcBKIHRGbaI+5SAZeQ+W2vLDBNox
QQ/f9fb+sv0HN99xL01aAoJ7LPzsiUDXymUJyr5nmNa8TGR2/XCTy69NRWUR1W4O
/3FGS3Jxqt8XwepeiJP5TODKeF4qv4rTFQ2n90pdDuwwh2G1XbYhg+LSWvZ3tCC7
Z5cTekutYlTj96T9HfpfQNCVhOhkY7NP4ehqSOOeKRSfJssmBIsFjEA303F8QjP7
lI06vHUfWq2STYaY5PNrQL8PggJmK+N89JaAG8DvncsNQtQl4+oZpXQ+MI57Gvhq
YtKVqoFZKcbDgUFKl7KqqutjAgD8pXpe+eBV1tCVsmAaPHkFgJXoimei4saFOgXz
Eg8QirvVVMYkKCSxGCbj9NdL8Q++2/aEbHuwwcM7u8fHnKVZpnIxVM+WRx1HGmg6
QiAat2izQhSzg7ZKi2C3xsbTkzU6H1aVLn7mzUDXSPbIWFIqO6EsAwA5qrK2ENdI
3w2MRCWzPMEps4Wr27bGLvqHpoOsgL3inwTeudkzlUOqApSlR2tHPYa02AZIHny6
4MJpVPel8upKIiSwZ9FdCyAhe+dmpAdJbQ914xdfrthzDc7zFBhWVFPN6MldXQ3M
22FjNpSULqz79LMXrcK1vihVwJNxxyfA3bKCKNvQJQ3vdXEojkM2J1ZfuVeUuqR5
sGz4KK8/5XKKxIRaj4L7mVJIESfIbjCooaQR/vdMjfTvxP3DLgLoavPsvvm9wcpb
boZ/INoLhyibcmWDzO7ISxJkxEMug8M8+EbPH//xsO06RlDargQ83VzRdGg5+5tC
BasU64FLcU9kT4y5mn3gJ6NA6EBhvpzZre8gCBxJ0axvBoSquQ3eXV6ZOAbVBYl0
PmwPz+RYR77B35UAQk0yqhtHBdd261u5eTnqc4wZBSHM4BxcSLUQ3fY4oOucczSs
pYRfAEh/i1q7tZ/uXvaRqt+doZjZP8ky3xgQKu8JcdIzIQ47YNhRq8GD0wHvPJA8
Nu4Ic7LNe7UVbRhdcQY99hJO4c74BHD4hGsqueifXxdorXAxs5WxsvSNl3aNpMpO
tHDeigmUU4XqM19u7kfmLwG3UzpkQxrwZVQtLV3kAxRIN5W9JoRVPoVOYtewfioL
Tr3cXvSlzv0uPWXRBIN8w+8faslqNvuSG3vAFLT8w71iIAxmo/FTTsov6fu/WkoJ
hSS5Z8ve9l9zn91Gzp6A1ZYFabmFGTpcFONNeUrtzd5s3wu6n1E/8MlwIGEt/Xc+
2bNhb0Tj9+7aF99cgSZTQre+h4+vknOVxCI6wdSNnq7N2LXOTO2WxXjQ//IwWYkw
Y/jnhnz8KJIxZFLTj71bNZ3jMZ35X47yEertISldXBq554e3URk/9mlOTl7TRgGj
ZlO1CqVLN3bHoVOST/QbRNrKrI92ht1sSTe63EoH6v6MAi56XP3L0UCQVH/1mRdT
zNuNxR0r6/IcW22LuqGK/uGyxirSatE3EMSI9Vdz9jPDLb8+ZDDkR+Z5ejz7Ili8
C0dnjdaj650XtcxRm/83brrFcOxbcJGIkMkzJxtl5WJctjhZssOkRTxyhqYWiRrq
eFzXgSTRGl28iJdFdE2xDnxxnQ/54OCDrhujBV4osQdOWOsQyCTT1abkuo0O7Tpv
rcyHJgajPTfpQnl1pkNVnnGx56ftLlr1strnX5g/EdITWwewfwkcfHA3C6YW2/44
yaumYIbTkRgOs5DYBnVvyQWgOMOsex2Eq8VYsuAhrQUT7Phbg0FDTDFdhJUIgxaz
edTABCmcwyCBV/glsOI3N27PtPNPoNmD9nBzxwLgVl0DJWQjVTZaBxUX/uNUzyXt
EHUkPwVqPyHFG5Ma+d2kmPmIbjisWJLgD+8MG9TdqmIWYHKNdnB8POLQMBDxSsjq
FOnp8Knbn/vI5XGBROYxiw4KA2b/GoJfUlMUlii5Ru0FB3vSZKS6cINOzjt99Qwo
S7yXb+XOXszmD6A3LjaNpJzes1nF4MqhhwGfVByXPYZgCBqO/Yt+B8Sj7axT/0Gv
VHDXVXAWrGnoTw6lp7N4QiUu98G2pGLtUsqhcn86UJzH2T/xM8cI21KT2nIQYrDQ
abGJAgQ2xaeyfzT8WfgjjvlAiX92a+1vzKRTif4N7hnNqGx6R0vDKbJICrZrhTzu
8gatLmiupdo7iThsqNS48n6ZvzsqjUC8FEjYWIkAmD/uu9cPuYAP0EyXozkOI6MF
e/yGqANEOAdatGoucKpLrrUPbipCRMGBtcByMptwxLnXTAWuBwriCQbggXWARTZN
ql1tTyF0x2el28jctBlnC8UjwwJARLSKztr4SuyyIPQGrFntrIHZwlGVmoyv7Oy+
rIpGToaMyXLEtN0cR4obwkqHBRpUfWT0VMrDf1CMgx8/vOc6MIZb03379ggGfPdH
sXlnEeDtLxpOY/ikmNqQpUk6U3hKKnV+Qc3iDWCYOsiPKSxaG4eMdzFirLPr9tkR
8sqA2AirdRr2H2cqmM83I1Ggo5k2zvmDBcdlTaNj5ddvuAsRhdI+edMVBJV0hEiS
jmuw8J4xuQ8ujC94LKph9bUP6/Yapg2N8vS5zwATEm73L27sWPAXnV5J93Myrbti
Ko3O9Ipsz0t6lI5TS00i28nhW8t1xzuYe4c7VPje2YR0DzNCeLwgP3OQ76G5gFRh
BE26Ucuoxq+Hr873wGtX9g2SzrVmj+8BVYc9jeTwTTnTXtfsTntxihws2M3lCayQ
LiN08DQXvAAo+jyNDdcIUnqoFZAgTKQP8kAs6cv9pCLUAgkLkcJY8URbt3Jw8xML
SodtTNY0Sy5xvPu9iaT9ODgWjldXz5W5vwX8K5P7+Hrdav+gf6FFJzNbs8oh7Vk4
0KdYykxHZmEQd8pSlFuEgbxJ2crfV1JqOrXkLwpHMWkrru5o9/ZLondcTTBmVrSS
9d5qJf7FBbBHN6cL2yMW/ypXO6UiynLCxDOPuD1zze0=
`protect END_PROTECTED
