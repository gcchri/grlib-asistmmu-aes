`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RbEW5BjhXwil12MVLxRj1k39G1kOn2U0p8OAbTz+3idZOPJFNWIMXnih0zHb+OqA
6FNLqafPxJ5SX28oFoPMuJuWmaxuYgsqxMWR+chct7aGA+jmsEEoawPPyyggn/R7
L2mZS9m6cTvK16teq02nGUnN/bvPyxnUMwDjDi1WDcMDoKPaNkb6WjrmwWMtdx3w
Vybx/28bN9HONyyXDPhmNtebQAieotwh9oqAeTUVAi+rO+uHEC8HYqCK7neRKbOM
9jxdci+DF2MCeii2rDri3glxuc7+NYoc5Qe75/ymx6R9NvHw9Vmp3WossQfhDDCm
1BMdYy057L9hXrFuubjiIkYZZpemrHuBou4VSLQFCjqp6en0YbQAmWRCr/1Y6O1t
bBW2/8746oVSsvGYlku0YNWvTR6FtCZ6XldNHS70xHk8/yg/fViidmsM9jo82HcR
IFx5KlB2IWDJ+MRMIioDQA4Irt5qyB+JMwbYTvgcmpfCoAQYtkHXOMCb3sPn3DMU
vcmWVCRGxf3vtRLtBLC62GJCksXsYu2njtunzUlD3IJQzNw/OuTDWhlOB0B/CaXK
YJGGR8axBHvo9Bhs9YkgUEv7ff1aQJOHDiBGX+WlkoeHoH4T3nZKVE7OZ/eLca+3
YnXRVcxGCYdIVLQrrfr9gSxq7I9g9BoPI0wCT/58Z3ZR30rtzPNxO9ahqMwU8sNX
MjUEE7kVQrQ9y9U3tsv8Y+szDzXebVD0r1j22dea9VqAESzSTDP4TnVDIST6QcmG
MmqSREXkOUtHMP1Ghie7JfgNdGnP4Ns+oGUXujh7iSC+JmXq9ryxnn6qETRfzR5k
32cGXbXW6feO66Hl2k2ybPrVTrIXSzAQ1g1DqHcYQTNh4XKrDzR0a6BGzZnvKGP9
JQpjT6ktggF4//CinjygXTqst0DlbWPF6dfIIw0TJGOQ9z0zyJLqepmsoXILY5+I
rwMuSxpXr83gJzuKG2ocTDNgGfINbCCdLzsF6Z+Q5rqO7iOfvr+pLk/LhGI6Llvp
mSngyd1CRkEKuNjCaeMAo+LAhz5rB2GhNWhn2+hQYRxYP3F7FWnI1BhmTooKmznR
pYlFbAMNTdjr148oIgQF6H/xpvZvlR6T9NnmPnevZcTBAv+2Hdjx/AOL24VgRAAP
Z1UjMU88Jsvk5rVCKE2uPHMG4x4Lz6nQUpZr4CoLeAqUP3xa9bIDSbEgUtNvQB6n
ksX843ojvrRDjeDkJ/R9/tdRfAaskbCilGAlJGTnl6+34ZVc/rn234MocH4SlNi8
ZgINNCCRulYRvlykxCV3xbOdHeLBegPXxWxkeiBN/zXCRx+lhr2J+0u/8xKpPsUJ
F5A+TRWHwDqnxLgw5bjWTg==
`protect END_PROTECTED
