`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lna+mJbbjGtekUHQMWIYyRR7RyZzb7AANkwYKs+tRZ6ygcVKj9CEoBeP3IhOEib1
/uYY9Dcrj4HcqM0S/b8/Kc2d30Nw16CEK5RiIcK6vo/c6yVyN7uFtx4B0YsYGnkA
Kr0Iow1HsrOiIoo92VORKABG4qY1lkt8g3vmYu/mhm7Y0P1J7D499h3McylyMAJk
0DzwX95amkKvMiz9bLaypCQetUhASW01Qn4pJg613jb8D5j6qaGQnbvDAVqCMWId
TJwL3F0nl/3cjgfPTUMyERR+2MCS6xHfZRgkXCQ+42/h40MyOvB7cPst7Lc6TvlL
qDNsAfOcPmytQw6fXwNWL2kPnJIwYRNzhEtc/ZE/XPdIdvnxXNvqiJHrY5d4vTEJ
ejIuvwzXPrbCspVAz5qEZ8/sOsCaf6SfXCLKIBf/GOR/xBjAp/9Ue7nBPbSMXRhn
rgladpfNqHr5j9tKvs9OxUWZAyAfz8FF1EOQ3Caek6cObUI4zgA3XAygGuHlbEFk
LVrgPXPOUmK1gDLrj5Vdgimp7KD7xN8pJ0wsBFc7ZZE5qWusHtc5hZ2BeacZghgv
caJn5dOX8a2qOu/Mzp4N+M1XajywCF5ACN8lH8XGbQK3Q++0d+GhsXktSDltZtd2
9hvm/xVl/HLgzDDynOr2PA==
`protect END_PROTECTED
