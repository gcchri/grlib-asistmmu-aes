`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOVP0b5cN17tcKNiW/gZ7mT8FGDAPa9MMELFYgQg+l7HbZtlmtSklINmi42cmbKU
f1KxOsLK1q4lqeXhDsr2I7gnWtl6BbuAOk14j2FtUKjPhpuNIglJlePAMGspCkgR
CiwWHyw0scK/2MBepRRo9KEkLbCihu9ojM8oCaQTuXk5oki5ETFzNQ+L8bNz1lDM
3VXVHR2PGJw8SiSoiju7L0e+rXCFEP3Mb74ONOezVuIaof4DXCDbKKDn7VZk/Rh0
R42446GVqZ5wbHWxvNNthOLBSLUSudNd5H24yBagOR2GhRFiYLmvJZMPXcAUdbo3
jJAofTgxsnG13Mvw1ixaTKufdDn4wb0U6en3QJMq/6kojBGbHcGOBk+MalGD3Z7w
JxraT3O+GLp8sLsi/CxqRSYPJD0fRO8bG4QqC6QO6ab8EkJFP0eUX3pH0BRt07Fn
/4fqaPRu8uX09HAysYvT8q9cCygz3fd4xpMoWV1efjnKiBhmdxjYmlF87VRAd8DY
C2FtBSuHodGzd1ixxWGz2dsAyrLB3ACP9bku8YfESRhZhAKb409IgfFjgFqW/6EE
TCk9jPBu8aeh9pjaJOttI1QkrlQfydhIhus4nKTWTww+S9c0/TCDIh8YasksAnF4
lfkpkboxpsuSWzE7lM8/vY5t29OHGYFhXHPAmugpYoLwDg6HMATma1U3l8NDeSiN
I1VQsoKV5V82IFYPzl2BwYRnDmSsN54iTDnxFADPDaZj4stV5robGV7rUm6MOOZV
OrVfU1vJom0xhwQaLl4jPBYRk/fSDRrsFJ1TKIz1dwaS8JBvbuGuN6DDgn2Zq9mV
5owiOmbpJwLXWYvy8kxI+s1eMA2iBvNass8fKMnYbqm0LNtHQv4JTVBRGot5zxdW
1TDZvvVg57ohJwljtnnsj+uX8PPQiO0sLmuaFD/8+OrmJ1yoZckvCAH+eev91fDx
555wI3rIflURJ8/wC3sSaA7mm+W9esjP4+2CC2AW+rkSa488zH2dlRWCHp3q+Y86
7eqxx/Fiq3Luiw2XQHrGgZ3ERUoPcW8r4P8sWVE1K2Gn9la93ur3HJ9kImwgVFRJ
JJAxx2OHoszxwKT4U5K0v0qrtsA0DGK2lBw7QQwsBEpKgCNKzy/7/Fue5YGQ6qUg
k3Uhs7RX1Q5fGZHH0m21S5D9Z8tOXJRrGyLlMo9a5mmz6pWc93ulEjc16xiHWf++
7eOE0Q9Q+3WDm2Z7YnVH3m7rt8ti4pQMVCaNn2YT5/4wz2afwrHznxLg8tZJdDus
FKPTtHlmqezky90xEIL8YzbsnV+62V32kymbHb2nYx0lVPg8iMT7BUMYuclFHKis
AvntsGTecTLW5wLUJg6HuNuhm1Rod2qOTJDuHwRHJlLRSLDQukCmla0P1gIrGlbU
+i6T8hQ0kl0h8GMdmoiCzw1JK/LBiE+/JK3h8753epX4A14lZZJPdrxeIOSTOGHm
GULiTTQH7GRKhYTLVEqDBJem9llypTbRclP+liPmG6+IitiasilecwoYJiS9sQK9
NFhYS7XgG20ViSc/U4kp4lyESzaTFrUcL7TuPr7Gur/aJyXadzA9NTd/Gdj/cYgR
rcUmsWbQdu0gl/WEn9hpPKXBRxIqwooK0JXNe4oVqqHfVDHbHTPhvWvwfG2fp4hd
e9q54gMT7TvUhvAkocK9XRztIDN4foRMh9j1kfiV1W2O45nIJr1+NB8INaOnvtmY
9Ha683x1wkZjOXdc2jzIz+X28GLLSoRIUcK5YrjfMctxIZLUyF5vdkduLupx+NjB
H9uM8437pDlAHoppgalG51nHDdfJ8SLtZCs4+J3QjW9I7qDoMSEjc/2egq4MN+Va
eR8x9IkteyVekdIMC+Kw697Ih8xpeGf3oGf33cu3yAi/141rUGOTeTUjlJ6jrbue
u0LTE+Prx9qQkeXefvmQHgpFI3sMzYjsp1+qHkjQmEcneX6b0Iqa9QJtQto/USQZ
cbW35lQCaq5nSgQ3xD6cBMbktwXWPp5gg1N1gjnSQIAQ0WZWo37QAX1BUmVjAAFp
B8hKMg1gpBX0SJOiaBLIEPLo5uQp4LXjHmgWvKxhe5CLkZwXANWIwdtG5Hba6NQS
mk/ttBGxorJ1eL8vagkjts/0a5YEMjzdmFl1Jm1JJjAOQk/HI3Ctjv9tr4xEf2zP
Ub1I6Yf6V7LtJ/35mDI2ru+yQlgOlfqtDNvJdxmZ+JsYG+6mpYLC1B4QFvc4tKi7
C0igQGfYDWOGxBBaTAxUUsRWKFJJpLyJmU/cYktY3MabBC/4jb2AFHplf5Tzl+Xg
aeSS+tAS9XSYn/uhV92f2XR1k6kak/M/cR+zbjNBxFMsyjbeU3DkMwPeEKyXX6gL
bc8FcPbmYMm6Usz2sDmPrKqA3eZcXWR+cTNX2EXdS3+uL8WmOEQMi9q63Zj5c89i
kVjikvTJ0Qp3v1IDxoNxhNbhhM2pA2sebSR/WGLl9ASHykyE6vCw6FkBy7eddC2Z
kQU8Rn7IsdmvF7j6CY6UjdUyNiKvwC90Wy2xSyyMNM1N02iXWdcAMf6yqP2T6UB+
065WnHsNM1gCC2LJxX/jVba0ExKUFy0haludOa7hzdVH2xq3Gaz4Ay0mCIrwLXpG
gqCcK2nURNlAwYoAJnlZrUoodN33Z5KMQHWf2AgWL24tXNTHvj5nvPrhysi1CK2N
xdrodW6EFwuZXZejWlRvrUZ8/nUVbBczr9qJhdD8HP6npHUcTW83OXXLSnYRImLS
7wv/PgGOL4PINQDkLUBoU5YsfXLB0CeHsLEESSf8btVR5jU5oUBCaVCffr/MfCCy
6SJaCvGHKHexXnxUm/TjX0ey0MW1eE3ozp72M3SyPWW2NuRO/hhaiUA4GuVUEBQh
nQQnL3VUULoDUwPkRRvYMN87i5K65ZiIHBXqS1Y5hpv0vPnMo1swBNm/5YKTRKLG
kzaVKciGmumxHKAYrvnUcLAGQdbEMI7fOtgqOVrr1/Ao7f9TKZPxPLZgHHJpUSaa
aO/DRYuNNX299YamA2wRuMkLHCxhTOjiGsZcAmhOMxakANeHf/Z0Ho5NBTLb+CT6
pRDyQn6ja9/aEDXhCPWlOyAZvxeqbrIVzTJ5aqJPEoAtiw7eUc5Jnkapp1mQpFSv
RIVJCSBx0LSxwVZLQ++Kw+5qwEJO2xtiTFXLfqvXDA/CcOB764Q1DRodzVt/q+ds
EpUnfQJhG6Wkp7tuyDPDS6f9tphFg3ALeIoiMstAh2l6MupAAhq3nBQrU1Xy5r11
0XRs89Bz+P3BBxDfnumJvACRRv13J5QEOO6aO6IJVJvEvHbGIkkPsKmQtFEroOWZ
rbKXUnwSegv2B7n9oMfrEua7QZcotf5Pz1HlWAwdaeuMCNVtYCRFzhZhkxTIPYIo
ZXoqZjRY2/vZhR5HMg9sQ4pLPNcmVzKASdYBKP1cH6N7qJ90QtmmC6W0YrAsDwe7
kOVLxMzllLxXPAnXsBlN2MmiZ4tC27xt6PRwoWmH50lJXqGdWuxJbEl20sTq3gc0
ezk44i1+Ioh5ejAtiIqPbByZNKbAHRDo9ekBClHgB2b0pSD5jFURkLxNY2ITTrg1
yJaNjRT28WiwSjy3rePxMg6MuRp/8zU+u3qgYGxHtZrx2+qDR5sWSgrYMRH41//W
kw3T7Dy/dvVsc2AiALYR3HAkQcB+bsG0J5r4NT59P4A=
`protect END_PROTECTED
