`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
llwofoILj+nEpMHY4/iuLtGpNAFT0eFfDZ/oJi2R5eVaY2afnoUitOHcJau9RTPE
HKJTqLz3qgNY2Tr6fx8PgKY493K2nQDSGLpYIot0Ay04tLEBGlUzaG0w0Q+xdnEG
C3QAYnkEL0jXqvTY7Tf1iYe+KJYh8m4wApkxM4Mr5wHbpBOCVv5hTlmCpxtIR1L6
zmqizoNcxwFjv9Pk7QQHx4RY/2wpI6FNbqRi25hLqX0cmwva3g3gkaqotJb0OAW3
yHHEOs8bNYrTkaOMl5YLkmCIClcUG1YYrQkCYQK/aKXgwXAKQpTzO8v/5Q4yBAKN
d70sQT6ts+iwsYHpAkJpsFO1WLidior1rDDPxFg4G14A2MBtMhT3oI/RSmmq8eAv
jfQ/gAy5muTnvQRb1c8VZT8lMRAT0Z3KFbz9nyUoMNMsGlso/HGj/TZ9SvtFRqWo
qY7Ru23V8pFBTAywg9cjZamsmG7SP7RtLLsxPlBFrfVYesI9g8TyJiBx284IBfWo
thUz3TtW5/sTH8YMEWcKGjQ4jo/3jK0GrQEhjxtnCPI=
`protect END_PROTECTED
