`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Oe4bvZjZOcyL8kx1WIRMUAcvyk4k6wrBYwAeZurh1PHsq3lI3G/R/PvQY4Z4xCh
JJFGlJefn6S6osHItY6aNiUTlNYPqM79wVPSxTCzrtbfWtIDgV+qGu7r/UaW6A2N
irqJd+G8J0ROWWRpiQsxmH1T4RreRTLWl7yiZMXAiZWi6CZeqdu7YfZJKKcsX6SH
VWrf/0Dn3P39YHmV5gWWhk9UWrjaCM9tGterZfHpSK8pO/dmE1uYoG8Kz1h3i2Ho
9VCbLxZn6Do5E2q0sR28Sxo9YUozC6D1QqjrEysAJd0=
`protect END_PROTECTED
