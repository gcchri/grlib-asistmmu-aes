`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DHsadwBJMWHVfGU/txoAdfyxHk8nKGWkXJH2zepqMppkKN7WsdB+FZTE2oZb4gY4
IGXntoh1YbJxCuRw6EYxgYc6jl+9PMg1+UU1GkzoI925IsstL6PBNBMMkbNmYD7R
kD/Tfh9i5Geip16vEv4w5bfetM9PW0gyoSTzlAKbAC+0UC2KuPBKrYWplmCzPNVR
Y3yj6AeBbdXlMOqnuL//Y903nFUmX1eJ7JVHgZoBuXKnx/z9xSydEOvSHs+zrBTl
OPp2QQpEuKjBz7i7IzkShTChAk8ZD4K8ACAsHzFJ+sDbGQVUO387+oALIk+1fXwK
wjXhG3qW9WqtQkzAiO5sUV/HdtXRq3bLJ62fqZ9WodVbq6HIdCJJA2jRjQjlHJnD
u/o+GoDoOpviu6YgwCaoLrABF/GWfuxBDIL2zQ1I6zBRW1y9SxiKJeLW4yYq9lo5
38kJJonTjiN/SfJSG+6wtcga3w7THN7laxIt3Hg1Vqnxz/sn0sW7NpH/j9uAOAMJ
XxsuFT1t0CgHEdA6f410zCx0Icy9jnyrHJXE2ewxBF83jpBhDYxBMaOk3fdPvOk7
/zf0EXff4kYJnkyR94Nuzu9/NM4hGFlmWsbhHP+G7mJciI0tbFqYX5C5D9v0RVtM
y5zCi/YmKQMsbLappuzJAo4Ls54AnNjJocIgGWVsgX8=
`protect END_PROTECTED
