`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4BqttiwvMadb9bP0KDVfKGlIvXT5Ey86TwVTGeWKxcoMBOaKYJA1J5durcg7fhQ
9sIsHo9qn0bjjJOKJh68FZ994YkPTdeDnLtljK/hrvhr4Y2F4A6rPu+X/luNaz4r
wF4V1d03r3I6ynUTMca9Hu5FoCbatGD+RUirecb/uYwqz8gtDv3qRilV7XJc2TnQ
sk22AwUnw/e9gAm7rF0aWGgqPesn/YNo5AXGbqjrumM7y8VdSJh9EGHmx9kgxadf
FjToL0c4L7jxLtuCD/Ra/b4n1lhSTPIgrn29jMsHltDXmYCd6YKxVIbbeIfSwZi9
`protect END_PROTECTED
