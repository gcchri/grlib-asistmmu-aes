`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9VFjH6y3DEEWDmmLqwyPft8No1I2OM+8eV5r7tFZZJyFjlbXKy3xY0zqgQ0c2azo
/3P2ukOB0uiI5Yc8N+o1sfUuvDVmhHbZq0UABBk5aDvp9sZ1fCrUCXP2Jzv5wyGb
cqDYu7QoCCuczlKhhH+9yf5KihAKLhiXFu51jNKE44wllMdMELtO16MAT6dZWYDw
x0H9u7JDqEsPyY68HghCbeN9exs3pXa0+2KhOzHHFUEejYw5AG2m+s9bJC1vRVcp
G22CZysbXK94qXxasz/Gl3mM0BwhLjvSWb3Eyw70OGTrv3ojIpnay10jWS+dcYKV
mXYqXEvpnEPfU4Wb9JP7RDtw5zMcjUpHSgFODIT77g+4k9gvDHvtCSn4Aqv9Sz6k
FErQkqDUPfHHZtrK90/UjIEtNUyoaNKDtVf+bhTudCk=
`protect END_PROTECTED
