`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
80Z6lrdfugXbMPECf6b0I2lJRkwkalkoS9wHPHeMdCfBMKOCP/fos18pNJGij4Rb
rG1kCj6tdWXPjMekbA81QfbcL4iKzR9yGMmmGpdPH4OlIH4X00t+pcqxpkke66JI
Pd6UVSpA7oLE6H3sqcNGE0KgCjzJmksEudBDpjBIIlbHHiYHDZUx007pAAhq1VSb
P6hKP1kOEmuDk4kmXpvWZNj0FnufzN8K0mv47z2lfupKmqjB8wpCKr5HgiCrCWft
eW89865LsyiR5AFuRZltE7eTP8l6QggXEXzuAOh4ynyjGyPcByMsodN/rYZ5rRYg
+d46iDTLXcKQvfaeDQc9Ti1lmpqiTzqPAH8OW9Uj48d7BToYZQ6tIiqz2L83TOzg
MozXt3ImSkUT8LRQ93XMXFQ5GRwLF48iHvZ2Y1T1UV2Vs+GkHjWWKYijVq0reJKU
bFvqxftBUN6R5Mma1NDeJMnKZqEHgqHpvgqXU3OiyIwHhohXJ4DW3E5Ei0DsZq1T
m1hQAC042IqS578Mo5t7TkbxWU3RY4H2+hwd3XLE/PX0jzxISCPeRh4FoB16o5Np
GTDlSTyqrxNsDJlopL6PJuV291ABLIbZOzL8rb0enwHuMAQrQA+DE122KvsHHvSe
0oGFeuZ5kRPVPsZHCyeS/kj3BFpzcOB+2LtLq15lmMafqq8d3L3NMKUZ2pp/7hYl
r8+JALQu0zgQLvIW9a7OrzWdSFY7eiyQFgScDaIjaFSLw/Swu/h8PdXQQwYUuXdW
T0cP8FuMBMN7yKWnECSb4T6PMkGCagkEJJJxRF1bwby2quOef83FfFwG/KQhSdTn
fGNT9d79SzNW55X1NaLFMfX2v9uc9sQUN5y+SVspZs+V9PYNmXw7l/BHfHOWCftC
oyVtPb9cLOzM+2bjIwn3UftioI8PxYAEumPVebyvwTp5vqm42Xux16UDM/nxHcud
LZva7gqbYBFRuV48SlLA6ktEpxOILqsHKSQiLuzw0tnQ8f446a8OdcxqXUMETcSy
st6nUfiUJxdTqMi3K8vV7YTHqDMsmwEk1W4qKizXgxHpTGCzQMyojoVLHwTxpVzI
bPqxLzUxl5q5AXRqJjvfRaC5eswOR2JTUSkRp44Q6NLRekD/CUqbkJJMCo00JUsv
KqdT+B1uJ7toPuuFBzg5PYQuk4Hw3jAGMo7+5zew+6+K+wgG5yCmPhmfU30uWGa4
FQRKDuVNVapz3gbUV0cCh/ljEpm2E2HaU5sjAuDt7R6H3p78zqdMPGEHgNSR9gW6
YX+Ep8Y9M+pHIsdrLpcOGn46d5e5waVbonBIvoJlPuMaXXaT9v91qOnFFFESIkyC
eox4A5pd1hAT+E0emp3Dt0JiGoycarHChKw6C1RuqtiMJKF3o+ccGh67qyD2NOru
vQwB9E2W1cj1CXbvYC4mkp4AFKdXDROdJVUspB/fEEZq7bczDhhHzbgVx/1UWJir
DOBBbMTfHc1Z/x6IysX3SUxlyE3f5ZUfIbeyWy6TwoDlxr6UJwADA9RUN40QqUTs
GU9rXu6ZzvJAiDfXCLpZMGpHJUjhvyuTAxyWWr7JnhniH14oP5P2qXkFYYeh6wCj
cI5DmiA+1idtcaRIMgQ76+xsk74UPbldlZVaUIjI4mzWvNGbunE05nPKvXSxnr2G
xZXPyCuVNi7Rw+V8H7YkRRPjQ5sKqCuG3A7mbHo8g5hDERJn6nk9J5/Ada5Y+uOs
1sg3uy4+CF6WJJZEpdgKLph04rnW2kfOstlejTBN9BWeqz0aMyTMrtHRoMebTxbp
iNAi1xwp22GawKEqqPpBZpE65LXKOUnVVRENxWfz3NnEC/5evlqJs2dvwskb9Gu8
t0a0lpITfotDjO8SENRyPNnNDNqVonH8VaRLoB7EhW5HXweDZVXtZRl9aUhcJWT2
xHWYwWkuZFRSFOXGofAiuOnDsDz6lfvhBRXHrFN8G/ihx7WN+rjsTGunUffAn1z6
St2Zadc4QrNb3MK1kZx3Aa9XtRt/Tx5G0lnF2hgPrl+HLaWZVYeKJ4ZxsFrs1qk8
vDwagvTZHgVWuIP7w/mbkoRWa9Z/qK+zOI2rY6ZJIfJKob+aQ2OkHqKBCMuSCfBV
nPGkr7R+Z2XFrVKwu7vaLWO+Z9ZidWLnmq/P1BDe3BbQF/ew0kgUc0PFrSCEq1Ho
qDlJXtSe1GcOc1YeX0rAnc3SSM9wbw+feLScPg2JAhMCySEKAJzQBEOKwEwaRmUi
OlQxVThSEHpIOgC+SzK7W5xlGTFvNwiZu2lsDx8jNkcIE1EkqkUfcGzYOqXhjS8y
VwOwp/fgqZ/Wo7AtcgEDnTz78KhRKoguTaZN6MQiZWhUylZpC+6rUweS4oM4egyd
bg8YJOWp6OJi7qfFV/5ca33vOIsDBTf2HvJm+jGhiBP/iLSmAgmPVQEODVjH424O
6HibtAnvoNBEkpz4kfSQqIx59EJSH9zeUf8lFlSohLBeubCKRhUsCfv1xGqrz0+Y
6J6Xdz7Yuv9i9zXcMlilZREBC6w2LpYIkpRZWRIBEH0sFkhSKoaJcoDdg1xm/EUX
pxYbi8hzWXlod9psCT45DmS8lUBUHNToNL546L+sf3KEedVx1KIqmQlyc56kcb4U
mfrngOTS5I/Zb87p3xKMhe3MlWMBEf6wuRHzLU1jp8beqIW9zddbnwPc0KPqZ71k
Pgst+9JFeh79XJ/g6haV57BIKpl2vcUapc+c3PuQs3QFRMd6d5WJdLsQpGaR/7vq
peMpDy3wyl6xNNoGwcmKOLgKs1qZCFLQnmzcu7HoLXwQpKVXrnOKJ5QHEpZhqBxm
9lD4NLh4PpwNsyRW+yHNwPYT48vIU0lvVXd0lZVR0YmUW6An7D2ut6Rq82rV0S7Y
XgUtsntGdfSltsbqRBZhwgzRLzFAtHCG7a1kC3DEGOchxcUYHqlVtUkBAtjBsJZb
ttp3g23q0Ji1UMi/FpLncZTFFv96CXtME6n5dSvcBDbXrk4yTO9eDE+pYYntbJfF
XQhkkJnuICtN03oxTCaIy9u2F9dl6UhL0YbJQ2eQlt0tEXVvHzNaBCoyDjoBlM65
IyZT8RnKz9IRVixRIKrZe/snxMtmyJSwCUgSGf+ctMZLctJsonfrZb6pj2BxFhJh
Hk9/m4lffjjuPmFdZTWzAGGg80yqn1dVb30WKlMR9E2duk3eKiMv6x1DQg/fSD7n
4lX10NjsBIWNJ7WwY5BFDj4+UYcwcYD5/P208Z3Pe6hYRTguXgvyen+9xIhkLZ/C
lVaF4Y8NH6WPF1JxK8x62eD7rm0YqxCFmel5AyApvDeHm+4QmI2BNA1srmvXSCrY
kE0F3JFbeDnUhQrtVSMU/lXEqcEPESSd4lUX0RgE0TFbJm4JKFwhlC/iZpxBfGCS
JEM9gI4FTwPaYZgFo3k1whQH/GwWNYXS2l3FrMb8p8XNfFIX+74ybfkCtWNihSII
nVizYfdxAj1zY6ncnIvBeeawiSxFCw6Rgx2gbARCKlMK5FxYxUSIlscyJcQI9Qwz
jZe9VWF4Tp4Cr73asPmEv0m/ayOXKG2Nw4bTYEzEYVzstb1aNgw74l6KM5BeBEZO
SxR8fsqpnky34hFQA5YE+8joRIZHzqbvJnB8+mrfpHwlh3Lj+DdtkpFKbFv76tgt
janfp0dG4qtXCoKj6vDf3ztM74550yiNX9Axc4Ivn/24JYuzs1s44Fws0sbqSqgi
qQ24IQkoL4t804/SYTPfy2q/8GW12tXFxJgRPgDUhYDrqYkzO1sLDOMXHHDYzzpV
gIviOj364ePLOv7afsP4WdhPLoKrktQrm1RJuAuUeRDqLBFBCFNTD3K6DgJF05gs
vzeVwI7wvWhs8rj65gWv626A5LJW4qjZkIg+cD0Gfr51wIE5WEBAUKs6n9sWqO4v
3JKm3ab/8A2jfKXsIVoWs3aU6z4KD5Ov5/ueirblLiHJ+fQToTY/aDD95g4FAqvZ
kEGc5U/EsXXFrSC8XAfYL6HXsdxVLurosCq0lEraES5R54AsM1V7wLtTEe6Cp69e
ilyXm0SK7Kf/M8jQWQm9cQQFbM1/lpSLx/TUxKItNVuMBzmHWl/Itv40KqZfcwkv
GQPDlEXUedKjp+Myo3VEYNo3dUNEBiJ/V9CTAIXMtZvU6R8xPdmXHHKMDqOfN5xc
/LISvPFB/pk5oLcK/Mr0J/diKtWpLvCGouzN+AyDdhbAX1fnuJ8J/sizJF7dRO5c
XN12nH8aOJEwGc3oySVTjYuY86u+GWhmbae69XXcJR3hfrL+ydnHBx5o/+6SpPRx
FL6scV92h65HRK/ODjU7i1wbMjfxZcNpEVkM/HJY8XkTioCCx3cKfZV5OizYitfx
UFcg9jvhU5zI/ZPZH5cPO/ptfVylOV3xvqH0iaDVorFscSGtV7ZKy2kYQteHa/LY
Oqgb80HIaJ5iiF9nWXFIl9WIWUWUUSGwrbj0YFqHtTucaWmx6nRTMw428dSIH3Pw
Z+J+m11wBTjPjzDeo6WmeUHMq5WH+ZZ8LV+a/KfQvHeka1djklcj5LYvrd+LC1vq
UpN5RA93BpZLS3xzKlkQrxEMyR08OKJCsPhTR13oLw2p9SX9Yw4ksSHcCUA1dvuJ
B2XlrxLa7E/XTLs2DDbFRMlDR76kDI9kLeda9EuRnp5snxYBvoMZsIUqsSQPyutQ
QCuvJZme0Woa7NMNCn8275WnQXqzGXoxoedKZPLdvSkagD/e51K8u7hCNXG1R7lv
PgJcw5v/hDJhUmc+W3G01jsCfy1UfYPqeHqusZnNOxiSzwgK6BKod8MvECkwC5mb
ibIZrMZ0c3ke1bO19avSPb94Ko+WbtdQLF0tVJe3yyqH6VbIEx323APXwcefUeHS
WaxRxV5kve94xBh0AdgL5/qiie3QzQC3BdlOagP6hj3PvIxCNuVbMwaIki6Tixhe
fQA569XmrvdHY8Llm8gtYGijkJpFrpy6ZzAtFMFy4wiiHnDen+/X3cRqUEEuz5B8
6LabQn4OFcP8ngcKP9pgqtoR5H7LjU9ustZq3SkBpEbni1UEhEGiLc2KvdHKPAlG
oy9CAEWKKxcpnudmh0/Dcd8Pr+A6WTE1oWyd6k53cqXJClERvZTSiLl9rdxPlJc+
Fo7XmAmOJ5YOpbhnqIBLMKmCJDOZNq/5zVvYcHNCH5wwQAH/+v6FeGE13+DIW1Q1
8DmPmNxedi3RKcMIuEEBMinhNXNO6ZpOwz1gN6I5idW6up06WRR02nUqCBj9cfn6
W2N1iU/HD1PCjkb/RQea1bPO1LhrgMXhH3uQbD2CbcKAMSejj7fyjDjX5j356PoM
hx8fcZhPjLG7S8ttH76YiYhiVok/XlITOR9Al/8mRh/3mQTpSOjHs6D2Hio8J5vo
mfUF4tVsdOVE7leRe15Hymf2MVXg8kv1XHBsZbMee4O1oXSPGH1bDAHpN1cEh65j
JG7c12A4U2+VCEpHtLjKOt5ULXfc4umWKYYOolpLqR5OuWtz1wQMXnapjsMBN6U8
Obd9R0xPFUhSxXPwjl4ltRGPK5orU+eHuK9b6naMZ/I7KJy5xpyMquyMLgAIA8zQ
BDD238DoKh0HP3pxrfjTcxquAyWH/WwG5ro5ir8yIDMtJotCXKVJPJkE+pn3KlZJ
M/BVNJWnwmqCtZmJ+/5tWB6gxmqnbNHUmxWLyyZG0rM+dS0SA6WUTOX52hBhQ6JX
bOinB8JE2QznEG2OMUKpRLAr53PbK9kUEw84XqpIHidPQmQ5fSpad8A9KgUwUWEC
D5Sp1+lY2vwjVFEWlFOSSFmM4CtNTSh3HLWcX6GrzqHaFFxNArVUPhg+SDUERzFP
f2KzHsHCD8VEKugwTANxGITJHC9KUkAsG3VtmiAA+DcNG1OZuKiNhOnbSYkurc4g
f8GAB06dzlfa0ySHmtAm6RBRKDqkw2RDHvXh6MMLC6izCZWDizPbXNpaaMNQ9wGv
sB7ECLDuW3FRdzNxwCnX20ONBcCmErz/OR+0SGlRJ8s9LEUa2y6TVwuxE9MBSoq1
UjrsQ0otroQlMbshxtuxkce0H5mFfCQI9dPmoyH2ke+J6xtDKthhrc4bHnlZlxhc
Vct9JoKiTOHZ8kv6L3biX0WbxpdIPPn+8IP96y9uHJ9mj3FOq+2y9jS0jGCNrSpg
EGdLF15bqMbzfjFnPwg1nbeBUybScMnmVrdJNrzf30hILwh3opTO2M704dwGgkkZ
OmS6sOoBgTuEx4rE1LlQBsbun42nygLF8RTJmgHgUlPXl4+HFOncZ0E3YsDoZirO
8IiMiz6bfq0ycIJohaSt3m92OiLelHeuENSVVQCTLHbJrzssqjtrWkfTJ72mPVc1
1JJDbKLO4c+O801QRv0Unl0CvONfw4zfUr63vGCVYiqsqUf8KoXZomXRc3t8Oarn
GVqA8fnQm1rtm0KNrnO7eosUVfLPTf/g473EhGmCDKZ5oqydveO7uthDS8/n4Yqb
4mUPUxBbuhid3+uH5hMTbxUqqVlnY57EhIALs2bQn3PdCjzezaRIe0Wypqi5Aqgn
QIUE0+A72YUyqkUhKouSWPE7rmHzoYGwpKKMTjxyFFuq5mxkkSskdoFFek0QgPb+
dTDyqu8CzHkNtxBXDm0sxvMt4ZZLF31ogvNy1W8bxuyhrcRwEPJEnZ8UwqvdKmB8
0LHwEg/+Z2rt8zzNeVYpFm8PtiB8UI1pF4gDNydHJfDCaqDWf4dcygIi/jTVhrzS
RE1e3eFZ/+7lF8bPcX/w+NtVuLWQaKU+4u1UkIp8T5Yqb6mpXghZyWtMPBuxlCpM
RjLhtbNcpsmgkA1DcFSZ9Zme3VaabFPY/7Pl/4aTS4bG6v39dLtuNDsEu70QEpV7
1anu56ifIXSTuTW6DyePSwPN6mwvXQPh6PRh+8oNuYxec3QbB7pswcKWQDDMs2qJ
XGKRVFii9FkRrBQ6FFeet+/Lxas38aM4uYYUYZqhCAE31xrmjlI2eabTNJ1nu72h
0Punf3nFoeahug8HSeaAedajYb5Te9rdxehRpahHReU7OII522VkE8kM9iBwPv7F
H8D99oqBAudgVXtXy6m96eFG4HR+5FHSMR0hd5dyVTYAHCG5mOMdPY7ACorqvGEU
QuY1yBug0850+2c/mvm507TqBd+z4H1FTMuDcgLhqi2FXuHExF8SYiXVrBnwQHqb
Y7lfcpQSmBhmn4/xOKSHntb0clw/WaIrRem6E6FkEGNqh/zpvUhU0zdVFGAH5Im+
EHlhKfE0vG1C0nIOTiHHR6AM84oeXQP+zrVnzd3p4VANsWULCCxbU5BR2fjAdNIY
lasUO82HM6lM1MBhe1jGUKM2EGrENIFK9onJ5dZIH0OxrgrBQibJDZe6ISLKMETb
cP1JVoIN8sF6LUZgHW4KH8CalAiv/zYgyO/0PMZoRTJ++Cx9q2jqY/nEQ2tlN8NM
z9JTg+V8zcaeY9+fmmMsz2uouKGWGvCv6cGmhBmQ4XMA/cTm8maRI2vDfJBfUOkl
6vu8GddZEYyuVpXGxjhFqZH2Gvhl8ZW0vGCzv8aoCEBC1Oyd6/VJHjt01AJWcSw5
ljea74Wc2etkv0kSVTWJVGf2QqlzkNWM7djGR4Ez8ehPT47PhHcac6dDrnKDB/qA
HShCaVhXGektQwLJ3hC7ONKw16KH/kLQxOoPs/ngaHs2N13M4WCOLYNg/ZmDBor7
9vZRbP58Z0/4lJbNyyubRMenVEUiWEzDysllmsueSlpabpyEg5qSp5phF26e7MB/
XOUjqThgUqepIxo4ZM4sl5kJ6qzGPyFWfxTS8sATVpFCWjRluxYBMuJVq8r0llEy
Piul33jhVQnwQlFVtD+pUkGCQq9DOXBrMwvf70fKEnBtM631rATpQE48kGSQvPYJ
RmwiM8qkWS1uS8ANCPyMbdFlGLgST8b/gr7HCXLHYUhsWzxfrrCXDvfsEXfwBoLv
ZI/Df6iN58LmR4WIt+fB7E7mXNCXK7fBCfwiiR/VZAbjROsTI8oR5J82/72rz5k8
mbmlhhH5JGlEbJ8GJTwt9gwHBRdZQUywP+vxJlB27y5HquWQPc0sKUglYccwqD60
1nnmgx3HcPh/fWMX1jPe0f45e/6st2LEEnbOBTo3ii/I2m9GQ7y4hdgL/d4nOWcJ
rCCOcj6jXQMhed7zECf7nrklq5Bta8XK+bf2qaYBKFdKwKzLUhus4MnV3bLDTGvq
7ZlA+QIJgViUggxPei4JonpCeEJNZLp2LNTMFmVEjxmMxOfEiQU1N8ultk/jHaKH
NUuDeBUwnjiCuzqeTrAjnAlL4y0LvonD/ojjzKAbTU6jxY0KJ+iHEVlqdcu9JnO6
aefI1fgGF0qbV/AFL03B41VH7rsDSLA2npgaT6YLcZLgSVLRCdY07AiGK3Lx1Kaq
cDMBZAD0sukWs4wHqwAW3tGAmy3MuUuT0hEE74LZZ3INQBts8vO7ntP3HbmB9u4m
0lFoCAjlyETQZgAkHqN0ESUWE8Hj5H3Jz/9ddWCvIxv/W42LMPgwvW/P/qAdyfIT
VUA1/k63DNcI6e7l6J5IOOI/DCXbXJVVDAEHZo7vdDqOCt4v03z4XOsL3ycJINAS
vAB9x2zx02xmDRTIkZUcFv91QXqHBfXkADqRVsyisa4uz4UIt6LA2A+78v2ut+7e
OWKY6iLEbVmiki8XMvauU9Qs0uZh0YkFvqrQyFkwt0HZCZq/+qYESaWYah1H9U6k
jgsPJ+YQONr7jqvDmmOJL2Ne6mxzXGQ8+FFm4Dq/LV5T6Z0iRjdyPNTdBPc2Aa+h
8/9cHwM0eOdmKwPK6a+76kPBS7KcpFP7YcVvU3e5A9BH2xKFh/lKP8RfMmG/H5p3
KCsxw3YsGwrLwv3G1OO5r1Nv6lNfkGWbY6bQ20VDJ6MHiRpcBmJnZmuC14T+tpzr
cJPFwzmFOw45Vezvk1Cs+3zO03zzWOWWr8a44QF+Y9CGSkV1KqZaeS10upyMd8pU
i94hP2zG6j3kmYjIPrmEJtbQg4VY+EVJE/2ex6+RVW8zfY/9iH6nSh3vb4PSGV7e
aouql20p9zTu2Wp5zR8yXmmEQsE06Kyak41aMqdkk4v8nWG0AJYWdhOzLULnnrZQ
7ixOUHzeEvFq+GeriAhJsNcRI7zat5QOlYahq7Qib+IQxwE8tpT7fBspQdCReQ7i
tIuy6Yg8Oad5n5W2Xa/AOwsj7JnnhCFuFAdNyJ0Hvam1OR0Z08l+vzt+CbpvhTwh
NCz9VcOK1BR3Crfn3TOcfZTMEfLghfmJcDi+zIFKgX+Re6HpiCv2xwTz3hogHw4b
eXQl/19RI5LXh2h8+cXVWNpv8lDHjpTMrtszHqMmSeTvArSTF2mw+3aRDNV/PwO/
J6RX3UWF/7HnmOMBiDslz9+Ja/cboMlmIJk3Zi6GdgRLJf1uR7MxngPxe+ZXczge
0bYLA5XYIsaUfzNsgDhv5+AXrUR0MKyp+UZCrUhbBYdoPlwmUlugt4Y2AjZEAv0D
6L/ZEsvx5vNTnAnfsjZUs3o0E2FKZUc1OhOpE6duuYqfw2qYqk+CeT+hjpvF9eqq
KdVeRXO8/WQBoQWblazygvAQ+zFhDVue8fV6YiQ8ZIBAbFWu4XliuMay/SEXWdP9
FdI3akhRGCYiR9GpofmgIxX0aLsBtdnB1gEBwV87ko4UPQalMo4SOrcDpCGFrAu8
U5zHHylzbinZolWEJU4hXVlbpCH7Hl2YFcZF6lmOahSL/IIo0PhVqyJm7LMNcrdx
nO2BkCcdGEvkxiMZznuLyonz2BhJR/FRoqntN6z3uF3b/35Rj0RDrLIHm7ifRkKe
q4Hq8lt3qkaP0CkBvypTc5NPQtjvnm4IGGkEFHrDw5rcjQldTlDfropm9DROtHE1
PxcoPoSF7Ma9cIg4vcNhr84eyRZ6Vjp7nS2ky9sGORAYrb0TWm/afJi6Bi+Idj1v
IVJYpcIirGLUA0Xi8k2tSW9DZB4ivBRYnFpCbwGJkF75UNpNMsPBLMR49v3H1ug4
9WetTK1egocFgKjk4zH4CW7dIC3tMXCy6in/lgX2ZECXk9mbKbnHAcA2fttfe21o
4FrizT0XmnYDYV83/2ug5v9wIzoKrVUZQt8c4R4GjuEAR7qaaESBWrA4jxgmgJPW
wvMJe9TL+WmZeFf6bZF3AnMQxlKm3AmgP4h4m+kyTh/Sli5tyDfT7dXlGCkoPhJO
37PM1A/CiiR6Yu5ap6GUKvLPkm0padXX9iDUTW95EbSQdMPtssf6V1RvJ5Lv8ZnV
hTddYmPgLQCZEt4GymOuPqWyzsabSaWY+otvLTUuCyod0sv1KH+8xJrZxb3QsS57
cvE3vWtYfRCd6ACdAKIfNHxusWy8DfpWq9j51nKFYJu7meXpZ7BfarljwWAvA9Yy
7YhHxyt0gNlsmJCfBK6twkWVzFMKPYsBg956pfZP1gf7Jl3eaHE+klmSzZTNSNcY
+edFd95r8lWW/Tt7xpLlKpW0kEI7f8XjM7E4BEa8IW/19B7qvS0WOeX+QvkW8JKD
XVU13OnqnyFV12k90nbsW1azUZ69u2TtCjn8BQXg8mkWwRGHL8eZvrP4DpLTPw17
zXGjuz3dPmGXAX27dxGb1FAAFXlFat1rBk3/ne6wizZ6zxz1NVnKy17T3IWZxTHr
2R4h3Qm/VNr6Vt48PV5v84LFrTMEepYBLZMtZOc26ppqsWm2tXU/Gh5E+O5j8T0I
9F2tP0cQW6+u6OiUU6XGf6bE+AkRA6ZFn0dWWXx/WTJogVG7zb/bsW7qhg6h2HTP
rcjdVKl3euuRZlAyT7mEIxLFWKzR4qCSdapAa62SDxrKCFvYoCuhICYes1kS0L5c
vma7XGn41eWt/19iaUoTBqmT1v98NsL1yf2a5M1rZL2mwuoirCNEwkp07SzQ8BiV
c4YD+WOxEKFrnHyTmcExoYea/nvZW2qLMJ85aDkYEhJSIZ/Vn623baSiyZBVJqCr
FS13tTuxaKo7GiGBfUJm0TJFiLcsQmaVsrVatHPb0A5qm/+V7ZQ/STiwwc+g4M7i
mb4Og3TKWa60kNrXwX0bMsGwPojqCOtpuPniTCvU/KKAYOV932KL+Bo4+qZQeWn5
9NqLvzhwTAjZmsFJDvFnSIqDEAZZLkxeuJnpXj8sjdYWwLrsLqzs58A8gUvlLIfx
jVLs4nObUId6Iad0jiH19r5F/7sfTOsHbHknRhjy2kYZXfQYLuWWoKgEqcCTYCYk
NgyytEhT0PMktWqqWd7Gi8eKN1KKqrIXW7q1t12pkudgR51zZH5hsh1jaw4thQ3N
kne9gyYdSDFH9hcCt6snUYkyzQ/D5jCsWC+iAe8RwP8zPDtqDPZCdBPrvBMrZGTK
E139r1Z0Dcss5CXzgcAkp+t0/OjGDYd9MencwDfk7OwpA6SwBeLGEjv+bbOIVZu+
7+pNGAiBtnbwT4N6jeB22F9JgITfjDjcqXOtCJRi80vsJyexCi0fQETFLXNBsHNE
ElzWAzcEsroltxdD6g3HhAsCSZ4J8MGyg/p/FdNK++8iCo3nGTr3M7yhtYcYsuHs
ohl0y+c6D//ZvyozDM/HrWbqd3kSHOFg7KGNyd2u4pLgW2NFwYVaFH42q5VLibix
jncoilHmztb/bJKUerOqW45F8DG/eci0SS6NGlHWpeWQJwjfdyIkIsF/41UrcMCo
bGMzS3Jwx6dnNFpVejouHgmfo89XukZRYWKQv2pgn/FBbBTZOx5af0GjRnp8Pzkn
xVYk5xxl90bkPa5wKdDlPK8UReW1/oDptUgwWddsfYJOUN7mUyEcsRclsbk8nq4K
nF5XzbHeIyUvloBgylWo3zuuM98xmU3MrmWJPr311m9nEJLHsrrZKtiGAjsIY+06
akfQT3NDIRCQAFpRrtSqATaXaAlxvUSfnW2r1qotpSzGJK+5amUm/CY94+cjhIHI
2wz79Y91ppqNvZ8ZW/WWZLU8xO+sq1YiKlOt81gHY4Nq/C1EZanvw3ztOB9NmYL9
DYDat8CpczR3MG/btp7IvFYQsXAQucKe/BSzXnXHgc8if2uOyiPaZDZFsd4Dq05T
E2dqQLjc3KUurKC+g/s0gAGjjpQZpq1U+ampyGpHfcGWTEkaXQgoKrlFRPEj2EqQ
BLH/g/RkNLh5e4RVOWPKcM7Avt+TWs3K5vL7hBqScJ7/dBkEuEbo9XfjLWOnxLUg
zc/fQJkMdR1lI8lQwyPG3ZkmbP3S55UyddDQqVXJAeyWwhnSyQv27YP9FMAYG+up
vAqtJxA+0lm/acpcnjvZ9XujjQvICshE8NZjfsB+LNYxJl9AWx+0WhewiZXSx3VG
rl1OjKTvq9GLzCmmV3nGZo2GwviORUOG5cZC6X9eCmhLXzEWVKU+i8Pe0FYKV82O
wXkXxELtHewqFBcMHPdoJ7J8zxw17lo6OLNVjPACwbTi03e6qk/fStDVBc7WwVXr
0lf71wHUhfklrGYcQ//gKpQtrlY1KJjUPCMTLhKE8lQfY+kRBpxs6TXXKtpgdRDT
HZBbadsLDEb7gZWB7R8VgjkbxnGbIw2s4WtyeslWsIEW/Ef1NUekQgLKwEpk61VW
HI/Sbx7C3MLwZKsQZTLrxz9tyxfjHo+LBUj99u7GsIUR1EiW05gfvUa8sRV1uEeY
DTAKSIpTCrTNJQs74r0qd+pMGIk5cMBx0WjjLEdt+3sKFyax950Y/4P+zxdPL1/9
4lWgXtn/cZaExku3oiCfWiOZbu/DgJgl6I0Cw49v0rsipT0xNxCdtYAuBuEm/g7s
rZjRAAc+EZLlbIjwAb0bEAfZWr//RNxh0sXeABrQ0VkluA4I5QhOjsNqlkwwRYRV
dIIBFZAjecEudpSSMCQrhRGvk6bSTmp4RZZzOnuHWvguFFiBf2dZbbEfQQ5ZcQr+
CllDHziAd362mzB4TmCX5w0Xe+081eXJMmn0EkP7gwpl+JM81t6eU8H7oVqvvRvA
VGb276WJ6UuMz0mGTYjR8Fg3NYRY+QJGBjjM/YuXRdxNX9XKo18TO0zvKjwJ60YR
oU4EGLUiFuvVsC6yB2fNUte7yPw7k7504aCDvwtygCEqoK11WxzsI6sNDlAJqi8Y
EDJ1gD8JNl2D1nW0eV88rytR0YmkoAqWahGn8eKnaY9bH20RIfdIt77IB19GEmH8
83JEbTU9uc1ZcQfVp3U5vzPQeKfjGDqxVqzJMXIbqmmEGD4OCISnmRC9YCj7ajpW
mOpopsZ98TRn6AkGn0btR00xftFujJJUJMLNXwSrsI9VNNL8TQRn+jZYfVrrGoKm
XCsqpAkCcA532cIgfCEVerw5+zDhCx7j8qPgydKxzdggcUmm3HSNz45W9mBrmUtp
cITLTf2IpCl+sWp7wqImWllH+02D7rnSp5947jTbtmiSe62IXaGbJUtBf2PnzB7S
+xAB5GoT+a7zLzMnbPwh6Rjoaw7PocGLmtrPGx3MIaHwVH1q7RKFrO7nzFDivhyL
o0YcleyXMLg4hTAqZE08FZcEPoZmupYvy8lLV0WvFMYneS6CXmEl/0PHPKkCFBS5
cKPqC3CLYlA2SzTeMqKqU5uiUeAr9SI0w+m2QhUtNlh87P/RRDTPnQbcaWV5io+o
+NYv+jw4BwFfAVjdkNqYUuaO26g1Bv8QcEilWJZC4Fl3EOx5hzv0M6P5N3XoTe8G
Ojhfo2RZq4TX90yaGDjXkyx7DLvTQ8+CE4dAIg4W0fJez0ZgaNW3NbttAYzP5+g0
gFHcUsFXHVTw/TbqEV98JP1yGHx2jPkxZbhNRqTMK/OxV8fHbaZAiXihWcCvyjZW
mMD5YerBVJXVdbdCPqKAG0rql7ygzyvd5iagw/zM82FJT9OIZ+uA/nIINloUQ7eK
XLBGooGvzVNvWCdEOysdetiTPNB9wwLNMFMBjtsnvePzCaNAzTYMHMUX/l3HWVcV
9n8okq6mAUe58m9J8GwLmFAC/D8E4jVgyhRdOsRJZgQXzglzMcsAq2UV7sEvcuh1
V7QBCIGIqUE8ZQem2MLfHvquYPG3Nfmw1AVd7y3WMYo6NlMk709vqMUaYYcz/qyS
Hr+2Mh7yNdaDH95NB6g7B8l3zsy/WmFd7JNbbL5UUwmM5Xty4EtYGgT7Jnxk/lLZ
XLmcHnJEPeRTa9GQIjH8VQNViWPuP+ynlFTreKx7ICu85dIvNV73xd3DzClgrZ9w
+ts9Z6ut/J5lTy2qQ3dKU9AE0wn1DO+4HyXYeePCby4eLNmTwTOHvMZI4LCmHLra
S74lMbDXkPLecHgA9nPyBxzmMKCmcMHbaUuKj/WYR1nuyyRx0/Y41OCkmivjgQMO
JW4IDe7JgfOfaIMmlvlHvH5kARo82CLwLoqt03vy/Z+JIDQpvVT2t4q/fGlukF8r
oLZ5uK5AM/U5wHICOXz0ocmgp4KBB/MKFcqtmy2vyQIq+m/m8OhYNKOHsEMRdiKJ
BDdxGo5eHGFI5NPvRlFRERQnMlWMo1EMDBdquOH2oxJF/6rwze7S+jYkxWDKNe3G
9Tu/jaLrgF6hNBEwZs30zLJLtwAeynlqOdXSeCSWfRpqDa/UxOu/bCBS5JnT7eDB
MroK6FATMAjRg4OCTsFuu3oYEvg3GY7ZhV1mvUDNTazNEePoVX3ydhG+uEibTMRd
oy2Iek9SqzFkZ88orWW2m8t7hc5Zv0jA21gwylERxmXUDp/vj8q/AixBqRElMbKm
mqeiP5l4MaZtU//Ad9+zIM6KvRxE9fEqUGPnj+JYj/4lmDNxEWE8SUCV5gw/84go
5s2DwNoIs01cPRVQLBqCxa3AlhOdNLbntTgh64JGYZugCQS6nySw8cs7Jhcrj2zr
dYRAXAqKXcSHInODznUOz2m/zGA0+S+3NGp13/ujmobylM+wtomrEXWY1ldGWldM
bbaAIGpPrYrpK0JHLCq6IN072EUNw5MobBJsI7hj/DdtXoPAStfeMgfOytNgsU1H
Rek1IotTN5IvWuQZo0DfRvUrDteHtbkdTDbVfCuFZ3eZJLmKSXxT0OoQA1YzKMUQ
UY1p1hntaTYsI4XaRaK2/Hjs8rNtenGREM4WUzFg61ea8HwPyKrtNURXt4PsqWNZ
dI13eRC3DdDQDO8wuO0/UaqGKa/PaoZ4oaYY1vabqJ6/WxajtIvB8+pkJVYieS8J
eYwpQFnby6doMVUDTJT0CwzLyJEt3ryGhfBovTMvWvI71YG2hBHMDXfnYId6Bmbs
ZNmvud+VwITpO4aN4uXXxAAuAKZksmfBx0STA8u0DxuPyiJiB4/o/7tQvL3O2MMD
HuRyQmp15emFGT3I3/hkc0YtbPg9Nlb5/RWdUKSuI0mFXvxuLPgDBifTd6UBQHzp
Wug/B8i0tGBNAjAe7w/mEkEgCgTYAiE17KyWp8Nq2AkeGRLhQUIRdlsN2ezG5WGP
NGLYF3SOzxqP/ALrnaZ/iZEgPTfDtEleO08lD0eb+QI2UXkPg8QIz8tk5OBtLFse
HQNBQNN0Bmxdb5z2p25qxFyg2uWTniXAYBxgZ5Qcp3X3rF4dPxTRxCB6qcz8OGHg
HzR2qPrJxhfQ1SYP11PETppzrA+asW6PeZFVhS6B6m8CGiXpVdI/F8k0RAOrvQs0
hzJmxeg3jBEyMk8JXR7LlfQXH2+wxHxhQmnBuhThJ8y+nLqJeU362IhwMwW9M8qr
HwlBB4vKnPJtjhhxFMJwx3LsND2inIj8Uxi8IoC0s4H4MINucKdDllq+NIf630Gw
pzf1uCp9EnQG4C/BNGufbd9erOexVtETSZ9cG8S4PK82JdrNTjtkG2X7FsIOLvLO
8XJmr6Kbw2J9W5syBtaZ8HbiuKtCMPLNUrOmrsdOxwttg119nXW64c1bhtCByFhL
fjoYYT938Vis7jDdxQPUFHYC6+baYxQaTVJPbBulQ9tCMYS9eaUoHU3AC5xEG+cu
DUa67B/qZ5q8mtanu9Z1jru3mwAsebCkFtaAjbzYABE/kakti9Cwe+nt5qquyDRn
cipYZU5dFdequFaj+IAGEr6OFFPWtX4cByoxLyvC+c4UkNzek2b5yJub3ZFLuoSo
UzIeC5LfqzqAsgH7cfsQzAsDeSy/ZKc55JPbbT7Ro2wi67c/kGv9j6hg0h7N6mKB
rQs7fJdmQee82FugiMhGP5Zrdq+9mId3Ep0hcrrxRZG4/I/PvLCEIrYRQvqQo+39
xvG5mXmvPsenwBhXBwv7lnB32VOoIgjkFygeiKEjE72xv4/vOVBFRlzDb8YRCnGC
RlPz4tbCpfTVDUTxLxmQVSrEbVrNrcJdhUBxtilYJGIBjs8YULOOBAURQrQpNATm
yHwOPBWOHA9YZ9+gVBJSWollN+H0GY+XlZwtpxME1VDLxgEEBdvlANRipQkFYHf7
pDJea9SLRUu5ep+/fjQYYLIToLMtHX9TbcGVnilBd3CNd2nBsur3PvTzD0b6Bwtv
AN+cMcnb8eluKUaobdC518+Y1AiwaIRqXsfialnVULkiTfTqPR0bGnHSaulNUhOd
sz2v06rBvYLVgT9t4WR3CBYXbq/sT4UaYqn+1QMwqvUbpIuvwP2tsmEY/wHJ4wva
v0yHVc/WVxrkaRCqahBGbDFVg4T3tdQbfDMFmDA1SLRHs89rEqsEMXxShUcSj9gA
tHTJTooyNjTO2VrnmOjQvrcop6m/Myo/cwgf9fer1iMCVnlNaBn6eGh8jTbSn+og
aAXQSwhvXAXnkoZ5Vfi24XOU3SG672PBMealNbEUh3BCkClj969cW4vN+hcp2D4e
0Wqtf/p+5/rCawHJL1UuDcwJFxsY9sFs9dYzA2++OIbEFR7Oei16U0fxTwyD5VzT
Xy/Cnyb+uWOJ3+H+cNHtLv4UrYRM5MLl13TdIao6t3HOUE9awA7yL+GX208DCjly
x9ZvVLXgfXyzBkiJ6VIS1CCY+xiyOK/yeUYHeaT4rGNf33wsTlhizCG/YE3E8ThF
VlRIioCBVN6nZBpS57UDSzamUJg4BwvuAboEI+5EhW21jX+RSsESAgYXdA1VWw8+
cZesgdMi6kAV2k1SjQ446pNw+3W89+gQwLjTcAzJOVlSuemp9HtQfwhd2/xyCfJY
ZxT8pL1P4+rOyUDdRvVGmNHQJSCVa9PGJK434scWtJJ+gzEkyYBhDXoDpoyTSbPw
K9aik/faVsPQqi62A0NPsbPU4nGCE/xStaBj+XCGv7ZoIOhwKK2LFt6hoB8fFL/Q
II5gFijsKz9Z/v5GdpG+Afen0xePKGK5nexTFZi9aq9zF1crlSNQqW29Xftel+gW
rQ5YULdfq06oqn+A7dX0TGZTf0yVn1y6oJ0HwvVCiDXqnHpevcXp3/zbY2dp6vcG
FKpYYAhW6FsAXA7DaYdVNpUATeyG1cqY5SSLlxF2zXk3ZPThEE6/PvIaDGd6q2mU
DJdOAde2u368wb7+Hlwv1urMvBPPHQ4kc0ePV8ydlHqeJFrNAbqXXcRjyxTNwj+3
/+WQYz9gmgXtaHzzVJmCzaE4HDQkRP6vqremrK0yEc2OfP7P4iNd5zHjQ9zpySU8
pI3kOTcury9oBp2N1oQ8oGqvFBMWfItC+yD0DBWQQfycklU6iVU62yED8SE0OH0f
dqB2X75/o8ZZfi4wyHpn00PZxYegyxe28OTi2jXEH/9SekpXuA4X1N0JVbQxGIn0
QxiTIzEQdkMlyHdFbYFDjfJUPPA2x9JiaX8ynYUWlxTCX/Z9ur85nYNKC0ZDHgB2
GSi0OiOrTEGRxLHbd4Lr73ouW+qVTosVCHVXujcRW8dwebAqagZ2DjyEu46jn9EB
3j8GamrPoL0ZIAvddS1NiwquXfdI/my9GXUpqoedJsAZIwvyxh+54F8NLL0CXvAD
FadEaWc80YTHfMQHWMmMbt9ydlQTQe1ycw23LKQbrKz3m4IozJdEl6m9q01fHqEo
6ZLcpBgvEQb9xAd7QU03ROwoXDs6FA0gZZLhW+OnlAFqPs8gbmYgKGvvq5T2s2RC
tMuLc51SlJsR3jbvime0qL8LHQsETGkelGKOiM2Z29X7KWhvgEF4gv0C6j76vD/q
A9vBtFt9Pq5AjsQEw48ImtGHoQWi+Vx127PRhyw+BdlDZbiC/GjO+6wxLBjHq64P
/Om5CNF+WIY3o6t8BS3vy1Vw9E6kkhL+mrHIEkDLbhpgHd0Jd50cLnHFseYrBJm3
xJniAeMIjGOqHx6H8N3eToXUo16IdNXT1ZQAyHXoHk20Vmhn4FpzGka/vE7u0Kx/
rbZvOPhKFJVqayQjAtOB2FaW8jqVTMf0ImV8dYCQg1fNVQy44/iMRBSCMrpJeWBa
T1bNRQApn2Z2ykMInY5BNdfSqt2bW3V23X1K05hsqpCvCaI4YaFsoJJxzT8BPZle
/K0/NtboFR7WpxWnl3tNK6Ho+rxVn4+dkBTIN6Df1NxJqrF2dhHq6x1KkDeopHFr
2qoP4DS5G7ID9ETU+N272gWXu+fm/4cPMerBrW+yzQ3/fGirkBZj8dwU4vYIlny9
fuJbkvSKKrXIe3M8l1Jm6RgSgE3DR6+NPTiEL7C/ohPWgGAVXd0aWkALDh7k24fN
2FDmUSMk2kpXCkcX4pH95fhE8jQW5YOp3lAa/4UamBDfWjiGZcmkvAIqUTDEhZ9K
dEJJAxSU+gYmNtOeVxlC9t3tiaKPMHdhNDpWAhptBzOm1woYCTzFwqNQGdWRb56Y
+Mp1zr6G7HpMzNQOA9u7+nyQqngSFT4+WSqdlisoJPCNrYI3kOysJoPrfBTgNnNC
9rxX8hdU6A/PRRuLSQvg7DGXSvaUU5/G8yOckm2Pk4B0qyCFq/6DRFG317XtBrRW
VZZlfdJnwzf2F9kmqa981+kakaRqwBq7LE/Tsf9NFKBbbiwZdYryjOY23eGwGOLs
E8WoMo/uirGDMvkD+w/oKmwpGtkB80x3gvLqCah6ZLaagE1Ztb14MhOWe4i5xxzy
fpQGD5juSyNHXIbJ9cnrpwhvoJ+05yhEG6tV3aIWrpRNB1pz1sAm/WFNFf+Wr+eF
mwhxdWYHsvNgWIWLocnwafvlOL5gWbNIwSyJZZF+MgXIzomMGjiEw3yATjEqewu/
bO2PuhNGT6xhWZ8ui09lQR682OnDGC2XEzi2P/tJ8kUoH+Wb5nktDYEaJ3MM2zKu
mAKkWTYG2y6L2E7UC+w+YGtQtQVND54iJATmElCAiNHL7A3GHZYM2eSUr+nYSPBh
qQaphplTjREkoYXyWHfspMJpyuqE1Jdw7y1qUtxQYhiKB6XsbaA6AWfvP7ZnubmF
ZtuoG8TiM0mzYW5gwo9a+PtMWB+nYkrk8JqvVjJRHMc+SC5B9D9xZnTt8uBUyWfo
+P3FrJsAxgGf3SFJEM2NvWMybR/LWEvPLPMPLt5+Nh5dH5bAU5JbB15qb2bJKRcC
LOrz3H3knvQipY9KbsnMID8vbuFv98qMWckI8DPhzXj0qYOm9IDIMXfGBSKSPXG9
VVzgJpwA+Tsa7BvrhZVu7b3sUrQoO6vqnvyYT5Ht4/FCTR+iwQYouWY3dCpuUWj5
DKoxUGm/e7l8txvHFN5no0OYHYOc2lafteOHowfIVbkMDAJ/feOyGhkTNT1eOurF
fTS1JeKXVhLPDO6eR4nGldrNTLAlgSZu6XkfHu7KFkpDMc0hYj1d1pha/IP/cFMK
XcJ2F45dz4a+BF2Yjt+RmGCoLnK7thhXuzcqgyr/gEil3DPUE9ocXvGj/4NpOma6
JcJ9bLZggnUdDBwzUDYxOMmSHKu8Ci1iBtGFdqJ1Pf89ItgcNVlP7lVlRiBwQM6S
kmzgxmWzPcNbZm/i1Oeojd90oKLSnVK9i1CeU0B4QRzxHi1TyWXdqjSqWMIOYydu
JKWd2tZp4H9wVybi2eAX9wQWLS2yMxs8CdmsBTA8viw0TY3cFwry02BaQRXorogl
oogYNE9WNAAchFCP/HBGzyiBAwdjJF9WBM7X203ecNH8VDJNBBT0Ax9m9Ji+8fz+
i57GCSKmqQPzU203MyafvRnbzbte4cLIEEMYK3PNWSmrQUI//lnP8iUGmSqpXwY3
AT8PcMmOihuEYlI9IZW7pNd0F9hFYSECt49t/PDXOXnEWjJga/yPN+O0Tw3lSshd
w/OKO1osfQTd1wxH6D3dgP8Rmv+ev2G2uEYABmMFPssxD1niO6ecz1MA5jH2VUUF
/cdU9dPV+X2G+nu0SecJnGGcKVCD/pWLXYBONnS4eLeYfbq1Sa9j84yWhDLLdH0b
qmbjBBSReNhmuangIp70hl7kGJ1GFZkKMF50T9/K77Uk5JcaZGG1sauj53z3aKtE
pCPnMIRA1Z3LngQs6wr59ACku83vI6PPCA/htwN7z0TzzrrJ76AfyEka8pIQpbdX
7WjLLJFJ2R1xkosHROmJlslAWtLMyb1+lLiL5ujYKu5DQj3sDE96WZtc32VxrlQ4
u0H+NaWNHqIh/g03CUL/CF8ojJvOVDeR6UVIMiDksbwkIRoTvRE/PBiX1zwCDmvS
EX0umgeRTlkk+xabL7DRr18idpbJ4gX5vQwoAZnZITiCjGX6Yn1OBMJdp3OCk4Oi
OubynMsAy0HH12Z5smw9ZJjaArDeAwkmYm9adl8rX9+63OMUgPSkhbAmT25hJi2J
brUjCwMQomRp0+Uqm6U8L1s6fBC+XpB5G3ot7epmsf0GglTj2ufxq5w8zd2z4wSI
ZoTBQrAEpNTPKREZwQh4L7w/tn6eOhbPvjclgyhx5dP89g5mV6rhtTlbp2gXZqcm
de0O2tbzcAcvgP3W5ydNhirPHKA3eHESPy2lCYkpzOclPm4nRUvpxzESNT+ZGeWC
PfnD1s5KSzYZycXulPQR3iDGYHr/8G/gnx01hX6IozjBfXpdfytIryIsd9TRJfIP
N5TgdYzNfY1Li0k709TVGFsZyWk5KEJum900teHl3ccjtinFyrHEYxCucWp5u5lz
Hsl9NcKx59GqrupynxJ2WlhkWkcJ6sr5F8NwTLG+CGcERX0P2PKBF/gLHurPhWAI
To9AXjwh0itMbChrgmBYDaPVTKOhs7nC269c83KcJaZnlWYRVBJvf0Nwpwk6L6GN
QKzKU3aP4IhCbo63KZ7sySgCdmzx5f0lgEBFmQWfQAeGc6cP5nPCSNVMkoeVIZGn
rIqQOG3vKHGht9QIAGqal7tDJjzCkJLGhVCT+yYXytxSfde/xEJSaIlVoXlomFuO
G03Ntf6PbOFshLi5Y+Gn8Fyts2sEDia6+qJwTOxFKHXmXqb84inT5Ve3KdHqlK4B
Ybi6V7JCqFH61rQLK8/nRISo8K7BuA7rD5LxVEr4bNqDoomaV6fzakAEvS+R31H0
evRtxOvhmON5k8PUQOSABKCVvBLX5FtOb1T2brEHmRQQRERDFlOWkQvjuu3cPzPd
+DpKJeToU4itnJWiatjT52iKxmoHJLBMcYLt7jmWnNUaf3C/YAZWurtlJMjKX4Dp
alz4qZHoDAChnjGotpfkv2RV6ScnbiLq0lIZa80zez161QqmyZpqmtgSgsVwpKee
9Wte4zquRWLFM+EVz54qe9Ov/ahwkCDNa7ScZU3w/GsxfQE4sabSCBUktG0xjy6p
QEvEqRxZjTYKg0FDehRaHH8UViw8S6kyrT4rS32f1/l7J8OKAaCyvstqFH3IGrgh
Ug/Uqwt/8AX+QRWf2/7uc8erTRMh6Xw3MXHjHMNgveODRc85NGPvSGUADps37Eeg
fQ1URR5frOg60S/nOcvJv2KLM1xmo7bezxy+LNnD2G0KZQXG3FLJWb9fOqv2dokI
knIqaLWjlZCBgC0q1PH0TfgGohcdSAIGg70Hq5nzWDDit8zRG5/8mIhou5fMeGzo
21LzKp4+c5wj97puqrupHVGGqM4ckMy2Nt49CNXd4rh/Ie6ExD7F3JjUTmiM3/b0
IaUBC1b3NMawV/2eDZx29uFW0fE5rEghbam/nYkhdW3NOLql1JltEnN4B2hcQHze
TTocmR2LD4Zg/xtTtbWG4h04oFo6nwlnD8+WRsvItLa7uGqAVrj5uy+tdcETVKhd
2SvD4OXkX1PwguXzput5849B+UbxYeAj/9y4ApbD8W4MZn2Ug/nEhVf46xXs0DqX
xtMS/3p3NW6gnCS7QxhtPxAY5+u4m5ORxxGE7/qVx6mq/M2f+YvF/phO8eJnBATQ
lHPL+IKDZmHZb6K/YucgIK5mzrtZpDvOnBIx6zsDOGwqzLd5ZiblWy9IGRWFprxo
oybVfvBGC6c9b6L5ugOouubB6JxO1dAPJmg8N4FQ7KflKDNkG7G5F2Iyhpq5vmHt
9SQtf8V4ZY30i/uMYQVlTn+1cw6x1T1f4WiG0crm3dqFIw/LO1A41DhQKoAqTzSy
opylk01f8oUrBWWbm36gjpe3l5XdteT24mYgRG/k3rc34WryedCcI/NYYu8rErr8
I2gdTvVDfADKijplrbTEdyUlnBUj/o4vcjxcsbdEAM1VukTOxQlghl15zQMWf7XC
QbqBzzYse9WZky+LvBAIfTT7ESux48nbT0fUC6FJ07UUaksYiAfuvHv7DgVIw0Wr
RPNLpr5ba91MmyYae8WQde5FHOw84726bRFrFMEJhTPsV90AoNkW9tJrwTqdPf+R
ab64IYXpa0DI0DrIvr3wlnkF395k5nSTuZauftX4x5Zd15iK1aTXmw6SdURtLCi6
Q/M0nAcRLpqUtr1djh5LGpzQ8Zaumj+HpQVRvwjSvxw8NumY5CGXCmYYaaJdRwOi
oZwJ/gcif9xrd6L8YQ6x+UJdT4CLGy1Ttuep5PEBEw02tVLJlYvmzA1oVDuQu7fh
Z1ahrLkEmC3B4UAUS3CpDc25a4IaWbnD2SHmFDv1hf0ZtM1GD0pAalGrcJ8y1mtu
XODnz0yKHnQIXuR3TAuL2HODpqv6v/trA2J4g45D6G+vCoaL8PpgPkp2uzKLn9I0
pTXmRi1wZd8SX1/h7NNYNTTRPfDQ1fADqY87jL5MR5ErB+tSXwxqLT3C5sxV7mu6
gqTNMu5s1WvRJA6ffINANJddwT6qSWwN5OIgmaqUwS6SJA30cvmcMPuOHyohW24O
Nwe54GkeRwDjZWzf9UygkxMbGXF7xEeLW+MBODuKtKlC2c6HIDA6Lc1MUD0ZCxVs
z1L64qHfaJMX5eMmPvuQt4Jw0pPjp9xsj3zUtp2iFf6tonW65twcNilpIFEWDDkH
gXSbEujpf97mr78X8+VyRZy+Gg+pKp9kX6IgdHR5NoJUIPjFF9smODmziuRJY0tM
YJl3Y3agLa2OSgKjXfNqtNF1rLFdwBSyJjq1D2/FlSWrPc7WWjqtFe/L6tr85fA3
J8rrVutXfcz7uVUOUYREeEo+9wk3IocxgWb+eufPdIW+LjrB+PxYdlIx1k8ABxZ3
5vEVfdhX44LanUqPeQ9aHpRHnbjmSdvtHCb9yqhA8XIZZJqc91lesqMf5Gbu5dpx
WQazVDzmwCQxW6NXqIr8EjbxDhLW7JHih6QywAiUVbvmzJqHbpnEKcwuk879K98s
KAQwZBxxPNjVpraQ61su3JOdUSvZd3YCi/YNcta429OLca3RTwYPUMnXSkn+TVr3
sMaQeIImY9QPFJuRjEdF4G1beJwIlQJXg8CD92P7lrV1UriLLlcScmOTLmqQDTvB
BLpVlYQCOtng1icqzplZaGHLo8fv02+vMktyotDKjjlUOMm+/V1B5+PXCfyHrt1p
fBj+zEVnobHIzIw/4wf2vwvBt6wuMmGJhu5FLx/yGoFUVCSqXLgA0samRoiJlf6U
EJu8z3Tq8Kfa5+VS1A8yegPIRtGjT0Oa20C2hj4eAqljVM420omNu1QPWTCyKHNd
+Ys/JjGYlb6SDIVRhrbMmh+2aeTtriCcc3hr+QN1wruU+UUwynBL+DnASQd2iAwQ
aOxRmr1FZMFDMPvzAxxodqHnSjtdXCDoZwuMq1YbQrjq/HPbfMZnePniSTqcteCP
Fx029Oj3yWQ1Gl2sTdZz7fTqGWClzHnzQvj3MQexSdGGpaxY7RDjNdLEmTLPFvi5
NA8UF8f9KUkAqDBjuqBIR6N0fqbzuWD4MH7XaPOL150nnbEBqlNbbPy6hj5hTvns
5NMK5V9ygdwUBUuDPnKr2LdeTGAep1aJ6gbQOkKDLPw0x/jX42q8vCTEMhGwmesp
aRrgimTZ+o9DHxstlHCkP44KT2+VUfPrnkF/vV8/RfYlJmACBHxjlVct+uWBqZfL
xDLejB5PkoFaCXqsTb1HGWBUEpiOY7z7axbtltUhNKGqKpQHIczz2vwmmdklH0aG
Pyai0heuT/cMxqIZJW+IPuQxSLUYUYup47XKv8zXWgAEaYPBUCOdJayE/onx4NF4
eQwcsiQF/OdqvelUeiULzSIqAWYA1RQ6wnKObiZhbvzMVI/110euHRiH5/NCE8KW
WTwGAnNbsbKoTUPy9duE2aBOk8KB++YQrdz92lwOE+u00qDp1ex9Lmiq2OpepoQR
Ar/h2ZrJyh7bPqt3dI2TC3Y+p/OVepSQa59ep/lRse6llIY4LapgnV10jQ6oaaQY
iQRw5Z7ASWSqpI2ergsVL1o5zbYC2VJ9iLA3dWi0sThqwneV99V8D6t7YXfokXc+
I89CODEZmTsv7FAa4+1MAxzJ/oNcTGgYUHBzPExvCGtyX+ikcfbBihQmWbyAfO1H
RSaCIWDegcRxv9e3TwqeOL7wPfsjNQUgWgrTGniOeOW2kkjSx+KdWHkMET6579kR
3CRSDV0V0D4mn8aTjPApzR6QYsDtcC+0OtqtKbPgI9gS/5EHxXic5O2nf+ZKJQ98
atBhODobCvmsX9MMYXYz09ANNeATYnVN7iue0geoqkFpEntAqvWqzk+qgA6ElN5K
nt2wIIYpy13lkTdoJg0J3MU4na93v/KGr5sSzifVCfucPl6t1ftFdH0cCdJ0EtR9
uAd/9qBb6SA4B8C13YTNNjZS36UjxVfzZA9QrocGQOHHJL+geYa+g0497jjjWwlb
o0Om5iy75TM0Ta6wI/FYa3Z8NWv7DPW9phxc6dvLD+vokjXwpQiE6twuMTk8Ic1N
nSio611lO2zcNPsYiH2M37yaFrjLnmfDOKh0esjjc0oleGXyHRZ1fZcMQSpYsWrO
r8Hj1TaPrmWjuPyrhM+UGz9DJBtoIF5zW+97xGP5WzzYSRjgChkzj5qZHmB4SOsZ
GHMjo/VNPsfGCYrZqQoIf6SqGgpVjxzNHhQEFFaVmT/GpJiCQzvTf3C8wgdJ1Fs2
zCb1RDGWZ2cG6T+fEC9mfxpeq6RwtNhhdPwz4DlpoNaSd6P9neGG8Kmyp93JYvpx
vlKkfhCtmmv1bHZSxOHkeOTKhu3BqLtPnBnUEmmEutitlNr4l1c/BIUzuq1lAQAy
LwHYzmn1fzCj/Wgv3aDo/GBNjaF/ZdlSAOmsy6vmBXo4Slnzo0pc/Hk8wgV/X8AL
Xlzwca5TO2AnLCgg02LYafURZfHwvvrb7VD3jCjvFia8BCCSxBn8pvE/FHKUyL1/
gLlxb6pef5bjICZGBnFnFiE8/eclUICbiy51+PDUMtcbDMCbaGLsVlx49zFpiVvh
EFNUmngPpw/T0kRj9z/9uRaC6rh7SrCVO7AAfthQUIppXEPmAwOWzs03zaE4cjq/
+gPXqj4ul9GMbclGZM8RSLz1Fl5LaZz1d5opIE/J2Sisnk1KMFAQDvBtORt4DfRe
UguLDEUpHk4sypPVaG3JrxSRhxiIFuntEU/rI+qPrgowZMlQKJBk6l8AXq/gQ3Qb
tMbBBNwDYiKW4Bh53gy4rqXc4WEC3oTszytTmiJJc00RBdXd9pqSMues4m4YlW6T
SNowSkCMcVefMf8NB4DmFgTdzSNgWB3sffrpGJS5xenFDrYUzHDNIjb7YPgxFY/i
2tqtXWK05doeb53pk68Nb6nNLH3gF/wbEfkCJDhm97Lc1f03M2FJ35LPclNhLVAv
xAx1qDbTH8Qr8JrKa7BwUQLIc7DDYE1xDu5w9+tB2TPY0K0l8YyIzsLwQPIbBTwW
EANZy4APP66uJAyMJHvSzfq1eAlUAxXGDdGDtN1eURXpHz++0rjPasOv1IfN0Zjp
KoZdQeKTHgzHCoWV8shCt5RMKwb5RVc92Q3D7Pjzus9T8Tzsf0uCT0nGCRh9J14r
JCOniEF0yfLP5oB+v6yeXsPlfYTQGnRgHketc09INyy9lilI7Ms9NwIEXzcGaoac
BxkwNy360kdePZ7xdmfrSLi3F6avM1RNltdopRWt/NuyOquiHkmUygh+j0LcF7LR
GlTNrDQYTdQzlISZFf5Ta3xMfj1gzMstxMn8SOjTj3pdwyq0Y/S6Is1jZp+LHoV9
o2FwkVH+0AajF+N8FKI+gdcSzwVjflg9ayxVRX0aOug48U5UMhPoZhw2UsvwYKBv
IQ7KDfE1an1eB5xPIIWdtik793U4scOKZyFMhb7MDEG30Rmwjh5TG8snDwRFDzyJ
UwM1qiNpxhMP55r/X5Cx7KKORhJFHqFP2huuWqbTMlNuijmrAhd1qtdL7AUMMcdp
nm+wiTjr8TQDSr7042tCR8nlu7k773dwV4s93f1S175ObI73Hfg2McigMBbOG51t
vY7p0s5HRTvMMsqpCQSpaLiYR5ItxqLxNnmqlQLo9vCRPHHEFCoBoa3E88OW9k6f
Sw7SpYW0FyzyEqIsXMkxN0YQmkpb6WZtTL6PxQo4zyqc8OX837lBlCosLMirHJye
9cmEGOpmDRBp6m5sI9C86doNCB8E3KhJ/PAVwkddA2mYE91mtqD3/WeH+wYfp8ZD
Ux7d5rjYi6qYOl68VbL8hoGeudwsghU5ART1AFfWs6b/9UCFaKLAhd1m0U2dfGwb
82nX+dqu0cHs8iotlp9YCfGhrHnOg5zjabvxYoLyDhqY1uo2w+8sUqCkJcY7/8D5
ZKatZlPe1LIa6YUc+KBJQiN7unicwNBTo1vq6rmKvGhPo9Orl2wJuNm/GrDm8zF6
0XStVBD+OKbZ927lT5QHc2FEbKQUIlnJY3mqhBQZAQuoWgdj/RUPG+ZcfFK0T3n4
djxPtt1aMTsbSDSprqect73Mm4zj0ecbsGh69CUluKX0L0IC+Sy4yTEkhluKzGIN
zk829enmroU08pzQEP2H33n1YcWIIy9f06MP4b4X53N6qTcDCyeAdtfszS2ktssD
2R32OUxRA1baEtV/lZQYj6Uy6JK0p6YoMBrdy+YCrKvUEi+P4BVgL6OeIk5VW/jL
e4lTrIEQCFmqOHTnGassrBiG1ChSZD0OZHJ711ejFl2/5vwPiTtoWvAbtYB9HI8i
AJcnbYkwAzpQKMuyXkoyiUrpR+d4Him3EbZ2SFkbFbm72/yqRG6nclS+jfyZTS7A
KVvL8paiKwaDtdSl+bC5kSOYsgEg+FgcQYVK8rkrGqZg3yh15XigOzo2LSwPHMPS
iCwQJxf/Oy7KLqU2UVV9rvif8bP0N9ILn4xsahloJvaGTRFlE1PdmKS3iyb6zoGk
5aHpfml9koKe6mGFFHKXLZQ3vYHgxpZjqbcYRUp9yXRUlAWEXHGuJyuOwgiP9Ske
o5XPW+8ksBHn6h/QSQZTmUh+FuzhBgTpEVzO8fCVNqW8V7Z4tKIbtP/Z10RMeJrZ
8KSu2VxCPvXvp2WrSLVfw/EjRnM6XmxKbGhQhlg7VKzkoVAKyXIkCqOrG5uxkLc0
NPaOdUurUV7N3cxX0TTrSBekmk67oeB5XXAqs0UOFG/RAEmKNDD2G30S6crRibHX
j0QokaspL46FIkDJYiiVnTBonUQUMc/SF1zjX+UzlGBizitv1pTO9qoczdtt6phs
MBCc54T9ubSceOvgT/1A/DDvFNUHVMI8ZU/R6KcqGG8LuX2o9Fp9nlQJkbxF+ec0
6ZXl82BO5hQI0RKrjRrZcspuhG0altdui2TCrIRk65YG2F8q3tLOLglxPMaCrE0Q
aNUtKN6PFPjGi0oqPsQnE2gRjy7KQwcWu61OWtzBmVqd7u1eJXnMrbw0qGPrN2J9
ilkbpF5wPTEdXr3AvveI05hcMt7LNW53DWJRhCDgVyk4LhIItG4/u/ffQFv42tWD
IN73X+ib4qut90B+EG42woDBMyHMAaV3li5WQk+pxBOqCbUiSKWHvtc3+YX6ARIw
sg2ao9I/+huUdsj+c+irN1YWwHqKVs/vX6IK1NFhFimpasdmQE4u23ddy469Bkwu
hwYTow1q06pGwmHLsK4vs9gWpm7cm+2thNa/YHn8peu7+eb0sOQ6UniLoP1Q2Ohx
ukxEsvEtmhGyt+PiajwBHYyG5uDxyZO1NbaBHi0XV+ammwMnt/Dlz0eGM8sOVcYS
I+HFwkF6F8DBc6dnCKUGvsn5pF58RkJZv0C3fOrdO9eB1gzGdPXj6vtir2x0JZDe
/RttLnzmF0xcrT/99uRnItdh3HQao3Ychjzf53RCYMKyE+Vw/d6Y+yDnAgtl3KgC
aM9LI6Zs+sosGp3Z/mcPpGxoYcP8r4S3kxSDAUmY+2QRJrj0Tsw5NegD3oq1l3mz
5UlwjgZ+/iHgT/5XvMdK2+h+Dme50Qge8iN2FgZ883U1WTp1Uz2eEy7904pUL86z
m4yxhly/4+IoBJ0a8V79f5dDd5LYc0Bf7tFlmJGgQXfE3EzDdV7DVAJOzf5xQMcs
fsYjcYeHuO6EeNLS0pfX+5Q/WAl/vpwfM+Y6mvbUez/sjUqUrW70YGuPHcI8RKTP
T9NsQVxS8oOkR4UqjgQ8HMTHidxA+2l1QzhbEEHSnxFb8YY89+S/XjxSXW3NKmYl
i27cY2JDuYT5TMDm460OlXXnSbY6R/7K6iTzjRAH3i5LVFw7galxsNUj/u6daeiT
IMDfh+ZnUZ+iyd8KRZdPGVVD1FpAYGy9VpcUxoyfWMD8DvYdk7Zl2+V6ktvY3qRJ
42HdPLTj/iyBhsUnnQgkiYcLPHGDYo1v4ik9z4ke4EKLgEyCBHMyKX3zRzgCM6eW
HXNJfcwP95wEQgj00VrNyRfm4Dgljyk/h1FxbT91Mnhn+BucbQCKCEx2ORRwBxZ2
xn7QGdzBTGN9onLzKn0L/bc/IiFXCbPkEnM18tQmIhmAFrGop2FD0Bu4iNx/mdsH
7OY9QhNZ91bQfR6B0tIZVtO0gMpcj7O4utxafDYioQjjAZmjWD0WdOe6eGqLzaM7
w8eELYkMfezvyyTHSc6BapjRDEZr8F+eqOKByX4EJfLJHGEpaLIgXQUI8HeDujPC
YiJ98B9ZlnLv2oVYOFosBP+9vAcufS1ReB0DEfIMemjHwlES0po3qfCEbS7rf97j
LPmCXwQZc4eLm1T8RWkiKHML1/fYBNcA6hhzSzCezkW1n91eIQ1KY16nnQmPkIxp
XhkVRFLzauekHoJUZ27mgKzKxHzjPJf7JROuZIZgU2elNtVBxEXTUay79M/6OM4j
ijY29+o4OATExWRx7yGpHY4gWy4spsZJwcKlwVoBJDhsrBWLeud34hyI2cV1+Qdy
Lna5URzxGRDq1ryeOR3u7TBJoCi0R92gzrnzhnY+9a46mUZxtpH/kkoTwjE3YzR/
5AVBLHZKIqMVFlOg/buQWC77Qsj8RrzL41iZOJH579zPjdH3MsrNL8ihD0hm/b6l
RVRFRTLqoP2Jbs9pk5ActZgGWWSgF+O/JJB925WgaLy5WjQrqYKy+NV6IR1vH5b0
p7ZjDInj7XOAd1zNSmgYwig6nUxYCT2ZCjdMXWNRdhbq5aXy8zz0DwZQxQfQfxa7
mp+7XyxB+oyh1AILEIAtS1J01mLH4dgOrisTrIOkoxRGL8J/26cN5mv58+ezkddn
tbZoazn6hOGegMp9h9KAEo8rftzmLoLhld0M9G1tTwxn4M5aUgtcQrXScL9Ygf3h
mTFztkEBdC/BOeH10EcUW589ZNAwQW82xR8fj0ULKPlbXOv6cpco3beC3jMAztLP
GG7joMnwxjRFFNGokL4kEaueBlHCzR/DDfU1Wp4x8Z0rvu68DgNrIGgjiVQ08xjT
2KKVpAJH3oSOhhiPnKX8uTPDrCRnCNNsp3d7KWnQiT01qDYnFtvzGS5Yd2qKQvD1
fl+GpikDRIKq2FAWIxVQUUhXPGdqBAir9u+sW2fYu1TjzLDdqNNi2PcluV1MTup0
nLQkgX03qAoT2bJwr8fhtiBTATyOfsxd0tAEyuhPWgpbsf4U2gq5yc0eZi9FfBpf
UkizaRFYw4+PNuIhdi6aheEHu2OEHd7mI6++N3Ncr+7rtMP0HLSK82QxDQODTZk3
+S/xFemVWRSEOc4EJfeF/ieAptC5hUXZ98GtpGy3qCCgp82p+FiLgtsycSWbsBRo
3qZUPllAaAMPfxnM4UY3JEm/j984jKG7FFZbGCgc1lEaHWICazWmIFoch4LTX6Om
pmHzyVf0F97ihEAaCxWoDfKCI0FGCwN+FU5kccDy5EtgLDHJPNlCfglZliAF5dlm
JPm6IzKgDlK0XGOiQ1fYR2EUoLvmGrDQ2MbDVziTFoN/RRQGnIqQ9soZUOWOWWOu
Cce/52JWsYnzDD4yCunyEz2qqsxaYd0J5WT5LyTO5SUG8SaKPMUeVJpnl1q5kdoW
3Ak6lS4F4KII6fsSU7DRHfykuNAYhvDTDTs9iZqyJ8tUbHrVMU24QtkDkCIgr2dc
IccBk0C8fx0cJWzBu8DoBIL6L0O5VuzsIIuTbrP6hv0a6jH0YqRv+oXbDliuQQfO
pUbAT5HufZDKEe6ySCK1ruMY9YT6qoxgaMFpztXPaMTIAGOsR19nrJwEllvJlSoz
5aG7QvBW3hGAeKdUIDc6lwutyuTKbFNzLMIT1wkQNMUhrdWfyYlNETgkAGsO7HGs
5LAHp5CatOffyQthmwTZv9oaVFRP97ESW/Da9odeWjlmqu3rMy7DQpOlr2xr1wKz
QoBS9u2bNyQ/RbDy3y3D0MPtapcsaksCyZZ1/VV0kUH2nbahvj054Ys/oul97ttm
kWUpWwdNXhpczVrKEFPFPs0l1NRgoBuC2iLxNyAAO1qCOBQOTX9GwUFeo3sgnC2t
XC2dogBfYpTtnCwA0bD6IPaK996IV/1Yo2E4maQYSmF5bx9ZnJV1iJuJGunMsNFv
f817AFtBrF3Po+OOaQuSVagnTSy54lN4InA2StgGecNdNsbFE9NNlCDVuFD6G534
cbbu/vBNgPYVkzNMU4pmz/+R7MGMGBt73npwhSyitKLrlVxcvzVu0M9dM8Ey0dx8
+x/hoKAeb814Jcz+lx3zfQn46DBpiIsy3lKhylj+HvIzLL8FJLsLSuqnB+0yA4dW
IWnIydlLFxSa6jS5henano3LLFHGgL4fj75rn1AH/4gudwrsdb6k/iJ2U99Gydjz
f+6hrNSMppTUdqyBzrt0KmzQ0z7hf80zB6pmS+aE+pyTzJs0AjtWGwpTV2lCHDjB
r/JSMr0mHXhWKLDvqGNKdEBI8cM+FaSUa5fCYoZU0Z9Vht56OeJIcUMSdncYfnSH
b7FGKnCmT8kquMNd9AeQfyuEQRVGtrg6FqR/VLcr2IVUc1ulOzNZP6STtUl9xjyb
QygqeGJ/TbWcL5M6JjH30hQq49LhJGBhhJooIGfZDN5QiHvjiPcSBpA5u2gReqk7
UfRAVVk7AbiL5WpbFlfFiLS/qbzUwLyEvXz2jw+1lYFYnh08VyGPqyrkuajRr/WH
4sZrm9KN3syqyZyYkLuLgaUuw+K4b748QFiqR4reS4ELGh/ChGqmsUSwv+GLqfc9
h7ie0Mmn41DiQL1T0B8UO39rSUqasM2BOx8mG+4mGOyebmEjt8NgD8k18JgBHIVh
RcldWWHQJZeMsDIfDrC+ZvU3bmsGiOXuTd/yUazDtDG8AeOegIlt+FA2o/OHrTci
jAqJLrmLtdU4F9cmzKFSvfLTf6HyjN/vSP+XqENO8RWw3c1ZlMHdl+9o6OR5sS4X
IAFpyxbVoBKZUZhF1NEVBseZte3UTF5wFNFh5EiW1pnsnuUhGnewwCJzTgkcdZEz
x5q5zkkV53Sg27C1N36EGRZkNyuV7efc2YdDz3GnsVrxUF4hLzD8jocBc2YHl9/A
I665VV/9AdTAuKUo+usQiGYDOHLQ1JM+uGaDRePuAJEq8q0G0skOKkkmVD2PNyxJ
maCPrU/bZoEIEhApwrIfLZtEZuwevrxVjSvfFVYewI28VC4TpSHgRvCz+/8zVy29
b6h5t4G81vaDS2lmQR9U/VUNF4Grv6fIk4IEZ5IfWO08c4nnRHy8hYhuTZ3ixl/E
r/vTYzhN7lBT2dsQUrpSsxtfFWTxjdALWI8LyrKvzU2zCXxOWX0TiFwRgjzDWem8
C2KNW8/YnoAcgP+jgN7Y1C++tWmAzCQLMon/XPZNfPZNpjQ5PZWrONlnKivODHwd
yTIZTtq7pB1TyRC5t0D1/pDDUcxa+dMCVsVX5rYd7yuOPhI2kRbKUJx+yuAo8Bhc
vqngXO0tna3mxXiSENjyj+7DrVJVgKlkY9Afq/RucvbSNhv76EqBpwfhFxAkkdsK
TFRDHH4lU+np+PFDNFus6N8q451H8Q3kytz1v1+5KNxwASPOmc6w6+MOZhvsYNcA
aahmj3NgA4HJqct1JnjMfdsLfNbp8XOcN1BSNVfwk4M7stMMqverOMs5B3NwgUkh
SJtm64vtrn8RpQaCrS0P3u4PtdCIoL7vyzPYemgT51WjjP4wwB4tpEUnCXDq31l4
FqOt+vdJkkvlcY1Gnw3XI6bHq1wWPttj/qkPYqrvEDqQk3pZUAXdEQZYjXwBoKad
lvjgzDZRPBALzJLUARNA35k/jqtC3KVL3kKQZkm7gdgYdaALcajRO65Jev3W4WsO
vZjc4kYbDmP//SuoI2s3SWUik8tMSfwT9epJkZLciTLHvslfuewywkBjVr72sF6G
/8t7ifHJ2Mz23fRaIqMuHEZuMuamC3oSO6JFt+uvOLwCFiiBw9wVInrl4wbMl9RB
7mkaM9D6+57dyBzsmX4qt4gn9IwJLi+a4sV5rhRbQScP/NNhBBj2ieDoQPLCxm4h
Xdw1gBgdYGoPOA/PMJ0QnezCBZ8VlGhbBLX3PttFqg76sy2H//W7zkXsjkoLUyDz
7dLh7PZeLQRh+N7YDoR96R0RLr5KAROllIn4If+U1YzvxUH1MUKAl6GGQBaCenVM
azXq49WE7vmmgrdb1sIA8GkjmePM+F+MdnG9xD4Vkv/8zjeAl38ekhoXBqKcH+UG
qGm0Qyh8YihXc7gOcMks5SkegASy27nEBYsHRflY+UAyhfY6eSZkwwOssUkUOLcS
W64S+d3Or5t9eRar6xu/2Hh8AOhGTiJD4LY5dXGMBUwBU092izVnYLpZyBkZXdLG
vxulDuY9Z64fjfM0BMG767jKc88qNeiZ6UMn/D9aCYAI97HxhdkMuxhgfsp5HRuz
OxOSBERNJ/ORNM7rmE3iBLg9Q9VJ74mciukFezcehKXzWM3LgKbusFVcc1ZlSLRm
EtyFR4YpfRQkn5daAy0wSaR3fCrRGSk72elReJyxN7rqVsxTw3ZBT2QvO+urqXrY
bmWSitGJlitxaheAQa9ojOTHpnQQ/yun+eCAN4NjRtpbcYwBDIPD2SM9PZ0rUehV
aj1Jskk6OlQBq4yav0MFT30MD9e/Sh+oECu/hugoUAieUHqmm+hMM3WSsM8suHT6
cgsRx3gt68TxzqDEpBggE3Jc7/k0V9xhHLhETDf2aJ9+UE2VVSQGamY7fQkpK6Km
/5Z5hp1SOHJKXhyAhCSqF84WcUpNUZL0uK5I5KBYqU6woWcD1y3gPaplY1LGnCgn
65sOlC+0XqPQCdNbhoCOy+xjrsSfkuRQDBGbM8Ut3gpvR2fMJZaGU7JKMHnYPdG2
Ielfjt7AiJ5VSAWIzFGn0jSCqz/jDooeya9UOuQ8TP9JDNrU5FkmiQUmT5RhL4QR
QTaUXbKi8kS2Z+vMpg/BaB81p+8sDFZm7NcnTWExLqZ9lS4ttSP49X7+ailpvflJ
sCtxnTHxQbp0+DPFeUcA25ZOEGg4EzsoM58ohFAa0GCP9d/4R8VyAaM3kQBZkUKM
kd61o2yg3z9DOIWRX5wHN3bDuwoHxGl7tvlq8o55eTnI1pplZN2kJ+Uicv6BLvh8
VGX4fggG9Hp3Q1qpygf0PMzARzQuhovMLomA9STNhR6UdjKOyAWjkmynqncxZ1o3
rDTZj17AFTq1dn1TL7fAHf7rVyDZKT1hwUoKmc4tR6+INV7ZK6sfsbJ0bajojJAt
OgoBuJkr1NJfNCHe5L3LNsrj8MFYiwxpiMJxZuFCnLNEo7Xyoanux1hyVCpy9ZUG
c/9rFCZJ4Jz0I3G68IujH7MYgrMqXdsofoCy2YSHK0mCGKlIxYMabjn6WL1miXr1
Ut784lKJdwPGpeNVY8zfG1aL1pQPUIw0A+o1IedsTYM1conUSyrtuY1LNwUD9uHu
wOHmecsx2ypXg94lrRkHGfTg+FBiFapV8g5AwZNgoY1pKFKhPysD2AZ6BCI/HFDH
/AneRZl2nV8fFQPtjSRGYdr9qgOWQOLoxiY0zI/n4aabipKf4zY6A3528OI6KjIq
yBeN1LBxH5YDslFiQRJOb/kPrLWEYwwGQIKIHsnWc7pVOWBhxAyAnrLR69p3zXP6
EgWoeYCHgX1Z23HVJP9dj+GNk+tAP/0HYm0WlvHBudpXXEwX2g5lDrAKaezOHTRz
5sQjuNaUqV3Wk5dcEloyy90Si9PYC87R93oGCVcFQyTEh9C3AxNokywwgUaiixf+
HV63TxjfXO9L2EeMTFXr/aQOKoJTsn9q+TPzLtPYqcHJDAqIBaBk943qwtBgfLlP
psK4g8l4fMaE5aJIolxNqiMpAyV8s31efYqSo16ewxxR02uA5IvJ4K4dRs+4ISro
c4vo9Q46vRfi3zNBKqO9/Z38SrwMAxKA09MzXw41jo09wTixjlqam5UNVTbLVTZI
19aJkC7eozUPE/z0bqRrlJ3p41G/i6GdcYuRd/HsxJT8yvOD/E4AES7u4bDAqT8h
5y9pZIULZbprM26+qBQcDsyzmFRXrI+KCLn86dLmEuaiVX3h/y+G0m+v9Y2YqvD9
ZZxVj3n8rhOVLU0ZIaBwTjnCmr7HEB8giuFuCiRXEPyjzwWHAIgEqxPShSa0+ObV
zBMZGxk7wDMEl7BeljEE2fkpe1HB1h9F6N0ooviBgnP8bxJ6/P6gnMGBIIyUj9Z/
GHJcV8WvcvUW2FT5Fpl/FEu5PgncgcadnJtQTxQ8aJF37ylDUaQyRwvRwe7y9UJr
I5bElAPMl7wdwYj3OzU0pLLLkY/WubC/J1w57FkLb7CAU+MzOv1mW0yTDep3uayz
RMxtLQ8x5Eh8LKp2Ain/HTgGGw7kjgSE2amcdMMIs16bn2LukSci2efr/xGWXdZ4
l7Jxk4J7EvlCI1c56G7pw51poUDYpJglM4axwLZ8b+wUK4Q7ytAd8IymKRc77+hA
9Fo2ymdCQ8ZXZ30lkA1Pqqr+RSe/SLytChvHuBklMWRxuSeHrKiVU1V8V48nGzFJ
9PfK6o8GIW/6XJbmNr24t3aS4AJEos3reLhpNOKrkps0HKI34YZ5IGaJkLMVQgOZ
U+iAe5m04G0+M+3GQqHRUrxw26YnSaDespdWBjMsWIltaSSCRLDXaSSVfXumrFPF
e+/nxcXsmWO97Bo133ktDJqMu2VJ6knkDn4eOSu/IPDHATz6HnEMXVqr0OUVKsi0
ur08TkFN8QIXe8knoKKq9iubduZRBqDtQ0PJZu7UQ4d31G1R38FFAsmvfOCYMyVf
wERDFkmpQNXiB1q0v5HOMZW4vSyEPybdn0BooMYbdiYVwWVeMt4HE3tfOUY+W0+e
AkmaYYOIj/eC35rojnKY9KggkYs2S9qeWlA4QIpQ8y2gFhX+kRiTYNhDA6oU7SYv
sTCwm/508FBSMZTgwrest4y8N9YqTj6KbwKXOGKVQfFAtXtGzHVuQsGj7BqlXdLq
jglr/Fz9AHZNBhG2D019czHiGzNHjq4a2GqvLVZ8NxLKg92JrBWMqLx9WEi/sEv1
mr21oE+6p7EYcAcs9BzlA8FcBf4PFY+KACaTpuOmM9MLxBHX+AtJsG3l0cUF5Fe6
ZBQS07AiMZXpU5pvX10sij9iVy0qNW9DIcS9HMsZIlvAN5+RTGWnRfm4wJuj7YQO
ntzfNwIPnPmNrEqjrhmAKWB0sXAorMEtV84Ez0ZI95Ca+Ar6xpxHezshw70HPWxg
bM0d298xYZNxgzQslbtSbVqAybgALYEXhxqqB57rVxZ23JGPdwtmybF1ljQc7atP
ZiL4Tzhedb6C9n0M14rBpDQbWzwNQRc0oBELSfRtuNxXLRHzgbccyjXa0vtB/W5Q
coiQxk3TKR0tzAorbm6vkXKNC9KWRQ9y3IyB8JrRaUOuVbm71gTxPFBOfcnms4Hs
Yjgiun9F+wv4LFjDvS+GDOyphXwUyBCVxapcc3g71vm8vFaJ9JVfqHpbHILL4sNO
T16I1KDftg+yyTbe2Ad2XfDfhHzsa/hPqsaoNJZLNGi3dEqPvQ9Rxr6+hHg6Bb+x
9ci8KNtMOVfo74/K/dh0MZQJhnMFHIPy/v/8kcneqh/iaC5IQBfreLG1QReqPpP3
0yGI1Vi8JtQYJMDfDRS1xzu7KU6H3IvWc+PgDHSa+D0/q5lfUlGwtXbaiRrWsgxg
LfzIVGmahtSwhwjxa4Bj7o9IjnWRm6DwJ3chMUGRgZjT75ws1bYx8KNwkfSaV6PZ
mbWtQSWTVyOALmGelc0WMrSTBN9NJiIjD1lnLvkf4og9BCx60CBbUI5/4SgDogzh
KYDbs2gptyYCIaLpa+UopRCl/vCErf2geMhUpVM33x6XQ2odnLXo3yq3s+Atiz/x
PCHItnxpwS7AUy4En0AHAQajQl75XsWTR2xwiiOKqClu7khaSrDpBeXUdZLv93MV
vkoYgNPjYfkrpXZmtRpKhMR+0FrL6vTnaAObsOT7vGOV1gBUhbGn8/bobVLz4akB
6Oqg90+KID79RZiMRsyFTcuNRUlXoy+OqgydHl/T8YStaHARb8Ft0cpWAe0ZV9AL
ptPVDMz6lEomJ0+Ga6zsUbYLJBTT/C8hLwxvoLHaldU8ui1wtYVrz9Ps35H9MUjY
1pdJcWRK7MijYG6Di7gKRWopQa99h9xjhXk8o6nTyEsqa2XsPo21gkfiXOaaQXIC
2kB3Y2PMoarJm1km4DiiTfpfzlLHeeALRUWEe6bukqfAZ4P9VZpFdGEcCq1D/zIy
Bog58BRkhuZKL85We86PcdkDI7YJXKS6o7Ft6LEZ8G/wtaBQuQ98jhpIbftqBHSI
l8/aB77cuENEo3cy/9xxSuzRjGApQlGpLXEzIjaJfDNtdjmMsSfYeFvbLb/aPaaS
LkM6cTREJiJtKqyRVMy9RCO4CpBcVzlnMAck1BtNbIZO37jC1zeNpitN6VX/aXXA
YfRVGvhaQ+fj5grrB0zAVo3Ui4j6LUxp5awk3aOzoM/y/vKxfcwPkkVndo4PG20I
pjz7uvreKleuWpHA14rpQyKLyHWMRCXjKg1APDg2GBISCuCLMj0YeRR7HT+8pGTV
tiLEE6HrkGuuMnHZjn1l9lF4NCLshBnGwU+R/UvlyTRBzw4P5j6nBBDFzEM3N9o0
ZyGlfOmmBRVcpgXt6bO+z5/8u26pigAl2PvSPCpi+6nlqX790dQjsHZt5RGCDENC
IML9A3ukkXSt6V0l1A/8vatGZkYqsrAgCSef5B6N9Ku+ieNOLZ/z44qKHIkX3mzd
gtX91tiRipWimxvpLzDQA0enF+cux0OeURka6Ag122xnSWBg1BNLw9J0kGYWT3qu
NFWRylN5Tcwptq3VwPCKKVj9IBoBvmhqBs9L/aPopS4I8CZWVBHxucLleLTIoLsE
6DaujKLBZ0m7OqfotB3yldAxZbt8lEQWLflC930npbia30xPAD+3LbJPaLOq+jGs
lmPi2TdcMaBHL8JohmprhOrU3VrusIK6iFi+zOVB0Cc5FgSOuX7aJkJGejIO7Esk
+jo7zlNPI5CsZd6lVeNqO+aEoyAV9MD9LdjxhYMSCX1FlvSozfEDg4+HYDCVNZWN
C4aYyL6nQHzn6Xo5czxnBh9JZdLATpvselWjDRGh6OXP4qEtoTW2DmEOL5k6rP/a
AJARXc6fdfvBPB092U/4S0OleuqkZ6wrp/a7XjvYjr4KkYb3w+a8H6KRNOL+pqvp
LxU+nj01gS/mzawpeRpVx1dZw+7J9MGSx4Sb5IlLrtGBSNGQyoTmRaBNee38SXL5
OHRnbMenSi162lFtvzdewrXHTLoODchg8d7YBoKybh7DP+v65rAOJrh6bVzjLO/W
LrXSlcBDFoQ9BDcr4P+o7riBjoR2+DRhyxQh7FWc1xy3DGRx97yYUa0WO4QdD7c3
bjluUSy39BEw+YCjyZSu6JeBxls88D4H7Cpa6v13FcVj0P/bz8UFAtdc3EAkADoz
neVQMcwA/wVb9lYwJTd2+el2hQ4v9rLsQT0QwYk/7WLNQaFeQ81pzXizv3HDnEqu
/08HepPlQc2AUOQhD8KhHCmQHbKhx2YWI6i6Q879sorD1lN2l4Rkndeo8QnTx+5U
UPr4GoulxIbVaondcMs+xYjHZ2Uz7mRQ4mvjTw57KPSqjCfMV5CVXmt/rJE1uI3W
KOZL/Ayqct3W9BGrt+T/OOKTRHAse7eO+70aC57AWprcJ7TxF41o6BQ37zDb+S/n
fBmZUS1NEE4h2e3aG40qCFb+sngNmTe4d+fvWdY0VDJlIE7LTpNfDStk9Q3Kz/Vi
8oXj3mgvJCejjpHRefZLDUVc25AOGA0ZIsbVtmP8lYo7DnH8vNu3HtuGDta2kdU1
TWtMQVlXhT35BTAdLxp3JUxtxH9PKHOZDiPybQt6Y5oswBa4UQsVumUWUmYd8cJo
Eio1UNU69qSqxuUnaON3kU9999SAW5JjG1UJEmvwKLvK5JF4dfD0M3X2OVZqFu50
wp3v1QJVpaOT303soG5ZbTm0wXNkTNHXM2ItWyLI9I1MKzrS+2HJAf3pQ+mnZdLH
JTgtWR+ekZashMu5sodj+rJHfyEYhYoDtBCzbhrc7LFrVHa2AOxOM6id+5KKcAx1
i9+tQrZ/ILT4VvvHob/dGrqZQP3fgsg25itta0KjoY/NIvrJs0Tkfrdc9upsbZlJ
trvPCXNYVWzNcCYkbbiAZtqb/9ZSLUF/VVL697BR/+p8EtQRrRqWoGGq/sb9XuVB
hBgu7icIm8sKukrC1mp+HjPFqWgPoXJqe3PVkgObEn94Md8vmIUyDqk0WIdzPzBC
8WAn517C6TRTJe0PgP/ZuS5tEASybmDvo9UP7UBa8Ygpau/hHGF8yVBzzA13IM1x
c1fSz2HJAXj0vOn0bTmz+eYDRZtk9crHbWJCcs9DxPT50m/iBzsjdkLdDCBDPUAs
OVN2b+xd/FP1NVONrDzZBcjlq7kLf4uMS8njk17RIwtmOqTefDF+Hbdze4AlXACY
Eb0dey4Hlxta837TPLQy5WantzLZapVn1FFtHJAnc0PvyPCelkp3pStNA3/+/T6q
8jn4UUN+d+/C5dwRlbDoH8HjmoTscxq1HLRSNSegbWqL4bS5tiuDr6QdjcEWwnv3
NQE59I81ymPa+NYVPo8CNiK/RWdviVgZzxmDeoCL4Bsr6dBydCGEYjrEry1vT2D0
Wd/8CuxnQhNaRUuo8swjJaoUGjiybSU7ZdqM69REYZvn9lp+sPK92T3n3La//gTb
ZtRYgF/+Yarxf+XPaPd8JWtQQp4KEoJ+7YRNnvQSAwXnRcY0LD83TZSihLTV0X0m
/G5HxHoTLXsBN+HgpOGQsl77w+5oxgAYusGjSm4RVsyYNUcunNQZDvJvK04FpWzH
ePd1SYbGZ5FV9Mh2TVQXrurcWeEs1HZ1jLHnLmCyypir7JaEcLEgxbj0InudIEjH
1xErtkH0nzO8qlbdmcQIyH+k42EJY2uqPyPDEJINj7LCjIq4eOoNNocAq+TiLN5C
QMGScu8K/7vSfSIMQVBUhT4Kk4mzRJzNtRKc5uLUxLHRjAXJdXUUfOTQS9KGvlUt
JfhdKyI1+YlOqDs/WVA1tiTq0dgOdVOOTV3w3RwwIJmg69R3ho81jfMgE3syg4F+
+eMc84Nv2MhaByChLwtA0J9dE5rNJaO4TO4P+OYd8vL4Z/MGcK7uGNAplncxM/r/
PCRua0DlQ6McSa/EH6fTUsbxjUbIP4HCzX5CzjmCT0DRVRjXRED4NeNi0jB0wp+l
u3E5FFWl5GafKDvLMNspZjZmqgfhwr1/XkC9oi3VaDQp92nrzpPRkF2ntz9mmAYd
BZsVB7aEJT2U8V7z0JjZeLAObBglLmo6cjlgLoKKepN2BNh+uh45dKN19YNcF/qR
0xYgr4IynbjXAhSwYCJ1WrmjcN/EzHdBEF1UHEcTM6I1uegmqEiVdqn5rdEcBbz8
/GWTuNiWOoT4ZrCF/6qDU9KMSL1rZy6eYPBvIfBWYFq0hwC5GLMHbkHGwd1zqZnP
a8p74Y7XGKgaruVy702uKQCyAtJUHczzlnsQE/on+rQM6q0X/MLY4/HTdSKWn7Yp
p9TNGzONjr6TD7HU33MNpee+U+JtO6yVklvwx6/Paquw+mtc6mL7FhNIWptFokaa
rWJHJtm7W1EG7BpBrkM6INtrUitvQNzp0+sN78q7mDucUXijGU4t+WB1wuGk/SCY
g9pj+Aui+yu7yMmlf0nLO3RyhSTDGuqeHk4si6hBsBjGibBABMsH8q66/+NQUOnN
U4o7JgQOsiXTOZ0F6Q8Mva8UO+xOc4/RkUC7I2mIQ1H4i653hr6fppQr6yFSu351
TVuSflK7gcM20Odu7+onxRlCJhs5n1rV0I6IBAi35tBee26yD5ECOz2pVR7H/sq8
S8BI+13b+/zxAwpyWOWT4ofcCS4sm8SJAmBTqoiJXoX/bFGAbDD84xKs+6a/KQbD
XmDySgsVBTyKeZgcxYNBU+C8a8RPLJIZSLUmIqCw4pSqRjK95oz4uCulwOu8sdwo
zLHchuf67F4LsMXFCd2dlO0wHp47qEIikUQpzVqQaQBzvgi0SWDWfQ2KdZyuzWBq
eBM56NfKjtLUV/oisytKKnD+G1hzOkr+Zq9uTSZcZ+OvWD2rSaNFtKAK2XsIqMqe
iU0Is54QL8AY0egKazjkBQoAIwCEPgHiMyJrGLuh1nfVM7c1YQTN7y7EGpcJd3Cz
eccdlsGInLEr2PA+4hWdYBT6ekmHWqaGZxZah2YEZq3Ndjf7+MX4v2NT8STtdQ0M
DXcxI6mz0RuL6ZSp9rIDciH/MP9Iyb1OgO6Juj0fO404ysqUXY5W4DqkxCiQNDhS
SMK0NjcD82onF1uuZM3AD4O4H+RUfCa6x8eZGhqs5Ky1MX1qohgFv7G0GEQV9V3+
wESU8XyVTBTXowbuPAYW5vkWUW2q9uTNZeKMQvjlpTkwPPocdiQgqD2I0SlJyN4i
iamcbvTK9pEa1uorlegRc8JedvANeQxzS9y1qir3XZ5hymgVK2bhRQwdl5Mlbd5C
fydFXOyHAxIKedpHgZ3FoM2L4P0Y9/hXGaFOWGcskQ/L7vZJUBa8MP0UC75ehuJR
Tq6tomuhcm4ub+v0ICQ0bKpUXW1Lpz3PfARSv+vBpz0h98gPsDvjWedq45etW2vP
Qe8IIhptowRgnAVlhqyOS0BPMWSehakb9dIq/JW2VIirQXD1anKMIbsy4jyMxCVn
jYb6xpxXTGoTjt92tmr7vO7MRExjbL81faa0n/tutyYLzvl2GxADTloaFy/bYvw+
0vb+Hu6fDQogoXVNqy1/6TXcLskLA+H6KRd+d6Dhn+1Z/6r2ehtnJGr4Fjw2V173
faVcP3ZQ7RsD2jM5UvB/kPekegvC3GsJyldJxuE/PoDs1oacMEfWjmhj3wkUK8bB
qPQq5I5HFsrl6O7p7wZzW55NznM3U0sDiRqxq9tg7F+cdFnpQ1qwty0F7lizhGPj
ip2+yeI14cyY68RgAsIhNwJgG46xGUHm2EFc3hrwAPaB7Umc+bvD+z/bXzds5NqI
La8HcxrsBOYdBdcG5Cuv9XFrBtKFNMyp0piUxKMjj21HuM53WLlzxn0lwKPWJWQy
ziMGACDNmAINiljzFkY0KEXiD9KT1AcTZyAVw/j3hL6qLsUTdUhI/Qnn3CtINf4o
gh1sM+SJG52De7JoWXIUt5PK40c3bNXwibyunSji/jrKPJYfeot8YR5mopQgThIv
Zqe7WHU/J8rR0+RLLw6F3eYNg2c7QbdT4hli//g8U8l7TBmWg6RtUdmxKNd9WdE5
vsgPf9NdHe0uTqluQojz/8c6Cr+xvDtLvBwDVzmJTTg6yQrANIgj2YfpGn2kVmsz
llUTDYCGaKIODPXHSTPJ+71LwLuuQ0Yyeq+VNpJgghV/6EFmvlij1uTI3MFlax3t
tFazvSfDh8MSpINnQfJl3x2c+0SAQBIEuzVuQDz9EkqRy2HQtUmCk5IY24mwg2jA
H5b6s9iiYFEHWF17PB5ZbDVyFJZM3Xw5MLiiCsCxE26eAuaJWUp5ZSie2S3rkiTB
ds0Dp9IpSCtLmzVCQiJweXYjq2WSTV1oUHHQ0osAlOZEOUgNH/2BePU9Gl6xvqlj
1tPLryyvXH64mcx5CwgO0hkuhZi9TLQK6YfLu6BeGvDMt+eOi1wysTr4Mbi101qu
7eBovXtbTqwRl77CqtSAY7KT3/RrJgdLJ/zl7d+mnAOe+om7I43nyjEID1jf5Nl0
CLSut7K6TGueQ/FXZEayYABs84VX8GT7Jhzmz9lwG6ro8NePwYAF1bFktWYYzkbh
eIJg5G8pgeVqFAEElQ4qWPlIV/RdKqKGAwnpm5QgWe6vs6vOpOVky8ttfeeKm0/B
KHeafi2a0hJ3q3V8uZWlpl4ygLb9r+Xjy/M0eO6eiR/iydndUrDaOooCMIMd+oR9
ltn9S4E+/QphI7eDVzl0+4t+/L5DKC3GuDHw4Vri6DdvA7mtPYb8q+1MGg/PjD3N
XEoVr+WVCl/KcTMIQwnpcQXpt+Pbb+7zN2zoSfxY1zQtnB4Ll8ClVp92hM2V7rnF
2rrkKRCN/XfLXJB2gvq5Wl9VjntpVignLhBGmpg7tOe4YNtlB7FJQN8PDMVNB2Np
W3XoPdBC4gq1CAJdkVXFDK/i882zKfGr9vXo6EFE3EKrQ5aGMAK747dDK+C/VoKf
0eLYM2XAfGy/hzlebSRm6CyAIzDe+MhtH09q+I1JMvEKkADJypctjZUFY+t74lBy
zt58aEjJBZOg6ItTV6oMQoIWfZ9GkJFke009aIb0AgDYUeM0vtowefJfx97mAGk0
9+ACqMoN4hOMkHkslWepLO0eyY69dY/VHl9rujhThbKlQEv9HElqXeToU1pXM/B4
BCFfKrul6xhBtUZ0SRsFdE9NASYkwEhIYtdtoqFD3FDRjXbkIf6Cwt2uF6TiIPI9
asO1ZuIZoR66IfvKzNY4n2qvO5ogASVg0JwAUx9zsqIOf6QG6UQi0SbGEXmqdrzC
DCreu9/9cRzrAAeKgnekGwBoXyM51GEZqvvlGh1G0YUoAUzN3Jzbc82NDyT84lm8
mvHkdrPwgIAasqeHtCpY52WZaCTF1rJfa2DmuNZBqTT6iC0+sdlGJbuEcoSi+K/5
GVexwGbNdUw2cZx3zJ3XA41G1khZXJ3Eqv9bYFQ6kxIsZqqzysjUu5mTbmYn4kK3
GHnRQBxai6fgX8ghcQrS9+eOB9hSox2anCLUR3iHCUlJc3O3Jbka6I7bv58cS1NC
kTcuIUixMmS83NgmoXp0isV0OZJz3vDXUQYy6ZA88kcON1dWFVCGF+k0Hc42WwDC
UgxdPKVW0z06+Sq7ESk2Q3gZ2IuslVbvjCN4bzRTtHhvuXeuWvMdK6/I9z9fudRp
uFVw0CMdz3EB7CYzpUDXQWGYaLloY3p/4fwdQ68HQXvY9efBptZumlvSNvgvYFfN
7W+RzNBaAhzHJsjdKkG7qslJspEdFeYTLRnxl/rt8OJ2mo3J6iE9pWwpiLDYt31N
ImX71/rAMik1xPqCuAVzVcVJOo9FKVUyry67x6MtO8A2bYQz/pAcgkKxLTufJ6Tr
i7lDAqzB2Ss61fMBVsgLC7THAPL3FVpHOS8qZPXkElyM5Od4ao+Y3T2Fz3x3reYA
bnJqK2E1b2ERVRtQ2FIc12sQxZXozbaGBa60FJjS9zXLvB76xTGFysgksXTmw4kR
oUIg9PtwhTvTMrcKrwf7WvOgD1xc0Ds8BBFZQa3N01BwgTB7VHe0MozAQ95pV1Zh
L3FLAwS5dbigblPIQ23bmXcoB6fGtwXikfjIRAbfxSxsgOeqdx/0jEt4vLWe5t7L
l/kvpAFi0PiONZOZ1ixLv9AMLBcNFT7PPl3YYAIABrijw+HKsarz89IS/BcflMlv
4rf/zctjtusXh5S0Tydc54HDMEJvIL4wpmUW/OtX2MXmt6tbdnMgLEQDNMVnfZRU
r7koX/T4Gvewf59DtUWKUdWBs+N3IUDCi69kGgfGzTI4VAqAEjJ7W5BiqUnJThDI
+8sBvbBUmT0ko+LzY3xb0JR1RJe4LxRibfF7Anwg9UTyoAdOb8EirKNzq0e51uE/
5WG47OeL9YLanEQqSyVmQe5XhNnevmfvuJpcCAoVSQQLC8yRco0Ef8oO6R3OKcz6
4gEOLb3Eo91NSvwTvurHWX6nytlbpXjjUqAPhw9OhbULcqVN2Jq0jy3rMu7+xBTS
cyoZUOpghcM47XBZNrqKKE2LEWoHpwOX0HVSfgyrx7KUE7BVNbNoM0R/6b+wG+cQ
RH/hslWtrKeTV52qY+b3m439KSakEK8QkZYkM9UxS0e/wfCW9i/JTqqFIuD6Alg+
MzO0UPoajb1P5yXGx+pMuOeQcJ38sK4UYbvD7/7zzIvTpDV4h4pV4tdByv3XzXN1
MhMjxmLMoGiZ3iubiw1AY8c0YdgFCcSsPYVhKgWfSTWAHvQOScZcOtI1uhT9hLnf
hxlWYPFtHx93CWM1mjXsl1D1xL5DW8tiC5hLWCpu3Q4VhHer9R617P5isJKUtcfv
LyPWoY2V6ItENj0ruigvA2KmcCXbh90H+b0jbfUMKnIY3mJYcx+23cBo6Q3BOsB6
i+iO+sdA90au3zVha3HpDd9Nr/ijd2RXKK9OYbPDc75Jp+T/V7WE6QwhZ5lWV7PF
qzTLjQqEcjxbm5XhEQObRxhW0OYb2ZlLD29RDI9havDvs2bp+mWph9FUkdCcrPi1
PaBOCOjYkQTVoxShIj4UQviBlWh0zB6uyyD+246sMirT8mYTTa86lKX5sLk1tOmv
6OTm2xTOp813j5cN2lIC7nFiGHymayhkRHlBiKvpv60jjxy7y2DKS0kfnLxahcD2
yoPiY/ku58SYlp+6THDOdPgweegGOzplEr9bbYbzEoaa9m/fGGiwtbaml4G+H5Ch
BY8MH8JhPIrQ5q4a2exewKM0+fOEvLiOd6XaLG7FuHoGIlJgtSK0PB6UT4wv8+CT
hUd8e1oR4DIC4V5obbTSrUp/cP6vJ073J4ia2+S9dtxJM0Ow0nh86ljD6si+WZmb
IRE6gP0NrUPrBTWcMpfOuskN5eAepZn3iFge9QtcRHj9ue4A00lp0BNyPbznG6Vv
ZdHXglYIKcyaaObuM1KpdWvliRa1UHsmv0afb0Bc5EP56J6fp+Xmn8MXrGOtB0eF
KM5sJiepcMO3DnV2dER0JLN0GEmngozWD8D4Tz1YvYBYNZ1+HqGPgwlpmLrBI+RP
/rr7BfHkwl0J2bQpRx/xIOs44BVEyVewQK0l8jz7YLmBGlJbsKk0855ePOaL04G5
hPRPyRE9nZQxCxQIdDQKU42SeYFxwr1nLn6SfZewi3c/5j/Sb1G5ZxDYFFp586Nc
yuW71y18oZ4RLH+Xabv0o4uC4FtqrFTBdn3MS6Txb/AAiGXYZlj3zszh4qJ+H/bZ
dNyAqDMmLEQx6yLBnrGA5ZIZSx3PjfCZ9I6qg1yPxibTxHyqSs9mQ/PSKHx8re/J
U8UHtC4vUgDciUyGdncbAjqyVcKbLukyZs2dTVpFM0EceclPxKAIGFW06uwLgTB+
E5erxwZUyUBMzZ25TfobS6B1Xt9PWWb1bzWqQdtsnPYCcwd/Etnmx4SmGoUoTRr4
zD0prsWh2Lwvyj5H40ia63erafL6eB2l//45UgWZmrqizAHRcVv+nYdjqX8m0Hl/
01pHF4eMN+T7iZFLFsSvnckYf8Sd9GgwxT0kjSVHy3KdPGoAxtS00L9Hc1keGMbJ
ndyiU7wcvnffbMuVzN0CgvEF9QbDF67E5XKqADjpTvAhdHU2XUuL8Gyi1IFh5ql1
ZN8KoDFA4gBy6JzRoU89lTgsv8HAlSdm0KoXdriP+TSPZPHhSxZMsHhJzVoequG8
iMajfTANpV5W+9biXzir4J6nqnpW1KsAILUJ1AlQtN0oWsZjT1MbJ34le/h+dg0z
OI79sN57JidPAikw+2qHRdWZvr3wiNnFhLqZHib5Sf1gtBgTK6UFzX3OATexOejF
FYg3dqgEIi3t1y1X/0mPOCFEUX7zMptIOhM3Lzk27Cj0oHfYwYM94lff1gPHxAo+
md1aH6JMp9Te0qpzMRNUl/qpfXs/VbEmmnHv/iuT0hRNgXG5YKJtT4Rz/uiQElsa
pmDaoL+6frkfU2Yy93F8qtgZ/1dTvS3tMvzo+QBmJd3Bc6t9JmHbcyDp/4TuRJNd
aVbGPUGNKZRHCY7xXOl6eW7iDQS7xm4jDlGKZf8BGr0hfNQ7JHhLXaX93DSyYeh6
W6UyU3CSTAf0CqxKCNWell07g8hktrK0+R27xN2zxSZ+X2beo/IGO8htrwmf0Jx2
brn40cAiWe20WKYpgTIjSoKnmOqF6XZke6/vJNmJBUZZFuE0ryxYTwrnqAhiTBXS
28N6lltnSAzyItGp3nXnl/op4+6U1Xa6zZY6q6Z9fHr0trkAd7twPAJi9sF/Pcu+
36vRT6bRV2DjCLiEktBXcl37iK11Rj0WKsNSO6UZ+pzxR0dlEcHWKVYVdenr9ysb
n3d5PTv/hS3jdhtYAjIbhM7W0igjGU+Fr6m2WEsp2W0hFnaFLZs0k0RQXES/JB+J
NIH9qSzibtyzE1m8fYCUmjoY80cEqP1Hf5UpPrq0wX7Kk4NscEdSewUhDvOa8sUP
OP9j1UUIjixk8uwI4F/FFZHE5Dsou9QuPgD+0LkTIM+Mx8I+hNZKmjk7sCn5mxjn
bre1k1vTvbuBZZCikYNOHwp1RvIZpkI5JaSfXf6UNZ8NO1ojz4ZE8h64eoNmaXrC
R/nSsjQBMeg+q2KUHvC2xdSzkK6vi6Vu0V+1dJphKW44wBagZbv9mAkV6ak5BR/t
U4WIHVb7ePMaN3/ddNImPP0yxuVR2icKuR2gKJHHigd4gCz67/mkp7RUtteSqHuv
q7UDzg6yiFTDdvb+EjPYzatRUAl+G0cw2d+1lkvhwp+wls2nAzltfRJDz/rSnto/
0Ml7btuq9OCZ7eWPz0OTBzpuNU9w+4yZs0bTz/X8Pnap2vcQgT5I6l+4HlkDoIzC
qBVJImLmbjduuwzirbTpZN5YzbMpeRtupGNKB42suPa8pW0ATA1bRl8imCqfUiVv
Gg2Bw1W0Z0Gh4/Yar8TXXoyz4EsjyX6IlCO8kvhVUjQfEvwdDXaS0lnjIXWyl8Cj
bjZbDYA90Yq6O5BO1S0/5YXfF0HYUpQr6ZEdwx5wfICJC66Kp0YGNtnmnJpC9jX8
VByAf+D2CC9+T2YuMgPZuaJXGVH/KWxyqCtepk4PT75cwqsPQbLxqZCDfu99CuAY
6aPmYjfzEyA5F/YmymbBKkJbWkbgFSRYc8J37BWzjg1nvuTFWIm/bbpyQ8wcGYXi
Xb8kAFhHqc7gpWKKclNEW3dLwWgWwc3BMSltNCMWFxqY7TDf3KO4wNBVBljGHMzs
rfbOueJeXetl1hK6vsi83mfRyY7Tb6pZ19FxT7kF0QkKMCRqSTYHQARG70g1YVZH
rxZ/WU3DHTB4m3KgEQhRrDOq80n5tUTVvsaHSGOMwSvchbhqBZ4/LG2otpgFqHJi
l9LBGrC/0V8xArbOAiH7fkACSFP2iPpVNk3BG2Mi/aLbjks1qB4bvNCDPU2b71hH
lH1td1kmh4VPLTXcOTxczD2Abx1D3xbShoI1KeYJgpXDZcEtYfnlV6+5WENqzI/K
1RbrnbmrGE5uXoh/rsvH6hawwjPev5vaH5415KnrqYE4gnbCUYyLFOFCEZ13Ye8v
Dl+b3hYGxz/iOQJcT1OBWnypYVGlz9PSJ3MqdfvctI6S4Fh+/x72eztGsMaGfrJ7
Vt2lfJ/EX9hE9cpKTkwTStRmj9TuY+IASYZ7x8k0DhMQRIbYshcZYkP6x6g4OGEW
4RBwsWLw0seHviKqqjRL22K64CKBlXHqQ06ggTk1pRfgJLkuDWEjxVkWeaWU53Nr
PQ21758OoUX+NRsfJRBk/hkPTYkvkIsKxgL7+elbGELf22TlCajkSou+1zvp1kFC
Sm2djMdeVYJzJB78pymVzjhxPrMjj6XU1FXFIBrAY9iCSSTRvOCTix/xy0Q2Mho7
NW88IMa7CCDDT+PnjBjgnbcvavyi4536ol2FaanCati7Gjvk1SRn4l8W6SXuEotA
GGOcGUYSQrdfcN4vkl0w7YNPnf5Qn4KZrLWb78f6OS7ZsJhtF/ABStHn9T/XHf1I
d1Bxh0UBRacPyP6b4bxv5H7JKP5PBQg34XK8e96egseR+QL+rUelVcHE0Yzjb/JX
OZP9JtbhI0ofcfonbVFMI83fsgBIrYZDQ1HZtDm9Get1gXIKehxCwFhV3LzaDJRB
dYoYf6C4hF2qVekpf+wCLo4IrP0cwGauAHRiYd1GtZTzj4/KbkbCtYodu+z3fxwd
nstkcwGytzduq1p6p5GmvBEXVXm9NjAKwJVq/FgWdmw/9RQ4akea8pncTQH5vm8m
0MJkRVR14qDT8Ko+LplJO0UcuSLDA8x4KGRnJHxGLhBDtzoWAYdwnyPtvcfviwBi
zk5piMpmR02bQSrODOBZN07OTn2ipYC6TuZU4u3qIZdjt1mgRAP91vv2Ex3JDmqj
oQ1gYMJk9xoU0SwDoLATF712X9ULqAZtv1GvepZZh+erzLpMcEJPLRi0NbRxfH7o
t2elSHEsuh8JuFNL0+19E64hk/adSINlbw+Y9+0h/g41tOAFlyQuYqctahV8DpqL
a9gdlNWtEdjSAq9TzlmlJQ6+4/OdI8wh5/ldNkn9VU2Ziw18hcu3mdWPjOY/hbI0
CiAgNLpxTOKVWqaTZLd6JSFImgDRp3p/UheJ6iXUeQgSSaDn1iTvbxhstqHn4oTP
JFRqCvLmjxDvUnWvqm4pNUIWoX7M4OenuDGbOwciUVFHGtgKUAwK1y6Inz9PRHdC
e1vyS9+QezL3FtMW3pSZ/ZnTvg/Qy8TKifEYSxSodi1R1+0f2BD9w57RPOf3Bdnj
KDRtlCK2Cqh3CvDYtkZXAs1qCvcvANXJLlMkKFwMULw2AxyzppqRSfC3E07olShY
b6IUBK2El7XFUqzMw+wHH3UQIAkLLAM9lfLJ6X7Icnm2nG1uhwTbFbCdmD/B1pD5
kZFk80z1ESMwcI1FXn5JQrH1i33WUh/fH4RRSyga925u0hLu3tlWG1tHeAEhpl/E
QROdy6QCV1+y0qA5nkorWlBY935gUO0IZXavwAGdb4DmB76jIeSae7sUCIgq/JhM
CN4cpwfjiz291Njlfm9mR62/+5z0a5QcmmltKC+DnTnTFY5RxAvn5NJuju920uGb
Y172QYUBupoMGVTVOXhknv7xQvz0l/PrcyPBNzVN4mSVb4+ttTqaXalvNbL7pDob
hdMQf6Llwcx3Z7DquOYgxrOgqVRJazQBKWuumsIu536hRu8Tf0FyTdTOY3l3z4Ae
3jWcQYhfHDU7DzCZoMk7mW9Fvt+QwA0W+s/gNX2lC0mwD9I6NzeIyU3gtrJ0/jYB
EPfEZ01uGZWwP4lGvxtGus+jjDr6dP7nz9s1+uqRCjXiBHj2SDI+cHgDgjTFqwww
TzOdgdqSB+xPIsCoWzySTug6vBAd9zh0SLVX928Px90Fh3OXskvNKPZFggIfq1Cs
6Hz7uLqwmWhLM9abQ0XjP5QGjmB6FFjWo+p5ZmvoFeGbUSfX5UXfPNogBn6yI2LA
4V8zMc6LFYevRxRE8UEdQf5uq4pNjALlfZU08wMRJJKtPbo95xqdYethK43ypl0A
cv5E56rR7mZ4egUnMRv7wFcJoRPQnAkwL+PbyzWE+XvGZHxWrvM7/X+HXmStah0S
YVpAw9nkMhuWdsZeYHLNajGdV0qFzVcbhs6a3NLAturP6fkKGhZ2CV6KPXvXTfSF
2VucLj2lg4JMUJS2sw4fIOFfd9p6cnS5CXAXAywM8FNlvIGfiS++HJs8jb6LzRVu
hzteNFwRx5++fmJLDghwhMyeqJl1tLZo1mnjoRmim90SDiD9BdgsPJFVFaQilboV
a05IaMbYUHrJgbTslF1T6/xNjd5tZ50kA8WVSuZ/WB1Qi0rNHlPE8VkpvhLxhLvy
9Ikoz2Srg7EDZo0fOHU/DZXmYPpRJ3TNlx1D8TfHAjeKZcEazPUeQVhGiauVF2bf
2WpP8FSMH0Ma+g8IkhwSH561yTSQZuBcxPHMQpLI5z1FdWLpClbqMdDhrVMilrW5
1OLXw4hpC70XmvC/yfKUOQkG9ijf72cMj9I6OeYYq4ka9/1CGVREmLR8/8QCxkqD
9enQJFcv3SJUF+aCu/os5KAwK8SFx+83D7yOM3iOuSytHg9Hb7pTG92CSkzXYxtA
SqwzrUhglq8W48ZoRP37d0KtsW17PrCB4oTvwSvN8hfnNqGyxsoEC+8OjukG9vPL
eN/z9qFKOeXMCuLrBIPZykePlHRHN9flq0PKEw7wKy2F31q/lRYz7NI5wtSsQK2a
3+QvV9lo4bgZYmlker5sQBjd9Ltv+orc+9/ubcqiAhbyf/OrccEzLKCjG711gqxc
x7ZA2uel7APLvpdAP9ZHbPw3mr/p6Lu6AfOrMxn87rWvafHaqXQ8xPg9h0XQmdKu
ZOeyrUMWVcWUE86/7seeqrNAfZ92tfcxNqRrVDnsoT7TFRfwbiYNvxgeutW563ng
7WJL+LTSwXJcHV/ezKJyEYQrF/MSO984xrLVvkY6Cd052ut3OTyJ8WtnuvARACsK
4DipfHHl56R6EwsHYuFUqPH5QtUI8qO3RXEhACOELSsMJJ+k+kwtYsJcIWXRUT9w
ZyyeXbuEpviHgk/jjBhNzazS/ycNqF/2zH97V5I1CjvJiPyuRcgOKdNZBYr+HzTu
BTNvAN4a8h/HDO6N3d+5mCVRX0GZgBESgxnz0/BcxTzuY0s7a7+5mm+/REFcn8ss
wW6y58E6RiemGlfKF8QWHaTfoeg3nog81HJAarsLV9kkQ+cPysrgodUcdfbLYtYo
kFXq3wlmc+lRGM6UU5vDtIEasPqBytwxLSQmBKxkeMVsaQ/kVp+LjYo6GGD1RO5v
TzoXcwPQg7TlufGFBCgGALuQ94kKgE5Z9TUat5nSB1/aos6Z2Pox/asXgUHrxKwa
MtBE4wS5GlMZ1Apvy9Vx2yBrHtw5WMuqGOPijGweJ9kr2Dcm/DpsIJskFOkS/RLQ
CQ9ATNLjiIzd/dmuKT9fBANJRh3MwYNrs7bVqcoLXq7hSCHsGeCcYY7AyBoF0Stv
sdjgvyvARCkuafbFyJo9ISEfJEXRJPkox31vkOklpVbjItjG5FkAaEkDPBnJxJZQ
L+BYKNu2gV4Z+QDQ3IXXvSqKlo90fobWx/ujfgvKE5ANnKl6fbJOywZsGuUFAcon
i6Dascbdbfg+u2R4HAYlSvV4gKzoJT9fZVSp+LLCjFnYrs5bgquYhwgFoI+V6Cox
OXJQXcVtuRD9r4vkg7uIrdPy6W7k2088uk6SNoZ9LCUtH6EOXwHh6ghegXB2uzLN
5S7VC0OVqW7XiAoMVitB25J3rCXCG6doxc+NPIZo6TVOpLFiEH+RRBcl+q35VXBS
/a+amfMsH2JEkhQSfLKiJhDcX0JU7Koi6tYIDN0gHhXzowlS2zIi8NitvYNm4OFD
eahXvMg6hfFRjWbMxDO+r7MjX86f9kU+HWM8usQ+UbJQvRoWoOgVUSku7c1hWjbo
sumSfxXR6xKdgJdMOaxx1lFxQ4BBx852JxkUmR/tqio1m0VtNPqSj5XF440ke6SN
1TeXqZiN25EkxPu3lpyaPcDgdrLdOlwuPIoh39R2MBGnrTL+h8zpSfHWcKXrX17K
YwqfCp8+eZV/syv8zAqIxne6x5ykcysb9RTXptOvFBRhj0JxeAzrfNS8roJzcd+g
iCGcptf6Wu5xoYBeKUGX5oOai+/iv/RnsSE1AozGM2F6w/+0LtOTteqVZ94Akg8k
A7XIdoFPT5IqlDLycUWj8WGFYQdObAVKGk5bkZemKdYWNyqP/m+/eez5eZPnHtgw
Kzkx04dL/AdFQqx68U+wNkDlQqRyu9+9A0b5wVnBB+QK/ednFgLBRgwuLmK9aWzF
+2EtljfFGq+AyjujTh16vsr1Z2r10q7Jcv5DbFjBDuqz0z0XEbP35u4mtgLKDn76
c0aOd3VEDo5PCA1CnMuZgh47w8+z9JAMVAIkOBvb+OO2hMdpZDt090txHEePgfDf
PC4GUsr71l+5fWnL6cDTfWSWuC9Jyf6yYsihRBpb/qfSvOPd6xZF9GeJ2mGAsPdf
AR5JsGraTyrfVTOo6vGFgTIfisQl5V1p7ACa0wllFzBv7nwlW5zEHKoWkXv7DDt3
ugLkVNr/SDnpLb3AJ3POYlgUFKQHPYp3O7H2RbOyVUFOo/c2NWHgIncCmP/dEp3w
x9TZ+PCMhgJ8j8G/seeDlTT4Qq1e01I8KdyBGQSXr0X6kiCWUH+ga/7+iRJE2+xu
XX+qaHgQ8fyE/2fiizTNYY7Kg2ndoG46zcXOIKE8C9HcgyZdBpOB8F8EfKVhjCMc
q924NfXv7c13OHuzN6wkWEve3uLPzc3KtId5CXsd+IRXuwIMSTqUFO/i43HZhmr/
4Hl8/8PR+a0DXHm+Pspwv0yuPIajOyHR55Fr+t9Q5jqCQKO5rrL55iJsCuGMUcim
xNajiczWGpgCeGLbvcKCST7yUQLfkLC/gLIIizi0C82M6PEh1j1kNw8FENI3Co96
2mqX5lO2R9sg63xztivroc4WnRVvcQbdX9q6AlRGB3wVcDtI2Mpu/hOPb/odW6DC
es89OtzHPrUu3iudjhcuwk11zW/l74hCbwylYhKRX/iRK3xamF/04C3WY/OorM9z
rzJkATbapqef7Kis9frNaS+iEsEI1GEPC7CzIp74TasEI7ztZTzzb6cee9AzSEZr
0LZoCgKhdCKZJTnCmvEiEfBeCHr3NpFjID0n63Ep+CIxwocDynm4GPi6ABFYV47R
VTVm8v1+z2cn3xbJWHEPy7Ls1l7Y+Nf5x3jWeLghKNZmsy2tfCGoGE+JBEiomb6+
2SazBeO/OhXeWgAfQDzE/vnXIO0n0LsuJf8TKAyL21WWSvoaBOGzZA6UsF5o2YYr
myKbGOAsETWxf6aamojmjAcohwxDPqCm511ulSEatTLMAeILN4i5altNQiRLitMH
wWHaBSIrmPnMkEW2nwPSzO7S/JG7YE9iqSA2VfNsyjrAJuvwhF9JISbxBwgdHDau
z4YbxPiMRcrsu2JMVLv2RkpBO1JqqihY5AH1sbMDpNf08qO8Q4XEQwRZFuQNrXTE
S9CizPQYeL5PJ1/kRQB0p4wn4eMJNYYXTBht6neSQmrIYCy25llm9dya2Y7A4vOa
ZRhZ6Fz9o55jQw9AFdWK9ck4Ekq1mQK+j2RVIf0Ul9mhXA6sAadzQBk+bAK2wMh0
JjXeOrxJNu/GpEFyySAh28iPpErxuGGuuggACIxgIql2i2w4zeYnuddGSK+tXer1
HcI0v9Uqdom0jL/R9ha2hsOc2uPK65PqoIbVhx7Xhr/nKaKQ15RC80ada38sTiYi
KTxKW+WPK47qzRtF0Z6RhJJxM2R9eYW+OCB1D9l+9cOr3Z1WzdT3l5v6FY5ZwL4E
t3pl/QQNb53Ubv0S2u3ih2/+e/tfa990TkoWk5nsXxhsxPtd1g7t8GHu1y/D17Z+
8rk7hIbvYsgwiA3I+oDAduksB2DEuPoUQGX2AOrLboVcwAYUlVMvyAGnJ3XT16Yw
ZAQ8kCG3j9vLx5lLd6RqiXgp+ZNt37qJs0ENqH7rtTWfsjmxXVJYYtOjateBCL6u
MZnUT4KsGtqjqHo7UExC33iXIzNYacjE0Rl/a2uG+CKufG32J9d88IV/Ov5vweYP
UViJ6XkINOLn0St4gmE8HdshyAXADGYyMCwnkDL9d6fJzaFvrP8LSqJCLuLuMnfa
MUugNi6z13FPCIjWanSXNpwRwpGbtWvVabpjzZF9i0SxqdBBM59gtSHfjYo7tGfs
gsJUQHXV7xar3D8XfOH1F8s/pHVK8bfvyC2rntuMSl/8sBDiJV1JgTJOJdi3DHEg
smaoOXqIKoB4DczQ6ypJR4AV0glgbwlL5MH3+OEyXnirrWWJGhvy4Te9AbnixAK+
kZg47IZDqWi6wNklIu2WadFFAN4um1TDIS6vljSHdNNBJgx3N6ERS1kep58R/lx/
+v15YD+Jie3D0slzDLV6cjcY/bwdKB/aJKH5m2uJiJX9zWpnxPuwNPw2o8nobQjm
sesKxv6RVXr8Wv4i+tyLDvM/cA4Osb55NRPqJx1kOhEnu4rSd8SiWBu6tJStWCZi
38wH/Q5cE+L/PwAGyEH5R4alRhX2QCid8WOq8gmjjis/RHlBSsF1kIcX2QST8+FW
yny5FU6CP4HRk8XCEJpNw3MJoZk6GU/dH9ycmMvCnRr9gD6xE+RcUehZgyJGIBoU
fq7m3F/JuTWZgE3oo4fOvibszsGDZnv8WSk4JMUCg8OaCF5WO7BWeWHQq0+QbQgg
i5Dy5Z2cAaowoGVPsybonCq2QCflTTph0x7zAfEBh1LZgQChDsiZNVniZro6qI/2
HD4wzbWgRa7pZQGusdT7aBcNPBEBUJ92HGDKA8s0V1a4Ifj042xAZ+mYDXk2QTn/
Bb0KDapn4m+0uAS8ux3g2MqLD15LSy95pQ5uj4emNUB2G7LkMsJ3qA4WfKbZpgtk
ALew5XdH5fAropd9BV0Lp8k4pX6snHbHrhgZn8xe7rHAqJRz/8UYsuu0HKt8wnT3
ExGt01aLdyQ0bW3ODSv3AjgonNMnLuDvraBnq0xr8iIOyCEoaxfetvXAcjFwUCGm
oCANLErZWybPDuauHSJyZpvoe5X29bL4XvwgnRjbunvQSocNWyI+ugL82Ki60M+s
fLdOxViYk8LnIHtt1CdpJitfX19wjPr82BGShfhXDS3cP1Z6AoVnEJn5w1TjRFzN
RZ0aM9cjtC/2npdrI3GscfVuJMHJwy1OCc5ATrmSnZx5hrGZFfagiHu2MKE4jNRI
+CzyKXM5qIWM53nc29u/Wyn93IzU8lfRM0TFcslQaW7m29DD7mLWb9yNC5r/7kVe
ceQHDwDnD7+HRH81kqvPOqXaa8mnYyFe6hItoMTCBePBv6U1/2surN1mkODGQ1hR
32epSujsXtOiJJEVJXxGY1LdgeZLwW33CW+bJqmWw6vjoIiJX0rPOuMNUss1LNrN
zKiX4+IRcyxDIx2/UPpR9ahA98FQC4dEBwm5j7IHqZINC/tYkAJqcSE1Kx1RW2BJ
L22IvCZKWRiGJt8AiMRV0JCfaq03LGRoIxCwmUOP20MgPUCJKKLhQBp8lt0Y/MAr
AK3CncpXkTmOCbgCxftaLKOveNvR5ufqw2xrOpbQDvf4IVANp1kkuzg1UDJgrKNY
UhCezx56Guxxetn98ptmdH+x/3VdRdchQtNV2byzEpJ+ecweU6WyoxcOT0mIOpWH
vylnwOHiV3utRDbx8wnY13oz4mzAD/Wau87gCcXJxxT8Yw9zFZcCIQItDODFyN3X
AOLTpklmX53YfBP1TawwV1qu+N/X5nlrkRadvEO0Tia1/HoWphf7rerRRYTKKPIa
cwcq/6fb+igQYU0chNGr2EVX1C8tDeUEJZ7lJ4ci53q/IrCVnL1O8FRQv8feZ/i1
+vFRJi3OcWOCv+Rg2c+WS5dTCP7vT+l+lvr1VUTQQirNt9VlN0jZA33/k75om+rB
5EO+ekroYcawkmokZ28zpn49dvK0a80OfVXFqWwtEnA+PvTfRpqk3HhjhPSCdvD2
cxhbfFqDq39ZBzqhtB7+QXDQFpLdO9Qxq4x54aLe31ZUGYjEo3eqUoUfLVEvQIOR
ycKVgP58qYwzm2GY6r0BlehS11aJVvDYpmP1jkeUPwrdKdPY3D2njizpc+Y6fpbZ
69hQzuailGelRXUe4h2nnCIoDjBumcxk32LbWxklHmBHBdqt95tu8q4fEiZDypSu
8lV80s0JAU4YBwPlJK/WCFDt/3ITsEfCVabANL/UUhWErw61D1Wxc3o9y9m8aO3P
dtk0qVqCB4OpTYvmYuGbIXpgAN0cmvCr7H5DQszVdK7pap+q/nMqniFV6UvUoH2f
YzWRiPxLZlJs+uhKYPSB2qwVcsfbXFldQatCSNBaN55BZbJH8UYij6H+cLKWz+gK
oTKN3tPZ9mExnndUcNT0XcGOhlVGspEWtMW5bjMlQ3qhH/FWBWCq6MFHjP8B1WGz
NP/AZEyGEZORn4RWX+6++psx741JqbtKY1B18RyCYItU+M+JTmGIRPfAwSq9Lc9Y
xB/CifxvGRbaawMyfFNyZxlZSavAnzB2xIiN+CKb4zfvByTwY1VXxtHLRUp3xKws
XLU53T73d78c8STbHPwGGQ7vpAtX0P6fZpHhM2FQUq1t2y8cE7SL4F9+aPgXkk2G
C3zDRILRluH/jooOac/gUD61oUv29a8x7BctIQKiqtha+UcZsdh6NDGIjKDsb2Ke
w2PyWIT73+NIMkr/6FNogUxRe6c8/QDl4SE/eDTJm89a+VeGcJghQb0RdCPRGNKU
EFvfQxHHUAl64M39eHa5vOtdv7XAI1x63GlRTvKHj0VZV6cq/cwYx3xNq8/P+cvf
ehMBgZ61F1pnO4rG/EOsBP/EZBV6YCxS6yhpRBT+LkYNxeUZVM1/ZPmKEv7lrxPr
ON6K5DPaYy4HfMHVcfD1mjOQLi4SR1e+1vAPQlRVT8URAnq8bbGUgZA6w8JcbE4t
+ikt4JrRsNtLcEIIwjWfP141dAaG4T75uOE116y/voa4UrEUeDyf1KFYnYQtV8OP
u0A13w475o/T67JNz0H54dG38NqkTRlaWYTXzNm33FY58YJK2Mw7468J7a5s7Wqf
bgp0XC/EJHnh+XTDHXzz7CA/UOubm4lZjyOa6XbHhYNSyLiB5IlcjwBYMvEpO9F4
lXKGVtqD4kMqSp8ZC1OF/eVXIFHJNXmfIol0sh0sejAp/iGPbkE2c3d1m1UuHeM1
v9/km4C4BK8T+Vb/IAJ5fhz2zIFkQ1Jd6904qM3bmfo7WOrZ8rp43QHjQBHnYsQn
3p49Jr0MN+Bvkar0LFXnb+Fpd5S9yeZdEMNTZ/61PHekCF9i7evH9pl9HxxEwWJS
02lOblSROPXdklUsrsbsiu3APw7yt5bUE6SxIuFy1FtyRxkJODSTPvYMTb7hneGi
aaUfBqmFjb9VSJQeNVbWU4Beoz6TRH5UxjmZAU6AtXfay2F+WkdhVYDaftcimw0O
I8eUyrJKa2DmL+FxVPgcGYp2rqquZypMsUy9KftusiNP2RVK76laqUK4KSe9AThF
WxWZYc7Mc2NbxLAlU/R8j1ETmRROn28PX+JNcpLte7DH/8l+nf4Ftjp0OSXb3KKD
9pyyjpG/gNcHhsmPbAg8cztp5lnVSgxuyQ+JBNlrlZyPHOA9pLxERkxwYDNLIRku
ELjvJEeuQ2OBZJCxdP+G0RdoMVkS8UmPktgyjokuY93PDudoStCgx0gssFq5u1hW
Wqz0XVr5dgTARqr2Uyl0zQ+skQqWE+daz6HPXfZSlKRjwqK5/bQTpk7XFhrRd70n
lSmTOCvF/2kDDyq1Jihh7CUBeKSYIh6VvH7xxNQxTXPHdZX+y/m2lC86EZp6EdYP
yDn2kMsmDsh1eyXCR1N3nvsIzZNRh6LMuD/w+OHjaYpedCpvjCw0viUMvBJx2sST
1iCRpO4+RGLDtvpNMOOh/t5N2G45PAdShkn8IB5q6M5TBU6BkF4l1cNnvlTBxHI/
Wo6flD0wZpF+3tL5IadKWQJQyHnjQnKRjcn7VJdn9yhLr7/KvOFJUk7jEPDIbaGW
MgyjtsAamcuuW0hcCr31WFWbnC7QBjkjf81DhusrAncl8Ngj++ujInkbCSoblhoc
bG1ukPB6DvuNJp+pC/xGHepodZ3fCDM5FFiSPmSJ6vl2Uhkq8r7MmgKdty4K5X+Y
ISq0tSW6wcDnkVi/t6Lx9yVIjqJOy6aQ4v5wfq9AtfjBE6LSqhpRk1CgxqxJk57R
XxaujLFfPVlWd3rFcE0fsotoUR7jglwwQ0atGfZYCfzBXrbBzDUyK3B4Uq8fbcC3
Y2n7LA+z9mnbhqki5AROJVGfJv17BAl5YZnpqQT4AfBl9PgDOcZZuwDpHexuTuLU
Ec9q/t8THQJXOcdDi/y6iQVj1g/HM4zMabFecm9/8+K8SJ0c+g1uXdFIeIH7OQob
1gAgOvgWHlYbgnCeb0BllB87IzGqfOW4+2JS9FwXHUBzJRNCnigX5uYHh3sKq12P
xHmJiyphWuagKrFOHQgzsaMT1+woHHN4QS+hTLsEOqdrYDM6xHLnhcRxudi53SYk
7LmvsUQ+LxtkMUiAvl7SGiRLlr7m3sd1NKR3nv/5A+DnmlX7n7ooCiNdtSq5Ifl2
Y8muWVpB3ivw/k1B8KgrmeypmwAwtTKqAVNk3KFVf7rcSA5b0dJykt5AkzjdUBul
qXUPkE+y0loc5jUD71CvQw7BMHy3j8JBads5fUEYikRSXFRcsEkziQ3cOCR0zMOg
jturq19fXR98diCmKx81vBu6txlRCD+lZtuwNlJhZBuxPCvxbEiTqTiiqRezx93l
OhO0MRIFGBtre9tFUXrF+ug+H0jx2+J0Rzam7TbzXo2ShZIEXNaUqJcOQPxca3vw
u25bD2fYiMooQEDXuZjogWr1YyyJ07Gg7y9+TnyNOX15raRqNdm+ftTDwsLpmGtO
9J/aaGdjZhE72KrXIBfbqmKzwRF/ZJaQHkCw6Q1cOF0cJQmh5ckxRXuxEkMWc6CR
/xu1zTruaZ1mUBkoDjD+qa0OWd1VMat4Y3H9Z1Jx67wZ1xScOdCfS58+EgLSBQDN
GyyKHfK5rZA2QdyMPWm0Oev4JYBdwbppcd282wBBLwV7o59KGzNBhpIjzHNZPbMe
tKMAIDqnO6X9qJQtHacHRXuAJKdQ0OWogRvAJU0SCXN7Ba1++ysQScF0dnUesuZL
WkaoUPz/slmDy0BVj2QazMOvRgBle4kYh4JFvr0QEwOPbzxb2Rm1OtTEvL3gSOo1
KaDl13YCfP2Ina2gQb7HGVoS7g+6xGtyhjywMlELDkzbx0SymO4y+yYnfJOn81dG
IiLljzg6v4GPD7Qk9BBndNTUIfrWcB3MdxGTV+rzCWNG1oT+LKz7LfmA7IEtkFI2
qt8M+NsC9dwOWIUVObBBD6npxo0ize2aq1Rk1+j4GvFYGcu7uh25d0x2CdrLP1T6
21w4mepy6KQh2ptcITI4qgXt6hIEYwnfdqQm53xXpuwzqymfLFsTqj2UYLuQhrbM
esyiN+bfu4I97YR4OjyinqXQI85mEYolwVAt5zy6jpfynjZEJwDkkVdzb5R12w1/
shebBha36MCuMnzE1fQNgwwiegCwQ8nJWda3naA35f6ezf+9tdy+V95Ahy0cmgHp
w3T6tb5hXSqzHU+XUDgWZvac8SuyGD27UZuGE/SIDRQdky++xGdxAtzkmLvHlq5W
ktauoxcCNqj8c9kZEdkkYSRcBOK4dP2VieggN6OcfhwDfdfY04fC96WJ4VV2Ppb9
zpD9KYH0lZFCOR1Un2dDzMKPopvIM52rb6a6smUI6hnwy1av2PWqPDez8Vv+/RMa
2oGOlQgUK4hDWeUBIJkdkiKEr/qRYs19ybj+aImRdtxx5+qG9WpO4WIOLNzWysG/
XcnchVyLUPTL433/mVSx2qQXOPQV8VGe51XOxceEh8TpKyso1AGi+oJPGvX8NfV8
J3ejfKWAoP6OIHyB3A3Hw5tXhwNlKIR8Q6NauoUNY2Kc/yj6QGPiuH2x3YZwnr/k
i1sjeIW8Z3drxUi3FdDzesC7pFYTlJeWoN4w5rWgTamH/8ClSFTmHN8+ROxj5nBl
orv3dBbWNUgKYdRltWjAEAXR0N+316+peh72xq3Yg3jSOwvH+fGFf4f4D1HyMFq3
uZE4fo9dz9zjBtCQC+YEMIwkcEj9Wa7B5Z5wnGp1Y8UvcZNpsJA0kHpfu04J93WK
BQ56OSmxeK5W17tOzK3p/ns3dRS/jxe5/fuLfeEVEloR1KCoHKVARjVhHJ6/eY9N
PdCAaDHEpKpld3oAQiwZXAF+mHp8DwuDJiamp/rlCq3f/adUL1DOJBzeGxXW6FlB
4E6SmswP/7sNuTZKfqcdJGLGG9uOW8HQ7ajdW4sXH8vy0dNAulCCpPygrNyUOR36
qKX1vvgWnpxQYy0W2lNjdFSUQGBGzZUbF9L6RYWABklIfZVZNANqPNW9B7CGb7pz
Ca7J8wG5kdwiP9BgNm6GIY7fh/ahdfrMjhUCNVXEENs9g7AfnhyYTff1x1XvWRvF
JnYEYHA+JakzYqgPqceBfi8Vl5Z3WO0AP9zV3BchFdLM88nnFoC3r/e3sPMym+xH
jGFugddcEiH+159XeJqQt+3YgcKaLG4aXJx+BIp6ICfDWFSNeE9su0Eono4+ulao
zaQpRPHGj51IaHJgZTz9rB+AseVMgO3/AkJvac5VrwYDWzzKmM4xmXb+eX7jBwsI
qV82xuwDpAigw6YetJcpl4Nw7jX3SecUTGp1h9vWWIOxhPREO2EwI7zdI8nhNgst
YMZ0haTwjyc64VmexWZZjUqBFc3bNLcordzyy/EjfVb5KRJ/SsNLWWligrMnT/jJ
1CKUP2OKze9Rhw1voqIUE5rubhy1sc7lOdO3r5Z4rfXud9hv09Rb7aYVjpiqdJkL
7yiYK6eKS2lr1zytMH0bdFJIqc47ktUzjYhpaNN07gFCB0c9kM/zgEEiy/3vtL20
Uj+88kAS16kJqd7vkr3hoSUmCcVyPF49RPe50lUXYOj4A5S3UlRRA1A5P9po+SQx
mQR8gxTsSi8s88qXyJL6rDBHJXnUUOJ4Y1Qp2aFKwJZPqog82yLS2ateIWld2rvk
f83RlRLVf0XfjkGdCj4yHR26hz5vhkBVhjVF+Pd2Di5hCnI7X0ZmF6lC+lDYwqOo
UuspqFwJCmq/4QL2ealwzefZr5qqkFxGfH+UhymdHrgEnvrQfqWl3bbRJ86eM5qC
nVUy9HOk30PsK+qmTEmyHsxaWIOdTDG2jQlYHIFQaS72xKkzQJuy6r6qeUPvUYcd
bt6kleuDpa+x4QMdNFriDDoo5zVvyNuPSq6xNW2E+yzsTv3Sv5GcuI3u0qKtGfMk
s0vnh7UNezxUn5Etr0MGcqUDmpb2xlcdTSzQAeQertC/VsUkVYN4pXMZBrUE1lzL
aYJJXYN9olaPvtDN6BTYGg5fVODmv1mD1zDkGA/6bzuWf8ix2kWzJbxeoXqPp7iU
1MXz6vD9aM0Hmq31PYl2nFlmFcETSFuiBIZKuc68fEjit20Z9HfnUk3Nszmj9i8p
TN4KDjOL0OSYtmDixVcTukLh4+UciZhCpd0sEjKXBJ2yu1bKeyiFGQpIOf87rryX
omTn3ch5OK/pYhEQUncDgMtHNVaY7f9sN87dT/gFHjQjIhv6ozLkPh2Eu1XcJzdH
He6WGtBpAzINbjs25TqguXkVncQl4+NiCivXrcpI+q/VvwP3hj4Wi97QGu+yVJza
UT4SkW08jJCspZ3iEdfKRVKAD6wjbjsgBzYFb0UTVbb2fQiWOUjxViKGv1l7jNK/
ocBo78Xva3Z9wa5GHoPpf/7qUuNa/cKs4EdU3FImu5DZosYlO3wJt438up3AQQk0
VkdCcauPoZr93+jdutU8Df3SKeJK9TQgiTf6SgC3HDKCc840plmlKIkUSKQLUr+4
7fHW66eUojqvNTUJ1CchLtoLmmdYSYsKbrp28miyT1GBCwrQAx3Fji1sPDd6iuCe
rQ9NKMVQPiSAZQ/NfUi5AI/W8QjgboxlMGUDZsUrRT1NGYEO/OFr9zZ6i94BZB8M
xUGWiH7KWjBVJ8FEGm44Nch3/nXewQkB+Vh8kG/xlaStkaC3eA6dBCRnn2jW8IOK
VuQPWjn0DVJKyZ/ICYNwx1V3dMKQyi6LcTnUDoy2V3f3W3SQN6Htfa7P81I5zqu1
BL7GLIy03XMdEL/yoiST8sm/nG7vNqBAjv2pZc86nuuZwx7xBEGw+eoGy/FxcoZR
0ZjjTG7cRJgD+YcWgy24kNdouan6fxsjOiDJzr3uAMF02qfRrj/6aB4P/nmu7UHN
OdsCz1jl5Kq2+s3283K7p9y0Zp1CdanXkoQa+0fOs1OHr598sMnUIdnFL0NMftGz
MT9Nxo6nFMb25ZL0/TpcOQ8Fp0xhOJotznFxrNTLnEqQ4o472nmg8q0W7WNd+E8l
DxV0HwgRKjqNqtDCmXKRXeRgVzvgjzGEGxdHIGHutthi4tLvrKWTnXiqt4ULBVD6
MdhTysHnuSHZTeumUF/OAFruZIjPHdtAHxtLXlIxoSuvma3iYQJmA7JM87T3HNwy
fpJl2O7Rw8YKR81bX1tePCxDBr8Km1yYYgCJEUSsrnbGTDmAOalYOGnaG0bUo5Rx
Xnv5gzZeRNL1aE9haGQ5Y2n+BwsGWqFux3gC/P24hOIh7zxGrG+2A3z2j0xBJC76
krMRITVrbBYiB8gD5KPFi6+cGdc4pE0tIYQ47AvO2Q5ngeEkkbTaXMXT4lTf36NA
FN6RqAOubOHelLe5J1577UpPVnmzVmTsS3czKWz/9OOUwQzIW7brQq6UChxrHMgN
IQU8hmR/o0s/SQPnYVAqeJNEqOW4DfY9rrgnD12TXUcC3eLWF7g94lwZKzFsCaZu
XyP5Ets6Z+uJAXHzWMPv9IwlW81NaFr6myWDCdKbjx6JXiqmXr4Njq9BTaYVEwe/
2wUfJPejDxpIrrenDATI1JrW0tetwyX5WnViM2604c6BpIu7n1fELlaOhnHlZRBV
QcLZ3JHZ4MY2tTjpVxQZdDz7kbhiNmXEs6lf8MxwNoIRIP/zNn5KD9jsp4JYfGmx
d/yOGSCCXd5NMHMn6pOz/ixjGXaSsRywAO/VD+ZIc9GNz82wnTTFpG+wUBwZgTg0
0/YfsvGNrVs/6ncKA0iSWKFkawVLBHv8SaJ6JnlCmnglt+6DH1cudOpq5RngfqHX
1K34hdzYttyOS46pPQAsbCQvbmM4Do2kQBsyiKl9wlfDGPr7eZ+z3AWV8Y+QWaom
u/YcbLIBuf0Xxd/gr1X1QG+TvmcxQmtprgoPi5toOvcysXHsSi/HxLXaGHOJn7K6
pPUI5dGwWT1ax1kxtSNvVHVYjaYRyzkOVu/ZZ5s/bIQ6BuwaLfZu20TVOatDUaPY
u2jwz4mzRnJZVlXO7JXUAQCjnUPqhBX2GiG9a1sbL/ukmZvlRpF6eGPL3GdCes3d
tlh3yDo5U7po29lF5AJvFqAlzIq3/ChTsF7tc3Cu/+rKsnRz74i9aTxfTPo5rlDe
TZq/kR6uGyKa3GX9eWnGEOdJnwQGsgMYUpZFSQFJfys60BaXD1NqnzsY+1lQAPTF
mhsPbVbXGs8NlueEm/qAEb9PeHCEvdHH0ggaQcrK6fy/bFdOBk0OlOaew23rbLCI
obZ7fsonfLXIzzOXiuc/qbX6uTsUMwFRs6mkBxI/U2db8GIVGEbsAKhaLY3evxBm
V1dlxAENLXCRQw2Y/20jAHlL4LGAfjUcH7WlHPzsSboxgPx4UYQPqMxEBLFhTEDu
UXMmgDkm/4xr50dDjUMpjKbD+7RhhcBL7xzgLjdJMSSAoOI+LHLAfJgaKSejiZ6h
SIwWt6kagbHHbG5cmncGow7De6jVMBGyb/KkJa9kXJqRBoJ2bktxHlTbmjQVHMgY
T8TwXy1tqY85KtAdUhTRBThGWVTCWoJdkYt+yGFhifhdXsFO53mhOYYYfFKFXbY0
qgRLLLyQSBj0h9GzJmr6So1N68tRSXf+vYJVBSmwead3J1BWNLTcB4pCHaA4ZyYX
ITR/U3ssI2AtqSCkmeJPhUCYgUyPMxueKuM90Qg0/PlCSuR5uy14h9GEAdSjfeRc
FH3EPAFEku+zKYQLB97A1VnvkiN3eqX7egGfn8P6Eq3lDf9OI/xCNCA2sJwr2fh3
dYjXqnKkGePhZzYaid4OYapPCeUoHXv8UNFuLdWCNWyiP2dxXWFJhWNZ47hgkEIb
j2lrsMqTrfj2rof2ppCAt3RU0Te7fkBLybFz76uBHP8uDFxuf7bVmN2jcqy/xOE2
WYNfoaTwINr09fejc1dwuwL//9ii+ZRVKSMs/uSnEG7pKCmDSKfGZsbfQGO9nR1v
l1WJtTk1044yjDwzWzw4FVSeJl0ywr4UIOBJfUJruepgQdS17fixtxzzf8xHz4Kj
xggLJSr2LUVBHE4FthFFSMt6xYe8BEPoKFonAd+t4R7hOmpdAciHWrZld1/Q+E3D
EASfx9ecBvePKbDVNlUILYTweFhUX6IF/3ofVostssPWYN4g1BfpFq61Rs0ZaeFC
qDUQ5lIanlNtoSEJdzL0o51S4J1FEKLeUcUUOhT01+ZxyPFpvOysh3BCgezuquD9
IYJQyAy67tXnFOJDZuXljcd1dqEMZWNtFDkaFb07IAqNYv+l3knL8xLrK4sUDs7W
ZfSJgt7r4+JsnnE94a1CMSo5pKnECCZLwV8qL1pTGlyQ8szSaxHFn8RvyPCtS8Js
Xtr9/Y1eBliaWPoY506EKlKnPxVaO3sIhdsyMeXGdcZWDUZnSd8xC4tGhwTHSCBV
QOh9auvlrCFXjEiNFrafPCDVNKiIsej6ikSIfYoa/DOG5j7YQx+HzIr3fu/Wb01j
1WcFcEPdqYZxJ1vLU9KciwQKwAdcqhmBHFJJLFvmCR9WjPNlFkknT+HNkenq/NSD
JRVj5Pikdtuf5qv+SpRKIAw0b63GMbqmlStjjB+JPebJaDfHqEtY2C7WKn5i+ueM
7ZlVd+6WCq+NBtO0LHvFNOapljjEdap6y+pbWyA48fMtfb0pwbYtn7NDyP7vtFho
GzgDCL+ZhNJF8ek305fVd8aVbAmSLjboy0+Oo2Mdf7Kc+YzMKsf+fIUsXkzn2iUC
UKxEE4twRxFWjNmEoaZHcJAvnP9mLy6GmWkGtpnbXp5dqkhEKbgyR2BlIcGBxspu
OMcOqTsVVltJrEewkCqA6SS4Mf4hn6QRWuNqccAIFWz9LbxWkGGFyg92zpWqB80W
zyD1RzzN1kEtALrRE7jyfkEX2HNIBRc58p89GnA3AFlk05fNo2G7WN6eXErTcr3o
gZHPWyLdMJGU3OACVipj6m170vwncjaUvzL4DBSq9ASpSiZYuZws2YnNlnQSihGf
iAUPEbTCQj55GhAK7Kgo5AjwJH49BjVuZW5cGEQRh7mvUsi+RfTafOfqIBLNWFLt
wQiMpr16RLfub8nscZryuGqV0FdO5b/+tyXFIlws6A7SalajfX2yyql84YBNYtv3
dqF5gg3Og5u4QbuVkBGvFkw7Qk/TMZOu5z6UaBu0Rfb0bEbvdAqsYAO3EVkvEoKR
JypOzeacVHAWegEfp1RRmOjwb85dKu/7uJRXd+rLTYyDLQDeNHukWXuEmEAeQeMK
3r/P1nJ6n1hf8cPd1T1uBAY0e/UiNsAu4UrRJnVck0EVWvlTLKZRKFVVGLnBXxwK
ar0ywZUs84/FLlnPgEMCD/845fu4uF1qkWeh1aSdpbCJDqvK76txpRnDhj1JCAgl
XZ0XNChrAneA7GMgVByS5jMIzMYzYmKe3BSl0O0eeJ1Rai5qrEjBKkWT5Rr8fxG2
jKgwT7NpQo0SynNiZBmPGW8pzcZU57R4JJlpr3CRsh8mb5HCBqw9cUXAvHCTCbAw
lLl0CzoacGygCOACQT8AZUO2IeCuMXALfD++h2y/JkwTsf3BevHis1tGsFQSWyx4
UGy5tZcXximHztDtvwkK1WV5CsRgqdn9Xn1XwSRzOkfw6O35xf8wXrY7sRZAh2gW
PukwfyDN37kYx5Fs7MU9O0bjIXyakhKyP4My9072kVNdYvPrY6n2+Q2q+/MN0ZJE
UDSbDfQ82lj6a8j0SDgCKma5B5uXtdXWhHWTbK+PB0snDBa+nam8uPGFPpO+POPJ
eNZ2P3z84wSU0AEFyZ68j5UESn8nKKzHSh4T3AqdWukH1F4F8IQu2AjczKkBG7NY
wYuu++qpMuaww7cHZ7nFEpHjet9XvPALO3TCTDJnmxXW+q390Tb7+jwCZ4vk3Nn8
cNJBMPGtubmbU/oUArLW8uUCtbSj/JawcckflFV0FKJJy3gHxKiEOpOg2Fmy+GA/
meqiOpITQVSU6idrKlTJbD15hdfs8fWNYbjcZ3Fi4fXKSub7uhdKyRZ/EFNpb6y4
f4trqhGp1uyGOyq91fJKBCJLI/xJ+n4jjQVj/k3N7mnkemb4efb6oAhhlE79TNlr
mNKQoWskbrbUR9k9e+kpRoFmo4tk3c+97qAfyZMDz/pxhKnlTsI6YHEiTt6Gs9ng
kVegux+IsSDXQHPAETXpGYFOpAGF4rc0DwqncjPo4cnxy7AqEf+VCJhAJBE8rKnt
r1CBbQ9VHb+TQyzzQJdMW3jIGeqCTNjhJ1EKXETIYtlaI2cqBIDpo0h36LD8Dszs
63NLFaZMLtzcYOsc3HF3fNEWK0wQt5p/hTPQiLonHeRkM9679X9MjXD7PPdGxCwv
gI/vW5I8fGgqVtrJlPCvk/5+FkEzytYUXa0yKturMpi3dZjxfPj1pEqwgmHuLQRx
40Y/Rj/md4FAcu7y811t2ri9pIqE3T/4TpS6IX1TIHj1yHNqKO8PxBzLwoxCbkyW
7zySMkEMa+c6OD0I5Y7ada5S+qeAs0TnUuFevusapmSQCceDf1OGNaWTllpF4mTQ
ifmfbNKhx8ix+MF05dPLdfYxLwifqdywkQ+vHd05L09zvmpdxKfhzP2X9QNLUXLd
bn94kiA3wZEBcq6jdViijiYwsSGG8I+oZBWNXof9km+fVS1rS4b40x3RkUidqNby
+Yy9MR0+VH8d2E5/eeRBLyI2UCnQtCw8aUssW3l/VKvK4Me26U687y1uhhO5u2mp
Dz6/0WfXyF/JOjyw/AvDBRgyJkbMoRcnGBOFXSvrrsFgMSf+5q0rBjxX/e38uxd+
xT3FTM3PNCXT9YEQPR8z5EGrodqRYAaSWizTUHJgLdkP+8rY+duN1LvhYD+FCvE1
jztfsW8TrS6ptnAl/tpHM75zlr9Tx///XML1jTL+fFwAWcUOU2p5xLhsHlCqgnh1
M7rb2dW7oAlFSXjAfKaP0ukF+liBLRBXJ373RbG5bN8GyZRHzxBqaXtBejKs5Hr4
BMa7dkFsNmIB0jJceRclgzSjxjLu6hQyvYa/H5UVZ8HCz+WSiTPlDwaGhyw9pTYI
GQEb/g/FcbKgt9HZF3w5yGMJtmq8e03RwgEdLUdeuOzAPpb67OgEQgygP6cxL3JF
ksqJaRWk12eqvDAdgcW2Qz2AxMGLG4SuNP7m8Gv9wG48tOjEkEen/6U+p/wlj0cZ
nw7GbSVGTCIzpotsn8wkfz70Pg6xr4SVYvIEEATLK2p1pghPy1unMsd/fuiBfC+V
TRbdMDYec0ejCZqffoEWyFHGI5QB8FJXR+H7C2TqKZLnTsiO1XCTgDuUtFfaGP69
uPDNp6Et7Ee+PA+ccCZFZwgj0ry0HOUw+ToHZkXkK/lZdM2ivgo8cGwAIutXpzHc
TlaY43cPqNS3uNWBthS05pQO7HheSuVDhvbDABjYx5BZbGbhiL6FLp5Spp4EHQK3
00vrUJI2YDLkHISaoJ9JMLt0KKNeI4y+51WEQ5pXtmrKmdcUFNqAjX8w5xMTL2xw
8mJ3yUmUsVaH5Uoj6+inU0GPpFnpWbm4KMf8SPtaNujn74mdb+Vg8KbAIoCL4XDp
QsmgWTVPEd7c3hWFr1pGPVC7T1bt7REE0T1Mi/lTsgIQ9VhU6yUkxuG5pGv0TSGC
zMO4c84WpMe3kOFdbUw7zTKBx6WnBZlyjsgNy7+OEr9nl3GbPIcA0I31ltxmSoYg
7EE7Uehb0fPfz7RYgmvbPvvnzh4Zt41+3Tt7ZTQeiE8XBiLvIIwABiv+4J1x2bcD
m44rsHvFIjsQAa4jRXOcTtP1QGlj7IAcYEKD2+RjqmU9R9JDlsGybHefc82XwwJd
uXdj3ZaKRXLshPSlos6QkXArlxsAqxu01puD5MLzD9kuqRMSVO9pxAkecnclN904
0vJlBraRZvc0AF/Di86IwnSS5ajU2Lc9WhYaKiwhOcFMb8HK/2Zqhj+GNjK+Ds/C
qTwZNaa5bCd2GKxb6sZYDrbmlKAk8gp1/0bK+Ii3K9+a/ZG/PK+HVEaoIotVJPHE
mAt9a/Bo13TPTRqpSNryCBfz6TKnNygCoLVNzjmEXUF2NA4rBVXGPl6QejLEgqzK
J+ixcnmvZbelmscdcGL2mtEfCECq6rPFUH3tihhqCYRg7+YHTqXw1RqrvojQbZ7q
9Gf+vAXSYa5zo6AssMg+nFySAvFgvCWrgSiJ5QOA5oeG0OhUdLFYjen9Waekw/iN
d2uViAy10AAfXnEIkP59F6i7MasOPH61UVgYMGlv48TidSagB9yq0eFgBAyuuFU6
vWgmc7IkhBJF/k/DNQj5qv6qsbOrLd0aK4mDj5wTxRkl1wL1NbKOFcaDmw07TgjJ
619sZrEnepcbQqGdCFNolwFjbwZ0GONTkPgSH1FVnO7RyeccHanPQ5rl+GVexh+z
XKsGe7HLNzCtaOXtofvdNGxNTkqaZal+9xEw0h5r1bAv7hcdDOpfVUCAkVKu1ehX
6cplIk3QiGPKGAZTN/WDlLmykHzXynSKHpUtXtSjtC+E/ZpA2cJM727/p+JHY+9N
I4cU5u4cT6f0ndw/A7TrXSUeNseX+vYGf5BzQ2loRUxGYsFmflgkcURSyWJXV4lS
P9zyqTuZwl0EyqrcvjHK4PA576DAIoNTpYQbB4+Nh/jpVhovhEJMsqkaf/SKccYJ
Foy9wwMM7T03WrpNIJ34kun5RpiYfH7s4uan9WSkuumx10AMFG6VRGhgOoUJXqau
tvqnwn2fNpELBEO/7d9r4rUeLMvx5du7AFbMMI84JmA+kZqRGygsp8twMNNlx9FL
4ivlSdWchGnXc/EOFlm5lpPYZVW/LEpoBW1P94TnZV4DBqV/Z6KkXWaep1ucv8fn
oFKJsVxHn9fH6ltf+ZE+uZVqGHVrnwqsdT0OEkp9Dozd22FQ2GUg+u4rs2LnZgSv
x2Fd1RfpXPSM3KLNT6qv3k2/4olpiNo2bqc2d0brQl1fvdAriNttRIVS7fdMOvMU
O+RLj3tpM972OAtmNHbOdqhvs5dUVQJtPIjOv13MukQGrQ0QaMoNXHQNQvYfHAHe
kfSAcZPpLixXb5V0b9ajGyE69p2m781xJ5TGeZY8AYtzc2RG4+fH0XA/BJn+bLU8
K6/Bva2YGAlkuCT0B5zIg+qKsFJhbwt2nyVdQ9AUhviLJhuhiiKLp9GnzLiaCoB4
kIJl/yXAM5+As2WCuxyIy3lK/YLrjbqPVAVJmDvj/vwzprtipsJYRiBA3F2b6w51
1bdwjIhRuhMnxaPLgmmwEi8fK7PqQ6xM7+zEZExRFiggIiub+iLlgTvQJ6GIUqMI
PF1IJR4Oa91Y+E/c+9wMUscFk9pOMmuQbN0QR35I6LtXIPVgfxjymFqHo67u9oV3
QpnK0nLBabn8Kw+2LB1VDIoHAnpRQ8WZNJE+ueqPrIG4zzD/Ab9aIRk0v9A/cDBI
wN64id63eDptNa+D27T6JfTHf2exhieOBVzNNBiwJ578ycE9l9IT2H/dnGXmGfWc
c4JphAZd/j46sRF+fj2qHKC+Wr19nkI2cZ5GWuWQFhqN+5VW/8hCzyt1EXN44HT5
JkEv0flZrBfF+AKT7gVrSM5tnqz7DBsEgW1xx8AEZ+q093gXMlr5LLFUhxNIpZVF
7fZwkEHBfENCrNGgKCxMen8sE05w7y+dkE/cQkujyNKDm5FJ2OSCnSAXeStgwgJN
HulK4qVTz7U+niThs6ANBQnKBLHNbFSkqxAUJ+kvV3WF+UjUXLhiL/MXxO9rYD24
ZMTu+wCFOBXR5XnqPgGICM02SH6snf4oy2SNrEX6NUxmpoNH+PpglqeT9UFW87Q2
VkojRlTmnAZukM7kM5jScLfWv/s9gdEUf1wYHUbidWS2O/YmVX+cFpSIfER46VsD
wEoaIs5FTIAD8KBubyzphbRJL6veaG8DDrVh3HPP2Mm/71JpGkLdCFA66YfSi2qt
0PvPdvdInBA61tuuWXwT0NlsQSQK8Zt/FMZTkdo89reLaBADeUF/8hB9YxjGHtHn
R0gGRB+kCBgOAf1BMLd1KJfREZRVmTJOLu3VjDOw/2DdxcNgbkcQMXDDEPWN9tm1
RNGVy2qr0mZhEAYSqsy8VI1cJ2C5TC1b/qof92mTXLaake6npIu7WXKCbZcUQ+OQ
MRP+inEuhe27Y8iiSJYjbNnz61dFdbppAl2aFMa5sUIcVDEO3f/e6lb+O9LWa/0O
payis0rtB4z07+VAE8n4NFYWvTRVs0i17obp2MXfaveNwaSMveUwdxza19W4RhnB
08kl/NVp0PW50y+GyOIBshyyGzi9GqSCAo0qX1YZOdYQs+bs7dK+pVXEQBG97vG7
PKX+t8tBX/iLhcUCtRmGkQgv1Xks5UkD6TCJM1V196ipLRkrAruPpmTc8eKLKC8/
CLSNMCTGXkLqdEha9B8k35fJs4o+Z0fIwEdB4ubmbiR3PDoP47c7ye0Yxk2svgvb
BqiHQ79yoGmEf8nZT/+HDTuJ0npMCTZf4Cr6+lW18QgOKRWgr8qc6zugZVNdd/uX
9WGEdyukiSwbFtLNW08PbghDr5hOwiws8Su+blCG1uAfw8iDVKVAFNMt6ol+YsxD
gt3QUCUkIL4dnElUkt4XU4PG6CIgcihLqJfY6oaAvEGVZvOz1vB3F1An140K/sU+
RPbJQuF9IVYhMMhCkVZ8EqInozKo2ikuKacUjgAIFmQa7Ori9USgzf5krBRdY/7E
VBnvu7Dhzt9RQReE9cBNlLgWEtr8in63hLeF8Bel0iJioiB8livto0sDe0BALlPs
CcvmhCM52YIIn2nK2rQKqZl/iXYdj3FeuP020dDuKt8+MSgoV+rVOHP3+2gHVEwW
+1ZzRAtL/nnAvQvrcnNR0DUWDR7bdffyHFL4AndGe12+x/2pSoLTIHmlX4XvAcxF
n+dz4d0u8HVc7xjPNZhPtkadBvviSDrWIcOrfej6fT5QGrA/HkCwpGhlzlgxNKSt
0L7eLaAZfb120KDLRJRt48Q4i+/2VoVYpUQQH3ytvVv9lWVWNo8LV34LARJqdU8b
nZkNhjcXK7q2wXD2qzwfEW0XCLbhrRsZM3bg2ZCKdi9eN4TojoWsBR3PS1kq3L33
lvH3+2/qdKfIjb50NVizBfZ+hYxJAuCvV4qOIxP33wGdjDg8sZzQYiNfcSc1bWxk
nIsQrsRwhG+Rj7s79F/TjcqmZNs4XcdDxGc3OQSYvOReVzumj2WLB4MyYrtUG2RP
yLAPf3Ha3HDqdkm9TeLer/OQ7oPTc64c3CuHjeSKPQzERBgVp3K/lIkvvEsKLiuQ
olrkLbhTEGxGEWj+yd+nOlupZBDiOwbqSyXFXXFKWf+zb8FQFvwbbLis10WsP9s/
3KV3MbTCVWRKcNXLnJOuqjUHeRiN3nLhH4Fu/k6jUchEzinBTIKvpqwEh6tScfvF
fpnM7CTvNY7j7wFVsQZpv3PQoIiY5kxocmh6BuTu0E+16h+wCAGqSpJ2B7bCf4xX
ap7e/gXiSMMV7kZrjgtu6vY6oUQnfk254cAh1X+Db/KuPpLRS6WwoUdB1FjcXuBL
9N8PVducjrO08pJMeKlrmhaNbhenDJCeuCd5xH1NGYUd+D/4cWc+L/2qZ/oQwRCf
U/j64fLBs6HO1TE+s9Tsr/s4aWDN5ziRoMBjK5Mbk42JOtJlqBwN5CU2oJwzZjlc
J86Dbk8l2d/0LeXJNzfHX/A0N3XR0NbT3EvZUaP7mqrX3xK7N9Q4l/PmxIdslrJl
8hBVV6Wk+Rbh4LRaw5cnwGq1BZl05augNTrck5o9KEi5D7+Ttl6ClGS9OMxgjL+N
IQooQzmpzvQWHrqqb2NXnGin3q3vMvBNZBgRZnXSRiPT/7deRCL3t8hA3YGpukpT
ypCAnpzZ/Vo7I5420KaGcC3YZTvY24f21R8al5V7fAct6GmmcaTn7rLpbgBmm4sB
PBmUyqbxuYWz9GqE4cCI+y45nwuSIEPDGi1caPM1f8Mm9SEkgxjXkvH98N+r/nhf
YMA9r2oH3PsLq9L8jBLS6fUsXt/ajoNdbu+MjLoHA7hO5ZQyEfBx8BbX1S/5NUjY
mM5Rx/DGKZ3qs2V0YBy1quQyf/QvKe+VPA5pJpbKZiFm3Qm2vWfuHD6GspefHN5W
Hto01OWXHH7m3vAePdgynm8bZlwfRv9dG0Pg/WllXl4/HMyQQB9zAFbox2zQc8cU
MeeD0pPC1oM5OnyRr9eSoWoZQD3ttlirgXPBThvvE7RbgkVtNPH2nmE90eOknml6
x3TJ7YfUXwcC88l8MYOqo+R9ZWIAiE+j3nClzGmq9X1NM2AdVnjOTQyRUNl4VBrx
oq7zvMkYC9HRd+Xph7ah8HyFI5J6zmUL52TRuRFc3sk1Okvy6TjmAnfQw8bkqE44
6p0LmIY5jp0uC4inlnsLTes1FhqS3ngg4vlUsXNzSUrB/f6FTlcawsuMS9WFkCtp
2ycwIo8B87S0JEg0z57FYLOMmG+WxIzuMYkiaBCv6lkLxX2OXP0UdzMbzC5Odv0N
lnmXEVJesWALnMxFI06BsosAmp/LqQFJUGfgI5iuK7EbchKvW2yGY4Nl1Mk8K5C+
MnoIQFNbmsDdf1FUNr6+nALQ1nRqaBas+ADKwm/8MGAbX0fO1YNEPAQd8+sQLUnI
oqgbR4prbU3pHmhPNbZoFK2R0OfjFQSe99aFB4BgHBOjtUJoeKNyHzNASNzaTer7
d2OpMGCwHVPW3IvybIj5oTUJexaMNYElDgjnUtdcx/kmtojQtn9Uv8y0pZntDhNN
YQVZeLt0F+NPIB3po5nkKDdYVHtFj2Cd8CWjmH5pV9xTNMDMMoOGIrEEuP4ufTyl
dH03ikX6VLdWEFWXuUv/X3/9YNcPjTz4GVqFL8JKEHiK+DJqa4Ys5aljDrT+I8I0
UnENzF0nb/RbzI291Gd5DEttcMgOeh5yKACe4HQF3O9Co4dOFNFaJpJQ36JtJTbt
/u/gcrM7Aj6luxLnAM7NKdWwMzj9lySFXP+CFY2vmX3mey6h++ZukuaeN6tHP+ET
FF3/jXq5kGVenbFQgh1WdvWon4LKrwPDoxL5bR1GlT1WpNUFQMPI3Ae0zt0Hvh/L
/9F07N6NHKzo2/FCaoiobOssHHWYh5D6bvXQI1EpEV8GSv0V4ufKym7ifqo34wNt
LQcY72zs8iwPfDJlpo8ahzdyVA0T95CGCF+pYGvJ8YONEIwRJC88CM5iw7S45lWV
WAz8NXgNYTK2dpJdLenDHg2hTdvrYymYQ7/2v9ER+XpxK20+thfTGNWz6ePB47e4
0oSUZdeKHQy7texa0GqUkAXMwM76p/moV6NLWJoCIGR7PoXO50qO2vXHeBXwHor1
aLc2VDbIutdnstge/uhS/VlawEVt8tqxh8Ch5/LNfUsSZko6h7J3LJMWilyD56HL
+yBH1oJBmFbOBezidVaRV1BPTmSnfwce9blf+KHGE6b3yUluVSo9lXLXshEjy3O3
xQFpGdCinAbVK8ni9pz+eY6drB6n9bBK/alnptkPdVhtL3S9V/jZcP0ZXOSM+tvN
RgPg9qZtB+tLGbdsu4eL5V2FpVTeHczUfmScpSLK0VGGCyJSP4guxAf8x9BxabZp
EzWQy4VQSBduocLdPmIB3pi6/AeU6jMCRXFOrKzvLzoxCADSwEIhQR0QfexUW5Tw
hJ1Lix0KCUi7aFaq2NpqR4mH/ZyhaaCMuALcTX+9yVlMGnCTzmcG/vACQvXkvSa6
88TEkuP6wfM+t3lVsmg9XOVD3qkwH2J7RnTv8beiPOSgPkcAp0g0oGkJeooR0X3e
W5pgLEVnKr/IlUaNmrJYgEo1Mnp9Uw+r2/eSHgxT59hWJ047b6I7qrFATZMczNF8
Mu09v/BQbDNu5bonG6G40XqWV55EZCTxKJy3T013eXIHb2SLRjDUcQlnsnPdLB5v
Tp4nHBT5lLMjPB2Sp3uwVrn5JE6DXycs6sR9Pc1sC4AEMHBF7LKH1YGjreMuGt1a
CmNek7KSIrCzhgladBA78unflwpySYbkpu7ueWUjuyXKWrCQcpJ2AV31R+id706C
5DWH1rJZw9cafark4fxDZwB/zxAFUEn5bhDPYZD9yA45jzPBZ0FnafNCXNpD9oxM
w018hhI7nfeMoHiqFhac5q29E1bo9Vyl29B/XCpHHO8dyaO6oOGMY0nDrE/obW+e
TuN4Fa6g8T5iVhIUi1JGan+ZPf+lq+6FkLOxEPGYld6Hv6d4yTqVRd2UtHuFcA1u
jpYJUfOMNGUC8JTcNEV4JOlaZrn0EvGKw9gLzSWie/RcEoqox2//UU4xI3ebFOwV
XVFMYsMHpCuqeg4ojyQlpWcDqtuI8Mq3Bv9Az6eO3B0JbIjGB6AR4PZt90nGKhI8
9GqEoVAfWp7kpKCQt4Uk/fhxEJ8bqF0LGmtslUEzTHwyBleZZ7cuQ1Ud8AG+y5ts
Lm0zDx2XboAxWt4iKR3iwtdY7CzMRwKA8msLgjTNt05TSZyV3uvGDp+rMsEP3dV5
ls44ECxnpjirAc1Czx+776HlHKYoJaHMCaDe4wJQR7YId+WLBoIZIlFKLQ6CqnNZ
7D90ywuaiKhFNLQ4mF249fmzJCFYrk0oelxlPBNni3RFMktIsptJsn3To4YDiU6p
GMHXdh0/P30f+9R5ci/qe27XQtzkw9gRD239pPpChXQDOfOt77Q/DAv5+NkMGoT9
3vP9ahdrWbF6MlGCNGNn4I82JXV0oR3fn94Qbv0E6zLaNXOt1qH1h2E7g2p/BDay
4+95EL1tpAOwHxsQVtswQVEdZay+txYG6ZRqeVjCIZsGDaY1mMtP1vmYXvkNdIMO
CSxfEwD9vpuQOYK4EzBde/WhoFpPt2o0PMANJqSCf02PjsXWi3dmP5xocNYyzPIO
If8O5/0W6HcrKD6epTDNW+xoLDE4eZNEpbXWyQa+oBSIJiHFneuIVgxHFmu/3qY1
mRCLhHUWNUcJwu87lFcDv4+uBTTYwMEz2ntgUSs9dbaflgmsaF2c60VQXGF/xBXg
UmEXr9Xyiekyckw/OyMHST3/lbVzvllBi85hUArFFaWIiRtvSsp1QHMd8O1spal6
qzRdMJ0WNVw+mtIRfmW0hlht989cmYgwIOmE0e/Aq+thAebUhIj6WGXKOYTNHJ16
0eGuBr5n1PzQJCwtTQWMdTbBNVEHTOotapM03Pfhd8GOTHRBfblzWbYNVw818Ypf
jmpbB8li3JDPhKUW84z/ZDBTa7o177X07WcLCIpzXvCq9MC3yG00Zjbp2lx2CqUN
68T7zXUn7/8V+HrC/ElvIcW5wGk4Zras/sDIikqxlq577n438PK0xUSvm5Q6q7oL
XpjwupQpCAP4U/J10MR5JgZd1bm2w4pZwAXVEztwY1JT3O1Hodq2wOKEKNPTMeim
FskoV5GfYDRVEZSvaZUH3/oatReX53/8VIdOuc3JVXGiFknQnYjktfmYu5J2choo
9W7MLOzbihEYCMLBrt+zeReWi6i27NmqJFKa2faCED/d2tOJK27JjXF/YS9gydFN
vp5LEYlWhbkYVjOZzjPFdLLJFeq+XsCnulPBwrO3Zk29lFPwCdok0RbvFlLHaxut
nwWkvxQExihd6omKGxAleUSqgdsfGlEpphKQSRfuUM5T8Nky5bcyCA59Xn9Ebpdf
6UhiraduTpRctB+ucOPxCK3NdWyc3dphAQa6GvnHW7bDZu5LaFkRvJsmAD7tEuZT
9d8BIFFBJEwFVd+aVy//GsTLIliA4LvPSGgHt4mc+ZnIi+Ver1AcgXxDqXQIeCp2
2fxdUfbc4EFh4VCmrjQPUAPVM6fCEPMmX3ayE86/7iLQmyQTwBU02d+j4FBqyIzY
4v5p5gcLIAxyWnfyr4nV6yYUxN16ummYLjnjNuPxyju+ekajQNbur/oaYoSKxxoQ
K2uaqwwHllKYukONZ3oszkRLuRatYtKc60R1YuJx4vnZjsCgDS9+zTigwuZS2oeC
UDW4JxwhalqC8X3U845hsNNeorn7Bhb21eYxRu523EwzimUucXUMB9bx6RzoQvBp
Dm9aLOincvv8ojtfVSxhX+naZPy2ai7nWv7HXYc1Gi4+UUlLZ2AlJmLHSgPeHtCF
rxEkx2FKDsDFFbWiVtQPsmNUr6Quf9lOQNgKmLV4ZmJVvaYNrrkoQWSiHDMOH5Mv
JDV0V7ZYGYLnxxkp8YBmU/5lFSd8ce/aNvi+uu4HVsf0SdbDP7uQ18sIr017pKSF
jVslwzN+THqNIt+esnDaGW5M3laxj77p12nsLTnevaY7LAYprohV0AExQwslUBfJ
YYdn9ifOlzI9wBheWxxdZL9Ojd9QylveYNAI9GtpCoNETxj3yqi67MgtV2vhhPvh
qB2okQOCvSOJ9MaTiK9riDmU1WHGVcNUg4a6Xy5uEmfFIFCwkk8sUwiu/S3s7GXi
3g/6SuyMJwEciz1jtzp52atEOBYHcBzzRqRuaHc85Un6PHPdrQiLKId6THC+kjOO
6oMhsDmtm8zqgHRP9vhdg5oZFx9p/cC2IYvZdc/F1s0HAPBuID24ejHbbiN4H3eT
wuZi/SLjy8ESwaNeFouk4HwRvQfka6GecdxCwhgsQdw0yYGF8LWYYzywN2mzCxzq
cxrtwLHTt2zlCxwJRSqrkfGvVa8Xt4bWAVJhcXlyAqRmcft1R6TlM0YeCD8bC1cG
iK8k7UHhCjv7s7mWzuO7T6ebBkLe+rQkZWq213ZvY4kNtUeIfom6W5mUppQnfH6H
tji1tizS5rnl8LdUPvHNSEdBboTuWCYfyP9e3cSn8fxz7TzpT8rojoryhQFsbCjz
qjax5boxHzRhGXltEQItfp4ojGjYItroiTsGKO/FoZxSRfL9Y8+xbwz2IkhrDezr
1p1U+C226L1TxgD0ZiVIHdbjD9ir5T+IJSQ/l9P57m8u6gwy/oJMG+xDLXlt4kGz
TXaYyrNnqPFaDTJlz0ZIvS3RxsY+ASDEmxDPoMzWuUGmyNtWq+kYNzKNZsmhiOBE
OivwpYsgPJqCg45mTvalUdNPhTl1b/Eta9Uoh1/tvlY/VdNMUxLA5M/5p15TfR5l
YfiT80ZmoKp/5REMCDfYZ+y55V4bW10VcJWVfayOcVY+MlBuLmpkJA5UY9QNPFF1
PAu9g/qvoKG1k5R0dCztHi2hX4unYBVrd8zjjUexsv8ynZszGi77Iv26z7X24xas
DrTLWZEaZ5BtqUf/LTIANOIxyq+c1IfJHtrvcyY9cQVgLJTfvVS2PFkWJExmxfWl
OzmcZ3swllM6OG6nYRNc8GK4ifXcUXXSYLsPQ5mib8aNibsCclTnVxjqiaXr/5wz
Zp7cd4YXB/E0AYVv1O3xp8OFTWNNlbxx+UmXTTggLEfEu2A5sy9RAEfAkuly4eEw
kI/WCOHOYor0CPFmdGl+zOICfIw+9SvnT9xdAgaOyZZP6d4RaO2AyRZBCFd4TXqe
tHjX+zhlqQWhumV6s/8AmBtad5Dv2T4CdKKztu7S3rKELvK2p6BdRtcAyUKAMMGT
8BuB+YOW8b4/sekDPm6fGAt1voOHfKLc5P0bj8262qcE9xtmouxYATsacQSslZEf
ntPrh+vPSrbwSb0I7q/uanb3uTUvKe7MCEej0yVzR1y21ylZT6lkn+mGidocas0C
CULOsbO11ewV20Zki8RXold3v0IxsPfqfkoZIWphBCypSfvccFSZrA8rXtTElqcG
GgcZwy98+RCis4bdSZs+UE1ul51zTr8u+V/GBRgNT86/Lq+tmePna+Hr4coiGUxK
EWlXEFOjNL4P8GvA3aRBDpRBqcCCzX6na+jgcSs3iId4yO7kbm2h9OtC7Xmq/y6s
T9uFkZhR+VL1/D9zpPVpWofBFMPk2RDe3lStAgiH7o0LxIE7GdQ+AKrP5aD9zGV0
LmHCnB7bqUcahgwHeCx9A+hmIg3/JiMI9ZRaJHkn8d5vI6CV5XqlySEaTSRGJ6BZ
0io7rjCunCxwzHmpUurrLbvsvbitnsNLEaNBSoO0RGKcyT3X5OJ+8CFiGZKIUh3c
1Q+EWJNI34+QGXcjWJwRwzcZL0zXHDHqMAcON0Pyyc10BdjhYBpDyjLzdVFEo9GJ
T8nMwLNmC++C9OqCeCNYax3njRA2tnRmzMzwwlHtGcaqS0lgvl6DR+JGbVo3bXR5
d6M+Hm6G3OUuCVpGACi6Ah4xpb4gaQ+h0Aop6TqnAfMhEBXBUsdTLo68kUICFT3T
RgffSWZHFvI4kdZiwmRE3dZuZZ4iCpW70Pi0VNg3Bd1CdzSOfL8HJSue+HFqUoyN
MoKrRmsnsRNfhRvHItgNv23GaEcD/kO42XZQfQ+21iL5DsqaqCrVs/6MmLVjoCF5
jrbV6YzobxpWc2UPOfFERH3BVicD/B1hUill+aZAFbqPkXFE2D5xVA+rpKbNCfv8
qDtZewRUnJRkDjLEGvo5vYFCVnGrfWHW1Pb09kHx95PQ1tj1ISaD0gHBAmINowkc
gyFGPwdNldW9xb36VoC0mlO6h3fsXCWPCeQTIvUJgE9FbokmNWTUm4ZfTbAl2pcF
MNwaWwAExjcd+1rj9mHENJTZtwBTe98YZZpLJjrdbv1iALplhIXCUMVirYQdQFsn
9LNA+wuM+xzOMFK72oYwKgk2wvSmOXBp/5iU27A2thHJxremzs0P8zreQCIoV/ip
F+ZrjsbInvt44iQusoW4YcnVWUyOZ7IV8MPdGCj68z6D8ud0D3niLyNAyP2tiuip
3d0OXDsOnzTipRNCj2CeSzgDRHjZyAF6onjuQnj3VVfQPPmg9DPJiczeUnJs6uim
QqtW7fMCHUgn3tTb4vHwTa0842lu5k4RvH+QY8iRvxz9zM3xjirSWuF4kkZhtmbD
o+iJCYeiqjibVCvQAXzwiZJrJPJ99yvYQDUfd52X2sGsK7Bfb85A8eTQ5aHLblsm
Nf2PojRDv1OIwOff4cY1QgDQVEv0yZJPKdqXVRDJaFtamilzuiksltKb+0Y3HiGr
sHI2FXXqL/ELyKZsXtVjRwazb6vbyGb51D5EzVZI+58jQTeI2eZH171P7xfAR6rO
wUdidybsgEgdZ+Gv5iFhaZQ9fl90EShE5gKCFDBQQkudg10ss+ivcC0CwnZlskIW
VXjyyLMCLP1j5ryz9s0qtDTsYnDFP7whyp3+f5DZAuiWD4100AQLOPxDUkh4nRHD
Z5XIXgpT2nHAwZonk3IrDSUhKR0oMSQDG/xK2MF0kLCEICwxrgIwJ2n0s1o+82LF
1drd/2gZZJP8zas1D+vou8B4KLEXTiszOa0E8SJCa3QxfcV88ZRAm/z3Xrsy8ky5
tkd7+28VFp66EOKGYxleiiTFvHO0OmKd+D+MNhi6M3lqKMQv1AXuJjNBJo2baQcD
gyGIyJYmvCOuN4H8teA4Ts/QN/3bIocPD20Qmmi+JxcvP54dRpYPw8w42iGcgxvO
qtVJMsJvfJRLSGE81B6RLizDo1OV62bf1p0TkKUlRf6ituK2sqRjbKRCfiwZVSlS
mEMVGzCV30NhORon0hJNJpe+5vx1XpNFF06NEEK8FDLi7VXSuEoHtVnYpqY0aN1S
MSQs35nl8zaAnuvO+/mGYLVjhfUzEOEJ64p7CSDJmuSPsUj9WS0aDLGk+jR5Forp
kr8GKe0T3Xb/6TYUGjGu28Zzr+qylhMtTpvowWcWxeCV2uoUyxGSHkwklPu3pa7f
S/vM/1GAS1pbZdahozmxsbpUmVoykLAFZ5iP2F+PPTUN8Qoi0EjGZaX4JakFed0v
eUS2i8pHrLETlXiH8rlPvEKIRkIFEweNeJNXKOwIUkXDLN1s7oCRLkGL00Xf259i
oEJ4U2/unJqNE8TjUZfulfTOsN77L/7yNAIWWceKfR3RbgDKG6z5Efx+GOLDD4J/
wgDcvvQ/9MGN+qKVyOAwQ2hjxVXBRGXrU0PJGyoGDgsu6k4dNRTRqbAptY8Bek89
UxfEuE/NuPCmZAy43OlhZlnO40TlituSbzRxfSEXXfK0SC2/mI7o9yofp0UCCloV
D95cdR3DxDkZ0+UbKaQyrWZ0QFkE+ldi7TI4+4X1gl7xes0nWublhP5dCjr/bkrf
O0vHUOrc8nQGvgnUlc8DXKMh1IH1tjsdJpfc6iR/yOuwaizMoXlAa+2LHc1w5jtr
ASJZWBzmhz1cRaDCgBf+/ZgquDuAGQHyW43nzPxDx5Dk/yCIpW28tPwYdillSmvm
9UDKzXsQ4iPsjvLo7Iv17sjigccbqKROdiaf2q4dh0sjTroF9a2BOGpg+fk55MYJ
lCm/kim+vYZuv+ii4NwhsaWfAVD/vfnmMF5Ab65+AujpR6xjajQj8CLH7D6+Jx/w
AvLLfeiVMwY+TMi/b6VQrFEsmBfhJ7OV7sdW+wDGUkRh3dPv09qlbvXdUP+Cl6Ac
gxVjExyMBf+pzqAoT+YekOckR/hpm5gnyHGNH+wy/fbxMzkDcWccmq03qGHvCVzn
nmd6/M8bF8kUJJ0RPEf/tR35N4G8kXxmKhZnbvX2+L+vlltzyMZ8thZlqkOahk3c
WXg4EUOrHpCESAzC9tUt1URssT1zOzJ06K8JIYoXNpOUvYz7vUoC8li4Fb4QynkE
NoeGS3ekACROUW/xiULHAkLsyelUSfKQvEXLYwfhBlOe8cu+NdrtvNOEtAPMFKk2
wt79XjJExI+TnZKF165Q+nVncON/O1gBjsG4SJbVVuHhqwzatrx06VK0Bf0eXpuj
OjybM5EigEt0A33jR3uw7PrteZhifM27BhsIJfe+HsOBY1H9El6VLEYpMeb4sMzL
NPh170cqhMjrrkfJNKx8Zgz0xYEYHsfzAP7rm3tMEv+em0eLRVAvLqVHi66sqxm5
JAg6lqOKkK7Vfauj8JodFgrqyaO5xsQYhamryVABhZgcZy7phqRIUYhkEMeT+sEQ
FZKJ1KlsL3Ad6VqnlOkR18rQAzYqEPRZJY0pZUu/SVq3/GI7E7DjfJYwuG5yZh0w
4mW7KOH5z4RhxpeTQHOjkrTrMENOIirchy4PIQDgBd47Rgzf+6C6OoECw2ibwjU4
qjdYXTOcMxpy61LjEkXJjOQ5OyoIDCGM+D6BTFC0CGEF3D/YcFHdgYUngjRYxRQw
p2hrkBpJ/+VUBkOCzsH+mLSrm1oOKBMzWpG4DlGOsqg8/PiMEQbZRePDI3k/RXqK
sMs9pejDIDlrSjrZcmECPgYsuXGPS7Drxr4Nyf2VjVIhJQBatsZYmKPABJljmmUd
rcdjpmlSH3Ib/piVMaBelY2FroeUGMit3zbNxiLTEPQxJptpTEoIjbtn60rybk4f
La5wYXsJAZAXrHXNKZP/ohE+9+2q9oiS/aKIoqf5u7PYAUX9D840W1InY3zuB8F9
CHfmbMen4/g0j1pKZjPLft0IkaQMj3oT7Urj65FSx5rC+DqG+Cx0uq9eUN7DK6rc
+vYelAsWy17HDhxirpzvWu4CWQkEIktAio1w/bGi5ms3isPvncoh+CSHoqn60nPH
ztHv7SGxo+5KCooD9H36xLi5Ndgqcvyvr2xEGofbrqyuA7pahlwkEVZAZxtkfqXP
ZZKDmf8f8WwYb8skumjIYw==
`protect END_PROTECTED
