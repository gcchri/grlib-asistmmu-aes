`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fuaucHbfwofQ63DZeIW6L5vF63f7GVNWgwd+y+FoYbQaJC7p94qkX+W5kiZ9APOr
xaZNr6gAlDuU/5rOY2FFsSmJTh0yEYNY0KhOlmS3SIjxL286tVfaOkhnXwvTrrVi
TXAVUgQlw/uh5iDQ4t0rD9gcfH/6ES88w2OQdv4EwswpG1Q9DK9qyrRrpZvmLTyl
tQlApla2urx6bELaPvpSCKMxsNED9wjbCnVBRsuAQALUKSd23bfq1msP+OX+Knzs
kST/mOEQ/74TbANWIfcgTFaJsjWv4iMarecu04b4qni88hzlOrezkDmGz3dgJ5Y3
G10RuzGDKEMWoF7Mm80yhCc/pomEKsLXV3bzHe3ZabN8THdJ1NkaYsaIJm23rTNj
x07uWA3MjYEhbXJKgLGCDbW+lQvWFyPcsSpYP5mHOxU=
`protect END_PROTECTED
