`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wG667mAdHEoP5sAMBaq7mps69pJWLF3524eiIF0TpkAhkPz74EfDuupgfYeFV9xd
+zedKSWC64WiILxaSLqZHuuPuLEAMl3h+fxlYWpDjnC/JKCtSUZuAVS+W+3w6nr3
UFfC9Y83XNebU1GwTFrU9a8wTJhDCkWGU8GJccneaZj40NOjA1NYm1Wo5luPxwaW
PVxTlnSjPsTsohKOBrqEeAXWK3q3ky5U6Ck/7d1oMSZYYJqiWTCQ1VqcCffor1tb
5CB87hlCSfcJxV9JGWpVp21Ozgz96gfHN6V4zC5IOGdAslpEzjjsVKf+mv4FlvU+
NIDFV7VcfgNa12dZcvtYR9k2cuhPFI9RMZfTvV10g+9rBMdfrkyouxdjXXfLsIhG
CkWxbDPPd6uKPRdGk1Ppec0tJU4jApNgD+AYfwhCf4w12imlp0w+4+kRyGgbBiXD
QrodBcGoe8IortQljpqBtLmZnC0auY1FhU7RwKLWgnbnMrwbj+0qPdptK9S9PfPY
fkc/lrsHolBWBoKMUmYBqGcHCWL+iuLnMaS7XVldFty9/vr0lzXHb7Smgkpp0Hc1
WEjGcYGxEbn0aY09gfXk7wwlO/jsrkjlttx2w9N1p7n1potqSqruRpC0MZ4amm7S
E3HobIVuhqnLMFsdthG1VVLnlIc4K0cO1I14eM7xOhqn/d9cJa79gxStxdl++7dM
2IE6LK7EsCzGsSnaPhTyXqFg97c3LVV/vQyI6yHIJlZ0w9ZtkisiGUP7HU7PWtJT
9mArRpVRjVRyqszk9Mn9tA==
`protect END_PROTECTED
