`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcO+et3sa0I666Ft9vEajISBQfk7yg0LmpvEXghzm3mUcehgfPYjcO94zdkBTVvP
Uy9B2fLeOdnLeUnA+0+nOSqQi/21gbLK8lmIxRjxtp2XM4MlFcH8/9+KqV/yImDj
0AzG+jcUXqJC+CqxWVQqtD8JxdOCbiMWpUIcCbC18KcwwOM9fU62FAP85DerfQtE
c68EsC3tRfw0dcnTj4kJjMLVL3keQVQS1+yrpeoD0CWyC7R8CarE2OQ3FGs3YTO1
lwcVvHGpU37rLb+ELD3RK27IJu0Lv3TO5MP2wArjazmkDztYUR8Cggp+0zcl2PV0
mBe7/2nztfEZJ+/ahuS2ASRMNF92yFCd89E2ZawQGfJDSM/6G+GPbtA3DFfUpd2Z
3rDZ33R6zoX134v6PTNpC5Y/J1b8j7VuZ08/RZ3be+1fMQPweO8AELopSGKgrnxy
wD6fkNcAmj2b/ikqpyWnMyH6FY/15BRI2yr/rBcrh/JcJtmv6gRK8tVEEynHI0Jc
`protect END_PROTECTED
