`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+XIvb2+0ZsHj1IgJsE0Wx+4P5Ebd+/l+6t2LY+Bt6N/83LGB8Ju9jLuMLgzgqrKq
2gCQf7RSq9x19WsNmm5DckiFp/E3IUKTpzFU1SsPWJSjgt6MZKRqfveT+wwLRr6q
dYfBb5GPATzjd9xuDxmWdLeGAScb01u1hNCFstcS8ETl+jax3lAoEZ+LwX+yQqKz
jKeC7gXP+evpzwsB2Lj7seXeyBMCyiH3uInuYSTTBPePRiw714mUFS/KI2dxDxd9
IU4tqLa6X+pDoTG/72UZFgo7kQhpLE58c1yT+95bGwinVzerw7L0CDRR67EQjjol
cg584zPUpmCDn0WDYl6jb0t9NQs2TK7aFXYwDlOiISrmO09OlOeKk2eUf6qn5zPG
4iLQj3VZUk21h5j7Wmg4Wq10elRotbM8ulGtr3gDQn8gRcf+JGYASv4l2zl5qgoZ
YQzGIQsYTW1uZa03QtmqWUCEw19G4bjoLUtkk8nDBWpo+SjENdGxlTYmmWW/CoRv
2ZosMxhbdJc8UReMjd3IrGxQ0J9LaRz805cd/q931mPTEIeQLfuiwuPNty5lhdfY
OLRQwf4mQmj3nD8aiErwlizboZYSuQMT8SVKNIsSAHS/+0ftckU2RwMGHrzk+Vdc
cdKB8n1Rpcotreh4jJjdcRjVGFwv1/QytAfPROUUHfmUYnJODMMBgH6lyNkPGtYU
vIfsTzJmw5nMnWk+GyIQXL08Hdz0IbTO16A2cGBxvEDyTlygPE68mIeXssDjgJiR
sXlBdbcy8pK+Fu7ziePh/31wiql2RWrlAGHXfE96JsjLT4GyPb8V2oRu4fH51TNM
sNP+lJ62KehYdFR9rfo7jN/hu/oVaZj1U+HqpGOoXolBKO123jlUUkvxBjTXwCNe
zU0pyd2ZD6MqL5eZFJY68HecpQDDGBV23o+Z7tUV2ZpxxKhw97E43V5Hf8S1gvxT
Sl6c2yo4xAwp/KSZsJi2rSkJS3emqPbWM0DsNr0dBRXLrhuNLkgn55xFEQQ1K1u9
Vk2wYRDOThep1sBdpTka7w==
`protect END_PROTECTED
