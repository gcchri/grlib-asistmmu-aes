`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iCS4fKGUbjoxlM9l2mut+GAge1l+TmVu/uLtMxi353ZsUGjxW8K13rUf3OU5XXGd
6BC/Zl/TFwBZAvmsawvmaB1dJ8APH4DZAwu6pAjnE15qYhcvYAfXI+AE+irUyB1N
mZLBBZIaAVD/0gGP3VQD4uv7SoYLZS9ZGq9uIoAafCr86l0zKkqh2EVWg52EWPcz
9hjauQ/1Nl5kUo72Jg0SyJCIynuexs4YoCyRI0vub8/rZnrJZtYGV+bTRLvN7NAP
WLXSHAMZ3J/vMmPssITyngaSaK7TXdk4VymWq+dcKqB+zBt/MwiN9xXBMIPAEUiu
udCS1C5VIZ7P3KS76QfBT6KYqf7wkw3ODEGUhY2KGe4oTvWRbag6STGuQhUBuMiX
/NvXcNaHQNS1vVj2KtxoJxcMY0Jd26uvOlYATTSXWETizI/C46CKM814c4kmQHkk
1/BLbf+tAaklxS6/sl2stF2b5O68vkfFlSLoEdg2Qj3QXWXOhbWduFuTvf0GTFkp
2QV+t8NR3P16w+dRXIQ0BT/b2K1sxY1HKLC98X045XO2RcgX2nO/SI8NxL08ut07
B9jmDhvnxShk0QbNDCwhbZmMaXS7Z8L9Ud9QF2fHDnzTJj3IFGsFp8t4nuKMU/OA
WI0zbnjo4c9ZJ0SiITRqN9HVbsiNkRdb9i8GNLk8NtRVsSgeonFoCsOgnstmDZs/
cI8rHXKbwFgA2oumF/jS9J60bgCkeyrzPFrmpfVS7+abaH47vN9KKSawtoat54DP
JCr23thTISfexe/SrU9PJaZfb5hTACrC9LDj2m1aNSwvlNkpHVMG1bK/b75ydNY2
aUqGsqbSlLbA2ZJCkdDqxMwe0QIHmcpwSaBkbD7u5FetD6Zp8R9m7gi69qHEM2MR
RpnjEyZAu4Pc+3PrGQtsrI2z+yyQU4rQxcCJlwL9A3A5VD44Wht/Rr8Mkw3XcftI
HsZbik+kH7ti5uYidCqVTvk+IjDlhL2F2EC7XsaHR5vnDLuqElMw0OAc4Mi9ncnH
HVGJvzclz88JrUxQwyvxz2SOagXPfWpNcLJTnHz+vAnSmryHlKzs8TXwYh/sO6ea
+CXnmyWKupIbNxjgerx7MsjWUt6vMQdDYiN/nycHXYv+RAmwgK60MIQluOKOWEHA
fMTckmGaKyzo4WEt6vBx2rG6oxyam40lIefC0XMe0OCL8NR4xHnSY3a2dR7Baqqw
FYQYtFHjGAwHsNiM9o9IYia1bqwem2rK1GBMovXujD3gWMeGHUttpvWdqub1jShk
r3EXZeZQ1sipzDX1Ojm7qw==
`protect END_PROTECTED
