`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZ0ceSwtBzzammnKM9xNHUUyNqGiGk5RmvJyKbjuQeC+p3V0qH0f3bRKhof2t/xv
IlX3CD+LmmIKe/2ZeQMYO2FzN+Sy9OlYKU10H8evVJ+bnp1IJtI/ec5A4CK1ojYl
Mjj0KkUor6foT6smM4jvQSQUclPW44WodkvhbVfZxlZ9+Gh1L/O+LMvLpNyZu/tS
8CoucjdfRFbZ6tfdU9GtE34UbytJrd1VI9NdHvn2xxeA2Y3HbP4NbADBtq2YcOjz
/K9fkvbxNsOfNt0SN8XbDVS+pDmJsQvcdCCnicWR/lC7EPtExHVPpOtZZ05o6T8s
On43WILwa/h3Z5pWntivJPfNh5bZskg5R2l2gkvqnG7cPiMSkYaTB52J9WA4wzoR
KMvqfX7HMw0UERWHfjwX/cxHvjJq+wa/sAVYZM8WHaiC5VWHJIdvoyq41Fcxym2V
xBft5vPvYMOvJCdqFOxpqA==
`protect END_PROTECTED
