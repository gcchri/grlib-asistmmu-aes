`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIlQNm++6/eW0eGlPie4t+Hdq3nt0bZ6D6hPq8tOINEMlIs2FxKJhdkSuFvm1Nc4
WYT7raQR8r+qANE5mNzAzGnRDez1TqjeP1IvnnEpK7rWsOwKeD4+mvmq5+cR7VjU
fsmowR+fQg7tu/inB3IGAyY+O1DoIFOdrxspA2GvvLf93O4YYR3wb2lfhEQCcGq+
8J47cG73YMBg7UcCmiQlyAFDJ5xya2zDjL04vkEBzVL+Ixd+JavVWeUsf5sKHSDb
`protect END_PROTECTED
