`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4HLXH/E9fL4NGPHKv/SSyasR+PuqlEh6hA0Djw/W8iK8IoiE001pq6De37SIXper
/8pJsnDY8douoR+xnwpNcaQGhOEDxrJIM9cwlDgKgpLeeMc66H8iOBG1K4kItnnN
CUPHb7M8az9s5j+UlM6LEgAdZ7qZ/vFwmf0dKfY9q3piRh2orTukuZHgKQJKe5sv
mtKiMhjqF2pBH0829E8UxemqstbDMNB+f3oeGE4AQEDSggGIkLXeLlor+ulsuh2I
y4yfMLM2aGSVkpLjBkhUU3ziPGGonrrL+C8Boy5NjcQvRLaTyaDWyhzz7vIyHPjN
klmtoKDlzdgah3pagEzkRQHArFX6QGlhV0kKItHv75JvWh7QMRSta+GOgF6BGEp8
c493u9STPH6vwRjUzYXQLfkLsd+azPU1Os3yBMVBehNrnswpciVMnf8tIC+sn3t/
FxeIZ4W5g6wnT7PJoKEih2zRTfZsD5V/50R+sTr9DWFoNHpppVSBjI1Wjq1sy+VC
TQD4tYCnm8c9z24XI431o2/2uqPwW8uwUUU1gmcPv/zY7F91oD8ZEW5NgZMWuGIt
OPb6RRofQpqGimN5yNiyLMmJW/WGIyjFI+gclo4dRDgYRLkWwWa3Z7Fji97tWSeH
+YJ7I/gir4CC4PaKXnfmntGt1yylNbH3SAqFqJssjdO8vSgY03RK3yP+41v1u4XY
mDaI3KChl2QFyVtJ1soGAkXVcf6uZc9VMcfX9h9w1HWpcvxN1MpFww2E7dOCDy4I
BhBeVTJuYru12lh7UnFFgaQFmcbEolGMTPW/TE4eXa7QLeGHstNrWU5s4vlPNWXP
gb3MfPtW36aCAO7j4Hyf3UNOISjSzprGCl3oYjQLxxhcOqcsyHTFRlOwHPgSBV+A
0r6q4ZqO/eCxIPYvSUzFGJ0Dz0gqHEYBzUpMAopion9PZWcJb449o6RRVxxVzdaj
A5vC11s/wCHnkuSYOmxaFnR2gGKivDB22/3ZJSEB8oKQZbq9yQ7LUZiLuMxrZk2P
wCpsEkgG6QZRk6/1WMRBXmW8yezajG9QOdeaECoFMsk/7iVqh9BlhRT8MOQExknz
PgQCzXsVTE51q4FF8e7K9vLHVh/DvIjwJWrpkBsHDcSrhu/C1+BQvfJxOthonNJm
8qptfswwWb52VeBdnvvYoG8xjz4oMNTs8knhIoKAIXBTUmQ3mTufm6A8kaeOfP+J
btUNtTzukEjFsGufyWd4G86Yz6ngbQKVqvt33sjcahdxqnJW63UVa5koE9pL1GBy
7rLPRkPa/o/0cMWtFYdwpr4V0Al++Pt/VoNoS/zg/e58YsAy48kCdPJjnsfKH8Sb
13WDHWsqfR0svzqKs1LPmjtPOyg30VruzRTFh9JuMGrIgySsSSpa+RDnwv1AXAju
XXmOcL2+x4QwXXJig/lv6iJm0TwaJTP9Z14XyJxj4TrVNC+vtS3qBSMW7cwyGWL5
Y9oJraaPejYRXMTutsoIovF7rV11u4uQgQNUMTbkcXd5ju+tmV+EYwCiDCxfgTxC
BVa9jw1Djlolz5G5z7GH0b4gypD14N5mqtYe/v/q3P7DC+fHVE8va8Uv0hrTAMTu
1RbNfvRJlYlzQ9IWXQPoIycTremHO8BqtiztCjAMv7vfohNBw5sQXeBu9F3cpTOa
yYx+6quKSlk87t9HJNdg01HQLJznbG0PBowl1CTarZ91q8Pva6rKJev0cXS+Ux+w
ofhGryoz3hUuQRhg9rNOUA==
`protect END_PROTECTED
