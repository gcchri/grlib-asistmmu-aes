`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FLrxqTvLX8wIzJ2ijICWgi1koHr/nOKlZaHB8Z8VBqRXlhvnGrPJxcPhQKb1H5+6
NucvbG9h5aNooZXk+EZhbLHfcz0WPfuzMtWj8zyDKi0fM8ZdocPkq6hOaQbhKuLn
L8Yd0gOL+RV30V9fL48q3HlZ8RmkC5Xrc4Lw87yR3ZgAAsKzq+Bm/Kxk4FJuFNLq
QZKMkVZaEUqyeZQcfMlLvpOgUW4HHlDLaNbYDy2POw5vB3+EB8QEH8eSEOqQHSsY
WD/PHz6fMD7otTuMjUrO/f22XkCQHdraerT/68fjVyKghRZ/dOfEgvfvGL/tWLPk
zTQFis6Wq4SaJ83+Iiy3F5IQxDAD4d0j1u+WX5zQLdA0Ed4283TV4tN3F1xb4fGO
YPAlZEY5OlDcm4VCQhWgsSwS0R3iOkjG49CTxG0pc0lmDl3rRn+xOoxNmG49jyo1
dcuwUwqW6QrrL6qj86024mzrNV894ekJKaY8OUP79j8AS4rLMxkBr6Cc4Jjmbqpx
`protect END_PROTECTED
