`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8m6518DtOClW97cP7m7ISWGW8cerzx9YIhMzBO32Q5rfX8yiIKYdJ+UBRZuPOTSF
5lQ9UA9cvSDb7KUBbr9iy07WGO5rY+ZrDEnFLNlpcNHKqbNTZSgugVvoewwYiXs9
aM1IGPU2w+y80ValdT39lanIyMJ9tBUVnc1aMZPQLoTGxloBwnXk5yiMBBpSuMd1
mE8Dh00aPOcps+T39w4dfXwyyVLn56CeJhnIS/rF6qIKL+yFhGxWKjR2arOWPql7
7z1/GJx6dDq0y9k2ZqUV/PcYigTDS6dathxxJkr7CjO9WLfVFd8oJ2G+aOygqMdf
EMWUt7WiQQ1v9DTGZvDmet/ouBTIhIuu9m5sE4OT0XbPC1pO+2uVZFapOYrVlMlI
e46RpCWfapHBUb5dPJCF7D8D+kPpx/WAsRzx5TRbZ+WAay20HWQaNVwKYydnHSyu
qeaA5icIYcDAGO6cJNv2BheAIZmRLK8CsHut8VAIhO8AHH1PbdR3/5kQllb27oBc
ca2ti+JjDIVKP/bHh5HTijlQs/u9TvHF60TvKdnI+WS6YogZ/x2q56MyqFXmfjEm
eQhcNUA7SjRz9bdCqxcrV/1htr1RC/bbAH5RPoB5lYuWPv2AkqVSXooymaV9a1lf
fU6S6GENHgeCvWDoCL+CZY+FUi8zc7FHMx59aNo+hIcuaIS+Hqa0yqQjMmrtPiIt
jVmnakwcpJKui4IPSnIRtamPAg5bXEPIF/I65pywGXTdiWPJOBc8l50QbQV68bol
p/Hq9XER+o2JktmRLqx1een0xEFv7uXNRWCGPMBTuQPLYk4l4mk/VwPagnsXDK1P
/DbKuSyie4gpz2IFd+QFtr6ZtyP4wpI6PmPUkS0kXE3F5Vd+rqvIHReRxRpzvUzl
eU7HQ/4dksiRTRXaDBwSDcA9Np7AOmtBCXKZ9bKMfFst11cmXLCUUKYFn5MkXKcQ
6Gllcy4tk1YpNMTdSzv+2i70pc2AcrLnNq64/W6g7J5xQHGegjBJIUdCMus9FY2L
6w0O85Kv3JEZD54V0ouM8pjo3SROY0ueJOedp7k0DAhB5ql4Yzk/pjw355FNOfoS
19spe0O8idTnKM0UB2gP/EFa4YTe6FH2A7esU8jAVtfd77VCN9Vb1sUO3hKHaufk
+jmFfhg2bs0WqmxJJ1VHoiHvkte+Jr7eoAgv3OyuqJg7QDQY4PNUVIOtsi5njA00
W4oPE4UifaN+RkL4LPu41dswHe9whE+RhjdXfnmldwyT2k7S+xXZd16dj1n8zZpS
QKpUljWpgN1IYkrz2BA1ySJJpXWBvJgJAFXplsL58wEfrh9EmbNvcaAuN3ipKqrf
QFBgYVbDwNy7nOIpYOJhghu+JC+sDGh1UjQMcSxsF9G6irVvLRBWmGxwV7zD3DxI
rJ1Uwga3cG9yj2oN12QpP1A0QIKGACQnWUObljQyMahun2EP5K8revslvI6h8NMS
WleJFRQ+f56Fvu5kGY7e2nPIqpRJXRIZWL+yTonKAhIxvjVNqyRDKxlDYWRRlcgT
L0gIoyOulFLT+rGdpXwxAl21QSJJYgLa9kK407kFRiDiDcE8h6A0bVtsnLO0ZF4C
0+TZtEt65bjcSLfYL9AbSNSfWOXPhhYM4e1lUtKmbcTm/VcljX0eShI36oLyVrBr
y41REX4S5j6ZDo8ANWjyVHoUtK/+LJ625ujw8xpVeHjFjRBDL9PeFQkOeti00DJh
HyJUDungGTKSu7RqOu3QBldpulfKGrDqgtv80GDl2nYavMoeFbi9GWoaFdfN2hA1
LrKm65ueDh9zPNp3DKT0kvaGh+2KUVp4Jy6iB5qpukX2yD3TQqrulGoeDSHjLfM8
cjZkeUk1Eiir0SZrdlPzagoucZ3tfW5K6Q/6Gv2ln1A+FFU+Y4+pxfDU8q6cIUyB
yCKjjlu7c1WyljNAOcMXpTbdyJu1SxTO9EkSdVWmnN38PCfDtTFvfQBgaudSnr2i
kasqVGIax1sbwmtDBLpIwRTNj4mH9o+aX8Y7mtuDOnv9O3K0yTxEIOYdFKgdDOHQ
dro2WbOLGa0TJF7zHa6z4AYygV3iZhp1yjJASaldB+41lI8Y1l+S7hmwsBtebVAe
1+z52p/HEgJxE67xpvTjM6zgUgc6twuzGlVBVXUQHz/EHkgnY/7Aw1SU5nK2ALhL
AfOdpjKCTev9lT/KxUVYPoUz65D2AVrOucB0neLIDS1y0cDWC4dH2QD7j/ne7Kms
NoGQ8BR0R+aoRIMpmoeYhidLvnHJktm7W9yxPVJmfTiOqwg3j/u+mmkUYF0du6Fc
18P0Ic9328HWpYHb+YdVeNV8xTy8kx0eYon52ouv84Y5CpL7EHggChR6xMlbK/bw
bKbodlwirnWbjEHAwY7EQzzCdFNeo0xvOuMrY5QxRhdFop4uF2wHE4QTF32hIz5P
HYFGGcdh1Q4lePs3SRG8aGtn3YAjZtU7kbxSWppLRRxy96ITwf9+RFVNNUHo/zks
Kifp3vbKS6xcWIg6trPHaLS2zfEQf4sB5W/dYmKvswtxPPS41+yFkL3m3XquzcLB
BE+YnO2R1tg1yxhMzPgY4T7A0PFdCEYQ9FM262Jc7l8eTaTPrt0I1n85B7mCsXDf
H+ML57rNtPOtxNoEvgNNq8UmpKY9iQAnnivlZ+Hl2iNsbivF/q6cLXxo6ZBP0MEp
qyQmKonxdOjVKmmYUkYBHR/p8K8vuaiVEBQ6ZWlLE/vk2XH8iarlnhHZ3rLif+L7
Zniwz7izqEi+CI2pN1x5U29FZrq6NnP6cI+4mr1uccxYWGs8puXRi5obo5/pYVt7
wU++u4xk7I40ob8LGTroP3KYe7fAb7CYNJcNOKdMnuN5vpoFAU2e4FuHFaSkbEQC
fFh83iy7GZdGs/IZdp4307x5A/tyjLSYdCNyFUv04e3yuAkgL3VJVJsftVimvu20
O8wBNS6qZ2YbkbeTkIZfJKbUvwYX/C8IlvaC6iORIHM2nCOXbvEe2xLzTI10pqNi
HLJSrB/1m+HfwErtf7Bctg6vJULsb59koBxANJwTputqigzv/qETUSzql3Ejync+
qSHRs2nXwqASFIX2kFr8cf1ElbBuBlnNZRAQWLrRFr5YeOIAVe6liENHBiS69Ulm
4CLcsyE3Bo3/v7VmVYzOGbJWNYPsK9bg6xwKb/fCuhCBLP6Ri3ic5PMPJ3bqZbYL
s4GOgg1jEDMnJuc0WSgUC0LPsKLlfkzTcdApejodAAxmJT+SxMWJB4s4OoW70kYE
3GoQFJhPUUkE+9YOie2tIDKpVJsFS/t3Bg7knxtvWv9rzdHPsgrli5HNmPaNmL8C
86HcuxN+/f/89lyWR2NoHsjop4VeVXUEpUj7/hSDXwpM3YFFE33c104r8MKlZf4T
XGQXaWxLTbS/srnycPG+QLOQve1Z/UJ2WSD9dH67p7ADFnvBTGPh4NtPCGmgdqT6
W74vwH0fRpRfEBqe99vYxkgZCXQPJJDaiuDbPGOjpOllFCHvbznhxeh4XEMD/1lo
PNB/ZnPvkxshfAf7QZ5Cy5LdKKFV804bYDEtTQSNzv5FRfzyLUy3fjooRAABVuV+
Xn4kWJr6054Tg2rA9dvUraZYvLvfiVBaRlnFo6J81dxBMNg4PjLGKOv11iQOOzNL
Mah/nc73wxedrkZifLlkykYwRLs8iAZlOIS5PsfcS13VFc/9VkB71cHp1+yv7GUj
+h6fxhY87ezHbqn/+pMV7ll7rkTDN6vhRpn8RZ4O57QQvGuqmKOxQREg7CoNKB5p
D2YL6Mase0TpfO8i6QTj8H0pTAwrJpohsaqPp1CsfWkedcWc1asw6TnhJpymddOQ
rPxydcatdil7oUf690NMjxBZzTHZWJP9693sdpZ/z/9WhdMfge19ay5lHgXv6PgG
WhFQu4Y0eh3bSc/a/aX5aSROsdZRcFLuRZ8oJPabbFOd5mgtfMKLSRzpznxDoNtA
TpAe+COiTDB1n6TP/NPRE2Xktnx6UONlgpgvOdCAew5EUWco/FmKaY3Fq0W/ZpdP
Xx332jMCKP6cJ3oVnhZLJ59lYS+hC16pmVFdrLIfs80KssEkSBn09omrcEfL6+N7
NjbtCbmyiMamUWBp7TAbr5N/8OH/Gkc00++qTdb7ht78d2ATXGS+I1bfwUlbggCl
GFj2+O1tMItPMl1S831j2tt/yLhecI9Gc3Mti7alllsZuzb3HrZP6DnJtz7DH2dm
OYi021koRUhTtzM2qxeNBOxs/UeOp9lJzptK3UQxHjsj68EfNCYxdrDclcIjXW8q
xToIJ2SEu8S1wMfYPdIzlXUYBdPqAEBIWqdmqpCqZ+P8e9LqdIt67xeNn+oRU+N6
YwZyXvysu48iIwEOQWsGROnEEdqsUDFzjk+/6DZQMR6mFq0zFLpjrrt2bL0IQqqB
qxsEI98tS8xY1OhGobpuJcffHzaWaR5PyH2FmjGu5O/tne2jUcnZOjCOZic+Ceve
1bCNdIL7weF7lmje1O0+6Yp98kRJyL6BllIYvYIqQFvsJb5ZepGOF3zo7vEDZvGM
ooJXZDq2PlFnyCub5Me3NEiMXLSwBRS1udmZGOdS/yK7OCEP+MnGN6s82XKVmmm0
DVPvmnaFoWas8QvdBy+REouQs+QFxghbVdw2P8ketE7WFj9vT04hQDsZpKdReiT0
TH4GkP0Fy0fsBh81e+pLe8EyDCUSBs3i3VrBmdaRfQYXA5IEsq2Vw7t6T2szalzP
M9Q3YlyhP0Jb03G7fa9P+g3+vsAnqcCM3CFEt9ALLxriaCoKgilbLM2iA0YXpqZY
+knQr+RO6nsoFOkH81B8zC0EwgJnXvvYR9axrky5rKvGp+D+vOeZw3fpJF70IRHZ
y6xxfeGadar5nkGtuqW6o0T3/+AcvcSkpDza1HwTihxTdl/EXIu/FfvsJ/twdu77
fuQk+duZ51kcyuDCt56TyPzHLXmFZM5TEHzrm8LFE+VVoe7RqCGR88p5euSKDj52
T0gDSYLPwRsixDcUk9BoC+SGrznDpOmlQqIXa6RLSTKdzGsbr7cTa2FymoaAPh+y
9IBkdbpxes3XGNFY8JMBerPVZcaU5WAESIFNJni8fNs=
`protect END_PROTECTED
