`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nhs4Y+agCX8su47lwpRtQPAvA1Ib/V+8UECdmxu2iAF9KnBBT1a2ylZbK7V1HSD/
T4Cmm1Z+3aA9aS3pPauEsDeC4qiBOc4Fs18BBc6VUpmMlkC1RnRMQLQJPuKJNyY8
Lfx5G1iH/h75+VsfhHTRTFleRO/jid+GjmAfwfcRib6iXE3HP5JEg5ZN70TluUiD
46r1iNKQd0v7iiSlndVprDoGUScRDGTC1YcGNWEqBTPwHIO8no/qKIyVrMWY8NAu
`protect END_PROTECTED
