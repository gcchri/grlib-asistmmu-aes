`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vi7Me27MZqkvIaD9MB39p9Di+zbC3LzGtFqthH5/5RkolC2nTxAUvSX8F6xgt4b
CYk7itDl+R2CWixqwNmmoSHXz8yAX1vZ1cgKFYkCvKBhia7vBYk2Hdy7PRX2Uf54
EZVAJg2uYBgfc5SOQsK5vqWKlDZ304kO64QPxPMIXHjROC5T0VjnY4q517CbBulP
D1oK/Vr2n13+UE2GqZ5y5+ts5gCKwzexPj2S3dR9wjd7zwHXVudih7Ug/jCqtApD
eScqjcFAiWtmd/t/yt2uNq7SjgRtDsFLfv2FKX3Pm/x6t5WyMS5NhVjz0ORT6Ndo
fs5teo8tNqB2B9LseRKr7I0e/uuMRMCoWh1xvuP5fiQcsmZF/H88PIu8LUs/2Gf+
fof/2O/hFAu+zrXKBPjBzoNQoZwuNgbfmm2zWKqw8TIuT+quzgkbuzvFGt+lPg9j
4thbUwc4zTSzefxwMzxIra3nCBugEizRdyBUCXD4wJgUnKqnnse4BWsjsS6Yhxk1
zFhQF3CCErdm5jdA5exNUq9fmTLAgrBk/k8qIQ7WlTuVudMNzVtKHGisnNV01jFg
9htNuCFg1Jb64PcG0qjdb58TAgObDkXqhzVnd1J5z880eZ9JUNoS7sIalFTMWrG8
h6KUXzc0oc6mmaY5mRQyHqkIm4rq8bYuQAMoJDst+maYvvVLfA3K99VxPEyA43mB
vY+1WJtZJBnp2jAanV+q4+FTRp2aoaY/XsAhvLHQ96ILQb36VYJLApn/rIv5Xm+D
7tdUNyB7dsy366VVzkmfaGMf4C6Bl1Wlem4ROK8rntc+fjO1vbVRTBCXGzAP4Ahq
GiWoGOPvr/X5ukYVuk1whA==
`protect END_PROTECTED
