`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jdhHuc1xxwpTQLiTSE3f9e0ixcIQDugno6yX35ZS3/SKQ60Q41dPDXJcVU0X3Org
0jWpOxDHBzUpXnhOVHLM2ncdsz0mrsoi//NQaElpJm/SEEULiywsYUJME98F8zBB
shvjTXDKbd7zVVxYCOTb3esa6+lk3ZYWEt7mQ899goU2R/aZ7+Cex25BARB9rq0U
pzz6cTi6onbLkQrOgE8G+vhWLlecpPJI2RyVypePHZ158a1zZObpnl+jn4JYtHIY
Us1bVKAh0FialSzofKhBKxBlwYVyNMvJvRW5AgjJYhSoizsNsB3NSpJNNSvyeQl+
LThrve1SF/1uYslLB+BlG1/RqSk5EZwWivbm1Fx3J3ba9vvN9EHyWLhn597FsAd7
CoMZasN+Yeafn+YfZcm4ju3xl0+A7crY+CkavxMrxm2i53h4JKAtZQQAgWfKZD4a
TBuoZEUiqAIoCJweCxR47dz2ZBjXzeFL/bXIf44O1ZjwUrNvePZxaEQ+/Int6VRg
aelUsejdIYxxe3xymdifZGXVtijrZw0zllz8+2jsTtzY4goZ3qs4Qy+r5vEo7FUM
JNEwKdZkRE2GIOXBf71eoyDtWXI1mUzA9m6oYL+SYYhvsYl3ftBM45qwWPYWOOtp
o60vYcz2SXboJtGUzu7T+HLcDwub2fGlCh6gVmPkYGrOxuLyHp8h2rBtqup3MWQW
LaHUw0v7zPUUGaXNyLZpwZZogxSm4hx2Broxr0VsOjsyeiQlY4VNJ0GSTxGu1wF4
n/apkG8DGU7WVwxJSol64wvIacZCN2xzgQRz+6mQvcodPsqmotcjuhNej06lI2eC
tygAyz7Ft5u3fCS3CgcbaRP+OjcciUC4b7Xa4ulK0IGxeg8fJLWNWpRZYSBzpmFz
AWs5Y4WeZotNQHrNIBU47BQozDnXcbyYQr+O3+EizraDErErxDekzC6BKBBmu0nh
t/EvDwXILdIHyVbWvgThAJ5n1jZWKk5ymGeMqcH0QmCMRAVzOPD8e0shoCxD6kt0
FOZf1VXJdgNbe83225Gnx5eU4u1R8xwmGr+cixHhtyFLSPXJli2y8oXKjP21T3zj
09826tnRsm7oCHHxSWJdjIzgb/g0hqQjKmybXQplKTcLH4xGr87fpd5c1ES1Gsf3
6AnzUzcs9aZqzb7CfofpH3W4HN3arLQwX6iYWIPDBkHBQkok3LRo/sNi9TsMWDoV
4TzJTQKbp9c8LfS1WaSUF5uR3VhgZkRwT0rDnehSU/9D5gfoMf3vL0Uqzgwj6P35
i88NvxbPIQK82KVIdtsuy3LQJQ2V+yKnmEYk9bid9GQ1excGSCtlsUEPCVGmj8rg
+tT0VeF1NVF4MApMhK8074lIOquKRFOthH4H00BglpyxT/pF4enKOQ+EkWg5pWKW
C9vyEFzhwpUHO02TkeWZyK3j/05dXIJgXaYUSZ7B4rWWCAA1LZAA3EsBCA+SOtJG
`protect END_PROTECTED
