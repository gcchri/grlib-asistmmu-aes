`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V0fQZQCt3RE6RNER16eUtTUSjxgVn/JYJ2XbsXeOnbUi9UmxieUAwtbeDXqRITcv
mSI0P+pf9eIkQ4J72utvCJc0f3v7VED6b9XoWA5TDFxvFbLj9r5yA1lsPmMwEoIQ
y538uYotfsGYAQsIjaizBGgsHtTPdfdoLgSPH3R/0q/DEAxuQqCkZENe2P6kCblR
+z0W/zr/RFvsBX4Vggl0PaHMtGzhqy1fqh+t0FMH0NJLfL0gbcPvOFiEVABVKd60
LTF7GSU8rCgRAlRDNPh+/AXIVqoKJNM1hvBRzKlz/kwQiY5s39LU5ncWqVSxqM3K
`protect END_PROTECTED
