`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1q7st03xfzk0rJAPyLUEFJ7Cy2LZPJMJb95g7j8vLATRjjRKtPOTU38tyGxp2Kiy
Hxd1T04d2oq3pQ0HrhK7vwz2VYLmib1kGSFEAsuM6Lz34mL/Yflo9E6K3ZDu6qMT
gj0r0cxN1IU2Qw0buaU3pSh3AEzDklKnUMuOI3aEsYSQiSbCW9VDDURoF2vaXsvB
fiWJ0Vs2mx3C3gif3rpz0nXE4xZmP/t/Ebf/gty/PnMX9S4yAlbA96MCS2sqI23T
xHLjFyyluJk0kuO5gkXFWSx6gXsBORQHhXX9bQnTikpHygFkSlKc4+wAfD2uwFKr
JxEzDMD3J47KzHUnHkgqhXe2lJgI3qaMFJPE8Cl6AbNUSNmSo5zOBmUAje+HOXqG
7mJe5szW3BgvH183ZGcXAuNU88aZmJS0FyeyB/QtpOF1CyZvVDBBAUS0wueZAIZW
xUPtAffnoP7XQIkFG7PpuiajoPzbcTz6oMxQWajVTmpu81UW42PrBFJlX73521Fs
Tzaa5u7XbIIlqJgMNjzl0sFwT+thBFbvVYo+3ssC8wXfjPbmdLYfqvSJyRHq/Inj
qw2+mC2OkE4SEhKcYHgw6XjTqnvZU3xDvHy0fiGtIadX2rDUwlWly91d8R0jBZ2j
Lb20l64PeX9ow1Hd/rg+lfpnnPnqKzxwGUFVN0oovoBFw2HTcWksEM4/2dtnz1QE
uM3Eu3sFZEVkfE63vL8YWq8Q4UMdMPe6A+2oZvmKrN9zcwK3xXdFxJLuIo0hyl4c
+o39yoYYynhfOWDD/saklDs5uHXxWAlV3fcU6EXiXqFBlvZ86sJ3VQ4lszCyPKLC
dtcuLJjH1Mu2JjGTqhAfvjhC9Dxo4/pamNaA1UfEVfwEf8ag0WRjTEkiykR1Dk0o
9ZxNFWf+ILJeayGD/AQ8npz4ZA6OYHfDVUjibtT5PuGicKdsjDz0rtpDccr+FQOc
kB2PTXXUXMZKqBXJbhiWfLqy92OQzpOJxrZbo/DS7RfvxwwKanGshIj/Ab0T3faP
yFTKxBpL5yLspk6KnNuNoBXQdoaDtWnzjpyHEM81pp7/jVzUM3iQL6k7eZpeHyFX
02302l9pykcK0jPYDbo4j8qWAHf4rf0/fs/Z22omFoaP58iTNSpt5NnigM/6hW+c
Oc7d5nJs4NdJymspD2Bkfrp+UWBukLTAwZpWlTl14wlJRG5q57o5q/LFSfXG80uo
c1NBb80+/pavamtNukgJKd9SNO8YuFh42QKQ2I7ZFA4QdzvojEqCPmk0KFca2Mby
5zYJKLWv0/d5Nz9K5CUD/JlWMZCrEJZKsy1gdx0NVUXsvkIoN0GDz0NwEh5SNSIW
POSjVyGxpLEZaQ3pa+xgWw54hNDHO0GElE5mi1cqoz1qGynZDHt3X+ZtZn7nIfYV
ETZb8v1CORW19EupYsOeKdTI56TdiQ9zLWnHBB/PTED3GUwp6N94Iw/KHWjQwP0P
q66D79q6/dBEvoajt+e8T1VbM0IbAUG0XCpunP3NPecctn2x3DhCaGQzvenjslnF
ls6aUb2TQ3U1ObyZDlmXwiv43YrX0n0obmL4C1oakMtIjPMsBC7DHVG0JMmIt9nW
V/88en+2usC4KBBYPnsq6dkElXGZEFPHWnoJrwQdp59JpONbDPYLKeHt6VGUvREh
fAgesEz5hXvLOP+AOzAwT1jWDiTa/5xLnPs76G8UBWYKVNYC3BVBIHAPhI39APJs
2gusPSSdn6PsyBezP78Vpa2ZIUkAWU2R50+w0fa2Q/DSjODX0LdQ5Q3gfzX4AbUu
0+rFcA+8h187Dwubc9Jnlcq7xtSYGm4icgTJPcnZTHZgSNiSVhEUmnL+BzPAtT5V
P2u2xToXW86HwZkt1GuOEXf9vfLI48VepAJAmSuCUmus84V4EQvPsyZDtHKco29K
Ixf8R/1bcp1yOB5p+HlImDP/o/Pxa3dnxNn3HHM9MOtqjofQtZq11teHEj5Iyk3o
/8cM3TcpyLlZ1YLEDFDfcVgeOk3e/f3PsKYNApGRa+U6Juihc/L9xIelL4gwkAQ/
eX343YKp82Z1+BSCot9t5X8ta2nmBLtRwBop+tbzAQQ366HyK0S6B86VDCNlw6E9
XtLIRbcb6he8zqcEkp/PKHl8RCZgyOpXplpbBSycxkam/sUUXpb5MCzcSXEgxHd2
09qcUplxKRBkWPHurYteRjIp3f0yDgMA4qp1MPBNGMRnvWnH5HnVkRknGMPExY+6
oLt8UWs14wbscRNt299SDY5TA7SUxvPkFWCmshFvxdOBloB8BCHi39f2wSfeBRt2
Q+OjcZ2lnQVLnn3dSTIGgD3p3/tBwG6zam3gACnru4F76hD+MQrbEHjNk1Emt86h
rLsuxBGjZXbo6niEG1lWc5byUGc+EN1NEcP7eu92mKg=
`protect END_PROTECTED
