`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iO7ezwOA0Vpb/JLkEQYq6DzoroGWGbIxoeR6ZL4iDSvj5UlAMKbjIbSTI21ZaY7r
CYn3IIV6jQgj6mRdhFVdMSYMkzK5DIV0zXTR6bFhixXtZDMbxZSvE8A3opmU7iQU
R0nX5+1kyrrywb+a4+oMHK8nYP3R9s/m4R3zcwud6/+Mgfa0Gsnak+BC4Dw/sz92
7pvDuQ5of0+1lYJdOidO7isEsD1zvsTweuPs2638axyIw74R+RrXX3lQLMzPIji+
qgsPa3ZXdmnDBvVoEZH+LA6wbpF1mPbMmpNtLUNQ7AR3dE6U7WIS9FgdvsxgkZPS
zK8e6WQd+Ezoqcub1kHPAJxvrVTBPBHrPRjOMaoA5Slsx043nOaWkckVZlU5gmN4
h/S0XGoVbBGofDu7LincNzeleF/8ox4+Rpe6KvSilQE=
`protect END_PROTECTED
