`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iE03rd3lfxCPgqWdKjdug2x9rTLyqoSg68XvSZnoI86MoFioieaMrICwO8eleigF
x8BiqVZD7WkTsg9p5DEJckSos/xM9aSgP2oOLaXrHm9+cVIydIjky4RS91WJ5D4i
aG1DLjsrWL8+E4Cq+jGSTdM+570sJypFv8/mqgqG/RCDO1bE7VbnxXstcwHRuNkQ
2DDUaGu4Vq+LScvYvpzZEm9CVeMEm0F7LQUskUSr+h37pCqCwiYewe8JocnsfFzZ
kLIcND2wetOAtay/Kut9De43yXBnym4XbA7N7AjCq1x+v4QxC/WueKSiPW5g96V9
CBeevU1n4QD+sWPz6Lf7FWJqNMWJJmQd6sksf2PPhyJsviIOY0iAMZivguN3Z6Ox
CLT5Y72wvMAzo3OrkeBar+IJkXxhi6ZSySSwR8dTpPgaigg9zRS/Et0ng5GPTCSe
URYdqjlqBgWfl6S0SSI2WObM/RGXDpJQjy62R74Jnq+awfCQ4X8+lJyPY8kEsWe9
AAZkP9f3D76oslQPrNxjRZLtOjYufdMcFDLsdJlD1BfF7/zjM3F49vWocjdry1uZ
7Saah1r08b6rgccnF0b/BAgH6ojZ/JVcZyaM+eM3cX5Q1I5HSynPeawmtACHFwaP
KzAXHQeEEAReo+NjxklYb+lpy2wNv8c2Jq5/Z7PtXrXQsND7gS8M1KtYgBCA7sA5
R/IZDoFxeuhModzf5OyuINPYbcbFft4feQJQOXCR8vsSuEOMIFSAsHarZH10fv6s
hAmEYD/IGkd5JZDz12aGJalnQU2xLLJNbAKGa2j+SsVtvHNo2lI1CKXRcrAXDQuO
ytB/qrC7JuEgIlXNkFU49xqdORxGLya8jfcGnr/eJ7xARmyLUaJi2PadAlVYVssC
Uc5m4Ex/ZSuByYKOdHdM0xjr6Vb+QYYKdNb7RjXH6ZVZULn4QWUQ75WYIunltp0y
rTFlBK2+Z6FNkwyRpGy4TyFjxG1ZJ+kCVF5RQAW8jA0oDkJBi0Lw/nX3RsmDUGFy
`protect END_PROTECTED
