`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZeHNvnopBc29Mlz08OSoASMd3s6hHB2zUXhjziAMA6DjYre9Jh7rGgg+0BsgjnWV
643ZYOYWugMtA3gzhD9t2cCavj+5xbp17p0HYcSyXt/V/oJli7xZZnLtAbqsXecd
PAM73JAtnh3+bVBHlt/4RM/7Hv0GKzSIF5/Z+JFg/qNzN4SqmGh8BrRBc4IX0oT/
bPyCeinVBvLSuZZOgg6jCoQ691HqQCWg56GULG9I4RWhwOdASS6Iwb59fq5YwZ9i
aTHq3WreIvekYMowiRgJNlbdh2mXUL+20FD8PFaysswufZqYEZ+ISb604bJKwINs
IfSDyhkB6oGaCAlGbQ5KpuoqFnH8CBlTnNHiEFyrzv8PeVGD0QKFsABNPrtC1/x5
S6P+YwWhTQRQqXgwmxw6Rw5F1rOakmXJVVmjLbSEMcjkqD1OGhX/gmZ11TeEUZav
4Kx1rkXcO3yPqJ69obpIQ0CmID1aspdFE+9JIcWGgOMYNG9HDPL6UPM8IKeIep66
8sUAwGUcR/WRcSoa/Zu+W733KoS3ozI+jLMSbticsJ3rroVKpLe9Ncua0k+/ZtQx
cTTnYG2o84M/Om4LNaila5EF4Zq9pDQ8n/DM7Ta7GRVGH1NKGKMUjmVtnzQpHeR8
exiIKJOkRGgZLa0Er0F297A1Bi5gaTN0eci2I5h0OFsEzVNKA4PRftcR/xbz2o4E
rGRm6GQzaB9ep+oXhN/OYzU+xnQ711tV6IeuWbk8930qJDHunkSbCAha3G4ni+j0
wLl8Cx1VHdiDJcf/zS1aZnQmpJNPvRNdkjnykM2eYziA+EqGIol/gytPjjS2Z6G5
xLbSbc1e4DotweTqmgzh/QWl2ieoHaXtm9IRYnAKs/du6y8+HqW7qmkvVB2gZjUU
xTgAP/8Pa1MRUP75aDivhsqOiUFxLTcwl2wAtZACU/eN6rnQfL0UC/CI1t0f7k8u
`protect END_PROTECTED
