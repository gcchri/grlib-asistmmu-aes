`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucspFI6MS5kp2tHVxrlqLen5j2gFElJg0FSGKU0jONHSKMxENBrUj0H80H03OSOO
LiirgtIzEIJoM8/6fYHVqYCjx5RA0IiYjALILqlX4lGEJ4jF5+/Q4fI8mGbFftBy
0tM2HLkW8gZpwx8nXOqbwpq0QSA9NFR+7Oylu5ikCnHcghoscABbcJ/mb9lpNtJ7
T3RpkZKv9JR12fb36dnodGvtDYGejzsneIpT4sbxMDICLevmTzrjlkhOXLVhOGvY
2EEJdLxDWDy8QxZgrw+TsPlsnsP3GfzGEiVrUCYxw4kCtZ5sfYAfZfroxuCpsfgz
fOw3woCD4/RcI4dy3DsGvbeKjyVBEMkiXE7jrcKdpb1a3AfzYXKNl4Q83r9GiBMR
8iko8RholjjFq1DahJzV+xU4Yq7R32sbcRZvNDBNNc/GDtRxVGkFwG1uTbD2rQnn
w0/mIDShqo7F3yvjUlaRgDmy2voYLs2klHQ0kSDkUlJSck9YgBcoXVNZY2q98dIJ
OPOACMgTWjioL0RH4WVsaA390X0H6HEZZQyYEf+o3oKaqXtJslzdHKINTETdvxeI
gzlewBD/9u2ogXHMiBGqpmWqqtQPkK0Tno9h43Tpnw651FTIb2M+dWUjzmpF10q1
1YHLR5GgwKFqQqL8siJJXHCoGU3rrAblaAymGW+mxFOKPtJKfDyNn3ub87+wDG46
HabXrgSa9HviSfv7HKjRQcBV08WEfSos1d2M/kDBQCt5L4JKlew5LsXieIQNytu5
BGTnFy8noEWOvqktSI4cbIxz2owIE9LJwUF1IuGaDSU=
`protect END_PROTECTED
