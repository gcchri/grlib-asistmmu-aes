`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
paRpndO54r/874nnhGiMlv90PCop7/o3EcL1yfF2MZfswaeYQEjSpzYKE4IvZt9J
Fmo+tYt/WySkpDIrbihVbnOyHwAD5yWAFAku9+CNuEnQZi4Q1SJQebMiRznmm8W4
AWG6ERM04pg87AR5BafogeWl8jgLNeNb6t6wDltC3NC6YUpy5n+Q8HxJWbsEZAnO
u8W7rq2rq0D5t0LFXar2bkQmD3+QN1kvyCNP93252UNWH36OMoOGuoMjQACaeJDg
F9mIAzNveE8u/B8K6C1rWvW/ecV6orZgozek8iZ0+cYUlGLVqRZCRsjynezRknAu
+PgohceEZNRrLheWLyj867LreSZT7bVEbNcEfAy+SKy2s6Y4INH23fdMGqe7/ESe
s98XWZNpOrkCDdcQi9V0pFIQcWSC7lctJ3THZ2+yTqbC2PcDgkT0CoSj0mKEsP0r
Lphi2T+IRDyS9G8oEf89GUGCQAM+tL6WZXDL9ltez0ZqMyUu9LhOtFXxZlbm/U8w
dW8V+/0WJTghSVS9t8AezAZNavJRKuonQOXy4tXbvlD4UiU4ra4a/dp65QGAUjkr
HoWkcgbAQoEsZBtLBdZmxleYC59QDI8gXJQYQOilhdHXGwQtBfGNjrJgsbJK/esb
j/dyMawF0XUak5VSCKcbhsJWh0Bw2nn2vRjPK3XUpVc=
`protect END_PROTECTED
