`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+41Bl1FI/9ICYYctMsGn8Yjw6kO5ASxRrPvW8oFQ5Nm6H+CWOS+s7jrlCPQsMBD
meoXAfDklnQ/v2fL8hq0dBzqEFyKtA0IijMBG6HMtmP3/6hwAjXCFZqe/T9pRzv3
tabucDAGiAbgqelhsTkNP+56YiLEWx0MGrI62xnIfTVHdGNSLliWHg3HXNjC+bgG
Ndrz8FbyHOesMISyrhmw5ouvbDT6Dd1e3HAXvNjLQzxrvYWd5NielPm3z144856v
2hLqog72+6GG7a3WYXZ2CvC8XoKmHDq8BeWKtNF0UnICcRVU1kANb994+HAbAJW8
puQlll6EPLef1G5yX9fvSA==
`protect END_PROTECTED
