`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+6PTFOO6xbpl4Sn2TbAg7jtGUZV4GuNOkMtM0H0xRuDjjh9L0FAM1f3YLZASTFIZ
CEOlXrzMMg0vXcp7t3MBqjuVvEpjfr1o+j9DB6gRWf0vAL2PGtmasopZi5QRm1hf
EpQPSNj9UvTH4WuGuQEs+dQe9A4u9neJTaNeiOG9rrySIenIxqgpnnYqgqVhAB7x
xu14x9n3nzzH8r7wgxwqZnJhx/rBmPTD9Gcr/snNhyYtDZlwb61ng8PqI6ffUanU
w/vKafWDKqkHJusuUkEIwJiK2V33BFHzuYfFs5WPmCwl5DuFusZ/iz5Qo31iO0ig
XsJBJxSjmZ2HL9SOV+yKdH35sC9amy99FhHZqfEg/zVtF200K9trABpqRbWFc1q3
oaPCAmGQ0o58FEk0x/4zFg==
`protect END_PROTECTED
