`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VE8SenmjKUO9a1dq+UA23kGpFe2fvrgw+xxj1F8suC698OEKlXQq/3ktoTu5wlYx
8ncxQY1qP6pv7tT8d2BRyLH1+emAoq2YyeTG3MEXUOqffy5JLsNtcPtzscHueMkX
Nj3X9n3Kfl3WS0U/uWp1sCVKCXBQ3PI1slH+06+H+eVCBiJVA366LOoVFHsXPGKI
6zeOFzaFgc9pYq3NcZdoDTctVr+OoUN+c3P8K/rzFLtRMSwlzMt71sGX45Oomx95
0otOha3cfgrm2YUUrJfv1ab65bfSq6pVRMTPPj/4L5qfQFQY1JJ/kCKDrZM9/gTG
XvxFj2tlNXW8cWe0Wf49x8GnQC9eFKakHv0jnCrlF/Ernn5KcI3bzet+ZmOvjzBP
Vs+Zg25pV6fs6tExr8W7qHPLrKYdQlioczqaJK1nodwUwy0DS0sP089V3VbUhtXi
fgO6K8Gy0wcXT3gBYzliTOsiANV7AaAYTfIO/xhKS48Dlj01fld8BNOk2ykAUr/v
vftWeJa/vph1bUfSJ5rP/x7rtwkX0m7OaglbYn6OLgMEZarNBUfYhGpz0TXBY7jX
mFxgAMbx0+urfgjpZKj0k7wHMtYI2bg8S5xVjnAykPCk1k0jNJeGP8R+8RPoL5fp
+PcmYcQkEG85OBN111imJdjU232LhEPrvrZuhhr41yCEfXij2T3olJhDGKVxoVwn
mb9HCe/n9IhIi0z8CcwLPW98zDYme8kc/0m+Nm+WHlcEUGN9A9tXA+Yx/y3xnfsp
gEus039J/vlnzp2v2qAolwZhul4KnKuSGuldLySevi+qmk1ssTl1LmX2wAxMfryj
H0yNcwcjaDqrg1lRSRxpFpDOpK+CKdjruXLUDWRuiORb0Jqg7TYaSkN/1JZnJk96
nwo4XDCij25IeulB1LDWSSADr+Zrz8ruqnD9jSyR39WfxOY04Vesb0mKH42MmVOY
umjjUy5PPG79caJsUGzTOvTZVr37aTg/7xsOBbII53DFl0mXFpaoiGZhpIafPFzH
dB+xwSosWboN+edCsXMHaEcWIkiTam/3O4ZzOk92dPcyBVyuQqJJpqswUlEXaxuJ
2iQZyoBPBjm8juC/Ufvs52JdTGQHcFdkMXFJ/eutdWzz4+jNbUCAcnLW8Ah5ZZxL
tHy4H/Zo8SR9pem8074O6seyDSaxauw6M6GCU0zDf0OC6JINkkbdvcSW//S+J1T6
EO/LM9sORbMPyCx10kzCHHs+4wt/5gOfxMHtd1e468bPS/k6DjwQJ+DXfpdhUTbX
`protect END_PROTECTED
