`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0GT2INAh5lbPw8U24667hxC6GEQw4UdJ28pSjhYnXNAioQvxJQnsvMyes+1gD1n3
SQz0ed/uugepDkPomxW7UshWJb4m0MgsZVy0R4NELxP/850ra7arGX+A7znI4n+F
05S8CK8d0FR3zRSpow2WB1M7UHv4+xrqO0Cuycyyz675FuPxG9nbsSjzgU8yOdDJ
VA6MlC3lOsKilJq/VA1VdC9Qla5atod1zvoq1hbBfkDjc+9ebDkgIb9HdCB+YAUK
0HNv6123YIdUieX73YLK4Wo9Giy5lDzjDSu5p1g131u/u06SIl3Hvx9o5V5YiPKl
M6lxHynN2GlCXjK2mxCrcARNz6EseYYjd3uSGcKk3PgNWqw9g15KvBx4D9Nd/6hR
5hZCoo/8Lw3XECavd3KJ4+rRKuOuyQrYHNDOE4JTFPrXNP8UGv+RrnR3GIUFKCu2
YgDa9MW1ERBIAi8lSFgTlh1xh4eMx6sKUmAoTtNfSP3zAjNbqp7nUyw6PKAYPyJG
Bzscu5eA9UktEhgm1kR7hhWWiU12N7LGCdIk8EwZ1K9jJENBhSlXb3k41Af5wxH4
5bZaSQcQawygoAstm3eaDteE7wyf0f2zcfHENe6XO0YkU7tySe9JGv+0d1y3S+dH
fZBTY94kYVpF69AZr8FRNa9HwW5U4p+rZ8NuCEWGFxLDYf0n4FmT81U+mgHgwUpX
FgX92jAdZSYYR1G22KrMYP+c1nY+0hI6ivyHoM9v9QWy6nN8aX1z4rRrQDaodXdz
LPdom/1+k6c/GThFYljgOzkp3iJHlunqR9kIVEf1jNauH2BAkaFFYn3SrsnfPJCP
DWUd/NjoKPf57c9ITHCbExUk70hiletfHF+4rWQnxHDj8KeVSr7MOJcHLKcslLFH
Z6pNVaDcf21NsCfHWUvS9m7ygFrEIE5ch5WynZw1lMvBPwuXTyYvE/JHLGzp5h2n
`protect END_PROTECTED
