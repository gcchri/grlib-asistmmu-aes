`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpZFwQXA+WH3P79wabjs9U5VGmjZ5sW3F+u8flhWWVAZxyxHFOjfP1wHofwncyzo
AXRz2U+EiJXQJ315dQ8Apcn3IDS/MWOES/NOuF4ZiIgGwCzQUDpZ6JukTF5tmxVN
Fzlg6iNE2VpygP240qNSwo9KyOlpupkC2D29qzrk/j3fhliv/F8dRBbDcVJy2Kjh
QcVuJYquJQYo21rCdlK8zSkMvKPD2+vRFuzJUDZejCaY53hCHKYzNSkdVvWoTZJE
wpkABhuqKLJdn7MACqGVaCtDr4PAjHIefdrq8qlubYPjm8MG8xuhNCtXztC/sQ/X
vTpCWpmBiv6YzWBcznQpPsRdfU7PwrVNxhaPtIPWw8D/Boroa8j605vWqdNWGDHf
8KC0yrM9cTpj5EYZiWlPTkeKMFj3kXRIsDMbjqFbFabgYb4FLC4V6CDFOZZOYo4n
26nkAA5Y8UJAcNJH75phY+Zh+pZ7Hv/u9AB3fmOMGVkOQN9p4F49kTL7A92uqBqU
A0kvIkw255jLahOtVserdUKTrnBc9CmEGuNlX2FlR1g=
`protect END_PROTECTED
