`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NGnfSnDXB5VI9towwCSa6X6lA59bFYf9SMDTGb9oN4bKY4WIes5G1uTnmagc3jQ8
C2elPwRfQHiYHZo4g1kpJhFSRElxIF3y/q/hCCCSyi9uwY3fGsgxTVNIytHO5ANm
XoDSdRIXMNjiOAyOlPtT2WHIT6xAeNssAouI1bGewGw8LU5Wg14XWH7Bh/6Uo71d
2KrrwVsOjLPAd15cIpb/4AwaQmfNF2lSPl6VyIgzStkwatydUn8arysZaydYy8Zt
vGqkvuusLWOZJfAa9FW9aulLHAIJQNe6LHBTMwy4vcKx0yRePoGtQfcdK2sLYwMX
0bjni4tKlQp+rKg1o+YRHKDbRz5c7XzxhEJi09458vUQmhYW8IrRwnjBVmH3X7cC
9rp6QOU/l7MxNC36DV/QOJCRjcJ0jqSm9UHKSzw3Um763yDzyTUJGVrQrwZalIe8
o1ZxdAy4D0cP6dSPKnfykFNEFexauIM/sKTKiZcZmMzy9VWvNpC78ziClgzWaLJR
Jpn/hC2GdMOwoBm2W3E5/WgwDhM66gx8r/AWiu6u4UAg0sea2KMwEBMBdEN7AeH5
V+RNR4VjyzZ0AtoQRnTMGy+lhV+AoVZaAmW5PzBUqnCfpF+T3Eo7XjldbIPWDmAP
1vy58e/AuxDnjJ14xBQ/8vfXp6530R7jVcG20t04xylwfpPApkV1TBgMh5klNlSx
DRD1nl1azEact5wjRynXyHPtS8eUrLqT8nW0Iz2ue6qcNO1UEUAhuVgaZ+zEB7pi
/wh7cS3lWNehSxHnehbb+T1w7W3+XcFw/1foGQNMUJA=
`protect END_PROTECTED
