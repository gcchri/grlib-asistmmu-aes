`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1+caScNlj0lTse0drtU5j9fW2YgySQS1e56bPOndIY1PAiJXwAX/jntUovsgorCn
ZObAE0AvIVkxSKvBBDav3mymH2C8ivqA3q52k8OWZinbq+PweoBa1z3w6C1dDVOp
jCuPhWT+yt44YfYMbBtsuI5V1+378MA8gV2fWYkrorkFcQMPw9a3zriMmNhZ738S
mE43c+eKR1K3MDtXj2SKlgN0+N2+c5XdFjWsUUuLqWaXIpAN8Ab/JczriL1UBIZe
HhTTafPQ42CeOtLcWHR7gK0sXLyYiwq6LVJilk5dx+Mj1TBYTJXhc2JVeRjAeYxW
9sCl3jDz+OYzUR6MbiRqTl9VBX6n7FWLppw7y1S3QO4JRvhoDpE9Fow4+U1+os29
l5zgySnTBaKFcmfamp0/6KI8t3zXUHOyvw1BVeE8RuzznoRiB3bQCny82Fp8tN5F
+eq2vY4jgPhbxX3COJtMcjcIkWKGxxCYulOjGl/X0kNjzQLu7+H0KgoiGgAlFu6c
hJJRtEaakevw/38YyZ4B12bytC9qsNorITss8SQu3ezI/UgQOP+/xx8opxBsB7k9
ojsWisiUmTJ2sOm1XBOcTPPOdhU6SjqvKT7xKpAAXpwZBVn/d2wipP+76l8xD7li
TbrGNSheNzXFkUuLcBzBvnSv7zINLMUBDQfzoAW+QkpAMpGijfY6c3KUGA10+omT
3B6SAbGdndtlBVZl0puQbUln4Um0wuZuZ+pZEO0y+hs5TJxt0lSfXaXWU2FKMhss
P/VTgZeOToS6f01gmc/7qXLmiFVlfJKyt76UiQv0mJYBN9DT8oUk82m0nISYw10H
Gnx93V3VR9n80JaCMvXYxd4yMWxKhafHQKNpaByzQXvobmv0Jd/nEEwyucsVMNl7
2gHkTZ5O+HxSziSpuEBOZO5z4AG6vpfPxDDIoaDGWTTdR4SIM+JM3WUXATJ7KpXm
M40taZWRwIhUDUkLv+RG9TL6cQOq595YFEUyP9SahjckBtdIv1l1YNY22w3OMyx+
hW4p+oiWVoMxp6w/BHa4AcIbIgMMyzAlMs/s4rAaBDODXAhvoJD4AIgbby5TUjBE
L75wcNNWroDuh6IQudzReeVrLd5CqkixQ4wH9/qvf18YgEhAJ0NvxO8j9gNqYKhi
AlsHAR/B995Alp0wzOuksJXtbSsjXL0uf/SBFZ3U5uJxzRcFBTJd1pvCLFFS3w4Z
Kz+PSJ1JGL/tdMhJFZp16+74l0IYZAz3cUFTFXV+mQXA7A5V+bKUP22nH6hCx1ch
L7V+BIDB1x6ouSQwTHVm/D5huc7Cgs69aPprH5sEuQQXMkbbET8GUYuQ2lxhD0KK
s4pCFiNvbFm9LB19ZMsSHs7zcOYt81CNPgUtEXN5voYZBlsEKRI0hYVEIdkFxQmk
KbAy5gRv4LPHsjR9blzcu1XR+bRroO31T3/6m4xnwrmJo/7xwFSRJ1hJYTuBabNR
kKrIbqTMooK2PmWB39EdCGU2U8O6w1/eJCP2djvCZVodEIbUvd6XZrBDhaxJGl7P
YX69Ow8z2CrFtiml5juqF8sBF4a8sFUMuBI/V4ZQp2FuNrFlHm++qxI0bmNSpUVW
Dy1htMUGacyTZZ3cZ3C1RqrAVnaQp8GapnojwHdtu9wjljo6L31P6mnk+AG2lt/h
WQ9tBIYzldeNVatKjU2gHMSXS+iQXFDDurj8VmoqKjguV2ICo+U6ZiA1MdjjFAgP
sigPSQdjRxcG/JjGBx+xgrFiaNtVWQSBJdvfiKvdeXyNAgUMJZKlJdkVIlH0sdRX
+bWh11XYQFAfbcuqZmFMEk/9bYKPGyUJxsDiRvfxHeEpFezyTHOKqc3/8mQAIUOQ
Kzq8qULipe6q13yD4TLXDFoO976wmyY8e6pqzJ6j5JemwaAFVvLpafAGrHHVaIDV
GrXdJINWpVw+Kvx6sSnljw2MZvORXDO/YDQwwpGhUvDp779ip/DGxeQqAeIh4dsM
42usWcHydBP5QEo/hjcQhVq4lnSgqEPQcmeAShFG/Be8oaoReL2TsiWne+o0UY2s
/uNP2aIEXa0/sYBjSoD/SehIy5GgRYa2bHXce2fxURjpvzynj/F3lR9Ee2MJp9s2
FsuGhcFCQ2J7c+DGBIKhEtftKDci3qG+L29+f/dhM8MCrkvRwGo/7l2KP3luh86r
A1t1+kXjM8HwzQSNZfL2JUYsOTNWHgc5cbUG7kSU2McmaD1O+VLvMaCTOgDXtpGk
h3jxtgAsMbOrHvGnezSsBAr5hBJNeKKcxHl+mjJbyFGa2td2xKRiHLI7CeRpMndI
gEzi/HaIwIbnI+Bj5maLHp9N87FooqfMUdnaTAroZgHRSac7G7wFeFoBM+QxJKa6
iENJRlr+2SQh05eB9QoVL1rSCma0fhA3fnf9hyjA2LlR6V5o1/ose7jOpM9bni9k
MbrUyeONx74qsoyYRnQ66iaAJAWInxfSKY4pNdfcv1rRCTIprK3tHTYGKOT+9+Nq
GZ6weZZLqgeXE6s8nxVbL06GAJaKXCI4pbr2Se3+sc2dInuT4jDMSXquYC4leW+c
IKu+WWW6hFoxfupm8xVehyL6tk8eiArYYvYt1KY/O7f6l2Q+DXpyoMTKUJ4M/VIk
9rVUQYrYP28tUmt5yfoxxnmMKbTMPtG8zgRxMLwina4YcemJPd2l0vJhiDtnkgcR
44Y0aN6ENlJRBzM1nvBjzk2lg/Svai4CZh2psM1xDLNzeLyk7K9A9UklInobFGBo
KkhRgHC32Ld13MweAg0hQHgFAW22tJC03azbf3rjPwlmGwjixSu0UgM5om2cCaSp
sWSdZbuakU6uGmrxfXB60mzIs3b94zi64HOz1pRL9GheJq6dXuMph0L5BRcdal4x
0m4LgyMZWMbLbT11b5WyznxYzbyLP8gDvGR6U8AjnAu7bVlzFzras1nj57znQvYN
6LD74pWfW8SFpJ3njROnP2viygSJ4mhTHhxTwC6jsie9Rbyh+Mu098vXYY2yyA7t
F8mjx2l6BkB5LpUgNHEK2He5R+wkuoyCoDw1z+I3xycseF8QdxNpHEFKN1/0nCUt
3J3jH88niGReNhHaYeFytmuZE/oN6wllxVep8edTwk4OHoLLr1lzEw9qUH+e/nmQ
/yXKR8RqUJwNkREgYLIVXKxsQMBEaeahGmo5WE94GV1R+sz7GrZofl4c6bApf6CA
wnNMPLkkkK4VlKC0V06/Pf8MW7j+MgSdrG+IjVYZzyYI7hD7EahYgG5WP0biXH7p
lB0lsw7Z3vNhbg92ymzMZsXSsV3pBDjoxVvASpm134pulYGX5UkQ7pou6IZgHgsN
GSKzzGPJqQuVcmaShoFRdOxy6ZI3oP13MaVWZuAAx6WzcvdNsrIwnrqSOb3GGbqb
ySFV/BEAstgUr1uq8EZgIByP1PgjKRtIOM0KMnHg7wudV8ual2qMWbjzQeI5CHYT
LbPZUwUBIWnhxrb2wYvcOXyDge6BAlZE67c0tTpQL76Etle10idkt1GzZvvABAfB
5KW2sLsQmM1jO3Ux9llqRvzfMGhUAu2gjgkNEDyfeM9bHkdXDyFvW03A6m2VTtJ+
azJ5/bpTQfS4mOlfIZl2eSSO/gdwDwMFtAn/VKYBzdrB+W3neKYeAG5QnqCP/njI
`protect END_PROTECTED
