`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
39CalWifbVvkzTlXKivGHPfLeqlrhSTz/FMNbIM7klrpp1rlB6/RlnGoY4pEA4RN
l7yd5divEPfI/SQi0m3xlnrpKTH83VMwoGDjrE/8bcQhQ/9pnEVs6C0A/1tpEqH8
20bsHIQiD+RjVK8ZAl8NC3wgO+HVYwgQzDLVFsmm5r+BKkGk44IJmPtUsOArV7fU
moE+MoUfqDgkFhfezYd/vzvSMgPhjThd/nf8oEmvirr/1CgrzfQ2oHVqsMHQwEP4
r5F39+w0WO+qM0UmAxK906SA96FipMBbxLWfVmyuEKWfz3DSMjG1IFzVoRKs0M7h
zDwc8Ko64R1GfEZZk+VpW0guV1jVGLYQVw5wJgySy74y9ygyf7QTXqTKo+CBK5zJ
3YbZ4XGvb5ZcWCLfPvo8+MkiPJqrFatr5lniGMR0slTE+NQ9hQXp8qKwmMo/Ep90
Y05Xd1cn+CF202qDOh8k+BsxFIKgIl+/xmdh8TMCszQq/DupQks9nQ8GlKymZUk3
sJybmxXg0zALLb5uFe8HzqHdR2W0sMxyIxsFgkYRKs7DoPfDt0LRgwd0yDe5NWwm
`protect END_PROTECTED
