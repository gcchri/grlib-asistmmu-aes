`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aGuJTtVjmHs1zwIuVDsaOwPJ85sqgxpdDY76CzOba/5yR5snDLxQfKqUL/sUv05v
eq3Ad9aNJrNzkqW5pUIWEvjEn5VK152+/OPOzWl8bAG5tuXFqa0gIQ/3Yt/mLIHv
a3iz0n0SEjCQhaLoWSARxzEVIZOd0P/Cm+df25lezpjednmR6ecbg4lfYXOP821o
ywe2Xb/sR4jaTemBywXg9rfRF01GaYVLy4sr1pZS85oJ1NSX/RnN8wmMhI8fCEbF
hLxW24H6+llXisybKyo9tAPcsW+HH65CdTYVov6SAe4ayIaDwMew6KstkOD55+x3
1fEuwvBr1BNkd2MG72UvWsZ4e3DD16xWBRI+YgHa3zq13+6PKTebP/UMdvyDPEGf
Jh4oc+fUGrGf289zs4iNNP5PWe5Umq6x3U5xvtDdwkU=
`protect END_PROTECTED
