`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5fo79We4wQeHs1jdUmgfP8CxDSx6rcuPPtjbOB+AWaGafPF5W+4jnWGu8nqibcw
OdAF8ueFGcaqBPzOjj85Yz77WrJO3Vv5issys2O9cgjI3+kqWb2HSg/XMcuvzOAd
tYeDuDY5jIZ5gRUSF99TPWs4FNbxQN8vPMU7AdtiuSX8zuY1FTziHml+CssVnge0
8g4WufmUgbLM3UQ9uw0YilO0Ev6ttV5IsKVh2CoRQ9uRj7bVTeorPLT0qhS9yyLT
BTVaTAx+CgdcZk6pGr3a+88qm4YJImfDY0yxO2WAPuTlVvWbjkwAg2nnIXeN4cor
WufYNDECJ70FzOdtBAQIH/MNuvURSJFxIIYvgCP6y9RdIkY0ZBFxk7MflqC240u2
8mJS7so4XEgQOGIoqpANlWVBTXclEDYnMg9UQuwtHbLs1pTUWv9nAXeUyztYRn5w
vGzlFHE1acLMyH5cyT2L9Xq2JFhpLD7+fBZgeSMBixQ=
`protect END_PROTECTED
