`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTQEPHyODawEKCx9O3vUg24+cZF/rG89ntjDZ+MLzWBze9vgIazQoNme3JnhnsS0
d7y/nY6tjfz/zGIT9q4Dze70y7088876ctnkc39vObdZJuR0DS0B1Qv1mTnQ7EP+
fOnVVl+f4HAioxhuXCFuBi4gblMH1meTChqAzuPnZ4/3mJzMTTjijlu/W3z4jSYG
ofYDLJYTZF3UCMC+MpLTYNJTBiYHLMKyZDqPsRcodLhVIK0e+9CHRKHfoNrXHZtk
1tz17Qi/JNcLVS34KpZ/5wNoo0R0dIQ/8TPjZWigIu1EOXF3hF6VInJ+PSXyTFnJ
1L9I6TcqDel5ZBW34R2l/IxiO87TOmh3iPW0WQkhYWbxpWJGZRFmWVRlJ7u+3hyl
nKLC40cWGSPkNMY65xio7fmwbwzwhFQASeFDIw9XzGUzb8ho1HcULd9d5X7WgsgC
tT4nfBLMMgKD9m1VdJflHA==
`protect END_PROTECTED
