`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LJtDa2kUdYfnyhnfAg/p5TAl9PSnJJklBCSrUEOqIUqCwki7+CxHfTdfCoiAOsV6
HZaTfhBUm2r+9f0Uw8GmbX9DOC1ksOPt/trAk3UcERKOT0QkQBT+JVC/L3Gy3Cwz
ngjr+1Rtu3KXcO7HWnOHKd9l6R/rEpyNE7219fRgb1VHcXkfcO/vSk5QXC9bvjvs
Ao7qZWKcqhIcv4DnjI47uxCWZVP/fG+Cx1b8Jta4i3ItRFyEDLyvd8TWOPEg7hQb
0Dx+2r9JtSBvlC3OjifziWq2JugSdQhhCYLJYwz/stL02K1BR+pzHBCQayfHvPF/
nelJc/DAAzcV0C3BPXmy0BjJeyWXGvcf9lgjqXENb0NhDT6JwXNJSs7lR79J/fYc
dsjWUEGxVCLrErUHQpH+5MLz0tt5mKshDx3TEqtqTaKxkVOQyGCTI3qzoo5Xa5Ct
QfVwwtJ/ADG7t7tQBrm6hqyguaBljF3YjzBKHcbxZeg1c3kqCRO+pJnQzCOjesMn
ZV2bbKOJeR+WhcW5+zfgLlp89FKPA9Z2IVhRErd5fPms6BfQVwOCe/ezp2mYBx7A
+kUt8BE+RwwxNYiSTCG4YqMUj5K9RRyWKtxuQ9NtI+5Xom4pgJo3guIdkTB18kNl
Hdz3Zv0oSa4yer/We7M6tTvhdlbDDH7fe5A5g4Y96wSTZYQ3nvrFJv/+Hk9RxxSO
ang6kUdppHXCK7bnwiGORRSb5PFnCj31nM5kIJi/3DRy4BaIR6NLq8ZetdG2m3n7
1oXFOupZx3f/5mme70Cw/x+ySyJaHCP8o40bHWlqIOxRevEnEGpjyJ4QsdaLnYeR
TjVU50ClRW4NRvEnfWXH6Xq391YsVHnNWkq86CZmn2Sb7fRXResmOMPuJ6FmgJn1
RZIJxQx2nW62CPLFoyTHjtHQzUlCYIygmI+SZXaMvw+u/85impXDrbEeM1ZKGpHk
vWXjGgYWlD7B3LgHsJTMNIIITJ0J0EfbppH+ZFqGgR3FMHmq2dWimgGD9gJ5xvQc
I0h4G3GuxXw0zpJsl59UWBRC6vzLxdUzTNM3esday+kq+iftPpth1lI7E82onv9z
oVZcwGj3fU3vI3xSKPdzM3HUijrsU8870iozuXRckQyDCEdO/J3PA7EA0z56cgtM
zUVOt75zuU0GkvqKccKuReto8c5XNgtDZ1YAuXdGNfjDXYXLk9lyvspdbq8g/+xl
iNEhUYkDvhcBelGhHDuAg9AcAEk8P5yUFI3KIFswGWA1ADIkmpfPdX3UKsLWioDo
9mUP06/6SiCZnRUBoR5CZ97yCiPD27/Gzj2QvNtlAYmCt6bQw+hAEhwTn2nRwwr4
ErK/3372qcw8kW4yZcnRnohKTyXQo43/Qw4b+zM+2ukCwVUGAT9duVQoew8bNR1T
L1Og36yIBYvHSNoRALOT1EW+NFAZjL+vXGu17PXLHVg4HJsXzmTNiIyqAPa4YIKj
Eo+t09WO3ghK2m9kDaGBHzYMTS9c4ZynwrqWpwiD0iMbJ83APIYrbqyDnCAv/dE5
sH2W/hvkfJo8EDN5CMRqLbwJ9TXVAMs5/2IpRAouf6f14KXov83gt5HtqbYTKbEd
fJFFtFcUXbzs2Qv6K+RQOdlqokrWKX8tXa/w/Q8FEcnht0HMFXwrDrfsQ8Ms5eUa
mn1DTsNZsncAkoNvygBq9k3gb6kwaE/HTRgwDrXeT0oqeemFfcVv8fD+qjWsYSCv
51hC03zwpM8Me+v2z3/XCLlNa9Cgp6McTc9BXhnw7fVOZ2bdNF1GIaKOLvPZGVg8
rJWjwWV5YnvQxriBx+XU7PJcD0bL+rMcMLtWMoF3Qn5p8AkX2U9pkXyVwTgxGOVN
mI6Wmy+g7t1qUOEtG/6AKN1Bf4HD1tllJFCp3DcLjlm4cgEjfvBevNVnGp3hPdnT
k3X5bXcHIC5Pwq6FOGYKXrxMf8oX8oznBxGIam+G0LmHBKQaYYXhDED+vNJJbcpQ
qcEm+uhiaJ70uEVAd3fjvNDMYjA/t8H1Jv4CSAx6t5KgZ0lry734Gpk+zPmTnS/h
Z7nNfxu9B+6GiixQq44gL3ECnJjQlJv1vw6MNfcZd9lEEF/1CusMZFc/uF8ucQ7v
1RMd9php1dr8FXOUFJ4UqVm8A/z6fUS95woQIMYJCJYnI6XoVWJ0A48gQl3l98x0
VveJCjoFsGOudBdK6CZLSDLXx/NoNrzKaxcx7NsBXcWEQPNOkbztsQoVrhozcTOV
MNLiYtNfvOY8rrWE+ml8/rbrJjA/c8EOTTitzNPsfjc3WwuqPtbZL2YtrHzNZVSQ
5Z81mi7ZMZ52oVdezpW859DRJzfDgcsccP3ZyRiReD9gtFPAtTRUlvMGbcWnMCux
y3P8AJ75DdeReJqn+ZWznDjrEpKazvIrc/OnYo40yd5hXm1so2ZsbayAMT7posYX
`protect END_PROTECTED
