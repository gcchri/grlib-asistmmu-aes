`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMyHuLNpV3OVg/iQCbxBWPPPq+tk2yAbbEA4xWZSPArFS2wqyWtWSu8cPutK7mqf
Z2U4H49A/lUJFfxi34P3qkcA0lRqD+b9/j1wskAXNn2NMLwPtg+qBkAfriL/+YPK
SqO2dz/VHYrpPsw7xnggTA90mwjbRqxEQnLH2VD21oNQGO17iTkdOGQ3CAc+I4Mx
aBd+oqIE4L9vBajGFX6gxjEHGi1dsdDKJQCxxbJe2qQRAUmDEmCo2leTeT7cWVtx
pPIZBQBO2nE+4A5CGU7aeQRfRsEMVc6rVjVw5b2OHcd7O+61cvgYtFt5xkxKi5TR
2I11h4jG2/iSrYyPipfU6aBrjVOvzaerXHLJgZ2kIVgPIOV7BbVl8keWJZWNgVUm
+8IwJqCfWhBI5sDmxk8Ucio00fCDNwhmin6wUeAN/iYfmaHyeX9Q3UiTIlmJ7uhK
r4M4n5hmats/jiCcIQ0jsECMAXuG09S7SwWZqS6GxSZh2L2q2e1noZzImXaE5ysX
eaA+9O0Z7FA0lA/i6Ws6fT7Qr0WGowu/ewNqwngD6fQFawgnFaJelOP+60LTWB9k
3NdYcRejrd6WVl+JGiRT5XBfBTTSZt0K6G9nMlPClzLOajX5KLrIRI+Y4wm/ooeY
JwNkGji0BIBUaceEV0e1L7JB8ry0294pBwgzD7WJXIQqoYXwBoLCvD5YVns8/9cA
UTAnhdRdXbHTxiTLSK3kBS282xWj/Q2O/GVQwcOi8mjwrpteYY/BY600eePzU/9k
dyWyZp3TQybjOCMP3oeMv7tw5PqSUia6b0JwFGwwdrSXeG0sn6Cp0KdUdX6gR7fx
S5goIm3eKyPFHeHO0W0YLxaD9Fs+kRF6Pzb5cx+A063W3PReLhxRyLM3yv3Xr+cZ
fIgpk5wN4xAh6ldYb/wa5qO4f9MypzpI1qOpokz4E2A++2VoEafDYY16BOf7rXpy
32iXUj+9nGcTmOvhmTKF5Hb9KkRHguOkwaXJ0RQcbU/1qI7rYj++lpSFsWGEFx+D
`protect END_PROTECTED
