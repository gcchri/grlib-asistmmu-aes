`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DP7Yh/ny9fnTqRhFrpvubz1uzk1iW7G9gfTDSnAGtEXdtHc89Y2G6mEsbTXPfA5V
tDllhBRNVHVxtNc+aWquCFg4xeaNLjWeBuRM8zULDTubQlo+7l9chnSXv+Md3kkL
05r3nvCTsCNWV3nOdmRdDuLAVhxdgJG/XcAlmF8tvqvD1k0xsQf1BTmerTPW2/aF
VhRF+17WvMB9OibWpAuO/oay9p27w6fPxl/Z8ghAspbqpbJrL5UlWHu2yl+4Argf
Lu+OSaOW0xHeAkpwhw1DGtFF+ZNrQCYdih/S5Nl/8/76fyY4dJ+Cl5B3KXGbQCHg
bkozVUXG5s8Qxlle+/H67wE3kZZiA34vmqlHiFuWIROIGAcUtKqM9sPg5vL15V6S
n5vFdnmH9iaBABtUNdcoeLnVcWyWpdhRGA/BIyuvjIMnX9iBn9JeafirNq5wFjfD
Ye0JXexrv85caKq4p1oeak300jCumNntTCvzjV92TvCHmH8vDnu7JSYq5K9mmqIn
bwagRkLzYiEgeoxogXQczz91YeJV5qSrwcDXd8xZc5Rqb5mUXZLfXih3XhoYZCBW
a6TQfNskzxO5M9dZcF8QVBBcI7TIAE2oGbv1gGj9FfVyOkPHpauHnGYABSr2GO9K
GDf14jcPhnAbmsM7LeWKFMZ5h5KyDH5IwMc9JUk3n1WxOLe94pJIzi34De0DqFeK
LO+QJM91U2TQemL9m/kdsLQnF3hZCt2/rGSfcQLgDo9zx3g/xtIDFkveuUtVlbfs
FsxSbcjwaXnipBdQBdDYnwrnsM1BrKQKbxV/AoQrDiQ+ZAQVPBwarBanJZ7ja2zL
MLxRTdXMm5ubGtZFxPFWhdyBN2zdFmFN3EjsSPCcrbMBi1Y/X8UXbJEcSn8Pq0nr
OPnXkf53AtaX+Y3AgYXYRwIk0Ypok0r+pAoxJlWN1d4SqcqI1JzSfKS6pwKKICmo
oPH+OB181h7ed6kVnzmQKU5LUERA8UzAigZyWQXsMkQ=
`protect END_PROTECTED
