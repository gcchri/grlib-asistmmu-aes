`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yw77YhRrKQddFqt/00O7UQ8nYsyJfeLBR8bbQtIp/OExpK4nfM9DKAuUljZOYNyK
dL2d4Bs1k9rvAYocmNnVUNqYhAuz+JPHbnywk7c14HzFd+umJ6BOlhPP+LiYrWet
7u6TgluqIstskrsviU8STtbxEAYduGMhCLtgDfg9MDhhEN2pTA9fwV6bvC75wKlO
hyO5V8VJ7STes+LUIBzpIonmG7+tDDu4RgPOfWUZ4YCvz0NajIm2ZGPcf0AwbmEz
OecejPMR91aLu1UHpkWCTi2rw0twCjgZaU0OEEtLkgQj2vg2f1WF0ZzDM7pku2D/
fTdRtLs5eeKT9fPt/xd3p58lQJ8xg8h9a2K6H5VYYoFjb1P9xGx6VbcR0oGVXyHV
DkIWtGuo8EZKuajlhBUa/JVRaRTp1BOQFM2IS41sDGU05p8pKhZv6/kN2R6E5BJL
fstUCNVcz3V5iF5Hrm8ZFkFypGpInlxiUdTJpyt3Kdm9yRyO3BDXvvU7z+8Cgtb/
8Ot/axE4+QTbyuPn06XJ22MumdxWa1BDn+f6KKkndKMRCkSemgoIkLqI1uC5vHvo
BwBHMSYTBEzRlFLvF3/RMG6o9dNNaz0nhxhOozlGpIqYU79Fu9NR/gdNuJsGMbIN
SbXMNjFxJ/m7TPHOMEEWqahpna/+NqN9XGKmEimUq8zVHLq94QmbhOdFHYaIjiyH
NypEXVsucbIhV2FiWYik1mk+AW6LTcQ7MtQayW9ClbM=
`protect END_PROTECTED
