`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1u5tu/QAwVdNd0BoJO5K7yCINBmMg3rUi2uuzwk2WWJws/XtuH/aCsIXJjdifDVx
CD4bkF2IbP10KW0hnYr++aIxpwG/gWt7lZ/ZEs/UqHTBBMYG86raWlIHN7ClQ9qF
ut8Loob5xA7LNzwV5Z/uyvi5d5D44oz2g+GLyAYwmEdjcM7H2fpLaNoh+xAKwYWw
eVKixieytfj7ZRt+FNftyUgMCnyR9X6A8LvcblSZLftr1baA9ynC4xPahAHTnmqS
Ajcr5PhOVx7B7tyOGEQwPy9a1AvXSJR+vUJ10KcF51qtofBjTHUXdjVTbcf+ua8S
Ia9lNuHS7/Ud2YHc0JhabW1vf/sGQ8E5NOcqCQ+iPbgPhThw/nB6/nkDFwH71hvA
3UR/rGRpFgBwB7BZ8AYNbSIgZuVy6ArB0To0xYXKPTen5v7e2gKTNAcAjcVAdUcR
v6Y4xp62/lo6gq3aSzFQHGQI0NPwel55wbAbiKyo/35pUgw2zhLi2AlsDlWFbWey
qmP8xQQ1kWIgLVTjY6Rs3dm2+8hJ42luo1XV/vV8Rhp5BC8Y391YDi+TtozrM9Im
ePBdLE4cZW+WmtQUA/gksqp0Yx5wJZusWktXNvU7BM4tqMwNBOQSDKyrf77xh1bp
smLfcZ+EU0Jy/zevd9lxGO0NFFRYlArJdPY2Zr9Sw7AUIq4QPmQre1Ee2X2KSRDD
iDaal6DTLJqrz2p87E+08nLIPZpcWmgQ0xb9EkFl7h6U7Cs/+znrA5mjT9O37iU+
c9+ZLG9JjKDaFiQPbnWEbT/+u/CBCq/kRlVB1bOsK+TitxhU4nCWT2cAeyqGt6eX
DQEf8/PTxtUI+tmC0dmhTVlgh2SnI+WipJadJBYM4RTy+APv7XSOGp0OI6OGlg9d
EnKdL9aziyhYgg7LyZFZAh6p792ycLl1/i8q8Pfi6BfB7yM3cirW14iGqx3VBmNV
ythal6lr+2xquhWvNTQ6DpXak4vGhgCg2KM9tLrVv2f+SG1ah3KCdONBnuCx2rYD
rR3H2P94Ihbu4wFX/nYJLXj2fDdEJuozErDhtzsrtGzqEXsezuROnf+2yF4R3B0/
uYAnwSCnFdDxlvQDHXIICxWSiVrhGvFWWaHYAQPHXbO7as9dKa4DQsi6z/K5mcL3
Mv73ni/jfMhREw/nze6uqOvfgbZQuWHtG89Vmt31k5WXbVuOwnUToyqFgxRP253W
QbcQYkGIyw2CLFPK2loMW5IKphNMzSO/CdhnzEYtnGyIdvvr6AQWqymEuti4LRQ3
jIBd5xWf+yrYXhRUEWmEpSA+zyvm9Fmogs2aS5k7bBzIi2SZsjycqWnAX8Y/uYyo
m+7NsQygQWBRCysruF7O/fT1pHt1lX9ptbNW4rcmpLqSGgap+w9VxBXI0zZxsQ7g
hCnTBCPgk+Qrrhd0JzFrpGVDmnxX01DDZpUg4hKFZ9GzqaszrKl9aBbmKQMaWiao
491wCuWtAmgvCNyo9U+CZ+EB6Gi/yfVkvR5YDFG2TNoy8iTF2nT5W7Mdw4rVuyrN
ttOBfviH1yTvb87QHAkwj4vMButsNaSWpRikk9MpFEh5zt0dMPUDwL/kT/rflUJl
/ZZNq9LNnfyaB+8A/pZHJAEl8FSpx4thMsgUu9F+Q43psH5iWkigP1rZH6GyJ1Zb
EDT7k3RkfypHIyHyLAyT8HvTovQZWkD6IB+arhnwHJESf1hE5d07cto2vWVrO/LD
/6uEYc0QOOWsJks3xuSMe85/kMfU1+YKgOOmIvPrDvmjYYL/hcDO7gHmqZDy3Fk7
4l58Y91LRZdo5fJuKyk6cys5WlnY2opPGJONq2mYrVQggH/3hZUWjsZ+f7VWtiKV
jHgQsmpClGbcUGIMGnxPCNNZux4SiHn5r6WZVaFpOHJ/sdtIYerfaD1rhE9RVOdG
qJjUK93IeIoV+6OFzVu0OLjkQvlcYXbdVFooQV9pzEaPf7gTK4WZTiqr2yhdSEIw
h1J7PGJmrUqVzlDD/YPqjqICw243M69Ax6Z7iedhJIAI4aQbHwZsCeW7w+gWnLYu
TnVniyeYizaaqXi5YVwJN0NB8NftaYi/YutcIzv18XKR3XRsl3tOtTRjf1g4o7Oh
s/0UrAkj8F85C3EypLjvTVTvi1rouW2SoKaVYb8S6WQbTrV7WXDuWorZdunTWGI4
j8Ki+R66DEVNUE3/zGHR9ubmi/KT1WMyewcOp4/uOqDr5i6oO6cTiuQlrA21fe22
/ufZpyutm4bSazTbAvO0viResv+me4DtwIUwWVBSbLo32ybLxJm1PLzfsQMyLqgB
4RxvZ8KKbWjugTVW1tKxowqFXhfmsvGRW6KjEfTs3mfWblqBpQ6ZLsGt/JRqSeM5
k/SkoTXElJ1XSzimd0gUMca7aywMjFk4+RHk3gkwAlOQU/fEvurpA5DnqF7vmOPC
lVc5hnWsWKLPEiWDif/uJYFsgvyeoFu2i4uP//fMnTYgFe8s/xThthAOv6CnmDiC
14vN0eBOhtuproqML7zP1nqhcgSYAfYKGVR5dEQNOY4aFOWbGMAJ5Oz68rcMK2xn
Vp8HfAg3xfI8YtWdHPdaV4cNhp4rCmbeTNKf4kMVb/C7y9cUjlh+mqaYCsl4vCaJ
kf/gPFKnhEOYnAGGXLTlGLj+M79/pn1BEbXcnEizncr+wepd81wwaGZUt5vk/D3z
YyhrCTAxuch2+Zlw6r2Z5eQ5Xg4cKWD4u5C0TDoHBO784h7NrRjActJVw6oKKm8a
uo6DOr7Tw261A2R+Wt3m3zWnkfPf8XB3QB4m/aytpgXna7WHt4eAx5RRttQZ9vKa
MZPohGEyk+DmWBBudT5ZVGzvlo5D88NGFJOnuCB9wrWZ7GkW6Fkt2wJYw9mcYaiW
qzDqPCimD3nl6XKfgbfo0xQntRSlxvopdIiG10DcZckuqviax6NYoUCBTqNr/Jb3
Rb9kqZKgGAHDzjkrgRmaFSmkCf8QuW1/D1XCc5OQ/sVkKA9hs/RwejRJirfc5qwY
rsaUlzsiQpVCeOx3s4JB7CCONjO0MJAWJfZRbbfABACU8KcaqPxXT5ueXaT2s5GV
wgc0Sijmdoddx0Gq+8rqH/jCP6D+OrxF/JUwRX1hQ3hUWIdf09C+q1muc02+I/fm
t/YvejQs8o9jqS/82ImqKpHVl6GOuGrbXR4bgnumV4bYLef4rnbra3Yeem9N0l3s
nfE+aMACIE5Lz0yc2kmpZHqCXbIBKoNflcCVgSu0DzsCzc98Oq1vvoViFP5TChQT
6LzHQAmFDi2ssauO6tj6ayOecinAoEyvY1eje4c3gZRQRyDGXec26vFXaoEUUweG
IG+xGTF1szIZoMQjr1zzxN3xkQ80nuKhqMjoPyYtaXckBCslWcWXelaDxSByTEAq
e4tiUmy5I3+GAjb3EljOrs7wFd31xSivS35i9T1Z09p8OKidcO2dTDuJi/tEZqrU
cVjjpd29NRWEsjvc3g8bdV9G2K08R91mT4qVzRJtSP43S5yFtjvC3yrNAlLrc48L
YYok5w74CDppBlSjlCjYTe3K5gA4C79FZd7fJ3RVZwlEeTt75E41Q+MfsIzSUa2w
ej0gPD8JwgQw3cwdLcBPjlg53pvLxcKDEtLN7k8Ur97ByLadtD+hUQeGOUSIkVLD
KVEeSz8HvkywXaFfGV9GMmGE64MFtRxSir1YRFZ3T9vWGMdbzM1QXveCs03Ru6En
nrrQeqSm2r211RYSJ+ZAO4rEaIw76uN2gW6qpt7klTPt1XAsBIOiskd6dNGuOxco
Wv19HX1FA7CrHEzrkaFr5gS8pEzYUbLSU07BpS3WQs/3V0GWAgfMiccKv4AYG5ZN
gtapGMCpNSjdb2Jr5p1pojG6tuKfYjU3noXWBNvLUkwREenTOfFdqfXx3LQ3WOpg
i8+vKrT1XHBMLOBJUZz7Tc6eejQxbX5RHbqUl/10cywfEkGEO2Np+31MbnWNBj2v
9PbaPNA8vlc8ITn5SjKuOvjC5ZAc+VWEMT2FcBjPWcWdoBktBI8K7vO31iIw0ZKV
P69CoeSHV2LKeQh9WcwCdGdaeCJyupnlJ1BSzNAEzQ6iahNqkROT6Ettsi9N7umZ
T+2jCw0ehOtUjkY4yizS1z/QASv9oI+5MBtFhIRxyIhguMIVk8+KeHvUjLig9S+7
uIcsGmj+bVlKxrem692U/j/wVin4az/krxI//D0Etk7D62oZXLnyE84jt6vS/Hj0
y8n98h8vliXTUcFBJR7RhH840EVpWTVpnSge0QDn88jbQx2iU+za0DxAdazlPcPj
e+dRqW+eW+pDYf3dzt1SPslLmMFVa5vUgLrEU+Nm3jY9BmRkpF1c4v7+poWjEM8+
31Z6aOmPKTwFdIpr1VeprsGZwast7pe+tHEb2jpX2nsEdGMrmUGUMtrqHyUmswSt
oCANij0/hW0BJTNExcCW/8q/r3E4WQuTCy0XP3ZNksiWMDp8Hlziyawf/MXeaOm5
I4kkqCuQY3lv/71xrcjIf0aEogiEWn75BRW0iOout2M4j4QLo3tZWdtC8KMmQIqN
Nn511Cwnz7Fe02Ta21JHEp9dZv4f6lIrwNg3DZlG5vRaeAjfuOB1aO3DYsMoEgAu
5a4cS0OliJWUaM0SqfsVjZkg9czW7K7j4rhsSQPLnyXk3mtgr+HtXf3BWmAqwDdQ
UtHllcdt1tUnbkrtNYyH3U2vDGI3qvXgjYf7r4gkW9awyG1COLetFOeIQv6TREFH
la72NfU/dMJR766+YGuuFPzvpNlFnwVCGJpaBLIITB+LnvEVBkBBezTk7/9dIS+L
WZIsIiXwFcJdsqk4aRh10RlC6256S4dyJoTZ7OMd9FZJpbgm1duHqjVCUkUvLSR5
aUrCa7gaZoC3Ks0p+Z0yG4muTzkgibDJ7eS5PdjUm5pX/kA/OLwDWv8BHcy4kWOb
uchouKAE7NQppoI4/NYoII0Yo8YVN8t/N1XRnzLTLGinpd7GyA8oUQlCTCJz9Bzq
To+KGXBQAmMD/pujO5n6EgWkLGyJaHIlqmTxmt8na9JuFS7uuTY1g9l9s36JCf6a
vaxkP9Y1PQecMINuiTRa25Cmbq84RbnkVwQW0IDWzwurkDFP3ASTW6+wudQtQO4d
b9Dhwkl5yYtEhMUMgG9WOYrycdPL8tRH/JbG2/sL0GRGMy3rJ8v87tbuJlZUeEs+
T1urLBlhnwRVX4ZFvb2QMbJZmzYRS6MFG3yI3nbvThGPFKphebbZgM7UwG7Hu8vT
9NOVFQW7HzufkS/FdSLGxq6wuJduUvpCyBo+HZlJ/ReABd5W+NkzbA/31JxA11fC
dqi2+WkMAzpbCRkkvqRKPZDqng3VUsqKG1z1LKiqNVRdvvSjrpONOTfg3Rj7YFpr
nnID/4PQiY9+DyUuOHldWhoMJP7MCzOehVTkemLmcgylb4Ztiaaue89/KeUEtGkX
KgaBYH5KBBDs6xfUNPi/CRbazQKeak2xBkQULHxQs73YPMl+t25BxmbzoX0mUM4D
9B0r3XCepTkUyEuf5AWQBX/z9R/5Kt27Mpt/durirnpFN26aSL8L2MiOMuJjwGBD
3FCmtVVndilQkGR448w1c1Fpyrr6Vx9i2rqjjR1w10O3AeyYVOv+aglbqSi5wQ4a
XZB0/jIgm8L96ixM6SdX1pydByc9Xb8ecvkh2I120+rvkZM+DxocqEKdAvSYhuyi
aowvBEX5DIElHHhEY705OWbJUmq7w13tKCWDJNgKVpxFFLQjYN2uZTHimox+cKKj
MfKek7j3Zem+Hm3oBEf/tDJLvQ3yq2jY0SzI2kg2Qjji4VsVJZqbK8IFkcatZgmp
xN8LCaj4nAawehTNZK0z4QP/FOBcga6XlYbrtrn8+TsQjC1rjZa7d1mxyGcQIK19
NdK7OV9mx/Jj8YHgDptH0QEXh2xtmzItTt5hg4uHMiw2FWgX6tUcQRgUMNLkpHmn
SXSOT7H71ft6E98QpBXVe/tvAPlP5EILbl3WfyFekNNz8+7APXTnU5nmleG6qOmO
Fyxq/yOeQ86uNRVmdmeTig0dRuTMGA2pP7qELtdzcq/W08jd0TXKHIKpr/IvZD7C
WkdlN2dbBEA6JxtAc4D34cN9xBZ13hO+AItaiunQlmOblDuAVKmFKOC8rUyymRUb
7hsR0GaiQ7wbHvWRRTvRedbJphifPvI95iBxBnsjNi5/E35+0WYgQRo13lmeJCes
QTaL2cL9JvcB/+PSKtC4wy/UQWeGr5gqhQpPXjA5890JE9Ewo3u9qi0oU+i3sAkN
tY2kjifGBkIVYrkKpBTULGxSXh6lmsjD3Q6tkyWVZaaEaYl+pVQPYFuheVn46+bA
RVno4VyNKO79ag45LQuuv6+D3bXvpV1Z9bpBwtXLNbAw+1BRks5zj+2xSqRO49ik
4vO0slBx/6jt6qv24cA4NB0Z365nqVOgNxrqqINDygFnD/jmF+kLDgU5a1aa21+J
FQts+MaRKuVZp6q0h82R/mONrKb1McccY4+SJOf3EsewFlR4zZwoNY0XGKCx+wrd
U3qssoMWNZ8xrJ8ajvOUh89hmogu8tQ+i6GLjuti7d2g9uXDCA79gisAAYxb/Ddi
AEsPNMOmthhnNBzmyvgwBHxUiCj4vSDvE3oPaD4PIUXRlC0E3zec8XWRoV6+sEx2
vU9lMQtjfmupFJIJV+5xEq8yuq29ilHKLYv1BL+dJNs9MgIEs6HkkNCmoldQEwA2
GKHpzSTD+VN7pzzSxl7+S+S3uIdNUsK6XyfG9vMVZwA0ahB1Vunl16uec0CpGRha
fEZW6750+6pS0j/L/uOTwSPwZzt5PDiC1/L5Dua00z7MeFYHNhVXjS08lvlK0GN7
JthX9/hYSvjfmaa3QtMLmLfNoo0lB6P/JXuiWkVLjfhkXXe453FTwogmhvuX4exC
2LiveNotsr3TlL0Au/tAeSOPj9VsUwwgiFrT9HNstMQcFoD3VycC7gqXGuEEAdkJ
aIDO2t06hqym2T4VVEUDRpedpzJSIjEF6T9IV3fnxLMDFHWhe/PBQAPX6xBG4mE3
Xd0mouON9BWfmmGa2ye/ylx6IOURTiwikRlpmAga/zraXRY1dTYVXPh3WkwElmtP
ZzURjO2/aD36gVp/wPsjdswdE0X50dhJvax7V1oxjixRZIO9FZOYfXdscjcfYJ+r
WUTW+Tv52JlhYNPiS/s41BQfaZlSZz+NydrCbqhqOyyCb5QA1qqa/4w7WN7lEPdy
oJVNNxDimWMBN3uajNKMXrc/vFbp2tDEGrdIVa4Xh0PMgvP8rZTsiauvSCj5Lqtc
y47iYOzHxFxCXTVaFUC/eNW3Lu4KGXnehKUOOXcTxTWAUK9XeReK2L/7JFu8QzfH
Hq9q1DbGaebTwku6XO7K35KD7eWlhANRfKxWC4KQq3wE/C/4o4OAlYDb/MlN/rGX
RxWLRDJsITEXxpqZ/Q7NN15UIQIfKOLW2JmdkNqpadkOEYi8vsb4lEexXr2pkr6I
6DvE78wSiQ46m6uOprHHic+MZAq9FHLkKqTUzbkG5IY=
`protect END_PROTECTED
