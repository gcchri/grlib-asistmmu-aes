`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zdMWwWs9LLMqbXqAM0tdJlnbp6fQilT4x2gzxwcfwZg/87iYerx/aQR0Bb6/e29
QMpcQoW430q7sJL3TIl85rqMG20eddm51Fm0/UP+2npkkjwpRT4JMMDdqLUGHw8K
ssM+wDYrM3yodAirfj+T3rgEu5h9+xdDL2BviOl2rqDXXo4IMg5OywkHi0uPuGip
O6xypu5/hoBKMDXDKlwyTKjSSMTaOrFVTCg+hkErV6+v/VpszE+BU0rYSy1Qtu/0
biOA7iAuROC/QSu0MFCKvHeEzIX3w2RA+AhrC3/2MnDPNrUJOxsA1CMeCRMOhJIH
VMBsy0KA+4ff4JKGpY/0uvCc5QKTqnAYnjV6Dv1+FJpYXhxfKcms5BpiYF+0cQ69
1ExTzMENzIa8mgMmsQV7K8yC+x0mS/hPdnH1e2Hl4tVQ+lSh38Wyk1vd2pY3J4E7
aAdK/uTTv88iIqOwAKenKNYR9pxhilBPqUftAf+Dj+7L5o+Q8/wJyCYTcLv59e6/
CGQFi+7ckBT7kLGwoPu4f0CXC6ZcW/EwfxenksN4V2bUsOdnUu+PR09wzTi882oc
7VcWdTqbGxqCJPATfLwhfzfYIZMoBdiQRwXvqBp6kkc6IZ8ksxIF2JRTFTJGnclq
5YRaaHDjiXVGRgwPAUO0/Q==
`protect END_PROTECTED
