`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjeTrcARgJqc5J0Nd/lgrQ5IOGgwRiqed0uv3VAgotwfwBVe9pwX2gCvee+/namy
Ek+pDHxPfOTeaeaKjZXnEtVdpHbMKvIcnrNq9c5goC+nd87YI739jf+4mNbql6Z4
OvvWjDk5wcXyYiPYVT79SNyqi5xN86jYxOH1yBSvQEvuYKHwupXNjp7NsCK5yKKm
qKzSWEKA0PafbyBvMhwZ/w60ZVjrISu8RjBuKP1HBmgwIrq182XFDWbKOPQQ+NOF
I7MwAa3Yv9DyrOQIGX11Gz1z4/VQGyhXDtCYwRzUBBeqVJ+eDZEaAkHgLNUEc/4R
MMww2z89bQ0WUqwjzgrukyb7ky7gSMToMNpGPSs7ihiTsG/HaO3km1BzIhg/SmOj
0bIzmVIyIG9XByHtD8mX1Ia4oqX9cvELetk8Tw9nnVoDj5qBXxhoRvlkryeA/btE
`protect END_PROTECTED
