`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTppIy+HDGg4i7FJyLok/EVrlTzQZB31mTAQuoovrJ0PWtIOUZbG+GtWQPl4ZMwW
Q2BeBFhLRDpgMno32udj+O8trvQdtJg+1At+V3zkqkTTHqunKd2peVwmDml4rm2R
pLugkOqBJb/wVYulRWeHsgli7StgQY8LohtSe1pSEluKTzrkgGgOGSTc460Pskp6
F5oIxQBW1NYvIisO2HooN+sE9kRE9FS8TreGXWcw+FfMvu/v8Jvw0ea8dULJxTzW
OkCk8bDbFCYnFz17ShL+9tHCAMFLi7eyRfsoExcS3kvtKIbtUQFHuBywbwHLxAyz
tsg04f/iTqQkeFSzsboKT0EDUQxAdR75JFcSkIrAbQiFE185SyCwDv0+7BQoQbkF
70S+IlKYRqEaLPv6Ebvm5HiK0L/gs0fAr9YsY5GRNqHCE0ivYavhJMY8Okf/QZvL
ikA/M7sGiYACCgR16hPPfOsD0A1O6lflUOlx+j0aGpQ=
`protect END_PROTECTED
