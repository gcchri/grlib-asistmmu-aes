`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HTcjARn37P8EJzKMI5bpRvY6GZek/6+xp4e+b9Z4H8V4QlTnJvTfGZY4TSVhpTvg
1Ecd8v85/3kFkXSudg9tUYTxEGuEdT2K0FpKaayKVb42iLSJUKlN6zD6w9sFWhSA
Gg8axIsegCFl6j+y0SYKIry/1KlAksfdUFCZWY60zWn2bl9c6ZmbR1PzQ5gqk23z
zsLHovoqIkaqkAaQbpkaLVaIKuYVBhJR/qs/t6nrKC5mjaeu9prBViqbDKhEd/v+
hZK1VDuY9mn1NHD/9tMCTcwzTcElAwTQ4DwH8lKzdhEHlc8dc04bHToRxmzOn084
kABAdlzqLJJttE7fBOpiMBX7LJ8TnNXEAptRHKAAIbJ37HgUtIHTuGT/YQ4lXdlh
UFyb/ZCfY22czlUIVRoThitbCBUdvt71EU6jlcQc1bl9fjTyzdRIqefmah3oBnh6
H0uYebQo59ZgNJMfAweR42MgwBbajI1iP5QbBg/5u7B4T2Lhts7YhTTJ5wJpc8Fu
q6crP8KNAdj159I/Ij7XsVmPZrTHlK84yMducYbNuBjEB/M7lB+3v3VuwvtfCCqJ
yfKKRI1LGl+u6aaT7f7YabO6vC2Zx4VD812L4+9U/ig=
`protect END_PROTECTED
