`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JxMIkhD78Kv9mDcX6iqkj2V8F/l7WknoktMCfmLftc82otiG7IpWUFIzwqbNC64N
aIjorzlEZeL40nXGIz6GGRXZBDoZ4zqtuA859kgV3UixS9Ddjgbcjv13ggMBTjJ9
ipYt2/+PRaI17nWPQEZoOX2SXvyoVrMYj/ojzZo75Jr9cIS+DZwe3LO7ggx0aRUU
71mAkl34rxO2xkKO3BIOP/hjShYV1/d1vzL1pn7RWFr+LioSz4W35EtMVjfSOTtp
luhFJhXRMVHmkmHuqP1d7UXG6mq7+nuYRFa+Re0aU6NwP1NrrVFJ9WOik1rrtcux
n/J8q+GK5ZCZdPsbPGJ0/fkNHzBKcbL9lFfKhQQy8E0CNvDkBB15s6Bjpzpn7KQj
QDTB3d5rWrOwfbVEtxPVgu3uKtmWOeQAStAkZsbVq3yZTCCsqu7DtZVcasuHhOPY
vhrQ2zK7m2rM8xyaxqdML/jdSohFaDtsVczMqXuR4dT1cVLWfJX0mIrziUq4z1Zy
boEDm4m/CDct4Z9YC63hBhs6gfRtVOYU+Njp48VFVQcwV36vZWhPrnUC4JmMp7JD
H7Rsff4GJ+JbcoLmWQrKINftbFDkbQgcc9gD9Bkz2nFRPu3IjU7OK9N3t2fxiqc0
dbrVzK55/uDXZOqMkDWYxMzXGrnOQEBP/Cp7U6pKJCaz1XUGLkWyc6mKeOncQEYC
FmJrmCfS64dJXOLCun2W/JTg6XvP0rnLYcgHUT754f3OztrKp38jQAE/2CQfHA8P
Y0S+Q6pG/UmqoMXweFXXHAtJ7leIwX2lScsy7/7vZoLOTTPiiXeKiEqYRHVtsi+x
6adOT0178nWfTAG2ZK6nKDZA4pJ7OrMVuoLxPkNreFIsMmsT7DJQKSwJawDAgis9
uuliDa5R3Xh8OTQI99OnIoSDfjxRes3c8vk7IBQoCLg=
`protect END_PROTECTED
