`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ByhE+92rfePe4VmD8LSwQp68ntSQJMG9lHGXM6H3kG1hTgijLMG6AzF7+ogOnkkH
gxKnRE/7UIFd5uts9OdF3rOoM69f2Si7WJE8mZ8KIpMLDIof+6Bfz+aUdeaLlvcg
Fw6yXIWyHEGdcefflBfchTUJfbWNGyK/CqzyqHpPcGoZ6+NissmGFjkRKtUmTLIu
F9k+/X3lUOq/4g59sGke9IXkZMnZR0iVv+60zqaht2HqyDeefYz9vGUvdxceCGmI
rXBGOV3eaRDNUOgfFprUbYyApE0pFvK96GEBqd6ycYV4KFhYzOoXDuZZYPqaA9W4
c3m0/2Q3QQSz8QlfkyHx/azKY2qluhiOvVuNCtwqI9CGPFNJ9r5Ft/j5Q106XbHm
/KNpS32KBO1Pd3OVXUoxYGMO0c4iZPCsRDcLf5hG3jF7PDtf6G7HjhdvNGvXCZgy
YyzLxwdlL9fCvOcNN0J6WMbuvze8xKjMzLmfqMsa/AfkCez5RFCZr7sQvAAsBvcT
EXy39SAcBNvWNAReKrFE1fCN7r+n3AUTMA+SOWBLq3+OkS2GvVPJsP5f6Zct2OnL
me58jB8vyM91ov1KbYv9FsG643bSvBCqVJzMVJIDW5hIYCDGQ9H80pP9TzNjbGqz
GffRoFWQ5ZGujOvAWqx9JLpNZ6zvr5dfiojVNNUavT10iPPHbhotqszE6jg50wnx
eeHxeWVWVCv1UqrmqRensFhOpjqmv4e5I10PUDCaihxFbyLbOFrHLZNBzS/M/E/3
PbIisbMj+Bopov3FMvvSNpzuhHSs8dr1p7Kw9k7GjBdQkfQRZHuD+BbyKdQKogg/
oLrg/zRioaIi5SAq7fUtrhL8KJIcL4up8KwTFNNI6V71xzAD8GbHiGrrW7q5jKwD
yMb8cbdOMGaTpFPEsCtv764safvaFjcPJ+p3NytqWNdt+kkon6hUizaROo9kG4vz
jQrXchEDfJcsBIoQ59ChQc0moqxHdZi9axNEvISVywwBKxDJ7d2Xr1MRvE/IWJrx
w4lEZNSjH6et1UcdeEf3xzInz9DIkzrLCUBpBn3RpeN27neW8axepwPwaHHxSQEM
D9NypAiG0OB5rXUp6dCIIAlIVIDc+wm4u8NG9FXKQBPh9DQjsqPe5Q61WKiZewKA
lGKIP35k/hIa/MSZlaVbjanyYAoBBOD7EjRxjT2iHMCTqLVOJUoIvfU3KQxfF2z7
St36hfv0AbD68aMREBjsiXJT55luwCF5Tu1WMvoXaGw=
`protect END_PROTECTED
