`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2PL3gdRfeQN8+GAGSPhyGy6tMidOWptCSIfg9YCBxPeA9cMMw2y4WyHDyFLYm9if
3+51byCAaSd931U46de5faG906KcGJHsy6+D3oqvo3zCKtW/KJ2wj/NNIVQuFtsv
Q7MgcPgM4X5crhZvfJ0woN0u1AZujnZ/jfN95WMe51lTmsPl+N8TePVcWfBrpMhH
A7PdqU60XQSk4Bb0wI/47AKSTR/ddRg31fqHBOFs6a9jxw3amqS20EGy1wepCbLx
OieRyr7t2xNGu2QjlNll7niJi/TgmlRmTm4DD+1Y0fhjnCfk8Nt/WTeUhQ25TGxP
fwA3xXiIKFgNGuKaVAWTY8nB/HgyPbsM5Lcyq5VGftLtrTr7cU+Zp6HjHSGei4zK
Kno3yJX9PQ435Ql0om7DukqWJoMaDI6Ii8i/mitweO50LHtHS/QoA+yL7px05/SW
1P3A5ZVSsK+KW6OS+OBaKrZOIbRp8R/iMkd48UOc5BEQ0gPiClQuJE6Xy4osmtyn
40HRukLslyKJa1imNz1EUsDw5xpTNFvabo6siZ+mLnFf4+XK+CJSYaHdrvUL2YQY
y9TaKfOsy7B/0V0siMc7bDAPpITdMqKp823z8tpZakhrnBgoyXcC8cJDtLTiVUn9
MxjeoZlRZ3Rhiy7ElHwBPugA5lQeYv0XWqek2al+2H/BhkkgvtX/3QVM6rFnieVr
hTqJiIwNAVlXQZGs2sdTpHiuDRVg8Ai5Nk/K5lnpPRBsQ1/LMI8Wf3mcHFMJzh1q
vKqBRHJXazuV0DgQaliQ2F9LCCivL7My2L3krk62VdTl1aYJxB4Yist6q2iknGAN
ntSssBSLjz+zidzSdGvR8uyG6VBgXbDWdabOsAPylwBl6FRMa7vhQjrWdKzNxAvR
jo/K1MlVIt0/Nb7zkolF99HaCHISuSLELIPV708TuVRnL+zborpXxo5hoVP3p86U
mww0mfyUFQSPc/md/RJfkFsATSsJ1q1hS/hB84CYF8+qhEKMjD+Qeabcp1zpSb+g
WPobbs1DhckSxJBKTgbBRrKIrjqLX8RMOaPA4aFIgc3ge4zsimAwLRQoRGKnKXX0
T3zNa5ojDAS4oKzfmVYc4JV4E4vNu7ZJD7/3MEy36Kvfx3LK4UJkeZpoJVJmGaeq
2/VCs0zAyCFJcLR/g0rUH99h/T1XZlNycvJj+SeOG93hzwqSGkv0IuNalHEIakR+
Ja0UW9ZGPUJZOt7+YH1Z5xtrIrn7YaoFraVsgcsev8MYN+Msakh/zKUGVmL2hUMH
M9i/Ij64v4vKjfD+OFYRqxy/Tk6mL74OPQIxhzAd1w4xNayIr3R16XEf4qVMVXeM
sVwtDg5D2uUPEI6vDRP2uXqaPl1RoRXSTQ/CkB8fVJLladr0txSkImN/96QelUQo
oWcfx0YjiT82IP6ji1B0ErHwcGdVOSYz1MHKF+vvkS+N7lk7IItlcO7jkZY1FiWz
GAK9+yPqMcItom/hmgD4ZZKVZSy2D197gMsCEVRzGTfRpBIzz7YnZUuFGEPs3O98
hccqZqoizLfSLlQ5kn5dvczLZx9NpSQ7Ni5mAhHBPa06aoUXEP3GWmS2hZr1qopH
a8o7HsavmyKen8DG5lmM7tuQ/u6lwRg/ivmyLDpPk42dqPgnSqVDTggnSBvMpyXS
NNT4KrPX1gyqlO1jYMDlJ3wWWaSlndbmFQo+RpYof7nBVoraZhh0uMwhHU93ow1j
YadefWj4XP4bDhXedZoXcvec2g3KSbWIiQw6NH1q8Qyuv9Ny54n7CXnfQUQinUac
`protect END_PROTECTED
