`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5IpnJ/8/r5HDkrgUjoQnEYjZw/INrWCkgjE716lLkbX8Fe0+KbMltMdGoH8tLdC1
cJxS30ZoUWCVq80JqkOslVLSvZgf7Yyqh5s0Q0iIm+hO7kKucNJHUQDb2/oKqy3W
o5b8dWKySLoExAcuh6vMYx75DTuFJ027MhMuRtqyP9pPVrfxH2VS7RceR7WMDd10
py+2kTpbZFOGnFo68y7wbQc4U1qYU9IVfBPpBGsQpdCMGAwZ/a9qJTI3w/CN1MX+
YJ2j9OnJPUBLOx0LbSdyYo7styNYt7rhI+yYhAhfJ9Tz23pVkbYd63F34yFIdUii
wzIp1TmmVfzy6nAI9SbaBZiMR7/fGj3vPsX2d2Z2DN/j4VRFZ3DBl/3+Ykip1zV+
vuWDaNeAJ02Ai1ShxzyU2JjpH8rC7KtwQL0i/gX60Ahjyg73EiLc0/Tqct4bpkDm
ZV4X1Dbwj3EysTjdfGhRclqfSC3mBfLocyJz7f63kkxWjyaHYcf2bjvCqTnkv9Y2
plRMONoDs+EbJrLM+JQnclDuALaM8qd0NlwXPzvZpoLHAkh4GakIyQzpu4hobZ7S
GjKiMxyhS0Lxp4uvGYl6m5hRHOOo0TfNiwV92spZhJdGzdMKSBMKwGIl2Fo4U31T
q3rXy0bAnrJHwI3utWeyuIq0oUeU1qQ1tprIfyGKmaXy+V9F6nsY2UgnSBAhIDpU
B5JvdmsMCC3+x8Pf+bmI7w==
`protect END_PROTECTED
