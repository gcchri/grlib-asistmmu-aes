`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j6bNQuXphmM2oTqSVYrUyTXGixrNN5upslFziOsAQo3kvfrnORsphc0lfBS/nNYA
4HCf9ahSLFEMRQvVf+QebsAGB7PKDzNnNW1HVttwH418vWcY8iWEZhLP0X+A8smy
rwB0ttrWf4hCpEocesI5py6AObOVzNN+Ex8eNz6loS5EWyzXm4gaJpJ1puOW/Q/G
yKvi2oIwy0KT2j1foO3DWEzezGLjOooG096T0kp+6yiratgIWCO6YyX/Tec3fEt0
rogMNlbbKQSDCvTNBz42J51hBmQ1UCeF/CU+ynrKiqfjBYV7HFNmc0w35UXHa0YP
PWwBoh96dwb9wY6ctrrqIBFJhsijIbEGkthU3hWu8uwxYcF1z2R218lGEibNfK58
wzTh2cD2j6J8wD+OMGTjgu6VsPBRnAYbO7ivn1278h+LMDUQOpIKnQFrszCUPSSi
cUB3ZKlGb8YJeqmH2Vn60WNB2YSOZCH/HsXl7fU3S6clOy2QO3xTEc6umEV6HDRA
ktvHXARYZZn43FIXIGcx+dJOBQ0wjBEy8s3rORhI8ZG/fHtpnvIBuVYkXO5zwcVJ
j1bSPHDQdP7Ok2+Q9FnI9gkjPc81Zvc2Fy6Od7ndSAmAHwmKgnH60lwcOFUorOl4
cCC2e18r3ixeJmA5128ks2vBJwyZ7/aIprWe+WiS+k028hGrJ/c9KzOvzeB1FQyK
nmB5sqO6p0rZ6YW0ccn6lOGC0HKBD+hPoKr7WXFrK0nzQfFvIUQ4SBKxm+ndpgB9
yzAA9ko3Fm1boDCGdblR8A==
`protect END_PROTECTED
