`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/VAy3Um+XqLPNzj7H4+D+/Pnb1VgB6xNbr7iLo1a+0XhK2fA1zkgku/UHQ7osjx
YolcoLsDUCjUAjzLMbnmpl9CmWHuEbKvJazI2lmXgLlQb7DtzwjBeO3ngwCcnWPE
KWAKGSPxqilXcizSNHo+4889DLEXtHYpm8ZxxZ5XSj1sOrXaU9lNTat8S9PK00G0
Wd5OdSDyliRAWE55snW+PjJtvbSNZ+S+3n53qhdMySX+IUbVX8WJm43xZYbYqIT5
8b/rzxgfObniHxQyt4RAde9bA3A7nma/K6NNagqhlIF3rwI8NnLqHuxCMADvqW+L
/9/Zx+rQAMbiSMyK4S/2rg==
`protect END_PROTECTED
