`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ceihu++MXUalMqErTfAYrFiA4mhWShMfiPhssT7eAUb79IGKox3AHHI/ZL0y6Nxj
QcSWGYALzW3lZfne8PGFRpPdh65vt/bwMIvAzK3/+UoYEi+uOlvCLxUAu20Guacn
UsNdkGhZH3DCDShF/XZYkI+YO+SMpYLEW3V84U8bX+2KVxE+e7qQVKwLt8PgyrxW
Rng1skMX7M7ypO6luMiuA/X2NDq1disMkdoyIayQXqLQ38ZHUhN6z+bQQaoAa6Yv
xBIkCiQo/qbi9G/HgtADAahP34wR+PAA1z7J3Y6dLFeSDuERZUz7AvtjtDbXzFAs
S3LkOc9KxPfT1ktXQ2APtFHynP4fdaEjBUQO3jSik1QPEskr1t/ZOQm6NAEs4PKQ
sBYU9QwYFQqec3GF+ALgiF4sqTg9aX0s7pRt4oY+rTQ6nR9mPhDctru4Katf1rte
hGTqEDtzY/uXJBLTauFxNMsXmsuNIY5TqcoFRv0Sxc/PQYx/NHqShfWxUmE9B1Fy
pJ+h4Ry1Wzp16SrKbCxphE1RZnwu+qtnHTPQ14kvDMGEJAM8wITe9C2KOWer/WFp
pJMDBt+hEyyKmfdSvKRliW7OFyvxY88F33QH9pdo3BDfyeSwvo2oOVtj6PVBy4vH
CUu9GzIpEjhUb30+UVI3Ld1Oiy+haxb8RgtgJl38GP4lW1PWcau6NW/gkQLVWIL7
tynw6AwnbLRSGvtHHn7kbzxdBl7GxEphtPai0t/cflS7p+R9/Lvko1IBHBBkoTZ6
5RjGgFROV24VTSLUPKoNTbDZMBewQC89oGSojdS4krXdTcV1fyhnuMpFO6xAEc2k
uxvgbZ7i9JOQBkQdmXnYdyuJPNfCTLWlHiMRU7kYCFhV2zWkdFQb1tQ/2a3MNSKu
mJ3dMrCTp8sVOgMO8L6q5QhmkM/QoE0sCyDeRUKfC/dm7Phk4ZLvJgGLHK6itI3u
b6O068R8qvhSd8Y9Rd3pAQ4Y0driPEEVa/QE9eQeq7JCR/Bk11mbXDwRunKildGr
PlXFuLrswj/mvd4e/ReNhq/uocVNC9VkGx6NH51inY+WWc824UjPxVZKPJ6kTIXH
kdH4rNZ9BmcLFdppx3Tj2YoECeyj62+kuYMWi1oUaMnIw4ZBWyRNyvgmPhwadWMQ
wjiFTT2XaXZ0nviMFAgLXDHTbgvvFT4Cl2M5NHJEWvBTd14VIQwPAbecrxyhkLvx
ylMEd6n2EOz18PzPxA2kNZnrVZYzOHChD/3U/cIpoAWJa5CHoQqgQ9RA/2Thyt19
5Nc78iItFt7QHIOvJWwF7qt6haPwpnj6nTxFeH7SObLKWmV6pl7bbCQwzq6Z9XYf
Ueb05otI2pV7+T2Hx4EYVYvkNOcyPqa0RSjMcQLn63cHrHw/Fez3dBEyQbwI83Ez
JTSgkkjPXjduQrxid0A/Vo/k1jl867wBGyI7dVr5G2lm6w7YMfqsH37PZ60oHSlK
clBleVMAuDUEZLMNnfxYWVfWgz4allnvFEbG07PLcnJ0hwWDwG6t9EvtYwwRcokZ
CwbNXkIQP3+8hOkXoEA+plbc5V/MingNKRJukXZnRirb9tsb24qWvQlQ4CJXFLgY
bW6yzZ2nmJcLp2tNFz8GdsniEb2tZlPpd0YuY+q4cE7vEorSQit3UuWIESTKRRQW
WUeoJCFwz0pRGgxIeAYx/cznK/FtP1nfobB9J9NDu24Fn5heMWdMilHhOzoRpZ+M
t9UCOuSBAmimhdi2wNPD0YuQ/9evXVFBgxBYX7ODqo8aA3FKIhVFUS7vE49X30yl
wnFDmyTNnPVH5MmjJpgHw27VkCCG1d00CxJJ1qIyNNeDa3SzgDqhoYGcAC1IPoHo
8rg/r6Pf/vIAJeQORAHCMoSS5UGig+O/vsRKRqivSo+pp40i9g2WDYlQJqcH/fK9
uiDHjYW96bw6QefElZHiS+T+PvP2QXBwpvsWwO93kJApKdbS5h0OvS9445VkAFmr
XkNyhPtMD+v32aA54rSLiWrTPhlcwel+EJgrbitzciNbfBBX0lBsT6ap4YNZIoX+
XlTDQA5c1livb+2yuViiavS1Yu9C/Ixb3ddvkX3sgTzEUdCuI4b1RkXJsk2Cp3eD
arVx2McCGETEFTXLgptbFimD9qEnjj73o4cBni80p03gAK9knSg1U7bbbmtk9lxT
dYE4OnZrsyWOT79JFQ2+6yL7yhHzaTl1c4asocvt7aPodn3hmLqAff3nw8XcDtEG
Tnhf9UZRAtCe5qBrRykr3Yr9b2aHSHD/jI00Ep3qrRG70EaaX8pMGyAllLUZVY2w
41+uiSt32s+6hS8jcPWmtqIboNwuvC5859wHGpkgxNv2nmAmonX6T2t6A1XFHm0A
Qj2DhLn5J6umqa4nuOIz36NAByO0g519SoueDbioS95HgIPPL+02fLb/sCChuY4d
GWCYbGCvgcHamHTgh+4wbl91u6zZW7a/OpdBMA+qj69ioRA63L24EKJi5Tx1y0tL
+gDRj0pkG5DpHIpbDVd0UcUryZhaYY0LIfPcLXT3gEGZbxjDObGzsodTWueOnC+j
n9YrYs6x2OacCY2AjaTviFU/uRKbaD29Tb4PzxU7daV6zsbz0PEu5lBvhBoVHc24
Nl4ADxkfic9/3f7K6clX6qhcRw97HXD+1XUAVxZdhGwX5ZtCER7qnhHLUuaFcPJq
Zh+/gSUDn65VVSw5ahtAYdkYvQec4RCtAqKPcijtoAelOX42ttTS6QKNoY3Lmj/U
O9vvXpbeYB5LdvL+loyjr1av0OS5fzBBGbLquBjKEjD90fE58p8v8unM0R54Cbxg
8ZhoCRbdRnIpJedxrMGS2UNXAWRX4Ml4mM7crHekgP0k1/fwu28Yu14CHRibTgBw
Buo4AkrIpzerhaIdOhLM2uxGeqq+5KWrizK0M+Lyl4oECrC+ul3OLSBcQtS2b+2P
Qg8kXexUZHZSOw37awiES/r1T2pAhz/XJM8qkrJw5/j0zn7uXvPIsyX+H9+mBR4I
22I9U6AbS3LItr50+Vfni7chjxbYWtOH3ixeeP+n88mw1ZOeVq8ehLrRSBOZvM+x
oh2ETEipkbXSC+3NL42WogKJJGozqlorI8sWWZMeZGdnpdBSrjAnHMwHD57Si21/
32aUVlwdyMwB6ACdtaAIfQd7EqcMCIlbkkFsDxoFeWVMjNIJf/xTaWKWi+MTMjgb
2SUawnFak29jkid4C5P5rJMXvg4v7KBR8d/d46So2ODQzzQP0DTjaSWgqfDxwJrV
pE7jiwpKlfyMN5ZJ9xPvhDvpVRlG9Wbm1Re3G9Lc+MDS7E1xgNd2sgG5GYiOaxCC
QyN5Y1aAb+T1AuuW8yFZ3z3KUD+h/MYRM0WEgQA28Z4l5Wh7ZgITt4jj+2M7v3ZA
VOVoiWK3rbe1oyeplaiulblbIad4JsuumB/QF/8tGTUcTggjq2rATg9cDKZ2/1yR
E1F12zhcZQpUIjqYbYaqMGQ4GfLlt6dzY2IZXTjkPMuaLvF73iwhseesa+jMAGO0
RFAqdZIDV+HL7kVs8Bn+WOeJdcdF3rqEzRwY/O8MNDkUrJx5fwPYsbzd3iblUX5F
vGdE32eer/DzZ4PXiX1yXNxY1I5JC1/jF5WPljb3kxhHD+VTl9iJpv5aeRB+yzMI
epXzMca35WyMFQH7iMVVCIIk+d1kEr+VypP1wnSbSo0Yne6rJ2+DSq0cI0Tlo8fe
edK1iw1tnmRoNqypRfD5nBYzLtcKD888gUJHpjFWVJI12NjNqeSa+Iaz6bM9gksV
Fs0R+xc4XlaNddy5Jh76qEZTtVNSktILJuddn9EvCuT7wONnD8w8E6nMs/0NrvhT
p0SuDOgmoLKx9qxlUPn1yufmx9gzCUYMWc8CGdRXnqKPBbocAzIxvL39LFL6+bAh
mKclpKDEDfdWcpW7p/ckwedQD3bp0e5IXFe22vU/XuE183XH47xqUfm/LVRkRcjI
kW8HEFlvrFWcJW/yZpqfG4akrDPivyuiUOu+rnrYLFahmkx/cQ2NXUw94wbL+fFk
G63/E22qZOXIr7RVQr6NmXQOMOeheg0C2Smuf/GOgujBZA0xyKYi6EAtXTP6sJb7
kUrUDSicZtkjjkoMLrmKXr+FBEnKiVS4KgedBvB8TJWWbX9XoVaNeaR1W5tIr//P
RhlcMo2Z1zgv39bcKuHZLtYZ/ZXmUe8FQ9CwPFPeSIYNpuKENAnGy5E49YCKObwu
gUVdMNS0Ui5hUVPZUg2aUk+4scW9eht8056puTe/PY94kW1xob5W3tKHtGGbFuW4
7/Nf52vEhgft3XTRhbztWwFWxbHfDqkn3+LFT98vHRy9zTcQanxNZfAmFOWCDz8z
Ud3dINjHrv+FsdEukHQeObkpE92sVbRHBr5TEF510rbdxQ2ygQEojAQl0cV4nI+u
t++VqpRej2ts40YmQfXFwAt4gCCpVmb2dmLCI+PbTklgyedDpLThDt1HNOsiI6kD
hJOWWPZSFXk+N74is6N4if9EuhDzEsyasFFUVUDvkd+zfbwyC/WDFN3la+Kw9o74
Wi0MhqzraAjROImYeXaD25eGSuiWNHaM6ks4y0MkS6jpRlZo/bqbvu8LDPiGEMnV
GQrRYvRwcTPx8EvIoHtmdO+b5yC8AabYHsqkROnRuK5BGExZjfhsoieDXSD4eY41
uSyKz3DuVFbW8y4yXzEUQlUhoP77odnD1mUUpLRHkA5/LQBiOkKxBibM/Z3LXt5k
76+/Or41JxDcA+DPGhahB6Epbu07KvbYwRrRq95AQoSm8WSduFL9XuTYyDO3HlV9
BjvYgF9sTxfoXhfE/0Yfy+4+jiSkdmwD+uQ9S6UKZ7TA2dpeEh8dSLKxyaW6PbaN
MCRHqJJcj9yw7zvJhhK2D0c400ed3hqbjHXMm2pg1msMN+fFNlpR/RZmDPIrJwry
XAe7k2aJYbFqesttdsLTHEJnKPqhvGOxZ4yGKPYThD2K4SNGbk/Hv5Rp1QJ8Mt6v
driBefaNkFN9jmpWcy/DoCgZscfKAfPWXl9+7hzH3Fddg2mUKc6K7bJaGiPbRPZM
DyfsdPRLuNl1gtrkZGlQvudmeFuNJfb41/luPDqrAJebhdXjDMRg0RRUjrn9sK+E
/5b9wylLtkoqgd1ivib6kGWV7OJBX8jzBWU0oeyQLntTUjJQ9I0dfXXpf30t5Kh2
B8YcU6p9h6waNLacBrN8Vjja6LEQgyacu3eMEeUxqpd0mBwSLUGWVAICsXKpYL0J
k/uFz3LOAnBM0k3sj2qNZtYT4tRy1d7RTRR0ABC4CnIq23PgF4/66zTNfdgPaDgO
ic121u6pFpQ9+kFHIPtrnk3BMPtctrUQN0CteK+0w1Df+1wbTDJW0wfqtDyjwgeq
Zm7+QnAeGdutG5iRzlOQSXWbe7QlVIjaoSK+Ydxp0WOpL4vRkPh/rybiNDZr8/vq
TlmMYT0PQiB5QpVE/6uAf0yM+tlduOO3gvrC3QfhoMksCeMOdH67DtcUFk5nij7c
a3dUxl6WVeKQkDZjvSV9QUqmEN9+0GiLJILe1X0Fek/glWu9SSDdZRFrOTubvezC
Q1qaE/xoYlwNF+wfGQPRvbK/x6ziI65Z5bd7buaMuDA=
`protect END_PROTECTED
