`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QnnBb3GpdDB1FhfcZos3uFt+GCAtJeFW7aC0V2bsgK8d2ZD5d7wxF754VvkGsATk
seHSX2CwAdYIEceNlfDjHXdxS7vvKInHp3XBRNVUjImMpzKnPU4CVvRBYoV81ykm
4/d8Qr1Y5PgqmW4nRO7gjyp8+RcwdMf7Ahu36T2uR+Tyj4BrhFo1BsyLVOQlSayA
nHCSc9eUQEyHsTKje46NL6BYrlaZbkFvKiUb1TofI+dg4xa1b+mZwwg/OD4zmFQM
nn6+jgKs8i20fD9Z6CzceyKR18I2ZqCeEWHF+8R8oDE=
`protect END_PROTECTED
