`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0BW7ttqVf4pcR4+XdiTIGbIvbQk8yIATxaZg4unMBHkAR2CWBcxL0o3ALl/YTrHT
DQyCicZlJuSAUQ/QB0uyTRatzkrmlbkVUP55Gr84Q6xUwNiCI/9qeEBIZnWP+opV
EWK31en5FpSs7mww7DU4/4RT5IkpkPJhkZE8h4fQPcQsWfGehSz4WCsZ2uqnlX+I
9wLdSxugE3ATupN1d9bMUGpX0huVUkIsLhTaokkl1xHvy6cTxDmu2ko64qAh4WCH
hqD1Ch63Gf9Wcx72sqKZFMdqIEN2DTKbZcEGQ/6bI/XdPGWNkXMekUrnAXb5AHFB
1f05Mx3IxXSRiQRCeHBKT2f3TgI5FWpGmOmg6oGZN6dB7KYWaWSH6+a7h3/qDV1A
Epd001cxPmFzz50KywifS9Y0FdI9Es5yLdbe2zcRSBZexuPX6wl5OjwuxPy6+iEz
P9iANMirbF3uiyKp9b664acIZVQx7KZQOuftZW80OKpO3/p5jZTRhVvd6CnKARo9
kNVVnLiOouN8vtfnN4Er2Ap+n1PfsYxLPMN+if6p7aKB9BOB5jwmH3+lweSOia9y
W2C7VtVC3zjeYyWQgTbom+2Dw3SRJiTAu8I/opBzRsM=
`protect END_PROTECTED
