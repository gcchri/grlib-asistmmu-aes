`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1s7oZ4A/+67FLkgjs55o++x5YNjQCBegTWhLd8xcnr6SLjM7dEWP33RedylXKhoz
MAgPksQ2YKgWnHqaQb9x0jnX7t8aEoo7JIA1/Dx+hPvXAceOIe3fHds/TlWxhVCp
TgvsGc8qlXiMtCrsqZfK+I15osgBZ1LCgQZbVoMl7ndwozEA/SxaIw9o11ZGnWhO
VsOdKGzduQAog9s94nOkYAkqETJZR6bGcYQjKet34XN69hAqOsOzrj8S8Tsh6rtn
ta2cwP4P546hzp8zq69kRr+8vNZGfiIwBKLMjjHg93lrHllEVtcrmObY/b1PnCgO
nuhX4p1SaeqEHsIRlFv2jnGTudOY4gkLglptPyi4d14b9SPA7WhR0F2VtMUl9l28
D6rbHEF7zcD7VXV57fgzDAf8xTROIMuZH9NqzlU7Yz7SH6mJi5KVip5c7bEOwnzR
Iv8jQIZal5tzbha6IM1/yg==
`protect END_PROTECTED
