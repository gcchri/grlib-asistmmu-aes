`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
01lBBiDRgLSOsKzqapCNID63GBiZ13GROcG9ha051x+MC52I4s+WoHBeNNopnaIb
91wQscdKbAA+hzBamIZ4tQ49uo/xYs9bWUB8wTXxFHidLnQgrIbAbI+MkAHg9MM4
GEIm9L5VaaytfflsdrORcZnizWovW1+bqmw8R1bTZBDiQ1ckyKNggmvbxnZKIc2y
OSvjcZ0k9tVGc8DW4qwAottmCgFN/MbyJ4mnyG+DO4w6tvy9TLXfRNmbeqwXI2UA
i1diZkJtbDiaOheNxlKCn4FO/IoPew2aaIoKZx/8+uYhbomkzfFkrrEJCV4NvcWy
xUFW4yYkSQ3WaTQy+4l6hQ1wghwi48yyXb4v4z3gds2DPv9jJ7T8LAVbU10vFXce
TOGFwBNnItwIPp8sigLVqAfjv0jc0fq+a7rLUKb7so58iJ+RF4mvlZi0BejpQilv
bK1gomdg5zWFaW8rtwu0/A==
`protect END_PROTECTED
