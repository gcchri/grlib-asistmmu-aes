`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OQcizVRg31sOJj1TlY3TXk3XIzlZBtYBaHJd35zDORsR5b6TpOF1u9S7xYyRIIoA
59y7O1Jzu0pij76IEbUly9sjQ4jl3ic6YsUnkE7D3XRRXaqiFzPUnvzUltTolXRM
n7kIX6oXpfrH7VV1VODRKuCfru6iSSUC1HmNRopF2bskr30ZPgrbnLzxibQL+VNG
ESx5eukWOZABuWZsnnraTMeNhxtXh4V353KF4fJyYKdpJUxhyW2sP90ZQLk9ZU+I
1Q67J8j60I1K0ixVu64OuJmDACorYaPah29DslwUIFNAshxX5HGXciTjMdDkhySN
eMoGkUPWQML/32+AP4GzH6mSKe78yElRhyurrDWlPTAj+Xro1JIZPTQEhF3oaIxF
k7i+E2EgyTH2bAuYL9MTwJUD5oFOjTnl3j8pR9tocfJVmjtSNf0ZPPRM1OPe5QMY
Q0sY5WmshgpgjIIIurI8Hm9Bvgf5B2J1YcBE5IarpE9a01j9t71FKQfstKeUYy30
Ga4NWCPdI4E0Mv2jhQ1hvkQUuOMepcusjhe2QAmRLwBMwcUCUTKzctxh0kjEq6rz
N45OF0R72Y3r90HDcJmsERwtWs3N6u0Zq/os4Ei2jZQ=
`protect END_PROTECTED
