`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tFas86bh2RbHmWReA+MJBBWouEbqdmRYfdPC/tTJRS+lpcDsBvEFVkiPvz4OzlG9
trOdzkZ1DHCB417yQ8S7/1j9Vab7BlzOtjS1AKlu936Aj41Jg5ITDEVqfLrAL54h
MB5l+VILVYEr52y6DURkhBL8JxiYC36fXfze4M5rifiem3KD2n1EATEBsQUFAnzl
Yvy1SONsc2Q+SUBurEJHdr1WspOHiucWMQ2+IU9eysyl2PHqb+4SbUSb7ttZ4/RP
6/A1Y1XfB8eI+0JtoFa8QYxJy80QNWO5Z4rAI6c5SibdJwC2gCJ/JCn9NpXc75/h
uawVZqRJ+c8h43Xiza7dPLSBqAkc/DIlRURMJgB3NvIRpOfHoOqQz/yhG/JstDU0
+OzIxZwHNgVyjsiX3m4dIneCx5dCWTytG8RMrp08DT2PvWil7Nfju4sMW09eHiDr
vJYkG/yX98zVIAQ3VDKXYg==
`protect END_PROTECTED
