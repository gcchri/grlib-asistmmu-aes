`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQltgO5yuvB1PX2vfWWckUMatakrtnUV/4ofupMoXvBeyXmzlMCXWmEg2B+KOBwS
ES/1u2Gh2TZBn89onWuVJlMXsQRijThOZqpWpjOyxrmCnBw3qSBaDhMyluWJhMaJ
XkLgOzUua9dhdHVBNLrgTfbDcDmfbW6HpA/R1XPZiRB45N6fMcvTQZB5iE2TuFmg
yHgXZCZ/rF4Aj2aqvl9IJsy+yPTm/VhBwKftA0oX6ZVXbjThNez8wgW4k2QZn8al
/+3zKBWJxo4D3CXfplV3CGahubQP8X1p/WfYUIyC1fEjE0RxLuNolm/lj7w4a1rt
YbKbL1rvfidje4wFh6LKb1OqLQCvLOiXUCpFAvTXi/uOOc8L+v98Ay7venbw0ii7
YtieMGcU1/tMTlq0+lg/+NUrJY4cFRVuPQCPvcwm+4P39wZE6YRu5eiT9TqKY4o2
ZNqx76Z49mQ+gUKdhxZprdhm6HVwbyTIi5ZtMbxpdNR46BJbn+3qO5btWLIxF/+W
GVkeXx16n+ltpwBeuhhRuA==
`protect END_PROTECTED
