`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlsKNOwNmXzMuC3BiwpOFJ3bii5EhFNXFEY7pwitCPmuT1MWrqkCs6IDh9YT6Rfg
XYaLx3g3MTHg6hf7hiVcsaoVlfMX/xeJvNi/GfW6HNg/zZKePbITJm6kJ5b7gs28
JJDC+jy9EnPfE0LF1xdUI6kJ9BtgTEXsKqEIc1YXW7DzFbX4QOBVGzlAgtyOQf6y
Veo4XtJTwePBuLN+OcS22BjIv91xAXP+Lai2OQ0e0ARH4Tr+czHzrwsfHDKn4X7/
8j35RjA8iMdAqvvytyj/3w==
`protect END_PROTECTED
