`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KH9CO34IJ4bo4J/Jrb44/6JPLNIYHTIGcP8oLsPaIOkwM/FU5HuwsvIHtBZHS+QQ
vMKiwvovyo570nIWSc31yIoLZoHsWtevPliHkVDdZ8KUW43vwU/OAwm4i2WV7xXP
brrw8xgTYCyYH4wOCPYzKU2Q6HUA/ZE6upwYYSqlw0DU7vzdnYl5u6jCnIrhI5X+
rTRV0Pki9w6vtU8vVEf6f40mXLhHsi2H9V1Sh0dYBlOCO46zq1On3kH02zCUeF4o
lKbCp/wMXXK9UBt2kFx7YTc4dDQ6Dbzv/TjxMtNQLiolf9MafB6J/J9GMbVOqctn
NX/aDfXf8WNggi5RHgPpJeLPUa8KdF68ch7vGNGY4hSJ5fy2zd+AH7qKrQ8zNrmd
dnxWkKR1hzF0KMsv3RIJUpyoa0DPn+SyMtlUPFQ9sZYWFvdwoFoPC/aSAV5pY7hZ
zwJHt+UT8PB00a62RSjVE5HESzu6ezHienoZmLpRZN0QDO59xvSns6Sli40NX06R
SGPrkPHhKYA1fngQSN1KkyDztGWhAerZfpzJ/zsSIthfelIjdu80xu68mMGG0bob
0PxE4NKDxx/WUjj1r+lBIrziW716mFK0hpWSdY6HlO4=
`protect END_PROTECTED
