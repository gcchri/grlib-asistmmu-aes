`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
slSRuCcHpfFan8Jms79JIxkR832UFou1tLse+uYGoqQYU6zCwvp6YRZViioah40v
U8tWBWxBpQYv5UFH1PunozZPxfCYpbF6amenjaq+jZZ5vc710192mKI52GXEvOHu
xzC4Uye/v9NWRQcjVLBct9M8q7pigVnws5nXw3Uvg9YvX7n5ckMVIltcUReiVwj6
2Ass+vp4rbViNWhML/16GDMw4ozmFnI1CA6A33rWJKOixh10rV4+QjcvjfhBYkG9
LlhdTCIUJFrgbwyjSFvyhzQGoxrMmW21D2GxBqoNur7pzqcQIW8Psb45AMSOHy2I
cSMk1tHSwmsfJl0L5SNc/N8XA+UTK13FZEakXxuk+xms5b9nRMnAO5ZTK6DvPbWR
t+CjPd7X5xbVxG5iuViAijnE5yxZ+9leMyjNJIfEE/9MlWO3fhIUaFZ1hgjUQ2sG
oCR2QI5wpDSyhGdV8jNIJ8urgtPtktyRa5GCTk5hi9x4GvTKYbeZ80LLy1wmnhxY
Ycwh3xBXyTXohcucfzmWcqmWegvDA6BY0pUD/Twf8k+bFwBeF0mNd3znxtbJ/WTT
+StnFQ0xCmKQj/Q8I83dekhB+M582GCmubjewN6qe6Otzii8qf2pTNwRqujxiykQ
mt9rqjUc2pbtwZrU4yBpnmefDdsBfXQpKcESGN/xe7GnDiaQ1MGy7Hlh4waUrBSJ
0QMLd4qwFQqpn3dikhfEwFuHvFE0KRxN4g+x5BF4Bxs=
`protect END_PROTECTED
