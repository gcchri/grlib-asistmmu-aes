`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fGW6VCHP668koM5WqxU6AoY3EyJ64U+bOAkyX0wdVQl2HYucVMW1tqL+pGR0lhIF
aIyOu4vJFsFFrpholoico5LLyM5b6JZfV3rEtUvA7f+jhkRR8+s8GSHP+jXo6u+c
v7KNKs8Ge9ttYyIKKEYuyUj6YyABiTiTbYdqxaarikrBuNUNmAapGeQ2nT6kJ3uR
PNCRWTMcsMtETggp9iExprU1E5PBMbgaH1iQE+ZZN7DL3crmRMEQk0WCzwZDjVZs
gDI1esOKVls5OD0l3kxIaFgz6tw7Bk9Y5kFSpzYHLSHctLZxJ/NQCF4u0rpUFl0x
`protect END_PROTECTED
