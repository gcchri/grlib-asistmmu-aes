`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KeuEHQwi1ZxpwevAbNgq3AA3WE5mkNkVw/n7mbi1uOmzFXhTIM0CsrqBfGPV3gtQ
MSk6O/9JP+Hc9UF3L7bT2W6lmKb8+Jj+7fUiYgS5pYLvhRpCLfNYk4tihda0rLZZ
tfCSWSRUbqRMY+802RtwUOki/SXKQ54TwJvdvD8Gimn42XM1umyOVHE53rW9n1+A
kPFlZBB2oLH0mHKnMCaBH8jRG/EK2GTnpA9Ti1eXX9uvUx3qylaahtBG+vP2QPwW
tqy+fauLSMDTWI2hCaY5CTUJcVyAu9ya0EDa4N91qVTNDAxKgRYaJbEI7L9RR8l8
DhPK2YaFs5yzbiDNGqiruD2LjYMtQU5crFffUY34ScbbT7f+jqcfNhy94Blc75H2
FhnxvWBr1eB1sk+QAv/h3+6lcPQ0+Up5DZ7fuIwSIdw=
`protect END_PROTECTED
