`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Dw885tSO5xgkLLejBHnNwPl+G9wCdUXZ6PS3CFVFo8t1NOIMoDsDu0qLA/i1jpC
xbEe2nNgp1qlHdT72mpye2QSuR6AocaP0bhzqN06GL+Sdi16e4q7fkmj68+yG2L4
qE4iu8/6dSJXGlPtYNJ4mSat7MpCCNuxhWvSKE1dWzv53VyXDZQbFEpzAPxfbfQY
8Zm5v2Sv4NkMBBgsdfTBO0uyob6K9RqF5tFOEbhPVbLhCRgF8ZMMSHskvORumO0d
S33cLV5JzcyVm7I5AFdt90pm3OSWG/QZt2NSzBfj78VfI2tbC0gy0k1mhUAR0ZJX
NI+g9MfBoZrgrOuBMVDZZ940l6cUW40SiAkHQ+IleZhU+uTL/dtg6z1cjYPrKH7P
ltfa5pPrFDtZ866NqouExA3+nKm16OYB6FGgrIsq49XKGS7SlAjrYBf/dt7mMPfb
qIKDPZwPITpWANB/tlP60mH8dyyRv3iNvXc1DmCj5N5zISO3wBG0sOQGbUJEwCJm
wiQsXRZjdqXmm2qfskqw33NQ6CDqjl6IL1ODskMPVUkqq6m7r6wfbSzT7ze+pi5x
yAxMnnE4BrRFwx17SZF0CEayaUEI3E3nwRecDBuaIMvA2SGDUSwFIJz+4g2RZGrg
L/X0U03AAOWD3cwoMjVnkbKbg7gNwdLw5ckqvdgHF+nvO9tRqruvpZJT2djWA0hl
fu3YD2phGVgeBjLia+r0HuFS+MlHFXS6QzWj3fmVWwYX2UQfX93BzN/roC+VVRTm
Gl65rAWLUVS7Do7folfhzA==
`protect END_PROTECTED
