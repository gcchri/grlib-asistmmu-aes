`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gcITQYH3kbGkYGBMoG9tBE9/zMr6il4U6kcWvfGr3uT86wxlS8MDKLMUssxkMkt
CiYQpTtBCbw/C2MnQlHcHE5bzKff9x6RfcTwnzIqOD8pi7PNXuWILT49pg/Xspb5
bjciD4XnkuprR3Qoa0orCaiLfi7057erW0qylsNVdJGB9YjnkJcacJeKIrypeoga
cs8M8Vy2ydBJ5wrl2xFAzleGJneCMqfsK//Z6TzHNAHafuDmAytQr+EUk5Nz3o48
vtSnJCSwLYHLd1mrVgjMQt5LFNuhcLiN8tAtRB2p72/Qd6vYbhsD0sDwRZlU4v/4
nOSUd8VlL3BDbBfP1TDli9HQw20Ordn73HNNYIHQ5HyKLHnyDynHPK+04+R2oQ//
BeC6rBTk8s0+VxGngxaypWA9bVv3fkjzwDz5em7JCuFJCy/xHvIzU68AzJD1yioU
koe4uxKgVdMiOfFC/xz45FWvKOzTyMU2BsrEsIbqliJoFJLFpjaZ6U04PJUCHFEV
Xq9g+xbtae/IgTArOmGsLzYuAniuRMzm2PTBqcNwnJ+Q538XlYa0Eq3NaqXxzPPY
WKptKjv8107A7QHr+ezlNgdjQ336BCOVfi/4xmtYZQUxdLnxJQ86jv3bP1ynV16P
EFSQj2kQ/RjmchwdJtW+X7cH9NJZRhKYbRRmrqvy+D4=
`protect END_PROTECTED
