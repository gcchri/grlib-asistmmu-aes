`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wq1WGroC5L7mwHyzF2PKikCRvBDxwDTrVE0fha1QZ9FlXZF8/C5KW6hh5rfrPr2O
xIyUx1vREA2JnvU7+nj1rBGKtU/sg6w0N7luE6yn446r9Y/LanhQ5i6egbnUg0t4
jWaNUteWTk5F1VMTSfkNYTqS+YXPH8sobQlKLB0GYQ7VNT5XEnjlQYZ6G1AA3T3p
DONHVmg8iI4k30YlKgCHyjNEmeTLpAo/W4TopS7LxsOFSMveh8ON10MnzV2VpMtP
i77anLQYrTgqBwMmIF6gi552JoFYMm9Ft7YuIEQ9z+HA0pCRQvQAUaZrFuVz7jdv
LituiCWfmVjZHrRKjS9I7MqZ7cOqcRGcXNGyCknBbdWs6kL81LU6a/+MOLuTvZdr
LMoF73eDeFYPLXA1IvKSMRw+AnY0j06JiODpUJwehwGuXlDlU0nl6FHUBoGffbmE
6WT83fheD5SbZAQoT48ZDuBMU3bGzuFYDeP6qOedtVojvlt253/1AGke9CdlTSlu
j7VH6x9LtfLeeu7UDZaGq6vw/Ypg8+O5HFTumARfk90IZrJknFpjbPaouMZjmRcG
mCJ+6AidxLePZwDRKd77pGwVb1oF+iQr2iKIxq7BNBaN9039hDfEhZ+jyjcxzLao
YDCnqztDRBcML+vtiUhpB3dy+j61kJDO0vG4+UI8aQo8O+ZDr+Epk8ogDjf4AEg+
5l3EqJwPOcpwMfpzbK5Ozc8kYrMFIrH+ibP8Lhoj8r8=
`protect END_PROTECTED
