`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWhspYRCCxa8XOUWWNB/+u6yktTCZ9JtIEgDz8q11eXpkUDj7/wNGH/LkjtbmApe
t5LIlfeinjAZoQxufltqJlG8ReGsTCdKtRkQVgVUDN4VLi97b7UyBkYsXJcgT8vd
rLfKZLeD1Il6PP7AOZvMFk67nMrAythRl0VUTuxAsLGPLwVF5TGfWK2foqtZPofd
NzJkw4bdV3GSCeJBWseIBJKrhlNnpV9/53bApF07tVHwGjWHyJSGMNGq7s5gAklO
7X8Dqs2MmAZN/Ra0q2jZ+hnb6jWVTvCwQgvQtBMGKQptJWYdZ0V8s0aLGsZ5Jd93
jMgRAu2QPSf8m4hqVvNwcRnQZmGLVGg0HyfY6pcrlleykO3/tlR/P0sASSaP1R2v
RwcSCSrfO+lL/ANoocJJQqgkdXACqO56OADNGHKG6IDMdlvLw+4gMm59wUdMcTyd
9NBu6BrPfUqRJQrBrboecOm3Tm8K6plxdi8oVGRYCprUi7pV8/ivTOxuyCllA9XM
hU+yTcNN2CczZEOOlgytGy0noql9YOXxiwZl0e9cyVFMfOUUohHCK7wh4J9WYuX8
hTymVyj2F9QhAdD6Zdr7VHXnp1G8Y+l1kIHdalDl22bf5gfbN0ozNQx1ylyDuJkY
S/6t3Ip7DA+pMy7aqweySCxmUN7spRg4cK37iRZBq1i+UJ1gHN6HaZhK72+9+lWY
gKxaci0bSVaVXXp/qgY+Wv6LgNXGWj9J0O1/nhIRMuOf73YAFz/BkjT3ec1CNtm3
xDd4HrcleZDvay1xYJbcmFaLEBMg8dhzv313B9ZAOf8M1BIqIfJNssm/Dub6+t3J
NFVkXVfSsy4FIxYIN2SveUVQeNSS8awIQKK25UllS6VRStihwJRSg5XQKuW1aDDa
NXS954SVVJx2hMaDw7o1FWr7+doh8ADznzfDGWaOvh6fK8byEz8v/1F1FYWkeKPW
cqfFo9jL8MY7aKUFwntfTY33tbvHGD3f0VsytzcEiAQRg/1fiB+6cYDgeImjL169
WvoSpy4U5hiEpkPFcwP9rskab3X1ZD8M963Yxd/EM4DBGZNvswMmlFDjfltK6BGW
/MikZUOAs8LKiCmD5h5vcMUFO6aqDAVJchOsysvWz6df+uiUkAFLIKh5U4j1aMwD
dAxtc+FZnoyMbG9ExVI/8G7MtbK0+Av+6NVkuIP/WFNhxupMYAf9tPqWYCC1NmoN
pMsZS9aWDCj3iSlJIGJFejCgOVe8kSHbQSELilpVtVfy7J+oeksuPHXrtt4b/5Qv
JBClx/IOqrt691jnJgftGm9/0npZyIHkhiPyI5vnm+Qc5uVAQema3Sq6hgi7swT7
Dz5a3Y5LmOrtBvYdw+dovI3Xt4bz9rh2T7d/irKdgbl27MgLGsWySi6wWIZ4NRv/
crj36RDXYeYvnJ3t3HgSx6oGYQ2x3lG/WtI5Ho502EliEpIgkk/hw9OT9BeD8wN1
IdXZ4j+HxBalXZ3KQtQWvGAjZcjGNU21EWErqFt8fxt3PVp2LC/kDF407TRkN5Vq
Q0aN6T2jwHFdQxbYsGY8V+MOqWakabCua8PaBHHekrwy6xL25u1v9E3K3Ftk+2pf
DA6CMYZ8TAqXwEhAQA/klOHPpVNGJ9UBDm761RxveqGrHL48c2zILvmLnAFqQJ6S
dU6CE69Hh1cWAC4iqS1gAn0mcibpd92WqKp1mLvXUWTD5poxp6jkLQ/UsJkYIv0T
C5hjli3/VDoQi5XWrzljOMN+EDzqPpPbSxVQpVWjioysg3ZfuDyTjujpsNXFKYXm
RzQ5+RsjqMfIPxgHbgGzRBeziBlfXkCi7XnTPQoMkuxe+Sjrb2EpxpDGKSvEU2as
F5SRNC1HuMV9LGKj4igEtJBYcXBYhF3z4xPDk5qubQUWs+v8zkCLrQm0pGgyp3WI
/TLoLkiGFJl4MKhoNn25i6J6aT/0PxB0IXmWKQksnGVQ0+cEkXDuLYnx+QEBffD+
AcC3gIlv6u65JO64A0ed9/KVoFCd57Q473UMXekFdSesZIYXQr/tiLvxlO0mMoAU
Ab6VdXI20+Fxg4/V/gN5Oib5SNR+TzyupZWXX1oAqQwLloNO/72uC8Mikq/JdVWb
nlrpZdd30+QkePvzTrIJblMNhE+uKFsww2623D4BGXWPhFub1GOeo7VtVVb87YMz
fTzd+w1MQ1vtvSfKh/Yp2Wkks0z4+bO8WW+7C4JZJxpZdK2zlbdAyJXdrQHizelL
4kxWKFFR0kgl3pFFU8G+QDT2XEBLu6EpyCssxT8OajfW5hQe8RSTZdXo/y/XELtx
2LmwS/Wt5qmmjyrHJSAhxeFpcUvPyzQKLNKD/Ss14/kFrVkzcv6XjeFM6p/KVTzF
siQgMBgwGse2erZq6/ieAGeaad127dg9ZHDBB3Fx2F2J6SdbPSmZ/wqHxjITD4i5
LSzclwC+of8Sm+khHs7CQMJkQBDJaMh0Z4Zm3XRyO5GjmEIxZadoyhjMW1Xkrewl
6ax6JuILgIKmqessQZxwEJZ/7VqP1zkyvTXw9T90IW4oUU5OloQZvOFuKVOf+9EL
pwP1scBleqtnO41Bclgt+94WSK75ZoIVVKhXnigVJ/cySZFKg04xaXM9SyxXRH9x
4woNbWI+Pp7sulOKeAxqlXiFQ9lq7qiJRIrdUNNVYXGveA8MrWOoq6qCZCClw1mT
TK1d/uSQ1AMxzxcJdHwo/SOfU0r5WgmxG5rMTkebFw9XyDKBgk8sZwm+ahP9Pz1Q
lref1+t7dgugz0a0oVcgZz7KEezmhbxOJzFRmLjPJiPnKhwZvaIswGWm2VK27M21
OdBIkUKfTPP2s7GRo2PLm/8xCDPKch+CGHd2XKUy7sd1dgc97VW+E027hSzvhYhL
mtAptGk8cnumN/PJFgXJskPB+jucI0w+Gyll/WFpXI8/gNTppt0U9p4NTv+zlwRH
jvm+McLtVOO3/WurmCPZtnjEPyyh8SpuavrDAmupY5l5fwEBd1KwUTPF9UngRiVt
w/W8ERADvMi8TXZ0xwN68QsPJZeFdn8DPjiwUNeuZgJ64JzNsmlQkNAMOu7K1F0l
mRErH6kq6Ft42cFY0q2t5VBquntiMXbocIQ38DUWmCCuSdUPAE46DrSwe0674mf1
NCmXQwd8i9doMYIV7WkCbIjGWZSGe27YJXNlzR3J+vSKRrTLxEpBry4MjqJVPL3j
IiD9UqvudZ9VCNyoQqcxpA76J7nnWfxXppAENqf9haqQd4zYP2DK7OyiK7fsCbMg
TWOSIsgucnQUl2NKLTFK1UfrQRmQK2updl85l6lnkgoV8wijZKh8dgJZXdbc62CL
i29DxmqAyn2LkK9kiwhzA4lHr0AqawNxEXKI137qAj/DbVm2ZOE6Hdk5bnLRA6NP
+UAwVDAehdC2bGrwa02nhh2ZDdUjg1FjazwfRERtf7Cf1d/gU6UJFrY4UohtZa8I
HdZ2zpnpj+aZKhQJ0qzjgBloFSAYJMll/BgpPJAmSnM8/EmBmr1YAx2FYQM8Mr/v
1oIP4+kGzdSMOavit37YlOB2OHbMgmHip9QKnB7SQz7xgawRCjUiJ0o/Ho7Na+ea
IeEiJCm3xS+feftjTvF43w+8uX0Yi7hEn5m98mhXzTrYuAjpcGEaxg43To18B6DD
F6n5Mf7VDdZsR6cBjixEMlU1jDRsEw9daFh0MooPnow98rccMe8Sy0EKYtc630Gg
ZT8lwFv+0icBL+r09S6pSs/Vos8mXWo8IG5yVp92L9X5SVUccHCb65XrdIcvA9nQ
GcBeHyFKAO7fdEGDPV0LVKAWswQL0aG4/6dWsf0sSlzfiBetaZaVejQfSY+NZ4Bl
9qvAiocqH96IKpcHlimfCLBoRaaonHtWLTUKt8HRXwHnCxUoAp5g3mD84csx8Io3
Fw41+AOecnV+B+6qlQMWnpI7zBG8p5/fSfEjlqBanU31lQMS6Z/MeKfTsPtb+IYd
Bw8VKj3/N7796YbBSxxckvDUY8qKvSlUaUaCq6eHB6tAYQZKGNQ4FuPztmdUROxk
Cj1wDsvYrlL9lHbFSx0eNECuw/hkwxaxVpI+9lj0iuwnvWtsE4yldWZelG2o5WIu
+9F2UraFPFOPUI0DEwHyKcqogOha5GMppKElNSfibzKNlFUagMworHxTjfyTR+ss
Q6P4aWR3dY1w6LUwUSzGKX2aw9tBN7bkfVJM3iCfDPGI6KIfu6qXjWOH0iwP8kiQ
Kc404Y/r2Ee1do0r+FhRzBO5rkJngWo5c3VaRyx3Qso9KJS4Ufp1N2UYt/pAc7/c
Yc+0euZkjVMxm7qeh2Vr3Y4ecFETV5VHkXgNwAfkVS3s2r7tZ3Vo4lc0kl/QVp5j
RCVKnn1naUhGba8bDZfv5T40L1cs3mSytMad/fjVqAua5mJ38yMeNwZVxVWJfdQu
cCcKr2RauBSSzewEOqxZb0IKUHM/XoaHNAfWbYbLP9SxVdx7DPyQcFOhDfaefQQ9
EomeOpr4QEheQ2yLrLza1vwMnXWOA/4Qb0jMaWhlb5sS8r1U8rVFDZ9bTNInsFk6
ly5R2sWhBGrS1obBlTtJVviDD9uYynK4rb9i6qmg6w7m8NfCA8MN5VKcnS6HZTqx
b991uJAr5YS3VIsKu5lD/LNICinSrYH+81DDLaZSpezyB4sqnmaUF4xrw6oBJZga
3khK/FITZ+jnJ4uvU49mLD7D33a5Ykq/8PmrgL91fjFwzasQ1E9x2J5A2RCGmcok
X2zfbLt3N472CZp6U5HMJnaaVWhm2uE+hmJqS8bDdO5+qhmH/pwgiDuvQQAvNh9P
BY7TMRAhO5gN4+S/iLOji6wN+ucBMKgg4N+Pb3U04/Y4idQ+cU03f7yolmYLU4rc
uukwnhqF1VWmLdY0FpoZRTOV9J4KZAzdu05QDrITLyqGfOrmTuL1IhY6gNgQX797
OP1j8rbEO3eHuJesHbd+oVFZLRc9r00N5xvAcZP0IXl16xner9YTM1V2wW8hoFkN
gUI0+DvC9qIs//Velxg0YoIuo0ZQM4Ho6nw2caWzdlcy4YqyLzbgZcE2xuPVmJoS
tE8rkhklY3mEUcrB9BBeURgyupE/VV3Bd6NeqYY5FKchqGIGBW9GhrLEJ7Gb1/2b
OSlA6vel38NfzDMoIb13DhWUiePyWL6oTUZZyoU/7aded142vYKPlLeU+QikBLJK
xHe+XGkvaBDVYSsL7ongza1+/rhL21su6g/8lx53jeM6tVlYIX86qToihSTbpmxA
fnwBGYd/NrMOlA9V07NyTUL9SBe/FoEGM0VV/nS/JgFORAgWm1v8lY/yximy9/uN
x6SDaf2FdrE3ZLevbSXtTXGwClV+IHOufyvXP1ZiAfsYvEKIs56aRB3uAXVXF5SK
FZXfbYwacsIUrl9RhXsMLL8ovVW+88/GJJ0Wt2lFuVgC80FLApoQtfhJ4uX35SVL
WFV5NakaXAsOLOKdtREtY2EVhLqYut5jprnUf/opd0ocTr8AvZvhPVq5pABix18x
9PGd78/h7meGiiRbjYM40x0DN/ff2fMb42xx767XoRMf6A7ZopXQq/u6H7NmiwlA
3xnXknJ2xvwgQBJy9pA6EzgkqfSgp1Mu08JOQeLP1fpywdTNfSf86L+SGIwgEbHD
LVk/urnHGopK1gVIoRnNbZmMYoA831+gmf1zYrex5InReE6B3aBU48sk3kJJCFym
7bSme3IoMxx/g0TGXtiU0d5jprA95aF62xndr0VgPmnQ4lDXcc9Kh2eqhDJmYQDQ
tYfZJGmpO5xoBVjU1Wm4WIW/72d7W+lEDaqWVG4ZzbOQWCIpNailmtkpqeyTPJN0
EvXj2AAcZEAonlI8y8vhU0Q2hh5onvKcfXtJwxvU3MJlzWJgJ/NbhSD/Jevi2X2S
447EjEXnhz362a/4EIWDoJ/A4mPDH6Wcvh98ReHgm1ai7SYOMrLUxtqRK3DPsKAy
Llik6q2MIXObsvawb/5QyTZmt0PYDUMopOYEtIRxIoADjNhYQZr0QyXSKAHIXJuG
glTn9J9QxF1W/rbXvPjoner64OfSJIGhjvFXBFxwVFLqMwU13JtVvyWvTZQxjf+M
R4NH8JaZnLRdXQt22dPPTg769LwM3j9yfmrhI1O0ACLVTFhzOQwTwz8rjdUVa4Ej
i0Ca/BbxZXXzr09TlKIZkzFqQLRqyPjj5yFpvGmFgdI/S2DybcqW4CFUWSflv7cn
FxAlEO2N7QU3QzoTixqQIin1xkMAtgl/ZWAo54DECXfLJxekaHWhTp+QjkJSlKTS
o51Ts4Yo9J86UzT0IGGw2buU20nQWR09p8+P8BfNHPzj7aE7+qMh4E4iFp3K8JNe
LnFsM/NQhqyXzmahBYddskj/8dejBEWvLXrYS1/PkBBTwiH+tu4IyosqwhDj1Th6
kypinP0VXcf6JEMe1MMi1ay7tGrqjEgr3NSNyUfJC3BAPr33vMRgox6POKmlHDNf
vsDwd0fdUR2JPT/c2PpnbW/0CTUoYCoG2rzbe0FnAat708UBY+QLsNUO7s+TarXC
4m45YrrvbBSOEmy8rHxMTC4jf6I1ygibd/FlZvYLqGgCCrNbzv1BmSM6TDmkH4pe
nRWBkV/5azoc21/S8dgbXgCYYOrZK/XnB8P3AxuyYH+RH2OK9PPUePXc9XWFEnrd
AJtSoKhhLb/cuM/U7DUk/JOFb0ijFfQ0FJvXg3VePeqyeszujSsBVHQ6Jc7h4Jjn
y+5DcAlcQrlbkaCjPaomLkizuBUY/nYXofyiTMEF05AmZFe/zVz9gcAwkH8fuXq0
HmuyUTlXqyWmTaEdJlrV70tW8YFETRChNU4dZo+FDQMDnaiDuIc/39y/cRcaPqYN
beSQElpAu3AheO1cm2rqBxnafQUe7Zhfstlke4/YRRXCrFvVTublg+esHN3ZL3mo
qyaNj5ZG53WSWe/Jdp0+MLC4wXpjJabDyJCLiPXNeqWCgX+5BMtWP7IbN3FMl0SO
Q79rawxgXn1h70IA34l3jlYG9Pbg22BocxSDlhsWDaJiBi5jrGXj7BQTX767Y1jc
0XqF9hL1sRXDsD1v+rgqCLqkXPO+26canbZm5MH2YlSSdt0372bhEdyAVzlZidd9
AfP1qvIBDJ124EdLlSa9XB0+u0feoo7MleV7idzbWezrBGs6zrBQrpqlWxUlAFLR
8NnA1eMogs+5H0xwRzDJKp/Gs/GMunFAR+YsKk2ZQpWdq21bR16MTLVko83bh8oV
nyAmwT2dyKiB3PSGlOue1E6HxVfme9g9txg0IZStadsLYKuffG4HDWCNrL4JBBzt
G9ysg1qCR5RRSsZMCQ5HV+NvAFjH9/X95dOMpbQNxvwnWRMWDvZizi0QXFO49u5X
8FIV4SY+t15jPxKvz+shWxkuVxjBYuzJE3PrrV1pbCGZ1vRY5Mt2TJiTJdxZ6Alp
qGntxJ1giaR9xgPRHVj9QmKsxE4Nc6I3htqvAu7h4TaaBODWv5yopPtf+oZRC6LH
tTVVVe35NYbLzKGDGLG5PWz/Csadf6g6P2+zhyUZ/kZUxEeTMlHnlxQmgPyp3Q6c
ubc5xPaNjzm5z4GNVudAC32mGD+4YE6RPQGCoZxjHUobowJLKehI22VRTgQ953Yg
H2Vmap2CiXuJF20IntcWeSamvdQ+9OaAxuwgd62wbLQZuEb5GQjO1XcCI7AcLF+Z
+h7sPhUkKGkeC+1AYNkO5Jf7kXprA1UM4VaEJItbLjR9wvVdeJ1PpYsXRA7Giw42
JR5t8hSU2PBc9s/Wmwp6M7h3C2KpSWdMiLxt1GC4F7lep3ITbSmXIlDcsxXUsIjI
ScOTguvJ29vyYDBbDSmmk8ET3Es3fr6grxfdHYO8m+6UDjXvVQadOGDiG5aBj8MJ
8m3v2vlQTMTGEmgNh0fRG19NxwWqC1Cx6n3rWwzaNHfI25rqowZC/u7DUkV7CfAQ
fyqi1fpuYCpLQGBnMs5J91vnhFBhtYmDL1MflCGnvOOQQIyT6CR+LO++p0PTqDyu
s9sDMXtpFhwmmJK5VAo1pUalsoXTxqF8WfDCSDhWdr6puD8hKVJb6JuoQXdM35HV
2VvV+FwUMqokOJJKlrH2QlH9aEuGvKNaZebi+dy2Q7Sj9abDhqCAR0rGM00PFCEF
80db4gVzwYA3KsywHpjtFplhDNXThzbHWD4YaaJxFbyR4/pMS1zDtZwDN5K3okRP
sypWoI2VPbssDanMWYtgP+pIm1kJrXqtrABZvCdNXDTdCCDNRUa0M3gdpE77F4ZM
kTey+yMIOTI8vVZSwbxERR1imDLlTsBkurJcf4hhq6QsDlX6axRHGi5yYbR71ELG
pDfkYOSFMRVy6UfzYSMtsfV9bRBIXaE5xZuGgfmdZWbiRtj/UQSO6boSPFFjrygD
H85dGKEGgLgdiLkeVHBxShCwRBd0ku0JHKKVZWSO0pHztbmerCBHILS92ze9/xTt
83C7/+mF6aboX9xvcfkNfbJZpgoYhx6BS5VQsCeGKV2NM1cmrMw37gofLE0B1wFL
7O2abqylzNpw537pHRjS84Rm6AKaed0DxGaCNSZoKTqAUQpJVpcgZ5zVHvBLJrYE
I4WkklgxhsN4n85XL1MQdm96dlyfCH5IvPx6HPnhfculrpef1avv7Lsbu2fN5vS9
3tFPOKVxolxgNIggbsuWuqio9OeMzqoEB4PL9dy7Y6WVUIEUAUsW0CQGEYzYaI5J
YTDIcC730VwgLO7rRumZSeys5Ed8Ohsbn1b036edLecgewhgofS1d/B2rGFStyxG
SUoPD7zomkqXsbw6XHKNBrVA9XnPA/1mdGF2bqobsByDYlP8AuWyr6pJHEwXXtQK
F/qJ4Wd1GvBTWzjuGWSecZMc1GQWJulxwwG7Q3Umk2vyHoqaKz2w5W9Aoq6KJAej
S2iB4bWjWV1l+Rrqn2d0GQgE5PDsvB11iuGV8C79bZ/NrmKH9R7xQ0dfAEqglvvU
YqqoLLJPQrz+VchWwDMxZF+ujWDr1yuPwMT5HccRgSX5MQzD8Gmp9iilHOTAFYTq
8eI1AdiWMWZk9XsQ9F7IdjbqI/D/oMLg1C6DU9ApyzJg5/VdASfB1V/dREEEPMAF
REr5eQawd6v8jxYgpDKqfKZYogasPnStwAP/rc+RD/1jNcKcNfKC3TOfvPJg5+p8
wxWxXKW7/tR0RG4weZ4OGc5Nae1get+OSOrz4dHKcCMLGTqfuB6wIOI6AtAehsIJ
FiuJPQPlbA+FuCqLflBGWc2TiB60n0hgaeAC1T5kpY6oQvd9516ki80+Aft9aIGP
mLwYzeuz5E0+5Ptyj/mSXstRgIofiUT5RPdFedhGusEB5WkLHerOCc9eMG3pmZSb
QILx07HJyX//UvFSlgPtLaaX2D7/uwXZSwO5lkKqoqNrWn3U9/JGnn+9L9/sROYt
3QVYSKS86IFZ8ql/lOR1c9L9IFf1znrUv7jNj/FUG5O2qUrenTyGlgvDfeQybTEe
QTCnnv8FUVQpBycRZ75F+vjOwSffIH64V6Fp7Ste63nhdS3AM0znj2WpZnYbqM9W
yVAwJan7bX8MOjw2mPu0Yaoc6TCmRP8mb4Sewdkjk2tiV9IJoR27NkEWtUSjNl8f
ZskNSGgM0HORzGu9jXGvqD2b3jS64STWZz4wWwkMW587/AvqoV17BYRSRLZvbRNX
j2gt5YLylNGF9TbxQh7XmOkb8YssIhPJjCM6A3WF4gL7o8svmDlgNU2McatUiZQY
FAiOB2toGjyQw45AhP3PKzV+hpgImpDs+/m1/lryrOjfwYQBdlgTK/UNzZzjNE2L
uC9U7OfcUzQDsGSHUNTaxmtqWowjKHV8ArGigmG5c/yTMC1IdI16c62i35Q0zY9u
GzhsuWzl/MIrDWTOvTj5aD/hMmWlE6zw8jvxhOL5j+faLueXJEBdJUS8gSyKI/mw
p+iP+1Sus5ig3XNCCaIJ1a5+V1Gs35zkSuqVuKUxUG8bDS5oUjMKYH1bGEDnOkCt
WVT/GdGKO2Bl9Css/8pESXMPD1Z5bkPnehBmLPqI77q5g5YYcOTiTKizq923vkX4
xjoKoiiFrQXuWZgSdWJW+R14HWrUJtnG+F9FOMvxcpOHos+tE0TyIp7xuSUc3Gis
e5xhVjaC+pCLiYRoQHTF0ixiVQPiBAHL4C5PUNdgzIPEQDBIXdyCbe7zoypef+fH
EHLDkF9ol6lZWR6lUVuqTbrmrAZI5czs8OAsfOUOsliVBcBmQw0tJOdeWZxjFbc1
hxaf6OY04OQ+c3GT71JsyWri7F16INW+apYIzNEtzMwmtC92Si2Ln+hr6c400dRj
Qq8ae3vlbpyXsYArH2wiEz9kbZgdqYGiaxzZAOYbs6nd4ISPSl/GpbnSUI4W0zlk
umAT6aR0jDxN/A+wtUs+CjAuv8RBZpOEGYW3t6Wg0w2Kxr8sT1lh1gYjOCPjqsXm
nuUu/eSrf/v0DPSscEpr85lLDP7OjED2Hel9zq9LLKulgMqW0ab/+NVVNxGOk5VE
wWp28us/02pKJjwMPjGObvmi3pQPrJrvPpHnSLgbNUEOOf4z1C5Sc4v+2vOj50fF
7GT2N55ri00tLJN9YLj/64hsDSGkPgQuDiwhvgkSAL+KicsPPGYQoa28qQOFd8De
2cLz3csV1e/GPDWL4e2KpIRXfN0rRCWVBl5qdXqhfJobMI3tHUSk+vdU04FkOQzf
kOk3u/MLxlLvffvpIlKk5USRADunhFXc19u9VemxVklNL/1Y7b3DzSlnBPf963Wb
7foJwbB+B8VU3vSqXAlcekgQIlY7vyeMFbH//Q9WE3huprVppmE7Cc1sgcOR+EJ+
ViG+REIyU5bR/MTjGWWlYoxsRYauoa03OqF/NAuatq+tud+7Tkj+DRiyWWnw8AmE
eKjFkxzut7ScywLtVMS8T5LcG+bRqFVtV5zSLMuM3ttq08lHcgT8JISxgShJGM/G
fZhKpESABFY1ZM9+ASAq9XFzEaRo7nHV7+07UVvvpEHovvC0CprHmtof1XLsMt6Y
9c8nBWeG7DjUPiMv2QTmEiRK3qfYaKOAeHx+MtvUmNkla4iVYZvQHNcQJL7VpwSw
2lq60VrKE8i1Gc4y96vYeeZJP7Wnv5j/MMx6b8E3sPXKMZtKw5+8Iwv59CG4hicw
uJdqnS8l7COx3cAR4I/Wp1Zper/VcrVEVC91mhA2CKsu+Izbk0WUbvGVuk57DUV6
a5hdIM9beNnkCicYWiqE0zRMR22tyfUX1qEM8EbbzqkCiCiPiIR8MJlcxDoR7oWB
w3pdBSS2gbCvbBg3qhIR0q7YAPkKW2y9DqInjVk5yjTkLEb5PMK9MZQ5dXCb4pjy
2uTtagU4n4QdXwvmFPi4mPHWgALTI9g1rVtS/m5i8IQ9mRoQ1gYMsYeSKTvnf1hc
lLDGe4WxZHteJcpQmsmCcK0RW4f2EzODlZQvxSVM+LS3uyfcgZcUXqPVEVim+KyE
9Oak1CpMwGzd/El45nRbDlivNaNBB2TLHHTnN3mElTfLmYO93X2QWOzbil0oMdFS
f1aS43NB+nrKJYXzjd52NwDGb6e473c4rMcABcq+eHN6WjOXjzcgh+KGfguz/oKe
2PRK0OTCoMJwjmuRh/bKP3ir2Si6cxbWqK357LcE2HEgLkrM1KMh0/kgQP56hdMc
qMs0lkqKUVJcSmH9zPaYRCmZhx4GYGjgI/tdlVqcM8ww2YFc9UotQ2GW063FHVL3
irGddrFOYdVMqHYxjeE5CaQUDBt7OId0B/L04aY72zVNJ1ldIDm5arXt1vNRO/HA
3/fDP3FCkrFWSYucrtXovKB+/KXsE0zXGoISj9CSfDf1k7H2FsnedJj9N+POabgT
qsengDOWrkRfmlPej+evhfvRweB3mRufc+vH4ZjEXdVmQzoWR1Fp1mdQgkgJIhCw
V7Lk9mdM0NEeU1z4tpH/A3T51Pz5sNJIYgvGDz/LMrFy+zATkBTx5Mr3Kxzei1k0
6fWNMcLLFtMRWlOmYb62NO55yDlImNjHfIwhvCxua0gBJQmcf0qdVn4RvOWVfJBB
kqeHTCPvpzPWquE5DcX9Bv5MquXINWcjrI6Yg5jqTZM=
`protect END_PROTECTED
