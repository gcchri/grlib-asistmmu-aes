`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9wfi1s2vscT9lngUbADAsIhwVfHQwGJInoHBn/bKg6PbsCH6rXqR9DRtOYptWg3
eWK7x4sINm78tKcpdbs+JRRGO+yYntMfcYMCn5TdS7G/hrfQILufZLEyFl+sbhhr
Utua+crA0IBfs57Kann6y6TKO5iWy2waBGsFYgZRnLh+yAEeuiVeeK5HVHcbtkYR
HfWpWKSE42+qS6RcPnLyw5CGbPKB9TWzjKM6OpHzsDccO5i7Z4ADzZf1+F0r6zkR
FiwsgpMAtRg7PYqG66rzCBAk6Oxwj+jTFb2KlTlFScCaUBSSHkdloqEAvzw1YgAM
lh1b8r0+/T+5LugdMhWY5Q==
`protect END_PROTECTED
