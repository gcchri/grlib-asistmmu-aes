`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jigo5hvymMWJf1R1zBkKH7H06LBGvEa5RsLAAVjc3une5cINAqtuDM7+3t6fpSXC
oSmq5lpP4sXH8FKOzMsIfHqEmbqDdtFAKFJOr5zNwhU9KjHIJooHsJQK3ad1Prpj
gxhbCdocbfdHuwRJlxTH8hjWWw8MSNfjwe9xIqWdnZW4WRhhBfgyKiJce8XyMrAt
0z/1Ge/5SQSMV0Mza8jE+7Gu8kb3FQWhKNz/ow+W+ErnbGz9g52r/aQZAHUpPUIp
VvKme+lH7nz7fe7iE6cwWWUyQGc5FfQtLZrIxB6cArKG1Cl5RV4YklkiFIM00y4q
Geo94B36pTZWLBCiAYsTSBH/zlP+jsgCEo44AfY/FYZKSiz7a5fOYjhv6r/TzkW5
3LRUNLP4uVbEvkHu8vFlfAmTb/itHmKAZVoaADYkwh9NycB/NTu41fhLIrxnmwX7
aGZShe8gWAmmyFj795L1G/+evEfCL3BDIj3kZSK/M7Q/L/SlJpB0oDZRFFvmMRGd
Y63+5yTklNVE0uXjklYQyWn6grU2Ue9WqBtilHvByDc6Irht8UupSu6MXpx4KT9G
PfjZtWHTYCvl5kMC79yypgD6Y/fqhBiPxQGTQm/JuR/VaXyTNxKAjJ77ib2RKaHO
6dCxM7AAJD4yxL6QdV18ppC93UEou4I5Y6A9clR5WrlX8yC+DUGkfL0gexw282hF
p7h9JcNasfW0csIpcA7LYCFgQaaw1htq5OAvKopf577JovWYsiiSayc/fL+YLe5W
2c4dhqWJDBKaxKhlRBxFos0S6uQK55+mt5Ytrh6PfH8J9WfAEvgdhn4+nBH49XDL
1OjTyJmRgavotDqQedBV1LxYHh2kj8UBEWsOeUZVW3b+z1btHXdgvo37ZhFLzXT5
6I17VkwwKJtd6UwzEVjBhyExP/ZhGzn6GuIM8oaL5H7j8tLk2nVYyZhcviMRo2vP
TPaVT7WUPHaahlIFXJ4W+3v4Z988E8mkAZuiorNrabUU1BAhg+MJXoT3MchtF+ox
puAdbK40xp1iO3v4MiXC1eRxyw+fXxB5VAAzH8f0jpxmBkmMD5DpXrr2Ot89golF
KnnwHr8PBiMudK84Er8vNJ9kBBFWzDAtIdhYvE3J9DtEuw0GUs6cBn/wDrHRVqVP
a9a7YVaH/FsirN3oQUiy1I0J9ghGj0QtbsEBh/GATXlgHYepLjMulO2SdHKdvu4G
znC/56WdfhTbFB5m+rADOInkpQHhRP80+sGRCmIpk+E/cZWinxa2RWLJJX9RYtNt
/KX1AQq9nc4SmbHxyHh1xFxNmQOcM54JLZ+jVEuQXf7W8Lv8VuPPEuKDetGcK4Hn
0yAwJOcj+FGAPTl6BLi17ratP7zT1DZ7r5T/95iOIHp8uqfkH4GqhLwskboILfTE
lYDHSmQsX0TYJWd+jxChE0DRnpqtKRkHLSC3vDGSCFXKf2W2lmPVJLwUp8o63qBh
+ZtV6gsjG6rRWPcD1Sm77UpSWAtjAuwqtYdr6k9o0HLWIFuhZTkeWoszON2KFifG
zKW3Mgr0PQ+/748tGFbxPRC0p6tf/Y8WP8JsI8TErC5fYMQU/PbU/UE1TeSeNaFT
RIunk/Bak+3B+vM/gXCFc+Bb8p6Q8/3fuxOqtl+LzyoAhDvAvYw7KNiqHC4e9iBe
ek4TD/RRDVxjlM9vAY6ur2Dnutyq8GICHZkKZNIHA55FJK2o42MNIXn/O9uVPjIz
cJjyWkEqRROWjd96RWOjPHukW3x7zBMNe0aXTx8mA/UNKA9yUYDhiXUAHnCLrpkR
SccZr8vq+TrPlD06iaR5JdMpeQLEs65qx8rJ/ABrR96noFTJ+LGVzNyzjGsYJuE/
Kv1QzEiCFrSeLhi8J4+TlApTGxor/bgu3t5c8EvQuO/zv4VJifouVf1LP4U7KJBx
pV3Ca8mfir/JV1nC6vli/Lsxifj6uTvwsEXPjpG6d/xr6X39q260oFFmBrzCMtCq
OArGoZasGuvutd3g16w18JzIACfDPWtJdpB3MY/eA0YldeBxj3m4pkL0tg4ypbWh
MNMRNMsgCmLtOgwPl3jvBaemLYWenNulSMErjmymKPtb22QPlrZJWWbFEl155B9L
t0AQu8A4JBi7RLRUw2hgYWLm9Dk+Jtru+c8zxNbTRzBjAdj29L0nRa43JDUPvZjQ
WkXEvSsUIkrApQkbzXsox+UminaYH9GEXzqOla1zzil294+BG990RYyn7aNmhC1T
+iiuxzaHzG2mlrJBTmGTrC99vcTajqLF0LavuX7CJfy24tTpS4QTwcn2zulrQEqX
HGx/GDdSvuBkJHgr86TtoL8e03rmMT488l4KGCdLJ5ffOTPqL3WmAf7otpo7irL1
lERC9WeFPLLwYOOUA+aSITdyN2ygoejySl3HZHqfeb7GGV6kVqe3C6/pFt1GFeu1
ywgPT4C3MGnNL+bZggfjZsB9uDJHf5PMlQ9kxa2j2LVz5h/VSLZt5OYatUM7eIE3
1bYLQUqvBIv+O2CyeH3xvHi49ZAZgPiEnQqtpOfMQmLQRI9rB/cJb9IvmFWcSaSJ
vB4UHohQ2pXRKUxfbfrri21R/OW1iRAEVIOGMVfwbPhnhq9LoPc1hzvVti15X/r0
gHcoc/Qs8D+i7izqxTlq5sWZdQMkk3JBAQ6zJWuSAoBKa6MV50R++GGqwmrTiI2y
RCxW+/nhqRIdElQKAoIXTj4gSoV4+Bvad0MBaLmmdbLt+eZt+/rYMiF+O9gOn8lx
SwsD+HG+r7263SlqUr6PGt8sDY8RkMyHsQ+mnSbzm5xrLAWowFmSFImX4SI4dJIk
HjW/d6J2+/TzYrzmAvN/J/3tgl0KUNnB0zICL2FjO37xrGDw/a1q1HrnNJColAcz
HCQUlFZSnSE3llpkO+QE4lCpqe+JmMEpg3X2jrCQpE0/KuT9BFZ3IBz9lAIKD0kq
9uY8BXWobmcSmfyqCMAIn1NEfhkWeDUQiuIz0hX3mrb66rHr66lfAGYDdTxEmL0l
PDgsW5HIzpnH6hOwc9z35j74SGamdR36MHjLLuAYMbCVQPaoJkhiQWtrSJPh3kRH
ng0qbFDdrkexZQr0PULoVbL5TD/yfVndB9ShUoOdHIFjb9farUxW43+tWvHeZn8M
lbE/1RXc6Yo8GUyN2/osdFW0bd25YfDByy3NIwLDIw/8wub0idnDwcLZuR7iRj2F
gHxNLRAWOieO4sr/7pW0wNQ4HcXraB4kge0fCYT0LYtXKmZsRNBhfx6BCIVwsPeJ
JBSIwvLZnR/yPsRTQTC+5yf9A3h1/33CxHW/UU8cAa0Jk3cRH/jKInrDvGNUrPZ0
RL6H/cEr2BTMWBvyeJD7ebjbLn5pXxIdMjFAHecjkA9zbqUJvP7P2ylnRIDCDXPZ
xA8WIKwqDPcGt38Qt4Fr0EinCsgftBifl3yaxWBbQn7x49mL2SfDGiWVZwUNI7Rw
m5EAxXGeuslt6kjLy02CNl8pZjWQpwMNo0f14oz9HiTxi148IGwBoc6UzuZWi+fZ
jZeVedVJfKXEgHQV+p/EbgthqY/nuzyYN82CqSTT4dJiT3ro8t7mauZUONuncgEI
h6a2bmDvAno1/V2QEWr39gaWxWzrz38cKaPCLCMoZ+eS9bzOXXjhF87TeM6tdJRG
aMNnjx87SkHzh7qPycRHVOnJ9mcfwUsFRAI8okZjecZJhYU2A5o9fHkCH5xiALb8
mLM4b2ZPyaLlxJlWcGVqN9PzvG9+QR024woUDbyjOi34M48yevM/rZ53fnznWKHt
wED9YkZEQtney1QySm7SENEdzRmdzcXtBiSVb1LJpF8TAGjpuIARgmE23z8HzZeC
gbwef05pFWNBsRXN6h/noszFWJeMIJMMMTek7I3jHlMIPdIjPTKdLniyeWMfF8G9
YfVM+6dXd7Tz/BIlzzw6NNdSq9pactIxJu/BfBpy9mf0w/hxD+cjM8z0CCiJnBOk
CEG1Hra1NwW6ifUouznsF5tLixphN+9kGu1s00AD01wDNyTcCkVCq+XBgthReuMk
gwTmCEZr9Hl0ZNBIe1WFdJORv/oaLpEqI4/aOH3Lnl9YTp7fnNZz+02HZ3zq5YVj
o18TbRqyLfScnmLfyMs8NcL1QcKpBCdiFvkpmvuprINXxe+09RiAny5QrHkW22ci
+7BLg5ffVhlsWi4SEinkWoM/WNEj5xK6ihcy3Ycict9dnfswrzk6vMkT9rQifEME
Q12KJTgN0M5PaK8X1EqfHE3gCG1eJ6vlb09n46ZkrTFZQfkVLEtP1uQotyogtcE2
J2hEK2WnArtxFr1jn2+zFtMxpcRI0iW0ndYTrIERt+FyBJRH+sU4L70l2jXO90ic
LEG/J9P4o3UwYBdjo2twB0miBK+ANchJA1KYCemK2QkQkiW4cgHw4mVH6/2+kl2i
uli2O+MMHY1vMau8aNYI/iJK6YVN3SIdGKkolLnDovlnieoKQL5wbHdsfCboepMk
ZyVfR0ErloUNQQR7Y6BiZB8rNncNvnlZnoGcxgcDfupHKGAj4YUuC6U1lyM8v6yM
4aCE8LzfPYHhI+DQsn5qvI1a0Qo7XDQoJdTnuEtNjvHm/dcvVFLKV9YdyBAnxavF
dm1KoOwUz/la8OZlgphYbjysS5OigLdMbRiUnBkXiwWzIQIfb3af6urFImfKGfvr
MCXJd/mRVJJrakTMRMoOp5D+/CVLkV8jJrFXmhhT9TDE1Ck9HTzS3wxVVbDAXZCJ
kmoctWmZ/ttjdMO0oRQ1U9hcmd6TT8DHxSUKljJbddcZy/H9stPF3aDSjwr2uicx
tM5yM4OObL2K+sc8H7AXqIqEARF8Cu29luCY3casypk3ihuNdL5REARcd/nWJUkJ
TcYjXZ8hnjP/scUSVuuRokmcRAnbYe2z0u2p9xiw1QJ2A/FFNmggmCa6eoemHNlR
2CtkYwf9DYcUzk+dsKgskykZcI0SZRV2Joa80TkeSQ0h7bce791xfdvBh0cM/DnE
aI9SjuSfF1OHq12FyJ0bmKawIXbC2/nFlRo4y98+b2mzGjBR/BOBVkixEqnRq9K4
b3qXj9sU5ygY5hVX9PY039DdVOhtjH/qMteAhXfygEP4KQNTh6iGalDZa1lDMz2U
vm90FVyZyDFm9AtN3tFJWcr+R8goQH573zWKi3VpwAT2GkimmG/dII/Y3zq/1dLG
skaII0nd4FHS4WMOTSttRy8g97nmQRIoZHoK3Qz3B3EWnFgAtDMLB+gUDxXFgm0W
FXH5nziOyk8JqGRDDhPI/9jDlYYpIgE2DBWqXQ8ahgUV03fS40dhRdgXZsxsFbCK
ySSlWE39xvLbz3r0ioOzsHPTMrSpatnSN8fnEvxcuhUKNkljYtC/I6Z+bkzs6T/8
hf4aruI/tTd4BvlPwX7SVyFFEleNtjhJRXGclWE8ixDnTfIFkXAYGP3CsOrKBjwQ
TUk5BuyedrKGruKfXA5knefVOG3pSKT4CGmArByVZ+ZBjxCFxBPGkJwfnyIMoXKW
lvQ3/s9Y+SFWnSkvJLWNAK28RDA+sSsBTngCtXGMu4zfi0Lm3CwgOpKzcdYzOXxL
+WVdGWSXdU4Bf/M+5RVWhvNSe8fotdQDSSsmK9lxCxFluHxkxnyqOiKKxD6lkjHW
LtEVXv9HtKxyZP+1Ku94fdpCV5aLch5lXu3BP+mvYdLJ0A5fJ2EtF+k/amV08eRr
CUnBPock/1cP5Gfe1ayqhqKsio05++ctq1vk3jDw3K/QpOzI5rBzmatlkS0Yij2v
TmrlUbrfSaNuvGXblOK7tjE4/k1DBlSBWJtLKgVcf2iANge3tKeeCgrWTZRtAA6C
g4fhWEw9JHqDWoskjbMHAWtZvaZs7me7lsnwjJpj7nBWmVuNFG4giwMsUfZPt8vN
qBTgkLFl1lQIhyTQo4XHlCeG1X5+w4s73TfuIJh7jp8qKITmDntOEGoVU7v9Ma4U
ofZR9OoFw7yRUETD23MIOlLiyT84989TmG8gz4Mk1SwyfTzb4KfCAy/ehkF18XCI
GdTliqjiud6IBlBeMMjVbGmCtjjG77NzxAxDWeMxw6oN3lC+yrCA2mEwDqoy379P
nUmVRR3m/thX7Mfc+ucrFPwiVeZzQ/oyLZ/QgYjj7gLAfQx9eNmoMhxkia9PdMOf
jB6LbRn6KLr757i5GYgFMacb8FL36SJ4nSNDI9SWohrS255lBBpRY6zwU63laT4j
46RmnT1FKn1FjqfyhZlDjaC7JKmZceL6Gvz1OKIaMtTj+D7lv5TQ6CuC1J3eLbBR
4G0DANngxO8i8ursEM72be0XVlRqDLlERCHAh84KV8SipPhSHso0ajV9dTuvTQzu
wIIPeR7KWA6uNgEoioql+PEJBgLshvxw56Lm/DbQjgPAr/fcUP2glEhncZDe+24f
FgrWRqGsevU1NOV1XqfKxl5xmIUYsxKosv/1YcyYnX3Zj3UwEqc+hjzuq4ZdGo0m
sh9zWLdwYYdBEPmTQSLbPe9QjScUb4qPEvJyNpRQue2ZTtjcU3mo1fQMZEfLSmUP
/RPVb6MnYlbTvQ4c9aE9E6UEFxHO43VdxCdei6TgKFSzwbhtrLGnKAj6p2s/HiaE
Y4xLSEmLLtAJFucnjyKwPMseorBBGJ5fTJ/cBqQW+Fe68kHQ2YmOQyPtKnzcoJ3I
Gpkt15uZkhp2QK5H/s0SwXOg/xoxfG9nEEsamUHvb37mV4tB/77p1Rt/DvoIVE9y
wDUBr4O2qyWwhq3ui2UmVZe8GCI83O6rH3a0s+ux7p06+tJZMDzy1oV9joj6ce9A
hjggJoQoWigy25cD8lkcbck8eSxo/nq9REGUutY7EhFeoX/FyCnpbiBmRTHbKY2h
c2D4biAHCE5UGQYn5YudAxgQ0yt3dg0qL/VBtKVmoxPmy7eaz8g8/qPgDjg/hfJe
21Sr8Revs7roOjwEn2B77NzsFJ2/gmpLoFGBM0Pa3IwmP1zgSjV9NVJn0sPaXJBO
SBb1OFK/7VpVFY/Q23/V+LN3Y9LeIc5iaMe+1BHNTf3E6sHQf/bXuM0F6zg37XVi
a4mD223bnzplKc5nNYW0sbQJgbcuieUwdopVIoB+Csw2dKirx6CA9VO3jcp1RfQf
/PlFdFXxmV+j5w0fU4KXOh691n2+Zyt3l9unRDs9ufZuMybFIymAZBYv1pLcSzZO
yEemGFLq7nex9x3MFAzrkDChm9xrkUrgLiX8C+XLyjTHPJQbjI133QnWW7jEoosS
Uo7oTViOQ3G5ywr8Q94KtbB/hUUypmsb2vMOF30o8g3Eta0vPm9kL+tkMsi55BUh
nxgh41wQZ6SknEXlLCfSYB6C3QJenRfyYjbUpbaAsUQFJWpnSh4suLbGcoQrsnw9
2rKxnX4edvkeVBiXIxaiqdJvHsQC8wdNj3wnmkwy2P9xfD5L+8JyCW330WL1cg6K
Us6XT0QmpCo8SnWaXRKT+Cl8R6SdbN95SgTbI59Ff6fkWeXdRd7KbE4BmN29Nv5v
bM6hQLgzgOUi/7dhgY07NMlJrz1kslDvUT0lwUtAqT1bXkk2HPwiDjGMnEVnsTtA
wYMeqhzbnQbq/ddjwG3206ym+iC7katHzMfAUjXkd3v/BC600oDGFd42b7c+JZx2
y7TT89dya4zzEhKJZqln8b283wVK2wXV+wDo78xBPdNm+3TZT9trD1cHlqK2oPlb
D3pTg1zRKeOmxBlz2nms38JMUv3xtx02rHQHiF/uMCIDcs5GwuhZbLub3y/Wf/lr
0+IJcqW7XHwM6CpgLOdN6mSFtzCkZ4Y2g1b6nI7qcENxubP+PVQC9rfJQKgkuwD3
+Gs8bb8kA92DBiRwoR3Y4AdQ87eSgSUMklgUIezgR6jjhzr8Fb+dVsfK2O+/zqs6
6i0O9RI+fO5F4po+3d2XoQeGguouq/KOc7/HDifAEnShcf6Dkp+EoHm9/LZ0AUDm
dgvTnRPyYFkGDZApA8dexANujuTS4bLeb3pvW4Tz/ky8k7r+Kympis0fFKgFGUNp
dOHbGHJpVwQOiFWRBq2ozNYL9mJlmNBFaIlCe/qXlwdoWAH5f88MZn2Hlx7SJ3Co
UBeWGCTeKrJfFegJB93wqXsoymZK9NAI0o3+/7cLZcu9CgoXQ3yp4y6SwHEiOnWk
fFHk8ucNWpa2JA0+FfVGZJwGPpZqxTriWAmKQYGjtR0dy9NN6gA/CtTpg415tqii
kQBuTzxzFVIT5VuflSpbg6IzJtsPAtIvrBlXBZ7nk5S/RsAAlqXg41elWTvo9qHX
5/RmMM55OsSfs7v9eEPBKRSMEIgv58In+Wiy2FpH1IgfH5+dZKCJtZqDjSk33NTY
TN3zmg0YkdclPjZ0FoWnJIFMoVY2KGY2/aSZqJ90LJ1V4nzYJnQ8J5gcSEvbgtj7
mi5SblUYGnZE4lGk0cDJxml+nFn5WxFtf++trUyazchfx7/M2Y1ShNauk1mwsdGi
INavd3cTGi4PNYhArgP6NLXsvbc/dJJj5rvUEr+p9Pt4jEoO8hXaRf+ixeI2Sb/b
2iAzLzBVE3o2u84+WHw6W2mFXApR64r8+Ji6yHsxV1blH6hadBCoTC6pLE4zg2FB
LwgoY73o3qiytMwu/TcGs6i8cwkmXtkLPLtHBPPIWsbOkRizfY6ktSwOOdv5l1XC
9HQFggbxi7iMc57mvE4T6q8wEplsbt9OmZXVPyWSMJw3YxC3kP2SUWfm/ElCiY2D
804z9irZD6meyplROE3eB6PRcrhh2j2DYKNXyJ6AhCJhy5bBX5bcmj1nqwdl3QXo
GjYw8vJl/iesOFp1LCxHjUxNH3Ru/t0lSTsk462fjliWDuLB5bm5kPJnVpXGpSSa
2S5mBdix+bmdup1MWttpWfz9vgbCfduCnzo9lYU+pU/RMV766yd7yJgABGRJwvJx
WZdo6h3O7iqdyqpm2hPJyEIf07slLKYwa2lO6+USRFWfMSB0/O+0GZhBdExJv3Be
GDyu8FmU4QHfr3UF6KjTzh3Wm8DCp0n6Nw1/20ofR9cp+5alx/bPXdLoq1Vnsu8K
vGagOiGab79zLrn8EkgTlK9usVJJQnYBvfbC/UzRzV2loXPjVi9TQ4RMIeI1i4jj
cqjcw6zYDXMjvpk+yvkybTvaWyg4EN42DRtOJZga3LPZx4Fm3Vk5/SJilk6N60TZ
8q0nJDPMTgBdl/N47FkwWsxPbbBL8sYQkaue5ievO6yzbjiNuN6M22L8AV6Enz4T
mx5pdmF9AXP6H/zACLo31NsJ75ayojkS9V+R/Ma+W1+zClLGj2hsmXA4SKWl7svT
uz7I5U6+HZg7WKGF0Pbhu95sbs4JAlpgyxq7Zp40Nu2R1iWb27LQ3AHfFEKjQpvP
OLwav4pDE388V/ujNZzbhAyzBG0LrYeNjehrcqO3k1XZDJ0WwtyRImFXR6of66W4
R5IfhswKXxVLxgnaH45fQstTbXjHqg3Q2zIDV/NQ4eTae/UnFM+ebHVrNG6Yvyln
/kDF/OzmdrsY92eZ5Yr/uYXi/HTHq/4RDzxgm8dtYYIDyZ1k5HdH6aBXUbYVEYnM
k6vijzabaZ7HwzdYY3nOX/2P5P78Jn+GBEq8Knklr3KVyxJTIYotucUFSOKjmHCv
bepmoFYjCk+h9g68jqKjsVHIGEN3dv7by0RDQI73uhrCkGBdwXFxqDXMLY51830b
vKaRzdXdeyNjMi8FGSFCr0sH66W5pYVi0cJaSsLbuVSX/LLQb/toXIhmmr5U4BJR
/lKu8E/tpoOU9WjzoJgnnue3AY16L3Nfw0nSUf/2LkL5JtZsoloj2AikIe1HdSHW
j5Uzcsf8ICfi7dc3PXmVSpsBYEoq7aZDHYEIKSKVFTWLMdOFb32zbJyg5i5WgqzG
gpGZhPxcI2kh8Z/m0gG1xUBWjwYSgVheu39FyQWEH6TSPq/M3ckP0/JpEvKZv4tB
uUwsZNXfpqSP576QRp3z2xxLe9E7RfvSSyUxo/v7rqk6jx4ZkHKTiLZaPrLQE4hK
JQ1yXCtULw1400tbmxers98AhprRj9vGZyKEN7Hx6W19jtx/m9lj4PgvnGNmVXbH
iT1TYpXKMySHGzKN2n49uF1mli63ZmYAzX9Un5swMiosfdNa3nW5Eqy8/I2Fb6A3
u/xM5jr+7XsJI9BNNyNTS/vNqNvUp0noYxew6Oq8s9lsqJh/nAQrUCgfoHxFRsdy
La2iR/ajQe9b3Vo/RvVqX9h3JQg4yJ7hm5ZjoITfMdLFpZqMBh83uYmh7Efpymot
hLYIK9Y1JkHc/ZEkkgph+xYHUolqCWHefTr8EpKJNLa8MUTfjGavFjxspjU3hRB4
BB9jdJ/FLhDbpIwzBqvcy2PgVmz0OtntGrtEXkUHnIe3pjr8MW2czSvZwF37olJ9
qY+tDBGsIQOZI0KUKouS+Ohs3V8CIWChX+Idanw7t5PcCAWXJKZ3xhiL3n41UqEX
IC3S5M/1ImsWyPODFguOrxdMmHHB5lMN5n6AvGVdduZI+xRwbA6wHkY2ui8gxfUv
HT9pscguJqN8NaFGVg6eU3zgGl1VY0wv5KisWnTcg+BBqKFtzU73TlcvdP4ejl5D
WE/120pncVQiVp8sstMIgaINIUbnIfiB/cZ9yBrVVdf3tQKR+jx+w9ySk9cF6OZq
H7eUEHkLrONJMBHym7rDUWjkOXpdQ/8p27UCSEESyB99U206Zh9QLo+azg48Cw5K
6Ne45VL/nyQ/mz+0R6Da9Blysf3yVoaNwwOjxZcsOd02ANpxgN3QLxMrn1tkJz+q
EwtCr+Ol7/XV+Ip9x60R2ZA+5eertFiU5IHPcF5GHA9LvxOmCwFqgnTEYicPs5Ep
xxSy5BLVkIqZLDtWGnv9CEexXr6lK5wxSSmIQcHIywnBW4GJBuoFKUax2YEZkSSa
BcYU1kN/W0fUeK2MDQNunYGK/68YEcVLVXfEuSFWYlTSfNQSQBPo4ZH7NKqFXtZ4
yqGZNT9d7VymmEp8vu7PtI2I3ER4qOdMQh0HMd0bokJ5PIVedPIFwph5/ef0Iih/
3g47pHgoIo+RLrTk2D/87wrPq0uoKBTEbwPj6AZTGlilPDgweKFvbiUDIS4G4I8d
tDKEBG2hMaRagErJSE8p9oO2yPBfWeMgMdXbE2kekNdiUa9ZfpAfVjD0ROflPh9W
Zsi6WySkY4D27E+XANJTZGTxjvrok/G1HQ/Hiq/zS0s2uiOjvYJ03cS3o+GHgEn7
1BXQgKtfnZAP/gnbbF+oNuTHdXWG7Hv0IxHBpMrH5bnt4/PCxJVXHhEn3Eerd03i
aosh/XH/m84tfp3k+wNxw3ANTIiAiyVczeUK9tuYLJxoekKCQFd6R2KlOkUg1ILN
s0l27HZhwR5dQbxw8337ExU6sEXz5mRntORci1sjYL98jL/aoS4V2hIgJzMZYBSb
y1BnHD/cKZmJm3nuveEt4/gy9qixZ6R+mt+eZ9crk1ZeG36KAV7KnCJFVNb4pIyY
hrjtCQN0cH7I+lNVNUgqfBwXHSzzUGYtcdywtnMB9I2GrS7B+K7QIqqEMEdxWN/b
KkBb3PB1zUn0hJHGD3Q3V2eo3mIC+smZ1yRW1VIXkJXe8wmskLEznhBtBw0LUs8f
8NxHUrCTIMva95nhYKiKkENtxFul5jyf9V9CEYb82fYN73HN1p7TDExKKZvEoJMN
rEMWe0jYkyhQ1xm4C+WcHoFkLkqSpHbdcOzryoC9uJaDsne9f2hFxe6n3tOf4NsU
k22xy4CQ9f8Oiv13B3UGWuCoyjBjL3ag7Copa2ORaBRWZhW9dczK0fDxQ5hvOWHt
9FD9dlNbc/QOO+m7pYogTyfAAs7ji1ExcgNMQ+wA63jQ9RPb7Mt1CqPTRehtJYNO
ZAP8CO1HNsxjeDHm0fiXST4taRL37AEfgdF0pNHVAJxgb8eAsX/viwrNq2Lk3cq+
hNCK8uLYKnIoeg/IOLMFDZOtypTI5y0LIcBCEsrbCoFMd09/c60m++myabq83eY/
N/7gX+1eNQZYA8/Tu2e503ZZc4159lCX2K6uauH7TZpDTzzfpfSe5CauuHQiTAOK
vvVSiXJqlpa/8aK6DlB7xzJqgnjRms1V2khGSf08Y2WoXr9eLjYmBdYMknnZL/HC
Z68vJuFroAKf8vwOcDrQ2MK14FaD4XOnXqIecU3bM0yh8bHo1eROCWK0vDyV8l/H
NYB9V/SAmhYpRtSkzpRmJKWbNTCx1t90zHpuBl7nKTowJEr2+lCaIYzSqSrrvl8J
nSH1d+Ggf37lCIWZdSXV2coHhkgEEngsEFIUSKG4/MvMv8gbKWWs7NMnrcSv5lTg
Y9dYMBLBcOu5/nHSEffI0eWk5MKzmwMVzw/i7OyqlunENcLYbei133Plu96VNu8G
qKWa+p+gvfwA/YlCh5yr60imNIqBbfCpaJOlleikrUuQw7qSz8rt2oZIFS1PyGQO
MKOfX2W7Lh4Q18DLvd5+oRlnOBXDbslb6thoeBozKG3HPpvI+3m3Obo1ss8MRwjx
gDPW6H/rhy9sUustk/2bSjYp6BGn3FzeJr0HxrVnzYlrfg5Q4jFIre76DO7qs8kv
F0kZDB3O9bQg+earEtoMdb34IkXNHWFN3HKLyVcd6j8SGeA8QJr0YT/iN/4cdYgC
oCW6WWkbyC49EjP+XUoUNIo4etIaKgLCIwsaQJXOx70Xr+xxMohjQgVIf/IzQ5Gf
LEyc/Szwhqz/0GNrwWOblHTu7xwa+Oc6aR7qHNhDcG5GjjSYYAF1pynp3VcbWHSa
bZ/XwbDn3iCLpgEfVglXsFh9vUC6xFg1T51BCS0J1wb+JSh+RC1+Ie6r6+9WGNb9
1HzN7ndqLsFNP9L0+ujIXkPWjcy+YHpJkD6mPOR/rtiSZDyj+ucxf/mojDLnEpAS
jv1hhWAfr67KozJUYDugkKOwCvN1CzGsYyEwWuhHAJToi0UteqWWNza10IPc/BWh
7C8caNHKgV3srmQl1J4kjh6z4DNNZf5c9f+Y+k+0pwdVFQ5bgzWqB+QEdLDOtIDv
ZAHg1PKmTKd5i71vmYR8ilBg6RdNgG+1zpphFIH4mmdXUfAm3oBQSeK1t0GjlOol
zJ9eFFJRNwFmsA5uYhV8/Z97Z/yw+Onu49uOQov5meDxnn2dPPmwHTjdJgJXvC+3
eOrfeAeF7TECqZAVJ4+J08YQnWtgIETJRmv/h7nspgQqYo0H/D+ViYYxCv0r3P4D
xcJCqtECXGgouXQjbrWza13FCkAjjLFJObNsqoHab/uVhLa6duS4ALtJuvKDY5K/
aVAOh+zy3TO1U2deiDzgxlqk9MJFKmegJ/UaDUiu7auRtvqqZZCyIU6Wbs7A4hFL
3tqoaH+8DChQ0AY65ehTq2dk+J3SkrnUY8iK7exjfx4efI9Qjg7GGpE+S7fuX3ua
nF8KH2qy7y3u7hFtvpoqmVtuEHafVWD8rRdQS9imxkgbGX3Pk4qzOL+TrwhZ03hh
sxyt6rw1oi+BLwSpYDHrY0aSpPz9SYBHdjBuInFwMWVWc/G/fvuBJSWOmsuS4VJ7
EbZ9T5jaQNIXu22xzfSayUt9OimqzOHFfNkkQ2Phhmm9K+37QqczM0h/1QhUPOIa
hwmXsOJoyLxsWlSHIuLWI+izpYhW3lx0lV+a7qOfuVOXSsLBHgMIRcASW9o5TaMh
7n0swUG4K4zwYTMti0r7/h9IcY2eAcjPl25KKpD0t6jx2RAaAfCbaBNrWbnoYC88
IcCed3CtbvM3H+XFsXVbo3Z3B8oSGv0a5DCwaTAVEBGYvDpKRWK+nJXIb4zsWeOi
2lhYuoTrebkUC4oZgjqkEYP6UaPZvmwzpd1UD70BwbnxNAuVao3l8ZVdGossZoHB
+hH77SLkri3kJKULJEBd8zEgDEoLpnDsdgfABCFx5LW6E6JPHWWd+aKkVDMWvuj3
zh2TZOlTdQ6keuMUTwJf0RphmOvqJXZbSCIVNnqXPCF2K4efTJSVQPLrTuiIXx08
ufgop4tGt/t5RLb/fDlMH9nQOauqF/1RFQPOc4r7CsgetTtaY1aXSOWXrKz5Z+WC
hYMO/uyg5yag8bz9aFNgGLQrqaq94SxqN6/cjceSc0xcuiBpFBZzZv38AGreBY6K
Z5yIv+zXP29M+j9jFLaD+mMwNLNNbokbbH80H+YwLrQHhYe5SyAupvncviNOnK/7
3jydsE43/nmvPiIAAfrB3Fwk6XZ5q2JDu45EtPyzCtOxeqDBDGkc/6KXGh/1ZkVZ
XMjpIt/AYF9UBg/9Np0gfg+McaDk1FnFuJK42smexLMDvujPnAGW0VjV0GXGPUdd
dgMzGeyWF1VvK63KS5NvO3+UmCixcGw0iLW5rzn2VE5pr8TlrpYv+oRp+8DupNs6
GRLKY2qU7yCoO+z23QtNAVsjcBXNtuT3jwzu/RAufVUe77jO6rJCHTFMIKwHTrcn
ZF9DK1JJ3UpSv4S+kgFROU8ShW6B0wUfzQl+/SOiI4k234SZsJGBYEN1W2HFCSBy
bbd4oibRk8mf/H3EGhRdRCRb+uFHI4AWTfYgJvYnPz4tdaHp+NIvlIQUlgU1FO6n
HxfTGJtYxPF12tKrMKKQdfyHySsFwk2aryA3d+OezNmz4Tfj/CaodxhfFVm52BWJ
nWQfxPxHhKqTI7cXWmgB81xhijvqZawidlMmaY/92corJGyQeKK+DCG2cKXdWa3n
7nJD11vUsGspca7uBtY44JU9oTRVLo2okr4sjYJ12dJDyGJGv+GY4IxAZHKMSXRa
fxtfXZlWNbil52y6LRhouJ7GmmxlHWyqJ2vHTSZwN/4Ev0LdzqHrRpUwZuVX9OAG
2xUuoTeDxW4799JPTynHtZU7MO0IRbG8YsdvdRQrfIgo2VVZ17KgQh1J8za51cxg
O4NNy6+XGKF/UlNRU3jWUqFhMVwEFqSw8UV05sZB7Zxxylb204xhsk3vxS7CWz6Y
YTc69sQQlqzDYYi87FdvAglYz95gVH62p/1+Yq8jW5ag/i+/giuOpn05q6ObxzVD
qkrbIhctM4JdtdEVzREqIo3TbdxZMMCD6Z79iqTSrQPEoL9PdfrapTZNksRwDfcc
YIu4qaV7M8PUtnu4cRMKJJT1jsH6VAagP5HlBUhDU9qviNoxVp7GG3682OganIQ9
Yp5LsTekPfzEeWtvtUhUvMewDPmiG1QlsBq2VATF6Q3XecZ8a4cfrqI6EPCvSYfX
vgxl0SoNaCFKJjqVnkr3TI9sJGkL85a68cFUn2HB2dWkuAvHXMPiP7MjjFclitAX
lW/t/qJRjhbJ2gZMxSouUHNxe6MRW90QvSBGJQ4Feld0pKPi5ufTl+jeNQPltX1o
pRp2XNY5200/8Lwjah8BzsjKpDiBXuecCBBpu1Ts5BHj3nNxH6UWrUWFVGapwg+R
aW6+C0nN29nXtOX4fdY06vuCy0Mh5567CpU1+6hVluCH1LOVnnYJUniK+xGTvrYT
5E8x0icg+N2rsZpViGTzLjSnyC6pfrMJEhmQzytJ9NjxW/oS0itfPFbPM2oKcDtl
xrvzCA84SZRW66xOB46aXvfYRkI8CFXf4tDXts2sxtDZ4cxFjuHpr+vRDoLz0K9H
TRslaJGJND/9f6Nfrnz8p3tg5RW/ZZDzscqTLtnM+y/eXML9O8AJcZ7CAJZvuqE/
12EuGj7fMJUV9du2iQEblYunkaRfdQ4kYpvUNemQlwcyW9l568aB9eBAIVivtBXA
lQPcCWgyfKX8ScqbcMVDURl2Uc0Zc263L3xBoE0o3nLEhGbCOc2+rV0W21tWy17m
DSPZ0DTOPHUyHWzYnMiw5g8SR0vCk8sugn73lB78tLPgqv5lKfOuYROu0E89bZ1C
lB0sJdZy848VI/QbSQyG6/gByxKJdp1v9WaJjU5RH73BUsxSrDXXCzElbgxaPB5h
Pik9rqa/zKmMHgU1Ha1YxBK35UWY7kOfQL/n/X8r2FCU8LEam5UP0nLSPbPFdoqw
904Dah9NrmfyRbDVTtUi/kGNuwMfmzz7NrgSMtauRAZ6uRCEauGkBInI3GaeJJDi
hJ+qUw1CgpVv8WHWSCeAcWS7oM1WnQj8PB4AQSkS4zeIGpYS/4/ON3fB8zB5sofZ
bLJfk7ktog+VpJxpMhpIDgspgM0exh0naRtIxIUpqUyEq3KfaA0mEXa2fZkTFGB4
b5Ypv8jUE1+fEwYowZ2Lk1v4+j/TuC1l1tvmHzmyAYODsiRd3fGnpLSsF8mSeNcn
Zk9/xDyjsEZjpizKqidoujKibElzSTWYDLVDb+9tAafuN0Pp4FuSVGcdIQl71RRp
vVUAjNXQu9GoUFZ28tOf2GaRTIyIl3oCSaE0mFmqd64aF0fksMxxq74WxLss25GJ
zG5DxFib4r1+u501wW52qWYFfuhMYLFu5UtNviA/BtvnI3s1N+JigGZmQSUz/WbL
dhM3w4Fv5qTQQh3/KXglhzLRuezrIhWFFJrgItbStNhs8yZM+7p7qmVhG9rclA6Z
8O3F5kXX2b5qWh/tQGeLr2XDruRWycntpzeD9xrKM4E0XOAlFsReRLd0ailohmEK
D8ftnUPWw6u03L72tU9cy1KsUr/zS5b/v195ddhMSW8hrvkgofD4BlklSjyYoVbz
fKjFenza+FZB1b+rXyVHpxoffUL6sgc1h2oXN/vtX5kxpQiscEo2es6HVkzso6ow
L+KeyJ/NmAsZNv8XY3fC0kXPcIq/QQ0jhawuuReecieNEV5bdEJSCrEMwES1AMMu
NbFY0EAc7iqFc8uoi1mJHwOqsdp2VwhCQkoQzc/C5dhoBKt0YkUgSTcTQE/W2nNU
r8bm/b3HmICD164TEC0OGiQJA9M7N05boUeHUse0CLBfaZ4e04PR/F+KfWMFq++6
mn8ZSsLg2BA1SjSd9BQjfUQu6XpaC1EhAdIwi5zWJNTU6olpCpxWchxGdT+CFGBn
p4ZRYqO9PMtKodfeml5mBpfhPJOepxmR6tXxaiJO51sOIEmnvOFdEvHlQGqsDcHj
MRkJa6bpuhOxUIsubNMK6PJV4HbnHJ1nNtX0PeiAfjhdVdrD9iz7J5/9DciyJBv9
cOKW12mOQXubnSd3fgUPMQRWmZV0QUvT172PVabCh/y2OBu8SF6SBVj2bvJBNRXQ
ZTHbGDFDARQWdJwQKj4fPFISLkmGMBFIvZWWpVWgKslhOenNak7KXSL5IqA/7HNk
87/kte42ERR2tw+z1Z/FkaUtMZShOhNhQiJkDuT0KJB+A7Gq+zFDavUXYL1eRG07
2LHOlpWMomYV+jIFW+pHTqcQErKo2mulS3k70/+k+9J8L2i/XegfsxZBUinBril/
z6M5t++qKL5g08DT8sWbOo4SGEJycD0g5Wem05pJhZ8DE7jbPrgvcYQkm9pkpzRQ
bjUqBWvBaNArOpMOtsGEOPAcc2NUiDqQKcVlkFaeNeBtEVl4cs680yLfMsi4xsIp
673rQv2fCozm0FS2ueC2uR2f7AXcWe+BVpkPsgzLh93SD/R+ClimWUO3b/QdbVYK
OTHWeeN34CVORUI568JRVDkfy7airxXhDaVxZkCmE+MYqbTyiW6u9Ajw7FFy93p8
r2LQZ7HmZqG/Mz7nb7I3np0vP6LlEJg23FLvgLygC8Rc+ucdlEYQxKzQ7y9TrodY
GBl9O+UeTVuVACc9fdMeeTnyQvYkraJkrWGxXVjMk2QiPg88SX7iPVTMLh9FUYh3
JCa1/3EQnsOrQmV4K+RfSfaAf11qbkFR4ckIBUVds9nDWfCWWtL/BbkFzbrxchqO
eyKnxj88jCvRkqXn6v+dSMMw1ADzDARhUFZ96tkqgmXArfsV2+qXUUR004ZcSkBv
yqKcp1PIHp6t8iLdDN7CQKBC9KbNrbFnGErQOpTUCkElp//x2I5pAQffCYsg4nZa
eJU1Y2Ma4ol9p/NiYk4zJGfKJSmwXueExx8Q1br3yr0ra78w99JaooOQrBPE/dkQ
avtCJnvpza8eM0Ijs6GA4jJr2hgGCuqJDmxkEV6FQ++Cn3NnHxCUkmKIqBpnCinz
onvjHuKijcnEoluGUSja9OU5g3oYN2KjdAc0Jni/K0QMxN8LzbsOhs8c6dIpvvOP
pjeBmGCIooDycj4mi/H3lw9fqSFd4Mg8C+dZYaYrVxrk6Te6k46jGx1Kf+yRX2q+
eOhORKC/O6vEVNqRHamGxOhWYly8wXjP33+IrvsuyvOyeiOQKfdcq+EVZdHNrzVf
hdUfEOLtOFzv9djtmuIfXn2xY458DJPNV9qbqE9V1HjkuIWPIPLs8rg4ZiYQSCTs
XdWSQj4Yqkok+Oxm2H3wzHXHvCR6cwAuI+kH4pnxVFNMu+Ct9egEeKhbc3UAY9b7
IiZMN46Oj1AX0Y1x21ad4pexiF1FZq45bdLFxCjkv1aMBhtoiz7h1vR0vC087H2c
Jjv+LEGYsoj94xFdiBVFHl1AxSCS8WJuduDfoTG+Lg6GiZRd91/3gyWzbPd6gJ97
eSTXA9wNEkB/QdTqeCxVKqyRPxyXvk7h/cPc77rMsk40MtMrgvstM1D53H/DxjWf
pu3KFTgxx2dtEPesp4Q4I/FUEmlsa+m28EQ0t1kbh6LXKhv3wRr/7oWhbNMnAfHB
NnzWC0fC11ttV7IYQM28H48xqyw67hLZ+eW3UmzF+46qqE4ojDigYIopW2O7f0hH
3Cn+0vsw8L4m6lem3ic8oElyhwlwESaydNGTq7GXKTZpzWUvS5dD0enGRHJGvDoR
j2PZmPGN8ZR1jmu/XwrsXCZZLHk+dOPpT2YD5oR6p+EujTvRuDEORQwXgFdNroiP
lzC4ruZ+DYhFU3FtJYDIvgmtt9UgzTsfJxtRxoJgtgEfkl1gwh9TPjsmLUqxJdSf
iZ2e6p2DNcjmVuyI9prRzOE2VHmoMq69r6OgTa2UYmTXrbOK+ZkmOcAoQCMqm9gD
rvnH8lA/rEngNSqiXHxyMQsYLvT2hFA9N5CAGePaQdLtZXXpoRCSZUGCqwUv8WIA
49aTqz3LQV+F8orGmLQinAJLkC69+CkTHSTPO3hdHKNbpVHkhRnT/LyoDVNQqZt7
GbbjlTvgHw4KzBb8hfjOQRlMFBRQE4IeHs8kCGppTWWE5yNe4Lfp4YQaH3egTzvN
INi+vU3SfMe9As6bp2+o6Q6ltABZNCXfzHe4PPIN32XHPXykbfNg1E5SYj8/Xl4n
iKzaQQjCaEcm9qnD2uP/U/8VRNrSf16+NG1B/raIfKcwvbucsgGJXIy0lrornGsm
QWlX+mL6qg4gZzh8WEQleQ36O+P7I0+nmcxNj+Kcx+xzqqo7F8mLU1UHD5g7kbLO
OyyeqceSIoN21Xf8XX45PWIX22mYjq/LhzR0a5y/HLVvVYTBNdpw+zDiEkvV9wcb
kohWGWVTzcrOPd5IIHpgNlYDOOmM1cngrtL3u0zSITUtbqlPONzqcyjpX/kB73FJ
2ziKzuw8u8bSCyg+x+lxC2VerplyvqrFLlS6BmOxwbzUH7sJvYZkoE8hu/dgZI0r
q5ERhfiCH7eB+YZ3IbEBVRGrtTc2ZznmWEet6Ct/qYrYKv3oRaMtVQKR2PtQJE9v
sQ4znuFgru1IBHwsGHRl/GEczGBpN/cdimWwZh78M7m2llle1jF/A5nQvsHFOqMI
2xL4/Mk3it8OWtvhPXzLmO6FWKdE8q1lF/3r09ZvqPTdBladBLcoj+k7V/3Wgb1b
MY3SrxIYM9oC4zw+eH/Kg7UvcnVTIAsCtGByWNgtYuN7gfXpsa0RXK1IYVoSQpSO
15uCqYvtjyaA1b+0L2+81ZaIilhFpJ0usBxvS5wo9GrB5KVZHL5/wmkDBHVOW/Og
ZYnZ1rGm3nmby376wjZtU5Un96gV9NWg/IGUQMncsSGIZoUWypK/22Hpf6irUd5N
CPH6xGDu7/lT6DLugGlECyOjqrdppMUYnoGNeO2sVOFO9M3a4OEsFGvl4Vr3Tw6O
TqsVzJwYv7KfTCO+a2NLoZHf3MZh8En94TtKa0OXdxuRZMqX+Z0uL4gLVE+LzgVH
1pVAQ2fuezxgZZa5NVHDczIIUtwY2iqGuR/T1+2gFBSJZsh5Tvdcr8JGm2y1T5f5
K1w4DEFc0G/F7KKBQ/ftfH+AXaxREkNYlwcy9z5KzoD+Bo6dpbOlQcQ/DrbfvV9p
Ajsprc88VXuL+xsO2NZKrifpQOEzJMyZgbqXNr/iBK1cut+g7AFqViyAo4IqM1vt
Fvna47zX61dowWSLghzrMhsOqsRlBRX7REyH+GvuKeRlDx0X+whmKcQfpyHXwUWa
SXUdR8pOWpibrzQkUgcnNPaB5Kpp6UxOOhGExCpHUXD+Ir5MOHFr0+5rq+9uFZr7
ltvze4Azyx0hemt+HBtOpQRUMyKDX9R5+VxxdpIQt0ETkGf/yAQC8Lf+jGtnzKcq
LRhh5FILCkT9bBxnnmosGkMjFi0MyA5Cnghj6XEA0reG6uuybEi8G+QEkIERm909
vqjvLB1a1Uu2gwMbRKUGvCx9vbJ4il5eq5LGTkUYl8QDS3JnuKH0L8paTC8KKqt0
sgKS39XUC2Eg+yFCLDZeOBo05EtaNVVHogYv8Z4Wur9+7vnkFB2dM0x/2oTwa8vs
rIr3WjOazA4ufk1DmuDdjt909DPVnt6Cub2RQskiKPZ81dGnPN1yKs2mOdgkO2fi
adcy69VGacp0dnLA5SqNvLQKeKAVKq8olub2Thj/r6HChA/upum+OF0pJ186DCeM
fCtqYNesFBNiQSiNXrYOCztH4QRLVKzuHdye1o//QPjLGg/8U9OD5MxsxKljtg0g
deiKTjJvQk8ORd6ybZCyY6KyHys3SolR2wcLNE1YPjegS8VmEK/yRT5kpiu2SuBN
CYs8/Mpap/pUv5VDcYohkCdtIQ1hIJFVLQHgqHwOo3esZnp05La4+aCcb1yRGE1/
AxBdSOD6KSKI3dMDu4T4Nym7bz/iwhsoVau9ym0z9UtgkXS+qDF3vlqI7rcdAsYT
dplh/ZbtmD0AY6j9EbiM4mlujcmhxDAVg517MPsQKU+uGJGOQtzPuNDX+4QBMx03
xaXnDsMaT40HLZCpdnK2Y4mIdzJaW6jR7OrPmwKs32hfhL+RLBYMKmQzfrRXeCq2
RX9th945orhwPhoxAiTFXLkCeUnYGEAZfADZHLX2xR5girP99TpJTH6NXi2935th
nEovnqBE0CwBJiV9vNaKge1AltggC0wQBsXAXYgQcKORPvARpivbktMZbVcX1PdD
Ee7bsNmGYLa8Pj2QVEqXonywYbuaNJtf9NJTfpn4o+SogrPBMtQwokitUUkqmrRg
8+giz1LXGGEp3Y4Z6IPkis6QkjrM76fUlHywm/lJ8YJJSEbsM3/roMOWWfr1AAY8
N+a98R/S7dGyFCkcUh6L5bCrWqXBCmkB/sq0d/63F1EfZW4Vk+ky5CnzRzw90yC7
tYbG1YfMGUcEGOdbQzV+nGp2prl6zUaI78V3gyGPxPjWSwGfCZeGIYbeNTkEEOV4
dN5/W4ucXrfFdVbh4lKP38V9HlUuX0HDxDxn13opZyojR4u2W+YDsdbXp9XHDA/I
ShKo8KLnHES0s3xv52CkgTUMwtB77FP8JmO286kaQ9N7q4etr8dV5bG8s13OL00T
a0Klb1tuiPZSgbBVOVXUS77e+9YzvU+N1o+9g9uDS4t7nThIKdo2fnEOHzTMLUZ5
WhVvpYiBKVz7AV6CjM9YkPZ6acLbHcHtgTN1gmWNEyWlsi/q6jiN7+F0JjRZnVyL
np7mjb9UEgAXT3K4aooOP6Djhl73qG4InTE5fWFClQSAPEmEZsTkZrXpNjroQfql
WR7Sj+tqaESohJsJmOXXypAis0h+u1f/NEOHaYJC+Sjh1ZWhFdBdkImzM/rU9ufk
CLIGYdXlCap3jAAjnf58zHdHW7NHz+F4CvTe+qsVGtSCczfDRCNfBET8MwZoWh2g
PSWML5/MJd/ChYj71ams3CvLzbCHAFbQZchTe6ck5ATa67kSEyGYpDHn1P4ltuzu
+YFXf+M4ZukGHTVQg74WBtAKEVzZDfb7rqRHFxfQKcd5Esk1+c0iD49mo3GHppiO
P6ouwlj2CZJHG2vaKNQv8niUc9kVpVEu4jntzcrZh4EhO5ZrGAr+Hlkyn3e9FUkg
q2OQX8MtTPiamkE5DTshLH8Bf+Lcnz9EwTVG/97jbjuv+iGzEWFgHCIW2J5BitDK
oov0t7KFpZcKKKr4bLb0i4FeNYnZBm4CfBNzt7MPSkRxSeSBpWljAkORmYFjeLwF
EM8hDxnotXMl8xdSw0QueVif871ZVYW8hTluFp4UPYZFkhxLKZhAr+xGYEJJeijX
h2eFKWb4ZwBBbVulq+F5T/PuXMJizNucRK1avEuDtMdtqfVJhGZfS3EXID5XWLSs
o5V8U+1QiMNzInVejt2MNVgtchidq4LFMwsnvcP7tkDhA4SS1ayspX3YAomOHPYD
pU1dMIJMX/P0BcibyY0aZnXD+rsz3Z0VxoT0JtwP/P/tAh/UnoVLmDNwFQujh6Dh
npbIgdGB3D1GmQl3NWOg95gehjh6AIGeWxuf1uGSp0EC43/SFHcBgxz6jVCTz4UE
UpdWq0r0cXt+0rgkY+qOVuv/Ttua5u6ujIt4vyqE6LKhNo4vki6eONHsS4XHH71x
VmkiM1t4nb8ML7nI/r2Ew3DkFVUla3z/Rj6i7HTx0zWOSKhAC5vnfdKxvyK1T14y
fj9anynpKCJwMqFpDFVR3gdKsEFgLNmRLa/C5bvXx7TpyC8g+RgVL2GSKeWSG7Si
Rk0GUeIoYmvgmPMsYfVQmorVo0QQB8B0JKPD5uwbsD0cpk7b/UyG9kWbCbYLJpjs
dwpOBL6c/xNx2RKjGKK2S+AhtBEgyLhSCqhIbFTelVuVehY62LmTLxkNI3M5P5gV
hxJMrAx+HAy6mCJ06i4343CtDnDk7rTNPiRgJLbkdHH8CV1HHFfJ5o12MqYSGtrq
fq13OXDm/2sRHnGBmkLNGReD+nfr+fOumu1pxi+9cfqP8PfkAufCB6KRSXnO9Tck
fzQU8qIoW5ymhQSDeqnqigNvVkRwRtJ+mAhyByaHLFaXT998DyheUjDu2rmDOs21
JmGNoWZeWf7+/zxXhJEpXPeMRWqJPLl0kmSxioFAxF4L6nI6EUku+NYBts2q6CY5
WHQFCMz9wlAO7BrDV2Uk+s31I0rtodeD3yCeUVBSNVtOAX2SffXKfgshyfpyBuMz
tFvvxaH5ECdyMHYWujx7PPwJ120cVFlWsy4KlUOwv1Kan+Qd2yff1VrI9o5I39yg
FbCK6zt0OYluC55IH3DQoj1g4Vbomcn8D+erLUZClS2Gon3/vsThBuB+usdyx32r
fVWwJP4Xgf2Ql71NkWIYcy6pXoyv1J1svpoTHZXgpRxL1eOlUD38difqaYoMGo5Q
Y71jNwkAnJmWZxydXnW3HCPqVKl3CL3jyN17javRhm899p6YXZXdMwucLtxkFtVY
377V1WuToB1upsuh3DQJIy5Wgc6qIPNllBCoT+MYH7aZDPuOO5nYQ9KkrL1l48TY
C6zXHugJgO+HrVr1prsnC90tN5/QdHOvKbp14TOJ2SbtxWCug7s/iUx+YyGBkFkl
0JNCnh1mS/XnxEkkD6bGsajQagtYufZX1du+yYyIdjQH1wRi2m/a1d3fVYZk0kpP
lNhuWio14auBJ2wOwCC5mIvghr/f1Y8f+0qSeY1iGPrxlmi9GWrvTUjEQMzb6P07
vSMtvY/AHbgcO0bnB6ZyuvfRJx6NCeulChPwJjHnzLDoUTC3dIerB/jZKv88KZHf
1bdxNcZ+n4z8MMaou8Z5Q3zvuk7K3g9i6jga7kzJOOhxdvaHj2AlmMBkqOg/DtT7
PTGqsoAAw1wJ6X/UhyJd/1ObyW4Gft82yheIAlmvQTAy+3wI+1GCYxTrunOjqMbD
kExYDrIaAMAQGPxFh/bb0SaGWI1/j6PIx2isR5Uwq68IRWAI3uJGm/6M/voy2t1x
YL38gp9RKmBJvIn6tmYRmynKY0mn2oQwmi3jBg3Lyq6YANULdEGFefstoFNI0anm
dIThVlp0Yu5a9Awytq2fFkrBKfAw5yaHDplKBUhLR0/ClY1WR0+VuNsLMWvd+1GT
FWLG6pyxPHTQzFRbG/Gfuqz+3ZXM2IqjtfpB4hwQrecK4o6N+yMOtdX1CzZ4kl3E
KzcY5Hvn1qJPFuPTGzdFOLQWqVEC/nfuEDbyyOgj2ugucD9YpPbYKsVlRVH3rEFY
eK+1dCOaU90FZPM4Pmb7RQe1jtD9hXJ5Xyf/HA7w2d3/Vx3j0mzu04yjq5hc9ZU/
A7yuXqrhLeVCw1xwJRZUs+ryr2MuVdWrMZ7XzoiUJDw6vYGnFO09D+XfGgWbBRxX
CX3KFLZYGqVqwOcHcJSuJC+aezz/caB1i8JPLONaLONJqCDcqRzXKGeRLQiQ7xz7
T2OHngFbqwx54QOPYtEhSQF9rBMhtDY+srpWSdx4olc7At8JvonUlUW3vIIE68YX
0dlqAI0N/r2CwzX5b7V7Wvywe/NiY8WTN/x5RGYl+TeniH8SToWehPvrVvPp8BrR
2b7yZEv12UxN4F9/vcKXAGiAzS74HFUgz929WKyN+DHb86t7vl+DDeStT+QWfSBw
3vthOtv6kmf4bRTz4SfR8nOLhfND56VCIe7W64YORLrde5lIrFwF/vcV4jwzBqme
yg55PhuXFAfdaOS6uSfafO52Wj/FkScpVnjrWNQK/QQpz+Nath+wwwuxeTKgDM0U
jaaTkkHMrBRjZDxFT1DTP1/ur0IaDMhDz+0vySjQa+Mf3HbyG7vquRvwL8vc4h26
axGIQah1izdiUa3AoylrGtnQYojxQ6XfOf1T4BDyAk140f1rXsri0GXF0B3KGgMP
fOw+JCt+vkLr+VkIiFg/59DoZWB2Sd5oiR4HdBExwevkIAYEuKytJB0iAVYFYjI6
vMk1l6mAWxx/V6rmaYkkLTTvbwZHhO1eD5mSk8aM2v9EL0H/QNfBVP443Z7qQMny
N06CWpOlp9cIgxQdLASnGW+mvGreWFq6vp6aZvowcFZHoku6S9Zi/xPa+xVHMhC8
7AUDogpWnOJdlc5Fk70qVPK3Cnc+YBAnWKvypcF19/kIr2JKRAWs/RsERNbkcl0J
YfViI8LwRS6nQRZLx5q7MNQkcRGH+XYg9K1K5XPzEkJLuFz3HsHV0JwT24T79rA1
jgS5pHUzlURgZCyLWcGTKec8iNBGFzdY7rTjwjI3d+5oNtYtyieu1xzOLt0ZNO1f
zLfgDK/lUAmb6ajcJ6dO7gqgdzqiRTCTkMVWuAipORiAHPI2NNy571eC4bVjurH9
wkkPh9k+XsEUMvfS43SCvOFWpZR/nTROz/cHN8ZeNGm3BpIkUaFdubJQcBuKyPFy
8z7G4GpfnpKfGD5jXnHlYpxdrhJoyEwrHyYmqARVRI79K6rlFOA8m9B4k1St+5Sq
i+mejohyVzBlbmFQIAhI2n47JWilpekpa+gU5m+pTR61B+J8FMn8Ww7FNK7opSqY
ryAJgcZJk2qN0vPDa6YgSAX9mf8H6k09XEG34sy7PIcH4G1gvcJzaeqyxNSEr3ll
rjmyUsNpVqBkcC6ltayMZXikox34XO1sw8t1mPaZcZfmRB7uMEEVKyWkZYKeXFtc
TD9EGN5g6NVReZBQBy8pf8fP7XT0PXPXszbF2swtWdopw5le5MRsslYHbHI69/8C
lZ263/hssPS5Yk+cJV6+PW1dr9wKrqkv8LEB0loiXBTNJbfTooe3UZ/flyA1/MEP
Sk0/QPDKRqGG5L2zT3YeNkZaTVbqCBG/XlFtCQog9jcAZV3LWj3UGLyhymGBzWQJ
DHGkqrrfi6SlWBP7yRjLYkeWcf1nmxsd4JrNs6lVcANM/eoYX/scwI5i2pGcHl53
d+p83GkY0olRjNd3LVIdufZv+u3BxDhPJ7zOoYrXJwcZ4hrM9dJtJtTylBxw9TH2
fIUdRWiFKbbWMMnJ0Dl+6GeDFQd8qiLIVFTbSWku+OphyL6F1QkugmmnTp868Cqi
GgsmLap+DegV0hZFAob3Q16N1VQtZkEl+iL5r2gBWA+7Kuq03QzTX2zvcJd3aN/a
tGFdZvibDXkJIXET/BcOOx445lk60bfPjKvpAQpNOhNMfFedXMOuXHdb6/eA0qLU
xgdHOBlgheNTnW7lt1MuViGwFwYOC4Na+gDsgP6j7qdJbhaLJ5RyPo8rza2bXXg1
areSWMlGAF1vo6A72VsHu4t13EKbzKhXmDr6hDFDwKY+S1RKsG4lKuXWbTcwIDlM
wqlfsjZCEM4xNoA8ze6t/1y0TTpCxFLGrN/cSpIFBiVUVdPtvJDBmN5UrNf5iz1P
bkydaByU8tW+Dn8TjyqkbetvpBYgp3UOxhy+ea20cdmF6XDUXA1rkdGJSu15+xWL
ELVaBI/bvXsXprMUE8jI0/okuvSdlUWP91EMszIW6+JTyGcfMWDP1RnxgACsVC79
3DCUI0mBWx8Q7HuS2MZ1vPjhoLNwRdfGMoqjXQXqRYGWCCyaQEizcO3YbXbjU5MT
Thv99ZH1ioq9dpG+wqRrv2Wg4kGknP4RQB5egSRVT8M7iz3cF6YDS8AUJxAheFC3
LcAF+QFIdU6IqBP4ZS/hzspRN7H2lXcKZQwFt6PshyQe+NSbiyzOviOFaxqOe2i5
1P9N0spzoq8OMOf+bytmTbS+vbAPV0kPhdVdT6xFmJKZOSQQH1j7K10J6LlF/yDp
73TnAhGEW0ZU2mu+oqA4pQ2XU4tVt1hj/cAIB0rpj9kCMH9f0JqukhLYAKtERI7L
rNzyzewonDbp59AoRwUysCjJX5M2IavDyUrX1//U2+Oognw7vTdn9tdZqpj7ewO2
xUXHNrMyIMC3U38fCR+vTWRuA3i3RbYIUNVKuHD8LHRAswRdlmYpARfRFhR5JNoG
vHcd2SS8d9n5ck9WDafnM/EbNCd09GO7AirhwLjTAZWb/j8OrxNz34tcxSl1bprm
Ew6zLkdpiEG4CFnW0T+wqKVTzRSqCWKEXNRNatZMeObMTlNkfBIu+NX9ydmw9to3
gjK2b+UbKaJ4nZtQrryMu17amWkohKi521kzGKnj8GMXX8VQw75nmyi6lbNM2NtR
lxvZAZ4iOhKn8WGm/c4dJDHd9pV5bEsXfLAqu1oWZzcRAF9CU5dvr4Md/tpfX4u3
1vJQufuC3JBRjqGuZEeV7Re/eguBR4/y9g+rPvMYW0r9LRw/zFDtucbIVm/pe1oN
sSx0smPfzKyoqxXbw8nciEGXPzPS0O5YnzUIubIhMHARLndoqKGxqLljSijiasU3
uYlgYXXhT7dAu5J2N+cuWoO6DzT/qElSH+LSCuH3ytPO7r4dM9FfFFMax9A4ti/f
TUGhtF60PbpNyDKiJ10vCqqPF46HPcK/U8xZD+1HqQYc55IpxyMDE/u05BAmxUmk
pH2QsFFCkgJ/FmWo8J7LJLrkoxxvGG4S3OO9DSVH4mEugo7TLaP3W+pJHLfH/F9o
bvx0GnHAw/V6vSWXUJajWrPzmKeVLaA8hk0T61FQFMA2MhqulQZ0VRBi0SRuBSAW
JJgLknUTMhtcRzAGv5f7H1QJmGGVz8of73HLuJ91p1v16RnrTr69E/iHufV8JSOD
nmEx9lbIgtN8sVQqRsLpl09sKqoAxYtrUteUOQfoe/yEEIEpZF7X+qXbawildaqQ
z5KxNuWvz7fhIyVlwZBhl/efROH4wSgylUPvnGIK8Qn3AjHQ+NSDoy1as8VWwdYw
tF2dyjx0yy5JykRdhOc4hxqKFGFqID6HCimwyk6ilfw/PbZA4X46pDLYcgPiQBwf
0G9MIY+l30taU5CMYys87JH87FPNLMHZ4sGIMhCrP6mHQxCKyR5Ir/0nStQ79YfA
MMlfkJ6byLbWNxvhkztL2kfTBZR8/vjWnx5AXgAfO/Ok3tsPgbAkhSFMsSRvGCTX
scKcXCiNECZeeIwgl2TykNhHE5PyZz2MQyi3qorlLdM/CwODhFhra9TWAbsDC7do
/L1KV2HDlEzGV5hHZrE2KGxXpCSCWF/LYQURy3I8G9eFrDkoXRmRiWYHdUPNjrhE
BQZx3mqBTkvls32mx9zRQ9Cas9LO8AYpGaXemMk2Wvcdoh3kPSveuinkqvwM6fnT
TiPOQDCM2Ii78BycfT2SndfOleea9NchiwfEas+tT57aQPTXHcyiz2UHSWUARSfA
Hw7C5vzOAEL94MibPXj/K7yO0OwJ+xOVntn3Q85oDEuCx+q1SRPN/vbB+nLbwxz7
ThMTXCU2sVzidgwomu2a9I2Bx75hay6xYgQKStAbvpPZqN4jxifY+Huh9YxsVsFr
TiPKzOXAIhkFQ47+HMvmFiqVvg0N3kZ7SMt5a/NukR0Lh4fsofrT0EtXgdv2hikR
IvLk29CnuX0cNdcLai6wNy6dEGcVSZBrTzzvSFNIrHk5EKKBQdJRbxaT8BgKKkat
H+dESA34zhF2a1no5VZIOrtu751IW5kf6QLwIl/+wl2g+fIokGdSAnEIexruiLLH
DPGu3NehyqrufVv5EEU3/sZSMgsC5e+gxNaxBFisFIdHBrNje7EtYpmOIubRxxpf
sSPWUxHWRzp/r/t33MuT1V1UT4a1Q6tR4z/eDLtorU92Fr4mfxCNSyzVzqYPWMOl
7t0ytmBznCI4YDogttH9ruQTXBelK8T5wh1JB4Y9gv+P7ffJuhAg+JJoj37vEHpp
hRfMNZ0bRwduNWn6qHHuTWS0ohuVcuaCXbeb9CEkRii3g7Gp2bmGEfyxc5y3MQFI
XL9WjEJ+SMjpN3CuMXKcudelaSOn1dpCyQ/EGpmdd1Km/yQgBzOn3wKBME8O88h5
3/G96KBsR4MMdj4pmQ61/7qXkHmWBtRNEafT7yX8KcYcYTcGS2j568x0kb9ylYoN
Bh8CALSA9UC9JxU4/224uk4EhXOwRGOzNkjOCkpv4jSY0WqMuCwKYcxdqubtPZC+
gXQ36amiy4gJtkf9vQaKKru6D1AFwIZU6F75V4H2B39XbiAldmWQXHyhfkAUWBVv
HuGIQnwE1JpeRo5WqgUu0kP+9KEI0ksnKFhJ4ys7JoH7j9xBolmQwklg3Qday6pb
ZpE3H0U5uD4kPBwHV6DfWqTMEd+Gbv1rf/hG7DBdo/ZCvqtyg+0RXXCKKHIHzpnL
WDQwEm9+RwwgPLTko2DF4L7ddVVjZDo96mA8qRmFKUaTELcurh3DE/fuPiEgwLSn
brt6irCiMhCwhD8DBeI7dgeENtHYsaUrVJ1w/TIBVJUE2p7K6WTqt7pMy0gHhzpw
FYs2WvcuE2ApvQHLVpJjMsM/7zhVIHpT7ZhkdnQCsbuLPZ3wsup0uBX9E4IpPV7D
XwGLrCyA1XK/A5vzcP1u4/J4N1KjvX/NXbjfJzMyY0XzEcuIkWd5Csyb5Mhu6ajX
YBqJxrqEQw6+9cNo30mg1ieThSJP+FMV60qP2cyMSxayM9AlVsz+tNturZ9cp+VA
3yN+YYst9IJ65+Wf6DwUlE2ZutV6vl9/Ukigd4Mo5L52ecLnIjJwY4ILEPz8cgU6
hjAuNAYZJF1cnM5wUp/VobLLuS8fHS9h4RMXk0N4FrxjRvBqiio1Iz/9qmW2r8Tl
MfLXco2GoViRI1EC1DS5dV6UGJkPP3QYfZogB2HOaxW3WKD5cJn4H+EvdweDeToP
tnIadiWQMu1U1X+weX9Uq6FRudDhcGC4W3UjIdtLZqqbgRuPeLJ9ZzFYf5se24Cz
3si1wHnaqMhqaWPyHjDp6VxkmrGBLmwhJbA8bPYmyY8yIekqdsJBFdAYqQrT5gmk
yYCxL3VdAXpBDkP5R2znAPgBRIePG9T3FPhR1gJLzvo=
`protect END_PROTECTED
