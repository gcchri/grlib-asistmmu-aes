`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
idFiK2RljX1jOUhMGOAVNQ8jHEt6nRIK2cML7iZMfCG8n8M4gNsE9V0mfoVoZAsj
0yXLGCywcURgU6qNt7RqeCpMx+OZoiHXPfGoc29u1Gi2xjuSz4pCk8Ar3DBuHqQF
XxqpDnP0bRXTmkAZtBvSesvenKAajzFvVFoBujr9YLH22AaBETVxqW6SNfW9+j0G
pileH4LmcYIR/VNgg/HmqH8g6hj4OeCRqK23nRc5uZWjwOdsUK0Kqmg61L1L6eyI
oRJPO4aoYB4kmGZ3ETHJXgzF1xmuvxdgAXWifyoxAYCIpO9gasHt/FH7u/gBtr8q
KqCwQGIDl1ZpWYbFbt13h1Llb9wA6rVgEKKZ3RK1jfS9NY9yKx3L+0/lPzxrQfUJ
4p0mvGI9cVAE47QGNL5pxXiDMC9r8srjd+ArUiC4BBQWTQ4j6acim0gU23VpnNTe
aysr10FG7Mc+ojoIGEjmxKhFil9ucpTgRnVr8+0vopnvXKLDV33/z3x4aWZQDMwi
f1wB4PFNDQLqIH78XD1YGzZ2InTljqU7FdnJ3asgcxetw9TsWCMkNAf5d9cdZwIs
MtJWIRf2sWnZe/XcBPcXHHgAAdXC77lTkkPzVpR5x8IAeHAn5A3Ul18Xassq8rb7
hgR83ryqJ6H2DtY2d6MfCU1Lh5s4mC8s64ZQOADZzIz9iZ0xC+t9loo0Mj/0dGZf
/AhBVVoavEWfu6CVj0Kk0y7TLDgnRxO/VS/cYGAhr7AXKGsn3KBlUrkf13mu9rly
JeWPcCdnMj37gM4wIs4jkTurerecPZsS+aeUSEaSQP+TIkejV73U9IRMqHIvQWvj
lQ7upCWS8WVUKVfoS+6cFVkknHYkE1EJ9WL8UF/Lwt7xh28V55D3SlG3bCC+2A2A
nyGVw+1rQMfTLXnnIeQDW596WbiTiDtJRssdeKf/4y6h64GTGf2vkHecNdWJq7Hq
JxBxMlHcpruqJPn+Blx8L3Uogfk7ib3wdHwdzD+XvGd27fQ0MnfLTXnpQFChUuxC
b/HNjAFKI5Vqmdun/IYD6KWk5I105MKWSb+i6wQd3wBMugmNiyp2YIciZl9xPoe1
HkxztJ4LaK36PyH9UxvOnCqyNFsQ4qVM89eNOqJ0Q8ovRb97EWVr1T8CVACuFd84
z/zLHDSnc3FS5v+H66TBfiVw7yilfR7LqBkjoKXi8oRz7B1OvOGzafApYbwmdpW+
b0I0ko7zG3UOT3heviUmNpnD1NndvPZ3FPuF2+eSHsbYukRvfeKu6g/OZaeaglc+
Gp2FUjUJcQdzVEwZbZP+8BfqqWKk5utAAafyX0YxE+cPdWv2KwsWVZ7sQeQSpJOd
ITfHg1xn+wsK9dEMV8ilzM39NpJkOrk8ZyIErj/ovHcAumai7eR0eXWlTUYtWAyM
AvGHkKyqsUh1pYUy8FF+kpUEN5WXD7M+TkjDjNKw4CKLc+flYuT0ZjVQzHiC1aM1
tCXbXEMwAUgojyD8Cf5Fln2+Qa3bwGaY+91naDyR/Rx4OTb4JihEWP3ADZPTzWer
mEME1+leSEnTl8xyw1toQnEJ6xwquhImu9zGnJavwfXSD5s/m9LU14lAiddnGYR3
aODq4ibSqZzEuF9pr9wduMBOznDKGRBIus9yPayiJBLOkQ2oWUOlOOc8WxI6b4tN
JUmgXt8RMtCpw7g5aXcyRm7tpRLfOOal0Wk8N4KmPxb5d/mG5bqJZJKgy6jve3lb
hOQW92iCSMctbHCBDXvMClHJflIJW0p0+l92RBN2kYaSYaS3hVEfVkcODx8NWRGk
gaVWhG9zd7MbNyRGyjYbousTdC8z9gOpaUKpmub19mLZS3xqsjA7Xoo2WDk6C32S
HOF9IMaQ8DiPv8OR2sqDIdJDFpYewoNsQhFiKKC2OxDS02M3+6bf+X/vEZBwT74B
86QH1LZJ9phdd75pXNPw3wIgvMq3JXerOCShrtOQ+h6K+Ql60qIi730QZJsu6VD9
wry/ZbeT98yiXNmf7aCsJ9JOqc+UPLZcPvGDJ72KR8kDD3oeS+aUfu45XVibce86
ivVwgjl7FLDbOjR0swLFraJKJe2wnHLqEc+r+R57wf9OHe86MoYRoot2kMYzWRsw
LM5g78bDN51qhFBZKPURULZOjV0SvawSJVzysoi9nqA2kCUbPvdmvVePznGSs90R
GwTZgL3z28kxr16ekfBDeDRWfLeV3qDll1GW1COX5L/UGTlI5d/X1f5+gBKrGX5f
S0pu43BvTDgPVOKpxaOKoQUY5XY8tzXnxQcQuzFOD6dByUMb/RwaP3Cq5CJTxQrE
bPtTn17EJXGrF/VvVHnoI+M8DErWGeeXa+fPRGfp1jdJ71RktAsNlvFV2d/JsyJN
gvz98IorPerVHkZQ0+hyi3vJbS23OaTWvbg5vmFmX6GiZWeUN2HJeFjKzQ9gwzV+
z2ja5V5HSkY7I910Zt4784veh7Mv/ORAraDDZ/z+ljOgksN1CQAnhmKIVxSZJJIP
4JcNhKpHaIc5CE1h+GMFNDd8N44z00Rqc+OeBwwHa9b1T3GDuifp9FuuEpj+uKi0
O7pK9oLZkJKhcvHVssx46/PcTlTGWZD/jDqeIByUZRdDc9wXtwfbRLxdC7Kz7dyJ
wNoL4l4IhNMYLW3IXkhZh6xGAR40WHPzrMdxhqE6l1KeOAjsJLSzT71MRwtoqs9X
IlNQ/5bLmZ7P9kOXp75Z5uI7pAlWF6LucLrL0hlCv4eIrkcPZ/o0b/Hxp2rYlZjZ
yzN+xgowviTZJfPO8VLX4oItU2IpPoYszqKy1hVpeCPAppHx3nXcjGG4FxjnjSv5
Rc+GVe2a6kYg0lj7Fkgo859lKSYYpb9Xkx9ppRUPxForrDwac497rSakgxFfUCMy
x0jOAk9O+IStXhq8thWh3/Ug14OTVlrJfV7FK5WZbD6ntPFYWdsarA4eyCD0sgo6
Na9W3eZFQLuqe/LTyH3ZtWWwcNp2ep6C2sap00HMoIR2aGryV5JJ56jXwbqCYG9c
ZRCP1XdgjY1oALVizRv5TbJAuSIaj+4M/M5rX/F1jVR07jxDQkNjImsjtTaVsx0V
NLTDSMhNFxPnkB8wFcryPyD7wnx3EcSbhuMgguNm9cvhA6HUoBmeo0PwpHPDx4ZU
APEp3yAmU/K5DPHHpJwigRXm/bpplh+i4IacyhswjtQQkYdL55eK4o+PLTu1vWkr
hgmC6o9laFZPLHY7fAsK0+A//NVjB2vn1fUBIlfCVjRgTTCLepZeHXbuxtBdgwDk
kQ52sC1wP8y0mlYn67jW2fbfQ1VlM0qkJpI6V16SNvIpInI4BAYGalZrk1rHfTaK
QdItEmILTPlkm7MUCk/1MCpNHpJ2EbRLXPuTx1ZCz13+gZ9+CYqlniVA5PjGOnHZ
ULsg8TdSZqPDupNbeB5oO/v+IRyg91kt7fpcsb5SVoXtKmMleifTNBIHiye3J8nY
B/D3WffnP8LH4jgXVEtNrpKWtjHPgbLU1oNoQZIQHLBgeFk79jaRyjLkZS0WDuGl
tqkhrzAJmnKhAlEdgIPrEa0GUWRDMdx1mSJjNUq+baXU9YnudpahouBJhS097YBn
U4QrsrHPkS6f2tLANy0ZLCIkjs9OEcQKrXI77PCHHfd0tpbyZkvPNOtPSIbussjW
zT0Q63c9SqZ+UIoMwMZ4KxFhAmxg/D06FiTwP2SefQczmf1GLbagl91gVdnpwZso
feb08b5JkjhbPWJ0+rZ3GMEfyxRK9acX8Z5knKnUfzRQgUHVubohPgwA9iDkKEZP
Sft59dosBofMSNinhXEElQn824TGmG36fi9eJYIZjbG0jO3uf9lHIHEMcqKkYc/a
LMqWdXKd5GN62etGhFVtbSY3kel8KPhuBuf+hD6h1tIZ6hRmoFvC06GXCSjG5JeI
Vqd/M/U4cyhmkIL8NgnNClGGQTO8sAHkEJwFklD/suBN9nzdl5A2IqkOryiFNZ21
PsjOLCqZ/jXAKowglEi7XHOqj9x5p/mztTTHi8JAUAF3d4ayQYw0ohEdExmP1kdS
P5b9kY9b4bFL+Zo3q9l6Lysev+NlbRAuknZoPDpKzBlFK1r5XG/t//PmDvXVt8g5
dOr19TnS5n5zE9kiALySZVEGcyPQ2Dx1J0yIkZxjSo4H5u6SVsSKg5VoUd/+F7uq
HUpq1p1lak15w0dBV92qbvs82bL+rBKw12YsnXTz6GiH9bwHO4tLniwq3u2Ue6Wp
oFS6E5LvGvWIr06pLzMVRO2bitQ+wKhGV5td92+uHRHhq9nu+ALwBXQtc/DsCtic
DGIaEiCy08KOpmyxa4iTLF3D6vCTh/3q6w13HX/o840Rjqm60mOu98E6KlibFbBa
Hw33aCkABtiD58/LnboXyykw6unidQARALDOpsd4p9pnMjqEH/Ax1Udrl37xJwwy
FVz8CGFbftwg3wH/itPqiOi6ql3gihd6WnKjOm01h9nSPiZOZOQPnzwZpYWNUdBR
abVKTftmaTQh+HsCT6j8iy4G5pyDy3tXmIKNLteX9yqZkAnjJ6ejxgL1cLorwdV8
zQpj4F3AuHopfhVppjOSF7qR8RI9jOC/vc1T/ZB7pzsHqbzwKS9ln7fstX8dJXrp
3blcwcQ04yBvzkmtLDFKN22xTLFGbG28WPr1+h1be8Z5kpZ7U6vHfkajhI4GGkyz
WX0iJ+unYTh7yKwmAQmVq7kyUaIKmZK8ADr8IYZRKeW19KUPWUs7+t8b9b7xJTpy
+lQGCcd/pHEydwwMSruJ+XTny75KeWTAKdyyyEGhPmEKCBW+ZPiMwaGVpKFTqfht
t85Qm+7iAnKLYL+njvbZqFzOqn9Q7U+gyLyXrBpadt1Vjto6Ezh3M+gvIFE3CWNQ
h921MTcUbCBcXj+p3JymmepTYYCsbPZFQ2/pTUcnQri+cZy+/F/PjZ8XJGpJM71M
DYX7t111LnwgJMGtIZ4SFnuPoPBAESZUT0KyVh6Q2Xdx8qsbZJ6kPk06+zq38969
hAKS9GM8uyA851HUYjRjch7ZVjoE3Mju0KF0UiucOmzP/nrjsveVNiymVDnjtg3k
jUfER0t82MWGKGKOGrJNvDtt6dHgI/w/ad29TqGHykpyaf28RkL0mrdrKJoAbU+q
9ndCBSmcQUrKEHuNu5YT1JR3RxZWCja95efK3Y+Nuq9j8bYu+zCmsZOsA0eFXblY
Y7qCfob0RHYKmoDiFIuEmxfhs1w1kOBodQpASKVIIJgXb8ceJN8VYn80Ux4EJ5d4
M2MdLhaepi6KpnG5DTO1KbhZkslmCA73DJ9J1CvWOrdJitRjNVHtur60MdVThsYT
JHxDQ60rmGw38sxm8N34bNNYW7OdK9m9LD7ZXjSw6IInXPzkuQsVTerolUtuxdNB
PVkTFZgfhyQJ9ILF8T2Q9lkK3r7B2IbuCJeRrOZAIn9dH5Qwy/GhAiRYI862UTHQ
IBkf1Mu4k+7XyJ1zcmI4iGvx8vIUYgVPeIoHMRryaH6Gokx/OnBHiEoFDC1tIOzG
DRuiJlTM8oihjgRWj/Lzf6+FbxMoBxQNi83WpZ1/jM39zi25M9WY7d8fjxaK+rnI
WiO9j7tF+YDUNYwvyE/uq0xClL+ZyI6as+diFU9PaJ6jsw887SHXTPjAtZidKUNm
YmFZKdP71ccSR4ZrfkUovEyoY56fVO+sldClc2SAx5CgHKIa9kZn9RF2u9dmhh3C
iLN8ct411f24jAm4WO06HyELv/PWFwtXeVcsz+pRa4nmhEn/hFgdYgA8rHzLJtDB
RlXvPrBQXUmem03vbBfeE0zon4KbBTSBl1+Nne2I5Krkpn1j7FTkX1qBeJXJ0EGE
Xgkj0+jC1jxFCGAl9XUtmX3KS2DKameRDjo8QH5miOjSVQwdTOC73tU4288aQnMX
2YlDkEUzzdZyWDAZSQq/rRWuveUksdulZ2CMODJs5NwMBop2oyOpJXtqSDDNLiJ0
FvdPyFkDVY/6RfrgakRJH554rw+nAdBJCuSi+znIdZfUKZQvJ1vUyH2IUg+YDRuZ
snxpOfjkYaQ89P/l/nncbs/odGfzzw+TiZ8RGmbRaJZjFhqVP2Q3MXCpDX4ZNn/S
VBrmRFI7MyHHWXaZjw/4Fx5FGzQAvCKOJCYavd22UZNIhWfXweM4UIdi7+KacB+y
8eDnM2DUC9c+1YuXL9FU5vEyKdsIun+98iKzvufdxmPEGrxxsGawtSCaLZe3xRZN
+KNjceZwcd7YdrBQ4pR1juBuqc+MEjWHveE9NQn/r7mLYwz5TjW/HRRmYBYeG8q7
v0hdQum4sfTuOdC+wJOO0xM6xoNN72/8J+f5T3bAch9B8i4TJgK4RQ/s6iYBvC+w
fxfjLDf2dg4X4+LQ6BkIdi/Ctydj0qr2AFGUpgIuwCMzuwulgx8DR+zns0ptRx/G
4wKvi3T4d6aqxo+Xa8SitYs+z3FN4SK5VfbDg4OF6Z6oAKzFm/tHr4VYkRYBfocB
kpLM1w2/DN5jdl0qMdpk2nOGuqWNNpHYqMAA23wXT2leL0i9dbMrYxCtNBAGJyms
+YQTNi/Eju1P0OZfJqzlAfgSeIH7HHXl1jjcwdeiZdmXRyYtGUczt06rj5ThpUtO
r3vZOQlCPuAFR2XpC8fajlEJTysucyjRM7jKaQUCh0Lf1bgi8GdvvCW40zl+otNn
9QKtAmEUANoZZnPiszjxCwjS5CK9Y1yvZhd1tUq2I3xHUHP4ztJNsfg3xEaGg0xC
bQXDHcd60GVlq72J2r0FclTIUvW99tondczKLtqUEgWJLYsj8IAtabKh+M6xna85
lGx2SKbiXM/b51tjGUO5YnOsFeq152nmw5fT2NFkQErfMaUEG9tbFRjtpytrN4Yn
oHcfSj19QKXKsTHPu0cE4bdllTr8xtg92MDPmzuHSwSp/2NpZmAPbLqxHzq6kemg
VCBxYLo/ONWdmCLR9Kv4j9w2s2NLt913Qea/QSypEi/NXLjr8u1mfyLbvJAAyePV
KfCJy6MqqAEMKg+pbZUWZFMq1Zvo0CKAAmwSznBDDq8LjDmoNnzf+9/pYl5ckasi
IalgnMHsFGgEF/AWke+F//PML9Lnv92n7pimkCimrbTfk8QM9fSLmAlu1txc6OuF
TxHJazhk2YJ4XSF+F7P3/KPhEWciVWkkem8zScR4nydO2wFODxhh1tzIxqKEsexR
qU0/tIUHyUPWgdIS7nCXDT7gL7Zw7E3pBKnVZqIIUFrFtcqSlgmckLJvxdYacxTR
LDHKApDf4XQdvqIjrvfF5Ol8WecPfZy5lveXRhupt+BWMFMQOlSxEwmHqV5OqK9J
DBfxAv0tAYdcbxISx80llaL9c5mui6bBULvxQYNu0dT57QFOnbwY6+cXCQOuE5Ik
Ipj0TU16oJ5COw3RWGCBD5rSJvJ+znRYbfT7OZ7PoPIce67ENM2juW55RS/o+y+h
cPCAdojwdszM5XAYb53unYb6YS2muv8RxYdJzbhrnGvBz6tjR7qM9OsDSyMSnJS7
4rcW/ZWDAnjC12/6xXM1lVu4X5VqChu7QRMBxjPpDoKBbEoI7hD7v97flckyIK9Y
rSl6UDMAv9h7369MD36/07887doB3fuoWtejkWvC8swtl1r46gcjiAV7M0y5QA1g
Mply+ov2u3tEzkS/c6IC5OUkWjZz8oi1Y7Qk4qsnSdLGOVjGPKBHBuYvw2notdwI
LIFAnRaCX+nsKE4awfIFG3ULCmCtyJITE5ezL85lr9B2BvWqNcw0lrviF6ZI8QXn
4Gs5KJt2OoBIQYKAiA0gieSUWsVEKcoi/oXWscbgecWyhJcXppPWCZMGrySniW1T
m/ggIntMVS68bUR3k+rmcpH/lpvcdhtgSdhBfqzHAtDRYHeEhiUxKzuqAV9ojfRg
YInOZlh0M0lM7pOEAXkC5nr8vuIkUrV7iljkt7SxVDY5+wKJ4DdMwo10sWddA0aH
+F8vQZJlC/ZAn2Q9t/PZdhsP4T5CcTJOmrYOosommi6yGWdl4IefGmhgI63kPqmd
q5RQhvyDVkf5Kvk/YcsH6/9qjCsR8jxP7vy8v3G8Yfqrf+TTsdnIzpulZPvabySV
nMD9JWnXQU2L4g6NQBZLgRZc+mkZiynHO6KU4v3/qKtwZdUe+Sv3EGPS1lniQL4F
VshMihLPnzFwW8IQxl3J2/lbFd9HhHVSStIzG6Vh+zqbs8NVmQGfkVM3+vAo/5vG
RKjGmX3w8yNE21NcEoXmVpH3UKnRyMV2q8SE2I2ExQRJZpiA/ACL8RFegg84OnhB
2ovFk/gJFEMm+zHK2QEBhVWeJw2lHfmdVq5p5KvoRTt5UlT9sxzBs404D/GHzHK+
DnV4pIfK2VQG6xK1q32s+EBS0dgRLqswzEgIPQOPp7yXbjLZLQocoup/ydEDtrc2
dXtbrCr8vjB56zuriAw/+gNIlAFwDRhhkV5WPHoetU/v0yz5bFhOGtr7o4+qlHSn
Uig4NEtTOnKDVQU7IQdQQhLkQ6jyhUmGxVvnBm3SiBsug8xLN/WZTSdacYonL0Eb
901BScfPC3+yeaVr9Ao7+SajmHt1IvEkiWN5ywi71WQ+8dG2Lea0yjStTJOgs870
hLpp+eK2xS8oLmCYlpzDzDXrNIMDnCP2szbVb937XNlrCsqsgq1u8oGhW7ITvC2V
C6g/eIdQH/H0sJ/Lp3AXvTmW6Qnow8pM/re6sQJQS6gT7flvsTLtSf32W0PVK+rr
MPS2j/JoBKfAlCOZu+Asvv5pBsiQplwADjl/hoOTbIeXZ2pCNj/JaPOWivkXDtAB
/9Gi8sYM3WP/WHgPa8tnjBLdME5BaR7qwCgOOxotzeIPWZhR++zmwTjqXqrUNVpA
SPtLIGcFNTZslgGYo5ySI1UdZLkvXhonb74HvPcxcWr4FFZbj8s+z70YLmoz0JXi
62FHYfT1dploGwKNVIajA2KGjhnT8CZucezh1M5QdO1ZNoODyglXYDV8I50z9Lkd
aAe613+y0guyxZU4CLodkFFD1n2TQBjW/0gAFvpnAGZ/LdPjYbsTNYq7i3uuoKVU
MGfyWdr/Vb92DNRO6aeojqsfJ76q64t6gRf6hC72jHAeXPcdyCXmcHQzXUTpyRrT
HPfEpg0yApuhuZnUcP2sO6N9bJPe62193uFu6is065xEeQJD2Jqtt1VluFpisS+f
s/PEmg6wPlAjQTnBJc18P/9/ipC90dWWJ2D7SeGk0hbKKnJejBBVlX+iW1Hf74+w
G66Kk4Ygay9MSoxiv+a03zgK69zzPjDhBaKmiOeZ4J+PV9sAxl0VjPzNAOrhdRnL
BXlzjR4XkfpBOyodfW4qnpEKz5ABoE91FtPkA1Bl/Mo3wxPp/H4Y2KqPaMr5+x9c
tzwJwVFO+5Q/QMaa/JC40hHaiwrkrcnYWiKIud2lmN3+GgNn8z4pmmK0uItLHUkD
3dwWyM+51Sl1T7wMZGebO3MKunaYUtWhVg5EcpdVfPi4h/NU0d6Em1MFbfqXnQ+I
OusDftYljfeEbdrKAxS+twfY6io9s0GCRihC/QUwIaYkAWFig1x79DeUbn29J3DB
1hWff5Pjt3VqBO5H6ZaTKE2M50QMIYRfb4EqoORnZN/+AIIT+qlYkaBR9Fvgi1pE
e5234bcsDIHJ7vZY6E4xAvp1foo4bplPVUv5yGt4UTddD4OCOq3FMSVGVLJPH95v
jGvBuQa657f2qgwHf21SwVd6YWspjw7WbE3cwMCMM8t/FCxEtwSM0lJeLdgcXVYP
b+DsPLdiH4b1Xk+HKLpbvVgO88BWAko8r0IMEVaQc5fH0dvW39mHwHyt4NqA87rT
Key7SkCUuwY67Isie8tyqPedY3RH2Rt9wtsjQ3gcg33M0M1XjvaSDMejZX/GGPAe
Hg1EuezrP+TV187c2Izk53ZKPgddDTL6UvmQ1zBSqpYA+yaitC83OAS4mpT23FWE
9PSzxFg+7I9a1AIW6eVKsZfZaLE24YMVYYW3ryI3eQXChVlEjlVBrqIsuhzwiMb2
Xx5/YVrlZfn/obI91imRxWTMrHdMtm/UTBHzVfTPvB2C2m8plh/9rkcqL7WT5F1a
njXdNnDoG30MaTClgb7eBcPvKD5G3a/7Y7fSzuW9BzGpggnYtQFEEvyCSsd+IXKP
Zz4dV3VqgdI7WPMtISkmry4XrmDh2i7o5xwNw/uYONvfRI52JNu991R0vB+fH9cS
gQxqOAsGaU+QzGH8gr76EKDhL8WFVeIEDk2y++VnMvOJ8RCm1q57x3JkjgV+pcng
pJbE/VZol3jTUFSTnOAQj8h5uU/nJ5/DNDmUQ6Tec04LYE9SdpjI7zu/fUM/PrxE
ScAnQBwMvWsNf8Vq6JpwzpgYtD20r08dXW9TfHP+bR4ff/zHjVlw9yUY+fPHn2wb
TeztCxr6D9sQma6bi7QA4VGJJat03USi5qMTcpaMmbt+2+zRiSPgJRDIzkqgxqFR
7REYbtTm+UDML6m1FAFQn2AEtwMkFkvq5pfUDpc9I51Y7ahYJXU6Eno4hJvBPhaa
EXc2ZYdO++RFNuKQRiZXDjqIPVM+jfXl0jVAV6kybFtlz/xRktnctTp67ko3oTX8
NDOgu4J0aKHcaB/LC3LV7zvcrYABasyrGXPJrRuheuqngQf9HqaEQs7GxdF6HRx6
fsgLTMHvfSpdpSpKOYeA+XBeqQF31UFOOVf1P+goa58+qQZlr+dsCX1fMPTR/va6
VQAz0ALJZv0HnXIbKX5WYCycRylNQ9aLKGHsoTyrebeYtyr/P/u0TsKQwEZbaDj8
0fWM/wwdCiT0Ae1+9cOlye3YsWo9/n5P7Da0rnHMiOTCpoI/uObVrZl70e1VWYoi
LjuxMeJvqIVf64Ww362doRGinCXunXgHUY3LvV4ndhgoj5cnh19Hsy1ZR5uoL2JJ
PKR19hVuuXsiHJp2oyDnVaTs8+2QivXbeHACp+O1MM6qRMAsiolxBt456qTRHj4I
1Sbel6bI7DLIupWsDK1m5pv9jTXTbYQT6+lZCvVJArmPHLB3zxMwvscXQSQTNVSp
wzVxJ25eyx8kV7ndYiRoXtlNGzS40aqmoDKVulJQt9t3e633UVX0t2vnTGP+QbpL
B+2F5pUdB4OfU0tlBiVriqsD0R8TgINfVSzTWcBG1Lz8WUewaaiJmSly+j92gjRJ
ngVag8nifiDVyY6zrvpuiq+ST4ALU73bEp4LXNvILnUzxgy4S/Tvh6QkfZ9bbkGO
u4uUChTYh//1pNmTTIBXXldKNYRiDehhVqED9tOWn7+QwTs6QGMOtWS9iVFvx2gi
t3vTVg/9BiCL+OwAIL+mLuW+geduH/uGvml3wjlQorfXGkpSMTIUELzTDj4ce02n
FiWuouFFjWREQ5WC0e1PN5WxyisieoURrIb0ovNkcUsNdh34etYdSUtuE0DOG3sZ
tEJuCVsWhfF9zVYHLsWJ+YnGQXGVIC9iERz/pV8NRpr1Eif0AYqm6UPpHzBD2qDT
iohKsJBn39DllAN6M14GeG+9yB4e25+e+3IzjJo71nsQ1TMH1/gmGQo7uRtCwIEG
LY49gPJkdEc4yIQ06AFcn+lgSTZL+UbPK6ZXNceZgtg+7T0Z+LLenP84jHrRrg3I
FFOBCt+2LouVbLplDKDVSiSEcUfpT95W22ghe7T2zrbhnwPRl7YZQGopC0QLJG5+
fSQ10gi0VVz4ViUHAeXFIO9qu520ZtA3Lg0xsHtxc59WJkPx+xQB8qxlX1I97O7h
48FoISmG4Ms+Em0DDeQH4ixoJfzQGqjNBvkd5TQnag62T2zT5rJ46uF3FLhFNVL6
ryy6F/07lKc9nDBA4NrcRVqn6lB3ItSaQseoMTPDJgVxA3EE0l9zc8K0CTifbgf4
zusyHRrtezy6Ku67ETYP4tnbxuuGEK/9gORRXMuTjK3bMpULP8qERpDIyaMHbHzl
Q/NpyCOqNE+TeK9MxEn7SOVc22SxNZaRg5Gz6whhNVTKotWxNebYzGq07FeK74EA
8GNs9DmKn+jnceN9KuAcHMpyNaKpZx+Z55kfoHlljVCL+IC6ZX9/8FoydDgycwlx
XamcoKNDDKctG93GF2NwA9lPri+ndVaK0XcMLSl3O5sqJUPLhgcbzS+y5NhkGGKb
Ig7i0dpb5UixWd9+7aCmZR5LXaHA/4tMXZaSPCrbPg1MJgdbDEXVCZLuxG29yzK5
FZT/0kr7SArz/gIETZbwzyJoPQL7mmTsfAJZC1o6yoEy9fymlMN52/Tdsm7sVQbJ
snEkXuJ9sHlf6lWqadz8MXKwGJRKgQnO+G3iE6VZhKi27j+xjNKlJzQRayfIg0GU
VGcsuqf5s4Cw9+DwQ+uDAEr60Jxi3tnh1w/roXec08S4HU6Vgg/upW8Q6rduWSwd
KYrEZ8xDy7aO//JwulWGg0Ra22Zz0V9r7Ba14Lsw4CCHw0xFY2vxFmrgEBhq2FdU
x1SPzTf/PbG5GBamXNJ22RfXhh7UJmZdZFvJ2gQ38/E8mZup9p615gVl0KkOKMie
Ldy4HUzbDY1rOII2EK11qGdC/9ngnWgywWGuK4UpVUmENTgApeEzvNjMYcmE/8aS
rpx7CKj7N7WnzdJmsq4W3aeYz5dgyA+yqP7B17YzfLAD5uAJZgdbBinvT3Ia4+IH
uTvKSjIxtYt54zoLTaQL4czjDlWRbbb4yPF3oNza5s7Bvci6xb4mR+qSMY3AbNLP
zoqif5luVgehSwPdE2B4gmmLuI/Wy9nP0geD9ntCT8ff/ZAVlhpUyMOHHpjNwywM
RJ3wNnDa6sCShggv9byLS6iBHeVjMFrN8a25Qd8JfucDJNfWMud6QnTZSLK6GR1j
u1g0YBH3KbO4kvITz3vBFdaT3vuK3qbpnKxSCAqeSdnFA4wjZEpPPeq7MRpDBwg3
I09yAtE8SRsbdeisa7wZqccA7Qzmq9NB0LOLB77TXsE/KiNb53Z0AtQuKViYiV/t
/hrFprrBAclnNsX9HS/02YEuxEUJOTj+U1cK8QXHyr7Ery2agNQFigl0olrFTLm1
hfAJUo+vb2b1VfqokHaOg6CjkQtQEfrLbgT+Bjphiy5YnY6L0ooLCxhS1LWqCXlf
52j4MVq+ArZ4uwy1oghpVm60TXrGV18HPHs2T8n/nOQqnEomfb5jszKBnm5VYuAp
tkXGMaVHvK1XhHAGxya37B8l0sFJlxJOQ5p2Zqma3x09b6Oraz/f+YSUxbXv1cIK
eBJ2RxyJ1HRoy7cb3awguyFOLBr90fBCgL82lyAypXJ1ajgcSuK5tRpR+XHz68MY
11ywupWzw//EWlxXnQvKNsYK2jBfJ08zKkVWl+QBswv0vrPu7k+z5PUIyVryx575
WFEUxSk7hn+Trd8EqpSVO/NEJiw7zSk5A/Hcq8g3T0j2wv2pN3eMGCuSyxhY2ZKk
2FSHCMnT4L7RjzsxA7CDd0NwBCoaQaig6QpdBiMqlt7Ak391u4SWqFTK8640NW3o
7pivxkoms4aKIydHagnVVNyS1R7OqNocNgzzDmxNcA3X7tELvEz5VRqMB6YybD7A
FreQkSWLCTS3uYtU4vJmEprs3MkEev0UWqwJ6sZNa2WH37A3fUXJGAAotApz85Z9
+7OluJkOaOaZ9pT5ziGXmYZy8uoIGr+KjQ4T9rnMFT/qVxZ5QluiiCvxMGOsOxza
bvxM03usGcQRoS18dLGx3zTFgsAyQzcGQvNFnHRh2ug0pS4Axyr4oSzM3qSqdfLp
8106AjC9EqgCfEabNfqmr+cyt0u/vvHbdKHmUgjS6KVEuWBSgVNf0SV7fwt8RImu
MD+YhGOxO7YHxR/SrXt+PlYdR2HiK4G3s28RntflqVboKlsiZRX9cMd8o6jVpMbr
g11lTxl2hoENH2MFNxnknsi/wY2LB6ZPYBXSDAof5tuV01gMch7MzWX7yaNzYmmp
BVSrP1EvCaFEEO4ki5T1qP4RIZ8r5WEcE2Fb1pXZXqxKvSSRk045uMBeIdVlonGd
IKVsN/hzqxz1nMFmLX7cyMAkmfALUI+A9rnTozxNkTYH8k6ZQUYFGIuKEDQUxMhX
YQjeixTeMrfEaywiEhMim2+cgt4LMBDCIfTIqmoAropgRs4cyPMcgdVKbKeTkRtW
AcGk9wVvhOG014xkF4dJbHiozTAZH0kOETNL0RazP64WB3Xc2E4/9pxaWRkBorL/
bgJPk6vSUYeJg8Ox5M2iv34sE8vAH4BaZ/Azh93b1S1crxWpCAnmnMc0WIJ5rtuA
oUeE+Q+m/xRHX+zWcxynvt7zTcTjqAzVYiYPN6fBRHtYqbJRiselh2s+2znFX+h3
AdbSf3zDqZUzAGK4UHJfh3oUtVBwyLVks0rs/lpy3v+tIeuU34MHdUzU3iDNoJrg
TXiUFTZBtFkhFlx5LsYTZvNhJvdRJebrMegIxHuM9/duACuTXB3rR9VH9+vIaBqV
gAHzt65LGbagC4FiMQIMGLoKEuK4JxYuSWmjAuILdtp9zg+MnDJTtAQWOX+11jp9
uwQxTfqWc1gHYYw+jpCVo0rh2n11P0zV2XTOT+ESR6ueGBO2AsD8zJyEUB66Y/ep
6mVoOo050QN+44YW24zf9Qmqe8Z1yF0zbdyWAbAz6uprvj1ddDgDMgGDB2SQrYlO
NBnbA7+7hIe2nJ0QBjAMhdSS8F5IyuEl8nFQyZs+/sXxzAjp/gQdJDZ31wNliHNU
H2MsN2IVpFDwyrfsynSXQHddz/5zzZsZ6y0Jo96geZMapYttCGFnbWee6Tu/8QrG
JK2R5vlNoKsIc7SWc05z3xAW1DqlEWWPLuC5m7M8OxGosUGOG8Puw3em8u6FfN/g
xU2NmFs2mI5LXDTKdpn/YSR6RPR9Rv0OQbp4e41xHLZYeUYo64iEZgPY7hoZ8s8G
nDrff3isFhaWeRmQk2gJj6paYdGblWoDZ1Mg0iT+dMpUoeBrd3drsM9sDy37UzX4
Ky+OZbJUjZWHHEXJAdfROqkIWUn88wn8Xvwu6lHr0XT/GBwS0wv5LF4aH/qv4hnW
F69gY0Dh05vPJ+/JpUrI4mb4u2wTjcmhBhc4Ibua8yhfunJNOowKigfb2EMqwNPx
LR1c5vV/v86GK6qvULE+Fe8/uQM/lRb7WtS/FA56B93peaesBdlw5MLS90M7xlpo
fIC8uMYPzYHO1IeCXUbnJXvfdn/3kLvf77hREPYyPfR+M3AGH7yV50AlfIhGK5ml
kTkPbyijydds+96dh6296eIi2BtF9Xw3VDfPjnQR7LMGqQGnF+XIYIckllt7v9wT
00HcYL69YP1D8c0L0dmM2DoluquHtD86lxqJ9TV9flxgLb9r9n9lvVLrDuFbloGs
kQmS0HqUfofPPbt3kFLSaBp1eUSNBwJ183hFH62Gs8kS74381A+drhEwd4+3ZQY3
zPSFhTibBId9AEnbxdjOLL9L22rshMk2zI2XV/vilNZ7abINC1b+/OXKU8RDLHMY
sYyQQ5385TjdtwGcnGNsIn/X41ogI3w+W7YtgY7NWwkOapys3MNWcbov2Q/9Isfe
zQBf5PXXFVE2YjvjbBgawuNkpBuGrdHKl7r/IMFrLLHA6DofJOQpQUAL3MDHoPBL
N7Yprkb226RJXjVQVsVx0scFvvd2kz6+dlbxNNvSDBkYzQ8TGsu5EIRyrD/FsFuM
0n7QRFUgIb9yuUUb8/dG02YYtb1GSGVz8vfw2Yn/ADJ3gG3vaWq8cF48dxTPP9A3
TXUQzMMtdGeT7d1hBzbxfA9+lvRoZ01gw+i7soWxdF+6GBOHs8r5QesW9ODNMVmN
bNUa0w0aR4lAR3CaU+Tf1wbCQ5XeTvp4EdVLqMRgFFRWsxRgn9mTpLsU1etV/M76
kWuHzBmcPEq1ZkM2ZgUaPYu6wxfLbClWLXdzr3KmBHeiBeQjJLCO9T+7ecblyhbD
IfHIKQ86rE0nk/pgre1389Sznwh/8OUrG3gfuucnumkKsa123wxJ0QDbaxjAbb/Q
m12ZVTB0RLdmTc7yZ2jCgD9QO8tGZP8Fe4MRZ8DP/zmFUM4oAdFdj95lch/tMGjN
l1sYfEn7EEgnbRuIAKXSFQGiyWjHgzekrt67cNLBfOshEFzDD0DJUo+UUb9S75AQ
tpaOXUFN8UZzeEOltyNkKF5iSLrCgb7FY7G1zxI4SVMZwmArcEFAGyy36XolvnTx
YcFiBetY8ueVi6kpV2t19T4AtfVzzKCMYw5c/fxvSjgguPA5CI2trLTWX+vNxSCg
EXH7jjr0jWhPwrVzxhibTEXnRpScU7vlh2V75N1CpIIe5nrok6m1ugef5tuARxqK
kFNmBSpyZXd+nthGfoYahtC13xKRd4R85e5IsA1accecoLa9hnFdVnBLldm8XurW
rpa1DkCnljkymCohxnsGIhVTHXXykB7szJ/PdFkqjBuhujcC60Wa/IjTVzTL29p5
kKqra97pc6BZYOAbt5hzMd74p5tPcoX+yKsr7yN9KEwJNhH9ccH7eE+Z13ablkfI
GiTfFrx2tUs1etn/pc4QGd25sRcEyJB1AJp1qtu/dszwdKD//EsARPMPW18eAcSG
b5SiWK9lq45PmURop3V2/Vk7TgTzjCp9nV7qhmNGNUoJbbV02hXZHeI5z1U9VzGG
bCqc7oSrqi4JmcdNmGQkY/4OpdmvGqAJlpXi9hzuB9NMItUL+wVgBWykyKSY2n9k
Y2rB1YnacQwMc9DOUcaysCHeKdUhOz8PstTZ2P4yPgoWC6JtET0J62S1d/85b8Ss
brfdFO5LiYHdzUyQEEGsInM7ew7leztOMLqv6W8da0wc0PRDSw+7U/UVU5qB2njy
p4Vz/Yt9enf3M3Bd7oLLN29woT6WCIgk8p+05K0LzSf0iVyFnejoxFHBXnxKrM9j
rLuWK6y5K/RyKKXz+HY8S0ehUYi4azVDSLHaFjjrJpOjahgCT4dg0a01MyH/GtMB
N6LKWBldrzVyBowAd+xwZzUc9R2tHHR+WUqtrv6zISDTYjRDScCkCuj/vu7x7O8C
yy7o4pYfEQxvjQETAoYI1xq9NUISP0XcllyklagkE3XKw25yS6iBXM3B8muBdx+c
FYJUReO9q2GLA9lN3uunbGOM0BcdSAIA+6mrcA4JCFAKArm+IInzSL5oUfE/e0Rx
voPzgJpSqN86peUJwtyN/86ZBzkAVp53nPPxli6It8TdRGjLX6wWL2A7OWaxCHRR
R4iqvd6m5bPSi2g+modflTx8q36CXXLTAxKBMD4jzlKRZucRZHkOrgSOi39OZcRL
1COVAH7hmdvnrr1xURd4o0lplw8aeu9Bl9gI+1VHudG/CvTTdtdF36UjScd1eY19
Gnltw5/5tnBiq6BJRG8SPLNkL4R4/tle2eMEkmgubMB6Mgh6d9NbDT8pr4DSw7dT
6g0NUgQLrFPKSUEOgwtxRf02vPOMLGz9kiMKcbGfhZSOu1UUcWfAJ6H9BIRzXHjh
adF/XQ0seYK5nHXtbEimlewC/HI/76oIowBv2QrNiwEJTh1rvIsqWs6XWykJ68Up
gLhUTOjkFRXQ2K4CC9lLTLApdkG0X/rTJqePLaWK9Wi5DdbD5CN1UCDLClOsskVt
UtoNeLdbg3ZYs24IwS7qWgnSKpu3nCwRTNhQZSuF8tXv0Qa4bmYXLAfpFplTIwHD
oZUrNpkGHIP2T1QAU1EZQ7Quxq2OjJy7X3UzOgNXoeSdd1pQwFO+aGCh932eoHai
N5NvW+PqOyVM+DB+LhLc+42aMwT/pUABZhTyh9uAIY7yy2aywGZ84B7TCrHzdruY
1Rijp49XjYij8M/OUw7XnqSg9qkgHQGrwEvGTi6U5G73LHgHxj7NpmNsgJ7CGLqQ
RU52Pp8HXnVddwfcJ+0xue5j9uwDz1aOAqH674akuc3Fpmdbx9JZnl28pDc1lR63
UqsHU9EDiKUKMict5GdJcfTYpz/VQbSguOMsxCc1L+SzRTCgzluMWmEwtP84lk0H
+td62elPQ301XFtc52Ksc/2nv68azSxtYOAyAhL3HAci3jV5MxX5ROeRirE01xKW
0B3/7nB7TAkLaGNSOlBDHgU+VQIlm7w9VjKOeJuzzecE1N5CQNPZt1d85ri0PlvC
C7gCDCmme7ebHh884o+bJlfvHbppvpU50aPgr7HDQQJAG31PPyQCIfr5c6LdCLhN
Fr7ri1zi1s8Z1eQg44D8T7eN/D+pa2KOzKnsqrgTRn/CfVBQdpPVtZh0hdJJtGDS
wHHvB47bngeCLJSDA/ywcMnMsILsu9aPUiB9El35TmAc24L8ijZVuuNbYl3shblF
AaOnNt4F6LZs5vE3gO1kRPHEQ/LsE3gqRtfdjMviFM0IRPZ+paWMM/RF3L+6JQXZ
Ad7iobXcckVXEmBltmUMqyEkKwDH/YmC/CONMZK7lciXk8WUKvopJtK8CKCCE51P
Fnv/DZso/OvBM+6ydIdLy2s6EBFGCTDJm0J1ijI78ZbtuwjqGkhJsbzu05vCGYLS
vbj8NUsV/gpTnVS9QwulYLFScaGYZ9GaGTU80Rte9WFCKHSW1j9mI6qaZXiGK025
1aoeHqTKJhy41F7i9OizpUySX81jgO+3OgFhyNkMn8D7+VO/tMyNzulXQ4Qy9iG9
/MQqoWaUtIEB+DeaFoC8Lg5Z+U+u43aAQIGpBj7wHKYpbDHnRlwq08RFdFuAe5HY
Qs/StciqkkJvswST+BKcavFU6+Y10eW+WoLBybo42JrTDCF1iHqO7DnVrJ1oUDc9
RfV3yP3r8xxdkg9iQVoV00+VFKnbT7XuXUDWKe3aGJdk2udw/tvMq4shIQpoUb7o
pjSve0fE1x6skopRgrOSymsGL11eZ67wrWX5nZ4siMXqLHdFzFt/+7VjaB1/wAt1
cH+LZZi9YTQyvEsjpskmD+7ZHwRnZUs5zd+gW4Pa5J9N4Zjx29/BGWXu1b0cSy3Q
qiRM0vLhvneOpT9q5YZUHpg7noRM8do5zBpW7ES+pRhrK6AjrE039SFykqTPJKKk
hAAnpMUq/zhrjmmrgyrQNNncqLWnCQ0Tpn8Zbawq74OdSgr9PDt1sVBAnbp/HFSP
mBh5d9Q5j38BE5A7ZR1Kj/+cGQXhZ4+B2U6HGGc+Iga9ITIVqZ8C7HLx1e7t6BE8
+PnrTTPlFEiPTk1II5S6v+pasA+DBQCjXc3V0jvjBZoajx9HrVWnpIPex5zm4LgC
HUnTjgsI5sONaxj7pKNlMl9NEeXMv4SbOGCt2dJIURaFUdTTSgJvMouz3el5peVT
pne7hRfVmkbsbOsOjEoRLz48Ca5qy7hbI3Q2kigV56/dyKYRVMXeUuRehkY7aopS
/1OZtf5rvWXAfDqlkgfoWBhDGkSAsUvSdwB1f35m4vsQ1LlREeASfIGy2wN+VBdN
cVCCA2kvM8WHBPu8nOFnla8qhV54Spm53uk0mv+1KIu1vqnosh5kUK+4UbkuzA1i
ezMtpP2YZzfTe9DBq48epZptdIXLml1K3/hij6HCbOwAWhRA++1011BHznlNZm/N
3eEkvJXmycrbaXUIqiw40BhQLwSw0DlYrzFioyUeTiyfJr0XXNGd9gR6XoSKYFWS
jGA8mXkWDHn32YiQShigdyyKbt9fJA0TieDcHCv2us65KDdnXV2CObeNuGCbdjeF
nTCWW8vZFDxvHUa33GFjBBnEdOeTkhT7p9Vi1yAA1ykvbBEmVRYbQA1ArMVcqI9V
7FKEqwY5HkkK5iRORAPARGdyjTgSi1tD3SiQHWiqa0ESRe9LK0drs/kU5P93o4wC
mXworsyFA7nS8DzQ8vB2Gvzr7YqKoyNrS6pdl3pxx4nZ8Gp3FPg8AA8hdKx+ABtK
1VhiSgUcZnoA05uLfHKb6ACLO4GHNqrXttNIivjshDzuY9MeQf++qH9nmL6RzytK
+WclCwnCQeOfx4hNaZUKsSMPdJkFVc3Ab4n3UibpXNYfZkYMvp5U0gnEJn/qzglZ
a8UFi5iafqoet7aDYk128hvIe3DRK5J5LD1JWqeXQihkEIQKlNQsu5H/5IolNdMD
ZgkoLNI2ljp0W/SiH43TKwGLV5EuouP/fh94lfErYI0aHrYCy1EbKUBBj+28UKhr
ATGyEGvxc1pem3LKV49bqydnSBmMFrfI3qFJ1JPehXUyMJzeC5aAlqnUGGvX2+XX
tyT4a+VNWx0G7hhtJ/DWvezYc67OxxlC16JUiM+Uk3hzrQsmyTshvp3ZJT2uJ+EJ
wnIXV1akRv+/aQ2U912xTEv4dEZLnDw9aRA9s8grm33pfHDJ0PDG1qFpj35c+xSV
rEsDwuR2zZFkC2wXi4em3hAfiikKzN1+LwXrQ0l+3x5Pn/EFhz2VmQ59tdFhK2M1
IVe6NAJllWLEcnp1fVjUPuSJexLU9vVvp0M6EUG2U8PPmSIGuX7gVSO94WcSh31g
hQ18731n4YfldBke60E1gKjyN+oGvVruw3SfP5Rqf1BrgaCccoJCnHm6KQMtWKMF
VvRLsyuc9N/9NQHSpg17Lnw97LOHzqbyWGCT9AMp/CHzTca8X1Ce9hcFjjFPbbxz
vXrHMgOpgFhKjk1S98np90r6tsAEl7XSZ4BD7qhtN/h+2ljibnatfNE+zbIjnC4V
p//AwpH4dNuNJTe+TYBo8lnSSxQ0T/bwoZyAgyIuUmj4EYEzCZa56lOWjCmMwcnf
KjdPiMbCVXSZHCtM0kyN6y4vobTvo7xhAOOkg9Dmxy7AoeTuL4/GEqNXPV9wL2CQ
uFV99SPlPY4aJT+b5QJJRSvntlNxr/1YWGeXqdzXqHcO90/eOc9MB+xdTbmSiv+P
XLFMarU5F2HbQu/zFRhgm/cIbW5WcxIZkZYK1Wl/8iA4cbJZnz+5Q6/oJdXAX8Ae
kvr7h+k5PX6lfD2lZf1OxfXscnoR02fTTvIWVx90sn0vLZ3ZBScHeVM/mtPjvc9a
8uCjbo1i5A1VbQTkGto1YXEb/JNkF2EPIXXNpKpRaSD+HbYwyx3bViL+/i+MsxmL
5lnLCzSFMCZtvkgdr1+wBBLqP9JzWvysVRDLnGx+o56WLhdgKX0PNKNKDhAtpJz4
xix+IrkPPqSwt0Z5t+aQ8h4yqIgz0sMsc6n4Px+2zOudhN2lL7TUR6XS0KlfUH7s
EWqzbhvXM8JLg30xrGI145M2w/TEe2i7rm6m6rqyUr6jUPaSSXDAL7yMSy8GiMWj
7e/4/+D8P6RPncRGX61IAkIaaiy4XNWX9n8JdUPUrRLHjtItMChtkcth22OsEZym
bW3huLxxI1a0sAGbrFPrB0nxV8sj6+Jfx8Ny/Hqgv0GX4rxrbxSCVqkayhxVraB2
dkyVCsOvuRbOG5cDPUOXoaZOp3DKjfG8nJj9f8G0hcXurQOz5RqjdHurAFURZd2s
/M1FzESqwPO7acC7ujSOfKlKs8GfI015gs//AyBsgXIORLPuF2BnEbTE7RvdGQ5o
a/HrcZi7XIJ4BOpJgqGz6wtwji/EEX6O62X/TOvGzwwbOtrQuq4gOGwj0oMSXZNe
lrDgzFsJeTjBc9A0IZKuvIe9tiGUd2UgAN8m+e/goZXeoS6Hk88gCWMkOn/oWJI8
Erg0lq4hMk6K2eDR+vvGUYx2UrZim+EOhpVFMHVSX+j1TQ1B0byCIxCcuyUZcetJ
IofE9GDOD+8s/DXtovh+3ACCe7qx4RVexgPvPdmaWzGszcWWooo389aUibPJoI9J
5cJNSYXbEA8uf76DpZcPYxTL05zYJdbkJHdoK+v6Us/BD8GPOf1HyPKDtHc/t7WS
dEDmPePYEOtnkCif9DinUeXO/BnN7s+GpYD3S1WP8Udv8jgKeISJcHgJAE7FJ1k8
P54ic/+NkRmlFATBNnOiUzgcjFtzOwxD6EobMbVkNjiKV9MIJLQrE3Fg/5r9T3+H
hgY2hsFugMUy0DLioA7EXetgLoUfxd5UycpaYo8mM4Je9h+jcNlgKpLO5wOtuq0f
0IoEk+AsiVIFNK5shhB6D8GZ5+fgzyBhOBHE9f7QLxPik7wSHjNsgnelmOZRE1RL
Qb+r+ofG+8FY7yGWpg7Wbv0y/Y5dkq0WQ1fhTGDsxS/lmZd0nF6uihVoPToski/N
iwFZPnycjoZ4Ui0mYkdYqYVnDGmQNyfeifN0ZMGBeFxnDPIjgeUzKCb2+5EuSZBp
6KGG8Dh2+yGpqn3Ykr7jP8TumzH63eUAjyBs6ew1U3kLVtMU8y5sehacuFWWCJYw
AzeWS0KKr/y/7e3mUO72WZR4kEOSBLH0w1BpTVWxOi4FUq/UK8OwlCEMEwsNtRGq
UVa068KLbifvemaCS10Vg7YeVV6GVXiFHHtHoaIvgFpIGOzn6grzf4cJmbyN/wGQ
NRLyzGk1ATBjC9n1jiDqKeTreMs9/zCDlvFHXGnQigkfvXOFmmgSYC+MA7FC4EbN
0mRRQb/yJ56UBCeLexttdG6IorB+gv35Attsh58gYY5Bvg9Xd98cq9mg6CnC3yCa
KcF0N1bcMciqQIXCKIqruIqzroCxG/fowI8UXmhU0o77TJRN8JrX2yBxLXMTAjhs
cAMAl3Tp4+Hc4tJ/KlMS7MT9v7kxtlzoct1gM3vm/5NPQQkLw4Zc7GfF9Oyp2EIF
A/lKyrjKH08ZR2PphD4DOEL9sTrRrv6GLnPkStC4w36xmGNRYhOi+RrZKnNcFl+h
t4EZmvgdQ4jteh6N0F5hsVky2HzUeqbqeeIahMFCH9iQb2RklosEnbmKEPfe1Dxe
p/k6I3x3jUkmEmv9DX30OjmODVT7oakh5KwzfMcGINEOgwQ65LAgkITl3PM5+DRL
44Ykxm+I7udsYrCx4AF2Gt4qcD9LvTmn/z9ortROpvT5+txd03/xdPl93XIhhLq5
GYBzsDHUdMjDQFA+9AMb4g5qr45rv+lLkVr/aA8r+6BTYJ/tb9jBRV6Cc74iMXCR
xza9Tardj4HyMJJaZexnv7WuNPwJRg+ny7gTbvN+HRx2d5OEYJa7Qf1hU5vzh4VQ
lrSrf5TpuEB/c4Kim4Z5opJsKBzbuiW7ySwMFXMjAyPAg4CtF3jzO9nQgzQF8J/m
r/LGfCVtDq7Nr4ATfyHKUCg4vEKmbzSuTxxynCfIBa4H7iomHIm/X57lhUpzw8Gt
XhMCyfNdaUUESnT2YxcMmOBQZ+bWT3osCWxW1yhWEDhbJeEB0MLz0mY6dbMMcnaE
qSfezTaWE1HDv6LGOU2iRnR6MRyJoplAuWOREhetLg3OcXimPOSBM8sft8Znp8si
E1Dg0wOM847D/GlpvhSX0Kr1LcXYuPvsEJVADGpKCLAXVTNAmVs4L1ZFfZ2PCRHd
KJ+Sua4v4CIFCDOFcWfNeo4wTRPcKUZxZUAESobYI89yIo0EhMr65QtjwxJENIxI
p5lM5S9UjRXIvQ8Ysj9p3uNj66dS3v7+ibSGd1PWk67yQak9SF7I27Snc+TnRERK
aB22iGzG6kJCA7Rm5CqIO7ilmPg0aNY43fQJf5N/69M+Eab26BAovLC4WUARFhcW
D8MXMue35a3GiwLjdAA72hC/EQj29Bqh+aILx/x//4xE7pFlazfCkJVkMjKrgLQY
dUbCJRrf/Ia8ZURyckgCEDq6lC4Ys03Bascjq0idVoA1MF0z5MLIPD09uT/ALX+3
4FoorZ53EjXeRARRJ4LWvNdpOpA5jMgP5iyEe+xdBjvuFLP1VG2zELw+f8QSqgxz
p+nxbc378Xrg6gAddVqgvuKLUImUHez20eJPXdrTD89zKVGYHQu8dNQyQOsIlRx9
o3tRFd23L7tIGZx/DZEN6jVyOLcQ+KKQBT7rXeoWcNxAZoSPl5f7dcIz85WBNwvl
iTCa19CN8mxTxlXlGrLPWbsZoZqYrlv1VxqxTKSK4iSHrhO7nEnnsO639NnjS4bu
1eDuv7ahiOpWn2dbK2NDRd1hkXzNTAfnQRcuCN4WZBe2AwWksuyM+Xa6WldM46/g
wNvTJQmalOuBVKUM2nb1d6hdxnY9G9Kdpda8T/jb+L5SpF4V3t7TdVp+ILrjMeMR
xeBLLjxfkCb2Ey5gKsuRWHcWSn2DiJfj78wlxqhWRvoAanCpLLABuDmDWFLC3DZJ
r43WXK8zJZuE2xPZIWbQ/gjcV8tRgeprPbqjyA3Yd9pz30qZbZdsnWLWjy9mjMLT
sp7zfzAMbo0zvH2vJZ1yxYUvB/9ahyFMIaplvJASrSav2A5d1glRLGTJjWoguIdf
oLD2OhFz2JfKfJRbrjDiGPWuOD7D7YdAzsQQ9BuVJw7gw1DVsNZ+259C74rBLDi7
AMAxQmI0N0ikcMzzGFx7b3+w2au7JqmGoaH2uF5IhoHvKJN6h1kZT6ham1nf2czo
//oonQG7zVwH7QaxvmlDpZda1nOQemwOfTj5T5c+gcsXeuG84BeFHzUoG8VCGMyT
t54abYdkn4u29RJOgffBrGz1gnxmeHDClHFgN49l2pcUgTa+LY8kLzhO17ptEKj3
lxBRl39sLkhIKD19m/quOMe0ukN8SZVC88kqk42Tr9LGEa2Gn/G5E7vt14xomucA
nZpubbxXPJi8iq6uq834uVBQzeuA88kLbXTmHVCAjOW/6FHjF2NlM8Bn6FYrKllo
lfrbSVQSjdm/Y0LAqqz3ySPfEsVXHxf7l9SGN3EjpZ7F/K2SoOjjU3YAVAFDp1AO
SN/Xg5eWEklnvT3CqAh5+Z6ZiIVvtwyV6vYf8C+cK3bo8kK15sQnFcXe+HtP1Swu
fBOKVA35OA1Z5La9R0g9Cge5ilUs1NSprbhN2CbPXrt5ZJvJU/bqpwZtw30JVPz+
QA82rNR+tvBUd5kDJFyROrcCLXRZ/UAmpeiZYaGTaBLEHVCDjJXScxlf3cKHeazg
B7xpj4PJaJVqskdDoBuMI69d5Mwn+LcVzzDSqi5hBqhwPoZag95vs7iMXrqaTCJs
VQau9qhMPbEmauYiv0aao5H22NR1oXMZew704/tzNLMTa2pkruwtA4rK+9FVjIov
vP/heZkdUlNxETft2dsdASCj++JXGv1CVWajejRNWjZjTTWtihTs64zY3phi4pF4
UV9Bsh5K4XlejumvFpNVJkx9qZczR4yf2M2rQ9XjmVAXp+34p/7YquMJRdb6JZZH
GQ31o13uk7+vb27qwlxAA8F77zEGkMzI7x7Da2PpdoqfUx8QYIHDEJnNd0XGtBW7
0K5ZMi7H2IPzKib3pauSQWfyvxafr4OXt9i7RG7Iw1E4SB2YDN+ObOLqZH3iWYX1
rLfmPucjjVdMxWKmYPJrZZ7OT59gMgP2PWox1Q6IuTpmkwnYPR9/e1Cn1DKkHzBz
ElgJjraRHplAkCT7TXJgQZ5fs2BG7Yh2pWZjlqNU18CAviAq6SVOzNx+ltmROBRr
oPV7MaxlYojsQGh6hA8xK+2mN4UVNHuxZmxdplaYnAL+moleIlUymhK9j6dYuz26
RND5yE2rG8cLm8G93wxdU4dwf6TV4zuILygXpnXnukwkZZUV6iaKKC4IqHMiRqeP
zbedHIIOx9H6h9HHhSGuTY8BslJ+v6VhSwProT+VVTCwrxVY9qu2k1stlG/WFmYf
yhEEgw0eZ8WMuz6CRk+t3GQD+Kfn7u1LOSvBiL/iqQgmkPWhIK4nq9NaptMrcr0I
ZAbo61eHKpT9VeU7zaW5gOtKRSWEYE6CgKXlcZspyXuLYawQSnOK3xCfHybe30f5
2VJbLivngJ79J/0wxSTG8Qzj4HFk84RkTPJ7qwnGFknfeTG02fe8Qi4gAbz03Bkl
knxIqtP9JulCr6kqu8TMtfYHCcBguX1eT1M9I0Cxj9/cnJ0UonQx5V+W5FNl8YQ7
Fj5lVx+hs4coPK0fPcntOv3USVwPZKMx22/0U4VdEXYhkHi8SniD7WHXvm2Slejd
iTvq9iQQcJYRsSA5++cYEaBs67uir+ADACcuumsl1btpjE1k56TptBmkh+eGTNZh
9hi2DrgBkRzwX8ebSlpNh3oVg7hOl2zP1zTVzntSp70NYjBF+GCDNng78K9NeS7V
KO/lvqTrmzAt/MYT8K4hiIwCCI8JmVpRutNEDS7EC8vMQsyRc7jeWayP0JVOY136
nm7+4T3UAphPU517uyGIOzJALwZ2TcPTZ/lh8olyK0Tz2m8uNbkgvNsNe8rs9pjj
xWHaFaY5YNGQRsIozH2FZh/NmcEkfZ2Dd5W3rRx/Hr4fiFqiHGAO2KPsqR8HwrT4
5qOG7XNIzSuFX54QVL2L/scE716ew9gjNLdmyUTCUAfLpHYcSWbvgFPPtRr050fx
tuufdgPJ2cp2wLVMuFJlAuuZXXBkvZfs5C3owj6XAc3OG6I4FdiwX8kL02wb3wz2
xaTKkE3wzAaRpFYqTuFCbbCmttBtE1IvH7tI7xuNYiwSzqomBKKkwaxHpKwaHIv6
4HDNuhmDdfSaaWVJ5Nciqrqg93YIlAep6yPVClkPVS8bGuTXe+CbqUF8Q+wJF9zI
3VuRWW9u2f+pjxtdYwMM7XcN2y2OFXwxScyDExzUe1NwAsiF8gHbURozqboKfbaJ
r2ZmCEAGLIFwVCjrdUQU3fyGLec8CILczgF0vtm82Qyx5/4DF3ae70mrcccETL1R
jaKtyI0Kvto+UAel1jxuMfKdLZXLNR7h56UaVjrL0AQoyGXa/6N/boy9eiaOV2s8
yoHe11IVBzmFoKz4yQCR7VUF7UaowX6A1XD/WXt0cmjgGVW3cA01iU16auAWXoKC
vjNE4SEk+ji8TECByut8NUoUOh92rsA6N6ONPKgP4zJ34uwN08uvtbfUdiKuUqkk
VtlDaRLuIuhqx0AfffYGRZqtpBsBphn3nE7Ru1XWDN1sPvuYoK3P5r4qWRTfSCXz
zZFAl/EM3lMmMr4I4xPFmwxX1zawI1HNRtc4HBzcgm8CQi0qsRefWOb0bfxVjJTX
KaHDxcbP/tLPoANbV8EqOUR61NxPMmdA9J8djaa4DaAKxyU/xpMQTzatmIfzu/wh
bwlA+Z9Qg/cnNH/Y2gKON2RfH49XOuwyMQTXX0m2JE7BLV5f2bNtjY8cfwSANopj
TAVvHyToswfwuCkKQsjNIVCaK40u0GtwDcE5sztrElOLTauIrhaXHZvKyEMdLasq
Rqygjg+Xum8bCyxgvcq7AUd6ND67BMVLGbSCq92gqyqQd4dyfHDsd+8Z9pGfJgsd
n4TAT4xBK+Kwo8mR7Od0GuQ22bRTFhminJaK6YUS6DD1EymlJl/852M2A9VlgVGP
UXMeFemzHTmNXSjm/o2bieydOq7Bx0eTwoN1DaZ2y4tn8vlTbxjg6ZAxT2dlYSTE
nnUSuYSLjwVUdP/8qBFtuYZu2ohJHg/Kc4lsLJUPejDQrBOrUvGEy+7iN+3Lg2dF
ORSa8DVngiNM4u4SmVSus5WoDvLmKnuUrQWf6gDXIHcN2GHlrnHNnBex/oQzPJaJ
oix6L75waA3ofCTP7Mr/YjC8C7AOMwnZee8xshpUf9wHEQIYlmcrrmIOFEqIrRZb
8NH3soJ3J/cncdLiC075QKhV6WvmkMCZml4bdDx3WYqVieborx/RVoZ9sgHi+Q5v
4bzzhwJAD63xydrezc+fZIaQkGRoO7L0yuP42ux2VjBUybQA2wf0TsZkizlvx3WH
SjUJ+3pJbwwJm7vEq4CceU26oabqq6AIGub2tdQd+6v8bmTp2tJ30dk6TBvcwkri
ONgWNu6laKMtZUCzs3gj9sdz1ggT0aOcOq2Tn+x/bH5F/rdkIdz3uxln/zkpfCUd
zfBXryu1Ejka6DbXkb19kk8E6eEb3Yt4GZAVNOAJ6NegvKxz9tcR5DUi1I0BpScg
kT+2sdWyuIq81dZCSG2Rujj8mdD+ExgPbMXJOdJ0Y7XQzrOpvLLHxGvr+33H2F89
LfVjq+x2nguLiB1pYjBlantL0+qYAvwsNR+ac1hzNpSFZW6cM2I+yPUnr8XOrFhc
c6D1AkstyuC1KhpVU4LNTtlIDA2WOxl8KxDsodHVWE0S3lXnXv+2fWAIYUxCw9nG
q6YlmdA2VRrWU1L64nqINVEglqPTIPwMz2nInMq11IQ/SHI8qEjRfuXUZRXoqWoz
o1SJHPT98NjtRbzMA62Eo/ZCY8fd9taLb0fnvCqXYfUxRv/9Tol0SngyFmjFT8Nt
oztjE8ZTbt+GdOMD7CZCoVFegHlK4pSKfevOZ1BGYactjJhsVabr5kYcGeZDiDpd
8SNhyiAG8ODi7ZFaa0hgoE1E/xSZA1V12FCumJg6qOAo+jMKS2n0VWLxY0JUDFMi
9egbXzNtLGTaSCRaeAlcDAgqW+g2Z12Y+AYtwUt9x3mRRUEDKRukx/rsF2F/al64
SC60bloqajd4pSmlXLoSm7sbz6d2WiKzPui0eGlW2933WDl2GNeJJE1srRYMXhx+
eakrvmEr0XO4IdtRX5tauD2Hv27sPecj4jeIh9oLHovX1R/vMBa1jftFswNZHz3U
8e0B2uchGcgd1vxqEn312laf0e+rrE7wv/YIPByFN1H++SH9GW4uuI3pj7nF1l02
0x/1NAFCljma7Jz2ep4NcUI3nVImmp9VT7oYrCSjc+zXafLp9xeebEQZfQMc9mFj
BbH0fmmzKybhno/9qVoWEGWiXWMso2XS7tLFx3l5aARoz2WLZguMfX5anT/ji7yr
FLdBA/6VAJoqCOQRSabSEdiJ7SurliGHYWXmeQqcbD1m2LhD29mMyeTqRsK70FIJ
yllNx6VZaJovl6niyHQDnQYOyzlf6PIzTVXBq9EKwBqoXgOCtOO4lc1kzcNhAZbb
3wp+O6minqM/OP6ei8I1ioNHz+1xwGfLlw2pRFmMg2/4SKvmUaJ1yxmi3EhNvLH0
HKggMvVsptVKCIHAviwClIoTQlWPn1wWoPaWTOfRxvOU7qLuDv3d+4QkYS21J2L1
6+NG8T0w4isM0FFOaTWYn72TlxxtEg2Epakuw0aGys4nGSWaRrhoBJuJZcwD6sUi
U/FkyAP775YgGrxg2Ht0s2dEAzmQGEWvRwGcbUY5dcLFSkRR4o6YHs62RRtJRAdW
C6pkgrqdVY9fF3ZHMvv7x5YaP8FcJFHPPT1a1VGJNe+LQQ0yRLz27SyHui69V/Ca
WIAR+9OAYlzmLF+PKoFFNRhOEAykJoScms8s3Iwd8MBAdBqVYbmASPlFFPtQu2BV
5AFI3zvV2bbJYdxT5qqbrg+jaUa3emEmoE4a5SAxg69gPOVkFz6IH2g63S0TMy8H
1ghgvZxFMlK0/c23cbbw/X2KLShiI3jaIEe5NQU4MFJk29YXJB7shsnL3bQIsPma
RbvBFAV9zPHtVNpIsagAGin6ub4/wfP62M8yVNv//651ag3vreKYdegXZ2A0JEt4
3SjrwjLDCN9cAnGWYsqAHz8X6zNdfCDdD3jWO+MArfZ8JXphFDSmvCLmvLI8bm0H
+doyJrBbHQtQZ2xY61Pnk+xNOg78PO258XVFiu1gEjC/YJNVgwHud5GHSDbp+SC4
nHbtIz5gboNlI+mFbYymUlJUQ7bfVowvJoRqB3m/iZSgSejjogZwGxCJvv+q7zGb
BxzcF+/ZQbr78bFpV2ZaYQg7LR6dsgjOsgXIapmUj4OAHm52SsFBIZ6WsZ7MvoYT
ArS3ni0IjLeINY18iyWZVdNVYehA3RT4arOPecYJcWCidgrWhT08xYVP53ZmHqbY
RczJPnEZxFOhrDYRZN2HsRBFYqc+39C/O8+Xx8xBo3bKWymEmhZZFQ70mPn/mfez
IO5bcCsPjFHP1Iqnzk+jnmdgrSYVsNXlafjlHB84URDci+VCNNRd0FnaisvBmocd
5RfDh0CLuWsSQNkFZdSzDfbloeXH+8cLOl+Ypzk3zg966DN0GPasPtC1hqYMZyWl
+IhPUaHs1MYkS64ErD0d8URLsRUANxvwlowWUFVVhIXegsAm1OY1D0X49izJCLqe
n20NIiAyA4ylGpcoX1V3QWyQEwx/YvuEj+um8Lzyx9a4fBOc3Nxox5bpCKdSxY2v
ujKVxC+nUID9n8gUWhfhu3x24UvbU+bC9X1Y559hPrmVsu1VE4qgpcmaq/6dETS7
HrPuiwADjYc6TupfxztLBGH4lUvEir4HkLxZWbrF0tbQbQ52J6x/eJlZHMHO3h3S
lDPLyK8gsQMbIPTk/1z6sbalBxLsRQ1QvFG/971On44Nnla1fjWydckXKT274PQj
qs/2AOFdmEskLSb+LcwvsSS+5KuwgdEbOWuUwSHgxUleT87QtCTeDzv6m9Tm9Yrn
2tFY3jYosYT12Y81ICXSUSW8VDgubs3a19DIhMCZErRX2z0n20odW/2pACb2TKBo
tKaHQ8NTwq9ckWbttD3jH4SQTd9T+PoSbNKfmrZy5kDaR3HEvLt906yewlAOP/I/
HzUOYnbRmCHNIjZAKU0D3lJM8VnHD9CjLWjp8RTCkUY3hn1nWYCa9bR0YilMWB/G
1XCxGkabzaioytdx5ZyMjqhVrRnf+IT/tpnIbeU/sf87PFZMYvnohugBPiPMy+n3
ws/SyVvwvzymm1gWuf1M/ooWJTIplL9kAwfNFQQ+F5d8e4oMuO6U1Jc6axMW0Gfe
D1LQ4X32vUgQV82QvaKJ8NXuVckM5DNBqVVlFDrnx1d0DkS5m+yNypwhHAaHDV9P
vZ8DXkO0QgkEJ/oYaHEmYLDJgiAUeudusvIVcInF8z2C1Puxa5MtwW9y+M81lLZU
Ke+zsQVffGmDejAzwX3o0NVU5piGnR3bN4c1Dn3jnmKJGOpWSFO2AiHiglPT8sy+
IR/+BWqVbUVh9nJPGqYPAjzqaUZneD3sbWPFzRMGXewuTJrSm6CMbJP6dAx18RSS
FsT97Lcg1MvFcIcNGVfYeszI5gkjziXJIzt3PjsxJe8Qns+hsXtmcvKdstRvMtMg
HrZsiKC34Rn6IyZtxmmq2eNkiVDBM8XaDRBJTxOjEJwX9b0fPzcdJVmyC9RSxDcS
vCaWmbmXJ4r8sVnQyB1fiUMdY/A+PjzU1ch7Rd5Yul4X+M7b6rqtA9mhicHnVWZx
n+Qs4M4PtpEJXLPOe6Faj2yoK20f+HEhiiv3I0QIGmV5SO/WIEOwEddbznge7FQW
FPAGV12neNUNhViYadIJ7Tx5Ooa4hauvlJuIv+2/uX6C7sd1OgwTJjzQQjQEmKUd
Qj2H0kiLzxGQyTcIyiay9WauIxy0i87O7f30mSIS6JkvB5h8O7R8faz7t+KG2Nda
gg54bJqTqy2uRD8Bvy9h+ScyX5qOTIZn1bisgG8WDbNEsaCfa9x7r1L/VXrARYX1
y2Ip9G6dSZNnJBQch3Nlv8MxiJhjQMSdOTg1EcDBh4pQS5YvEXZVs2Gro6nyI3Ss
6FSDt35tKdJGzOcG6ZzDva2O8FmBJTaE88fz97DjBhsPNZ6n6VZk/2YM35AWCWk0
MAdU5qyZVHmZs+oBd0+P8iIKLqkAbI4IRq3lTOpPS3KHsabvb2uuWPB3yVdKfrB0
x3bR8U4btrBVefkpVylYsprFJJNeZrlHyz7Z3ATX+wYYuVSzq2n859Stosqqkfd3
h0sY7V/ZVTQPaO0l5DpWj4JgtMyG/OI5VdF/okBcaPSKE1FDE0m65/hhsKCwcPHc
1JysEuis1N6dAmsQZBTiQjByK29+OCxzbsq8Du3sj+MjqAAs6jJCQJ2prZUHvmjy
2KLEdirQUyZt3LcEf5jl9ES2oaa4Xi8iMxPfnS5Wm1voy9Du2gHFDlTcvGHD1O/o
URQF9QQT9qe7j76zJcG2R+R5ed5oATLobezFDZuJJd4ZsI4oSBDDWbjArdVSfEyK
BgCd8T4jOM5aC9ToL6vjt6zkrPEMESIs3AcWB3xgArwCmHM17MmyLfxCJcQd029H
0yG94LwbDjJGSZIPH1b3nIDlXxxkGuRAUHkxd3N4iYsbzL6syH/nmyEFJSN7Hjly
l4XcZ4lsRnJ4gOuY99anL7U9Op5VjkDkajnLd6OdrZiUzaXwUmix3h8+Nk02YRMK
mIUl/Cmlvzfw0JFCTLfQ3AIZxDferbHquLZXT1lUr+rxK86drjdmRIt0ERZq0R3w
8BDNMHRmuWw4Nrfwq1u/3y5pH+1/Ztwn/oDTPgZcNp/BcSz7jI0u8cXf3+EkKzNz
Xwy+sWqNgGdGDKdw2PXP4Dq5zbleQQ5vBPoRuJLs4hmnAJu+z6nZbhg90F7mm87F
PbIt67Ljb1Y6YQJsshb7sOBqLDCFOfNHPVwR/8wP4v0LY/IBNt1g3h+9oLCT4XBo
9ADpAF/wK56nWDX/F4fdhr/VBVBtuW1cH/ZmAjnnP1PGQ95dqeNQH4FBpo3EpxDQ
OwkoVQAOaWEM53w9gdH46gVJ+RuNcHR49YPIkZS2SE9r1042nKuWQs3EA1RU6x8Q
UhCm80dcZgYwBLY1//IgudGtT5dtEy883kZ1pXDmpIMoLs4PLZ5JimGicXh/DZdq
HWJ/dFUOISBSWFo35sYiTGm9dFEtiLQRz5M6+NUWn6SkLC5dZdyq/tERmaxbIZei
fvxRRtScu9gfiwAf5k52f5R1tq5GwGCgmhpOJtWoCAOqU0RD3kYRMQPjGLOcZFki
muTVf3EwslI1f9eNqCGo9ddrS9X52Xhl85P3GghL4SJ+Eh+H7VN1HYJlOBX/5oQu
hVK741RIT6UQxurkP2f5la6Lq1ET48/tSGDkzAJAgN+bShZVPe+rPgfcBqLM5ap2
M2ll7FRnlZjtw0SRaXWsvu6BPfSecU0PLHV0c5nUnQWNyCsaFceandcbWOrw+0Ua
YydTmlgShcpOmUnNtTyGIJcFhwONZDZTdydeFIGyjlJtj3QJqyoKctl2n6oKJMmJ
DK66eaUB9CRz8HqDHdCf0+KKlZr7+9mDhoWQQet3DfhscD+SFj+WMBOMZGWi2KFc
E/R4bZe+yKt1xpPsHDw9c/o8EWqWwFpT4XGQ3AGN1r5F8wN93wnW/ZkZLzzkz7+V
MgJQAOF2WZ6mIoBsDkdDzbVT3OnTw0LL9PUibN4XgE98Vy0rRdahjCwwspmPy0v4
BZi6GajtgU7PwbF5TFF9Pu4NDoesOMnxVakB9jQaoEJ+adUBwv6xid0nipJuLiUG
SjZ5IbXc7yidLcYCzP9TolcFvUoZTYPREGk9DvCKf8JJ4X8vDLKp5MDOxyCpWQOQ
DN3qgiu1zSYWL5I/grlGyTkbqbb0rNKUvhYPg7rQbQKCbSAvtDlO00MdVjg4fYxI
kpx4SwWM7CK3ouezGe52dEl7iEcigLRxFyOucjWSdIKHyct/l9a0e7Wj+JHaiNVP
KRN9roHzY453u5W3eNEbNDvgpPWZs1HE0XTYwyYPIvzwjKrqWJj9m76HT81Tz4w8
X/sJVucJLSuGJC5MUnwSSB327He1DjrU2fOWokw/sL4tGAlZwlSNcFFH7lH8w8uS
g8K4dM3guyt5sRJn5uPQNsBCQpr+A10SR7T4ABg0OBBhHPvtprJQNhHA0jQItfWm
Am3g9jIU8QtTc++la5P1GaW3ebwoChRTiTJIS9qDqcWRPMxF+QfZ6FzU1KzoC/tt
5PI2o13XfF+wkMPeB+CBr7D6VuXfa1F/Uhu2FSwpJU21YKm9hvxgapHwIe0+lSEt
+bhXSPIdYuch/ygHyNKINwxx74R4aE8pnsc58RIF1HApbzDovh9f3X9ddoXPfXWX
97NrcLbVoHs7d3wWlzI/5dMMA98smRX4x1/Jm/cWJ2rE2+G1R7brSJMifFlXWh81
dugSjv7Ut193BX4MH/5jZFr86sOZ5mxbnvm27IeX6Lf8ed7dg6eysTg9Bucjn2lE
qoyYpYzj4E0PGd6OewquSc5xssev5qQRokcwh7xnXDBKFSorLAL/TCLxeYbRBZ73
BC5pM3aDhpOTB5lcSN3RDnILonRwA6UWaL9DUJZYr5K1Cg5bWhF2KWz4ZYL4mToD
Cy20LLJ/IiR9GGqD/u/FUP4s87QrG5SKFtO9g1n3dWVGuHevz05+xf98MMS6jIEI
56aDgBBpUcctLR19BLSslF1kM6ys8XlEgSBw+oWeZJa2NT5Shis2/CtUPdda707f
LieG4OiPcDt+8sKRrAAEcxBtBbsLTNf4kOD35WwdyZKLwE/BDCg+NqC7m+Yoj+1S
MCYEl/mcJAMXPfRrckil+Jl8ToAgnzAESJvUv4bgkoI03qV2fOdJzLA0ZVZr/+Vg
opRNwE7fXhufCoVjx8pQKb0nNRILWWkJZsMSPi7lN3UooN6OxxFi6lp7NfrK7SLP
XCIQ0SMD5PiSPMBXl9wjDs9Np4yLMKxIewothYybT4i+MVQVR5RbqKJlqyjZAeZp
1w60cVsPeL8UBa4I5lEHtYORAlnxyyvv3Pwbj3iDiTh/VWB3CJMNI+ns8S+hZ/TC
FvrqgnxwtJiW9Wql0DkirJH2+VcLnRvzmCaeQr9ckLDvdN2WurMOjQzQAEvBCk72
bYJykm80p5ccgcuWw0WoiRvvntiwW9hJLeXghwzsytb7CqG0SE1e6phofGIxQTVH
6S2AycxC+RisN266beYkZQAIIrw9b1juD6rHQrw34LiADZSgmeigDQOfS9RIVH+D
duyrlxaz2qnr+fj99AJ9f1pqtb1OLgbvkqC4VoK5RaEMyork8oUu6hbYrxKt4Xo9
C6ucFp2r7EhUr9JbkBf18h8qbjRV7gK+1tfIoj1L+P24X9t4gtmEEyJpe8hd+1nZ
rHceX+/+1xYfu1x1BwUWwajljms58+kQUyE/I8y/xjV6/IQPTpxkoYffZ+UNtIoY
9MyXp33qEmDDRluudSNGYtNygC1BsyBdziPaU9m72WDTMzHGXcxB69laCgQ9n+f0
i8jlXg+hDEqQdVl5sma/bUJBbvw617a6NMSdGPEmr6OHrNVUzDE9JUEMLJN9NGhI
Wtr6BcDgTCNhzUsHYjI+YdkszhRToF9N51B20E+13snN9/wbsSO1h1haiImpHjmk
R6RzxvhbYJyO4O02KcdnTAvhO4xRuvrEGK0doU+WqVvJ36ZnMLFMV75Q2g/lGoyP
3LuIx870ne9pzdcSqus/s2Jiox+4ETAYHDdNfD9sTjWFM2CcVDZ4fkypRj2FFQCc
X2wSlZuyBTGVIVDkIbTs8wsnnHt6SAI5Ja2nIatmexeoPfOt76rSNhiNxhzp0VkO
BcfK3pstbq05jt2MIKG6k3m3ySZ1RqvWhPfDBWY1MrBXNah82DoeOludBuNSoaBZ
fnPwkKOuEHd5iSCRhwUy+pbhT7HlfnS8YSkl/s79QkkW1RbTTXTxxru2Bp4acBQV
XbvR+rJPh1DuIh6S6yvroFJc86FbCiWi2ciRkO7OJOIvl0bilIwml2xy/Y6BcJdf
n3ycTvcdh0c7JQBQDpH+5Cx6Wh7rLZISLVARRAvG5JKKnGr0KB99vWYKvkKeqxiR
icl6/I2EWeSHxg1iolYaKypZ451FgZhtiUCTikX9TRxCjT+xEI2oJ0/F5lDyK5Ci
YztGd6ysT7lhlDlS69CJRVZPgtG+SqGkLPZGKQU2nwKSOHbG9jNhyWoLJj13bqhm
6VIjvRQgnnEb5BAuLmxKoZPjksFrAjOTgvs7uSdD37mQD5BrBS6q1L74RSvDH97V
kjcyAOZ+hrvnC2A6WYW+hf3I7wQCXLrMrRbHORHhsV4JXi+8ggH4oWCvcdPHL/P5
UOQrgfT5VXdNEI9GCJ93of0pYQLcOrOK7QgQSJF7SyfTHvaJ2LXCfxnA8FKG1HCs
Box3sDjH4xurRo1Tt6ukIkpwV2+5qBvALwfTAQJ5KIiVVk9nGBsEMym0V/e6IA4B
7MQg45AZllVykcmoD0NAvXFHkvCpWWMlzZN7N6zMKWGPci7u/ymEDNTjdFNoW9DN
jPZzsHLmvmvq9+PjUhTmzWMrBTwSN+kSysO87ssejjZoR+H78QFajC7pR3qaSN3x
b199DjsYWPebqgM3AKTllZVirgHEtLGqXKFnOY0ejUbb5TLdE7gRNFccScyz2kuv
0nN3MqGHywysXJrSjZcYBVbwIJUxRoo18QYDxw/glRjn3gAmD7rh9M5eDwnnzexQ
6CC7ozCqwvg8V7Q33udv+S1b2D5kO3ExLIkNLuOdC3mlDFeEdZO8G86Hja9MAO0g
UDSTuar9scvgY58zBq2MuA+EQOFc8LTctpRTttJFkqUyvbaJeIrhfi1+JbZ3AHkb
727mSiQ+esI1aBonw0P+n5SN9594Wk+1/UwxcVGT97r3AtsZ8fZsnDgm4Wbz1z+i
sdxTzsYInviyOQRzTtBzWiN8kfszRjAFy6peJvg/jMlAIZtNxKUVo7tz1ouop9Yc
aY1b+lvEHPBS3cAIOo2uAiZTf8tx+kewDor5bg0k0nt8v/twc/+oUV+a64YEhXNW
+6BaYaGwT9a+IdTv0bI4LvsojiAn30Cu/HmDiu2eGvlsEHaKi/10YXQZZT2qt8Od
BFOGdUqUnsmY9+r71DcTfCwIJKRv3oTykHPyJpJtFutthPFquhEDiNgy2zDNI1hs
74Zn0CQXU2uh2w4WSI6Z3RsRjYeBAcUhvI3KmXt4XyAZMbxlPVzPP5SIcMK5hglk
wE2UMIazAvk4P1pgEyLh+MrhgmG6WlnjXuss/Ilq3rRhBZ1/uP2+ilTOqhxCio1/
jlKum9tAcS5DrtbP/aFR33YnwFnd8MjOvhAEX2yjQ01zhBieJ6KQuF4owU7oSOQT
A4hnB4HsvdQ6CgXoORLz9ju9EA60+8y05zdd20HVB08SvXmN+xGyJPGAlC1yrLFK
azVVmnAdYVK9zadEN53ke1BqZarpi29xP93O8rujnJdGBaO+nSMKzfDQXY/7qpUI
PK2Ms3wl+D89w+hHVVTRaOnHus2IM/YBYtorRVrf3nZC6fxE0SyswT0u+zE1WxVd
o6QKmEjl3yZCEkYIyGT9SNnMQwtGU5jIIN8phgi/3l7X9ikrJWvoGwml9HB3lKC3
6wU/Dsl1iP4Q4Ag1udJBQjSn+EOQbUifa9uPiioFJsjRw477V8cfsHzwxUXkWQ5f
+xBlc1a6QWo0BeOLTjjSzTaPoX/wrX4oWv8vdcuk2bk/6wp6IkqfTcBs4gkYcjb1
Cc2h4Vvx1G337GsMoQZTJ74nZnr1qL1fjLcGyUaZr6+5lrQhHOAfZoqJ22QM7b1K
ASCEvD9YYXw3DmUtRKyih/fyDDVWKB9sq3pqUCzyvrLzvKOK0Kt+8kEx0JHkpySg
8rOkWyBAb1QoERf4ECqVbaA3r2WAalnxfXKxi6rF2kMCNMNBCc+z9j1Iwrbtj88q
1ckEuDaBD9OUBQnvLrM80GOgnEAK2/cWiE56OwQApoMnlfoBIm6OJqyfTK2uKPLk
1o8oAH/qorg18M0s0t8v+6meUSO02DcjwYhbfvjkvUlYR9LMva1DiBQUwZg2CG/w
Obkh5Fik8uYCEcKjHjxsuXb3VaW4EC+KJqp0qSu/RoN/dRWt5H1KI2e7wJJV2g2i
Irjb67wA0Iojnj7DoxmAI7OrtbDppBXH0MlsY1YRCoAlNXi8PEMvPVlQB0ItFN9a
z08nw1y+91cthBFRW98C0BHx5ZKAiFRDRdjLX/iAa+dcU98YmoscbxM/oQmhxyLn
g+uN5mJohCKaOPSDA0drTCguy3xx0c+HzBxBnc/o1D3gCE0ZqyxauaWcHIS9Wlhe
EBt+jzLmbqxchNW68H62nZCwCKPHWeYETJCtPRcSgOF+uA/A6A7xWy6jFeQ7lfbJ
DbCI/IVYnqRvddaQKCLl7pJartr2f3N/nTcW0z1BFrptFAFhc0opIraukuCs5sHa
TZNoR7aiP8CAPxAz9A3hIhbzc8HA+iX7k3R8U3I3cRzXrCypHB7LqhvKcuIv0g27
CUdPaSJfY9XXS4vteOPFzETJOcs82pq9fao5iF4Ud18rhE8xe9md4kXh7GRxrbET
6o4ep6ymWWJfoX/06j9YUhA4FEE0QoE2lc59wFhG5wfmgDbERQuI+uQW6CUHqDhy
Khxq5g3Y5O7vmtgDxpFlTLs4qrqXTizDbjudkEs3Nn8TYk/LgyU9zK7qiqNKBFP/
RxakJxl6a2fVrpVJA+7NRu122L+V0uGvKzzaSzD9yULeZItz7n3+GxGliE0xZXbR
0kaCI5gpm9fxbMBPFjdg40zB3HKW64IAmx7kwelO/+gWNkC0XAAWGNw/T1DizViq
5vkdafRMD6YeH8dVsoF9WR7bo6j1F0Cad0CJ+DGq0MYzS0HquI+HoTVi5K7ZEVkF
J7syLbmeUup++iGIwqKRruJIHftSZxGSZebR1bqyAje6PuR0HF+yqZu8LE5CmFT+
JxPap/uideXxg/5LBL4p+Vk0W0isugpCIurjGrA2nO6b7OHhkcRIOtPvlpTKbquj
SlArxYmUnZyAbmXEwSleSMN8SbfSCascLm36ik1sqFRSQvT2L8HVfg5GxRQ+iBhY
jIq99HQkR+7JekedKUHHOuM3pe+LMQf0jPzQbuohIA1iHGZhFWFvqUFfw7dV7vP/
eG6EmByuv+rKZbV/clxWnVd2/971eXK1enE9FXUxZyouB9JHAvx68lF3oZpV6g7V
i7dJVenrXQj6zlfvmmlbC1bGbOimpellhMSoWt1t9kqHj6S1p1DqqaHaiJRVZ9h1
pKNEodS/VR57HrOvAK73OL4yzlQGbU4r7pGq9n3JzqRYM5bpiEtQsbJekWh7NeN/
8duPwvGY9HKFhT0oRsbXLnTAMkq7ue9FNaRRoYxTb27ir0uDSqmEWS5CcA2BiiOu
IaYqVAE7QE2CIQnzJrRCRrafdIZDv6yd8JiSHPNPs0BNtDQKhm2kKqGZPhFcygQ7
/lkJh1g4+KNhDwp7R7rsP+fzbYQIIky7sUbHa4nvKWDZQXKgFe1JUo2oufJNzZ8l
2l4UkKZ4lRuxOqsoybveVkGI/5nWa0Vq47Sy4YcXOWnkkYvPyCYYf605WUx27uOa
XvyctTOotwdgWv1dZ2ZiupJYwF3DU6Lq7sPnN2iHc4t37STIrHu33HKHXxkfRJ3L
reLclNhKT1tiEWyFcRZN8cXKHQKcfI28rNX2VFyGgaQwCbqJ34h0VBbQ6FqKY+RJ
9I1v6p07grtkX+0c+uvFBi68EsJuilvUr6Lcs6x+aV5tlhCIE7MnqlAVVMg33nbp
ua2RwQ1f/jgqaNYztx5MBvd7Jejtr1K5Nzn2XrdlnaoGTBqVr1Xqb+IRCQCqh6ye
GwvHtXIzPriPN99KeNKMunmGsrp0ynhFKYtcI3NuCHb4qse1TXQyTB5XGhbqBL29
fM4VYkndbU5Kaij4bU/V8Pny/OUuw4Y3qAQqrJqqg2IQ5Qvwoiw/nciIul7h5RTg
sZImGF+NfphWXBFiWUNEYT9qonrU1yAEPY2IEUZlyH1aObDnLN2kQEKozF0ysza1
PRDFYbrmJeppKn3Ia/ehtgJNRfBaM2tQz7JapXIgm+eWMXbpRUW0t9xUrwBDfbXI
SetwYXj308e6uXgeknLbaL9EWeI07idvKcfrpGHIkT79K/KiRCHgcW/B3vfg0zIl
RBx4FrS4CddIPr5cwWyxRivNbMDTE0tiTesWDs/3q3i1/Lc+ONBFXfBSEjdoolqT
ON6GVjAp/x1iT3xacrlJAWdHF05R/KHvPX/XYhQRaKKTMEepRO/PKzQ0iur4IKD8
qH8Sr2CZNcRRBsretIEoXi4puM4YphTARcvsD2kHFOd/NUv1MOYfPN+sCL5aJ9bf
r3uDWpFuOwhlYF2m3nkjXY4IltfbLzX8uerZKKL68eY4htCJrPuoJEo2fdSVPbVm
vAVuBpv85cUK9GRcP3O9jAhGksEtwIKSZE9Wv6eMy3HSuwZYvmBNd8taKKzU4yaJ
1VxhQMlUrQ2PK7LPZsYJLxlduNkAV0+/h9QMPuHKXzsvta2dw31mC1LWq74E5WaQ
WYqErezMFLOe3vO6o6D2jwgbulx2iinIoyWSx7yX8yvZAxvkrf1m+5NOWWVYZ4/q
8D8z+VUs255lT12cKVjtCOrbXaaYCKwf0Wb5XD6wFGsvwTN3fBOdcxoa7JCwtBhR
lQwF/rCFZIog7Bx4QJ0TbzwC/dYNNV1VPU6C65Ay1yXRQreCpI8miHwUNAetKgEI
cx99Dw5UCoBFscf1rcqNKfsHLUDviYBWK+KMuALV/8qt2VKM4FVFqEiCDjPXFDUw
cs0imhCs7OVKK3s3OwU293qcrnBSW0VrFuwlmwDGTTRL1RKGztow5FCqtTV4iKT3
653ECXzhe2Llalwdb/dCkCcz7sfSo6b1a9VNGWenoanAHK1TcOTR7abhwAtb8pRU
bF8EuXlou5Z+b+NKXlYQbNxSXdUnTSnDa0mWBL16/yZ9obKijkon1ZH/WZHFfzMU
w2eA5iqtncXKPF/+yxbK2dZxi1IO+ymW7ak5BG6XNBhVizddlBpsgdCdFJ/ylB7L
mVWzhCvfxYHSxYKodLgox5cAcJSyAZV+ktqrhBxz4Kut0Xlr3Vbo3WR3tEAUGj6H
UftWAMXx6sv3vi6sCkzfsXD0WJi05xolKkLgA1N4xvvWK+KJqsHkb9aMHOHadvJH
VsMzZjYRtj+frMTzkvToC0n2KQiZlzzVZM03HIQ2/M46UyR3fjqYPsXynbCCWBVs
DzNxI7vcthDO5+Oc+JpMnTSJ0JEi4kxXDmPLO3JnNXjnBqqpQmS5Io62LSj8cgSY
X9bYcNjYXZY1c2QBkpp4M/czI8lmVgf/0vkP3hWF2yJNeCDYFKK+jH1DZ5KPr2Iz
mzG4nYRQ/LgXVRgxyKxzelCLpuk2pprCHUXcyjQ8GNz18fG5UwSBK/JXUcfljoZo
inMRytV+rKVCcZr1PpBGrH8WwYZOl3ddei8YGryEBmvtk9r8nBRwIPc+RejpjFRl
qdN/t5HuKzjct6sKGmIKkbOWKYzmdbmca92yQ5Q3663hCq37HPn0pukQ9d1H0Quy
orsPe4NL42J9/qn3JR4esLWfEOHaDSuQWS1z0SPwBG8AYDl6HjPSKR1m66XpDNiK
N7rYeVeG5fhaTp46GW104JE3LgsC0zXe95czE9Y4biofEDO56N69OwO3foByv7XS
zXmVyLQKjXtcaBh7fhl/qidTCKqUO/aLsMAU3vOPCc7EYssSjHWJ3E2n56MqJzH2
E85lJ7Kpifu3gEY+ALzosU9un0363uRZ9HLZZqY3SR3q9DX7K9E0DV+n0zSDvxjl
FZKo0xkYcaDCiCZAL2ND5+o0XCKkMvZMm8T0k+BE7Pi2lPJr7eDzn921cETwvmNE
bUycDxn7K3ACAs/Tcn4nQX4DPMlSKKYz5A8lGOP38bq/mTwaPgem9UqP6V9Ub9V6
/HR2Ph9lPAmfYRpJVJZuWAcFdqtqqyWHmpQcdGvz78BTrbdiirjXtmc7ezuTBn5q
Ex3PiIzN2MSYx+BLQxtZ4Hvh0Oun/659uEWiPYACoJzox7aSB3fhLQcngw+Jsbv6
SED0EUsvazsJKue8a3HvtcOeNhsY260S4avwj9TSjzr7aVAwa5w4QPd4AXQAJkrz
n910OKSugkbq98NNo6ZUyha0//x7aOYKcLtQ+mbOlL8KID/nRvJrmtddA3QkO0gl
FKbIdZnS2TLpw3TUVVom33NSWpVXtuH23Mu/GnLQGnSREMz9TTeVVdSzaQIIKdjU
dYixqRzlfwMGhTJ9HziADRlCEYa1D0ou6eUcWu/yJTNBfQRVoqFKGMsi3PgmzdAk
8HjSIgSNO2jqd2tAHomx15xK2CL8CNOdkicz9YsB8BISSpRz5WAwNrIuFhztv5TO
8jffVW5YxQFn5oEO1L/J4hQB06RU2xnB3i7Gu/ANHqvHTNobVaHQlVpcXVJC+LqD
DDnOv3fkOG/t8rEsY/6/2iBRi1e8XVkMo90pwlaPVpBT+8TsHbESCRFVJ8LcHgrD
aJiJwn5XC7ZVVGtQg/X2smIZHOtI+LqZyM57xGZgO/YTjaVS7QruDEU9FNZ4ayRC
QjQZCx3/o9Dn5pZTZoAAFWAi9798aGqTTO5/xtSQ3EukVGjt8EjcFMeSzHuljX5v
m3Fz5E/88iMvsWsrQWIE0WZMjpUXCDOSJlb26u8PK6DYwTcvHuY/XN78WqtPirFq
CWMLu3jeECiimFqw3iQDxtjA3S3gXk8EgJlzEKLzjZLve2ChhRSqRiRLtg5yHI2i
aPdySWFbV6TlxaU0616m3NsXh8XE/keMZrMaIPZrFZy/cp7TUkREdfytYgmd76Zz
5wIP3JptU4VzMQTLK+5hg9LDT6jIpZxiSLUsBoMZh2gDxSqk2243Woq8FcqxeAzi
oBPwPl1DbpRSGTmlHzXqHqpLFUm+Cqg+TBLq4/iuIphQsISzbLPAIZO8RvmvTSta
Qh/1V8Olhe+I8sKBBbOmDedyGlnDAVSyRtTcNL+PG0XKBBzeQNb2y89Lc/GJmcKR
yBDalZzOqYgECdYu+YnaBpkjsXLLbH+rzAkn980oTeCGGg0oIzi5TSDH8oWjTdue
MGV5GgNml9g8PDmODEXsSkjhxWNPwkL9VjEFBLn1TAktwc0PqFFMrWHcQVjG/S3S
fawwS7vxSkgdyP3DxM+yOhByNXsLgs1o3E0MqU/V1xw7cqUvs4EVm36gSWHkC8pV
giwzZ6x8prz5dsorytXPlKkox6WFU2EJNYNCh80GcwoTuM1JKCeFW0HSZ/mmHVx2
bNKGQbq0wB/q3GwYxglzwVhUee1OnaSEwUuZE+3GHYjdt7+VhgJdhvNcKGRF2MYX
02lelDUcS2Dc5sR+gYaqbCRlvNlFxqt5psTec7L4JBwor7aIROX4r7aeFeXxfybr
7sJyXr/580RvQWW6sQZhP9/IacIdy71473p0WUWuckMU40BOzbGzF1p42+R1Br57
EMd3OAz2kGSGDuKCWkNCludsAEEA9cA1AGiFSNsBXh/sdQ67csDR4I2K3W/I+w8l
wcPXgJWJV/xEL1K3a5UoVIBvT1PAT5s0xT8bI9VuCzZEQVx9T2ANWw7tlwDe3CiU
2Gf2bY4KFruSQojyj0ox/NafpJMrgEbTyWDTd2+uIdtzBolmk3toCXUOnxZg7rIF
QFibNYbMLq+yKzG1FPAkjXSnjCkaCXuuH63uybVDUZaUOjg9w9XvKuQLqGYIsO1J
GFX2aJbi5cozWffrWqQm20yO2szXe48infrKTMFBc7KFkwo7d9ZVmtluoLqn4pbC
zae5wcAGfnFQt8CMhM+0psZO4sP+vkc8Rnps/gNrMHEX8XQI/GBa7/G3q9WvgdcM
tsiejKbsBnZUpPHARXrr5sv6Ww3aL+ifIigLfpuVXhjjnk6hYPerrcLb//K44zK9
QiEaCOM6sAsgg6TA78DfGf/ur4+OqJf7u1Uv7pAWV9XualOuzUkhQSjUrhB4czP1
iwDsa5V9r7LLNnxMcGDZq69fcHd7BTlrzKs42Nc4VVTKQoYjNL3FjhtFIyT4xEIw
+bCRbx5ROzDZ1gchqVjkkZ0mOJ1RJ0gt8JqovCFdiPo4w3GwTEeqEHpqxEVp7YfU
heRJLYgN4/phHJhwb28teJov4quJfP0/DNUPb2Z6MrK6yqeFZ7Ywdv6SEWKkZTT7
b7hPUT9Owbo3ZRDy9PtYJMw+yv5DBO/pAbzc/tzZve+NPUgO8OSGAWNuDDBY9qxe
QTBge3CjXomw4RBVRMoRb9CkHTfXyCFIbLtpSWEWODI0Iqoeo/ef4Hi4Zxv27ZXz
3beboszTHt9697aNlCVPRb6JQhtfHrLSXxziep0wLCEct48pI15cCWI9YnY0A3LM
FF6AoYCKq3AIOmjun/NkXwtMUx1INu1DzsPZrcu0D3w4e0llaloKvEl5HnR/zDH3
4N7fM3lQ4YXLXbSuRDEXR1kogAAoBRDxRN7zYP1+skcceVGHwuy0sHdnsThG34tg
0itgAwyeURacXxDGoVhlbl9e/xc5sBu7iHPPKyNlDuKzu1q1KHdo4o1cgyLjrQ2l
RNw92/27jnEMePRWP5IA0LJ3ENqdIb5xbQVDg6ft5m1Rbg9ciFW2eI0rdlmqMqUR
GNAgsA2BpMxDhu36P8E0lBocY4iC3HeeRM1I70D15tgKCPw4aaCelqPHGImIvwe/
KY6N9PRGq8gySbG9jd2E+B44exerOka3XXjVRA3iKihu02OdNkMmJMmF+u0tfyyB
CHBgiVZnD9kEjbK4KpBaJd3N0AhUc0kqDu0tDoxdAy4R4T1QZTUj0EKo2KOHDJD3
jFmopmGl1vLw4UvPrO6vr/PMZMJrqdsSG3EiPBvR64h0JlFP6wF3KcKSwAEIvL0u
JTml2ePbgCioIX+cN3LlE+W5Je2MRZXufzx5Q+hn1rNpYzs/6JZOJSmNBcTiQIYI
BbEYPl+OBlueVFDCKcD83SrjKVeUi03Yz62gHx1N7s23C1QnjpWlWgfFBLuyQSd5
4n1oPXY9z0L7QVvipBKwZDafQk28Ifw464VYLwutbJ+9NZWKF16R4LYlU3O96qtW
Rky6teEJpj/xLR7ms11KNFswJb+Cj4gJ7hJZC/YDHABcb7VCGqMr9YFSzRPybSpa
2LQEoHkocHi4erNq5SJEAn/7Jb5pdd2p+t7cGhILyxBGnaDWb25XxtT96xcUqYyC
25hbWCAAg9po1PYDMnXX4fx3CJT7C3ZJhFxH8E8HSj3o13Bu3jx7uQ1cu9oZIvNq
tW4fpy6zznDgRg4yOr9vBbt0SzuGMhuiGHyPwdpl+T3IB/bZmNQufIkTqTc8RO3N
xytliCkS5tLRxeurLHbHREc/YmsNs87p6Xvvfz7zgDF8opD1w6juVGDkNpmg7qV+
VIJmgT5GwUXroXyortJectXZPaDd4vdDpChwq6LGIjBYvnQMhqtQ/RmzpV4UrCwo
S4aP+/clu+Dg5OQYp8TZboyx+rrU7GaKZBj+G9hvndomy89bNwGN0sTv4n5/rbp1
GOVuBC1OS18nwzr9SY4VWch9LQ/fB6GVmLRiCXKtQqtz9qyV545lJGUbpiz1o9PE
8WCVF/BItVDyKQ2Hmpi7N/+2EdkS4xiJipjn2FPxhGYp3SSegK7yal42dYmr+ly5
GnCYMq/NJljJNeq+YzGmK3hmHaVXTJCS+EA9wjCvRDwfZlwq9hZOBj8zRKKXXgzt
XDEdcz3UScNX/pKntwUS9MV2Rjyrkc6GivoNOta2bczYx06qD4dyt16JzHr5VTVQ
Whno2s3ka6wd+JbHdb6o5UBCZqGv0UKYa8yMTZcXLrZPqxmYsEUpLwxO1ZnT5ljW
YvdCbd0AnafbFG/7slpxXx948Y+q1JCo9ucbARr3COE6xLcsKZUMxeHQvGGTWA5x
vXG9VFPxcFfpcFXXfU4zqZ3DA2LHqsE1ouuas0ASJvkeaheuVmeHbI6Ce38yw4mq
sMTAWqz+6oltEYpJwAPKSIAQ8xH237BGYSUMThLiMxUMW98IXpegye79tq7oD7A7
lluwBYw6trVjPwmUYWO7gJdKkXTJ8qdaLdvBX9M2p8h2kaSypAyLcVq5fV3sqp+6
GgKQK5lkBXNG9k+iJ5R2LG7ZKoWnVG9Fk/IZ1wzKP/of6hUDlDloHVpxfxMEh22F
zc7ldS97vjCpFGKJOWsiBUnXTycvFhk/rke3kFKwPBVanlzPzken1qHig1PxRt7e
zlhXK08WZAG4APRr8ssHN9fTPOHEzjhwlnUKigrtFvWfzP6nsbaqtVA+1C0Z+lfC
queTfl2s3tY1/FtRG8P9HzEdsBcl588YuKsoxaNP8tg5DWIFV1dVdQb+1OW/WQOG
1EK4t2vHJFcMB088L2+sXEuNiq8ZT31P3B63UmPBlwlkCDa5FnXBPrzGwbFLkk7O
iMP6+vF8AE1vq/mO8HNwm6LwPKaQ78nwedlGA/F8rHn7CLQlRb/a2BGXJBD12Wk9
IygeY3FB7wcItAZ7WzViKeXq3kj2uc70+znbYayOIs9FUKA4DEiqsr7xAf5Kx0Ur
60FvjXao/ySpHD2TTKLuVGek3t8in6XJjiTXFNf3hkCBsx7ga2CHFTgO1L0FLOuQ
h/ysozssdzfkuIg9EhhcGvAPEM2+/r+3ghkm+6jkaRntCaycUvWbAM+u6RwKUTq4
ZUiGuMPIUg5yHf+MxNxMV1YNl7XQa+5YGpOAF3Gq9UF4NBlVzFAm+8aFRV37+TCl
3cIqJl02cU4/ccPacVSAokk9Wb41PcyJUm7Hij5tL97WIaMO3dpcYqX+7+kziNkf
VovFtzNSEgVZBdUFIygNsW+BzfxKM79XZzUhB/bZFEvR9+ANclXkFLQwWaYWgu04
XnFtcqp50QF7VZbSx9yY4RYa2aPaqbnUd15r/U1k9fWY9J8NcAjDWPYTJs3PQm7q
xKv8qAwU8FLh9bNxFJfa5C17MiRE4wiRgkzDi/jNFXdbLuOllyyCId/bZPUHTMRE
gADrGWmCsSoAkBDUSXJ2jIXSgpiYcz+FILD5G9+BvqzD7UTBrkGvJBEcYMmzWy/R
wsQrFwR1jxVSss3Na6gMEutJc29WR+VtXm3vdceJQMrAu8yPbFN4njdOEiiqIdnz
ZR5AtHPYiqZzEPFWn0a/zs2iVbtZUvYJ+EXwvkTlnBjP5Yaugztbi/d/2tJuBn3V
knJelzkgEeEkS2SqT3+uf+AadsDOrm8GrW29p/CMfJJp+7YZ7zoHp0UbQ6ShkQFx
djIIM1jSv1PQPTYeDwW5gg9wuSenZkWd8LDFxNc4MjrARvIf7OgU5eW/RT5nR6w3
m0U3BZCC5S61Em7jISzp8UvudZtixjnfMxk5tokt1fuC2hKValn9mbd2B3NZo0ZR
PROoZtCr1ijVWRyC1mYsJBV/xr8eFSb7cxZ5SiZdxbD/WinSYYQjXY/kEQgd4hia
iXA9CGBrZBw2bSRLVacnw6lebWOahmw5vFGH1A7Pp3O4W8/LXWLUm28mRv+boZ83
V95Yzg7h3YC1SbZFQLt840ReAo62sKRckseKTjdRSt94qMAif9b2aK+s1MddbBYC
SJnu0KXVNBNAJQaSS4xjT3+l3v1028ELcRpvUMlMrAb1vQCehJSgDC+A4IyIUPw6
nIHM7uCYDfWW1Z6rz/Kz/zCqAu7dRXIubv4R6N1TGQP/JUOywHSpY6lx6S/PBS/B
76lRGeVX1BLUS7bFYJ9EWa+rPKJx1ZvpxyhsdAI4wJF0PFXNTh38P57eeSkCwHUM
DeB0BXIml4D84LxuOitzSBa3YSp5DKZeiO0WIvvp4dc+oIERbLegQvqSXQkzNHxS
loUxam1ry64i7NwppHeXV6yeK0gaHPqgz7AebG0UB4T/vunJ5cvf1EIqNqSxCa8l
zjx8mcy1SWuzOZpaumqRQbwspzKcR40u7h2QjuTHZ2y249bZEgb5vqItyVpLE08F
uvJ0Nr0oVzwVfYZDQu96byxyZ8Vp9TrFAMdwegJCqWEKiIwUdZwYeKu3P11ij0vd
b5EWIBmIF5YCf3QoW7/zvfDhsQZaTXUqiqS3AfbeMfCIxhdwPaDYv81pqVjzOLEf
7MSFE3ZPIH2BfIjaCSFx1UpwDIARtKLEd5Z61TIHqVN6D7mPwzaaMG4iNkk19a1Z
6cWDgIlVK9E3tEAScbfsDpPcVPhc2Ef21p0VRiW5iGKl0vBkC471LLnBRllVCmH6
MVDuf135EW9IU6ET/hnbQl/NyoOyVSTY4ttXft3oeAuViaiWG9OGdiYdZissj+9e
eg8pJJCkz7LP8jpPmmOnVaK8AKz6hiqbF6xJuDhEshEd9xiXXwfQXC/3hyy2LSCc
ZW3t0UucdGXFkL5U0hgtz/bOmqY3rcoWFAw9EqUZtOJByMUecMAzyFLhyqy9MumX
qDl+Ru/rW1znb9IZj1IDimm+Ph7+7HkfZdnhh6lGZ9TSrYrloSrmdBaO6btaLeBs
/c1irAQr72FY0FnDAhXlr4UbunFTgojmqFF4eAEFWYVJ45xF4999qX8cw47dKkxh
y0NT1lCV76mcUfRkFfI4q4Wk/YqXvzBNZl36RX7jbppFJLij+nhrsrqhAc++koPn
icSQP7UyVZ08jPetdpsUPdpHFforPTF43C7TIUsydIS6xj130W8b1fmdGKA/D5oi
ZSdmVBbIbARGn8uommPNIVC0wapEmW8KP5jp+iJVQ3o3NqFsvli16PtelDsVJmGS
NEctepvpPWiUcfg1rn2VOOY+owBWojiolX9M5IPHSq9JJD4Eb992UCBAgdIbo8Ot
EN3K+na5oFaD/Nxuy1G97xhiWanWrH58zih8jq6kgdtSt1TQNX3OvDGbmg1tkt+P
ym4vKq74ZNORzAkBjy+Dk+r0tE6BKG3mtkFYEv1jqxHgxGu3/5Cd+nKuKI9bjFe1
1afYAvcaMyV2i1ssjU5qnHExlEzpNNgUYErL6U08sFWsccZeLP7XsA3vBvMMAN4Y
4TwwG5uRBKXVk8tCGqqPb8K5lBk6ErSxyAgb3eblGg4elKZ2OE0VkabFTTRX1Nee
xk4x8ePcv0vJhylIwaQ/mEkrP+lFUZVcXC1Aqu6ipL3LvTtGM3GHI1VNcYpvQv8B
w0Pdu9JuypuJm12V2Iuq84TIt6OwS5ujQvbdIwxzX+6jtTu1N+q98quWr5r46Qy7
bLdCI64ZToCPzf7tkuvE0wnxNJXzw9VNZfqmb1ts0c+WKpqTiev3QcR1FZcndbRV
ASJgGhJDVFwf3PDDZKomBdn3DYwkg0qqLx3WWjK9R2MsDr+6t0GjRuXjfVTeb91Y
V213+9Fb7coDvZAH7QrBR19Dm/RgT/uaKQc0X3R0IcaFo9kC8QCZLlhU/kkgpsrz
SY2/fL1dATPyhTLJnvFcFTWHCQZL9BCHA1TmTHzVrQVLPCKL+kCYMQqUTrsEOExe
X04r6KfMbul6Lw2j5duhttKoe2F1SkNPheBG67UorfAppVzN54jLK3C4PWiImwnk
opaW3RVdq/D/640UhO/vMMJ5luQ3/S93w1WyEVNcWJit9HWP1KoxrMKO1st2bWj8
q7pAEm659jTglrBQv0YYacrix/5IwecB2P6SufJQWAS6+sPngx8Ol/fX1cnk3VdB
oG+NxQIQfN7VxnB1rRf6vDejIJFZhMtsyMQn5dfrlgJPNlCMolqXlOBIeSP2D4Tx
PpksxcG9TO95gQ5DyoffyTuVT2i575pLWvupBpKQ/LaxajH6MBVsjuxSqSUjTJ/0
1ZE8SqYvA34igm47ru5BFUB8PcwGzAwm//mlvD6QeEhUMjRk3YeRLj0rza7q8kET
YDFVoKsXfX33TYZhKnJN4RKFqzPDmllOZ9Kq9y1sHayP/oVX8OHIRf1xrhlBTgkJ
31s5/uZM370G2MZFkbnSOtuzlm3yJg2l4f0H1MVS0EMtzFS2wLZypvnpHbvVPfef
0ttWfilmNi8LHicOAwYVHaojqIwDQNcny/BgPxCJsU4Rxvlq0t3pBsxT6oCfXE4r
Jz3FlXWItrbpkMgT70pXU4JSwufj83lpL6WXeZHJlXbbDudhRA8YnWYBmN8ZBb65
Z9QY1CNc+UtgMG77IIqOA9PfclZh1ccLjxBxn8ENFVAkXYuL6HmdpAdvG0CcBRz+
DxLtxysXrVCd3a4opzqlmRQ9GpmHF5ZZcIG2TIyQP3vgBAWUQOOhc4oQpfNL2e1v
sW1VqumfY5weVv86bog+gyc1TwdCAoMW4MRlkDrciHN2eEOcdxTf7F2RWJ9uYLDP
fNeEpDshfdylty1YNrkcxAK60r7fQu+0nSm1Mdcwwphf8tmzJrOdMDZYzf4t/Ow1
mFfMCw0RM0twEDvH3+RG75uFOL3jM8r9oPvkxlC7KwApF5o2etMzUl0zI6+ew8oS
W7/RrVJsyPc4GKwVE3SpgDZ0LhUW+jnwqDsJRfQajaejapLQwDx3MJDwOjbLtBBZ
vMiG6+W1GiPq59bN1UiNg31guSFHgB9vvGbcSgcjRDbIzM74D4SROf4mmsOPAUKf
iWI4koOeXdygK605mTYq24KZL5SIdwzQ7KORJVO5fxpGatk20wmmBLBnsaG49mb0
fDh5SW5QxZrgTzaHnpNhI0z5GJqT31b+irIfMbgMCZz/dD/ybfijf/KbuYKuGMuN
Dlo82yp5uVu8b5Tnl6XcKIcxuwNEFNrMf7bV9nuKuKPQsJZKsj+gSQJhPlxcZu83
cBFNHUQ3M4KbqL0Ehk/yoAH7pUIs2Lc8Y6G0EUrSqLeJIq1nwb7Wk2+67P3VNnm2
IO5S/n7LssBzRdFvzP/dqMAwQZz/L9f/SNDBnmCpYjfoyoXed7YJal41S7lV9AO7
UHRcdGxCEgF/0mFbrjWM96sEfhUi8tD7qCiSR76Bov3PB4OjReNdGcKqSW61fysJ
5L37t6Ynw+HZDNZrMRSfsRiU9UoCStSjQ/gmQt8VnQAMykBBG4cIvjTJEOrMPZn3
9rDNrUQ91mURvydljmXPdIsmPM7k18G4ZE4ILJcojk99Ag1jbs6QQFkZgJBG8EGV
V0kBP3KOeUm7tlQRjjyk+kqtRHZkXDr1rgLzkRbA3vOEWco78HQnvmy63lWvP3e/
zYMpj1RnvVon+w1Id1MJ3KpxuayYqv1yf88HAEhMQAyqw5aNSVPbrix9R3Djh8Tv
KSEiC0hQz8DWS+rWMLjUTI0jhdIaPNaOgOisNZFKovYZvFtyYr5YD9HrquRonFkx
BMU9gRzG1m1x7rbMJPwuqZZX/2P9kosb9jOOjls7J3qagc3Z1iX4VaEbB5K2VcXS
CP7bUerx4s4oHT0+EFecZnaADR/eFIoGjtTy1eC1X9es+XDQ4b5AB7imYj6PWuaa
JhqNmHiOPhfjPWz1y1hx1YhCRkZ+fAW+w4LSsP7QkysQY4UJZR6f7vXLN0EBtf3j
vmlKVj+rULPKtLE1SqBAUw5kX2TLWdfVpeygRx+5VTAdr9CyYHlIVrockrzykfxf
kClVGE+Ke9CDZ12wPT62iS76ZErQDfwVD72uQdezZIQdYKatiFTfVmYoO7QiIhV+
AqeK3FTr0YQsSw0ZDWfczYmewB8t0UGmMcthZj+8Dxbk2NibCJ5C02eThsnDWL52
ZaG3Zq456K/MYnJgSYNOweK1bZQnvFgylFD7+Vt5iewuheq4LowAU8e4eNiJveJ9
tlqxJMEhnTR8AF53lI6f+rD55U2puIMJJzPIJAkkx73HRuAemX5XsMJEOPB9RKsA
7kMVmHoJxeVBdK6E1s8szXSE9zGzbZPfQ0rQRhESvKGAmGbpmIzy2OplbdTZOztM
Vl9HI8yMAWwH5LyWlsswMS53F1SFaq4Cp4oWfY0CBKe+1dd0/VlGufeLqUlCen7l
A8K3ZQQwODr2kcgSTs+eCBEwMDLhCwtJFRGb6vue/hq0am7DzWkzFkrQaD2kTa8Y
Fb3NcYLqA7aj0WbejW+ZjMcrSHqyrmVT4GVyKRr0JYN+Md+u8P+sZ0rHijp+fhBY
UuC251xGbF8oMj3Kh6wKkiVKD0JOd8SHHpkxeNqj+htPiq5XsJKrwR2gqupck2Gp
grsS1GcNCwucFOcIOiOm7AsFMRsG7CZC7hOx1DEsbwvlHFc0dNn0XlnIE1nyCM94
fVchbCqKSPF32jy7aCPuN8Z3WEvq8sJVyNLqbQBoItLAdjVz4nKcxWySkirdQEVo
Ue45ZFYtj8hbkbNCyrGRPob01JQ4bNKbatPI6h+AR5fgaIcWFT9V/AuS4TO9q5SH
MYCRwF9og5xKoIQk+U1SnQvxBGfDKPfEwT84E41hzvOZLN6AdQopPobWgUvDXS4F
y77+NNbMKI+9ciB6tnChiUPa+YWYkCROQSJo9qvDY6IQWvyvCLbTiJW5DWotcwEH
k9pBtzSzWuxA2AW/PFPwor4zF8RAMwPb21k2zwTHjteLpOiFP6DzG8BzDYC4oNzv
bvJZDHSNlw1KSbnU5Ce7VjAzOypXKBMagp0sZB0phKJZLvfgXbydnjxMZkYwh3dA
GmZJ4sDEmcwsfKvhkxc+iaXkutTe2bYPIZOlLBu4uF2LIprQ6LZqCHFnSUWdw8Uj
xvVBpKIzMPzE2iKLwmVOhgaeKPTyUOEaptH23BcaaI93ouwIyYW1HBRX5LYpxZud
xb0Zn3fxeZ6sTooNaaWxWdwDn5/NxQjaoMo2TDghCevzp+4T0KnIL4go5s20jsI8
QAjuw6dnQnRRkkU1F/b1K2B/usbYWy3t/fYUp9/WtWHc17magVSCn3CkaSjaxDpO
NbvGZL+vtvJKJTsFhN3hDHb3Xm70svVmP2JsLeThQR1UeJiVgfFGhgQdYTawHmdz
I9Aad5qbVNvn2JOUZdwEhkr4WO7BC9HNoA+l1/m2+wAmswsCKgAcNtcmWe4Plog9
BLqh6bu7HAp4rwfXryVI5eBZWnmtVwMrnnnyzGLeR6nMbD76w04Xyq9zheIxN2ww
6oRvjd4u0npUlNDRhv8Chfeyi0Ty3cWCas9ZcJYO9gbH5V6CYLVEksRtLf6j47ZX
T1/UEhglJwiRQtCLYgHC7T921OnJKMG+ww+I2YoJQSO4L2ob3IiBuWevGZ5ZS7ux
ZgjOyD23dGz53HcdBEPwMpZ2n8NNuSQ4nb1vZ7nKnjFS0oJvj63f6AiyrvHhoi95
eqAswoa9C+k1S7MypeWJRgjeVP1UqLF6XCU4XBVqUoI/NyFlTv3Nps8FdCJco2zB
qd6O6LDIOJj7No8Gc6/gqDMbiIee2Avw/bZpbEW2noi+fcyMGExiqxeVfoGNWp/G
bkU+8syFovMb23+hQUFnlnfKg0B3U2twRjQ3HsIO4HPDrl8kjw8URTJYm8OGWZKv
ghgrC8Cmmwtmn3L+uFByrLznBXykJ5qIphu5fmGNPUoP2jNvMYiZ//nZLvkRdNbe
2pfTRnlLm79kdr6a3ZjV146NLH0Ydg1BST5R33fcL+Nzt3Z3B4eFNrRlqRSCvHcE
n9Bw9zgf5/pb+zN9qGv3ps/OtAowUAV3kZVqfIUQjIFI2GcqetgbRpjo+1RUIotB
TE8WQXLcMDtomTzWO7Q7q2r2j2M2sZ97JiKQ7z8BNO0F8pd2MMmnLewHnnYlPAdR
UATEmLM2/1N5Rdczhh/Fjy+34Jki9bs2ihy9BXtjXyBf2JQpqhoHDaIeYzEnuFaR
6I9uYFWL9aKZg0AngknksOjo2TyyXGFjAwzermh1VWoFcmgTVdzCME2MRk8PycGA
Jasy1e00gDkKu/iCZoekQuHibwshg9rRnWgUw97fdb5g+0XU6/uwpxrw7m2fvIz0
gDslbKGXnIKZJtYiYuj636Uf6rUTAMbhiKlwSAW+GyTCeJ02yL3deHBeX2wGb5dR
433t1dFN4W1nWHzj44wCol5GCTB/UtjHl5q36FwY4uDmZ+O42Wf30cfHOH8cbH44
yIegn125iYWV47ycpDHim++4VHCJX7JNGzevg3X8Gw9NyK1jK64hD2uzquXzU6OR
J7ecoQHb2pIn4BCTEj0+m3c1IvvNgyj7zQzmS8J2yog/7YusbXKziXeoOVtLmjg+
y4IvpZYcp9y3lXlTEqeBEBiJHP4bwpkDYGYx/aip7+kavAR9o2jZBIWcm1CRtlqW
O2e675Gb7tdsNRRTbSb8uptUM/QaxGZ+Ntk1aQH1Kr3rvjm3lvQz2q+S/o2jluyV
aozC/0fCrBRsiGu00Xi+JUxcZWg0VLs/6cd9ETc+fuyIsLlqN0aLrTO7TOj1//O/
ryeqEQsYGJanIzGrs+kgNuDlBuVQsuVrLuaOesnH/HIdFBuX0PjVO/YsuX1P4pbw
/Sgc6om0NLVAlbRiY2s3rncMZFEAya5qRTkHGHqNbF3957DulQpHgbRRriYWgZ4Z
oRgJco4ZI4UEUSMqps6X3OEdTB0QmR2TeCnwYgP3YcbbzJfQ1zx86200YdHZDzKW
jt198+AQQF3UZvTJzUEPEHfNzPHL4aoIBr2YeYZUE8JZClbrUmUQr//VCLFCxAEv
CnJ4OikdGmOyd4W/uF4iRB9gVA8LVvmaAb2Xa2j9fsNXPYj1Mcyxh1wLHzvqN5uM
z1eDaZ2snufBnRWkoo8XCusMgjeNAikD8Bjo/Z20/YG6Z+wSjqBD9tqptqOBC4dU
qDCfH14Aj/SpM5AJC3ciWjjYgoN0JhOFhLjzKE0sM2OL4Zh8qFJGnZaZpFBnkt6O
sqSz/6OGFBJe4/ZhJ7wuDalepKPU8EXxEXu08wvku9bBBA58nwlMmvIcjacwZrlU
8PRf29jqdmI+Ecw7hjNB8OjY8sqX8qG8/RAzdLKzwD/EXizYmRbvLUw2AvXGxoKy
PR5cSjvnAvfM7IUbj6zWWscs/fu0nJn/DDNuhDKyK7wIVhdeVkrF87hxfTeeEOKr
//B99Jbl1CrR3v80t+2eKD2AclO6kf1lVGr2KJIgVfVJn+H/sonsrnBnfRhUV0yC
bZ7YfK5RI3JqwVYcCzt8EzTE3PQwTIwx7Lvf1VZXIzS6Ol8enPdOEH6IUs7tl+Ae
gMtPkOIoW4sspHeR9Ghb5c040doCXn8pu5C13Je1eSBwWa6Ech2jiyPAR5jf42Fu
kbrXWI9/xzfvO/7Oz6B355GTsD91DY0cZRxIrR2KQ0tRn9PYsCudufSi/GKY/RQD
QdLHJHDEyITRxv3schLhEKqM4Ym9nt/8NyCFXIC4wZwcQGlK0U9i44pEU9VtXuqN
aj4F2r71xLS7ZlYahlGQ8L+5qPdp89sA4nCafSFJzxYaYUkBDoFjw7EOboJHoYcN
IsNqcHEI2GlgP+6c9e4+x8VaQ+9H68LtXur2yRacl0iPARD6/fLLSKErnVb7Bi7A
PbgYKZZEh0ZODVuhJSZumIrwDny8XV2T4X0dJLrR86QuZGEYH2zwQAV56N4RxSGh
OuAzpOsRM0jxgeJwdMXrirybI45MSVj75CuQ9MFXYAkT4thTdp2q2pr3RUC1w58R
w/qTfHxLep7+MxDhpVBm7XZgFgVXEsUUyMXDmvcVonEyx2j+xqEQyqHQxKExDKSS
2j4/nSZVaeFvF/l29hOdMs/R0D860WfQtMZRxJ7FLdB3weevUoLauNs/qrW6jqQH
G02pXqDm2dJ+yGGcxgMTAIt5cr1/JjshXg92OO/xxTe6h+s9+qHRqKExfZWHld0e
wQbB7Gz06OdozwEnNvzu9S2FSPAHHNW8cb5GGdcOCdl41Tj3J9fBmOypZKZucM7X
pO0zxFxkWvi/NoVsG81iULbzKWooBsJikmTU8ep/WzyRGxbSU/dt0Pm1CDKRK/AW
NBLvsE0EvPWmiEh8imn4Br8ggfXuWT4/SgKtlo/k0j3h0OwfXW5gTTmTU8JqGiBY
PL+0VXPXtY6w4IeP9gP5iPLSj359H0RFr90WT3iO1vUYaMef81xBjM4OojeHx4O4
mvKc8Tfw9XhbB6YOMZnVKXzCfjxxgzrXJrerdtv7owsIC8/7WujZcacZaKEERWIT
1Y/2yl5uzEH5CVlNqAAiQsDaATAQXo5FsEa5mQw4jjncknomXWa/d+HUhkCovKAs
/SoYZa6+iDP9L0Xif8/QgAF+qW2M6tHh5G2RLPPyTQzrNmR08YaTkm3+tdDEz+1W
tJEzg5ssfdvSbi7TbPMjpsFBcv7UqudFdaIZaF/Aq04ETyjDwkVN0LLpYjF/Hn4+
yLgR+uQ8g3/3fh1bUnZb7Mg8KXeHTG62MabxzZPq6Ow2aENYbvwfW+eSEmonK3vP
JuA/6sN5dG/888BSsUHKURdTPFvuKgqMvgbRVA67uxTXp7SX5QzJFdoe8te34Xul
IDjiZ+m5ECgSJFRcGXLNGieGuFsfUhKSqOaU5drfrESLL+aupJA+mkooI5cqdHLu
sKE4HXW6amU28kwwWH9YV1cmvULN/hxgabgFrAThKc7YoEgAD/Wgf1bdI+Gn61JC
6XmP6IiMAQ1rI7BaI6tsQVc2bK6Fi0ZSEgVE8zPFizZpjv1eTRC8se8+NVc4mMwW
DJuAGt594S3z0F1MmJCWl0qq/fS2gQq7J2VKDTfzB21uRPbNOTg4XHvGfTGszzB+
ddyxjcJMHpcm4V8dU8xm66uOfrELfFuBXDDGXW1WGi6OvW2jvU9y/uRFmlk5JdGV
13+mzTCrM3iaJH5wdOYkd/7cXZxQHqehlnm9Vq87+BQe8WAlexhBcGd6bmcfcHBP
JXJ2AULSUJkEprZJMz2Iv/CbqdS7uLJoS9oH5bEdG91mNTRYZMGoitJcjP4Pwf1/
FmbPEEQDhY8FpUa/jSi1usP5USXcpS1OcZCSsSbQxpBztTanzZej2ZAYeJ49j/vN
LJ27IP3cpPnqZPZ1iKplvxRIlx5zA8QQCcnkhKNNsEK5ZKfMjIPdEWN7AqbAAHy3
zeT11u18Ekb+Zfc7Gynou0EUTdTyo1c8nYK326YUmGaOsB/S5H0JVI7tm0NncQU+
qN6gjr+BUR68aPdOXdYbyjRFRANAY2O4/I22aR8MslWNyJdNYx/pB9wJ2R7MWvsw
ePNPTwFzgM1xw1KZkiZYFKdC9E2FBEE6oPlM47kjej5cMrqQslGAEajLG4BhrDfM
eOs9COvDVNvnDIWxv7enJU1kzMjeoggAFPS/KTfmyl6nZ61WeDvcoUO/obsHDoML
CtTHp4H8XyZ0LSKO0dJ+P+jYWiZ/psUfm6qDP8cMjlMaa56mSRQSQDGn2xW0+wH+
UcE97LsUaKRhOAIY8DumtVxs6k+EsYpxkEfLHA5wdodl/ReQkf6fCVz8Onpy83y1
TzBaQyscdLTzIAa2kW/HNq8KhJXc52A9pto+1tJfpKHpAh+iWsx5HQUYXS3+TUe1
OKjB+ZtFtN2G6eWSF/xSx2tbmPtwaj1NvVgT+ugPsoykgAbODRafkTFUInW+sy0v
QuaE927HFXFA8epThfKFMwKa1pW4vZ85Y7XdOrXMXWELQ7GQGd6FI/S7cpKL7tOi
TqZGf2mvNKYyD6o3c5gXdSvW3MMhxKKGu+V2tg2dZRUknWkvkTxMOZjEo+fpGSl6
OlKyrouTjISVqWeEIa4tJMTGfaCg8JQ/bcnKCF/ioDKl1bvPBH6OXcPv9KPyJ1zx
Fv4vfk4RnYtrRmx+0/7wVj7Khng69YRDfy5aOM93gicsMfqNCSQqiaDWcy5qYWT3
GARek5nHugzpgdNz/01X2eIrBYubQk6rNHmhmnb/yurm06QWunt5XZr3aARD+uKE
+BqbURtqd1iOuAhWKS6h/Dp2kGXASma5ztcRwOEAV4QvooOWCFHGI4SM3G5yzpAa
xpbSxNCJs8kCDqbipPnpT8luOWPSfKBXVUI961Hsc0ndeOeKgrJNjkpfa2z9xNi8
NfqI2N+Zl++24mku+g8aHSGOeXAl5Nhy6JLtJ4Mbmob9N38U5By+7QA83facDuoU
wBjHxQ+K9PhK7ti7iK5wo35/UCrGO33o+FLF38QgsGFKVb437E9mvVn4ZNtA6zTC
Q7Bre48UK1AKngkrD5W+HE29qRSyk3Q/wHjUNPknjVPkBVae2tzjSXvEzCArtVsH
c9DjgShnucsfvQvqaJA2P7IKjb0LG3Lk2gCnAdqBapUm64eJMHEddY0LuVMFS17p
Noo6UyxEGi8NWW/RP+O/RTnOkmy2hkXNILEWKoYIN+aVhAfefthUNfgW6/2Sg3O3
0kbUGaVmVzOB3gn/GkrcIOw+7o9KiP4H9VuxjbakU2MHI7yOodjEyO5dNmYknmXV
sJshlgG1R+Fh+v0Fm11FqxgCs4Q27zj3CBqujWTKewWVV4O6852pWGvySDdEWkB7
Q/kWqymDqKeEjgQ6eu0CzjXyjFutLMfJDnpQX9dOe/s5fnRi28sOl4vQf/lD1EvS
iuYDLGTCFHp0dJLdZ+VGKV9ycQ4Oeq6gEYsepPBIwiRDrxMoxJ82EoK4Miwl/EYC
KgbyOW/NwvLpjIInsi+0fwx9FDmp7GhnojBIK6Sufk6dTl2dow2+oM8PPSPBzTjw
zxblFoXkee6MNB+ESy9ZFIaIdCQr2mrpw2JPgmZSG42k2boNAQYnmmUqOS31XxJU
u+TyGR7jgFNhiJNG1dLmAKPTxUD25JD7gsA/l5kcIpPX1FdL1xkBgCstM9A96h4j
7kVvmRJbuCrRSp5DCfG0M3yCSyF9//pMJEdJXKF2WWcFTrO2Retl7Cy4WJPip3hR
Xj0G4J2EWYRMuRcsPHrDKO2oglVGb0BxpV83lAzaxnxYBZ4mHf0n00ndOF2jj7Ko
lt1JrMI0rLXulGTEnc6pN5doytifM3FXeF3S6VWAuZ7B5o6d84YYw7md6C4t/j4M
nSUPI/4oiomlEruo80Ix3C0z9USuTXhRD5JYP+e9CyIryvce2glR98K/epIDzq6H
5JmG7yMUdGQskoxjgSAPfEChEJZre0OFir2Dd+MBpYqCXfNu9vah6irUqsQGmY0A
XDBd36kZ/0SAF2JMSC5quHF6E9R7cXEEnShf0cQAjyz8M54CYv3Y/GBpbtoEjobn
mwLQ1jaSHghv/8faZy8yGH76JJ6tARm9Fbh1LjF/w22MMpyNttW2FMqlR4Y13W/4
XrH9Zh3dSeGSnbuigd4WX6wFz6zJvewF4i2VGBs2Ct7Ajvpa22TgwEiR4fKrxQrJ
b06bOPmlbeSgtekLOGK9D6NjhQhcBlDL0zjKtgAYTBIQQnlFtlLIiPVSnm/prHnK
l6tHwYmdwZppeQhmwPh4aZ2ve2UMeCup14IJhrRKzKE3XXIcBYzUaIHNBaj3XVGv
+9VdNmgFETb2II9D/i/JnSuWAjuBQzTiRCPO4kIuDNiDab/sn9qmMDteqPo628i+
S1zi7BG35cvaIbHjfxDbPh6y/aRtJy2wD9sgcBzor/lxusEBxSD0bKbQC/BqaPgw
lioWJDs7jHIdGSwVffmNPU8JndELjT7HvWC0MyG6QrL6x0teGVqnCoADzUv074Yt
6CMloynkdCBPppQ8fmt4C4vRZep39b1ERGWOp+InlU7O3ACeX6yNta/W7BvkC+6m
47Ql+ridSHQ2x0nE6HutZu59LSAKHGG1f6L/BfxQ4q9X41SwDoxDIxzgcKS9glwE
DvRk+a9XAXMy4wENEAfhPXSdOeGpcRoiYBXBsOcTaH8Kmfd/7MeUs01bH0cF3tQ5
CUfvlFFtUQ6z8QAWqEKCCL6aoHOHoQODp5vnBwB/NG893LK6OZ29muAqG78hi3th
ud1Ch9ueDbyyYKUOW9R8JNvkYopnecR7tduC9I+XlE60xUmJESOHQnpjlxP6audo
NMa8hORg9tcZe378fAVsEFBDKGpLwy0G6ysGXHO2+TU41R3enRT31/YOYaTdNp2F
O6K5qTkFA61lfb/mm8dcvOPmnKSrmDTkdNs69BKoW1lhUctLaufB2hpQlLH6ewIs
u8uIsJ6Mf0YmGJg5P4qciq+6mkwBId1Y/55ykyII8ylE0ew1VgGMdXdZ7+3vFKjG
97TOeqyhrP+V8K5TFDSwZp0BTKn8N+nDRt1uaqdYLc3RdsqhojJ/NdQRhqo51JyA
ZEdMwR83h0s5iO74W8O9UAlLmHt9Q3tnB71ceQWzTsyRKqe4EyPcNqxPcHdXSV1z
Z77xXWHp7l71JGxKbXlpLpzGFe++0qpPmTRdhncgdDUI6irohxCKt1gw9xXCmLGO
JjIX0evypqBUaxYfK9iv37C4p+mu7/f5v5iqkw4YNVIirMEorzpWt7daQKhrs1WR
tWaGd0Jk5ijmf10EQPspfKw2MCZLs6UVWlCUP6gar/FU+HMb4QH6aBQ0FFvvIyp4
i0knneMT3YY/CZpxBrSr1yDZpYlGBkwCaCLnapya3PuFWL+emXdh5q2/EsM4s0UV
9XxMN3gzbCWMjv2mVamI4FW9GeiLiR0Mo5CIH4JxtvLATao3VUR054N1cAIl6dGz
+9k5EubMdT7S2oasvtU1ZuViezfEJ8tOC74K5WBEVvRafa8FXVEdj1tv6p+/Yf18
BafRmCX81mZ9shVtULkJmYVw6RP6ikzC/g0KOEfx6Nm/1p8Zkh8mduX0tc3yKSOG
n5/3H9PtDf882aiP8FPBNugGw2tD86jk9leqYNOuCc3FhCPssFtfzlxOxQ0TK7I4
U8LIXUjQ3aKfh5aRqy142cdZPJ8MXBU7Vk2yj6sDbQ+550TxWu9VLkUKqmsryiMN
MsmrQcFFNUxU0KrwIoZ3RQ7qadoMzdFw+PHSzCyHdfGVGe7VGGYqZl86HyeP8rwC
mzGeF03H7HibKRFMJe5hkXukhQPg0me8lED9e3GnhaZ8pghEYNxt3raYx4zGdQRJ
dEnowTfND3w6AKqKUlWyz8ctDRcTUIC9IxjlPvA1jf2SqxoAivL6ByCCxHl1gkAU
ll54TIlOPbZoCM6d4FsagYy95IMLnG0wta51CHEfwCNduLk2DOxOghFyejFrigf9
E8UpWJlP9l65Xyj76Q4M6m0Uj5dONDQHt1TotmQ5WpLdaJQ+qmzrzKQOZBybFmXl
PkMA2t+16HJqfzw+/C+wGUeP5NcF9H8Mk6hlLslAj1wV7FoLFYHk58TMmNJiM7Kh
Jj2o+7e7JOw7C9XkbX47+Sfd+7QpMNWkbcBk521hmY4Fv98JoxqKX41B5FJqlTQR
C6F0i8VPiXqeAm3Shf56qFNsiWxqYM4Ti+nwPrDnBt2/z8eMlY2M/W/3rnR9BW/l
QDqpHngK/wCVUMOKX2E0VQTma+YtTe6Pstoii74ShR4NT83BJB2BesBKffAytynb
CI0egXpFZOQ4vlP+t/fVtdHjTKxV6cWY/HgM9M/EmCtV4ffl25MQ9fxCg7qMSCK0
WSLujmIlYHE/5UAcosmr0yUw656udeeaZzIfAsc+6W1HnvlHHeQ65ikjlWV1CJKY
007ViLa67jd7RAlUMfopXP2X4tYuqHDHWtxw37igaGyZIgZOH0XfpQM4LDABXwwY
W5okpeOR6RX+RfmtzVshRAPi2cfDJMpo5DKz0mdTIkzqgPw8DPog0erZNYuN4d1C
BkBKX+eVyjpB84/QTsgQmsIe+0ffyHEZke2WK6oTBPSDGLf0pPLu5T3770FYfJcZ
lk9VqP9IdTNea1Jdjs9qhz8TS6nR+Ghv6215nlR6prdGzBFfrVN0qNKOwKi91Ep3
T6AbbHjqiE7jjBjAg1eUIvePG42+CFq7hDCBNcAqAIbpMYfJTnIo1BPMWXqvofL8
un96FBeFP2Du2AQAsuOQ2Ngu3PuONGx9PUDPBU7SrkueL3/TJL9EtBXP6um3ErOv
5h7h1yiB2GWGTqexZeAqzI4FP06oXSdx2WMBR67zg6EdRVA+NOoFzvD4U04CGUn8
/bPwXKkJ8kCLVesbQJNpYvUTE0AyTqqqtR9BCNeLSoW53CB8nZSp9oIXuzkD7ILl
FMI2E71vlk1Y5xh87+u/tzgs2kJv+SREFZdX9hXjxGiVd1QYypGVk4oJ1r7OVRVP
rIHq/9vC1aq8kriqwlc0SBPQ9/BcYbUW32rlTAVrRY8CTkXEnWOq3M7Fkl011aR/
UoPA8MZ2juNiDyJdyeM8E37E9wSpvowzvJGg9hGUtIMVqBBZrPmnnoc2IYF5Xlu2
F5iKg3M4osFOpQxy9ol/1Zm9cz5eKACxu+BtUqeFyEeBh4OXSzXn2pQELoyXPHoU
Se0VLLUY6uLTlBGm6eQjbFp18VTfKuxPjP68p34BQ1/ZLv9r6EMeQ+IXMrisK9pg
kLSvuhmuUI2r7A9h0FNNbhbDWWRs5jeV0kx21HqP8UGEm6Ndd57M7MiWvGIWpT0G
hZAJUhQob32t8Rx5nJf3b0q6ONYfAYBZrK3UUfC6+R0qEjuovrRzvZptiiQ7XHYA
BKSiU560scuDf05H77lwERPYx3RT92G7vx4VPST4QBDzHjvNan6LnRvQPbdYwcFP
GfJ8Ji3vhIi9qcIl4aIjeaZbn6gKzrzLCEzzGdktnkyOVXEWU4Jrl9bAOQZqCjzC
ubhZ4Utya8jzFAb3KxlF3ICSZq3qn+4s2czrVnjyX0J7nm/pKBsw0c9llG5W4qpP
AiqNitC9v5U+bTeAoUOkV2yvCUvT0+0zPQLCyub6hmvtXiIxdzWsvsA4uBmzZCpa
om+M44CGdxNnIEwi/oYkTI9THYvohVOxtiuU2JnuYFDbDJW6lauV78L80qEuGB1M
KjO6WYMLVK27Ny+B4t3fnUcR3dCK5jAP+QGzyXx+JYm9p5nRNK0sRB11DinLKq35
K68qjEYHtizh/par9qAKBUNEkqPqfO5Iub42Sd/AZulbFFAhmC2Xd4fsK4VlEqvL
I/tcIN7BKjnXlaEqfCAN0r8BtYyPXI0h3V9Jtv28PKAz82hiGqbmP0n56gA1cZSd
wOXhgnd6b7ysWM8QRRM2sWmi/n661MprWrkFlV4VwEI4G5X95Gx7a1rTXCtZrJqM
4xhkvI16lfb7mAE99U0dbsi2Y2CPr7yLub8PruO6aBi+YhDMv3g7yE4pPufLJh2E
w0ecM5FO4ndaFlT/ZCwNi8NwxG5GmCbtKYDVvTvtU8ApsumltI5g8Wv2gGMuVqwE
NwP7fxBf2Bj4jksUkgWDNGw4r2A+4Jb8hHr7P00khTf2PYMuVsEs6uKVYvT4F5mk
RntR5VY6DxMI1sincC6kXkkOBprB8+sxwj4Dqa/jwJRGyRi/Acbs2E54K98Rv8/d
y/d6rNfFbBMvmO/Icea4JRWuGliBPifz8kS9f4VvP2rpbWad5pfTTph3g6o5LyuH
dKboIoDocQSahI2oivhjmd1ywvNgV20gMb/sELyFCYc/Fo7R+ScTCfm6k7F5JUX2
GW6cRPVbkbOZtN7yEtLWFLMxe26w8PKkvHPQsJQ60wbCz/3We6FeBSZ1FI8YUSJ9
gX8AXewlrEKEMjbCZxjVst3pCUW7n5QjV0pDMnAUT7OChjDXC0ixe173ukzsOHZR
l8YvoJGGIRGjiYjC8zLgXltAMmmxQVnCgYtCkIcQ3FBw9HFN5is7s6fyXd1sATAQ
OVu7yqUN/Hc2ZishVWbY0z+vpsa5QsV6o1StUMxMFqfmYogg04GJ9NQehj1zmPtP
15QIjqHka5jwTh0Bgmd4QA1nnDLwGXgwaM7Q6GuUbEWnuImMn+wx0JowOZVkQqMb
Qh2MoI9wm9+jhqZBvo9tJ1Q6PMzyNDc/fuV/VpLPPEBHB6LJBLgtyAuFfccTREa1
a2eeRKD2PG3vqA9IF/4jmibAYnRYP/IqyZOzjucBmRAhxVgaWHJCN98oLTpmaCHn
r6DY/mNYqNTMpO4FLBLlaEFHa3VsUXPejYTdng3mK6VRcY/AsdJl+WNfxbSwbG4Q
awLWmCtUUBISdagwNJe369tqw5G3gsEkmKGTVI7E5SqysY9Io71C5In1Cy86Jn63
o8momxsvwSY4mMYjNKelloui3+FbO4w2xZODjX1Q9y2AThbdY64cZ2LisctdqOFA
mi0rrM04YNYe4oeLUuijEgalFpPXylk6RUchKZbZzw773WCRElmQN2DZBJDarAkb
Y+7CTaolOyy0D5Cj3mc9SAvxHdRUAE4G5Mf44SqJSnR+9ALhM/qfCkIhcb8zaRQh
agJV1A+TlEjodhZ/OuGa++NY839Jyq2SRTltRIRNjtufOdgtHY6wshFBzeg8ehsY
6SF5txT1FUYtVTvsiKpUvzQ3bEo0ShcEKhL7EiyZJc/PTbVjPWJjaSC6gfDSyyoV
krrTjNyCH5mpg8uTaLGBUTrxUK88EPzLcPT4OwU27tq7aosk7RY5tDQqlHPrW4Tv
DuKl3qZtXXRgR49h1sJWQRvZQ/Ew1Vl5zOr4274QFA5DSEsimjs5VCiG4g23rbxg
7NsngY3bG+cb++UJpt15ckKkMJgn4gjerGxzcQfu6ToupNgH9fXxaGEuYZcKoFxX
4a/hDQ8gKZyRPCpEHiXj2zG5GWBapDQGil8JPN0zU5teg+CdOUZeujdNeEshiwMB
WmMxMOP/LDq8+DFvA20pDeIYU1gWynz+twSF+av45YAv9uhkYB+Rjqh8St3ZSyKr
/DW+dj4ohV6dnM7Bl7DVI3FoDynqYR/CIOhgRmZueLVVJFAkFXe7Pwe31D3P69iV
JbHC8t+7RCMXEfQCKcZmkdswf1jzxuKFTgEbE9YRiPncOK3xOYoNV3qFWFkpIsWK
UYnnnZSfaR8CnrzB0RWten/MxUSmH+gUS/tKk4ndqzMmkIY6/cVjoR5REqW9m8J2
Hx/PWZ/wiYnkxzisjN1QrCkbk/vpVLt++zAmGxDEMlFBoJyJVY9IjvpthnNJsjsR
8uNwJHQ7KJE9b7OxI1VPKbD+Nk3Tl9wojvKoroT7Xajwtj78tteHp6CtB0Cs5qeC
ZQONcxSyHYAL6NJJkVjfJByZq4+042CuvEDXXJoJGQw7kD98Yci/4JL3VFlZZpsE
fGKSSODERMiXRU26wa9Rc3/oq/K/7JJhWLJFAbiNIMrBigxx+SyWGxgHF1mCC94q
pTqkuKMXe6VbdCtpem+kGS/nG5jHgRGB1cNIMMyreL3X+ctxOKxTQwiNS8AUXdXa
Dw5/Bs5CB5JtlTdr+FrRWluf38c+7Y+Y9Pr75buHXtTHK4qsRcjQThin+xDHu13p
95wxTbGwJPjKzMwQ9dOUqwsY3GbT+e85lYLTPthJsVl7oRtTyKQQZcTmZe2BiDot
k0A35EAi0pjU3kEf9iOEiizKJJBHzE+vQ8ntARgORN642Y7+Hb0swANbu+B59sKw
FyRY6DoprN8AwP2AbKMX9UhjxECWw6WqSuy1N4q5j9zH8hqBDf5cJEACvfs4iK45
EzhIWKdzm7nBJnieBolaZn20sMvvmeW/i22pypfqYY4Y8kEzaR/DBw/7rkX7b0Ni
fQrwdp//9HVCqHs4Hg/sb8v2bSh3PcqzNbYG38RatRsIhGSwGfZBT64XavIbeZ2X
zgydo5OeMDoqGmhDQYsUZqlIYpMM6X0GPK1PeSwds8RMILsSxBEyfVRKLo/t/Auw
eckxVSNfuQmR2kUjjOcv12LHCwflTbTDV0PRlZK0shvpOkVmfzKFlzn8Kfa+w0u/
K7eVisy0QXlFysbhmvaOVypp28NwZfJ4Js2HG5QHa2ofzH8xEG6GXLP+e8A9yhIR
Tml5EMtSB7cQ+SbSL2//DHqgYbfq8Gcy6HhFVAGnHbGR2hRBSeN4yx3YWxWTACoO
U5KqlGHjJp7YEcI9IXDXz59qpZ6HBXZgN71X8LHGu1nQzOo23jZgKyBfgyRNdgm4
frF4syOBP4UQogO4bwQOoD6180CaEhoOHlN8s69X429595sjiKusIFuspIoS2IVQ
QnrfHFpxBp0/P2ydf7CxvIrC/ExRjoD7uqLZ0a3LIayy4/0YPSQNckqvxVKKEtEr
8KQwTBQgXGpt6KwYO0KS3c9KB3h2m5iMd2wX0dy0P0alZ6A1EUJsCfJFHKGhR404
T3qtM1St7TrbmKxYOtZtmESzbxGnyXNlu+d4KkZo3zXeNr/Uk91UUJ3N4VM+lVdn
WERDuS7O9F//MYS/JpTlJpTu7Fs5jm2eyvUEyZlfFpilCyvISKFx8Tb74aUO6qcZ
wz3Uz5g9GYjKwdA0UluNKsHKC9Z3hHDFRSzmRU7ig6cIjZv6N4n4AGDywhmGtcoC
OXkFOhiaR0pishxjm+mwHul7OrRpVtCgeOYuuMtuYD4Yw0DeRQNIF3JE/abrM0T6
NK3FUuxUpLH0/vPM1bWwxzRmMX6sql/XR8mhojBYwxU+1RUM+fD8uVq4RTiANjZv
vubpbwzb+AYtqFAKVjX++ADj8n0he6LaaJL1xgvEFS1Tkf8/2tcIP//sKk2UJKhE
hw8pVmADdScX46e6opOuaw7V9usTH3aMA7QSl553zI8eDdig3l/CqXDvz1uNEDm0
qjHEYdW6W02aNhAY8U29ubVjdkY18Bf9CNyT2mkYbFopT7Tmn9Cvob2IDqnE9po6
V08Z7JR2QqIkQi83LAJyh2Hz5V1/ZV4G+lRVokV9zy16yt03BPvJ8pHVcR3rSv+Z
Ld5yFH2HzzcGXhGsq3kw2MVProK63zCIm8EM+G9PndZWV4755zwTQYonPIRg8i3Y
9DnU4gmkYAdvDrUQ7jLZP5vzQVuxh3+IZ4F/0Q4+XXOpbu2cjeB7jxVfGGJ50iyn
qxOgxu7Yb0XygtXwhQyFjkAZxEQVDo5F6kMJoh966g8VTc8Ys/esdTE1rFEVR5Q+
WM6ZN/ZLYllNB39fisd4TyIVCy/2rT6WGy+y2xdIBgvzSIDTlLKyFhlHJ/zy8npS
aYSKQSVfFJIvK/QWgIywpaNcjCO+pMhsOzyyjD4fNFhjOfHI1fARBE6id1fs3qoB
kLQ7wxkj7QbkUQTQwDzoXU6EU48xorlT/LN86vcEFSh65eECQIfLKCtRxLQIkMS8
k3q2aa/tXOYk12QWtX7bZPB5z3D+PsuvV6JEarVLaCa6OAqL6SfHGU8d7jsFH9N5
yJNBj3Cp2IU5OeEQ2DMppYJDHlBNcvETsSpUsCT0yNBAnPNwgmWGNxWL80HKh+ia
4VnRRntLnaAkIZjLmJo7NsdKOPZZiReikVF0JoeGtNG00vzf6A4J0FoUqPnfqbhc
A9AFSa62/dHBtErBgTb8tuBC6FYtfPhSgmCaWIr2lMNEeoUDWzcrt18EJFUwaAcH
rWm88iCZlOanLECGbWXAuPCCakzj9l1fz1YK2g+VavzYzEOg1owtLD1gQe2ByxyB
V87Icdf257s4yFHQFjFTpce9grJFs5wzlsMZYgPofJ3K1ZQCA9+PEuF1B2iXk+Hw
pzK0QDsr9KE/av6GCsnR2Lu2HGlsCfTSWGGZLhGLHWWwsGFvtB0R9tjKdp/Cmj8B
k1goZd6EUZWQpvjyCFdrS081z1EQBxmWkY5uSMsy5wxkuOyejHGfwx1az9YqR+8k
lMB41sATqZmG/U43BmKJ9KX8KRLjoUm8B04g7ekcidQVct5aD369+Gj9RO+kjL0A
t02ZegH9JANCZqfnpxEYjRoHpfD131O3gi9J8HK8AiJxiNCo3IsAp6YnXTcY6gg8
4edzCZr15VYoiCKB3HhYE0pt6h0kbH4QzCs0p5NOqq1SU1uCGfSh4QuR+dsFf2Ry
ZTMRyfAGwFN83DWOoAyGzN40eIV/wZPycKdfZU9TFcTzGiRsEVZ4yADCRa/C31J0
8zJPMwaycAUNA+i3SKb3/uss4QK33M4PHzzsYcShMbyQM0zd0DWpynddj9E6lNmm
3PBLk//WJ85UcE2ayWR7qKWeNdAQt0blyEJZwyg8/Fww4YmaVa3ihpJoEM6DYdtH
c1yrdB/PD0t02ijzesDW9DiEKWPD1K21NVDdmOey49+gYOnOLLhzwhucoQmreaL1
4sJxLwOfXxutO1AQT6ZkGzzW/zxsmbseq60VjA0OIVuTRNW6BbVMOm2flgHbVXDP
MwC/beGkQGqz58g6EURzXBeNw+dyCHW/uuFNqhyoi6QZtuOqP4iUOFto//3EC2XD
n5WTrZaYLWOwkhVz7duTuflfVuDCrO2pthrjBCDQasCe+3uCzqxdE7cWd8uGtH8s
5WqTj0GlZj6Z1K6Mw0d6H0yUpu+M6Jmy3cBqL39FIKEdxXPCzLiVvUkBQEpp82zd
4h5kft8O25HyioPeZsigp4QM/PmaDl/MX5NQoP8xlXPbKl6i+sEaoN4AqDxCeSdr
L0KvpksOsehsTRNyzrvVKeAC94R1puyPACxWgxO8AoXd55jGCUrj6H8fyoUeDXwU
OIW5qzuYf42gUHQ2/XUHIPx1NUADATmQ55Fnv++j0eXgKqXIQ7NlegyEmouvQT2j
ixFRCP4RQalfUv0C1Dvu18mel1lexPD0EUnwC2dAgOpoxIUR66EQgT/jYZcAC9oy
QNwQdpdPZ+SsjOdRRjI/cQzfbaa4ihvWckr4tqP/AoYmhTRD2qt2iwHQCLWY4Jnk
mRNLH80oZaNWEDzm3rJ8hzejdfWaiqJoephKWo3kZOWnzydSgU2Y74VkTc7059wM
OJE66f4xxZLVAVGivtDH1sD9YaLXpYhfJgCpDsf+z3Qjiz1r1D4VBThpsgZlq3Jj
cj44o60tQ/hxpPUENV9VQOYtV1Z+lFGeGQE1MWsIRpZexsNPUGdrqapsJlHHYE/z
gct9HzAUsC/D3vgeNHq0CbqOBW4UX+3Lke2/g6P1kTM7XMgc/2CWAMDEN+upoOqL
mihKK+r1qCYeswc5kjgSLfBM+qFC7N/zu/C2Qold/rG88LJO/KiEiHRo/R6XPFNT
KfdrMKosBbHz5UzDmVbhqpS7UQXtH0KcZwepBIXfAor9TbrnsS/Jg+6SvMl7bWNO
8Aqx0I96FhSDZo3EYqsUGI4V0xCJeURpGpQVh4/ZD2dmlNN4309nTrWEKdgmpxY2
1uwimXCeaIDfxGwnOTvLGNjEigVvmJnLUqHIsOJ8lqlHppOrvbOLaI4mhEYPsj7I
V14RuTQ9p2m3FMRKjjvD8aZaSncW9e6zQxAch2T1ugqniLW6jaRjAwVT/PxhzjF8
wN1kmGC056FJBPHzyak7POf6oIRBvfu66N6Bl+Qvh7hAKT4Os9YBLX4WXjDdKWcP
ge7IFNIRy8UEEkXqoqlRceVPhwBCYt4SA6cFxsmxExjBpt165sqp8LzIdYGSK/4K
JkdZYX06kIQn4ZhpSIwdK3vNdk97gIXBuBIE5JBiEU4Es9y/ZsuxpgkVwkufEJhr
wgbCs89vfSh4v3wZwSyBJCgN0EJfgbj+ga4jSXy+WLeaEO2rj6/OlP37lrcVbtK4
kPfOby2/s/raENKSRfnP0Kz3SskIXxRkuAXbamNhlxbAkNMd/s52jVsK/SP7Sjf4
aZlB1Ttmdslr076m7YD97qZgMBxSiTd8eR35t2dZNmdra++V6PxbD6SlbhAC2lms
Azg3ngovCbY8bc3IE7YzX8yoNnjaXQ/E4zcEIXlxKiQTlr1hEWyy78d3uoyB2Tyb
XDwsq4H7MzjaKrk3IWPqU6RxSfiCr9P5ewzUtWsCsHCoH8zj2DDt1Ahuz29QqLeI
F4KGb1ov5+/4vDj8ooNXcf/8PFBPPjl/TGQlVHGFG3gUmIohz7YTL0cyEfU+wlMu
duo8wo7hMmZQLf0AHGu1NHjoz8/p4IZYfu/NkQw5IFON8DTCBRfc+vbtpKZfi0eY
j/JuCgXCxohK459bfoF8MJoFmpYAXjrKed4tbJKFIGycENq4ULC0DXw6hYm4VGix
VQzEJx7QG6mKZiqgsihO/th9HBwzeQ2v9c0XGPOCEm/iHTQBVljRVNJA5UUXtVK+
Q/Se15V30/ayZxH23/wUkmALJjH0umvzqd9NrJLDYMxNiCyLPpByJepI/hkfQjKE
yhXBnn9PnirJymPg7hEenVJVGQiLOI0JsE62hJXFE9rtNwisgMGLmencWv2MyV8A
tZ3oB5zsv1htAUrfJ1CCCAVJQRX5sgvEmH/V6SSzkdXWBvnuOP3PqJxPF2f87nSA
dBxVPNI58uD8KfDVgfBs4JLOL0FhKdpfx7xIW2Y0VHd63KocTjuzU4HQqUBsMroZ
j0OZrx3RzgxBuXKqeOgD1BbOsL4C26rvlNGPy0wbUIaU83Pme13LvKEXk1GAJtM7
m52/0RRddfB51gZnch2K1ct5f5rIuFCn3TT2odDkH7tXRfcvLH7bT58YRiSJCcH/
1e5nJG3LKilO3GcjGXxI9Y0jDFhm3MJ5Fwozp3cUP+EF1usO+BlmbGLu3pGjYmtf
EsMqTC85YTVBoAxEIhhy8Q5tTHmEIPA93jmQiLHIKk7xT6c3fyG/BzMwShNDPKPJ
cTZsRsBEcn/mAXMtkddWzDnnuTI3DxlaO4cLBkErP/TMuk0y/4TAhcN+pumi41ew
fXFSVza3LqfkcnnbWboxCFWg2QYSif980Oa4vnJCejOhfewGiXVo4frqQl/bKjfZ
uH7c2ZbbfYZM3IYtSeqbJGlNCvRn2hfgL1lWPEsqJwLS9+T9LO7iRHO7/XrGP83t
LH7Btmsz0+mxTpq+lYh7FUYFe+/JslEmX1uofgW8anw0FlONRKzKU9OzmPdwK4mM
rJxuazHC7a+WjAF1N3haIb+zdFEdpB0HGwvdSvFjybhQyujVGU34I3OhyT0R7NwU
qHfGNH4JeO7QMdeGjgSjcEsQBGKVOSmartXS3cWkZlo8wK1w5ARG22E/hScBX99d
DbWuSBSJkH+5LfINFMbey59+qS3lr3EutBp7dhXK3kfw2LhuzQ3/6s+2RoDLqbUy
ZCJAIKcfVpLIHon0xEBncME1JfgDz/M8XRSVctkN5XiAlQoMgSKIW4rUASiiJbcX
m+NchIMXEP9ON5/51RoGCojzc390pU+FYNhZ+qk4D5tVq8CaGboqxXfDUZjfVus/
vh/B9YgrkO5XGWk3Li0Lso46DDS75MhyFs0kM5VQ73czvJnKKPnSTqZJPYqvnuFi
GZYpMUpqx29VkNrH89qy2tQyatv3TdrNR6u8uy+iXoxIBUsAJFOEpzTwdrUiwAgI
M/IzqE5/91GbEA+1hF3YKIWdddtG0s2HS7U6+4fX7+dyKh9bGsbat8gSxMcK9Tok
11ZfK+t/E5k5yGv84OyqlwSNhDI/4ijJWH8CBqtcjTc/1HOg2RgMCr0xxnOObAyt
GDtVwiCG4oH3xmmzJ9NRek+uD/U/3YOFLW6f2zccO8ZwL2uoLmcgkt6gIKpBpsTJ
C4wqJi9/ZOdf5CbTs6nfCpUM6sV2vRygQ61hNO4lho7/7K301kYLbzcdPivirFvT
SsfRiTQniHqFl/P9+o2tojnQjb54RCK3ALDRfdMKzQhExEAB38gsHK8adma3l3EN
TWTeoY0oNticceMQ7EVC9xJqaVJKB+oeN1/q7bPowZlkfwcyyfdThKbNmSrXsD+l
0pnJQ3dskhhptYTTUoJQAx0DEwprtpVpTGU+ZZHZZZwR1aZ5lJwreSqDsqRxkmF/
XIJurmu3lyvNA3eHA8yFojLgJt5KONIhysAj7+jhzrIjwBLIyyq3NyHXJ48jIRKV
6r+BwuxXrr8IVkz/8TXtnwbs8eq5wuhW7p7Feb6+OVRR9on7Yco0beCRhyzKkgj/
F5CUjmHVUUrSw0ChBYo3c31xVRMfSVN+cKtFiy2Dh6TKjPOgfWRF9peAEMxd562c
D5skwbko09+9J6USRGIMZ01lY46kHbkb108/75XGwGzmDdyUVXpwTtHQI/GMrV82
GeL+75M+8fNDJf1j5sr/yHYE8vJfy6/aGIUu9XY76q6pxCPahJX0m0jOHXjY4X3N
/r3JHyHhNBIln2pV9EZdA8rnPcCMe/5R0LINThJfm/XyYMRIEwAA3nNEEGQQ8Z2B
XKlcQQU0o1NvmPcSahKp31g7g/z+hkubJN42ASxOSzjtR1uwBioWk3z8iQDLl7Pi
vcQURSSBGjhkmxx2tfoCphP/oC3eayHZdQVF4dpB5CMhcc2NyVOUReQu5eqh1Lv2
eAAdJ1xQSmMwkEkcAKQgIoSi+EjSQSlrLhpQR5sbBLVlY+DdoAkWKp8ck855YISl
UJwK+uo9gizP7XEii32amggvcmXa9ZGcqcQnzFaJMWX0155Enr88nb5IXJbuPpaI
Fy7brEN5ykx/sOQeNPkBYDqnRpIOUtAs+NVxhuC2X5MZhxBRYCAoc87MaEiFzdHn
E3oTbkevFk1/Hn2mrWvYEiOlEpHSVLbYtmukSpPHrTaH/sqBA4hXK9WDxUdTCQwB
wfmfp0SxTGnARiQwIfihKv2y+MJnabdEKw2ZdvQmo6a3YVAfbnxX+zRVG+arzCM/
/nNklNQV93SzBmltkmcwxaEpbeMOajoffokMNpUSi5qn5SZKsHYIsGFu336wFMGz
+TfieDDMjw3AdCtTwkHI+CIq5rvJq9iyB4oqzuplJ7siwfH9lkueANiL2AEvrhbj
jVId/4sRO5GIYieKC7q5BQRU8AalG/qqsfIY5gUF0zRYwzMr1c29UCdPp/pOeGZG
KwothGTfSyZQpyK4EU3oppfpuawBpTrBP2suf5lmQjqtPyy18QMRJeEQljYOCw9/
D0AVXlel6RlgZF7dcBYIeS3hwPpw4n1S0RYDDl9I0os8aB7DmyRq1gd7tip02Wyl
NNIIXYlojuFXDGkoKoHI4w9IYYi3mOSvfh2NDXXUnrave9RMKEiCbnuDCRBlWfoD
GpM+qFZz5TsamZ/FB6XrnFjNmfHt9l5M30dD7YNMKIai8Ey0svcCuXgIq86E//mN
bNHBf3bn+uMwXPd1BFgkD1phnL6s57jK82xxg/ZedVBN5PLbmM9o4GF94dMRWqRQ
0bijVg9o22PFeHu78/VkHSqf4UHjlJx2uM6VukHWk/kTej36GhgH2PxMKl4oF4hY
PrUOPlqql9IrLAv/D2OWo8BrbojfBiRD40WqyXQaasYHpxvnt+vvXx5mSVTjFo+A
xENdrOMTaTlkpSryaqP7CHjv0UNe74UibuL56Uv0hOMzwTPf/A4JMeKVxc1Td52C
Xb+y2fCXJqBs17s7/dWOa77KJR04hI8CvoDTsmG0DxTCnTp319tKEooP/3P1kiMd
dBdhwwwTuZKjQKBLZYiktTFnOipJR5eNljef3iG3sozUOzKbK/GJtC7O3oJGEaqM
vwjXwgAuFrZJ4A3McdtSiENPeB6+DcaXDA62UyKEtQ4dnQKw1pK0+boBqIh8azP6
RRZZJgNL1ut+JL3kSA8aggoNgrF+qDnkC3R/lr69rY6ujHoTMp4xZ3IlAXJejf0V
mRImRFUPaLUPpUAzs5/smAZe4XrYyW12rZBXXtho/OwO8RvA8diz2s/31ERvMewT
DJph01xiVoBzLmhCzZWzHnRvK4Sh5mR4sYCwKZJwmNNirj7JPdVjwxUaIFnTenvX
/5pFPhXUeFQtnrfb82lkddQQ033FbVMRZQuBVRxIhaVRnbvqehlW7QXtMnPFmElp
K4eNug+L6URCzv2NRyga1L2721FOzbCKShJeGCrFTuR/Aw6SLG5E4uM7T5uNHCEp
QKEbv5OoRava7If6Jd+CZW7QkEhy91gSGWNtahGDuQMS/xOG5YkJX3SDukTjt3rg
Yr7JnyBnP2Tv4JkWPV13vxr6dYIuBqeu/UXSB3WajC6/e26jqf5Di86iV6S5CmjH
HMbpBb0yU8TMKiTlaIwgPjj2Oo46mM80VPCiFYibqQhJIMgDBxQJComPApKlWuZJ
Gri2gKU0YzezIJYdj6xbiKhvCJyzVQs4byEfCXmQYjGdqHtP2Ob0ak3NW+pnhuxk
krBFbzqzPshE9GZxT4XIJNX8y/aUfSFpSM0wtgslu2tslOgrOLB4fG2k0pd/DM/V
7BmjJTtYPU3rP4kcUDKowB2BgAUCes4dCP2TDiXVU5q6zo7ZtXZMo76tSfpp3Udk
G0fPQ6QEIqrtwkvYbVFRgC5y/XXXOGCDDtwtP2Aa3J/fZoRnJKSyCFF9ik2kTrbC
VA40MGeWyohWRCqXtF9xvscg/S4qH6fGzhLOFX4iii+CawxSWs7paPcgjI3uge56
uCdao+/GY0a3Ub1giNWF6neOOPCB86G7Ulwqy2qvNxpdJfh6xtZ9OgwmZOlYuhyA
mXqLDSh2iHdg8lrfkkP8T2rvf5T0b6LraPNENabj2LxTWUmsxlsgseYe+AauD/vj
h2p8JpEnsofaqKWJSk4c4kdbBNiL70vfz8gEvMAO80pFCkuKaA6IPr3jxugEmTl0
lEnKx2f3FG4QiUck+IoCwPupHzk250hXwWukvMZr74ivfNIf+7WShKVvHTWOTzWg
D3aBmHKMqSvr6fBhXtbGFHhNdxFis5o6aL4TqMKX+lRV0FgkpCz09nvD9NTVDVIA
2v67QbdV9lBAi7ZDIpVZKRmE+BMk2h+h9Y4LaFtZDRu39Y5DRZc459qW2/+8mZqv
I+Z4qL+UykxpIJowj6mmjwtKAmnk3nTqDEdXoR8NahiysCNxqd7+mIvnSvoh2wr7
yKlKTWo/Zuoi35DWC8HgNBdL6jmcBnsd9lyhxDBt+Ms4st+48F04fb6C0/ftIwJJ
JtubXu5wiVC3EEo77g/kZpJpAjX/sTuEBY9L/nhg53KO2JSGy4tnNtiSjHWYVqch
SwqIGY7rGco9q2Ep+YChiniHRXapwg/Cgb8i74SwhPnP0ZH4BVnULzk8SGnCmCLr
vm7Wy2MA8oUBmyYvcMT1Q4Lnk/tZ5VabJ3K/0nMSLCZwKQwSV5TqO8q1FaSHYzco
erJairQ87H+dY5qTUG1xn9rKh1bo5RWSoiRA+N7/4t7nrFj3+LI+jOSazGBCYkrA
RrANlCaEw3TPD6OIBvkOrOHfpa+EVbP1ehmxL+/4C+nwlrPslCBZqlLmZW8q+QDv
Q9ayWQ+mIrPQqbwPm97RIbXNPp8Hn9zBJ9WQhiIrDWyxbL6QKcoHFy+jvnhAzJDy
1svqa7rBGxeM7kUXSGTnwUEDlP4TD/Cn9FYaMVD7IsKvPB3vgUdZ9gUnpcSxSiOq
gRnsGnKKhCX9aSaTiKxP0aMV40URZs510ijBvEPTzp0XvE46FfNIRsE/EODL5x53
bsZbTOtBr6iIt2i6kTDCQTc7tP24tZPh8j0t5zdMCZxEBENCCM5AGUz35ucwttMg
qAk+1ywsgF09rxKp9Mr3KLDkgreUDKEOfOtz3sZXhyOvnAZiqgJo5YH3fjtBoXJU
TWlqbEP2MGZp0pl5fOTuXrMHzLZogz96xayU/V/0m4EbWS1w7LRGVMtszEbpdQ4I
9Alq12HBDJeEaV5mEgmb5JhbN1n0JChKTksmEILoLOh83C5PxLUL6pbC5hgUWsDQ
NMqAIvn+BOpv1xS7Oj9YMhniywWcaw9jtboWOhq/Y5phiig4ftfLdvXl9GZi+K41
KqsgbQSgF4+/MBJYg9rGtb90E8ydsuCatmTjsX547zK5T7SPmI32hUw9W/NORGqF
zF3pT7j+LvdZaLrowrWeMMGR++8GLxRUlp2KIb2KFjE6qIMDADEMdQ0cJcoc3tE0
FDi3ZCe9AbU4JZzpEfFHh6qBADCTI1EPRwOfc9azY3G1a8EdgMb5kVAEDLcXiqkn
mITPbB0Fggx9rE5TIForXxWo4DuWUk5T07K7kfk2vrdJpQeJe9yfdIOA7Ulje3Pq
9z2fhkYLU+cuqs4tU+vZ7FckR5Zv11NYYdCJO+5EqVxyGFoOqS1qRuc/fQ8RKgka
MJ8ui26YHc9p3m8iyGMj4EBILFdYFzHWoFjS7tN3yCUhpEECNFDb0q1iTY2ldz1F
E5u/TP2Ef8UZGZTOLYdS5dWMbQzYInV0SPx0d5mYhpeSGmEHAsMBdQ1n7j8mtnMj
rSAJ7p+0U8KdsIPbJ+0v4O1yYbv3rrt97Ps37n202zLNeTE4mjdkpLSOyl0d3E1q
kscEdDsL9yB9d7IH1JcC5IzJJBLNUejOO8G18faeZSXzg5rSjqPhhc+o/rKXHV1E
tKcpeTdnlwRxAKKiigjDoHcIveGzungxEaOae/B29rNSJQ92KNHAln3C5G5bsk2W
F7/SLrVxzEmEZ72UGEkvS6zswPS2nh2+OllfhOfvjwLjLFOSedofVLQYOWWU2xbt
kKCchvZ1Yl0PaQm9IiW2U2hyQtc2zaofzqP/xX+y6id7wqXL73nR9dcA0+twyipZ
QldIDSEMAn1U7oq+hoLsNR5HwURbUDh5naEU+Qx5ey7OwnZBbORij8PECaAt+0TN
47WUGj2N7Li1pb0E8HmiE3Jzp3tP7rX/zfVpBKMI9SIwzZV7AKVvbfvutn27Wp1J
IHFJeoq2tiMbZPH2vHFNMibOEG6lwH2eIYe6KNyuOqz805HoWikGOZA4Rw8tnIXp
pSU43PDuXmGBS+3yfTIvXv7czDj/zCxj+XjK+Mau8r+thcEW99lYQBSQhrPwnSfm
bcuH1x0qnijnqdRoCg0vN+MH3Georj9G7bqgN/vmNmPsn+VwJzc6D/BtW4rZUX0y
mTftroljPCzgyLxNEWpsfCRgAXBmTUyT7hMgy6EWs8K24mA/h6lwdZzCMwgR615w
w/U/9GK8hGd8zXFwkiyhAHbSZDfj/VYubgNLF4e/ZypLZTUeWtmf5DljJ2/+R3it
YnbYSgiL+QHrVYUOkphnvnoQCIlATqBmDqNAUoMoInyGjoiOp3KapFW09XihqXzO
iXDBETv/TCCRVAQ73RVh4vPYfhF5LvUCC/2yPhPN2geWhVHzAKcQSbRffO90hbmL
Rbc78vBQfZVt+tV1JUNxzakwaQxkx2/h0dH9LBqZ0Qqn5PLVOlQO4vU3rT/4aGFa
x1HnDfSkFS70c5cR+O+eZ7Q8W3H8LV7npK2/8DCrLbzBrdEWvCmNXbkZWcKR+U9q
I4OVybfNagsQb0JbatylhhxmQjB382MXlmcFna0+O/cerkZSm+04SOaXXd6UtyVd
HLKl45MfZ29Y8x5RgxujIaSf0t8mNcuqe23IKG+6gIcXDtpj0vLZ+WGwJbcISdhU
Ujhzk/N/VDhr/WFLGZe9iPVUGpD4w4dzIK9tXp8m9W5nDfVs4GT34l+U01sT0z4e
hXlpjfA8GVLtPAWlU+v2zX6Gg0uyuY60khSSrGeswQRqd9CzYqPbiv/Rp1HfGfCi
3QtFR3BZsm1ut0FOEosdH/Xv6r1VQnOs74+9vr2CpFS2jcJfrIt7E69EaXngCTEq
LGneOTkhLO6E1MMVEcs9fGaGuDzvca0hW823bLByngAgEOhByqIR38Kh8H5tpgMT
pnzdQWBwWRNjst0nNNj0cMJdDrqt2Zp0GAof8ZoiD5k5MPTATvhY5hCVJ5kO07bc
X0cb4obPvfWqFxZ/bR3QlWIM/f07mdNs+rvhPyIkwe6xE8xjm0KqYH+9VwfUyp14
JgjTkV+rN2co6lNFrRTvIrphtQFngJ2LSVheXBZvHu4ZER7rlmGcIsxbPuwAIunv
pzWhTvuIXORAUDV+ZLCEUo672WgZh71MSyOlTWqqW11Idt+LPf8+uVJtk65ftLGu
VyQSFaFIFhSdTe8m7PtITuBwavubGdKnxqXZSQtAqv7i2tLJ2x/LFEZoHRd/Gw9o
WqtWRRsHlRPdRz1m9JhCeuDZ3Fyvf9gKklTU8/pHYFROCGmxkCuiesxbgsPLmgn9
M1T+0V2lLVdstcw//WFzhdWj2jFv7tAcsj+U4oU2FydCDUQNOVvGfi52fk0+70D8
56d9Pv+GCQnURY7Bs8oZnksAt1G1MqUpDit6PjAyFwK3XvS6IwuRB6qkbq+AmO6n
wEae23Fa/Nq/IQO3CPgGefOQ+3M9pPcGO4UVy6tlCVhbn5ge6yu9qEs3gBcMWB9h
P3eycqXNEaEG7m8KP0edNf1yZgtD5//bZI5HEM6GFeF1uJx2mD4Wln4snulTIQQY
sPYfLPzPgUzHwIm5zVy4mvRFThe/LXcifyGR2nFyQKuzYLOwl6nvVwqUP3yDUaw9
e8bMuA/VqiGVA7V7eWZmIDJu/cZm+eSAKdDw9xc3yS5RqLlcvf6INmM92viLwT9h
u1H4IqqezeKun4oRP83o+LV4JasWvREb5C/UAJ7mfrsDhmnf9Ryrph5YeQqXvULJ
Ya5ZpIFqBRGeLD75eXp+NZHr5pPMo8h3dXn0W6hRwy89iUz5d6ApqhYdILpxAze9
LICoJKFjBNglShFORVkSt06qwmzCmwtPgQeKQrV8yAzp8zshD5ApMFb03WOWanan
WP8jHX7YfSBkiHFlZlrBWmUhO36mj4wm3wdE7LmkLiGaRNv2c6RPtABJ9Z3vVP/2
B8NvR1R/EdPrbgV/SBVj7U0darkvsKTbh1tIPBJCQQCiGd+FgsU0MKr77P3FGlKX
cuWz/l6in6nAKzwjPHTFCGck0FIHy8dT1U49g+WcndMEiB8KBWbWFBAkZQfWbTY0
XgWq2p3xhRe73SzYya98t5e2ahFm6ite1n4Qou+JdlDSwLlAdeeipc600JHR515A
N0qi2rfoNoP3nlfYLW/4/YMFlm0d5rPWPgIj/r17lBYE1VI2Hn7Dx6iZcIguRe7W
plwaAEoDJISPTbqduuOe+H1hHr5mw82s10GRbMANgS/GXk0xLFodv/S4SExDLLqs
WQ8EUrX1KPqxh21EL8WHBiDW7N9S09YnY/4iCNAunwhd/G6m6B6K1nzTINPAZY+F
Tv4R7EvhNWE4ShTkaZqz/N1LiLTMfNaWcbpwZ5glP7PuDl13BJi22jI6lCCQ+piZ
eErErXMngS7OJwkgrVEQWmvrQ0vzmNre0CS6iJ4dY6MtosR1YG/k+4C1jdHxXAUm
slgs61TLlJNMEr1+6WYALfCKJ7lFdpPyV3l/m6c1jvnJY2cCkoRJ7dJImOpY/R/4
ZZhp+al3QTWucynIXkRgnjEEs3OZLuxf68DyxYwXywFNXSd5D/96f4jrhiJdqBUG
t4UUi7KCuyhQuLOPn54Bk2iSrkJ2zdAJeQwOqps+mlNw9KDHc+4IpwiOiV4dfp+e
zMtMIdlVy/S5WO5hDqSL6Avpl+Z7pu4oPsWWh8Hrhvip/omZHGuOPnCu6tGPTx7T
LNjV0R2ztbhhaT7dVvwqLjVHmONamvb1IvOZKRTbGjR+k2Y5ixXI1ddz9aQ/BPs4
miRfUY3tbyf7V7d/xiUfDLdsyUJRDudoPdmZ7X2gP3zw0ECbfu7N1tLrCcpaZP9p
xFQ9QTet0BttxzLX1CUEKT44e2KlcLTrlHq6uzeglBDBGNGUH4yLNmSill0a9Ouz
7QhnuVzJtS0a/7s0TZplE3+C6TRlMxqGCc2qdiNSi4mLYUWruSFYlsODvJOt/uH/
LOBPbyQXdx9sT6tQljNWIQl4ckch0gosOwA7p/g/EhI84CM5C/JqAlTN/XXWaNIg
1iDsUC0opElMAIlR+5kcAs1eZLjibk42RfIgCneu7jB9FK0cKBy+IJQJjSBNeb+W
av6kxmrlARF1ytDDm+DtbgDL+Jr7YAUyK/7lkV34GjD9K+vCfkyxJ2deOHaIDFql
4K5d8SkpFZ/XYPn7FL4A3bO8EggNlWKlGLfioP4EYK1xactFHk3vbQIwSSPDw/HW
zMsyn7m/CkZuKRl6UCK3/ZTk8xKgwAI5jqspMudCK3gbuMiAFEYYMTMVOnLCTX+p
uK6pYKdo0pbqWW7Z2sbiABTYaTHggIFZg/IB6Kiz59uF+a2lrraJZVcNvi28RoDi
Ub6BGiLvlXPsejwBsd09Qmj8+V9N6b1c6Hoil/tISgXyMWlyZCnxAso+0/yEAIJb
0hAUixWy3XjYGnxP/ObL8XuTK3AiU0yNWaSIVxTl+ri/GW9Ctr2AYFCDlmngXAYE
ELwXCk4YkHlI+lG97Og48fGcNmoKzuqY8uc0neujSy+uxMfsU+ThyWW+lvhG0eae
s5kxB2woQ4LZNqSfdIml1JnLHXFQjagqDRD/z+ShdK4rUyb+GXj7riSMqa3NvjdT
FN05nE3VbyAqrwTkakFgv2WVa/j7nM3ENceaxGXmcZmntTda7QMvpAL/b0RGtfX8
ZsCwIc2jNjSxNFlBt0zNJfCyJqeBys9CoHQdWTHTYvBR4+DAj45JRP1Ks11Mi1/i
YfA0R8mRz7C4QDfsuyPsFuOxQrfzGOA5X3DB/ZJ8rodZemP8KaL3flWxhLynh8wH
U+RVEOtzE4J3Xi+h+ps7yO1ij2fvIWHbdw6gQXTeCyoHf+hmjBSZMRwWZblCCQrC
Zg3ifqqin1+po7iYEmyyS4eh6w1I8YpTDQ6bIg92Zel2qmbqAEOuD1RZh7AozGLa
ohyVgtjirlb1fWsmZQYxDhToK2YL3TlyftH34h+DZQROKq2fnoQF4O15CV2CF5zD
UmlRCr4dIPs+4wOHBrUg2yoCBKAbm2TOOxrF5VxQG9X4vjFkHTl2scX8BHOuRLs7
0Dveg+JHDNa9CDn8wjgdjZDTk941w6mpXgi8WRlnnhoVyo+bhsfP5sO24IqSWkGV
nDwO9qODViEOtzrnF2fJpZWZ3dSa2OO8aL5jlvr/7PK+k0DyuAKxcIulV/gS6sky
sINiNW4gpfX7yHF5gerY59w1Cu0cvvin3Un4nsbw7+ytompI03TkLak06kzBF0fF
ledcJu518U576VIGJ44HzRhXxDwVpe3KBZQc4WsjLKWiB31Yi3VD3WajL6LNCreQ
8J8Q4kgrBg+wR3LkTT8ODcwtEUrwxAlRFVyX/t9aBeSlW1YR3Hg5Od7rVbv0SRqU
7vmtEmWBmMl8YSzGSgnjK2/iZaRUiQMLokkowGCkAMqZnJcgFU8D3H7sZ4bHHeUK
vQf+y+hmzg8BrQpq3AFJ99elIlZNHEwFDQQiWpngPW/x49Z5yEm5G6siLGMZ9Y6n
oixh2/dH6D7y5VOim5YSB5MEFlSLdrE9uWjuWl3xCFYnI+lMyjTg1itjbgFQP/Zw
nylzA/70ioZ5suVlbADZ4JisJ02T3uj4CBHFYCbJtWd3jXsWEUC7JaQGLSNHuFn/
67N4gjds5tK04atP8u3IxqsH6DyYEdmQKr04Ds6+CLUdVthpQCHRhmAQPiHrJjU1
ukc1BnktbPRseU1pUwtohQeFVUIx3ArSp9MAAHkVSkaFjL6VoMVHGFha4PcgEMEc
vWSa/L9VW8gknB9wibWmCBZ/W8DwvCo9kOmk6L3M+VfzOqFapxFCgBnmZohojfX+
0gZBF6eLdTx9XyTyQLfaYhJqPHpMUqC0GF+l+eBd4McaFAY7joK6i+5maV2GuBld
tXSJcEAXgro0OdngUpzYfcOOp7hF8M/6bp88hho61mMojC0NyKne2Xg9rBJFHnF4
1bgOx32aKnbXJHNUrRaviF7XAYNpEEEerVhYI9yEodyi9OL/RDbLDn7HmLJjXd0l
EcqR6Q7njR0KHVJLlPv1MaE4Hyk5d0Nvrc8pnWVUUreiTWSFLIgysl98jj7T9IBT
xWpAzN/SWBjR8aGbfy+VrVPa7jtGH2Wh4XwDhDtcEhwTwjuWq8v1ymZawUs0eVYw
hkYrf1W1ebPpEGY8fj1s01fg4UeJBadnIFRnURway9Eryb/5AOuXkL31PapHroXk
QFqOyYiVIw/oeTBoAvdJJYfwfBZ+k5jmafs0T8Xmm1SLa4kwADUb/6OVHcLwxXCh
yhLhFILOtXBuEmiRQrx/x7nNQ0vAqqJIt/oHFhUW98amim/uyOpnQrVNfviUzEW1
zyc+G36fvPbNyfRIN1fl/7Ar9+kl06wzowkAgnKcmkY9fBYiFCzL9sKYTait3tOp
RYYsJV1Xfy62VJ370rgrE6TxsW5H7omtb6Wb995IghYCSkyLrD99KHpRI4sdWGHs
Y4eZNF+M3aRCZ15PlliSgnmRfXHGV8YY5qiG+fNVx6KHKish36Xh9TK396I12GqC
k4Yceq832TeqY0pjTQ4fKtDHM1KtnIIpUuMvha+HJUlEknyjX81IiPnERMDngUSf
MYcZSAfBmpkxVfCRCZYp6zAZGE69TLyQ9uAweb8vj3EknKy6DwsLVoBHLU+K2jrN
PNsW/1kGnxbjNSMVvUyGCjMgG//4UQgc+DkwPkuV2BREsJo1ANQ9spLNn+SnMcJO
aQ5bfDCVVFAsi4O9UFjhhmpC6LBE/Ye99QwU1mK3EF5Kon5mMWBvKLnW8OguVxRj
sw/gYxTVRl52Gx48cM+DPfWE3nI9IhPx/YtHsmP62PntEsUX0s/+TJOaSny5D9ZO
kEB+YF1lS5eJnM9sf00KkOX+TUCkzkI+9/mGMR+q96FxxwzY0OZ/55uWpcifOCpF
zKMObPnDNYlZ4qGgojJVNXQdr7JutAda3+8AutuO7G3PYJBFMcpeXor6k3pS2+lG
20yYZsJXAm0uXYqU7xEM8oyZzOIjIgGKSmB3ZbcabHhrUj7s+icLjwDP5XYm5ikP
vKoSH15cx0Gh/7cOyM2IPEHqtlkGGAp5uqW+HPLlD8KBHZJZO0q+W5CN2QL5W6KJ
QKTHo8f+VerReYpFmB2/Du91QchF7HHRvz1s5og3e+pMK2alWwC3+qMOV/VogS2R
+FLT/hvORsuR6lN8Kinpc023DYSNTl+sFWLOUpr/c6uHUujpghJqf6/5hlkSKnZx
Mz0moPn768aUccPHKSeHBq0Qksmd6FlwS2GSH4eE1cSoEkNAHL9emUMASuikfsy/
Ef4O46akMXRq3hlXSK3OBpFGyWnTEzrHkGqEpnPN78eQ1b8kJSyESR+bnAugSQ5/
mo9VPHCjg0Xy5HKipgAwSuXeLU+XuLSfXjPR1wPxgaEG4QGpKcUjSDcRWOOyM7D7
+RCV/k66vxPqqT/tlsuOHm+y0niDLMTrf+tNaL3eBt+ZVWNbU+y4tVkY/dHG8Hh0
ZQGHaNbz40BLrsX4ocIgtMzLWhbNseI2e9gTs4QavO5X6Q/TUW91vJuFgyfkszCi
duncEGKNNuPsDWPSNdLmc4msGK7Pt3669ktu0DEIt/VrkyFgSriHl7uA8+uk3JC3
EFX5+EHpVJfjHVz/v5XGt6MP9usqr539X6Ryg/VFmh0Q06WU+/ZTaYN1hO0M0WsD
W5IdSr4Qw29pW5468mYpCri7Rg4LHGejKWnzII8EQwc0ehzJpY87PJNjgF8ecVEX
SRF9utjcZo/Mn+GPvqWuvUxw6F4lS6SRLhnNqpfCVCT7h1aM0upy1+3GiE6VHlXl
pI9eSzBCRL9H3ofMXEqLcHoNGTZd7za3pM8TL4M4Q6UgpwAQIEjPOJ3T4vQj8sXh
1k/AP+n2qOAwpJ6iJVKbjHKZsnPFl4QwhNlZf6sDMvsEUmAsVL0/aEhpENVX3mIT
Mu2OdUUU/0pEmHViPi48vA7jxI1Wr+oRpda/QRPFEW1maszGjdNNf+GYrZTFFdOM
Nm7PMg/dNF5cniQzTCrJ+l+u/4+mJb1CA3MpKZEwzMNuyDrxxa7ejeG+c9a8UPpT
4wwfK8DU54zOFuIbwWZcIdRiM9Byq4d3Y0MZsiU3VJCwTwY9A+VQEIufi/G4S98V
qnpIQ7ncZ5EfyxHj7xpLx5JveBjJ+ZlT6DYuf8P4X5p9jDOdRIM8kvQctw7l71IQ
DkfpYpKgqw5ihhLF4MPW/kJE1coS8JvlydNZBsBi3IKSNX4dAsmMjwfMbfEVn9qT
9uEP42ngqImSjPMTAgLBnqVSxwspzj58qIk06ri7ZpQ4lBl0MNVDHk1Lyd9ra1Tv
UzypmomXyFlApORJjz7UsIiUkuazou93mPkAk86N+7+tvv4qu+W9f+asQpfJhDdb
bQyvG/zsILGMYta5pEDRv1jHQ+P8Yp3nj6LIOoZy/Ww3ZP8kNeNYU1ykD5nxGEhn
Z8bW4jOU0OlmXFMnLHcF8cPrgOtQPeW2XjO+/sFlPBsL9H1Q2YWwiYIlrnzegD0w
OuJQav1ZxZz2dsjut4Lj6idQtaR1rAuHxUbdk9mefiTCoT9LRZwgPbqrBDc7sV3m
QzA6toWz938/4HI3wVwY8EF767gpG38sBBqXG8D0Z6JLvxuU7+FMPp+Edu/iBnqX
45vQn9eIqdkwbB6OdO9HLbwH26KElUOzity/hUzuxP4LonX6/9jwDMKjTlTpgFCC
tqVzmeIIlvEwfo2rqnKTSqhDoFBQZxZSFKg4MD6SFhDhi9WRLit6m4tKYpEs1s0m
l5lRiWIUoXq10fpWrLB9qMyyCsM4uKOpSJfXQtLWKlPRXd8791KaGD0kk/X2vPXy
Rh6xygJFMMRcnGTKtzbtNGFhet06vCYNokitp+W1msprV52TOwz+PLO2Ld4WEdsb
GmTctJJsEVbE9wvgKG3X2gCdiut2/OCCJgTs8LfSc6Y+tJkI/DKgLOntkPu+Zq7D
mMku/xu8lbIU/6d3qoIsFBW6gdj/yFLIibkSACN+isu1nbo+fHnbytaDcM9WitSX
fnAuH7uDVXY/6HHAtsI0lvdXHH/b1Lfe22vsQBsm7i9L1TfWrX2JVggMvQJ0KAak
6pAFCZ/mmDokN63e8aa2aGJEU4qYQW92/Bif3tX8TZKrJEZ+XZz24XOovpGpAM9s
c4CBqDyoV+5tKCvjxF/XfPQOUYkw+jaqsHJkGw01gu0+K0wjk3GGyDN0Kz9Ja1Nc
KnfoqfM+d9oB13UPq4OhBq9+Ykiyd8Z66uZP6qSFBsMBUxxuzS6hKf51+AVyQUJk
ScGTY0wmCQoQQ140O52THoTpGwrazcZLNJ0hjS/Vfw36TuvlmjjsGJoUdJcx4kY4
bOsHDcA3Kp1U7T1/4MEeGirCbrtDsWFIxHxG9ioBmKrg0IRwXa3JrWmuiOd+q4T8
UH3Eq6GneSPDVs5mOpf4ILoX1dh88ABEoXrqOwwpIuClF1l4ZcNfDw9iUuf1WwGW
ALdqnTDeUEXorVjl5X0fZ9PyU5svRMNs1uOHqv+sWEgbLqnj0rAoaJoQ4kWZDfpL
oV5vueGq/TRK3Kb8My9h7bqyLBEm9bIeSjQOt3BBNrkGv42v/sU/nyv6wIF+Higp
rU1V6k2Dcejg0ULghAHKEI6c/eMYpZPQLFjXvVwzXKZIJt7huiSy8FUtBB0OYJwu
z7hnsNZaV5IeBOISEonTY7AgJZvsQczMuuEqYglkGo572RBJvan0mvULI5JTirCm
B4hDUUWwB49mAS5JFN1SSpe5yyy9mkqf6anfY16ANmvPKU59iBL7QLmv4GxeOZFo
jWfyAyQg2Cdmd4GNXFTf129z/xn6jLFwwMgSh+v+zjEh7dn5hnbiLGeOXv3dLPFG
QpCNjYePcNjKd00RQC5dC3qRHcZozAc/3zYXgR4xLkX34m3VsFv+tOiZ7300FiRZ
6wDGBXuRzgP86UUQlOGLvZ5dw/EdYGGNx1B4L4syF4SiKb6S14odTzKDaJjQGbiQ
Qe9M8QyonJb00oz+ICDoBkgQskB+AciNXlNyhQWs58YGEILrRWdknCZAzGjEWOGU
cLcT6Fzwf+bV9WoGBEe6a299Xa1IqttDmXfnIWk9gxGoFlpoRm59Vpr9VscBe5zW
yl8VYjiDE3+8M8dVAvesXjeia/uzsfsTBTV/Ks3a8VNZygRk+qjbcHHLd2mt9Dy8
zHxzBobF3nmEorfiqOr3REPBnxYU1GeMApa2ssiEOlUFCVRbemCrrZB4BNzB9eAr
mLipWczqkCaHyq/kAW7jNPXgVeq/TnBjdsjs75B3CNpC1v7S2PGa5wYlwQhBGYDI
TQysJVx3Mmb7gQk/R8p6Uiv50hY6HSwL0wdRIk/MY3/F63w4V5xMvUJj/HF++a3X
GzBGCzmP1qjd4friXhyqpL7oCQo9oAsnXHKawM5S9EQe5nYPnA0u0KisT1/38/Ib
kk5+KaorEPPyN+raAH3ugDhrp7QGI81QX4CSMI08A3DbqfUHIo5vAziYRuIiy40i
BLFJ8ZPEKGsHzkAX/yIl/+pvQz9bldpxvpA9EVHeau1OmBA1wYmNi8Hzs7VEDfaB
vXWoxJaN39/VN1jtOldRc3BWtNL0Ig1it8/2vxWAR9RZh5Pv8udw0h79CbB6olLl
+UPB6CaDm6LKrWsx4JBsnR3mRLSjiWgo4t4DLfna924DCunJl2hd4iqfpE4RnSFO
WF+nKyNkrJ3DgS7pjxmEUAPUKYhw+dEDkgmfOLyM3gYH73mZTZ1Ws4Io1bOz3COF
UvSGKlIUgUEwhkHf5bfbJEwMe1Ipaf4LJr5XTy7/4bQO0QtYcsCOHB92UMDdYC/i
W3Auxj4MomxRLg95mS0sjX1DeOACupyVC3fHrmg5QkMuTLRz/Iay/RZYk6s+4J79
UhoiJ2ftCMN2T1WyoR9W2qQNHX+Z/JSXyGTNY3DVqJErciY+yEh+o4MWXOaO5Pb2
Mxx+06X+d6cwkS/yW3EwfN9MhuY7MxOfl1jwHR0/QJbCexxYjoo4fplVGIZUSffh
hWQTEB0sTD4bUeSzGv+A13612RZZ2TykpwQxWw7oXKGyPddrFYoQ0rIHK6w4Ftnb
7i/LRgw9j2dUA5mByjyy4UPIx5YqL6Nsdi3XgC19KWZfz0QVVyHPllNhkVis8rfP
cYzOqLAADTWgwcSfyXfH3a0gGu6QgQ/GX22dXjqaZ72kSD7BF1uuiysFY9ifsT80
4Ah4ehaTlrk/S6OO/e+rR6yODU3SSjbw5x11ID+LSdeF33Iyegm923V9rAVWvVkg
6XbxiMJk/H9cCyUewMnPmDm6JUG/Z2m5HMYo9W/AHCt4V1ScPWu1cHrdVbLuURKA
BW3Dz9l5/sUfbzOVS7SlmZ4acx0TzYiM83pbGW0o4Tjg86KXNb/KjR3d07YIeqbr
sslKSk4tZblcHyE68umsaYJ9ki0pG7qe09aonWLuq4UUtLSHLB60UkbmN8CQneHM
r1qhzMYr2gtUnsKAxG13LjU48m1Kri1q7AAZ4HgIw39FsRxITk25SIMdtlmHdoQ+
e2hoTcwZsYCI5BUzT/rzXvjvBUdeh0fqnkIXq8wEBf03UKejpKdvBWWCeixsHnLO
aginaxFOkqH0h9M2jUbwnffzGvbZmMyLDo5ajm5KX+n/Avf/5M+w70/e8wBVPysn
YbAl9T8zEFHywu9bn07Io2+GUX24BjYWfSWvooBwX+m4jUYxUOekLaSpoC8RrkG1
XIZAcutc1Vj8y9nO9+diMSpnZnCcGxbc7BDjHMLX+RCAhRFVKqIF6vagz/InR/gr
HS7te5U6QDypPy/szl5dYlqWcWGObFGR7mXbaw/dSi0qASrvi5xWJ6O46iZNLABE
oi6FQ+zOdjbeGjhaX3Km8kPwBa+UlStNNp2Z4saBkPxCxtW1iQqaGtDxdvzPiBdj
D9tsny/DSjr7hptBGTYDCj3XdQNllC63xLpH2RQkZ211ZfNYv3u5J5vVKMlSm3si
Fxu/9wwK4g4G/7ouYIuDGTOjBruUo5+AuAEXbNtZ44tA52zwJLVOQsA+ghuFKPaC
U3oUtX2CByzwS5TNdxOczhRDqfk56/5Q2Hn7yB1+yxJjshHxcTfkaTJrT6aoRzEN
E17kAb8lEX6ChHyAR3Ix+zJW6QmkE8wTcJzc8H9J54bwsVa7CphUj5ocsRqRuc0R
v2YGLPGp8BI17IQlLP7s/YxgKYYqDbeK48rq5oO2iKq61Sd/t7RNs1bayZbv5v+B
z30bpEr3sSmsXtTwOh6GRr38r8rPPCBoLP3d4kVy6Lb/Sf9yQCNU7BfA3upJzl6J
n3uTLeNI1RV55iJAvuavL8VeXf2QxcFRdpMZ9hwM8cfNYR3zdH8eVat5ZG8aCgVf
ZIRkC04pyFafFj2nzvXN+z+7h3+tSJ2o+V36WEyWXELx8/DS3vYHD1f1UvBhZtsn
9I4xp3iELJt590ySpdUOIXH23/76MuMQv41gNChuIzNGaYV9uNUvSntVhrUeYOHr
BTLRvWyxAAkFN2m6OlkiX0+l/USomLWBnTYJkEI5kfpRo5rdVoZzraQcCeZ5V8kO
/xm+bfunn2KaFE0iTBsspQKZrMbXdAskp5JFjr0lJt5LKfNFNfVisWEl9ljcBP6I
snFOI5wGUTVP3fQCAkfjIg76xuhBN4g1bUv1xihR78qeANdwWx0H495HQP+bPwS2
nYnNn0pKxUBAaUiSykXr+SX+ZKj2NP+Dz/pS1b1xZp4HaV+MQBeTWVkhvS4CnvOr
Jf5iolz5jbagaGTGh6i7vjiOAGds7tNDxgteLqc0I2lgYAR6L95MhUNMPJoenaZ5
aOY2KnU9viN1rrjzLZira6TijMF+mTcWc/SSKUAs3R470x2ng3Wh3SJ242QVw4To
bNnWvUzZ/Dtp0TpZlDx/UDu5iaxOKPaA0fge5kWXFiXiwRXQhTaEC/HuHLIeVyuz
2LI9Jd7GwU0doG88w8+FhyV6frLeo9Wxl+d/BIR40sTSb5O81ohyDBlHRl4+1S2n
4subgSY6QhLt7erFRFx/SwT1TbZCa8TQg675uzRdw84k2cVjfkWBzRo6Yq8Q7g5j
vMnvljLfFW3Ta/9uu1hADTqHucMxxImvNiJ1qYxecR7rGAjrEU2KEGyfBCkuG9vl
xhZMF3smdN9Qo2l++JCnwppyFy8Mn+U2KauBpdw6tzeANjOMyk9+olHktMa+/Xhn
oCGsFgVGc0KC3r/NqkyfP2f2/5BDb15CgSA1714r6v51hJ+vQ7QNIjTGnmIzT89C
mjhedDbPG4Q39WFHZQJorFdU/JOVQxTm2Y4Mno1//Dl9SAtTpbEUGr+4541/a0Je
3opweUSUvITEbQDzXhlWzjiexMZgN3fdL/jnEZs3/DC3MqRHK34khQ777lVU+wyh
KltPXMmla0eUU39GfSZwmx4KV/p/xiyabvIo+MInwYZawDap8rwodL1XsHSU6L32
PaF45ESLFnR39slSZVRVOGffowhW0ljDnWWfq4cEc6/JwaDF4uysWQ0Ynl5wmeS6
TilQaJmYKAv+MbSIm0t50K/HSlSJxpm5CQw9oIMTjzaZgpoZBYG4NGXKhClYr+BJ
E0iO1h0lmJMMOh2YqL7Cc7fuYY+aX/Byy1V00JriljLB+x8rTVslyWSPCP2roWPU
fqWBP/g0JHLuxW5Ju41eSds7ah1MDd6GXCpfaRivYRY95m0Sq7TLMvDSgpMI/ug7
OnBXXxHaWnymu75BCbB4HB+bs+pRjDi+YJG7Pje6HZjT6lRW0/O0/759ue4fYD+7
FIaIuTqwGquiT1SAl7FfxFRdjGtHzZMQVGENRt7mQUyBRhFSx40ajF0IJY2SV9o3
qMN+vYp2Xx81QjJNc6d5/g8iuYHPtpAgaQO39APLpaX0yh7xh7FyFvpgRJqQAfds
B1RW+txm4/D45E/WszvwoVj3lOKHbKT+toEKB1EAAdgFMcXtlti7DupcTl+TkIQo
+Yd5ZrEFoJW7E4BbaMcps7RAue9EjLD1+I0Q8g5Q8GUTDuxXOeVWUS7RAFuR8E7x
m+kRM07ZH2ZXZIrMf4RTRz9GEckv1o8vHD2dX9PPDJ3R80zs7LQLcAtht5LFsXt9
n3YbE8gOXXw4QLVBchqDsXcksQF2f0kqvKMOm1dQJY0delkzWJrkVuY+2qMBhEvv
ZduuQyNZ34OmxIBhHHfQxBr2h878KJjUA0H4lSORfpU3MUWLhNrRUQ1adtk2lF2g
OxPv+2HEzVsP2+EAP9486Yp7RXxgTT6CAl43Y8pn/6GX3AKMka62NCcL4IRIy25q
UF/USdbbAvq3pKekQOoMnC+Kvo4XWVZi2T/f/s/Tn08e5o+IfSbbcKxqfcM+ee3Q
LlvYnC6IgkelOEOvPJ3lHB7fS+AQbpllMptTMSUw6gSAjtNOgZxyl23pzgRUA2ut
Jexgwn2Vj6FVvTe4IguMppFN2vbiuVM2qn5wMEBmmyA+oZVENKKoBjsM47/HnZnR
z5uMU07aH3fe4AV1pW6uf+s80rYwhWfYzcJnMoiQxTdiiJj1NIVEhZUs0jdzsWHS
yVbgoieaQblgUUaNebNEGdUhJWGh8sAk9iY2Udofbq70O6JybIBXk5bx9AI46UHx
ndj+81PYDdP8oWO3RLzib6GGtW8xzboMkLZ07zRK6qj3VkglwaGs0B4c7C7598jt
augn5X6sX6StvAD+bx636hxvRwfn5x4lDMy7+R77qz8HKlTTirOBJKLY4sPoaeyC
suze3SLM8sEzWD582w2P2qE1PIx92QqsKKrq2EDm9dkwZMhzs3jGRPZL2GiAmvCU
S3KoJzs0ewqyzeXbw/K+5No5w0/kv68JyYyVE5NjqYoOyAhwcOXhotF7asLu0E6T
AXTx+8IDwCvkLC/X3wBY3CUg2Qt1x46++awpUn49BFQPQ9CGfCNGqNnWZFxrodZ2
qf87Q4qhqE5lghSD9xsu4PISB/fuvQtxjzNQ6PeHUAzQz8rBnExYN7Sg/UDKtDLb
ELyq40c72shY9xiUokyG5ftu/9wKRZmjBr+Ur/3utcw0ZgmCDmXJDVd24JUctDlX
iGRpI1zOCjWS5GOSgz14GNv7J6zgAuXbt3SLsQs0K2z3PGuy+V+gEI0yE4tyULpN
aj/bOTJZGJbTMCTQny4jq+xeWVjWprvjumz+QPWxVf6fO3Hq16rEOgKKlXHQaAI7
w8IVc0t8IwCUEm2G1pnHFj7jQ1tlAIm95YUlRh8NtW6EIiR4ubUIVQkE7KigBC8T
wJYnmm8GxcVJ50AckWUtCn6tTQOaQaLzEgUEBFA0UZXvAumZQ3udiB0GHDfpHDpb
UEm6NfA0Yz4+Nn1Mfi/U9SsotpZVTw0T0qR6bSmIGRz4RknVrtOCg2GE6xOTHwjC
BkhLX0SeOEbqDkwKJQTe15VSTQe7gXZxa579UHGwKlpNN/fHAfbcywYvf3P68xdg
Mw+j5u4BcRx7AltPPH+DH5lBS5Xs4LtvYevpk21KtoXSevK1KJAPchjdodBnKgVt
skWrbKFz8kuHxKQIyRoNdW5d4AdW86YyuW1PdLd0o5ZY3grMnBh5GfkDZD+CdIbo
jkIneWUBBd03RW0K9JnpcQqq5VMaqFEV78ILxdV4OVn5Cf3dwF4vBCvwpMY9cHM9
cJDTlvUS7pZTNqKtsh111F0Fv6EVHpvhfBcf4kV3BIfv1XU9whPhWmafmExYxbex
n5CmQWHagNqaQ2U4uK21hdDYPcqnI/Ly3yBZlYwybBQWeCBFAS2Ypdf8WqESNy2Y
EPj4YnrRPwGJqiAyErd64Y+n+Sok7gC6hiX4UoDL8TUbgn1Jp8AX51eR2Lv7pfVi
/MyISS7qxjGdCCmLx9hBvA/pBuOv1aST+mVvgZPA7d4HbK10x0qmQf0O0dh+uL4y
kpKQ/cwJx8qDxoTuE4GubM8hwA/rWR6D1bBnIgz47rIGNEfr5RaBdjlh1kF7JclO
JqFv2fFDGx6zp5fN2vudixqsXBRRJZ0CYyH15kbvzxsCUVIinWzOAPeNTJ1fgn++
GtzSkRMBqGRHhLVcZJj1w4Qq3h8Ec3qVksRmVw2qG33gpeOGifgblnlhdA4knDox
81l6G2k2xZ2gaV3v1J6nMOSJQMuyVS4QfNyZHZYmhhI0Jmr1JzzNXwu85katI8Uo
9E6y/35lsImRnWINCqNg0usJWRV+EYMslkYpJZ2kAu6NPZMEgHgNpYuMdYOcRT8r
L/m8CR6UYF7CV0EsGbpJTenWXLwgaRGs43xyjuCe1AIr0ERmMcUNwEfm+jzUkJFj
0aRwqC0Npe2/gGi9prRleH9O3iKBY+X/r67aMxqunuD0V9OmkkA+HPsvq87BYI8A
UY/sXomrs1E29JnnfN8VydLmwcS6h0tDyr3FMC+vfO3DhCC8VBG/KCu+ARsZCWJQ
ufKqtjHiaIBFFksqY+nHdOERThAYqebO+pFYr67ylK6/GNETA5jySxy7HIyM1iSV
9f2rJeKkHhG8RNIEbM5UEPI46p4VpoekaDG6lbz/7w+WDwyLq+jp0qEYdPJ2ZV+e
Z1MHzMPPHriZnArytVGvq82ed7p0P1q66ZDX+a1zNAVBgyoNv+u4s8rITEJ7xS1g
+scKM+KnxjtAQPS5RrUMoLnDm8SuPNsTiN9U0d8i3yY6XZYfFO5PeEy9Syr8MOXo
1yD2qcYXspP9pwKpGobDHd7SRG3TsDpBBC1CqKLlSa7kjHl8QLkcfKe0hq42x051
6n1bCL43GBo5ACuA0vmVlfH1kRkK/XPBL2hQopObdk/4O7Yrc1Z39yRFO37m7KEb
9mPpC4uiVi/WQPUMLEyWHehxBVZgEr+Oc1DpfMf1ZBwflVWevN9Yzoah0bIOj9B/
mrq4yXuB+Q1FLSYL9Hr0cvKoWaXtyUG5+tqgNMleSMw9pKCG1IYevyma1a5ShrSa
K+VYfAmixD4axVdAQs3NMOzbBBvRTWwZDvLwbl+Bm0sy/unf7/v+VgHvCmxnljRT
ovV9O+5J9YDYeUFAv1/t+2vUc/H02+oOgo15fIcDUPjyDB9g3N/FTkhYR3o5LsyX
QUGh9bcBw4hLk+Aes1Rl5EtI5o0lNuYJlvuSlAm7AkWRUcXFfF1VKTjfWN9Vvl+6
hf8Vrr5zDhKjU4qS9DG25ZNGbR6qxXsrvJ79EJ/UPMf/eFR5Oq6hmFhpVLn44/qa
bLBY/vFEA9UU8uLuY6F7KHcU9TWjMbb6ShgHxdRxQQNwsB9Kz+N/W7PlS7QUJuFk
jY9gA0NWMDzGRjTj83TXyZMqevJDH2yo3+ixqfP+Rtw939XlSjs7QjnbqI4jsgyQ
etJsU/dFlszYaL0A6ggEOJGsnwcUVQFSommHfET484R6dev03taxpCNN0egpBbZL
kI+nnWAUcbRhUg9+AtOeyjvOFUuXchJSJGtdPRyqAFtL4fM+FPjTYLxqZv7ChepK
E7uJVsbBSRD7v0xx9uM8botCM2TQO6veo87hSAI6h8W5aixoaLGaskJrqLolJDMM
H4KZI1xKua0h5wpjNceoRFaQnHslkX2oGn5kSJI15PyMWEwEGA8/GjQlcZ9sW0x+
/bFJ5O00my1Xsk8g13ApIclCGGWl6CW4io/drPCOjCPhhN7CWwbUgHx+JWD6ubqx
Tb5TMiLrixxpl946OfP6Vpj9QHJ2kOi63rhZWRixAnQZ+a9JntdOur/81n5TLVoK
wYxI1JAUR20+K3F3LAXWBbmFzAC9tjxVSUHv7oW9/hlD/KECmUtaGLH2LRdR43lQ
kNUL7SwWcws6LTQlcn5b5dGXELWANnt7XUSCNqo77Zoozuh5GXoCHNp1c+sJhQ5s
8h7yZ9jbV/Htq+SWctBg9/fwUIII/xar4/JojurDnkZK6kwRM9gnaJ9c/xlQtJG8
lF/P0ZWk+o9Pz2Cqt+v/J2CoOukEe3ppSKkW7Npi+YrOpHTjBYiLh69Fa6y909qp
etzjjSh3CoMLs75ESUiACoaWUL2iblBqVbDRT5VAqGncQdYpw/JmhjHXflhAOmop
zcSEBif/6BIaXPY/kNVmmYffCJw6LKeN+p87cLgwXNjqCjxM9KlTJGkXbzb5n9hK
dJKd1gLJp1TgtPBYAMw9MkyvxP6xwJEs3nzhTEIzxGYz0EjXMb2zrhpyseBy/BtZ
FiIjqlDWLh9EMMEASspY4Wua0mTT3sJI+v0tob3qC9Nq+RewgIK95nR1fToungYD
Cf1AkchjPeyWmwvNVmscdhVrS8qG0lKH7ALSQmqes8ZUblckfJK7zS+CF43BikZd
5n+WrtU1f0OVe5gUW/6v+NuYl87nrdPrUMUB+1/3sxh2KRtz4g2PbCUOx7SsJ/UY
40kHhK8EWnQx18M+NjTjyfKaaTnuuUZD9m6ozgL9JfxY9uHPoT+WVOPioetQ9Wjc
Nyzp54b26z2deJV+0ey4VWck7H1bx4k6EhQ4cFSIXGQ0Lac4Rc7HeubMRCxD0/A6
NBs7x6NyE9ks7DwTVRHW+2QXlwdMOBTAxImNuNYSfJnrsNkC46iZizSv7e9T43Uz
xIvJM8qRgGw86+UGQU9Og/dB6K+ewEyFsSVXy4zsPzLVYHaqp4OK66XEZHVDzWaM
cgKzz5WB3woJZF5dJm8jEPWbgKAILy2HXeCI/QWzsHK7Cy4F0LFSfB3mgHuMzu7q
iioyU/NVZGxvL336AjqevMWT7ftgYWPypFvTqo50LETmFc+aSEwrW+QiD2QgVrYj
6l7rmKLz0HMuGI6ROIM3KcslbSyr0j/FIsWZFURjYqa1b+paSts8xaiqiv7nOkyD
q9kH07mh4Tp/hylquTxV4N0/RY9ZofxuQu1O2bz1RIXI1k4MiiFuvxHzhIN1qurN
Rvps/y64C3GUFhAyPxhBb5/nKRFo2s6S5ue39ttE2feU9tEKH9Sl63sDL+Smlx2a
MjSrj6d4zbh9rfGbNj1uCYoBPI3PF1jeTAzOlKJ8s3wMMjFOCW8zTXASIykq3/kO
wqYfg79RV7M2tjpkoady7sOYbTbHHcWx2jGIxTCVFt2IL3xzpCQZ9Utt/2bvFzzE
6GldXQWRTIfPYUfvycds3vdSuzzi/uwGMmhMgf3jiQdCO1o6ug/dvck3zEKLbclx
tyxD1Ywzbni0Ff1uXHTt48nCOeYBlXu0oyeYA5NBGnwCYt6ttmQc4XlixAUecjAU
BRf4Y+4yqy/WZ7lslSKTCYOXfi+R6xRK/kACjhvzwxcbjVOYEXxtndYmyUK6bSYm
gFABdSwcJ6vzHYSFjsFh3+tIu+6J+klO1Hf5xXXeba8tFyx22FKNR9glfoe4PtLU
6XyVtw0Aw/b+noODusEsZkbxoA1dBQiHrjXtXc2QXJy5Dv/ARdJfT+FzMvPQJzpl
LNlasl0zxC5Zl3ZcnfaBpPd7jG6ACQ8EAEyuYfX0aD8dMRec1BANuD+GjC+569dR
mpfOVXAqmf8l0d6wrzbkhEur4fukXu0muEWUiEEUwTxv56YJ38W7f/fc9JaFx2sa
UyYdHcKlLiQjJMEYbPKby75adLd6QrXec6Z2/roYTDjhZLUCXSByxwiEk6OwN8eC
eKXgje0TCPDinyRJ86Fv7Hj2849r2YgBI/frHTQnI3obmleKWOX9yDyrDSoq4IFC
t7M0b7QQq5lWNn7uW3lG44rATaBgFOLEs1iTGtw5ZQf0VnNImqd++5ATirJE/rgx
QVDjpVYN8TOxm9R73RKZSSY8znLmeCf5qPFgNpi+envq4PIWKg1M62L6YE8P3QkT
qh6dsMwxnlOww5/9QZ8Lu1AGvAx/JOO2ke/k43KvLgTzkB0CASGecPiaVjhb++Iz
mm4LiKaRuk/HkO0Xsd6+2vjw45VBBgpW3xOwC2llYd2dB/87lkX6DJ1F6xFraZMM
mIHjGlAw6wRheFjFNw7ucKmkpJJ4207QFmslNGYa5mW86nwbJxYxnse7KGVbkI4F
KiEG9L9S2ueWnX6JEmtCQfwpW0PWdDoziKcI6k5pHbOcwJvUq1//DLL2DCDSigrr
GqWdubjp3gokYITm+Mr/VWffkrYw43D6bC/4H5NOUSFyEjjVCr+GitEjqxpcZYpE
tfz6308zwniO4s/L+dzQVpUgQ2nptm7aJO7HB8n9dngeDWfYlNG8zJ07/hz2bZYr
xiimTonx48vIbZBnciXDhOUS5O/fV3RU9XTl5XfChpbZrdPKNrefOzCgQaBfP5af
YH25eSGu3WypiI+eUoY7yVYhmrvz5gw/86PXb9q5uk6833uZMvYADmWq2dIu3yNm
EuYT6s7d7ntEZkTSA2GmOfo0QzFhlRMTWr1g9ebktjziS2QJRk2CIb9t/vUkPBxQ
sJC1dtPNcMMRmqRlE62EscrH9WhVG2xGwS+QYpI3Xm1tG7z7SLcUPShKy+xaet+8
I/YTUj50+YGh0GSSAQWSVidt4kX4/9VcspaGZeSzNguNiEnlHt/h2sO+wdH+IChS
hsavtPlNFfnat1Xy7hWkaAcdDTZZjVAhfXwfE6f+lgMdd5aKv/al/HtcEH/6acFg
c8imB9u3NYw+sV8P95GLv4KdYj66BjL470l9B4vne725iQuYGGW53mYWpAhhrBfX
42A42CrxSOk+qaxVET7jln8/lmZHKjMtmcdkBxvIAg2zM2yEZlxETZMg0ciGyS6P
6N9J+X+lMtgKiM2FoZQnjtUmAmanLQdgKAtxsIWhyczFZHu3DnoqopKyldUCidwy
NQVKLhGbLown6xagXiViOSJoLp23JDhJjTwNwbivxQivTDz9nYNtLMMXd6tTWQWQ
dBesRiLtMk4kC3MfnGfwzPaT8qc/KFCNTrd3QKB1h8wa1XWz7z2226yjkhKYH6QQ
JMWDIDAexLMQlLBnRSc1xZTkCfgcvKTgWH/nPgPmgz8tmYhXK1Gkbau57jqsQ9u0
2EwXSzTIpxDGRlQXUcyZsit4iGm3DBrv4ZmtZjrYXZoN6qa1y2VyClFPkKQ4wrJa
B3hQ34rojVPzVlwHs9jrp1yLUzUQIuM3JGxSqgZUK6yE89NzT7EUOfKG3ji8wqRd
3wk11+d/UO26b55CvV29HRoldNa8EZFwxnBtxIYzyw6Stleiw5jN6sZLX9Ma9HKR
T/7uZtGnRwQ4+3Fc0YceIiLd/aSLJpZtTj6H/4NMLj069foRgaXi9E65L2/fVwB7
1wypHHTc/UH+SBe3un2H1/jjpdQeLKCyl1n/zfyJ92knN3IzU+l3OfQCLG+OWrkN
OtGjW7CliEpYM3pzhbaMCzbD2zdxCWACvwSK0F2x+6KxEqMC1180tjpylc5l64Pd
iNTLvbo//09sSiki3MHml5UxiCz+chDrEUVHGVdHzcKA9A3Inp0kJmnqQKbYEGCW
JYY45Qld6zoBZUBEeQBTvqJv8H4MxfEwQr2HFPAREJ5l86wXSAglcpEcBA86f5mI
QQ5cWi/j94GRWHjVpI2QtF77CCjH8BifdcknXHS6UmAiRRt/57uF2lH+qvdMLS/u
MJ/8uE0/9ELoKcLPf5MSFRVarS6+KqZlwqISksAcr24LXCX7Qa/8fO4Xr5kAB+J4
fZBZM8/ODTrc0cMjhu3ZCAhyMJZ2ioATpMPVzUuT11AB6zAXAE4af8CH6bnn137X
k/UtB89k2bTOvzlo+CdQ/3/tqT0oqL4amJaBgxJ1y3b2G9HUIMirG1CZCRP0GklV
VJ4pcGyeaGQVowTqtoMw1XThjLa77URQHaKeJtq/66suf4QvtPRSkg4mS58dDdOU
qjSHCI3sYVbIA9qNQyb+kyUL0Tkix867e4E+E/rX8H2h+EiQ3qg5W4G4gxaukCGj
e2UMR7BYGXRMHq9NKjkuc6bN69jJ97KCL59AkR2ycgtAMQmc96RPiuw57PRaw5xm
82XkOiunB9alCptQBeK2cXWipJWIsnV7h0HgvCnp6n0tdNIRhdkjBBfGAeqgGgOB
iNG0JjlQZPxqgsn5qGp0Edj86NpufbWkGF96TIWUwuYLRLrya33Rt0RtKZSL0pz/
mkYpEko0tF5zq7c7x618vlg/yhzjWPOVgwq5mhdWJMXhsbQzxVzLIh2dZLPJ2otn
n8W4TnLQEzl7ZqrX0Hj/cEBFQX+KxDlORjy/wYd5UIWsRHxNWHF1VC6DUEwmvSq0
AipuNf3+SWVedeYGaN3VhmYlTnMNXkkjQcHqS7U5UUgPcmliJ62o7zXfS736ly0p
O74U8/k67iW7YdbPw7bAhHw4ZWYkMuOaowNSE4fy+2UO813cCifPK+pfqvHrXT43
6JHnwQWfrBBwz5IDMuwZ8QQwuFy4cLFU6BOPFIb30Ch3WuXNqbiQcl6cDqCyBmbg
3R2/EJcMMEKit33wif5jwJSjApwXQEa7kGr9uEMaMBrOnnZnuWmvbKsHiQ+KnkxK
mTBVR438dOYceFH0N6+7dVUn+c/GtABUgOWhAMpvUfvp6gB4ju0t0ZaclXiqF0x8
IwBzBHRpIX+Y8apujMXx4FimRLPwYstBB1+Fk/ffAtjW/zEwyyVCT/V+3QnvjO2s
6MkK+4BQAjDNFpKzhb8SZ3o7Yda9XjDzX5MACSTO8bS0KtIT5DxLEnrHVU6LtLpE
w6PUEOeDX3AE1DVfCp1LlaRJi1GYpMOHR8MSPaCZ8Zh+4NVYIfw1B178lgGRlpOD
KT1r2CtzWs7igGwue9g90/m/Lrdr38yHetfAjfoVusr9fp48KYbBDaFVb/6ZaMRv
u8AXxK+JvRUHt+Ll7ohUUq5GENwmsQV5YAXGWm/Dpz5g2rS4qmSIPdHBV4+rs8aW
poDyrctSS3wog1w2/F4wIgRHbbsHzwsK6bibbzDK0yRZv3sQiQBxyz9W+lztZJuJ
MzawzOq+ooIFgh0k16UpglCRH1gRiSBe0SoIRNvBSoYG/0ClmVFbxyVxw1Zot8Sc
N//0vw7FksioDJDzupe/inGZILurqPM+Bwvf5YSRJ4M1JP9VSAppuF79Pbp3GPig
YgczIpC7v+7W0YdU1oPakoP37KKrnJHhMNJjv/ANTxWVZqm5ap7KHm9aaEjqQqXv
KKWMk8DpMRUx0b1Yn3GYMaj6AGyM2pqYUtFmLiDnJ5EHrKo4BAj/CP0Z9pZVSGtx
KURPC4kVWJZB88cCkvESzGA993PXrvnW1gRnccHKpXBqAPAenX83Qxr/fx+kBGym
/v+t7FQ0hZNVZTZStccT8BTfjvgoNN1ZW4DBXqikwX2Gyl6yAKXVi9Wpzh0s4UAp
uAFSNoECwy+aJlssGNpwwdYDLQu0S5FwWfoEby7rB3Xju67sNJXSYEo0Lj1yd4tT
lJe36UKe0C/TFu6NupYq/OVu9GMKPvmH+vRmBBEolAsGSXOl/G4PvY4fpT1cOZmD
rM70RCNS7R4z8v+s//jP1l+SbbeY1jc0JdaXmVBKN5bJXpwSTANvQNfupUBMJrst
QYLUbYPFKZ59ZHxELs9rzyr55S9qOre1VVB27IxiQZFM6t8sWIqblizrK76S4mMe
YJ+sK+gzoMqxs2+zUsvJhtr8opNHgoSYp+ykTTrRHMZ5Tr1+QN+a5VMVcLgnyDy+
0Q8Wc04C2jZr0MtQdDyql/FvwQx6SSxjaJO2NLmxijc1+aPjBpJReZNWY7IFlcjI
OONif2n54jwgFCadFuf1uE2c6GhXZ3U/BpZ0K3faGT2NCdywAr8nlEEwv1pJPfqi
0qk5m58gd5HNVENM6qQsdBLM0aaFmwCBHgokQdmi8m5B09ZM4a354qGu3cv9UhL/
+r6rW4wXhcobG8KWJmNrjE16oNtx/MUoVKQlTOGkigLJATjqZzazZrVkOyLlZEzX
iXrTN6miiWLwWMVYh+pf9AxAz7eMTkRKQb7J5rYbo8R2mT/HURZSCetBcZT1pYIF
gqfVfGCGb/5pyy+R/YWNCksZLx7RcMYYsYDPzpm7xMymt2C5vw0kuNJUlKPAjCtD
cQbxEVyX9SLCjKF3yTUhRg41iDO2JvJQ7+p8o1YDFYMgm6zUjIBY4XAeLrz7/A4o
ywQ3HhjjJxnbXqAFPuiA9CI7Jzq6OdnhJKA+KpcueL+u1tM0NV3nVSOU9vAZd4f2
It8T8n4mmQpcAQ4b1IjaZndDr+t9oVa1R7t35m8O52/wMbB7SFwN3g2NWmS4No7N
JyH5sf7TSTlcToxX1rzKgE50KfDFxdFkrX9pkHKnMe5rAOfCl9sODKzaUzXdmINU
T6QRVnb81g/uekk0Qps+MJpc6NbhqR6sjiJdP3jvq19g7UZIOhZGvUFPt+EiYd6u
7LHZNYdrzVcOr+4ukPUaI65Yr8TFDUbwhSDFr+qI73GP6msFODSUHZjAE/k+KQbJ
npLb2vrQjNbgEzZuBDsFWY0rwba+61banYaDk4eBieLLJg8Jvz7SdoE6P8PPU9lh
0tIWgRd2AYDCnPbY1Kn46js6ilw4NGzszRBMtMINBS21VItCuHQaoOzcJhGRVpXm
YiHjE9uCD+bFV45JwITMnD8ZSH/VyNcJWYvsahm4HGvbPf90M6TVX0VDv8RSLL/A
itbDjP64Kck7/84+nfDbX/27nfvqtSJwjOAUd+6RX57ihDbz2QIePBA7IPD+5RA2
+i8dNxF8IIbYNXnnzeDMwPQoB/uqrwvypCJEhcUucx/opuOKW72kAPh7MZaUcVCe
DN3/gZPoN3SlMkEaRWFMnAOhGvUUu88eLIsKmpCFxPeZIBFytEMspmfkJuntjLpo
4+RUzkXinofQV0pu5zLf9Pm1MQSWTiC1nq+c4boBlZbnMDsRT5X/DmHCawCsSY8f
SLS0BtovzkH7SvktwHpP3B7jR1kLiL9bDPHfLNEDkVsqbvGEOIoIGt3/rRcfDfsg
3x8L09mfbLbPtZ7LBy6bpM88J3hYIaFMfTTs3BlTukkHXyzeiH/dKYIfEJUkG3CC
x1djj3nVwIJ1MOVQakQl7slJzZ6bmzSgb0IrSuFvf3W+nwJTIpsozUmR8W8y/hv5
NpjmLbH1pTK5LVRb3TKZMQKPmPG3kaHd12/TAaZRTxIPsX6Qgio9DUKZ7ZyCgqlQ
rskcj0GBcH3ceOKldevNwUmbcPZ514fPHzI2I29cJqiqW1AcHsjUrGoOqsU0kiIy
kE5LLHWUchr0YK8D974z9EbCaHWnHX4SgygNHwGqx8kcSI22JEobS8FCwnQ4xsxu
j5Q/+c2xZzcV3wpzU4YaRfcFSh9ZyLaHsq1KoyLweZeJeVHucUkhPSfabtRgj/zC
/GgvLL4mlJ3o1YwTWCG9iTX+EjkEyxRhnWoknQPg1BIRLHVN4DwR0BIYl2Yn6Abb
vkZ1YDsl2ee/PuZW9eCkrusbqzrw5vfwW/PPMbwC9K2t8WdRNscoC89/8cMUbBZl
uQ4kv6rLTuykG+r0+JAAb33VQn2Mk4Ep/WRg3C7XksoeA48XAOW1GUjlTYUdj80Z
a0Dws4vzvx6Ej9aDI75NLaL+mV/ruWeE6Deya7MGmgWvPKFM+cLfyTmvJhJceapX
d4AQ/ev2dqTogAd8xGok4OJTpsmRRYTbFRx1uZ4mlZudY1/dMBUv37OuXcHq4i6c
AHRg/4L7ohYwtaUQvO3GeGE2eOjocM4W7Xd/UfXPjWBsBB7EqrzcyGH0+VvecNYD
E6BZb6jznfbcLeVVSD34y5XZWDJCgCzBLOMdTnQVHtSQ7upCQT7BlseXGg5Tj+0f
Y3aB1/sLCGA2IUmDppzFd30VbqLlfBqY3PtiBswfOh+0Qi16CnMIYV6yqL2OZbcf
HqXFC38lVNRy63tLcKTcJTMGTJ+wggWE1rTeaTikQR5PcVoU27Peb3+AmXbI1k6K
YpgTLqM9Cshp20XwUciilaGJomAFpNIaBTY9fSUEyWzUahJSGRpxqUKqySvTToUT
F3HdfE6/AAedXK4VFJ93knMZ8s96clYsoodl0KIBvv5yTRe3r5bJfd3ZyUBpMNre
6U/ke9iw64577IYZT72CS+bwfGBZmZz1GNjKRh4H3t18b/X8tihUyOOLOAU9WouL
IBgD8AHUst12AKpcIwA1o7oHFbFG+9TUN8pxqx4s6D7q6lI1iN6vnp+SaERCUTlU
6k2uytDlv3WuqW6Cq5boVRyHHn6Sh9JDuLDEKrcUWA3564BYRLZWrcg8ed+s0Ocf
CKJ5iB1ybuq3Mfr/ytUrtJGTgFM6uQhuvHyqUnUKuFvoMylWXXLc9ncN+NY2c3oT
gt++c9NLVotdIRCNfC+IOINbu6RegmfJsDa+ndNQl8RogyhOH6nurlrNMY23lQCV
t/E0fEAdsmVQusUj2TACB+2NmA1aimsu9B1/masCAbgDrrrC+Y+2kD+b2tD79ke9
gRmxVZckCE8YLgrfyp/reQpmS7GYO0L9+LsxGxbjoR0fD7rYtL3AHbxSznzr9YZP
oSgxqSZU7NCG9S1PEHyck76uyVkvxGNrtiDy8K+1vH1KqMrtWdtcM21lHiPgml5r
8P2Bev2F93rijq84NykEDQnbMZWLjWAAQgmM9JOAtKJ7/ssrSQde5+BuluSyb/Uh
Z3Kxr+vqX+gge4EBRXeR2F+5/79uDBkSAjmw1kpC432UxzifUT8+sFEY17bw2BWb
DRqGyFM+0/EKsS0LgR2s0mSJ5+l/r1H0ioWtKwWdZcgUpDDrgVkUoAvg+P+exZ58
SqveNRsohVCpQ46/gE7Dn0aC3cu/C5HHzO3C8E7MUSbzHNFHFnvYEU1X+2qZwMwP
bEB484n0LBOKgVaprSfPntG7lDj5yOZl/kljtqpXWUb7JvKMBad1jOuzCMS1Dbqp
/Ewrv9vIbQt+ioTDHwQJZA9rlwb/VMusOCIZ2tnzn6Nd3xcpnXkzYBN6+w7zuzdr
voivIBIbXbhpYyHMI7IwE78HSvXarVePfv6NKPRISTmVFXNgRysn+0BU2SDTdYGD
liPaRx+2rE+UJnFeDG27kjGm5qYhI5lCNgtDjKhYXfxtoPoXPxEnUtX2lMWeF2HF
/eoUtMpae25RVfKGlOOyNiGtwxmbqgrkShU90vJnT4sVjrNUy+ZoFCUXGoXt88rz
tZao67dp7CMVdabDu13LFgwWG8VDUldDgp2eVCz9CuygBfrP/HWWnvVFY1Qlr5D2
WxyupQZ2YI3dOAhbJALvSgCjK9UWtr7OSY3ZgTuPVkwzHOPk9+RSAcZApSDYAIdV
8XH/aziuFBKyVVQbR+LRIsEPh90hiYWK+x7GJKqShDoVlLoal18gM0GcWhYxYFG0
Qnc1UHwK1n73GbnjV5PuGx2ZDo61r+kIT6JEoUvf5zDALo3Jdd+vaCUZqrqUajeM
6L1cKYZwDuqhhYIbMlA5turJ2bI7r24g70HifxJZp+TeCBHk5SRuUteGIwQMPHWS
/+kJW/23EVQ1vy2zkG5D/hK2tRO+yUKzOaPlnpDYGggy9wmad7vL72XbXyvr/kCg
w7469sV22fNY1i16BkrbgjXpZ44kS31Kv38QF3NwzivASxLndbjOdBt9A2oZJ5ya
Ti5mVT7gZNrEgFra3R3VmOnWiqdZDSpgmLDlZElTEvR/hrv+Psjql5GqVNWBBPKd
r9kVtZyXOwiYIfNmTOG2/rXhDjr36awhmsFKJGSxK5JkwHopDGapiUUWu+9LDyh+
H1QjxCH2igNu8DDoPCDDMiZFFS4PR/uol0b9N5ZpFw/vGUJpgcRl/Y2I5LLnA3Oj
1+5hBnTXTVHCqzR3RSGeBPJ9QLo5zzWiAMqTRYlgVRoHojQK9YPcBYbMmim7D5l0
7ZGGOw1iEdOcsdszZh3HQnRvlXMdGFWaOhcKvy1WBebg7gsBNe1XWxMJs/4D5PFP
8jpn7iMxec9h4XaajidaQj96XAP5olMWcc2Z+FhK4sbTKQP+/ex9L27Z9FigErue
BG9x4mlaJF3pQdYtJsEP/PhhSif05jCpocVsXA5+8NqzXQdM36lcCs7rlIPq7UuP
I1gbKCsvNLEFg0Ur3ALc+Xeaheb7bX7LgXB547ftlzPfcZbNNaCruH+vwU16KMgd
+lP1+XfQvtfiKE2MrR2pcgwYtz1epijYNeTawhl7gAUXP33Gl75wVlZ5lBa2rDyB
XLgV5ZJc2bRwXWBQVfAdZtDcpcJXmLyJFpsEeyhAbwdY3jGKKOYx7SOaoYtthVRY
pDJViDBemwPYulaBm8SaPJRlSvcBU+x5swXctcMH1zfSLVyYdpbC21IOtN9S637s
2uJZnRyY5mEQ6NH3FQiOT/eQmeL6ATjtxPk0S9mkd58JqxDxYZ7U4PE2CCWrN/aQ
d/lvBWAhUhlcK1UC260r/P49RfFOMtB+uL+JA56e23sasZ2MLnOg8PRdcb8cDxvp
srctts2Fg5Xx4Eelho5sAo4hbmYMDTCu0bk/lZbBy69aWMA+uHFeXpfqkZv5aJuk
dBnqgA/53q2MvEOfLAfWOfDzzRwaU4hcGMJcD+fvmat7aQhS4lpWL5iljRZl+723
nQPCW07oCHDh44JUyKnCT845cCo+LLiFrBcuLqPWMa31EKT8owVoFrrIN0T5dM/a
PYyTwhksNbiyYCW3PXMdi4QK0sC/wXnzzVRR3BXt9oJ0WWWplYkjp7kGaQ7m2nzm
YVzzI/ayPQ2E/46gxYBiXtZ2Kcjd35e2+V7MFI46ATy0tnyWWVvRgUWrAvdPvV46
Bg/UNBXZWEL80a3KRBsttgfyr+MEjhsknEmDHmj3b3WVm7X+8GJAfcBLmT45DBqR
qa9g+wt5vKM4lL79x1MTyk6Wl/aIAoxMke5z+H2E8GmxkisWQ0wa2JrzlSoXGug4
ANmM6XH6q+WipVywXwNem4N3XEOFM8cZbjnjp8GHezkWeOorLSAzJKbiBnqYi3Ea
O/26bp/1uE15ToefjKlD8hdwkizB0mV37ADBYn2v3DbQghqAaZ7kMdN9dtG3ymDt
o+OOXmRGpf0Bmj9WnBMoMtMNJXhQhyjSyLQWV/Pcv4SSHGi2cnxqkQq57Uske2di
pZYacIOzFXNPUIRi/udVUnU9oupm4J2nUiaCBNryy9pVy8bKreoRwWqnNeiuKkhu
UC4tUM4mNS7dPXFbTEzwUQkufRDQkbKxiWArVL5M4LUQWYjeL9/vXZcw7PIHyA8C
kky5zqGCb8negqJu8UZy52idbC0rkzNmCZxAAUcqqRFHFTlFTYA9OUDavdu318oE
36mLSLoB8HMFnPKkXLueaMI/DIh2eZTgaqhYGozamLHtLVF5n6/3RYqkXNoR9ojf
n7OeVkECfGJjju1E7GNMLRMdEAySmjS9r+2nGjZuYUpcLy2/4cmwZc0qVD9JjRCf
kfMNnNPpGR/2YTFJrOlWR5+JZYlN/Xc13CKX10XZwUxne2xMhNRF6Zbhyn8L2UOA
RhMYw3vtlKQTmGLl2XUdWHbt5nHjWZTi83YAxoRlEeo80EpxlDaHxl1+bF54d038
66AJQLltc55NsRu8QWRRysiCkV6zpzljol38JWPRGxvsOJohLoF1rdIfRqflStvY
/8mxInPAESzQGuljqn1Vrvc0t5UKvTlfO3wfsO1pZM2Lki5GuI2snMsQ/vfAUa1g
pzHxP32Wfgt3suJv91to362KugDj/w9KbQUmBKa5nTsxltTpCRCaACcP2Zeg93LB
ntnVbhw6v44TS7tooHC2Hcp5niEPVEkCtU5Jo6wB/7CiEG/EkOdapREvKWlFPhmn
qKIPksToXiIPMd3vbY/uakasL9buIWJ2kDdwk+Bhes0fpOsuZSoBub0CyZGYkgxs
ud3kCe5zU/CGtRCzbuIRqaBA5/N0cnyIyyFiWwVhWTha/B0tGmAWjMaggIMwrr2e
loR819wN4hCgdxHKJotq9raKMvbPK5gQXhlY9V8AjGClH0JAzMkPtH/FNoh1C4/j
/VPXEtTf692qGhSEl8Ey+Q9El8ZO+EM+7NKDOkOjKwTkqMTfwZ5Wx2fFvoCUYR6c
PpzpK1spTiWxEuL/MDPGS31mLPKNCGuneQdq15B8vFgF3tH70QfXocDD95SlHfTp
U41OBNIbjfZF7U1L6zU1fVivNUN9h+9HI6BVlT5GMq+jgBVd5AQ3VmUNZSHHCXxh
TChBvzSowDgOzuQfKgL+qBCOYTp8tcTvs7WrJLKLipfKsNoLcK0v0LBdCFTbjQEG
WB2yk50TG54XlTZ0vM9eVyMpI3TZKrVqLuEVkVfOSEukJ4aEGEvOa793orHTcmG3
hhVjDJn0uBw8XvSahYaWT8ocm6FNUSK/kCTo5OW7Z3LqE5bb69RRpfD33qIMecnP
eo/Owx0lh8K7GG0p5UIk2feukbXC/dnlVj0hSCncrqP3rc/k1R26pNa45Cvmty3p
M/xNAVP2Bh+3aDcZQ2Eomo1coKnk/2QssqvlSP4wAgE1K+o4qReZPHB1ReO9oFll
z7jzlqav07eDrhcO+Kjjh1MlB25cMJChvbUWCgenMIfKf/Ko6IPA0XqKawk84QrL
lJ83R/HkjqBbQH4agh1SW7TJwRizdRjtgyhzTfeDWHATWPpmvzDBGKZ2/gA1PoaY
MeKdm+bTAcYBlsll3NelF08LglDIe+aiwf2nRzJEs31WWmOHsS+tSoUDAxPFrQ+U
FnCWi/BZE4Vv757BKSfxrDy0SIPqhRiTdLw+BVrbhd6a9kqKB7raqwzkitzsKr0B
CVJHNrpniM9B/QYbqr6wwhVj+YXBbFxUp4oB/TGHQc5ftkyEBjq2SDQyuafXdTxb
B9Ql68JTqroZHAJYiKAz0XrqDX2KilSVxfpHkULaMsMpHYa/P/u5TAP4Q41uXP/2
XgpVNPpzBj2xRF9KoBN2YqncSu0UDhvjXdjztsNXvT0PTPct1XXKoGg3rThy7peC
X3d0DFyM3Sc5X7gHg7f92RRPwLoapbyEawVAWyPQWR/K/oZoMI4pKtb2Km/ZPHB1
euV+WVVAjvQR5W6xCKGNFs5QXM02+XOG+uA35ePkigpc1vHQuKfAc7phRdhiwtvI
vaxwAenfARtmG1o/UKKa5F7NLAyJ8vdeFQPv4N2hGSuPtHEk2Z6Gj7ACFGKVYWB6
DsPkpOJW/uDk507TYvICObveV2IMfxjwrRzGApjdiw4SSo327DaQF7IDO1u011F7
HdsVWHUrhX44deCW34qjb+fUQZ27myVZuZRGXrq/DQyPP5bi0JDAzzuagssW+G8B
e35r7WyQfWjJMYJA76aWzg6fEFNS+rMt37qNZlsI2isJ6Um+eIFHTnvk8gSKoHQh
MXos9mxFfLuuzSvc3VOntt+HGkss9bJim0tLk5yxthxYINWi6jYhXwJ3oeZtgot4
Cex9xRaNrSvFElKpVsBC4qoFegUAduOF5jgm1qsMRfQ1UVddGhP9wsrPRBhtoI+u
Fv19X1yx/ejBGqhyDNAAKkYxnfkqmfDLHP9cZajaVfVHUGT1vvHvlc4q+Qqg5+ZL
CftmgRu2hhFu6PKXtKscFiyIXkJM9Fcmc73o6n5naaRkSaZfQruBvAVmI9PC1vVm
kTFPMpFAXd4JjYUuM91btJhSq6AGgbFCLgmBtuYw32ArJyrp2yy7CdMq1Uuh7X8h
U1bRmW6YQocZq2Xey9fhd665RtnFWpUD/0+jb0s3rl+AkrloWjJf/80Hg6XIGQhJ
DnPEGSIzR1pv+yRih0eG80QS7ux9X6NCIc0w1mMinYutptCNApzcvxhqYf1AJ3s4
1vWwVAy+JYZPGFGqC33MnskpC6y3MoLe7LCsQfvMGwOfAv66kz3O4NMrZLtuo4bQ
mHGOXcOo/0axIVmrWoHXiEJQDzN8M+cHcc0jg1yTfFP12u+LAVnn1jTpzq1PFJfl
3lstO0jw7LQikegv38Qzg4V8haxYiXkvuybna42Gp4A4xswQssG49YiucFY9Hqbj
QkjTiobJsG9BpCf1vIAWrMVJogeLfRx4gAfXYWVukDvhW5imX7KBsln112gSMyM2
Kj6OITKxivRvax3MtFtudXUuHaJNdyhqyu4AwDlMWFuT6mQ6UpgK4tbS9v8JtXVU
Fx5iXqJ2CQ7x4sC3XPGX3epF95Pg77l6jUI6wP6pMjg6RGB+uS4+rGVTkN9sjH0E
QYi5s7QhOjZJcFrNIs60gUKx4oN/GuokZwjPUbaZmcyp2jn9SbCaaO/IBALlI4op
gNYrbtM1HHTHIXPqylCWhJTZKLg1yg5xxSCbYbSgBU+PB60vk2ns1sTwT+SlEgoO
hht7YwlOwgcISxJc2B+ss+AUWt4vS5FGuBKNH8h33LAdW+BLYdd+w18gEo+mBpvY
8/ib1yJdeay3eoInR4QJKaa7ujy/Xb5CrOWCD/vOzYJr4broSH0OHTq0FZVHP8SB
DlNFurIDq50yL0MN/a4WO4qtO20xDDxMNgh+SfDRKghZlluX8z7d//fLtY/Xtzlb
L2tMFinaED0vsTTbEJMcr+hyNnbLkWgSV+Mm0rQsOMywjxLPza1VT1h/RU0tOuBb
72cjq98rlc2z8gei1KIyvV2SUM57OWHvQtWjVWD8pH2Nc+wIwzmZ5rydX6uEEtzz
PeAJi3Vtl4h7VEj3p/UINTxQK1dDlSqiTMBn8eSUaKX2+Vb4yvT6eLK/2hWDYEU3
NJ1pCLVF8iiWTIV1tu4R5ctEMi6fZVakn85HDQrJkXB2COD9KGc/DL/KjpLzM8Xm
AVff3Jo6MgDIwIPd1Z3m60tUvvlhHnLTu1hDTAoEC0OzFsfg7OaIcSXQW4QEWiuA
ffghZOmfKZOIjlzNOpsCuIWH+Hc7rnSJa6iU1iY7xXA71hkUhK1u1BTRTrA3XWTE
TFNQSYG9E6Bjen4G31MNdnxI/HriWZQepuCU3+W55qYaXDN1UbDYKQNZN90MkOk0
nXjLxJLPm2Tk4gdADHxjoZmQGy/CfuutKkUbwyiyZk1Tuy3RQRLnGXcEXBLskewh
zT2Cezo7ozX26OzhRsg2dR4yYH+EnP8HvW6v4/7dnWXiTUJQiW/xpUv+d1VT53QE
+Q8RgAQ84oxy3opbP4JNccCBUm1zY5HfuGwWZjzjlW1EHpKLPKbW609GiWFrxtrm
oxwE0QPCtylaREGDTNtIlbDGyTOe5vK8GmifSmUXv/dqJ01b+qHF2r9MF/wdCfvP
1p/bpGugmdyAQe4L8L41IKUc8rCSACJQlOYya8BeHfVgWtGOgKXZ28316laUbCEt
UEATnaWaMlH+IM5QQmr2fGtWmo+vrl6+++oIfDa1/YaiyPBV1jU7BTX1QbpZd2GO
1pCAASIUAhm3RNoquisH7xLzKIVVbYnE0E5Awt/DcbFbXn5lvmM5nqd5oXYD+AuA
tmAXouGR2XcltQTFt2skRaNymT76G70CDoDdgAQd5ibRmrpSHjKGlvnq1wEAYBNT
myog0My5SeIlZKcEjQObYQMkSjbwR8EvhQD6JTeMcqbvcpt0DclSVuXOqcCCTbor
/+dp9SkPLFGuuagQDiq/66xbT3s+a9zw3K2mk3iXq1uLC0dZDcQEpvDG6LChsJRe
0SzYq2t8r8ONQR511LLFyXQYB/5FapxKVaIruByfepMQdrQpeAS265101Ib4OVvN
PfoW2pXdrvQMBIWUTvWyxvfKEs1iy07FVEaVJD4iJCAldkeViMoxDhBFAfGDNaJX
hIpcgZBwEEaMuAf2VvJcPdigT22roVaYXDME4rQ8x5aBou5kDMIa9+RWV/hxWklj
OyIpF44mqhJ1wYlu6HhnykMtAYuIwFCzqvocqbsiWngShtPpBgUx7YGR/mpDFlrO
7w2r1FoUFnA9bmw/X+apppXAuN4q5LjYQr+uUW0OSp/gN41KXi/Bcp0Q6rqmE9op
m8nNV7CSZRN7iBbijfW/WlHZ0oCam5bXcDe7Too0iyyuk3cxfHXMa1lBAbfGhpqr
v/4PuH43atZDFJwthpAiha7SVhDv7AfmI4qS0owS5vRRM+heeenu4b5U/6H8+v32
7I84Vrm9XG8ki+hX3oLxCeNlyidyc7CYdjcOIY2kqiVzBSvtUFhyTNVgnF5Mzix9
O05a521N5qYX/jEAbqqqHNZVPPuZyqU2q+IgGaGcp8Dsnu1Oi8FdnIJOclhXSSL8
4qcPXLbQ/0wCMyiIG/6EM3Kmi+bHt4pVEc40aCs5e19t4+zfxmZ7SWJpms7ZY18B
Z4jHMmFSOOHIVczzyG0I99ehqAwQoBNyFkoXbD7VohAT6OUthNO6zVD+Pw61aBak
yYaW+yG1stFehNy9ViEPU+9ggvgQFUq98dZGbAgErB3JszbJPazTop1cXraEHHB1
EE7gujuWOm64wtUnEOfOrH9OQoH5xeaHbZl1LiZggBKEFn+idfD0ojmYiiZzAvxX
tYalPqs6UaM9pchY+vjzZLTXmkQ7NfRjwiBmKXtA7Xr5zIOT6MKXSL6708IXxSPW
OIWvmqSMj9uPCJdgZLDH9lTlRRqjQBTMzumDW/n9lLwSfE/TDMAYRcPC/hYw90wr
3nr4W1ar0XgXLwbCNgHn+j7KsYgTc++3yCV87p1j/0NJuag6bMziVNsTfTR32l7D
A8B4UYRDuZfCkqKwmGltKNta8yWDUVyBQp+bvj9mTkZWOe2B1Gx1OfkckCFQZRX9
TBkcjaCwFhsXxEWx4xL14udZJte/nLxzix7fFzH+XbgCdeGvwvL7HP3A19qy7Ini
jNWsUfepNyZj7LBlkdZZnTSZj1/Jq9clholV9YiQk9W5hPJ4+CpXS/aq6q+sF9Zr
t4sh7Kl4WVwjlIPoVl8KEnrXTzZe+H8v38ynFPsg71c0NUW+2MxEyp/xtSA6Owh/
Xdm1H8O/jbyovms65j+QlECsV4IhwFICD9WqoHqqeMya4plgkSslazybOr+ENbLx
LAnz2Gu5jkblsxNJEaNHv4LLBowcjkdKDAnv4isOqJlIFoUy/7Mo9YRifyPNh+Bx
h4Fx0rfKlqp0I91uEAIJW/9usa1aykfOh89MjfnuwwL9yylVNsHejani12Weado4
9hHy49oGaL2dj5WXXeVlNtnhrhMnWNiwxN6sZ43G/8bKx8IvrOGDlRMC0GTto9Rw
sYtbMeA/heiA3JRRLFJxP8N27qrDyZt4EPPFgmHHwtLlEXWvcFLOmfMYCxjv6bbN
yfW07RGMV588mVrxTwVxpMKLXEQTlZHeOJWKNkycvxKhdGn4kxCnBB5vkNHZxiUE
RBjWIoCR4pO4RbJFXMPJQvcIflricYcjssANHoG3wytyO5ySVgDEv9+CxlmDeg82
Ycrzt5InYTtjDhPjoQveLkMFpgW9M3PAZzUvoFbXaAKb5yW3YGRrjGAJm0Hho2qe
4o7xvb+zYh+lKvWiRvz9z1CyITwF3u3btymeEjJI+hTgx+Ao3eK7wRIZrs3Q3nVa
LvNh0PeMD8gDcCDaL7kRVBMlgQ4o+miPCh5btpom6zSHVtzL+i71nk1IbkhhPY83
fFYzl78fuIeMTfbcN5c1n4LM6Bdwgm+ZQMLjLWSLS55sLdZA76dz/F22Rcxtx35q
yUyI3dEVQjJ6CLMEYbk6912kUk+2n/FzjYE5g7GJL5+FjvQeL86e1xDA9zE/nufH
KY6HnzEapAUxnqMZv0+fPazHSZTSzxo8FyyZS2j4oPjgdFWxevT0OvxA/hCyOMiv
M+T2VCkqbXoNz71FP4vXz2auSMTdlnELlykbe9VA1Sx2hrtSwQoDwMWoiDX0SY9g
NgHlO4kCr6JPltezncz3Gr1KXUkUmvyWnTJHq3dUT4+PZ7AIhY1d742TdxRTW8RV
O+D9Fe+oMbqhN7sWVtFdNvtv9zxWUcqCWJnBDaUwee+0bIDD4Ze/tYSDQXjZjs9y
BO4UrmfSrZmQnCUqwh3uPkkJgs4gcePJQQ19cXQqayTqSNqRVDAmhO3jya3soKR3
JiDRLXpvR3NJ1BIop9jKtfhYFxqQGhlRVylopjOmAHLsZeY3zEEqt1GMF+nEfPfN
D3lD8BHiE5CJtKxX5MRVcar8IPGClMES7E45jUh5Kgrj82bT6nXsgh2q+rg09VIX
y16FeMVNsuRi/x4g9xLvcDnACF2kfEC/QJjmSBq/XyquW256jyZ06tS5t3AqdT5T
3J2JMyeORIs2EkKl/CSvT88l0WRpIxOaQjq1anRT06I1kLlnIEbT9XZjmS1W8VSD
4VCDbH4LNdpgywzhrJb6RnIoPLS0g1Dc4GlZY6RB9vhIgbFmUwSRMkwAsm1Wc4MZ
6h4ey4w2BVENZLIMvmxPLmdnwbP3W6NvK2jZwoLvGvPeLyUJxtge0E2VA5W6nWKD
+fv399I1lnZ4fkN9aGIVlbCRwf6n+bqROq7ZDZ5NDDhuXMYNnYTzuD74vTyg1zDV
ApSeExIm3vnLDorUaILTImM4Q30SEtrHuuG3Wl996KhiOzr0Ffz/1IuZL+Z0jVe1
qLkDg88c49gJfnitrVmE7bkRmRKS9j9tAu/cqjfqBda1p+3T01iZciQJNDDOmG7h
hfU7Wv0mB5wfYpE661JyXm68hsXr4P2dZPzYd/jdB6h9K+kJkw8xVbfiU9L0Isbo
FLLSXEWYCwKe4SYtVaCXJs1uIQ9iwaTRGkv8mm8CaaDagQ+8W2hUyGOZ1JSMYmml
tYkqCwZF/eHPhs33k9hXy8DwSQOfX6itwPX35hj1jvrORHYXfbL5pKUPckfXO6wu
r/TSIypJV0c8kZEL42jB1FN3BW3G2raLfzS1YxuoSPAz+8rA/GpjokryTLPb0h62
LOexdvBtU41FfTHVMdwgEjtUTuqdoHFVD6yVF1aoJNSY3wzwFei14gTnhN9xWo5p
eEXYUXuOsRq76K4pItS1UD5vKm1u8FJhETXFpoxIDmZs4GUwhNmjMjiuLgSWuDX/
nSfhaevCJk7z2ApoVfa3qggClL8QYnn7BOe06uaLdYB5YgvGKck3MFJ8OcFby+Du
AyfUMqKzvzmaZCCA6j5zo5V6mdlARnbstF7TUYHH9akGULjZQbbYPJ/cFHlOP/ND
LgbC8fOXJP8P7yPzMk9uKpBG60DkzqPSK76qoRDuABHtSwTAMHQjo2F0znfXILgt
QFkHWiatmm+msPmdRXnEpx42KVuWqGmC79EqL3pJUgvuzf5UZXJ1fYlp/fXphvEO
EqIWepELDz4E7tl0edi0g46qmANq3H8SIIwzwcatBGuCKzK+77RlX0WQ/olwkHh0
+jRX9kP5DdtdLmZZupSLGADRSBVp8G9f3z6Yn6Zjr+5Z0h4BngoaYP33ygOAVRVA
gZ5oKF40IrzYieTe5KEXeLp3SGlxBEMRk/6GewKer+uY8yXzTMllvTiogVdJdiCo
OkjLuI8LkrPXu2wgXl1jvnBCXYL559lvmnqEG0jxWxmU2KHAnato5ypfZYuzNnJ9
jhkljsfUiVerGEUDFjxiV3BAWXWb8SWISeZQ37NQIO2WWaewirIDTix62OC10yJc
X0ukSDfORVFLivkxER2pOd6CDIeVFOTbpXL/6evwhzxNleJCMRSp08+mofE5LsGq
gPA3cdSyWGvFZ3BW+E51JwHZJi/OzWEcg+nDg0hJRQJT9Tq7SsX+qfzPieuymNTL
romHGLfar367zpossbTJKXQtaXCBblonlHhxNiC0VTdraluX023P0xNt/QbtMwB0
pX0lRSk6TCYhNtRlFfIXCddg5zoN/hpGlgzegSmK+TJ9zoChh4K1JTcJmYzwdPsl
CuRnM8N1Z2EN4ZODJQMtppTZBxDGAJq5PYTSPQNa6/uxVpG//m87+hPD562DIPlo
MpmlV9L5a4huCmjhvvZ/0rxTxkG9UA/3aWcupk66gY1XZX4lw9/iS2bQPIdKlaKi
eDur9tKdPuvyzV6+rtkq8RatPQUSdZwYaMqF0aJ8vEVjKRPfWSvIwWVpaOKx2AVu
Ik6oWiP6/1bzeGRjS3eoDMUB8JySE5PpqFpzSwwYtTmqr4KAYPATuwPutKoWhIcf
8yJkf1z8nC+j68uB5Kr9h1DlElD+aPATwXlO8nUlzMF92h1rhX/65T0JDgd+EEoX
cMpNZDP34iOzFuUf+Hzwqi5XIzjKQgQjtuPhHa7Bh8PaLDvQ3ESWfHG2mDVRoe9Z
XH/Bknr2fbrCONcHETDedsDyQyCTOBJYhU7TtqIkko/n/d4MSUmeuaD/7l7HnNKC
ox8rXEULBs32GK+utYwY/M722l69AucyLxrmmHw92S01S+1+gNIaHFIAGxW9ttEX
cbA/+Mb6Sqwd+m28OnI6IiQfbk/3OWtFnNs4sHFsrq/i3e9D4kvp/wnqzIo6/gox
/X4VhwQxp4tkBrStzh7tCsPHKW8jn/2N8/J1TF8iY/98kFcjYxwpTBpyAtuIVN/T
ePvEaJZ96/5JRIOzSEqDD/vs1E6ZSGwBNrJDoOoELt3L7wieLID4VdpwAydyiRzw
uYXKnbkKCEe7DxyJk0Mt1VEajSKxA8jbifnNzg4usD+Yiz6zgL5RhjYyQ6xcynYH
1cVmyM/0VXOnuRrqBjSIAbPzBUHheagvTo5+W5OVJRfxba1tatXsDO37fNwDKzyW
LBIK3h4JKodj/FJNz/MtDmgd3cZuuimskiYNmyQNTBhLkmiz+WTj3N0TOUdKPzDU
6CfM4T2069F2dYz1WPXt1gDod1o7AVx1KXQpWXBAJyFVFhphg5v5kn9t1661iOZW
m20P4G35FpDnsNu3WnLcYi/ABxZZt4j1U4LkqJ7yxVPQ43EpaxmjxuFhhs84djka
xY7QGHDOS9A1t5KD9cyi9u8eujQD73I2k3ZvypjOduuOBdUBcm2E4BWgLZup+lm/
oKkwEfvgCf9HXMJVlRbA/8u+A7s6LPQAaQUZOk3gh7ay94QUjNUQIFsf5GE4uhA6
TU5wiK8+RAerFd+qGeeNRi6YNGx2S2LhLY1HqbRnPZwGR2ZQbxZA9VUPfURVEo7c
HTeI4NJPy2iUV2L6spydDbWJdsiURgSE/dhgXaQx7k0OzNmuoSdHiY61oN+YJwj9
neKmEu2I7TpFxD6hUK4OilAGxQQ+V4r5w99gQxKuF14/w75f0kHYdFS70TL3LyJ8
3T3JE11BUS4JEovwCcgM4e19vZ0rWrzkYPEDVs4Jvlvx5GwOHU9pnZO+IDXnxEQR
w3H6CePLDqLSEh1OjvEn/ipmldxj+SLHZSpeCDI5Ssk2JZeymSrNgp8c1c1WIiP4
t53EGKVAlbocyFJOzM1VgeSqMmbVsOQ30FZ69/nPs4ixpHNmIKEZ16KRgJ1nEsY6
sHarU+MBn/JTFFCgFJgm0UJf5rukxNB/SsPxSmNOU5OZ/jMXOI2Y35JszkUC42GP
GDKF+OyMc2slr8yuuFQTx4X0RajV7OzqqwdlV5ULs/VzfOl45p9bFwbY8jTSSIrO
B1KRw0iSkael9s2IK7v6hNR9iyv2JcZKqAz5/Wwb5kcfc/IG69x9KSRH2gbRQRJb
9cmmHLzi4cEPCxKTnXp3cJkIk3c6HjhMNhRMElEfQ43B5yxgpjP7VfGFqvLxX+Q6
+sQArYlfpGKCe6kj4XyO4POtvR8/Qee2+3Rm3KmPmU7HCOqaVeXdVvXbPix1Z0vy
HUmE+p1osXkfKqu4OVMFKENL0u904yu3Zm+tfd7HU2nD7B8xgKcwafhi0/a6tRSI
ruoXTO+MoLLdnTAY5Si2R4qEN03gYYR6R/diK0pb88gie/k+WFpAPCrl5fJUpXuo
PzJ09o+DB3MKazvTwNLiFsUEaO0pqyRQigYtrn4eI1kIWkZRlTelEkJNl5h9YDiP
Oi5S6PTIilLhFZQ8NmdireWYULMwFW7Y9b0pEq1SbbYVPVG0n3Yrp3bFTdnjksHt
gH1THdB6b3OJNGhfe4l0PiCBkFlop//WcnBvbVzTe/MsMQdxhrNmsO5Ybr8ZB6xc
PElho7XDtIdvAGSqwR6wxfmou3/v6r1daADPxK4TXSw5N2x2Ihpm6TNbAOIyW58n
j389YUTaVNXXYeB9i3LCnTmxljUtfycIXLCcYj1FG5JWPwbQmiSM7cuYcp9mh8St
xIJtjJehxz3Fk1fQnqnmJt1jk1caE5rub4PDGMATKnNMeK6QWiFWSc3A7LouEhuO
dEJ0GOo0ymAMalMPF+fG2qiet9OVWudt/b+kviLY3lyoGvuBf+J3xXjtVWJlUFRk
/EAKRZ9udAFdx9cRmE2AHi7uc99UTyExWtDEITmJR+WeAKg4aH/kbxl8+eTuTai3
DwJteW2JoAt0AjwnGpJ+IPsjMD/HXxsLraBVv8WXldlTtU+eZWzRftP0h8uG0lN/
DokU3HZAzZtGbHp2r4Xg5MX9GK/Lr9O9AKq8cri87vfaZssCMGRX63K6YhnFf0qY
YFz7w6UPwKG58/ZfxcrivcLxJfDz4O9LQNGgI41VvB6zsbF5z0G8deZxmzgmazcs
5wWukkUMWXUnf/WJjORe7lKZlWvD/dtQ3+UdiV+lChCcBuBXjQq72x7TQpfLZMlF
ew4mvVgouipxIaLponhi3QCV4sHeH4xxuHNQCILrlFC1DBFtF7BjL6H9pOEWP/E1
TbJCUD86yjAfuF5YRx5oa0xRXO88yn0uWkDV5+SCDtE7xoWyvzFij2Srs7jZuVu7
Lgvb69+hnbPcJRP2gf0JAxI+3v3qP+9jDTt2hK/4uk0/Um/GxrwuCodmp4I0SYyS
8tcRW1RpOiQDc0D9jN/FMOeHAbH2oWg6QFRmWNtOwcGv8/mC12Iz1lO4QUIGCIDp
vl/CnwWrW0wczKnA748olCOt6b2v6G9dx1yYWKiolmpqoFMNJn9QyUILLVg4KqBe
ivdsTomQTzOETKs8LI1WRnd5McUqO1z0jgOb+mKQ/bjTCijKlye9MTjauc0p+Sa4
QrX3MnpuS4lBjA1PCIC5pW9GXnsiZSzBUQwZZCMbw2NI2how8pxkm4WZyE56cD9g
egqEWzJZKNJUlRI+6gjesevvx+MDd2HzvnkYe2J4qCTsFfvD6h5g4LIfWohcEvVO
Dfs54EY47VYtgUw0GtbZdDwjxkVoznxGgX/xJx/eoNMiHxr20hGpPGn3IKIShlgs
ZxsjGtJ4RnLEUn16RdFMZG8iJPEQQwdFYcMjuyGuGRqryZEMetAVOM7WBo8jLYyD
Ic5yFZgYiFJQDmp2UCvkrwVFj6JqZ+ID03qsoKXcp9r+HPV6FJLP0ZoGRlwd+Vod
Q1UATi8ZQwCj0cjDTn5mcQqE9OwSLNjGj72NeGLWvjbsYvhF/3gl0vMF/BpHxGEZ
+8gE2/sm7JWqE05YXvPsqpiNas0+sEApKzwgbAvvD/QTgN1araoaxfNXb1bUAITB
ZZrSC57eusNj5wH2BqbkUB/7Neqx0C3M3K67deltG2JxtIY1Nj2mTaVUb8rWaDwM
ZvIu2LkfKiiuld0RyOAg6kECaDKwVmFsrqwgATFklKXm1KOTld/1fJfYLCDg07ih
ra3KCX6rxmomCwMZUg3MECd4oZC77QrtCIz9yGna+GKsUuq1zihph+7rkx8Yc7St
G4V5lB2Yym4vSzJF0itaZHHMJAO5losismSyn0yt7vdt7IekJxks2kYebICX9h8S
hH4knajnE5oF1Vv8kGt5wYeoCk/3VWF1eQaZ8DICtGWVPRtn64TR8xbATgWdUOcv
la4kcL1uG30W4TqLxKBZ4F2H9DxNNwy0zdZZls83KcXEFHEKO5RZ2nmhDUeuRhni
0J+2nrDbAy61Y9Ox10AZ4O0hlXkR0gbBvtvbBrC2E4b9dFJU8hsdkT3L3D8ufEkW
+uWaWtY6rybMeeWa2laDJCa1gTqxS/gprYse8irgD8rT2dQz6ViXQlQMPK2yF+cM
UL6fMMOlRCi7UD61f5scIjZQ5Q7tGHBI1K99XvmlgcOD61dyO09ZpapyY3LLSUMH
z/7YPT6+I3BVrOL5k6Z0YJo4odwg10R/z0JFUjBQAuIBWoG/FeTpQWH2GpyQd+7R
m8mLUrRDeZZQlI3dbnwHAKm95npD+y9BM/TaYbj/N8tHmnNUsTQqxiK32O4Bhh55
NAYe4E6B+wAZYAprrRlLDOnHw5iFKopdHByrutXsGkrvpk5UjFb2LguFKzYOBiws
RDdX6CsTuVjPrd2sTEDWDE46yp+MroZZIfn/DZfCx36XIhzrcKgRMRiY/nf57Q6E
7cuMHCZKfmaAb73xhxoPd48gUIlCgYlyBElpqPdS+AzmOwntyMP1lDDjOUA+e10t
JmEcCUrVPVi2aNjdpE+y84YRLhq7i2C/9ItdDCv4NSgavofJFoKOWKfPzdL8KJC1
Rrhhhxy4pvwf2qJWa5fhb0qDlwHvqBli/a/v5egZAlQFziklPXqNHfMWm/ECzZR5
JVdioU+E7lhD5Jyv8NECX2ljVDAEf3pGZYIwudLKByl0LqUR9bHjV0E3ooHLOfcx
t1QwvIQUJ2WT5vOSVoLlmXsTeYzhp4fPjnq3oSPXswcsIdYZbz9rWJfAmguQcnKH
G0jHv/v66d1mXt6YTkrx73J1s4n0LR5phTiF0U1YEw3ZsZsD/pciXWg9WWUPYEXb
RlAO11HvgMnMaI7A2TRnVQmpaEDhzj2e7hWO+28NLV7v+13uAXCr9YJDlE7f7PVK
9VdOLsLO11bFyQ4mFhmhOZmZyn4yUe+uW6d8pV/l2mfw94pR3urb8KFr1WEKFXwR
RhQGPDxTfO5Aj3q9XI1OGp13EhXV5P1KZxm69RRzpaJ4bDBD8j2/yzZhPNNda/7U
is69aaKPSxZjNlKoC/Kp6wjVt5+6lurrqSCg69OiiWCs5lL1Rf4bqntI3quqkMoR
niLGeLDYkANw1Y0iRBxHOkiOZrKTBLgchokbNQSDyTyg4IMLvnPy+ophUnWEHnf7
fXWcpe4qcelPD9jvcBZUPJnqt5wOhAgAAwYFP2U8B/+oU2xYC48Vb74+JgqoH+pU
UgKQibRGfSwLIL6pWTrfwZ64QA5bNCobe054XXkP4ItTIoPzNHpHg0Ry4z5xZ7/t
v0YXvD+fbuNUjvgjQnk1cP307cpaMo8uggGfrPKSORaa1U+KS7VRyNOkwUZ4o1Hg
ZoxjYN7avCoTVCjzmwomQn7AJawI4Zsj9P1ZYVH6pvp8dKFv2x2l+HCpRgjBsoy7
vuuPPvr/Fea5SLrY7IQ6ogDiOxpw0r2Tqx76hmYhHjtNly0GfLB5Y+V1z6+lhQlX
6l9fFB1eYfetugD85wo+9oB4QHXDLi4tk/1MaBODK0iEPwUItiGPN/DzzZkdqziP
g/3hvz7O+Sy5EcECNN9WjYvEDxbpX2//10oKFiNDWpNs7GZGXrqSddk1kIm/WDET
XyjeMea9P8AbidmkruwR7BmekphL42TGTVrioA7IJdBvh8ETV1NReT3DQ5/1O9XD
W2IlMnv0EM5kKUlI9PYvKc/lB/C1Yxk2Bjx/WDFnDpe/sOVBykoSb72EW1plD9v2
94te0Edj5UQoPYOjXIvrnL7CXSEkB0DfDLypjKnB3dYVq1ELwARaJwT7VrcHNnuT
La4F76v0UpDmC1o4zQ3fGclmNqTnFB9NSCJ+dWo1WCd+L5wO0dhbvw1I9BWdVPtK
BPzbJrqsriP0fmzHT2MjEdaDMZkUmQ7OjOIeaXKnnU8HwiDj0eSLnbTFV/AoSnbP
zlIz/4sPuFqg7DkdgUlCGhmgjI5Q0WwClkXCF/c6URqn3MMivyp+ONCbgJ+Nf+d0
KHN0Ev0tKFAprH1M+YgMy2sSm45BRjmreRJk4cf8fYNbKfFASQ2y+04ahtZetth+
VJDA2b6pcuuMYmlpLfJwMWLYMVBOGdZGchWsIFjUSxikFif43CNhQasc/bGznrT2
acYw4Exm6EG3PD9nktP/3RErpJpUai8H1xTcVvj5Sp14hgEOALubdME/1FdezY36
IxzfkcJSfQRJLfEgwydtWx55TLF60UkKlIb8HV05VDRoxUjsj6ZU+6y1WjxpOQto
biI8rHwj4URNLQs4PUy1eBx2h+5EdzZTNN8tZvv1OORNBNcTu40XRjIGASAbg9QD
+eUHEtGKV2iu8xNiQDBHWhk9UFkPUqqGWKYu+G6JwS5IPGerNbJj6GzqLuQbYpfY
qGAnihnsNswV06QG+Bl8h+3n8KHLfPhyQ4wH5QY4jv/j5xKzGq89ifWRtuRYytNO
WkmQ8Wl8wF2sLe8SclMJBI7WYc0lq+ZZDw2xci0TBYFM1uyHh32o+kVueKjl4pvu
Pgm4HMpZuqqgHUdGb45U4ZRM8CaE3J/JFdp+z6VDc4XTCbsYd3Ibh6eoMa0tFaA/
FdioCPvAsXsoBFp5rTOnJlbXhOpNLtsIxyUVwquS/qCo9jYplZpEQNkasv/BV4w1
IfqyMGd001Ww3e7+NVfJS6Z25UgXpR0Ll5WfILzEwkocMie7eIMPgF7lRsjpyMi3
Z879GK07kd8G+WYDXFk53qJVV2wlP5MyIhdHom139CJoGRYvrm+ONJ6EmNQH5NlQ
o6B7aWxgAHRg1PWceSYpXohQplToFyRaojfR53oZsTnUVQO8qjDe1dLU9t1szGBb
Vy0J4zM3olyydwiYjL/lmKceXcO9MzVtgCEkNtroq30ZqAosV4O/u5t2ULlf1lNy
S8l3OfAYwECSvwa3GWqI1xsGxs1T5VDO1NlFFK4dEVmzLcYmoYsaS0aqyZl8dnMM
Zuywvr2pwjdm/+G/4Cl9CSS5OIFCciu0ko56HK7qByEfCg7RAX5Gq9l7HMvQTT71
Y0Utl6zetCEAK97f1FQLr1M1ls5qp94eJ5TOL2klFav+MlT/mxbqdlmhhxZyq6H6
DQHSbTzlHJsbjxgW7s5dFDdmEVcY7feOSx5m7nOUmB9IBTJj3LhKNSgtjmSAiWy0
RtK8tpobnuAy9zRFOWJVuItCw6uHxBvBsk5lEVe8xq5ctLkI5DjynCvfKin6MvEX
pXIx0a/6RQW0tnxxqqAWh+uIJc+qDPBGwk852JE6ZgnNLr/L8YbZVU1Z4oUfu/J6
DYpNNsuGXZdhi1H5UHd90yCIURQfVmjzwTUo7G1Vhmu5v7will9tuZ/3cPNW6+UR
ASpITy24EjKYQ8LJ+DNLPoHA98AM533QY8CADvfbXaFLDxtCravnKIrkdJt4VclH
p9LJDwyTAd4tPHMGG36uXB2AQ0MNGsHWRcLDMPX6DvMZVM9GzATXFtgeVZJ3O3Hq
DrC+hvn6pnksPmS31+7HJTtF0MYOOHrCmYT0TZrALgKSYICOIK1rttA5xcMK5zj7
2EKg0+N9jc20vKMRqPBj4x23N288jXUUjg47kFlG67U4iP6dCuDlEWMZMbNfugIj
qAkKteh4f8KuDnQHfsWz6V5QwoBW2XNOdBF94BiHSbCZftSHwdiRF9ENA5DdVMOj
nwIj9nCQ59Iyx0mhSIF45ZI887q4TFFD/WZsdp4S3PutG+oC26VxFHxvdwGXI7eE
qEwy3GKQJIGMUobEDE9owgbSgV2FdqVJYgd13Isnas2FS9C+NkqxS/mHvnnS6myc
z8uEdrkIHTOFhreAUonPpGLw0dfaj4gsrFTpFsfnD0qZO1jju4DJbFeQz3umEbcp
Nko0owuRLyBva9sExUlA/hqf9fHevIIui3sKLATk+OPZIRksx49JG5JSscpm9CBN
mdZijAzh8JUTLh7ZeLHYYN/Ao03KZDO9Hs3IyUORemWrlaAkwLLPsdU59t52gZfE
x8pymaANAiH5M9PDVwiYyvRUgtyIAOKIAuwxUKolMSc8a6KPL7JqesM1LNX5WyY6
az5uQYh+cQSsA88OujFkgTM/zodCBOiYfq3mLVgAstJUW0yiPG9cP/GLB6E+3Iy4
gdTXiHVSvQ4vHB0dRKGRiogU2dhrTJAPfzj/Pil8MVaPVrkSOe5EkRrb0a/08YcW
6YSmHpFfvnHRZIdb9rnlxX7hzzkEd7YUkUkT4NdRFDECELPwXEcY2wLnFBj077vC
YsDJZqDjFVtv86kck6SA6w7b0psSMNG3EhPfvWCPiR/5214/GvVf9kYiw7Vamhla
eKLtrrwShvIN8DCmOl2KaQaLmd11bQ1co3FGBxH6Z+LAPFhT3PIr617n8XIXauyz
M/azZUcJMdntmolFF/Vv8fBA93TSYg8SMEBHZKqyVzeZE5kSeewwGCI21IoUGV/4
A2dAIrqDVY/hwPigYz9Yk25P/omzM78ZWHh+r6uveHcPZlFm/kgCKLRRhqrJ5no8
chIi/cA5PYMIRqvX+aKz5kNj8YUIXo9FzHGH1PkglEqEaSBDh2EBCbhnYETWsuIv
lM1ueAWzHow49ARq+a4KNWk3s8KgWkExLl1OIZFJk3zrIZyJuqXr1SNyp6EK1w1e
3Cg/HUbuLCN9MPb2en5uKRdnpisyAwzBA0dh6jCRoyf8ruB5NltTCuW5MCKq6QaB
MAo+4+Z84cxwsPhw4NXgtf2NNuAsxwdfJY5S90r61rb35wFaZgIkz+sfwPUXRwMX
NsSQGVW4E4lXS9Jp+ZUbaJSQj9pSTzvL+PBdKsPp+T+xcI2TPiTOzNheSHGHkVCM
7OIuRxRwjB2kjHMP8Vl6nKohU1wS2DoTzA2g6IFC7TtaA+qhLdlfIWcfKtw+v/qN
JH24AVa9yiW9126pyWpQyIa5OuCnNtCg243Azsd7sHq87d+bSlsHTv/orUgNoBTS
SLl1RgejwFAEnOhvrCt/JN9NdMcKfxBEm8dMa3DdNwycBnySpMxnO5gRWNjc0SaY
XaEJfWxfrdfcYIAn0DPKZZhMlBN2QmZuhXpG9bdcPyMwDkNx6zgd/k3Lg1VQWZ49
0DZrcfAfJQTk9ni6aYE+SJJ/QH055ZPkfhoWrE1nFJEGTWAbS53OB8IqLhcrWIu0
3+oUcU1+HXxWglluiLGLFS6Ynrc2YTUskkky2jG6RJGvSrLBoofoz0ylwYdR2WY/
HKwupszzj5MtvEb4xKpsvEQngJkhVKhxxTOSP6zpOkkRKClNqqJDtgg/Wnj93T5S
lNJqNGEXboyDUJgxI5Rx4w7NJ67zh8abls1KkORQb6hHrWFbuFd4KpfU6CA5/FoI
MAzo6qp0xUni5IEjZGa/XhQBKNmWX5BiIwkoZRIlwnjtQK5HhihMvZ6N+N1qeqvZ
ulBLsiFJyhWdFNM5YD+COkLS/mrsCN5Pw8Nz3TwSJ580ndZGy1q4DEa25Af4j310
kFPd2DrCTeDADdtsfzfafM8KgIQSr2SKsXr1s2mMBiS1pPlDQ3QloYDnEPkYiUXr
HTWk7tUR+bPF4xqUj+XlZIdV9/ZgFKz6JEgxCyyGNj8Cj+ZC3A+O3IM93/Ya0FPj
9Cjke4SRv2VNqW9CeFfjUKRGw5A0iwUCVmDG/aKhw1U23AZHHMA7FLXvjHhyOIi/
L/5IklwojelZOzXWtEzKx9/esEzSDSFFUTC9zKEwruVf0kcfHy3mEYmP4Y/tz8ED
mEiG0AALH5A7X+hEWcujIAxSJkHHPIxxl6IRwBd+YlhuOT2AH6vY7uvWdBf/DLCf
41fPW9QjzyVlUJHsOSbJV9NBYeiFDniLwtwbN3BKDvfgGnTW+bhW4ifkkNja0vim
sOwfvIzUxfPeb9P6K5bbDA4rXZHJPATnHiKxqPRZM7fULSpLIARvp3bsoyMY1DAF
8nlDs9PX4poRUxZdnM0cALiApzAPPpCJeTsUQaPRRKdVjN3AFa3uc7mFp1uZGSe1
XEUI0lfFMlcZnZFwpxoHpQqkoV4AjZaeFezzMg9Qeuh1iHEog4Zskp/bmR5Sqy9I
TTMZNoUmL/OXWqrC97oamITuPyX23INkspshMu3mM/uDn3hLStbLEHd8MMLLSTZq
YFJoBBWUBsE/0eubKvO8XTO/HnFgm8Y4diL7QgYLGL6s0/h0J8RsYINENDN417M/
4HKMXuCnRTVzB3BAH9nF/FwpTODQStq0lKi3Ey7p+k04dI/Q8KzLLH6ML9KQ0vsO
bVZ2ddD1JFI4nxXNehhF4Ix7o5H+xs6jivfE7N1Ax1hKAnP/xWqQUEjqpByli9p/
+dpNgiM556WksL4jXuRIve8uqFwtkq5slUcxgW605lNPb8L4X1QZi4yStSFctLoB
/+M5Me+RUZdwOkt9/HzV43ql9fzR7oQowb4ZLQuN8pN03090Gr2Wwz0jUbR7+g+T
luQBSXDIdmDCV0aINV0WIWeJkQP7O7FTiAHBCx2aCCQsc1t37SCY54d77ow5ejMi
Zfk7yoCgVUy9aXeVlQtMeba8RFvj39gigw07KLGJ4GINuc6WXsy1qYPBJp4WN8yQ
TmggM8V07yRHu2uhhMGPNaQ2UXFmfCLrBkH+Wfr/A9mJFjCThPfbGCtS3UxMJd3m
NQSUTereHM8VKzsvKICTVg/n2+DPa4c+0vgX3adN6RMJPbVdFSn1nuX52B2jb5DV
FwRsjpMpY2BlC7zCVUHwr/dKDO1AvYlYzJLOszLqeaaVEfRdV8YZcVSzG7+I6qul
2lW1jGnr410hzumHcEMW+DeHS6/UJJx/5TTslIHr4Ca+B89/y5e9rU1qzxhkJ6BH
T4zsNIeWrMPwZIE/c01JmnjDr/Se2JVC2lwyrZuJmUeWKgT1AH+DAYUXdM0g7qO9
F+GD+iG0i2wbMKZLtpfd6//FCZ38B1p4afLNofw0YQ514BE/i45CqZvvsRD0BQIx
hG3vS7lzFm5zad3UFe+GbOPUED5BzwJV7cYxt+s5zMIzRBUBfu92yHdITwJQAxRY
RnABrchM+JBdsVgthn86Vj/nQiSixXQuhTuzUAOYQAKtrRRVEhaTUOPvDz4Zlcm3
0V0prq27iWnJ2MX/c5C2D6IQc37VncLXpqCCeDL1Y7nJqbFBpC31Uy9dlsgP4EaD
smTpOMQO+EU1ZHFrHCv22Q4I4n/2psWlYJKs65eltYIfP/igZV/whC/u+ZGaew3w
LEzv7v/sqm2j1eFyVgmZ2I1Rapp7Bfa5SfnWnlBGxH3VnTHrSZV+G5JNkxKpzE9/
/ITgS58TVG1DbtMYtVwX7gk0Gy+zSMgz0e8dZEF4/qqU3+clu9jo7W1GajPDOhpl
zpRnsmaCeWXgw4rMYU87hxuEBfa5IqgJYu/F1sf4Bye77MX2pphH2ziMVUlCcPAg
TOeqsZocbuLhLKgOXfw0OSEJtx7U2YbHpAN75qAjywYNEal2V9Z5kEeMp66IBADn
zsKKuhaPM2oeTeD+H2Z7yIqpZVy8w/SoHnVH81icesgeMKEFTPzcaHz/17AoD9Jv
78HMiN5Ljl/s/joXUtztuH0CE4gNnoFPjadU95zfgKSCzuUJbmtkEwPMzgQ4Vat3
V2Xw85SRDOm2A/euMM7+a9dgHaqCn3b9wOzxgHXDA72hoyNyVNDR2JEnc+pKMCZB
5vOZkufCakW6uoiwuW39vzJ+h91TUtVvLVGf0Ot5ktic2ZzdeRPLf1ewaZRnM7Yk
rrLiN5hUfijq1VVywLf4bhvTprZQKU8/2hfWaGDGUY0/uvt1uDybJew6g8EaS5b5
81hs5K7AG78t0nSl9X+YTinNa/x710nusY+4KlFuMHllVjq9vtU5eY800jGscuzt
V6JoHmC+V1tilCElJ8Fq3ZGOxwiaAZslNv+wqNJ+yc67YAM3KSKiLKlQ5WiP+8VS
HrYQTYhXKfwcJcQeOunEaA9LHBRNDyR+eK2w1GKUUF3klEQAvgGK0Yl9XVoEnQKm
4J+2VKvVb7d2BpN+6jJmxABjKnv6m5UJ+fou8HOZ+N7mLgTd9eP5yMWFxyWvwJmE
KZGNfMMRYn/jgMO6aCcFsuVO9shmEqLrvKGf5RkgNMnUCpioHuhbYNLMVFfUROjO
jhaTdxfRQ2M/5f3DjGB2pZx0rGZam+EZ5kL2jZ30Wro+Ckz03fbtn7VBgoQ4om4x
6amH1h/AqbboaqzsbZBg0SincSa99K9V0SIka8DGgcmk/7cIz/Cn0oPEOjaWI7/X
dSdA+tdhzHGX86kQDnzpRSx4ATF5M3zpFrQmc7o1Gp2KK74EIlDpEjuVksYiiATn
LnQW2QR2t6Z8wI1CK2BVLIO+/9P269CqFuKeyAuJ0N9YOhAvbKWM5rssrcQApLUm
ugQQwc4NkDF5sjE56YWgPcCEUGo/acLncNufpg/I9WZBfvLU4w4yR34291NgIzTQ
HdpGsgRzFH776zwtzDr3eS+rprCepZliJSgRA5ybbpOLS7HY5ZV9SYVx4G1ywH7g
F4ECBMmJqVhaIjcwv2DHGVHR5zrFFN5ZBx1QRTM3okXpQxHeRFLwq0Xg064aOhFH
OiuHsiX+uGoID+oXVDrIoZc2FDoG08hJK0D8kOWX/puZqIYQevjt5JfMYQd59ife
AbsM2OlNOQPdnjjiagPMZchxYWW6bcpOEgPeAU5iPslEXFULbx0NSliOMiv5mAg3
Cgaqsq9mTmPRYWFf1PCHTXyFeOETa+Spmdp76P4Tp7t/e8lw/uZQTmqG1DGzaBTv
v0I++jWWnGalLHqk7YnKxktsuQ07b5acBe/NFzc6FBt+lpZnRrS0BOWyOiqWker5
t0N9dzSE/uk364nC8uzBgavc2p0uoQ57V0JBH6rvh5X0b8HdJlx5ZkV4WcDkCt1I
J8i96hOfMfta280Lf1d71SXG+gYH8iLGnoh6plMtINSuaXzQmOuMVG+dPL0EWVVe
oEpKPQc3pZEjSfCEqPHLNqbZPz1ZeIkp7FPXsilQcow1/X8z9MxCOUfom7KVMD+C
wIcJ9xtdjYmPVrJBroxEck1GRSHsoeI00FrFIXSw5rCcMgB0Zn9Xot67by5SNcFA
Fx2nABzhHwpSfS/AZIXi+xLZu8mlbMta6ZcgkUc7HyRL+9sH9d80uFVv1VNNRGP3
naJtqGTX+wXao3o1Eeh4PmSLUzzjugzVSqdazwbZdCXmoGHjdvJrrN9ZQQOt/il8
UVVJl+jl2CeXyN66xJsX30cPVjUlRHMUYg0H4CcjUkjOD1moVbOV9WDzlcE5Jkl6
BiaHjdRvcSDkOAtU1cGHOn66dP4lGSTMRTjGuNIm/EWMJREp1uMCac/i8gpCktRy
r98mD2s1t/dClNXdD7Ux+xB8omNsVzeGHojmuApSbUKO3ELH7ttXvTGOxXULqIWm
wmmDPhEg5zfn+BSWv3/vUZ0ZR5FZ6i943Zc9AWqc6WCOlvVKaf4pC6m2skSo2t0u
CyMS4VMBrIZrgo+HGS046h8UMPJDRbu+0G5U5XQ9nu2YL5gVB1yymVIuD7+TiHDI
p0pl2Kwkf71e5yspRlrx7j+cBs2/FglQjP8hIPKPjaNZY148He3G0u8y6OIbKa+Y
q0NPHdXLMxykQQLH82Naw0WCBsBdjjQ+1jNBbkLThf4ecdEIDUAvOQpGOBP7Pcvu
goq2wQEXLI/7Noj9UJaTmpPR4o/cBbLZDPMm19ahrrslotXFDhQNSgnPJp2yq/ic
onN3L0efDTv8+PodBRxN46YJB93J0p7kVa+Em2aFY0vAFP7kZZ6s0HArckCZgYnC
2NqUuAb9I3t6bwDVInUS2UG3w4PrlQhkk5qabb9KUHveWScVfvlLO9ogvCtgqmI2
suFZYtKyfetJl4pbT9lV3n7OMVzbCO+8LRvCS8DDaj2sOa+uO1JUpVNBmCRLM3uA
BdBPicNAivkgBFpxwXEAdDqof9p6fhMOyhQKFpNNgQ/CdXQ8//yi6BuPPRK+d/ou
mI17dYeBuyhuGPB57XfmxRo0t8gUibo11FYEEedcBqx3hgUEHROGzCy9lGJO1OZT
cZ3EFw6ZFeeH0kNv9JRxMn/VFsUFf4Te8guSeqsI0tKmq4GKvkQSLv/CYlBHIxPl
mr3HT0oG18+vuRpwSL7taOfZZsu2QVTmuQtKwBNr+L1KLcv8QaIo5WtL5aHGmHCo
U5Uj55T8YJ3UXiA2JcZXyqLsJrvFSs/Cc75PjU2b1ETOp0ivxv7alNAXdPQ7KYrS
rjyI4lLxC7VfiROhqbMLwXVf3DJCEM1/MWIqUHL1ddiY0D5GXxD0Ql2fhkOURuIl
eqnQvHgCWrFH5Z8odvjB28vqpTlxmsEexoiLIzvs8v+FmD3HeE9XdXzDOep5v5b2
Cfhos5AOZP8vkFRob1ollxZJeb3OKF55+I/XI9tFoDjQi9nagu/D+8oVHdpaIU+L
5KZGK2c8YBZS9rr5avnjzwiBzv6Eo5OQvK7sNQW5tw0VfEGR/86oTJoJ5IteU/RZ
15e4Kt7h9bVJAEKY0T+BSGt2G2wKwt8PduUZYeAvSdfnK5xCQz/Q6meGe9CMc5DI
CAVCt067iL3wFkvboxxfPMXcthIzlmnFQHNeJzuQ2R8Icj+IPRfdf3VJixaFwWrm
N4XE5zvL8TKkAh/X5rRo7u+Zd3NVMr/ZKxdb1vta8bzOwQBwwRB2mnTZ5yH9a9J1
MugJ0inihCP2hfVk/KwcyCSUqFKHgNc6p5vugv8QqyyJFZqCaJeh6wb7Cwjr+NG1
m6C/igAZxEoUdT5eUOFDalLEGMRLQhjrn4ha+NhXHJc75uibMwpovbl5tZEUojza
EfUuBed6QRKrpuSpylqkT2jV3SN86hJwcUaRdEG35Glfb3uWc7xsdXRWsRBVjwvG
qo+SBMtDuQPRj0L131oKIPUSrZq96ZKtWnv0ws7RfjBEmzvFP2y40U1s+IOeGreq
AXssrN+9WrOcBSf3cx/uQ3ijPa9uTEF2YAVilcOCdcmsRUZk4VSkpFsl1euL1Q7X
dmc7dTiQn8044ijMutQ7cIp4cgmt2VChUCr3Cmo+hl1qXRFOoqr8QCLxReBX99ke
GsjbwXeV7Qd+F3y29owjbVv2Dhp+NVNMXs61BrDXj58xZ8zBqJhhhtuoQXMSZN3P
oUtaRjCKKg+Jh/q+5mk+dSXadD2xA53SDP9Yb6hFPcsleZ2vaFtXqN+hE+Eqpnd4
2bsB/2hkOc6/3QbQabdvITX7eJLX7SNNxcxdUEnTlUOOb1XQHn1ZS5O/FqjCATgx
JHFXPv3kEWTUpCQPrAkLulzRRO8rGFda+c+I5wiBd9PUj3O0zARdGh4IqT5hxirM
9A9mYIuzfhOyBc9VjJz1VWiGABvmH2ne+3FiHMndW7jzxrNaxcptpSdeLQt+stR9
+ucs3cBWnUwhieo9E2uULFocKZ5u/WYIFwuJC7J+805evS14bst0ALv7xV6UBORL
O69VfqjRaEn3x0O9IoEIUG6O6sdHVeEyHw6F5xhNxUapeklp2vL9Qtq9g1FjJW2a
GZgi9rZFWDnMxYIk/iosqjPOGmIlsXvhGAPHlJuHeRXN0nLFV3Ek3COXDH5KCYap
/4SiKaCWQ6rLnhig2q6SpxQX6s8fgnhApJiF8xJZaeLcVpqSX8MNiWihFY64PQWL
9SGaCmLtWUCXSZ0CQByNDJPhEzwJrRyrYjEc1OgBlxAProf4nilQUHd+bfzikUjN
5II3t4hqrfAlrSEkpfGzvaNn6D2lno78WkKjgvsZmu/Gj5i4a1pBldYjA/ylKaNu
RwaTrhwaRvbe0506nfyf+ZsPKrp9ya9nSr5fCky6lMAfFQ4J1UlDIiXpxvYaMP/Z
wbT53POFCRMiU8iGqejTsYRqLDtcT9/93JwAVz41b8ueRXxaK7I1aZykDByb+pkw
CLT+FsUB5MPzztAlG/5lvzR8OBj8aSeD+SfmAYnca6KlETGl41Y4DoSvCJjsgYT7
e37RMG5suDrD5phX7gYpG4BndAkHXpD7VMSqtmBK/SWz9wyKb+4zCGKnf2/7+u1d
jhpDMq5pRYTWmcGaWdZDANk1VN2vF5fDR127zbX23/Sit2Wq3NJGAC0l0A6KcemD
xfjadfAeLxNHYvnLyv6UTL6AfO5ibDY/kOZAbBa6w8IM3MVZJ+Uq2mtM92vykQtD
p3nV46V9+UDi4jpLpp8FTiCoJh7XgoXhRXWYf9Czy25I59KPygIRLSKvWI+TZcn0
NAOCB3t6geX2olhD2DcAUZoCQQcE5rcINPKBqyTeUzQ2xMZi+3Ta52Q5/SbhIprr
p5AewucrekgPWrXbC/L92YDT9fNvqFabOSmbJPDgoXHSTwCxI0ZbvDjdgJDA53Xl
BEu44E7+8YFmvMPfAPBk7efuHCh0a8ssXO03rdsYnV8dpVS93qJE0Fnr9vBJTpmt
39q6Oz+0Kyq7KNjFgzQYvzf0YfMDR6O1gpDQuSajyXXqKTwIYSw0T9HLjGEFgHpo
vIjBweFQlEtA6qab3HC6jqqEH92KuELoFD+KlbY0AzXIAGmu/dajxQHopbRf+ryA
G00/6RE19ee5qLFfoDSulL2tdvpl8a/NQDsL4W89EUKpCwlQGlYgUMw2ajHIYIL1
oc2KgH2G6Fq8oyywvrPMOwkHKpZQkQdFvfDE1IZkoF9uqadRxg2DDYgLJCB/COnA
iY2RVcV95NwTAoHlKuK1mFb4d5hAXCk2dV1FLto+ZkT983IDh6fhTXIW6oBJ2iYe
qzhYhJZVp156GhbA0l1I+h54DDJHcUmRDtlKNoev5MmkMU3cDVJ9iazQYVIBYPsJ
sEF8rV9ccphYeh7duD/vnKh9HS7xLMq4TwpIQB6JkEDFWQ0hB6prrXjSLk1xg3AB
hLRWOA/4KIHjDzcRfLJEYmurTsuvbOXrzdGAhDmbQNWDv8Ie7oFXcmNo+l4cGuUz
SYVARHX23mUG2RNsSj3RTHwpuPOjfv84lNcP3sCQfjCuVgMNC4Zvkey7aN6IkOow
5EjpXjQD3ruVs5QcuJ0sds8F7e2AZSE+Yhu/lOkjltZAezTYyVZtsJpnsOqg2KPi
EBqw6comUh59aCr0lEanE+cQIOyURmQ98JDNLqSJ4+CfXG2RSaAMzAw1fISFy7OC
L2OoATwQx9Ef/xgLvFDNOXebz9FdURJUXTv+LsNlgxsSLS0pAvz6wTFRDva+YODu
v79XZ4Z0tvMwVbMS0ef3krVxMBuPNkSjJleXaFD8eZrLVm6lW9NR8LHtInku367c
fwWn7ClUc9XnCzRyszjIoK46HqWQdIJKOEJhU75v4/VmJQCD02csZ5GrqmCinuKv
/c6VO7o9lRFbzyN6OFD4sRdJ41TPBKowMaN15he80XIDvdIP2lXNyj09ohsuR2DX
1n+aObO8rkyDx2NUNDUL3Bh6iURsgG7f3ZelYesuAdNVP3fRw1qwa0PLkD6naw2T
T977niXPKjzu5ZzL9WbRgrnMIxJCuR1EEWtsn0AFiK1ulytBIzKtAMc4/EP+kH+r
ZtLAfsuTGpOpW6Ah5g/bd7rsbz6TxFihjRJafY4DWJkGaPoYGrjFaib96NsLYBp4
yMjduyzW3Cg2VoHR7gl+cu4lk/BlXQpyryeHAO43OP7vWG6dPrhW8/Cxwn6jIyG+
fWahOdi08Sqzb29d2Zy1hTCSXr+3nBiFdzUAlT7YsD/O8u9hOA9MO6D4KfhVqiFc
7qtkXvEnZm3WXBnKbGjxsFs0HV/t1Plku3cOwsZaXfk/jmM35ypL+i12xk7GMv0K
1Z/I3CybWYj6kBwaJmJKPnGQj84Zerw02dnTrWy7hlNzorSPw54aYCTfnBcmt79b
jEln4ePXBExbpWlnyZH9dBA0U5ImSNgfBtDgMuFdhVlz76REJAYLputGxxKqPZIY
J2XwWPisu4GAVzhPu66gMchmx7dFD3xp+1xAU1NX1KkveXfbKePK+d6JxeruyUxN
+jGPMfJZWr1bje2y19lRreHLal1wZV/YqW8eAtOnUaqqPjPIVU4CMDzRExn5oMBe
iW8NV/JTQ+iNTFCyVeWfVw6KgPBEhSu8egcxmeUj/jx9sWwwDwUmlMx8LeCfvxTR
nLBhNiAmrqSwI0URXpJ8+OQxMQ8rEAYMOY93DqsWCeWuEmq9oNXk4fRGTGV6qtd1
9xJlilCuZrdg6rn6pq8GacuiU6Xh0vxN5nKCpmeJVnurKgUVSI6pOZjWK53JcDEY
ad3opsxZGM2McsszjIR4Sa4oNeugP5cJVNWrbuA02Ox0v0+l4yDehZ/mx/PUo09m
Qz01RQdxfE9T3HYNpsW4JXwhk6Qml4HOirJB5fYKNbtv/DtKtzO/R/1GvYh/hf2N
o7cEN516KIPn9KAOLXTbP0JYhTWClwpxZxST2HyecDpjn3/aF73JKFdokmjrtnt/
ufOkn1q42pCUEJEe6JQsvekECGTyWhVWSbjmOev07njGXM5Of7CtfJQ+4fJWobww
639GnRPIg8sxQ8i8xgMBm3TxsdoUHNm4cb6KvaZkELKz+nDk4MqwA1/RWqKzfGMm
FDHW7TrJE2cKUyq9eUQJvBrVEeua+wxKA1dNflz4Vk6aJ9443dAwtYMPfAFItR8Z
ruUNc2snQVbRgintQGl0MmsyEWBpkxbNs3iQnjLfT0j04o6AcOTenFQSh1ltpb4H
oE5J/fzCMbVMH2zlhc+PFw3AvqRXj8GdHT4e9dZn2Dkq7wGhATDRzVIN4vBDP5MO
vRcwjsCE09umI15WNPPgrLcu/TllGli3Jok3iADNmusjyGweVfMM41BEJXMM5UP8
6+3EwwDus/1MRoX5t+Z1xU404kTJ3Z3yi4Orp0iRepyFPZUAFVxrpgJa374qNB0V
dVHPob5PmMXsLBJsY2HF/SPpEwd927Y8IkqLN0Z7HlzKkb/fubAbLSkqex9ktPva
ojo+oBbTGENy0X+ws8of9WhPe1vFVWYvX3xCW1Jk3kcwuVsOMSGuqooLxcy2legg
5qvvjLw8oRR2bWEIl3FNPzSCZ03IhyAUPvKu99b6XGiRh78Jc4bLv95RGfIf0GmR
WXgbWsFhHfRNG0MIltpZZh3CtFnijWJJp0Q3vUbv8ZCrPShDLNPqStTcwSnr2Zz0
4IaJyc86eB0XwzwcqCqQDmtVVtgV8+6OJDB0b3pMnC1hIYm+4GiBFOuTRyLuEeF0
Y6p3niPYqIHi8cUxdWFMMWegOrbATN9e2B+vCNFFRIWvxmOnUgA9d0Uc4X7zpF0o
NuBFN5OUi6BlgMLXeUbT0BhnJLtm2x2igiNubirRosjlJPMFCkwOj5SsF6pC4ORX
tZr6lYqrWLs4dCm2WZkqU6E9V3RnysD24dPpohH1gABOzQ/fHymRMBHaBhStZT8g
wVtvPrEYUR/RntPQNs7uQZR0jeGYvUxTjQ5rgVQjJSGCzsd605GDlkPFRwpUmTUa
MAQYX0FkCx894JGJzEpCZIVJDh0M5qDDnItFsWvqzui4ZimGeaurYbR/bdKnMY1a
l3P4SfvC8FZ5UVPFGTHo29WR+Kq5mGxvCOFmBs5Xbk7oab4sN7OJwQ4dRC6mHOU1
Zfvn2eCSf49uCMgEBQTTs80pDyt80Zk7a0hzK/yGHzLc6cHdnm/wlAAD/W9V7SqS
bskKQyi69NerSCOyc5xjL9ks99fgiSpuJJlydQ61Qg+bu25TVILuZyCbGuhhYdq+
eJM1svUEFSmPqTygrn7hjkHxrRwmZmLz3JT0O8UBD7rOcHnwX+Sr4q/9PKemsOlz
d1kkbxGyU4SayNSOWRqAWrl+3dciiS00289K/44IWjXcJsWvd8TDFnHLxcnCo5hF
nNWWQmcEMEjorIkUn/VI5J6ki7qRgxZ9763BF9+KDyMw50Qxp/1IIrpKooG196dp
92gWI95FAth7EiCivsRIiWLpsjfpDqjQUPcRYsq4m0JU0o9X66LXVUiC4v+LXRcz
5S9d72aVx7/LvqGxdNOtwKcjnygPwC9N+8WfssJUSgivvKgNaWHb4JAdi1XHfSsP
uoxXUdPPsUgRnivRY1hqKsdYNK6HP1pSFSuN0nd8RmR5NbkNUxlXxfsUchnmhtB/
RaPNtTKEn5EU5n+8pUhe58of8wVJfAA9zOKUi3R5mi34csZ1oiPTRHgzHDq6gtqP
yauAxYnUZPonOvXKitfrjP3mmKB2nd+WYW78sMMV3Tmg3JJNHw2AbWYTtlC412nB
wwL368TQUQvq8WZ8RmTCevYysyfFgkZKAf+D5Svq2OnmTkGTZZs/ME0Tr3AhFJX1
k+/Lt3CNy+RB553GzafPoUsXM9CatdyytCdghRxe1zHRn34pbyb4f9UkhPqLaUqO
Eyxk7jbB/ofNci/7LQb/P7o6F8sr6GkUjwEdGvIymBpx+44KYu24gC5+KeTPif1j
vgZMM8XJPW1AVsPCiBSZWLz2sk46G5okI49rv8wIVKTMLsSrvZHLtDtkV2U1JJd6
TlcgVfPtQTF5pIJ7Nk/3EJHsSBJP7m4mXYE4EGVxAWgxbkFwiSUUNoXdF0DOZCXx
okyI6fm2YKMraMjLLwggO86gkUbMKWSI4Fmins3JVpk6l/YTCVicHQEr7DSWq6WI
cxP+Eq+BIrz7xpySnZXu2pCzo1wKEyJEI12vCRDYaPm0PVtU4XCI0wilRxZYOlOe
nfoyI8NJO4LVRM+etfj1ig4gziyqXyczp6KRngQsUVhEeZOq0/E/fltoP8yTnC9p
G0NNiMiaiKl5HJIdBUnPZOv4QuKK1ECdP8r5sXczf7H0TpDxga6C3nL+e0BbGgUk
zVa7yQ7oJA3MjA3QORzriZxcuCF3wzxZ+GcGbrAHP0C83z2uU4VjMLcfQefqjIgE
NWWHEkaxPJR5a8SdzobLzu9S4+cbl5xrDSekJFSSt2M/Y6HKedbLVrub2gi7e27m
qV/pu+3X0tO/e7tHY4x9LYw1PhRwYF145C0DASORMUnwpqdEtyqo4KXhI2TDkvpB
HbkeNPz5bogX2u53qBl8WqjompAgy1WuZzt8JLRS+Y+QxwdiJJ3WIQD2h1Ub5LZR
TfmoHOn4XUFPw6/N/I0UPu+jcsNNci261LwJfWfj7n5WYu9Q30I6wQfE7dC2lA2a
jVEGVt7LFyJ5mC/66pWABHlxV3NotXe4MJTD6kNaLX0yVXd818/Db70wBS2IvduP
FFoJY5K9IGuyE2r2mpCgAhrVlU0zVx/AMB6luF43cIfn9RRlVo6nKOrNgAJpwKnI
uxPkRO3rCxhu2XCTNq7f/bLX7SjNByyq+PjeVMPp4OKNb/KxtG5/rNFc9cAy4TY1
TIuG16s37kudJtWstil/fY98OhkmhdhVKTjXgnyTqKe3anSTcar9g8wYC5cO0PBa
gULLsh06heGffp9De6DZ21iVh6CzTmfkfOvFEmO9jFqqF95pOIvW8w1c/L361Cdy
M6o0vZqPej7GZpPIZgeiW9beW/1tNMRKQwuKb/2PIK61lovWKjEf7qoq9eEJk7YK
uT7GB1NSX3Ie8pDiIAOgl1KZ+LuKxmTS99xPoyZtc67Tssjazr6s9m1roJ8Y3WkR
kXUPxZSpyKCcWcmqvInB/ZvkUEjlxzB/Fq8boR067sMky4epyUfTciiL2u2reqd8
aK6cLOWL+ze+j2xE8ZUAV8PNHtYsSvfE0NT0PzBLlVL0MPS7+CPY1cUhTofrMKjd
VP/xvSbjNe5UT9V69WpPv8XXDA6F2lRLgFIAcnVGwgU3Zu8NJoyAQsAmKLdmM3qj
dNfc+2cRR2cEbEX15vamVjgHeGFicBOfQ8eR9hurn2m/gQxo29VfYF8BQDbbVvbH
k8wixVgx9MeIn9k1CLopzTWYWqNum48gGigJJypx1Cd2FZygzKch62kyfVwiiLpa
`protect END_PROTECTED
