`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1XqMQ5GWPli5SS9UjWw8SvXOzgthkPyAeZ/n957sf6GB2lLQuyUAsJ6+XNqhEZ0b
/yBKmlQbRjYb5XknLDW9AzLM5oU7VUNSPhzrbLZoA1sPSFUvs2i22nggVAklhbCP
eADv15saeyC5AQEiMk7ewFgbJAl+OLde1xQDtXPHGwCT4QkwTFauu65RYjpwC5oO
X1P4+CkG2W4xzHyXpeXLfqnUAmZ5y05vWQ9QdL+F7CC9yR/qFivn9m94GR+xfwSY
IB7CevZgl+eo2l1lN7daaaNSSJqRAFgofifTls/LW2vNXWoT4J3Lb7IZ4u4sYnHx
Ow96ywURiR2Jp+hzJBndY+4h3nYCy0HgLGivXl2JtR1oCNoJPa2XzhCxSbGfL8a0
l5fS6bNBn0+ufIFK7Bftk6R8NrZvSMqI0ttdI5sQF7FRxyP1nyXb/QM9lOAm/J7+
q8QGqJotqI+suSAFhpKaobreqFs9Qmy1Li8t04Ewu22WbF/gTGkOCv1Q5d8HdCn5
OhSbgTf4WOxdgXr4fG+pYlmf4+xRTz1RUSe5PqkOXowIOhLoak1UzIeklwCrQ21C
DODKhJ+ns752Oa3qD9FjSkZ2MdaiA6rg5zkLJV/ovDMrS9de+R0pLEygKW5L6sD8
dCBimzjni/n7YZLG7eeW1g==
`protect END_PROTECTED
