`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IaRApFH9tLDTWxwWSw/2G5wxFa6/w/NJ7knjvAMcwK8CfIHVYT5DGYu9tqVWN9ow
PjPXVj/Dj3cAjjZiPpI1Tl0ZCCX3DVJQQqD8EXnMF3hOygutvgLd8UoflAxOT2NW
ktVEeynRTW9L6Us6HeQ0DRajc63Q8p+ueRhXpOMdu/LpS08BCM452AsuTtkA7XNv
AR5P1gaL8sdP5c7m106A+ENO/ZHTpJCE79T2ha0cVgeXTOYhMxhHGrWp0mswhQ7q
o0tG7PbdyDexLOtxzBzntSX6Yzr43Mwv01xTYAsh67yR9ngAuVNMMLgrbGJYWSXD
rEE1yymMGFQ24R/R7NNN1JGJ6vXL82zCcFHskm84ninoxYQd92wVk2kERBM23y5E
6A0da1O5ZrNEoButeUn3EsLesDqttAYNQQVIWn7XmA0Mla6HMLS2UaZz7Bi7I99X
hb073IUR79OZqHRdZ8rQIpyAawBhu49MR1gleRPe3XfORJ4Hk4Ef8Q3GyJLfuHuA
RpHXRXJQLN5nZMRYkjOE8JaKc3kMTpXoVt2U9OYtsWWpr27K3WNADV7tdBhFPbln
EVVsL8fpa44rgTdtwnLjZ/zDWd3EsA53BwWdR25RvJRKRVsyl9cs2g45C8c4Llgd
hgNBz9BYSAbtH6YKsHfRXORuqC1c5+bvEOqfpYEU8rYCiqnDLVijBlqwH/s2tFwh
KxSnLlbzBpQoRlonuMXJd4YNuO5ToLx2Yp+CzunL5Xw0BlmqgxCWXRQbVKa+PUtb
OJraX8f8dOrtV9wipfeIdtwFZWHXzBwN7ohqZO3989iPnRU8oGTGNOYy21MvsDtu
TiYB2dQb5Ddm+Bn7r3Hg4yUHg9ktXatLFVRqyHrpwWf7O9L7qNflRz8IEDDe5JwD
F42GetTC4Vuc+c+5awO9sERKXZHQnzWRAiugjJH4DyOrN4PUO4xPg0GJDfxL8lzc
15EOAn3idj1Aiz+lKlVGagiOhUf4LGRZqrBtTNMuHFCxC/yHn+vPUnxXfjMlS9oZ
rUTX5b7ELsId859mFFNbs2ukDdcSJR5RIhO+0bb9ofJSC3qAzVZPf8VLo1rUzXM1
gwMcmPZT5YxoV+LaqjaX1RL36BCTLIEL5xQB3DbpAMUGZgre+dfwAn5zcxJoO95l
/0bvc4NyYX8r7Cr7byH/Agz1fwU4dwYXzeM1LbGbGXr0hEC3ySO35Wvp2AWga1yL
o2l1bLFENs0xpzI7mnR/tYcu0GTGgn5PaWHcUTGYFztffK822TDkJpFt7Nvbwbpk
9H5OX90XvyKCI97LjZuBScrAffnn1YNzodAHHi1N0KN4BZ8BgwIb/Q+kTUHj8BrX
h6QxxIGYkADcuXrcRDetww==
`protect END_PROTECTED
