`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YNtAMdLhR2YY+rpGbjhjifHs17CkfOJAK7lil+mD3AYMkg+8gDwq3AE2Q8A0nO2a
a214+sCc93BOqsJ+d12nwI6BdpDGOfaP/clzA188qg3wums8KqXSjIXixmsZsdql
Nqs0mDnDheweoA72PZ4zYTmw60kqtOb8KsvTaHX/kKYZ3U0wuluEJEdvN48MfvyM
Zbsr0+L6RYxnvpqyit3AWk4zHbsmnUm2lbIheEyf/HJjQ10xaVjeSu25N/en4WD6
nGMkpGJnBWUNL++gFfIakhhE7xmveK/Km6RB3xRjZvRRvhF5IFhVbkIIr77JYeEK
qs42Pde9tVol9CR9TEmpoWiOYjiBwIzrngUuvp3Fgzt4li3NjdlJ9JL/1H5gLZqo
Y3A2bkAKmUQ/lnHYqzBGPOF/caJpNBD6aNx8Pkd4IM8=
`protect END_PROTECTED
