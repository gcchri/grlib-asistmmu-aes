`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OS1qzClNokcvkAE/YY+08RF35wq6Y2N/hgI/Iwfh7UsNNm0na/NB3A8mNgLed8PW
4f/umRV45w7qfbpd/rZJKH23hZhTbtiLADfbaop0ut6FOBU0zNzNamAht9smwVYb
tanNqtFFbwKc8frepbZOH/0lYJB4R/rduV+oWzaTmq7VqFckwIIp7qcgMsRxaHVT
Ujnu+XyDw2v1XmPLLVEq2BbQw2H4ZYXacT6p9eLSYjKXYhyoz2DZU23XNnFQX+4c
dzD7oNSPyvZao35PuUGmsQzcM9OklnHAdhWtxCAnIHB35hgUZE8DYF1gn0AOPhsI
l1bcTCkUwIU0aoxOpGfUq4qLmCxk5rvx8dvN17Xo7MiOiDqB6rSZsCtlM53XZncK
HoGYkjbdVN508SGLZnTxMCfn1NQgtJE3/HkBhX73k+OI1ImGhGDFWb5a7dBBMY7l
KEC64bn6aSz8W1YrZV6viDxHdXO8ik6YfZhCBZd5tbyve7/Ma9Q67o1FwueJNd3e
Um0saDUKOKoCGlhluzN5SBfn9tZJMfhhWvnwT516/+k4IXEUnOqQWVe8ns5JPfm+
n4kbjf8GcPqHBopOZ/WXTchTxJFhc9EwtxfYzH10vtGkhSIbyVad8yBnGVruk08t
N0PNtAExFGJVYtxryNnT1j0jgqvHNySdg0lgekOjzcegFwY9jBslmii2375JuCs/
rRgOiLGKBX4cvaHS/KO2s2dTNticev+ftywrXxaslizpAMZ3Vq1zqbBZi0wRDGr9
nUOaTd4eUTFkKHRGRLMolemDO6u/skCUABjQWI0n8y6k9lSskwCVXcfiIZX7AjAX
uJRW5dipgA/X/hqwnn3FAEOXKbsAlcyB6RL5oXYZc8mkBvL2xPJ0MoVdbEXxmj/w
IsMbtNBDCiYJxXmBNV4X0Mz/qZOGtlJ/77HVVIM03hUl7hbOYV2Li602Z/flTNvx
zQOsP6lawIhd0/PlvnhhMByE07bClUI8oEXWxCOuLViZu/CD42e0xepxIKcGBXG8
dKswiIsHWW60r5jOYUiFaGUv5H0Ap3P9A7Kdi8SYalE=
`protect END_PROTECTED
