`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d5WAb3vdoU9eI4e0ETHUo3iMqy0v3WvxkqnPmkPmPtfXsctlw12W4WcgZAQNUisb
jFcvZTY+o2VMXzh5BkSY1m6L2fjrYWPtzyq9pZZMhMayz69GG/UxllPqNNMHYLbO
K97sBoWu71YZ519V+zJ7I+B5PWJbHNbAiLhngKdzJMLtyJuLY9x+oKKU6o8vyYsX
T/gcRY/yfItDeo4d4QXncmrfNomSuZ4wbY4ho0WqPN9sDrZ4LUIZeMFeYHZDpaoX
kLdTMYs5ppyPTC9qR6JfUg==
`protect END_PROTECTED
