`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k6luMxLmg+kA9CcqfHMEDjNNxfPii3Sf8g8vALz4fUOQ23ZieX6/u90OKpH8XivH
8WwElqcFSt0VyQs35T6IAfvcc+FQwtkNW+wkEKKa9B4IsrONoZLH7Hggd3HjvQcd
q1At2UaUhCkcw1XAocuX7DiX4BMFUmjPsr3no9BPr2O7Gv7bjrvsMH9NcMEAuuWj
YmbO/fkgDpN064j3FJ+opAL42/BMMwbh4YeGXF8o0B1Xzw48d9sopUJxP7LGyp5s
bFPO7XK6tC1PTbqmRufy4g==
`protect END_PROTECTED
