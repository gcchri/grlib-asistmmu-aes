`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Q3ETePNN8SPcqE02y/XNm9UilLR1Uly06l38KfRIHb5KUNcapa/A16MxnS7DzPx
ybxi0ywCFqMg1QDSSUlerLjlykPBCjrUIGBLym1rc8eX2hV/mhGM2RkucPFEho75
u8ecJQFCJHIBLHvfP1oAXX1OvwrQmeOHhKBLNBjbvRIKrMI98EM8omb+rgDHtDgN
Rgv43UlNxlh60PSw3ocMo31Zo90FRMKYOwUpEYTmcdjiKic/QThwsF0+TdAzmEb/
BGoX8d33m9gE4qZvn9Af16udm5TO7Say5gUo//TjSaD4SmIA2qcdgT5n4Pi1Hn8e
xVst9QEzh9LFR+Vf0uF+frbojO9ULcu5UnBIZxMVHbt/N0y3UQ3ghUhV1pDK2cKE
l2Wo49a9IiaWRIJA6GgKjZhFpOMgBVnldUf/WqpDIeHJzqVODji4pXxXbBJ+Xcph
Ao5hS6HP2wDXc6tP6lBLLa+ln00nYuV9XkHYEW3HhRYkjpdNkpaxT5HqphtVxLtW
emSeGxIeVBQ93IzOBuPz6VHckPxeTgQ62oIdyxtPOZW+YIVmJ1rp7pwBvJzMEgpn
692WpvOQfSJFDJGOkUsfwPNVymGf/CfcOrDcJhXImaDvVrwrLxh58dUqCm7XGKIO
CGWHaQePHbsPCWVST0a2vCmdLuPx2fJjJX5ciTjtbFTN9BE6ftGlhFI1VGhJEZgx
d42xs5tMksLJ2AMa5yb0yWd3CwvqmV4v2xaUAw6dT3ABVpRNh29Ij+0OHFf5Q58Z
vVL6VudQYYzHMeWHgO3h92/iIZiBR0M3J5j9oNJ+6DKyafPo/iV5S1w2Q/DcjnRf
zy7wD7MsRFh4y2Pke+OsKWZ6+/QFyNpjOaXjBRylq5pt0tI8gkaahLG8Hc6M4Oxx
c8XL1iNSMDs85tdn6nLpS7c5d8Qot2B7z+RK5CocpqUpuw96PrkeV5TXZXPtVfCx
IrQ4QruLrrR+rzABlQqBng==
`protect END_PROTECTED
