`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SewNUAFiH0SbAEJOnJNCQMrvl7gr7vv3kVZiN3sTfRiS3SpqxgXXSXSEqY6W30/d
K254mpr0AwPFOv2pkYNBOdQxTm+gZitmjGc+Yv6+Z4Ov0qrGFkbzhKcqPytCFbVG
X+bSy7jeD0i5QzUdNJsSYHeCZ5rxHYzKSDqpIoVWT5ofDbvuxCm61v2/oOjuVS0w
DwFhsrWkltE0bDiABB9RYPRYQwEEbOkVChUHm45iGhvJOtc+LEsikf6nq3bP+hSJ
fQbz4ZKF63yNVGJgVHwlnaQevStFOb8rEa0q26/9SfdHCMHmp/2MM7FE8s1pY5qO
97PkGz3WtsvhJg/9Y3IVu37z43XrCd4yr7kHIVtTCz7OvbbPvmVe8eATIcMdQjwF
JSqrksmtLQ6sBmBSiHKajQez61MryXTRvo67wP9LHyGdODdRJKwboVMHj8/Kxn8u
aFT22I6+cZiF/Vn8yRBzG2WG1+4HgZnRCFcMvwEtwmbc2HJ1udYaomG3m+u3yjKS
`protect END_PROTECTED
