`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtRfnGhgTaa7iBEaQbShk2eV65XNlB/UPTanSrXfDJqaHw9+fGCdYWrkmHbelEaS
kxgfhakFiYy/FFHHbjZeecH7WdMD1H+UMLn/UHhPOpPBDqXjG47/slXaJSzadkQO
yqYccAYqEMnepI4VRVXXnGmclvyugj9gISo27q8X+bk49RiGK4QL4Y1mbjacbBgB
1ygfJwTew00SLa9lo83sh/s54gXGwFEJP0uxJQ6g6Q4RnlB7K8T9Uy0K2eqLa4O4
l5HV5G3X2tZZ8/tEHiWPClUmMT1ph6dbTRra1MQQEuq6fPNqJKVUTHECDweuHEl7
BMMaRGjB9EqPNGQUL3V1F6ikGG1QBtegkJejIVxEcfy/QkbenBZCryTES2uR3Jn+
`protect END_PROTECTED
