`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aOViR/AVx2lAAGcN+Ew7ucoKwfGNVc5kGP0z1EM8CJeUNCK5O9uKsdp2nc0cfwHd
cuHlObJ2jvDVy9agH5w/Dvgqy6NYwSrvB/Tw135KgmFHFdVbXVUjyZBo+++X5ell
E+cVyTpCBDGb4PK1oVuL6DErpKKZDWfGB1Bs6kBUYrdH7SreA6Lt0ja/4ZfdFi7j
omwgx8Z5R26vnhiBV1KmXgB24/50RJqxKgWGvAtKYtsh9IEbF6RAdpPbiMuEOrGm
RmxmQM5ThlMltkUJvGNjrLXCxAEHLII/BzCVkB0EGmJjb8qe2epsDqhqhfjLTIct
BSDa7Uh9GlCpnkZYFGoEAxhrnlVZCzRpE0J1QzyQ2e9dzCG+1T4DxK45r6BFXNQZ
WORqlktLpqpHPDwTPdhshscd6z3sfnZZTAi61N0Bn7U9EBwfS7hzQsxeAcu+N5RG
qd6MUxYXGrOCgWXuL6Ce+YwJOCy3ClZD6ns/rvYEez8GkmxCkx21Xq6HC3+bsdGE
jQbWLNkbFZcwCugaTYpXL32IUvFoTcUncgLIv/48QeTsdTcv4RyU1W8EcvPzICwm
ZLjA/NyearkWdI3Ps0V4nMk2XX9owlwkB62Pkxocwmlr/V7GAVmaHI1pz0Hbzdqz
UaIUVZuH/Fx90J44FDQaIq7kIHjcAyF7ZLCYe0tT84xM6k2Ict2rOksNJ+HLfc3G
ZhELwJxrYg7cofvwpaDs7I3uavIGpBQmFE7BIjYhDukYnIcvXrDD9ml7Pf9WBONc
VWE/DwQPQMOHLU/w61uH4g==
`protect END_PROTECTED
