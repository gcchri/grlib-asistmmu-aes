`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tLPYOaBiOgGIRMJOG5JnrCQbnWhjtfvmb3eVu4CvTV8VZ5Yn+Zhp740C+3NyfnVr
/7WCzj0BdQd6Dig1QXTL0cIIPYNhGfqz6ud6jQbJq3uHtHwQ5IkEM+chJoarNfg1
dA4EQkG6lAfqiteakcZG4mn7bKCJE5NXnrAG2jIn9vODBeDhPFn98vPp6kL+EXbA
QL1pdrlOfnoDCpf7fbA6VirfnIZOM6j6RY624tQbPy/eXznXWgJBlMF2n+9ww964
APKt+YutXClDJ2ptZXwusrDulmntHUPBlZ5Pg6bD5KzSjbmhvacETJDryUp65pkL
4nbrDv1UJn2f3tR7UF+i2kQjgZHer7LywvG7TRs8UDJc5bAByicbjV7+H5DGey2H
CBALFJfE6Tq+fnW+Y9oOy60bLmow4jX3XzN1+UWtIJCxjhCYfq3q0DuK+G1V3awA
+NaqppCQifNrg967ciShIxj/QL5p4QXrJQKh9HKC+moZhtCnA2GS5+gBmG0WeQbM
wroDz0lJ6fAUKra8OmT7jMpAZevoTki4X6TcSX+XdhRo/qp9UreHC1IGgKjMbxeN
qjPCp4/L+e3YstKs0zeIlqmdtzl249E2wL2RvMTJZRrNPd4SFFSk+qe1xXwbU/lt
kSVqZDHCsg8yPwD9e4wdocxvPlXs9QHTJlA/iZMX9UwdCgLjNeE620JlSgReo08i
AY/8+NeyItKeTqSZKD+iMXKcxIQ2VTDDz1GUUTsmPo/uPhkNkvuxIKmRv5P56BE8
YR32z9dPwayq2jov86KNBVibiHz1w4QNwcMqMwXFJvLUlZzzUgpeg88dtwBFPlwA
hxgokPKh1HiusJcY0/+ML+T7bUHI7yZcgI7D+BDRzQgphpjipEw3cGHwTT5R6rN0
V72KgxKGENl4HJM6gX4CUruzb1rUWZBZ+cTT5Cpk2T4YGftenj5ZcNg86RW97hQb
/j6YAZHsDkFnYR3xW942J6sjdwSpMj29CO63BSay8Xt7BLSlI2QtZIG9ilxv8kEH
DsfT0SBYrKYRSRyZaPMCW0LFZMO7Mj5zu5CUiOiU7BK/K4nRyqAx4s2bx/SqEwwi
VKng/sTwHLrXhtwgHwFBVXXUAHwjlWK0NihgGmdLrypGiii5p4z3CebEzlPQcoHJ
nhV+cpJ6A6WdgAptMDlnWHo/uIQgpsKNaye6aKwneZtK7lZAYvb09LJVJNqw82F1
PAU02N21cGF/cKf38S9YGuQcOgkkAgcf5CwPzh8c0Ssb6viU4tetkQhaPOO0eboO
WQHLdLJ+3WOsQv543VyRXB/MUXsq3vwcQwyEFO1GA8hZGlxJdMRmCjbUulhgCtOr
FuxFeKI/bDJcJbKmZTgtLs051V0FvH4QGU5wK6f7FxAtu+euzh8DkZLIavfRfkX2
XNLJSfmy+CVUcMOofRE/gJ5QztQ6hMAv3jzkFSRwwuBPO9KjA/69hhjq6WyPOEYF
+DUXEHK5TO0mgGMDgTUlj9I7PEHAJskPXaEWBokdZRGJ/pzLCNL/GrmMrT9jcDH3
IDsYfy/oNqveTL7WRwgJsBIgZ5+v6hUZ9Rrtc91c1r/VcCVqBp/g0YP+alYhCprl
CBQU3UG5g/9Ptv+lgciX+cGXrT/kSH7bd5QmcE8HpRm89/yh+SVczLMChGr5y6l0
v5vV+GesqMe9oc8Af9cZEMRdeckXU9ALC3jvW4I/0cFXA7XlOTiS9g5eWcUHGCPD
oVoQng+1EAnYwc3UrB6ief9oXOg62KMvQxQdR8XCRYblpkbEhqfTGSXhcwP/WPiz
9jjF7+QH2pnKJIep4e3g8wYnYB6jeXyvLJK2z5MXOotL2MXN3u6TySVBbsxblVPR
sypc7Bhyv9VZZavymNgziITUKuzAHnEjrdqlmXMM+iHCsZ3+0996ZOPbl1rTPObJ
ccWEn2oYR3wtHnZQxB4m4fqeKcSV0UuAl3TPcQJM7sJK8Sj2jwhLvusqJtKURFMr
gIesxqIxHfGB9YLvfEWJTOsR+0yQFN+veyG60MsARdnUlWChVVZnrHvozvpDqiJ5
aMFmxK/5a+M7UaNMhJROu5yGObENpHeN5iHEUqqwIMxrzjbgb6eqcIQoGXWWg8cF
3KmEnto3qWvlvn5/bNvpesLt46N8nUg7D2gEB7ES1a909x9DRvMzmVbYO0EX8BRA
TM/q9F8PgO6I6R0ynWhamNZg6ISD2lCcwlZeiTIyBZxym+zzFBJ+NH2x60Ki5P+e
Whym9YL3StU1YMp47S1OF36PO2vm8LjMFfWOzC8KoG7PsYnCWe9Fdh99Z6Q4bzya
9wd7Ed5+jwRh8MCt0iIklEDcHFPbk49ME4cITiJGGWR9iha1xru7nDNi2DdGXVIT
hb1DqSEC8OivODY4WsRdgtKgt3XfDqNoRCM+aT/15RddxOu4C9FrjhzLZXbKte+F
c87Eg5XEfaW4S73fhsUtnGBah0p7ahVn8weQlWru/J6tks/uE9IwX4eZozGMeuty
UGSpxgVq390XcgKproZI6JcOUxJZ7dLU9MSZUGjU5+vcZbd2RddAqmzfnGllkXT0
XXiouO6oUlNobwYk+5KjSFS29AWn9RGcb15JMFC8s0UXr5qkRevXsy1YPOzIGKtJ
SLithItKE8GCYtcsNOl0JJjtBqRl8mKDo9NCFJidc/WEiJeTfGu1lzaIpExtNRF0
htemKIA9TGKxXm/TaOqV9cj9F0q1EopoeRLEI7whgCAc8cDqfCiLjGKTlXuWGuqI
u9zEKdUxlNWlBQuASEi3E7UhTmVNr09RnPBQ6gN24JYJC/kmu/cXQ6ywd3/qx/N9
tGC0KCDZRr8HncSR+9untb8EKRFg9au0b3430pugK2VRrGHa4M/i5M/1NFAlwZc5
i5ChO0so2iJDB8jZOe/VZ7PKqz0lYM+aQ2EDiiSr3d7uZuHH8qaUW6tAZL1LUlAA
ggwJoQLlpaV+xYFSaB4y/B2aH09Bc1GP4sbc10wm5/iUnHH5eojJnU5QvVgICcTC
ItD/gDfZg9vG90hETG/CXbQ1OY43OKEYuuk4inG2xWaRXZLa8rMWoIwsLM/tJqRD
EBguzWWyo6eAlwGWXgVCz5XeffEzKvbnqAPzgKP63T4Un3cgQFjBhka21cUD9voT
E1j2QooQ5Xi9FiIId0UnlxzS05W7zumUf3T07XLkVpMmH4NAc5s1sW1kKhggQ49f
pE+PLK/2SFUNYIavr0Twrismz2YETuW6bry1/0RHJBuTtS956WTGK/TFUvcgSZjS
Em9X5R1zrPpaevdlsFO1ktgbMCHIi+nln77aqpxGeUm+pvFx4tHfEn86KUDwBS96
9Q8H82Z6bUFpVVX4Rch12elwV5pN+9kZmSMUb0y84RE/WoOrqf7xs4y3cDM8oiyJ
2ULynIAg2uhavKqQs9iJXT+6Rbx5++KOEG3fBgy0ONilrNoY/Ouw8Yxl+3rXDi0I
lXE1IZYpAR//TIROJrsGPwP6T3IJcB153Qq8NWXBJXPdecdgJYlNzQwFrxSVQNC1
UdWmJR5zpbukQjiRMMuC7xS7YM0qU6FMYtePA1xuKtomTo3uGeiv/Ne6c3F2x5Q1
ZwqwNL6zI5IFrpg5q3VpF7IvxM+ZjydOZ1jS4yfR4gujT0ohcfiPPybDOgjTbNnv
3TrCfz09J/FY5FbKpWryvxW+qjxZc1XBP4pine5L97VAm+Y6A2tt34D4LC3zRcPN
2xJ6vEkzBVstpHsQEQ/TPODifsWu7shn/tniJF1m6XU2XWKPyBu/df4ycIZeTwKO
Ayjqk2mZDn1CQBzuVyX/Nt1fovrWUpqvogVC/cthnlniv9VitnD2sNaq0rG3RaId
XqOv9gxQOs7pMXzKdJhjuWE8hYolWiLDlQS9ZWLo9gQ8lHfAUVoDrgMwJgluoEqF
qBwBrhiA5BCuAK+Tt7NNoGIXWkCvUj5ihxDE6FYUL929lanT1hFaYJ2hy56Au4Vk
n2ToZaW67Fis09KyAn+8vbzN0BuBkPdxSmE9k8E3b3Hb3eVvz2/HOmla+eGEF8ma
qI4tTIYobYLSy3ygZxMHFysl3MdQZa138P7zVPemS7+h7a6guksf/qOf22gZm4Sn
6Mb98/vymNnV19o5VJp58k3J1xb87ztqrigfta8Ubdyd4CZrh3GLNp9GBoZmfxFL
J7PFX5eiLgGF5zjxwya7+90ZB/cErV4xvI9EmR1hPQlPsmhrkgH3BY0WPwGvCt1O
cqccJJSCtQBpK22A2WDgFp9Xp2SAa3m9M7PDmGWFTs+hiKMMjBQp6mUpDDSmhsR+
q2XwXiwYv9BLUYyClj4tfocRWbDzzu9xsiNDaqYSXtcvpXXFH2POW4tMij+AcNI3
qXjZhRkJL13hRdKxY8VsbnH4p3FkrTEtto5b6eIi9U2K+SxpzM3g6iexg+PvcJGe
7HhE2bV9Z0tVB11Dj4hIKBK686uRGY2miTU8qBt4JrjjsSv6sGy9VJJncSxvWYCP
GZJ4G0V3v/+SrGenml1lwn5b9xkuAT0dG+dtQpeehkS73hEFiiB4CUmw/MgBREXf
SYJdloX+77CKOpNJ6moE3SFAuhwo8V/4OZzK4F2Z+6bVqsT11ttv79tQnIPbZqGu
+afxGtwwfOM1+A+V4jb5e4HpdTi4T8LgwLTNB3u2aDnn5DHexfXdNnF0zZ7y74Fc
pI1MgxHAsSpYomGJ87vvYPEd24qRIgN5tAMfgddsjLa7t/5InEowvhHn/0ZTpNrx
2AtLS9WRP+MELM+bOOWZpfG4XSdkFTSd41nRjneYNF6Zb1e+JgP+tuQEpmAHbTZJ
XNOZ61wWRA19qt+d58/wmEnzqV2/o4F6bfmWwIldYq62KDq4wg4cw5pPme1KvT1O
nLacKUE+zCijJmj7Ui1V7tNelZFraBDArEPHhxd+btJwHNm8m3eXRAr844VQCV9c
nuLFec2JlN3bq46om9pmu6lWSrh0M+E6djelaOONuc9h2k2ZmEdK4376uiATIbfe
O5SH2kD/nSMVy15k0Voc1RUT9AR0/pcrvBVf9BXDEv6rEgOWvxY+lfMzz0W1ktVS
9gswuXcmRiLe+mlU46BCEZMzhzNMvBkOXJvwl1c6DvDqmy7PI/vcQFSSr5X7B1M6
cqwa7eNjc/AaViguPTECeW9ODkCbA4BRzbHQ04vAzw0/1cPIeJmFYd8krO+n4cCn
aF76ofbyCsgBzl1XodnmxqWu6oB0v77NRVqHZL9E44bOzJOSEGq4YWyzluKaBCVj
yKhIT3mlgUZOqSFVYtDK3D6CiGp0f4HHml+EkG4fGfogWR4jE7h7Rsa0CmMO2fH+
/NAmfNoHNJS2ieynbWh7MpGHYsQRRom1PBqJtK5q2Gt/3jWauuSFJumwGvV32vZC
1vVMk9MDvMXlhJUXJGChnL3t2hbZX1MyqJAj/W2Vp4cIK5HJ0TwGDBNfgczlDK8o
z5ZdeD6OHxvh0KEwJEK4TvsmklxNahVmxlTyg9w611dxPKOn4pNWzitTYW5TAkan
0Yp75EPYlcjsJoP1ZZFRhnz1Ahj70rGlbBuqD7O9NkrT5sj2J1VJKdCmgR4ydscZ
MH4f//U0gRILuuwM+B83Sq64j00rbvh5w1e9DxcPQ7lxUM0xFMSMFsbgjHgjWCaE
d20VHs+PyKwzkKM0InlX7JkfFG+DRDCjdz0ayUbXxb8sVi106U70uyTpowZjo2ob
X+30aQaf0+22gB/FNiPNxyL7//25Aoz0p1xGKnGxPL//Wc1AaEMz9ctzIiTXiKag
oFARK0uRelwiEP7TteaJuqxZhTYO2qcRYx8VolxLJkhsJtx/QMmm9zmz5L0csCp8
P27s/m5hNDqShhT7ZChTMMW0hRqB47lZN+YnVEchrtZpJLXQ3ECu8N/BmB2cZ8/S
/6qb7ZIt51d6CgF0Wm9TyKiFBLw0cwxuY/MO6OdH75/eBqkbW62bmUpfOPNxom/f
agk8E/G0cdGWF6AH2NdTsck9FL2HywT7b07b3PJSyczCqtEn+rkln/l1AvsLS0J/
GeqA8uPZqkV5JLloqjtvTEXXgZ0IKhsaUpvPLZCTB0YnN+qkcVa+yVMmYzYtRfmJ
fN+lJZ6AzsTloL9EmDshu+mLmEnLB5Jxt/saJleaOylIocqpgPSB/dNCdZAr29OP
9iro/Tz0yWPNhuw5O+0PMciq9XqtnmHXl3jB6gmgEOsJVAik2W/vz1j/8YJTPE/K
rRl+AROC8mduJGxn2O5uJNe8J3Qi+q5wYM1YA0QKRbfsGOlnIAi3wjlILKbWcFsM
TAgH07m0J0283AhNr88ektmXdZ1gLPOL/ZNv9kT4nt0qFU65w5oWgkljKsJgcsmn
4jOLH1WJJROjUGKISzFARbb/lxrggjrIO5Ouu5Psm3Llpd6WwViEtAasiMNZ90GU
wfDpe5Ig1Ro6Dk4emiwd/IHst+JTpLfeXPvWKywR6RYn6Td4gpnr27em40TQOM6p
Ujuk+vI3Zjodl2pVp6BeF5XEx45P1OZrDLsp/yqFYEMiTb2ovrfCRb16VP0CPOuu
XdSnVCVEQS0wewErMXw18w/F+LyPvujzk3A2xcRFaRg1U44NjZ6Ys3GmVwb1nLS8
2ExjNmh2M3NhMQ4FSLsaAW8EnJT/jHwJLYnTkIQR6i/mPPgesU+Uf06MyTy/vaTf
jofHYTkph7hnsuCdnFzYq0EcmQJT49k6tyhYHoe+u7YL//OOeWPNJ/bd0pes39ax
YTlbqf4fHS6D9ZjQDT5zksM11Z42WXKisnbEyHmrml3wP/htw7v5kEkJACJ8jMz1
lQazThJQBdWCx5bskeFMY8u4jtOw2hVyaBNOGK5lrPF26oZcaCq7a1bbieVxlx3t
nX9A+RNMWxccNHuySnBAyzSUIwJ/FmUYcNrWyx+F3SmE9UUMc7hPC73usOOnaUvD
KhclUJR0BRUHKY3F3q+fE04SXerokuwEXmv6m34jSAWDu+mpgQYEWKgtXY6tu2Zl
pebmWb/Nljrm7OXOXamrkTBKoTlTxiGbNKTbOPWWTIoWlfFm9GqEnD1SU22nZO3Z
oQQ5nq2rx6MqwSSlyipJ0I1jgPRHxV7Rr7v+04EDu2ucnNwsXFyEKGERZeGjdP6U
YXA7wYLn8b3LOB8ZoHHq/GToTMAaMPu29jbfpy9nDtHV3YzREHJhj+M22YA9KZ7/
qwhEw/w74T4z++q4wNoc1sDr+TwOOdWIkGhp3sSjsBfxyd1BX4jBU1NHzi7Jsoe9
2TqbVNngHWA66Jr17C6KS9gdYk1oK0OrENKMZ12xcK+cm+jPy+El5IF907KVWLqK
bgRzZcLB7xZztLIWWIAGTIU77iQMpwfckt9gvsW9Z7kVmTSCtXBLnfDNHnBNUDyM
AlMyBhYzjdKw/eqzhN8Bd2vtpv0Jx90KJ6z6vTHZdBrowqBdqtgqCqxgqpzSsCsQ
9LV0KgHC1Xl7flRh2lwHYsr3xeBmjbX2+DPBEbbbzYxtwtn37nRsH8P/gimq6em6
/cQlO9NsZT2DRIM9oZZwAxnbrCfQkCfrvv97roW621PU0YMfkZspXjQbE97GgOpS
b4+VwaAo5HXdSRgyb7R0KGyHeUwWVAY/3Ct9UyYznaVzxUxriyA+0apfPkezQfVv
7sT+sqI0QPMIvsnFD1cQMVozw2nXlCx6b3a8yk4Vl84m/xqUanbU9/tDWMuVkoRm
AITK7WBnS/+1P8i/Aw8tg3iCBQEL7t6DZIuwbzWYbBeYXESneC9iW1hDJoyI8ogI
i/d8GsyhsASQlCugpST7dD92m3uEbe6Oyh8EBDv5crLzuiuWdVEaktynvKA25lKm
4j3gDFbe6p6a7iiAagLSHVxyChOTtHOAbHaJihpxAnxepi3+jWV8IamMIKN1LkzR
upziBOIDA1q3MPTbZUHjx+HRhaO2NsbRjT/h4pc4ibxGPQHcIy7R4SicSXYnvHLR
lYgkMXeUG/c/JGiFVM5kF2CYuHNg1dxn1cqiGn653PKDKw69Y1+eHUxvbACaNDb3
wpJckDbNNBelTzyQNCTl7nr7cWSTOstLZ11Ho5QoWOuPhHi9DBylO/RXAF0KEYF/
+CCBNT8dGMnnK/8OPhE5m9aBX4Jkzkjrhaq/XutFUuS7MoI38NvJX+uqdKuc3t9X
FILBKtIAIpsuyBllVZUsShK9KNIrO/pEQTNnDaaBW37256V37dP3est9pI5x4a1y
Q72etQeyNqxJtRMGhX8k7pvlTL86k9UwNvfwx+5Isewn/mluPaysWPX0RzI3vas5
HHRLVRnR2Y2GNiBg2d1roUaXJ7MYxMYaqiPb3rPyj5BO8YiLiBtJCYTIKSwdyRIk
Z4gZfdtf5/ESFrIvunUVwgQn01Jx0xGXH05pwd6wilfQNKTRRENB4mGKgOa9pSsB
80IIYK1zYeq4G0pvGSENT1/S9kt5g+Mce6eFhfWN3aqQZmxOcasQX+9qbtD9PbLH
08IC43ULcZG18cSA9Fd52M4kOnRj5IuugvBXF9J6gPY1/mF8EBtc2I+QvCyiBG5t
1rKYbXCT4q1wvrzsK0x5+FsJb0nEsxmLk0J9FS3VxiHi4v6OVi5hxd4cr046XaFU
LDFIZ6JlAgA9VEs9BtnbU48xfvR32VBnimYcY7DHG/KG1un6IGvnfHmt/RKeH0jC
k25+7bzJQVZNIL2b+Yl6GMsEv4TK3wRF9325cDxENCUSrMZBDAk9sr0Mkb+M/km/
ox1pDg7EPOzKNaGVDEE7XUQlOIqQ+YM6BSzjmT3oX8xVKexxWdg+Lp7p38RL7Sx0
g2umBcPFWrfVJ8qrhV6WoHkAsjXb/QZT4V5MLbD67DlBD5XH85QYxLsSMm1Th6Kh
tIg5C6UIv+v34rf7rfXn4oqUZmQbSs7YzwU5LDrDRjK0RlIijYI52w0G1tuj0EEW
Ruv85xSlfAl6ycHOICRAz45xn/yoU+gPIISQqcC+l4g/90ICei++R7kVVE96G0Fk
TqcAJGYRR62NuZ8V11Ab7LKpMtE6eKY4n7pHYRRMtEPr9Iqm4/1jWK4tt3in7c/J
G1avNNWKa9w18UFdoRiFffRSDfxY0mTX4XhwA785nm1jAplG6G7c220v4PJnNFZ5
Wf03xOpmOaKW7ZZr8IDgLuuxalV5YzMyyln715VNdbUsBkvVu1VS0XUw7zDhMMee
AQ0qXZ/FGeZW229jtAsFZtH0TknjpEXZOaH14g3vrenXSfw/lE7b9PReQnChtnvV
8zhgtvMNs51R41o0RWBi48RiPEvA6aykwk57vqfEddA+uK/9KQZ+d9PXN4YJRvC0
46l239l3yNybExh6toNvgfFglklDlUAJIFv8bJj2/PsBBAKGVNYX2WgqeSn7/G2O
OtNemIwxTUeJEPxif0tOai9pRCc058JPltBcz+dsWliq6iSPgm+B5TYEii3eqUnV
IG8ZyRaIbMS/8BATPwNr1tTjgS5i8hA3g5WfjW8DpwbGVPpyOjH6z2sDZoPz1Mg4
LQniLpN+ozlXaFyHpHMHsN6o+sO2gk93SVbnUdXeZJk=
`protect END_PROTECTED
