`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2GPZK8k1aFZUd3yPowu982+zhnGTy9d6QmQ+mtxICNMHVAQ7pizlVJe7IfJ+wY1Y
OHtN/vCLHbdIYpCrSBwqZEmrH2A9GetrrXFJ0wDNe/fZ0hhAXEgcB19APi9Z49xQ
GlEheghyhh9Cscso+pR+y+N+Z6Sc7Be3mDumRzECp3cLfBEB4IT0h5tXmKS/iXp/
dv+1wp01xrQ7vM8AjE3T6s5BfloO1BcqM0WWpURA4oe/usc0zImBIf/ykpZRQYKO
+8mpy/5FIXAVbeyWwjFmpzc891KC8ZRyO6SV34UVaIJsb68glrJqjAxCYWDLG5O2
zNUUOIQRpPbHWsl4C64VdKnXx0emt2O1ExJIlAWJBQRbWUAeY6vUAXJkUzsrPBM6
GpaUqgU4V53Jr+cnEeSAqw==
`protect END_PROTECTED
