`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
poeztYJYFIE9P6ahfpncgxvyn0rpyCrFrEM2HJrKY28QYf6cQ9upJHjIbWjLLyh+
QELDi8SuepXNNK617Aeal11N/bM897gyNNLvnPW6AQdc5Rqk3rtH5xpROPIGTDZY
4Xi82lFD29F2KwjLldvW/4nzV8wAVeo5VZm9tPG4y5WZeIf9kdZ8AjR1Uyg2W7w5
m/BFGN0dxjfI17WekuhLRNp6HyBqxqLtbqZ0NvgdGxDTg+TE0ztJvk54ZPvyhUte
UH6kPvs/seM/2M1YIMCdqeNyXPXrs7eN+HbgHD8VML/X8SzZ0uuJ1w3GssU8WN3E
PUQfj0NT7EokAk1EFCVKemmnEi9g+zK+0gn/MwrFGkakkbsx9r9v5LGlESk7f0yA
IG7SmSG/skfE6guabnp8xBgGaL1fvATQ1YLx7qm+LKY68XH953C3OAkGkFREENEg
BnYJ4xpY/N9GnysnNTfajuCo+vI+ItM8vEG9+xvjoXFBWeHf+TLt1IdKJQ9pcU5/
g+UPLnoAMv/tPdfu8gmyA+RNGqlrIf61Ty7I6pCA5AtIDfVq9KmAYP30KYG05lFL
zGcztOa/R0iXxppzsXMH3c/rdplGs3Dh/2xRNk6m5DnMr9g0yOF+Y/f944nRrN/d
xUqDIbYTyMWXa+b/AwYlIA==
`protect END_PROTECTED
