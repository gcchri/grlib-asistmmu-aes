`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RGhSZjcZC4c+mJf0pLKFQqewSvoP8hSvDXzNgjX8urg6VFjLWCvbTvcCBOfTSNFO
11nalFG+FCEmG0EqYdNNWJZQlloIvZ2VVFMZWVm/HrN1td42gAxN8e/zARmZkrmQ
nEgVpks4yotypk6Ghi1ImIrgip7FbocYMAjjL2F3z/nzOpiz3xq9p0PU77/J+NDY
yddxNcet/gbyuLHaXoi+tedcfvY89iG0W6l02o3yKi/5T9KT2KyvT8Uwzcw4oooz
tvTsJnX1Mqkz1ILevHxj3RZyxhvuBkV7RDqkUilar6TVPKcxT6pJShJSVq62wCLY
8mv6LhlDd1fD5vzpRmlkK5jLb0Jq0sbdwGBu5sLpz70CN/gSZpvxlbuap1Pyttt7
7djJycKe1Fahp8R7X9+l+vehSl5vxlXX5fiXQKMHK6IhM4s8FPrpVk7qXB6RAZhy
`protect END_PROTECTED
