`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bFE72BFQ4gxd1+mEmfuXwM6kWEAW3FMA8aL+VMoJPywkLzcGJXR4zxuTYO3O7o8S
F1A0imhKUcbBji0wOg9aEo5BTwYD0H2wC6SSupmRa464K5+du8BnsIsjcxMHt2zD
jJiGs1HNhpR1/E+pv2YKHv11vCiXr45CkbcUMArn4q6MPSckdIvQPcMGVlKJHzBc
I1OEDWCQDmbs4tp4AVCJJCg0uOA5S0eObimjF2+4Difk4kDqzMGvqGG8sL5zDAJU
VMeg3EoFuP6N7AYBemneTSN6yZfQOjxffONhdIc3utNIpX1L6VGkxGs/iXkpbgC3
U1lOmhLLzuFOpzfB+/bE/OweZwLlwBsD8IfeWwsygfocbLQpL1ILGfjvZ5p86jha
cbaqnVWZQakHgCCwvN6TMQkXNJnUsUPZG6E0RN5ubNJTMzZtejLNHT3cL02Kp5p2
qE+S2XxUENw+5/l0TJwqGMK+xLY4QAefe2fZ/5pcqHmCbjTcdr0b5AKwyENLM+EP
QXDzHQ2qjDW9+68pfna2hitoE/IMvpdYaMbNIQlFiFboTZBs5LTFfX4ZeHoDdfNQ
/ekZPGHNGRRTR+s8b+iJJ9l31KPSxBjcFxZw9EhgF9EMvFpW2S55LS3f5lJ/NHb3
BhMyCcTCfIg0vQo6to2QkOD4/olpfoRwwf+4zbb2/TZ98xVgaQ8S/BPgU7EGYEhy
IPZuvLnq17WBwrqrHOQ3/+/aYrs8AK/YM0b/qtwAipHpcW86uttO4mL4wHVZ8CIT
Tp4r4rlMOg7YDQ41Ew9bu28sKYBU3S1kpnDKphGWOPVAiUfNRb1ahY9x+XSLWivW
+1fR9YAn7vmTUFuXISjXSA==
`protect END_PROTECTED
