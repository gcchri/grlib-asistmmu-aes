`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uzE6jcBA2NAfgr/bzZG8nv23of4w129fT4qLKrL3wD8sJLjDkm1caYwRckoKBtO5
CVYZYJ352imxYMWqh0VouxYSAIA1HZM5+uHPqWL1a82xs3FOHhOyJZMcTeohzXYR
zYYndm/Uon1TO1vspWM05NX0eIJQeXZ/fqrIt9QeTSlYtDzAtXYetd6UiuYgOUNi
G6X8+IK4BvZFcyCRrCVAmK1CgKEa8zKyDoQLSTRf55ZZUi4n/8y9HlfdQWkdvgCC
2aIfC4g9AovOHZIz4t16ACil4PFEsBO5+X9VGDZjO5un4aBPLvmimCJviFmJlOgZ
9WYquWzkK/O5COM77xmQQCwTeDFvfVSPMta+GR/qA7McEsJU2xu32IA7fapPdMZp
UnKax83tWN4e8WmajYNogvmE+vGeZ8LBIyaBVw470MNfydVYkJ7LHKssFf9ULflY
a95eRC+BODIZcRgpjbDODxX6YtBizw3Qs1x5gAEON1INMmGO5FFtTRKg/ozXEpSD
GZQn/ovyFsC/xYmWlTOeQDYlybEbseLLsbLF4ubBkMO8HXFa5+/zXccAdX8kV0ju
FCIMA3SFt1uthPaPjUTIUePYeAph0/Kq+MTNXn4Ow6ItbKo8QiCGKwQJWUnBFv5V
QNmcW+AR2TsZMV+KHcCrfHfntKgibcdnbw/ydUx0A+XoPfMkwvAW1m9BrG+BakOx
lNePyfx/3JQoZN1REDKaxSuUhmpn3dJYCqHVgDixEVzKkRpJZEczckaPI32l2koQ
B6Ha0e5h0hNfHfiQdpMN4StdQvLJKgmdmyqtmnPBx64oUjloSi/Mh62gsp1Bg5QI
3SLsB1aut6pjRXGZTyu3smuQWEzPPL+WeuLuhPYLlPCWey3MSdqV2yQFIVhu8g5l
eksm9yw7o/kK/q5nIKVz6YCanP2wuxD5ZCdHSfAjG0RrQqkvWXJeGw8Hq7t8P1s/
Dgt2StJvrfGUpf2yB0YfDGOn1SWc7I77QE6IHj3gKZw9CMy/5El9h5LDWniU6ffR
Fsqm9XBJAmrq6BF/QepFCjgPPALHMSeCecDmXay1trajJ4UjPrmzYsTjy08mrZYq
lomIMSfMso6d+GOU1MrXAm44spkkXTAsuo41qQyHWd+228nvS2R6wVSxzZbUNEz2
wsYk482LsuzLcRbUnViNjwTG2PplG04KKd6Izhm5kqVFC6ahzmU7BRzR+QfYux3s
BSKkayahOdHSQWKhkJDrZF+2jp737IqrFXoDynPLq087m907g+jB5IJxlOCRQt+L
32natoqCrMEFuOGDGITtGRlLXMbnucikhfqQ1Ohf3dfmztArzRrYsCpv1LhOnj2J
9fT2h/ruS+exv9TBJnUJmvi00RZl+wIKrG2hHjyfYyGOlwTrVEeFObq9Lrtx9MS3
/pI5frXAeFcb07/fLo0wnEPA1I19BFHxRsBH/IU9qmMZK7fc4y2s2f10f86bKUB0
HSRFDzn/lZrpkOnt+uQP4Zf3fSynkPo0CYq0OXHHkiPjt+hTMRWWv8WBw1pgzhcr
EBemp1avDn0MoAOzYmwsccHqlDzz7KFlzOBCpvab9zCoMZyF9I1E23ADyxQ1ioAE
aLXfKlq8PfAMXQpQZhmhIHe4kL1RQH7qznqLU0xn2Q29xTvI/7ZT6d0bALeTGq7+
8QsGTLn8/VZvxXVz1qnyE8OzN5o2tM6+EbfD4avysqnHGU3dWx6bP65NNlfInbZ/
gXVle4iM++nelavLEkHDJaLdaoMTNZGAOlKgGkD+cj7qnmoJIKtyGglsZaOnIbZv
2pXr4JmVXFpUdddk0Jky0wHzSVBrT6xW3Ui9MN1R2euAuDVBsS/fjD+/5KnTLjOP
EUEMQj5e1TYXhzhCEsoERmDB7HSDVpx7L0bgIFVG0nVnbHTGsclki8lbmoeUOZfb
`protect END_PROTECTED
