`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0a/Z+k6qUD1dftwDrRSSXfQs3PjDsgNc9Lxy/gurus+MMd2/iqRhLOs7ZeqW0HN9
sLIibnXDKNIkh+DwI2g1Suz2EUrYvpM29HEjlmxXxSLsBFTtxJHIOqAuPrdTluUr
2dYs4/iKC8YYWDlLQkFB/BWhS+wN+8rmWVEoJDjKLuy02AJOwthnvjrlfxSLIiUt
/yic8+O1gfieynAb4G0mt9LZ0VbBXdPQQEVkmdw30/foQoWlMZpGWYjPFIY34mSY
zNDKBo2Q3mr1Vtd8J0lfm8caLRrJHOKLBkVycFo4dIVOG24w03nVmILloVQVmGyA
2DD08zQ5QikY31ocMB9nxNeGna4SWZiagEz/xH95HphyMeG2FaegjRyYkN9HScAJ
yG7XhoaTu6WudQyzPG6uRg==
`protect END_PROTECTED
