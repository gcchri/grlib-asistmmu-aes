`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+mYdKlnNO4GVaw7xAnrHS9wwyd+MhjNULhQQDMi6SkNdwriPo30HBBH4IR/LSI9
A2z9hioISOPyU3s91JZxViXlnMqeWCETGDeOY91oMzCtRT9Xok551BXyuMKJ2JeU
hGb4nVts65vYLq7ICPTFNnK3zv6xhfEtXT/8zmtD0s106MoIxCdDDqkNqGa35+9u
KLPbkO5BO+h8SGN54GPsY7zcVT/m9IHdztx1vG0WPZGNL5dB2zfNJWjS0AKzK2vY
vMLeeKVrjf0wyGI1AnzyZsy7JGMbw6fLzEeieF8dFaMe8HGPLaA1wmFUharMslCl
beLXLe/Z8nT35ZyAt20naKDhru4npQMXm925RftH8V/EkIOVlzRzvwi1mdpWI7L3
h6NZnCtrHjzAlP2GFxkt7u82WF4dt50xtpKO9F7cwXJyVuNst2fiHpusTXNr/n8u
WPCIlU2Uervxt+LGQAohzXlvneYrPpY+J+cuVQeCfYc=
`protect END_PROTECTED
