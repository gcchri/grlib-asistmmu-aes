`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69VJiZjzHf+oj1NdWs7GeKc8vvmnQIOiSxiFjAfpNQrTheR3RjBGvF/OcdVjsVZE
6uwWCWW5TOiwP3Pzo3NDtnFZ6MzCXujMtkZDALqgPz4lICDbgtw3YXWdHR/FwbED
BuXc1G1ZSF/GI3QeLe87wAfaoIAp5mYC6/exQAhDLcEqdILqFi/jJZxMl6syiJpQ
ikxA07mbU5+HvXOMQiKbJ/CjOpMniyPXe8MUVxf3mC0lJfLDbSB39AELDgI5D/Y8
fI7Nv5XpncYOa9guTpLt8cQH5w/wCwIQFP+fj8Nqp4y4L1Pdwj/qfkZ2GbURgbI1
Y36BZ82W4SbaYZ06vhkg2Q==
`protect END_PROTECTED
