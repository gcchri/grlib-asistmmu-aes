`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qAquZIm6QeyDijTJ1Hhq2P12/llp645TI6W/ejfUYI+vj8oh3uLJV23XU8AN2Ym5
IE2IrPiRXd7MCiNO/aGCJY5Ew4Tt1Ank9VRg+VcehyrDcaXx+GCHwD5YMqJMwadg
lL7/oAD4Op+TSA9rjzJSpzXO/BT8TIsBeBgwb6Ip5RRUFzHvWkP4+44rK4khFOnj
TBrDwlojNqG/3Cvr91uNPqgfEgWOYL5P9kuEF7AYi3jxDpC+MNN8EO4UnFcc8vaQ
ljCOdNP3xDvLbfFTQstP9p9yO2q/sM3LzBSgsC3sINYl59ehKvp8FcMWxXBh59Q3
RvY1ec20zITZCnG51RQJa1esv+J+4gifweBgtNsSh8K2woVI7ZiS4IEehSgtIrYk
DoLE21/XE4DrOX0K5YgCXw==
`protect END_PROTECTED
