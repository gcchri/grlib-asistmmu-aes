`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPo1QFtE57v1+PgR5zE4LzYqumUl9Ldn4GetqXHarZdsa0Jy9MARjkeGXt+rbGrN
aygLsRSuEzoRkMjLJjGXTLJOqsRlZsvkAP4xzD6kkjX7EzKaha0oQ0GgOWLxDT3m
/TtW3sN3154FyMxrqXCBvfcTx8V6mzqBMmas/wsj+Y1poHMCVk+pQEbxawaO4HB3
k+WRyGj13SBRBjlDlJTBb/ZKgUMsEdUuDXw1qwM2OnssevgcHcGI2r7wD+om5c6J
BLSxUKilN1qnDcxnS+7RYdmZVeGtMH85cVy7D57BLR+D2nkmzIY3R/73zV26zj/D
DNsrRDpO6QZEfI9sApMDtVNNOswTx+22GVwMmasKVm5xxyAPsKoQgiTWkb4ABlBg
/LJ4tzlXtFDmstij6wcXdiD+R9ltRNeiuO0Gg5DkUOM=
`protect END_PROTECTED
