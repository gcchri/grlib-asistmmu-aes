`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09FgGpXp88nnm7GkUtzNxEALinjtO8AUMc3Q1B2AfLYaCChSHd/RvArn9V2W/Xfh
rVUIa8EbLvYOzoAKLLN8sXIZ5qvPSKKC/lzrMI1EOCOxQ36Zjhy8Ndxb3FZWoTeh
uAw0MybunCeDUqU5fw4ODZQgdJahUbGMjWdqXNHxZmZJDLTW7aNF6Nv4BuXGYPNW
TACDTducV5g9n/LgUhOPjV8BD0YqBRlvV4WhCWwCmUnKmSBxwnTVHXX9+0gz7Jx9
eNz4i9m2a5NJVSwHxlY/lumL6PAJTz0qaDeob/i8iwc9dqdbjDi5YqnMqw3hbzFO
TieHik/BxJkTmJikqeaeEOdmVEMkK+st7a1wqcX3n77WODru/hMjmC3fzqnU8JFr
RY4pOukupYyX04j64M6bqCA7y5xG/GAtb/QXQVM8wJqYB3c2PgxVYTocv+cdKcxe
Es0o3gGg2XfxSF47JBh/07neGAW7gMAryht0VmVhEAGt0WRTOioCPWCJ+XVBZ1AS
AesAozaduQIE0Zl4sPdJruzVN9fjglgH7CqYEolHERk8bHky/v3YLhTZ1k8Az8/d
sRVzoU2gd7TsYW1UvMDTQeGhXje+tEbAFYl4TmNOCiDqRX9Wad5+NVFTNwRdtamI
3lybeS+NWQ5lK12dEv5xjoV4NCR+NgJULhWa2kJ2+Nk=
`protect END_PROTECTED
