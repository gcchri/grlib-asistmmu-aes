`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DYNbrdOgj/fUlfqE9yubn54+wcXIIbZntiEQ19YtsZJ9KzNCjItIrLnP9ICdtqKW
iFSAZCZl3qXtGaQ4dsGxMbgLGlz/sE+UwYMyWD7aPwyXzfBhTEYAZRko2XexF2TO
hcIsf6zHXU7OgQo59xWKoVQK53iIAeTxL2vT3XB7B+77kLE1L6kiE3HrAzdZPK3/
XxSUxJEUHJgIjGp8uoiQ+gDpSBNGQ0q6gkLcHmQAa9gUZgGeidMiip9ujR+MNv90
`protect END_PROTECTED
