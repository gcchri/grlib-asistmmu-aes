`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xc9za3fwo05Q4CcntGFNtHZlC3jA8CdqklYJTcG1cm+OeE+k7FB4JuR9nyRKwq4O
XR+lcX1J/FzZjzOU4r2LTUI5QNCKskHp4U1uXYd23JWG4ukVka8Gmp+uLYqWZjbF
6DFYqSHz9zSq09WIJUeDhEYwqNhjvmmzdoZ/w4vXVvHrcnW3oGGw7oxuny8S+4S0
VaHaoL97hc0ZyFyVm4iXLebxDg2lv+Rrctvi9QVPXUMgLCqTV8GnnykvgkejG3Qf
2rAr9e5ZFic2k/5C2BR695QbjRnCgVsxtDxnIkcn1+ueAuFFIuFUdm8ubqB91Kp6
7jxlKssJZEaAvaGIqGUfC9qLfq6BG0IQggJbUnsaLnNNNALJkXdsRsS2hv7FT8wp
DGVSZ0vHNBMhPECs8HoljA==
`protect END_PROTECTED
