`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kKr+21J51gEzf12gKNkiNUf7FbxlthwWfoBJ7usyiDquJr5Vj1LCIKkqqjlppQdQ
tF14zw9RRwLxWyWLVVwa1eTtcnmoG+yY6GCN4Q1ojlRdG7pcTrVUk+g0pW9oTAx9
uXJZZ1gOett/gaRgMPFrezpl1v3dwRBj8VgLjIjrY+NzMrJoTZNsAAxgu7v0VsMT
UaH7VxnBCa5fZYLlgQJfp0RspSMt5AwYON9Xq6JJUkyay6+9oCW9i4xJd9v1/7K/
bN24HecM8ZBPaJNcHskAOgu2NC7CBCM604eOUKFxo7h3HpEjBHmC7+oxwuA/AyxR
p6NU55PNiRt2NuiyQl6GishotCyJbq5Yr1j5wTJGNkjjPgfkGNjXKQ5BZ6Tvo5v5
Sc5U7N5S2AP/2SnZdeJtjA==
`protect END_PROTECTED
