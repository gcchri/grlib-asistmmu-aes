`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0t82oPAVsehQUwwMtBH44WETQ3MO6bAewfBJmgSzH3mb46enE2bTENReFVNU2gQw
Rx8WvGdI0p9/VeWDXUyJTf7z9b+fN6xQrq8f0ohCGb4fpi9LWW+7FVJYk+rYbhgO
qecw8VhbzWBCxDrJWYkcE1TKrGJlrRABaxAjWPITddjmmVSkjR5k38y/oG2XzC+d
I3SD5z24D5sC5u+zqIc2iMspaiftMrHlvXb/1usd0HQOM8MrZhY1nHvwB0O6GMt9
uCVnHtQeiN5lnAFY0nUk5d2xX/7L+/f2K/VY+PW4ghKHFaGv1njfWRaZP+Y9sfb6
xFyn35hwci5N54cjNpyYIIMXr6+8bqr2a5ew0bS1Od+KYNdBWiw0jTV0sx6yWQ/y
n2pejmoV5Ziz4L+oMYQkHjtyOo1+ygLl/AcgoL31718kEXJe7ETtlHsCPogTcZHi
FNv7C7dZWVuEMLKY7sjyXL8Tw2jHXQ6m1zdc9jt5K1RYm+jLKNq0Vu9cr1ntoncm
83nzXwW/DPTSSYabd1LHrP76Ql11B773J96b3tkvASOb/5FlzUJtbtB2XPC5t4NX
ClD2xcek54/STBSLHavMRZTwCLs6BfjCkv0E9fxRVjwWUAQQOB8DE4PbOjcPxZGw
49Toa9uh02i/U9US6ax1FC5b9/zMNfvcnFLhPfSKyj4EeucTTNcnoCPrkgfjokq0
tlTUAv2tfd8iK4lImV79l1QWcvi2VBqGJ9f/7ZNLmiH+acHz3eaChMrLC/Y27POd
kuE5LOJZbmMwLcizhIttMcCyJPuYyp3skmufk9zWOfiLMFUlDj1EF6GuqfvmcDx7
Wvrtj1svH+iuy6zNc09XDgXFkx/E4hyrOxEtBg+B/LnQQvCScMaV9iXlrnkCCGcr
dL9grXYa0zvIrLYrxl4d+ZozKm4op8aRC152FbhgiXOn7XmSbcKYU6NZWITSHtBO
MTuPdR3Ieh/kQR8Vi3KvrlJjjIScoXNDzwqTlXJCCc2Uo5fWNEPibdkDzSCZhQJ8
OBZseH4nk6rAtLq/nYDT+ejNHURL19mvpMzc+O3K9gWZ171ZO/vC/PZ7QXqjsxAD
ZadjqeNoUw3EYA926NRHvypCXIA4nezIrt1r88XhZ8bQRkBXd/xB7a6mNIjo7hvh
BY+mPLDnrHZ14EGqFT8gDK6UnLS7EXze5TIAMR1TBOAmBbsuSkEoG8o7hr3C2wit
rsqjgJ6wY8Col3HCERlYhOmR7vTtN6PSmagFULeRTFGWk2brbdVTYgslJeP78Xpf
d9rbd9sl8XhoAysWaw94jBcvdUfbVQnwFbZoSQxQzCcmGP9CO7gr7W3LbzPLlK/0
MPHJgP80wC3aI1eoTuDQvxErSxJEwW38hBJoglcAnvIvQ8iF+H1wKSj7iFOkTq12
R2TGWiF9dfL5Du+zdab9ClyJQ1u852yz2vqu4qF71SeQbifWpgzd0+J/mhUwSpY4
IQNGzRcQLFyK7DkUfXTew9hA6A9yC+dh4MlYMdio0MhA6NLEAHPNXvKvqJ5w9Yik
eYP3VfucS+dTsKpoVqfriT69LHSuNLwDqWSZoB5lbdRlUGGew95bXonU00zGQKee
EcZXspUgk1YVDD+5Duo8hfzChQEVn9WrhpOcerMSLzHg2qjaV0hZzKPEsvD5FCEV
sMCglxmhP/6+DoQwJW4VonNrra0hOhtU0hv9Yg8Vs5r9wzXpfe1FGUf6y471sagC
zWz7FjU50g+i6fHOPsZSfOvwAoEGPLAb6dkKn2vhKNADycqYotglgp8ROFHhr9S7
XR7eCMKpDtcqs3TnKFyw3NufrKTJoAvGeQv1cyO9YnuuSIL8CsqSCqYsc7nroje4
+Sz1K551bnw7fUydwyjjoMQy22hQs07K8YSWvVwyB7udv16fdBySgg/5EOePE5Qi
PjtBOd9VnZ57TEUd8rHIwAgfhmLPyy5qMSTON11CyxsHeSnN1y7K/Q4OhAGdPIxr
GR0qlih2r0jgmsMvCutcf9nZ6dWKI2xj6z9qsnVESNyTwFb48PgYu3tSVB5S/0Kd
r9PdbpRDUbqNvylOZ0A03Re27lCpuZX/FBO1kCugMKamTROVGlJeZ4w5Kkw5XFDl
qThX2YgJz0VPaZhAupuX0HRFKDmRsL2KnJW8osj5BobGYIcJQbW4FJcyHRdvOXLH
XWNKt/KGgjphWc3GALvcVKhQY/V/43WKgVD9tCaswNVfAmkM7OLUCDgfLCUF5ULD
j2Y5eh5ICOtPli5PejsVmpo532nRJt/zXYpL+0Uwq44SnsfVHbPMx3naG5LqOp3c
7RCbUdY+NtXlSqU0m3ck0BkPCj+/s8ms4aclvgoivrU2d7kmy4PfMPaksLMv0YGI
SHwrxPUCOLJfOo0q41JOPo84dGP5/8UF1HtUlFX9hUIo8pTPNfzhjZQ5IuT+yUWS
2ZM1dIIh6/Xlt20WycjVLStZwPRNJBwG3bw/NrsyoXUgBOMDglFrucHs/vOrJez8
ZbBTTEoMz4xK0bcxzew/5XceAhzyvpWKtZuZl4PUV4RyhzTeJ+qYZQb4OX/mPR+/
lkda3LS18yAtXRxZDExsQxOtLf84NT69SctNOklvWhoIfOV1eIVQbsZ1gvygzCQB
+sc8UKMZSjuBgkhx4EtBioIYkWUqJrG+/gjMTP4bR3cp0oa67PsXvwvr17gugppg
SYcf7nf4hU/3xHcLq/1Ry5Cx7nQdH9MrRRIvOhK5ywoThxQWGrLGR2+ZZEghwd37
/R+OhpvRiFM0S9pL9PR/EntdoOvBnW0i93dqkIhhR2azPMgcas6IxXyvOa1pB6oc
JlO7yebxAzy/dupV3QPbb+K9FpzB4545CTTOquY5+vdcOnl6c06V3f0/zYklq7AG
tMVWlW5YCksH2vKb7KEngxor8obE2a294E3X4/A3miZXgSJlAuJRLJvU91KgJxuX
6WYQnnu3oWtv391NkB/9XQCW1L2TawrVTr60mCQfZuYoCBUNbAXSt4cm23Gts+tl
1hVkW7Cs+/3c3bOUna0UWY4TmoL3AW5+tlasHhFA+z/BB4tG34FT3BdBwCHjLwXx
yRReiesYCIVHG8Zs38c5ubNoHuEnxgLDUKUmHtehBRy/L+EbZeb7LIqHESDoMlp7
+667oHMRVlg7Ucr/ULHIYytZtFxOwi7IZKG+pLTzzm4kQKOU7n2Z1qQQLUAUx/FX
RvNN3wWNMcN8uxjIruVA+1CzJIp/oF4wr9M4uvTJ9ZkEVFSQPsp1EYErmu+vmzTT
a5H6FCgPWKIbQkPoTyCCvOy4RPFfEo+WxbpfXL8+pubhsBTPgXF49ghsCvTMIuRk
4Xl2SfACIJ7VYUnORKtkwejo2BXkIZCYjTrwOKHA+xPc8Vb84ZHu1Kx9Lg9F3pn8
bZMotAidYguR3EVp2ldAMNvnwgm+6qjyIQVEgyOE7Bl3DZ/hpCFnOE8QsGndBI7/
yX8nLnuX+YNI9AtDDAO/7XdYFh0b3TabQFucGkolRVZWnY6ThXc4RmkfFLE477pV
ebbghSh56nHH3CpMEB8EVWbK/3SCiRAFj80poSfuBYAxdupeiyWeXx/e8lkZD7WI
TxJHcjFCtCjAFN5eM7xiviYajMP8kCmkak7tNLGHbx1LPlc55WYv7j+jZv4ikKHL
ZKGkxYBu1LC2pW9NUYhAmiTcWVvf+3TtJS4A/wVSqzhmXij9cIaFYoXAEoPEsyHz
WITSQb9Be6Yg7moPrbzDC/fR0yuEZD0lHS9hXjGCc0jVKRqCcVWZqRkGmopFUVVT
ygZVLsJ08+s04iICcoWl1F+NW7Wd3YvzI7LU3bv2HS3OYCMDrQ75dROFdSShwrfD
5L5Q2Abdc3twjymtSNkRdyBK7oXgsdlq3/Y3187CUIq68aFUhJDck0Hk5Zfx6sCU
tAmIM8P6/7JMbQdEs6eR0IBWLwE4dDYjE5amOKWAa322gfqgiVot1yioInZ9F64O
v17GGfuK+y/m7sDfRU0NW7nSJC4/MebP6/my3/KiTuhGF2p9uyht7IvmQ2S/YbR9
BASb+ugoAq7flwXKMGoUXtf/2KT9Yt52h7WuHzNAlmRKDmfe0bZrgifLiPLwqZxw
KZpFG/DVq7oI/Ca3u6LkTOD0P3UlcdFBpXTAGNRUTxOJd70QGEY440t/jgD3pGX8
iFihRQm4/TUMLccrp7pOyyHu/v3evYOrzNlqfNyh9QUvzwPyJ8UVJbk+fOarjbat
bcB++MYIwqRkVKxV4BlDWJfBkeIYK/YrUpz2QHKP7qBlYt/RHMKjzrqgQnSD7LNf
EN6hHuE/oFtVhW3ANyWNtKU1Tfg/2a/R0Yx7EwfG0PJBuesBgkhMzo7HJg/w+bIB
F+sS9FapK3v5tDr5fGAJa2Wc7oShQHHcA7tOuubpjb/hxCksL6RK0qHZeEitGo9c
1E30yvKl7DFz7u9vEj8363Eh2FXhGTYKjBHcceOG09SF9qXifcpVo8ZX0+75YoeI
R/SzUHUWATiulUBPRxp+wRmc4LtbHE61+iuJLawWQ+2lN6nJmxvTI2fyHdOtorKs
ElBOFMTRgTPp0TKZKlSqu5qRfG5NDzZZR/z+nbb7Z/NvOI5xTvzq24w1R2L+esRt
/6YJ1dETM1bgvfYUrauXDJ5NpZpaGqEiLVOVQHF6TW4LcWfSfOQHGpRbl9hYe6Mz
Zce8nIs12J1jAeBKfi4+CNs0atz30TmCo+tPQqxmf/sqkgtTKfSHdiOjpCbvgHqM
dgvPZyTCP/iNfYz5lnV7CC5WZzX0CmwDESfZpQFcpG9Up5snDHl6MExkqfcgsp9x
p0QCcOQE3TOCrgEvM5oScDRjC/PVzNAxwq222iNLva71+SDFT82/eWUuYigKxkWR
USlA+OHzCRTSIG/wpYkehLRdWUpAf34srkyvhjynLj3KsO+aSsIbkGOcFaRgqs2D
psQjf1qF/DsFxDPm20pyJTIjrPou8E6UiTYVwmyKKVZtrtvysyJ8N6UOvd14+2Fy
JHzx54eHcfRfDhsEQuvUeI27ItSLlKT2rQXB7viLc2VhLqeVulzjYmmMmOwSjN2x
dsGVUgYSmEqTriZqah+UVMPSJztjg4vYKD0QHZ0TNZxXZU8asMqCjHaE/QTH6niw
sm1FCtvL6oNR1Xj/pViSMB/OXi1QB9sNYoYiEkYVtmt/rQx7B20ezx3ggPkWzOaV
TJ7Hddocglp6e3ukcI7Lz7JUCYbV67B3K1CQdKyKvMScMz+jDA3y7F6WVD2zK5UJ
wKCnLVYEw6vmixTlxYP/Wfxht9RgaEoAGM91ZrpbZFKjsMteUnFdX6TxYbqfVmFq
e9niT9HzsF0gJ7Hz1wkRGD4PqnKU+UUh8tiA8yYtmTlvUDgQdQOA2KM88ZMXsOik
5/uKg7gpofLq8WnoCNU5aWhnSX4SY1vEpUWh2pMeT+Yd56iP0TbTwcY4xFKwpIrQ
w3YOT0qANRyRZrj3tiNvsveG6HNDiwwJCSoyFcFxMZtZ1urLjjqSvtvUxj3tggC6
sj/m0FEIXOifGTWS+HuWGyQ7uJd2+bbxaDUIILw3oQ0kWGO25IhdzUxZ/kxX8P6R
3bSQC1j0MQzwfLVoEDZbSR+fnPYW5wpyjM34mKBCF/3NfaOXNULswHGRisWH/dnr
yQm5ixgWJw2umawncXRfYrk56ifuvYlJkbJUUUK7rW+aREHvFqgHMkMxS7LO8fbL
w2v0LN8I0ZwHP0at6TVsIwrV13UeA0XiGvhVXh95zKRdQdeJcTGd6EZCo3oJI3au
xfmUdHYNsr47mLqkK3Hep9LtogVbPmkwehhj/WraB1NC67WmGLeRLzgHTsK9M7ed
MEP+9Nli45IczKVkpavDtlFKmeZWkuVA6JqKpQ1Nu7H+ZUuxFH83golupHf0TwqD
2Gt34xeRVHuETaLZJA8ywuk5X0jbG6OfQMvnJNnZjJM89926+6cEfiYivBJq7uqs
Kvo0F5MyXiaqL19IZO26twqPLU21kvlFSDsuwGy4Yya6hG9AY1KmiuSqWGn3zRfH
nZQS34WKrSxXQAOdeognMvEVglZ0o5wJBBj89ieRhgTQm9SclQdcCiA5wyVm6TKp
aM/H+5DOgKrYGHpkwkWC3L0oum5+tP5F9tEEcFRy90NwCgw8iRqSTrd7s00u90b8
VlFlV6bcVjOygf59FgehWQ9gqQRrcD3XfVJ+4q93/60XbVZwC21xEikyCBHRbIN2
u6F2EQHZDFkiYTYNTm4+e0BU1Zgm2VsVtYwTYVbqy2ohV3kqPmHQFjtYpXB37dcs
+QY3ekXGJ2DrkGceVtj8deUtxmGdoL+H2VQBTSDr780VSw4Sx0AgmF013UG2qN4U
bcMYeF5zHNUELVvV3xLIqg8lJKi3oz+jBbLalTIQXVZjCm9K7qa2Qzaudj0wUJ/v
6GuDXnJYS1VNPq1xYtYIfvsjVrPCgo8Wbpz9cmbPdVO65BrWg7ecgtNrU5rRzN7j
9mpUXPkkkE0uvegijXfIPOtB90AetvHr3PTmokTw0PYK7zb0FmHW6OI7W+cDNO+2
JSuPul+Ue9AWtEIyZVfOsYXnW6lKLopLWZysVyBB+mv+Qu1N+zYsZyq91W3vvbv7
QlANkb7HpGxAMwRJuP7H1HnGxNJhg8sVxxfNitddnszfI8ppxTfnjgFQIGWlSHe8
TtL0AgQhg06TfNhwavvmmgTEJJQX/Hi8mZjwLzbazbHdK4vhfUt96rTFoqymjB25
H5EtnntqeuAws+TOslaw41yjQ7a4iZnGjqB3B1XK8B05DKRvSIJc1zc5NmtuGCSx
aSsB2PH1gCV0vaVFHOo+4/fzPJwNb2xiE/yRZTqG+4/kjsjH6g1yFHYZoobzVvuS
VVXfJiPUAZYl0HJ/ve3EzGfm3WE/AnK1MA/Yvhc8zOfcdU+ASHnI4b00Uneop43h
4Ew8uGMTKQAjpllaxBNFlfHvUHYxBBvacCCEOtn9VPXJDID9XFs2s7gyiwF32PRk
RC/enKqASZ3X2sLzLN5j8n4T0rY3KfZaNKjl+aH3zKysysEg3cgTu9MVwLpHkMYj
JRy8nDXlhBTdJ8lIKm0xFFVkB9GqdbP44NtE9OcsavZyUUWkKcdJVcBoxTQp1kRa
q/Uh+Tj6UOO3eR6mJR8z+SyJ748GszfQMxo7PToSsIQwatRJD+EUEfziZg9i4fty
3UGF2bTZDPpPoMRt/aNnjwF9bOK9QOxvdsVXImoBwblIfiP4o3zLHOD10Fo93nai
KmaZQES+L4sgAPCYNx343WTEn6b9Z7/uRBKqc/ETTUbO36I4FeGlALkG9K9mdGN9
4vM30gP0P6gr4e0RsXXTEovv3581isLWYiw0PMXNDaubdJPtm7f+hs8dd4HVFULq
17I0jYRAbtPccNvfuKTipDpOrtGwRfDItc6q7AeNJrYXTkwEc+ajcE6kphSP2sHb
aWrif1Q2O5HipSEqiUvS2wSx5oCQn4UBkqT0lJhDGrEvcNIpMGYg/Usvpw6FsL4t
3fpLyJzPqHxBXIuKDWR5QLTuiMqVnkFP45N5c2E6gV2QsQAhygsLIvOQlfsd8k8h
lylZGt7qQffauPPzwyMu08w0j6PlQ7H2XkU+oetfKGmJZ3vjbjb7elt/rnZSpw3r
eoHj93KHNIfnVDdQ7m3reT3FEK6JwuiiZfVax1j2y2MgVBh9uf7+fkDAgUs/HeA4
dG+laQ4XwFjK0sWp00sQtjgW47MSWQ0HyZnlyiAiysJDEjOiDVvJkaWu9gBF6bzc
8AK+uXcZyOYqptV5yjtz8qXbS+tAb0ytd0CcO0Mc8LtcDK5i1eZ8K09gN7ZeOH8T
j4QbzvfT8Gy56/dNUKiMk0W/kzIIcKdm5nHJacJUdqImdAWfupeVtMyr1WL1J+Om
bbs8CKWEZbBg36tybMCF6Pl0uiIDAKgmGqUTrx+gp9QKdDeu0HL8hyF4ns9yLVId
mGFg37pwm7iRzYddAVYP0kR996kw7dc/ATytInga6u4RILaLDSEX7ejmMAD4pOYS
4Wof00ZHw0cG6Ozah/7Yy9xAbvdKP/W3CuOh4o6WUFnHkjhRpY2VCTsQpb8Ohq6J
AcbM65zYvcaBRtUcZsmFbu413zQujyMTuPGgetYDJU15xXF/mskSHnJiGdYJnrC/
GVSlvLIgqshgUpVwiDAD/3+5cDMn9E/HGWONqOewrRYQWUD23ETrKPrigUqUZINF
U6bQN7vEAbYCjNgPBNINwbQYTnLftDyY/3CVTU0niL4uLbrf70A3xkuYz03v7z/m
WvUEmEe+RWQyCAi5foGBH39jASmr2dwe7H3QWckW3m6gvhsll+GFrD/Wua0eTcLw
IX1MVGxcUFTNu0rWqytSS6FOyOBJgLgu57b7mk5A1Y/SKqKWhwpLjbd9gmxI+ah8
v482xs3Xnk5M94zGdAsfJfHZcmA1wUN3lbxfe6dCszQB9z4t23OfBFzm1JAXFP3m
pii5oqStLx2/v9fnagUknTBLliq6NyG7otjZZI3q0pIEiwv7szuzWQEAr9iKMVR8
+V66iK+wcStwJ8R0/i8I5/TCt4UePVIqFZbea6vSUaV1TAW5GiO69b3ziGliL5jt
Qmb89EpMpPnCnVI25naDAwtuB2BSX6tYoABj3c0APrVJ8O90WhHOIcBw77mlDLKV
gKdf3yjYs6SbmXZkOlWWQVU1m7+xVv1SrhWY9g6MyCoVxtKnnYyoFmt5bsAWin1j
Qy3WjmifI2IZIDYOeTKV2f93bDE7lz7eNvU+DcZAPKIiOW085yIp5TuQJ8QTLS5s
oRnUnzSzQ8yxvvRUFp2VR2zNCF1wWwbN8MnY7ZPpRYhBYfNfHgIQc0fOAYLAnIBH
Tlw3V7RNX7oMX4bLQ0Qo5K2tiJf1PRDllFTavds5bIK8I8uEqAjNbL867tBDhUbX
nhkBfve2nyLpoyJC+10jykdVKeB/cz9vBrZUBJ8SYfIXEj26GyPYn+uBa4yxmCi8
UhxoiGKVvnw8M6Qy2AxHP05LOwB6bbzhy5uMANXV7Nn2WIJf10JBIeL+5YB4Tza6
wtNAL0AaAaR91lTqEou8RUP63VZJO8yXkwMtk4rc5mbrxq5RtvEHf9iwZho5jS9a
qIWbSxoPZYZX5y0TL0PefmwTE/95lNiC9wO/URQ5bcmHG41bhVoqhqrVspl7aBPr
cqY0xCyhwjKG5Fa1kC/rFIMDh2xXCTyoF1pUtb66OnFiTz7TT9dUInspt1QPsCw4
LYuh70M5Uj8GYx3bPreERtb1P01V7Ahlh/KJfeo2VbhZQHCdsHNxp8iEXuPAxX8m
ibD3KklBrinXl+2DCxZa4sU7CFB2AHXrj/m3FkH61gfwjJyb1z92BONvkzWB+KyS
wldAY7x3oKBLHM7PKhY5bAqdhouWsiX95RLzubkectOeo2xZV+yQNR07MoibVDGi
xDJZHLhVOUrKFUJMLv/K7uqqJbxU9tHMDnndmkjSTBKqxxyQjTffJcUQMdGsV27g
v+C8CBhrR16WsbJXCIXPkcOA933ve2SJDpfASLjTk+NKbbKMlvBYli8FDI2a6JaB
t3SlQbInuEG2oahPW7tUol8WdVjja87ZLzA6DJUUipuJfK8DuWL/3tse2e4xLSAX
7fxOUXSErQJ8wbRSduVojIF0Qvs6ZHYAzUD7rpA65+iqfXvIjs38HlkoEkG1ztUb
a1+d3Cz+mkPAPqf5PSAb0NHAEy/94v/OiN3l9NPp2diP9mXZJ2tUIi5hkvsBQlbz
EKjPOa+gRlvhmSzF7KC3AsGkEomYEti+LGjV4eEDtAvoj1PEuHGI7su6j+H48rHj
lzWlFJ7a2+nAS72BO+PzQOA2xkBSjwC/TfRJNsBNYlbIxzVirRXNa/7Vtn5yU/kM
lu6UcY1oru2OhdfgKhfT00GwQ2aUUDFn+VLU0ts/r7y+zljJk3tVRsz5lbjvGP2Q
iNkQQnG+97a9mCqIb2+OC9cyOCntPOPQdAWpqI83kAnU7XSLR1DMBknKPV2fOhVv
Hn74M31mAjqz83FsGYMyHJ74QiJ9adcV1fhQpo+a3FroM/8pz/b62cBPgvU/NIO/
UUV7ExTV28RUJqAebMowloMgqRhNiR57ym71n4TI2hr788bpWtfguv3LoaVaqVqL
B2qcwXj2YsTZkSmi3YmZzxtc3XdKHhv+nUN0npqQTGazT8LL+gLO9u/BP8OriP6k
860Ak3/T6STZWhSmKi/up5As9UeMAXRHX1I22Hb13xrH7k9Z9pX00jwiBY0eBVQO
/LKEoE355UXjUF+/XIaYj6N2CZKCyNxKtCs6WSmZWr8ZTxKM6dL/IoRurgF3Aj1+
k1kmJo8ZqBjI0W7mvfmDeAlJdQxr8Ive+VqogwSICyTVFPS+CYEPHqdiA6HQH+Uz
tHAkEkEwstdLoCb47IX9lBnXRKrBTRkZ/IL59al8hF+Bt5uDG4+lxudv2R5QqPtp
DtEstvMt7dVmX+yR7Oju68h9Knc2X4Qfnz4Zz+jZ/p5oJ7qqJWed38LsSKZbLCOM
QLQEnVQPTRvQp/mLIcWsimAQJCmpi2F5HNccWsOesvcS2IShVp75Yl0y9Iau8Zkx
Tira3I/IfJ1yNjlMEXMHOc7V5wNVz24vLoahhKzArSD+zhz14L/SCk2VIaJwRUGZ
5g2xoInAbNUNMgkTwYWFffLUGRLXynkwjylNqSfYF0KCxKA74xMEVk6XbYvlhiWs
Plr9zZLP3h+Uxhbk358BCEl9HH514yY9YejUBmo9KIZbrOGIRnFFSzgm1ruoiZFJ
XoRIucZHRBiaZX/L8M5bfBpgNifNc59799aQkkgGYLEkJeaORsnvKSiPPyC8RXBu
FyGdPv1f8+j+Zmpz2c9yz3vOrnY6t1GYgkY/VtoZpO8sZAiLXwrG/qyCeWaTSwJb
TdxnTpeFNQ8ni7dWE6Vl13pprAKupwd+OlRKMZyGHsbpyG4ZmfxiOCD8IzLpfc2k
zFv+JyIsq00fVg1ACz46vYrdnyJ0G+aD9y6pdMqsgMwiDPOHdIwvE1uhRVN9keac
DZKYFUZcLyG8ts5iZYzsIWnry2SsAk0gkuHZgpeP24CpQmyaPHPAAOqz33B7xBn7
xD2WGY6x4zvj0kqpKCHz9krb41mshk42I0m7R7shlXqY/yQYaND1FLQ87tv7NaK1
exDb0lE45XyUZgPx21gA3MA5fuFY/st2nf8L49496wER9Np5KKZzKyBO7JK/Dc3X
iDFXbMpTUYtF5TLMrgIiBkCjRPByo9mnQPiJmpdPgGNhcpvYZpIdXsFUR0dgtW7A
vGV+oadnzVXb5wdyUX6+JjuxHR1qqWi89vVfpCkEXpvQ0UP/QGmJKrb0UpyeCiSt
7F+KIs0xZHiBTa2tKG2RuP9zZmv7UiccTRL5gzBWdEgfVwlmfRfCsQWa+XWSHka2
6SUrQlGSyrmMth26IrM5Np4SDcEQIrmdZQuK23qNfei3IyXGhFZgYrAkbu5vJ4/e
4bOAqPD9TacQwlrNaqwbWf1c8M10skcXOjL3nlJctxk0gTzfToPtSMGnTh+2PU+Y
D4ECERra1bz6S1JH/uIL6LId5BE9wN7OeFBLTz2Bk3UfLoJUv80hnHjuLNXhtZCk
OGMW6/XzQjAbZL5EvtnZbOU1j6TOnwntRG1M1OoYUm8B5CjMJ1432XvYfXaR2HT+
w0CPtIJEwvWbHTeq0y9SFWQCNwUBJxegJX21zNfo2ndWYsjMlek2msrWr9fb4R4Y
X2SyoovFS+E+AtqG09gr78dDyBSZOjCJDtpF3ZGuC9+trePW3ItvktTzbYMAWk9J
CNm0RPNwYQiZ/UvOW7NKuge+ZgAt9we25kv76166bQ9q0VxtLYrGQ2WoZjmaJUVd
b4VDXNFeH7RPLJnt8+rLsgWmbilhUz7M9HpO0GHOSqhC+JLQhQXGrudb14Wc6CRk
93i4JaPDUHG8024tGqXMGyKyQkm2oGo2FW+iJ94l8t6ILFDoJfXv+h5IsmUvA3fm
1gloGuaXemy6XVQHGgm8ppPSygP28kaKf3/sxhFtMuHnlwiLcvpBrFRgFD4kXq/L
TV2CLYTTG8RGQVp7Ca/K8FeIQykCqYSZndYwmCLPxnTuGvmVanH4k9E1pJ6qxAZG
CE7L7pgix8pogiULiL84UBSG35yMmzy6wrWvhXjxieApBxHbGRgLzzR8jovl/rz+
ciJqBkN8FZGxSNtBmXTkfNqpEyxS6lt433/45KzL/8mrxXkSX+pXL3d3syjOUluW
4G6HAwBtm+y47TitBS1MJxvOWIbaW/uTYqJJzveH1/x0vGn+Qd7BCllmbi8w0We0
9eyJhJEKuK5/BkDhXPOD5pkOVlEcjphObOwFxDzr6spXl8T9qU9kGrG/tdtbiS7F
4EWgNXyRskiX9/9swPResx4InmCz4t0Qd6G7W7D/RWZj9SZDO7iL8u6xmXi/13SF
EaKIdzSwA4bp4dHfrPQWCC/o1zXoiQnzm9GphlMcV66cvZmgSuCW44t66G/1bR1b
ZofiEGNQ7aJ2QWKZNbRCWnu6UpFAyQvF56jPSa1zCzDCJlZ/0Cxvbno49pZydDlw
veOa57aB3/iH5FRBJLVIx7wmdc1x15jFGgAi+YPnK81gnfuNNrGPQ9YHnVRpafBZ
3qKr03q0bSEEg9mkpdI3Dj/4Y2uB36PjRoi2rzbbj/kgskHwCA4UpAmX1LCXmGNK
cvxuVTMYecwsDAyyjTrB6TDOBo3LbhuyLIdqD5IEK88rPb2WTIUam/fOyjPDPGzb
ipsAApv4BkpF9sxp6mwWjA1stFGQDyhglyoAs2pvKW+qBvXvjNWqBqUvFjNpByam
83i2IiMCZhM4Dcfk96LFqWwYOAnTk7Jz1Q77uEeLzT+9HQ2a1jh7YyTWHYs1X64X
iYpKfQYnv0u7vHUbjMZUKKd5h8kO9+Q+khdQsgA/i7A74wS1+eUCwldY5kF0tbdM
/QyeVkXMd/MICn/HDIMh99T2aX9804D5PzYC45OLL4QlN/4dMxnL2MHd0NPB7Coo
P+1Virk9Oeu9picQjAQLKn/vwWG099K0f+wkDHWzWujrRPyhDXSyjWjLv/WmnWQv
R8te1YfXTVmuRUfihmAFxUlZyJxtL6Q8CwC1y9+FgIKjibBdhcaDTKquqXFO6Vev
xRkv2lFBvOGyhamixj5As/hwT91zJWQD2FF/wVumzO/ZrliVldVZeTUH5fIK3Q1o
YdNlcLfrFMYbO/khdxjaxnAk9w4kP55OI/gMGUDsz2xxJdHWDEw7cuw5ct+eJD9h
OjRi3uqWnLFnheRaPiUJGorAiFD16vSry2UbvYm5wH6C6HBH6vMGTpvS3Y3WRiCw
3P2D9GhY+n6fgzjUJZbvhdouP/UOBAvGdfNEZ/ScwTI8cFJ0pijUM7s1LELh1Dbh
nJ4AmNeEevqHlz6ZN7V8cVKr2i7/0G03gc6ft3OnNlikRiQchTQfU4yZ+kkJNLGy
kIbev+MKLm2olky3wo4fGJiPLtdpJXoqkU1k6IUz7mm4+s9P/8KVSnRTVA7gnQyd
FKmsJbOndH7stY8QiLp7gZwTWqhI71gSHlNffVZ/HlRCIcVZmm99yd+wspAoBmNq
+Q3Lxd6q+gnjtwkroo8vFsd7ti6bE7SCrtMqbF0nCFKgY/TQuxjR87hPxNNLyHQw
zrqSdA1E8xoH+wm4aiM1rg==
`protect END_PROTECTED
