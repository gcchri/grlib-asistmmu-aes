`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
365Vn8gM1iRO/OwgwFKNX1GwYxQzsDe7Houw73p4riHxkt0+lVVKd0ebuxW9bmmW
A//0e13l0TmYMnfiXGak9f230KYSlJ7J4LQiwxvS15/foNZQ8aXglZA9ctuthxvv
4xrH27nQ1E45lexsum5R9A1Rygq3XVH1d4oVtNZsc4Qzanq1euQwJesvs3hjWkt6
D8hHGCycAzO5BfHQqwG8gRL2viu8mUxyDrpQ/cd7JD31uG9klizv/UtipjcFJ4gW
qz5Pa3ECOsr3McdUkTwgaSYrigOiyekccPaYIloe8TB99fqkckW8piUE6h7Xen1u
fqPChEzFGZ7MFFXQ7l0jD1iEes38A3OJqLdumDhi4eF3p/cuJnzx4I97D4z4oF+i
tmdPK3iJ/Ii20NYc0FnSgspP9H4P5mLAcnGlqJ2tnLdW4vAhjAP6yjKqv7kWRntn
WROg+impzdQR7iW38RvvgTsMr5p1NKwJJzDy1VrcXWPjO4ycLquR3fk0QK9F7wkT
ma+bzktLnhk6F8T+ERYZRzvvIOpR8oas/RHZn9n9wcfIfU1S8KEXYDG1Xc4t1n9x
dluZwDlKBMlu7U/vmZsWWVNIHM5BG5dDuJJoOo0nntgFzQaNSMTTCROId12bXpdc
clUnmy7A3OKNNS7jacZx2sTE0N0ZPKJz1eTk24YwyVI=
`protect END_PROTECTED
