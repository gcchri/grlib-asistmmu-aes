`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZYRn6hEWmlYG0F1EtFb1+d5YTC0nBX8x3Kiqi5Ho3DKR6MPnbcpj63crLq1q2dk0
4LpREPHJPrv9DJUjYt2jQNoqdgkQ7RPN4xOMVxuyZJ/SXTj5F9tgWvyIB/08cW4q
sMrtLVceSoSSpodkdXJy12Q9b1At8tYNYn9IopmWfPGIKzelH62U1tWRBmsSMLJg
51VzHOCjAIq9EUh3O4n4QeReC+YJxKsPW0u26KqLYSjaGML0LANSpmKGEMNqMvw+
67hEHw3hrZWeI2MPeTgRnPZaq++6I/fRKHSdc+b2Rv0hwns0AikFNDpawSi3IOWH
Y2VZRSAnP+3e5Xrol/SQTO3mQfyX8M8/W7aVIRRAIctqI0lugRlQWcNzcgkCrZRp
WOpB5hV/LzI4dEhpbxX0BUfHrW8e44EIK2lviQB2Bvz3rlriijx5XMZWdPA0UrMQ
1sWSMP2iJnWZKhBk/NISPXJ83WClx6OuWNETFj8jIYGyqgYQlZ25Ig0phx0rTByk
Qfpe7lzyVpwBxgWhaQe/AXrsLdQxXhqvyui3bY4vqhfEk1tL7jZPq8Yx5hDFBZUS
52k97po/+Tmuc8poyNmK+g/CBCVIDSWXoFSB7gQxBsK/2jqOtbSBUw3WyzatT+1n
M5+/4qKKpTkSCSX1zQiTtSDg85E+GFWCFHbc2FCU8D1FlQLJik3YwZ2TTseuGxhN
kj/tkX9E4o4+ghoX2JhZjo8Fh281eq6nnu4m6lv0pML1d6mkh90vSMbstcTJfzlZ
3Ie3fAbqGJYvhJUbbWGhR25gfJfHIToKueI0SAeEuGHja9tHhN7OD3iHU++euKLw
fP1joXvgMUzXyDb5wSzo1jpJG/di814SXsXZisafv0HBFyQmnfund/UXg+IZpbkV
48EY5t6ex5LWTmCF10wRfdccd3yJ8EkUHDkwZq5b9BCVcfBKz6h4INj4NiS6Ldjf
m5srNo7v+wapuvwX5RNZGdElJbYjg05GM6RxV+rsmqSfhn60xJoNdqFHdcRZ/big
gXOdRIzwXNLisO3Mg/DU7g==
`protect END_PROTECTED
