`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AjAq8PFLJ9y3QuMoA/zQZwH1frtfai4VSuw+p0jvrvN1TSHpkFF7HcvmUBDH91AL
C5sjiz4CHasRznoXY0mSUklfNyqHL6ISdAEuHaeHSbK/7tRpF9xn6UZp2LV0k6sS
RcY8aXi8XsejfXOIzr7y6bqRVjZzG5du+ngaj0gNwVNhpGtwfHVo3UKP9Vw1tzVg
r1TJct28HU3YneyaH9QuPsOWwsvkpW19H13ByNRtCxv9ntZO5qoTvrCLGfVOQ3lS
vHIayHnDUcDOk3tV0rm4NnlezwWMOBsm33GuZeSE5T+gLouTe6ST02Vm7aWB/2OL
NaxJI6tnb8Ctjzue70pdh3HpItRD6wGTaaM+jyFvLck0raMIdF69NnZcCmegvIWn
5t9qOi7ITWVYIx+WAUuZe3lXG8d3zbnN8uP+1JfBue1pcq/lSSxWsyKDJ8jcC95W
KPALTsJmNNnYJlrFcWiXiX/K414IQ6+7aLCpCcr4gUs=
`protect END_PROTECTED
