`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xMGqEC9rMvpQKh4zxkfBDawFQbCpogIgyLyDxdceFtq1A/uW+l7yysbt5fxS8E0q
JjDZjp7Bp18WkdyBDlgyRCpVMhlMD+S+W8yV7yRkhVw7xSgu+qO9pB0dN40FYP6h
MW5ZRGFFchUbhxbxwmBuMi6tFepgkoMCQHZbcYKGgMbfI4r2gzxKKTwIR9XvdaEr
7WK6J4XC0aUY7RLj3aWjzDPzSn516T5GuWPG7RqR9IW8PN4oS1TGVbYBssGGNwSx
QubhVGl2wRMsiW6fLZQD1fYvX9QYb6W0J9Ne/JshmBLttHt1QEpWV/dPQgGv+5/A
ZsKkexYzUWZgwzpCdq1iTY/YInyRMNtdnhL+cj0G6cpgT2w2bnfHYJMYki4dvahL
`protect END_PROTECTED
