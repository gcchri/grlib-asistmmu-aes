`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HklPGnuDq7ViwSfteI2UPuFeq+6CpM75JgiqbQaz87nwKBH5rXl1QQhXbgxrdg+I
EL6668K/DmZ7o6IqhuPlPC/2CTw76ykrLnt5oMgXJv3q7ligLaoe3aZgkewJP71u
4EXCQaGC2cY9GLsAYfe+pxHHG3y5+c4WrrKo1grz6tupVCmWCZcov1u8ReANUMnl
A1laKFUT7Yu/n8wOl7nt811QH9uHX5lfcDA4dfjuV5+b66O3JmOadrTlLKv+Dysd
`protect END_PROTECTED
