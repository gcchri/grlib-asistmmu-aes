`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dCPBFaItfzvICkZhLsbhYPt6UDDwwj477UM/kvzBS7hrTIx0ceb5vQJ7Ec2y4eFR
FyLWoXz3WX6AXfp8ygM7ebSDAGEeNvUCsusf7PG1SBQmaeEVpOuuiEnqpzsuUFwd
3xeFj452SfwEhfkfyQpNcLsbiqfv5SW/EcUaDP84BNFY4JABw4spK+KlxzJQgbvv
or74crb2YgFaO6UxvyjNYICykJ+ke2OV0QxLLU2EN5Ki0NviYWdhT9xaa0DY3vFf
D4DDDWzm5dRgVUbn1HTCTwFaHPhfyszfTRKdOwAaS5TW1MOY0/n1dMHzgvsdMfQz
i13pBXGisojPYkhEOP4hbBfvxrbWjPccau+RR8XG3r65X51bGhLAro8t1N7GEzuY
Adzri26NQapl//8WAV7MpayDqXc5Fr0KpdrnBrmlHGFkvqs/Ax2yxbtkcrSRsL60
rkz/79chT61IHEgrIYkKmXDfvk+aRUcEEpj0GBleR/MGPUatbLmIyaXkMHjFHZC1
ZQkz97CSbPG3dIsdDiyLFH+fHN7rnlPcsDF4fEXlWeOpusqkuT4jU7UlXdHOzK5t
WxV1kTxSt+kkafEbqhfjokUCa5H5ev/g6bRROOraxteVqIQEjE4Tn3Iq/DTdu1xP
jXYN5hZjzXDIz4piI6f66hQUIdVri+1RheB7R/I4/gQ=
`protect END_PROTECTED
