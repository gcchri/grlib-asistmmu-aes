`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wejLY53eWnDBHaCj4INWgrF4xkj5uqIq+trugLjd3pogSWXE+uKO6wgGJUJ1rLcz
d5ksrIixRSUFjyCaLXVzN6pEEkIcIZnrqjGq0LqcsZ4zuKEGInw8wOkVXvtgVwOA
xs4phzjMkwvhZm3xyrYu3Wi72EKnvO3NlBdDJaEFDOm2E2V5SelVAfF4PGUNq0Ao
odNpFbhaLSdTGbMlP5x75NgjmaS7b1LBh752NNrbMwa7YDlnXYpwzQO1oaJeS6Iw
8Xesny8pF1Ry90/mFF7+MtCr7/feEfLXR7v67TKj89Uyu5Fke6uAGytFbLGOUIEV
J34HvsbB0MvU+HJiHJF+GFY7cCoa3KQYgXoym98tZiSDwi6p0WSrNiwWB5SC/VDv
kA32HgttJC1lQ4i6P8P7hCdn9wuRIeGprScL4wfaLBkqsEiObp7tvVpLb/gAgFzJ
M1F/w7GLGzVbSBcQJ2NozaIAxGecJUos+PxpyHIT45w+CM5LZcEqNzpL/na3TcOg
ekRndDB/PP6vWqmZSp9ygp5RbOY4rTvP/mDHTm7/WpT6Xu+O/2AF70HAE2BH9Veu
Pipea37PBHLvSYcOuSZfXg==
`protect END_PROTECTED
