`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pKkvWQXKtushYMf4xbd8LoZ2Dbcrthu4NV/9yl+m6D1EQKTXGFRMM7MD7bcrglH4
TyzRZAbXkvDLYw2o0iNKkvZFUjAqhiKEaiRAPsbkH+D6iiop33O56ZLVYGKJPmCj
+dTu+qkEyK1Ew1P1/bmWWIp+nPTXuWvipZEANjnImTmcGjLmxF4ZaCKePqYkP2ET
HTvVZcIBf8bR7xjXtaBU2Nlh7mv4BRcF+VzTl8TGgJ4kqwQqaFFWnAB0+XZCnWzl
HK3yR7XLS/TlLRKxZwqMSNbxO8G4SCUDAEB3cEgeW1r5Adf1LK7uB6zNoqRXkcRE
3/dFJmfkZHxxUmQOt1c+jPlq/mzQtFOxGLpG7Rm7TaXrCeev6I9zkrvkVabeQiKA
QsRFqpiXuQkEeLD362WN/x/eB8UjfkpruTlWT+8InH1ZW2sgMkMIEdanMtVEKTLK
OtTdZ/HJ/D5brWuqz9CKcmP/WBQJpE+y4U6mA27DtFkIzNfmSdCmYrwrvWIF5ksV
+sq8CdWwakmEAGNyDwc+IMac8BtRRL1F3uC5yV8QIrKbn8fr896enShkorrC2x+H
jZi72mt+BNPAqJlTTSdhQhwAXUjTM8Zd17VYMKuWK0j+U9PuasBw+DikgdP45P+w
nqlxwix4LKaqi6WSmutYFn7Ad8uLyORJdjvDxkXi7H7fzhcgpm8jv4+Z9V0fIkzB
3+3sASsEtwfIi3llynLLECVaURjrD7ETktuJi/tCAdKqDWWsXaA1nCBWS/BZ3cse
ljuC+OwrJjPo2Tmx+6sAH/VIQYDQQhEIWiqgVKY6Wsu+wuRFvApVqTTpwsQDLYq8
L5cqqnHMGmqaRDFxGcIfHtQqnfi8DmXh0keCgTdnZ7ig6l//OuXbvWkwX+IYQhCL
X7H2YUXbcHYh1518pLFQoDTs9oIkToUFgMN0gaik0b1Sk6Vmm1GMYSnyLkVWjFQX
`protect END_PROTECTED
