`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OzsOHR34LDa7x9rqlFhOrEtCDfQc+cVXcTb86PjJ0RCMXjrwcExoL/3lOl33H+hR
xQT6CQL6R01t+fRxS2HOyYenFHA6diSbNmTAue939gKTWYpiXFD/8HgzICEOjL/y
IpmgAHEFanE3jg9DBj4FJ5paTbPeB1W7sDQql8LBZcGQPnXBBgwpyZAaL8wO7PAe
8xlSw8sRKeUdun16g24AN9+StZmXXNrkxRCGysIK58ptL+BupDEpm01twW0wJzeb
UrisVZMo/9eQiLbW00eFvVC8F8GumtQUeGKJAPhrDZBEigAa1F0XUWT0wZZyLJI5
1Hw30jg3v1LCrrtNVcd7Ja/RCvOsIXbVPUl9SLaK/axiayKJbr8nkg5QCDmKzu4u
iD1707ePHYB3/RFjKS68vR/C+sRaPDbTVG8RLuSPNS1zHn6Oo1vo72rvP/CpQczm
+C3phKmut89NcobQcfN4eiFxU78IAjlTDVMy0xf/tVQ=
`protect END_PROTECTED
