`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5vSj2B2z2qdf66nkDeUIpyvzr+ZqjPWn/jDccZKeXDyZKwbmAL/d4oW7kSi0XZF
PRU0cD8qlFpyyaNvNkrxPUaCM+PricbEjVM9FK5EWBFP1sMDkUGxgFVCJqCFqdZN
b/3yezPFsERRjUb8nXslKoGwdhYgztgs36y7Gw5UFuu390xF+SW9dHWadhuXxqpt
ww0ILL5hCxDoyoc6UgAE0A+gVrbKSHGKQhLemzvmDPVUKhIwFFzJ59CPiQNGGBwc
9AVhSP3PEYjXNOjSgGqvAR01Xm5jFzhYYQjm5Ib+27dE1diL4yHXIirB/FVJ26Ga
J34GdWDf++vzin+d2DNQCeRGuXJay7eWQGwqNNlLW82pSJdZdixSyNW3k5hYWrFd
ZTw+M0cSy+2jtBZVr/sfDkaf8pADlKJNodZs7wddu71xQ+8zzI25gFNF7GUzPQhY
CHFEuoyxKzU3MDG+LMi1lpac+iqTJn0K4znupUBrASzMZ/rbmy9TIRunJgDWhU47
`protect END_PROTECTED
