`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jg34C7NcIteN9n9t4WDE2FBqcPPuhv2wEINjhzIXTNt+QE5oIaB+xhOvvlKL2yKW
d1rnLL0UwIqKKrW4Dx86YBUDHsgSUaRW7k/OAKDNGnZ8SVfgM3aflsZwctcr2nDR
hzzaIbg7KnwSwlhEhZxkPCfGLlP79yWKS6Ni09GIBzeExmAY0Sqot5UtVXLafppb
N0HAl1LvIEj0E5QuI6NwH3uuoAqWhn2MBuJBL7RiVflba2p/v92QTzoTH2YUVNuw
`protect END_PROTECTED
