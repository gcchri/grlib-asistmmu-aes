`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIZwMmy/A/dibe3/uJMpZInbKtdeFJqoMKuWInbOVaAtsGbQkOJcO2/hRKjr6yIX
gk0r8aCXq6u0DHnYN66IE1jgTwM9p3KWa4EGpNNlRdYMyEr3JDvhbJeyC4wakkxg
ltRZEZ1SBJ+hDzvR2uHFKc2he1PU2bDAlnn/bV5eP//gLUpbZjJmMyixdjoh5m2i
xThevny6Zfr2vwj7S8zyZy/vs3FWKvshcT8UEC8vJZU+vGN3L938sVWCjXTaLj6K
NYjUPtmUHYVnOXUKou4AICwMksLKAXIC0N2bG57/QcEZRZRpSRCPrCPi/jnNTXVH
wuRhGva7p0jdMfaOcDZpzXnAgJ9zqPB54Yl5zdyaCWAfqkWKW5cYUTNYtKNsbgdk
w+/uKdHOWrf3xUYOr6GxGHgJnsrqDtbXcxvbKf6Jwn2DGT8mqzgZzMvuCU906yqH
c7U8xBo+0s2D+nuYm9m3V7xIevzJ11mdpJebBevbyetVgzU0YTv2h82XVyCcbt1h
XcqKV/NTGnCG5BZ3OQtSPcrfyh/JGyqUncDDGlRKd+/P5eoEgG0Sm3s6V4un74/V
DpGP4cfdASnH4vI+q6n09fh93boKIFv9KNA90iPpNE+rsBJ3DNw5VMyNnhhrP+lk
C7zQB6eclg3lUtdYFTPcpT4+ccQSW2v3z3VYyuAsAG3B8TskD5iBtmiAMRiGFaj6
`protect END_PROTECTED
