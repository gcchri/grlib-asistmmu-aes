`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MMxFVu6YK0lpjIvYSaYji5Jp/fzHNAUz2ZNGuW1XU0y5a8dbF84QdWck0s+xumHQ
0F0CDLlI++VnZ6q8KINUzuDJVwijUJ80o8xRRmrqXrOfDkwykoB6upUzny5yJHvJ
CtFitzn8eCsF1OQ8QKWZWH6ojijmYM8rVCGDA7taQc4R6eFClr3sYOxIiC4GLytf
rQDkpNu9M2PAaryV+fZEbREdTTkvJCrmSJgdimGpm6SYMPsu8+l0WZd+wPB60gU8
n9zNP8MqNzwmKR2g38nqpnMh8GUueY7z5m5gqOgPqgNdJPBcO1XoxzcmtGTeg8Pb
W+QP4+8Dy8t1hU+MZmqnRKVVQI42DqndZLHlJ831c7XP8wGRcTafekDLdnNPF6hn
KaNT7XnI1c0W8Ly1AL5mXlDRLey5XLGtmexO8wEAd9iU74KYCBQD49x/ajjUoa8S
3jvrxawH6M5tFKhSdEkkkRleC5NYmNBrHPc0IDh0FKGVV2VFH8n5/IGWQRONlZ94
RN1CABptf1qQdHj26NemfgSGOY4jbU//oSWfDx4lrdZL5CwHAnwdSuyRJtrg0eWq
18Uhb+SnWAeSEy9l72S5CQ/tXj1qYIy3zCFcauYJF0C2p7PylGzVZYkTEUwyHrr3
WC1mnmP9kiTvSHZpZI+hKAKvCOE4KutbYTdYxDQVmXxKi9po3Lni7r/UedHyYtt1
KWO9y4YhpgQzggdXRpwXXrkjokvyNOuaKgsDrkOl5X5J2UEQidQjJxXdBckgH2xh
QzJ8zGlsBZO6qx7hRozH64fPdKpuqhM7v7gqQADew/PBPFwQHZCynByBMBNpsyDd
Pyi6jxxafGiEY2UmaptdijFljzYXanaLDX+PyYOlm/MsP8SN/TkU69D8j78Sm4kT
nu9V+2UL/8HEzErLzSsekTDx9E2wkHrqURjlGoUCxWHNmQd/ReOsNgY3+VNr5SZf
nM38PGcshbG9zPRk9dB/4vwD7/ijniu/ZXRbXgYrWnCw0oclc+BM+5ZYSLs+mpbr
+AS5IECBx40ieHtglqycbK0ZNaeJBmRT3xOkIp5SYPhFUfEuxdj96Xo/ohzCegJU
yKkMjzBtEi56cPo0M4gt649SH/Q1zYwv9tLGDTSTVUOU4gJalC0l5Bk821xn8fxW
jd7ftkZberQnXQmbrdTG83i/N8R28I+rjsiIGjqJhuOZpO3+NeRhm5ENl4MVWa7C
KBUKQepkvaamHoHEsOsELIY+pJxDL/1incC5n2IooNcYUh/CJcER9zNLcZootyjC
9Gqu1oGlRpSEY/ecxt4YtdIyTj8XOG4/EMn08/RjIhjbSy38HY+4yCkQJy9NQ2DK
U2/fkPxYhUvU3vKeujypk+IQKJxHcHGMacZKZPsmsVGGzGkR4e2cyZlJvRGgtmD1
DaHlPW6TOTABEGLOy7GJf3seWfbpwdnv87PIn4gCu18mzAnsXwBPwuQ1Sby1S7Ln
ZF9PUwKSPMMyFVFxBDUnc7I9MnbfSCZnVH7Rt1jLvEPWmrYZy+667E2k0yRM+EpK
Uwu7IlUZcII0IgqtEK9SYCa+DWIzVnUZU5K3BMGW6CtfL/+VUrCgAt2NjuQ05Efl
IEmjpxCMW96/zGWgBY9yjaTlX2Cp9DTWZaQPVbmY3UoRzd6DNcMxHA/tZ4bx8f3E
/diNPlpRo1rMx1dbgzFvBNnXwoa3MTGk7sWLuvJ0Gbf63U61pq1g3XnmQ3SKrPfz
+OSnZZpdfrdjIgFc6pEkIf+IhqHAUCmVEmYEOn65DqngGm71asopQRfh2z2qiOFT
PN/DZhM8GEyFWIOEQByuUe8vW2kreVNdsnXehiAXlnqtNcyUuZB/4KhXJoR04SCF
J4kHIA+DobxAhaqStiLplyFASlot5BQxyuyayEJ1r3LZaHceflTvOy9uRLH8AsQA
A5jLU/p1EJCEpjAW0Di73TccWxAv/37SyroBmbtu8pIWfr8XDYfLpDzaDAZvGu3u
3dUo9DJiSDlMAdY3zJXT81Mwm+bnS6jxRnv5zRkUyj43fxXqh38KTj+nJ6Q0af5O
LfyYpsDCxXah9ZTmJpYNfuwGXa7dItsNSfdAhC7vnfOIlE2Sz6CpvDnboulUb7PX
HKvfBRsHk4I57xfU2MR1JO/AV91Bt6Gdq5ql9tG8VLGR7qp/mnE1Y6is2Z5kDrgc
NAXo5O8JH/CSFLkacra2I4JipVteFlQajV0UUA0DSv+RVNVq+Og9PeCMzFyfwYmp
Cck3u/XqmQQ2nf05SmsRLbor2RlqJn9NuGKq7sXkMHSUD3MmZXLWbCdq8iSaLrkn
1gmSu9sA3EDKPuf6WUkpHkMY9pSz0UI7bUtF3RUU12K7dHvBo52mIaPuVLGVqXnz
/fWHHHtfPvJ3mj6eBmhPumtIMAm/zLuJ/ieO79RdGWU70MTI6q7BJ+4W9Aqr0esO
Bl7G3jsRq/JKENWgpIrYnOTM9t6DfH/1ANHQyCEqyKF/PRhpKVuDfbwvEDK7ZPcc
eqTReO9a+zio9Bt6SjC/0rPgSeh5K+oGr+V0XjUGDd8MGxC1uUWUUH95BC+lAjFr
FIfOCMjmxeAKJuSS1g95otIaoyc0mdgZFj5xEfzoblmDeinxMBirAah5EqJrdjNM
/9IBm6x4lh+KzYere2CxTienywH7HcN8kWFNfDx72HLJn9GRQHEs4HWgzPk66QWp
4T/RYRz2Lr88qQpMbvb5fZfCTjFV3rKMHracaDH9E0Q63zdD9qPQbcfWjnkFCTPi
W8iONX5dJhzdYZoe+14KW/b1mUmU6E7KyCVlFEolb/b4hzGwrarueKhKSWpzN2Wk
xOPK6vd+B6hQ24k9Pc9LHPGmlNqsaopXsMDP0lM4+2RWfMvgnUW3vx5C6euyWQlC
yKZIK1ZHxxJReY6QbWelfzED7dX/Si/uIdl+uyf5YZGeA9Xku1R6P36L+d71porZ
khuXMmnjhHghuWbcOE+kDIkppI+Dv5YrgY3b96ygHwiOmNn8+g6PA/DmBa5RcXpA
EkgDaTNC8beEjtwrZCrRr9zyVV1kRIFKnkEjan6kGhzi9gvGGc/K/zVybEHYFBLQ
HzpWEXpJ/HySf57aOi98+3CdCfPwBdE9hCk1YPvUXMY=
`protect END_PROTECTED
