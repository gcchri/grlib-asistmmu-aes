`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KakE++KCyCR7CUKLTlPWl6f0MTs7GkRUj/uqvJLrtf29v8FpuLSGtXQusozEV72+
Zo5LHh9l0zfmofTzGFxmril6gCYDYNhB5/okTicgSacM+2s6HvA3ZT5Mt9SMkZY4
b/XNY4MCJ+rS9u7ByTT9AQ1YHXQ2LKpkcz6tGexWb6E9LnMEcUvrsyekXYZB/pEn
5O162+4voPHm9D6i4vWXi7iKmEMkU3JMX9mbK8bI5MkPpxJoACAjvJ9mx0Wya0bL
wKjxwvlDQTzO/nyd32nMi93A/Y/kxsdE/F9J7SUAsdSMguP4EuDmCEBIht4xiEoT
TGF8SUJmRzmxJZMVnt0C9CJ0ucANsNGefFBpCAauMfIRURBr9VhVWVWNfC2tZZNw
`protect END_PROTECTED
