`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gz8MN5/bv4DhbZxti970Fo97LWPzjW8lGPwZ0K0OpEGGJ/lDh2vHu/TyQK2CX3hT
MdMJ5uMfJuxnE62seWDyfgmmyLVZ6CgzsarE51U7gUges24yBLooz5rXjDEFY6UB
Kr1FXiM/DxGkWglUssjaHEFshz2qHo5TGNC8TLQRqMYBe8V3tcyM5ZmbCSEBzLME
f95iU5A4WL4u6YNgiLGJFiAIf9x7esA5nI2SjLvAvZq5H/tKoYpyn1A2H8Gzz3f0
sxKIw/p3hU/QyTCfNtGK4FV+fX0qfZeUa1KVRg2pLRzl8lFZTxVkmjqOw/KfMX9a
EQ6MCxD3JrRRA2yXisaAR+SXv8E0vmWENhqZrwb2ChpgpONbxaBgqWIMX2YOh9Cq
p2cCllZLWZG42NkzjVJskdO2snMpKHO4SSTz0QDH0dm4qI9qu8RG0/cqJPTAUm0A
X/OSDsK9nFacBtt/xrESTorzoijYIzAu3Nho5ngXBuDYTeMyI5qp1B8QAHXCLzgM
JCrjLH1hsBdNg9C0bQNSUjuoWtMaPgTm6E1eMSdVmuaU5iSEk/nwcdp7x0Yo3SDk
qR9XtR8VrJr0eVaLZ7YKOUh1Ea0rJPVCrQdKRK0ms7gcM8xAh7UzvUCVsBqAYEuY
/tczJh2wz1t+fqSh1kRAsZ+S8xi3Y933LAL607matejzINymaBCXTVIfamRTEJqH
sWfrU0xT8MLe7miTy6lO6KbLDQTpRfTeJOrBO7SGsr1H0gU4NMkX6ju5eXgIilmD
tonVa/CSBbOp5X9EcGEr71dNWMVx6GHjXsMfO2FOM7+iqN06ttH8leuEb/VctSZr
0V69mHPpE0kTKeNkRnObacL0yMuzZC0fmwVgdDoYge0cqFl8GMVyhaSu+b6XMJr6
YBi/K37O0tlZ2dVYLy1tImrP/BS6G4nONMvGDxyHnEG7WH9UiFx7baMKcusgog/h
5T4dfSvpakdAvv5XpsATtAcWo5+fWKl9M9SJoUH5obgV4oAziJp4BR4xNnZtq90U
AiAbiJbx+5I2s3GgXmcDYnPKwCY/BzW+thnmTfwJ3kD5bgmWrcO6JG7ZpmQVIGWK
mUiGeh5QldA5hwVscfSXRmVCbwSEriFizoEEAp6d799o5hJ5LoBFcO8FZ1iSbP32
ymAmXc5e4qDXfigZBryy2FtzcC94lNIb8GFTc7BzhU54fFTNqa002CUVUd8ZDhae
apGwGSRr/BZezFF4AKSbtq5mR9zD8CDgePAuDZ79wWZu1/1YSMFDIiyB6DTNDzFk
5jwixFFFF3pUpSsNJHqfJzBNJck0e50WD2gnj/SdbbVCT+VxV/HJPJDFdIksSIzX
sGp2iRcNOshteMYOilWT4XVIgdxCSFjB7Y37xyx+jq/36vvRryz9+r1BuhwgpaDv
FOqqHxET2jkjTddl3p5+uUqM+N+3ItmUB2hq9Qaa/4kKZegqcnj04Agt6thuIDou
l2PoCVQ4iXDdHqhanioA0jAUq4rtTYRFPK1+XtTwbA3Pc4WdrXZt4N1v7Gxlc8+t
Bj2gtbtpTtZc5E9XqMFfXp0sLM7O6CgtGHyqrPNmfOykQdLZKhlqqAY202LWFnz4
f0qMYyLj+GfbqnG0BNt7Bcb9X1JEVqoRltfP7Q7tIKse7nrVz+aNxvOID0wf8bXh
UwIJ+Crh18HQ4RcDla8S1rdB9dpDGkVHfUC6nkkOEBU3aWblL3E7qRo46P6K/NH4
PSISLXEinmXfkjZZasnrmmdlwsor++7H9ph0foESzwr0VnQVXPvfj5x5t8ZZ4sel
l8Jqq51iUiUYybAWKqOcgZTLojHQt5jBcTyNOohNvMVIfIqGsZeJZHBxG+xwIU5W
QYK2JeSQmIgwEyyMORMlkqODwDvLpRhKkv6AGtdEKkrQ82zznn/6b6Lx7p5vpp2s
LIsusdno8hEEhvMmjnXyLt21JtIElxPJmI3mdJiCNRamNlWJCrChsey2z88GriGm
rseQjY8Uel4ktBF9pPHzmabJDIN+xYfdTqSMKi9/J6/4aatcAX5cTzSRk/E67qAT
eo+XW9Kcn5ugxesH3FceTzsnFfYdiJwyyiBiOY5STZaBCSL3n/oyyCYWNrs2MFCx
6wxrcE8qu7pVhvgSmbrsnchGdefsXnLtne1ILs/eDMi5Gb+a4MT/LI/yl6Xfjq2K
c+9ik4wDrgxphrM0nkI4oY5qnJmMosDa+dLX2HuDhmV0pssLANktf6eD/UBNc/7N
WC6GwFBkXkKp254kHlgFp2nOC82u1Wt02tLve8/Z3cEms4rWSpXxj88uB9qRnS4/
eD2UvtIp5GGm65zvZudOV2iNK+CGhMBU/AdnQoPPGpiPHDPfvTL8lMaaRw8Pc9S/
36YlHYyvJXfyKa783jXNHWfB71DpS31ryZ3jRkqOZ881NQXV1tHQmX0mbINH3Er7
z2GpFcOjTCZNfZfQeumHM/cCulT2EJOiDx5RPo8dak3wj0NvAbXy+Ww0GnfuNmht
6OxLgHntgFSBQOcBjdyU4L8AKJjOdKFj0Yjj2BucSC16BO2Vln65rXioeqWpTDBP
NrfD3AQojcS0VA4XJGUHiAMjhw/ZS5J0DzlWEhgU5GNFDga4wPs/I08PSaTWX953
cef/ib6Cf0fFJeTVABiKuXU3bLEdQ4RXKrsv5CRoDqSgqexZn2NmfvxNMnllZfWp
DoMgOGRoZ/8NEisKvBrZwxO6V2YsSVc6K4Ur3eL4AwTRcig8brzgLr+MIoeomnOJ
EAAFAcQPPOCln5LbF8guslYD6lYxLU+n/63trlsB3Darc6MJxAhBilvBhnCjmGG5
EkV9QYDDVjhWr7L904FzKTwI4aWLdwoUAmPsxc+f5mjGTvr+wtswj5iNKxzmJU1p
aW2Z8tPUxe1TjGE5weeDx48mVRNJfbOP6QHvdZWPkhE+y7jDJ0GBsMeUQRAG6nUI
S90Ou5YrO5PwJDdJLeEAhA2N/Kag5JbsQvOBQYEAB822AXWoNqn3eh9xULjD7MMU
1ErzbI8PeCnJEqRxNTzjOROCxBZlfj6C3wxp9lwByjzHwcM+IxAufs9PaWoel94V
RVqdTAnb9rmDAF7gSVrEQmPDMUDSfQjOkOmijEPPij6T3LA3ME1iVsvSlLL50MdT
S7LHzuhc46SkLoxlHBtNfiY0frQIeV0blQJLmMbeMS0s4/DcMhqNhWjRVAJRI7G8
gqFGBid8poJ3X6LnkD3BMgZ/l4JfOhLGvNZrHKL1mc6XwVdKrvuCawIypVUJIGob
XQcFCr8P8t9N4ERVNZhWMXS+qJakGBee6dZylTbzAHvLRcB9roMcnTvrPf7Cif22
++Pkq1URZhpIwgErbEkGSbH0wZjcSbJmBTeaMMbgCHjNmwJvwm1LI3TYjvi2ElwY
9bbGGeprNWdO00x5kEqVA+6Zc1kXauRZAa4/+8Wg1IBVKbB8fCGaNnEWWr3NpN3s
XOFBUUww07qjfrGpyUJdfBQVLeslO5qxSJh4H3rcjv5WXjjg1IfJPjEeuYtqRmoN
OB3DJAQNWCXuTlhFA38E7Ygom+NipWfqCsEeORRaiIri0whFq2939/nBj6U5nXpr
+WZVSOWOjgZWLyLtOyfAMs0iReq1km1vWWagaFHGfJPmGrOSxY3e74RHOlnycQee
Gcrzv4qJjZlgslQmtwC4JbVLVa2s9ZhiXhs0DCHqx+sZID5djx99hTMLNwem2Qdb
49mI6YsgJi3Ej3nCnMPANbyZ3LZYhjxXNS4lN1nIJlMQLpdPQIXyDp4/SM9hPTGb
GhKVgnCAQDvY1RYTmmXQ8ArVZa7OtWYlGnFt+MKSPsjZRBHbqg0ew+eMpn3+himN
5iSn7IlnJ+/mY4InuiJCqfh0Ffml+r1JUblkTxcKpLpPnlu+3LMEgjyyc+XDN9T7
5U6CuLvv/WK8eHLhMYFv24Gyr40wstwxfffsQkwYpub1VEo/kccVxZht+FgiuBj2
ESJQKGTjT5/ykG44w7IR5j9vFiSVTvFRCSDK+ENmzbi8G9yGi1YBTLPOgchQfYz6
3zZNOtQO/RpvuLMFPBZ9NCM/pCA+igaRzoKMpxhDganRnZlY76/SYelffWPRR/Wi
PDAlVKYt5PdB5RMhcHsMPsviCXc3qz7TVQ7x7BSgBysdsEbAXXvZvrCZxXePLchT
XeAXPqxlUwfKZXvIMVjszdk8PHky94D/B7C6yFQ4K45FBjp193b3LW3DQgZ+EbH0
MhAkNvav7SbxMY7sqYBp7/LY2gwWHehZuIQLtF1uUcT3ZZL1qHkUMHFOBVfiCIu1
uTivzRk9TiAZD9BWzWB6R+Jc47tMnU1S+GP1GR6FVnct5fze4L8yWhFQtykG7r/K
kdJqmYu5BJ2adaPk/Jq68dMiiuQSfqXovYI4rO4SnY3RNw9Iw4Tca1QLJZKfxbIG
vHxzxGt0yMUY+JFRn4mDWL/b0AjMrwCnTEF7OTQsEANuy9fGrMT7KiOr5tXVQlSu
/1Yw9cw5ZZf9VObVmkef1YJqQODoxn3jjNGZz5sDUK1MsGbmOfW7VBqIOXPjS7LI
rfARyCW6ZQRXvn6+4axsQND8XquQLwN6cF3RXcOYpsAFe0WyIlyrLmuIFQWMKAk0
9l+dbjPrUuo0/1AzIGj1elyNigW0rF8jh3z3Y2oXa0fBOXZ42G+OwZ6JdPEShPZR
GRZOteFU6EM22qEBvYLAh69rGXlxZq5duyilHAh5rs1LUZYuc5LcD7ujcXc5cjGZ
CwbwQkB9GgzbV8t4lJPpVQFbTxrOnXAyUGnFeEKX4BrkflluwFfJ9aj7SVbLQbG6
5GtNQ1+FE17L1s3mZ6VOAz2TlkBLv5JqhRCnY/RUPS3j270v8k9HRMH68up1LvzQ
eQ3IqwKRSifaLZum0d9/9Qugy0H2REvirwGTdBeNrhv0IFNLC/WaRJ6IQQSFVyEV
IWJdhX33j/1816GQtZ5yUKow0AFBHBklvfbma8mv7PcKHFygtqEVTCUFMXXFn7/l
ukjKV/6LGo9IYdedVzgkwQcrPgrHRAOgN0QE3cnGr5uqWplzFwqQgsKGHNPOBsjV
9gmY1PTR8tdCm87BPzQR7qyRGodJ9r7NlcyaYlKwepMDNypiRKnotzPMvWnLn80M
JCSEzwXXSIDSDt/W6SwLad+35zJiniY3ekYLeIXWgTbTeAgbZ1om7qQV0aN45P42
qLezJADc4J2+UfIzvSMrO5FjnqHBr0KqNbWrz8ooKHQMhFtlQRwEJ7n73B046T/P
N3hev8IEMQUeszBkTmjPlguyVpDWKq3AXzK/nu8unP8uYfTXfOmsLsHVqt+8Gj4F
4ntTMLJXJvHED6vTP0MG0/gmemFlls6Pushr+Wyi2ZJxTkmMy/lWRUI4aBylEx60
SWtgpN2hPIGzQtKUTzfpTLf5PlX+v7+cPhdb2lle0H4qAQ4FuUFfVttvPQr7elQl
Z+vw6XOFTVTkRgGvgp2X1bZF/krvONCvsIBQr6EWwG4=
`protect END_PROTECTED
