`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tf9qePNaRJFs2m77UptU0Ko0J9GzlkTck5K156JjB/G5j79lGrC9BL1Ky0nakAD+
r5lcEUJeZJfpZ0nGzeb/WfZ/fP0IIjNjPnbE+Db24B/BZBcYhdtu+hvsFUf176YH
AFPOJXCgQvo6rUb9qOh9F6VTF3sQ+nYr/GvfiD6dJiMVfrfFSleXqBnv2b99ULYU
AHsi+1IMhMxlj4/lKKm8NKXEzXg3W3fKr+SKqDCB0cRcnXLcKfDGnc24ZrRiV6fK
hzbs5bkBzXmrcMmaY6nw1zw+ztlC8a3fIisXWyg8bj9djrhw5iATh5JqnugW7ycd
LucUM4zRaisBmBRwhtSqJwaHJRwKtU4okL2afdUDYRG7lrgsg3jNt1tZzCNIS+cT
m6UttulrnNMHdPF3R4eYxTi7DWJWyS5VmYZh1+oRmkaeuJmCtpHjksvRYuefTXQ7
yx4ELvGz1df74EKoCg5hs0DY06uqTT3zSMAoxNdLOVIc2Zsn0GkHV1V/aaErvkpS
FZ273IFc0rfapU5s4sXUIvSfGZ7RyxQFkGEgROUF4UJbSWw/HP5Z5SfxX6Pze4SD
Tpe38Qc6A49ECu9ft6PWMX2USDlGEXTCncqVugX7tOzc4u1XzIYf9y3aQWzeyZBN
eX0YZfsEfStUklFU92J8mw/tdZXu3CRZfbEsr0SoTUkMdkleLZezH6SLK8TztNi6
TPQf0CEK4naNXHrwMPa3WsnNMw5SDlk6Gp41q1SyDYdQRLPaMyaio8m4ESx/7DQQ
pJ3Pvr7LzSDzxqttiUyHk6XBbvVzVq4nLcbo7tb1SXgSY8owjiX55KbSZHtRMIkq
EDEIJ/PYZOrQbXSJuog4ZW8WJBIUcDlCDNueMHkPaFmpgQhjCHd32VR9dI4FmS/W
IzyvO8A0M2Fpu7ayNsR1pnwddMgoCpbJHBopDwMYLxx57bllgdowfUiRXEGBc+Uo
0pACtBpTUSo71x44auYRRxEptLitUJI+10Tm6Bl/2+Tbnoo6Jq+pHt6ki8moefVz
8ij6U+2CqpPhHA2D1dDqvUq34xuTDSM8ukiDnwiZOjp+yM7C29UBLhZl2tip+hFo
Qig+uTy9Dhyexdo+mkiVSY+wgnpV1XS6dd5pyqEo1JouGRx2wttwfNTHEuGc14ja
Dk/WfYkeYU2UotP4PZR8iPES2jogks4lAUF8q+wH03M7exy2M48zfCBByRePYNP2
8VtH8JGIHy3CFfJp5UjNe4TFr4LJqicwWh1Lb9REdnjtxOd3jOPCkY9pUMBgin6Q
vdNRb35p8PVUXCl6PhlCq/RTl2ZjV+ycGuQNoqD1KLax0SvW6wX7dg1SId0ERujg
knlkbHDBC5hoeYPK0EKOXm86HN6l8HkJilnuXH3VbCftffQTsXblv1BTI0YUgEnN
bzUK3nSrhl0yO8VWGk2Mx4yjAMTfjoY0c3cXde63BLADGGj0eZC44th2cHmZKljP
JAujWdX8ij4bsbxHooa0TZXcx5PP+KiV7BcOfb17cUZUvOzjPpAY71gdaLYVW8uw
1ihJWVxQgIEZp0mp6T5zPMStpzhiBs/rUfjrRbjPS9joKTBc/Bi8lIpxq2odtVWE
V/qvI28wOcZ+R1plzOWuvYQTSd7y4sGBq54ytxmXBKJgb3oTUeDC6SzZq5Nx6kGZ
JCR/ZoZEKpX66vMazhDmWQtQ0GJNjpQcTRuaW+ocz7RiunpzsCEAOrN2JMuQmEa7
4byH+gsFtWE0Jxu6pUUOzdJGGPlmu2/E+3EmHjw4eRK9A+QOIY1lN8/mwGJG9FYu
Xxvfek1CDFbN94bka4nKegq52OdO4yJ9IFsaxUMk0expM9EZSi959isI9NZkruyi
CH1oLY8u3cPHaVS0rRNW67SmPCIfWWptgsUco2F6sndikfjyw/D1MpsIs1pC3WSs
RgUqChw4EKivu1eZ6FXZk8jaVkb5iJC0BWmqHM7OGnCJjMrxKuMpu1UEaqiae7A/
wLj2GMES0Z2MXTYUzWx6ithaznYPSvtuAnwtO6UwxzyMWeTPTw9nifjEJkjM745h
gLZjG6mh907UZXwrDqzrbWQEkc73lUGTTn71P71iQ5ZFRakm3vQovYdIUymbDjiT
tU/FYXjspc+WBK6xGUaB5KIhBRLdyl2fGPkqUvyFc26wa5dzmK8+phxIv1QBRJh+
zMy24Pc+nbALP9zPlxwoHpP8og6vh8f2s9k0rZXy0weI8iiPEJ4jsBysqP3hECs0
5k9de/OjW7XvuCpjAUYg44aMQ8u4P2KAglum1QOf4nb0tsxDDdF9KjHpcEgsXT5z
rncp2lq1ALXMGkufZMGosLeow3kHkppDW7IKaIr9QelKPox3fMPINgAB33TWdPHx
89cteCjpy8/MtiM4/wDnJM7fPSGRsPDpgaqITpmNZcKSRfQTARSgKudPE0eXTOkZ
8X5jALDUa8eBVFx4u6k9n2Mi4BVQ+0Vo00J+HMUMQcV9iQ/dI3Zowy+uoGnhNcf4
+qcLjOTnS0LDdpFSjM+Tiz0gMDwBvQ9qz3Qnxpylwqu1PYJt6qF3FZ/SDHbouYx/
AYYCrxXAUae3j4IE48R2pJkB3uxnsC30nVp65TEghUOzkEF8U4SOIn834zbHRZAc
2HN9COj8a5eKyfMAc7G0s7EaQ4nn82moMkMbkuIcZZVt3X0GpMDBdTsVg02ovEtp
Xigbe4dh/BlIxKxCux5CC/0WQ/nkq3gbG2q/qp0cmVt8ThaWcmZJ0OfWKntDONDv
MPHRjyshi1QAF2v7kUGT9NSNEsUW6VIxWbq7CBJ8QLGYAZhTCsV44QKgYX8dglJ8
XQAtUC84h6vN3qXb2R3QGcZCh3tojSyfgSebaEQfnLp2cQ1T3twOKTl0r4XOnsTM
J/fNq/+c+MkO76SkD0YEbxT0dKOidd+gDEXOx7xA58MwGVRPvez9zgt+d5b/Dk5o
CamrsUzwQ2nyyJ8Lu+csJprAxzBzIw6AqcFvISTgYff0D6MRMx72ek9LT/4tjixY
EEXl1+VmtD414jxtdGLkQOaLcojRdo5jVaNsHfb/XU67DmiZ8X8R1StgUfQuYSKo
0S7eRiNu3wxyc8jVdbVH1Nua5agL7ryjJkO+AQlBN3YXYf4BQUQDdwTLGhjLwKVP
J5hzIi1DCdJt8+JRA5fQX45jhyalAqWFHy/OqqJoLNYMhZKBG/34uRWXXDWwsxEk
2KbDnr1TsX1Zb2zeN36JhogHwHm1ZAvEhM3xhLaR/sqI/u0mqkC9caGj9mL5FMN+
rJhPDeG5yYeHgUfbyyxmtQC/NY4SYvn6IzLcH6GbBDr2tRJliciEZVBV9hmVOOMA
xYm5bv0bqjVPlqrbnJ6VcUu9nXrqb4u0FskUIpMmscN5Aj9uD4u+JLymZgW2txuL
TXdOQJJhVbSmik+XrFHEm/LHdPBl3e101wjRVcG5ysxRE08ODacbWe6+F91Gfnw7
rJ1xmT0tbmF72uKG1IgE2dSanMJKds8i40rYYTLePVKbutHAGjmZ8uhnB0j3Uyau
k3+nQPSMbUlza9lAL6UjjXsgRqwd2UthVBMdekEh+4slPycWb640aANCbOFg/lnI
Nkeu+VGe+odNcml/C/AYNCO3qAhI/aGQHJ2Foe8Y5+ElVmwrNzvw5uN114w6b5n3
5gOxxpRBqJaneXAs4vxmUziXinlcibWD71HNxiy1YnpGYJv7FQmwrbTMXkEtham6
/bnM2LtCNiv6KzY5xI4D6lqX9T0vvzuorGD+/aQKoJ8HhbF6ieV36nPx66hibBHb
LND9DKAFMsCCMLw4ANaNGR7vti9F2GnEYoNO02Jbuxkvqa91p1cyHDQuupnBAbhP
yiSC2E/pILOqQNZWna+lHzsoLunHODTvun1lyTlUjnvMBEEl9n3bsw/0VW0YSaEl
Ie5xSCI+7LFzUEnpixedDy/LEShHxczbEBK/o1WOKYC9nfhApuwerM9sZxq59I53
DN3tOPAa4i2DOh5C77H4LT0NJmDnTVComiKGjn4h51ckTi004FTEAaZrA4Jm8rh8
aRk2q1LpL4UjkRLynglAtX4PIHfMsm7UbpoP4hpg3j/iJO2ZFccaIkhwRZUCV4bT
lIeA/E5nnd9A0iW/SxnENmf7DREfv/04iF+kL0VzkjTXokFrTmSz4hBYpiGYz1Cv
2z09m+cRODVRBoNagEtsatJiwvUDVfslY6I0m5uU2Os0uoWga5sutwXNbhGMoXkz
L13E0qZfvhnkyDYgIeOXCVYhVEp4hydUDWMx7cUHVJtoV/OYmpxYpbRrBhzdAwJo
71ppfuIqHNRb2g2YmTj9Q+ACJcqHWdWVjTnJhQPTdL3kz2Mzu3EU5HfuGk4XhB70
rE+vRzlimgp8yWLXq/E72F1eWtVYMtEi6NrIhCHjSBgAG964ukfAMhQ8OnvTRezj
WvA0+FIWFWafS5+YQotg/iEtcvxjctbiD4uV34JNcFSBB3J2JOfLPx/YZOWS1Hfa
slaJ6ZWjhtU46l2bsODU9yir3G8N8rue583cl+Aicpa8dZFT8NyLjkijSPmB30+Y
2t5gjJY2JYdoQg/d3qmQ8B2B6byoA7Ia0TuIG18sGSChKjPArLatZlUL7kmAM/kU
b9kjw4mwih6lDt3B+aK9TdeJ6YZ9bYKuVV9j6AyV9de1d83ixlX2PSC1i9sQuCYI
ZmpB+sxOLGhEWeo6TlLOpdNTFBb1rpP36nQNqfqmtwleANIgkfkW89DfvsTQGwnP
qkfSCbZnizGiRM5j1TDhuvnjivgUOGVxTDVhXaPLRwsDx2MXmtdel4X57E5o/gQu
NSjY0OGmbuhjhFJVOIwuGDQCFt8QMM4PTqok6FeVDtZf/OAh7GaddPIIGW828Uw/
hBKIoxtPXQeWY9wy7N4V2hkqMHHQwVJNu+MHi4xbrORTUYUKerdP3a066e7wJ1kZ
ZN3SJtRcvOqH0d+JA/JpZTVpaCmaVm5kvMUO+jeU/Hw2Q6AUc+aWG/tbMJMVItmV
YaA9dgPnIRQHCN+yLReICW8S4DQjkGITGevGg88y2FhpcbyQVDQOStOsyvd6RNKu
f5BhMQ8Bp2MU9OW1Shhgte4oppB640QfbjDvTbJ7FpiGXuH/74KJCJ2llGBNFdQ4
MtuMJct7YPRP7mNXQSQ1qiE76KBlIQhCGcE+8U3YN7u3m4+yreH4f4AxG+nJEIN/
3RZF41lVTQeRqNlwhbIf00mb7bDH0+WFT0N3LMxXUJQU4JI6mtwbVkflYqyhHuKD
XHc/1PRZ4Gg1yG9spiL3j34Mb9KQEmwVZ58b3tjYUbMIKc3E/ErN7IlQQW8VM9cy
l+agS6EccHWEvzpG9tWHJUsZ25hQ3w7E8nyPZ2xdUmHHwaq3JSxtGxM1rtFAkIJM
nTfOE9IPH3fB4A+Ls8PmZzs40skpbgEb8nJ+YropR9SJ4pZ7essXjnAt/iSKmoeX
VdSLTMA69fBeDmZkiq/I9CTRB/s3zZhCza0CvKLImFm5B32oJRkXXXRXKTZe418P
KCt/bidmyHWqfb+9+DFNdBnO7HPMWpMZpHw1kN2T1AYy6Oa9P2lu8EP+UVUAdSFf
YrbvTxgDXQD3YxJOPEYhV/whH3wZz1363x1ZIVV5HwfZUH/dhPbZRK4Ogh/7lvGv
r0XCSY59hQiHHdOQfFjSlQy3/tMnAncnslZychWZQpmbIWrncNVDit9EXBuFp/n7
nfk+Rjl0Q2ak2TfoFvJsbukDus0WZ18vTwDkPBy0OzkpQIPab1fPUgDJcfzRBdW7
AEKfHmtWtYgIj9xRK7229uF5uZNqLRtyHJ9nB6bHhEyTwqkphimOE5jY/FqzKG+R
35t46legvi9Kexdk1mljY4IuvwSPKXnjGojST56zs8fsS4vugEP2/JvsgjVeKYVL
Q3MzlZvemCusBi57d+Pn3FNqvfan+9ovUnw/5pd5xT/TMNVFY19S2MYeSPdWmFHS
re8J1WoiWtNYwGMFVEnwYSkcOzSPztsETjg9WdhevL4W3TtQCbLm6PgE01JBQhFC
3Hn+f4piaI0m9SPMzLZJiVmVmR1z4/pZ9GmmwHF+gxkgeI66FNQpOq4AmHOKhNwu
Xb93136WB3pbowlVAqVMoNRkyrYbtl92516ik8TvTpYH7ev8sArXgw2FjosKPJAS
lBKCxQ+3bro6FpnNnOY+j8tssxUbVzb8nKR29Hwh7cTG9FGHspqF+t99F+nvvxMP
FeKmbGLhvvCqjMSDVrU19kIlaCHUn8ALWzfD9GFCBWPI8a3920/ojJK8HFDdea8g
Rra0PNDXU1p94LWe1cBnIqI/DVnsLHKtAas4JDIX8KLal8ru5SJrLE0KPjcQGdpW
pR8mfM5EDx0guzDw72V7WzDxMBeFdmgHohQbh0CcsX58tseFNUtjot4MzSqBsWKB
X2jKRx7/sHjJhK8Qe28C+LbpJsOVPp7vOt9bttMFMXR3jSvbgFQJiJ9Ta6JvqqwY
TdCvkiJXWRahfoSxHkwATy726SrtEGceJoPsadnHk41lFF/3j4Lju5Rb3tL+MNOW
dI+AMBHJtwyQ2y10OT9GsNqQqltWNydL88v87VLDcJPJDR9dltcS3vcRNVM96BO7
8eZDmLGyu+/DEmjyLLkGzpFQ8op/40hSxfZu2XH/LZkaVbKFATpM+tHsvQIQOfzG
WMN+nWvgOBls1X3Ng7z1gkkhliyUVIxEzcb9TqiTS8ONuG5C9a2Hpx3uW1oAmFg9
ZWxMGUApfR87GMlHJ8mbuqa/OfLjxCA32UvpHZCfGm+cjQ0PkcIae1iZKaMViskk
1vKOarb9ue+rcE6DvLlnlF2eyDDuUIW1fDJ/JI2bBGGBuC68HkZEBl3r7ZM1e3BI
ZBLP5Axb9QPf0xkL7RnBcOvAo6hg01FOhc7W3zkOeRmmNLlOkeArBjQMs/maLELh
Pmvpr8S3rHyi2TndxKDmfGHEPvLfDexGDT+QOMSTKVilLeZRIJYUTOeBwymqpLsv
VbYgtA69Y5CPYKnptNUIXUSQRVMyb/nXe5fBkUQ09Ihv+tVCQzcEhW1aH07gsAFm
Hmyt/03i2sDTuRrdXIxEX8o8ZE8BzGkPDTVz4FoiJf/bdQNXZLcflqyLx6XsTCPl
SCm2Ehzjyvk4S/COq05yCTvQ2b0qeyWncIlVLAVX+RxbMXqEHkcPA+DojQNuR16Y
ieStm/pwOZVCe6b0qEcoDDa8VLGoMvF5Jwt4mLek9/Q6Qb0dz3YfRYdfVG9R2T9G
ftAfq9BXCLJFlOgdYKB6nrg77zoq+dntZyVIJnFZXJHlMd9MyqAUZHqJ0WAPumYb
HQLikU5Yb1Thwtv0mwYp0XDb4PrK5lfZofffBHcqgHqwSj5yIIcUTF3JxJQS9qP4
Zu+01N+KgJWcPispTuqhUw+3X34OIWc8h0B1hIzyGGcWI3wVA3Mjwc5voTH4N/Mi
Lfp+94R7O9p5XPd9uW7p2wOtbqCjcRGvfrqCI5LzQSnzkGphDe/UA8ZuNQsYBHH1
nuFJx0nnMmI3exH00je5IS/ZER9ZIc8mL3ncX/X9cGl0DilcRikCcTSu87yapYiN
tBWTx/81EK7NK5iaCqk8rIq8rWR3MqsWH1/QZA9sUASVxS6T3H8JFpNCWVZH9hvP
6oaePtBtHVyVqO4Z+m3peQQj+kOTDjtSZOrDQfWCtVN1WU8F6XzI0F8WjOVmJpPb
SGsE8OJq3izBPBU7OMVWtS4o1cG6JJkNpontSrkqj0bo16Zxc5eP1dKvWWmmMseL
R0opGKt9MyuWV3ViKBpo0kgnkILxENpJIPgBQ5pFQimooCA/EYsvQKSFh+hTN69S
qQf1hQ85i+dLyR13RncZIPZz6uuBEc3d1LcvKXjDitBgZP+qpHvh2ZFm3WXTMjQ4
KOo+U1Iko/ei4zM0VM09lUZtvTrkwTStNm0N2Wk/dfhxbc9ukNCzj40Dp3BrsGQP
GhHuXoJ22bShcYE1K2S5U9AHt0xewM1AZ09A+8UKCitAvoNJe9dQW+hyCv/hyTtr
W2UjjAPvOuk4KFgcFX/lpe4292nbr8FO7UCjgrXmOIaWGlNJCA8bVumoVxZxN1lf
J905chxb8dNB3RvNhSnrrSGqr4A2JaAhxl3RQtDEg9QkJ9LkpPs1WBEglaFukZdB
4um2PtlHujLvX9LPblZRsLLWRS/E3v7m0dvrKwwXHYni9tWL5s8bV6QCBmmbmt6h
051oLvG/OYO48Lc2IRLaOMuQUDTawQ3oJjq5Gi6kftXN/EHqeHBwrq/nfwE4peW4
Tpuwvw/rD7n94hg+gXilzj+xgnteTtMzfcusRlqO05qnyKUEn5+meM4cW+OOzSR5
c+G7Jii6bViV0UjNyHoKGgwcxrb8GhlcCSa1yldF1pMRm74zen8RfZo58mT09wqG
4s/saWKpDbP8+ZZHflJ927gAzcC8vlwuldRozMVx6MDZxk1cRXmSeBwjC3nOvCrE
QMZYD+NoNasMDQ2Q/ITq+vHCFWSIT4gnrwMM7JGYqWDqZAa/3XFz8TooV3JeC5mf
7gC66+l79aV2A6DE6mWwPFqAN0Rf4Wfx4Qf4MbQczWqhd1MczHSgF55/jRG5vxmq
IRhhuYGbHF9A5wXBgh8tyw/tf9tHN7GObYWuPmRyYqKU7D2zJh1ulqpj/ZlhUtmW
oqkwuHo0QpgcxC+6QHW/MTFrLvz2xZdr6OkqUPrILR00lc4XM/t1o0GvGktgu1Um
oulIuYwQWvAOQ1S4GXTmL2byWWSsZj+uR9SRcgdzTXM0OmVt2UP7oiDm2LOgLOjC
y9U6VWfdiU90o0ZBoNu4yO/Jpic9Svl08QdOyB5uYUvUJvdmXbjlM8/xacr9Lltx
O9tGSBjyl0JyGUqIr5TgeF/LuDwZrV19EL+lgTksSSECxuR3fVhDTy9bfjwLxBKp
D0kGb4bo/cZx39DDozPgylTjaJZuusAzISoTHp5pqoK8T2RIk63X9mANOnX9zH36
zVj3SYDS/gKxXWJJbRLbDhUTOip98yrU8PKzGw0pHFoLd+p5YZyk0fDp8YTH9L7c
gVcBS+Q3aU05EIqTHSEBKL7excoD7MmkoO/qnwUFJOZn5Ul/U8dxTG5Dn5q5hFeD
vCy2Hk9UtUTHJ52te5iP5EOzgZk6yXTKB/IloprA4nbSciDSPmjeLagIAlHcLTqg
PmbQJNw4g0xczZaShGxoSPN6ysGO9hpQFDAT6E0yfOanNNqHyfpQLbfKZX7ELA2n
EnY4r++E8qsdiLTHAJ32r15U+Y7+C6TxZYdOturaAon2EaDIohy/9pMlEexkN7bd
ULb5nzF1VR2n3fYKDqAynWnInd5FUeRNTmFHXM9h/Zx0tirlCHw2neB8ecgxcxSJ
+5wBiTdjVBxc3OeMApnF62WuoySm1Ocvn1MwshlXxyLGRuxcN8eg/N7GF7Fbye8m
bplU9FcMlKI+w860iyMadBibLTrDkjAvmw+oTk2MReWyhl9/e0lK9SzTjpNljKMU
vdZP8Wa4vPXAmB3KlFvDhNL3rrYrZo2pUYbpJJB6sfZg7296OnR2LwqkYNGPFQy6
jc50zES9xCfE1Wi/2uB5hPbTuHxeSFsyapAUmdYMeT80MJHuv+/YWx1LI9jHl2j4
Ptc7R5peicCKcnFpKUU2J/Ir+Ob6xs+Dj2nqppIOSG3a1AZyNgsZH1cbKQF6T5Nn
tZ1KmWVHyAi/KlqGxgR8fC9BrS9qr6SmwjMevJzYWjRLFVqLbBcryCiFnEUJcIaJ
Pck6JhPXzPP1/AOrktL1cpL+YpMjq847AzgmKrXifpJEelbQL/1om93N1cPzoagq
hZ+xYZxOhTtkPgt5ZuuIOxs9OfP85W8q0t9rtdTylR7QRfRs6qDZbkR5KT6X7IPt
jDEu0Wq++0yWZMclQmjpAfKNVt6S7S7HdInG2y3SilYF8y7JXArNYFT4bRq6iFkF
8CLHEosAtYRgePV60GBzB4pLnUfJAsxdsQP2bL/NeTbgNfMTeQP8nbt/VM/pPIIO
ZEuLf7hfSShKUQ6+NPh1hac9R6XUFbF7gzEXSwo7cn3MSEyKCNfcH4QAhSHqLX2m
+vVrUlhDd1iuoseLcPMaeCpu9DqhP6uHvYEXTpJZepQ39E6KwQ6vBxX2gCxWvNvt
F2KjIaCwkDw+kjNLscQwSMvfjwv0fS6gszSnA6a2XFfppWSXMUWBAIKKPHN0XkcD
rVXpyzEg9Jaz2c4ZtvnaUhrfPxOPmRcYAiot+YVlh5aCgFcF/XKB5SyDcf8AEASU
eyYSQw1EymDGeU/aORqXnQG+ju5BzotpcJnSrvR97Y5gGuKZyIOrbKITDvWuYrbY
nhMV3W2Vdw/1mgwMgAClKUSlSOiCgg0mWwyUyKeBh3EmchZaBSUMDuSzHZ1GW68/
K66UkK6PvCGY/byYiOugAJrAcNoIyCKrgdFfcCOpQ/8doT1NBWFypPb1lY5OW9mU
mop2gQ+EhgaS9oOeqrGm/J7eJA+JBVG4nFqirrZAivchmCMrGX30OoZQhkL0HUjp
YQSg8ypdFhBCKjS068lg5R6hwGfFEXb0Gm/0ICLpaABVywKSPa/4AIT0HjdLLYbU
G02+39HWSm7lwbbxXCAOnoXfcS9STBraO440UyMlhXdAKFnFkYYAkvhdK6JLCYTm
axBs3NLqhDcq5mC3pL4+3aCDz4StH397NsDt68CDZkc0v6Ryh3Hyf0CoQ5WSCYH+
2M9JAZrDR32liWtsDvtTFNnpTmBXoRm+AGsq9ZheJP96m8MkxAWjoAHzWlnhXZYL
71sV4nUVbsy3k64ERI3hKeUa6SX+ayT4Mim7gXsEdRh+39AaHnfcJo5eZGtYsqvx
4rTSBBrKE6AxAeiI/qn/EcC6XwO/1V20dpfpqQjiQG0ybRn6WDoklh0SGptc/+t3
gTWNQ6jY+9qLp+bSrNE5IGhhmuD3+Q3vbc5DThiXeGnGEBzD14SJtEbDUzffiZP1
LRcEf1SW9gKGJfrR24ulqhn0adYG65uOydNC41YGbrp4tpHFLw1DYj9Vao5oEaTB
Qbx0M+J59zhjlUQCEnomne+fFEyTC8zbc8Z4MyshiRxFwkeqMBZ8BtbCOWktezx7
x7g6NQcO9IoSruB3Aa+uAmIzedWj9QIfWAehH2n2MOxWGi3XxstUw/gtro5ExlFQ
pDv7tg9C7rqP5RiYCIML3EIauqrUzSemYt2MXUuT197cRXgadx01hLr6NkboMSBd
MTO/HN5Q6Z1Vc+biW0CBBkQtcKUy0z2wcd6oo0YFDn6n0KXpIkMvSv6arejFGQQE
8M2owP4YmbSXVMcL3iOP+/+tMweSp0gAAsmhO1AEGVDrCHRRZYY9KUIXqyhw23Gz
JENeHaaIOEQpHUKyHMMuOPdd2J35vQSRwIBjWSXg0QYvxCkeYBoz2TPeNMhDBx4k
cuPkFdLPBaKyGQeD8HkkqE7mHd6ef5O9iw/sf/FWofL9OrXtVoyrW0zByV/xsf83
AESP8lLraCtGJhhjARejBtZEfXxuf3GlvBOFP5L3IkTVpG9EVsTqTilhifdrNW7b
e+XyCKJ+mWHvHbcUg24ciwUzraIaNbmsLArdu2+zU/6aw22jUpW2+6vAGHevqGd8
m4BEQr/hdEJ+sSlAq9IuBTvD15I0GbrQvPFEz0Rds5WHRSv7WrbE1gNmyOR8yYN1
GfuLBoi+AxZd//RHvtnRkHy68q9vcWbDKCna2sRC2hPzNamDjV9CZHjVWa/sJD0c
gD7WEJZ2GaU+YZwISeqOU7w6zJxbI3ty+n1VPKlWG8vc2LsoSl4ZXiGbeImHsE4D
O8RvYXoWuSuB5FQHR3dt9fUl1vjzpOp4q+pNV90SGr5hfI1UH/n5LWwLZUflly4t
/mZjSswB4SeYCj7Xn+7KqkvteRVR2TF6gfL9vCs/1I4JGCI4aedXZxf8n7EpA7Y3
0dwwNI9+6V79cPD2P4bx6iRc9oBTYOwQcwoo5naE4Y/DUbMkto9rZg341D8PIXVN
LujFf0fEvt+SOREm5CJKenOBGvIx3O9Uoe+o1n/C4ajuFhm7ae2Tk7vNWJXrCAmB
mTisKUjx3StekQSzV2aeYwrv2ujb6qX5FIr+T1bslKxZ58AFkQTaUbOA5AkhbB/c
S2eQeDc++TaahlnUVt77VjdKgj8Pb1det5PWaJu7NdaedOzmQWPTX5c7Y24rE7qn
eB2EBqZyQGWSzq0UXZ0GsqFy3ypT0NeI9LJw8vpCRQOMwhfuddq4cbZeCQBl1Skv
HEDABMaNH0gtBWXwdnJktA/MU34Qc/brGh1FyCZPOi58qzP8WOiWKbisiapkMHMA
jIBDt9YRwl95cf3upWPpaUv6EM5PnVKtHBKUGvxyNpSHNcg/4spRDxp+vgyrZ7tL
b/dv4jj3HkYSwCaqVoPvjFMX8mZ+liJjVSYRJHRVf2GwtTqFBYjDjXLE1lvRCjUs
8K5Q9Q+3CoYBMqHOhTQ643AvvZlifwXRWbOl2VlOFdmf90vJU9+e0XYD16uJVeIC
QFY/d3ibty7b76JMUOBPF9wrrE7+NKWAOReVcnFoHGUEzGW9YeGuQuVhbdrmGBgh
MxSAwbaWe4rbAIGyMZOMUwCT95KDdyWaOK4mrdfVxScIJrsjuUY9Ks3dLZga5sw0
HyWx52I1kQcwxjVRnL3Zgez/xebHtq4Nhl+sZYcUu0VXYRHVqTm/zs4CDFrd9CS6
3l8Le7tSSaNkEjebnEELQ4QuEy4cJ4Lk3L9RfWv+sYHMYHPMmxUUazSfzV5DaQ+l
3+jnppH/vIZ3ADkvs+Z5i0pe3IxySOUOHS3qJ6JqaP0DpXmuTlOorT0QmI5Uuxnb
0tjaug1rM69f37ncsWFWUZ1Q+kKiZrRnajUeDURjOlmkJy0Hk91JBF31uymgpBZC
iE/EMyCoPVRo4g0okFwta4v04Z+VbqP1hAfYbtggejqVSgZrfxyIw2G22xR0hyMC
EDCAG/KsL2NBuCjiDFdOfM+MBlhDgwcnPh2W1xQL6E7j8/OJ+9nu8XEiWXj/bbC2
yTR8R3har90gIcBAdcYRXZlR8m7LYYX3Wjb6GGA6qv3T3a8nGNs4Bn8PQ72RYxhz
qGFaDETThqyL2oVbBrRwiwNbR0wugXAmyyrPJeE/yOYdzjfNORReqo5XD97VGPOD
qd6VtZA1eOkkqJCSTljsB2do4/TghALCCy93Y3BYvlneZzVGnUBRmSf5eCup2BT7
661iYwLmZs7WW2p/LH7RkzRffPCw2lLWWU8t3GuP/J4mwGO+928L1fJqLMzRdVpZ
znMl/pVzqzgz2L6G7oxvuwOpsEpBA+vkOtptStGrfA2liTX6LXmLW2GroAaQYKSZ
rA8SgmHdBkRenu401SpkQM1atkOQV468jCtT3Q5cLo3KaifkyJ/wLk593t8PfIxz
SSBg/+JayH+LDSyWwBHPujNMu2hkpN/D9XFNnBzjQbHOa/pdCTspePyp6wyCpNJQ
fpQfYuel6I5iNE0sDB/7fCPpSPiZZ78ZGBW/otXcwrK7HLO5ysEsItx07bhpRzIG
aLLXI/Xmuo8oWUKU0KQM2gE1xZZalCltniiafN01Ekrc+DOZiu0BAABJQWmI4oBA
KP2srlxene/M38tf19MZR5rbFbJEWUw4YOkIEO4bXH4TtOSv8RBTyurPp7QHlCVh
YgeWfGNUImwHnl1qJyenHS+s9xhtmDg4EMyEGAIvtDCU9KHUZ/phWcttlTFS65+k
kgNX//X1z/zytm/7wJo34lu6Fw19phmgilDorPcwTiEnZFkLr8mugVALtA4+ZnBz
bkJ9q2tXQt04AswHoCaGLSFac4a17QE4bY0Udq2vBTdEMRRamv7adDC713LP0JaG
wvZlLOQd3i8gxfzJKPDxc+UXm7fRLW5T/woQgwJGeKljEILXIRmvpSTGrwqzY0nL
LalJN2A4y3rP/hID1YORoPhTg1Y7qiq9QDnd2+AA3IwkOyhX8Uk0go36Ksi6y+qT
35VOjFV1kCISfruB582a8HbU8Sy3EmvnZtMypE2JEMLZ8NWG8ucNjYajVip9M9sA
PzQmt+qGoWuhw7vYEeA7CRyAeK811SICTxGD2uN3OGEg6MiiU83z305X1MrkRiFj
ed4kHZOm/kMBrFjkGnyvPnRT0+l8hF9begRRYruqYAE9kjixuvU3JURQp7KXXQPl
uAtrBj54IvOnMTfRvs+DbJzhBOjmNuXFwj1FIAH3hfduth0csLu5WdrFgd+Rnci1
RXdZxBrvo3mIh/tyMN5wMDsi+xnAKj6pN1KonOcGIVtnmD0h0Rg6LChmYhZbkF9J
765y6B8y0LcXTQDfpVsMYWrB0ENdhJiSJ32fpqmnVYkgeCcUfX7MzOobZja3OvJ1
4EFsiz/kxPLtxIrQjyIa2KclzDXdjDVBQQjCOap53TSvP7fEvezH78HQCStZQT8K
xQmM6whljv4FLSD9NvPZA//Wl9kLNOzToDi9qOG5DkVrWBXGumiZLpiNUA+5CSIe
thxexA/Un+lAtMNZsb60NioCoOPU7HQ2n3OaQ8wpX/n92CRr3pm3BX/Ax7hv8ptm
IBVsjMIoJANFMzjHUavTh9wHGSianARlxie0j6P6LbtFeKOv0iqsZBFTkzwvbqkL
JGLz3vAzn206/8g155A/Hrdrv4xHQ/UI5YgPoNRu2kbR4FQgVemSCqvc3J6R9G4b
NGZnKtQVOMf//q3q+2M1l8kVIarvat5ii+/fL/Phqd4YRC4Ryk9OauL55uDB2Vv1
RKkuNqF2gQ2pLDoVSsT7jvMBXmwVu6uwLFP2AH39rXLkcM0pYwy1nehWqEipWH+Y
v8+rHCpDK7Kkfy0flb/uSIf1j2fYZMVePoUmeV0SMNhEqXlOif1LKbaX6oz8MBau
Hs7MYaYAUbGhxVfMU1VsDudiCYmiAjjx5pCQLQRR2Bt1cTxln14X7oinZ4sJdsZR
E0CZz+w+iXrZ8hiz3R/xi76GiiIyi174KCZy7m3SzsORgdROPYLNK3Cm/lUDRFaC
pPAJzHZ3qHq25V/XLdCx21vQqrm+BAbuIcWS+0SFPnh88dp3ysolc9x4xfjQI6IV
aiSYbMi03gbXhKCvrBZnSjeexSijEMyAEGNtHdvZTW6OGYRSwy6zSydSlDc6S2vl
vNdW+G9LotRPJwOmz1LQfx7uU9Qd/oWvZpPoliaSiIF39BJJV2Z9kuWjBMMLr/Zc
GCVjezbNbUBUsRqlZIlCJfboqVEYKTB63ky4xPEto//QIxnBEoRLz6YybUlbxvXp
iic1zKQJqS4sY8fSmHgm/H9Uz9jOOpA6cfkNV73G6L79r3iGcN3LOpKgRdw2J8da
Wvnqy5I9cZUlHrELgdQu27G2JyFAB5RK3KLVBBuTIm7r9nHsjPkG4zNV/YDdLWiN
hXTM9Ea8Dwr2H/gb/HJ405l0fOlqohjce9AiRjCcMeeseTzTCHqBynNqggqMrxay
RbhnAk8NJjMIwsGZ3nAHGPGfqKL6dbf1S0sSIfjah7GOO318+/aYBcMdWqWrRZKK
OvAXJBPMTy80CNbFrxNMY2icNVEfQIxDd4lb+6A4m3xoacKK/XbfaqsJH6/fxXoD
0+Pk2G2bR1/9nuHJmK9vQK8Y4Yd7JxvIWSNFqTxY3Xjf1yl8Md6MtLAKK2ObYk+P
vod+poYWE9eDBOCIeipc96Fan6dxEGxfIYqW5W3SiwiqVE7rS1grNG22NW6006VB
JnpPBm1+8RRMwXvjZTtXxLfbbVZ9ROoVYbPXnzJAditG5yO5p5XnZTlhEKqEp4zv
GVjD+8VNeQzVHy6GvNqeyODbYsx8x5icOlFP61d48kwqd9XJ6aityUjUpXXZ21qS
CE1iZIhfzmmwdKCfR60YtsnPCXhzcheKfGyjKgc+nkxu1mvziTcGPk2T/rFbcex4
bZekS1ltF/9LVC5X/Go3rdFfUUmTRCFVFZTeFGd5OEBrXkOJ9XSScmL45vcg13fx
2+tL/b5wJ/xHYcKKBnSQfF75pnHmcrJy5kTLGTliH+KDpGk9Glpa+7/NpeA5tXCg
NrXfoDgCjFlmLPpvvv55si2ZwIIwCm1SbWgImMB3G5NmR5bS1bF7Wus+SSYOgRBa
L1aNTRNpizP1yotrBeWS7X/Cq/rpEGVdsHrjPC+5YMIQGsVr3Qx9zc+DBqmiSxLC
VnEqGBlwDp3i2A2/4IVyGViFTZHDjF3YlMjsExhf5D/BaGhmsbzWAfn6Oaa0b6tV
iWnjdP2J7i7KIXPKwIbgLUalohjrOPDHqPlVqjFoCf05AEIPhhTdeu7HnKaIfag2
rvJcvruEwKb4Hd90KOEO9YeFczHrjfG2O8vkmSdCroiSftY+sfeYsOPm5hrdrX5m
z4falOdau54xvzEmUIXA6He8mKYmD9mJsTJQjq1BjOOTyT/BgzI8eIDDu0aMrtv0
fRFC8V6xNHiQUfkL+wIO5q3MGJekF5aMf36LeSYEtfVMCFuemqd03hOVMLpTxuYM
ytEtejms5jlQfzNcuXJJR+NN2KEJxt0136Nd7/bIRFC37EmL1JXzpFAoFB1SJiBg
D0Y/QNzTSqalAM3HbhrimY7A/Cvg7+P/M1gD9S5MKQ1lTIG8bngSLKUjlBDgTc/O
nG45MxNwNEUQqtpMzMsBE+P75n/95DpCGVA78HJ5waed+EICnFazuw3UlB3ySeha
zpkIJFAV9X3UJZjH/BsziiXV8c5erp069g1FhXdeiuD3N3P2hH4ZpZkNLQGqhOcq
AekPL9OJ0Juui/D7KgfaTA+WpfV0gYj+F3aC0KFs50xvPo0nCtwVRvCr4zHu8X1n
KF3L8UgU0JwKjvnY9Fa7fypX+akYSNXl8vnU2OzuLV6ZK19zaeX57+LSjjMSFZ+p
bfpDiTzIkwXTRD0YBByvoU6NGThqZl3AmZvsr3dAZ44fSUw8/1aSXrOaR27bHVnv
OgPcai+cljwPnNGvDZNFaYWN9Rhlw4jYv3e2OLP5tAdGAZZQzGM0/tn1Z9ptyIXH
JEGKX0/hlIBq97kYrnsukULOgvFruKq/Qm3LYfuO93LWA9MgsLI6woNkyi2U61rB
HnjXi6SoeOJrrcIFTbywGw3sI5iCJc0OlTOvjmcc3u3dVg7kXJ1zKqKNYBWi6936
939EXviCPjbJ35zyU9B9CXf2Bkt2Q5yVlIMtt1+ICskIFJw0KPPYzRyMpZ1uxjRr
LyWr7PwHmpBzykd0fc7oZdnI5ZipdR/ar3P34hZGhmHucLO9U0jJO/X0cMOgQUHq
pYDjUbcawBJPjdTXeDRcgwkybxPSuC6hf0eHZWTd96hdCRB0NuGDHtGkd+295xVP
3S24cg2l5ZgK6RCdNYdjnu36azdML2RIR5GoAGPQnFrSgIaZn3CSYfEyqKmN0UzI
JfF62o8oVKtmXhG9dJXLSRi7TT32xMK2KZZkSnfsfFSS8Q39HZR+2nKm8hULzkvk
WOnfBMwvn6sgfHgCgSdDG4DNZy0HjWkp3FninEenX2Y+jJQH2T8kppcs+nROjpTT
8h8EyW/CSc+Q0OHL38Pv+U5NQ4Ss5MYqUVcisFdqY/I9urQiR7OXFOtYqsUlZmoF
OtMuNuvzpNIANfAi+7y6NL4pNGMkr1/j6IKKurFGvoUPXfdhTVNYhGjJgV98hqa2
fisGHrdtiYf75NUSEE1RTbC35Kwj5hUiWytUbs6g5HQkZEBq+YuIhd95stcQnzQQ
O3OU8FkemiGb16KwIcdVqscfhFZ0qWtokGSvTLL1UwEPpbfytc2YAxtW6uM/4OU0
aNvb7VK4dPzJSf+BB9PDdeKKYyDyEbpWrSO3BQvM/tjWbsHzTKau6l6HC/cEcAqB
dp4UqKYxBstEfS1yNpii1cU9dcqQfJBuloBd6K5hej3ymOxNe0LsXFb8ZmL9IQTh
+rRdMHIkWuVQhqcEWUzaeie48HQt1NQe46VpzRjYPINZDfKj5HxOPF/FALHsx6rz
M2Rzxx8UinezEsbF8ePaG9iDwY/W/LRj8QztOH17eQXK/bvzEIvwxvY4WAUWDHin
mHtndkxVbGeXy7dYgr/2jIM+e6GAF88hQRo371GNz1RF9IAw29MyHKjSqBRN4VH7
p9gCIV2uzUnIG9iew8ODFocnrGONTKjkv1+CddYlKcFuJxXVrJVtrNcFKOcB8U7j
8vTqqVGj4hepicIzQF3VPYwi5xq1jGMyrkTG+5aWoNTu63BVqa7Lo/9VJGCwm76u
CkKszLqk4LvnZbkVMDIX0d+zWompMvnJtDzHds6/9LhDLwImkgeL1+Dr5ARD7/7g
WY/SjBmflOnJs0HvicZzKonzJ8UC+QTWITZgZO1276iLnCss/yGHEf4L5wJd25tQ
ffVZ1yoUZxZO7DXMvueLE/4aUYDmnfLpRXqK22XiAtaTxE0wYe8e5zHJa3vPFAoJ
2Robi5p/GQp2DtCDrEe8aIDl3/L70dw1KqJDYLxH9+/S0nKRS8Dthd0b/yls25NL
vTuPx74cGzfKgu+OIpTAtTzGbBGeWGvZmw02hlO54uuduN4uwoMi7knnNiM5422w
fFWikm9fQO9Mfp1/4mzWAnCRYkLxm68JFwpJeYZitO+2qZuC3oKtwIA2pQPHhZfY
NNK6rmyRNCq5qFTIzwGk93oJAAhyGu6AQkJE+vA3c2cpmpZ1v7+9bl2Fh2vjtHcu
CeQDE2vMcirW+PsJOqQGKZvgXAzmeWb4uznTbK0i6+BtCtSmmumON6bXJwDJl6xE
gBpfhh7BS8ENBUE7tHdYqZDnZT77mkIayiWSVHz87gJVd/NmsDwh2Wtt0Kkzr3L9
gwFIbtdvWjzvDyo13X8fcDqQTLvReIJvhZo+LXax4KbRSrQ9RGPS9R22KSzQQSkZ
r9LZ9xm+c8w07of+wKwBRDYVoOAicxDxRo5BFOq1sgotTmLTFkqJyCN1DyGRQSO1
ZSUV2bjzJiQ19/OD44FlQ78KRSjQfOWIajyKaqRBEiiRKmAPwDDCAKerjofpsaf6
dHz5jjwe3sAXYuxFOvoM/ct40ab5pcR+x/83tSUEjAlVOzMi10EO7k4yhb6uzarq
4WPd+QDRWCqFWwJL5xUmJJDcHwSjoNroJNs1iXrrbcaWk8NWqdrbJUgNBxBNzsUN
6Niu+Q/IQ0/5OgdmOZXOlSmwXlwsjAGyg7jvT+rtzk11fL/ZyViYg0d7LdWT8jqz
FvtkOwGVWNWLfdnoPBhBO+Z4jvC8DpHA+WHIN1SZKP3Ox9kL9DtvR2/9qo1nXYIn
qsrneuqpjdALnjDyiSdP0bBHL+9hrRFKmt2WGfUE8duoZOpoz70v+V7FC7DxQpSu
G/naJ7Jx3j+piDYLrdwdwlfNzk9w6GByHhhzkTSPJJbxaqQS9v/pMMXIgsB72N7Q
71oOB13GUoDkJZ3GFyVls8KSv2O4bCAdXhP2zelIyxsOZHWv9jyPSX1HU+eNrgX6
dJM7/BFdD9Y6suyl2e66ZBIKmFCYfPU7uvpZVqUpi55qXd01pumq9guh1QlGXa93
Yj/l1Tg0R2H8GViXWe33b5QwtriuNS0CDIc2gSZ6i1GOs0Vf6vhbok93xAi3Jr39
6xGG4BjN/cQfSgTjm6LO3LkGGrD821UcjatIGsLfA1k/RdthlZDi1qi4/6VbJXsz
N0e8iSgXVrx/D2uhCMfWI40GRjKC3fe8dyNtr5+JeOQ4vKuZ/4HPGve92wWKMDkN
aRMhNPBtFTAGQevByvljr4ft8KecD07zeqorVEGpGnwtuD+sOWqUKmSznFZAhyhm
sRwfBOIpAnNahs/ZvLJS+/gl5b3PHeSOvy06xhXFEWzP/Pr1KMUERe/rekrWgQkm
89fW4FlJhFmaibkT5kfeRbFBUu7KSZBOIvtyejLAXK0tQKYEHdW4hE4SZGXtj0ZL
C7Pg36fjStpSdSho+aVpT51bSIEi3LbTqtLNF9gIOh0pDLCFaiKhUzXg3rinr9Ps
rgtGsxbscsoa/BYL9XpvDIUEWCba8KblXzZI+Mkf9NpySyrSQUCIdbRa3qcb4dkp
6NyIqo3tqd1GlhJVCM2/LnM784GhiFUJCHkzychygfTk3+wS8HxHKsNO/vtm61nd
wYF3yCyfp0wD6VneaT8FgA7np5Zn7jcFMnhJZNDphpo6ku0M/w6iWtm31ofgoll1
oTL1xeoer0j4dR9jYtk90bDB/UZp5tmWN9C6ZfchFKsaZFeqNkFF16KLRyO+KzBB
qHfOwZ89I2ugrRL9YR1uQuTi9lj+heL2pmFmWuS2kW04W010WtEBIm4lHbaB4LRm
PymLEq0E/9RI6Y9IP5U4LJi0g1ajjObgklubCAFlHhHgELuZ13cEy6rDShtEv9/f
uin3W3OlE3VGfw0mpqeBRUEI6YGSeQez8b4flyoWAcfZhkY9JrdOY/r1prirtGxt
lEAlvqNCUe1mh/kdnikkX76skvTwAeWDyseKvztgOGpoiuGDTpyqfQdqPhtvEqfk
vGgjS4QHANgWksGCdXi4PVHaibOc2Vj5EHeNNDmVpm8QBwK3IpF4VCbFw2lFirwX
`protect END_PROTECTED
