`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+/PatIQlSS/nXkYg4sce5C66LJGJDArzcWlFtkcgql9P4MopIEskQvXw1KIB/KaT
3AOYLtPe3PmhlOD/3FYC2Q6f6aitMe8/f2nLidx0Ng1p1Qx4QLy4HF5zTpVgNbjm
I2CzKvifTW2tE0YXNJ/ECuRUOYREyIE5UJP359GSgQbM1ZtNtrbf/H6W5N32FMi9
c7/fTwaNne4MxfXAhh03Hf8mkAWzotL5+gxHSuLY8vPTegRzG9GLMU8ZbW+oYPrn
3vnWDCN5To9FxeaaLsmHRFeSFJ8458HPAWaq2ssMlxA0F/SgM66i26jRTWPImJWq
2LNf3EPodTKe7B1Vt7Q+vvNhX5nvpMWqwxvapz05FDYicKShHeon/awPzF/IQZwP
oLpL8ET/ZDXDt3Qz08YON8iLHEOFmsGdSpqcpWMBTeH2dJcqDkVaJI5c3P64opiR
Yla7EisVvpegdCODI5EJUNnFKSxhpBa2QFxiDHq2ZY+DhTL7piXN6IOmgUMEMdhb
oyRrcI0uUJU1G+FiQrdSVR53/bjevM0DtHgZ/iazgdVtmSCAySCfBnq0iM3ftDWc
1awn7Czgj/uUsylDP28t6A==
`protect END_PROTECTED
