`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CqbZrfKfTuZar6WnbNnu8Ml7+3f2qua25F/QJZ56TO3GLjixCP6NVytGhJp+uva/
oRiYS5ajmYZ83WVcnbUL0g1z9b2ol3OuuyNWcQlwuxtQJMdd2Ma1RHA+x0HJHrEz
876rDJrOuIlFUfbTSaDgpFgK9wXmKSYtWYnr7JFlk6D4bbEtFm6MnhkQX/QgrNn7
9LlEt2Ig9FIFM+XortDOxeXxaOgkYppJHDcUZW1Fm0LV8IfFofIHT8FqwZALERs/
dJWNULW+kD7IxAUIbjFXn39/qfudQLNA3jT0vjtVe2xEyNuSW93xHhFTPkpnjrFP
QjFFFzlftiousvIqInEXuFqpc1OdXtjkc1NkAOasoBWB0PN2gNksLKi7XvM0pQTG
5sKduABdKlN1IlXzgSqAvbkxq1cZbRuJpr800Bk0wsiDdCOe0f+tPLEafIYygF/y
gFKU5+LdYX07wWILOloC+l4qV8JxUIshEPg6Qb8fKTCVe1yIAz7FJ6oAvWnKcnzj
tJjP1dzQ4+5u1pSJ1i0ka6Qe0delM58HHUdZk/fBFgTP4aqZc5UquICv7P2VtQRQ
nHLW3R9IoLWsVLF3FYuU5ggAuYxi0WdLSyDuRL2sAt+2rFweuqQ1MruN02U0nuYf
0fnV6HeJ0wLH/h2w4vLVq0kTxtsxIjigD0ZQCPN8W+7e2Oba3HjPaQAPYWgobuQ7
s6ZpPdan0jf3hlPtG0z50V/17WVjrwY8TGmzfVDTQG1TJmTL8DoWkqRM7dLlstym
tEWOYYMyFX0kxlvjFKtVPru6AVb+hYrpLOwBzkBRBD1FefzmCJYoev20iCxrOWf2
ADE3oGC3Qs3oYetK/ytT1ZqhHufw/N0Z+LcnTvaBIe+YDlemi5k8NIjh3wZzyzwP
ToXqb19WmkO16xlMBUILLgm7g2OAFlFI9XzX1Nt5pcQ=
`protect END_PROTECTED
