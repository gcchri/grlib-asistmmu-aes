`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTtMzhSggjM2OiKM9IlDWrGD8EjMG7dfjravTNLS5TcZFtR0u+6xnPIjqPn0/F1a
tG5F7Wr8VXKFEil1weQO82ywlwkgCpT7nRpKcZRO4HaE39rGr2DEv5pK3xMmRVYU
io9UJYENSWsV/TDaFyOoX9o48u4De5c85XfZSivSs5C7lG7BehnwVUAYDDSI26hb
hUIIwp2gyKgZYuL1OJgLQD1LU+8YtNLFtkL2yJvDyWq6Z2G3FTZaR06BrCJHBxR8
UxnQsc1wUom4LmIUXOYGtZACZSqzjTElagnEuU6ECHnZhq1sPToL6poH7wUSZoyZ
PpQpepRL0dO+HfjGIinfO8tkdlYQC18d37GOnRySPDRfOsm5NzhtCl9G5xme9C97
VaLlheDnMqsNk+6q2gJdtMvKQ8xG3W+exOS9E7xb6CQb9mTBTZZSrWIpBLaEkw3s
6IPWgqfEXtaB96/bTanyJkohRKOt4a1ZPljaLvi7hrjdn16pG6C7xyfApXQY3cXv
5xjWKU2eqZEDB5bjBcnRNnUJzouKiOhBJdwLAEAOfzpSATArnTsiQ08U3EoP/C7b
6EUWopVSQRSu4ESALZLnFEzYsi3w4vCqGBdIOKs77gCcCb8lETg5pf9PQ/6dNyQv
xK6GmUwzeyX6SsBP6pFg9bG+nIopYdz7oiEcOL0RBozhqw9t6h7eiYZfjbEufjZb
kDNzhgfo7bt6FM1bP9ZRnRjt/Bk61Nhnu2lJUI7A8b/uH54Yut85OxGnyVEKbMX6
qrNNu0xOyLY5FZxmLGRf2XHlUViBBOR5NaT0c6q/gSQ1cF6KtpmeNC1P019M5gRP
moaHBvWKSBhWcM3bryTsmqq4BImicbIR7e8e5h2uMSOroCH+AoxQRKPb6hozKMoX
8ATC4Aqp+O0LCSQQ6NmL5oi1jzpgxjl5Hup5lVC0Fa0mqP1F5KAckE8F/E4LHZgq
2JSKM5iNjo8Rn3KaF9i2B5v4PhGFcTQ3UhRI7Adzt4f9SQeDZlPXH7jrqCDGuWNf
5JcVgnBehFKhvFPo3FYitqCHuPqaeDw7CKHoFXOyOl0Hx4k8HcAKsccakTHCIsG+
CyEJEGeyQZ3M7jWa1aa9m7ix1nXGR6ULveTiwLlaQgCrP3XIIjym5NFNCdfZUfQR
aJZ3S7UffwMhF30j8j2cGIHQ4xZpcLlFJ23lL0MEiiW3Cu1nYC7tTgYzj4UxnLxI
CIqb/73UwnQUYHvzMSmoQg5VwPlOO2/TMD6yC4qqxgMaLPysfk5Km41uXIo/1Vmx
DpwBQdwcNy1bYkRBPFW1/DhXMdo0cgZ/aWXCozvF94EFGnmaJzeLB2f5Sd4htMQj
TalKrrlDhaFRIUfBaQrnqdpYJl4D7OgBukKWldy3iH2ym/DqdgM+sxS8JQslDy5N
q7HqtdPA+PBmFBKMfNzKHYoSf/pfmYrOSpp4rwjFDMnF21JLLAO8zaLkGzFa7h7s
hBewtUvBSrGLeeX0ogNvOCnXKbCnQEej7NJ2IlxE/mXYOOOBOTRoehpj+9WNytlj
zEyTgSrneyKX68u91WTBZWrnk++sUyflgyblopeV5+5f2yci5fhZsrVUQivrn1wS
gfI1/+SnOOHD+qAzB14O+xfALHkfr8yhx0byosJu0SZCLWI908roBvmck+Wge12b
9ruC8q2AH2VX3op5amKlzCAAGC0rCUcXK9Q0n4araW4YJYY9gz9i1+xDW/+o6H00
ijvMda/VzM0Artils71a4gPR4CcNJa0YFpzTsuEcP/vsqk1BfgYlBw3AvDrh8aWH
Nl5kgRmjJE8J4SLvG1ZdMl4Gy8zvIz0zPbpHP7wOvOe7KSAoTg0u+3X+jzFMHO4g
Ze5O93hmSatSZja3Gs1O0D+8ysEPaHbz65TsQkL3JSbCHLv13f1uB1A/8mkDa6AH
im7RfIArA2RjQhW5Z22v/cYRqlQWCYQY1AzYuXAljcg2rYBUgZ/noy1hoJ/7m5tO
XUycieHKIzDEeHhvqwtgzyjFdlFOrbFujswbUMzU2TCBFq2WHH0aO1n2ZrFrKyBY
78K18KtvHRoW+ncLBm7Y4BunudC3c1njhTq4Wae8M5EnEedcfvHZUhWG6GBE4O3b
cSpj/+oAFs/cD9Klsl82s4rnu/msOwi0G0mblJnlTDF5iNAgc+vusYYLiE64ZzkR
oqQtsArvIYkgFAIvzrZ9p+maarfyYx7Yj4hepPTWNzDN/UOt6K2EGPE+unhqFVuF
K8EfHpe3XpnECa3j6w4D7rs83SeiSL2rA/KN/MB1xuMZSilCRsLs312/TXOICqrn
GzkkRKJN4wloj4A3M/pkvDehk5n1dTdiUx5ZMJ+gwuOS7WtIvEtMW/d4zYMmgfoF
KVnodhXl8wqXeJXf4YA5F9zujwsS9n66QsZDS1HcEtt+wmfn4BJQtttcMEvRp6FI
SE2U/ogDsKkuXveVl9n3e3UjJs9Os4zlKMGU7/j4CgBlOOGjpLIxrUx5feXRc+dA
sOU9wnzbyUq971hZ7YOqlT1U864l6cGMbxAvEfA1ce/spYCbfTq3CgZvKdwih5MR
HtL1HlEqjmwU4aUmQZto/AJIdqgzmR/BChrfEjzvo1LAnRls2eMmHK6Cqea2EJ1Z
RYMKFMMyR0SLxcNM5hXU1l66AuAh5ml1m6n0t0nyqpmAA+xz19m44PBH14nA0Tg3
Dufwn+KSvhCeMimg6eEVk2+swlRQx5Z1NFhJFpzydWSHYFri1ZT3Lzu7NKW833e4
DhFU3+SykQBmX0xLwo+8W+DCkqhN1oKNz2pJ9O9lOYvEsY6xm8jQvIrw4kisojbt
+Z78YtXkycskNekvlprN0qblR/QgPKBR13X0t0fsX515n8LbcvxCkDxYizCWr/Az
+U/7VQ0UO5Ex+/8xeSsvLQn17uh4nb5aQwm8WM0BjG+RLuHW9mN5YIItLgQJ83ot
fmpMbiHoBm8lMhiZrvqMkFCcpf9cEKBzEW9QFG3HLiMyJmtDd5HTbvtLPX+qecWp
x25Ojttmt5wTTeojJ8FSfRQKfJAME+fcgRkFs8PAnDcwp9aOMp/WInxUGtm/gldH
VO2GKcwiD3pAeVryZK6U6YRaLhowLKuX9E3DF+UxbC2LC3Afp0zl8JdbSkT0jGjP
gOQLZGbtNYk1TeGQvBbqj5k8kc/r+lDgFc41IhzRGvgq9SqwEaXMv3mCNgdbhTEh
k2tynnjsSTNKICzZ8WKz7nSGGW5cuD5mVTV6FjQq/FZyco9YVVgiqo2Jx/eCVRqj
xoVnXW0TqSoqc/AMYTRsb/53id5yl9gkOmKl87eL3iP7577vQQNpy2RfE4pSxAJv
D/hqGA4Okf0oEpwpWGv3TPvTSuJMqb7AVMIadLQu8cs6Nz+S/qWxh7qQqTqRP4wS
LB09p/GUq4ebhLd98CpB+yqLBIdngj6rF3O/VJiyLW1B/OjJO1KaCSmV9478HLQl
jlsT2ccgyNcN3QZRpzbQk4dZsdtVT0XXvbQfqmWLW1EmPAr3hxnU0xnLqmHanMMh
7EHxWB4j1Dnyv+Hh9RxQMYx3kynzg1GjUZT2b2qFBAPWzgYARNWdfHJm1o0f0bqT
X2IK5ojzoTlrOSnwU9aVqCzAVQlxfBBEE/kVShC9x3Y4dFyR7/t6ApU4Eugpxkzk
NW+eEQ5pggI9kUuZDAMoDogmnV86OBErZRQv+EsqW06XMyacvppBH34EXQKwiJRv
SzyEFukhI+V/hsYh70wX4tgPqfH1+3pbGFnKhs1gu4mjrX4oqpGw9qSS5OHBBLP2
0OjI5HQboVnfHzkseJjwNIfeDPLHL4js584l60xeuDuUYYl92x1LHUCjvBpLuKsg
tbXzMeEZ5/QOw3SJq91LwKhVTWpQhtCUbAThlWgF7uNYShjo/mPuiIWzBnSgjlVr
3NUzpJlkd8U0A0pchalVj2rOH8LV+MlS7HE/Wm5KvnthqH8/zBWX24QXuo5XLolT
XyqIcucDWY94cPJQQqQJPcxG4gRUxne+B+zhaDUnDmp+iiPO3hEjMTakUTTvabim
TYDn1YuI83YqpDoaA7LxxuT74+TcXywfHzpwSL8xmxlaDly6plzo56eprnTi010z
OnRiw4/0InGEqttx+Lr/bLTK9oHwVuMNoZbB+4Pnl9/3ORaYqAIXSjvNjf+IWpGr
hUBNDWgHL9XYAk3C635EP/hSXfVM48Wkvq4fs+qtiXKzIpsGAtzqjG5GoClqYK1c
ZYNlo9hA2evv5x5NeVMZVeVLi6jiJuK/bIPqQW5nKJa7QFiquLngOREn1mUliPjk
AJp7n7pufnDqwbXJozgAJ9JS4P33QHX2XjPLSBi/BDC1gniz5K0htX6EFWR+2kf4
FhCdygxoVq0oPPimkrAgOOWolyc0UP3+Bv+zMYTU4TzuzPyW3qjQa+1ouHPi8/yX
/5UuNKWjpPQUjXufMafeLvLYAYe8niruCSel7VIfgCPwOQMxufqaeHV0UksjQwqp
datKi3j361njux/vUN8rYJqx5s0tiQXVDxRXMduAjHQAOlfkEhplscoqvu3YGSZK
Qypm+u8owlBDc/ju2yI3smnGEG3l9/xV5n+ESubyIvVRj3fkHSr/Wl4loWJBl0FC
GlquzjTuy/PuSTeZj5F7p5nWM92DoI4d7tC51IOFCktEnoiZscxP4++p2fMxQ0e9
HVH0Jl0OuBbkAsMRd024hJ7zPfz8Brie/7bh1B0wyoK9H6R3XhROeQFnjPGs4ker
SR4w4H+BySAtTM/ivUOCfK4BsFH+Der8G657xIg0RLYT++0U68JlWJl5KGUDIyeg
N8/XDSXO5S++QO2toBdzt/7q22BuO27Jnd7lw9mgqrg=
`protect END_PROTECTED
