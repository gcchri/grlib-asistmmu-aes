`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e+AKsL+KrM78QBboEuFn3lXA8lUy8B5EU4fRhdh09ah7wBPK6r11NoOs41SRPg2E
g0wqTqNz9xrMs8naNsMFp/2rx9m8Rm5DakaGIjy+wiG3wEfZpaMCI948X0Qr9OmR
XQEV2+YQWRrKNkHVF3wl/gvK+YW1NPIXpZFLR5Vi39yHXLouCODpVOmP29Ypn/ZL
0v83+ZRvPOpFFQ7e+jnUwwlo0F/ZAW5MmooxbvbmhOPVzkz39bXXOB6+dEP+0QmE
MzfruqVDt/KyZo4mEQ+j45n5YQWTxmwUPM5o49Io+GCDgZtRp8I8Voky+oGlnX/A
1LQOiS+cvsqF7gA3lCwK6vCHYqcrF6NLd9VYQFV1t3/etcuq8jtx0ZwCyXk8JOrP
`protect END_PROTECTED
