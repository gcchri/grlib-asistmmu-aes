`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJxrkz/AZxQuKlLj931usRMb6X1x4/Cj6zx+r0hkOAAaQSSPhSmk2MscYPIvWXkE
r2zAHI8Gm8Lg9rzR9eicwVCoFpk+8FSbLvef42/ZQnXYm5kn6WGNCpEUeLXgHDrw
Rnap8JlSonHMsHZlvjHKlc+yfUA/lrBsBOjCnmbym48OdFPDUA8ltGOgkm57yfHZ
z2/OEigV4s1rn0bXTTsXAdlqh6H9TWSxlYpgBZ6SmUiAIVCmdykqMSq8cBNw97J3
oUgHUl8iSCXdjtKREtDN7HT8bmTjVUh5ahdDsQ1W7AFbLnfPnJWVPAcs/Eu4LsOw
x4zfRlgOFbpMOWJVEcznTwk/m7lAGuy7Qr2NGamvk5Gaazn3ukPpeg3kBSkQ5+qL
qwFnxsqzHMomIUKgQREkEk23R9BwcE38/vEs+DEZzPilDtZ0SftZmeQFMFbro4Vo
FALJ2GXHrjytxmf7MYNO8SMuKgJZ0XWCxwiRTE70n3Mvki+aBuwGcbxwyESqwZEZ
V2obuO65vC5lZskNlo+3gv9liXHZTIGki/FNi/y8ahG58rFt4vqR2wadADndb0W8
brsOybP1spgnzoZJWUZf4OVqJUC47pNbkV3kE8pVkjW2IJdNPOma62g/Goh53cf9
dmqaomibtGw6LIV9vrnBtXI2v4f7HthvzTMDbq+LKCMFYMqS4wVo/ZIryKiFYwin
uEkGKOAHksdprO+ITjjlTCcbDpHUX6KH7ivtTnOevVnZgyjoAiMrgSEfAAbrk2Hk
1K5xmuWwkkeIcU61nBYHThkz3MlXuH7y6ZDcnWmTandeM5NmigiYCS+yl/q8jwTv
eFFL3Zbz3GyhBsf2mkYbVT4HZDSMYYQY7nkMmNkHGHQruDq46M8U4q2d1Rh/YuA/
V5ji+Rab4HniLBaIiYCB6IPZJGeZkUz3OM3DF0B4Xy8Zly1RU7WK9JDta8JH7n40
c2fXE/tKd+0GIxM649fyFSB8W9mmqq1qKV/3rc+vrSRASDyfVgZCxER4osS44PLR
Vmv8GkGyOIVoOH2sqt6cETW2pRGARQk0VwdBjOKnGK9Dz0mxjl8XvfEMkwPHPZI8
v/257IUkYmliOrXzPcb6FVd5rYZ4Yh95L54anBox2IxKBFoh+TejlfNFUkfLoZBw
S6t5/z6J14qYZb+WovYI7EzmhWr3D2l0XUOeCZNZfzorM0CBVgrt4jLn520Rt04O
AxqfNJcCMoiOcGc6YgbZ7zTiWcg0EQdBXsrD+Ycv37Qzv19ptwxMp7TO05PydaZK
CuASRdrLXQ2XVq5gsKjK6Y/ysFPaIoU0x9KfEjOYb37Q6ntCL0EhVXAaS+GsLGFW
K86p44J3FLJ4Z5pDwShFWnhmBP/Q2xLQw6zwN84qHOrpCO8haOktSBc7BMX/v/q8
Veli3gYKEwY4WvGiro5OKwTKwhg4ZGvopYgLj1/FZhsCpK4A/7Mp+sLbmObyCkFV
9kesMqonGr1bNerl38QRssdZpjhFlUr1oKP16ETIGEP4wRP1Re0JtxvjzufQdgdT
k4WluB/cnMjwKbXvvmf5Oj8YUQEPsitLNKUjpjbfCMsyRDqZJ+rHZ7e3rV68LdQA
sfZXTMK2HjvGIaJ92wHrMNKlwTm5rkqdiUgqJl2pvCefT+a1pNIMBow4Omt3DGw0
ESqNZZ8PAlHt2HUj609/33Jb3i+E7tIfJxyc6PY6OqUCDJn7ZmD5yRUSeXC4K+Vy
oFNSG8b4xdyi4tTaLTmYK6mWCCs4o/qQQiFdKQnnVOYWrEvppOzAhFtbax1075Gm
IvpFmD/sTkdw1c2ZV7vf3bfF+r/KFMBQKBbkwtnCeJBDGFrgTyvmtgZrpYa3PLbu
lUdNkODNsvVwVkw7HE+ndQ==
`protect END_PROTECTED
