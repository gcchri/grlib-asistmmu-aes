`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFUqYSgddaTCXFX5FUbHP6mSv+Jy2WbtAb+hf8amc5Zbul83zrWP2QqhxY5U7Bqq
JiIMI7YVDfMSeeXWFaKnvgG2fdCkPkIfKELo88cHrSyps/yNgDByCC/0tk8zybHo
EVN0HozQ5e+xUCdhqbHrX8rLpY6ZOyVbhQwZ7BUc6AkAEFvPeGI85OmveYFzDHK7
pB/Dj/MrqW9O7SHHIAGkQ6Br3NF3Lw7CX7ShHJEQqdmYrSrm0uDYMYn/8BxjUis0
Y2YISvSCFOzdVUaVRRby58ZalLPu8XjOTMV9Hm4l0ZaRt9vJSmmmF9X7PM0/hHBG
nHxYbsb/k4IV/UF0iePt6NDdr5atcon4mLu5TGI9dF3bV4o0OXz5UvPSounwdBL8
zXEIu+Kr0r6d8ouqYldyu3zhOx3RR+gzspV9v7KGj4xFQgN/js+CjKUju1twOsXM
h7CyBKRXdBTqbKqIRoaV862zbNr2JgEz3hxTFLMp7u4yYDnxBQjLN2qXhG07AZMi
vnsVqBgo0RKiZ7MkaWJimTmv2MQDCiXbWX4YyPcRR3UkA4Hgr5qHPAPfoLAjncDq
5D824o25a4LFbjbNri6UvJEWHavJrPEkPU4pToIWBj0rAyVwiSo6blSx8JyEoPOS
qF5+XS7sFOLBdFmCz82DvGKqGBGIH9RaZ05UVq0a2XhdsIiyoJr2DD95KwHOPctY
uUdyfeSgTd+WVMWtb18cQ9B9goSPV/osEXtkz+W7nJfWV52+wjMOpqkCfLb2EOg1
g+ZczANRORl86pDcbjalgAT9Xbl/EEQtU0+dcqDEOItq8AdmI7YbwD4bExwpOId4
sBh6tr+uKN9Ma6zHlNPCub3oLX0fBVSkLEIlTS8QkMg1i5D1wp14KDoobUyNQWFx
a9a21Q7bM6vxtCojBlzo8zArXpErurvLXwqgu47QFWPp7vs1Gvkj/AImo36A/ja8
cWYs8lTtmoywqCeGUnxRnjUa2pRydBb9Tky/J4/YfZnvZnqtODKZvqTHMkc4RFj3
il8Ye9B41l1dqh6cvDuHZk58O2nL03CyLvEC09t0K2U3IqJaVvFSm4WpIEvYVE2g
UMZCoLLBXyqwOQzq5LEmir/fqE3QlZFDQmKeZ1XPx1eWOUitIfLTr56vWLoAIi4t
rz/WzII0FiiofIAdCJJGjUKRWhVA4NJrFMBZtCANAiNK62F2gVHibs7acl3KMk25
Y2mU4pEGYdyBvEsZeZldyg==
`protect END_PROTECTED
