`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pWI+9yskiZSE6sak6VDXXXPpLYxuUn3267xFRXF5Vvs5Ar4fOjsOYd/sh8QsYavE
zFwzbIQmoLWp1/JpSyOqSFKQWb6FOiNDznPT5F6roCgFXk/WggeOgF2ghCOm0/Vg
/86L1KwGYhlrfJmyYMKQUvGUx/iBuA8MiPmFEYcwRNJjJa1XXKTqMmiKFTnkN4y5
kPcO51lwfWjhZoKUaDvVJY5Gj1/BCWIGM6dzNi4s1ujFNPBfXi5AFTssqcQZjxm9
kRWR+64BnyzONlXkUWDyey6MO2L6Fk8X44JpvxquuLCgUS3FLxa7Usr8N3+OPwg4
GjagWjrMLdKXCl15d1YHJ4HcIhetHAYJV9vbYCkvErTt2XVvHK/GTVqE9e1RmCz/
DQzj9lg6AkuSSYI2rUejJEach3HTp1oftb9g3TJuFIMHE3gQRbnI3hwgcfATR6lp
l55Oahkkr2YweJE1vsCagPPphb6Fi8ms0EI2Bb0B1sHSHw3TNIcK/IccSiG/2uTq
FOmSFIyYNfoJQdJ6hm/aoPKPA71ArLvv0lr4mLpiCeLYCLLpg3mPX14jhWFjk8/J
Hrrlk7zSjPQ7lumCEzMkC7YYkCwnCRnKZugdvHQSKWo=
`protect END_PROTECTED
