`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYorGhnMBVYiBDVHzkeQXtzW1eRxKmeFRZUElBICT0aajRuZhskQHj4mr+3mrme/
rTyx3xHzdymxBtSKVymS5rfkoM4ntkokduAZNuy2LanFGMn1SiI9FG6Q0hJ5LbU+
il+/tB69VSAH032XlMT3FE/kG6YjLOUrab7QGsza4lNUwprk/4cpnSMb7gtKT3ck
y1sOYX7kPLKkXB1VvXNYbHANYlwriuQYB9y6K538tNTFl8KMot4z3ZZlaZqGFsWm
J+OZbmovduSFqGzOnbO5qyxNlWMWMwADFOk/vs6fDeigKrp+Q8T9yZaq06fr2/QO
5QXbC/M3pU40VrT6LqyiRZTTouMMDJYWgKuSszdoxmbBP6KNEAXBeVAGqG8Nd14N
3W6sbLo0PHkLNFAF1HFvGX18L+vFskWO4imahpkWYgkV5o5kHv/LnrJTCav2LMkH
rlgcPlZai9YQECFxahC/fZeDb1mRba9zJFXkBT4z3/Kk1oKif7BQNKZngRI9wl6l
USyo2hEWkq4qwULeNqgSepHS49s0YeZDtC8VGQwibd+Cfc6s6Q4femcLsmVWjXLJ
n5+i/UBz1MYHSiFvNWSvPiJELteuz3YAHTKTfVKbBjYRAEUEOxoKiNM0J/9SJVgK
L1F9DBBTIO+5k2PTokThsDoBTOp/VIT1QabBPMo5FkzgnKvHZIwTln+LIUM1P3zE
ipJIkzcPjyZT1bb63hbT6k2KDKRx4EPHHJL90roNMzIOTU14xKWyhomnbaPP9pHj
g28gFyVdFMp5ULiXrpasFcMshcu5WdqSBwcHkc+zY79cdsk5AoJHp669+sAWUxPA
XDKjW12ehUYRk6mOxMQmsBfokkISh7KvMr4Z71M5zZ2Na2BJ//L8CUdtwaUqxtPO
/hLtmuqw6YzSrKRXByRC+v8tuyXYc08KhBp3Re/ue4oPKnQuONNO8cE+oW/FlYg6
bwH6z2gi5r6d/P6Gp6F7O5uBhK8tgfYvj7VejVfvLNFZfW36WRFPxMDP+wgtJOTW
HcgfsBhtXcCnOsKYDVYbKqqD4+FgN/e1VSKNRzJbdrKWisYTQsgoAjK7XFx4efOq
O2iySLGCi0S7sqdIyVii9XlMBAKELEjMQB+INMLU32PtcytybTE9FSRHes7pyVpF
ZLFkNdvAuhwGyBSBkENTTWvzDip6CoBpouoNLhKX9Q3w2psGmYO2a20oCbc+5y2w
vunHhuV19OcoEog/oU16grnP2qWnIJuhSYWIe1zsGZfDjuDlZ6iXSffYe6XPnuPb
Sogs+7aAsnbb2cB1xlzoY/ctOCu3jCiiI2r0sCRWlJv4P+VMb9sztpX9prf8XOBt
sH7HeNWcQ6A8fc5FJHiaUHCizQTAu5N10d7I6c32u26ZUVuj51XICG2fo3YUbq2T
QUJovkq8Vod5024+0kBk3FovVj3B9gWBJVzh/DOO1Rijk2nwDgiFpqevlL/JRncY
Bb0FEpl1Yb64T5I9IaD1vdbVPb6bb/hAAfif1/uEAv5ViVxOl0K+KoS0fSy/dMCh
Lra4YXn8a6hC052dp+seo4uksxmTHM9LUYJGWx91AW7S+iByOs2ByejUWU7h9hOQ
H96+iSfyS+hAHN2rYR4nem3HMkrlC5nmHWviG1bkj1RGBz9cY/RDWVmeFA18LFLK
WbQNNQ0V0jE1/9d4YLzFzo9SjuRKghOLVtCcx923IviQaI8vmot+bC9D3ae8xK9q
K3ZcLb+uTs3PS1PgVca+8u6RlDQY5zCqfhe9s71WjK3xqACsncB2A1eVse5hYwRq
/0IOazhEGbg52TMfh8Yk4X6l763DOrssUM7f9K4/eMTs7gareSW7287i/jD3yyMa
QrA0kE66uqrV5NgdS1Ai3oS7yS/ZqZc1FXXcXmyFxY7RDmY5Eyvd5+hPQPzbDY2+
ia6Hn0j6mBb9e5ppcGgCAEq19YGnUmmqC7WBH4pbNosXsz6LCZTWHPgLg4bXPcLr
DdM3lVJRJD/Wa8rIEBd3BPN08rU8PEYWSifJhYh1OCkMSeydq0xhgX1suf3nyK+5
oMVMWJv0fEOmON9WkswauBbgt3pVPUqg2jyxa+DInBPFpRLv2Bm5eQ+Vc3WEIhr2
bsMk25OwySrYDgGma8Ah4IodDS0VePvOPkR+aEZFiiHBDVKUEDpcV//S/Xk+0Ujc
D4FdkS16g5JEKOnXfv7m1TbsT84MGXaQmGUK4pf5qrKELBCj9XnYPAbhR42IjjSX
0Wu0DxmuCdNn9WmID1/Ak8akiMDnoN87SgBwH83mYLOG/j/4O7+s3nfxXMBA2Xen
hXpJzaDivGl/BCrqGfKVd7whaDLj25AWSa05+itocdbA+ngriG7X/d1eS2ZORgjT
cn/QP8UU90FDkBeIcPV6cQ+bas1emUBR/hOnCBbXQlaJn3YcF5NRwgw7Ws8b3mmv
yPLoQkYYSUcgJz6Mc/kuGxN85tiEp18hfDsbYcWdLSrEO28xUNq6j/G7qdBFW50f
dUv9RfvSt7H1Q3m2RnHSDQuDvs74dKZFjXZ7tduqthaTZXyFu8gmbi7r/RpMipus
NsF6zbatRS4Q8Ah09Kac6Q80gnPvsCjYbVMF2TnvUTc1scPSjMvAsvudEXgIdot6
yoUkZfBEoFCd9v9iARDHwyIqvvyoqHMSPMcUt7wEN0Xwz8n26NvSrox2u5iWQ7B6
6LufG5vHU7Zjft7xUpPKbceKwT6ZjOj/18NXn6i32ooMCJ2ydJ2aHSd2hFyS6/QS
FUi59tzM9zKNEtHGbyq+EWDfO8Rh9l35Jn1kd6WpvcDDgIZI11QnlkVhSY22J8PM
PZzIK8MwmAG5zvGDM2+9vfb8n/5kSRSdUjoa8naK22czO8G7V02Nwj0qWQg/12XW
9Ru4LI900Bp9PprBmxm8z4NzlgcgyR4alV+xXb1k59bInjIn9ZIs5yWnV8Au4Esc
Bh4vvsbfC9exkqjO6dFz+eSm0bS30yVaFMxAT3+Xjq9aSVwJ6nhLHVB8Mv7dZHe/
/h5EZ/cvbiXA4XL0iPz3s+e0KJjqgtfQgL45EWiDqFcvWFEqC18vz5YXe4WJCgte
U2btxJsQtcSlFOHRaEHWjEzGrUS+mAlqT5vXa9Gr1JQnfGK2aEX4zmFmqJS/msEl
GIKHjynsijJmPuQZh0hf4lilx4zX6QyTug9WSUhOzVZX67j0uJy9Y2ZMQA7fF1Nf
X4e2I8XcIMv3RRGBDDH34hGwtu05++hiSCe3tlPc0u8UhQ8ODwuvbv7IG04kK6BM
u6wjt9UwltSB4MMr7sB0FLjvPLaEXTbK7/avzyxwwskcQWV0nIN0Gef5uwnAzX1V
Nc8mfjr/PaRQVZnYgqsHCnN3n/QyzU9+H1dEfWvsmaA1YrlaHyT8arts8j3fOgF8
1wovsN5qk38HeSkkMXEuO6kbpAjOuqF0kH7WXxlmNlFQosjscBrij5v4Mxw66iLA
y9ZSl/uG2Ug641zBAZITne2UV0NoSdRA3bcKSaRJttwxcwMFktpGSryqAJ+5QdLl
faTtJZ1POpbIUdfnroaQaoRL7eImwXOphqoxl7pvIIxUEFLvqHA7mlR/S1CZR8+T
wrATfBqQJ0Nc8/kIrVI3OvNoEXoBRjYcw+HD9HYeNCMzIKe1QSuMwswnk4I5haui
fZeR9X69DZ2lbho0Kc0o7eXS9Ywk7FC3ZHlvWnZ2+k4sig495ddOHrxPzPoKC4Ys
RfkThvi1PNM9fq8d7YbfqLp0qeTsWlEPmlS9B1A199ksTKdk0HKXN3j1CPe34RFi
hvvEjKyxCBLRwfQeiSeVY3uOZUS8Uf1lWeLITp/GWWDey38WwLJ5icpRDcoangac
wG8ZWkAHv0jvcX0qDf5HQZh7aqLojg/isKOqKlst1qyYkp0QKUcNanFonyGKb9z3
X9F9rIkk3o/wz8SJJrHIaLLPEJKr9lYuSed36z5z4YmhGJYsGaMcrShMUv0Y+Rxl
qVNMuVVZ5mohzgRcInbCLLGcZ1DLFPtSi76R/S+TP5fGi/6bAxGFdpCvwBvWJ2wh
tj5kIxCEl23Mlg3eU+JJnjivykaenISQSN+WtF3V3x6w9fcVyDdJ96VhjOPTzOL+
HeQDgtNUH3iLTEAMMw051B/Yc0cgIyjHZl+1r/SmtpAmQ+FdlXQ8f+5iW8qVtU6Z
VYRBTmSt50DvrvumklTYSApC2i70nVWzjIQfDw4eYDXUZLFofoCpibuwmj8Oto21
tIH0RH4BX1frplH5/Hr0DJV0+9CLRVw/4btMAMSKlQYyFjCmrulF2uTzq53ZufZx
VdganypneMDQ1ysy5CsMaYNJ1AmG/3BI75qbFB6KOru+lETIO4e6P/3F69sj4NU9
3VYU+DKLf3LF8W6hNk0UeGWlwjc7qzlQmwJ6dWXDiRvMzwoUmYtTX+UaZztkajSX
0AEJUfvEveR0fMOFg8o6OM+VdJLKzaKp2fTOzm4NoREtsEofG+2n2MdNf50K7K37
KO1T8khL5T3TYonRRc7N7AmdcBG0OF4ixtCCfsO9OYWs0kvg1xcjUwP6zofJrTQB
4UL5l9PoMqGjhU6nT89RXFwSTzHWZKfscZ/tsuMEilwk8sOewFNUmpdLHj17d7SR
qd9YjC/Ttzw2mmividLonDrRk+K1c9Bpi7KBf9pyW5lJthQ9MApb3aAq+/cLQTUi
5Y4j+/idT2LESOTNxj1/APPs3cuW+Hp8PsEvfByTO5Gx7/p+5IkQPvj7DROl/WeD
L4VMBd4gJ391IlwfbCykkcc7r3nwwQZtv7dfY0dLbqlUfpYKIvNa7DcksiG4Ikk7
9/GZ52brLMyHBNBcEpmBPFhQMzENSnv4Jv6V5c+LNcdH0tKNvNM/LVcv2ZPbhvGk
ogLo7t89uVEgKH1bo6gfzPrIXISb9ynq/hwE3aKPh7GMjxdJESKIhuQBHllrWgx0
ultib0EGEOraAF3Ldmtg340QDwHxwBkfGhgAPoUhBaNXc2tAb3l28fAHK+5TFtcb
TNk2p5MEIjR+8JST9LaenleTJpRBLsDmpmQovdOSbjwxkvD3ZxSVpuuJGsuzArCc
0f3keHoTiGBvh6/0CfJo3xIAGWEqHk4ug7DwRQrkgP4cdl2CL2Ilxf1YaoJ7JgeS
KUIegoMoK8Z25jUPWTx5JqW5eTPskXsh5xgGM7frmnlpfc8JSEtLeIfTvsljVzgq
UsU0KZjIF+KZCXfjln5/LwMdJpd1Tn62MLQ3sGNcnUW4fEqPw8hprVp54LQ+1A5Y
ojvZADtANV24O6IZsKzxE8quMhTGo3kM1nY3D56/dYa1tO0xQMTaCq4BZhlz9qUT
5p3m1bBInpqHXdyJhrYHPo8VCQZ6YBdruoI4v+wN6YUi3qr+civKdlWigMsdlJrD
0BG5Xua2j4rju3prfSzrckpYpycxWipbX1+h+zpQxtJXypdLKkPwZ4ODQLek+3O+
vjCg8P02OUGBEzvH+DseB/ZFnh6JZVlFrg/0rAVTnNvZb5SY/UBr4Tkj5WIsCL3i
8yGvIX3/3fJdyDho5d+8QznItvHqdZFeZNIUyCJbvZ385+yb7R8Llf/6RFfOLdkH
41D4G4rFd0VfSpNSUpmPtucVZH2Z2luQjtpyZwGg5Dup8yM5O4FvRGgujW+Uk/L2
qmnQndkQ3sxwyT2mw4LCu3tQ/n+FciFLf70A46dAFRJi4hq9vQjrVJ6LMmnNjrAu
FxxgfIw7A2jO58WeToLTE+rNSgTcKKEgqwbuEmCWvjeSA998PK4l+xcZfEVyrVzB
JM7SxTGk4Kj95hOJQd2Nsiv0RnNDzYsy4MELGcprMYjE3xYrM1WNrXhDqISIdXRB
oXB8arE8mrIGz1RAL2pN0GYfqscB+hFUj5fF2QdOb+ztg26s1vf+ZREDzjr+M7yl
/GGC3eFcQ/Hkg0xab6TjiW19YeSCSDtebFdhzsrY+rkSQb+dhJ5YLmQaCtkJdKSD
gMmfzo6scd3eISe60uwJlygKiEk19zp9CiMEpw5KcxX2zPAXV4ihhv1UTpUGak3+
Si/VOrdQYzPxHSOaaaKiOP5IuxhPq0B3AD24ODdAeQTblyY13ViybLTwre4qtp4B
mH/mvq6LgdoOG84+4a3g0zaFd3W1X0AfsojOIUu15NAs019iKkE2kSaEehEyuLgL
uwKW3CsfCzCKa39rvJhHf2Xs5x0HKCOI8OEUf7IO9CwDOqeq3Svjqs3tqqlokWr0
BmyF3Htq2g/h0BhU9RfDdnQKOHPxtRZexZtcyvCUxTl2dhlUTBspckU6q7M289me
f3R+40Z4rJCTR3y0LZgvzOBBE+gepMZMGpKEgLBSDcabzbwxzbFzltrxeTPqCg1I
WAZAU5lQp2WvFVcZrSe5mCLavNy19bC0ZJFZlfao6mmkuUHlc48Sho6qcDx82tZE
yh9LOgRplzW4Ngo3aO3F8QFAquUtSHz2mUcAglLXX1kXpqZUxV3nnzD5tX3S0ZtS
6oo1xKUMTUg6IsaU1y8aRJzpF1/tSYShLYh0tdvjYKzg0NtIoBD94CICQFC0z0j0
WVKowKunBcK7a1zPB+5e6ZNYue6oCFYv+BFXFt0Stufh+30atfR4WrykSmjYz3rV
rNVCcP2WRMuCUXx4VX0UxQwzV5mrf6/WEf8R2xZOTJeD5VhceAto0n7IOzSYyNMo
jmDaqNTNdgP7t109qfb9nA93MkivXXzQEzn/Rvj9s1j5inldUx55SwClrFh0mqbb
NosZ0f4GyW6lHbiJ+9LUEaS1HMAGG+U6Vg/rKRmtPJpSs2WoS77t+ehnaxe7vwoV
JAZx8bU2VpUGLX+NQaWlSQ6d2Szq3aFwuTwxGZG9CjM+ZLwhXU9++GbTRXg7zIQP
Um8y4UzlsYJzISkoOKN4cVeGXJudXeD15Wq/bzJwIzdj79Xl5eoHL2dv10z//umj
PfKcbSE+P8yB3SZIyBY+hSl34M4VfiHA5uXhZuKU+ImTTgIp8R8Ie/v5JpKNOwhx
l8YM8C09Qn8VzO+7AnZk5PbIRG/gCPmRNstLDfLP1dPL2GKzhvwGmcILnQly0hQV
7VKNAQfbKtjr04Cz3OfgUf3frls7U54PW3P2M6Ip2euQMY2lK/4/z4RfgUZIuRhn
DA+koCDnYNYnhnvxK/t5qy0Po6yBHkNavBAqapXo5GS0tghTDVRTupKkcJLNAmza
BDE/icI/eV5ZZE5LucW1R0AXuZyMkiwsLXJXSU5oPwQJj7ZcxMYn43pZ7VGKjB6Q
N+ThYwjp5V88fZk9BPqNXmBe7DmuleRhWWuvlRwIrAIlk1dWrdEcLKnuNB2IbI3+
ohhlcQLL5Ou/M8AMsZ2FvmGUSTAtNCo1nDS3DRv0ZBVbYl+g6smQfpMSINFEUcWE
IrsU1SCplX4+etAaDVpH1m4tfFBGDudcHnyjiMnt7rB102Ln9xykBkiQesBnl+oZ
WB5VmhFqemvQNyR2LRBx6AEJ/2e8BumXZ6EttSRmglZPqL1hMam0B+bBETwViRED
SRTfkQeY+ZKp0Z9x670wj4qXEglcuT74QbH8VpwPegsMDh1PnRiAWWL2seodAtjb
IQh2+9+tBIsaCt1kw+UwkrGFmIItvx5kkcftk9qGjHpCC1/qgbuvNJA7FkycauNq
7KEmZrAsdqHUusVSsPbkXcZ36e35qOIL+9tAmMlguXAoGg2fpdzPo/ws16GEYuF+
JUtjGln+dG/rEL3lX9Ge2Q2uUCfSUWIOPWgVPuYlItNe2PdBkwUV3MoPdv8hpPAp
FFCNzOXUKvCqS6cezK6ebOAy1iAn6gkbRaefRnuSzsHdYFraIzgcK/0298fcNdH2
fhT1VTQ4ra+sfl9I+om9vlt8/dTahc+kW4EUiL8iXjcrhEYVGcwGEIEmls37NwQj
3mKKzBbyetjGoOdQNDXZJBv/VfsC3ivd2UMWK0L3Vk2Jfiodvxl22wMHu92Ii4ME
1h9rGRkTiORyllBZVPiqUzCFr21fhF021PvKzANB0PoyA6zcr1ch+7TwKwsGRrwR
rd3tUjB5JrQWL323IZuq2M5jBAaiQjQMabh6uIt0g+xknN5dHg47y8eeNhVQkVQt
PrSACzGX8sKsJvnG2mFb3Z6FOfKhUrJu9xynvFs5IQBNtrQVqPjqKbmaRdbARL9h
r7484fFUOsBvQSJuJxyTNtK4BNI5XcAhe5PMSJUUxITnjuVid0/AaCL5cR+RMcCP
c38/KQLHaQAjGhZmYC3cV+7mm2WFlphHh3J6GkIP+yc85UB/3xej7aqK0GYVdARg
VQvEp/0cJjcQ2IZu6ezDncYoceNxQbFNN22eFAtUtoLiIuCTdm6AxyhwIAL0BBxP
5WF8XGllaJJk+KKxl3JnAKsieYJo3aWeAMiJl+cqrYPew0y8BzvN7z0+7n0Zbgzm
m4pf+j6Ml+kpOJaN/U0O1h4jvhZzepRc1ai6WoGrf/YqngixjSO0QBFoZwBR0rPS
XarPn8Z7IIzlAFQ/unej3evKLLeAfNbBYK5KcQAMvph6hylzoevMOGV1qjOfdzJj
6DmyxnVnfVjIZb2Fpdyc+IfnP8kOv4xSUKUIET8SQdvxGFCqaLxOxmGi4JnljwZl
fvwtXxomXgBr60IoP1djCfc4kKsH0hOJcB6g6iQTFPQYgLq+3XPjsS5aoIGqT2fb
dym+WXTZZXge6YIun1nF1+IlKBf5hrNZGYs6T7wbMDZ8egM9ICTbJkNDJVKOIWrj
uALsv4zevM4U8+c76+YNMXPVGAmRsMdSroryh6e4nu+jAA2jcbPFO5vFpXZih90h
n5i4ZIGEOVPCnTYeSOVC3SHMDAth9rDKMo7ky7DfRnodnA/Wm+CCbzfMGZ6X5gP5
APFFcEr6wVm+vt/4HHiqyhtxWhMAX+GKuafM/+k5ttJO0cZVEzkvvriTGZ2hViNr
h3C9nkcrgEa4f6ntA5OxuZigmqS5egxrlcuy9JPTj6OWw7WiTzD06umfBekKsdR2
xkDArrjq9YgMx2TN6lNwe75T7WzFdreW5ZUg1BFr4kg/kOqstCf5hoer5UVuYC+L
MUTM81+WxTn1Chvb7eJhdjaAgM/ZfnXhZBIZ3MVdjA3GEw/DBVYY10/SF8iF7ZcE
FEmYlla0hohsR6EsCL0i3V//+sUyIILtpQtSFQWxr0P3UXsU1VcQXThkCN0z8gyp
7A0xIqlWFhcwygqTXdNk8Qgfogd2EDdyHrQlyItoJwCiHeV20PqNSlP5BnTDOdSc
ZMbu2G1BoGOiw0nCs+2mObq4121Cn5iuJRqlWYKqZcdyZUS944VOsW0VPZrrkC1G
5jvff/6D07pmM4ltsu359DF2NdDy+cN3fuAf67xJNF7+hlCH5pWiGaK2ysd3hWe5
4t8+hvemLhfL4I/tWFtFG2B2K+fwfqMTy+S87jvn+wuQMx1ey0n4YnJXouEqWTtd
03/4lYZJ5X7TRoH6irY5zVghURJCu3+CwN3qEEqsWsCiKPKgXMcfFuYwLvPN8+6r
NQjOELV4V8FkyAkShBZn9JmwkeyV+6TKW6O9UiufF7bhiOoe504U13t5GQtSFuoy
WZbn0tOnGk8TOLwfNMfAo1aQGljZDn9CRIjuy8+rHG7G4KikIu/noutyfny5Hpeu
1OBOnnHFVLKevUeMfcPUja97easnXLFSLBfwSTJGHqB5YbS86RQCETzBAw4nzE0E
DXOfMVvrfemIwQymhvnOMb9CF3MbViSlEHWisa9tXRnFF4/+jsfduwPP4figLRrS
S8YEJfrEh3AJENs3erm7e14pC9TzNips2K4aHvatrqWrg5iEQh/pbEwBCCoKM5pp
`protect END_PROTECTED
