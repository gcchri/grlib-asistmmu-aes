`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZJQmff9BQ5hToS0VREB08wGrnglJHtpHaOox5q2cy4jDzLy0Dk7qbauXUiht+Jn
Vb+JOIPbJse2ALIx8ssJ4H/Jx00VB+AtkaalHlDIHCHfJQqH8Hcla5dkUWH91nea
d65L6D+j681mKjbizF5u8Idsft7cM/ghpomqYbzB6uJH30hjS4i4ICXnYa0YTxT6
Wv0OscyMkfkuXG2rzUlVdecVcMNss9nqZvA0TVdrJBPhbMzHRDMu2j2MmeE5kWGi
dXnkbBo7DCkoUmdnUc3Mq1BxV8EskSfhZPw7rDFtK96FdTVm3PeeajSPpJD9Y+39
BH3YvsSrvYl8gJHlnCQiTMK1J5WffhLZZ+muEmWrND0wyAfrVfT1ViFvjk19HmQb
TqBu37GOCnpWL5xCX8lqUjqecPIUsz85bBoHe3Q8EADOxv8t99orVVwZxpIdosb0
`protect END_PROTECTED
