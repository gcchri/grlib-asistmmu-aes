`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHwtxVvRXa6V+s7ckJnmST1a3D00hMr2VjAd1z1pOe3sQ3xHuCDflUoylyQTmRYC
36gG8yWPgJrFz1NCJBNEDOTkIjb4V/yd4eHxE0WuIOqNWNFiSf8I5VP54ihEZEeE
XyQC+KM+bOitxufTtzIgags1AvGteXnqbL3qKrn6symN+mW+YX2Cq7wtTVU37xZQ
nso6pudYOO/MWLMeMv/twB1ey3PC8vSFXoZcqBfYMzhR/l57o04veJZaJMjSsjs2
6KcjprgXAXvPWQMipZrCzr/3cMWqlMETeng5DcqwLWU6F2E0CJefL3bhBIM/ggVW
OiLSwR58dGbkL4K6YgC8nlgnRD9FgxYaESQNp3ZLEYjeHiz+8Q4+eocqg7SgeYyS
08KVMQIlLv38kgfdTlEicOTI8SDtv2Vq6vaRGMQznwD13rfK6Ni+c44xC1rLYMsY
PxuJ2WYsLx5bgGxhWR+V/z4yziQcM0RA93Bas5PjrhCocN3htTR5v68J5jlALfNd
E+8JXInuXTAmq+umYTtwUgRRsV8YYO4UQ+G6dZJGQYQVdMsdcntV3ch+STpStJiw
WuIqH5HgrDyX3pftDA02PWer1kWlFAxFYbsC6SQlRsyKug5XfZeCmuHCUVMZuWXv
KkS9/rSYCI20dEWC/SOzFQ==
`protect END_PROTECTED
