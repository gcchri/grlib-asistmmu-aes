`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bg6nitVpn31VXHXzdGUmcO7vDygq3Ky8SpafCegOeZHrMEXIqo4GdfwJyCAdLpci
9YUMMqRraLRjXWdDuytC1wHyUtonKhRoISYBu39qmStbcTvowHEVjU7F0FR0XKGG
oYzDvv1T9j2uPp4tayo4Yo9D0V/AbhXlNLkl8+RqbwrXQkJSCW5P6JELbvmPYD/t
3Eqn02eYq3mYE9izfv0XyLMtCII+bQuXLjfk7Y6stpZkRSmgSMlgzBFQr7onfTlr
CEP9xo7JbkMazb3kAdKuHfUAblaLu4ch5QXXqfTXE+9hM24h7uOJMCaKifJPHfbQ
QYrBCztRNkDCsSEHQDB7yVJeYtP1ym3UWATdLm+RRDZZ4JYRr1KD58+Pha3mBp0P
WroheIMfB7klNGXOjvdrA+ouflkuYrAMws5IyQQhVdmR5B+OwLsWi2XAsLzrrup8
doTCtaHQ7y60PwfBHT2kLlTYRcyfBR8+Z5mIOZj3nAPPZOKBSEJf2C7Zaqf3atfT
yq9WxiYycQVQEPA+wS6uwhUdcfqpIqD2fWUvWAtFNo0=
`protect END_PROTECTED
