`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
urJAAlR052VXleV3UL3JjyHYkJ7HutEfq0b87k3EgsatZ3+8e4uzW56ljOTW9Srt
3XK0KlKMQfUkQ1hsZYZzawwDhSrGf3AehWVFGAZHGqrW2/D1qcdXMYht1nrt5JlB
ZzkzAbqGLe75w73rJ+FbHGUtRUCIYpVFtAyMhmQqNx5a7NK5DjQRbEC0oZMk4njW
RE/1qtzOVPxRxixpxMehirvF7l0jw2MgHfVOe/qRRuqTuoOEj2LvyapVOy2X++H7
u4Z5fpt1QvWUfLsZaUGZX3dIO6vSOQwUETkDgZ4Av00kLlw/RLNROuPET+emIIQM
sgBq+5slgTOBeKCBLHw3+dbCjJwlp8MOVCJkQwNjvu3qX3P4PGtPPUZ8MNq85MUT
v1VawNCIKy5i78q+M7SEv8pt4jGFrsjbhmvkG41vqRZzDE2xRq5IMRW9D7ZMkljH
BVo4PumEt9SctmDSY8WzVreQfstjY0IXjWKTjYBFFBVgqwMLKmTG4J8s6Cp0WGTM
JJIULxma7/ZRriQwBKkwpxsNf+4b+eULQNBIpM5udrO9VybGxDevIMuuPHvF7tH9
ngbukPBsUuDtfOV3F/CNVxKgsozO+skK8X7RDb7e31HBsXBUQ4TLdpLCFjPYP8D/
2tRYrlmwYrGJCPr3CvK95uiGRFuc3Vd1oun6ArHNnrf8RAoFkaUpoCGfIvhdntVp
aL8FsvsMtuuX2WCAxZwQm+vZtup3BdCqHkvXEqontB7ilWeCG9BSNYXTiMvQqHfy
aVHwRMFFcjvvceBEM0MIoB70FIu+EtgOoIxywOY56XHSa1PLGRetVkl0cr1dB/Vp
FhtiaZ2wIx5YOXRnFO3nCo+jH/AGg6jZzBi7SDS6h4YQttwcRc96ge2gVpiPXAfu
c0LNcGcBDVSyOkoKEeh/gkSVi553sOl4IWZAKjEyPGZKrE7vaslNPRYaVcvye2E9
+7w7RnGKscHwxrde0qv1TlJQ7CuHLY5fB5Z8xY9AnzeyhksIbZLQUvqAr+O8qCWj
8RUgHSH5AxU9H3j9rvd19i6G0WA7Krlu/H+F7XrabWnPk+ZmSZKhBkeZWAc4cXK0
z8TmUeEGg69v2AUn2AVugBS0TJ19JDui4JWKh/riIEW5IwqzNNbsOm4FjtmtDsUb
WpZKVD3cFMjIqgCMMFsk7l035Z1hmiMg+XS7Mvi+jcO/G+TKMnv0XOotOViXB1mT
HsrNOke3dbB/vFMvBOpou0vhEQtG+2mKB8pG3Nam36NiEif6/5UNMs6Cq4mLtUDe
u3MD5zuCMJxSOox3kVEJpq77i8lAQrVdRWNvQb9kCiqb9GbNqZRYBw4/Cdfg5DIP
5IuPDSsTnprp0EBByJB37CKJS1H6VDGPCh4IxpMiQEPuz3yHvhHUVxQvZaTDhT9c
lKQTr/nVF1AkWZPkYYYWtY5we1mK2pgve5s0sJzUe66c1SSN0+RtzDoYjnA2QgOb
5aJ4mJTmziW3UcV1TYDurCLEAlZ42wSw9yDvd78Kn6TaQvWwR4xlzjWU25uF//7t
Z4h4DZAGG8LrXgiNOBPX0s1L07iH1bFVaD6tKYgeoMi8MIkXreTePLf50yn2sGdx
6cQQhKg4L1xJtmFZ/xcR40W1W/eeEIhAENuRdk5IyanwFmkjOAAqzmvjmSCLJCuy
Yq3BWszKXJeDiYFFEthBLj9aoCiS9vNc6HxhxHRPOCFMa4geAjxTlMJdiw9QETY8
P9fWQb0+Hh3qBT/RsI0elOGgPd6vBWHjD/jPMSdRaoj4fIQ4MGVxBhwNwj5cPzM5
ncnniUwBfsLvMH4iniyz7XekeFKUMTFw4oPyoej5uJwm1Mp9kFOc8pRO8K5UbMHS
suQ6xg9fjI0nqAFE9ZMH6vPXJBoKfyQjgJmtv5CR1+OxfWoYDSibjwTLPVNdcVz1
Bmo1fvkhxZfO4QUNv1/v7547fYD7Jz+/e0qPGyJI2RlPk7lLm+crKPoFgGN5wfD1
s5Mz8sJjvfeg0hDR6nZ5s0X4IcSMe2NPOfurEWGsRMijIPaJv9Xb1vbCLoCw+ybj
O09b4MzfXYuv/hKt4qd00NBkF2J3xeAVXGSe3yX8GATeG4x/2hsD0Yvs5yPe6/gt
KnuboqJBOewrJNBoaYEUWcmvTDhxLosPfdU7SgVJRNA=
`protect END_PROTECTED
