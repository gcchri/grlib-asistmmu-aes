`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GcMuzCXeP62KJxgZCgVerawcPdmCpNvFoMpjIg/pABPRsg+cgm0osQa2UELDb30V
vW5IS2e1iRujAjjjGoLkec7cJ8sXfim138B4VfsZrjciqeIVMA+6n5YXIr/UC6nr
4GhqtQEmSh/qyXcZ/+PKDo+8W3MEzvo9bKMN1WfUE+1qdovpqT1kZV0QBxH3K5pC
YV6x7v3ri1Q4ZiDPWV5UrW3EuBPCy1svVL5MXMYTMrqCcXvTwa6tqTysJBbGKVnw
XJ/8gzeMs20AKX3C68AzjVbUGyMJvUna3/VkzbOXkqYCbgQCiUHSUbhoyzyXM5pw
F+0BMwf/W1q3x0yge96Qk4uxCv3AlvpAvoT5o/pX6IK3Yuh7sih/2xjkmQW5Y5kJ
OoJqCvSDEQIpz4oGYFH8WP+hr8nRwnsUeb3Pi9m/ShI7F4d1eqYhwmMcCqJdgiKk
Oos/ulKwFF65cxylzGGlXRd4IYXNbvZDou5oBkD7sABc3s4C8Scl0gB6l6RK+B3U
XoO0U9UnHVNKG5hSwj+LsIQug0Ggyl2YTYzz4Wtb9qBywpLKJUsFghsl3cnVmt/b
7EwhFkTvrjypEaN0zhbCcJRwSCntJL16dPTJTixjBCsS74tRRfHmzkSvx4E9GopJ
prZepkwKin8u7OkUU5PClw==
`protect END_PROTECTED
