`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i8bjxRmW0aOc7gEEHPIfIXRgi995zxYKQ7xdDF8w4wxE65qojeLKt6xIPPmExQXI
I3xZXd88bMAqes5qnAY1aNqTk0iUUDy2umZHaBEdbQbS9m++Wr+NWaPP39Os1I6h
sO9is/D3bE+o8KT9Wto9RFGwFk60wCUi3af8gDdKio8lzDWM6Nlh5wp3HUiDCmCg
pLFQBBmJCTpk63sgCOR249dml1hgyCzfT6adxg93veO4XqAUu8nicmAYZmAQaI6g
oR9agSgbhOKiX7sWpoi0hLV/TSEG1sMMmrObX26QXTWJTGbPY3Gd3Q0Yt81UP+uH
g/EpTS4kxGgrTmMM8o23CyTTSIi/KIe/etsd4Lzq/gRipEcYypTbmS4wBbuhsZ4V
/qvyJND+5JwcrT6b0wkFTa1tdObrLZjEyU6qcTo071q/B3MsU3br4hkBitLSWo09
4lhnrHIp7gCjeWx1Sptl6hpuCb23tQI5VlaMQy4A88O1m6X8scZ+aZQrv0qTZLXo
LYjapL/CFeIGY1QMAFwojYwakTVj26mAbo9naywd8O4OM7MbFJFfzdJmRs6GTi2p
sXMZm+vk4u902UV+Dnvskq4591AfiXyTz9DNY8+Movflw9efHgBtk2O/8ttJAHLA
jISrxxuH3KM1GnLj572JcfhswbiFTYUXNoQGmVbDLEYrRXkxq9LiY59r8WBeSacU
74kSUcf6hkdju2Q5uu14MNxu36uwLbvd5l0FTaBMrw+yJkqciOQIlEYrCq/wuEhA
xQklaS69Tw0FedbD6mqtVSXzlMSt3rG+75fQgxm2wEk1gqLQWhlRT788B2y7eik9
u3c6nOo2/2TrOcP3FsTZlqNfBSMGS2hxbZJzt4Q+0yAzwKIiUmr3X8K3GWkX6OhL
DP8I9gyTKRBBtWkvrzBv0XC8uCaa9/Y8wBKqVNdMKMxGLiRm0bMeJs6wPFKpLz6r
UiwWkFwnMJUKoqllPFarAA==
`protect END_PROTECTED
