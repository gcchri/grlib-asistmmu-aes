`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKNyWOh19VmU6MfCqGzn+Z3Vhll1/vqs+Od49MLejMPzpGDMjmSe19RmlB6ewhhz
jJ0F2fBLQtgl2DLwb0WZPC5PqFwZQ6EEJBKj2YunEg03o/mmDBMLoX8Q2EaqbCE5
ueOicdxAmHwgBFBWV6gUbCLKQOqI16KAst7oXiIDYY+pgeUTiO+1Y2WUOgQOIpyp
YphdG07u8I+R9W3zqHWTYKMNYKk2XLwQVyoYv+0Mwz2ogD2Afw9EJtRxj92u5//X
4Q5wKyLjB3i65BnMf1zoeKa4klTH77ldR/tMly0PfV7wWCvtr7BsO6LjoifUlw/v
Py1KISLZi2BV68T5VO/RKZ4wmDFie1CNK8ct1gU6+wLLnoJLkg72cQ9GTz1bzmqI
OSTz/42VQ3d3opHR1N5h8Q==
`protect END_PROTECTED
