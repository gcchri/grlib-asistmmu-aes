`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2g2KKUlqjSYht9hEmsNCxut6oUzftuKynmU6TfeHkXtgnb+iml2XG495WMiAyGJ
1QZVGY2elnZ9JL30gxqKA4HXt2JnWaQ2HPpsH0oLFEBhw7RcBkqBHgxaURAMQmOH
zW//zMC+cZaYLd9MFsIDX6s1YtEShVfY1oBbDl1LTDhxiLcm84PmuJlj2lD6oOmn
M+ii3TwgSywQpDTxxVLvTSdzUh9L1zCiagnFTSzY6LEekr3ar+pkVoZtvzBeDiYC
ZpU4ndfaodeyaMvXn9Wcbs5I7ETHcjrz1V1I5naKsoWns3RGuIlZMpj7uMESzout
B2RVHgeZCebZdbbyPNG1QfdmAUBs3//CArZ0XLA+5m0qI3qbbmvREQ4Ql4hTl00c
atGCatH/DrvHwvOiICmDBPBS47GBKW9pxNqVN+d3GopwwTVrE1UR1wB5Q3ZI9j9B
OwT4SXgwgU8eh2BXnbTYE7ydLtD4tXgydav0MC8yLWNYXTo80RYZHq/SNMHUtSb/
dk7DQMym+7oEhNcqf9SYM5AKQeK0TtZwPfGZ/NyXDzr3rQwQOyDSDa6hKh5vqzUd
hfpXbW66aIsvOD8JDvbM4tTe+U4a5KBO27jzgrHmH1+ViVR/7YyQ6WDNse72Byj7
knEynGFXHNCNMml/ddxnRhVpxYACX5dT+V2zcukg9KqD6suB4SokPlpREpMvAajF
tC5iVhX6IXKVDuZuctdUAGX1BICWWs5+ji/nZjPkz/LOuUk/TzAXXGTn/DUB/LF8
yKrxCvIG0LDRegIfkP12ZBWvngaBRILOPJP89HXV5zBUyrl4rhc1vTkvdQXV/Vry
RkRisrb+V6rSZgDQf70+WmX5ms8Af1QZHrMz52Biqx0YzKl9qA05IxJbCjEUWnrz
PE75GOMqJBJEsBTB1Cktl39Qx8PO0HGxnbMmxafIDnOHWmW6a3XJRul4BckAuI3Q
vAPjCoE370/jaPJBVGrlHN4FLsdUszs1HuLGU89wpCAMDWiFF/lxIJtBNOm9DkZq
TFVYPpGvahj44AMxYAg+vlOFvfTJS8vBG7VAoIAqfr6mmg8MePhsEEnIxi3mqRu3
9r8tzrSsyZQDgF5bp7FKlh7IPsBZ19YPtUtSaa0rBJXqt/LS1eFxU9xmAUGArBUD
0XQh1czC0KX6sBeAw/ZIBg==
`protect END_PROTECTED
