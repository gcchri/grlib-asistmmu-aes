`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/fkEZsfB4bkOXbLze39rLWRVFnN4c1jEGi7sMyMYSwPfgwh6UW/yWrxX06t++DI
Q3T3IuK7wn5z03GnUGfWKbuxelPD+5otulVtFcmi0retcH7lNkVMmJJ2ra1dRTRg
WExMbezeMd2D4jogMTlyWs72rpkK725IIxVyPsiOyOgo3uFB4ndUgVS12Cd2KiRP
VwlrTWml3QF/9UejWOELFzsaMQXScwC5IOBiqVvx3323PxKjqG5WFiX8JFNLB0wF
nhW4Hefr1N07HZMeskkt6vG7jcGk2//dNNe/6jQ3OlcY1a34Dlme5fC9wVEYKsky
+zNQlmX1CLvDvWvGumUanSD+HBCqMOnJZ3yrGQClPRjrIQAsz37sNFBun7F2aBm/
kwkzknDevFHiLNIfW2i63VQOker2oWyB+zh92lF2U/J4xp7EIQu2+EW1YYlcr6s2
TkQ+BOTqwfRCN/zShSBIKDo+UFHgkJ06Bg8Ze01BrHM=
`protect END_PROTECTED
