`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LScQ0Y0v/blzBxzcT5lcMccqc1h+kG5TJslqR79Xid883FNxITK5J1MZPb8J/4c+
31v8441Ura90uxJja42CkH/q6R4y95IAcPfk941/WcrRKhCszmkLY5l88ErXhDE8
owHG2MjcgFPIIWH6Ab0rhM3RRJjERTcpdfPdP/rM2WzTjCVJsBLGnf2z8wR/1FOi
vlzQ7xROfPKAaBbis7GWL78ZXVSsIW7Kdmy4E/+rSa2Cs6Od7RV9hqZlBw8jT5+W
4ezo9orHvhiceKOKmTdgUWXw18K309A6B+D0U+UAYBuIzfEVRFc3mOTSyn9WQXl5
j/G90Y+wvUGU1/+di3yC3g==
`protect END_PROTECTED
