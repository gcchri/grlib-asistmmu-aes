`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hs9hXm6hRQYbtYroZnx98Zw9DLoxsqKKH/fLtO5TeiDU7XSf2qRqKrtRCmQiitE/
a4ZvR8Kv+Bsy69xcOfAGXqfXcc5oJHAB/1lckJPt7PJPGsjikPaAeWN59BA38/eP
1UP0FpzyAYK/qdBeK7clMNv66aLiLIDfplTKwjPUVfPBuIxtoX8eck5LjJr5/bV4
gd+EhR2qZHyugvb9IjbXV9S8wpcmMthufLZaUrBtMfC8zUh7zmcQnre0rSDed2ai
OBdM/pUNNB5rWIX1h4qu9TSUVOHH5lyO7b4n5ey2QaTEN3DgIIY4QworlgGnGcO7
bSZjxp/BJTkohWvdG1VjXMP3emcy7s1bwHsCGW4Yb52yRmBYRyLqHNFF91/8q5Kk
q3ZbfltgmYt4CeJJLKxPnVgRTOh1VgQ6LExwa1bBpAbbS5GVT3y+hDbv+gBMyZUm
lezkWZmNtLRQOumP5hGXLdX+lES/C0Q3I9h/mdOjp3uFzoNMWysgw8Tl0MehO/Z/
`protect END_PROTECTED
