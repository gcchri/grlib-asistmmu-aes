`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ARZ9f7BxzVdNIpJ9T1XJlgoYauW6MqVZcNnYQNfO6AFRXKhVc0dwJkatYmDUyJ4C
FoSdjfPZEEPuDCLxV1H1yUpgSsPiGFscOVumbxt5rIqoy9l54VGePzyafscGDhYE
mf57/AJlDWgYeC0lKqC547fNFz7lYNM1pCTthOP6B1MrCMucMxCyzRTBbrcw6Pca
yTAZfs/t91rUUaB+Ezzf7giPE1I2eET/37BaqXIUaNpLJBFBBf1RN6MTHDivCfLH
4gnsLIeUD2t6NiWUXD9VkK4jA++7c81iKZSVgS4b18+XOhBs1BOG5yNs18c2xxVn
P/IReRW+V2RNiAKEFprClxjl0nblCG+GG8XvNPU2nn6f2brju9HmvOrdOhdVAoml
jJO0LBiIiQwJZf8xQwq+4dNkMtoB5BjJTt9FgF1nIISwqfHDAjHK5C8ZA75BLDeR
`protect END_PROTECTED
