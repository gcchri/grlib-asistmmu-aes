`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1cxrxXSgkBZ8w9DE7Rse9ydrAIwO+vRJpVLQXjTy2zkRh4TteM0pOZyTfM667yT
eIy1tbM9UcKXHKCwYA6GrLb2vM4iEg7zDhL9YFMSGqY4H5O9/F0NMZrzMNmgSDVC
27suZ3djDZsZ8UGpqER2agh9L/AvSpwdHfOjREb7mJfQhdZX+rNx219JbF3+PF6x
j5s2ucO50JhuiKneYv+GkFyw7RByRhvs8eH+nhX3CVME4C273en8vMdqCCOs8+yx
xDp8dNOlcbV+qoiJ0PmPJvBBFxvsqaTTeFzLOdFnViQrYgR7PTUFDR53Kh3o7laa
DgyLkUh62BjbxkbtIx0C7gYbmopT+qKJgeA5ums+Cz/ywm/YXrvYrzov6AAtNNF2
bdRjh6Aj5YshUGVbL5prs1E5ByOXItColp4c6FpOvrQ=
`protect END_PROTECTED
