`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jKi8iA27sVMefzoh3+duiDKwJec22EiHO1uckxJ/Bki045lcngNod4xrR36YvwT1
7G2RUBZ4ISYF0Y2UHZLV58o8hESnfJtnueo4Y7jgVoAb76mg9Zzwx8kUkBH3Voi/
QXLdPR/fARZqIEpSU4O7Cc30ErDnYoTlO8/2CsVPbE9+jwZSlXKymQtJGLrSKxoE
iD66h3Sgn9jWqrTGcb1eYonR16RkGtTiewGfA88biGJdC+QuTm7R6ZNJ5k0dxWAd
d0/4baAhwGiMkEvcybSYj1sf2JWNjRfQ+c9Ph87BMkqBKy/t18pJhHzxZYu6PK2o
N8273AX5XFte92AlRfuienRb4Vk+whadwlvEXF7QHFOCCvBpDV448Ok5mIiBCOtn
bhV1JWWen5zlDQCzRUv7QS9ZEy+2jf3MuQKjBePLiMJkCtWyJmtHgVawb8xrl0Nm
pP+J29S6ag5kx9mo37cig/+BNDYnBV9s0BInMNAS31I=
`protect END_PROTECTED
