`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ogSRPT3XQkf9TSO0OqNIAcsv4S7JYMeDy9cAt7G/HIH8Kg1FTV7eCWyJi/J2yooN
3Fz8JmBYZmxvhIMl3m6kPmTBOKe6ZQ3qb2oEom1UurVQvnq3dcye77hhir2WLTGP
izSf10IB8qiQxkgF8vdIEdAW0J0oR6AP2908sjdmjzIdigwIyzK3hJHkeSllg8/w
0Es+uiZCbdXhOk8dpZ/QX+co87EbI+FTmxQnmpTVx/f600vgLbCB9B3NBg1hOXL+
`protect END_PROTECTED
