`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2A4/MCfzxQ7SQT0arTrcScLWFhtZBMCTP3P+4Kr/GHn1wPkyJPwMqvKOg0kcF8c
kSLvAWdLyBA2JAvbxtMx8WkRUmWr1POS8hYAyFpVaPC+mQzITdJ24XxaL4/6Rtd2
6pMxGnONeOeX5cIT9imcOKDzRHRVHUrdUIDS2f9cUhezaKuR8OX3NlZ41OdHh4/9
qhUlxVG6wxiYWwXgeErRqy7sOEh0ShxpVRxbU6hgm4JHc7wa23N4acPwowIhcNdU
PPkXr7b239rin3F83WoQAfd667V52uiywasG/f7dGNy2v2u/wpcbZSSo6LbfDJnu
tOL9FXg1elBX+R2NlLQtv5nEMTsUL4FN3zU/CqxPMDVKTe6EczfxdWnBSbA3hKP6
KMYDOkT7JGTTJ9JN3KtdP/tW34UJFwCEPMq4ix0CiVvK1Jy2Rk1COlAQXz58LnfI
`protect END_PROTECTED
