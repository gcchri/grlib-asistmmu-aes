`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wWhC2HmHcZQpjHWqaZD7heF8Y9iFp6IUskNnzFQ4hoiiQ1ykJGlcRhVgQNtyHzrw
HZg4WbO+b0aMbm2pPvWvCBiq7yYWc+hoe6UYJnOd+8v3IAb8OMmrFZ5AYBYN9YIQ
m5FJZsEOuffLaTnca1RARTB01Y3KrymOTKlVETlOIb5ZHr6unXMk8iuHLPmUTUJB
x3zuS7Zhmm4BXoehVwb4HtKuk2zp41xEoDRE1NbPbjQ78hXodmbfx2tTNgn5pobs
3wC14ocZAhnCU1Ho3f0UvWk7Trd6zWmgFlXDoKObiaQqImxR3zq1Yi9JfPDv1/WW
IMkS5KouZ07IBptei374RTnSqOzaqho78hjkKDVMh9A=
`protect END_PROTECTED
