`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwnVZ9+mTlKv+DckLoB/Nisx9oqX+CFlitP73akp0aFQ8QS+zAdq9fRsUROK7kYu
XmwEg5D8DwqYJCL57ChYOZlSG3yl9QDMtRUAMaB4BWzmpk8yKLUyXDKkHOepTdr2
AnvFEFBM+JArPgkA6OiEgSCLmyyiz1bTPPdAjSt96Jf7R+KXc1SIkJq6+hybf/Fk
jINIBnWRuDHR1uHvTbA9AQgYjGirMZMatdPcwduogifVdbm4wZDSXLK1gsCOL0Sh
L8pxNpfD12sIFJcVMzVPNBju3VNWD/dxM7PlrNyncAb3zdloPH5lG9QTDgX112Ai
Mti1ANQK8E5NpikwLYauzQ==
`protect END_PROTECTED
