`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OOKHw98yDudq1iOj0U8tkvVvXBHZSBc3cNhkRFMLgjgJEX63dfUHR0nGRtR8hpSy
J9xfGUD4RLea7xiS+2ybAXMwjqeByNKXBUQjVvqymBo+snOM+qaOBCEVCF9vhSAH
O+TTEEiC1XdDpeyHMzGJfCy+fzVmSmbm6xPHlukxH4u0sPikPkTOIJY0aT1i4pIj
FHVXaozLrDdCFRa068mEFLoF9vHRxZUvu42Xu5ZwNN31Kd8uwWfsWBqcOiAvtppg
4TnbnIsRT/cWx5QfUkNTmm4PVwE6TdY++xagbAud1QPe2/MopL7QWuNQucGJwgKn
fxOV2ASk6unGeNO1CGF2uVxyI02AVROQIrjk7Ha4zWGYzB7e6xMTZ2c2PFmuRn8f
kb1Ss+7xGpAorsIbfFveJkskzzXzDiaH3xu7k9wNhyYMfdP7M0MnlbI1MWB7mZpx
kKi/iYprAK4wzSXhQCYQHu+314gp2Pt6x4DIKTMAFVU=
`protect END_PROTECTED
