`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wcSn/A35E5cF2rCKTbquC9yGPXqOoQRscDue9om3DEVjz/9eEFcOo2XBEIZDFVCc
MfvqhxKxEzhayMNjkk4/kONxnC58NAwV/slj6xD/pQTyXjXqO8PaNYtk/MeYzdNY
kfd4ESyxHiiU9flyvLlW/fJlTkfEoT/pqvIFxu/HhFFuNXA+MCIRnV6uOUHk5QTw
dWCAo4ua02MlfS5U/ZchKCr3YD54aahWVZVJ24KrcOKTbAL1sVbzI2tnnHySVDiB
oPhDNWFF9QWNHSs/wHvpZg==
`protect END_PROTECTED
