`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IA+nT8jREpdzRJ1w/YB6vpbEbR0I7CxIICymbpOmJifP3KSB3Jymu3/vv81U5NyS
tg+T7mTnm9Qdt7TXxwvHAhkpZz906Sn8m/d4mmkdaSHt4aa1HcyRSu6QAbYOKp9v
non9PpSzvYe4arcA5fFWnoMv6K9aJzyIEUV8EuerS4148emGU49dAkXWFHWooA8i
51xknQDYwscd0VfH6fTAr863/67qLe2O4mJEH6cbv6u3Tldem7Q/Gxe4e59F9zGx
KDoQuzRQD0ZsELvUZp2CuSHyL5tfJK3hjqVhq5I4Aq2s8LbKy8p7pqqJ4CzI8X59
EWIlwvpmSUXQn4Wd6DcXU6FjbUhIoFPQ1cRs4iyormK19apyr0dTZPPo7ZbqbjU6
Wml+hHbyNT1M3QTtoIUNYHndz2dMd99FOOUk48BjcyLiP0MsoeX2XonmRyovFPzv
XCxI3RttP41YSu0SWAX1HTgi65kZshe+NNyRO3+eb2I=
`protect END_PROTECTED
