`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ClVl1OiKrpLDvqBHHM2f+SOQc0yaaS5jx0GYnu+o3x9Jvl2PiY+S/Xj4FbULdbHi
oDlUO3bKSnRZYvUiJAGDADdqGbc00l8si+flTZRoVC+uIJqDW1aMOj9GhkJ1hchg
PmZdIv5ULY33e4tkQS7bxYhnAGJb2ixWiToeHX/qnaeUzsnGcHnZq9mQRn8Wpx8k
lnlK3hRB6BablSO6qqCLXBGPuKC61dVWy6m0QhfQWW/e8QT4xSYWY3SSkc6vwCWd
qFNKkcd+8x37CqvtcvGj5vmW9xLmFMSg9CADab+nkIh7cbdBDBiwFJRNXWlamhYU
zHFe14ToCyKv/rVF8mj+1Z+s5HixngVw7jUcQUmaaHUlWt7vKNIeUpZmls+N37mh
S+6E3TrDP1N0MDLs13OFbOuvfOMQF8AehRUELFDR9Hs=
`protect END_PROTECTED
