`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/t1n+5wPaVOA1U1rHdMC7V73BHEfoBfiDkid1t4JJwZQnbiEcDEPWQp9oOapGQ7m
XgUzq3RZ+k7isU5Sob9AHFoM7wQwqpx1mbNB8wyIA49JiuIrwkWDf9SqmJe2byoo
ugBa/Ohp1i3UVDOf565fwDzCc1XMp7/lElGWYGsDyaGcGb6PjoZqJhU0Tql6HU8a
0Kkai4U9CU0SsgJNVljBWY7RK15u8Z0/zf5sF9/Jpv4bFCCXFfUqvkZ836LaOw6N
0OQEtnGfrawoKAB7dtavxxMLjSZExA8eglkP5u8vhJ+SMPKRSFmzti5KkS/O+LbY
3kPDHKewhwlXRheaBxT8y15sK7ty1WHcU6MnNheVx58nCLFbqHUhc6bfC0oKxVG9
`protect END_PROTECTED
