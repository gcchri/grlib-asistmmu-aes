`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAy7hPneCJq3twczPL4wEAVkYb+zqWJgYkqLxpznSEI/ddcr4W9n51dQ1OQ5vaW1
GNsVMhq7Ef6J2LbBvXGBfL2Kh3ImzMrdEgjEtyIj32QwM9ZPvblvXtTr0Uh2n/Ex
DGX7I8Y+wzWadlMVNgULrTEfV+OddbTuUJRovGkSwL5NsAKqXwG0X40GgO4aZk+R
xqhKC1asF+JoHMIT0+0Jf7q4P/LLeTDA/sI9g/uyZ9N4Kt3g1mK+BeAcfpGASYCt
Qcu0MENaVJrO13Nn0UALFA==
`protect END_PROTECTED
