`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qYbQy4uFr2j+eQKJ40S8364Ve1LS8R/FHpf4vm0O875/QPdj9rP5gWiVZqiz3CFC
R1HV/UHY/0PXxhlUtmD+xEhbLC8TmI6XhSHWLkkg34iSlMswIKr4fQZXo9QVzubY
elDgAEEo7lFIRY/x7IPYdzUMNFm1UtpDGKxfVtRpU79zCFnCEnsA39MuAMFPbowg
tWMcCgVxs2T2XSb2Jb4r5OsSIxYpeHFCwA9K1m2KAgjdh+HYs7M5U8ss4lIOLDqO
ODZ6Vvo86cJELHNQ4RfdxNKZ/3NAhW/a2JcegYQWKPovHxZUXO6nJTfV00+fddaK
a9avdKuV5S1GWA4ZnqtZ0w==
`protect END_PROTECTED
