`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xDs2/Qk5ynNZlUYkqh7ZgPpZnpDymew/zDr3itZWYCh5YB4C97SM1q2qNcIXE7M
tHpVi8DhbNspC4JXLV/KrrFWL0Aatsqcqfp6A1WJz4/0IbPf3U2Q1t/jLf3/yrmM
31GLgbIIU35PjgikIc392YLynjJrqLrCRccZGrVLAxUsxI/l5yOdyr25JdKe+v3X
qNytPCZ1MfLfSri/k7Hq9La/fP/D9A4y0adZJbrFxXWoSF8Qr6ZSEnmKHm/HOzvJ
tle80B8oTULpI6fqjL1e+Trlg8YpJ6VhS8tBdS5sDyJAOqZ4wpc4fQhg/ynxtQXm
pVYQid1LjaJCsHlngyB06gbj1LCxyppp+vPuDWDiZPcpdA5y+Xbt9nkJBriMFPkp
3zEv+TZiHeN02PD9b8Ccp8/RQTcImppMAfb6BkPGd+dfgclgxhN15jNSOD4Kh8gN
NHzqy9UCVbafdJ78FPuGyU8/XeYt4BO00c9byHkNAg/L5gXsdXzaukp+0+YNGftU
DpUy9/M+9Uc1Z//x1M2hhV6wOcKwQXYNrf28SuCIhIaYRrFSHaPb/aFEKiVyLL8d
r6EEnVM5QUi25EyDnnqzO67m0vKSQow1Yl/BFrwZgIfbYWl5Ob8UrLsjkem9a+Jb
g2+xh/+yB6b60pwsm6WNqn8mYjkNq3kphh8BPhNf5JoVKl5hxok5JewtiT3ZBfN/
EKqQ1apWHNDH7fEAoeKIyp8fFGLfnQFUKtelQdvo4ugOi9xPCfZCDoiObDm1gld2
EfRG+93yGH5UErFDdCVFp9wf9CjmDd00IY3gOxIgQPIbyavOgHKI42iu+Efo0iMr
H0jf+PFqb+g6xkTCGH+kOcXNyuRTOeJJxUrttXOvP98=
`protect END_PROTECTED
