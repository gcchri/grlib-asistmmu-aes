`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ktqdEmouQkFBXegix5W1y8h7BgnGEaxK3U741bGv0Mf0eNsIjWgrHCx670YVxQL
7tPNibvqymxNjD4f7bzDkXh3YPGceVK38fpxbkeMr/Wxxu4c5bDQoYoGOd5LtLXa
cNvowo+pbcRxUttubMbTJ/O3rU6/RUZtceTLKKVz4sdpot1pFH2QlgRZTNR5t8tX
eHnjMmNeUxBgnVg4Jd9JvETONF5F1r3fyUKA4x4FiZNfcze3dh/qsIklSUQo3m9F
Kd3ORnkipt4YGwr4yaSBH6f18VjzGWgevPxggZSL+8JgfS9i1Iaxw0bLHvW651qn
QUlyk8m0lHUbE4YezfIn7AYg5TJYQXX/VaYUY12mk2ydylSlOcthlT7NCmIMxL2R
2qIjP7pf8xDjyyHtk6wbTE7MsQkknWCZQXwTHzi/uJkZby57R7peWgw2G75Iq4+s
LbyCFMJTiZKR6tsMo3NIUKGaEcuhVtZh4taJm8UDVkhnNWnI1ZXkq1brvvWhyfOG
S3pp/gJKWlohj/ark0IvK4eApFv0bXlJDLuJCl5iFCHkd3PsCpn5l2Zitgg1jjoA
MLbghxMe1kZg7eBfZYoYiUfTf5qK2/TVSGGtJ5BHjh1ULu2eDE7LTSm6kQmJj5co
i5l24aomg7AZ9oAlEsxy0tje1U+j2b9pt16PXFCS9xXCpG9GwwYME+oFyoaSRckB
2DXYoftRWarXqFaJdcHC1uvZe1vX8NJDxhhiLfIRcY8=
`protect END_PROTECTED
