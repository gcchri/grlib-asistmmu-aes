`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GB5/F6pmbKXi5ni1mqPWVuqqcir9O0UtP7p1qBHxcE0B5F76uAfI7EnCbwtnQ7WU
E7BxEvuJ2nVsWMQh/e94fApy3ymcUys96WQEAAtNQwW5r/R1KFl6XcIwNVFH/9sO
lmWXs58rOJz8N0Mo5hJHf4rvlqvnwYzNirzn8L9F6nEvW/btr3Z4VOcESgX2Cfgl
qEt0FRuyTfyKowpUUpIxEXWofwCotUfxDMsjjuj6SaHCcn/NBIwymoNcpDidQHJS
8ilMzGbLI00F65sKO+EgR/d5eV0fKq75ceGyGoeJttI5NIaBuiWogGH8vnTnIK2N
UVoOijNHBJGED/plsYApGlyhHwfghDZD4q9cAV/b1nw=
`protect END_PROTECTED
