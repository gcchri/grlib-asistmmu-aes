`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ekH+ZuRFa6hBaN11MHbdv+5oG2vygthopTKhmwuWLTbfRLpXkwE2bofa+7Yn4kTO
kr+RyEnQmvv0VUNM8nPfWh50i4rug20nT6MtumyWoFwwtWSAcuSf3F9FuWFgmmF9
aAiFq7zIGxrroDoQuX0vIN++4xpNUBFvJIkZ+uJXAF16TE905P99BF7V02fOFmmR
iOYS9jre7+tH7K9Edmw88All5agzfb81ubxjtynbA1tZhyUHe4ZTzvMntiBtVCP5
EdqXEi7faxNAKqKT1VVn25poXhfTcD0iZp+XGjiRiDc9212P6bE/4vlgCIJoifSe
pCt8SQA641HaK0k7IiYfKX9bPXSlzwTeaGOnLT3+h72zS+FIVpYLySqh7V3Ej5x1
OqhEFFvP0H/RljkyuQIYCz8mRloy/msy1JbyWGHmtyPkI/Y8a2TCFEvis3f2m6Bz
ITRMed/xCF004QgTO95jqUId7fJpE834HOngmhLLGh/USHKQ4K5bLs7nxiAMWFQP
3vp8+dJF//btsPgGvorGOOHcBp346SiIF5yKWA7SSjKBqlGQ5gYKHWEiKVi4T/Qa
oQNqnSiYsODkm3QXcs39I9bL8jm5EoOt9SNEJDFBrQgSYxYsxJbNYI2w1p+IB8PE
XG7qbb6eUiwReadtF9sO/A==
`protect END_PROTECTED
