`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yKwXoT3vE/1ibjzCTRlWpy0dRXBOip4FnmhGfmBpefTO3sP5oqjAYuVv+rbix8cH
pmtHFMrhkvjYPkHPd3OwlUuCE8rKnEq7pdB1gQmeKfgElNxRPRtYOIq7H/Ca4rRy
coUOZXyunDQoSMQVYtqdkXKG2aUcGAbdzKgXVL2rIeyjxPejUq7BEiQrtLcGemHH
vx4i768oEOaiac1e/mmmD7xMqIlsugAmHp9hDsN6pw+3TVGdni4dy8cqBjAFfagP
zgrgYuqfVsWu3lgcRgIlqHjjvaq/TFnwKFvWsAFSfiOt+SYzP4M3Dg51OjjVMgtk
F389qgWVJfkazfbubgc87pPQ4XVh1gvQxG8XEYGGsvZYYGaqoQOX5UwoTAiTmNYA
OYJJyJTKfcCFuiZ0poBI4JhunbDML+VdZ3YsLAAnfBGPdhNauL0g0cdA+4cQY190
Flq11s/A8D1KDx55I5psrrtng9/WoCxYGLL/nGY+h4AhoHQ1sJ5K3WVAFgJTOEem
`protect END_PROTECTED
