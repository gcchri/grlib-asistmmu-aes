`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L/ISc5PqDhtTympG23KodH9oA3PGuf19QrxZG3eSVI/IouNMTebdLgUqhQJQvZmj
OHf2M3zBqNF+v6XUXjf+cNHA5JLfQR8Q73PEFMiOz4zGsrOv/Eq4JUXK8US/wj3g
yzoqaZ74SnrEwCPOXl+G1mzLblsRPoQvqBjZtqt6LtQg05bIbMAed/IjBXYMp2Rd
tUIJUw/NMqHhu+mGdeJuRHSsNsNWMQ0Xb9F51/zCiC+lM10EfCYzgGrUk1ubUDD6
Q8YV9Bf+E8ni+oH889ZdYTyJWtRdFVG1C9JLmMjQnIJCHMR2CFwwi2ur/9inZXGU
ApN4AELkgDYspQiylhSuksw96WF16cQTllJ/9LZAHDoFeHF4wQUTjIzajWnCB0vV
QZp14/71BzRktlziGjYcXqouoAFqLmjgSuTuNUmX54fmpkHYkFmRI7zE3NH40SHe
Jycp85F4Ii1iQmarVkYBfzksCUomO3Wvug7ALndin/0mPikScEkG8iqQiFUSenRw
npOO7uB4PG6BZiD3+1O88a/49dv8C95OGEJpwX27c++678FmricNIq3LjXDCUL2D
KbwLZQ4erDZAqEyfC9ijtNWBN75VXGRnalytLVd18R6OQQeJuW/eMkY8+L+4IgBk
0czurA/xAwiSgnI/5F67m6NmFXTqNzNq8+d939FtD+i69USDLUNvbke2Fb7gWaPS
q9OTeaKZPxdJfq7USXO1mw8SOopnQ9RI95w3JvJ5/RbZ3BvOB7PNgvZ4yDWeZ4TJ
XY+CbyrGNNY2ZmBII02gG+Gri261EpLag/sQcgX3e/KlyMNVkmma9qMNmVdbRNA2
QJVseMF0F0rEWK7v9uw47Sm4zOQ7UWx5nvGcqdGtpcUl+YVID6zPscMfgvpWXD/g
HQwGTMyYJ7s9uS+yVmnDBdgOK9Qa+Jq7siMsZtvzga31RVCosRluAgNY7w2J48E6
75uTDKkqihefMnjZllaqLJHtIR0FSS1jQsONzkG5dNUA8Rdqhss+96vVgKr7ugmB
`protect END_PROTECTED
