`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TRNUt0e53rZv+D7MIxsq8j8r5CiP519i4o1tfkFHpyqgaBmfFcNumJuKENxCCbam
b3Wtlt8esc1UFHvFWKGgIg2+BAncCQXZb1hbd0Segr+pI+rPqE5UO4XIDDC2LCYq
ifVTnx7AuragAl0zfI3UG3dgRLIggu5FYDMPguVZgIjDm8lKKhFfX/yS3v11UhkF
2vgDYKcSqXQ4iNY/+SElVwk3K2ycuJApzpir6ThIjQAcMHQ9ZH960kTtqfsRiGkQ
q2tR/83lqnBuOSMdf1QKK0R6T8dO7dgBPlbLrO52CXvZPvBFELB0q1/VdVP85wxz
kTHKnAfXvNmAxTff1CMcF+xLi44nfcDNq+w8sna7d1F3ABolMB7+CvFn32+meUUX
2QW9TKYYOrld9BEdv31EbEJy/K822MrGhhcxHY4j9olN+69EPnnk3kNN9s754Aj3
5RGL+jdu9tu6uwwTRZaG2C/IUYWbkfj1jgKJ/AEbf2E72bM5k7p2pCikn6rHz9qs
`protect END_PROTECTED
