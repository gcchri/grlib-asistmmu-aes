`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJRGWZMeHTf4Z5Ts6Sm/ruJVXnSH1YAs2pdkXb+3FWOCJcTdy3ztdvFuHy7/PNYh
l1AuBEgj30lkqu6Napw5ibOBF4ycwe1y7eKrQWJ9DKA7/X2lXfEzyZR7JlDjrk6s
CbYfuTMcBEj8/pemDQfwQllto/Eq4qUZgfXXBHsRi1cf+j4joxHb31hSARnqDJ2+
GzGnmSXrhO9SsEzW/+lMtAmeyPJqu+Q5pjB9w659tSG5EBnKoTBfrfkHOi07XPn5
HxXWNV0gMgInIsIY/qt0H5aMHD4xoaYsVkyPRAkI1CVP11VFeMkvzXZ0VuwN+bEd
007r41Ss5LuItHCN1ld4s/oGSV9YNYWGSNMk528A8jpt7I2MWc7PogjOL3w9sNCI
IoZfuRjiwcoqCteWgc859E4JmNrgIgFEaP4JWxbG9hQRMHALRcXSuJ9cLi8tPsYd
T/w9Nn2tAYLMX+BxZA03fTfJeLSUZhHnIWK8x7ji+ZE=
`protect END_PROTECTED
