`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JI8lyXd1ndBkSdiGFD9bCZU3HJWp93FijpeFpX4IJ68FzAaC+ynpBRvQ9HWPKCXl
KSjYOPWBg5S424lBAQYk0gs8EBIicW09EmJ+08dK50yVWZTHzryCUXhtVnPgUaKo
EflOLMoFqHefE7gJkjx+R1/5Z7gd/lNThF8/aD7R4RKmp9a+jfTm4xgzTD/lzPow
Lp2GEm82OcPZqzg2Rp5XDF+dECPYu4rt7MC+k6gyL4aNYlndaA3vAul7lCHEVCbN
IWgNMHoxSfH6HvjYHhGROq09XA23aG9xOF/V5gFWsbvSbkyNgqcgFahVzpl6XyIg
a/Dt7oS+TDkeZWyy78uvTriX1ON3vcnT9TuNl09CYMJsjs1/ONnQYWr2Kj1Cuh1g
11Zjb2ypjQV5sG3pZn/lqvwWeyfAMuU8OT0vNG5F2QdMY8UQtqoESF2a3fH/7X64
Axav//Re5L8GH5lVl2BIT6vCwGWv2IQjROByOv5khmW//RqvpMNqTuislyUo+qic
`protect END_PROTECTED
