`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zz99oQ/5hypKAf4ZKiXNqV2qu0y394ESxk5kovglr/c2Oqz6OzuLaV/29Gn7b3sE
9n9kxEmb3I0f4ZKTLhR99Kqn+vb75uJtHiGHzcsHOD4yiqGjxZyV/IQYnCZ3Le9f
8iO/RFiRVJxyCJo98Cwy08pjprK11zDq5LTzI+/Pogn2titlLxAUQmsYW+Dspbvi
Kt2HktUaiwqXaTO5G/DPHLSWpJIRBflMHccuJDQSpN0tjFqGlq+rgVnJJoc99c2r
dO0OA004XD7OEGvTsuKCB1MDM66nXoDa57PBWjuSmuBAwAAO/a64LC2vMLhwWMit
1xVf+yhkVUFPiC0yqFaIDZptnGSNI+Wqw9ZTG99AxvujltaNeEx1AWAOj41a5cGu
`protect END_PROTECTED
