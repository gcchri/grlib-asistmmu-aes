`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6F/Oup16edWvPg9EUMW/3k9y5a4Bg8tdQeZh/qS5bhUtURzbktHagCTnDQtzlTW4
MCwKz17351tv7H2aMRP2sYej5G+X94nZW5/ZJxEWWRCHGWH7baiQf4Pr7zTY33zz
VdPOznDK1JwVJb7HrimtW6XnlCn5WRQLwDHCPpxHqH8p3CjWORwSDDYAK/GD6h4G
c9yBpnWQqDguyy/H0/fcY1AdP4ebiiYpRylKGRGa1+rJ35691P2vTt3/PSI4/bcE
HuB/A2Cum9pqDEUbEeFVxgSEJqHJX64cJKoK5Cr284XF+E8w0cwIn4fvAm82lVCS
XqP/gS5/UJZ3eOej2b5+SUX7Ny6tKCwvymTFlWmEjS8uQvv3dk9xwOlMzZbF43FT
K9bbgAT0f+1EB+e7xqN12qrflAc/I3UCAQupubZIZAOF9ThkTzTL6YX9PiXMQiN7
`protect END_PROTECTED
