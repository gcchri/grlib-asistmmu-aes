`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDcL0TD+JBsPXeLBa0+cLLir36+Z4LRtrmeWpR9iO1GMm3VZ++6rcWZpZqr2M4nX
e4QTRCcZb6dDIdmoQkGNyJS/ltS2xd5AVSBhuSjAgDF2Jfc95XrzYjmxg5kWKA7C
Fvs16ldiaQ2kpCeTlsStnrQ+VRFUfdntyFBEMn925Onae76dyysD5imRRO7sDTEv
iQM/wD61SBQMy26y/YjESaoJj8Ze7P/tuMJIcrEVBJ9ftQxlsqxsG8b+CKVmmBNl
PIKReQ3wAgTRHOsUdft1hZcMWVQGktBcjy7FpcH39rPm5mBkovcLsLxOCrw5xOrD
pc3D5Jh9gc/WYSN+an4Ozgj7Jg5qXaIPV+9KueAtQZtfa80o1Z2/3YwJE2JDFgb9
O1+bYPQXj2DATVvKm56vOZAcczQQcwMQTi0gpUk/T6edLf0xxlzpQkkiLneCf96B
/a/tdwcp7EbaAElDR0NNWoD8mT/MUAUthw1VVIy5s62Eh2UR/Vd6xQGVvIu80obp
dCxCIWr1qgeeOiIv0BUB0uG/V3sDG8ohK3t/AmmbQSqtsvccabi3vHLg8zVHuN4m
xMF8vVpblQqMYDTPAzw/hfVCJ+X5wkHOz0gYMdwkl1PZp2zcQV0Qr1+nZbJYKS6F
mJeEdX58KAPfgRo3KTxzGc6L8qKtQ0CDj3ySgvXO+MMcVJMiJJtREKwFktVSdehp
sUVdi2zmDONRaZpyAgJxYgVPKCEIlTu9CbbK5aEJl+2G0OQ+iZjR/qM/L5SL/QXh
Xmk4fCqcFaLetR0cbMZRl9gPakWZATzDXJRpYrCcQRErvUjo3QSKAaKeW4YwyxNh
SBFlTOgyjmJ7U+Axncz7iBTLAE+blQvm2wk1K1BTTftoF+101cFK356pegwKZ38E
CxltuvVd9AkfMtt2vIwGp9N4MLFziiCX+QruKZG/MM15To+xMRMyMFOQ3kBX3h7U
U+4kQXLqCj1SKPdkLHgBL95GQa+F9Fk8ptvbAEA0aYJaJB3d+qbUYd5Hibke8pn+
ItYv8TeSdp0mjBbvOPUNTVd12EvLkjUCAnD/gzCdLX7/CMyKWlyHyR0hsp5OE/z/
9vLQLtRlufko2LK9rU57NMclHp/yWmaS5CbkR55uf4PbowIG4UbEDXYzTNjLt67U
PUjEMPFspgsSZBAHQHxty1JpHocXDt1OSRhTlhuRiszt+yfr5NRYOxsots9BhUEi
R5L4QK0S+Ha4SxZ6o8lnVDJwTy8aTzoJgQR64swMJ+vBz57mrQ4HsND95nwmEPif
ME3MG4RoXT/88A1ueeY8air8ZVAz39oHCF31qrXS5R1O7+7OdEXhhNS0XtdsttVK
g9e8E6dyADZjiszbFrzu3QEo8s+vC2mUNN/Pixd8BE+XEyBQk6vPfUNq1JVfbu52
QUgbvwRZfKNi9IcnsDYPNKZ8pb96sQWS3xM9OsAc7DE3K9Hi3ZEZd9utHS4I7R+b
eBpFgPU+etWlmPXLj6BiYxHMuBmgOCycxkhMMVpkH97MMBMTKjcTSBbeFsykXZTG
67CYDI8TtMS/kfp6FUOdNHM+bzM1N3PUYOovugOVK/Dqyb1IFlFNlWZe9tQgghtm
HjrJIfFN1H0SFXgZytkum3O85CwilYk44JLeXRiddPCwyFaC55tH6IKRDqI1DbDi
ypdAV+mk+9+iRqT6JR+fZQzvs4LlD+ru6ZMgCwyFj1aTNAu4lULcKtBTxyvitorI
2VCcfshSwAdBK1qEQD7v5RvYkGeyzZj67OO2hcrn28rD3G+Vgr6KeaZjxXgHSIIx
+Yi4vCiHUhN9+he1FKX3VBJxHQNakon5PqvfxVryMV4EPri3PcHcioRbHulq+BlP
cdkSJjVS4jCIH9ZEEQdWXYVrcDalew1gW85ssmUtSCd4D6CcUrsbbAK4XpseaMfH
0ObTJ3NZz0tKOHjOTAJt4YlWexR07TjpqqbgN6NpEoCYi0XyRrIEQd+NSBebYDZj
hL1Ll7cLh40aILym7w96a6pBruGkhjL/1KGiEm1e4YMgCCtFuno9KwgysNJrOUKS
aOD22I7kkp7dNyUQsXOyM6wEVdoRFQWu6dS411826KuR+2ThFXAtnTQIGz30V+FB
eeQtGvFOQe4o8urC4I1ZZ6Mewn6olSZ5/kAtKX07v2R5H8e7mg1sRzKjtrEk1Gah
q/ebxc/BbZQcI6gmJCF30JhPwLS0w78HGbWR8JxzGbX8kf3EWMt3KHufLSnaqHR6
BiY5UmcGOR6T8/AMvUiTtiq6XCxB+CoKt1DaQGH58jdDNIrshG1Cy3AndvUTFmup
FCN/tzJlEJ8yXqY2hUBV+q5o+aBXXYBBrxD3lXysGv0FjEppPp74apsB1wfSdi6m
k/VNUyiaSmIcy/3ywwCMK/p2DmV6QXAMmOY7195IfSWwOcgG7/w7GviXr7YsCPOa
Z+ZDqL3nSv2REw4iymlKtJ70W2AJKIAKf0olNi+Z08m2sxJ41WzIIEQG102SsnUq
np8w4xP5k980WTulmdI0hM+Nv7OlXf2tBeocm7BAdqrOTIsW8RIvqzilBbXL16eA
wSesLefx66eCwQlkm7K1lgryBWUlanGDXlftp8o62OEA+WEm/81JxPuRpaGNhqM4
DRWmdNDltLvbnrw3bCI46gZQ+bNI1RAcZ+nWcdr+f1T1rlyg1qNiWnPtCsbAt2s3
9gXARncr5xm4NeuXxtbw0mOl5AyNLM1M13vHaRBusmEAY+T+3CcHRzslvYAS46+l
p/QzW1jA+qneTNuqjE4XSYVbJajMaDyrwf6gGb0AOixEKuGO0Pwgli6/mRZLud3r
BMDriieC6QTfULX/N0Whxn+L9H70/O86g/KgMTlbJcOH8uarO1P5cj4/PMXBP7wK
bchYcaWMv9acW+a+jg9VEdZDzyHAXRzC3mkj40jtxSOv/c3pYOjxWwAJb+TU3Pf7
KfC7//5kQRLj2h6PYifXg5wfJi3RQdTQrriYNKU4nazBLsHcnrneU7ZkzAvfExTI
CUnKYxRnwOyaBOWvIv0Bng+NDuknORll8xyY91uigxcJOxD7HcHqSyLOJsyixuf5
kFY3JLlIlNuDD15P2ceyDWI0R+CTej5LINrgq5BPSg1N0UE0jOy8dksEraOJYCkT
Vtv/Uz9Rsbx8GeqPUDC7qabyKK61pX6wexwqYc30rphY8Zw4BdAOc3KKC6o6VGrT
wIuVzsJieC1PgC5zLxEm9fWLbHA18XjLc+MCXOTdWsuCZTQdnbfUULjMWDcMkRVE
EltU2PIGtsHOlwoF4JIadlKPSr6N2zk3aSVjo/42uCaLV1qxEKJg0LFoB9a2OZjB
a7t585bONvHCPJUcCWz5Y/3zQ7Rx3KdINRkyRvSiT3aQSAmhjP3pRoGdcZyPG8iq
cHM2S4dYhi+e9yvUfTrdKxdi9A6U/R8pq0QlQD0wviANlPZQfRDnmXIW3jKyRswa
1VyFzC1/eVCzV0A8oxv4q6uT4SqsaJLwN0TJSkYWhp9K6pfd2A3iDbReETFp4Zxi
3PaHrhsZ8HahdJ4sB55FzTaSMPIXn0mudj2Qw9NocRj7A9sJIbw2XNJQAf9XTmb1
2glq99zP3cc/7PgaSYU8ZgPFYcGJKuMFnx0/F5tqtREqHslM330yHugLfSf/Nb8t
3l984GGHw8SNG9eRdGUagEZPfunuERycr7q5aIREsOUQ1/S2P/MpSiZ/RIbKSmjv
lDeoHRze2hHDo/+L8+MD9SRmEK29DGe9C0F038PnDxYNnQTmBokkcF9TUD/nSq4U
nooRfVdasxSHWLHAYpitUrMO9gzBNxdSo7qU1UkeHY6x5KxHVhN9/yBY7QIDqAmK
p9oKEfr6CnvmUmnAwmXYki2fUH0z1gXcn1Hw2dbx8tzGqM0p/NRIs/hAa6a1L6yS
m8mmGWRdsiNE/r79j3PKY5VRMv6ySbvsGZF/9c2FChXazu2CP8znKYIvpg4ADLtT
xz15ohNt/IU68rJO2ovw8MaQXWjZ+WdQnOjAOpQadw17CwzvhBIMBo7BHFZ/URaN
r13R7plilVU84gsqSEuz474h4e3R5RDL6yGK2tTx+gJu7kCg1JjaBs3c7UTFurdV
5a8kcEGYUh4MfVexW6JzWrphZyvyshuIWkBJvLNL1E19GlhqaOyZZc/q0zOThVF3
Va2A7LJ0b0Nf0Pa89YabJfC3oElI6ci7a45LYYkX6y8uLBG4cWpotw1UJ5s9nrk0
jLHddhO5qHHD8GaCLAAcXNfFZtEXLN5HkWvh4R/yHSFsV3oRaohRr2HOWE+fzYem
J4GWAYo8a9s5k8AgstMV2MbT76pPm+ZEVf2/CfRq0oHN6P1gHbOXhv358Ni58NpS
iEqtkNegjrVofBzi2JopR35RTBgm+07bRRpZcrTq3tardgYaxqSj5UakXExJ56OF
ctKwAA9Pi8KLsJY2tJ433N8c/Yu27COYwSt8f6f/GoCWv2gBXNo1i0zf37puyzzK
iMZOL+VbxAKaYZp/QfPRwZlliZY5oavbZX7ul8rVJU93wD4y5vWxHRIe3umMUBhj
HbKVeL9ZWzalrhv3W2g7cWNjnXiWzV1uytAenXqZ0pwhWyHUU+jXjmbfKIONrbiL
PlxJZRh0O27nYvsU5DCgwgI+jTnpmTxE8ANoBH29ovwI6n2dlP86JHmi3TXqJL49
nNRBZJufmL2rmqtE5pcFSaYdkTczVo7YGjyaTBGb0otWXunmBj2FonYX1g5cq735
5ttxleNneodDhDWO1eXj7yfdbCan9lQ/QukBZh6EcDP5Hahgpiwk1pyyIzGmgjIL
vxyhA3Qg/U/6nkg7XdWwXGikq67wYVfIcOp4eM+7hQ3mkU1AoDbGKdkV8kSYcu5V
N2igJEaIJV5ElwQIoBBLFgBi6LXacb1IMhSHH0hB6kBAEeKfFzrIesqhTM2IQQVt
E+Sqbg6A6vO6/ozZt1z0TbFPKuMz8AdXN6fK9BuzJlSGDaS9tR5WplG09s4Utbx/
xVQJ7NwIsBxzlFfnFvJ9EuJZMIM04cbmo2grqv4zwXOKLzQFlZRkGgTS22GoSyzm
DMFsdtJeJrmuDG1ofWnYL1/z5yTWKsrHAlsZxnMICnfQmDdHHMdugzFlfK74vOWQ
tN4wB/9DppVK1UkBKw44D9g/1EX5VvZWonEOQhqfWtHupu3xqcH4MYNRifp7+vwB
5HGYpqlNhRw9RfRobOcYb2XCHBT7B2ktEa3FwkbRiI47XsV8DR5PvDo9Fkq54whx
YOLeDjQkzXhAmdby7FxcjogBVn2kSz/L8eolTP8UhnUVK/3WY8Z8FsyEFIPdFH/m
wA4zqb+53yp5ZgHANcSYZjby+7fEKZnqV8mgNVv5aYgm+BqiPKuQSAag+UvqjJ/F
yDKsy+ucmX/pBlkNNlJLRWoJuX7vtXacMHzmPUxTJO35o+pm57p6BnuEv3hRfuxZ
sDAek8+RR0MldONafnne2Zu9OCahzVB56H7cHg/uFVBaanZRlKScg5lmtcvxP7g9
o1rwUlTejbC+mYlu5/Ns+drEKDIBQYlpqOWVjraxT97mgDMs8YARUD55gpTW80Mq
lmjauueN8Q5QM9iqLJ4htElRI9ogFtyXBrgYqcr7c0Gi5l87I+kR98/p+381FDf2
GqafFiy0wxzH5falY166pwuKezZPIC5kLcvMuZviZnjqr0mLnb8cMQz5OLNvZVff
Wkg8Iw08rBKzGf99EP7qJBlas5u4ppjKT9/zFb2bvnzdgg4/NxAep5Ku2ewDOdxS
+5PHpeM7Z+/NTMuRqheQ2xZY/E1uCIbirApZj0fFDeS3KrEn8qcl/gP3vhOWqing
46quuibfMnz3yZSq5T4EfoLdeBPYCjiRa9F25vyjr0ZopMJQPZ1WG2rg+NJSf5oT
k+2ZicsSfMtU53K2l7axzpn0T9iBopfmmUpIQYqvrDWDcViPxXJY4xifH1iKOF8c
jquwRID+iVLvAQEbaIP7kinjZ36nCb+LpDPpHlJGUf38+zMj3LA6K29gAXC21GR1
fyrw9uK309Sz6CNLOXjsUyOAloFeXDGDy5eFKKl6E6crnHeS/CuMFxcsh6fN1D9Q
vCezjKCZtTjZjVwSkY05wZm2t5u3YSNFvDntXQINPGKmm5Abbfebg7cbqrMlYqV9
1RnhXzB3QlzEgY3VcWKyyZqYIGiXrN4ZNf+Om7r1DCEfBqcn9Hi/LU2DxxLN/QnP
0qXTlB+1oLNAZ+uqEqKgJkDeh2wZtlCtszEwUUsnaESZjdOgQIQRCVkHfFibNDw6
tkEsmMdSVHg3ERnzFdOKC44SunS8JdegsLGSZ7pRsj/QQ5ANVXMtv51aCJRzrPjk
ddr3FttGVbs6KsQO046+ic+5gSOWJCS2LhyDyXJ2HYqJdV8aeofZImYcUtfd8i26
UEN2x0D7Ia9t6oZys7nsKQZCfVwOnui52dd1IxlhHh4CeRkEkMCYkJ5Sq+CGq/VL
yvzibtTlSwPWsNSZBWWnB/k/fthBYHYjqyHAQDLiWDsRdqnMbb8la3gy34ifyKop
tm0U2jBPLm8O2RZ+2f2GTpmleDSJVY39vYvZRsEHYuMd3m0jidRsUSS70zyHw8JG
BFDPQ31ROtdUh72+NDXhz/6vbj0QutXoOgUo/+Ej/GlUq0g4haS4t9CdjXWZ8XbY
qDNEQ7exzUkHmninJOe/YimXEBqybSQrhtkvVPkylQccOeEFoQX6nrPuvdeU7c+3
2fO8+omSs9quJ+2slhKoGBv6LUjPynLdIGTdYufnpjgyE9XaMMxdV59pDg8vixkA
JmKLYIHno3bIK2d4PHcHPfr/UOFNIhQSjbjPgwoKBmZjnEE9lxinlJoZ2gOzrkCz
PO084kMadRMKxDslLMgEP3ejPdH7hS2L8WaoJbs7mqM5LySWfq3gE5AO7ccFC0r3
FJxpOcxs/4g5+x3zbvc1dXIf90ytU6TJesJ/NcS3esvsPjR+e7CnW0UzLtm2z6U0
mva6vhEEFspBmLo5h+FxO9fJFz6iOMoxW+POfWqsmR56wc2+hc9GM7mW5uAAG5s1
r3QAazUJcX+M9Gf9yTuEpr6wDwHcfgD4ABdvjK8Vb2mEwPNa/LW5ss9daRQfwQ5y
Cjtwifrjvp5A9O301n3XWssSaQfh4URZaZmzRD7pzkF6MXOvDLM47LiE6T+t2kQX
WRrutUCb89n0Z6Wf4b02QOoo5LKAOeaWPQ/GM0HD5+cE3Zh0orfmTy+uMIWzyooI
wbUTm9jvWQAhE5BLt8A44KBQj18MGyOCVdAzDJ9nW7N47tFXQAJouF5CpyQckJBe
MPHfwgW8s5yww+UG8sHHWtuJg3/eLsu2XK5lRHabB/mKXzLNtOi/BNfvdtJ5yZoU
GysW5oUg4LSp1RZ0Ccn+yPixODFFu6VYdPhhKceHfyIwhRj8HvrtjP/EKhHNPiwe
E/S7292WylyGHqTIGNc6mUKkxAnzW/WaluymAXo2RNLAYpEKMYiNoD+LI9b+Vr5h
jvu6AuAaIxwj+wIj62Lkb+jk1Ts2CxYg5q93s2aKECJ0IUgvcHLqglPEspDmO+VK
xUG6xRvzENnF3JaWyXlCZcUAcmB2gy4lXdYiAY3dqrKXseopjeCffsXTnVc3w5Dx
b8xXFQbpmW9xgYyfwI99iLlPCGcly4ra8zKTchOyqv93EdCS7eMJWZNPC8QmBgfR
mvFfDDsihpm078cx8RdqhMslTzhPljwiFBynTUISjfk0doQTE0x90HKGU4scvrYJ
Tg6IUzZw1gqXknPLfVQ658vCUAnWC8kgut6OUam5W0iD37s+ytu+eaS5XrDWDz2o
R6hTt18JU59lftXmJGWy/v+0xmjs7srTZKHZbdMHCxre1auhyESUt/HQQSguR1at
7FEa4V61GvU4GNU/yRMseR5iEF7lP+BNadTS2x6Jb8R4I1WVmF66bTVtwVuDbY38
NELtWcCkgXQa+HBddGMmtj6lAE6e0F6Qy12KJzTRpnhqLstnuti/tKEuX+5vMCDK
80w6pdrJZ5UjFg4xbwjcAmaP01VtrBAUILhFRyGPPwIispijUuJBVEPczjEX4wcA
HZHdOIDPixyNElxKGn2SF7d8eVkSnunrqDBvXHmrH9BWuKnSwTyP9Dhr4A5Z3rDF
5/2yxN4pPWKchD5U2BYjArfOhcIanjygODtDRqPOHoKOOyIfwkLo7lItwDp8jJ0w
y1Wh5FO9wwH9X9tTEFr558+UUSgaUZO4iiq0McuMT3erItEssv98FfkczXXmut6l
ohYSq198mL9+cDfDjtCZtRVU2n34udCa9L1IxpjrBOk4IKkowJtER1oEczY7QQks
MYzMpNLEpOzKrByQnVC1Y0jLj+uJh3ES3qwuqkJELjD77p6GwoL1jMNpSPANjUtU
amgKok+PgvmLPKKC3AzgUUXwmDp4JPC+XeMyD2fLmegmhNsgmD47YCvU5CAcYHmo
OXicTjL8LpBN4V/txxPTEVRyI7TbM9OjJ2dH8yaRULKKPIuXt/clYVbZDRpYVPEx
kPYtn+lYoSkRWqhATeehHWeOrstURRCbYkQiJ7QDSB1RZPkaXcquQZMjwZQXuGqp
TKPVmeRRiBSWd6EaYpPFFZ6StUhHgEW8Y/VyFc7Tz9DVdzpghU9+OA6DzkFJLu+D
NbQmIxjKQJv97BkA2Pm7PVPdh2MN/DsFKxmIdZkQ8hJhYuF0GhTHg01Ocn2FT276
hJNbDm41v5yHB3WyzPmMZ7Px3HnsKPGwY3MAKd6rVo3RLsF0OdETCyokyAunRAiK
oQBZS8fYEnDXRQ1OzWbAlxryNGS0RAdTPR32BCNA1QFo3Jj16UnYnUJPcmQU8qCm
2/8CdELIGQX6PSzTBx8tFVfkvT/HzSZXPNl9XDTVc/0nHtuOmnRzs23T1gE2EoSH
nEpRGth+U6Ai/FtTKHWNjMrSl9R6meB4H4mu/gmrE6+76qo7aVb5uICsq+k3E7dF
wMZbb34GI1RWPR6xiSbRW4QBqHzgPvhZPERFyZmL02pKd6YmFtODOPD4It1CiTSw
WosaKnMpz0tYdQsz/vdLJu+jXJAbtnaNT6+0wN8eXbgVdUkTUlxWg0d7KQaL/zAA
nt6FjvPIl83VrXgwlUjdyNLwNRDbGtFbWH2Dn/NVA9GTF12+kG6qYOrJLUQc2QSE
`protect END_PROTECTED
