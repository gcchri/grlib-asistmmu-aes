`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZeLRnfT7XnHWr/icBUlIJb/e3V1A1bjcZdf17x2IRkdpm3s0bbOChhM6PU18pOGR
FwhEhlOI8BiwFoS+6loqIR0tmML2udPo2NwG1Se7i9qbcfvC+zCYRgpPJUEfZNFk
JngC0ko+k9Io17kEP5l+02sd/ldP8d3ob1NeUAVTnhvyNe00ds4YB7g/Ul432ey7
SPe1Dr7D5vTSP1VJ5bn6EIGtmxU4ZCNhm8zr/iOD4LOKKUQUlsCu556Mi7ePKYvq
FiAfEWcixkDze13ITc+hiA==
`protect END_PROTECTED
