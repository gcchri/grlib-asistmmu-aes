`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gNQOk/kOseMWpVxhs1X7g3zzr9ihO4awukCpKRd2rcNk6VzRONf35nbyvZDe0lQ
xjYllmG3uiDKuUiz+/jnQij/V/QRQAxMXzSXDFtPLLYWvEFHY9bfk10172pOb0cA
r1RMQeUfBv02rT6Po+FzUZ56hlFWTyck1lyoYACD/qMPAJ4+ODfaNu6hACz2b3PL
f8uEV3vkO3AAIQ1l9DRRxybeM53rcfVYVh63Afz9trkFUayLdIt2t3Lcz0rH4dIH
g9V/dCgFoShjaXf4hYhq4iE2pIU5FRtGDIq2q2J7pGLom7cg76TGHeJE2NDozAd4
B8GHhBSD9EkDh/M9chlnEohv8iAjUnLZOZDZ6YOUjaO28ZKm45xzQLjKMDtLXJl/
B8moBIf4qF4Ym+0+iLzNKB/59hxlF01QSXQdK4BoJ3xJD774AndThiCu47yeYpsp
5oknjUOeweyQ3QfBtZ2FUy74Z9NnZxNUWwPscs/9hNG4o+jHsUJD53npWto5nGG0
devfV62IwyF+5Chw5ZHzI7QpHofO8wjWwSm6BiWFllDcnNIGVcPzEbLsb3lyACf8
Qfrc7XWXrtXWBGyW/v76B1C9BU7TQVAoqqOIC+bzXQUEFVhMZHNXL8ueUrGoMX6Y
G3c1ryCHEWqxd1vq1qgeiCdUYx8nPIWuywkirYae+S69bpxy+5KJsFk2gdplcjO7
wisRf4Pw2HwGpXWvlj63hek6CprCJlfwKiZ/d2DZbdX9qniqtzKtLDue3Txl26ll
xZgj3w5/h9ZCQB80g7iX6tbA2/UfXcAsD4RtIMoWgh1dHjAqXw97vV2XVii5I3ku
iiVt0KQGZk8N6kU/Y/UbNX4acEbUW2U+jgZjYB/Egdf8V1JCVyQYfEuGQ0OavvML
020+B6h7RObXivgJDpzXFq45JjvkUMU+CDPzxNw9b4KiDvPvC6mFF5wcSUKb9gce
ZyMDKDnH/Wose+gGiDtE6yt37uwpbRgP5TFbTe4n6S6NySc+Qvqv197AoHByTLgP
`protect END_PROTECTED
