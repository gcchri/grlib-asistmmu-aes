`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ADXyyqUJ73lckS+XwPmACpsQ/+9VlrfIl6UImn3suehx5bSxSyzSoWVR9MNm5FG4
VKo/KiA4cZyxsAPfcMgGjvdGgJFsAghAhGi+FN352zVeqaQ8HKC4CZt2gK2HxiYL
xsJysE7dXIRGdjp9/vzHqo+afqspYfSe3oOzE9XmGRkYtc7l0WF43+0Yw2WUrx7d
BzokZXzvKoQT8srS+GEpwbaS/XdVQ5GQvhCYwURS69DNrnh+Blf27Bv1JssoZw0Z
baubPOtcNvJ+soFAJdfz4g==
`protect END_PROTECTED
