`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Vilsxd6JGXB3VuqzvMJAnfvhjbmvAPGMp4MmZuJxPfWFPKrknu7KuJcIUQv/hju
2CwET8HAp5tXA+p2I7JBB+9bjQoyFIfYBG9Br3N7+ZdT2CzuLRAXb8pv5vZG9icj
fPEMVEJXnKaAzyDzbqlnrrc+nyl77+wx69W0RP/+AqOnmACsq/JcIOoZn0f7Fe7V
a0j/G9DjRsN41TIGf68aqhXgO5SeS/do5uYb4AsjXoUMHQxepc2HpmpeumXeuX86
WQgqh/QNo/muI4bWdfOk/d5iIcH7EkTUCt9eROBwog0SVh3jrPT/wBgjvzuSLiRd
xBwbLsCoMp82ZZideecoGJx/PRKCfAAWGGz6xyQMUsm+X1Xccwxqh6sMiqJMv892
O8WtvunK12IF9DlE5UpV/P2xjfWGmqLeCEp9+wKfFl9LkuNvRwci5Pot+S8tEamx
KAEDcRM/UfahAZu6G1IGACBH02Ed2pxqxNFrhKv9pmg=
`protect END_PROTECTED
