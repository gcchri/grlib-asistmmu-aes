`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GQLSOqaVDhJVukbCBMXmWFKmUX/3esaSKX5/8qoNEgHHqMyyA5AAwb960zNy+32y
pe5GCm3tlYcWGthaJ8N6LBVBSoEsi/NGxG3WHv1PIZWwGNguBbiEKtzBbB5+4kEg
CW4ywnPm7gC7bYk3DZnih2FJRaEqOEZoByI60TSCg2eQRW78rZJnfHy9Ffl9ksZd
pi2CiworiZKZy2EzIQsYdbiDKXxZU+53/c9j9vlBlIPI6jBkneeC7OsZ2DFGov0B
Ay3mCgrnZm9Ue76QxTBHNPxC9ARNiHePNqldfA1GpPNwErCGdMVVAEjmfTUA6ZVl
KKuD8PUeTOAz83HScHklcvhJg7o1X+oD9R2itXXiZilns/WtzHtgKf0ZVJsh3Lnz
dZWpOeZc5ERjVRYEWcmBpTN9r5GmZQjbnD24LsM5gzQKdymkAjAO7yJ+ZJIxet91
XSR3+4Pkcw9cxy32ZVNGZkR7CgK30G/quqEnL8EpMa63/n0+aZFn5YYX724h8bAz
KkdbsDrS22xHeKNrbCxjtsWLTNduI4dPwgGRkZfTnNf6sSGhAXSnWqQ41xx0xVBO
NbrO8I80fbQdWH4Q+1jX7qAPSlB5Iezk+lycFK0AXorizrzsSkFvTYhEwnE9nVV/
MrGJ1b5ghp7YsR+eTAMM3w==
`protect END_PROTECTED
