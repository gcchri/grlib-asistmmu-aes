`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Amfxuu2xaTF4GxDmNlnSHaEma1jMRhWSdTr7IkVmHu0ImHmAG9d5cAMX4Sgpetvr
LbAqIoZ9pKtpJnqqe5qvnV//UIisuEzcD8H7h1WgeKJQXjdi8DMDSB6IYHcVUKgq
ASjOVfBpcFJ/1OyefvBHQo1rtza2ipa6XGW6pXX5GQu0KO9xfNNM5bgqgJNEZ0I+
5DzqUlH3BVo6OfgoNAljOzGVacdpgFbW9rADE+mrgh2nrAhtQouhgMFM0cFMxGfo
H86nkqbQM1riGibi8LoEUORmPrR35RqFaZKCubfx7UkdGm4weYHqIrVJr4keT+rL
alCMP0PuO4pZ2aZrMvEAC10JXVFVAlPKXbZm3OmQElF9nlDkIDaa5Iu7xod/i5Vp
7Pu8xyP9eb9m6xVuCDvhxAJFVKQTOpdwOy0cd8A5XvCqIGUdyBlNhyMnZG8oZUfB
SBb3+KMU5KohzKNQ1+YGKs8CFqTt8R5EwLZuRpwvfHUVFycFE5xFQTH1JaEHMvvX
K5AzboQ+lWFZ2/xVhMJtR+/fm1d4jp9qqgDSfHHqtXwW3fvPx9z/dDEwrCjO92aU
Kv+Z2lrlUwMzCLIWg1sp3cSnw5ZjZnpXq25k0TQM97P6JGjn/a/QALHNx+yPRaKc
mQCdWbOvH/SG2zuWFRb/4yI/qUpz06B1qwjg6GrTuMKUdaYOkedr+shERMeKmDTx
1/ZiO8Wpfyxd4m8FCql3GBY4x6g7bQS4y+kRfjEXM3iSeeP41V8QNZT93cztCUOJ
3rFfDBUuGGHkGK9uZBbRfJSjTYmaETVoE0TT0K1qrO6M+uBLn02P73nDLYeEM1Wn
yO5LjfR5DGKzTfXgIoJddvX0MGKzsjQ4tfHd/dqVizUsvxTuuPEXTQ9qyP3R7o3Z
9KDyvzHLIBUjS3A9GdLffKH8DGqTzhgOIcSsPwfBFujAXgcyga3MmGzDMJensTHP
u5MoSJ4cL+zyq4LW9xQtKCnr2OyReNAJ5Z6H4oDMB6zXyMCgMGWbGokfs+6I8BPa
15MP5b5ULE5+SuaWWTrK7+beecwvZ70bfbCDPiY7XLX4Ug3RFZfnFHyYBY23GvZV
BqeZZadeTprZt3LdlgTFtQ9FSqdRTXey9VBZRMJdohKgdKiPyxpm5ngx9tnaAbLq
9ul55xQvpGe6g/f1FWZNRSN1SrOBIkcLz+OMC5hSt+vGZtW9NFpvY4GZabqgqR9T
xNz6NoDKM7jdED2BGRd5okIb45KpcGrl36RHfIgyVnNyi8P0TrFK8dlNLWu0m938
`protect END_PROTECTED
