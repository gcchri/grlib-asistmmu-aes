`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lBT6+A+egOD5zLAa9x2YiBsQQjYgcOI54jA13adTmf2J8ymO65UUTpW0PIzKur8Z
kFG5BWAGmSKROwuufnvmxKeomE4lfIVklT/PYDEx9+Z94Blq2Nyv6cVEML+5XTII
tQbE/TQfknTTGpiaW1y3EhWs7Fg1PKqUbHlucOwzvkiluTGwD0T0BWwS9m013hlT
U6ELYcwQzGMw1rWPaDgxNzfE1MMxQswe1N2yfIkFXbCCiT+uu7VtBiXau+AKM3qM
ZVgfg3Ft0qyIDbwVhY2b1rE/+NswUF9Wldw4T2NR5yz5XzBKl5tC3NpOE2o7yFLq
BwESz8wZZCthJ5Et3F4i0VUODMoHxBsBcHTriNTvED742hyCjmVP6BsTVQ2hbf7s
jSyu+ZdgkUZBhtIYPLzqWY3p4YERnxuYieWhzCGl0D9Wlkc2G7JwG7MOiI2wdp8o
5vy8VSHg1j43qk9LE7JyABQXt3a77SExLs4RJk1Etn0c1Uz0ADAaNRNCmlingsv3
F3w73JdLo0Ned0ZBTyu17LQSo1p9CN19OKjQnxp7sa+8XGe0ezqNeZkLBC/GgTuw
5kisdph7f8lUEdpKJwMZJiaxFR0Q7N/drJsOfS+0HEPiLvOD/Pc3G3Ns5gczGpX/
d2AzU8ahqB43tM8NIbJlEs2fzNMjVgmaQpQ+Nu4TrgdZiECSNda6e8bPJSx2wL9o
zpKGb/GoRwtb9hieri91bSjwjAWq/SZkdbWT1bh5ctJhITGvvpRYVRYG7nH5VISg
5lM6xO2QU1YypQWaG48znGtUp1P/7KOXvHTBMNt1duz9KNdvnSTF7HtEx+ho/3fc
yLyt3HMNymWGpDkeeD7n3vDwD15yZu6jG6reODzkGXNMwpzYcE+lL2QLt+fTgfbT
RyYUTuqJlIGpwoVLXJvk/eSxeYpwpxQbEQMT9EiOiYdd5rRuwWHYLWbb0QvWespv
dcVdGbJLKnQpKyvZY9XDfEITumTZOZkdMCZef8dRg3cwdzRxS5k8nClzbOLaJbr4
KAv0G38oIFf9sCL391mRQ1qK0CaegsrNTmdJniDvRxFndQURvbyc43Swivb0rO13
bfJgMbp8rzW6zyRkXBCOuOgEngRFFyVtw7v4zJjFxzyihfmh02iL4GWnGN+BbPWL
v+18d1XUJ2QXRM8XiyUm3bsLVQnjCXay3zpOgfpM1255NOM14FBFE4yMCmJnYyuv
jx4Js/GpLTirOj6/6xQZ9eVooCsWUBgV6gq0dehSzJXPRyH9sIK9Xodbs5Qhhf6r
LHe9I30fK9Mm+gItcdmXmrargvPeDIcw7STc4M1qyYwUGmZ0r93Y2QTZpmgMgxs9
aCbTZPQsKq7jv/t0RiCCtNzYdW2bCqGru/mYGb+cgER0XiM+UuDIsz+VU9ilAf2n
pdruC+utjCkKTiLTE6MSEzmRg/mlL6t9XgRMeD62MoplUWE4iTwQWFYpCVOVF3lz
6cvvQzmXEiIAaXq0eTPdZA==
`protect END_PROTECTED
