`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7MZ2MTWn49HKa4VogeXJ/HqFBfZXG5NBvbKx/l+Tb4rUDnlb7v3eTwD5l8d6tzf
YFeDvBrtAIcf2o1WOOJvAc/3t0qniRNQgkhi8ieHkALLqUfNO6yaeeUm/wMzNmmw
Gc6HuU4UXkd7fzJI4IZ0f5uEdtQLMf9ANY9mOUhJn7uPCcPnflpXDcoSvf20IsIF
SoM58etxyNdcRyuh2S15uO6y+ydGyNBzF5dAN/3Z4SQjmCoODWj4LjKgfv1JMPKj
zSO2Zq7jtEk5gogxAf+lQ5XZmLdoq04OttLC831UzMMBM4qx2AJWwJylloqU4fJ4
y8wkllqDooqfRMBWmE2QH72Gxrga5jSoRGj1rNIXK/eEOPTs8MySbAH1OC1J1GLY
w6SuOHvZH9wwXSSzWpkWl4AsrtZ6x3NVdmoNSFcq6X84yaZEOiryirMMIpMmKai2
tvx/6XcIZd/Q2uN/+ih1ow05Jd/rnutytN1eDCF5CY54yrrn3hDYjnhAAQA8P0jj
nWnxaqwXi/hF6PPhdWfccHTJZgqXez2iD3saimy18JT6ZMeshTie5pkHP7LyX2oT
mStdS4R9DBw/lG8GRZqfwtbS0uiyTTKg6vNGVoHO87omsTojksrNU2JL8PYWwt9R
Q0sizcsnb2fJQOvMPnMTuOYTmxnmjRKUSIx9oDiCz36sQodjDiti6G8QENxAK37W
RYXCkfJc14+IZCjiEFudVvg2dyZzTgho++kb06tZAt+0q9riq2wDVjPUWAGmTEfG
ituFMq7kcD9t/jzDDH8TbTnvvh6hzSaiNRZhZQNZPAl2Rgm4dRbu4I2H9Y02J06c
v7dUTmu5Ii28YupMchd23DpoMMQPnrcnUskb1Ftbbuc6x911J29Xqb+KEVZ38JZH
kYCWAMV+HTiXqoa2mWjfWfyYJT4uVnJVdKb4040JRilRVfvqfdrJSKxIphWOI5D9
raesjZLL10QfwjOeN1U94udlJ+KcqGr/I8OdeWZQLDNtYVm5B+Zc8CJxA4C6TwNq
uj+YeJ7uk+bmHGWbu7LiOfQIQmXt1ohZ2iR4sH7mCKIv3BtCJNFUsbKOQNK+QMI3
5XocD98UC8LwV0Ag7dBqGvZVLc3nCj8qWJ9gz5N4GZeKB7b4d1gA8CyQELDbVSup
PBc57wkDNMRd/zUq+0hU6Ni6L9JRTmvBDUu5KewjwN6SEUQm3puBRGWuECF0TO4B
LpiAX6vQCwl9PmhI0Fg9aom3qn1KmIYNn4kR4xAbjEIga3fa+w5Xgo5SxuPcjajR
QD6aYMU5MLyRWD/l2tmO8Blrh2CNQG01RGVYhMqdPbJv3foKaLbgT8xATDvwBQBn
PztpG6hZYsTS+2Uu5+S4CNCB3VZMmK/9V6PXM3wJOhmVOYBBZypMHJS/xYIvQ9Yb
F2NgsieTULFoRcIdhi9Z84XV6reFhKGruGAz1NqMLvOPIzpV0a4GWT/67zmJV/N+
G29EH+/3u7xSdYQHk0BO7g==
`protect END_PROTECTED
