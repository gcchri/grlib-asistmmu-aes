`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jzQIrMOo/JPzM7lNbPVlfWkUIvHpChjgNKuYQxRf5IxIFXD4gC60GAWDfo8aYlxi
s6tkKy++STwH4tFY8PPzo0SFIlWYc2o6gMh2/RUboFPfryVIf+mvl6QL++8S6j4a
ZjGoHTJAHttHrenWRa3/pCVqsCInXEi5pRx39z+kAHw5ZbLea1gamS3En43YH4tq
dyGEQ5YQpq9XdKoJSCYJts65QAjLMzmtZMPXOyz6eEA3zuOMhQ37M4pS6zMmRLvO
rsxM2QyVDAh8L4QMGt/1soSEwCz9U+t7ud9I2nw1gAk=
`protect END_PROTECTED
