`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D2aLgJ99qISbv4o4Zfg/3rFajjIBVFV0QbyLhQ4h6fgoKmCTBY80FS0s0m0Qb2IU
DV4DPbHulmhuivsa3P5BYuH44gGVEyRc4nnm8d7GoUNN6O+Vn56b5NvuLBOWCf3k
TVEvkn6uDnt7C0q5EVtLQcG5EjyjTEBWhvw6eC0EkvWTfYV3j4rxXkwUZdjdl2Fz
a+FG87zUGa4Hgy4f0LkF1tXl9Vz+6snMXMc+uSw8ha8t220MHNeS6yJFQhoJF+vR
kDMVLy/AN4wQtxmuXkkxKpfLtHctOexKkHIlTso53auKF25HFRjLBYnOel8wpr/i
nztGjXDcR48FOrEQvHlcvlD67QBzyzpwumm3y5yWUELnbflTa9utR4NJVLth5Y7W
bBu0iKnTnkA0VRJVXECcmSuGGpkWIPYhv2Fy5vBqV85RnVHPMrBfpjaOmjPhO0h/
p608Mdq2dff8eBB8SfdlCsJWgUBgTlD8cDYgJmGMRSxPnt+jbrH5J6JzQ0KDhpxv
4hF9E9GcmHLQwli1vfs+TQ==
`protect END_PROTECTED
