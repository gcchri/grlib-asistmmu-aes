`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zi9exwkuM7tl9m2woJWWshr8bq1hPD3YSsX/gZlNX0Dr7mGN8HcRiHrVp3zpqFCV
BdhEsZU/3c8Lar/8jNMMa2XvcC34fhqPknOANFjIn7XJsUCNu+jW7lUhRB7MAs8M
k2sw38ckIKg6wJ/wKSKWxSEGGIrmUTPxA6mouXGeInVljjeUCEz6S8vYNgmzroQ8
E7rhS9fTgX4SK4uoDRLGmLeO9xnHCIDHbrd5Z8eChhVDPSztS7oiV9y0qVqYiPlW
9GlPvPsloEWrgY+nbQ0kraMRNRb67l1kk7NqXrqy2M4aCqetZ+tbTL+hLBk09kGP
2hc11R756LmpWIuKA97C0g==
`protect END_PROTECTED
