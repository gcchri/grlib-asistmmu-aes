`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NVfqk9lC4ytL0VAi1VVyP7PsRL4WgiZDqs6/wO3iJPPrObUJ0gQcq3xcx6NRiXFY
jGNMMa+EWPENZejmiZxChu/Lg//fEDu8Uz2/dsOJb1IuYwKiV1hAJ9WMxP8tjcT3
ivVVqg+Cqz9KJ0ke6iKbryOyExagTFT2jlcDm7DWPI265LU3+SUVLf9IS2l7kTVu
mJj29wCCizr0/6Ixzrm/B6WIW7PlrtJhBWpIznsTIpOJgaJ1vDbxuRQKgLeqbRQX
vOVF5uUcpv8sOviFPiSyrB2gB2cjxHflu8LgOQc+o/Grs0U+fko0P9ux34LXrRFu
nzbrAHUuYOHazF2HuitSegH3xmD2MHPFY4YCRJ9vsmKGUUGGOqifB7Ve8Wyoeq9l
8zXE/n1T8+bOiYVrf+yMj6UpAzrmmLt7WD2Z2IyT1rOroLC00GZndgLp64ckoJ5I
4TEZmNhh412lqC4JtIFhNXrs+pdpmkTb1vRkYMDJggES36pZSOAdXAf2XSBLeSpw
8kFFUJCfUeVUjcHHSpvzSMSujop3rdlnR8NIk1oAwbmvnDFgFwommphIMPZyYvKF
v44KYpHFZmGKXUkqtwhiSdH+59k7jpmMTOa5aDiChgUtY2I92VnOVZGZj6pMSjuC
vHyGJjkBntiItvXV/wyCDwCmTwhVDbVwKXRusxssIbj95E0ppfkAEaFH9valma1+
Uih5YHUOpyRf0mtfcwSCnBU7SPHkn8lmO0vzwCboCxMBQGO+ZvyAAMzNoaTF2YFe
q0BINtuV/FW/Xoy/W63lFGEnXGn/Mv8lmCfHKjcjaoWPybsHcOKI/ykumh18rSRA
4CPiOYQPEQIO0Uy0sCDWIiupH9kvuZZrBvIIRbuhdSwdG3Pwws16kcoZkCKkRYzV
ocrazgBmYrubZhMIn7+5Lr8BghkkvKHmRXD7d9hHzgrQqTcGHe1t49MzJiNGP4DD
BAfjJ8xTPpLE/SAJwnb77WJxct4pD0PA5lHkVoA6kcM2Gnssd8mLLyV/iXlyPCnE
+Vrhx8TbdghUuuZyarVkRCBDOdzLlW6X2jc6JxcKkMd12Bb0Vs3Lg70le236Dqs1
J4Jnc2MPHeoQpMcd2uiNwtqKcQhjW47L2Eizusgsh/AI39F08D9wMZgjUxISQfcN
kn5zmtuAiENa21Mxj0SBDrvuhU0CrOaH0lPLlegMEzEULIhfQMvqvRiR+t/jsJG1
H9ip4ho7KUG8JSwsckKUDzojQYetXSCK2RmbysQ9frKnHM5ULHIiCuOUxSEwmYiv
l1Z42JMrCBnuuI6YGybsQN3GYn/VQLmZL1nGYMkPQZj8jSd6wNtzLg5g1A59FoYV
vB0AR7Evs+QCkdoms72xJLpfHu+lM5FWLBqUJsR6OuXskX+/X6e/T4WsnmbCJYSf
pFwfWJhJzTipV5BZje0x1IPA4LMQoesQsPnkdEcPSSdMoxGfDGscHHfAFh9Cq9Ay
loRuYWlvr3sjCpNrKu8ssDvEgUirfkkweRkehLBmpowkEV85NuZsWFQ7ETx13hGo
Y1SoMIV4I3rD1vm2vVLlT7OX8HFnsD6spgjIjgS5yxiaDrqTH5gNVVs0Rl0XAXVS
biFQqsShzTBkEUAYZ/cRMk+TVKU+HEik0Q3JhwtS16stnkgZVnPbrM6sdly8z1wO
mNs+6zK6x0STBrRKRa2zVSTiyQk0oIj/EB2Uu+vnvExaVZCLOVs/ODoOgL2PbPlA
lzvvKgueDeKuJvnbTE8Udvx5BpevKDNNwP89zAMFyE7bkjc2Fayf0d5gr6oj1BIW
etwDNbu+YSCyHunDQ7g0P4uId4FTHHHmax6KwV3VMgEpO9tFtYZU9/co363WIZOC
oMdkTiaDc/RDMKvYX0vB99JfN4wLSH2id9RynhfuojMtabwueZXzFFh+/ffWtWNt
pOgja6JPUV+VMQKLL9vWnq+h0/ZttWFd1B2o3JHHRNM6gJaNT/kD5WPqOD6btQ9w
xrj5LiNX4hZ/hhCzogZ+Njdwr7HSI1EjfjwzjZI2k74A4LEj7RKb+XYRyuYcZgKO
6fvtQ9uyI4v5nOi1mZSEFSOVqSCTn8eWse9iPJERNksctiYIVZ1utjuYgo38ULBa
jWJvbQ3okg6KUnh/M/DjkIaRSvCDRh2sFTqhsJYhT/R7GQ/TEN+KyjzmPvm9V9U9
BAPimrRhG/Z3SekK3cbUUgHN4I11Nrs1MILrManvNniG5hkIF4B6tJ1ko7a0GcnG
reEqqy/Ww3jjgPaVm+jHpO/+aTC030lvATxZZx2HlJaXZMDrzrzgzJhC8A+bE1tC
mca7tJGuEvXkUFRx+L22BYlMO2s/aPF1myUomKNB4QIUj2nOLqRpOKvZuOsPg5EX
nY8EdUMuagECETpEBz6gulcKsr5ki5a9WjqvK/XAhOU=
`protect END_PROTECTED
