`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8vDxecY5zriircyouR0hJ/4eR3wYKINxvB3rt7OMKIJGArgN6RO75Ke3nMAlI8f6
C7UiiVASJnRw6O91HxkmjXrYUxsj2SYphwe0jmx90Rdv3DEzmn1YhkKfhPX6O3W6
ZIwTj5ifdQUaR+pmGKtY6HAhxFQxAPIpvD5C3ad42qF11DUxnRgULJlrMkd/2LtS
hhTOk+M1Hs/O6WSr8lhQRkdonNjv1wLjy/v5qlicdQeShLIr6HWn6p1wKKi2EBXV
oMbFbkx2dxo9L5Ufy3Pyk+AiBYUBqts8BWVuSdtbS6rj80G3ugwQClb4zOafYdMX
gizXQpg978ieiJSEl31Jk9iVywkUr8dYZrdcp//XsdRotNC0XZeSLADbCh/XYrCl
CWum8zmkpt1Gjgrf4vFHy3fr2y8bNMeoSC4q/ZPb0tjGlfQThICpVcGJK3XXUZsR
B5yHjEM0nYne7IAOGDeimo2ZxnkSfGcre+jdJtskYGQ=
`protect END_PROTECTED
