`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Em0ifLuXZxRT7mCCbDdIvpmtAVC9HAbvzY1EDWYMXRqlH3VqbmIGtr7p6Myrw2Xu
fafEwKZ5ZAABFSqmVbb7KMzVgG2zGgCipsImcbobnG/Yc1Io8wfSr15UzpjfutjE
98fq6zX4PbSJxeoIvSC5MT1jgaTBSSVny+NlzjVsugWK9TU87RmgS6jMFq1+0IiZ
P6z5GPyUjcbxYHRqhlIN3SqnH0ciQCuLj5PzkVhLCD9/OKpZqwniVRDFAoqKS8OJ
OCoh+C3tBEKJ8KdkmXIcta/K1VT10/zklDH91kV37tHGU1L+NOc/8zMwDQ8YhrzO
3vW6jFtoep8eIsM4mdMPe8WogOnrbV1DeEUz+PwjlEsx6PVYnWAZ+EbqqcgLXVg+
gNxdfRcZgr3datYotEd8pxENZVAcb04tSVI+6hBY1UtiCQ4Jpx/1j3Hmh7P3tHJI
WMCeqqtTxcGzKSII5wcRwrxK3sLjmCYPNmobpx4cTs8DrRnQ/kH5qY4mFFQGhKuP
+Ate/tDxNl1ZajUwl5MnSmhcBffXW5OAjXt36TP6U90m/7A9aeMCqaUrXEx/bN3Z
4vFmezcidZDRUd8hG83FOk1Qnzv85LtKPoy3SyaEhP1wJpku66tia/QZnfbFnYUX
7YrbvxK8LnC6p3m1njqIBo2E/pVJNu5sgihRtuTWmuh1Q4mrOTxywBJORYfEMCJ+
lengd78ma36cZynRrtmp0L1VHUJmtGPj8cY/CvuZszyWv5MuZrsUhk9RJFfwkRlg
rf8Ds8MrrVrhSAChhb5lc2XfRjvPjTrOtvs+OCmc/MnLH3BWBhazekSKdJ3cMnUb
7qeCs9FjmiiUq+HLopKLqUZHfbgvCkF4A7sC1TkK38wsdpt/sxiOqOZ0WfHBzN3h
BYLeya7qM6XZzqwA00TfEsqtMIEZGQzbBH4O6U7qGmGqrGO972vr71qop8DvYvTq
XkvEZTguHuaSWBI6aFfzQaKEu04uqd4b2FcCu2V8b4Yz85c0VM7hGe++SESy/Vdy
1QqFl00uLPaJ39axU5tBsGBmP6Dm6Ct6RnPxz6HQeWrxkZuAc3ZhJviPX7WRLJmN
b75wyugmIIRevtyAzXeRW/ytpl6+jlsuqtQYBXdZNMxalf6M1DbEVPKm+pJrl9vY
OCIhsyyvZCpT8FAxaVD1+NV2XiI/RHEAIXO1rFGLOs3ozX1QOBBwJaO7oSTQf4aZ
a2y3P3YzN4kcAOsf0EJ805RnY/R3m2PgQsZ1UpqtUYR7zfEY3EvDGKBOO/IQyNVI
uAuF5RfSrQmJt06/v8BIiRl7SUl2hQlbcnDNBvquCyqXXUsDLL6jyhHN/8Dwwvve
FcE53Fso2ZkvuxqYJGI+iiMcrBi6qDUBvTUaIC35y0GvbmMW62QtcNTn3l/iIXH+
hswo3zO7g8CpkrAof6ruSuIF5i6NiHO28ovenHeDOqBTGLulqPmOAvDdelZcbL+1
rUFIvF+BIH06RVcbZx3IAcsAETSLjs7SeJDA+WpexW2D8QExQj3NFAf/LeUoEv7v
8wSauhsqTOyWSg9gqTQXDRX5h7ZdOVV7UdpkQEkDhU8+6bPbFfPwhz7A3ooYLXPd
CQOM1uGRhspfB5PBkT4MSnQpzvS0ZC8ZX6pgOarPvRsF3VxDpdD7xm39w2LyLbPv
VlhsyTK63yqIidZKVNep9F6GRjA377OLcZRi9Xjx7Z0GE4pud7moZamToqHPv+3I
h2luF7rqRSg/d3sSAvM2hqti4nOCi0azGyxkpUHh3jf7+nIbN8rbFUeOAJIKO6Tx
qp5GMuw1sBqg67ExkM5gHjVeMjTVYIlLX6NRoHHO1tiSfTFl1veY2fg3uiuurizZ
6kAti2Ljq+m9P9jmNyAbQzUHOM52/iem5/Xr1KkQXAsXy5mSlkdVCNcrQpKDXEKS
EGSStWOj6duivhv+hL43UTLFeNPZIdhF6K2GEAnve2htKB5hYJv5U0BvFeVUY+9S
9l7/Chcy+LnkO02smRpNJn9iNpGG2Ka8ARIAkambKSpFcUkvVdvPWpkwkXQO01Bm
1+iMrMk4VIyPlpCEH+8eN/nz0EQ22XOb9U1AhVZy6ItiP9ie+foSRfCjbo1Vo/hg
IoKV0rNxTmjxaTK1m+z+yCkYrE0eRETpJNj9JXjkycMbbghkdiFP9ss/3rCPCBdA
pK1gTyvO/pa8dQoM5PaJuuk6y4Q+VWlpBn9b44MMDZDLZeAca04hp/eGAyWD5EPB
qMql0boWQrESPW8xGYfo+k/5cPg1b51FV5yZmRrvLbFxGJJPSdWA7cuPXePgiwQx
UiPYOxpHIoGv+7UsL4XssHWb9KbarKEnS92zxdSrFRv0had0Co+TfN/vbsJ57osW
Kek1Btjub1I0Atk7BDxv68Xzd1NYjPf5azVW9mYdXHquWBSXVMO3U6fyu/R+7Uy7
rsejPVwH3lCr7+LADcgZ5uGwXrqJAVUXRPLUPl7F74hcAggh3hrLbxZN8N+NE9Ns
QvlyHUuVkWdXOYLx8g6AnBvQdDsFDt20kGJpkddQUoCpxk4Knn8+SffMEwGjafvg
+01V40NWAeNe7Oh0oJN8VNKt0KfGfp9kMH8Dz8rVlUptD2rhudPicth890ePBmbL
AY9iLCQmBCZUmOibOsLaTeuf++44aiAfNWn/VKHGnKANVvu3tPaFPS6/eLd82T9Z
a4eXBAFN08vMGWtQ1vxwgASBt+ZGGQabkzuvpD5Sybx0mvTAwyNyZAuAjAsE+oQe
ywCUh2kYePDyQfL/qHk+h/v5g19cH6Y1ZzhbSga259wnEVxgUHloDJ19hS1OSx5k
uXP4uJRdaaTcGqL8w0I6RPLGQeMPi5s5gyJq9cfAgOLNV90SyjwfYk0nU55XWvuq
OthZIQnMViWooqKbLRojWV8Fuk0WtFhiD12BXuANw+gLCqIEKD8z0YyDjHjbO8KV
Z2PgGyWRVaLLFLyO05DnP99LW4Jl+IDCYKDT8aFJRz3ufLAP8UZF81ZO9ruex7fz
G2QjXe3SQKSX6Ta6fv4dGJ1bG3tyPzfrKzb49XtQ+QU6lr8n83HQ6PW+BZOnL1fc
ST1S+Qwta+nqv2zstOXtF14hfXcZm1CXn2hPPR6OKN69RpuYygJD+NMmykiDq9ZE
qTAEVOvR6X+mp8zh2X8ENdKAaTbsi4/mgzGTURkrWYcBnhPUvTRVsSTfFfOn8XYa
WZ5w+GartDZwQ2UUlM81P/vJ741vKSCTB8UYRlUh8ot8u5s6M+nbFd8Nkys3azBu
puWuKc0ocbBma6mxjPfRJFx33gn8YARnbjOTrTHWTSz9PhcWjR68T5OmnMu48V8O
uwfvaYlzEhhlkV8Dxa98M7fQ/j+TfzPUe8fvOaHVNop4TkGcg8iDCOQX/c1caolK
CvsxPSoH/g7wW9FDBH5Kf/vefNJKMI3Wpg1y0GLsIONf1kv9nUrqBY8zzqrBCgF6
9l2CoiIUMTLCcs6iZf4G3hLHZJECkdxJ2/7EAB49Js8cuNtYS1rKDkNdx4Nvilga
TxJw86A2bSrynu0ecKOOPrXBcZXyQZ/8wKkQ7/RM+1gJDktDGSp8rtRiLbiDy1+t
UCRP3SAhNXUpmmqHUn4/5K+joh5AgQo3QnyCUacea+fO1uWXYyoZmMtIXd1x4fgs
mW+ZaOetsWVfp4OeQeRReoJj/TqaeH/agcn9Ng9PZR/MhF+DK61s9WX9GIieAUsG
E1pZ4wXyGthFileV2zxXHnIm/pmj5eiSKYDks+tavjz2vvMg3KNbjCReykxEiVK9
4m0XFnO+9rUl5xjFm0732mezFo8UeQ0biMLDOTWG9dbXm2wbFgEBIKa2AxEPpxBl
uCwWbK+o8dWuzpGKw7A8HxaoJV97WAcSHbx1xfSMZdsTjq7/qhTJEOBx+IJsdAWd
wjcSWAzDVf6Vj0Wc8DC9OH/pyi9YmvBnN22uK2+/0hULKiZp4GtFPxzJCAN2VTKl
YPIXrZEvnluKdz3/KJg4oWxPaXU288HfhqxiRDTlzeO/5JyfViFWUSjvp0r0siPo
/MpPYYOZk/z2YKRnFTuqCvq3lZxTINmeLHw5BxyEgwiz0SkGT7SmzuPHUNQRHzbW
E9V8AdRoqynGzR/6ch+TQbzBwNAvTzIBUPnnyrtTvT9yQPL8HcePoguBeUOftMfy
ctBBnUdx45KDvafpuPSz2OQs4ptXLdToVRGGsEaMY3XCKWCYHsXR9NM0ruvAN9le
9GqviM2Zf1prx9/Zkj40iedQsI5n50vR6qynXzdq6nATq2piiIIcDpDCDgwNVjOb
KluyNA+FO345UJxT54se3PtNFx2niRc91t3YNwqBYndnz5KK1nP9fp+PCujo2l9f
f2F2d43/1HGqWYwXd+1g09ZGPYMCyOZ8HoD5LITDeoArEGa8vkXmdVjmWSVxa2Cm
j0eUa9tSL5QXPiYi9dxcn03f9gfsHA45mPg1WLXgD+wiXXJft7TkqvE+qy3UHAMp
CusF7A4+gVoi5gOSCkKeyIjnPsxrHD8Tzr3cW2vM7FPMifv2eIygA3jcbmTvOYKi
O2uFe8OZ6QX5FCAoVA4W0JG9etw0i3teUCfSinXWW9Gy5jNAKlYH6AM6tUgGsexR
bPZiv175M4BqIT8URZqCRVpqP4q+2hYVxrp4gsWau4QIgkAL0cHN4LMN5YE4NccL
gXllDUG0Jo4XtqYrgOYnEqWI03QlRoblfPrZUF8vVT71eRMjrIZay+Coqt+QW3ij
2yVtnqNsv+RVqdqP5Cn5dV7Lt0h275xOCEs8Llh+P9DSritKm2nVbwMaVEXIdR4J
CjT4FPsIGfwOJICApLeUPzaqfqkuOov3OjB1rhpSuEceGv+sl/4l6zxmgVIdxUtp
0MfuqAiJrfemm3QrDIFRCahuJC2gkeg2e0mbmjLLYad+UF7IeO8hvOEITozLSc3o
kX1uX+RQGfshva8vKccPiO4iYxDvnZqMmnsJda80pG/M5/S1ZCNBNGTkiHsppCq2
vQnO63lTpuM5KOrkhlEmlRyXDOTl9kiQvxiNb18w2/yBH4fMCmESjWpidvho5wI8
kjy9caURYYJoqN3TPgiFgJ9UDuazpxcioYu5+iO4lfecF58n5tXUHkvsza+4GW7b
WgBPB118uYo70ENaB07/qFFP/8KE3c91jDvdwFBo0GO+em/0qDpZ6KJZlJaXB4gy
r93IlgO5G3Mk60srvFRErHB/+poodS2RtS862GyGi6J0BOPAP5zzElc9mfLEnA87
0b8RJqIsYMV4aItQvN7IDp2LHjn4xOPmrLKMHbLk1HbHuUHW5yOGlNZDymV6fHLC
nekFlMlMqRspxV49CHpDCSQPuTNppNvJeVsNmph0VKS7B8OJuf3SL8Z8EJWvQ2bA
ZlrwSPygAzo7igZuDxLIZcuFSc9YBMiYeinYbPJnHNnCdquiYay8fsIrgdgFQf22
g1fJJeZlsBDorLOI08LEUzkOGIinEREW/I5QmX5j4U+3WqZOi2EvSopsF2EZag6O
V9EeeJW0ZljnevbaYG7R6v9GyEee3aRMXI643n6E72UEFEvp7s0QOS777QVrGv9u
4kpeHR3r5RkzPfEVk/z2wntt/sXSAmGRlFi7cOof4RaGAV6RXDbCv+gXmAETVPxg
of6j9czoePGO0HT/W7tfjANtW1vpugDZEpETbegotbMdsVScLeRNamvWBCCjLrte
bkFsf0AepfLtG2tv3qgeKEiLArnvu2BdLM4nEb2iksuMTcJsLdLqeBoxP7jPM+TI
Zfzy7dKgHoX+YHxoNd/JVCnl5pgDob6Lsp6ukSF0sjqzIxzz/emhW6FsUpN70pnz
O6BdTcBGiLf2y3NxKOZ167w1ASrQ4Eq5F11IOb0R3mUvr0k68XjUF7pGWD8iMsfy
7cCeiwXzfXcOcaohA6BteGLC7ocgXThqSdEgjXqx+FzJmou3Eq13KBnrRRzKMWNu
6jG5YWTt/Qsz1cag8lYF6XC/0xCE+6ejkEE6CwKf2gVHjbG+gfL5EOIu/NYegJMM
hw1D6QqMc4YVLqKMEFb/xtfE88+gC3aXakmxo6WTUFvnqIEsNuDM/P6nhHl69K+j
3rWfiSbPQoYcMJEaO15AoEEAYsAG84bFdl2rBuEDb7XOvker3RPIch4I7+4pCCN0
aiOauDtJZNZqJ9i9fx3h4smp+0cWyNfKM4qEUuqdu2lQYnTOQFc38NX5S9Y2rnRc
yi93YnrdSw8B0cNh7VRGX6dcmdW3TGI1VAqnDeWanQsY2PKcY25Y2hjPJ7JAV+jg
v95gRi4YRANC6W4G/xGEg+booiASZw4D8rzS398hTIi+XsVY6krSTbbPxfsAu6RE
fBTql9aG7B0+ohklHpwoMBg8vVkEFo4fom7NXUlJwG2fHRXjD+RGW7gFy0IAjxCm
vUEEvP93iawNj10XFz3o70UY00pPvAgWdHw91ylV76pen7xV9aCfPZAeB9C9+MT4
/HS+4BGBtgPqP++ax4T/fUpBq0x8Mc43Yvpp5wYVzs6G+BTzuO76qr43SL01MQOe
fpUyJMF52SMlsmV51B71yQFR0Y8SYWmcQtgEq4EHuv9CT5Fh2mqsm0pZV8UTjbRZ
FKsxBOOeJTD2aQdb07tmlSqrAgi2u8K7JvcSUTEY9H31npppHa4bIjDhENqTO/Rf
UeT4T9sMBOJ/LT/DRYF+OFQGjhOKmDJV+qfhDvzDPZh5nPVcgnMGud+GnPaIiOQI
hPbA9UHKWso6m0ZdLf0s4XpOXyycizsymoUd8oZIc0+ZoM4Snk4adX7C8GW7GflC
BOmmiBcgsmn9SW9lYHKp5L4USxLxMSHwzmr/cn5EdT5yVTf/b8L9tPcTWZgo1RC3
UB/hDgIMraDf3NRzzy3m0SkFx82/SS3rVmM4oUutDW8+7e+YMrv0w2wQSm2mzkIn
QQtS5yYsmxb9ZAmgraPwcM7ZrvyBsibFnDqD1DflygLtoGTPb5LrBPzYvMEnqaDr
Bs7UQxhjShNAHXeUYBB06HkEHS8/oQj5sTWA1EROSPYpaWLZt/6wiuhauKv5iWL6
uj53y09xZeShlcLgtNllOOfUveo9RmhPNTyW9r3+qrSO8NKNANKgm5Nhq14gOwlS
hjlL8K4iUGfS5CJGPSzWiJXkoACZ9RdZkeUv7CS58E79fNym563+Ce9hu8f+5bad
y7OIpPJCfdWp6c1Cl++tMGW/uYy4I77tYUVPXaA6IXua/wjUoL09enl8Zk+0SNOn
S3xwy8Rk6ir05uWatud/aYfkxVa2AtvWxMlWXdo2RI/rObdbw6Xsc6TwfsaCqiAu
n+8JXBIEoU7jLiRGL9d/Odv+Vjh+PwauJxfhmcmro8LTGySRJLOUwLwcDxqkw4pd
yryYxpgswnJhrDhcrzjsEc5x5KE1Y/A6v5uVZ8Fi9l/BiHhiFVUGpFzjBd+yUSxY
ss9F9xdx8VdyMbLFWemJfKfSoONf1c4KZfaF7dypunbD6JGJI/WSLT6u8m/o9HJi
NEPsx83RaviwlPUtD2kkIvth7NyJ/8l7zK2ssbMbMSjhUzBgpfbrOJnob0JFDYd/
x37isNBiIq1NqlmbWXtiB7kMbpGUkPzWkEErf1EI9VlI80SFETIqdckQww1t8B7T
AwT4VrtxTTLgOfFyZMh8BHO4E25TXpFtPnqmQLssQYMC0UUF49i6DFDclVRS30hi
A4eU/I7KsiwyPFIGsBIAWEM9DLFmU+U1/7hW3RkaPr0rWCW2Y0Gu+vwT91WNvSL0
CwynrXyntWs4DB7z4oabIsBmsSkiwC1KSDllI+PfTRQT6F3nbH8Wh4ZWunIsBc3i
g8ut0qu08PMZruglUeekPiuCU7rT2jADBqVl2xHq+5mYBtdp50+T/puxUFUb0WhX
bbsCPvBQg0QV9ZTwZTB25JzWlq9FLIp7mvq8DvEtWX0KPuL44gBB5cN1BTiLyn/d
m58R9FGg5J2nyC/JtzjDssAdMFjijBx5ITmVJ0H2V0HykkPxe7OpLrFMAuLEoJOu
m06gLtrpzb/lOcOuGE6ld/Fo9kiw6gp9aJbgcKzb7jxz0QOuPdTPJrkn6AGgTQd6
VHQZG3SZwiGafjBbbROv7m03Ve9i1iujmmZzAqmd/iHlqV2oBCoDfqIdYv/Ahvs9
g8aJvsFdDu0vnlE+p7lKSVSZ3xbiqUDwQmkT+CA4bk2S/VU0ZWK8Llo1caY1yKnN
36hZplcnLSQA0lqep/dd/z7qYZPmX2j5Fadd+1e1f2DG4AVkmUlL4BNTg+CjQ6My
174Km4LQD7oxz/reiUkR0D/oIGXJCRCiKtjmSVKejdij1SpHu04isUavLFhZ12ZJ
vUcCNQB+3poyPVNzyJY/UftTiWKzUkyDZLlayYrDNfs1A3bnfpy56rI086SSmFRl
9gHLiAQXeacUJqwwXmW1NdCvephJmT1PAc7Ee31NPggCPR30qOzOQmRedeoClXBX
qbecA2cO+v+5TSup6OdzsIIToTRePRTl5nmlesUCdaaytVGFPBIxbE9sjNY/bST9
tvqGOc4ymj4vPR/XmyZhsBtr4w1jAHSpVdeOaaeXKhjUS+DjFjijtRtNmqFnom9Y
soHikqxFccob/SYIItP7G04US1FVGcyP/2/2pkEVwKpyW6O47Q+HA9I4QNyM8jPc
9mWyrtlPf8fIFs/OiXRWTdk25aVu4EcG7h3Zmr8T1XhqUwsrAlO/sDJ3WsGq9449
PInSQQH5QCfZ6QsDeRGJRN/wl6Iti/SyLy/Sq4GFZDZXXO3G/pwR4L0f7bzKi/rT
RgIX9030GKGQZlLszoOyqrS8Fm3SWc53xq/5pypYfMMYcvvzA8tptiz/B1T6N0yE
84MUMH7bVj44v0ZfmPvEMzdA4TPN0ztaYyKlNYgX/bqqdBVaBS52E0mq4zM4lJMi
0Cvd7Pn1S5NJDGoFN3wbAfd+CBuDAUrE1t8GwdxsYgZfpXHa2X/Tn/2G9n49vJe6
03C6soa2VJ2VGMeH1q67h5BQxOB2dYXhpQiEiuDtTQCbwvZ3jeoG6x5doyyCNdtT
q1JJvZ7P1v3/9UfLCOJ2DAVmCTGy0qlKlS993Ax8vg0yNde7KEVZ4uW1Y5bbdCsX
E5fZFP5DpcfkIwY4V44w0vjmljXV6rrfCxFHF/N/B5ZQdM1g9w99GIgyDBSVXf4H
munjbFB+x+Y35soN+0P/yQ8IT0bIXc9gsdufgK2QdLPtUt0YKGGBTLdlqJoNcn6p
Dz7mdNEVO84IIVXs1YVdpmhGZAhdxnlGmXAfh9kVzExmfW/3azt7fXsRJ4D6IPwR
uCbxHO9woojly03M7Z8nX8l3fM/8cLCaCVbPiOIeh+Ihq71DVXq9ftB+++/Lt2Cc
0CrinYc+PrX2LuiHQClOyJPFTDtS6OULzOSMCOnODf1p+eGZA6PS8fW1WXo6EXa5
67f4LqyP59FBy7eHUCo61Zd7xBmFd1wAdxSUrxgXHNdqQOH2L5/ymqsUqIIx/x1n
ms/3yQnVDt/3UTi03gtsbVXXQgpWM7q+ziEJqcoqlW0O9PFGbp0ObTNAo5M8x6OZ
CuzFJrvHG71/8yHD/knmWenxRjYBBCJ4ZhgOI9lH9TORNsh2rt07nbDhCPC/M3C1
60RDJ0epI1F+g1lTvMhMuKnansrfqvfGSbsQzhgei0X1r01846jR+XQ+CIp7FtUj
2drkfcC5vHjucF807qxIGD8iu+qlHNDqPxyCEmJ97TB+oGHhFwmvqSnQSL3KPvWl
PvLkj173EQPz1Ow/zDqLFvfS5tvzLJTIoaibSEWNoG8fbJIZt7bwczfV89Htq6OI
29xsNfckxEzs8TXCW/yXQoRcM51it6tUOuGAsYk+Am4qGRjqE0ikMcOZwOzs43D/
jtmZtEguUjEpKbH968yrH/QwVLAt5kg5mj7rBM7eUI/B90XO3ugjAWU0c2UNS6c1
QvOvK5X0WIug+kVQNi3RpJonVJ+nQ97SgM/qvSTIyiP+JrnCwepiPGcLd/OpRaQa
3vQW1IByzgTevSuZWpoEugYS/heM0b7/ertjrURN2Rn7TMX9dVq8vgsrk0a0xB3K
zSF1sGSUpgM6N2jUaPmkrr0EmQ4EDDMwQQAsnW5n+FsF479L59kyNxPTVswr92dE
ukcv1YBjf4tEbsHX2Z5se6Htcf8/7rW0QSAKY4OmHnTRv9T8tDEXgMrErJ+1ywE3
Ov4klQipJET0xx5yXLsQA5iQDj4OkIOGI6dnTtOj/J0MHpnrxBJm6kCq+s0V3rtf
lR4a8gd50nd3m2zd33zNSXHTPGvQvN3hxHFA54MZEjN+L0RHBnZ2GgmNNaesorOy
DyLZKTgNBH+PfxtKCEI5jq6QBjMAY2tL8+aW4Ce1xG2qc7+jQ4ss4iiMsXk38BOp
UOZ4PEhdge2YGeNs2OEkL5H5uuK4Oi4+CfOu+S056bENGgS/ls7DKd1Hxtq7dtPP
SdA9CLxv7qKSkEp5XrDJ5yEzPHqogcvDD57tEefk/rxTsoBhbvvZujSH16eSXeoN
hZmS7QxD7ZsL8k/F9mndCpR6T5QoNp5I1zvJk1AGW/OiGD7zvj69ZXvb8mEN4eO3
YxSQEJE70sXZf0u0EsO+zmvVmBQOJ1bjTQJwR2vez3Mo4K0aDsTxdoOuWChAWf1l
4DMHWr2P14YnpFs0HlgsXgmXg1Qn7Hjot2k8fVQ6f0khMJU4r1soUmdjelcDK8Vh
SeOSh8d5fHesuuu40MKVf4xVsb2SXdsp5vnGVLpm+pp4axhUlOIXw1GeSmLMCr+R
yKqKEl+NNLLQxVdrUYIBhtF8hcHQWQpt6dAmMI1x4bJmJUzbqn/HAGBQKkGgEZam
13H7+YswpHGfnCu2kLU5Gq8o+60WU3db4aC7v6Ge9uUtL0BlUSUfDs/zhMbyUwB1
9vqWbA5qZo5QgiVqS6OpdTr1s3GEC+LUJchLXyxMhi6Yg8V577czs1Im0TI3557j
GDpgDWGhdZAq1fhXeAWxe7V9eIaiwbEmnF4Hhj6u4ETJCViIbGgXuDho423A0CaA
oeNA+lRnmBSfEFS7cdFlfLVJh0WouEuAYUCqV9k/cvE=
`protect END_PROTECTED
