`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SdtmRsS7oYOrIpdSuV9oqNxfY7aP79rcCrbWvJgeZLdkn3HoQkqAV30MWPw0laAo
7J3KQASPNQnOzL755x1rkMWdZf0g5gk4bYNVSg71EgfxpgGAZAuM/EkJkBq3jLRB
i6i+XR5TUQpespbbISwmUdjmKsdtAjeYQr8jDo8NF5vjWq2TTdXW0cZ3WGUqtkqK
O28s8HZ1hA2naydD4PKiIKUIpR7TbLPGltUk0iogRZPPzYS1fFBMxMKIUNlSmx4F
sBECWXcjvmQ+N9QjCSQo+Lr1Z0K9KiNn1ydIZW2fBgyFt5kxU4zNyuwLsHnIM8lp
Lb0F+VhWytrkTk0E0sg/qwD5spGkpMKwTJUq7ia6oGyAn0rxAbyE57XnidxUQ3DU
NdmqYKNwY/TsmQiJPR9fi34/mk8yCPJxXRX2MbCUl9lLFB/FieIqqVfBFEhFc3cU
g2RSYYihTHsgaViPu3M24etbU9u0UCk364a48w+kWcmz463PbvmVIBieeJa7fqT8
sE8VzYy8pG74WOqLmNKF7TuAe5BqQGHsNJVNOQfCUmVgBxTftFolVDPWq/KmirYN
BAYONwcE6d7mMVh7PwdMje2TTPR2EAxWwoXkFyg2q8wx4YWdhdgcgHaQLJH8PTal
ipot2VWj6K1QJPsqQ/c6xlxr99Q73Ymzg6faMAyMa3c=
`protect END_PROTECTED
