`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3ApOlSXCeX+TqP7rerWCkrq6UssfY2dBIO2456CLGNum02Bvi4EC+5wYHS2W1YX
e9rcSQqxU3EW3mpqwF5cvu5ltIDJbYnr6108Gl7uvn26aPVJE1f4URjp4Hnu0tXr
z6jSZD7K0B52u7WJbJ3qZjIwaUA8z3buSo4buC20rdDNIX+SKkiylaiiZ2xLMLr8
9F2jtSfROLJS8jZw2+JWqc7oICbFShIUFSmew8Z1UEmWIHCxQGl4j6c9T3It3aGi
k5nDOSCfhl/gNVE4z+Vzk6lFkTyjndp42RInT3b5PepYQB3UwydZ2p/oyul+GAXo
32DvSVpSRCR/sdeF6llgnY5XF74JL8qimtO6hh2+Mil+vMUy/w7pU0xyVpktTTPH
sh+geinkPZqQ4h3SUbcZABIy8LXOa7fnaCSB67eZBixu2L73Gg9XLCIDKjG4jt/y
TOzxdi5S0/JadS0X/ZOIVGmh4ya1VdnzVn0ivIXq/QGZQxQyUvY25HLyjfgOz9Ih
NlNlk3M6UR8b6CqFkXCJodq8hOXdUjng+KrbPx3+TCSPQfd/Tw8zWXSR2GH9Eas0
lG/nP/ofzLvod0YsukOvuRZImIzrqsqRhubmJr/7rq1nLM/C8cQ1rIASAcFN/N6F
V0JFA0A7IAooyxXWriGUhI9xzJDUDua46nN+lBokrLQqJzgcqnXCC+u4Fyc2WT6p
E9US0wmM0RVD/DNNGzLnlBpA7MnBpp440HBLlZaWueug9IU9x8zC/+m/5at8TC9D
n4eFRnBWfQOCvxgxzQXVEwYlkgQDGW4SPUCrhnKB7arYU1+U8ipRJB7FvWVv+gIq
Re/5762Efqr/v9h+xHtpAkDo8OWLhFAITFNAfH/HnUtZWTFEfEeCLyIQBOBvkV30
rkz+1NnWIJL2OYf4nh42YJks/vS7gzz0H3LDXkDKAaEPpps24EG9TOZZ8nI5Qucv
qQY62MhgWeCEk4CwjLGGaudHqtziuN/RtjCJgp79MTilUNsrKnCZvg21cEEMZFzu
TAVTDpuitUHcWoEHNqAf2cYIzLEzRxAkGM11T2M/yR7R/EykV2jL9Y9kMaC1ED7v
ahw9Rcl7Jw8dootwx4APB69bq0uTaPKkgWFXZDD/0RoC8fzCNL2CLe/AXieloRbT
69qDU2M859iTbrrlZRQzHFWhwx+vKMSTJ1+u1uMilMRgkYr4r9tVeAZORmAdZZHa
MxjIIkCCIHptfaxABh8Uwt7fat7NVh2JWD4s5fBOq8h9iAK+c33UdSVYdGuRvDPJ
2YJaXuCKgvsVIKKyrPhu3gRuRQq1b6UWDDNqIL6yXW3lrYk69mdFtbWe2LHVoKoO
Iy/PEAuzMvG50iiaK1cU4WjSps7xDDTa6vV9RT2RcRhydzgRkTFRz5PZeFslifqC
lwVF2LW24h4DIefRmga2U0+DAtUbJRMmO50283SS1wSz1w/ouMDQ1yzCAYyG3fuO
z2DebT0vNSmb3LBJgdsIo5w5wrNFnf7DqXjsAnISbMqJgqGaCzDflE/gDgAsuinq
ihEcx/V4oRbCyUYKvDy9c+E0+PA28p5MDrRg54BSZYRB6Q78GpNssFedbAQpjJxa
RmBKWy1b4kaNBfUSUyqGPuIb8x2nGpPLlBnWS5kC6e8JA/VGW1pe2nhzWDMSDgCG
Xu5lzOFle5yeu4r2Nri5pZy7WBY4VmNowL74FR8NDbGC7ljJSk4VV1JwX1HcWcs/
58k3SpU3vHb26WNhv/OUqRrOdXA51mv7c1JQKQ+ODvIcfO63z8dPufVAUgRlT3HJ
ks6NBNU+76DWobeyXXNImp4f5k4QELrL9//ZLLwt6JiYok/EWznpCWENQPfpY3lz
/PsGexuO9iCYS+8bqCT1z2tloAqOLF4NKuDp6loejxN2DqhzdBIfOA/TieS4igAn
hfbD1DwNawgm8AUxui5Sms+2k5lxkExX57TmyalS92ghyIOrYEv+ReRlaQNUmQos
1517QBC4K4MMGYOet24yOt4BSUfbt3Zou4asQ0rCdHPMD1GSmZpGlHtjDZdyWkgj
osZVuY2G3Ybd97RbcJzZF5arY9YELjElK5zVGm7EtNClACxGspRYaNguwFDB+ysB
d10jk51XPmb7Z5f8Xj0ebAwAxbg4/nytstGBikU92kqlVSezzJKnHDM2rZ724EdP
ol/k/s178xqHtwX9iVLzta3OdJ7UY9zX0EGGc+9VzNDNmawvMH+erVoJ0mYn47pb
rx/XrtwwA1mBbD36QXBO759UfitTxH8ZO3Srm1oPmsnP6ptQx39k8IGLTMTwAEek
foKNW7mAOVPqhvxWIXSdNboDHn2xQcBlrvMZyoj6JE5z8CYkiZTX1LHzNAUQDHRW
rGTblCJ1eUvLJBurtedC+ddZY1yW/hm+hGGycz3/eflo6wDz0agofKQxQ+w1jd5s
L2B4OdABa6DpDGFk8OwB4DJgqme/1s4R5xroltVarIx1za3SpZzblo6NrWF74ck8
GJjaMc0PMYxn6IILjLNwbKNB3aJdB1dTob/NnB9ePMfThurTUKYUHiXeWevGOrOw
OduGjdMQbzx61pwcL3ju6IxTSj+hUVUsoqXdEkqmxlSifFp4JpJOvrCEZKCxvf+f
f0KLsSEP2NEAZ/fFJal6++WhRrtU6lMnsYxqFX9BcX7g5wddV4w+gz8ZkiD0VLlF
kWVdn6AsIaNZH1fDNjqGMvAWV4Unxz9xHlfxksCBvBJnmytty3rOWijrHzWzJgjg
jsPBJ36BulWUKRioY6akKfOYCbam+k7MDcc3EIJTICpwG5hWDkybpMW3mWUSeR2J
u/D/O8acSYKF+ocPOvFCtjWMEu1DTDfgZ0uwro3fkvDjZ23xfQhY7LDAAfGppm+D
gHqFpvagti5quh85PoBJh2gcPU/uDhXX8Rmip10J6R4DDbUxEn4ChK9xWzDDZb6q
mPwrA1EjrqOE2F/2vlZkh9EF84L9XF8kJL5haUZUUkDvKO8nQVC3BAOT87UpS1G/
UxeYilHs7Z+pnNQhXpsdVPWaqnuJuD8HmZa+HBtIBOPLARmAoWtK/swOMj417xmx
w1YtP/KlyBeWWt0C5S9rzhmR8lrBE21L82JoW2DeD1Z9jSqcPv16idMS67x+0P7+
k25v+amlGJPmF/opqY2vzkE+eyTnEAV/Hxdliaou/mT3BtrelFZctETykD6xkdG7
A4JpD2TZTiKqgYfDhxOYbRQPJtJlLe7bDYI5niw/bVVktnUWVsjg1J0dE/U+R8xg
uTN7/IF4AgD4AypI83SzmZRW1ju6WwgmUaCrn/bXGDtd0nx+OMPzwj9bWUBnrtzh
4JllxCDTltrQ/cU8HBKnt90JPyJwO/k6LwNBAFhRec5pii3dll4UQuuKEXE9uSuZ
v+VoaSYZqf9MqjlBEiRnOhHMVdRUO8lftRvR0YTO5VIhSiHLiKmP24YYiehJKIYM
esUIAHFiiHjG0xnE/+KJklC6P5DkqH1Nh2m3udUPa+HSJuGWMxXFQ0ronyJC1lCU
Oa3Iq91HhWoPAooQhs+4hrgSFUbd+UMMse8jBeTSE7ediMd/nCNFuZAMHrcuCDYl
MGu3E15/7s69gn8lbcLXnfXa81LKmphWvPNCV+wdRbDrYXty5g9KNlFa8/y1udyQ
GbvenaZJpeodXhnCPMDA61G3Nfc0EySGgjLcg1eCbvpo9HWW7JQjA8ZQt4w8pmZo
JvJSuf8d2MpHf3eUFBUoW6R78qMjn2dD0AFsar0x8rCes3y7FbqsqFcpH+5+OAi8
xFJhP6vhOzqzhkZ9FfI8O+yrHxokb46uI2Ijsc4Smaspii/E1u2kWoqbbBnjvM9z
kWw1He+029A7MatJztM4xKvTj4wxyh6i0vayHgSAlUFV7dOA1qdiJbIq+TD56Gbu
XbYL/bSco8z+8xsmDgkjMbIA3LdDDIbyeZH4GJAY3iIpIql2xo/XmFKmV91mqk1c
5iKLAe3+ARVpcl1p2rXdDmU+LPfMN+eZ3USo5evtwQpQ4/O3ZslAC61kcFv/hCsY
aozF/0zcFwnEKfHZZQTayzi04ZVevQ0SK12+kbQKLYHsThQ319kNyPRaH0x3eLaJ
MNRvufxa71JsWyjNjlezBLm2GT0se6/iiCOxsWBn4xZVEcsBeR6dt7bK4/0sxEqI
iA5gA+Fyu5gsg6M3uGd7TwXkEukJbBmy1AmIJZgrlSG90Fv6OwAKYqGp1N3E8wxS
xtVrOWf17upoTwakT47F8gvtbFtK/xn7pfHoA7/zovwpKXy5A+vtEz3zzyncG/7y
sxgqSQvzUYDpPTwGGmyBsou6hNADYQP/VuwD1n9kh5a6x+hDagl9qRWl0GbD8OHN
yRSEANS6T7K0SvVRgJsPPQUChWQ1A7sWDcOseVVB75CedBSr+vZqZQunf10qLPnd
Ms8PXqymk3YjcryQxBCQyxBRHG2Wl4Pd1PAIruO5b7iWIndIry3Mw72dlyd72+k3
d7DE5VRfR9+EosykBWngcfj8+eBaxB9LUwfRlSWork6ORIek7yIkchDqd+wUR2GX
EI+oYasXobJnxgB/6WFWJgV7v8De7Yx6reqv2GR4wo+a44LaIkeL5wQLMJtH/L+r
sARnugwVqvA/FM/5hiDUTX8v2hs2AqHjh54aL7dzgedUpvmOID1sA67H/xia+vDK
tPOutCQG0jLc6v4QcS+oHRyv9NHeL/37l9AiEMOFVEbs0TgE/0kk3iiF6ttOH2x3
xll5BY8VLX52RIuBbEMqjKHKIYMb0fYcyMKXpa78dfAlNJWBhu4hZoF+hvY5F3b0
WgR+5ixagrr09TCz2hMNu+eBnrTD5b+BhqDuu3fo1gl0xzTVYiYpN+5/sum53rcQ
4Wbx5h6vQ/mZN8vhoF7JBj3N6jUzoTbCOzojmUZFPM+wiZXTYDTiXZsnJcJQwRPA
N9RVPpUiD+8olpECuoABEOqbjqE7xUtvb56jtheZ2S7h1bbuJhVJN34ODU4DKzgd
+1JYWhVTBJT9W9pz8j57ZT+izpEtTXmlBiYQtRrUL3DpcXjjXms2y2Zy8uzBzCti
993UW7dYy1VZ7XiVmWe5AEINu5zApP649Dehixq0DZdOWk+7Kk4yCkvAd60yvgzH
a6EjAmLMNO1nqtnFd81aq1ACevrXOOwUtpnIL2YWjSRnqlWefQ2R7YsNEiYJ+gHa
vWVcVYjECfwDYmlBo7CdU9AhngpySlAirltldML/WkBbvbIg+YEQMEbv/dsdFTcM
pGfnzz/VmPEPmpX9OOpw75eLbVVDVF+5ovVGdjppYnrUIpNc6rdK9FoOe0bvYYbE
tjfJMWdueBGJw68TE3gIR6NRO2B4a6cO+aAcGV836iKhIf68ROTQ9y/tzy8knuQr
9GnVkVIGLC5cpHJm26kziOxqzT8OGBXj4hESwcOVR4ROl8Y/EZgssTWqhQ9kcz/i
PyaAemnwPkaX9mMNTTel+dgVk5xZbOphjKbap18CCDmsGkIU2c+l73PD39eGtuBe
zBEaGr+5ezBgiIeQkoLOOQbZi5aT82KOSkWErnynN6Jpcdh9guF6/use0qKpuxxi
23b/a/zIqSHGMmlP3Oaq5gXltEJPS64HjxxFs18r92ZQIF3rXTWgcRl0GusX73g4
Eqt9vMyWag7TjZDZVsyHHpIavop1RDQ/zJzSTHkyMDcGwVgROXs2MG++JOzMzstc
HLHDJ/sut258yGOwFMKdaDG681AeBelM/FPDPd8AaLKE0GuJ6gKT6L/ws/f7yJpA
sdx3XKWGPbTyiimZ3jlkpVd/79vvtPUaHvyhznGG0ikUeJDbyoYEcwe79p1ak3FR
6LHnLis37cQkExeKTdhSx4sW3TXP9f25B7dfmkWEnqiE7DpdCf6axrfK7o3R1iAS
ESAOC1hyZAGbkjU8xkPG0a52GSRCZfY+xyUsPGhqomA6CSNdXMk0wghSXHZbExCS
QIofoufO9P2JloKZSqNrarQ5OQeV9/kOUBORoHmJZZHek9TkYvbu4EfdXrYLjuiQ
2rP28PKU3jQl3kJwJDeYl1UG0LanpqRp6ZMGjKLvSabUB66iffc0CcRxzlgKS3pa
MuEyBHdzrBV8Q0CrOJvoZwj2A4IUC95TPgJfifXVbz3PbTcHgsI1sh8Yci6b0Xlt
TmBJsCqZu9cguNDka4YTSgqLxLGfOsEGoiR168NNBNDLPKY6dK4QylgpzLU/9Gt+
moW+d8kOjuQ/gRf7M3pBhTEoOU09ghAxlkCTCgBT2J281Bmsit8dcRJunK0I7BlZ
XbChDhXTa5zwnkFQpSGQVvlg4jBMBIbxAFy4PjH/Gl/CsnT14l8CFFEGfoWom1eQ
7cM/lvR0qkpG25I6RIMmVz5CRObL+eoNNtZWEQpqPdqjop2LPxJoZ04dRZquHn4G
jUd7yiKmOHkHxkjZUWFMG4mlGsL4JUw1jHj2QdGGBRQ3DIFtWikot3/tHdLxqVJ2
hEkSwapms5RkfSpkPL/sUzsGsIdynDZt+0onwoBnakdX/A2uWhAQ46yjZenpfcU/
WHnLebx2nMrIwA01B1ocgoJZJR1o5J0cAnyjOqRv4J6ZqS469ft6fAV/JzZQu/VN
+WQcn3rISKdKspkifqwcZbivvTORWjZYg9k4FsRwkknKTNPYIyFPYh4QRmSE+0bg
gHfH1bsBtu0pv/cLbhZBduO2fztciAfbo2H/9M0BgKzicn3mlUkT+l9mws6DReSc
F8qOKk6n/LwyM6FpSoNuqZ4eRA0IZmqk5C0W059SHZ0Nn/YZd7mw8xAuGL9+0U/6
C6by9H815E4eDtrmQMSDwYsvpIEIgIKlDrxuQIeArx+heW3CdKKXxyeJa7cJEN8I
hS89n4g/s9lWBBTZrn16y9TdZWsfirOGcv3/eQdDsLsyjNXTa1/ztnix2FU+1rBi
VGdc9hiZvhCBcriEP/AFtYN4SsU4hXqH9Im6ygPMbVQ7YWZ2tMw67lDSIrkD5nR7
CZVUUIwlDmiUC7dNLmDpP1OtZIcXO34vj/xNl46BpOfv+ZuL4j28bm9mRu/t3DYV
N4ZHRtQei/HU0YFlcw23AaNt0uUMh96mFAim2tK4vQvJINohq3nwm+hnYKWuVdAk
XjdZPFOR4qLnnfkBXHK/pUsuzI6pdGcgORRI0y0m96VPOLyrU+xLImE6ht6uadjU
+ZqVHy23IFDV6jKtkmiY2iksv5gmhANfTfLgz/TewI0N3wQbWSr0cmalq6sHJCVo
kqZlFRlOrUwGSOp7w8HicvnIWqq26Scf2qu8ADtJpaNBnd6uCx/hONbP9iWFqv48
IyOewIAeMeBXA024ERZVxX4guCHHT6jK42jTFqjl0fVEicvop/hsPDNMgBfJZ/nh
2P4rJNuSfNWILACJapifwyLx9ur7wg1thA4r844oEGbdsntB4f8wikeM7NXXjCN5
6vaYcAk+RU1dT2jdUFXVOsJGfze4lLKSg9LaWWpHdNLGQtuhbeZDn4HRgkZIYt5x
JjPUVqFWQPwtgXw4P3IsQv6QlpZmAxA44r5u5AelAODgDMAz5YDNJpMqf2VO7Ec2
s7CFppFmtSvvV01a331oD5ZnXXtG9oty9zrH1zOEx+RXwjkN9NmXrTwaO2Jdq5Gk
saG22lzkEpLKwHcxf7z3vcjbVgyzZpLHT1CsaawKL7pl2GJNNdkSf2YNTDl3sfdM
OdL5w0GZ4JWyI3Gezqzy7H9PSizn8+uhKnWB9oCphUEbXvUycDrpZk6p0oSZpBzx
xBCrezOa2+/BEKlwVwGemvnk++Y8u5/Usqzc4VzAwGDqJ/xqrh0BP83CZEj98Rg2
28RNXinYo0VBfcuUxAcR+COqNPacTFxsvbq2BqZPdC7wzW55Om6k+HD/j6srbCbj
juDVzT9PdMfai/vHxocG0tBaPaIuIE5jMN7KveAVngaSxp8qLmWCZPVNFJy6HEvG
Xq6gJtk2yXGoEpMU878OYl9VbLtdSSpCSgADvy6b+Lxq5+E0TG6YsPBsDhRSYQsr
CYeM+cm/f80wNtDst5v+gD+QkKWwFjRcp8kMSuLDdcGcAqUqRaqCZm4Mzzm1BCTA
yBqO0mrhJtkC91VqvYnpcqrO6tGz+whay+lgt+kqULMAZYBsXDd65ihtI+gqbUvh
WE7ftqYsLTxuX1ixoYv+sxyljne6UXiLyE3YPHiweEKJRayZpXbg7rAm3GY2ivR6
hdVLbr7/XxspTyco+WEBdbV0dsMWLN3kSoIiJqq4H18I9ajbKj96CpQy+8yVLhQx
ZDKikvvwOdQt76JeBhaQzpxC8nKstGIbClxcp4fquzJCUTdAUfyk1mLaUptU5aFg
yxv7pJpgHQdw28UAWS3gi2DbWUOT3rBMTWrruTPeHoAdLLdWYv8kAeH083akX0DH
k9Qm2ZLFnsz8acMYTMqKaPnRzkzNMw9ZeVizihIX7NubXtzTABgsTMc+1SiAV53t
D5RsT3TlCOCGB3DIQ/e8GZwdE/72EEo5eU+AJQbxTlnRp8Sq3fu5rwkfMfmpXtiB
ni2UXAD1h8tNU9TFBPYdLDJjaxBQ7oDYLhRMxfSpmK/GUBtNwDXwpERnFp90lqb2
zLwAD0M3dnG3RHcvtx4tAlghWhGgibtJ5V7P474U22hjEZUdMmgnLyhjeQwtntnP
MlXDrMc5oxlLEfsklOuI4Q8U9fj6TeVgIIg7hIWqbpyQGD6u6LER9VBZbFKaq4K7
+Q0JKY2hFQUp0Py3tBEhG5KsnBU1u+K1hgjRrkdZVx6DitDL1pPCzaMp8luJnwcr
Ewj7djG3s0t6r42AvW1ZvKq6R/dxJrp7NRDWcBWQrfYMhg8zp8Gm2mgwkJuR0tZW
MQqHdUWt7+PrYUiY8+lZj1bg1TXtqPIeOBeBtkdUHCSMz4vojtEkyAypeGRj9V7n
auMm57GuiJrwvJHNUQYPJRbHGL7I0uYmmGXPmyga3JMfDE9Iygmu9bp4XyO4Pu9Z
Lhx5ay7thxdV/NZ0VUJ1KodCui2jWX6kwYuHzNYG81/WTt3iBAfU9GIKVE0m+M4B
JMYMffygA6InTsMz8BWsezHdbUBu3MTZQVNxWJ5VESvki0UWZ6W4+BJR80WC4pTg
930eIRA+giSndslyHrLPpxfUg7gvNwz3mgxateAIlX8UqTC6tho2NEgAJPwv1z2r
EwJLPeAqnxx+KnkH3MAri6MNYh3C5ehi6Biy5foG29SSiE9KRoIHM6HBEw24q+f0
AAA7s/RVXyE2BCyANMHA8octB3tsbPAjS47gzcNswqjB0chKqfIETo8kBPE7Nuqt
96oW5RuMa+LB6areyUv/OnNe1SnMIV3Bn3gyTUwSFF7U5JAyqfhc8sUokBB89sxd
h34zE9PguwTUT6DlKS39X2J3fU0Ai48JLUD0L0Qi0gPWJyMjdaencWeZno+J5oqU
TRz4Lg04gQXhe6SAVf+BnAGe4LGnjrtXps5bWmKoO1Ksggo4UjXq2IfHKhPLaTTD
NRVDTWRn5F6Q6gBWztxW/hBgyV1UoS+5j0iL7mo7wlVJEc+isIUnEUhAxBPgbir4
vcTseZMOFhDeHweTzuhyyBoptR93etR0RNxv6GcFoooYjlgW2vmH08ECwTd+o8Y2
NxvecTBC3L0EH+7z1yBZ8ZzixRu9TBUXJJwWxmCRuhGQ8F7Te7cqglHOh3L/O9vE
C4zvlw/7dJOwhOXEg97LVBsGJS9Nb9FkMJfzymFbZfVMxiH9URLuqDB6tHA/Vwzx
9Tp9Asv2kkwKeazi7QGUmZqyaCmKvsdXtivWFS42CKOTtIMhOfZ+Yf8PNKMY6Ikb
tQKHz1JokLeklT6aCBobEeoUrp1OW2FvPx1fFhTJn+wAY3LaCvJjLBxSdTOOf7g/
fM2vbPRLintc2vJe2DMzkHZbYTNkBe5hNNJswx1mqwhoRaSmVs1cRUM901YElUPu
BkiKZE92WP6IjT6UgwNCKNEqpZQEg54bOrQfoUJv4ElarBk3PC3CKFIEKZy02iID
0o2m1F8wprt3VJvO68JJ+9Wd9E7n+TqYLtmcPWc+3vajpf2mLg96Ayk/gmdUH1Co
7wLCJUFU2vS+/+d1Drz1fiImCNz9WOLnHCJxltyon6YQtX5OIJS2dV4+/Fz8MRtc
n33LIATmDD0LQTGPKOcg1nOoDY52z/u2SwHEGQrFrkLNGgsrclnjwPAO3jXHsIsN
TfUIxHEfydhXtWUKaKZVFJNvdRmnTrPxqEQXP6k4p76MwNUiRkwvh7tZ0cWPfKlv
ljzWUTlyG9AyvoKFO1CvM8pLMU14yaJdZu97Y1TNmHDWrq3qcyL3UJpTN9AFbEhq
XXJQ68TA/qAOQLn0svpnYMouUmqWOOefoZ8IsOyZnyMpySgCBNTl4khjYJJxt1h4
J31rJX7k+b24JsQAi9XrS4rnCsulCb6FM/v/R8cZULuF0j6svIhHUxZor5GDtOPI
EPsSILkojyMXiuvOq+pE7jLc6zpDsh+53mT80zYQLfLJJOQtXvLhvmkzxM0DEPMi
WoWqI2YKbAj5QmuYIGHOYg8nwVGlWoSF27j35n9UAf0u4fEbOjnYLlgNP07t7kTB
MOB2bInx/oaA7Pg4zWusXEK5dWTBz7DMWNisutJC0EIBI9VtBtcuPKlxPtDY3AUD
fmBAj55B+nWEHnbsxdgppM+9yWGsFbz+34gztpKdyYIcoAWFA/mkPp2IY29AgmMx
RREMS24X/+A4Ku23ilp83yblp5pFmSnUkBwM4+mw6/68W5x8AOVA1YRgqcO3Bv+f
sZ1YDoD8LCTpsq3ASpFvmzVIzGAGNtgstvCmm/QBB1jrMr8053Y8mqWF50ZAsyZM
Z3WamZO1eFmiybjDI39wsPmqMyRYIDuUbUmmjDR+dl6k0mx5jzlO1FHCWnXwXew5
2RheZokbl1/32+exZ0mRzt7lZhocibrC38RSfElvQ0r3dwUBCx95bAP0/1p/ofwj
FMO/7pP250F2dTbprzyWi/QZj5XBRthYp/ahaL0JQraDZs6dtPwVDR03vxwNA2IL
2HcS+zTkRYBw5Yne0pzsBL7BlugByNGI4INfMitvO65q9tkx2Xw7PzNPJiLB+mqw
6bXfbNOmGNkyyKQRCRXs4scrkG/G1fRDZZttrPp1MogUIjs23exmZmTKNi+lY9I3
ujgnCiCRiQ7KI9RbwCOZczIeCfY0ucCw6WcuzsSv2DRAGaWMFugzZcYIvLFiAlyR
ZUPlZ8gIHECUWCEZJnXEehFeoG/FpKIjWQP3JMmJUKC/nZbbJf15zBunD/7yLChU
J4S2lllrqqBjaPHFTkEiCsy9VC2iCbGKs7yoW5brmxe1Go3T9ZeSaKT/XINo49zt
+ho/OCEGUBsvqceaFRW9tfFv8Rmjq38nWdOb0BnUvOYCQOmsEZJIcgZuQn7KjZTj
gt3ZB34aWSCtgI0K8cfFlKbP4RwW00dBQ5oR1ZVpyUr1wmRCOABQn38NQoUKJufN
kLxQaPhQJ3lkS5Nz3IuhI/yh4QcmzbkRxVErwbkiM2wlVzDB9i8EK54opmSCdtWl
Zs/cds23fYlreo2L7l9SlBJfWU4U3LcU0v+hnhB+oZ8kArSYxE73tGQQk5hE5KJu
f8nq6KY6xHdvxq+AyWJeuyuh7IDzGqV/COmLrBGs3B5WGsxUHMG69r6yQy1YoX5A
DwwXxFn6FWfhIY1BqNjKPm69nMjDQvZYZX31tniHodQ=
`protect END_PROTECTED
