`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wtc/d8FAvx8fpXNQZieQS64Dv1EPiEzDSQ7GgoWABnwNXjKFkdv1YWQY0FsoMO/0
Tmpd8dXLLKYuZaqholcQG1uhbkw0HM4VP49Jlh5DW3LGvmIwKpRU2SYdv4qR6Zsy
zxGCmRTLdFaPUTnfS0L5b+HLKFvkKgup2Ef0FKRzz0SxmlQiMqir/mbrvFzfRCp8
k/GCctlT9g8T+t4vh8FKttRpa04ZsUzThs5pgp5nh4kyDZNjzMXT17kOTtD7BYBY
YKmhm/4ZsWTONOY++Q9et5SS6S26+kDhrNtrJJGB24uW+3upr85h0FK0CZZlQHaW
SN1sXGZ5XnS2wSEQmbvo+DkdNdOZI+KgA3mJxQoLuxcnWPZgE7MM8+qPV0BYqeQi
cO5VLu0eAjzRkA8JcN/Uo7wZWxw4dCBy9JvVB5jvhw5kJNJs32XpwZl+kPrpuuy8
D2NAzciUkGad9Sau6m2v88J/vnNCvDSOJXUcm9rrKfyEILxZZpdjrt0xzXsEpBaL
FUfDw6v1BagGzio9t1Wl5DzCLhzPyCw75e8QiXPiPYbWYE8fI28j7mFZBzh8w3Zj
TjhBJgb9bfyQ21TPjsObUSMxHq3w9l/Nl52dWX1TAiM8D9xS0XEr1nHMQOYMkfY8
zi7/XXsqq6g6/pblUaMtTtc3kIhuD1YVK4HF3RX0/tRT4cpHZBbapAJf3bg7ldv+
bg+tP0WWj5+3jUeIfOuEDcixt7I8Nc3WNPy22Vdf09RHddsgi+KeG0kTkxPRzbIs
qbuaohzw5NwnZKlcv+F4pvnh+zDNA4LU070kpAe72Va+kAUkgRYU0Gu0uqBHBerH
JiYr5WZ48PoDeyGIaOw4jwRuJXtk4PHAGU8rPjry3WdjmXxXz6clXIbRsx9mSUH4
IEO9ikNsNPCSwsJ+hfmtgDh2uAA2fMknJaatPT3YYkGG4JPqlmv66Ok14W9Jlf2r
VDxTFmS58m3eAASizFQe+zqNeCwZPUitLcUmD42IT/xOqMUF3ymwoqX1S1eKBy+r
fMXkvo+VKpMhaQilAAlKyR4yJBN++iYz9tOfxVjzWLM=
`protect END_PROTECTED
