`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rmB15tP4VuGDkYJhTouswX43JfmkySD342G8+zuXuhswOwBCwO4kXkMtA5F+Eup
I+91zJok6enhc84eXwnO5VgvSGNEDy2qK3FRxsWWMV7BMPMen/aA1uanpxkQaf7z
tVvNJNrnue3iALdjt4fyM2vi7e1aeHvc0qzHQJOAY5E5RI56sKXyFIkkfRiOcMTr
GJJk258T1in90oknKoD6GNg69fHNP+e+x/jQGocaju5U3K7ZDf/BkjGFbS1kypq7
hyA+nx52XMlhk/IdL7XmH3u4fDjK2gHVMh5sdT67gBUbXr9v/LeelFqhQ8EyMNLZ
6TJmFiNp+sBwie0qRXZX81UcewJ/y9ERT8gzcj9oqZLCBeiZ7JKCBnEN/WiUihDe
MfHAW9wAY2+YYWORhGQaLpS5Ik+t8j/R91r9CUFdZnxuuE8gmjx/0Y0mGMYe9/Xc
p+VibM1apBub1OPiShc4oRUaVvTSx3rPlMLwK9XNdoB7elYBS8h/nRPb0QuGB6Dw
/3mEZ3C98ra9AiwIurAVStm/NvUMDvLnUwiyMSjiF6YOg8q+poV4VvEKyVAEYkVO
ZN7sguL3/Ldt/ak6tsMzEUB8no2UbcmtT4/7VgvQRqeQ1wb+gnI2p1eIn0Udkksc
+Cr7oNkebZr1/FRfULCmbjOwPDO8Cy3ifFASsuKeDtPyGyNWyLxo5UYR3T6m4wdN
IAQFF6LfAXWNIaDci0wwio49guTrrlw83mX375wwVDezrwb2J+hJfosm0dlu06Kn
5Va8kToScBIaCgOWsEnZoiLVs3/dYxZWYJHkujkbfrrucNMsvi5TH8f+JWnYJY6B
qHp9f6O0Qfy/xJPfIJLByfMt2CSozC7ob1/zTj6MyOYw6ax/DcN6YV6NFuy/dWe6
b7cBTLY8BScjQ0qk1430zJXUsNXPjV83+BCllBPxgfe3jeQKDd24oIr/HqEtzEm+
ALEfvb9WsjJZNSUIuA9olbRN5uAeBxQQ1ciM7Z9cPeYLgznC/ozCfvaqYUQIPUyj
nblmGOy8wIzL+6wcbVN8xw5UxNZ4MxSjwWuoQljdFdL0ozmvtJo6au0sG4MIBW1+
vwrPG/b21UZIauDJgtcmvg==
`protect END_PROTECTED
