`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJ7ruc3/mfj/PsA7vv9+/Z6yjMbsPAI0Y1LJMZOMj0/9jqKNJtMdH0Qo0HL2yFUv
P8eDCUVoATSrQhERkS30CGBf+DmySiYTYVZZ/ix8KwTTgPeXZSphixe0W7wSSwZt
ADd3ayiybalFLYG6HM0Hn4fVmqDS8HnncCixuj5sN15vT3okEc/qmj5Ean/T1+tv
OC5ruUUWu4PwaXdppJRy6VW8ODe9hHTl1Kp9oTYBAkbCB3o48i+OAYJK7TvLhPg8
IEL5Q9J3oT7Rq2uS04TWrDon3zqjkHPNhJ0ANO3t880SyZ109VXTSVDBd/KuLveS
ypViHRcSMx7m349d2eS/saJ2uQbcZIIhwYWLgHR+uIwGmYTCriPBy2kx4rWSPOsz
KwAXHb3wJxM/35dYSiZJdw==
`protect END_PROTECTED
