`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0SCFO9oUJgREa12VlD74GVyRqAKIEpDaTiEdY3KKEzWPXoTnfUbH9DvRoeIpMIqe
zo5SA7l0USHKba+Po27P7U4psjRv0pp3IzMirZr8eGNlWXg/7lRfooYFkA+LJoYg
+fAsuq3tX5VP2FdSmeu1mRXqN9ibmbRR4MxC+t4TYWoLp+WIwYpRgenUeXoJtOvj
9WLKIB+RqIFM8AJjgmrcwu/+0vpR8WKxZLvguK3p1rApRiuUrS1BgXwGXjGXHp+F
Mm37SCZkR2SvtDMIZsuXNGqG/yzaZ3ppua3Gv0sZ+lOd9Vfx3wm9RyVLkskPOSDk
FU6GptWmv9WXie1os+zdecjnJVf4JAgKRn6lyZZjPIXZITgh+V2gNlYrisdlahiQ
PLPnJjto4U73Xtzg9BH3d/mKbbrb2mzXaWz2/ySb0BYnT0KNVA1IjusbX2jkBUR0
BklbR99nJDlA8N9GeiZQsA==
`protect END_PROTECTED
