`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nm7ediCwt8hF4r6/h+2egQF3oNgEXyjKnES8UearAMXUGdt1nwrkj2ZLuv5Cfw0i
UaAKUMP2E6bsJRf2DWXHp+N6fGJl2Cs9DF0p3MULFMwE6rHkm6A2kaORb7+ShY/V
ci/Jh6ZaHDl+6Zq29YsX6fJOJNGwnE/fz4hp/EUi5h1piVbVRMgVtjURf6VdiR8M
MASgMJxT6U6WDKp5QNIaZkdalfGQcxvd+/aFoA68koiARmOwK5KVr64BZ0zJFIeR
JlCfI5bhDMGOZwaYvYZQ3nmYsX8YYt5kaC/jTLIrzZfv84WNZKa4XeSZjmLb8poo
THmNHdBdnNNBQAhSEE0lYw==
`protect END_PROTECTED
