`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RC0YSKL2bDruAJ64lamBjbP3/s4Bcv5fBrHGQ0FipTJ7kS8ewfjymIazHaj0AoJs
qota56YowIhNiG3CwRYv8klIDP+rroWr9CNbARbzd2X/gWLeMyCLJpwsYEGwM/nt
RrjJI02RUTIiIkploNnd+b+jnJ0z1mPXCyWRcDxRnYlDgchDRsLETbMA0hcsshT9
Ppsooo2XjQxcEyzZnWWxojP+xB9McnKST2qDcAgY6AnOf3Njn9g5k6OikbdUu2hP
8/eLiBhuXvRgzIVMDKKMsdMsbpbkuMMdst/e380QBL7hUX4fJY7aip8t79IgP9v3
weypkh7+jsqdQdRVtUJOO/EwGZDfcdMwZ0wulqgz4jy+Z0uGMhw4XPHzZ5qo+OLF
ISMgMZd3CRQXLn+bk4m9i/JN2ufmbXC9gODPpda6TNVKqmheTRyYtlwsbxU1Z6nH
RSWX6mUwtBApUrMHTEpG0tWP1/EWWtYxZEngB7Pb+E8domClfYNwz1mGRYyrNTEy
51Fe2oIyFBHFqUf+0fmFxLCP6BjxtzmwgHyheOCftJlyEbm4WPhyckIELulNLMD0
ewlj4xddc6IKAuVsuTiB5w==
`protect END_PROTECTED
