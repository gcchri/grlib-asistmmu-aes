`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5hirg4F3Vp/qyFkGvKJzDnwWSanZDcAGHLaRzWXMgc+hrlxoBHLATrJlEPcB60xG
HD+sfsy7u5Bx1EIcIG1vBHa+FJDQ2bzBHx+DeLAPvXhABJXkz9my8e5kJ0dqYVwb
rAUhoyvTuiRD2k65hsbkXmcyAmM3jo5PHfDPIF/e8DteROjiE+ClDemofNsMAoLz
vrHyWhCNtKrxW+yszTNu0/57T6b2jVUy1NVc5tVbukncv80C4EmzbC30kVwLGV15
0OQupdAZoEZ+fFxAEHxTkJEOO6jDoULC/3LduxJhm/Lp9dM54JoMeUdYyYJdESZJ
QkdiwNeCgKbbYYIeoHarEhiNZp9M+XQh5MCbT31a/2a2EYJNjewqyWzKRjrijO6g
ZTHm+z1QRU/PSFQ/oHnuxGYQk9E/exbvxjIceUPWfkM4xiIB6KOBST7+kJqQgATZ
pUqOp9jURqP4eOzUqn1/9kDKyP9flrEUumba5E97PEaKOboLBqbirJcU4R+JfyOx
2hdL6eviDfZlHD2MVL89qRczeEuoxA86hpZNO5shv9CPRs2KozbEl4h8jaQPhhuE
FQqD0v+7g5PdHk+83J5/WBMqyPjKGuRAyQnLdSEJqo85PN57EbhvcCcEzZnEmyTa
qjnw2h5uKNK+LZDJDSMZYJRRh2j90XJOkQeSF8obRI4YFqLXcmXzc8nHDMjhwkVs
kAbDlo3TjsMXmXhnVTEqlV8LnfEfPsPPbPkuC6VmmqiE4LReOYNntU4eqwlimCKD
aygUVpxyOjQIrDUq73mUnwS0rcFkzyQQamnEXOich5xgoRyRMXbu5jOUwIjdYt30
v+evItCBQZ+l/i6Zwuy2mWAtTcHroG1y3EKgZwqG68nsNelLUC1aAreIVLUEZrpJ
wbrOUoOTG7lROhYOi4dqPFgK5WEYr+XlgipKirSc3M7BH09zwIMxARyoKIZgsdSs
wBLHdP8P7XQ7amK6H+XuxFpvItJjgNU2Scm0RC593EX3F9wAXrSG8/ssR9gD9/uE
/cDKvC8N8n55C4CWG8t7ecJnC9ek5dcPDuGBvBqE+mAk90x8nHABmwUUrlju8bCe
cacGd/xqNGe1q0slFxqqaRu3IlyTpemdEDJxt3F8As6YdX0HPfHpGckhzYEuppNZ
okZQ5tyRaoENvuYgLoC5965XeM2AgfuYx1iifSwNekUwOmdURCslz2IuSKl6TLrI
`protect END_PROTECTED
