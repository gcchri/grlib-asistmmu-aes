`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNd6wQc5ohgpiktD6WPN8wkf6T6bQrRlZYQPRtMD6h0bRRZseCa9CXpnHGZqDGA1
hK4aWRyoXkG5Sa+g8BcRe2XJvQsQQCaJJQsu2lLsfSyXZzE1uDIiXzJRrDMZlbXm
Iqkp18FrWItUedXrMbpmF2zBJrK+Z1xZL/F/BUuBet5yZIuxG98gluE7D+PikIH4
Dw3O9jgvdfs8rzNsFdogUDvY+OUR5vi27uNL0zBWR5SHzxTNR0oaf3GgoLGXq582
Q5mi9PCwk9HAeP8LSSkJbFynZx8VbzdoN5u2dEd4YtV8EO0miOCFrI8apWD5FeXJ
DcOGWtoErz86QEe8PxX+EvwGfRHS4d431JipFxr8s/FCyWLL+91rQXnGsWPmw5+s
GeaILJI64B86KAQycLJOhw==
`protect END_PROTECTED
