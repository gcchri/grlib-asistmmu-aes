`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QNg+Pa3k+kjgGW2UOjkBDvCWZ3ZUII1NYQFq70yB0aCoD4RTdf8/eNmAb2d+9EgE
i9KKJ9GL2L2o4jV3mlIBrPrGGzz7OZFp6dodhYWayBO5bsWqLnjsDwXAu76onVse
nBNX1YfzHnTIn+64sAzcRjbYhzh7hr7v5NpBMv+lB8XBe9j5vSj7nED17Gg/HgJb
WizrnEr77kdYwh+woyEn5VpIHKzWqRp3tIK+FYMAqqppzbPkUlKr52smfU5RtOCb
EdyciDgsVzjH5RXhWEEWtwemqKBNsoVE6DOHopb7Y7K61q7Dysx9qqQFwgA1TabV
wVBheNjJ+I0puu6HGNyEfggbyDjjSn8ptI4vkLJg3pR9bns1T3iHwo+zb8H8C1vd
qRT2cdREBWc/YsQ6MtNTzHJ90GSDdhaoYtWrzhBSssIO+lcGfyxPJpuBOBSl1LQS
goY073Ofl58hAe4FvHcs77l+DiI5BiePtHKpKTav5WtvxP6aFMysN8vFLNN07Dqk
rWMoQ3YiXGJLJ1iTmrcZ9TZf0S9JV48B41f9P5/It2vKiWABbsSiwDgDnVQv1ybG
RlEZUxIrS1BV97DO1Uxw1XwulMKF4ik5YNOPjLGEu+YvmOJNl3Qb9+ZlOA2ZMZWq
ldJ85Criq+7Le/lOBMCCCg==
`protect END_PROTECTED
