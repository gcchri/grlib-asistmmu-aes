`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mjGlegN8qzrmPKpJpq1nZkRzQYYxubGSA5nIrcJkv4K+xO16utcsbzdtgZU33vm6
z42C8NrTfdpg2O9V1Ogn1frlnbG9Uy1FKoQA55eOJ6/KJfgSgyussQXloJJTlA/v
4XTRczl1o4Kl/+GPrbQwkJcH8YOGrLckyTsnWt+fqPRbNYOqfSB1+k0Gw/8dIld3
i1wzRiW4QzxLsJMgDetOsIy9I4pMWSpg2Rd0rbXhAk8djJyzX5OK9BmU8HoT1fVJ
Ty3CJFlqgUEiO+ALO+19bdPEg6SCeYEYrY4CdcroD7k=
`protect END_PROTECTED
