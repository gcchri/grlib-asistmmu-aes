`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y2/Bz5SnP8GIZgl4B9btkrcO3HzMnKuUDO7cxjgHbhVtVxwGzuDcwdKZqCmIVXk2
S/WguMBSFXgZWg7n+hkRqAvWppzYdhWyzjNdQ8BRSfyR+UTLeRwOSvFJXH8KdYZU
Ljr2X/by4noUR+JEODNRg1eUFG5+BOKv7ah/aOOePbBT8XfbzK/eOvygNOAIpN3L
sHInOIZT2lJMmaSkfcS3C2R7JaNzZQmTjVk4CPab3HaM3adQizBwoU5/kxP3HKvc
bs1kjflvVTRyFOlHURLd77Q5ahr4gA3uMXxzBz13OuKD2Y6imXWVGoF6qvhscdzf
UVDLiluSmm4cHoO6aAUE5ZMbc2yMquwpd7A9U5Zc61MGS8U/o2X4apewap0GT5+z
GKkIU1dZOaMcXZPqEOkkFZI7lRxZmUaogZdAvvp9rQDoQjA6RNwEr9apTAZ9n/OW
`protect END_PROTECTED
