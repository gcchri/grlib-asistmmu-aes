`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dObqRt3dgJK3SikCT9qo9op1EK+b1Vtc+14ffs85W8z13anLJA/s2HY1PnJpXg7L
BSOVnBa5i/zPjIIYACLLAinLFfwYlpFGRU+jDCF5mvDFihv902l9DeLXSq6cJUEi
DgcdMkXe6XTFkFLk55WaXXwS0o0nuZDaF0hByLZY8V2rs1URUA7TWHEAL+j+Y91h
ozIqj9KqlYnmN65bzOg2M787KEUanmfHC/gwb6ZlWAQGS3UigGTsrg6IFwmmKLOF
Aft/3rO5drqdR/2SfNWS5IX8oroyQGLQGFfDu4yu+NKg4dU3XxZcmkre77J6bXzi
JWb213xXx/iWtg/vZPZnLx/926+9RbmdBZeaM1bPsN6SsXPJ3dPAUhgAPHlChpHC
hplW8pm9c2mp+BR2TlBvp7TIOg4+v//3gnfOwb4dJWCi/GxFe8h9ELAPXRGcrzOd
SP2ceikW6azR1pl0jRZ+i5UtgNRm1YzVEVRjSRdnvLAvw6bBbsg5r/nX+hjLxeTQ
DqcK3/OZax71wnbh5WLWqHMylY00ae+6ME1Qjv2WoiXZAwne1er89NxNEFjoHV4i
87LwJp+rS23Ssz5AT2BPCBO4ORJxerFd48K5lZpQuMc7roHcIdOs3k4zi9UdyKAa
ldd/VBELjfmaa4IbmGnDV+cLmcGM8NQQ8nLkkcgbrUN47eMqcWQcT3Ia2EBYXDtu
LQgQiJnFunPB6mygqROlVQbig4+QOxwpC6WjFcJcPGwDhuqtEWW4ayIP8UVTlg4c
VVm2OTxc3Fk4E0jxwGBtyg==
`protect END_PROTECTED
