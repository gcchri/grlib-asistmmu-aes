`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
owssLGNylFiDqXor761tpBYbsg9+U9hVKY7FR/UGzytKOM5Kwcys5dYDWCbvQ463
cJsT4IWoMqHE00yeD1NE0JyGB59sJr0kMduMvkBvMJYP/Zn3VWHGb2H2RNVqZYyT
LYWx1SDoSC1oyBQ1Rz9mOlpJZsF3cZC1yi2HQxkhPRoDf73Htqq2LT534BkbKkQX
UUKaWQ7PWRf7lditZnU9WoMvGeT01pL0PkCMB3N9JgoBo33gaPcvROXShqldueBz
Z5Cqh57g8ceHOoUBk65vbsW2BZoMId6Wpc3S085YbjtoRgLFQFx+2CLb7QgeTDCI
RppXIRGllKdFe04fOamYC2fAM5ijNFw5e9KRtCuyfEd5caM/scnIeyO2MlEkBFzJ
cIGSGEgtpDWSVZvuMXdanBLIdgiBUj3J9CkScF/wcAY=
`protect END_PROTECTED
