`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gWqQj3ndNhtul7mOQjPgfny3zJRLgURu8PeFTTzcuz14uvcoZv9IflN5M3pJbyP
fm0TJhEZ6myhZuDppau4dfS2gLQVt7P26RlarDwLiq0HAd+gCfeohnZW0YbtSewt
MRiC/ZjCqDqZkbmqZ6Ab3OxJS4SOOucp/VtRpGfn9z5PMjLVLOsUEdBM+SVMKY1V
mcF0G0abDMamWp+UVgELVmWsICD97hJOU1xAWliMv49zuLL2r36BbyHymEnmyOOi
bb3pnsiCBOGcocTbDWaOM5zc1oxfmCOssN1DOAqFjE52AKMUdrYxi4hcB+g6F5IS
WvPrIzcD+jwTQgQE5LESiC4IUCGPKYGkscBT89wKRIFjfrh9hrD3I/Q7lSr4NwkV
ZsT/A1UTL8M7c/0KxQc/czKjtxNOLOMYYe0ioH7wZmJ2GMOzbMX40W+GMyJcscsq
EnNxApkLGxv0meUOtOSb4cUwgWsR+lzyBPVXbEPpVDA2F8SVZfABMS/3RKq/GMwP
`protect END_PROTECTED
