`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihLtGnPKHtv+/YCjw6XxLcnrsb6LBF1NfU2ozoMbutXWKvpjnY+8gyBCEuGiAmjZ
B1NE5Y28/fULNLaC68gqn/Jis4uS/HytsgaOq1FC1OaFmH18vnWKZj4GDMX2dwAa
7SBgeMpF9AedkQ6VQP5cjwtKkxWxebFxgcC30VEjwP3gAOR9OKwK3we4fefZl0ql
zTk5aWjo+bTwoIMTU6fMHi1JvvnbnWVNNKQ18r3SzAoCSUGyXA08fu68eLew31ls
zidDT8Qf5iFkee40BSyP7j1u2f5GmsNoQk/jv4X+t5vFmLFg0v3O8W2+N7QnH61P
yHqNBJBd0KGoAcwyDpjBzA==
`protect END_PROTECTED
