`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IDOywqikM3BTbh2COFJ7TGadnCY9X0/5OAzaP+kkGHtotZr3azGp3roiJ/HVPqS/
FOEVcBGt53yDLdZB8rYDzHdLlqXYv1nARFANk0n22SayKw1zuTwiylXeX7l6h4V7
ncpEFBJbT6lP3dfVtFglQb6mFnPhoKRn8XYnt2m5n08tbT/w6Xe0GonDoEgvxat9
Fin3NYcaHtdybZW9AvO2Ya8+5f+sj561508UvcbbBztCXdhh15GWvyI1g6CXyOGJ
KhBGiR+yE4vy+IGXF0W2hYzblYDwwBBRP0Yw83W9WWFJlLr3Au8zGHcRIoIFZ1KL
NEUkK07q/WXmSQFyUcIXsb+JO/S4DZz4PPHKThosdt8t7EnMT/aZEounSMJ92GZ5
xr46gLtBkUZQ5pY+VNZn2lvNBcwd1P2Wh0dw+L1P0M6Qwg0ZclJmBhk9XWQ7DGzD
TjLfZKgehJBTc8elyAzi6w==
`protect END_PROTECTED
