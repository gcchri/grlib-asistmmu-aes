`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMag47L1oLBinzdgLUAekSvZUIsYrkRsmm3u1wF7tUzjTmwcwHIIPWOc0zIzTnvZ
OT+MoRdH29dwS6/za3XEpQCMStrRLUUE8i/2pg5Xvk9wFxDZ0nCn5E7jEI+qgcyE
vdgynFU0k+ruDarFiYsn9JsgaJ+97TLNM8h8TDxmeGCt9hx3H1du7mepnCVpCdYu
RiVKpmdaLxWpuJNr2Ong78A4gCgNxDkYnfKhpX+ncOmMnwXwrUFCOXPddui7xzdh
HYvW4ZAD/GaJ7TmcqK1XtlosbEsx3KqeIc7nKMNkjMvIqBZKXJZcZ3BFaUYuXALT
2DBSsXsUU8pZWmvz+q2XW8hlU6uaYF79zpN1Jln/HpxbN3urEtU30kIHJVeSrQjX
eHrX/R34V/Ioj40hyQu+l347KnkBAMntIeEaE7kTgft0kpPRUEp8d/m32WFaB/W4
falfbaadz30kB3u1YsABuej+HBE6lUXuAKR+XyeXQaU=
`protect END_PROTECTED
