`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/m3S6teZ1TEiY6LHwZLIBXB5lDopkAKAqzaxioVTA0LLIKoEqGyfmLx5rqdASdWH
KXorX/CYaFOkauy4Rz/1SvljOmB4pNdqc6qWgHKebsk7NEY6MOwSSXJ/+L52ubkM
18Xza0bgPwk/ryUzW8WPWVvoRpTmyvMPtpKCu498c8vmkqRtY2g5Ev1G6H/Gbc2D
1sDr+VZa9rCw8fGHno1UDRP4O92To06aNZ8j4Q3an2hxN8uzkCYQzNb7izM7Q/mJ
crMUMgJFCOvnuAw471JRpVhyyTNDRXlka+0+CeK7GNbaunPrMbYxPdAaJSrahjdz
WZv8DalwqsuwEzGFZH0T234E8HQNXQb6n9GXo6slgP5NblDec+ux4PTbtEwoo6hJ
sjMTxrwQFyAnjWjaH/LKPIfG+YDjKWpFXLPJnPFf+r3mAq5MetjBymBzB33qJnAw
`protect END_PROTECTED
