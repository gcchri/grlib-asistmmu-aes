`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJDNUrFwqO476WZ1kKaeZvjrjJ1g2OBU9xL8QHsegeuRWdqFtjUPZCCmlJ0degPn
MnM9x/AzWTJjy2HfCWdxVTE1GhBxnlfEB74srhILUawDqH1RWOWzjmtHZDk/UgWY
xvKCav9FPp3gES07ZvrHtA2Ee9/7+QUFkhG0byvcgVIEqpik+dF0LKbjYn6NxFp/
SICXAAti3J9e2SYtFMwepSuwkKjQObXWD6QNfH5LbBdN3g0lnwtfMSCJLIDpGPgG
DNxMwdQI864VvBqiUZmvMAmEE7zbJJ+TZWu+EI71pEgrDNSwCOHsHZ0Ys4wGvvTV
UseM+KaxtFwtG6WtB9YpJ1Y5KQtaAegbtFQaWbmGd8XvpAxbirzRNmsBS65U4mNH
rwgxSqSoM7uibRBZ88Z/i/rv8Z0YFdhCmWkk170bmUutVFGz1ZJQftOV2bKbBtJU
D5RZVCgEgxIVt7nYZeoYh3KNbKXgp6YcPXWZtB+xBG2OjjDFb1qb+84QCcb3CH5N
rzGzhlCv8wxCthKgm3fiUg==
`protect END_PROTECTED
