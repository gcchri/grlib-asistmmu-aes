`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gee85Wjx5zSbLfnbzjCptfNKeQbM0GSX7FrYXOhlJ2NDj3jijmB9VZhYmakG2ydi
3auQPq2tdOfh2+bVnEh7ealcLOmOHpta/Gxc+0ZPH2H0r2qwTQ5RXskeaHvu+E+h
Om0jQOGQdvSNBYB01mEGE5vlUpxLcTzpqDuO4mum4hYOjvt6yLaPFp93EOQYBNID
E6uMVG9WVaTUEbXCojKJCckfTqS3HEYfe8JiPJ9Z1R7eTgItRgOKTZXNfiFcCK4y
G0Ui2JK+3rEy18kVhZR3DKWtJqJUMSD2tzJbi5H4vFjOPeg82M71V47LAN/Loqe7
bEQ7w5UrjW06nFTn1LdetFIwYS/+EnQzNlqZR31Imx+F324uzjYDrFGD+MD5dAkW
6OagKv/fCDXxk11wwNZ4NZszGxOrYFjQToqD4HX5wxU=
`protect END_PROTECTED
