`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jl29vJqGr0COv0bSF9vCIrzbhyJs20236zGoRQqHNqrz8unvoQ3YXSh26hrNQzl6
L4lZymBKCeSTHQ09+apZsLqwsEzLOITzzHksyPAJjjZn4qZ2U1aw0X2gqe30NVsx
ZL/9MMdlBKxHrVWQdRbyFf4WS/J6jJrTw/Kq78fWwNUrA31MCTpzoSiBJxXMMjkq
KfjXS6w2xgQ0V35EUD8AkiZbbrdkNdRZlHLFA32vGJRTQweB0i9nUrry/1GfXAwp
Nf5kIeoZki340qCtZIHCKzw02sb8wRQbEA2uNM42cOk=
`protect END_PROTECTED
