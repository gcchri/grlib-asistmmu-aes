`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BoxuAsv9nc1OeDQ4vkCQy8uHGdlqadcNP4OQAYoNFVkndfkeHldg+5Tg/XZg+362
rXXNEG94WzcskeS0EXx6N0RiqGmnpeWuMTQPEYPO68PxeHihmCLuRcsPYnBFNKRc
51lfYPaeedqQLdGZV7esC+BYv5fBMR9WPLq/dDDr+YfeoVugLIg3Oimwnlgpt68y
TOje2ZShDUlGlt5yIsSib59C/i+TRWh//kjG/ZVUWTtIB9E3DcV64UIuNeSS2wh/
F/gomFoL8PH9yNpXq7G+uP0RjkyB2AIy/kINHeoms1LOn129OwgjRptjBKKkhYFA
9S9KfwN8KpbKDvx432tL2Oni1SYgOFvrDgHRD3+fDgJnOqcOyNlFcx2HAmB9V5y9
xIRXvhrNZEsI5Nvj2P5y9ktcYUeQYoiZGFys9syOgtn7vntE3Jk5Ba75ixYxdZZo
T1/uUHILwim4ZPJs/s39VVkVMv+LGviUmnid1O4HPbXq4DHQTGseCCjV5mbn9Z/o
3a5XmQqvmTtxMwSYzpXucc2+Ed5NpYTHGPrV+KElWlqDbVfCyr/kUoQG4rl0O1qG
`protect END_PROTECTED
