`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AwGc+dSOujDptF2GKKuqjpf13w1IrYiT9vhtrCed6luDcQRDA1HNCzbNxTkg6ibB
4RA1eP82xBuKmIm7FJmNRD0Hr85I/H2Erej7mAN+bCZiUMr/4/H+bQIxE3TuoqVq
yjAPj299l5gxmAoZx3jdqmgZ4QAAqCt8I3YXm6D/iPqlAW1IAEXQHd3XbxSE+3FJ
gDIdmaCaIZ4IvGybiDDIyKXH8NGz8d0oEou8xszJphQJIPhEXKyVvv94UEx+y5gP
mKT3i/7rpoFfqJSppnhLE2qAeH72TtSjM+3SBw9gR08=
`protect END_PROTECTED
