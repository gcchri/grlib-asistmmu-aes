`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7EUeph6/WJBdLpFx2qDjCpVesPp9ZEKjAHxLgGCW55inYuJiWgciXA9qtMc16Aad
q8m/eJJz1cmDFuiyqC8uqBnXCQw4uH+J8KxRMCSCwmZ8f0uuofeMpAi58rtQPHUJ
7bBgxOC4jDg1xJToDI2ITcr33g0c7E6KfIZRDDnRLE5ioH7UFU5pfnAoQg0fqRI2
ris+13/TWln6AUNWycW0o5qjJXYPut5YQs7njMCrMdn3f4eJSl1wMhmQn5AcQTGo
/++UU50p9WJEx8CbmzoZ3L4ISN20laMrDlNscWDRRi15IF+49LY17PYmaj0gi0Hi
9G9UTDVtsDi7bk3MDEVKYFzvbydoup8LNIapU267Jz1+LHqg4eSdZakP69pJB2Ia
5qRyo1oucrPWWl23N6HkfQbIxbL3v06WK9xng5GIwVC+SNhZ3ZmGQOChI/Og88Gk
m2N190ZMQkDSXedrNyTaqeodicY9rw1NFtDAqP1QuFcKOpUarr6q523kb/PoU1II
7lvEqe05wbR6eTEFIx7dQnMMLXztDxCHrfFZLFk2LayP//QUxrrwYueCOlo0z/dV
GGo6NpcvhUfFesP/c8KQRnaBoZ8UkAuwCp+oa4sAOk8Rf3BGMoy8IcFiOWFU9/5M
WWjjbNKInI+ayTaMZeiXZ8xkBpl/QyLQa2R9BwK1tJ1nzOYn4C3dkdRxNB0PQ1Bc
urVrdRZAh3A05vMQsB56sTCbKN2biMiSwphzoUAzwGDEP/YDTlaopFnHGNcKcYX3
dTJv2U104I5sCS9TVhIpQOBFThVmebNMchzbLzwBt5oH9BuenG7hFUwcfkC+bkCa
0dj18zoiW4L1UDLph3aUhy6bDq5DdaLfj5tnlIMNAVc7cFfCNTyIZA1QdKD5IzEq
E/hLs8U6dX6tg8CzIx6gMENh3WYJqcVBFgq1ankCVOSJJ7r+IllpTWA+rzOrUksa
pCiHwZcb7pm38Wjj2u9scfxkVG2pBmW2qT378ezSe3F3ULBZvBn6Wqt4K2kQlmi0
5txUyjmrK8/BC7AqJ9fW+Iw1nzv/3VUI+yjPd6oB1A33De0+Hx8By+2rrFCN4DSM
rk4RszHl12VMyX3Cagm5iIh9LMsn9icDUs5c9NK2mOSakkeGl5aqa8v8tRtDmWsY
T5szo+U5M95NW/OR5K14yiXMLtaTx57IrS7gQLZjpk+Cnolz941/mmf68kln/S/x
spZPmeJxbuITRH4CWpb6VAznihAfKGYUt9vCZmj7pPK7sc4BH33hl/5ML8qgoVSV
TLnGvE/3vQQV7Pn3r7VZ/JQjfrzzVTSf8kqjcE6aQJsl6nY2csfG1Q1Uhsv0Gm3o
NN045pqzs6Zy3q1L2Wi1LNdq87V2hhxFOfWvOjJMJp3f9MosjYu5sOUfsBKlSqdL
HL3lesnrG1x5FL1JUHOTH/BQ6WJ4vmqH8DU/Gw6DJI9eKKMQK5f6Q8mYGI+llacD
MpGCJnDjTr9LfsknUhhII8nedFgPTvHucKdoUuQRbcv+YGqzYI/nDnlcXNwnYN8K
iH2jV4eR4Gi0FiwzlVVy3GwqUJ1GxAx7ylmFxYNgmH2jYmPvH3/iRYdQSZ8JuzNY
Sj2eywDVumpYNO9jc+oDvOS1b2VJ7niwZjeBijuWdInfQ6mj9p/0eRFwKTFqBtqh
+bd9XcZnAd4qIyphMu8IcbnnBCwQq1DFIY8xIFgNVLCJgIpnAW5LEl0NXcCxqKD5
cML7fKEvvnlr05me5Bf4mnaPfLr6YymEkt4QXmU2GXYfrzkR4nyT0/lxAPgfZDZ0
8mmw739JsY6guBuVSOa6ZeUHw+udXHbEjDZs1NarCxJVwlz/PB0EbTKLJ81gYDbW
g8R82WWGQOjhdOyVLD/qeW/MdErEVBWqO8QDhcT94lql+IA1idkWnI4+0qheRkiW
dFM7/govGeM3a5soSBm9ORIRTQ2/gX9KTh+Dx/XYu/M9jGCbY9QjIPVRjz8VvGPT
y3TQPIRoI4pDwn9e4bpT4f/kzHs6BDVaAFv4RFb8tqs1sCyAbN635Gtv+RIN76nz
vmEfZmU/6CZRjdxaNhZCLkbyKrT7tT4CafzNaMBs5B94Nn6bv82wetzAmn+EqrZG
JMhd0iuOh1Ze4CfUUjfeMQarOmIh+wDe3B3SjoKM1KG4Ptc0FR2YBlH9yBdow0K4
EAJCnwP6WquKsz842+p3YQnP+l1+gIjhEOGXqcL1HDRTXz3kbik6PR6PXxpoaW66
QyGBSddCGdaE4bwyfTnDDmTzq/wUXfPQb99wbJmOMqm4nUHsDd0krcxHN+hI4Bs+
famcENiPievdemM7GSrOVenQbqgKx0A3n5Qb9a3jAIjdbvA94CczWdqPtwLI3Urg
K7LmcH0aUiyVQJQVQysVgbqRQ2Fm3exhnaSOBsVAz3GH4FWYTZvvaZxttoRMq/0F
OagPfU9sYgUA5akr1TLYLdgI8nT0iSBivYtT15dxqV20q80D/HPDQSPbaQqxRr92
4Y7MCXGepnTBzBqonDl9VaD9l8DyGjB+Nh8IAX/+e9dlH2KHq+qum66wXSdNM7w6
qxAKC57HcH2Z2dRzN35zxKyvPVJ+LU2iIlS4MnkKKGDil9Q5lKRwq6r/jjLe6XFF
pQiY6NPMB1hTxDKaQk/Irzn/NwBS+uUrJqZ7fvsZrPKdsFQ1vP11G0sOw/ITrad1
hkojyhikQrsFwNV7IVbrDpk4w3PHDTYW8hPJLd2r4DhmKFEcqRy9+Tk1Dh14b6ok
PKBrvFlwt+B+ikOkIqyhwYdk83S3ycPtdQmhRPHx+KHrpGCks3EjdVTW5anu0als
kWm7sMZeN2jAml4dJy8blInWO7NIEVHiJhVGiQg1Afg/xuFisWEha/Hn0eklfkGr
yW0OmghLT/Or+veZIjn4PIwQbVqOTfRt4XFXowXzNCWdfeg/zaE8cApanUXqU48f
FG/yOlUaHeS+XBHb3oex2Q==
`protect END_PROTECTED
