`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A3W4eNv9BIOOCsB6aItgEF7kI6SF/KuMWUNgV7K8rvhI0Juv3UvUXd6ycUY5cbUu
JUMYJRfVAuzDpmyTvQhgz1rpY96O5KgmzIGHj/M2LK7nRsvy5kzKYNGvB4EjAQwW
W1g+3PDxLWgyjLBuRc2r4/tSLgWDWgVmtEYAVx4lnvfXWVF2WOhYPfm2fpVl8qdj
5jeZ5fItXfsHPryWyoM8Wf2M5JOuA//v381KT85t1fi6AWyWkUdPKvIRzgU2WF5/
ddZaoorT8OU7d9TGX3jrBERz+/kCQdcZtykQXpUg1ZZwiJ2OoNeQczgDZtkfJ/6z
hRaDLCRXmZiF+ONjeR5zk57Pry1AVQmKQGMHpyuR3jY=
`protect END_PROTECTED
