`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/A32BV96b3Mv1tGhLoZau9HIXb+3oKaPis5mB1qheHrCIkKxJ5KouBaNEb4FwS5V
36w/3MC1XjQrNLS3pKgRD4vkOo8TW72z2sxbmcMzwZNesOIl4VcOdwbYNRgOwYna
CmvSCnRAasGOAUEvB4rcOLY8bQDazhSkHijHDzRyO7QPAITdst4UbxRnDyXFnLtd
NW1YYdyIWNjjXRhml6IDJs7aO3uTbuIka8KmiWSHKVcZetNRmFujrVQu1mP0ACOx
V981Klu/9eoFH9PdOZFem9pGjC3O/+fM9o8fUqEnEK6IzZWxQqoEv7amsVGNIG+t
jRaoLkfTsyR59LFSHdJvlg==
`protect END_PROTECTED
