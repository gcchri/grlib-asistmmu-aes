`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6iKbsZ5mp+YKSjWkiFXmNd7fmpJ+1NeeNnNHppWDEACzKThl9eyuGEWT4DiFH8R
xt6ysR3LybXHLWlEQxq63tOjhENqq1JVx4InF5AN4h4R/iIoJBNSICqLYlR+XlpE
oWy4U3kTXBq1lZfaP2KrPo2WTET1QNsNotpLyFExMBMmrAaVPnzBv5YsNgv5HqCs
WRoz7TTkgcCIZY4ROAZzXg==
`protect END_PROTECTED
