`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fLf0kfHpnSusEPCpYU38We0KAVEXoLlgkygWuhNVL2bHa9Z29j4nbUPI8ym+vAmF
WFOHqb0SFjIk9dbN/g26tw6qcaFIo9zlybZ9OG8Ox/Trb5NPRXCSs6UsLMxeOVpd
v4NXynqAyFNVGFDq9FnkoLkyOV35Kxt6XlxM1QfL3e+flK76+iv2ewD8RblRLQb+
JTrvLVzotNp++ipgwa0Vw/2CiIv6HKfttUagqJjNarCQCwaPFmS44c/KyziKwWRm
DdrLPKmEKUl8+eYrnT6tgiCpBSNCv0NfIKjH7jSayNehKEdDuwa7wnskNVuSzup2
knakOWKyGaSlL8muoaR+FKKmC/zVvX9fbJK8TdHV06j0nHe1oycPUQ7ags+kJ5Fm
HY8+PRO1oy8mC8RxiDWV33FZ77x9e7TJiG/3GapWJxjpbD6rfaS25JkTCh2hdwY7
ulM+hovKnN7IGA0u244A0pE0jLy0FV69e4p1musrgb+1VM9lUp9ZXExqwD2WAshy
ouMSjnyS98Va1+/nxM9cds9O++uEuLW5opjfLb1LxuV5zkbwkdPolPUAkLszcRF1
eSaDTaAy4fVfuaXs+/3NNnGDLC6RBTvokAS2qpWMMSv1bCq9hkKTSij2wnCx2ihU
8AILwzCN6de3nGhoVWaV1+YyO2OPsQ6oYUywDRajZNNETa234Z4A5wsOkyUVVvLx
hy5/OPcrJKE27AvvGn2FJLqTvfFG7ba0EPE1zMmk+eGI6SW43Rpt5YH6R/GBdqYi
Rs4/UjMv0iR0Q/45haR9vTmY6m+pmPKH7GCKtcWaTpeAexFWf1WM6EjUJtWzkyrT
KBG8/3h54/mqAXQsz8KoDr6wlSM/YQREea5RH4oJH7UcHDfpQdTlbR3c62KJGRnG
hYXB+EosSGO9ioHunN7dZaLrNjaAOIqUg9JRNWeFG3ivVielzpmgrVTGLdOp7TnC
LY6zBeP2ZLz2j2VYVDcAnjSyZi0Ssm5V7QS6zUaxCFt7X6U4H0IRULCaccxK0q/k
cIexcfFys/tT8ZuPAlM9Uw==
`protect END_PROTECTED
