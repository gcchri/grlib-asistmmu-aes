`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7awN9D3snBfSS/KWhUeXB07RZK9axLl6x32Lart6roUwiOvY/0SeFzeXO8zU0SYQ
1CjQiPB6rVLCl3079cgquGa6MKP3UW8diclB4orGIFNBJbawfQy4eJWd927TZdtP
u9dymMRGvod5RSGoUYKREnF1OUro5u+btqqFNQbLJ+hXFcT4X0jwF/y9GNWZ6/8N
X7lo4mY2+/hZH5Qmy66PYl916WD5xaP51AmxY1v4NgVC9kr5O/V06ZV3+s6kDeZp
k3DoKcbmtTLVrqDpsMZkb5FTC5vZAt0IW/dgH32F9yedX331lWrqXPkP4kQReniJ
1A+C9YCmw6jrn1P1e5di2WKxM75+eWZVn+L+kkjMrJxbGIDDN5q920dwro7q9sl+
7lyWRR2qhKe/cy5V4vCev7h5+hYvvFeWlfTKgbwPNyI=
`protect END_PROTECTED
