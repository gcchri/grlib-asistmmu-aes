`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pnTU8hK8xtWEyEbgWn+2gV0Wy3k/I7mFIPhoOmhwDrVR0MQGKBk9Sxc112rNXB2e
qPPdZsIKUCBvCrfpEc0LJ0lF1fVrnoNUCEz6NteLfamPxATszXlVo3yzQGMGIIX4
l4knWAPdf7csrgA+mY6n8hFImEBiDxPD7lh11MR3Njv417QWBOoj1IhIrnjF5bsx
ZyHnE2Z0aeqtgWGckw3KQkurJs3A/Z052yhMJLJCrLQ5kVPav3hCOIRGs/2cIe6w
vmfNZ19yI5oGcRPRkRuGtA1jQjqcnpGmitE2s+0Jr0kjbJ461lVU1qc5FC/IvT5o
k6wqmx5kNgypZ9PYT+gGgTB5t1G0kIpbqsleM1qhEK7d+G0p8ql6ZCHbgZYNwPJn
`protect END_PROTECTED
