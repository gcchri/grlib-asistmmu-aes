`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GfLL4tW7eJ00Bvb/rwQdcZujxvw/M+OSV6npahE0g5NtP7JOPiFlgV669V3lyYTr
s3LdoGczmh1H/Bh56Pm2GX22EIITSys3El3sOtIfDsvVNv9ZvS90mWz1MEE96gZz
DCBusKwh1X77+9sTKITNGmn1egjbfSfTPFaELNQ0QuEG4DPcmBkYZC8BIMznLBtl
+kKfB5kjRPRarZ9mzE1BTv/4+k5OMEGgU58r7R/K1lNd8zZb0YFNWtoqVhS1a1D9
bAiN6opNZDZuzwpsJbiYF6Vft22f8QzMNO+gnQJ9OqPfqnM9oHz3XrMOT+AI/+MI
Ww5NVhQLtRw5thydIx8a2RBAWUFObVkb01Vu4H5atXUQp3HQ8BwsPq8vlD7DUAoz
Edfd0kuv3fvV6D57nEFTYWfaWGoQLwGusjp7mXfsrYfg1GV9G1s87GAj9ZXLAVBj
WxXS7RjMvDnRrJzHy7h2AQIG8R/WbmLLv3nHZiHXzrMJZltXbJB94MaQZyMpoZet
FKiBEr1T1bbNrbV5Y+QUgxiXNAjFlMPEKiiKx0OZEgAJ7+anYGGgN5FS0ZIjV1oH
FLJeMdH3JhQ1ePKl4oDD22SH+DUwR5HTIc5FwIjqws8=
`protect END_PROTECTED
