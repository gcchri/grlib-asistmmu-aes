`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+EcBLRCrmTC8beVvUCfZ19ew6LYuncx+2z60mRfHE4rhqNaxjmhlo3qJWTE8q7UL
cHATcOx+cCiAEh7dSsj4uumfvdZYbCOJ2qSF0x0yk0o9fHj10o3++X8M2gFvl7U8
UJZZuHjZ8u5JkJOcUdugDcZ+4eyitmbf0XfawrHswtSG2TY3tT9MzGTzQyWzsGfZ
V73yB4q18lPp5p6iN/9hND+PaIVXH/wYCn9jz6Kj59SBJLaiSaz5AV9cpIlNrrc7
GOzkzxQIfedublv/nwPPkO7sG2SRZ2z+07mnr7aTkpuj6MxJJ12kGPC/xTchjESb
FRTNKO39sTM3dt7WxbtER7UD2D02IW6eQyI6BfA3A4UoIZVJCcWuwPICVQNqFb8X
99LzNukxo4wfLEfnMePx5k29wBIU2+EQ8SIHRAtgCf7R85NXb5R0HeUC4Umn5rAa
`protect END_PROTECTED
