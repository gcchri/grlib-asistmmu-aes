`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IR7AEr5hvepbsTju3lK5zMUhrpONG/z7SFjYzC1R4rl4KEKix7yWo+ytkwfrbUcu
vTVMEcFE0WaA/OQcNm42Im/4O+tcxJv7vXKtnR6keBI+tE9Y2mhnLogLCv5lbVnD
YnxoBD+Mz5rlm2Jyer0nBEWffai6fh9cBadsp0iVU87kHeERRjxAq5R9P+FtKwDR
ojKIJi79zPJ/oSaFiwc/ATR8zyAhlbMQz2dUw8KkLCWfYaDtqA/W9J7OCggK+xrx
JYURmeDWy64t18mi6+zOH739TefD2wZ94X0xDZPsw2bG4GeNBzctBVRYqw8Nqzmi
3jn4Yra8MKM/s7SXYlk1r1R1QrKSNnPtWxOqG3sS5x/yWzoTYMBQKufKNx6ITao+
KUL2t2m4/ClUAVfpMKHhJfRT+sztrcrjfDS7zI1TchBVjk6valKwpWpUd3ZFAmPP
Do6ALFelNsK+s6jOcbUJANaqYHXKC2758pP6+VHWr96DnHnqggLpF5jjhK1PYwZo
jU5ftBJcgsjC8mOIoik2A6SVJJEADilP2sooNUoYmvr9wIshdZ7aRbZ4YL1NCmpC
QH0YffxdSwKenUOIjNv0knp3I+l06K0w9kJVraARpFhyeSCWdKWwfhlGW7HApnT8
VzX2Kg5lJNxOAQs276kzK2mWY18P0KRH4nIvbudRWi90TDjKo4uegY5B/rap//RF
28RlloZvADBUq9xngnP+JdhWdujUThmjaYDze8LyBX4eu0sjCyBBnYam77xtCAgE
pcYhonlPxnIkcoqGmv3ry5SRLFc7Mb8Vz7mtJh7t1Oyc0pDetWa2lvciWdAUJSRL
HRXhYEI2YXpaBWAfTnm4UwL9sFqcYgum+/NKfdEtcZRV5UiOgnk8SnaDo4ekdIql
U9euk0OSZbYqbXpU83+oda412u6UgWNfyQ+mqVGs5dt5SaCz+YkiTvpoW/HUL41L
5LR8LgAmMq6aWgoHN57vAalcxejuKL1CzwoBWlnd00bF2utbkZ2rTMKRv+aqMFXg
Ubf8fyUfaGpSYiourbnoy+RBf4xhjJyrLB1UB8OQ6rEr1rG2TtpGVU85jC8CSgLT
h1JpTM1ik7hpFUep8cxsbDxFSkLvXGDR3esa0fJfDEQM3txO63Oq2Gz3d/P2cQUz
ZsLypMm30Pze1oZDg5G9zpeIzHGHWyRWA1FsMJ0XuXAxvitZbqU5/ouPLdvAPRAb
SniDP3VhL517sELKtiuC9BhGSg/Oj0X6W7xCKKKOYvnXiElR1TIrZHfV8pruumpi
jrYke01FmCldB8EGHpe7DvGswyCqgSYvnh2s2Aid8V1Iw9QE0G9caJ+ofX8PYxjG
py6aYXk/wIbGJyIQZ5xFVsN86N+EC71UimEr5w/vjMc+Y5ZW4AY0DIu+t45cUoNM
WPyBpysJUKt9tbRbN8DjCwMD/q5u/J2N+ChLar2puJAmCm6OA5vnBgr3uGqKsS6F
28lrJN6wqi3HNFKBx+vG3+7KN95NeeYnIyiDAeVO9A2N4F4TOPxmp5OVeuQJMfve
CKdGON3viT0915n59MIDHYKOI0U651UQjFw9Tnh1a4+mkbG0KXwuSMkx0mV/nPzY
juuWNgv9t4RBwq2wc+8TnupgHSlkXjL2NffOnJStXm731D527nFJHcbHFnlcDB/N
BN6khMbZTRI/KSjDI6wRpctR+N05sAGqdbIEJKli/bip7p0w6OMeuDRbXkHDNfsy
G1vOLYM9KXeTLmzu3UUEPDAKzDg5wQ90D24Dd+1P6GxpXtFDgc8y1kwG+T3GuYF3
47mPJKXGFe8ox5jvGY2TFzesBiKnkaSpq0Jg07fmHXMvUh+YK3KGZkxtB8c1WTlv
dkThzFwkDqsUPDfs2HhWroGPRMrDvtBoKmhvXir8ut2ZfHVewG2iSe15xXe8qHOw
nrIqi30cjNV8Eimhon6maZw7ZCPrs9bRK0q7pP+sPXj/TqMtTtFy3vUJj9Y9Q9+s
PmkV+SccYZ6EEyyRmk1QhgbPg9OxfbHz0JoXH59XuCUwAdJCCLUyYksP4OIqHBlE
3wcdzPLBH89QvkkSoNQtncjNQQP+bPpl43hdo6HYlwFORgjZgnUyrYzLmIkajJFO
9vq1uyMqYv9DjYX9xTI1q4LTe3UnozoMwZS7mFFb2H0=
`protect END_PROTECTED
