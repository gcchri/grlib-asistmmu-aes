`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gv6RfK3fVauCshHuNjeCncxMqOnSJjlCQkBK55MaD3qLuKBtOv+/QvO1VPE4GZcl
7XD4fktdbBs46A1KX8td1yFoGSSf56Hhu+HHb9a5XdMQfRjlNPXvECbefi+AGSNW
TDLn2dq2iNpAXKvmEncJimzUJ2ApwK2+7DZpHD5YDbuQMCXbaAcTp8uduZPSWTgU
ZOOB3aUkfp7rX6YHgWs/W+bJjRxu3UXBU9hSvNLtLevAu96VjOu/n42jDPnyiZjD
8qboRalbtXZlEaJZzo9VOgJI6o2eRiixHqX/WZNNZ3z55qPlhqvJ07+pyVb8Sk3v
GUe82MtGDa+mSRDXohtMNCPT6sacrQ+0CQUxv+8117hC0ClbRFtJKEuClXib9RZQ
DXDIb09OS1eq24cEmHCr6I3YseIUcK1I0/pAHClCCwNxcXub2UFllDRBAWlzcYkY
LWa0hj5qqffJdN4ZRc6e9n4XnajG+pZGIJA6DkEjf4+n0VzcRORyOZkMP0LVFSV2
4jZno3Relhdvq8yxRamLa33yi7sxcMNm8P3lT09lsfSr6taDk0lIsa4It47C8OUG
GzZ8iZ64eUvk33nfrh5dpmJLwHiFB2jeBEQrLevSZzIs0z2BpQN2pKpRKBIHLSaf
Vj41VxI/yqIn/9b9dRj6ES4LZIapYD02uf0Vs3DKemc=
`protect END_PROTECTED
