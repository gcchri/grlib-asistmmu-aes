`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqq/KsBUs3uZYmci45CoOHnXU0XKESjC334m7TD633AWeJBzVMB/RjilfvFFUxpd
FjSfSdlkD/KS0vUITeEMZu6ImuV70VBT8GnM6CnY0m3td9noum0ujGPzDvqHRGdQ
6AsGj4HhgOhc/ZzyB4nker741vNgkvDvFoNfZuwuLupMakx2b+3vCZ9bW/ZVCD8R
s61JzhBkpelrwQa4L63qPC0fq/BmVhxP7gWpsPzHURHDKOhq4ulR8RgxRx3eVW6M
eFn6mbl889Ik1RIZxyj1gW932PB0gw9NJVQ/fMK/20xw6MOYGlr+sDfH8a/K83UA
xjg5L8uijAc7fYtIlJT3YBR9kCdeRzBLBqvo/UnyI7KDSYS00lwHMGW2cImOEX0R
Qq+Ju3FLT16RTuMhgNABepKgjL7Wuu4vmC0EL4Zgq8VEkdJ+w4bPvFLeC9uz/gGU
WqJXEev8h98RGCRIlq8WjLMfoCef39CNgKIQaHjByzLOWGrVQitwCUaR08HW8/r6
v8zZbhOuT+M2+ppZmwhxg/1rz8Aj1Ia8c42Gf/4HXl9Axt9mGj0rG32Ttiwz7O+5
8qveQpJwvxNfk2eeEjQylzQbZQGXZmbD5mdG3SAwudsEW5N+SEsG1RmxOH8Lmt3K
54d5Yqlcj/e3hBR+epFA2w==
`protect END_PROTECTED
