`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t8GRmBxflS7DCST7fcXbXYm9MQIloVeGxw8F3rm2i3jM4lNLFCab2B7eoNz6Mnrx
+0bSnvVe7F82nw6SGE7VKdKHuGNodYX4yhqSgbgG2qzaW0FDVi2oAtAjhSgSWAUd
WPmocnXPJDbzdyV26RLLRSMo9vsAkQtYnyufSPBiWCOepG9SSKZ+U9PpSMhDSHH7
JpT8xPF7wE4WnyZrYsRLVkSDLsI8fObDdgNMa6gdO+s00bADnxurtR8XrySTAF/d
pWb+Ws6Z+j5Xq5I2doRdMDRCpkUhV4We0RYEOXo349WdogQT/s2yu+zyy/BZQxrz
h3JN/qLpx3U/YpFVfNijtXnO0ao2Pbduq0ct56HpfpDmdmCTukM5TZRr8mtff+y0
D3qNgFlqDNF8hW7Xjxr5qjsEWCX2GOVYFLSr4ykEimUrmggwEloEKyskF0yD5r3+
1yMlSerIk6M3Vz+rwe4Jk25j56I164TFGgRAmyYE2lQ6IA+tF+Qcotrjno1IuaJR
8KLbThatekUXW3OxWFSIbjAyg1vVSZHXbSsGgk+wznvv58uyYBaad6bUX+UGKSih
4aR6C0dSq+8kxG/gxr9WsQ==
`protect END_PROTECTED
