`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JH9C08Jxk8eSFCMWhaZ1T+2W5ckLzAV5GWPuxiHdOkq2oxaVjyeW0PMnCRIMRqfD
i2lMAYc4ZJurGhOQ34lY69VHapqwkGS7UVeSD1EL97IyEwNdrtm0SW8q1t0u+t27
yKULLbO/FlQLoeRNqHwv4yEa94H748P2m6R2ieN3coCoUnxvTxaUX5F2xqFILB6V
bkF7WZOg3bodg3qKF66MnK0/+rfGtDLqSQRjnzCGJkOeDFSSzfZX+2DZkSUuKgJU
87+xlUvfgDDNFmrQULKqpUvdfnE4Glli3N9DT5K2LIepE4jnWen654YbunBhRpfM
SqysiiHamxKLskHHsor0KAWWoA1WDpFpPvhI7uTsFocal7wBg6eBuO3GeDCgmvP8
J3ohs+XDuzcZnbQCP4Oj62SJJPVW443MjcLtphA8N3xjdYNMXDPQnDd3XcT8zhvx
z57FJEqfIMDah/rwPrPVXNiwI8bKSywgSPz9sqcJ0/pxcNK0Oq8S16H3niNNi/bn
jM97LRfbbs4AHQsGmtvW2WC1wYp0ZYgnbvs6McmFpvYsb3IveBaxpi144EBC8aIZ
UChYi0QjtzZD3zWSWCUV+cLhCh4xypd/+XThwvI5YH/r/nr6PjhC7/x7JftBRGFL
uRDOat9ZRw9Bq35KUfhWf9fryKg4F/2rq0QQnCtk0d6o/FVwpEyES7eytlxTP4t0
zjPkwRwsvX+qPXkhgxxpnv6tHdWt+IXNJvk287zsZlk=
`protect END_PROTECTED
