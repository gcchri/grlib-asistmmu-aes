`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AX6AvQyCJgDVzq6RAlxryRjEhHW3o/Gtqeqf/YPAfPjjxz58dqmwtpgJoFavze+b
NSHM6QeEqzaluLneUEan6klXW5uR2OXfJIsvCwtj4q26YqAokvd6D/UzSNdG5WJ0
3sfywymQjHn4zSyUBLMkXH1DAV1RLfdjnwZ/nGa8Dkx+diIhIaQTNBZsYvWnTDvY
fUzF8QiJeXVzWLxrm6t2zim3TBdXDU7qf1C/mEceApRX6ndyFbxNxvjAa76ZM4Oc
+S/9m27TJ6ilSswIYt0JTiGRanxmbFqiaXNlyvQ+YTm6HpQzwQkp4OrfV4ohzOB8
md/kq+nuoThegPHjbbuLfEO8b7fEkhsSjtKMN/56TyBNJCNYZEK8M6yWeEMlUP2C
e/CATNI5G2QInGrkdmyfQUI3nXeiF85epAdkir6Pzdy/vwbTFREZEadMW1lz+6pC
rFcb122H8BFyIIwHGcBiEOhklEVuKMjkoyAa6FeHeAs5n70jGHrcRSr3mSmSeBnE
TXg7MaCDVQBMpWxSX3FIXuV+krrD2UOQvOhFete1ncBsi8F5TMaAGbybn7fj5Chm
d7JUo01i+ZPcsIpWwtESAquyEpNT79rReb7mOphshych/EOHcGHuWbDvxJoWqDfm
E64dNpkixHD6BndWRh8Nmac3vDR6N6/9aYP10HL6g00TP2RDCsbiJchTdJvu266q
awCWRSZX4F1crH5X4FjvXTRjk42A/1sUmDMOijwVEaZXkR4A298LAHWY9HI2VkTf
C1uN0eykvpqQoMQAWU1eAkSlRP+nior/giaGAZEiyxNHi3zMHdjmrnlGzE5fg8Rq
wLynP5oCAoom6A+So1qH6OQ24LXuD7WsGgixE3eKPcAmvsEY/7WGjnSpHY01O4UR
HTwKWgu3PpdCr7AJl8DQ5DWlMrWRz9qa6GdMRHWlc7JrpaRRpWOHOPk3j/8lb28B
6JnO0KzSC0LFE4wz0DotsvhE0e+cbLZgq0prxd989uYsd7zRGTfPhdgAp9wCX72i
8AuT2C0B5cmo7pH/9qzC63JYnVf6ji3I6NUY5peJ4n5jxbbC7zpm9DNcVi70u34M
Zv9Um3or9j2E+d4tkunhg1WCjgRN8gVnmtRF6xV9e6+/s5rvTjoqb/mthg7eSnLF
keBFdf7gSH7f8b0R+bp+3wZlWathsV27+MkH65HcBO89h4RxuOxkhTY2McpXoZbM
l69fVJF5eYB6nNcP0IPYw+s/QD33Z/U4ViBWnE3eHJ5jRkPTakrb1kEPbMW3u4rm
J9w15gXKk+87uraF1uYZ9uuUs4GDMpBnq4oa3NzcLpEpoKJ45JZyXHcEyhCS31A9
5KMfbOYv8zBdX3OuH6kqUvEm8+GIR1+Zv7XjYiv5gqIj7a+zSnBNoPE41syJRiE1
5pwaufqNNY0L3R6Ny3GbUF49z2tXdvy6CZb4cETg7LoagssVUxNQBVo5ihqIXD2N
eMdFoiUfmQDNzfme1JwzJldcIqtA9pTu0gDxqQ6AzTSq63dW7agkdKHOSFVa92NG
poWKOBtWklq7ZqycWbyZtJDmIEjzdhz+60o8sjFrBHeGWktf6A/NHHj8TEFXlXle
rfN4XFxL8HigR0Jsk2ufoQye1VKdIAjFmhBJaL9zrc+UJEIPFCjRbKiIHUXjn/is
j38yeTIjdsW654iAQESAKDaGohcFHWNg/UMhhw0dSwSrLaOSIbF0u3PsdZ0kSzos
LkCcUnAAi15N/LG3J5m8Et8yG5or6MDlw4YX6n3GRPw=
`protect END_PROTECTED
