`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k6cp8ljRxrSSiWn0+tJDO+dYTJXqNjDoVKxVLh8ETu3jCQZ1QdiUmQjhsZPu7EGx
U1vlDqgH352rqfX2xOZlvstQ5z0KsOPIxI4oBs+ABntm0j5/WAhbnITdYo4rW8gg
vnaN/aT9hSR8WsKYd46S7jn5Q3EnwHQYF1vfD1vPXe+2AI8WuipsnI6jg3s06NLM
z00KrXecGHyCYYXJJVdhYLfxGHqRsWpaXM5K6HiVPIX/pcDzonRt4znaFVRgDDw0
V3qinHN5pg6sk2/RhHgtPJ1rQWiytvo0GzhHLBL7cxUayLmliban/maZvpbqRJha
Eh5FigQg7wxCnLmpstTjXqRRyMzsbeXq4HvytcwaT9ZoX7/lZ0cJBVh3o5+nk/cw
1QbQactdla01xhyTAdSYQawJFL7Gi92R8IsB/XircZxfR2eGYYVUah8IZAtfPIro
FdLW5YzfQbGgqp0yZjn2+lbYM1yEUcnn1+AgthLdM2+qU8pd5NCqhSZLQebG9CGn
JgiZ+udjpBxHidLJGnnDRWDLVmoW5DrGNMgbKtsBqPqLJyOqUIbE2iWjD3mQVuJ/
Dn8wJlTmj8SUJlqIktui7B34t0Dsw+t+wf2NvCNHlF4s7NL66vkCAbDS4+knTCho
w+o+kiIjvWo32h3HW+BfNOXRFaDIJ7FNhF2WQLOLBZf7AtSi3NQ6BoVJdjHAncGG
TCfIFmt0HWqq/kY9/ab0nUv2H8RJc6l8ggULTTqXPw/TkNloj0cji9MEnkkhMpHf
wZMRNgMM83s5fyckodiK8pz8WB3l+FSPvNTlgk8xxyy4Bx3aznIQ0nRc/W+2GLG5
KrBfWyyBrW/aNHcN1IamP0gbKOrUcUqyMcXiB6VI9IvUZg9z/SfDkmvg/bSHULTl
qbfCnalzbjA2zqD1wbvDgrQAzAvAWaRVCAmf4z7qo8bUVZgFs860guoMZVNF9KfO
cd1sOBUyBoC+VHmaxR6ug3/dxoLORw2Vg8zc20GxIlz0EKzwm0zFkJk1fvT6FNZU
73lcXI4b6A/y3O3giL5mBUKG00JmK1Z+EZei5+WiKON8ZYwM8Rclqv2c2+QPMaK5
ghg8FbhJjYs9FKp6N/1i4XUb45QGh9cfagH+WbE5kIVhyGuuniBS8KmZKNJS+9mo
gSrSHmlj+l9GNfH3r1Or/tJtp1mut6tq9ON1Y8t1N10NunEUh55Gl62GuqDxRlrF
V+PPmxA4lx0TXW5i7IUDbRZg5Ntjr/HuPQNyMbyRShJfTFmqQ8mRxmMEUIp3TCBT
EQfw6itHzvG6Al9wjANMlr9nIDVZVqSLKhmY5TQEtvjCDeVaFUaVq+rJIkWbPdmG
cZbXtZae8piLuCLOTW+WEGBaIzgs+KZdaw9bzoRmyTePrE7ycdIWtf1y+yMy1iWa
RIYnO2c21KqBLtxFBC/3EfBC1DRbsL5WhecGBf4W2QjefO6IeaZ//g1r9GoB7FU8
c5NNTyXRyQDfuNUxN2xdBGJCGFkTH0zFwFPBsSVvvD7OpqvJNil/VRBuiiMHGIC4
U5DwxkHbBCTz4e0zgNwpEoGWlQv6mdmbtYY5jOmZQ98gOYTpB0G/gvaAvzvQaJUH
INnzQ2euxA9LL8H2sY7ajMzB2hZkZQnEQx04yw3gcwhvHkbR1FJyZurh4pHJWBFG
5FaYmByi6g3HuMgxt04RDz5tNTHbiv908r5BhMfGcm+K0PbMx6kNbKcyBzTeA5/8
OfM+EuJv3bV/9zLt0wRcTXeBhm+LIFK9bHi14fCLFume70Im7zY31bmXR1W8wMTJ
D/ZPGWdT8BPPtQFar69XO8E8cxgvM2iD01rIxiKTQGnrcZMC95TVfwW2wM1mORlW
OOCGAR3I9czDrg3YLTmwRaHYaE4aYaRMQWmAFDSIqum2mWpajncFE14GuWXzGDOC
OdrQ40U+GhcAD6PyJonp3aPTPLSiZTyzfkHaQe4IL52aC2LSndmgMWc5PxZ4cWaL
Q5rejTsdvO/L+MquFoIJ/+8HaAjHKeCqgK+DqsALIZ9z6sfruEigg4in7nOD6X1A
4Pwm0xglnwU2ooAaRwGdWKuqlYf/ERSlcQkIjqxDR3mbuyz5uVm+GHUothg/TRxp
5vyrmU45D3XoxBc02frzc3fhRJxzgwto+l81pGMcB8dru8qKWxDn083epEwjNzXa
gNQ53TijoppVAGBx4KvE4GZxPnCRyWNChl85GTRO5OPTgdiKrXOqZlciXH/Q6lS+
Xi9QkuSYfmNq32c0fLTB9E/NJDGbeamawZWzFJ8W1D4gEQ94XDNryQtFjLs3np/p
B8jWq2/JJcn5Wuvy0NCz9JxVZ1cDe2SOW27OP4dzQp/jFld6Fn8Vjt3zMRnDPC0j
DDRlsmRBhVVKyjP/Zi7FI5ZscxK+oxFheKu7dGfEuUc8Ax5nSaAARvBIPPFKCrSN
8NC7akoYoz9fAiP5ZXa8UzYIuyOdU3l3n7mdinWS4SMWiYwJYZhG4/fQkeIcGUFj
jCm3zQ+qdA2eMDbJG48oDSUzfm6L5u7yUxqaNlp3CvWabTpzkzOEInmoiUxsGnsY
Dd2RxvzguENxTEF7ozRHI9oUEUDpY5/vuHZAsmIRoS2NSJX6HV5z29aCyGqpz2+q
nLBhCWsgu6iB6XxL6GfwZg==
`protect END_PROTECTED
