`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
18m0YVzt/Oh+gHpfrxSFLZqHqyVGF4wLWtfujbmzOWHXXICxkZcQL4vIsqbaC1QE
F/yZ1u2ezRUn5c6rsced3dCPA05iNZ9gZGmSLyFDKoVSQ9jGT4R58xTyYlQ6oa47
xjjlNnVUGfuOToIRhbpbRwMDJhBxN3jwOUP6WFxeFhcka6HaAG4OyFeyqFwL0eoj
uOtKeIShMYz6u+dNfWQ+5elNLv/MzRsPqjnKtbeF1Cj+XbCpFOEvsaD0ME674fi6
7Ton1QQDErefoDn5FiefjkTuaM2hzq6vB6dbojzs3xx3qhmGqbDpsjtVAirNdOq4
2G1bPYS+Ee0GOKm9az7oNyImqxjOPdlY5QYW1CaGkOCMjUkYb5mU6U2dOO5e6Cg/
mDwVZSDwiav2t1EVOKHE4EcLzKs6savRfWki2OgM3yA1Uv0vY4AUwTamEQCpN672
`protect END_PROTECTED
