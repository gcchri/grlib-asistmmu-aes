`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kldqigSX104XTsSSg5RknJMlRH2WsK480zoUJDyNjQ9F2LgkM0nw5QlbjvE93DdX
GsU+3st3wxQMS5vunKqyLO8kyIDrNFIAYBFSwIFL0apzpoqaQHAAFKtgHsAsCbeU
B+uX0rVQr586pi1MS5Sf3z734m9jD1MTqJVLwVfrR00N25vMaIFz2h8vSfIh4RgW
gHT+zDpwx59eH8vZY9kOIhwrNLh2yD5QwWVt5vHbd8vznYTiE6P6Y9bXu+Q2+MT0
wNnq7sn9VhKheaQgYh3ZGkGqEd/a9fLKSA3PFULyN7JB3wHExLT9eMkOybQxbc/1
I4UC4nQdPCirRudcCPvPg+G34T4ooVGbszQBqEr1vUC7g9TPB4A8ZxpqgIaYc32u
nB9CFECY1i0LwVFzbb6ufLMpVe8g+dvzWvjJBnpSx06pRlFaXgcMoRW23oJPu1Hn
tgYV7EKqSfUetR7zs48/tf5evJBPu1NwzcreUo8PFlk=
`protect END_PROTECTED
