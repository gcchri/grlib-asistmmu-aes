`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r/lqfQEm+TfyEzDUpOuq3JXDgaDsbRnYQ3LjkEA/tolTtVBpgqmCHiYrCMvHYsVd
SO9Bx2o7WRvXAUAWCCZKlfMRf76CchQIum5v80HeJrmxPeQH6YDBPa3Z/kTxEC0s
rdJX8Sm3frsDf2mSSibG9hQ9cDCKY3P4pQV6iSBWMgv5fXIJKzYLOFEZFZ0yNstr
X3j3GZ/GBHXQmUInZOqMOpGmZcVtKb7Isi4tOpR0SOlNWEVBl7d2rLQ+hYz1xlnU
A1Er/g5PZqd8F3+HYMWUmeIly2gnbdLgR1+W+54C4du7+4+crWXgC2hoJdrAs6nq
8+7U5guOY6U+vAcamInyTEGMEVDVF2WJY7Y/OLIeUTHereQjdxvHG2dvge8ooj4H
qyUGnhtfQoGd6giy5uiDeE3cD0qx7CxOgfN0VtcTo8YSwyiokmOSRbUqgpI2eqVb
El5VkcCMq2IlENPyPJ6UQOqbPEFkOPNVKwwtIypteH1XNy//3YH99wHin5krMEck
/e5oVRPrHUdpQ7dmCUiq1CtfUbQ+1+NNat3VZpln4XL0f26+jCKJ1nrlzXf2bE+5
iKUmvsSh/UzRt3lajCd4xW/Zqh1VlN6jJuDP79N0CbsNRdcyq4So/ST3zLNKD9Bm
ieHv8EqYSBpCB6bsTOyDgCP1XbatcnUgveWAhCREoRfelVZmO8Lc8hQfoV7tzzer
9oobhQURmR0j1lIimI2VmtJ4GMxSCh7Ao+hwSXcHybCA7GKztD2r+K/yS+BQ5ytD
KShATTCTsSosgxmK/r1ZgQ==
`protect END_PROTECTED
