`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M8w4VPyHU5kU1xTAmp8B/l6kRCO2B8VaOL5ENIoOcNkuLLZfNQhs/iKfkoEvmoHT
iWohQksME5+Rjok6oC7v4lNTFBP/rtOb920DkK9tTWa/GC+JzL9m3UFVlw7+3IZL
U72o9cq0GXm2chQvaLWtPp9/BQc6WyEGl0hkbieKvJu9Tx4hVFbPaQtvxdyu5Lvj
fl4fInG0DTLi4kyKxUlqbehuFpDKUaElnKaZLqAf3o56y2BFaMDeAtXTokuJSuva
pZZ6rP9hpnTtboUBc2Xy8CZjx3QPriLseF7/z4/q1JmTHAzO1mx/hQF60+SlzXVv
MjbOuQ/BH8JaF+Dlbit/Ajle+KPWKkQEjt3cgyyCBH2TYRmKoIA911ARRakHwb5p
vkrio0rPROrvgJY191laJA==
`protect END_PROTECTED
