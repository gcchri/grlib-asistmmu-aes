`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNZEeujJ90NEeex+TtUdUZWR1EjBKNM04bZs5Glf7/780WhjFXm2cAEgS/MXQggJ
SmHGpiZbB1KNKdn1C3YZ3kp2lpZFid1P/own0Jy6ERYWk/xtz03g15xf9hUHojyx
es1DmUJ7vUgadbCihxz29L2jdgeYyvS51Q5jshBMk/b4cK6Q7+ylr0OJg6ia0+AI
Aw9Fcm9HpksWNuPVe7FEjJQpQg4kwocL3Is1zgtNpougduiAN/jMVaZK1Tq70c8S
r93ALfvLbZRJ23wuFraEz7cLWlbtYYYZS63g8PBiAAAugcMU4ghpNLOn7xyVl0Ul
pCw6FVU1lxdxJVrvUtgLiqfXMkELlsqOaNVO9fkTSI354Gf53+4AFq8PCmkYSbMG
253s7z7U8eEyrSLV4Lw8jwYl8JYKj1T5bh5Kze3pGLqM4Axc5l6XCS7OPQyfjTdl
RkujFVndJeIzS7XS1AM+F6sHPuuLcqeeAum8J32eFFXrfcPG4ahsDv2jWuei5KYP
m1APCXjWIPHWb4fipuMjBAThtTmgPOGBoKOigyWpZgLSepy8iWDgZk5hPrVgzyS3
aVRogKcDLasDGrHsisUG+MIfSGYa1deffz1GKPBYnq/9q74RWsf9l08xYxuexBYa
1zBF6FhI3xS0Fm+Y1U1Yrcjste5He8sP51amS/hXJ8VGj5wxV+p7NZ7Rk5K9qtT9
udVAxrG22h4Zs9sf8/gIki97eqLU370xnlsp/FXadLqvcbU46wqO63avIFckAED4
MIvgJxmRNeUU5oN4ezxKNjAm6ocxwT/TIAf8VLM39l89GLKYGhNPleWrN/RG250i
q7ql7YT4z/4KPHtUhOgYAk7SV6ekUIRqroUg5FFKTEMdjgdUbiHHa0a9+eIDJqgB
bnGJJSNzyrrGFqZ+7AC4TFLsPgFpsfEKzgnVhj60YSsB0UwpsApWT4pNCtSgjTQ5
2p5LlE2QTYeVT8jRbH2mBfvO4A41pB0RUIJuf1DgMDnQmMMPvj9bATtWdyYimKT6
xGUYpuTkOCfXXK6wqOXo8uQFmDjrcWm3n72iZo2E+k0CGjgfvyGzokp4SJbdvNK6
bAKmyghvPjMvl+Dmy4lfenTmtzPzYYltR1TonYVkWdG32zIno4EiMI2SyWhiWL0I
pSaAG2mhMkVRDjUqX+DTNbURl8jPTt9y2+nqnVbiY8HOHx0RtaVZFsexX1JOrOAl
Pv4ofMQt1LdhhBWA+qUKCXZMJJxHnEZlGBDfXEQXALlq0vho2VRKW4g+Rfhimrzb
kIisw18lrKlxmA0N9Giw+2pXYyQ9B5vxO26XqSrzZx3S06RaAMj1k0kBeWfFUZhv
TJv3+PgdygP7qqUgwVLTCtQ+8iUl63J9BcOAKMiWG4vvLqBFksKcVOYFXA4OYklF
B7WEfjhMlI0dsQeAcMIBDqkYWO4sSn2Kc6jd3zk6Me1s9qYub0W2FhElCeteUvcD
vo1+0uwdsf7m0XNW5ElhyNFnBB6vqMz5X8gNJNj57IDi7GaStsaM175bx4tYtg/H
HsOgRLNm1/p8/ZdOULaPT78dYnZSF+3AphFMUg6BxyHT8bCjBSPaIaL700ac9PjJ
I6050XySz5C8crX6TzUQlR0FTvix9ZR/Xm+eWdC5AEJEY84etDBL/3a9v6gGoPAg
BUtXzp9lc82As8N+vpfUjBL5tSKeF+Wf4QGEPyaxbNOlLlwqfujN2dnEtgUbNQza
sKrGJSaqKOMGBEKwwcrDyA/ObahhvKLe9oZmlvYMbfKlh97+fy4gDovqjBtPMB0/
cFqxH3UhmkJ2vIYMpDyd6X309iJaYpVA82z5Fkx80fyQxb0qR0DrSe9PUV/s3412
3/9F17rK5+WLJlOvSmcaezjRpW7Fjl5asMiBfx4M3rtgsU+gURvede4vqPECpMyV
7UhvsuDqRpeneH1ne3lubienH+eWUgkmxIyr8xUG5FXQYMvzP8ds9Cy13fxo8va3
Wy58vkAv5VZBaDXuq6W2KB01IOlrHmLc/bIoP8H87Ja5CMgsnpNTNedOIxyEOj2V
fxwomZQsIWR9rLDUoHs2+2xqRkaCtNcWS6g3Fs4bk/2BLFkAVsZu9Q8sYmnSjkpS
qny1ua6Tn1PX20BITqOJ9qpmGZUaYR0Q3y511Gkj5WRk4MQJIko7uPZsgZlmv6XT
PE0o3lXD4P0NCp8JPCR9RK5UTR3WTugTh4PqWnEXxlsmpTe86cay54lBxI3V1WeN
u/1+fAVAE6gPWVtjAaIT99dHNp1woUpUC5FW6rtOKXR6iVTLeE3UZWn22Bq87Z5Z
G0JP5bWKpetp6x7wpUNrCFUYr/FPhJbw+nOkjIujGaq9kQPulrE5PpQiQd3cJDF9
vY+aHV2FU1yi+ps9J7T/20Q36SIqRYWbDvEfauY8R1D4/F9TgtjsrARBB5qNBTkv
w+hzQKpQbXuR13RXIAmg5GHPFLE1GVo79FbIkQ7D/S7FHq5eBqJQo4J4rm1UU5YV
5e7GH8bgJ24KCCxlepzlM7f4jtKA9pe18D2yUhHqJ81mIrlzjJsh5Y/h9b9Ho7A/
F9NnvGLYavT8ZYHAnTrveqiWyhVtpwtK9CDNYLaUr13NWWy9Xgpcab8L72vKdJLV
EDKa5lPont27wCsVzhQXZWDYr2gBNIHW5Re+A/ik6oyhiG6kFP1luedyhK3RqIxw
HNXG1V6BXd4opLzjLMBY1FC0zZl7LNx+iGCQe8McsQkwydrybpA681fw5yGzLlvY
DdiO3d4IxmXKujYUbNP7OWJroQv4i5wKwdKabh1MhdIF2GmDjjOrB/3r/n2CWGWa
DV35NzMEZZhbyIw8BSwX61Z+G1eYLS96SlaPX+8vMX5jw/zSOtwNtnq3JxljOOPL
AxYZ9JgMi/XdWaSmwOlRMA==
`protect END_PROTECTED
