`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61e0nNIuu4kOrfWWCDJ7Dyv8DKkZH7THPGIHV89rm1d5R7mC9hBqUH4OWIY6JDYH
cOu1A4b0EuZobwR8uE3das5M7FGO6ekkH8taqBUiUlbAbhK7BxiMBgTh2mqDU+iJ
yk3I1iRCHaG0WI6LcxW+A2067tLBXED9CvVJ544IHJz2m3aboBFqrCLNtfCcGY5z
YtexY0oGsbPQo4eUk4+WcEVJH8esjCBDglbK7kbGU4TDnsAMPOGAPcFih3n/232g
KPhiWxo+pMO8eYzePlTXs6wDGMi4u+WHyb2X5HAlKaSzOz1aC/iED7OSSoKXokyL
7eePkq/EWkwt3Sk5tLlCvB6CaME5oz3BpzWZORh2jGGw86Jin/wbOrQQreJRnx2L
YTWCWLrygKBG61ZU8t2Kvpi9SrZofgbIEfiRiPkDfNAsbxpGcqniMH0EFvaLAT5l
aRZB7GcfPdIvKBFErgPHrt7u3XubqVbwqy77uGRc/aEWZ1VqqM06d+1n8YIKbtoY
fU9k6ZzJy2y5lUwpCom0XnmBwdyPNwg6n15/oYEnwWK8JA3kue+qpqJylnB3Pr6W
R+wCZe4hVRl8YOuI9JswriHRK8mZCA3a1CuGL6VyDaGE+MJp52Yxnh/gTKMSmPxk
J/nfe+3orHh8DD9MtN+SlzDQixi24BNiD0Oe+BNsJF7YwBT6En7S5Z22spKixTIv
R5Qqmr8SvP5Sh8IBvoolZwPD3YwfG1rpcSurl8oGxHfCj5dGkbMZaQJQnoaj+R4P
ZPDTQ2n5mepTYGq+TQHReVUJS3jSim1TkHhaHd7CNNyVrsrBqh1sV72ieHjDQF8K
u3fNvPmfMvJBfuC2fffBwZcHKZ7WfleaDfu5AbKHr1Zzm1tkFJdtjwCxGfiM+Tq9
LlUdM5RoAd4GLIl3m117NRuzCt0biiz1/77uR4uZYvQHd3Wyuc54xBO4AT6/n2km
Kf0A5qFj6epZvMCSC5IYkVmb1Ttz98YHGoVX/9c28IDso+PQBBoVWUerhwyOWR/Z
X7zpwB4TdZpgbH85WMh11+JnBWD6qvu7NtO5Wzj9ImMF72CiaC9pj7jZUJNlSzk7
bTTLZrU8cVsz1QTm2BI3MD1+mbZNEzrdOpm5HVJy470W/xLDMi612ME3mmDXPt3H
io87rwAUrvOAXJXPrSInirLIV0UTANVrW7Xkw+n1YC2bPSc+ekQPhypneIKMr2mG
McFU+TUJ71C8AgMLqiUer4UQxKva0dH1gSYglyWo4MFyaBST1RVuxYlHqb8FFV0n
AH/bVuP5IjXF3xuNRjs+JSa5kMrX09Nsfg84G0nF218tsziUTuCQwth9sJIsx2AT
XUEyO2ri3gPyKXD6qz/DPpoL93HDgRAIdvl/6dyPeOH4MEhQDAALVnbqG7s7K+5t
AGe/RJo8cWwhgAgMcqopmzNDFo8+p9qCvJCYwyPD1H/cGCpGjwQRGc1U7Nqf+QFd
Xr7+z+NV7HXoQkFV8XQFLtjzjAULF38NlKPI5LNykHe6KFg7d1yHvRTnwu6hvVmd
fa8RPM2yn78mZWaFdopOklblqIqd2IS7EgBjHd+ev+fkBX6jafCoDCKnUSmc2hSz
06oSQyy2IyynLE8ecn4TiDcbiQqv7UNycmZR2UZYCM05tomffnKOc96Yy3MjYnju
A5dy5MoJ6i4fEVQHpmf0D8w9M/WeRfoY7dycfhooTkIYfpFn/UjMEH1Tb+h7et1B
BE/j2UkIHIjd8iVgRyA7tx282oc6+al/OUwjTwI0z0i8bCgOdDAf6Nx3tXG6BlWS
DJ9m8KHfHCJU2WJUWNcTqjab1cEk+Zu7LXpnbJ8mzx1YLZZvL1ZXmwTr+JQS5FQo
1eyYEuGUzHGLEU0wk3J/ixNc9R62O4MKjz0nntAxE04Hy1vnO80uty2EuAtwJOmh
cPWuMWk9PC/7tNjhyW0olGuCuIiNnj2N8ui44Hmk48eZvHhp5KkUvnzkErNH4JYq
is47Xmj4M2r7c54ySOVcgBljW4ksTXtKaQIM1hhXQ4NOi2YcG7k75IdZZgKLnDBJ
2RItgvo4aRY+Jn6zpd7LIC3MUo6WLtYDU3nuiZKBTEr4nPaasvKJvOOZCqGA7Ulu
3XOIxmjFCh5ur4KSXfl1k0pupQlJlTOS5HtIRs4AzHP1OWQDtWMu08O+ZrJ9422A
VrKay1FlKc2qa3+Bfvkb6kZe6fGPWwN6Tv1mE616bILCkQzSpUcrU46mxjrcN7XB
TxPhv9ZYn/s8TnyB0oVVoP7gvZ4mRzuT/aio61WDzMDs55SGwhiYJmX+W9nRcY4g
gIRxehl9BDa/iYL6YnQrdDXWTo+fxQpktGtuaPHRPbp35Q0xvl0P2hY/shUtnAdi
MFpOX25wP11UGrsMONUxg4+a/FD8gYUl1aKLR4BDVLRmnBbxi2yCOM74NfEwZl1i
ezHTf3UhPvspuITqZQzwaGEbagDRPhTnuIbL+WvZ/xqbKlYCJ9Y8f/Evil6a8LlQ
bFPxt9KbyuXcAcFnPXMQBEgfaFRpTap2ew6WBbfYTtupss+KDhK3iBFz/ACMHMWg
vDRCuY2rljshzxL7+ntW8AFcuqRDMxClRdwlgY4qN8OspVPhakr1UmFG/3TF9UZO
bWr4gKkNko2i9s+4tf8qY62NUNIvLqHe7nBUN2f7amx4QgR0866ze2meYZDRu1bp
pBu+u1MhMyjuSo6lMqIgJx4CvEl14RF9Ln143ljoh8uP8koinlKhu0125BFNp8+g
QtA6rQ6xIe/JA6MQp3gEzXiJkYAqTNi92vPxBnh0aWZOCChYnYbL8rObjzAPij3k
b31k4moRn3zEYzhrABPIuhrdtWIOExdVBNO4iq8NjZ7REJLycrKaifkgN94WZPKN
1TrPDTtVYe50CurFgDJ9LYflV6nwqZF6L9XI8YVbFQDGh8UAaO4QVrIzHkxPFRHO
u2DzM4Ulzfl7YG4eqhH1SDSbu38RYIzqKSBzQ2WMWnB0fghtjZbo5Bb5xVhBAPlb
gTsyaTPCzSYbKgIoURQnMie8ET5c8P6h+0G/vex5HjFRGnhPUPCG7hhhgv7N7NLE
VCA9NNPZq4EzL6xuQvSyv17z/WT1eJ/ZC0jaIyBQahBCmLgzJmczkKEm12/hUeW5
td4Cumscb/NUeLDz6iO5W9dPo0VSj8pG+SmZlApIe7F1qZ6zP5LYy8lZKYvhbm9+
jU06rOPoWktY1aipe/S/q76IRoIeEKqnhraJmsIXW0wt1K28dSukTvnXhQkN/307
sa/o1jKpbyOwce49rzTwZgSol9HQ2GYQapnLh+mf2pp8uXRSs7HMp1UD+Xgbgz8V
a84fjMfvhAv6QHB5tJFhRSpG6dL5SRv72EnkKQdBv0HExZbFpgUS2UQtG6wUC4lv
Y++Jz+fltPU5j5fp6EDvirp8SV2FkW4+2y4A3ulQ40TeIhRyrUlMwTvjdnvMEIf4
Rrc0kCZHPj5bVrwQLtTtBqd2liHZNYBW2Q6Brog4RqZRnDx6qNYQT4b55HQ2NJxE
vmK3vW89cRFJvobMLe13/Sr20UA4wBy4OJ48Shioj2HFSbZaslZLfvJJ4yDM1l0b
ap1dr3w8EsgBEQr5us1XVpfSij019NozuhKy63TW5Z/+MgBSPuwOsze9YJRpUm1W
bGu8AHkOnSGjhW22XYIxZqhReHQ4kghocdaeKav2AGmx6egUPIZSy43OOBtVuMFL
oWe0Prtw08JwAJkMlZyojdjdO/j5Sp9750t6IDFjgkEF/8g3ZfpbsmKyiWrdcW2U
Mtc2NCYDfi8uxabxjcTqIJRjef0RPiTwVigBkLrApnkC+1ucoiWKODnI00FwA9I5
EM1lDJjfRGkdKzNOE4erg5gOas1o+Hsyy1K6VC38QmK8F3kbHMb86iwazEWvkvb8
PgO+Sj/tllvFYCfvHgf4psGXEP+jKrYtsD5ynsulmFf/w++bjjK2XLbiZX+9n/u7
yhYIkcRtXBFkw0QYdMm/9yBooNzr/Yb6c2qCpTWMNgRj5C8E9xnSxlWCeRPvuolm
OZUGlzMV+6JUGrayOhV7enV0LseHQsRFm6DWSBxVU9baIghadooxqVOx0F0SgxF3
RicB981vQpkrOyvRRA+K1W66xynZ0paRn4dOqc1eq7weslVrF1zkmA764XAx/2/s
Xg9YnAAJNG7/y4tVaaOOlqMMPqOz2yvM/+f+W5UL6wzDkrsAXkXv3IVgA8ITzAym
jdo+qKQInI+HatD8CU4p6xmDPO3pCCTLt7lVDJwtexdSwNCsb4xem9Vd77wlF/WE
JkJoWGFG/3QZQmtP3H8v93Grz8Hx6+Gqi6TxyVgZYzlouBCur+UZ9O0II3kPFwED
IliO2kfmFHUA/XjcLSiuN8znT1l/X2CUnY/ks9v4O6tE7jucN/10FJudleZdh90q
4m8yGGQdQw0SyNtJf/f/PeBLgTTRmG2ZoudXVVU+pnntDnxsql0HPjp90fIl4hwj
g/qJ083oQiqC6poWyD+y5Qg2Pqt6zxbBWxpx4QkZTtkkxZ9HmSG+7R5C4MO9PNzr
FzWp+8RxNMowy4bRF4zRe0xa3qAXO920SLsufaZFdlI/Wj4ztsihxmyUOmgvlsT/
lvUn9HUyA5qKHjYfB2EohUKf/sETG5MsaaexG5k+OHA574fPeqEOJgq+be9mkOkv
RG3GWmwVFhUhkJffGI2rG/kF7ipmBh/ClOx2Hde9C4LpCUFlssFAlB9t/nDduP2i
0T7tNwXgquRTjob3WUYJLgociQuJvePFORK0IXPyuDuiUUF62rMjvfkmQYFuN+/d
BtXolLdtADp8A2y26VC8T80VWrmuuoiRICuTzSF1XZ/j3FTEOxeAYHzJ8PluK7Di
ZsUHnsiy0LvblbJurFyrBurfQ4cbCZk1VcC4chdvrV/e2z37fyrXPSYoJTA7yNER
4Am+zJe/IHyKZYpLx/Z+USIZyAW4APMOJ7qU/mFOB7TsCJfp2T2VDfmye2wW5a/+
32Z097KmeLsAq+OUCiBbk7UsIUeXRngwOfD+/WP9fin2rqlFKSkYXSP7fGGHZZja
LLFmpS2Dih+pamSjlaaQKA==
`protect END_PROTECTED
