`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b86KxjRqimue2aD8qiz+xXIfp2PGEAJni2wsvO+bDWavedEZF701tPYK7pvejnaX
648tS/C2y6fHmioq8L7CSsdPiCOfJRL4RgESSOcOU708NtPDgA5HV5/irWEcdpbn
cV7LslHifx1EbGJQ1bBReTBtdHra1K+DtJUlCrk7eBop3dzyr0erKpsTQt0gFloT
6SYIOIEeRfab0HY6tBolo1g5Nslph/WltpJ3J+oTvAgeLAouY6OZJuWc09DeRiYq
lb8NG21NBoX0nVUxdR4EVItUao2eeonxpLtVUgFboHT45xNl4UmpbcXFumMDBfwg
tptd4QRs3nIcOGmTlVqoF+neyuZ/u9oj60XwkKGyXe06mGWWhfEIu9nYh6U/8TQo
8RRC99fEOrI5GyMhoDuRK6/IvLCjbbKduMofbng8A1tr8sE1pP9HtpHPF1p+qn2t
dgyBOr0PZA+djB+QcYSvyebU4G6xMcvR+tYzhTymJRE/YzENnDyBfrB08SNTWDKg
E74ot3Pf0alcBiJlj/80Irwj0wx3q4vDev7lIhwpYUgnJbEjde9OXS5N5reFfr/1
RnM1/bYI4FZkYYT1LxNzNoTXgb+QHfyaQsGj5F62bv3xeB2baUpfl1lyXoPgxuU5
B5tGFa3+UkwLIy6xd9Ni1xFfVOiuQG+fv4rHUwqB0RE1ESSOBxG2Zt7UShLFFD/t
iYmifYB6nrnQbnAo+rbkylMZA64GIYObpmH7GX1vMKEwh9GQMSsF+k5wEHAs/1c/
gGWeppnmqQ1wBh4Ag+tyqDPGKjPfuAb7h1Iwk/BhjzmjFQELNNr7/7AyVf6YhjTa
pRzvWufALLMAp3/uPdjmawks3nvk2t4e/dBg324P0pVzfhLNuS29uFQvQGlja931
lJE58tpuI9X4X1Ya9nBJeQ==
`protect END_PROTECTED
