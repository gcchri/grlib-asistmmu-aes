`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yGEnFr/VZ4U+O1Far9Q82DLyayQDS/kMAYOWRTj/3JgI16uf1oeOzF9YU3rxtZtJ
CZYzHhqtmgRepAEwKN30oHU6N7qd5THVdqU+SfsD4T/85WFJBCr1x+kV0pESAaiz
QM3ApIuT8mBuEBOa6FmfNfJZbr3q+0m4JrJPQNod1asSaHTjuN2fwkchRNDOVgU4
+ZojlY8hpTNLMz5GzszRyvz+yIkz3KT8wmnEZ5k4aZRiBFPR8k51Fx9L+lOtt5G5
VOzFr8/0s0sdetpc3F52iCRXez/rYMclClXsiOyiWFpB6hit8j/2Xqgd0Z/tWAkm
LguAx91iaUw04xTKCOK2ZPp8StwwICUbHZqa1StldxxpVwepYkZh7Th43GuZutQ3
YWs02+eobcHOjFbvCbja3gGyDiU9j1d2TlpwoTpKYM50/OSGkU45aP+BkFW2S0hr
m47B29Blm90YSS5LLnteAlwo6I/Q/9DEHug6REYqjAyorT5DHIFajEOoU1sTeo2k
fcHeJDEpDgjODw4AMDCD9iUNRbCd9yS6f33iHxJwmRuC+NnwbSbC1eaPIcYg1I6y
qa/oGQfJb7LiBFZjKvJ36gDn4iAgQ1y+SsGN3LUnOqhMKTB2WwL4CKO0yDEk3i3f
6ZswlLxuU6VZ5HPW3AQaeJKEn8XBpPZD1ptyWiLi+CpVFL2eww2oqCpE97UAO3Py
M+PR43dv6vLfX8rLsze5vUaHFM3vNB+WaCxl6xt7omMNv3B2ZGH0ZnXITUPjrIIs
yCXtN/ZbZI9RtPvlGEQybwHPOcenUVGn16Q4mTWkvReDXrq7QEEW1DPMC1qWTF3l
DxSmEgco6PeF1gzHJHsFlewEDsStBIOW4m1mjX1Wa9yqdqNqvzdjbIEs9KuAVPTK
yiPCDz7INwld/7HA9vS9BXFgd7Kg4A9eGu1Nz7dWPsMJiXLHuYpmnlYc0Z1SMimL
DwU0JSeHbS9ixRm6UTB+fIsKbOFSvWDsm67ATUr/f50iSDnHgbs/m7RoNNqrXHZQ
lBpXHaEvCu9RVn+8yr1rVgG+zcmGIG24k7SV8v6kZ3DqyOFhSbn+gt0y4ayoqp9g
Ixb0Hf7yfB/972YMOBkB1NqybBIPW4RJ4ykiq++2FvuWHtyhh19X+Pjsa7mtbPnC
rm4mtmqmg3A3QAj8/gpqGhQAuiM/sgfMDerZ/bB578mi97t+SY+xKQAAjTScpeQ0
E/D78kzHeHy/o5LDWpkMQ2gF2zGHfApraUR01DGtZE1mysTstSoT/DGkWiIF7WLd
hr8LxdJsMOYFB0yWghnR+kh4feXmsGg3pFTVKX3W7OvQh7hA1FeaIh1Nppmpo90O
pDmGT8TmUwDiR3lyIgarmjvyufVcN8NYDq+ntGHgeGHAHg26RdqceC5/14hsOYTH
njhaDbfNou8jP1cYOV0rHUisiEfmGj7s6fVW663lQP57USY97JGqTdGpYDgNPm9T
dykM/JNK6caDefCgQnjy0W78Tq0rEjApPsPVbiMv+7HIraEfKlA7dm3RWHThcevd
jNVWr/Z+Y2Xm814rmrO3lKpsxECMJeALQQVBeM0BhpsGhNRLKeCFK2i2AYIhPMY9
0FImnoAW5ZrZCKObBtJFuURUHm9kKgKA0pMRj5voo73IVS+y8dbMxF0begj5lZgE
BWo/4tRGU1NofycYmgRbQsoxJz7IaXKKmEoL1cJtvC1Y5vJ9NFYKM09JHxfroyYb
TkGoVeXmN/niaKTI/lb8Uzae/Oczxi7D/OLFUIjKhq6JFr4UvRhHHc0nwDNreIFN
P/eOZbw4gwcKswvG0pOWsskcGlCmb1IbSJhyHEUgnNWeJwLnQP9ooAH0m+k2DTMf
YpKDydf7cAygx98iSPmVkVEOhuw2zg9Dk8q6wBLAhlz7Yqn710+MwRxOCpbiHtEQ
TC5CyNttX2+fJR3+ON/MdmPpeH1k7iXftNrZmmQqCRwSC+GVyFmG7DOFLmPAcOBi
V2qsSd+dIjE1qq0AkQvwpO/yIW5eiq+cUTG42ARKMZx+98UTgFsxioz+V//ZXxKP
XemcQTYD3vDCqQU5ID/lMb8VVUykEn3JPv5LdINuVxNr0c42PGbXhJ40jWEK7ZCj
0C2o5yV2RNGOvAxtBBx0veau46gNOn5aCz1nZBJx5nq9NP4IVmYMeqzq4/urZ/Pk
bX++8R/AOH/5Vo37ATpUtp1n6s7DbGioHcJ98Xec61k1b8kWeYFPnvu5HGdXJi7M
nPApNbtC4RgSzos3ZTk/ron9TmpD7kbbR20FlYrCWlPKlheUt/5MVwp7CJjhwNYQ
amNP+Gt3ePZ1/PNIhuOgbLl3klTI+Z7LCY/0sC5xKXtcATymqxaBpOhetSdFFYuf
BDzKOX+gDc35vGRLOAutEEXVhdANyFTAt2pP2/m82+yT3X1BREb9JrtGl/eGNoNA
Xzovs26Ja55VV3xc+eWSMfl+gOslv01wuox58Ovo3rLZvS86ziJ6J7RnQlUTFkZx
0K/uDmUBDkDB9WhezeakoONTxAjmIE9cuDf+/Trh1hgd4X7o381+YE3BWAERXvks
lHJzZpK4+V3qdE75+wMRT7uXHxaZ3tB0u3dMntHNRj5veC+VgY87SZr6mco5yY5F
jcZ5JZCBRL0qMftToNPYZwpKMMHLqQVULdywRNIJ0pW6YgtPbanMqj5Zrk8WEqY+
My2TOy6KpyRJn275cBeNj0/0bwxcHxMRwcCgcyQoKFFNStHJIWd1PP7zFqEQqep3
ELX8o2WZOmnqb5ZXafkaBa/f4p7foRWVtKY+kG/kg3eIB7vgU0LSN74IpFXAN8Xy
Z3IPNOjPstVs/QgoyaGgqRlkE5K3DX5tjXXhdv0GaUGLOkevM3+TL0q/YfnsXizj
o+moVNhaM3pTdj7rXyS8S3vY6wRkoHG9iTPQE379+oGn/HZp8UlAHNjaKmAQ04it
k1iBdBhGBbXRlgfyE2ofRJif+RwtFxBfDRrLON8Um71Rzr2ofFH/HE5Z27voQJZK
kZNsd2MoPAWNSZIWj89IXQxx2j8P82f52d5GsLz9Df9uGX7uSwM56QKf4l500msl
6azLFNwpEODF/HeWlccEUKc3i61YsVATFDP4tLuJMqkHh1cdFMn0yQFi/F9Gse9i
fahWug4Qtk9uEPA0RHsuTvfPcG+bWd0SFNTPqCj+y+vjhUQxmifnuYsWPL+V6Tvx
keRmO1rrAlqli0H0aa/+nciM/QlACcfrZWZYL7SAZ0VIZHf5sm1UYl78HDmqZ95J
4/ExT3W6vmWe43l6LWvW1NHCLUcCSRajkhoxJNwOEjx7hJUQNvG1aip2NCsDUqKV
QV43CNhCMjmEJWi5NMFWyomTU18zlsbCyNE1w0PnfQULrlH7S2awcpYLXOPbkXfd
x0Al83/cIJt+XRUj22m7WerpRTbAJs1udKURBApv7B+U7U4a/tRZ7MfFjGEK2PT9
jid0QASJLMo+dpVhHuVC2gQ1edUhRSN4jtbhLBpJli2q4RWI7HfszuljvmY4bjP3
zYaNmtoD/f1Wj3C3HwLq0N29vpN9F3s3LDy5LOWIe3AVp1pPGSsq176gsUseF0ZU
/kKrYYzz1zeQKti2wWNdppzl0hdTK0hfH5aND/FuOOpd5OmJQ2ne51NKm8Ybl+ZM
BXTTRHkUDRy4UklKvD3+/yEHB8VjPkHiUc0l+t+VRUseOTE35YIqU6AoL6JCMQdC
1l7y6kp5cyvYr7Xd/lQ4ydfnT6EyYTHF+nSUCLXx6OTlLJG5G9QwL+rMGecSftzT
yKfZtPr2UCeKr4mgdlDosASIUn9X2riTpqVzur1P52xOBA93/gWyd2Rer8Bs5xLm
EoOinTyWBhlmU+5EthJfe6wK1zuLjx9MmzGw13T0eScZ8DAr8RcjI8F2WPFkd4PO
l59lmGNEkXSZBXIrRfKHf7ZrmYd9xO6E1edaVdjZBK7uRCUDi9CiZtXUY3lpvc8D
f56rF07wP6zLsQHNaDKqo4VOQ0dtb0ZrNGkm1mm22uhg/JYltKL65XrzTfUnBUSC
M1Seu9KgWYBxM70AdaAFZAqiadXb2fuk9fTb48n71pNc8zbrpRWIXGGELQeCxLEF
2ymalbSGTUlC4bI9c43WhVblk2/PSV/cgJfiIHFzrnyeDmZKevs2XFgSyAXj4Dt5
qP/tHaKcqPSK0D5ZSW/GFZl4VB7fxhbNf5nCztMRwhe7DrQp4nGN5+QVOBvj/gPJ
26RiC2IXQ794lQItkyQ3lNayVXlKaKpDaWJN4pgOKUE3EVR3isfBIsGQDtEnefwc
xspiO1JybiAQ2TyJ59GqjyFHIQ60y7D5BF2LQ6OXD9CPt0tSmL0EqVaJ4YICyQPn
52Cfcyl6Fp2Mrn0rWMgUKkTDCtBVNlz4drum99t6NTA71dQfJsF3+UwUB1OGFrhX
Y9A9F8iY4va8Lr6n+4KlYxzd+jFk1LrUOwApdsAsQs/ORWKalroJ5Abi+/Qgfgmb
HbjpGXJ+coH0KmkEkwrDe9rJ7v1kPaoYCZA8T3ROmdgxVrjuzx5ljNP35cJbUYYb
hl52tKSnOQs0Lj4cHIdOpseodhLk++XiKcYTdZOhPy9YnQr41wkAR30aImXPyRZD
kkSqHjwlLskfdEaeBulc6PxioNnaAcAI+3YAtkE817AiJQnfZ1f7em9ims4gVZDr
5Sl9/ql9tht+Y23EdOWVsIOAhD5ChEadmGW7F8jWImnbVAYdR2dT2PP+bWhyl60+
n99jdpTGGj5OGajmDVSm1jOlmWbn7ZBiZ39cQOKQwmWEXVgGxaTCuiPVQhEWQi9U
uQfu1BT4x9OrTYjKwwuaG6m+axMbeSzhgvUXQnlkBm5snYMaHm1HcJi4qJtBVu8b
dX9PlgyBaqAoaJE8KzLBJFlFrrdnWNlXBMYqzjWL9hqa0bed5YfmuFhNJMG+KICi
lgcEbncX9UwVm2RztFoxfkgBvh341fpY/R9/MSGVfN3Qb9LbwtfmdLtMUBV47O38
ezCZfVJ14zj5il+Qh2rvmLuEBSbwRl7GAotAroYcqm9HqX0J5rvWw8COpT+Mnmxo
5Og7KS2GUCI6uHU6n1BkbGF/b/baSlo9RVH4solUUbV5X46EgNgPsbFVhBQYdo15
DD8c48CqTYQqIbeuhnkQO7KvV6NEJ4aB53PCSGS9/DMoJvhKpLmKzWilwpynGMs2
XAywmL3WObpJQuwyXw6Y4uFQn0b/1Ypp1zeIee9lHKFnCwRydP8QKrpKwUcl8wxZ
akEz21BFh+ZRnMGF+Pll4YyvKImn5HVYaOuz07DBlHcLBCJY7bJ/GuYbK8qyA0AQ
`protect END_PROTECTED
