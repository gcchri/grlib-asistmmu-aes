`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jNepWfzBYG/EXn1L7XqwG2E49Pbi7X5mvfIrZKFf4w/Mwl3WKaUbIYltcSxPbAlq
4ohpkbAvkkL8rxg7tN8lBHhIN3KA91NbaKp62KQ/ujc/ssoPz5Z9j7XVKVzIldld
P/+M6dWh2LvGD/ZcOIGL9nsynh0/BaeR0kzm5lBDFnUPwQCymuI8f5OykUHEn6fn
N4SPCohxc0J0ChFRCieOo7OOzePLKz4CpDcKkMvLgIk3POQfH/APwFCpX56aYAQ1
EKdLQhoVVo/+5nIoRZpjigl4Rr4KOESP5X5Wsmyye76EXW6nZbDEkeTver/IGR1g
S/Ve1po9VOLxVLtNWoOz+Is5ADB0GI/u4HnNdC+KVA8/055XC2bP08c1+xQ6pbfm
jf/8a4/UhLSOoFrIGPVXGJR9bnWbFm67VuBrpATeRmvHucKG8UVV0P0HR53JCbj4
kTO6Z8erCfS6bDkoc+9YlMCYR8nqENomElPZZtOQHXpG6iVavyZ8ZWTqqK9zOVnQ
7qR7gBWKjJazyZncCA8Nmv8MpoJ0hBpDrxbnP4ppymOunlYSBXvo+AorvDpeIvZG
wUBiMgHjUC0TQVe4SmPErXJyWnR2cjlQ0Tx+fnz0dtP9lZrg0XSvsQ6mZEkwy2To
W23GLUYWMd1jkZANWHtcnQsBo2nvB+lxs2/3DTlo/ERUef2OhQkIUj94oLz6U6ZN
B/QYeCrUkzXOiM2KFdridBr4lOJCVJf0Kx9WZQtXfkeBGUXi7xy8c0ZxMW371I7c
V23Q7PtVd0+6B5pzrDK75foUZC5ir2aPK61xvJa/rCIEyF9CgPvrWw8dQFpOMLLS
XsNZbo1nahq/qGVPEyeiPmZWT3t4pxRwAccxEbjpctd3knEyOhdOu3vQqmEST33O
EzFKbNuADdS3IqpixnSFwt9FOFHjiClR1vTr9iv9CCUHcAHzMtiymQ/kKchSuG+j
lz2OiXkAlXMym7TdDoZCSxGilaGhRI4CUOeyVuql7mlIQ6aCnQ4HQOlXPH8+a6QS
xPjbLo5vfQ/s+DaSQ70feFeT5PiKCSQt8pvwYvF+nV1i2vOqsxOabtui1DrY5l7s
YoZnSIeD629FCXm/2urlbQn+9OHfZ/Vr70pMtUkebhOKrvwsLxEsvWuy/574BEUX
rg5nBX31SuGEEQS2Q+9ZBbkXD9CK7WzNi2QNsoVIADDJkhAhE1rMrNCnTF2NxWxE
`protect END_PROTECTED
