`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQP1VuhK9VhsNA5MnE+vOQ+Bv9Mn2DpaxnKnkmWvz9foKY7cbDTsAGpLAE/2wsMq
xhnViIdTY0qV21PMqcD6as+nkLWNGEmDiS3xTUTglafKQpr6T/kqRIm5eM9FfBZz
BHOtN9GQJHjqPVk2AgXROPYHhhG1AYFgO1dKAYBo3Wbgr2zrW5Tg8XQt86ZntXiA
LTIYrg652bubygoJ9X6KwVY0fyPRhl299vz5rbMIg/65GABrt6Vl21VGi3Dxpb5c
1yyo8XME3hwABfxHZnkuRjAkuj1SbVwAhYqa8e6xNETS+kFy4reXb+NgablT4VzG
cpucx1Nl6YExduE6f40NpuA7aE24ptobkgog6bJR8WERfq7h5pgOGK5/3gr+iWul
4TGsDGvdzQ++ajwU3Zt4f5TsQBfM8c2JsXTgUPIrIUw4OVjcbkpcOONXNP83xBP4
qvQmwwRu/bfkiAES9kPqmZ/PM/JrG/i6zt1t3T26rI9ZwEK7cbBtIuhE25S4Mp6R
p7mR17/ksDnzOTs2+13j1FhQXa+FwYLCzlmLNx7iNi+nXCRm81YPGj+uu0LyacaX
eSA1vdqTBzWzVLnNALEMB3x9bm0y8EMePgi87jxVIqVqaG6Mj+HAdjtFOWvAyTJe
a+isiqfZl/r3XpauncnhdA==
`protect END_PROTECTED
