`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPaoQr21jryWpeh5X2sRzMGHhXNeFSLwJXlFlikoDS8lRoHQWqhoS9fz/P0FmAmH
DHkP+W6Be6N6BhC5ED43ojeFXIGNnie36JuG3jYjr4wjdUrQMiLz5FHNJwF72Hw8
fVRjwDfdE0uP9U8k/MwIcNaWA7kWXACgEleWhg3RnW32Bk347vcawh0o4FbeUHfQ
XdCrn0icwtWVc7ypFwlSqkCNYrwOcLyjKEED1W7HboM8nhpbNrvrExJA3U7AD/ig
PoJZIfZ4rJiikmJ/yGYqVCGSOXNXeSuwb/vi81kiTHfIQCm+C/chGZvnBKHcg4Zv
92uRdxAeBFUhvHwz+YD8zFYaGRoQMlLDhQc3+eD77WLYqw4+7/gi0eXfY8bJsZE/
rUyBYvlQikYvj/91NgmixdWEN95hkSgzB8DRAZ/XT1ZGJnQTlTAEpnvL2QsLF8zW
v+fY2SJcceRmryIc31bCw7cbeJvApo9ASAyK+j/jnek=
`protect END_PROTECTED
