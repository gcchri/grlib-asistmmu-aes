`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3q5MSd9fW5h0gLJssjam503dZrZR8Oo9/s3yHJbaA5HqLRicchHV/BPEUoG1puRr
ZbmdBmH9ZriWFiAJ2D/H6GcpphG+88XR3U2x4ilPzlcWLZ6ClYYlN5bpEN0bmCHD
+TXW5X5qxoId1aiV7v+dTeIaz8SaEFXc6HHcoiAtsQ00j1U7Fw1wqywWdvdTtsfF
Bb1mQLq+WN1VGg8JHEV6JCno06MCXIwPc/0ID/n9b8At07Am8IpNN7p4ET7Xx16i
9xj8lHK0cptF5qwhFXqVBVWIZo7dlX1jOWSKGsHAXLS0TxZSiIpupc8/xugmEP/v
prEVHEQdP6Fp2C9/i23hRnGcv4OGSmQrcpPb0A6ltm7zMdTumANc9vsbOcauuaoC
`protect END_PROTECTED
