`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4XfneYHyTl9Ay2Go97Q+vWUs9BGIIrFsVfwkosHCo16TttpgWlGK4uxrqWbAnBQX
Kb+xbmusAKhQb5ZItShKCsON9wVpTGi9DqCoF0mNfcpJboVdpDrGjsNg+YVh/zwL
JETry0KcBJYw8cjUmhotlANeOcvbazkTvPqeLPEdIA2qtNQUcetO9pkrsKgBbomX
9sp6nVb3tqeaSEE7oW6CvFNP8CyHXXDVyYCrNMiIwhZuhsiVIO9LKlge9dmNFYbF
lNL8H5F10AwUjvjg3xI1IX4xINNjifmpYUpYU4uOGrx1DvzxJvNpPUehSWl9RWMm
28SWBKml+AZiKifvaVOAoAvgpfPW++t8XVvMfw5+eLoGJ9d8mRQ9KnvFvC9n/XzU
NGOk07j9iEt8wChjrrrM+tGSEmPHBZta2pN4f7c3+q/VEgjqHOQb6I3GF2kHLOXE
Ui+T/YYRh4omsyQmq3T8CKSBXWKuP90uNBBi/VyHfu6gxWEPNLHAJUvfcZ3rWxlg
Ep24RHxvctVwsdTbe6XRuTSd+yaX5IjyK3uXfH/fY5+HxnALXFRmWY89PPsVeksn
LjlaAxTswn0tlWoZTpkEblf9PNRrg/8fEb7V2SFJpIEiyUQAtd/Os9zpQT5HGt6K
o6jDGl8LCpiwbIRTPrRo6cZlAy6bTvS1qgoZ+jFJAUxLjx1Vq0fqqYlWjzJIMupv
eWX0xiB66UMyg8qKB7vUavr03utPtluttVP59wYsGYtV0Z/RTxAGsrvCoyHGaPhF
EJoPb0DGAHQWgznO+DaxEKhsFTe1i4/d+6pTKWNE8QFxYi+Mc8oKr96v9U+8QgON
vtVqrOQ+pYtDpo3E75VtRkha9bzIX3P83gxuSg6jTfuUOWQ2qFtGBfVzr5AcmXh7
vW29rHkcmTNCFxeudzB6qsrpSVa+j57Xp9dDkEcqVcgHLvfXolbIUOPb52iyACKB
49973+HwVnNFpkrlSpdzYmwVZl93Mbgly/0Y/+fV0nYBmmszQMjt4lqVmZofMw7l
0hVnHy/+YDU763DNTVOXZ64wNGp3hivP3048+jzYC9mGhQ4o5chS4CfG4x792Nad
MlRgh+WbQGD9ztNnsxq7wuEiebmzubGUJH7qgqH5esUD8exSMyt1trfEWqQyZwfo
e3fbLueR4WUnuANBN8xBIMGMZoy85NJYlq5mFYIdlrhxcs1pT5ir/DxEGkKubwQZ
2Mu+U5SDyxyUhxbXxLqFI0Zwigyy/6R3MVp8OUhA+IStxbUGsc1YepG+MeGzZyyy
5ITjLh6OHlE7GL1jl36CPxNfoikL1Zxwng8omK6hHrD4650g2Y/lHWCE+TV0MFHa
Aq7Ue5zts33uJpdaYEzgRCDAS3cnwc9kaIPrXUZAHMCJQ0iX62lhb5NOFfHycwpZ
PwGTs3p5nbKFouOMw2hpIZGnb3Tk+qLPRHiEAaLnF7dkzOXbdbRC2CLLnbChTr3q
Rl4YQtrDZDk0xpQog2yyRUDmRw+BcX+mE7cGymQr2XivuPNgxZ3HMrVFVtguv4Sg
E8YzkhN1csvuZwW4dbP/V+w2vxk8+6xfxVC6yVDLWi0PdSK6xL3FSyJqQakA0qF2
eVc1um79hu+cyxo7WTSvv5A9+6nRNyujKKjbMpnHmw33bGCnXVSblT0zXFZJG6U5
GRunheY+Ts1DSlOsiDfHw9HkHKJ6JLEewoPgcz9ECakIQHTl66VgRhGsZi7ieyxR
6X86LQabFY+SCFFI7IVGyyRtF2WJVHFaxVm0rg0sypFDCPvQ4Z6/RoBp9yIVpr3E
XiOJVJT/ikGlUjApzuKbh11C1+n0E/9CRWSHHMF08VkFZqsJibnedXJIDxg62GHy
rJqPBAPg9rWG4VMMIaUTl8vgFq+WKmF6Gb71Va1DNEgKfbi9bO+0/tfbKpEw3xOO
iF5cU9Ab7s4AyWFkWDIzyiLEFJ9vdX6Qm13DPmDg95lQ5iRFZpTlZ8cML78C8qw7
iA6+zwBhSYmzwyPYnd3NFaFv08S7K2Zqdl5JneIocvjID7/e0M/2YRajO9hs5A5q
9u9UXkODN52l8QAHj3+Db+Ek62XZ2iwCfbMGA20jsIE=
`protect END_PROTECTED
