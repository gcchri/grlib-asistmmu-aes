`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISfmFBkzVAmZUD6XYYM0Nz5Bt2T4ftwrFINAMPYbkh6fughmKWr9XFQF7oHjW0Pw
ziwZuK6g9R+D6/i7Ndpih7NUR50XPqBF8r9gi/wfADlnU1ZRsmbBGhaomyv2Osfy
MaykiMiOcXKstNg8VRFmpd0z20OiBcdmnVYx6Fv7cH6RZoWQ7d0sl9AsZ1QwWvT6
7PzwtOSylWusx65xhsRExnbBZ31FCm4TxW/sbr5sTjti7ywwpZro1vFXBiSFHgr9
ruBMTfAtuKYyQBKaJKegvT1TIhE4nuPW5dE4AWD3lfxWSx3QaZHNvzkqO4OsnvgK
NxA7PdZ3T+Bwpe8dSmSZ1GshSrkoW0jsAInst7swsrphzIBc+mwpiBO3WEduqtuA
/NQybPpvKBGNFlw5rvtRMrvSKV8RBQhMQBesc0vwWxvpKRu+PS+eWVO+jTwK6Cas
AyJIvfDPdMQaDhWeqPJzxiw2EAncHr5ihkPaiMPAQV4LdaUBmMD8ElqjHG+Oq61d
y+9jMoC/sd9+ep6/5qxMUaDi4OU8CBd6zAB9mqLsyGzoslVfTOmjbBqjfofgBTj9
2CvAxY7E77R6ny4Hw3jOeaEo8YupUWKYQ22RV1NSgdBjartlHZEEGE6Hy1OuCM9/
xMIlyfc+GXxtB2aB+C7wbG9lIXw057xJfohPnUnOjoRd9IRvrqhFpHYOVH5BlCgw
75wds7nqRaJH4I2WuYJNB1I6W9/5K2Z+jWjlQ39FcDg1CkjaqdDjvpl2xJDQea2P
CLHRgtcz4SuI6cP5R75K5rZcsaiIyhbTJ5n8vXWlRz9THpW5kxC02zwzrwj/lB0u
M4wKOBGJlYobaPwPP2qP4dfQacHHGuQIFTfgpfTAIoB+sHEQKKhxlfYd8BlbfnS1
yVQpUh33YHgr4dkoX19stbcx5CWeCqxKn3vy+FYPvRnghCe/ga+uKbdijiLXid3E
ZM8WUsh9mf32KuPpF31Sxnu2FW2QjtO4Z/wHJ/JT2o0XQFHoI5y3/lmSZ+w1yTBw
sH3CwVFTviCacvLmaLOubhgvwgJdcHI4yDbDyZcpgGhmYEpm0OrJUO7+xZ8U4hcE
c5LnH9ePdzeGSVBpWS7P6UYOcqM/tCXERXvbjYL9eTmfi7oaFAXAB2JRsdZFJnYY
bwA+ENcCBE3rZxwBB36fZgZdPZkZJLwrVEKZ1Z+5R6zMCYOUQDUcdyJC2ee+XD4F
K8XRnrWe+jsvo2EceBto6NPcgv8OAFgbn1ZH+WI7Kcmu0OJdJzZSa+UDF0TbjC/X
7lsq7yu0owZONKB8eC9kng+t/+wrAq15nL9Z+jmB3KFgoHe+oZAVGNdzjjhFCW5Z
l48lw7zg6vZTvjYzU3LXmJkaPla9lSpiq0jKqZzzdVlt2D+0/bd+nwNIu0J8TlPm
/llX1SOzMzHMKRFr0sHOSqL/4xya+vOSzRjOOgAw/g9pLRtJjGxtxTxhYOJ6quaB
rAsRJdnla8Dtxo7Ld4bYlUr/zjs5lMUTN2MQIlj7Q6l5mqsnkM+Y7wm/95VyDEE4
aGTWqGuESsMsSFRbXm64OyeDHPHSXjX9yLN3/leJliyRk1PsCsIn3j8d17blM5WV
8EXNx7OLGw2SOI1Mu8n1oX+YEK+pHjqo2QMvSzNF/FsB6XYzuCx32YnoHDOfHxU3
tmlcFiwJ4sdZFTt22zz8NDoTJqyDwP9s4UmGAZa5j+YdA3zDLZ6tyvAwonzM4lXG
G3j0QN5H1yZU3Av0C0Q0xMRFIPxCqn9g/GAMpe3iQ/bSqNwXrwzN0rxoHQP/BM0m
9aoPElzCDwou1rbgd6SCK5jTuG1RGug6lHiv3WXg62hUIpk0IeE31KaZVxnbDzby
0QoDLVmDw4dLZ1YsGPnb+A6qehh00eW8vB9GnxBTTJooZR24yKxA+ehE3b8yfbWd
8e+CytCmtCsMVfSx122NU9oM65FdJSviDBtFRMNb9xiKca/TX3DlasGti9yzXpSM
9FMiUTkkBzl/ZSAMoK7ZZJVMRYrxx5qraOg20GLoSlAbVJkdyGPKo34LT/eEuXW9
zxSAvoOWX13iLpTOGCUDWH6ZGpCvkHGWttuD54twVHTDELQr7rOW/h4CCV8wpTIc
bUJGhp8km+dcxq5pxpX5b5l0cPrlSPdVraAEd/LO+B796qjA2sdGfurkh1gvublh
WNMSYvReBLjw2b2O5p01/68QuJzSVmfp+2bwrkxFoyyVCDRc6BDYUQ4zouDW17qi
avAEuFzbsdkO8qw+axQCJC0B2YIjfydweKtAqBOoV/x8RasO7zmtK02a0AWPfyaA
3Mm2Iokn5a2GaTkrw4eLxygD5dAOCN1369URjwYHubleanRIDJPT5nBKvQgDIsSk
/cMGHly/cwiSpkGRyWYOXNy+HQ/zuIGTAQUe4MdObbRhK7RNIPvElid7cI+JL3L2
xYREeOYcF7yXgrNFWHZpmv3OXpe9vmOWQZwi3p/Brt0a7nvS9Vx/ZPXnhmOQjIa8
2OegsQWrhxqdusSH/XV0SSE+d/D0wgou0V9Dp9tsTZI3phPmKskQHVIGrN91VqZW
hiXWXLXeTRJqBjN1Of82mefIKtKxEfY+GkR6a9YhBn5Fn2vB8UTV0iSGzQ+BaIYH
/vIwwhshcnnqIfgcQhaTWFCZ0mfgULaDpJcPA+ivgAAvtkQ4hKBtJ8C5aMvTTvHX
YVGjATo0eQzjQXfHuuWov5EKZnPvy4ALPK7wAlOmwCDekJ75/SnwWTt+YjznooHF
/9rln+fSXbLgzaX0ZnS1AHM1b+bKMxO4XJuTygWQ7d9Zq1ZJLzyIri6qf84ZtVVG
2q6UTzvpdJZKoNdN67g4/TpTpYwZDKmJRnqbAiJ3dydodqTbC/mnnENphUvx9/2Z
ioCT/s5rnB3qi5ep4mbwfpkj7xUEPyNUKOO1U4grhqzS3vhBJxwBW1o1OTC22tNR
JkXT9TYL7RLgu5LTg1GkI++wgHGqWMAaqx5OTF0oR+qXkaUYCLoKOfW/yEvazWac
79X1Bi33z1s+Ok+nLVnu73lTNuO+xBM799BFxp8uHf6Yxd6CFUiBpeMKxZt0aJ9Q
JY1mYPkXnc3BSien2LzIFs1sen1HnhBGaCEGV6fWOpyFE0qKqjNc6KPWxSRQGg1b
2UaFpIYq5xoghm7/xJznk5G8kApsRjAd9zUxjmZSeexD3QVwgWaLQS/QuxrxYEvS
PZm3sI0apcUZoaSn3v9JocqZL512gSKC+g9jrGoKZJIMgGWeYvLw78IJDILEjRvV
LGpZTXo27TEbbvmLt8hLw4LijPlxt5L3yHPIatoGAmITO8KGKPGaYxKauP8Qn7Lo
N8mP9YlAiB0AXA1yG4iwY3OFkVdkVZTp3qe+T0nm3I+cG3kkzOXyicS4SufC1/rj
Cx6hSD8dvbbiSeJGHe/Yh8p/SDSBRnR3qmybFL58DdtfpQt5pzYnz64idEGMTtOa
lGCdcvtC/7IZmCNvGU2D0Octtg+g0jFOsMO64lcktnCLfSsj2MdRLsd16m//cXrl
z2zdxuMB3xwU9SGZcAZCzVFijylV5mrbEBcycEH8PUziURmFUj0MjIu6eppcFFej
UMQ/geYK+0PuAoj4gxpzqYKmKK+lUK0JGAuXHqUH5IwnIPCCGuvwAuwZJjeEFcAA
AwshSmO7f3rprzaA87TkRCHfAEnROMirbsD1SiaKIoU=
`protect END_PROTECTED
