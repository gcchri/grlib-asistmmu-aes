`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A1Ew630OTXErih4MKWB9HSzgIx34LvU0/AVxvKdj5EAbxSDPhV7zjEVrpGa4pGPv
T3CsRIT8e4iA+m5cjYZ2MHV1gMIvp59veeq+arCzhKNyxzGg0EcS3qZSGJWHSZRq
d/wmMp+IRCDMVZEWLM60T83YewMlPhSYEFeHX7jtZlxiZu9IdFRVGWI0HP64Fg7A
hSRvRFdA34gn2dNgKIMvCQMLRMFvf/PgHT2BQD+EPmW1qQXWr9gs9P96a9L6hMqt
EGGW+WMjyRR2pZKLZIu96mB9J3O05JGEaMBma1k2GA9/hVxS3arosmO0vTH1/Du0
RofF98O/uv33MM53Z4MXPajUV0TfuZtdeSOsYyRDeje0QOx9GgPxKqfaVQi1WH2E
Xu4KiijAeQ0tPIqFkWd1g1b8MLcEtHcV7/QVA1zBfXY0v8yCE+GmdKbXngKIi1Gv
y496oM3GP1XDcSvVFNmf1+5rDWJiBk09b4VPJeqwWiiAMJjoH8RrKSPadT3+3Rix
it/swGU25bTVMd4WYF3SoeMbmZzK5E5y3cQqPrCz3Q9fFTODTia56YdUYHm3xvpS
5M+Adg0/e4ggUo/LCiOwqQ==
`protect END_PROTECTED
