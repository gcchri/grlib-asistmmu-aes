`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Yl0eXQUAbavmB9TADfpR/H9GYxQd8zzpKi352h/DF1BXb4ZFZIYxN3avq0Ux7Rb
xQiiUedPjfz80Iwi9zHqBkmhYZ5IvESEte/VSgcusLi7TM8pQ8F2c2yiHPaJTo8w
eiymxmCX8OYJ34orkHy1+VatzLYThBobVbd1fXY3NBI2FAvKhQ+5K3yh558DA38Q
1mjdURgAlwmdh+fqG4cmlpP2rfB0sMBlhwhcYD7Eb6SzFS6pNd2FIwflY2N9XmYz
Y7VPZWr604wCy6UyYqINi5vIFG7oowIxSGP8JTTEqdRUYAXi9fkf4lWjQOe7n43d
`protect END_PROTECTED
