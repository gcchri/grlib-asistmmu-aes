`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H7wvmOITCOooXRr6oUOA8bcUWWTfmIXlpfVoC7OY928aTVv/fIhxkgl4mUd6SH9q
VS+Dw6YNlQCNEslYESWcLqJSI0i+CYzDWyeuH2x6JrY+y4A7Bv5mzgmRoUBbnm/b
pcaYjpyqBzpAAPt7+NXHSWiZb5YyAT69LdaBcXagL5YtIkmidJ+G41tzucB99DPo
QP6V90ReBeCEHifhG/trYBdN33Cp7bOacjyyiIdqtoaaWnkTPD0ZP6uDjoZ7h76Z
p1nYhYa+MyExBvAon0g4cCeiMNkSfarCo86ALONRKuCthrT3SwVrv8Ahga+sXlmL
KPSx8KnP7PBjBhAZV3eRQVWQhz0BYpZOojeGuZQ1m0oV+AgNiecsV8Z5kuAk02KC
FnmJkjgSriKL1jZ6BnWPP0SB88EypLONZYijpaP0QhY=
`protect END_PROTECTED
