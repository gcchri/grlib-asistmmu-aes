`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/hk+eym8Zy4zDsPenmL2yMF39F9O0GPftQ48l05VKLfZMuoAhZ/30rnIvML4bUG
QlZUnF66StIUpLOavOiIu+WiYX8HjxKKYYHcN+fOH4kH33RVBK/G+C4y/EpHYrsU
RzCPxFj7PmUeCOBynIhQAhPILQKYvtukb9Aa1KL5gGdObxFtc6ELPoUZNSka9xSd
3sB0gE0BqHj9QLr4JDS1q7RPmQx2HjVF1yrSVfBLhYyqh974ayaqdR02jbW26fLS
8sR+Z4P8go4NWWGp3nPCBqLJgxTfpw9EwThvXeIktTuSAz2uc0g/sqMEYhWU8Xmb
AglPalMEOKN7UrV8Mu8ubhu4MyHb4ps6TOHYUdSSXh83VzVq8kawBw5QTXFXEW4r
Txi4YnlBad0IotE6IkG8cLv7AHwUcg3rAC2sccFg+sj8FIFSxTc+abvt0Rjrtj/u
`protect END_PROTECTED
