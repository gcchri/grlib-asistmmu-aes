`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DgNCuWcQowofQ5vcfwN3kOwXEEDfokEdDdW3bTFE66mIj3YHJjokb2p3Ek02HbYg
1K4Omgy8EjHyvlwOI+Vbvm2whofEDOz1peyv4yVQXgcR5WuYq2jqhmXgpAkSFDN9
BN+GUqzclsNepY9XP8NHarPHtY3ho986Qc1lVISX1qnaZobQJ9NMT9w2+AXYw4nV
7gTxaf1U++MhlIbST3qMvrVk393RPoexwuGVtIatkqElk92RNTB1d2SSiqtfitVC
uAARaGVhKn/dt60YxFEt+2MCpziACwTAxzvo9D0JqPC3q8lv9TrtL3b7COdnTwAY
oxdhLSd8IxYuGBRl4LXCRqrBq/xDbjlvrqUVqLjLrqMpW9sbX3gKsl7mesiUGyUX
dBb6CwdOY9owSO3dpnp/VN+FWTOeA6DWNNcOjXEQ4X5VLOzwWLV+xEAfIB5KdUji
oYVsXR802PuRWLDGhM0gZVr3ULwQ1LqD8KkrwlYPT9xP2AuFCOOdwUrLHSWyar1a
DvgvYs0ZmzPwIxft07QsUUFV13GgV9OaP1igxTSQlN8MF/vtSWJw7oIEl3S7Win7
1aaFqQbw4m1F+xOjIicOYD6ueb9Mb3UbmBInVb0hJQ9oRs8pLqIgsW1Syd26LyLW
vSfmkiJsxwx/nPgyWKZ0UL+HArzS0ZUcevGKEFQxOK5inx8WtjK12FArf3FcXKoI
EbPreCl+2cwa2MhmdLIWxLwsIm+/EN6D2bken6UTODnFHeDUUGYPRK+DCUoSYmoK
v4z3nkWhFe1VZSr3AfkLA3hReIvW1sqkcilEX4eqAZ9N5Cbu+SuxpQ+4xUEPFdN6
OpRtZN1FZFgFTNYy32GE5BxV31sGP23hDNPGNlHOQbMTQ2aNh+aAk07e46efUDhK
X/TWafJj0MuhEDAhN5IdqlwTpkI4iicV1efNE+zWWo2+oAT+YA+ketIU/ZzXo85D
kj/0xuwyEEihOwSVVrm6jVzNUgZ77NRcHDZ12urNTkQPyv2x9m/bVuT6hRmkewDd
f/JmglVLlpUDlIMSi1bavAr0ypgI7BkRIy1gKYrkfKhqRZ6aKfZKjiSEQOnyWpXL
S9cLBgiM/bHw6syGL1noiQ==
`protect END_PROTECTED
