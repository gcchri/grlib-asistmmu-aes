`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p5pdpbWDdzkCI4KnaGW5M+ADrqfTQ11ANefXRdH6BFvqoX90xLApIhd9BF9oIvSc
bFgay+ceZf4EKWcEbdO44x2TB2pJQeSpwllDv2uemoJ4qKVCL60bgbQvzyRZryAr
qZAH22WWEDcolaxKcZNIcoaTeRMIRltjPCxlNtFvkZAXoroknm01AmsVGwvvC0+X
EdJZgboAHNEYOkj9z3ZlHIsQTE678akbwMDL7I1v6GwG17pH5q1wT3e2BzYSBoRh
uq7E+tarQfLvcg+hFK3uji1e62+kI7kAGw3KN3bmv6ppPhNnPe+TFV82KuXRG3LN
`protect END_PROTECTED
