`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+6X2uKJKdUh84ofGQjKhonmRRN9dzE5tP9XsZX69Uts4skT4Zjo3qXE8twHAv666
8OJkq7hismlymhdOe0MmBjJOhKMgxlQrgdz7VRjrW3uSyPISuhh054iwZGDdZYL/
o6xa0ktuNwtoyvlicuJcVX5S9SIxrHO5BDsIoj4BiS60PfEblXlc/up8NjEbWqaA
HU5krMMIhdoxS+AylRLgV1AMAVGdwC4AsGoOXSRgr8ENKpr7S716VSVMeBQX1Aud
l+E+GIDYXGN+aUsTEVz7AG6GeXcI79kI3ohy8s2zpTvT8mRgEl/WYmJiv0JbfVwc
HzxkndotKz9UA2KKfa4MtG5L8f7Wsi5getS08+7PLxc6B6J/8o6DpaZ4kgvZ0/Y8
kFlXDVwtfcWvq8+ut9hAw0el0JZWbLBVwa1IIM2sJd0=
`protect END_PROTECTED
