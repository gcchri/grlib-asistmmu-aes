`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WeKvooB98e5AY79XJHgrHc8iIgxyDmM5E7nAyRLpmdtzb2vVt4Ulebyv62XINyYV
+NA+UZuXDtYAGewTIfKfWpH4l2nhYOQ8yRHxzlJ0urD/t+GM+K5D5yzyrrsxDrYv
767E+7/2J/n+GIINdGPs3LHkZHzLOBZhnvRiOuiYORw88vm7bQHXG3CBvtbGoZuZ
OJkS5mmXcbV+y+ronUV6uER6vsVizqjFBDJhl9q2qUKsNJb6c0IUMvaxRf36cqHh
mYfh6iY+AKuES1NZSasG76B82TkM9tbzxf784uq71iN8F3dzi/Xu1U9PCKw9U1sO
P2gjwiqCjMPcG2zFZbdEdh7hwonWtBQkK4xBoW1azBUi0q3CLy5FCLpJ2/DZhJyO
aKd6cdYs/zrAzE7hLAbBA6jfnmg5uAs/XerqOEPBDHBpj0GH7GGHQJOl3G5vM4pe
zkii54wcVF3247tGmUH2HLE0bKp3OKr/kfFVlS0zhXimjZHgVuXHuUpLJ0BCvOhY
GTZeaptOMZErk4fJCCw7BA==
`protect END_PROTECTED
