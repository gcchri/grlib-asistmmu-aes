`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MrrMGVyD5yoCKPCZ6+ZGfBjknfU8SQ5d1kMs5y8nOVcO1pjJuGlWp2hnFxsKCY0b
99ygBtDGjFTEbLyWqrR8boeKm4e+Q8ldGjd7kIDxF9FmqRk1jwx8yFrdW2+gMN69
y94dZM3Kw57QddCNRGu0SGM88P4A+Hc8z9UfXspYLBgUEQjiVRzSHYrabZnG5HIK
FNHj/D/3ENHjdeKHRbsRc52Wir3aeOYetNLxy52f0bcRX5NSDkWMc18kJe59/xwF
azaMFsob9wtfQ2Ftp+VPnuUypKmwhmK4xrr1gfmYRa+/b/mcVtbYRLP0y9IiOw4C
cZf6VwPYP0fGy+eIH7QclnyAmoELSQnpIHdDt2Y4WIYCpkQWMzESqhUo/SN8xthK
`protect END_PROTECTED
