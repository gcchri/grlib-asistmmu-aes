`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkTQXoj97szrME/hJMMp0ZhEKybE+FA5hRTKbj8m/C2qx6vFxobPXg1odOXmWA/i
QWabix/ED4X4ii34UY39Wc1r3EdXWWMDBnd5CqcjmUNzG1A2dh6a9G1n28BkFMQI
bYNefYpW7vT2nIJetuMN1b0RAx1OKcPxV6UaiGngCNrdF4mWprHM09OqfpciWCwk
pckgjnSYdsKdTVsD2Ed/G95y2BLo7UX2WerQVPGqhUqQg7SKgY6AYTi/X1qFFTmW
AQ7Tb1eQZDzWlsz0hJdhL+lNsilpgtxHixkJK6q52GhQQP3f7rYgEhM0O5zZ/FSl
o3TFG30cJQUv2gwhFmJQ+9uixaEzU2ZUHgorAPAgv6Zm8TjnB5RFTp5JG+uXL3cE
6Ic+dLV4bdplMTgS8wWeoA==
`protect END_PROTECTED
