`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7smQ9BReUHaS+yXk8P0FJ1hGyE3s6/SOTW0J/0SX8GZDgjUjoI1T2TIV5rno2ON/
OPWewID9pHO4p98XYtL9Dk5WXiZIhf4YkH/BDsAKI7kcorYEIwO0yFOjLJeYVzXr
OiZndovYvXg+A2Q0a0gj/u2+0ap0Li7kTRmuhWGn08Vfg1m2cjS/NeopFa+FE+aR
qjXdsQylfnKpgvB5gzdojA0pGKduK6yypqEW5dN59xD/dDewhgCJnliyoY3CFQAK
diAl4ORSaYf4dU+14oXd48Pw/dv1kDciKwk5QmGSnOAJzwEm9owC4r+4yfhhnZWw
jzArosKVB7zFrrZzelkJ/A==
`protect END_PROTECTED
