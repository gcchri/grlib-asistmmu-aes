`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xePQxU3fYaqCag2/P5mCSuHZcEt3wqhviKYux7QfLAHtAoa+s9h+oDKU9p0ClKEP
Ke2akFVnAztlfaiRJ93FUxevRlKUcqYMZdO76IUduLu7lcKG5ItHnW2lf0mX17y2
wh6oOHY06c9UtYtHWuZ62JcsLLhBC64IYq7HHDeJoE2+Kp137mjV4bXLZ8T5iMm8
VoWVS4zFxScHfRAa3hyQNdRAjhQbf+ORFjBlHbm1S0+UjuRrseGo1iEkdK2mS+0f
RSFv71ala1gV6maot8QWV/g5x+rD/cAyUrqxOIvt3yQLzTflxw7iogia5DCUM0bM
BDDnBRrVWKndIB+TVwIizfAZ52LvtAFLNfToETMAZQUEXHCVekRYZeeIK3B1d7+l
zj50V/sONsD3g2CzZ25REz2l6DUVu+ZIEzxZUsv7Ndbfdq2+tNVMw1EqurHld0cq
iJiMaOPnwTR2z7LXfbwVoiKCoyIqhbQg1cOZsEw9d6fYt3FBSLvgRaJ8dxyghVZM
hbIfFqgLTCSto9hcfmda5pB2J+Ucz+LOUOg51pcQjzLVKn3/wEj41RHaLUwWKOoL
CMd4HZ6YiHpdEs1v/gVGAtUu7tyeIw4xDGQDgIClzTqRA2YcVfJgNk90/TbPbmw7
Hb9En00BK7iJZGcr7s/pw29hd/umVo+b+pd6xll6HklfU6P16i4MwmCmX6FCu9x0
uMEh4QoV9TluLdGbz+5Z7xjAqIRUgfT4XQdNokgLPWzuXflLoxX+pA7rdM9qi5A+
CnmzO8PcEyePb++6V+9in/vhLTK79O1l1kN5GWqfJ6stBPII/nAYqnosc/rY/IdL
XskyJOmcFkzwLDp/pAxaua4cqO2Da7m3B88PxHaLu9AXT3xSiObKZT8/WSEuSOPD
hT2JtmyftYGKkkNqwH7q3dyr84ZmqCOlDec4ObZRzehA39pBOY6U0BQDgBATCMbk
W30WCdJ1dQVG0Zst9ptz1r6AzZxKh5CncVxcMMFiWZVnfy2+aPVCWmiPaOuI13oj
Xm2/glhoDi+/smDBhnD+dUA+Sv95WbblyG1mMLClmhoqiPwDB+gy1fqEfKNlZIU6
ISQmWSb5uyG99Y7IDiPzIW6kNAKTN1r73Xomhz627QtY1QNcfQMy5bGEUidJJQ7Z
H+ZzlcVxZjQpigRhaaUF7jikNBoVGJD6SpTbelVtic15+WtQjikYHGoupHM361PD
ud761s1YfcnHA3sqgn5nLc/6jjCJkF9QHJ7Zk+CIRFvlvu8VMVNemgUeZpSB3IcD
2RcVTU+3+xPp+IZsg3Dr1GUQi/CCa+Jr/u3TTkAxzokySYo14uxOXLbqu+lDr2f9
Ax1j1iRhv95sMf5TbOURlKY34RZkai1SXb37fCaxkv/DIjWehEgTA5QWWmne42hk
dw255zzMe9cPVHHc3aYZ8FZffuCTbbE7fnpYllXT51Nqn6FHZeX2o5Vz9SP45t2g
/u0RcnHQjKn0utiQdRoBA8r9/kxI2kjz72hhy6EBYUZAUyYxaATLKXPXjO0+Eubi
T3EpHVvA557Vw4Ye+ciExoD4LxZw0dflbMg4Tr5wlYmQMOSrdhktrgdfQP+bEIml
I6ipHmwKsWe1U+suXI/wrCirwMTFlUUmu9siRvnKLs8B9qRDTUS6wF9zc0FVFKUA
80J/aUOI7vBPmZP3Ln/ha6pe6Beto34hXxIlpkBBdoP8ip2ee36AP9Qzcd89DqHI
wxMjgD1vzZTsXp+XhNFlyVvOFUn5Ladl6akaLFA/x0lo2xNdqj2ay/6MHQ4/36MQ
dNuFgDRl65VRZyUuLT9O//pb+p2+GRz7RlRPNgCyTnJffmAb76pMjMvmY7xeik9G
zLxaC7FOCuYzH9YTdiWM8oW6UyL4oq6Bb6jfgQSEcniRzA/Oh1wmHlbrkOvLODkp
Mu0WL1SPuE7U/PojIrcuYJYMWtqZhSyeZCPhNopQ9jqSzTEhcq3xdgudiViJC+8Y
vu/2oWOB6H1LC/rbvVbXAHBkqGJn1VwyCekiwKgkLhbxJXtmyArA377wwZrUZxYC
Q97jHr7XECiILxZHjFVifuHwHgsSD4fiWW3j5kIL/JmImHP/58pNRoI5B6LymJwQ
oTvpxQF4O/aNlRiojRoC6xoag0B2LnsHOGjNDHtGVk31H6YfukfTxym72elKY616
AS+j9bn7EK548H3lWZJWSrdZXYiIXcm/Vsiig+HY64iAroXuZsCo17PMC+9BCMwj
AWYQhMW+94RNIkCigllSPROQ9K47qf40m/KuQVeuCrUWmU4O573VAagE3mMOHIM6
6hJXId4SAvwYgE1C/IldNiY4o6NoN+NqfDHVHc9N8s9IUuqrkxg1eZGa3pqqwn7v
2L+myRoXoCYUB4ZH2lqM2XjOz2cs2iI4gZSx8ovGnpcJeI+rSvxxMHjSI2XnF/nb
fwHz8UzMUB40ZWqpAnunjdufXgP06cJPaz2kDTs3nv+iuCFG+DWm7cXKn6hpQvWy
r+gdR+cycQe7G3OqCdGIC4Cu+tOF64TcuCO39uUChDuvTTw1NUx930U3xQpdBhOu
+y0UNCr9dNH9c3qdOHp5baGUxGoSboULVjHe8kjdyvTYW9b5cCDpXeiL2a8J10Nv
nj7t9TyD6CqQ0fdVbiNX5PIPl3cxISn2MltZ15dNpcfF5Bui97XeTU2YWAW/Cu+Z
HbdIxJjTL0JJCUp75do/X4R0TCGOySbFFKRPM6meDCbx7PNtBYOQw0bcXMNJitLK
vWaovAVz4gDmUczKj/vL3xMf9JZ3fG+LJdKFkj1bAL8u6G+8AdR+QCKTpyeR0T03
pnJeoXKYMDHVi3y/RqZrC8hKVa7KhA7ctYeQvmBXI65IoKWJCQVeY7yurftrP9Mp
CJo/6Aioa4fhonD2Qxu4P/1a3lBD5tvJJXHgOYXLL02az70tb9CjF9PF9Fm906dO
KxOnRj3aOgYEtBGvt8IRrs/gA7yzRfzloZuoVnktiQSsAC7+mYOn2Fi6CLr7urF/
C4vQOMgxYG4kmuH53jLT+1skkNvEp9zwNrysz09MiIBgJORoSbRMWpStcS++NwH2
EtT5A/vTyDt99MvzPchzVCkiAG8/LYv8ZbT6v1J6DO0ke7H23tACZPR43hJuYU5Q
hQIU1GwtLF+OG+LvUU1lnMoEFs8H8i3dgh+KQoGreahXe3THkOO3D88rPVvy6Opa
gu+zf91qv3PSi3gnk+ikCUJ5AaV3y2/VH5EtAJC6ztK3P+mbIBEPUTEZltxFV/MZ
QBQ87ORNtK1T2tPKWnBk33uC7grA0LFnkn9QgciHL0uzd67vJ71s23nuKEmQ0YoL
WEEy2Rd2j7IwNf7q/GkHBFfrgjbs3J7efed2bG2dlRtuRSbIRs7L61ci38PNerSR
+JXW3ilNZZD+GxOmqV5c0pGULojxweYy0voS51EvKI3PwCbGFZwuWt+7ph9UQep7
eK7MZqMfVLB8IrCpA3EpukZuhmGE0suR8TWlBHpIyxEUxijfeOBH+uk2jjKnI26j
1E0BYDJf4om/2zgUSQSd72pfEuVmEzNzmRBrd8hIhV/xz7us7Be5OvzxsWWHWiXQ
h9xZwTyEZC6VdacJBwTQyDt9mp4A9NYjDlermMkct1zTuBfBMkgcaD9iF0NLGN2v
j+3PBQefHyFXASoxhLO2i7AMshE6KyLjlyRbL6VIrhiJfpaDzcrudoqveQ40/szP
6JB3fVRdGysuOhtJpEzi1Qzv8Mv+saceheu0YsxuxnOCo4Nnsa8draoNcbdm7Ff7
1ObeO2HtnUjaPTI1oI6wqF9uNMYGhwaIhP5bmBlbEOW+HFSdTICDdPXnTOgzJMlA
Z041lQmO7Lhr+EQf282tRjJFxy8u2hxMLwoWEr1qMtPYvdu7K72PFdbmKZnS+gZL
k3pimM0tCLUZe54hc7h7icbjJmpx3Hxtyxm3b/Nn1hsZEfqs1CSNpo5NcXvtvJMb
jmKKLnKitZ7ipoeBfOjtF3AdlhoGrvygoFLibuV8C7KIOyxiH9eWIyE7NJVZ29wi
UiuXyWfD4aPIXeQV/xdwC+z/xxe2oEWdTjQbhGi2HcnGo/lHChHYfBiCPGBp9i2H
kTt/Q8oO6Sha7nl+UpIIl2Sp2AW4Xt5YpMqWB0dzN0P9kq/iBKyRXN2Qxn9+xeV9
+rFjFmbuQCb7BoGbBEb1bAcpK2PRf/E1nAu3MkrOK+FPaO5LAHoJXz9vuEF5QbtB
vE4KLgQon5wN/csTP5oV7+j2EMaMBLC64MmKpeulotU9oZBmV7pBNI14xtG5jgb+
/sO73XzcVi5xWfrf7bLG8w6zFebIZevCLKLwX83dqizahhqAWRnxO5rEPW0576re
RysQJs4WOCAtKM+sdx9A8uwL68xRvjU6UhHnCqyNuOBj1h9O3SEGNLeb5C7EIpGj
+eaWx0pG+dnB8O2JllkD7rwi0EsqEDwrru5CNrWb7ItWa99P3Fv1IW3CQF8DuBRj
FeblcHuM7XzAoCw96lE4+FYv4qVuSFuqICeBDU4tDeCZHQU6tc3AomV21KCCtbRg
EQmXW5ik4/8K/6Ch3uD+FUlnLZsxA8E+v+MEKWvh5omUjq6O9rLRJIb4zf5BAPJm
x6b+awyKFYkYRxRREeFmGjXFXlpXEiJUQk0nzTj1zneoUDqok1B+n0gRR6Brhmbv
cA3AuEfK4dNbAMFIIqHYqgzANF5H+eYym2H2GlaEmDOm7nGnAI87mQkCQObg43T2
NlZBvgeoYbi9uTkvo4QSreJc4u5NbddCmbVoyVr7wM7PQW4owv78VERiKN+Mnk3u
nFnNTyuvIJEgWoM5u+AJxIibQ4NNsIp2A1gDSHL84gn13iTBIVmWc07+5G08FwTs
KcLJlZYzvZja01kMi/EqAOZ0sDWMlJseea4mjiwkBIxLk9sFhbQwuavy9fj2exA9
tuD8EMAC/wPdTwVZRV48LanOOegvNKylVY1D/Q6HS/VbLSWi/+bb/Gbkw36Whj8v
3yFJGZ66bXjwISeYUVRToxVEg8za0f4WGKi5FGGBcSiZeXW5TQlh7At4peYi/aI6
lS+XAcFiAMtObVMhfypQZM/2XMttgmKyLkoWeM8wj+nDav5RpA2IG1DhiXkY6RrI
5nAFSgLyXSxOpq2qMwc3aB2qlF1+oQDDuyB1splHKPom8INOyT/rNdf87vhxn12Z
Vst7otsGZ0hQQ3BmwIOeg7kp+iqXqvVDPUOr4oTvpOFLeWE1kZfFnt0rgN2n9ZY6
9nl35W4vDxLnWnvFqC0FRJ6JVp2nDrNmrCoYLCq7T2P4HRTLnafQiBdQPThxK2aQ
6LC/bOs9BGKR4v1a6wVJR7mW6OQrdljhoj42OHH1G6Hrl/mLnHJhLeqC8Y6dyofQ
7e4cM6O505gLENVJN7u1GsoinStG//jqCX9yaNATjANz//+NtD//GaJJ7QsgMYjn
fYWEkK16u/oVh+aknSjiuub2oT8K9SKAB/lO68oBbcyfWsw7h8aiTZIiT/EuoY+a
e4d2Ty1M1Zk/Xxl4+v4u9dpwfGoLLyz6GKBhO/+9TvLjih1HN7KKE4aJ9q1reF2k
mj9KOSkt+NdT/R8ZmnSh1GpP4lvyhm0o9hdqyQNbeLc/xqVgyqN0lRj1gKB+iI07
iS9p7qpTuWMp1xmruYMNLnugOOES4GjpQhzDq6sOgDp0TnrHTQRADh6slRTccOiu
FRCKrma+lBt9+4REDjTzT3kgZ2H1vBJxq74c379An5xeT2KIj76uAmhlD8Ao7QhN
XKgZhc1wqDzQNQaRIX9Ermu6kk9HImzATfusLF+lAC6oOriKbd39rfp/sFOeJpGX
nc1FvOZBaaNgem8S1ODQRx24IKHsQLZ/rnTk863Qk2NMUsnSjZLMYSe+o8JVBaQm
nbZQN3G0dfhC2CEQsnCEdnzZkRsvL4w2TBDIAytejZa3UndxtmtSNH/MeXLmwWwQ
OMo9TelQDbKOWSPxz+S0BmV+WJ+kqy5OPxzKcrcRk55mw6GygVFOGeRHkeTz3kBi
+kKeXiKWzv9dcNyETM6T8jjOc34AuIJ9rMFTyGi81egn2PSUjtqLkzWanbw2htjZ
YxatR+UUjSHru3xrvrC+cRK4ST7vwsDuzvS4+UG1BnkF/hBtp9Xzn9oeyLeGGhws
yzM+PFB5NWtAA29i3LircMqZD1skkVSmzu0Daqp4AzPwiTgXyFaN5xTpkEW7K74a
/AlDc0FmZLw2IfB7ZqUqmfFOhMP+Ml2u+373lxuF/cDdZosiMqu4PTRKLu5P9FXB
b1SlDwQAgQVmN+MhxTqW59FtbnvBx4UM9OV6vhkG8SAP50I1kuqB78T76dfKWuk1
9j5ryZLaovuiprPsxmwvFv3lMtcirQ1RZ/jU8mY3+Y1GHi1lM6fLPJ3oz+DZ2uu8
e2puMRWQ2t/Nl48/WaNLGsnttYJzdOdqGK2RavFz5dzvP09P+4lsFLDACq/aZZ/2
epK1cSxe3E0bNaLxe+Po6BEL4MxjmxN/NJAyKS+sRj7A34Q6IxIKZgeTnbdcAv1q
qLPmLan3NgKJPK3I/tjXhWSH+CJnUua5TDXCxa7/zYn8PUp83tdjaZr/uqHLNB8W
EYCo0Mhyt1Peef9lpT7DXT8k8LkZIAHgpbqtEKyfbJ3FP9MNNO0eSc0VNqEKfPqn
H5hIdi2OLsGH19ivFQqEncnt8sW565kAqrJmt8AMEy6l7UhZbqqjvWPpYxx/IAPi
mYv7di/N9MMGghYw/RDr7DJ6B53Yw1xYLmmtxUvDi3Kr0cY7taubkeV2GmliAz7C
25IJFL2PjS/oD1UpnlqYwWGEWeOs9Yj+42dG+81jInnjiJ5B29MVsovyWVvsP+C7
5Z7Dbh+nhZqsS+8AciVIY4Hbh2UuKuIqBiEqaSvCpASBSQu1Qs54+afFdAJJ7R+U
8TRUxzNUWC8sdNmNbTw/zqnNI+0T6Gto97xeyLU+RCzOyOQxhOglrMsW0hp4R6m9
kRGi1LDspwMVJLTogPglaHaeV1W73orQvQ8ggpUvmPQybRrkiAq4iLN+cRTdLi5A
xHqWrPuQwSCbUDOKBnFMaRStWU/dN845sfu23HTXMz3HFd3w/x9SppFKcsiQxifi
wirkZiROtmiNmF9z5Yl2/wDOoAgSX7QE7nCha0W5wTxeBjt9N8Cd/UZPRktBfreS
fie0gBjRlrSviyXKc3J9TI5e4FuFGO5S5OsRn/F8jpERSW1TPv3x4DlPTUyM3y8y
uzy8u7KrNQMGU2lT+0D/dVSC7zFIc2OuRyVIOAxfusnhVSU4NfXtah8CLyZZgilv
vmhbCGeP6hsDA9dRHSDjnCxLFp/Z33GSEev7YGUM09gS0fkByfFb3/YwJI3vdxEE
Cg7E5H9xErXBxwcwYhDnQHMl7qJ/uoR6Esy4DMZOHfmiiLb/JMBGjJ3jlCDBPI1B
hCRZS2IMkzpAtG6xz9ZKif+i8dotHa37MVwSSSdUW9o9nBSJo1OnkaX8nIpCXX4W
EipP8NfPtImrp7l4qa6vyOZDylFxIhttDRf5MGAdVDuhUAufBeC+p2ws181k8bOQ
JgvHWwQDOkQ2RCDw+9bYUjhEh3EG4CrEzabST0lb6KJAr8VEdGsO+ky7vv4vvozX
zGAwnk34Y3Y6oXZ95Z/tGJ7mEGv0TM30HJJLOK16y7cVeVZ5KB2qVzt+4m1lI3Xu
RSGDT/SsGGQmnjJDOW6M2eniqtWUgADefeoKLi/SdQB4X5/pMU0q0Tc/NPiWgj31
FniHil4t6MuHrc+efZG4X968gOTq1R8EbstoXBjztRHT7Bm1cakum/jy6GK++Q9U
ls7j9BrdiMp5s8nrwBgVT4AyUtf94SkkH9J1fcI+QrF+oqV5VT9aEzP/pVLmxKam
2/A7cKxgv9i+RG5XPAOhsvJvkTRX2TqCt0pVLGL9PvpHNm1+fh4ODkFooIZa0LTB
aFdbhxn5eHBciygRqU5FrbAhQIeKVHPFZb7o6/C0BIjxbnuwHWSpUnle/soJiQe9
BSGsXLBFcwzEBvXyalsBFA1TTKScZgUG0Tm2/AhRqJf/23cufcGkNW1/89t3K30x
QFIYkC6t3GMaEX3cjmtTw2LBr3EZdesOoQVucRSBnAqzw9rJXy8lumwS9cZrRhEL
9GXqGhJ4cx25UmYLCqmSqb+wtErhkpZszFfHt5tGG1b70QLHVmAAIJLNO7SeOQ5Y
SygoyXjg5vIqYjtMmxLU4y7RT8zyLNTKm8kQPM2zVm26FqEmSKGku8nOUaWHSyI4
6PT5X8dZ/qDiCVUjW9i4UBWAgpZeh5BQClq6Egmjx9i0W/FgxWCmVip/CTRc46cm
tV5TIpJGg+9HJBM0oECuCTlThzsQz8VCP3S7+f0OUdZbZmIs2u+zKoNIdCWYOEzI
sghbsGIQO1ZCzn8elDkXAonwyioV9cEYHjWr7WsV/3due8uScZbIRbdbR8rTwbar
KYetpWvGM5YRBNPhL0Yc96kO6LnsI3UYSx7wkCIf6w0JrkgwWqvAqOIp+yXGWxDI
m/kJHwETeI5qvchdq1N9AwdRq+vEfoxeOg9nin7rf2eDH0idBvbhZgf7A/B06ui2
cEdKUPY2nHmIMRc2v0BbwmXLpJFM2JM4k3BnpErsVMSRsXW73H0nEiF9X+AblOKC
QjbaDr/ocYu4L/0zaflqdShJbv+pTgndQhyxBTmRwNw=
`protect END_PROTECTED
