`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iL1fotC/D6IzKnn1UnlvXdQLocvwfgDtM/GbECfxGktB4PpotLCSjI3hoToKUdbc
y5Dz6HS9pPbSToKI+0puCfuO10Goxpcmc6G6IOsbc3Cjk29Xm4y/aZ310Q/IbJi6
w5j25o9sz8xIq3q2IlJV6MmUH8m27diVHVsGifslG6kRnvVN1AP8koQOVB1VVH/7
8+1sYqrs+B9RXfyc8ey8yCoQqNBSzSnPuWztKGcabgvUzNVwMdtaORLtu4QG6kZ1
eNOWNIGeewxNFxvLGzgQpabNs1tRIOYCC0KoiREnDeL2/hu3FvChZesVRlwNEPHO
+0IClcOvyjftjLg8ocvmh9F3NjhGgnp1W5fyaH/LSMz3nGBVQA+kL3HYzXx8pmGc
oK5mZiA62BJ1PfVISPEYqB+taIB5fcnI1IFY1v4H2au6bR2iQtdxEQas6OudugBu
yQtsCidzP7Oa3pYn8ijys3BIIO1Yk1FEZGQHXtirFuIPUBvtTjnrSW6HP+Qpg/xF
`protect END_PROTECTED
