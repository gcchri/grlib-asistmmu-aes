`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uatHiQCKDSQvwc98XTplqzWH9+DKf6dlLCY6SMJm6WBVk0PRmLjkuAvmFtDR/hZG
PD9MfAISoet9f1ODEGwzurwaKTcPcqY6/anVItJLsFxIXvOaRJkkS7ylKe8x7/6w
HyfFItAL5cgsTu1zqjOjwNVzUG6i1tmdcJPhtAyRi/sZAeqG9ku9i/lJxfX+3BR3
UEZpQX7bFJEgc257yj+xMWjdwg6HlVlLPCsGfSS5lpWRhsHaLn2rofA43Ow3niDz
bd2Q8u8wqPWFU57fuAPBYQmcu41hfKValAlef65W/cQ0a9O/z2maMiOe1jD4N5Ge
i6JLdODMm3ywnDiE5hUz5FSNc53ZRCkGNlR/LfWWlMX33jJ0i8DKi1KxJjFmPz1T
CccYTW6c5BZOxKXeM/lMvh6NYqaoS2XrRkQzgae4Al1X+63qUf9bGOFmJ8/xdUC6
/g1/6BQHDCiHoDWbw1j9VlcgopUbi6XL7v1CA7ftGvWyWKgBZZXBeJtWDHIIK/nw
`protect END_PROTECTED
