`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRhhR7Ude9LUoWNgqAMCRt/pA2e1RsYbAOXswUH2Ikolmh7AclmtYP4O/tRIsYSW
LG1Xfl8HPfliCaLZzWVbw48A2M6zFX76TgHDJ/5hICBbnd1c1cPLE5eWDY4EHGGA
yF88G9BSCdAXXVf7lZBEvL5TZX+N30gS9Aj5YUxVh8rkGx66wBUKWsy1xTHzdQ0g
vcW6a2vren+i1Prr6toiaPWXQSRAr9Qc0NuE2LP3NbxuxtO2xSrVPmwg1nOyBhv5
fqY8Tw4fZCz6tiIM9Mw05krjZ+ZyLQldPaa0da9ydpe44M/7IJ8AiEmqTUXv+hbG
1lW0ofOC8MX929y7UzhVrA==
`protect END_PROTECTED
