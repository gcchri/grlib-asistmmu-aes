`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
onubKmLnGI10dI8DI1pYx4XdR6HG5RdAkkUwX6MPrjdLptQxIM5KFcJE0zx5P2af
ItHPcEdX5Fcf/2cjbed3Vka0+mZzaV4xeY++TBFZuGdWPRVhmtQ2nJ3J2EyaCYdp
NY6jodL9Sx43vmBxw3wy8zXffPqG/9qQDH35Aof+z5sUqYGWPPwwCFe/H2i8UBjZ
DmutcUuwpFaMspfV+sCtW2NPOG/5RL+1CoV5ZGq2OUSy9yHhmrhxW18Ih78QeU+o
`protect END_PROTECTED
