`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eG1Tot8WEwtwyD8pFL/G0tNYdzIS80MNxMEjyYdu+k9iUFTEZYcztq6kPp/x4km+
dH0/e9P5ARhxH+uxnFwkPfGIO/+jWpSMcKX2Lg/AwtOlQ4kkZUBYBwcyUIx9tsPB
qJomrrnI7KohfQPLaLD06M1C9ntUnQx4Z/xaj2M0QoHAnKiWf0lscnvQm5uCUY7F
68VWkB45PaKmGIWDMnpZ9UDI6KbJkXexmpB2tPHOatLR2WNHWuKAB5ChWQQI2/Py
dhUVVmM0bw/zVs8cnxGtVHfPQFGlh4JUEJin8gK30WwjUF9524Ghiz265C2QmtyT
LaWQ76mjnMkf1wF6H3ispA==
`protect END_PROTECTED
