`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBf9qGZW/pXS26J4kCZCJuODn9EsOQj5tErsEhMpR50Y0T1uowyskVNH6q32VqqQ
ezt0pQT8ZoieAPezmEEbkcZ/9nHGbR+k2WaauYhxfXkZk3GJzdQrFJvtdKtGgdZM
vU83R+mZE01GamLVPI5VFJ4CCIJozm3lOByRGFEE/xza1lcLHp9YSKmeoUB0MPPv
uy/S8Sli83eRLF+YslO05BQbgxCdCetMEmc/4HhQVOMlUhIGn1lllPkEbb/yOXac
7K2XOyzU3Q8BOGGEMr5Qw6icbpdfbHW0qVCR+Ez5sMD3Ycfl4kmJpYCfnzLk9w4V
LFM66jxbi+f2aKMlp5K+L74KUX8Zdl8Aa6NkTFSzJD5JniP3ks+nsw08ULSqMkvG
YVdzDW7Hold3a1TJf5mS6KLCuYaFygsv+M7lNJQEOAiLm4ZXwRfInsrZd5DUozVi
406qZJcPSg6d26UlGrS8oQaAOIgn+ud7VP4/jK//XyL/tpiKHdDsmoGOwg4exDXB
GPasAab/lYPm3xzHgg5t2HuYIuog8JNrox7FypG/Q+24A1Kpyq1R10MY1zHuNm30
e8dte8kavUL2StLo6jG4TA0zttnE4mHaaXHAbRXOZcxQuq9qdy8GF7ZhSxyBTxot
`protect END_PROTECTED
