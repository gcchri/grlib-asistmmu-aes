`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9iNvq/stNhy0lMoGjeHRsnw+u2cMDmbKFJ8aiHeSmGBYidJyjhr35E/3Yw0Z5e2
WQfgS49eL4ijDLW3wQpufrLbIPBLQuxE/q546FI4XYDPhlr0O1uxvCgjNl4khVbm
xGxCZ15ywSjwdUlxQqxmt9xxRV48Jlq+Q9oUBslUi9/+s6zJtxipc6chkiylYIPX
Q7n6y9vhc3v0N//zK2bG/nTcLD3B+bU5SfModzGeUjshp7qQyDaDSn4Or7JYQoRH
fxxIDypXgXl6CHVDg57OUusyEqpujmjJ/vLLtX/i7DHFTeW8JUk4PUu0SHM+TORQ
qLCKtk0K+8YpLWsVY+XQOxQMH4CbXaym/wVXO5kriHarRbaRIDzdsfUrsrhbWCq3
WPy/dV2QXySOQ8eMdZ52NmD67M9eSXSaySTV031qihgzqbP3OUwM6YyK5k7uKQaq
yST5yPfWfKVMNkm04AJIH5Os6qRfOfcZDCrn/CbjI4B440obbJsMKcXXEtrX0gE+
zIizqBi6VGvBXT6aqtfgPOar2mdMeejlnd2UI4UuQvLJQTOb/iZ4eY8hN6K0FGpW
F6PwW/09xHKItQrtYQi+8qbmJpbhPXKlJD8JyCYSvTzMRlRGfCFoS9eMFKXWAE0A
HMfANhLyiKJO6zyxT5QYtw==
`protect END_PROTECTED
