`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVqlB5X1RnWU+9+oeZ9oGtkLYuLanDIJa6/rDnWIWHSLHtUfkpq6REdzBpNMP5ri
2veSaX8FS3WZas3lwCXSAz+ZDC2zYQXi5f/WM+v7cB9JRF4CffDCtypQz4rHbjRE
YXIY4PUWg/EYiSgv8LO+J4u6QanQUzYd5MSYQ3swXwTOwarQL1hTOjap6hORpdkw
Q9mSRWLLniP5VHoMgirCWw3a8MGmAXdujAaEEv38uPyt1skD1SjhARodSEjlbZ9r
0dJdB3UNrBdMJDYlEgidwwPDoQLppEaAAUGoeVl+Ysg=
`protect END_PROTECTED
