`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g097WQBkLkJum6/+HJon+306sMEAJNXqsTex2U3UdwQcRHLZ0EpmZ2kIYuXCwR6N
tsuoAVtlu/ZqKmh4gMSAyboX1S6Na2pfwUrUurDu7vh/rukVrEoZvC+yM3lXlaJ7
ydH0g6zSReoSFIp7G6dnNulgJP+8wGBEgdTTx8zVkEYtZU3Rqft85qUo5hV9bksA
j5ZfDzFkJnEZmOeQ1U1STOzMJPDIjgBHSs/yM1Kvr70TrxHWUomLZqOFnoZsxWR4
JLp3kr/OXTY95z2RowihjT6vZHl3kJkD7/u3SNFCCV6Rgd2n/MYLcwN0PZbFJRXX
iKpZBT9qmwZTBx0KMYz44yT1WOG+FJ+juuihc2SGMML2dTrN4cFfj4xqs68g+plj
HNLqA5Fo3vjJtXHsFjXpBfuph9bsLGC7Do9rwop4qoKmEA5LsW9hqwHgYiVenOE/
wroiNSNFsIEXkpuedEB54/7njGZE8Pr0qkYvthACElLicPi/Kocz8Zsr1q2sTCsT
cDwIUtSz8Ayn34UPwZnCc0v03tpUguADNrhTv7qd2ImHgqH51sHXutD/66HURdqu
GfJOylxmdO9fLpendssoOu5vyLKntYapOWbz3DjdzWScXQyGxHMOOR/Sy77YYdQb
4mznra710XQiNqkbiNqQ2bwyh2mygQSTPIP8PiH6vbKU7eRXTkuO4hnjCrDVGEu2
DMOqqWWhcnYDthsXb/KjiX+4k5dPC7XNFPuyyhzQR90C/cKOa1GLCxR5cg0gMEbi
`protect END_PROTECTED
