`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNwFshluXWD/ftyin6v+bcT48FaqvELD8T/9jy9WuYFV7CFPwepHkBa82pAMPge4
u/34dWvIMzm7evBr+vLfzuev54rKoowMILERDjuL2LSPfhu2wWmRNLejhy4JpGVV
rUrQQAaQpxiwkJNYjYHrJ9FfVFs2hWavdI7u0FuBF2g2yhrBHwJ27N0wpVaaGwxL
ot+i1yUJtULZoQ69zSHBhhpFmekJGIIUH3YqWqjrw1h1qxbbpVgkqCe6GyXfu/x9
RXAweSBk4izjv2w16yuM40gN98x8jfojmXz2XhzGLUV0pCO0IO9NJf/yS7ciYe4d
MCplCw1IM/EL0dTsX4wO4nRBc4HfVGJ9HEIKlDxK3fjQT7l4VI5bDxfJwqF9KHr2
Gf/jUj7GNa11834kJ3gNh0FNudVognMnJR+lSExJZeMXR8FhVKbXl+28iHDtdHO+
H990c/hHTsdOtenF+IS6n7MQCXMDLIbx37Qfv7hpwKNYMxzTiZ1I1MxtwoUlL17r
`protect END_PROTECTED
