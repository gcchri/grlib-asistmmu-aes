`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
31DJJtPURGWNRrfOzYwglFY8s6K37TZK0v8qcDMt8gU4sGU3OlTjm/kr2QAaaq1g
r8pJOnmiuh3hrbQcRF6qyrTajTy9YI0oBGkLcOW711kpiNDMPSU6vggDotG9by24
7KAOJ9HJmkOYKZUaPUJnewdUISrsc32c6kjYtFtaAhnVxAO9ovx4xjxwLsfe9SLV
ivPuar4+fyNQOtfvTiaIeAXxXZPkJGmonqOam+v185lOdrYXNMIG73WD6m9fhhc6
MrxYpzD9RToJ7TvThJO1ANZ41dCH61LvH9oqcBcP/PL7N7pm7zG4Ji15CfHKaix1
UAj05ft/1BMS7tHSFwnlLcvWv+gxLcr9T9d1RoT+ZJAFVVI+5AIv4YW42kbJubu0
UIhHGXzy8vSq8sICnMZrdXMoCafq/nBVAFq4Y6h/UZ8=
`protect END_PROTECTED
