`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5MGNZvFhi6rwBJD9YNYRHcERsfhkczqJmb00Vnl36VTn5/xtCIDD+gGfp0Grnf5
4GLwdHXXF4A7lM3a3CeF3ozwOkltB6elapQBnoJBNlpfqcPckhW9mCJvz5xA2Ouu
3O6tKQzuaohiW2krC86dEmcJag/SNqLKDq3/NUJMnRxYV11CTC1X6NeRvhxqRLoU
wbF8Fct5/kdCAa5XSL5XkExbeBubzt823qK39Bk0JSAEtqjQjLL/3ESxme5ik1P+
gficsYJHcP8BZcYb2uqEP0lfrU7tbZF1uTssnjuMG+N6UE1MVDkMvHDlpJjWWO+S
15fneSrCnmp3i9ceS3muZwanQHd+5Jsk48otkrzrSeHMr6mYQ9n8KGzGVj8o0Wdm
CJ0m85mGIm5AORkqUplbtF4UXvFatdK07/0aWi5MJP0XtxQp9+o0Fo3ewf2eR0AN
84V5tIalK8XUxoFNJQaM63TSjte7pstiBbqNzRKto8xJZbRo5lLO2ExCVtWry5Rc
D9sn+UQJPl7Z/JSHYidMYmcbVOS8gntNh70co8mQBOOlQZq4f1PqH6mUkgVXTmSR
oXNTcyUaLh+70jgXFcgdrH61MQ4XSe3CQOVA6xO8kiM8c0Idb7wb33sNoPu81AjC
KQKRohdgZxb+PH7fmSA0Dg==
`protect END_PROTECTED
