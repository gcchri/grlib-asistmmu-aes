`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n7eVsxAeTdYF22CadcjIh7BFl81UCWX6OvQSXI+sneqEdyUU604CoaW3kpz4FgLJ
sLxqZPnXIDhGgfgnu1NsoKOuKxR8bbLbAUzByJ912dr6eZTKMKH6tYBNk5Y2ICEU
wH5UISaxZhmXNioawv57HZr1HGfHIOnB/oBIzvdsbnL88+HGx5ZhdAGQkXQ7ymrV
Tp/qI/M9ZoWgh+WgEAnLnqDGeJo08N9ydu2/LUoGBSADBfsvtL6QB+P7waRd7jDx
GxnikEuCizcIAAC+EgWq6il1l4cpt2+MLtUs66U+05830DkPd89geLMd75beFI7F
4BGhdPJ6qc9qdyGcPAuxlpvbt2xfPoAMHBFpfdRbydgvne5BrHA//a/LkqDJXkUP
wLh4wjoJUxcQGDnsGfN2wXaW+/oqMlPZrk7+M+kCppKvd0TQBacTw/43Veczdx9j
6lYB35l1PrC/7Gw4JxhvOOPprbw41QeS0HD6pH+Q/u5e9xW14x+Pn7fbHrUsvaus
9Hnqu/1UPh9Byom3DNnLFzHyZf8+kzzGKgD/jM2gmLMlTgnOISlFXt7xt6B2Ove8
aiCakFKEumPasvfd//F9Kqy8nU7LfctlC8FKf/2sya+fmsRSXl4V8OAf5je+Ecpj
TCxRGMT5nDXrtZlLTyOgS98p5umQi4pn9abfw7mvQKoQbm+YMBEXXXNO6t7N9kGq
4xu6/qpYQXFMjqXEeKiYoB5cdVYmYVAAgNW+dLcDWckIYHH68XkdC+hU+hPpNl21
Bm+1g2qadUA/mRGVHbFKtikmHCOlewdhjH0fJODdLqmc7m8jlu9/uXLgE8qfeIm3
vlLH0t810L+6kWXtxHkFrCPUBcP1swMywDzcCD3eqbZ9iZE8BjOClhfo0LXHs042
8riPu8n7yPk4/FfkpkrRWirGGsF2FbTXL6UETUCLPhC0gzN6D23SSHNmul6/w3i1
7PCRejz48LjxBPrV5NR+GpLEy4gG9YZzCUk778Gw6s8LAQwTwQ5gGJz0JWeU6SEa
sDKl5xxx1lK5G3RttW25dxvcsWVV+jvegcRlZD3Hy4c/WY4JX4EiZzK8rwRPgJkN
5snpDjmrdchFH7cm74K4aeI6jLod4BV4dF8E84coM9UdKqdOMbkUwQFStGWe4w0I
za/eSwug7yJnZMrO4NwgMKT4oAEofyd8L2Lk54CHOcIA6Rgg/l0XfamLYLJNk+6w
1rX8eFvcDzDZJZAbGY+GKFd16DZNhOIIqAXvE204Gz8lxQY1+216nszm9JZWjxj0
ahxCw4sAQx+L4uEcGz9DId83n2U1pK2OornjyXovNNh1163uqM2xA/18mZaRmDjq
LP7NIhs5II3kYp118FUwEw==
`protect END_PROTECTED
