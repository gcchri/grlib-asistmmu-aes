`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YaHVQ3diPlqPhxR7+c823TAEipkhJgqJijchtDcueIAxPFka6+rW4+0VoxzRhE/D
jk/vB6ICQ3KB9NlwZpXkjHura5hqZ3c0Tyy8enBz1nTrEyG+n1v3UdFl82DBlurH
xmEroLd3UMI2VOD64nfN0vrb/EFFqhLd671siZjFYMN2V48jxOlXwmTzG3RfOFBK
pct0nCg+RdUXjn+JVTsieJn54ulkxnoMJ3SysF3YRqyYrzFMTnZznETpl+K7Mqpk
C5hXlAII0OHyjZT4wGNbDjRlWCWykGaYTEqnT2/HZHc32OYgfEw3c3EVS1HzkiG8
WcBZMX9RwU1Ew6+u8OHOLQ==
`protect END_PROTECTED
