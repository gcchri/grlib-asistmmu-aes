`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSv8t7+zsSre2KcOgKGCKxFPLEs6q1UPJuSFKmVIIx/tM7AQx4yK1AJ14VtWAvC9
Vzp6knVbcuu5VyduVGqJWMN1G0fuG9I4f7lbz8/V1YJLE9Mbbq/1meHRsTEMsdfV
Ye+RGFpxbzCp+1/OMG9EI0gkU9reLKD6Y5stlyYcV+MWR0mH46wuGk2zfvh4jOY7
oO38SQ/GSzvq8bgfrczO5IC1tMrTdr0KGymhvtVar+JuSiQ79uVw6puTjXVS9WPh
/Vb6toq4R93vtiI9wPtnxVrAsammXEPHgpiQIt9aRrzs7gNP+1gaVRF6qrxU7m3B
BiwNbx/Vw82SjCSjy/8KyC+a95lGYRKaTEaD7PxqhNadCe7my54hWAvBoGpGW9Ev
arDsYi5TWVi4ZhwvgVTauw==
`protect END_PROTECTED
