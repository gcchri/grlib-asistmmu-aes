`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pe3LDTKC2nuSjntIfmntUtk6HnOuWIdw9MToOA0hq/dy2YIZDl5NGv9PANs0/aSB
2DUlE+1Imhxs1ApHl2V3YXBsMl03h4wNGsx4y8xt45RRcSKTlJ9kMAl51vNn9Sjd
M0FDbMAsyLp4o2uip98HUZ6qTwd+2+GZIix2OdyJFy7o6djjhaNWllrQEYTFbfOZ
mey8TWe77cdW/F4MJyCcdDXeHJFH8cDXQKJdzFfvE4Z467Ac7PafiCdNKeaZzzPr
2TJXNKqpSic1lAbgeY47ca+axz4PBQwRDEJFIskRGXdO+NX9V2yr47kBlZeyTaTI
GvAa1ho3Tf2VvBDIeNW66YKjKGi6pjAoOmq90MQQLSa0006sHXyE5mmtp20B8HsP
OJPSPvOqXECE7fn0BasjBA==
`protect END_PROTECTED
