`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oRAfpE5uJKNTs6kaUfsxxWXWiRCPHkrR9DcYzc3DTWalpJ4WpUGihjLyR/GfSNa4
qaovJcKuk1y3fCFbqnhmKiIxC0e2PoGOu71Eiyef9olLJyQIALlZ/Jr8o//b9B8L
w4BOt9m7LwVRqg9xWQvGvVwydNWmZZDLQb0LWVWBugTviXyjxc9HDSUCMHMiMUqj
G90u0koIaYpsIrlJiOuE/ejk15HTq+PANQ4ToSGrW9aNIx1VMOmarfj2FSg5OXOQ
l5ipBqLRrN9EJLILP3yf/Jte56yhQJe+hlgyZnTABTX009BCJwAZfJkUp/bgEStO
5iU6Mwh8ZZNuqtNoaOooLoXK2TBg4mXQvdPdbSw7KhNavlTmuevIr1YojBeYL6I5
IUVnXWSF+4RffqBS5TER+//yvHg5gHCAMmyXADPQBFTwBqa5VgKcc2q6olIMov+T
nm15LfMP6vPUXmErxpIpSWhbtrkPrFgizZYR6vUMWoTtGmzkENgetWbIY4299cUS
7RTKd1jpYWf0bruCVwQpgUI6Vhr67bYMvoVr0DcvqPAJNYQjuhG9VEbbbKdfDIKv
5JJkTENKuOVmMmEDZwW61hlJKx8vyjofFj1503GM4dE=
`protect END_PROTECTED
