`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7aP3g8UzcCYQhQYr79e4qMhrlnr9Vaj642OBJp0yKSvt8FjcHYXNxgC7LzfemPiO
9iI0S/6mfgTWEs77GcjY/c11pEw0ja+AP/xpt7dfr8Qu1twICEU5XFb3XCc+Vfxv
84C9dYD7yIITaQpUSqceimTVy83IzUoRvl6DC47sn8j2oo7IQMnE/1+NyT/w1aY4
wmULKaThp+ht/2HwOdKeiToSQO8PnYDNe8RDjX5Zh6QbduevHhQahYANkW7cyM9z
Z5+AnLe8fSt4IxZxi+cumjz6XruBByWkyziK+JLlymreb4uHsajJxmN//zjIJQ1Z
XT3zAu0qI6SZgETpApHFN8A4BpYcEPhR89J9Z6rPwmKxmC98fExml3UxxzJ86yU2
SwscQN08/2Y+yMfvHbq6kofcwe0pURSDYsuuoJGe7xPnbt+wN0F4aywDZrMymTsk
faH0IQngc0Hm4Nu57H3JsZWIHKmQMsXZ0QSZ0Wl9JIwFLzEhUEbOS5kt9n+tSwBp
GU+Mc8cLTFZurViDMrYr0daiX58xFhuQMpvjbeErWMk=
`protect END_PROTECTED
