`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pZMuKGzo5q67L9f1Z54Y0GazM0SrLQ9K3+KPaneeRNdxyrxrJdEEZLCGjkPnMCi
pZKRT8QcQ8xCh1LdJQ0fZ3VPMGa+uwF87NchJwNY5lHAnr4zD41TFxN1N4YBM/ae
028emvXg6OEFnpaBBeE74Wy9IngqAMiEXCKG7MbCATSGys0jCRymAv8jiD0IBUA+
cfGd1nWlXXIguMM0EfSYbjozLYp+39AYQTLoSCI7WSk9JSz4PntC1fwmorrL2YR1
LcMc/joFYbXTFJ3ahpbV2NlvYiEm9x0VoKpP8VLFE6yFUFAj3SmZvoa5i4rXl+Mf
Z7I9fCwSWGBOgaDAhtooGUFPonmEXp9Yo/BSyjDJPzyXOOYMZiN7FrsONp1Rmszk
`protect END_PROTECTED
