`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qAyMJuuRwrcYu6UwBK8t1o5DLRab7VbWsGN7L1mgsFVuGEjTILyR37t6yZBq5a0
iRJKOPwz5h+G4dO9Ad4ltexv8ReK1KXYgIJo1fvvEPQQ65EuCedLaAW4sUEftJGO
5l3VpLOC22Vq9QLlOEOLC8zl07TmIUDy1JgjyLIPm632uIZl5J93LmOiNgUp8ZGf
664Ci4ZiSeLrINGWhhCfop1oRhe+/KhdfSlIxYUSWaHJrhPloaiYlebZt4HWknmT
w+Gs19d0eTM+Q9O9Yg5MV98G7oOox5mI2KBnVfwQERV+j/d9OycJI/9asncI7A/s
pB0bOGRBK0+hgmMkhuGLzjZeZM8WXXNW+R9cyItv3uZ1XYjMpcG27/75U6QS4zf/
nOLiToGZrVqq+F7fYN+6l+zUVpH3KcQ4ZO4bZQRY+aVZ/KZ6mVkGVglWYcINf8AF
Yq9MtFdpTzGDV7S9wo2FBK0cE/U43wRN6V/VXuIDxNFUIob5swIwIl694HdsUVu8
jljXN4nOgx6OteYk0fzK7NDnLM3TMhrdLUdtbnGdVSRnlv7XNs3ZJM49UMQNa8Ta
wAInZcANuXtwtU33h7YDjMJNd1a4PGuy7ObYZhxR60E=
`protect END_PROTECTED
