`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEOR8kL1Pa0nDrZvwGNMpbxNrZkJLmdgAVCq0FQr92Hjcbx5i1lcNdQYv5TdAtrl
HIie+W/EyiAbTdHeoOxjoDSXBb5v4W0RpArLAG0JKcR0aeNmkoum5WYdrg6ughTb
+K+H3LaHi9qg+zj8mgA63wN/2+xBv+rzSqjUxhepFX1K1kVF7OVADaBA/CzIkuFM
USog/7Os4Vw+0BpYV7MPy5YnDPh0n6cpBK4OFabGpBuW5rcDgDndOQSeBmYz46uC
`protect END_PROTECTED
