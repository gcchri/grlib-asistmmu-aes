`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0osnDk5Z5vcLHbY+CDZaPhE3acR6ebCSb2nWZ3S4sFUuRRg+yy0LkER1rnwaqvp
frz+haU73CWVyXjTcgcKuRHAwXe7RHOAg2jndhhuN2RGH1sjQZJAQ2pFI16vePNL
BQrAGc7gYko/jbvzszdumVYWacWKAdgpxvhm27OmmCwKDcy5dXOzEflKkqM3RCFx
XY+3GWeL5RWK5gG6eemF5+sYvfXm020vOIio8nM3OO5x/Cz/RuYfMPtUDIx+ZRU+
e6LdGhzMqY7rNebxaPP24Qr/Bj6GOB0Fwx0B/7iSNTZ2a9ghntHTYp/N2oLw6jfX
iWWZpTWHscZFG4la6zrGeoJ1m0YfYkKp2T0GTgrQRRFWipPQ7/sfFW2wk9RG407l
zX9lcp2lEi9IbkxnR3c1S2Pe1GeUDRaUPCXClucGnEpWKjFQ9yFN1XOa81z/AWvJ
uYGRyE0aZfRmys7ZgFPRAWuCQfIXsHvYnR7e8LPUTV4gNd1nSIHAlbbzv843XRo7
zzXZ+RMwvDJpn6eGBHmmCnf+1N7CW0bt4WIlMzMPBxMpJChJqKSF3wfCM/r+1m6h
sRrL4fo52I488/DYAFAm/L/ebyodrXIt7CP8B/G0Jj55/m0R14JQDh7IclF2F8bG
g13mtu51atxMgOa/xQ/6VA==
`protect END_PROTECTED
