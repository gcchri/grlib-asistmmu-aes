`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zIAhekyVbaJJDaZU5tAX+H7TmtfBVgknbiLOiSUFUEIrxpl8ZrhZ2HB+yLCGHVIO
yorV7ymzMgIAo+4tk1eGPBqxYv86rXg0xIVMF11fRhbLJhS1ny2x51H+P/7xnlCY
FOURWXh/KxPnc3YO7W4PJ0LvQjGbWq3aNVHE/GLVFjn2Vcxzh3m4nZAxWDsU2Pg2
qCDsrVHSIyuW0jo3vBTz+zirWVb/NPQ5/gHowxw1717eHALqs+KTZncvkxSV7sZ1
+cjrO2iylJTijO31jp0E1fF2YqeIlQRJK0uV1IcOmNbQTZkh97BRrVc7AuUaanTn
P0KrcJVIrkY/K7mAK03GA53mTftprwL0CImUABVP6Dsa1kvB4+K28GaSztGXRDbI
AMjM8xsYLsox9i6/1VC/viu3tucly1orHRotjJYVJr3rF0cGSwSolpfcqEVWN37C
uSvODj53BE0QWab62l9mbHmrGXGJzNB65tTw0LgL46t2bMxMXEeN04IQEKQ9RSew
ZC9LfgUd83AnZ4ld0KsIgnQawTqydDRHl/AhOkr7ItsmZdJZDJ/4QjYI7my9yoyp
puM842+U+YPih1LMQkcfsVwtsDSSDIS3QO97KhJLkR40rSjATIPNY/GKM1uBazSo
JUiEZCf5EWY5JrbchenD3b4YtWcJdvYM04JBvRf9Gzd3l3lG/ebSnM1ftX79DrMc
3QKALXeoNMolLYSM8VROerxd6BM/U+qbl9Ds4D5wN51HvWVaBn7Wmkx+z8JjRfPK
vRBxmReImsbQgnMHIv0NQnSaZvDETTfFIWE03zy7POHgsQP80q4KAFJ0dckU8IPx
6Y9Hn+A85gAYpb8LZWuO+r9/6v9jflDsMzdvnRvkCn9KLkKEsnyCx5jOc5/spgV5
WL6l10DyKsvL4RqTcf5LC6o0Rd7ySeyRhKEG8e1h/aEjRzeUKMg92dQ9n+yzIL2K
n4CiS7VtRrtMVeUf/J7JPTmXTn5z9EMWKbCtfeXxgry9aWsF/N4wsWlgrhAxNcgv
ctvCf35bo4rJezruGPs4ENlHb3DBrncER4GdcP++QUd35JGHuKuKPCN/W2be4bTD
fUXLsQMaksKByNZLdLFQnEgznqgzqG59mHyyCoHguUn/aIf93D4wqH9Noe3UoBPD
JFpIUaIhWeCP4PT4wUxBUIw+0miWguDHS7zxTZZ2N9I=
`protect END_PROTECTED
