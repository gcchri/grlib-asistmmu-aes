`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4brhrgBWT46gsG0tuvggmg3Sog7+RvlPpMph3DJbsMqA7kRP8a64radXCLGEzAAv
EowyAJPBsQ0FoTq1ppfRLJtTsrqm58FRH4ZK5tTH81taVFW1sQX4W+pM0x85fdys
vG8p5Dm3lUA+cS3WuUFtHOIBXoYPs2NjNgWv2VTeIy6XyqwZOZhMNL9cjWZRZAnY
/zpCvF//zNchkqha9kekFI9B3jjAgyZlm3knP5AiLDZxiXkAXk5sR83Alcj19I+d
QFm4sCuCM5Cp7Pz9pdP5UoFKnoeXjphSD+z5GxwrWXHQzYeoxV1U0DjCNJ0SQBY3
ZagcpmnEAKpkVD82BM2N+XMv4YZC5jx/nh71QyZ/NkZkNLP+OzznonzHK374/DEn
7MIOZpNC67XVpA0PfN0jlI7lZNJ2/S49HC0REB6xvltjJzQ9H3NZMMwPIu/I35jb
TYCCvh26X7qr2fz64dp61jajFTLJUvs6PBbY3Aefx2PlXJSP/4d6NguRanQHLAZa
O5ARD5qVtpAuqA+Fj3oU6EabhhgeH98oFd5FktNFvGjynpgX3pHWBtVM3aYj3v9/
WxUyagBpFy7XVsNvwGWChhTAD/Y2W9afCu8Swk8hsAFCIkI6A0xSWRKAVPZMD6HK
EVbaGyqFfwibCYRjrSom239S7MYuY9pzm58ZqYfaxzYQp62fdOKkceLnN+cqUDh/
zlwbmrIqu1hyTTnAd4v4ih9kHz2kOjJgZ0nNY5WxNGTIdqvK1wY/qsA+7HC0eTKW
wcDBYE2ACfnnQCF7UNep7+byEo3dX40KT/XIuNeW8o1zDXrbEdja4RrRjRxORpn7
6d/F+qo/9W++4IEhMtcR+MVt8QFHNLg9k5a5UL4KwXQ2ePtmKFUsIGAW+A5zQoj+
bAcePGw3drbrkk6wbZLpulbtVJI+DHwchvV0LlezC99Mh2xOTl+e+KF2ING1Tfmf
lgj2vrzv1G7rCdfrYVcrA3FcICIZGB9KaIe9S60z74keLMyj/MkOYLe4DuYra4N8
LEbwawarGI6IeXYFGC1vQW9Rhjws9RLQWnG7a05ZsLv1rOa5U+Ya1CjcpTtdogLt
U9o5XDMEHERYpWCSujIrt8PWKVx/W/SgA31Y5ftpdyh5RyZ6DzbqWoIaHgCAmbsm
jFC+HjWL2PGXwMefWqoviRFZP3Ac2TcA3pZqE2vsSuN9Aw9Q6cuiAQoZ834Ld4yW
jiJH+/b0yf6Wx6Sy21VaCWx7sZfR7OqOJ3fnaxEdsX2lpb/32WWx24LvNX0b8iVi
ilZubxr82cN+L4Jpcj9gNaUVUap+PrgVfIuaIgBnMab6EzOnH/ypp94vvqq7sjsa
ZXOAtYR74HPCMCaxPTSPBfSH2K8uz3d5WQsrUnV8VcHErz44DG12a4NfeJafWcEn
6fgfpeMCqpcYZ34Nwaqnv7TdusYb5YnaFaaXfIUfD1jn6J0bP7YkXzQ9LMf2nJAp
BkVrfWRGoCvwgQyb7csmc+OTAXrjBy2gsANpU+PGk0PdCbYAFT36HwnyW6ZGIoSy
kGcsGw4r95qT1nlDIzvjnGfa5OxXX5WCmhSpZXJmp0g=
`protect END_PROTECTED
