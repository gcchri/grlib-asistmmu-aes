`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Qig5Di9/qC6X+cHc26x0FXv3JLGK1YgFWf2uQwEgRud+m91WLrkomLt+YrBiz4M
61ouLjueKXV/zo489l+4aPRFakyK7ohnvoFk+nBQFgw8W0hbpeFtZBKDW+sknhE0
Qmgx5eRK4/IelyZZA8EDYv8jyCmDhfzXRMdKWJo4T1GP2H/7LLtwvJBNa8xZSwzm
Zmhx0yVq0ra4Sgjmts0Fg1PhNzcmhAaqx2WR0H54p2TYh/aZ1I+3nJAkF/a7u4Tf
mVLfrvdi+4TLLCvVo0z+xWSIyBf4AWX+YhYfRLm8VEK3bdkk1tpLyXJOmIdnvXnq
9F1wlK2VsxSO4vzA3FEETKpch/k/yBrIug0l9E5OtVuFQ7xSMEbgq0LBohN+nle0
jQS32F9SdfWNu1l+k0AKAU04YwvjZZpsmkGMb6HT6Lszrp1HMIIKSgaIsLEB0uWk
ZyhFah/lbkmWbISecfis666tuWinPbYlVLYdWqWNQuppXTn+TIptm4fDjfkh8+h2
t/bvNxH5PTSDgBWpksmcCs6f6iCTfniMnKitGTzoNBTNnjrPbqb9ZRTvpkcoA7HP
fL1iyxQeRmEbRdYOXOL+9jasTZuXsq0lMSuhuoLPcqTKnreOB9hu30VQVV6wFoVB
XVGjWoY58Zpz0ycA/AMnHg==
`protect END_PROTECTED
