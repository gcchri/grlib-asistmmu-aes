`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gxPqHY5GncjSeiHRfU3ZgOAEdVR872nFEvrjUBLvGLrD0iW2OGGG8gjXR1+scrn1
UwkgediRFU80pZpNHEzlWMuqNwg/1sdQqjKN401gyr1mc4Q48TQxuy6Bma2bVpax
AIDPAeb1V6tgkyAKA++OCj+jriykVFf5lUM8hYc7oMnKKo592Mx5V8464YGVsVkZ
OvTIEgRMRspdbMqubUPVkhuW3nyOR1IyON8+rrGn8F3giSR7WA/EOUzkB18w6xeP
Mcp5ojKlIistQv3jI7RNU117yXgKgRKy73iHoznJWwovcz0lJmoeadIe0WGCOxOR
IYEssNP3v4qhJzC6+gXzS6sSrBvgdD8vIpD7JHC7t3cl7//m3MzEa1u6Ga3ePqad
aMDbKz6Qd+wKIBqk5Vc6u17hxwOW7K2JQXUPYyzquqMB03J4al6M72SfS2b0DqHb
qrma4oNC8OJp0sbe2QZrQ5G7xlK4pSTaceQFqy1ZXtwzglPaASv3J/wLwvgM56RH
ZrTrmV8+KDZ17Esn0txvfGWbshEM8EaPD512zeSrr615/RXdYnPu8vlrEXLTvduh
9nJNpjM2dINPMmwohgPnn0GSs/hkM89XROzym38WAlSDgPrY5wqJwruLXCp2S/jo
f7pa/0EEt6pM2hI2h0pEJKOUpRvVyAOrRB+AQGwuh1Tv/YHxdIfUwGEWB3HJg0kd
JiFpsSfgAHRrNoLtqgjgzwsqd43r8sQX60c+/2TAAD56MyGDZmImGjkCjaYm9Th4
TaWHvSPagwtqU9ABPHrg4pEHXxTjARu/jVGRVGfP+Uk=
`protect END_PROTECTED
