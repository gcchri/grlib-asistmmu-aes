`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6AOt1JjUoydL/syhViTGCCee9ssdE97uxtLQbw9EOth+W6pV1dQKRIzaQsxjY1c7
wOHWOd+ltfQsaEYMPnzgw66Atj1bD+aMvYIFHq2UnL4/UIMsKY995nY9OCWRxu7+
vqXgXWzqswC3evVcore6o0oFv3j/AT7XJtFSeQiIC0N5JvjObRnIhug918VcNM1D
FlcH7tHcvb9fjEV6C9rVr1ckKWLmXG6dzHOTfN4E4RyGnwm+1Ic/QhZlLLJZYmBP
iEjkkZa5gIy2MSZlklPVqKimmmWgNrSH1Iadg0eQ/H2LWGxa8cqV4R6lsP52kFdC
j5Q8nuKrLWIBwwtM5s6Px2fMeADaUfzeyk6RUEIpyV5AFhShICA5K0WlbmjMBzGp
FpJR6KaKThQDd/Hi3N0JZnVBBCErEbdvpgAjhhWrMGD5EPt7nYOEQHt8aGQy3/mR
aiwkQf2qJG/gnkSA4IFo7Tw50HgCuqhJW16Kui6S0oW1SGVbzV73Fc5CNMH34q9S
AmS4pxby/WLLlMVRgdpej0c1YotRicapMXYzWj1VOCNL23ZAKzt0QYEpwHeP6r/S
32o9+DIwkw21kipblbzVeQdIHR8MBw/hQtAL9ZOee8DEy39FLDuaq3070onNUwSt
fQKK8aK5veVH7UGu0a7EjAVefVMg3G4wYHHFNZXOic5TG1C4WDBD79Zx5Tcnny7G
gtrWbmtSSoYUCWQDY5SprGDeh77lLqJWVqF1v2fCojtmhHf+bgA1iOI6baUa/BL7
GsaMvgPl+mm8o9KIuV01lCuJXShUS28Vqt58slGP8dy0qC9joBLysnsmtv2cJmKm
lwj0H/KdJbAxM7DdUuAft+FdMEVTOL+7OzNQrckXb9JTgIcV42IsfzrWZ3cV+vXI
TIej6mViw5nBt4XStr0sCCgRnrHkuFI3//GaDUmSTZyfGolOHEnMYPF6vjlOugaO
RURmJRT0tF5I70ONu9402XixN4rZhOcXp8cO4v/lVIuU/LKyE/CB9lOCk9Xpy2c3
BuHL46cBqOpqhLUkf3h56C65i4w48g4aUnX5j5nTFmw9A42Oit83ikKxhmjSO4cH
VqgRV8G/kxnWryhtA32EntS7fxILIG/Nd0OsgKzgf3zHt0KjWnTl32mAoMCY9hj0
hmO9CzasNO5cuqVcFxpqD3qVfON1xNGHVaBYuxgtfELQJWdZauFKQbuk2Ko84RO4
N01mrswmNQWr7VPyFlXYuerRWSi9SbCDqAt1/7LSb3547rIyPYfk5Np6nZOhGKjH
klf5LF5du2paCUJYRkZmv5ylBDsIIjAt56F01ObZWynfLgDBjAxLsu/BaXF/MeYE
W1I1zxHWaMGEsUoBUCsgevnGQPnKj2vIxyQdqzE4aChHt5QFZ0zL1+weVkyJjCZd
b6hnz2mSD5llbn369F/GGxMux6hrCSW5+R7NssVS6VWcC4PjrVJwurar/y/s1UWu
VsMZh9OIDhx/o4xkNFWSBoTsfPyGHX5TqDkFi35WCLs/GJf+1rwWbR4VXhpVquf/
/npF8xxLbQJlRhvlghmbZ1Rmq1ts7W5jJnYPbvdLmFeQLYJSc/vYgjUUEbtfFTK4
YALzWmpRxLpPl9lYZS48aTBFV5m+CqqyYJD+uUEY7u5mSp4z9LvnZ6GhNB75IPN9
VxFkdXXWtVD5/HTCAb3qDsGKtl675Ewr3M87Ya5hRdBAqJaNxvXgD3bRJQaIZY0s
KSmb8w5wMM9YZdB3mrSga1VlI86He8CCCpeQ8Qt4e1AYe0ZM7RZpd9CzUz9D/56t
oG70I6/XwJkVAbk1Hx6qWwv6jGGT2p3eeenzrtJLAClTCbOLGOa5eE+0N6MxoLTD
7DpOrPI232F2w5G+1T1u/jmF6HmXkLf0aEyPVOHwgvGO0/6hZgUlq7ayFo/DU2XC
mPHMV75IHcsPEqdGcezUdb8sojWacSPqnmQK8zXgHOGR4l7VdHBZu085mfj2Ziea
M/CYthAm/2ARm6xykbJRMBGCSDw8qxHyyPJ+7cXZ9yZFHDOiXK1P/kvQ+1MmB7np
VnrVPTyuwyU7drfBVHQXj7gN5dQ8fAgMXfOoP3PdYnDXK6Ygcew5A0DeVY7UoVoJ
tyA/faifi0q70o7C+yGiM2a1fBlsrgO0ytv/o1ZLdI+o8OGlWaXk3Sdh0VfjN7/M
rDAAo7JwNmEYlx5NDxmDRqwn7j4M5sIo031n9RcmJZjFi/1q0zqIonWmm8We6Iss
Yr3b47kGH3yODdm+Q0H1XyXfUBzatq0klOtk6lyLBCGVVM8CLsz33uAiW5PlTtwP
Fk5hnhCnmwsd3YKMi+FjKSzXSTr/oMLewSTcKofRmCVRMKoQVnr5vjrlEBU0Wi24
g2EC1MjbgVAfl2A0mWIy/9oRBTRhtn6ahGAmOFHG+Pc4uZCCzrnWwtjq4wP5oMnL
YX3Pj8X2ykF8XLKg5z6nEV+is6k+rrz4kuLIONbm2LdQho3gad6/u+aY7Db7SH3k
`protect END_PROTECTED
