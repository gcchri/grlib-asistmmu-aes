`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wAiQjaLYnWxy/HzuZxod3w/9W8C8nnyRfWWouDzEWeKdBhDkfH4smy/NRX5WLq3I
FGol5QHZ+j6Re/ZOPYOqfBU1L+cKc+DR2yZsveKpTfVDO9goJU52JXArJbzThVVR
sdSBpsmhZGNnkyLXvWN1KqyrHqCv6uGDZRtYcTrwQ99veYIE+zOF/rAo8T0GLd8R
ya+GilX3lQwhU3h41lSHmoqp8mUdcceeYazqx64QCSS8wNIyDnrgCvPHGy5fJ8LB
M8thT3Mb/4QyDPUDzysh+2kl6UprJ6gOjW5yWQWJOqE=
`protect END_PROTECTED
