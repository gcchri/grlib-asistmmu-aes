`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvbbdnUWdmTnb/gSuj1RFgBfZ8QFU2UeupnvZ9FtnREZgvzxe0ptE7/Nd3WP4J/L
qk7Yui7+Ky1990ua77LS9unjrCnJuFn4+YsQzsrKkVpj+rAWCHfJTNARQ2a5p+Eo
te4uyDofabK+v7z3SUoN/ZkV4Xw+dQiEPJN27vygaMBAw5RL0KPmTciT6hhF/w3Z
xAGjTxtk3yjRPlztosLMmTMG2qWrhjRwzPUQt9hmrRTT9ezO3bc7069OLU/s6XLC
UNNF12USAszVk0c5AG3Vh2LCx0VnLLij1/W5fbCuhiv9FULugDK4LndixQs4rTYj
HDWEY7vPLmbANT1ivWgpBIrL8BpdAL1mVKBuwGxZQVJx8hpw6dNH7UsIPc4HAKBi
lIqqKb5n3f3fezexpKuBvVuu4N9lilxGpRRy0Z8RrgFNJ3Cc+ON103aNTrz0RH6e
eWdRda80LhKT1cfIWjk0PL5r6mKxXtM5LumpT2UC8y1e9m8UlwTC5/35/mpajtfC
QZNbqjDmFjZzfRucPpHOLMgdJf/jVmFK2H31c4WhD/YnPjdAoSVnEn+jtpkYviVS
lWUDBrxsyQhv9ZfWdNV/MQi9j4ylqcP6Q1fihRAp5WHg5AA/aed7iaS0/r9DVHGB
Z/TRyl4vQ3oalooUy4hlGiHOyuCoXypbuX/REGQXqHdOR5Jt0+J50zBJpaLMC9yy
JvLh4rDUdpwhVsIEoEqWIJ5OoMLTWCSv4jQzksdEevMI8JU3d0PVoYmRrUTy3d7d
bOddZLYJQbrUvLqQ/TgL7Iwux55DNIaDyruv3OFkLhDb+0Usle6JOlgACPWpLmsv
bqIA/wYVjImAHzEb5gzR5oFiQeHxaN78okVc+GSWTwVocIOMjHcu/tr4/E2oeaGm
n4VuE+lguauG/q4dWOwLbkIMN3S8BZ2nu8w9CQ3bUB9/sREyeDISM1Gyj5Yx9H36
JH1lbajJld9Og1gsUM051jCdMBEYzBQv6dgD8yUsAfwW3lc9eNabEIc5dj20s9pF
qRvDNTJ7HuCzpPkp54dme0e7tFPpU83sUgvBRKZVdQU5K2AW3cTmch921z3xOAYh
Uw8kUpgad3ek1Gei8rRhuxH90T9J0pZr98e5nXyaOwvSwBBsVaIkacY4ABvolMSj
4hcqFo8rxb7Ga0TiyVHRp91b1hCMseJdoEvLonWOZArY8p5uCLc1xILzp3A2D30y
es64EQ+qG1r+3GjwQo68XOwCByl6vPXCT8HNmKhosyt6M4xLGOIDTKbkWWhGKi7u
4XYhtFYyvPHhxWQEZ8NHO1j+YCyW+JeKNverZ5UYUZn3E/jVaUQG3ClrI3+wD55u
KWISQrUdKvCmS1ISFjzDV3Kx6NRz0G6A65YjJLG25tiVOYdoTwRKM6pMPtvI+vaW
ZVYDj9WPT8Wasx+UwJbfxMC6Daj4ez2xfkvwAarU9Gq9VTCnHbd5DsxsPWKfX++T
qv4kkbKhM87axRIy7O3uIhbhOjyVi+SpSvqDfnT73gJtptyMzDNT4YhPZyhgW8Lu
jm5x5+REdEtNQ/rGjqWPC5raoTgKqwEHIirEBO//+Qn8UmH01RK1QPa+/gfczZRD
+u0uYEfSXNL/7go2WXUNFbj33LX8Sb7Sc3aD2b/lJum2j3+NdlZh4E0X/mTq5JmW
2lvzlB062eZ5/3BdAaFJuFo18U8pGhv0dB5GwEOhbHFY/S9ufn4tnEbo3MVx2duZ
Sr9F5Wpsv5QjtjA2hWJU2T2wxUFxskmx09ANimPoOBDPDhXS0ZsxcHoTTrCltzgR
E03/m876IXegJT9Vn64kr9pakv6gOTq7YgXlC+W6vfX+iJqldoW9GDpU0z7vyWr+
pRIz6Vx22V3OY8HF9R9jAIn//sWoshLDOOzh5ZSiO9Hb/VVRt3YMdq279QtfN5VD
bEJR0zWp9xBpiZcjbOKyUT4QXSq3HGkhCsJPGX+QSKmZDhkOYIXmLEPWydEvhZk1
vOn1kqOyBu2pe9QWsqhlqZXmWkL4n/marZifiadxTBGtA0Byduu9IDvd/8MxJJ+x
4fvLx/8aaHcKI593dceCftSndX5HbtCu7wssUBYDt5nC7hRRHq8eGIA6WrkcYoTg
hQEaOR76yT0tD9oP/zitL24eL/LPrnSkWE6uYXyeaTPZnLgVE5zrpENsOqtHJjZS
wiFPjtyXm543JLxdMix1GbOK8o1x9lSm4l8fJoggiIsfQn3MiPC8SU8EWeOSsLvG
HA8KiczGf5Jzfdbl1Hmlt4FkL5GbpmqmjdWIuYrqHpm7spYnl50JwcrjNIVwnIRj
cxDQS+6Dmwh2O0yjLLledaBqtkE15pzsPGvvRjy7yT71mYD4hYUbZMVBav3BzuVf
uo8rrzqfRseSAtsDLPladrtUJOS1LvPfvumvkuqU/cy25NWk8QKI2KHPJ4Wni9g6
y5xKwdkGTvUy7I3jWxpPq4+xTytVqSC9RjaDD29HAGkyXdr2fdtOYVsMWdnj1eEA
QvWl6zwV6XkZf9dmU7ieFUFzFMAPTUkTivaw2sUUPmEq/BuR4nMwfO/Cq2UPnAyR
hWiauy+kfRV5yDF8UszSwwABKGZv0vx66N9Wz5BalMwfU3M63NLfsch1F6sxDeip
MknqIeEbOjBBSm/vTIRRifPo2D+aYvvdBPa+qhas9RsdbM9LNbyHBlD2QxdcNeaP
5KZRpO5eMFo65nkNUeORZ3qRLEzCgykimCnbjo4I+YRs9vUdcBU7F5CNNfc9u6an
oLfm1v0mr7guVtXF2onm9tpTXresFSWcnh0DiB4lXMZewWz95/f//t7a+BStZi+r
ru/RNgwlto7FoONHpyKfqrd7ibxl33HBwf6IcovBhxHjESvOgVxgrAKIk7INtI97
4EkC4UMADTyeLMm4buIEisuBeKkPg/UOyK98ivCXiXfWZBikhtf0p147c4adC+jq
uf59sgLu37HjuPzXztZMseRifcpCqiUx4Cq7u3DTJT3Aj8gVfvdxcxjMh/LobLu7
mOGs5L0pnm8NSgldkdH0Cw/cW3jQCRUhYV7h74UlMgBVlhiYbg5KCB4AYib3IT/y
2xujBIL5PvO06PLa05z8prHIkJUcabvDklHTkKVtPuH23AYQI63PDzH5COey7igU
PECJy5g2u5/eUDRGRM/nLfast2BEeIZxYuBGIlo/0H9ONrFcJqUwrmatNWKoaW98
tmWVTYxCxZVrn5m67i1L2VPVUsPPTEfAKj/22fBFDLmfwy6B2S0aCLKfO6NoUvue
4B27l2NswMhIsWsdHxRijomUyFXDNXLxhVNIIX7ko+t1LooQiCDm6b51OGRKwCuL
SU0bhQXyLMi+ltwInj1Ag8TLohqSlkpB7YyZDdc9N3TQxjPFvCpy38U2mdIkJQTY
uazReO+RqIqCc/zAVi7yhY5WnfCjh8rP40JKmH/OAxNJLJIRoUMHo5/ljgaK4NRs
c4VjWZN6mtNLp+ZYHpVM/7KkSE7fdOJZanCH3y8RcHGG1a8N9fE856ihUYRe5i/S
M756K0kUVJlxh6gkx0O6pbexy2Oi6G8mdKqHkl/zIFHENNnTcTvGdDN2dt298Rsj
YEgM6/iq2eaYQnCPoiJ7w8XPT9tFqlTMLtfuDYNsQUI=
`protect END_PROTECTED
