`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lWx2LMs6QpGJL9RTktvae3I4om+z13t/8X8uYuNIkm6zJcLyMT3BmLY/lLbxRLT8
jFnjsbfSsxo2HmmL0Fnpyp/5XV31ec9HX3HsEVpSOWlCInmGr55JMs0Ojngyfa6y
X+LBQMO5EGvGfMajaPqTg7kllQ4WY6FrlXiwYqx8vqRxHMSKFyoB0F9AvzUSMhcQ
FYYqMK2r9LfGjTvnEAhtB6LbkYF3/xL5/w2PSM+gv4ADwJqARsjh6tMuKk1JDnNW
xJaQblhDHiyZ/Zv8zkuTjOUh73YblXJ7610BI1702XoRRqHhiN5OoWk8DSDxEPYb
26LKYCGXS6JjONVG4xkSmwnlhvEcgeSigVJMEU1p/dzPSHeLVxNj9y9OxAQximCk
JX+A3TPGUPEZZez4aNwjrj1WiEjyGmUU1mrTXMnrL8v/B5ZuHWOITI4K3JHDUB6I
npJmHfs8DwLFfeMnX9meDBPKG9BtkVCiqc76R/E/2DE33WmFUriRlfeQZ0vvzga2
gY0H/J4INExAL7lL4p01fZf0NBkTQO3ut3xHkJQfw5hPpadWzP4JcHnPSQRHyrf2
`protect END_PROTECTED
