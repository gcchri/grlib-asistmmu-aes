`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AUkEIN7kcG7ET8sFJpJdKj5QtoCLRKhffvWq6bGS7ar/q/cWxe4tVGTI3VWBkPXP
pqEFR/uHkZvdwpXolr1tkNzxv+59PhR2wMPAFVyZT6fPmLfRHnNFldrIJjY3l1U0
xy7yMfl7rtMjeYZO3cR8DUOOaHoPdhch7Jko2WwsROpjWOaN5yfKIYzkiAAsDl12
bk6qzQTDh1Dol1k0e4DGrw==
`protect END_PROTECTED
