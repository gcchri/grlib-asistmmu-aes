`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3UZ8l08Gewp3pxTm/axk9ArPgZ+LqWnSSPYOxRGEv9o5lBx9eZMEIcRy09XTzVO
ZKyQyIRnfMUr+Monb2LBjHQHQlggA8Bm3QOPYCDam1PnnVjzreSU806p/bmzlZId
fg2yfriqhG4PkCf7CBfLO1OCIK4gMcWHyWjkeUZNtowzw4ZzcOOcnpbfttx5IoLQ
9p8ftxuE6aWXl1ub+4MaKuaIw2b6iLqhGC34NDf15DV2wMWaoQK+0wJjKpqxaSvb
1EsbHT7gqoKkpeV0uu43p5XIrtEVDtnBkF6Lt3KDGUk8DlX/I6NxOGuXDql3WoE6
TUpR9cV7PcekyWRPWAtPK8G9dU8bZK2xJp4DGiwa4fc+GaNx79Tx8+GDLxNFMHRw
9bFFPtfmlfa1/npcVt+d9kcRr+EVj71oayPSCAcY5Ch0sO7dmup/5Qf9aUpg89Nx
bZgROpS9YK/EYaT8klqE2d5IV4qj9uPBmuoeFUrE+QaNp5e4LIA+TniQXSeJfNsN
`protect END_PROTECTED
