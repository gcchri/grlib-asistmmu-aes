`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wXQC9qvgrzpB1g3A3ZJjdc/nimbHxxy80tSCzil/utWNQQEsTRFfSytK5qQYRukO
S1SsG8JUq36LIsjlBko3I79j+QQxwjHqHT+3wEaiJLIEV0SzxqQZGwJ49oU17mZT
RFEY65YqVhsGgCaISVx1w4X+lSqNUkVQTTd+JlSFlL8qZ3x6PeN7VB04YEthBO1p
6+JIK2cb8nut/c4yEL2xOCHvMvQla0Jy/Hfi8pATy0H7KpY6AeNAX4LT3AMlVa7U
XLj/Ldp5pcw2morisHFo8jWGStfqD+uZ+tWLNuRNn8tIs6JrOZJivboP+YUYDA9E
2Wswsoa98Mbcem0aYFq1Y6WS5q7XIOr4AN1vIPpCYzwyYx0wf4i8fQWdYY2mIU2V
oPr9Y7xTV+Flz492Ew2n+K3XVeFhJObitrbD3LM/A7AzOCIk1a9oxN+t8gKQ+/9T
QNhice+oynFchyPvckN16z9yJJPmc2YsbDqd+rah56QHp70ncElJtQ1ee1mrdYu9
W/EpwwNnzXll5B3jV0TEQYH0qMDJe8hT0g4a2O4O5FU=
`protect END_PROTECTED
