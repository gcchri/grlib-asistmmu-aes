`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LIG9gTHFiLbaL+mkvozKk0xPtA6TSVbWwST5BLJlYpZiL023HVmi4gv195hMoM5l
aYqXE+MQXWsgWOHJOisIPhibHZvstnixgPAqCF24h5FT1guJXFkdZOD+kJsNJNce
Fuj+6zdnIGdE3hfA8vbrl77d/8Ol1bmt5AAISp1rxHTEy6Oh5fu6un3I7QDgvFxa
q9krJpmpJ6qVVS3uV8TVgjxERYkDgxLQIRhTijX+r9u4SX7GCIfPKPeHNnQAhj0/
XLdzusJZJJVkkpKzyMfedljW+kIA0nshFubmlnae1OJkxvu1Slu6ABwH5JNno2kF
9rTNsZthxWfBApX9z9bFyNxuDDSWEBc4pl+afvNVmtTEOpl/cRmlAPTvVALv72gu
QCbkKwfkQD0qGOGdNrp7Wa2N1qU5QTbIkj+nGIhni45G60wW+YohuFVgnWh7VRCU
5LQ/XmngJ1tNfs94A+AUrAYhuwjU6rQ7hnc6+UOdeJorRP3DPKjfJLmfyeWbdcYr
`protect END_PROTECTED
