`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tqwz/8S9ZnCLn6F2bbS/PdHEHjIwP2QcOTufexW6QjRHABXDOnjZvUSmeKfg1TGA
INlsQNmvO5gf6yWtIUl3PNsWpm3eG1DTnfI5jlH6e0EiVfEbWywigmQ6LEeFQFsW
fUTlBauU9lH5jlVkfW4sQSUyvYJWdIAXMxrNDpcGTXvVExybV4rCnQgxsYze+y2y
6QwZoJShicCxDoKfcxsuF5XH78/v7hOhs9JG1Y2ZVYeDRtnZTXFjsarRXGi6xnJ9
X7auBMgLoL/xx0x9CKWo8RTbbZ9JVlJFpZw2ocNnQT1dE8uEIqQCIQn2hLkPYx6J
aTF9EIraZ/nwITmJPTrm9fB+kWQTxtKeA1J18rHjQsQ4GhrfRAgOptWLryLN8bcf
ef7OBA+2zH7p/7RQ00J/7134I5yRc/HiLmSYjAIthRQa2+cshBj5RUWn5vFhvotR
V/XgxuFM7c+vSvMem7kKng+rAdx5Xbvd3UDApwVx7b0U8IuphNYHJ5Yz9lRxxN0r
KNqk0wyVReDcnMl95b8dnJy2vKkL2Tg4c6yTJ7Hk0+ozu1IgKpk+5+LgHZcMXohp
zX++3c5jY3cTIrFBE5+5St1hO16aWFZcBSxDLKzKCWg=
`protect END_PROTECTED
