`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b3zrfko/lA/LamZUpJv/jfqy14/PCCwAz5nZHoNyNZ5+ymoJR6E/jMFMLHtZF5Gg
deRwIvCc+mkhZmDa6kYmv2k6mBww/zTwAT1m+xoR2+myyYHUugwBxdBt1pRW/xvv
Ino2tBGO9ql1BPeFqabSxCFEFyWllyzeFs+VW3mc4SZE6a7nS+EbDx/dZptNiajY
oKH7PYbrJS2JcQTdkey3/Lvyagdo6BuxXIb2GXcSnjAVMglm+cnaLwx91CKEVM2K
mWoGEo85hdR65jQS/PKNO+TT7vpR93oOijnvjV5nY1IonVwEVa6lv61gG9rPjN7g
CK5g5g6UiryFyLUUa+ySRtGtO+2ELeOKHkLRTkhUfM3UAQYTUfe3F/d5/juZ1in9
XMG1sCKkLPmcEGEdhOGH4V462VaI4CuFn+UneqKRGs4yXsYgCZWG9mr9br2EgUnF
HCiAnLg9LgKmQtuCMmTBufbAIdO4hgrPqUA4RhkfiW5EH9PpUBe3B7RubpFuYhwJ
gRQW4jiZFJROTIdsmoYqhH+osmQVOX1EblwUmhCJXoc6Jud/JyiW5c4rCghlr+ob
Sq8iDNNgRMnNCzQ4K5eMQQID9aOsfs++ExDt8dVkqWg5UOoEuHlx7cent3GOEyGQ
78FpHhHZinEQXIRwLcLipRhxooSmRKVd7wdFrhr/diXZpqCWlbEZp0NwldnnpZ0U
jt52jUWMkim9DsZFOohXWt+wrtJgZFZkyDorjyumvzJC6pyLEcRa7Y590SRa5uOQ
4h4pdrvhmgWU7SF5D5ZXiNf+9oxXLnhmhr0J7f2OHM8HlRAcBLvSNmsTV7QmvPqr
LKxe4JFyKbPlF/8OkNakTSMig0N+qV/2EfRh62iFUR8YIy4ti1AhgOjqdbzr/q0A
5AaJ4cECh9uGtkjUPH5/Pw==
`protect END_PROTECTED
