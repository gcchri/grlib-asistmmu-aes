`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1cFwE2znlPq2NqKy+r2xrrpoN6gkMsdGVC46veQpNh3G06xnFiSfmBO98iqDche
Wltjx69xpV+wdjOvEf76gca1vFiBvmbwyPzuJp+R55v0JlGNNFfiy5BsKZQUc3x9
AE5Bgq/L67DpD4KKPwLm73cPQlz0EG4C5idPTeZKCbgFExnQcXo2N2dDTajEOxak
ZNwEd9imIUg0EiOdBqdZRLPEBvznaFuLVtSFIdGfQO6meoWBt9YUcF0GmORL211w
xg3pjHJtdHCRK5yixY2zGiwdYsr9H1dsdU6SKmI+K663QNboD6Tpd8FpLDQk4KwI
WmQ4jBf45OpjGsSLZ9boOncQiW+NvbDvHKUkz9QVhwDTQRd7DqlQA9Yr0ycRfEIg
KucuFk0709Jd8m+78s9NBJzreSCvmcGIEBoPQ1jG4NCoXTpdzF78uyJxhslWeoJ7
WoqyHPXfY7553GIdkWeoT5GfPDLeiSAUeDONOBhqPUdY5eWuBQ0qIkw/4RIywkjn
`protect END_PROTECTED
