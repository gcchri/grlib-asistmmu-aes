`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWYw4LbVDvhh0fxQRddAvTwFJd5YWbKYKMZvOaAI9qufrLUu7xGkumcLtRf/A0+j
EQTllVVENTNbOyJJtfzTNrlv45tlBe4KcN73iwDmc9POtyiYngURBiAIWAhO40wu
mAfRDb+iNZzbXEkWe/jX+HUdBE6RyMkybjG9CNfS6OsWtxjrNkxLVo5aNWp1EY90
gbecCdbW9D795NkMMfOc9F+BHYoBsMIyFNDbiTwgArfp7IEGCG9NkdTti76JR8wN
yPmmfOP2YQ+xkSs+8s3Pr2feXIU9IG8ejlOGb2B0xolO6k4vvVbnApOTYtVNrdDG
9yMRBLQ4NNfTJEx+hr3EQd+4bCdxSCMGvgl75ewwPAHNudHHagTVpwYe2/l67Yom
0jcqCVHBM0gYMVH+MqcWnIEp7FF0d5kq3MdpSoxlItg3FKsWuNXCQb7sBMlLcvWu
mjJY6L1oRPnAB2rEHxcvKB0VbdHhYhlIoySOgU89yf/mbGj0sD810K9F70aEjhNZ
`protect END_PROTECTED
