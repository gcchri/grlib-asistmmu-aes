`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JDLbymqNUg5tzyQI2Rh/9mYHK8qMnaKGTpqQAK78xCATKE67YHSoEM6GqA+F0fDY
WFjwNcyTPcH1XgWd82iSjjS7SEvldue4DYmIYPLB2QC7maoMTaVLIlk7+ehhcpR3
3khwBwW13DatvgWGh7X1lS+f/V8Sjf6F0vnyt1jvVUM0FB2SCnqQOpMX5N45wqeH
dDQag3QuJ4aYGANl88G4E3Gy4xJJRXnUPlj/rwEHBugJsdsX/hQVR/BXsqQbdxmR
T7pG+DZxd6TROugIKGQlDiVlZrbGKJelbrQ3lZuUdeON36zEa9pGm22uNDKf5/Ut
HjAEXLZId/BvGslJYftTkSCfnlJ2kd0whR1Zt09CaFw0clED1bi0aY+2ZLWNLqeP
X433Zy0efF1UHdWKp5oeUguvRshhgw6gL0LlkydIpYU=
`protect END_PROTECTED
