`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vgZoHeulpjWHKo3V84mju3mMTTjD8zXck+Nfng5/VRCxEAk870gtQuXENoM0pMC1
TrjIOEx1em9u/O6+qECc58ZFyaPdo3RA3JTc6ib9wD2U83RT96e2YU0b0if1Xafx
HGoAwfsjXlo7vnQpMvBVe/lF8KZL9kuJD9YavHqgSPfaEgre4bqGrQOrgVmlxp4a
ei4klGYBgU7cYWFsu5hnV8ko511Wn6PCRHCLJVuk0tgKGGq4Tc7bJT29KAOpm7Nv
qc3IfdfAj0Sf0lyoE8eSHI3Aqlb99ePE5bdZv3K6DeZixmRmp6I2Z5O1fmhumjGZ
+j6yurAk7snTtMp+uzH11I8v/7MemCB+hAryEV43hIxG2hjr9wVmDB7IprrGCvJP
6kSyvaVfgIJHTK40HI/Mtasd4PQ8MAQfZggrYbdkZosGWCHa9aQ/lB8pPzvVUtNW
OZbYNQoHpqICi65HvAVb9QmUiswh8fnhURnKQw3ykFUml2x2/86chxZjb1QtPaQZ
OB+ABN1+7heBDAUfjtpsYmK+EO5nqeyuWanh2v9F5BGTPB5cu8jfVJTl+oPi9YsR
Hsio7F04GTSuks3H2p9m1+HiOJFZIBRDuxbTBhxjucxewsLl0NfRmiZoYGCSzgUS
Fxqq2w9P72MaNyO79+aXb+PIOAeXOIGfBuD3ZeEQQBrNaykGXmL+Yz+AkTRoyk31
SAlvLT4wYVMVauIi5MHcV0RyLKiaBfPrIZFb3y+7BFIQDso8IPoTwcbTcU8E6N8I
f+GR7AVf6ImZttGN0NqkVM28Dq7dTa/gI4lx2pjx0rcpXOqP4NYJbTHh8FIczP7L
dv3qsk27yWNGJUZyglKe4/r6wkHWTOZILOZa7QVqOeoZQBuXp4G2+XV3AayJCqEK
tRih3R5skheoQtdm8gUq0MT0C3MDVY6zjC8N7S+6F4MtKFbRtLuhrj9fGKTdKKLy
4/I9du05yuVvygNIFQ6/oo5m9SmKebEX5gwQ4d8ZImc2iRGFsOxWzy2CXldGD7uT
0YfpT1y5qHByoOzB6ue2Uv/ZSVaruTXK5oxKtnWDRHrfaaCC3FtVmgt4L7IyngdJ
EB4gAky6+k4mJ/jk3tAzJQ1lNjfCAv83j04WBo7hVgqClmT3jSpDJmOavjwn/RBH
VoF5770Hmvs/P4r90Fk2NS71XTj9dAcScsCiGiiwv46o0L8HLqPSPSyIFRwzW+tU
cZdwnWw3G5SoxXtDy5XS/rIKXPEIQN9Xse8VcLaEec/zl0dASPZLaxcInPaXD8CZ
QR+/rsCLTprfymt1G2DselUfpUBT0N7NMEijBtHcpGyGH0LBdMo9FRTD08dcd3ca
gRyffSwQEc5hF5eWS7NmJ8s07CcLLggP+qv/mPj+yuxumREb2JJ/bEAvfaKzbQTJ
FJzcNS4lue8sTcQGqYvwLzNWFQaHQtTuFI+PKE0l7iceIsl17ISIymk8W1TLSKDW
tveo6ckTd6BGLGbSpUJOsmxXm5Rh7awumr0lXkeCfZRk1v60/GYFMsRwm0xa9f16
BYKylXL68UElllTyNhVUNKy1imXzy8YNuG4+AaqKI0u1QDwoXqkfKo8h9tIYr9Zw
TDKwSjRCwy+X5RjmvPYq1DXM2M2i5Xd9+oknvjbjEYVTAUbUb+QnZ49Rkjl8rMtm
AN3iiZnydQvnPnporcxl0T4cquIFSPb8muOWI9ocEq33SRswVvd5BtE3f7/sm8SU
SZmcqu835ye+lJiy4PWvGKRuAt6Mz8PqY0aFc1TRjZrmwn6NscQPx3CDX/tKsbHS
cp+sNEUVlq4yQ5wMDBPO8jU05AuO4IaJUE001X+Ka4k/axdJf2MaeB9KYOcSb/KR
cTiyRWEODnbZFI3Ptu36ESnepWrBVTXUCYkqztYr+jogNGPbXFb1ujnMPuNWaXLi
6tRDvoi8AV3hSgPsKfQtjzwC4fdRXcvqPHMYKD4CchakG/EKcjsCmLs8g32enkR7
3FUdgfDPdtyorB6uFN+8p68M64zSYxWIRaGQ46lp+4Rfk+kl4UDUyAVhCnFL97JY
o13llq/nZ15iMIMdPj1q4Wwad61Sgk9BIjDFIjCB98QFzr0yrxfGnbA4WdzqWXXG
CMCLb2C8z9Q01eBLOYdoXprWlO/byN+E5wJ5JJIbksl0HWsA/CqGZtH+n90gK1yo
SjaVSkqqYnfFnhrbRADuRdRyOs3I2a/eMWoWgOlSl27SfEOsRW1Ly6453Ax14cGn
2oDq1ZtcePb+LExnAarobUeyZVVDR5UD+Xab2/otbVlWQ8w93HjlfS+IUj++4OHF
EedW03LN1FD4UrAdGxS3w9wbk2MqcvzHxRjwLnAmi6mREgA9rkmT9Fl+nKxv04/d
35SCv1GnMqeygWHIZLOOZ4y+n0cKMYJx6p0/AjBoeIrrz2SYfYJVym+/QL+SOFfY
m5Sr5gJKAJi0kd6Gz2jxRQs7nabN1IehybYLWAzrmWSxtUa5XyYbcaICyfy6gmD/
/VwXjtTFS3yJgO2wEUwYn5snIMRdxEjt/hcicc+BXWz9NUCD4j3cY26rN+jikoIL
Xnb11Ul3OzQAdfr/ok0L7ZtzH90Wjtb+rsXTxHl6gue3SMqwi7ZiIbVG+APTtipY
IxektdbJD5UNRYFZZ8DJL2/QEVSQwjmOyVOmnJiRZc9quDXtswHD+K42m1KVd6ug
BS0onU82eUg1fGnq/ecE7UcgiW7KPSYLp/CeOxCQIpAVfqEpV8TBMSj/qxu46syO
oMw/iObcY6k5E4VQQxhLDNHGCVlDxN2j4fnOVHowXShuU0Mu5um3JjgAyx1xOCQU
3QI0Kybdi3h4RCPC+8POelzITEzw3zBIxcLLqMj6mzMToMGOC+lH1Ly4d3ahtjaU
LCnrTS2sJTFEZr/bhhxMKOAzYI5v5DkqTRrARDd5T0MKh3TeCvXSip5yWV3RZWhs
pZkGuBewgrYYEZX3jMI4qCC6wBgC+1r6phUCWk9PBzCYe+lj5FT03o9aA6WM/GvP
Jz8Pc734f4KS8EGVvuV1Xo1iyYhhOxcbHNBmJ/1lO2qUo7/Eub8vGh6Uskt/J6bh
uMp7YtXISOojp9VQJwxHOEznaXOqL7HDweImT0z/JSIdZONVJt8uNq/O+AAbtKYQ
kKNSxO7sC8cGY0t3u3ljzVv5qqQhZ20pKTseLXPwlMRURoIGsJkK1UWP6qHkqL3i
F+4P4BzdKqvR3gbnPuxAug71DQSHg9CV2FXL1Uxi1+M6nhLkzLHDjshHhxTPjPAw
3Lear3jl2lKJ/fBULF0fO3aw6warlGizHkqNFcE8L6YPZvI9Gclu43DhYVImigBu
GhvmnXw4azpHo/koOP2T/mmuJL6lHhrvi/DJs1CoQeFFmShCE5uGRlA8wxXNoV7S
57+j21afjWwvgenPy5gAP1mEPOEC6C1uFabUf7EMpCOJKLfRsOEOcZvl0jeus852
akOe8Z2ck7aM9XVfjolzx5XEJdKOvsu5BO1f3jn01y1Kr1XHa0eR5c+Ic1NZyjc8
vu5kNAdc+ZzoYRGwDdMTh4FAaMTDlp5dDJlrKkhki8Cj2SHgu+KbiZXoFy2t857q
p74hSObb+ZgyZ2iidmVUC/GWdRqahrLRmqgKswzA7yC2q5xnzexHp6JqfJD2rZwz
hyMthx7AuM3iGu5N4imBerHauMw+D8y7arO9Qe//FUnQMK0m2uspJDYsYJeVdtnz
Dywg1PDSwSWsAnC13xEfA4uC2PcwRgS3FjH0S8NAa7zFzMATDh89/Wd5C3avgN2y
pCQl2QfmZ5g+sB+Z08jc/GMwpADNQcLuVXeJLxojm+yuapy7otAYC3HE9L9FBEpJ
0J+5lc5AZv2lQDPWcD8r+n5+l8BKqNUlXf3UV62MND/zWgE2B9aoWHc4KUmxEKKu
TQSgCy6wnuOp25WRXFI7oMxsO5YzZuFYaOn8Y9ETlyKUYgiU1+jo4Qh2CZRd5hdx
fdc+fA5/GNcj2+P9ax5w2V4bpVZBZNfHAn+MgiOQgYI+FJ/of6evOExvoW3ZHL5w
hPZFXgI7TVXlbuMqQJN29wKpIuYzZuFyvCFoWLihhRw1uXZZbzV+nHqrOaj8XACz
k8rSSWIOWrO8ilrd8Ad+kkoq/ADl5izceKFcBEH5eOvucLE0hsr24kMkwQNomtKm
M7BjRIGSN5htphOdwS7sHw==
`protect END_PROTECTED
