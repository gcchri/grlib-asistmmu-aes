`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v8ePZvO136M+u+ZiXN+vmNC7vfNSgjO60iBSnwcXUBkIMqr9KOrdev+xKBYWdSET
MM7my9i3LzsKQ5PQJDwjVEetNcxSA3AZPpnj2xGe7UizsrZb9KT76dBhxcaa3m48
cqUAoPeyEvqwaZbX5wqUJhJtZlkdSCDgz2CwjqMSnrZZewYxdaa4hMOUZMphcZiV
k1RvJzeCmVBKV+5Y1n9ouo/v3XpeWxv71yvJ88AZdoMLEPkUbo8+e/Fr65cfZ7Ei
vUspnv64CJUA/9o1tpYWzhanMycPUJPR4BWbEBafEVwcnUuaF0m9RaHhcwrbn9M3
7N/mPWXEkOF+Y3BOCNFzr5JcLFjgoTYtb2OHzjU207O/DqLFJJvGbk9+Me7wHlxK
`protect END_PROTECTED
