`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LcjBIyMtfEqIK4n85sCd3a3/d2gy5E2OU+sWgzKpf23XBeo6PQ1vGjQW++1ADJwd
THasjm2bUoNZT/IlvP+a7RB6/ClIgvEDwZjDP5LQzRHlFsfBpTkiwc+N8kC+47Ci
kkk8HUUbEF8CJjJNdkrCLyMfNrY6MuGPBOXQGsuaGINgTBn+9ocL02GQh/RPA8GR
5qTkQzJkllc7TVMlsJtOdLhbRTj0XxzF9bUutwMbVMJLEijjXuGExqu3rTnIEoN9
SwAebJ5ZAYsu7/z4QEDEOKb5awZZmxTIb7qHZhL36ffB+ZlDMYU8wmu56ScK2Hs5
iD6aFWCAlgxDa/u1Jy9htKtXANZzpDFPuQwCPOvDuge9FzNU9GO+B0Zb+SXPamNP
KzyN57R+XAwfa5X0TsP4o0c4F4xSHXlIcCX3/ByVTyWVOMdpxzpHAAiCshbEZc9v
uQPLTHouiwarwHGXqzX+lhezr9bIQQkYQL4NyUu9SOk=
`protect END_PROTECTED
