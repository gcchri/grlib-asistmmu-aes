`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IKVMcgR0XrQAj9qshyU1mH9NAWynCLfl+ZEMulMGEIk5y6qhRsDw4JZgGaGIughh
em5uTxTUMW4sSqMBlnRqqFXtJj+ARLMGSBopdAC4GoFQiuJ/l/3Dxj8jMUFprKES
kk6iOyKZMygccsLBPd5S8YvELNUgg96sjNS0Bfu3zmuBYevUiDAdju61AWWnIdd9
xXnYtbCxtkzq1md8eOqRHStGqnjvoX++xrAKAaQPulXOPMn9Wy0yTfkCTg+ydT6e
8BPIfOrXVBJymTFMp2kED+oJS2ZkQaTUp0TEw7T2pJhykCt3/jI7nTnd6+7HldMm
MzMhE4LfnCNEeUutvv2TWLwxUzDUPfS0fnQOBOoDLwxQ5IH/Wq5/dtigG/vbYVGL
9E11Ms6MGY1dDZSQmEkA5R0P9LeKF07ZENpPgSJ+I9gVyOOmb10802brNUreM8ho
OPcHwt50A+I9o2RFkVgkJU9P5ywuvaX8ithQRcJ8ZFgzBYyM3D/Z5EBuNkkUCJ8Z
`protect END_PROTECTED
