`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XLh4xlxyjFiTBdfsJvKg/50OffqxtPowDM/WlSlYB4I0dg1IFjokx8TvJ19eSM2C
8uXKSZUaTXfhgtc5cfjylFZHZzWaMxy/J6ypVDxtjfN4ror3bycsbUZcLok+jHuN
BAAznuIRM4T033AvdERSogArBR1JDk3TRO9CjXm8ekyGiGgrfAVbIEfWLM5D1SH9
gyih2Otr2A4uuSl3HDC2aTPS6YoXFlgrKI7W8NNBLHriF7y5GsG/on2w5NQGuxys
7DjbG52YMz5cB5O542Sbb1cEx4Byo2oUBCquhMtAoH4XE7fyQvHDnA/paZU8ShEO
TN2jYipi8qGdJvOf3+MIKllFoq3yEVlTNJd3FGEfJAtU+4ZW5B2G4yFjQ8Ls1x88
/VQRjQ/BoU2my87rt1MS861pc9Wk0UAKLKWtrExkPc5/b8g8+hwRvkKwsC6/IP20
JQHXFVLhpk6PPD5WnpyxCIZVqDLGuaG851lM3tE9+A4ZERFtkArCUkfWOa2X/67b
vapbbJXVapJw6DM8NggUkf9qZ0bSvUVb2NaCPsQFMYr1cykIIhds9vjfgQ0CagY5
rMpjWu0t8uaaA6Bow6iXQAnar6RP8i1b9WdF5eAm7PMPJRDONhZsqoAJnaa7Q2Az
2GRZjE4OPBhmEI8hSkbnOUJ6GDdSVFUYPrpEhP6A/NSlclIElEbsA85Px05e6Jbb
RG0OuWoFRjBQ58GvZycVP9yxdokXxmxyawZhCA2MY/XB6KR0EvXpIEGzVRmRNm86
ZXHSxzJLQZGrkzC1Ja5Y7BAfIqOM8qrfLN0eHda8aX7uQRh1vXY0xSCE1pfupCYu
uXQEs1SolEyK99vI6dkH26uH7GA1QLb1sbOawU8avHYHFaJNouwTe/rDySh1hNqZ
1WCGbcAnXVkqbQCrxaRDvhsmgl4Tt+hc11kwpPZdQe3WhZyiU2Yuf9cr1zdl1We3
VSM4Vp65MJp0CE3nan69ipaLMImtx1+7bXkl7K1ymHrjMgEc3sOn78pKuB913d4/
2GbsYp4U1rL2E3luJs2IsQ6ykRqSFhk8c0L2Ex9zqVF+59NevYv/ufHZvI14tM9h
Xi3uIS+qde7s8fY+niaHR4M1tmDlJ2VRRHnzFJGS6Oe7Ts9U/u4GgvIjIP7w/UNH
`protect END_PROTECTED
