`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Miu1T2gvt/KxUjVXUpAneVCWVvxJmQ92oED6bXD2yisuOBehXTqrkcFHv7pnZIq
XFUzDPSAmEEUfg8Kwqg62hIsQkGspCTeUL8HVTPI9muPT7UrYmvvpVqHv30tvU0d
igW3T7t9ftcz1u2Rl+pz/6UU+dYIAfgTeFhkmVIpBAxaeVitL+MJ+I1kqXlJYhe1
j2BQZ/qXmimaxncpyOwpDILdiG4J9KOB3FJut3Lhsmu0yOuuNcDCyUgR9qLiTvMV
QCbTSr3TjwNBmxEzMDbisjmJeu6b6on6qBAtHk6K9qdIkK6CreVDxW5iGY4CLSjy
k6McqhnmRhnm18cvb10VC1944VaO3m9s1ukDb/kGqJVFLkoUVPvwjV5pz4DIN3c+
RE5ihJwMDfSjwDdA9Swj/JYYaRAIo0rjCZli4NEvYCSOKPISOgZ/AIqjhcmifXtA
v650SxyIwTjZz6UYXirrcePlM0GbPYEkMneoOKm74TD9Fk6Vhnv3o1F4I/aTN+R9
BoGZJ5xT33qrJzBlusouOIGx1GHhoosau2KttPpHTLNHYJZ2KX51mT2K2YhyP3zm
cMYQkITW37Ud5vlc8/GqRbyHE17XaWh5axTilsw5v6niPx/AkLxEAwQETRTXpB34
dKCMKKVxUBVTtJxAptwwkA==
`protect END_PROTECTED
