`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bN+8wX8wH7Yzh9T63Vmiwq9ErthPfUWooYy1Tl/j1+Fhz9Jnv/ba/lltlRq2NTN4
PXWl1vT+J1lYPIFfYeiy8n+FA8fpCZlo81A3Q5D7cxbz573Hbs3Pob5M69C9XKX1
VxA+hSzup/GmKeSzDGE9Ndv6GuKdIjCKDlF2FCGAVRRsGuZC27cx1cm/M/j3wXEO
+ZGtKKv86KV/Obm6iHsgEIdaox/QFLhvp4immjMtaUUYP1eIMr8IRRqNnLtp7tmp
VpUh03HKz6oEajjfAQ0jOKWUmIwkBO8oXvLq6o5aWicu3rvgLokmklRMXwYVxCTJ
anvuIOIJGlD4sce7oIZvgDbi7jPEfc4J734+cacJ1rI4Uu+9TIvW+XG5Atq1cYio
oFOdAsaKCwm73kLcV/vG8gYLWrqr/P+/p0fmW2ACyEezfbdjq13fDXBhG9UK+iTZ
vHwdnKZTTBzoklvv+f7Ntb5eaacIU05aht0fnZhsvTPuSM8nn7mNkPtvaBJpdy4q
xw3HbWLvvfMSxoX7wVePRxFL+1xAacO+YSuPuoqQXnNOB6SQY5StcQZou5Yme/Gu
g1BnkktZDHmIGW9uLFbfKwXpYv74dZaEQ5FuoF+UFAbCqtGHIigFYJHMCV+URYKU
Xwd2R1rGVbO7wV585HDEUTFAgtFUy4EGaWXOfGd/dAoF1lDoylVS7UMXhDeZyxEu
E/x10k4fVGU8+GKbJTS+Uh/yFv6n4C6/eJigP9UsxqLX6pvjxCdPiAPN+Bw85Zts
Jw4WeVLjfQGdN+MKp15gejqSe5E0STDrcXas+cP4PVTmR3HSeJDf3NdK0ndz7GIY
Bz1l3pDqkQcUBIsee8TuqAExoQMwOsrL+R1tLngkmkSPnDwf0iEKdZA7+CCOiOJ9
qz30jJdMzyzA0Fy5OwH+QvPZrUU8dLxAdRBIRj+kwSI02/BD9HhSXlK2hhgh2NDJ
`protect END_PROTECTED
