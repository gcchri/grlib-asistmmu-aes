`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBzQ0uzdusb67oH7h+UCEAEPNlJPnCKbhzbggOP6y5GtfAI0sUBmUYTOqgzApKPo
vpxBUkZTUtrRtAZ+8OY/7hvbQYOZBi24BYedZxgymBo2f96cRpfQX0RC45ZrcwUg
rdZfyMEtOf+O0w4U3HWOuHAvmoAbqrB5caeURdDBOtVFZ06kspcDw78iNxGirtHK
ZbpqPb0jd/z+lVYhdJt022dCM9UJs6Ry9QvpiHqhI8ai1ctFWkzPfkWEiW1SSxqh
aXrHmFVcpNqaP+Dggi4E9akfWBdNmTsBZKPAyY5oeyY/fGjbiq3bTIPnvnAuOois
LJoSBKySmh2U8D6eJM2TL+KZ9aMnc4vhVb3oLBczZUemM885jDJmI18JNr4Im+0i
wAGPTvNZS212p+A6DyhNlYVnciMrpzcIfCnMYCDsfdSJL2uw23NUhH3F3OVj/tx7
`protect END_PROTECTED
