`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OQ9kfdxDnzRa9j7+Crq64cjKIBdl9K8HXFsK+E/A0wX/XNFJBjMTmqjLpUP0pFl
mcnAEfAErPJ+wgXy8Gdqk2JkALTy1G5JY8y3ro0gOJkE3N8uvueBABoyqJuPCqhW
uFoEFqxTZWcG4yU/2yMcQkTN9SfPj8kCocD9spxOXj3cOx/KRpl07/kAJ0CL7Gvb
IPvc6omoEacCrtLAqlT91ESOzTH88icVJ5IqsaLqps8DZuLQFJsgCzffXQgW6cwm
bqt4EjVuMpNfFawDO879QkNO27NLw3W5BzsMd9iP2IzrCmgERhUY8Pk5RaCr6zhz
P6XTeXRWteajy6251ByGECy/QmlMLZxsJaye6p9kx4wqCd5txjyfixKEHZdb5aUn
N2knGgAtzVwss9T7sl/DmYEOhcmMy7/WPy84+Hcun6LyCZd2NQUfdFmJJEEXRicm
K+jAC/EU5a+lzwqMkWSglmXV1EkO6HYWNoQFuNo8jpSoM5is0jeHdu6po3vB39tX
klG4sIGlhcf19HcoLUlZewnvRIcQIXr9vKfoRd+AxQVqzgwB/k9gdFugsgryg8Yf
`protect END_PROTECTED
