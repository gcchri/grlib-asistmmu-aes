`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xbRxtiwSAaEeuPAi/Xweajh98C1Tb4pmcIw1aDtlNTlnk5Y+5CQYZC31vG8KzDI
WM5NOM5xh0Sgfp26NesKDzGQITWHfwOLoMzx4Nm2F06Q9Rps2P5XckHI42gIdtc7
EF1YlnhzfXyDDsoTdETYuwiIg8ErFymV3yfdZeaAc1oUMlUuiQ5amYgv2/I+9zfK
VPZeo/TeXhC3ZH+dROgpIU1Zx0fndKbWjXqG9WWoGccTFPyRkVDZN2ul480vrehS
fWMhnw2qrcBxBPB6eWtpJizpazt+sZ7EjnwnBtKmTW0J50rErRRk7SAeZmaYfEr9
3CWI5+UGOoY1LJLt2E5lQux5qAnteHC0axPwR17xOYUEqhNatAYRjNr13mgWoh9B
w2v7jV9l0uWjXewha2PZJpw9sz6PV156vHz9yssBOMW9k7pVmqdUVVAnnw2ETRTZ
2eEvrrYHb7MEhSnoIK2KtJoNe7DxICVTeoZrIoy8GEpqROAKzeSjqcvvuTtWNr8w
pMW7zkzjduBVADkk9rFjo8+FYmr2cengJjVJb4AFkFXdjsifJ58gCyNBZbE3VT9k
IQxgutyMt5aFZ2dhQ3sEKeNQcQNdxhHmN+WhkInhlR+vIO1aIbyOKl5TT6q5GEcN
Wdb8DiEG9ipl6UtgtELGmUqzy5v307lJFYj1wTNAFm+i8MyKF/AyTRitvmcKPgag
LxngV++BEMpx/iruBFbIsQir/ZgygUMyE4Sx8NjM76JyRfWoMv9xTXR6xXN6cq05
IWF8gXbv8CvhNWTHKqurziK1m5vYSHitTHMAjC8wYYal2G48RVknqapyHK2R4oXK
MqL6s/8U7fNQKUT+R3OBBAjKWAYyHBEM+3DUr2oj+8+zfK9KvUiiTgpa5hQGKAcr
ob2HtvR3eCH87M70YOOrRkahtHAX0YYmSyo2z58TsZpK4qOUgDgG4AnAsn5JwsuN
k++7izMa3akxX3znKHYJbxDsrrpcy1RKZ7ApKIoIB33wKY0zjowhQAmYpuwRPCpQ
4Y2jpUN9T49Yb77P2FDE9CY2fIM1UbwXgOjOPSA2ujtqQXOi3IIADqq7HPCfVIzr
FkZexVYouNv9qgC8EXvwk/QZS9dzAirWnBCv8aRI6ndnS1N+kp9ptrdztl4KmH1Q
zJrYebrmkZpI8Y87nRmejD5++7lAYB+AU9ENA2M/hQefimSUGS1YcpXBA+nC9mNE
HcMWaIC5N7QoTqYS0kaHO5RgjzetYhZwCXuCaX9w3HXB2oZ0tDiNBIZM+lHNJpGO
M41IfDRSApgCqQGKkaWN4G1GfL5Wvq2K3K4asbLe0Jw9D81NCwY1GEUpmnA7rNth
B0nDpYf0MzvFqlQo8OGmXLHlOTgak61cMDc97LP9BMxfjG1Ye1I2X2zBa6s6aaj0
Z+b1fTSjp097c6twuirYrVBijbSebaruCXQIKr+uEaUpZLkpziOz3FYJyyDHPNfr
VXxbjFSkvo/xJ2Jj0krIy90Mg4wIPCT8NyZxequjtWzZnIIBRexnoF3lshTFWaTT
BZlQEVOGcL9tjHtiO9/xzxutYmVKHrH8mQuHSJyP3teOHjPMvcFlPloHlGlq9sxF
Mler2SXnX3VwTeQ/CJXqN0aQm+fG2rqpJjy9fkmz0UQ4KXQXE1BSm1LZo5ZTvLAh
3brQekAY/hMx4UjRZLw3ZQHSDtf59iBVwKQmwqN9zllx1lvobWLLEMwiwXmgxnuF
uHeTOn5qsWpIEDOBUNADsqRN3lwvWxsMrssvgXojt2xrJYJ/DUmkLn1RTScNN5fF
pzFytlLMlVnhSrnuZZcZnOhikAy1+AgxQPqmR0NwBLcv/Tr4QqAlQ4h/fiEbR1TR
r45XTqhaW1xmwVGop/ODl76wsNhpRNMiqWdQdJKS5Je5EBDRM5L2107oSfk6xtZ/
fR7ThCFiQ+q7z9z8gn6a4cvaJfI9mWZMSLRJHCePsJUJaCo42/aioVPDhjGAxF5z
216q1UmUlOQ2DjWigWmYy7ZMvGGlS5LxrSMkHjwahRP/T7g431z4oV691yFUDfuk
Ttxu4DYkyKchRo0IhRRZC+pyRB1lGRVCgcAa3SO96aGYCDSHafpg7hCDSKFVnb3Z
CDAjqdlChFTpG9idGv4Pu8vEynZ5imjgDDC+cRJWxBKqbYFkvrEqGqxc4r1F/yMz
Iws5X28RQ8ukTFNe7gsQkxy7OwWo1Dr1KpTvYYo4v1NyXpcJaJyh2DLAOBir/uL9
MEYaQa5M0bHUu8L1xHkVy522Kpo8a8Ah2fF4UMAUNjAZTXZi4J+4hWy2tN5HwKNC
asLOkeneAG2pM/9/+c0da5VHZzxdzbfLZp0lBnepd0bxXEsXlln0rZJbei8EpUKM
3nUFOLxdRn76lhW/4oa2PCnlROxl+uRV781YdXfbQk3s23xL0E8M+JZRbWxJWJKi
yzuQXiV62UWDi0o3T+ESdow3fUuADYdcTpCHZEklsLCpof+VYMbGmVs814WsuIN3
REe6jYwORVEk8JmCaKSaznkNdQGmbDHmAf5+jHcahb2gJKDaKyInzQ0j9enTSBp1
0OkWKHfcZhhtGUkBm6usG8AKgjbSFwTVhC+rRBNK8k21fWRlYUoUvKMYRi4d8ktM
xmRwCha7fl2QG5/3sskjly8Og/yH8OE5bAam1iAkZM/HSL9wrNf5MlShoguQ39Z4
JMvA8jWksjJhuIx7TPEu4PDE7urhvpdVLsAR/Hce559DDqSV7AgsyYCkO6GICVjI
5Omhv3XRrgEiEzUSI6JvhBBFK+ejGe+Nb7jRNFg3uNTJVWqd+GMX2qaBfgRWgbcQ
49AT2NoDsqIHSTC0LMMAg1Z9lXwWjcE+jcHS9HIFBnL3m8IcTvw+jR/J2+XKLL0U
d/S0USAYgMB3Y/R10+g+KWP5xVJ0qJfFf+9lasoDdvKyaVOMBKcQlzwDBZO3l2pU
RPhhPSsmDMWXeOTMk98yRTmuxExUR2p/g6HoXFDuaA+jaOJBbRIbdXcYq2YSlrko
nVRodknoJ089R1oPI5vu4eVfocd2IqVUwnbeYywlePWoRFP1T9L1wv/tq1sKVuiE
S7MVsrvNElekS7sG/4Ha66oXmNoQMOHAdj7RAk8uif+xA9/hvbewdlVs+XqrSGfz
3Mw7ZVd7YYikLWpBnHfFxty3wOOhVi8Y25jGm1Q8oAjHyx2Wxt6d2sWShsRaw+6O
0VS2+w1xlAi2vrUgX8ReaaQxw0ZcbUQqdiG4TTe/x+J+nOkjWnKdvKJ9CVqQbVau
DABONjAmR8hXgYzcMMV04z0AyOwjJpmHLaQ7l1iBzbXg/abr+w48pGtkj6pFN0Mv
ybErRvyuqhB+Jl9hBIxvdx9DbVjCrL0RCX1bHj4xZdMe4dQvKUqO7SNYY/BHDYyP
Oji8cir08HPJt/xeRsiA0gIOKob0acKJiNkDNSXB15/FUD8flbGMii0AuU6dbEYG
Rd83EqfBulNBY3kGMJ3+flVLrAEPTwxyLJqEP1+j6a7Fdu9PlkC+UD39sXl9Om5m
W3XCOEPeSzNjDi7He65xEb46wwqr9dWVk/cl4HIc13zsQ/IAxS9EZo1oa/yCvSsh
9c/Luj8jzOitX9bEpiPU0mGGNe1EFEwP+k3flK5gm/xIrHMXS5jgMi8iaKPGaR3A
ns1Ms3meo16PfANVyrwrNIx1P4nOVP/LWOTEut9vTkM1pDutJk0sESlnyh6or1zf
xvdp5GiVSDL6hrC2oET5JIURPHwHEIICU9fgWCaHE9BCKLuMu53Zi9Piw6C2xUXl
aXmLyDPTOqb1dGmqxoH/1K1pfFMuVT1792OZwrVaWRNekQjoBZyT94OpvtF//67j
7AOd1T3ejEPzelqvVq/gbw==
`protect END_PROTECTED
