`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIjrtqA0h3YRNS3VizTu2xQjQYk5V1mt+5cqv7dE4yBVjkKgcMJPXEPfUCZYASr/
VPnmBr19hqQIxkUHycN2kcTy1HUjYZM5cj95Dz0MvoaHCl9+B1UPI1hysIejCyN+
GrZBcNpQF7Rz3oSwhQD+LzR2SU+UogoiL7Wjrk2SxAhx2xWzvS3h3Z1nkszaFjXr
RC1+O2ARiguLu0BFVgXTR3ZWIgTljVbxZJZ714+nacwjQes+iKpmbzBmLRnCPI0Y
nKQHZ597iN2cC40Z7MbmdETcwF1QVuKrtxFnXBerkreUnVEj4//KgK8TLzV5uiHf
CxhUycSTxRsswC+VNOEGR0JHCVahG4k8wDvoC+DvFghir2HEij66D3tqjiIhReRi
QO9OSdYPn13HdFL7flLEbB0bZVpnIT0z9ItULfUnL3s=
`protect END_PROTECTED
