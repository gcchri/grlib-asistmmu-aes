`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BrXsh7X0ZpZrm+gY409rwcdGbBi8iUJ0Ty+pmvTQmFTbcR1V3XnFU4SEagm1nLLl
PLI2GbXl8XmssqreCcUxZL8XhUMWi/ge4OyHu+Nd0PKVPX2WoNPioE4jSJtnbmP0
XnBT3o/Qq/kAVsO6KhFN0UwA+HJBenHKuN7Ort7IqJR0nrwTPkdtZHS1KLpaOBE6
WJcc6CD8cJ418QPiQAGqqvVVBkl1ok+EIiRbFzk5y6EjQn1PApSgQNJVr8zhKDrD
OWZQKYKK5TRQLORZYhAsSuSbJ/R6YINj8Z0YEiIfH43pELPTXSNHjly8fDF7+C6Q
72Sc+4FQVF54AhoHlGlU/X92EZCUfQFQ3xZQHGjckb9kTyXLaY3jiutDcwrYMXX7
C6YaZEVvFKKiWDkD4K/LLAVEclFU+03/JIhNVD2fSwblYa9MVl9z4/N6+Pgl0kuu
AVnhiUwyM5hgKa753lwJ4SCpHHKe81cP7CQxrsulsjXjdjPOl+9drHelKfl4ihtx
lFO8qmqXa6/dm64jVFn7hoFUWn+RVNVNVEa2D8PoabyuKYe79FD+qEV1izWHwf7U
OQ1T7rvZguGOIUsUCenlu9ng+gxig2Rt7/bF5gjIfdlbhLADp5k0vSYbPUKBRyML
DK0+i2aOmWjP8O5G6KF+C0bvUvfa8ETfr/x0ygWnMJa/Ps4SxXAm1NWY+a+OsbE8
504/wrHTzIOQb/vbOE1yLVjtvx6U9j/F7sFutQ3pimkDL9hFzlTSwM6IMwsp2gfG
hG2RIll+g2v2u/AmLTlidBfOdwPiCPuGoLLY1ZlMK/g=
`protect END_PROTECTED
