`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RnTnU+hhXo6SlzCnRIJItiUpsxlQH5/xgO3YXz41UMkftWY5qIiy/da8goANQNu0
Gj2Ptxh/Fw58xnZ0U4vJD/6s3ZsuK5NZmdW9jXSZcSAJnh0k36/N6Ulrng4e3YNN
Wk52e2Lwk64pvAsG+ypDgAmQRn8j/UO9Hte1UR7pcj+GikhhmuVrmRlUNJHm2sCn
ozCJTzQhXtBenoDOlTkgpd91WlUK1W+RwjpFiooUICpVqqHro9YrPDj7vtASCA2X
Vp8rMpWFXzSkXTGiU9MvrLDXjmAB4FjewjobTjt9/dWKGNzepXjCp+uJw7K7ra/3
e813SrMvKsLbVt3iDo1Mzn66RqpxGKdsQwQtzSRUG9ey9XfCuqogcF+RnMCPuujp
iXyQIdoqUy7ISZw+cERjb3XO+hGL2DMDAEmltBATOyTsmOXCrqnBcK5zGLph7EXU
QMUqautbrPpRaKqDWAYWmZQc5JSO+WlSn0HVauHooBkkWtp+b+sAYBhyOK7940/B
l2c7SsbweSQcpV6zpeUqRAiScBVYBtuU+I09FxmWkN80387vgVPvPWK359TelDjp
gtiXTV3E2feVqgLit+dr/5afCcjPXU1ZCKVDsDvQNXDhWNVOfugfTEZnNzvurql9
5kGy2iuoosVDQ3yPZDRfm8LCKrZR8e4p9Hqh66b4uBnQYLMBXVR6fENX/xZKCJ/Q
GPLtIW3EvAas6YYxMN2LwF0oH8c502MIcgKAENO2X9xXWHOeW4EmOb3GEILEUgeF
I0cfZl0RcU/Gt4wQL8NO4yIVxbua6mqtWh2idHgIPHeqmuLaxtqf/Cw4YNjYDLsN
XmfUlvFp0Cbo/u/95wtLPwUM7ovZQdo03WALtL/pL3Tjq3nCJpVqiypd+AJArjlS
VijKlZYqJMfA/sXFZECZNPnbVZtDGQzXmcXD4rKYN9zxA+SGiQwSMrxE8nqCh6CP
E/46OBm+dMAmQp3dm5i8dwOfgnGkbj7tX1e0tyOFYuaIDkRqU2urK8Dthz4nWUwd
QnYO0z51k2K0hG3mTtdoaKwkafEpB4TUKhQGP7uc6PU+kpEgaSJa6UZy9IOYEmv1
OZPZTAJvjFS8WMwbzWTAyYQS2A+Y9L/kNXmuv+S1a/PiJDj3Bs6J0W2lGaRZAfKH
qcxNgJc0PILK0qFencW7DPoSu69wVGblWSbLmwRX4mOOhR8Kdfv9RANUc7RjnGJI
TXby5M+Dn6DOiRxJVSylwwsWWqCPR647guPNBho33XJodyyygc/aZC646Zj92YHY
lOjqpB56qM8rxKKPTgGJlo8yZAN5fw4BkDo99VtQpqEJ1N1sEBdv1+r8Yn10UzbD
oO4Oi+24C2XoahlAXCzi1telkztw1d2IiazdiclDM+8/hI4ZEhWoWRTW45oCYNmv
ti15rhnyxg5u4QDXKxkilZffE6ra4e3nuA0oReBuV6+b5FJ21/u4ikcYHNj4Wxwh
5fFNtFrBnGNOLlvjvCB77zQxIJYyPvJEH1jUIO+3fSLPaROspdjNHre56jO4Cj/b
n0n/8MR7yk5kw0e6i4kjHcNZcbjht+wbbMe3LknAgax22cjFG/rqFg65yHb4Tfed
TF8E98NwYjIknZIxK7P/mPBLHkLHd27hJaFzuKVMpa3Ga2A2Q48f/5zjzPxjEz1+
J7GiuQX4pxUd9+dQ7z1CCtCNEtLh4IhMrGtymHOnURtRbFEb2dy+yRnCNQG3ukmB
cnfokdHjpSAS1ivt1o6xI/PuHO9oVPTqYWu21TYojdMCR/6ddp8tbOY3sQFJEz7d
tAk/8N8BaJOCI0xYLXmP8MNCXJ0zOs4y++hHw8M2I4CJDMDfZUnaDB9mCeFH8y9+
CnfhHG0WKG4Syiun5+IXboA1bHUxCzTUmsYP83bSdAtFDNK41fE0N3ul0YEl8/H+
pfqOG8Imx3hOJqOpYMHn5XAlB8+984bArxwESAGAamFY/uOlAV3PiqBo/9GpeRrC
RkDYaJqjdv7Lb/XTb9bGJfY9bMTiwSO51UU4nFNAq4FIXeZI8GjeXyOWLAKt5R+w
YMnzZyyNFjSo37coeXN1mVRGf4eWV/qz6esgqymul6ls+/CveBUgTC/jjJJRBoa4
BYxnd1c9yhQTYvXMpmn8HcMr5CDFzmrFtb4nm6i8gCg4oELIg5NrD9BgGV/jBLwN
pTq0bYw3ClWVsD6d0ZsI76MhMf2NRbEn4t8pH6F7PIogrUiDTBRdSj/Kr/FPZP9R
3wqBWk0UkOek8mD1I/H99iVboNqEXZdM4f2bWedZKcoT40GtS7IeKf+HAhUMKTch
VNAh3uYl7PIw7JGuIYZ2U4YAwmwiVb5VjJxdP7EA3QXbMh78CayKlIjnH8Tw+oGv
OLkozALkZrOXctQUgAqhtkEGE09mEGPIIWTvyw1I2LKr9mppTuXbPC8dl+6jQrWJ
GTfk97Gx28SAgGdQDRP2T9GaavuTVx6Ntwx8mD5SSqaX4ezcS9CVMmA0+Ym+YJ1O
V9pWWmv50jDnXCFPAwU+yJfTq+opP1RzCAd0YWqBQ6WBOYk2nECJw5RxzKSFPc0V
Rn6uD/MzO+PCSH6gacYhc7DGUw1xcXMmPJJOPOExlVEJi0eJWBvi6yIZEnYx4QCk
/PXMSleqPYa/YsXDccoDKuRZYUidn06r4w6j+kHLHD8eiTW+GMACzq95bGtL71dU
jCvfgZt0pUn79D+qSyz/pbQbIsro+v4oliabOpdJ7MzUJsWJlRPgVpPYMBnIcJaY
pWfqobADlb6h1hlUwBW0oviBsuroBfVphyACtsuI/BsjnhgxYe5WMQJsdc+p1zUv
zi/nBpHEZZWw/gDiXkEYqeFVvE/aPzsLNfXz5iSK1tSmQ+QH7wvu8kwkkpPmiqGO
Ha1h7DB16Y6bUMXZYBeJmXmzWHN9le+v1DBdGSmIPsD967X/bFiXR9g+1s2W2gHU
XGGU3h2eNdhx6yVjNO5/qCqUjamEIDNBO5p0+sKyiITvFGhbFJpfN7HPM0BJg9N9
2poLmXaBa15PPivbpHbogLkO4/IemCmcNoaKsrKd06XVaecF4x/jiZ/PkMhtJJYy
56DxN3vf6/Mg4/kXtCery9gphI249Be3GvaJFsrwEoo6NkiWkjd5UYsVehkUv15c
R1976yi4ntNMOpDHDGS9YEitvuyngCTX+vgUKEnrzbNyFSEt2i1/D7wLRGxFEPeT
2hWYQ7U0v2Vk4KLacboBJNt1aOE/MTSeJZ9oprMJLg1bB2+IFEJUgIYnhot/Zqvh
zjWDO2T2jrHXdcyy4I2gkVXtu7cx5PhydJL6vdF9Mt6Benuo2bjRnQjW7Q1zD4T9
1/JJU+x1oCbf3hTAA2ESU22JtyHy7XuWfqqF8gzMXA7dkhSrW07V2AyQkShJNbON
0qyhgZaWFvf2x2vdIEj+GjmO/RgmDTYWG1aTLT6GLiYLPanp+9sgXkndd5bOHo4v
ac/U8e1BQgaFKF3n5ICZax3yyqSpC5hT+54GFoi05+ir4BFYde469hsecqsti5Ml
Sc32Gd66X9z0dw6hVbfHOJDmDeKDB5oBW+0hesW6h/aYjvyIW3Ph3Cy83K6VK+95
HzNbtzwcfcsJU/06cjliQLgRCNArBC78nN1ioDgaBu3Uc0GRQeaa/zKeuHMiwvpj
n0h1+jzeJw6LiA+eji1dGDRDb2mE5oyRUb7Pd9zHeyCRPV9nygq36Q97dwjVBVLO
JadPrQh2WJdbTUIBngJZWhNz2pk9zs8uCg1iAdjAXKytJzwvPzmlIVaUqrC3dN/Z
ZgDdQIJ5fWdbvJLeFJ6JXt6FKTrpV3TIxFHGDbI+AwmnYg2BKta+6hHGcdySgc1D
LE6m23uvV2Wap1WHlw0FM+Y6a/yOYYEMY+ngWH5lqt5yoPwo4pLYWdWcZ/yRjsOr
ur8P7pzxUvja3YitrQttDYX6Vu9Tn6E1QH/ZU4xbmiaaLGdOWzp08c0bgWt62bgc
rW7y8lq1JTdC4+30jRjnZaivFUEqGVT1K1ZE4i73ec0NTo+cR+vDUKed/mwiSUqc
SpBWbdWF4oIdX1iITSwDZ0F8UtBm6ruT+JKlAYOlVmfdt4qfVXs0aILdS6hEvk0Y
uosgxbqSV+8SPC3wMDHlal/VR+8JK7QLomzByAlc4YIxRVHI64fbBwZ97YBJ2mEr
VULi4kdqVMiUMsdQoxquEOVrJtJRngvqpWSmqRu8vYe9OdGuWXYEIHBTHWC9ccjF
c2++zWKSkEUc7bGnKVkKhV35QDh5gek6Ycr4KZ7xFAcbQA2zvM6BoRp/SNv/sKe/
kyHqx+oe2oMb6d6p/Th0S226exHkkXt6gtmdc5yxBMOQWqXU0j+IhVMRyZ3eBHG7
38qU+yeh2QgUipAbTjARfRUBkgTpbYWdpIX0Nn2PoE95sVOZp8V3JAL0Y1zWZVNe
FiXNsJzzooVNLWB8USKdqO+bEawF6n/1aXieGfWjmGLhN7x5FU4M5y6b95WIdWoW
WCL0ls6o1ql9y17PPgEiSd7pzK1OfIKeJzH9GnKeOYSf5xcKGA1Uk4ja2/qAa54B
nKEvEwoCo22KS+4/qeq1FtUbPR1AWTQpCS4/FQw7W/qZuhmXwfJB6bb6wneTnOC8
FoGXsMTTxCRrydTmXPFbj+EX8+uzUkUNqIPVg1By77cX3VQraGiDH5H46Vbmq21+
EED9VjHbw7fv4gvfBeEpM9zgG+9HvmCRcb8S4KQQJradW3qV3UaMjRkYT0X4XNoK
r1p/Gf6h3/gmaQs3oySUTpXFW4AG3kVoEN8dMHHnJkkupY1Oo3zTLWipm+UknVLk
RvjJEkrge8sJZ2Kfz2BbOU/L4LdQk6jP/MqZfHZnY8e/f73FBhEYrvMMMl6BtvOq
ygh7c4SiQBXzqja6dd86sJRkP7jaKDYUVRkJO29c3acU/CypwLkJ+PhPIHQRkIW/
Ca1jH9Gqulq44rywQNLj58i6z9V3tHnLY6jbFPFm88Ycry+JHl2TBOFmdD9UkRbg
Y4k75zZoNAQrABeNFwcMz9SHOiTtifqjFAq6SUESE5j/kJYOmnOVx6+czhZRinbB
OHGEosmixapVmrHZLdZ52jxYTCDjdl06mSRRL9pqBSjBHq/X6+pSOVRHqWj5fTn2
GvMMR1sDsddxTZM/0064AyyOaTofLaDlhEdalZjI62omPdHsnL7k9o81EfWglfHl
bJ0ecn3Lhh05HvXc2xcw30RGjwURJ6CiJ6q9HrOHBHQaspsj9Yz5hV0qqaO9w2RO
xOxYukY0Uy3DMO6Y+OsDxZBJ+kH4jjZQbjRZLk8/cQEf3wjFP5eRpV5D+O8S6yA3
/l0rV84TmVdPQvyX9OtCgIH9G2nekKD1O0rm6RCMqim9lZirCBsSlbawDh7HhhOA
0MR4F8tPPATbw4uYZsGBoa4EfbVI73ecSnUjFnYw1kUd+2vzcB3xtz5iiq8U8gLu
0sx7T2xV+XDUpjgk86xNTLLelwJKMV+hztZmCqSa5jNWZa66X9FA73LxwBskNF07
0MdlDmq0S5uDn/5VEbOgqBaFDVSHBPUFhsRzF6Dk14Pkj1fSRfSxn/KmtjNNwjBE
ili6Q9yUQdJ9ih+xAtHKopq+c/sHeuW6btP/DBdkOHo59hiLWlmTFtdB8PSL8Z67
L97DeygPb/6+heEjXOUXSXAXwyegjfJDvYVHIrI2mRv7ow5szFktLC4yMg/IZhk0
RcKbJak4E6MYqKcuB9yV+cJjzLtsImaiYBHEFwdM0pVU2X8B4GP5r/ZMBDwHx5Ms
EmMEfEqVhsIi6VztEVC/7JbkOw1a1ELhSaAy5gAA722spynaEQj8DwIGbAWD8jPV
7yRnAErxb7rEU9dpiOirtI68mEPPx7Jwwf0mmGhzjsLbLy2wmFdOPRXLCvQr5MQU
Wt0JTJjcFbHmB00fUNyRBAHV2oQzV3xKqrgkUrbgMlRIsSBvKYaEP3rfyO9W74/z
XKTdByTA29GmmqHHeTFsJIZ7UhFDdqQy6+F6pornBMXOPbMNP9/ube4q4K2T3xdf
haiQXicvL4FFWAHFXttVW3y+Fi4rHRC5aciuQZ4jj7nci82LoR1ksgBRC4c9kJfy
iYfxjtcbzQXXG1P5EnGr9s76cgmip+4bo8qjlj6KsT605lPDF1owansYDIS+8DBw
WwOT84ydv6bET2IXb9AmpgS6ky94r+24UB1yqa8zxFZiYalZ26PVbjqw47aEIjWg
Tk1vl2CbPOxZ1jL3jdRLr5J8varPFbW+dMcaHb+MEsEz2ddlJwfoP6j1my0GJO/f
0L545NhhIGsZYmyunxITmee6B54a2ZTZY8HWc45SywEnbncJ64GD/c+MqxGZcBdy
ls+sciSEQBfk5rNRkBgM+AQHvkSoI2VwdNXwCrW2fM7gsgfRAPSwm3z503xUJvRl
+BOi9Raf9Fyk3i27dJC04s5ORa9xTrsJc6Bs0S2P29iKtsYOtKX+lKk10D+AXHGT
3ABkF4+7eQCSPqJPbcvfTZL+hh1R/Nkk6JU00tLNqiCebW0xUPWdFhN1TqdCzDTb
p19ZcdjshWKyvoRiN62+3e+r7zYApsZeH5DE9jxUUuD4zWK/CAdqLAZre3v6gwyS
vL4ewiM0L7n9bhLz0R46tyB4tbjbrpvVFG4CgnF3uctE/ntx0CC63NpCLbk+t3Bs
r2RFS5i7yq+xq2W+6MRyOlM8G8Lvh1J+SvHUioNjIgujs00vwswRN7lyjK8QTeMX
EdBLhdf49CxdBTwELOb1Yr3EHiUh8Io70HX0yppeWFeG2X0HQoukb94O0VaUogMS
YEoL5TKctntFXblXG50Mv/GTbnNP47S8EX6Iys9qlZJTg8krtdWCy+V/uhANft4S
JgVp4qUU38aa4k84Z6m44wIp4+04ZQf0OVO3pd5PpJSZkZvXVa0Iy6Wc8obfra4D
JVgcNml5c68bjPUNXm2/KlG4B+5na4xJ/0x651eQEKR4e2NCCKc5GN6QNuT4RM9f
U/q1azAPRKMd/OaLbu8EFgDCGmBurG0p31GY0lIinjfQYRo8oY9El7O5ErJLnkcH
9G238kGdlQQ9um4fcAhEIrvKP9NwF2fCYLMjemtBySnJLOYB1omDfk+/p9+RkYEb
tzIxcagtV2FXcgdzG71YBrf3XztQ6iX/V2YTv449W91XZcA0a4PX0yjo+oQRIAU8
BOuHsc8zryeqgvAUVzNlxWqG17RJOFfApvJeL4nx+A7bNXpBC6l05qpqV65rp+87
k6uIrlp3xuLDbLOLR2ZCVKKIidZZDaA9Nf5F0wbF58V5IOPUjoG1JPajwmy0UbNF
gUeFnl24PgB5NcMbxq6kc05KvNDCKsVx0yMTMtQMD6ufndHql/Q8LK8QqlGTRuOE
J8qHD6utlxljRKoBK0nuG22lDL4gGxCzhpQP5wj8MVeZQdkxvUBKUh+LmpXP7Nb0
Rznp//0vV674v4Xld605Jl1fvNPVJ36yFiRt3y4ZMPOD7VSsAN1yV3NOQ4MgYQCF
ZEp29UBL8RRa+8egmiy0dtHhE0qoE0/e4ZtdEaBzbCsn+A/nhETwxN5xet0ePVVZ
G2WwkJMgC3E/gMoSDNLWbkAEMtUNsj5CtRwyuBLk02RwDCSBdTkvGkREcvjj0K3A
502qxdqPoLofJPxuVXKi+0yLpaU4fZxKV6hf3XUkNpvZoa53C8sQ7jy0zCumv3sJ
+VBX05fZjNe2EHTWXro5NTRF9H/dxMKf4MODrRVv8AWoNoLnWiSvTP4TtifL2zDa
pqAMYs5wyS/PRin2BkHObOuTG3f+hjtZPvuYelaSy5ybPcgAWfnUDPuyVpyXnAmQ
hauydiT2PeUd2VVKutIh4g0nGMme6piguTyfQ14rzC8Oor+zCAqCrYxht0Qe7NgV
t6d5ImhMj5nJCnVEMvdtc3iQhbbNxG54smFoS2+PrsRZlelj+JYgmFV090qnftaa
ZFyhY9x0XlLjj8ghPpUhnC4KLQeAzpp4LqEnRNfH2jfvoXOMweTRlF1FdMywzO15
E7zX+9yeetjM8r8bPIlXq6JYvaHLEw7G+oyHi9i5/8mgz3PubrzpoMRH5i/2+/v0
00Kxwm+6ik1D76mWjNsx32cyoE55BgQIo/v6FlgPjUoaMZYnINcdvEtODvBiRr3h
KBO1t4SQAelIq1eq6qAW4y03MUbcf7Xo2flCVl1uCJyBM1Vrq3VcVIIHcyB1wF/o
t60Kf2XcrUHEEeIMkxYu97VfXA/2Ny4LIyzzH85vm3THSHoDjP+Li0I2HEEUafDz
FpVfd8t2SSZ6EaRDefxm3aDNswXjmeWi7HGf+PidK4z6lorsma2uoNpn8StKoOpg
tkYp8XFGXU0jCTskRNK7/aw+ExhSuJTUf6zXO8GtdI5jnAzV6oKPbFgqf8mqE6Zb
3sUPB1LElsrZgUJfhYJs4CnB/YG7+F6A8ywL5aJprHArFRyJDotJuXL4uWrrJ61R
m1l2t3yDRJhB9Scl7X9ISH8mOMmBptqVZBYCNfoP+TpNHwh8azPiaOys9ezfXBXQ
oSdXvyX3mhIpFJoxASQNxM3FRgdeERJ3LgWur7AlATvE2zCnDWNLzPRtXGCkChrG
MRKBE+jmcYWxt9a3POE1bvUegm4ujlN7augRzAQcITMkeuOYQEF5CQXJ4AGr662y
v1Knu/iXFqX3YwD9n+b9ksvttwW+y2Gd2QFHzLVl92kLwLc/gy+OjTpvIPeFWVO/
9gGVsvDaetaAgAgIpGsxEveJEEJr8mxLGUMPVDWnRxAwLe3I4vbczTCJlcsSjXGH
wF4myy8PRX2iQ2BO5CGktop9oYDTun88DfBbcbrCBAaaVngGYcEPJoeVrT+hjhN0
5Qj/Dzvmqn+WPUT5Q5UsVdK9eGt8ZScEf1oUJRH6rpi074aLehs3nzuDaCOB6GQM
lgpbiEYWr59aZVJK9dTrdmrkQi3YzvaZiOeeizF18eO1MYavmiz3Pez2Xgs3TAKT
RBu0IAMz27bURfm738Pps2Idl544hul7Z2X7gwkhMkq5Qb9yYDRILqj4tptAI6Ao
jNX+Xk2wR2bt+qmW60qzErVxC2QZHGtsB3jPtbBTb0zccToB+5AA8skuH4yy20DY
RDNPf+thhtVUpqTDEIJJCjQ2WjYJBdd2VXtu0Uy5dgWEe5JlTqRl/NcBxge+qDps
5TFRAfJVlUnaREasrqjrhKWvQLIL+3y32+ls8rwtZE62Y3TTkeSg7dkpAI0FN3WE
ay3/xNPVACZ+y/YH9TjkKxjsyEpqEnD9VUcsnV90ph923/UPuUhRWNhwKZXhkBZB
CFaNbhiQDS0QzV/gQQOxSwlSpCm5sNWI73AQKiL4UPu7bZac4sGyF3fqc0u3Amep
cMsj+nGrhgftk6h1mAjQvuTpJ3vo9UGwKS1kqDMH3Tmf/GKIkoNvAUVKxAbQtFAy
/VWy3nTNZV20jZxdtGMu4FF8qc8Oc8Eua4IFW23aD5vyF2FQPbVQytaJbtBaObd7
yPySYyq+L3qRu5CpKkRSu0mHygAwCcImYOKMApDm8xwM+RIOdOuO6srXOrHhmq3J
tGKLXidDCD0VXN61Z8wvCSPVrgcmMp7adwvN248EPhBXJtzk0xTZttHtEJQTk+4J
5+kU/pjstVAdLgZehuJUB8ILFuU84PUaTwXl3WwomtLmTZCuXBGo8xKRqpmVjhzx
9TDzNA08UOztuQ/yowWmIa6KRTTfuyeiE/qFn9XNh6WjgSFUPDghEHgBgNNecunw
ECNAFzRKYHkKck1gpPAChiwXIJiOyYH7ogvzTLWR4GhFyG2w3RNmTUFJ/peYRmS0
6yR7yhW9vL0Jj16lwYIyuHWY24lAqiKiQgpWvSUYLhSCyCRhbJmdnJMo9hElJED4
97WHk/soF29Ae18TtNFS77m7v0oCZiMDJmeOF9fWEpmSbZFBhRSDkJgfAmRxUBnx
WhNGy6hY49hdeWiDgNiKrYxejguKj3Ga0r2JsPYdgCSysdv3pf9dvcfazSxbZuFs
uc/f/HEhr3gyCiawPmupqk0lphed21R/QQgUS61GvoCSMYIw+gjXcZsZF3DfVCCq
PPYU0c0AijShcNTysy1gjsNeIXN+BhUb+7r4dDwrxRI7wzoQ6agL3+fWqvbglY/7
rAaDzQrQBlHBgOv2xxmmz3MTGMyHr2FgZT+Pf25rgAU/euLDTBa3MnbwWLvrRd8g
90Wo0QZmuUWjOQs5wGeLvyaU+cCeIc4JkUhDt4UcuR6uo3IiImjjctxVuXJg+RmY
Uv/21YqOhgpN9zslAN5CiTL7FRqQqWLbalcqctYKfHpTvJzs3znlKJJxEeBzONkA
Gy2aRd3mFyyGq8AjnXjRYhjl8GOiH3Xej9whdA6hFLvctE/wvte4JweiYTAAGBjf
Y+bdpp5oc9q2ptO7DyBRd90JMfsDi96SMsQqJkrgxDC9cNuS81UMSqNP+oiiZZgV
S1lAo28j+PKEwQNvE/Mew5r34owk9ir/EDXMRjrO+ZDkWW7IQpMS61al7bMk8i0G
Jek0PP/dGZe4jeuG8M4DXyJq+ASHgtbJJn7t2txDl4fMVdPsxyppXcsykkTgD0L7
7eSxSBi74C8ybxRD8u4xzLvqWpBHR54SwVt3YWLp0MwevNumTJDah1z9KgYo+quM
UwBE2u31arsuXRIVPGBUID0ptS9W8XzieybFITy5xzcr7Dre9zspHXV5b9Ng36ib
uFYLSxQ2OP4ePK5q5MdPWM6s/wcMqaWoPI/2h9KLwh+V3/GUWmFUdpRrztuFo+oi
zIe+Af3p/m48ycZB5R/QsOOpJZQ3l9YNPYOAdWOIxoDxRLsNCuhRH8b/vxwTyyBn
A7zDlv7bOvjZ09WUQUbXuesNJdrJTINX8Ysh7YxsNNmfyVlYbHw9pazVvr0cdysO
hUv7mAI4GAdkuVY2HVgKkNMcw3/5XCKV0JY3DQ26ZunqXUYeEQ/NSMxwXQ0LneEN
j4Zp2/EwFs3ftHHrEGIvVqqsuZKEbfr/NRXVt80rtrhOy6//v9jDGpObu5dTr62o
d5ytp2Ki02frGOODnGcOLVfD+Ixo4PFbs1XwJGVURgVOCThh03DwXsUOIGTQb96q
pq1NIdzMSTRrceJKaGVG24PXQIGdGHr+ij0B6OeLhpNCvoaFW/WdNfF6gIw1zgsI
CwzHm9jdRLg4wIi171KedhS1kWJtEivwc3ixY0zu0HOdY3kcf8gKcMrHt6H5QFSR
kCaQIacCQuESg+nMghK3k37zowNyC6oiN8Uwe3UR7nX2oLyt68M64pBOMHYugEXT
cyVJ5JoNZwc6BCxf/e9Kyp2+MGQrz8Z/fhHJ12JZo9L4KkSyXJpEggJYKJfcex8n
LPigpw9Gf+wVSEg89lqtB3V7FgZXMHRe48BEoiCd3G3zk8jyzMVxPrOUHHU/qW1g
y5ImUlKYNCKHkbG13CAgzGZwsenRlhvpdIStYjCVry6sIKw+UmrT3VqxFTwf5s4e
PPKcoDNdZ3DTeYAtjlhq/YdlBLJOggC66zOj+ul6NUVXjo4Ql/OXEt0DzM4sBlSF
CCCJ81RLroY8OCDzPfHA4hUWq2BnyY8K7sGu2skGm03HukXrggWBDndN/KvEnaQa
EEZam8DxooOFa2V8oj104ZkqpONI/tV8e72EwVCf8lXTD6v8NBweElo/MF1AlqEo
IBylzvWVpW/o7T6qQqxmhg1urtNyqewYbDMpsu5iYfXjXsU9RuEsnCAlOBQ7K4j1
kSPr9S9SFuHQlvw9B7/SwRT5+RNKOXAaXHjx7YaVNNOuvDrtfPuBAd9QlPtHpF6M
N8DifXr8QieU6KWEx1bTJT9WWKlIdDav08q1wbHdPtHWyiElD8xkke/bFZ92bx04
TKs2vpYUA5pNI1NFFkWfsy5gXEPAQs2ttd8ZZKychNtRa7BFgW74edgha/Cohii/
1Vy+VvD0PdTEGslBeb6RjaZ7qtPs++AuzcPvkvesFFkX4rXB/4ezE9UhyPcGjV7C
zEZ0XXO9NJBACDw4fpu5SaAa2ukh6vbUNh9vSSJye4TVB/tkMLLgm0p7c/Imy1hr
ySrwgYotfUWcaBBUHwWbgfCfhoJgJf4Dw7W2gm985fHIT1fdiEIsddEnnQYrrry+
mWkiytAbRcpjeH4Tfa9ayyFkao3jcJGEEAl9kY+d2pHJAl02YVqnzait9kjkYDvw
YvBg43IcLJzehdH1Rbxr6GVSe8FyAiclUGpy1Qu7B10rz14l6LhwXG2z7Mgs0xum
OX8MdeTq8OT2Q+3wBx2gVfGzzjuGEhjs+UjQBLU4gX+LUz6+BnFzpVCfAmiRKa45
R8FE1qh0cNWzJZ+ac1JamH3AfEm7DAV6PYJXo/sIDTdmsp8yBOU/fkYXVlZpDqTz
re+9ce/6gSx0RbjHFwwDMl3VaYBDbIoZdWP8Wd/JtpaELAO9+xSDinIbNBNpNwau
Cf3KA/tEIDLDlYIV0JlqJIckiIwDQfAw2/gyUT2B4D/FxJxoCope3o21CI75q3k2
ARx4w4GRQ+gsxWrro6fTUOVbk4gu8plqtQmnvCGVaK9nX7ORqJTOZHyJ3uPypmCi
lVxQBI0F7mio86CbNEjq1kyegqyWfWe+odb5ygW7/UZLshhRLFK9ak1lMttcCtnQ
lXp3zoDOxvOT4cYS+PMFOp0CzEHJYWqUMG3xC/G3wNIjFv3NOCZ/tPSFDFssEl47
0AqtyeqW/UwZtWHrbWxOjckO8Jm5cBqHHsq5UgsA5lBmp5gItBqlChd6rgX/LbO1
0ZfxrD/4pZ4de5zn+aJ2msg/h5F10VfJWDEdlPxe09t/+76ueUHbtCUr+YY0vHRi
IIC9gJhcrAJe4WQGGXT1IY5rUsaDyFDqEyvFF8l7CSP/AQ6ZsDM0v/ZH2hVeQDDA
G+XIcm4EWdM+h/MgNYLPUaUVe2EuvzFOqcSghjBaEgCHxTU5K6kAdlZU9Ri2hC+J
KfiJGppaYvcfXmLgnyLEcbQu63/092zExvsymWEkrug=
`protect END_PROTECTED
