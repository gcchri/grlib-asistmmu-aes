`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRYkW0od6VcWiFTcMd9cGhyflXP47w7qC1SMQps7N6RX54m+akJEgesCnBlcVu0W
WEtYBfLGAtj3yJUotAY35Jj1Rv52RzAmBS4RvlcQ53RQa8/W5aEyHAN/d/6LxT+r
0BmEKapqLFeBLpmxmW/CLhpzfjW50hY8R+UU3AYraBpNYRUu8/1bZ7V477mMf7EZ
jpA8z+qD9fYrLhNEZC1cgcc9u+oUqs10oqUTpN2dYAPfFAGNOa8WB4vTcW0g3PSV
VstIoa6QjFEeA/yTY5F3Y/JHA1Q6a5JNGF6/TwR9OiXQzF7Bbn+j+/8w0O/oeZTB
Gr+Y6EzUplwRjOo/iydbLh3ufVYeDp0sjsDpWaJQSabonhOKfzbOdylRlEHJAzgq
jwGOtMLiv2QOZO20cfto2IbiD0lShxF86u5IkgvwiFl3+yKjdlyhhYtAAwno0nLI
NIY89SEUHojj+FkJcB0MoxRX6pUAVbvJ9QUKlq62Em5R65KG2+2AZVNCDz6PDsPB
94Xq6OShniaiNmWxDtPQZlxzOTxR7D0f7yC2ElUn+4EImjV8TWO26RLi/k6WLxi4
D2mNflq4kC6WG2ODWDn6bmunk/NNGS+gaSZ/zxxWrc6wHyoLlpdd+1FqZuY5blY6
bXV+Yb0l7nG2dM4Zx9Vvzh0eGs3lDhs3EVt2x4IcVpUICq5LZ6BjFKwuZ5DA1O04
MVwajpcY3LqBlsxGRE+KLb3XIOOhxuAMa4RlslavoPtzK/R51VJ8i8NFeJ9VFNa6
wgrTnblvYslYKsFHLzB4OA==
`protect END_PROTECTED
