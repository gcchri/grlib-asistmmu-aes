`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljDC2sWWg7P+7cKvpbk3qp2DP3Lj23pFC3hgcBHX0gqo/V/3eo00inKRUona9LwU
Tn3P1ocPUWvCNLeXAobnCVMq3M7ID7u7VO3m8zLTLD6i2gW9XkQ+qLbAe0Bh4Qd+
v4r/GkH89ssS1q35aNi2X8UmbSbKbX3mCtvZ9rLOnvMgBIjT+OOTARxKic2hFeoB
TQToB3QTc3JNHpXD7+KfKLoixt8/EfFWHzRrdHqrLW+zCttCRh4ff3A6vWlFpy4h
ExGKPd9Iz6LecM04IZz/1kM2cIJCEPDlrNwPrKaAOk0tC4qgl7rXwJ6N0qTHoT8O
ZG1eEpAqMiURUz5dsvhlk/E1KUoV9bOvEoRLTeT9RMghPOKMasKVt7FhcgKg6Efy
8Nqhs86LMqmwT7B8OrKXxs2vMZOvOOVIdN0RKb2BuGAxLTA1ipYfqEriLqlGrgE6
EW9ySYzO+rFYQnAZwZgd6CdPxDKVsHdYGk5e6G0Ddhyyej1OO21wCPcOWWMcigbv
qJIpWruGHABJ0UgaAkLQrXqlCDit2EoHjV/HtSeobgJiZbvE5+yXaDmNI0R3xZfp
y4PIPI8UWeL/q19YwAmtWLg9BCMgp+/AbVEmxlQvqn7vh29UnlIx8FG71pWtKgS6
iuNZnn9dXrMFFR6efstX86McNpqmFe/JXSYzNAbbwnArR9f5yjomq7oMWpBdE0Ea
ZQfQEYVdnRXpJP3bnKjpLHo04VZjS2V5yWF+rpZH8BxARLTrZ1/8A8yV1K1+occL
pb2at+Yepj7lN/1IV3Suf4t182+dsOA21w6dGv/a8hTnOd8PTSAGEuYsz0N7bmr1
mLv1jI+itvVGBvGZ88jTgXrw3jFQPRrifRWRQBQZ3Ex485kCKU4nut5gUcBiMKwK
WhzKSchKnFMDf3rwGrM1l3kAW9BsXPBNubMqxHOlY4ocSKPuU1wAh0TlU29Ud5my
oTLaHgLDOW4/htLK36aKOCZDDsQOunBDM309JPP1vHpv60xK3SEey3hRbcbUx2Be
LXYnr5RIAJrUQjiOduICfu2Ic5BzByPiw1KP0YO27MjIRNvvBilrFh23StMKD8KI
CxkkijJ84OStY1ug3Bq5e8zoCVJLlQXIL/8itOfe22dlq/n9aHXO3NtL4/4DXI/P
2I/ldABeMaEWNKUZzGJGeT8Nrm/7vFyAMP1oO9C93QWRcREx+bUG2jZHwplJtGjO
jyRPt0zP5XBrgRXkP19BBC8Z8fZfSrOlq6CF4Fj2iyAobEsMQszIOyztr8XgKvVL
M2VRNW+u9OHPtI/hMccEiq1pdnAL+jdKg2V5H7mjoykCPaxmxYIeDBPr3+qBcyPc
BQi16daZnamSU4chCmuqwkiRaonwoHFJs9sP1hmfIyrpBuwiYi7wfDLrbBWTN/W9
ijwVFI3QAScqhgWeRgCKKr/cyJGWmFXC2HdCtnkyhHnVWhHO4fWyqusk6vvgpLID
EPWdynCAxFN+EJddIa4IEUBjvsJ6WQFoiq+ea8EikbmwUyFA9RQ7ZKes44ea5BIN
38QRP2g9JSq3sQDv/lmeDG55Ui6BURjGSwRPkitgwb2KfZVJQAZaWg4MdJGkgf12
m7pB/Li4Wxqdvzf6l/SsH/Zm4DCgXzadXdmqaxDBADyBvTQaOXlc+nCQtFS+t5FC
GTBPufyzeRPqb92A2/21mMlvDFszuoqpEbdDk7tcRtrj90lzHv1rycsqTBDqHl+F
lzCVJry/C19s1dczxsXitNEgjxWy0LoTApEXGdxKi9vlRU5FxQ5uS+xN/bwDz7J+
+DWvU/ASX9fsr4S+WHepMC7LkVd2UfQF8R/7+l09COSfHiEnuOPt10/3N5bOVEWj
mTJDEAy5cfA4rjexUEEi4dUy6S65a6xp92dTArPY5CWg8WlXUcOxq0xad5JrOY/C
5UKxfA3fuJ1H2xGtsfNzjH8kQAH3CnZp9OxdhaebuC/UqriGw4dKjLOAWsAszu8i
7/Fr/SJNGtBlcLGr1lrHZmAnpIW1l0P/RX/ksKG0WgAd/gBdnwQQF+gMrFzsIefT
hIUvvtpEDGxQoEYZnkngL4p9//Zmw6ti6BjcGo16rBHbACLoI4o4pkxwFRKbuCpG
afJiWa3VEBWsBYGNYpBal5ZbIuYdoiv22FZO49DQOkCZgC5ir8AINfBcF9ep+paw
dorucfHVz7AZGSGt9Oi/LDOkGoAxpuLgP74qNxiISYxDm8LpQT7fPf9vp4yYTkgB
iQdOp+AllQFbjQiI2+r3VejJ1VgAJsjb/tSnNBJ7GtI26+1ikAkL/9e7wUktmvEs
6YKdSL0hW1WVyhpTNeOu8zx7ReN/4t0p3GeVzusdHCJs2HYx9r41arAm6caGf0Lr
xLycLad5hbxWbTuk+UMR4Lkz4BH3x6eWxNMRBe2uon5m4KvYLjhcE9ymfQjSQqNM
hvBjPjMzddjoP1rTv2xCTeh8bs+BW20pglYUGyACvWuYl9/4NiQQcXItVj6ccMFu
V8p9py0EvTVBhU+pgJTR+wiEKIrN9h5ufF723RbMA+ZKMVp/Vxoj3/Zn5SfzF8e1
D6+vGg1G41L2o5w+HqMs0K2UtnjsydH8LXLBxMN9W7FUJFVJj0ecBr4hMVH/3hs5
wcU/CNOcdsT8eY2g3pHxK3pGWhYspDeRapqQoJFGmpSRLJzfil97FNko7WcN6WaV
taHY6UAUZf4CiryVtyNN4DlemqKNd8aooazqGCzFTa/jWl/b7SgWNyiuSm6sNlz4
A783PK43jztYWbVQkeLtTJ1P8C8NL4iAPUeUiQzgNzer7IrDec+E8sott2Ho9hBo
j7Q/9JHQwmNBPGVa3gu95VMIb92mdUUBU1H1GsHCXygu4nREiaJdq/+VCXnxec8c
UDPbkFhyi5oWYSao4acgUsgzgpqYjKv2VPjz/RrVdVLqwi45y8/UjlTO+wxldGfr
KiQK5CKB6ufc48TYUnrfT2yZZxm776Zdf4KeQ9J4XB3NQWIVjTYsPWf0o8Jp9Z5k
h4KTEFzwGNF+yjgtwyZKD2DFcpGULCW3rDQaHShUwhvXc0w4TBa+F3wj3J4NHe0L
mkCuzoKrNLjwHdah9gIJq4lJ6pwu/g73gsI0nn4S89h0lbw+E+MOHgFXM5Mp7hJy
u50NjMwJG0GWk8vbGPKAmJFnINdrrLZexvIHNigZUFVCOLinIBBFwDII9sMkJFm6
v4rM+Sx4rTE1JxV09V9chgyr4jnjr5RcgCZxGi9cD4CDpBF1UrqbtuTBY8uMvJiT
5aZ73rdYYXXv4iVWfMXC0okbgMH7+WkJNxyzr3vhF6KtPAOgqgYofHQ+rVqWYjXJ
cMOZo3NOc4PwAme0XKg7VYp+GJJWa5KcmydSB+pSFvA70EDPtWOXUfOc9KxAShas
5bzYbD3HxMuOd3M6Syg6CJ+qVj4cnod0lnONx8HoSGb4WqsgqwNB8cFHEuatp6s6
tmr1GdlE+d82DCn5JzDpdc31vX5RyAgGK6Mc4NpP9c1J7KLtSLmil/3GGqrMmDm/
SLSXlxr3aZxGN8qDEnqp9LzeyRp6ZuMTPF2IAfoJPWcvUQtPVS84z9PvUrRPnE14
9mvVnvGZfSQ91MUbAzQ4DI+/ZCf0ey08dPS7GlUdaJWBXkyOfJU36jj4Ma+MqWZB
0wwB2jO4JaPvrdqp+/3LL9ti0H49TxQKResVQATffj/miO2hHDnBDKq+6oC+IouO
9+D8afoaqRU8PpqQo1RRvcR30UXklxYkXKawOTwvuKmcxXVXYlPqDgWTx+1oVqrL
`protect END_PROTECTED
