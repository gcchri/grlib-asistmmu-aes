`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgKVMsXVi5ehL0KmvGDAyVnbGWdEw8vmgPVj+1T+MWWC2FHYG9sm1tx2ePCffRxW
3p1VE6ovkzx9bX7mJglsnMar8rkhL6fSNu62eyaB06veqHgrvIWKiu7aEr0ImfQK
WyJrF2wcrAotW4gOg1m8t3m7lDp0anT1Jlj/AWymWASjEbo3crQx7qwR8Jk1ym7x
hDO023rc7IEWnMiP14WpDACkfbyQ/8hkE+vm06OpJICHK81bkz7UHuvSypUtrs1a
g2TJp1E0XCpQhkJ2ECqE99q2H6Q0GqInbZG3oriVr6Qa7y8VsdhGuSnz3+liCPZN
`protect END_PROTECTED
