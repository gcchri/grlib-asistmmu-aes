`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHhCYBJxegFtuEGcKiWbdex1v0JzkF5b0DI2R12L5oXyMZcSgS8EV4fYg13G6fMF
eDtjmEHjtzd5WHNLf/tAuqPTDT15S0di0/GXb2Flrmd4+gQSqSyFKSuhC+aCIapi
6e0fWmriK2wgl0O1vRkf41o0hW0FJ5zUGYv5fxOJItsyFBqIWRrtDNKfo0iM23YJ
ZrEgmrSxWmHbvoTVEuPVErh4vHqyhP2dds1NhfpaaMY+xAy4WdnKoROGUADJkVhp
0Eo83GiWv4/5VpS+iousKOUA850HDgmLOjn9cO47P1mHcF/fEKu5JKBhCoFXE0yO
bBtOGxwGylmvF9jCGYicbA==
`protect END_PROTECTED
