`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gljFQvIT5ve/E3TpkQE+kn/cLOvfYbW+NC5Ie0flkZGyurxRUduSTdUhkS2eAtw6
z3o4/cc+CIxkLelzUc2ie+T0BJwH+bDS3TMXL559RBl89XaPWOxkXrlsU7f4Yz0c
O7yhUNv7gBjGLc1HtieDveX+gw9+Wmer50wpFrhyjOePcv7gTICVi1GbG8+Dffgm
ICKEw6t5ST01ljEDm0OpjycM1OJ8L9zghOI3vF/xuSy6fLaSIOhQuSbbsaaKw6Oe
ZO0ZjUbc3U8qRrw+Ks0hQvslMJxKrBbfhDvom+KP3POiLd/cn0E8dN7tWy8l4Q7f
nMxHrX1flCW9GMIG6R+Bmiyt3Lfb/HAeYdzaFhBqORBW7bLPFg3occ05NoQFFmC9
qkbq8G97munJEIhmU5y0iqwJ/vJPry7DC4XIuCQfsHz1i96KWZBBZ4BM//8Eub+p
q9HT242L7W5wnlLHAg7luA==
`protect END_PROTECTED
