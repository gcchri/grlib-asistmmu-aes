`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHDm/PNjhm5KXWncN/HgLz08jwaqOBn1pmDGpDB9QxlTO2n/Az2oQBFmcU+49Nb2
Vn19t6QHb/3sSE3GWSSX9vrMzEw5dNsmW+N88Qx9XfzkxrGPehPs6ciqIFvHc70E
sSoEb8cGkUfkpNZPX2M07GGlnZan7+a4pCEDNSjWYilJycaWkxeTQjsmQ5khGHj4
HvP7I4LBYURELsZrLhjqqBL2ZQEf91zzoYG94ynuhori6Ez+VQ1sJDsO6l7GHk6U
2YsXa0dlst8GCYUHKBCxzIDVCyEl+vLABlu3wTBWIlHj2jVqwbrhVYe3VTCyxpEj
hSgYOijDV/1AlmML4SWLTBzL3QBVM9jKOt5b9SSCReQH0bGVHi117UQo22SjtTq0
YqPJNgyzoC7vY6jiPIqnfQ==
`protect END_PROTECTED
