`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MlaAJUT9eaPC8zH7SrfJ9/6/aGa8Zv7vMxPH/h6wEIbIyhxNF1iCpQtlBsKIq9U3
WbYrbbyEBgyqgzxjHxhUpKLV5hvaEw0DFWqyOqieZRklaRezYCqVh14a8BC3vnt8
JLU20qS0g5rggjyL7j04Lcix53iM5u9Hr5DdHqWQnnpR95rwa3INZNupA/Oss6CN
2ivgtAFPV741FbN5CAMYzSIXPDklmzk5gdkKVNts5osciVeb+zIzhJRhVNUKKrBa
1Y7DJbU8DZzXynRh/IvlKg==
`protect END_PROTECTED
