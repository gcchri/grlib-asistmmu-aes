`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rPMaVjvg+Jpk+7HF93Hs3EXzG5lQQ4VFHJ85/2LkLzG2PLt8+tar9fNxIC5ml6oS
Vo+oQL7REPaorrsBLLf426hgDvm8haD3c8gPGrj26LSqc5OiUm0DxlP/EIyDZyai
PKFpLJ+Xev3NYGp3FgM4xbUuc1Kz5K10uIJqTB54smYLttyGLDJzjOOzKQ2FgbgB
TbrtC/rNIjTEQajpeP/2S9GdMFBhTTODpXJwAnwX0+bpgleLaY3rBfyaCBP3M+Lc
Hc0L3GA/YbYij/+kqcqGWkann3HY2b6qt+DOdBz060Gy2UlvhuZok6Z3OshB7pDj
3Au1QE0LK7xn5sSnRs3eIcVDImefSvJnTIaq9LdipcKwYKQUR4jl1GHLmLBqmBjr
fTxvlcnh1f2BvLwhls/YRtkG6fxu+nQ35svpOWDauN25evhLfFXqE8CImjRMp+MR
oM48OrVwLSn/c0/5wFuw1Ap32hXAdO9KFdwaqoAc0OgguQQqPFPxl/zYSDBF3jg0
Ue1+7lyEzKnNywIslw1hEMI6hFM25Q7orMt/FbMq1d9567ijulnOYRHoEN3zqct0
jtvLfJ1CKUFBzwy82eTum3UOzGSVo5fncvZe9upW8Sk3umKIY64KJPCCb7pFysBu
Vso8rSmnHg39sh5lvFlz2jjOmh2pWZ/7W3Mz5plPZxTF/GSOaVJMu/aC6sroIBDz
uOsLDHCyfTXBf1NPyvMcol8aOhHvEmbZxzxlfBgetQe4DrubT4N3qWBfghjeot2i
/KDuQQvmh399rmlq1QIDSSZMWFVAzK7SMqsMVPnF7q+EoXag3zk7GAu8vJ0jodYC
o0GAUcXml3HtS9pgYdjuaJWDfGmziw7gwYffPy/671TSMIq/Hbcm6QHxwAtf3Xmz
fyv4XUX7MEMF6waAI/NMrWwy2E1oDd+92h0b+a3lF9HD7c78vGj+HrsAeS9kd/xU
01ymYwNZ/rydzDDG8RfFCgvDD/bbppjwc18y+8hpIEWEQs0+Qfc7Yur+JxuI4MkN
dcPD3LJJYLI2irS/ZA69UZKxFltowHc57me6U92OSQNEEOvDDtzLH+4iqiYlyX0n
eTjQHUStliakSWrq6UVciraHUDmPsBJVuPY3a70rbxxWTmFXe2kdscQrD4MQCuEm
tXAlouPVBSmmKCylWR0XOoOoK81mu9EI6brXPDJWPAxONKaJsN42G0A+oYoj0t6y
UDRxYxZRohFOEyEPbR6DgH1uv+bJAG/lxmQ2alIDRVHI8mgIF+WwkHDWnq11Mf9D
4G2KHj/ks1HXa6uuMD1aGxBYUtrp8e9rykqdJCY3rkmZ9l8Q7mcSeOAKnAQmbfrE
4fqBo4R7AStcK7PwxoGUX06VnzLkm03gL5jQfW39MQiQaa/RyYFMb7Xk/ZOZIi46
UeKhVa+dSPA4cjf63H/RXT4whAmR4VJnm4W/SY6AYfg4YDg+Avi9rtczkLV6xeqh
X6+FiaN8qkJxj+8YoBpGiTFVyGL1j5nhI/UpwPND15j12UJRwpooZp2/soRnZ0nu
I2LOVVQOGzd42GQIbN/pTc2+JQGSgixsM1o+YEVKYd932TyhXAVjRZ435P7y4A1I
FtxXKUeXA8pXxIByqD8Bn4kU9QnKaVVZiRMhgs3jbwDsg9SUEBcE7Za53DJ2XmHx
rRSnyaoc0Y/Rr7V9iL0GKw91HbaqzYD8VqZOWib3cnYPg4IElfZnL3qtumeTesLW
zM6RXmQwXhegDd+Hg7XpgcInawhbAhAeUQwwr4AJMipyUsJ+nhp8h3Dt25WqrvwS
B8g+XQFJTbZnloRpMGrxDQbo7zaFGuz15Yk6g5lzkfALocRkr0YvpSOQUaa+W1S/
URKljl1RqsfA8rfUNYHgmIvtlRc+NnTbzCvDX+rywnbdDUpIADmvxvCG6OsO1WVv
3ewJG8baKkcgv8M9GXmNlA==
`protect END_PROTECTED
