`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D1gyB2fN2+Snizi+I7i4aLtlr1XBs/hluv6+KfA6F2d2uYjdm1PR7ZZ/x5uktSKH
xgm8gD80ryDu1AFkd77syVqvDyvklcx3iwwCGntEITXe64SdLrhz4N6bHi6zpB9B
+73jHN/89mhWnh2uNAU31HAorA1JH/lvlt7ECzWTUA68p83edTJaTZK2sca2uwgj
Anl6fgt8PVOTuh+HDgxS75UAEpDdu3OGJz4JAHYIjTUe8KFIncGgxuwJOv15sKQ8
x2qfStWez4LDzZmd70kfPu6xJW8xSF0gAPQWF/JzoKXJqhc6WEhee2/EeMLDwTMi
wIYxYlry6A3P0Dwds/E35F8LVFXc2T9I+GcXL+6uReZ4t9oyVtkTDbJ8kDOeLL0k
FpSKM9/rh2N9BGkNB4oy2Ww3OdjsRnRAgMFIvqQ+HiOzA0dHrPxBoAzrPa9mJW0s
+8h4F8qUNnHqXj7xrDAyfVbwIrelOPN/lnqXxZKehr5j6XGCnunyf8qhfmadxBjC
JpCeoY6WNThQu6O8E2c3zGFoS2Q3hB9ashBuxJV8zVR5hAkN18JA7aCs9MdTM3mW
TJlN0QzscMlhoGAFdYQSex28pMLmpAqbpjPK5yQnveVqOgI5sMWhZ6jYlmnjkQmd
JvnotrF9Wmm6y70NC5dQC8YuqYmNQyRghYH4VlK821HK9SGxBTrGOTfQzwTs9USx
5j/lK7mig1ct86v2ezCwyeCD06WBzeKCV6C3dQ5gakr1iLAJd3wPgSb/RBAHYtBf
ZyyHQBJulKengEQr5fI+Lg==
`protect END_PROTECTED
