`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HydFNxepbjBx6QdPOKkgnakZsg+BFkyN1IHtc83jcVi5kf1gNHtGhLyrw0gcdRBn
Le7VR2CnwaSFxOUfK29YtwiG8VU5VCySz3UJ8PXbmXIuBjEGQHnP760evizRtfQo
VU/gFLSLB6qCnhzQbBxZlcH4NJ5vX499Z1NA724P2/5gOogSPUdn1FgLIJH2QsZc
odTFUM32jLm9BRPmeNb5KoegllL7QY5eZVjwQQEajFhUBzvmIsmHoPbdvkEHapOg
YY4o76SpOH6nfTCljvsv381uxqOX//lIlXOEpJjoUILo/kGUkiculz6aKdLzVcym
viRV/KtsKvUD1aJMdv6VKxVgiwI8BbqUprCJdAYqgGHLEEL1CxzAQQnS7+pQWp4f
wsEK20dL6SD8QFB0QnxcJQ==
`protect END_PROTECTED
