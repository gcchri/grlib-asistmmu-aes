`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ttdI/8ovfaLEnLMOFtdQW0TdtmqQSbeg3H9PuhCizJA8/d6j50paJWvRYXLAyp+
gXFw9M5neYMgiW0wunRZl97xKEzBVDWDSHjWKT3JPuRMyJ7HfetVBYwmNSGDrseO
uSn/xRdcbCm0ywxwHX7ST9AIuC8dqOIhcoBDuuH/pGxGCsfm0n3189IsTHym5DtV
prtHcINZY2pZgMxOUPUJUizbWn/6uHfojPJEYcLVrloQFGACWhlEm/Ph7HzIQ5CL
psz3rWBSmAaq5RniqAqReVpKbVWiWsrbcBO+YqzhrcDhVLtxKNLRJwIFjcbnTSBZ
I0YkKRAgX7XDUtd/qLDj/kHiUP6LGpHrUJXbsb1uy+awfi2zJnZpFbQIkF6hNaY2
UI9+hw2bdkHf6LNoFpa3O5gHRyZODxbSILL1gp1yRYxptwZHalzXpnHNbGIut0Ul
`protect END_PROTECTED
