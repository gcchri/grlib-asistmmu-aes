`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oa0cqFvGFMP3pySDovPr5vgyCEd33ImMnm/fNvkU3+An3/+tPNwFaQZjxbg5jmLM
dLBdCGy63uD98xYZJ8xmH77x2O2byj/GeUUNXtuvXLQdprOqCRhuTlOEUqTiIRu/
F+YbJY4f5SR/puLb5Wrk7q+pwIkglZ8DzUxKQnKQZHueDM7T84QYjxu4MoDNFDu/
ANAlPbWi11e1kd7PXbrsnsdOtirfiQ0kaYlaPf3jngiL1bY7XWQmIlaCdd/HeM3b
3mQ1hHS9K3h/gtZljkNhirFgbhpsyknXudeQsDPY7PZbAVzvajhuga/sxD+0/8+a
p5xqdjHov5Fv7XdxtLqcYmQkI4Z+7MZcfjp7oanYaJptL3xfq2LiNfwoO/To8Hx6
zAmyP8xB7USz+9D09Sc+jtNlrV4AiSeCTt3ktRcdKX4zU5e7KbiMdA0zv2LG90lp
eHEGfzARRrieHcYpb6v3DjqpIZBN7F2Ce2j6+9wfhFdtl894Yo0hqiWYRdnvG2r8
ffUhGbgVCTNvTOtN6cC5fbU2PAUzBthOcw2SvXeW9utaK3eT2EBhSHIEUaq/+RKA
tndrydka5QTgxLUUB/Zljb0GC72zSDX7YVjIBqQvO9CHNLvpd9i0o+GYb+xJtlQy
nvDydgo1FQiSCeNxAICqdG+eI8Lj7S53iGgt14vTAgMTAp8flYaiyyk+o0KjSKnQ
hYHg5eSA+W3mNvX0EJYXlwnhKqLd6xZQ8+8H59uCpRnO07I3QhNM+LbNTU6q8bJG
a5k7tvedaEPjzDGG1UN5539UqcU4Vh+9qwyi/JsGggaEQDbZi2erjAjNLSAf0BQ8
Ek2ycYYahTD1/mzdaEelmEGmsjh8u6qRFegtKlxZ2xIOCqBCu5zyxPLTqIUWuN8n
0GlkRXfZYnsx7d91b5pcJqXe8YmZrdhSsnckwSn3gqdvpTXJ30NaDsd9mfPYS1ZL
QDCsuwYE+2w5nwP8LY+UdnFLjxrxfC6VdQRHiGbKkXUR0XSstst4vgUPIZ0uWGHn
0pO1OThVCqYvMKVTu84QFg==
`protect END_PROTECTED
