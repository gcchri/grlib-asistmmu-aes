`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n6Aat/vuTNDUsNMnDRO2prAZa27Ek8hxdDpAmlm8cCOce1RBsKldapYWwXUP/Rc1
yGTtlLv82dkAj5qzhKcOPBQVnv02xRHiVHjlY2ytNt8g2LIRAEzd4TgJdtQlUBDo
/FgSMzXu4IwzdBEMBiFnygFp0Uj4pd6SR+iTy7nmGd+z4xBK5f6aVLCYU/OMggpV
5G+mPj8vzLdYc70CW4U1Uc8O6gbKOohZ1V0mMhbUUT6TqreroMOAgnHJ2HAedcti
z+Hbu9STVd7A3mCM5dJAOyg5lI+xq+3OOSPZlcQ0JQtrjv+aVdxU0GPJivjKHi/5
j1m0Hgb86NCguVPmnUdA61wD7S23SdKGWHHEVnoKLLWIf0elSJw1iAftzLX3D3A6
JqTSJ9zTRlsyJ+LPSNxaeS1ID9Wbm2lfQvvD4Du0ikhIEvsBs0jY6DHj9jAsa3JX
fwIwY44yzlsga24fasMqog==
`protect END_PROTECTED
