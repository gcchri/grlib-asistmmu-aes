`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBUNDhkEbXHBdqDG7E2jQXcrQ2HUNcUmdU0GEbAD0Ov+4P3gBE9/uOWX9H34EzsM
x6brWjT9jg7dh8riNUrdp+A67KLDbChjt9l41NuQHn8oobhj30BU3zRm4zA92+Qa
3qqpNNObGWtUTT0d+U1fKAL9W2l++R9aMnENQNlHYWonsXTgxspVkO5bcfdvKQKI
W/A2MOSvLMRiA0ziWD1JX0bG2gw0cHH63m/jPcKC+0R9P7L9U2tuIaOL3+QAAFXg
4htKROv0N1zfax6FRkBGITbo6zt3m58VJ78MhLwqPQzk26nm6FjldvNCdJARXtz8
11S2K6aNJLU/IMJiJweJ+m30Ez2Z640S/mchasUu0Fj3VFOHMJ3c43BGigm22pOI
IZe0k6qexcJV5abTPVc2Kg==
`protect END_PROTECTED
