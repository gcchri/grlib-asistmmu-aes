`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7fmd3l9WevC79rTd+SS0z05u0/Ll6fzMyiF1bruQT++mY28AS2cBrdVmFnFUnPNN
0rmr/wuH9y+cpmJgkIoCQOWtW7yKKDJErWQhjdgiRHfkiaKrr1VQnKBlfobX/c3X
LgA1RYPOmy5CHk9yOEXTOgO7i9aw4Z8Gmb4MFvgIVvUzjkmcmxC+kxZu/eNhEW5V
DVAVz8kqv1d7/5qYGRyEnbtVEqbzyj80wu8PIBAF78SOuDCDlxj5EVxjrtcWN65k
f9rwReYa7eURNo+M/ybQZvzQKO0FRMwUKOEN2x2ikSLjyLFMmKD7Q8x7Am0ys1Wl
UaxyXSlkLEeObJcSEnsWPA==
`protect END_PROTECTED
