`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9bNhjahu/ktWNLasKD65hwgQU5lEz3ImaKuOg3Am2mzjeDMOTAE2msy90o07p3l
G8klhpZsZ9Cv3zaMRwfxE+vrj1HOYvDc0ImzqFAdaJsjdbE0o6s5TJvTQpg9J3WT
p89UCDu1q7jnc4zbFb0oEAZm7KLM3ckmPdLX5PAXAWkQBYclRoPRiZNNYrhig0z4
5uJQfQnqCGHON0pXTmgBJ7m/ZAOL0LGC8PKYwYtUw9u6Fl2THJtfmffTCzd9VDjJ
fg92wZ02H2jYLyWAeSRqshBapg7KOYRVXwLkThdfRZXGk0VQ0H4B9j2+LX6CVFHd
Zac3DM03yndqHo6kewn8AdeSe7/8ayoKVsRwaR+A1QoVqg98W8q57jAzP0qcCoXR
jY5twR5UOCJdCZPt8hX2ATfE4JakXK0wmWm00CSeIxveguzlRUgtd5AiN0HWsl67
IkMtp0sxo2pPeOcAMvbD7Dvd9m6tZv8iYXEmUAW5biQXPX+yD74SYeUJ8SnnNYJK
v84Ll9WV7KZwNUfmT+6TMFP7x1PS5oPUwhF8sBxwg28kXRlrQA7ONHIodKQ6h75R
15WwMPj4vQIfwNMPMayY4Xn/O9sKJhee7rJ3u3m1V+EZ1F/CgfefjonxpG8AtZpy
oCBssOLvPZcEuDsgEYItbUQh4ihr8f1WBp1gqdJLvaXMt/5F2iIVM5tBSXuT4FJA
HDGUEUErlw/Rd5Cwz1XVS2UhcFkp0MfZglHxUJppHv+RPk2hDiObfRFOUDC8Lr+a
qZ0J9isTGrCfDuG8sKUXqeIWawzUhWF4zVWe5sLC6tDPgWQkRN4pfSdE3BZLYIMy
/1IznbvjERDd2Da5VcJOgOaXibObxD+G3INkwLKGbalC557RmIhHjJ88KCAcohox
Zd/UeHvhQp9DcJiHZ0CLt7t5K60dswQck3waTcAS6aWAtNZnguwZpIjAtnilu98e
S9mdeaWL9dJn45T/EWB+ZG2H/BXu0isQ6DT622YsEzyKQUqsOzaYpEQEan+scJqf
2B1gpgU9eI2ykKzQg2F3mddkozr/h3k5//V6iL6z6EU3vTnrJzYSu8BwfJnKvU/w
Zy1xFU4hGGObm8x0SEvoqTLJWgqtDSoWeFzAJowSpojJdd01x2gQGWOy6CSdb3zJ
odD9NNwSyuq7dawtuF6DVkJHOgh99O6oBiqTyElnVb/TwBBqVtMdoTkOGQ3i/p8F
nspxLq/+7eABSucxrxeW8cT3R+Xufj4WhtW7cxxiUaTEQKgwxS4M+71v8mvoH2aJ
MiWw/ih16B/CM9R6mC1J8DGZZxiZqppzxfLr2UryDYiZxZN5hLgedrprbUBsZwWo
2rtOTubR6wMj1vIbSeRDy0w9wD4jC6DjAXiNS1hcZbYrCo9FqflgoxXhu9EAg7D7
75TzdFrJoOaPhojJzaLOViBIjeYl65epgsXSeeA2jcLM2g7OL4xE4q6n+Vd9sNlA
K6ACCHcnWEHG5N3TIWTcA5T1wTolIB9oQnMaWGxL+Op6tlN6VKy1HwPXhd6rjai5
ocui+IYR0bZbAPVPrzAsHcFrO4YU1O3mhOitfruEiqRnAeRSCjEWcCioTQE+KzL3
SDken4e65jL+R3Xo+z7g6Wkz4SaONFeUUUnn3ifWfJF+e5xlZOgb+Gqhp0wzrOWG
Bsqd50XrcWxl8GWjNrZksnxVab37u2i4vispEC6oaHYAcXN9j1jDnU7ClSK/KkV8
czlJ8YzZ7DcKC9U+p/QqyVJO9K6gP5PEERL5ICLDpXMwbfia+YCju4MetrybAdb7
Yy1uyrCH2vxQvqYl4NxIHbCtTUwWI0eBeplzWNfbtZakp0USytHwtWiVCs/yHK3x
VRelIw2w6R1Rnxe6i+LFF8IJQ6xf3ohRm6aAQJuf4iMji6dPwwGpqAoAN9/zfe2T
4q03tGZMP9lHem3mwj7mUXd3+ItBgWunatGevaiHn+8KhVmfdOQcKjQfdjJauFuc
z5QXy9BRgE8MgxTpOCJvGL85lzq+awAaLbvnyBcVAGnBqusWS6zG3jxLsevBXum+
YwIUfo5Q6NAXTEtA9EbRuMq5OEBb1/BqDCcmxUw3IUnJLXTywyOKCbCpS9w112T3
6cyhM4aZ1H7pA7ESElZelXQfl862H7GU/HxnUiAy7l51+savHvfLrc5DrAg4WJ2Z
4wXwk2LBCz3dddT281YEC7aVLgNTDe2IOlak/l9Cojy8LAKqYXugzST9EhHSutSv
92JNRJHWVeCysQ4LreFgeDtssXrWTsx2KPx0tUH2WGBEck+f2/nYBlOvqoa4P5xS
bh2NAt6Pc4wd91Mr1gAU4x0QvklyVUlyX3jdZgRv3+dkNAIXYzkUf9Ua5XMUrSzg
9Zv9xJ2O6fQcOdE5FnhIavcQFcMfgYA79A0wbyquox+33ADI6WGoNC2HiK0OJ4Lx
2DbOmTALQ7JnP1+62imvX+sKXZhNT/aypCmx6tSfKzfIjLgrgEzidyCSUXRVtflX
7tcpZNN54oWXcQoFE5DMZ/eZxv3/gHt2R/HuqbJEeR7wfTFpPNy06nIFKCGk375L
6BupJXr38Mswgp+t6v0cOPVlKFHqeGeDSY63NXUYQ+uDfJmtoCx1+okZZwzcptF8
jchDPjJsoArUJVfLcKGLkifSf11XnNwCizoNssaAISOWHR0hnphyN4RRp6KGCtgq
y/HBW8bUWYS7AYOL2Np7xKyQ+Z+oNrUQZajlXmmWqUgqJty8NoK35sl1REeJQ5NC
auytPnThVdMd+CXPsOjii1TzpT1feglFjT9DGgH2MbZwaQ3aPF7Ey12uhVxOOH+Y
oqJh7ev6GWwRxy+8EVGAHi03+vp169IHtlopB9KBZlpZDMIs+ZlNAjkhXhQtWEBV
Tof3RZl/Kbbowh6k8rx2X1yj/OPJMu6CUQ+GAlEp/8bf7/m3TKsEMsBcTbz6t/J0
z4q86L5ZNppknq4+MFTvRHd2hLatNYu/XTHjikyRvRh0+wzVUnvYMjtvF0RYxU26
eAYkQDOP+6iWQc6VTCVg6ckgdYfyD1rXc2W6s3+XwpO6TH6DtF+boN7ZaZbd+7JJ
TQ2h50bbJx5DGZ4jrS+hvB5biaNmlAI+vi4CeL8/u4jgAWLYwGStsw6h5yix1045
opZTQcZJk446DcQBB2Xq5ul20DvdsT3S679L8BvKXUQtYA50iT95G2eCvE7vKOgK
tqTq7T1lWt1HIa1psuvToSzpjf9Zc7d0U7K3ARqL7jJA6eh2/6dWI4/BOSx6KGb0
au/zV52B2b6PzOfeTktLUA3ArHdC/zYUu8nAMzyd4kgc6uK+6jx6362sPDYgVWWB
dywnXb+I9FPJ25llgEf9YBlwmYvoeisBCZqX4rAywwdoZqUx576/GsxLRwn9mkHn
CXN++aaJE01lSGxBdJsATOjHdEnMNqutLvFq8N4XRI8Szx1l1xgOLBY5tbWe3Pnm
ArorM+d71BgxZ2BoXDiCXyMxKV6J+dh03TCV+P02V3iSlO1ZWwtSyWlTQStTPKBq
3fUnPSqgul52qYtG9OtaoSkWomlNGdj8VDn3etPyF4LcbBh7dhTfNRhwT5XoNVW4
N7v/hXBghrmfXQsZaazwshHsakhepFvv/3fhUYCf/7SeNWX/YCgtV797nISt0YtR
a18okT/NUVkMjQp+Hmpq+RhLVy4/RFjKYbe9ek5hgcBtF3L1c7FHeuCQYENafORf
KbMtvqDMCpYcwQ9ls2/3dGdcNd4Wea4duihztAqhIclfA2swR4UaCH3Ui9yAVL+O
Vyd01MLfp3UMKKN+m8rmUtTNEXolq/2GcY3Fs5zrGWU3oyHmoFr3Ox6UglEp5kUB
nB31Qbu0YxBwBd7hKJxfkH8W0wl5wUbvxrpCxhsAOxovk6472qCEZiUYOR/dt7r+
ZdwYz/2PT/UnU582oggF369/mGJlacHTMKs9cq+OKu94AEVg03h7MbXLMUKibtsI
p+uXY3dKJolJ+EeLKEdkGzVD5jk9FdOU9N85KTrw28pJg9RrNHbjiKg4O49Zkqih
o7lgMS/mindyWelgJ3BLxTwIesgZtx7o/xJ+H40b946jFT3/p6Qr66UinP0+NRRL
QQBlKCfriKV8NR+if9psWk2o9UI1JkYJr0bb5QnFuf73s3lCvcWBRLgQVLwKV0Hr
onZBKU5A16XDW1WpSupT2uwjYwhhezLH7MInCb6wCuyaFqJ1YBhtYZ/KqhIGr6VK
TB93HPwWbtlh2vQNwuF/mb+Mw/35bXAtVFfOIf6sJLYppROJbr1sprG4dOhLre0D
cMH0NuCoVAZ8LDhW7H1UhHczcQHCIsaLDjpd9dtZLIYQm5wK9QDhU4amTZpD7Hwa
hUk2VodzSFWH3it63P3FDQdkwYQtr/rAxOoIYMQZjXfY7g84afgSaGwyRiiK//p/
PALIm0ZI3et9tTnDDgDD547joODxf9ilwGM/X/NU9BpNKj7sGk4f8FQ4jpo9NXBV
Ne0RFdB2NeaJza5BV0clk2TKCrev59c4jR+SCS3YFRwGdWh6Im89z/lTyq746Z6r
ZkUjbegZIQ4F4yQFCMSwmyJG9M51s742GOCumjFE+jtcwYj6twhG7aW5BdhIpJly
5Rz8/oTq15QTcCsmSVsddng7QrEK5E89GPolUiHuHMpeIOURbCyQa8DDEicWT+g7
0UXP4j9Wqb9VLd66eabtdvxtGIEwblfO1UtjaNk1EAALq/Gg/qk4l1vat602pWM9
WQooEvWzrl9KLPxLK6pjos2OmWDEIWwyf8GYHNwtN/Iq2nWf5luCxR5DJsSyut75
M2QoRMv0FT1QTr0QPc0bljUV1bNqp+7Hx5W9XHKwHuYHOaVhQUOLmgMz/epbH4q2
i4w1ylvu7cO4t3crLec1kNafvwLdKXcCPvpizjqWiUkFUOE5XW8SsJJiy6pTg55P
JF9OhpaOUYIAue3k+jFrpU+IY83wlyhqN3sql+/cSHfF7ngkcbEAhqTxX63P9RBS
rx3K6PLYgd2rWGKEtp17DgpIhBzdNZnJVG6BkgWv1zccy8cBS744UQ8nd76rX4/0
HZZdYtkYBoBlt/TO+636RjGKIZFL66FsX/XD5AVvATWB1keeJwpQlSpROBM5I62q
NqO0mTJW+HLLdhBhF1fpgzhSjub3cnWa3GjHQhFAiyf+ZHuWSUzPE2JEfjtcDcGI
cbPK6DUpNUHyylXW3gD1OY70Vwy/yb01LVWLS83Kvalvfy2gP4lglw9GhqAq5KKW
puF/TdoAZtRjeIliDVLOOGfUscGnGA5Qde126CXIcFOI+uBYvR3v6rMsxRJ7eI2U
8JOT9idDSOtdDQCkxm4lK51bxQPJ1auHF5CI//uun9L0YCGFJuMzQHQOFa39U/O/
EOhIHFpWTpj1oO01QKhX4cYRfWwKfGEm6NJ0WuHoVbEQXKo5uL+VqB5yJlPD4znV
MpUPFpq3g8duca9NYkB5yss5Bp5B+QyeIRMmOvN+oGbH0Iv6M4yomphYsilC5YxP
mDaUja+XL+b9YZ8L4TlEGERK6h3hrZ7K0iOY9qCrGX7u2Mnwt+I/wsCq313KgBOk
2GAYT3dOSt8AWI5ht7ng0tRniHaGnEiII/iRoDQLI6i0jqCEisZiGDReqW8lz83S
7f7dZogOxHnXAfGZNgA8A9KgOdgmwNi5i3a8GMgW9EEKo8BaUhqPdPnwRF4thxxy
58piKfgMqfNYIGd5ShTkJJLJnF8OKfacTWM6hQE3Mmey/js0/Lk3E7bStWIO2ket
Eb5Ghk6YWywDYvDChzkPE3InH/e4SgNltX7I5kPbPM19qBF2Oledq9ZSVHafJXH2
UiNv49a9LEaDLgTfwdvvrWVnp/DI22DNlLAXElqoPpdRJ6p6sw8/XlPqOHHU6FXq
Pooq/iNic3qSCNyQ3T8KDNUPLkdTXlTjMRx6wJGWU2AD/dniR4ZwTl+xBDyhOWtC
8RhsTeIKxwevpZkIyjE2/q/LG9LA++UgnkXaGD5v2HU/Fly3g3gwB3Se+3tOZ5z7
DW9y98yxAXdEzrveoIWYr+4rBf6VNWUzFKighfpNKrzjTBgdCA45vQ3tRS55B36L
79+9yD7Ai45d0BDEVcSty3g6eL22X++w/a4Ae4T8bEzxruSoC+Mp2dde7I+LVr1W
BlNb81SjNuoharESEzGaaZ45cW9vuCfGAFJXTS59IYBX1MtgvEQ27C7PGK8OOZJy
VBPuq0jfFdGzUUK4oozzi35tREZLTwUoCMmH685hJO6ZE9TbPPQfDXe0+s/s9sC1
QXACMZtShyoBN45vN5Fi/mI+p9X+XOiBNMA7XnjoWQS49mB3rwluyg+HwxWk+M+v
ZSMjL1Vqd8QeUxlGuqxh4S2pWNryseYnVFZ/eUw+333IOKsuuZJPZWefxSMRMXHe
1UI1SQIsK8O0b/RT2ZgR+OuWT10ondbYASPRte3I/wNlOjONM7o67djFFlhXvEK1
T9UXlvI3WOhldgxXwBq4du4gv2ythxm+s76YeVdpuezDStHPC0jAXq+qTpI+nDeC
YEyHZw1GupWF0J+MwQOLFLyFtk8ubFkXxgeVJP4G+K8IFl26cnoJV/qSMa/48Ox2
c681qNKE7iXliT58t8CkEQVryPqxl2oEjUr/83dYcj5AsMRuGP4uGq9XaXmGhd2K
xrTFHDgBNd/sZhz4DfGKINlujTJCYkk7Ig/QAqnaTAaWQvmL6wEkEZb6DfXRTo7q
+NPgPtKsHsxHbPnUrE/le4CIT4fCdlexBi8aN3OLShfUrz6caL3Ro+ms+DF1aiPJ
sBOqycF+K9/ruYHJcTmAqbkdun33z22keAx4xQ+N87tkMvhiJHMtyWuYwcuDl2GW
qYT8o0bhfc9JsD46LVNXjNovBt82hUPbhHUemUDZX58Nqnwav9TXFwiQPeVKns/u
BKNDsV3n2LMHN+sEPlKsDfYb2PmBl5MxjllT68BtSPAYHQb6YW+k1Cu3s061Gk0q
9hu9jY0lgnM0a1YKTZPEvNO2zJEgVlNKOyM6ix6wlSQ=
`protect END_PROTECTED
