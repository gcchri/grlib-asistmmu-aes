`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qIUIz7WeSa0NPsJ7InBJGwnZaug88OofWLMp3bMllzz/wkPC6HH1BTjqov6t+u0d
KbK4kLkL5McNNuuQEF+2Yz6o0vnc862pYtSCbTR9Jmf1O+JOkndRZxu5Rvektpju
T5mynZurUGywQIqtU5WuZA7Sjw7dwM+5sJcnK6Y0rJ0YqTXLz6KVz+ijSTP4q1c3
7Ev4XYYe+MfLjDqgTEYaH+EXBYLSYaRMms5udZsjWQHAATX0qDQ21AuMFiLSr6cK
ZE3VjoaNgJIMqeBWeU7IRJCsk+GVYWYYzEf1H7GJ5JVna4BmXE4tQUBUJepUtck6
g8FguXaHW340/bb9WeAACuyI/Ok7iNw+qJ9gaI21sPLJfrvd19ZOrGVVIufd3h6v
UNQVzQq/+8GThymqFa3rXsgNxtVBFiWD+8awvWik+UU5piv8iW7cTyihB/BCRqxb
Ccg7tIvneFsjRbjJ3bQ/bIoF5zLHJkmVH1Ghw7/HX8vrnSP9J8r7EzFOZ4tm/NgT
RgJmEYHXtF5vlooyQQvgp9hcy2caGo5D1fflWdNyKFn51abZs1Rw5pfck4jT/bJd
q7kI3DTczM7ggJTmKUU4IRJOPFwOj7RHcD+/AZUCBnbe1rqBqmWfNgsl7OGLA9I8
ZqkuFFpmLg7d2N6BUvr7edJtEpAvW7D7s54a4Du+PbbwxY/FWv3FNoyXZ4WHXsPj
EDk24FHM5L9GqrVopaAzs42d6iChl8LaNTMAs69JQELQx9DcRnRS3f0BSlLZB7O8
69CxzSJhototD2Nmp0JdS7c2NzH1ShZo25j9zauQEqxy7XGQ/ZKa5TKnZMFEW6Kp
DOgpA5hYhYwTFd5Nz1C29eNr8C5r0u4oxnVNPlgCXQcle5kMofjpmZJCXEF21ZIG
yO4GDVqMw+e8/u9UTOLI3vxkB4WQil9OJJ1FvkNNZN6fwCIyIPcq6qdClfyfMcPS
`protect END_PROTECTED
