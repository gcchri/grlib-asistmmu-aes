`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DhU1Wc7h3yNPwpkymZjHuxBO4hhSc57cMJanKWPnqlCm8LQezAz2NzFA2yxP1sIV
Xrlcrb1GA98DceiWSeIm3x/RP2e8nK75Zg8LiWP9LF1DzPtDi+6wtjHQXvafzLYj
i8tGUzDHsH90BR/JkEmizpUcYi1iKApgQckLh4xcLMVlDN/2z0UBwZjzfX9HOP9k
0iro9N8Qs/TqXomD7+nu0xiyuFnvmFCxdqz44hRk3hFJdE7OJcsBttzMMRtwCoCs
5TYRTS+ACoz/NczCBHmB8DsBcTZ7YCsKiQL9zqKUd4fk1af+KKUTV5iJISRhdCrR
3ESx1E7Wki+Gt5J4TnY2SZ2mfqeTIRGzsNOZOeN88NzUAflmzKkP8kRVOvezRtNC
m+29AzRIqXdta8ne91nRjbhuDNFa4JJWMqgIz1+9ucDEaKaT1jYKJ+4rdz6O5kTM
prIgcAUSfx8o4JWzflVR4zlGnuz5UYMpQtYoR8MimcZV38WH3XjnIv5rqlc6MJnJ
DWcB2azWxUV8fGIeRsXTjUeIUEvznUsSMAPXoMWE39o=
`protect END_PROTECTED
