`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UY+mUEbUw60WIH74pP9ihYjBgdUFhYeY3G/xH/XTOrtIYRXKIagu6VvaggYMv/VI
TT7bTRu86sFyMsIlQ5gbG8UkoYny85Mt3yKV92v1JF9bkurnKS+AkbgC77OZWGwZ
QnTgnHKfInSZmTS1vQXM+qt1SkqdUcRTAVTloCw95R55kDnqCxdXIn/LHvbSVh0i
ee9LDnX68mAKNDZ2w+o7XfHbymYmTaD4j3cx2a85lO4d6HAZgi8JMOYgLzqCXWbn
Wak/4G3LNcc1EQcrA/zzT9b0GvHX8AZv/rPC2SAZUDA=
`protect END_PROTECTED
