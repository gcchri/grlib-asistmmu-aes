`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ov0MEFJA6wcnR+HcuqDs0gz6HsY9INGlH2g5pHl9V7DMEhkQg4/RYvQXDbybKMG6
60y83nrhmXaJ/3G9RdK7Im6Alv052oWdVIvFAGeV69r1/JJITpl3NsHMBjwlhrQn
3RACJx/AGbzXzqwVV1u/FUudkv6W3hGVb3OFgeIixL4K0D439HGKxxla8Bb8eBIC
qFJfv7jvBtYOV/ucKbaWpmLLCqG57u4VTbRG5v4O1B1QHSsHeeNiD87AMxbyA5ic
bt5cYm6LthO0bGiS77wp2AlaVBRnwvme2UEaLrTLExTTHZpMEyBxy841Of3KAej3
YKoiHXrnSkkFZuicK1iMT+BN2wN8ZSQIpNrgj4s9kODZLoljK2mpEbR0jb+JVb4O
TrsjV5/L1RfgvH+EsXPx7GzG9kkx0HIm+gYmFf9hYtNs/zuDJNNkLF4hi9Cq5nLE
v8sVSvJ5XliF13U8loiQX9DWMlBLMI9CCYGt2H+sdNFrH8YVYyByY4hYpeJoQc8p
7zm13T26Mz1FrVtgmEAGwJzjqusMSREYMybFHg+ueR6q+lsLAQJKVkn6oNmRdxJj
XmcIPo9nytUM909WEF8+mfGArSuW3w3ndPVH2TjkKAr2aZNSMl11EefAkTYJwmK1
/kbd83o2fFkZPSLmK4BqqzGzJ079yTi/kMtSF57ub6PNvyxQ6FwM2sY4SMaah7vI
ziaF9JgWM4ZrxbPF03FCqkJBCAEaQ/PQP5psBkCYbNzrcrik1c3YvLqyv4Zw132b
hDXuykZifJaQeAMotvHQ5hdHzSwLRxO+66ljFI5r/Xj1pM+3LJzdMxUyqYcg5Z55
lYQiGk2NOrmojnfK7Z3JVtS/cY1ZZzwmFZZ8/Y4/222HevLcGR6sp9kYPIFT+8Nk
Je2q2CExZJrwZDadvnHDQaYmB7H3aXoksOVjQvGakuXQpCUEbhi7jPn2yJHIF3PT
18nCuqxnSHJVZwEav9kxQ8s2UY6oA4KZm3L8WUf6RQHvcfYDOl1UHlNU9/xsKx7f
7BedjZHRMz4WsvqHnOrSOsVRcv07frCbi2BRBkPnUgcMy4IirkJaAHTdbnSxU0rP
IK3Dcf4i878XmLxNes+vEgnFrLOMIiCbzqFXCmgqJJzTSqo7G/4lHbOPndhgGuET
bWQZMYvBe6LdrbDBhXj7Q0RUS77jWUR9vUrZT2KQHncZ+gg5NWMl51veOtUSjd3M
jCxnlf/qPBbikZCCMkJLd4khgtBP57nz8E/NxW6r4d7bLFjsC8TAdYg10M4uiiOc
iki/S9QevXuB9HpdNV+gJBTTwLJwGiElSdONPzWeKEr6v/ogRbVlyo7wNaDlfe6I
UCObzfj9cfBWRRlI7BN6/yhwzOnCQ5rrgnITBFK6PU5VsuWCv98TnJj+zYf7/zI9
n10HODERgYHpinkdfw4HPSpFoxDerIBuKqb52X7OHA26UwgFKWNp+53yOgZs1CEG
OXiReToCVBbtqP/W7f6bC1FnJUx60ak6w9KNgNq+lwrzDQ+Lu4RcFbbW2eYIWTC0
SwUjJbgQq3jxLjWD/6ZbzlfC9UmtYkzNoC5Wj2yIxYkhGfK7VnZM3IqJ/Qh031Zc
D4wAsBrDz8BuYT3YmmzNYVs2mCK/8iwArBSeIZvi6O6n92vBG2vxFsi0H0XxpEM4
i7WHrbxZwJMiNroydBDw2bNdc5z3Q60i/OW2lLgFuAG1xqWI9ANC0zUaDycuzed+
eFMU/59/rjLmfwPa1HV5DCYYnrq2sUSo1aZ+knTSbpa5xEsl0cSoGj8Awuwx0Lqp
t1zKKw9Ip4m6239UiV9MlKpJ9FIlQb5KtLZSxVmyLJCJjeYh6lhFqWFhvWLXquhz
miPBqK9E0hCbVPC37SDlx145AcprtR1g4FawBgR6oW+QqawmWWaEc5J23kjk0aAN
JQd6WhC4utqg1h6HOk/eBjrylqn+SpnQTSM5JTBkfDeLvlNFpN/qj0IK6JCxgMZh
3WLItwF5t+RKB1WBhrbEdWVGygf/bTp4KOEsvqfVjn6CEiUD9tekJTV9Go+b2W9V
enXA4nEZ1l62DRoNOQvitv64NQ1EpgDKr4gfW7h5Ce3Y2RTgt2Asvoktw/nF2dEc
anUB8uYtIVP6TaW9BjtLXm8uGi5Tkz8F3svt3OmcPypYo922rG5Ahsu2HgtpzRXX
nkrfHJWcbRkDGyRtRpJsRFB9dTMrT6NWPAu3cG0yaAZz5ndglcrRB9Mtx3rBCuAz
`protect END_PROTECTED
