`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zeY5iMFqTzEZRIJfQ/okLG9dnorPJAWkTJglX6/qC/H2bDmTgLx+bg3vzopeXcQV
iAybnbNqq73GILfq6i9nNTXvG9opGVKHx9G7PFc4T2FnKvd+timlT10JahFq8Dp0
cqBSBu/p44Sqopl1fGpa8fBqDGaCK0p4sZkzgKnI6wXFIXek/tXUkRD4bxNEnr+S
Dqgz+W95cEDi0hcAMahqzZC+yqwoCXhmwFGDTsfAqPzdwmBQHZwZjiRmoWnQQTHR
AacqordGJ9QHbXGdVpBKm+lIbqEsff0UJVFGoO8UD6ZRN9teVbXMH8gFpPo96PsM
dCstcKhIbTSsfrgEtJ2LdcwN11pBcNetLT+83uvGj5MOcISMjf0oG0bpi70lgpdO
CHTouVvCKslBWqS9UzQmZ077DWpGYJJu7OJnRgUYyM7c2n7GXmcwzx+OhW8gCycP
gXlPC/K4ilOGkARSoFo0lcwodw4u4gT7f7NaDmjcw2LUOI8vRFGjwi+dFiT0MuDL
AQ/8YfSTSDiFpJd5YytdcmNqL3k63MteIiVafv+ft6TpMkXNjkzsWwV8oeVlDl3I
0OQUS9Ujq3TSw0aa0Tw8hv6qAkYFR1l95E57B2yUDfOEC9Xeg4/98nr4iuHV1NqM
cLTMXPFsZDMExfm6BUKspKoOsosYAldkge3Yrw2Szksl5T1h/+6v9HFCr8noqIiI
Tfown46jsptDgPcDhnunyREjx+Ic5EnpYozNyfuz+Z6uCHouMQ5eKyaWreNTKv3A
QvPgpxtWtPDyBKDYH719gY8OARDjLIMu5TG+i/NzGWUN3u7drpWM6P5da2E2o1Gh
/92tVg3LldcBU/F08nZ/h8OdHI3gXv0st3+x4gHWpg8VvzOi93+sMqWAQ8gz8nmf
dfZ7/xQsO6HO7a2Jn1ommm46Yh9X/Qtxxttiw+yMcH87FwG2MGHBaRxeWaKOE5qI
M0NbsvZFuXosBQPOW2BDCdXI7sKBsOiRuWTFpQIw0hgefvANpmb7zgSbcdjFmbT2
iXFaJy7YqUhmuMRQnJ0SMrw3BipyE4rtEBo11YYX9ZfWaLOj18LDqwG6a4KLupdG
EPtFJE7dN0GlfuMCrWwwwBHGS996j5e3iJdgx6yes8EHLPgInUdlbK7KTXrTXo2D
1YVqUmHwYEpXITqQ3j1Wj8nPxx7dxTkhk4DcgrasYW0vjUFOHoFRP90WChkpgGYy
VDTexivuyC17Nul6LMvza2ighrzkhAVHc5QoAQk3iLLqyFnm2/gd1iyxOBQvF2I6
Ukenaczjyr6LPBiwUKMA+2j6ei29xCndVac66sVMhI/oxcAyFkZjNnfDGUMcmHR/
NH4sAFFZgvSCVkeujI5pRITXH5gDR0hbHCrE684OdM1Ilp1CbQtY1hP2Oq/lhdGr
w/q6GrGDPUvixNRK2abXQC0r6DnfJSHyLIBeCtUBdLTe8rSL3FhKXzvf9w5qxtLJ
gTxrIO9bF/KyQOFQDcTQwfKM6XSg2HtVGpGo0HTIlfqZvO+4gL+1/M1F3iLOJVTN
8mB7o50v25Bp0TatmVHBH9IXcPG2UpfHuzxnx/LpRtqGW8JAzR6jwAqdSVrlza2d
QfbyLZp53YOLmSSb/q8rYKTmrjSMoB/umlcWAYo4+zdJwATEKFOnzNoNB5Eu58QS
8AQEGkN4ElEJ9W2oTOw56XUtrzT6Fh0bq5U3l/EElex0lrHVfLKxkvOYqkiM24MO
+FyzzakYcWYirQh/ug8USJKKvI4uJtJw2hiv/sUVG6WBLAjJVnk0u16MJg63eF//
PQmQ89F6UkBVlrk7ZzUYeGAXHuP0i22tJC5PpGzMWOKx76otJRFmP/eooc6trGBv
mScBQnFiPceEFQ3BBIekTGG6br1WKk6aIWCvGsssvmP+jkmDnYf7fiAtGGVP6kgy
+WwIvtNRzpwQuda/IzmAO0RtEBG04XWYvtWUKWZq5qTlnELypwE2Mahpmt6h2/qm
lE+Pxpa+4mW53ltZCjj88LkN6F2WY/UZYYlBocNt73G0DSZdJ/N7g90oZNF525C7
/l3ujip+KNwnw2cy+MfVVBxZuet6xDv5qnVvir4rYKP4lAWCbQOPjbdn/yR3oOeK
NHGEsg3mWqdXWSRiYgx3uET+fCCYHSSuNf1OPd7oc3oUsZVdjeiXfWcTJuERUtAI
/bK5CYIU5J5jJc6jIH+gXSeHE3QPgtm1WZQeIkP1woJxyamEK2KOF9YNpN2eJn5I
1TvYL3V57sAOWSg5S5hq+3XSTMIH9sn/+LFSyoJ0bC0wcYR4HjpOMrayW56F/uAc
74DqbRVP6wsS7bU2Fg1eHObNV0yqyY8sCmIu3xnF16Y5UayAag5Q6CjSmhiFvUVA
9DzLyh/D40oVu/IVM+mv8B5h2qDm5wbCN/O63s7mAm+EruOSD/w1f9WdT6iv/Yro
xYe9aN3T5dk806RODAKQrsCz2y7z7PelSfm0fROa7hQPGoKZ8c8NUsut32rd8auC
0K4PdvsSt1N9PdptMn5igv7f8dWk+gq0GTeQpLZv/L/TPZIsYoxz7jT4Y/pPkTxJ
RSyhkQvBKusBWDBFuq1877sVVrXlDPYkZqvjScLQHB0EZpyPdKvyarn2SDPwOxGU
2dMco+Y1u4TcacGBONWI3w==
`protect END_PROTECTED
