`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFJOGwKK0JD7gHDxqp1ySZAbAYS0izFqWVdyLH8PAncFGFrVj/BpFVDiJT8rIQqx
Zq94iO1WpLkShSmNgiyhv7ysjqiXrtDvWamnk2CONccKX2+QsS3KPVe3toKwPNmc
+F4k0I0oMSetPNshR/XaW65cHOf+JQ9ciwmGIi22upvpVtWDWW0dmNXxlBKmCLyF
+RXhCTGcMgiywhX8vwV0MAD/MDdTpAs0PTtqtQNNTioETiJWv0+rQMmwuwzpnsQf
djptNDKBKC42EBFlhIBX6xdtFlnxhOA4WRKAEAuQ/U8iBeQKcjOA9mkm8gzPcv93
hJItpEP6aqXc8Of6sHH3Mw==
`protect END_PROTECTED
