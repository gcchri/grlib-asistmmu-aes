`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16iKc/qK1p3cl+xDa0HWYuYEDkJ+fVspdQ6BdmIRGKokGx4o0o3CosKqhDVGYAXy
7ifA4VvTeh473KP0klzxHP/D+Ns91pDeRB5DKQuTzlSd9NjLg4qSoiZsCVHBf35w
rju8P5N65oB4LQKCjDFsmhfWYVUIuN9lAEQNTLbDftwLJw4XDyKLE3TpDTzwgHs/
UIHZNosZq/LBtVZCebdxoN687nqV2bGH6CgPoSQCngONomWxUu+/Ll9dLmaqB2bS
Mn5eUuNly5OVX5u0rpe/D9BIb+9ObSN/xeUqigK/aQbr2RywQgA0EBHfZMEJjyLf
1W+Br4QfYnvmTvNRQBIiBA==
`protect END_PROTECTED
