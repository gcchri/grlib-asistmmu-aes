`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dlfjRWXuh1IidCwZkVwSWo0hVvxEuhSjF3qaPXjgEzRQk04Ut2/1UkWpUj1g0chZ
/gQ88S/38Ti6jaG3aP5hv0pJUhSgMZouYbKcm/4Z3ztcWckGzTzg9YSPdo9dFjzm
9hc5u4X6UEnpUG6cZCpOXJM/YY6Adls8NEPsFxyCuEiy4iGnK+RIxokFImTERTmM
v7Z9tTxkjoRO6vTXm7bGcGMlv3j5GCY/sMclTaskzRh8c+Je7q1QBRyszlWs/tX7
I1kWjDngmUuuNlCGcH3NbWX6+rtiu3sVfIp6TN6iXlAgdQNOeHINOKO3pnGv9eIJ
CSLWq8uAYbeTn9UG06A9aAZybXS1fTWrmAZtoQJfkv35SbsMowYH3/nu+6R3Mhnf
H9y0LGFCQ8ijcEdAA6cyvNtOcCXTMgCszI6YpBwayDQvcPhdnoUP3igyiuoy3hXB
nQwfWZ/Pe1YO90oJnOaSfzWhFerx/jHRbGt+n2tDY0DFaXxVyM5fFE5gXBUAb5Vx
j7saS0ysr/PWn23qK0+sOGAjCJgPJok8Sg7S+SLhFD+9HQg2Q3o3FEmHpwFtWD2T
Z9N+bA746R0F6/uZOf4Y486ZgWLs0/MvYnyDUUVQbGw=
`protect END_PROTECTED
