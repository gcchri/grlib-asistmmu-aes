`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDI+YIFvHHJGUZV7G+/vwDJwkPMymGvxCYWF7wtT5vf6+Cac3zlNzg26VLIJKSOY
J3bcnhbIkBexpjOZQYAGfPhwN6jLfOaF5zX8lZdOcc+8niUpcB5m0sRbe69cd0Mk
SJI0KzpJbZUoxb9E510SKz2QKWlNgiET3ZPqADE3dmToQYwg0iie+ULJPYBTWzCL
uYTM8A1yosiRSkbuC53/b1UfoxaOPd77HxdIvXvACAkXjQEQX9qQzGetJjXiNPN+
BrUVYa79VOmVjblOnuvOAtbHsE6mYc5MtYhXMLHl2RLDqO52H9V9DhiRvrkj0Jk3
T+jf6CJQCF1HMGTyJkXL09Ap3j4H01DTWJEVQ0kpB1UqdpnuN9uuO4i0Q0Uyqnbr
ZML99Qfb4GhGQ+mc+MLNUoTrbPs/8HlAB1aB4hqVCw1cRHwbsd7oOTT8j0wxaR0C
4+6wo2WlZJYuk+EvndTJefbqeCig2n/7pEIRNCW4ozKXP7EYTWa0JYIj8KExgchy
KlrpxaM/NvpuVzbcVMCW7R79dbimRkhrw4p8Hxd1oL6YZmAbFdLEcJ4MDIFnIDTP
8cjneXHEvXvF8/H+O52278t8GT1XSlz6c2yOapQ8ReZHdWY2vSLukS2N5M3fZx75
AWUdtS4VsAo4R71hGlA70TSryKKPoGHBhQaeIlMJmfR2+vqB7GXoDMcfiZpVUxUd
wbOEEw63SXICYY8PgAMFdp40LGtLFPM4PHo/a7xZ+Mn3Omx1wzZA3ndqrNDFSNI6
TvE7xY4PH8ONz1hCuokc/NLQcJxDxApGBowJ9K+UJxoqKHkoMQa9HOBgnxDwfjjv
1OZxUVifhR/vhuhh71x0ZWdR8MQYFhHZP2pu/UJk/PKBUkPT1ZnyrGTRpHBK9ciI
`protect END_PROTECTED
