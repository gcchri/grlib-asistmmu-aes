`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eDPCjgBtzuaOGbC9Xv1ZGqhl8lGA+eKIX1XU0BLBNNP1SCPNn/waFlGBVtXvlDsx
sGp2A9x+zbJUatE8O6Wr3McFnPsVY0ifXMjliCIwOC8ZI71gd6LCqXHBGeezOD0m
Atz1M3E8SHZGqb9zqRiWvRxh0v8iKipm7yrfu3w9VYTHbYoF5u1yCBegODy1nbRe
gTZuxY4mp+2/aB+iVuHMf7zY6PDGDBYXp0w9Yk1aNVKWF76sptQrHla14nDQPFUB
`protect END_PROTECTED
