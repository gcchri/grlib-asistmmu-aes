`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VnujA/AGiuVSWLdVHJxxJyKDv9cTpCWFJZupdKkGHouGTm7015Uc7Jnm2NrSq/TE
V2zgynV8aycnDnQJNZURMYOT0Sk3Ze3pvegqsA8VuRvDVbEiOS822+ccKPukIdFt
k2v0aKtg2xO/KVAwS21j96IjvAJ3oaEHTKG5OpyfT9MY4IpRSa+bMdSPYSecQBG/
TTAHxKs0kSWZTXR7NKvQYSkBqCc15BeuFzoxgT+RzEsq0GYJvB68Q5ZBeqltucrf
7QA+jqtV/bb+xD+hsKw5436razc1TJKJhdiu6t6T8LacI17BRtUMQcOCvYaKuhdQ
LL3HynXisIlNKDQGrQAhySKTu/fuLfgZfLuzEM9qhcIUQr882Z6XHJc5OElzHLQu
FMFLjaIr8DAKbDUOq2R7yY7+bZhPD3r/I+MIY06sS/uK7fweAb5zU8Hl78IaSP2g
`protect END_PROTECTED
