`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XhU1OPpKO9Vtw1g2YIK0kP7I3kH56rpWtRW9li9rINZ30oPJvDNweUmTmptb6mkW
wox4m9NTJZrnyxvbAEDasQA7r5ixo4yMYz/Cp9QJ0taWis8ME+jrWYNtHuwh4aZP
uy68/+rnlM0A4uo/JCi2L4/yqTSX56dZdydwBIZsd2nJ+7lpKUyG9fqfpFvKa9/u
ctSzGFE9iawbpPRgz9Bp7SAet0mthqwScVBFamoVmBsoSZ4TELIoiCNIXBJsUTul
VBQMKKYOOvtc7UGQOxkGOQ==
`protect END_PROTECTED
