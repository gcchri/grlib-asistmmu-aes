`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1ycHrehNm6wHYbQp/yYZkJvLUBnJgGggUhKXY8p4uCRP/S0m5C/lY4xdglovZ0Y
fbOO+B8e5whHjaRr4cSamXd457/YztWr971TV42CszDk/a79OwjHjzK2IAe5sQ3B
ThtPfkjFLNtPOSHj2qy16LCr+KggZKbL9SPXeg4HFSIOgeYE9YUDqbjgH2hBqBdz
rEMrPq9MzL4ng1Etiq/ZGjGc+swT5CVIjcc5ib10Nhj/MjMZ8aW0kFARSrk/X6T3
J6RxLGExp82FhchEK138csP41wgUsmty3onjMMCu8+fEx8G+oeEG5ubM9p/qDWDr
R0G09efe0vNWIfkxUcGhk+SkySRSv3AvPC1qZe48fjFXV0uRD0j3/hdF+dlVpsLH
MeGNxI7cQ6vSGoDPFicRyDmGPUgeqPeSNAbSjje8JqnDyIRaWyEvaVUxOjDyDikU
pW7lAcRo0rY/sAIdRSL9RPVRNPOJgerx0xHZPsUryMdMYEf2Cjz1fVd5Z9rUn1+J
aCmOoKJ4aPRWD/Mqz4k8MwaHS//ome4wFnNVs9LZ5+ErfP8XYw3I7tRT0FHtnVYe
VC8NukycLTamDJ5P/htjWvSX1QzkuG0ZMw2ldt70TmsSScgrQt/IaNAEVSeeyWMn
UK9r/478alLEY/BUVAcYnzPDu1isRYuZqcOk23Ts7rn7al+rBe309W9ky+0UA2mr
q7NJu29WxPlS2er71q8Lu32YGsgopIokIebx+0rorBYzA3Uc/4YXOF5QVbd7ZmEr
sKj5BpmdJzayX3YL3i+YzVDdygunGHLDqiPMYlCiJ2yLu1/EV9L3ecl64PpD9V31
RDOnSJ5X/EqllIptqdTMnieWkvHKk2PK580innEsHsFeDU/W5ipA4mk2WEjEq0As
SYAEIptqmLR6Qg7R/I80OChwslV7S/GYF/2oF4pvSK15NkEIM27JpZwdB8yIq+ff
2KJr/rGHGHEvEa1oK2COdS5UT14+css4aa5Fr5GahA5Vw7xRSMSr9cniGBJ64x88
ddtNPwNLrIeDHtDTHJOkGS9Ed/tPrMC1vpBLjsHXh4r/KyWv4ksFGu2WmdN1raJ7
oN151CGanHyoIH1a1TfLCQJaXtAYXUJ/7bvhOX+8UC1EzVrxH/d3dohK2leDb9G5
+kOQfmNy5VBG4dgzGCdRW/EKujNxXJ+dOwdQJ0PDCdkHSy1trOWcdLQ/0x4AuzQT
Dcmn++JvFmHMYIHBel6UFFVac7c60ufJ8NME0+ZaeIESHH2zSqP0Pab05ufbIMZ7
1xG8PAz0TmC6tHMrl5dGZQsmoF/M9aHHrbXbah0qE0hOghG5BvsrVG/xtEGgCVb/
R0JBkxpUtNZRGn+M+aB7LSElmyzUtlnW+JfRTevxwiqS7aG8PAjzMTVtJrG6lfIx
A4MN7xF0PXkgGYoLpjDb2EFf28zahd8deoLrIC6SAqT6Xb66mM628RabqQ2lC+4T
aTpuLr6yu1Y4ek1vs4ujlx62eHLZfUnhqx0MwjsaEO9657zwDxDlvB5NF11LBLxS
rLkjeQR/Dem6/5+Z3PswAmje7UzBx5r2IlWADrGlVUxotC2XYp4ik10eYZxLbb5+
bsxPHfwBw+fPDuKjvNkLw17XO24EoIsgTv7EzY41XTQ1GYQ6qbWtluoZGYfwYAvg
VS//D7WU1oZ2G25dFxDAx9QXQy22gSIsw0fIsrFszLT7vOOMFktSWsHVMDM4EUu7
hCNu6XWU9arFNUzbVfG9+kRZdnVGZCsj3GfcRas6E3WnmOEFHV9PjikOLV5xxPHi
tOhKk9C3XbTEp4fNXN9yfrx59z4/hBDqOJ6AAo5/IcOKGf/RRVt5y3s7W3sCW4jg
n+viEglmmWjnWqni+WAByE+/yCRqNufS30BJzohvrDcIYH+eXF8MfUsFH5B5/TlD
jW7eBS5bj6vSnXD9lsZIwkuUymSUalJg7iYIZlJ8nm1jFBVbO/Xob50ku2vHetP1
JEiLPqYhCaomgVWVGvpRLaK+1yvkKXazBcXMdtPw28tH/CLUar/tDSyA0I9fmSqD
M+RB+atu22Fp6DY3VaIjzGLU/UbnOJA9eLnWWtrJf9V28Y8Vcw1z9CsP/5NIeU3L
NCfa+AuWQ3lMSC7mfnn1ZX3imeQr0U+eR+7ymYP+8eNBrGG981jGAzCLqfGgC3wS
jz7gIfsjzUsU/a5WTyxTQFAfDFVzqGjd7JxWNXFVq/V18NC3sYoffO7YAnHZW8wx
85YU2jsy4UqTqrg8OeHZRoQQBs4e5xnf2GlGBn5vnVrsy0MUIKh8Uslg7EOf6lvc
2sCR53ZfQKyXvOuCn8J2JgoA3br3AY+qOa2nnSyZydJmmP/KAIMRzFU2970H/TeM
BqKW6Vvq9ObGWi9DKnAnJpJFGU3B6OlQ5aOG7espdqVsCnSbAAvwAKyZWR0KKjdR
VJlZCKCFSvYTF96alQqvAWPNltkqK/wbDKxhrab1UtkY0GQgxIdHgp1WM5PaKIpZ
K1dEdEei18nmWTVau+V6A+aBtW9FHpZvHR0eVuP0BzPf2DE/Id1qnq3BXSded7SH
232KVT50eGVEn5urVOIRy/Ucyyo6COzB7Ubpu/WLAJ6pThKJn7aegJQmWG3DMyT6
Y22LJKYiZsTVx00OFgGW08SkV58fSsnZclC7tn4eZkn+RtST57P05ld8KlKPEP+W
PJaYFfMSA5fEM6cpg5puHwrpo6RoaJC+LolrROFivhJPEeXHjy5T6tCPOFcy+fCp
I7OwZF8AdpgvC7sYYgt6FVdakQHkNWFzNb7p/Q0Oe9ROX6KXmqOCCEPyUGrNRW0x
njNm4E0yB0PONEj5VVTImFmJp7LKmC+tOscHX5gvAUS8lBUp1ApQsOMJokZ3PBXf
r9RcdhOUNPXYyuZ5EhtuTEYV/4XORiHVNm3M14N4d43xE4G0c79FOlbGSHnxKkMn
cxVm32n7AEoOD+QUt4czens4vkQrMO8ioeJrLWiE/9xuuGrq4woaOFXy3t/iZPmJ
IRzadJdHsyoPb8NLCtxzB1cR5PbClf0WMpCas6dH3gtFd6nu2meb8jkxhyo/Pjd+
9469HmQqVytNRMvM/+AckiYKKjyBqMRcdKY/j/IZqP1ACs65dIEy6kD0Ijw/bzeG
Nx3lTyLevZ/l4Wp+mjTBuq8HjN8b7WvkxPXENrnSgdvWol1j9NuGHRxzJVf+rOfx
KVXlv7KZ0fnL88gc6uls+bYqBmNgNu/idLikMahN2T+aJq63dWTcxpSH/ufD+S36
hEwyqYv/XM5VDOryIHT5Wvt7FS7KKje9GudwH8UjEAW3OysBfzyhi43WhkSFGcdQ
hY6Nt2DY6zFVzEQjyfRiAfzuGxNgJbXPr15ivZbYv5dCSQhhN7KSu5OYJdpqsE+x
TABIuWkRG2xqpwR1rAQvR6H3T9kQcx9ids0dbkF99PAof0vCCPMNJ2DqmI3E1pwe
px0YCWpdw8/rtUsrcsWmV1mgNVNcfVtCjQ4wklKEVE/ta52WElSOI3fWEvlo2DhN
OyrF3WNRCj880n3p/APUzaIr0cUiXoh4+toy34pECqsk/YtHQZiTrwHb8R2WfFcz
+pN9pyelirMkmnuajrRu8RmZ8tId5etJ/tk21rvSRjeUzi+oAsKoxIu9is/SPInF
mpLOTLoNvUFbEoesEhiqc3Qxl4wiXByO2uttItjxP5G8H38NM5Jiwsw7ubUzrEMw
D1sOrc8XWDnuaOViOJSqo4z9aJhNKxZ7NaqOjJzxDP1PTKT3ZA+3ig02cjb5WR7g
pUVLGDMjGOxG3qWAcrsX3vrb0pj5bUjIicwDsfiCl5/glFNAGDvDwbhQ7o9Nq+WE
sHPgLilYVZP0KkCLk38giHQ/4YrSo6Cuhaf/SyfAsv7lCFYgAayolRHNawgXxKw2
TnwhscL+Un5mxx6rsJzU6kQALTsS9CEnc2COJ6sVF5eTKY6UTwulthP8To33FD8+
GEFK6HaHiXX3R3J7+LM+vMtWzU7UdOIWEkMYkT9UJxyRq8kuMTahVq6UgI73/k4R
2HKA9N6jp1FsiavfS9SR48YE1pAwOiYbJQum7uNvr67zLtvsPo9hRMn2m/qM23qX
1g0bK6fgj3yjltWDc0e/APdebhjoUnBaqVVE9L9UvahSSRQglPb+7uHxsNshsRH+
i7AupyXAVQfgCtgfBFdBHiHwSUaoORWzRjG6aAPDwPhPQBXL7W1vH2eLN/qWgP7s
GfTMeKPrP3hEOX9lAxoI+RejFT6nFuiyWN7BDvD1mMCfeoQE/+ddYJyzmHRkIP+X
NoXC6Nk76+j000viehslAWUcaPVRPnlJ5FfBqUPSr/1bZ6XVosRR5GufJemz4duJ
H2KsYSoDM5Orv4CiafyrMTNKU4VKq1UBIr9jIJF8dLstWqjaC/U9+xYR5ZVlXt28
YzXm0FNNlvso4qzm6tXqwhH87dCm+kB5dr9CdbpkdrBmXog9Gt3Bn2KjryuT9l8y
AGSCrPfY5q+LSpOTv8qrlq+7X/VJkd8Ttj3VHlKzbxmR+R+OGT0DdafHMoUX6Kjg
zx+Q56e/MEeb+9OMLbuXbdHc4keLlPcfQY50d/SJhuEMltxiS3ZVIk6vQJaYtWbI
MTYSJ7ZTf+2ZrWpHHOe+uqKy4gVKkvAY1fnXm/IQCAi+WjTrbq1BnkMIAzLoBmbS
YpoL7CZi9Cluy5P1roEKvPs2lSr0nyNfpFa8jFNVT/kF3ybBi9EFfYo8pWTJ05DN
DccDTUx3IHpfw+MWoGj2OnOlOcrLHj7hX+v0dt8B5L5PEYrgvSLGS/4PTdNtruS6
aBtq7g9MgWutYwF4/PsuzbmDJmqYlD5d0Mn+jvQl6A4=
`protect END_PROTECTED
