`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ep7xxLffRVc9rwT+p96mJnV6L9cNss1YqpjCRXOmMTuRPnL/IAWLQ5CY/bFsI7FU
dYf311dHEKmY5Knsbt/MctcsB8roFA3RJ2jnmlB3SHL0wDyCYyeVdIAi9TGasGgq
i078Hxjuc0VhM7YlMAjJ5EmaXmQgheD4EHlJQUcRdnSL2RwaeXtY6G5iXmgYhCqo
rmKKise0slEFfXF5sxHgAPvt6Q0+Gs3Mj8Zm9kMwCzrzhYxyO8Y0CE1z1peDSou7
bd0OSzfTjJLGRQKquaqbWtFvYQ5qEdHnKOT7yYxV20+fuDwhAxBDGyJjnnbsFXOy
/QFulSyP/ztiMrthwYUdyXiJK/dexRQqIKLHH+M7QVSJfoPcCQYyvGdzCkKRcIs8
smn5uXG6trVkyXs6CNqmRw1YEZA6faNDKvDn5vCD+lTSRzf3lT+yycraYOfsr/zE
6jp0JsGVHsvVkXy45y8mEIE04iycTio5eyVVuaCM2IZ4vWCx+idby2dGIIprt/W6
L56M29WZJQaXKmoD8UTb4LO/4X/6dKOhThgi8JoFb1IBBbdHOrWMm2TYiwfYTdNi
2Wta+4Bu97cbmtuzUfno1hqYrN1gT6uO1UXoJJIRifZ8PnI6wDftureDiEtXkIwE
BrgAW75kwIA6WNiBQKS4Ng==
`protect END_PROTECTED
