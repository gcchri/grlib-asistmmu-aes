`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3wvmUGx/0wDL4IHNvilnjkykmc08pIw7JUO4ITBDvyBzGX0J4EQz05rKiYcM6HAo
tMAdgXhbXURbnsXZfxOmT8DhfBKoRFBJ6++oXqqewhxBpJ86s6JLJZeXz51v+2w8
R8M6bQ1zXnSDw1d4TBmKKX9BOYDZjVVNRqMfkiYrjAvK7uDPh1IEY3uX+ufMP8GB
UaforooACARDsqwNnsV03Qu66QG63S1c7TGFuqFWwWrXgpRegA0W/8RhHSQBGen0
IacDSDBWUykhu1SukNjrCbKBQLYa6YZ7rp9+yTnGn4ichUwFvQzRxfGztueUGSV6
bBybhfwTuiYQ1kOLb9G/FINOFCU/2LFxNm02a9fdBrWQlij7uqgBFK0+S5hnOZUm
tXdXIfcynWKCGDTGlFpYm7jsuXRK0uKwqC84dOtBJUVswpKxWZBOIiNXD6vUPGW/
cQiMmWFrkaLpe4PTWP1Vft++aTSZ6KNFiMWmuM7R4Fc7QbRpsGCNYl/w/WzdOmhT
CZQfeVeaTRZ+GUcRTZszU7wzrf+ksPm+/mEgX8oZENExNcwo6plSe2Svs0q6OWru
emzSZVAYC4c+/FBUTo0RtpACFEUSxJjkH0WDFgH46MmN0ST/t3g9kCw9Emr0Aqc+
6KMqtpFOz7v1kipEiR83xADMTPlYqOkyhackUGFCXNN/w7h1WcD1xEqnmV5ynG21
NOVnYgYiucOwOGY07b9lSujhVDsrigervfEQrMF6LWGcPzywqvYy9wUyaK9sCfyC
jja/ZOi8mzA7omOVZ0PQ4xaVWzz8OK7E6J+ZQIb4VYNz1jnYGON8A87XeHzZw6tB
OUT7T9i5DxBn1BUv//h+4xZpfND5KXPxtsMtA028xH/Um+5eyjVioB0oRG1XTmBK
rVVKfSl645/pPOCIJvxeuqMw0Gjcfpt0qzF0ZiBiqSBFtEiYMcB/OBW+hNcYOxhZ
xGFoExPpTp0YcipSN0IQb7kGOMqJbBSbyZic5NJwpAbn6xD7iHdawCac6QuIakSV
4MPlA1U+pApDujcuzw/GIDpeQPhZXOZCnqc4Pz2AsHIMoNxp5O352nQnwz66vfVh
sYJPrS9qMj8fCiFVyFbf0CvdT3VN9HxN/gg9rC7JQALtxpODwveQ7cV+G1ct38p0
nko2V195oEVNQopuyOl2hy77wRuC2AXX2VoJ/0z0hHRL4wtDbOsNeKXoysKhkSJ0
1D+X7AeWM78SfOF8gpNbh0GOhYVMP5tbD4eYU3aOjamwctPmJuRbHo7XRPM8QD9w
bCLeX0Enu06jdqasDq8XuJEXcvszxke7ifmmHAPaCDnwHoN0iI3XEeDO5jvr387C
xQZ/Sw5fUErWYRLOFcd+vKU20IKLLA6QP+eRIKwK7e32lcyzMHQGBI6XDuqjRmhF
1b4SXfoK90y6s0D4iNpW0wUWmNlINfHnkCMgsQthiB+X6291meZEP6RgWj+6l8nn
DaR5gzCDl0hDJcR7an6n2o08KTeczW1l+u+1oPq6rM8Axq1z1Q8U7cA1/S7P8rhw
5beJ+z22hH7pIVqo2D9wXa2JNggFaTmwrFIFenUg2aWTLnceC84lwMyCqtcrd5j7
hCL4Ll18e7VK1uotTzrcDba/63/amEYXZNDy8bLc0aNniz5UkDHr2K2eT2+JVw38
cCIr4SnowktEH+fQzCbDYcagIGW68pFNxdGHzoHASvPTivA4N0M6PvsRR+VkOjw9
yGz/w2xp77q3kKURQ9RLGT8U2L91d4SO/CbJ08oeNnujkXnBfOUtERDbk6l0MKJD
VfiklW4734uGK8dybWnDKlsJUMccDgF5Jl1Yf1VEhsdlixhKyCJweb/khA7WT35T
U8Ql7F8a41MkeKamgIVdlM73YBHa6N52JBKHKORbgNFxP7BjVA9YE0dlQWomrcgM
vQvFJPmVqQ9oW48rNcwHiLmiNaqwps/JWT8jJXwLLp7SEgqIG8S2LtM7fGI+2olh
RCwiBfjHQf4uKlaIkAjCcHuACkX13Vy63hsxylJ0RXUh7nLQIqVsN3Ut5+oBcUwr
WkBQJiCpnzR4z0g8drEWbIxKtI6njbjprCtSWyxw7tn0edMnpYfPt0Ryi8Y4heBC
e+xAPVKKptLHJnZXhpOMNlhYcs6AbRV6lHvgc/iHINP6QEl9EvjI5O/0zwuv+30V
eRzIcNOpezherzXjER2Ea3bvariyCEdE3ZZSTKDRSPnecL1uRDnddRSvTBuHiqgC
Rb1jlIZnl4e5ooUob29hO4kbNJW5uTRpPrpLMnD2tg1cgI4P/Q2KkIE19+1/PlwR
lvpu4TZcQYadvVWCLjDf3iNdfR5R2W39KIA+e0r9HarRla8ewzufVqTWGJs3frZq
pQc3lGPr8v4qGEy1huL9EnqhUYMUO6WmlOO4csHsl5hqacGSABdk1TRKeUIBdko4
+uiX08scKms5e/v9I8JCNVTghDkCNgDQjodOtbX5N7i7wGkSjKmbwgkiYJOmrTG5
iih0FBAIAIblTpiMGHu8z/vO0RkBB3axC20fAEXH8YK3Z6gTD7qFoUtdQtEk9EZm
CZLZqxKL2fSz1tl+AAcqW9QhTsi6t4gmWmSpBozFqXsKA57OyopOwMqIlTXzmb+a
w9h7Z4UpLp64TazxJaTNShZT7CDb3nwtdSvPvTC94Mr5+AiwgvFqhPUJapeEnPKK
n/AGlcQhmeSoNIh6Noh+0KUE2wmo/oge7PloiT49RYhs9sD+n6u114ZpDV18WJPs
Bl59WI4sAGIkc6l9NayXpO1KAmARGMuGedkQhENickPnHmfekzOdu/heTBD9El7R
VEngEqW24fSqBQ/m5kzGFQ3bKHrX6Q/QvKUkW/mGa/jo1CzRucehRSQ3BmS3+rYt
f3ZvEnkKv/+2UMSL3oPn10UYnRqPzVH1DQHgANMJfjAzDiqQ4zJHrXezVldI39GJ
1jU6r/Z4NOZZqmqdtxGCG881C0WYEn1uu27zENPj17uoM8hnAyl9mzLxFV+Rh+Td
/lY6luzXhxgPK2bzoi8hiNNiak4f0yhxjFjPeeWSnxqcIOADrKm20z9CzjwLD1UF
3iIN53hhOsM0yP8e78tK9ila7FqThGqx1FUyZIv3HvZfW8Sb4RGIyOPbmBWv77Xs
f23UXfs6ZBe8IuJr+AGE2coeUpMpYcKg6EPgph1IYk6ISmSi/spr9NnHpa7pqKly
emQAiZi4FiUHrA49Ppme4EbIqTBEXrISWKFZK8NEFmPHj+zqcYZo/h1jcDj0AX2g
xJj6uRZzG71G6Y4nYYx3J1Z06iytlkAl8h7Ju2rK5kvTexaT/cEraujpg394j4VE
03/UnFEGEEN6h5sqHrnxQHM1We1dWVu0YvQ8gAV5pfdV8QDqZoGcoU1fpaB9rL8w
lAmZzR385oRk3ZYarndmUMSosi2w3lRNZFzk+jJJEwSavUNIyA5CpDgEezOQ7S2S
BAFZyHUw1G1+7gJXEdhPrYYfgzLFkYqbmAw6GWpgSbZXYJ6pnhvymCHVskRpKej3
cEbT6OR2n7sXJ+gMLbgMTvziV1nF8ZTHTn+XCBSchLbl/BuV1nQTbxmV31V4Gls0
oFHYWVIIQTSm/GqP906Ca15JZ8tjizj92c7jJC4O8ntazVcjLq4FrUHcE5Dg/CCz
RXT2eg8HO/qBuejksPC/vyJkq01lNyfLfX5x/levllsa361Ama3w+kZ4E9Hy83aT
n0oRZuZtD3Td3cIdfTJE0j1qBc5ZE5s9fAn+yCyrEOgySZW6YULh5NP0zccwRMjM
/CCKKwE09nuhk2EpdaA3YgPkZQQJi1WbyBgzGmTh2jsTNYJpGJT2dkZMC9L10Y8S
SgW/hRbbByDmjSkzpAAvmK2Kxvq6AV6Ivrs4VIq/o6SulgXFqWKYGK60VC+LUowd
cyUTE4pe9ZgGaz12Wr7jIGjP/r/CMngqEW2WVsxSepyVcE4eNSvRZluxaw0tSnQL
v/R+HGCu4qf12Ke4xXlhY7FlJstUmXi9Ho3gFU7l5o0Mme6JL6XZPDH+nkOMhu6s
Rmd2APGPSPvz9NJrPRb8VCxNcJzusRd/5IShhKWqKg8k88aNNuPAe2zh+9f+vFPV
2xRFZ/Ix9mNePQX8cznZlQiMZw5Nihf/g0TsBQrjYYJeo1935NJXmw+ZgqPNxyBv
l4xplnMpX7WxHS5uQH/DkWWNqx/1EgjWzv8+nujsHp0a5vGKezJqIz5hXXfbODcg
iJf+L2owUoCojTZW259P7eyTtSqnKZDcztEvOEIAAeBRIwdbAvHI+ruJ0G29AlqA
ds/bkmqMgh1piUhGEtJrOF8/IRgLYiiHYZrlLqvNz6YJDAYDDDLH4LHu0u25fSwe
a89VjetlPNskkAuhhkghFfAZJ2+VAhL35WIBMBpXhGrSvtx6sC1sAk/U6jdT29bU
O08E9Ym5Z2k6En4MI+lpq0QRQKsq0Ftc8jZMEGw8TM8T4Gu1mccujqrDlElQ3Zgx
4x3KL6E545ouyfWouFUqtfSIBaAvR2XpIBZvfN1mIJp/b6IQ/tlF5vayrQWypqUN
jGgZn75xCLFI9zQTpEftMRxPwUi74l/zlifyAAiG0iJqeuEBiCp06aZtteCNxHAO
GuEM84earxQBLBW9mh7bynuR2cur34tmViHj4ZbB9EdUeZN1NHG+s7Ggzd7TEbxb
Y6wCR0iMilxievqQIhp8Y3s9J07q2F4RNE0O33//TOatvmSYzNCvByP0DfZVAYuY
5f05RdLGlVnMPqBeNQd/omtoRRlfg+FP2tiD3HhLU1snjvlIZ0wdOVRy01wRqeJK
bqeA55PUe3NC59XCB5WbTj5kMU/El4oZ9cR0cFNmD7eCSMFS7JxhuHQ6WiUeSa4T
5p4yowe5i5oyxNBXO3nXI2FaSv/nd6M6xHP3EPkbuBbNkRqq3LUad0QBlmG+H5aP
Bl3mQixkYgm75+dKXllYstCfGTEqq3oVWVff2Fgq5XY9t0SZLEbJAKwDM8FETivx
IiKuust5z0cc8aGX7Vw4vKPHrqpyO6oMljDWrjKQortwUMzypoQUE5zZ17/P3XwB
PkhLN09vfG7gqo/TbNaZUtCnBzOxWXuVRWnMM/ifhV/XsHd7/GtAfuTGUkGf8zun
e25ldXOEeWcHc3FCVCq1T6CZNf9ijvsbtRrktTgojidikrLMl7o+/fQ+AuKL5+4d
XMeDSN6cHHkVeaAG0pF8MijftdLmgbWQBbgiCEL7iB08F9gmhz6PC/pg70afQJx7
OnnmERQcGRfipcpeBzKxVXX1/5EUCRzIERGDtGJ2GXSlkF6WRMDR8hUZswpibVXa
nEuqyos/WZQ7AVCIYK0kk1hIIBSnoS+BOfztNNa7W48Wmc4rcEs5op8+h6d7xvO5
Zb14NggxwxYvb+vqS9Z/8jXqACCKYOxujBEGaPu0HIRXbd8BKTrgRzPXZdXO5B/O
OX99fjeyISUpGUkum32LTCTqOge9VXIn5m2HwRNAb1ZkQLzQKfs7Iagy6gQ+GVxm
AaS/YA3jtNXmYu9ECKATIHnC3jeiufD/cZIAZQKowevgFw55jd+JffvFUCCGgUxp
IqCZGwx1h4yO0hTiSSLAh3SUhLxnmid8yMXhWUlnP+zJY+KUGq79DvmLgt3ok5yG
bBxTg0kIP26JlRpLQk+Vjncd0CD0ZINMgXsgYCnoEG8LMc+RpU26ZN1+lfXLeH/7
ru9N2ACMMrgOwsjJGJzVRja4gkhZA/jERSY731OhVxu7If7V//L+GeJbGAnJPpRo
OMWnltAwpXi7YkR02kTUVWPRBw9IIgKXyJweUvhqLwwhIvfuH5prypFSbMtCCkmi
xB3g7rA88EcNto9CRfcDd5FdFmiV60vuLbxWIZypDB2Yb3CmZFoodu5CHjsk0UAX
4Pr2TSs9jn9YcizSAWgsYtyc33JLjWLlvdqsasKrD54C0CSKTGkIdOHjjOW4hGVa
b7NOYkAK0e2fDhRnWzfA8zUjDKLAHro833Yj2y/d74pbAd4B9acokh4owfdw0cPb
8eUW7ZM3ubXnHOSLUVl560c7dq4KJompo0iWO+UjSznDVmdMh7VAQNNpZlkmLqG8
Kv5VQgHNBi2uNNcGdmrnr3g6aeTqCE4dYtp61IecgwX2MU6q7GqK4k2uSylqtmMp
jaViiRC8YjPJUG9wIP3HP91JEH74MgOOGm1FfZfOmRWSzoLab+5QUg0P1vDO6H3P
+dSn3VBx9rjwoGSDa5gN+h8su5Lw2NMfpRk6r7Oc8uX04SzIsYvZnmxoMhW/EKBn
gsTjyIC2x0wA9hTuW6nFRpwc1AAKYCvab8NhiAzWrYVyR1aqu0GnBGTD+9MO5zE+
GHwMQb8mNcNj1Geb7qVd0UidhUeKhK0LrcQ0ni6dvm4NFX9J98t4dE2IycIN/hB5
hF7C+E8kprXQ+jEAx/WP05ISh1Yer/6+ezxH90jQXj2YWOAmytydZOQrmriaTQuP
2r7X9kskHVWO/doAGnyFZI2DoyGJzeShQXr5y5v9gt1tHzzFoMIW/5UQgazxcBHw
VjRDv/AJHDt49E+5RYcTDHP1zvFoYNHr/zompWWuRhBoJ2tbqJGp9w7+PJ0RDmHP
a1xRBBTTLhJI0MEew+SbKB1dcUP0SPWWZTDzN4kPHjNxEZstZMOOhDMZ0r5WbCwA
bU7MFiOgP9H68RJ31YBr8eVu7bU0+h3AntmmAAOpv1ETnsRLNJGZgUBUKaTAFqaC
OQIjNkuTay672HSa9S9lAgY4OgXfU0S57OKOYfAyBb/ITm0nHAGtbWU0ZEde2j4S
/+2jNYvTCJ/sHSrgtzdXJ7fKaOsuitPFg2Puy7eUOtTJGWy3GOeGTk/+UZIlwKKB
tJ9fWf5n6W/VW4na2zgKjPDXClE987oZtLZgibUujjAAGFYlL5Z2f74d401axOYy
6yBASdQzdvceUS+VE90MUd9vKJr7B7A3uxjPY+EHGbDHfIGChQoAWw8XZipxj91Y
3PjbnTYOZvPd1DlCxCR54r/8hk2OEaBAnkT1vvIWC7P/k6W8VYwNBMPdgkXGKZHK
IP01qEQ7J9OhfMILrQZn68ty26qcHN2YfB0PeZIkn61GiUdyLZfRGKOe+3gsLwp5
GU6m/qLJe5oii845udoo5TFMkR9fAm8AVTspj8SyCCZ4lgCdbO9FFQWCe/msvHHT
wIvmctH1rr/Id0kR/WO9LzFUWznZKb+/ZZX2rM43CZHt+nluBw6A6/0Bd7NpNIhz
V++MqlUU73wZkRGHBN3BOVHY7zu9vhB9uSU+M+TcMzsMklT+Ad1OAbn6LIVvjTJI
tRsSukJhlk1VKMkxBCxlu3b4NIOuuLl0MuUFAwXB7UptEfpOne85M3R1a3A8qULT
ChyFapYSw7dv0/Ne7YFT/l2nwqLG0H7rmm1Q7M1OtTwcD3pRJMY8Ola1tVyNKdhg
9AK+tJpHMljpPARHBOMzagspfjEhhkEB704dQc+tQSxU7A0MkQhheGUyscMIc+t6
ZJfmPysFSsRM+m6TsaCpoPATsBTEAK6yhDInNsTDZD1b1yujHehreEO1cSR8xTu/
DQGXuFuT+G+V0ZIGUvPB2HSbDfX8pdGVj62Hh4hzG5WwdVFMN62DL5FreTAVk7QD
dqV7S2o9nEMlbAx41zBv/PT2HsVVUJ+HM5iI5eF0EywMzJS9eyDi62QwAXxu/DVK
7T44jO6GfFdepJqfMH2wp/OyNs/Xhd3nwozI6FMBRvrw93kyiYu+K8UtkyZVzIro
RXbO0h87rD84feImVPLeNx9F/GaA5HA6KhXPK70Ih8teUQJoUgCztkBSfgPClHuE
N6V5ok4rmQ0TflB246+QInoUMYQLgLQ9k++PUGeagST8jTeqU9OwrQn3K03sM1pI
wV9iBM4x8KSrba+3qLZmYEYoXOCQPQ22In2KS/xbwYv4LYXb8G39AnOeBy+rY+nE
0763iGYz30N6kQWrFzOTrQovZzhEWf96tybb35tIKv7LSZ3l6qDvgXiWiku9104h
bhr8szHIpZkZEVSdc4JcY/RzjYDCEjZJ91KCA6j+ynQQpcC5KxE1p5kn+jr7jEOB
rdV2W0WJ9lJwd8dpQQblqHpnwFxmzXIK35BPmLWL4TQzN2amh0o0L5qMHLv5LgXM
qcbUvAEi3/02Uqo9Oesh0K1F4na0F9TgdQlCF9oq7Ygg4Erle6BIqYPFYzq2jMw7
epIIfV0uhp0btc0DvHhUACDSuVlElvIDPO19IuL+0uNc4sJRvEbxb7yEY7aXyEk9
13+YpQl2sJbtP5B8SzDevrZptOD0jmq6b7ImcNU29g+nkFxVOG3wZs4F1ZcgnO/d
9ODGCIbSPtEO2Bed3G6JuRpyxgHETFL4NnISmIB7Pxlo1lbSVFmUKT1Z4Rplnxht
Mdxac0BuvsCc1yJX7g93ZqdL9HemznfA8V0uTto3DjmYRB2Ok6n89/oWYuhqZxA3
pOuA49xSXfxzJ4iJMoydWzKKJRr4zs7qOoksfox2e3yiRTaHIovviPgbGOcZI8xA
9miEvoybUy8xRWGNuz3L24O3cYjnvt75s4NF56K2YDiiy2+tAEcky35u1N+XZEmm
Kfg95RmkQhBMddrHnZ5i2uuCq5fJ+2kxJ83/08+uNEY2R6dy6MWyQ/1agpGBmWEL
71adTQ9msd7M43w4U2uXYjubnj9zRUxuZohvxBxZfoV7oer0GL3a+I58llerB3/G
eSzbvMZSqzRkjUwVvTt/OPIoU8AMq0cjoiPUvqNT4i/9a9puSZgIxqd3l8881Vsw
yFIreeUudOz6DM9oh/4cPOdOR6xcImq/WpKfOULFYYB4iqkpQ1anvvcS5+xo4qXs
PKu7plIdhp/c1LrFaJLyFSrwYw+VG7RmwUDe0FrFwIOLOzu2MEmV+naIz5zwDzLD
iSstjDASohKELOJA0Cyq3NFWaUUetAbH3pEdh7yLqCVRDKZrCYiAV0gbRsRLofil
x7RATBc6azY5Q4+m+A4tOWEq0bItwG8Xw1jYxwztvbytLhY21YuCbfUsjdPLnCmX
pY47W1opX3PaTLbmKev6I7VmgiWjL8r9OVm26u9bJ6O3REvVW1ONqdsDfZ0aOPzZ
Dp1yv1oCFpw/WG8/7673mJX0Oag4uG1efx6dm228cwkGfaDG1eGJfDYwUUhDoOYR
azhMFiAE9y9WBF0N6MbzAsRHJM87MHrkYKuA6iUOXP7tGrEhPkGHJkHnOhcdMHmN
6p4bvxYq4thX0cHwuxKE4LSjO0WmAEDl61gILFqbvll0yp9RptintU2Q6ns85hWP
xxTL1BEb3OqcXmXWMcmdQLTFCieJG/Ule9s6U77BCfZNM/V+9+IzLPYQPo1abn9w
VS9DFDlragFeNbcAdzIxqBqcJPpQg9lIXOb2w9nMbgvBiqc/gBDcT5+Bx5yhyBT8
l02j2PXXmBrv3Q5f/SAu9YZEeslq8X9ZHVlNXAQHuo/RbtaGo9rAmpktpvWfvj6+
8LNUOfpEvmAIcO+6yJTl9MnoKU9gDyru8KYgXUoiM3+aoP4T3vo44D81g9X6ESh9
IcWZUYYlshVqDVR4g6+Hig1Eeuct5snKVQ4NFGv5ELZ+1B8C9EPxPwWXpEB2+rsM
+HioMJbSWXiG6eKP6p3JTRtJmi1A2bmWJXFG0r/QAXjJOGRJr7teXJyq913r1qEk
daAjbt9wZMxbl1wOQzJK3/dm+Jgb0nJTQou6Ykn8sFxATmyIy51C+FyfaturrJMd
oENYtggJiJ8uvnVXWevyFmiB1wFB0Sjw4KI8GWCFXLpNA+deBRAzQyY7nlCjG/+M
v4eeu036Eh5W3XNas+8IFMBsX/iZiQOiTXf+dnWCzaHaCXuestiftQcDpDHMjklM
65msIznR9XExyXEo22wf8KrJsfIpvj4SvNsjmgV7GkX1NRTL39axfjK3wqFHDto3
7ZC3mszlbX7nxtW+pSOWfLKh1NaNbEbRybbbKW0Si3G+ykPfsykLSlVPmKrYoHyh
5m8gQ/WV18zEJXTjzvodb6BSUfaxOzpX+dD9cYhNjfQS1/GwBb6Jk5/lgmPpzsNV
MbJ7lLKmFOXCyD9xWuKaHZElvjAdTio1d3bG76Ew78+/gLIj4Kg+Zjv3MdAud57m
wTn0HsEXOmLMBY/th60mrjqk3vcVFKaKHFuWOSVqd1m1h18TGAbo72V+fi5aLO+W
c1vhimwZyrw4P6HAyimKN1DEkNHSLtsf0D3/oGK5GZ46NRy5jNPyscM0L9Woq0i+
0ZXZLm2jpyyMvZ/FQgf0Z3u5cO3wpNtn28cykqYjy2EQ/mFeHhGrEq+NiYhdqdAr
6+mdfjUE/h+J3/etbKK8zd6FPByVb7GFIgwd+Q0k6rZAzvCp9wTF209Mr0yimO2k
ap8gxrsf7DmFEHlIoV/Coeb2CzNqDhm1u8wKpGxLeeHXIAzbaGdWFmw79rC43yOW
Av4CpbpwZ8uCII9fo+hXRZb1BIAN1XRjvXqXKFrXsSkgsjHKn2CHNNnMekrTXdHk
oiNmKjA79RabK00SncT02D7x6cg5R1Dr7MtAT2nZwtdX1L5pwqrvDc0sQEPMXOLB
68FbPrFDvbK+oQfykLHYO6FU1JwVbxSKZyDWmYOcGkgoK9SI1iFfRZ9YvLurobP2
oEqEmlcZHOj+G6SC2j52KzcTALHlRVU7ozj9jOA0b/ghJ9s3POVPQE1qr4Ss+GKK
Qc4tPT0AAH6mq4Tv+tvrM+wS8PNhLX/7+EfoElTiLXTkG6RcO4aivMZUTCJNvawk
AWSI7iOamBqI/uEtYrYSe/47n9smFW8XMBltDispthWr+2/NZWEMSLEmeE/s7IXa
cbWzzfGB+riYA9poYYwzDogtAu9+aAdI8y24P05dCxqbAlYwqmVOTnW7Ya/PEV0p
D5boW+5dNAom/hOorRLZgwfVH+2VfbHE8y71Z0a4CIKgbF1w06Lmow1AKkqDJPV2
2RhuJd1Fipt3ih7NWu8BSYp0LhztEtFYkUfY+M16/JsGk6UV+EaZvBoXJ57Y1qkw
+bz64pfJ+poetY7a363tDtJruiL9w3hbDrGxtqYb7++mVsYHOje+MV4p/OsxcMHv
OF0hxl9qS0rE9fh7FKv/FdA+OH+YD7Cwzq6IHO4Bx378/gx2ZPs1Lzkyp/yGzIwD
tuCa6EsdrIU0KmQeoQc9DsK9jSulOtz7sMSUfT7Ov1pAU2TYST9Ggak7qGqZQSwO
/QZGoCHyUvA7yD2/g7daH/PLTJcnIplpCvuDFRIscc4mZWi2ZDBAs4817VZDZ2VU
U5Z8jdf7k31I87tYbfw0i3YFU9qkEM7hpZxs3zoRkUSeCuoqQYJgdDcgzeVqbSTJ
lRJDjEywBpPFpstsdpOcXm5jT0KXcGXSLhMytGBZH3W88eSGOuxnMXD4EUdX4dfL
vNfXw4J0a/ljl78TgcjSTfsEWvdn56uBYG4wpttuDp6Y9S0edomdss5El284HGBf
lA7IgCPBjXI5OufiM3uL03rrOt+0XGI3Oi0RPoMzU0n1Ad9NgD2UNdghTGrK+wOp
2q6p2fOgVexjYxk52rMCSbGs+Ek8LrfwFcdZ6PB9znxyCvFgIBq3ZAQPR4vEIHw/
8lCJtARa6O3t/Gqvfzj8HFXAqMDoPGbGr1oea+5MWuHRZ7BN4tz1vs7W9K//ZB3V
m2vQZrw9Hu5v72TMMVkDD4d+0DM6L8vz7sK8z/9qHou6UZkrYqL2pWLaA54OUiv5
4wHpOcyJKOxGjzcmqo4JcIu2LpgFSqPnJvJeN+yZK8vh6YUfzNlaYxzAoUigS7dL
gRnq9o0JhkrM3HBSqBf+Llgv6KUhI62FIJ+f2YkkjRJmgUg2BFrPVN0SBYJ3fgSW
wsBYNzyEcUE2J98AecIx7oZDkReftgzpr3fSd+chro0aTIsmk1we24lBOaC1Ircq
OHLcuQPOJzRSA1QalnNfbuEmFN1Mce8kqZJHAL9oMoX7Qgy8bL10UlrXKPeM9PVQ
P8AJXlTjj6T3xPCZ8HYMNObKdWNnfwSSLVkDXz3iD8vhEaNbABrLbC0EzTuFkpHl
MEpYnDt78HBOfiQ79p4Uc2tEh/hTreje1RKrbtItRzZMLZXbxJMJiXBVIcq/ED6X
4CF6Kb81pq6tEle2H0Dgxc+0qSLt7xzR43ZNHtniBKYSpVNJSGMp76MlfqBBCGFv
24JAfzoIj2G/mW5UkxRX8Nq7rwwnRcp5D2EciV9GBWIErdcfIuPiKe6vHGFd4Loj
ILIPSMVISKjAKXCysBI2/RduhGN319DOVrQgcnxcXe9Qnl88SWNW7y3sOi6cGnv5
fqxuAPS7TPGcoCDAcY4mAk9njOgN7WsCk3LC6ErL3r/DQbep72NxLqzqJtK36YAy
rM717igGTtDruwATJ9Kj95xdyIFHX7Jlqn0KH8aep0NsD44RpjVHg2zoL4LCiLu/
TUtzI+BTJhjjCd+EyuOMjWNk8XFZhMz8gbSA/Hzn8oPJ/eLbytNrvuTb3Wz0qlno
DAeRrEGhpocBTppDjQ9za3XglohjRY9r7cSr+m+ludEMSmbry6LpU1aVJL4+o6A5
8j8SbG7eGOoc9zh8GZEsPiUCgaq3RQBy1aMcUKk+KkcamFXbWlagjwAjTVNqYrkw
05EEo/qCn1gnyb5KDU5+tikyfO59gEfO7T7Jgd3FJzwpTkdTv2hm0meFCSJ690I0
kCk96BiyCW3ce1u4QF965rMhHZqC9MSwhxjb5iDv3WLJDxOEFcWjYwFp6cO5+Ayx
VdJQbffYXK88Uhma80yjCEhP6b5lOpdPlKBS83+W0N/w9s2ly1V46Y0NaZ4PCv4c
XScUg5KEl04a3gMn2Q3cop8rYhhC+OfWhAtG1yFxXf1ocoYO8kif6+0JV7vKAcX4
1WmDfsBApply/ntlLMuA9OAUkHXdxAtv/+gXuVlYBp7izxUO/hh15TXppnJoS+9R
dIJp6V9ED5jVJS1S1UOrqyTg9vB2WvJTAoFI7e9eJ0xEoXE5EG8H9/ZQgi+vlkpz
ppsct6XuUYJG8Eyeu2epn0z94dXrrcPqQzki+Sp9TSQxLT8UdO3yljvl4jMH2Ara
iOgk2VeCCkbdT8egSI6Xc4sFeoYqfmrVGuyEA47Ev8IZBkAAf05oMy9CUM0Y0wB+
lkYZarzhj3zteySqyZypB1ZKUGzNbhZsN1mID3DdBzvwiJsv+5KQZzJ1vzjBxS1I
ld2hf9wKTgo1WUF6tZ57YdQmpBBoWEV+Vjtqvn+so4Lc2JfGzAyensClfhftIjav
SlQxjKzrabdJrXFAk1ckp8Vyulo5dh78zpysCbcMEvAYwQtoEZq1SXoZXY7CUwWz
2bMqY0gasIEMQzkF93F4WwlOCfyx4NCnFpWJ7dK9wWKeMjKyYJFNS/rfay3KqFX2
uj07lDqlKK90gb+b57HTxAhr1vNywtQRlzJdmtLvxu6Dz1tTjIHgIquTaqftGz5s
pwS4VEQ6oCZp+lhqoOES73i/JEGz1l+sakrf7lyqS5hiDREOUiSnBXoZnbiw4yLg
`protect END_PROTECTED
