`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f0Oh/kRIT7jtamwsY091e1kkRI/+UNayAbLXJe03MwsbzxIJ5rahiQBT5PjYnmeO
cd35wdRCUuZ6Q14b74rHwSISKGU8eEBqMpjdAdGwWXnrnQsrXaCfrDEj2b1ByGRi
g9t6h+lJU2prKrH4xdPvvK02GgbRlXpQ3Ee15ROjf1gNOGMoWKA7P9df6iPfI9nn
j0mU1B1Vlfkef9WtRMk4SBMkTZo2+4eFK/SxqprPDsQCqB91BVYduQ6KHRIJZ+SO
HHD4jNg/of5IHNSAWyoX/0Hikh3RLux8AdmhePI9yRtFkS1lX5Yhfe4O0dTONBQ9
BEK5mkkfpb6GLJXdSK86R0osCeEMf1fcQoreuKV39aSY/O+IzWsi2hY58/iBr32W
o5lf5cyj+sByGOSh/sHJlUD9ObL2VxDtiiLalaWgyyPAzBhyBPVCJDlm89IVx7C1
NEG+e/oYI3tfJNasZgeAQZ7ejoK7JayW0kynC6DBVY65W2FVMj5c6o9ki9MhdNVe
RW1gSfCMEWXbf1wtY8C4Prjo1wTeI+oZLCl3EPnmoJ6i7/SDrmJ4W+sgJ2dlphqN
vMiRUNrQeEaD7xULX+AoJGrvq76A1MLCNVxz+d+YfeXhwQVem4CyDnsUCwfo5UKi
Ov3sh+XUQCAlTr8ZX4O8fA==
`protect END_PROTECTED
