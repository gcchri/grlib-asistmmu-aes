`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bc7KwgS1gj+SQYoJ+SKbhWxYAhvqxg6uU9OFkDRn6GYqrb6LPmXtD2HLgDZO6ejJ
6vVloN9he47+ekTbuMzp9HjubpiKHME3qpcHHHhsxA2832B5ncISXxeynkP07zMR
OIqV9BinF8k+n1wA5U0u82gz1xLhg4AaJyolhPJn8x3WP4rSCLpmSfOeuv11bBv6
djfHFiw8z8ARggnWxc+mim5t/spR4dY12jgO+rh4kP0MLzaMJV39hVG7XxWFPWKS
I3lzznBA1Kip+g6jA1xr0Fb1hk+gl51xiQvMLyA55YFjA5To28VRMt5zcRq59qYx
KG7VN2tW0doPyb4whj3VNy+q422mn9RMsr2DzIsmQas=
`protect END_PROTECTED
