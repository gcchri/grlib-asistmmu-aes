`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJQljaQX1FpuI9HviXzPvra/BfPGTjzyzydEvBqs8ludC1DmSrsXbPkSniP1ITQz
uFy6EkKJOEvoeq2aWMVovyWTrLHdrsYdfH53KDLWWtBNW/oJAiwN/E81nUuHsKBg
N9svHb32j8MHtcqANqXwcpKGCKo1pZ/CBFaAODQQv7Vmomgz1S5wColPILnu8jVN
eH/ZBtwawy1zo8uu9A9TaJ5w588nateZi4OaigXws5Ba7S8SfrKtAcUzD7epOWtX
GG2mEmiydpNeblInhSB/8g==
`protect END_PROTECTED
