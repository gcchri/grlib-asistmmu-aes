`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2SXPqRIGGNRX4A9uHYlgAQEbbJqaFrugYlv06QFQn2yKHge09gxXEznddmxrfFLC
2ie05YNMcl6MUxPVExEahqRHTsvxESH1oBNHVEVitlWITT+JbOPH7+5v2lQI4dTZ
PCM99oR77nxYm8jYUHcTtenIbyip/If1JC7FOmRWbQrrtsdtKpEbnrENbSz8o3x8
+d7FH3KeKr1/4uiHttIK0sUKV+F7F12H//v//1wu+iNxCUQwD+lIImZJNkXN9P0D
8vPHc5v4zU2TJQjOleM3IsAz/b2QR1g7Txij/NA50ZBFFs9+kxEeb9OQvTYcwZcJ
MosueKcHYt4IYPSrqGzhip8zO0IvUddyYXnqSLCKZ3PgUrXmC+VI2JoMZwwuNgm3
durZpc9TXR1RbKbrHHBziVlVqaRflkylhnAfKw6MGcx8p1E9LexSdEvx9ncXCpA+
FjDBp1sKoFcwL+9pvMT+KMdFBhHBP+BW0joN35PEWMvjn43HHKhIVJU7oSInv8WV
`protect END_PROTECTED
