`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRmlqYDpKgtIzYnzUWoCxTpVfK3w7+MVALdyCU5FdxOC6vzIMyq0fv4BhkQP1KVl
oIWxclWsaUREiqD7qNwAHGKCV89cM0j76ZbRxxJHFi0aN4nxPOM2uglO5rHrmYAT
nQmT+d3UkWNNLidTjHwwTxNGnr5okqmXwTEA1psV/BUQ3nly/bJHJy5VLPU9C8Qq
pEF1QpiHJ6gz2sjNLK/MkKxTxDqRwIqGdzOq/ApyMG5qFW0hdgGo++CyZMcczMUy
dqJBPO/u6O1Xc5LUlPhjs7YKlaM6B/dtWqt0up3nMGVSnJ6QXTRQVMxqTvQ6dgcZ
dRYvSiNCYdxUMSxRxYAcu3k+ozG1UscV90WmHZ9NhuE2Vghwn1+OjMMw29bwQws5
OU7b3eeuAqRk9/uiveJMyUfY6MLs5y9GoEDeFQoTtM4=
`protect END_PROTECTED
