`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1OcHSlfu8al+l7bF7pmbJQnFVC4QTA2B0ZKGUk+Mw2pvngMRNxOQ5NhKDqDStUT
vTaCtB2AEL4thCkZ/4StC6gFrElxpkn0+ooVJpTubWrWqpGd2eYZ1g5freflU6eC
GM38QC25QIZAs+35Nt09KNfj6ZVM+7LZhefyHCPQQUJ5lAlg2JIR2VtuFXfpEIus
wn4uqLejGQVe/3HDOlSdzCcCaxWLZdge7FS0mS9LmXY5I2D/Q4XwVPB3IbxLo5ZG
vuZdbUdN/U/13QXYs3LYy/Ua3s+4BvBohZy2AOdwhawxw3uRch5EXllBbQihKEDc
MTnU24ZNdFO6W21CwfCdSX2RPwYv17vhspx/olhOQTFlwXdjrKv8QpTpDsTvAQUT
Fzp1vRvA2NO+jcuMArrurltRJ1CzGJad2+flDbrgxdvDOzycpA23Sc6A35oOV/4i
`protect END_PROTECTED
