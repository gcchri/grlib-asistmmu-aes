`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/5bwFDXBC53DlT5Enwsa8Y6GsRKe26RuHAPhPj/j+B/veDsPBGASINDI6PUN//6C
o116v3ynxdfsUlwZz36gcGWHV4NdNLXFs8H1n4Nd2/puh0bpusztpUJKVupXE5uM
2upDK7Qo9YMqcDPLV/O3bwjKIREeXfbJth26PzC4o1ocegIJCBRNDtjFcfJsCIly
f12yw+DZsxZbrSefTKCuVzwXNDosHJ+O7iKmqHR+oWQLsswiCYvs9AIbIezDy6/s
ghpkDCRo2B8vXOrN89oyTVBdRx5KQuO5SoCDuKsNOOChpkZ5vSw33eHuMNIVMsq5
CckYonqHZojEcim8YozAxWi/1BbzjughcHRSwW3TVZyU4DLZzIM6ddEk7Ghn7zWQ
MacQowepayaIoxBQ3Tuin4p9HbFMmbJoq7EY7WfE3huqQWtn0cSB2YilMLc/9+zX
K+Q5RixaIKfqBAlIiy8hP4l/228O0uF+SVgcc8MTunklkNMnYD46kO5Ip1swyFiW
iMctsevmsxc4e6wvxg/gE7b1yWfAvSaE7HCVmQCkG0woHRyIpFd+Uhf0ww2uUxmV
x4gxDpb7t5iKuiAkL9AOJt/Lvu/ecCW+zgUEXFSPZVii/rPDl23puZe84YucAEb4
wvAg8PLA/DzPu/kCjtcUei5Ae5u+863c6n2YorfvELBzEVsRM5Esuebq1FoNRvQY
CkxNZJnVhzUIH1XKKVAimFNHW3tg7tlCC95VZRcL8NdfB+bRlknPL0g6WZDx4mWM
jDRWdcufczkOheI/aUhl/S8ihLGjBCQFlRGAkhHxMKpcrXpfsWy31oLuKP6laG/V
Gd9tkxw48/ekFN+zjvrACzMxnURl1ZuAjUB6hMsXv182SO9sAKIFBo9LaTDmuaHS
z9sQ8p6+HW6zXrYMG1mAUKmYJ3ycA4pJTkSXXfldIgTFaPCP4eRhB5kD2d3k4Wni
fV79QvK40vc1OqrdlNeiWkiVG1Tu120pNizP9z2vIWg0pvW0OwmtQU0ZWi7ZdVSC
Ci4i7NHuG2H12GxA4zz6hAoWFuMqT0kAc/wWa+jpZ6XS5utTtP5iGZXufiSE1dNk
PyAKPgGAC0CUDneA4ARDhHEsICFU7xy87AVeKip5F6qd/uID7pCm5nYE/poYsV0h
8Qa+XXBdrm75Osd1NHDPIHETFJqV0Lz91oL0fwTcggP8vU+hayuPtfdPkEU1DZfO
UskePLTL/QhTNJfL4WoAHmhYJe6Pcvqh5OSUK5qNiE+MxOt08Cs0IYLQJ9Ltm/qD
rWVLQ+xYLBEyh9s+obAVTO7nlz+v9DKbFbmmAXsrmwYA3Lul3nW3MdMNTMra3f4m
czmRR4BN4MJcA8BdgofH+N1/9pLHe6yYmVzkJG3vtQAZAsefuAbK3i9lGPkrBNAL
tfVkcMDpcGRU9A2E0nPdvLLsA2y0lqo61mnGNtYcx6UOQ/7XErdr7w5dWuYLoeaY
+j2jT1ZKl9Alc9kNhs0ET7I0rsjqyVsjw5xCRYPH6WkF32Dr6LK3UEex9obORk7A
k6O3Eyyyt0kBK3Sbp21LL5Le1DX8s6oeiacc06aWW6dankZw4BA8v4LFN7d2QftR
LMcLnjuxaAG/zAHPsJOWMvC0xESVyMUG6yqikAwOtU7Jgs5sJXACRoNFRp53l+tB
32MVJyS2WnxQyMxKbtEg62k0wI+UkVy3bggyCd6Z0YdOyKi8iSFPxOk0r7HxR4nn
t72QPCfz631D4R10SS6n+H34h8NrgWEA5nGDkO7mLymyCqxHUIF5JPOUtFxBlIG0
NB27rN618kTJ+BtbSoBx1+QgVP0aCKYQFxYZYRGgPmBmZjmDYeAz9PSN7OT6vwZd
bN+sh+GF3mUBK+Fl8kTm6dncS1YfVznb40RGHWlfZkwQk4VJkdtfGGBEIFCfNwMy
NpBA295L3RVvotUMK90RikqSbc0sGF8Lgo0YZm1wQ9wU70P9Cm8GtPrJH+rZmP8k
eH/v2Jw2cX+by7fXg/RCtKrlPqeRQhtUw9QOvmoSia54Tf/SLcQLMPRFoNlUbVKN
HoeOGmOFLYzlmWrjUWfwjZpyJ10T0lZzyX/Qc/GW5azsnXK1EtOf4/+LkhP/gG23
JWxn34ZRAb3KvlzIjl1B5+zPzwcKwDubkOqGSglmwRanDodYt92xkQgeL6Br5uqw
8L82XF55EhFGIyjO1WEcvLB252Na5C96qfed0jvcAO0lz+9hpgLNZsMyqaW7j1+f
McTqdn2ZQ06FJ4oxs18kd3eMGl0k/t4i9JytzsPli5KXntNx7NOvsxnUZG6Sghm8
KeOb0paNSPHXTp4lXbrxHqm0+uXCd+nbyKRD8UpOrqg33zEsORJxs3Z9AEkLrYi7
tUs0p2DfEx/V6FkQcO/PManDPVyHH99cljUtI0Eb1enHidnOp5s2hHNm6itvMLb6
OLgHdgsfv2YjXHj5l/dYDIdup55BfYp2vs3q+dXm7lOoZvQkbDObHUyU13VthjT9
vcjmVma4upkrqPe5vS36cXY1eYAQsyg/SM8bZFtHyMSM5Jf71e1OyVquftsdKGvk
66V9+LmRBff0sncYYc1xz3VRBba7ZAh3bgac8ZlrwA+vp4x44xigr4zNj+PCeukP
fGWgjOA+tzbTjcvHyy+t0AWt+An0hDSM4AKdS6vs719bTZeClQE+6DXTTqBPdFQZ
BBxgEW8ayXjmJcvi1x36OFnythgFsq6RGi+G+Eik0MTz6LY4A9TOcLzsV+mph5Ny
hM8BxuuDXRypS+JNKqr7TisGxzpuQBjeVxROiHX5P+51FQqRv0F7kg1O6zpbvc21
gRV+R/SodHLCaOp2ypCAMJvYSHIjLwALaK2m04t8haaGOWOtiEie4Wu4O7Br82i6
NJTOrxKuO2m2UtYXyM1q7zTR+CJRIbR+aH8oXT3yhsj0FSrmcuvzxENCwDxBVJXZ
YbadH21choHn71Y60TnsmaMh/3mxVwZpPE8+SJtORwmsxwnHQfvjmwrXniIHfWg9
bxDrOIa1lyT/6C1DLKrinayObeGvaqznF2o1rnthDA4CxHDI/Euv28nuzqfNBoQf
lBTfRE6le/30ZJeiAqtS08ZCwXQZ+aJmcMzGagMGZ4fo+2GVWfxzXUXo5mFXhIxk
eWtRby3uBf9cQ+7n75s3weizv+NGlaApRQyyQhyfOo3mcqzPyLxLt7HQPGcWYZg6
Zas/CUnGNACSroVPfjoiQAsQ9pcRC7Y74I8sG/l76myviaF6CrgGfG5jXrl0keXi
kzffwdzQzFozzBhu9ZmAUv5W1U+KCZZKrfY6+rQgsL7rfANzJ2Lq25BoJ2XfQ+cf
ZZGAFTwscGWiBbMgA+2k3D2GrQW7rbFwCt2I9x4EERhXea6hrdJhVTt8NRex8gh/
kTexIMbxX5DJXBTl6b4c0AlzYwtb0VcuZzdz91Ei8KB/VrMuCe1MzjSQ9yv5xpth
rGZxeXxfMy3n6ym/J8rpII+H80E+2smcnSN4vuAb/l1tgbSqNhWmAAecEKB/s3p7
nd+Xnwdn0ZfjidahPJK7iZkCBYljtH+E3v9zHL7jhfdXYjX4Aog6LHmePjEEuuv0
VcamGbms9hKcwYC79EA3cmpok0Jopd8xjf802ePA5wJbArsflQkBT2G2lL0cuLD0
GW3o/XAkxUxXGsRcBP+bYwetuTHbPVAPIR8cZmJbKI6PtXA54RLSfl+AtO80dfDP
pkw+SJLVlZFkMa7mDrCOgk6LEweTfjUCPw9BUEy9UUzjYnaexdbfxv93LiOXFOM+
a0JBPdJzudyCwxUqxmwk1Lke2rupDQRA53fSvubuLmKb2UqgN4eEYVv+jC/lC/Qo
EOuzZCUYYFDR33Eadqam2yBMbC8lpmFeLSmQcyAksASPYAi09psp/AmjV8o94zrK
YnN9jXLqjB2M8Nw4icQDxXrnfziAJDAwRn9FjoTje25ALtrN7RkLGQLK8fA2T6Uv
o4i6DAkTYFWUqAvYcsZSsVsV0iQNovJuFHKj3QgKi7wukRZmBPJHU4nNbAQzAqtz
oS9txOZIVyfTcx3Fog14KrO/A/ef/lUGN7eI1huMjavisWF2JtywSpGxLKwVmPy/
6+YI2sl+Hgb9JurPXBPayBFq0EfR56a3HxMGdQLbGzqChEvMaJbGJviivcRuugp3
PlvPF/Afpf8a2y67ehU41ksAdHTkqbO1lcI0kE2TvRiBGIu2xdogPYeNLu+Gkzp3
LRY08XxCzt32GF/cs4Z5Ow7zV29cH7nz7gM/xkH3g5YTHYFnEO7aN7A90X3qIT9+
Ir8NlRBXyf8clOX9hKidpWX4C1CkkT4VR9TNsuU9mnK7x4j7vHzkKyI1LmA9oDAp
AArYpYhcKpFpLApEoM+tPWYqPn4W2OlKFny3B1AD4Tg25C6pNp9Fwaxdd2bphBhm
xdDZcsHaryy5YlWNvMhIJsii7rOYo2BbDvES55qQyLhB/x0KQGcU6WF1z5aQAp71
e7EzFsrrklFtZOBwuB5/hM2l7oYGvIIXqE+o5WA+qRck/nQ0TKTAZZ9hKXzFUANm
3jdBQJJYUcMeb7PHKHaAyMU6kV6e7vWyYMRNH/Qmi4Kl5/2kVA6QtxLVSCDAudWr
ABxB6U4CGullNCep6UhdW6xA1obO3iwYCXS2Y16dyFGjICZVWa5hUq1qCe81ttfX
kAscivaFhZxMTJI/8o0J+OCUf3U2ndXxjJPTyZDfN9CBGmRd1LwLgWA3mlo0u+TO
gtd6O+5A4zbu5UNKo5WqsJ4UIzXc8aXntBhndHwi7+KbjLN2iVCaDZCboOgOk7g2
+SgyJtZUBAgMeNLBVFe4UwmMSa0G1gzIWlteCXtkLjR+MuUCD/Co4vr/iAnRO1PH
AWAN2CFn8pZl1TqYBtBIljpBeLwDbHatDf9HYmKC+ko4IEr4xrblfLVx7JXPhpYP
/GnL/cPDHrYEeuFjUFFIiH1Un/Pe/nCj3MX6f6b7//V9s2eyx6k01TQjjwoXFnrU
UA7xQ3m7iNpa0FFCRcUrbeE2T8MCRAHHedS/S1fSX4V7gyJ68bK22Z0DB80G9HZ0
4G6vfPm9MHJaMY3cAWiqlkkkq+loEiaU/82ZUDomedxytQoj3Ilsmahg8RRu7QjD
FCtMAxv6bPCB3Gb/SBEu9QjkS9U2Wq6AdpTHJOfmbAnFfS0Fz5QYS5HRxw8MfmUl
OT2QZ8wfKHJ834p+nC6iN7qVOJJ/HwXy6XIqokmTZOmI6m6m9O7b3lNYRWF7Fl7S
VbrFRvfKLebBgJ9Bhp1aNUFo3f88aZkuw0O/cViZinqBGwoiD63RUOMB5mFLIyHZ
6hvqh6ni7y6ObTAXc0WDL04QWuzMiRZaHU8cmKpYF67rJu5GJBmkEI4I5dkxTMpJ
bcu9clJeGXZ7nmX9ebeDEBN8dQRgepUAeXt8UfgcfNPNZiSHNrmfrYKbhUtXnBvS
SsipZZBgJBfY+7xEzNacZJoISxZ/K5AOUb+Vf0Ome7aKWwlAbGVuHAddhhEzfnsl
Z96E43WvSDu59Ofta1zUNyHr/YhCojQl3qWDaHf2eay1C0OI5LL4jW9A5+bi6qgu
EWN7pu4ajEvkZzuSVItdXjiwZM7bPB0gWxjDrtcU0be5oQJeiHSYYDIjtLH/8s28
4SRnSNEVxSrQF8Hgu/iiBCIQ4ThDVImN6qMtxlF88qroNxlbUnPEQGF+f8Yy26Qg
Cll+gJq28SGG6uuZAbt1efHRhWF2Z/5Q0A4NgdE0BGGK1w7qn37g4wZdRgYOItJU
INdWFtagPQop0I39+xe1fgfC5asC2K/WOLxuB6Q9RLg+MBeLQ/mQUXS4zSO4x7zA
HskeqbvbyLg5XSb1pXl07KqqIOG3rwlRxRKbo8QrF2beDV1ynlgc3y/DGDLFLA1i
HLf6cuxU5L+vRLI/w+KzhPtRoKhCPUvRwP1xH7/UvyT/Vr4CGbEHfIzgn/aFDni6
TTCdfHj5XZQZFPx6QUBxHkfSmtlTwoeKyccfrB8uxZLm/5R2mTZYNwYmudHsYdj7
fZ3tAf0iboAeemm5IYXssfQG2PGZrLUY8KvYdcgw5LvDTNymKrIh5Lkh3GyvRCDs
/uNpjs9P5DgwKY2/93vXmsdx6teJh4DqfugYY6yS4yfnvrQF/Eal4jlyNYCDU3ai
/fKS7ZoGkBpA52Bqv7oWoldG8M25qemHrDJ22ufHLa3qkresVdVQ/5YqCnwDPppv
l7+9Ec/KILSdfG/NEAZUe8D0pBIFe3vmxxsSyo7npBztgMTXISWoncIagSU/C0yC
Q5rOYAt0Uw1p4sGNijotMSqlS2QLa92k+gvsUDpSj5/sUI8ujknVrgi7/g6i2FvG
GsEmhxy+lpvUwKQ5me5ig4+jzpdCRmcsnuCeS7GA5Ce0ceTDeUXfkGYEuaeV8fY3
k7gwBY+Yo1mVE1fKZ8uNOMA+eT++fXtR1zZDAyTZVhLIi44UCnYu/hesHCUKSE8j
1e4Uf1Q+kRSZoEhdzANiZEa5lykeZUecFhiUZDXfNzCTpo5CTsyf61JnH/G3N0g9
9mTI9+gTzjaVI3xua8F6/TkJjPpITJlmnewc5kgc7+krnLMsXw8jAE+p/xpnbiT9
LUSKi8ZoG9bIy4FDTC0kXXkxpTzxAzHUlF0S1V5ZJlnQz9tiaGiLems+wXmwfCjg
HJ9fGIkXUIxzfwP80Sk1XSa8uGIuTC601L8c83YgYVJNWYBTeK4rYI2Y8TtPYn+q
szTwTE+wCrl9o1CyqNQRZ/Bcg0/il+E8l79q+SsEAj7FyqFPARbENKz5lfa38MRW
5Ye/Cc7Qr3tqwQVjgtPMxH6koEh1m3PBto3V70ctgZvpV8TUhbZP4JrDu27wm1Jb
hd8HyqbqUvVMFmVWodV/EGdYdjrseIw37nNaFqONeFZOIDlY9LX0d5apqqu34S5g
yGSbQ6t5iIjd/W3qTBilqbz1YywmJE1EC/tJjeZAImKyXMfIbW6iNpexIbNozB7A
3S4FkfGlbvegrmLhXuiS1umzlAz0BcO4DcYbCaJkh+amHITcwK8qN2noWEHzSQrN
uSBdNn2Jfb5XHWwdDj4UCs9t3Vdzqpujw9DBI5Q0CmNkUtQZpox1bJIJ7EQab0Ev
FlaRn1UYp1aqSo0Co2fOpMgsIGK14wNz1sl3qtlvstJmT1yPpzOlymjqUaA471rZ
AUnzXo0AhROB5ytlsQsfXqhZVx4zOLqCYKQwYH2MCb46VtYuN++bDjN1f+jLa2Yr
8tFi1J5PsymUgOmBlWz7jew0QcdjB1ulMGJ1QHpHAKWaaY3wcAxsXdEKi5Oeipur
K09ZYTzktFIVPKiaHMZmK2xO34nuHLS9yKWIkFzt/dBS41HpaSlqhbn5/WM0pdGk
Xj+VQfpvyjRkW/zhKBhhVMXFbmY5N9rNfS7ZrP8vYE/xMaFWYAAILPVZsOizEcWM
2bwHvHuFy+fM0h5buF0iwRnRhyjxxamUCkBQ2XTrmgBqq49lNxG60SIgDzXHUj3i
Kqz53lgThq1Shk9JWKW58khtEgSDkaTf3quuNPuaM8qZonUtowReAEqVXS12YgUk
fCMqnWz/iMiwUa0bQiK6KVuYeME/m6qHgjtdYhv1bLkxh1hGhWZmpzorACmhALTt
Sf6x+/+zTfWDHpwI7qut38r6KqEHV5NtSL9djlK3EpIMIesLPUYvT6UNd4OnpGjn
eDfSm83aXkPt+1klRMbOQKXwG8nRJWVLHhZ2QnhGdKLF/qSVD5uhgN6W3SZo1V9p
4wIv2pNrL73Qf+pKJzXzHQh2oDaL3q3Jm0Xc7rwrGPYQVgq8b4aRdTplyOyv55lT
Vh9X73ZWgJWeLUMlQjhvULYVJjiThGzsULin/mQfGoc5AnTGHwbdamZU1MVObi4C
gPTVLlStgqKPryFWBb+YsOYZ7NfnqmHW276dp5NkeRwDKc0OgXGr9cOinmSRHwny
CIw5xs3VXzTi3Fw06e0TvHnMvFqZsesbJN1D2V9nr1/E0a2hNq7/SNCvHS+3tCGf
py6kwdi+lCt1Tu3dZ2YiNJiRNK/zBo5Dh57RrJrbnPtF2L7tl9XWZokQ7MMGjLqa
NhrPvSP0sVAAWfPMN43/NaHnRVpi2OcsR63SnMMNfF8KDKys/NrSglY13V30XMtB
zB7iWQI0p7hpTPlWm2GV8zPE03XfythwjQzYeTwyRrD1/rhrjnpRpqobH0u9oXdC
iCrpaAXdufKcv1iFsFmNw2eW0vOyjEjs/5pXoyN0VWauTACENF/9P+GZPpGw3kLD
RyI+cZR6ZtxBOcDv0bIQVqZ4lNxESLVTYzaDtRDhHZuG0h8Pz2dhPnPg7gy0V3nE
mDPFriE9dXt9tg2TyoU5J+M600nWne1sum8igDVKn4mUIuh6/xjS6bvasUdJVha+
n90Xfy4V+jVPtB8IsPbmTWxprX3Dg/IVw8ztd0Xl9BvvFyIYpdkUNPxiMB56WLm1
OkHS4hex5vrCjpBHZyxNtIVIg/wzDIJvkO6tp2CWuA8GImLZnNTmWfMe7/sZ2Sqo
kRQNwxgsB5C7OxwsGpjtVGnJTC1+mnalXGXxQ5kUQ0uxb9+kOO3HcSv6zW6NrMc6
HnhrqoIXohdptI7BGniQpCNzg+7ldSYu9qYOiIXox5ckhMzAYa9jFb9T8r1wBLA9
dJLzDTXhojQNAr23MHOVXq7N4QznzENPGD6Jz82qco8hHFcV7ICZq6/FmKUqhv9V
B9nZfF7mzgiKcnp9iCEly4cWFYvYtFKDvhWLX7h+SciGOnxZY0HMcuzgxR0p7iiV
VoNaoLw/MzpKO9hZWZZz+TXMVqw2i9LqM2D/inUs7tzYz4oTR+S7LQ5zu/ZIrzBv
m3zAVocA6ISZfPzMCdkRzc2F1O/tW2yXGm9TMt46MipPcJh5mv+X7lFAeKE6lgYK
RqmUX41WDrfQwbIoEGA7OR2EPDByTg7hpotPyHwCVJl7Av5vmH/lyAi2lznN4W08
MpA4HkF3EvXA8X8lREx3AeeVFPGy0NFD/T3JHD/jTfrs6XYvJwD1h1lNtmbR4ZkY
tLSMtX4s08BU3Z73Ky0JLvC+YV/IDrWGI7BIpefly7UF4MQq5tr7YJQpSIQzac10
M7j8ikhLeh7rI7lMv32cedRv7QYmu62zed+yd7HAHQ3GwZCr4MKmXRlCUNuhg1Eh
b0vc6ybPdZ4Sv4Oj55zl/mRQvGXjcuwB2PNhqkL0p2GulelC0gn/aTAKHdw6s2Cu
y9NEMPrTvwbYE+eW3R8wOg6EJmd6cdq8AYycO84tKjJ3daMmBryfr3AEJckL84N/
9PGlvlEuJwWKnuMtlk6/jAYg/Ji/KGXoDZ8S77TlgMcUC9PoT6FOqLyGKqJVEAkV
xNyv2B9kC1lFK4PyARUgE/RG1I0UlLkHQD9RV7Ot3ymmX7iEobHPZ7pxhmxDpiFV
LE/dYjjFBuidK+vtLezpAtLAk4bWoiVR/3perez8a0sRMSyglMQuPak9ghOCYbi2
PdltlITCaKxLpkEOq6dsGYWE5CHQF/oLNcj8Gs3xYlqx3ePU/bnEq21Vz9Q4515J
GeBvlhFPF6Vwo0DBEMn3GPCssxWQljvy8wwm0c/hy3hHIV8Ea9Rs3vHce5L9udrD
+pKCgMZKnfHdJE6IsoWYxpJK73etMqp926f318s+kuwviq8gn7TuaeDWO5qSum3b
EATF2JwxMl7Ysk+wL5Dxz/NqjN0yyG53LGJstZYMwgO5DJYslTSWlQgM0hcfz9ax
gbO/VjNu4tuyHkpLeIAC75oOvy8hCiBKh8cf1qmCCaC73BbtD4kC4QT3UN33AMPB
UFZR0jlW8RhW0M+64pJtZsEXri8j1AtFOHYsOJo0s4HkfFIJXkxiiD5L6VZyIgsn
C/JmieKhzchUaFpFUM4TQloR7tu5ak/JL1yaW+ArbqrDsishLZguBlIOD0o5QFaH
z+iKzXkfsxW8EJAMS48ykTpylA1k+RzdDyo4DGhFW8qi/+RX7MVbrU9/1pmpDVqf
WEnNfIQW2rPJbswch2FCfzwTKy3jz1BEtGD2b2PlLH7R/ALldYQQkawsHwMrEpWX
hzz8q6990ISwMiCKU+M5oWyCZU3h2f9yH8aS6bm/FFh/0kk8gH1OmNjy7Bkcd2nP
/xuftqzYz7WsJoVY5qhm6YDqMed2j6v7z1jlijcTfIW06wIydJ6NXg1kdmAPEVnk
h4GqLobZmsNBtujyc+BqXlvE3SlRjA9SwDLmIgmjYIQGwUDX7sKbXfuXUheJZm0L
/OHMz3ZL+fEjs1+5tLt+7NqVd7e4wUh33Pq/ste6ODOckyDPcSLybHvCDLE5hHvI
m1t/jgGy3xd632ycJh2g+CJNpVWNSKIA3LZdTnlITZ6bHRQ4/UpLJwgc02gehxy5
VGfD4erRk+phvPrVeLVjCmgr9Fl631F437PhDAie2+M/g9QLlXcR3HUeG9VW283O
HNwUwXwZtfBUlmbbac3gxIGVT+AR85e+W1OtFbjuz14dZT/WFBYvf6CVB9FxMUlD
lczJUrInWr2q5v9dF3AmHy/xHAfaVZ6mWUo9r8gsy6F5yZsKXITZwz3lMa5oqI4t
caieuZG5fTBR1L2GMwK2QXQdUgdB8InCU0ObAN7VulgZDWm0vDilTAVmowYGehoQ
Y9uRefRvTk5d/8Plx/CvMCrbTecyAdfpNDYbpUBonnyRufQnoqRKZgpPeX9wKBFB
au8X5N/jwH0LytR9CyP1X0kvhKzQMCag6Lrnuichqd3N1Ollx7mkj84GS5CQidRH
t2pqMw+Ao0XW7i2pLf+A+H+jpOaKTsl4Wxax6SEzfoOU1Ixz/2DVntCUfdO3BxMs
4lEVenujorK+EKrrgrWqpgx9kWe3km96rgIVU9/lyYH2ir+LYijzw07kGA6k5LT3
xRqpbuvCbtdozrukFsfE58QE940blH2LlLBpJ89t35MF66KpbVp2SOCG2ipHmlEd
`protect END_PROTECTED
