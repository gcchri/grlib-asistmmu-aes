`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
249ha6GCqNa4ehtoT0K0CB+TB8X1ip2atCC3Yp5uhgxRkOewKKHhG40WOgUhUVe6
QW4tQwAPd/9mXq9bpAbScrDY4IIZ9aROeOQeWvb0kG4rpCAfR04DlZXC4Ui8Ssb+
6Iu7s8W0PQOY6aOy/DNmx6N1le89gu9ezxYyLioeD9AsIQsKYdP88qQJ9wYqDifZ
DAUXlZtQzY2OM6ydCWMFwyY1Dg++HEZu53MFzOx64JijT1Z2rNWbVlRTGa7e8N7N
IQivyo5VNxf2JgRqxzUha0XQWUASP5Bgw7F7wZLlTewH0LK+VyyjWu2gj/iDGMEB
Hgww49j2wcZSIL0MEWfVqgFrX4aczVsJQZKVceAjwIHZTBblToAf8e2Qpd741bmj
IbwAZf9rV2D0FSeziMhdibdaAvCc4tfFjg9m/OH+NwKEE4vTBkK4ckOEo5Et6e+G
StS9LuJ2XcqBHqF2o/krF9ZMIQlEEFVuDCmOTg81txm9GOhcbcv2Enn6kQ0GAU0j
zN1hE6ZTj84UaueMmyc7oW5hSDfcw/LTrI3fsVhTB/vkAQBApQ9aH6IJjahPw12m
CyNZ3DWtn509A1xFI3O5hM9VJcVCGWZ+GB13J9MXQ7+ZykqmsTskKvGnJ1JHDQCB
ZWpq8xrrqLDdfpQ4eEkvbCWDJFi1RFOGAZajFd5JcETxrETy3EC0M/WU4vRvppya
jhNmOcbHf3K90PSXJ9WKv3Gcm2XZtd777X/lfDu8cARCTKdrTjwh6CFnMRGedhtl
sMqc8QWWM4ryjbwfW98AsJsMFpvJ0ZHkTstsPtx9egJ/en7BkS+Io1WTLT7RZ/4n
bLPEAMk4MzrScHh57hBrHYyc6ucAywW7zuTn4QV6y3H2XnrwkU6yONQWgyu2UK0A
JgXu2i4iRLA3I8ExTVY+lk7bf84oInzesaJsflv3K89gWY8cPtN3hbKXXQRG5U51
KeXatYk/09+9JvFkfv4oOz1yxS0Veezo+zCFXp3onDEl+DA8pLu4Ph3v523YmSa0
tPh8IFBQq7oK7YttDYEFX7BtNee5vfcqhQFkhKXzhki/8iIG83n6P+qp5WELe3ZU
mTfZ2yy1IXAWS63HAGS2CvuzGp389tnAPKkS9EvlA/ZV5HlAXojS5ARCGGztw+ti
`protect END_PROTECTED
