`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p1/CpV5/1H82quU60yuNBIVkTYacLpeblbEKDtllmykSvs+skL+t0cy10vN/dewZ
vMikkytnC4Li55HaSXyXwL97Rge95KNqRJ2EOvFoZ+5pYInhMenO9abGDYCcYILN
57dd+eblQNEJZF2s54uc9fhi+CfhCu3MdScjNIsXLc3cTl79cko4MYlX7TKwVep3
39sb8OO3Erbl6CJ4tJexLwTl0nmIqNl4CfIwBXpthiqkrg/IZ5/zkD26d5Fyf1jx
iqP5USNE4gOedp96rQuNNDfhG57OM1s6E1bGsQiJMtJ4BXQlNHD1vH/K0SKEUrd0
skzcyuQJW/LbDj++taEe7uMCNLToA7XcUUqPvsNibGfWHWrJYPPIbzchkSgwVEol
fbQqsYaVcQAkPOK5Q6N2lSjRXLZAhqqbbn1tpkyBBkfjY2vDv6Rj4FIqV8AtEdnK
mg/i3xvEM99Ep27JyZ7qSR9zX+fSrzYbsKgQ2Lqvwf9TxQhaFlsOsy/+Dxj9X7zn
BNZdaXIXWrbE7c5W+PruRiGQpVsJpf0AAZvIzaH8sAgY8aBxoLca1+p7pMmVPomd
Ni36ZYSvqbuLrg0OV9GxeuucuRqtr1FD/N9Jdwdnbpw/Gkm1LErXnmtv4MYadYCv
E75KxB8gospcE1sPZijrqcx+ZlxcncGW8WWtabRGQWqtX/5YMY3UP9ZVViDAkG+d
3HVZfhBZJdRKyT4Ge8yOJNu6cCGvxIOOHvt6rLcI1LANjDXIWSVPjh8cHmi6718W
oBBsSwIUEgJnmFrX7CbcWEQ13kaLY1J85058rZIhzetL/FC0rKkuKwTAPGYw708K
lIBTyrn8exC5mppuVlpKMxCVnWo98IIYa2FuLbswCNvOlu7ENBFvwonpkMDxO6zr
V8G+i/YaHc0FtLaBSxU4rEHakuZDgHjZkrpiwsAiQRa9mnpGeONSuSZfWPZsOzTg
7prrNngD2RLJpcB2ZmZ/NipSByE45k7pR53phfCFXLwXimuBwzhOPcyZmYyN6XI4
tsdVO+FPDg+HhzDdwmsZ0yK3e6JhgliwanLiBu1IYYwI6xlhoxaCyGgMGPryh5Hd
H3JTwK8QmXa9UDH7xNYmzF0Y3Ja7kMcuJLdyWsG/FX0WvjZlegusQVE/QrGEaCS1
ch/kSfAvMnV8Y1DY2pcljeyt4iUYr3nL1iZBDn5rn8bh9zc6eR/OKB4z8VaLhSpt
Rt6Joto97mw4ZaQAbZNAL6+WFlgczBCdUw4AVByICSZRZe6OzBS9WfWU7VNn2uGY
o0X/CN/D17Br0Wbbr1lsHHPJhLA0dYYW19c5Efj7VgxfDIc4WTZvk96Rr0N64Mfs
SOlbSa4DHbQpeJ/f3fI2UVoxEflohOWcKouPcuxjf9ShLi0JnGL9fCMOl2MwnvNF
MgCXe21JIk7IlHy7aRCeNrALeIRqPKs7qg1SyUqbtw4Bgz2XJUdTLTwUWxB7rErn
fawM4nYwniz5YFwe0aKwtQ68tCWhIbSPZJ3wMLVbTwIYX0utWtwL9xJARnRtMjwi
kNaiqf412hNyDEbYY7b0QHYmCx4jHXdsFqxaZLOhipYnn7cBEQhD2Wb7MHNcudkh
1FuNg5F0NgVUq6d+GO8qXxZJZxkOyUjtulMWnxopKTCVRwa3CE5PhBDaTsau7VeA
OlcpK4iOikV4UJTJy7zG3ZGS0F8DRKMPkC91oJgHu2HnD6XAAl+Ycikb6nYL4dO8
oLiSOjPWFOz3jILMmHdBbnL4/MtYfEMlcIPLDKl8MBYV2rE9mSSC5dlZwv6g/JAj
B/07EDh/FgCqNr45RJJk5sTXz7qogadwBl3HTVnZy3ReUwRcbKZ26tjHOgedpcvl
5qke00hClCj3ipdt0+hGVPIKLrgbCtAos2oOXiWFkVchFSILe6ZLmzH6znmvbP4Z
Wy496sjPfQy2WBPFlRPsYQ4U3BzXP6bgsAXfOFrcUEb7GI//Gzp+3lWKe2ziD5hy
aImqjKIfxUzmZSbQ6/crxABRzBOJCbS8e/SphMjFnfNeTM35L86dm2wH0YhXj7Lm
ihNy5SJeKMeSUKmucueBe18StUgKADszJy20VzCBtK4cd8LoQjDzh1l9Myvh90Eq
t3W3g0BfQYPEH1fUrE3V1wTc4woUY5J5YeQ0pDYg+n/eQfmlLREdq8ZzTyABzewm
b5oE2rYAkeSkZ5qP96iub8uic05Cpfj1rtjQb1Ye0dxQPjyCIB/Pek+JHZ45gJtk
m2m/zvyl8uff6RDGqJ7NMy8LpnwK2RwxZQ8ZH6M2MTMt+eAwneSkLtqnok93LET6
Lpo5tWUbWBqaDe2mxnQulxTeHslNqwbF4I79zJGpTOB7C9JKnWXmAzUcCz19RGIM
TbF2qnsKewE+H3PPG+tN8aSInIRXkMokFs77UUubvO+5GZzO6/+M5Me+s/xn97iM
xE5kvlPFHPItim2NtRDDowCwRmv+2dP4q0vyAJPVsPg9GkbO048gE+mTNfNsAtqT
eR5tS8OWMFgs0LgFtxIqvmGEdiL7enPai9gGPV+xyL1Hqx9Q4n5JWrXhkBGsKGVh
HtJNCtqvBn9iQ1Cd50b9kki4AlU/1KmxEpWH65Gz0AJR7CD/dyj2ndYeGCxpm3R2
rOjau0Xf2/twPWPuCprIWbVy2W1x+vQ+BaAGdPhImggHikeHT2dGboV/lGECTqOM
k8s58Q99+hCgqIOkr1T60CmGGTfCEAbE7h7c6xIsP9VqNU7SNn2BPPuxB5HiR9Vf
4xu08TqBATF+Tl7Wczs5VcYcQyKzC3ZwnIsW7K0cjYCM6fQezLlkWT/I30IA7pnM
UNUp2BbOaClPlZaYwQskKAmnuNwD+Nz/dMcn2eZR0HDpfkPqBz+sA8Zj4SImdJqB
TMEv4SZraYy4CaQqkBSU+QABJL3jwEuuaIOm9JIpFRzOnl4TrD8EVDIrEblGkUFA
p7uTVV2M1ysU8iQ7rBuBSypy0UAtjVEHQQrqp/mOFFhO6qHQmp9E+ViEdrDpZvWQ
gaDXxtkkVdOvLhhUP6hP2AvKAxWbNetqkapbTyn1MkfWVRjmI9N5IlSTdCYdIBDF
V/u8DVeP9W8gZE/dzOPKkkzBwjgi8YKruPOxAfOcbBQkrLJnW4URi8aTRzVVWnV2
aReT5H9zi9YFKBJ2Aou51HD4gKG8BGYrwkxZYZ3KydF5MiD0n4Naxe+PIbX30QId
C02F219AJJvRSKmqIbJeFVQf95duWL2tQ5LjZf/uBIEQfOjQ0+FUPg27tJpJO//F
ASnumBW4wmHybFSafg2Q4xstIZiIHKF3gSEte5gbNcgfV6dUBhN74UfVMhanVhez
1MLYBsGxMzh4jiUqQe5H7V/NumWVhkcViavfQOj+hTpClrMVzdv/tiUTiR0m0X8/
ad/MvpjlKApuuAoyVNM6aZxrx342M46fn3t6Yav2mU51pZz44Edcg+KdW1KFHpwK
nmvR9/TlTjWgi2I9xKjn1koFiH2YBdJpKe62r+9wB4dlgVu9WGLJ8TE9G1HRmGDT
c25kbcboW8OxOlcZvok9AxxSjz2m9t6jAvCbmj2puV2478WVJRuwwcpqrnVyXY2H
KYthh2eba1NMShuQfEhQa/1rxwPMYpqwNXns2DDB1DtmP81+fbBA/C8A7mo4HZ0j
uGACIMeciWN+pbOYg0aufmiSG+twpXseA4bgyYxFfn3il/HqrbQA4Iit4X6zqOx5
3JgCB+r1vTvReboDqdczwCbdcQJkHrPszsdGBpz2EIYmgl1yBI3jblIMSdG05EIu
tSWW0OdVVYcl7UOi0KKdWO91JyIFEviPf3rkQbB0N1jyLOIzhq6RbjlBudzVFyN9
wUTSCMtMwCjXqh89NUmxEV0rAGxde92coeF9A0tc7s6O8HSqtgNDvK2TH4peit59
BW85QwDUfrJns+2fpi4NIAILPv6TJpvT6336pILd+gIi7j7H2crQ1c2liUkT+EmP
zdi8QX0A7DLph6TGOtaO5RAZjMiPkJ5OmHfppZZtHrX/Ct6usPaALJnwlFsqaWWW
Fxh1Wjsp6ca67ATzceqQp9r2Yjn3p0x8lUX7+X499HH2YlvEw0+JnbCRpibzrwtJ
FZHK0cpGyAEME1GHn+RZwRj7pZAx7WR19hSHp7aDzuWBWsBW0ADpHDnU2S/zM8Qt
1taqYsMoZPuty1EdnbPI2aHfji56cvcYvTwXqRO9zuLxwnhQ1ALtxz/N3aSXfepz
HNRe4ekXVGPrQzr6Nhxv8a7O87g8h8dySmp1cDQDvzo2CZ63DUjs31pnvFHF0TQQ
icjhkZWyKAlgsfBNMmZgDTtLegQdEizHMWG0dueZWbkcaC5uZViPtS7RBzDLvUGv
/n4PR9nFA3/5XiWz9gAwqzzaOkGK7QZW+WASKYtsbWlP6mhE79K0HBsNbTU+LJuN
GORv4FQ0WSWe+/dfDEZeOJYiGhjoaWmFonTuf39rTLq6e+EYbMyXaqRHfcTB1RVQ
n7O1nlC0MUc1+2HaNE9NPp8TpdFzfx7skTCWWYO3JAPK5jzaE9nyrWcTag/FFU7g
X4p6SJvhk5Fs6xdRQcOw59ui4zCGClSHlb8C4/bo7sxbjVtakXTW+1luy68EwJw9
rUJskUKtZs/fXvWhgdGeWSMEvQFIvecUNJkC+1FtKWDiGQ4LsbIyXxDOZhsI4XgJ
dEmTV1kqDmWTIXLYbnpycz4p8LQtBJdkzc4OoZ4tI1sFEExZ/+EoViKgkFHMRpsD
2+X2Vq2UoH3WXw6XhgdpU/wqX586pvRtpSshBb2REVrwkKphCKd2qyCrd3ADzQC1
LjO4A7L0Rta/KV0c37Qc9n0grk6KbDSsMB4upfsfmmhD0DLQNECdQWi/GllhTtoB
ie4ADXWlN6KiJ6ZUpc+QyaQ3JtBf4Rn1s2r9IPg1qJ4GEKROU0bLAmZ8NRSLuljT
c5hGEM1AtPFi8WRtEud2XBI+ml9QiY7z0UV8erUm7BHBwWXhb5RL17ep/Ha6JQ1S
m5W2d1nvNimSEn379I7AFwN4r7ojc4cO6o0U4lMgaUQkMBWIP43NZCWv+arHgvi5
4L2Z1YOAAEOgSd1S9m6ADty+WKcfE3apEe6FBwZbIZuQUDk+qnEOwJMrrNt4SaSI
YHnJ1JoFq5zytC60N8seAdD7mt0Bc1A1WsI+28ML6owQxsY7+xBDFKqlWq435xbb
joLaVUhUiaHtmSknjai9PBgxy+RFWwuf1Drdto0MN/dezcQrGYEP+hmvO7WDJ4Vr
36ekJld0CNaHGOUDLLPt2XIxBFWK3lhmtYHj6cRzP1NIQPwUat2bIYg0m/KhxbM0
0k4pfeMGJ3LJ8ntLWBr3nCm7M9601kIQz6JQ6yWCXEmqdMD1G2t+2lEP/JTtGNYG
vvASM1eCEoAxmn1qF1d8sTjZ/Y91qCynU42bfxBHh5VphlO+tGhyb9cl5JaOiiOD
JzwPHym9nouJfM+KxhJ3YBmvx1OVXgX4gaTyAaUCHGLoidmZbfwyTPpGo0EDrN2y
ElHKjWMrTZlUPLZ3OgapaG92CBQ3TJZ+qosLkiN+ZchEDO5h4O2SnNIqs94aAkrg
fKqB3jMV+KOz7QclCsJKhvpSMng6e/rCDsXj2lWAMAl5ZJUlfaO07tJOgbucbNoU
2cTN+M1xn4V6SW6tgKmhSJ0q+nHgE8aLjJMgzFI3F/4gqeUTqU5bxFYAOk+0I/iL
DT/CtmmnI6LX14RU5iHiou7eB7ZQ3Fxi2EBj4JmGKOER3KkYlRl7rpDR3/KLmZnP
U5434BuwcQF1bkIPCQlbLZnm8CmD8/0wXXWY26Z6cExw8j7bkZNhWcXkilmxaKM0
FEH4S80y8fvKrNycCjdMJCOw+AGmAI5TNTKULU2WRDwD1wu4HkaGC/1W3gqXaBP9
WOoK+S/zvQbc4RJ3qZ/DxqV8KeuRBuox1lmbQjbrhqLD/XCPsDIP4pXRJuXWwo/0
jbbPn6rAxaK9ningTj25BB+evpzsS1C76YaN88vERAMFCLLHLhNKcZ/P/zEd/P8O
tUgOw+GDUtSwJdMvO/VMgBFOTK5TSWDo2jXHc2UAKOoEj9BUJnxojdEr4zFoMtyn
9scFpMHMg4M2tUdLKm/u5GTgFCyLMep5xZTNlVeo4jP1Zs8WXNaYSNC8notuBGuE
BX5ubpNnQdjQVE6/8gb4LPpTyA7usW4hpAjRqbANkzVyovpjN1JX07QTzEuBY2tb
Krig5XK30srGMtGxG/UhGAxb2Qnb7sX8sy+I0VuWgR1scKkHeuVsmEw75uIxegLq
egv880Hn4WDSfpxYSQPMW6nnqfevOKB9NlPu/ax/JIpFHCiQwtSM9R1wZ38GKb8W
kNdXNJlBsvA9sB9iIhTds6nXBT/wz8wc/bjqq6n58z0VtIaFv2OdbJeTXDSPwE71
M7vaoX6bvvyUzmjmF18GTexBV/TJ5F++UqxF3b9bTJRK8SKL19q9L1WDVH7Uqgo3
MZcQ0dabpbNH9L/pUkHxWMHAma1J2Bxmjpm3BhyozGLB9vfDRfOSf4UtVpnOJIVY
+y0LjRVMA1r4zcXvca/nXtzdieBzGKpd1PlqRf/0omsy+yTors84kO1nfJ+sHoDl
aTuw+nCGROWtPU81ST8HeuEMF8Qw8Vp++KYYZegzuA78YNCTeWkMyJCx+8YKUznB
I2gJZEp8Sht14tDwrt6Yi+cw72Kp9MecKDnw9gxSCHTRrPdwhbJfS6VrpJ/Tne4m
EYdqsdxPpmke6f3ikzQY4PTjbXVf9SL6WEGi9xPJSTzFabXnYyHXCkZQyiREH9um
qrjJmCFH3trX9Z0dpUsP6fvjN9MnNYg1a+n76JPDLjLLE1kOR5f0A5EkWwvPN0D8
3ij+2kBzyuoQhwqx2irOzRE+tlyokMAcq1ZDH4S1YuritWYD2zkYjut7hK6U/Kz0
M9r+H7JGmdZkRPdbypmxNrurPSP7yiu7VncBYbvbmljZJotdsTveoK189xLS+ehS
v1GvqRe6xpZZ5qf5cgiAgXtFMFmi6UonaSQU6CwTC/+HyWXjNIQU33Ams/Efplue
ttjH0TNLy5GiyQ9B6uOL6ED4UHFdjRvzlqetKMqssBiGcwdj40sNaasDqgu/C4We
/gOu3vWkxIYDE4V4iz1mOEU3mtrVUGpSZMLbwfHbxjigOwwnCrSsd16PQMjBU9MT
l8xcqsvv2HrWvCoKV26UQWACDRZcrkqWVkyJqCgly0+2ikeKWlvMk6dZLusc4R94
uqvzntgXUSI7oMqo0VgvtROF9et6RJalYjtehxtPJK8Zl5ttFI0I139v9kT3cdFj
SqXttzi3RaCp0EEmZM0wbQTlAeYP0uOENWkxqtPo/e5sw9+r8EUxN+kMSqux8Ic6
u2n2VETS+BDhJgoGfe6RxxbngHZojbQ4CnbF0Wfg0/PanKH1Kc2fhnuykua45u/N
Abz7y+U1dqnz65KU/PNyjhfEznUS4aT0nO8O6eg20qYA0sNVDeqW1JRm3j9E9m9U
731XEUa6JWL4n1Oc3HchGKZVg7Sc4xD2lA4Ywkkwz5ZAI65Z/cAWHENOQIa1J55m
SQ7XySjO2B2RilhX9zli3gRPRNEQXSubftAxt9fPSkSCAb4g2B1PXgGSj7A61ndo
J6AtAcyhZRDw/IjrTvRe1eUExJfITNEF9BHiFBsJyNjs5GmIM6wmgn+jQtJI4H86
TQ/4ErtwRLoIj0j5eiyTSSeS14bYzlNeXFgPgERj5RnqSTEvQifTQ0oohzaoV0BV
yBhSgxh3fsBMVaSZm2wcVD4beHFi8qgJe9eX+1PQ51W9470yrKESxQaxK6vw2PwA
5vVVQKnWUHPYkDRHa4cjafUIvLsCaXmBxPxbcyeI0iWB9PWT8a4TH30TeolbI7e1
tIRIV5CU5iMCEBf3SgpwksOOgaJNM4E7teRlLGMCgIptaCYhgDBpk/08LqF28MOm
jbWLPNVdyMY4U4nOpncX2tvbWcTfIx2y0rEEHOUC4VFRY98fuslvn6QrOy1HF/8f
fPeKaRtOscEq/saPoPqVeCt6BN/mCjrTMWwnp5PzcCeGSBSE/6N2pAZncAx0Yj4W
r8nFHhCWLWfd+Y7jpXFLexrAL9fdZejAFz9mVU2h+0A54FYkOatBNLFcqlM+bya8
z50avaG96l/H+vLJxGT1mAM/DnWbHwjGRPkhmjodIrMkBooYnzRo6hcDBQIgWYL6
O8u6kvHCfn0/IJJq12iqtYAZazuavTFd5a4kEgL7xU0rjrN+ehFap4IJckfgo4l+
OwIhkk65oKxMagpZFITD0YMmVU6KNssBl/eNkpzZMsCW9cBtXWVBTJUO30q0r3Zf
3GoDYa+Zx0nj1XXxck7A6B/xqTN/o2W3xeL9NXSuKwV5bowzKaz9C/w+9ypcRGbZ
P2Qcq4GZztpnENhGgK7SNiULM3jLMLd/oefhGemS+yI6CvXWENXQpjLFm+6RH9BG
GnK6AVFinbsZl4K8trSLCOeQ2Kzq0Xu0sDdNtRBFLYp61mS8ApPQLBC/wj5CpE7h
KYTOAYZTpZcOglBAaBBZlMq3Ku+sa4qk8gOHGr4WeC/yxQsSjcS5TpOWJZxW5lJT
yKrGwjCMaS+vlgTJKbKG8vfkDfziccdHKjofUL0F3V7BLtljovkPz/57MiGRdByc
rKFwKIQvgIapppD9aMs4dI3lvcGPL616D30Rr1J1uNUhGkh6l0esO9Xu/bVdR4wy
0puDLV95nSUTu5RIYc6zmyRpxbrnX+Oee6h2ePHxToj+EsjrLRjiW6o6TDoXb+wu
GGFoNZqilVDCaUlvjiOqnB1v+1fhmGB5AFAJYjC66EQt9Juzd4KjUi0if/3lk/vX
LNvfamq6822S6qlOzxtNIr5OV0xYNgsS/AJOLQ8Nz0mZTSxnVc8wNjihd75ND4Kl
dhsmwi1RKTTzMoW42NHbzU2QQa/nKj9v2LVnQA6B1Vq8cyS7t0AkTbwiv0mTBOUq
NE4RAWIzj09YQVmN62J+6ByUESzitwjNQg6OJIpl1rTH7tw0eIcOlvu7haaayc8u
Vs61OV6UBee0mslDMu2H/gOHQX2cWK9C2HJ/zDclndufrlyUYCNSUmS1sN++7UCf
eOc4UCQQSMaIZgv2+tTh09KUiRdh143ku8d931xfRSUXKKyx9x06b9hJPtRVVzv8
SzWfcPApwF2qSUt5bUZzX8T13gCJxape4XWTql6S15cDhs6Kzybgq0nBi489CSY3
enfmPdczE1uVn6jja1/v6/XcTg9kjsiLCTd1MWdfQ4lJJPlGIla/RSjvRBBTzUYC
GgTgnCe9gFiErRdenu7Kwy11q7TorWYkT3aWEckOndIHnSpmXFqXldRu/IMC0yL9
AvmAZUb6ZCW9iByxQ+kDos6QVJQwwtIdT9eLAWqP74xIwaZpwezTUBX6vsl0KNpd
oJB1Yg5a/3yZrUxxnZE7Ix7insAu84FessSBT1uEjKdDv7gEj0vCXLVssFSDVELO
moJEezRzWmLCnBiy6yB/MDIz1KXV96UW0IY9aEHXkOi1tCpOnI1L/aE49bPkbyqY
YPeWG5sEHLy7I9wa0gy5RlfdkIv8yNpN8CqtkiypafRIO4AHc6uTx5OTUCpEqND+
mF4EYWvu/2kKxZN0L2QTTpynNjewcDHXlv8iNzKJ016GJkEtMN2KYmwdJBg/s0Wo
nLJbEUI36F7lbznguGpr1MxaqrQ+BwdIrvA6yoJPr5B1mwzyC9GOXPTyZ8H7zV3k
n9LevQlce7kXORu7BMF3FT/W5q4H06nGXhW+KmRDuaCqetRjpOIVPjKjIpQ2c9tC
9gBc9CJDWUQXVsAvGTiDGegkftnIiTdoKoEGjqrSW53CvrAVKYCec0voC+kltYSk
28CG8kdQmzwpDWIlDYXk++YxZP2t8INz5ZdzTyPZtiTupMtK117eOaX6cDb3rJ5g
wSX3XjBqUv8yaH4/av8vMhCfEE5cNIAIQBjFHFOF8kGH9BefYHFyBCFG1o0iyE9s
B4JDXfb/k82CXM1CqX0T2Q9dKzce0dUgszEuZrsFR2LD+ap2TOF1GT21wGmKp1O5
Dm6mpx9q/0ZfFDICkVyfq/SF702eoIeeSa+NQAhFcQEt1OQTTI6KmtuKCVjFPrrI
fTMNUSbgUvNe2dwqK9kdBFNkF1hqfuNKeM5chy5gBI8zOmS2MbabgWDMj/L1sFwg
GQQfme/eszWywUIn+H3kJLSW0CSKfu5PdpKOZEzdged/mp8+CaJcjALsxCkMt4JT
rtZ4ZywIKSNYThByaTkzX3/Z3ZIHAlvZI2k5YMXazb4VAr8++lWhhhFXrVHOG0+e
FIh2OLmZIQM5vZBZxITX8AOqLyp+JzWQLBbF4OSqnaB97NTJBtvTOWPBmGrA47rh
dPMcK+w2ivPsL1T79RaJvlkfZ60+eBQWxXm1yPG00pG6yPRsGP4XW7fFSduQJrfW
PPXHDJukNbuEHAkIlc5AMiFHLQ5kwDPVPsFEwDhdtKO0HcgLuhpMEGytDf0f5L8a
GxK9dvlPtD1Z+I8PH3M2176QG3mN4XBeQ3jvBNAHtmFamAgdCyr5foGtYT6l4irl
tt5dUhO6k27MzfYC8AVjmiFcCXCGWfdK+JFiAg4Ta0WURPl/tC3umqg9fPUEJhls
k9LUhKuUSiW/T3NSPwb7ZMLo296JZro17B8RVsw09JPCeWKttNBC0VqtE3GMHM6r
/d6of8dWtIhdqc3TR15/KRgVLS9UjHRx/fQUVaWUu4p86LZ2ylmUtx5AC8ZdbnJJ
v9fIZoFT/gUS/6/w6Sur2alGMBI53xq0JPCnQ+Luw9Oq/pmUTERKuwhHVNv6F0JQ
OCA2fdV4qInM7WnXewEczgPcN9SR0mepEy4UySb053hGtQlQz8D3k876o5jyNZVC
agwy88uHsHlNCXPqkH547HW06SQMYuKN2v21eGEXAOyro1HjXv4PEhgYErN16BQu
p7z0as1gYyG87w4BAs4x57rd2D3yVCJ9g586PDrvasYUyCjWQH1oHzF958GkyH1Z
UHY5gN1JsHxftc0rJULLG3xxXRKRf9Shzo8+a+/DISoan5R6eFjgvzNltqiEVKsC
l3RWX1ZfxRBDumSs1qxyTJ1q5GXFSBiNHEXags0+QST8GBiJvrX+iEsbSiAgQTXC
569G6NjOA+LTNRlcsktRNYcultswFRQHubidpB3PkHDgvhL9idreUVErkBjcaQAC
S7M461a0fUebbFrE8fY2KrpPJxN0Qo8wQelrd6ChcM582t3ipLhz5cRtQS8BDZGi
KVgijAB6aTbsW9B95wS4A9z7EB21Dq2x3UkR1I3iryo33RzTxi2x+eywpY50tOoF
/V3aDUm6NXENohrh03HDcLIjcVlDAIOdX/8dGBmOtxhcZ/xgD7fxeal/3LhcXtn4
KFisvSkck9MM19cgNDRIR3+I3HdWvPXPzg4IzPlLu/D3sZ1BLoUtPtzjjpUXSF/r
VB2U3pREYgd413rZoaWQkXk/f9zLwkq7ITt1ERFlCvsk/qpqFsUfU3oZd5jvp1zl
R5X6dq8Q7vdYloPZx4aSTHLbAL7ggNAoSK/pScC78NrMqn/7jN6TfD+agrdFrMLR
/LdmFcOJt1ikzwqoH+7eNYJujQG9wIngeyNnTr24BhWy0J3zQdQmoB7SSCylRMQo
o6dzKZ+IsW8OaDur69d7+zgpgH+EYp36K2b6X02tdCTbjcuyV6v0oQKRuxWMQGws
FqO7XKiwZ3LhMk2TTqUme3WLbDNs5SpvoVdgQ2QE2mB/i8OaR/33BCBbSCTlyHOT
H50iPboz2iA3MHd5bhaqTIA9LmxmqcRstnuU2dZdd1X0SyhUuNIAVXBZR5+gJopo
mC0UWMT/DrSzJajxsWIIxGH9OKLQyPMxn85GuGnzYGkXKAUADqbs/ebUdAkryJ0+
hxXstAgqvPRgk4vAlmZG3prZqSGgkgmreGo10yu3GaT5JncBuyESK8dTb84MzjVR
Z0wZI8ZZiPsNHc8BSC+gCsNBHq6LhIlAE5OcmEArzZdMybU+X+2K2MAcANplRHrF
7bLD5L4/uD3XsJBakZnHp0G1QmIPtiuoZ6xGp6VodJ77bw6cnkNoYwi4r5ekP+jQ
rmRifY+6zpb7mqt4RSwIbSQpEv3y6PUVW1a2dRiCLXHHfBNCo4wLo/sVcJhn8fFF
bfqM6jKvOg69t9nD2frwXLNUMJ1wpdL28PuMEnDZ2w+k4jNWLIKGfT0/kzoUgl5I
40lBvOMZ4L6jbCuD5GZJxH5tcUMY1JgqzmMGGiM5JgUFmWKPXNXhDgJiCIbkItXT
5dS9Fh/b0FLff1qHIcDFqasmWVvl+fvSV2b4z8+f21N6TXw8d0Nr9ZcN/88+WGVg
84DuOe+OETK2xIKcwkGeCHTVJAdK4VV+34um3YLJ2Kl9fBUS14CTJ1llSKzehWGZ
PgnIHxE5NH6U8YoBMXMDfgRdCsPm22meiNb9M6tasOYRwQLMw42TIAJ/fz9Mrgf/
D3hsFqHr81ATheEX/mbsqWsBKMgOKcLw1xU54cs4lam2hbuYin5DbvT6h/08IUd7
as/GpI4zUDzEFu7F5GuRenU6vSjeq8JxhJL4+SIVBsywUcJlKkMIdgh0z+DLRQ7K
QqCMD7GFrqk7kSGiYYcTolVD9VHnAEOi5qe0xZF2u/cJHkprWHjd6pAOLAwc0aRF
AGMDgqP5U8FWrX0FgN897ftxnl+mpX2Q0hrWGeATUisAGcKTwfY+FmsGwg2iTZsw
odRhLc59VRC8AuBiS6QwDWjt9zrFhsXJBxn0nujq+i1ekTZ34nc3i3n9YzakUSAp
Lov0fKd6U222rJdW0W2CPUgNgKjU38jLIblEGxw2ns2qiVsAg2lbkKxvWs2P8gm3
R4lnqDjrwZ4cN7BYbyUPMEPZZUsK5M/gROlSz0tCfqAu3WKzxCGBe159ACkxsc5O
9PTP5j2x70fGOqFTLJ0sJqXQaPMcg9w68uj6qmF6MHYnRe5mO2fLlz3Pm5QgNV6m
+3G4I9wMyLu5Pyw8sgy84BtSoweua/l/drv5m802k664jNp9rEFYKcIvehmS3fps
vP17+ICbHn/fQounjn2zDtiJESpJYj2PiWN3wm4EsRvenwNcIjSRG1cqhLnfRetJ
IC1+3x5md+A6sdvCNSPlW7I81znYH5TW9whbw//Emx5dUoBfEwN2PuoKDjDfuJS+
g0IJbLxbxgXgB3WU6VVzwFKXTzeIBGgqe12vF/XZSI2VVnGKzhW04g6pQV7GxY6y
3jZDpvlvQ3qfVQ9WrsWV1e3yL05O6wkt7/ZXhx/aDC1qDL97ZFymmm92JCVZ8Eg/
z9aD6u3VJzDEy3TO8dPKZ9g+b86FwHwovhd/1u/Fun5sgna04AQLC7iVQRMBaqgS
9ByyQmifn4pLxtBrGrjmGmh0QiGS71HQi2SLkZMt3phDmvOB6qYnRUeNuqDPDFz7
PAReEidV8EptjrCJdTCP9liJP3UZM0SgHG0/SkmJazipIa5aqFp7l+W0BSsBy+2m
quSJGrRInh/mkXmDDWKbZFXyAZKis3ha5lmFWCr/zalP3NH8kMSXcNZrcj40Awd3
7E87qFSPSL2y9pHd5mOhRyzdobM300ssBP+tumPB+8GA21r7QBLqOM0hwusWspuV
7Jxao0dWvLtjt29+Dy+JK7zrmnqC3f3EEyNorrgmvz6mzzEEW0EBCqqeWS6/LjNe
klRc5JEQjoHGVXbehhEOX8ZR8Kt8d7C2LbYNmNjEeXTdhSIkfscbtGoxIYXKawv3
iv8Pz7R68pyBuKAVh4+oQSudY7a9nt4UNPHy+E56YUFI3uxVcoxtaZffIUZ2dy5C
TtxAHRrzCrDhxaCE3NpkPFN7qRmp+x2uibW/A8QQYZvqgWFJ7OHFB8U5DUiC1qX2
BC0tPCfxQ9Oi7z+XTRBcHVcj+smQ6H0Vl8ww7ltHRy6t4h5Nuk+IzTZnjlhTaFw0
IcTvbQiTDv4m8PHDyYz76USDqk6SrzWVwIFcCmoLF130P62If9XKwkDvBiSS51Lg
RYMQeTEaBd7mnNJDPo1sAtfPhoGvsbwxsYyCMAYB/z29ctU2zFnY2kPL8iOBcG81
ntaaM9n4hIR1IHluaEobl//VuQVJUyDa1VMWwgIsUHRlo4nbbG50T3gNhnBYc9dr
5hoTPnpOode9X7sI7IfvTKIJL/8ZY1SU/0BLY8iEQaVjXWLXJLeKhYxsFpUI6bGB
GmUfhwqL93XSghgGoH0MjgOPeZ/PszKA+38ha25Fwps8a7g162pQKHHyI+hVAeWR
n0S82ab03WFiMJOO2hcSHaWCjiOGzJLiAfYUvVXi30eoINUPDVE7afDglcesx5q4
xfdwKLvK056IcOOamHp4aBNt/ozxrCYjSMwwqowLbtq6C4Eoi77lKnMlfj7dZ/ah
OPhvS8PxM1+s498M7KqKnjKkVrI5qki9fHRdHLWJHNgcI7cTU06nJ1uvzj3BVzzH
ilF85MC4HDsnMkDp1byNlEghh8dWq30DcQT3QcdLA4afK/LLhq3oPJnX19aFtZeH
PpZcnfuEIaQ1VRazVgYhFz5fMvh0+nAHr5nFAFqZaHIc/hDPv+I1QH0h9mbr6gEc
jpEC1V7Rq/Kz7zCEkfn03V7W+9tmjmeYGjQ/bcACG5yco69LoE78UOEbTt0F8j3x
p31Z8ibwbR62RMyu6cMqaIwafGv/4hySymvDG5LxagVOA0RtM0JUHLJSAzc3yTcQ
Di/z6ShHhnQgqXppPB2eSbC64PHGzpNkkrQgNF75mcQTy+VjAl3mxifGkWLGZ5O2
AkBB/F673DwSPfkYq3GHbxTkfUmqtLDYaWtJyM9/DtaTk9qNGN7Fn+odUy0BRc4j
PG78xT91BrFEYc7dfQsoGueEiRJipwpp8MzV4ll5Riu2XAuAKxQQP6cWaR+GodPB
z49O8/QWpxLoq7xqnIqNmehx0qmJCW25Enw9/EkewGc3yTFm8c7Or6g73X+GNMky
IAB1AFdvOf+QPRIi8d+tmwMLHGWlAuO4Z8JYyRDgki06dWRGaq/DTRtDp8HOkEwC
om2HERxvfWTUyjSWNtIJjhBwLhacjaKpMuxpt7M9PIh5gMEXvGas97os/0GDqWSm
q1KzOoIIHuYzJxX4GrLBLG0e++iYXWFBXD7DQ21Hl3z0PtuctHaWpzmtUap1RJlk
p7RStce78WNH/7jsd0dIgEYV5Mnh8+lNjPreghyFNsbd1xt+ZwXEN2F+1XW2sZWp
1Old0OiXBL8CBW5b4lhvOBko58MypcBuLPUpaCcz3WSdUqMNMRYmrbPkRek9SpqI
aOSe+Is0RrHCNgnYz4F0lEQnDe4aT7yt1CD4gb910UoQjKl6NryPYufbHiIZZo7a
ZORNcnZ1q0mBu77utltirHcpAIv+B8LP4A7vEcXkYozEW3iWuTEHA4uzt4S0QyUZ
SAb1tyDpTHWFdbMjK9dAKw42E15cqdncE/VlYre/EvlcyiD5ee+0T6XMg1eslhDM
smIIKB6X0zgAY5IdGpUxPP6u13KqI3ExTgtz8Qg4+mygydVDsMhpm+uphEOi/Re+
UYp9pqfl1Zra5z6s1kc8cycWfAi4LJnljuitiIyDmjqRcpZI69U26Jrv3de8hSSM
Lf4qRfCcye9x7KbsTG8V8F2uzdhlBrR4gST8y0eEd3myS/gMhylNXhROxUlWH1It
1+uU2IVaiMMqqwuWJ+xWbH1VuZ3RArhGDBR9HYWHHcL0UsaPKf658w236S3hkpIy
WGRI+UDOzYWfkvG0t13HhzzEgKD4EzyDrR7zVa2SAaj3uQ1fwRVGsohDRnhPsGe0
nisiD3j2rHxj73kcOnOwsjmDS//ttnWyoRr3guqSpOwiZHnlRf59TZoaNur+WzoC
EoIqAl3XTqd8g2iZ16bqATG3sTo8Ssfnz3cVZ800o22bAO7+yD0UI+3lrFuIQDnC
lbkL+mYnkeC2utinB/q5N+pAEsN0QJzUG8Hl/7/D0K8c59sh+RYeJr3wmldsHX33
NRDutE+o3Mw5HGOjI4jnjtN60EamH8DKAzsherlD18LFKNrDj+oVgPlANI0Fnnxf
hZGiiQxfu6AVYzZCI5j/V77tH7S7arNJMlVOJEb/FZ5GYS+UP5z1lSkPvMXU54SE
uzLrlQ/nclFVNVdnAelCzoLf6N71hyrJaLuhJ/9jUvI2CWC2Ar0QHbdM+jfSOSeV
cZE2SHos76qWOgOWXsAUjwxYYBYjBJcJ7LFBsSf75cawoCyiwenvyNkMgDctZH1F
aJEsAGg0bNiDMbzAwi2O9fo4Xhu7nFE65gG0SRGxVH5rnO+80k1dWojVJbAjaRR7
irP+z/6ZYnA6zE9nty0I52GSraqDxG2QOg9CKL6iZdusl138NJu8pl4xnHRpOFKO
Two4PafGIr0TtPB/0GMJguXPaaDz5WuL7EdzofIdNN3SX8dFdBqSevc6Kh6r1WUo
tDvvIoe6OPBZ0hlhxZzs091e6lSjUV941InsbiBinKYk6Rw+i7Hwh+k80ydgCFP/
y5oUlc8/I6UcnKc7RnzL8Mq0Kjj+cqZxgyDcGKgheV/qq9Z0GU4gfSfb/ZurIghP
uZES9BeijUZoqTUsqq74mwMuwZ4e5s07QIdgnpXECQwOZOCuHDBjtnccgUWg+681
K1uTKZzRkNx/kfu0CY6sANs2pgsnxkMU0JIA52h6BcB3PzAQCmxildkJ7iTjUHL0
n+iHR9zqSozcAbbVpRln8GOd3HHy/a6dJHjSu6u5eWYSCyKiowO416GXXMc9mGYQ
K46Du5KNHoZcncjj97mWR1zAmIYz3eTsftISKRlsQ82/9V1MwKjq6GzMTQHCls7k
0yU+7767tV1BH/3LKIKPd6X6hzMGFlO4X4J8+dpE5sIJxBCqAOBWRMgZYRV/XRPE
Ld26kXTRVDa1trkk4Z3EokTH5FiLEozMMJ4kH2m/8FfHpfJIADIPTQWcv8sjJOPh
pvYY7pc60fhwV0xS2tVw/7mQz8bmIAXPzRhPAj+nzHUOs3jZlGHj99l/ukvFvSGW
T9+QNuKhsDVtSiV6Qd8NZtYzZsCQU4I5698QZ6my4yQ4g7tsYPv3zCm9DtwbCUAu
CTT4U2CkpjrWo2dwwUdycEUKSrJVp9HSGR5/vlPhVJy0oQanokgK044Gw2xBJJt1
/h37ZcDf14PIbIAVEhEnMtk7xpwA4b0KUjYu8GQUUMV021DG2jefySnjr2RMjVs3
DZNljve696gr8NCr4re8jdlVYQwNSsm0Jnh2ifPPX5TN9Nz25fDbno6/+kaYuEC1
X2FqLkxVE2LjGnPVt8UO/VLubTOpKDXoByUSRl3Ylioo/r13IHQodjgUumzSx+S9
DUp0GT0wtNHxGzxUFqNrAobTDvgqG8MRS3LKnT+TcZVJPY/0eoAaOef6lSx59Laf
84E34+MVV5XZFY1OcXuJ1N4GpaC9xr5Or8JN60ku1GavXAeuSCMBRjWdwQcTmAeG
awItv4cMHsmZ1bjQF3f5gDLeR7Sg4y5oASbq5Yr39yMZOstiqgVUOYKHaSyLidkL
5Vjllts/D5II79dYX+pTVFOx0L39GtPmYri7JDH31nMQq9eBmWZImNHxRZOtE2wX
vYQZjFtWCcGLiCD4kKx+MB7Yv4qduxjOpSEhT0wpiFhTfTljm5nAa22pRToAEUCA
LK6FmtCuysI9A2S2xS/AT6zJGPMyKR9GS9b/i8sbTJthAral3A4uVB9PLP2R75/a
Qma5UZCCVSslpCyDpTSWoKv67m5kGedIo0H4wCc2EbmFlIx+cz63zcZBR4E9Gx4Q
4XI7LobGqTfbcaq3GplyJX2EvzfiGFSKV8SDuBLCsj+D23UTs4NnFmrKN5kgjRyf
hthW29uLdikyEVqwn/GcBKgNoiixQCBgGZ50GhwCcqSD+gf7y7w50CA0OAUJql+y
sy9HHKZ2kMy/cCOB6MbYxz0+eOxwFyzWuCrSvqeWgsK5B4T3M7Thtq/U+kJsU/du
Yx2dF8PA6DtbQLG5iGqcCtdlCUeGLMxZBHGsR6v4ZjApGbV168XU7C/TCHEH+Gk6
k0dMT8v2zeZ2SyXaZS53Tq4W9MWC3Jc9119en5FR0eJf+D8BNpQ20vAfLCP5aZjB
h3VXfqdbgF1XJi5hYj4AF8M4mJBm9wfhOOQVbZm7lCLpjxCwtxUYTzzuiA/4BdjT
dY8lYgti1yHIuJed3akY0Jg+9sAPfcEqspyFtirdKrAipU/NEedT5TQF/QmT8geI
r2D9kQVszomHv0bbN3kagJ92BEvGDn9HB48cJz0dot6E99KXLnz/tJUkxTOFA8c6
DcmgKQPDqI9sas8h6NLvzFoGUQkOlpMmEqgFtz926erPwxpApr9+bTjlhmNqT57o
RBKT10T+P//jrK3Nf4ZLNj04vNRZPydJFmh+dXxDDDoukpq2H/aPaqCMwJtZHXZP
X0woT/cIaEp+vM6Vvba4O/qYiag+ZD/0Vw1526YlfN8JLIsunwjVnzbBD/B+/wb8
vAEnsxXAIppgIxnlGv97QwwwuAiopsRC+3txFZ//ZAGTqk4tCEAF9bkFx6VPhiGX
rdUBcFrsw9Bmww3sRF4wqpd35t1pbOtuMSS77Y0PRAaC21ZLYjG+RXr0kqYa/sNq
Z5rhC8eg97avM37JfsdkHHD7tqMO3jRv/XqrxqAuK67V7sdwGYBgUkHgy+mIitbR
2YSU8J6RetB+dO9EKH9/GPoTfgoC90NbdFn3mw3IZAr8e/E+qWf6yrYHYz9GW5oK
+vWZzVG3wFloABHvhCDotgTUc6ZihOgicKNpQ3Fw9SCFaT1NetF8ssjiDfAPEDv4
vnp7vFOVrLmj/oCYLWU2MfiXcAFJ5IJoJ7ag52IaKI8LyldBXuuEPIpmlXBMsh/Z
mdNvPFCPCpLlUdPiqvX3uyi0U3eIBMzFAfnE9JKlxdy9i3nsdETUQdGAjFdd1fpr
R2Q32FK/Rut0/ouuqRIFLHCORcdVABRSI/v+ZRrzoInv3Bpf/qg9ZcMbY6Wb6Emc
hBS5Qgbs2PEi+uTCs5iJ6CImKqPsjjiAKftMJ0Flgof3/PT/i1lihs/C24Yb2UOW
6yYKPxJ8MiNBIT3L1vLdzdyEheIOHBYY8cnxk7cHrMvv+lkJTRP7+ZpbhxH5XqN5
JaV0SkjmzV2DKsRns1fELABhB4UHc9geHe5KWajSt1GOtz+8S9sZ00svXu7GnKPm
TGRQi7cA+xhSvcJ0XlCxAc845ClFr22quPZQLyo2+pVdjHK2Ze5Igpd9wCBejVMv
5dPSPkK0ju4rvK4Qa8r5kn65AlMeGRIQ0hHVM5jGC0T/P3aVJmgJBu1szNs2QeSA
I0ggSPr6my8RuZmOpFiLfZxB/dNmFpTsXtg4D/mulWFaI3HN0ku1Bc/P5MRX7ENd
0/IQMY+MAOEZmyaTDcMtv9sevEF2snzq5hO8VY1j9/nF+Crz6QKhUQccTPI8D7Gx
JgnB8h5HXuMIEPoVwDkLDhGHIc+6xJNt566SK0QDQ/uVxLafJsOXByzA54Mf8nDO
WavRuWtHiMq3oouqRL01tqYqc7GwilXlbaQDwh5gMN9q3hFnRMkZAHRd1AV793jD
ouWZs5fWTGcSO4ya/RQ/vIDjJOFHvX2zyXuRYSYB4BvxLEpe0jCZZ8AnGte6xfPV
SH4QaGZqzW/6RSeCq11wblJj7QP+PFY9zdje9cZPgKLzJeAWgbwJU40uHdjhEKHx
zx6bfd1b2dOCrxYukzfUMj6v18fmnmggKbTkatI6HkdMvXgCzHCuYnKjodm6K6JU
kzrHvzLIChL4QSK1aV3WPEFL5Bz56hy7AQ7OkW3lhmsfaOxlL2rUGHcAy1juX3sp
xRdcuXaZwaXsllHadqv/8BKwg915JzhBtYoasHcYSiaiY0lsH26PgVecd7oG6+wW
/Noi2F/88vW8PYg2MBdCTwzfRzaCKIOFTZCRzL4qfhMsGGIJ2qewVgAiRyArVihw
GAZ2uFLTdH5KW1sAKFAvteULoD20OXJMtwc19O1PkQYNvU8/EVuiWGqFqFkavE1o
6tKpqx5hMf3jL2dUYyVkafQM3p+pke769VC+iIB/OoVskFaDCS+S5fosH1hql3SV
hMtQCqtvNOIIlTXLR+wM+/X0lVt6zW9pFuGYoQ3ViPGZa1DDP3aUbv80e/BgVr/+
mi67T9/4Kmn9CX4gX713I2ZS12DCJ7oRfJxPp43TVUsa/RNA18+ZZayWsPEdtwPz
LxXAArMWw3xSQvJ4YqHiFG8tRgNP2jm+2XQA8CrF8Nmd+v0i2ZitGfDQXKg+Rkl3
GODHt2BWamlJo6RhWV+Rg6XGscSXxjVRkSm734V9GkaiGMSt2XU7d7hdO/VWOe36
dyKZCZ4e6Hp27yZ7h5BdlYW/BDjluvKCmUFQf6YuKjO3zHEsYvZHV/ZK7OviFvt8
6xj617OWiQCdRBUVs7rKLsqm7D+pYbedPrLjwYw8ByhbWmEoDmXh5tBF5FEj2EFc
bT9fSkGkFUJj5PlS2AnnTqgWJsy+4s87cttRLG1zbto5hgizFEThb+O9mngMr7Gk
XYSvv7oM6OT85ICLXADze6+rAwyistx9vx+Fm4CehviIqZ2fMVZu/CmnSWl6QyTT
2/Gtxk/GvO0qrQfYGKmhM2JzViLTTyU91F1MPVmFegcJmRle8MfnPN/p83uMwKws
0SQnT09pKfLEABDRw+vMiw/9hlNrWDqV6WpMjQpVhsQgNChIM0ISNE/HkBPtEhcp
9v0psM6OoXcTaR5msUgLKXuufOtpD0hDW93oTZON67usYL4Xh5x1qzegZHrC6/KN
7+gR7RfS/9uWGdqz7VlCtMR/fK0oZ4Gy2LB2WdBC55V1/87gXHXRAkYakJsOwAWF
U6pK4C73czTWxL/XVWBDXVcuTPaQo5KqrwxKRNoCIzIAepA6QrekZZegVRY5rkAo
p/RalC5iDzoY6iAyyXEvCv1TK2XbfiEcCIBdYNTm5z2heIitFmOZxga18E1rQbay
3GU32Nm1uuNd4iDkimUJN0ALP5RpYswWGSnCfDxSIwvYjUUiaQ7oapmfNhYf2zTc
53YaGl8rYpnuhtdU6RN7gGAQ+eZBYFS5xzu3skyc5oqJfOigVNeCYUs07hxEoYvD
EitfYQz3gH9uc0+vfNMPWZTyKINQZomoMWrHJB/50G9WymWsc6RQXyOxxs46/61y
0xg4czNPJ50Sjz4/XjOHBdlYD32n5FOAGUQZqIeQqB8iJ5GE7HI4cYk/0/lSHxA6
Nqb3HzrrTTp26/4FSfMmBpHg78eQL0kFfTgdobPoaP6Ml2h8mZjn/OEvr2hV7cER
d18/rdpPgbb6oaNRHG5yFeJllYLGm1ZAap5p0PWBgoZ0jHBS+sjI/vGXY/usjKB4
YRIyLDXxRB33ybs05sXDOivg+vcSTEqOz7LNKn/Dm9+GDyDCLZ6kHkpgPwckk02A
isKnkmgrGmsg19d+REmtZfTHhxVTUj3+IztkvZ5jD/TZlJe4MgsEBgdwS1FoXADQ
ckpwOXHBgd3qMPmnbNzKeo9QyMNodMmKAjCcSvvmQ332WiL5FicQBw/NmHzo4lop
bwJeXtf1LiMRLHZ1ijh33iR2hpr0jR1GqSE48UcDJ7kfzhFrkisvM4nC4QGPZhf3
SfHeEv81ePQy2N0+h5XJDPB6a+qNf5xzKWPQ/JUaXEyZ9URP71DqEotggdK6Nsa5
S7Zs/AzWYNBrv2PRblbq7gj7cpTtcGrTvKcxESRQ7EHjxjW53oXZDEtQ3+MJoWrV
BgrE40gupXp3BE1kgC4OnLF1a1I6XjLaJMY51B7EjLNQvGWC0aGsni9XfMI7YooA
Va9xGeWU3DzNw1xTgTS6j19pBw1LWWZBTscO9gd94yi4uU5b23MV24XhmVISDHiA
IJifsEv+e7GsAjd+daEdk8h89ytEdYtFKkusGb6PYy0WMh0COi1Nqt68bfz0Gt4B
RkjaoFdiub6QJ/F4LtMXdsTIj9XcO1+sV1Jv0/ChEOeqGEih05B7tOkpKp2hQCHF
bD0jjZn2maez9vx+sRVW5Xd1saKGYVYe3w/K0+zMiNtkHyMZhYKmBKPb+fGLdWpl
VWQYvEZA6+ItcmFHliBDuS3IgocCXehHwbK86jRS0aiMojPRuevHl55iwue6OcRj
SjGVLeyrNNZbeeYbWBt5l3KC0sducfa5V/OnAmBrEsnzLtvfCCuZx4KNat2O3OlE
lU8MhYQJPwqiDX5ZO2TzDKy5I5N51Ul+7QCTOoWSbzncxP5AuBNSSChCwVaGPAsW
Q/9hn9+6ATLeW3CqA+bKTV/me2trytSarYvPsPnVEkL1r8D1VsGDjrGqK+kynKAk
DBbZ/L3tWkT5hBIYXindK3uDsW2e6S9T/qY+hGQzSaK6zPowwJaKY4IxD7DUIG7S
o+DuctgI5EriEFQgqdnAiMg7Dw5SazztfBUAtfjMLO44f2VL2HAAGrr/NgjVTkbh
yVR1M+/8MwkyYApoavkcluy2+V2C4RhPEO3TtQ4MpChGLQ7e2MMIrwSl9P/7WpXJ
b7EI/Q8Ch+tuisaiVws+5jxSJNXw19Sh94deKBUTEKdIq2Jpvam1HgvjEjXEWpQ9
YxLYYehQWBMV0iu9R5xS2sX9wXGYAYY0TCLNXhD7gkReoruZKakOzIGWFIq4nXbV
C/WHH63f7nWwSCjxb8/OxFNKbWcWqu9kdmzbuA9pvFcDpxpk87Xamn1KpgQLvaGT
R60nRMPjR9pLhEfu8GzsteByn61YxaFvBgGr+1fSTST9ONHbjjUImZh/gGgvonbM
acJ3pR7EedOyYqb4/yQ6K3X7I99LRLZXDXLtdO53SGcSaoHqhhwhyqkXPOK8Y/7c
JNDYUgW58JMfHzRKsZOW9nbKBkJArWCsjOFuBbW7rkx/ICD5ZOgKAp5fI5rph5uZ
FbMzAC7jcDrDSrDOvPVz8bWW2sb/JJCdlEPI4f/EPQHMi1CXp4q2ITMXCvpIgVxT
oITHIwrRwIJc9ofeIWJuycYUsjRoBEAr1Sj5VO5qEA0ZEg66omck727AmdUdFzST
lIkwEpo/EIgf53CudjHq9d9Rdwn48a1wJt0fbkdJTas4Q47x6w28LHH0mwDopMcz
s0p+Td+F3AjfiD0xnGv1YY7uiSmQ+SwsMLEaFP5Q6/DHCV2nbyFBC14Q179gyKlD
CSK1PlbEutqjVs7EozV70S7rHoh1eB1yPmE7b4SERZmjU6U7/MGO7OUcCB6TLSww
2XqRI0yHLk7GisL3mmGR/6q3TJir/vvTy/Gq4EOD0nolEH3iL0a11qtm8l2A/Mwl
xLpIMy2AI+jadJbjUQcvHgOfI+ieG8nGbitPTJL6PvowFtqehWy++VVI7E8n3amw
fcSRk5SgOi79ByrUZyBuEn9PYhj60K/CqcoQvkM7aKRqZn/HLEQu+2c0soo8uhil
HQln+QtubTvvxJQZdckl9UhwelHFLff6M0P/Mzo3sW5rF45wEVLqnVJJS06OykHt
fRE3ukwy+D7Hki51OgBRDnFw+thhcAUZXwAKX+qiZc79h7uEmSCuHk7kr//V/YkD
Q+1tvnt+7SW749TM2NihspiAmO2yw5/rjRfDBkNLMvvhtqqZGEvpzrWwaQMR+Eao
qIjiMoyx2vexHM9OlngQnWZCvXlMFmI01cBdOLs+AcwZrHOA4A02Ihw1gyku6j4P
XWdVBFDGDBNYFMF852Q8fq9OJxDTmgNlT/MepkHNb4J3ypOsx6Eot084DKVUl1NI
b2r14N6NNI9XAEmq7wpaiRCGSz9LV31s6k0IeGFg0P1Qee+GnGyJKjbeaWOWP8UP
wQABGvyevhOHORoXiKMq5CzSLV89ZceM8TVOTDTlg1f2rsYUtQrM1Hf8T9WMdIrd
3yerKX/3X7SlBiGsPPZb0eymNz8iFR9R3NZC5OiTZj8JJxVz92f6PWtmbdIsArHE
qRBf0ovh7eQ7XLsF0MnKqc8cG+bP9S+JMrw1YNYdLDBh30kwQUEQn/2o6DkSn6gy
tnJILWpecsWr4/V3HXbWAJgh4/HRzqwsvE6a3vJ3spnbFL0ZXEm7VsIak9iD27c2
bLd3jvzHbTFtp38+yThHUn9IiAWtwBlfZlycvMuaQFgsa0pSnd6b7s6hstwMV2Ey
8CZmVCdBiNYnptzaD6nEwDzTikCJIHeJlqI0WE8/2avUjzwubYvcj9SWrWPHvtXh
uWaNNmCnkCI42yfp1xUMEKjtDHcIowBxIDFC23L2w4kRQ/mAFaz09mVsSurZlzt7
xfNvod7CVgMvOdAGoUA8b4dFo+LA0z9G6UEKX5daWG3D6XfGzJZZVA6KZVHGRjOd
zAGj853yJnDgHF+uc1tZvd3aMQzG1RHq0J1qm5pBbLPXuBtesWRuyTUJ4VKu6PI8
x54t2JVDdBsELUmKu1qBNRVslKW6KUV580D4AIpz9M1/HBm3tTY+koJosaJhWjwz
T0A23heHBvijOUrX4M6at/YFi2J/D+tw2PNzyFzW+cQyVOXXGY98UprdbV4D1yLG
fGyVW5V4c7Oog7UUETJR7ap8lX5/Dqaqz90907fg6oFW72FEvr7B2bBXsCxeYyPq
or1BJqwIZJvnmTEgLbxuOIX1Lpscs1M3pkCZdCZnACTinvE7rs1gJK7LmQPKdqGX
CulcngolsxEoJIVbaapdQhgZXyRN80dZ8h81L/YxkCkM61FrUfzHkI5it1bQ/UVz
rolizZVpE/g3SdQveLhWP6LBM32cSzz1oclqCmUikSOGPlySe/l0NpNaOk3vRAK4
7DKZ1hToNaYUwdHIMKOIqRzLLCnv0JWqRHZA7ScpWnlM6iaZQHRBFef15FFB0DpZ
W+cKbsNMnLWlM0Wt2J35Ibe4EFCNGkgrQjuy7oWgqp252Asw+adqZb8baqsg3Km+
Zxmx+iyox8Hk8P9bP/fUQ/k5+m/vw84vni/01LEgSoSJ61IdA+MBmp89w95dHUHL
Qa3s12d9M+CUPHKH8s0yW8zIC7dN9nPAKN6mjVtPG7w0pirzOXi890fNndQAhU0X
Bmc2nNEdqKgMWL1hOaIw9t21yMjEMI28YKRLXLAJkUWpvjPR3kwn4Vj3W7Z0h5eJ
qA8V1GgmuOZQnaQB0EnePRHKqC9JONI5UTB/oGnwurDG4S//vMWCY/ANc3kJcpf5
BDgPJg2ZMDE1BBbh8YFMK7oLV71wUtWFjOclJmF2r1DIME7+ZcOSjgznK79TEkUP
3kXqe4j4vvk4nItxDIFNRhndkx3SG9dCZx27jIe2NkgDa80+o/MnlpRCia56tFGe
ZWjNgdfG/u+wuz2QSn18wqC5YEG5Zx6bTMtT2p3te6At65uI1bezQo6lhGciQEX0
Y1JZbQwXs8I7S3AXF3a0CTiex1pNgGe1dI8PJe92vH8yymCFJzvHk7TZcKghwUkq
RpoBXOb2xd1MO+jrIoSzY9BJ2Hr5iKD77dcNetQZGP3dasBzhtRA6EKoK9BXDznJ
KTxc3FuWQE5gpbqilszKUetElSRNmCsJtUJLUZlfjoxfgexNWmcUquMAA+xzSo8+
vVxDswAzPJbHRoHy/AksTrjVz/vI+wtxowAIDH2EQ4hwc+AwhHZjNzOe3SZ5yLbL
dqyTEMI+qB/3sdtz60ujt6BDU6753V4oXCsC/6tQh13MllyilJDRc70AvcOE95sS
4l1hNx7ABtllh2RdmXZ1AJbQM19s9TFnaHApyZRrBysLZYh8H/JGwakB6sUUGXDo
xLYYrQrvrkWSvdVWDx5br8FeQG3XxPqPa7YtcnAtOE1TJoxaEJm5IB2bTpkwC2Ht
LP/xuNcYaJkR9AiMmu1yHWC9kd8H0aZlpUwbC11J4EI+sCWADl9Gq6YG3/1iLkpW
DXTbViQ8VjUejiUtLJNqobHQOwYu8FdaIOre9Ub7ceE40sfP6kRo0ca58jJ+v2YZ
ky4peuOCwWh4DhlAWVIgPIiCbJ5LfRenKgrLB+B5eeg5nQGfW0CZ67edwl1XD3iN
xuQni+Ixas9hfw/S/xOGcnz62S72OsoGkcHZl5knPQQdYseZOplP7xXfP3EqF/Ee
lZhZHqw4umHZHK//TGBfbdvaNsupSfvqnh+5tDi5e8M/QcCQT1qq6RuGGKVSkt71
ECKYa7lkzbBFoXOy1NsX/pzJgFs7j4l/SQTtDKhZSXYRFyctu/JQn5nUkaoe9i6f
/GaF2eApcQ7lgtZ+KZE4qCeiZhR0wphay9zjO7iMu8kDIZYxP2Fmeixb4B0DFPjx
g3QJwzihGnRfGkS9Cv61mhe05KRrTEwTdhWtGPDPj4bI/bo+Qw2QjVSHviHo5vfc
Snc85RkJ1I4DuboIuRPce6dt2CWgJNcYBBZHxedHPB9N6TAOkEZ0citGrW9q2gSG
/sZyEIEKCNFXTyLIdd5Ef5n5iOYPadLjuWvMGlI++66/z/9J3VDkmjQlXaM+9JXD
qcz9FSIx1Nqv5g5fcLICAn8NOYusfbrgD+6oy1T0Y0/GL+ImQd2SocACTSkeep6C
Ml6JB6QNXkX9kAQbE0ad1rhxcU6sOm8yp8JN9hs8gh5Hu5YpNyHFYrtFH44ZlPav
23F6dJn16ryTS+CuY7Dd6mWtVSLgHrMh9r2QH2tw6ZeuhUdeNdC1rFQVf/T3cm/w
4MYEePH8oVIqHTNd2qlQDveJ7Jrn8y4XGfu+HCbSeEgUz2WXsiejyPAcvf568IWI
MXiCZnNxD56EnjKm2/NI50rIA2Mb9qVALTunu691OQXNHmOKgMMYyQcn/DwMvfbj
PwHjNMcqczpqhI10P1KI+TBtHTJjcZCSLCQhSR5dgqikp4Yd99mQVvVBh0kBfG3X
/+bmXLFTantLWYRnCEcI+KUhtIXP6DW0626tnZ2ZL/MSRpiLag9buYRfgqVZfaJu
ZkMu6xt9Lfimqu3E3wVCmiF6IMp2f827O4mdOcknx1k55NtpxF2Wl+YqmGYjdc5/
dFGJ+bErOyYYdk2045Vlu1mg39naxUf3MIRV6RXoDSax1nG+htqylb6oAVICSYNO
h/ET1FKsNE2EJ/b0qa3a0DKQBxAwu4MqpcKZfwz8ZuCdgBcjbYnCk7JrUhCTvFY0
2WhMfJAT2XocongP+lkA7tZjxLJfEnbWww+Zr2rF+9uxOIrm1eXjvPhRrGKHRPe1
5jdTOd3Wa/HdHOWhhGW1qj8artTFVKkkQC6EmA6GJCJTXuyvAA1vkUW7knnw/PlG
hvREbkLCnkSwqzzBQpBaufmmLTr9aqOnbug12OKV/6XnU66WivUDwrQulqvrhB33
hcMROk9htFqB2yP/sz1sGkQodOIJOMr0d7gvdc9q/cgpKunINtZ9ZRV4z/YCDIZS
nU+OR3E7azdvHEyeKWIWSwURFLH8+5fvFgTrRhWNRZ8B17Ch+RNgf6bDDba1ZBn4
8NPIeZBy3jju6pheAIKmpndEcXKMVZYGos9Tb/ykrb+qfHKKXSvSYTqhClpCVfYH
dj5fktKRxUJT1/VAEpu3sM/zCRBsMVz73QV5MGcMV1KXEKpb7rfSU3BrcpI7/Tde
gZSCx/JRRYerImW9efQ+ksiV7PdmrUBChAkExnJXhg5AZ4ijwkyo7VSWP7MbcPKB
0Ld0kzxJu0Guqnb+Bam+ZG377wqEwC+x3miXo6BxbeTqNR7ZNLJvnzmE4AooSr6a
gvpck0HeDiZ5/4F2QK7EDKlO70DL3mF6h+B1yRGXjfPH4/rH4yHDTZEDRp3XKrw3
f/zBX9EwemtlYndDanQopWrPwzhI/N/FNdsn5cg98MYeAPNTHds0DeXhUQ1rVaLo
MTqbFZ3BSGElDXgFy9nZPao3A+0mS/3lXecQGk7MgqqSQznq9B1UiY45L4dBIid7
NMLhSyvv5P6YMiQejijKUPKDQSweDUK1XyYIrRNcO0r0FQdYZaS4Wsu62yz2oAXL
KCj1yMKcmBwmupuvsLlcIH7tftVYvAhkZKJi9iz8Z0nFOEElGlkaGnhe2csEOkEk
dRe/hsW6TNpDTGKCNmvYE/j09M6xqmhJah/S7QVnIWXLp0habBODTlwTBApnfAUo
PxiD4/TtgAkwI+DsHeGR6Tn4riwqPXoTr6TIkNgo523QeEkaFcHa6gPyU8NcMGIK
Iuzsyi1b+ylC/xTahuz4KfiZ6ru9SKoh3pkr25K+zWm6XXd24H3ayGa5bKsCeJ/A
wBdw9Ouu9643HdWv7r4iuDALJUVlf2WS0nXeFLAau3dn/y+p3CIC2Xcd800HNG9r
Z3KMBUuLS3E+3of0Uf3ted/oSj4MFstR39e2a3BKtyqKzyLjiXaw2NtxBHh97oJ8
iVqM7lw/eht3DKlndRdBwqGXOAkSTGu4Ww2PbXhmGxXF/sXOZiDMcLUDgd1KHtqL
2lKyo9EY0/tZIh2lPcHI+zkAkdTq0Tm3v5wlXy8xNM3XQALBbtB1tpWBoBgv/cVr
ElpUs9146mCp/Uhmg6XVK9y6jy4VtgAhY4VxhRxO/S+wz4g3xNlBPXvZy3JAxhus
cgMolp+qtYuvaeUpRQsXqqp9PQPgkFholLPE5yMOenYvvblSTS7Prncf1IA/gw5O
PGBroxfBI4IJ2Ee7QUakJz+7zEsMka45ixO7ArFAbxk36fPVyqazbGKQ42folOCU
riR2A+bZhxBNrFtSqXK+OJx6g/PmzqJael4yIB5bipBdKDYlPNqhi4b2GgTt5fFp
hxPukutD7Fjq3FP1VNuA8H4iPWdUwrVvI/tXIS7AyTXsI6dpXVZSTzpNc259W9k/
3gQV+OkjId0N/iHh8VNS6LSBcmsWh8yBVtrVKaSVwTerjV1C7UV3ThTj6YumLnM/
K8WPteI8MA+Mtv5qAmqSaQAufU1BdLa1go7Ohc4YB5SssUvla2np5aGERdMN/PdA
fYaZLL0MvUK+i1rz8nGCQFFACpz+4dbrcBYNmwp4Q9VLXQiXPSaebvX0QlxBdg0F
iBamPuFB5DTob8EV4/nZviBGw86W0OAZVLdv0bXzP77P4JRW8Y5QY9kgMVCt+Kwf
Swu/j1taBjL9fcDi9feD7t0l9SctgKU8+zyh9odAcVHk/9k0rfu6F5OE14GMU63p
vW3UiNCLYpCfoIiy2lsdiWlgzCcO28cjpubeHb4VSFMdUq7zMgdkuUOyx4TE74zT
pRe/RyjwVqoVeFuB3Y6sUuaT926+I9t4mwyDXhEcuZFPwuCdO7BONB13A6O5l5d6
t3OhKjV1QQ2Ba0iZLIMIySi/Ux5DvH1D5sVbUKM0HX/RZtuEfv8GMP4gjuL+c8b4
EHZW1/V0+BFc9JK2jrjq8ly9XoqkQz8U3sSTpMrUV8yEzfGzJ8r7llX52BCO0Hss
67+VVTslrdMNu3LaEkWwQslgIm/GEOJf/Uf837u5RZ9diPfWnTsKvZhu1wa58yzJ
WLbRpKnSJKieDWBXJi8TKHAghAwmOaw94xloHczw1r59I7kopGpU/t1E9rriPqdD
VL8Xn7m9+YX/O56SLHBlc+ojEj16UW2rA7VIqz4PqZmXn3wpSfBKaohTIvp3KZoM
Deb68qjp1YfElRRVAP++u0SfcR4UTFPJQaYrGBEKNWB9USCy+E6rlG11V+fM63yx
fm/dffmBZVPRCnSNyhDSuoeYYC0uGLfnvzGiPY1iujfIC99Wu5r1RqKyk/sAiSkH
QBreB6zUCd2xK54DVmVKCP3TXio/GtFIs2GnETMrtbi/iKF/WlEt3pAAN2H4c6uu
DRSjztNAF7p5Ls5qO7mOdS7koID+FX2yhuajRcl9RrTitkDgsJSUnAEKAx7iTVpm
JeHmEqJekTSNeJ5mEOOIy1pQp2SM/DGhPfzJWmZe7x+pXeyFB8ghChE3lqyMpI6u
1eFqEePjrtaVcyXg5Mz0kKRSSZELuMzGR15Ai/t6mQy4pmVE3dXjqORVmmVnqzhG
vZn7K+mXQhIdd7d1TZuiWwhj4gmrsdSKQPRSw51HdKnU90HDwp5GmPRqv5ujn7VC
TiARqNDM6kQzHBg+jupJnhCAqiKq6sKOD7x9CYErFb1HczsCS13jmNFYnfmzw/+0
9bYCUYwAf0HoPU2BrSXFvl7HYwwvx8d2GKYOm9sCHKKFoEpucfu3hrf/S2gu5M3h
5CLgsEiSHTLm3hUUkjVpSl5QasTqMA84hd59Rs/lYb5Q5mXr+LpQG+W08vEazCW5
Ql9Dbu7BZHnvgrPAPAiaCAFDs022yqYcr+/l8L0FtQzuBG+Np72YTAhkFq57nwlj
ZtFLuqbZnO/dFvOc7MOgoh49CUOc2FzWj3YaIj+XYsojo3LjBQtH5j1OH41rkCTq
Ya8vD9Q8GEME+RkYbz+xkxuXWu6VY3ZbsAKdyhOGrGx+34Aa5ImgiPCJg1E0KupK
CHGxbo4VWXdXjHWESUWPWzo3+3ligvVHi1t9aR/xxJ9njwJiNUkbFqx7s1sJCznU
+Uf7Yuj1ax20Wq3QU6tyL2CkJAv0mZ6mLubyW6xWx2Y7aQjdOeJYIp44xlqGqgEb
EtrTApCpWgtvRAVoLQLQ8kAOOALW+dRi4n94baxpnpgW4dqbpbhYhJPc8nxvg8gK
nvrTI1rPSRSu5/ukaGLJUOrhQdOVuNNcFJq9ujQ+gdMbnAhVhOugAHd2ot35QfYu
7NflosRsJknTyqKC9AWEkjGvj3jA1EMS7ED0HOiYKneAZJ8eSbfJYojYLVuOA1rH
//nSmaFZXaBKexGVlj3DpAR5yY4Y4XYpIZDwsGn7VaMYPLEXi3meBfGVK7nCAiI0
v3uhBkhv4jo/qebgmaryoo+FuwgR1vVqWmLLchmIgjlzksjC4ESdyb1dT0w9VHb6
vxCvpyOqwkWsRJWROAuLNwmRi1K4pxPirxGiSr18TWurqtkZPuAyT08DI69Co+GV
W6IoTjRNySqAvJSYyIC/9y06aEVx5UEOe/TMR4w2Lcgh9YbYDrk12JK+Syrkck8+
3wJiOPk+nhNMzkjlhoW4x/zRhAoXbjf3W2c4Vw+0kDE0r05VDY+afrW5sOtxnEE3
C1mlFlupeHmX5yrXiySSKz9FPocHACmTE6mEOpUw9mDWXgebN5Q1HlDoR+jbvwWY
YyhwygTwqvjxR2Orxw3uaC1ZL4ljQ/n6axwYtage3+zHH5WuFqgh9rceCt1JoNKQ
tzK/aGwyoKxPRPJeHWWxAH01anQlu+Rfb2QXXmz8VgT3Loh2o2DRAbLrbxvle/Mm
CTyp1oiVYF7jMesLzALqM2MyBYEIbaNZA/XFp8JvmnEqkwQ5Sg9cwen5QSJUNM0U
TeaVPXY6XcfTbgLg7u3ao7F9zThJEfCev38YrKrTjwJUSW9rrevuHEOGLdSFOOF7
vWe9nCzT6aEZJxpBBuATgmFVk9uHrR5VrnlVSaikE/jrRnbb0HLxAnxUyxzrPsdr
Svd1zdudYmsOZwWESeYIZ0LUgWbnBwfarpzli2X0b0oPNSySqTi/k4bYVuYCGBmg
nYE5M6cgUO6au4yrtyqjY+/XWLxql8hF2QmoAyfO7YYpTX8azRlev2HcFkoVPnoH
9Z3cMZ21OQI5KP4a2d4Z00NbJeessAMP6WNpSPOX6vtErrVsCa8fQ6YtvTwLgBgB
kK2PZVTXtUDwJD7fn4XpeduhqkwERo6n20mZToQT3u+QIUWovWcKBcEePUfAwK7o
kWHnKaP93yFpuaK/bGxD/GfhSbYDUFUdCB/8wweW7Gy853gQpq6EdELeQCpAfFw8
dsliZojial7Oy77PI+PspCYQFBdgs4k3ineciRaAJo4yoPQ0bkkl93qslqoDpVwT
tayvwDEc7lk5xE7tlzreQgw1Go8Ic+SNN62NIDrh4G6dCd7ptIttR6MTLKqx87It
PPrEUTczgBOafEnd39lZzNSOLVfQ9ITlhtUoXq+vCDmuzkTziezKrKPo9k8K5Je9
2hNpCcfyYJx5hxu0B5zEcdIL+JzyHaiV2lMcL5n+Qo6ugqDiUfilABBiv+NUUwzs
Nvef37HbCcjMFUxAEU6itgBcuV55qnvUIDFpLcdbrJMHIDhh7wZ4I80Cuh1/HMDL
wc0QcpqukzjTqks+v6WBPA+Yqy2dw9m0OOoyAFPCSAGHOuMBKiMmZVpekE7We17/
eNkAb+Wf95kAZ6eeQZISIsbJkwvR/Sr5ffnlTeWa6+OOhaZ36xX4gz/fGUB+XtKL
reM6cgWeLQNQB8kitKmugqm0Jv1a53EoUKxI1rsMO9cxysekN3Ya4bwG8M57irPk
FL3HdtmHY2+P/yqsLLdfWcs6iDNh8woUL6TflNVgXvHDePBI/CCgsdEE2zi2u9j5
YHRQ3kHhB3Nghblj1xL5RYa19YnetarztciFAy6/KQbiHTrJ1GYkt+ZNPLlyiYkf
xy+8XGg+c3zcuqwuKqYGB05zuNfShVUqc8pngVITvjQPgxl7sX4pMr+bAsoIE2lZ
19DEHA8VEjR6gWrH8iNnuSVzQ/w4hB6PSThcjq4lXq0uOHAqqIuweYbtrecmWRFi
T6feK3E1Ph3iD1LGvGQFbEg+4cyN1eeVfrnYuUZbJ740VQYpBdBnICf+S5pIJUoP
PdrrEfguwG9H+whusjeZcD3A4fefaRz2kCW3xzk0qgL5xQZvpqdmuNPAzsOdTFLj
VUF+v7TAmEO6x5fy7SDZ6OyxXmHMX7cLKRI38icM4DivtPhtnP7oirdpw3lEFfo/
jBP3k3+J9eQEIIq+vQNhfpoqOgCqb6NKdZ9Rp18LdQe9taO32WseJU3V2mHWhl2o
1cAIIRi8xnBRZyUdjlEC2Fn+HmmbqgjgcHpoPFwY00YfoP69SiTTY9klKuS4+Z1/
SK4C0YmmDH72khyizb3BZT9+unowWisGH8iSIw7d5qcNzZ31BXEczoZtk6CZOeM5
0j6dWZ27k5FB+9sToXKEzxfybvwg9+y8+uPHkMgBFr4pJY0anOCMwYhLT5sjnGeN
yBa9eha+oXE5iPxMVZx6MhEwQYBzNOBKoftLmJBfr4uuELgV8RT427Kc8E1QoWCi
NIj3kFtqILAhCJwC026fRqA2pVzzGU5WhS1eBHae60F0KXMFCs3JzjIgrbeNWRth
Ba9MuloCLaqkLc2OyBBP4H9BksE6rObSZ+XNxOBQX607yXUvmuZfRwZAJ6LtDu6K
cBhUEKCodr6HNZbjK3+2uu09r5GCpKJ2PDNuVj75c3Ro3Bp6qTGd//ONcakCQ9CG
S4SI+wYzPdpYt7cjjSxDZnDZhvieB/1rbGnrAKvSYF+Dz/ItGuitpnf9XzQ50RMt
ewOuOCCrEYZu0WbZqSe3A1cN/n3U6o3pnhgXK5VzgGSzvIk6dGz/10dWsDGpeUXk
n1bsRLYELhKto+9SvIpDHK3Xd7Ug8ghPNuA+Ee9w8lo5U/Px7Wwz/GMLOakME5Cd
d2ohzGOXFhah+41vYe5UYrhiTQwd2Iiy+GvZ+oTTUp7etWUElvVnEXndVwDdxfBJ
FGq6GFX7Z5ysP3j0WZvdJ787I+KhtU1wGQ4hMP5oWh7upBftBIn0otHZlMJxORjC
KWJrOb2rL56lucE4CVhfUGzFPt+WXEKjAk/q8QWDb+LnAElQYt4aMQYQ29MVzVO2
KSmYkXhORkeH9jsiEs5Omkgvx57JQADuugvfHH+szAVA1uKmqEV3EhhyeN9MX8p2
BB09ckFLt8M5G9w0OT/id3sYX3LxqWgts8cgx9mqiYCdaQAor3suO9mYEzbbBAqZ
iFpwjDIvkKa3fiQmVxpNKDJBV14VKOpw6WYlGqvvPHHeA4KtFopQr7WeJwzgOcX3
Ol6JG3wytPdYhWFZlesSvtUPDFwjPkR2umyucgvtN+XrJ7k71gcEX8Dwv3cW6y/4
wpwAU/eupUJGd9yVYRSL/zFIOXbqi85TLfv5Oi39v8esw9srWmph6qrLhYWglYbo
PA9AGBxt8FRihkQvrA6+jg==
`protect END_PROTECTED
