`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CRu/q12037KHwfUInuv0v2Gr/9hNEQXks5RYkD0K0XMIgmqFgyMhlVpsg0rlVxvV
zYhhCQ3/zw45tkbADSX6GF5u9fPyga3IyFfBDiEwwAHphFLVrXCxUJQ6DFTHdE6q
kNG/YZYHLMQpH70iDOzJmvq/7gBEgJxIptCp1qdV+chDBjrjnWJf8vuZnRc2FJcY
dB7voFmtNsmomo2PpPEGECniNUd6BIRxxirxgCqgSehivOPHDf14CsTbcXY6pWZc
Dsg2Px46TbTZ5mIg8OTWTCmI9gk0r2rv5QEC/1yQarqpPxdpPfjJ8v61q8MPK60q
W7Es9n+vdXp7XVe1Q6WSwEod7uIRRA22xEmO0TvEwP6tnXJyBtXDpBQaOeeNRIZj
FGV2yLpSOCgPNWEHp7NV3w==
`protect END_PROTECTED
