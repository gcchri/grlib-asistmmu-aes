`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FFrT4rzn5YO3OAqGh2/59d2afLRXBs31nG2F1SWJwfIboriJKhTs5uvgk2oRm5C0
rmENvH/7m8Lrzdo5lYwZYKXElOvTY6Bo0r6oOCZTetx183Jvo3S7GHD4LBqKGI5c
Y9f3V7vs8gepdNi7ihwh13KQ9aWptFEe9cfBTzhhY05MSgGP0RysXDQ5k9B22saY
Of0vLkbuNaLAAqQKpbkMck07uN8UYsen2Hb3iH+Iyenh9wdBhX+62DpizdKsrF2O
m6y1u0GaIQLn0uW2ZZeC6dr6F6BYvyTb+GoWZIobA7VIE+vDG1FL2rtlJviJSd0X
UjDSE4w4TC3oT05EbW5kC3UWIR8ZbkVGT0g49RofITzh1BXORQ5ph25XDcl0edkc
GWzin/RpXAP3IPIA2vqjw0SFTUi+Cx5UGIumJ4AjYf/Oa9WeTyWPXoOeEzU/BKT6
oyA0LIBDkdr5BXFrlIMaZuzseGEk89U8Lsm3YaN+ZGfhaRepV3lctsrhTeKXOGK6
8iyAYdjbZwnDzGGngmPP920f4UiR7ROOiRZV+jbOFpt7dV1XXoodjUpfLGFom5wC
72QLM5OEBerbG53B72hTBfU5KXphOYb+YvMMxT2ZC34=
`protect END_PROTECTED
