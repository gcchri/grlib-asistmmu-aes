`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wt1fEVz4Y5WNxfT0gKUcQgYqaSNlMnfvRuhyX0ZD6gwsDEIIhoOaznJOBhR1c6r
U7wgxqO9rS8XuQpXGmsoUByK3KokOTA+IiyIvmzAGQzBItZt3C54L0xv6oqOE6Ie
BMcbnMjOZ2WH4dFQh+q/jx+QjjxlJKuBj5/JH7781ihMYkQxMQ+V5uaalvfJ4LA0
aqEAioGrWxB7+z481axrYeI/XifqXieiwVHLwLEEAVfEAAOGkZ8Q+mnLerFnzR1j
yI17yFeSRjkkttAsBiwmFDsSwhiFM72pivwr9liqARNCj5OyVJy8cKGqL8sURNQy
2KWZBiSwWzE0+3/zeVWzK9rTbQ89erGidrGIbJIYnaErVI19tDyFLosh1RMam0n+
4ebj8I9q0rsBpuXxCWmkFv8Il2nqsm5An+ACYRItg3I=
`protect END_PROTECTED
