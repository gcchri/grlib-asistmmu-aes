`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EnvyiHJ/TIxGySLOXlh0k5bbwErtuaGBU0kQ9vedFZB4uUsyZbkjmt05IpQ71quy
TwK+BTUh+cDUWS0t0uQuUXTXQTg8FZQkvjJ/P6b8WvGnkZxhnNYhBRZyFOpl5fZu
ygbHSTWKUu/+Ha2S2bSm/rAUmN93MTDwoSh6KoYKg0xdFNKZy1a+5uiETfhPONdW
egMTCZfp218EK1zfS5u1/hOwyZPgxnLFIaLd8GeX54Lvanv1rEf5IaNA6mQiHkZX
ennfZ73YLygltIdZ4D7HZLXPw47Zf0i4Xk1Ug+tLDbsWmIxZqp9N0fVBmDLpxgZ+
WYPgCxJva4omknEk5TPJpw==
`protect END_PROTECTED
