`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVRtygrkcgIatqTY1fPHokH2CHYanCt3CdKdmQy+sAacY6p769ftfzum8i4ff3qD
8noZJ5y3kK+p46gKHI0dWtTwu2XmiYiCNypDV59FVxYiSveW3u5Wl4pCviJsgYLJ
StiYtp+9H3CE+qbVNjSLJ8XH3YKLqrtz6vCoVFITmvaIHz83mGcyGOnys2e4nwXF
zdjQFIu1Gb9kirs/N20sxBbfaL92tWeKCgFXpmEEFApYOhzq044CFBezGvJzRGnz
sJdBgNDAdsCswD31lbC3ZVs/9y4dbYuygG0iM8DAWHoxoxbgmMj4gU/k/IL+OIOa
H7zKb1Pt7eOrdG3QZKsocEqTg5mG4JEdEiBGE4lsul523FQx92lowLX/5Wm8fwSV
jvoa98l9elc0FgjqkKR8zA==
`protect END_PROTECTED
