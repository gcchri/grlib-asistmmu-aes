`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0WQgnadMN5L+RCLV/W+MNd6PL8JfKuMPNo+betqpfDLE0iuOC+xZEAdLZO6H4PFy
jrZEk/82J6orb/+XomluJ58ea/8SKw1lqDQ02b9w9QN9c/EMnIUg8K+erBjhZzl8
nCehocXP1C3YKacaxzPqUZRC6Nt2jwCF0uVr/VXpBBPz/52NQ4yHw4L8waXOuRW+
1BjWW0WXwFJUPwrW7BXDWWJCa3PAuLNDmbe+RX8lAMAyVlpnH7w4WTsZHDZKH3kr
b9rRwhUwx5kVcAXR/B+UajWig95DCvY/lauo4xgd1qekiwQh6bmKIAQoByyMf2uG
y+K+w4mInKj8IOznhckThiuNs7fM+SkjjovMmKu/zHPPPndhM+mGavOc4JT/69LK
oOq9e2RP6iJ3BtCzEYYuaQ==
`protect END_PROTECTED
