`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+hrz2DsYiam4LEMymUW6GdUUm7WmpgggWfAmPo2zfec4ge5OFJ3ffTlBi1AaHLs
gPaQOrxuBNUn0PW9YD9NSiQjb5F6BJCZVQJHcvmT8iW0dSE3IQa6n43825iaBGtH
UH8u6qB65JmLTWRrh9eE1r35epa44nUzjS/fzfSWqdlFSf29USJSUYc2GUl84JYl
OWjMtunp4ELTecqrKjr+ui5Wnv3iJPw4eQy9NvS2NzhN8HzOkizA/bXm0lVaZT0z
bbMfxfMXxHNJrx8/jdgMaSVMMqjF8j1CbWAI/8qTt+eJebDcYwPuGaLKU7lu68rS
97d4E58BIQJzWZbWaPaBVHf2XsOmO9mK8lhxoHJ+GeHJvshKo0UtILdStA6U9sGd
YsPeLRodN8eTtek92H6n3oiigsW4ZVV4IKvgOaq7wFx0+iB0567hyyK081MPYO9m
vIYLhgFs2LAjjLNNUBy9J6zagwn5NmiV+V7vrqNsanSvGElcHq9RwG9I4UjQQwoR
2zz2gEIWccMlT4JlIlQCsC3TbmrtS2PXWhjLFHOWYAlbqNPiPBMm1+Z8TMvmfYfO
vKDbnxKFNybEvedE0a/ngBIC0AVH7JFPiqVE3+OpQadyWA0uN6sux1guDeNrcaf3
XfDH0VmqEwkPZLzoiaIZl0kbjooxYtg3wxUyKGjjBc+rYnxJsfbzGvh8Mop8t6TI
XFVRk6a4oZ4LIbpxCGW6nUzSBeCw9idjry9hWWDD1i9b4nCrXeF9tEaQJgxIlESa
2R7fAEnFKTT92wLFEVnpdZ1lk0/JSVuQ3cL3o1JBXRiy2LYxrJgbUrnLzaXV0W26
eVbAdQKCet2JIqkdqoHf7W68W1W7rutxDKuIx8WtUW7Egu+5pw8UalGZpq0n+/oQ
4Tlx15xCSHyRwAqhDnC278lkvmRcOjW3rlkQvMc4ibygZBiMRsvdGcYhAfHkTbE8
ph1NFcXqduXX9noth/bqa01FwIDbwQehf93Mx9j5g8L3cZd9Z/71shQ+2Wthv2/P
sDH86hYzJ/p/DEp1IN/z1HSCMnkX1GdnmQPJ4RNtFrPbzkLTnprl5ZXMGD1amAWX
uNENVKgEIKlIE2vae7KHhEiHt/eU68ELZaLmHZyU8rckZQ9rrYWEPUt/L3IdYYeA
5/49a3sZm8cnv/OOhhDu8/YDKHkLOHIJSU04aSJCQ+0rTBXnX7ixczdvqCdbERxf
DNOgsWmwzzRxmGXSYFNq0EizMcYLamuoA3tv1pvZgMLbXfIW7PkV/MPx0na1jIrl
g6NOeb9E/4AsxTsKkzsJI9MU8bPWinP0v+M2s9nM8EXzpdH3xr9exXzIyjTy/c15
`protect END_PROTECTED
