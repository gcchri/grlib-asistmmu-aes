`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LIZ/gOaiblv+CgTr/0Klw0NOfvHfuBbaqifAxudzRxwTA49u3OU9ALN21CviY9A4
d6s5Qz3Md7G/Z1kL01KAzAzL0BE1OtpRFoa0kV3VQWXj30gk+VYv44nP3wlvorhi
LfK/AWFiyZJOpJJ3mosCjPxtDyNqKWZ9oWfDVhOqvkgWsrHlI6ahpRlxnGwLrXmM
7q2gSltX0Y61tllnGKno4wfGa0ge70gdzpbueo0re3AvNXVnCtW0NtZ0P9SW10Xi
Yn6+cwpbidAn3Bpxz61CnEeMaEZLXYsGn5PwSv+bCqmataB7iwg1LLPu19pzxoi5
OVymMHlDVB6plRWoJvaLrgayDLT0hDejMlsVxjn1+19BGbwnWHuXmBsBGjbfqnpZ
xtnMqFzFTfccZGW0dV1K9eDatVRKwcGm6X3Q4Q0DBq8rEAJJwGyUYJ8Reo+AM/sZ
1vGahSW2h5ypMX8NTiCFn4AjeIwIASkepamWiOSerM2kk9tVAJQLB32W0B1u1sos
DmjHQnZAQXXJrs+AY6RFRHsXCN3eiScIl5/zBVQZcFoBm2L0zxzVmq6EYFCa8Age
LOvtrM0eFe8CIpB6X6C3mw==
`protect END_PROTECTED
