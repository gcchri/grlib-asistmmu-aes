`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMffqWbWxKQDlaW+DKZN8JZBgqPXJc/m587AnEVEmcyLkY/++mcJWkUSN1riu+ID
YwYcby6He1g6WRHE/FflPdd6IrXYoFErchvtJ7WbArDbSfAkZ1BwHrjcViTyuLjO
TnF/jr5GpEVBQ13Aj0qpG2IMSi0OAGxcVxy9xzyNkPqXYlKExtSt6FkSRHXOcKJu
crLUD37dGrDEtO4z81dQDIGcDHm6X+Tj0VwMfQ0XNT3um/LapRvAkR4mxr/MIqBm
lFG1OsSMjq2ggfKs2aWEYzaokBc3SQoekpIj7G3coQfUoVR4lMiwetMEUhXkZLg8
aqqRTrPaQFFktbFUxn4domZJfYrt0zFpZCzcqjejLG5vNF2xAIiLfem+Lf7/P/cz
5Miz0ivafE0GqmMR4xEMNdmvspnmpkZV1xy5GM1HnPCVWL9s9zf8zJEoEPQVWiuk
A7fAPFnxIN9O1jtq1n1+F8rGe3YjfrS0HBSE/ZZngvSsDH+M1gjnAdRocx+GmTyA
a52IPKzb6pT8R6xwkMkrnrKYpFYhr8JrRTi19bue2iRkrvUQ2ro+7uhWbIaanIr8
`protect END_PROTECTED
