`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k5syfxbsqnAboR7b5TCAY30R4zgMJvcMG+Ok9ZGoG6IIeQULwP+s/vBEtWLFQOld
tY2x7ww0f2zj+uteEAwQM90BQf3BmVl1O318mR48+F2qbeI+AEPIYsBwOa5tHfYZ
00XYEYX/FLtlea7aVbVKKZwBIyPLMo4NzhKy4rjarGP68P4p4QBtgD4ryXRrTe8R
isLkXGkTfNh/kpSjupNpj5NGfc5/fmHUqOO0deMpIg3o9KGW0spd0wrRBEZB+yNb
P2SFoj7xtmP2ppzx7flMYFbQr6x6T8I5YFw4Ha1W0a8/TSPkxCE2XTZqdC7JUv5k
fjGGgf3rUMjljLHFy7WCQSPqdzGFGXAB4LUtYpTFMyq/20cfK9nTEHSCmk54T4Gl
dXKelHidLKw6sSz1pFtIjEM/YRES8C5HZFf/c4KdRbh6XbymuRiwtz2TDRUxKLTc
flmyzgPr03y4m8Y833GCnESQbiOWxPeb9JY8eLespJZnxry734NiE8he3t03NGWv
xkYjQvFEB3avVO5ws7WNJESoCP5PGk4ndxy4kLZw/DmsMEaeVXLF2A7PWR1JNEJF
EZ8/0oXx+JvVcL1SCo+t6y1AzwaHfmw1eb6hxF4Eqo89AcHpXHHyYgK0sBsY1TVy
/MNhC1YZeSeApXAanK4x6UbtbovaSX++U7Dg+yl+bexZfNpzqGFxLuy7C61etnIv
1IYa9sCwH71kgY7yigObh/6CgaTQixzcnR7dn09ALK8ts1Cv6Waw+RqGqkFtCjOm
KMc7ZpVhiNFyC1W+j2SEFyxIkx0ZQzAN1Oc1tYhb4GFrkpAU2J7IgOll2KsmUnwB
P9dS1Mu78bsAtranU1xQ4qTNvRh/fSVBxPnAUehitOjgTe5owsmv0h/6YKW5H6pP
YgfI7ZeW2CrFotZaJQ590UG4A/ngkAIpGKQedw1yLDAPnBgFczjpYyYH0T661kbB
4wt4PNE2hl4Q1tScYwvSMgsVtGnWEAYmhjNXyqB0Vl/yXWQFBaNHHD761Gynjwit
RTxRF2rutn+qWRG+Nj39BZ/m4wRpLYVBhdu4e5VfYYVQFJli3moiK9zV1py0R1bp
L3tx1ovSon2VvzYQ7FneM285/XR8zv973DIlp2+OGQZQlX5iRVkpfJU7+8U9ktSb
CpBSReA+0kw+RAue/AC0K6jYHn+9JR7sqKmDyYPtgddTW1uvDdr92y+HVkQwQvAp
yZJhJrsuSWjTX7GbWab9EjFKYrKEeuPoKOzSxAXj2lgQIE6zbWqMTCFblBu8X1io
81tpISi8+DoWxCr2lTuIB9kX/2OXNzItu1B9zteGQ9RtnZWtUal/FNRxFfMeNP6J
O03E7B9INeU9i/HOr/yGEoEehWGW0lNaQj7GDtmP51F2qHvY9L06UlLlouVINVgH
pPEmv67lBoBxe7DeCljC22366xm3GrHR7/G+NLd9OE866/dlOKxrXWiP44y5yV4z
KdtaWrhxCDvAvmmeF1xuJBksdGUh6rGFfrA3D2qQfPFB99orUyTlApLBzOEw+Uzw
4w0oLNsE5IEF2HQ5xG0H9lqQGOIhxbmLM+LXSwdzu1a4csvYLqQOrDBVxnwgJVGH
77zqfRQeecmhwqxbbQVYsROUxQ8hABP2gyz99tq+72pb+LD40T7kwIWTbNFnLv9F
Oz87sF2oJGUV8eZuXtHAeR2jNz8cbjvD5v5r7apwGuVhWVFSrmKJfXRFXflpYU/B
4WvFlI54wsS6OrLpY0XS8/GxEDCyFHB0vsjqSi90XRknjrt5HIOShB54wj2gY2MQ
bw2WYG4Ha4vY+OKiiu4GM8dKjJXurLnmxLDOMXtdAgn0s+RiutBhCCjsMGRgtj/z
nQmKwU1LR5igDEeyj6ZF/axnBbEBze3UZn39d0sbTM9jnyqZxHUmhFhqsb9RVZAB
PDLYTE194c2YOHcBEv8FiWORluoc238zhkzdmANCawxY7pBZSKVDNtkJGYGhMWjX
R5fVALqAuTHLYvGTBXMYcvabwS5kdyPavGSN2yEorJBfcZQ17S/HWMAMUEJfRWo6
TKYnmUHBnRVwuWhegDqncg//thxb5WtKnzBvEL+627kNT8MOfRwccm+nbl+sXAal
CS/LwVQk/ZH7XZRyRBtAO9P7NVyDjwWqeIscbDUGAH73heH/FUjFVRgSZONm2Qv0
I9GNF2ioEtDk9rWMH+UfgeIgDHqoDJFktAnTBy3Ss/q/eTkH+gdGgM2oSSBKuWRo
+knmxHD2MI9IYsyfT1poIyg7AGi2tzTVpkGXH/XB/n1DUItCjLJz50z1FYXHxprs
io/OZvT5lH1EHEufQejHL6t7Y26K3C1QeKsog8cpimkDxX0IdEOLbqPAW+I9UZWs
CYmFtvYI7zimza1BVWpgzDeA0/UXNBmbkpuYc+rWvuYe2JHERg32DkDB9rl7ZDWk
9J6wr6TE8njXXFUJTCeEWMRqVjvWxnx+ij2xElDjf4hLwlYALdPRNWz/uWYdOf7L
4Udjim2EyZP1AW3FZMp08ty7cmdSW7a88I2l9rq733qDKL2dBKpQqj1+z4Wl4CPa
wHN6e+NA+gMt/IERhYTWAicpTVNM5QrIj9saHnC0a1eTHpegiX2OZfMbD7Ys2FUl
+sWQGRGcyURoMeRwUiSxv+FUfAeSUd9MXkv97HQjMSWsRq6PUhr82AHx5pnppRDe
uuF6j3YOtwwKBkwNcOoKU1SevN2gdcbvUScYsQ4+praGXL8jvUR+GK0NKNA1NiEI
z9c5TTnMFxITHSNZawDQxWoJ2oNa93NnB8gT6CGABqjiEBBsT7RE+C2yHsXEFFha
GM1h47gRoq2JjLD2N+9S2zD3pTUAyxBd2bWrWhjbU07dhBhmgOArz+uI3MNWCXNq
I+KKjOejRwjXuqjW8oTuw2PV4wCGjmgkp7lf+twxOo8E4rYPhcHbz0inicnRbX7a
Hp1WHCERtaCZU6Fyty9LrPFFMKMcmro5CCKnIbEbnH0fhpr5vQs3tRBKpn5aQ1mn
Dx5jVqXOhB5WBBvd9+QAAKh8w73vYukoT9zzMkBpOHbCzDe5vm+2Dh4k74d0ryfH
oYiJ7u+1HqiWDpErxV186yCnJbnmYAcBHViv+3+AykIr3QG5k3U0B74uagsru7S5
WnH8bhWRwCnMOQHbxE28VE5jj9cQMeA60j77zp4liudQRLkStfKiCCTmxXzP+Vdc
Rtc0RCVNrxODh1vDf+jAvhWIRwkodWwxAz++rTvV7Ba0crfNy2TFbtUWEkqCaaVy
jo/i/IFR5Y9RQFkaj07NVCvext0EQ3wXWC6PmANT6SJtqJ0w3ON30AnJP3xKaSZM
26CF6rC2GpgJ8sWksleKQ393dYyOMKdFQlZ8j8UpPjRhEFxEX4ou1TA7rRAorYz9
P5SMt48vH6wl1lPoN86u9jylF0Es+BKn3O2wzJAEYzQscC7gaVmfj5aa3z1MTpGd
fK8359q0pkQ9VSTqYIEtSHNpojlvWVWqR/PFG4aXo9gZpSFGHDFJv0FIQKKvBzUL
7mXLqq60i0kAuuyR+UPGuyCDnDV2+sDEgaMWeM6asnm9FDOm0nrCz08gQXvUc9R/
K0dIDL5motewgLqEEeUjTOkr7YVs68eRhsqA0v24kGNTvv3P0F9AWSLa1xnBNkKo
MA4Vq3BNN4R4qQ8AF9pWAOV/F6tDkjGax/sPhTPqDsN1p3cz/w7to8gdVt/CxN3j
QgQU17oOBlKdiZ/htlu5Ns7vGTWBSiDcKKw+x1NfjzxPHND3plldQkUIN+h8tPAT
lMRY7QjENoSGV3eHYOm5SxfPsM2kQJDrlIjrPiohsWUPYKiFvZFI4iPy+BWwGdz7
C4R74p16TCOHDMTm030qKj+elisLuPe3LlK4z6G3W4cy3aPxLI2+XDqSY/i+pYMO
igunYQZwFOQmntGNFKp6tUveSG/xwvJ3SgPlTttv9SuVNw8EkTYG+L9k4YvIllzX
hvlj/IkIs8gOG8j97VIxQCYqUQ2ozwIDfNR5l2DBWN4nONVYoCKhXVlu0fx4Pr88
xaR8iN1OMGxEbpo2AB8VUakbnYwS6B8tA7bsWFfgAFjsab86YLkYzQ17q8yuZvXx
SOW+MDr7c5O1HNflGP4/GfuyqNCJ/j4pY7WVVrxQtVRZT8J5g2WnRLTdu48YNnvA
j0Bx6a5fWfA+bqg9L501r66kbcounfRiM98ebpe54BCWNE6krLVBmUrNZOjOm6QC
v6G72fPRlWEXTINCWiQbZ10KG56Zh75q8QsRsnWiDbWaXUKu98OwjbD1klWx43EJ
ylWduWEWELvyJxbZt7SZnObHaKvOUlO+lJPRFqpF1JwfKJK668BV/GXICtvleKQ4
M6JvwO8/TlkRVF1YOvOw0PzuUblsPXJGoMklLXvFzMBqDLSZAdHI2wQxA/QycG0h
y89XSj32m9r7KEJdzHV0xyjuqKNlDRk8JG5L59JLFNjJiTXXtaW8RH7pS+Tw9ZrD
kKo8vp8WUMqGM88ao57WQTAxsMeQn5ARVXM3PGAbb+4TIzAvtrLLlo1+KX5dzHT6
TeM3M0rd6rTF0VTIK5WedMkTwuMZh9B1+R3JHbFuJlSNeO7ztX1IHiMBm3dpKPU2
+6Iffl6gWoN4DjHonWXQJC5Ty8fI4xFfFz1y9lDWxxXsVduNMEc+9Yfz/flXyL3I
yucwDdeTNHxih/eVt3B63KsHc96aSuR5/T4qziVGneB25exA5vBbUiQaWv0NmfAq
sRqzFCaQWGl7jKlXK+ikFxOfPKFx8kVKDslK517CyDcAw7ir23pYaCNIJdArga39
4ju5CC5jJGOWNvjR57PykvJ2+ACgIrauOLDKdzHWhGSr4kBL0DLCRu2faeH+hchY
H2nCHGQ4C27DOarTh7NWLihQQDd4pRHg4/16yg18CCwmBvn0seMz5KqWRD/2gdTf
vEexcprkFfI2X+TEk/DNytvUO6810zASu4ZM6UofWu8d4Wq0EaIe0cvkv6YQxgE4
Xms2TrCXJRhYQAED0ES15w==
`protect END_PROTECTED
