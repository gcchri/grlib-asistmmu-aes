`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGJJ7W3HhQ3rQfwQAm7pAypaTNjo1pTZVW3aqsj/ZM3ksR3Vnx7Jp43acsZorIcM
iA4PlJ0/D7BbjSUHmcu7s7RNEsUnbZ2BIWQWDIqZuYxmXBBE+ROisbyxxJWLIIN2
XHl3J9KjaoWEchNcNNnFqphbNAwp41CIpDBQsIaAqqqV0znJbs/jeXXLz/OXZWCQ
s+ibspwDuVwFiDAfmDLh8xTr243D8t4dGspEToiF0J1z0WhmISVxgt+1g1xPyTby
dHGXtXFnPHymhio4G7pcTaPsXOV9fOYIfbj2uZnudVau62Z7rGXwuP/MQ5fLjc6q
t/c/uvIm5f7MS5yUH3UtYLVT8pxXXy6Z1rEtxfaK3iYtEsIchsLuurJ8GOv0Nyew
nNKYN/LrvTZ2aK6NDPgR6osEqJrLTBP+s7kYvuE5HzE40lWa8iQa47XV4QlLKOqR
cbWhfT/3WNSY3/PtcDwlIc5bfKS8NQzjhfUEE0KJI37DzsNyrqPnZaSSbnTWZq9w
gxlQ7Sugz/s+TTCEIP/xhQeGZtDSFN5JcQ/ski/ld+FaSpM7n+Q/0m0ESgCWpaku
WZaE4DjpNQW2iJBWGxgvHmiI/EcEZ6v7m5y24yv6ABjyQC10WItgyEtenxqT9dIu
M3FBkzRD6dGkfkaF0AOpcHDC8WhXHMQpBDG3fCU0r3QA/TWwLUak4U98WpN0S/VV
lMSBBANZQg966nfAxT9ESRFh6sSGqXP9btsQtyyFgCs=
`protect END_PROTECTED
