`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CHqGPc54JODvqJWXMfBr+oxwA80EYQVq5iPbZrGi+xQD1Wk6IZ1HPzeE/gVObagh
YUYqM6BJ5962iKQAKPMUQIjX0oszDTKBIsv3dG3Ic/5xWg75llsPxPzqs9+mDleE
efpUApS63u5I+TRURJff62j8k4ZeT9saj+Puj5MkL642aVRQea7jYr6/CpvNWk8m
kcbMrzwKIYfhr9f/AMghCa06NgiY0UHUFRXT2mYERLbqE55hrihc9i1IWi5vT6ed
7YKLpY/NtOWVnpDtKvrG9hL24Vul5VEPGesbXDDTbbfNiyzAtpGICOwlV5cLI5qq
Rhe4GIkR36R4x+GMufExTjXjeFK9h660S0XQR9Dd1AArhJuzwofjgl/JDpQPO4AU
q/rLwUbDzZGIs23tvkVgV+fpDf69eIaNo9+rwH6kZHSjrQ5dOFSo9Pbileu6IJ5L
h5wRCLMKH8a+1OKl0HOWfpm12LFzaQOVODSg38j6WNKZwMEwWKAyZtE/YLuOrE/A
PoozjCO7zBgy595tY/5dfyWcmIvknaNhzNrSeJvYYu/MABb3w+975u0OIOxihonD
i85G/53U0p7zxONQ16dJ8UNIUi/Ck3DUZ8XPEspv+i87KLfKIArg0cPet1se20XI
Lubv/d9pLk7YSKFpPgW7jw==
`protect END_PROTECTED
