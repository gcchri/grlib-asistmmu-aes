`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0EcJQ1J9XGUNEbByktZ9t0GSma/CRNWgu6y8SgAe5xRxmzQ4jGYf+AVP3h/hGnxv
QD4iOTPG4zzOdolM55/OvWOwp3eeMX7rwd3p7fQfCl4vfXA6H92eYVjdkXqpejbv
SFufCm1j2rxeVYpWAO/wr2TfcANMKcw7RzyiU/2NzO8hIrxPXwo0MRMuxZWO79x9
ERXSUEJhRD/T8Fm0/RfZWWkpH0H0zt728j6Xl4Uvjqw6kSgv9nBkd4Y1nXgH/l/0
wKbLK62w8p/DlJ6uSnhaSZ0EmvpQ/r49ndfGUOPiGKUnwSmEx6BEl39sx9FVjURn
pV8k/W/S/9CZBHB9rmNmDpi2xIaE5trtvakqrTrVnygPIXuVPNN3WPMhWQxVw2Xa
DNJNsvGwgT1t27tWdM6as6F2zKN5r6N/cJ6q6w4S5XsUxYOkJ4jdia1YOmagaWEn
zx4BjfdedqIQ1LTBUNdOPq5rqxgvO5IboeN35cjR/hB5rjq3iw7X0MclTLE9u+m9
`protect END_PROTECTED
