`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sk/3BJk8mXi9tiNizl5hlPvK29Cgf0fLepQiTKOI8aCTc6ohSck3lVWdLifkmDg2
QBqCTEwEFCfwRzSDWVYUZG7JITIRUohHLV2XL8j92cRIfUkCzcHlk3ghIiATfTdC
7MxdfwTklRrBMg09vo0VrjfhYIOZch622ji19GHa66fZwvaFBh/+hJxEBZnEZKM0
/yDV/3ZFFsdqq5BvK141zkCvYQY8ePSJSdYqBnEifou9xr+OW5UBqcUUIJjy471y
O7FmOI7ZGRLfUYo10Ae0rc+jkROcQpIELbsnkJMqw5GgaEeijSJkjbaFewftI73E
TCmO981HUc4UoSSmu2tKMb8CFNVR79bQym51TRTsgux7ox0Nd2o+ITgMXYZYopUe
jszDtgVUnqO1KKAnJjk2rc0twhHNqqSalX+jU2xo9u40JpZmWvCur3MxZDbcNxLz
Bor0103izG+An4quzgLrQWWHkoVlTHEIp1av+LxVx+cY0Ud7clx2qNiY505fullb
fjIHN5P+rc1RFIV8DMV+OG3xIuulBcaqensN1OBhUVNgvvzP3oWjyDaKCbB+JRt5
knoaeuhB+AwVSIa6z8KoA0AN85Zo2Kwx6m1kOL2/HbL3Gd6rhvT7cmKVr3jm9A6A
JxwuDTboj+hgvnC1MQ7gyeTR5PUMA3+xXtUPVc1HMJR670vshqKcMNYP0arF4IKT
ISZP9lUHlcuSXuXAxwQ8fsvF28kvQ0whkCSkZwoI31KHAXxG2LwomlO2euHM0SXK
wEQAZS+AbGIR4rJu13TGYOJwUoiNP3vgoZRHISqz5hF8fN7WfPokFvo3klOo63sE
52jMS1rffxDTQ3T5XFE5MJK14y6rUp9Z+J50HPFfJAmtl3wd+278s2+4CE4gLqJp
ohQ2UWsgg+RXPlOnZM3i/DD14fBDfzCEW71LbtrkIK5TA8+YSya7FAPwnuLQOPee
2XmNgNI230De4ux/yemFjGMqW7TECe9rEkfWwjVu/twpdtvVaPZl60ILtR/7dMZw
aNKdybkN3Bxh+ZEjtKvG5AV4YBBpWntdxCjOIfj/TGhYX942eXrIQxjRb53NETct
33qpIVw4VP0Sx/dCX/Ty53m/wmgJ710LivEL5wAZXNDaUnquzJqhR66S+3yIN74l
8edVfYok1+1T0u7DpomNiiyDJ1MBoOg+ryl6XAl3Fqy3f/ag1EdKbANyiEwGsbqx
81SNUIMqHCP97M2a6PsxLTnf2PUjP3Ek9NnLEeJRUKNjEqPTL2uoMxbHY/Xe+apb
D8vbjPPKjlBdINTLl1wQRyJ6vN8Ug6W9GKj3GEBLF+jYlqMKzZnwLBkDaOyrTK4v
K3qTdM7rauYTiPLHx5MMfQp9s+RFrbxoUACkBN07HCIDt2yov4vcGhs0D3nO4Ub4
2vwi02+16+e5r6ZUMWfCjiJy4/PIVkRaRjRTcyVlL3i4M2HHgSN4YlAI1+2RZ0fy
hfbBgzLh7WmKFIMvySNHqeivRGPtwlW0Z/h5wv2W/HCUSMdTQ7WTeWnk09qbQ0mI
i2TcHIRKKzRMWNiihcSiBCM5Oh/XyXZg8W9TiRFkD47sgjn3PPsMedEQBHI741cX
vklsogHPnBkgK4se2wigfFZtfv7lRWNHiPDsbXazoocJi5PepL5+VwjWGbxDDN6M
Lt7hZeZuS1fR7ohrOgfN+OgoFnUJncvZ4Pd1tSb1nY2z4QQxNwCERKG/PY63NM1/
+v47QcKIk9gD2Fhhu6kN5NygJgsjpLQobrI4aaRk85zPhw9QHGErLozS/iBIWcFV
/2+3KKO8KSOX/bNIoRpsRIWfVWlxDIocPRz6DYDTY+GKTm7ozM776guW9Y6WGK88
ktkLbOK+P9svaEwQlllCDSnmoq9sICVbdlTXC/lDWp4Tk6vT3/KngMlxETowSB7V
sOdx70T9Lt6B/y79PwNJhDMpKrB5xguzx6WdiagLpEkFmJZ/oau1g5euekx5LqrY
uyU1c5saDizRJXhmmzwyMNmBOlKrN1sHlOt5u1xGznC4xn7/FdbhX1P/YdSVxFMq
tx5kUogTss/bwQTGK0NOogyEJ+2LC+JTpYscDNXt72EWQfDa6jSfUW238FdR1QfT
IDzNBlzXhqGrBzy5jWdph2jgcz2+5/0Fuqq+R0x9fUs0jH1UhlrZ7pS/2dq2b65P
BInm6GcsuJDns93sZ2/I6NUavtvnww7QQ2H/Q9MPc/yG3RZMoupTww3sC8IB2QrY
hBi8VponGK82okTmg+2EPfzGMWDp3IaoanmNXNyc2h5XaQv/VxXNv0374TzGMIh3
yaM35RlFF3otseX2KcMPTw+tBGFIcBDVjeHuPJr7M3WBsMQGCOqFIHzLEc7PNAAS
UdbjjCYXfxTNVDPafzZ/4D8WRrPlDzbNJUS0izWa3bvTzqCJNR3VJUg9FHFimQCM
f74pzPKTowi/D5WfvUKMpFhmqPA19xDTt1PHGqafE/I819NiRu08xy2Omo+rKnAf
djRZSnoCjmiw0JfHrhF0AoR8YEm65oG4vZAatGo/dtojKc7nkQjiV4LCsR2xgm49
UwShGXJ6a2WvNpLQwtjNwcoeolOqURu5fQq+pagO87Bi5d9u2dhK4sAaVg1JHTbU
/fDyTovwH6lPTdI1nBhAgBJMcqKE1PZixbgzJN6RDe3cNC6HDciExkBcFVQbMePs
m5MrMplWq4h3CU0rWOGJEkt482nYRNyiimZj+Dr0KZSCZuMLXO1I9Kso74ViCKw0
Ycp62Rpv0r+U6CEJt0TQZE4qj2wtApplYwy8sw6Mpnnnycls9Nb77lrMJcTxqqUm
exWgRmt2KIi66q227dkLN8lCjigVTaMzQx1CEVCQ1ipFnaCzrLgzb7C1KbBYASsv
IVXUN6Y6Wvamb7npnlFiQsAHEsIse1+esJygfR819dl0Tdn5eOg1Q7pZhoZfnZY6
8FsMeeDvQct/gEMCQ6Pn5myXMcV6tR2glZoEs2PRCSD3/V3qppLh7F80eYcGaT/r
Y8kjlnmtpxWOIsf6NKb1Ydt1wUL1Sj2FFsLCztxdX1JhLnqHyA2eg04hVHpnpTLP
jeFefzGvLT/alshlixiU0I0U91L8s8bc7I452SG5vUO3XgIYtrM27P9fvHiVJpMV
knu3G9CJHApZ9HboNl82dtB/g5fjYRT30MfCZIxrqgRCIZBWPR3bYhPy4KNTt28e
cXZFBdGdZkQ08yOBsChCmqbhDZ9mbZWX4WCbljcDet5B2L+qQ6FHYQ4mDau8f9oc
usidZ3fXdu7rw1PC4XbBJC8S3NGvBJpnHAPXBywg491JsxqzK56Aw0uYtBHWy4sx
zg8FvqaLyoMuQGwHKUotrL4AlIp+UwHr21+HkfNY/UtcW14egUZKSHlsIDEL2Xux
zkyRpHDoujvc8Zrzo0y52Q6duGj4yzq80QEe8gidLVs2oDK/5SbeCBMSGEmBS6zU
QVxq+668hRFBG0hl6Op7G1jE+Yp0UowqIG7jDjuhPNYgn5OmIGh+kJgfrzUo63UO
wmX5uEKj4pbC1xnLzL46U8Cm7IKPL874YkWyQbWuLxqssD3xKqe4Gbj01yC+ulkk
tYy+h8OuDH9jSW0C21SRIIRlQZ94FKOzhB2NaUzlXJafJEyn4hWTajUfrPpWArKF
SqUR7vJC8+nAE3sQBKXj/FDi7vLVcJBzYQteEDfmjiGeO+OUx4qwGzptzIr2mGNM
3RX+5ot6Eev0v0vwx6NLjt6R6Nw6NYA7417KPM++lsFSdoBrlvgrT50g4NvGhGGv
DHRhOEqByBqambTgx0xg2/COAQqdYfenzcX+zO3POzbWVvCIWjfuE8ql3XBjDf76
jZpgPiC5uBOkFhTp00FqrMYw3E1X8tiCm4PloJsIDXOnFrXN2aTzBBNTtVqSO2GM
Z7Q7inmITkYsHcuyG9LELbBQc/z6MqQ0OjNn1dSQ4yqi74xbnh2MGGg3G+NmXbMp
OW0+RA6NJHD56CjvzhyYfBDrktbHQtG8wzX3E2B4Vq3rTTztU/oy5VeY4I1eTn1e
FO2xxHL/Sdu7vJGK713/nGWC0HYDyHhtLRcsMI9k3Q0HAyeO1CjWLOMQkKHhc4Mq
+HBs+/nlZxgp5XN8nZYu8sW7WvPwXzKCkiSbbATNQvNywTrYSBRo7T8BY3o8SY3+
xpLOBGun1QVl3e3pUDO9QovJUCXOM/pPE1pIE0nNmXgADse9bjxAGxsTBOXxP6Ru
gDp9QwzIDTKDKRCAY7gDkRMJWSr3UTcPItS/+tus611FfZtfhWadoQFCKWVF0SxU
b6aPbV3wAIfNygVX5wJN9lPkzlEx49nwSnqrLhH/lk9niMs0TKKpGKc0EhNX6mBz
iB7wN3C5lAh68Pa2JfeWeGg+7j2UhSiydKhnreE5vNgJ1ByZeYzq/YPWwyTTJjTB
hs6vcCBn1pSHd4HldJhy6cmY6NyyAU4W9ubT5Jnd0pPoU/0/fRb77e5aKNF0+4VN
i5UhfFbO8xpxhawLHGK3Qhw4awNnIRCM3O+SKLJStj76N7EX544I/y1HufIskibu
mVRWyqW59dzE+EWY44Z9SNzTTzHbrl4jRrV9jvCltrVzUToh2i8m+Ssix0wEr5li
BzKnYXmAI1vNhTCpBqLr8PQdPPmbt1hV3EHjSQfRmHIxEkXoE6esUVgrOJ5Kl546
mUe7mm8MyRnuj9bBzOCxFlZQTWXM0PJ7qaKDFwobmtZTKXGIecs4B9B6eBZIJby3
VdQoVT5IaQOIA44+zgxX1g==
`protect END_PROTECTED
