`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50bfqtomJVUZs9cw8jYPGKwGX1ou4Ks7pSrbA1uPGT+f0Fog6qReymW0ALOE7h7A
eQJgU/yvJjZXoYSZTF2mnIrnUDLF98DNWbxW7nQeSy1SaWEUtRV8MhMhYxAHPUed
rXhl/QnuDvI0O7sk39ZX5FnrWQPU2KP0OAnF/Jvs1HHLxAkPC4URSWfI2zXEdUvy
qz0j/r34vHL7+sVjY7DVGTAjgYy+gspm1N8yKT2yyPmV4ULtzIYHkVUO+LKqBqRJ
ZWU5X6w9sjNIy1JwLnyGOW+bpr7cpsaVTQ6WMJyTtYHhKYM/LFysAGgEu/l+qDgL
o2P4f6fNjtHL8XbPZqmrgYf1LKf8ykRHK8rNUBos7Zj/4Fp4Dx3jPjm9UuiaOJCZ
3mgJKukVMgocH1o4w4R+njB2X1l4DmF87XjtFZvs5al8y2nD9DmiV4nmc97Pqc+0
7jZJPROxASqQGeuNcC1goCuJI/A9ZtdX4VRBDzpq1lOZR5YZrwn3HUoNVTt36NiQ
a4iib6D7jFf1rG2jMAINCJWQ1O0qu0c8vP6V4QlnuYP/iCWg39ZYgUipGMdoOn4J
laG89GmD6wYCpkWRbgJGiDYytAfmx5JjG1BvmS0zRcxcPI4SkNVLK8pZR2Y3J5AW
XbSaguPayKUbooK2QhpS5o4pbdx7vZd6kWWX5duud1L491pY1u7JdmoEBsMxX1n7
Gb81spItrTUY6YP0z2vj1cLwDwztnkeCjlzla1A1ijQSib72POl9oJTN6gig0JEx
qVPTune7AhSkZM0fjrsrEu4eZ+pW3oepHl7symPUbDecEOChGSyxWM2H3d5gGEW0
RYZrMtz24SmXfBUGT+VWQKtblyrfKXpDFzLclIRdmq4fztk24rR+fTjClaxRlz/o
y95C/bCn3ZpBx8WrfI/i/O6D4IN1aJsYj5qQycYYwbiFtE9+vw9W5X5TImTps85T
475PeUkpfUqK0FkFb/zV5cEMQ3OExFkxQeR5sjb7IFuTCKMmkKCEVJDNcZj06lDR
dVQDIuLAQo286cuIsB1Z090PmNU1xp0wt6m13zWRJoSzJ4oeHJjRkZYhl+82uzes
tLUmxvY5QLBdNhKzrRL2It4vgFXztChTuGawhDUnKMZLl68zlGuDpBQBA4yPGiJm
p4QFjVYEWFJMKXgx7uQUCfW7byfGFkmGCZ3/gnfo+HAH8xzCx3Mf2goXVF3k1Y4Q
XljfJHS5MtAUh1++lAIARSKNvI2rUPwLFgQGKkDICn2ej82FqC4L+OaTTP3WEeVB
cGAJj9bxa/ZvNk/bXbm1F00ubNRsw7/IuFyMuvIbNgzx4/of02Hncgx6jG/aot05
JKisy3uzjwB12waU6o0aSW7F+X0npfUojt/zhw2Lb52DNXg7a6qlOshepiixR5LV
kBDQpP6E/Ztmx/vOHMsWdIiDHoU892ZyPGmxNCyNnWMacVbv28aKXbEr1XPNku22
b1/GXu2l9o6LOtotxd5NO4u0jVb1TiaKv218m+o/X4GHtLhHR66lGcImmeQHlICI
t03k/LHZ1hQmGw+02OAOzucvt1X27PmcEEgFBd8vC8sOlJfcj3qTJGDf6IEN87vX
uzB3f2qr1AVQkju/nEg9gss7vSLe/iNu8ziMeByYXnMskc3gifzgiPxJAS85ulTe
4ZuqWJqUOIE2DREs1wmxLQ==
`protect END_PROTECTED
