`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNgYQ5amBsUchjDJ3QfykFEysR+whynktdRBrHLfvbATCvRfsac44Bqoydlhs1P3
IA9MRogeDOt9IeZFtWl9teruoV4XsVydB56DliEYA1VZUXpH5ZlRS2xJ9+hX313H
lHq5TfkX1SbOgSmjgje8manEMYeveh8UyS849zWrVOA8Ss9GBvsj6MTCLeTwaWON
mybbYaq+42kxg0U+zFJs6t0yUjdkRHwd4xtWP8RFiWPmYBFYfGuiPx0g1/iogVCO
TgbxsJyZ/qa/C7dpN6J/AnmNGzTGEOPiUkaQc4VLprGnE3Z3EQZf1KXeaNSzvtRZ
f2YPnrSAABOvcudA7AZ1c3D10l7liOyJ9Dp/kFSkE0BjCa0A1yooLUDenO0U5+7Y
`protect END_PROTECTED
