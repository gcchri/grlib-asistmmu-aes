`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zKGd2h8Q8iG1dPaYH8vmNWMLsBulAWz+HU5c1nj+m1N3G6sjK9tub8rNmIW8e8sC
b+3jl/OfELiX4AUjPBDk9xhk7UuF6pOR6ColXUPahdJaYvRXhErO8NKtxEmZ0Y2z
isu9iDO8lyxxb1s0exja/BCX9oVLRUjU07wpSFeAEeyIK/x2VqXoVfooJhKvueFR
ahQXUji0WMSXKqzbWBgjt0SfXPVdHIUykhHLnfBoA3eDyZryHpCE4q5VSq+Vgrnh
`protect END_PROTECTED
