`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBKkfW1PhiZatIg2mr658AV+Pfvcx6iC+BdmP/jql5ftoJRiV3i7pSgx2XWRfgpe
iOARWa/fCL02t2klOXtenXvIF6j6bluH2CD76/e2Ip+Y3KTEJyj9TvmW+Hj5EZxw
cc8vG+E8sUFfiocC1PaUrFhIopwbeEhLi8mklypQj9WOL/aXmkSlTHJkAOOOwhnR
2O7k/T0ILZVphUWUKTlM1W5Cew/Wpg5dFVMJ0Ps+LX5uulG9I5gWcGqsHRy7vYAI
vgtoNLQsEcL171po9ZQsgbw8oeyiFXpY81KM+0hcNnYVsaQceTt/K85O4dyGkfyq
Qhm2kUhDptje0DYfVfjIDXTaPwYwzdxtMMSDwVSrvleNtsF77oTb6z3hNXZls3tD
gGF+7ZTiSHPOWkKXI7CBLVhq9J3AM47G5u1Jyg15N1BO+WH8LzNNEgKtJrwqI6gb
iQ23Rh4SQN1y96kXaMJTN2ZQNuXm24OqdFu3JAWJ7xC0jvHIzBXwoJkpJclnOe4Q
P3pv5cvEiRb9UMZIpm8mtXcUbZr3ZBRNNWe4eMcqmduAwcL2BlkReF5xXrsEECtX
4ddx6PIOqbgnBLYnZ9ijUwJxtNjtHpVyB8SeERcOI1rX+tngJTIYlEhRGWCRiUC+
7o7wc1AI0//3gi1E33HUEP+A45WNe5++F0D8OQC/mF0GvRuX3SUwL1N87zvzkmZZ
`protect END_PROTECTED
