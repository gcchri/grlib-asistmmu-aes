`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONGixhxRAzpP+Vbr7luUnhFJhAabFA9s5QsJhhdwS7avV1F/7oFYEM3gMh3vqWec
pDjScTrUtb1d83CdmJyT9LnompeGQEX+VtICRbnmTGvKcmMK2EJE7DhHSK++gwhq
du/pvUHzR7TH0NWjpcKcIUlWWlE0m+5LQMCsxEuz+jMnKHdr4wgMNBabx+rkWHEA
MHG8TiTKiUoPO3uf9ojHzFirbJ3dwxu9PHHRbEIYeg0I2JNpLMMdBk8o4UVhc5xP
LN+Q/dbKRGZQkQVS3IIK5Hg2SmSf7D8Z+xYalRjKR7xz6Ek34KTEe9ipVtGCzIVd
zh+roRPcMutdfMq9vr9eOj3L/b3eYeQz3/Ug0G8BFecUMYDs3yZva5YViweuAyIH
xWhWHCnYV7XQ8sBdsvUJ6MW6SWLyHi2hOUcTftX/XALjeUpCKo1FeEyEbQh/Mtpb
TiIJqFN0sbs1Q7MVg5DyPp8aGwg8pa2xafN0kyN/RVI2FB/kW82GGNVmFfiJOEsH
52o3kX7JZ9HECpVUlZVRz+ueBgBsX4WxBzU+AGdLTHFN3l03ChcF9ClS92Dos0v0
ISMGN0vVEoE9eGK2tWbo3qfLpamZCHmHmUuaAsr3LSOZDQg2UNM+cBmWMEMMqStE
`protect END_PROTECTED
