`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZLLCPFsaJy9awL1KGVEAuMEBMPhcjZBiBsKacuzvRyneSNTi/9PiqCvgMkvIlE6b
z85Wr2c8JP+EkB0O1lF+V9VIh32s8EOpUM2ABZu9CelmYMWpAqQXS7S/jEmwpl9G
vtNHntT2RjT1/JxIb6XodoRkpnIiIdNT2dzNSGSt4E0Y3k+dcrLzqDpC3HvJDyFA
+pZggPypkuvUYsy1mbENJhrAsrQIxqJtED+Q5ZEOWWBYpmZkHWDPVn/VEocC/uKr
jshYwbp+V6KaFbOqA93IE8WlMskib94sJhbIpiB3SlCyDMOC6JOVGt3LkByvJVF8
rNJiq29ZC4jnmvhp4ynG2cUCFhh7C9oSUfSQV25YEaR5xMP+b2Eqw3X6U31ZcRFt
UQH/UqXyYfN8K2KPzXWblA8C5wtdWlh/N/LPiGJ97i/Czj/+lqUmTwQu8SKVE+bm
plw+q7Vxj00BblWzX5j9Yw5+EQLmnzJnnsQe07ubgAxHR29A3InXtYcY9wSHGXm/
ODJ3KDGFj9rT17Y7LbBfbMoA335X/r0sr2mJkq1vD0GMrU1h5eah20XUnDqIJ3GQ
eRZybcL1WkV662TcrL9jnpVIvrXQ1j7nAdjO93gqWBR83Aq/k6re05/FL1PxFvpx
f7+RrxkO0/8mcZp88/XTcqIONWP5Q1CvYRyTX2PKv9PjnX1k0nplF1RBsmVPEoQG
JY7z2A8KEM9Go6c/C61SLEMs3HEHktfikQEdRjC7XllABFuyaf3Vn240OFXIpnkZ
Pj3txuD4oTwtETJNRD8B8mrf2e3VcLUeWvNq+Z7LdS9i7D2kTM39tVUknV89hZoI
1MPTAi9dzboHKVrIpPYYttQdn08VZ7AqFPjhLRJAhnbKNbNqns4dEQ6qWrylgRlT
ES9Zwom9Rym/T1o6AB4OhLKZ2cwdEIFihCHbVcruLayYkmVPorbIQwv0UXZV8t2g
AvUpXBRPn3U6LPLay0pixwg8dmAnCanvyWQH5VlBk/5EDvNlpZlT+ZCwHlDNBkd/
QgB8+UL3j4aYq+3xMHJP7G2qib1J0Nxhfqx+F+WTilnfQolc8qa339/kuv5mj47y
gO7XPkMI1P1u4X/bveXwpDRUDJitJw0+62gU8sYFHYGWbFT0vlW0o8zcv8xQ4yjS
3/o7ujOlc3oISizW5ek8S116g9psVoyd/8xVh+/XNCt5QKwrJUNDPLzvJR+mRMCi
8cKjnV740yKnDnpi8ymU4wBvyKHexKT+sc6YQLiBNctTdh1OkryUt3LjQbaUyKpK
MV8FkNFDF96eGoMsCEBCb9qNE7sy3r0WlZOeRB7kBobjy7MWDLPWn96jSbv8r+yn
jlTe5zKtFPgvhJ/M4wffVKMrMLnbW2HbvRgxtUgAINNCeZ1hW02KUCTh7mXQkzCi
K6tAdkWLRzzcb38kuxO0G15mtt2ilGNfUSYKVo2fpHXJRJKLUkVlFR2CaAN82rLO
sbrdWng68j38e80P7uOz6KZoldjHgh0OnFEvkSCgfvqb7umaNe9a3uYnk5Ii1Zfz
kd2HlUQnxZwmM5jVfj48AIUqUlk3eB00ppcaH1HtI1Ap5E5PDBEOiYyVfgClVGKR
J4+jdVXsrS82tE8Kk+qxIB5aVQovPoiOOLOt6T5wWgvRoEXvNltyXNHxumwkMAqR
H6vShbDAtBhJNpsZySRGn5bulc3+6lzws/ywFUgbBiMzHpbg+RoX03B2ivaMs3Dv
qLYoWx1OdbAgqXmTZoZ+PWWRkvAk6vw41bmCW0gQQaEZZmJfqPlfKBkTnyaOc1Sf
rGcLzfmMD5H1mJOGq3z5jWz7D+o5V7rrVpSA1heUlSWK5MgH0GD8S94kveLHsczQ
OkOPikyWm87JyZRjw0EYjWxB6N7ySkG7ej6Qd978xOjUN3SUe+kwAkluoL3D/Uj/
jn1ZXJnxaM6rfUXhsZ/Wjpwg35NwkcPfbODmW6NAZG2aLqnVGs3wnX15h0S3128F
iiVxwsLZSkZwqaHPS0qoRx4JuR0OFZ8PNBkN+tFLJEL6nCMHnMMh133A95cPMpHw
xqxIpZ9YPzg/ntkWPabSfA0hMMe2ScgRWrGtz/jgdtrNdt2LwprZ6gzTT5dRu3E2
PCILQhYUAL0eOBU4FRWictmOZZJGsL43EdxH4y1qOmlro+TgAnQCV8LI7LCGM9dx
KfiKidGtGnyZ4R8UNF89h5EBkfwQhLA2e3PgpvEDmTs=
`protect END_PROTECTED
