`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jh3JDAW22l398e6CDsOVwGeDFH22N8BtdrLsl+nJco15ikPFpLuNCKdvG733OuMG
y8tMqMVBHEEUbvkvMl447rfW37K9XcmJ+YNcfJz/aFxO2kzCzrf7lL999GJTqBI+
4zbn9voO9TNoVbomIYY5H/l4xXhIP0IOmUlh+zJ2WTAMK79nMZqqMI666TM/PJCI
eFdolj79FdXz9uqYxOTPpuqhaDTNHiSQl3ekPT3AqOS38DiL+IRFTi7cIKMGHHFO
UfG+5JL4l6srxTAMnSAYrMqJi4hO497UDkEqLoHcwr/0mv8g3x9dWrCmaG9tH/tG
784ZjlOfJkC9oSKbfy8ebcorN8xtNNkFgvsbQt4p6ynZtNBtPvuX2GJiHQNz6ubu
YVhG5ckZxkVxvqDJCrt38GsCRBSGLqdb3vj4wk9K7GVw8NIAp2z29UcTIYk678O1
TI8cbFenTgVX7sqPQeOsnzKZf6l1u51u9PC06QH4r4o0XgqoYt5xY0pmk0y+jQKY
lwU165Z+PKK550haMRwf3EygTINY4zFcwB07yrt8nI/1YnW4pjVfPehuNhc0PFV0
4WBJUEHI58wSKfv0x9EbVioD28Bzqgy/vymXtxc4yYowxCvVPk4eFpD1X4TdFCpS
hBOs4fDEYIX6BLS/QRZNGLcypAxLz0f5Rl5+4X/ye+TGS/nOOZ6NnAqVONstWG+m
zJQgz4kaAxN4fR17YE5In3AIb4D6ZMS4qhH/QU4mD+QbIGF9syJfMVbCXjgHK/zh
ItPTpYcenze1P8mDv6iz0tcAxuK6l4MPvnblzI8kFxx9YFRbVujPrMNeEty6bH2X
dvaBurFweF+exPVXI4GHzEfNOLSYKeMEAIU7RPtcwDH0RVMkI5zwgRR17mSdb34W
hpwgS4Va1gFg8rTSsVURC8NBGc6n2JV0m2L68mCBQkydqcm77iswQw6mmVdIJNcr
Q/xPzDAxgJyT7dD5ysXARW+fCk8kMyOZ+WSwy1NvB2sjRAt3fGh+0bKRAHzHG2Rt
GEjN04Em8Vba9lLLVqncLziH3ZKw7m0uLHGK4QVED7EvIoptq3kLF0SnVbnhJliA
ny4MQA5SgN3SYxJYZIWdTPWqFdRwyBAIiq0484tPzgMYF80U/NRTxEyaNMP2b6fR
qjnXxjzA2LEMMVR3xP9cW9TnFtZMjzNu29eygiBvy4xCY0ES8YGfOPK5TSB74dqD
xw1Dbg5e5n3/cCYx/TK3hf4IhdvKHSrzlQt7hECrHLRoZKZJoe4ZxQvmNoMKW66T
NZry5NZGQ1OgBQYOjylIOEhBopWhFR9H+eHoIlHi6roVa/EYP4S4RfZhUgR87Is1
TXJuIxe220OOjbDukFFjBTWLnAYW44QIG/GZrBGcmLZsPa2O1R+PJPnxRtWhMz8j
6mNiWSfPjOOUrI85ZEdz10m6FoWVlKbh6sZLKIrSh4lKNDO4xONOr0jQ5Qe/rT6y
JeQMh7aghEAFCPyoCMfZACk7MYY/uIu3aSvKqMLOojtnjqYEz7+akHsitUpdzFdr
UUETGiO2W+pevk/iDhk0y6qqH1CAU+pPpUFxdW/eSVR3KvkvX8e2FjM4s12nibqT
Ai9zL1N/uFcwV3QnTmRvzKdUgd0PW3PwI/2FVSTa780FKDItkG2HbqW3yvGfgzLV
Wg/xCLK6hpynz+2IFWzjxo6cAZpHrzclpxzFq0uiTfs8ySl94rS1vU6rdvVnTL5j
ZET9vrsh7pXTUSNTERFJGGFwtE1K/DbOa74wSc+onZ8RNTTeeE0Nvny1+dfMbEuj
gdlgG9xuYxVb7vt/jjO/pkVP2VNf4zh+g+ozHhti0t9Gs9wx44pOdKCKaMEtZDnA
5J10fI+pmvNRgeJ9fkwXjs8Xnxmh0ePtWsDbyrSfHIDlSX+9qJBiPuvhdNJVZhzQ
s9VQTYSPrX8kR0wSdvbK3oMaDVK8+HBahePjwHWF8fG+kYCh0lSvr3Us+Q47AUdP
3PVsitFUyujbemF18jP2qhB9WRR6YB9IOrxDNxm0Hgn0mky4lfhuXKyCFwB2sPW9
DmOk0ONUMvmTt89fytGPvtq4DMaWErYXpJgDtC12cWTsprXJuX5nbEKGpMiVWovi
xc0uF55lrVDG3HSI1OWioUfrG9+Q3PH2d2wIm14fzd1Y/70M16tUkPKCUzfq8CdL
xzzIIGzEpRGnEzJOOPMrp2tv5a88fn83pCPkuVcKubBQ7qX+5nWUGgNKoXer+OLs
Nxsf8IGHntWaYB4H2CFrWxB3Ppk4yRQsqMlVNuW1DWsxw2QCjxahy6jRJmD9p6fk
MyWA8fZRGz62H0lgx2+oxloiRIa12NyFmGCtK6L5SnwhF9Mc50j/YmPA9wKOPpv2
n5Yfh217FZ4I4dZiHVpOjQATrrLKI0rmeCQgqnWfsn8QO/nL2TvPlRs+dsTmEYy3
01aYFaYHhgO9NJ8cE4qXQQ==
`protect END_PROTECTED
