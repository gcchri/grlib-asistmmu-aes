`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t6Aj7CaXvZNa/auwjX9GncS+GvtjxMlBm7WznNFZ+VmfLn36vEnenvo+hf+uUIdo
M/0lJ+21Ek1a7QhvRpPlSG1nJCpU/AP9J9YU/eILaY5O7PC2yB/Uyibx33wOI7Mp
3J0p8cSLsk9e7vXGecJ1xldK9E60h0BeYgZ2eaAxsSTEoT6Ch8y4eVarm4AuL42S
42GVTLCOrdQKh1UpzShwsmj1gjlhYHwQaldQsDLYMlKHIYIqt/7b5ylKZgrmF7DB
0X/3YJdlCZ98GxjBWJNOrZZhdSWcwTCGZZnK1nW9uVTaAHrK2jvYCDbOupITulcu
Z9bWqocb8S2QGhNjTorayqbHeZMMh5/55M2WehXG855waSgk1UEEpNhCxuzYV906
8Mel8XPl1nJ/8qUAlQc82DBDdCKhWwg2UkGIOOQ/McGbhCtBuoP0EN6+qj7qc/SV
ahGGgOrghHHFUUTtr3SKzg9jEw2jUQZcg58TIxz7JMPLPlYNic5O+oM3L4hCcT38
ka6jCvX8xX1Op0W9kOAG3cQQKPGIr9tNRY5oUtxE5CK3j99ftxWg5fvd938su54p
CM6PC2QgH+w2jAiWSSAidQufDzBDyBsdzjW8jZ3ktmVNJa2VaVo0W4eqXyLQ78go
ElSsc/AWpXsrIqQNIJqyICiXAVxquhv7WFFtRxg3730sXKNjf/suJNqlZf4VzaxV
sOipOIxuQQ7uMOn+gsfbKehCqM6PIq+v9zV9UMtGCtoj8K5sHJnI49o83MmMwxC6
iEtlNt8bYRUJFJq5yd3Z0gwtDD8pOuiB1zTTYaDxzt3qnea1o/HuxVA6fCrhzZgF
aAKvxnNY4OknrFH6csLzF0J4xqoEl4A6UXER1pq5z4XANJ/I0Rap/9KFlGTeqOzK
8Vj2nr7BysRo8SUgJMkA3FnHfnrUfiSMNEtPl9KHR849Ggu4qPGkvqq8qCGGnSzt
uj0j/pU2WGLPFAtJX2clDvfxTlOwrfs9NEyZ1npzalqes00D5CXcPi1q58bvrpg+
V542mjdHsFd/ywuMqyHOtxVhqMJO/N9ye7wirszcRkljDaQsLKsn4WNPjk34FshA
f9XCcnY55WP61hlCnVjjZReOWm2bqv7Jh4O6EH9C4sc9r+3+rgajO0qmaRiDnG70
K6aljF/NCaYbZnXbareMEU6MeylT+/rCeFOj70JgV3/meo053d3O8TyxIxf0c0Va
qvjc1KYKGoNrj0cQbfCFtzkuEv9RVP9PxneIDFpkS5Je/lWhn2SnAcl58z4km3O2
/xSiXuE3yoYWircfOED71xN4weiGoiI8fHYZ/OmDZ/0ElYPNQZMd+CyTupdDHzwd
MEgrvPsCYF+nWgLAMF5rLA9TA90gNA8TIicpkVf/N38=
`protect END_PROTECTED
