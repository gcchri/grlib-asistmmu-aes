`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZmSTo1kHvp+SaER9KKbA33t0j1QF8sb5w260NPCur0w/Y/qT/XtJm1KPhyiVA6d
A55R3J5Nwszn9sBRnqr/jnk28e5OWyG89W0zsO0/WttVB1TjT1iNxMPWrpVEOiqo
zIks7tqon0QQMyUhFHwBlBEc9SxU+8TZFt7YK+IwvG5a+qinP17TEHsAk5Ss/7MF
PoWycCmPCNtRz1iTggzDUTgYsu4s8sJJ3C7IlZOXGh/go+sMWHV+W366WUNNPybn
38lQ/SZA7UcYcPjsnQb+zsAinm1N+emFaGQjzQvMKr6OU9L32/iy8geASfnHgvGV
9XDBLs3WERlu83XniLNSiPkxsdlEsSQrkLhBla8Cd/4xKAnupOdPUC6zEfKMLHH4
Qrx4f2ePljhgPTBtgYPN+cxZZzxF166Ywi+Wd1Qd7Ctm4kWQf/d74VnzftANqVKV
3eeEzL/PkI3y4YAXMqUH+39F2RX55leVGuJMjaa8u/XKW8cPpnhxF6735YhETbhN
bfr0WC7oCGDSHm9RcYiudchmgYw8rBEgxxT2/r+S5aY7L3xT+KV+mhjL/0bXE6zX
eeQDaNV2g3yhh9vxJL5wu3P37vIf4L5DjoBDDL4/+Bbd4MmuhlWvapN01grZNze9
hkEwcioSdWFh9ZT/FYKsG6z8FoYuv/QGaTMlC7EeeS2M0Zs8thCZAy4QIDnuD+CB
q9mrvrnG5mPjwopyoqdsVlHxwnGW2fiFJB9tWpMTl7EIDHGRQUdC56yEgvZZePdg
j1qHgM1JgLSOrQq6y93W8qdJ23b6pCGtv2/50nNnsxQEiSunirYRfNFHslR5ODQC
z3Wjuj6XKZyF4eVRG/DfdY0ZLyBT1GuQ0PaqXk8HcX4UcnGTMiH3BL4CuYSp9PB1
G2COGdr7GvC+l9HYEaJjDM/yqe/lBQUL+S9kFbzjXaKcVzw/N4HVvIphTRB3mIlu
GXKNw/Vf4KMB6EimV8YKjI9qWw2375w+jBlJXANJEOPttLCXFqqsqy/c7dry8aad
J06UPMfFbEa+spmQYuanGq5OOhSjuQ3OeToTNmO0wrpHuy+cg35IWkcmigClyW7l
uScu5Yj6Thk8Lp5/KPg5A36dYdVcACm6Ljl2l83xBr/WvgEVwMPxKABIW/qKEKep
rMco5CTSNmQfUWL+d3eLfQ==
`protect END_PROTECTED
