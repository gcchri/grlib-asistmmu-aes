`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lECwhXa632JR7XqHV7Y26sxhJi0ogEzU4xCRG1Iu/pOPjPNxx5bLxsfrjaVnBBsZ
emFuaBn9nJAWIdWijKhVkLXgjfvHdm9+vGTGPyAFmOt3PWL1sq5MwGM6EMVTgUWZ
uYBsY1vepM82nCt5jm6O5gbZBS+lL2//SO6qWVBff3C9cKZ49ihmlhptSreAIkFG
7L+ios3G0DdhImPAivConNJOy+osovXEh0aOhxh4H/FQ6rx/FWtlH3uLBZe17OQz
TsSDabM1FEfCMWn090C4xD1Q2rtR6/69/q12dHTWCKLukEhYeqTyDyXOpzgWPC8X
nkYWue+4JcE25HF369f5Dus4LfUhwYB5HQUCQKqmx0LooK7yq6pUWXd/4S9mBOoM
`protect END_PROTECTED
