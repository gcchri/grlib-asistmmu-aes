`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+AY+ZPj1qlg1R04leDib2QpewEKLUuV5IKryiZb4Pb03ShMoE2bh/ZXnFCmHk9vk
BElaU7pH1KP1TkpPDrROEpJnHw2hJe94U4iXHgWftA4HX8pyAXe+Oj2QHthS9AHW
uewxG68nuB8Qj+sD7mmc4u7sieTqTBIw50fOnXZ1wL3Os7JL+wZCc8LZcch4V1OU
i75ACV2UbggCYbGBAaaIHSOTbk81NMetZzrHR9ZTKSsltpsN3cxXHhJUUnFO976Y
959lVQS5iB+/X0cz6x27Q47llo16fSw8hmzTsrQ65vOiFf/Rd4WxJpFkiDDysIM0
hhuFPJVF8fmekVejr7v30muBT9Vw9LHpMz13095isGJZZG+CcZr8EyXmHl/J3EhC
djzQrICzq6XX+mKKNpYeBsrPdGKnTZXkQ73OPmBpIWWQ8Ff5R3qPvKLihvp2hhSo
dRgau4A/EkWikaP/fd6dbkvJXx6yFDqO8lqiZ/lvkiW8wu/rDuBL72WmYs19RUj6
VY8nVvaovtw/jnw0XF3CTg==
`protect END_PROTECTED
