`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rdc2MDZE9MLEswAn/a/WjiH6yJQoR0hNp81LYGSFTNhL1ml5Ub9XcHB+en9sSxic
aKQOVlVAhF8Cnz19RGK6I1BkKSs6NJoJtAOGuSLTUnphDzFtHGhpOcnj5EoSJBod
SniCs3Mstru8dfqUdKz1RE+Vx1kVxpf64a8HLI6v0TrCPdiG+hFlCNEIdO5CQl/k
d7sWAcBqCUv6Cw4G7VYnV3pfu4foRUk4bjGidtvp263McCj/cqUu0DfThDLxAbMR
+Fj5woBx87eBx56HO64BT/Z/oamo39n9uOS6XUITo9MTqProWh5frR6qLtq2Mp4q
fdTgXrpmZcUT3zYeOxW3rnFD55mML+SFhxcDbbjeR0OZ+S4OlYrsKhECd9A3058j
tM6RAItSQh5cgOjP7YHcMxR/ARU03m9x3NZuPzcoyGBArEjIxYbfnO/i8r2kswR4
MZWVXSiexNwZPrVwddeeo3OuAu3teHg6WVIs4EQtTMyfm31KH3nxAjTAjDv7mPnP
R6WQ/r+oHxe6DUXPe3AeleaJLFmroVT4451tcQKRGucHUcxkswyV3Miv7sHvanE0
o3RcbZLY0qbPVkJSkV7BGx8rP5qJH2wXLuRPr3B3cqPwuh+2pfplJmO2xO7NZGDV
2ykpZE3q6NVPVCKSVSxW/Xk7z8UUMdPaeIgvWiF5FD9k1BSQF1z7Xm1ViothiFE0
yyDTpJCLqcPqismfCCRGmjE9DpsAoHCASgmWgDFjzECYrS6k6LoyMX+apqA2uBK5
EXW1WaYCz73yc53gllM44QHOIfI3Xv0XNib9fOVHfsb+k0JxvXh41CEm2ydSD/2T
pMMZPiMO0gUMDPU8HZdrwlme+Z3RPMqf9AmM9LtBg3AaMeH5+bGNS7d2D5icVqwO
nvuugFIMIZ5+EYoZ7ZbnnlvdHSjjmfS8nHk3aUFXrVm2KpJknhD0kXVQchZG26cR
lwxeGq8jXgjXA/LaQa8WigvtY5eejwk+CmFAeqqarw11nwl0GDmUrelYiZroP8kS
6v4wnbL86lwKea/SZ++9EF/BSeT3p8Cz/Xzqg/mluiItCnpd1E5azGIUoFldHD/v
KinthNNGPN6yBVIWwX2FojelGPqIM4gR+FmqKNQGsTcB5gvH+94ZFLhz5+WXOBaq
8+Nfz99Wg/issXpr6UHcaWze2wXWbN/W3Z3PRWcf1iUORSG9l3nehXWC8U6npCLV
eRpbiP62lfGAeUSoKK91baGH04Tx01MxeOZNZhAQ74e65lVubaXmy7V7mrWE7N/C
G0o48bWV/3Sw5PVUTeU1ikIwCYzCEcSOctHJ/jo6BMH6vOsvk7UW6i0MRJo4n1a6
Hs+t5gTCCNa8P2ItTWRTwF+VIkCyyLgmg4zKrqjvBplDXzX+WBfe6fPh1UoZo3jl
I50vdrmCxdJnnGwkD3fwjGDiB+foShWCZKE4pq/Ggwn0yIiv/2QwLRNnxP4bH0iT
TYoqxAS/NZEN0/j1O30rwvmkiPY4uN326yYRLjHDVCZZtKlJrBPJFXYshdGSm7uj
PcAgfR/J2pMv1iZrZizUxTDk6Yn0I55suEzFeLBifsszAjQeluyyaPNObCImE/fi
`protect END_PROTECTED
