`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4yiiEz52LaefJRO9YG9zodEa7aCYm2e1YIWThuu3KCHqgHvRedFyNUY07yN2A5C
Ar1k0vMYpOAYJVRSKxknYJb/SqtPgv1fEv4hCqMhHEfUgo5/A/OPFNVldP9xLzoI
p5HtEsqU5f+xzeUFHYtnpthGsXyW0NaXAk4/TMLNRMLadQuPpgzUTdq16uaQaVvB
73A9l/UNnYttuhEl2fBP6h8VZcxnaOHQUHdxdr42eg7S3SsyYJR24pLgazMXOiKM
jqocTx6sEP54CiR0Ek/Wb8Ry2sxFKfVoOYGYhTpul4fRvgvoWETu9huw1ToCr9KB
Jt48ZMPLzdv72iOlzDI2K4wWOrdzpgQIE7IxNa1Z6BRLULEOiaDNgffKwKFxlq/y
rgsPi+zrzKcyBLGuCF+WHhgCKJBj4zzh+4oAg4OF+dJ1hMR2rd9f6re6utIYs8JC
25WYM/FXVkxxBbshvqbOj1V/V8VLef/QEc3BhFMBEBKM1mVX0AX9V6oOZn5iLeaU
izTkjPBLNhtkx0msUWV/K+dTTUV129p6V+A5ZLVYstVDj4tJKsNy4L9Ms718HfAO
vcrF9oWaakdH7ItT8kHTNA==
`protect END_PROTECTED
