`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3PrkKD3yU0KE92gNedil+HESaaUnNww4yCqM9iq/6HzckUQHNqnRX9+PViHcSs3A
Qu0ucX7W3gM/b4dslbIxvkvNWkOkUzu53wqXjiaBxeRXlmajfcL51XBHGvlLPdxR
wKwZ3zRYP53Y4bRH3IljffF+uKZ+Rg+LCqru1REn1bzrtOfSjK667KKb9MNahk/L
mk7QQG267kbXL2IVJGRAPrXXDHBO+WHcqmZo0JefAuRpXRoBGovpAOB8xAOzriGu
MsHb9kMRG5xpVAlErLsGTR/bMebJ2xv5GOpOy3DWRBE=
`protect END_PROTECTED
