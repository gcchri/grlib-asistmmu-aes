`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3rVtU0NJTBH1Tvcg8bgl3g3Vr53RCmiDifUm85lviRctMkIO3MNf3tEoHCMdixG
XQh6shwidBlAcev84vDDDvb54n1TriscW22J59FVh817+gUBXnj2GyTJteu6+Xl6
TUg5ejzmHXS0az2Zds+vyRhK/8QHpU5MTPU0PK3vhDcRR3RwO3RvLsgYLKyYVc9F
58JZmNbPz7ZHMb0u12q31xrqcDBFYJVsSKyArqJeqoQZAvGNI4hho6s+d8LIgSos
Xe+weZ5KWSBs2f5smNH1ZY6+c+GlPMXcHW7UeMGs9hP864NanhTNikOvYTKXfjhy
P0T2Knw/NqgohxlQQFI/NYmIEaXCRka6SEj6uPfgjR1WPE9tQJP7H6kYmx1nZMrq
T+SX+K8I6ec2F81i/HZfhRLbLfaK1bKJAfWF+zeEYiByvvQWr8SSmWxvwIa6eQa/
YDnXlXIdnH8+vzOMJTeCPTxFlO9gCVWtigh3Iqo32onftOtUKqobDqn4iexV7ZdD
IHINnLxOOocQpPeJUQy9u63bjKpGEeKA/zzBX8BeVFcJyR+wijXQD/P9ZGJRYHXi
wWlUm91zq5U0kMCVeNTNjRemoWl0aveHV4bBJSysCiZly1yyiFSD1pVGwY+VEkVg
iC8TrDIrbU9fX3XYWc8k5G5T1gSToo/0Bj8DmvtaqHA8gXfkM3YUJfJ/UYXP0W3O
9YCtgH1LhjvhY9mC4kH3f0/AyDRO9yV6anJEd/1GRnlEBTVyKrYLb5vfHaWm53xs
HDXL9G2AZRoBYKJm5wjTo1+lVfmKOM8kvcRc2AOjFTZqLhgGCDxHqbmbMPfy0TH1
8xkcngrBuzyDTKGAHx5W87AfsToanhhfGQlEisuE++KG+mpOX1l87NEG6OIJmC3Q
r/wtGIh5mMGsrHaduKJJcT/tI2CydeU0jy33s+hvhhsJX+KWd4spI6Y7rRp0LWjO
yqLVyUQN7qNR+t6NTaj9AWthVcMM+48B8JK5piITNjWm4dCalMMb4VeeYwFiEMN7
cSzLFt9HzH5FlUIoivORTjFwWTVgF63p/APWONjfpQgDS5+CN7J2wPNXVRhwhD6I
`protect END_PROTECTED
