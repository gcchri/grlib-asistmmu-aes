`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gKiHSFg854xMgynALyMEi9+IbzXV0BMVdGK89cDeWqzNcCaRAvvhGdoLZeqOeSM/
5KNxCh2rhwJqUUEM9I+SaemYaYh6L7N7S8Bay1G7b/uONQjDVQL25xO2Tr9DK3V2
jBKBgkHeOaWbnTZbZTeWza1+qDINYnrPY3YevBZfUs7aSYj3Ns+hynNXG66V0fAV
pUPrrV4zZfQJMU2qv2s3CjjFQl3yThy6rrJAybDCeASuU6DBX+e49+r1dG9FBJZB
SXOOmflTZQgWw0UIQym84YLt8LzMX3dwD+EUNm1AyoI2EfrXj+3wUBJoFoPuhNRK
awfvhzedZkpvNoYuJiQy1FqTnl4mluzlLbnOcoNV0Nd1HDXKsxOKqvagbJbK1VR5
wJUDsLsDv0md/BGbRN041YWVvZ2Zbo5fANRV+NvSmeP4orvwF4t7DpdckEZUtpDX
Mv8LG3UcUxH4LCMXldSWFGmbuNCaBJMKHxvD/maPZso2eNkW9M/J0zMVi6THOj9r
SY8k1VBDa+AlG+9eq7/20+Y80JeP2/zX1aImsWItL6DmRtbYWwus8cDcWbrk1e6H
zwtb9i+maaB3yrf5idmwQZ4YkooNGcGzba4IXvAJPTXPGaQ4fmuiKcQjv+6ouSYT
B0jjqwLV/Tp3lmAZY0xSzg==
`protect END_PROTECTED
