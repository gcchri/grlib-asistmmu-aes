`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bP8NlVtbtBQFojkz0gU8rRLxpRTrLaLgGIGt6QgF6Ma8/dPxyyw0kEEEkqlIvg24
LwT0pH3b8u1emqSJ4bKjpSiT3MeyRzic8TLDwI5LitiXXWcdlHIo0vrkmbQacMTE
N2zmBBs9kr/mI0M9+JITn8EKXbvEcQOhONhu0Nie3jkSC2l0PmXxxahdu9W0lr98
wZRcNIo0CQn6ia4w5dkaw5ehNgc+0G1dyUosDX8EKkNGh+c/HqGOGGwtcubwW6N5
mHwFqYv2fHTtTs2EnUfbJ+n8exFVoEKFK/HkohDDsPl5csQDlGd5jkQ6g7v2C3Nj
1J3hZosemYwRzi/EMdJamQeJfY2J30lsBQ2uFSxh4wgQlKXG6zj4b2rbN2UkmRfd
BlpkHutxHw6ihRARFHMBdaA8VQ32m0V2iyODFKS4eKwYc6NAnxxJH4zlZwH79U5f
`protect END_PROTECTED
