`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frFaH32jspiMwnpIEd3Qmfs9qsr1sueAY7MUkAMjDpVR7QMUpa6XKmAnAq4SIDzh
zzKkrHPQGNKhmjPUj/gCvsQy9oRYSWP2QGd4rrFp6fgQBgtM6OyObKrc/ktJl59B
1EMsNe3L3xOJytH4zfUA2rceStJMqY2UTtBVwrb4cKTD0bKZ4gm2RfbWOc6Wi7DQ
PPwRTHfJwKizgJbNOP/eK5yNM8vFTuPaoycOtTNgalAw48xynNa+HhT0bC8+JBv7
VJLenD5lwWSgSkNlt/8lQh5BvLY9yQWgjxEkAD3XKZmWlMalyCLAlN/qiqYIuvoS
A/aHjUWhi9GmJxf72boCPBo+coGQDbPUfAmP2AJmtNMLcC8KgYpTYCFWjseNefbg
LDUdYUlDgf7QIOt82+PKwdkgWRZWJlfso6FErOJXhZHBEGKvvO61eVlA63rl05Aa
YIlczDVOdtOZX9PPKdSpPJi775wdBbXcKmqukdxQI5Py1OuOAW7G6mCPFumIdxzw
qEbNR5c6hFST6f3IR/sN6hgcOiyGnsF5JBPB9ExP9sSXvhDxA1amQeFsjjC+D8ow
NheE7o0K1u+tRLjEnP36du+ND2tU1pbs9BCOxkKSu9hkWy7WQh1jM6eBsOSrjZzK
9lmVDPub1E2Zn0Bx11pzUg==
`protect END_PROTECTED
