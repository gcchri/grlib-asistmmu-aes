`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMELAcMFJrRwDtcUdTKPRMr9dDtj+oIP3h58AvgOIFWJNfjilSFSmZ5dL6kQPjur
ebwu+ixTKJOfMvSZo8GxtDqrWVAc0SQPh1AVg0tQJlJ02zXDzf8HLenCSTuP4Fhj
JSGEoO7rDQuKuIayByvJHOS+0FDBkfCNmwF29GKs+YS1CWySeI1r2OI1yhh9iYT7
bIP9SdPluoAfMKEpE/3WBgyThHii6zpwDwwmAQkQzeM1tp2bKmz2wnwGxeFqKftv
qMLa++vNUcB43i5MJsmPKD4VWRtMWWmINrlygknbDK4tKxjlkMjZVnBpZUxE2OoY
kjA0mVp/eF7Ew+vA/HOYj3MNXxKvj04S+HwsZhpt8Rkt+RrVoObCBZYmaQvb72xy
4330Ds30dxw3H2DRTo6xIqevaDMhdnNZ+NM6x/n7Dcp/w0GQ+hM1+AeFlAOAxdzk
nUMwOtvdJCcSy0+5kqsJPDxohzvzHyrw9b5HrQ7UWSjH3bzFyOgbUVxCXk0/lwmN
MN0Qy+UzElp5umRobg9nmEeO4S9o1VzVtsaFqpO6h5cUgkBWsnCnkVUlF7Cdk0xZ
aAuzNtwaEbW75nh56wt7b7NRP3pjI3Gl2My3b8FAUw/ix5VXHSmOxKSU3nj69ox5
/G9KKh5AFc7EP1tP04Yj4kcIWwgL4oaTLNpuS6q9yXkJf4LlvRr7KhIXaztzpkIx
qE0knwe93GOYocEzssS1fZJRBxOQPRTIiQtwFF7WBiUy8wmYH4rMBrmaQL0jyC0v
of/QA/F0lXGWkkuALGva6HPkvQaLhyNHbIMz611hPdeCgYxa+bYfZ13x8lc1RSc5
lggVzXgQgyoGbpe25pzWw/9qCIqNHry+1OU2nyQaxmTfrD80/axtp7Chz6AuSwSc
sgAbYMr4m8RulNTGBPtbApcpOgOL0ffQ6UFKXhxKZP4+Npq3J/v9GvrayoZems2v
10L6WKAXsT3LOBj/f3V7WD30jDZf9eCWHvjqBUbETeMZOA6HtGmZ/klQOBD3hgvl
XRQtE/ByzWBa3nEcQeSvYFx7uq1yKBnr7zNcdWrUvEYCdytDjdUiNDLbES3hErK7
cZyvNYJLLA8aNFWn/s9xM6BNRZPHOxiBU9pn4PyY2cajGlb8cvGSRm3xvFloj6hb
TLoyTvkydrc/MGYeHxWca/8THnEzWFkCjZMt4kRWokfwuR/vEPmRr/uws3kVM+UY
AyRBf71S691VEbheEVRr+nTqKosQws0H/4zi2SVMEqqXgOdMceHngBr6AZ2dp8Jl
RVlMXFRh13qxuycmrauucUcHyc61E4ibN75/rtKE7o3aY5TBvA1k3S1g/mOua8Wy
Ec+SxjsZlZTT6iOLO/8eJ7ZS3Oswtrrw29L2HVsFrpNkhDr5wxlZstvCm0yeIot8
8wf2SZdwGBtcO+IdoDvA9wX7ZsVkp656ppP6CkBhzOoImafhKNMlRijorPBCpdec
lDKSfBqzJB6zYCTuuIBEDhBXrLp3PTXcn57UmY27iPwh5LXystjg3vMSfHAw5YJi
pL7F+TB0OXDDjxBdoLNxGAc7R1OyjWz5YSzGf2pqxpIOP8DKGMmbeGsewKAQzrTL
0ZmMJA8qBgEec+zcI646SLfhgkVn6om6oa7IXxQLeTntryqO/PgFYJ6avdFsBNk6
Y6FwQJeLf+FmRNAKwtcEXdbb1BnkPkCI+ged67i85ZpYpNhagizvbihnFAj3aIky
pkVPpbur5VwLcqYBH5Ts7j1J/AT1NMOuitpD/M9Rk0KbIAaVTMaFQvEVrlvQEt8h
vx0IZE4ge9lo+tYXTM5b5FHJ35RJJm+2hiMHCtNghI1KdWILM7Y+zUvO6lWzY/bz
f1qrOlgnJsEOF4ftY6wxX+d0fy2zxo2e52tsMqle4tGWjTBrx8wGlCayFNYzkh7L
txOAiXV2/6cI7p0s8XWvs2ozsXmHeM1eJLczEzo4bM6bfcHIu92r0Mg2c4CUAQky
0aLWf/iWk2VgTc31wI/mCLZ8JSISWZhzzc8dDynfThyOIxttBEHnSmuPW2WCSLNi
DwFkUkdLg45qVIdBLXjdhaG6WLyuXRZjHwfyIG/dnr4uxhgXyr0otlzY9B+yHyvA
sNIpcsbNuIspxscGa7KYVvJgvhiBio6VPXMI02LNtKQrUCsu/eQhFqVaBSzENWqi
zRKXEFk335h1QEnoPSllViWjHnSwn/F3/mYxS+4O4YVCPHymHfZUKV8C1dhUAveG
kD4hIblmwT3liQGCJG0EBfbqe0Y/TaQZws0r+fD6p6ISDabtQgZ7y7MHqlca20iS
IhrKlcw2xcUNjsjwoU3kPjQhcR/+9vNdeyuwKUCDXIh3AKM+H37BBkd4sBD2QkXN
d2Z7+UBeuBCgw8kIHgTLSSpl7spAmAB1xsSal+P2VIlWNEhKtRvnRrhijplm3pUK
AqAGa7gJhhzgRcJ3PWQ3vWud3NVbwBzyvQuCnXigupnhb/Vzz1A5WGPw4HNz4+5X
5tAUBtDREB/ZlPjtvj8ik5EBd2z7q3wPr9/3wnpWOlaRZo8gi66xo58jAkUcd3dc
azxvVGoGiD/ieRi0zYGtTlZaIFCoP5V5xSBUr86/0IegmPCEXVtLrdp4w+3alDqC
zka3g+qghpLlTfzWFF33jcl0vFQ78BN+u/0ZpTA0ZTL+dm1Nfu89rwypW6WEIuft
vo3YwhGV9CJz4FqtWFdh5pu9aQuWwtJ67nfthvMzr6KJ4jejpI2vXiiBA2grWzC+
z88RNv5uawXWIKmVQkuYF5h3a6Kg5aft9wfIuE2JL8CjP8ckzFz04B4zM5DE6h1i
RlurV4F4FQskJJQIAl3dZVsdmolI3xt+ovX0NOxd1zah4D/ACuPMeQhKmx6prltz
H2cUTvvDjNHcU9Iapj/ittjn0t96Cr/pxs2xxt19UAyy80mZ8UwnKrtp2kDzRCUO
zbiqV/w1MqWkKAvkVmWI8o+ub1kuXzrIQtiNTbNqGS/IDv8yvjKQefeyavbMdohn
75D1BLL4It5GZ+hWQXkqyB3hIISjUQP6obR8p+zPjBCijqRPpjMonZv+nBt04dqY
sp+NSPMdFRt+fqZKk74eJgWS/kJYAmi7Ttgr/8rD8JNvB0D8kGwWWjC1i5LCa8Ax
mUbYKJzfMZ+8MFeKea8RBTuuMyxZfntV5kA/GaEc5jalbimiL+7a+pmf8bj3OTGT
FObpD7D0tk468ukSCK5k9FphPTQ8ZqJ4V+tHlBuXt5tZJ3W8fp/yqowwRC1wFi2l
e7/Eb6rRfNmBRy+4PbHeaPguBSryN54IfWbM+L2H4uW2UK3SpGpT3pN7L4BSt6zD
1ZuLYJW/y8AUlzr7HZu6wyW/bH4WbfyLe1Tzq8ubwtyc9cuSPanBfO4zy5I9ghfo
jXaArta+GahE48cBB/Q55wXStHGD0+4MdHhI0mh5D1oO+fHcJDpnO85iCwwYXDMV
VtL/OgU6WLzWgDZI65fmB64eu3qgDiTgrZ25reS23yO7KaUPf0G2vmPOBa45o08J
SiBtT33tf3dKFlUO59hfePdhFM5ApFQrCn2iZhqw+l6GMtQHz53MdlZplEbpt4LX
rQFdYNOLABj/rNJ7EhYUBOW6FvPODioRajKj2WwA/FMcsJejPc6L4EO7tdMEYN9Z
4t9U1RX/4DRiXlB3pEsjmjQpgdFCyrQfIu+vIq3xIRHaGgAYXFWiBLKoPl/R/TJg
rSHlnIYj1M7JEmI9DFGCEjBVojgVHZPhrfSO1gMnKxUoqwCgSp99gf/hBXUHqAGg
W4sxvIIJzITihZPhEAWjSxLqv0hLq9g5oC+9+RKVb+u2cxzCjLCnrDwFInbRlC8G
HCgqc9WuZWdU/DoOqjvUi3gnHv33KFaA2BT4wgdYQ2hB9ZtkHGBU7Mx2Nd0KhGs5
tY6gkv24g2+vQq9fzwPcsfJxBiZR11sXPL/dxv2CJ5VWu8aEYZVN+Box5G0SyUsO
W2+s9n5z9yTY1BvZmp+EHFlBtk56c1rMztUKLANQWgaKS8z2XRnmJvmlWTCUCuSj
WlefIZ2vj94Utvmkl5Hl9uAg7Ao3KtwqCJvrMK4WlT1mvxWTcaLXLmRhanyl+jBA
DpchwHEI/KsItYOR1juh0eGx2+PxSio72PFdDpCheFUrWUW+1nSVLhUoX5tFrHv0
kph9D/GMuIIX3a1p68Nd+M9AYA+fhpxNLXV6HmP8F7mm+REmODNX5vVv2LBJH4zx
LlAIRjD85whgJSUpmHPxCwP4mwyoDnGD50vuBbuk90FmTwkEG6bT0f7UGAwl6yRR
RIpbr18VwzVyrnWR8oyMUXsd7d8bb2wW5S81jPMdt9zjx7MlpAdHuwMxNDSDlzxY
UT+K4be0Q/EQFa0jfd3ZW/A4awwHII4vEswMv+/mQcR/nj01djki8Si1W3DoADiK
PhIb0ya8WK5i1GQTgQ3tRwhAgk6NbUPGSaTh9E9Ul0I+lZg94KB4ljsX4HjULdmR
5r28oFJOJF40zqw5viEwsp3X6/UAteKwH3jYLy4Fgb0Tj8VDtksqoA1SNpmAM6dB
ZBSfiBWLz0EOf+j81+E9QjigkKuFkHBxK9K3ntG1ebJkvmClmwMALPuR4/Sz1Uj3
PD8DYSV98uoFU1TjB51cdv9GwIlzFSlB8phjrajUwAGn4eby7Pj5EOSyoVMc5QuF
tAXyWytmnluuo6NaM7TDvebVI+k1IuAI1rLREPO9s/lRcGsb2Sn+BuL4hijbmAxL
yXrLhQlFcTS27TNtITeBNSbrGyohxHITT8B86K3+ftY/uFtsimS+CsS/EI+pS0QY
JrdIGrhCrH0aYhhidJjzIfXZun9YnlHeEgj89L4JS9xQbuQsbPjS/+3Ltz4Y6u5g
CdfpkBt4zTao8AImIbPUFKuCXfeVqh2bhfOKL2U7yQFhw+UgmW379Hc2oO4X4Mz8
I17G4wm/tp9C3bMS62Rw4XiYaIQdFQVBCedghBtMEAyUt7eVwGuc9slTykqplkTK
Y5XOBa2yjGX3yMRUFvRmTZPnhGdo69SLbitvz0orNAB31leMe7dj9mHmws17zrJY
SEQYWbMf2oP6H0z3IWq0S8zexXq0uN3nAq9qQoLsX1i8NX/PVSQ4g+jm2O77IFyO
fObW+6SAKJdxa4pG1hZwPtZU1bGTfb27JY67G4NZNVrO5Gzszfvte26s8lk9Pl4a
Z++EGQpO6kbBPba1pC5lt77Mt1ZC0b6483PGdzzmqQKQYiEeE0AlHlBYTk0KeczK
AqTYeWqWV8huS3gJCvmyTfIVGIIMhqPncEI2uyb60VdJxtl44HCE5ELprEtey2k3
Vn96gaKtRgI0+Jtezp7WX8vQGC7gO+VBJN45Ivs9oUPXFkzUr4nsZS/G7qinlufm
5gWks2lWdTpcYNOPY0bpOMB49YQj1zLEYNRDFAiWYJXCt6Ww35uOannvaz8M6hJ9
Oa+WdWKUjHi0SwpEOi6LEZPG7S5BtIvwALxyUMOFyVb879mefkxFIQYiTtuCXbHw
rXa2L+M2Mos/8gIrWYmlClG3KJKlqwc62TwT9xC2kZr/43k+JjFVyI3lLzIp8SFH
bB68GZKOQNtaOk4hT1FqpKoDfb71BIPDWNtqhhoEp+9rjErMHB8VTDMV0In2dtc4
yi5OrgvgYOZmxTnmGvKgvLOa8ArOH+E5sJF434AzpUTT2xeCNyqALzGYWwII0cFR
2r5zmfA1BQ7OMuUez+xj6WAB5Z+BH0CTAyDmnWVOzv92OMi3ClmjZVrP4KUr+fX1
HNN+zIUI2t0H2i7yUJ55BesiduPIM/UDHZxqWULMVgmckD7TJcZ71KbNSdsNe+de
nOre0iv2oSZKbezZq717ViOXUyYAKdy2VZ2+kJQEZJwRSEtg8rmpkuMiGBCYsYNs
jK5mhxZ07hITC3pNlDW7Lmzb4n5PnupOdV9Zwbu8Zhl2JmnynNJc0ito4FHIzEPE
PRmxU0dgHK3nF1kSlQhvwNQG1FNW374yJDPFj8eVhZQNR7j6iIhgp//VaCgI0FE5
7W/gXOodJEP83ZRwHzDOuKI+3Mb4m8FmIA7ZRVzb+LysFI8xW/bkwEgIgzZIKS+h
UdDxLo7CcrFoGUrFcGg34JdwrTtHZdUP8Utp3+LWboyoqZQexdg4gI5Gg5RulIxC
GAdXe+3s3GlZw+DXN0QY8D8eDo80Dq3zPBau0y+lryhxba9aXAPqtvfcC283ukFn
iKzS+lqpLIa37aHT1mnRw4FNdE/RHjYd8uTJ7NDmnRV8OB083aidQcyL35HObm25
hcyU8tMLHscz7VWB8CQ+1nLheNMdtFIUvKgGals2VoE05H0eHMHFBcICmgE5TAJW
ehOPltHjl5deaxMirdN9nXBCdVfj/6xN8VPap/RqQFguXXpT4ye4ArvgOyFZr3MX
Okn5pLKtcb0oMCFmF8ajHI1JzuLm5ijs/dM6/D9XNxMzzjvFAkJ5npcw1y/V/2sp
FLNx5e5rPuMlqv7Kvspr6UVE4qlX4hWYWDyRWlEDcHO7K8GHV3l3qf87MhKcEfG6
15hb7bWoEsBTqNGtT71PkC0TZVqoCB9p1GddisTHYyqgWiIafP77hXbdNxt/Ay1l
oWceWQN6X4c9q1wvNVUG96GKSgDYf1EIJB0l3WCJ/EfpcbETOheCjEN7rk/QuvHM
gF+q9fFpxkC68cfwMscEwwVv0sC+m6NOMKrTFXaJO4eUW24vMZ3FcMQWfWXW5G+K
rN2iR/FHtGijAjErPg6jrHkasPLJjd88SbMpSizsoLiSCXo3j3tYjPALhAH1FdYh
artjyQ2inn6risghBMSUsexerKoboul+5Q5SiWB0dWOKyyLkn+lP/YWhnr95OU4F
58GTqvwRCYEKf3qmaF3W5WhLGvK+GGpVN5gww6QLhbDrkqu1laWciwcmnduvrP9X
MSpZX/970c69gUf1vaD6PUwEQfiGYyVQamPV7oG6NChdLkTmjAD3DBhpJ7oI8SYf
Ee7zt30cDjbyoN/mStEc9uJYmXF4FIiv6ZawhpOBrxMaaSjwP2bSkR8j19nF2eRf
mrVADuHNglvrnwKGIl5UWKDsztywzRi1lYz/7At3dzgs7edR2VhycPOGnb1qMiAz
MI+r6PGjhKEEZvR5G72OHjA/Iuj26KEcLIYlBiwcZX1p7AXSI2o1SKEu3p3X78WS
OeR10/cplC6b+vrSf/NDPvOxuYHTzQiQXvs5f8GxvzPRAiN3fbLlexU/fh/DtyeN
6e8g7f8PpP6HT2a/rEXeFdwVS0qrNggHnlzQH8SXndRAKpjbDYQzHeRbdpLAOe1w
JQGuPzCWFtXiblZmllckeboGOPA7oPIDeSIHH5eZr9FxVZ2dsEN9ot4+Zmz9c0dC
WV/aTFUz5L8oaEQF6kyf+vWoTnuKVgeeL6cVYBVbMhRvCc+c9rbjRjz2J1+xYX9j
NYUH4J9Id5YMEK3E6KLLpAG6JtppAVltPjK9GbBBud6fsjDTeSmx4yvNoAxY9joL
FLKNeB1kYoYv4u0inpWKyXfrVyZx4BsSSn/ht2bnJDIPwz2b/p69k9Fjs0xDXk8M
i3Ho6zOE2hZlhxnDhZq3RSce2ucVwWPLZ/D1c3QhnJveXQS79YsWYQUKuF0kcfsx
gdAVgMHu3yhiw1u9DZ6zrO2GqpB4r1OBEc+aaxFRFpIYVTzthjOqSkbkhRtZj4ia
CiqfSkC73W3Hbo1Rjsx3eInh1+920iwTQZJERsCZ/pxywsOkyb2iuXIMZlVs398N
4/xGhWjqk1fp61kN9OWrBDSU5mxIx7k/9/4ysCI2s8MuP/nrxzaIFC0La7gPixw+
eaT1AEC64Taaxo4bndE8a3wukRegNjPZgWXCAxp+VXQReHL6jS8bgYj24pNDXwkT
KSIZWSrK0btFIl9RBRd+QIfwrXq9HWANhpc8/nJRIEHEcEFquXYasTz6C3EkIGp7
86Mdi/5G/1pwwol5s189aF7gcrAaOWCsFfBOyS28Ldz2POTON+A1deRhCb9JT3Nx
nd2crxLu8CBY3naqj7TJymrZKtv/Rf+MeMFQ9mBKwuOfrlFU3h1Jukikkd/7MuTC
PmOeMrdAmWMfLzohs9ScFfG0+epcpIJDa4qPQzByXGB+km2C+2oZrDbb6HVHhIbx
+f370JG85TxJdPzC/2EFgDeMPNWP3IB86zPLw8+KlLzkLiZ8ld7smTgVJqzytuF0
TkPTvvJP/Mf90E//sjrvm1+aEA0i4AXSJdMoXhXu743fzKc3pmNDf7ej3dS95F8h
3/eEfbQ+NnrelhvFRzMYIkvR+6paMRdVWJnxaqb8Dju/z49cJxjT36ZOhfvGDwKQ
7wpAMrrd+Zv38nm5bSCFcyYSkFG48C/tp9yV1P0R47XTkca7QmIkn/Aoov2Xz084
yRNH9DD1AzjAEk7WOdQTHkJDt/Yi0kwCPd1Df39OgXncQsxzIF3v4hEP2+CI+Cni
5wsDgwdkI0Ag9CTqBWJ1DICUxBbeGrBoj8wqwz43A60BJxNKDczpjROa5R9j9fNw
Oltqsy6lbVGhEycFZ0lisKKpvk3QOjMSrQ7cNgLz6TM47vE8Y1SG63PP1XtZ56Up
hLHoOdnaNZLgH/3qM/9xjoOeTjzXSwsYKCSfqm2pwvk5+NYTlLCxKLF9qrRjLvXs
vwMfuEQJUW6sSZmgz/AygdDhQgFWBC7YOMlkT5TJWbzce8Q63Gwx40FAatVWNnMX
ZeuF2i22znB2TsmMYz+D4aRunN4BnLKaoh2Gm8TW7YB1+QXAKJ2CLcFPUaYUHYPs
Rp3N9WjVy1a0FynWzMnnJf//3uPBy6iAT3mAYv+8iTmnDBQXuYPlZjTMkZu3gLSF
O4/tzRH3HwQtN1/8qo+y+SKy0jL6doP8/xtAL4uB8NqzPd8l2HQZDXDHyYtdLmJl
bDdojtTB+W9XRYNM57JmtZAK2S2uJ1Di9Nb42gtyBvSmbzUeKNS3EwnQAYZLFx3L
DFXu6INVKD+xI6ABR0rFg/t6pREVqvrpJRqvGTn9roUeknbc/I0X+Uct32gPuAOJ
5FASyo3PVoNrU/0V/shtWboeu6PLEK3pdqoWPpCJjtfKy2l/dPrsRw9w65O8hI26
LjDdEPRt2CcfFVtdbbwTmDPn6fJB0iAiW6umhPllBEHwfFGUQffNxQGzuA9ef8Rf
RQhczEtBsiiUintnXFHID16UiCY4kAIESr8JZXoPTv7FA6HAJTPAlfOE7TZY5ppz
62NW4TrkEBCmhf/Pnre/TEruiUG3bb3ENIewoq+ANs6HkfIheeWW++HOC2UYdLSA
CpadQ6ZiLn2qEc6wNkFtR83qXe0cOuhK3JbvCXSx6oy9BkCmqm5YPK5Ic/ScwKaU
u54XO2grIewe7TT22NrJNlIUuGWq8PGVJg6qK1R1YYch1tp2Fo5vgNWz9Pm0KhUk
lbf9Eu2eOZJ6LT3eEcGH3oGyUlVHolERCgyG25WBxu0UUjN//+9PM16q0PtbpkV8
0WhZZjTO3v/vx+NBhpNYZgFSNmLgLMRfthGS/hxYKATh8MfZRHM407aZeckbLqm2
gayBWJyMrXhKxzUtL29xXmiiKgOYdVXNl9cLGf9MJOVr5UYWddHViCZV4J4E/rGk
d1+B/LcWB3cki9uu99X1D1HDslWh8FUfTfPd10YFE+oaDhEFQdWIBELvKxYSW6lJ
/HWedotvdIYEf3kIhuKeRTSwGAJ94UBHSIhHTymD+rQj/HWKav2VnuLXOWx0z+E4
z0h9dxnV9XdHPku+adXNByMZKMofdFTKpVUdzHk5Xg+3Bgio2vZSjMQbNFm8Fyxt
q9nkge0zXOgm1uj2cLExuJXCv8OjIP+4Agi1U+06humJZkLuuyVxMapmMnqRVobm
3NOM/TBfp0L4h3xolCfkPBX0sdoZMVPgwmFwr37wUMy1a/655F63MIn3xpsmJP6B
59KoCVwcFLkOqBAiE1nmRSxjwuJzkDhRa8Je1P0pIQ5HZXLbSKXQDga9cqYQPeBd
9ZtQuid3/mjb2kTdk+ZeuDuyiNpChQEu2fm+qJpF/K8f2SUo30EGsKmD+lSJvuYz
WXXTb2kYCauYIImxMzBDE9bIXRSi/FAfqD4UE85Cgukb7jx+xu2zwM3WxsOeDtEU
w3FFqBQAUVlsFW/10p3OVPe+4+f/JNFynXMWobkkwZTqMRteTkPn3LxRCSg3fgRW
bSbkZ8Zh9mRnYMTYTGv4f7sm3JJ2t7O6ByN6T5lPYsvZkXhNo3TzXKnHrpqZQ9pC
PE0lkiN19orwYx2iaKUySH0HxApHSvyaaDVc3Ngt2/qvBWTZqEReVqaRMK2Y8fPR
yzb6K16kueR0TNCY6aZldaAotuJYe8hVLvWk4zcF+gMe0upNh+BjVcpvssfk2eu0
SdildHif/s1UVOe7u0CkI64bz4C4UTT5emMcf+c9Ja3uLlldkHGfPzdh7WQugDJ7
JU9IG9E+n+L/cZ0TfiG2XJ78KHaQzUK82wsWaCRBnrRXxXyhZpCC37FnTktK5uHF
R7p9o6cjw16fJV22E6IJF7AOrPjX+sveO1OoOV1qe6HK8ApkyuvdG3LHpZnpYZV6
r9i3OWS9RgrGaGF7VV4qu+uohvEbZFUX2FHxpXUpLiLiL7Q9cCHpm1A3IIjkPFQz
4ARr7bCdrQ01oFaN4R0BVKwgGfiEyJkMCDgpZhl3Z91H2zN5TM7Axxp+a2YkgLs3
F4x/XZscW/zeZB6Lq7xmsf2UibX3c/UR0FBtunhGMBRJ7YqeTfk/6R8fKBUU+P4m
4il/45beB/kGMoPEGQA4ctj9Ht7/wLo/+FN+NpEh0O3+bJ4407BvMeZYJmFf2oof
LSI4/YryqdZ/RKZOoQjCDPAU7On3TtWgQA3x7KK1Hgc0ydWV3/gVVNAmvhjDBRdr
Spl+VAlGIwnqvGjcoAu7lb/NOx6cbv9eRnuUvLHONUFNzH6buSlKAoC21tbrdW0E
ncQjbq3xo7FdKS1d/apjbUUY25TBxywESckZANcMkW1lcUO9MK2J4/65ku58mtpf
mzvgnnJahPlP52uWwqtE+csnTDZxuSfkIyK/2QLR2gbCV3rNvp6vNRyS1U7a32rk
Qgr1l0h2FV1FAX6PFeL2yAcHX2Loq63XvLe6YCiUVPPsnHVBvmW7fN2u+zDtqfpC
g5BtIQcddLhxp299F2GEBgKnqpuICC/1BhRI2YWm1qDe6efQyT40ih134s8cvqdm
I1WWSwy11Ku0BknitBMOR99VEnX5sLTnx5vEnmCIzbt92tNieoo7hJwDVpbWT/5m
SCRpcN6gBdZV/NydpCTUBgPEHmppKX9Dzhl+0On7zncFDZlq2P+i6Kp9aw1bCAWb
Co8OFH4LOp6vmsA5fypmxBMKsQi7UT94CRza51I0W3KmBTOXoyJIBp0r+wf8fAJh
AboONM3Mhy5BFtzB9L/2aAMu2IAIwmhlNS7MV8kKyvfbtwjJDjq1uMu0n3bOfXFe
9acAhFv2DmAOhnuK6GQC6RLL0dtd/4HztZZ0EMlcyzmjWaCUDwckz7G9HhDpeGfv
CSPXp/RPAlMX6KtOSS6ZYn9MMKg71owTklbbgtKU9hQH37KJHi/eRqXVAhxv7pr+
LiQTSMQNpMu1oiRazNLVkORhJWbXaaUHmylWeB6yio+iXtpLnA3j9Y4IGl/Q4JSl
93/fdo7Ol5Y+RR4PEO4bxUC6GFj47ESryvaPZKXb6iPPKJaTecU8oVexxnO/hwwo
Xxe7SgGkaY32bgV/rlG00/VpK8Cc1ieAIHlZhfGMtKLF5yzTSBuWKpJHF3Av9V9P
NR7BiZBEz2bWt0on32unAtYooLBUVUM+aIOWs9n3Nq773j1JvoLLgOYs8Zd/uqEP
6bJINq2mnC65ZJymIRxj7H/LYOAQxgIT25s/CYIET2yOcqLYT4dIqw4/s1G0a+2h
zCa4yujG+hQVssZIyuUoEuN3MENIFiRi0lU5+szJolW2iUkpo+PjCgn7BiJwGOfP
6U89vV420PNaC+z9TIsWX2RfaIuw4XxZ2uOEQ/q80QgZqVYqwLS7G1XzKBBvYtan
3NbDwdJk9kj/JbnoiTVL5dRb2ZPJzwS7nuLrQKPqMp7mRHrJqdNlxOioa5Ss02Hl
qskuQfUnOitN9mPjCq12URK+OWNrvl2pwMfmZlvm9+EhPnNbMxbkZ5/42H5N6f5L
Q9iuZLn3LwwdKQxl5+JsTq8XeBnJbOkzspIszE1/eRdKnhcGpDbSKLrHbPGKHrF2
Z5PmWlsUzG9BG69PWP9j7K/DxHuSKB/AaNGX89I3JX9ctecpu1RVf2ggG4TpJolA
AXyjG4uMM2XE96HtLnBv96Y85oj6IzKf5v0lWbW5B0JeOvH7+qE0pW3u7NATKwBH
IiD0IGZwpmkqyug6VYEZRO3bGkH2LNJqMyxvh9AYpT8NPKwEkHQVHHbfQkkcM+hb
74F1Bo6fDuCIaBvvQrhKm8Do3qjpeKNqR93tROLgznEYjJFpXd3EfEIn1XoRzeXn
+QZSfYCHSsbpJTKHYAUTnwAXl8R0+a1MfEyECFQpncR+zV5vUsJf4fOKHh9uyhuk
jVNtGV/CbKvPBcEu+iqK/59t4iLOf2St/HsRcJX5MXpYhrUlLSJ8JSL+R/cD9PGe
C+sWtVwYkYtu/21Oo4Pz42LM0UZtsmdwXWUQz19lemQ/VpmfftCq0OmAJiZ97ReF
za4Xp3TPyD0VJdAjgiBi9b7Dcb2jgcWaTX34ptwFDcjGq1Hq1M0nNSwA4TSNNxeK
u8Z56lyIMuZqZUTu6kUlt46SRPmkQ5e9Y+1mPHjvWiVtb5jfXI+Y7zsegAQZ5oka
DUQGBWCHPGcarx1j0BgG72BeI7E1ETmMPgEAfjJ+QCtYoNRjvcAbvDIIQqfrrf9X
GlYJgo05p5P2RloGfcvBF5MoodKlAXx1gx8hQgoOvu1MlgRiSb/soPKfptUmqlPo
67Bfvdrh6AEr9XpBIiytKEtvNM2yUECGkcgtD30Wc7Yc8UnrmM9cAGoDUlSG/9LM
JoIeoIfPuO+oCBJL3pfyRhxIR40B5z99fziGR/6lCbDfGhmOTI/sGeeY9aHVt1xt
zBboJKohgnlm5MOOMb6EqQwUWdIqTRn5by1JPUYN+hNghaURISgrQ5F17Gud8LHr
1K6+l8LZd08Y6+es+mVrwz65N3Hiz8M2UW1jx3315VZmK2mcwJptsYaGinnBuVJ8
Xy9JJ1VqqDaTIA1krlRoo5NjQ3YfA6IG9lHaYUW7oIZu3B09zmko1Qis/OK88tPP
Xdjm8oheBSenaslMXw1z28Hgq3abtAQs2ZlwHocCsLylqFCAT3isOGVFwSG2m4xY
TcehzslyboioM38ZcZO+QvcZwOZ/U2QkQZBuzi/g2ZkZphwslR+aXF6gkt6yyroi
gHu2g8V0NgOcdt/zTLSOAaeHh9zTz4VNu40e2Q7r+9FZ+4mjYhUYY60Ffk50PEV6
+srKKFwmDSQeiprMH9A1VgxwKuqTQkDLwvG+YjSALR2vxXyxQXNuzi+3TPh87T3s
CASdsN/f28xvYXFigU8gjjmpPNrBmDY8dgcYCgEDX7DPYeaL+EbsDtef6HwVILI5
VQX31/29+xWTqqSPTBMZI+Ep93pVWE4akZF3VxONS7b5VJApY/neGxO1u30VblaN
fTZ3bCXIaSd+8+rQNPL72y3P7njOME7VVTpA4m5BIQZ+bL8qv4DAGVKstN6cu1KL
OWCkswdT4HDndr0twGjwHdO6XWTvTlWrG5+oQ2MRQ4FWTKmg3tKWs/JrjZQKB9rc
4qxQCpxayKs6HIJP1FhW93G0iQxY9aCBAI/5i9JMBI2cFlDO59dzSy3p+Mo9zPj7
ak3Tf65XWUMN3bTzsNjZWAB3ExPMHpb1i+HzcQ8k3I5kJkdqFWj9Pxxr0HoBnh1Z
A8pCyL8ip9tO6Bk7DITkfxii5so1G+MzYJ6PeQYrElugB+B8V8IBGW9ENs9wnHmv
izcfO+4lEjyVcGIftT3ZeMTiwlx9Nk2Sfj8M3XTYSl/Ty59Q2QssNIhz4nNVBf/L
fBLspW31kyBYDPRsAQR4v2WuHIthrZqRgPLvRcf3TwvOJlsCsDgbKLN5evfOgEe/
yEY6rrNP8nb2M0WWe2djCdnAllVuCSHJCtXPRkFpvmEEGEY/Qe7YcmF8NaZ1wzCe
UbMZE8J/VJiULxG9A/FnS+nfcDp2pBzpYHnQVdCKVib1LSNSOB2/u0iQp8IjmfpR
VcTRwIp0Os0kyoiXVqbTfzWkDbTxBTRXJVZ0FrKXUfEi7m4C/iF7pZSyOWUo+a35
LG9wvMeCdWn/g8qFP5xOZ2WC3Cgbp72CKXhFVkvcOUWxFb/ayNvcnMMNZymAoHcY
XOxVfp21GEBqSAJSkr3RGWFlQTCpYYvI98kAFjMOgbEE7rH12Obx+Px8wrUElZ2M
kXRt8RTrVWC4RmhpG3c6yRR/Uj4HXTyzM0+N6wQkuqrvhBkaTqS+NqzYXy76W19k
ZXBB1eU9myXQbUlmzfl4t7j4PpQFh8XEg+ijK1dX5MKk7Xv9RTRX3lhn3H/W/hF+
xI2r3RR0uCoxR/Y1jqCysvlQVwQvE9NJZGe2BqEzLiOHRdXNyyVdj8jtpiBTVFjh
0u24K86zWl36DNrp4rdQU/uU0WUdVMiCvIrwqNUwXgX6hKlPvaknnM3hm1Ls9k2v
RlEeiXfyAkvLOJDwaa5hQvXxWa4KQh5c9JGE3ux0Q5/rTDK4Gghi4FRLbBg93dZ9
uE3WwDvpf1BbrvAjgXucPJD1kR/bVXcHl1zXTtUs9nszxvcSpfv5ish1Yi9+NgvO
l93LuZxDvtyLw6vm3K1CTJ+a76HZmw3xe/GX6b0SOD6alAm/U5f48QB25jlyOJNf
DWwo0l4H8Bo8fNn71YECiuyCfud9oEU0XKf+qpFmgjMcmiFe+0j6V9f1VczPlaaB
E79ubHSzNR0Z4tOXwAHi8qrsIu4ZVTwKLA3vQDfpsOfR1zTavAOeDHOuOh6i0JvM
tHvZeK1DJVUsEo1die9okvjwnFV3yOpk3W/limREBykANkl0x1utsL3niHkp7xB6
/guNLpQcG1Up+j2jyrQJc6WtlCeuayFOaqL6RT7u8hN7plRqi2KyVxv+T3rpVV2K
ky964U6gCI6p2nGkHyiG6rVF5WHsu+aTWXBzS2P294IQ0iZbt6l+rOf7WozRAZ7Q
JshvMrI12O0s61idsfcZSrv4SZSvL73j6GN0ySPJolgugr3KB0v36mn95fsE3HVM
RWadfVzcB8lAj8b9K19Fk3ecexnZv79lXP+/yhJcQhhySzBCt9eE/apadjSWAziq
4sODCHn+t+wY6L2jqgpW0yCfw+YC3uydcbULDyuKqPR+taMi6rgXWspZNac6d1t7
2c5/dvD0CNiU4MehWLetszrRlJ1h3WOA6jfkUfQtj0JSDsNdSecqFIBIj5oUExGt
2v66XoKkxtMgXJ7K33g/8uBNPf2LSe22/Ljk8pu5fVLfQTpRl1vZmlu3HCXIBjSb
EPEvoAx6wM/HgG5lUdparGqISJIw5TvrAF1qMsWlaGLm2OK+whAmqKGOcdigGI5x
z38r6mxmueFZgfd3W1Ui/vQgdAZYGRR2gLbbR624UYKdwKMMdQpHE+re0GOC4FcV
dDxNGFQPqqIY0l0wbqtEM4oR7Bu7GL1cgaePFVbcDUSgKBi9B4yWWuQFkzKPu2A0
fbuyzQbCDoWmlrD48jLJEVgTfv0zNAimM5L73478Md8cbyVyMAf1dx+sXohKAYFe
r+wjqEeYvAhmp09Yp7/3hqZPmeDJJh8sJ0S9g2ZvZLjKBeS3gKYZ44HCMa+V1sNf
5n9J5c1GfdUViLCqC9SyltO5VOFLYUzrXynAqrxaJ4fvJ3rBVn/iU1cHJCiw58DB
IpAEGwRUxP9E2RIgClO69B+pjZYtosPagxRC6OTGzVAcD+IpUodY74es5PsfpPdO
812O/3pMaPylhk9ucH+t9eYigFUb5uYBrnR1ra7x4ONgKirznD4RMdGmbnTYGsZC
RUy7oSZBtqcPdTzo/IhScXvXlOfrYoqMOtphq7nzbiHA+GPgNtIn3cAqK0PfHskb
qIGSSKsdyyZGlnxuj5asm0Qua1RcygXl5PFOAe+NsoUknM4JACBmQeqG6BoxVnh6
1NmAF6hd7zuMj/tYzhOYE15yTHY3jKrCzsIlPUTQGCMZxwWtuTdPjsoehE8TB1ot
LWqp9VSUV4MLlXaLuwdjVoCqu4RbBPgCNVXTQd6LxdIQUZIU0D9f7YEK2iPXlNAS
5cLtw9BUrjLwRTfGOrSUeWckfrGho9+7QkGll3x2DtmVW2koUBJmeiawdVTDHvmY
K6eQ5aq7BDyIHr0L8NdYzWh1gB4vIhYyoCAM+PKvFkPlzmuYIOMZ5m+mqFCN66X6
MuKNReZq2BbOoXHo6FBl7S/JyVwEukER9JB9MhnvXGyHE75TueI2XKZc1XELmiXD
ViwRtFNaQ6sJzGNHstLMMHx5hCX9gObXl2JDQCRF2216RTA+FEoTu5h29AKBClQQ
wp/2ZR0u7zpZJ1bykFl8YRig1fe2DnuthbS2AIQ79EaWd/oZ2mdYxX4ucf43XT5l
k67fFs6ec7sq4XudS5c8B8oHmtEVaEWwpvYWyiw0p2I6cuBv0l7iKUudP+C3k45/
xxhQnllUK1MbwtQn5NfKel8Wm7fPHltBgzd7UFUpPwSuEiq804aeLK+0NgYDTe7W
CTLMpYjcjL1ErTfzFv2f7SFvc/lVAvhluLuj0VvosyREsENHvTjsEskLqDZmFsbz
9+sKEwDWz0OVUwyyqGUSk9o2bRxKg1VyBePo+xw6QxDAiDanuBIGF6XFIble1hP7
OvxEJX4gC1bFmG4MUGOh5pT7he7WhUgPbnANU144HhH+3zXMZ9mXCX0LWoC4EAHu
64/fcJF6fCAr7IbmHjyyE/CmXnGUVNFa5hPrzynQ7BndOO/kkED+p8u5uo9rGJ9C
SaIXXVAvQFW7FoqNI6zTMbOEGqUO7NygYd7MneGAWKZ5lrgDtDV1at0FGyqitNrw
v4RAq31XYq1iO0jQ+piy04/N4fRScHTbuCxNCsFUZDGb6cA/Pbhx3Peo2ItB07Ou
+ZDu3zgXvz7mhKmsh3kAwh/qgYNrOjfn0CtmnKak616VsLbA+/POmdvWYcYs4RfH
BmrtA2jshJ83P4Je468TmGzSA07AJhFCD6CkLM3Y5SFn/cEWnjfEfWqoqhtdOioM
2FKs2Ei8adU74+gdXQW9yLQ5m/wB+DprdFbaDqFHa6lY4PmoInjJqDFoGbz0UyO3
MQRGM0rgwMi17zjyTCF93WaL1ws1j+JjkbhW+vXh9imwGRal2f6rd7mdHBJUjFdC
Ee6n3tYdG/uyHw4Ov3A1/+jkTa8vgghUQzORCqIhoqe4ZSq43rzNmErfR7Ys6d7f
foGNf3aQFHnK3lvvrVld0sgHodZ5AHjCSie9OPVgq/jzjUbESPayDKMRikk7z4AV
t9SFNv4mFId1tlmM80eWBEQwBWZ4+eqhHRsH35jFAE5ddVrFr0I0pRz3455PLYao
UD8kesLX1X5CqIt9MgBpjr1gH2a+3Sb1C1eerTRSyiwPsimIpHt5kFzUdWjCKt5k
PcdYvdvr4ViuKWeHq00TILKYxjMLMFcgEh9pBMWo4gmj44b6FqE1UIQ5DdS8ND5V
ML+OCPajiexGcDWQioULMUCKTx/i1ifGKCVMpZ9RSUhI5fST8g3x9oxlqdSfDpeW
GbXopMhqPbxDmTUflQyA7iJ7aBi4TLj0tTFHqjRMAI62IL4vi1P8ftDsylPUz/+9
2hL64JLtN59GByHN1ymBBJUol+9SZ0dj+WBUzUHB4ZGPgEz6H5RHlpVM7Kx+pPzn
K9oeEK04kczg0vO/rVy5zlrIPx3JlRMQCREgGm3/sPmNJdmytJS3GBDJT+aNF08V
9+ejUe1UYCLiXjUt3XVEtjH9IY3MJ8BbPl0Jz9Znow9zgFpMugD6Qrdqtti3ljgJ
FmSBsBD2HkBWld9EbmQjh2IblTxX2Fhwviy7KBZnxP7OCGf8UXNz2JzzDUBd1n4+
WSdSOQICoiLwdB7WEnbaRLpAyzn5Qp16bHSq2YCW5QKcN8KaRttd6cujYDDeTpaE
y8z5Fw4bpOyCf9temV9xf4xuMmpQnyhrTjMGg2fCJp04sdhHT0//rQPxTZ3SxJQe
9XbXctUM4F/9joEe5hf4NeyLpgvAoYl0c3VdWNO0BdI/sdGAumRmyC/8tHV4LLRz
O3CoimczAaJqGvBn/cVy8WeGnuQHlwKJlfGwg+ldPTJx82Ume8jsDPjdElpG/AKW
NgWfHnt8Ysi5avO0x1d/6AtuYLfBj+ttuogaetc4WU1ByYHE5IJ8IUMQn+Dgue05
Zd2YFLmxR7EwJtE20yQb9RViKmbRG+wCqUzFypV5kMVerwuKO66l6zwX/oFRjw0y
GArhMkvRmvQIMaxCGtWFPWiBnK7GLSkHdhoFIPD8IxGsgODd7eKXoVDu/04LBLiL
pWUOH9FN2dIRCj6lFZO5sdp/T3zIUsJZ2UA09zcn3ir4Q6DGcvWHSPAWj1ud6Ldr
QDyNzItAXFJkGqGdb4NRHmIQinqltJXuuzfblqm42CHRaone6UTDDJKfgS1InB9o
CEpGYZhusJJdd7euh4ffMqIA8u49iPWQ4kcy40wygZpiXsiz//REj+NADk4g5RIq
3JqkRVhC+V3sSabVYv8QkpuNvf4Iu0gqEu8g5GSuY5QJ631gE8rOxar4HOxByTVH
VUt3sy4/ACavs2E6xsm7g6VrV9GZKU7gMGHcvDsiC/ZYqbdbD9hV27Zraq2bLZli
7bXeDBmsdwzu4Gi1kFOxT4Lnk30QVA5jDlnTNWCSq/WUD1+8u6pRihFeduqZ35Vs
1tL0IfAbKl9SAqweCSDQ64H4a7U9jjpIRa0mWWQMBUIzPuT4ia5bxPDLsG4V096G
1cqFNrp/zwWG4Yw+3JkVNdgLe39PaKE3T3Lp6e/B0vRH7FLISRFizktZe/rVauxw
+oiL/d7Q3Eh4fX6mbUmt4k0SiCa78i6GFUjpXLiUSOouykN8ycObeZzJ6UUg5vnv
UHAn7QW9rQNSipgF5kh1VgZUUWBa1vW1WrLvots/eaieZ1/5oXJjYYMxuBL3SSXw
i0kzELEYcwe0YWQGPkkSxfaVscbFKENjTuRRd43Ea5hNAGBdqnv9Hl//o8D1aaUd
iBIaoyUBM6SPv6fL4ixfiVEpdX9h446C/xAXcwg2zqGBQ5nUz5wH3vKj2QrRhlaB
GM1IUXImLbu9IDjF3LViwUEyR2YCw2kQB1ChsFLBtatAFpodQJFVrZgTWQneQpSa
zNj7MVOvSO1Dy29HFTpGSihbwjZ3SGPvuVKZGPvj5Fq0kSD/p0iuAfDDypUtQ2ny
onx/4DNHNhzvdf8hCgtARqHMc1v2CxRmrCdlALHfUaulNcNKJlnKXOmQ1x28Yj9G
2kseJXdath36RfqWfCe5iKJT2g/OlGe9C42VZSc0NInY6D/F5sOrfci1/XGw1Rwh
y5yDJEbT9zvN5H5eM/9HHdHxvhnQ9c6ClpZZ905IPBr7oz+uPNqxSjuD9+Mpb2pV
nldh0umO2z6NEWxhjF9yl2pOMmoq0Zkwbv+m/PYXAgwBNlzd6YQzoOTnDNOnFJq7
NjlHR+UIpAmAH/NJEb+fg2qxI9iYp8nUAHxRTEF1O0MOottiXnzyawcnRDfw3/G/
aNwLe2GU/cWdytve/DNbKOkNwCojJA2iaroIt0EngBMgsbPgH4s9twtas3nIQFwh
DVsASksndueZQgEwH51wyMnizmTJEXhVNav0ZAxzv/XBncknMnk+3Ix83/SeiRiE
R9F/VS14k65714ZRbyJ5TZ+KWQyyryA+HEgZkuJWVesCUsVdgkg+XojjG/ysgObo
syWyPVVq1cZacjofA+MS17X9MUNZ300pWINxncSvbdXvH81ejPDiEjZNdsNxjL4s
DBiNOQYRUKnjmGhPH/4uTtit97yR/0ueh5tmyincwjsuzxn/OpTlcvvNz4DEUx1O
jDNiMIY7bUXbk0GKyh+djIFEoBtpXECzm/lB7YUZyPIyy3H12Q3z6+zTU5VdOlI4
fAW6tMPhysoKk4SlaHEtlE+cdHeDyOM1KJoRg5kT5DWyIDCEQRkDOCHfcaH9XguI
PhUMm4tHAJgYjtKGbbLBuk2XqkS9M4WmcsalhWJMiRzoF/vutoFznrf1P4fpNZ7o
yrJsqZ+VdaK6bUJDAJx3J/kXCv4sEKydz2bDJNW/H2s115KrnYtPls/GZFtJlgG0
fjscfWOEDAYEwCItVNviwGy/dkplG9ie9xI/jS//Ja+qFW6IR4Y1BLsrpt6+7W2U
d0Nhf7j5E4kfKuw8Q1eAl9BPJJetFg3CX+RVpRrBLKfWlviggNddYhJ7LRaDg0e5
gteHqqSjsViBCazxI2dAeqWvVJEIOH9kei3zSAUrXwf8ikEuLC2uYZlX/dHpMOXB
Xc7MJ+5dwxaVAbw3q6eEtYd2el4oh/zODTkChw8pgFOTvfSecX4yA8VIVTf8uzEP
RlJ5LlqNpEs31F6ppUYT3cc0ezvGGwR5ZTywZmE4qvnzgCmHtKDr8/L6CmUizV2y
RVssQRXoOZQoTyTeDx70RS3ld3EvcrKxaER474smBCwpTLgSGG3VDSLltmU5MJdi
aHlaxsPpxOWEjcdGMo8K2Fd8X2w2MWML7OUAHcbTdZph8QS9GdkP2e19WOH8VPfJ
dDNutuTcfvetofBs1THHqcnl+FY6Ne2cRn/yW5zcihcib8uLFX+AJUptXNd8shjV
92TcCPqHqwKh1VsV8jC3+4FiWT2yrj45LHKEDyKUgCzABFGzGnAQJFzxDRrGFPxl
BRn3vwkFnguyIcOkfIeUcBx+PHWyikVgxhsrq0nWIdWqGMIITwrFgF54Se4lK86l
noC93Eeb6LxbohsUlpBuzXNtF39gFknQZQ93GXCCuAaYSyj8j/MxX5R5+EHvaF5z
wdQL5+wXIsJ1MNprgUVI9b9zkgbSTzk0Yb/B+8naHmRxX1P5Bej5+uIBUgZbiWE7
/QZoVB8xmqwqUDQlELxGYPsvJxO+vvcpf3pq329nUCgFe1KmjoHcZK07cItOGs9I
Gv1RG1h1AveqJVL43VQhr3xdKPxwxToCPMrMcWYwsW+vk03sNXD9Gx0BbHU0m+OV
9DFnDf1OI6gb77Li5sTDwUUPJm4jVm3TZXv6xmcGuv73vL3CnpUGnqGh1emdaNzg
oimni1wyYqNFrAetYdZLlpNpX7M+RaQv2+UWkXkZNhsNKSXic0TiIlFnx/hWgh/S
bR1q63co8VO3dWQP4IaGHLKqr4okCqhXtOEOkQtXYi2IskljFOIYa8I+7PTkyuMZ
Ock4eXo7J2oNgUizFqB/rVIjETKBLPyAIUgLoeSA0M68eYdXjgXiDV2yyhwRVe3+
V/3/OVknu6dE7BeqjktRurI5UF9cmOiDKh+bsfUgDal4tBCQIzue+Q+hwbKtz9cm
e5zIfO0pyCCH1nhjdL3uI+qEB7rUlrYkWwxN/LbsDdruGnN9PuGgmiZ4bw9j9hm+
cIiA1lB2qxe0YnoEXglfDQv9hfD/MukIIpZdovI0E/cxuec8KpMUWA1ju3TbEHOn
OvswuzuyXwJyTjh5jgoiwkaBy8tSMinOaNVIETY+AFZGJ61xLIw6lbe+hSmgWsCo
WSqGdqdV7HwbJRuCTrESkqWVg32JrRVRS1rOVAiSbgjdLHIhr255+INJ1ZntHatl
K6/8E+mMu1qg0Ho5c+010zTKnsmksv1S09dgp1vduZ09L48FCCoJLIv2ESFuja3K
ko/Mkd+6jXTrspWX4ABTmhSCjYfE0iulGTypXO7+0dcr53fw9BRW9LKGsWNP4qtn
99x2GqfYCcqu9nDWCroY73q+cO3fTNH6fKNLdODIKaXKmwVPn7/S93K7eCpwPLCD
ZLz3RdC0HglvQzuCa67tORImBu/RwETiYiGuBNHz8V1R7fybsrMwDAKFVAbj4VGl
VC4pVxlswftdWfTtjzs9jR5KpsjKJ1r6l9W3l0zjvBT5BtbV8hwsDnaXeybUupSS
Xc9rZYfaT66VA89+m6xkOq/HO3MjUJrwlZ2+Kfsj9tOynzxfTBHcbjNEUCCWMUDg
NpnSBHKJE/SAh7wTp8O7yUyKTdLb4lMDa5E0WMPmIRdKXLGI1OVQfRaSXAczKshn
i87P10GsJ5BsAJXrxwCAiVK0VaeippEWicaqSgqUG0meXbkzNflXy8mrxUlRTWbW
BNJZ+72yxNv1ze+NPBzOfzXWl3MMHC5LmgsbmkU30a2bRAEdjlrp0Zac9uiPzpWI
NYP3ct5llCvZ5g6K1I7N1Oro+YoEsHIvZpuU+fopGFRn9EzIFXbPupxR0HQ7a6As
2shZf9hMZOW2xnKwknJklO3ms3wT0j3e0Pm0iErQtsG1HMCQUI8zokQVCfFEEA1o
7rhuTvNiroW24H/xVT304aG5ed42h0vhz4wcR1BBzDMFET+lLiHfj3y3jyW5+Nb7
5hMzYHlBFffZK4s5IkJI1oLTlp94hYnd21HnfkFaq4feI/SAu2+qLEvauQh1DvHy
QaOyqdfjeX0SYKDWspbZT09vVl2uyYcQ1CH02YSq303+z1WfGKeABaiCxyA+roEG
eHR9Se9oUWAeNjocGpupoQRTBkn+or9KOZtDN8ScJEnfEkqxzlA3ugdqHUXz1Lgx
/e2CYZ+pE3Y4fcsvTUrDQKxlqRESO1KQKHlQZhrHAZ6DA7Pk618v8HVxg9CUKvI+
zcOivSdXr8cGKMjZueLFQqXQP8C7eos+SIby27nb6A1MRCdwF8tuHMgqfdeQCL4H
9e/GYjQX4z1LNmlbXK+3IklTGzsk15+e0JiIJ1jBwWze+ZgIQ0Ez/fWQOXnJaRGU
63HvcTiZ4HxUtlAo8tbppdn4zeNoNx5X7BymBaefWYC9ix66BNESpOJxgJ6vTEqI
ucx6O7bmeKVuX6yy6EhoPEcrSITuBWejlTbhO5XFaKmKzsxXEnWi2qdRWLV509l8
ZXOIv3GxZFBal9puAOn72mGUoMATxsdF+SNPfcwu7jcWKh6ADrNPAeoa508a+/Ur
N65AYkyG+4exnhnCmCx8GFGOmn+tA6vZs5+Gk2NvoQABScYYjSilHY1SDjuVSfWd
EYa4dRs70MOWkMCv7Ev06CIq3tBvmxdCwZAs3OUUH8Whw8+QL08YbJ/Cbwc+d+cw
ng9h0mYRwWHE4dNZM7F/a5U1iFXAEh4nORkmCjRZN8Miwsy5gnSIFjF9H/xgPJTO
4CTi7kCtdu2A88Z8vD7cf03kPK8iuQAclyNN/LS9Jsuh3Xv0je8b6OLzRrQttrAV
h5VPVHgxZauWNxf6cTxrha30fh+HfcnUATYYgZrY801N2kIfP1MX3Z0cxQF5Nsdk
TGI6E6UtT/wwLke7O62kd/33MpfEoqAMZcacE/UTpkr8ZZViZQZWE56PNwQF483i
iP5qTFIr9S5ZCBDNFsIZL4Buq6h3/qkJAKeOAiGCSfmx/PDOVjSfnE9yi0Fqj2Lk
hYEm/jSrvu3t7ja+b1Ooey0pCc/fTS/PRWRAo7YAmSoqW7oTaYSYl8bbRiclw7IL
BSwT+Wed9pU9/BKuisXtkyGpJMjMWLiYC1NqI+in4OZoOY25sC6clegw8GNQLOz4
jSv2tQ8dr0zUjqXYvyjXKNGV7CGVuncE8qOofx0D6v412wUn0XJNHGPJlVe8Issf
IG+hD9A/Vdua3ZxUu+4Qe0SqJ58zyXv3X3eYlh8Xx7iJ2x3z2SunAVmNrmRsFr1f
woesHQq9paSUoDPhouFJSQ1bEWZJ3ZO0dfOvg9ZKc7pxmiWmPCtz//ZH8/d6NFKA
IXtUGDsz7lZhXcW2x4PIFkI4dP8+F0lFqWVju+D/INEm4xgq9Wt8YWYkySKmbsGv
+QyKB+b6gotuw98Tp5Rw137hrtOr+LExOP0QmM5YmGX+5ZW3ItFTRqJCYZ+IZ3e9
YAVLcDUoHSHc+UP4IcVpJYG7iAODpMHtopQ4uZxAvcGOSxr1sC6+4sEt64t28Iim
oaUeusiVBcv2OOz/roD8uYVvQliujWpBDqwljMdo+SvqoZemgP1YTXzm+B2CFyE8
KpqBd1N4l+IXNJ8/j3RRrwac6Gf4AUcpsxDhddcgkaQ6egsQrq2D8KihGpfbXOYk
bxLyUl7QGjY8EjiQEt3Jf7aVCGV9Xy/gr6X0J/b+eWndRnkrK0ybmwdWJLWPCGiF
xTZ44f6zFBPcfrnlIOR5RId/NTuA3ApX4AqGdrewbk00zcFMgmudhy5ZeduWRQUZ
LQYW4Cy2j+XdkyxcZvJxsV2hPF7+YEnOjoi6JlOCIk5m3LEwXZR3ukpbV1DL8TbE
jAejNnZj4NIX5jQE3sxBQwKGj+DyTvZ44LDITQg4lRoZItJC/am2Wh96YsKdet1P
W0OjYFmr2nlGuSq3ougZ7SSfl/zbKw03aubiHCqHDZMsIdkiY7EOB8vq+Uj6IUkv
FZ9e3xHQqbnPtyPApe0HRqbVHV7oSrU/auh5pvl6f+Db0Yv0+fMmeCdwAiAphWB1
72uiqJZnWCtO6DT9K98RcIgGExLxTvoyuefNlwyWkeogU08gCYOVZMQA5EYfWZXP
GDL/VtmGzDxQ5lrLo3obXKHpoO/Z4E/mrgmQq7scCHCqvsVSKZQjrfg1+RIxFy4B
UPMUBT+8fasywjrZkArxeH+RIRH7E/lxX3h5VmfXv+aNQXZPyLnk1fpunMhlFNuJ
mPMLfteYS/5PUB2tO+V2lGNesmEIzfNflWLXfMu+IcLTe1MiKMiGIUXoTQogUdK8
cO760GNAzqq7mJ/eXhbypiIVEIMks2ZkC1ZUOssnYluJmimpFng1XI0Rglq7pfd7
RILO8A2XSwQEy8UKFHsn34RfAIuXWMhV5aiUWjlbJ/13nzerPy4pUw3rM3xIGdNG
TBbzdGR1jwIUeC8GyZhZ3BvNXwN49qOVaW9dT6fy4yGMtRbDwsFxCOBml40OMJjh
ymsbby2EBrtyph2LHYYNZl8N4DVKPzPslFBlBlh1C7PGK5qb/ytSSatfSsLWpnIm
Wbz4DW/0Ss0PJRnul5VrKq59HAE/2EZJBqmnb8s6jmOf4jYmm/94ljsPlNR7sjdd
JrdsRLVx/da9VAU3yWXoFcWeOJbomt5YfBlgTXyEGgR8tseqLlaHIx7oumu7Uk6E
2zxicSDWZDtqM8wIZ6fsWby3Nrw3EDZ0jKHLzzW6VkeIaWCK8rbkH5cJu/gePO/s
JV6Iy2S/eC1Yatnqw4ho5NJkMvP3dbfBSrwpGytD8wGhaG2nrxyk8ssj/qRL6ZLB
pn2zPkuuacdyzVmdDqQ/FvRWKeTlVCOy3tN4HUMmuNxHLOGWPFVvk2GDSghH9+W/
Bhl2N/BiBg63WnDjdnH0QaF51PuR8bC/8zsiWrufAicGhF1lGbC4t71YIDN7H5PV
94+LEesScYKGXrQHCqtDcvxP13zNVy/X2CfEyYv53ne31Y/HCQAfZqghIlFZn1W5
AzzOFZ9fmH/E+fSbkLGa+P0k8/dodBuuuQm3BE2z+9UDXdvSdS41hgsX5hm0LMIQ
ZXafTDNmDM9QKKWblhdh9wC/zik7WbNaxS8vXOkyKyVjvOmYAeNpNnAGI89BwRf2
Dv2onZRfpNAm3yPvqQY4ElsCZVz+E/WPgQJ7nymN6B0JWGAo0VSpmWRf+sIyTPS3
fHbPHbcksPx4eo+212pEf9Ey5j65cTQhe5F3n0nsmuF7eILHMhvQC7ad4E2xc+0P
Z+Q8K8iJ+b3mR/Yy6C3vI7Fh6bkIktx5ydg6Hr/gQRwv6ZMxPXzkiiknLOL2HdYm
iOFFEpGhwmK3TuGV0iQbpdTrVlJAp7/+bVAUAN450Rjma7p6xMXYAwjAxnRxpr6Q
TXla1GndjqPfLFGikBVdwIhR3IvejC5EXKUK9Ei0/lw8zTWXrZf304ouh4AOBmPD
60KwcNxNXH1XLNxODJS+yhtnz5BsMunI4f1Gp1DG94U0OvYjk5FktGd3TLYFxUeP
Ftl9hCd6kgP/WbpKZqPHyJ2YvxY3q0zzqoBkFcfoUil8dYpr4t79FxV2HowsA62W
joTZfGIh/MAJCKzxQa5Irh6rMJP5PpA+ZR8xavE7FQfFIGNVIuSUMpLgpexH7+sj
AGOLfeZYWcl2gXOcTCxpmoiLV+3jWU8j3uuZVOw+0bWj5nikGZrUucXuE5JSV2hQ
rTxiCjHK1nu8C3is1guxRrh287egTEXkmZPWnjgnnMgeNQNP7Z+jNfYdYw2GCyj6
ryTF3WafSC+s3UT7s8duy/8cvsSlLbl2O/Vwm0tBtvSvd1baphhObl+FtPybDR6i
9Mn5bEMTNZ8sWycnQxT1ZuqquAeFZSK+oaJ2amVzEUl+fZPdL4DCKKnVh6ILwIsR
aPMvx0/osdOtjh2VZPOFEyNx6OHgLXVK11D+pyXXQ2PXJUUfCw5zw0/E92ahqyxU
/enc6n2O8vsagycHMAVKsuXb+RgKS9f0t21zh3kNIUjlAAL8mO7Qn5+FO8+lrPeg
GJsCQh4Bynm9mlWjjtWCvpr8QrY9+1kkmGfi8+jMuRb6ZMoQ4ExqsCK66Rr/IjTP
GbvkjRNwuHtJgcD3yce/bAVXYSioIOpeVL1oUYoyy+6ehUSemSdz6thAt5/VG8X0
1mJAxlwHIU3VYzzz2mzeJOWGbh2Gkk2yf4HFfBFfsyw9m1n/qD6RXWZqyE02Ufgn
KEa1n4egMm7rVSZ7jI16rdhlaQLTZuE0A2UWBfbOjpdvTK0bxiD1rZDXEApE2Wjf
1JzFRG8g1WQGggjMBU3hH/o+05kWH9fqnNrsTHWgdv9xCLOj/K/2x3OYxcXXDRYl
/5GVQp/iVLxLVNG2NAwzqt2kIcHTMLhx2xBTjmmc6pQsdy8mekAxrpiyGxXnTU80
aecVQaZGv2ShZ4wbnL/7KlLtpq+BzS7AS7D9j6PneVhhDATyP3KqmqZrwVh8ufNt
Yzti/sbpsNZl5RGofxv8h5pjwVKTdjgUEEfgrC2Lj4ZJYMQxOJvJ/1MUVdeZNlNg
uPahaTp2hcvbk4ABNNRiFIXxGe5W+vvZX4WZ9ehmlhzIh+YaKlstilL/SA1MGUcQ
rhhprJjVeDePBC6pSyoZUyx5Ul75Tj0+5v6f9HKJtaISEbxXYgcth1DYh3iOEjj+
dwSUKLPhTZGm9dELSHc3V9X971G2lvmG0VFbRZxc63Jau/Er46qvc11nwqdwS1Wi
/1hbtQV0x3iVPtFdYtOb5WgDeWeGGuA9NCIFgq1COh1CIYog4qTrvPt/FKzHlxio
9AlKSd6znfhUM7its9eN+4H7vSOkst8ulgnj2ezMf7dQHMMvG76TlxJht0ctfD1a
HztuZcuWvn0d6Q5ARCTcW4RdgcLF5ml7Xv/XH8gsSXEFQvSzNACIeIeqFvgZpKKC
3CoEnS7l8I5CKfuVonaVphnpsV053XUcq7Z1SzZw1LvwQiJxDyU33dUm/GYJaivC
IWfj0wBsDQ4czhR9j7KUK7hHhIXq4WlxSuDh6hBXYjgTS6LN+SNjP7Z2Vpc6CLNA
VEQxn3MHKf1gejo/Y5Cnk/jUYo0Pg6sDgVfiDW8iq9/f3BaBz5KIwg3MG/4FhcWU
1Ht/VOI5351SPj9JQQOBIBEzvtaOFA0HwhedquJX52eHLdbNeUIadAz1Ygtr/Hkp
OpwhomoVv0kXIP2r4YbSwUwspWBmDPJVkGEODhXZrzsrR+Q6nqHAMAiybYWH8N2C
2yqV24HobHY69UDRet/ylpFTDZoXalQXk/PpzDC8N3LRtAkdk24HYqhGsIdIk+PE
2WTkB9Tb6spvm8ZTeaTPq3WAc6nYhKV0Y1He9zJwM6wfbTz42gJR/noAlgOTQIAb
bDGCb0tvua+I/MLtdQjaTLzD4LcWQ224A04sM4li0CQyWs/fy/AagZ666AvXa8sz
7Tbc5khDzgh7ZhI+R7T+sj4phckFWh9j9DLrrQlhP225fVLM/lOBZWyTSON+qsib
P2QDeDDaKYEBKGN0Oq0kjbHyU7dms0nOXoMI+lTqxl4TqXqYY8ckhlXk0gUnAxqD
93Z8OvGMFwM8W7hSJToencQsfeCWSmmR+3thgihiiN9OyND5PAhWmBsSiIPB3lau
Vci1U1BqQgGP5Yik0NDyemQYM+7y7OaEbtluyV3a3Lqd93q8OA3A6S9/bly5Wsyk
qJXic+jpbeimcnge/KQuuOOHYRPysJzBwJuCmjlEtk6a5eBKzRsbb8bvArjTLBCM
CJBsn0HiBiJMaPpYUSU5K1rqjA+I3SwEQ8bRsmaAJAUSE2L9qmPVaEPg2OVEIQKE
pRGKQ6AbWApT2o2+b2Cob5yFjMLlBOfZA4Cjl7HJGGtUUsZBcC4wI3AkaHv6ve7T
G/YC8zvbbEwrP7in8lilFDZ+ert3yckSn0tCpISkI39PejgMwrvFh0wzj5+5oba0
UVpDUxsLmVRMo6G/AVkDXTvUWXrvbZkh0C/7ytv0BbexIUWKd5LBFY3YVHWTjhd9
ZzrUaEGbYjckdaW8ZYlN28yliwGopza8bcJtT6WDJIYgqyrK2I3i58nvlciAes/G
DIM2WSqquBWfhlvxBLO4RAZ2RkQbaqpeG9LVHsA8fTNeTjD04RsVdLCk1WE8ibI2
yRnsdg21SPWsmTFJcM1pydKGAkYQYoYPeu1ydmvU3TkfpM9dv2NrsaFRXvimqwBp
mrPZhJ6thh3ENEKaXQd8Cw/GhlFNr9IOtG71zMDkkbjDH+pLS5XOxEZ4/ajx6KUS
2tQ0/T9EquOXM62Ld6hvho15rektDFAc9p6Z6UVO+eeUBYlnk6b7l9iUtm1M1nwu
QAnoxcjGqtlkYiy68fHOl0WDouKdGjAKkGxCWlrdiMydEfcPxm0WRmy//jmUs501
IkiFo6c+gqHhgnEm3bpP+FQO5xv5M3ITkDKlX6UpfYBD+pLUAc4qkWF09zq9g16X
HSQY3AWcdhUunazoWIgsH8dNBXh3N0L3vvEjN0nP2kiiQEYW5exL0EvWW7KpClS5
G4M3rRwFLkWOEreiohX4OhEqBpmSkN2B+jG1jud3gNmTJimRwDfNfGwQKE0e4f3e
KepuUsLDDPv8zXVr9P/iNGyHizmVqFD0f+CMOAa4xf8NtlFQQq3t2py0PWaSW011
2kOqN6nwkWp2JLEeEYu7rftrGaLteeSsFb+VdJEVvvgWbpoxLKGnRbzRVl99UjUq
2DXAEr3eBKeZ+I8DNnnTXGVnbARyH0rE9P6kilwNlNYNio1ahq4jBkoZ4aBRlDqh
Ggi7Ghkkp4maNM+ZSZv50q/Fudis9C0gT/vr0HRZUZNz/YQhsRT2G29Iu6YwAiEv
K4tZEh0rYaMOHmJBTt1X1q3ILS5S6g1o53EZ169PgeoorBqi07Tb4joB+gi9gaxT
Fy81PMVriLl2M919pFlScVOAW/COU3mhZ2X4EyTxiKXMkZ7qT/w9mN9VamAbTyWj
yciK9VIbxjgxzPyIskRfaMGk2OQQiCVBGMAU7mkTW12K3IJWNrUa/jO2QJhVf6rF
zVk4AqTNQvrKrtwfkeQdXIJbf6lWII1cLvdSPpZvdNRGvPjKfCFftHyUwD0LkPez
nQUccTh9jdh5pvstA4f/rPUffLSta3OIs2wbg4vCxhpANz7N9MpKK2XxK5UwFXX6
m7jSKMBkNqRVUs+T2q2oGyfzmLK0GObLjzFCkdu8oHFoI3I0VTYXvNAkFkqhPg8+
C77STv3uoP1I7pswfFYXxZkSfuTVaS6fqLvWVyw4fH7waoUcHU236uP58J638iXu
zLYNB22dRIS39nwOaXYCAtSqW/uyzUmqDT0bIe7Z8kMrnSHZW+9XDEZOMt267A6l
EuPi1l9CQj3w43k6AUTSM+ONKRZ2xUcjTuFr4j8FUe6q8y70a8TBdkbfa/5iRFy3
sUME6i7DlAxw6TKKd2TuB+0EJkmw4tVD4YLUOkIWrtvpnxNxGyMXVNouKwq5P+Wg
9uyAMz7EYVTr3Z5JqIW/kMmp009B9I9CLN4nZUDdG84W6NnAtYDBwP+UHPRRrxn1
C+JkmxdK3cceGhem1GhkgoNKmBcA5I0EfW2lphYyE8SeTcQbKMZPnJuTzEwBdewT
SZ1Pus45i6i2dWgM/hzZoldJvs25z6GNLnUYPYc1dUFIlvLfDliKZfkTzFSb/e8M
8C0wdH7kTg6CITt7SgnWwS7bCGziZVfLtDogJTWEEFP1wDHDM7wTOIx53mZWvbku
Pc5nU3/pmThe9DdlMCfPN8xRU93+IlD3Vw3qWwBqRNdj6UfGXhCAInoaMNrp5r7p
dXoD32RtZvtbh126xQXN338ZqwFIlTVz/gFjMUS+9O+TecC/iAAk+mRNjn3lsZsx
iZr08BiyDVak0p4R1YA/Mr7iV6yqeJ+kqkby9H7MkL1uae3YmJek7JG9fJ8UVhxA
3OhobEjH4qozy4H8UUhzOi/0ZyPFiCRbBDnA6NyLNmF5eFWWUuEpCbo1FawcpV8T
Ol0PNeOFnMGLUHfTwVbjgHYuaC2c/s1T+1VWDe/QGqGu1TlXZ6iyAd/DONCL0W6T
kyP5FNmgtu8KVTnXSXXQFH0L+OWeXIfdzGFjwnHAer0HGLpYc4cCJWSfByW6IfgK
B0UWKDgtXxRzxskhcl4hi4G/cyBZs3VxE+QAqjAgy3ZHSYdEasui5uPGh1zD4VD9
2ErmqHSh+BWhHBx3P54PVHkEdvD6JolGXmhoxTthKOEf7wg/r4nrRL1xd1L3Eper
NhCSc0RzkeWrm1IHWhFizOvqSdNzWFiqiLcnDzkYhbn+GVBfd7g/wa3JZOafh1WT
O/YzYvYsFyY9bgRb+qArRjZe2ypx877/Fqw/gyZJzks+9KEvFs3frNqU2csRohUq
bVGbX0bFJnz8KUWnFshcZZjFUCbO906xg/ypDcfdVxo390lCzlbCpmc2YYEMwFeP
R6mAEI+mpHzKAS8jIuE9SJ4TQ5dsITXacSQHX9c/QQaCtqa5euKPQHucqvvQVWKX
wwhevs3rUr2193vrzQ5hfXKZ9uff6N/62r1K6mKONQrn4AsVQzhB7F7y7FDlnrmg
YVxuKqBFpEtHtShXdKKhiXbzbEpmRen1c0YSSjoiWPzLPMzuJYSXzsUAO/9igulJ
W0kW2xbwgB+pCM6yfHHlDCa7Ro8KZOKOneX5h1YVk47uLVVdthYw6331eNdEDYjU
g12c/vU5TppYMk8CRTFv0ESCVHwJmVrEW50Evc93+PKc05XW8Cl9hE1FT2eoUldi
k8kPQPi2EPQhsvHSGLNJ4sUdPaxh0l4Bk0DcHflhiqWhK+ePfSFXVEf5nkMRn8hb
yQzJYgoXDHsg4mrgZpXWbuc9n0qiAvaZXpWqySP6VTV+UNm7m2omaGp98e+fJqj4
kSv5bpZN+OPYXRYt7tugPAPdEYXBoAUZmrZK9yrnRYmQYOvY/pwjRuB3YhTFqGtw
tMh8hJbOAE3nComKlO74pycTj1b+b4zJecIgdRDcVgX4Y1U0X07xpVvynT1D/H3x
H32/VW4jdCjxrNcCgMGXbZfN1LpEO1hGzUDgGNHkxx33+DA80M1FLkG47VnAp9ny
pxwu4ZAe+CPguYB1EH9aXfVP8YQgZ05QM+54nj5bLuebiL+2NnCpt3wzBDShYib/
aGi4nkeRJXqb/egfrignzF5ix1v79w/Ny3gj8l97M6zi5TIPZQlLARhCygQZxBel
MYQC/EA0KQMoKvA72V2QCosOaVdqDiEESJJEzMB6OojUhogGwA26rcx11lMhn1Oo
yW0wfyZFlMpklPwcJ/jmGp8iG9rwiUal1Po4G1WUmoPJJtOwlIPiwHUmaNMgnHu8
iPjq/zDODR9fC3surdZawWpe8YE8zj6nmRkAOI9DRTvYDqQIbOQg6r/aXBkLWkFo
oJodnTjaiareL3X7LiSyWPO/S9UbdfOOhb3QQzETwEKwXRZOL9cY0/yIo4B1BzE3
Dip/5VO2RwFMhFozmH/hJwfHHGO4cBSN9gaRkffRp5HR79wgh9NQwSn8GqcMHEKw
y9tJbHe7GullYFfojpmi2VDkweaQjutcP2XLUvMzsm7hilbou2mNRnVR1D+dxxyo
Rr4Yhgph6EdTfEliJtRB6X72yBASLAQYV0rUpx19301JGa6PB4BK9+T2ls/V+YBt
GlJqbz03a6/iXymVfrqQGTxcTzNoPZsOiZSWGwH4yzDH39FV2SLAKr0NvI+jCvus
5G2vX9tNUuAdRGFl09cjvVVeZfY3SCiftlE4GtdMKZtjctPhwTRSvFgYV8baTRqy
07DjQnAqg9560mxXhclnxjHNEnlyLUjP+fiOw8dFGs206h7raKuRoF/W83F6t4Zq
9bOe/my6fTrOZM8dgncVNSbAqRIIOjvwSI7oXvEeOKv+ZcMyD+PN9XWlsCnc1pS3
VTixU9jIlmEXWt580p8Ar2MVawNewY3MiBESlyHiTN/sKmhexga/s6iybbTGOuYT
6qPtrUxzeQV9OMjZJVEX4h4B+0x0dcvZMavFhQ+noqeHXGdp0bWJpub9ldMFsxoD
GAepSU/1swIA171K2NSZJ/rOAEnh8HxoJ2dCezfNTBOY/rmXO4lbbV6vGoz2oqE6
djqkBCSx6UOMLMIB3Uf9pfXHLKXG3DX1vV3DTfCcokhotMDuFarcRO4mQdkwqw4g
SUC/Yh86dal+9KeRZgmYMmcToVJ2kJiXM1IYc23tdFplQIOTRZF2C79Qe95RR1F8
M21x+5YpDeDU8nMBeuKXPT0A0dEuHKgTR+htHbb+6jm0KhKqvfk4yIbwNfwqbFqb
tCSkD0jffxGTQwIBl0t1FzJClSCD5pxsUA4W46yJpdOPtp/BaGGddtu345dceNji
Qavo9AJ30KjIy2P63BzM97OYZnFF9jjoeGw0SntKNXMFPppNu3csgrWrBv6MRosc
1CbShBycm/BriYsJuqyhSuH2CGMHSxZKRiAvgBeJ1+5+MKB4fj7r9IjMrjU06UQn
MY851ta5jvaLiA2n5BgC2dn6Ri1tcX2t/SdzJL8dmQ5IR2Ztz209baa5cns4nWsn
Iad+d0pmE0gSZ+61nIXL/pHsl2osGVBEs19g0NSfhVp+xLV0KkSO+7p28PEIovl8
XTDUfOjVoxYyL9N+/keQ6y+dTAJrPRRrBS95fyvzOWPW5pUdoRtSxopyVvUHpSXD
txDvZGAK7oNOwWx0EhJ6pe7mP/H8yLG0xrLV0G97GrgV+/QGTUV4CzWawkdITMnF
kXlFvTczbjj5qwu2AzTR1Vds7oULiDVIHJEg25pNy/7isr97GcneephznuZ+QUSn
GfGx8wWWiZFwrHuFYOy2WNGai+mUftkapHR22p9n/sc11GFjagK3WI4N5NIW4K/t
PvlJPQ6D3Cmeo9vNGXXWDqZUfoRIE39YxSV2NEa2G1k8bZQhq4Hxj0nz4Wm+jhTY
fIKJtZCrRcL3otK+aHECoQLfrDCGqnTw4NswUagvr9s0Pys+XZOsJISuMNNoA9OQ
slMqTZS9K4QaoeyVBK9VxJdePg/94glCTS94SQyb4EarILEJ3h+9ktyu4sadKjfi
N9dCIkOORj1QzunEOoiTqsGzY+3whMWabLjiXZCZAmEf7v3W5oYBo2nWhZfkMB4M
SZVCjXY6I9prFkcPLzUHIWT4sR5x3Zmvj9axSGSVugvEFwmsurk8aevmTrkp28MG
BMur5XhutCO2rES7tId/5eBQ8/jhjNfkL8afgbHedaaIC7coSz9X5D+7Vg0SMBjU
NVRVywchtjZFKk1b4z+td9THFVFqRm+UBjG08sHbacsm8f93ih1r//f973O7RHWm
KjdEjWD2NsHXU3qeXU883ZDQI9gxeditUNZkYnUWu80eEYm2ZIm8JbzG5k+P9RtS
RPcOgAcGRxTKm7WNhxabLFFLeRbCvKyiqX89kHgFIfethdaXhyeiSPwZihf64RmR
xXTUzEFmD0KyxHdMwmDHqwGJM/hbnkyCGIup4ya/ug4DUTX5jzsqtoW4ptbDH3rv
5YcTsNOep6CyTiItwpTT6jh/WCpEEFQ94FAJaaklPoBvJwLqCOtLIRkWkZJEhI9p
02TK8x41JS0HcYOUjnkZGrcC3PGWCHQZJvRwEF7cPg3MB+DzqD5J9eTNFVXmbyRR
NLr9FmJkihan6ooqZtdiVT7dLQim+h/SdZShSPs0egOuMWbp2nVQ8E13z4MVNxv8
P/gWHiJwmcCMjl7EVwjKKhp0wWckccr8/I4Yp+Po+J23U7D2ujy+xr0GJtX4Lo3p
pzbosdRN9tHX8AH+RGFt+zaypyCApt0+tadem5tlJh4ON4DTnRfSQ72t06cTlGTU
VOV52v84sRwrlH4kgdIfKfsoJ1DCLDTEYbym7MZHSPi2pu0Dt5ptxeiV8Ijoayfc
HAHypuVKOyYKXjDvh2M8RzIbcnRefhO1ai69rbSFk7/R24KPZOK3El/nFRkw0MVC
66WTRu2rJWvA7O6yCzFOCxYT6IAS1xt1t+RWeirAUF5F6XTfeGSQs/PrrrN2zAFy
hAAx2zaAK8nK/+JWXOze5q/ZBgweVigMjX4alGA6swOTwRiW39JsXTVLcTqSu9Lv
NpS1fSHn+HpCin5Q3nu/SvKamngONQJdQDM6emfGBYzcxtJ5Edma/KuX49XcE3a6
CvAmRuQRC++uocgaj7yBWU3vDWVmid3OhkI8MCJu8VuWzT6eB6i150RB+dB4zbse
mMuNxQT5qFb5QvKSvWzDqcbs8LL2bVivEmywEGCkMSZb33cT3yoWt+i4he34DhUK
KEh4F0NXAJ6DJKbX9xeHuuPjhoJAZlndJNwqVVEqKkLdnOxT74CFtFB+A4QjzoJz
e+UJ5UkjKQ3shlWLz3Assmbv365tL54haQtwTOKASXkzNt4Dby305zRpZtcr+k1k
DPtnxLlF7YyjKg4hosMyagmBQXpc2hPOno8CDcBz/YTFeeLCQnOFqOVBP8XJm3kS
ICfLuvt3NfNHLQh1ybOUJcfTcwjzmAUUJR2MPyJTL3tD848BRHUgh6S2pvhzkKWY
8OoK3kMd2sPPNDv1mk8FMZLuPsNsuWdUIZ3/CSItrxl5xGbJy1pKllzXZbtWJIH6
sNY7+NdlXSivSgxK5y016bgmTtsiUSTZHwLcHi3FY+78vG03vSgMRGQ67ElmF360
Dpcfh7/6gcsXhdgSb8OYr4J2OMxOfAlDQIB5gWjemyF3DomJz6UpWSDqSDc/hFK/
u1uXp3z+xh1uhNgSnR65lKtMwVYy6prfki3o5c7R/3WguC7IilFOvgTW0OXR6Yhj
3HBvP05ehsuMwrJ0/PPO8GdC2+mzaVcb1gJ5v91aJakJLfEvjjg8mQ6w69NOoxhs
apfylF2sPJnYADPS/s7kmJDq4CQpLPvCKOjMjtP/eIEigBkjsKuet2CMj1zcNuYP
PO4Vn69DpPNNLvuurI9xRSxKZH+b8gwliycjMlq1H8gXWHfeK0eBqWdq7Vckm4ba
sLvT1GHQ4FM69qsCr0DAE+df7Q+MVQekftCojq0XKjy4sEWfMQP2bOXDEobflUlp
H1zvF4ZQnPR0f1kNeaKa9QrXjdodYGiescTJshd4nxwXdkjZrc9wuYqoXO56iwSZ
Qju0FYEbE2DOmbKhl1SE8yfzOOCZFaOezqPYbDo+NyoSbwD+i4XqBGk0kxQDIPhU
dpKbnD4EQY7XCMovokFG8ONp9V8UXBHKkXNgNb13ShrkCIb/E5hKINooWTqPpoWC
2NEU5zUbxQfVbkEJvUMBqTRn/9yOaWOmDhftyOhYFwB/fONDNQA3mq6DJ5k7vAMi
qc197x0f36ORs45Sv4tRCVbTV+3dTgA9KKshQqzwRzJdta/02zFjXmsCP5RrNS3D
ZkR3BDGiz89gs0QWPDLa0m+jR0mFFRjYsMsDxmzMUKbCYlqEk5wiIweiVPi9hlCM
R+QrTclp/BOKkw8oArsCwNZOaPIcDZyD1FCvwJzOjvGi7XinPPUjftwDviKcJXW0
Ki3TGL5xf6szb5hxVrsKkebrsCWHZQSAOKmgSN6t9Zm5iuHgaJnn9kidAi+mxG9q
ZRVzfiYrfK5jDsDVZhlATLBu2q5iA1aN+tRFavh4CLwWuspSdpkLDmaHDLZS7oOj
NCMhMpg0WWpOB9/1ZZySKVH4D5Z/1CHZglcB8SBiv5oRRzkhoySrFV4HBK3kVTfr
izIY/JHBu/XT34YFPXdIoL7iqpuawLkbzSQX9hQr0t3Mi3z48xUZQ9Qd6atxMCfj
tJY/Rn6s5StK7Tc0WzfiZahj2go82yv9Fzld32+TLFhsOiwXCU0nquHrJ/MCuId4
sDFMLqFgOgyqdGyzYy7PGbF2tJIaCD064Rm5jQyrRGvXMPGJZWk5P/WDOhHb71tB
1dGodBhxwfGrVly4G0OoD0NYSdvG4Ra2b0NFpufIhSJ24EGkzg6jMI7CVbBL39EJ
XWp3ngaY9K3C9qkC8FN/jpSGjcLka2rXSM8NCHQWYIPg/t5Zqj4ug7qEUULM247P
jG/zMebV9nruEKU0aUB3ol1Ozvh3VyzxEpjrx9mr2NzvZvwxzmRS/hn6pC0rwpTb
tw5FAHbQ7QQndyHk4PmSIFcMuB5yovcqJhEj7xWgyp6VOBFH4gB8hBh1dUDjVPpA
H1A1+ZLmvhzg/mSsU7sEmkQ9wwoAa6Drf9kAvOeL66Urtn69ASMfM6K1whGnpOXp
D7FU/gwjtI0WRIuHb9PpKbBSBh1zNFHc1E6jgpkmbM8NOo7RLElW8MYVYYz48wz/
6YG2kjq1R7xXvGdCv1duvxLAEu7hSDf3xje9TH/oGluUeqgaZG8Wbz5/0HnfcEsA
jHDSUzuBRPze4bRXmam2UWHB8TJ8e5N+G9sRCtV3m50mS4dEaZOZypcdMuSGKrJ6
xd/JzWL7y038EQe5l9JTrCMH2UBqGM/+XtEtJzulXQAKWYS1hiFop6yQmRgY3jip
iNqv9Gho2aX3Ki5b0tZan5dInJW5VrMwnr6HFjLdGUg/qRSyhSQz1r/Cr+TJRzmc
qhN1jNQCRe/TsveVqS2sK1jgjnB6AaWHLzkEUDaeMQw1ZMqx2qbSYVQsrk9iyCxe
HOOKR5nQxoIvVpNBfOF815NvBoFiO+QdUn4hN2eLXThD6PdkIBuN3fppSF+i3aXO
z+ghjM80d0maU3Whcqlq0RD7Kk4DelZWYDqgo5VDezwdRM50hU0VicfgbgqaPqYA
AQlTOCGs5K3KoNv1YpDL7VuqY00rpDY03Aab/2EzGjNld315nFLvbkf6rwUlPJpr
h0b8XebDBSuUeQ1RWcEiGO8OQJaMakKm/iVXLdRrlZXGW91TZhMgJK+xLFQ7aOHV
vLQu/ZRv5SBKIjadzH9nEZkL+o6NclkDREoyE84gSHECtc+XHJykBV6NxusI4YHj
2LUnfJKBEcZECp6blZ9G4S/SsEq58+hycrxOKiAPPQxbJoQDIHWvS+Zw3LU4UZgb
NuqCQB1qwUI253RXASUXCrVm9fwsuXpvRHOMZBrtFaW/J/Sz7r8eES4v3k9ZaOIi
zx9SmgDvANmbP/Az7ItFaw6zsqbhsvSebiAY0J7uS/7QkwwbIv5fnzi3ojzG+iml
F0/HLs2lRV9LcAsr/swB3DM6iYQhZ64pNY/x2a+QTneO9R8DgCSqgay9ATJRDJIS
g4vvMfO3BScmSc622xvz7RmDhnB+uasCQO2tVyQc31IxXRgemDzQ5JSLoNNx2n/d
8fIDCOaZnS1CGnqA2ZkVgg1HN06l9r1VzIFYKKi+9AincgsqwueOH0fxGdNlRuKU
xx52LSCfAUn9CGVb/Mgvwcr/zFnvpju75xZG7hKSb87w7r5Fs1DdzQCD/Hm1Nife
GLq95Jdr7zgZgY2tF/lbSe3F376UAilsrrFaBnTtNuGjwKiDzwA9cQl9b9oSsOhb
zPR7tnTs6Bxm02z0rleb4fMvPO+i+U5d58b3mMbcLFc0FuptoqeAHYf0bOoh92uO
7bVEyVerfgJw4KXWUvkWxAz31gao1iG1o/bflnu8bIHtmB97/6RlnnCKxgXNuG2j
yS5Q+y0NyXQ3dic8KNMWoOG6TGlDwICYYNSOznIVN07AT8gRiK8ho+TUl57SL76f
2KDye+tkZIQ02TcMY0QPr7L5M6TXx7lseduXfayriPv+deFmP8jcfyAj5DBaN60+
X3hl3GyZ/4ea9pBhp1XuqwsV3zu63IwW3vWHBzBjTazm9CgA1zpFJlXJCEhd0us9
h0YplMjFApKjENMYJtN/ESsO8GeC93LVwTCmdHNlCd2NizjEpJVEd1urxfHYNAV6
eMhfGT5CbJ+uu3cLDGa9mjYnwFyvtFJSa85x2dx2D+75PqjHOoneas8InXG4mpED
S7BnLFwxFQcZOxKY8vl53iCKUCCdsKQOIUJ5dp/SRIe+nebH0BmTNHolER1j3Ber
hpsm+71t2VvVvKDGVQgur3SxRS9F3vniQEt4l5IJgICi46aoCetTMTDlO9fdr8Wf
FMeKFvfbXHvE1GYIQ2Tq+U6o1399JI+PZ8cy5Iz0Yn5IuRDAGkTcfA9YQerFM6ld
RfjZ7xPWZVQ1akavzAxoXlr6Vi1eerLa/HEk7sCOIt9UhF6hg4P0Bqo0goAlFCSx
VEfYi5pDqMDZgSlci/OsKOCo3NK+g0/VKzE5klJPL4aRGcD2tW5gSXWd/z4lTUNg
f5OYVBo6aIN+n0pXc/1rkPnuLJ3/oOahDgTLMjZDXFujMvfjiygDcNKAtG9N+ObB
KT5T2NLoJembQctMi4DW95AAA5s5QQpxlaMQ0V99gyH5M/mVRRCn5OiUtKU13N8g
gpw+GqVL7At3bdWEuM6gErUaPlwiNX7G0X5VJJCcowX9oG86m2c39xFPgC06x8Fo
x4/IMwCICMuMtlxGeueI1nqiEaVd3mysMuoioWGU47aGSEm5NaT8mYnD0j2hLlb5
oGQUr1l8sFW+iBnMTVf4iT9q7VXUqwOxW5/ODe/DR98UrRjoNzELYUZ0K0hEMotD
1pb1oxFPMSgY9hEsbPnQMsLVcMmgfVEydmQRHTZiv4tCDmrv5b9owFd4yz5rjdqw
3j6J6ZgOKGmQ4TItJxOREsN71G6N/VTHUkq1pQm36QZ7s+CMe04qs5WtbkKYMFTa
KvQiPXRdxf1UgIGXx6bFLTaYu0r8gDEsx8vojvpWGbxLntGlzIWM96Bp8kIV0/jh
Iw5FiGL6uSvM6f3vPXN7bO4WaI58sPG7y/xYkpURjyOcBUYZeI1IT2M5FA2yQn0y
n/wxIm1whUDUSwI0sYpP2RkbqPjTCA4z21+Dn6T5q9jtNY3MUwXO7Ou1V4D4B+K1
0rMXxHfx/rhM+xjZd3sikYCoHHhQ7vMYf0EnMRjlHvkJmq8kPya1JXvuVw24bJ3d
MX/MpF7waT1TXweW7JBfbRyX/tCFF6Up7yEZZK+jvxHyIL5JLayvH0qVZgzYYZtm
aB3jh6D9bQlgZJ1XZjjTV4GBnPaZLKhp32/gZLk917spHW7ZvZqRQqtcB5wVIbDV
qjWl4l0px6ekSSlotvOPdWpIzjg12lZKCbN5a2swFWWUILJukobOmDTTKOAdjMtm
yIma3iuMPqew5DXJ1hGbEHmTByaY5Ol5k4P96AdsEQgRet2QGNvR3WcOVodT+VsX
0K1lUoNtbI7ajsApVnKqcwIV8nG/WC9DcslZKknFrCLzRCNhZ5ePzuAbwjGhhw7+
i9xq8l2AuCc2HY2YI0MaOBbFn1lSR7gYbVuqPQVvEOdqlvcyAzVyemj36DDpPCFt
zkckJohE5ZlbIePgXZNuR6VFgfF+eaF8FH6jqLlMEQHBGOwW+chfZQYegeYohoNB
S7/qvEXXCC4QbjyZp8RSTPHDHeu1e/1tAB61QggIiPpvlHQpCPRlS4wuUaDy3cs6
rEUDJS/Mcokq/T9PuLSmjBzdmPyhFetF3Gf/fNYoDAg9R0tm73Lm337XwXKlMN02
qElPrN5U/+a9xZiinTah4/KOHZ9lVnQ62bnwi8VgIgIqvMEl3NWkYEUJ6bAVkRuT
STFKi8ZSEG4DsehsFRvzkfM/8v1gmaETz52jHXICAlNio+S+j1ywC9Ap8LCfDBAq
4bHkCo475leFNQ5iUAw3usaEqLTVToTiPMIvPf8fb14Nlq9EOf1MRFWSlpFMlDq7
TYy8eRDF4nVKAT9QjDMZbk9HZ41bKizRvrRZ7sQFOGySEkE9NfuLnYPpVW11Hgvt
A1cFVAc8stBtn9xwFQL96IOPTasIktDIPt6zZt7NjrEG9fmBofkcA3EWrUbbrXsW
/WZEWtd2/5Yw5AGAt3zCepj7R4BtILd2MPnP0JIaYzTUjlPKCT8iO6ESNOTatKE/
AnodLL4vV8Cb+gnkpEipz8iFZNL80QFN5z0UEiUygCJBrOwAWQg9FkyveEVBid4U
U/JLYidXpz1h8U4aca3Kp5BSDJsV6diP3/jdJLzr2WHhS39UZa1gtkKREqpn90nk
JRA3diUvOzf+x1vBHoqoF6psnGEAYq+jmWqPAFZ7RbjThYvVCgNiumaD19DeVgO2
nOae40ot6ALADPfHTb8YlVpUEN3hy2fzECY35chl4BWORFt57BrHsOimWGVTbBya
JTdW1Wg4eSngyyBbUK6PC1+V7wCzmXlzDroicuibPZMqHRNQLL+gVmgxS/hFPsMX
deC3jxvqohWTAavenDxwRR4aOHYP+AMU+2HKHNlV7YKgeY/xg3Do7diY6BGL9iVU
59CpKF77vQfHjZ54PMPV+/mRqVp59VU9gLI/TMmMh/gm6TuSnn6wPJC2khPciKRJ
Rg2vzn3f9nBz1atuvHUK9kveQaxVh94PaGKhvqm26DAnlFgGRglD9XFl+mJ55Oy/
1L3HS7nNTtP7u01W1Q5rdaWR7/t7IOGqXusQibY7mBL7LX3egRpjEfslaVPBLYxW
HbyR48nK+Okkv2FBieIrILZERNdgVBQcKOQ72bTpZQTSYf/l2dPwVnP7NocU3i13
ADM12KxOw6ZTX7tw7nggaBvmaXTtB13Rza71Ayadj0nvsb/Et1MoyeAmlVpqLjHm
FJZyYIAf0VgI7jq2WLhGxkRG2CfZ8zuIkg6r6ijVrYWY0053jmugQiu84vf27LE9
2L9rE+mWTo3G4xYVaolp99G71j/RFiTl59HD5BKP+HqQzamrG3MiesszAl/2GMnT
oS9oXq5OIID1CrndocSBFT43jO8/28S8KS8y9YptRiVl2xWWGv5+OZXwVsurTbbV
LGouUODD50PS7+3ivX/qg4pv8QPLW+ytKTz4vkV+bd+cYPvz0pliNeh/sl1ZrCHm
EmSgpeGtVWapBAVbXGu604LgtuCj7ghBmOp672QbfDMPqAHN9WxXAe1VMbWr9I2F
AsdnR6KbD3hfmyPzcOAKfuMzf+uzstwoGiENLIUsD5z3jYi2N8VjGkL+ItV52k9D
0wwuAMCQh6lPiNRakMQUp0pDSQK7Q+vHf5UKFMYZb+tbJHEceog1IZk70aIFd2Z1
VbPCZsy1hMJqjuvqaYhYz7rPvnxmwLipnxJPsRw0bGZUnEvfzRaIyTvs1wrytICX
UpYQ7V9nhp5zXRRjB0Lft6TyZuOjhsLVLc74q/s17szNl+ICbAM1pGb/QAW0oPSz
2fZF5fhIi5DcmuS2wXhhTloyVNkH4/tplNATcK+o/z6uyJNu7uvSCvjDnlzjZGXM
1UKslLeyyJGb5cSYH/4tBYt5kjHZBx53mb3vhGZw1koTVHKhq9i5eLkMBkrs3nh8
BF3mZ4dGDWzmCwxmWmLzAYuZM1ykxMQGjbanxPHDiyqTyxS4s16yZgAyCBMRsu/r
guoef+87qDAfTmCFmFSgasNkIGPV88dqOLhoGf4cXXuW6R7RffUSh0OlkuYPTl0a
MlKJFxMlqCH+Np630lE8sgw+2NaNc9vkawTU+B+6/kz9DzNveb1h0kRRe2Suu5nQ
C6xOH7V1W/uxJL3LfSdSv96cpmUVsOs0zzJub4JfqrGQD1FYcrlW3EJuLC0VAjVo
HKplF3Kbk9lwCkoR5ev8T14Oar3EtV62tTaFaOLNBjXLOLggiumod78pT38C5p4t
TX80+B1IPgU7KcnLvf9VK1sYPIOvmNzmh/NGnPQDJJUCnBY6aOqbyZhXeFl8Tqtb
8eZzU7IrheIHGkPxN2Z8Zsl59kbJQHkjfaRmdD78YAEj2io/LT7JdOGoKWZIcDzP
nzZr+cqceoGd5N7RV8KXRI2x65DvQzaRSrLCQxHYZN8Jt3GvFi33GMdwUXOvoklR
lG2uRQPyxhUYTeX28K4BAxsUKtmoL6Gyozc8IfA50AwgOpTanIxqryAu5H/8Tnzw
3SxmeZIlC9wKbVX7t6MgFbNoRgOAu9Ls4ZRYZpYFsPRLG9hp7a1gUsiDCn8tWxVd
YuqRIokU1nJub/1X1hlydDyqbxtvMJCd/DgToDU4MV1+5H3YIYSXA/D5G9zrArjF
FvbLrrbUg14bOOVMLtR+heJNtgPvsP50fZjPe2H9hcOKjgi6pmItOWY5b8PaecVW
qrQGV5hS5xBkmumZ37551kzmWAtqHUZO75SiF4ZiRSUcqYm88t7HE45WrUK6hSMD
D6gy8b/KGE54k680eZF6y00qoVlmQNTQ/lvMYcd4xkZz0svgMDpSODev4hBDCpsz
6L270mejRxltibEBVgtTzqmFd19I64LL1Jm+9hi/99qT684lOes6VbTxaeEcKxBS
+mhwIllhjxUDQDFLuRZ/09PsnMIWCVR+Vf2E1SCUS03ojwTHjRzPMYtEJTrFjCmv
n+S0ifwTRM3ic88c7o5u3wDl+xZw2jfLx584n5tP7Ru6MTCvsIhaJDPum521LUFi
XqJ07UZsAP+tr4ZqQ8KmiwhoJhps0IQQtcgoWfaUrfOcwyWHBd3XH6kAkfxVA4nA
yP1QbGHn1zkc/WhdmimXEosPXr/7ayPijYHPwyhR3eat9eWmbfRYpg88n5XY2M9v
R99fGhHnNdQTWB95HHHR+vlh4EoqR/TrNDbz5gbo48502BYXmIuuIjys1GOfwmH1
Pi/RYjZtH706hecyYxaLG//8TVlWftcoqVweijMTCZ/WwwRYfo9ADAENgcfpUusF
8ZQNm5F1ewNXgq/gik7O39Dnu+9XZB9ndf1jg65iRA11Y776es12yA0VM5Uluim7
LTaS68224F+QXy/lEv6NkEbet7WYjnW0D0fv4aj0YEBoLLCKdAdLlDDY5uYMOZCr
IPAmXikJWfaHT6gQuUREJOycxtejAyHuUoKPQZW5Ixwl6HbfmUYDLzCVC9R8kazW
GkFcIX1WwU7lGgBKrGhXWBWg+4m6EcVPuwV4rdedRoUnk6nLnO1H8j7EsU9X7POt
GaJWcGsb6C0+cbWHa4lVqcIYGWVeOIumCKifx0cwWLLqSBy5tE+qU5mhOFM7zspo
OMN4K1w3vTmDjSoohpqi9gBoVcls5CFhzklcgwIW6vSX3KgaUcbkg1PuEkUBZkrt
By5odyhFMcC1Wv2TjAmQnG5BxHXT8cDhpq1SbWZ9zEyIlBXDSfidwhH8M42Ju/5z
Zb+jgE6lqojZdNMvoLPHNWxOUI6NpFi2fM/cEPfpUlqvZY7RXUCF/EkH5VLp2Il/
jE1cPDkx/yLDNkJcNjn293OnM4zUch6klPoUG86NpomiszrksxmPifMYb3Jj2yLN
k9mjCGnvS0RV+H5+KizN3nHA/Vvn/Y5AzuXpG2CHe4usKOGopyaY9AcaVFkXoAal
nB537e4JbvXKVXr0JXWaNEwhMg6jvveO/qBH4U2+yPFUcm88ueCrKqLcZz7vYV/p
LUnFtZuCMCHnAubmyLhYTNlnOZqFMAuxnKUuRg6RqtBUs4eVngky+ibV4xyKqv+Z
lBAOPjHMb1wH5ykwPlw2EsktQ+u+hGuFVoeXn6T7kyJCgblmlT1FkXNIvPv5BKP/
o26YEeG+0PFx2DbkFaYR6TAZH0m/BX4Rju+UD2TXpKVu69v34NxCjE4dhmLGETT8
nYphkY5JtosekFqvyAPZmkh5nUV/h9/s+EhPLg9iPRo+dTpCipRMa5R877x1j+FM
ugSGCdwwHvEGK3Ok4oucEveRWTVmEgf7cEcgFfrnkJ6V8VnSns0i75O1t3B5HXHa
coOpj40QONS+ohGx9iJftBjbDP28G/XIFu7U4dF7I6Czqw0zi6zG2W9+fy/FoZV8
KRuXERIxVq8VRGrABc+tY/6fJlePIERuh7iSKYMsBBraHwpPoljklyDOctL7mHMF
Ev9M5WZd7RVuK/bgWZ66dMZqqEU9lRDzNYdaKhFWB7B3WQNnGCT9gnNYcTq86x77
yycNKaIhxMhPBhI55Gt6a9ra2CuitEaw+UwPDZnxtoKBbU0AFNNJMiD9nCP1rBk2
OKY9vRGg/kLDQw0x2cUgW73XeCxEvi2lwSmSoWHmbOf9FYr2mJ2Ey0xbb87+F03l
ELZQuFUegWiCBRZa4EPK8teOW4kiTK6hVmgsayeyabBzdjULRd8E/aZGdX5aP4FM
I59/xFt8CaTCbnLdvTZ2UapX3WKzlPZSDWFQimWh1b/1w01ZzWMOtA+lJT1IUA5p
Hw3SLVHN65gTMj6jUU1kILPmTDSje6HIMy5t3O/yZ9miMvwcnEc6O55K0pvCOvlb
t2BvIAhBJ71+/k5FjoeuZdRGtLkrfCNe3A2CNSe2r+g5xjiNUr9e80M6jJLNoa7+
EjmmrKcoOKG4QY6dmCD8p2Xr/YPt8E/9L2otLWe/8PW2w4Dt6nOQBIFswEKR9x5M
3/VZlgOGN9WGAmlubST2o6AmNtmZJ7hRBdNAdxDZVGxrP8pinvk/f/pg1Stm49QP
n6e0cCMyjDqRPC1anslITdw2gOM1186sJBzKI4oPoZl5KNkuuMPejTmCstBuNRdt
cpcZHR2GzSAf+f/rmXcgE4DgaVZIMJhE+LdW43jL3QbJFp0lgEZQBR3TYxYgPusW
V2uogq4M8/vfOFUdTpMoIQfwtoUy62f8Zts0Ve03UnnWZhNWg/8EiOddGUlAICy9
dqJdAL+lui1tdcmJT77hi3PtGLZ3WNYRXdWcg1R2X1aKD5PJnn842pVowEHuiLGj
x2fNAyh5G61tcS0Lk13Eq0kCo4lW2IqWww2bzpMRTx1BdHl+9H+BNnukuedDaCsQ
mqfC5xugo1eGYz9Y/AdGT4UYefzs6ze9tD9SJGL7zBG6DZzNtYrVX/jM3mTktyaT
QRgkQBTLcdj4ZB6/W07iveiskUQIqLcy0NwtapSPC8ffwPzIgrIqpOhOcEifh/Ml
gT1ppzE2J9nk/0EcJ1ajPr7M3kRdoerMGeu01PDqbme8AFtnPssSfrdwdMjYR/Ft
YF92rTz+8fMoYi+EjA3KMPahxdyBDn23f8r6ugTuJgPmMBumEfE/8CQkstStiJYE
63zCzfgASJJ5ZhYloXB14Lfx96YrT3MfaiSBS4l7SsKgOdJQM4F5WwrfxYZlh1fx
8OlwsDND2auAdeMpfATbRkcltXzlDwj7JfMkaXMWZyC7WvyyP81Zsbm1beEm7Vvt
7Ut8FNl+IQYiNv3Lm5ZI2LYDq8v241eZq03E+Grre4kOY3IvxGMamoT3JJhrMWVa
U9RgVyo7CDKIAfhhcGxsrnr7wmukVWFVZK+FbPBFbxhb92MtNq5fGNV5bOeVIl3d
ZjSf6h+pR/WDtcNo++gb4lbhdSVdHvUK45lyj0GpDSE+GhsPEG24mlPVtItoVKra
uUwZ4xKle2Mmvs4KaTqEOUW5TYGAEqBqcb5mYCAeCIPVw4f00JPP2u+wXB4OPTno
gq0oGqDR4p8EF658TCKNzf5w95Qk6hvqOqxN1er5LJnNxCGonrV4kZIawZabbR4G
/duEENC/xhoJfsBPxKjM+W7IWJ9YNu4n/Tpff2g/8UbVZ5jf5F7xIglI/hpGeVBb
45fpcoq1nm8IFDC7nNOj/lDvzLHcgS+5dvfS485kldlG72NVah+MfY1nSpmnQwON
ZqwvXbCVPrgFFu36AjIWuOEzuhV6gMNklw5YnA6HpmH/7bd5mzMyOGDVyTHRB0zB
0oG+xCW5wij9GMD2TORoEAC90NKSs6ZTbbLtByCUVf8OBsoRfQX0+Grdy6J2/Ltx
QIxfVrxMkMhkE/IOusuP334Yd3TtE8/mU33iamAwBP74rq8rg2N9SPkQWUV/EL4w
uWSuRvgWLm4o20Ucm2wqk+PrfbECOXjByzFQ8w/vJ7qWZKErjIECHYUDxUDx35c1
TiyvGiHS14atKejMhxqqCX3ppJNhWtHrAej8udSFCOcdNG1IpDjiIOL0fiLxVMuE
2smo9+AdzOHHeGiGTKofI/Y13xpANJArfof1j8WHq+gJRXapApvfSJvLgZX5OgtV
yPYvONh1ZoGLSStqKtWD9qMus7p4GGRTuOJQ9SN3gjsq3IG25DyATSgF4KfnlO84
/sBDnQ9Hj1iVhgXLB8Z6xXFs0oIiIc9pATgL8fOl6F6cXA4WKuXwtXpfDT3/Hd8w
3d9I2XZ74jHFDKnI9BRVLg/cszFWxmkpeQpgokFSTt9gc7QbuAE0bkR9pDDeiz9l
LwZNk205fPDK+QGLGqJfINVqDomd5dgteLQE8J90v2nm2KiB0NthZaN64BQ1Ugvr
dnnkrYVwzX3F1ED46YAT8AebqAWM7onOULpwiwTs7kUqcWPH5NHfaxIV59H1I48O
zeJlW6JdhmN1Mg4vGlq+54y1N2/SUjS5OxGhkolS/G7uzdhC+f65GjmkOz6pmQ0G
a6p3P4uKs/xJWkXqa2r/XRpiWga947G1Zg3AbLVOJSL7+o5dtbXGgLYkrE/fb0Ku
FFGTnADb0mvbn2/rm7qA4qDM4+KI22Y6bB2vY5BH3gmltpXRz9bUoAdpdB3kFt6f
Uv+Vu9Puf7c/GzbhAYcZAVOfmGMG7+pElqT8MfoeX0u+2dmeGhGo2fwRm6hsvGI8
PZbzXoCZodKZYWGwPv5kro5ULp+43r4CR5QyCFUSACICxzaOOI8MG+zxY2XJqQUL
doMig6+12HSspN6rpu1syHaBnGLHpRSs68Xy4o7+Lz2Iq3S1zti7TfwS+pZ6tVRy
iAeE90E8CqPYBMWTlvGw2VrRTgge3sYps0Jedpf+lqSFGe9sliqDoj7Ogj1nMzMK
q0sI5j39dM2e//CDzW2eHgX5H95biiwUabzmOUVT9brx7LHFJQaG8rIeu6eXeVas
Vtq02aVLN+O8ygKqPHjBro3HOMMsETVUqCgIdXWrfY1zsz8mIepiGLACoWgbie16
QCU1USlnupl0yYIqxHwGs8TIUuex2dDvuyoN9Iazb/qjSXmZdU9ij/aQUOhujlUx
T4kk5YrtR9NMLMMZWoOmAXdPgpdKbWDbPXoN10Ck2PD6cLPP+tAEvDvqpO5MYcGT
aMlB9c03DvcKGd9M0HEMcrjJjebE/wM6AW3jW35/X3m/D+MQX3b39NT13U8Ka3xP
EbygfbDMFidtPVvypjhg5lpQNg6zAlEdrlcVqw0zKNi7/UHuih2Sjm7SISCVYY1y
7VTszbDJ68fBtpT0BhUMmzrinkaQRphQm1GqjtEIRr7LKKfWTnhOUZ1G8LbwJKmQ
zjsrCb5Y/JIZLsEN3A8yEzq/IkpW2O+e/01rF+jPbMBlKlpcY0ouQfS+vtchOLTM
JMt0+wwFnhZADXQBr6umIcZXUekDg6I1CSwqaSdWO/oyh7aqSc1aqEGyu0kDflPS
DwgCdF6dieXAN9uOAbCwNc/j/Ob8IvtaQnDkkkI1C8oYgfmOIpTZDcVY7lhyP4jX
YFE4T2qtpPd4RZXM8gtJmJGJbHV0TdriOARmELYe4w8q5UwmACZO84c0D3PEkzTO
Jd0zOI6dF8+SCsIXTj/uKGblVaQX6jy0L2Wi7lNzxvWLVyOVKil6ejVfRterzJXx
zeD7x8/E8WziL7Vts0W+onHCuFWkoBHbIia+0iSvpdCVtYKdhTHy7/fOjmSqNK2f
lxP+LA3UoTJpjiVxZzEjUNMe5hr0Ax3wcDGPVRNQesAjAtWVERrE4xMnRMeCmPWl
7RLWicHvyU7HQEg42f4JcE7PGv0KSHkf9ePb+QYUNLMpxR7NQ3PGtpTemjIKUTzC
nClKY5f28TYJbI+fdOX6yER9t/9S4gBseSLxc6uppbBgX7m9OVKpLoW1rXSAGPgt
azh/l2KuDmeJ/+zaXZ82rhzAMuJNuDztCk91EXCHtthi2aq9qwYYaVTsf6wsxdBC
wSaGXE3Z3SgX4JPy7picmdAOxNkUQd3Q3k+s7DloSFP0UQvSOdvS6gKH3UVPEukW
o9iczQiWwx+KNxW6coa6tbL1kxWxe4GAokKirAWE0VWhFzx8pZGUGRZUtxOlG9Sh
y0ejPk5akGMPgrghMq6ylKUa90DkV5u+zpCgaLH+sedNYEFI0dyfJT34ey/aSOse
elCOrwTzHJLbu+QAevOTGqjbkRAD9DX13BP1SKoxbrEiv6N2w5BcJi+i/YpS1Eqw
Y23lLDqdIVhHI250mOmoBSSEqL6Bp2nfix0W3wwbiE0XEwgf51S0mQx1Gq3gZDXQ
uGJcjJN8HjaFmhPL3HFM0NqKCePI6QVaH3dKQ3PMAovhU3iOD9pMWBd7ymY1Q4y/
CfhXuV1zjKWTxELYbGCTwoFYi7H2JVslpigrDc2spZyYKMVuIqnAp35gl/XCMgId
8xEa2v19vW3xIrGSXJvwbmlvlIVzcHaWODQ/FSgckFX8+lbqlAHB+rwvrDTXGyF9
wKSAl6h4PFkW7dmAJA0M1zfrW0rARSvOC7pSGlSSZrfDPW2UTEROBHCF7dJyJHB8
8VX8vaAdU+jcoB5gYnD2r2668DblYXhFGzT8eb62+Hv++NozeRDFlXfYUxurItbh
VhRKqUFjJutngK0QvdsXLjQ7czfdlLKELV55uYoSAn/7lJeQojnymVQYte1qAWvD
NwY1pHcJyOOZ+rdjMYN8xpUJ9B0UbMrJFzSvJa1FR3TL8jQy0ckH+JD4e0U7Y0av
ibnaj7rkIrMGBWoeCNvW6oKCZAyw8gKgQZFJwTck8DgPrXpukXYJavGEr62X7sa2
8a4AxFOMUyf+dLzajmSxb82uFbD7OACZUQPZ9hLx50RmPso9u0US/z5lw2nN9BHs
BISqGYEH/szachxqGxANNtqvwBVTdH+p9+6qL7A+F9btz1hP1xRl/nDgXNyzAnVK
aW9mbc1JGw6W4CyB8Qho/gAXR6IHGJ3+53cmJhslVqyKhZJP1EBw0yYi2mrQUGwn
L0A2dSs6/UQyo9GK2AsUDD/iJD3qgm+lvEZQGI0UwKnELv6GusMNbEDDlXUWUXSC
F1j+iJ81aaCT0thynVHGaRmtvBvrukVV3xrKIrKRYeG2gR7crAkGwTI4Fim3v6zX
mADvMMIuKLXQWH9HmIyV5HZJno/f4Mi43vWgdsDLYe9g4nvom6FKxJq1DtNZ/lml
ZKvi4JS5v0FDMEyMI2DJwErk4RVy3Ber5lNAVdB/3FN4AMxo2T0VIxD1odBTCORS
BZ4V4dnT6aXJr8OVsAlVwE3g42AJHB/t+eebbRAwxqyXhepS0DCH2XPZwGTBKjG6
H6HT1Zxpbb/I5QrUYcl5TClIb+UNoOWju10tz0SJ+3sq7sdnYbAx9++uLBAcTGDM
8nnRcm8cgBEACxjlzK5Wbhv8zQFlUs1DEG3P4Dnt0m/fMQkGfEA0dZhLcyCFkfkN
ilBF9ARLIjOuDZlc5MI7j4i7cuXl50cVA9bM08qEPojjbyIVoein8/Denk9GB8Qv
IsfO5kitc4g+32s1J4Jq70d8AbdqvAiSJ6GuqY6ku2FVMgKW/DfkYfuL/TjaHPLc
CIuoJoO9tpLT4wbBs7n/7vLERysT7SJI6aoaqC6nWStxcTVCAeESYPVSaHPzSiiN
xiZYm/TsoQEY+P614L/xwkB77WMuSI9lUcLcUFdYc8uscCpyCz3lPHl7OWDje6Wb
Co7ngmOLhYOcCczNzZ9VNUkCM3A2KKIzqvwCLEe4XzmV0l1PPJ25Zw/LNTaBhb9c
1lG9ivzPDUAOBPYsIGlAMxv7p0UMA3Ca4tS4EysR83BY829ruvO7V+pEKzIwFhb+
spN8sZo8hyDBLApzHJ9rxCsqZTyv7Fyp7egWAQzZNyvCwtujGsCksVWmpwmQG9/a
BVseYcxX7TEc1Hu8KBjgs4Pbs8RH9Hz5xc5+d+IgHO59e/3viboEIpmW/XO7pWXt
UKu1uD/8qAbTa3BepxjQndTp6DqVS4vWIjbVT63tzc6ahNF/q4R8Mr6p2nRHkCDr
DTb7spYFipiTx2vvATmAB9PQzf+qrBdlT+6PxBUjL/USYnYu5qcjcPEypC3ZhhDI
RFo8RKfUzLSUWjnNfWdL595tflu1uff3fz9Ua2X9GrwjkE3SRbvQczUqZAb+fM3F
S62G7cBABFNzEmSy99FexJr4lr7psLae/PVmoqvvahs/kXzXrPpx7ghy71uOGEoR
zrSjjnH07JrERd/D6nPpiJ0gwPQu+LA4Ko8wtVY/vWBrZk8e1gxr2rrI0PNwpaNr
b9zQ7LVVLGkFZIOjm9q5e/rtTbRbbSlXjaWALVz7hnwz6w7vsXeSOCzYkSfth89C
810tBLe2GSQB5lpgvMIVGYxHxX9sSLoFOIxDSLzh1vwhzksKULldgM10dCNVxGUZ
t4rBCEO+OlnALDkXh/qeclJzF8GhwfB7tGL5vnePB3H8IensjmhhfzYXKy3D8pnW
BolWtIi346MO4NldfaGIGkNR1hLveowMb+rgqJ36Tqvpk03Z7canlsNnoJiXzTtT
0cMSZYP5ysXlLM6FnxI534FPoFXeOtFcQpXk+UVzC4X9L/YUofw9HsOJLqs1gkzx
P7SZ1nl2N9jHfaGGn7c9VSu3Wuy4yVo7xpJYj2peoqfed3ISd2r0LojU2wxlmyGK
nSkGfJmgyxe1B5N6+vkya865w4AKZEp4H3iT2BE1JhfDXi3V1ARK1pWtN0SC4G+j
6ho66OIRKWvIw4MrMNzkU+BGYgz9UCdd1lYd4QoaFKoHMYj63T8jRzJ08yX9eksE
I6z96/DLVGaZIHD2ceAcNZrBV7qr9FJonfxCZtXNsi6AYaABoM9YRT+npgx9YOTU
BV91h+N6/UuuUYDri/B8Fr6QXRgQ9nU9KuVB9+0ZxnkxGNAcpnEtXAU+dYtRzHub
s0j0v24+KRdKaUwXDvauDqI+nxhOwdi2eTZ0ZdulZc3qB3yFpu4ZG4LGXjK+YiP4
nrmlIt1FGLubwnEP1TGQ1Zau9XEiuXni3+yChOVLiiYGLNPTNolvNJVo8vC65ddI
PUHFITSIFk3BNdPhQ6AnV+twv8WcoKe0yMoFjJI4pC5IoENQ3hdk0OvPdovjidBR
1Q/mfoIZn1++rIg9g3Gp5ucp7vLhpoEVqMBa6E18yMqggTLTslnoB5397ioZ9W6F
k69qy4722IQumvvBy6wW1SRl7T+cnFFcO1eSA1S8xs5mz36hm26mJsXWKOe/fHvf
SW2nHk4P4FViLYUcz9NGGObSIAgdpvxjtmts3LIaLlXDknnznFn7WHOFGyCQH+0q
V4i3fyZQU/bLU2wR2kHQy0534Zz1TCcQbcvNz6FFYf8zB1tSHqJK3yFcyLI+SNTG
6jyq6Que3lEjm4H/Hr10I6cjGnSNW/yAKYA+PnF/i2Ll/sA61Z2Kr19XEDGr3U/F
sOAlSJNLNjcoxkJ8V2sahSczSOKvMIFzGo7EPZDRjfb5QdcXL3fUtE+8HXDO4Xba
uM2BR0KoNPFeyQ9QgzOhtL2u7TMNZkHzpB8NjHQJ5F23f7d/uvjBi13I42Kx4Hrc
cCmlT18jrj9AqFLanPJWFVRf9B3CkdbpiJ5CMZVaXEd1ShmgzLNHghx3/fccamNN
5wpDlTmOb1IhFDKCDvwqCdmpzHzLIcwiJHi60ARlm2U5SLGzQ08KGD6QZNI8Q2rH
LJdn69mISiN88/SysnKJbeSSKqm+X9CHb78BHsLg3RfqSWrFlWCcH9qyCWTQzvzn
LbYBhlyI3E3xvOmiBS1vtRaM83tJJBdebWWWd1g0M6CCL9hiJnct4OJaQomNSmR6
aCtLsEWqW+04WNyS7o39uUIL9Vm9uJ6GPboFcj63SUIqV+JzRZpkAzZI9SlqjUAH
3Y5AXxTxCH4XBw1adqbmhdalgKiqqa02+gMveomlBK9tm2bAl1HZ3nkOs6pYbSWR
lF5xcz8MAEhZf45t8PIO1dHbZ7GAIaRLoRWzSLLPqoLeKdXfm3soKOO7lGY2vCuS
M8tjjOCjyqknOsQbr0XgUTCq32jONFpf07JD79qMUIklJ6xWADUiR3RUfc7dx++h
VW6eZFnbu1GQTEcTxLWmQ9bSph+NeffCGiHZQzhdfFxoEjTqzYFZyRMKXw1cvBvX
EZ+P8wG5kouWkZIkJg6sCoHPdqul9WKb4cla1rXEVaU5heUIBx6Zv7Ov3PSjUUOJ
blpzIvIQAmGnPQSNINaaORTkQKav68Sn9WoByGDmtXs/sA/g6LMrgJCSGjKKx/NB
GLtJeufjuZiQJU0KM1zVI5iQXon5dlWBmnyUHfLBQcZhGXZf94qfviC5auOJ0+bH
zFkpszvfMb5NAiUcAMX9Yi6MD6UHvUKa3X6UbG8UETEhGk6JJeQ1c0CgYrx0N1AE
d/jACVazgnmnzwi/51lrH/6qY7SSe9UWtfJLK+gr8SjVA5Z0t4pKrmLoO4SYDmVJ
cuOdItSKwC/a9aVTbQoli2TMsGwnYvCmUxwbmhy+TkZMXL5shF5rT7CiRbF7rggc
ILLWDiDmHjKdzyER+Pk2VHduKeWIPfhzxzgUN0QbGXN78zpMdnFRpx6JRG6JzqMV
W5HR2y3yC289cwxMQIEEIPDgQqiV519KbC6BSGdBJWxLj5xm7erC9m7oLNiQHJIM
0dfcVlX5ZyORWOivh4DmXLfUBxMOFj+wQYOTdQYjzhjeiwKlrirVkQOgx9kZO9lI
UK2rS2WzXOg7qrAeWHXvshav29T3PflOVJhOUmSOkZ8QaXuosiPDfcq/9OJ3wBq8
QZvMcb5z5TQPGoYNZ6m4bZwP+m5BR4zlngQluJCoZ2cfLrkas0j4UIjjmEUTIbe9
48/E+VXKsrqdP50ZxyVHhBWZGax+l1B0ZhVbrXBed1/Dk87ZdMBm0BIxGX/Kj+5q
eS7ppTlMMxETbNbxL/EbCs+wmM0pXVSvHsVv7deYG1GVRRSFJ8QujUFGEv7C8dGQ
v8Gm7fUxnJcut5TluxDYZC8GcPNLlPyPUBmL7I+DSacNRJxabNVDuJ+addLViDLV
tpqBMriTjA+iQsGrrqWNSHZo3BuiJHJoannDJs4XnMrVDGbx6dfy2PJ4N9+cuAIv
IAPMcsPWZYquSthBm0tOcAyaa4NsoJ6QcgeoRHRsnixg8XY9JLsH/tbi6YxUILKz
jb8RihxyEQjpHDkHBPYlK3Pc4hFdrs85cRxlPHWM/HI15U3m7Yq2bAXAWbd5hXu1
YYHO8IyVUa3d7f7jjo8IIGt/lVsWb2Wf4GeLyc9WKV4P4iBSx5SYEjAdQIhDCi/z
tbXROXReaClowitRQ/zvZ9niMUx5NrxQldWpv5wubLp9lq9pzf7KDqfe7dHbQ+Tw
b1bg8KtydZXFNc9Sx4oPJuQxRMtBgq0lS2Vv0smX/BV+j0vw4aS9CD5Hk65YWe2T
b9/Q7fkR/FgTe9pdeZ47gwOWya72pfgZ2f4Axi2ifGCXBoWAtFJiV9mxMtejFKUL
wooqbCatu45EZaMCw1W5Wp5TkV9olSwWSRT+9Prtbn3ix9TFa6VNUW4CVMREK86N
YDAZaRNA+3mB+Tw20VGhYcqnMRPOBuGYhXlWeaYuZdD0vRmKqWlJzCgR20c2gkVO
XpEvI7PKSpejvo5eLEdz374alxZlltACF4c+tFZYqSFNRArEPSSST9nkkXGaeR5P
a4vt0Fmry7jmRa21dSDYc5ospXvqOZfGMhVSTaR1jSllHqal6+Mbi9u6R5dX9ib0
7hOOamiX7ssvGZRyXy6DjKs0zoTMweZZimaler1k6xOoEJEnQfcFwzeIn19F5WED
o8IzSUT5DggVCm4YUZIdurl1fdRW1L9uojvd34iATPnb2Vb0Unm/xUWemheb+phE
r9wJeEyy/8oIH6DQ2Kqwkj4V8myINkEYWLQk/uVTCautGWrtp2vlc7zV/LX9PvPe
nTiGEb/8t2J+mBTHKHb/SmPQG8ipp4V7j5DzemNwqgzq08SGInHkUGXLl/rUofyN
rTtmSuXBjIp5K93WxslDtNl5J+DPZ+S+1O0Cro6Ev7yWzkhibu/s9nfKSOuPDFjs
YCNOlK4O+Ln4iSNCk/l15/jOT6Gu+6TbzOcP8QSMHW+LeiYBYWgSi9zFL+GCdbeh
qGJ8OxLAHsPc/X4KxKLvPVUuR7VnULs6b8bETJU6XQ6+LFV2T+5j20dOfS4ekDiD
LfLzoWk95f7nxU4NdsdKJ8FjEn7cltDejhRFCIzvA3l8SV4Wm5Ugf8POjF+gmr8N
ZHUO4lLwajGLNpkZVIsQrb2oiE8IoDyVXX4VUagD3Q0eP++sWcjHhycSj2GOd80i
iVrEfYDBZ8T1CYh7oKrNUq8alzzCv+cHGidHdmdo+PhWl5J6N+5cmTIcCoa+UEbW
sX1Sf1VJTbBofwFXuTrVc6jE5SpMC8plMVE0mqFxvIxJPX5Y0RFaNzjpd4alPayc
6uAOm99ZiSG7OU/pnLizNNE/pH28xKHV/APAOkS0iUtmJX6oj2rIRNTuLSLdjZQP
xNkGhLF7IW7nJKXJ9724yucB/MLO4MFNqPWts66ZW4ZrQFprn9U7iwS0yJHCgQHk
kdC9XrUgr4g/BiwA9Ojv0xazvWS2cN6OsLjOalhX9z148PHxzFRWEm3mrIp2rvq2
hyJji8LN5pRbgKZy31GrgXxOCsK+/ro6oewZ1nvQqxuAVk6lBMs5RBFRhuYfRtll
gVceJqBBq08Prr0/8WbXFoD/crtRwMkmnvgdjP/RkMBWzSe6vs4JVhn4OxE3GwCj
xMTvurbR730AW5+bpDXeqLfgxfIt/BKZWw4tqCJI1N3cU2vQd0b5oTOo3mLvX6QV
LphMe8D11lfOEA3DpO14WWUm/9vkkB+7MgBNLI5OvojSfREPwdXXBUzeq6yyXr1K
VRsE8VQE8va0+4Ql7wB8FOHKKcCyrM43ZP3QX7OgNVp93QmWbz9kZWES32FACg52
pAJKZklD2WtUS1XP61xTVpD//f1aBi891TLP3sWI+p66iEcl5jEDFCL3J4DGwk+U
2fvc53eoCMiHux05ZD/2FJIZs8MivN+2hX4Qj5HesLom75tBocSLVDchNtygLV4X
HFmuxLsX7A1JarQczrjqzTQzk0f2h4otjvrIgAachF056eXdnea4akrBeoWlfhlY
H6OppZyHUI9aKsus9HjTIwbICRnXwNIx11PmL1ByLHMinuT227DKSRo6MEhS9MEV
7uhL1wE0gBi/tv5kDXQCGeAI6RaTUcWqWQsDNFeizKZUGWKJr76QakEbiQkfeuu2
/xMcc8BUyWJqd2ISsbM+9LQk24nTuNsdX1bNYDRi56d59721/2aiu/KQydRowfx6
bWVZ9srjVDQyCcOYHPCXgUgjXAXB4S7kqvttltjGxjH1n462iBDUkZysiJ90EehW
V+8ZnrAIa3u7zJYr8VjztrvkfwOlUropCgK4uN5yMZwooLbMAf9juhBSaimxfJ6A
1WSdY9wuUk/uFpDRyBl7oovPscS54jmj/gxCrYQfZMoLFSPk6q2bbzwwpi8wchpy
7/lWNJksq0y2EwmLrbXGN9pRzfLIEZtKZ0uduN277h8tjjGfKHa4z/wTVfLc6kyn
AmzrsvneoSSsx6LtXG1cJWKUwqkmJxCAmyTkoequ2ISf7zMo40r4XuwBmbQdOoPb
W5qAx7spGoZCzE0I0URU0NeHLZYVbYkqn3gpDjc9uyJ8r8AirMBAmoJijid7+ZgN
EdmvROxqSqRmxtT8kdIJDXLFLHCaewj+QeXRoCciX/vN5BGTmn+MmoC4rPfdj9Fs
2cHTF1A9KFN3gex5bmf6dYn331UV4ORKyYbFipu4uqI3IWVMWv8S8BOiV2cl9s8n
RIRlpStw3Qa7hrZYxjy2yDsvZ3IgcuvL1a6hqNJMkaTjNuAxacglOD3yOZlFhG5L
EQPasBzOY/2FxleXb8mFqj8AzG4QVgwFo6cR6cAfHsJiXEkD7nxcR1B79l3LJU39
elQ6TfmYAWV74ifDytAYRrsv6ENzGUgK0Fc4gnZ/VBA/7mW/55BI80HjRC0dGhvH
1LGzotgpUTVMzHKkz8Iuraaec35rCdVbhSxrhKl8n/KbipjBy7bhNnRwkjtl6qtj
sQNUPc6/7MX6GII9PEvf4J3ZJxg3jAJxt6KuvmOrmurntSMUsRLj5W3QRp2QZ4Da
eqGUHlJKTOXASSl6ZIutqWWKi0ZTuESqhc7tAPm/8OFFeD5Yx6keMTlOJuiEwK15
su0jix3s7+orFXVpUBWBTsF5iCNJGyvqp0Icf5ManNlMKURtTTDfcuRJyiIxLzZd
GtGshLzVCtYt++H5nqf8P5gwkMslvcyXZjc1lI3Q9v6akFi/vnB6ypSD9g3ALjLF
fI85xF7DvWGpgASy9WBjwdzAfULHVDu+6dwLDOaMRz7yzYklD6FWc9Ag2jgNX6s0
VzBgG3LUkTkPMh6cSsVzueTznYPD0PxBKnWFn+A68Db6pQD8FNSX0MakDh2gqSsS
bHEN6t0l38jn2FGbPpdaMNMKlec4K4t4o+3EkDqgS+fq/4PvulLDcDLxfhAfWzsN
cDy9AEoPAkTDQXW8kpP3zIP6BKO7mqlRB99/1mzJKDVedxqFaQrQ95rboeNB3Ob/
HIUf8R/OK38dQ7gEzGID0phw3SMTOZKJrBJ3hQKTlSsP+V2L4tG99niEuxpY9Mqq
iFDIsUU4TXY6sQGeMxqCBKfAaBygStRZf0xjuy0dHF/Ji+8/2b23ywB/bTPp1ASr
uzwtaGSE4X3bU2P/ffawxbelfrVodDDBMMUEqpD7gZR6rHgMLWooZP1Y42Wk9d3W
v/LjGlZgDDqKHWLwV7L1KIVZwcU4BWWjvQfpDoGPAr+m0Zs2hSOzh/u/ZC99Tbh0
BSxwLXYc+JKbWYuxtxJuYbiicN8JSdVfVYbqQ46E71NtSaZ7jwikh7MXqrpogjQu
55G8adUPIIrBjWG5LgtPzGKqCW9knHLeCP23fcvdh9wAI3KnFIuFADN083vh7aV+
BB/amyPM/RFp/KkZHh27vokea0jxraF63zybiv9+FadH2hkD7CAbCiUkR/IPzcXx
0SnhKsMQPE0V1opfxVWvO+9WEHM0+3Fyh3Gw2fGn/SBdoMvH4KCOjSz+kCxIwHDE
N162W1wB2qdYtx8M29P3NxqOe3X+UeoyrYdfcXSZ15kr8VnE6vYBEgekYzIxIESD
nokg6EetVFMtV4lrwKAEXeuzKURwO0Bs7FhsiDguV61Qqwd/fwd+5GZK53+TZSDT
E++c497IEuBKAiJbdywnjoTnBL3gWAGrTkRXN2zl7NxnhhTf9xBbND2bB3aqVqTR
0p75wIo95d1m/UWOHuvz6QxDJJpKCLDh0PDeH+rqlpBcFLqmilIoTiwiSPz2ktgB
QG1yexIaLsob8V1haxYsAKboi3nc2rA44UA5QnTjlk/A17mA44qpb5LkTrA20IOF
yk74QxfXi2Cd2Mbp1pmFglG+c6Fd0Yc0gFLx4FhekH+CbwmgxvCi/ZZM8PyEKMBA
PYgGYRKsiEIJ+1bXb7yTgjbKGaCDg0EH/XCoX859HPktBP1r4HEzYqKYjwMiYLtY
dXlZElR72t/aMw1F+L22IqIgRaW9SkDc2eDVuygfGt1pMR/Vqlqv3pVay2r1nwQq
3mvs6TvE5hf724Jz5kARjBDvKK0F7tlWzLLhZ+YodidzlzsC0LbQ3DnYzhw8toJ1
Ks6HiarHFvWmnP3qy90iNyuxE2HSo2mXI6k+nP0NO+qgAd2rVV9tr8CWTe0MyOtx
dKuNv2Pwrt0QvU3xh7kSoVEIx66wutXY5RXo7//UISPsiSMbI2CFm8r+Jcojh+9z
Ze8nyLp6mcSvq/yh0EDVSh797qs6+/I31DRsMAJBOhNxDidbGp7mD3jL6K9F0km+
yiNaTLNhZUWHJRXMzqrbOxJ2/EyuF3FbrH+t4B0Pf9RSaB1BauohIXptljo5OgLi
JBHlJtt1JcJDhXGJvzVkCkV1IgozHRZclQmrCjWDQL82H7VbRFewC09SMUp12so6
WPk3gKajg9AiHMQq+OuVPx5v1cbLWQukcwX08Dx8KpR24TwP/wlfvk9N56QnT/yL
6fuzZce+HUgg7keRDhTAVNvghYtsqp3V+GPGfpQawB6qFp+Yoj4xVyJQ9QmavKgv
k0cCVTxjdnzBIHZnyIUR7C6gUf9moaRjLc6J80UmzM5oDpz+Ji8ewb3k6Y6s4zdq
qT2+qEkNVZTHXv84jT3j7qRrBMLQKXvmE8arrm37qifggii6G+B3VuqJwuUH46GQ
WcFDe4eVCmtU2mojCIv/PbIgFkavAGPhDSjbCMv6Y4uMfY0kfoz7G+/rdATUVY5M
HleHbvMKHnjtXqURLCCu7U8/HEYsETgju0lZ9dY9CFJE9xIS2MktJwKNSL1N8pLF
inUB8cQkM7EL5TmAH5eBw8lQKir/49ruvFa0FUtK8xaEu9QBXiXprri7usiN5poJ
bYC/hbMdJ/k6t0lQXmjMWqWBtLQNflSYzd/vf37qIPCxFlPTKJXiH1eJ0WJffWFJ
62WEH1d3mmPZ8/Q6H7G1pJDVInc/2syP5dJpP9oYqwbWSzKpasrAc7obSFpol05O
Tmfx3YGGpKvdx6FhfeHkjCRToPP5JVTSRRadE5cuE5RTtXR6NVOSMfdhwBs49gI7
XKiU1j7peU6ctv/vsDYKYlwj0rox1pofx/4nSmOG5nFUJZEG8LnYg8OMSa5pvjVI
MRzRaxtASWXFr77sy4/6XQoz1B4aUsSk0D8huycNz/r3PhwQZl4cUbG0yAaTD4a9
w1J5EaFv4BpYrE9HUKMGhLd0Dfqz6AzNINviVj7vJ9Sz0miFIr8E/Oa++4jNEEdq
6CuPpZL3pfHe/wHt+tIYbToN1qnRi+pBuRJa5PBp13RQRsCr6yRl7PgcX+DY6vGd
YdFRa3LL/GMUywWfBRh7rScZqkG78Qxybni6ujMC/r3DSw5imtydLx08boDorslj
irDmJj/HrvtCp5eLo7gLiODgUuXBH/bm3WODhJ4g4XTUheEPjd8LEZDvb6/ztt/A
VIQwQI3ru+PrZoqYS/rh6HVE97CBK9QYNCWZm9SpiPcSL88wo7ccIHqxQsxAXptJ
0fTioCGGC5zhqEHqmI+PwdGswKOVy+mmGxcSCXXI4dC1WDJiSrsXqJwHOatMJhwV
3LhiXLXQGTFj7JmVhi4icTkbpIggWcNDqIou1ALQeDv/WXsduZDsf51871dZgLnS
BYh/Ld3vpAWZ6RGYYng5tvxfI8nMcEnk6p+/BZMfYMuPKltGO0Knpfq8vAlhqb9z
WUOElzNqT23QCv+f5cTrbokNE73kVEQbEdV1z2AE4U36qT52xPO4OhOqhyc6imsB
eSJ+x++4bP7z90SM0egYvrEI8w/RxDse/WlYs+nETdKwT90FE7miDn+pkXlSDNFI
FWA1hq/G2nzOzzCaSnFHQvIDpE/BpK5KLpQHN9gXZvfsE4mtGP+ewWRWS1++sgyg
xTxZpyjvjqGlil44k82YevJ0GFfheAA0RhhXRDzuvzYt7v3NaGBJE+ytwdjQ0vew
Gqf4pB0eBfedAMStwcRo7HsT6jTRpZgEiCNR9ODfQL5Z6F/PJAxy/by3IhtA7NEl
cN61O6mZRORMGsm/3VaTBBkIA60Oz8m5SCfii88UR9NyTyAhq21FlesonYNIkdar
3N4P8JN4eJHzrzFHiwZm1UbRPZ7I2CZngHLBwrD+kyEifiXab/3KNoxOmaMgCR2A
nodXyhx8WBbudpruUxL0IZR7FaIo6sg6ewjZvJ6pT6SzZesVePgrzPUKpIJ6lMZ8
bVncBW2/c9YfIw5ySvEQRrLYcYsRSpskF/4H+Pjyg73zQHSpeLk7eeE1XwwoDq5v
S8DEchUhbkkOjG6p1mXy2+d+mdUUo3PJIUktA+RqPQauWMtEvktLJ2jqUgj9ed2U
Im8HQveFTsU1y/FLpp0JZ0IVcQUKvrlaPQvlMlEM/iy5GI49hjwH4/5LdQxvPg8o
AmJnCZftRBB4Weq82u1+zfmr/q1SCJSYDu1wYwtdGQqK8QWDRENSM6XwdDEME/pU
lYHBBPRFyKkR6sGGW1sLzDZRRj1sIM2AJnlBNTOKG/BFAvUbhSgO32kjcbpGx44x
HDQ5yC37q6pMcr94U6PRJa7fb1a83maVIDrD1b8LkNskS/twUqHw77hXrro1i9wB
78RY0zRA2FNAiJUMfm7sa6nes+hNuEzfKnDX658CJ5UMgFbGPgy6Bj5SAUkCHcZr
NFhocxvlPxZz1cwlKSZANOrNfK1CybYKnOYJIsXEU4YUe1i4n4hnoRmCeIb9A5Xp
Id4/6ethrky6su3Lv3ecLfGR+YpV3ihzzufcRbWRCisgxph1hQiM0refm77ZU6QY
/Sbwp2J4l4fPqnfWM9dGpitH+MGDOniDO522ipWpo3qX69F93m2lhyoVB5vOSNYD
B0HBiyJaHLBe04ABm40h5jLWRgtabVnLoqE+3kUZIrko8u/tHQFStdEvpr+62fD3
72KPAgfiYSKRZKs1SotRRd4yGJyD9qRgxicoMAhjPfFpDy7wBGv0+eTKD4pWT6jy
EYtTMf/H2NotODpcJGBliiSFY0BTauDanmrSC/+ScCUDn8pjdlzCb8GXwhRjo4bf
vj5Xy4E18eE9/zZgkyx5dNC7Xa/AAiGbdXiGtsULACkOKLMDkjrDHyZJA9OgoU6K
d9mEfb/FwS58Az6S2CwR6JL1IQUFueInQGfEtZlIBS+c3iWJ1FsSjYvy//uuYRTf
9fW8PpQmAXw3Jw60glIEaaX6jPBHVmTQWS+d1QrX7qtWOmEo5JuSaniIaMmM7dPY
ORgMithf8TzkxQsiRTASxyTaDCXWlBIIeM7LbE2BeM5orkA6r6gs9E5XozpDrcko
z0smjExs66D9ro/OpC18QXXHFhhbSjjjFNMQYlsaSx7rUXUiJgBL78b0Vfqpo4/6
beUKlNrw60KmPpKjaa6mt78LgatkWc6VyxvJBcGFghvMkZYov4qlznf3J7YTJE3X
iDCeeai57fRU0F7RPy/Vu35aFfpcTUzbnGTulsqzENlIBHD0Euc8qwFMjfoCNZXO
OqdilnloCgejDteyUzi7w5w/fuy3i2d1xaFU4Z8h75OOejoT3tcrxvDrCaNS93ik
9dSynnhu03SZxNKGVPmPdAJhl5yVb7eFElQXS+fEIj++nXL07+X1ZkrIgRebWh8T
JH3fngEhHfoA22/CaRi3rWH9woIr/t04pA26IEpCLj23JIWBcWSrj3LTym6gbms9
aQIWiTXErEMVVOwb1+dnMMbWh1LinQSwcYVa6M1yMxJXT03k3JFMTHCXQx97+7Fj
a96CzI8Q5Uk4LInHH/GTgL2L14IVP7LzsjY1UdOArhF8biGOu1F38NC/y1XXN8bK
eAOzuKxZ7Z1ILzYK0pmM+BYQwC7LXRHTlzTZ/2450+XBbtLcR54hFrn4pCYjgq8j
mGLHA/deAlpRrMqm684B2ZsSjBurSc6rj1G3Mp7/EKaOHqBsm16BqLqhEOYdhJO8
y7BfHKqaTWeCrTOuiiPHzil989OuOHdq96W032/RyY6EkPrDeSai/eGT/D0MzzUA
pTkrsUZs2zPmQDhLWxwVGQe/QmcwB6jfCJJRFIGHb+MhWLBcbrk55d8zWAh78ncl
jLzeCFk6FZ3zh3cbnMNBz1m3yGiTsAjOYWyg+g9eF52s4B7Gcxs+zjFK/U0P8u4b
/I0FIdfQbyHlruoMFFnYRRwU51/4CKtX6oS5Uo/thE/QeiXjh58Ysy3KIIcYntb+
oLXDkm87c4S7qbfieOhPHiw+VWqS/cXkzJWlQy87lhwXWD3Z+6SzH7BCBlmCQTg5
WzcwImjgurUiY33nvWEq01/gWPEO5NdlwtofLYtTyUfA/cThKQvHS7pb6Qrv4DOE
BkXDBdZiEW5FutF6aK884i8Nm//40E6CeSwL2jjgWG81VxWSJRV+f4FcmxdQJtqa
1Ky77MpnPodAAPOG4LVawfcD3Vb2WW/mNLw5a+xNdfhovivtQtu2qgVpnnrPCRU8
yq6nIfzqbEHOw8U61foRgVKCQdsfUsoOnOcBDkxW4iku8RPLfL5lCaeHjF8de04F
gd5B3oBdffln0Zm0OFmGcK0hVT2V87dh1AVPrwEAwVhGABlEnDev/krwYN5glZWE
tUxurxHoo7Wcb0HucZB+JD4dTmGfGTbS+rqvwxzCkf+R2MtPlZjxIDc77p57DSR3
RLuOLb71sSqL9+mu9VENt70Dbd8A2JIfc8rnrUYWn8zFFfePyTCpEmBwisXHsnJj
roMmBNtbsL9XoKaM0LQgQAg/akTKDR1RTkFfEg59nRRgB9ihgN33LU36mZH8PHr4
T3QufPR0mrtIzW276qOhpW8s6+0nzhexzY/hjcYKuFJ9SHVKrTmraRTheT5+T7MJ
utGYhKh26Ce3OwrLZXOZx5DHd1uTEIsxq1zMQPn1JKxBssqNrvhwzZFoBo6bFh2F
ZPYBgF1ey2bePq2LJ7iqsnDzuHxTF/I73GpSXTW/Mrr0RFUdoOJhN2p0HqeTm2kN
gCsH39pNZVxr5CXEXoaAXTRbCp7AjhYVrvGihezUrK7s8RZYf+mcrZhYGicYug3E
dOZG3dhcXTSoLsDFIT1yqthW0Eyi65EP7w74qMcdrcBmZtCPPdvASBVoa9Aw+fTM
Xn2V7vPWPQBsRU1+Lthdjk5LtLEXAyJ2VWgVrRigN1fP8lk4ICH1DNWQHDS0kVTM
iSAAGJ2SA03kGWBASjpwgXGuAUikbhcMIvwRP+058SG/0tjxWUNSNerN3GSC+OW+
7mqWYkWSpKx5pNHKVkOsB594QUTNsFMFalJ9vE2Yr4ZQnaJBRnn2DxeDzEPdEaP0
8E9hAe4mCwG864bvDvvVB/eNCpQPXtrAqwOpD1e9vrqafEfCql+LZar3XegTHplD
6NEvPlz2Nqzq1oXWjVWJVPi6jAhkF3uLTH2TL9UZkBYk2qYgBz52O9KAqz2k7BRP
yMkvi6aIVg6Ju5oUpiWcH0bhY4aI25WFUD7wtBjYJ1JYt2LH7bGUsBA4ggVCH931
JDtLfVMhhkdbQ9bu0my8bi1QNNcx5W/VQiFNdvo7I2W35CN4viqkdDOBOHJQtp+q
IXtJohb4hNvwW7HBNaoBmoqK2AEJ+3rnbJd5Gv382f1h2lmV8PZEZCHWwNkHDKbT
U8KcMx7erHOROUcwwHKTMAcj87yKMGH5PBrtsNw+S1MKbSR6dFeYntynbiWtMhGd
82cdtp7lgsnzC/P8qgEQU5QRUfCNFZTBfqW2W4OD6XoS5/oPL4xQBXFWfHg5Z6yb
20LLzf0Bt6CDFXFUE6TRvhO6e5AHUvo7efrKT4TTHRhLG1+tDJcRI/okJpP6euLc
9iHyeJF/FdjRy8AbPMoL+izFI8UhbFm51iFuZHbqPRFO/rLJ6msyJFukuQRqLqvK
kziOyF5dnVR4g+lS0luE16v87EWWCikz3hVpUXYvWPHmSE/kSnCgVKVLQvGLH8eZ
djjBnOfDb3fLbspfqS5B4qC1vLyV06npGHVPnQvfEu3xHWQIHzSax62IsSpQkcA8
UhIGpeEBpg9+mq6XWNaB+z939+wqzJusU++AJGDoFSHiO7R0t96XZiKb4PP05cGt
BIgpI8t2QjKwM6tEbyRIZC0qdMnUUkpZ0KgT1sKrSfHUtHEHd+6oRmdiKgbGRoG8
/mPHImW8QK68d5XDDEVRMPuGhn+hinDQ/Atlfxvp5RpEIPX7RLQB0JAt/S0dO9DO
M1oaTu+sBGrweH7pFOU/JwHYrjzl0EL+VuCVA/OUmO3l8Kq4Xnv9YufZgIreXgKi
eSOkZWp0z/a0+olfq7y19tE1w6a4m66W/0HM24H4qI2pqbqoVqmOtnWBuo8WHPUm
r1FXz1lLZQXINj4O0fkrE+KiZmllK/lAAEBTQDPm9vfulnxlI/VDKSA/ooCKe5E5
qjBZ4yhP/2YqUQDA6IeHpEXLv5MvOUC3251daWZdamPEkcmHV4eM9bxInA3upZYr
Dzxp/ZpjHQ55RaCqWyd3Rh40aj4bPLYe4EwMz1+oACNWJPqu3t/KeUJilgbHj7Ht
sO1WnLCyDUOKYflh+OwqFPWqODredlBNnul1CkFZJNR0QihIICN7TZGQXvnM9w1s
sD7AHmBKLbkTH9KXHcTa+JeZ6nfLP7ih55l5TvzixzEXpvreeEbqUG4+fgE9uzkd
mhHTgv+AmAhnvVmR1sBiksxibZ3jw3P2rvdUoaBb28s24QS/wAeQHWmfesBVBVlv
0pD+ziQAwyeMCcoKsqBEDO7539oYbgjcCh7UOEWYZelYm5am9h/SA7RW2ki3rNcf
mPu4bk3lHAxOGq42+4Podw2eORPa82RoaAZex1UvAJ8AW8rRmiv6i1T4RqC/VvxO
ZkzGSimFnxczWvvQyJdZpxO1OLHpnDySHij/BOzy1MHybXGY195Dwh4jvh3CiyZq
Cm41lFhgU3cZ+Oz0KuxqkgoQjcRwf4hbopha0qyxaARFuzDOzSU68zn82zn4bP00
rczhtUXgvydXNyAx/dWqUSeEuxj7KrI1qKy2Nya8QarAXObNrX8d2z45nIe0tQRP
LG+q5wr3utQN4W+eBp1oVVC/lIdSrYQ7m5pX7/6FpHo0UM6a7zZknGIe+rcTG5OH
cfeJtvTSTGlji3bsU2o+MhXUKxBF73zfgY0KiHYNLki7Kd2G60UiCK5gsp+OsfZ+
ARZOyusHGd6UvkI05N3jVeYyHPl/d9XJ0SiBmDynk0P/Fwxpm5AOzKrO/CJYBPal
8UaLlEzucfWaxmabgjxIUhYQ+Y6HzpKo+nlpGfLgh7ASfQQAYHsC02CALfuojqDI
buaL4APdK75motj1kaadDhURkdWp0Yn7egXRnl+Ay7iOm8G2+4TYUboNTAjnT/cs
PVWC49m3HwUc2gD88LA9vVx5iFSpE0s4p0T4LF51ozcu8EoiNrtd5Qld1Z/hGtLe
5IeEJm8DqxX0d2LK1XtNlpujW2jCjh9vIAxdR9A4DI9qCJKMYaK2EuQ/pftocIkO
VsJs77gsbxu0GhiuS0/BTNLJAvSbRfeaoN8F9LyUTcS8fZ3JTWArEVgbf+OLz30U
1uVdDONaj8XF2XKYbynM8u3oE1IADmFOsNwWZLm2LPSSnAPPhhcWiheZG9lZHNtf
2CtUZjGR2b+NhLz/IQtWowVMQdhzJZhJmIH66Dm8FDvHTShtZEKeoY4TwJiK+nyP
Od/nPHzmhMtnbTyU1NWEPG2QeRbSCGgwQPNlKjoV4CFPfOLKzM0YQ9im4EdVnUjI
7PshG2Y9jfOiu0Xd7eFOiK+qsVsiEXDIb6hWgu3iy98/2Gc+2jhKj3h/ku/2LBi3
et5VZ/sziQ42d6m3R1K9fNrV/Bc62A/2Yid9kMPQMzJMGF+cexZDs/hhgv9RdvSC
t84Q6+1coxDj5O6rEssLUcF9Lx2siACpQXeyC1PcfBST2rbeEA3/oSPpd7UbO3o8
laU20GwUmtu3kmRBSPsYemuk+INaUCHo1UmgwTE3k+sJMAbmXPys6ffn8WrYF+sn
RIDYxqRcwgg/Vrqh0EXW8NugIEjBQNWgwNPmxmoXxhusaPuhQJpF7canBaoz9x1P
MyeNZ9XHBXyIL+7w9y2al5rdvUS1lNgaXrKjUjSiOFAoQzrP+zY0pzMSR8lK7Nk9
O+d4Nk73882uJfDcyMwWBGu44CEJD1Z14ei2PEv3evpmbkm4OjPew3R3JK6BLQnv
K8DjRFYXkNuWTCgZ3h0OPa0OeY6JDwC0CercHvoL4OaXbz5eBD3tbetb4bLr8EQI
Lswg0G1aeFAV+JYYbezve3ezcDvspAAqrOGIcLXKOKGOgBE+NerpeyJQARRlFqej
dTQv4IQNapdVjZLhoDqL452AK1UBMSqEeRUiBxJNTZQkccOOQsFGojgdblqzrWyX
u7bxHjpQmchiVzZzzENWaOZFikUJR528yVJh42mwY/hcsTsLRNyJRNbd/vSVXb/L
Yw3UgCAwmu7mdkC/l4LEqhvHRxI+UH987bApVWXO7bedM8PwYvaQCb7WBQjVm2T9
aaWp/WCiAiO78A+lOUDfCYzg6QoB0QxljCkCRCQ1TxfdmPak1nDvk6yMGGSfUg/h
GCwCTgBh5bkdUE+tdAUhSJC+QQJD7rYtlsu3ieLtPv3ovEFyaOI5WXOocodgnIoo
OpVz6Q2OsyCnAIDfAbSbgEt3j7aukSwxzHzFtctA5SkHwbs4l/heu6SnE0Sy/ysW
JZ0xSVO70z/FAaBHf6HTiKLR6jvZI2Eb+R25GDqBQqZD6cYb3x+edkA+4CPXXIig
ikHqMBR/ykzyouHQA0SEzCFRW4mojDwwEbU1LJlKafmH3zM+Hu7lffutTy4vYaym
DD3pfugARpthbGbw2sEHtWx4yAejp0ybFXcgYVTEZErDAi/jMTXzao51WIYcNSAx
1LaT0xhFFpf7M0HPrunJUdL3QrYD2fmzeQz+tsjL7Ewb+veATIyRPsC7VQoB4HZS
HNq70N0q3dZZ8kIAcJRQ2IGNyRNqVbk3ireLqNlMSGCEQcQbwnBoJx+zgsL7mtWB
Uw5+HU10pINONrCfCFcaReFi7Nd9K1/zokc1H9AMgrTpauHmaO09Cr6y5BstFJn0
axShwj5J9fc4ZwnZ3GSGmkbjHdmA3ko/8MvodL5kmVEubgZkhX/i+WaoHF3zIgcg
2X3zE4vrbtcKV4wfKRaqQvtb0Ed+5kxQ587ky2oKYvLnJAa0RS9fA9BVaXBXpZKM
tBasXheqqtftzmmsJn7BBNxeY8kTfs5eL1XAOOcpBxbvlZlj3ICzgNLF4Zwwsj7H
610SYkTTblO6vQ5uGkHtMI4THlFM91csbKZl3+wwWiX8o/OOA35f2KgCIeXLSw+t
YRi9VdP7a6Wiu2HwCFRKkRvncIfE5xDNoYRMOKGFNs2JeNWZnOndq3zZv7cqpUjh
6d2BcykrBROBoB5SPhmdIWb5gPaGxqmD299KCPoXkKk4dIOB46fys8IXH5kdUS0X
pt5AjE6BBLVu245UrSGaZuSlEGFyCx293L++oL/E9fn+GuEZhGkQd6kBARtQUxmI
KSNBbkQYn4OFQjVK0sYnG34shPo/JPVshL1uXwTi32MTz0KL76X4JwwhH5fXxv9Z
UDpAxe1AsrQiD3PH/7/KDDCgOZ3Jwnpf4V22n8NTw62MViCtJ5fuA5xuSJKOEK33
c/StnRCaJKiXEyNa6/h3FnhIampHBIv3/pU5sY2BhghdqEnkOw74fMuU44kxAGZ+
QIKMbLhA/qpeAzwS4VPQ6goLTpz1EfEcyE/bXgbORMSlntFiRfXSVla3N+MG9vga
R5iMdsrt4v661oHXFxRxXlja25z48xFaYMNRnryjWM4P7zlhRlOX7oHYgwxEU6jg
fWv1l6Q7wEz/E+1meCaOiN/lLm/FO8YO+XMnvNCxablPlCfpsO7yttcj4ZH6kNw/
DmjA8zQJw4Y59ZoUS1JGZjmZi03n1cxkjnTLNb2/C7Adtd2BWSuJlUJo4fVv2hcD
x2hGSmxWVwn35oRpJobAzhCtE6pyrS/dgX/SksRA39GsBxDqne4rDeE50cemc9Pu
AjfWoZ0K0vEWARPnwOVnDcOHLhB5zbXpbZ9ItlNKXFgWTaPB4IV0y09ELe05nPn+
3O9cpX+NgAARBbj1RJESHfUlhbp3Q54MnW5yetBLFaMoy/rL33CYoxzBrzez940q
437CbNdlAGfD6R+iBb+AKO3NJlx1+qRD4JaOSmuxjdBN+gYm1opB8IFyRXNL0rKc
0bUreTa4yMsytu6nv2Imqx1mQjtnxGi25sAj2Ko8gf1nun4dOxzJ1HguQDOrkuQC
pV+46/K0dKlcJIlZPPbVWvlRF+IjKSSUc+4cHTBoBFn/GCEE7bcs1pcCmDz7Fwc1
Z7NlOVyJcBEZ7xmAUGKKRjRWr1yHYC76QfcbNhaHUAGbp+vdjhHZ/uN+yC+go+N0
KrD+tZ4MTt4POTFBLwdu6JaWK7uYSvNoIjrvRVhHtI/LoifONqX+AaLcJAX3uejJ
nZFBW5EGWawIs7JruC1PaAqshXTlk+5KvGcKMk5Vf105eqmUmssBdcWv+Dpa14AC
JsyByYvFhaWUjhhIWFmFlUjD21b6quihMKGQxScVj23jP0kmWj1YnHT1EHD4AYvH
yWqjk6K9AWQ3/8yUC68uvwOyM4nQc1FcIKWIiW3EtObUqDUNSyCQdnhNcs+H4tUJ
pfvEXBv2UHyvq52v/guBPFiffQYTqbSBN97GvpBUvfvRA38VJTLZXdIf/MhPTF59
gYSnMsN5xMzDVadUh9aJly13jOUzGKdjpMIRqkH/2k9ZJ3c9PNtkBEHJLTY1e7zz
0YtqWuU8XOpijDvUtkDXJ1RLOZgMHMpEfTkjDtR9S4BRBW0bcV7VSt9rRbCP+1Zi
bCrV+q1M9RlKD1wgyTne6IQbhzkqkZm+ho64RYYnXNcZqPBKhDSBeLqQFtzgnjHk
vpEel7SgiGcI+DHKBeo+t8hpfJS1RKf0C3ZgC8YUwttMHcLxzNTPdX++5rm95Jv4
7EsZDJ7UCwD7Pw7+GwxN0gXettsSqLsb+JQGnVi6l0x+HMUcT0W34VjKtD9AhNXK
dLyDpcLSItkInYO+wEnxxl/BtwtKFxeqeJutm+K/yQIWYoG1KHY1m6C1Fo5s0sD3
1+0wCz+jZA3YYwHCJRLYeFId8oqsoi/v00/dxyuA0flHEBjRWsv4XCU5qEdy2zB4
pFVmFdXpMdLwN1jjnzo9QZp/fSGhv4vEZkhakqeKyfYZ3iZfbND9aaHssl93EX8N
2w/grBhwit3VPrZB1CmudfdIr+fa0H8vAlLtC8eHrV/E5MRKk3dHKc+xGJHn8vJ5
KbMqfMn7Ca6XXuURJvMGPKOeuFGe0oU6cN04NXh42ZXqIofFTT3n1mQr1AakFk24
Hcju+VW1/o43FSESbJs1ekbxIBcHh7HgpbyTbUE95b4WDG72eyMsz4W0HYliUeXZ
GdSdjvnzJtWDDHCIrxBN0WXQd6e53/XIQnATTICYLCMoa+z/Z7LG827BdGlxHbEs
v+udmioDGC7E8cVKxgJ7To1GjwnDCj1kQ6oss8CGutJIlwiQVHfDIY5lf54DaP1u
XyqNjGoYwH2WAlFczt5Qnfu98IIuyhb4DgZrwU57v3Pzn+dwj8luKP4uM82xX1uf
ZscopuLimPDIjkHWRKIGTW/nHLN4bqn27dbG/b+sjnnkM3JSuHK7yTXaMeVplY1A
/dHUiB2J0C3zxSuWqu1w2x6XhudwWSYFhfl43lSkpqthvI4/1qSdCYSj7jPvLeXL
RM7QhbtFTzKAuphDl/7s5ZFAag8exqoQL+dxsriUe4iILOg7fDfFqhLm9Jx1lnB7
16GzHKNfOU6hhCxPQ6DTB2jfQDG5gB5gVutYtwawcrjz5TVWZBnDOWq2wby7w6uW
FKa/UmCRpThrEN2upSqA5HfR1HC0k8kvCB7Yo/NlPFocLBYwISfTDPov9uMtBTaH
dCynSjjqqbWWKyXtZz/XNXCWBxC9hP7lrPlDWc3QBCxeOR2oIVfom2lFy521K1xv
Csire6vd1HDwUIAtu0nOd+I/090RIM/sh6BnX6a/74Fl1esB7eGy3DL42J20koIX
lmApREVuwVmAbBAb/bZuUjXgDkLue50Djw0rERvjrX9O79GkIg4KilgAz318o6Ba
Gc/6V1p7wyTYjjaWEQAFtueTlg7QWDP/4QhqBM2kCFLxryDxCqnmARQOeNY3y394
HTC08aqmkoRysawAZUantNK1xHN2pYnyZv3wv3xGohSho+B8HwDnD1hL8Pyko4X8
j0qTsvgcedmZFd1dgzVwXAtana9DfBDUqlin8ddPuu8+iaDX2YYMya4Iz3QetrQw
0EK6Y5LtwkQ0agCxHXrl45u4rCTQ+NmveTk0ar5bAcFuTe1clNXGqqw5ZQXwAast
KkpfwLWYURaBmYf8W/JflmF0ORyqJrbJq8FDGiM+wF3q4q1w0O/0iBlOk64V1ttX
Mh15QLjr2PxyS+t1d5aHq6N5Zq5ov4n4FZUNIVGjDToYKq4D2PVRYQVCD/pLBVle
6OcYEmhGL1OqiDlsZNhotCTbfY6LFrnWAbuZhTjDH+iNjLokvZzkBGrBaQpBDuaK
7XF4TfWCFKNX3yEv1nY63NFnJT9n4nI/7Pj4sJB2bQjaC+7zmNi6RDBE/huzzmnP
e8wYp1GcTNmBNok0r7v6fhbKysSCvVeK93vMAD+U9WLMrdcXEUdubD0w2pm1TcSq
t6odZ5FTe6Bfl2lgP90si2MsiXvP+Q+lDuhz0w22Po7IL+NsJinUtyhpKZyeNfab
Xscs3xcrmKX/O55+Oy46kVYfMk7uWy2EuiteqLZPLLLlLfsuoYn6zT0ODZL/1JY6
uC5DwE+lO6sVH/F4mEqicE+eu8Isa7I+52ity283SEI94Rckj2toZXqYQaVK2XDF
8MxWOt/ZERgcHxClUnGnOBLciEvLwlcQLtolAvyH1xGrrydwxtPMGkISJ3oEYxCL
+U6pOCgu9RF8fWkQHirRROZ1au+0stWmBwOoHbvfFjGHyI+X5mSuhtKjYOY/XbJH
QYM/V2SMwEZjaAaBTeZFDxvw0qVSgU+Qg1wxJD52sQrCOtKN96LdrHbj24cKuiOg
/ZFV11njxi3aKfmp2UO9f+hSYh6SzOC5mDsfOutHPp0siKAFXcb9HY46pzeNGOzN
pN01g1gn4H57/TGYBl8NKH24FJlXV7jb9CBt7hAv7IP2E/qRlyXRknikztMjcJDC
IK/aF3ILvav/+Pg3Vqawziv1fv5NO//g+t5UzoW+xkZWNfOHN+wnJo+wfqpaG8Nh
4oAMds4jzRMdcpT+Rt0rxjwF085VFK1BASNfXODY5CLscTUwg96RWwuPQqGyifRN
pvXaeh+lBy+MeWb58qxprRQCQJzbwjqtftP/QCUqsvaxP/QDFO1DbOfvqb4M5zy3
i2UqUmcGOXqVChtmT4NgQAQK7gCO07Cvo5VvXJ44rh7WvQx0XMjsNoxHbXkYu84Z
pJ/9VfaKeX/vkRaaKWKBma9eKzSQ6CBKM2gtSh5OznvSz6W1TrLpMYXK2Bimuy38
78O8NL80u1/vEcMx5nPIAfQT02JaJSa7xeHuiTfluK5Qb2/0DT0hph9xIM+pzt/X
o0j/ElKvAvGoJkpDGgItlTPBkTgWwrIDmattvDbyF62sq1YbGZtq171yL4Wat6Z9
Hkts56HE2180KLqmr+IIJDSgnpBNydcaXhoX3oFu/qVn/dB10TcFNLccslkCsYNC
+HdtHFeQIZ21zbyelQDtpbxsdpoz8yDQsb6trabWg5lOP7Y60U3bombTL5miju80
DfNqjVvpTEw6XgIqdHY81b5mQfGyJHmdaN659zWUaxiWixMIjROYLM/wSgMFu8DW
zsmEoHf+ZDtzRHXLkSUPhiF3Ou9s718eUrtgxvF/UoYl3gKoGTQvXDToOrnQ9YVv
x5cx0UKm/qhI6/CFYmwzzf5hIGInFeDMVa2RuxN3XaRuik6fP33VLblDUqV6o5o8
bK5/TgqsEbXLR7eIAx080CgUUVBIOG6zBAiJ1pZ/0/jnxx5n8YFdaecQazfw/dSm
J1sygFXrd0Ogu+O7Jh6t79obuRBXcPDwmtAk8Rwpt+NC6PHvLNeuzHih3dJOCE1t
zP7CqRlk0ooCYgpYPq2DyuecUf6hdm9mojITx9nC6u66eBmwYSMSHFEtLudXwZxp
SNVLAa4SiW59MYQDoZQxPEF7zdfWRNvjjSaU+4trgvKMT2yGBIkkk2DQifVMVLD3
E8PnVI6iZRJdJ/5OMHyCF0vf/MxPdrso2RQUL24g4AoArZ8Fr+sgBF5jM5mF+qNv
Ux7F5bmwxih9GnSDih+4dMpPv9DevZOaVuCCG/pk+0prGRa0Z6zEcbnrqM21VYRg
9/anTNaJh02Q/gadE+IB/Tq87eUxaJPDZfwiZeV72XECOn8T0ns7I7v/+Zau74LK
jfRtlMz9kY2HJNZCznFaUe7g8j+bAYkKtCBattNWLoLAA4L3zfcGc/1KXcU5ZwBT
jMkFY3XzX4RxjOOm6gq/OzpdsJV8Rj06DawERPKOA/ePAEwPYjqosUbLRzyklhEG
I5PYvcLrPcmTyaUZnnWVSrYdUjbOGOc1mmk7fsLRXjwnTuEjLmtam+elbgEt2F2C
zKTG8v2gRqUe0gy3okHO1iqp2c5DcGG6plFLUQ4ae3R1wqRIc5v2sJA0Q1yy+cmt
pP0ktV9NYYYasC4eyGaKaadyxfGjjYZZY2VizgB/xTtc9r3/r/QD68Mh5lJRf3tb
Oyw0RXSRU/wjRCqNuxDpIDtb+u3/GEzhK+sEU8IrOQ/rbNuR9qURzVWLKiOGuqXO
ZAXoXQ99+Pj6tN76h5PvC+cLf8FKkoUlsDptCFeNVwJL7ujlMxca7hqZx4aoHaI+
ZThCooQ9MxGVbV8y+2gkS6/2ML2spmF0STcq/UbHxSclFHhExYf+Pb6i+U05qRuV
ZlYrfx1PQXVgNG7CjPq/1U07JFosWkIu6AiBkYumMfu0A1J3z1wswCVcq9vCLxD+
ybNdjHQLbYe4Pwg2dIPjxtHLXlEim/CH3AMrBnJi1Z2LTFPTmQ0jkqIturJWhOou
muTNask7jWOosW7x5M7+EilHAgkmqCFBSWzcMSPnWo94xxjnP/lRaSDIcF5/o2nP
KaUM6M9HXH2EcTryKZNwMG+DoBSOEKjdVEWz0Xm5t8XZaK6lBX80yKuCU8mt5k3e
OGTiwe7lb3KpzMe02ze/RkfqitYJQNbasDabcBuXXMxofHYKZ5Udr771rMrU+Bau
/nvMqo3sb1qrl6l+ufANGxFO+nlLuaEHZq2U0ubECk6AmZLDHuaTsHItsojoTKjg
CWYfTUaUwvYl6V8VGEQd4PSR9onKdpTMQmxAblvmhsbhqJF80eYznm4zS6Sh474G
nsZEfjuNWRe5eRoOD2v5vSZER8wJTL+MHhZjvmlIQOQsOVJ0FMovtUyuvTG2iQtA
n5iJZSUuw5Yy+OsZ+c7cOitZeoAYM50th46UbMMGxYaeWK8C1xUtGIu/TK+M2U/3
eFfzqgQzGJpNybGI7/486trco24w6+OZYkkyleeE70Kr+8tTkJfvvOKwcBHdb/ao
EjSPWSw6x8cB70M0ul9MC230pJiDetl0koL32raYSVENf3qnDCrBTu2ML5zgZVHd
9agsAL07K67nyddbr8jzVTzmPUXEZRZmya8F1sm8ghXAgcpB+ZLXXTi978C39YcS
QI+qTGxfH6xYbYqJ1DLedVe5qlBOqGeJprrtFWMlGZy7VP3LHFcQsh1+J49Dl6+A
2+9y9QSj3GZIn73g+a6n1kAdwbp6IxSXo1U2Hlt+UKN8WNyJaMBe8qTxHVF8dxMG
0FYK7Osni/3sD0fCnPalySU0luW1hlkXhHQt834upeHTErE7mBzf+NRRAxZJonhC
BLPIoF18ppOhRlnWE0rrYNRbfCEVDCgUUcMGQsjpbuOzQ9WdrzBbMJbuXdt0ypR4
FudQ0FBjpQrbv4gh7UnZy9PEzVUW2AMcyvJq5X+28+U2XNKBnNTIXwDqnEPdpa0+
du4ODe/IjCUs+j7bXi+aeHyr1PKvvRP++EsIwgb78hcfILC0PuQSEsrDU4vx6/hi
RyljtztC2vx7O3y6WNtiCt/LViEiOAv4/wjqUR7t/ZI/7TCjFfOj+Bl9qsaD7FhH
K6Ifqhpx6jYCWjk+6aWWugcX5t1+YuNEi6HeaJM3VJrluW38ephApugAGZ9fP/z5
rQJNL2XhaMJkDMwaxXyFfm317FhNl8W04Hd9em4zYOYwQmDvYUuTdBQCOzVu5bJM
ZagMHST1k4EZk/+k30xxS/R4MtVAJxZEhiRuNitAQaOIBCI8/G3EZuw1TaBSe0YT
nbXXOpekcDDVY7RaP1JqAG6a63qp2LQcPRAoEOpzxAihZAIp8ZrfpajNK3bv+0Z9
a8zWB6aLALuvuZjbUVhE9R9CmfU9hgVNExnACeIShiekcpA5KZp+EIrCd3Agf1w9
Wd908MwYkQiLMU5VsJiMrRPXR4mi+h1YGw1nlmzidyhFdFzMskKFQpJiQbgPZjvA
nI8LZ2jOnxV6VDEyI12Dk6tfgvDtvvUUJhwIiIpUQIupybXWrhvnpvsi7kjxMH0f
oO7FRD3DAOrAEYz8JQODVPlTQkvjguF0Fl/EXcZ7Z13Xej7KB6PRxE7trL+f8c3w
HK5HdeJoip+xIiKZn3indCK7vLfzh1XHtb+NtTk5cgT1vviC60Hxlit3lLRKq0FW
2bnCBQaIQd5Bm/Um302L5OGE4yPsOM1biajzIz0zvIz1tyZ15dnCNYM08WjUJ/lN
HPpVcX6sbEhbvOmTFl/mr+uNt1nSdppp/1osUQdek6cEK0GKKIzBGMbOsYP6xgXx
bE+omTkhYe41o9QhvA08pNRwjzbiAqD8PIQOAuLwENHWdiAsVQgMvJ34QrUb6s2t
Xnq8YU6RVvDerQRLeZJ/deXY42Yq9QRiG1zX8NVzY/SxOMB9+T0bRAdv3+A5EM5h
FVZ2JVZJiEtVazufKsNxYpA6htgcC41LCjb90Z0u3qJJ1E8hQunLRrzUrcnC+QDF
9vrFErkDxGlwi1mMr1gQ+lFjshxqeOZpaJnmsw03wxCSk7/kkHETkZ2anukfhYG1
NQQXBSepPkCQovYm5HcH/isX5POtG7FDHyD9v7yY74Ddheia1U5OeN4XqPZc6vhK
wDiq/bd48Ra+/EU+WrpvxfoYqtXSfkedogmmjDnP8RLPvuCGceRaICJxd4/KAQgu
Zh/NvIKICr0ZpcSoRTI8nOB+D18HctzRofEJBafON9I1ygP2hiY8ImN6LwPjdIIy
M8vy7/jwHb2PneMg2M3ZivTbabpAgQzZU1CSO7G+67wOhboVdcasFiRFzCRricN8
6jVM+vHAFpETZipCcEAVc/1HLzTSbK6wGNJmtyQkEJBkAMIGeNPpOZuSk6CKU46m
us/uApgTb2BouLa//II3XU7DMa7wVzeMHxcPZCb0AkxDMVUM+V6o8jDWKlz2/eKZ
fDl2rzguPeXKKCZ19jM0x4tt34VE9KH12FdI3Pg3Ket69N7not/ogS62N7HtiMoi
gg5hC1U48Zg6SeO7XTwQ9pNVv4g1dXVTrCUlvT3X9j5Dn6tlOO50rTGZkyuYPKS1
dO4EqrFNvyqJsGlwbpaFrue+tOxowf6s8PuyQN9o9CXIkT0Jx8EBK4nsd0us8yvX
vAuG5kMJ1P+ZoSoChvmSheaT2LPRyTwD7rHV43QJYLb7ajuN7K7N5j1GEBuPyUwk
Ffl7b4KRbneaBk3Z2fc4Oxa/V+/66/4JdQZSpQP/RJqC6irVx0169zO09NTjwcIB
mfpVwqhN8ImJ60InB7REsOD7427pZerXCjYQx4f0JGgc6iM5wdrbQM3ku8T9sDT7
55XYIcyfl4sdbiIpR2X6V/Gcng19X9/m2Ex+CR/GVsYZd+TR4CUBujrZowQCcfoC
YuTvnduc6rHa3mieX00i3mtZ/Z1RaPd55CoRUhRAd0XNKa04fNXRKh8YO82aqiz/
VeCan0WqyE7/0rszAInnsGghAG/Fx8NXMYyFkirNB1lqh/pkBhtf0Xk9UTGfhTLb
r5bNUdJDaotdKnSbLa3L0+iJwzusllF559ZygnU4EhDVgMus0yqWsXPInchGGc7i
kkSMe1mrqxdxFMVnjyp2TIcNohtUDeqQ/O5DHnEo9NfNHDdZi58l3huokZzjm1/s
96wZyuZWP48ZxL/7/ahTS0apT0hz/E64M4zbFlMckUgE9P0TVVHk5WqX346wsCOc
EFuxiDfdt1upgqAHtsIumBCKjaaq9hjuyprsHEjO2rEFLqvFfmiCG/8Ls7KKwrL4
fXd2w6K+66uvfmvUbKcS2GQMQMV0AWReDeDBskmi7ILuEHyQMMm0XSxjS6470S/y
dPvwphrPcMzbyKwSj//h0RPBVg9HJuLGScRU8AxdNJX1b79pfSqRgfIau1pzVXDT
0AAxH3lC0KcdtmfGdpXWE7cKE/x3poLwBkXCcnhL7/yt1lcBQtw+mgvc6NljIVKP
sINiQisUUvoLXH+ry3yP8dp0c1afgw9MPBg8KIPuoTq40vVsf2RL97UOvtuBfXzM
e5VW5LB6Y+98dFjAQacrbf9IwlwRXYPNjR1RjxgBqOSWDZvU7WLjsnt3oPwz9zoB
BDZtt9GmpKNFsrVH6bQck3A9dG0wMiBps3CDcZCVdHL2PxvQ6UQPfdFMyMa9z7K4
HRNtx4+PamnS0IAFlJagDjW2U+HSKS3n9VFNvj225ZKtFGEjIZG3GbMaq2e0oZ3U
BCrtbnkn8zKLJrfl1DtAli373f1Nsj2WoDE825/eAEXykYeBHdadpIVdtBz3wxhc
m6+JZslXeyOpQayuMfLNs6yu9kOlLvjx+kRQDeTM05SngITDzlJZIpyl86bgPGN4
WYEhC55MTTwhME1SBr2iE3Z+lwnoz17+6GTBMgRLINMw47GPTvBPklxtuIeNJaQN
tTcP9F+5p5IizrQdFRqrvsrtJDu2TfcKeLlyYyAhbWIqYak6AHCiNHg/UXNe7rel
BhgoDzYIqbFiSKWCs0h15XkgrTyFTxcGvliSMND0iVsBEOO8W4E9546PMITTY4G8
ao8frxYa5Rw1vPCJhQXz4uPREVAUkCF01U6pNdhSH6fGq+CXj7wRu+XobcvT978O
huXCGrSqL/+i1WJeee9j8seT2kIbdfpTzmK3YVru1RxsTCZY+OQyV9u1749O1/pN
aFwyG0PtQlS9hRpP/bfg4krs3MHxQ+A4M45vfmRx6h6XVm2vs6Ja+z/B8wHCJDDN
IWbP2hTnAn9Yf/2nkRe/Se/cq1OJaMtK3WyGg3l+wYEIsRLgqzWkG0MsruyMYvUd
6FuISriaI8gRBqDCfAR+rw4Zux1Ooiu7ElVn2Mljq5s7fHSj0AU1RML47VLfDg4x
1WhEXraKkHsrdb4pBYSjv7uvcuqtqHgRgpl6E/BphTXCy4QIKP8uZ/vQaFKDIcK4
vqT9vxHcs8ok8i8jlxXdJrCYfHNWDVF+e0VotP6bXGqHLxubIectdEiXFlFdEEuP
aco5IV6Ly1R/j3m3bliz/6LFxg7qJk1O3zQkAFPCuDDWKyN3ET07dKBMq8jxtDmk
RM6wytDz1uTwt2bSx/pq7DkU+qfj5gBWBHCe2pL9hFJpix57hPrgc9BQr3BzT3A7
boh8u0wlPLAyPswRVBC3zhgYYpMPDa4xWxYZiPgJhquTfeE2tLS4HN6vQnCqqNRf
ICtCA+6bcCy/AD066qdFKG+HYkDDct6U9vkhtz5OADUF9xCl15LX/wJF830UOYq/
87j5/BI+tbr/Uf8j4xrg+YrWY/G4Ljlb5O175R8sWUvS9ymHyLAfQukeePWLwoLf
v+U6mlf4+KZQzsweT6tjmIQaTD50PZySak3r0vCKdZWZgtD5/jTG5C3n7vbLk7b+
VZ7UMC1DfQpTuT0mZYsjyARIPBBGM5nKtBlxlLf33XZk82mn06tYI+z7KWaZFedz
/QRF5Wg3QZ6pNKcZuCQoXZqnjMQMHM0eWkRkTv00qTiS+33ExJ0Hd9wEG9JKJbu8
fVyMLtAGXCw2d3crkf1bpXc9MR6Es5nuZPBDdZ3BbyBEkecJJBOiroZY3fsm/Hmb
MZY85ghjGb4m4rLNnJP08VUykV0B1SLvm5pvOigeDY5V5W4X2UVjMgJ3/yKRO/4r
FLqLpTvS0SlYLIiyrGV/Imkrbjxf/L+qNIMCavvFYYsJsQepNYXhPsq2XkLV0haZ
kecaw58x7NNUyUJJAbqViApM+ck1r5r39xC1Bxv+WHEMm6zeNOZpb9bZRZm93H61
KsQCgePe4aH7Q0HLzjHNZvNgFRiTjHcF46TNYDAWlI8dAbII04accmFHOJmbL6p+
IsA2EWD2XqYcwGIWJqPHCWdpegHGgYmr3eDWkeTEwLGjh+YSQZpi1sQMHDXc1Spl
+47GZKTVi4DxM1X00t23o2J0QTJSfRwGAMnbTT14zDP70oaBVmPpm2Q+dPWNWH5b
FBrF+fabvroyNWKZRDKhsuZiijyWMuWFFw3HDKPQPK4CnOe9EXzPusV9phxm85NE
RVsAffLIaM0xCP8JaJ9bI0ne91SojrXMUUfbMXkJE6Z2I7d8hGD+D2dfo8tKQu3l
ESOuRzOqorGFTVuz2Euu2UAF/mOZ1KmiP7mvFaLC1hyvV2kb1o8+oKzMPKKQipp+
oDdrRrXYn/VBtrjJLSLKe4qRbvJncBDspDpLjzLr/p1epJ/qJMkfJGhz06fAB8cI
oizZvhUJbodeQj0nkLXS217Sb3eADO1eMa5H9U3PKsAa3+oVlnzyrDYIdAcdiigy
QjV6bOhNbpCWskn+kklgDpTabTM+Nt+CVwZgx03IwdJ+ouLnJr1eVnPdN37B7ER7
1H8IOCmrviqstSqbTYzN5JpXrTi94zMsLL2QFJoelCNY1p3mki6rQxbRnFJBQ8jF
CU1AgmQ+cHmNHmKXwOTFMj091cq0h76ezaUhwUmySVQ2R81km4QFhTWEM8nYKrOz
cq92QHqgLhedB+uI0Jym20WGq/yVCZ/+mrz7P/XP4le06SyC9jttqZHdob51fHnG
+9m9S7tEvs5LEF7phV/ObhksPia86pNy9S8TPRpBOnhJ9lxBvDiT84Y6MJa0bpvO
YAnLbQQw2UKJJOQRMRSV9hJS0ZzVjuixGYCSZAjajtyY8c3x6tMj39V/I7NKfh01
n9l81bkJKfDpxrHuHlyPkqfmtfRRnquNQYWH0wVERnQ1bp/jrWMqO/9exIAS+9l4
qeKt/f+W/qm3DcScZi/hecbNpbR7MdJWo3iUYvxk8tjj8ws2eELEsWvj/dXb+0+W
3OPSM78xbdib3gnBnWWIOLaMAglTdCVbNtwgpQMt8JmUe9bxtjRX6cGcYCb2YK0E
ehQhRIXCGBDZruBgLHzf+7l3e4AqqPgP9nCNDTLRYZWX8GZa0duy5yRRSxHJq/0g
KP7X29RG6sUCkcl8SZUvksyYt5E7nRE5uelJ/F5m44qZosbiQjGhRwSdEwUITkDm
/yuHJRuGgIfcb09YGmvY2pdADq1BXIilncR/ornnRju1pkf/oXQ0rv39uKoTsj3z
0mxqS2gIQH6ojo4/gxFkb1G2mf/gEuRPvpooLyg4P1U6/ExIShveGoxNDurTTPbI
MXDR46/mz6EYjvO2ERT7glyfuBIK65S9ymmfoVQor34Lro6a/BepYIyjhcqGDiKy
YQ8JOkFsRrqADuWboL9R4B5velIELAzv/9kDN4B3caz3t1C8MX/q8ArGHhQuXFWZ
0LedXvrlSpuRQ65N5kpkyCi8BALGS5pBS2CkmtEqgUaF5B52aZ79utSBQ6OJtZgl
tvoSTVXFDDL07LqZB1n3sKzICdMqFcWjGu24ux+TPZta8yudRmHuMvZRcLTeRE+4
IaIvx+x1N94wbvKQ4kvMCvlRznsFn7/2dvGxkPE/Dte8KId6TUe6gOI5Nx1K8oDD
5AFyJAfYFNdAdoMX1o4OzzyfEuDWjSqGEwt9FmnXdOZz3sGKfnlblU+fPW6QRrYa
VvtFhSUM0z9/UY0QJAawhsO72U67cKEJ+5XIyVDkJThyJGhUeuAnZNoKfdGSjVc8
SgofEU46/9kQFUePLUumihLzq+wQtRQoh0uTh6RADIiBj1raDvUUaum0Dq5aDlsC
LBNnt3P3W3DyKQxH6PztaG9D/cX3hPYGVbgaKeu4VG213aBKoooWqUzzRr3kMBVW
qpk2JCUogprkoKtoyj6M/Tf/7lxhVkyc990ZXRgOhqwHQBADs3LiJC9bbufTkCQ4
Z55T0mhNdqrUY60mWd0GxaUpqoipPif6RXf7oKFC5Bh1erS6i0PvQA8SPh+FM1b1
00ZNvVc/fIUyFpSSLNSbux6oRlrwQjkxPG+skYjkEb5VPiqD44EK/D0yp+laaLZq
jMTe59Ijrs2Tfv+rQE8nofcx/QjtZsY2UDgzK1Biv1fNAzMjZmd1QFMRgW2WJF51
+bs0seotkpbTZSWmlmEWQYxY8NTOi7nEV0bEdz+K7u6mhOiz13/xwrmnUkLo4a0y
9SY9LFiYAHZVt+9RUlBCMXsLtcDmqU+co3PdVBadM5ggnuBgKBBkG3C9qqP42a9D
u5kG+0CoCQCQl5qOfTUM2O2GbrWkNWjmeZp9KD8oHCnbJJTkwjB2keew9fdKlG20
Tg50DXIfjIzr7W/b6cn+kID1f+CflXFDG8wGZ44nZdQhuUBRT9VUdEfLO2JkPGzm
vRP7bsAuF9vwGXCmM4iH62Ibki/BjDGCyOlVCdRFlD2tJd2daKIj/pTSLFZKFlAY
syH6rTK32ZUNr+ImPnvpLNzDElknKbA3/lf4Egkisg61b3adtsBy24ql6nV7BZhr
8Mv+PYQ48MZ716SMD1a7lYGBNNCn/mHHP0jLApk0EuOe3VqOeISlx4kWLVYLr17z
5gS7NVrp8VmrYZnkQbQ3QMTT5B8oPEupl2ZXwYCvcG7HenTCXvSlZUZn9wXMz/zo
Cof+TUcVKRGtW748OMVpfsshkAFl7rspaFZX+7u7G1/8yyCPN4J48GUq2memGAKc
nxuVXFp58BK+FT7mAggJouARxAgkYveiwsXnI4VwOlYniOhww6qorO+7GVJBqdoE
CApKNpAn0w5HoUejRyb/XmTpJc17OGVE+u5957OPny5YkGrmLY6PiDubFe+hDJAF
TA8RYqXQRzjsdSjR5nbjqe4sSYmzP8SvZzjnWvSl0OsjgiZpBGvb/8JuehxSzEUO
pUb1YReSPQ79wDV/5OJgMn/X1UxTbvl0Z62j0kM44uKVWNYJZv6GLoPo6FSyT0+I
CwbmT7Zy/xp6CK7g7u/73a/9nQkIox1BkXojdldhelqLbqZisQhqgZxyxK/gczBQ
TM8mCNuqK5vhh0SN/FSLrW3i8HshSPsEPHQffIlVjRh26O+c4mWHJjtNe+SGVPDD
ghw4IXsfbI/MhG0QDygcOs87mKQKe5NwUo5hr45b1HsyCuzS9xA8GpRsgUL1X6m4
fNiSLpk0L9CV9mpCbV9+OXX/QQaKHxf3rSAmAWWtaHdalXqQpYViHLTjL7U4b+We
LxaDTIRUN1TP7v4UkjN/i6N+sspDLCsNSD2CmUBSLRBsjsI2YNHFctzOUkfHSl4Z
/Xr9Ru4t0vsaZTW6yWmklp6jwUMuyAqRaYDbtvZToNES/VpRhtFkTP3GezW8ynJF
q1b5U7gDUUYnErmVeO5ZB5kAM2ZX885tXuFIiWURdJiih6Qn9RMCAPBdJHi/T31I
6iA73sFJBNCK29EK1dVqr4ulp1jv5xM7I9f6EP2/QOfJKtM6yn8v/y65ZIUcOLt4
PkIbet37V2nBk+Tp3iihlomoNsqbEqr/3+/ivfYu/b5nWhF80ViPYOcoAOvMJtWs
F1lGw6sQM42eZY/nYfXYOtwM6wR2+iD4TGEo0vckl7sMGIP78V422e6Mx9SYrKIt
jgaF9Ax9C5Whha2CBKCh4tFRtDVuxl2b4a6VfUbmv82nalkbnkTst3gj8Vghc/uM
wfElzGL6yZ1eTcRF8LLpQAwN+2r7iscDjc1OVxZYh2EOtpQtARibPv68zuoO22q4
kqMoPRbrmqS+Ld78So6GWPyuwS2Eb/g3XFqgrPF3b+SYwXvX/AE1/I9HPhUEIGWA
OffT1EY+wEVX6N89TVHGvQqEWV2HnklBm/DRCt/LQHNKcwBa20W8XiEaMUT4pNHh
190PRMHFKyCnZg40v2K4Ems8rDaXQWJUKSlmmsphXYQpDAb8xeJxRhnv+1oQ099V
PnV+XJpkrKbWclw+WQNSLASP4rYK3gQlLYyKCumI+f0KuSu6wxgrqUBCy/tY9ax4
l3MvEzf+Ui7KU60/PMBXKAP5QvImTytArsmtXsH0et9w6dKu8DXZ/v30hYi7/ulO
NxXnggJ7QSe87R5POysw2E/frWhS2tlXrnsj//Ou89YsW2RO7od7j1JFZT/oa6oM
16r2F1AL8jocbPHtbhC3rjmUYFMwiDi6BwguFWZYvVJoYEql1jbqm7agpiPWju1b
RW1/lkAUOhqM43Y9YcgYOs+z1KV8CEV1miJL/YWPUw2Ksk6FBBttV39LI3FBhh7W
ihBUArIemR2NFyfSTYfvvYkgmb/931IpPzEYaUVpp3OrxqlFFfEyLT1PxcC0DzbU
cWBBu2J5uUBWgcB0nvw4M48BqZV8dp7XQyLbquYUHKY4LOIlInit+HJXrMigfuQW
yMEPtWQ8pxk41tlMO8LfoYMuN95IEZTYVZNbv8KMhFMOc9PKSdaqeKmYJQ+rnjlK
3TaZQsiorGfRz2SvIPrKx/0M427o07g9cIGkpY3bRx9PTtHhRiGskXgVHcuB6LHE
/bw1yFv8oKNJx/MtqLHrABlUzXkCKVTW9ZY1cqUFuhoPlIrrcHArBj5OFSXGosX6
3u7xMxEwfo94hybvTgpt7+vePvspMv3xCwGK5DqmOZWwJUxml2TE87zVCHaQvfR8
IYaC+w4KlHJSa7HEfhgJcysiARNBOCNVuw/w+1dMwnv92RMF3dW4rKTgzTnBbCYm
uqMaCgocAcQAKZIfJt4tnaPnAh94+EWi3Yq4tk4dawLfOUehJialcb2CX9CNzaxT
x9Zw3A2s51YLi9CGsMNasomnJeIShsfiywCpKGpPfIdtknvBV5zGoZkNf0mB/1vQ
d0YA7Y5w8W6JDMLws4kwWwJrH19HWNGuRhE6+xKsCMUR5nqWjQkNjJVACQUbO7JG
C2I5ihl4QX/CKKvrjOicT0d34zZrvcMOJeCpPO7KhYqchLeWvZMUyWdhL5gpkH+G
ARPEatMrakjmpaIBhxBrsDYjRNVxqWS1ayFfDI54uO+dMwnW8sRoqbSKepY0Euxm
URf/h4AidkHdIgoh6+q6OQjF610NRVwTAL8C+XZZO6fJpPsfS3ZaVVPp51BM4UKx
39A9L4MLwsvsACEXnNxJ8aIt1owjmUJT6caDsxPX8HBEDZ0J/0ireQD2VMURUOUH
dRHX/yFmEuWf2Mqz+f8Dq/GaalL34+JMygRdsDSmwGAiQJ2mBplemJKO56T+dWuQ
rymMBysjjvqBAOd0R8E9h07PjZLspv463WJGPXSt4LoKv5+9cAORFUQLz1TnIB75
AQnjxDUuzDpOC++1MHU9u2lfhmt4Pf42A3prLZScO0zGioycyU0jNHWR4cKVypKh
9MNZeNIDDWrrRWfX5Rz0JfEaYukgu25oh3vq9VgUGAkc+BCQgh1L9LksEdcC2cfT
t0b5xYBZry/6A8DkiO0sPw0aCRg7cWZShy7+cMKiETKoUkFKlSK5fWsMy0q1Bgs+
LHTRLMokRHoj1ZuLvPkDiGzeBUQ2T5Tfk89QamTJjbbm4CgvBGhoi363HN7yrvp8
XdEB/RyzW9yXLJEZpjPW/f1szJiPp6CZxwZzrwLDkc4QKGMDYPYqi3QHYmv9e3Ar
ysjy4Jd/P/Mw/wwxzaWD/2KTdYwGrVLDWXcFbuALqSeR+cwIoFi20kB0EDAoIKWM
Hd0CDYIdNS7X3hkToNK0E9ba+66uDCwEVuL15xcvlaCB75QuyilquHG0MMwef0T8
vMm8oG3skj/ngdxl8ohULiTWc/Znu8v/25AGnNHMDHO69dhB8PGFMcmVBj8mpSlT
30+duh0IJWEiWt01Rgnlf+CpBSVUvo8SU7hTr7IcAHxnDmrweoMJBZ1j7zdbmXTl
Qw8apL3INMQYkJUz4IjXuM3bHqcXbZkc/StG+tT3T0sdi9ShSU8lJM/+PRCT8LmH
RSdMryv4yrqPE3WTl/iKXFl8AjOOBjZC15ckpR5/93X8BtI8QPuElw/CPpudjtMU
YvcUZkysJRKSyiRNPP7mlFvLtWiOYHg/UC4WL2zi7J8mOx4Q+gIeZiYwHyBj1DPs
yAVhihd8LdD2mLvZUfVNiO2SXhE4dJRxDY99SOhhw+IPASgraCcIXJPstmdUk6Wj
xC19vPfuoZj23GTfzol14FaGmSMJYDYqYoYnWMjBW2amLjnHYzJQuySR8v+Pa7YK
JdYilXb2s7VGa0Sh/aHq0tXck1ADtckHBbqXS/F0rNcxOGlmMBOB7g1jR3YvA52Y
czvwQEM627D1RnVaE3f0mxtzzexmbaoS076uFNnhiGHpzCsyeJJlZKE+hsSKu13k
7f+aSlPdKQGRK94xgarOFVaiqaLlYDVlP837dyZwjkLFVOJRjy+sXNNaX/J+5zpJ
2rbjscsQUt7mncOWdE/2tLRaJy9f+r68uTAri1RMXFahqQIqEj+7sPK62pH8WsC8
knwlcQkxnlrw7RTOAxM0xMeml8pF3SR1tBH9qXqJ/vqN+nZIsUGkKzh+w6vywdlP
GlACCnMgznxZjh8iTdFDYJeVy73JRBj64/+s/FgtfNcNbdRUOaiC848JStF7hXHn
5s9EcypOK8KO1sp+jEUgwEEztwx5s1Odx9LcK1MNYHduf4FA+gC/cwuWzheAZONv
vnFsHoVAPWNpHLhmS7YCoXo0vEsYqJUND7XNLls594rCw3uNvd/eqJJZyv9IiDmQ
jjGasDA1YpqCddvk5cIBaRj2Lu3iP+qKkjD6A2np8OO2xE5pc6QpjWRr/Q/gAa5i
bHLTSza6ruZOfCNyOQnqEt3I++TrJ3xbB4n0zP/MPtD5tv3lyPHoXJ/Fz4fMC0QA
jjm2/daOnItTnDFRibhlHxQnrwnQSknN6iXdD2Ykj4b/OjUTKBEaQasGMoo5hR/7
T6cXRTR/GzRjdDjeghT5LXTihFOsVDsGGjue5ZDgqjplYMmULfGPnUcPIP1Vbflz
QOOKWIVt02NdEqSQH8sp+YeMecMFgqY+r+1/7t6Dt3m7JwfErtBzMFAOCoC8k8h0
O1VtKT7l/B9kd0OUB9XnpfIxbfhM4gSbeyl3rV3JF3NTcYdf+5lo5XYmIO79Bny4
3tUz9wpo0m57bxvt9ywx+uWkTTOpuIwHtDjpbBE4ldkSZ+pwFfXmkDV6kBXuSCWO
ipR+ZFCOYcYwfwWz6OcvE0m2ivO1azhUKS05rR1tdu/rqovf/Td+Ks1DlvChOiqH
B0siqQGewUxC8zAa9XLn8KeepSD160RPLhkwZViKUyHqtqu3cCDfa4y9jV3Oil4h
iNKKU1pewAILvli8uHBbnKxHQXBvMmqKgSLUsFjVpnqTjnQmrHLTv4fcRIV73Bi8
Y73eLPgQ7ajqmcK8U7NM2wjpGEhH+13xI5v1a9zgIgbYsJYRs2mJHh87nZTW7szh
h8ZWRczjPIMiBdWo7u1u0uBS1WC8ZXz6hGTFklTv3wDPsgO60CRVhKo7SIRRBfjX
RGyabM/FqzKQB6JZ4ndK+eDWZi13TZ8fwSXRC0b+d+N8BtKx69zCovLrL7SCmTUf
g72phWxUZq4HsOMhf0mMuKgP2MvWlxnkxPBxk8QQLbCswxFVESqmw4wzzTO9ndF6
03z85svsTRp0HCrb7QXAOAMrtLDxFK97lmVxfilZCvgn1eEZcGd114vNhTVuEb/k
LG5fwhM8co2yicwTEoDfrBCsdDYaZmtcPza3bMmlA+biWB/ZJzCTwEVN1bqIz7ge
fZpLPlw5hdsr45XrcQccSIqan2/Cn4jiaGSBybwuVFDia1tqHPFhdLmpd7AcMFwD
/kHQeV2dh0aa2Z0tPPi8eYWGPco+yrlae1ZX9PqI7fvQvjiM1suU5bWPJOSsvowJ
ZrLTmQ8m2kW+47zZw52S8RvadjlaEs17hdrpORSg+ATFtB1O9QMX6WdC/0WfcQ9W
zoF9YZQT+Cv+U+YcbZ6RECApOuEAwpleMKjjcKxBhNQod37UrRsu2kn4bgFOEgcn
cmvu3TGSWCoXZL7dQY9R4XT8SoGgy9EYeVQnskeEMEAKkh8MZWoad0DhT05rxJXf
DzVLatQ6H4k92T0mBwSJ/UMe0aLCTFwtYuQE+KOmGJH/0t37fYmpcckI/EfCxO37
bP3hxnRNXkilYfZ2L8Xza5b3d6Jpu3jIb+pgO2jzoA8KhxMgBYxUWiQkkszZYGEs
cW82nJNBrrQvhgkMJ/Ex0v5J9LXyC5dFMJ8wunjGe6bhetZDTL4+3MvXvudS5KjJ
kN01JmeaGwPcYsVg2pATDaxPAQg94LoKHN62kiYTRV3HuhpIV0j37fXqGi+yTenx
ONmW77NzaLcedsqahd0ukduaXmKScwkIDkhynvehMaKYrOa/4YlF9cWYCVq2MuaA
gpEOt6souoZkSN3J4xta9w==
`protect END_PROTECTED
