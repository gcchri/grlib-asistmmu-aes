`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5NjX4odZSDN6eD3ufb3WAbUuj5GBjLQ1XPfqyhZ5lOMwdXJkeh/wlIX7dzMJENzg
LbXDJHSp2ntGB92hQ/dOz9roAOJf+v2d7ixrlkYRAMIFLGKeP4jL5NHtvawJ/yRL
WepNV96nsDt2ArwA3CTEkEqUSOLZCHe3GZmvd2ma0UJ18JjQQYYCRcjsPT8fPHJG
quiRVShQDa5N829/X342jnoP2LH5ehdSfwAvrmeuePkYv98NXmG5q4SAHKyOapr7
VaJUClU0Oax9QquX3Et/i0DulNYDm76cqO6iZIqrdaRNut+01hfdL53IX9iZx/j3
htjxn+oQVOfrnri8bkONZ4SV8T1JMDY5HYLHl+z1HKoHSE0d6UvVkjqKVEIaoRAM
l3MlGc1fQDnWEutAthWf9wKNR2TuzCutfoe/08CkHQt+WZKdFuaNVtWF07/YK9/E
p5RD3Wx1NuzWCHJEA9gSIEt3WoGchLk0JTGxK+pM00Hp1iVZPgZQOwe6mQ/Td91g
GtZUGIiPpc6+CWlp7CZcqdIs07lHYqvbT/5pvXRdtlgLkQr2ip6FBN148dgwH/aj
DYGIlLT72ApiKTaKTV5iI5mUMnTcwWwhPTvTbuHiMk0bPurdeO0QOhHZ9ctU7lLY
PQkOnnwQvx7JFvKUQZDC0jN+/LzZYlPuIzJO05rUSrSAiIPFTRJK4IJVQSLKyCkq
WmiFqG8NZDCOEFOeCjkMJrkKZVf+JbXNlDbdtT7a0EZz1A+hrsU2ycFhnpeWhVJ+
BIHqv5X1azwReT13K/n0KAs6YdTQhOFmpZ8DHhmdSYcO7qST/tpEc+cV2EFX+uCv
OuzTtO70x6CBKXSRUJFUw7v/APTuVMKPe3DXiNDxJTz2MLtyW5dZMY6wS+g5R1Dj
v5PQFW3ragmbgzT48Cyb65zf12vKamrOhDqCPe+1ocJUFEF52hyFW+ZF+tknK8S3
`protect END_PROTECTED
