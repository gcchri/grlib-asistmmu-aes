`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64vfVDWZg1NZaoEQlobqo5uPOj8nvOOTlu6ai7e6m5SRcXSaiBqHp2o4O6jGIpgF
4Y5+rfPgrDUKac1Ri9d211wCJw8sT6ruxBrq9VgRC6baxVZIwwQMgUsUAedgM0is
74JIH3i1NAjFSYJM/so0/rmeWnIimzRnzjxwWVxOQhqB6eSsrcjgNcVcOosIBqtO
OCaIMCeEsKMHP+9JqSVSLZdWn/DqDf7SzOvbi0KNNw8EPBmc/6oswYdeBMRExlje
GldMfSxCu7+rAcQb//OIGgkGB0hQ/qpAbdK2vVKiiY3GUNVFxpLESUeMkkkVGAPq
mSno4dL+ELRyNe8FngQpJhHaXYtMhKHVJn6GvUCSHPIKoBels+KplQE0ZNqG0zT1
F3eLWRkRnWLKhJ2kpBY5WJ16hNZGHlce8RrGbfO2xYGn7G9dU3jn5DI9QEa1J13J
Y6S9c8MuuKEUQ+Nk8oj88OwxMJdjEi8MzGN3nkazG+WS9VGik4HkfY3JXBHWYbHb
ESkoCDjyRp2/mnRnn2IB2zi4gzkdjPtsMScDl34UxUV/Vn9v8UgXpxfXMsi0nvnN
GUxtfzjdvEGHkS4ucfdZOl0K57SnHMXLKwOtzkSGAoEzHFG34DAlwryE3T6aZ4KR
Lr8L7mmX3BaN1LF1QHhXGlyBBrXgpI+PL8HUm+jqsAmJwGuEn7BefJ0uC7A718pQ
ye5hiM4SZeFXN+IfXNB13lDxQUzup8DJmHUajJSaMu61fbMou/F/ez/WYwurpZlp
`protect END_PROTECTED
