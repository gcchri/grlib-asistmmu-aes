`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CUCutX1Lwy3BGAAPo3xfrnL+qxMIhVk9BTD+wjgj1Vz/TV/0QFevTxB5h9w0OBGd
lLiqO9DWWGHPkIoNJb7pWeW6XQMgp0y8FnZGqQWiZORL9PA3mkVTEqFw/lkKXkP4
zqzWDsitSxAbT5j+fKdo9l/B7yERbKe3wNf77V7Ku5vmteeLDfLvR6/USljKnh8T
jdTjmy/Brs5He5PyxNum+HWeNY51PjDrTRMGJCdAuc+jny/K8zWQGy6H8IPeELSu
N9s8/HlZRlHn86cBEKZ9l1yackj2DIWO/jr1Q2Zbtol8DcWDtnLJEktcoqrQYRx+
YIzmL+W81bKGALYrgMS7fM4iWlqntwGkvgPNOCaKP56IBk63H798fnFVqgla3Qmw
PJ1pz98YWJX2Kz58oaD2nzhLqr0htb5h/Vb9exEAO3RKPNGJavlEYIziZp4on6CZ
R2Z1sQNB4MZopRVX7PPDkjYvlxJj0EJo8lIsqs2d4T45d9SUtd66eM4sMTGXFM3F
MQdXUTfgXG1NMnmQ96mfyC6wKi2t8IpcFwKAnIW7K4mVD7m1gS91R2Y1xdGRMrHd
ziF4cvkjMidDtbiqLaLjYS8namNxCY95gdbSHRFd4teLumS/+2HK3NPBAHsg0TYI
J0QbXxBWDAXQUdZAS7H2q4tHVHl1Hdz2qtjnSKxi8TBdfSDfrUKBpM1qS2dIXT5q
Skayeblr9n38Ln5xQxGmYaMi4IvJuP1tkCdDJbOw6m3CyaltpHbM+ktysG3yNEMD
ILAN33HwiHCD45fsjgRknwZyjaROzOGxBZeRvbuYGy9hk5d+jq4FX8zl4QAWYml3
28nJuVPoKpgncPZCcWvPo+PyDqbLHPJtNu3O7x7vVu3WnBV4XiTj5+RHzSnAiVPE
oropRlwqVhmvrgBQrXvQy1cJ250F2NRfkcQhRKN5SOM7tyiiifbuPtKF9uwNZpaA
FWCRI2Somtxfz1pLViKqWa6tM878jkStcB6NqnB4FfHDt0iMeF2F6L6O0BSHFiQ4
6l82ClrMO1qi0G44AMuOp2/B88plZInXmWZQo0Y6hoKVg6cclsoe5m1bZfdoOXhF
Pv04IrNs18wkshwxN9s/dWNq93Eg1tdvqdk+NvkEFKJ6OuuYulX4M5/OfbEBElmj
M//G22Mw2wyHnKGX35u3gznDckG98S+Jw078Ab8eO8ClehAyZETjdJyZzbOPO0Wq
97lWXqDwjYoPJRP0tyQmONBJkYq7mBY4F7jJD+JPJ/OEWWMDk4oud37ga2z0Jv1u
dlUmSSuW6U13dmbUzXHOAbtY4HEFG5SOsFU85sYduv7J3zdOGyyfHv+DvLaCdU7c
I6/s6791BwdOPKbWXw/pOK/KgqRXMDPzIZwIcP6ePYlIfvXitEwRvxYTKBzjawNe
JJC8XsWuYb1VtipZxZJJR8n/vQVmyXi6QK7gEMtfK39hmiKwQqPBg0yOBz0utuZl
3345PqENrwZ0pTdSzXCwToyVgmJ+CHu61Ts4YE+0F3Rn4JSZfIFS9Zr6tK06k1eh
QTsA0jHZhHRmCFzAtLKohXqKVsgQ1coDjAnShCg55FLCZHHjckKw+Z+F6E2a6k/T
+pzeiDalPmYXrpn/0cNKAhje0ShITXZp/HwmrIEvH8LcN6OzhN7xZobCpSj5CGvd
MTbsUrDtySP/wB8u1MkjO9kk35IgNFphHrkdCxuBHA9z3oNTHfR3xpyo59hRZiwa
033bI8CB/Z0nCisA9eMUq82V/1TWN+eKi+57bfvzYw0ULGszq0suz7zcFbjKU4JM
jhfhMfCYxmGpeeExNvoFBYhwtyhOSFvOAfRtSRtJiOr0RB8/ksO1Ic4cWNV8v1DV
7wsVt98i6BAm+hLe1mOlMv36lxox163/2SzLE8+Xzi7J+GTh8o4emcov8HjVngaZ
`protect END_PROTECTED
