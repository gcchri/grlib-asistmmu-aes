`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5a5a4JCrVcnOt72HMDSGCTTErzYptkUqQoZiQsaJRz8u7+rlBNP69xMlwMVWsU6U
tfSOUaTVPh8VFHQuNqIGbPXpRl1AP1uziMrSMSr6tEdJOQu2b6TTMffXkI3OHGT5
LrwSe74Jr9JReUAtXiW30DsOCaMS+9AfId2lGXmQiRKMWCDm2v+qVIny4qUiQbBP
6Hcbv5xcfKBG5YL7dP/h2aLsh4+XH3MfTxOs+fa3enhFSQFR60HuzQvJHxO1GfgY
n1DyJbD1tyzqQ7aOl3kJapmsVequlk55viakixuJJVe3VLwca6nLG5AC4qpw/8Fa
NZouJDWUdllJp0esH1GKYHNxuCuinlOlSsYSHAuy36K5k9Y+S0DzTHsfeJRn6wjG
IH+brRgi+qzHtgG/66SJyJDdkhjbOiJeeiMIQb2HH38X/ObUm3gORlH0jscfjtZw
8f7Gr+/l+sYSaJF37BAaxVAvM4BW+GQJKJmTh6XhHi0W9iej4jvIthcHlNb+Zw1X
lPbxxMaXMHgLCdoo3uwhKUpiEfcC450CoiJa8J0cIArHsX7ZTOr7+nbPQgxSDRZx
yUwHtOjWfsPdgDuWE5tXPxyrxQPtHF1BrJ8lvNopl48BWQKYIZw1doc/MvAYQ0Pj
gkqIw8vgscZtF0Myt+vCgVRp557IiaD199NQGJ74WTHfRCg7LCgxV6aV0iP/mdFZ
fKmQAo9HhMGFgAbepZ7kHwGuO/Kq/7itQ6/blJeBgpSoT8zduNcJDREvjRSFONCy
xA8tajxL8nfDAj7Y4Vt2sAB7IbDs4sXveXztvW6dtZ7JKyyHh6o8X3/B3odKM0wS
D+cYRahy1KqT1gt7ypJ+1T5PqLZnZCmIeB3li+70ISyxmOBALCFexuoDoQiFE7SM
qMwwkVfiaMfgpKPLqqQFUEuMwWBreFUrYOL8IK8YKNjZTfZ6GtnfqZ++0LrUVkJb
BKtq7plfUuf68qMobxy72ip4G9krSilIG6mRfC7P3Kz9yIR12kWnKVtjZJIT3kFx
YEZxUlnJCz7wR4D2leTwGA==
`protect END_PROTECTED
