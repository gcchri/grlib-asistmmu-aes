`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KdRttjpw8cuDsZMPuDTljWXxt7KPpvyJmAMrfYPyYlTPLxzq41jyGL3C1BiyhzAg
BJOg9Ri5D42YYd4opMPBIIH/mPg6/w5bjVwG1/ebyiUxnrhTDEBPiQ8vsgmWdB6I
L9cLEGzs8v5FBhKb5FLD4ngKI3J2KhZ9ishubHjFsI38KwECpSZLSdi4OXdhfOPp
WmhIpIPEyagrapAAB9Loc/VHKuQ2tbypoePZNGP93bVpRTk4fzn5YfFL0mD68tYa
nfp6LB+w9zeCBXAyKlscL5jlnNctYM02s4qIW7/dgj3aFZT/pgOvj7NQwCjI3D/X
+9WjDO1RAH2kjc1wz3xaMaXg8qFsRaBcQiB9ebQmM4GkIAU1eqoxrHwsxFJyF7to
7lCgUU3eg7xcBVre+xc8MDxhIy09y47bqy+AWTZFvCvzq5rWw7bwkchC9CiKrPtG
0I3UiSGwp8DNG3KOZFum1x7S5VWxInsgtnTdnoofWLer27CH9RvymmPf2vX8fK1f
kw0F01tNkyHqHheZ558zfsynxQWwIhCcA0GEn9KyBnZdZb6Yo2+BIqmRU4bGDYeT
z3vzUlADsNY2+wi5pFkG4z2OBLKlL9MqwkICXqF6jh18/Ak6Nr7ulUcCqNs8QzkD
5x+umYZB+F8GdElinfay1zFvySk0z+1ibaFuMjcE1EQn2YSZYwbBUoEihkEOikEY
U8d4wXBAxeNVxvM7uMXwEPiXzOo9IGrfU4M0wkSXGTXVm7YsokW/oL9v4ikN00vJ
VdLhoh2k9YErSRPBqTECc/vIG1LAMn/4NGkNo1mlUbw0zNuxFnoOrYfbatJpXsYa
uZz+wjCaNhmSjnZvBSXB8A==
`protect END_PROTECTED
