`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6oPchwLvCjIU95/wUTMmZmum6ek7Dy0rTlkdxpUhJJ+kAUG+E4LX9+Mohjn+Hlzr
k+O7unz2xtfmrrt5i3TXjCyGmFhjKOL94+EkuzPicWJAWxev1/acIVdEJgBdsWqD
8mwfaLbSxfE92XsSR+vsyfdySEiN2dJPSYPqO1Q25lopMPISePNrwIRt2X541mwX
snu1fHXUwnI6QXOPqb1J37yTusaaQmGjJ32AkeZMO/+cH2klz+0s9BE88YAqP+/Z
uNpeEKQ9qFZXMHfl9eldWI4LF6oSoJiooWbhEyrgAT+D1NSBqTHwwarynfg3kGiv
YtQa+3oZmAbMh375XTriBbgUWpuPUW7trHB0tLl6Xe9aDpR6HgALzFqtD07Jt3FB
Bc93ibRVNE6K5XgQPUYKFA==
`protect END_PROTECTED
