`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eYtgTDznKS+syhJxQk64gx2k7RIIj4E6fTpa6mb/PVpL3ZWwx77qwzfBq/+lvIX0
pItMIQkWVOvtgJL/qsnUDhXar8bM5+kBiTjQJq9BI9mmXN97Iwk4jHYwQlk25eqD
10KdHYkcYKcsqaL1jlR1AWFhr2Zo0SSr7jEE0qk8KG3aZSps1/ZQGWNwLp0YrE8L
trMNvLiRpIqs6hH5PhoUzgJj0Q0+s+OD1keFqRkuTq84unO0clt9TKrIIL7CWdHH
F+ps05YQqsDGnJNoPX/wMjHLnfDXEH3ynS2Fe/oEFpxMW11HR0mimQBhyOtlzGOX
K+zToI95fbG+sFFVTeTidkdH5025y4RHQB9ubryWyhwVl2K8/EjPon9PvdkgoUVU
9YiqXp2C0o0ktue1DF84NI3dycW0nt9ryW6rTDkDxYKDkgK7lbB4acWutf/q9vH3
wapWFkPBojVyikeLxOF6Bt9ScE1ylE8xdQEKO5eNqsPOIo/3UzR41FF1fPgSXKKi
pX+Y8Wsrfvi0zcZAaQLNi/yiVrfsQe95WqPA4ahwECymvlm1HHzzcSgkBwL9sg3l
wbTG6mRAFHvJ84jrAW0Q1QPk3SQjGgJ2xRNekNDMpxMMVknf7RtUPqZrUyRHRmg7
vXq4Ksjq4j9zQmgRHr+BFoagN6Zm5GPFbkzvvVc7Rs5aIJTbdfC/atECphwjuTrb
m3pFj6aApFHvWocgzS1iZQ==
`protect END_PROTECTED
