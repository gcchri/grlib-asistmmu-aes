`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sviDQvJoBBIM5khzFZEkEgaCdHUC+NOD+HuyBz+s9PIPQ5l+xhpuPgyZG/gQyAUT
irnu6cTzdBiEwz9QukWxq8sV4UwfrwCMdGyegWiqQlthZU06wIKPWDdyvV6SwMeP
7BeAHK45etDA4nVxzeNs+HWnErf/mt0qtvzz2KJgDjX34hUtKYl4t1iWivKvrN85
Mh0InwUUAs8n/NcOdm70hc56xq6wUcw4GWxkVQwydd3hhtja9uNKndBoFfmlPm62
ct0Cr+NuAk65mEMHYlqY47Fa9qec5p8IqfBIjQNUfoZKcQNf753PR+dLVDNAyQj6
hgRD5Vjs9EHcVERBCmbvBWttT/1FR7KKHlYTPQWAGRZZ+5SceaWIqevUQ3Z28rKA
d0aZq/dnlJrrmCFN2cd5KKMpUf05NA0D/lwOskBMc4wA7M7vyfmHGUyOQocrnOe1
VEUSH+sTTWES0ooDmktZjtReFBFFWrRyeFMR3JV9l1OM8q8YbrQAiznq7xb5Wo5t
bNfOmCqX2p9E6lmOgNgJF0NhqGSymukrs0ukALtOC2pISkmijhuW3+baTAXdIf80
rUucFhalTSeEqv2GJT0YDmoUX991iiXIKa4dEE+2fbYtO0tDtfWrpf6JjbIFhL4H
FWYxD0sUM20gqQIWZd9A6kf8QW1amQ228hXCs698yZUw3doPbDSZJ4DW/qbP/AaF
TRzXaVbwZ/r+8OaPlnI/B6IQUMYjQ9PbFNeky0Yu2iiF+iLk5cDZFDB+mA6G8t2p
LwqRrh3+dm1NOXsXY7yBDW6OzJhPjx7ckCvSpzfVoiRE8ulMHMXG5pwmfe3wwNnj
bRtvsH87EbfLITGsiitZGHjxlBLDQ75mHGcj9seUgar04ScKGd5h5uY1ajXKMjil
NJgAL/ZlWhIiBH/Y1VWUGXi9KRMV05wRU0a/9SyWdDKvzJ1K9gT2QOhnC8TuT0M8
SJDgflJKCz/qvAGV81AmcHLlQTVqpnnd4MWE/RFfv3L5vCBoadm6RwEFa8Q3UAMY
IkiVrOCWaxLc9kALFeZc4Nqp17IIxlWtS2SyQmV7Pudab3rRk97PyiCqjzoiYZy3
vItwwumbgrS1UH87qsHaRkN08IEhZZoQSqRJfgdoXt6Nz1QLfC3fd99euNJDWGKw
5MT4h+EGH2oOVwXFxWolh1V0JczolX4o7fvpGLyhnz1EYVHCqpX2IeLFGfc8bM26
Z6DK1iXq2ZQWWifnQzX7NFd9XWgRSiaJKVriM6RlQSviXEQSQQUKWq9mInyUd7iP
7qwJdxdLyY+Hw3s0pQDLdZj1vmMzvBAw2BhXZMgolBfwdnFXkB+XisC8ZYq9M3u1
EJn8HC10vGjW2FkSn29VV+A8hDVceyNCOAz11GxQO5r5mZpVBSfrjfDEJ+XcD2WO
ggSDoKd3dAVhKb3U/OivsRgBfulbvOleb0BIA/wuZoYrlMprR4kW++U7HMn8XQAl
UO5gPnXMT5MwyqVSB7d+95xyH8EPjx8TSHvbrOf4Xnc=
`protect END_PROTECTED
