`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Rk88uSQhnls7HVZVHo+8DEe6wZ5fzE+wrxSXcCJ6nS0pDPYhU67VzPko9SD3O6x
+CmgJ68jV82FVBdrseTiUB0X2m1l8fduhVGlrRyw78HXVcyUIv5z7JQh3QpMlX02
Y96Mqrpwbing6al0l9deDJRgIsJhF0OiPJMEVMSjGFfD7jApo4yXzw3TJnexbP/N
n3zbkLipPymgT1SypwKs1pRoN7b2qTAYJ4PSu1V3qqup0iwRz2wU7OqJ01Ux+nC1
jvT/6aZnlYXh6YtkduBAHZxm1bFvr/4hhcCYG4FZ52ksy0iE17xoMoU4e/EbUAiL
MP7mWiAZEeTxZB8rLTAWTsKhrHwQjfuykxbIPjRvzZi5s/c4XGVQpDfykx3e7BTL
UM3tNOj/znOkP3i40/KKAARGlmRI56HpJKTVBC4y04S5AWJ9z/jZtKRQynnwQS1D
NmMBmj6LESpbRpkvV/y9Ee513DlSOBMtsFGKExS/Gxp788QY5kHRIfocAPljkQew
YycYxOX69r4dNcch+asv6wnQ2ZWY/NoJMI5Ufzu5k3xnCyGhBdqJg+GRywmYtHZp
mnpD+JcyuvbnGn6Ly773qNwLf/48R2oZYEKbPQWmICo=
`protect END_PROTECTED
