`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ft2GdV1XvFERRZqkSyEJ2wqM6nOKot6dEfEn49sj0B6C+6o/2zrwKnqKuSERvPsN
J2Yv29EGN8DuQXDfawbBZJua5Nl/d5T0ku/uTqjqEr4kMuRCrUaQrH5LPnvg594q
snLrJNI4yin40JkLHopz6guczkmDZSWhqqt5jDfNs4pMBkyLxmkmcCs79fDcMadZ
E1pB+qPmHGy4wkqx9xsZsfTiSU2yAM5QcrwRHtZxAfhB1/L37fYF/mvWtjg5oxKK
pPtc2lkkSLBAUAKfvIpjqNWJYU5vyqrMdRJ0LielvZWRUhykTpiWtagmYEGHnoKM
iDDymlL8iHnlS7DRQlVDqTDzSsQcy2yfnLs8SB6ef9/8g4D5idenIWkgReQaoyPQ
+MMUrK8h87+/sBtLrdshZ4ucXrlV/kyU5IqkhQ9BmM4xkC0CZBrsM/gQ55fx1RkA
udzGdq+bRCUsiaYWhUox+BkY2lctcuFzQWut0n4DaGS14zMlNe9NWVUuHOf0pQ68
YbUp8/nXBPl2DrLiqR4JjGnp2udiHs3/5GOfvke0xXW8eN3QMyK8nBr2w6O1Gz+Q
LA4j+aeMibt2YSV6L8R3JY3KQBJGxQllDDMJzccNeEU=
`protect END_PROTECTED
