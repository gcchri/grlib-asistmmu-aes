`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ax9yefJLhfbfcL85dh82fI9lvsDEnJF2yjvV2yNZi29cVJK1HtVWHHOJ9RrpeCS7
OxlSvnuVSvfrv0YIJc14tbPeqXNZSiE1haYKDZT9Is/hwHAaNhHaKOU6RdvihMVx
tfLC6tNAszDLuPF6ylYyxyktvVNlSHU1dhI8PnjKVkvnSUuco9CgN3QseqbcXF6r
Jvu6ATPu0bY1RjdKmDcIi1px1cJSB/VJdi0Tk8Lymet8taApif2SMY8clttv53QC
C2hofgxySrkjV371rXNEK+6djMu24nUoxvzQP9ZNLD7ac7d9W1ex38h+cGASj5TS
E9ykVIGoFFAYP98+zR0GGQ==
`protect END_PROTECTED
