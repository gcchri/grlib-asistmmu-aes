`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yR7PWcfVInbwoSa+VBPZFTzYDla5lxnkmkIpfn3ZFMXBYmFql2W/4tInRcI5S+hp
6QPjpzHaKOn4kcy+tiRtj3Cvu5XwqgdvjHvIPABzkz9YC3OdVvQzrktTQe2YETsX
d8HtQHGvuTzDiQYIKNqnbpBaOY+sETG9wRsJhL6Ru60oXs+9+vdYBdvQYUVNUfpD
0H5svX4nB8p4alzT0qC3y6HV3rJufMcV8jQAsp1MfXVxLN1eJThUAETUE1vwtoJU
lf2wRWtQg72NPQGpab++UBPEDGBctTaNi2WhU33hroljN1BuIetAX/A3dHSIYNrw
pSdyq4/hdyoyPaJI/RfzkvVfUmsZUdUF6eT69FPUNSZcvg/1SQ6LsDtXJYAnPyca
dk9Zx8WGN6fUGznhoDJQf0OQ8dxkDtpeq9DA7Av2K07gM2AZuA/zyH4vL3Fg2iPn
ztMpIr4gOeNgL4YvZMDFOQaDlPQS+rhjloW6onye4LqNICBCXMrF78I498aEqVsi
i1CfGgUsoDciZ7tn0CnCJ0ybNk+ZRoZuaKzO+nftgLRniMopU8BDXIM+uzqZzAhd
TGeMJ8kmSMNxJxDWI3FngVzVFjHOTetE1ryJl5ujx530P0i4bFMsCGc1pMFXHi2b
MXvUSjLJC6UQ3AP2yhVZIK6im3DMtZOU4ZqDIOSFx2uTB25LNLI0fqWuxrB1Axfw
voWjgOpf1GTW+Zws00YzzQ==
`protect END_PROTECTED
