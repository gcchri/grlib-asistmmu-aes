`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFbdgey2ICFOXTx+8nH5keMvi69w7AOIN9v+7TofR0JmViCobXiE7/lGC+MP9jY6
C+Uc5oz2jCTaGtz2QOg7fJWLOGwkbrZ1sGjHqD+1LloluglD6AB3a0KBpwY41IT4
UmnVHgNg++bWzb6UkM3NLGVN98tXs6Tci1Da4VkOSXWVgJP/FPz1QEaKd01+SoWj
YSZA3Ue5o+Uxt2F7tAvoNhyBjuCXhdTi4XDiO4weQhZhIKgaMw6fvgLbDKN/yxyz
5XKjzVefPVoRQX1wOKWWzeS5d0aRbPGMDBfo5kdwe6UV6BMEN2CV/hNk+CPgxNKx
tpdvYCOJBCKoXLhAV6inys/+Ra+3MYP0AlgmpdvSF1y3TBJwlt6p/VU+QO/0xaqa
CYRL92Bp8GUuUbRG2KckNz0ZoM41g72bwFfcRjySClIzK/xyqjlHDBh9VqtXYBAe
`protect END_PROTECTED
