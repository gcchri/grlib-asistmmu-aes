`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVQewETQMiBkfuxqeT8/lzUPbqZV9NKvvPDFaMGkyMkH3f/ds1TPnUt0ARvL/JOW
09QY7TQGz5+qVnKeoG1h0nhD+9HH6Zc0Petxpv6IGDWt1TyM8SBnwLcpvrK+SDgB
aDkVW5Bu9QrWxAphPz9Fsa788mtTzQFVGf445fQ9YZ2TPMNKOTwTf82ANe86CO7O
NDQbGXBBFiQGqG/2KOGgCnwNCk3KBzEl2jHN4siM9H5QeCLXNPccn4vx+3sDqUGO
QkItJXBMSjUv4NophRXsz5etr/Dnw4bDH436kqId9Zg=
`protect END_PROTECTED
