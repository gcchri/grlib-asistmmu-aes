`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvAGe9auBxvaEnPmK+BWpftJ/thK8BvGOVczsVkV27QM1RTbNTWEG6arExAWNmTN
VvHoX0w6fkVKEjztWDiIL5+ALd/CR2DfqnlEZ/fAF8vUky4z1V0RGofuUAueBL4T
Mv04KH3eoWSaCK6pOC4kSiTjm5n+beOGCAs9hQO+q9CADDlr3mJHK1kx3zs+bxNm
8v0FK8QeF4L5HVygMko0e9u/z8WQoYwl/eYgfX9aLk64uYXJtonCOmyKuaTqOX8q
LX/ciopjKBy526uZXsLR8xnjLviXdOg/wch6UlvokVw+mqajbJdBVbZCI/ZM2zJ+
alcp3oupRATDaJ19/mP42n3WOxrdvnVCk9u/JIE0GBiEPiMQCvZ/gBLHWi3zmG4A
sMAYcfIezrUi63CJ7gfsHIknHbCplMrFlAO41LmQfv3BpxFo3X7HnHgJjtlJDio6
sj/0O9ZCjDzGl7UuGIeVHvALSSfRLsuWi1rR1TIw+nQg39KkygyvNo/kX4ikY/Eq
D6xtc5iyQ/aZr7MO9fKoJ7OdI0LVSrFcy+fc8PWs6JSwksz7L5bN2eX9YvRW715H
xvDhQE/ifzKMVO+XxDZIavuEjyjOuOGxozMCoZqbaaIIX2x8wuSbVjMjK5pgx4tj
c9h00UFqcbyrPdn7nMjHIPxTAAb09AvEeix3geWFVBYGTi+UMz3iZ9oZpVYIYIsx
kKtwxL8mFLEM1Dua5h/jnWKujweljxXPOOs5tUzKo8KcmsdhnjPKgkRmrNFjly1n
ftvB51ycAHwmUAT4v3mXalysAfV93UNqxDwKIO6wRYZk4moFMmGGMuQbLN9KMIag
QgToczG+jCKC0LskVAp9hnVjHHLBlbXyVZaM86nub7KfAjC6lzjK2eJV09E4G6r7
1ibHHojAYZqCkk4TV9xV27JrCAY4kfLS7xjqSBEfkKWbFED60fne2RFpKA78PMzL
62Ifwvoq4lOkvryqOgJSa+Q15Rfw5ye9kgHYJjRJyDh/SQtElal9KGfmZzqI4wTK
ob854TQ2AKCj9hBeaU2UGEplRW3mfKT3ljkRrEnBuwl0QxW2dFyVDPDsGE8CVcQj
iH6/tuSkGATJyuyxbTePIJfnzKqV72Zv4pe4f9jaSL0DYC2m2TSmUWqkrCIKxbsw
GWkeqzxw/7JiMiKRUGa7ajjJLEzbVSW/94ZqdUyx8skAfkYMICIsVtwVsvxIzHxP
tBqv3iFW+mG/ztZDddU/NBywglyg8yHNL7EJ7Bm5qe56Y0goPzANDuc85D3OOWjY
rTz9t2m4dgC35GbQg6U6mYRBKedtXrgMf51OghkPW6sx1/3ZRFrYLks0vg5LPwIy
INV0ysKVwXdO0JlEBWqhSFHifTNGSjlQdvanCNinZBu68cGgXJ7xX9WJQqUcsAN7
uJbROYDqYfkMD1Hr8N2nTLUYXDC4upTqhcS6nDKYzLcmgfzw+3XYmJ1R9FFKcgeE
qtIKCV3YseZlkKkCNpro2WQA2dzyTvQff8UTM+PQgIYiefambkJ9/GtikazIGSDe
Eq5jG0k1j4qMTJSUgHVwCgjKdU0yBG6249JPf/4ewP7WPlNTlY4cJCkvkmg9g5t/
GkYgOazJJnOSTJWVZosq/FPMEjvtgfKir+jRj/UxrU0Euya+u+p4z5ZWX5Tjw0J4
4nJLLilVBwfzL5k04bdhOd7m2E+HOZxCKXcX3nq78aYQRIAtFoSOtdNWeI7e6P6W
0Lr6FEI/h6O7qzWmddnNo5TV8fTPx9cu8gMtti9w5XKX3fUEQe9nKURqh1wpbGSY
20dnlExAfrxJ5pU32kxIsvcPvllrr7kJQ+4aIMWhpHv6fwE82InfXRLM1kpM6Y1W
GmNY4QvUwI0+HBWs+LE4LFQb9zVUFQyMubENiWnNcgyHs6DWsfPc3SvmRYbYgabt
s274kT1u0b2pBneUMAZRjA9ZLnd5mpvzzrxBYugGws+BZ5hbv3NFaJeemhjd5byR
2f2qxX2ZlZPv77e+77KVuBZY7vSQth5CcP73lHjx3duspPe8d+nk43hBoFz4wJsz
WNay1P0UB5/fCiCDMYdCU7ew16u4y9R+v4Zs8L2eWYBAtBsYuL9My74Z8mDD5z2x
2mEGWDv3YIJZ8f9ZNjtCJUJMtn1U4CdQYR5H2pYVMXwC29fe6mq0VIENlpb5/d2j
7iy9xVifhW2bCaf5iNXEGBzKW6DeekQIq8hyFgVgG9UIQbdXLxEman/8s9BI5BG4
4z8xB2KsTcOP9h2zG8N0PvruNbYHLE16/RuboyNg3S1ZexBLYLtBX3MW4mA43vTF
Bnkfy2CfK0tMi0PYISWUj7RSN9uEp2k5oAK3stpraiPskrmTvue24gPEJAHPHX4J
XxexBYf5tk4AgApODyXHYeKjADT0/Fz0YWgB6fWOn+qzwTEto3H/i8sUUerhlnTc
lUbgHEEcKhBKdOyJcDLQeopFz0yXOoZhfVTgIYOQx5lU7bV0rrYzQnNbPVfyVA2a
cUqB84JFvoOT4RtcKdW0ybEdAxiOQtWLkRJd/WH61e8pvYjTSYbttfJ4+Oxa9Qxm
9VE9mx1g3g/sogmsJK1KroEFouCZQworkNPEpYyTDjrjA5bCULXa2Zpc4F0UmgeK
bYBKy/VZDF3MakTFWmPyI+Ki0KvBPqgNvksKsB+Sh43zSPcguDoNCeVGCCz1D60m
v6Y4KuDGgixrIX9E84FCx84qNT722ZAhTTXXWojGPAT7VKOyhsjX8NMyHw4NRZnD
JXhDjKTjHx7IiZ6kqhTvoTO9D5IjLErONdcpdK+n1vDHJo+q8jvCInWv2O9zqaRt
vOoklf4WA4r39IAW5LXbFCwuP4Uhn3MSkuhqnTs2Gak3LqUkllPgHonuYHNv93fD
pzvWR0hovNc4J1KPUTq6uhXcCNLtP36ge/CC+eQG75KU1bxb45s3RA6OO6I5ps7g
L5wN9LFZr/usxHPs1iAY4Om2Q/KmPZYS1gun+UCNbOonxK+Q4okDGVEs9USQzCIz
rMd9NbMi1Gqr8lhnGJVAdbnWp6lrtH4saccvwVa7BF3xZG4tAHiQ6BgyHemQZFvB
+gEkvIPa2K+x9jCmQU7bcfNaf2MLGuGaZ3xEWRINko6HdwkzlCkgz347diSbLOgu
D4/vrs9CMAkLY4NRCcfr2H0Ln94YfiAQzlZA4Rzm+0QkXbhgGZXCHSyqjKn+a8y9
Y4iGgOR2yAjk1zsjqA22zbbSR02+t2TNo+wXQCajvLD6vLK/aqWQMbtB3dtvEaPI
8cGOq46Kjo+W2Xq4SM+SbzPs+YW6I0O3/B1qoV3i62rblrFyPTmOgaHYsjFOoFVb
TQSIHx1mdsp4cucTXTN2ImGGNUhMpaDfS8PFa0tYrQb8MjT82T0L6nMmZsCKEP+D
HydJeIjngLqVGMAhm+ZASOqAz0KNn6FH6Hde9tj7VH4/Dsk9ZxDWe6wdhqTV5/iP
1G9+mehdwTiCXRpO76+DR6KHT+sMJV1qaW6IuliJmFTNSTxpsC/lIsR0J7g5I6qR
H/I+gSDcIITqU98mgeT6FEeFShMYGUZi+HRAHLZADzigspzH9A9Ke6Eot8DZ24KF
BBShY8dBggqbp+nRStcSpbduynM+lAWYHel5hOuGqr7EgfweGjW+nyT9zXBOaYuo
3zOxmZG2vJzOJPlGr0LFcVmbcynPLjtWsgWYNtin8NAZOs3lDEyOX0or90xzzpqf
HqHI+iYu7lA8WYlDtpzSe0XaQsc3B6fS2nNP8CPsl4UbJbRS7exO0Jz//rTTydwh
9kpO9anhtbNRhp/xQMlSck5SMjSznljyoQQWqhZMHtoGOZAOp83oazLmPXognivZ
5fRUU2Wxk1RsXpmEghuMjzVosSCw2Bo9Oyy+ECuRrDK/x7RITPGK+Vybfn4z0hZ1
bQvJOX754Kq1CxQiSEBhIaFGpvueREwQID4Iz076cOZm234igNIU8apXxNC8p6y6
UeDwPltK/H3AueM+i74ri+BvSSoytvAdFHC4duw+iIZdOPcSW8tAbbP89aYXbYJJ
wg5dqtJxIr+8oarBzv4h+10N/HFINJw2izbpzXttS/riCvkipch+gPBtMVNdCtpT
X7HLDgteNRyZh+iDLRe3ZV6MYqJ0ZcXolBprXcipQeIcDKTrfzLuMQNdQM72quyr
LlOO5ZYH2i3Rzy+vFqnAcW2uCi0F5vUosg+odG0qIlPA6IK4cfzawO2XF+fq/ODI
GOaDDFAlurz3lyHo2uy/AT6wjcEhtrx4rK9xhO+bGkNNplF3NKghvgEApS5x/Ffi
9AJUXYT5pbwVpiTJJ5rVXQA5X0WcqvjzAyo7tlueNXgJe1FpacD7loKz1wHTg0Z0
PkuNwP1Yo2tqn5E1sK9xYxdt8J5KO/20Tv5MMD5lcNRitBtpTxpHfMMk9lyA8HZZ
/ofuFKmrzBDdfGnCxN85NJKMXVlXm7LILAR1AzSXOa8c/e6GqaM6uPQBnsKd8ycL
N5cGZ1WCf0ZWojZ1qtwIZtDYrL9QBlNn3dxtAUt7siSmLOCu5zfW9ReCHVq9h+/+
FqIZw4a3GaLl78MZ6MP5thAtQ4Dy5K3UQKCWYR7DLMwsvXGA4oOkdQyY/DQnJb9S
NAhNlkIeyXnfUs9Kcets13Zblvy3ds0BbdEMf1njp9ca715gM36DucFeq/fl0LmS
mgxqtdzyCx1ON7ciSYSnbwaKyVRScOQyK6TrKUyTgsGNl6Tj5KtlqMHC0LlVk1OO
r++B0pjuIE4atnqmzfiKOFpbljuOImI3SIu4COBphc6BWbsSpuUe3Xdjmlt8qE+t
a692ixPH2Dt5AazsOpZYpoudDQEqxgRcPdk1bbsn3G/jct8fYJ5yRJoynsv03Nvk
x8SsFINelCuelCk3c/LfQigIw3m/YxoS1C9HbiLZMMAL15sGQpyGViRfiUQKvWvZ
O0LhjwfyNd/zwNgSE7tFDn1+PYlA7DiCc4EyRcGVgKOaXQWEfNlblKdfuVx8yfmk
PUGxugr3xTIh3jm8PCB6uLloU9vX0jyaGolGvpICczbQXGKwe+Rx9pU0F7gWoWfo
qRvL3O5Zmo6MA8QBcF0YlJcqPTZ3LgvvE8swmYEvKL2xn9rB90+ms6nY4L4V8eqY
QHY+qVnmkYxuOUQ/HBVQyY/4fAPry2ceEidmWbRjPQ6iJokvUJpLuln8S5os3Y5S
dJAV/j7iDosTEhNaDPGiYR2tNkNb7I41VU7DrLsDGtdujTjmOGthF5POwgu+OgZg
u3VYxbNzvfMvAS1wPtIZJlhWEil5zvuE+sfGyxmweRu+hhxci8RFiW89KGfteG6c
CTgvuDpClp7/jwtORDdDGvIHn86zyhn+e8Dms5m9bgAUiHGIiy+cN2vH88a1WfC8
W4Nl87BNK85HGBz8aYPx895fYqzm3Uip1i5LQG59dYuFQUURqgbENPCxNzFqNHhm
vbd+TDg5ISUM4Q0B9UQUv3tUsBQoonXkBojpnblWdepYhgASNUFXfkj3ubppgyR6
U+l90VzokrnrJwRXsuMRA0mUYnNfV3AHkHxc3nWuFUUX1hFgJ2bqOf02XScO4Uat
/e7BwnE4zgCVT/hL8biOzoC8f424YGkMJXphZkS/sAu81BPDIpT7vr8eZb7vk5BD
BeJKZv86578r5+vPi+ZoDqbfgHMAcjwnjH7LZxzcjInXjZaY/+ZqJ2XSp0imYMZw
SEwSkq01gtvghCiRDizaIWv9vwQ/DHUkjXj4Wv2+hSoQBu1JOoCwOQ5sdbUtkjOB
kQW42os614KxnVzBCnTaFi2eATwazIa1HLvUtrDM6KtPdUKX2nw8iHRZerq4N5/b
oX78YuVgRsFdps3cuRzB3aknYjtPZzDKcrE0l3NE8tGEJaLKZW8wmYwW1PCYmvRt
E7iCoLqKJWIMkQfDrRXulmcRWRsSo/kH9rD0x9xBmeIb1IXR3hTtDUkGl1w2KFiw
hWrzt/W0T4MH9xyr+htdD87Cz+WIyos4j4eNcaPxqVW1jiqKMbEKvryGaf112INU
+mghHJPtw6nk2hs4bHEWd8mrDglvbGQx8PuoO9kI+izyL4IwIZyTDf+YKp8yB1Of
TIDhp7almatarGqZYzW1MV95QmodA6mXXUa0dDohA55Oz4g0/Al5DWg+Gw4wO/ez
v0IQR6OdRXoMmHd6RYil3LUo0eFsx1FiGSMoQb2goAz+7dcGDxT4h1M8mXWUkqjq
+3g26+jbArcqLTwwzfJDfFd6Fdzzu/zLrtiKu4wtjX+eXxhXUO9+rQ19avpqX5zA
gl3Mx4lBd8xJwXN1b0n5sLCtLbR1A6wZtjFCP2hWgA4zLIbBOAeULs7m2kWCVR1S
+K2kBZmkbfYW21UYqIQW1+GW4zbsTzGvYYck2F3RXt7zxaKt6pDKhGejeiAtPs2t
xFOPCerrI6m0FNu+JipfeZXvAh1tJy/nWu79h/1fRNT9r0pUDENX4GMyh2rF0xzB
7GOWjepT7HqtTi+0gO/u10YMkM+U5qEH1dWtwaJhpwjy9nDb05mrhgzSEcFV1/Mh
L/Un1eHK3FyhYivMdcv1D8kf94mLlf36rp2G6O4dQJQMbXNiRKLjOaghoviE3AK3
mwJhLpWbSSD/iRa5W8Wql+8cUvoXxBBNaLRXC7jjikCX4VzF6pK/7tZIM1UTbKUh
1JCom3mdFFX2uS61JXWb6SPRyhzE86s86kgBrgMfRCHWeMGVLw7T+Gf3E2QhpXIT
m7GR2lmdkaQiHW9cWzJDbiPatRmQUkaZAtE03+eairM06nf4RxYBqSbdSYpKXCXs
4kYaCBcFKTKrlKCVXNIBDDiYuGYtKZATUw/dybViL6NvIcejTDo8JgnlBBbrEFKz
lyt8pkEVlNvVxamqY9cIcocX1XW0z+zHdDTM6Qj7W0HgqsJi4F0XHLMz3Q8Lf7yZ
ptxbrI+QtFWvqGaGilUTd9ScQ/2+A8fcePKc5etiBJG3pRti1nrOxX81vrFcEiuo
p9K8b9PabXwo3PG5r6HmtBceuvQX5OrsLtanw7CHoI4q+EQVEl//k7TL7wdyyI+i
82BmiYyimRiZKc+AVORRUN7xTPngqk+rrKQW2eR8GsqRcbldGhSf87fiCBHm6S1u
E/GqhyR4xc9Qmoc+zPEkviFGXGO7zVxnf+RFKWSLdBQSDLDscTSSP9rjou3Y66X2
ssPE4OUxgirqKOkkgZMjODDXm2W+6mppixlXYCKp3CSlkIk5vyIs8rZDj1RhYPg6
nBV3rmQwIqpfl5q1t36g3Xc5vYoyzAFF5H760wMAaTYahx3eLvx61IaX8D8nx9IN
8W5BgeTJau6YpUFVzeeJPkc7EHs3FotnzPacwD8VU/etCsY0tltV+QDum3q5hO0E
QNuDPD23MhO6Zz8GWoxYFwbCtPU+t8OuWmqGVodpCp+4TTJn9qbvasepwGimJ+Lf
TQXxiBk0Q5fx4gF9gjIjrcbsG0Lf6R4o9e8nE2h5esMRuoxNFJo6w0MhjQ7EScFQ
qaM8UW0xS8TilZV4NWrnBuApGumdK6ZpU22qormroTih9npMqsAxzXZoQDWeRcb9
e3GQa0ElG9f9TZrpGhioV+PMqA69iX4kV7394XGtxwIxyxyA+VnYnp83cznp9liK
F5OE79297RcAHqrI4LnxAZV6jgf4dIpG1oeyS4HITTWs6aGOs6gVgEsosHKSwz6y
1VSF1u28Ub52ws5G4TkRQk8ZY1DUIpw6UkV5HfKH7E2WEP/gFCmttSZwFRBQ+wi9
Fw/O/gWInq1AIGaeVVcs/r3BhqvOExVbH/WcDV9Uoe/bMLVcRzZjUjNhFIfofORz
E1BEvZ8q4m7IcWhmNP4BfpMrHXmJ1iMvh3qeGvjH8YUt7HaaAfx/y5/3CyWfyMF+
2L88bhgZEMzLx6hEiSZC2iB+rz5SzKXjDgQFheVkwvzsQZGrMiPtqp9l3OpUpZkE
GAjmnr0jgBEsklJBh4pcXVSQ0V1DHUvEAG4hFx1ZOEBrJ5soJBbWgssGQZwgE6g0
01HPw67r74bBG/13FF/cFmjXKV7K1rVLIAZq/UtqgR+yvEbRQzJmgjWllaGbmILk
KNDjZFJrQoXVasJCBYovB+/cv9tL4dURPMDjYIk8YnCo/2tEL2h3IKauJDUsKGTV
XvKJwNQuS90RSBrx8fU7Gj6Uq2Blq+fzYn4A5tKPDvPWgyZWmthiBHdugHOUCUhb
wtgaRJYl4bI0p0Xhl1IEMXozI/+pCLzUPrJbNVn6caFpTvoyZQ/xEqgx3OdvYrUR
T2lh/ciWxV2g0Ihy8tHzalob9I95t7NRNps/+bk3MVP9X22vi/IE2jxj2R0Jh6e8
9IZ4jU3G+b11V60BVqCZB4fwf2ujaMyj/XHIXnFjYrrnFBgah5dsvMZacdXont7+
9YcIdC1zmXlPvbpvvk5wPYN6on9S9q04SlQIa7tUf2MasGVExFNAuLr7C7taEXg9
WLe+CMAIYSROYK1uas4AnPMI0KMdhP0rt+uUewcmsfQpljaQAtz/ZXaVKcboJJjY
OQPZcT6qUEknkZQDs8tmbUT0hzdwvCkU+ZZz12pXr8AKN3Rp70fEjWMi694L5v2t
do3GRTQybLNFhub6d9PYthZz75CYF7zoPUUoUWgSpo7Z0F4A7T+KnTywCtIgpFQo
VOHrZh9Wx4nQLdxtqEs9KAklnua/fuvtPvWwzfPvJc2WXCeHK9T/fFVg8/aL/Y6w
2d4WbZSfIG2nXN1JDQj5hwncRgVM/WdZhIERAcs7RZLfm+OfqfBwubEjtpzEpb9M
1guemCtPQ6srROAmmgluHsDfRwmwPlwKSJa8VSSA80RW4VFhEutnXguxDJi4DMR+
kJ1NuMttiWhhnWpIIc6rkpixwy3wMu0uvjGcmPmgs6RXBBTgo6QmZzGEPS/SEZz/
sntLvQC4GMOrvQgUGVpiBQzIVqnUqEaMJC+6tnrUBJGS8UKsY4+zCkJrvhDQAPlm
KxGWDSaqayeswJA+kePd28kaRmFV4dA2OBUJLB0blOBb/shcIifCRHR3Eaaxm4Hl
2ztiwMpSQH3GrRsNaHcYTAlfXzCXxnJxVKVmKpGzIb6YF3t7l4y4A8SauPaRyhJ3
c+G0CBp1rRELbCgCIbNYyD1x9luDvt2WNj2WF7qoWwjVAJb92uHWpSQ91nNwsPRA
l91BZt8QjcqCJg5nBQTHslwdtEOMVHJX7ZSAdDpL0PAyRJO4Z/FVWyPh1PCK3tfK
QK8rcvrPLmrX1E905OnRMAADzlp0VZNa4kElo3GJ8s6TYxzzyQPWfaiJwPSgkdce
v3H/mwQ/+GHLledmZL6AhZXXdpkKAWxiLXwHhs2xU7eUGzxQUYyP6NoXdF6eNLSB
LRRGwrBqHVAtnmb5uq6BPvKyAwbuP5gYLpIOGOHRyXdsG7ZnvjUFMJSAgSnKNvG0
OcyGJRjeLpjTE0m6ONLgUAwMvBSazvqY6AlPkveW5G6iqBtTaglXg6qvCZJ92yZm
DJFf8N3ZSxyQWvXYMPCbW4U+W10YQcSWaw9qbp5oz2sVXDNo/8DWfOP5T/ywQPbU
ldx2jCtbz4bZOOLQiBWJD0iNShy8dBGDW+dYrmLb70PBgRfG8oDFNanbwM5Pnxfi
dmKvke4ob0S5d1JJ4kWlEYFHR9AnPXsrQ5u96q0qoEHkFsSVgXQG9PERjWoVwP5O
MmCd7SDkwpejx02zTZQaAOIT76R8QC8TrVvAwFHrCSx9I+DP+veVug8yOBV5WZtG
s3zuM60a2hrd6vQ8QpJPwQGqvE4JQhuN6IFYVw7YakvLRgewAFty4v8LQGaxNBN1
fEyXzIRKYSAK83xHZhHNgHk6Itx1GnGGFAWiCUUFvv/5FNJ/8WXlR27kRLQs1uOr
TMN8XZO1WZKR0iFezl81g/NmbbX3zOyM7x8gMoiNoHQpJj5IBZDWcLGJ2Ip2KnU/
aIIb/n7fPzY1KuCDFqax2hxeWDVFgehmlsV6mKfKTjSj9MeqevmX5U82VnbvCM9A
fRJxgeg8s/RdkfEB8Dgszg6evzhE6IdssrI4CG2gCjv4qVfY1IVA7y20zN5JbO8K
oabe0Yp8t9kJ7agAMp88vX+8mwTYy+wqE6OXmuePNbwjstynAaHtYkBbk/VAuTVa
Ph9k1XxxcdP1yV25nm9AkzRI+Ge4iSexOuagHUbC2zYb0c69mEmI6fr73l++C2l/
duNu/HqibjGw2M681Tu5QdHWxjdE+gOrjCEb46t3zXKo9i4GlatYS+hHXRJJyoW+
Sh9xcjXgBi1dMHdO6qF9z2E+zfv15qxttLDDmYyt09/MFovllLk1hjb9f1+7pnxO
yUtu/Kb+U6llwC+Z3ifFpW8H21k0qd1en/7Jwy3wrYNOWXDKXpPjBa2ivxVpzgBV
htiiErFFPuUU/YXtzf2rQEcLBa+/UE+sTGLQFGQG/2GSN4xqjU9wkkNOzA2GRb0y
olqrPAaGtdQXGg0SUTiXUX5zlAj7EbwxukcMiE7XGxlcouGXZIEEEcIKkRaGTCcX
Vrd+C331lloowSGktkuqkWshTdL+9VjhIFdirSH+joWsj80IL7rRuUNSsteTKJm4
wLJR163sVXZ17E48liTzXuS9/S3SdnE+G3w4NcsYhSWboNfXgw3W8oKFQOVX4s0v
kpptLJz2DaSBWhU4XP1xxiLc2JSYFgsO1+gejN/KZd2vKvoO/MS7kB7CS87D/wDH
wxqPl4KG+Z5VIldHcPWxdAOVmSJpNun6rmviyrXVJrjyurm+ioxDLi+rBzGGA211
xo3m2rP6yjlN/NsYg+7NxzXCBAoNpysav7LckhNMXxbxONRzVM9rP5QJ5IMiF27R
3J/F4tFitNGxwMJmtZTHmXqeZCojUZIj2lQX29DsN4274w+mSqoNXXYRRChOXy62
KNEgPwWEiaqqpQ7dHEebKxijw/Yj5a/X0levRAZgXWl5j1JtA5pNWZ8Yvl0uHdu+
`protect END_PROTECTED
