`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTI3C4sNHSUVI68Ii4U/fccGDhC7Q0ZMRr5lEZX2kQERUeHiqSaRJMTuteTrUNr8
aQa6D1LnIh2IS/b2BHUKQvLwEeprn1PTVckoUOOJm0AVI06lCmSqbDcntQliB9PO
rygRNpU4Vph2dkzEGlDJTn/iIO4N//RfCmYskLBGi/FOsp0mGqR3eQdTM25IkZNh
JqxXbv5iYGMqqUSau7+s35BUS8nDDoY6tYRNX0VA99dl0xjNdefRP/dN4Gorzujp
gw/Ljphy+n/nbz6rj05TTOKQ+Gsb44sMZ2sxseSD35GUz4cOy4shRQpU1AX9rfcJ
5lpk84ydtepTQpesQWUNXqv9ZQBCSAxJtfIDnqqNL0SzYjgtloPfkMSdX6ORtGwC
/3ABeFCdAnp7DHuDrMb0QWiTpROBSObnIdwa0OHij0/9i52XBe+2VOp43OmLr9oG
rJ4ruIMPm+5hbI7j6tnuDS2qHRL9+wHns3QKLRcXislc4QOdEjk611kSFeaJk3t+
39852meX2dlhocYw8ji/LEjNmAs9MAhyVID4tB4SnfulfR9ebOHQIoctag+5hcmi
hi6tB+JJ1tEQMPdqxflKaDWDLWc0/lWAI9X3kLP/7fT8f0ohtYdhaCsM9tULArDr
9ubwqZBKAFDXWReHz+NKp2iHb39lFCs2N5ZcLI8RggHzC283VCU97g3OkWeK14GI
H5dnXMwlmZEms/ehNojcCMi/g9cWi9Bw1D4rcg8SJuL455d4d+3ZOsduGM8nisyV
eiYfXVq2qdLPnSlWSYMi/L55yaEeJ9IZqRhV9qiRORQyEqSh2fBDWkDhs1sahHVA
OaBiBeogdUNmjQYDjCGMZVEsCZIfWm9FmRLLLBm0LE48qE8Jl9aV25ywosWDLcjj
Y5AcPGJ7zyw5sajT5Jmv1acqwCzgFsVQsrmQJj9HOREywRCHh2cgIZXwqywOwqp0
rAOtN5ftBu5/PeC8US1IZ0feWXgPFtKKiqAKTgDNuqtpmoi0vmAbZW34jPb/DMa8
CmZY3OVobRlU/2IgvwXj9lN8eLLrs2RmZhnB6vZetf8ggihAEnyMPuOHv/K4CTl8
L6neo4kWYHLezbfyy7VtcKjKRxQHHxJ5bsQdovCu0x62eXjiAYdL+QCa2sX4hBAz
/uLutbHb4im9/wStdhjwzsfWqkgt3tMveBZ9g8u/afMT03PTeb1k8XhCKzCaz9Ut
Oted3HKNQA/K4eTC6vYIl9kE1nnVAfi7+nqOpSobHOwT/h2NPUSGzJxRmHNoAPfc
6aCQXB0a9KwerWJvQx7Rzj9ZjewAZ6pOmdqYV49507/Y6FdBam9daSYjzMN5KaxE
E+/eLPUfSZSUsjDE934k4qlWTTgF0u+M/XiHoBABL5eO9KvAtO3src+VA+2EcGDH
+d4lSH1g0yvJ7KOEVpuDpVmVdP7v1ju+sT20oY6VA30y/q1NlJ8Hu7/Wanic1hRu
itoSztU7C59A9HRynbOCkRVtjVFpUcwC7yOFcCDmWlhA1lNM5UVPpVwt/X1lO3N8
+MGmfzVxPk/5U0eGs48j5kYQgBidXWuvaKefeNc0+SsMR96VUl1JK73gvJC2jIAn
uMjX5gUfpSPnYQq6NGIw2YMuaeWKPyZ4od+NevjjQ6jlzC8TMJlz75ebgK6ayz4k
TYwh1rmSMspsZufy2CWM4YYfXBv0ZZ6ZJGR6WSlUf9I=
`protect END_PROTECTED
