`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P3s0Mo8LouB8/OWUSgawnESNRcEuuY0Sn4srgMD/+znwxMNeWmGie/LFxhtz/Qk9
LivUYP4lzGybYMai5t0kVFptlh/98VGf06GT5XwTOqnQoKEO8qRv6+SDl5wOE9A/
Rdd1OK+K736TtjWuIJSJ73k2qtKtSLZ4FLwsAtw5JSPt9hKrfg8veNkyRLciFtHi
b83arF2RebZw66cdfdhPitWc7dXwUl3TEfBjG3JJTc2+QBpsaIyt3P+rTLxo0lwY
Zw4jzXzOnsJY/N/H2NsP4+/KKrqsqevUnbVN2/477bX+4wbAHK0OBxB2tjb/J/Go
uYOecBXeVMScWXnfWoRj1Q==
`protect END_PROTECTED
