`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
otvaZmbe483BmiJ/luIBItnCtpuCYxzvBW9ALVORHmqhQWnifEYMRxGZ1Dg2hPUx
oB0LGk5x/ohJrS9vj7hiUI5IvnVDiA70fgWwGxXd7+NuSzzUZXeCiBd0pK4cjmDu
/WHODmSJqY7GT/FK03PDQT3Ci+DDcu8bj8Vnb0dLwJ1cgoK9x1M6gi1paXWjCsg+
c8RtPcgaTQ/M5IvW/3X6CZLFm/WuI4E6pJt4Vb+t0QRpe0xiCroGArTKvm08feVU
rc7X3eU3m3YkIpUMcyjy8KkXi1ZqF+5prKztpYXtFCO8heINbhbjqUSKyWYprIs9
ct+3i/HxQ18amRC8K0iyGUyqOpql1CFpwElC1DpdzKNewnwELuzecGWZ2vzyVx2X
ltBfJ2Tp1K6QehchgmyPqJ0ieYo2guO3DGGdQ0gaDEq6gQyvMiN38DS0A0LcqkOc
LyRy8w5Fi0sLRJMl9v1v6GFEfxfocVcIgjsObxVjt9E+DLfdoQ9gAOHuc8w5Gk+5
VSpTvLe9614jWGvH6ilRdtR3ci7oPFZO7DXtwxX0Obzuqo+FAM3oxTNXwyl+E4ZO
mp6a1zhQXb/+4noBOHlrbcbmUgmv88Qro4KW+JTATy3iGKPKvK8wy8utGaHjNt7T
q+mz0zVIcQumRaX/rLdRDWaH8mvlXLbjPyHSXE5+0NYW9r3UfxzWhfYMHUz3JD4s
ZRfcSXa4tgXVWpKdJS8RD/SYiqbDeizZD/hrtRkewsr69/Fs3WNYix1MZc6l1V+M
yQRqG3eoE4q6rl+q25GlZDigNXg/aCcZkjT5iHPZ8RuJ9hnKqbbtqAJ9d8CMVdJd
Kxznup8caygBYrU8Pq4m3GR5JGsxGMUwZw8VSnlME/wfX9H3wI+J8m/Bq1Xzkwdv
LqSc7RRnkjWpDuGZumw9UZ4IMBzJenup+/HpONB5jo57IgV4RkefFUkU+bnLSYS/
2ZNs1vppX/ozbPjuX034WvpD0EaaOV7tZq7S6dhCmYWVNhgQwz+Zed/qR7R/k+RJ
b8pCq0RXuFmf9ki8LkYgx+AATW4zLOs9e+8xfKP8G4cAq+CDmPlGgRQm/xLeQjcl
kbKiIhTgAaWbwGVrRdgohma5+dD7O7RG6zA7btEC7XQtwX23ebUcBpE7namouN71
SnCUVRxeK9CvLTopBbh5uiSiZnihI6BhpX/qIqP4A7kliO+sXyJCaUXHgD0s8D+5
m6GdN6ybRl+RWKlP3mDA7GNhjrXMOZzU3C4xP6FwIZdTZxB2d3m8dHZnbNCF1dr4
IAYi1MvtM9rPqX+AHZtmeVBgTxuQPMaFlfovbEw6kc+NKUs4TlN727gwBy7/4o2m
2r6PsB0vHflFxYkfKRLRpN1WG1HbwUqhbgLuyKq4Jfi8/ZBEnAfucF8G1R5xnPeq
Z/9f/6ohde0wOe2hupnSzhBzegoAPb3W0hhUxxQQIE4ndA9nrrMZM7zwYbCrcNFB
fj0VpFY29de/QWJJ29cwSis6u5HIIll+TMkRUoe5IlWOr6d5+h0wHiyn1GzbNIR2
KJ2XW+auG4owlSwpMhHbzJZT9FU5UOlb5eQfFNAlBLmUb7iITJ9rSrrAYTRxiMpl
yUYwOnqHh/VGKpmYcuVIlYQ5XP9eYKk2ENbt48ZHqVsKCPSrDcHYQauNY/8zEkjS
FhqzBi5vbRPnlXTVBrlU1yzoypmniCivwsReEZ4KZ8J1o1eUg/q9pAd5KcM+9xU5
6Zq09H84pMZrRspCercUkHNAfwZ61UujpPFp4AIfAkCqcm2aSSOjOBHnpVa1qZU2
`protect END_PROTECTED
