`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVnLybptWqvexrlPiXNylmA2pk9eAZWdDGefh18vxL8m5JkSA4hL1P+9AyAyGUIF
DelAkZgKMlZFdU8xhEkybE5O9u8tRh9SPygBEmFiyWp2ptYUnSxqsrEoMOkZq0gL
WgmkWnsAf5wikQfW84YkPnaXSYl8QIzRxZMJ++HO4xfPidEvAXymAW9x3JI5VIdC
hSCnKCFiwUxrTdTG3wHbAQujuYp1J7lW4EsrEpleURpiTRRcapsmeGvzpkaC0X8d
K6O9Y131xEsRj2PrTlbA/9V8O7pPLEwIgYRU6smLX2mxiAlVPWcet0T2eBvt6Lsm
ncY8TvcpeYzniEjZSZws0Us/m4vP/7g9v01UOnIDxpK1zSDSmf1tOSBsXoGbl4RR
gFCXe+9Br6PbMqm9pXvm1YGVq/8+hFTgUp/XUGsYUGRPFTbfWU82H9dlwX3Hb1g/
YdBqx8oRIpWIJwbdVU9OyMLssKpAKYQQtZq1eoKZn3UqoP46B/P69SzwxAJngu+k
DCLjCEYBcOpFBG8mMBXiUi5I3pxQxrSkJeGdGoYPEfLbGR9RcxUOhG512yy48dpg
CI9QTYyxOhuYHt+4rsotOQ==
`protect END_PROTECTED
