`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p878LloZ6MQPzOZUV6bfsVFsYBFZ2OtTBmSLR155GEwkIy7F5371wnJzzrn7optr
vAo+2NP8gOAng/PIbfL40RNpZtl3ExWV70uswoS5qPMrCRDw4ehYHIY/AL4ADwPv
DWEdILhZ+ixIUpF1zFInFQEbHi24L6k/iof3JIV9JaO224nF51WlMgaX1VpQH2G8
wiMiq+9rA3pHpqaaoOx5ydxAlcvnbjq/mGxjvA/5X37NXsCIH6zLo7JMAqKaB3r4
Vlbcu9MX5NP49RZ9Zu2Admu6X+HidDK3DLAVXYSvrJTIIjDzGsK3MM3yj0Qtwxv+
jE38jK7CrRjj484FGAvhdyT4EUkxQWQNCIBASsbWoj5PpSgmA+eyN4Dla4Q3wI0Q
HWiJEAhA7yC4II5p64c7HvH5HE7n6+AeDzirYn1+QytJdebtShqFW3P2bR/fHGqM
ot/O0aRkWRIUhL2RFa2DWQpdZ6x4V/nhwFlANOqqn4YNdnHKH0ye0AGRC8Xc7nvn
RMvP5ADsbgdbT6vJfI73ILUQgG71ugumsZuIko8HVyldDFapLlQzYWLOh6pgKdhb
ErmDN2XfctSwiBl7Z0X6ag==
`protect END_PROTECTED
