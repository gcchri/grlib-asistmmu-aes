`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrjseZHLX9wkwsGZZ3IDHi1lqDFfJdGGZ69DoK0RoaBphjCO44heNYwBPH8/2dvL
WxiUe2LWEdWCP6/1Blv9NGujIGkKdg7AfqxUkjnoUD1PhJTIGHKx9l5JxmnlSDJX
z3Su3nBEduZFaOcAI6DWDuC3jpJftzD041/mCiDjzaw/cn9q4yB8gy1ANfHR04Ha
8L2YSbsWN8+G96FQxIeGkZ28cQn1rqLLqoSZ5fgpU+n2ZpSHmvIIF4seCaA3jRZ5
Zv3CLKJhl+lmfhWWmiOjjYFqXFMDH5GnS81/TA7ARYzcKg4gLl2i0RXZuO0jKrBM
AEyfMA4rsoTYUDZu5fqM74dsi/HQ9mazw5JY9eRhJTPLzWFAlGviwF4LefWIKiyD
`protect END_PROTECTED
