`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZZDfsp9OEPrAURIgICep8KH/AKf0AxdIe5X/llaEPnlcffECdx8M3uzK0JmXsrSh
z6C43NhjrvqlNaZwVhguZOK7OwaqGKxLhv3hQAtam7V+eimrocw2Dp6anYmidMgk
4odGJx4vcDXgQSdlAl+g8mDuQmgJG+r70OuiQCdG0/Y+tiqE7nkuuwwY3aTwDiAt
KGFmvAfQa3zBB0MV4sFCXw9E3K5tehrc/tP7DpLzAzTWZEzVVqN1Izc6TQFoRurq
JiJ5xJaA4+MCvhVC8f3e/LXRs6gyYS67+UQg45hiXtEoYoC8ZpOQevVcSH4f97ZZ
DRUh4dOnTOWAAgUkOlZ1s17qKpujyfTk4eKXH7AgD9VY4FhdlDYgsutYB9gmT0x4
ccr5zf7xBEbnbS9hIezDPAbhtmASFwuUX7uqDrrw5XZVCV2Jrew7lYLOPITLf0tw
zEhMlHRBMSwOOUF7iZaYrOtFP5XVIfaJuqit6fcOEVSqIh0twsxzT1a0a2D4qY3P
CloDck4fFXk5F+u0Y9PkntsW6cazwEcNtVZgVwWL8lZ55TQ66xVdGiRGqC397ZXP
/Ho10s455YawBn3zqpN58J8K1uxib4f1EVLj7X+mUllwaTxRr+GefyAPOp+pDSQq
DfoUcym/k2ZYZXv9NeOMAQ==
`protect END_PROTECTED
