`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QcY5q2qpUdalDkWAiP250V1MQwTQYKI//jqiZ+xiyP0JQ6uTS4pRh7L1wCw83n7V
ES6BFjjhNwDQvrjzJ2U+FO2P+evlNzuxseDxiBoAguQaWnlYdxn2iLRg6Uf80OaJ
zZ3T6WqDB3T+ml7FvXGydxTn3qM783BKt+i4a1Dv9B/SHt6OwYCM9yDWQWKOBnuN
AOkEN7KOLz+T4xr6jwB52k6U+vO512WlStL633Av476ACXIRH9lKAzpDB40CLZB9
7WpCFuvUUIO2ve/JGlF6PW+6Nq5DEcH+fSc3LBcnTd/7zIfBkXQNdEuTIJ5qMOx5
7QiwHAc1fasNehQ1AtWoxL4ElamhFbz59sEB2Z+g9+/NI/4WY+crmKCBZGQGBV4m
neePpD3YHy+xdUzV2mGI4au+ZyGU/G/4CKGVwO2EQCvtHwwn7ltL33Ld7znB59sm
`protect END_PROTECTED
