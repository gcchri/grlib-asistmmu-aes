`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
87luzjITCCr8Pu8IzqX2B/bSchTbUwT1yjXg+uzFu/UfBi/fE8J+ukziDpPzN74q
xdzsxlz5idq3P94rji1MUDsF8UUL4Dp6wMtvnZCN0gESNF3ADqU2qgavTWsVGmEj
ey0RmQlJ1dC5LM0D6A2WHdYRyHT4u37FfjeI2jy58ceN1ECMAPLOWLJxPaoGbzu0
aABJbww5LuZnHVo5zHk5yUT0Wzh+qDIMsWY2anJuj6FSuM5FOXxktu0lXEj7SMLo
GdoxxEpoxGnCL3XZ7XdemwmaKr1zVmdBPtrfDlGbvgiwPQFj0luSRvFI9M0Nqol1
giSe7elVy7dR5GDDwEzSYZqf4WSFXfhQ2x/j3IND9bSkNqH2cy/g2YIBkTdr7xgm
`protect END_PROTECTED
