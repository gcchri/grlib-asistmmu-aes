`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2lQSz9/h3GBXpWicxWROdUplr9tBz0TdLS12ma/jXKdupoA9tYJU3auprLup3FQ
3RcIPidUM1RedEnJWOOJOwVqpVfxSUGA5kKqZWTIU4cepJfAXOxTHZPrRWVrf6vX
YPQY9cj9oXkh+OjtlYhWxPVWf+Br+kHGNyr41zgC6n45oLJeWrcFPOVqnL5nvieq
Lw0Z8A63gT9NHz4UxCMFhV3MAjNBJXaacdcyjMeIUWPEUb9WwmqHy6kF/lVmXzHo
Z/aUg46dBiReZxBWt1SQNSyqWRxEa3kBabsP6lLuZCkdM1Nhgm4y8UuptC1COrxa
6TN7SvQEf864Vq5K9yBUCcIKW4/l+YgPtHVI6cIW7BI=
`protect END_PROTECTED
