`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kf3nChAcnSonK/hLLa2eQmLpZe6d11K/RppKZCuR5A6CW+HzAL59D7FBOrgoHi/H
SvTV3qKWcqGwknlEmNROQX4eamSy3TjKyPpK88awiRQmP5Uc/KiTE+Oix+0H1Jc/
WIVvJnwg531y0kRTixqWWWmgIxPbc9U47Gz2JdCe3KH3uTwuUaZNqX2cOMqX2sMy
nKr622nldoUCFsmpHtlkfzcCMP5Dp1HF8YYSRqHa18GuNIExSCCSTqcGF1PBvYfq
qWanzk0ByrI35lw0bDkdbpJ8ynoRObHWYPfmsTtYnNXjHCWcEb/4bbQeRoOPxIPE
lwmOXTBQK5I2f0ld7XeBmMuSdA1aEsgdpJK3m5JsbhTr/MtCdDglXqdPDzRlCE4g
KytcnpsTFKGlxo0jMN5J9wZzR/gwjNR94zWlZV7sa7GD9ewEYSi3+KykoOIcRN9U
iprgQn/7m8LeSVXTla9cODylv8JJtcya5/a6XpVFFWQ3wCqYByJZFoYWwcboBXrK
ESqEFDUY1Uv3efeLvCWZkDc2wzx0w50M0whkCapuG9NDsbBW0rP9TRVyVGTyDd5r
sjfp+tRQUjk6DBu8ewq/nwv8vTl2l1MAHEqRC2D1FVev3vZmWqdTRN10qO+hZlBp
rB3p8CY15rDjTFe0431N0hwsfdjp1s8rloSlIbMIM2cKYqzmayjxlEJsy6evypu5
XWH7TScZOZJVqk6/QbXJMj9Ik9q1B7i8t6QBNLPP1MBIW5B2u0kLVR/3tzlxNXiu
GzNyo3SkAMXBkTKF6O9los1QhwqXbzgalq0yBAI74Wcc1UIFfpsTVej9qYQ2AhsJ
WbLUvtT7vAua1dF2XHMQR2Y5qZihJ8+iHHzwZ005B67jvBC8oju6Zdq98kOsZRwJ
QRkmPwG7MtOccQVzIQ4JsA6uKFFpdPT5X1k4PffVQj8oM279uDsSgJq6YG69llh9
Lv+mH8cU1r+IAydLrQOXN776/tvcqeDeySD0yzIEQWoQecK+ADpRem8YWJ4tBEoo
vF+M96PRfx2LRlRXzUpm1b/EI5qX96DdZ0VTtxLBB8Flg5NaxuIZq1YoI+46QSW3
CwKxtcCcjHO+BannAIQmJ0AHwq2nzu6TR8w2MGUvK7alwDdiVk8bpEkdlYWOF7sx
duFPOqfsA+GE9I0gsNonOQ7X2tQH3RWgAXMo4JZ41eBkFHvdO+yFYuoY6tavVa+L
m0s9dPNAL85RRgEtAxosZeELG9gvpfPc4xog7Q0N+i2Jmvv/mhQOFDFWhkeidVjv
VJXV/LQ/njL1mYxRUr74wnx+LNYL6KxhmwnVEd3nHbenu4jFj6AF+yGI52s3FmLC
de18AlnMGr/upAF8anx+IMf9zSOf2RPYX+1c5J4Ce/ZoQc/Pyf95hx1T8X6QbFMN
aDzmdSWYO0aGGCgIPYQX6R8vjjKhsruJQi6U3PfJtFgQg5Q6cVMtrrPJ77FECzXF
XbRRhkvM+GQaiG51w/xilv0bIo10tcOEn8thMmEeEZ6SxYf9OiQA4B9PnnS9QpqT
W9OdqHzkWeA7roqTzrDKS9h5IUCpeBa2U23tsVv4OttiSOkBlwBThnUfQRJl6omU
72vD+kvPUI+n7tlphgivcbG6c29SwTpgU8oPQNGKxLU3YmuFJk+qUOhpH01Cjwsr
tMHMQz5gxXRxG0iJCPy+MI+1g0yWMGt4ScdpBJzVph5yGQ7v6mSArUXBEeia21Fc
rJj3XJi/9Dk0YRI6jBh+ofucURvf8kyaPCYG7ljaPHBX3PSUne9WZ2Br+Ei6GtUF
Z0/SHJSssEiBK77rExlBYMPKQeX8E1KdYlWJmf9QZC3bQ0JPNdNs8MTT21YE+5eO
Rwzbsft3sDiDK5JwM0bpUE+BZTcjT9BhXjsSGN9wd1Nmx1Fwzaks1amh+u8bZ6hr
ngGFcpDZdGhmrJXth/3kss95vX3ysMVGlACIhfqpBPQyOkKH0rsj0TEW6apcFLrX
JwicFcDKYVg9eWQs2CbhlwUwA58NTyRzokZUdW2vVPtUYjpdkCMr8wlL0cxNjVuh
677qAp5JdKJiwPwfhYva2T2eJVo6fiW3mgnyx2ySyK/L59l8IYkCLTJoGuB0iFM7
QVyuTj80I+3tp/kRuOUPyjUTqUlX3/RA7rj3Ylqs8e/wBJNuucmWiMmnFWd4KuFe
LA434OVggEglcqkBu2n5ALOn0WO4NnXwk0iH/KuHDO8TTsBhm0AQEu/MNXknCi01
eT2RJOCFu8b5sj4oMb8Vy4T2rXV/izOuSUmShF2xVbnBqkUGqOf2GA4z3hW8g/oV
ObbsOmnDC0LCjaH6zTQpsSRc4pG+wavDxUo1SxNOTD7hSSJlDPNjyCu4wxabGSXt
G68Tqk1TfyQUqYBkMw27+KM7thKklQrKO8M2AZ5KbTCTTCwtVE2yYRupy2k53gCL
mNkCbE8G8TJ5lsQDHFBJcs24r2obBCrhbKMOitH0A1rgFJ8xIb6FnTuCQcfyudos
1i3tWYAwNhdHMyd+h4p9FrcH6duipLpAAP4SMKSVTvXdW/jg5zvof3nHyl3AEPkW
I5Lc/ak2jDAT2KkAB23T6Vy0O/P6smrHT8+kcNb+XraJvULb5uo+ukEMYCk36lU0
zZqLTM+CelqO8u+/nLhs4rui4j6vwPswZ2V0DOv2uS2zV7IwDp/KX/YXE4BCvOnv
4nou1r+xhgwoliitBl01TMEpf26s3+iKR6BMebZQpSRrBeDga3XclypR8FjhZVkL
oG8J4k59vgveJUB/3etxZhGVpUcRNPk9AagSw11p6WR2yzbhNaCA4c6E9+dx0Aic
E2jCfTTIZsdNZVAkYYNI+tEgzfOrS+p5PlzRQzjgtF0B5JJRvoikKsOamIt8htog
eSWJuSOXOmi8/0OKZgQ2NKURstn0aKzNQEIaffthCYzpunGKZkssWUNyqpvC8S+W
3Ec1pPq6Nifp9fA+56Dy9eTvw2p2DGV/WtwWsiqCXFMCW40aBjogrb+4MgTdO99J
zMRtSQu9oiEV3LJ0T6OvsAEUg9TqhmtTNc64BV5ANRnAXjcbaKBbR1LBRuZhgt0P
DF7rj6BcRcQnIQmEWRDcjkRAcr+a1LLsrvlok5/w3+1uVyAYX9uK4iYQtK9nm3UP
oAk72LyU2VKvRzSporoDdfF/Lq75kOnwJ1LKby47RcXjkBEnbfvX/vk1Jn2z3cau
fq8eK5XowRTpP+5dH+uy6VqkfzgU8mPp/gyGQydNtsf1tPjvIuekKbTFRnx2KSQu
LqESWdJ3EHhPq18Dnxh0dDcbT3c7vmx4cSQ6ZoZRwub7PNiA+d3FLhLRD38oqoEP
8as/vwUoh7a0Mxp0RbS7QfSFbkKduNzqXYN+UU4zcTuxkQ9VUMYtN3sBMtWL2Vq6
xmBBseK2P7QISUgICb8Nwf0fPGy9y8Ic95pKNpZDRuppyM7CTXX6ugEG2YGc/6+y
OS+q1Zkm1wIfFa79TchL0rVSyhR0albl6UYMaDGGIUds86oJNgqeA6lZhnk8fCyG
fmRmH8vcF3lkWGNox8DKzKL2QcFdASwxt9h25K69JX3ZQ4sdb1pMDlnkjR+z7r/Y
DA5eu8AbnjYfJ9BPEfbmLbZOlQn4mL2tvsjWP5sCsSqk3wAZRwCamg9Udbv+myiW
PdSZn/ZQ7QbRUfcRaktgMLaxXtKfbQ53dAiXY01a8BLeRVJxp98++882DjXEx9MH
oSNvm7wH2Bz9/pbZQBssf2bvPNTBmDgaLh60wXACfD+1ZyK1vPc8NAChc16w0O39
lWe+WFdeu33k7EextvjNb9Nio5OcQU3CGWDVcNuNr0kW89E3W1RrKEsy1bZs9xNA
60Btxjs8P5bxmyr4eRIVjPw7AIDvuO2cA4FTtlFcco1K//wnPEePlZCCaYIUPMw8
bFSDRf6kpgVHVt94sQ1wHZqKNHWycJ06kI503JIdXH9dkDA30vOksrYOSJrGrq3L
PTqFftIiTwGhLYx919NtvfBMpxMeIxWocDyUdnuv/wMFzFMngZZY6G/3LWrjwtRt
H5vGFHlEMj0ihc9ro7WSjim+MTa65WuOcXHw56ZCNWMPAqM/3ecdsRi6UW4Mxj+u
zdrWXT6vfH923fk6Dbfu9DUxUOITVh4OamGu/AxXDn6NNFCJAKXWtAaf9T08otqP
UtS3B7NG2EOv81Vl+1uUAWnNI0xNFY8OZ/WG4SqE1ojsIeakS5dFXC/z+1zA2PN8
`protect END_PROTECTED
