`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdXlqy0927hQPQahHqWlYhtl148OpgbJ8dAu3iVCSwmV/Vhx9PB6RvrlfEbuT8Xf
ksLrpuULLpP4lSAlvQjvl6+uDsk/qmARkdzbiIsB1MPO5w4RzJlawQsdlGFScztQ
uzLZ5QFpR6CIvmU6ub6KNC2aN+F0pN6DoYOCXykYHQ3O6HbA2uYzwAcK7iteNCTJ
dMbibkoeQVQ1GGS4gSFofv2Kvww1D6WN+PDaJJz35OutOfYwlEuZN0ih6vi88UwB
PmYnWf44B70jSeWqzQqO63QBfKDP0UEIXy8hkc+500ORxvGpGbImVxeWEeNbbCil
KaVeHuxS9cqjvPAHItGAiAkLho7R1GDE2PHBD2lHZWEvjJjG6cOFcdpq7Ei/u6zR
FhRG/lgneBvFXJV0QIPpPk/87u4aoyccoGTrrBEwkVPtqaRXzhgAztFUajiUZtc0
marALo3JBFEWc7CKVap3TcMivTMwOn23/+Maj1W0YGHQSnSPBa9dmrnIFBoK/K/w
Y7GebdB6crgufIDn+TASoE7eFZavS8Ih5i8iLkxyk30kz1kQdCAwM6OPtGVszVIg
z9C1Q3ApOrdUVQA/Hl7uPVUCHKuBlEuo7VX0UpcCsxZFqWwXfiY6E2bzlZKAXs0F
8RXUcBZI+GoNee9zRZlrErB5X7ngMGXNEzT2dCzMGQLUErcnosGdFPgsI8/OQd8H
DBU0tlCi0kFJrFVHoAN9gQ==
`protect END_PROTECTED
