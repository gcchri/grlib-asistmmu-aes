`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ohEK8AMkPNkV+fiEsaa0odc4hn8rWjnFApHBWCuNbemkQnMoqDf9z6ADL2ypKhQy
flEFWI0wd8KebKCrfgum26jKcrAxFc3H5ienSzKOpgAySrPp6w+ZURN/AVTci+Sk
NhNbeqpQA4et9gcmU0w+WIYQL4m4TCtzxSbP6jF4ZKIOnAkmZx6kfH83eBqBNK9K
lYRqhtgjWe0ab9jD2UscFYSMKgdiwxhHpLkzZBgGXzb0byAt5hrKeMkP+1NqJwZ0
vVGZm/Y8j+2dvuBTpHWojppsEWJj0lWt9j0W2AH/VomGouF3JlyUVR0BbfEnMs7D
7O0O6VngtoiITx6i3BECmutB06B+ADy9EYlxOcDB57m5xexyrdEpGq8RFdm2ptEk
CLsPWfJgOXsmEJIazDCJm3VtsDT2MDGRrsWIvaHowKBAn28zdU+DdavjrRv4d0Na
RvEy9VTZxYuuShnmB4zghVvGB+lWaC7eU7St+mHc3WXNJ0otwBL5tkmEYYjaTNuJ
qI86p4tAI3f4FBbdoNYDOgfCkwnkjh2+n2Yix/ms6q4qjNpx1YomIfKbZ9RqrOKB
k0xWk0qgKMbk4r6WeklfFQ==
`protect END_PROTECTED
