`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ha1m4RhvlSYDjGTn4IFvuxUPh+EM/MnVuT7W6P9xt6i86UZBptnXiaqBAYu1iAN4
tvRFoSAZCws3C0USKu49j9oXJG+uzDuamnB+z5y+PKUjejyleW+OqPlgdtFuFpU7
itX/LwbkfkMVkpj8LvSXJxlCPln51LyXJMUW1DF46mHd8Yp20wvgBK/1u06TEF8G
j2kSQPUPvHN23zATdi3Q109mfKrzApiTUA7PSkZwSDtBe7Wmr6mj30ejfE0nLMjr
JO5N3vyRRSwYwIIotfvCQWVEqbuNE+bZBlADuejMJAzQbN3nBZxbT6pAmD6beBRg
N4EDpB6O/l3cXkhxJuLLmJQKE/9gvcCCn/85e3ga41/P5dzNztEGSN0Y+rpBQY/w
u3wr3mo1KIAoQP6aOofT6ThbOv2AG3pMvwkORQvREqwg1Al6i7dhzqlT9cv/RP4G
irxh1IuNaOVoUnsCtfX6/fSj+Ip+aR0hmiF7ET47OPQa3ua4WVSFyRtEyhzu7Q9U
NyD9ty2Tg0pgwfPP2mRfBjfMTKYR4u5a7zMCgAbDEpRj/2Fwd3in8O+Iz+dzgL9p
eyMPb4/f4+cJUdy3bJwT4/DyrQTxz1zHq5/rDYvXes02Zcav3WEoBQRCGLvuGeS/
DpAW9yDt1ihN8SBb7OzDM3hbMX8yuQ9afbd0PRti+9CQ/SFvcgBPj1+oYhVKOSz7
rzMtv4LjhzYkKHMIzZ4QU0Mwx1GdeliNu913+A8TD3I=
`protect END_PROTECTED
