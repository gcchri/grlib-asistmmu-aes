`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z1H9bwcyiJbvyw2qaLctwc/4toBVFeNmXUnezg3ILIWJ8ZqH7mB2n4Se/wDpDmV1
zcVrSIurgW0PtU/ZRoXcvFfxEANbgQL7+peRCWXgcjTw47Jf9vWajdT7wmUvuqDj
RFwWIXGL41mhBFQfTBGHkYzgpuu61k2IznAzgfFYLHDx3ueOP+alLRar+RcIsHe1
/N/fRye9AvSTm8L/HC3r03ifbP4y5Rmwoic71F4b1ehf8Rq4wmDOVtE25ZDnH5yj
a+tmqVjdpX4XH2IG9yZke7birnYIziyrB3/O7pFx8Z9H+SlJjdnIH33/3U3wR7LA
nF0tzjJ7gRkkdoFjJNg1cw7cz5hxRbG+TxIUGUgJNqZUwm8UiTLgS5pEhtmMzXRA
TBU3pNpyjb8cJEqvzhaofn8nVyeAbJHpwq4lOWGW2090nf7YXc/46kIrqltg4rYl
VhT+3WBkPnkgp5MATasRH+sNdWLL3bu1dW2yPWLvN3+NFUaK7e5zcUieAKXqAEle
epbPD9OICNxZ08Ry7WmcxOl6S8Y45li7makwMsHWZAtyDpmL4SBQDBSIpZlGjnKr
6QmwBlksleMOuKYOiknN8ZPjwsBO1K0MeJozBXhTzhk3jDFjs+rH8oE1pWzDzawy
T49PTyYtC6HxqM0sK5dU1qZVQCYF8KUvckpJf9PiTJ7hk5WvX9z1mcQKscUqmXNn
XsREk/EIWAZ/bAPDpj/nwgapUVJApINRY0/vnfholLsKu6RPNS31IKGjyezIZrRW
NDRbQ81c4YTqworeBqU6irobBqnwMgrUcElBYsVUFzLYkHBlrT9tTcGJu0VTycBH
3D6yJ8BnOA4IkRNi0ru1wGTkLlVRDq8WSC7qCemQYRMmID6vsPp60qZxwHQ4ScZV
i7YVpalxnb70UTpsB+ey1bZROt/Z6zyWh0dJ6sQzkVA+9RiE0robX7eXy0xTGixQ
K0Hu6FtWR2Snk4KSyUN9s+ka0oLK3LiNSJzO88aTZo2VYnx6VUCK2uLxI2jXwv8o
h9wijs5WFXbjEz8f9Uy0iw==
`protect END_PROTECTED
