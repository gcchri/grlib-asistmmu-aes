`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0FtufQMFJ2lMLGCFO8gPkjeDBtMt1Sca02tLGIaq0bXdQsScYEugdnh7LgzGs3Ew
LQPFJ6IpCvgsiktJdr/3nkCuua4FZKbbawXcbGHnCnXn3awQBXhbrIHKqTOW3iI2
UKWTEpgDGm3pqkQmluCGlNJ/mDVNBdpN7zO6qXRfRBhwA9EWtVmM8xuYaKCrjcFM
lVaQsUuZkghuSjJaQdUUkKYkLzXvkwgjY0rosrCOh8BNxGIORIZ+6b0zW+/yxHbw
GwpweUfpHYN+3/tA+9JK4vwEuz37Rbpb4D7kZnNJ/sTYLX/wLmZGabac5W8sjaVq
6QZl5q0Rqp6gkeIiPWIHd5/qpCkuzCOMneGmAo4MiQwybdQWpjXcc78zPSveVIae
vSXKU78ytE9R1zt6LCbGOPI7kvK7EVDRJQskF/Cz3z/3Pmj1RmU0BvHM13uJ2EJb
`protect END_PROTECTED
