`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgxuNP0slDKlFmJ1PwsZHcG5l1zd2jJ7Bdim2EE+OoL4Iy81nM9s1oiSsvvnyfBG
2OV+K2GbhqachguP3ZaviDqMtlMvSovyL5EAcdRjtp8j4gphuib44Jg/RY9stwuh
ufftyHmh67+wPkss7n/ixEHKpfOAFUnhynpgMRnr0DLHXSUCDzvb+0xTKh5WkF7C
L3w3NpQ12SyTEOQ9XWMRotOCvp8qbAy0g7ho1G20szV4UzzRMenJtpizg17cwAhp
7+UHKrXYsiONvskz+CsuGeNIB6MMGab3z0qTBgCri2kVokqLdu0edop+Z+2dDsHu
GSUByK3IYPWw8YE2nH1wAgt5C8vYh3HnOQaD1CnLgvRQO7U0cj2K092kUipbVlji
RQEL2TB57YyQK16ZPcuELJpjs64vpU/VFnVN9MvwmLqQ9mLlvwS5yx5dK921eWZh
QwixaaJuessDz+GTv+hpFvqwQTrBTrgUsc6xVh/4yvuZlGKmarQm5vn55rw+sQs2
gPSRy5Fs+Dze+XMLy7Rsx/E4j+h57VkHVWJhj5oOGYGu20EfekuW4m4rYYzHUZ5G
jFGEA6JyiycX2mgW2gitq2E8uAQT+5FPZRczxLMm2xI=
`protect END_PROTECTED
