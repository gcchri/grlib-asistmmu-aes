`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eeTCHgXwxIYY5YgvPTsqiRbbzaiwmsuAN6oJMDcjw8kUcTLz8qG0oqDpga3KHrT0
BIp/ePAs4y5IxOpNT6yug9BOLkhiqRe1ZqJAT8OXlyWjStKC5N2Z3O/jjXeJ2Orf
cis8ChJBcnSUcFX4DHEZOQVLa0YQDrITHydAvDSMTkHMQjDQFLde8XCJBgL+U88Y
VRCLM/zbxouQV3uYw5UHXFkV/1oCw0s5GfJQa6MBHw7pzfFWHC7NSWmRtjzbnpSd
369bj1RGrf9Qs9nWBmiPFg==
`protect END_PROTECTED
