`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1W4H3jdJus39OI43ehfBJbgRinanK2sTkAKGKAbzP4TrIBdH9zqmfg04cX0aECrh
XvrWiUEq3XhbvVtgikHV/f35MsdrZfw1XH2xwiHpCNK2vLwkbrx76rQorFojlo/Z
3LtVuh6isaQuYWJjKSwFskTwxkMjU2Cbx8Qi8vTrxuxtbvOczdhyg+fxxY1FWOk/
knhuMHRaBjG3tM51rcY9gGKDEDcXGV5LI2HdFUU7MnjVItCnqSpVeuBx9jqaQJEG
o2HKJN2kNxJ77DyPrxOWI6mEIvS9OIoVcr8Zc/KzxsFqakTvHmvJwtHPAfBbEnaB
rED2IfdauHr8hhIudmeDwR7o0pXZb5wSaTGoybNY2fDhW3ANfpo1PTsQwDqZkpuk
YI1mKqU2BYBYjW1bu9+FQxNUNtbRiGIFw1jkCAPX3ERpUe5SCclUNTOsQM4QbiMI
z72fVRpxX4ZlMamtszXdZLqJhW1qKw4AjjGxT7ZTWZ00BDLmfyMyPwyHYce9zoy/
w4QabEjo0dxDs4jx1FVFaQ==
`protect END_PROTECTED
