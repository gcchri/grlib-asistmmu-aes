`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKdeqsUuTQ16uMhmKfXwf3x52UH+jZ7VkQiYosDlWiOPhFTDIVFGCghIHVd77V4b
zJX8PDJjJ7qxSfwl/rVFVoMUHxVPShymKJKy6VyMNe/iWI76PWsEQLIMbH5iA8iM
BVcHdjPOjqNoYixxqsO21KcCDP8TG+4WcntwJDgWUw5o5XUCMbclDsmZMgLqNc8l
1gE1CiFqVH8+00XYF5atEv/PznSXO9/ytv9tPkIU9Zfi7mKF0ld05U7GewVIu6x/
61l7aGvrYsCO4wHaK9eWkBE/3P/rVO53wPHXPrkoJIG4WsbWrsYmToko69lQuAdn
41y736/H1kK0jKdL3mgl9IQOvfp7UNGziVrWvqNhfnu4y43d92gm1jVBZB5/C0V6
EF4EIuN0WCNZsFXA8Odq7KpAMG+S01IsMaDbnVC9fUTU9PcVAXIKH59NPFQhLWbj
u6/qPttsPfjDkBqQx/QlsOFvEDJcXpYh8Uk/n61zOBaX8TEAAY6mksxwclb8AACu
f1g3ORGkEsWi4yeOEq7XzNtSQTIlZ507ddWga5XCbs0v262nisuCe/aQ0OMZxBx4
AbkLO4OkF6jhVC1FykhlR7Jk4V+XmeKwwNXnigINyQo=
`protect END_PROTECTED
