`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oQDLa2cWbp/tdns8v7aLD2DL3OZjPtR+u0vqD2hWdRd/5BDuU0tC4ba4dNH4tk42
LWpgY+7LpZW0gNL2g5eNdOgYPk7kh1mEuMiAcDfu3ogf3gKQg4JFIXMrzc68oMn+
m0OnRSY+Yr2hYxSL5CJ6FnP7OzFePKF0O4JdZbYwDMzHLlpZlJZHs1W44bHon/RD
f1m/rCfs/riAxeRW3GOnrcE3cYY/wQpj0oatM8pohakvi6BRty2x8btunZ0FlARk
`protect END_PROTECTED
