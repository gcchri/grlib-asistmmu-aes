`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zc24gDBRyW3pq++wIWkLVo0meAECG06sf6sS1RmcAN9bVXMB/panqnddngwRVE4r
EXxZOIaoaHlmOCuxk7/xrCNGquYVwrH+IeBm/aPNO8KZFUiQJKaZb8IvDIyPsRyu
wP/DlX5s8Bp+0K0Sj2DpSYndoiQJnx3YVVnOUpD5Q6ukGc8rngmIqcMxH/mqH+Jc
7DOp6oA7yOm/rzvKZ/C0rbl+JYYUEGN0SnAsa1wOvZm15SyWKGUpKDc0Q23YHBdn
TfHhcSrFHPguGivDx+j/UA8wMF7RpQzerQLyRBq8ormH41adRINIFzEz478rHwF8
snFFF1z03yIoXxrcRet+1rlf8qVYiEX+2Ugw1MEqKVTGqISVY/pCPW6NB+nme23I
oJN7qH1suyIsa+T7uTDCOgJFqaCD0lorPuGoHdIbFe1VBloIEKkaltESjmMjp6iz
pHulhsD7Ys3htpiX2+bZHRCC8K8Tj/7no0npvXXU6/OyUEAddemGYGcR6WQRcJae
6GLSIIN8BgOlD7wC5vHZ0/Ei8HH3c7BU2w4nHCvpDAstHRwgOpaB618r2nNAN3gC
NDrZMmHlYOAjLlzrmbkuvqKlx7lT6modEp+egmbkSOvCQoIH6W9LtFU0AqvrAgw2
Y2Q19JeU9lk8/ptLkX/3r/eUQXa52Nsr6+OdiWEjT19c097dKtkw9sgpo4PunKaK
GeUVhmvL110m8SYnxIhRbg==
`protect END_PROTECTED
