`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gpt8ZmzOZkryY6mfmQpXLJ/UcUIlvGLQ8u9U8X+Gi8wFp3lKBELwrGHGo5LbiSIN
5Lctc32Kb1KH4KMAeLpTwH18BP36W9cOVc9vePcfRaQYdidSHE4Si3/aY/It2Rkh
6JEjMV004pufmBJkUffPBpCRqi0kJbU5ENPf6utf2gIRkSrhyRx7xe3PJsQINSzv
jSLEbJzS7GVrSdLuMP/13JnYWNMsk3o4m+M56kMLawDvtg+sh6Xw7sz0RB/imqNv
OpnIxP0i9QIiIqnZHYi+YugByau6GLERfoqVrYgr7OUCKBEWG5c+xuoBCSCgDtHC
NuO7B7NXxXvG5qv9gNBUPLytLswVCGsKCzLWMuAanj6ZXcgHIsi48bzfum/37feU
1ftK3D0MySsQp9zkHDQvjxxNfR/GpLNABNni+h50FwD5svC+fRNnXp6BPa5pmIfZ
vaDDVbHX0hmxx7KLVfchMH0e4HWMh1e15e12PaUk8j0FcJ5CiMMteRD/o3NLXRwF
LZfGc7zvDVIiR+5aPg2jEEuho5Bc7fhYCIj3rneCz/befOsL2wMpnQDxkV4dABbT
pXEAPUP7OiENq2K0YKbQclZ4Dtw6KLisnXC5IckA6rt03T28yALoNnrN5+yKy+PA
FyEA2mfhtCfRsObNSI1xqaxw2lZ2a9nsuJJuTZtjPDjROSELri3Fzcs6WhjPuUON
MyzpDElFp2/2CDcRwU6reqYyLPj2U+iIVVRoYdrFucPO37O6UHcJ8KqwwcKGrpfY
jSru6u6GT6OO0Tlkq+PrGiRZE0V6bMjtbc9yJoxbCp9EB6x98MPUHgBLDvekUPTj
ldYwR3pd/iDreO6oKVOKW86OOOvMtrJ6rFpo4aTL2CQZlkzi6+tbIqkq0HdFVVOs
gUwufBtGtkpjFgL7npMBg5bs3dBJd50bd58ZnWKeCQbYeoyWLmRq3u2UiVZC3gKM
3OB1GiAOxXEBmdpsF41ql0EhoTZdYxLurXfz9NP4sxI4fDMdFgh7dbw/+ciCl78s
wpja0mdEqEsg8xkFRpFwxYatxpJWcKx7bQVKCmGWhkHLVgV/Dttya8nikBQlLFcU
tReUEXxiMw1kd+2tRXouFReI1AgVlM2T2ORVAtQZmegfX4eZgEMc8dCB6eF08rv0
wTaqkW6gLiRFYh4EfrZNSezBRP7WEiXlRt6wS+k64vrzBHO8fGF81c/BRhsZYhUi
mrf2Xe4G1P7bb6TZBFz4erJgVaktqUIiY8c8bM9uZMAClURu9brCMC9Ko9T9Br6s
BjgcUJo+5es+RSoR47qduChcYzD+niV4xuzvp1kxwnNOartM2N52zn7I6+M/J1CG
rQnPeZFqsdLQSWCjy++iwXKN9ibR02jwsXnCqEJ0YbFlwPbD4viO4fJJ3tByzDuk
4MpD2BQbrGmlnHq3MQ9IdRo2NIEPfTNOj5ni5OuBmdKuDfusUxKon4rcNF+C7N0F
Cofyi79HCeZjcSpanVV8c0UydJHafz1fTg069o68zbvidD4dsIItdddG5HfYzm4l
g/wb2GWUvycFP7sYsPVGmmgyxHN84FWx4WRxXNXCqN0Dgfwjl5Pc7PNs0lO0qe/n
aGVCLTxFrPpc7PrMf2NHzrtbKq1V/zeyeuplYZmfrRqJux7yBWkaaunXQG1IB8Nn
jXQfj170V/o9Ts6DYb6xP86G+/VxKvLgSLI8dR4ubfGYgBc608NhLx7AzdKrH7gU
DXL8vep9DKNrXvQhbBuWi4vh6GL74UV/7+OdUBzaRsZ5cfocqVV5R+dLgEWUSP7V
Q2+kWhV1/Ykln8TYgoDP7Ad2SC+lyICUNZ35KVJcG0EGqrAOG1npfGW1/3786DG2
Eyik2HYSD90p9pdfTSQlDVFU4uUHF4ct9viunnSkumZRc3hq/ZC7Z0hdGsgXYF+x
e7ta08Tkds2306ORWFUPRnmpOAoIrOofd9nt4kNnYt6o1XO6raaeKenniCvi8BCK
77wAPqVC0sm2otXy1xmPRzBvZzmnIwmUHArFv+LwNWYf+Fs35IoIlsTBv0qkEmcI
jZSfCuZuNNexWsoBk+405QAYgUtH+fVG0VnZvavBGfgTILbCKvMntKox5eSS0jlj
AQXgGKqW3N749PB/I+cXJwpWfyC5RQLd1s82eyODxUAsFHigeYKAnW645sYKzPRl
FgVwblPy2T69zELFgT/qJYrxpzC3168XgyrNgyQxr8uMnWDkSr19pwuhzep5TJ0r
by69I7RMw/1kjA9NdtuuRvZErYTj9HDvmebQDrW2Q3/amAdZa9ojV9CwNidfoZLz
y/V5uvEM0VGoe4XLGOysenD3/wzUVFsWbZsR726OPvKA5/kyqOWQEB8pePImvMaa
ScrL6Lyp68bRRTexgaEkj4ujthlftdLH6oPVGdo1li41nvmcXr2tzxH7cJMk/JQa
aUk5yx4KRn58R9ClK05cVB59YozbarH2X+8c4z72H0NRkkVRWtN0Jiv15VwsbWJV
lbuUVziwMcSAEwwI2I+pZUpSokvJ0rnCVnXduofkHSMZN1XTaeGTCImYkK1jAV5m
ymwKDJE3LsKKF1KPIvDJKBh914EWy/YiHQ4pZVDu5iahsl9WeM3kAq3MQzriZGUQ
C2D5BqYZCdvi5+mDWAMnVEnc85cRxA4D0pg96f8Xu2aAwOjj3YoYRvDtJloGgcS3
`protect END_PROTECTED
