`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cHAHhl8tbT7wu/anWl/7PKNyVD0FUXc9LR+W2Eu+pVphwQZaPtnkdmV6XqKvaSMO
qOkoLGDmLBHHe5aNxIWiPEIc3kuD5tC5qXbo3dQLgoxKB62vi7K2Rz5Av4Y3vL6Y
+y4RcSu8/AfuNtr/SuduX4yNgWYjf5GSC4zzio8DgxkSbpy0z0+7E0v2gO4svUzp
6M4/xQTaaJM0VO48A6NTZ0q1aokXWfDIaDk8eMOeGzgibKgwDgOIfHvRODfmHxfl
6iQvR3zeSzNqguzZK8rA9Ov12on+X7Cj4PUZRNWt0eq7Tnp+1gk4ZpMMlk1+m2Wl
xGiuhedZI58vtRfDkvjlTjxNkcwhc6yNuXx//p9tfG/nPEe4NTaBMcWVMqPBewQc
ZwaCQErJQRSWIT3kT4oOrbmhm0gAifTOxhHkFoOX5G022lf1ZOqXsaF3Jct8pngT
`protect END_PROTECTED
