`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BwKXJKccjydXoM9XBioANJCBj3HmiFc5N6whOd+XjgJW5Y0GyyXeAFjA4wMfOS2D
p18HkPgyB/V3dk9/SdesnJfhXAWdbP0azuGvh1UlmDcC72gIBnLDo7MpYGCldUKi
XOxLrC3DkuzHyVaDx0J0ANbXUshREcBMmWW7Mr5iKJbOGW79U4geVyvdE3/+rVhZ
1WYIAAFx2VJCGZi4Vx+DpMJrqZjXHo+2sT+fkMhGi7uIvp+3ap3Plp2KMUE9NSJT
T4N01jl2TdWIpqbakSTBtSZIQNEHG4AW/edrJPXUvdCY086YuwX9mLpiq08y9cAI
DEbmiEvEpxtKnrnpPRnq8RAPZrWAqVksy027ia69o4mKKBR0AZHb7L9e+qO5aL88
WCeCxlB1wuwTQMpaX4A/GjI9YGk4Izf376BRR1FCqNjSOJprYXhK4nLBIBOle6gI
AuKoL9b8uSCqEI1YHL6iokFv3XcOhyROywCOF+Gx4iqj7ZvIca2S4e5IKn+O6Hn9
e0KPQUQ87fdx/xJbzsUBRZr7c4wyJ1R6R8vQpMY1EII7WsjfuH5S4DxrRT1NRiHX
rwH7AzCMTQn5vJpllrfNe5J1Uf0uVBOP/W9koE+ASDYA6nR9e/qKgNhbFKLAkB2t
`protect END_PROTECTED
