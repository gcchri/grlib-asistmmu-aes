`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HtFxmwpS9NfRZFt6lDUJxOH1g2hrqbsTtIn4P2xWg/5TaJEEWDUwsGpDDylkVqcB
ySBS+6VFhrs6l0Z38pOYZkjUEQdf+TH8j8SadXP/sxY334nPpDJ/qFsFRTe+o9fm
qWiCe/Bm2Re7c943Ix+a9NibBJ9PMw64AzZ+QC/oyFnEVlKws9rnqyJi1OsQevar
LYmK/yDaxZK+jBOzmdbcvDc16GZHrTG6d9IE7V9v+vW7oHIVIH+qIm2Q4VlLGLM5
ZbP02jWJ1ceKpEmEkH95BxlT/p5b55ZtQfZJt022NQsNq+J39G8CRRz91KSuUfSe
TMfEji5JGJuhK2SeD5RyBSkUoSNtyEghR2p/1GbODA6P43Is9F6hIGhMxOug5Gdp
H8MadfVhxf1oJJOdSsie+A==
`protect END_PROTECTED
