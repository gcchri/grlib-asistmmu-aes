`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gB8pX6pymHBtS3VGL2oeO1hy6nqxZ1vZjNfB9DRCSGpJmyBYRRN+ysdq0QNWdHH
mq5XxL1bl6Qc8DKiZHUqTvpD4QrqEzei+9TFVRouQ2Hr7wA3wqd3QWjD1+6Gnpbu
pP857DTsPp24zkdlQn1opGLBITV+q2oeLyO/rK0iTzXf1rfk8UG+hnwdUfHn74sK
9TnSqAh4wFTKRGR4RlGk+hPoYUijxxn7rCDEmUo/ez2f+gTQLtocas/1hwfACKnB
tCKrKPR6NSwAkumK9PvUxIiOSn6t2rD6owTDpKntm6F8XOhYbxV0rA9zmNe4kKKK
/313A7/UcJ/z0Ji9igTyAyGPiX57pyQlQVxumKN+BGzbCkmFwUt0a281aFpKiuLJ
JFjqsipYtdEc6qO2h11+7mi6ZzTP/6AWrAYCow360ar6Fcv4YM8dqRx1Zgqh3AN0
96DO4Z0uyTFft6iMXzmbn1rkZoYlo8zTuRKE9TQj8x1XoP39qa6ecEr8nAkaQDZ0
6ZSNgygE550bYUfZulnhwIP9baXLWCxjDLRafKb3rCfFKju7QQ96/jkmBMmcYfVR
rlNFvCULJxzjY8Cv+nBzya72ju6AQ4UvcoLNj+GtFVB87MU4gWNz3lxeVfX8okCA
0uR5Z6dsgIBxTeWy6NvazE8w2oYzOYzIoRVmMfWg69dMlfvGSFOtec8C1QgA2cAH
MxwJ0Gi1Qs2s8WUMa98wumgBA9cewo23HSObaKS/hSKVfy4dIqN9Xil/Ejj1bGbS
igy/k2zT4QgdG++yx8nTGyphwgvvp3xE6CuwReBlAxVN5inXLKNhGHlfEJyhakz9
WCHmTSR9FwZpKPQ0E8gX663ZXPbQU7DLyim05PsdbuCAJacLFSWEQ9VVBFlzaTCm
pVSjU7RL1z/m0XE6jzqV9jN9Ej8zCxmFXRVmcvOpM+4T4kKHZUkvqIfCHcd8vyxJ
P+MJPEabnZtmoWN20tUBaw==
`protect END_PROTECTED
