`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWmARLo6KTrdNLh+ksMzpRrIlPjQMP+ojfc3iLO/QgaR1wGAlp+tEmhfnPj1qmxj
evZpyqJUDnAASAUwH8/PGLKcXLYfLRrlsNXGj1ux9jgOeyIxGIMJ6wlkgD3L2PJ0
evyC8dCIHlJW28r7jyD9S4MigSeHUV2kWRWDFZVI6fu/jKZoiSGKiC1ncH7lIs+q
fndy4vIjGZbXV1ZBy20z4cZcRYQ7ASQcHL3j+sbsYxFulxiTOxwlByB7PJDIyPzn
up+x9qYV4XUkAjy0voktKe0Sm82l2OhIJwE6dA4cwyv7bueusSfJZBKc2ySbbb3u
zqgQvfR9k/UjfHS9Q3FJf+s8d+Bctsg8yks58Vs2/O3+BX/g8EFyCqHBQwQ6Pryg
7waJukKIHV1k/EYpH+vWZZdssTbACJRpDI/HmQCSDJdSdxGzbr600iL725+f/o2l
W0boAFuOfGLPsBChhYBsPpIO8Ew+kStJftapULiarishB9ZEtx1nfsaDwZEW2YPI
7Cgp1qQLOF6QlUyBW7Ed3GOBeNDiOHVCGZkL/lpKSKfYjyuiO5lpvOkWv5kz1mbN
NGG6bRt4GIPjppFuyBBxrT59P+lwMpPvxQpp+O6Tj9A9PAuBaPNWOAjdxb866a5s
EgKsKXxJlCjvr63Z8FLt9FP+bGOBf3gG85ZZ9fwIMvdYy/bjiZTNFkuGo4kr7SQx
N9pXWvqbgmsYJ5sNetNra8Vw2ggTYFhyNYC5hezncMCmPX1qmkZ7WmQkMZQK+Lgp
dFhQhInB6FIkCeNsYxpGrD/hejNI9VZ9DXif6mtwSLva2gtyZ2NHFrE1nTLOL30M
jvK0miyYK6q2JKOSMe0N+0+GUftDfb9muHP9YHKuT35uxSM8CpAv/s0GopUEQIOf
aU1vazxV8i6M/WfTyq5wkqcsidFQB8ofx5aSvK933/wcYtSFeTnmp+/QVYGZli/R
hXp+o1K/A/pXL52MLnXIr1lX4VyfGkwsl68/gQ7Wc+N+Lg7WZ6SGMrROYjdK0RRg
csv2mitO/vMJBHyUoHfDDq4CpBoNxoDExrTqQQ/Ll1Z36EOrtlZJfyELvq0guI4t
a/4mZLAsv2l/jjx0W+7uV5tADzoa9xXTp7dgms2GHkSM1lpy08In5jn3GKV8ETmM
IPSLBOZsaKQYyyifoblvWghneHzvBX53HSnMB/xqNwZsYSnSa1gqXcJf1ZPfXEyf
keheTUY5Uw4f1feTklw4Jm5jsIRVGrXeTO0KvIH05f9w18n7ZEop/T3ko48iv19r
qqLCQvcnV8kw7C95xjWfN2eB+VpirmUqNmBQtM9W5FJ4/0USQwqxO8jcTTiXY54O
oCNHXxkjr3owXlZfMAXWGWnytlkaHk5ScVNemqXu3S6fdft89wofzfHcyDlArqN4
Xn7HZsYVmMOLioG+kcV9Bo5stP4jS1hBgz+eIAHF3WcP7a2S2MBRQXDbA0B6lycR
SkDc+iVypIHEy5eRZ084yla37h4OXUiSVGFUJqvbgTA=
`protect END_PROTECTED
