`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bRIjZv4hb55Szfo6cQ0K7aduZTnNeiKJ3z5s1lu0XWhgJQ4cJPZlCb8EkjJU5kW7
AYTw2pTNlPTzJKTsWktdW7kVFNhJGP7qr0mjG+y7fxewqk6z3N7AeT3hGjIUVLBw
hlyCawvgk6J6og37GLQMzj2Bb3HmV7j6yu6CI++qN2SFz11ROl0UmdIPbEFdpvdY
I7KFo0PKiPS1fQeV1rGsYu8xVtIeIxi8bbZUaPRNo9ckm79KcyCFZMrd/orfDch3
8Q8Tv+35kO0+Zg/cbzmP6/VQehyARfmfsBYZMR2JZTC5tlP/Y5Gi6xoaN8OW4rvK
rlMvcHmitXpceuQfTuZZZurz7jyv82oNarzwlx5PIlXhcbZGLjE0DDiSxPm5eRdQ
6QKU/Ett26q0gqDn7Wv+FMCjmbGx5+EgL2CzyMyAM5K3XsbAjo4crUYOF3aHNvyJ
8utfZOeR2qswEy5qTc3brx0YPhL8zUbEikJR9LjX3ix0voQELQ18b/FQn1Hh0zY4
`protect END_PROTECTED
