`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y24xoYw3oJG8HLl8Wq3U7ddcNWBSigwK8KNqS6lOrrx39yG/0bWZrOjd+p/oRJ0W
bu7UFHLkyjf7wkuKXKGrQ/c0VzIKRYMjagqO8TKEVancORbhCuv+DlTd9xktfuAg
zdw4ZUf9V6tTSHS6ShWF+uTCoSpKbuvYWMEfFqf9zTV1Tc3HSzQ+NnsWXIK0O/T3
pEcNoK0i7rt8gKjHftbk6wKuTreEC5bBraVnZZ/kb2jRx0gJU9IAqE9MGB37gxaj
qXn9NktX8Lb8i9X26eBuhT32YRnlIB/0HhxMATHTGlDJUQYoBcWlExbNr3JvAhUa
kA0fdN/FL4TFh13Crz9ICHa/Dh9VOKQFqYEJuXI/S9fSQZlfJjJFACkk6x/xecW/
LjpzDjVPlz5vRJFEueSG7Q9NSIbYqUBNhu7v2A80Jpuoa7q/s4vcPchJCKnRHRvN
oDQAyneYTKWYsnlBPhkMEMfmogFiXg7StsHH+xW4BOECXcjQRIDV9Bg4COkNDaXR
`protect END_PROTECTED
