`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GUFyqCxVewVWBxBplSwvw8Vjl8GZNmayGJR+LYzEbWhraJCUrDKMFyI8S2xduzX7
7bQeq9tjX3iLy5o7D5OEQC5jubGUMZFyd8NQslXumVN/nHbrQa8fV9W9rijv8QMK
sLDcyFWIAx3DItkG7FIQ9o+kFIu9/ebIPKfS4pGqCwsFelRxvZKg5BYanYHj9jI/
UpefzpXvOIcPzLyf3l2MtaH9sB6/qKokeXz56M5MV1UoeT7eW5I6WX7FjnZ8h3aM
qByUEBdXng+WwmFFcu4oZ3KXvbxrBTeu/TfO8V6IyG8BgVglFE0ayj2lTh6lenGN
ujpi+88bbdn5NfCSFJSesA==
`protect END_PROTECTED
