`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+kGKv2E1nXqCRemOSiY3VIrou44iO2krCzVjPkCvFUlb8fEcx1ehJCpxWuHv4P4V
3i3x+O2uFqvmCFA1WRzGijkKaPE06UZFTL2ucvRyvDNZmaT7lBe/YTvHiwz3uj+E
Jq39eb6wPhveF30WZ8smpmCShFzei+dljsFeL3Fx8rPPx+GGgX54p/NwAz1D/QmQ
u3vJH3o812yfVqBkSdjhlLCq5ZkW3DZJz+wTMtAm+A2kvly5S+A7novgFxxCiQBO
wCJCjkUgyMfU6lUjy5issW1KeuoMnB0QnMaWZvv21ZCLu8CquS71HT8fn/v4HlLI
LlF6SD438F6Qy1bISofj9gXomsDMRaJ8Fnqc+prdj3Fao+7sHUt8N8nU7ussznEJ
2ozoJa+1M7h+oQtT3e0wTsd3PRJq2LX+U9pxSzz/09zxVlQTMalqZaY+f6WKMJEJ
UssSlo3iFoTbIfGDnZ039gvaN+GzB99fv/lh8quVaRAFtJBxZfpe9lnk+IK8KsLY
OjeMkVYnmvBH4853Ndrb3czv3Cp0qk5+8Ci1ebp0JgJiD+p1lvVbjqfxwI2vxuUU
iFUG3Mi2P8UgPZMOlRVdggAI3pLqnTChlGZDDxecJMbl2N6w259u+PwHH1UYNvYd
9vZYInJd9Fbbg9O6tfYXPblkiFEhc3GrcdLHjYCHh3BGQSqFidHJ7EcGljpRQuHq
19y8YgGwQP4DT7LWdvAeFVa6daEaFwdGJ2eDlk8plnXkzRMsTNWFiB2WYwDy6bDS
VkNIBtFUgi1NuSR1iPwhIeO8BGBiwyvsAAc2eRovvIBrwYcuTl7ZMbHVZFGEW/DK
BvXjUw8jOjJ8xqOzMLkatZWvWCJ9wwrS5ypGzHpoMAeUFEHXVufdh7TI89bHJuXi
maJVFd7C1yP+RGFHt6Y29uIwj9tCgOoQ8tfD+rYBlLVaAW+xJc+VR9z0agbqlAvn
P4mBiuHJNi2BGW/YTEwU/CwQqB863al/T1bJbQWLsLoH46mqH4NkNZQmGfx8E60y
a++gCoGr1SK+5GV1bPRaEy7tsW4eqDm8I3btnblIPKkUTH8JLn31F0SWKr7RS5qx
ew9t/iaH9CB1gklgl0yQRJoBFjlmqxPJHsJSTUV977lKspjQ2FMdPhiKkIZhEqif
RDXy7JCVYpinmWnE6QW8gvr0qxNlQrch1iBL7TXeO9nsMf9YoijL8o80XrU5PLBd
`protect END_PROTECTED
