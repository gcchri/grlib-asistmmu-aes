`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/zX9loR9U5zfvgTaKt+nI9o6EncgRffxJXoSAEfLrgaEMAU8RMnDLeNa54ywUsF
tn2tBhtVy2vVjnpuZ/9nkEX/m6Ft4na/WLDy7qcnOlyCxA7VoBfVwSIPL/xJlx2C
Xcy4hYbhCjvahobH/wQLXZYc4zFudkqGT7YBkuKD4IESfxJyuVyhNZ4Sm8yZuMU2
0EBbPQylnhh63SbH0BxV96w2o8Wf/CfLRTvBlWXQxPvu4VfZwJF1NGtNw2LVntjJ
vRsOFDDgar2RZNh0MWv7U6g10+GMhdvvG96N/GiSVGM3w+jxIUZm2UIDhdOLrcUJ
minqTwJMUQbtsWRFtVECTPrrXqXLPzTZE+YBZUhL4aoHmp5fGD50YyNI9/8FmKEG
`protect END_PROTECTED
