`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rp9T7jhaGjYXW7LSY+m0TYcGU4x4K671JoOlzVBm2WUGhMYVoYxPxt11rMrnU4HH
dFfiIDXP+aeQwTJTh/rXtTf80pXXYX5a93XqokvvTITsqQ+hZaBueGyY71tz7qNo
cLGWIwfooGC/GGNE59DluXnfCfsMWLrvZKksI+bt0woNeqWAaqZPzgJcWpM5Vv4/
HKtbRCL/4e0vgQpnZOUkMCZhBI7wKS0muV2MreGpy+y70nyvsCevEc99TYhUlXkS
TX1dgSrvOIYdKjQRnkNGIBBygYHm0pC6qW8i4dKcezA9B6GnBzhjywH+SWY1V7kF
UWjS7HouZvR06GDGwZSfnUH3anVMnivUwUgR+mmQMWmp1EOv1iq9gJxk56IiGKql
hfImmCAo4rs870XF1lsFcwvS1llVRI78QHhzS1CUw3nh3z9UXFwN1Y3vifGIrZ0D
e5WVM+r7+F0Dl4A0XTiiU7+Pw8O1zy/C9w/1q6dbt06WNN62yv2QPFMQf/vqqvEX
jSFvw9fUUPeZp6uhZ1r2qfHym+SeeTWi2sdGbOBNbpyXUMyJ5CDOQmCQAkDVRKtq
`protect END_PROTECTED
