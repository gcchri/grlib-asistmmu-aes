`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cd9V/yduw+CtqIBQU7PTWh0sHKidfrwGC6y+00aYeehL/7v00mXFgsASYdt+e9Wh
79UMEmep7B08OqvlCGY9eDLXy+dcbxXRCF8X6LXs29H6pfPDMGAkt8XjT+F71KJs
WPZVU/8fGIS4Dt/we/FOWAIUoZ0paDEXvZsCgtB2Q4ZYcH1hfzk6MqvOc6Z6rq1N
wXk6XfCqKh4egtoPS2thSXfDS+mcZ/WpM79XpYUqoADiLSsEqma98DTEz/0y8hBS
3f4ESrVqK0XWHBMKiauYTPqBJYk10snIPDLlPC76dB4kc9YUi30Yj8WzbMzMXD1e
9DRj8g206BWGVJP7r7+2APOnHY7mO8THlHOvaTVBTsP0locC423XIJFnHU99ksuf
L1AspSkP/OY7MfuuFJM/qkw14rIEiYrjvMlr8vL46dIqM0juynVoN1yuZfebClnx
GYZFV5jmQ+CUprwJzaOKM/ru0jaitToDUTxwE7dLJkFzQw+4KEDVw8kBNANHknHQ
8TdDEQIo9gzm/HcqgGLqu40xisoJdmCqrU6JNmYEV/wFgS8U3wpAU9fyDyOj3QrG
t5l8e25OuBRifwrZUTs/UWwgx2Psc4/XzfnayhGeE8vbOiEzd2XDQeL5FuG9YJ/3
`protect END_PROTECTED
