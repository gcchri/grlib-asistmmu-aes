`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7tbDUNIzWsUsb7pRgQMqUKPl7W49tFytlUpT9J8LXGLDE4o7889g0gwGkzO3t45W
X5mHAME1mDaG9oyMCsGTVHTBfxXiGA5j+Onxo+hM0oEO1pfEcnVP7O2LeoJHsybt
TIpSUhB6+sZoEDz8qF63/Fg4/CPTP+dsNSkpGt8mZP2sMNmr+wD43pdorRUlcKt+
4D9IMn7Thkwb61js73++5QbSJt+ftYm9A9bIsDa5axQoLerX/QC7Clh4UHkakNDX
PXWsIBnyozVABbQPiyNSTILh2ztRXNNaX2WgZ/aRrBiZvOOYnn0cJEwqOekIN2ik
/UGrIoFnkDsVBHjnelKI4hSrKXv4zyaWy3wCU4NwsWOsRq88wKBmQXXEbLMhnVjG
q1AnR17vLPq3+0fvPEswwVgVpc5ry1K6rwFIcC3DgpNT0/zyhq78LXjje1CDKFC+
KHJFFERabCe7apsRh0WJX56NA6yP1jIEzb8pYT8OkCCUPIHm69djK6gC0uTOmgZs
IM8iQZEW67cPYz81gLmQ6g==
`protect END_PROTECTED
