`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24ZRnuVy2GGc8nRBUTlDKmF+7Hatky97xNSJzBrh09qHFkBjZnJxLfCotg3vUq8V
9ZL1vinLf+cJUNs1R2S+p5Xv4DyMDlBfC3RSbkTSsRCAu2QVvx047P+1dRQD35Gl
Pw9YhKGTD49+7eO3qKSdYsrz3NIsFe58ZvC5PtxHq0LzCL67OZ8WaM2BZJkf8Aqe
q+5UV+FUpSJVH4JI3lgsWlTCwLteXFHzsxHVuce+RU/xE/jr/CjATLRlxgmkszS6
0aECqW4mDN2CHhqJgTi1GvHj0CnAd42x/xICQlII0JIxVXXd2X9ipjpBWi3pfy+K
gWGggmN9xo1ak9C4SV3MZwfJIf2jNVHo51KdUrhvhzRrtumSw7vWlJ4e3yGsz5cn
Q2xQkZ2uie+eU4xmk833UJ8AqPxybYtgtU3kcGSXCYLekVzpKfxPxuBXyBEnC1vK
C8X/O6ATy3GBxXrWn6XTg+Ddq+eLAOyxIlTmMJan0kmKI1NlysFSZLqkBCli7xB7
bttqETnOv70qSy+HSxuMdljG8LbnTVMStWZl2PjQwwA=
`protect END_PROTECTED
