`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DmfrA2gy5Q8jtA5zreXR37+sUQRohLRQL1khGhGMxaMY/g8X26FN0vOiW3J2ZWUK
3jL1SAZM+tSXtPrwozcgzmUB9ebFwYwaiGHnVggU2NMckwalzMy0yJKGsk42/Ps7
UsNDNWkWFVCBxiKpYAOJF8NWU1SNxwOpRnsFWqkJKpH/hZkZoejfmkbdUvkIJsUm
m7nJBNhvbpEdvNfzford6R0UiRS1vpnuco9x2FY0hIG2gGYb83OM/kwXm1hduv1j
EeCinfNbweCA5w0cbnOsh05FeedNYY98iv9tFlVmOZJI6O4HluxiSbiR2mJv3d9J
Y8//R8QJOStc0ZG9rT6ceMZuZX/z8vxkdYJ+0K3hkn0OhqxUDmAG+sE0cy2AwxAA
ASScR0ZyNwZ2e0va3DHvx/So4x7zAVnoGf5rtJh3ywnsUNbSn+2e1gzAl2Kon7QN
3Ryly7RJYXQ49SkTspvls2xVd5csPDucbP+ongaRPRrlynVF/E/IMK7d5Rl8FVIY
hlpl1KQL40L4alVu5bi+xgya6B6ZusTkRxvqtjgvraxC4aQOS3bBqIiLnpxJe+Dr
7xzqQqKc5M1v7qrMMlzOUcWWOLxkepYBPACw0DOnmEGNISY6Qt70AlT55TwqUpH2
JLB0fRtVEI/Aad5KW0M+5Tlep57WuxbjfxT5kGrwH1vwRlJcYqBx66HQiqGrxq0C
KbMs3jilLf5qXF4PkNQ0bw==
`protect END_PROTECTED
