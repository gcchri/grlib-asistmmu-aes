`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5NFDl4G0mZFY5VTpyR9QKvtJmmuyMeMoLxfq4No+6tDchuyiB43ik4r2FfNImlE2
sfBwwWDC7olHHqAX52NtTuU3lRUccIlnkgqXne0ArlI2YdQpPUuTIFv8os3gMNf8
jergTuPLxXtl56G625Dvm1CLkeSVFK2VZXvfrUp1ATXq2JBxmY63zEGJh6CBmYtT
FjxyX2x7Kkw8IYNDvOG0VMbGTTklbZzgvqTD60crPCt4cYjJKS2MdkrP7hNfLwUV
0qt3os2LwwVqoPhw5P+e+xCq0KRQnopk70xhy7rGWq7arVd28ZFoH6FBQ5PvIrMY
lI5RcsZYqkKxy2ZmkkcOMybA/ZkkZ6t2eOQMAgy35x6Kpt6qWi4UxQtbPPXnDfGY
BB2Dslr+UlQkl/lxn9nuVS17PlkU6aa9TOH/Qrp+uuGEu7VRKFidILjtoU7haBJN
`protect END_PROTECTED
