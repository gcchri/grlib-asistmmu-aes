`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ji+8/pQlXQbGi1sqDK9Q1hg7oU65rXeiSv6Kk85r4MqiGp9vRjj6TRWWdPMWgN9P
Cp7llM8VK9yvCQ/7vJuehoc72r4N5OibtpqTBHqiH6k1RS1WdYVkvjn3yy6Gy230
RAv7uq2X5+NUbcduNL37m4vBtj8SKJkOzmg0j2k0Yv3V1/xnJmQPr+hrl8RP3h7w
V0DzaYeoT1aV0/jdNdqaZHOAieKTgzYcHmgsmFVjPaREs/Fjfi+Dj6JgTMKrdCAm
OYyIMOhKOOpgofLEmJ1ipevbKIQH5W7G/DYNbBcFw4EV5xEnsH9pwnVlDeSbB9oN
9jF3BUSmewlhzUIUsaj/CzDCX0TabGFPzx9FI7odpnMe4aLE+Y3SzTgVPxaocwpy
XA66Cd6MKFowxOMFpVPFxQZoNLELwlo8qQy8P2bK73AtRSyJSAOeikGWv1iIrOA3
fJ7tTJw2K3i6aRpTWQnuLQU4aiK2kk1ouNafUJ0PFmf7fV/7mju39Z4bLngtS+Bf
aXRNRAKGtvyj5sn3ewGfoSk9tfTSgNmlM/X9sTbbFhvt8wqLV8dUr8Tspf+dLhL0
Xrkjztb/VpAgrv0Nanb1mg/Mq0XeRZwOLBfK/YHRVW5YzSDmlYoiqb7wqV+DLCvL
m8ZkHAjkodWnQ7Bu7sVuRkyRRVk4iMkE3hDy0fuoi63qR3dGlqM+Fd2WXJchYAGQ
xuXVpXH3MhE8zhOLxHd9SoBQQb0OeWCORxGmW5chWLnnpQkqSDrLEaagMSTc+V81
a0meyWW0/1UOWcra2S6D7zQBGTExJvWaQ+mESNjFKGoVgkQb1c4ycnD9nHs2hUER
TqrsSOQ2d3Hh56DbNl8jrJiRj9UKQw3j4Z9sQ7M6A09FoF2SLUZzg47JO71U1A0e
7+QkinP+Cy1rdqpi8mEV34X29i1wepTMzJEB34rgJ2sySbnriq8Ko51u+kBsi5Cf
ZJ6zA275J2dhgXirZN2lA6WmLwdCH/mufE6bsegic2MWMo2Xv18+qJRBXS4SNEUm
t/ByY7V5G90zRhhzI316K9az1RMLF8VQxRnH9GUVD1wpFywsTEKamVOrOAEz67pB
WtQDH81smG9b16cXShNt66eMIQNGmgKwS76b3yjZRf3B0lrv94cu0dQQ8E9CoUgl
1kLSgUGxXmZ3iwB5q9WzWRbSwEPuI5fJs+Y4CKfbmk7+bj6VJG+El3t9tVlHCmrh
sZphzxeu+jee+bQT60gLOGzcIk33JmJvtynabO1RLwXCPOvBcecIKdQALyDsNzE4
1bedYhVIVdibY8MlTC1rDOJFdJeHQJGEGNNvfDMeaWSWPiKq9MUsZovQZ4KKTpXB
eeQdUzmQPClQSoqwtdxcIAJpgZMDjxv8BZqDCRT88iydeCQ5UL9azsoY5QPu2WeG
U5B77aBbo8znQc0RSXyNeh1GJ9kzoDhoouiBJxkY1L6EbHqIbMe4Hhv8akqBXJ1p
4rRlv5jt0nCrzEf6fWFPZf5qWwrk0xx4LPUPWD06hNFmVoVJ2qocIQllqS+dPLcQ
MD73fqilwJdMJy94t1WGYCvwUmQLTTCop2w6ejNdvsX7eIxsQS2ZlXIYJ3m44dsL
0U6J4jOata7x8q/Qjrp1XvMhw/WOk1fRbeVQGCvawm09EUUIQMTboaLq/fTSc1Ge
meyqxUkYa1augxHdKvanE8l+sBhhwEa7YJ9xu79ZUJR0eJj5pLzKf3XNIaPVQkNJ
mCFqH2bzvhE5Pd/sGjsDmEaP+haXB4VkTyz5YAAaOKdVmlJHHTHrrBYyHVW9VLAG
qKkF5pEq0WUbIFOvIct6kGTUsyWMxQME+MOi59Ll6wkO7S5aZ3GQiWp3m0zdokxD
BkTYUE+yrCK/KUZwxU7fFuHQuiKkTs1UR4wiaHR4VEN77wLb2L51RjK0VGe9T/r9
oKbIE7x7ljplGvw8WgBPfc1tv8k1jGyFh3jxzFCuFzEHoXexnAicziTO+hUBZHVO
0QmO/P3YqE8rlnCmoc6NXrziHXWKLpFCJe+m0aWfuB9UKLfYQfrJDaYKDMF2Dy1X
Tj7tc0EE5MvZ27lvS2g0cA5IWPkr0gKj+LM8+fOP/h2w9KGZnxbSwixrPbx0gOAI
GK9z0FeiP0qy+bH/zyJ0PKn61CH9oE+4y7Hyotf1VtEhmqdKk4o+YsvNlg2y/WIm
gdhb7scBFAUYNFLVsgXUiCf9sUaU3aF7Z++f+1/0j5sZ2FjSAvmKKMMidG/wNQ20
aDL+Ly13UfsWEcUBIB5MGhLrnMIv3nEQbowKLkxJ8c6p3OtvxeZpN0gWB36oQQ/B
Ve33XjPqnj+ERs+Y82DjWvflpvYllerPvH2A+otpsDw098ezZAa7sLw9Wuyin/hH
Noy5PxzTpfvvLjSRKci0BBntV0E+ovYDai1YykTav644GE9MRUUcABoppwnK5hXi
FGf3pgdx3zAhI4l+CqPdX0XmcRYlNq5fmRBtmiQZ57um5zJi5JdfzgkC+2VQhAyO
z3f4bV8Gxk809SC9QQcs/E7/kbDE33LTtFPXUkXA3sGZ1vDFS+JkrTXgHYKAGSL2
HNvUr4dOTSr+V1GS8jYQ+7Px8MnSMVgtpUAsfkdKon1h2PgLznsA1lKrRiFCWVV/
x1uwN2Rrr0ynS2YKiiRJenruMag9fTu8C0ia/T0mhDNwdYWPToAVoDlnDa7QqSNl
2MbfvDdS0zw28GTqF+m8dfPj616SztBW+zkxJiDTkRH+BM32m7dscKdP+FGPE5xg
2SPOv2E85wzm/wUb4fBHwqbQOVUzNe3Ob8aRQNtYeo1Dyc9XTJ6iechkxxkEEa3m
36KfE5TeCtE94ROtJqgMJjs+lduQENw74Z7tQp8sibFlyeXF6gRSrAae65bjNbdw
eSg5GVIMlYSBZWofqwHDRph0hT8Sn+5fGMypKVnw3mbyFuXlCciAbwLtRMItWM4R
nr67jc+vpGQmB2dUbbWszh1Wl5hhAd7ONrt/TSpgORn+cbNfNultcuhLig80b4nt
W3OAbh3u3eHCoRANIw+WeREZFXTva7Zox7zaCiFTNa4bhGSwt0prkQofZXaSwkMx
nQitTZJiXSxToPr1jN2DN8Nwa4Z55j3wflPhUkzMvTspYLQWUp2riVmLshmfkqzu
7dJMzl5UBdjSioMPJEZsv05InlyuyjO448xV/yWs7Ri14RhGp6NXKJAMxKIC+Smd
fhZDkZzQmAY/c5MOLcfPXMzPDU06j0FFDFZl+w6hoQkb1zuKCS7u20fDjklhl1IB
nMt1PuztNzujFa0xuTxDa5Dp8uWZ22r4eD409EB05kooXKj+N5JPw6IWht69U2Kz
8casIxPglNhkgZpBgXKdcAmaTHoMF2TXxTIzL+c5e/SfJhCdtzl5MwxInqguW+rX
Ot5HsQWnCcCJ5/PC38pIqew6XE5bNon2diP3FaanMGzTE9Svxwzmbvn8Qh9JITEr
efdmcYGbibdGqdc83ADXqkxz9fyon3B+PgduDEe+1LfXtCqWJmaawpKy69zGY04u
DpEMC/0/X5VQHQqThtOUq5ySOpVuLa+EU83ioiYLZa2N3BtME/qEleSpNiilmd1g
8h6YPSZzMHGojlUwQyv0c3ITyUae+JeQ3bBncNTn++6Fo8yRz9tvy2CTMZWZnyCq
v011DyJf98/33gjhzgBfZ9OUDoyvQEbR6k4LES8yQuQtnRUtd8IFZvC40VgJkU4c
gEW6dLz8XYYPHhmHg9id9W00Y5jMHqY27ytd1EdzQbv5okwwcLGhH1o1pKFpD+5S
xPl8hUeTTS41uRrYfcyXHvSmGV6PUV8v394eAcEh78+Rpn1CrZ3Du97kwZbOwrig
wcC5dZnOPrFroGREyrPunNxKAaH7mRnyalMMMRDHpjD3UUWZzADdnRQK2x/6r9J8
uOS0IFgIDeGdYH3h+kY6+W0mza/gU6QpZ209ex1MN1ggLf8zhasoN5YBYWab9d/1
j2XSt0gFixCd5ZB2aVhzeXfCwr245Mok1g2tgPzNOgcyt3FaAvjsU+zTAfUe98OA
Cjzy+vLIkZtQpRHKMO/7iVxDUvVVQhk5vXmy6nRGZzPC0HcGsc9BOlgt2QCw9Bm/
0ixMr1bOIXhTRGrCTMks41iAwkBYNrRnFZX6x7oKvG6fFf9E0/BdHQfnSAgzaBDB
ZBO5JzHxxZYCGyYg3Vwvt9mqbUMsJOx3/JASTI1WAWzzYRlr9xB9HFPGvzJ1N6TH
cKn7mfv/9HTxpp/XPH+8sDHfxl59LIkkVYlEMJ8lQPEsiK9nNsY+poS9sVEiefCo
yr28nPGDjLE8hsO+o/+9jUUG/sbmz5G32OrJGbZqjqEtDz9ospMbLMPw8ah51ID2
KXsJnklDg4sIPnIW06PvrIx8bXsad/v1yZ+tP/we7mLfwAYyKezFW6YcHqydsHQe
Yy+lM+zfWJwSXw8p5Y617j8JG74aCG+WDYfzX3lFq/AkiCxHwq2qWnsWqHYiZi0T
hI7ppjF9cZOOysyTToq/72ySz5m3QCbvhetSBfV0ElMP6e7nNFxHktN5Fqn29Rww
+eNyQQji0msR7bsj54R4YUkFKEYP9NiszOHwIhwXF1G836ECee4ObMc6G1oV7Brg
7wCrCTGfGZ1PnB82Z5T48fg6R1fcu0sjHD2H7xrDmR86Jz++u3BWrjcPeoet/wtA
teTNAqF01/ych6HWo+jzhNgJLt0tj3hzeVkGwutmb5BYFtZqC+vyvAa+ZG8QQ9du
/RbIgZnE5VCWjPSA8TE+AJaSnZoIqcfOpUBldlU6GKobkAD+CCSzNRFOoft7KBSa
05K6algSFWV8eMOMoUj2rbrjYrZPVRG4HhQb7AoFEHTqt9Zw6MXp7ETwDOEavb9u
vK+vuCB2QZVZz7eNv2KKZ2VAnBt5VW/ALaB21zWQqEqxTpzfVDIvnvBq9k+YQiZ6
zaNMK4RlcuCvQmx8Ek6crku5W9Fv5dg5yiSdwaqRXQ03obOuFm90wNy+DiKCleZo
v6q6eEfMP6p0/gPIwUwq3TPVILJMdTjUP6bFvmRCHXUkAOdVRU6yOmH4Pv1GfUri
LmYUuj2Z+hMHMXZZ0vhNm1G7nQThqTeDjnMcQP3HKfCt3iqjf2T6nki+rKwYM+cx
oJ+hIZAn5r08zJgs824GF1tF5JRhiE7jO/9Nh2WocqNVXy5+0x5We6D5uxaT9klq
gELLWJLfrZ9LnZ8FPvhEYLsTRARpyw1RliesTqWM50QGOFDPWyf+SDyC0wbPbt3O
+ZmH7hY3rrTvpo8R2lF0h9HLJ25ZwTks388h0YW380Lttx5P4sN8q6PB32L+qYIf
wMeXJ3e4FMTqqrhO4jnrjrY69AedBlNUb6j8yETeyXdkapPh7voHEaefnbw2/Gt+
958GZBAGHtddjEeBPq1kvzR43DYI1YQbKpGanmcc1J8hOkC/1ycgxePUQWwlGwRM
cHF85e6UqJlDEngonSDp5WoTWCjZjzOIc2a21m/ASSoTDnOQYbTGOBkCSl1X3vIP
dMGHkHdM+Ck0hl3hv8lSRXsnxhbPcqJLPuNWRYSU/DpnATgLm+EkRdX2ifUxVyhh
8gs+6kmYUuUGN/NaX5EDQxYJWr+gCdcvGWdsgjH8QEzc6gEH7k2J/cUbn16jazhh
oHQlwkYvHZRqkkTu3GLURiYLSQnBGZ8v9M0/Zhmpo1Yy4An34SzdcRQHVGgm0y3X
vGO/4Vfex4shD2/nBxYY749e+UsbBQ96bjDE6o0Ul1WcFMiwFEg4YfEERc3U43wo
xxlteI+19BDhQYH60eOSIJsNCakzCy1E9CXXxEnW0PDXfii4NIbKoER4MpuzdDpD
Jpy/w7UfGiKngcG0Ek2mHeCL5PczGhaud1D/ukaHH9J46fs5bLTjmQL+CTFr6aA4
4fODqSIiKPEiHkoPXkwHQy5/AdTkAVi1WwoUhdHWNQM0GbslCs4Xi8Wb98cKs65i
ZyCoe4g2HykpLkocN0b1q8bQNv9R1sAwT0D22T/ixdcQ9l6L0qV8uX/X4EAXnX7R
teSw6vtokpzAWqMjyVD7uhnXoMjkmEy6VRBdPloFj+wP5O7RA/ZeJEkMb1v4E3ZM
bBC7l5o4JEOZsI40iuuW1YIPc3EixgJu38qKs6KQwY43txMeRCEtvlt7IfgJm9jo
R4q5EbuFws+FgVV0hzsAzRMkAjlWJLy23VgYlM9hdYBWbW2ugC9tXvgRn9KrqkxC
v6XHf4Q1DRUivootIJYzt3jppd4fePcf24tqCs5+jwN8qSRTwSo1EcRsjzwX2lFn
nrrb0ihrjXZ7dCf4uARkVvF7BX0qVMLpT1rPYRx89xH0rQHnbpeZnt3XYZOLHoKB
S9B+yDrYDvGH7+Q3l1v79vKvkbrzbTpAdDMHqiiiT1ilOfkiX4EyR/z2d7qm1oiO
sChTF5pIvTQvOACz5L10Dq3/xQosXtzzHLZsxWZ4D1ulI7eTDDglzxGS6jHC02W3
VBTsi/q3MQFrHmP1u6Hyp+V9LsfpobLWqNjZOpfKKy1CDaj6vmUyXryFuOzHrHvC
JhFRzU+6UgCVsjhDesVpwF0/684TcfHWa20Z1G1mldIguIHz+Qvh6yXQGEtVr/lY
hWHjUI92QBE5qPKAOn5SJEduJMQc42vlpGsfgmjJs77pY+HHVLYxulAqm0S/cx1V
fx0Z8w6okK/NS4fFvXJIJ3cFrIQjGIPQlVexC7bStYAvtwq8TjhOoOENs8iJEFat
YkNfh52sx3CNe1wnwIfalp08piDwjAktr7532CqafkdVhm5eFNcPKC1dIdIWfLNb
zLJrWavRFByE7ObNF3cFgsCgmZShRkiVpjdYwfatOf/VKGXK4YsO/RbsyTwnRMSL
Tk8SZC2F+UQQRGHmk2u/7/HjIJSRANfdt8C8fLrU6COFv0qM7dz9KfHgcY2S9rai
fNUap07bNmlR5CaVLXfeXG52/JeFuD0NjY+SLi4cDXfnGKpzwuYcID4sT7LPbAVr
UQejSJObXeBlDmx/cVRtLhaIiaY5UCLNdlv74SSx+GXZaWB3N3GzUgyCLcl2t3In
yvNvEqHjZ3yDqlI/yixg4GtxT/vbLGIk02BdX7YxXXyiK9jVYVwjzzQXqpi1BT9z
s6VL5Ess8ih6DtyUr95JXUrRT+0WzALbQG4oceZ7TFTjB7F11cdVSyApUzJazpfQ
U/15hVtxXxqrXCz47/JJErLZI3jtzYofGWH4nGnqg6iZGEg0Ic2cbCSnlwoGpcqo
s/RiLzbDv7fIHs/YsUGSaEC4GS9m3L5GWWyRZQ/x/TQ7r+BdmXTyulUBwxFYUmsY
khIqT10u6iLSrufWYBx9lfSNPD0heO1z53yDa+ugAJgSlIic8gnMCv8lvyScYPZ7
+hnd6tSpWeJ6+ANS1l9YxXuNj3BQVE9Np2cKh361Yy1eCY5vYFG40sF4bWe3pQGs
XbOCJWqtIn5dH18mIrzv5w6NWDO3rSGzXuuUggbUqZTZVYaVzqZrOLFocwIHAlR2
goWBhpXWU4scMs18VWq+Gn9QN73/92redB5c8328U/KMBwJrBYT1Vp2ca3wsKLEL
57k8hZWwCs3Se7nHj6kp8t4Yl1dsvQuzzikuZJYKbqqVMUcXYU0vVn2JsoODgWw/
PAd4jS8snIrWEAbL10uUPjO/xjILy/87wreioycNGCrR0JkKmMUdp7qEDMVKmp6i
BVH/s0b3lJN4WgYr6s4d/0nDtdo6KtCr4GdzTwmKIzHfN6fcnNpdcgZxTweFfYUx
pKsHnvQ1MUbLKZtM9QAEaltOS3TVgKc0u7siGluahQ33rCEzFyS2nLiN2bA3EnZb
69NDBFBKbnIKB68N45Pd4K8XCtvYMWISjQo8UlAfyH2N5SN/UdTLu84cm2A9BrcL
diVhXNalhva7UI8RTL5KwRueYABzfhk0Cfh9pV85rd+TzKMIE4MhtpBmOMdW7Tb8
XM+CIjjRol2SE2AJje8hC7XU5oicgRSXZMeefhyB4uHQ8KXKOIVrctzGDujT+nJ6
Vlo9Wyh5lPunhPVxmtPHE1GceZcPdvWi/CbgG5/txxo20lW+wHQIEzUtilCykyKw
7WaVy+hB5l2XpPglYN1hUjU2dqRbqSufoYXZKjkvOvRk5+BWQswFj/J3ARZWZ7ye
pkaSvON1rKWirLS3787LP7ZpwDzxD+nffZq1gJOcnEZrl6U3yZ+q73W++MgZekM1
sk5tdDIQXOSlhzs5A2a1zYImtYX35m6YqESzz/VZ3vwcWpZtCtCEaIfEeX+pl0qd
PSuEwV1bguttJc8GBqcFkD0YsBXO2e/5hhweQl3GHp6d/R6S9aTFFZRjn2zPXkkh
/eUbqGg3vSrfyroGVG1ZdmlcQWCZ1Fe70gCS/K2TBhd2czaAmaRW9dPqjsS2aOpM
jqg9qdrBTMIV4JUQsBEuLECExwTPV4OHZOPcW/6Y3k3boqofQ7oIkpdbciPbO8m1
jr/MF6CeiUCfchkKiwusQc56NZCKJ1iC8YSD81NXFqauNjZ9EC88X1E0G/1vVkPs
4Z7lQnem7Y1MlUXcogOU0Me4e+xToZu/Jzbu9tEYxDxk1DGq3f3oo7hl/tRv0SLD
5wVFC5LAA4MZSiZZ2qFpmdyelx3sROlYRG281RqrZpk8HY7tsKhbxMjPQKX7dmi1
0R3FQpAYjmFbnNGQe4OiRvfREEMsedkXaGVRu3ltox7aioINsxDK4CsfEmv1Klct
4pcJ/3HDi2JksmK0nCuBGiH+YdmEVPSsp00xPD1PDmPSwIN7EoFDGrRdoleIhsEi
jWmhqySgJ+7TGChw+99UCNn/r+h273h6n2/FqpWWiv/VpNRh9KjR6yozTuKwJHxE
yM7wgmzhHWtGF6icAv8iVrKelKwS/hevzT/2rqo268Pqs4PeriIuWtC7FpLFjrQi
G6voXNTUJmv3mM/JzSmwBVJi1AMbdYQjPgpqN79l2pE+2XKAOVFCAn7nOkj5oYDG
cv6CZCgMoWkvh3hF+jmsd3TxHsHT9TYI6Yttec6bT1wXyx5HTUrwVDmpkZ/3TVln
W6eXHLWMS6JGs2/xByzj/L+C9l/OydZ5Bv7gny8Ib60IS7/9fas/B3RyHYTZWUjJ
8dyTJ2zrxjRVdpNgZ+qL5i7OJvPGn+MVqvkjp7zouT879GyfiBhqJxqY5Pew7WHr
0S5lOWQYOSOKtbYdq1aAUs4ku0cj1sHGBZWSVpcBy3w3Lx7UAnUF2qrr2ZXI12/W
uCXdIeKl13KjAyEd5hcH2BuUtvqorwhgHmfvtS+87TmVU01qLbqLtmB8uQ/UYnFT
xzUpucc0ddR5Z+bxlh9ZftBR1WWqJpQ5jjjW3HEvJpVC8bZcQZaRvX7oXIRRnTff
UXtG2OO8jsxoV3RFJ/j8md3ncvvf2iBwtvaSKvbCN8JW2xEfLryXOI7yHauzfy/s
RQKsgmhlKHBbV8R+JnY+qC+kUQWHUMPZA1h3xjaa5wBFiQJ5c01T6e2J0A1W2QPy
89Rpz/QY43JKqBN/3/qXo/RHuh4+yR2Z4QUJEF3H/CtJ98puWvcZo16TGdZvW2ZM
VJjB+z/TZLLWierYVgJV7SyGtWTDZrgZIpC/SIIMthsAOBgxlZAZt4HnUVQrf9sb
2sd7f/Em4H98643WJtzbVf81t4suGGhdIvK+IH/1aHnjjFtUPzaw1gZS5JIdWD3j
xUcfAq5nLk22v+CN1jW14qOCc8ecLwehxmzYDiw/ZjUIKSx4hZhGFleB+ZeqJB77
I+oggW7fmdUChyle6uvv6PGM0FljhQLUjz6BZbzfuYOFcJqu+niC+EUKlWNNdDkX
VMEYaPtQX1YzEvx9cIbFEcMCmGTEvgkKry8ib1sRxH7FyC212sJQDiuLX+rGsOch
ZKt6MyVAvklyGZQq9+Sb8d8FS7mX/WF0m2b1CIjGOZ2ZC6tRcrxx3qHqkxyIvLr+
gX227J15OGORKWoVjOsOGcta/afdm+DTO4NjiA4mKDiWVTFma94BWyW80cYPLBVp
eXcWdtcyjXaQAKsdW3VMle/sdZQENHKQXjZ6LKUqyjKySi/cne/3RqeWRTWMyHKD
Nug7PQ1mrLgVyYkBZ5gXRk1fDEDSnfMeXrpONu2MT3LRPJRn1i35vY23uYrEvjkp
4MpRVDFinikiK03DdNb+TuqIdvsf2WipiRREZKOZolaPoG1cYFNyp5VENoUrF0L6
fr0bu6tjiaTe1f+bMSajwnuv9l/0Eg5sFLSdAwxgLsh/Mg7c09kMHiTjQdIMyqef
6kVP/qArfdv3nsghmbDdz4dyVbNcw9L7Qeca3kNbE6GYfRXiBITvGcg7+HlEKm5i
BiDqd2KJ/AHXUY8s6VuYMx2CyhxpM6YhKy0cxy9U+iKYywv8sdMuaZHUN5w345uu
l+MLbAz9PjUFCG//ewuiHQBNpUxePPq31Wi6WtPMANOX7oI5AZIJzKOHorw12Dw1
pk4vl9QoQfxq2Kv8HPjrO1Wiubyfdqra0lSbWS28RK9ZsI5CQ8HLSxMO9+HxjOl5
VHL+1jZCOs0tqXxuxQplH56bcWnMoUIVHexIXg+L7y7xtFr5OqpfSq4eeP1IU4lh
uuYZ4OA1opUrELJAWAnrsgZgEr4CkHLroAQ6dmkd7qXUgsqwlAetjEeoPCF8ny6l
WB/Mxp+0IgSlWZyDE1H8RJWyRiQxwMnO4PnCCkYPVWdNnhIZrvm9uzz0yHLg8geI
leOPST4ji4bJnTu/VDq/wQYXqSblVAWhYaeDeqLoffjmk2oFWJ8IvhELBZR464Ch
Wpp/U6frdYHXbegkA6/ZVg+UWBC+VD8Cgx0jiFDjAf63ebDegDi5hwsCAFMRijJI
bRWe4Z6JX7jnVSRE9I1/XylNG9A82TNIsTNupl4CFAlMd1kDl09d5LUOiZp1reTV
Eh9M4zsHYGM7WMVLyYN2SMrqPPcCoesbPISpONjNLjh+KE/3rMkRSW8HzeYUvjEw
7w//WIcblwGOvzsNVL7kos1xpNdAvE4DWQvjKmTHuchW8LdTe2ITC7Er6LcjFgzK
+tKHXUiI2R96Vt65xwqdEdhG2D515EfBkq0WwBbiFbRqbm/sD/6GR4IDthzQe3je
EVKiiZiBrXIaO0719GLtCQbjeFsUp5/pGsNZzLyx7+lnbeswcBgtmA7E7LdvLZuC
d8vqwtSVzaHKJHuxz2nfXq78CSADSsi97FZZIAqRFeY10TM4H0+WWmsQugnBiT+b
hCnhMBHK7oGqDAFm8hIcf3HgEZ4L6TNBGgkIO7g08CIwwUawKlpFCs6rvg9VojME
YXzdDbLrEAxHWqjn/Gur6cXWOltT0y94URh3wxd9/0drqv3ggdaWMBqBKfQtIEvA
oLnCEyM/ONRChTrPNy/qfeUgA8sKX4mItH37ylyLZUNQs24wpGe6qls0xtniXkGV
9Ted4Xrk0DIthuJrZUKIK1bngaifkSMxVXCtdcbzFqEFf89Qb5/MsQJ1HwKxono6
KssH+nbjQocBOr9e41/Kb0ZQ1DYwT4D69KnigPVhbK2PEJG3QbgW1cQDRp0sZEyv
V0m0xLGtViUCXNE5bW/dtPdaxVPUS2y5sKxqaugvcCRpwY+NeC5k6QIrJE7ypLbt
XO1u9flUqh236fe4EIQay/3wdyWwNFlhQdLJYsGDKAo0H5403aYAX2mkLky/eOO9
QqZWaQJ3HjaWZPFf7XmwEaAfxtSCEfM1KRoNKj3A+JOxtI9HokGsSWuCUjdc3Xe8
sJU4VsTdOXXnZBgv3mypgoesgQCbXHhT04fSR+OT0RVP8JiGBccqMc7S23Qve2Sr
zj2gUxSjnKx/azb87gp81qYLGQwVZocCbFNLc5gqhRXhY09OLhq3QubTxQqGoNZF
xlfUhKIoKPL3c5S0puW6Edk4IOWaJTj7gAynAsuWol7zQdjabJjjSIbYGuAdpIgo
huBF/3QFXYJiRM4S9Ch9mQ==
`protect END_PROTECTED
