`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4RcEFg2f1K2QaYLo7b+JqAlh+Ekg1bERoKKmkQ2CCvHjYn6WQ62QCr9+YhkKdlQ
dc+R659+P32Xu7/YmyGpL6wTVLgvyEcx8Ou4IQKg47Pl7Vh4mmgHTbM+QKACoMYT
aMWZaTMhvmwkMs5K3llKGPF8n/drAvmOHrqTC/Vg0zmNhxLTik0rTZF3CiNTfTaJ
hj/LeX7e1EkBOaafKb1zkksLdgDUJqC4kcPMZ1ELGuJkjmvcOUGilUTOOVwA6BJ1
PejFnh9HnZx07iUHZiq1WFH+/I5IojBw9Obe7TgLU+nbp+lwUpZR4MXr5ZZbMZBs
E+YZaMhDCVax9JardXJd2kesYMCnUD0EgSMN8Ey3ZmQzfuFBZPhC0xZo21Q9RdBn
kRbrRq3YJ21/CIOiE8yaBkEd2ezquzti7tNQ6jbZ3h5CTd2Kyzi3ZC/pkSu+d/+n
KF1VTa4PuGjW6Wn4EmbZJQICSVvgo7NOUQPZI5wk6op3W7Xs9x9VpRs1PVn88VM0
x+GBl1SEt38DzQi3y8RPjnaWWXz4L0C50alrHl/V2ver9xR7qFXTAJLMCbQ0QTYq
fWHeI40EUZpyp0zRtygOnJ4YHQ62AyCqrHyI6AW/H79G9E3l4JeJjKxTTR9W8EQf
TcH3sAJnHYSeUMhJRU+AJCdE1zigYiNjwpj1X2nIdIOzbZAJRPpsRCa1C5ZY3ft0
/rImj4W5YSeaWBEiQiX+GGeXxd3ByB8EOOia61Io7sAiubMA2lStUCweyS2+Twod
lu6JklFtgoHzRkKZWZXCC2foPGGgYUo4GWPuRuJg4uMii3KZxq1dvCnbBGRIlIO+
vGeZIep3KJu0UlOxcIFPBdzGqtJKGxO50WRAXduaMep0XRvOnD4bzx1eQUR9cCLu
fBFJFdz6Kz+5pYoCC821X6VSrgpRn0wm2eeHKwINxy4HHUfPgwiOh2tdOOJyU6x8
yGCVziI1rdw1mD4iG+uMXlWTRhkkEnJrgUJTibScsVIvLZDPwwDTT/kwVzU7/pL1
xk8YreO9TK7+csVLHLC+F2HBfJ4FgDu25cWxE/bNrDpKqNIVPcWVAPm5ZMGVHHTn
Rcr5z04XcaEgHg8IFxeYksZ0gRoa+dXnAch0UtIvpIzjCp2ZR/I5AYQRjsyuHzgh
K27ZZOQCFdX+QMO2Mqd1BtnY00tXrgODqcBk+WcH6GU2Y+O01kGYHSLBZA18anL2
VFqstix+2vA+f8DTJZX8vD3YzhZ/hxFRpxgyh/MnOIuzhiPdVqqzqlV3fx9CSbUK
+y7OYAY4cqjnc8UP3GuNXHKGhuVoSToipBDIfENBakENUGbW/GgZqcHYGa2iPpk6
8n8Zi1u7mLwCfjbK8cj+4kjneY7VyRWauWm3EWkBd3RWc/r1wqjvj5DdJx8B+nPX
xyqLHyvnXZCW0yHpBliOY82RncpmjcofqwtfpYMlxpZjr5SQZNrSDzxOlAjvhR0k
EDkj++GYAA2+mmDyTYz7wnd9iY8APq/dmWNwMeCWPb7fP0BDpcP6+9Eh4Q5pzHTk
0h0bac/WfEE5CswwDF3A88tfxBkcvv6x35v8prS9NcwC4oetYM6aArdqrsEM2o3j
v/nACAug8/++LeB0aOwo4qNuf9qVfaiyXmr9SoIZwAYEhQrqm2GrTRXxhiy5F9th
sDA8364IdGSw2lAyaQ34nsJ6LaCMf4oabMP6PsK0gb3wiIlNo5QuoPJPOTRMtoHI
SVIWSgmVPiMaOANB9+xT9IzmYH+mYBKgUoio1CQjbNvnEIzI6Kf9srs88E07XZeT
SzVa7UW+wUkH0jqinGcwyf19q3JeXcL4RW1jeTQnlXjHbrNshMwR2T9WD3Yo/Xy8
MBrQkwbSKhSbT0eooZeqVQq5wJA4wb6AJajIB1HBEEqoMlUORT0o4gw5IGiGdefp
SRp59B4skK6tyyuTyqtjgbCagcZN6X8fQj6a+n1drCjbvktTKLZUPyjeUOpXy6dI
Ur+JFlUsI86hX2P5dMyaXAWvvdFZpfw6t+lR8mtxxD800mqVUEJf4Z79aFqbwo/B
etC21l1jyfxeOc8maxEO6AEGBQ4OvSHvBUtZVaWI4cEUFmMT9bgsUacas1OpmUOl
0cAsXJahbHUM6rhfMOq56IEt+O61hElhDXzdDRS65+yEuSen6dLzYCw0Pe0DkemT
8oeyS1jlJ/KsDNYD4r6JmcdybdfD3AqbVg2TIzStsYeaYIIe6fWcWzyL8sY3YNct
PAP3zpkp9BAu+uvzHmLrlE+DwinA5We2QAAXOWnysOszq3stczMXtavdKKvjuewn
8DxCTVbGxI/1NP0Pwx87htJSVvZ2SjNk1nTzEw6knWuB6F6cyzH/XxT9hvbsgf9G
eEhO9UoFINMdl2AcZDoHafZhMCdA3nQ/gA7sAVs2ycqkIsfx1hvdscGKKb5dwDgV
Anb1OStz8UwouL4uK/AC7PXOSlBKl02K7LK9EA9H+d00mEHsh0mPbqyrTrHFTjYe
`protect END_PROTECTED
