`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBEws3SrQUjh9QcbgpBct3krnWX/ugG613fBN72r1CclV8aXQr6+IH1Tw1TFev7V
MayzaFR26ztxjPRjS73lcYayAAQDF7fCVzSN9VaJFwpObMuFS47EhrNS/0LQ4VAu
f9wfenCeItW9e/K+YwZD7IeM/HVbUTq1VzZ6LQvC8UoAfTTDL3M+dICLKfbf44zl
fidzUqlR2raQT2N0SLWok6C1+zwY4Q7gm+mezuMET+stU1pmwnNu6hjIB+BcLq0M
lKRwAIEKu4fipB8TWLIOnvtcTUA1+4CZh37d6WQMkhMXxZeZvVGpJQ6v55XAugTQ
f1dIEDbbqEQy4bI/W6UaOHNbAXW9KY9mCQH208fZ9nU4REtQk45vVS3nW+fs3KOM
o5CeYfb9TAin+lI32A8BY55YIvQIkwFC/RGH0ntJgpHZLw0ilPKTUyIDIc4U9pFl
7gQP1fwXhCbCZ1GZa8fnPeP1S0BKKAwp1F0iZJrORmfH83ZGjChDn5h34hxVD6J1
`protect END_PROTECTED
