`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iUavZyXhiaCP9JPfZwUeaX93q6nWyinUwa8aC7R0Z9d8Lcp+DUjuSJbhBGlGHG4E
zxzr7oIi91u0DHs3/lcGF9hfYxYZJuNQKyGIg37+rujIVZmu2s3tAyegXFM2LBc/
MH6Cjx1XfwoiUzYIRH3KLqH3Zwp2+sB4YkFBpMHgURVtQnC/nE/VPVhlc99vTiKQ
ijPpRm2iTIJq+syI3dIgOsM08baY50kZE9G/JnAvOAXRq3sWQUPxmPanOKqmAOYy
zpGBZ4KPRAXsfs7pljeOnk/BP55+87otdkkqdbMqjVFOAWVdBWer1rnUzxaqm9tr
hcS7v5bRWKQg9uyo4GhNd8aZGGgW6CCjDlFtbsXNlG6baoUjH6xR9WYSnqUm8Z5v
KZ6IW0yqcSu9W0u7HnN74heXhtmkCVzuUX1vS+pXepdy/3wpJd1eEFWFzmT3/lrS
DDww9DrGqpSGjxoWJtOIuQYdBXC+CFu1H7Gh+WDCvDo=
`protect END_PROTECTED
