`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Xpymxc/y7o9JoHvnyfF6+HHfYLueLcXTfrnaGcFHtdZPZhxQKSwJDwQtfCQxM5A
PgWi68Zb7X29gSsR0JFOj1WC2ddFhMqlL9kVoHKcl6fpmKKtU6B3K6fqEAOPqkmq
3ezHNglHHV3yivFQL3AHLJmNmJKoz1JiR8+zPbNvPtJVD0NVCMqFCGygI82/Nu8e
Zgj3To2zK1zEqG+zNkAoKy7Z5Qs8+JsS34U9IOeeqKLGlUdUwT2dpkb0kllZzBw9
RtiBXCNBGpBXIe9bmfmqhXzWGMGGtkXofsv3TWok2y4dYKJ38VM95Ia6tMiVc8eb
GTzPTsYGB+MSMeq9IuDNQcclzOt7oACRYumJaBTqVJTi30WglwOtFrXCBv7S4hW8
6a/RtpWVSoQRTqBgtIgC9fnYjtARfVrdMB4vbbTimx0KeoQYYJQpMrTEGo+cVmix
XMLKM3nSmwEGO4DJHm5r9eAj9un9/fAPWfdQcvjKVaTFpaUlC54KeTuhDbeTmccd
K9WwhdcnZAM7bVQzA8wijYg+wwsLhXhidU1/ARphfBD/0yF32i9d5hKmUguP28hm
Fly037n9i6XIJamuAnk0QNWP51SqIfdxnZQ03Pl35LVoQ4CHxv9b1smK8btThLBZ
cefaett5WSlIWLLWLji/npoAJnZBR8G9xtaslL8TfV/2RGEljDM/6KZcya4Aigbg
7nsS8b5V3r4TZplkLTlP2+Vkk/5iPjmr3EveGKDBQ4YkLGoyjOPmKSDIqlAazEE3
2PVu1asUQ5a+c+u+qq3XIqTMoB8umEoknvVLIrh0sX8K1JiY8qkXnQ96ffHlASaB
bWUUuA7y3tFVrQMq8p1V5uyMgmG4EVYrwF/RqOznA2z7sWRbBl+MjRSAqj8Z0YHn
fVHVexh3wbEsOECwUaKhA9ub+0dq/1CMP6XucYuOZUI=
`protect END_PROTECTED
