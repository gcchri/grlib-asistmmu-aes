`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v9mgiwJgQbvVQiSdwDewsKT/BJFe8OR5aq2T5Nb+kokj+F+mkBjKFHFqY8H+sBFs
rHKkRyKCiNcjEEbUVbhKAPL1Jn4UZNd6Jl7X3hlDlVrxE7ENC+sCQxGcTCSYsooG
A04O92rmtU3qOWrmQFKQvVZEoSDuc/3oFNRUfVtmoou//EZqVwDi/2Xxw4Mz8u9e
aXu+34dLNNqWF2DDHwSN+EUk/PMOb4QG6aJfu+DWHdUgzI0uRCxelq+2z/e6SOx8
Wv6cpvNDLs/HveRm7g1aCUhMaAf5Glvjl/W5Kd3CFU3Ze6VJr4KQfdsSxjflwuhg
3XwAa83xCxiha7cGdEFXp055k7K4VB0ylG2fVm+8IZOgxy/NZRUMCWEgPs2yLESE
JdJRJnfIYjaoD8ST7SxxdFwKOBlzzHAIy8fMNE38DX/NVS8TTvCIcxSxmA2b4CTl
RoyFMLufIYft3IP5t230nvgMBb8z4gd3mK2Vl0+ru9EdQc6427e8T9K/71cEtRSN
adCW9GLcCN5c8zIsBFaYmt2U3ZyEYuJTflPaq96mHuKFQkMxkP+8mRJuvbAMD8l7
e9Ux39BViMrs3MObtr9hAanFSXeJmDwN6qFuFE6jP73MS1cOdXZ2NYZ1/m3jXJTH
FZjKUFGxV0XHp4BnS9cjJ3j3tcl/NrgZgsYkwUiUPokoE2KsWONYq4tZa0OWadlc
d4oDREzM4Ox5CuihZjFmTw7+utRqS86UkO2RNq8O/v/1pCB2/yunnBd3LawvtQF3
iwJVmueyOcpfv17nu5C3xR4Buk4zoSQao3X6PEVhAkHuTyctgl4fRXfuqDIAnOeb
HuPIT6zeuabj0Ggw7EIAdxUZakBEVjbD3VOlERWEh7sjit06nR6zp/tHfrsjMXlH
jnjok3uLPtiNtcOW9gplsxrByfO8CH06Nm2WGpsX/VjufEuFsseRIygzOW1c3Cm3
NitZk/u3oQ7TOAzZ+3bxCmiYsUOB2/PK1OPnsgDv0mt2j1zhSFpz7CEWoGMb3cSH
hTHyRuKJPlW9cdtoUK1r/VragzXt5ZJPmzyVtmmvZqvRUmmInISq6QEJYjcZT657
JMqvUnkzowb7UvFDEDQoYarFvwzMWq/jbTLpCFfJeuOeLxTQNjcb9VEuwZfDlYf7
xedoIu4HR7WYNfL+vuBe3T06luL7FpuaKH3O+is0L0XC2ZxxXB6Auvar+y5fDbHH
Eo7OVclqWLZww5PPQPEaLgghVuYDykWnHZNI4LR/2NSv+tJJS+Z0JFaq+TFSeL3y
N2jwGJdi7bsbVTzEydAe+0/Yk706VczVlpJ31744xPJ+EzSM5k1xf/cEmAkGBbhX
6jUF0Ge3ER4ZXE2MN/rlAC+8RqceC8MLZlX+gaoDl7g7S3JdgdDgyI6pToh7FEcz
`protect END_PROTECTED
