`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O8Lp06IaJnwP6SMoMKazZ8sRiPmg8pHqyjoDi0xefoag0O0sDlyPNLJbUEdlZ9+L
1ScjevUvuG4Ml0zLI8cvspQypT+UAk8GbXjevhvgNoZWbSuD0/SECiHZi4JQKUgH
33OV07jjAD6Ik5wt50AaU3cUVYEQ84mjPxTl83trYyfP4INXGjFFAQiuRTipZZuw
E34si3tjP5idACZm7OS4kkxH0GTeexq+wAEsUxY5MVuGsDX5pgSFT8qMhHfWOt7c
LgAHopo+dgFGpWoVUKFjBs/1rQy/WW1sII9f/SYOSu6332Bzqx7D3Haz9CSGsaVa
WwVRDr3cqVZBeKY8zZwMsfYA0bL4IWJfcRvHWkghJJiXiJBrLKxMs9W9NiQZwODk
7doFtvFikmYI/R4EBP8PV8jdeuZdUoTzZF8Z+/5y0TiHTtgsWh8DKCfjnUL/WIti
9QuvyVu/bthrjgrAEA9Xhx9KZL7gzJPEqNzxuRLXZ67CgumuHuUHnm6y8+keIbLY
d/3QhK+afyRfR7r92t/A8PRodmmFMnWZ5GPK0I6BRMq5U9MoKrdW1PWcdprvj83q
hIge5O4/zUfwoYU2yxW2he+cWePSvKvUFwcz829X/fCT8J6gEQYN16HcV/Srv+uw
JqVnLGXyYtdpe61unOfl1sG+3R+vRJrJqFC2Ou0efwooNQsHUgXHQEykTuTHTk6A
s4+kI2qATJaIQDTqrWfRwIPaHo87rQv1EEARo+IcFnRtVOxXFTiRQcjdmAs8sAib
apikbKoaCXr4Tdz5Bvew4zOlZJNZZi8Kkj2hnOM0NY/XA1GvsqkW9HT/O98Uk0pK
ihbcD4hwe+/qLDqUXDsrWg==
`protect END_PROTECTED
