`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0orOQWo9fAXrQoNAb7AXITe0G3z5Uj37S7CtLsIVffDS5LIrSxOI2qzBhjjyMCTY
PDtHGJEwmxJhtHfm/6cYB0ifNy08wFMDYli+V4Qe+hidoHyc76yorqWi5B2y9HJV
MDDH6coaC7wCln8lasMtXzCP/0sJZpmWsag0o7SN1gMyFcpPlVGULUId3a0GWWC0
20b8WKEXgFLDLPOgt6Vx6pQJRhspFeNmWB67B+NSKRLaHWVOefVXyrAmPoTJ233t
ei/N1YWjfjN5Axb/DlZfix9Rp3hdx1dJU0Bx0ZNdeyDJwvfjPy0fSxiI7zAqRrmV
sGFI0GqaKC4z2r7vfJ+j2fdJV+kCXJq7GIcel/IAl/h7AXq7NEEaZgzJ+z5qd9Gp
leNub4D+kYNK7/4ZzUtlhKu2Lmws9gb1WOPAggScG9cdMjxZh/OIi2GP5Mn3OOvg
Uq0Y7mGCZtfZnsybFx4Ay3WFmTlfgUkZhTegxaKrOYY=
`protect END_PROTECTED
