`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HVpG4+ReZQrlo73wmbW+xJz5UkTInlOgcRi8NrylMVoJdoNv0ws81Jt35DoXqSZW
CWAN3iTyYg2Tut/qKKuNvq+hfgHFH+/EnZ4Y1F/Xuk8ynjX//Dr2B6AsDI1pYILG
sQub/l99x0i+UlpfkW6cUU5upegbI+UwDHjhce9LDxUvnVeTFHflDoZyjmY50lCS
98ySW3N7I4oarz8CXBYk+1cws9fDSQEJhW2QFNgTIx8q1P/dvj0Ie6wDDxO14gsa
NwWANGKDAwZtcgPedXoxXVvsgVjsemL7UUHghCecOY+PabN5n5JG+a/b4Y2FOjLT
DV5K3i+KXpJvSw8zh812mB8Cp1HNyt5fHVtN4EjrJpwStWPTZ6K4GHO/sbOyHsgm
QVCCfxs5830Nfiw63Fh7dN7KlR2//JWw82+98DOE4JWLaQNkpARaEhwBhb5mEEDF
SXdeuhWzdBnbMUoAcYn52BX6fIN8SzkIJx+4zTO7VZS1Ay/+nylIQe1NCbjGF+3Z
8fr5YvVsJ8jK9kaT4LTT9LMGD0hKNXaSvFsFHArITFBblpGWQbfJQNAoAqsDmsu0
F4h4xmrxAyuNhnNFUnurpw==
`protect END_PROTECTED
