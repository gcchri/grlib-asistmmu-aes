`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZHU4GUnbSjcQkOGdKE6VVg6tp5xBet7OvfnskGgZdDqL7paNUSHCWgrEaJumrI0
KnhZRKusFGjBSh85IRQNweQ1yDJdwy9V4ImaPxYjuo76ycieUCG0FQoF+i6s9yr+
gfqFots0RpU1kWzPqE++T2s1UCbLJohMs8BODaVxEmye8N7v/kNQupJgVexXgk+y
N8BPYtdZk9m6ap4sMzZyh63Ahf1yqnwjY4aXcn3eDluTAwDJDcnYCoRVLAGN5rXM
j0OfhpoMQ1IPYZPJE7a9hrlQ5e4bTHAQ/aTLdLCVkCdEKggiCAawoGagA/acBl41
9TfdgXYku/CCYMjsWxnyRA==
`protect END_PROTECTED
