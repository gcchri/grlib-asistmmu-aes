`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxXkuidn0zRtHt+eBqQaK3mUz7pYgQjakY0n2yQbPzVOXVp3NKkLWHRBsd7+mxdR
O3tBbx47dBBRmvrw/6P0wVzkCpEpUK+P3HclDfjTW9BQff84iuX0RTXBwmUTamW4
I85w+IRXEF2iSreofmrla1NbtbAoJtykMXDWAC4i7gA24j20zDr52jvEOreO2cVL
E0XRUr4mVvnCK6By3B7Iz2JROQw4VKjiMaXx2qYI9LNo8PF5a7NwzMeMhDAfq0G4
tUjKY06J3BKAIMVTuHwuplVG2haAXgyngUzJakz5JyaSrvEr0M1l+LiHR2EgOPgA
hxsDAB3Oce1O6QxDDoGgjefE/MQ+ItOC9N668NWsC0tIevdcRofr7eergdIEWURO
3Pv4EQz/KFFUZFpCZdxJGO/t0UV4L0UUWw08qrhFNTs=
`protect END_PROTECTED
