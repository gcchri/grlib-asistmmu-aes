`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKBhg3DxhxBpI3GSpKYD5D+BLNZIn7aI6CUWrurvxI4PtIvJfJr2BhkqXGwqtJN1
usJYmyO7fXwhs0o3+tlPykhxmOKo5VlsKgQvTcSfkywYU1Z4IMn/nGuQ+DzEGk17
OrlAhv9AURmQ6gnSWd+eO/pVXQ4E2py8dZ7iXbMwjLJ6cUnT48KMBIWGCKe118b/
1/sRDemxSrTyjlzqhCgg6Nbrtfb1u5W+kQcLbaiJo5abYCwhHuogl9wH6LYeeFlr
YeiynX3NQbAsCL+e3H9FKGxwvGYdVx5Z6uhoXJ39+ixHDCTlYzbjy1tQCcJWo5Qp
b+4oy6aMrxMvaIpZf9/O3ON+1OZK6025LAPm4QVW/DyLygbblDdNbToxwh+eLOg+
49FnSesykHc95eV+0YiaXar+6+c/uLoQVXaMZtnWSWbYP1K3KnSIpXZB4C1IW+jB
ONPUIn3WpcDJ/VbyQr7byw==
`protect END_PROTECTED
