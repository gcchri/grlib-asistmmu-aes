`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HqnZITzLxfjMn2cJ5+HEpz+xFXlWasGlERLQkjYZUpTHlLdBzuWV4Qe3znhJVU7y
CWcusCIsE9+94yGk9m8K/6pkMXQgVtP1am57zZHLzYx7/BCAU4pvQyRM9MkF5xuG
I66ZTsuPMBhT7UJT+cq3Ro/Q+1ggi+t/RdivwfxMHs2a/hWEysLKKOmYMACj0iv7
Dt4V/ibZ0tMfoNVx8yCvCpN9BJg3vPZd6kA6zzkIeMJOwE7jh3u0ZT0RPrHD8Z3A
g8vA9IcDgvJHVEzidmZ1SZIUgQ8ch+OYF5gPGnVK+ccWU+umBYLxY5auTHJfk+mS
mFabgywvl/yw+qt3Ij/pFq1gP6yg+muHVqPDJ3UXQTwnWkCNFBmtWYCbmNPPFZjy
`protect END_PROTECTED
