`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7GCY+1IV4C1wx2RkQV78lQ2Bja/v6CfFZJgWxxTqY1hrCvly4X8HBZaQKHXGBsxd
nCpNS3jSVCl6Zd8sx2Ixsa4f5qSmR0qGkGI07siKlz+sYKTY+2qSN7oFNYg2wlTy
Ql920K8Nc7w0VMwJBG6SOcTwNYbbNjgCubnAP8zVauwk5uBlg5Ipger+qQQMo3h6
A3AfjoQXRtktEBe1GCrFtxSsjyeDuQpxrlUTf72tLpiwE749Du9I6M9CFUJ8x7o2
L33Z6pG4KJHMFW95eFzcdeAdVa6xVzGZG+Mn52vT+Zm3pQeCbvHPkBfUGTGHV1Xp
H+VF0q80VNPKHVATCssSB33h1JXuoNFuEYndSLYT04E0g4gcprq4gQgmbulN7hsS
0DqszTyzRFbexCWl2NnmGg==
`protect END_PROTECTED
