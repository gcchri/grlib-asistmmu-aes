`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uC/RnJiBIYq4P4bus7jlRaCRqCBQJCtJrkrr8rmmBrldIUfr/AoMUvzmKTk5VqIS
SwFqx8DCuR5+fsfFgM1MFOx3TVzh6DS/xv/1Wh07CWKw3zvPq5EswJGvWokjwMhx
ZwnhK+yYTW5M9xq5UH5h2YbAmlaJZyLzOqk7GLrZTFTLwCPlFAWfUwLWqIUQSYjH
l+KAfMMgcWdQK96yhXnbNKAf5vqDhXzPcwxlQryGexW74OW9a610FjF2MXEjmLsm
ZQAndaXkyZMMXt6vNw84bA1DZUCrO9V0sb+3vxSDf9dQtODMryHnbV21mnGdaE7z
1GtALHBPlulWNk0AaTB8V0FoafPa9Mc7D2u68+AKM5sm/JCtdIDkTFld88h85St8
WJB1vLa5OJ7P9UsWwlAN2C0hUCvzIn6Qk8KDb+7BI+nSzS2wfbVo+nvmx0GCDnMu
0ZchbZ/Vmh+OBG/jlCqNNuntkXJcZObo89TaRk4jNapZKdLGrmmWs7RvDvG3c9Nl
PZFy6VSagQwekEMsMk7nJYfhsQCUtsiyExSqGTTn1oTNI56UN82rAd5ei4CMVuck
4zmRh2VdO7CxI0Bm2KYN6h8mm3PldIHnKE1E8lmJw113mpkIs9zX2ij4LHeG6/tg
CaTWvEQnnpZul4gk/s1HeHFoksMvEvlFT9650Qn98LPjDN97LPQuijVLBv4+ZEHm
vRlhfAv0r5AJVgTc7LGohci1Zorv3sKBVT9ntM7cDUyTauFGFf2corFMPPMgQjC3
6ctmgJw+jQYXCSXZb4R6K4z1uQxlfZg4n8mR+bbn2XFsreyNcoqVmpSZGCUd1Rpn
Ni3oq387QiGwrBvvaq8svCny9frSuxbKJy+WreRlQ54nKnLgkxUa8naC/Qt0oz6j
b2XVNDAefRBgiQjPH6rrmJtygn8Bo+Y/yJrpnxRUdTf7XArUi6wTRnBeqgCR1gJp
DS24Oh0fL6M66m4PhgKvkYvw6sBIH9J/8SkiKOxaS5JTe3VI3za63GatB182fwq5
OU0/jgVeG2BTdMfL4/TC5AT1S5WvVrfkQR/wAvF/Ju5ZPKCAhb0sAlSO1rek4xa7
XXdcznrcUxNeDrVOaM3Nyyet5OX0eAlP7OdXrvph2TMo09TTCYUJt+WIa1u+4pNb
DBNxBJNIaSv2b4z2mwkjcXYnMLH3tZYY/vP+LE+E7su3xOUNKSSaoEoNL0Jm0Hfn
bLlN8MHVjeBDRUllxA8LE0O8ZZEDbh+RpqTtuQiP7miZPsx8Ae4d/iqIiaOmRY+H
AuIo+xWPhQ+OfSjUIMk78YqCEIAyjwJwarJvwcwfqZaTCsdmsXzG4e4+hezcvD8i
ENXQo9lsFJ+rDJ69InJAt0BPiHtYPGWQ/JyN5/4eRVyda4GO0by2WXysMHj/sHnJ
2D0alRTXsF/7106WLQEVc07IVNaTgKFC6aYsWfLCr3i1O8KAsqSer+e0TsxN5Wdm
nfeRhl6pg5bVc9L3e89Z3CerIMKNdZHWSrl5qQMytGepTQmHANvlNPq+hK5cYys7
CBKQJBBRKmQLdEAEX1cPS3Z7c0i0yurQhPCdFmYrp6ZsTaGTcpTDt1WpfZbxxiTi
5KXaDFTofLyq4zms5wY70wWmSA9wm7O7dzQxt7R/k30rlW+91f0e1ffZB/4yDUBT
RdxBQAwoSxKQNzMI0k+T2iSwWilegDtZ895XnKldKegG/sKf0BTnaFEvK2A//S06
mgADAImWultiAx7vEpx1OohW4PDlCzvfpfgEvs9A4qM=
`protect END_PROTECTED
