`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CtXXthMxHUD40C+5/27apFvogx3WpWuHotBFsdFV4LLK/5G3XCn/d5R2nRDRByOW
GpKRuK5FiDvM3jMXlfJmqwi7ZU8dBqIj28YoFCzFZrP3NZXphiJNNTPS7jirpAF8
lcigkQMKqA08WMPcMTNcn6aSZGOxRikVLBWPUzF1TqU6npYTTtMSEtvPKJ5QsG6A
oU7nrWXzcYLzhR/azYni7AZ8OowRxRI0O+2PTfVLly74ID2XTZYFyZ9kD510hPy0
ZtievI6ine7p33tRXQ4wbmabqu0yr1ipmW6j+rQ6zzVvtxCQss9TcBDPv8hN83Ks
duTxtUc596yetJvseahwb5aDUg6bhU1eVmiBUiUOkhB+SjvJ9bpl2JyNzjcyum+f
KvUvsIRRzjskaBZrHsMTHSwJPlaeKOR1mLgiIT7sZsUAmkSZy4HJOTP0++RiXgGI
vEQyh5IfurLdPpDBldFwbl4bT560LAD9dz/nZAayhCI=
`protect END_PROTECTED
