`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RI8YNhpjMHMBSoZhT84vUZdePyj2x83WzmdgiIooXBTPlc6h2SYtYq6ekodHlzv5
bPvuXF59DRfBV4dBqV7/4gKFSHLkRYjJOkBCDUE3utDTgjV0NgqirJJzY+NRzjKd
2P55g5JIl4RJ5BbBrFJrrwyEHcgCdX5ZxBxoV3Ctfwg/Cq0R0UMmH6iuN1NZXvp8
jPJq+bEcPJ/+MXmiDum2c2UL48HZbwfMyK9WBZasVtpxHjrLlmh0JYfvzeNQlNI0
6VmwuKkbKJq0YmAs53RWM4+dE9zRSo09SywtH1Bl4mP642LEFzY8eKSHYiuvB6kk
G9cUBMhuWHXAsshV88a4UEnONNaa0kk0vt1d+xXf681cZ5fWgXpnkdq6AiXzoptE
oqasDDkzYplN73ayq03IFiV46my76AOhIm9eGh+k1AZSbDggIX8otFjWjYi9MQ0E
384Siga5wXc0lMdNFL2bGi3MqSsrjHjoEvq8IabvELkW/I/2fjZWMaj4XxK2TUMM
aYvibArDBTRtcZp/HaeNWlpUvUAMpaI7laC9zIeS3/ZhzjJxUf2VM2IhEuP1n9BN
xQh3FY7/E3MlTSIFG8A74wKhXV/ltX4QLE/LFuxD7ddoeM0fVdHfa/wbZ6oA+0Bt
DJc4NkN0YLV8rarSQRo0kqbz7/yFNm3odJEC+4CCeOp+k97j4pWxZxg/kEHmyzW7
Mn33gcApcbDwR36FxonmVcdJ/Hsz89asyCTkZ0lxSzdt2PkNxM7hL60HLCteo6Ad
BLI0kMt/Z4F/82p25dP9EVyPFe51CV5JnStqcA8996DJAMd+DcUyajy8b2409JN/
A+vFUQi33j4V9ujDC2N2D4dySrqm4IDrJWiaxD2Jq2UP1EVtAEtwFpME7UAMTs9j
I/hSASavcWkaOBT3Yuxtl/EayZh76m0IYij9aJJ2CmGugn+iJjO/N9GJlEdhKNJO
x694XOfjoaow7iEp/KKRHd/IifL4pZ1RwSf2vr2AFI5EJDKRsGTOIQ6+1HFFal4m
`protect END_PROTECTED
