`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vu3THMKrQAnmjKj+JywCbaL6GU/Hv9Uv6HflTB2++upb27fwDa1S1I8grK1aOE+g
Sa0iw1weN68Y23Qnp3XAY/wzzDwem2CfGAR0lyZg7GST/Bj37DbOZUyY7ppLpBFM
hiKYFoJpKYll4OD7YKn45Kg7TiNeexVQX7hYiw4soCNrJ7Xm3Hq2tU7mtRjdBypr
FG5ZVBq8UXY6Sw6JwfAVQQJAkPcqBpWNmER/j5svu5wTzuEZLTL2MsF3FrCSZErS
Reu33vo7ALTzyL6JE5jDfUWXmNmzlJwiCRFkZGIuoRF3w2d9e1O7v3yqnsv9tSrq
aIQXXOeZ4Do+sP2FnXctTZf1/gVDU+ok+c8Px9kv298=
`protect END_PROTECTED
