`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OTft/Bbw6HhJNxia3Te9n4evNtwCSafSXzYJ8VhDiE3Z51stR4+Kviff9Ln9/gco
bLQgPx00wjvsjOSUlx3DIHhnn/gqDk924lCtU8DZLu/dT5qZEfVLd1XwCOiQ8zPQ
gmY/GQg9I9cR1ZSx4cjsZ0Yaeb3rj2V5k2MLkVVDyPiA9VBCN6+PdqfjHBj0iqQ8
fXlFdSW4XgBkB9Epb6vsSunjmZlcIGVYJANNGtCLPN8A4/qe0yVKF1biUDRSAP8C
7F5EYofSbIksSyVN6Bj3mjY1AshahE+dlDQI4SOm0NCH4HOO4PZ6TxO1tCfuVYt7
BFPINRykmLr9cL2FYYvkvvqYwMIjy1auU6uMBqeXWLtleYCOv5BMGMVvXwIgGsao
YwWPvBfBuPE4P74+27DsxBbzTWfI+9qajN+nm+yHGFpH3qNc0s/ecBtjeoCtoLVR
54Z/juQ+bInkR2k17Ff7SpuTt7QMVCgilDLp/eHGQKIweuoKQmkPXc/gVS2TAs6l
tge+C3+eXFq+BkBh7B+xaDwPRPRde0yPqgZzMjFsaJiEIahuQESm6JKHpLpA0hQ4
fOD1kl0NTedRuVR9zUeDuTDCtA/aiRtUteZ41xfdJo40JBQZBcmGubQf5gErzmSn
Y/T+/PSVZM9uqpUoxyRaliClgAY7asvJGSY8UO6OAb/QNc/lH5Jc90vwUg97SObg
+QeBPdQLdiGibuzPstT+YWJ/E3/3mSWTCorEtTAtPmkm8GYNfLazdCOyoTVwQWIm
10/HAZurNXHTgp9kdNhLug==
`protect END_PROTECTED
