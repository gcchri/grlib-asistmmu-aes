`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KW3Skq6Tnl2FE40vTdu5fn6sRYwUoFnV1w28b6T0e3SJ62X0C2g5SepGRntO35Kc
8Autmlxz3jfFJgjcXSWcSNOa2FjIRAHhUPpq9mtwMjZbuyDPab4jcUEOiWUfnkCk
2CjPsAcinkcXH0IUp0ZCBmbs8Gs7e3p+CzialGUMqtcfkMpxeppFxV1qdy0nMC4S
YfoxqxyEJSNVDlMhRZof7lrq4/1jhord9fdCOknlbOZUAKksOteT6LusNtC+2ch+
aqTSMb4MhXM7R5vqu+mubh0K8iIu7ylc2/im3PnaMzJu2RYuKqlYp26WJOfSlBYE
GT5GYaWJIz3d/LWe5dgkbmGrwzJmpI+p8U9k5YIB22jhvIwNjdz8yEllcHB+V5mN
57Vz1mg/rD2kMlMimkzr3tBoNUIhVV1cLHIoVUUOmgjBlWoR687v4F/Bx9qez0k5
zTHqFjBrXzDB0jRc0AyUaVWEZ8OjINn5g1KzcJuAstymwxx1qRhjQ1/+1zdcC7nU
4ENsrFiTFYSlaEoGxj7+MLeGFh8i81/ywx7W2bKS2xnwAiJymSpnboie/KtJu/nU
4QgXfoC5t+jGwv3WVUvyZFBox7//mu44I4ex9itgB+JDhydTut6w04fzkW1HuHPS
YAI2ECrpjOqclc4pfUxVJ5sSY0NbXpBfBJfufF572FTv1dZGhSsA9m7avfYvzov5
gDzlV1eajxU5YbBE9GIlRh8WXbdGtnf4uXsmao9tsE+TfCbeN5AWHL6lqjeWCe8b
TwX7yhF0Zu+wngV3bEFSxvx3lYxeuV+upr4rcKyvzLO53Cu8mUUuhJXGvYSBajGs
61gU4azzJG5zI56/ITZRJ8XltW+RD5W2CqsRH0jXV4CP6VEJMRkrSiXvuzMoTTgQ
zmx42u7P102GU/pw9uwxAXZr3c8SZValGQAbp1sH8xK3dYhFghI8jZFYscdky+ck
F+00MCQ+1G7rj0lQi7N+32C/cAqvMfOHr+ti7x678pOYDY2XpOodYNmUKgpF+54e
3nRmsV/aak8tIDu2/4oDIHisT4HIJJX4EbK80kuachBrbqTaQP24Sx9HfXyDnK/o
hzonSsJ1LP0G9QDfzjnc9jxES7FM7altV1+V4Rktbxrzvo6y1h1/7iraCTe5touV
Fp8Q8oNeDItmP7WIob0T1eRKqvgBktYWgtqT+O7I1JmTyC6xPvnozNpbjWv15jLB
gq4HNE//GPjCqgbHEPM5SJsN6IfyK3TG+Ta5CLJRTyMTRQFr6md3bOjg/9zL2trB
3/H++VNNvcqObtnRqkIl4U0ILVccPDH/vpghQF42d6NLUvwxStGnpTUYnh/1lhQz
W8RyuZm40fbiZhdgM/M86m4wVieRK301wY0PdK+ESuZiq7/tSnpNDHDh92W2FMHf
whRkAPvlIkIdV/DKYfE0v4YS4vidNA5JymHojcTUt3YJkah4YmqpHmXYHiVtDoEu
`protect END_PROTECTED
