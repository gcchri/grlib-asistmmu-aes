`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJWH9J6Rh2qBSsOn+ey+PwZaUC36mpQeI3YhBOnn20QG3EFFt40txbA9rYkg8Egh
5/ZUrHWzzo4yah/XbW8snLZNOdbw8+T3DtFKkWn8f+6TUZRhXYkW4MXMwGmaS40A
gDgozATlF571T1S7lUrzeKOy9QBgMqQkRwF2/V9z9i7HGXxWzY/aloMtLbsSaMvx
v5FOK0+C3Mji43wYknU75y4+LohW7unaTj9EKcGzK/eCTcT+0lFyNzDHh6akxLxy
GqfYN6fsj5Iz91igPq+aCxvzbAuHAISkPAjxHAtfvFUy6hy6sh1kLcnAVkm6cx+w
1x6XOw8IY3ln0RIE5vn5B9yztSl8Efr8DIKgsP2hzS1WrDs1YvTi9y5e8JdHKHwP
gmj1mUyWl43SabVKcGBXji1MsNBqC+2Ya6gWr2wEbIc4MLK5TYY7/K5k4J69OQSW
/443nhgPrdHaJOksEvwgk6nztzBocIw/hbPz3wo90wfqSQwcGHl1/hxu8xCjkPsL
`protect END_PROTECTED
