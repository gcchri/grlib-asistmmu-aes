`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gIsR20B+DU1ZayHm1Jg06MJU3Z6cspnRmrE5Bh2Z+u8UOGm36mFIeFlRlG8gtOXK
R4SaJ8pmJd8yEZHCVOFZOJgHTkIBAOc2dnpWk0dpXngjIYfV3BT9CPvY7IsWmimv
SkTjcWL26wZ7RViCi5+XS7gs4Aj3xWnbFgDLoTU41hQ6an1SRDZXMxCkNy902dV7
g8IorsoU3z0k4+tZoQytPmPyF4cRvRf+6T0wawoh5BiLlWSDKETFY28liyNslcMr
w8rDuwzY5TjDCMGn4o3BmeAZd7v1jByA8XEBwp2I+vihQQ2+CckkpVgeV2KvC8R2
doJNA4eaF/Xr7shbEo3u9hRtDuRH4cFq0+6FxMx/o2cYqLj+r8fsJqDFiIp64i7h
v4fahZkIjGRsj8j6E5E0nA7JyaiymUXc8I02pnwSIsUvs+1oy26dL4vHgnSq04TI
MjGk2DaukebvAWdEwFFnB18jzHwMEOa53i67njdxVXmBGTpsuWQrHt0XsQOHzYY1
LYtdt2Mp/quaVt1ENRwr695dnXkrjKo7aVTO7pM1gaIP7EOX7svu970coY4CfoJK
+DVW3OyiwBNROUUFX8QObmEIyeP4ZMzIkRSNDy4h/TX9NHA1ZCNCnstoUNoFfuse
vlwRwOpr9yH+3xyJPL2/T8Bj+1SU/Yyv3SBVeSHNUJtkkej8FRY+vYPeEeVvZYfI
ICYfKlvK7hknptQeBgZ7I74SXcOmJu7lHOuPFKBy6WLm/kx/anO6GzEN80jXBS7f
moWZYuSqar+D3UKHY0WLgjkFLNigykklHrcA1uwxA0jbbiQ2FB73wmfoOpwkF4s0
rtPlOfi+dMf2LW4KI4SyzV6mO8J2Y0xuBq0bylRzQa7vBtUE1Ci7RVzzKnCatjfT
pSIg1X5ZsqST0cVDkAOxem6Y5vZyWVE9o0hJeshGXenMdGgxcSBlKIHh6WdGI+Rr
Wxx+UXsWd5STQOVkslLmMbVFZEf14XgdEes3RifyGZbgE1EZy/Blqml80yup97LB
EWK0Q7AvwB92N7xP3RRGKjA7q6f2i502Gc7Cn6DbFmi4tDfmOo7lQKw8ydVsdSuj
NUJw1OQwew4cl44elKjAvuObwMEVvGgRpImxSgmsf8ztxe3098bbIKN4IESujTEH
24RGoJLz3dfqCYjuK8Rn9oFaP7UCXFv258iLn1I1zghuXppJf8fq49fJ5f3qwjUa
QO2LaeJ5mwzqR7kCoukrIwjiHbhjTGuZhK5EXQgjO8YA0ioMl5oedmHYqoxICRaz
K5/38onw/vWP409YuB+QPH28iPF/UAb0pJ9cH9GBhkSJL3Unu8BHZWgxsXyR/Qk2
Kt/d0cb6xMk4wFR3KEl3q8PNcA/IVVnRKnMyBWcpfLYSZQebMFNKP/oV8Y6JydB6
Y480zpQym6S+Ge/WhELLXO90QpMgkMnwrUPXL2LhCnaPIKs6ohhVmKJMF3LHWHQR
TmkW6hnFjLJEjZqxjizHH6jCQrBgwExl1PxPajxSNMw6YZ2CGUMW2jn9R5eBJwwE
OmvIvUaOWPwwOwJGNOv1+Hksdv2UHmN8yng4HsBmKSArbeXkC8UmiigsUgkpRrIt
2J+aUQYPc3kXj4K42YFuj2OZsNAI8I69DMP08JPe0TOZO5pkL+AuZK10FYCYvm/A
GpXlTS9Nj0Dw2pYL66NF8DEW0QL7np9kDHIe9tmxx7AETOl0MOoPG4lkTTkJFh+n
gu4e43zgzKIKGyPh89DMxrnVCHaTSbajm8DY2U1P9m43RB0Sss/hSuaQFFXOhQaH
y6tNqXqcxzmZdjPQDbty+lU8j2h9Wx+V+zN0Ou8JRpG8Ug4SzQD/NBLCh6fAbZ5I
nj8d/mCDjCXAxZBmhjdOhFk42pf2vbPdaW7fXMAYJJBaSVjG/wnmqUmBUgEePzHJ
zl0jJ9jdCfMH6UshXCTIUyKOC+urMMQ9m3sQkXgcpz8WOVid3QWkFo86VdyW/aT9
rfEIyDtjidPnPvolcWLA5dRNrgOy67lIYpBeTwVslgkPiyCD4jhOosOZRm6c0MPo
cw0AVimRmJhNs49AmMPjUoAR/Vw9/2BylZWbebB9LsKJ8ufOqC3/+NriRM/pgbAC
FlCKmubw12l5dA3KMnshfMlx+ytrc06NQ8TLJnaSp12Ta2/EHXLAliLyRQ3vG3sI
GlOwRVpYDIKJ5J7SEfCWKQoVk1tyuUyQ8xJCNmEvKDnEbWw+XV2rU91QGeHivYtc
dVKiPOjF94N2aNywdjCOucim3u3f3ME5GN4+zpFhvlIz1jJtnUTASErEQj1qNUwR
RgceDLUzq/ukB0vrWW4UoKZwy7FqtCDsk/2IuARMhCpAFrRe7QzFSo0SK3LLPBe5
NhESUoWtmW5GhgdZAkydrBc6dvrXaNaweNZ1+FGH7OzPzYAXoeZPb30BEti6C6Uz
v1yYbEoTXTWXzZ9HQwu5Gy7InDg5H8c7/qpgSxNMyXy23iLlzrdsv1LpwUNdbMFR
MmELZWcf91vZ7C9YP7VNfWEFVM3bBSyouL+pfxUvIq9oJsh1FYRfSNCdvUTosLz6
m1ZWzOTT8BReTMKhEnT7pUdntq08Y25czYdZ6qkMtBNim3Cvh4p1DptJ6Ic8lpUM
eufaM1NBgBh7+dDxIUuKDQ8m16wsJJj0sNYm97qTk5dzQlAV4syQxA+87lepqMnV
0hT3vT7gac8sdFbdMZ5WtST059g6cDpc36+XEVHe2Lk=
`protect END_PROTECTED
