`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TluGqinut+ydSzrsyuLQ4jHu9sX4aZnVWVfIm9xbQvJSTDBsKTyfHi0cJpKYFSBM
dfupJDbNv41ANnIK5mBLmmK8znSYb3ybLp3c0IT1D1DCsl5NbmIzwlN93P7BFaWQ
TyIUodwDZrkiRNZbN0qymjGc43Q1GvcF/v3alsQqjnlElRvivMnM4U8qb9T7G74f
BTDCA7NBmO3wMjj1rCoOJB6liGxixqQZIPKu9SOXZ4JQTFhvoUb+Ttf/SzTceiKl
in74/bqnJhdZq8BI+IjmrrOW96cgVZS77IvJBndUDxpSbUM2SEOYl2vIsdRe+MD7
jRxWSy4V+oSfhh7lOCP206ikg908ST7cC5em8nAuryXG/ie5VCZGSPMCUfePXkdR
16G3VHSYwA2NPhQuPsNlWibaE4jCuICdH8Zd/zKjR/rZkMazApjVuZGO5U5YPjho
mnZaxeVIUYXxdSbmGMuq3SfmoP2/bjsgsC8VsX8EXpMIN/jvRlDs9uozXtJC+Q5Z
`protect END_PROTECTED
