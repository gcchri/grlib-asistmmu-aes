`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7z0LoQW63paeKPUl0XZwlOrw4c3quIeJJmmQRMzI24ExzdCafWkheS3+WHK0fHOy
5XxKmNNjeAJ7VIqodiPn17S/yQuhtSx7rzHAVsinl1g/yBRprXvASLWX8xh65u4a
7TB6WGLrUIlDNYc3hQeAzN7BfuJ4rWR2dK8/YBhE5aeSGzlJV6965lmagbZgKqOI
qRvClg1IO9jCFwj0LrpdjdZUrXJPek0Fk6L/xxwJlT/BypVkt7Ci9WJUJDvqjf+i
thrVBehSmKXfsXAZzzVzjxwlf+uozW9QTlwIQoDlOm4pLw0Kiej1NW8X/qrc4gaG
NEdZFGPsAn8Tf7jPtOVXiblCe3eW6qOCko1OMDGr+KcMiFlpsoA1+gR9PWR8jsH/
xoZQ/A2qH3QrjTCUs0JABee6b9j+dCYKjD0DNkmfO4CVHbrVjq40G/65/oivK8OA
WQIbaKE06NRz/0Y6Rty3cCCXKpet4MLCzaAKLhVuizW0zUbhZ+I4DB7aJ+7umxrs
tadTm2rmvaeuutQIrXGwXszk8pUoCXt6XCoOgrF46awqWe9xO7qv0zFs58HvdJLT
vxjmgTbs8VOklW/5v0zzumUi0Ce88G06ztPdt1su2+OC7l/shdb7gEhG7dHbMKeR
FtY1mrYv6WTboAgqrT6OLUx78HE0XuHZHn/jNG4EIATpGuZulf1ilrzslGC4ky3v
FRinZcEok5MeWlNkEWPMiO2OwDeQwnXoR8Oyc9cdE/rxEmGhOq5ys1EytygI1YBh
od1GtDNI+Md10oBO/2GbGJwxhhlT35cZ9Ay7ZTsJNw+VxntXnzqQMoR+yGW7ocsQ
`protect END_PROTECTED
