`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SGxZ0b1tVD0YsiZ7wBkKel/UrbijuOrcB8fwm2ECUlRpzNcvo1hjLgBrcLKXfIvQ
4Nd5cuzzIsih6Uj+jmjitZ+JmP6Q67/b9QgCQOT9ySC8PW/ALalTE5cKomHYHi19
Ib7ngahXsz+DqXhiu5UHiecC0lRIB0TrUPh1HkeaRVtM9yXS8jT5JJMbhksXA9r/
JUkspbv6vQAKJgvkzeVO2lVJvw7ouCtuKyPQ52nGDvESbTX9QF1QplKXBAmJ6JyK
p5RPFHOZFmjzcFu+jTt3XiaOWdb0UTJR6id0P9ZqiIezA9WEXdVfnY2+ojkN0piH
8n/jEOiyMiO2TLRUgdZCMA3Pef9zr12uszbL5Z2EDBa63zANT5iXSGupJ21sgeQ0
6t3nKXsz8q4ZZTI+nbehO9bdL8kr35CJCkmPANxbA6YjwNt6z6Cit39OmDDAL1jM
XN5hUEdmK2FXVdymnMdaVb0ohk6vVm9i4GnoYfBeilnkC4kenUgTtwZFIo8vCVLP
vTsM3/k/7qKc6iGBzqHWUz8hM+tiRn1B3K2QgIKUE3D0s6WslBbe6UNkv2txAGPY
/T5Dg03caKwqpN/MjZZPCimwOerx5kOIWEqxBUBh2JL8WfwhENSiMiXbJVzmcyTN
Rj7Q/3JnjbkDEq1ko7Bt1PRQHU5T2IsJr/MDhczGUi/fqsxDQkD47TKo2lSgxIfS
Z8a0HNbMe7MPP1Tk6P7KYMoLwXgnvMISdtrCsrPHbHyC8HK0tCXizj096g59I8qC
3a4d9MScMLzNp6fC4bY2Ns5oPztwixMID580hJkByjDgQRGwPMeJ+OwEXyTmIz8V
WcR8gBYrWUssgLGo853rF/VQ5IDWUUOd7LnzyfY++SzVcxolZ0G9A+AftaGuxm0i
dFXjttdsKbt7VJswIanxfdu00LA376wJGvuO+rhHwaGfwoO9Rry5fWx6viKTClaL
Ac1FnoxhNHQZrkbJYtR2XS5X2Q2tG9FJdt2RU4EYgpZNr7y7/1YzNwFoSeJg/ArI
6okCd2/IywY1czGQ0mZJRPVJ0wDyARcIb2W9Diu4pp2SnOHaHe6R9VySxPW69oN+
k6YmITFjRUt+O+kIyuu6fRWosfsAO0r9aiwPaRoCQD0hSzXlV7LPEePp2YDQN5Yr
4Jf5lkRKSLPbphildpaDhDz4A2+s+Hjl3D+sHKiZENHDw5c3c0IqZYm8hiF4uiyy
IWsyuwuiqRbgYUL7eEGYqdUeJ0F6Dww1nfrME0IWqHv3PjDRIWsqJLS1p81hVols
q9owpZl9Phdi8EY1f72fH584KguSVmfFqt65xIZonZwnxJOQSqgiGzLN06wPMqeF
cpkQadFUsXWR9ydaD5plHxVH+cvzeh20JZ3XMIcR5CHbDlcvsI1C7/CRnFHkizbr
/iVY9md9T70IpCTTuvJCuuiw5rAdq8lsTwfCzvVUbjKZk9Cq7qvKzHFDfyvlmSLf
JiKLdhOK0SV1FXeaR8WkaulWKKB14n/OysVClZOKo17uHkifyFUhWTt6qkwjLUkY
/yFb0An+P8mmJ/FCDCMuv9gwLznYGEew8HA71/tVj5cz4rf3vuNqL8tycKDC+NsN
S8iesf91DzojU1u9q74eeF4LylEtcuZOi1EzbaCKWdiGVqevVhDGqH3ELZ098n3l
+RPA+a9wn//evalS3iFHPmP2bFW4n+lAOCTWa14ftLY+F0k2XjwYb5wp2CyJE2uX
m4bAdPMolrRssvd4MkaaGa1cyyBUPkpxeXuDfL6wTlN9+OUHeb1H/kmBWSuVxctw
RRKFiV6ouMtL3M5wiRvr3SgQfmilGQaWTt+35se62RNZMKdzo7iF46DwVbECdpet
OdrWa9OIQViNLa+byAYjTfHhUQbfigbAJmAXkRlmzdPB4ma2MfFpHd7NncGE+CO2
YDa/ManrT9j//LqbACCbYg8dJtKjdcGhmqq/orF+p4DlJMJu9hHMoqtrmIKW9H89
GzC/pOCnW+Ja2s08RcvXNVgwKFONpEx3mszK1hgE9Jzj1nDoSSW8hP/WKeJwUTs3
inBUFJxB3dl4yGSAglxev8n/vVdI0AWNUYJm5wX0bOyfdDgFFNhsjLKWKQnf5RvL
GA3BvkRvOOBaLqpKY2cYjXY+pboje4A0LVe6ykK7RTd7VnZvg1BXDB8fK7N65kgm
uuKqOAIy1rrx7DQCnoPngs8Qp1PMhnsRaRwxGzkUmzb2nexRkWedXEtai0J+tDc+
v3c9j/YRyK3VaDnjWdmveWR2qlFVeKxBGjWP026+xy0mPVUhTFGWw2ArgOJQuoXk
`protect END_PROTECTED
