`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJuG8C8STgMuKHmCcvtu8Nc2n8GfZS4LMBjIHiTnQbBMuH2E7fvb83Xt6Saw1mC3
ASD4LmGRI6Fnd3U+E+VuzeYiU4MMbVPO1tXC+Ws6cSyMJT6FKm6I5cCXsgutIMLR
P/NETxhRxsSuLd/KgQjBMztrIHzNqVJtjn+C/YRp3gqiYMOuRL3RgkeLPCl5/GcN
F1aeMiLuOTC1h3Rcydsft5ykUcrvF1givI8sa0evXpEdjMJJdzPi+UgKpq5A3Zsp
rHfagpL4R96hFDuXa84hTAEgeoD5FR/+j5OChDcLwaiQCzrADTxvC9XJ8lvgRt8/
6TKOq6r1NLggQHZsqUy6MMpSCo3oXkGasmV2uIRpxz9/J/9foAH292zDQsU9jtZC
M65vLhUCBrwlbrejUSKXgP9SPRsSqGIWjyhoC6cn6k7N4LF8MleVLHqOIdYJM/RG
`protect END_PROTECTED
