`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMkg1nFZ39BxaQANkZokvKXb3WE8jRKRr9+PX60cEktpqgvER6CYEfRG9WpD31VX
UMvuZHFo1Jy7fwlxgRwyHj2vRvcQaWo1vXN42Aq2B5/8fiLbx3GYkJtND5DVSvWl
aejGvH/RZ9b/diMEKskk/Q23nnuEab3gAALDJRVIfaloSwaiJg3knCeWq3QB0hwL
Z9fNrevkpjNC8BFmWG5Au/V62qGZYjUTatl1abPz903zWx7K8xXEfEpwPcRrBhj9
2Xd0u7Kj3cgAbUOZ6tu5wdLWGkMNtA7I5TQrCkRaIqEX4LW04qDaAfwjn4Ii1FwO
PbqjFEualm2pWvgbTw40ky+0XVmOAe7JUZ97pAn3QF1/BSPcux0+rGoMvizG3rV9
IMi0fVvYyzbNBnUjz9ilodveZgWvtMpuJLbA3AN+o+86xnTjShYfdR9LqEbkQJxS
S9iTMm8qMlOcE8NNtoHe3heorZHGXAuVo8gK48g5PcX5ygKlQg6MYRj+1SAsX06x
5qOqiekQ5UQyIB2exMCfngHb7AGEnQSBXxWxgvDSLs6XKgLYPlHaKPUCKPZagUIb
6GjokT8NO9VvohYXX1hHaRrhnKGD23nm19yXExdPXMk=
`protect END_PROTECTED
