`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0iZOWIU4Ge3oD6v2xUtwY8J2Ff5QI8BsdpUheoO6+vDtnqLozaWVrmDzCrK9dzw5
+WTIhXqxe+0tfSZFP/Ar8f34Lgat4ITYfXcB+MttKNfb+FRdRBJlzPWdprkN6zIO
D7pGYE4rRizaSmsBnszbUQL9NeEzhFxgNWtNDMstlRcyG01g4/5FA8ZSqJb+l1yk
OasWXazzAY4t9buIjw1COOtYh6wR5b5QPHWqw2EcWkYSpkM+CZ6dwbVlBsm7rqT/
6hqmJwA+UdbUljn1FuG7/b5we/5BjBu0XRM8kZyjyrRzoyfqpdhQmRL5JA7C5YBy
OEyfdvZKUjbODptI+sEXC+UnlIvJJUBITuCcP9JyAGagsOXxR8pZHa4SBNrWDD1/
BXhLGe4RSUj5s2i2ofLAMp2KGRphIVwwRQ9paEoYm6JBN8C2RB4gzS1sN1GtDHVJ
IVDzh9BTR8euzSpChIb+vByfRlhjIuqr98t/u269xXUPDAY4Jm+Bhukac7S5IQiW
BQaFO9+0H6Zgl18GMeo7OYaTmPWd0kTH2l7NisxBPvMz/T/vv2UmfOHakFq5MnVW
n89TbhL0vn7O9YbPGAYyMejxoUfR58KPHb20J8dO/Fw=
`protect END_PROTECTED
