`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eUXJHopKyPAmUiEjgZK9NjCmJYKlwUMgGPrR6PLYmkVEGAKw0VxW2xblZgjAP5Tl
jhQT5d40yoBeTVuLQQMKLjU3SEa9LRzH5VC2P6HTJOuE65ytufqp0ygtmzgyTVdW
5uiQ9mrhuRqA7RL+AG5N7sX9twiNGJM+t69A9k5LT7aA2bM8775ANh3hwlMMQXTU
4i3ZqrOkxP8IDx2SLmyWwsBjwQNpeUN6jQrPJ4bHBmq17Uf42Qz81yjQp2uH6XND
qaJB47MWcSdeAeZk0PC5Cji4WNE1A8ldP4xF/Lh+O6dHb6roy4mVGaGRLDQdWJdB
DIqCwMVnhAxQu4wTPduglQ==
`protect END_PROTECTED
