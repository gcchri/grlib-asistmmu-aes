`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2i2tgewrs8j7xXamnaKU6JXzDhD4Fk8reuSJS8VK5qLtd5CC08Ut+su8oHWsIMzp
VQAYPQ5C5C92cikuqvmNvRKC584T2ZsFM8KXQReXaBHX/MmHQNEoyqVYA9FzaSS5
1i2T8cgJjejDveAIq40+jgxH2bYrNHxO/Owtb7AjflIgx1gqs21hKAiR0XLg5W4T
Y68Yiu6qTvU9bvTZanzyORThrgNyF+RA2vCAwBz+aDebYxumk4aHmh48n+k01+7s
A9zNOTyxZ+Jp6tx9Dd2TekrlneJSwMj2COL1wwgNCTBIj6Qo5D4MRzLBvWv+XWh3
zuUBY4IE0KuSf/goLGwrGg==
`protect END_PROTECTED
