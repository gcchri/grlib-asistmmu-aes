`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
87yx4dzag3uOHAvMw35oIabrLZ6FZQpTde+PBXrLewpt1uWRbFrvulgBXZT0DVHl
IyoO52X0Mv1QqHPznHoqurJnpLy60JTyEHm7Sv7n35kcR5JzZRyGQCUQcJzxG21C
g19QOR0WnBlwTb+NJsaYiW1zbITlgYGhdZuEPyIVv+dt3pvXi1vU07BsKxTYgl3t
ue3Ck1gjdCtquBEsLKb/NUD2WoZc0KNSeqkjm4cetToTcczQoD7tfDSP4ug2jbR3
eBYNuQnjFYPpriiD2qTum9Mvk6rKcG97CO3qTdAVatx7TfpkfTVLz1jpttuwzWxi
vkIrTNCzhIUYMwj5yJWnnTCho2qLb2FCSGGFhG7Xpzbh6I2d6beYyndvOJuoDMGV
MJGN6qvhA0/8XsKpsLM5S+v3o5jzmzF9/Qcgg5PdCR3sj5rsYq+Hv5f/qY0lhMKD
ptr+ePkC0ykJVSw50LpZ5V54IDviwwE8bjwHVs7vktnABu+qCRtwT9raGKoG6GWZ
/p1T/Y9Ydfo2Z7twR8e4Rjxj4Bxrj35t6b6dhCfPSDpJpCSRFZORz61R4higms+j
B731GpV1mvq5iNfvBGJ77fDHbMBVw8vhfdQsqKfttnvp9Y9YHTuEhNdOBSd+sHi3
zt4qXkZbe72cmrdAKnUUnorJzGjECvMUpZ+qbns1Wg78VySSQddzcfWhYbCTA0RJ
1rXm27JZp+cdKYdB0ZwE1g==
`protect END_PROTECTED
