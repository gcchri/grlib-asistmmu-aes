`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OOMPjTeX8B9twvXLZYxTUlV0LqcFweZqASUa1r7rujV9YgHuNptK8KgUmMOVZ4aV
vMI0KLdxYJ+ym8RskuxeACpmz57WTvfBGhjWXMwSCOltRrjZXbBAnW/y8I+JYmci
QprJcbPICPLA0UpnC9N2UCWkh+ZVHzba0iZbDBZFPrQUcWA9vgY6zj/f7q5kurgt
DKZq2K1JNuA1Ff2MmCbZlRgpltHGuw8u29/utHrvd64em68wqQGoR0jWg19X9DBj
aCA7FNlR+Xy71VIIfvyGQA==
`protect END_PROTECTED
