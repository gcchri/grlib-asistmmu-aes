`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0LLw4kVQ9sTZ7miKwsZdPyppwxpEGWYzvU2nuGCxy4uzTTSn0QEweeu2R5LIu7wx
GnAD3p5Q6n2ndEqvdFD+TP/sq/hoCy/rHpPCRxfkNkCNH/rOo9PAtY2cvI7XDqex
6ysPAz0U+atOqCmnwzr4gQGD0TEyOwW5Fq+llxJAbBx++tJf4c0TeqSITpmq7DXa
Jv7l2VWPb5q7S+Qp3wYiEB+zH8pRZqv0oq3KLO9/w5ZlH4/qqbBjTL9sSX3C39Sq
zczLVYGUAqVNr9shtPL7mjyCf3HfKIqM3pmrDwdkETkiREsBw2c6ki7lpXsQwcYY
kejmjvE8J72tR2YPOOhDoDecmNhN5unQUz3YAc5VKbzKaJKkr+hYE0VyeDOnP5tA
BeVWuTtNZSDdTopw1AyZc1XNNk8mVi0qRKJN36gc95dsZJRspl2vqqdGNP3jvHcF
1OWt3nQ6QUG3u4GZGy0L4dpqQBJFV8GNA1uVZ3jOyttg5OcgQFtn06TSop8pbpbs
iHIPkkYSRPtAdYO513scdJ1KDO98HohzK4QKbzYlLtC7rYo4UG9jG2Ad6s9dLJE7
vQfta9YV/UG3jDClv4tL/sA8b9mXvFOhaIZkYHT9uqRYM9gJJ67jnrnzz1/5kl3X
DsBKyi+TB8Gsm3zqZn892YEj/qaAJBQLzYkcSNsPLE7HlAp+4R57AeAb5lgRb/A3
Zwt5dnDbuXU8exL6to9pbLWoUuypdkklSQzVHB+rOzZTKtvhJtOqLB6dnjcOphvp
/FTpphdSUmKgwMqBrEP0eW7Vn+Q7bBrBxRexEtaBZfIDSLjhoLp8HYvoyw8y0WvO
629FVBx5UmJ5nDUfkNMUrnh1H1akbS1GuyCbcjEXURPDpi3MUFtKNqLFTG4vXk1x
tVsR+OUalp/VJ/v0k4u9AYNnFwrEo+MUM8/vc4PlaqNMktQIcgCOBF8anIjF2N93
MdRTvGXsAJIv4d4oiPHom+6DDRPIYKKPctdvQgv1TiB4W2GqOzBVugyOD5IXCiPz
PMMojZ82SLV1YDIT0Gc4wv3dtOT1PVV0l0jUdJuhq9D3ZKoxdSj4ASjJHcheY0Ib
5uTWA92NBGBTOtERJneR9N5qnjJoRCU0cRCsW4WNv57SRLTeLCYi0KWdbc+MYDz9
7Aeme2NitVKiHtEerE7LHQ==
`protect END_PROTECTED
