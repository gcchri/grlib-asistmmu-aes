`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/rQIEkRiqcx+xBNhCqc4wirY/kc/bV6AJO1cBQGaVMd2afIMs/AxmO0NRh/3rKq
14IddCCowHANqPf13gMVsZU1ujI4NkWnIQf2JrWh++lpX7/aD9L4cjdldDjga1UL
LZl07hLBvcKUCJKDipuSzZBF0dOlWDTwQqiutMwipsH54Vx6ZexMg5PexlY0jogr
rTCEPL0jsLxeAaY0Ay42zcQuUNbdlrlImVr3+R5q/mvChGdhH58oL70qki7Dnkg3
+Y0cmBDUaGedTe8J+2MItX1fF3uvGoNLdsxvLNIe22QcVhqSbbylBeh6LvE6HbLq
LuxF8/txkO46shVmE58ic68HorFnTWbN1dtr7yaYXi4=
`protect END_PROTECTED
