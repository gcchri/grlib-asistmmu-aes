`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbRKpLaHYqdvbJXLqvjzf+sYmcMt9C6YFJI/R0gQuAa09zSbh76V834NK9/vZjo1
07EUG5C6pRxDm+k/w0zfSFEtypYwDPleLoAoCKuwkKo2zz16WX7nO0vWeJGZFO/h
/L1njCPRw0gRufhXgsee3dn+aik4Iwt7yXnUHrnz7vcILrBr+Ncw7Xue+ieUsIaU
xMrlz5y/cGu9V4j7ueeh6/JZctO5bLecsosuTNHJzM+7J+2jkYVmF1dMSTLjuDpq
/tp9PtbJKi3Fiy8gmBjl14mdzcvNd0HW7WLGpcla0aocIMN5TsKAeSddq+Jl63Wq
ZVqCqBdKyQrh1x5ji4Q9p+riioBmK4QUpjHvutFfc2udlpgy+mgV5Oc3TTkOArRl
SSHVVW4MP2/0x4H06uHspDRvuE/k83XyUKMJl8JuO1RYS/HULZw2XLIZwkncOUY8
JdxUkGnMzTfzKUPKteV/bNCii7BTxS9lEegt3pjd08YW7eL38NjGlEdqEYrk680F
O6ZmEuir67w/jkl260T8tYw3lpw3aOGDFW5LEOu0Eo48fcQcX/UwYjLvT4iVFPu3
c/6GVUqgTmVpVBqDsxH+Y8YYcbceo8w24PaYfEvuar9XiUxbvJnCGyCHF5ot4Wik
IpKNJheEesV8bK0G9eu8k/OjXR7FCND6JICpY4wqO8ZIkZsqF8RW1EMRfybGE846
2tkPjJig2wl2FIO7ATVhuyuwEDcPNol2kwql280tYw/n+u40bZ3fuLXeT2sMuG5o
3HX2t913afXCsJtVY2t5u8dRbI7MHN7bYfX28eZ/m/LWXir0Vqu2ihRdb/r7Pbyt
mn+rLKCQ+iWK2+/P8k0ELUZbwGqy0AAUbabJMUzMW4u2LHCo5vQoEOxHQXCrMSt3
FvOpRaJ2B3dcvQZVdOcByQ+tiLkfIS1tsPtSH0j01wU31NIiJ+f9lPnOrZu/VqCt
6DFH+dzQKL7xx9HgA5o0fwpVV2a5ZR3xEuqDyV8iY95SeE16OSb6ucQ5oNuZfeOB
vij+zd/wnneubDOxCiMWXg==
`protect END_PROTECTED
