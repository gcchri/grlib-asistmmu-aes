`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nbd7dV9aY1BaW4BkMVwb6x9/XL29S8wetdC2S3mB/GX7GANG0xgYL5oTW+oapoP1
c5Eii7ghvTjNOm0se9tVToURoOmiZfPm75TYJRpj6KfufXLVYKVYTkZ9cgGiI7rZ
fcJqjXDYEMDc2tS7gC8YrloD8v2KgMn3prPiisUTRtcF5nGXOta8bExV1RdWWv3O
UlmViJAuiz0hzc9fbI1UQ1+jgW5pnugnZJzypV31kY0qY0WPx3MjsVAy9RsLfiUf
yGo+UQxKLUVIzltQv5KrI0fUbC5XVLbrF+l3gUg43mn+RsD7RvY4v4l6ua66T2c8
4YzlLcVMOZnuye1ft/+JBKRKWsjhXB8v1ZJpXW9M0Gjjy0XmNT/oxk9CO+8cFGE/
Od01cBPDZE29ARAL9Wri21bhxpNtD8pa2kBoRD4AgyLU5QWtMzjgdbL6D0P6Wwvw
iCZPislYrj9eTD5Op4rqjA==
`protect END_PROTECTED
