`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8MilKy+w2DFuXCr/xm6R5gT5iLNizBh5HZBdC9e4qGy5B4JF3LTEIlOSy7jPdUR
7ha49t0NQt/tJOf8CGDDzqEUmvh8RzcQDjBjGcelxVfOBtgpa4ypKyo1LRChogQf
Q0fDnHVjNTobEXNnmKyZ+tWxGDJIc8xrG42WQg1TXydMf6N7gtMYU00Iqc1XjxfD
MOSuwfDfrhOBxwpa/HNuVqY7ptzeGz9UYCLQhLKnPLmfFDpqwh7BwXDNxKZdvtyk
Mr5mLcIuatmYn/xICwmL2UGlVZqHtucXvAOzmu7Y+dz1dwD3XvWNWvpeorzxsCiZ
NgwKg+Kb8nLAEDf5LDJWDrHnFqN702H5lN2jyXCdhOObbZzX8OecGThoaPWDnrGY
BBtgO+UF4+11N4zNywnNCHCxDSTdAcaL6jZlN3zFaCctDxvfML7X1ElJJsdjRXcl
LW4Dx2R0cGsSh4HDxQfK8uKly4ZCm5DZZe60LWPsHd+OKf62zKTqNhOTgkCb5P8R
Q4noD7k+EmdabagLzZGYoqRrNEnCeOqzThcKa7gJFEIa97/PZ5Q8DP79Ta8h9S97
pjzxhnTg/jOkSVVk0cx1zPfARBqxlpKhxv8bJ7iJdBzso7K4DUrvK2zH3EYq0qhJ
xU2kg97Wpr5vZCm+P+ztMY2kfn8u/ubmSiwBVh13XiakkhwQxqSIUk3MavzdiJAq
lWTF+Ki2xs9o8yhlCnlZwaQO+ThLVGM+RLVKgE563HIxrLgKu9jQli4WVoWXYqqV
FVuCO0FiIG6Zfq7ePQ7a/QCjrzbzrx3zz0AgKsv/RM5/ubVVyBGNzuCg/Go7TCH0
nQumo5Ut3idy9C12t1NP/e5eBdyHZitkdjxekjbUfcnzZ9z0ihpEBt8YxXCazys8
tSUGir7mgzgDegVHAcN6uWxDKOexvlQ36cgb6apxhQ2sY7+HJKZmFCp6I8jaVhN4
MB/IZPq9CmLAdGndu79jEIM59SSNCtAdNL3+Y9XJjX5jWiGLrZsewL/iBZZsmOwl
1BhcpycN0XGD8H3qNp50TgkG9QGzMsyOHirLImtwhkY2MF6i9QkUZ9vhhYAqcjZ0
HCE6NJiASFa/axe98q+WWc8230/HiTTkdrDMSxTW48GlLYVut1RG94yxbi3SObBI
3aMsA0evVOpmn9a6OFPNo2SV/+reSdC0X4uD3LFCkLCOZRHja8E2pVsomKjo77FR
HCDZYL+F1XS4bv0soKo81+iKQJ+by1dBlSr+OQKmGUyBEP6CXCYJwn597aCo0hGF
0V3oWYw1B7+TNL/G69GKm5J5VK7wH+CSUHW4gxMrRHIp9+ySeZeRVOvyE8YAd13+
36Ujw1+MaO1lSfZMaB6njuvRbwqzvErNO0UM0XLtSDgLHt1Ly0n7HNFowR6Jgh43
7H3OuS7jVynKm16nV9EtJnyGh502ipPR5XBBpImrIAJIK81x4Odx4dlSXGRpwhM5
2G3Uz0gLI4tSNqz8i8VMj8AEjtjCpx2m4zwlFIY2QioCsbg8eQCOzBoSdaIsoXZi
eHzF18OHx+/VzNjLp09nCBIducRcitbEzMgX/XCNbXhUCsYDIXPMZLoJod6CffXQ
PsrUqiGjDy0VWJOfP0he9bKfQ9AD4EOrRr50TXBbMk6Zck8r8sNgAZwJkEOiruDv
ZGYa8lGwMKiFSk/isfSLVomE1v3Mqvlv0zKa+R/besTmi6EZlnLkTxKgKm3UVCz5
XqqvQ7P3W5pIGAcGUQc9g1irbQqWlSAa1PY1q63mnnYgTUVlx8vFDEIM046x/By7
MiAqVLyajJpRM1e53DdpeEwvBXuafWOUp/bTX1z38okzQkHSNec7IfaJCRhJ1wKV
f6e8bMnH0Ybr32jGg/uWcaLsp741f0SpinKC05Lad47PVtsJ18EaVEMb2+lSz8Jf
QXnkD2lc+oi5Np5CB5LFFRbI9/JfR5joC9GSQHi/aAbghK0PBJcQFH2ppDQj9sGS
nKCcEaNkA32BIWFeohLMRQ8NDisXBiqeTKaiWhOmVPk3lMwbUjIrhtLhC84Tx7k5
mjnnUoXVnd/G6fKou0hojgFB75CiuObiy2aO+posuWmRWkeWbyJPv3IsXL1VEfx0
0wGWc8JO4aDHFvnqKWPApsV/2lhmDuQ6Et+SXGSQn15G2GeKWT7pI1ux0ZNIntgz
81RxMrp18bf1KG84TL0KRwvDd2fdKjxOX9bS+hoA0QtA7hK2s/OYPjZ+P+cCTKQg
+WHlQf+8zEY0EQvssNYgkoqAnFqns3/KGlSh+Ou/cY4cFJomKIIkEv6Ja1SXdpVp
uUR50+iX48Tx6HSgVy7tqsIGc7wGSnHTjJ/KZXLS/UAyJDy3iR2Em84IxjDzkdMC
0SyYT+PcEVje/VE2FH4hw9KFSg90K54NNLoq5+MIGV1TZNmqxl91VknrRUnG9Gy3
Zp7mJGY8kCTZhNFjQqUM64fs+HdDvgSp+SmYW43zD6YIC1Ivk0spxMTl5xUX6HTa
ykaqzx0ppsC7Axjnm4N51LseMIdgqm2X5ZwBOVOp7LJOxCpxkcvCN4N7CYNaB4Ec
KvIpfoiSUB97HF3BjQ/L2Q==
`protect END_PROTECTED
