`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QVLIw5LyIlkBjqfnX6ZQgDpkfnSTNiGi0EorF4v+JfFkFKY/u0LfGd74H7jhDP9Y
DHSUPHI3YhEbeVYFmYWU0bwc8BRGslpTo9ikQXaY1hpDt6m23EAKxuuhnj8aGfq5
WJ4PXfDLlYTFUjcLuE0TMJzkoe9TqKnw5i1jem+zVFdJLLCy3/lIR4nOrJDNfV7S
G372m4GjMnvUgQve/Fwk+wsfwuCCv8hFXTlrMg8E+LBWMf8LIAuZnqqAYpG6kVWI
b+Tkqyjx/Z1X2yXjz+3TGNOnvzs/dBtZbdfJonxNqjYWFrkQYnbXiwlyUvOJn0RM
wSSWQucVGEHhr416pm0acpXM+IPiinkpm/XvhrQPRe8ka88U4duXhCM9sayHPHac
ZVMnRXiVT6hTdK/lPqYTaCKTpi9kwM2h9by/r9pFdqSnoDzp1o8iCttz6a+Ge0HH
oslFCVpDdrXAsDOSYkv4+48DhRCl4MQjaganBbzayKorLfnkiarhIGJl4x1KsnRK
4uWnUNiG5YEvb4xgu6qme2K8q03XvpDS6dp/VI3HW/FhvI5ZBQyRpTrxfnq0udMq
sfAfndClVoOMIGOjD6Wc3B08KJWQBgCvf3fDSUJAjwsHwYugYzByd9YjLne+Nie4
cUmtvZmpYdd/zLVzACfcwdV4iuHCcJmwpNlv/wE1HcTJ5/nfHrvNecrSM55kQO2C
`protect END_PROTECTED
