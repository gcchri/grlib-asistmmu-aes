`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1kkUr0JxcM6dWQHtcBRbsE+G9tpjPg7+7CxIMRRVd8Fm8aASKyDdPaH84EK1ys+
CFeSDVH7VRvmbCPo6qfztlKsMEye7ky9ULoKrNqc8nDfUk8qpXSO0mEYOOVfaRTv
/a8Z2f+5M8gPE2uHrVzqxm00dpy0kicXMerPZQwe+oPfk/foZIrCi7KUQwT8578D
3dGO/bXXsPttGgJjokv7flkUlLhClv8Ms2P+es7KEZEbDNvZdKJaS/uha6deRdh3
N4bhlE4w3YDQaKEKrrqWoUnN112Ose78R45gPQnuFOYFUWBQkvLIkWUOB6HCJXir
1WGGPkM0qQU22WlW1IyWeSfU6hOi3Ch3B9xmkUWQQxtdxA+3knH4AQnp/dSzxIzc
roR5IhVZSKXPg3i8/8F17Sq2knK9s7T4Arjhmgz0hyciv3qmk0n5a9GHWDl7N3tU
1w4JNfzUSWI9xf7yjnfgJ+cOUkpTLqOtzZMnb2JRVUk=
`protect END_PROTECTED
