`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5iuzRnioWUURjHDbKzkt6CG3UN4gyFwM0DF9iC/zqRzjyMcHpx5IGhwKrcu5ywU
DvWXptJ0YdZl8ryfLkRFDa0S0eWjoRQsTgjJpyBjzkrifgF5IxDS3bsOHQ2MNlwz
Ok808Ite9D07kZu6vV7OjlCm22FuFLszXTZuxWOXlnrZBB2UZL36OPuMl8Jb6unv
/lJs3ma5mr+BIn44t+co4OAUIS7Xp/ZICL4KRIUeYQgqqgS0RU7AKns37wWPUQn6
fakn85nWgnnp+erNm5IAreX6RV8C0wIWxoSrzV/r0TQD6NK+qjYcm5BsHhLsLlSh
CG12KNvwTPf2pAFzjHza8v9FCzCiSOQhDVVKSZZBsvE4lRLEKfEOqOdTtNmkZMJs
GGTmVX7+qoSd/O8SqvH5tUkbSKRAqsdBdffFNIWuTjwSQiV8oT38TlHzQpLyDvDL
mKgYqWAi+M2OL0BZFKXDAQTxO5CuSQ0JoF4iXbSbTzzjBPCPeQgiQ2JUGmCJMeUz
`protect END_PROTECTED
