`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cz4bHMltU3CZ3xr3SS46l17ub4XuPMpkCG68x63HHchr52S/gDCerWRKM/fiZB0m
RKjGKV+gX4qNCk/VP+aVkiktqN11AL28LLuqnU9mkiXPVgEjSCNcOTtQRltZYVFq
inunAera3B60LVGkUqgCuiXLyCq634hytg9G5X+2thCUEkPJIRhbYf6yhOF5N+bI
RJmytyOFidYEcvufYU2zCKHebDmBQQXhFCB0HWaux/B3Mj4UdO1RwpDpDmlQxWMc
eY91siNx+q+VNLsGiqGOpaqz8lFGI0Ayjt1YoawrHKwusLMt9pabkKAGnwynH0Qg
bd1Ji52UGGGjoGF+3hD1Ga0ujOu/xQNt+bvu9sDxSKLQPBZHz6TzTkGpWXJ7Dfza
0tK+W9oA0E7LLAwM5pjgYA==
`protect END_PROTECTED
