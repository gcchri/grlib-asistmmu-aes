`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bG6ZaJUODJ8P65/q1tsXOpD7UCke7H9DHbtC0V7hpejmBJw14j+dRHtqTc69tOAd
0hoxaRN2sLMr5YUhVGBGbKNvZFRhUlsiO/2jhdPvMK6HcaZG8hhjnCC+HXfHhc2l
WmieJeCqflhrU1xVI/mwoP+hZEtvxv+8+3xd3znnoUDxeX4LteJ8SwKOaiYrxd7k
MdMJTjZWBjQ+54HZAEZ4vK+8NyXyEceTEAKZm2kT1etk6H0hH+eyeuNo8TVZ2SvM
OLcWxaOgpNrKdWuFRB+Gkgo/Evngi04idZ6wZdur0fDBnYqRmkA0KotwyHcH+O7a
sGWVwGanypH1yDLV61bCuQG/r82RiRwmZv+tzUdv99ED361N/iJ6ln6P/uuwEBt+
Tuq4ttCvcGUaVkEfHn/uanXrqbmYxY161Vt9teQc167WUPx9lKXbWE3cVZyeBmHH
dSXwWbEQciDoJrSSrwreZQ==
`protect END_PROTECTED
