`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+T3yh1Tg2s+PsKSp/bZ5t6J+FR1th40GkWGyxh2vMsSv9ASVCr0Uz6mcta3aPgH
Gm+FlcraHHj7/e3VfM3Q86Hyu/CxlYmGNxlzEHDUplBTS3Kgnh2RGFnyOxF+V+YG
TvR2EaEAyX4zgy+jzLJwzkXRGJI9Br3cEb4Nqoxk+YpIrIoRUREKRvW81LI3bDiQ
vutB58YSaPCBSifJ4sf1PtnU+GjDARIwAAiNokootCOaF89C98H1d4wwHyNAlzCj
n3benon2YBTZcj8Q0O6Xavm3Uns4LmgwhfIl2Cej3Np4tnvvGnNnN/Wz+IOMmPsm
nFNm9Cf8TYabCaTx/nr1zg==
`protect END_PROTECTED
