`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Th9TAUku31f6wIxvYQ+wkrlm0vgk2sHrIRd4DLYYnO2X8iVHGp32946vYDa1pLH+
0B/n45eNSs6HKqwhbS7cZuX4TvGpkiF6BKVAKXZoim+aGBXUgviEMQ90PHjUCoE5
Mx3nFMxXRxTQOvyXCloo72wFy2SdkgemMv8mizb63r2G8JRicgY28Cm4X2usB2br
AQoSzduoAb7h9KiF7QC94/WhkORCluaKN1SKi2OhLouA6xRiiIheyj5/69KEdki1
3sgJ7zARy8nQrrEzVxmZDm9KoNeQCO2M8gw7/8Se23Xq9QJuTt6MyTWOB2NQwR5Y
iJd4ePNl7ZbS+XyS1mJPHJbF+uxOfrqrRkea9jgUFqcfTYhFRIaE4RjZt98eylDq
SuaumSXP23wyl4fB/Or+skanASv9NZEllVmPZglTtu0yvgxOlUhkYm1hhx6kOfsx
EPx3MggfXQjzSltgoLgdF0imq0fcyeQHjwDyEExb1Hce1a4siV3ifHhBZwOQ93sP
0IDvAuVZGZVXwLFh2gDqJL7kfL4Siso6loZZF7TnqeE=
`protect END_PROTECTED
