`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZwOmmik/l7Cew8XU46gKuJ0j0uh0RT227InKfTUjwZM3e1kiMc8+1MkUKJxZH9/m
QRXWCuw/EVyU//BveHkqinfTdjptKZMeC0AhGWIoFIMXochNcTRFSgfM68XAKi4r
iJNSJQKtUNQwEBbKSeRQvOBF1IopsRgKRK8d3lmO/NbmcIhtHHVgTEncKjbo6OWF
9t5ysZcF+BEhS9Fanh5GzaZWaM71TuKTkzSahXEn38Qbo7af+1PLvtVajk0OYJCK
K/2daMysiNG56UjP5rTuWNRC1CT9L8d9eefyww/mNS87Do+HcZy9wY8ClbVwgw11
w43uv5V8E8CdXgntOgxJT8xT6gnuyRPA4MQ+P0AlMZoCQIZl/MV4NEbGAsdOpkJ9
B0ak3zGPbDfJbZW/EEQAhw==
`protect END_PROTECTED
