`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zhsPaCgFi7ZNIlPr+HoKPFe42UBOzTAgeHcM6qROtjF/Tu7Ovsx4H+1Z9m/NnjG6
k0FMxGeiS+UgSDc4CKAyf7HeA+BM+wHJtaH+dxDwtuZO9XsDbtXXB48ODEFiEpFr
/Z4bHoAHY0IL0p+TKPaD5Bt/fNxO3uaguvE8lG7WZ29Gj276Flw92Y2PYMbMkxQ/
650/VE1+YsDwMKV3wxQcjMbkoDpEvFfOgGwSGUZ/rUptfjLYeYXZXKoWSC5EIgRZ
YbUe6VcS5u5gwSMRb0tv/MIUEBP32QI3dtP+EI/Kn5F/WrJnuNWhMdDIAZmu1G6u
GNa74x/Vz4Tm8bSXrVofN6OY195+7sf76NwjZwJlri+sTJxazlY9Q8X5lG4Wdifq
sBVlFi6ftvMeudk9xluGpMzCwcp5FrdWbORlWlWGYbyMthE7lj5+6gmSfTBdCN7Q
O1WDn6GLy/YP5pC1jwO1dGJ/9m5Bex/CQBtm1ISeTHi3UC6MvbZsjlWXme+JtnFe
fXB0htW8VWC8ow0shDUkOYsRa9oaU40r6d8GAEQsI3CV8FMNcPwaZR9ZnnBWq6lU
LvVSogb5M6tBd+bqK/1Iw0FePOPoTEjuVjpbRms+2E2XvlMM+My9EFLrblCL8PLR
oc98nfLeablHOrf3iUF1hDKkYu6t4Hs9GZMhLmVeSSNIlbNwoShgJmglLkK2tmME
07FiFl6WoSIkSHjTWYBvuhY+h0AXjEgtF0nAfMz1sYOv1SEXJTuO5EpBKzquscII
E4V12K3By0TyBw6AzbIyCTiqJafqdPhhQik3Mr1vvufa35wMFXRPK3WKXLFz6dLU
Wyhe+ZEMfTDs7KmCOwVjB1MzR7j8mHhJSiBREPn68Yw=
`protect END_PROTECTED
