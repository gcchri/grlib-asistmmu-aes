`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFeEsAC5FQZuqXPa/W1CI9GIX3M4yaODTVKp1j7IAC50hgWYBbWIwTCt9Mo2Oo9b
J3CYjfYtE3PTlMqaJED61YH7ki6ylPKaTLjsmWE5UwlUasdUcujagTsAGb3mEHSk
w3yVagawZ61VaUuK5UFSCFqIih2OLz1m8aqt/lCZMIlnnjpkYSFUAyX0Q4J1dJTX
d6Iw2ViBeLCn7vcf9MXgV2Wo51/4C96q87MkZtCFaqYqLDQkMgU/YmIqqzwqgM+h
67JDwy01yo0eKSOFucB04oSdQscztr8rU0hgQd/AsgGX3fiqNheA9ttY9q4XyEKJ
0ec7g1DiIyD7JoHQDdwAWwLSPbqNw+JVVNldzstYAiWS3fbe/5W0CTpzRHWxVQq1
VYAgrBn5/ACuDnS/XW0epzdcTnjowWjIwz9TDGV3/K8ihdI+jBLlRQP0TKDfZfIE
YCvBxD7ZJWtS3MW+Lbj8tjDNwRxcQ7AsELO1dDMbu054AD3mzLKfR4Fw3mYMfFxv
`protect END_PROTECTED
