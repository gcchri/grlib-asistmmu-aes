`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npJj+KsEtfxx0yzfnvJqT99/CfiB4CC1PZ9ua89a4uYg8I7ZueUz7RhgkhGWHPde
+PzAM2cdiQwZN2pC+cYz3sRsZf46pzsu4BT2pV8cHDerMZwJpiJz1bQXO6p6Yicl
VMO+zG8EXcopT6bkeu0mdJ6NzVYtiVh06j71OsL3+NLbvam8Xyud+YsGUJpcoY8n
lbLh5kWmuOHWbcgVzzALESE139dEOKEJyfnMm73va9pyPcL8ln23aDXGm2+X76IK
2yxLJRnhCqQ4CrWtCqxosFyrmxi02rKv9SYiMjnxNkDr/6mnDSpLxnTayy3wUrnq
pgeZ4COWq4dB7lYquBhtytPtREeOafSe2y+ir8SrGRhcuSGnjpOuTlqLig+eIZvR
+0YE8DhsnBWL/SCNgploJVwpBfc6WezFAx7kg5PCdCkZLU9Of1wp1y5iTrUOZLZR
`protect END_PROTECTED
