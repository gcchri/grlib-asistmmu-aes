`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bvt8TIXWfc7D+N+JJv9b2kSp5Tp6PjIsaf1JQNV9+Cq/AFjZkWi1wQYtBHB/igiZ
XPcGQoxFtywagzbId1PRFHxlawohHhesq1fLQo4LMEP2XZ0aXzy/Qg5NFuZ0YXWt
cKIYPwEw2frJvS85LWSEHXrE0vWAoConjXyIfU07BoArhHICMIIlwcTdS0IZQDXk
+HpvuB0InGLcQQ76kMtewjwzKQKipjZUpYjyHrBJkyQ1HWzsntCLDxAlsDVQe3gY
Oyg4c6cxFrmGYu2HczmdT+c39fY9p+NubTsTIUqs5uTf3cvaz3IpenO76GChcRvi
Gikih6pg0UaPWecuIMdNwnbhp/WJG9cAekTlxXWq0Rr7cSA9lFz3DTja2gNyFo59
EsWLB7fkiO0H749j+h9EIbneTwzoF+E2HSFbmrKR1WwcaQ/3SF0o0yhMWvRDoiCY
VoLHhrmBNVKSViRROJ37erb5WNNCAeKQ3Fmn1XvvjGhpbZ8JNpsmbVCdinFjrvtm
`protect END_PROTECTED
