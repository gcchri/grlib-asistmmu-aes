`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mE8q+09OfkrLJXWsuEyC5MoBtuQ5k0s8HI7Cqj556pFBwoPaKyZEnaBwwxx6CmTI
n1ifQ6hYkpGePG4hZsAr75iiWCUfd42HppOW4x4NSd+ZQlJdWzQ9kSIOLT5FTuqt
ZTcN7ls9ZxJZiEAFtgWxUCmDbt6DlySGE43pqLAnPfYxxRFGYGux9q91Uz+6PLUS
q2R6+ZVpyDd5QN0gRv18ByYtZGu0dbh+PRijd5VQ9+V2I6q25sAmQWVHls0IXwu/
VfHzLGamQmWvDZxtiSTpLdpCZGumvVkliejqy5/Cp10wFYWxq8RENyBS9hZ+5y97
9CfoCNaqImnlKWCB8EnQh0DOhyuHjYQl/1X9hpcR4CvQqiS6AdJopkDUDasjcjvv
6fkNfJFauH3NAxt3YOK5+tBURN5pWcz2rXkvrasDyUpt20NaO1ejFKYtOALeWOwj
dQ/S1vRiSkqvsTpxMOUoBxRGKoJJ/xvYVNvl5O/W05tJ/pyL815AwA2pHspbpIVy
0LQRAiSr3QJLQSJLkjqrASBcRHMdU6utKn/Aev5wAbVWEClhOHL7KCvu6CCVFKz0
kHDmAoAzpTeDqzAUl4hnsTnlH1T/hKsIXiBGanwXOqhoFI4c+kMyrFfnr4/B280n
bT967bULsB9wtUNKeifCRi0kIycajnF20rHmoEQka20oecJtnHDqK0ipbahvziBl
SbkvubN1zS+a29TSSrWsxSnoE+8bOrD9kfDdkbDiWTtlh7YowWQJj+hJHv8DUAUv
uUmqIU2AzvY2U7DZP6/Pqu9btUHLQcaq/WQq+tMKkMG8hINcnt+pOS0XTSZR7RU4
Zv3Iocf1+Ir1dalQSqCIwTHzUeRTt/E7MADjm7SVWjKnLD/+InZQyFXUiTSWS80D
prlb4t06GhAFyd5KNi4bhZ3TfYcaNElSmGcgY1pHcauChNQE2SbvAojlTurHM20p
Maav+TtppfuO3GEtPAvudCvHUKyLHvpinJDuMnm+cM3a61PyShHbQ5vKWE7OhUPO
ctUi+T1hAX+uVbIEpNV7VFjUB9F6qbeaugxsSbezd9C5rUSjuGtewQKgxHENMRyZ
gyDso1d51yLPXq9WTHGq/Dgnm34p08fzmatnT16lYykDBkyYzzNHcdNz3HDDISO8
ehQin7FE4gGeErxvSzjuIMHokTVkCdoFvA2CR9JWNNFPhwqThiUhz8t9hyeOXKRK
ao+fdjFSz06toq1duutImywmvZu2ZkScGYJg7vVO+fN0+vgBKetMI0XyxPFRRGq4
ZkjMHLiUfvkeWdk6mdfDRZLvbz/IQDqqf5F41QQrm2VOwxQNMjxZ8fVOOBvaktSc
xlr2BuECijllrdFrInwh8tbPIf6Bhvap9r77H6/aiEsc6BsqGemWss85bpzmN0UT
xodwrmOSXsF91udWoh567ssoJh8E+TvSXPyAd1vJOu6CvkNwN9dgoKmp9BxCslhV
kh6PtaHCY+g9sFgEnUVAWXpcPzxCNJ73vpD3OJ48pCZIJwapq2ah+eysCR6lU761
DueyD4VjhVg45zr0wgItMgWjlYz+E3rhDRCpLycJW7/bgZoGbH1MOFtlTnpU34Oj
J2pU/4Bw0PT9+3uAnoPj8IfnHdqjgn4uByQqhtONRMWCzcLNwEmGA/rkwGofY5EX
5Bt9Y7PjyTpUI2x47wzcoTu3FtrINBoBEq+JIc6mFRQ+8NAJRaqczBpFZ6Bx5Bp0
qqV31u1HIxHyrlex2Vb7RPDLu9SK2WZDl+bmMyrcNBVKIV+3GJspPhp4zD2ijb1w
O7GyC5SmX6GpXtLEN2965JsTRjXymvAAtgHlGaf+SeAov0oJs/uhsItQt7Uk/JAc
r7Bvx32sUlGjo0+BfOUywGOBSv/Mrp/FVt6ry4jgn5xmqlkvDLaQ1+2oxlEx9ZXj
zjd/cFd0uZMMNfE5Sz1L5h/1KdbjKl221vdN9bCVBUl6u/Id1ZH+OOZhXxSrQBh9
7c4FoAKWSORyAN5St1Af8XMocH/Bi8ZIAPt47RiDRGpWkQXnrGVQmJlxpdjoNjZM
u14Nv8csSXHvradOZP4/as7ua7aFvhbebJEWrZQl7d4U/Scg+MZ31HrupHAQniza
KSIWZrP2L9z7J3KzUmfJXWDMCrncdQ5gTta86SB8diJR14geTMrPt0wMlFNy3gZK
A9O514LW5/YPR358SPVPOnBN94KWGNeY24nU0jzne0tgEInTCOODF3FAKERc9cSq
m4ZFkVVJQBTjxA+lHpNXtELnAICGIMk/nD5LoV8cW3b42/309MfZtH8v6adm6/w2
ClmZtUDSkRhsHvsAKtBkHvGJeb3XV+yVZJaDHlVyud59sUiCTltRMUeVKuVpP9J3
0NM3Nh7o56NtJNIPhS8zx2ym8CEPIEyMGqIHpZ4xjyTOMNPjerc4FYgRRCh6a1U/
Aacwxeh65vv2wPvCISZcvKCOWX90aSOPQywbT2yS5Af/eOyHvyVR1+Zi6X3dviw6
VAhwmcd0dV0lLqR5ANfGZc41bsfJcguCH/7zwdjdKs23ORznoHskvBoRbZIT0MgZ
c8iioFGMDW3OAgt/DZNkC48g1TEYohalVy4fLGtLHF6p2qPfQEl/powwDqfOTPAC
+VS70ISdjXTpJai4psuc6I9v6pbMgkdI+jfUiPcWObqmpGaZZLPMvMhvk0FQDO1Q
ypEiKTiiQDFDDSP6Vm88q/jFkdcn2WNxdTGsAePM0cQAEkL/sAvGJR5ZDxjpZJd0
2p0rsFx017sDqZc1Wn9bxOrLXAs3sFFzpZg9IY593EtWSP19yP4RbiR8xjROt2UM
vdBuhs47hhp9MM/eeYKdD9FJbfNwVn6UDMAXRx6MwN+CRJywWMUylK4GMreHzyzU
j5f7w5bKkI3roq4hShDhBqs9ZtzPkXHPB1Aaj7zIL4mWw8WiyQd7yOiMw/Gk8yoE
pWmmXS0hKpoRRYEUb4DHY5E3hDygvenCPIyyv6q1WakbNOW3a8P7gGmTjBWY9+r7
8NmFsQOLRkg3vgisP9/JmSIF2TvLHf4N6uOxP/UP+ZSJShWp1wy/CP9UyW4MJlXI
cl99Z7TkHC1j2kf+QMrj6rCJUdZi3rXECc3meNisQtAt9+/qhlqCUTFxt3ZSR3iM
1hlyw5r7c+wleK3K+xgVDt9p6pMOs4EjEaRiidLKg5SHahPjZyXFs3gWSMPqjDuW
GWnXXLntEvQrW7GLF9oxr+8lt150y8gAF1iM1B0tXgVRQ9iEZ3C47pQCBMDEWXhp
ocIxdStqZaTnXrSo5yMGe4eDp7PkfMuILdssa8C2v+4XpPQ/d6JAImgxeS5m+Xr6
i29FcRYaT73UtBGQDHUcwaR6nNI/h6rFLnggXOQ8z/CkL2xXKeW76CQo0pHya6Zc
FRs4lsWlFPGMy74dMba7VqkRAwEdXhJLHnqTAVjGQSEMtg0asDC1uw3Sqrzhptea
j8tLuMfl7JGhrjbp/b/IrrrZLSi4mgrCzsqePh2obtkQjyNmqLF+Y0gtRheogbJj
VZNY51Bkx3Gci5psO5lQTtvkJLdKeRtOL2AyBZK5G4uWQqRRWhUWxcLAUIegDrD2
Syd2V4+pEW92SF/HEKOSMOHJOJPYv0XBjWGCVwLk+dKmrAhwBkzjBYnuuYCD6CUk
X1kffSHof+10qxQdSBPwYZseajQ22hNh9gZsz41njiDHn+uymJXPpl7pQJ64VZO5
G+7LKAjBQkTObwHcSZUfyFQ+kbzJbW62RD6m4k4fvB33nq2vgPf0M0Ewe9/IQ+Kk
Gkiw2ZYyTYPrQBAhk02FX+9yfAfwa80EylO/YFI+THTX+Jjr2OBIOXkYgdalfSAO
hO3YoIchuwaCsiwo9BpqJAJUnoUQLQXTkpG9y28Mr0iWYpXCffDs1fcVPWTDl9uH
etL1DesPzozrfh7z2gUBq4NDuCONAdTMUqmWq877yC/8AQEO450XgOdiAlQ+XCHK
7OOSWZDsRIrsxJ2rFf1c/U28wbG6DvLo2tGZyZNlSyGttqBQGqbTJeI0KKD2vUc5
F7PFZbZdyLna0R/PBf3HLIwi1mQ2a9atk4DsPbety96HI2fAJ7E7HnIm4ZeX6xly
V1+kDFkdSiEbPGUnOvmiO0VdvmszX4B/68wrZ5QMxxmmE+DuB5fSxoRLqMfrFYjt
QemZrI4QxY6qxBWm1uU9NKMp61xwZJDs3UMIeJ2UH2wJzA2uSfBl9eQkEoKa0QUE
3R9F6FuW0pl+e4oQZYW0gwWO+dfAu6TqITaKtqzmsBQ7NvyPCclYV591rylyiCYg
jwoqC+z1Hmm3+KZ6ErHPBLbzZINppYY7hsRrY8hpUIfzTHDiX6hJjMaLbtoy2t7f
zsirZomjhPULJVkpMYdW36m6wSmaYoLJqgp46fM2X5c3UKqs0GWDERvWTbIV4ews
iCku5wweUOez7GNoHG+qtHy7zMTgjJWc/nczAPPgj2VBUf97hzLGAQtExn16KzWU
OzelvVsHNJbSfc7uFhr+e7Z+ntckvHLDcNygkaS7hxqY+2uXSnJeAc/rcmNXyxof
+t5tc2EqBvhs2PO60+dUj5zIYOUKkbk/VmmnCUHNUVlwKMA1QK6XSeBm6Q+ACLg9
oBh20OZYDyDC1zX+y8U1x2ua8g7uPNoMglgmrgxbbBRe5t4qIHI+oWlKTeJ8Ki8V
jZ/QuepfJVgkvTHPoOBr7D+/tr+YDsAzNfeiAZoJBO2ApxMp74q3SpFY69akLj0M
15LOk17htTL21XgeU+BZEeU7s9Gq8OqsWWS7+UPnFPu67kSo3/5HYPb46rsgKArV
KIxG8+FZeGxFjWKvm8X8zyR90gD3MxvFkYqQnzDAGy6o3hAdH1TKRb9mhjjIqhS6
JsRJ8H+vzlJ0UeiysFIO9iR92J4M1C1o5u7ndyZNr0jikroRqx8aQKxCj8FMsfm4
ah2/2AV5BXdf++FRLNJ7Cyw9hLUTNWIjupupNQWchMYUI03On+SwDTr1MIeFrX9H
/vGnnvITpPo/qkgaSO8NpzLULOx8a6GUN7QhwqCb7ERy7vMhjhF0NegkOSQBwph9
11lVho1h2dmpAixbXoWalXRYOt3ymtu+rsLDqp+sZcFUy5hVkVXYb3ea9Iv7leoW
bR57s7/OsovE/4ApvdkRo3+4qcZygRnIUjezVAA4uuhF7sIR6HmAVPj9d0B1lDzO
15i8bMZs3HSQEegx8O0DpbvjiLJzDW54cYqrMsQefKrbcutvN8BwijY3RWmQjLN2
jBscuO8bacn3xv9hdI/O/T1XV6Q7W2XSKeAHbOHYzABPHoSge7mJ0gIsT5b8nI1K
5fKuHO5t3GxnPHrQL8M5vlOPaBDIHDZXibaj/eWZ/7xKZK15j0Ni2cGh2tjnd+AD
doSs7Qjjcc0PQP3oIVIa0LKR6TysgeAaGeflUIRaMydYjipPUjDub/YTMrYCw6tC
x1tjoRB/VRdWyRFPcm8vRq0Bq4VHGLuGzG0ZZp2G5RJYZM3fTfSRn5u6A1t2AexI
8c5ZGwkWhIGfGoYou0e9xvQo1C0JHDddMlaYiB5XmTcqZyT9A14QHzg//0ZLEGVx
z/WvlO5ViIbQnwAC40bxdP/bnb2QlxkQ3xMZm4R2Jcr3jxEq+cuMlEKWLcyDLJVv
TndtX9nJoojqL8iqUy7djcHXzYLN7xPJnriyYWAO63njz+V4Bor1ftJTaQCLJ5QE
xmiEGTiMnSKI6aaRokbw/2DAvrIpe4zE4CiErZ+T4jXpvnjDjARFr5gOMDem7w7Q
A4R+deEusavit3LrCfwbMT8o5CLqQROx7gEGc/II9KG5H4k/sYFzvnvy+ur/zVJK
KDWII0nlT+baQl4i8lKkt5asjF5zhigotF2IAlhc3jg8FFY2TT9MYEHOwzBzHAvc
6QLa3TRlJ6yORfEvefOCR9e1viftDuADPpbnjVA/zC3GahxZ3PTUojaUK3ZhShcB
YK85L0k5Us9w6VBjulAflMX1SpXRBu6JZj0BW5OH3s6UG/Yb9ohQUUQc5GjyJBM0
tCTCD2NpGeUb1Xd7nFximWv0WdqBS722Iqa+Mgu7Rh0RHZIT+vNSEf2D9QOQyI6e
VLMIYFToM0anArWzvj3S2Hdou0mJAVv+6ZfmRQuIyoYGnuFHdu7F0uRBqhuZEfu1
ERgdMcZL48efeJHXz2S6h1Uo/7rKo65tjhUcCJw4TnRjQqMfish7+CLfjnexTnRr
MWV6fxtaO1av5dadk5Q/uz4jX2CVJEZDvJjW/T55nn7dQCbC7eWTMzx7r0jHj9eW
YaXwWlBLmlnssweFi0muFrQQBbfZABHFsxwWlc9efZw/y52OgABenmkfRu4TlKK5
OrD92pOSlLDOdNgrNbvil9u/56kpElPlT4OC/BuhXLGSjkDNR1zXCWPEhYXKu8To
tQg2vYZoXqQ+pJv0u1E+HfgivfZfdw+H6b95zuf3xA3rNoN2cBnZ/ArNXJWFQ93T
evHBui0AR2bs0sBoLV7oP+z/OEsXjg2xwqhWpXKJyY+KkIoelcJcPCdTsplReCIP
uUrFwYhUfq3wpDq/Gm0VntqHgF4m1lhSsV3xfi4OAm16dHqVyDdsWsuLYWbIYqDi
SRjSAh8uDYVK7ZOK6H1sU/lFXcI+dI83gfrzG9+SQtFlaaH1StSkT+JDV4CL9QHb
d1+CRi2CacnBWM+bGtPUttHTaJhWuAo1lKIZ2gNOvd7IfXLDEHe4XxeB6nPSR2Bg
ezhBHg7maYllq1aDNdU+cfvNnc4eg5kSJ6g1y3zlEYNHtyAR0wM5Fg7G/PQo7xHa
pHmhEWAM8GyoeO3aqcVdWCAfhYbNl/ztA84DgyND8wDwFxFl1sK65fLcuumDRdlm
5hxhmOnzxehqGDvGw+B+duidAGGKUnFXF9KicqleGNNpb7k3YFpBjKX5dN8bn6ov
L1nvNdg0eddeK7AzEbkcYjFd4LMA92EJsvhWsbuo0/1Z4ZlDg1nAT2wCFJgv7p1r
Ez5pGolSxL6f8Rzy7wA5ftzi8JHgNlBFmhAjvczfnDlgYeyCK6R10GA/g510o9Mo
WfKbYGJJn/sKvQbfcV9mpn1afYGCImaD4o5uiQwaX4b9rmSiiuVwjHH/6a+oX/Gp
JbOp2rp16/frqW0dLZ++4+J3gDvOg+qGs8VSV1RrjzBtZQV0VZVYEIMYiKGyDRrS
xzitWCveX1x87rTHUNnrKpbLp77au6JoDrlspAG+Jq+EsjEyngHLRkpOlcJfF3h/
QXqa5+g4irMZlOUIYKP0qaATMC2mpmbb0XBEj6UAHc3dUMDpyZBcHdkiNxm4Mlgu
sPEbHEPC/CbBdLRUcoHnd4laXHJGEbEy/fRj+rd1vxTwBBvnjItKqPZ6WCkf8V0x
CxoSy7yjteyISfCLz1etEnQ2lpF9XTWev6KDwV3YDf27FOW2gOOkMAKtmVeudx1y
P4tGo0hCzKNTEsg6qgFF2zy76qkamThZFEi7mCUZPOP3v4t/2AX5hVsLNbrq9Pcr
sogfLi+hWI329yG9Zd7fdstqu6x8sm6xxv7s0YdyBtFXqIiY6h3Qv6aTIqgjKy1u
/A7zLwf+099gMHrJrO3Ly83UUTT5wsvuFLIOPyI9GMXcT913LjO/cURFzR8xQMHj
w1XBfzAfzevqEjMM8v0m64GYn9h52DOHEJgAx3pFseug89wNnEs5b71CDZEX11Eb
zqpIRp2jnuZRTUupKmyPtc4u1xYS00MO4dpLs8aNpviN2dccQpHI1FKMm9UjFte/
Dq2ihJgZw07A12tS2gEUUtJiTOFsXDBWCP5fUUa0ZxcnhCPYg8baZERlBr+apWZ4
9F+CPupBMeh/frbfEdagRgq+zHsi6/olchA1ZI5PpQH7iF2Lg/GPESoDTDN6jchL
r3T6g9QbrohqBJrwNOy6pnj5zEVj8/Ju9umVyj6o7rqjeh3IOiVSC9L7BJMEYuFT
1+Kop0Mj2Bdzx1AiQw6sh+EfJbp9ERXteEVTO/460I8rMVSeqxhIfsRitmVB4MPV
QL91naBdc4r+G/9MIdr6EvKo5YXwMTPa45UxqNNr9UtVFgX9hN9jHr54kAoq5f+H
z3Ewza+Qsgv3ZIWHHtHmpBrz0Lke4SOr/585CrlyNv37oAjq6FkxKMeJlF8D6O7C
bi7NsFcImKv0Lg0C2naHV+STVNPsVmdGhij1jUDRAV5x1E2n3I5UFcsh/fLeRwV5
b/8Zz6GU4Hc/T7DNSu2omXOPNQhaZWvJRZLDcimMwmDrh24+2gYcTP4Pab39HHlK
jbne+YJgjrnnc0B6W0D4l+647iDkuuxWhXTpIjyGHQJ5A/6bibRbVnOb6W1iuNi7
AjeGpJvIxCHpm0rZwobcn0STgfMM+wwhIE788bkoon4F37L6Dwx8pfFbY8nnLaZ0
s5LaWY/YQ3a+2lzxZHJNUgT/k5zpEVdPJmizrjtt1aHAnj+aULauNnUaCB39wy7v
weVfgNS6dC5rKKZsdS1nQvTHez9VXfZ3HmCTRomciCEYZerBode+4i4aTx2klzXz
INvZyPgYdXfka6EZUmTnOfwK8Y6pebnAvfCneVclojq7rhq/zXiV6Rx8bfg9dZcc
4dyPHgbnLjxqfdEPTLdoUB76tONiZ9sxJIFYqAp1enTnRZ3Y2tDynEMQZ2IMegSY
lSexDGyYNMSIxrIQk8ydMnkkouSxupYjXkujipzhyERt7MtkM+j2ktsxQyp0dWnd
Ahq5QLQKGTmTmeaaqy2IcPwkYWfnulULfA50UyCJIGb0YbshCQBFL8xQlOhMIAzu
zgMm3G6Sdy7OlGX+RSLgFSjpqSaGjBvwqIY7Wg/pPgFwPt+IROLQO7QvUa76rO9G
CN7qkArCAypaENXw9/1qQkH9oDCdSitrVqQQ4bBImUM82Xp8eA+rb49kzFMQS1Eh
oDAa6bWUq23tqY0O+qPGE5bz1YK2i/Utev5AFpiHAEnbCF0uR/qo1yZXlNiOpUV+
zs9+Bpb8muaSlRZpAsv17dCYK7BXWAg7eiuB9v8kXo91Yy3W3L/b50Ir+AaCEHuO
gWhYm5jmzo27S0XroUeJQ1YNFtj+Q4j8j61Q1Zy9G8250P9wC2Ph0orUObZAu2MZ
Uak2zRPbq+0C5kMZS+TqGxDqJPCsMX2JLpna7e/1gtI8e26eF0bUz/4FLVvzTfCc
GVaeyDtvgTzVnT9EckmHK3mdieIrIGPSa/gwZCTY8sCyKf2XyvlfjrALYxov7lry
GC6BIj0IjY10D61eVEZSeoa0KXCHdAJjYKkmSQ8zRQ/Mbse8RHToK70lde3CdI4u
D2I/dhotHXChJzBIOldyymE8qqOvjakm1UKhelk3nU/SAwmk7sPnCXfsonoY1LJx
8twZ1McUJtYuPghEAc0FEFIFvU4g8fdkOaR1PR3IVv1Dc5adpH1AsytHA7PkinZt
s50suzdhc8ajVHZTUTkpJEeCh/qUn5dkYBhRXeXXoMgeU085z9LAiCX1bprodSdZ
j2s8OYhZHOUsj+kZanyBZD+FwBM+xIwoWBrtaWddIDkVxwf1UF8XjvMeFrdKeye/
+o9HgLdkNQEx9Ou0jZzSLKTRwN/pZu4fd2yg4k22EoEJ38a/nv3ngqqmdUPVQtwU
ybiIHye2soUrAJ7DeDibt/rFJfe4DrnDTuWpe/2x6bbF1Jgm88iASO0xoazSO49A
AxiwutX0A8rhOZpPfnLRqQ74ONILwGhmWG+jKvO5GMzJGlr9cqYEPTzixUfq4E7d
qoY3YWmES9wb71m913l77d+wICiFP/esojSSyREawi+ZuTkYClNeQNu/+uy2rKSb
iIMAqTMNSMfcZ5mO+iG4IUfDORpxUyFKCQ6Ye9ZQrM8RcfpYtnoYBe7RzXNfNSPx
YxwGjsiw8DWFfgMeoGON96mYqWp+vv5FByVpM5MCTAE7HH5iYp/EvXICIf2/5Tf1
7JST3WJDyVKR5XoXCTwXG9rOZYFEYG1OuObdS7FdEaJGGSWfckW4A1KK9B7AGSnq
kdce0D/D5fk//KahqczIQaNTCpIREWC+yy42Kq9PqjhBfQLjYXCGej7AHG555uEC
HqHCpQMFTwXQHLG1vgi/GyZccnbN0Vbi0B/00fTuPONlu+pz9vw1UgRANZxvW7OU
nmk7ZiyCojkIj5Gst8MjIX+1QNSSsmntLML6zrCQ/kRPXOiGQDtFC9L3DxknotSU
QtFyaKM5vHz/rjo9GinrSUjpj1cqQcAda6RcbNuWu4oWxxcqGq9dJdytm/1N1dTU
VqHOSt4+sOja2XCt/5CuVejtHA+WCk8NnzrRBgY+5/42VOc55SUIyrdzRF8hcQuE
QoV654XwA7Kof8w+stT5WErcbVDsj2j2yqvN5J4ckli10NrO3yL4PMFNuDc8WBX1
sXFDWyjACFlJXCyI2e+XhiECtcinRxr0z9xLO5Z/MLmwWNsIPvvw6q+xHk7oGHwY
xbMvqmb6jmPN7M6XV9ZxpRA+tSB2Fc/zUsuyWSUJ8o4AuXPXwnqpj2PI2ldQ9zw4
x+G+JRX1+4ZHHz/Hi1/i5Wq0PvVi3ucMvhPqWHelemcIuUqtE/pxRHb0Ml3tnphI
K+dR5mFtgTkqCZifz8fjUI34B+BrQV3KbqatZV3hLoy6cEt8PJZZDgbEUPo1wsrY
b47RANePbmNQ4OamAa4oLfhIuHrcZxB6ZEDQiNVuxybwAtvQkvn9dL1WoeQBDAW0
pJFxE1Nml3EbdpvVIkTwcjgv2Z+XyVJE7etZE9XVOmCL8Nh+rmIKbJcKeschaUrG
eLs1gt77mHR+of6iNrXxpsFJye8uSFSylam+AyOSPrQckx5FWhrsHOrOnYjXv0tj
7kQPmLz22sY8VkemA2FaE0CicJjwdzYnK+f0/MsqAKuxfGNKVB7c3JANjh3gQTR1
TwlMhHP4ucOV8wtnUFEcv2lQUUEyz3GXSgKsCTb2tERFKNq++bHFXfSRbsXUSDMX
/a1rX+YqHSZ796ioNhrzbgw8DCUs0E/ukv51XjQgsRZCV8zndIg7dJA/W5Vye0jO
uTQkaRxB/veT/y3PwG6bV7v/2i61NUPGELjbILrVevb5OO/PjPb3Y2auxLRha4dg
ji2g/Ay+/TOx4mkrVTA6Wwq1f+B37XAv+UdgX1rW5t8Y8mf6Y8DAW/zwfA1Nkl3y
YiF/BA0REB62UEJgyNVHM9bUE6o986aPpXQNxr97chBUoX1pKXwkn5CCz3EE4kqx
/fFYVxg8DaZZJHdWhUTkVHfcozkg2MCu8v0T5EbfzRw3QdrWOpGVgi6Icn7OvIL7
I4u5B0h7jWR3hohb82YxiNeIskkOIQPtvrJIRuLZKeaToH61l9dRoEzCAUCEokzZ
9q0CVQNAAw2CDVS7k1aWMaThSE9p3tx7XfRD4ZLnbfj5DmswcCkTTZvYnD0YsJrI
CLB6MuwdaUehkYmgSciBZAyew5sJKelAf+aoeW3LW+DU/Sd4mD6qT36p84AqaxVW
EPO+hK/bvn9+4/pe6lwj7FYy69hgVSjjQjM/p9jI9IRGW0DvoZyspu/gyT6xnknp
vtHlTwYS9gpVOfnwj/7bKDhpJS3YJkmabxHTU/usFC+RYyFPn9o1qx1IZhpV/Jx8
KSk48Yve3DqgXEBc5G+s6g2a1gfh1Exm275EcIhUCFKKVSb3NCnowcC8id34WYJ9
QTyonlEyNKKoVQDtOH7tswOuRsNyrp4Bhwr1MzBO4a7iq/kxhna1BW1MUklySfF4
dxhGV0KPiao81Tb+FhPx9G0KMscfdoSKLTqVfDL/rJePpP/S9UDQoAY5d1JBDn2J
0SKJl4xh89O6yQwQf9V605eWbTPtgacU6AqlZL4Srm/JeILmcMk5hlkx9HLzjTki
2R6dEdisfyzYVyNPgolh0gleSN8As9IPT0Hn5tgE1OyaLD6YQRs9fcW9OoCUaO4D
TMe68Hd4XeOMlWwisefilbFOt6RjlofCxPivn1J0rMmoLMNF5XJ0kNGyRggbykoV
3SJeZ4K8TIXLr0j0/g/nhFslLUHPNTExQKeP9E/ZFVxYN6S8R/0ZPdVwgC29ZLSv
nTOKaXlbGreK/5f4jJBl19RjL6FNRj8ar/KUryHhOntm21pKusSc4nBU3Imal4eo
1KhH4+I+i2Mb/dUH6Q57ie8IonykO2+mRUfAU7KBVF6ztd9mSxwfvMYfVWWTsG+S
`protect END_PROTECTED
