`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ncXOUUlpZorpTjFcSqA8ldPmT6qtCS6kkb4q/PPhH+5lZM53HajsuYg2Nti38tJ9
ErDgswJM/uRCSIqth8sacR+W2X0wNCaQ0J8SaDu5ZZMfRmPcEOT1AP+QggwIMabA
7u/Faac+Oo66V1tWAbdA06se2SxKZGtTLNJOFiGM1CwdtLY8MJSUAll/kvEHURcy
ldqHWElMuGU94whLnCx9/DbWf0UDUMcTGE24xbIJ2WPbKst98ObPjmylWfVCAz2f
UqLtjc05KZPvr+IIu+UQLMN/lscQG7oVIzjACYs+9JjBgG/ZCMPxLtHY0qpnzneE
jQnjYh5Zf0UfRbOsHN/feeg8reurzt/OZknn5I/pW0k+pfHKvu81IXr9Qwj7UMJs
5E87ND7TOL2zF2v6+///sfVzxq4tNxrMf6fN/xSKOguuMVgzvL0v1wWs9MUCkbaA
wHWxei6z7tpJGjvOSkhJaMoud+EVF4O9UaZ2cPw7Q7wew9m7vwI75yMqkaT6ra7z
vjlcMOTmmH6SuzzgWJktjWj9+/KWsvNIif7sAhA/NUvnhZFoEOQdgyM/Ze9F+Yx6
eWTOAiuJsA4cBvWh/es622wBuTedIwS08Kk8wVsN4td3AHA6DlTL0mAgMoqemvI2
sKYdWsLL2NT3CGzYlo7vKkg9daYoVGI94ag2DYZpcJrTpdjxfLATgIs5/rybRVUW
RujUj0QyX/kEB1lAFNoMrA==
`protect END_PROTECTED
