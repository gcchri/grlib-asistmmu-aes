`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPv90VDLiJaQII1Dkd6blntdo8YgSXLQgvNrJS2lVbFVQ10lkHmEjn+Lv+i5qEFc
bZmuekuTrkH+bfnSIHiwjgKqVJxmXRQyia19AQ/W3vTCvBzTes/3K0nJGUnH+eqd
EEQe83FqZP3NXkqH+UGZmRIhSl1f/0LhnTYe7b97zZHO73lKtIP3jWjPbS/DWKrS
63zBN+4Rv7wsfhWOmzEzjtiNpXrFzgQQpXaojkYRS3maFs4idrC1fK52Cnd0CDK4
`protect END_PROTECTED
