`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B82f46NP0IyFV8a5bFPrI3hZ4ZEvxvWAI0e0KufqgBkmTNl9KMyUEhsnXjmCYz37
gwBvzIPrFpth16gUGi+Bvurf4v7TfbkYfUWUx/hWy41IL8vKm7ayMEtPSkuDdpxR
1VaSqlMhFM8jan8/4IvKZFi5LCsOFT1P27RUWkW0x/tKvYkhBkDmtL3lHPwZfaSa
jIBic8WQfuSLY5RClxj2tXKj1k8FqvZxGdk6aNWtO8ZN61K2anCJ6X3b/OrwLpTm
AwOBAevvlytCUrPLUFNZ7X6pB3LADubCtrmeBUTMnQYz6uhhtZJ7O6w39UR1xASV
20GtTTp6XTUdUdHmQOXUpg4+hrnE9tNenOtwpOPA/eLC6DkAO6X237IUzikTV1FL
xEgkQbnHgdpqe0XmOSEiLcuucB/boQLRURwPyeK9q40O5UGPK/ThKtUhSSzKYyvA
SsTqXWh5vKmkzyFQagL96yVXFQTG6X7CzhJHz59Ao0U=
`protect END_PROTECTED
