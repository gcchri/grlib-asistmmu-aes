`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BkLv9lEuj8/xyXrpzV2UeHruHiVHbch4OwS94Z8JK+VGM57Mj2LTGrPPadToqRbn
xd4CA+pxB2BKFnZj9D/ua+bSIYRY42gdI6IJ8osVGu1ZeLpkvKATbzRzknhuQTQm
/vRzX9DL2RXTEpEE0mCmURqqvGJA82d4g/OuwsUo4avWa1OTigMeZTz3CoRu8aML
xcP1plfY7w6ElFB2id/MX023dte2llvJuZNyNffKzOHyk45YoT0U/Ti0MEA3i6Hf
tNLb+WxtAj+AtNezZC3aucrFa0RahXss6Ibdc/y7bc8aza2ZuawJ9CC4TycEASzq
WW9hX4KBOI3QX0TN5D6SHedNmkUKbTxFMxFaz2nuJHv2p+sn9Cm88CArmmysTEvc
vVdqhja2uFysMDl5ZpRgJKPMVKeg74z8ZFLBHrFSmy5qONbr8XDWdHClOdwwcRqQ
HOJ/Qx5QL4c8bBU7pT/OwsztcKEaTJXQqIcy8gOeWRnBuG4zsxaUT9WlHbNu6A47
GYiN2ga/asD0LVhoaVrEws29BMzBzes9CyJMVUBFMczZNxO1hJmo48zOk83B+eg9
`protect END_PROTECTED
