`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4INZmo4H4LTQ6kdFKJC+ecMNkgbqQqtmRteZpSTj3Y5JcwvaqE2weqEYbv44ZfjS
H34vCD5fuodRxOsUph4QqFvnhF5NX3YqylI/ACcpYxuURTG9EtNNWL3WnhxrIGlC
j+MUHal5P/9n107GzYdRRHEUegPUHfj6Pw+Twu9gyZvuuJwNAQxTt7abT9hMaw90
saY+feivcmQrGxYkBq9lD0esaTye7Hbc833pjdWXt5EU/wbesWzzea8aMOMVAF6J
oh3CY+yIiVVatqiqZp6H2IzoCp1GnmNbZFkg6Oyka2MJ3W/gIKmuvr37t+7WPMXU
t6wZ3oRPK1KjgNxn6QzYgdAlATUfkxQoVoSJsu4gZSVRUjYtCKbTwWWcsvn62/s+
gW+tfdpia8G/a3g9JV7feP57B/7fFHHr8WbNnL9PoPGUUuVXFuEaf0Gb0SuBg0dq
sqRaCOedUqFsxhGgJ+a8P9G9p8ZoAz8OvUvyWAo4jbObgjPIaDeVxgLz0FnOdBPT
AZqN65i/2YVIo5hKhPS8/dVRARnWkR++j6wP9hb+MGAxm015ZAoBf2sJwgRjIcJn
7uc1JwXGOjxplDBrIqTHmVDL/Vaj99HCOTOqVG77bMT9Zk9n7njPoDQwhfYfN4MR
`protect END_PROTECTED
