`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6rKM0JMos9HqCQ4vcVW4H2riiAOBBNxmzlIoEl2QUOWIyjUzQF9oOiViwMyIMNcL
DN1c/KrMsV83g9/zD0QWL1aZzTZQxc7X09Fd7LMHwvt1G82l7OfFe5rnUhOcmNzS
0OMeeqcbTdXjv3EzM93n+/6r1oriadk9NSg7zPHldxUcJbWjmJIESEOKe2rPzOQ0
qUsfTbHJ+v05RVifaqCUpG4y9+407WCIiMmwuKJw5vXYYQmmDP1QtGoMyOMLejdC
jmSXIX8gvtwuxTY+l08jVLc9kWjlrLpIUs0TdKThZ8mKyN81MPn3XzZ//CYRHmQn
Ow4eij3kOzeMFyeXtUGsQhR+lsL3aJsixSJ2a0iTS5dAfVRqrOGeXkqq0PGKbanY
G5rUl1g1ilsXfByu0rrqwMR1GqwZR5UXF8Nqw+S+7O2PGquDyPNXAxcVU7YTjp1g
B4DmoAISGmFp4tBZEYuy9qqZHrhT0/B7vj3Y1Gon6wO1QYCfTVl2wCW4P//9FaQN
xEWnrjgOcO50m7IRcab4N++s66qBlyK7g//Rny6GXMbxMSjD4tE9LTl2wkuyGyJj
`protect END_PROTECTED
