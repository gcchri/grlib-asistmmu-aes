`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R/ncdJwwYIpiqpQGnAPr1vy8toMyINPvkCdTCOE2+QX9seQL2Fo3FAccv9aHQ2zF
k2b9E93GWHKrB3j0c3meFQ/mAEizgpyEF9F/BwXWPkscWbc4RnDcfgYtd1WnOGyP
W9kEHhV1LzitB0GETY+5+73pcIx+QjZ0mAliYbYvQhhZURO/s432I8j0kV4revjw
tCTHTWMkXHfEYMDlnDUzaLlaT5EPcJxNQ/eYAeby33HcTbG3zU7OWWboGO1n04L6
41QacHCEBWzYdqkAq/K6utUMmMCcdCeyuVji5aNdfmWAb0BmJqBBJbwF609/7u3B
`protect END_PROTECTED
