`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e274JwpLvn9vvYpO3Y7mMseYZOV3SuxDCliNijmlDUawddEgFV7TqlUKiN3fxZoh
WQ3XC05f4dX+1u2g7k0iUm7/rspymdqVji6LaebpIw6utGupdPXhLWoTfSSlNRWG
ERLzypQK0T//ahB8bmVY9m390JNbS9TtfMfvMmwml1/9iacdRnSRPvEY02tGLkBm
TpD3zuIR3hN/OPYmJ2rmFAJnMJjtJuLDjG/EsdshnSzRPt16zRy8c3Um8SYOP04v
zK9kKkJ3mVUb0npAWloSiWOR4/DQayJAU7Cuh2muTURCU3j3iuUJ0tLYUVdfQJbN
5V0HgWvxjB0+P0CU9JnVueyueZZqs1gmsp0KC27npzl0hsg209emrMcGKTcbNqjY
QiFjw3mQ4wlnoXKLW52CmsnHdWj/zO3RnD+sA+HoOxT4nZKk4A3SdLeChjIVZz01
NMe9v1kE7Cyy34k57gPyQW2p4e0VPUlDlEVfU8v9DaASosoB26XjSEMaGyH7M2zp
A/ranz210ZgOoNqTJPh6a59zRhtJhw9x04XsvbPr4VD08R5roxdtOcpePGLWxRxT
OqXKkWlfT7YCOp6bYouNU+i8/qM7xmx+zDMeEgHrLnLC3nnLrj+7KZf1bXIZJXV0
vSHrji6C719luu8jZY4EJukheJ/ZrvNQ/Rmg0zrGMaNAyVZt73Yqc6ZKZv8zzrI2
36C5rgTYJ66KQBoU12c3UMR3htYgI1qLt/kFcNfxJwenY7n3dJxCtu0aQqo8nCZH
HUvBsJ3bwAeJ1+GPC18INeocZDrLed4p6XCIwhO0soAdfpoDOhGoQfQAkmqcTkR8
IiUhqFi7ilOFVDLgZYexQwDjdONrZTykV9oaz9DDuxOrdVeG0uTx0ATQixLzhMd3
xQ9wsleduz8cI//XcXbpon4KJGcEjHBtkbTvkRAlKgOcIRYGDT1JhAXHE5vYfc2Q
pTtAxvbo1u+uRH0j79m/FA==
`protect END_PROTECTED
