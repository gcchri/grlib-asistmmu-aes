`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hONtoC4F1nfRuXKwc21rnTrmMppyXfqb1rkCHLkEtVipr02AM8YXwafCKTxTI/2E
jndKbapwXOj3oLc9hQGXReS9cE28x8MmyuO0aU16IZvB95pHrzz94OoIpBYUGzSv
winZbE0GaaaDFiJ0Rpl7YJ7mRGZPOycvfMzfHbNF09cd8Mh1lbX6KvA9Yses1Gh/
ScIExfKaSmGVLXX0bBjlXvK04klZzCgYbFx27B1eKt7n0K20WdX94JgSwtpdl7s9
rd6MQnh6JYWb+L67Web3fUg/rtGfTNh9mNUyh/mAaXUpIT46mlzZU/01+oBFrIwg
itqT+lhYVck8PHdQwCsc3qLZeguxDC6IUJwkmiCcgvKEJcbNQvNAdvXC6L5FX3gw
gKW+rAA9ZKHrKayLRydGH0eSUXWnX3DYwKtwC494KPNTbg5IYtRAX79GgffLHD8+
5Gui8ePxFYBgYAteakEGR0y1q3RNQwVB26A5xum//8dDd0gTBuZgwS+gJKLBK3GA
Evw+d2Tzctn/Ohwyhk5WMb+b/liVJnv7S3fZUkAIyJWMHcF9zYAOo66UCUkw1zfL
mAdk0bPCGHwW+R53mAcaueFadzadypVJUfWDfwIM2giNGpkPDj7XtQyQJQ5vBxj/
21kXXStxloGVvWus56YQ+dvNL+5WDGvRpu0DM8Ru8UB0XXcTlSUAWcOjpU4/M+Kz
5A7/vVcBhaVU0YqxCG832MNns0hmTFcUmcDymp/QCOpL8VRy6PULehekEyhbw0PJ
WTL/CQw+3QbMqRD1sgsatB7T7TGSF2qM5QDg6m9EGq7LWInmNoI7KmSghleqf/Ib
zuoDQcf3xvud0ClsfKRHOPgc89Ea0AiaN9HNqYFAcw5QhEDqW4rZoh+OE/GUL+jD
psk4VzMlrBr9gTyqxKdgm+gRtWyuKieCUzdHXGgUjnJsOWQFgYr/dLrm6OEvoKDW
+uTXtrt8vHxTgHB6qCmpMajdf/a59wrWzKwENlaP/WYlQLkGJ9yPhVghzcX3vee+
tBEgzx4eEduLNjdROXlIl+4StKFXhF0FfAbAtbllM1esM6cRqbZ/2cKYzh8q1PfA
ZIC9d4axF3sjqHy7YbSaDh9G8KHV5jocVP3nfEwDr1XhAM11VuWUf6kescRWW8RT
UZvUZp9LkEhDb8r4yC+XzUomUO2ZofviCU5qFDSclI3vAiaUIuLdeDp71IQ7wSd9
E+9SU8XgNpBj+66RxhxhkkWVC0RnZVTd0aYYvocxvP4wmPF3U+AsUWudJE0vD1hb
5Jzg77S7hDa8L8/cO7SGT/tjDoovvL8YSuwvBqexoJNfAn/6eKYcB89e1m+xTTEB
6c1UJiN0qFN+dCh22uHAwtv62KSaPECu33yTA0bUhJ0Fds3oL5xWg0E6xO4p5QWi
rbKmb8sIl2QJJB6X7pe5C9e9aASqyi37WdGcoiuFfbaj8G0wieb89tJTuY9SlWad
9L1uTw+S4Y52xTcx+v74MPc/2sav+xkyQYl2NKWLvoEo+aIdGInV/h/NBe13yDUU
5sK8bc8XE5wnBfsz2xrNVWZd7RtUvO8122uPYB5RQtjtV5aPGUkzT4+O83H/6hsd
NVdvjrnLM5Y/lAND6ycUoD6P+aV58V9Y6z/VN6f0Ctsvoo2z3AkqZzHbHp8Hge5D
kE+3ZDJzagTXddTxpNZLTHBmrwzfCxBat84wssYtDqb1PzQw5r0mzpHi15RFjAxk
S3eV50UxyEPUWAbIA9Tkmq4sg49MX0UwRFTqkFCN7dvWKd61FrHr1sn7Xu7ub9Ts
YihFswpj25lSnkenLoUnAK6lE+Bp8dNuqvk2NWtyI99vGsu9hGOeNVT9eaTFhjl2
pHN4hQMaBESsW51rg2rgopdmmu7CjWlBX3FZ4X26dyKpesW5E02/7+vyMtRzVIMZ
kHH7mnUf9apij+MCNEmgSZ95Ok/OqFJSvLNH58GlxTBFCq6F4CY8URLn2qhEpdzy
FGY/jWK7JjiZMrCsNxKfxoMHLsZgtzw0WFrguS2n+W1YdGJWz+UV7rGdMCU9Ayrs
7TfN9EKPIlaz7YZcLDlUffyvrz0Dy6TscmbdLrKAKh0O0LUuAJV3iUCL9pmM3PrM
mvoJIrEMFtBV1sxT/tx4xb2Ljw5LECoZ1S5CO6DEkELwNbX+ItkhWqmFriwg1VJH
oxGL+BNH8DOl7u47ijpodeTwyNOX6/aNQSq6R1cSSHBYhTGdvuV6njtB8yuUppb3
OW2wvpk5h0fa3zSag8IB3hCQTP/952ljubwAKlBqNx4dw67Cws1xnXpnQCBaM3Pb
QFV0V22Nf167Tv02Kyz29lUNEV1DJUjoK1EHtPt8N+qhYbJ3a9XT9kkq9AnBnQAN
cCpCk44sKmj1lTPe/kK32oSlR781OJkZGwaKB+14H76hbWY44FrpUgNR6R73G4Zv
AKImxnDoXr6Cegxg+eHTg/r+rclFSve6iOsR+OhTVi3SrX64Yqd+Y/t+OZLQpOcu
gBMqVzyrixo6xBR0Z+sygBw2sahmKQE9ZDb/Iu7D5T3tNExocdIU8yfmUbyuZEHX
cgFfoxtuO7B7HMnEkbR3dFxU8xCKHXnAwxfz+ltO1MG1ul8JQ0jFgWnjPUiDgpMi
UhHakBpniA8CWz18hI05wx1c9eR0yiv3UkDAS/PSiFbz3X1cSkYKUh2Dauj5oIIc
pGgiqUmgGHngg+1Nl+d385ukT2escOXCwK9lu2vT9Rx070EhkEfnRAjiLTfHsW/o
rINTl9SzJI2xRYZhhskiI9OtLCspUdEwI7uhCWUFDs7N2s/KqTPsbZ5RcIzT79wa
IwXR1Wcm+qnwemEz62Ncom0tcHCbc24JV7x597eTjqeZ6qlW+V+arDaNhFNaqHCZ
++hZwnwrLSkGpmik4N9Nkf9GFDSSazgLHJCN8Wt8N9mn2YoYFwzlFgHU3LcVaqgc
WQKCpqSX+4ItA8W6PSoUvnJ6aUPiFP5jZYbuSwt+W3CPP5JZB7+HBJ0cYTcRNruc
PIzYoHOjXeOv1QIrwkAEDQ5cgI+bRa1VzMSFFQkBeSIpqPaEzzY5LjUrKin/s58w
Z965vT+nEJR4Q1VvIZp/dreVxiC1GaE79tryTc5sTDElFNp6hsSbsMFUGZ3TctPl
4oHwkNKvzK6Fdjt3QasOQqID7+nviXK0lkg1LQGu2K47KGiDwdvFhDNxt3VzXBmj
UZTsNRZKxiArMKOqMOvH7bVN0JBXWT6tqdcZPAu4XxcUSUJqAz/NlZJOaaTDy3fD
IMbBj0zwyiZUsTf9J8hr3lt2pa13oMPeDkIEZTmSGaW+tQDZUzq7C1Q0+XheR+8b
rBmsK5LQ4IP3aIn0SKYQqFnrqt0rz2lJXmae9OeHLgzk8jGDDa+wbur5xAuOHgon
EMtQvXo6bmH8IcBLEhuoRYsb1EY37PpKhyf+S9reX8IALalv+jcUw1zX4QQu0cne
09s4P+LcVPRVYZ/sMo5pRcaNUhfsBadtSw6uxrvcIebn1CYxbax/82rZWBK59q/B
KBAzDk1e/ZnlOmq71P3rvr86UdxJuH2ssfXpkiMFv9cQ1bMb1MPuKcC23trRQGL5
QUXO0/ldzsJFPdE4ODXQ1UD8lERAIgzjBiqQbidRVVAvk0ZuFJJw1BVYzCWfxUPh
F0VWubVGQ6erSakcG/IAjQWyPb+QmSDgbc1o3LH9dTutvHcEflOpYjZ6o1wSb1Nb
5xImjkjCLQ+NxpVms0tZ8TEVCZVHUs6r5aE4P8JABAJPPOoiuRo7pGfxoyDJRAiY
88pgZ8K2ERYKBwZE/6ddw0BmNns8PS+p2o0tTG5FGZpcFXEh/hyxNLzQNx7FDF2I
r/3JqR352iKZIrLlXoZedYx04P+gzwCeec78R9IPHCed49dV6MvCHr8xqNXaH9H7
/ldDN+BQQz+rtYcndHC3J0ak5pqXok5NkTwZI1LVN/BaeyD9qGy5UhxRbtgXVfIK
/GiN2friyBhqxAu+R6h7CaOY58/o+g7ySRh8E9mhXO5/k8pkIHqPESnNbWQ0JmKd
xVvyevC8mTJ+dRZj7qu4HWRX9QNAJwjh1s1TlLV66wfOKnVkg/51IvanVFZ4Oqzg
9qsBhNvBhaK7Wte9G0p9vrJ6Sm7YO4BiFd0k0ht0MJpgVKnzVRmoz2SMOaUMNQfO
RsJRR6gSgIHw10pg9l5RNBQbGQ/XW8oF/VCjTZVBSXm/zmbT1nn1zmArV4OCTn50
YeVMKZ6w3PcuoUxRoU1dKV9dFMKtUxFFvwc1Mpx4EHmqclc6ZzfVITPnD6u69pLz
ZM0E4csi48Bt+bzElUu3zD2czTw4xXZBIcCxwnBcdIbD0bUPyFH+l4KM6nYpltzc
JK9/NUG/16KLrtczusTebGFJ4iUDCnQVNY1QYExBEOH5gWVV4u6zvkjVoKDPipfc
BkqAsBygOb9/CqVRfZxTxhp2Ke9JQPa+KoCyhp9JGva/iKYDk/d/68WRYI+3vn4t
2KT067uRM/AbBq0xejrhSGkA56yYLR4KqPhWgrk9KbtI24YzvvrvcD4f0fSpiBaZ
Lt+vhwPT1uNKJBoCBYsGJyYRBluwi/wB8xDcdBLIlKzmREEyzZ8/7R0ADPXWhxTJ
5qyAeK3qIJufzgMAXJjY2R1iYQsQUOd0EQQWiy3pgyw8xBkL+fZ+ajb2kny6HlOp
zl+QsmRa6XqWBouFtoQoysn/jVSNSxhPH+U/Hqshzrr/jPydztlkcRwZXJbliu8P
VvCADTcJZngJg7fbrRDiwyesDbG+FRbfyFBoquGZQsaOjmXjlS4ogHHup9VeBr7W
34sNn1oeBo3lmsyAanznstPLWt4ofON36c+HlX99KTgZDr/eSJHDgsquLHobvMvo
Zat32NyOLvg80o5PCUUNGmiwlEkslBOvoEwAxBJ7JoFPk8BdMfqdCbEsj72cf973
Vcl5pLGxlRct7Rctsc9FXwbGM9bVyv3nIKVEU1qutDqkk4rHBzFRzOtRZKp2HEbC
WJByUo1WU8dw+mlVM4u3+GhpAhuJunpBpe/mA1WO5vS7bwxLo4NqDdiWwxvlRU8l
GI1Pv4+CnzbV3834QZGvcg==
`protect END_PROTECTED
