`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J6IoMIGHIxwnxrMeemhKo4yscCTdKgDO3TdcoCs1vvoKIZW9grNTGrD7q3wfq2wu
qVgySSCRJ8ZJ8u4QAoD7Q+/JufML02Zd31+4dcyU7fe1zHMwjVndxlTuI5dsgx2Y
Jih60D7VkHjS7DZEsDYIV6gYbfE5OIXODYTxwHwUJ4KzuNuadR8UoXwnU7N3cutC
sFbw/RNzG3puty/K/PCgZutHmoiiGUm3M7DMvx3hx+OdQIFfywrbMXpnpKKPJqu+
37MF3/eKiQTSeVOQaOD87iCdWt838Hd8MyWHAFXwkuzcBpluBMpTv+aQAp1dOYgs
`protect END_PROTECTED
