`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMJ/1NJx/KT2+csC51C+juGDHnmvJjq32dZyWVzh//CwTi4ofC4TDchnd97V5tiO
IXUU3VzgIY9sRHFhxY1wz6gTLwMXbuTVo5syB1/Q/p2R2Y88je2EBZOCd9DmZrOb
Y5wYvfYvOKSYx3mHWLb2MBG6zZ4gcmbb4xJdDGP2z1CYmlVWjH3zc82VeELyy6cp
9rQOLoYPSf5mYtVKjXXCMscm3GANsUyulVLnRSFebsJjl0fDaq1aCf44NkaWQlnb
04sRXVLAQIe+KlBF2IquYE72xlx5H6xhGNIwYu7mQK7YoK6ZqYH6/3YcnlextXt5
Aof7Mkk0lqB9rp8MEXxUMDxEApaA80II2ihkRMzC6gQd3SYOJul51FIOJ0MDRwL4
BxjhfrCZbPwAKHgRKdt2EV7CuQQpSIkOzD8ilB4Iyu5tlELxfZS6um/FGukl27N9
PPeYImVtVbZp1CmEbEJutxoJxRKWv22oR49T7saQvRUSQ8xrxR1+GuoAtzi5Xyfs
6NSTiJYoGSmdOVpFwZ/pVlbC7wR9Ev5Au4rJTanBbJ/DiBlfLpIS2bUKyRD+ho7v
cOPv86ZCcgoBMJIzno6Zb00wpTUNT3P7smwe6uEEXyurXCHIz6/RV1HhcuLSmKJT
G8voTWdG1de4wdmLUCqpADfjwdqeU1kN4Yo2tb5e2eJvhgCaRzqnsFJUyFATOIQ0
ocEhPS240RRq1skD3LaDGoQtQJ7SNmhln8JV6Sal/n5HhkYE+JUp1POJtuqoNgLV
sXhMK1GxaIKDKAXwpq2cmVyGe72WTw7lqnH3mmMtrMVqxiubbLB2K/arrEX9mk6X
IskjYXKlmudJIJMGua3NeY0A6vGonM5auZ7pIuoNDduJ7U9aTKSUJTyfuiI01fOg
`protect END_PROTECTED
