`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pKdof8phj3sA5iRMZhMjDLLBHTgZHcFdTi9G1xbmn8y5nxzU4R+tmUYob8aRnSzv
CCYHGTHe2sd5C/K+aQ0MndizIJecP9u2AL+KwlYl7m2j0kV5qlXrWzJcZ/lrTdBX
CMzRLmhV4RBL+TUWmQDnCNlnF+bIKg2BcMwcw1lJ1Qt3Io8q/cDRUL4hlLn+fF2Q
w0ctU5063XmdiDzU2zVIEBf5IszwK7HPz6gJUeI4sz5SQgTZJwwClZO4gy1hAYCi
8QdC4S8YzMGdOkTJ4DwB8445bmfAI9M+SHGOmLyiHRjS4CGYJq0K9eMUmzLRhCiU
Ciz8n3jLHhFqmyTpo7yfW8cfjB/63/ALrAhUVxektA59/8Y+Gq9LJg8CyulBxHcF
Htj+qXa3suhqQCFW1gPaRLKi4bR0l/QOLjk5mlmnW6PIxLmS9yJZcL6Wc8n/Z9A/
w9mL52znB20a/w/lkqcp5MdwLMKR5vmJzq3V7O9PWMohZCre+IS+3vK4ZCd/mw9Q
PHgqZ3g7F16PuUf5mIEB5pvXV7JxUFfwdHIxzS/fExxdXN/B6NtjqVVll1kehGtf
5V+vXFI+r8biHlKp9e0ZoOoKtd5xMVW9iIOqwt3QVZG07BQQkrDEpSq7x2UtlLnX
P8e5hL4unk429cnrBsRTzc/3SXlISW5osvL4k7jFPV0=
`protect END_PROTECTED
