`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m88Xt2yKml0H8qLJ7NZ0r0wRi1mVY8Zex/WTAkIRKjfWDeg8yQr8R5kUF1VVbEdH
n2R37FzLO8SFeFlLkp6FWcfjPr3FZOpCuMt9/h43X7Zbr4Ex4fTj5V0TPtU9IgZS
F+jzUOYH9S0w2SuGU885PRwcJoLQy3AIbuC7enNCf4ZKQ9zpU2ZKeoVZHU5unVP5
93woNVxUZXNCqyMAMyQENQ/bexA8yO1DdEEV5O6o9dAvpn80tQajxWH63QQEIiC+
x1wa4XrThMzJZjD+zSEG+lnRheK5GrNep3IZR0wEILqIEmCuz+cKG9QLzRKIwkVa
6gUnxJ0gyBdwSc7Om4K12HoP86Iozol3BRljvvvN5m9fFNmq4Pvs77khmgtFqegB
pO/e70JAZRR61UTfI1iHFU+p+ZNLhXOBJur7+zsT+XxgykuQiRAC+kuSp8Ps61MB
5Kslx9+uP06J7zrmGC0+MovHLVZ48r9825U0ExwMPVqWwOPnQbQgv4DxBMk1mh+n
+FJCHnVuJDDfdDDT+7npLT0lLyAjX0NUlR2J0T5Io1xO2CY32vHhRf3ySSP6c0wa
siZzOrApDVRdy5UrulYrmRkX+SbiY+0vZn2MaYuiIWXDac63ha2Q0WBxN8ORENN3
QprjvkeOH5FCMDB1Cjb4VDrnYPpV+vqRvign4qoHR+d05lGN9fltCMLRDEzVy3Ga
HHD7NrEJHDvRlJGNrMThx//JLGfkguRcCmYM9cUbpsfbu32oYLkqqcvD1VvWrgnR
sG+hN44zC6npKFe/dcE9VOmU7CbFlFTBunwkm1B+/c2N146QEvJ7t1Tw8/fkH4YX
elccLuEjNSuXyHCXGsvFngdHPvnjpye44FeFBI8buFaR20WQe9Z1Y5uS/Lv9ayz2
pLAfZ+E53eh2ZYVS3rGlcWd4EbrLXrC8UcEEJaSzMz7MgnIPqwZ/dtojJOXibe3e
8m76+198jwa5oJMIo2hrPsbciJQfg+1e9/tAic7r6SAaE95fvIV5rA6KkqPAb/fl
/UNk8igtkklMeitYt9WPxnWjaAf6FXsykRq8fZj6ZCmY8nY6Pxmmejj3O0Qf7NEi
YGSzO335AyygrnMHd+EWRp/8S4GpwA1ZRME5Ssks0519FHaaU48TmmOt1gWFyXGd
TV35zt8aKn8AF8+I/yDW8XrmS1/Bn6sk+hmP5MxpC7/Jg7F+isfDHJuoTI0zsibA
EC7ggqbmaoZrn4+GVh7evZE+4wmE5eDxfmERb1LlO9fup/dHAAoOjJbKye1GDaAh
hiAd2CHEOVAZaGD80IBOIp5U/9bjqkVsr64qzXpwYLp1vzSNZ185FvZwIu1xWRVs
EzVP6RIARVF5sU3+iT1ZXix9NkrFC1C6Zedx1jSqMaxAKyIk03FcFMu2UdU0zAMi
H4fdPkwuzeo6QBrnuYvJ/s6Wgqsct3PSs4tYS7bCUyUkM1PXe5J6zzELSS8TBx9W
hq7jPqvXB3iHq6eyCoxboGepDJD5URkRlIsaqvLlXQ6AyfubdgeV/IBdr2mUv4sB
4O/KeRf7b0pv9yuO8bgAPwsNL5webBcg4mrFpzb1C8rgx0dgOzbjoHqyn7z7t1Tp
+ILJShxXO720IghWoCpMU757pGlWtORu0lP5Cn8U1uJHWklp0AwYcYZZmakvBN1D
RCa3qNGpbWAebI1IbcjDSMIEb36EXlttnt/nFZ/SBRoOdna746i5rMT8lO8cF11G
IkY0m62Q7Xlp6XrusjiHvBFBjF2PUYxRXgg6z3/CwBMwSs6cIqs4hF2xsA/aDhMP
DC6H88oGGV74Xsizph+fUWePS8sl8VmzDax5iHL11t1lSQ7gPbfaSCx1a9I5pCAc
HD30cGeMwQIVjgqgD4tyjpGELSstuw51JyXy/B876DwM9yP/CcNcFb1wEOdCuwAh
mlqoSzmZAu+4CdEf6kimjEhZXU57Uzp2gvoRjHJX5nMsNH4xqFhc0MxCG6f2E3D8
5ZsGtY9V68ni6sYX4aqZRtCmGS4aboBzvrqZb1X0jXuArDkaRBzj0SijvBAowGLp
qUR32BXurrLLVsVAy/t9p6kN17jaZz3GAKXWjQcnfNg9lyTT5Z75j0QiBfFiqirH
22lmHhYyY4WTvHyYuGjB8ux8i2Vn8+A+iENmmfuRftx5cX8sxjP4NVnlNxA2J/rP
NbpjKAG8E1ST7ImPbUR7HmSZdvzbmeQxMsYLSiTP7eaSNu850yZhcW+/VTKsVE48
bKz/thiMxoj6Lu0tP09lit0bDkIVY12cH1IUwCeTtVWv+fFO7Bf2mFlrQEHkh1p5
PCo7LCKPMMFpT1caOgjc7Ne5IQiiLRgF+KNeho8SPmJ/ew/sQ0hEcs5Y0fMsMOQD
qRSrABg5VcYg+yjEsDlL22RP2tjz8BtbI+eF3dfg6UZ6bVJOdrZiYjWrGfXkUmfh
CTVZGu11x8Z2I1lTO8ecsjEaiAr5IFHoV3tZEu1FiV9trjuBRuGbzI2lRdnQeyeV
RMkAnr4ToRDr4ZUgnEjqeODwvpSslas1UOHs9ZPoVtEQpRVUpcu4dVT3qvwZ70vR
WD6+2LoiLYV8+IPZDcbX/BzTZvmO+w8fjmo07zMs/J3RFksL5S66GrLDzH+5mUIO
wT1+acgua0Uyad7J2aLHKf+ij8XsAKeckSGAd+Yxp5aMMakRTxAL/O8C5qK2i0PE
A6p2fNmx7x0Poz2+wSAmcC6Uufm/FYhArYykfR71ycIFmKszfe7+AjZfxXRQruLr
GUNq7fiiYi3qIktI16aGV70Sz1zFxtq7GQQUPPQJlHRZomUVbWjhrc9vtpiHSJUF
qk7qov8addFznUUyizSp/Q==
`protect END_PROTECTED
