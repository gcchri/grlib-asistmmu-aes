`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdIKzbSaLm9agOUp/SJTqsoKCRax6xc+3rEoSbE7HcnvVPPmB1zBd2meu2RJ/unm
BRnNdufokfVgp9Yu/Oaf0+N6kHK/PvTN/d+iw57qIdabIUw7TrWzF9shQrAO9IIG
tKHcYh6el4nYP9n8CcrIDB6lkdeR/1I+5Wa/tF19mCRMMWlufrM4AAsardNdXUx8
r+GnyUXvQNVIuiSCafxy0uqvNJz58qgvQJCe3qXZT/9m81ugksKMnT0g1+iAR0Ov
mkhhmySxrJuydzptN+tnIA==
`protect END_PROTECTED
