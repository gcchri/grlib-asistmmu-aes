`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DOBxOIIZNE+NXbaz9yCo+3edCxVto2nrdGE/weDpgq7YreJ0YKpbvZDGW/4tug0Y
d/r3iogP1Ca97147xNsOhOXOCbBRBXDPyDtMGt/yI5QuGfjgCI64P0Z/qich9OnJ
NDVtK0QhJ5w8ikfE4+TQNMBqc1eA1vtBtMN6Bf506vihICfbT4J5S8WQIsFtGhLE
ZD1HIc/SNlF42bvtFe/hwuU4h61QXmI1VzX6HyZXjxOpnko5Qh8cxbg4+R0pZ7bo
zObdytsUzbbReflKYTCpEH4LbgfyTbY3E9iVnqJBTU26P+ObbOBjRfD637tgjG6W
E2/xUyweQbeqswNRZgD2lcRMj3GwLRtP6r9Bq1zN2AjmeZLlCzW+1I+3i3rvcS1M
eN+h9D0EYNWih5PayfKdxoDA8ob9bIBvuyl9lAc9PulVvCiN+l0GDYZObe6zTs3F
TuUxQDalOIzJtw996IuFUfyLVoSy3q4IfvrAAX+uzHD1QxaX5YAu7Yq3+TQo/iQ/
w2AbNm5a4Z8IQMe9ffKi5ycEFbrO7I+WxgS5JZ2tgiG4pTBUsXU82KcMkZBw+7BA
uNQRsIIaRpUwRHtyQJWuwY75dsOtvyDFffzG8wDWrYJlRuku1mbfyfYBBXf5wPcl
UMmeQNuVwbt2jezbuF9scBVs+wqR1epHJf0JAAnVwGxmO2AX6IlgAKkH/YzgW9sp
ZDqy0WJttQziruhwTSl1T8AxumO2cawVYorrqDRbfduYyNaqfiIIRx7KMXUjvrEw
ec0Pk1dYeh5KB0Imvyr/fgpdJ7BrWl+h59hm0lsBNHSv7/j8VkU+7rQ990qBwYBg
YI0uDUmUUeVHGFvAVucQVzWo7EVeVXNwEGB7CJtWJ9ZHtDGCO13k8Max/xgkvFfP
Zs034wv5TiwtnEw+e82pupwMugME90YXwEmHKpehOfQCVkUblVfV0N/MhD9X7kaj
ZNS59vEmwaYPS4Kl4kO0gu1FbgkbtREwk1ZlpFzdnjd7qyXq/dDKj7X4atxjM+NK
h8d+nQKJhfcsGvIQyVdFaLoFP78krznkcXLH7/qhGbbMicjmy5UrwAtAPnDyfWTm
EoiIohJUoyUMF0ffr3wU2UDTCjRvzab1ytMjn4SO46+as7Ez0MZTXPzJM9bg6Rpx
PZk3IH4llWJfNXPQjeMnoyWUYv3QthxfZLqc0ZuxT+oBaQ3DzBb/SF+otQtgxzrJ
xZQbtTxLSck80OyWCjzG7V2T5349r8Cy4HzJzrECkEva0+p/DAtgSHP5mBPw0Lwp
CDVADSpSxRPB5itOJZipf6UDwDbLZaDdsj0A7iaZluy/WHOjt970wzb5j9LTHttj
XJ0XADEJI+DJAeQBlqpph2Fo/5MiRiXFbmeLk0PcYO9FMz0PDnoVrxS60foZw0Ci
aOLaIiEpC27Mgj5OHX1OW72feuw82/Pr6LXhxRgZiPfewzidnbOGemK0L5HrdSnl
m4q2b25dBJ3yM/i+wtaGmjQ9izVh20sZNhtgpTwA9QVswt6vZc73ul8MCBhbtpB6
6yNRP7FhdKfCsNybpsvUF7H4Uwi9eyNSypwIlSXLGT/+cvLLuWUFK+hst9c+gZJ+
CLqLPJ+F64+RG3wePOtDh+o+fr/IGDKjWyEoGeuvArgzyhLNEEXBUs528+O0bXxe
cJpMN+22GrKhuNCARBihDmRzxeHTzYDEckl4lMop2ZQLTbooMem+brTu5JA4VxKq
aAW8hiL8lx7HLrVfE4/NIDZF3z4nVBbfWHpSqjv9AepEchHgrJcG5rDDlXWni8+j
uAlyE/0Sor7MqDXEXTUdZKGF4O/h0nl6dDOuCf2PCNk1F8o65dpX0+JrutK1h0/l
0CaI+rOUXFSMEMK1XVn+cN6OnNR4wLOdUqp+gdRM8vQ72r1gIBTlEdBPfWOpAJ4+
lhy9TU41b/XHeeIvDBUWtW1Qj9F3Mv4729j9qJ/LJKyYrJsyGHi8+4d5JyB9qBpB
OR/MonTMwLvvpstHt+RrHOnXeWRjmJ+dTXvu5j9PQWTY2X0pONgpCkjCclatS6LO
gbtKR6opx3MC3/C3DcO2yHRyYMY5S4XACpxAZDpLt6NwybeyvClrmMJkLlsKA1j8
YnTO8ahTxdTvfu7BO8aHCPQyFAbxD8IXgUIjCKKn2MY=
`protect END_PROTECTED
