`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LHaFjDhI9nPF1WN+AlhNEvDt+AWM1rFbZQqwPqgbE/WstAIKtVYyV13Mf5Qqe/4J
EtPDfnXXZL1KFbsdpy179MoMlcVMWjIUR4jSiOkaow9qpLOyukIoE8iygD4WYaLw
4RgoZ+NMBwSbAlynGu+R2gPnDvz2JQnAqEnmoSmi0WKb6bxr7tR4N5BlAKU0YMBI
emfvabvU/ze7jPCE1Zs+NGHtlDWYJwrNqc+NPbw/YL2rIQOjEB6HGH3gwmTqCLNQ
2OEVx2NR+CNmNIH3tbnBroKphiEFK5SUCvjv3mKkCwTyaVwa8oGf14yMgxy7ifsF
Jk0GUpENDEnM/rDl/foWVaEzNvLG7d472+xwlsxqR47kfovcvraP32f7sOgbhhx2
yv4THAMrgFFaWTx37OFfn77wdpYKJOttGqee8pqbNrBxZ/Iew41hq0U/khUn5Rw4
r1cLyvybiOG6iduqfkhwiq/FBZXuW9bY5o3ipP5e2/eaWjnaDEcsUwNT+tGj1jlE
9bW2N0LGH45ACm0/iP0qK7qdgg4K5fJuIXM0yPVFxJHpCAhH21KouAgJxZaw+ANY
IDjD6aUS0BP3axPv/Z/xBQc/VXsHIk+UdBeD3zPRoQAIVYhyaaFwcskauMnXDZiK
Ej606YeCHFVA2ijI9BMbgVP8L22MPlTQLuuOpDc0RLjzmNQmewsPXQlYOA9vVOzK
tQ+RvFOufGuNsTbjB5Q7crsruV5jW9TBbXl6TmG2NpzQuzYZZKOZ4ExHtRiuafWA
IPQZvYQyxCO0rjgmhMC0KMpycW+zH7noGRuEoW83yclSvzWj4pVfN3dHQMRyYEIo
HAGTO33bIEYLhJjhI+gkKO32rhlua5WbiJtYqMLlO4/fxqtNSb5h4G+gTc9i6v+z
uILKh7i0pncnooq/Wxk0rGmUA0eEfb/qJUrVTB2/aXGyFMjLZfWRGQGTySyR+v/X
7Ow5JERhrhgj6PGZCw3BqkJ9zdOo3oVhwgnYqRkIe099aGEU3LqT3JonhivLNDXI
olKZg8b990ntHJTzxGO6UgWohJ5wGITaIbl7+yGAfhVyuFibryHC+tutgiJk+qsM
roCCHFdmi0Ze08m5FogoHFT7O88W//8Dt4L8+2xc+dIGbddnp1Ou0/+nOAKSVb5F
Yz91P9PHCLs6FbdzVW2nfqlQtmt8ChV+Es1TUTDdztSNRqPcjTyY7i/2R6dtU000
Bkk6pJkznhofK0Ms1YrphfUTIgdqYnNu+XjDHPfC2WTVgL5FiU0T/bUXZFRkUI5L
GZ1eauHPuVIq/DT258AXzly/eVH6ymSyCDxMzJYKP8Q6z32KK0ZlWG5AJVzsTAiq
LkIUPrqPU1OEYvdNf4D23nhjQgQzjHrdIrSrMHA0ccqKJjG21JM0SK6OQu/Kwn8g
q7Byo8MJDzzIJ0vwE1XKiiCtawayOoNU0iYwow0Wk5mz8OQ5v54PRPTuaUeHnrUb
LzTNTd1AYbDo5pZ89NfVZx86NF4lyjXtx2zR62rNciYqjU9jfBhqqLD4PC5GwcE2
1qLnAKbMAG509ei9YF828njw3Emy+/sc6Eo3Hs6r1lSfw75ZKDipTMMkYwYB7PA/
Dv9ViLzdvZCHBgXky8Pf4WRRo9VCtBsnSzQLEMPBx4PHx44OLbw+2xJ3jeN5mJGg
TSXRBH9wxnQ/sXndKu7gskllcxI1NzdynnJgWJAJtDQ=
`protect END_PROTECTED
