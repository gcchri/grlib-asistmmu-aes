`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3sqSYMs//Vkcg9gfs+P6OlgUkjbJir1wzMexN03tVBAQjJC9yrdqJNKg5qZAwNFm
C/8Rgq6Ap15VKaU/+FvWkzIJCM1se4/0+EnaCUa/v6sJ2gd/mxEKlV0AvrprtEUf
mzUjNOqrhv5/GabNG2L6IrQImX5N7t4lf9hB9INNYY2l1+SNONbMP4vXOIJqyW9h
SL6qx4FYaUk6PhmPP3diFe063gkl1HmrQjjyhUCdByxRAB8/Cupj22SSEgE6le0+
lTcLpN3VsD5uEepRN4WOo12cbCp49IXarE4R4jFKMJX2uPODVOV8DnvC1IOKb68K
B2uuI1mFz4zHp4SmPzGgROoEAUy7+v7ROxZ9bja5pIAg23G75hBiespV6rvdmb2f
AyNB1kn28njjvPPZn40xCrj7UahomG30oIW+b7p2DRkfCtlO395P4pW25sdUMPHT
dAQGxm2lPyA7laEvIdMUHglPoujeqTdrjew+1D1d5pNbU+ph//FQfyzHCAfeEtGR
oqC1d1KbHZ3HhIlFrRsULcAvpjaL+2jCDT7c1wP63haXdv/WyUFczcaIOrty8/56
h0/Y1cRsFJx1/g+rWJoF4u432ww9ppoOiWyPREsNlq3P8VRp4jkoTn6hr8VC9Dtj
yMJyHL5Sfu1PL8VzihANadIi1pQTTLRt+B9JjDeNkhUZGz8BW9yGfnbuYYr4uk9/
flO7EdQGjcFq3QFA0YseWQ2LwoJBJqKWp37grakozVd3v47H38yLCBi6QlVcRFWg
GRvZ2mBCDJ46pfjuiSfBlprhYyAfO9cKPhd12T1iO9JPg945tkuOBZjgdxCoQVef
LaVkU5zGPDSjOwk2S2UVV1dx3Tb/yGlYy3Liyi2WmcncUQq32x2gTxtTZlyE1QWM
2ntnfI7gaEW20a38IbHGvKtvMRYCHG7zbciEi5r9Edq6Kwd8zReB6cShxwpXikV2
`protect END_PROTECTED
