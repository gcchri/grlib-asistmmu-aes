`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mTLqRqbZ2+6df5A2h72jLkR1eLpa27q31AVWDyX/7nAYbEeDbBLShA0DtOr8j6qU
7cOAjDiX+S/iLoLVNP3EiaAVBYr+uyILhdKCmzMTuMEc06x4Q37mFJyoIyqIkbXa
J1vto+VLE9L11l0WHEtPGTu5P4XBoTvWaOg0XdFQKnW30pm6wXBAByIgPmUcLSZY
+BlM+d1pyw23195aHwMa2IT2GcbooiqMTGXavNm2mq0f1V7vcfJJD+mRWguP/MSZ
6n8UX1iuqKOxU3wRDPBo5Q==
`protect END_PROTECTED
