`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uAlgT+mfim/W2GhfCRlQTR/rII/wdIvrVDuT9YXjCbBlhbXDvEs7t3TVuDHU8mnG
lG+LOdL/9fGB60oQMjNdjT7fapLIuwbDJrJn1HgWGizQz0pU/hqZD3XAq3izwX4L
JCbsLp4BUZq+gX5dRt/oKYy1mx6THuENd2NY1uKAyoyH4+0HW3NY0UB9VKe4cRia
5j1aGh0cg+GB/Tr/8UzZ28+fu2rfO3CohghL3IcCfWqFtIqNzG9qs5+k2qDtAWZ8
bSaVpXVEGkyEgY2Fvce7S3XU6WCkcxIsX1sVPh61s0mjEJd8ZNi5v5ay9HbSFP3W
Wt51SjoqSHlSn0H2ibHaj2WnOA5DnK/UqmcUZvW8W7anB4fidgdZpUzr/hcCuB8Z
KDBpxOzYoOH7xSApoU227g==
`protect END_PROTECTED
