`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hvfkJBqc6x9cVoWd13O9dREUCbdGHm/0caygrtm6xjUTXVKisKHtvPJmqyfzwO+
7Pkzd694FRuzQ+WBXOusyZpmQHBKqVDUT1S0S0eIs30J+bsShE2E4jD8+mItVnaY
A/eUfXjO1nXYvBavdwbKeL3v5hD5R8JjTxfgegFs1LK4w6AXxAgMuM+2xqNPZcok
R2YVClf3xwErYOGEnfVdfMFpqzkUHwXLpY4f7keN9H1nsOtbWf+q2vqaRYpBmhJ7
A05dFNpj92Rg/xMoByd6HxdoUiwngTBaU+CQNJmhf9eftztk5kDlzAhDsAbY5YTF
k4tGkAIIvHW9AaCVsO72PzxAD0NuznKxEaYAuQWyeA+VXtgkOtrvyr23vyFm3+uB
xbzEtkP8JLtmZWNFSk1xsg==
`protect END_PROTECTED
