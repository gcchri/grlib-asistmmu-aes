`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOcP5FTPIsJh4kw8NghcSC+NTjCesl7hJu+eLFqJHbZm32F+u4Ebk67maL1TKl38
jc+law+n8ILu7M+Snr/VU1yXCRlnH4UuL2G0UWFfTJ4I8fgT8bds2HbBgh7qBUrS
e3JU2Rso3+apszwk1OF/Tbd1/LhG1fG+oJSpsjYxBufshtQ5vSaLZVARe0DG7XkF
Jn0WObUI3jutg9cvNa1JJ47AuNQsMY+IqY9EWSEVgGEiELQQ3GcibL9Et+8NP9Ds
WqqJ7U7945+uxvMiWt/uNUJk+XUPXDhIzt1FEO/2yhfBGcx/kYyjKh2j5H76oZ9W
7EZmUpqXAIvAsD7PZVsF36Do0welsvtA+PsRlWneMbrBWhuMHa94u79Jzf3W4YFB
hIMbFWusdaeDVCO1VUhtN29HOJuZO6AwQ+MDONYluIWUjk/peQs9Oh4LM7F/hmzR
b+7OZQ/O+LDJmH/ZJp5yDJj050lOUeXV6D9k2j+IatQ=
`protect END_PROTECTED
