`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/CQPvuVh5bTM2yoN5ohTGE8SsSSl468SoXfUf8u7iprc4YziCgx58iGyxRzq3kn0
ZxvXHi+Da+P5/o4y2qNXdMo6Pyd8hBNelwZAVfpyi5IejehtewzX4W1axjbYIM3H
+YrGWTBOHNrod3mZ7hYv/zusIQ5qogQfAKQJ+YTUoInk+eukJJt5lGYjQj/nlFkV
QOlrMhWk9V4VH1uWbiBvPOgdSv9l+AI21sdiZTOHAL9zsQ7OcYBBBBWOcQeNyPmk
517ducuQiOAepxbDxGPjYECOGDnPTGExGIkWmaRzrpUvdv/YGlcejpw1+G6KKNHV
`protect END_PROTECTED
