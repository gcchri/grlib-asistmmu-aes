`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lzjwFDhoHdOVXZxmD/UmWnxZop+z9JJNyED3rPtt7piOAnyBGol4UfPOfxtaJz17
f8HBDj9Duxig0VtzXn3enbmpkgaQZ+swz1Hn+4fd3svytLSW1RTsqMKyILFanDvH
XE5KjweDZYj1hJfNYtSZyBk7XW2CTvTgBbMiy5cq4FdeAsHP6lk4VIkitAun7ZTH
m1TJ2GFRRNtqlgLGUBXTCyzkW+1KfeaQw811n/rlpLx+LsZaSM81p7NWe8jOTUWa
Y3jUMobzniNxSUNlI+EUO6e0yBicdYW+Jo6LECp0KoE+Fg9r82l43bvvu4SOa+DY
PPFs3s9mmTDY3GkhQpR6LsIAiKDvrHuk7eqrVhnAGyEyheWpMrt4kcrOZ5bWbQLK
qwMwDbXoLSbY4lCV08ypsshXiGjTGUhhcFFG+EVRKDCGbrV3UDLFMwPf3oIAGZ+m
qASpr6gDZSDival5PwVPQWnia0SHTId3a4XOXwQWjiIHmWGK38C4nYfqQ7u9YmTC
Hvz99vBT0WIxfRLdGtib6MlqQv4RXPli37VFqWRGiEDVbfeosMt2H76dgj3NgDSW
t1mum4A11odPKtysda9gvC0fS0sC99gm87+RBVxUpNbcJ/yJeBcYg2s1Hmvz4txk
g3d6uYJu0Jd2leepknt6EAU/G+tr2NWnD2Udxr3vmyTQW3vTjNkoFPQmOicfH+H4
X/SJCmhCf4w7ZiYxWJeqJ0gi6jUmrf2nWvTAO0jmt3i8RB4gyrWPdfD7NFdQgNkx
4ODeychrl81hiZWY+d+1V23KkL1RCY6vp1DjVM5QCPx/diOLwjcj0UXDD3D+cN2v
gmJ6Tgavys30bwFE+W0xVw==
`protect END_PROTECTED
