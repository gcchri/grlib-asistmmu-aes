`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P9GX1qbPmPqMSyFpuVj/lnOS8XCNTudkn38gjQ0Ms2UXRREynJTkM1pnBHWE7ErQ
NamEXPdaflThk6e9BEPPWQjF2U9FHKsPwgRUSVFQFP1L9ueD74xTAJzcNPx9TdXx
iWDaa+ukdtUILm2fSiXVkhpCeTnqU/FileyHCiRMYl5L7dRc9pjyDbh/NeA6ESnx
U6FxOEh8pG4p37CIIVyJAEbKRIeLarDbgn5vxtZyLViyakM8iOZ3hCHkzilwR1Nu
HkeuiiSIAViaI/xEDqJs0VCVQEO9o/mAR/WJHiiXMUS6Ki4WrTBb+ETQ56xe2EK2
nU+hURwrf6v4383jnY3u8s1YOyuFiXkclVsbuvpLxt9yQvBW5FlKJKKdquz5gacQ
`protect END_PROTECTED
