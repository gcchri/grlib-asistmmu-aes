`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INWmwSh8FToKXR6N8Lto4wqdDCg+59Zbu9a7MdfPNh5PnDCkaTvyHfqgVUH2SiE3
lb5hEtBT+D04hH3eCaEEURzmfriOgvhAimq8I5pg6p2OcJ2MiCpDUxZiEEA0oJ1f
vH9xZ7GL6hIcHHuymRMB78+LdwYIdrEN7xeUbNojaOQSGdnWM6Eezmj+Ri0ZPLHF
8qqV0VwGiBsqYga42WSk8NBA5XDhRMC9kRdB/Ds/EfbtXdYPtPsoRA6jd6tWza58
ZP4Gjlqpu+v5OlAMEPNA/g==
`protect END_PROTECTED
