`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZEu/VChDcq7wEs2xyeAzkqVOOjAAvaZv5mM1jpsL1I9EQxj59O91sTNrd9Uw/Tya
vXIy+C58+9Z0xfncO/zU2ISdew2CxSL0Isq4VbjvB8YYDYWKxLTYmv6bjl+KhEy/
5JM+f9g6lnSYBQQZoVCqZbXJVvMY96piU/A5CojbBJGeC36yCDwNZPlo1B+45NMV
cujb5NdkHzI0gdW67daqyfDE1+865gOAOJNh+mdUZ1WL9uCeZnV157m1B11nF18m
35luPbSJIasouEAoVj5cjBNrTngz+vF6kSC0ETOp/6/TL947Hu76Qo9nAf0QnFxA
6TT36eDDwoUyoGypcayB5Q==
`protect END_PROTECTED
