`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AnwJzId4V0JBQc67NXOdzssqWZ7QzJ12UkX3OB4pKb0+rPuBo2cNGABTwT7kicC0
q0/7fNzk/1Yho1YudBDk7gw3ZOj2zuVhG9NUeuTY8HD3vn0qUM1SWE2wukDAO/4P
3GqW7/JhCaa0sfyalg9h0hijhbuJDzsJElhHCIOObYW1MjOFJtA78ynag51U8NyT
o78kKVdjLfayYLHVJzDEf5/USaTvqgVfW8gmvPcTisdG0O4dIQBw6PKGMOPWPnTh
Gx6vK8FIz0H5qMeAXcOFqoJ6RObLomG8ay0OB9xd/zrVAWSs4l6rXXghdjnEZ/+I
2by78Ea62waIB8/4GVm/Zj9ljztH/r5mgVMQf3RXL+RBjoKoRLSjLTR8+oDmfDzL
iqPSGfOLXNV/4KBaovS7BttvwA3+H0Q8a4QogSpi/chmZGbSUssQ43qaM/sWODjA
oHW1uEzS4NvLUywgmvRiNky9gku7URfihQqDbk2Rj4H+5EfURF77V9rcVT5ifCQa
N145GkLjlkJXobgRt4sbKLiqjHnwe86zjWGdroDiHGgsTXwO2NtKyYwol3kOgQHC
F8MghXcc9swADmhmG6ydKnSMrO8EEx75dTDtfg3d8K3+X8o2IHRtbaPxPEdvZVEq
yXM6MQ8XqeKbAwmQbjJ09A==
`protect END_PROTECTED
