`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1UCTeetJ4HN+WPkg+RZVwpVMNCFXMZsHUt1qW4qGeV7qUa4QFGWWH2LMKWMFOfC
QtLaRjTtT26+RGDE7iYCft0RKc4MdVz7DSLk8ig/F5bCCqvWvq4vuRrf+bsof0Jf
KttcsvmbAgtxQiu6NmydH5S8RPfkj2KlLriOP2ABfK+fi2LfeMCmKFhmcchyZZPy
mV7oZoNWzeqyOZv8ZBxeowEZNd2kXfOALOP6ilFawiWaYMuVVAqsC05NRGeJLsSE
qOT1OqEsYZySzoGWd80P5Ig0OGVk/HxUZhHhl2v9susm9BBHby00iLj3ckchaS2H
863UEm18/ANj43+JODipZmvVaG9A3q9vXbuoz7vnMsU6TuO5xlMUcPDeJ55njTZt
ZeURyXoZ6T0KCE1TBU2y39lBFsAxFMVTPB7lZ7WIbpIZKjEMvG/1sw32pAFr3eyY
Gl9zJURcNHpGf/8FmBbfWtcVUA2dctT6nnVblSCQ280TI7wwFDUcnvR8akFRbrEH
Q2jR+krfxSNLwu9Wo7haiFId8qX2NTOVnk47WdNbQPXLEh6A8LVZbis5V40lJAWm
Vfpjc9DSJR+ev6y7bKGq9MwOvwjI3vfxfluUk5ioQLGK21Q7VgT/OaFarEAysCtu
ZHN+BUpDF/0oAeGUBcyPaJuQnBlBkahE+Aeg83LoNEquBugDRYkhOEW3gwMMuD+M
qQWgcZotBkyA9iM/mgdB6TFwIRhDQ5JwjcIVAZwCG0Mf1yp5jc93vlBGU3BISJIP
AfDSk3fCfN3SB32RI0mUuE7S8Up4APm6FOwRnbMKB5k/3Hg9nCkkpvHJoBzMOvnX
Zaw2WKoklvZxGGICTx8s8T6s6dGAi4MrH734ph4uNWmEsPkAmjDsZK4dreQvtoyH
hKmhe/aB5B/KTzK/xDlKjJKR+iHMl5bA6kO2bYeeOSWSDs9Wm4EWy52K53O55zlx
HwbCIRtpGyMCjcgtK+3JWdyRqUMfDaCrJpAzuqBOJ047OkxLqh/2nJsPtMnYZtYc
`protect END_PROTECTED
