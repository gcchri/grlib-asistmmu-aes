`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+2nXhKFv1pERGZHew7kSXFKSmfdhJkT/x45QisYZK3zkjW2A/9kRBhfm4QfVti+2
xz6kK8m8zS5tsJDgrPlb1VXRodbvXY0b7616kCy8gT5BvimTSoqxtTh2nUC4HFvj
UrUcaXspPgR2rGhaA8gimUoOS3/em3Nh0XRps0n4rmqVxRd/t6SrSlz9R+VL8li9
QOisBBVPN4oLNRsYA7BwmTqYO48uYsGbHbIkY31Yub1JQ1k89Uwb3J7u2D83Mi65
5nqZh02Uc9vwbR/nPb8Knc93kLYZdrK4Wt4Y4SIJ8U6RW75frM4aVtrTcYpBQshb
aFh/CUdMFRrKUUnvXg6KhGFOOOR9YCimoV5EiHqmUWnqdEgcQM1uAIBLju1V6owO
dKiYkw3JGSyV4dzLmJIzWUXj1YDwrQhQt32OXg6Y+z9xZ3UErfG2JIbsXwSq75q6
1mSxEXvgJgETGTnnmOyuawMSAggjgsqVkZ95xe0Q5YNjz46/i2Bh2O4pvL/FV+6/
ou0dxJJXZVMVToozsGR7S1JnztIedk4dNHWX1Qn2dUHUMvp0RuSx7pQxR3bd33DG
Q1gQVKYGlLuf4Yot4y7J/oGqeegMaudGcGAKW/bJ3gUKIy5DOTxnkFmIPwOfbKfY
5Uk1voRXLYhY6NB9LSXkYPiNo+5wOSJBQWt8SshvdQO2VT/o5MNdWyTaua6UD4Pb
9HQic255KUq9VyzLiodJ1LPOmqmdh1WYiXfz/TrGmaU6L1P2ximosOAXgAyX3UrM
XvIkEKuZiwRE86aedbPrFxYyrjZ8b0JRBD7MTYEgCcwIQgxvpvEr0e6XaZJq67Bh
WTqGr3fpq1z72yommgRz+gB+jZqxyqK18OigdtFGwJp5pVczltXH2qKOoBqOp7tH
S62hpvUKjEw5/ei0t7GF6falAMzX+/udPrc4INkk/jhIYR35nOLhYkxOBWOeuH5t
O3B1owgxs5j1ecQf2FxneKCMI1aUl88fJgl0sK7zKSpRzdDoqsa/csg3uPKI/Zmi
U7EyHqxQ1Dt0JyKz3LE2W+PpBz+JasiKJjKjjG7x4IZEaLbc031M6aFs53aYR8Ta
7WOEW79KIqeeUNtVYA3Y1p1YnFJdJzzL3V/7nCoHv0VPjfgYPwx6KEznzojONn2C
4AbQfN/YW12RQqjfrEzKUGTwOBQXS8v4wHDWV87AAN/AkYXzZKb+oW1ZpAfBxnSb
R8zIMdKhx/Wo6DClcngYm7iw64x+KHSd9Zr41RQXbgJaTCvHCHaycUNAuHNkArwF
tXl0Mrju4jvuewGpay5U5ejMNVgvzxhHWk2/vcMHitoK9CrqhRDniGVk4hyZQIeh
E0Gcgd8GCImRZwzfCzoaryctt72yaAJbcifYGMePdn1paIIO0Lu0dJaGTEnqGNC7
hnbPjHOfNNyTc6P8a+CurWUMohtNek9iwGKYv/4mmn9HwPPn/rzxjAL36tlGN9yJ
L/BkpJ8ShYTshe6SwLxKCFRKS+kIu/+tphhLrDnEnfa9gkbgFcVjnPWVi3nUmtYc
iGt9HqSNY5K2rFeIv10Nptt9JWii1iCyYpDRLrZZNFDOLy6WRlmzSIZX4xiQZAke
NOlgLie1NvhI8wVXthCcO5HOnyjJf7qiy6nx7Q2yIxhksk7RBPPa3LIkDFacDwRI
zNgpV5vnKU2cmFLmtfehBGu7JpcwzO4P0nr5ua45Gmo2K02f2XHRpZ6zuAZI5LE5
GrmWLuA/w7jC4aa2zyLWfUDB+ErG1FOzbWRUd+ZiA8eny4PGot2HUnuJ717Xr8CW
+c9ck8gvvQXD6NaQmGkNMOrUKZtI+x3w8YQUw+UhgYT7fQX+dBMTw6RKJ3767aps
Pl7hQlnx8g5+4RHtxo8wrRiffVMc/nDrjEvth8nQOJco9sXX/zKzHd0YC6j19iz4
wxSMBKtw3PR5W5MLDRV6zMt26zV4WkddhoTWbOdrxsOSQ75FbX6WEPgPPRXODCcO
6oyCQ0sRxDA9LWnsczL7ER+/SmIjVBUxYKsVOR+cHOY6ilFtrO1biF9iKE6qcS4c
YXMt2dokaCIxIwMv4NhIOy+IraKik9kiRxfM1CZguEyGQxKXoh6aNMEsgMC255vQ
9bNwVo7c3WyVIz36YM081zswxFj1mhyY+QCYEON+/vzx9wcHY8oh11pWCZxiqsW6
AUA0KY8mYdVqEvvayupyWSEEpMZU6g/L9VYKL0ZuIgdcdMncxnwTBS/WjW3gyZqF
Li/uAN2Doz3VZxX4+GVgV5LXRDtBxl2zdhE6pY+FRjT9440JI5VIMXHa1FwTMEq2
olXk63B4g9HrLg4vIcRQXGqjsfM+eKAa+5hq+jaffreWTBbIFXYAXaPfqJzZGb1D
RhT+59T2NlGXGcQAEVIhaGmbrycbL4tc9J682nV362V2qNGp4oY/ZHHPrL2zdclj
8Xmmg1F3y3wh4Uoc3c3FCV3TNLrbxrgLeN/zZSG0xQwe0iEe+a3OoUMr1flzXhJg
1UQBRFSu3JWvu2nbRpyR/fKU1GqH4aAVeWKBIecLVxazFnxu/F2yySVJNV+K26yE
jIqBy8bSIk8cSZGmSHy9lLBfa29cIkIoF0qGmd7lj4XwekplWZ4TybLi76G1tsAe
NFepjk6nfmSqoALgW7uR7vD8mW2PdJT/nF6V0MJxKBM6MmnKhR9UGwpumlOJeKrB
ipEYVwNZTEfc+GQn+iAzVCqEBrUekRFsx5GXW0ryYr8dtfoDuNhpcs291KSmWkG0
/3fQzjHQsluaRG/viIqls7XDRK1N4BC6oIQTJlqO4cbVqjt3I1U9mkV4+gjPh72V
Cn7kDa8UKv3IEEbsEiK+HWPp3+8ZXnRxsY/c+bb7YJ9e6oG5xlKMK2chaONCave3
A6Xd9KK8icHPJWJfBE5bv8OAXJNeY0G19UEv+IY7odBaBe+8EMHxzCiP0E0f621O
sGXdWNWv7BGwHMzPkaJSmkIIeZYIKuJqVtWEBujmW3d138H5GrgJ9VgDIpEifg3I
Ds2i2dWRVe3Dseb8Z9VW7eHzJ6FAkopfXJ9jKp0l04ewmlUbZobVAmPFjLdiDMEy
er0uDkLJsHaMeL1OFE+xTtj33YbJZ4ySPYK+4TfeQoNju7DQ6xJJfCPP5NLQH3IK
KQI0Lr/C1p96gKlH3XhY41Y85y2zNbxoyojBU+ZKHCEyWIBlsnU72t0blTuZG9Vl
62knIVucHqsZfZMIT7WvMKE3jlvrQ0pyks0BJ8sFWznSgqYejdTjXmHhe+PZX2gG
uSzeLAZwfmPwXwMbX2MbZzIApt/M6MDirqUkrUQCUljojj2s/DYnjQ9LlCxfbrvl
6zq7TW43QNV9Af613SYSQu3iFX9qbeEJNe/vKJUSMU7jdC6bbJYmDCbPZiv4ax9H
55xDLBLJfNxhQ2eEjf01HBtiOMMbgyOVvo1eL8P2PT53t99e+xHTzQsIzSuEIJNi
5mbV8h36ZZ5VPjknUXZQmEbp+Cyj2w+gIzHDOe464XTiF8O+nH2AomQqqTsiSxfV
KXSqReKBa3vH5VTF+8pdcKs+puDOfMROt4sYW7lsJgvGiqx2urvbjynd0mLIAdVd
pDwrCXjfXTUC468XO6XYq2ZBpZuuirgspV1ltaEoVmT5n5I2q80ywX1L7s/yaFh/
0kxhB+GUcNV/ms1J2F2QRRDdFJGiRuJ3tomMWmO3C9Zdd4VUrP2B+ohfLcKJNSQE
emfZSxCmutYrmf+lPIJNpxGOROT7mJytq/pNx+i2Xr4v0YSj8vX3fWMB4l88RETQ
V2wW2p5MEMBVmwtzvYxVIxdboXoT1MQEAHVYePLc3mK4mS4LCqwru7A4CuLnZzCZ
wJ+PwvSgwsQAhzGvdncPA8mRgsl+ZWT4uKVWJat1KOQXwTBcGu0MPmpaIMUOoUYZ
6ebS8O3rl+lcsc7kbzOq8rbb5DtcZwm/9jgzhaVjM0X3Wz0ZS8lZID6vAVRlYSO1
ZXVEsTNgoRoAUgVDSGlenrR/S9uw7SwBuyceXQTkGaEay1ek8mmR1QHT35WMDkMn
Azn/IqeqxllN6LRBCUNxMEDRv9P76c4bhoAlPyBb+iJgDD8BG9FPz1aBfm9YL6ls
4323IxXF4PB/KtvcWGEnt+vRav10gj82RhplVAQR8Im/UhEQ6vD8AgWyAZmQYM/x
Dk2eoVVgXzSlSz5t3svbQDmowbtQxSi/XDQO/a4uBY4fs/sTnXwN001Qo2H0YhHe
DtQdVChav6SHocobbHKx9ntINawc3IQOhfcLLiagydHmIs4uA/RDwknoDKPMBxX6
74quZW2Pb8Cg7OO47kIsyWpXaVa+k1HSA8kimW6+SqL5DMaKz6utrtkt33Gnwkzo
Ek/zSVHU6nLb4DSzxXiKAollhPqnGBdjK5QDDAtLEsRUa6VZXdVEcabunOiTwcn+
NUBOca3A3Ei90H0mM9m2N6xiTx6K7SF95u28Lct2jWpqRrWt7rJyT8me1OUHdq7W
bRugWJiIrA442IvUEahFKhEQeC2eNOU89xrfOIuX+KlKGjH+256U6L+2bVhvA51+
mPmH8D+aWEsm5wt1VDj/QH3vTwf/gqHocEetMHk0tw2udeq1U/s5mbJLjBmFrbGc
4918eHESSmC8m9NlyCI/GzZ2HlN7LMMnIOU3r0Q56YN9945pJqXW7jOoBHaMvvim
vPR1wCl5gUxOIHY/a3JzhXXgJGe66hQS7DNJO17OU7hXV3UakrdcAdP8KFvHI1lt
uMA4s+wohjApmFiUkyPifEIdMZeWBNCarZ1cC860OA6W5qtl8QKWZvzVG36r7km8
XPLM0Nl8nkxfb5bA7zFFaXEoPXNArnudR/dbJ9LhLJfUFqGaEj/4pToUBl/mgz8z
cKbP1ibcZsuGBHfb8VwhPQ5d6jweVtVrootozX7vXORYvAeMRtiS4sRKLWZHGApw
31pixu2ZJ2Ym6aOZNqsiEuJirA3Z/deGYYNpdnDE2fnmBUjAmVQZ1jli6qQtAX54
/7KaPTUVmztJhQuShYvuep+hZZt5fbYlkk0hlU4MFN7YFUC6J3YLra5mv868lrgg
ETRrnb6wet1JuIim9hEPisADbsNxEjTQDyVEb88QFCBPFy3ivTuwAcxSb6fKm9aw
oWM3HPWI2skmLzIfTwU79ul/uZkferpLaLCy6xT3e+gq/QcZGpQimsWibkkmyzg4
e/vMBtoxETokfOipoPb1DnY0xy28U+E9b2yj7qT0x5lxUGkTspk5A2Wn+00r+FA8
1Op1rOi1x7bURJCz/mn4lpU9hQwimjEjn7W/I/NRqDztFZfp6V1S58HNRhxxeOVc
MjC3OpENHZTK7MOFaAoj7UaH6MBdpWucTHMyNjO/Y6zyC1CIpQOa53o9j7eWXwln
vWDvyUWI9/lUrf31Y9U/MjB5t43EWVoGer/dRgyFWOhESUk0FRm1hWYg8FrzXmbM
AY+nBzXDkoQDi1erILmKS6pMhYN7zC3suHbvkEztr07AkKO5LF3taDwUsC7miJbq
spBEZBYTodpRpU0WoTOvg0yNvnQwDsSEb+hlmmzosmpUBONDFwkmQKiiiwB6d4ff
e4ca6rI43IgvVgs55YMV6WL86LPXcT5b8NmV3jhO/eGfh0JxVt/kZm2BO12iBG5G
hZlaTrKRMohrAsRYpF1PyQq6+TO4bcJsl1LzTVfShQsy71lanr9GVcsUSLzN72Pr
UOPBH40x5pMEJYBZmbtr3cVEYU4FPOaMAz1el3+W4y8asYgdoWv/IVGkc/aM9PCU
dV5fD+JRt6GRWdcfqxFVztulAwE22zIabsMyGc3F8DbiKtmwpcdQIrp4aERkfaWw
irrPHUZ/0LPKqdYsn+tIO40+UJyw/b/M6tUbm1GFclHvjRWDO97A7mj5WxaP2wYi
QFdrOYYF16C1nmNNBJKhYMX+ojXqiankTdPzXHpLBdx3u0q70gASckx9ibFrqKhS
1eKhMhvyGfZgT8f300St0vwSPANIt3lZQS/rZhXRPjKROorOsFOYXWNTVL6nOBnW
wIVhSlYA/gwy1JuelBAm28zBzSZEDaprnjds75DHJBPvbXxjoiR+vf7keYIdOrcB
9mtETG8rdwA7FPFr0eK/HaWuwtcgOquMLLYDF39MrD2e9YhydNd9QDauvwn4nfpZ
C6ldcjEpP0zWiROu76g8moxVmTVmczy4xA2BXUZmw0eS4tKWlT7/TsPth/2o6A65
Eu1VJ6wOdk4ypIZ9On7P/9dPMind/Nx/ZDSJUhiyfUY7iQ9f5HkPbJQdicnm9uS/
FKtr7o3o0/mC/2SRT3lmKIxQcNnjou62rzv96ozTLDVcGOJTVi0SPJKJr/xyuMZA
FLxv+aisjCH05x2yblBHEdbwVlOoxf/0X3eNsktUCTQAiOqMAK6d57ci95q1UYjx
hpErqUIwnEg/xDIq95+wkEo18sUi9vlJB1TIV9Xmy1lqdCqrB4uR6bxDJlGJX9Hq
Z7M/Xihfa5EPngYlqNqS8glse/c7KpmBAdAr/4erUfD/fJf4QwVj5Ze2fI3m9rTv
D4X0N3CHN2ppV4X5FIUmiFwJjON3cMu6QYUFhjRqc9orwCxcnI1SUgTm/Mi6x7/R
5QiumTVQ77lQZWOdy3T1W8zdy2UnU5q9jqJddXG8XmzFOd1Bp/fOMB7j3KRk8COW
1Dc67DOsxmHF4AfiJ54QxO0UOHMs28p1wDdASsHqos4gP5GuUaDpbENuPhfblHHY
cMUUifl9MLxvJKgO1fhfhn0p32xeOsy6s9C1ISRrquuNmo+YstVuLWJmShq0X0e7
3/NCeebppojo7ZfF9XPC9DsQXvmxXb9Gxzmmt1ztpNE1UeauqWOvrjIdgdR96nRB
Qq1dXT5PdYYTCDZelAm48ZV0+7W+WA3WPSpUEwOkGllOCs3WRxsqd5QUxfs1bILF
dodh8V7Mu0MtFpGcHj7IL8swvVOXaOKqUD0ecRgnqhASrZjFMtQ2VoZwQZwkXV/g
JwH8VHcTmiwWMiwjOG3i8WFQg/5739CRaWgkB8qxvQNZiIeGK4JH7SYV0ZYfKI7f
OA6pjNJMeM/KC9ZGdUFtRoG1KG5CWb/Z5CQBLgsBTQUlx9PVv4xF82lmsLzl08xK
hneU6/s5qeZ3u7sDfTDTYBYqDFJgf5IkOIvd/XEjzlRCjNL0KiqQJg7CPOov55i7
j6M2MrAmNwfTDWB1Ws8sG5c9uNafKLKOpKJOKMkBnTLtxpeeE3M7ix9IkAGXblq1
qpDLsQfpzHM1jy1Rt4b7L3hhRVomivGfDhncCZaKyUbXgYsDFyoY8dQjihYcyTDP
WEzuaL2lGKe1jJVoRM00zpwiPDBnvGakqDIRTyPpXX8SE1hpgzMPJZO3EZ9bdnDo
vuE98G4laRSerV8tfukvakmp+m3O1zuo0F6Fyiu8ZQAGTif4sfekoNb+aKTF8968
AIVRnEhwjSp8Q7kiPQtYfzuWlvxtCh/Gy/F0RHVMO1XRMOGo3CA+C1lu77q8qOJ5
+Wb+lH96tH+6/CgCvHbNa7e+xEe48uQcJv/27kGigq4vo5xPyd7tgDp9VDk42471
IS7tiK4VQfA8WF3no8Jd4DkuvFcGGSLgaP2DN5kgMu2mPQ6a+eNzxXMi4NO2QB5J
bj+wY5Wde5iktqsO9VQqGHz590pbTzlkqOON3sgZf7fmz72DT1p+xdmnDDGTurGI
46LC7OVtyR5DqFZ/9IEtrkAoNIMNt4b9uLbcZ7kmvDlWA866HHOybhY9ZM8WII7j
xnIefJ7MgO3bfwfi69llDLJDo+EQUQtxVUkfEqbjeUZpuEpZvQk2P2kL3S87hc6B
YMVgPIzZw7AZVL+xNpQSAVp16+C5SO86dVVao4LL8CPG6ti1ii+udewFFZbH7ltg
+QVDI8YQGEkgR/oVqGtCXEfF+cqPw3Yj8m38dzKuFUW/gYXRfexcT27Mv6cYzyPs
+HR0ZePWVCRoZLeuppmGmhzxXXjou96A97miSufKYIjEQNRyxcH7IrIbSZcFXTjY
Uf+sKWkgu7/hfRrQoeQQtn0Jk420K6EplktbqS/KmM0UfwnRcAuTHTRscVStvHzP
MGztFe6z0Qorqk4b8PxC3QbSjLRlGLJn+4QMfk/jZdQXKnKbf8IK8U5rL3d7l1cJ
z4egAyxjWwN8pxYIAuTNYmIbe7dOgCGskcRYD9OGo+sleKHa08yZ4Sg20bDhKGZr
dvodxT8eWJ4ftRs5xriSH062tkZt1M1DfqDAQePmcyLissHweTML+bQN6sBIAZaQ
eFZTaqp31WggPRyA7Xp2ifspVZBjalj98w0rTAYSIP4YMRnDmVmRg1BCP7DMaFaA
jIaEcQwakhXBxgPqVzXFY4ingGHoAvb3IaEFxBVqDs6BpN93edplA2YQgxkG7XuE
7uAFVhwX0NWGqf/ORZFUiGYb6WQR+r5z9JdJeEIPdA7IRzIEz7nLGyYtSvCdetcD
E8rXiI75BqKtG2Mh4fMs/xg9sxwScnVHBEWSx3lHF7WV1p+LVhsMRjbVc/JUyDdN
U14puhexsRAqm7tRWu86gwOeFGyPYt3pA3dw1KUZHMSCzWOgCqRUsIZF3TjfsTBZ
3bpo/gd2RG3v+PTJqmCw460bMnxDgH+6plgPHcGGIQ1k4cTZn/DeoWyDLtfGioVe
lqJirR7lrGyL//5kjJepD4noS6YO7kiIf//7JEWNti636gLmGMiYZrbkeW3UPIzy
nu5976OnabG0lZLM8y8AgA2ZHZ6VUUG9S8xersY0amIWz/4Maj0NCtksGGgaehIc
gQjmygsA3tmTIjTF0JQegtWnCFL7itAFk0MDDVUn0eXQoNMeIGkLR2u0NatTtkfz
Ee+MtvtnvhbFzWZALbviFqr4Uj+5FkyhLM8M9rYqWPopFvEE1RV4xnHxpFdUfPFM
Ps+rVqAt1hKc6NpxFEmyShiXk8OBdXHf0NMb9QgEA11ARJTh8S+hNhPiMtVYmSak
Dvc44PGcbOn2LdLYHPUZLtUszVoivckyf2H2DZOPPtgPVVrHhLJ1/mxRlLTk7kNL
kZY5+K2KDBmL+WEkW7agVdA5wgal8UmPL6H2qrRBReskTYlDNJD5RWKirtuV1HH2
WQOgnNu/h4awsOvsrFZS47x6cKM2LQhCSJduDWeSsImZhbjSjsChyuQwZN+dwmnr
aYS+AaFQi6g47tSE4cADijSIiOOKG8hfLEI8qp/tGZ++RMphMWUrHm3q2v6aW5MJ
r3GmttZgxIxsQRTtK8sRJ9vFWOIGiWOMknYI65QWebFtec0QaGnxsTIdvlXZvQlU
mcQWtYKBfGtxBZu29OX3VuDwxDY7rrOY1NkCzUjKEZkPfcR9b2KPI4ZgOC3Y0QUM
N/s1OD2nNtmIzVxxactU6A/aK3xJWtlzIKQB+czreyZW/AnOGrU06TG0Qc46LJGl
/3RGSgat9nJVy6hI/FVl3lSC86JmQLfJYVl2UKJdZdsvHVZwBuYWT7RUIS/stXxS
b1M4ebr/jCCrHAqunXzp45J0Eb801n4qX/+O/dKWsDGmDZ8Yclzq0fysFay0lLA6
sT7ImBSAgy5dHzwcEyzrx67037HgfoyCBZyIque1mejbSycl3wfizi5W2gIRFxfP
+eA7p18UE1DTGtLlI10uM3weev9WjCSjmsx8TGYViEx+QY9lN8ehyt0+AOX7IGgS
qsIKXVpGMieouK8P6EdFsMlZ9PKSfa8dzNhyYJ76x7jG8A9KUnvX2gWp17SCt3oE
/Q6/hD7AzFBFnZ6ImN/zombWZ1+/arbkYSluaQdj40SAQyS2Fh5TscF4zi7Gu8S+
1MjUuYKik/0zNTRwBK41EcKNN6yziOw2ScnU3LtCynWrBhACfAp5zG4qen4VyBq9
lPQh2IJZ7elbREukUz0aDyN6wg2+BO0rDuBd9yk/qVHNaDRnxOkKExL/lpqB0wwe
`protect END_PROTECTED
