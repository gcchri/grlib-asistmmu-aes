`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cLjS8nFF9fakt+TpByZCi3chs/+CGsz2+fTQb5o6KmpAAIEg1KuZ0dz2Xya70Kcz
hI7UmaUvDfyy9xJYIqVQeypgpcf7nIwkS1ZL0HfMyeAD2s4EM95/McWMfxvM6YSF
5VX4LYIsNrMRKQ1JzXikNdGzl7M7pinaMfYWkECKqkapKjFB9OMJGHMCtbP1Gn1e
xHtnsEGroKBhuz09W9GTHFSzTEFR8tpD82czGl0CHcu8fvBHLQ4iUZSIzHE0RKTG
tqp1DcKfvEuJPH4F+B8ps+9ym+3QzsK5KUfWCtnf5qpexSnO9lFHY0Ov4EwpVRQ3
LJ1dwCSMYI3NVap9mhNirVMagQr77MpFZm9tnVHjy90yn1XfdhvlVyxmo5Q9kuOz
CcwQ+dC3L65J0MNhk7VY0Q==
`protect END_PROTECTED
