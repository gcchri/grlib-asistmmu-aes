`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1xyxbbxY/i9eCTLIQCMNICV8SONMnDDcHqoVL5VlRe7Jj4v7o/2hLHNH5xKC4u5
OFBawnbPFyE+2S1aqkNr/w0/XjDXP4ugCiVYgZeFqXN6hQBeugUHhdDT8kvIeKe7
uCEMcizNOxnCqQ8T1NTF4vzNCbssesSzpfwR91v9Bl1biwYdizaac6sTVYrr6Uk5
0lkvTIF+4SeBRyr4bofXOvUa0rGhYl7QdzeHlXEE6jf5aPvMR9GOQ3UC94LjGw/d
isgPfBnVRfp5GtSDl4oypyslv5sssxhRhniKrAAtjZqMpIK7WbrbjaxYheh9ScSN
KFI1CKo1DFtMxADzXYt4N8eZaNNtNqRyNQwskqTasXHCnKp0z3BZtcFYle0co+mr
rdMVnD8DeNEFu5RFArXxzqOTA1TvQUHREmEuPEgiYaJhb4Rfj8ZYq3EFyej6Ri44
xCBRQGjg8K8Fv4XXqhRo6bzv0R0M34vpXM/1/6wm4fXbOF5/O+h4J4TGutrB/pnC
`protect END_PROTECTED
