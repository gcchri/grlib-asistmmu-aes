`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uajUaxn+2Vwydknw4dRMDi9Lh1Vdg51P3Vpi2NzSfuCTOPR4CZlfK8PNZXhUPLp4
ZtUF1NwAKoS12rRAnFWrbgYuqLbxeZ8Q1cfd/YzONQR/gXDrUo9PqeXdABExZ5by
XLY273onuZtNFu/BAdrqEGGBUZ2fVY8pwXdcbVdChFsKRYFiefp7+mLpMRZkLlwM
J4EC0CetBpkfdHpFZo3zfpIli/IDb1lFbcfxz6wBo5RA8T3T+rjUeJcBbo75bxwh
BZplS1bgCewP3j6HX93Jfq8aiSfauiVB8uHVPhyo0IvT8ka0l+SRK4kAu6/1lJLd
zL5Yos7OLda/1KumwmJPAwjkQ4drBKMfFbAvu2yiCU8lFgRcUL7i1JfMac2sKMxa
ARgFwa2TVyWrcVi9+xwEf0t+U7TV1s7lJARe7zzKTCenIV4GNgXb+uNx4PUmnen3
+jtIl56vBK8lzk7z3C0mjtoTnUKP3u8tEGNJMaYKC0i32h6O3cJE6Jh+pVvvMcp1
0RcPjGfsYyoPgEQoDBmuv8j5G0K0ICorumOqxUNHqLGKKd56SujNZdEQhPZwleM3
Vj4YZL31HzdXOJDuihFXXKoS6f6eqkZjYZv64U9jWBeOEezFTy1O3Z3N//IeOeUg
oQY1I6jz0iTYrLcT9cGIYXAZg/2zDutedR1Ubt5UM2ucSdmP2Md3Bo2hCZjz04KX
oWfdgI88MWg2zMgwK06zQxWc/0z3+oLexsxLppUcsEY=
`protect END_PROTECTED
