`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiDv7Hy3i4DVnhqU9OkmEaV4n49ee/2EVrOHVEqSF/yIDCwYqCzi79Q082ey0eVN
SVAubmXKOFsGf8wXs6DcbI8XqZoqozDbadnWmTqBAWfcvf3cKbB37VlMuyXuNvUr
CaOBBu/ggc7M0lmZfEl0dzuuIB7QUHbUubRbDmNFj7VCz8YQIjHwEv4GgipsBra0
ha9QIvPP1z1i2shoqvaPHIFH0TBZIkvtayXnp8YpF3rWHjdNWU9dNGYgVXRRus71
GkLFQQdkPHsBKIC+VhfCEOkKAlkG1R6ZvC8GXXLyQAW/Hb0bdDuGaGTCkoUQhsEB
6MS/CDau4VexBssXpqTTpSQ5yoTTYh4OCvoHe/593t1duUrmyZLE3YB8rAdyq6/L
+AJVU3Q0PzkmJyAnQUXbHRbw+hsCc8bzatEV68tt8Cqu5CmRkfXUYsIHQsSem6qN
TOWbG4I7CGFZoOkhf5mOkXei6PIAiDPrQD7o9FbBX0YKuuCxvxL9LEiabKbrN2HG
WH04u6b+P17ZmFHdQVmF4w==
`protect END_PROTECTED
