`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L3JVo2qdal0qO6B4ufrt+ysMVjrjKf5+9TObvercY9BYQNwA41LIXbN8t6WCCisN
77fK+8hOWeydZddGz7Ko6lc6XP6Q9cGTwGgCukvFZqlaFtad4mgJDVD2h8wRnxWq
vpRYbbGGqwshTkJGCP3eEEVhVCsRbAFonJZFrSgT9SqHz0a1MFSTSe3/Flrdfx9O
ZFR5WYkuXWXYT/S+LCjLCRUU1OnPF1Zb/UltFa5c8bAPLKEgzdjFx/ZjXNa+Pe+/
uI0tKzOOiVMF7Z0erWkPTRfs1YxVXUHpDJ6H290+xK6BaYYbLFOXyyBfHyfDrc4C
+ZfYunsV8LvigxyPWMgh7GiLm+CW14Gd1RKJZb7qmPnhbg1nKgEGT83/vKzS+Vsg
rfHqJsy9fZMYhNfT1yw5/O62ckVxPgldYsnbWD7UvZcKQGOQkG0nd08QB5jt0vNH
ETwoPVaURywVd/WChrPTsjlm6OyjE6iU6JUvwi9b6alpx65L/xB4r8uYMw/93ZXJ
pXygZrGPxGda0ZnYcoZpfaJGoxM5NiEgEt+YobvZtibbuXVzMsu43a2yivGTu/hX
8YA1YB6z3CTWarzQJ5wuORAXEKvJ9oooxsPO7bVpTVgdDlddoHX3HEh7z2gltvRl
5/PVAkzWN/PB87TUKvSkCvaSUhlrPqgHb4mkHJt6/oadOqUegEAop3X13qcnYQDA
cROYjuijw1XgKfoNibzT7uEhidM0eNfPH9lvTX2dHGSniZER4/JDVObKM0BzsdTL
mIpXRzfRgZqmiDISZYiebQXzLeMp2bs6QpYj3OOEpgC3A4gKTOuUin84jYKMqy16
ynLU2xwmQiYY2fxDyuGlyVhTQkDJ2hsghgBbjrFufFvC20tH++3LSq6jNQBFa6RZ
r3h/UQFHcxwo12bKOu/FxNQETb4qKGAaxeHBtPDiNc/O/ghLDIUaHuwg0stb/cPM
ADi0Zf70GDRvJldeAkgDSMlMTjOOUK/4bmqp0Hrdo9C1PVyuHSpM5ExOsrkAhJYb
Iy1I1/TZ8m3Ij5TO8F6mwZ1XTV7R3IcfQgEiJK9m/dIaFiQ1vgKh2V7cEsBGfvBY
JbfKUFTeyD5Hd78AFPI97aDv1+pgxk32LCPz5yxCZ9mIj24WmilwFE0Lao8jlKL1
hfLOkgG4MVR4r0n38yonCNorN0mzrrDHfnq7F+PWDFQokUNJBq1b8Z2C5Qc/CPPp
F0OFGRaJRzer8bAjIMPBKLGIvYfgTbFSz0+dT5bqjIyYazaWAlEYsv/54sTlzJBb
hiVMBFqKuQ7EeoyvUpxPWftFC/gqv2+O/aObC06x8rUOfxJbt1cLaHgMgWG48zVB
/yavmcw39wlN6rq9ZB/jRkfi9W3MTstl7r3W7pxES9bkw493mzweem8OUVKjN2OK
wPpKKK1YMhO0IAZe9ClRhXlq8iYyS8uuAp4P8H6Bz4vQUyWseQ40hnU0wplJXJDn
z0U/2xA9PmgOUDQu9ebU/1vbAOrJ4hQPDraEqx6z1wkW66kgeJVBYMSL6WuEBPrq
v+Q8SpISHZ7e9jiqmK1AxVHPy5kr5x0CZyJN7X6UFYYwgrBFfn09WxUxNaOgVbmP
Llx2kUJ6uYa3dJ01Vat4zOm6PY4JF/SdamqIzFRrzQQhhLHkUOreMHdsbAkJpkSI
H7dDgpvVehLEKYKPeJ4002D+5aPQ61FEzaoWMo0Jr/akwx7m9q2C8T0VHymGKgyE
ywKO+i67oolxeWQlL+Fe8UB/Kt+fkw15EdS80/Q7AXs=
`protect END_PROTECTED
