`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mgJH8vQc8N85drlCjGmir3EQxpynPSjjM6n85vAA02Ij5yf+o69l+GT1qzwGjIla
H6nJ1de1u1J4HkBK109HmvITvBb5YxNSTTyY08ObW+8qfpoeaGwjsbRw4oIF2ib3
+0ByKN/Z3mg7abxVY2cYs35SH3thtHf+mGo7IczxHvaKDfAA4jge291KjIy+iYiD
rb448smoC7urO5qSsok5gGHBhpQGNxG5HJ9gpmDLVgwnWMQqDLhtFGtLEvtUHxJU
iEOsSnRtUSTTn9W7cKLB7FZVVfTtQNWZgMgdp9NBQ6T01uemwtfsdoKp/3sVZ2Hh
3uOi61zu6nCnh6wFaYT1r7jmyQKoi+utiLvqh8Dpn4xJRbudL8hdZ0x3zR5Nytf0
Vd16OqRhD0Nlk+9HVY5wWISDH/6EAklLk0XEr6637SbjUpXK8Mg7H1vRffbA35QG
DaU4Koi93iGXAlMACAZ3o+NEu8ja3wAkioTxYR8moTsGWzlYYC0bYRpf2LYWG/pr
b1Ygu69iQ1CfEc0Hic/4peoTnjzHvffW//5cK8wSMTIf4JbwV8UD739FuBiPgaEl
ASeab/UB5nJJbX/ENkMCzkgr+NOzk5JrLYWIxpt4ULd4w4z26+M7GhNZLaSnp8Vx
AYO1pbzOscTgwXffQHt3Xs3onPk4ueRNwhCYvDBF2w1YEcT9hIK75vbAx/l/G+f9
52o3A5SvdAHCxVelpDQgJ6aAMD8SEdJxBBs8QFbOnH1VCNWLxdYNYchRxnLGRIxE
BEMFouiJTRyygfJJM7FJ/XMLMD658HEmyz+7flE8GWZXcgPwFYkyH5a/UXt5YkCG
pRJbL05TyhrNo3/5moMFu4LAKmhgI5eKPeQY1xK9B6KvLfOXrsyOKHBIZ2NrBr1i
xNj8YHiYML6XzzbMvFQml+Hz1F6SOXg0IMBwYOllD2dBe8MAQTf19FXgIZRpWD8O
GJcLdOYUHnhkhpgfdZjvrS/apuQGSc+Y1jGdxeY3taAkJpR1DTtPNZCoLi6ky6Q6
UT16hMqbzMW2FrYhF/9h5wa/SyBgjgBfqJI/T7SFTQWWsF08urTQ+x8Cd/EGWu++
ohmiJ1/8wdZPmI6Me0eIOxtVqYGChsUvL7CCM5BRJSM76SgAZ+dgMis+Cwvqu/eW
JIzxNmT/6aJ1vhRVLk7sDmAZPMChrccEP37k9IxP4UIJD5BnKOWfRqnk+hgolr3P
F/LM675lfQ81wNMZ2dJnY7L3gG/xM+gVrE5SzlcNmNd1G+0sUbNaj/pRwm9y5hR5
KGnhhcY/6sGAJzQjuI2YeWbgAHLs4+oW7Mz3WgdzLkEZsS+Rlm3+WpltlKk2PTbe
MJ5la4EM1oCywpukgh84oRwHzP87hkKKB5uXV872JRmg5jHuhWz12tNb0Gpt+nO1
snuHSorcWcPHd206p7lWRuZvYnXd5bwkRUuiQrMQVYosb4mWfukhkj2HHt0q/xmP
i/GTT99uxFG0uw+X5at/MRSf1GERIUJYZD7BZqBgO4I4LcDYLoSQy/9E9iHjq2iA
Yds1cCKnBdj9kdjG5a19MUWI7rB3B1jjwNE9bUHntOtiry6n59awmNiJB2FXxKaV
V8l7gNlclH+R6nA8jg1HtZK+J6g0UJlbi8VftWDvEJqw4IM3F2MOf6EsmsmMiMkZ
jPaaoyBNgyNDIdndZ13v6eTwzyCQdWRxpk7z+tF1HG8/nHrRBuiiabNfnT7NNup1
508EGrWvZtdQ+mc4kmRKmtBKXvoS07/8fd7W1lf3F7opGSWGLqQife/Znq1Du5oM
wCGpy0D63MMGm2RY1DuLh4I3KBR6FJzBOt5wnnj/SoiGv2SUqMjy63MTJ5/0OQG/
8lqryulOMedz+usKV1zPPelhMPgTiWqsLLbMy/n3rf4IMgNXnInHlxBSbqCqklah
C5ZbZKKo0bsNQUF5vVb12btcg1P9cwVilID8WxJBhIsTKAyQLaS+RncwqlAXD5kv
o3V1Qwq6TcpCWYuRPjZhE4rQxVVx+Ac4e8Yk+GAncJRJOeZdOpxT3ObaGz2acZ6E
wC5FJH/vVO4Xley4yKYy5COqAdDmr4Shqxvcg6z+WmKaNB23W2XDWkZamLFpzqw8
PLG/H0cwhh6x+qPGS1Io58j+whkMCD3+8KVMN/PwU0ZYkzT0zItA3BY9bN6CedT1
7/TF1NVPYLXc3JCV2ih7TMMu0iY7Coi31IHTkDMbWZIPt/lkDnz1NwuCQb39F422
vdid0b2J+YYzG59yYRvHEb+S6lCxZunMKmeaR/afX6z/28Xdj4ZmeiZRiJTe9hBg
ObxHfXeueH5TBq2gHMINZGJEg5PIKw9nctxZPMiKFBDw4sfG5koaHO1pl3xG3VHX
4HM1AQ+VzprKM9jfKlHh8SKxc12KT2Et1h28fepAFNs84RBFPHkocf5EUith7qZE
dfTPMWI2rLBpaD+P3/gh4A7k6TgyqaE1OHl4J6OyH+ZVc1BgM8Y2XjC3/AByFwBb
1U0Zb9MByTtN4J/RR+S69tD5NcVOjZpy2cEqoosQcEKom6Io9htoTgXsvuHloY9I
MfeNMSDC9UuYuVvyqXmtJKb5B5gVqMlidu2cmTIdgZ7JR3wgrwoS8xJr6eYYqt1K
nkaBxVG27Yzjj1tUpgBtFSRDyyPjh4GvdlhX65FPrYwgOugSg8AeZx3oP7+SkmbI
AKd9rXOHClyWFGcUp1XX+bmdq0LEXt/8sIb+a92Yu2pR6xgx0Ne/cCTcdIpQHMUI
gqicEhlon7FfpbZqSSfn3Ny/tbCLcgwBgXr8GQe6QcFJa8rl2bng6y7sbg4ehY9C
/aRTsjUjuTzMUXs/0/R8kUHexLzyOcjOU62hScAkQhrGw/jByxd7yg5pFBE8V66g
dK5jhJISXTtihypy6OchJDjM67yGKlrmK76rPOCFatIfi7IGfIy2l0/7PgPH4uqN
ZE4GjXNEC1j1avf+gUzv22AZ4PQBjR3MpxmGbGa/mlpBMNvEkQr2oApecWQZ36nD
jYLcumYCW2WSnnopO97lv2YQYbO41Z10lZzX5NPYKYiSO6zB7nJFdTLToRF5brxM
Nm+D0Ib/5zuTQVICYYF8jQ92K/AaoybP81Bc1NCcg450n9w3fgEnt5tqJWgo3zqQ
DYMRmDPiMc91vy9YA1SH/eLVShqsl3jO6XEz2mWSg58nQAWIiGPMfVAZxeO9dqQG
/AmoQfk8CCvpoW2xaj08rjaXj9T7+xMqO/HlmH34KhQCqJ1zNk5KOnyWaJ2oVobh
81hiSaZaq5NVPLvPTDCxMbsTb+V1llA6WhR77dV0l7k5Y/A7lEb5uGK6AuO4qAUA
Weye8smaoeEi6FJhesd4oHQTWJjzPSGscFCxwZSWpV80UkvOpYy6bgaQ3ZCqFEeH
zlPmgxQMv4PgGP8NhK5YfLzo6LPUWc+Km7SFQx+uZ2PoUrPuDrcBYaqjx1cOM5iQ
zgN6fRopJqqPX8/ijeq01yccOfdXwTN4+0vR9m2Uqr5VM+3b6P6xIk+qUrvkAElZ
gJfpAH+WApIFKFAk9hM41qKK0Z8p8WXcZo4kCqmN363n/5n4dbLXfh/QfSiL68TN
CxTryTWKd5vvMdoXSLN0rPRUJKwlzAX8/1pxzYZvLtdiE/JBQtM2LipI4EjZXRFa
0kEMLWfg5FIaRzXc4iwbf4/25k2b7phmSs1IdYqsL7G0SyML7tpz3bZKsFrqX3Zn
wNXyi1MlGxUV6SYckFNwUV8OZIEBDO3Waxfi+qKLZFBh09y8c9735xKvHNGGlnKF
hhBnxlvfEp3o0XEw8cphjXMrfLKD3rFc1Ig2kExwXfR7ThyFQmLUZna41v/VIWU5
6J5F//Of4XkqvG9B1a49REBPmanTqxWF9xAoU2Tm0MgMSqzNs8vS63Ah14Wj1iaV
ss4aVvTAL6ls164kpziBbb847bCQ4nuGBRcxolNItgh9GoEaYPiQQVjs/fAMC9r8
xhM/tWED4R7IFxYVCarwpNRaCyWSbIj5qPjSvZ+EauFtUmrO2BFr2z0663c/L5Xl
qMP4Ob8QvIe7+Ep8UjWD8T8H6bKDvwKZh0Sak8gVf7GaQN7o5mi5pwpFMh8QiWlF
mPhzQwadsZlNFSP+NoMkzLbzcThiolqB/KiW6F20JJEpcHbHt1NryMIA5TvE3wu6
kDDHzI1BA8YYm2lFfcoH9lx+4TgiCiRIv1jqG+18MCGKexWMApGXR4xVYHjSpSRW
sn4uH8Tp4g9xMNB/ocZ0px2X/dIh74q1fYciSDHr8Urzr1WDhrm9TJHG+tbbNtOG
hVsxGnH4eUO5eEE6By6+Q8xaz1QA/cksymZWAUtrkXW9wk+qU28Yts+sFrjIB1Zx
BvWkwfHZNNnOGOzJQzF5FFfVT4yVfDQPZPB14fxJidBgUEhyKSaDus+Wo8XUp4YZ
hKbScnZzQvYSse936Gvw2cNVK9JkAuhwUT0vItDT4LJ9CUL9C38uyYEhiRpals9W
0d0SpUkN8Gs05OZsBtbOttPFB5K7uJaSxqNx6/X2+jcNuGsldopEieRsMGKqlwM/
HnPTAnkJozwxdnwDt9SLp39TrSeRIomJZMJumYaXjYH7ITkz1ALVKoPo93UShTSh
AOEP6PkbPd7E7pvxVo/xovmaEvoH9r2FwrPx9VAf7f+m5W7lBHydcLWNAYouJ1Ds
zceqm2dsvNg3RhqcuNXAISRb3ERRyHHZu2/3BhjVeZHfcZz2M9/iYK8BTW+oL+yf
8FnZZGjShyY6bpMzlrGrFyzsXL34SgGUJ/18u69iIewz7+JXAwX7Aa0hXBlQrbiB
noAI5P50h+DcPwuWF3bkr6sGcLDPLQv05Y+pqaMTfBwJQ14brHQqaRYWt1+8ZElR
7eeC41rcOXt57dc6ltCTTGms3Ba1YhzvXn1GowvWvFJ5QmatpEcyVCd2q6k/k9hl
CIfDzLqj2YDpmS1xoK+1OM9skGQuniG5W/SDurh+rAmsqUr/VjVJirU1LOTyl/V5
qMP3gLpCTXm1Pws1NGBZ8fvcNBL4qzZ9enMraOM8fjRu3xgjOxfTN3OQTNN2sORQ
LlBj8Qer7A5K+40y84RHujqrgUO3KP5X3F1VDgzW7WlJ6UyBu4g9FOkA6asED8Sb
4z3mGS8Ekkhkn44ftu4n4ooHpdR0ZStGaTG4Lwc5BAjs2ssxJEgSoeXNwxDgJpoS
Z9bn7Ek2zQtVJNRCqdYH/oKoO7BJ4dkBplwKNPoHV+eipYrUvXaz79xvBvFkNWV4
P/IoKvClEbNfO+5rBn5P8BeTrigPtcFYzDpsOzPY8oKWwIZ5oQAjEPREy0UrT23b
Iy7AWdBI+10uIrXXoEnR5RAYWCwxkyeBT0lSjifSsJSgxzPs9LbSuKkFAyd+Snx1
5NMXnR0x8BLwObdaa+Y+rEgEZA3FPJdBL8/LDdiFM2UE/P9x1DLVMS3veZZTy0VN
77qDSFw0oddmElytxuMKAA72ZIzJQWL6bb46wtFWOgItMuUBV97afXXPtz/sK1ma
jbVXtRPHMjJoaqpg4Sy2/LroUu/0bcnPLskVdGTvw9ilGmi2q3HI1lNPlMUw1/rH
TOAa8twPcbJ/i5QEfAAFr0q73BvrJ+PctGQdYkBQpFRSAMw9Qw4dzIX7fIR7jLf1
jULAzZWgsrx8ik8NdaJZO+FwUJXqkn7effhz9auBiI9Hbt/Dzk0DLeSGsgji+p5j
yTW/FSzgmjWjDyEN/zoiorjZTBVVO7TTeh8tS3S8ikS/rLHwVdHxKMANRGPqBBo/
yjvUEHLMsiR5W6O4pADnMXKfVIKDLi8wD+0fq3zRWMDKCLB8VdNOxEFhLjwD1sOk
AE4DVHs5zA8kHDQqPFakL4eJyGENh6xPpnhYMGRQjeKDnfC2UMp7ppXZtLQQhP3a
FWzupsnuPIEX/kEXnPZjP3/SwXrUBLtt4CqwlZvpzfaekSzLhyE9QacaQL4cGBPM
t7dIBAfFm1CpUzulAzXeLUSQ1Obt4+YVFel3kUkMC/5Fz/d7PM/3y3JpXBFIe2LO
Rp42Ntv37egQMTD4cm9XIWtaZ1Vd5jFMkOokoW256rIld1P9/bsLon4WjYmns0X8
2c86yO82YzFJ5iG41cZfmwWxncZ+FAEj7boNqLPITqgPzqctJ7dAaDjGyrR3jgFY
x7gXluIQbqZbbkUdaprwdAVbAViU5l+l4BTgeItmyigSb0lizbA060j3WnI3rfHS
wYYqhAtsxXCJTqqLZ3wMpQ01yMUNdMmKALDD66+aDlaI4IgxoG+LRIN3fgQD1D3Q
YCY4T0c9sRFMoIbdPWkJefGPS+z+4p/4uO/Ye4LIdkF1+MQjWV3v8KZD75haqmf3
NyMsNvsY8MoDgvWX0M2PvV8NIxyCLKA/+LN2iEWdQpsvaXPtvOLtFxZJ9IkewzhP
1GcJOyMdUGJKOu9eC1CKjWmJp1h5ZDgpHvr8nrpDKbDQrhAHLGTqk7IbBHXHo4a7
v8BZKVYyRkS4hrp6/ze0w0fkMOCMPawjFKj2ILl0yybFXAA5YzglJjxM67CWFPM/
wJUn0DIciaIKFXLYR3umCPoVIq0crgUl/ARG6o4KnqF1nM99porerjqAr6YSSwCN
a0gFNJ9AvwF4lI1lylouPW4pFnXhD1ODdgnSbT3VaMB2fQTVNRTO+pavegg0c+kr
V5XFgaRoon7m/nkzkOlYY9FKEB27xP+40Jc07tVhQ/52ehSS2StNy8wocu0F6eQd
NRRs6dpcLOeas1XEX5aNMcPvyondgiBtnqvVmemYDLa6y82LEPveqMv2UBqXnxl/
8kii579O2fGCMBIsiCinbeYJ8dSscBuDfrZ9QWWIm9/llDgpRFtoA3Rb1G0XuL0n
FEaiCRY1BJTX30FI3Y9c4PYKwP+0lF7z+FSs8L4n9bPNJA4NpieUPCNREsbQM451
BGZTXa6hVjyoNo36wO8ymTpxJmv3AxkBBe1rT710mgcn7N3L4bUyCuaYseUtMPvb
kLe08KCjw/EJgXEGGC2rT5pr7bkTWipnr4EXKu9/haxZmnaAQoijJWc16NiA6I8L
bNEinDRAnxw5MYfbUqUapCivj6eMq4AsVSVzzrozuJ0UfHb8FD02TYzFegE0WjyJ
ik4SCav5KzMaJc7KLVKuN5hFc3RYLfMPWgnHPtcm+WpxjKdlMcvmIdJbzO5A3+nT
UFO2RM7ItKSUkd+YDNthn6NsFUggya8FTypXlBfUTrL3BBZ+nnU6uw7akQNgvCi4
9EDYKrqJ01jR+Ify2VKX2A==
`protect END_PROTECTED
