`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vlOKjZBrVr+i6BqbrHergCb37DVNLXn5B02pY4cCvh7atQcox1yvWRhobjSWZbFO
MGHnqSan68fHaCxHu1pQYsMrgSxpCzcxiqQZYi5fmfir+8BBnheFwR1HHdG4z45B
3G5bLDlJLov75tx0BWc31uBXp1Z7mkC9RR6GaF59lGb66LVrKHeRWlRL+ZPoyO27
VU2qirm/FiwLHKLjKsLBGByzneeXmp23IijP/ZALr6FON3JsJiFnGPy6roWCKJj1
rEt3vVskyE1lRSOxXXUmXS7u1cpZ8c07Wll+qU9hjm7IMKKLh7EpaQ06QXq7vftl
8IrKFgWCvx/qqU7VkohA0mpF+/PNjUAy2t7gVGdkX+g=
`protect END_PROTECTED
