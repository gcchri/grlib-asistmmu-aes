`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cKuEwIPPhLOWTg8E064L80PobZuN4YVP9na5Xxs6pvLLIZmu6mmYGcnAsDGYPEVf
8tt1E7Rufm4tp5IL1RMVWZvwItZJNwyEXEX+9JGCeUb4m4ZKdLky4r9U+y+t5RM8
+cg1lXnz37t1HXYOQPU4ty7KKEGOniu+MZbqn1pOu29e4ptV6SdK88ne4udmCP2j
Cph2I8GWDce3YLn4sLtrO4MzXhxVk1VVpPtJKMMe0R3g5goFqUB8Y1xv261bDqdd
KfLv0SrpCAoXivewRwDEUnmE9CakadvDVRDVD89bnk8HMNuI6raYKVyPSwzowSIP
lBGN/eodSFjnEQYsH4k5fTqtXrHvmkQA6zf0HUJqSt7zQ1SuvhH0BzFsgFlyA0LA
iH4C5EvIgxe0JFgILdYEyYkb0tzr6XJ+osRZm+98gug=
`protect END_PROTECTED
