`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMmxzrKOdBB0zr2Ot17XyZ3eznpRWDfb3bgry2CMGinX4Qsmzw+FYWEGn/6pzXw5
rUzgI+6ue9QZjOVCs1lTmGvDEaFA+cg3jpDfAIpbdFs9sQMdQ7Wb+yEtGPfIoooJ
u/JgIzPZQKK2C/fuewVq5WgS5Rjue6Q70p7X3e1TEe4WTuU0ZwB6vEZry0xYHXVf
kKeCBXjh9xJ3boETfgWU9edJwUmNNwqCvm63a+/lMAP3bYoz4lsqqy0AO2xmek3l
Y3IcwVduNuRHR2Hqxst7dSDhhjzJYjO/H7t9DPGJGxs=
`protect END_PROTECTED
