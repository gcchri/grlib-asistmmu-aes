`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHJ7gtMq+FAp/xeDhhF5JOnr2ixLbQzSmovZHXL3tprYF/jGjW+bYaKbkZaDCjWk
IDsoktEHapPlRQeAwgPHSiKUr1E9nYBr1yAfmAKEpBilT9gT+1m/EefsPNwV08as
TYaYo0RLUgBUh0ZSQNJhN0JB49Edp83EXEygzisUUGVbu/mQ7LCZJutP1DskRqcY
q03+56kMV82Gxn1KQPQKGYZJCQh8zy+wL7pO1kKywvtiUnLW1JDqJdDz9dbjyYHM
R8n84yDJk3cWb16wMOulBHXZ9qK1DUfRg6e7vn73dVoPSYBa3d1KG7SrdgGWDLh0
oup7N1tPsbZk1aEogppJ3LN7alpUM+QjbUU5KpOW5f7Ss+T8evPaWp1zXL/jsL9t
j+bAF2sr1ZHhxNFP18PeHfJ3R5zlvfFMFdnmvvtNRaihl5+dqAClIun2tN0WpPX2
iEHW2hVlD3sRtgQis3vC6Z64/OYeWmGZ3kmAusK0THHTBl6EFZUetz1HwW2UuvEK
j2Lm+4ySV/tt6voQ2Dkz0uozEZdz59u9i8QFeg09XZYL7RVy/PWtRWoLqArsLzHi
pMAh3bkhf0qMc6F8bqbXChwGCR+AoPsyeQwkEtR336Fw2Bkrgt0wV9hVVbU7AoeY
YA87wf3G4vxrIPgYa4XeX05Hq3uOU4DiLO/PzTf4fK4ulOx3s1ztfnQ4HFdzePoP
qY00gzlw35MR4y5RiBih/ewN8Q5HZtSpwU4TpfoaMBE=
`protect END_PROTECTED
