`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhUbl+mIXoUODC57Or/K4Tuop9E9RtgyoOU6IZlI9oYnciyj93BFJqUYTtF9GoDf
2Pj2H6ivGmUa8cwgwSdaE1p/wkVaKzOnpkfZHJE60A0H6ChGkyC2ZTKg/NYkElKJ
mrg4BiHiJ3055ZAeRKqFSywFZdnLIpFNt+r3WJYk57e0Cy9j15hsRoL23ZSxx9LJ
GitAWxWIONQrGn84PApYwpTli7Nqt0FBMb4vcXXqdjyzUP9Uk4yMtp/SRd7p+N6A
`protect END_PROTECTED
