`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y9R3wNvfPs5GQ8jPbmZq1X58IvrOCIWB/SUxspACSNUOOcps5VHcZXI/i2mRm1Xv
18PIApNZpcrlz7enjtbdRX6OmTVUInD2mdH3CcMQcUtoMlVvHWInO/CDy5Os88EY
NGht/l8AngfzMAtGb7EjHhNb2gEHDez+aDAHcwAuDYVKtTptGqXam+Vw3JeTMPiw
jhsOEUSwKivrb9GnKZWi4Adc1AnyZr2SAMe7eGLr54veMDlSqhzmffTNrRO+Vbmi
5c7N+TRPebvi55tJTXjvUcaOHOyHBtk5Wr1x0WcIrRN+KYrTvM4S7PrZ6SFNRbdY
0Xw7ru0ZaOx9eq2Xip5PswNnxVPhV7p0OyjuaKe/FnchLrOBfymN4Ck9NtwLJBR8
05jQe8AurT6NRUeNarfpn/xMeUVZzJnTi2EJnzYmso6Pe86PqNB05ModW5DzI5fa
VHgXrQR9egyXVpYN85z1z9vIcBNkkKz76DpjUxrC2u//vFwlfsf/sCirq6ma4AWz
jAYKiboxg+PeQqHtfjn6wHbXJzmgWfVqnrcZDP61ZpCAY0R6aVP6ZTSHREeADfUr
X9JcpbMLAzG/K/kkbgsCtvr51IhreRPLkUBZci6I9ChmIfLZCm7rXaqFUSiFuXpF
C2qhU1OSZdE/GaZfaVeWGKEIK7gEOhRkl1D2OuOBL+Qnm6M1pT2W1AwiWIxIDtE3
Qlh3lH2R3/TF/THtcV7MQyx8GU8hXggNST3PNnTn1aBz+gH4pKLRThEylTXAwYIK
4IhfI695whNwotzKluBGROE3t7kFtI9ERRFGX1PRtEkTd+bvwE/yRG80tfr4MJa8
6yRtjmZeAUBVCo9tUOUJ0Y2jSa9cBpitPlPqpHaghJg6hXjaqzE3jXmiWreZTfWd
Hzs4wWHr4vI/021uaqjPITsBfsrJ9yldivl9Z68Cc7bI/gzr0PMr4397QhBMzGjk
2ND7AXKwDRCeXoyNeDn7AnrOFvZxfWFnGXM0bDQilIZENx6i4je0jY6RYFplTaAD
QYc1bQ/Y/oeObiIFZSBqdqthpYcpdgVLN8Eu+JAn1JoMOYE68/LNOB4+FpYIWMEn
yKrXPWq+vJNI0OjMBoB0rpVYg1J4l6RrIxm49XJ0w7qCk400+rogbVSBR+2QethA
Mhq1NLNXNzmDSOCiZQlLYlYf0BHEHbhDwvGEI36Q9OXntFIaOVIzcBjIapVME+0F
1ZWAEHk/sSN4fBgPm8C8TD66LlnRhBkZgJ6tuTqZ55S1P+uHgxarxq/Jg42eJfJX
rqQkIT891ymLw3P/7el60qpt6tnv8AAUqdXxybnhRQfkVoXUXadFcInWBK0W39jp
F/rstK2rW2WQ0fOq8tz4jeIKF6VuB8zK+/BJ3ijct83gdBULdZEMSu3DE6TmmWPI
y96cMIsIHQgSHTB8ldpb6ulVkmIEkVDMGOytEdlBguMXpm3Hz5Ul7KZTaTR1+9+b
7LivXd7zawnZHyKzXzOraoOqBTzYB4DnVAse0dpw9Qc=
`protect END_PROTECTED
