`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/hXMfruJ4b1d1ZxVC4G/d8mlReSQrUHc804fV9GrG0yCo4ZlWv7y3W8IzV5lzfS
HmFLqR3i9YnmJbXeCsYQLx7Njwh1mOp2DBv3NkmsmlxQn8rvwb+y/JDpAJRtpCXO
PDR0AfYXa2msKf58vAypHQ6vWcxz0DUMqzR0D+JncPUzcC5HLbhCUjzczxEnMjOR
12I8tTEl6Hvxk2oI3tiDXZ6NA3FTxOXLPrRBHbAi9x9LlaMmPUlONl+g0pBqu0He
lPXp/nETCHiJCm2PjbHnConBta4kYPko0avbFpFoStTQHq5URrJArv1If1+crk/G
mm/exogrNhHobeEngN6kP/cPemu8FQwsnT/THeWzPcCy4ESeRDDaY1wq+3wZ9Amq
wRjbB6uH3N2hjxUY/xMvLQ==
`protect END_PROTECTED
