`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10hIChsoKtj2GH7cYP3uImU23G7yo8Rr5SWdFRwzcBAczi2U3CdGnaVGtkepigk2
kG6GN/3ALhfjRjpjiBo1ZMkWXxMx2oWBS7+lvaYQHA63wzFCuZLhdJ3PncmwoCOi
Mj3vbSgaREZAMc1nG6VesNyd6TD3FPqFBKghNEd3YNrKD3DAs1sW2tRkVX6oyXGn
ZTuT51SoHxwwjL1mSt7xg1tSZ3O2I8NpDO9e+QGut92H3dMATj/MZblYkHmnqeFl
KCt9wHP+mo15Z9l+pROqkl7XL7295yjTO4WBmjzbmcPQ0MZlALuIMMRLQpcFphxq
rL2QJYf+O7EhiSCasWgKusD0+p5sw37tIaVzStn+Hengej6eKk+4I7hlYOSu8MXn
lkPfAlYk8MJxb+u1TIVFFVbc0mpNqxQLig8Jn2v42GA=
`protect END_PROTECTED
