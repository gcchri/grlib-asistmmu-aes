`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y9Lyixpvv03k12zmzxzB4VXB1AuyLl0iNR751bUZn/sLDRgMqUMkiKvzCiYQRlIJ
pJIYDHST16ylIgwdImMhFl76YCxwnKpl1/AYUqsqsQiwJNzo7hDULJ5FK7+pCvOK
Hyq10pcPFsgUUAy51a2agP0fprSHY5toRUm47+bjgkjxyHDava+pzJF2LsEn5tCF
evvaKeCFXwjNF3/2u+j5p+Xyp+Hbd0cAbCzYN0MvIZixf6xpSesDmlYgcdtkGrOB
G3sasREZKRRpOFDJXzBrLQ/8xNE/KIeOV3oHz0FepNqwTNKOLLl5Bj+BbX3Bk+sF
7xBVEKZTolovLNQkeyqwJgMuJ2cMopd56RSePKoY9GeQzYLLrWNJy76aMpYPAfZ3
h4NRhwDrdRlupOZB8hq20BgF9F7b1EyRrGlIi9pzt0S0jjDIIOYKs7ewbxqPedn9
Hy0ppVdvMSqaXksxOM/ytUYgsKeYs3d1CLj1bdXIp3E=
`protect END_PROTECTED
