`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fe6VaZKF3nemIYYDjNRTDpbgHiYcXjChDyTkjr3lnIOUqDeCmKMFWoZE7T1W7lx8
EDga7YC93lVF+c29aOSFkqxcb1heQKF0N0JE1jjjkM+FWKcmzsQlwGeWsWG3ZsV8
TrOiV0lHjNQxmIgMzj5ZXtWOZe1ugh7sJrxDSwj+pXoi71ZLXmndPucvCfvhBA4H
/WcWa4BUvgeNj28San5zo4ls6D4h5HcDTCB8Ful4uzv8t44HnombijSl6DdQKzA9
ChCgXeJBkPAwbQaB/OzlrrHxF7bqS6+eiSr4EE/tNXoBK1VJq7wWihDfmOMtvrk4
USERFbvFQwmS1Aa7gZ5qeXfprPDd2zCMkKhdSAUwci+pPGVgff1leYe5MD4ApEap
XDoWlr1/Ly4FnpQB1MmQWaWwsgLrk+h52S+hRlx8cNbN/Dx/07phjjnVjyujwN02
`protect END_PROTECTED
