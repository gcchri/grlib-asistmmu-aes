`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDsJSdlH7eJkpjha97h2t+XdkkdfYNGIRe3zABXKwFK+rkzuEzJDSqM2jCu6n38D
gJL2yxYAlV/cZvG8foJa4IpmZANDLsa8JMbh5jI0PMh4kKmNTQUrda9z6JVuT4Uw
uxIHjOECD7sHqyi+b/PQ/M8TtDE4oerNmEe+LVvefZHznQaMZIGBEMvqEmuxDLuK
LudHFiKe0a6ctCf+PTdOo9p68aDeMH2MLPhVh1bUgbWzddWdFlDo7nRep+jndkh1
KR+tfEZW8ny1hYp6MRFWg31ulkrbliAXvbQgKao1hNvZAl9+HC8W+Iicy4uuiv64
exZ0E6HDAPSD/x45dOeiS92g+ZnCoBMIYiPSe08iLOE=
`protect END_PROTECTED
