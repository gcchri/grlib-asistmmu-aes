`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YdDa1LRIKhWkWeRZgrGW659ng+2yei7/wF8OHCNI+xNrQVn2cv1NUZbZr4qyXK9y
mi5iuoPqSdS4joGh5bwfWLnqcdSD9165CU6ElkxCVe1qF93GhTFbAyr7maDS0lNH
uDlyg0esP3+7GnsWWvPQApgFBrQrqTD9/vXvQqeLtcmxEnmSVgDnM6e1qs9OcP0N
kzv3XCyCaf0jIJFULw+ybc5UFV40CI45V7aK1lInU2ujRLBaEHFdHyuJexrZ60ie
+Db7Z0YPPF++8ZZlyApvCIe00DDoS5Muegip/YlTaaw=
`protect END_PROTECTED
