`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pinLdQa6TA7hC3VP4oP5OASCyhAHb8koq/1moMd3bXA7aFPhQwYqXQ/q7PE5KB68
EzXKCglRYG3AaYEWQUESPMPhumUDTw04mIY03j0t3f9CNf7POvT9ykW6HlXpVjkw
fp4AMHMjm7dYEQS+GnHlFGaJD5MAPWqE+ue43LXwGprpHJ9Qx2GWUcdBaaCTmJ/k
yjtK6xHdLVwcLaW3pjZWM946i+A3GWmDew4STiNqOX7+Ro+G2WIDvvxFBldQv3b5
K6jM3aNNUGU4tezHhVoN1EKzerxXgw19ZxafOi8bJ8qybdhKGRBro1OpG2LLOmra
LXFikK1dAT00Ovw7w776pAHDSyR6Tkj+WrionKAI0O09J/gqYRK2e8vS112kwz2s
S7dnfRPDtkKNLieWRhXjAExafKCU3gpqWie7fl6Mx7XB/axuAxRO2o+Jxaol58wR
JLA8vwYwFa3NyFfZs4BppyJF+qIOT45kXRvgdZNGZso=
`protect END_PROTECTED
