`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MH5VDBbo5/ORXLoUDgbSnN9Y3UlcmGxQykLeG6vg8H4t/l2Ja8NfZAxPAMSu941o
Fq81I66HwK/kwwkwsYVjSm1OkottFwg0Lg+MFjwWV1ulkHZVdgdoplTS8Ya+ZaKS
6Dw8u8izUmEgghLPKnDnjqXLReBNK9AI7g+yPoG5duUPa0A/eztgRtq17bwP9liN
5WXT1fdk0nmN/QliS2uIojutsvqSAS+l8LqQvfPfTufG/Mue+H/QksLq8njRMDov
nZfI+ReyejSq+PTYf0/WREtd1ZUweBCNnRKaGYmJbJlcjM1l/hn5pKCwySlo93t1
Sg/JYrVCq1NfHvll9xxhu4LW3ASJ8Oo9fk7iL12WnwHJKjKIb7IjM6rbyeUaZ/Zo
KE4ivuUgZpkLwVBZ7YX1vuzLDQ1iOCrB2U2DutcJVUM=
`protect END_PROTECTED
