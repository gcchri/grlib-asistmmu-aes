`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OChjF8XyJeKjpjOe2wRTIE+n3X7aFx3dWyyJ345+2nmVxMLOHb+Y0mWA0FkpVMP5
UA4Z0709Sfk+lqKIYhILnsTqRJuP+SDVh8rMBEOE38imbL6/aRuFX9OXfZgq3gHW
m89iwpiP1GwqoOLTIBDUg0YiLWYFDd2ZiDiJDgpBdontUMOhgoPeGCRwvJWzIV5Y
IVj70EA8GDhK4eB91pVu8M3mlqEXbQB3Szr6Fxu9wZiuj91k+9fw4gz9C5PXIMGk
oIb1fV8TtOYTlVnj6ssQSK/AbozqKOtDlGFKf+89BdZ5k5E//sL80zaKPcDhJzbN
T3MpZP6dsNVWOYFlqgafVQ==
`protect END_PROTECTED
