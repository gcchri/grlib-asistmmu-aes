`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSuttQS/WGOGp4UQn540FBcUWD+DFPh9zh1kMxtoAGsEL32vfquzkUYYh8rqHPGN
F7F7jRCnd9lzURE7aWmwA1oo22cBvNWRTIYRCx+OjPQxGovC4XSeZSW9agmGODjB
NKXa8CLhpYg3GGdre9n6huNIKi5olkLyA+gpQs0nbutDE7beqDv44I+/jSI1mbZg
uKZ9ziDN4VmlMc7e55AT4sy8Sh1XLB1j/NmldNT+USqRBpr6DAZFtFZ8qVNZH7Fy
iq45cOcdzDqSXUJyfQLquU6CcN6VdZfXdv9Up0sgbu9S2u912YVu6fj4r9fKpLwM
3QJh5w1C56h6OSlRjv0AKviz0jCYa3vB43cR+iTzlR2tMBmXlBThWo4Gk+b4l0Hy
+ZxlOkBcKD7Uc31w+fRpafi/5yN5tEHWV8frRdeO/7n/enWrxgvnxGlys/Paweyt
S3saMJV9r6E0E2enBJEWmg==
`protect END_PROTECTED
