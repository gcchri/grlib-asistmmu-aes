`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EfLqTbhVC0jGA5Nn6aip8Oglkp31lBYS3y0U+9ZtqygTlHAmLe5K39difr+ZRZvJ
pGigjqZBBa/a95TUfywVWgCAsE06axaUa0xqW6auUvJXuTU/V4OKACgGUQkkUxHb
B60rsvrEh66/OesaeFblL5ZxYwWUJ7FD4HcIuHAHXKOJg/edrFrW+hpTef9V8APl
lYmEKxqW+0z+/W69Bh+iCD04PDvdD3KfOGymih4SXNzw6KBDfLq8jY9IRl+TAwsH
JzHvvREl0HGkv2HfKs5t1AKrP3AEM6HYo63PhhRiknd64GsObEd0Dgq4vruMwL7x
3Y3ncA3t8VmUcZFSTrVPJBQ4Qx7iHyE40W2LLPmVCjl6oG1xKzOE7wo8b45lN3Hm
GRtB784vkMOgooswJtWQq4fEJOMarl8eaatpNCK2WhGzKEXmI8VXS1KIa9x5RKbA
6UdTUBxX+aPdaMGAbjkbRa3gj2rOEcjcYYPmOy9lHZ/xw+h+vaBIfcHCvv+HvhzW
PTY2dcRAJf4irtto4ptgaanHBnTT2XrcFohfrOSlNWY/HFrbMQwV25xvjVcN5UAL
0X6vmXRw5tp73PwWcXnFhT3K0dlMrQ/weEfVPn4pr8MC7L3X8LH4elXpdu9rondj
md+WSXcFD8m0ma0nu1JcP9WV333EEbPkuG77cjlDj3CaP9bTHNV1wxKYOjetjM91
MEwX67tDjaMW2MoLP/b9neKwfD/3FVfhNSQS8rbPvyZrhuUVEGq8mQVapsEogOSf
Jfhc1JDA7e6W3QLOGrlFTDPkyDl9lw5VWCFIfZ6x0CWafIMSRBWFbVEhxmESW+oj
11duIzwtiR/IwFURslEZDfwYgzba7vJzDqFRRRGJs/xO7tyuCqW8wGB+iqbhhIDv
Kf8guxxXTzsKYOrmKlcdUJTbAq68WFPbjrd4ogP6lkZTld40q87MdQemrvmw0tDF
LbEjreF2D+7Tiv0kzU5VsDfhsVJMYVFdX+cXw7WY/WxHk7bv7sEUQuKnJHslRZNS
gQJK4wYQ1BjfxLiqyecJng1aH3Om7Aje2ohqAkT4RiMBD+dcjGxjjwhnPxFx+7tY
mw0JHBijmZl8cqTENGmNop51ZT23En7msjr9XacV5cxb/O4ZtOceTASnbI3FngFw
RAXk4Ckb6NqKUOgJIxtbXA==
`protect END_PROTECTED
