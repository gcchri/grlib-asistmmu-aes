`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ik0eq6z5j111zjX9sPxWWjtGPdvP8HM8YRWEagRg0Uw3JZoEOMtPnmmzwR4ihcG2
LN9/gppS9mb6GWLFWhTIsgj8mIGiHEgxlI81Y4Onna4WeTMe9h1tdXPbO3KQw/Zf
3yhpoC0A/CoUJynQ+0UGta8tfMrc8l9nMS/1ZdJ0voTK760QlXveyoglbeCswfHn
pD+NL2N2uQEUr1IdDMdGbqNaqeZjkkAAg2F6xfd7l6cAhvMKSJij1D8Uxu9n8bAw
2zqElJNcYd9rSVwaXvZFpTwpzKkrnRaKbDGJOb9gzereBK4hucdcHGXCvzXXtME4
hyL0BUiPh6t3nBgu3s9Xi93G6YM4CxjUIbwZrFo4qONIscxtJ4sLnbi36WedgKhG
T3MNMfVO4VaeL/TZbNpPzUjuOf+MUvc1vP50YW2KBhoYo/Iu283TGuxDKuqxMT2Z
4WGnP+m4sjZvFSsvi36aQcfNok4fltkuXnqfhhBsVZ2S1YA174frISLOQoKRHCbK
O15LJyhA8+SZHU0eNsEYBSYJEAadJ1j2UHdPGBhVUNKp3fRf/M9GiWhbNQrsxWBT
398DyB0nwbcUjczPza9VzDVqr1zcC0YmP5ZvHdwGDE8=
`protect END_PROTECTED
