`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
es7OBa8AuyuFPT8ZGWdKmK3lEt6Qhn7j7ooRMDOAZiXbIK9T+AABqmjvp1ps9V2K
fz56GEkEE5tMgoW+K3Q0b3hefSNiRKqL2znBhQZa/QkH6FPOZbm0P4cO6GdPDKNz
zvhMY2/w4d+mdLqOhslFz/h0HoW7NijhqKNDPr6AOV6VMPUkHvl3754Qpx3tw9Ea
9CrdqqR+WPtwq21HuXHYXfFrtQOL3FcOfSW3L0ZpDWLvBu6S95atu8to3Ml3Pr5f
/EbUK/PxBSg9c/oporHqYg7Su6rGn1z7erzZWGYlBJUZoJ8OM5qclJHXeL3zF0mG
Lvk1ZwUxe2K0qeMN7tlDEDXDU1BWd3hYpDTiIxbCXuH10CgABs+sTsBGNefWuQXi
X14cp1OdH3If0mGZxrK4NpyTZ1XKzzXn/Gs/GJKntdpbUF8djOgqvxYLPYDWZ0C6
vclAxUmOmI7LYVbp2A9zX9zi3PiZXRLqXZbiBALcPQQR/BZbKy4JUBYS/llN/dJj
wOfpbxbREZQmwlJ0kwmd3jPuSkh2td/A9D7z+unBaNVbLzeWfawQgK9jN8qqVVLs
4iyNFwmLZqVQhI8YJJZRu7Fmub2gdZB8kKZ7VFWV4YM=
`protect END_PROTECTED
