`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AI6IfAX4IwlutwU4DhyOm3RJxBv8VE/Do5npqxpkT2dZ8lJ5L+BVjUng7uhsc5Xe
5LKWB/u7XZSfTkDVeISDqdmykk/WZI0QJExC5qrZggxYB1JKyZa9OPiRmrZ5FMmQ
nnaKuVarZ0JOxvpqYM6eEDQ8reqauiWUNWVKp7HLWEpQFxj/IV9UsXxFdvCJfK2p
Bvel/rF3o4tu1GcpKJhyFeULahkASOxdBMeE0AEeIcK+R+UqauUoM72OXCgNbj4x
KO0kd+1WpYfumH1efbNyw4sAjMrP3waug6mjozs6tnkk8mrJf6EINTGCLGb5AUvz
ybMgMnBgm85m/wb+rl8iTRrYCQGx6xkJOR5vyh5JWKDuz4yzx2rzUXGmtw3DWC8T
ENnmPp4pYJSjR2/ADS8qs8IC1UtvTqRIy9Wmiz2Bg3RluOcHGe/hUpCWSmRBHK24
8D1uohghoL+Kmgs+4u0pqIxve41VroxHN2/cOGvb6F8b7rrsrI7Rwpmv+bg6QgWA
ZFqeCZPLk4ChAPiE8rj3Wv8BxuL8Ld/5zKlV9lcG9Q/s60JwN1ouiEjmAFTL9Ao+
`protect END_PROTECTED
