`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UfvuocD459iaZCsfyGlL1npkkyKBozUxduDdSSFxFnssw6VC0HZMuw7/4lZufYuk
myWCOR4IwiyJcjFQZ3wCmqGUfVkV3S/hsSfmTrov+FJAug/IQaxcwJf2fxVD1Ggx
sVYPg3T/i2hilbmB3c2j3f5mHYbZOpKBzQljeHR3tLEniw5S8lmO0gVkKsqrUITp
fFHkJPf3kKC7wjlY0UiMEOkm92JWOcy6KkiYR8QtzaU+/E6e9f2FdJNLIOjXqXAu
1CZkienl4IbJXF8sXOPHZdliSKZRoDv4KGTNeBp6ZHePn1yUsjpZdfnOJPHWiq70
VR8y8WuhKLQDn5YjcyEOihfaMUBM5KVYp/wDcidk3fp73X/AHMvJxDSrYHQrcnzp
NSPOQO/fuB9IBoEqcAVbEUkf/wPhZ0dmB2E1ChlnuqY4Tj51nzlLOU1u4ooR65O2
QnF5AS5W+wjokAKJVTV19IZd3JJFJws91UG6KACr1K33edvq8aA47M736qNlzfwS
PxvhDclrFF4Nom+vRn2W368XseSxK3nnuglDQ+f2IjXjCamgKebQRLsjB5WXE8MR
Sxh+7hlE0840Uwi+xa3CXlkH2LYiEEKjFmrGuQa2hRsH93mXn+LW+GY8QmS88YaD
6UDAx0HlVnhEmaXn7R90c5jsI/3LoRfpAsah++p0vY0=
`protect END_PROTECTED
