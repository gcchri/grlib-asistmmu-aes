`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z+ROzT07uOGs/eK8tZ9ApYTWxDQCX/dFOJHkjjkXQi0TnQVzpuIxoulGOtMazBPE
j0QX6FQt4JblZQ8sRb6L+KU0IaivZj16L6vzhxYDMRUIKZfQJZ7dIMuQ/l6LRBjK
ArlfdWqFWZUV6miVgZJp7Vo6JYuaupBEYadrakppeld/Of2JZ+rIuQRnNVccuaS2
6ljXWLNBLOWCFb7wymE1EaaXHlV+PgbZltMqoRJAPxcfr5iNY+Smmg096Qyjqdjq
N/414WYWuQN/tlfMdINEeGFK870SrVhq+ru6K9mkT0f9pGoqzA51i/VeblzcOFMd
3VVK4KO/p5G1WM6EQJbLPCQ58N/IjWOQO4oz16pjOq+96048EBQvQiCdBxrLbKPn
tUbt+vpWG4FkVNFIUj2ymeISg/dfDUvAk2E7jPLI2JYEj4Xb4kFm1iogD8+eLSVh
1e9zvgUih9tUP2VT9WMt5RmjoWfqnMw6x2MCNuDoLFAqJ9sjIFSXNBzKYD4Orp/p
`protect END_PROTECTED
