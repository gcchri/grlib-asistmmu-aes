`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYhz5Sl7JvdcVdgb/4yLdba2mScDR1IIF6I+D2md1395872/4s130fQ/blnaQ+mU
HO7YyQSOfpXTYsod3kZfSH5Tlusfs11hSYLaN49+zte6SqhYJZ1FmaFIT/AU61UB
+3HKGQW3YPipL9fh22BOG7IYEAIihsw4nBNIt+KayTbotBcIHPCAueewnsEtn4sm
zsoCmxkQDB84YZgFkKEGv4BrXFKeL3qcHpHB5st0wWziuXmwSSrh8KCq0sYuz+Y9
xrLjRgAyqt29KgKUVJ55LUYzQCZZVSy26i0pjJIYOhfp2lZLnjd5OJbUYS0boYmA
J0QknNQVzhTVqt5a5cNdT2Dlsuzxz0jT8i6HLL8oW/bD7ufXvJYkHQQT9i1phtTo
C9IAQIm5T8Coj7yGe0SlIuIL16ridwFYmtZtENHbapiFykj+j2KO3xQyLMQH2BMW
n97wfhTMoYWv8lDVEmKV6wCOmqJL8YFmunNiU84yreotYAyz+qsC87vSSR65oQqW
7vLBPxLGke+xSjAkOeGkeGJ5us2tNkbEI+dQJtVDkHBdMcSgOMA5WjTH7S+znnMJ
fPlyHl9Yi88zD/n1h/cZRBmNADv7bUqNrBnXeWBdqqc=
`protect END_PROTECTED
