`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yJUzOaw7eZPbbDZ11y1yPJn5zJ0AbazDxoltpvPSZmwUqkA4LiPb5cA1+fFVveF
vpmHLZKf0zDSXN5FiByyag6T57nA7j4M31H6+cuN4EgFvommrruIQO/I6GNMoVen
LE9hYaVBKxInXiJRAiV561ZSxneyN0Lyg6InHI09KVMLjQ/1TCMeTcmKTCklyML0
OVFEsXiY9liUh62oGIKDoTjNrlRitqtQhrQbMw5ci8Lusqxv04tcBuXjEJUkPrBU
jy2QpSe9FXQ+Eq2JCjMmboQ8AT54pnDPx+cjshmb3GApGSOnmI2u6hSH5bfl00qG
GWMa0QMGJYPSSFDHz84du5K9iQaarG4hfVkfw//eKpw8nPIFV/Ds1aCHIXOBpHCO
d3IpgDJrmEYaFnIOOCxdcClC68yAdANLq17EmqC4jQNW2D5aHxylD2R0ZdzR20cJ
YNssRjK40M7x9WSu90ofzcqIZKSEKEKmv90UTSzp8/H+LHFJgvAVcooqFL4LLyVZ
kRaHlqhTGWMkdsQdLhgtl2IHwHnuClTIwegapdldOfwE5JH86pfn5loF1eDamtZL
Sum7qexLq0yEgRfBrA1XIi5VYrYmlsf/x2++jBA/P2YR1fYIm4Ynek3HrNMGHRQU
vsyNeo6Thn33utfTATo5iHJrri3eBc9xa9dVUQT594Nyuksuo/1ECQ3uUdsb5H2D
w/NLzUUd02byl/63YYqFHUaFfflepuyamOirjcq0MpM6OK7QqdAenLEXucxMNWh7
jfxeu73d8f2eupVuYrYGhQ==
`protect END_PROTECTED
