`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gd6xOY+4Bb8BklYjccRLjsNqJZi0GxcQJ+lJQqf0r1SyiL5SAJLx1LDZcd2HNqvS
5vCUeKu3VFySR2d/zJCJxIeLVmRYNO60/FcQwIPDKo3IP5OCMbO1yYqulzUhGsZ/
GGK9OJvzxCop0sn22ch6p8IFFc6s3SeE2RgAEwKZ48GXGzBqhCC4cG4Lu8KbzWaW
4CdcfXhPslvS9nrrFRwB9QL/ZFIOqLuA+Dk3lfTwPmI/vtd+w5zIcr6BBQPrBYef
DVK/L13inMCX2UJeKE4W56C5JzKzm2Wy/JSK1Vkv7VCEYv3V6IehhtuSDd2zizpq
8UNOv/p8gwYdpnU37SYDoWW7W1+ddu7kFPRhCK0i14F/JfJzPKcdp6UwezcPT/Pv
6a6dpV8J6P7cyaukdNxRrbLUgOuJl7ompG5XfxIakY2VNAc48Hh493atDzcMi0N8
E7Pu06efrgP9N+hb0oLo90afR9/KwhsDIdUCkwwBaTwsFNlvtb33zjxWkvYWO1h3
+2l7gYmBy/AJOTvceQdEYIQtsp5ATSxepUUlS315E/rCKr/V312YPu63qIliRJRB
wiKP2n8XJfPlpBAA+T6qaUxTaWKQGzDqPQNjHn4EEjY=
`protect END_PROTECTED
