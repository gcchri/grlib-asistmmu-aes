`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BldRdvR6Xq43xdmKywts3wQSYfrUwDxS2izM/v18qb5wzAckycC/icE8tVOkzIzF
GoHCNEiJQs2azdEOmrhiztF84X0fW/dIPEyJ/aXuqVpTrJxCZa0jA3njK1PeEjSA
D+j7wspefULhKmtoBvIFy02NSjkLAVKCtm8blygjaj96+shUztc+7m5745MAK340
55EAUqebhzOd6b7pON60cj75xtysj73N8eXEzP0DIMjpDSXsC8g/gbZH0kVBoZnc
uxQYBesnfsBcZgZdXJPHoxBfurbYovZH9bQmGOK5IvtRoSCtWMScqnmaUuItiBZ/
B+MPlOeCt3+2cHfUrxuePqCF1/xWmwve5VfBrdg9UCBIjb8gDiQK++mfDe6lK7TI
3mYFHLxIqUx9YIHpjN/mEm/NK6kH4jMrU7Ao1uidVnmUwBS74CRWhGA6K0wbdzUO
KweLhDoFJv64Gky/OuInrTE/rHZshTsbImdJY3ksqK3mmgtdPEUkGq+osde7K+F4
DxDMJ6/T+0E7W/kCpRBtNO6m3Q7ipiyLiPTRz00eUyVKNRS+mcjTjGFnmqn1QuTH
iljcTlBR0z+arXp5+BH182j9pKWTgU68WhlRBR3EEseIzSL4er849VYx0JJFtX5h
cVkFtlMOwuWKABIEZuyb15sMkVkjPGxw7Upc1CIEuU0=
`protect END_PROTECTED
