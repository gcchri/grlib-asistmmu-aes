`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHLBzzaekEx6rb8lk3miIBY9siWg1qKIhnlqs8gvvKKDXfJx8ndf24wZk/Qrz4tV
jcjobg7Jf23kNBhvsQWne0ApIBnKWY8NxbV+GVrWst1sq5d9CyWEkc3bQk0H/kLD
2KRDh4qlKIEJU3FUuI9e6UEvwqN3+rV62XRnU0LIs8EBGWZPSxXhnA8r3DJE2hvW
KUI7T7VO6HP99JqTNfbU0WvH/TZrGWvYK10RV85DDaWqqb9Wg9JGwwjgILWi5WZ3
eTfIh4+vOZenB69qsDhMGKdW/JS8QFXALYLi39PnuZgbHNSg0qGyqYCbVtRkyJ8z
8KelSeuaJe3dIliMARFOHw8n+rbzkdbhI7Ckl4EQC3bL3Bw0T3izmro46yexV8Do
wMi/XgJnKXz7GVWGalw3aSh7a9++XrscXEA5RcsHYE+NiZYmxv+EVtsfTpMWNn+p
G1rhdtdVmW3JiIe0IuHc7SRCGbvbYTeULupE6KeKIk/P3tlojjBtqg8BdSIijRF4
BESP+WqIFpSPu8oBW3haOCyBhwMnmYyy2eiiB1YUV8adD3afCTxWfpOpkBw6aPX7
CrBTJQvKh1awYHOFnQiewjsM1Ht+5zbK8CFGkuYYXHv5KrOp6MYC3bJq6O8RJZDs
LxGD7uS8mai5kv/c2jQV2/vbUj14/NdRE7Y6JmgHOBlsG+ygf7Yh5PwaaStUbRV4
YJVQJXsqq9JKB57sHAHuyaSrPIKO0Y7EEvnqFwbhZMJ6SNorD7vevfjaM3ARRCA5
UyxCT6ffsm4cgUpvGN1NdpeXMEalkGxTLUYAyOFvn5FqvR+UBjcKoGeA7kAnpEvf
dKCy3EhV56jbcTN+c1ES/9IbqSic/kkdiabIp+MjLT5ya5S0tH+dIUo6ktioxsvj
G+jXpEwzWQGf1qfdGweeNOs0/Bo3hRM+AVNLg3qG9syqhmEw2Vq6RhajS61G0ipS
3UxObtJVp+7QscQd2Onh4ckJFGjvEqCbbIth8VYTsg/NvStLVl4ZkXFg8poyfVQ7
hiMOMiMN9cGkgoQqa81NPvJkQtgn9gxohgCvfmXkmWPfZLhrm+6JOHf1WbyTqtIE
zZb40IAh/KGqMTPrPAXceMnqqtm8AX/Tvv+wf8BX0n8Nc6MSz2Z5o2oZ+ACDNohB
SjmZx4uMWsndKSzEb8wJzPenmvanx7UHpJkEjGikhvU4VvSRZi3xqA2/jIsywncq
cYkaB7Kb2mt+1sC+LwLTl7BF+zZH/AULpBYhQDQfR6U=
`protect END_PROTECTED
