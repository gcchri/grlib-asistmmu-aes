`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zp6dF0v+y2oHWrWrqpSCQHDAvuR5JwmCAKxUkOnApu5njtql5361mz4y9oq2lmRF
DTaIzX1iwLYtk3BGaN73JR74U0NpahACxJD+6FKfZWLoXaMEHP40cZcVQDZb8DdX
ZwkJ7dFh2X22CZ6PHAMYqvY/fdFXoFPxyeaYq9Hfmqj9i2leAZaoLSvc1kZk9Hzo
QiE+yDWkVYVqkgBHTtA8l7s4tojuuuKamPfkmYapEbOK9eixUhCVN5u0Bt5h0hxv
9tg/I/Yezbr4G8GTpjOLhVCP6YcD3Z+zw6tHiHY6JPYx8w9YUSLbcQK7ExaEO9NT
J+ha2UBVSWaO0d4iIQ/GmdOjUTD++OPmxm35Mu+vDybGJkag6xha2ZKvn42OOneO
KxI+AQiyUtOXnUzGGxrzFqEyxRW5T2tUffVkl++t2UUBsYxiIYc/4TvLVyppkRmg
r1Xqo07knAcjDBCQaB1yE+JKUHyRlCZ+PdLQvEDGmxUkaFOeu5X4wo8lzGSXLsMV
vlCGQWiQLsihhhTL3vb3AV6iVL9dhSrGivzV4szIyi6EEiidkKaZdDtPppBKZ1HZ
`protect END_PROTECTED
