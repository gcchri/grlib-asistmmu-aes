`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nSG9JgXSdsjAQvUOh3rFV7LyYJI5sCkZHZ/9BAjttCpDfr5EHY2QePqyE8DprsLn
Bcc6+ZCIGqcCzOTv1zW1xVLqAP2oNdNS5+ghxx4OJhL/Gww4mH6/wx1n+ELt8mnj
avdsC6KBAantCn09U8ic0syt/xHJDl+v++FRFlPHURCUPGl61Di/p+GJPyaRg+Bs
O9NLxk9VwF47YffhuuID7bd83IfKeI+iJIInvVWiDCb5jl+aOgQlWok/ZzkHP+i8
vbePU0kxaKjp+HtSFfIShS46TEcZ43jJrNu+WPJ6zjnsXvs97RlkvUEaJr2nNiIn
GaZwNC1oB0VjsC7vHIS+YT/E387SReOMJnNtTU2/VFc=
`protect END_PROTECTED
