`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cyFpBl3f2h7l6m/9vMedhffBSP5bSodd+V4qnLeFCAxCDtgvyGuEAJnTMb1Mdvju
0eSbGqQHm6R0FryJksAK4ZhnRmwNvjfrv3WG0E9PDwyquhm+u5i6hnGs7/HIalV0
rkXdL2GQCaLsxo/NX/ky9C0zZN1U75u5BX1UfR3C/NGabb78z8p9SAGJyUL40juR
HsIyzoV3IytiPO1T1KOoeYOU9hR9xfzsAsN6vX/KToSDw0UYnxfvC6e11gdz+1JI
29ouSKwh/cflIy9q5HYR5qqdVtxxmQc9tRDeEMlUG3Gff9XmQip9cV5x0SPEXE41
VU+urj9zktBH8f71z5GSiA==
`protect END_PROTECTED
