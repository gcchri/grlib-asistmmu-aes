`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2bDQ0dlw19Goqj1cPFZvebrlCKnT7wJbwA6XyRANpA4mIujEEXcZH9tGssYywu1v
eLF0t3WuWDrPqOgTq1EmtARAmZJ+feWU2ioLhUZS+ARItBqWXq1HgnMf4RCdKpqA
W2GE7635uXd2wNtKkI13lDvAJumiN+RajgrJorRR774dD7fzvI50rnXerp01Wt9M
Oig1iYNu2gtmTpIwf8QC8JCjBpnLQo8aTdEq0QIkA2yyz2Hp3GTqh7G5U1sDYJMN
QbwLliVALAdkewE4j1SawnrxuFuSLzTkHc2zVnc+NARWb15rqzoeGkoTMIu7Nh4X
mlJli4mvW08m3Bh0q5e3SYatTLZqCC8HDJnKXHe4TwWGQ1qKUH0uhLbRsu3BqhlD
EyYkRHKLyPpSTy00v5fmW1my9Jj8zg6bTxWk9V74ADHXOQM+IBuozUfHajM1mo3J
djW4lJsgf1PtOZ/Pcxu5+tZIqXJKcYSvjNj5N+1hTZwUiliQhZyg4E11PupD9yP3
zWjGCctu+/9Nn/1hWweVXhLEWXPtU3V/Bo8TAzA5SCE9WU+U49sYaPDvY06AaxHO
+T4DQ745t5VtgqLrNVvtMKs9xESCutMPEqMl+dVExr0hmIuQQFC+10vI10WmiKRg
YGTHHN1hnCCeNiapbC+xzaWK+GLoATFlZGGXC7S797DGlHpAIvXpjRSgVGQBlmJ3
U6nrHStcyo1kXJ6a8R3SQQ==
`protect END_PROTECTED
