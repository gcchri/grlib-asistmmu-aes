`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRz0AWT4XzWItdUBqjk1sZpZR5a3KTOJWyj8Ehca0y9yhRRbwrGlZV27l4kqDM05
89ewOpCssOsVy5bHgKFYUXMuzGHCn31HU9Q/mkYHFutbEnXQ5ZVGI0DUEKbllk8J
MEUna3VJHz4hpdIOsv7b0KbhS6xFotNPcLbYGgUTND0YGQa/R/L9bd3+lVDgH1dt
72CeFbaJye4Gw9wYZ+QyMzRamAXFKfs6QPX47T3V6Xdbsx77atHugFyO6Rhy2kOP
pa9K/AhuwEQ1l8IcHFsex/ZmVZlQR2e7fXE89SnnrSsZdzPzDokwbjjPi8VA6I5d
FNNwFQ1m382b4tAqSczq62KqfQQu4zKcNG/LeZzlzN2xdkkq3hff+2FRefHwxuTK
`protect END_PROTECTED
