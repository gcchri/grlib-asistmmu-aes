`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/OUSOdHeYSwmJl7e1LR1R1DnGrnHeoN4eBtwbFLqZRD03OQudjekJp/z9TT1OtL
SZ46pQ0j7hYyZYgHw2BTQR3NgkZ4mq8ak5gC2nlBKkSQIap3xhbFzBMha+rtuGsJ
E/3PkS8VRy1A9H/egiFfkjQ9z+ycGIGc1rfqq0wvQTMNf7aS5ZB90aj9ZGo7N2ZW
uQnyum8QnRhxDjy0DCLAHiWS/4zp8tKB7mZPr5GOwAKbBJ1vDj48eEdU9UFOwVsM
IFEwooo9VGgpELYaQzzQw5YoavZMxeqgRRndU5l/MCY2YmQl/+1qHs+ZEeh4LSIY
bqaWDUarPA0JnY4ZGtVFp16KsBI1JS6RFn6DSL4uI5tiR7JKi/NmlZNlFLYl95xN
k48HXrtP+LdzstVGqklCQKSVIVCQcZ0etn35IILKbaB2II4E3hnUHzz7Oqcpxy7Z
R81i1nFWxqnNRVLTqeArZyWKn8VEBgIeOwlvM10CudiW9+USMTO01nXGhIwfLoIs
`protect END_PROTECTED
