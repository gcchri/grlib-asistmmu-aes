`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JnwC5+eBCaMZZqVPMHQBldAZPakX5dK9oZ6hc/s2hQpMC+so+m/dG5NW/sAbN9ew
hp0vKOWCu2XVo9+U76mdSpA7XzKP3a8njL/ukgmV5ESw5JBQ6PvlxO/hLfzBZau6
zCI3WMGjnQlBcAMTvINotZg5Azz44dOppLLMHDPL6PoFnDsuRFgfvIY8lwZTQyan
fh4fmIAE0tBywlQB4zGTI8HgoCznvqIOckUj2l23JLkhwOQ3J9a7ko7mFdxxOFG3
`protect END_PROTECTED
