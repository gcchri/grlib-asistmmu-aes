`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhzkaRkAGzVyCvDgnrTxKcOww6SPwo52gffL4jX9e3a/iuimGNK02zUon6CtRi0h
jwGT/eP1NwQXWjID/YmsfNTXl8knPx7HbfL1aH1DjIKur6YIIpxqw2nI4iAogTwF
er8+JypGdJEq8SkaUtwUpeVre8bqdGzi156tV35vBalaoCHWPEUSaFJhJe73Aa1Y
fos/inVdlPeFwF+fg6d+g6qzr2R/spCagXuZDY7buCHXE96sTvdiPY6EVoKHbI50
x3FJ/d9vy2CKl/FceBxcuBjSXetpCIMSF13kpFPYux7NFHke0B22XpsOxmJpzpK4
2bvrZcEJtVGabNZUGaNbxrtWTIpowdCKhTM/j91gIEUsMqdKcsjKrkPZrhZQ2gl5
9/h+K4jLxw13tNvps+6umQtGZyYLOaLkE3Eof+KSPXLZqCIC7vSCg/494cVlu9CT
E4eR1FfdUVl5w9DE1ieNSq60mA/5ZCP1vR/T2T5FyP+bvD9HjBLGUfMI1TGrmDtg
d8xZs+HkDdeTCYy28ytmd1HODtryljK7vPylGwCDlkKeFdS44DEx7Ae/XEHafil7
uKLh/ly21hgZd7UW44pWcZrQ+F0W8E/i9PXMdXyNoygJpOe+L0BR6HXDFLVNfuBV
l6A2LtXGrrFk/xOeUSyWRwZCdas8PHeHlhJPefPzqY3ueirAMF0lYxudJ+YowL16
OagQjLH/TR6g3ZVxsJPniX1vp+0i8nC8y1bZBg5J7LBDNQSWfsGGbr1LgXuqmO+J
YUVPx7r1OlDJ/B8gKaMQHuYE8fdfEMycxZ8cPzBx4k/XRLai/WN7blkduR+8+16f
nlfqXLIrwN5SN7mz3FMY3OmzkXeHV3+HKBR3XleE10fQEEpMMOjS6zCQtuqUyp1t
ZrNrxFVgeT9HUh5ZQl51bLcKuPnRpT5zgyCL338R4orD6H4dOMJHrcT1yZAw2X9F
ZzBtXUIDret6mESffhJE376IyFbupB7QRiQXXVXCA0gSLZgdG6uHW0s/DQ9HVPbJ
QdQWvQ0kQe5GXSnpUzPmCBUaImGwdXPrt/tX/4qWoj6BGq0tB8SYmO/0nhR80Rex
WIfVepavxMiGs7WKJSA4cHp4u1epcI281sKrxJmFJf8JIvGRprUU+mZZBmqldJwR
AqMCYDfUu7CXoHDGc11Qhz4JU/uI5odilkTyJ68LPhuMQYSnAswe9wPHhbXOCbjn
dgxDgum0lAX/En1OiyxBMZOeaEbPEP+LWEea2VWsF16p2xJUN6PE7EvnFPacDhX/
089UKuQbMIwNn30FRTcURm9stnRZQvAJ76K3vFuDYKbcbhMXvTY1RUugPZ8EZmrD
zA49sW+q89pLE1DavcasXvN5mcB1+g2KeOJLWcickGzbozRgaoKtP81rMeYVEJiB
G/3FgCaEwlauCJrPUTDmDA==
`protect END_PROTECTED
