`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5JRtTHps0BxPXwm93i9RMOA3XZUlZYCaWKri2B0I7H4zJLVU+TRDTli2HMknTAU
m9d/fi9QnhYDVJT6rFPHMDW6FAPBJJGARaI77TaVolrYdOhs3jF0PuAg17fju0ZH
hzaXLua3eNpQpNFXnLggkmE03EKk1iWHITuaYpPV02Rg9pwliVoy8MYB0aAz5O+9
zrJCf1fuC85JEqH6ytyapV3Fbe77rlzHL9oUPHJGApkx1F7k8brOsfdNotDZviAW
+ikIHzTcdpuntaE6DnEkujRVIfzwyhImujC4osPd/hiyG01an8TcZ5nxdAeNjREW
VP1Df6bV/Murfz27WLzEU3x0aE6pRVsRHV9ghaVI+HQA+584glwcQ9T6ehvuR5ob
TIf9MLIQySEJICYR2m+4lXcxx5bEe2+OMdqepku3RnxXsAd06h9gvr8mYpjai9Bv
ST1ZeZsh6XIKmLZKSDgrykUvBFDTrCOZrQpWoIbODH2FphPOM6ZcmU6D24CqTGSR
hYd0mqCS0a5iJ+aBbbZ644i5MKe6w6h4TdPJ2GIMbPoFryIpZeTvLQB7oOhxAX0p
ieQrdb7+/u/2uCRGf9S8akyF/mgJW8FAI8EAcLPIaV/IAhN0SaK71Bjd9kzGolJ/
qOj8aMWwGztz3MLWXAlb1SB02jXN927mu/VrvxG7RDCo7QSD4MhSpv+6NX+9IjVo
GM6ds+Cr2SrwJb5jDAJf2vbanNw2PO44ZDwAgTap5MzFh1MywX7j0yHCvI0syg9W
TyyoJ5GOZuB9FF+nsFc/++GcgdDf5LIlQN1j416CDwIKBOW3X3FAmNLk3chdr3JB
hCjkie41RlXPV+GcvALM3F4AOf5+07cCyKfWVSKeCmj+cZGi4ZhQZ0ie+8S295qp
FV59mCLmnQ8wvAq5Jl6+6BVE+WUD7x1fg5O1lWAwfl6KSckDJF9r2sRBkT5CkOgI
P6RnXoDF1ibnyHuQGLBwziInfkiyw7O3Z0yFi4TxPc/RdN6ZlolefTZUJWc7TEw4
mb71f8aUVx6cc8pGPLQFE5rNxEwYRHzqDjZje1P95s7rV0htFn6neq85jAtNCqEx
Nujh1AyQBSthdtRhrETHaFVa4XQmHMtU/ToPPWqHkyxCWBYY1HzfKlmyrF4a6Fj2
eJLc8BAunFSa76IFaQmEF3/yGtutJ0gdYuWbsENRbXkuhdTyzlKNzrEiMH0NSWwz
AVTX6h+0HW5F9990oRQ+ZxgBTg1lsKnONu3Kv1dkJfgVV9iGli8O2FDQjuv2pFHw
tIu/t9EwDDbcku7pg+Uu9q7sqXLJvT7I0YjrDba07KWaJAbw6i3ZroSObMx0zS5n
1hum9h8SCCcGs1KliNZ3i60PwHatAe4YM7sjPjqUtDtIOxkpAFeS9ZKWMmDCNhxv
V8xykWhpMVUErwTeYsaqwoBgBZ5VtWBBCW8wTMVvCyUofj3t7SH4hisLlID3G0Ru
I0p+KA8L7k/YRnd7qy34xn2kRDTeZ3/C4cTX8A4Z3zNuzoO9u/MkxGGpgVcciu1s
jUIdEN3oNU8QHiXquMwtrC9xXoKmor2aVgsIOYwkI3HUfwh3JQk6kzzhQITtWdpz
qAqo43kGVCiy+osjcJga9L8U1wRp+jUD6IHTIrpvSeVkSPw92ivU+SLHbi8HKjE5
ZgoM1nVaHqTDr7AvLM+2XWMAMsPeJZHTlGtzykJAPFoZ404j+kxemSMEWY4omB0r
s4DIYWC8nnVLXnZx/oBYimWvsAkpi/IiNCW/DVe+R3sCcuP3qFDKf3KnAgJZZCVW
e1/V9t8DW/fLIi9+fhXnaMT4zqcVAwXhMTQj3/IIoRegW+ZOin7Dz5dbzpAbmku8
Ajx3D77WuHeYpg6KMBeyrg1CeC3skMCTQQGHcldHS6Da2bZ0hn8g9/yGR0SxZ5ym
E/fWV27LrN8assaACP2343qrpiCANNaSzQ9SUrHXFweMlu28uNFqHCPchP0Jn23g
XZILqU5SruoE1/D283ga6arVvrWprLZN9GznHaPpQhBSe8n8f62odABmKVT3V2pF
wwqKpdDn3ABECeYXWwo4nPf+Eq2boLWGSTFgckzMH+zbQG0v02SZy1bP3C3PqX3E
R6Zx43OpSOZ0EOHw0poC2LShgpxg4KDHFOSk5TFtNRRkp7tT+qkh/uFC0mLF+0rd
Sk9dKFKRu3M10o4+RjXmwCU8aKT+Zx29HzVjKR9wrL4S1lIQM9wQ8QxOrIFlmcbS
E2v1SubGH55NUNEe/NA/MsNv8FZmAN1Tio0lwc5RNmnC6a4TNpyOP0H0xwJakb0F
xFIohJp7cwNBrK3IeziWL2zmPh/5dls7kiJGBYFdfW432jcL2OSy2xUuzV5rCdaH
t9/IX6nQ75PEreuFzhUvEDR2xhQdBKXhgJmn3X+oWdKJQl/Dtcu/D7rATMgdk5xS
XO3bJ8ShpVpCmdwFZpS1Is2xnIJtZfddi+vEqpYT6tcNRyDmBMKTac0Zs4Y8Z1YY
gOjDhPyivI6bUHLe6Dt7euKgWG2ZBB8OSycI6qmdoEo2+fjHIuMwwztIU7pKJQZj
NZZanmhPSmlrkDdJvO9cpBFRGlhKPkH8dQLws36qu6P0QZkb1TvtWbGbFxkizt13
i82r3PrDwLwVsH1KQLIPTKNJPyxQK6ckAWEI0zkJM7itphUsHrrSXYFIUGhH+Qh1
smzFhPPLxsImLwUv++slFC/1EfsNjU//Y9BTdK44BU50VTo9Jv8QedAroAI8YQa8
RYUuxnvu9YH/QaufWuMEHvCU8VvipK7G5YH4W3vm0p+VhSzRBHnFfmGSS8cL6+vc
1ybpPwLj+hNL7cZoTnjkmQHvO1/Af4JtT2a3+dSjBO09nsWPElvqQpW7GK8KwBUL
M8QdlZdCRNKJyqOdK9sEu0nO60lnbX8U2DO8cbfILrospzteojUbh9eoKkkUJdet
Dc4sPDIRga465coF1nPN0dzK9NhouflDKGJtKV6mot73fREbgqWALdiscPPQaI8+
8C4vBiOQa8Sx9vB04gQ9fjxu4a4ZQQuL0J+t/O7020FVW/e0yLUqcF84dq47hOng
121PeUt1sbl00h2EjrXX+tvhw7juJQyYBt1DRvei6Yq4lMLH+SvSe3SZ7p+st2yA
K4FZEz3R/7+9nX0AInzQ8A0woe1X7Hp8OKcXQSit1pfEyUNUKlRwxDj/7zhzt2YE
fC96dHRe6G7Hxi8kEqRjLKZrv0SYFKbnC/RjBrKerx3qh/dEtXljjRMAo7dYRTyM
1U0AlJVZ0fJSIfHeh0m22A==
`protect END_PROTECTED
