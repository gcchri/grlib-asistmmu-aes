`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DmF12UB4qYZa4hMsPaag3oDopWQwXMpmt6M0PUtcUA0h0SrjLYnjLd/bMphah7b
bcRQkrZGXXJkqRbZIpu+Dfzr/wYpALfgu9ux7tD8qvAUJ6RbQeFZ+dXr9oIf4rgs
twMUiVBZggMt3KX73y+hfmnJCgjwDDDeOc3By01HM5VLLgbduN9lmxxdef4K1xDb
WrnNQsY2hMx8EmXoYTHkgs6cMzHNlVP24wp7sT+C0z36c/iN1VJrW2Sw8mfyhAqM
V/lKI3CeQJLWl3oa5apXT9l4dBtFC4Ype0At8jncYZaIe01iHMSbz7wxXynPd10o
zn+p8KufvE6TYxat6Rua552ll0l9isi897SWYQKpL+xF2PXTYtZrx+wcuVpHno+s
BlCYA3gLvJ4iIN8mptUPjmRONaNDrcj34cKRB1jzMVO0ubVNAv//mI1zbDa38G0a
PnSkJpMnfqR+fWJMfXviehkAd9cXt4/pzNkocBfuDYpk7sNkJ/7RmW450oqPX4kB
MwKJOndLTfWcAzdna6fPd/dPV1xrS5sIl/MZw0LGZPv26uOETgzxETQ8bJgxqLiW
nFFcZ1ukgGIQZ03QQ0JHNfFaeFatHLklFvUUR8/5oLXc2CCutPhbpYb11iqqK8fo
yaQr/S0OzFfYp91L1urcNqYnv0f1+AdHHJ4t2yYPLR8vEW8Gql3oo4UQBos1iZSH
2r35yxmRfiJcVO1PnzGNCVQyOxxBUjesjhdc8qd200h/SGSn35ew8y0sN5rxFQqP
w7mUAGBzcWgypALoEdrcY4jHG0JTAVCaRT90xGuLdPRcPXFqBZF6SdyBx5Vw8F1K
ijuzMsQrk81XvrHTFYw6COoyw3iuv4OS0BktR9N7WENzg1mYnEJLmVvfPruFa/7y
rQjUQvs/t1KCj2WKfqbOHn/xdExdogn7NvbXPlUr7vO1ABbPaIwophYtmrEcnv+v
QNLe8BEMHWAwKEfUkwIIOGIpebBaDaeeRsB/OnlVZh8SxLZ3Pn4ySTLf3KzpRRSm
Yb/DnD9vMsyuX2BrI8bOWFFMQZZypoH8vJ6fo0zoo22moiJMVxlD87IUm/tK79KS
5Mg3ZeUkWA5csep831XPqw==
`protect END_PROTECTED
