`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/21MD60Wfd0XSmX//6AmpbOya5LM8qzxtZz7DaUhV9HuM/+14YL1U8jnsrf4zy4n
CAW42ubLW7QfCNk05h6lScUBHWqgDZOue87pIXE6OwVnzq29iQniVobPXXVVcrjn
LZPvUxEd1btAfNooEWRrOfll1yQ8cQD5fJtk+fjoXX1blKu8eW+U4iv1kOXecSWT
s/4CiX2qDipC8zkxahACJIeDTUSRcdq9w6RXOmLVnfQONYr8xOqkEEKMJvmrNoxL
8navqT7aAup05jhWuQxhyl/kGZR111ul3MLCChJRoz5PESNeNuyfVZA7ETMDsg/o
EktL8PfVzwILgV6UQtxuw011TC3XvipH57MIp5FjQBvtS5aKMlb84t3klslNGbWo
pFn1OdSoysg/gnogV+MSD4t/hQ5Dski75EfUoT9KiKOUmQUmKMXQNrMefTCrz5v+
QucgTB7FIDiNa9CN9+yiM+wL4kY08yBKuCTw5rR+9VA=
`protect END_PROTECTED
