`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E3gaJ32bf64mPL0Ifguv7/IoufX7CEfLgTP4SLLGZ3oqI8+zLXrbsuTsdLOB9dgt
1QMf1S5x8FNb7JknTFmh9KvEwGU/Sx8f2WDbC4HJXbSTF9iVQCSrb4qD4N38c0MH
fb7aVWwR2UL8rVdrCKHKibkVeAtzfhIkpCb9EDwyyAOBTJVHUROmHi3BpGY6DCRY
voVVWHdokMtqA9X6JeL+olt05erUsOD7tKQPq43nrnSg3CpIgxJMKi+YTWR2Q+El
o+l+kpu9xtrpRwK/mIx4ITxDJT66Ejvvzy7C1PflYMCOHpnvgaWklFlgYeYU5zOM
afEDFKn74lTxGLPrtkBDAoTcfh7hy+nWzSj4mZXJvBaISHNYgz1jbs4CCO5uwsxH
wqpV6CQWj4BZ+jZ3VtVoHIR8C/gYC27CCEXUao7L+qStedIkI9zGH/nFW37frzOD
ZBN2iv9GqdZrzOszMF0HLTkBORNLtrYPDDW9eHyRJE3JodoaxdxHpTGmqZzKfftM
BAaRyI7lDEeFjRe9rjuadVOf3a7BXZK+HgSpZHR4pPYrveAgxXyI9ri5fEZvFwbG
jkQsyS1bfNlg0nlOF6lf0kI6EeIT7oupH0y7EiUInkA5hWCmoR1G+4wUUkIgZgFI
xjSsqHo8SEvgIHsqMNW9W6D6yx/EzsVslwpxC3rGkEwFaqM0TtZkpPNm03J7Cn0z
5BSHRx5ck6n6NGIbgI/YydiPUydAxZ47OgeoB0lHoV1nuMsdTYDgfbJWyr75VLcR
S48KVvemuUJRs0lkr4Lg4ka2YHDRLaEaCmN0FQQWHGKJxcMDV4UmvSSbbFPdSpId
Cdh+M1pOBf6iK3KI7MGf00rDZknibPXO0IGH+6uspJpE03gavwS4nEFtVsD0hP30
yyAMkIo9ufDDZmbHqRBbXpn0X59CUy7DcPasAZgoTGp0cvF8ByHU6ViFFC5+xNd6
`protect END_PROTECTED
