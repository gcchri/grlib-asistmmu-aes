`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZqTX9hdq236RLr5L3fvbqKpnkhONoF67RW8ZIo9nc/i5f127OQzFA6vyasqbgz3S
vsHd0cm0JwIkueWdFNppUTz5R7XOXV2zUn3sPE3UvEfA7cLUcIp5lMLs0hggGNL5
HRdmsfLXkIsFLc2BnP1hsO+SOuR4npHIULECWJsChcMyk1YmyfQ4W9VuIJ3/MKkI
mX1RL6F0MrKwGOZwc2jSJp/DQgNxCt+v8ClVCaIn6i5v9jLDKjOIxYUV+l7DOI2x
E5W0dHRH2JSmj5EIVLgi3vfD6L5YDsYVaSx9BvAKAYuAncxu5bXzDruvG1CSwztE
Hdfa1FzkXkwreXU/X8ZRPdxDxhe6pPpURBedPAM1QzDmD4IHc0Rk4VJ7jul2TdMf
3F/chcaLv6WEY4fRgSbJsxtxJPn9DxOcsJbZktnQqrlL/e8W1u47IWPpvkKGYGgb
ott1TL5oVQLZxu8Tjkmo/1qjoDthWmyz0k5S9qtgApcIO8PQ9A7lzCRoIOPSgKEl
W0MRI0982M7Tz4Ky3IHfhQbBV7rGLEo9yoEQhYsepVZvi0KSIYxLXqUfLvQEweev
0V4JOhRshXmiUqQqUHlLu9JaFO8yZWSuofuJVMG9bGaV56A5tH840idsCP3XhWBH
vQWK7GYm1a2zowp/mWliaxIToMsnbRf9cKzlnxgXLbJBgJOZ2YUmMiGsdKZP8eOZ
60/1Zsh6TiRpIeQfnsiI9PMdtJ+aRgTWlvzf6HBSubvP8PmEFuOuAzM6ACnpJfJY
qQKgD2lAx5sqUr949G8mzGa2LsxSJsmJ2wFTVb1boX9TFijcTSveIRxdmnFPY86c
5YRzP9Ao8F/73i5bkSL2Uh0DWgIWF1rOTCTskiQKBF+sFwyLF+xYaLvNxye8PH58
JUUVcT7MbS8nyR4nza+IWivLPEtmQ3JC9wCA2t9DRR4HS3RqHTD8DJNkl8yzQ3eZ
`protect END_PROTECTED
