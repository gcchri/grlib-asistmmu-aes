`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
COIN7RmI2gWedHoq3Dt1VvolHu6HQBPmNjmowLrbKampchk8wKhCZjbnwRJQwCra
cWrpOUvdAXvhICvjs/eqpO5tKLZIMTU/BCyZXznQXRjnzrPcxqXcHRL70YvlP9eh
7hHJD/aiY3V5pXF+Q94sXOj+rb3u68FvAeglCHrXm3JUwip3N7vsu5zsnpPDaboM
TpSblwPhoP7Ig3SK97qCLpOYzeBlUQIoDe1bDLUyTEqPegMfYTHrFUFyXgTQHCje
Z22vPmvB/bZ6+J2Dcw31wzJajIkQPl/FMNASHEm0g+8hpwEAIwMnFME4kxvmqCsQ
bzsdb2KPJtkSURJiHMTJiRRHzrLveGvl0MkCnO1gvxndAH58n0YTMq6riDxgePTq
BjcqRVgAYDistOGBP1qoR9HwrdbgaEkx6mnf6HUstzk=
`protect END_PROTECTED
