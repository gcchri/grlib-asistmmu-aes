`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwjB6x1LrT27JR0AvTYagyGjohKsjr7aHtrs1cpC836dfW4Ad+MXO5tScFjsT5bB
jBZYIji3L2yz5dRKMFNDZnYH7J27Vz3L2ct3aI/+EBpsoVB3TU27PbKQhM1oyUWP
U6+LVYDKR++j5XU/X1vC0AvZXE0k0Dk8ZL3rhhC9RPpoDApM5wwoG5dlvfUW62MM
t70QwiAIjiSux7qcUeW8AedxUh0NSLXPRLCyIHSp1L7c1uPvSQuVcqX5krQJPH4I
lUkdEbi/PPMpUEWkOkGANnnX9N31GFdeaGbQiUjCI8x5YJQweHsiYP5uUGsWsTrr
D36kDn/Zv7701qJrA2Ng2uE3fgg7Un/dnJyiPa2ephZDJEovIu9t6yKa2kINTFkE
baEA2fZVw7Mei4W8tQ+CT56bzl22NIG6gWlW/Rm6SjY=
`protect END_PROTECTED
