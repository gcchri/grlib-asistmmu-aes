`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nZtNIPou4iFJbo6ZAiwE9ol2Xv7TdwZCJpPLLvUgZ2+m9AtT2/1b/Twzf3AGwecg
39rJaFgDVSe10fKU7eKvQ/Md+xwF2LhBCO5UjXmuoB2xHe54C5nipAQ6Q25HzfoH
No7GwbftNnYFW87AroGKpr4kw4pgMzG2FZElq/9qYVUr2/XYbZ8BLGJdCjecdt0k
JwLXaNX1KGnL8ISf5/zSdZbqc3lWIW3Qw5yLwpkAjnQFaUITTVAXyLIFBZdZoi6Y
di5wGtolXsLVXbuIDaRy8QEHU4VoIXfBeIRNB7iCtrnIF9kIQRuFZ1u+OT/pydAw
Dwjruft3rHgPKpLmS2Y791Lg8S+XeefT5is2QjCYfqKCFtb5HNm43tbVDTrOscW2
7mQQePDYAko8o2Yoy4WyWCpGKhv2BRgOMXBjufq6qe0Akr0j4xvKP5WNgG4FJNmr
yHxwE/I140ukuzyzhsEzrZoRWzgjPbQQyb1UZaA3yDmIEJmhMLp59W2bonwUqAz2
cxYDqfZEoIZ6xrqM/O9N2fom9XVHORtkAEUTBMHSjjn2PRYLPYhAmJvizN6Rs3wz
+uMD3EfWfCT9P29JaDAiYo9oJNwk/M+AoxQ2DqYHJ6rlMVIvk2U/tDIUrKEQbMMk
oDEKhnXp6a4OUF6Bm2HNGPhSiZjUoV9JihiOihhZgtPTDgttA80jdgZfwTM51hMX
JCEJVH16CNKsXbPJjiKo3XR0vpDbcUVZ9RW7Qmif6H+4EZpsh+uMxWQI65ZHX/vO
SahL6KHDbvLtAvsLZVjUNQ==
`protect END_PROTECTED
