`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOBZkuIQ4ABVxNfDsOPORJpERYw00IYYvVKQhj0sSvWuVGNMKAq/7xhMCyD/OxbL
pNubk7Itvcvnt1xDvrBGlgWUv2tSReyCMXW1qMifX6dhvhJKkCFN2E00xjMHyFYp
Aee+GWIYp2X8+Uyz8xgTt1RzN52uG3+2ifC133tVEhLLOnfq9hgCK5B71FzkpFVs
EngMdPhhHa99duZzzBX7nehilflpdBnTU83v7b7KDYUyVxiFpR0RmQSlZhtAbeh9
1qvAXinQUEdbkGPDdQc4nf48qmtQSRIH7k/YB7N7a2POaq8YjP9AaeMnAwd5oG89
`protect END_PROTECTED
