`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lXhwkB3zpwbfl1f6zpzdOQsGBlWvdLkTpX5gBcYGz12TVATYopQ711CRwDFqRKSn
+00Pft/Fmpl0XNBO8THc1cQRQYH4WioIfnDrQ+rz27p75ReN8rmDvEPht4hYZFZb
cpkDrrVKV4O+XrkrbFSgGvNZTzGQHZYy9yc4CbmcWbn55XPxekVgoxW75cB6jBxn
mtPUj0n9488E3BbzQ9QblpnXNqMriAs5UUJ/NZAL6OMewwm14cnYEHQvX8BUchH/
3mwtP87MrrjnMnmryP2vphGdK5EPFZPZMbjTQ85+oj5k8GUPkVtmx9RN0vSZtW3C
2vt92IpBSFKPGfvA4IZ69abZiMiUbKzDdw+MCjYLdeytNCfJyan2FL38UnR0J36R
qot09J+OZCGvzxLlMgOnqtPfZV1JqxkeP1ODtejMuh+yb0eTwghYYXdHLu2Zco5D
4iZFfiOyEXbE1XD2aH1qug==
`protect END_PROTECTED
