`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uu2JEG65dlCiVqMl3+qkGlp/5iv9jh/fK4uVMbin+Qz+Ga2k0e6MBwzcG3jMjDCv
ar4xlQblynDWV3i9KyiKj6Z1A+nQS6euoRESg6koTgTJDDEvOYa5lwmP3KSjAp6a
56aZgU4EcU7lZJKLG6EBLvE8tk1bq4NcARji/glnhhFOk1sp8majX+ojaWBXz606
aZSd61cTc0B3t/VvyWDSNcTbWrjOtgZdjhKpmzZECVFTOMkMp1YOPKAkkAXNdVPf
8ZLZ4Nele5cwtSwO7HyfqtNmqbjMrjizjUZsQVI1bTBXfUOugKCJVLyqr5KhTmgF
TTXEe6i6r9Y6C+LvIsF/wNNSZfIQzYN3JtSMqmKFF43bsV8Rz+8bDb7nIxR8I/xE
eC63O71G2DA3bfsu9hL1r11qXMgqeAx/51g7TEd7kZ1xf8TxOyl97viZ6j3rvQkZ
lO8tDCsIt4Hdvh6ZjYLXK0QXRv1WZgycrarWn1fEP4CvCBjVcdYMDKzAqytVjZWd
1vhn8djND+zhoMID8Ao8sGgIcWiDrk5Yew1Bz5/0Ac5nGyYwL+m4DjRUitPLqO6Y
y4Nixx4+oh+f8JGTVXTNiBI6LTIX2bMboOnYYfhWU43UhrocV7qD0oc61qp1tRJj
2Tt9trsk4hMmeWfqZF7nOSvhyEWzs7I4qiQ0tNkY4gqkD7AxAZH8lglEmzdv9t/R
GPofuV/e/s2xk3aAZBgRS+/nxelvHSYQoK0xz782KKL9CRvO5+s7hvduyw6TNq8P
30/Xw4ZwvAepRs5fFPYAbVdB7jGgNcoS09fZvjjFCWEKt99cUH1TJ31BJinv4Bds
H4/G0fE6++SKpT+x+1P6ckvGWa8nfgZyy2RnRMeeQEyzy96K7coSO9kUmpBxu+zm
`protect END_PROTECTED
