`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJK9AHBJnBloyI/sNMhG7tpUj5N2tlkyn7S4ksPY7fLuWV8D+c7blbik9V72lMU8
e1OompENiVTrAbQX2t/wcntrtSHYbzniHPk27XDc+bJkJLAUnW336IrpMmTSqsVq
cJQSGe65JHTwJ83PjPaxcM0hS5dQyQ6GUzQt6mSUkEklgxmpJDoQXG09DTqTmM/9
ELDd4XFJmCWl3Yg51LMIhcvNMaJ7DNIgDmqEGJ0HVeCY0v8n77Pzd9qiXB54VVGN
P7EEwuA0toksGqyqYRKIkUE4WOI7FkvUqUhmac3I8pYaEDHvtO4fPaIr319dXsTY
g/0pkGj7zXPeq/jAETA1l5nhBgxljAodelXzVNPmrbrxObr+RGwbXvDvOsNupwT2
aRhxXFQNEbN0T/f3Fm1WNPs3xQD3MInIROOPghZOGtPmmdoZQwBqfmAIc48tuEI3
uTEiej9uOTcvts2IPaddZRp242oNngNSXtuS+dTOGM/n77QCfdd0HZuAcW7JewWv
Rs7cSyHYbHnsIpCIwqSnK/RmRGiCmvNQP4fyItfU5A9Tqxz6kXb5MvuSkWPoKhA7
5VyFLBgtvBKukW4RPNeK4MAAVvMSk1vd0LFC+ccd5uDRz1V0AX9blCRuHS+lohZp
daqnm8joLJ4MH1XpVVRW/A==
`protect END_PROTECTED
