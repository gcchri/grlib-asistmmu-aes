`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dqh2TlkKzDQMOIzaxpb4N2slwo9sO4pf+IbnzJL/u01JrNHpjwGoaZuhJMMMon4X
lNRUk6yo12N7upU8EGJEjrLT5ZTvoyb3OWBerBXWrYszGLEOZWRPbyhOawQ1IshH
L46Kfc7sYdfl6ddBTpGRpffiJzsFEW4URxrjLPs/X0mF0cpFC8oOlSt4/ZO7OoRH
bCSDrhatil1tdNTiYFotpVOVFBiJLRliVCDxgu8C/i+B+Z5njWeBFwoRNn0rN0xr
iF2425b1I8rO3tH1eeyKZFCvP3iZvHScfZF8yHrCVYM24D5oWO+7cJ6RHn+TPP0t
E390BeuNgiUWCKPso5q0/ZzSW4TyfEdl4ScDhWwjSk80SXORu25jkxLDYLZKPmD4
qCArw+CevEJ2mdXfWPEQb3uTmzuoNj15VAY1I3nkCG90MQbALYbsWP+E15ubowBo
uqT5aEO3fco0HwfzME4ZIePlnQuTHTIzvvi8wirKItAtJfQLiqicIBJeTMhsdO3l
ltzU3g7wFxTWMhDZR6oGtgamswXISQFm0lRC6Xe2T/FkSwCgjSVAyX+cE9RfHal3
vG5Mzye0uBj0aP2um7cHAaVU1JCpZshVRDF0ULGqo7PtoC74Yrp6ut2BtJmDmj32
l/tZ2GhVskoIJttmThI8nW9RBiOmeV5vMHL8WtNCWK+ShdzpME3TXponF3+WGWea
KhA3/KbbPhxJcgFLaHywlH7UjXqWsKKgIHDmnHmg2gxsJA8L3kq5/oLXz+u9OQ4a
2MtGAUc62A9hQx5Fdl8p0WnN5Q33aL7GzZIVFe4HRWK3904tmzuBFKIgg7+75bgI
aIh1yJgnTQZCG4f8zZDfmdExxjqtWt625PE+FsTXohmbMUKhB02Z5fp3IO4ywcyS
k1xGBhQ3v67PpBrN06slLfudIyTcY90eJ/KDnq0P0z5eAx1GV/UfhJlN7rIN+TQf
V+EgXlQ+HWOLsvd9NW6V32gK/FbdapmuDKdFqrWdAshfzMEoNna/ljFkJ8o3jcgv
Q7XujDYhFwV5be1+uBnu6+XGZLIk0VF/aLPN0oZzWtNQR/ExyL+NkvfjqBc09f3+
vBs6x5fCP3Jfr53F8efry4jDeOxwVAVE7NK3NDM27JRutg4SK8ao6fqQrfIcFLQg
QF/PKI4Q5cIaDYcpOsju8UiJ0Zxd3HTSuhGK7WsAdjU4T+CT2fYecsUi8hogHRQ2
TRJFUgNk66352HWiGmJ9Khj6BvLcCrWUYmt7uBkpJfCWGYBCw84pW4MEX/oNc3jr
voTaFQpY6eYkVpdkmn2tEzXdbO14t8DjXvhti/jKTzbgHGIVsYhurf5ff05URv4B
mH1Gv9y14yl725nQpGOzDX0NggyeyIUc1DcEQPbfbbsAQ5DBJAPAwHHbFUy4anmy
jfEhwheqJs+kxJWZpsKtE8GehTnx1R+9QO8yqdIn42M4dlAbEoVAC83VZOn71Bwd
PYfkCrQktY0fbQNOKGMnV7QQqaE665xO1sYX9O3MlSwEVqA4WqKxPERUvno7LsJC
X5nKnfe3oR5lKr/+ZrzenfRy2tebJ1EiMAbRyUcGuqpcs8xahS0GlIBto/98VMD6
+qzJDwuUo+0q8xeFvUG51ZAW9fiGNb0RVSDNKsA72GAZHiXZCDuVtXaFFMeQvYgm
8yboimb95WCU9RAz1NQACjrQh3lMug+ney0Mwd4Sck8jAI1g0g8VF6Iz3Ygvt/lD
NvwStMRvbdGXqPs1wcLFqG0/8Y++b3K35Du5PA3xoZFyiK5882NnNm/cuH3SWFll
PG9O+GSn9qn1l/Tesbyh/kO118AlrB/0+n9FAOfey5ti+477VuC1eHjNg0JnLF/9
m61xnxktpVa/HkYCCr8fpB2fBAIccmg0PCAUGwj5N27dkbgNOSu6IwcNvcKzjj/1
Prus9FnM9JPiN8QIlEgnN61Bhj23ZtFXwQ1Y0mZaZEHR4Os5HC4sgPyxb6yQ8Alr
FhX4aOt5kTs1bNZ3TnmJKqvo0GTBoLQ/Gmea9ZRy3VERzf1F6LGFzGSM/gfwglpK
gSjZ7yZdmgC5SJL0xfBi5K4ujQJhTpYl7bcTzXRmLSt26mYpZFoFDYG8+TDOsxZA
VMhX1awOeeRGumALhEp1eSL4vYE9lfhWh1JJiE9ysPxhPrIIhFSDXWvFSQaXcmUk
MlnXUufBDuNUW2eDv+7Ag83JvUqvt4nEQB4BzuaFMnBZyCuDlbPuyquWSou0lgI3
pLPCP+xEXhDkpGchKhIUsTn0nwZjC1ZIrnk1Xw8/HhRaPSg/drLbD7hnKi+pN6L0
kvTdxzgraLj6DilNP9xhD9w0efVA9RAJvg9/6FRSj1Ll+QRtbb5SUO3G9LQpFqj4
VZm+YZsX8ELugpBz9hIXw8NGq8PM375AfH3LMJ2Nx36T/NTB0gV6qz72ayJiLjil
TT+1yKZnTIEqI3gbvyQWDSQt8AGQKPTCslRP64lXURrDOAtCLRc4ye4D+NQ2/N/Q
5YVroeULxh7rvk9G5UmmgKpLdmz5gzyCw/hlbRmbVQDXhWTflRDPcR+YlzrUEiMO
K6+fHLAY20UUE/JtvLB4zX5YItZXgUquWEtWXa7pjuD41lzd48g3P44gnxLI06In
IRQiUgcjhsRMWXi/DGRYbZxqZokI7UvfQRFoSG69z+0NAmns0OEGE3nu5+RbEtNx
gvhSVawN3XTuvXyOMXfpQdr4pBeNOExKz1YT2ROcUFc/50Pf1tBKAJC0yWD/nOGq
bWgjmNxBvnHXOUMFmGcpgFlrYC8YX7wf4Pp8aPJMq3xP6DpjeB9P7fEqitWGOPGn
XE97Zj7T1IBMcGgHSOfvlTchCYZRl0zlL2CnJWFhLz/Qqffo6rppmTB8KniJMT3H
dgOr6SSrav5jRHdPnHHIsjUYP2cb6YzRHTp5N95w0sMOE0IOCM/LF0pcOdI4jRWh
uMdbmVr9iZkn8aGDDqKefsUksip8vT7zFlGLiHEffcaWrNQS4VHQNYiyEdotP5tc
zeZs1ywf5RQeFWjU8RZWNTtA6D2z0vE2ZxwGlAL4UURCtRSWQ+rPWBlwx+Dv/U8c
3U2mXCgy2Tzik20Qp3voKj3ZjXiywGTx+cPzxiLeCuCQdYwQ3pCbO5+e/MjZqhKF
9RrRdwy0eynIIorRje6q0XK43IQvZ5ILrwO27CXUzrHF9lKeVxc6xDN+reJGty+Z
KRakV5+994Mgg445RHbsflE9tE7kVmfJp6pxO2ezrVk0hJjQtXVM+/TjguEsMcRG
4bdSeLvay1A9VKC4jWGAphv5Ch30StVT/0zN/0JHn/Q0HN2MchnfBOmhxm2RcTYz
UbdoMEUEtVlSceG3Z9act11UYBizhVSQ+BlDBodGtxvijFCCI2PyOIHPSw1igMyp
UnMx7mv4Gt6TT1v2kbjnhQmeKnmGhw2DGeW4OkTEiLyThGjDieQBH0IywEoN0/IB
3tHc6zwnYVKTrTk4s6s5XRx9nVOttJw+mpSnjDU+da0YFRYBJOjd0ihvMoqKNjXF
l75nnJiDV/vMXxa0ZiBMA/2Ug7IDabuAjTjUVcWCG/nen/NqemQ9WzaM6Le3SP+D
ux+O5O5E1HacymY2gjZDeaDYHDA03gVnT8bwCLDOpRJYx63dgMsIm3BRVPDUgnuG
P7JplSdykGah2SNv5169ZZGwN2lowUEXZ87gJlCmuJ8IIzT0zL+bRpJybsiN7+Dt
jSjWD/qVC3JOjJxDZ+/64iRskRzd82lRPQkGQT7J7Gt9O9xCQ2L8yCKEVAxGlfU+
nValZrpE3fgexBYKePkf3PcOhDMO0EdNHV8q9s/gatc5ztMsBJySA+7AYMwg4PGR
K5ErSyX1zj80GPMI3QYFHjoUMV+D4A52Cck5o4FOTCpKSdByS23EclM0JfOjSf7d
Ma8bJS/kLmxUbEUJpn4mI8sopwpFW0q4uWZxb+Z5IdbOqPxM0tlL+a640NNnQwZC
FYgrbWDxNN+XJJxLkB8ocdnnCPYy1xTAQs0oUpR+Bgwsiad2mtw1l3ukzpbl6oup
c3DLkKNyRBQ6iC/rLu0Ke/kKLQhhEnyd6dE5egcuPK9FR5c9zx9ag/hCv+Du4w6/
hO7wmOOC2gSbCFQH2AZZw2n2dC52+ZyivesCJ8NiGQk1DmV84DlF52cSnNDEoxbT
3mUzXkEnn8hCJDKzFe05Yn8xozHQVBN1gRz6OS3yRkRaNT17ElDrBQDA8asIAjLw
vx3Wh1uVJeX8tXrFUmFO1u0NzPra4/SsbRq8wv18EMSp30k2vGLwuVscli3K4dyM
G5rDa6vIkhBciB+uXzlBNoraPx9Ho8Ad6oypLq2RcjoJ3pXzta8243CeYVphiJ7e
DMngoJZtpK0abUJ+5/xZdR1mjk1+WLsPyEMM/BB0ZdLIt9x5dbEjPOYGh8Q5Bja+
OJfVO+nRSL4GKOWDtf8GtxUmsIc+z0GhE8Bjv7ywN9OgX58lVX/9f5bM/PgQyao7
uMcNJJAof9IZbOZZ54DjpLKv+QQtwfpUewJ6ExR/7u0mDC4H15fuDyruxFjp7Fkc
TR/uzEkxDX2kDoFAMBQjZMqNRqh8HOZVANh7AJ3TSoCsVnjCcIejVMCgSDdVoZph
74tGfEf+P0YAjK7g33gu1aR9/0oArb2Ac2CTDiExDQfRsySIXP24HfKd0DBCcCU4
WV3KYvIWyMwJMtp3ZbHor+So6ttAFmgiJ6O84akoz4xwABV8177QbHiL7x16Fo+Y
NyeF6dzfekt0TvOk67KcOHONDrz4hgWz2JVeSRt+pReVieVb+LN1jS0fgQmjX/GU
8/5TX+sIVXWgTG8KCgb+1Uo7l8YxWzaozHF0IvJHPTZGlsLUnthJtBKpRYEC5nFP
mohCRXudgzaMyCOuXh6y1atfC2glfBwpXhMdcdYNpi+xtVONpnkvs6Fo4oxP8SQZ
3fo5SlyqQP/dZ7bESBIq3xIknT2D78Dic9J4O5ASzY/6O4D/gbqpGER1Ws+PJ8bt
QAVYXktbGRFHmFwJ4SYPFmgp9FsT3TIsKMZBFGZDBcwGii4GvJqpoSPv353WG3Tx
UqP0Ii/S07vZE1G5JW6zvdCmHNmQXyhdAKsHt75g6ILJ1FR1nrRH5OhyGUPr2gJq
scJncz4Db2nsXtJgNBuHtCVv5nx1uvzIqLC+HUlseEtBfHCIRyfysFcYJprBtyMz
c6OaunhM7Aqp/kKN3HWNUF+xG6Q9ArIICJZ405LObvQg51RO53dXgi+I/mN5oEcE
FpZbySqGGCGH6qwA2Cks3Bi/vRDh9RnDJvWyxQVzyzrFS4Z+r1NE2bNUUoXb68pW
rCTBY6yvEHmJqTNMKC1K1mfuIuL/5VmH7qY8ZeuGMsRCsTRF/dz7bZ+u8St1OzN+
BMFpAgxkGr3qKPRpYxxJpSsQ1iY1dMDTr5X14wuJ2Hnu6B3HOf4tqQbM5LyIWMCm
rLPxB5Z0XiY5ExTVemEkAqkJk8tZTJ32eThkBDdzRDv5U+hSgzIG8ASR16Pn8+SG
jO7aW11OeEdy0VW9c8mLIzlTXxYzL5ix52wh/mnxyYmxJJyZGwPcfQ9sQJYick+F
0GNC/AQFTwZ+MtlYP1I5Jlmb5wfEnEpvEgKErnRN0KxoSp14tJrLCxJ14jALD3UJ
NBvSgLSAumlg0Q+IayPYpqfxovdVLjbmB/bhhYNViu00w7ZlEgiolZuhLeM/Nuoz
Ouo/jw/BzR8kJcyWmLDuv+WcFWWbYf7X5o7DAH9q2hUpRzfY3sejd+EhFhLP2Eoz
8XGgVEKm13fpF1n5oAt2sBXfpRL+JBbsVpAxm3bJu7rV/+4HSLYiZnQvdj/Ckxni
vANEFsxIIrwKociRl6RPVpkkI/ID/jKhYZFk9+mJE8ywLOHJl9ampxbsqLZCGry9
vcc9nvy/tdBGKVrkXbEo4fzN2uY5aXZXTCx6cGo1V8lnit/xWWcnYDoAQXDHb3R2
HIvfrStzqc/LYH/8u2czFgdcG/nQAosraLL8bZQ5loY6kofnkkEC8KaT/4kZkj25
B0rpwBnGx/NzmyvolAY8Wzz4UN1QhTOG+LlLI77TQMOXDp7ybMWUji1tsuA2M1sR
rfc1CmEuuknbODuyOWOBQTNXiQKZNLLUhiFmwOjvsNJCNdvuaJs4YEGmaXGVRNCo
5ZP2su3p2I5eTrhyz10MAAQAvJix2RPApADbvNce7ssbsfPJSdg6uhuF1BNo458v
K7YfvuYaUrdcU2KWmyNoZ7hgcT8HpaY8Tdo465RtjlDEngN97lphyy5q2Oj1lSPz
aFsV93dt/XWcsx8T3s5hOpPYZvQrP1f6+2+z2jvyXWtx5ZSFg0IYgEBBKTMzhJTG
jlEVbFj9f88ibeivo7KupiQ73capNRthoK5QUYPIEYEfXbYLc9UKVp0BY4VjBWjJ
gRuBKbsnCP81ED+JM2Kw3FErbAwG27ntctILA8tV1gih19eZZ53uOwHpa9L1WUci
+fojurugDaOxyzNnpKeiV311/6XytLaKQ4hcl60roRosTTVCR2br+GG1R/JLvcbd
BDNAGQsL5H8JHKJzdyZLnizpIDr5DbBZtxV7dPMq2S+8m8sqy46uT0WESiMatPEY
xgvyGcGv7JUrKA2Mlnxu4h2kG5/NNmda+t9DH/rD4wsHheTZUQ9KeaX60m/E+Im+
JvkJIYhDyACFsaFE0rTgGDTVOlx+Kl8QIoxVIn9EpzwgwLCiJCCMI43HKpJVK9aZ
MsZkaQL8OEr/UvOvxky3W7y9ZNmimlo7ZP5ij53+YiXUggpkmL7q40haqRCot2bS
WZnD61BpDr6FcDZERk17h8Z8jGEGtH4jfstROLHBAnYM+FKYTIVRtC/thnHci3xD
T9Ue1ObMl0XFO/Za10/ApV5r8KqmZCotM5U3vljf2VmBKrmwDcwHq89jNo9OwNoL
3WePu4brrtVjPVmSsYJFTrqenmavYpOMEM3R3+vDCoBwNiEIMVZ02edlqJtgQ8tD
FJH1+dWB0m20He/WjAlYWGV5rE+Bq1+YYs9yATKPEDXslXQEdAWDPWL4SU2ycn4U
VO+hzun3K578ibdD4Nz5PPalUTPk4rJ3F5AeTEOCmkiW03GXJYAsD6CFy2DhLYzO
Sgg1k5diQZSBVIsiqEKZBz+7oZeUl2+BMNeUvksXzGbp7N0MJK54aVqTMayDHQ6w
MYbcI4jmWRgQpF9VFnd0qKvI65pRLyw+kpt/v9AJ6iZ0N+4z5Ni1K/GZf4ip97gy
4NTtODF1ByeThPourA2aK0WqaxOe2ONsfXopOyJ6I9/CRkCXeosfAGIczY83ElY9
vqpY+aX/zGX7P4ZTFnKIuOe8FQ4xZsZpKLj3EAQuddLYaHffCyDnOPtmqSK7EfBD
9YKz6oZqHZf2ch4oPgZO3tBvc2KGGoM12BDJLPl4OBesoLliE/c8ZjuVvyeojWIC
BPl7KOR4b8LQP3pRosA2DlT9qUjfAXwkWhEh9isD2aD9r8Rngb8jUD+rRQVzlPwy
PX805hHdF2gYbSrGBDnuqjNUxPr8ulNNio3QvqGauLN9ptq398PMuIqFoGIMuQG1
gzUK+EN3cgamF7rjsFAraQGBXRC0znHP/sbHdJs5zgm7AbdkceR4qqyQu28sbiFy
lgx7XbMMSgi1fb8jk8JcKJ70Qmsc/nH0KyUxSC23x0esBM+XQCaNcC0MKjUDyi3/
WyKdq+WAys+mHJ8onXwPeaxS/URKeY2xhwfdpDMmHYSq9RV4RgiJnqqeHMhMpF1d
32o2Dqou1l6OfMaSsueF2qiC2nlIxMMioB/heNrdCMQBapif1duacSpaZjsxqoEm
9nbEGtsuKB6qZOG7jymqLxEJG2jhB9pkHLZsopA1ku9YMMQ7P0AdGiAQHJmC/Eg3
8k6XuidgLUQheDcZJzZTN/mgiWCRCSFDuitNllDMjVvyq4DW6pzFZtkSAnXs4Kpd
mmaBFTKvBF2E2J4ZuQ1c69e31ZsyucCBRu0bS1Bc7UOHGHIUgCC+S1auhaA/sp1M
A4KKF3VeoFs/qSfpKTrtJ07vu0ZSjkZA1Zy4ZyRRFnvPl/xjzAmWC+dcf1a9sbQg
J3664BhR5nX2ZjFH/zLexIgBhM0HP3uNbluxmFqU8XwKqRdsQLREpiogR4K33SZu
b77UgMLvBpEpdbsU8R4OcvKePO9QW3rq1WqRUKqDigsKWYs63Te7Hg7oZC8Kz3Hg
SXVsN5fVLvQfslQEmjrwDQ9JttRIKzFDi566rzyDdYpZ1nzzyrCmbTS6bZ/m2viW
ibwZn7gMcb/XaygSa3sSeJxFiQdQEhNzztJcQFQih1ZNpAJRmfde2OoEuNPv1ymp
OYlwAcxKGvimhFN1BNmyzq5pEiNSIlUqO/sBYXA+1Ve5aspY352j15kCKfuNyOwc
pSl4SxCmpZ3gV9NvSau3Xj2NhyRoryDO1dVrkklS9nWhvx+lgXofMPwyA8ox1wUs
IM2/D/tziixlEKasa6Xrj8f7xxjyfIt54rWY4Dt2Bxw7iJopqv0h/WgKiwfTtq6r
B1kmRN4d4DHORCG44W4/VV6cOrbrKSJdVXKAXiqdmRhidBnuMJGG79ad1/vG6YFk
g5ESoDq/C/H9qTkB8W+OuC2aK+xwG9bM8g/DpqFnr1kyZv6bVkaXVQ2McyQCSjGH
9vJmfmOr+leNxWk9neutiifLSYk/iEUs0lBrtLybTbO5uk3I/yJYk5MJcOwh11GV
aduq+4i40lW53tYjJhCuJg8ilzAxNSOY14SsvHhsAM/dk1S+Nmvy9Q6mTvICpXyW
SkREPZEFdM+gQjObDuT6SSoQsJgOxPx+c7G1ABWo52p8CgQWPHfifFumczCfnNpm
pbPfcZSOS7XiNm91PkeWnrfdiD+iR947nqAet9u2rqEfdXNLKe+bvXYOtp9ujjA9
+1GLX/HZygkaB1/1SubmZ/OaIR8gkm4nxeF+8+nfRVm4itM8YUcSM6M9SO+21lvQ
LKQ+JI4pzzKDi7NnykG9G/SRJdCHPufiWKFF3et9rFhvTTokt5cuACu3njEtRJfo
pRFWU/+Xdmkf5WYLqYAORQWsnuzDw276HGvDBGU5sZCSXypFmbDc2ii4NYTls6MS
P4PipPFAEV5gDH2XsKWxSLlTEOgrCPVWG8fvbupx6/VnjMI6zA3RCAvd2UP918TH
Gkx97AwK3lK8pftm3hkvYcjPhPDxmob4cZUekYnH3kX932PElfs+MrkTde08BFWu
i8PGyQPIIWY897g1INR7KfFJrXg+pAeldhh8nbKiTwY/Q1ShQk9FWY2rC93mIqwP
FPrNLuiVltxDTBajal1e1Hw+5jZ1L4DDL2w2PrBfoTuBRS0QJUQJfe8+grGvWS7Z
9gL474m5cuUxJhbsTn4c6p2JIXSHA7gx3q8JwqfeMl8FZ973232yWV0YRtVox3T/
vaLqO0zBHgos1I6ETwYhXsn8qkeRC2b1XtGYKkbFghCgSh8mgDEc0w7/nulcwB0K
BVx7vqS7gbO/DV/9+h19yvyJqn+J6jieDb3M2oAMC0PWO1eJ+Nu2fq1kyPSxld4A
GY0TOnq7VKZPmY1F1/1lV2LiQKoYUyMCscg8UViRMK2i6vWLJwi6+Kn/PvNHGI5D
pUA3Y0FwRUkFtE+zfOMxk1SQvF3kquTbLaADHcuy3Yb2Mdwm50QDkdgyuL/3J+5B
tpJpRdZcYHYKpxbtdeqenAeKeAtyQ6lFEGXH0FDLe/VBvGDqurECh2d38Y0p0QZD
1tyLVVdkyocYu9dV8UbUMtz5HH2eqveedhAd7UIqSORn742quS3VNdfIwokXJb7+
Udzr3Yxd8LP4G4LwYyj7Z/A4OiSZ7QA6UKl4ecjjyxd46cjooBXfhTEXk8HA+EQ8
h0A9E3iblsZD458mlQb0vB/a1IL7Zz0a7A+od9m81e1rlu9pHhOVMrOi9YG0GgRg
7eT/ffjVpj0QtYZ12e4Ac72ahTScZJjdgNuU/yfkL8iqhX7uSayKqL/6YXy2gPLl
FqnYXQMgH41Zu8bRDGgA05r83bGRbZJ8SRUhUTwuRtqCX+++ZdYNEvC2AR2O2cYZ
glwVxkR8212fhG56Y68W4k+wctLsDlwJ1yslCDMUYqQJDBjrIlzveg6kLuwztVA+
/PffhNHZenFyqgTECE7pjzlwcXi8r2cjApWewzvtO2tqyMiTv7DTPW8NbuXLXMXg
iKfMmkP8k5aYL1ys+W7hWzu48H1XJ8WsaqMomI6mGb5w1/0BPZD52iBVJkMGDRy9
ANGcIY4NNjk8DutFwg0bdHpQQ2bEdGfpq2Gtg0Oc/TkshMWDicB+qsUNaYBR4SNd
euKBbL8qMTXLfmSi71kQc4rfk399ViVOk/Cm5ya2DFO6TDyNoRTVhcDUFMcBnd6z
hJXxMgJ8ravRv3MtI8C4VhgvE+QdAwUtAYKB9ibyHJqSuAuS4kitBNhi0T+/Eogc
wf3kEXqIz+jAgFqAswYiLAKWjBS7VhcMo2PkCudZ/8Qe8ym62ejFmjQ+VV8RCVFL
jODwtcCTDLBndYWImFUqpG9ayo7x62234fiLmI5i/ehfx0ue9Yu21savpgKD7LCW
Z37O7vzBNtjB7cYKOkckCdEA+xGk7tch5xpSkVaSxGdPA029Uawzr9ssNF2gFbh/
mOVTdYb+qtME5HC9agh0uALJiL9F5apMMerb54B6TVCExm6CSRbavAWgRipv1dHc
5zuTyYHYoMnfkjXU5ORGMRK4RQGwuKmi9giIcrr/svxeH6FSB+wKWH6DAZkjDOfy
xFDnaccLHej0v1yVfktxG2yX4njZLkTANxgBi/W843I2fT6gw4ZqdcKht1yQSV7Z
Vousr2zaD/WEJJScREwqLtuUdncUkkbTrokzqf2olbi0F4fIo3UHKeuY//qZAxtj
rJfm5FXtHbId6YxoPdL9IwtnXlGlhP2NY1fYQO/U8+ULWPWTgc/dpVEpBMkxT9mh
WwIPrqOuLKDmhvD52Nq0ITIsrJu81Txlfi/7ja0hiXATl/PUOITKF4+761xFOSba
E6oX7cVBsnFT2j6UMPpKwd2LlDMolKx3icWLs9as00LbAkuW4AzRUMmaigdGc8fx
i8facH+NU4ivpVmJru7KNWfJ7DkfNpHfSpV90fSIWlqZ8mXAGGt/kffhvJpSEKSf
u17UkPCalMusJnGABndPQcLwb44DmQKv/TckDvGd3t6EO1y91MOOdtMFHBLWb7yK
jZwOr+zVfapQZ29UGZ8Rk++MIxjTBSrn2LOfrsHpHqa+EIKsHf3zH9S+k3CpNdWQ
owgj2JZ82Sppo5i4pxzLutQbPfKYHWfmNhJv23MLcGnErdFYLEJGsftozsMTZHxQ
t8wdUwjAIMSEb/XDpboleVR8wib4sh/mnksJZJu1A+6F1VITYDIVMJzwxPYEnhgK
bcgVlH9C4+iA4feapv9Kjs3jJsXu7mQN9toIFr3TwOHPg4JSFnnZID1+kMpcPtYg
09MwRHEwCZcs/SSyE+e3F3b+ZZn3m7sd5JfRdOv4CIHDGQeBovEQw2Ge5ZkCWbQB
rfgnp8HMCWncgq82K7U2jOaxW/w326ARg0LkXQ4xf0lgc9KqAe1M75LTG14EzEIT
fTl/aQZwowSqPL6XuVGdNfueuj4KSLjeXguUIVMT9h7MDSvPfXpTbLsCsLcHovbk
MzgnPXWCKxWUen4fvZ8vNkgLPPuReSOh63anaceRKLggf/zGM3K9kXL4nneWzsl1
qCE5GWCdpbVRPkSWyVmjS0BliIJwUpk0x2NuyZLbtjBtwHXB0kl5NjupYmGTdxMW
iqtoidIuFTxI5KXNh2ywznlHeJBNyJoF1NjdeTDESTTPh055h1uT5+KxDUe1vspe
t+pNedU8fYkzrkG3LzMU4HdPnuArXgr1Yb13hjs5AQw8cHdRJFFhTkJ/lJoDqkzz
k0GahRBZGjjnswpyv27bcUeKQM6a7TF1h4A2n/FjKyuV7PEpZ8H1mPMDBwqt5L72
HtLkXfxLvov/IMASoOloXuYZjMCLvfIiYC355WVH51GmwB5d6Md/5qJpPftYo6Yg
ALdat3ysgGkUzwGRb+v4hudMNJOaoIXDG4Qwi5iqCKKG6sDxu6oIxO+fyXKBsQRy
nIXkgpsR3F+HvMPLHYkplVn01NRHFfF7OhV/hIHZ0KL0ZyqOPxzXnVhaWyYY2Fdg
zVOcxFMH28XC9AUl28FMOWY5lqH5U9axwj5NR+gR/+Yy4H8BkjONFzNf5GRlfmAq
v8zqUJgZvSPzZGU8ICa4eP0A+rO0GnyUQDodZ00cGj4fy687zj/RVIogEJAn4WsT
qJd4V/BD7kY9II6nCtI5xrCkWOulCBsG68A9EP3oEegcSmZzqWu0s1ZEC1OjpkKK
HlNO/16G2Zv07XqHauKwE/M2SzzosroI9qDcrMMGRDjscjS87uBATGaXZ7rlFj1U
JdbYrf+iYBfhfM9n75otBj17RPW1r3G5mMaBuiSnSq18tziaWKIVQzaGs113yvyi
8i8bkpTOrF5BtKrH7X/CzlAVIThaDoqhcHgTsztvrldO/o2/MorwK6T5eKu08sE3
hXC2m3Q/GamVGpckRlQU5TD/NKMbFgwM5o2hEmzBE8prNa+RVu4EiIMGxCGnlHTz
l1hQu/Xl6dJkP3wvQoY/cQvR16sLWe7g9eRFtiNpZY3X5+WdXNv/t6HyYWxN2WXO
PwVESNRKLtEFeTIU7DZ0g8nqMGyu4gJuvpvRnlb3hOKdKAT9slbrGRJ7gmweGuum
AuZ0xM4Un3QkjHiwgQFBqNfwgX+c6qgGgDPlWUC0q+0UGl30MKBc+i7f/ihIXlAR
0GL4bNPbn3Nj7i3R2Tl7woxQnak8oiMxltaQ2iqgGYGW3kdbNkPTPGvXbtkhcXUB
S3y1kZmiADoqBq7w0KUSenft+6MgRLgyv9XDvLqabqMPp7ij3sMhP/QWnIvBtiyK
cid0MCVP0aq32NI7CW5eEYBiMQeqJgktBPf7KTAEtb9dTHe+8EOp7t4Ef3re0abe
qulRI9qDzBQWyKvxNu8go39z0xteUab/FVp6zX/x35ihyNNP+lMNmPFk81ynca+2
eyiN9jmk4OKsJFrk9HAGvk2iQBcCaHcbb1+rbMa0rob/Y2dc2bxFqBHnkVZE8wtS
trGmXGlU1DZQmfqskXegG2o67xBHoHu8aLuqXgsLOqK/lv61qtc2HkA+ucFJRqK3
2c16KkDRU3VGyZUV5q77mc8u2k9cM1T9KGo/DgWgXnZxxanmGb0u4kmMO+RZDQ3Z
OdZQqn8oWXcWteSmn39QQYvN5AANLShPtMqqTBTALdUiBA2JWJf8r5h2gCh1v56N
aIikVYlHdZL42NixSyOU8zbsKHRXsx1vfMuUNhXotmJ0IepWxGvHa54TDcQDgrtq
00l9opx1rmb9bHbjyTyuST01/7JVTWTCxbuEMMVioGlBfMMGJmrS3LB8K51i3nsR
zZgizo7FNT18uCmuhKjP4jNsNmMVwJcFcr8mCpOXIOKSZoj8krESkWhr4ATyRNUX
fjrPMWCTdkSRA0fyUwCXCPTNZMT2Y0WaFaPVa1XX3KwDp49hE4ApX3VaS2QIMW/c
2om/fCG9USidMFwFi3+ZSxDfK9dga1U0XgeoA/O/fC50DT5NSuFi9CKPLXfgqMaH
abSnBzB2ESqg4MLccY7H5xLrJMxBE1nIxx4zDoUg/+6oBeo0NRNEdYUK11IMXGBM
2o8VHtl+CIDnV/pf1HrY468ZVqiZp1Wxmd/3jhg70eM6IcIHZcbxiBdcN67BRJAg
JOsuShUGBGYHqFqCUvQhC5xvvyVed8IDccByCoU/jXHH2dOuAHZvHrmNcMNXUNRG
AR07+lFOi6tNk4vA58QmJ8yi8pKJifL55afll9HFpGA2t4v7+BYXLenYCDVl59nI
OlfsB8z+NxWztTTAIu5me+LgHi1+9Bd9JHS7XhOkRBUOOe85SG1mLGBSGhJEMKfe
5kMRmBSFzpuzDr2alPIO72dox7ojbf7/5kGybWc8SZ9Y/pmKEBh5kklj2ZtKZfDk
MUZQ/jOlyWgeLpuBCL8qGwZkwyY0kJeJklBkuVQGniwaeLAotJsAaO9lTOFnUaIz
PRpM/GLeKyjO/bTHh2WqoL5rfldwbPzRLVvuKxybpT2E02rVEsClXIN2j8Ww1J+z
23JZEHBoq9c2ONt/uIUrAvH3wegPsRLT9DR7UeXabHjrP0VUADNBuXVv5pA8TYij
nWPMEMG56QDXfW/RcpysXrtH+jKu/ktFfO9WsBDJbspa8p87MMhGgFGqxEFgGwwF
5MOiKZmkS92i1DEOBLnfpC1M3JjlGNqDP/brlbYWCmjA2DSfqis/647UnD8N+jLH
CSlNJeBRp8PFPH6abmBS1wWvmI0HBtuGmQpCGwtIOvuWEGWYYAS/X0HB0qjCdhgW
57Y6M1lop28w11FvL/BOCnr/jrBJOdmZwdiCduCX2QAhV5rxWNSrG8ZWhkngu/+P
Oj00EyC/bSK3rOP565Kf9SrRMBRBfSOp+RvM05q6iRpr620NiaanAfIv1OKP+tUl
IQeDiZcIHxs+c8bpy1y2461SLKr3XiZxFpCC4r8ABH7gCa8Z2E2TfJXWxrCFz6BJ
yWcZzxz3p8KefFUaW6RxN6699qBSLOOUXPOwqk/25XeIfYJhukPJ/A18ifcfcJsx
jsaL1QtqoUFPAw+lK4Nn7UyxYvyZ850MDq6AmpdHOcK/mYSzumMPyWn+BK+y5duz
SvH26KG7wgr2Nu0SXTuWChv206MOFjz553Dl+/xel9CSZAOWq8J+zMxuWjDJPfO8
X24rWVS+dDCbH7BF/xO1vFxed/oEOjXj/kObkbayFsr6wLP2zMTxkULpOlm1j+dS
3LkTz2+A2DxjseuNwIYJTC7MnogiyBON1HntoGvY4tJKrzguJ88Jwn4Fk8FwcSoL
qObWaL7OVH+ggvEIUBODvAU6ZWSAZQnvivAKHnBDi79+Koot6soXA+3SELaYUiCG
6lPdFnduqi3lBTRsAeB4rclgS5TISVC4naqf9Kwu4dqtk8sADMxz99lDeNFrcEo9
VcaPxp6rvPw67GA316WhwKj7EilizkonY4yQ9SrhGAW82YK51++OVIhljcztZ2ig
7UOt6vChORc7W7SOikOiQvRs+cbvxsfYptYP+HjcmTTiXDqmXVIEKGsXLctaUFvA
a8BXk5jNeiNkvol8iQdDwtLjA/msOVoE3wk3p9OOLNUXJS0tsDXSRjFtwnN7WwZB
NJT8iHLHXc5+CBDZSGB2t1vTBseg+IZVlqetmNV4434nfYQP8xkKoi+UL0CD5zCH
1dmSkgZ0PbrD/+gns5d19L2ihImM/tvn1ishVO2ivjh5ZPlVMVKaO/P8t89qXMF+
6numqohWVZacqoO8SD/YOVL89Yy4SSCsmQvEbWKxnitgV6h9YZdF78qUzDVVSI0I
VViyi8Es3OpIMsrCM2qW3GjH5WLP/8iT0iB5GbhMsfkDEHejgfqN5KmVJUQXYZ9L
jRHIT+yz9iabMTLyGQwicPtj/BS+nKYhASxNHg55otS1Kho9l+1c6tAgZVVyHLcJ
1SrmBoHGCHJuCpfmxSJaTd00FUp+/xJ+UvkhVUhC4J+4T4vCJCdTr2VYpB7seIEf
+gyJBhHknKELcN6gkVJa2UUaxHvkMhSeP979n3YrRww4IiCema4Y8zpdInCo42nv
osPuQs3D03tIXT5b0GxkSJJuMdvJxdhowC+ShbltvrHGOLtqF0Cn3SvkWB+CmAbL
uTHYbidIQ0k2kWFzMon53c1Zns8kkvvsjZwgPFv5Z54CNTHpgt2bhQfW3sTqyPki
Zlb2Oj8Li2RjXVrlBoHze6MYIWV8Bh+3UEpYGCQFTdMjDZieikNq8qI9v8D3bcYx
x2ClLEE02rSPjwpxoezTrwJLU5FMaVsmSfOSfxMKrE6DbsoXsCrzoOGXyAq86V4a
xMWEmL+69kDhkYNadPOjJNxqUOpUekqDOYDLUyljquDOT6/913w/0JJCSnhFgRcQ
CBbvCsIBR+QcmOQrqi/kjMZLWAKoORI5WG3xYVdzxE/jCpn09yvjzBEn36zOQu2c
C1Vg2MqMXb0fwIDHN3LNapkaoMwZ6M3yurHLF+f5Y/ud85TrlsTt+T6Yq8HcHL0P
4bsKqqSNzEQEehIHBygOTm4XIAtdz5UPtNCsESnO9P6Ag+M5rTQ0e86ObcfDQvsz
pCfLHsH3/Rlwc05du3VHlVkEh0DX2tZsyx2E1mx4bDlA1ldJDp+EWUxc6xLCkzM/
/KZC7B3oV1CkwYK0cWUZrK0wpMrB7PYdtbTwX01B320+MGxIfZOOX3ynkoxqmLnV
p6QBvVGGbi8iEV+qLiV63wBWyUQhu/9CxwtJhaJNcSHzM0557cMrqO3ShICXmA+S
Nv4j0P36VOno1TMYacS492ns3GTOoiK67UwopGV7dLxfLcbCYMQMshv446kgXSpT
xf8fNl4w+msgy1ELrN+sQeM8P1V5VsHnAtwhSOoRLAXvu/XJQJhAuHJqNmpx5FTV
fVfrwkyVPPSShXnBq0EpCDuJJTRZizFLWplg++voH/J3exp9Vlncxwz/kvcdp2RX
WPa0hjhF5X01bcBoAhp6genB6no9bCos0NJPSCn1B1Z7W8Jqy4Mb2HF4p84HwYql
LOgIOAvl7WaVwRwgYobCYQOLnih71FXnuZfQYUvIq3RkF4VX61hx8xU9WbvnKZGu
rdc+oyFnWRQUQZWz+gEf7GfGNm0JNXJKTPtUN5U4z/9pdTPFALDSGSSYdz1CVrUA
hOcoqwtzJ1aoUY4kDv9Vk4I+XSY4EakWTCu6Rn3KduvWmVS+Ar1lVjoaMhYitzR4
++398uLvascqPjDi8MlPl0QfvsxhLSpqUD2Z1D18gpZxPP8CjqbICDHotlR7Bt38
C7Ofn3qPwv/vsFkGXgz9HgST2510TePa5P+vQGDovCj8/DwQFpjnE3GsB8V1ER3N
jM1tdiVUFYiGyZJCFKkK93i+Yf218l+4/Cx2vGRrgq//CGXuLKG7Wu971i4H3twN
Q1N9AzuLaTN6zESf66daInouZKNBGvLxPXHL63E9bca6kbHgqQaj6is5/n3oxNtw
r1aEOGIhrxhTunnsdKDeOpP6ycALkDJhkcrBaGObUK02rlCEG14HNa4OK+HfMloA
82dlPVOpt/HIvtm9jUnzQKoWTi/EHNXVJ34qb+SrbeUFa+LYnqC+xQXGTEY+LkN6
jSHpDI6fzMdz5eSxsOWfk7qyRDk99X/1JSXL4dzJ6aJcNMcBAviBG+ayGFSEaz4V
WMu3VR/b627uGTSSw0ePq3eQxXJ5MlqtOwEFd6mpFI8/DuEhLVrJrdE11CgzEcBg
8JDOSqotedCyIdLVABEwDZrZnCWvrgG9QpFDIE+KUQCA4LCO5iH5peYAb8+Sgkuv
H7krSelEnro9Nof15hbvXWhSLsMcN35Gq2zB2A5DW/SyXTgFW/QM5drEvwNeOySm
ozyH9NBjGp9Ue26sFQjO8Ff+ZZF/c66ZGz+3s75kBLtOxbX6rWBta+45Drj8NWwM
ZFVKxDkDDXpjK06VnIfSrJPj/iCabBkOBh8Rb81TCZCJEWk5UKMbkNuIcyanj8Cs
QqxuToou6mBWORbeHmERBAc5esYte1pcgcOLT7vHHkMwk2/DErow59P1EefdRXPE
4nzJvOttRCmjOxgSllx/MCjxZAhKsS9nZx0BiYdZrkOWzRrY9EKX2VzFeGPPxBCK
WVhxG2nsLnEGBzyR4v+e1Mu8n75KTM04soCNX7WPt032ugs1YK7Q5OA87gVMNoVh
fMUvzqU1vxPQTIWkkLzMX6Y3im/DHL92PLWNWdFP1MM2S5WJTjwruO+a+N54XgB7
I1DeY77b1kQk0/QOg1FDNwZdgI943JpnmSoogygS0UI/LE05D2uHU0Cb7g/cf+cS
Qjon+fNIz/H6dZFrJbHbJopFc96uxkvMg7FmAmT3oJbopilwRj+Jb8GtznFBNL11
Jbz132e19xaaYSpVXW/rCbidwEtpsOA1L//1NE4inEemge70J3IiXAE6vpntrDKW
HmKJaBR67O1g0JCCknADJjQ6WbIeWkeTc+Tw85WMy3hPD6IbTCHKaIXBKzktqNx7
+4EFFyBcmkVsMBCoEBoG6Mol+oke8a9XsgareM60Qp/uceXGFTynExZf1yjs9tZw
ftbi/+9MDkL/TorHFq/uY6dDr7WOUwoo7AF33CjHTKBnYaOijngJxI94TZFwgd5U
aotlSyOPQGJeSHYj8ioh2dZNfApZ60vyR343EzpMXto55fd1oci+VPNn3DFiWx1+
JNl5SG0TizNDDBYLhxNeV2KKmHaiIKrMb4NQFjdAezV8QW6+G7zC5bpRqAppHJch
0cygv6Ed0lANy5+A582PxY9XRGr7ynlWPYcPrVY5ifc3IyRv3ogqTmhwyJtqNwWZ
FBnZVf6e60BBRYDlBQzabYXNFPPzbnaQNRJML6U06DNNXr5tCfHa8116HqIRZ64T
oQWePBzhFj12YKBSrEhcRf/htycCdAdp6AIausS92gSBvyEb4ebNj9sKFp9AXu0b
/j24GI2THZKbfdCOSq1BRB6uAS9Zxe/jHqcKvJl7xJsH7SBiCVUPZFiq2vfPIYE1
0TN/atR5Hpa8P7UzfLBSaxATcLfBfuVbxkxKLPGlniJYTBr//78SNy4vY7/sFw49
zQ2Emr3yfk1qc2p9HoAeeMjecddcdIxPXBAZB+dyEFJHyoQzpRrn7Iyxn9Lg1aqL
V6kM2b/r2DavuHzc85rFc+WFW4ahwpwlpRjL/734TyGIOsNvOMQSeg0aB92MxY/2
DMRHQYzb1Nu5Ji0SjQyNeQ3smDu45VsJttQk0cS2CkyBf6crpSgD8sax3UGmONTm
uM+DogTT2Zx4bsdrkm6xJbp/C82ZnHj70yJMlb1l3ciwCrZwGCB95tqOf+5eHn3O
ip7KJ1NZSr5qxeMcrQlOQY0gQoVLYmYb20YiqxyikvQ2dcseTUS3JBZRHC7lsAaj
Zsse/iefH8Hr/m+E4OeXuFkAjDacfldXl94SmAGCJJBz0nOF9/oMkT0ltcpBh2nF
Yhz5a90m3oMWSRW2rEh740sgEV+aJahCXhx6eQkEQVPpVZ4S50EpVuzXRWEicOmV
5MZjpE7ohUlBnsPcKCL0Ud3gvwjhXasfzYDCPoXXRfyS41YUeJaviZjLeCechYvH
o37G09nXdO3O84ONnMIIkU41a4mT7t07MD9rO5x4kuDJrOuvlL0ieSuqZuBEzXWr
0PqOL2PwfnxPOr4z54cYnCXVZznnzH1ExNqTrN4DQsmlqZYb1aYtamlSv/UJ4AQ+
bwHimfMD9BZBWTc5AmAmjwlWPCkQ1sBNM+l2nhIaEVs8vftonvWMqhszzTfb78ng
PHNv93tGorYSsHGbzKIheG150YegRyKf0XsygwOWXtNS1MBxaoPvgNJ05d1zsRx8
OmcLkUxOb7eiBMomR7mn6G3Hf3koIFFSpuLiUeX6Ye0nwGeRM5RlCQKL87xLM5b9
7qkse0I4RedRU4zVbJe1M4WmCMk9WLBE0OUhzanW2m8So9QIMA47djrIgX9Kes30
fELnmjnIuAcgGsTjJbC2BnarRLeuF1pmYL3+cbXR8ZhG3IcpvgJIm6bqVCSCd5nw
CJ7pWyA2wJVKnKjiS0MFWN4Gqu3Q4TkLZfbb+pdPI+C8pxS9Qzikl4uBoQkmFhYf
O/mIZs5RACcvPvOincUfRF4aBf1xP8S8sKIiwbBbiktEod4Ldiz2SyycVhBCErzX
ZMptzqfF0Sw9tc2x1KbZ5t7Q2/MuometbhfoDd8WmNi2U+01ohNZzEg0XjF18N++
hHNDPeRRo+IjWQlCMTc7Raz2vji6mPpJ/1euYOUtE4TJ2IZYnQAOlBZYsEp6/7qA
+bBp7VVx8hLgTIQKoxRRoXnqlaBPr16vntLdw6Y+1+ThZp0VFzznha3MvYiqL0JZ
Oorps5a0yVGHfq2SBZR9I6ckCPcbI5kPbDVqRKgyz8pMclQczQqfk5WrkvS7mk3O
UIg9m1VLydO7kUIxwDp8kzsr0QIc1pmF1Z3Qz90tAfZVisRGZTmlVyXWJIu6X45w
t13lQxKBd2WnBSWBDRxW3AFSnZUA5Ei60KsUoU2mKNpFk36p9kvdWDeTFInJ0QGC
lxze0vMsFynZBKXbsEPYUV9Kxkhic7EqyBGLA88lc3CjXHOTcHMXMWUuW9V0cteO
AGcuKbkG8SKUrBXEA72nBhZ+HxLkW3LeB6Ylts4t+kb+nw77vpPZ6j/W8dUx9Xn8
p9nwY+JcG1SFUUthQDx998+g8FSHEA473XA/wUiTQxHrWf/Z+6HnHajB6Kh/Z4zO
O+dbd4sjaF3lPZAU8ceAgona7ABEhzTKFXN1acPuGHFIZH5/IGCiViE/JA9R+kWR
mNp+3fitgKwEdyuvBg42kHpe/ie38qVYPw3yHbZiBWt0ficGRsAU64kPk67yenX5
cezX/Wh4zCW3o5ba0QBBMagRR46FmImCLlgRARSzPO8ciNGb+/S58UYgOORGHYtJ
GdMAGhy+g/we342uLV44O3xyNKqGOiCrKua35oJmZtMTWcc3yIZyMtSmyLaGr9XX
jsIMnnq7jtsMNvyBYPauXhHqg3haniROQvOe3BIjQX01Ew/WLC03IfEYtoFZfDxV
7Rp1iJhf8YefLiXeVZcI3nou0n6n28TEZPtcfix6aKJPfmVUfB4rJVhdbHV+TUNg
hA0JNX+yQ+QFmjEmK5WC7WzD47JhC45JITcKXyeqGnSgt6nBaQPTILGevDAMF98C
rqqANxMdJgtafGtreV3zZYYKXM3lpub+RyKPEeq5C1HEuSz0CZYAYRXZkrDTjIMg
Nc9ZI9rR/fs9ZpkEwlzrzzRybXTviP89e7kddt9jxh9v7qPJhQrt+sE1Ejlf9SOV
Zs/BXQH4A13xQsrTKPJr3b/4CNZtX8Jo/NwioippQmjtud86UmjEp0KTRThdjpto
Uc5BbeF7ROyI1ZiGlB2eWvCRg+inQt5xLLtrF7jrOIxjJUuZ7eMayrSM4ewu8YXQ
9UgDt8W8JlesolbUBXvIuSpenfPb7P69qDYvediO6D0hv/FRJJndrAB1DG/zqIzS
s2g0hVOVz2TF0crB6CGPZCP32nVrvc7LHv7rEV/VrdxYqYZcJhnsbTueg1RXv5VZ
nbTXBGiwV1a6b4pzlJe+bZzXZ66G/VP0DACBlTXdpkIHn6pQCRaT1u/vPdOWiAHF
DtnQXQ/Vb77fvaWhh+22QwTKBsST1FnGfCp1zbe5XLqGqrL4UAek6OvJX86T4a/v
3zp2xj5PhNhm0DNSHet4BxbiV+ujrokiyc6i483CWEBpl7lyr0JcObQ5cu6qVBHD
2dK9bokkuqeOy8Oxl4eSP+wgmExZKrbbh//znkcukZp3zcwWc3ryzxl378vBoNou
wKDP4+yhuKwCwNxivtXpMOiXaQmnhiRCluO1eE4563YHkajN9r773KS/GwraGZQH
L9Ys5OjAULqBLEJZQZEx6noaYcgLpBnlDURoe0qTC9WaabnPEP0N4esk1+muwphh
CREV3rugToIs4s0KIytHlxmETgcQtpuuh7BBA7Jy+QqfSWg8ir70C4uFjhfzFyTc
+CcYU9eUi5ULbt+bdPw6GijrY+VSc31oIm6bEh71SplBYtcbZiXaRGfzlJkDK3Ca
uLT161udZhL13/gCeEH+KDbeQDMwWYImRqTsPQIzQ8t2tp5cVQtUgAwMCO+xYP4e
BzHyb5ZaRW8XnvU3uW3S3I3cJJxax8n2F8e8FENuEzzEFHat19t2GERRJr9Yts8X
DHjINojyIJcLYdxZ6nJFIL1Fwxl2Df7eUB8uqI8P/beJqGyOpHZlHkFEKsnhLd5r
zyMz8uelvrftL+fau94hp/AnH0rexY7kDf+N0ll82UCEfMZ1N+HISCT0DN/0sFRP
WtGbbQfSq3lKz3PDcvYcRDi0/uRxTE90M7brUAzRKqLq3AiaYPL4xi6ZGmygJmfy
3ZoAiLh+9EoSlj626ujSXk9tbsiMsFDCMv4Sj2hgIidJQm6aduav8yqUsmTVD6us
QM42TFt/nrgZWIwygOvmvdx8x9Dnq9rKsis/rtQ2SYtQcQF1jehMv3njpOHLosUS
RmTH1lxcKpKtEP7ADljFiSM4mvDh5LG9C8sezGSiZi1CbkJuQItYFOE5/CCGqOH2
eKMJ3HKsrbO6fO8QRk0yvpHn1cYDSGskO0D1Ub5qNPbE23h1EYM97G+oD2Zwb404
c13UqNW1p0dFZiO+Wr6Snu+6Uy/VPdiZPFbLEioNPdSelhZuWH2TfITL2Iux8ueZ
nA+I/6a9R5sgUU1LaWU7RcEPei8Em15zj3yc5oKgd6aiA9Tga96HUpgHg5/sda4P
kRFQ0N1XCREKMzLEhQF6VUa/fFngxaPmkl82ZCAII83RxVGvKkq8troMBeT3wr54
EN6GoEYKbbcJPsu+sfUpeJU4r88NC6qqMu5co1Ja+yMJpvQ8/nX4sRqdTBld+6EK
muuj/Dj6cX5WOutS3rBxQreW10y2l+4FVCdmLpwWfXe++fPeA50gxwqj7r6SMBT3
gDn7zQhP+XXje0AWaL1hm4Q0QKTkzOPF9Vkfc9h/JEj3jW+05T9QU7aF4MZ+AWg1
kQUVXUePIyHF5rl4PXM2uKb/SI4/+Au1Cb4s+kFe7ax4KQfAS7heqJt7z6TG6d1c
eCvqtPdcI9g6Fh1yw9jJxf/LaQaWjaNA+Au4LSiqiemu2n4DaUYblnlU8P7tc8Cn
8tviK6AgybHBHokq7HlMp8ekIT4Jrcgq6WT7WPb1kKLrTmmBFlABSM7SSUkn2j5j
N8wDuPOO+ZR7uY9Y5eFssF7u1eZ8YgPY4vSczRyVheWC1uv2Fry3siwWsODK6QLK
ppA52GXjwtcd/tYm6RYTAoLeszMQfmzRl9ls+PnQ2QpqICp7IjeoCE0ZFsg7O8wf
3zCfusM6x/nHF+N7UM12nnpQ5Jptr3JQvGtukMwOJxNfoet0xAqDC4jWs7//c0x/
IerGXuGXGzWcv73Tqv0fgduCj+/fx6694Rb4HChILDKig1skpsJBVIRMR8KTaZTI
1MP6zmHw7AHVrLfAYowiNbafFiwzqk6r0irf9wQpk7qGZoliE/cw5a89eWXSjKp1
YxglL5xnYSO5pvKMzzueyzNlFzvMjoH86DIsYppnQIhevLxEkeH+QEudWt0MAZEU
Sw8ArfUawhn8Ew7s0j9DcLONEdJpnMJrXrV6NWxjruM8lNnkl2GkemelpIJsYEHJ
yRf1Euo8dUGiH0MxC4QRMgD9xSRNd9CEZKns65hVBs3zz9LhtNKDMXWdmA22go4U
yChzvMtPl6VVNTAyZmEXxxGIoW45CBf62J8z88l52D70Huir3wgi7tbIYtHPLuHg
JF2Z7T2kPKT7q7Rt8NMnm5g963m0jXXJBa2+w92SejN6bM/4yzEpO0VQJaQTXpmx
ofINs34H9pu4v03UZi2zNzw1oF9jtirTTNSPwWxjxipt401rxRzsCf0k67CRbalC
ToCLHvz+lrNve86kZd6WYd1r14FHzuAee29O55W5m/PzHn1T4iKwoQGAwcRW0665
Oi7Hoa8NZ34Gmu4SI+2yYXYkjgzKz1zDEMtF/5nDGsopLe3ziLP+ke+deTRvft++
kjhKKIF2pIwA1IZ2TDKd49axV+4AY7xN4pN6YOVzP7D7+CzdYP2DbUVu3W7H6YgK
Sd1pf3zY4UEjuquwb4aKR5k03UHhPT0ZDPiSEz2zq8Xhh3C57Ca3NptI668TbYZd
PI/GGB7uPqspKV4Cf3pz/P+hVL+s9Dvh4m3M9uxnqgD2ZBcEXA0+oyFeTG/f9Nib
B9locnBpMwOFHlJ+dwR/hCtd7Z3uiF8EouKLe4ZHKsOHUT9cMAqMpePlt2CE4ycO
F/v+O8CarNYF0FJBZ/vXJM8vfDYRNTx4OVu05gK3FfADvYfD2YbnvgqWZt+GL04L
8CANsLZwR3rvlo3dYkzyvvA9hiWRjdhNGijGnkWqsQH2UNifTc3WYRqf55QkEq9u
X1gjoayub7J/LkixvRwcTZ4XYgRfQFbd0Gd8yBnQCgECMkrC0Uhm3ovPETVz87QL
/ICM2M8Gr/y/B/HCnoCIzoWPqbupZ05IZbsXTU4HRrli/gVL9uz/mjOOj2M2vMF6
EHhgX9sGaDZytWWP74NTL5pqheNYWM0d+8+tTFNRQcjNAEPil9a9QQlO/7teXUKg
KYFjIzMwsM7d3gvAbxzNtL+etDWVpsRQFRUTnXk5T9eer42+IRdS9/U5l8mE+4QC
sSSZhRIgBB0KuPXItbfXGgvueDzAUPwEbetb6snMg3CQtS+2SYbtPIg/1lhPLjDC
Vx52S1/wX3DQdQR7yogJx/OwKFEH7CWinA5VstdZDfjpplPQ8w/zWAwGab5doMPa
eAKjjaFpxdqZQY8x0sF+znLoMor7IU/gQ7/OyaUk5UZrO9FMbYc/k6g6/iVEbX5h
qP1SsvWyJZe6pRbWLtHMRYU6Al48r0qE/DoPerbMIMTBtlmzIw/aitT/ryDwj1fY
m4G7yjJ8UMDRQZUqTJdeAlZEfawsKTQeH+XMxvuqmIUxjrm2YSWrS7n4vdgf58Pa
ScK+49C6z1ad9eBmOeSdzaTiwdjV0snwiUms+WooXmOW3tNGhvwidc6GCBLygJJb
v8wgMqCtP9ny08jryTuP9qYqtNvCinEHNGMEb/VgG47jCDIqzmfTpfHGJsVoiUYB
CdkLwo6wlZvua0+EvoeEl3XWwDDImrZ7YDvKYgEv0Lkphce/ofHyUJz977hHS/Wt
Gv1KQQLEo5FSkmdOLsDQFLYRV+LWZQBfvlddwnnxB+9GPMmy5gKejSloo8ExBvsy
q7aHcZruh05/LO9hWO0KKMiMa9qKSc5IkATcIzsNBaoosPPVxIm95Y3tj8+MdMtD
7l/c9o7JpP8lUCSzmKXiln1iE6uOJHDRgW5nyNYG5MWQo30iHyXFeGI4fPflbcPM
G6OKXLMDi/6N/bvGFa1MG7/ghAJeyaMi4SqAqH/yf1Td1dRIElA7xgDo+JH3Mvmi
uiXhRo2OnE6Un4bOHs2BOzC98pLJru0TtmVaSRNbk53J/wfsq5S0KFRsnZRjFTLH
k+Nz5q6BdVXnlHNokZlQWJG0ks/XF+NNIAR3pqmvk1bTqzqNU6srB+//WUbTPifW
rFqzC0N37lLoIMakoWmtQP48vdxbF+xaQ2GcrQnIOicto4OOdIvzhuQw0p8Yn+Gx
yVufQ4BQ41GLkbUeEaGEad+j9Ap6B1mjVjpVGtnDi5xRQ68Rnarstkz/7WP2qMZq
qHftqkEPWH/WKLQGoTXhXS0LmwAwiMirZpboskNgkMo3/2xDWLT3pp0+ofjHjkhz
lyYvRMfeJxJfV/1hZ53zJJDq2q6CfFNdXYL4dmP7eGa9uLG8j+9VFa+7XzAZwECq
KLY5YIcjGXfAP/U/Ypp1UwmkEscaE8EiV8XFnXrpsAQH7IXlL5LxxG2Kyxk8g88f
xmzKWcZSVvGJ2RhosDC/AR3FKc8t2FJoj3nCl9fiiYSwXWvWrLldahA1k5IwQncn
dckyYvbM3WDR1/rrzGO5zCT/TYywwjJiIzmVi2nBh54zYbZ1gdj6LCYLsMoJfbIy
RPrgu6tYiIqomV/X+w6ruSC5I6JhCVUxgDafgqpuvHwLme5F7nCH3bPX33YMuNmi
hP1GCr/WLgU+58M79Wnb2ZLiNJ0ngEZeYnXlfL3kCcZZW416drQahj1GD0Or08H5
4J76vCETRq69WhddEFCEYiVfOyQ/gztstJDcwHI0em09cDw+rkemGUki2N9U+ngk
xuiHED86bN0NV4XHjmZ0xvu8NxFfq0JaNhbXwR4AKuwKz59a1kjM3uh7OF911hc2
NxM9rXPNAn/2X+2+wRud+frORELU0qsYVYs7X3t5AIbqF2/w2Bz8LA3yCXZk0vf5
DlqBpCx5i7lhPBHB96P7R0oXPrclSQhcGmpik3yg3lu51niA14DAo820An22Ou8a
p539gyLkySC2FGOco3QKMpxEmBOpBKFaxfB3gwbfU/LtKYyc3ukyZ0rnyRBKvUEE
UP/de9yqnY+plteb3D9hxF33YY/pGNF5V4p4nTtT968bd0weZwaZppsnbmTOmFCz
9rQbjj27+ys94zw7PsNvqCRh/odQl7nljR4PHhc64B8mgpDxuXk9XZaz3LFcjLxc
yfEOkqC+aYheEiFD3+P9SymH/cvTnwLUTfpnt0M4rYHCmVZ6SfgSlFn/ROkCo4wB
/SFvdud38X53C9a6Tmg8V9tE8f0TIjq7gyiHRktrcJzqhwLO1TEdftvhVmkJikAn
LVGMPZZk5FwPI5ZaHH4DXQnB7PP347mGMniW854dzzjvGWwSvy732yVb9Limwyvg
TlQIndK0uyeJ7nkM1G5Ue30YNRS35oe9dHUCPbUWtaOVp0cGC41Sv/iXrhdGO5Cj
nZlzUTY0Q55qTzrU0wEqSqw2rZmfmh45Eg/+G2CjnqQ2Nq/A7E2X/vBTiHiR11/8
oRgvdIQrrO9X7dfSJRZJZYRtMLz92OTQwCSV5T5/zUEsSNQFliDSMq9LWOwaYoFM
kwISRbXns1bg9UbHn2zwozZMb3bYZvtIg/W1QODrghWwEEKAlFR/pqYIBdpbHMtU
ff9LufYYD+c4Nnrl5BdJi6EbQr5xwHqHmKaduGFVZqZEc3JGWDj6IUmS0zLzNlkR
U3dXr/g+HbfDFkMHIKBijkc6748hYPomvQSrY6QSZrvWSiSsnoijzLdwIfe1nrYG
qv1BdH1JFFZcF5IAgizmVHCPwEyhGBSd41faHJgD0KnLTHhrdoF4h+dN2MoHzxdx
z7d6Aeq4yrcon1UZTVJuBCR8bDsidbVxO+jvkuK3BNnT+SWt7n4VxqlKwxcvFXWL
tpsZq7zeYeG+5jmoubzL9cfP7Ph+GkOZXrBxz409zwML4Mzk8aBkZE9uT3Y8J2Bm
FGTji8nJ+fMfrvsAkzRqNbq9ZPEChrJaXb2TmSFnMTFS+PFxgwLpyIYMH1M0vS0a
3lbScQm9jZKcPzqD3EuOXIlA1pY7s0gNvRcWfH2zE9s4JCZXqy98trpip3SVkzUX
P4wM80Bv3b7BlIIYtat40F8Sq3OapfQw1eu7dd1Ko/A3KElEW4QW2p6dlr7dFP3N
KVI5UG3iecamu8gKWdp1WKyavItnU4T+uzknnwC2ryEgtyzl1GqiWopinEcNQ+yQ
2ml4FtAnXdupYbapd67trDF9HEPYtCcD8psKt2zvbSumUwRkP7o6NjpbYx4EL/Ks
QETw8xsSzfr3kQ1arECPDLiu5HNxYYWKC/cmoQLdXk0K/s+2xlJgu7mY6CNW7ui3
aXpbAsCoIr/xIxI+VCwjCMLhN72hUSr3u3PxAShOnoY+hS/HHGJdXgZH+raHuOwX
ZxaKmwbAC+8VfG9y2orSoJVPWRmHGUcQsBUyFivpQ+k3ZDyVwoXoXkEb0REGTMBy
v4fUJvMqScmcTGnmaSLE5SgAv5wFxENjpfjKQJaWrYmFYZvQ2qTFtcQYTggsVvaR
Y6Dt0xNMclfJXfWMcoA5ZhZGADC61jdAVrZMVcUBkNpSGp29rZBAuQ4vMfaJy6ao
utbRiqDJ9DmLGPP+4Me5tFhclb6uP6+WlK1wAuAP+dccijsClGwy5lwWAanAtumB
DBZJ1neHk7U6DTCdpN/TUb4PZyGJBYXUR/ZSIB4ckp6F4Yiti3xRBj8JOCo5IZg5
kei0Qe4Q935AyCpYZrL42+4x7UWKtNatnv01Tvs7ASY/NmYY7Q+iuGcN7/XsxGa5
9M0QNz62sSPnNNuN4eo05ZNEcpnMWu9HqHoIz6RMiOmTZPK0Q/8nB5ITvRs/H0TN
mg2Jdar85yI/5ppp4azJIgHuMvxCEh+X60GkljwZRY0tdh0e6gOy1pFo+O2uLxBa
pQ6g7g6rVMQCeiGbBgY+O/tdAn+A6ThN9F5riGszqj0igg4C2qtTp/0UEf7kpIwJ
jf7pCdqmEw+I5mi5prhCe3I/oPJS3WJr4ZGOGd+7U90iqikpAh8chDIom5k1HOla
fTYj1TXr7KkcEZAlMjWJISlVQVq9Y/PVzyUw8jpO2uV11fy82uDYFp6WEfXnqc1H
QFzOazJbaqN4p2Gpj/Eow/CYKMUEQ3o/MMH0/7fOAQ2lJoY/5tVTfjGnLrVcfGRn
UOHkD/NxOFladf7sTaPHnkA+jU3dxR1HQ0Tc+cc19HclIJ2szXxmtIHBRme8gn4C
qyvHLrAuoweI6108eBXhqj1XFv8bwjdsAR9xzTf9Q+fEmurePWSScjcF1p8XEv4I
WFqn847lzg9bwntV/6GNkyGxl0bjzm1hqiImFlsi+6jVRGPIU7kiocNs+mXZrr6v
s8kI7Spn8JyWyCweX6A2iiiSezmXS8JCatjKJDnx2I4hlTszTHjGijF7VHR2ul3j
TtjTogHXBIPjKgWy+pVSkpXEib427eQseypHsG7xT1n/T62MLoQWnJ9jWoZ1CYC9
/5zn9DIXSi3TFt6g7aSkx9UjGv62PemSGFaJmg96TiHlKc/RTbc3Vi8ziwFI88hO
NsXnu8JWnSfwzv/HWTZA5MEVW9zaVM8VUseSJTK6ppf0hC0kOn6/gGOocmgj30PB
17ilr015oX26B/7pH+TP0t/6dRcBWNu4nxHKDrHIjnj2BwPS2lS1oStNL88VOi4y
8nP0r90PfiT5hgL2GegYGciisw9kOF1MTbvJODZAsNVerdJmqZ6le+rOhALk12Uy
m4Rjz+1xio0sx/LNgNI0EKiF09AndvNL8GMWMrkUDPc8bTZITAfcSYDPkrUkwn8Q
tMkUOo6fJCiUXi+uHLrvqjC2KHHX1Dl5SStK+y4FwJ0iqxjSnS2MzXs1zHGtlV9K
inDiiGI+lLZUEHQQI4092PgUhA7VQATgZ9RHzCRvB5eg3+DWCYbIiNGRJirg0qVY
5FC1LMIh6puS+Akd/JfXA0p6XOVqfU2BE+vrabnF7nlKvyNn7iREG32Gu7skd+mo
Ppm+gmVscEuQuJJipQdmHCKh6bEqgNtNWCeNNBx9eGll0FKbCmldNPszPjtbRAKP
qvOrw0bsemv39a/Ao6ew3aKAahjxcQ+Y/d83MXbQE/5ctGMxYUDg2xLFUIC1M++D
/SKd3ythR3fpRWU+LAxZqdOKStvX5XAWfPaEd/HVTxHIp9p1U6/s7XJqYq10Y9Tn
lp9TA8tAiEBm6XeNR3VEsU63l0hy78ScLFL4IyBq8F9MZ1sWhjRXL+0UHTJm2z5Q
V8tba6FgyeynegrmNENCE6YIyZxIFmiQXsBqpX2OhbpUCq3tNwTcGYkzIXXYN+I1
8XHy6tPgsDIFSkCTk7sPxMMIzUrUn6HKFlcEYownOZZPHh0yDwABI1Ft0Dpdj4gr
IGgzyzqF+vnXDClOAuBNCp4n94URd/5janNj6TnIEQA8NSMVIVM3xIs8/EUgWxEF
I2boOZkkG/+rLOtTqf7p/OLwz8g01AgEzGShqTlx3E6tu+Ci9ZtkjAQ0u+E+pOVP
crz3wsgUTR8pMCgcsbGaaivZtz0mEC5mTuq9NURJ+WwWc9jxYIL6UQoGinFkeDEv
YmosqjNDkZbVcFhIsFONl1YufbmQjlIMPdRBF9Ex3bCf8+Tl2Jc1P28d+2HM0Wml
OZwB/1DOI83sE2u1GX8xSpRbu4HpmTkR7l4iovnpKj9cWb3b75tLtOQ8F1uUq3fL
VP464ESQ5t2a5uTBlHTX2+p5SedWh/Qs8uk912Wp7pVk3eSH/nYQP78hsl3c4PP4
v1+o44lvHhTPcmOoF5Wd9ls3lnGeGgGhrELSTE3H9B314A0y3vlkvVCbleNwcIC1
10rPwFLZgsLsTgs7WFRpXypT/593AQXQwxT53Z39DTjvooXbNs+DS3Y7mNCq2rJ+
3Z505a2/wFI2CAgZaRiN/wbOIo3S6Nu5/kuzmIjxVdcDTxt0BSGyu0LwG8OxRT6K
dUjXQRgFbRTTwhkDZ1OabnPm/89vtVt0g7wkzVidU2wIRCxMcgidt1/+sNR98Z0/
7nMZlgnxVGBXXpQzatSqTeYiHA0Mw1nn99VN2W9cpOUBzSQ9sI7F+8V7u6uI8S5q
cbTrQV19LVPve7QbjrDZARAr/gGjpWLiL+hX64LlHcHxtC+IDkenhv7rxQA3CeJD
hPrnreV2HJHU2iLL5kvshQh8ORo1i0asKbX2UejpwWPBCNmxA5YkuQTNiG0shngT
1jMFODelovLw37M5/p9DHlaILdIuUzXpFFkCjr3Jgkr24Sf9i0aU9oEjqMVjsHuw
Rb6sEK1W4yPIiOJKrLBia8bLcZKkYj48TvM9IJGnXTrISxBMgn7zeVEOOrATCeIE
O3gQzggV3zc3tQnChD8oWkNcz8FRX2/3q2qcZZcgGrwBqToUrT/+a8xfhBQjCEHL
N06vAB5C21BAuur87/7Q0nXQqTBmxeQ+uKqCagP7anS5qBEOjVD2nGXC+ugdBI1s
964P7LF0tzhcxlx1Rsqz2fxJpWxt3gsW3XEwep7cHeqPT/BTRlGrX88l5uIsRnhF
gU6YSl9tLJZfYY496L4kAagmM7vXlHVAiCeVLiRxoxSsCeQvXc5NY3nBwvKNwgnr
2/CdFq/zO/TY5+M1qjIYpGhHPxOE2Z4MW4KmBsWGKzri1tIMAoU5c6cX0pam4whi
9maLB2bilPxm2rV3KKFrNokAZsTG01hZ0sFuycdj0/U985gVGGAp1PvEBR/nsePI
w2KghaJqZdkI03YUJTY6+Y/zZVCpE0cIaCf8/e+YQQvuQaaKV9ZfFi026SstX7Mr
Gecbd0uV25jA1dQwyW6AZaBQhS6mKgCqUjl7NetdsoCzo5Np5gb1bA2efRw2enKq
WRX6jxNAUjhfH+3wQIGIyIPBJeyX0jO1LXd84nld8kzX9tzStCwz3b5H/Z/QWRPh
co89GZIljyfqw3nxgnbT5EghhNZ1FnWkpnvHv67SJd7HXe5dEv62SSg+pEZfb/fH
DaXtkhCQHt2ATpuzw4xXEcowCx5EWO5ASRXX3A1V5emxnJ4YPyKB3wrRS+HfjoZf
X29vJ8DgDs8k0hUc15NsBPnD3hpuKbOs2gWgvo4YXYBbDCRveCE2R/kmfmr3OIin
U9QvP/WbvYehmYnhzRJcySy66pQYwIYYHkYHP084JyZBe70vL2PxYWdyff08dfDG
wGEFnIvsYgn3/8Z/w+Pa5i0/W/Xvw4KATyfvJk2L/Zi/dTkjosMGtNTFhpH5Qawz
6zOIoSTm0kPOhnzJBqZkcRW6jTP0HnoCFMHbwWRZYGQoEgZS73+ihL6DWELX1cRS
GgNA6JmlwrhsdZTTlZGJQzw7PnMj/YigiJXAufLobCxLO2BJkWmyI8uPFcMektMH
T9KBT5QdSD1itD5df0/CSsSBH4j1giv/gtrkQNSzWZ9igHt8lwcA4ShI0nPVwP87
6aGEbP7WBqaKcsSAAy9cTdd0ctNlUI14vu0IfR1PxDVgxC8nOQFWcvZP7gKP9xI4
cFVoI4mlsVX4cPC7UiQf5jj86JWcahOWClk1pLnHLLw5fGr5Z2RaLNrOR0O5L5zf
g/iqV3762pMdbiT3GTOlk2XqEtZQvk72t3ausb9T5E8nmn9266uCREPykNn/q2+j
RvLocjbcJGO7BjVcnptJQHjt4SJDr5rU28AkR0aRU0W+VrwhqeVBTx7y97on1wht
PhFgvsKO7Qsh4O7TvmJ6ypeqattRR5+4eagxy2ySomL8IQdFMbsKlq7Un0yubAqb
6ueygpHUEvHoEJ8l6gFjn1eAuDWnA+RpLewL2hvVc84vIkj+jJgPHTRGYa5MGDpZ
7SqlK8YXIgf5+PRpOn/Vuw3EUXdNA1IjHLnvfr+PQgqBJhedI5kx2eOdTMolpghq
hn7Pu76ltrPZMb+K4akW5yqCMXQu5YXlIyiiK0xUz3kloED1boveau4W1edU7GVA
bH9yQq1hFV5zGrf1hEAY0cf6kX6BP0XH3Y2LuUguZWEMDIlIPtdHp/Au6shrNX5U
+14uhCIWwmI5IsgV/TgVAHGuU1uQxMMqR0MFPdC6Zdf3FV92qgb1jdsp4c4QweHx
WEKFyMltc7qKccyLDHLtBwtPFVJ6JKcfPDQNzju1HD/EZ4IMPLqMxp8NmkaIzE7G
QTtWQW8Wnsf7iMdBKGRD8edTI9DUSO4qgKZ/cFeLe/FMw0GLXApXA8doP3xRnJs7
JghlSC8uFTYTyRbvtDWt4s07YtXXYvbKbTU0Beo+ePzIOpMkd/oGFfhidQUT73OO
4JjuMH22xm4QTdUBhMRfkFzt0a06lsfP9g1pYteJAzCCw0ZOsLdRd+TvjnVj8+AH
vYwgfAGSJ6M5lV+6U2vFrRB/LovYXP6F5l1C9bLDsyTT4ma1NAG9pEG4hChHuM4h
MzV6BJsTJbHLqWIkXOWjblxRf6rDYIVDXwN/TU6MjwDIwEUCvr9h9IAvWEpElPqT
ray/oeI3nLjrPYPEf2YEDQLNJVlYy1WbJ+1tO724gBcbNbUBokEwihL6a66PJOZb
DjTsLyT/d28BeOjuPfamQ1QQXlGPr90dFlulYYWnpiJKEtWnymL+szVGIzWADJqj
cFc9wOIFzAbAd+xJANNHuvmv1nTOOs24llJQjCwUYM37u4FuiUXx/SWgqWnPrgy0
E7nD9K5VikfQKQwNecwPvzvQy/QITNHEW5ATpoQVNePk+4N3lN0qyZen6BIyIdPf
eArNuwIDFsMNEdLO2keykn7VY+EeF0aOdBpHxgbHUypwC1KO3z2+QLwlcAuh+ope
q+fSNxhvQyjec4S4Z+E5G5GuwFy6zDHTv72ukmAqGpmnur9pswZAKLbOyzfnlIU+
tlhEWvPJF82vIieH4vyIv9aIHxT3dCj/218TAVO678ZvqeLt1NMLTnCWe30h7Ol3
HDoy85NL9dT/5tBWsK8NJx50S3KkAfW/9p57nM12QYlanv6nguqAZ328C5iRTkyi
gwuYfXsWkw6Q96vSQZJW/z67MfpKKbrq7eaySh6I0u6atCdVAsFGLhg/HZ0B3dbU
gTIhshy0HMRvIlCb556R93WVU+bmH6iSCmJgFICXyLBMED+zqQXaKl8GGJCv4imX
OMfHC+OqvAh/iJ7fYcPKzmiE7S9hF+ttKB0O/mKuRzn8VEwGJoH17UNZ2UIzDlyo
Jt4Fyb3dQfriVBpTmmsjdzPJQTrlEuVM01i6e6Qy45gXjiDUBX8rIVhCahdFRz72
WAvHRU1D1yDoZbunYbq27IoxsR+hv6Zob1RBWq4JqdUwUsJbcZzJxUjL8Kew8sfR
lYhAVUuYVHRRCCJK93K1WLb9aa47OierawuIhzRXxl1R8FVBCQjM1YOp9IfExXQT
3cjJlFYuExW5x+BZtgqKPh97NOnGB68pPAqPxmBBPTkWNbHRX+ZiUzk73Vz9/pZq
gXYEZ45WL72tjDa+4wKGBs9z23ZvlE3ZsBZ8H8BoBGSDFiRLjhss+HvoH55QpdED
us2N2gyb3jYbNJPOUG0vgXz//u1Zajr4h6awM9R7TVNE358M6deFlBTZbSlvLX68
8vOZMvXM5x619HHH+TlZORyCvymoKif5SJFEB6IfZdtp2qsx/2ThUON78vRh4iMt
Rns5MLPImagxEJfTPzj/ABzsgNTrE8AY7bDq8VNeeKKHq98NonBaWadU8xj051yI
gNLK9z0FMfqPZ1uNthQk9X5hs2W+3qb+/aStyJIi94kF+u4gR3Rp2/mzPndHKOxO
En5Ei3zvjdkPn+5jHPHeVxa38nOaQrfGSnslSXVw2V/798XfRDKR6shP6pzv9aza
YRqacoP0FopiqRtA/KOQzVM25gjzw+sxV8nUnnXiBBExsQ1Z7Tu8T4wOy28vKneM
mwD2OxH0aKtWipZknDkI58jtUDr9nUBWTr0meABR70WX2UBNlc0p7WhFky/k2N/t
OnUTPEpXtULGYhKEXNo8UPpZdwxle9Y6vpK9FU/PEILxh/bkzQ9et2rtN4XdvW17
3Z/SzESpoiiE0Yfiqqbx88eSWCeOutmv9J0n2C20hhIqhrKWCyMqZVjqEZDQXzfJ
w5M6ABuDjA2vkM2G/lHsv8ejCw2ZyhTzLH80zeCN2YzRxWoabkU2f9zg8oDGcoba
bt2Ok99x+X0OAOsPwyVE05fslOtlUooyO38Necqw6r8JT/ZcEhRaXIXPgxmLyKhW
wpwGfuW2+QeryOG6SKolMEMFJYxK1kPPrJJXNbwbd2woMQHB0xq3rDpB50/LrAzA
NxvPNci/i1gfK/0C/JMnVGaYyX0tWjk4+hHjoVchpfwciJ3TRgUtQja05Gl1Hce5
200lSj5HsG6jJmFF88ZNmJDGUUHTTA4/tpVf+s6pL8+FkFxhacFRjAlJhrf2MaXt
ogl7EFpjCZAvYKZpwFJrIfMppNX+tm92bWdAF2REhaeE+cGN4F/OqzUgF0Gmvz5r
1dW68gGmtZn0XAqSI9p8Q8iRj9JfyAf9YbUKdpdBIx/DPfxWhPnd7izPiZthJNFC
uk6DZZKG3p24Y7VCiDniz/wBzaxHBKjUJQIOqXXLGVmw5WXA0+W3oG/kqmI/KIJq
5BaNK6aYz15CsmWV/6C/oDnFWFkE3h4OcY6PP6/Ddrsj5606TyroGzGgJ9WyAAp6
WrFDjDjpselfU9JR6kkRLkycWFI4WdtHfao26SknsxObuEN5FfZ6kpGtyNG8AAyf
RacLVVAQ+lmSwsAra8zNOy3CqdkUkijkzG5YZTApVJl8esLh6h8ygyqgQPz1YKzb
iqDJmjmz7uTIcIPosQVRrbnV5j4+yobtTdzQ2sVh8tZUpYU9Do2QUjtzXQqI5thp
2vhePEEdNdnbVr2ZoAkuK1gB4UjjoT5lPJ7h3WPG4XzYUtmnMZDRyHe/DVVEEP7g
TUfCqgMo44p/qH+gdvJXAd8hIypyLrtVmdcMryZoNrsxAMS/8e72MhG9ZH7iU9QQ
rujS/EtTmjFgtmqOde8udg2aQV+ZBmT6Mf/k09x5PgrA+cZq4brBivOf6E/RvHqP
VhBdpKRAwYeKyxR08drAfBGhsOMpSOKj9OOW3J4A59R2WLGRMxbLFbpBeVwOWldv
os32DaOK7qFArX2Gk5gQK+5LPk03T27zdRAouZp4RyXTdM0puJ+fbbyC8JDPrVbX
fcNK0BMiAEVZ9NzIZBh5xjFph6T7HXjAN4OlKwS0q0GNEJ98l9cRYKp0UJfgOtVT
PsAEZ+BMONCWJYQqNOWum7SOgKtSzFOqP1W/sOznbm4atTjyNpZWpAIcBINfrfkq
8EuT4YZIwfbJ9XD4SSXSaoxnfoLa6h2am5q8VJU1nc5SSS7RHCkgPgUDqBDjTYTw
Vr1CL1bGnDtBOs/VlnxUMQu8IsTIJtAuhBgwo0WJ8fJ85BO9sJhkX/n+PpEXKWZz
uMSn5RrxX/CLORUZUH7KDCO5TMFwMn2H7T7frsLTaRZYLOeJpmQ28xctvz1eaSAG
EAN9DjYO0iHFqCeESqrBRsW6h1yqrKqDEDuts09JHaEtxYxkHSKDZFRcCYzG2zRl
nRAk6RCT/awEawZ5Z2eAxI8ZyvCx2KqAnQqXRUQdk9tSjemvq/M5jzkKO/a89Wmi
e1iIqGUKB673kY3UQ5Dyqv+ntwCE5fGv6nqz4G5e1Q0TohterAdVQv5cTaRfPb9M
FyZoeQ0URhAZyor0QT79tR33/rJMM+3Z9nSFx3NOXM/Dms3pMuYccsHg9Mj9FyNW
moH491nu0IZ11xof95EXBIc7t/1Zr22Lx0Vy+C+dWCi01CifF9cY2PfugkV3+ddY
ll6o2fm31GiC7dvPcJF7NJMGLe272MD/pmXZUICJuF9bVZWX87CdnDYTASJtCJva
vREOryEs/8CWnyMVQfRotegXRtegSXlsyS/Ra0FUWigGQBNb41FfX5JVfVVV2jn8
gRLtgY9X844AH1qwWmEMqEUSGMJp4hqppsWOpcRttQBgK/M9aoFu+Jau6Xix4uwT
2BsPL9Zklep6rFcUR274l2diWeeqjW8iAiCbLytoDyUpX1Cy57Wn3yGxmBmZaBy5
eA9Ei/IS6G3L8PBmFyyfcmrFVx2SOklLmnI+KfH6nkgsTJ+mBomJd0qaM1LtHjbs
WpLZAobhF13K0LNyclM8KL2gvSadeMsJNk589V+YEVXzOU1GVdYC4MtrGy5Aekxt
ID2xg/lmTAi1oZBrdjgbuD3XGnHYh3ivCf+z5IzVcHRsOqEtDbS7bniLIfbv39lO
CNh9QU+0JR0gSzhaB/yRgGD2slpCzxHRutsd2ddoTgVoMzuoszbgiTmFM9t6uz+e
ZX85zwP+uJ70ey7XSC4EjRAx1aX9gW9q3uE2EMHk2jslGuA5Ac4Gm/w1F1pLjRwZ
VkQGr2SJb0mdjAQg0s9yseDs4af6tGJ9FLIhm4nMsf3z578vv0PDf2KcPCLf6A6f
1E8yPD/IJGWqoJjTzQ4pvjVDGqVp4d+o36SJoK95GSMu4F1iySb3x2YRT8U45+DW
QZlygOSF4suNFMFKG+EbA8paMNT94d48hXVAshnuX3XinQH+Zw6cGxG6NK23ueCx
JQP8Q7EINMRtbVoKgcalfC4B0M0aQ5WpreXvIA1fxhQfmJsp9Oc7094IhBVw6EUf
b5OM7qhVVrK93knh4ydyODzko/K5Os8wCERqL2Y1v4cNhpVuBt8UMhMeqm0+lkK2
cDlVRY7W4Qml2kP7YulgS9nB5qbaMp112GcMewt/J1HbOOYOj4bMPWfLIwzjWNL7
1Cs/My2EKA79YI4lKxhAJvN8kBTsPgxyD6m1radRElJJ/ouiIpqv1TYiXZKz0gKm
lfTAMOA9KBhheZiI8Oy+9xooeAEvwUs+Oq9S7in0UIGte7JF5BAUD6b4qbLwAsGs
2UnJFnly6iLEusppKLwrElOUoMaiNeQW6nOyykm9icNPan7vs+gxl7RxPyu8QnNc
vAOHIwmdf4yvtkBQm8d+1GLVAUOedAmySxYdLu/k3re8qxs3xooaln2Q+Y9gAC49
Yew0G9u54ByrcuV8+SqER0V3T+vFqq2yquP/0YAJYMUqUSxwsBoOEGikDCwqVTgy
xWQuIXDAeHxnRpulX1sfJcnQkwpCc6n6B0N6jtJrGysREY+pi5+j2irmXx3+yHiR
+F4FDeiESzSxmjudGJ3HC0g2Vk3LUkmEMD2tRd37vT8a8KeeeMaCEYf1XYGXtfbS
CSbg3dj9b3jq4i2I3ufYpLQje//EjA6eHDGS7uIomDEN6wxrrUnQ5rQyQihxboly
o7zQ0OxUzsyPU2XQMCoFS7UQLMOr0FcaBGaMbNIu8Zw+F7/vBKmuBOnOOBqw3d4w
ryP7+8kc+XLVdG/9ZaxQ+amVsrkIHgk9m2r03gPdzb1HlsbyGJVHC4LsYvUELOHA
Wp+S7b8WgLkxTUVOMWmQsn9LtevmVPZxbNN793ujROSv5Q4dnajB1ZiywsjvBa3F
QziuLb3WeBSWltA0K+MI9VGAZ0iHZx/MnCS4peARtqvM3Ouc6w0U+kQjkSUoUOhV
d2BebUYhZ58dNVggH7eNosVIWWIntB9zaTLytdyUKrp2eoC3+cjvkvKmk0XRSiAS
6KeZjhO2BpUbHcr6ofMaN/2P5HBp2X+veX0JVBUq9CU0Lgex10ctIE4aGQbbITus
M3du5PrNUZND7oQDXoPI+94rGJ5t2IMIzfmm3YSEN+HI5KY0z2Wct1c9ZKHnfNPp
RznjoAG57BmaAQsn56J4EvFqYd6ND6piFCSv6Zhwo4Co4wIknGCqiQEJXOPaR4V2
9ehDjuRoa/LSNpiQcu5NqJuslPeyKxPZYg3qCP0W8vvaU9Cj9/s6GKjWmRCdAifE
0zWgbhSTDTEuMquBvd5NnA2pp/EPrSRKxSt3U4+mJilCYZRPJH1wAIDFRZhuuf4G
1POghw276NOJX9DL9gckydpTMCvsOrrUsfZXjpxC1YGLmVVtC3v7HVsJHegttZrB
K2eMYOkdaVFX9CXA+5Akwt7RfXnYwa3buaY3wDJDCjmN3rNp/XGhDkPKD/4X0ecp
Ahfep8mSF+ECtTSD8B+sQCPY2rk4YR9Dpo5cD2iAq9eCuo8aZdp+ev3PW2QsRgdc
hv6Zt+7TkLXaH8MK91uIBBqU08GKzzFU915UNEq5UaLyvUW39cdc8let1gRVgeUN
QhYcknnw7aIhP2kdU9l4zXwnaFhnqLkhxGYJ4Gmhp/TZ6MdMTS/Mh+O+5lBwvqHa
w9o9idHmaDtS76+oKYYXQvk1y1jydY/9TNVXKIiYKqAY3X4bBPF4GBG8LX3TjQDe
+Op0KGjuzSrqwrw1MLml7GxWmDYTDPL4pEgJjCDUdfSfc4lT8Qi6pWZ2WlKn+mgD
b08iaDyXJw2HDg/sl7lVtmQ1wEsllmpgfUl63dukLsCAEgKJ58fQ2LaZ5UPur4zN
xzkhH55JtSHgKLcUTkDu0Q3/mgbW3dU+LWUJ9mA3CldLRz0ozdcpqnTODNwv2Kl4
lMEfISFiCScfJHwuhd4q943yIsq2gFgq5OZQciqF9+DUJGjudImkWSIzCjCRI3+c
cJzjUSvLrsFO4hUDMuyUY7AWIB+Rww4uRA47aTfKmrAaHraC0HjGn/icPg1zSG2b
jMeQqtez94p8b922UFYnXAq1h8/ELN0kCbZlzCJ6LpenKrJZT/xeGs1v1FZ7VwCc
gCS7Ko1ntf7iw3eI+o2R2V1euEo25z2zhzkioJeiqtscVR9dttkcwi0/4Q75XJCZ
/xlIL2aPPnWOhey/WIvghhAMq+/hDNiuQic6YiaQpDj4Nve0CrZGNWqq82jAB8lF
Vdwp6riW8Z0XnwKgdjHRoeUZFOzkU+HoSQFZqq/3B+h5BnVv2UYDCng4eJXcRZM1
41jJ+nXRMBxQ3HQlraIOQPEJ64FekORcbzuf4lpt/GMAN4os+w7tyyPHiQveFbnd
/IdFaHlIBgq+LpmtzE4/CkpMty99wvn/Qim9WxV8+/rRrwqUt5EppSt1NnobFLdw
6NQxGx+qz3n9HuZ5V/QWg3Q8HGgNH2X2WZvzENB0Si2x1af4CRG4vxzEcXtuWCMM
`protect END_PROTECTED
