`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B3ikc046qnRb7uTamthweFr5VO+S5dZyXzSwjrzpU4lFCwEcEDrYUhWvCebAg74z
Bi3WfULYJNMX8npeJ4DtpSt4bzP+Z1SBEMtWLh7XDO5e7t7QMIb6ztFc6HuNrmIq
4IYwHcG0yZe/u+rAUy1yfraK/lPHWz5WZHRB7RjCJYIUVmsJvLJnPIymgPzmtLSf
rgrbuHEcieR38SqxpB63AQogR7M1bevGSO/dvHaYCqP8Zqkq3afPT2UyPwug8x3d
bJ/iNbtmFJW82YbRaPTuR26/m6Dgwmk7r6N3cCq+oZ+mHSrESYp9in44rNkkwEUw
Wud/9RoeWRgyr2+DdsTrfVds5BbQzbxKXHubYc7+fOvt/QMC5SSoahELcPwg9lQW
RTEuTxC9DamtTQP+7suOJNhDXd5uBw66ZepXnJ9Ur9byydxtQ1uz7mS9+Bp4Az61
8TIZKFm+imM1kwPA1SP/HRQ3d+gigDq764NMUakCV3Hz/nrrIy0B9iwq6QKNb0j8
FB94ivZUOcKm9mv7DFFAfW4QhUY3L+ry1cyhulVp1qJEWWKt6+SycrL1A2imz1AF
nXwAn+WQ8hIWbS8Q+e73MIy0FVbRax9G0OrFH5WAuxQQgZ1VE/VLAOOhT7livFdV
44keXCpo90gB87ym0X0cQx5eUTc6Qhq/cuwIN9l1BJDQ0pEMTJsuSLKkuBZ+apAd
f/UyI8HDUf9/2Gg+LaSMLWuTC1nZfULR/JBJbX2H4xU=
`protect END_PROTECTED
