`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s0PoleEND7sgcTJwGhTBc/AE8Sm3dsgJ4YmUdlC5AueMpaDcBs1a6WAZA64GS+Rw
JZ9BFufMPOjuCxeAds0qvr/TZlvVnIGOWeJnVBJZc8cdpYqqB6cfecJWE5tqmJox
aisgvFF0Skp6rHOJMvum6qvLjc8yGdhfg2nG0djkKtdCH+CcLAWBjuhwLuFLish0
pGXZrHUYwNagOxfQb6HsI7JBahMTag0XD3J4/b+8QvpQH7i7u5RALqPWT/1q6br0
SdnUBGxJZsO9OVDiCtPn/KPAbbWiDvuF7Ucs241OEmrqWEjVFGGpMaOL1WPNgaff
JMq8cDhBDuoZkFA5ciYmUZxezsoNimJK3RURZ8yfdRYwiK/jzPpRnMXNDAIH76Ok
E4tVwatiFXutf5PtqZE6Sl10jzsA5U624Xb2Rv2RlzfhFV0elckYmF3WVJuskoNb
44BWE2ubqmRvi7e4Ex+x2LXn95NfJUdS4J/66FbJPV/b5HkV3/CUQth03NuX7xD9
snXLOVdZrmwP6hch8xshkqeezsDd16PRjFOJDUPE3EvCMAIG/WPR5w/3b64syQZt
VqOnNeLGnbnSk7Hc+qe5+vylR5CChmNvte/GuqyaX/TrQLVp74zVuoZu4pY+9iNT
WRLNedhkhTjoS/YotlrcoKD1u0ZZcue8UI+WN+p6vUG3BKCjwDOBOF/y8RXL6Ozj
2tk/s/2k0mTzidsdkcM/wxXgi2Z+8UuJFrdsQ7Bc4DVCsTVaW1ZbGbvgFlhWqN1e
CxB+i1g0DgoHauoC4OJmeQ==
`protect END_PROTECTED
