`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQkU6fJSq+1iMYCOGKR+bE98E1+8vd6q96ae+YoPiJR5Bk/HY28XvzMfYMB+STcj
Ye9tXS8Q4RkUS1a298Jp1yXfVe4AcuwEYM/R82mv3sKdF28tQOnwJDaYt0pWig21
CzrbChrxr04aLaUyyVnx5TgMHdhyDPvL6xWnPFYjawU+nT4/TQmr0Mr0mt5pE41w
P/Scc/YoStOZqf6LCXGdWfVZgop02plI/XQI3hRGNyGtEWXBaxgZfFn1k3EUxB+q
4r8rhItY61Mxl+xjlcYBb+3c1NeCRsSl/yqteyAPkHmFdIS71QujWaJ5qhiignwK
a2HaIEXJE1T/s+k7YJ99O7llu+PLsxcJ9qGzBybUsbBpG3o72T4ZY0ar7Ri7Uqra
bZwM0ZK8sm47pH3g160+zvZoKpvECV1+38zmnTmXkfY=
`protect END_PROTECTED
