`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jr1mM9R7cDM10JbEruB2LXx7UxOOwhtkhUcH4wfdM8pq/1KOBVhUTDhMvZB1VsTF
/+0KgPrY/tu5+P84meioIkBSMzc3DW/LmccgOnh949BBNL+HhNI9MTtKGDUWunUu
aHlfYOk5T2EXILkYTKKROvOChLt6BbSUOOAlOjV0EC+L1SSKTJJ2+5A8GltdyZr4
Eombh4etKkaDS/zXYZZBOyBnzKqi2az9A/AobFlhBWtXXaIQfa3yM5FD0hlg5Htw
WhMY15LM0HRX905hrZ2fRisB58N+Oz8JTKjsiT+AYa0JN3h9vBB8DmDgt1BRPaSS
Mx4FePi9UR+yb8q8bz6/TCnYBY1Mb4D7MdWTA8pq1hL0kJMb/mxzBO8TzfkLNT9i
SJrkMM8DqfjsJFbVO53CmmH2j2lGl41YpJ96MyVlkMVLgsld2oQx+G3dd0/a4sXh
CctNzyDM+iW5ucb6p+L+YgcQ4BcMS5LYHh42cQLe8Ti0924ny5HWJJ8wcmEY+hjC
rlFJliPA10eYuovaF1/2Q3ojbdGm4Yr0pyqR+5kaXjJn9YT4RzZVaeMJefr7dr87
`protect END_PROTECTED
