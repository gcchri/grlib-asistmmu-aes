`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXatDRvWD5J27u93sDptfdIl2tDrCtcYyGrQc91axH5B0W2YDnAD4bP1oQztaiVM
6b3C5K2PFHYtJ46kATGqqXoUO+X/vSKx6blZGnnBZBVnNY8hJMPercq2izz8izNu
ot6Vj03AXMcpkFVQmMl6KG8lSK8vg5HvJakahxGi72rWM1KM+QquthnTGZh9JQS2
KiPXR+4h0K2c3FBHbCxzYvkMkVLvnpFoHgkm8TDDjZPgLB8OHJ3SxtKlyfd9zlZa
CqfnGbPYWRnS6iU1u+rGRsOHtCGWs2l0yYWunMw3c3XctxlmIRA7BYgX9tIEZ8QP
HIYWq3UhNXZ0ImlbHdfzbJAC+Rs/z89xYU4GX3YvvicWXkPTlviuxoD8NW0FDqSb
AnF2q2F8aL4rOQT02SBI9i5zN4RupAIWEIhlvluHK5BYtXBaADO3hHdbWbaG84MP
0wSDUI9WfPAykqyQs2qKxWytnGNUDHxsgi9NfoaHA/hdlZlI9eQz74VqCnBuu0+T
Kfb2diux9laAgrNtjSvpMIp8SHE6qKHFCOhzgmEErYKEUkRjl778o9+MCzZ7ynGs
Kq8ZgyxOnrvCEGIQSMJ1yaeZqSFfxy+6Rpzgd8WvWI46FmjIet+bOvI35xlLnC5w
DwDCj5oEyxpmbwLxRn3UwdFsNneSUy4gCSAHNhbFbz16SiADV2abE2vW/hacAHnF
25+XWQwSxUSU7GsDu8EHEDyLYPjPQ5Kd6R0I9aWB1IcIzL0wlnHxMxU61Kp2lzBA
WD41AaSq/LcaHnNiSm3k2fQWlutgmMu7Z55IqbEeWVSUb51MjamzbADm68SRYZEI
kyxV7N7EXxmvDqGulloMKaw9YWC72LYO5V7dJdFH9DD61z/SBOdf/YhYzQx0NPAE
RXys/c27OyroDVbgN10CkJvZbXVvK7pMPF+zuI6evQE=
`protect END_PROTECTED
