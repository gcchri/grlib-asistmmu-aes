`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
If6ZCE+P4uFz0vjCXlTkrOiJV5Apm+jWEvoMWAEruioYkpve+/I7lg1PUw+ELzBo
4G5n5E4T1nlP66SqE9jNPEiq2D1JqBaoj5CkaXR1jDkeN4Rhae0ZluKzfJCCvq6K
TaoXWCKmV8FVDrpQnxXxFxnjhkrhig2FANUqes9sb3OJEIyLVpagHZk3vZ6VcfJn
QAXWCi2xS6ZrHp85Mqnzp0/MRzCcIUS71/pgeRFzET7AKt6YV1MS6oYtfr3OFFa5
mc9jLUMZf1j3IL5tv1flSWupILGsyci7ZDmn5nKDOHxyuRwgXKV3uFNLlzI9YLHR
dfJ9jDpnQORQERGxf0tbB8PwJeC1GMwF309VW5ZSL0lJUOnr6M1m3QJmyAjfLJts
RTMhcozMfiXK2dZ/z4+MdZitP90OD2NphLevzNsvdltf93yrwpvukvpPVPMHN/m9
7QtU4j64sR56yx69ile/YLrizNa7a5dmBMtVFSRJMUIa6BuXTwGwKHn9f6YUojp8
jn7XJrTuxs7nsiqX0NLFefmAfbH5a72JSSGySYJ6ZADcRwJU7rtc2JmhIIWs6SOL
qUhDGtFgGnNOPQrnwkLeWikQAi5SR8XOl+rrcYx3DyssSIwdg44lvhwDPOeDS7I9
UoHd3h69OQFqS6wRs5eBvQ==
`protect END_PROTECTED
