`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/NpymZuat82N+25D8DMBP0+vR90i4TTfQK5Ktc3e0liovGUkYndUDVqqP4qIx/GT
P89nUNH8vdsFmEHtCtr3uXJY6LJigzb8JbPNnPKrMMOn+NkWPTy8Hc/VrqSbo8S7
0nO5trtwADS/UdTT/6MayvEcZzeBnZ/3acQcx0zBYBqlgfEepvlrYdX4uamtxx0Z
FeRlco0VBfWZ6fDwzAUmcjiOhd28gSOMUdFuQbde4SKdbqqEQh/NJhXw+7pxOXjk
gygKCl1Xf4EsfA5aYBT8QQfLg7n/nHOlFF6Yom+0DnTyeqH4PJwtYoiKyzRf4p1H
jQxZCvr2iSbsMAkPmuYXZLBGWiA8wWW5XDBVrpmB0vXL8W7YG1tW9AExtsK02wPO
KzfLRlORwOGwNG+VMai68YjzrzPBdRRgjfWlUKV20C2mZZFS4bnhpGnjFW0stMpw
ccROYUcyrf9hzYbCeZfbfVp1VnaDoZwSri2or7zl603kBZIpv5Q6CKR20VbkaX4Y
EaZOZGzd5F5X019SAWx8y5YsaY72S4RIc29i+YJqPZUoQQMcGxPOCHvXcOK47PB0
1X24gBK8rQKZdOJfjpdz2Dm585+Hfu3oLjQWMAA0+d1/ZRH+/PekwDlPWgiMVJuk
BiYuYmd+b50pqPo5EsGUJDSykXwKkwmlulgE5K4XMiYU2rvjsF8nbLUY96v2K2b8
ASggay+fASC6xM2/Y1z8gZ3tUX88bQV/9MNPIBLN7s5hsanfagNAkXczvUvpwAH1
50jFhbhr6QaKoc3uk29Xx8EB87AcJ6Zvm5L+NX6lKMPV+gUpnrcVKZBoB6X4+y2e
9D3SAOmYRgZPrTRF1neSAOZZ8zUIKTq8Ue7j7s5CtjTugVPpFSLkwhThCpPyoNz5
CMvQhG8yZxv8Zh5tHc79Oowrh0HqqPYgcwwH+TujZkqCX3bnty+gRcSl/d6RBh2w
i7z41S7qbNgL2a4LMHvvxE261IfmexYh81BjGUeivpgZT4DHFy8x8nQzg81+p9Sx
bnQE3mgfe+/WuTWnCBIGGEQmElZpKagLbIixBFTqvSz+Uo3Psh7lrwjA+aeZ+jLC
Iov+SAydP976AYTB4LRcS6TUr4UmX5WlrJKa3XySfaX+T8Lfn0J1Sae6yOLpi8P+
xqCOv5ArNv27jpiLN3s9HLjftmhenP0yemTZUso4/U/b8pi8rHicp+unu7hlYFGk
j4BxQovhouoER048Z9eovZHXX/Nu+g6XlEb7cEfoSX2iZgICeRo0LOOpyG+/0Fw0
GhAcbrnY5HRnl0CKA5+uhs6xKnLH8eg6Z3/HfyeFNJcvdmj16vjVE/93Hp+Smgy1
bB1DvpxxmZfqXItm3wgZD1aho4CoANrYZU29h6DHe5ZTp5efc5nCb461cF8CdRRJ
qYpbpHoSEKrkWwrqPpu8lhh1W3++Jtek8cQfYKeUQ7pcoAQjAZncwBUUFduzcTn9
1rYYXkpaCAB/RrpHwnIlVtm+aVI/iqBu6FrYcY0CaraFXXUJYBjiTGkDsPT3RuhB
XpdTq8caFCc0gPjQVh1FjgmckMNFQx9HAElsFrcXJnv4OoHbwJua4Hl1rky6ZKtK
WuEVnNTeRAZqbFwUlje3/Ka6Go3jdTaatoS4QPBeSOfxDMUCwTB7WLeW0lR3FKO4
42ql804Gkwe9radIRCcSerM2433x6+HxQa3KUVjGKh7ZUEiJHhNJT6HI4c/C4u4W
9+PilkZ19AlLME9itTiAZtzJjE0qk7qUlDnYxTdVSs4vbKPKIDOwO4Ui5wuZ8Hcv
reocfI1Fl84etKLBH/vUGFoWL8DE4mDY7v1vJXtek6gSTgpAmQc7KDBsCxt33U7v
/u5iCbOBF3T4Ej5mZdlQcdRBQBG+kVCaRnS89OIiudLetXXaDV1JAJeg5M6xPQvq
wQV7ngzUL2ez+Q1p5yliCzYwzgE7TBT6dG9zGqiIpImeTY3k4H5wr/DsXq1oEG2q
pIQ85i5qWw8BiZt/YzJ58q4bvGaN3zGKaCxrFTG3TsTk8hlDY9dyjau29F3oxMpd
gNeNOmHtELnhp7qa4VbrvLNvNAXmnf3wBDwwQgBDJuz0QJvLgde4Nx1nTvM2JGvc
YHcDl6vkNm9yxtmqLKxyETEyVEiDOf7Z4PqXnSXf5/7wI/hR2sPDsn0upYiiDsQM
5ujimd5oyrZcRnBkmH6eUnRg1jBo/O71Cd6GCDcbV7twqLxWLnaNwOZszH5+j5is
RL8/3PTHOD2B817mXzXLNWZ2cpJyUoIJWCz3yx6AUJhhCdGEn1FgFC31lInMXOI8
`protect END_PROTECTED
