`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMNj/gX1fwOuGInH68KyjQMlc/9Ki+U3C4DIztwS1ojIoLIm0MaetiZTjdRge72S
LrJVnTUMxIHb/6U6h239jyLOfwTUSO6TBRYwaWjZDTCeJOu/C2HCmn2lUebJdgTL
ekju1lcKjkU62GsiyJ9iAq0EghnTHvcuNFo8nypSsGbEFKG/cQnvzhcQF0GdSSOx
jHGZcYiIEykRVo1Aj4y0ODdQRcY/fm8D2Y7yVVm39alH+e/imozZXc47rlfMJJDP
N/eBpDkCYqxf6yR2zi6EZr4mHL9CwwfyFePqeDbcUHQ1DOFYs9oVkkFO2FesX5y9
RTNhX1E8QdVx97uAJcHgHfp4AoWsii225j4aB6iJSsk8mmNxFgg5kWuNym4EW+p0
6M6pk1fE1IALaJcWNL4EhB4ew6qTLrmorqHUAnyHTq38XZLRSgfkGJwBPayM0Ccj
T29efPcw/UBmYLlMkT6JiCMQGbhom+eOwPUfbf4YzXKVf+rSB56zeuiOETp0q3NM
s6hKGTspMLILTKHRaCRLQQ==
`protect END_PROTECTED
