`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQP1bVjN9noSlS/SrjYRa+uQ6b0bz2Lg8UpJHRF7dizHvIEUrv2LhKkPFD10T9B5
9IgrAgddfPn8LcuuAFAyv+twm4DnX5eAuIgPR3LKBC8ajDnUH6XrN7Cj6s/J8McN
hXdsG7gca0rgkOpyzKHM75Od8pYJ7HTILsQZiY0qFigDEYi7alKWqSRCI/N+jBsr
qxrKuBssa3gFSBKNYgj+I5I5kwfgWxFKmO06ryKRK1avc8frpm8AyGzK07SUiChf
am2Sf+7CDn0E4mSFu6O1q+yY8Z0Gce7K37S1DPJ74QNCiizU1z0qI1v5UHYe8XN9
qzV1zOszkxtoLpVssbExyo55oDBfuRff23XY6KxXbZCl2yI02lN3mjd2J8OCVWv8
q+DIV+lUK9hBn+P3f8Wf3dPl6pC+ZK8NEqhe1LUOWz5NCPDDASK7t6d05R7vUdHQ
Ev1pmWofhxME0vxvW/4ie81NqcLoK6USUyu1gxhLm9ASFDJ3TT3JbNY2O7mM5RpC
yyPqN1ndd0l5YiGVaLwWakvln8kY+LYJ1+k+arXjZLbKWbux5TdvHjaMd4tmjBES
r0BA0rs7YeZZPsZLfWtaof1LewODAtqGjD5Kx3Np0M7xOGbbwmbJ8dXK5uh1u3mT
V155ehytsfD118w83+UeQGxl4Z+e8ehfValAWXlPVgCBVW4RKKAX2ZmcVkn07oeP
Q25Fh7EvS0POZSpvCUpBFd7LTyQb+vmc7F+k8qDpUlDc/ScUEfsA892F1LpJFPCR
rpfKDr//7xx7gD4jSJOZzXuguH3gSSvwvBPwGs3+CKY=
`protect END_PROTECTED
