`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXWPNxG/qvoSkvZkuBs/KjAAro3OuKxSoLHJK6b+cFiyH61u/p5NCuqzbHs1o3QA
TpMxmPsxq8iGJZy+W64gdUWUktJsxx1x4L4gcbr10Va/gfFN2FTETkw/F8zWqXa0
bASpl1NKitwPxSAEGjl96NE8GdTB7SdL+Y9umL1ADPd7voEJXQZTsr/fKgeIfGvA
LiTIlhSnYu9LoBSAOLD3wJkTAN1gnWtr9gF11cgRGPyZRx4Per6wBQG/C0jugF2r
bIqiikr8VzwxaP3Cw0hXglIuxgI2wj/OahCFYDPXLT2q9lvT2x1K9dzAFpXoiQGk
4quLmjbnDshg2A9ZYEue194jbeCkF8O6GEIAXVWMb1f3b+Ru1MpMVoxMDAuz4cK4
UtP4STqeYRSiaUe5ROV5uacdfkbJU2UQxfAnh/yVftlw0S/g5mI1Lld140EgeYsm
33MfLQeXwIIszFrwQmw6UstG/rh/aqArkUfGCTXZHVuDDIN8PIAa0WWFwb3nHApt
Rt+Vf4Fyv58TiVBtmvFSGI+6rjZRJ2u9rTbzUeShxTK/xJH/qnxOGwpR3Q39BqyE
oNVh07GbwqDThC4OM5IgZ6xzOK40UDj/ZdQEwdHUhin59hQRI+6WlCFhCBNy3P+3
Fz/BlY7jT6fjLQQu8zYGJ7IcPaCBofjD1WXFrEu5aNHiEdGh5ha/8HU/MO2/GnKP
kuDV5sNviwNhQVA2tRZ1HsI9Xfz1n+nqkYX+H1C7gGMFwqOpiLUc14u7RHPi7yOp
vhFsFj51201kvRBDFm8JQvIP/gNfnNs+qr0oZFn54wzWn+xUOvxR+HNV3Ql3FoaP
lURZW3oLgzv8o/HZgUunD8gEOz8mgWkIcQUY3GNqTuL8AXp8XbcO/WlIn1luUMNr
0LbAuCgjRQePSRe+y51AxRQKMWxN6BJL7xN7M3GPuVtReL7LZpHwneiNnjhXjNrz
oy4ecmLBEp97YlXNOHKl1J4s8+5HBkC3+fG2mYjAkT41osPQ+a0Q6lwkZxhsqyey
lExhRugEhrhZf0riDva058PjzR7Nr1mHXk62Mz6vCFINb4rh0yfXuwwmFhHINH3g
T+hhh6h0AamEz+sVOle+GZiZk3MG0j4q05tVbdYDTE69a8YHyUW2LJPauxtXvoX9
7WFUnBLs+nYas+46qrrOjgWfp1WwIHv5cGG5lRFEhPjCP+eNeuWjgcp/rLaT4TGe
itHwvYmfVUASthDh9dpjBrsMOb4VXMKDZlT5pcUrsm7w/H5wJx2VG3LWpRY4NSUr
2JeqM0wYkktG583B57kRzKCCv/Cv5k3I4BO08Qw0SH3TfxHclgkBQCw2tTRSBmA0
4+npXPlSJy//Yc4gC4BSA+lIPfejdHDE0E6T5iazLtn3xk8wHLySP8pklOgc5WEK
XGgAGM4O4bfs5AuLB7NuKPS98dHmySUqzXEPtniRhBSNI2mYx5KDiGwPoK7Bk7cu
0JfBNIFi1ZICby9y+IRNHuAqxYMnsX7Ei3/G0NmU0cOv/HkoTnQb1IC7QtA0u8yX
kkzZW91+baOc8QO4m7oBq4/KKNsJAXP5NBGguhuuAiVAaj7UiUel7TWWq0ImZqVf
RBHBnwZheTO8uPp/zwxHCXYwf0X3opERBiF/GISlG66/OjPbGFrq9u7+BJKOpxL7
gMvcV1/myeITpCMzr6TnCcX1QOoFpDWheEmQ2NPqf6LaN7jxyDJ6Io7ZP2R0hx1J
aClHd38ABWWQ4dpVkrBHpyDqWa//Cr8XwDoFEbYZQCWTd+Owo7szxWteOzeah4bT
UBk5K3kqwek9GJ4yPduBvRC2s72xoejcG0yGYr3MUf8i6b5llWnBt/mRxfkUfWjw
E9ogY99BV8iZvAncjRjhYCrrgHdMdf2+MihsFpI+GCbMNW7I5kAFVvPA5bkf4Dls
l+pRNkXKRDiZ1Qxe9z6K6+1Dq2IBpj1Pk4p3wzljXbA3bNc9MZiH+/VHDOJBVGlk
jFql6vW/AmDR67aafmAkTkpXU6/Kvg3Vc4Blwj12YZNdPqX7yzBZgv6K4aFSOmWA
mGv5az7ez6qoHMFTnW16dBqz9MqlB5yk10kjFiJlP1JaLV3bgbGlCLgmAurWIZFC
E1pek2oiuTHgje4y9aYzLbvNIpv16JoC0U9agXjrFANubgGqBEN8r6OjFGO/KKMH
fZhVdR8M9rUiWzNaTIYZXFrZ1+yWRONs64WRgEe0qBhHSyy2/PJHWKJ76lVzxbD+
96rl7f7SU0DFnDxB1AjiYlfmsVOKLcV9sqlRtkJGvdd1LZ9sLxd1OGDutK+RU9iI
JieGo09UcophLUu3fFOyFY78bgeHjQmwva2Eg/TcXClPLb3SNW8xtQUcVeEF+R5H
yGUPRTi+BNQEzMd4oH5p0jj4A4AgUrmw/vHknhD/jfj45QXVfYH5fUUkRB0nGAQo
ttFgZCkAlR2TQTRmtp20eXoU/KX7HNLnlvxZ4qkQnD8ajQPOM0TZ5yFsBhTBgs3T
Vy4o4SqRHsqI1jd4Y1XJIvocYxoLNQhF/0P1QjFX+VPibh5sthzwWGC5IA+OY5Y/
1Yk+VKvaVKo4Y90yFIQcBzL/d9R6OG/6h4KawIirKGc9ZrjKaz1Mn9NIx3P95V3G
LBC+gaetLZNUhjPT/z/DfgE3jGx+3rS5G5fCTGhl4TrJjBmc7eHBhna+dBpWcyJP
ZWELXFpcpXRJEhSMMq+GgHNPdjdizBvQx2S3GT9szfH2I5hd7wOU4lpa+IUfVpst
8ZTDM/CwB5srio/+pnyL0Xz7QBpGsHWlsXzM9w0071BeIL5N5yC6KvukZyHB3XJs
tF2rqq6pOArb2tBQe5eQ2if8JQr4w3sjBceBkxqfLYlsf6Pj6hevHaGjNe/WTr4p
4ss2h4M/Nsk1kdFQY4T/T0MMY4yBUdw2P72v0wXKaCgdurpTqFXd7hQ4ETl/G1XF
5r6l/QvHFfq+n0KbW0Qnp7ivGnLmIg01DBiBDI3AVrOG2FO01/p8wc5gAdLGe4xo
EKfoooit3ky7a+RZTrw+if56GoJIBMJZRXkkfiFSv2VexhFavsgi29Iy1LV0J1CL
Dxeqn5jc4C/drsaGDVYB8tC3TFaC3etv66I+aHHhb/lGq8s4bQI4A/4f36MGWP4V
VezqJDzeja2RXE2Y4/l96MNyKvasJqF31RBy66dm1zw83Rfpwa649Uq5fIbhkBqX
VC85Nh0dzb9kPr8EIXSocS4YMtb0Uvknd1EPByXintvplB/SByvw2GqiwxGlrKs+
s0CTPFcnIbrEQ0zjmRR+xZRvP2t53GO/xAW/+Vu33Mq3EtTDJK0KUlXPxF7/4KZn
WE6exdAmPI5zyP7wCZT5/pMLrW8w78Sq2dpK68AQEAn5cx83JBD8O+lYVzE6+B0v
xn3eTZ9+dvh/efSnnm1cEx13jHgnvrms0JRkzxLUmwtt4ctFEwPNVzjpUSd1Z8RJ
GiUwkPt4FTFebVwkzRaXoWhhN5nKt5MvkY7IlpLJi3Fyjdz0pvaNtYB+aUOWtHOy
0c7a9w02mGgyFE214V07j+Ro5oT8qXFRLFpxnv11IF3ublVGEPuYYHpbq0lUKNxQ
A/+4po8smbOuElxcmDji1rPvdNWkXjM1erMl3z0qm4DcGLoYGqYWJsW55p119Bfu
nDtCwZIrS7epdAwb/2HlDN3lwu813ejm0BOXTnFAGaenpNu+lyT0Gnff13q0zHjG
tcv19Xs4t1djIGy0aeUKAewI7Z2m3UC50jTjof5SCgPxqqP8UyVbJZgCWnGQWaSd
dSkYSV/mvh655a3ubkuD3j1aB+U4jsQ1gHQKY3oEjjrjIp7+LzMoj6ILHVWSaNu6
rtLeKzx3KWyTNeospcYhbvY0trmxN5XhU7hEhbEdp2GRf3YUKcrzxHSf08Taq5j5
gY+hZ8DXZtt7OSRtC2IWXi0ne7mdCtJpX4qC2wTmJhUBMQn4BdxcbldK2XA0gvG2
YTN3UzRTRcUtYuZzIWMJVUOp8qeF2Lfnw9tb7E2lLpPHifhTlEwVn3hNXCd1J4ju
BDndumZ8tLL1INvcKYQpGvbLrc8J3d+RctALEVdTYQp5vdCFSmziXtdntgLzE/zW
tUkvsBgasyzsMW5JBb91++xyZlb49KoWdTgihDDAi8IziroualCFhHnKBXFnlrOl
6O0xzA+J4TdEC9BcYu3iwHjRjsbStxJsuTpnhET4v3MbvGBg2hU82GdA8eGEcLwV
rCbyccbvOLNq4Ta9zn3M2DJ8tedSamyztqwJ40jNPF6+IRyoKClsCzvllp4ES8lm
FDHuT58X0alzQKIMEh1pjsoncfMddZHryHkC4QNeV4CX33IYYRVhAISVeL5bQCUb
fX+wzqyl57gJzPdED5NYFCv042JRI3PlacUNyRsWdw7sY4RmLI78eYRE2CbiK05m
BUVcGOMxLXHDrTov9mqL+GunEWRpmBhHxh32txrTjKmJxJ2PnQZZxCb+Z8SwNxaB
oM7l5xMDFYF5giK08l58ybtLuc958lmwJSlFrVstonpvVfXgj4JBkwrX6Z/TWix+
PlBJjl4TOmeEOw/E+hM5OXLqrQlO+GPf8o4mi8oLhhj9aPmEr61+EWxFkaKp0j0S
cnsELU0+OtPxiPamxjOk7oV10lXien5adZtnJ/dl4xPrQAELxa8LtdUzMNQzXiqT
mdLIZDwMxY1hPGbyX0CWHnRZrKvbitJjYv2VEHyZDC9NpfrWgGkXD+TyekoG5c8Q
bZX71Yl29R/ijFsps6Wj8bT1dDXILRw+r/usHTqu36/RXFS7SaPS22DaZs4CQJaX
1NP2wmwQ8Bq9NA8qeC+PSDq0Ns3hLaCmtca2/mqVvAFTNPqH85BV3YGAmv2tqlvU
onlJdGsrJ5swDtsDWyx35qr3wYAC39G/tGpJXkV8L0Aq6sy963MgsqfRATcHUMHC
5AS8J8tsoQXz9wKvIpOf8kQFHKK0njD9zdKOGEvEieuiKoVOzzQJzHg1oZpwD6Ai
PgnBz3xEX2UJMqcWo2DWSlk54xhZlqTs+Uapb3q2k9EdA+Qh16U5ks9TBN5hSNQw
HpWerXk895VR2rdtkt8COh1/jMCJFOsHW1kU6+v4Kjk3ClmIbIR0N10Nbhu04Ah8
sEKLUYRdMnk4E4Mk93rSPZ+aYLMI95q1l30LWvV4UJr1iWCK5GMuwzlGCsAV04HC
eHrD+DWZBZ33cNhn0cQ4xvaYwbPRiSsTcZmKc/T6CYLhtNEpZZqer72nlgmKhyGW
m1FYqP2XkZjxHNCAF0xm8OUH7zXhoCjCwhKiraPGzUjFTQCOalamXWDq6KscXK2z
6X6Q0XhejpfAlP2ToubhdTEUtFjkollEHp4yyX6LCiucZgIr5jJMUUgdnd/WdLCr
NPEXrnnX50Hl0/ixCmiFFDtSj3z3B7GT9eespzwqnM6/Igl0joI5x9fgq9C8TRgA
uZSz7sDHpdHuNVTf3Lw6VHdM9+0QlF2XT49w6xPZcvpNwKfd4zZA3ub5JALtfQaD
pdOh9PK45mGHzOLgWLT7CwPksrqmyqNAvlYB4qv3UOg0B14NcC0thVHAnWJZ4mwN
W4XiOWpqQ54Qvv8Iii+GF+tibwrFyBTSO9tBFpKdM2yOL9KHQxXUvpbrRMZv/2Wl
sNaTCVmxUKB9f57BZHtunvJ6l6iblVgQoKRBIx+N4qBI9yi7nGBuMksU8MuCilom
HilnF2Ob6dZD+lQ8ReJCp7jIitFRI+znVnrXTZn53i2u89EOO8QBHElOPnKygnbR
I3rDMUFqA5l/uSoVlpi1poWsEVDzgx/e+GxYgz1gajCy1eft9t5NP4M7DRrM4X/e
rhoCExd7kNw7F0dD4ENiIap9z84lZzdHpfK6qgxxsK+8PPRqNWI8QiqNd8ZyK7V9
ZuZ/w+VTdHMvKa7QoYtbrVQfSEm366CBnZDTKqLn1ADweCWdhAJaZ6FiWPbHnXka
Vm3lS0L62ndR81fycT1VCNFdENmnSFM55gV3IkJGz7d4vYh1sLBFbHqdlftaIPf1
Z87rjJMmPwW/Kgiph47lrFMDeRYoXGPRWXS3038syWnVvtxgWDB8Pl6gqooWzL1D
knlguLDxnAwyvMMwUMOjaOdfVzfk31RtYl3PKr4XPsDpxuJGlg2FNMyPfhK9Dfyq
sZF5YWAxD7TXhOUK+UsqflgISGsQ/WxC9XHnbfpaCnVNpPScvqiSULL/jIOdEMrL
HfIZ5FQBmf7Qz8bVmxzGxXyLFj7msHL8+b2Urlc0qekZ8khSuTIE1/ySQLoUsqNH
TqXNUaI1d0jcgcloEr8n60zJL8CDgIWELhwN/Ofdmp4k12fZOg2od+4wRX2lxve/
0wI7YzSA6EyIHk2HCyWTA5xOpzQ4C/g6g7No5Il5XB/cl+e3LvUqndBsBGkhIHVQ
PB2jZG7lswVRJRfUYf2PdfynzNhonNury6hCRI0XV4IdMuTGt3scjJzCEcc9SEtU
UbSnYBARfyLhttce2RLwDeD2QX+HLjykLnSA9qsPQj0UiGwFFRomqSOn8fcXsr26
/YfY21Lj0O7Idb0ZmAoaGgbMRsbRYrtFHFtShsVjQkTu19jLqEbkIN4dp3+S9Bnl
HVkCiV1UJQMnRlD7IarX6nJ08xKFbrdSsOsmEkUy6xakyU41RVnm5APUys1I0ckO
e71IS66ujwuH56LX4k5IGTeyd3eEGNdHNlSGqxO9HqekU29j4kBdBvA7dMGMSDbj
VmPM7t37eYsz6zC7MM2TstDyGVVPkYT0lJ7+9KKoSj7YBB3rHpeiaDIvyEH+5Tz3
5r92I4N5IfU4uJjlpFeDwxilgpi5380VSMAdJC49hVMPeoG/UAPxbhnH34SzwNPO
BDBEhtnskRoZ68yCRHB4LbgPxjeAr7L1O09Pc5mvVadMRcd40bRl6OA7JL4eWpi3
8KME/YynVJCvCsSmGKOGiHyhcZ+E7D+iy3cjM2SgLk2eNpXTfZS3CErODfuL7n9J
IbNquHyIaX4MXIvBWHLY2Bu6HkcgVMxZj88snB3xpZ9K4mCqISykbJKrLG44Z8W1
/1PnK46vz5pQRaR0dTESnawvE4/VC7l0OsO8QFEw3ga3zX1LqsBo+j4nWKupgNs1
oWpHBeZkQdZjB+8srkS2Tpl1x387H8LWZKf3eF4NcJQEocfUOphcZ7TZax0oIKNJ
CzcrB9lqtktiLMmYEF1Hy7v7hnwI3xxy0h3hXB+2C2KxwjQS/kSwgtp5dBI5DqXw
iSWe9Zp+rE8uy45u9FGO8n304xhbIduSW6cRGLXmPAHXbHLjD3K7mWhOz+gRfZd9
TUwj8HqLZI4IYOdXN5MZRrOTlR2m8utvH8abrQ4LeQSWfm6zn4AtP8cH3L7A1K52
gPfCG1gWMKfNXQueDw+BKQmSIG83s+8+VFD7QPJ0i4jandsbe9rZJZKVNNcoPUWM
DaDQvhikEMMTuIRCXsUWwYBMl60DIfnde8f1sxuJrM2UguThdcdvo4/XEUrboVDc
xd4LaXxdHBs5RqH1S95uji9cvkGhsW2lm8jd1oIxrZrvnilPFxWjYiyY3HPyYx7N
7UM9vxYw/HlENaGhqB5636FhQSDbJG8Eb+pjVi7qqs1ryu4FmCiS4dD7nRsloGFg
HAmPOkJ6YSk5z71v0o/tpEd78kkaw1PytLMYjQhPuCGZ/nssxtfR8EdLvIF0HHaV
WX4tV+IGwHv0MhtP81Op+wCigKc07+Wc1l8/MCjrqKvtyzFt1GjSAN+4uSTdBSwO
QIN7+1PKDp/rM1mSFx61BW6uhoPn3J/4YOgaX1ZgrT3FLlbonFVnmtIatdmGynNk
ej6ox9Xd2zkzymlVIv5TxmO2GhnSz+ZKHGa7ULln+VRclXn19m26sWecksvI9Vqo
YLku3TxbFo8OFryFR2fjbsoI8TVgi336RpcjiAGbzGzjVF5Z0D/r+CMjVJB7mMV3
C8cuNCLcPEMAcVS1XBaaW8rz4AbnE7dB+8STc+1Y1FaVMKJnTeasqBMPi0E5MFle
UWQSPf5rAU3TJZN4kVsUzxSbW5WTWTOjIZ+KAROfbJFvufSut9KjySBy+ugN0TdI
VxmUiDV9E02Jqts+HpNdHQFVo0fsfjDb9KI6pwa97x1Nona1l1IUQO4LzL7GErxk
hZ41g3aS2HHMMNiFEoyvvQncQXIiywkLrqnx3/NT9OV7eQoO+z5iPJF2z4GkWwxA
K6Sy9zUsLRedgbFpgIGH96jlIZkpzhBHIPhNk6WfHdJK6sCmGLA6FtlR4gci0Akr
QgbgVkhY8HXgGLISpusGaXMBzX7+cWPG/jbok2wmULOUQ8cZmoTzaP0Mgj4SokMC
PaQBpZ6G8uCklaOZPmfHqM+cW9aQ2u3JWZAmUijCxr66Sn4FIH5OTqE8HqWv5/Y1
t07Yt8wv1AzIpEkaPEJV7hBRf+dKNlVOn7T1oR+XUD+ZhIvvdqkHUm4giKSeoXTU
BN0GIPpD3EdYAkUojaS6iSIWizk/gZgHUPfB5W2dFT3KNr2GoSqLW2PGRZuNuNX6
hryXUJ2iyKhp5Tc6dFQhSnlVWA6kUwU9SNsfdM7SdUV0smrRtcxdt3iTDzBiEjRt
vF4mmidEOhNEzhya9thTYEO2/EcJEYlbPneAzfTWO/RRSuFma4lar/BEWKDlE65V
zkmESjtBOrMS+fDAN8zQkKU8NQSttEHjYzOk5ZTwJdPYok5Js0LzoeMkbUy7X7Cf
iXL9FNnqe0RBjk1GtD1biGJIiE4mJ8B4IHXEAMLaU7xSV91LZmTcRlI1rpo4pxFx
PsO6rUpmRdOtn/e3/NrMxB9/9gIQp5Fk5Vb7OTacx0qaN64mNbig+XnFeIvD3T/b
9JXYI42uXftxUqwIdr4gHv2Ovf/j4xiVjXMqK5fli2f3RJMl39KnTAlPGzPFVBH7
sVvqAUygh4g0ZLI0O260WAF0k6SXGDPl6B54MF07ib7UDiWhSbb7eFvzotlfsl95
SCvCqmwvdg0iYJaaouTfbe+x6TBtuJfawQJNX2/+G5PCkqzrjzmO/na17itBgzWL
F0vbPEOc8+xcSU86LF17JPF5ZRxM5RHqa09iwCFPBSFwgJptK7lcfgtJ37XSHIb6
h8sa2sJF5RbuKkFQGZpXuA66d0FoDcF0/rZDuoGrD3fTqVO8DYYPmNGBbErvmBJU
YuLLoVpSugi3jBmShQoiSl/GwHBqOGEklymOq1XcXng7vfpEPU8pB1OSDKRLpCN/
TV9zvssGyrToM+anUas+qDfVz7nyazbL6ShEbJ3csIG5Gz/kLSanZT0D/+u6SpS8
Dy3VCAYwZqqAhTFIVP5fQ1HnyMIEyDYBlFDJkKEyy033MF+j0wYGkt/dtmI/6anF
6jGs8awnVXLw7+tRpf2yE7XsW1juNxa88vDjwNRUbglxAVgGCoD27kT2zfha36zc
U8c4c0gR+TwjcK3DVN/36u8bBKBaiHfz4TrvvdL8ZsHJ76m9t//Jia0uyDbRTUGj
8hGWr+XQl7wFil1t3ATk2BV/u+muJ3QVeEGGXMNxmSXne6D3mfLLq9wTijI/Rtis
wGbQ5cWIw7W/wnvqaU2jHlBDbbC9+mP1aLeFQ9gHoMaShdq0JMQ5lQ3LQrS4O0Y7
FTkm9dddZswVO/afxK1jWi0wJNrorLpoEQ5B62paWa3dWw+K66YlWiCLeYlDUokG
rzCtJjMszBJ7Dh9d1adeeYpeYjGXjxzzXiuWHtzmG0jXN2D8DfLPtHutRn73y5Og
MRd5THSS4BPqQwGANg5ENQa86iM4gZTOEtkXIP6214Fz0fhlolxkWEVPLaEyfKSr
sGmj2fWC6+FyQOR4qDAol/L2ZkH5G7G+X50VdNrbTjsb3Ov9xHBIaIIAqIm3ej73
cQVaOOZ/xQCG29rNZIPp9hMtR/G8OSetWbFzCqJ6+FR+R4K0LgKWY4YwxDNlDVtT
CzNJlifZ10IoyMMgSvnKGTb3px/53Gg4PZQLthZjqYHTBr1W32T2INI1gfBkWX39
R9MOlAYdcjM632zkcrz4El93TpMMPN7CO4xBjIxznapxiQMlrOyw0CnxEkyCaols
NEsw9Hp6aRwHSutGtfdRRLOGcis5sYx7o4STEPse76cxM8NSS+faRj4ydrcZpMXW
2YpqBsDp1e05LCwKYpinG6t2jUu8LYJOtS/lvI07N5zIUx6jIG/0ldzoyd+x8sVi
XKKFVzfNwH00XAXmDcKOu30RyZzgA0aFAPzu9QaoUyQ/YYQ18i+ufbP/MRzaihEB
nsYcJHSg+u7MfA6DHdicfQSmH6X6oWgMGBd8nfk2u4CIXF4wKZeKkVj0scHfl1FG
cDAP7N+4VKLt/u7gGqFcLZ3qu78VIysBnPWPFJEwPhup9vVdO/0V6GvFI5lzsKc7
vItpEvGwRlpY4PwSr0ItA5LKw3zotPoJlmW2eq7XOg11/3nH90b48nizaTEhCgM8
PatBco4M380qxROcA+XZsVC8ayNMAjV8jys2zU4xpoEFIu3wzQQBJOy6+IHauqQn
hYCb7INJ7QrnSvhX+44pHQmu0N0X10ytUTfBkJ8Xjk9bgtiuS7EdPNOyt1Hid0Ss
K6dhU3oVX+20bMUT9LEm9JZ8TQuhcJWN+idTpqtp3UBWrdZlkiyZKS801HxyfL6D
ilPGb60J8IhiaLoqHHf3oSkymRG/T0oA9OqQPneCqfGtXfW/GyvGU5eP3JK/JMeO
D67QLKMjYtGpCSv5FeySJZPy4mLXlQHjkTtuGxp2RuKGojnHtaSCzdMPCTVqPCKJ
NI3AT8PcIz84ZONmC+pBi5MxWUwWr6WlQDrA/cIsneMSz9OJ/9r1x5HHMlZgN1oO
5bcU2AuuvcfwCJowY+KDawXG3b1PeRbcnnBYYuY1fyahFd/jtqzR2E1txqz+rD0l
VLuj8eEWy/rB+yG5WMb6KNHzAmy1uj5pwHQrXQ68bOxZVOBaEL4MrCedbj4dPopy
FprphJ0s3g3y0+bXWzIxGP5MCF+fBbDGaA4yczloUuqpTMH9mICm1CBQULOuZnDp
L2oLUmqzHQEjGYVfuLM5PqsOjDrVC5t/K4QohDECng6Srs4lmmU9GOFmjMjQDUKx
uIilJupKMGP9wJJtgZgoTeMoAFMh6Xme6+TxmPW4hXHF+8P0AOihIvFQbMTW1ZKy
5/0YkBJzEWl0Pj4tQx3FF3rSDg8m5Pyz4lCTgkLYrrwpOfre6HOvwmfkUqpMEUJG
hwLmr7OWpNnFnDR2oBEW6r00jjZSLbXJCpLMAXidtJ9S+D+caVml5YkaYz19EdEP
fnhvsn0DN0+vOVjAFOQTH13gc8sa9rQA/hbSrGOBBvUF7dcESn1ocWSUzyRdE8oe
aPubm5ipFG/D5zt8yQF21wd8rj3YJaeNri1pfeTaL+BrOFs3NjEAH62jv0oykC9s
4wJnuZky/weLMiFxhWghUlOYvJbIw0utcmZjWM28RRWmlurUX5RPRG6JQm4d6g7H
SyCHeQz1gjU/cBl3pj5cDVMCScrZqhYWT9YWjRr7wLw5W6ehBjlji/Fkn5iQ57uK
bgICWheBa06oPZ4LRBDNI46YPEWqT7mv/ICWtaPKaolMGPPrFO8G+cDJAIpTv0cc
zjk4vg2H7QGyqo7xuoiTvD8Eqk13HVElkX4eRyAbC6IW1ftsqtR+nJek9HZs3f5a
Moj6Kzn0ARWH+9/5TKG9Xt5YTokx0ZvAiNUaVyKXnkLl9Vg9XLG2+cjBrWbk7wrI
7rt5d3fOu/CMCT4uB+lEW8DsfED5T2V2d0x22V7a52uVKHUq699JavXhFdLPgsxv
GJTDxigJROOIM/Fimj/a7GYsTEaxtTLRXNeLmZLvV/NAlHgfgNN2wwWJnxP4sa/T
cqAXAl1dL0PymwkVS6rGYRMoosvYbjPZKshMc+C0mxLvlo18RNTaQ724M3Skwx7k
LCA0eDBztLaF1EbcAA1KWUAIjc4k6jGPcVpT1B7Z+vdEhutkdnzmWT/8zYbnO5P8
hmOBE7Fd9UEyE18Nod11BM1RwJ76a2tMHS5nzGpGMuaKY9hj9VfercIcSuCQDmvR
qgdTNTBagkXgoybYX+kG0GaQ0X6v+AkQOSlnyzqhLLgIYgR6/wLoSWGQhdeWBV+r
Yh6L+gDhPQlPY1sDoTX2dSNkCh7CFLE5OMuCX+xuT1DSg7+dKCRv59aK3adEXlqM
wm8lp0gh9hp4btiMeDgk8VopAldGGXkw2QCTZPGQkyFwQNtIuIunf0K9vKirl/vT
AWlV05UYF3OFCWMeJl+FLOgWbvP/2pkbrxSlq8fsxfe0loxJm+0pb6j5bXnqRki6
zWwfY7Hv985aYXFqRvpeRkgg25z7lWMOc49vazLCuGYLktVXKAverISiIqFvVuCr
Y4SCYPCtDo36GPAO3U8ndvIcWW0AUCi//t1Qo07CxdxbL8M3YdRXXi3PwgP44NRo
DmByM1Hntpgv3EMOv2PKqddDGtkq0bxdHQWf8m2C7HVZCmvddEWmi3Qc7DTgYg2v
50pva37Sh9K9fx1WI1V7H9KKp/sdlRY/P6EsVrrDv0QIWo4jMsvzdbqZKHz5Pk+a
rWNu9MH45lFGAPOCMz6+YrjOIdVPWQR0bAmXjYm3uZj1jo4tV9A1mGHfYQMMWX2f
exG4X1Dr98ZB5d0SQKgHlfqRAMSot+G4jkZqkoG+h38qsooAGON9QMCz58w6QxkD
QaboaCKEMfZNwtklgp4EfBjIr80aIa1mDM1AXXpQNRRKvspoiZIXSywydVRDm0Bh
+5TlgbkR8Crefa1apWdw0Oqh42vgvlT39eWMWCDe0vN9raFKlbuZgtRvdLOcFbIw
hKk8UOM1Sa3UxuYq1+Gs89r/S4KdSywk4Ya6aRJuGPa9+kZfP8yFShfKQBvj3CDU
3wKFKBonP/jwFv/kl3Yxa4z1HWKm6nJqF/Lu1Pwr3IUhcwiA931sS4585rgK2jde
SjXsW0Sl9euzqqABFwmX7E1Ot+a2z1oErPi+IrxIhcw8T5ctRUg60cxhLPnxRxft
+cWkfPR158noE457LQNHAA82h8Ibd02rXrb9dZi40TUHG/E5CnYbdWaENm6cBhWK
I00rZBNNvJ7mhxGFJa1lP8TL0L/q6NFoi3+DpF1OUqS4D4oP6QwEAyTYbRFGtkk9
qNb8Y5t260zyemvTB0qVZ1JGQZswssyUiwX1aHFZ67Nv1ihgsg4qVq/e8ZIU9JfZ
AgkgiGlgMUDAzwUt5hnNWQMvL795uLgH4fQIdYkMSATAc2YVhUhy8JwJORULLI2/
w6ICGEqV5EXZajRnT3bx9KpzJyho37Tct+gUuVk7sitmfR+JoALfh4s2Bqwq7E5Q
nMyblEFhuyNCM0wAcOhg0uRF8d2FN+tG93MfMX/5iFIcz+bxbm5vzju3HTe5iAWe
KdB8FzBIMNEEb+VuP5kWTu8vtQ/bhlyjj144BwgXVci8HtuMCGrPqhEtARMg5mJt
L3bbYFd2mYhB8yyZjQ0b4eAc8Wsqya5dHkwlPpmx57NSCj6ALnrqtSUHqv43Okt5
+qpQXm9BQM/CzJ9R0wtbr32OzMlgQfgnhVr9LsdDEcltWWGt15OUV+pbwCcSMhSE
8bcYtDIIS4sSx3D4enONmQ6n2kr17ZMCqbsGsQRTwXoV71dWLM3KonhdUKydhJ2a
oUTLvM/mWrBBsgFiLIV1fmdSKsNRstkX8EaDKsFu8p2o9yeQOUypzfQYfAdcdby6
aOuqOW/H9dQylpARF/v50lcuz/KbtAguI46sRr+HBxeOROb33o3eUcWDUTw4Y9Vh
JBzuPL4S0bTftw9dKAe/sdhSTHMEyY9bWAFSEEJ8NrSc0AY8exyxlzOQOyaHYrSN
qEhmE7VnFPWUHlpLUK7qqbzvKgesVi6bm3Z5jS4jQLu/2TyCcl3xZRWHqOIVnspS
ql+IR3aVYSY2dTbsFFKjBWzVD/QyXyYuRUNKn0L1Fng+TMocW8EQ1iD3V62UxztG
Aw+q/9mhrZ8kuIPTEhYRPNle6FxAaJRvdWIhzaLvo8sP7h0ypiUlip9Gqzx6vByt
SNzSqfYtE25ORahdHr3RZLroBc4qpmVN7CO0djieyevnuWFh3F5eyD4Pgp1TTcHW
P2Jxj1jzkX1bjyRxZztH/RNdubyjiHTxlawB5eUvxpqvFyxN4qPrQMXm6U157Aax
wmmht06Zk7Ax0Vk+ORl0Qa/1dxsRElSKSYYvz9Nz+bjJCHOVQt+kM3iAmrnxYuw1
kogzdkqTCFXm9EUTmomOmtZ8dcVPzwkEfHgQXxZHEg27QdnvZyIN0t2qzTKansjl
n2kdwS6h2vUnQDzgRcToBXgG9Th+WBzT1Rdm8LLxIVbtT2H202tRAMd4RPmjD0JC
sCVoRJNLdxkeNgDXSBq8IVWC+CS11VyJxK0yj2pdJDNbqwJpttmUirt30846XjUR
3Dnfxwo2DyNERF6oFL9/TEMD3PdwZ708WANOO+ARBxz7JcOCnwVczBOky70GCeri
p5ya/gCHGApL2fFl1raHIs2VXDxHh88z8Rqhy1iHxwb3ASrkYbTdDm+kvkDmfTjL
+q+icvWWhRdDkXgktFAglOq8xI95rNQwiXZu1vocqVhMiQKIk+oKHprj+vJ7r05+
5ssHAzx6S+HvoICwVc+9bi74zKXJQyDLm1CeX5npbqaGYAka8AEDdZxxnRYx3sgy
pchuO50T6RouQ0ClCPfZGYSR9pQ6ogpDgvNj6wJ96JWppBg877JelABsIEbGy5So
j+xSNX+FykM17h639/H5DCDqYyCcnimS//KyWqY1vkYQZ9lSe+JlEQOaXRewlEpF
NR7ZxeO1hnFNnESmcvu/YMrYOmujEZodVjBuNT4KkTABKWGpDULXLI1txHFLOYi6
5P45IDCqTeYDX/77cvkXwAoBYpEjpl0VdJ7drhjr5s5eE+UBJW6KgdR5G4pKbU9K
O4I2QJxLR2W6iDr4CIQBc6ubeJt55Pq01ssLkWyVIWeHbb9f7jEn7b0PYk6DowFI
3x2ynDgsl2o/iTl5B96fe/qsa9lmYSPy7Vm0Oo9e2g/th7IrVPVszfnqTsm86/FL
Sp+5yv9eVqgNKhHnAB5G53tUoLZNmmEBjX3tln94fn8cnKnUgJPuyJX0zbq37cCs
YiZDau0Dnn4JAYzOOV4SXkQNaI23v6xgclv+bctJS3LIckJdu3gfAemHofGdB9xt
nhiThYXHVL0JOlFmTQ4syrmHtKiH6YfkMWMMFMZ/ojR2bf7asj8E//Ke02NbkrG6
QrjAhxUhkWzPRugTikCMCgGNlo6ZfGZem04NbthGGIoxXOjjpaYWTvGSMsS1cXjQ
2mjVZ+rX0jhRcEe+LOt0oDNc2zfvfrLRc7VbH3doSaxxeb8p9hJBP2fH2t+wTcg5
KmatAsP9fnrqrzYIICWLDbOlx1obZxsTL5Gq9P6gzqYI230jxlDETzX47ZQYSr/4
zCe4ZLF2dER5AyZFChNVbDPJCVcP7Swvv1POIEEtrG3PZc12OgsLei+wQUU3skU4
w3nOnwcZXWND1HmYkj/sZR7Hmv6NXERmmc/p9nM0Erj8EhscqjOpGJCZ/LOUi+rZ
jGZne9dws4Lq7Z65VT7MKljcKqEdPtNWF6P6Ou8e7HyNS+C0bBDamABwUS0rTvsH
dlO4Bdjqw+ELMuV6sCsgFzOP+XMXOinFUrNyiwc/aZQ03B5lp3jB/OHFKrAmRDY8
UgEdnBcrqInCvZKw+fSV0EQW+P3wUUBNwlSJ9pmoVK+CgNiHyT5zsgDhL1NTO57y
QYxddDXhHt5/6rT13PxvdP1GEl7i2Lr7NuZO3f28omrFzkkzmfb26jrtU9AD0DLZ
h0NyTUdAUyJnCPXXbmrxhqjSkw1StL0ITMSuf/iec63Z7c6r2Z2gwy+O6WEdGBB3
kIikvT0AcTd1ak4tfJckUESNx786JHKlqWVLpV0wTV4/0gdcIPNfSZbP8fx545th
FV2PfjXoSaWwQg3hpHkHaW0dS2Rg+RFCtqJTmRZEPZfpVtgMcG1yX5w/YjlLdgu5
xbNlkg/QKHR770bCkiuvxdV8vVdVmXCbkmnq7BTPbIoHj2/nIq4ftwXE6QPr7Whq
7vl+l/VY8Vn0xPkxI/+105rWAI1VtKthrxFxztJqVx5/XMWzwsnbpgzXBvOSnuV9
qZG40SOvZqAtkgGz6KRoI31GQVYWqRHt+tBmoSbU658Un5LunCQeZdTT2gLzYjf3
N1tSdd6NcAik4HMlNlwVdORLl/v3Rh7WVrybkQLq5v9j3FCgpxQFBWovb2FtE3We
4CzuASTvZ6s1jVI4700FtU1TZWv0bTiDZqkd9A2VGqgmCog4pWFeoNqdDRafpTz+
PnALLA7GKmU6f0ImnxlVt7/1MJgkpsjwgquf/IwWkP6XDWLmkgUaxs/U3s7SRS5N
gi5iGPAS9WugX2Bi/pRCqOOPZpwFj4FeE/msoFdprfwePP/4cMt+g87sppZ4a2g/
7bZ+j1/k/5mFTbDjbBysxvliiQsjaeGreQge4KJCh2VkJw8NhUVbDUQRpuSqwPkB
fYb4v+VMXvNWADgMjdo+zP7TLppaG/blWj2pjkKWCCGzumdfgf7iBumvRtapegvn
nWlth/TOE+gNMC62FWgiZGqtsdRVGQoQGcK+KCZOXHnU6HDQBp8xe0F1oGoyqnXE
gtylDwyOYsZsAfsa3fSFdtevZAh8C5XaRHzRgc3iTHnfqnNUWQtleD2lwSLCjkxP
cavP0XzwPCo2ScgIBoTt1BuIUqA7BDfs2J6HrpU3Ldofz+N9V5u68qbSBJmqcisy
iERV2ulu10/mc3KLtHd/d1SOuAau9wpwf139y24sjgya18QIEak1rJJL3Ltk2Dhe
nQz7uPpKZaoi+logvjplUhWYnHqZhML9mcIxAFBnBINSPZXB/JGr3wW8BTrzI9RW
e0aoPMTBlGn3bM4zsltt4h9qpapXBYwMI9Hgg6touQJzd2keJx0s5JurP4J7Ka/Z
5plREo0yooN2zrwqOt1U5suVYES/kKcdyipOgSc/qgZWj89v6lRzcumYmiJvmxcX
MzPfMv3b80Y71wNvC3SdmlL181XjHbr5P+ihGG5kiCn1Hz9iD7lS3iJjHx1Z6IFz
G/DoeFosT77f+CZdOMpa5Bw4g3wos0a/RLDNnvVVDQmiCHLn090f7xuZTw9JJaQw
WV7w0vSmdcw4qiNvVNJe7HtSVp9SvQWyuWTVfTVWGFdMgEoGtfXJYVd1plTIsnG6
6nZ6cAn4eKCx923CmqbK/xpzKx/vZF62EP2gdasoqN0mv/Pql2p/SOWwnE70UUzi
xRbCUcTdOeIgCHHcVeJmolPoqV/w+MGqsk6m4d04Um0GURI6aIjsR/+XMVdJElSM
GL6U9d+7HCkw0HT/0O6rUPRCD2udFV8tTeZbJ6YflWA2yLjT29qZZnKeJeABt89/
QBKaQ/B0Gcb7iFAPTLHRHo5M7ZnO8FRIq89G0mZwfP1AUSjx1T+ga/ayp52N6jDb
if8OdNDPQCAp+ZFHTqpnO7jGEe7vDXnVP4EWzem/GOyfub6rzLFVYJl/+GdIjXlF
ZdHPJ1+vX378+doYJBHetkePLqOUSWyJ+J82lHisxUH21+E3IbWz26yhHwwY0ZkZ
L/Xj/xg4c17OHuqSniTjScWYRnQnRQzbpB+0P0sw/gyJMbxbdH2gmEzTrfM9jxc1
3oa9HjBWjmpiKyJVNoSfH4KpiSDAKa60UskexdGQxlnp3vDPi0W6zMAwXYJbwfbI
48L5qwJluCNpdA0JMgPrGjHlMEFJbQ8FK1LtW//3X+ldtVr0HED1ukxn8x+iJwCn
phaceJU9UXrFXzixVtGhzHrHZrvoVzq+RRjbf+cBweQ3tHWSz0nySKmnYf8rMyDJ
U+0geVCdCx+NOkDDl84sur1VZLkVlvBrk1tLMpz9u75dcHIlFZdqFSxnk50H7jfE
2X2pApUzCiXdRShhvKDRyHErdrpq3/n0K3azm/aNMCVbNhsk0fOftk2DiymkD/8Q
BFOw7g6Qb2EIH5SCRSGi5WGOHnxjqRxTmCS1Nt50//SDFv5cfL0ZCyilCZYBFNza
K6MRkChYezI5Y247EiHBzmbYN9ooOVcQD8u9jIe/9S0OXQlAurMG3EZHI1JCnRVv
5KnklWH5SH4kV5rgArFNyYTyveL/ofOwVuibSSeYVpxK9IfVbUS0l6yOJj0E88Z5
/XOayBU4oeKZVnejf0MYT/u89UVxoBMsMPaEC03Ant63Xxp5eh25T/QJUO26BHL2
0fh41wWCby6YV6pY5MKgjmK3CzgMDlTxwB1na/efsyNhBG/MRucueQYz5P+c3XV3
w7w1maKktdxaqUW5wQGXemtOpAGWPvv3DOcRdOZjpSGrWxiRdLN/c5nTGvbSi/Cc
/8V5ptrr2Wv22/N+egIQY0h0heIzuuoL8OfbW0EGX/4yOuyCDphviaXReS6NyqMn
WFN+hoeI00jSvpFDlf6x5bujwfwUaIsrLflrpEx3V5kTcleC7mW9FbLUxkRF9i2u
/ssjlBO/M5J4JbRTqKhzfbHkc9nmG7Gsd4Tyv85BPNq/exdDxUXZp2HU/+TPrJmT
9SU854oemYpKIvQvNysHMf5u8O3q9oOGR02jxxn5tWyDxQq6miTZWlmNdoiwFWOz
br+X3unvbhjDmDMAShP0jKqIRAn4pVhO+CVplIYnJcxAcwk9PoEccmxWnqwfbqBB
J0CX1DEdvFMtGNf+vY8nmKhmyo/CzJXRW7qQvso6Up6ObpCO3UmZ0k9YMpKhwY8f
gIY3C1Ka2MGtpsGEX/7yyxPP8WCvv5MpFvAOhV9orZuYwmfBWDCvYkdSVAtua9Mt
HsYaUKX0lvcXqJ2ZOf0PjGY82IT215dMyTLVlMikFmIVmStp5P9MlNRRbBiqHaIy
Yz8OBtIv0MJafj3jXIBGKpncdhr6JybKSMupLOAJbf6w3wjoN/0W3SN3L/HPj6cB
Nwy0o3JCtLHY0Opr9thMOy7Ia75bdB/SBVohpjySl+PB3y2KyoLUBhsG4tDOqv0l
caW25RwhdTt7Q41XMsUxZtm7EJ52buGalS42I/PFowVK6G1ICDvVkJSgGgeq44Ny
lFXS/Q551zghPCgxTyVdNThnvPoamMn85OgGx5oNO4j626OmgT6xf0twOKea83PH
TsBAGkYLo0VfkfwyjpaAuD0aUjXJanCfzfIsu769AA9Ud537moSlunwRQ1BeZevb
HLD+Vz+5B2u5Gj7GwK6bZB63fFCoH05nRMQbTrn10Xc1/UtE2YIdCviE0CQ6W5O6
JtHCnUSPkM3d8V7vElIhAxii+Qc7ux8n6migP6vb8Cdb5G9Yx46RhpuT92RGuJqo
q6WKKJvvSRlMiKRk4exBGVVIDBLdB9+5hUApw42dGqJu6fQIQ54wDTSZ4BhyhzDz
KgjD/oqc88YGvaAw3BhMd9VkCOReHAZWw4KvmwcZ8A5Eylu9uREKk7GDqJfSSHFd
vwulJV6uPkMLmWrVxyjoHpmcEbzWwQueCNTRblI4+tvSei22AcrHJXwnyxXu8o7R
jw2FGeTguZUfr8cVrYc+ddxOlH3b8w17JqybVel+8CcTmuUDTnui+uZggFVI1iG7
vVuUULzJMTWITbaVKO99CHmEZjIQKaxIGlaxFgrVynDzzzzUCcGhsBodH85xIcCk
qhzb+DoHFJ+IyP7vVS7GMZWsT/ru81Htx3yAq2gz3+7xgaZFa2R4QeHkVYmy4LV6
Wjl1we4HABb/fiqpkUJHDQ6/ZFpsOxsGdejH1GhfzRuuUc0dJ3D2gBvQTDRL1vq3
g7v4VY/GKDawKqLgFr5VTtC4vWEhY12B1OmSStsPS5CqJIaMg+bXbvMSbBstc5gf
kMOaomPZWm2ys+GP6WSdfcyiPzC70ihk+acEhWe4DiHlJHUZSiUt1H/jqGeYzSt6
DczPjpcY+xF/ge/13T7RkNvq4/GKegXTmIEOM7Wg/gTqABWMXxc+68FeV8WWASRq
KJqkO+r7iCOyNDXtwaFFLrJNlVtdGZdYsUboAM71+jMj2265Xc+pcAiPEXANbtiL
WfcdgqgmUmH9GOlRt3eG7ZNI6Gq8KVEdoEpodIGaah7vTOb9MC+2b8e0oqYuw/Mq
/CR+4dNRjRx1ussnVTTZL/wDSJi7sDY8WLN9+RGSIr9jmnhb8uvOMMVklyKpQvPx
RkiJMZL4UOUITGPZbvhLpvWAK7nq27K3gQ+IN4PSDqwiAtku+MMqy/Ajf9/ZBkYq
UKgEcGypnHlbWkdVC5/AxQN60n2EyrbrKDMR+2+L7D1TOqd7GoqUFzzaqYGak8kl
/ssGc75rwhXbMHoCWxztEHiQNrnBp/y2UN+/hVaRkjac5tMWMHGI8UfdkXsNlMsG
RnozxUk2LT5uk+sAIwHUdZUBQ8TA7Or15w/LrLDC7PirXyo/QRNqmP7iLV89uiLR
qG5YBBpT0xRzB8g/eWU9I1ELZEqKraM75lKw2b+pZvCP1EQkJos5cB4HJPga0a/9
QyzRXRUPCDl15Am9WLhbVnl0M8KR8Td6u9EWMDi50qi8Pxsyzm/hcDVDeAG4vnX+
op60XF/k582+sFPGlSOh1APHHX8b2lUQFTS84Ol6L6k3wyOij2G0zbCFOUSuaFfM
ijD2x48OJhJ6y9QUosNFn8dsMKlPFANm+stdVOpUEL36dzsJBJ5DKCvinGDr7ROy
yrIcdmTPLU9BiFLNicXy8bPT4FdvRsZLKIj4LVzVIXkYXcioL2DRfU/qP6GbEFEG
Gz262E/PERAac2j8Si0aZCzM2QVOTSAJ6sz2NqN2VXOxuNorU4D8NvhF/6z9+bPL
K8Wg2SGF9BV08HkEBEEHIq73TBphWAW9HwSySIMVlYMN22MpRirIvhXQt0GlRzG0
Wi0YDQcNabexXqeYVyMxl4QmzgcOTrJMUHg4/GiZY3+Z8pNRm1BsSYWHOBA/Jr7q
y684OUiM3tBZ1ZneHKKIEAP8rvKcjkNo5lsI5fcSPn+WtLTH+kNocFWbVq0/ogHQ
SYOkNxTo7kwbWF6XL88NnZicRoK0t8rA9tqpZgrdKLUsC1a5AGIrhBXeRJxsVYLg
+0MZ8XvN66vjDBug2W/l5vevlbom21ygrLMgJrwyWJvv9RzbtQU+0W3ZZeYJNUdE
i1X0QUPuuN8Yg/087GyHam88KuH+urQg+6Z/1smV+D0q9pF8FblhiHHwgclR2/2d
0YqxDKV63vfK7/kaSAeIUvQtUV7zaaumvD1hCF6H8/r08/Y02o/piWEDpE+w5tXP
QTrHr40EURdpr4Ey3sWxO4Bwjkj30NTCbuKi4oidbycQdSXjJkNUQc1hN3oxDxnB
apdGIQxM+h69cFK34yaEI4jaTGrPvUn319ad30lbzlRwFs6+FiKcV5E2R4d9XwO/
XbPaA+JT20P7dIyr0Tv6IjCzCiNn2JO65iVk8E+yLepTGrVa5h+ZZi/eseb8RAgE
bB5QBFugg0qdlB9etJ+36OS2mcxCg6NNwM3fI9Oa7KwFP72Y6fHDX5YqRvcxH/pu
6z/bD3YgbqPk+U5DARY8zZ0rCEEwTPHfSosy2snAnZpsitL80W4ZUVeP+eLDvkzV
7BKXhe2UEmrQekT885+xJ3VSib7HTmu7IrY3oRyx/B5Jfv/scwEyG5h70DOwf4pg
qs8UNjbNqPCc1g0k8+L93LJiI+cwkLh4lqN977khqow3o3QAKTrdVf8oZ5Xhp0oy
SwNQ0PI/iXqY9A1j9/2n4QpGlCvwAnWg1Tv0KpJxiu1DhGT7D+8X477hBm96ErK+
C8lFJYwlSY+e8YkM/HHkRvbGPus1odayxZ2L+PvL+0TyUYFaB6tKDlK6yzoZotq6
DYm7/RyzlfXJ303noIGDZ50rsVGADjXWNQ+D3J01aapkHysBfxuovKA9WYaiHU2h
uszMgljNeSTVfFawL2Yw9R0TkMuzzuQmJ+LBPUWOcpZWcIpPjcAapu7Zw4tOynSA
rcXPDn9kgproU9STYozN2zPGQGJ1ZD3Eoez7f97q1IXe1jiy58/luDVgeQnOMqcD
t3jcC85Mi/3ThM9abMULue47SnuDQC/X7XWhsVl+2qeZ/HfN0vmIdhP77377BhbB
mDBapXuJmhGZiG3khbZkuXjDerRezM14s9K3vp6VIriPFMeqHQOs5ZBrVHAl0HEQ
YtAMNBB1vgLYdaVpURdwZ5BuFu83n0PXXwZ7LC6tAxIIzvBJMaTSpHoHeDSH0oe/
Z+XLdeseVqF8l5SwrK1HlXrhyUZLbVvusAw7JE2ijhsGajQiCV8yDHGW1rUshhrS
pb7Xb3bd+mV75PVAGl3klZfgEHmmItDc8AvhdzCsYfJC6XvK8GOGi5y2B2TEJ0Em
oNDnCyVC9lgOnpuMmD3mz3DUB4ndBnvO17zMZdQqQudOv7oDAbjBp9GIskX4mNEG
mylWwBehBFnnTOSkw5U8lxTpeg7vHKpW8NsMGhPulW+WbwwGgZsOYOLtntvG2QZs
5X+xaC6LtLiWDJDaqysV1m406azu5+ZLSrbxtTHcQzaXHzkfMVxf5k8zj6DCqQxv
sTNDd6dNgGF/pBfXiNlLasrM9e4N3gIxDHQVASUhNZTLeqdoT95/OupaeXvBhSLA
MrSx5b+VeqmNOJksTGmRIW2n5xddnszQpQBFtSIkV0fwAjSWWXWbYDaePLGy3Ior
VFeZccctjIPog6kYORON1UvEX+xttSxDVL/ppvj6GeNaF0BXLBxE8U5ADzjwT3LE
nYGHWAtQM0NZ71FM4tCkK3b3v/uwQpqp2xEMOnnnSvykQUSswp1sgdMLT66ht0g/
N1J9QV/fmdHucI1eUcRtoQzbAdJ2rgzWANdC3nRjxbODy3uQlw4dtj+CxIB4s8D+
nVA1s1yAzkGa2p3w4Nep8w47wsn/Moob2x9tJ/xzDwuIfMa43TDIqYaAC8pK/aoQ
74PVI8zzJOjuHpURDooyA+I01sYyt/iXNMzQfqCmHi67BZx7MCC/tsT7cUS4QNvm
jpat7NLXh/peckI2hdwzUNyJNNPCu7+Bj3dAKKMKbBkM/zsfrkNtm+lBBnn4bi08
aAVzrTFyIcVEXQYbFf61N7gROvusIPEXWm9zStLqwXzfEsyFFGUo3i/jE430Sipu
oY+tfXO3Gyk6pXQdYpKGRe07ABveR/5U5qib/zc7+JewDt73SLiWPPuht4x8fm9s
ypzV9RhRw2MfWaxICUYJAgE1hAfMV1kR77vGaXQf3DLFGIG3rJ0Z4I0/g1RMc2xd
xuni1BwI0n94JdULsn2AfKWhzJGN+dOVfsOPRDYv73gDJB53mrxIkuDSYmJA8jER
qi12p7cfYF/TeanH6UlmclXSiXkr9yzFfnkE7puF4VeWMR6qi0xOF1RKn+ELKcK7
O/TlfSyb+LlMspO0ZhcP/8rNO9SzmUDFKdAgdz97wee0B0YMqP361D7L/JPjJZ9o
urHlkwHrG/nHt6EhUzf9890rYSYF5yB2bqJZWgobNWIcOQIh3Cp+vs9nREkBL7hT
+vklR/xJ60D1HCnpv79PlWRtgBt6nDeGS8E6e2dnjOfAljWJzofMEFFx32wArLJ4
erubZKwx+QIK8E3eiiExXhJTZm2rmwtfdXUwNJv8Yd1c0hMODYKZ18RQ/IJ/9zdZ
/3dcJPRncPSfTHG7uk9voc6o+hD4OIuKOHit2+2MLdUhqvyFEepGHEmy9cPdc9YC
SG2lggGf9qdtXPV+mRmr9C8l/KHSLRkrO2DaySDnRmQo43sBjZhfyTY47lDdH/Oq
oxOyvhwyJic6RwJ3zuA3tXtxTWJvaFP5aQt0WQOPAL8dIgYh2NPnDjMOwWf6mjZ+
cUEktFc7PeXL+znsZ7p3ottdFTed+z6MYYDY3WZOVYWWE25SXdkiWLnsqV/qHj77
bxTlIuUa8HD5wuv7vrSQqGZEWwe+jzQ7cEP8ZFiOUIpLYwoIt0tvgekk7PV0VCwJ
ywI1A+A/KNlLWK9nyBsIk/aPK/qCAnBS40Eu8nZFvctC/f7qpvbK6ciM78k8UkzE
Dbh85luC8DkQ8pIAbOH0DW6WYKw6IbZRGkJ3TmkzsJqAz78RrJUnq9YayBjD7+6b
iGFrpH2fB3ywFExmKT29KQHTrWO7Tzmajvg9tEzjcCCfgU6cJcRKvGX0wJ/CQlX4
buWJ+Q/OJ66FVRyy7/QWcGN5QmnEmmMxIH3Vg+u0fZbbH4DTgT8VAchAQ32nl2H0
QBGZaDyzgBwXWhyib+2KqueEo6cpAOmZLU+yiPlgdEcMYmbLV99BTyrR1FVzWEDa
bdlm1Z0WmUrIWSfs6dB/Dc8reTG9sGWalj1VSxaeZZJkezd7VjlDTE2iKJnTP8M7
J3Zc/QsBj6CnLwssbcMYM0VIZ0mR9pKgbWj7jrmoxXN02S5o0lxsUHxgdGvzVZD3
6l63p3XiA9k+uQIByuT4TQTf0WFhNDqhqmc0rgaTyUW10L1LetuPzBbwMJUV42mc
PsSl9KdnnAscgeWjzrtY8kmwuxSfHuO3QwV7CT/5348crTaDkAv9CPpRhxga1e1a
nqKGumzrBQJdHQNU3QVciwTSE2vmrTFBOYLyXtAq6DjA/fFtt2semlECEU9vBbmZ
sSsCtuTQpjne7OpTKlgVGAETnb5bhXLKp/LWoK4jTmnf2C2EmpI4HDhDEmaRwf1a
O6sRr3Yr4jzUjl0ANfnm/iFxXUpbU1Wsc7a/eTiLCPshn90Z8iQC1n8A3EGBM1QI
hYuMJwj+yKXzeALImdlyiKlJPNbwblKAah/abl2LsD3Xe/m5l02keH71dsHLWgLN
ou/SkFsQJIbilO0iDiPa0ZbS2EWIXCGI0GG1K0h2yAgigL14ua2k6gO2S53Zq7tm
YQZHcL8xQIcEJwEX8WDCJImyOd8uDx5YwtWpQ8W6bLTBMt36xAlxKhSt5hJh1RBY
UcqkAiRUut2bwtjryqm0EKoKVtapWuj/2B4nj02kZbVndpZX8ulvxVSOxc+Nrl/Z
upHjhFetahCONqG2fgFCXv4e+7Qjrp+L+akDg/uPEn3EaEk6cOGkDlzdHvYo4TC7
+mQLymt2Adc4NG0apcdWIuU8G8GWq8yOwOpYG5OTKX/r5PmjEZ/OCBdAYgQ4AzTl
B7xXrvDK9KQD/kTC6/z4weGwwz7foBnhjHmeahXXMUQKeCSi9hwjSZsvt1Ae5IAW
pZY/YfPRLXKnI/nVPDbNOtmn3JEC4GikAdPOdOZaAl5Dw7GEWGrY4j4MWni4Mcg7
0Hs7iV2IjSe1lUluEA6u1s4eaVkxcP+WLDwl4dYYb8K81xwp3zzvJlpxyGDS4EUS
PXDZZsU9ess+7TYttOBE7fZ426psCnsp2C9631Q0yfY6OBsbqU1zSHjcBSZpGEBs
DPwff+HCsD14wUSXwP4shO4PP97EbFaB0BBNiWKpFziaiWoknjFZdfcoMl5K2Afc
YE/opkPQ8O8JNICVVslgyxnrXqb/Mmp9BB3ghTloTzqNY/LRQmzEPNtnCWXvjiqg
jdN82io0TW6Z7+gXcIxXcKjZlg8SrQWiGyZG9hLKcPU4F5XIivwQMKEzwllX5Fhd
SoU9yy4KAX2YIek1khUNTNRAaJozWplEnwFKewcmTeqOKteOfhVkSOsq6Z6te/HV
52UovrfAHPZ2S3/lK6pD6QnHH9MXDOe5pY15bJ+JdiPFdx1zhY2RNj8qTk682dPe
QpS04jAIxKsEJzINPOkusFay6VLHXuukXzbABK6uzY1ATNW5AEZHQnr977P2IxZD
unba9PVpRuaNLS1ReoClBtnXalWaouXO+Rw3JX01GooMS1Tb8CxxF/g7qSeAgp0Y
Y6T4UrPxijrXMqw0P57JHG8pzmHBMGhz9Vy88a2DmahJOzeBUhmh+cHQWqn4ZOqN
0EjlnYfEfS7Ipo+d+OM8T6LZ/fJdRH62MsjWAdAyCpjPifkCUGTQJRXKoPtLZxPH
LXj04cncZabGeLeaMUVRrFBH4dB786uSh2WsrdXnDNxZEMSXWltLXyOkAX4D5PI+
/lxCDa5FRjUpYVAgLO3CMHHlZyFbtY4/oAh7wU9QghZhZbxfGH9lT19ReD2ExSXc
HfGjxuxN8scVGxhjfDvi2/HVgdtY+c+x2kbrKGk6AeTFADe4VYi05bSxSMitr7az
D62HO6XM7JTouxMF5TfnOnu0dI8q0B4zJV4gQW34jaMkptit6XRNaQ9mhl5j32xg
j2FUeHjaSV0v3qtCYmrhf2/HFmbxeWmDit2WxRFjJ/toNeWdRkyxe3nSRw+gmOEO
w78D2Zu6UVjKOQ0ojFq4Nc+L2tHQSPKw3YTIy3hKUQKAiwTdriFTBKB73pQU5l6f
Ia4U2OyH2pLe4UooLiVDT7qv+zUeAP4PSAYHTfVcgaju/tYclIsqk7Sh5n/09VqN
X1pp5dPc2XaKHq65VnR2gOuRdWxgvUqGwVLtvY/CthHUpMYai3lx2bseZW6kyGks
rDTqgEkc03JJ4GN5euk1Jdzar9eddI79nWUQ6+U3AqtTkqhdyNAdk/jmZivNjhUk
7gEi3YWq8OIlGxQjFD3q2Jqi4WtpeygzidU/u2j8bCNED0GOA6XLtB2Rbmvaesf8
2VgZ6UA6RFPzBTvsHjPOhQm32g+n18OcQ20J4AVVPq9rFIJ+l9+iGFZKwTr/zvqt
u2KeEPn9jEGyP8T2TTNqCppTRye2xWMtKD54cS0xPmg/irTCYEAONi2f/UdcgyJq
rNFyG8FjhMhz/XCuR8gotpgYaW8ZllSX2mE0cXeQ90768ygArHIXSkMMtxcImDAe
uqf3gXRjy9biLwDMx2CIquIc4wgvqjDeR0zp012p0pCrFyI8s7D2Mg2H6PgnHyG5
qOjoqTaOvCWoQOGfqU/jQq3O+qVb1LdTjg3/fGw2E+aj1vYa7xulwah268C2PxFj
r0kBHGKVi/cDICGyzQW+C6JGn6pI/9ezUgOwdkR6VCgrJQ+/yu8hdBx90jFLe6ei
2SuSvtrpCNSaEkPa0KWghCcynkMcBO+UKJ60hQxTwQgBkPCoAo5x7da8M5Tg99xx
gb9w933ipnaQ1mgkwvDvztnMGHlWkXzYZe6Oz1Kpp+T/kxeQOnwVSCBNfG2n/was
QhLEO4AV9FuKVbK87EAszId3ch0xtQcmzEHA8tSc0UMUUQVHyewtPUmajoBhCAB9
BSbnJCtZoV6enC0nwrl1eQ34aBWnaVCGAXUAkcUymHExgMCDbIL0BELZtm6gVTY5
7jauBDkxROngBDzqOtQQGoc3OMUx9cOWRJIN/T8+FSIKCzdznP4HsitaFxGo0LV4
wsPapGJErXHJk1xd24MjsifqfJskEUAYtX0m3HUF7sbkk0sAKr7xL0FBvWzUato4
Q7N6v2qY+kGu1z/9cLH385cfmKMXdz1SamKryvNbqcRiTApPt+8IJLt7Dsh8RY4H
2fiGHV+cwwhd6qmq088tVEkfvMvuq6B/xWaksNQBGSCqgFxuMylLVZwdCXSYNKqG
BZ/T+j0/S/SOzhjzK2PcjBMUkC9RZQZSKGGlcNRBSX96HNgMgPInBsEqkamh271Q
BiZurnF74Uzi1t0yPTCMdNNgBUNNa7HnvshncmZbdbQGPh7tTkMtDCvgeX25PWLU
dSvb9mapCnVe12DTWJ0iqzFL2h2NmjH/gfmr4y7P/FFiNbR6wuCWRJ0XzlUDfYq1
0n5XDcbWda/mS4dUyrcHOmYxj5OAumQVzUcY31DS5z4N8kYhz9HjgSSR4n+kdMS4
OokAx2cvxt1hx9ytF3oOgrDWAhcKFdj+AMpfFYHeJSGTk7Bor7B1rwBWs/tPvozM
1IvGxiyItn033gBgmj0McEisQQyCyo9RdT7efp/j+x5g84ggwAP6GQg5/FyaYSlV
pL7kM+rzdHkdBG+P4mb+QEyUbjWUMMWvXoU6dJNfCl41xoNSY4DZPeIJxtzyXcx1
xqsibVWkxgISbh952wfO0XsxLPEIgRbvNbqgA+POudrPUvaa/67gji94psQYGA1P
DnHRbQuShVq5wOfTBIDcLTBKuB31tVjCUW46tCcG919eHq8K8WYyFwt7L7V3oXmK
to2PQ3X5FpBjYddMIxhW1tundyKM91+PEcCqHBuscV4u8fPOD9OzSvzjS1zTxoWB
bEHpEaHdMhQ9GUszMxzRRajiTW74i07sxPBZSKirA4SCxcck2C7KsWt8DJUBwiV7
POOH1VLWD/Npblf5/RotAOI0MSq7tcEuDekiNih5/QwonY2cmDNwR5YeHH9lwSpv
qXMdT/Emn6Ah7mQdd5ZpcL3vQooChRANewrhL/nu+QuCbkNFnentDC56mvqKm/kz
ZTJCwZnpXb2OK2Bf1XQEJZiChOKsYq4V3T8cjMqCoLs6X8nvzN5RQxhfI4g8SZwp
mJ9MhqHlqnhz5Rw3aFD13h4z8KYoajCGPTdGh4hubDlr79BkZQpVDJC1f/x6BZ4b
6EkfiqfZJAfntnpL5OFctPNaBAdSAwzwQYtDjXyFSICkpDkmsE9SBg2UJbfu7IYS
Dwfrphvs4sPrqfuB6PJHB3Mcuj3Vr4PMdSbNy22ocZ4d0RPEzZfP8PqXW4pHI3jc
5R2ykypYoYBZjFLLuQ3OvsA7/4/KWJ01oqZdSD0TZQsEnzJPQyuLCqGcjIu3y9Aa
OVjeETuEOZ56F5QD1Vje/uTa7fFAV4SL9XVtZx+kyzltVO6cj8gVmA0SkzVM2WKO
K6v4sNNjxU7JgPhkyXZe3q3gn5C6K6QVCj9PguVnUW9JDPzrkzGt+nylbImAsyJM
bAGHTN+dC0Of3lL0zjQwR+WCWdvUfRb1gl6msTzcZSSSg9vxUtPisbEz4yoSZ8Oh
1Y5iGCvYjTlgsdnNdMR8TGIiUAoewUUlfaFdNDEzWHZTT1KzsbHuEaTFSCCbjS3F
JMOFmJ/P/987Ywat4w5imiWtmKUmvf5oDgaRlnDhdP2QpdQJyXeh/jRv1y4DJvGy
6VRr1pOwiTWYaIUX7TkJrh7mBUKBILQSXgli9qVAXPQRxdlxt56smvsFIz7wBB/B
V99C5udH6Nx+3BMMgKJVKSDnF7ZK6FNZdQB26qSjTPiJxLDk/KErpaVUCeH00xbQ
sDxkSNqtEV0bJYKNgH72VhzLcGoe9PrvukcHdhukJUuhFzkYeNYnwYmuV+ktyc0w
oO2Fmma0AqyfaVsH/5wb89lDAHpYHeM9+gQCQfiOykwnv1vD2RGtO7ZZRysIghH3
60VDDIifb+fKoYtrELMGZftWLEzM0Cq4LUKR0lXF5n6DPRS3oneH3p/bSE8+ZIak
BfvpxX7jtjaPi86oKl8HrK9BtMNysT1CBa9yn56kdcuXdfoK098MeFxt29AbJ3La
Ou7q74X41wUhnmPxym4sE30KUuB7lGFzF4UIQ1e0BpVOPYYzfaKhqhW6uogG/8RQ
WSXquoi5x9sYlp7eplOl+9LkQROM60m2TOQAI4NfxSbZv0YMdeoftFF826sZxQ5w
1r+RXO3btscXyNUljMTzELE9lp0K8fMOAiS/uO2j8T1xAWwonVeCrex9ey1cV1VL
qKNjJKXDmzznG62I4OruUZjw55N2dtDPsk3nyRnj7KPjs3+ayNk3OIl/Dyzv2Jct
nbNuMx+vE1tprJzky3szTP+R2nIsyYXjPOCviGAxgpi3BFyOjQfYLiAOFfLMFGsN
SpPTbI6gj+DViGqN5RygB1D0Hmr8BFHDRQnTKmxwDIz1fPsWDINN6A3Vm2Xjy9DU
H57tr9TB+xMNKdHF5cr9HVpkRpwzpxNAMSITzbfBXXjnAwWV5b0DlvO3Dax4vzFN
IFfD38w+n1gids6ebl+uPIgUVgfr1nQ69v6EkQIpLvaiHgvQH9UakqJMpbehJ56J
JrN9Al/8v7SguyoNukGAXj+ifXcbfwKXzacpYdUIA2VieQXkRe2MUsYX/eHzeDcX
IbxiiUh9sPz0mdV1o24lsDX36wws/pkH+hFI68PoCnDnoslYYg3Vozms+AT4vAdK
go8tkSgqgYCtXzMybDkylfwbjaHATTV4TsloGsnxO/2dEupDXVhevR+FdJF3Xqur
Z+52WP7eVI4towaaKH6fmeXQ/ck1SwZtMZuUelEpt5XYM8dxeXJ74r9/G64kEY6P
HbTOyUeMlBfZg2r0k3AIt9OM/HoU4Uzq2L/B39miHJqQ0oqbG1r10nS546Q/8U+T
swNLNz2SDi3TdkYVJE49l93gbZCV7uQlGkXJfZM9Y25OSQhNUXTDHQ04Ooe2bgai
xdi2j46B7xNEUicb/+mJ2zZ/WSGElqdwFZXLu5wlV8Ol1dRSx7fBIBqpR1IMoOjb
6k8z9mIDLTnVjjxM2HV82sRRNjCMq0F9SKgE+TUw5RGnz59WXMQhrRbRc5k5DgFJ
FjUw7wtWV0McxaaJCz5RUUUWRUrG2Cd48Ku9+37atQqJ9gLp5MHuGpsLsgWUH3YK
WbZsDL/ReZBaDcNbOvLRilePt0NYCDE+J+8yDTR0hEKg+yGsmcBY7mOAzxImxGi7
t1Ulffsu9Go0Xqo8qxD9hx0jRml9VvTAOmi/mu5B4ke+MjR6fGjq1FyzOwtwCeY3
aKHXicTIAT/vd7cVPBLf3O3nER6uWnUrEgjok0oqNPZOTz5exMnLOGCyzQQ9Gh+Y
CovPXJ/d8c0TOGklVzUqvFb5zLgngQQgnMljGLI3d/OKPhQDh63TEl5jBsDMzL/r
Gzb1R5LH8JrOy2i/a8wCTbdlsLTbGudHIv+e+QhT9P1KPTA4uC3JaLPhba2ElIMT
Fb7FewV90yinWq6Ceetp0MpG1bCjZzxgvJ1upXDwL+v8WJCt8qhUAKSB34dWnKWN
CB/9MGU/JWdO1W11MB8TXcJNIwyvoytuGMndzxbrUWMP8ezyUiLqLnziE1UEq/7q
Oop2gd3EvVxVeP6uXNY3r7fhfI6cS6lebyO0AA5lHtK/mdbLpy06HeEEIi83Jixu
wai0O5Cyul+j2ZuztNxFRXtyE0wNMK1zKp+TWJ0OuzBYJ+4dIc4vWKGJz5ijtYQk
2dHSj+slvFq8YrqCLWiwcps75EQx3Aiy+kI0KJT+h5k7JA/34c7a3Z+ddSwjrHUY
fQJXn7ojthZ7bLvJ6PYE/AaBcqR980DBezsQa/M1FGsDbs1tHYexKii9sCix+Ihe
9KcKjXL/x1+7XjVucYXHvQNsw45Y8gQrmheG36lsU9hRm7a+l+imK3pwqbmLUDrL
usqpB9hJh9ojqx0lGD4ASvPuAoIgJnTklvWatnzM9vmlUWPVWnQ31VzXsK0iyFo1
3n6NxPpLrUOWVRIt8hH2tg98CEHLxtq06QkP84x+Rj6B80+PS+zEYejLyxXnzhqd
nC9AURNljRfQBknwcUqsHTQR+tg5tTIuCGFN71+AuqKBIcOuNh+8cfaTCf8ZJ/a1
FhLcftfkrWDlqojC/wIMGxde1Y/GFEwTfV5ldJtZ14vwHMuQ+uc0v7yk66J8DCQi
qwsjjc/GVe50CJvxFw524WKRG9AIxEYWxlUAFLfiPC+B14YbZ9a+ixjDpBSvozGU
WS0ikX0Q8btx8s5BxStUaecNtBEBy8yR7eot1XlS+/RBh8UuMYfggJIB95fZknYm
j0EJxP2liwlJFv8NBfr/pb/njMKyUseC/EWg0Ek2Giy0hgsbSQ1Jk7y6h9sY9dW9
8bE2Dco+VcPa1QZgaERSO9MCN8fbTlLSFjmew+cXh6DiXZsajpP+Z8dAVTnFDmy2
Iv8mViZZfmgLzv9M+XxynAumZyYtHgE4mJ6EUf2N30uzPYX+8fZB6DJc/rknMLyQ
v/LU7tkObWylYzBUIT3jU6CHJO9P7zkvq8BsnpJA4zcUYGM3T2ZcUY3OAh7LqB2D
PAlUbfFsGltrVnSsmwLhsBBoUWRrSundoTRVOtg7SNfeygsI1PTHgaYWI0nPT4ui
tsaEHYGldqxOSeF80oxrlGKl99w1nDFXtFgw1YXgLdHRs/PUkTO/vp7oT1BNLCK3
MCg9Wih6G7MQMmQVHbstCeWQW3vi0LfkXuf7f5yvb+MTPpCh8I1AC2gKaQrdOKJK
SWlmNXw37mSbB4+8RRHu0cPLsVIfI/qYHkOD1w1hQBZZ86lNg2UQdw3tKPopFj7b
ngPf86lNULS8dNfA97AeMVZ8B3xmbhDGIigSoMwfVrSgLw6gODDMCQh23F3h0mqg
tEq5Pj+gzMBWMVHVbEuthhxnDiJd4p/XkINpfvmFeL6s8btKoblezaaiQQdHW7HF
WSsBbBcEOGgIAkZmLczEf6Jh69pyE50I/BCKx8ZTJ7dPDmDM3Wdsm6Y/5BgTNFBU
q+mb7yphUo39I9L9fe8vBYcRgIUFG0Jnf67qavd09w+3rDSbH0eh69FCK6FT7cJV
QMAMhMUUAbJLJma+YWjzbhjYjhNGRmuyazVwalhCbVZbT0pzN53AiIhT9YK0arsZ
ikyxB8ye+//NlS1HXlgRfp41uAL9Z5+9HmlWKMlEIGVIxHMx1DgRU2oLLjw2Ml5I
3Nns2Yq+ZmMUoOFhMykXCn8TxQt3TEzKRrl9pVMOPqNZuW9zfK8PsWJRnafJjVNg
jK0WKbgvgsf9ObzpvmBfBhDRlMypaO3pHzDm0B50LxZuU2MJaaejrpZZco8+DZc5
V3Dzn5vH1B3MPz1Yl1A0J8SKEfW1i1iw4j2nZG94eIpItR84xeg3097jI/ISDRNf
Y79lepGDC9TicGgM5qNEeQRjOp/ZxD1mfxGu/Xzr1FY0AGtRdyP+a7msTOjudTse
GEGz+AFtpK8369MQUqqAQxoGU4Ut0R7huV8v0qjbRgsp/dGD2MtqjZjTDsCuAYuW
ZzVWmNljEsJ9HVB9c6swSoY7oOtWt2ehsjpX6R+cxTzyZdizKGw/2e6YQYAL+gz+
Kdo539sPgpeq37IXrZcBQLFZa11AQvaOkqzOUEhEP5XPxtf0Kt/pLy5Mwuefx2gC
aStpjfLfDcMcK+94ua5INN7z0wrwU2Ifg37DKzwbf2SP0H8dSwRMfrfa03IrNYcv
Api6qYjCyiur7sLpsICx7g==
`protect END_PROTECTED
