`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lElEaCffiDae1GzLeHWdSGabeV7JEgyX3VaB6QM8fAaQn0kPb2TKXoImpN1m5tgA
NkVa/ArlVR3VjszvTdB2U3nXZzw02iFHQJ5e8NSi3Zosc1h9ssdipo95w/F+mwtz
AsI2X4h7/eBizNyp4I4hS0+N8nXdnIQltcJppxAOkIPPOuMoh+pSA3XUXw77hM4N
cyaGr4rejj/ZGK6riAinpyEQhGQXonl3I1gL+WUfjplAtR+AQVH9rWl76m+TOhcd
o2VcJDCRxZawxdVQUWBEj1q4CibtxS6duRLHEeD45Oz7wfNIAuq3r+9Z2mJZJ05I
fSdRRq63u/QZql9wu5JcKdr/+XzTmsWDUhFqoJQFRpr2h8XBlTwPetwaNOzDPHIL
UlhW52Q4s1nww06B+jy9m0MbloSQ5ql3ayAY7+C5Px6/VAuJDeUIUwJPSKBa/MqW
687ZSgWuu4RUAw8y5KPwce/yL0AeXz5f/WEnPxg0gb7RRsidPRp+FXnEYv8Zaumd
+A5ITXnJ6iIGvZaZu2QSKDSPEA6HNayQFyCYKFZprjIMCgQbogdktBebDF4F4Uti
n9o29D2iAvfIE2lwVXCS9yJVRzTadqddtV7eMt5ufdEeAJkRPD6Yym5o2ZMi6ILq
/fe69IpuVxSiveziPlJspmLk4jm1H+iQ6C8POL7ZFujiPoww/U6KO+S6QqnF7P5w
3NXaIImvPXGbFbCuycbq1V0WyIdssm3OrHP7iRLZuu2+O2uCqG1TtfvtxZRTn2xJ
BrVDLk09WFq6KoepRPjHrFX8Kz0a+HMGPFvnPxoT+UgLZZBGB8jvkiCwiLStupGh
g1u5l2SKWs3zSQyHk+8W14YmuyVQN/PM0AFm6wSjB+HZRvqlgWmX5tnJGMsGcM8W
5wMeJoUyFt38mq83v/qO6HETATCKFwFQdShhKL0xyQs4Brqv5hcc10uCLtcPD1Rn
Lu3rrqA0D595FMi7sXJf4To0b1r4KdAASD/t6+j7TwFF8EkCiOqQzytWTd14RbkF
cAsdsPN4XOzuqXF2Y13jLRUnWx9wQM6qKJD/Hx4OYqETHCZOhbI4CAmeIEC/v3/t
lgvvFw9fvDq8kuovPYGmE0DdXKo6xgFD0gXQHpnHxWEiDwQssHNvSne1vgioPXa+
IEiOoAY9QX0BBx49N6FVkZQhoBrcwZi0rfFgArCFmnxH5JfP2BetArZJ8l0M+ETn
pldDeOSbCPPK2FYUw+1naPV7H7yl2rm2MYBaH8ApHE4J0bG6VDl7Pfw1gTxnvPs+
ak1O/rF2Xu0btVkEvlH4i+x5Duy8GNCq58UJcvypWw3++9ESo55xhSAnJO2BOKAO
X1Dz28BcpTRn0oSx32Cl6NT8KU0TB1GJntoIgo8Y+SjI+DEh0H+eU020x/Dfc0mM
LuY44LNGuXsVeCCidA164s0e1hz+qThcdYm5YPj/QA0MQ8snk7i0QKOytxEEMkHT
WEYoIM13a2nqGcbSyiYBCF0i5TsY695tjkbMdZUE1EH0pR4aTgkJ0VtpclJv+aTK
C9YzzU1+Po2lRkYqmNx/0ApsFHrIRlO69CtTClkPTou4PoXktiuBh5Z/NSl4lkmH
h5/9n9n3h/+rF/NTHjashwjNPLzR0MnI7eBQ6gYhY7X/YBMe4h7aUb6+dyMcr+Aq
xxow3c4f7jJbii0LYLk/xX/Y3RI1aIsVp+mJ/k/c+S3Sf96Ze4LYE4Aw24tmaz4r
`protect END_PROTECTED
