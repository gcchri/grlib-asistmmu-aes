`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C1Y9jyzP1PVIF1BYSRdyi5OaA6msgkam5Na4EIa9QeEBHX9b/Qg/ws5vRC8vxIgU
cg7jKEJmg2ZJ6AQbg1pcWxB+1jQBCk5DbcxwnSIYrsSI2SC5M7BEHIuo7QV6PxL9
0Bx2UkDH7zoXFytD8Nms+oyxKOBIOcNmomlU/qolSIKEmEPl4FDCW22FXyLbxDRo
i/u+umIjFAws80PqqwyRKdLvbRrfaXANauKrAwsASFzFObLVOjZqtU4IGdlZ3zq9
LV5lRvCmPGIkjjVIemPluQR0cjE7CEQo0IKSPjnw8zL/n66rNstttX/6QQvguXpg
LrRu+bgGQv3zbQOpPstqYCfSUOnj/O1O1aVjBtLPzDzyjwOGa/EzKwO4CQbb3B6I
egFz8lz/RYLNL0dIX6dsYyzfSGAkvjjZke07qfeyV2REyk+kXQI/OyH51kKU6Iik
rh3UZv29ZNG4jGbHKvkw6e+ghHV/bAx30jGgHGxQd379V+/UUPUmPEk4UE8tKDpp
+nY4Qlxq60loKAJyOKRqx6uwOmiB/RMbj+kyhA+21L/dpm/P1fIZFeM0a38EAbH2
vergnNTi7CBGGKhlOz+O2tQJK5Rc9FaqUBu0JgmFl6TwfcBo+odp/HB0FObdzZpb
LfbNfc3CiXg6LGU8j/uYIOYGFmYjGI3sIfF19oeoJtRgRfMZgIzoKGjOXtR5UVrP
Jk+WRNTKy3L/t4dZghnOTT5c4SaTBEPijw9Z1ApTcpfwnKBqR5UHt3N9ig9f0rTR
xHtJy43majQJXdVyjyN7EA1CnktASD/y/pWv/5ttP+AqfnEFH1hinMPlE+Ex6FFX
TvCVRbzsVXlq3HaOjGxhUtACZtV8BWgbX6n04rFlGSp81KFpgMTn3Shb0UXOgmJj
xGvFQsC69xzcgZPBafD1z8tw8TH1JalfygoCZCCOq3sUkFN/X8gqWbH9X8swtgPe
5JKLMBFvK98pFn2gNPpeuwz2ps+YyZg6ufBjcmG0Rnw=
`protect END_PROTECTED
