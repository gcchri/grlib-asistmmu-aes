`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2GcTEzDbMcxK2DbqTpCPNjeGeKl3WuSlRusFgkAV0Bkmh858+1nXSVIG4NC3w0LN
7Q2ETA5D5v0OtRAFbbw22B89/MEfBggxBi+lCns68atPhgRUflZTTaKwAiK8AZr7
58Em0ToGgkKDWgpXPSDaDDo+wkf+c4HK3pP55lJA2evAa6snYc5zdGKWHbaorV8v
sXdRhzX/ISnP8KL0zmlGKjSZHwogRfZtxJuVZNZSKMui64w41YG3mvc9vdqDLtcE
b0JxAE1pCvO8tRwLeQlWsVO8bzT087RAFJDS2oTKNPUxoJk3LJ4N9PiLmQ0LLzeQ
Ml8oLuBonSrDLsXoCl/O1AfSpIQ4qXSrf5YqOptG9wy/rqztWfB1+FWJ6epa/HKV
VxOCDlPYdYnKkOC/NGea1/m3AGyOIZAWeDVxBaqItPQNsRDknHDr4EljXVD1r7wn
YTXwmGaZs54SNHkotEPveUOUmN+Fd0sdgrwTK/2a/v9wnMupbq8Xf8DPXAcXjs0X
`protect END_PROTECTED
