`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILH9DsXYlhJnzmiqnxv3AxdQVtd2baRcx9r29EhMmx1ObhR3sSxH2LInB0np7JOw
ZrAws/WqQhufaHvgL2gVXAP2Gf86jXMNhE9vjsOLVym+7O2ySCKCIv/IHyjyCSc2
NS/+64d7UKx7dImILHl2w0CnFLl3UsTKqapUTY+n/qYLqnNWxe0ftbLRY6Kpu+ZP
3fnqHI/3YUB3E8xxuvHAKbNwSJ7L0dIA2FZtoQIMk6WHX4x/Y10DcWl7cYD8nOpG
EfHuSEBhA/V7eKeXKRvwSsMr7XZdmx3xi2WWj343VEHtjb9Q89BpUj59JWgJSSlZ
MCKD85izxnZvlHtxheR+imYMiMy5WNyadkTqIskeaionvydZg0weJembVOohPdvD
uEgykmDe+lUqp5/u1fO3RQdZ+ogoyAWe5AT1p/1C/lM=
`protect END_PROTECTED
