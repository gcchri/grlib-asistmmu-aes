`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jB3OYFRBF6h/t1r2bsYNqQapVpeZybuYtkOyYQBUIeyfbD9r/lScc/LBCf8p7Kq9
FItgn9vVwBqClzTu5HQEDzMweufJAkqZFnJ011aFYm1cC82GRdGygr24rrTmC60U
qCSu9Pk89DWKT2zhqxWvRKzAJ7Vy5PbZg0Z+TOJbeIYZalPweq5a0Bo8c1aZOWlG
WmsHerDD+oZLAHrmtpWBDUymHDxONOt17wPlCoBnXR0F9KV/pRxcB8ia0A5i1jAh
uHeS8xZil9c43B2/WNUYfz5dPU5rLOKaZr7P1n42QBHhQST2VhsGKRb7eEdPcD5q
xrrDIF7xwX7VNwyyIQqgeiTU4DlcApPdgCEX8GhZGzxvjX70MWk2xqgYdRqMCdT5
AWBT6PAxWjTMHyZTHFBOr7B2vS68YzeDoAUfIODvtYZtTAqsBwwyYe5E15fQN0Mx
gmNw9UfUFuHKHcEPcMdD0shLnmRWR2WI0f4OV2Auck1PnKWZJbVU1MRX4tfI02FP
H6oNic300qHhdnLwfXlfxS2twj71eAos/DVMpDUSvRhHhiXwpuFhWRYT9OLIoXvg
PLSnWIVKQc0zrn6h6fInWFYoDQRQKB1y44cWNab1huksiVv0foUzGWIR8UKdkCnK
/dSxGSGnKD8+fwLIlUsOsIM51Cx10jSO8Epyp4Lp0JIA9RV66pPyAvWjKPniixY0
DSJGAm6luBuk0WjHETaPQJWS/CS5ICsaNuds2W7+ELWTOyda9e2azJ9XXEq8tAuL
bY8u9pv2MSAwKbu7rLVCTvMQ6x0nNmg650p6ZHU11lNBcT9DaWYtb0YG464WGaAw
8VrOKxZjOJfN4atJ0VOssIfq/nGschK2wVv2QEUuCPQw8pw1ZLLe0BhjCZTXj2Xl
hSBo0Z1M9QXbK3QT6Z9kw9XXoonF0TIXcL0Pt41UObcW2rEOTboCsbLD64pU+GQ4
jFJ6zBMyNPrxqyGXH0wnNvyagHgvnomFityLZFPXAL9VautqEcAm18pGgcpJ2RaO
CN/UBSjkgLDZdKTJeruD0AVksVcKl6F2QNvuK7R2jxVeT2h7wizzM+i0sKzJgzMK
qEjEDy3Fw22rad51cyIqtIKnjh8cp0qTdaZrrU329KtuPHR/pi1XLIF+Nhz5lgPs
NqYlT1nJEySZ3aQHFqwf7jBJ8+cAhaQMqr0s4paLlEpNfNAWwdesYfahdIs+NnYD
D6pBoXljIfivzPtJzZo72yXXeuek/GMdZNq4DN0ZWvYjMaIz0rqqdds3jtYfdsUa
YYLaWFTEm+TmU8wQY7irEQrunFPUHjGPs6WUoYa1Y2qgPaEl8IvEj5Kf9zhHpqAa
FtYlkY59UWK7Cwr2GoLemgCOSx+btavIOjfLCqqGtJxgPCAB3tT2IEVVLmjBzKt2
GCzyAYYbdVHfafE8NYyEyFLLduGRFFKT0qnglfVRKSKh7o7XC88k5qluZ8DiqwRo
1Dj9ZPpbXS4KC9ebkTxA81Sp0Op+2FIiuhzaS+WqjrhiwAnB3tYlYoyY61L6qJWH
Uy8yrb39RRLhAgyrNW/cv+wV1pHvODpj8AyriB9PFjfSwZiW2ql1Q5mqyEHFt/tH
C8zsSerPJlm2BHKOW9ineJnVRS11+TeEwtyS/q+GicwQDAzGei7Nv8d5BKYixCBJ
j9syzN2RY5weSnJEAiZ7Rq+6nWONmGoWeQDRbqdWkuf9iEyeUPN5MbCLasvfwt20
Uh20ozi19YxZKoLHy2KJ2KfQnz4jmWLtdxQgzSw/hMr2SNv1lrjsUXRqKkrCCv0a
8DVYmNcfx7NTbLt5dzo/dUSuHsWP0Vibi6WyC20yLtTTFYKWUJopPKaKQL3m6Pg0
p7sYBF3GOg3940F/zt577nbXjYvk8X1WixMY7Tqbwg7PXI2KM0G3qUjgRD1ioCDu
S8UFl3n0w/9kzSNIMS3YCVLqZdnhOx8J13DUIv+WL1xT+cV6TPmuIZcVtx80UXHj
iXbAkZxYZUHgsRS1lF+mOjUGV4P1sdGG6oexuHDCSTnX4EQlsOQoAnjB+s0oN3lO
bMHDmXCNMshYsU8yA2TuJtVptJ2bRWuWAcbdAy27FWIGV4uR78HkLVdr86ol+an3
ZYBR2w3FlPldyBuYVwMK99wDdk7vMk5ZL7i0foNavaJo9agW6mXX30zn0bb7R9Ip
xFMb9qOT6502dYJHI6pEs/BW/N4+v9PzqH5WiNFZ+gr+OwyAYIbNdz2mg6kxkc01
2DlHlSKeAQk4HWbNLDnKBVRfE3DwtNBxHcf2oeMA/JSrzrCiZ91hoduniZHCdImm
tz/2tT7fjwkXuTQlJg/jRPaISyt8G2MxqNWcTbbapXe6M88CA8t3+XDM0JztKzys
Cnl2+W++mmCmcMG5E8ADG+Ii2dOUYW+9wvuj380da6SjXhoMIUMKir5pxvZleo0T
I0Y6SIycBtC08fTjpGd1VQ==
`protect END_PROTECTED
