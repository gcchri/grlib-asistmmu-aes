`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DNhVi0OzEmvf/XrBFg53BygFplKAfya2KBF3dKeM+btsRKmb/XNdtWFQ6n/nTjvZ
SwLRSookSp4T/ZxTBNlCAnXogJCkc3XfRsZN9v4Mmt8yXp6xXzx45NrqjHZk1p7c
C9Do9ZGTm1DGSJUn7/Dg/yFHkRyyd3pmldhq/4ZyHS7xGTEWumHMkegSEs68uKaT
32hsj5zlmCLCkczr41qLpQ2h1AXNbwujuynCD0v4+OdJc440L0nEmm2r93ugBdng
r+eNsndNP4R5xFhGdtysAfixocB6F4F+7+yuHx4yZTJbeqZNfDvi6GbYl/ybtpIn
be+LjqAgcpPmbAnqW6HdS3BV+MJ2XrNaIV30gIYACiaQyLxxNg5mHOW3dFwRpRQA
Z9IvpctMsKwilfZut1QwQw==
`protect END_PROTECTED
