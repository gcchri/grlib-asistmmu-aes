`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfu2c4dbU84TdKEgRaBg6hCf7/kYT8Id7MKNxdG5bjfOyUZdiJAHzawX9+ZYwMn0
NwHtxhHY1pmSwddDkyi9j1OgZ3sQyxvVXMjxRteXN2nbYaGY92QjotUMm83UqU4W
YWzJ4vw9dRvdPgtmzP+zlOijAZvS3Z7u+hy54MaSeSou3ejblS/pwafas0zlmtUN
I+UUq/Y3oNsw2DGwD8RolZL4j6z0vyAlfPEmPFzUubtbe7otdq4jipCBWu0ZS7ru
mOTFpkTmg2OFWVxip0pQkCccqTe3uKtjRHq4ffA6wroc7796gD5BxCUjYHD23Ax0
xTwk4E2HnPxBOoZkk4Zape40eGUc7jR4Vt+uqxTEStI21fa1Mb6RgAjvOWoufqLP
bCB5HHX6+NtV3ZyIixQnfGGnY0xW9TKX6jWOdVzujaRt8O3BXl76a7AM93ImDjsE
+VQ8XVk/EwBdxGNLz2n/yVEqcj5QO849fplanPem8OXR5S6Q2LyOJldl5GHN9d6q
M7jcSfZ2gB5VdarlkXRLJi4fsef31Ea6Metjhqag+TUJ1uXYJbYNUGN75Kd+vcD8
BKxId0nUER244D+DvMrrjCfiGA9mLxy09GwW4pcYr+tMDZIOYBybSMJYbZOqK/dd
49sE87fPnQScR/RnuZAlNpGq6ylCDEVAZtLaDiB71P1+2w0S6i3KYPe1iIae/Em6
mK9NDMJlQp8GogFwlcxmi8Gt9yxQ9/ZTozd4KC2+F3Y5sRh3t7dMhelyeXM2LMDY
JBSu8r4IKKd5SNJtILfnLvUq63DpXAJrbduEvOXOFR+Wo0WVgF/RhZvp2uletwHv
PfsZX9CufbDAUqoF3RXc9ujePm8BMmWEOk2cZLKbIrxJDxO/ThaO0+sHs3Obeldb
gedClqIw4D+pJweqVxf7CtqaINk3yJlNeJP5bD6FxUz88i8zUta2pDSL9yZ97Ghq
`protect END_PROTECTED
