`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8tsXknvXXsFeagN+L+cXpwh8NUiRo9tSgQ1QDEwiRgeSV5FcMRS4fqV43M1WXOF
oY2V9xz+md0+AmkqKtjZ8QPj9IZYPa6n7IufW0Lt57/eUEbkGltw1m7RoHwciP7A
bl90lvmbp8pitty+xwLGx1DsLnvuclZ5/4H0P3jjilRSMXCIBeGcDCy5WMuxvSt1
hoTFavvl2RUhXrGIAcgzfX+noekiGCVs3yE0nB+uXro2aI7A9T7owI216NIdbClq
0GOmj8TVUYcB1sLG6Sue44I1z9hnvhHWZBVlELX/A3JjoLBYBnuXHOG/MIW44Jhd
ydQq3pkXJU0NsrK/Tv2LRQoQ8YLja/oy0hjz4KcLGQPSAgUZtQO1IcCWDQQGAu1s
b5jlCqYseIRU+QvW3sHqch5B+5htzqr69mFwTwsPlMxyTAY7peiKH0ohNoY28Cwk
IVTrRbetyYBeZ8WL41idu2WlPU5qUwKETjdFzAdIPoYUxwzVyy1v4pMAxMNG3GFR
`protect END_PROTECTED
