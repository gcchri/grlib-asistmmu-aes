`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+94/I5HMekNprDGXm6cCcJVaI1P/ICBYKMIR5VIOvI0BnhCqamOlZF/PhDv9bVWc
c1RGwPJyDDf3+ckgH5/Zv6A4RmQN9Mjt3kszySlZv4VNp5/gAmMejElrN2MTlV8N
v/T4HkZgCIhUWZrQvAOQ8M6+5fzqflhfJeChKmkx6b2idbIoT9+5hksgBfJLSktj
hLFBPEsQlidn7PZfna2ozdCU1jaRmvF/25X+vLxLOoX6ngeSJC+OlN63vZe1jRXM
Csw1x0Gir2yolnEqdIrXWQ==
`protect END_PROTECTED
