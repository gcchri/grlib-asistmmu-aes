`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ezLI/H3Y6U2MENburqjPMqYzKGMA0sFxNA2Vi+w9ex1D8Pzg3voaT2VexEoBlu5S
rKa+ywYnBbEdKOdiEKnXp9vUBhMslo7MiGXjgJILGlrANrAqjimxvDzqR3Umj8ks
8eQybXCqPfk3WjeAuBUnEg9PwnvkF+QHYEN9CT7lPecdobrxzTYyiKPMsUFlYrlW
2ED4UXH2ZwJc0CZ/GH7ZPBFo7lHpUR7zn62yI2aMi3UMqm4J7bgN3FAuEmeQMhjA
7PqOGkEts7kqU3x3yX5rzclOJFbOZhiaGCEKSIMsK1Q/Wacf9dXg9bCPsh9J6nb4
ervD0bGD3P/ozwZyC1KFP7sV5weDr1V1+ZOuihfzkD6BPpXsd2BRL++7shgAI11l
`protect END_PROTECTED
