`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMiCWlyXH6ap4SV5+I4PoBfTm3g4B6MoLmiO/5q3EeyjaOTCmi8e8xTCKe365nMR
OBm9GO7AJC383ldSO8EsTNyzcWRG4mrnhdCzWW0cGApxoga7X30IPBQo/NRXhiSc
vKlOi++zH9x5R6YMa7Ez3JeSt1B5oS2EyfSUCUCh7n9P+5pbSS4NKJqeefOk8HNB
Si9dD/OmsQ46VYg7NxVUNjt9hZVJ1bw/bDryHh/qFrgB8WR7dqW+6m5p/MinJ1Z9
xIBBNXrLyOA5u62ArOiUC5NvmZ+IZnbmVVRofaMwoQy7aLSGmDvOULAS/ViMAkXP
iPMmZCdLIwBTskICvHg0s8ulay+tvFQh5cEXnT8omJnzoQVYsEAHKSbGr1CMe8xB
Ezk/OVRIMZ4fUrennU93gA==
`protect END_PROTECTED
