`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wZrhBpKE4jykiAXvv5kX6rjKq4FVVB1mt9IMKuz7r92O+GXdMeJ7bhKzYwnbySKQ
QqE5UFB4pwsy0wdlMRe+4eZ1LYnuJB6L0hgQkk/9k8Mh1pzCogcVYB6+OCwkxZqK
exd50au2gDs6xXyLKOOBUqiWAZ5+yVG+TD+xPDZpCbwKQ+MCIaImBtd+xEx2wgtv
f9emqSUFzM4FuVnC0IWCGsEmo/b0QXikR5prPmmCbnZBNZj+Li9Q9Xjz2KDDc5Oo
OTr986I8qZzpt++wMJ/z0arPpywERFNXw2ONLvB9n5dnb5yDHTNCCkrO2qY5a0Ku
gNiRyubMd7m/z/1kbKvJrhqE+xsG311OhgRGt9GxsbHcI75bC+TzgGbHvPGGU6Y0
`protect END_PROTECTED
