`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOKNdDAKCHK/1srXISsZ/wPsGZUAUkjohc+bLUme6fFgnT4u8viXqHNTQclCqHaw
8e7tba8LyqUfGpGCrze7fGAWGHf6s/NyeQ3V4YFeb/rL9U8m9P92VIfN9ozyac4w
EdPRgUCNO/dABUS+OL5fXwEN6H4M13vKM/niZanb/QxWxFeXSOJrC5lycO+h3aEd
eQPryOauNc9L7ywIF5gIYbho1LEoQyH1GPndD6F5pQ+W7lU/AJGGS2C3l0SwZacY
wdA1GrHB6fvFGKmZ0UdMDoQQIDyvlkIVzLQQOxH88cA4G+F2e9VtNqnt+j94TOo0
rYd32/bQ4kUwWlFTFThZbOXj9hAX+Q9Ok/tZ+Itnmrr/wshD3b2hMXE/aUue0O3L
zIrr6b176h2F4kwbpdwaQenVUeDQ4O7ns4x8saKJvn28gI0D/i5GiOmgdiaIuozN
QnqdbZnQUttrfjssxnMcFl5ROlelxTaWtC01dLiD3t0TrDL9/+0WfbGtEzPWCuP7
tVmH/A86ZLwJRP8z54aZQu/vTMP36nWZRhFvrXylt2pClzYFjxzYTRv6A1fJedd2
GSiUfdOIe+KRJSP4wkV3y94ugKurQMabKxE7ItkMM+/7dZaapzBIzp8xnh4bot03
knLunZPCd+K9Dj3jNS38c4Sn3nkDlLyFTM/XvX/W2NiMpVQs8Zsqt7TlGJOajHN3
/Ge+0IcD2yW1bme3h48iv8I9+QH/eDhn/gRbExsgmA9EWeiw++oaCqU6uDJCidEC
XtPPBuTNimTWRwMDXimsW4B4OX3O/XZMKHhd+jdbHlHaHrTYGneIUiTJZpoGvhnu
tt7HQrnnQjAE1sjnrgGZjJ6WTSfIOzMl3wX5p1caFPfysCGORIbj/oRfI6WLMfM/
Sjw0xAErdNWww2VbT4N77O70TbOWdSVk7ygP0FIAYUZ7v8OFbjY8jbTY+B8zZOG/
v5+ICmCe/MWuc0IWr1cGA7ZXFcZBISOpidFLQ0xm4bMqtqI3Z2672LEEcfQLsvR6
umBoB6lx+HgIAhjfGQoV+9K8H4p2ahRA80ULGYdXChNb5FVqYN5zrJqFyzLndJfE
vvRibvozLQOizLHhTH3BHwWZrs3lO69nJJvcInDX+FQ2+T0MMKldILfVATKP8akf
g8wEdvPbWUDA/ZwZNLWIr9eJRKNiGeyYy+WglBjT4/HIXO87xcfXaJMnHqfOjBj8
9biDlEHi8pH7AauEt9x0rqxtUJiM8nyO5prMkg7z2mK6NN+2d/mhioBzIAhJeWxQ
1AFTTZPDs8zOfEwnZv/aFYc7HaaRKHcvHRvRj6Q5F9H76OUTuTCOu+lzy2TSsO5J
Zc3mDdZ5+WRv+8kC2YlTOJtRkWSHe62N9Ztt/kfegQm7460/I+2CpZVp0NyjtvPo
UTtKMn5IvvT/rGfzqgEnKUoe+PF6P4/cO2hmHAq5A5LRqkU15WGWiC4T5EL5vFYO
AjJ3Lca5vXD5qm+VImN7WdGiTibgmU8G8qKKLqPFmSB0PKXyrYtgInRAfTWBSujz
tRa8OA0hZTs63XoEYaMAJdWsP5M6iWS6Il7OopKQgwlFnnUWjI307L5GbxU8Y6Mg
Q/+YOkLdCRQ6NzvW7aUHn0pqVUHg8tdNEFj5WxuLSJDbyRusIaiEcF5V5lCxL8ED
+kpzAI0ohNVGsBwq+hI20MJZYYxhZTcNyTgosm0Ok3n5fBtn29ZdOd6g1stHC+by
JLTTyuAEK7o+dBJbIX2D9s8zygkUWIg0ESSD90K1MJrCIMMO9tXOG5/lxdSnMP34
W2E4kwz1AMXhn4GEgAp6A34bGyMITbZ58tfA3scdLy+bxSv6HfNSVzbxAv7TUVgT
eUKB/626BJflIM7rBdqSCyglq6A0xVB3QGVYB+yebd6sv2VoR/UHCulURFIQwhVX
eqH/cfCSRW5p8X5U0+IiXRpO/uTj1NrbDbTtjxrohItHInyFbIV2m7fmoiR1W2ML
o0A+nBWYHd+GC7kPcLmRopGw05nv/WnmkWs5iBdfnCghk40DsYPcea31ESF0kPyD
UB/u+xaB5T5+4Vn/IF9V/uLQMuZYUgdiRPeDLnIPpAzT3DjEHfeNQmHAkNyp2C8E
+JZMqOneTMSqcf2NjMcU2BrIuHZ6BGEDfRkaZKWb+b/jrJ25FWpXPWVdN9YgC2Kr
pG4ptUGydm3sT4HwEMaDQwD3gmaDfB8sOeaiNKfqSLCEN96FxsRbcsf9AfkVZ6n1
FGB7LCvVc9PU+q7q/uj7er5CBYCSR6LErvFDqsX+Lw0gdUYnM+Seje+KpmBP3wrj
K7zIlfUvS6cDR3p/MTRvDGVPVoqrXhpHPFT+m7ogkBI5Yq/SA6F1tT5wYSklsPbw
NtWGv6/hKK2oTNA0AnLun8Sco7wqo+Q8DGjW+jtBLKHr60cNwGHUR3YkrRZ1hQeV
i1kfSQnWyBhyU4jDGFe9JnzBmpDaYpgfk9uzetv3aqsOeSa9KXylH2kyxNuZV2Vu
3BzrfQDZcRTPyPvQGxgbqTxeFPE+SfQdC7JLOypmcBYeAEcUY6zktAQiEHT/KphG
9VJtWFxCX/KW3W8xQ44xUbN/813QJ10GV+Rvrs9k1Jc3dY/b9R8xaMdr6K5nOw96
/knoLkQgO//MLq/EkHmlvxk+7sFfEE/25tIjKymjL+s9k0SHkYZ7dlexXE8uuXeq
t6IthHGKSGIb4lZvNsPreoF1O67T2RLRxdcjmVOaj+BnHR55Lk34BWJjQfrK0P5Y
QLkGkmex2ELKketekKbE48EOI9tPACzWOMeI4grfCAN3XX9xabUKWGxrfjkpg/8E
rTtC30j8eA8c6UN8YDIuaXKfzCctpB7mzC4rawYVG0w7W2Rj/OaAoLhNRstO8SDD
E0DPkSZvibp2cUaJSRveCZL+433lvuAUDwTZf4DW+qms8qzCYPho8P/DAyqTuYNG
Z+0XzAYBQorBuAWUUdGoTJpI7GJf9xNb2uQaQ4arQJVnTyYVktX82NOFzLKN6M/l
S4QRgOTU6SpuyKG5LPItvcAoBF1e8cVl1xpv4cSi6vpbJ1DceMBNQh6mvWSp2d5F
CHzZpNrxuJuy2OIRFUGsGr5Cn8b0chUG0luLrGduqZK/XCk3twD9joofu/jOt8Yj
6fBEvn8EGHaRtLv8VlaBaK2kDiK7avoa5qnXaFEvWiEPodpVjSy3kInZOKOzi0+k
BY68msEz3jYvzDeyeGA1xc9gjHMF0+0NtwmV8rBEAjzLj5cdNgo4uxL0jTviU8la
dea38LTH87YSJEVO3Z+culK4k9G4ee/BktxeVsSrjL5X1NA3vti9hcik2dBI+W6R
XpDgro2V4XlYXcbje2M7Ai7vcDw5mIi24WyU8F2/eX+NVhspBxpm0ysJLijI57ee
vhcHmFwf+7dPO9WOqq6RWQ==
`protect END_PROTECTED
