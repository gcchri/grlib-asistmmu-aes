`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eNPLuooyIbmO9stTYZzukA0IjKuwxtNAvU2Z51L+k542A/WOVtS6/b6Ym9gwd8E+
pZHGmi5iuG6TQ1kTgHG7wWi93owRQqogZKeKG3pymtCe1vBYzMEEhDUazbgTW6cv
b5R6lym/qKPUewv/APGolYJat4bycgHGxfVBpWZ1vJ4PDZXu7KzPyaXCYgdyOKmW
iIJ4GkHExnH/a7FFN5qAkOKTu41Pkd60VdPz7Kp9zSHNe51iB/W+bbsXVkUajGfy
9yMZegr2eRWgbvBE1cWwXvmG47pvblaeT32wj07Ld+iZcCa6AXTCNKfUQK36Grsv
y0Y49rpwoI0hHMiMPGMoKZpsQhcq03Zd8SZNy0Y1ZALwimsy0ZTzI7Krx0/+ST/H
0ymbuDZd7XyiWUPEc0bSlczJ2+0B9zNyc8rbV7DI4XW6xJX/5SKB3lfvhky1Jytw
MLdXK3hwUIgE4rBE2CuVZa2f7Ph7RozmKnU7VBV2R2KA2himDpvVSnMX16SFcGxP
671WZJQ3U8z7dmXCGNIEc0HntsBgxYcmsevfDnFPhPkS/+RhCzT1v+PqoxL78Wwg
oDIIWVlyP6OcUX9MiIFsiI0F9dKGWgdh66Oq8t7HrxsiNx1aYY5qnpkHJsboJd5I
i+bwswmuiprCnaBba5n5V/ZNZim4sutGMfDRsgVEBn8/bdVRhPs9MklX1vYs6FCN
OBkrwE/X3oByq5o+XfkQE+nCLODBQeheQSICyfFJpdzxPGCS4bXU9s0JTholTTIn
4lQiZr5l5FBP7WZt7LBcxEpi5sjg8HVYcrNxCz3PuQIpKDiSkpFHkZbLrjLSchjQ
sLBIZqrRrZM9tJLN65yWQrc8LzppwAvX9bMh8HctNYsGsepiDaElxyY8FcizjMqo
SyCgGC9q6cp4BkobiydlwMvVmVFH/HRBUJ9ocPdRg96Hx0hYwcdU/FQAWs7D4gJY
9QSWEv4cHLDSVIyUcKd1Q5804iL1hpG89+KeTseBcvmR/3QFVDLfcqVg6pjQg211
`protect END_PROTECTED
