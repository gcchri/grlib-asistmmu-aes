`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYz0XrO85HWsqlv6U/E/aVrjblMrQA/k11bSGmucYpsTEW3j0qUUZThcCHvB2VDl
tXvYN8mQebsMDqMmZM7J5fHZj28+TtMjNjYSJsVeHMGbb3re5+AVQi+sLbyseyoE
05/npVAem4VFR1CF5ONoS77TVNVHo37GHRP7V1TRb9B39xSokwNp8Q+owYvPG3rR
YGaVD1hJduHArGJTufWsJzAp2pipvS+1k5s+oI3JAkOPU0xEbHO753P5VCseXZYc
PZSufiEG3KOHeV4jAdMxq4NgWD6YARAHiM5Iy0+046eLhHxGN8eO4u9hlrCFODDy
5vTozscDYXPEmeu1mmi2DvbhZTEm8YJQ9rEfTS/+XeucX21S9dI25q9WnTaCccmF
lE0foHQTYn+qS/WaymJLkG7gEOegUZVKEjp9M6EnIt4ixS++vNlp9H3Byvwh2rif
b8WQROpJ9Ai9X1cldUXa8JrSPb5Ej1sPEGs2La3c9adNtQ6WoU6jGhMW9j3U9KAM
M+Jg26AVsQntSgiTrLNTdsfmupyss4OgM/aY4cDmtCv1T7IcMKuBKKG/yQTr3/+B
`protect END_PROTECTED
