`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+fip9RJNAPyrUOuMJAd2CDWPF4QjfnvpqvtdchwDAeqvRQ0P3/W6E879HgKBmy8
6Q85nIcdKYGlj/nbLJRC5W66ymoeypxy0B0Jq6eBo3iI70o2JQZtngotVl4ozMrf
5tY4hO+Y82QPRe4ZzERFrhF5JyEQSIv5srqsEikluI+2rh4ZDIQ9/3Cu9d8sfLMD
yHlPynnZDQNGJUDQKrdsk597EgbABAyv8bT7nuIwu0PK5zmU5GtFeueJ1kQkLSu8
Wky9bjWgC454Z6ioHS9NMG6haitGIaDf9J3aEXHaLK2PUMv9RqjiWX6PvDUiaS3+
RkPtSpEcvKH7HGbXhf5q7O8iCj5sXudO4ib9G0crmx73q39QMvMPOagiX/CQhKkx
M3xLS79npKH7RFUxv6tNskHD72ER2j9J+Ra46RbvcTmJjLZvMWWyqEG667bW3BUr
4zj8G+hz0JZuKfhGWdt5dkhluqPuMmmq6jICvMzj63T2BbtX2px2o5UBrdafyGrR
GAqYLwJoxIh+sDeWYpK6cOHEg8Qf6oR9RzaTIw9TK4nLTZqIPQdH7Qg1gbbpNR8n
WqaIRTj8EG5fTzXrSONjqN4yhPMI78gcWL2kjGQyWsTtqA7/TYoXgwFq9DST0JpJ
HKcR3pwfon/CHQPr2sDlsh8fTsm8Jfs+cqCRWv8DqYOJIlWOZfodkSi8BIkW2jwa
mKA1NtsmTMwnLCC+dN7MjkmWT77HQ78Qd5jUz36pbLtNhkOpYXCVxu5+MG4+EbE0
wEDLDWjOw6W825wiE99TVwgdzja1040KFnK+iA2Ep/c=
`protect END_PROTECTED
