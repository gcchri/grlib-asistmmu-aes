`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T1wRTKZFJBSLWjGtV9cnPyL+dqLoY3szyuoRTKd0z4fdw/H/CRMR7yDKaHKPCD08
po46XsXSjMwjTceEiS7GPY21qVcCtiNQxYF0hD4jcrUNGgaGYKyaTffni0GZS8ia
hD/ixOv+KuBJ6DYt0KhQS7weDYS/DeusWyvQjPjeyHNm0etmxSeBE+pI6r4W/Bhg
w5NcqpoCKQ4QTu7frl4dX3fVS4Qqx43vOyAQkaVNWYqXJWIWVWxmolQJzgdoEDY3
lNozxpc08NQlcgVvpSbkww==
`protect END_PROTECTED
