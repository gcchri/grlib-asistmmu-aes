`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ala0gEIFhw11OpsLVaA5uFLGWidozZvbRdupGQtXBKqucG9ApRqE1IyXkyeVZhln
YZrsxJzURhNOT0vtQEdL3Fdo+erYHXxzNidqegP+JlAQ6VAcsMjUiroAGVWXP/9F
Qp1ZlCnVQa51pri6Mi3Cr/5Msg9b1MwLtK9qdbsnERz7BqZB4dArkIKqrW9rKjGk
cw0++BKq9kSWVmXkh6Unm5vGAccXyclpi2tS11OySoIUNHzuTpdTxgEA+W0RHP9Z
zyNW9+9yovMyVzWgnmGRSg==
`protect END_PROTECTED
