`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eyu9Y/XrwG9mP5r584xq1MqMqjAvA9zTdOXNxrPsHFD34YHbR1zE0xQuY+H2RtA+
PR2b/e8ROZSx07LCNaDNyesGwQYUYvtX6JD8nxlMlg4ykL/uRbp8RxfUru/nJvKA
aqvwq1y3WI+SRuhNjRU9/0MkoSXtZJNJH3zWAqMbwx/3K2NduKX5yl8FpEy3f/A9
BdOhJzQwlM69Q8WMD2hjL/uumGmyaSIBmDg7Apq3FXgNB8PFKCcBtejI5gsU6yCy
WFOynrbTUbnLrHR7O+cQUGt2Jm9QiJ9tluyZRjSTYmBo8p7T5FGDax5z7Py5qG0w
OxiIi9p6SkH3+znxHWi7frsgGb4lS7lLEZvO2fkS/U3URFhDrEW5v9cMqc8nZQNs
nI9BmPf7J76j4soVw9aSey2Au6KF66L8iDx6Yw4lIkJCXQRdNNH13ud9w+41SgB5
WNVHDQ8xOX77oGfPpbREl/KRx44Hg9Qg/SGPx9ppKVkjScyLESmkK9chtH7k5mfn
NRyNr+Jk0R3ReZ2Pg00ARCZyDUBKHOm2G0eNMRni7AlQ7BJXG5fgdhhlcmknvuXj
j+hK2kMtXqhXzdNUd8FrrT72xO3iKmZwY0gVQA+vyv/r6JDTdDFX00ppTPTv0e27
bxA9fh8aAqAEYNG4J+bj1g==
`protect END_PROTECTED
