`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yaUdda6f/wDbylDmEK5Kq3jWHo7vz6A3FLIlWvI32/Nd8fIJDMhsrtpLWZtsQvhu
iPh0EkQSqUu5D3Jv9r0d5iaHK9SXjCyp+xwUuG+aIcYHR1urJPPyfU/9sSmczqM8
4wf4ednS6dHP7RIF75QZ8K6rsadAav/UHdhUryfiSQprNSFQ2caTciHjGt6hQolk
1ivGJcBWQ5rryvhIzKsgCQYSh2fNEvO+JWAzcur+85HxRB810a+dM4d9VMwZMzlP
sNTW1MmL4yp8jRwbgXHc+HPeLJpYQvwg8v2HsRHfzKwMdR+SvbGn0f6wcVSYFovc
I6m/p1NCKjF21PWbNKfyYjYOwj4O4JNAYnRKw/F7UAZnMpuqLs66PBBUPwph7ikJ
p0lzX+SM7lvb5ETXulzdG1iyPYxzn1FXqrRzfbYNY7ySrYnWUN1QQW5rzLIrwyWM
1GF5lAhf/Dhgh+WxCnPwEj5+COXNVZcGE5ZdOaNwhgLgSijtVvBQw+FfkCYR0enH
90D9M0mfosp+8Zie3RmY+iHestftrVfxjZJvNHmwLOVxcrM1t9ymqgYyhtxb35cI
`protect END_PROTECTED
