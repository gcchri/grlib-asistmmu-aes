`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i038Jt9tSblIt3KsZsnB7Q86KSriWXmzmaHwjfeDb/rlv+Kt1cIt59/Wx7Fez2FI
ubMFhZxzPu4OGFVMqmZ1NdOTdA/vL3+V0/cjXj+y9Pyt7FqZ4X2i717opTWe9xkL
LMWQU83vIYPlZi3v0bfiu9VABFTIoRSIRfYaoYx0EZWp9k2FIchCvycRlEVU/Z13
p5Gvf8QYUjl2AV0Y3/KR4EPPLVjsltsBSC8mzRVF24/rIlZZPzjhS8Hnz27wJne3
kJqkhcvm0nQNWBNvPyuCcai/fkRsQJZrFKNseupF1kgUL+Tt4YhSmruPmlJccAXP
k4aZBrv0HrWmhc1awjVMZcmYBDqPsBuILRAzjNTc06Lvt+g94shY+1xuOE1krnNL
LPBTt54D13qqjX+eqWwbEpCLnBX10PC+qjSr3cTL1c7wQFDDnpKNR5N3V3GXWuoi
vaQ7vwhU3ud0InehARU+afuc/DiS6huY3whEuSpUKjKyseBh0TQVYafHWGU+A55A
Jwikb1Z/LUCiV50sETZteaE0NoLoHTOclfsD0hjZ7i6hHbMy9yNLdzr/zk2mX9c1
AR6p2PaUkSRCqQPeARfq1X5eujKs/Sg1QUj9LzTTyS9kmc66JCUeT9REuWwKscsa
bulXHgVpjrA6uPD3VbTKmsMpV0yQVxVajd0aFS2m/P7BYf5ZNy2asesd9U7Kshxz
`protect END_PROTECTED
