`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FFnPNBwHupaCf8Gm75FA+tvaIu4HJWYoXGprFWLb/N63dCL3c7Sqq8FFnv0jtIre
91P5NF7Noj0qgzkpX906/7NPbhXIlHQu8uwebyS3lJvXfenZQnY6Zv8Rt9HAa2Vn
AtPZRwvIwa99Nt6j3RXX9DsCbCUOBs61Rmq9Jkt0rlMfJJByeA8maeovumo/JulX
ddh27FHFL2VUV4M0xqlIKLxGypztJ47zDVeRo/VVvQY1iWp7x9Jmf/NILWriyLPN
IWRY5l2xVhxvz4t6OmKW4BwR6SeMD4v1zYuwj2ihTGa+mN0N/4WqRmhSQCkiXmnQ
AzzH9MAKHy5MByqLveiER8iwZqDQyCSQpvBwr8+lp2hVGGBA0I+LBq3zQmu1iuJU
pXDATwqRIJcebbxfSX/trtF32ZRN4FK+RSK1ubVlLf0iu/zpLhdRyIWIAD5IF/bM
Xgs6PVfpC/ClDMDc07A6D8mBVUYRRsheagIv5YZh5tDd7zm5qwpyNJP+E6HGBXg4
aSuOa+AkCCDPEQuoHOVWEYIr4Bn10v5uXV7rnE6W6WPiKj9iJts9PQAW9k65D861
diFF1A9FhhG7bm259JpbNCVO6Xmw+VfTqFFYy/PvQoUMUi4DxzmdgQfGjjed4teA
`protect END_PROTECTED
