`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eO7bTrykrRAyi087MnA1Lg9q/y4qu7tfqhwL9g6sxIYcvuLzo1/3RYbDf9F0S3jE
iO7vSifbT2klxJ0v3GVul3bU4NClV410w94Rmt8pAwbBO7S0g/g0y0LgO8W1yu/z
nEhDqyu9LhHCOE3cALk/3JkOa6KAqpPYJyBJmFs13jcXm1l86QXhFuJ25jfFJk4K
gnDem9xHImgwkzqMKmr8Scy4CxBn+Ad3NiJIvM3A/ph09xqedAhGMXnrs132Ikfb
FzS/lMc5zbDPZxHlu8heVyjZKCloZFgDvitP2W2xRmThz35Rkmj7ptrBm+eB+iPe
gnj7RVuST9pWBXQfIDFmFG5ARFaxVwFZQ88zRLidXPNz0P+rtyoIgzr87SWISNHl
Y92fHOv2QXGT1cczInIkTH3dKXWTnSnAZMTJTV3BorGHpSeFZ6sTLYspecGEJOtW
7L3l+6B11RM6pS2bNPmMJlyveBFdicS/WWFs9MfZUXmqJWk6RZfk6luz2GrkqgVP
yh+X4IKn/4r/PfDOt0VESQXlkcu50Lzoqe/GScjkB9VZ8NN4wXGrJMGHFWGgqyZt
aQGG3bptlCzWQJgT3huoectBpD3+GEZ6pM5pTZPAj2dcAt6H1oihUUCQEpE/b564
0+GUdWuHIbO1VtqVzoo6zRd/j3VdKHJh4t972ZxLZuI=
`protect END_PROTECTED
