`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WOOxdrLa/ux9r7o/0LCjH5PNvw0ccFPanLbrNVqRB/yRkbqfodI8EdUbVmUAykBZ
CKjzbp1KIVw58g8fn7n/ujIyb/sp/BW66GKAutEniaJV3MUDg34UTrzbXw5vGYhq
uxYj2lTQhDtHAXVrr8/ha7/K8MTQAXSUTCTYW9KebGxXDwcb+nvGW5NyIydzyJE4
4kIhciu33uw6iQ0/eLSvhVUVK9iIrbXLWC77MMByhaYScHxKF49/8GiBEr/S5FD0
024A+Vk1xeDjIH1BnjUzifoQbiZ+sqDVWJPvBDxfGn7JZvRkLwHAxopP74CXtsp+
G08X5z7+qS6SdTK2WHjHpk8BAmHw8X++kBfvbl5eVngfCmgLeu17UXFTD6NWhC9T
dLLhwiqhsKmxeXK+Q8tLQ3jNGuoAEho68O4IxEZBhlybbKMPQtNLUFHuRIVgQu9Z
42jEZGegiZ+2hxAABZXsoI6+3ftN0mR83dyY6Ad6RFNLrzvM/K8cE8e8bXrptoNH
2Su4edIovxQIA/JommfkFUCLFvJaAlJi+g4ELng1llhsn/RNFnjIKg1kk962Jtyh
/HDAFEvaECcWyTtX/K8Ue+r4yBxqoSanTGsM00BLO7ll0ucMZlUYqPVpZix4NLu5
dAJ4cDKl28f7fAogIvNPOf2HEUU2lGpNIT/lJLQTpJtifSIvGg1xzzYx0f5TkNsx
+5TLwvSko1+rsaztosoHpobLOHsHs4cUT4vZz2QKsncVjFnKCKHsbfIyk0BjFQGK
9rKlGYCLE5lqChZz9z8H84Y5rPfNNIJFsWCOgFxjBfrS8Gl0GN5Sesv9nqzOIsI4
GIiJdkkn2dbmqHG+t4EZBny0Dpe2C46uv7O6PhWzgxKQEekHXQaPh3e2/nUWpcKO
x7aaUKZbe+K6Z1Is0boovzcrsocpWPNntC7UxKPqF0eJYBTgN6z71zCN5MvdbMay
IgCKrDnXYLyUcKqsI1Z08xKP6ofAdzwjcAB0ZazH+USGCNeJahNGRL6ZCMfodb2m
LkVKBn7uubQNy1FVuHxsm4aw/9MMXXVqLk1P8T/rpyf2/8M5kQtNaZrFdc0x0WvC
FZODkVbw3NwFdSQhL0AQ86Ni8VTdhcWbU9AOetGk7q/sUleT5+Kf8Mt7m3FT1och
J+eJwcbo83qMHiLdDdPy1bjLytIJiTEh4LlJUrwwfw9LYTwfJ0d56YqQG421uIAk
cS0qc0ydB+Kkx5yDqKC/T+OtHGWOJAIgJWezBKnqZnxD8L7+a6FOnQcs6dxESpZB
WTR5q+gvnJFzGAVahPE4BGnXbqjh+reOg/ADOWDJ8QyaqaKfaGhKnH7A5DEbOKN2
gOg4QmU9YT5R0B/5sW13+zXPIrzKZR8mjeCziKJaEgSuaB5PfhS8yVy+FnlvlihS
ZBh2wyvgcUUDv7tZBcLcm71cM38x45Xap7xxnzoPUkh/v2m28QKN147wBXLbXCAA
1LbZ+fjgDE6k2AobSzFFzOh4GO3FnE9RcUy2r9FAeecQ7+VPU2IWRiqCGLJaPU8H
KyTsYHLteCvVewTPa5qQR95IDURfIY8l6LODKtlTtYEILuivXMHU47J95/KM0Cgl
vWHIOBXoJNbYbqovP8ofZo2NztYtxikF47h21kWtnYPrg8j+WboSPVAXC62wlSWP
bwpzODZZbVWIHSM3qlL8zRW7C/JuITThoJPRan074InS8neJwfzaU8nh8SvV+Oiq
h4jFClKDmvZ3gnutM/lHaZqicSUWeZfprkXjTPnD18jMbQwdl/65avqQFrYzqcOw
rec7HyQeCOjRfnpjnhpBfxGvsAoz/IWMhH3G2eGleXzc7aB2ebPCeT8WMcQf0VMF
y2Q9iLEBI/1J0gA4jGgjghbLuO5FrGPXXBSg83L6RdAmuGY4l8/GkVwgcw/0jznm
gX/Z6oMKFExfTDOTMrI0Mmy1Z18UgcGw9T7LGQkKFJRXeta1gtI42i68+hE1tZ6Q
1eflWM/yQPmf/jij+tmyLsLDIT8oZOmdrmfxhW98ETysiKna/BKFbqFqLasCVtQk
SxYAAPqWwI2OTcnEFTPM5i7Hs4eheF2EiXzlTNJeLgObFBXKnVFhCuyPVBR59WGW
KwNnQq5EmImUQAsrFyfrkORfONmZMz/k5KbEhtwLhPIed9oQar0BzVa9PKhiQyFk
j6ut8vEnlMSAKQzdqeJvFuPVJBWVFLuN0Zj3d4hKTvowDnKcvsIIlvegXUd4LYmw
HUbfjXJYvihFksH8odSUUoSuYzc9lhO4JdIyuQJzEjdP+2BrhPpMKvb9ewY4t4ez
hnNKJd4SgdBZWBjBK9oafV2Gxv0l2HF3aTwvH5IQdyrrYYmSYG5ckwCWE/2g9e0x
jb2MXmkpXAJAZ4AViAkF6MH8MGjELWLoqJ3rhX22N/oNQjGuXx4yO2Nopyd7eXGn
BIwHDdtS59SjsQIzGRVVXAiYPziG+oNY2hE0oKvJg4g1yxqDaJcqgjzGZyCRrU5k
+biPPvg8ug+7DJhW/MpvghSy2XsE2IQxXaVf54LQRO+TsVgup3BZvaNLMnYAThlG
Cm37S0fjBBoAVhhB7TFLOYlOpvsnPWawxOlRJmxtcr5vl7EzZTvYfRgicKlG+RBf
xFR+PCZRy6za2s6bYY8PF9Kp+cVJbZjGSCT0VU+lZuLLtwfnRjinoANdvf/K42B5
z1yKbCECWN4CPs3b/qG92udBvgxnG5vyQtj6sn94YhOLJribYD7PVIha5zXnAiQg
vpHXVs345pb8iJo3FTRf6/DhMMMmlU4iDQ28vp07eHTUBoIjihBpvo2A/m2sq2UE
yka9BGnIyzpvldmvp2a4XWwjlLlo2bEnv46LN9qPyyV+Uq64g/oQPm9DAeUG1IAB
AmqR5fZaEGSPFS8U5B31oMypW+2uYAa3UEbyCXUvHNF8vWVsCR8DWUcdxZ1C4i1y
3nQIgfgpunq7ewetx4gBtf5mbhRRsJJJL/vL0usyrwA=
`protect END_PROTECTED
