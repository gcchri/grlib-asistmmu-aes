`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WiS5cupjnDYNzqOfcnHPQW459t35ib3AdxIVISGXqdi0P0AnvMFoVqV8fftLB2q9
HoZe/SzIM5xJGsDkGmvex6qtxgVroDKDz4T2d6x54z8iL6Kee4Y4NnNQy8MOKf3j
3UoJj49RVMvOr+OrCR2gVedcsNVIiYhx0/uYZ57oET5j/ZJ8ueImSIj8z5pfB+7C
LGNswaDt6evLU4KUY3t769vEkIAmcWMYZgcdxc4iYuwve4CHl4artj7PdOHiUb5I
+MGZJdcXg+eTXMnlYA6yu4m8HGd6ETY4YcR+VcY1RPNGveelXvbBoO5pwjJuYi6P
/8PmJEfWccouW3GFMx7VbLBtZXFTqM/WpBbLnpbqbbP7UzWQmb1IU1QxuTIKTXr3
bjlsdaGCpl2ymFkTTCOcDGT1tTq7UGoFkoFeiVBqrj7uSELsb0vjTlEOGe/+1f/L
+axcSvS+gxWhz9rOuY62kobLcIwn44cohwpxEGovzK9fr1ehA+z6NnXnzv5bwOYQ
RZ+rNrdheupB/G8nmEOdF7GnFoelgCyhidQJPg8zBvi6FNFrHsb4pBQP7fX2hpCS
OSraYPVU5a//OIdP65G+YxSEvo4DYpMO2JUYkeeivALU2QX3yi1egF59McxDbi7z
NUNTESkfWwiPl2aSIzLFfzIicK6v9NsMXGLR2GIdWgNDjSoeIJp4a2IwcShCqpj9
w+TDlMckFidMByCerwiHrrjT/p2826B1fthor21t/Yw9W2zt0SgatpfNks8b/vdg
MDGx+PIWzzIBR4qElQOPi6SqCoCjBiD9wqpflXkiJIhxmHXD2k58OsPrHjczd7g2
VrM5CcM4oXXm9HqQ4fqMXQKoB1Y9aSsa7RPWcW6InWs6qYkQkqka9eg1JHukYyaT
5t+zoAGj5jY8PnsaLck92rNya9UJMbHrpbr+g27GSNBEdwn1MVlnTjqRIqTYHI70
DdR84nL6lhWFjpZQvs/CORPBDrsNVcXjL06WAzNYfy4GVPidZ7D3mWi/Keu/QmKf
cnSo74JPV2li41YhztKdCxMYjIbvwtHgsukqcjtjsEYucCX0rVsbRg/52VkMjUoD
SwXRonwHvv8dYj0BMc+YbVjey0V0ScXHw7Xnwf8PXcSt8ln6C60aTf6tiMf/dYCh
25VFkWW+Kwkk5f778LprvSGC7dMMsQ1XB6j4QqLPU0G3usmuWk5T1UwT9J7P3auX
7e9SOdpYiT8JoaZPVtcZ6rb23aDX61K5rvxgydRa1j/FgNOfJ40ocbJvaPBoqRhL
hJMPCPx1vXnr0sAm1ykcON/u7vi6nPUeMezS+PNZfL2KjnK9aEXIBK63fw9g1v/5
fWOo8DkxWEB+/bOxhcJTJPbeP9zKQkJqtUufgCIB95dfWnUa+k5zRvBCiFKpk9f/
6yyKDz/m/Hz5Jm+mUuQhmeZlTLA073fKKHMtC8z1eHNbZMKIF4bX37FBVjLsUmTo
zxmmwjHpdNrb6xZrTZql86QuuL7TD5lZfkUXM8EclTwxtV20v3SBG04wOEufMDeN
OHtKWRQZHuh7G8c6FKqviLpffXlYCqx+SeetWQm7l1odyAUb/kduNcvkaLQ9hzmQ
rZDl/z61ihguRIvEkN+8uTNH0/VWhTM1xJ8x/C+gmSHUEpEx6FpHae8TaQ8qkjHw
tiByrjSqyOaKZOdLkGLm0gO0kD+KUOdZsxLDi5M521+QJLDPRAFPVjpjbzIe3S9i
PPJamKiCkX+dKSfrz86elVVhV3bq46G76tvKLTLh6CJRATeJI6Vfv39fo7wUq1Cl
aiuyGFutCyMVyN/ywBMNPvqKJrOcB005TQd7b577y/ow/fTaBbCGndmQ6lYgjqhI
cS0OimV6OQvj2VsnbNNsX74ynrAyC/U+YpQrSuP/s4qIaxVzh/GniPEwjJHsJbl0
FiO5dbjLItTl+V8yFEZY+nbYswjISdLuuSsSsOEXgCNmytm2AMWEci81vE8pKFB6
Z5EOVreEZVAggI2Km81zxJd9FBHy1tnZPJ0GndDHJn8UgJe8eIFwCU3XEnbK54xV
IBqPmRbkEpEjNhndfQhOjsy5op2qMP1JnosAsbxjHxKOB3kMjZsDk4d42ixZfyX8
VuVtHqAuq+unsWaKmk2fQCLF1FP31QgXXVmEX/jN0O0uPDOTxZ+r3MmhIJtQMwTO
PShLq8sXP4rLPHlCSUVoAvf2GtrINTEpeMX0f7evHipI4XPSeopsr3/48pRKvCNe
lv9wygbzf2FARyuYYpAZGzv+kXoRGTpOBTi35qVniu75hxgJH6+2F9KEuaZQQVSd
kDoKNTwhYo73o2ar/4GfUDN9ryE8Eut+hoQECC5bXZWx31561l98aYo838YFG0TN
YACzC6aFw47rPt3dk7+N41HHIQqK9vnbd66yYmOW0Y7wzhyeEQr0+q9glsCR11dR
ck9YyDjlKjwlFEuPufMREnFGF2rq1yty2KxV6kxb2N7TtpxdQXyIm9/TiIaUOf+M
f/q+LRdcoVqB+c1HWGjQQbavKaXERUwC2BMqDuKniELZfiUoLDG52lCHbJM/x1NZ
NGdLIdNLB6evzpRWSjcKivZaxc9CE78aKyHdlSp29PA24zX1LxWgq89TigRCOKRQ
hc3bdUTB6lyl/AeUjhyMvniNlI1cq1nypUTIIb6hJ2F0Ytk7AU8wgJ5hw3Pi7Oop
Q8Vhtq91wBNhsYQo1D6ur+C+FCuTl6zqR9wasNkwRCk90wxfn4T34glV4eacF63J
OgVvcJiwfn7SGLagXqSIXQrcShEF+S/yBf3Yghjx4R/IbRtZzfRVAGYKGfSBA8Ob
u2GWD3hDHpUNoS2RN326Azqji/lNJATyjWS/nfmWzCGDITggv/gL8M6dgLSpw/RJ
Np1TC6E2rRyq9tajqvxI5vRqqI5EdgkY0YmqByjmeIfvJSaYkxD2YPh5K2wLYRa4
iUYtt50ZyEdAXYmLvCmwcdHSh9EFQ+MCVjaNpvU0EwcQxpQxIC6q42JTWOmS4iE8
iDsHz/sUYPRYDQpE6an9owoiSlm6+Kh4HhaLChN26c4fv5+Ds2DM/L8m2Kvf2SFK
xpPPs06j90mkxhJsEKCnmVxrJSLRHX2KiCQsFdbcvQb6YlRoTO3HH7TrR0ZkzBoQ
+B/jtO9DRu7/x8Ji5G5JHn5IRjOhLSl/SsEMXVDaakxjBUrZttFCFhTNwKoVBR/8
YgkRN6J9AxLuBRvU1go4ivuGm+xgEu3yPM5bq4ccJJafmoVQQdX3P/12NOH+9aqH
19qWqotnDdFjwEuyzs8GoG3uImBSRLTG0siH8weqdyLL50xdVo5K/1VAffkO00tP
Gg985p4qi6ctq7fKXqdLUsWu4SAqcC9GhF1PbEJALFNlraHJ0nl4QCpDpcoksaS7
G8QY8Wnm7ncUeM4fW5FZ4plcsI/ljEaNpfBqUEh8GmuG2vmgnZCsOsGhR2usQMYP
ph06OfiwJfIPj81WNowvv3Jf7QYs14Zb8qJOXhkjo/DYN3NJesJ1N4axPDsj1Gia
tY8oGz9RXiUO+quStw3IrR7EnVOlcF2VDYum613haN3ze5PPDVTBQwNh6cJQT5zo
642wME0P4GU7urIYeBPDCYA9RLH1lJd8yrSPpIh5VCUH9ZP9tyX4awVzhV7+q2cw
`protect END_PROTECTED
