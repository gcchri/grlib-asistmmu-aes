`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bx8iJNjqNmKaFNjnijMzJNkokZ3/evD8KXLz8qUGzzkzXaQ4WUEgRyt1OnxE6lHz
IcZsxcUR9AFFGSvxjZEfBh1w0ig90+MkwGzAMGEcGIIKT6HeHuyBZMu2uKbtBGKx
Qyl2M7yVlgxgIAj4Wp6Pj51rX1bF8ijN3WKP5pOKolTG2G3vkfv577+kVjo1HiFK
+tVwCgLUvoJCPgaRdwvXYjz4+GzXzqiCDPZxDh3VgW7eHPxnT30O7J98BKXVuaWc
z0NJFoGuPiU7YjwFhkr0j0crzj29BX05Ht8tFafCKQDXEYhllI/vUqB3Do7oFlmF
`protect END_PROTECTED
