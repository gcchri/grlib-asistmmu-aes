`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VePdVYxS+j5K2v5wEpj8rjMI2XlyV0GT8qOzl70IomEWrJN3bqKXpt7m2aaT035V
KtWS39WaxpfR5C5VjfO5I6U+/rqJELner7rRP9rXlAJMqTkR99VqMWWK+aKgC0eK
sukMBiXcK2vJ6+rwM2YP3bg/uQi8JmjZAj9MBsdP9yTV5BwzGxUzIa7nfJuNKz40
1+qT96IG6CjnfnScJ4jmd0351gGl8oRgGLdXWu8110GZnsgVUt+gC0biTNwA/TQr
uCaKczprmcEDHMNw2OsjbBrQX+yX+c7UMPDnkFQ3wMGSHy0Mejrk1qHmcVgWvJVj
B00PUScl65+oNfJ0f3Dh6z0gWTc17lPZotwGEZ0V3YQoYDE/XEW6M7fu0YRmGDtL
MOH4Ppy9I0qilaCvkHsCsI9taswTlLhgdDAQDFfe2rBc01Ep9jRTWY713UtUBbC+
XrIH8aBNxAVHvCDyNsr3TeNijgUaJVy4elu90ACw1hqZirkz9amc54RjufTk7oJR
b9qTt+CtXa69K6OufBhzNHAbCHBV3jllDIpeAuN0B1G8zDqytkfsOobyOMhcXDGq
zbZissMbsPYRFKqqvdDaAqqVULUj0o9NIgoLAWOyRu9LZE/RFVe1Du3JQQhLee7Z
m2QCNLQtG7s5SW+cCmoKoNT/t1TI44b7Dh4Mhvua41HUuz2H+N7orwreON5yU569
Eq2AEza/yp6bFilI02XJl4xE40yaKCRxQFYWLGniOR8cwxSakd6su4Opo6IJW/WZ
n0CPCxvD9KuOn4whORIMJVe1w1xGHYb5nzDiKmea8QgdYrBlemiXVMpRk9qCg25h
6omnichlBnJrEu+OY2RAT9QFYSoPZ41AKWaf1D10HQyZxva0nOllvaU4z6tYNDME
dOZ3G2VUdbDWBIqSFvlDV7ZFZ+ds6WQ9Y4/0qHKfO0NE9lM4NqEjcieYdrlsQDLy
DibBuF1+5TZOVJu1dLxTWXAqCr614LdD68VBqojU4vbv4uSqjP3cqA1IlCqs2gVm
+J9ttGc3LeHjh5be3wbQKr76+wMUMZJSnGEno14nCxwPqy1M49xIGlmjbYyXl+P2
nCJO6R5o3HbC98z9Yir0uRwhX4mY+UEdJsJoUgWKTC0jq3i4Sdn0ISmRm4jx/mHK
ohkeHZt/NYeY+eGmHo77epHd96nI9/aJG6gLFq9itKFE9NCXf0Sxz99UiqHSghoy
jxWTguPEVbIK8zus1bPSRTurww0tyzUljLWPfx01CZlQ3p3zfZw5NT1ODKS4bVHK
ypykB9z6WPY/bE4+tKr7gEPun4iJiR6CbEykWdeHmREdRTReN9fbSk2Y9eJDUNHV
HcYlniOPkHrpA/4FSognj0rIcMdh946TqEwu+xfSgsSZA2rxYWnkggiDW6CAGlzs
wK5tI+ZYThjeKlNJwKtO4gdCCQj8VoTV5ai+mpcACBCtYxeF3n6nhRO1yhWWEXON
K+9MSRzzKl1ZF3+VRP8SAaYNFkt1Ce3ce6KO2YVH3k3wUHJO78Yej49Q7Gy7/f5E
AEdJgKRPrOjvdq12qmPKVjp/3+IzDYbl5lE05L6b27qPpIpfCpXQa+DPWww7WTtV
NZOwOf7/ueXwdOX0BP3nZ2h2j898Fb/Ze2HxynsykI/OYQ0gMDvMFZ2gJ+F6Ou1O
FZDJz/hLK8b5altGVWUKODOOUCIglwB5fwNJL3MKP/aHDwbwdRP3bGa/Tih9NTKD
g+HIZtqWp0iYpMEtbTPBnGh1McSkqoE1NP3uWpjEIX76qLS7BsQakuLODaIZDRRT
2uPZXheKpoCo8/4tjxog+25qC632Cq5o5MKhLSyHXVGqYGXImWaa6TZixzQeATuy
EuP5Dj+1fNbERW8JE34QkzePbK0QDA9zHV9n6HeIke87b859hcdt6IzdM2rbCI9r
PwAx8OEgfEqnN9qh86rLiO7sxAWcf0JG3i0fqC3OkCjOu+/KLbKqx+o0SxGJ5oeI
GjL1t7GiaZuwaFke7T6jaWPvM4SwuK6LdS+DFZ9Hu6/TCUJwXbvepqMouJxfplqS
xq6yRaMqbUv+j6TGtt94FYyUuUjSWtTUwkyLcO1JxwoZZFsd7SPy8LXtGMmcQxhm
pH8jvNlXfbaViVTx5PRM1wXtIwQUejSveU8j2//k044VzgxynzPqdYr+yz/jyNQo
Z+25wvmDuRYK9JvEWnrMjpus13QQPYR9TGm61KRI6PhzbGGoExGyPfUsPM38btOq
ppQ5r5a9+934ikXoR2hHFN00cop3+AMf15UUsSdyObBy+fWwhgrJULJ54JPfUus9
HLGpLhfwP/zSQJGs0rQFlnLev7pXkJLjnhAI+pf0WMR7zU9Au2vWWhXJXRuWw6hl
iqyKSaW/pZq8oJOYILgr9f/OAFe5T5ZZoQuvlsOddFojEvwkqXjoFDcmSIYHvbPg
PgO3VLMnLsh0/Sc0d5xwo8DyctR9nhQ8FR2tEeiKUBEUty06WBh6OeiUu8tCVvdR
uqnoTLNvDW9t9Muu7ymZWA==
`protect END_PROTECTED
