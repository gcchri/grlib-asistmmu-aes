`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJuy4eZuCokTgB/gEjBbqm/x3buxxCaD14jvE7bPA1Nf5m/HHywBGbj8v3I/ztjw
SfhuvKWqioUso6MBtjbX7LhHte0fvCEBw+7o8sXIyFWkCrie5mivQD/N20GC/dXL
8mSlyP4Za/PVMfyQlgdu4X+IGJ6YWCDCY6fwokInRsmYYtyHT53XoyT05K5JSdav
Azt98qkMAVbmonp/sLwfhP+gjEMEjY4tWPNU9We0tdFtrTTiRwR89QGrsl3C+pqK
Smh96IAbDYjj2VkPK3oQVua6B/9nQg8t1SrRZDhmfiI1ye44lWKApBPmitQCPX4B
vz98eG6yutQV4z9k1MOtOpMXg39qXEiWg7i57EFATc1bjUTMm61QeW/cS5A/uTxC
QIMTtcdNIzsDHDZRv4n3RVWF8hcJqIYg51pTCeeZdQ95NEk/q9R/nc+Mf97ad4Lf
k3kgAma6d0IAPTAqNvAD7EGo0f45nnRS5bgCENKWprBmwQYw+C3KWWeBJdFI6G7q
n41pM8Cx+WudWYebeyABut5xlcOOFHR0S31yyyNC3AmH/gMSAf2RMNtPcSyQJb0y
3mLdLjH1IultHxSNXTJ38DMC1YFKGZjt85HozwFAI3aHDfDfc7cP33U4XaVZRnEu
fyvmBmLTu/Ei0SwwgApmWKE5zgI13lvcpZ3B4Ei5Lp9bwt4YRergK1KmBkIul3GR
NGLHRp/HSRyvMx5OuQa+xWwdzAPX3jybgPAzJHK1DrV44UKLINjPyXEF81gPJRrb
BdeMywbahrXV1Ba6J8C/MopmqRIJzx4TVHgUhehp5WY4VkK75U4PYMcKQkFZmlDR
+biRbjA1pzjWznKl6lGJ0xlwnp04XBLCMfrotMPqE/U=
`protect END_PROTECTED
