`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
msrzjVpEFpmv1MqWvx3ZrjXNxWVu/fc4tkEySNZVjhcHbtdCwp4ODLANo5CMHKp6
4fHWDB03o759tX26RMCI+pVIpLwXo9fNgUkVIi442/hFiqGHNlrPS02HEYOaG55i
DWIomMbRWkR7wVrzfBS2khEGFNa+PNSNj16hzf7VIczjSMA2FLxb8QUxGzU6CHXf
DEGy0vpFq+1Yvjw/bRk1/5Sd7t26Yt4xzmUL2hu4ociYQr2iKHKUdOXuafu0BDa1
fva4RhTGYneXK5tuP9ZXusGqPWb+ArHB1/TlIUoriiY=
`protect END_PROTECTED
