`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0kKrJ1/8f3XzOO+C+zwqzI+Szm6gXs/sKLVrOVa53dxBWxSv81Dtydd3TmoHSRmm
ofKy3zWUvwlTahBwvlgl9mq89IXJMZwZFqXfd9Qsgcy0wFWmrMSyIdoSKvkkQroD
SzQYPBP1ObQI8XfAXOg9Rza4dkMDgUC7yvKHNW71uyA6BtfN9WE40oqyj4MkS3dk
K3dVlVti6spthuLt+iAHfsRO1f38ke1e4Uo/fY+wgTSMJQwLyxoTJin6Z3YjIx7l
MSNpdFNY8fpxYmHEnzHfEF8r8zFM4X7V5URGmEVmDzaEBF+eTw3szDPj90IJcpFC
kabmBfsYkdTFWhFAz1CMwpygWYMxe/QF+nmh5iuT1fz3srml6X1SHQHLXZ9urKbf
WutsmsV1EFK6ntnBnyuKxJlJKEknAakTNQnSXmV4V6e6tkes1Su/N8XL+mugaPph
TTw3B/ontnQV58QH1EeqAPe2SKehhANt437md4NjEyLh4ytOBSFL5CcOiNYcfbhP
yTcDi/efmuKCJcxDY3yMAi2JAhPnXfIwXi92RPc9W2jXExBMJvUud6EMBXpwSixy
oDKpiOFDPGRkhv5qQQTwyGyFKddmLCB23EM3ftyhPr317KOdpjVnOwZnwltR3eAo
W4sj96qftqW7/Vol7QHQB1gsKXKS481smmrR6J+Kry1VkmdszONriNdAarT/NFIK
+0F1c/0vFbVVpeXkA/WE6WDCyoMqra8MJPxS9UYkwF7SluyHc6DjGJCwCjjhNns4
Kc/lSwTXkPWnq7Ds1xbKNbUf7+d23Or7ZbL4TduBTJYrgdeKiTbDUwA2wWY03t35
TriKaEfxsemcXO3tFaoXr23kbt5TQ31QRPXBfkJR9W6Lhts9/its2YeYg6UpC/V6
X+h4UiMWAHE3bXWrRL01aA1bqcZciq7dEb95g0aY02/ONWrUkV8sVeTSnoi8rpwk
E9z7Hcaaqcdk619rGIS4ltxWtrTCXQwHR7tKqmLqgIwMhs4ZTBoUVVyoJ9H6JrAy
MDoVp8XhST8OhYDJJvePv+TQnW7ZCVZ0Ejyj2sOnIIwjJfkTYS/a45MithxVSOx2
UYzxWsgGq2Ed/ye70YKBct66sPzGM63X88TUd1WqWaYgqIRnm+lT3oT0wAmYYIag
WyqWiRj5rwCKiziH8kF3B+OYyfC5HpSV2uTNg5vAlw6VuC0kT1/BbBapHhteBzmv
TIm02lF0YiiL2LRK6kbvA9HwjUX3KEWEnz4qB0joME/beZesdFZKm1igKfd3GpO9
DVIvZ9UsiTsyWeJxcRO/Y7QDbkh5+7AoKhhHNxs9R4ZaLQ9SrNgWM/xkmkjhtteC
8qyxM9DxRoNzS64wLoe9tANKNSm925aUAoMvx9NEunrCOBxcDjb6crKqsJ9o1XS+
IuBSjOheyVg57VlxxZkdvqSC/2DXDdx+SB1weNaIehvvfgPRXGiFpjYvcjtno9Tg
1DDfYM8JgwoFAFWQlsS5gg==
`protect END_PROTECTED
