`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
izSLtR5U+qsrQq5zmRJp1WTrstV540vP+T70yIGXMs+wVWGSDwcHq3e7dattU3Ld
IwbNsnZSNppU6+9+PvwKhKdl4btFNC3t8IWj5wHluCZefpJJD7leXIYnSuiy6Ryc
Vc28s/9/1xZj4CSKt/e0SpvDopO5F1wZFp6ul0BmMxLalNABND6axkSrcOSg5qQy
oYdiRlaax4CKtaX+vt0H/L2Oq7PKnPDYwDyA0LUntFbSLuFhdVg0K0xjevC7pzfk
VxcIll5AMKyD8BrfvvH+gaSXfadUJnO+gVcM/R+Tmtmsw3itWGQu7PNKWoeIJuel
+xr3zHo8mCABdtuGOvmMZ7Id9hcgrjjUVaywRqmFYQ6egM5F6/LMcG7JI/UO+crg
hrgAoEJMH+lanuVJt0agbN5++GB1e7a49y4rhwh0doqZ+LttDVIwmKkiRWfyRhg+
0XWv4hWYpEcEy9EL39z3bzVTZY3jR3vtzVniR0h9HB1oaiF+vxe6zKeGrYAbaVvX
tgkpUgd2EVtsXzbJjHmlcDU+4U3pcHqbJqibulf0HLh2skuGVYy4CFJYIBX60Sju
bzBKW7thzUwMqRxvYeA0NnW8q4Lz/bFR9kdygvb4vOJ7Dq8r7GCPMKbfpzt38hoK
0dlsiI2YgqwknWWE99hMPOz9TpLrzN1vagpxtEPj98/JBVMWQ5P809rbSJcuG6J8
37hU7E2xty30WQmhlCGAF2JR9VhX9MPQNP4fBJzc9Bs29jDbPfkWYs9DDhvFwj7G
KNuyY7E33fy8hDdk121Axwrxjw6dmjOEH/cKBe/2DebAd8pIoR291QxFPlbEsoSn
skBU1XHbZL8+e2/cKJCFKRBWGPm6hiLtChcCgJULHaghoMD3tbGqNPxVzaZgxe2K
`protect END_PROTECTED
