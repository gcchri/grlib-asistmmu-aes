`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Niet0GEtf7QJ3kPGoMfTKvG5yeQM5FHVITzT7ZE0UrtgXlMofSzPAJXgtuThqqRW
TmZUFS6R3ZvyV03ngbfMKC09BPPLSDVM0X+KUyzLVTsCKStmBO0AiU7Javc8pGhB
mTJOLAyA0e+XhNvFjgp5laU/APwosTnc6Q4vZQutXLtPMCUxylsi760FxgI+tN5L
/VrYuxiVzQY5PQXaIu1s67qyoz6GKg/bce7jE1KzOVPGnA7nHZNzuiWhOEkxOjTG
YCDnVsNlVWgDQXqvX4ACpvQybgN1NCW8voOTmx+QtQKntQ3v5M8RnnqjGTczCXWh
HQoRL1sCTsKIN+IBk99p2rqNmS4rSRjfV/4cJEungcR30KhreLiSaIsWR2/58+PK
buDKlMqxPBK2yH+LSl8pF8IhlMDIOS21IdLPb4an7mos3rnJPRz9cdqvP3so1Mnu
OgpEqZd4wiDRkC51yb6pxFqfWmTsAdIMycjykifXoK6COZ4gwKHoODlSCeKf35tv
NgK4RwVYG/gAyVaSCEUjp74YPiUVBrW+FRdDG9dGcro9r6Rgu1k1McLCepRba/Vo
P4Wb+GNXn0+aOGnCMlgRZIiVyLQ3QWdQRcjHtcxYGJCQollNmWF0ShLY140YsF8f
U/vXBevQrW/9BmP1phcu/CRDXaMkTXW5qlQEzBTsY/VEpzgixuK7lpmImAr0bkiI
+EyezSPSl1G3X+8R9h+YC4BOWKnv08rPJ5eEwN8Au6pnW78ZFKLD1BAddKJdCEIS
QiHNcrgsaSYmK5qnDW1z5h7DlFm/lvhPmU5mtH++i7mC5EHsm7TeuXCyt4l/2R4y
tnAGTEyMKI8llZKerm7WIAQK3G5KDo7Vz5gk2Aug+kpa8htzx7EQnv2Cpzqz1u2Q
/3lkBpcmPO+Ee7zvVIbSFe/4VUtwduVaeXuAMoFPE1Ov770CTWxgg8niU/6FangA
zStZlf3HpIFYX8JukyINWeojPEuAZGirsWd0JzsZ7JF0VotOSIijYCEVecrrUq9J
vIUZxnIbO1sPAy0GptS37x8Vz+0WhhE5C9pIvA/iG0Lz7o5cfir1RLyxH5Vy/hU8
mjkTuS/NpW/VK62upEujXcGeGFRx4C4qDkqw1f2ZQ4r3sVOuVjAknXzcdvGDhFLQ
+b02hdAnHaTKgUyAlPF/2laijZrMC2alNamY0i/SxugYARwNYFiqZHZ3kS0bCG3t
dRwTCeBcIHBpvC/whHeOf0oDSpPdiBcE1esxryizoRAp9uxL7Kkggm2dowaWII/S
qEhL5j4JjSluXhGt6BAb7gct1k9T1P8F1wuJJcTmgnRKgTarhACMMYXMPXZbH6Gz
T+V5Khm7XH0/MSPmc59SX5VCETb6MFwuP8Wzo5h6UpyIxhbqoEplUD9OE/61DdjA
20FZt6iSoece5GaePKoAP5zGW9/3n1luKK+StbCpmTAUr63tZ0P8mVb8Q5mzE1G5
HH2eLshIgy9EkWgHbswg3eCzWDu55nU/Jw/RVlK5wsNlmMfZofluGfKmh0obtL2k
dQFzf/d6jAWjZBQ6JLVKwpMcOXokG4lMH+tWPdTIyN+vcwoxWOoeNJI58bEhm8qg
jneFWoCSRkN8behmXOwe3ZzujJNPpoN82hmoEUqP4wTaOCtmrgo7PTAlpatmKEwk
0b6FvqzMAPKOw+2ZHB5BdBxxOPyRy3kq9SgJuNMVYuvSQzSFyV602cO5wvcQU/eJ
iafMhG532BO6jgqM6pOW18vUHGzgTLyqw96/QUP1yyGLXavi2ccrxz+pbXkLGfwy
3A+18crtm5Udtc/d6VYGHkk87rjf2dI3OBCeK3USsCu0joHE20vzYO2RTx4Ej+wd
3z4pdUmeioPGU8oPkPkvMygtmaFidEFXCz3QR3/Yab1ninVZRtF3gscjKXBbvDhv
WB028tvAY4iT+bw+1mIsa1axMqCdYIBRT7H8RMzFB1qAfWIM6WpWlhnRKKyNtcY1
sU/QQ+GJ7dcbjbhceE+ajHXfK0Z6LicV2BhuY+j01E5HIanx4fx/76vGvSCSkcwx
MVY9Qk1ok7F1WQb4SY+/zYDzY7s/D+CDd71SoXHqB2lnPJsN4588dCLTUsWzhah+
RdlPog62HIzKqaoOeQU/cgPMadyCtlPfu8tci4AYoWIWgXnO2ANh1IReTlOE8Qzr
qh9qtEL5KNoTB/rN2On7IWfGwTcw+PHOlqMOFC+W4WFREyDOAxv+0lCHsgyLO6al
9TSJQIjJJfluSnixLjNyCVGVgV4NGaYhhcSwd6f/wuN1PQbSTYPh7FPZ4b7TqEoZ
6p+pviMm9Xm1bNfyujXVXimiw0eKx1I2urcvqqRLYKYHWvkwmxXts9K+/4KgL1VO
P5goxo3sQ4+VpmIapWxMUxiUFEqPGZoCvpkDz5ixYlDj71LXuOW5LYrnBcew5Ofl
pHrMsrNvRHhy4e+UcUugsao+0SAFUIJzmKhcZ8ymX+fZ3P6qtCi/yiiHm1blg5hJ
2U4lFFtp8ucHSJy6Ad5K4sgD+RFwtdc9bBrNMgBMyqj8IHkqkPrLndMNtGuDD406
XQYfx+pva6Sqg9Wq+UcUAzPjdMjE5uDbHTgraxZ5x7ymfybSOElN+yQ9sdbXrPay
L0VK6PpAhb1/oigZHnr+ocM+kk5zMfDyvEZfc7aNarTE+xrg5YmPRGFvI2ceEns1
9iNSJCFA5q+O4SGUlocyyOhjqe+E5gG3kJa0T8NCHyBnabiIhtJLtW2WEz4skHJV
Ikx/6bvZdsYaUGQnVRh+rGOT2aNWKK6V2ReW665NHuetW5r5t5AgCcRlhA4rHl/G
IzHW8gwnBTn7IYJ5ZfnsJAKTPrxWjiIwXCj8T/vgYGalCZcRdYVFUAjA67VMMps+
zKG/quCMLsuFXcy4xFArp3J9bg5sd0bQRUBo76xvrwqOipcF1j16ZwMEGC1IMepO
vG011ajPX+yLnXxW+cCIivt/+ZcqaYZcqqs2L+qQjKCe9xs6hvXH3BFk1vKpVJ1I
LeEBfPTCpGMInel/deInWVqd8RsPhR0W8y/tcWQZCqqChNfnWzfyQCiMzFoljavU
sdUrt79K9eZjyfQFQH4A+sQy+F5FlwAH5cau4my0ld9je4SvI/zlFB17XdM70jKc
ZH1Y85gbBLEr1UPcikS9cmmHqZ8bVc8qZ0wWXpWSZFEb7msJpnEYJ0ym8wePrh73
nWOF+1Q2VE2BlGaSYeCpJx4HQ8SSOn/6ZTKAhuQ6p9aCQOCQ0ALMmt3mEZvcLZnF
b0kISMgKq1sKaFGieVm93qyQndad/D0uthTdvWZ+cdHT9238GXDZjDq92aB4tHYY
nlJLjNtc0BfqZFh5R8dGo3WG21h/0fhvBWLaf4RperYRVa6vTwEdn6tzOuevrhG3
ViXONKgnzwB/tAIBqz139AFV63pesF64w60PbMywUsgngjjpVoXLp9eufayYCeIJ
dioOueQG5fyEZqRwmcVZPb0ipsyiZ670SYhyH3qqf4u0cZXW7zBJI2lPU3rxMaYU
if89gayglG2TL0HzJ7OEzXoBPz6anxX8g4wIVjk7+aQZrQA0CEX7jabkUHfncpnC
mRF/Xuu1lOvXNW7l/eZNIjRHRtTOil7XAXb9/D7DyZT8jfeLCEa47na9+Ogbv9F7
oWe3/us2iHBy9k0a4Fbe3U2tGPHOGenmC70UezN3ePNmpfeu+0jbRVSGzGUBQIfZ
FrbaCLgrITJUiroHklN7xQhy53ni+Sh3a8JaoSw2QojK5cjzVLlgHXsLW+E+H7WD
KS7Iq2csAWgqHD+TGyfyv5YtdH6b6GsQ6w53GIYoJsE312zkWpfFn+sh97I7QBSw
A+h45p/bbXBnnLDTtiyaWKAMYCX3yNRsfm7xevIbAoA5JyjllGoIEF1ZmTYcfE64
ZVomrnEeUDKapIotnrj05zgtGqjaeRpMv5KKiSaKVI2+7INdCFxLHtrePOknAe2Y
XuvMgd9HFilr+ONgpY/w6KjSIws56Lx7zJpq+6oSFIfcxdTtcaUtTu9oaNKWQ//D
sO/iT1sOup2ZDSHfowM/H5oyMz5stri/wPcljfOrAxLH00Ssa0nl6hBHiJVZn4W/
93cqIKUrXtttKcQY571YcsZZ6Q5s7agnrsMH+GfvC05/bVJ1/UC7WbubZpri5G3e
2rCGPNawdVnoWtssLzUdeeHocadaccUoB9/m2VApJIMVUesZMG8o/RHhB3F5F50q
HYo4G19/mNWTVWQxSiWFiPR5JL9RO2sN6wIRzsDlxo8QL4opjG4FfiPcPbbBNkH/
P7b3u7Mlj+CpoKujrwAf1MVfYpRNkP/q6NfY5opUnFXOZlY7NJvBnHQ1/ON/ehdf
8wb+Yx0cKPDBLVL25Uo07o76UOSlnz+FM7yHlqt8U7IHmKcfp9he9c7ZQhPF4iv7
1K+V7JvL8aeGCsH5iMB81R0a8SB21BJdHXwbmzxCyR20AdfGE5khyl/YbsKnCF89
tB+XMoESlYIId4C1S+zc4wLJwfk9e9iKhoq9r/jkYobpWkHtxdEZADUuvoH/Y4lD
pPoiWfTbQqtXkELgeHY9Bc+fNh0K9XS0WyLzqpIW5GlKQYuybCDV2n32pdWLkz+X
tm1WYW5PMR7PkYeqUKzYJNDHmVqRZGq0WVWIWcNk8EFMA/7PgIBoOI76xGcSu5Gw
Cug2q7gB9oCwRgUfwniQm8+hI2f14cgLz/SlBkrih85SbdcCqFAV2Wr/tzfAQZcf
dW+ktaLqzQlo8cpADdioUTmRudua9esF00yVIBUQmiUO2OXwf5w7hsz9Xa0CXYD6
VbsD8qC/CEN6j+n1VR9sWBiHgdDqLF0rjsOIVC4h4LGdvzMxr8LDOvYDdzbipK+E
p8m2/kzfX1IZnuNnHJBxpgb5GmNjn958G6yK3xFO0XNpHKrSHXlCFLRlj1fihUke
v7zO1nM6Gsv4DMVAJHaFMH10T3NIfAsHYl9TGeml7cJyAI4ThGEdv8ljh0rqnqR0
4M3cQmqPeXIHimbjPI1eSkVDCZGddAEU+aEaWXjkugHbwmjmNrQL8BmmIfNxHu8g
mZ5a0dCIVol1T69BR75Psst/5zHaYuoiiDKBf1YHH7umJ45EsHdjYMZF6tUz+8Hl
dcdKoepOutb8gDUmIZVw2PaavVim8DC4yScEYYEMQ8Nh9fZMxsQE7y2qPg0/CmZs
DZ0D2GCZKpk+LIDv59Us6juSd6kukqwNgVXY39kuGnYBbPtQ8QtYAoiQHeNNSsaM
raa9WfZOsN6Fgk3RKaIMeCDuN5KciTg4Hf1W8jqcgOfWO0KGoGch4GFrq5YNv1/I
gc9LDAycTvm7YuAlRXabTzMPfL7qcp7NDZ7STbJ6UOvSK+OqtosPrqxBtsEBnLcH
PYFo1pJ8U1fZQ4yndXQtzHo6TxDcDWOOxW7w/sUaVoDLV7E2gIs9bzHGw98btTDb
1V4XyICa3waYRchmgcY9Xgn3c3v+6WxMig0hP3QiCYd5ySvboeDPB54rjAursJLS
I6u0TEfPodk1nwbfo+mEX6rVR8wcAL0HIM6/RUeIGTIOtwTOq6nofbZSw/Z0pcuQ
UaeskvkArcKwXtdgxzYMdgiBtRiCh3/mf2wOCMwy0Qh0ajIWPRua4uRYRREWq8/a
40HpiDXfZ6oybmuRYZkmLTYOsAcpawBltcLstUJnVLAwdBwgu9fFczeNyamww8pu
4tuE+LRi4v4YIubDyNMalT2u7/tnAS/raSAQcaZz33TQnF460baU0E0s916KHPx7
DjihcZbBkzuFGRbTgk27wbFbdE3kKzHQj+MsiGBrjf116zMbU2AZvaZbAhEiegaL
FsuZToGCoSuibslvHjW1QrQECyv5Y9rrL7KXpqL50grMatCmX1u2fmQBFZMV8XNR
xwyiYnXhiBlADvVxJ5VTUBT7Fj8lM+BxRV8oc1mn569l21sPJ9Y7Wns6zHilCfCM
h0z12cmaKuLXI010glxtUgG13AQHs0Wz+ejgT/PS/PE7tIY+HZW2VmvKfkIEHMzJ
T8bIAg5BmVWM9OWQXHBDaXjkBJ5hzuhXKML73rp5L144n+1O8XREFlWFdsSRpQXD
w1yFA6opvdN/hVEQKcax1F/n6hnZo2NMTIhklnpLPFMLscUutI/dQg+QTT5Q1+Nw
LdaLw3mQ86PocHh7I5Ftjurf7r2BHcreb4F7EChpcv82mHTHvWW+ouDJI2viVFb/
8FnItW0f7x26p9YYXmBXYqZ4V/FNk9npToNPYora0ND/ciKftv6P9ThamXrcZdKG
IAFl7EuxulkADhZS70dRVxbCzd2HuAIPph6C5QWZMJDTh5tREhrz9fjKvOJZgCgJ
6SjGQoCc9rqbV7Rp3fglkq5X23uIx2hHT8G3TmRCSkkUFm1CXKpwH+Q2K3c8jyNp
6wyoPe7NdaiqHTm933T9psoPe2etOKLZ71Nf5ZWtdpeWmybqSCB4ZtCFR4B52oH5
pjCloyLuWvVLY+4QQ9H0qUco9rOMAH/TtmAbNbP51TLl3bEphGZ30EUp+lY32o8P
p4rfFrAsKpujto9AYCDdol+XgRFaViyPjOrjt+yTO15WV87lqvfRCAWdpZwTmwqS
0kKICai0z1ss9BMTEhAR08Y2UcbOq7j//+IomdDOsqoXdNTagbtjmegMsZBts0Ip
77rxj70v/dWSp0xo3OocyF8Ys5xZlAgkDUWqSmNZRsrBTc8O/sDauMScGyuIhs/8
+s49MVGqzkX3EJ4G2VqBSbhp5rpR5uWtv4vYP1r5V78f4LXCYM6saV8kbuc7BivJ
Dc4HhtFnD8avl4Jq32TnM8/1WlC0D1fhB2mOkELUnUBq38marevcVf184gARIsh7
M9d1aZ3uHTDUYruHLxPgkyxJiMqmnW39Pe3LoXGhl5jq1zOK+uQXl8g6V5DQgra9
xaWCPg+10wroPzjRNOTH3ja2qZN2zYmkL5G7SZyAQ+7ktf9ayMsUQq1kduIsMuP5
Pww37dtcnL7bvgZSUrNksIePgoM8KI2u9+ZVrKaMW9AaYPrsJHzjlfYz2tJQHaZT
Fj5197Z2rO2K/zQATTXhIM220zM0+QFpgsPHJx2Mpcdng9FCUZG8wfEc8pa2T1dp
QQ6TWw0qW1oGiQc458LjwY26g39X02W4FH9bPT5XC3hOMVr/B+8JyW4JFIT1c2a8
sNClK8nmKJgFFTvFjNYk8zSyAPADzMycbD1SjEVsrjvubLJMy9Aps1bdlxkGX3Xt
3MByWtmgFkSJh4UHfpKQ7zDJV+Fx62v+co7VgGC2cYPgnBtWyTOPlFkfPIhEHAO0
gd5CNeBWxBnmi1xSaolhrM5ziOWSem+GbGZTURxtBCxtnAz033x51sS484+RFPKf
+mI7uF89tZhb51Wn/JerULrJNZ6/KXp6PDBxUMlJ3s96pO9D25pjV9JwNHOLQBws
gYYeZRLh/XuGQBVmf6aTIIsQAFeBss6MAW7+9jJooF3Ma8Mj6YHaUvUfj5n8xtc/
jORIWeuZXRJZyLlrD7LXofYYlqCZMM41o5gQMT+GVpvSH+6vzxlqKNW5KfV6hVXS
FdtzRaytv5zYmnP2v2CBaHGyvHb+TYa51K1MCJLhOrKARxU1Nqc9ywnb/4SRb62f
MV6h+XiFR0epEXl9zyaFaeIqqp7gCozEZzdHBzgmiJxONjmepJtIANf+0WGrHJfb
/QPnPUNvvEVSj7cD+T7R8zsSvluh62KqfnEVlTIYfQqQf3qBgxFWepm9sAr9jofR
Mwqly5rw4Jw+jZcOaZSSn9t/Lcwq3ZntjSHpvOEThpYKezkKz9xKKyU2r2BaxsSE
hcOmfduUwikYLoamAkSE2A==
`protect END_PROTECTED
