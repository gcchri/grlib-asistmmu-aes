`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iVlQWAVjmseXv7aowNKRtX/GpKAp+2xreZ92sKQlep6suePG8rMcJ3ApUkyXS9R3
wDxmShfxXIDBcUoOSWUhySvVisO/dhGA5J/GgnZz3d2/MXTQu/ZW2LqVkl/jfEDb
ADNlMxh6meAOVr8oZVKsYNrI1IXd5IpqjtjJnLoqTRZZlWRMqohi7cThga2Y1Zae
Y2Sko/SFm2ZfVhgdXKXyuI3ByTsvG0tYUYAjHnWaFu4tRd+ZHFjIkFLImfSGbsvq
Kw+cKxMHYNHYhtLwNap1jhO+RZjQQarK/EqLPSLJ5YlhlYB67NDn8mdzHPXpO4E4
y2ZJaFycYi/QknkdC76VzBoCgHjLmHXIsKioQoXABrJXJCcpfQg7z9hSo2iuggSs
Yrq50jBktOkj93dJp8erTH9Y6MIr6nTkU2ibWJlpJzSkzCzm/yE4W7T5XjhektEm
VorB2MbMYPao4+Buo6VPfha7+3V34pposlSdegYfrWc=
`protect END_PROTECTED
