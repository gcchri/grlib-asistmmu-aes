`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYq0S3JzGlUMzkhcM1RLvfwl3JngRaAFgsdD2PXK3t4NO4MXiL1aYTEddSLnO8/w
k4R6fvrppFq2sa8/edxtOjGHPCO3fgTqGRuGHCwBLE7LEofde5GabpZi+mQY0swq
hhYfxrKUwy2cANFdM2D3QsLTlK/g7KOAbGgn31/lZgdbqYUCAjz2IJ+XG4xoYvV3
lCwHK49E1oWaoURryJdPh1I2y2CZhW9WlRZPNE4glgrbTYC5/0BQ/JrynLPUZoT/
/wkv6B/d8gBRX5Ujuq7susMgs5TlMpXYun1krSYHnJZZ8sU0Y5R/vi51F/xAmf23
m0UYHgVWgwZapAfRP7a209GdDAF/eOBvSK59yle/FE9hA6Gwuh+QubLoGLvfV2lq
uFf0uCEdu67eNsSri/bNnOgOGO0Iyi1xxdcbaT/mxBNHvVl0TkueovvXHYzafOQg
bF1aDZkPwNlkbq+PB3hY/gIwwi6rN5Q8SbpQpKIYXN8fi/e9ZxNCVG+wJ5AVhlII
`protect END_PROTECTED
