`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yj34uQBYFkLww6NGAfXruSnKW3LhROlGN4LTDanJrovp69KVIyR+x5RO/7yIl96
oE6aW/AATrXUkRCk0CBvLUkbqvak02A5Q3XhKUUranQNU33IZ+JxWYfhmzBPFIQa
qnKkwR8TKvmad0u++gAh5CDCKDVHiOYbkk3OQu71+mulT892dkFf/DKvXEOlJX1U
jwO9p/Fymrn5KhOTHc6He9Qn9ZxzXtQ3N6A11q8Qm1Zae3VPet4QkwNz2FGPFr9E
Hfq2gnm2bQlT0Ir4emlSptKgiWD4RNjfW69U4Sxl3rXvOKLhrSTWCo6V3qzpZIrG
8MQA2adGkNFUefIRnpkkfDpTc/iX0tg4LiNoTID3hRWFBfJr0lJg8tnf7qK7ewH5
hS0qfncTl4hOGw3gL2+6qhocNslPP8B7ydL2Yhb1P1EJsKBoWBkA2mMupnbazaNX
YQcEDs48mg3UUAwgo3voUvBJGco/OXfagf7vQMrDEXRAfnm1JxVUneixSmJ+RJoU
4h3AXGsn9aI1wONaJECuLKCNZfPSqwDxz/h6jkAk4nUE/FwzNgRTXNuW6F79CR9H
t12ZuFmg4FPGQ3R+uUdQWvTODROnfzN67PYRuNk1SxRgzAi41knHp/pLfQE4PHHY
6jvL/PWXTkiMye9Qn4Af+bBZjIbDm01NMO400nBL/94=
`protect END_PROTECTED
