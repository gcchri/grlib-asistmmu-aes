`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDnkMcFTfl92wE95jX6y/9pwjE4hu0lvfPEUYBCcCZVgCz4mmIJ4b8vbURHKYmV6
Msx/oFfF4fJ+/ysFOmvWNtEYqhyCxJbYCYCaBAvFNbzUWdOSJBwNFZGLvKUVaHd4
Wl5IRuYnHRJrny8K4Z/TZzKzFMPkV9QmyHIX6wuGplzh2AavhWx9rne+WKtCLKFZ
zCaVA6vRFcVfsvpEzKt/+SydqU7iq8mGOkGcUgO/ctBk6xR73gMGWpouSHLunWcA
toMwkTfoGwcQSrJWbgUnxXpxdmu8xsPjxKWFcvFylsJgQoRwMS0IvFWlFg2pPmdk
yUVVvfeaRSDujncar5m/4JHev50P0k9LMfT2UnnNkFd2p0+5hBZMC4eULu7RV6Vd
4fj5Rk4nhSQPGwtgxqJZJYfYPTx1RiBTOjQH2vTJd+FrZbzmy/PGA9X23MIyjR5A
+r182UVz8R7f4Jj9lTlQ7pK2CqCJzRo9D5K2a+aOF5UtFI/pOFQHWdlLAbx7Ftr3
3kMLX2tlzysH87lo2JIb9csqTSLL78rqp4o08ItCy8oAZE4GmWUBzs7ApYZl3l7M
94/kXoGjfTB/hrgUxjmR9kXMBUAM5sAxS4jRq9wWvqNyLNB89GndIXW+QdXl3bAh
DNFn15GnUTsSyHQYjGtBgRx7cmHD8MrYBn6mvyT0k9e9pSAGH6lrOR/QQqkpNuk/
ei9Zqg/V2kSDVApclrLvv3Ff9Ta1lp8aGh27u54sIgWJJryqaujSKN6d1prJoqBE
HayDLF4FXyLepl9EagvUIzuXNVQT6L8KxGp/C5Ne1zRnAjU4CGCDNNte9dqikSbV
`protect END_PROTECTED
