`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PcBpR5jnHwehfdp6i7E7qBjUE/bQNhKaZl90IVncrCKKfQXHZhGwMlEeu27/QKQM
3Mm/zfxiEgsj3OtoKHoz2H4CUjD063V68tejjklr85F2I6khjlp1FXX5eg8cvD2Y
+p/e65uwiskMYuhBbd4Nqic+4WifE2Hw3tHopv1TKcXDRx5s14CTq9ckDUwcqJJI
4Oe5jFNU757C/vtUA/NcLqiYzG62C64cJYfynLh+VEGQ2oD+lNgpaUnBYf8RD87A
glt45Z6Xw+1k8B2yM+GokDpYoOP0+ujJQT5YiJQ8cccwn95QiVUSOU5rKs7xP07W
hPRe4KVu/YtV3Vg20eQ111F5dU1UjxkR9zRNWd9+4CthXp0Y1k7OsGfVVnuT41Cp
CmeBLruGl/WDU5N/NXcYGG+CykuTWrkaOZmsp4T6QsG+H8Lhq7ABIXgVE6eUjCPF
uppI/Y3/UBZjZu72vdstWR9VnG2HV9IYOyBYicSg4KYGMVl1GLuJT8CrqAJEGKfP
jcy3aitCD6VHOehdQy2iCarIwpK3dVag+vSvW5JGXNM4oWSqEav5sA6Jl/R0RJQJ
zZoenxUUNTcEGfREHdrq03vj2iFJA2LQ5C1igX4Gleg=
`protect END_PROTECTED
