`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tTdSNy0d9lBKdqMvxY/X/PQw9trOfzMfWjjhgQjPR1jehMVSw1ZYzIcI5n+9Qmo3
obbfb6mhrXFwylT5YuxRgYvh2k+iskctSvXURjILiUHPDOjxvZgnTgCCqoIiNPch
u76Z3rjZ9CpPgm+bVo8+05Ta/rm3/fS2FXASuAE/EcoBbCauH7PDwA5MBgeB/CGS
Q+ZOs9kDsWNT0B+ApRpl2osbZdg0/JCk97XAUmSD80LRGkagx/nAws1t88zGzGtr
l8EoHqT8g8U9MXOWqhONbtEldVCjkPneylf6+hTcOCEesyNlhLhqtuig8g1lDQnC
8r+vxxKWvGPP69xE0NJ4mEwDm+n49P+n7HGOetzqJvPgqJxcKBfCPPo3uAoFsvw9
0v5dFCE3d48dWgOZS432A/oyj/2IxQ4gA2QfH2Tpaus2hu49kHIt/GwgEiPE4o7S
Ky6gt8TsFJfrYLuJTHgdk7rO+HJ8kcm7RZvyjwvaYDUjXwkq4klyUxKAW5q+I0aW
SC5KDSO3XIt3cUEHbgT2R+A6v9Xymxb34EDaeblWbIxkRK968FBQ1ckhj+ZEfmKf
465k+wuwJFMNEe+IbQKybU0nNjcmQao1b9CgzAqqcDbMRz+eX/JkGb6+o9aXR/Mg
hQc1uCNNrFalnUFc5fERxBW/JID2e0DPzNJFFhTEpZt8o9NMgOZet1aDZNoXkzSx
ljzL/aZMsRR63pdM5AZUA1v19yhO6RLJ6umP6VkJsIm2IetXko2x5QaH5i0YCgug
SxEq5uXNl42hKfKi6sRwP2cwXdu16v99oPnddznMn6/hfofDCWrhfOA4VH7MKA+9
HoVukC4eUGHQYToxDRMxl/9+UzwrmelCwAZczqdUfCzd+ISX3YiyVbvF2n5Eadyl
WXWhvDexK9RDI/dXvcw3T7IUT7tyl+qSEDVnrXkcDQi+ggrmddB2zEPE+SSQ/cGn
I1RoBZyeItPi5/IdQCmf82M4uu9S3Z5AUaU85vFTY8lhOcwmFK1OnjaiaSAwfw8b
DLSjAIXlSOr/rIkGLw3FcQ7DmGYMDb22iM3/wyvuS+bOIJ/J2s4M6UWJTTZnqZJ9
wTSXWqYAZj8652puLo5WAHDF5ujnZuMrtzWeEHzS+h8U1V/TMiEGWfzZCJYBidjY
fpVK1qGY2o0jR3B438ly9PxdqDUUCAU2A37Go7FXuLBvLk4TwNitC2vlu5M3Ogu3
tlpV1BOCq51mj5Vt6KE3w+Tv146iWsesGwCx8Tv9ZPwFzyxTeIdP8bhE7kItNsBM
vHCMmXoKRYczkraNJ+RLnUwS2I+0GY3jbVmMtXC2zyLObU6qngPhQGQQe0y7mw9C
FlTAx3ceZ0PxEX4++CsQxDIiY0LhoSpsqo/d7Fl5AQZd0O+42LPNRj21mMqOpR96
N24tzWPguLEEQBg9KVYkxyn+9qzIK8l0akSC0RGY5v7nYob42/riE8xw0lAaltWw
XFFjrRpuopP6EeEpaXWVzBFh14XBgA3+nUzrdoBpK6pEXuRn2jmINFak7nhEV6OG
VwarRGosc3jRQCgpCIJKqatQKmpAh2QS30tRsW+oRFXk+zsZfnI4YUY75i3bOb+F
xq/kenc6fEu44KfDrSIduLO+jbrp426BdGAcxovbLyUFSq2V1mn9cpLWctpFBNxD
+i0Bfud8eeAgLfdKMb6lTYg4hlI38QI1N6HwjXuLuh8aDUBIaAilZZ9+qiRThmFX
kPqnZcqXphFMw78jF3D+awb7BobxLk0j5EvtuVBPbFabZced+bxAhqPI/uItgYsf
+egWuU6QV35lXcl+BLkI/1J5iLll4rGnF/1vPTVR1UCkPbjbgCOIZHcPbdfsLkzv
wbsk5SHpoQYcOPW7+it1j5ZIjQRNcZKPohylf+YIYT8jZTjcpC3Zot1MPcJBc8ER
eXALF0Ns6FLUA94pgrzqnrh7kkf5jFk5VmoEJtT5xQFFCW2zCTLzX7ittS+63Zss
3mnqWcfW+Cpazs2DjhuWwoDKZuGnvM4wUuBI4wJKvwdnx4D7rhj8en6OROVp9dYz
BNw0X4QFSzpgrY6mDQ9fN+zO154uIu73GMQuh3gbxrlP+E+MTmrm3A/jvlRxpLWg
mW/rjGTDgR3Cx4S8r3c68/uLxhRI6GtrPfA573Xj84lhNJrZMJIb7o9zzP0o5QH2
miOP/HUQjUTT60Rq3Bb7cymunN9hZty44MgdZhX3GE9HqgYq8O3Q95La/pjIQjgj
RY9UD9Al5JgPg9WRhqiVpU8e+tPar+PU4DUUf8En1ci3Yy3PXSRCjOPunTBWzh5I
EqkcHfvysg0a3/LN8kACJDhLJv3YZujTxa2LomrXJd7xfqaobTS04tE/Jl7ce3la
tRQAAEe30cZaaNQExsUxZo0//cteh+EyoE4qtmt5LRtNzCtJdFoOGNiYsQr6Kw/q
ReyzKSSO2kBRdi4FE4/KaFlePI+NYC+6wABN1hQW+zHUVG8bTVrafMw7Ng6yylLl
8OIhpt1x+1m3YhO61zoAT32NUQnIk7b5+L4me4vKjrY0jEZG6oqnZ+aIaYqPKYWe
Be0xfHsvD3K5JwIMnoMVwo/yHdu0Ns2C6LVk/65089GcC0ZETqInlvgWEBkX2SXc
Ns9u1dMlRHZHH6cpk0MyX11n0ISXs4gIkJ/axTK7R4YqbCJtn9DUBj7L6hTFnc5x
BgYWuQzBnfjfa/mI6FhbWlL2ymWjq5PeO1F9j9dMBJLrmQMt4WgddZ3+aT+HyfCc
sKGYtB3qaA9yZpX8fjj9xR6xYbE9XWIlUqbmrddvwAx2tpD+Gjl/42acjGy8Snf6
NCiwzbafOimYR0kGg5y6SoVcSMvy4uvY0F72+CYwE0lcQNIZ9iz+JtqkqscypmDg
ygdzEKD45xG24B7EKNgEpzy5De6QmLAhTbDBYWl39i7s5LHLEmArMEXUHPfkJlil
bYauA0f7t8IbWJZqpWAooSFXvezEpQRBq9Zpn9nWZPD2iRnM4USyxKDrHqjVHx14
wpwOyVOzr7xFGafeBc9XCl2gpjrF3tMMFV3MHZvKiJm1P+zp+kBF8cpQLSdmfbuo
PW6gxksFSNP1jEU4TdXzaZUKjpkqvLlWYgiVcistaUNf/CB4ujpA3+qMbabQtbGb
nVDltRx6DEzAyC5azwGGGt/df77ozv2OOlYgRg34WfgZVYVat/RAOj+mxTyEG/Yf
+3vUYjWPQxZtysxMyYVoHWZKrU7n15Nnn/c0c02jk+IWKsu/nZiKNGHAsPUDXX/4
508tl63t0THl+aAjZjWfd1CEojpZTNZiWeKSXaR5qkKEAM6JU4Y2bK0CPm3okzpA
cgHczy2Q2uvVzllVJkpOZg66sZblRrO1buZyKDqyL8r5UvV5Nvr6k4nfssym6i2b
TjNK+EI29JggAdaJ9yWZeesZLhdc7E0D0hgoxSvkvxlO/Ut2OIX4BcIDRtn4nHaF
egpr6WH4j/R8wtYD4o12wRf8O8/BcVcVNCkIRVCf4dcsUx0Rv8obygAwfA4LUh5/
A3xUzWjhPSNGqZdMrnbZuxhD7Svf32cR6kKDuoaxq8fSUhb/RBmowcUWMyesKUK4
KPB7NuGidTCOKfTXxmPY3GNNHfd+EEyyImYDzOKQxD0z5jAY/e1R2X1g3IgV0EYe
Ub6YSFfTQANcgmEJ8YX1CrwmBVdgb0eWp+AKVYOxi3T09DPeTw8inqa2qGihUqZE
Oqw0LVz9Q97H8p7AXSwhrB9w381sEMu+XIYDV9PZhOBHp85vmQze6DZd2GMauNEJ
UamTkq5wW15JgSlGCjmbhht9xzuhPSbOepQ6DXBLbQzvSGhte20D5oZcq7tvMXqq
SfJO3uMwKO5TO9cTJUhPwJpTfTmDZ7Wbe0hXENObRB8mniDYw3uGXMaQT4yXZBd/
HV55QHtDrlLnO4lUVFaKSlVnOwl0Pg1WzIIsIDIw0+dcEQDgjm7JDo/uwVIV13Sy
ryJ16bU8oKJz1+LFq+YXsBk2JojhKXJE4rBK1VN5grd7XMmTZGqOJmkojNnRncPi
kTDw9xzsSJj8eH2AV5E3jTT6V5QzZ4aVqDudm7MJvaiVCoyfwdZwD5mteYWywzir
6yj5bKRcBYE/M7IdJA0SSW6lZtXVjVw2c/YMLuMPEjir2ceGYdaKhMKqxYIcQ2mZ
sKqRBlPaANZT9N6ckS+FH1fZFtUKP8HlKXhaJbizZSrr78YJeeuBKoMh4oyUEeJ8
/Db1KPW0j70LVndF56kOv0B6Dwn5zY37PoSDsc6liMMME/sq79ySTbRjHtRjUrm7
+YswjXkafihU8mrDd6qCLpGb+zx6VhAJE/mik/+vAl/3507LURkCHlEwRY8nNLaT
EapTQPHUbKRwxORV30lhlivdH6/W8uIj8CpT7iZwfeOgeRYBNWCnwMGZjT1l9mjZ
UM3BQ+JAKF/uyqmQ3dllRLTGhdFGz49kxnODwqy8r94jI8Bsl7yXp/DEz9KzoNv1
QcPHQdaQs3t8aCf1InTTkjqEp8SWnvVs+rnDh+NpN05ZDBPWRgKfEIIlLo1Uvv0j
Kp7zV19941P+RLXoNA+dKNl2Gzp+Y4d05lF5y2gQa3SL1su735T4UZKAeda1zPQJ
R0tVAZd2tYj8Z8ayXuvqyu8tEXekQ5pKglT5uwPSUQEc1kL1Vo8RDPsbH0MLdGNB
gLqYfUgbMZ/Ef+ZV/x/rpsWPFJ4JidO4pvHrQhMCfkhEvM4FSSVdjcCcIiWPtAgr
GPDeSaWJ5fz6YUTwnPUHlEeZEb9JLWw4USdE4qSHCNHyshFov0cp4kKfOPpBvjvO
atKge5WYKM5v5zKof+E3uSIVWoHD9XHSoYGAyAqmHeLQNFN75+DdBSLcxEXqyHBX
8d9oMoDsrmcLmyrmbxejTsm89d6vXokahPcWfaDcxcOEEUeLmTp79nOdzTWT4GPV
XDAVHm7Saq/a3m/YN/9n4BtnalHHpyddD19jvbPgVM5+vcDa0EoqmOLv/SAesdgH
pkyps2LofxNDD6IaHMxCWznQBkSVMvq2uhXj/h4UzWLNtPjTZzHFbVJaAMujPzrU
g/Lhu0WCk6k2N8hsQlvzgIeKCw9O4hpU94OScT/KB9OBVLFC70EXNIirgQrVRAqi
ggV9KTy6lgPRlm0pl55Et2q/DLxxb6+3xf2OOnpkGO4YCRE1U91tGtBD3C9tfOz8
pThhxItQloz4F9BrnKJdxVtQg2hVnBqm81DHuJp2dCgXC+Y9v+RQBAHaGCoGz/SI
1+CTfHvxPXXqfd3PGL2sGUZziWrnjnuws5D0ODSyx84OUK/8sRE9iP/YdxGSZpBO
pA6zOdwtFBnMd+LcINKJVmB/0R/dO/OhdAt2Tu0f0KsDyn4f1bYFeQR0OnOGIFwW
bdVnlUOQDpMRAp3QOy5oosy+DLOG8XeRT2gUQVAcobyJphym5u4yhoqKIxDgJ6MR
0aZC1G/A+a5NbUsa7+2Q0XHIGMHhR69cbIAgoYsYkCRw3gpq4ir9694UqrjW2jVg
YJdfmYAP3FMA1Q/224y7QaoOFCoxwkpvr2oBwFKTm66QSA1jN5/2qGxJanAchneg
2HF16VXZobJXAYX94Bd5z45if6DyoG9oJwdaUiitB/uJQCaTRYfpmEJu/O0sbi35
ixhKKfbHzKIYhwcp4qqt349DdC4TuzDJqzu+NzptUe0LwAyrFSfp4A/PG4q58GuR
`protect END_PROTECTED
