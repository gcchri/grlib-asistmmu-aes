`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oe3/wU1SzpkB8HNUnIY6iOOcBGGyE8QTp+g8o6yZ+16DklwNuuWIDCYw68y/HaAg
AsKW0szWUXB5tj68anGOgQkQwABNf0K/yAzeXGRd5VW5N+7yi38ysVpAu2xNN0ar
QwWLExu+Fy0jz7UF5TvXZug4j5KolZqRT4kooxiZKbmpdeh9GtdcykIff3bBps5G
tDdOlVKlroXpPAfgRn00nrKpfAdFJSru7Kfe3Dy6K7XRTo5rJGizgDDz5OWkOIF7
2iptbUx8klbQYRGqZUSgnK3Cl+EbLGZS9WMT9c4WBkzPHNyAmLQaC9oHGwDXC2Vx
QXpoij+Th0kDj3SbrenH8SHeq49pmQiSTQfpZbIHg09ec+O4Z72O7SApxdRZqKDF
EpupyK+n6GOuK4rnTsd+5Q==
`protect END_PROTECTED
