`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J+YUxig6k1eXOM/zPF49mAzWvo8BaDpQWTPJpoZ29LyziTM3vzZ40sxxUStr5eMj
qwHPPyu0z1FaKKGbQBihuzrBUpZtfWOetQbptW7+DzCMt3AG8iwQ2kBssdgKlM5s
b0n5bR5XttzZNkOisui55p4e5r14OhhVerLoHyYp4izQVlXQQl7rhMxtB0Yyc6Dd
hhFBEKNWrOhQmlo0rQNGFrtLXwZ0fxvOLgHRP+ROiLqJxAJ64PUKZnUW2niZAY0t
zDTFQVOOiDhzOB93CMoeYwBGnX6o3ZWQcgIA1offmcPuFLKw7LX15dnXM+L4swmU
D8xEMhnxPvbcGuxIDfeFbsp33tCFuFOSxD78aNLJ6F7it6Ggv6gK3RHaLz9UUBcT
`protect END_PROTECTED
