`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kS0IV+EfBVlShGU/XAT/Cwo5g6tyed+GU1PiPqpxRAEveLc6xiY5jKx2Nod8VjjP
1qs7ClazTmXwQ1mfyHnpxY8GGJ6HmqPLMCJwHDJS7us1yDzzwaLw6bXZ2Xm4BCB6
L2W8AdnbLhBGV6o9P0nAa/YAttLf6ZQKWiGWiANy7dLNs2/R2zD4qVLmYQkWgMDj
NaxqAlrjvtbyZqflN8ZfBCnDb/H+kwkWPtTFwjcBixrP9NkUBzASiRx6wQMvVUtT
8Hzr4w+iY41Lx/LZzxDgPg2Y2xvOPQzSevPW5Tv9BYVYFyR/7jraVPxlJEIshjfk
eOO9D/oTN9RPnFeB6yyJgNn5XadZX/UrsNRuot1oSFRmI5k5t1zf39rauD+WIYoQ
xe7osXrR3Cxsp2YlTQeCLdlm+uk8+zT5Rp2SGhWA1Z8=
`protect END_PROTECTED
