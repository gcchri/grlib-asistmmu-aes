`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Ss2M+0lf+TBCefqbGR69uOz53OGJdm5vR7blAjfhY6n29ZYd+1dIFIxNU5WUGaR
FRBNaZNq+4FtFSZvq8leWanlqyA7yqkt/RaUa2SL/LF2jQWphSwObom2HKy34AkY
Prxog8bPx5i7bbmZ+BZqwXNYkyGwYawnhAO//xFaJcOzEMDxcaCEXKz7UhCp4yLL
rn0swBQYd0tqUfjZOErjaIhp3l/m7CUjayx4YNGUUfkPD7YFUMjObYEXh06bV9F8
CBfRiVBGCZzbcfiViD+BYJv0EGejVqjPIrUcjFiqID3uLl/d7SdZ/+VvuJPWZ64I
lctG8Kbg3Vy4FjgtB1nEeIy6z3a+g6YxJTJNIXHa/M0K8AjdjAR3/jeoMMgoP30C
krBNXQOXo1I9Fxwl5kgvs5T1RrMjRk5/05pdCZq7mowy5QLgJKl0Tai6Nt/qsGED
AnbGCSBO+8H+910osYbBvk28w2xIhyHSljbfG1MxZEXruJGI5SWDgmud6DGT1Id0
qclgRiDTXkLxjQoMNO34Zw8Npr42HquoZuofU/c5ISzwPEeJk6H2hSYM9OlqhgHW
fNq8KvV6Rcmua1rxZFcmizY8FtjeChUENxCe+OSMO2xe/tvq/xcRc4whyJMNjfEV
zBlR4ZjGBiXvlnSizkmMAyHVUB0XRS1/ttqcnSSE4PcY5tF2uIh7KTL4FK8RcAHD
kfgHYxfuV5W94R0gx/m8+OB/CZBqo3WzegbcDBVXjMxdKgxSsqnpNKJnC701HRLF
Y7dRNctbTdaJx7VPKs56kRueuc8W5kkwSMYh7eGT+euAGuo4MHWHo50p43CJqEe5
DuffYJwQlXIf+u9q+C7ACg6Jd2meY3WFdTBnmyoPRCwCm4rDBZQwRQ0HF0cIsw7m
EHwe4bbO4a+76wvXZAsKu+38lZaLb0ieQTKx1sMLPEPENtZQdOSCdZoz/7sOHqVS
dv8VSm4LMtrYY2LZeU6TMKFMQ7EGYVTY5h4pjgWNgUJQJsSUCkYwJA1ISpGcvE+y
0QOBtQ7ksakdm9cT6DucQSLw4RirQG0KeMV634pFHT0moRJn3xS/QqGOaQUG7WDH
JhbFXDHTVM8HR0AGCytyZFnkY/gpXO3nwmMgh/v9ANQec7DpKsaCZubQhSO1RITl
`protect END_PROTECTED
