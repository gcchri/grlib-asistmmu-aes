`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzZeu0ESDGrx71OWkPwDW8KKemiTW/udcCfoQd/C4efzUcMLb1TtN/jeYpInq5vO
i66BxiQDHHaSnCT6LYFP4iom7KJvfRreWnvNCE53vsq44T6XunUyl9jp77myqvIu
QG9h5/gf8k93hs+S/bCrdS/R8qusDwwayIVJuD8DeGe9thMd3BAuZD8ZBQx3OWs4
GxhJ4VUBSssdwkYm0uzT7k44FwppmMYW25ITuWiupeoNr/93waayq/iUcRqo9ICK
rELa5UQiOShQHQ8v5SKLFy+VcBKUqgJfmFld9eKr3gmy3K4wJWv0bWSYwQOJQcjn
HQ8AWexXkWwz2VeckBQfbxylwnRStQLANfQOLLx8N1K97p493zyItVTm2wJtxxqD
lw64B+bbQ8iN/8CNWp72MG7J3XShMxh4bAYi/2p64nGBa62NGxaZh9DahDGUxvz9
ceHvH/sn1jx5PVBVB0R1X6nCbGdmmhY2SNNR0JpSMuOYa8N+MkL9LMhrzTt0uOb0
ugWCUaLR+lcoBHgLCO/iRnj2YlbnjXQ5n1gcqZOVTPHMvLocbTulUQYR//62gnTz
YvALFJa6ed5m7HzuaqClielSpI5XY6hKUHtnPHS3PPOl9LZy0l3BjDcKgoVfZmz/
0+CcsXYgDy7uhw6aT4EmXVGmG+OIfYL3r8MQ6X9Z6KW8qIUVW8C9On38BINzBo+x
8MaxPSb0Fbyw1MrfcdEaZRa1rzAx+StPA0fnZL2GlIEM+/q+Cl95zLfdj7BbyEKQ
gV/ynGK5j6meXmHXBhor4G/RGvMiCoe0GmBU4BsZ88XBWA/WPddfvl2eKvRS2kjR
EEXZnMTkyrT8oMtFkuIIroQpzXkfKYDsJ1htOqNLVhQjq2/yjKh+bhoIXUgasmvI
`protect END_PROTECTED
