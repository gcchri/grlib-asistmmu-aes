`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKdg8UJ27T4cNGRHnSyf95/VLcLehwWQVI1S24GDutiriGmenggMLSyuq0soNyhj
M9nEHPm+Ts8c7kaaz8VgTKNX5zn2LkzqyL4dNIMZA361Ka4l4F/Yj1wpiFAO1a1u
NDOMxF0197kbq0CGZ0QYZlrUF90XHGnsCmGdN2XKPiOFfi2oPXaTRavgnHPa1yKc
DCjtswh2a0TADD24DfW111YWEUCDl84mRXbt+MLGGFjDeU8yekS5hjeUi+GMACoS
Xt0QzOCV+igoN3i3pzjz3Zw30uriAwdqvDzI9xl3Np0zxiL6RV68ckJDdFP8PwFm
`protect END_PROTECTED
