`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jg6SWaAAqmV+w60ZBfolsBQTJNDVPBTy3J0S3l1X2DjRd3/bZ6qLrximZjjiwGbE
thge6I3T+Z2aad90DAQWqQKgZomRlZ4HWn6uLdVjnDZVxwx/emPB02c9kaTD5vfJ
76JSWcUCcWhHKDhQw/EN/PhW38k5CZfsWHNsHLIydm+nv06TnAPMAtjDiOqjCw7L
xyjfuufcRTMj2j4K5svv9Phs1HwVt+dbuOyvn5KCknmVNhAWbdWnLxZJWi6+y0h8
2Hi2GZKLkgXooa4I1mBG0RcN7o7RCdnXAHdIroR6YAlEwCXtd3n/Z6QMSn0evT4E
SYZhPzZki8MEj6PLSTrTd1sapa5GVDY29yvQIHnkodOERqbdMeiRoFOkg/WJKfW9
6y8bSpMN7Z1thij83YYu+0K4xaDyY2d8+DpnySe4f9GRNtXgDW+L1brVQP+XZwfK
WnpvyHRZbEFeyHKoCnIfSCAiV5iXhwRbGidBWjH134MOXZEl1pBjGFIvKEywbilz
O/eQ9A0tFgZFQgLMKR7ATWCqsL3fifqsqbCjoFPg6XdckTB68FeHRiGrBoqfevxu
I0EjZSUKQa4L0wbZoAUrZleRdjfJOBm26GEFhsKKd4sw7ULhFGWIRw/VZ8g6lU27
u6mqzaGn4TSsWJcZxLWDO4lEzdyTJBB7k9k3UChDWRzAzxPHNMlAo49HSha3CLuk
91xkWWf8UIqV5Cv8/8F+/fWuUlDdNdyffzT+FWMQ1j44kNsZN0QF67DiJBuRFvG2
9nf0viWckpSXhCrIejqkQ1by5nULxxZ8n39gK9lr90etS9XOLwgTGOeoPBfy1O1P
fDyv9LELRR1ju5nR1DXUkhWmgpb9yznuCDn+EHrXfYOYHn0PR5V7YUL8xYYdcHmB
fUs4b6HmApwvyaIoOagDAmdgYTYm67FSy6NE8wxvdlv2uqNC7Qj6hDjjpOgMgYiP
PrXs94QZLt3Wb0ZZvNGj9C0gz/0Zb96LVT5artWuVd3X6mnaE382EQbPFVcJxRdd
LdJrHE8GuqeBx9fxv9PuWamTjD145e9R2y1oP0V3b0xdwnwl4LVbZRI0qHaiKPQ0
Gh7nkkA2Cub7Qyw+m9kJ+Pvb7b1etxHWlsvkSV2qC05kAtheQClSSOTGIr+MYlrJ
nqiqCczvEJDG3Zs0cmPUr3fOnRxHFhgByk2wN/cmMKYAi/QIKWrCAAyr4FS8eu3w
AHQOQGyKd+zLvSJLdERYbo80fnTZySGKXa+kTHDzqth61uzfGrvjypIHnTBA3c6r
YmTBaPClJFwgX9MHnikXbtuZLlxckDUZjr1c2WvnvFY9Xl4XmnU16zzENgBeDDc5
dv9YhGk1xiZ9Sr79VMGySspBVT5H8lTaQhkKiulfDzYMNWS1gohEZHg+N7nhwkK5
xjl5QpGy2fRZceqWV2/pNlu4vkjE3d9Og9P0TiIBC8PaoB2L0RAmE/kosXwx+n+f
+GjRNq/5orcmpbvg6SA7j/wS1r3OB5gU+IhX3rgO/z5eqhkaenDaInOdtmVsCTsZ
bbuUGPuM8nT79+daAGvCKnsLrPnw95/shnUrcYUtVy+03eGuskewdzzyUpugMEuk
eSU9c2ht0ePu3Awp5QkAUq2TCR1ushnEdsvwX17Xj1mBehqsb6lHSDwBEFSM53GT
qFvg5RUDWNIJy3waut8gX6dUyRYTPHVLB44V/Eei0YVRNcTxiZ6Zjo1+vU7fkxLu
uB6vPHhV7KjU3iqaZ1k8Dt6VaxpYb5D/VVmUWjQGor/n9cde1Xie6aK+gjjcWtaM
RcMvPbmFC0YvqFNqfOK6sEhqcDrw2h9QtO/6cLydFyt3Oi9WRy9y9Jpo/Iaiw2y0
1R4rAsPkV1KIMRsqtBV+wzG7/0oua3ViLOyqZ//QUoiDTqfH+qrVkNc6+IZCls4y
Xo+vFsLHUQeguARJy3Uj6Ih0vwkXc0HfWWd9MJCGwYiHdPgtZ9t6i+Bp6zytuCDj
bgIDdZ3fQzcl9lQIFzx5xeaiVJU4S39/oSB1xGINloRb8u6HOmnbpjgfUKEP6r7c
d+JXmEIvhG+kw8TSaDrJo2WVlfFQEuBjIgwnr5T771sFhU+lbvATMMx2PqysSvfY
PciNTvo6Q9yiD7moAj3jfA9JYq0rf0yyELBAAUCavwckpPm11lig7J4i5MelV8te
0x2jvvYwVhAdE4eO0njBoUUj6OBv/l4rE2iMqJeoU2NIXFPyOd/xi6KSGK7E196r
XvGdfQMoXaKvqTHmL8zyMYeFkbVVt9hpzP3ar7E0csHY5ZfLeYFoESQkgGRVOy/B
ctV5isc07KMhG2lDDafXfpcqy13btvLMFkIk9qKFyy40wRZShOzJzsZ+gMi29Lk2
7HNG1Gtpbxu7l7QcV/cpkeYEHxftOQjaX/Rii+bAOGvbEGGq43JtI3EWF4Sk2jPP
joPBYz2gKx3r0MDvbq1vEDErkzmKsrvefNoDuMHz2rmLuIjqco55is3w2veO7NIU
4HKSAtmFptTdGwBD2p12HemqcREMnqkaUJzGNCl5mP8gNWqWAh8DgE3PDSfLgzX9
qAclyZayDbTUZOYiOtv3x1sNZLAC1oTaAJ+Rr4w46ZLRSmZTOguJ7E5PbnxF7HMF
yEd5UOYNnPIx1b4wPcCkuhl+GtdaIMpDb7Vks9gxG2tY2iBdSXtVa58d/JnGH9JE
84nfswXfmRy2JddQEGbHi80pws+Rt5d14qZlnFBYLoH1/84W6+j6xgZNG33/2zsv
yu2j5K22yNd7cVTUyaT9p/tjW39Q3CIZqnaTuf09xzS7r55NwHxJTFWV2UkfY8qI
0WnWvET/3IPHsJrRVce+d0fkkFAO14gV08ZDiBSo3WY4GH1q2js7Ph26p90XckFo
nPtstsf5OctbRza8r6TPK0UDIcUi8V22tYNEch6IXK4LMqgpL9Qgk7A0/HUjLbjQ
aCg8U82KEWyutk0nWWcOaiLOO2uvmAEyB5/fVdFrjZyHRlChh5b0CM6voiNiCrO7
d9vbhxUrKjbCP8qRPxH+eCQdzhltIvwwRuUYohkw0EKr1ry/SAOT508Jd+uf4kV0
Nk11H5A+85WsS3FfIUBMh6Ytk4nQPdq/gVvgFN8MAiFhBv6TSC/+cODAIxveThjJ
zG6X7DnKXBqZ6BXPXQepPHsUVNTGS1sFb38wpg70MHFtB00nf4fRzzKwuQmVWLBi
q5C0/ojSGh1qMe4j+izlP9TtRO4hK136/x6BO66nk90TLWYSSSd8kb+ePF2oroCX
IR5ATJa9QOKaLLrSdNqB6QKDaP23FMuVZ/+yVWTML1wWYoyVp33/Pqtr5kq4b8lE
aYxuHw9mHUWtKUMwQovAjlUndRbUPRyuj+6WFZDnsd8urjjdw3FJnwxSiYo13xCT
S22ap0lH+uzuDiPFkgZHpppqF6av3nXZhb56tvx+ZgKSXeRlTbTZcYmYwOwqBBtQ
PSmLCEhl22dWJqIfouma0aPcQ1b53+QCPPk8770hqfEP2OoypW2V/z6Rv7TKvJf1
zpSN0lpvwVsnGW40qXCxI8mCtRnMH9mC3wMNjh5+AVsWOLjtmV3c7sNlEFuCRhKZ
jQKAEzRNQx3LLARx8ipcL5Ajn4SRHElXanL9n0Iz6gUpVXOSt+p0MBGkpjcoxIkS
KSBgCWKlEZH5mT9Jta98nTEXPNYoaRxeBkcD1NGOdy5Ms0UsI/CIL+6aRdu0F/Nn
+VwRaI9rqk8cVD5Qo4JAZknYyfI40ZxsrY0zgRwcqOwsn7axL03hGOx5XvkpGEx3
d/yNbOGzs2pDdgGtmQoXCZGo2TwX9k8XUUv9WbBXtjCs3YGuGQh8hkWB2UekmzsU
MSb1iJ1ca4N2OTmJzwpO0vgCfKXOztoWxa+4ma/sJfWzZRMvi9T6grb3KM7i05+t
P7VmdDcUL+qv5brAaIGO5yzVElYU9v3JHKUcKX4Ej9py7GMIUcb3D9ecQf3nRPXT
mGRTArHtZmkaPD06D9JC65qQ9oLBesJSOLtAWJjoonXnh92DFtzwJjzEt5EpoNmt
Gz+kJjfEXsR23E/hJz8x7uteb8xK1iCS0c0Pi5Youn4l8udYPQoSHSpCOFLInKkn
EbAW+cK/Ds+/rLK7n0Gli2Hkyyj3g7cKdLQF3kySeTlkUNn/c/7TlbIUkTKa6mnI
AKaaT+tXquUqFlUUCrnb8ZVs0r5YK1LgKhpgctPXh8crbzDLLtXoYnne9CNLd7Hk
1lxQwcspXCAhKTdKe/AwJKGbdofXnQxdKL/zQ5X+rtlaIr7v6YkKHkMUAgupqIU/
Un/M1nRLq26wBirJbSmXRrbn06kH7x6WNA63fOnSUFXZRT5AP7lEqZ7JFHlomFnC
Ta04yPd3durPBHeE3EC61UV1cmcyctkeZuzrFUBWIzyypJTTUjLbYLMowa9x8gJ2
r3HFGpXHcRtx00qAmP0WwEMfBa8vx3XNDKZVznYtAIpmhNeMaEPhJBl+Upkds3sS
3TpasYFqzvY5B78a2MpgHyo5QxxM99lbRo4my069E3oSaEMguxhUBJ+EpPCvMNuK
9vTxHrCMbWWXf0e1LLBBMcl1CMJdDU+R1bFM42eMwYhTmJRlqYIPSWcaIViKYirC
4c6NCEo+bJRJPU6eDSDOiAKYPUHcUUAdE9s/2cWu0AWdyJoP/LH5e0cMNf9XjxTh
4+fHm/8YeaoK08HRANpVFpw8FwfOLgINYMeT0u8ojUVob4zEHDVboTheoUN3n4dz
U38xRT8QPuAFuKwKpV8cOGfznXwp2i2F2I+UIKSIMK0yIQ8Rb9JbAc8lTpUepcoX
XbpoFstjXy89Mi4BhcPTMW7BHWK5TH3hPJRiUbueczzZ2hAIPostorpy/c8YZhY1
Vn9IkiYD767BL+bnTGrcBzN2WmHdHq4JPu4RYe8HivJJq0B6BPzi7/3lb2ztTcQ9
ZLX2fiD9eskqKhhGI5GFyhcND3zu9y2mAopbwxMPVSfTDGXa7PyGruIvq5hjXZ8V
gV8KYJlloGVbULSnw/YtgWkTsd40J805LOzewF8PJjHa4UdPA5YXmUwNW/uXMCd0
R/nXJfHsuClkfbyo4aXFt4Nk8lel/4sL9/7s8BBdxaRtK32t0r9f9xSRy0oKp7WD
LtQI1hTgbKHg3gLIGUKKCtc2vtqn2BhSEXqFbPE4Lpzz/sp0zWA0MaUA2qDlKts1
XORT7g9axHR7djb4CfFNFxhlivj3mymf9ZK1lu4tw45+bcI6qKgrky6KeLX2pKhd
4ZwcEIJF4u4KCBUCVmiYFd3tCYc4ZjgXjebNaY70av7+keo/cXo4BtN+OY1/GTMR
+BcMxd9GgSnLM+GXmLfNqw5bt/0PRPUys3XnjTKy2DvefcraePwA1ucrSNM7TZk/
h3ibbyIVx0tbOB2LYkLZ+Xem2exbjEYC68KexsTlC/1qYW1N5mv7l5g6q8RGcBhS
LZXDLvjGV4FtW7JBxJ3QeAQDiURBqShl7O+mivqipaRE+960H1QvDU7iXTfFaH1R
j09mmif0LbpmPSUI9yWMt/g1GeJ9IhTb9x3ZhSEbdGFyCkqRnXmU3+rVMBX5kGq7
S1bFQ13KB4mfrRIJZoiEMkxhmjp7M6js7wu0ksBPosjRLXSRgs2/MCtKzkCqllLy
g0EK6rVmOyXiAapEQPSGXKw4Ps2tvjodDanpX7RxzAFZJsioVd0SCUhT+AZlDQQu
d7mLKa8Ex/YJTHvRRsKU9FR2ulxJNYIqvsX4x+02vrlhZ9tgPQbV1aMxqy2Sqex7
2gzNy9D3DXDnpU1pIIP2qJwUkO62AL2p94y+T4eWy01JxkKYXYG3xbc7eX4EEavW
VfaN0vC5rsHZbvFxMY5qwBbfdfJ5nL1R1GfhXDtg1vTBoy5tkBynjUH7i3gRNYCP
4TpQIEr7fhoFQG0FlfU67FK6moxPC8xNDebX2eic1MA7NgBigvmg4CAhZ2Ltjy2i
wPM96nqspnbqy2DQ8mXBrM2s70JqQewtl6SbzrkQ4+JNnn3YYE6erNmU5xJrKXCW
yCTkpAOvuQQxCnhNsSJoUBfxexBeKZ0SItwfLEY+v/5EMdVPf4KeAoauSsmp596s
SzRftoHAZ+3nfvIe49LJ2a8YACm3Y2lmd8WNv3sDeTlFEolcxV6+O6ilz9h8cbYN
EoBDzRgK+kphKjtkm9IahTbW14iZeYYgSCoaP3VHIrx7u+78lEb20SeZQwolvRI1
f0GqVX9MQ/RQsFhs5zQ5kzJFEXFrCEPeXIKE/wGdXAdCwqebNay4O+zTEzDtVszJ
YAOnbAeWeOPA8yfjX2ssUz/y0kY9kxMy/6B/IHYgKVhwI85oMZ+VcjS5HZg6A+Og
OBgU+fn2knBR4n+n/Cp02YxLR5ZFGeIRCuFC5FgCUJKkXO44yIUKuv8G5KGzSgsg
2xhkxTz9W1z5y+Nyu1fwbPsV0iAKtHhqp8NDg5BW4CWWRHflm+PEn5zeZXkM5EbO
7USUmc9YPtD98d5ApMyiouC408WZoOdXt4UxT4Npw9ct3BgTZPomnXZsHRjNDU8U
Nw444SEaXjEX2mrymQi4bIiw+EQcUyYd4wrqJZ5fPDeQh5qALKtvlF0hKADkKXZG
tNwMnNTILSxO/2MH8tvx+XQAF9xUvE9royT1UHkUdxGUnY/i6V5e6bGYxZ1L5SDQ
JAeOJ8jUWasZZBsBytRCIrcEMbYQ8JVjHJGCJLySx/hljH3bfR0N/8+oNJ6AjM94
Nkb+T03e9tj0od5O8IE4q1OdcXMo08zk3ODUOS+lVMLHq8wZNSs3BIywrCICeNFV
VhDSRd5RpE7MZwxHc7dySDOeBrRBRK3x8Yxu5OGmmqJgGV46/S35fKDGLo46vyg6
D+xEx5Y12nvoGXiY4OloDTGbl7aUEruI8nleXTCFl8yAW3H/eE/JXNtF3hZ7yvq+
egVaJhRylssSTcJKbgeo84aVU9lF5tW81/pXwRSx/B/UAI4a4TNqR0gxoP9OAXym
m0GBI2iDtavGWEtpRvLZj2+7nl8/9Wk7+zT/zw7V7Ni0W4eTjkiGq7TRzvLikIjL
KljC38aRhMioFts/YciKRP0PpNzZRHuXT4kOz1nkHu8xGGKMbVfBL0hQkp05K32E
DvWK4oAMRFZn+6Yy1auOZhiqCKDLh1UVcyFU7rYd+6TpwITzRqXTbrn4hZ8e+JUY
mTogtYE10G1f2LPCCCDxUqskjfPdJ92gVhy6wmLZYZOCtFJDuNrY6hnWb5QJvnKs
iQo3wdqajJHdIc23ElkDE+eqU8jFqBQ7BXmHWH24u+MVxV/gy/y6kk8IwUI2razg
xX6x4StAPvm0nqSor011li5nMghwTFPs8SPmMRC+N6KO2NRHAiLBrTMUXOGfzVHA
tXf/cY+vRjh36B+zeN1phMtDwkEBoYfPWsJWQiehgCMuCwucwl2JtM5v4XR9SjbE
u4QMkNzueUOG8hsUm4MWJ7RckvFLo4t1e9Mpmscwh1BKs/H9AYvx72Iol2FraczK
alVJbM7JPqjL+oa6NRT0LfoHERDq02lMXFsaYTqBCjQPR5zZF6VMcwESEvGytv1+
qKL0DoPtUCwbYhfl4nJcDiOhk2VWATtxWFNKpjXm1v9nMbAm3/ZOgJ8czyLt5rGh
W/LbPp0Sxf5+kiAf/rprWZK7iQ1+NvWNyagtrR4agjekpvdLEPlsi9UH1oZqpS2/
ofDP92cw4wd2y3PePazaNHq0MVbjv6dLbqfOuL3Dx6PiU70q5DYre4c7RAwBnOKE
2iJCdMo6ewaHWM6gaMyXuPGTDDBDm7dHeDZfWf745m69TDaoY8VxZMvVxfcP0MWx
7LO8kWqwILCnuPQAHaCNz2ogaf5fPAFFcCr7omHFAvN5BV8wD7TXY1HTTt/lK42/
2HulU9OhYknJQFns1hXadXKLaP3y+d/OKmgkM1AMvNmAomhMPIuE57V65z/1ViE8
F6yw0S1MFTVYI2L4Lb8WMnlAY7o7+pGnm0o/yJCBgTUL175iDKrOIXeJiJzh7q9Q
OTk/KgFsLravfZ2geLaWJYSTPHmReZgBG3ll8DZxfeqTYJ6UAIOb1LsMy86lc4Ng
sQFCaVBqAZT2H8fjdh3YomiwhIkn8q99RSZUevmLQf8jHZltjG/CAKTSI6rrHk8o
DxPn2b1FWk2B/3JR/gmSCL7z5uEaTAJ3EbSyZEpMGd/3t1T64rUFwU5oXhZZ3feM
lOlMqYlD5Ttuz2nIAa4T0XkXcInTL8gY3aPWd7pMKA2ph39dqdT79y0QhvP12ZsY
Jx9+Fi4yVXGgTYV1BdgI/JRo6RhI+YLDbXy0NuurUJxxqQK2rCpsGhl+h+NXPx7t
B0xltz516lIymys8ArJisB60gcO2tkUFWpVmCNov6K8ZhrTk6+59dq1j4WJRaHGO
25fQdINxNruD71z4TI3rT+CkrRm9+bTrbsSd+3Lae+pzqOhtQSiWo+Vo2B2/29fo
c55gbzGBKyq/a0Di7nMhE8OSfiFWWUfEnZFCrVN6TYw3vUI9gFXY9rF2hyvUck7j
1hct/6WNeXVnicWsmmGPnsaWb9zWPmhMiQxmQuX2Xo322cNg+69I7T4r8PwJy7sT
qns6ekA5D+d4OPOgvUhm7UFUk/mOhs6zfHsItFe6/3XEbTpGri4IQU6SLUocBar9
uooOMjBQcIZSZMVwK3YzdEK2k8EtODSLZX2F1vB0nVdw5/46p12RRBjnxMbha38D
iJJDrmBN5w4/j62zxY2vH1g+XnYDN4EaRfT16QsgHs7scdMDdDEe/zT/vhuYH7q1
/mzqbsflAcx8DyPEL7GSJLAKQYnjffqdY4rgXfNmgItPIl1CX70R4ftbNBYemlXq
HlVVhZzLVqvK47CNJYItxLJKcx0+t+CoY2JKdWYGqC2Svo6PntohoxD57AE6/ZWT
KNEAgU1Yv6d40pbs6qgotAcofadM0Y01pSn0dqfj0Whdq7zjxnO8pxpUFs8OjDHD
dwgjynoOmbkI7vUYRqj2mRoK933Ese//O7b6EKgqgWUz2v8frTf8s/62dimAEAHj
bDhB38QHT0rjtjOeNoLKeoefE0fIGrTK0knqbSClq6mZu53XxubO1oBCEYfn8Dsi
ZsLzhfk7x5TkkoIonBj5qbN6G9KxYmNTXw1+6Rll9xk15gHzOAywt4LJEvKbADRu
C8FVxfyMM+WRuka9y+RGFUs5cKW8ipntiyKza0xqYxzgdny8X5VksT791NW1Y23C
NlcehgOe+d6b3F7B2Q14nATGwjHKTaqYFhRTxl2fnz9IFpOLuz0d2gOkkPuzdJNf
rhGzllGo1dT4ng/8EDCkjWgnjjVGQgmikCLZJhC//e9JK0o8VAVdcDyw5e0y+W5Y
nYV8cWptPHkMGVOWDBpIwU6KfnBAiMd9Hrndom3rxeUaz5O5r5f2HkGKd34K02Lr
pOvkg5YFjZL2uAANtzMM6EZvoejkf067Ds9t/lR3xI6lv1ipqU+32pYk0ZVlQ2/i
C7+Z15GkwP7S4v1m8wqgSlwU3WbIvocEOGs4Q1aVRCPPLaYl401whZJ0y64lejT3
l5uSVaqtWa3vBLgPjV+1oTkSAtLW95VCKXZlUQypQpmd5XtIBF+RqC/TCQ3hkn0s
03ib+2p1F7rY/5li9u88ZELFPsc6nHRmVfB5gE/lXIxsCOB+hJGuQCXYWL8EW8OD
9XmYu9WbaoJsAOLTfccxa1uuuAEGiyYY1sgScCffNGDAdzVS93gLRcd9UPkZ025G
thhhLwKOCLt/uVKFqOSY0Njo3QcG4YCGVwutO6+3jvuEWtvOnAwMF7CIKzVkzBNj
BU+gGwqfwH039DaIdjf/EGYv+S+2tQbPZ6ahMGNwDHaMlAOkakSvfORqQD+efTPv
g4sU5wa8W9EK0uZrMEOmjzcGoAo4kNtJx1i2Vs4oh3okEc4mV7tC5LNnTxkJeCV2
rDEtsL0CvF7JBGMuWiFjsbTbE2LdCXt9cIqr/g6CUfi9smAHIIqmDspz9KouMYgZ
9UykrdwT1eiUm7jnSQfH46+t6vX9qH6AZvF9j0+CRBUkTye8NzwMmToQqVsb++sA
gJ25yiRc2bchtxTHjCmDYBTL9s8dtUkt9rAl6hgE6VlgkFAVXFIheGaZjFa5TZW8
CNhVQVhAjTGA1yZ2pu0Ck1iaKkEfzORTH9JOe4BdklqkEndry/ECkzf1Anqt7O6I
wArxFVJ4g5wfhaNhGm3RlM3G7gCZ5E1clbFgS77tFhHH97bMdnnlQ49IXxMMTaQF
HF+QF/67ted8+yM+VtkPiC2xKHs6wRZiIRs51NgDesrHt6b7raZtHy7XsMDFeD9V
boc6yyLxyEi48ab+5il0qrIJfKmQcDaDig5iVGTVsFNyfbZ24Vmb8ViH9+VM3/GJ
I290uEjSCJ/EMBjGJh5pmBjZqs86B25MtaDqydHBM4C6ivPBgOreI9g0Yp+pq0hw
H0dnSROV+15y5c2W6HaEvczm63NHsT9By2BaSc1AB2XI62943Mip7i2Hdfpqv2E1
71f5/DHf9EYdZDo/spul4jgbjSqGQsoehfwIawfT52CfU0DuFB0yHoek95Q5duqM
mG5S11aay376w2jPFZ0tni/Q9uFvSjC2xe+f9TMLv4tquIiv0+ikjX80iWVhPf0V
zjdaqqWlT31abdS+U9kYejLcn2s08FQ4rY0ki8HxW7jF68rf+8oDEau8q90x0tuI
PR9zCfT/xzeWkORzPXYzAiW7tRz9t8PkEBB+RchQxpslGYpLYHOVmdyq4nFQ6mCO
XEFA8t59q1Szl0hAl/gJbhBrjmvea/r/MW+dYuIIUcKAMwssDAQvCDDrnrRVw+Pd
6MsPlUggQVKjxZ1qUIwNuqAS4eUhG8NwAJ1Ks+Lpjuat8XZKoCAC3O0PC5JkQMfa
7DHFhI/y0gK0bmCQFhvNwiRPDphjLSjUiVKql8E6MqDl36eKJVpAIOxh4F5llyyb
2aAwjIrqVFOus+IAh9cTwaos+MRcxrGHzeN3UuaoPOYYG7zIU/V+qIIsMnIhsE0A
0NeMl+qBckqubgxqd2E8NBrr6RMyjF2WBnx/n1foDUfqT7KbIptI1z3KgFtb+gF7
nbWBRt1IrmJXj9D5JmJPQa2JQTZmRR5Ve4hkWbS7iBj90dmxjXFcnzufNDYKaqHC
kt4JIlcURCHnNeGow3zi5lWR06GVmlUOLuZkXMT+xx8=
`protect END_PROTECTED
