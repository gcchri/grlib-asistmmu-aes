`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ptIGarqVSREcS+1aYfnSj/+t+cZWxutd4F7XgAPqHB6Eunyvh0X7WXtvy8w4TAcG
xgVV3mW1OeOITVRCyFI4l8MzwD919irbsIhqJSfrerJiPxeoHSaY9Boxqr78ZviV
+iMO+Cq4CIK+pJhkEP7c+6Zcnm154+YmFBFLYT/CTRqBs4S4DS3lJXa+PwJLOM2F
ZBeBJ8k5N2oqnb7ZnBEXLgQ/uHiBrMG4sxfF+d80m00CKzexD7mTpQs7jIQllaNY
lzfVqkwpkEmxsEb55PVQ2NrFOS/EFRRgzhvF3tZjVTmUQjp+r3zWsWtmu93OMXds
FLKge3+qmk7iIRT3LNIzu12IBcXqjQMNfWnUTGcDRutiBa3HwO48HXn7UC4pmGUu
RsoIQN89gUODvy/daJ/BPPu7BsXtk06QF+S7QqVagqQgLjG2KjfYK+lxpdwWhv5v
FOS9bnGhS2KQ3iQ+3o50YqACH/lbyKoXQQ2oc0oFRi4=
`protect END_PROTECTED
