`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cbTepWLvm8u5JnccSnC0yKFWhd4TrEZZp4Z+GtGXgKJpxon2Cype8CCvAZictpKW
tSUnBGVMQRjricAsf6lbtBSAlFsby6BH7ibmqTBlookgXocdiI2AGuUenYZBqyG9
sYDkS/U1r3VhgHF3K324zmnn7rAiH6AsW1Z6qvyYamRtELeiCyqNNcwnqM+qRXG2
vNJ5DcKWHgrt1qGZdKE+ttmtNg+1amrbhYahN6JXA2LCcdWbh59IRqtnjLv4kYcw
vN7MzFRKsH1INMVLViDmulojyu0JybrJqTpQ0tV/Qe1Mqh8aMTDFGthD+SjdSkS1
UUZXEYbBjppkfiIry7zpf5wvWL0lWJenc3SfroFLNN6LikQJfMFf2kU7nyG6zoYU
uyfXAlXTvRIkULzq5f6hmkEtq3NU1TPRFCcvB9scGlcmrYT1OkeTqXqhggENEZj+
rrhUx9NDQOuJUB0IMcuXUJ0GQ5NDwIATIrZSqdCva0uQXeatsUDhOT2lSuUktA/n
49i0u5zCbV5Rso51v5d6HzIc5i5GMBVN9jWdtk1x6x6wtAZYHI5jbMleQKtTb4Nz
Srmp1Q8OmRBSa6LEx6QqeGMU9SpGNIH0zDokt+E51520LLvMpug+PCzYmdobwYtX
WP2byPvGiVxP1s6kTNKbzztowbEdNMYFQE1AajB4r6RXisHn/2dGYwgyGMbR6Rr8
HyyiefUj7ayq5AjweL6YAmprszCqgK9SxYa3LtO9CMWhCRVukpu+OpWve+Oq9F/Z
KmXwgnec1QcdtXmL7/oUWAVafvX0cZrReAe8nu2GDcKWgtdDlBws7EHn1RHcOk2+
q06XgjggdH6fMoPYU3CAbUYG1U6m6gEyK6ikZ5KEl9nBepDckpr9g/GN1gxeWon7
85B+aXH8doVRAc/89DIJTU3bmvQYo3SdoVQvBq6V7GLCbVqfVx3lwKq7jNgQYu61
kYfzvehvTEmU3oVZS3s3lYBwFGrrGF6G7e6V0B2d7HjOnDylbmCeKsENYbTwAGMA
LcQGujwiz41U06TWdPtcLkjl8oa9xY+bzeaST8SxpnenlKL4rq3SwNy/P/oG5v8C
3rpesVN9em4baSJHP+Ii3m0/UPu5xvkTSZNEe5zfIZweqOGoZYlRWI/IdOhUY+fW
y0glM7q8+zuQ0XX8ITizT4LCYsanva+NbPkvggLBxUGHJumqcPNJJb7ItuXSQGma
lt33+tUyoRqrkxxaD+Mp4AwBzk70/rZEIDVfdmt3VeJknVPRvFXjyhd/pEonpeH0
0s+yR2WkJFGUHgK11rW1qeMLIf8yGSKwWKiIaP5vaCDQezF63CnBmJqkbNqFQ2Vk
RizRN8M7/DHRKnFq5a2Ky89cunSxeuTc2wzBK+XAeirTALdoeA+UHjzLi0wHwGoq
zsINx3UbiQpp+Ig5VaMJhTYiLiGpzXXNTaqbTM3VYJ7Xh4nIP4FMggVe4pZHKqXi
xnFOn9O7d5be7Qm+bacOA7oJLkki4u/rfcRlV9qOpCeqO19o8QN72RCdtiG6LZt7
2Yd+cX5cHYbo8MHpeupZuiE/N8tclR1J4uxsWx3Vel7kiy8IKcW7xHw/hU10bYM+
l/yrYvGmqz88SrD7zgCqj+ibpt+eNYs+HuiqyBsaqlRPqTXMMfQPwejMLec/RNtL
1mH705r/8FfWk0+Xb1sJVDRbNERsgBItDIMwfflMwvC+zN31sBnwKGVSnyVME2nC
BxwzwG/sewMOglhEApCWl8NEMRdW0jfPjSFGgeiqOOauQh+mZYbjOKmKGZR6O7QQ
R1zVSb9++fSa4wdsPaDvrpqI4irw3qHiZecXGA32AhQ=
`protect END_PROTECTED
