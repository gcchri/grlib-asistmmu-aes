`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pL+qs5gJRlr1ullExleAmXJfgWuzDDnsrVT9RnB0CQ/2nSz1IT2Ve/QvhvVbg6yw
LL39KHAtJmZqnzVVWehKkJs3br5xegzLEQNBlcDapcQw7ygWFr22laO2Noxu+EkM
vAwHHQgOfSh0CNbrmy9Tgsq8WDSKxha+T8EjDsQ4HUQNF94ky9LEZmzUtDtreV25
Ocqzpy2pBvxJQTPbpLoOkEG+LoaqL8e5IvjGjKJXUd1D2oeAq6w63pfyjO2d6/So
qju4eUlo3AfJUOOhRj24TvQr/Y4v5AagRZ/MuKUNVwd1K01act75HpABQHtI25wL
R/4CiO9nddnHAVWnOAzZl4CbPd+6FIRCJC0AfS12KegGFCv970tXOXkomJyItrwu
qZ9X4uRde67eN5Tq9DLoT4T5Tb/p4zZZMCfgcIu6riw=
`protect END_PROTECTED
