`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RhXrZuMq+AADVjVdo0deX0wYVUnqfnDdgLeTfk1yMNn1nsM9JMKyECRi60m9uxF6
uxG0fNkiHFYj3mRqxQrPX1EOnlKypFfh2n4F+x/r4C3aW05nUJ92KsYHZvqGcMJn
lmd3PLu/Kwae3KGz15ko+nGYVrpa+pQepA2Ors0F9XoGKa6Af0neoppHyVp5S0Ja
oxfrkE3BCTVESxFDU7zICYb+IQp2vMLaODZaL36VMxzPzsUyk7TWo9U+LJriOJ9A
VQkaq4PzyqZbcbhEcQljEbFoZiN6hMOgtnyfOJwy1gjNf5Gb2XOZvg0vP7BfjoUL
e22vVkN7HAjKa74hmStMxkJB6FW9fEDmaMmnuY7Lapn5TSOrKBa+iwXyp/fT1iJI
9ptn4wEU+CIdNVtYr8EMiR1sMOkGxeM0eRFG+zuryrh17tFPBVH5Nawiyx64RDce
S223mqyV3sHdww+qYIfGhZyd2Qg9zgYddCt3AgRpVXoFNy0O/Y5AdhC6599/Xf8R
VAI6KD39NqeT6+bdHBPLBJ0bG4sTTsOk2C+XqrPUohGQzYztwuy+bBSDENKbrZz0
7bMpx23XvV+ws6mmSbkzSOOOatQn76A5BbjYrTIQBQKkjjiI+mdFFvpVYZar4eCB
aYegMyeAkqOBXEZLhwx3LUDtub43MYvT5eoT1E64q7aivylnZJYk/GBgsq0f0ecK
b+rQlEiHPV/t+6U+4ACer6ChSzWrlw9l41IhOZ/M/8q1DXyW9JiT/RNFJmAs3TPF
S4vn8OwA4EtWqKcsU5iYfQ==
`protect END_PROTECTED
