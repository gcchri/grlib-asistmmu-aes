`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GMVb2dliexkeMDLobF/ZeOkeRsPY/gFrJE0fiCSuOIkqdneogaLyJEzt6bOgrMnX
AZ3dirud9rye1IyDoQ4dM2ERY4nnbGCSTaPOl/HQdF0nvjDciDbU0WPDZA4RBL6t
303HPshJRRRWiP56ZUepePS8jW8z0Ksq5gFbi7HFVz8E2kmwCEfn9QeWvocy5BHA
uL2DdCENgsbEUgK03HR1NFi1QaWMDj4QH+cX8ithmrCXtNXiyoEPlYsk4NDY5R+P
Pk0eLtSg7Gwu7cbrhFNFY7ZbY7Go60ROx4GpAHt9UKvp84v2/K8CMZorJ4RvajK3
y31Z77iH82E8ZqvK9kbevG3az2TU/aqeziN5Xavm/A+Mwmrci2m84+qDRxRb9cEm
kwy+EQZayuBEN9mpiLdHQQlLUpnqHYrO9IJVLRgeP1xzNdi3fH4Bq50WtMLLOlO+
fPId+RAXWDolG2t5q38zK25SyOGxvqIgtmJBOA8WDVSO+8ZEzhuZRlMBcHZFItfi
NVB/ADNMQgqYyS2YRG+rHP1svsb3jZRxTP95uKNn5KSnx0/aG44ogugUVQ9D5aVF
nYW+vTyHU7qjnjC642spwRMyqetHFJtIPh+tBCQUrwq8j4GfOYXawp5vqz9ujAx1
+rICP3H07mAxcruCaO4mk8h/9BKCcVVDE7MP+jEfcl221T2ULVxGZEwK3G3evg+D
Q0mNgq7qzZop9mpKSS5+ELVUO77vT218Im8KOB/0D5MrgcxRwlbZuG3HEIpMBmL5
3RJ3Th4LLET2c2ss7cLT3QTbH8sA7lqmEBH7Pt1sd15A9SubqmrmFDf+ZBwL71BO
LTB/8fG7a6de2/DJp02cZqgtlObHUSd2p7N+Oc/IHS2m2eqDEWow0c4MKNzAAhKl
tbqsM5d9rhI/NQZe2xYsVXInQ41zwwoeNrxvJWJcg8DV3ZhtLjD9AzxF5GuOdvUC
oi5JE40fHptphUncysKuvTvWLozqg12heap5UXaANRqHUJBsgveZXsu6WaeRDaaF
ubHjF/1nM4FlayH2AC02XIFkwM5Y2d3i6zGJMXdrS12jW0SqMoJ6bXF324+iYd39
skuFolTzZyT+QeY41/qIK7xO2j9I1zfuUjB3BEr29mZ8RwdcxwkuJsLmq4UazFOw
fIhU8m5roKh2k/D6FQY4mRT+WcOX/AYb8K61MRT0Imxp5HlLFlgNfMoxNF7jxHHr
/G7KRkl/f8GYybZhtAxFPyO2Ngzd+3muUYgZRbCKbt0BRpVuWYsCb4pwl8SSUrb+
j/dMv8LAIvd6z1Ty4nOXSL+pwXz6v0HHoRjeWrxICknAFammct5+nWMJGIPNRGEF
s+VGeBT7/gakpB0C7MSEUvd9l+Bp5M2mqxvL7WABUAeRrNrCJ1vOoU0PowdZM/Dm
OgOoYfIhJbLY5S7HoGcLxZygrs5d93039pAtqZEac4y62QZHcbCCaNfO5B58hTCM
Xph117SmsTW+2BKZdeaY2BMaCBEd3x6WtCd1OIfevUQw9ZEXYyr2xMpnNlAmAkeS
yKRmKSAVJUgy+zEy/w5o3wHdVdOBFGbZCu4adVS5aGe4Y/95vSzV9sXonwmb6T/3
zPgR/9tYmde+SOJJQqLCN58nqeGxExGrk/3cSIRHasZ1q5B8YUesvW1cbGRdUhvr
ak4+XxErbPpaUQg/DNn1z5ForCdMkhYczqEqgf8FxDUH7FmweQnwn/zjLKVDzkgM
vDW0hXMxRF4xRkHig4o/ttBGWC5FdsCRdLPgbsdvn5lZf4o2TuE9SZ5+ebmG7m3W
uieFByS3QQi0/w+WnxklSNT7GodSv6u17cbOqrfIeFFEmyohkUAlWl6mc+uBWAqZ
ZXVDAjgGEkDYK5g94l/GqnZ1LWo0xYk5wp5LvE3Xjm+tcurqVG27AM5b7x7VB+LS
GYoordr1bM9Ln606diYYiQA3fKn0YUT9LavYD+vCLtEfMhvALKdMm0pJ4eqU2voK
3IJdnhxvkgXPse9Fo5PxoIbn6x+vLYfg04wdZ+Ivb+KyhjBEpwyPnkxy/AhYfsXf
To86DKEK2C7iNg+hlTb0Mh80Nm/Fi1sHhMjWDRefxN/GKWQ7Dcv9aqg+4q9C+PDd
8ayky3ULYHRmgpy7j0cV+z2wE4b/OBW7kHcvm+0U5R1ebZQNL/E/COuctrroIFnJ
GBb4rUwfO7kWQuLGMz0bFT2oCDjgF2/wmpCAUv2EI5IpF3pmQEAzOLpd5tgzW7td
3AKM56ir0Ku9XzzR33QUUHEl1OAg4VGXJVa9cPkOKe8RnURnMQCBAmJH+7jFPJTb
PvRwBYppaV8Y5K3LC+F5Q1yg0+SjjQHM7f26zyI6/RjQ0seeuBuIqwQDdO3vzX1K
Nkz4URAT+cYYlo7JLAz38njDxlG1IQ/YaYzWaMGGPyWZGbM6c35OxWp7z4slFuS6
6OREXL299kAORuEXLKQLenlnY6h5kTEiRlr5/4+K6Ml3A8XMieiK0F3EjSFkx+ij
STfIGS3ftiMPbeLzZukPlEK20+uwYv1YFjp4cYrMIIfcYNI7bZ+x5PAtrZKc2fAC
Ic+SCa/Xh/O1YFcJcskz62tUHkZj4d79GW6Zo18b+MNvZb1uQWr0qi4SsswWhcUg
nRCyf10HvqeZGYRVRm8TvPJKGOat1nWwn9L2SiX23mItRkyiFdRr60zAnTQTItzC
0a2GdhIYdkQ6DkSjfufrIDosPiBN/OhQwcRGlooVqza6xTm0kR5pnLmMqRkt0XaZ
vT8ztS1yObYLYoeNAi7cK7IphmQsCkRAnLcAKuAKDFIX6EY7/+zJzzHAdkAVfsR/
rRjPPv5GEpOFjwTlk7xf6Q6kR1M4UtNQdju5LM9+QqHG0I9Ad78fPvcbBwotExfq
ON5g75VFQn0rAygVq6EgBaELb0iCWrxBW7ATCl/6+FvJltraFww+SzWkdV60xDQ2
KTWOUJmzojmxhSNa6mx3MY9GoKx2sALrz39G5IsIfAIXxnCeDUROaaiXKo/hBClv
h/xo2Zvn3D0+LlgabadBKfutD02WtjZRZ++fVPozx6iFPXZ2FfvGCx3lDLvjSCEz
uhJ7B/q+j6mbidVy7PKaqXs0EPr3JUwyHoPMeu2ukzlfP8IMw3y9y75r9vKYSebX
KhUQf4yIJmcSUFAGQ2OGSwRzl1Cz7zpxGOBphhMEe22lhHVges4TJkgEAYvHgAd9
2gOPPpmvDaaICzjLhmd/L+IBsajFEKGk5Mix94ZJwXOT2pzbojjDAygxaoApbWfk
YNflvwAbZKxvHmUqpHoDvxWDmsfCBJyDHBuAgM920jkbkscV8oVNtOTsLHUKfoap
FrHSw5v43rGr2c1bwv+gV6V6Q/Hefn+eH2c8Mx0KiLkOdm4x8s1qUB9N5s8rKJD7
d9nl1db/Zcaag7n0MuvQbT71YEeLY+jRrgJkN7WQ/qh5AyJr/3t2mWWSiI6pyLtL
kQjmDVhUFnemW23G0uYxMp5uc3+uT3UyCqk0kdLdyJ8z4u0PZtv4Up0bGlb8ej59
N1hGvhOx86/2tvSWMQIUJrtesIfj3ht7An/bfsPhlQA7XICUs+MtagJNaETt4J9B
UXCSkKq5K28z5f6czdxPWxsQQt/ODSXb8Bv6GSlBLnarchAE7szVc5cUOviYlaq0
3aKeJ2xYlkwDocKtq/7I2uHBnZU4ii61WqUy8sfn3vWTEUtEK7GrQRPfu23y5kDW
rrjigQdaQQduTrQLWi1To2XiWMDP7pPXPdIypFPw7veGHH2Zfbd6xJE1bvhl4X2n
mwXW1ZdbNTv9v0hipg59ye5jzgN6jr4zo/q/57QoGi9l88pVO6QUwFWmCOWppFAL
CIPfQyEfy4A9UtFKEuFZrHrbdAEAWYSjK+GMSWIK1C4VUEsrWb23oK5BhRKsg8DI
w+yxjbJ5lYRLywHn1G5wrypJHwmWhn2MeTcobTyMTVSOj8Vo+gvC/euGFjtpMfMh
XfjKLG78s6saP/Du6NjoJAS51qRcAbrKEz5ihJ9g5XDdE5Ai3pYbe+um5kyq15T4
bHmq/HNZLxCKK9QusDlhxnTRX4xHpeWU4NJf9s+UPUlrzOJp4SbsUZHg5O5WUnFd
qDhk5a2SKJzIDFhdFRTCqww5A+VpxIW/C/I1LdG9T6VvwrSS3vRtIk5QkRgJ9e3h
7nka8wzibC4uS/zTxx4lV0GdIvWZuhpsH6dLBj0HJAgzaQebFajMqWP1Dn5sebcq
AwXHnf7fPmgEHuHGYfEPlf1y3wdvaiMXuLDnvGN0HhyEW+8rhXWuviWgjcrR6pYG
Dlh0dHEukC9upB96T2ZLYGBe6rpToNFJ3kZaUYy04qnRM+0paqb8L2G5xE8/4Hwy
1k5goOSZPdB607ce9BAcGGki4Jsw/n8JS9Oj5A29ONUDMU1xwp+Wbiqildg/IpEt
TsxRbcxaixkjXoLwgRpcw5ZereF/i3SFt9kjPrMLqFRZH58NHV+SgeLxTi3wF4or
UVD2G9BkbAvVfBhqGelxfMPNoLI9Pyjie+OlsVegBB6aMMNts2N9ww9nQuOlvFCf
Ccq3pW+8/ImkBMTAmyyqNZr7lMiV1NdpsOEe9B4BOMl3g3z/PuKuOzF8gG0iExE5
6xPVbVwW88KzdISmeWUgi7tXlgmAWyEIVCgXHy8rVoXt50exzA/LecPjooJmowdv
FRMIz/4hAmAHT61fPHFcbZDNh/Lg8bB5HvoyOqkYdLKf463GzoOBLAKWoUKjc8Cz
CoZCr8b38Rf9Rfhnsk+T24zC4gMQc1YOYy1IoSeLVTbZMocKaO9XvQHve3Ng1Wq4
lXQuPAQqEDjO8HI8Cfzqas+cFFmpF71FBosTwFlUQhUQMIF/Kqn27+E2mbYNfOfY
Z9xFVtClSwrXdQPzN4+taPjnQC8xnZHwSnMBzZwl7YKX3KJRJQlRDvrc8R/iGXMP
dCxF8qJ8EVZ8CIhxlCnJ43VIFNuAsXqLMeAmffThhvYX0t1st4+w9iRCS8Dlqh+1
GHo/2AmAJ1syLxUccnGbzu5qm4r4yraShtY1nVPcluiSeJIb/gMdTRpB9dSeP6Lf
3ypHDmvb++sJHvBW63NmLXNLadxCp2Il0yTlU+gigVgzBabZjz//nZkfuCtxoPKf
rhm2UjRmqZguWDKKTxu4J22VFSJOZ8Xk/VAIAJO7F1zVu29OyvUBj7c535VuyqUN
8/toVpPIOaik96PRd9hDq6vJt8d6ppXE0SdXoaWzSgALllTv+VJOUoh4WHAbzP8F
vkEokHWqP4UVbOtuoN8nKYwOvjOUlPnpdnWq9BBrsSZCqMb1+V+8d9IGND3hNHZw
wR/F77s+Ofg7Livjk2e9TFdCMpfTSwrbzKeU354WDoGlok3G1IHCd3aAydVZdGab
zS3yq2jVfPcA2bLqbnren5PSFvxHo7/lgxSdsHWx0o/8CgWSxsLZoMy5WWWDjWLD
pl9p6u7UitOvVLY1lgJEKtfCKik45IgwGhmOnW8Vtzmn14EtV/QXRNzwkHRm+XtI
G5+/YATqYZwxOZw3PCurZas3sE83eSBF4Z3Vrj/cGAi3zLGtVrLUYSDgdEysVQLm
WYSKlvJxNnhWBNB1DXhBCkRW5rd0dMFGYgoXXyRgk3ki4pFWtFXUgoI7naBITTdv
lq/22ucLGMDIF7cuHvla+CVhQR+awlAO72FMzbp1QjMimEztFpnKJV2abug7uaiV
0IFg+LMKZhSIKW9PNNdW5SHXd25kdHcLcWmOXc3RbRpsRUBypm7b5EF8f64u8wLb
Ea7ah4fdOKJpAAj5/+MBQRlQBWMI7acUXXbpjRokvq6c7KInTjF5ehtYp0c5r8B6
VDP3IXxc8yxDzVf0gMPHdx57rTfgi5Ophgr7YviwstTNXfw96vhapgIrbVyysD4Z
IJ35q2Bo3Q8RhNchb6PTbGNBnAPioR0BamfWZYGHpNcsIKg1j8PZFaud5P+spA7f
3qP2BZOVk3JYp7OzSxepvCEEHWQoQIpyVVwTssadKwUK0X4WbqByA2R89SdXBz/t
iMf/jvOznLGT2LDks678NJOgtwGWGPjQsklMCyByfGVJjmHKO0+Oc28EQvdUyWut
v0MfA6dVdGaITo5IXPH5JslSPdVzfiCpIfm52vOIa+6/XRDc7kembaBhVIkI08Ua
zirw/9SGziyaUlgdX8FhtUezOZTYEQmU1jyIne+m9PCKiUOHg2aw8yE7+TS7D6la
hqusQrqwAMAhFuaacdw3nKKzo7JSjhH5u1Kd+TMqS7mLt0CfGB43ymgVBIKeT+BJ
juvWqxv7fqOGWuZpJwT7rBDucQm+8x8J0TYLC8W/oUkyF11cjktGTLk4AJMMmGqP
b4y2FWlcSGOQT2+kVVvlaPRtVYK0QRpaLOylTXq31l3QzgEnBi8rmH7CXhsB/Fg7
52wKQGAu0ZYGB3P1rSq3PtDHwqvOahaG9yo+dXvShPIPu+Oc9bvkLXT99dA67VKC
qwappJPLnnMzzfV3pASVdFgHZEGTiE0hwlOkuohF52BRgdpDioKcVx0/PVO/bO5D
TIYyZD2SWijHBUjNTl0m2h/ZBudtmhNAmYW/pvqO1Nfeaj1gfO11nwrVLXM3GwpK
fWfSbYbLSHpPhE+/P4PjhEYm0a9kkUMeB4OZp3jKWFjqI0J9TmeL6Wp1crvAtGJw
iX/JS7hh+gyZ+UgYJ7EnJqU8HXjklYjiZGS8d9PGaij3b6Go6ErFgcIOHJVZmQrg
ffHn6YrUkqJi53B8eQHPpt3NxEKpM45fculzlt+579LOuMNZjhbEetHVl1VCJRxA
ZnduwdItGTwMA76AoSbg/IYLvWgYfcLnKf+2+7p0JaAj8c83/LnniAyVssCKOMlB
dmsIYQzEs2H6nf707j09wjRAAkyRvkjtgHyW5DLJkC629RNglcD2aIZmwPsWdgaF
mv9RRcTKNKRpHLH0yzHBuG3nygl16fCxJOs4LZovNXwZBM/ooiBDaEusLHw5loGt
Rv5wsn0CHChlRgFfAL569qS8NWJgY4RAxTfEE/sHlESMZfKOCUj5r0awc3mpAjGc
x+Lp0odQEDDYtBuVUPR6FalMjkxnyBt/SA2j72KFQU/puK+Tkw8xcTqiBB6Lrk52
IvQ2KSyn4It0k4dZKB8ga1SHnT0neupglSmb2P6rQdVcJ8D8PnKFWBSDgg8+V0L7
ecwt8uePl7Toku8QcRfHHqeTlzlnflTO/3F4ctj3tOExhku0Aa3suZOT1Zde02lL
AmBRaemDAdPZc4Q78llDRtofDyOPVoGNS4t4TsPbraDC61s4Aaa1lMfS5UEdP1+Y
XXqrg511LONXGvyqWha0DGBU5LIYqNGslg+2iwuOvBuZWETQwvGh1sM97bq6RRJ8
zHjYAjpua0UF7fFJ/ilMtIIfhBtDPVRu0b5Xn3Z6WjKZx4q5jOvLOHkxwBKpKnsP
AQTxL1jL0D2Au79qVmFoQGwP5pxC2rvhbppyPZzwWieJCEkMl21vG5cwY74dXiyM
xnoJPPye6eWG8UBJFj4O/qUUWgkH+e5JIzFUgzmtGEFE6lMttdHsq15T2g2qgFC0
qCuaXiS2c7uEpyjGyNVvee/Sw0hEoyRbo0fvkTYQn/Ci+4HbWEKZ0U4FskiyEI7+
09UjNSBMZW5MMK+WdTipVb9kKHxu2/4OgK4IcvllEqcGwrf5qhkSpLa5xiN9xFS8
t23UBrTpw3jM+8O6iKLk1fRvDvI8TR36mrr3PMUIDEV3E00A+altvLdZ7t5AFZ1w
WCizb+pU8fdpXR3h+vJ1t9v/JPSPaSh7LwTHzsIaAJ4=
`protect END_PROTECTED
