`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AN7rHRvMfzpLG/wqct4h9Jkn397fTSf2QCYepMoS313SO2ejjdD3nQR6mkdi0Q4V
W6Dp1is0tEN5VJJhBgfK/YsIsjw0LhDoF6yhbXDqprXCcxyTNN4hLnvtEvmzHdpM
q415ceQIyBaKrpBD927pPtC4S5KptdXcZ31zErv4AhpD3tipOScpp+4VIjmy86j8
2hEJ6nq6cF4VVhgZ5mr9w/E8HklUXhA2OdKCt8cNMWR39UMeRG2E84xz9TXtJCGA
D0yvdYhfm+RVSmixc+ufng==
`protect END_PROTECTED
