`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9xo/KLiHTeQ3pnxg1IIhe6muHyVdQ1tYyaf/HSRXvS5jU7NtZ9yB9YgaIsnGpVum
9bNKWV3jDMtVYOoXXSiQeKBMAc7QJhCc3F5vY6bEdAuxCZJKHYskO3dbDDCZfRBU
AcD63HTXUUSg0msEbJCaGd+z0YNIZ40RLJ3yJT5Avk0Fau1cC29gHl6gQCWiPKri
tMLsObwUBmw9Oybv6O77AMa9kHLt7m7k6eGM2zOmratGUQNn3EpFs1zBoW3JeIPn
9qtXw75Q2978JDTWDalVrA==
`protect END_PROTECTED
