`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wTb1t7UtOzJPVgX2olGU4n20jC+Ghq1K0jKHCiMMlC4KdNpYMTGzMcRucXbgxYQe
V0c+k6twaoyf6WabyoRyA/rjUSrJgqT+hxbKW07t/zNgyNCm0y/CQs0FpuMleatE
h1p71labSZDqmo00KCQRV4SiRL/PCPhzWDWv6J2/nSAbW9i690y9bML9SXvcgpbQ
KzbZkhmXKl1SdOCHkuLZCrh50wJSeDjiU8F6ahXQDMrKGHoitI/lUs2VZGHmQPP4
MxTkZ9n9SS0KRx6dhrO47+2zqNkAvIc0qbawYZ0ejZ4dh7mVe88jkLueLZiG8AeE
JGManr3+fIbm8DH3vGZPwZZreoAHlh+QPZu2TbrgL9seeNa/QCpKj9KWIWHr+3VC
Zdihiznr6fnz1nnvZz8PIMAUfGsiN6sEQa0Ff0SxmjgDzdXOFLbQIQ2ojuSelglX
epFcPtA3/1p4b29d/Ch8VNB2oMo8rAoxFe2+91iWEcNcly8lUBVwi+zYhQZSUt9O
hYFprjH2naOBp04gB64dcgwbvLpZ6dGgrLD0W8jVHK4=
`protect END_PROTECTED
