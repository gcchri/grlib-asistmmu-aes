`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMTXF0H1wfHThPAlFHJDwZT06miBshmoHp1G1CimivAzbUSCt983f8TBH1OhRaTv
4e6N1GmvgGv+UMO/WsOZ4UzjTQvimaXtv2b4H2uwFKfao2ui3WA2kELQ1xJ6kC10
dw8rTW2JIvi43Mjbv4avUvrMICLAfDzzNd9k2dT3hbWRxPioD6BZHA4eFGxx9gIE
UODbUnEK3oYMH41S3MYmVyIV2TxWsrKadrkaRom86yYQmzb6uM3BNCuuBejUiyV7
PIwyL1shkGM9sR6705VCHC3fkXU4v3TGRig84piOjmUKiGup5sbeaVZkU6x4ZHYm
3Lzl7Lo3rVHaTKj7kmVXTOe5GFTAp/NihbqXipQ3nvT8oxWRd7FPRmadzpYpT0YF
NPuOWYloP/1yQto483R3PR20tsh93flubIyAhNZTM5kKEZRjH6Hp54dai3MKRokq
8uQlYZk4Caw/x8+LUNqfR33OBjS3YCrf/1zBa+I8Iqf2ilhaowF5h0BNf2e7zqUJ
fj2EIwaFWKzCo+qyO9Ohe7MdbRUbkA735mDY1r3ai0K1jzyjVXTpV61aAVAyKAJa
Ooap9SFcj/g2rq10UCLglobOvxxoW5vher1iG3vHPXQIIibnlvaP5hQGdXtbLN40
ejxIm9Hlr+n06NxFxUfRuiYmmmfA8Qz6mR0/mQ6rOaiKT43COvkHaCZVpHUmK+Hh
jwP+VuhyqYcovH2iF5zFGXtRNJWUa9xeNh0M0hhGxANkySU/XG4g9ZUVTbziV+u8
tOTWm0t9y1VLWrZbaN46nDHB80/GqIdgcPgEfOJ3+sgbWwhLHk6Xikm4EuxtF32C
B3QLth0XTggwKNcmXT14zA==
`protect END_PROTECTED
