`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nhWbDYH9LL1Fwl9wYVgWpd6i11XF3qjAQaqtjCytkSLUnEWvcg3m4GsUxVyq/ArL
2l7OCKuK7iUA/z+1u1RU+KhkGC2oaXcdgz6f9y/N7r4sLJH+l7xwgf8+ED8349hb
hZ1gjwF4ParJfmEVVZ6bi2jtT32xwEZ9s4rSsGeAa1mT1rYLEdobVpQIseFMMaLj
DDaEJLZTgEG/2iZvBJXTwswDc14enaaqgpwUfZsf4S7W1XiUsn1GOOQl4NdnXLcX
7VnFTsk9D/XuRIyQ69YXm9ecuJVdAeeLA2Azpo1Vho91t9gahMCem8tU3gc8d/f3
o/kP4bT/lRS1DjHeG3tDFA==
`protect END_PROTECTED
