`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G1f1g8xTrENviEQ5W+77Miu4IUfDL+nfePkQ+5IEYA9gAdx6fVkgg+7v3lGrb/SG
vGHxjp0DMqQcE2bRTWOPplRvfIgFfnrnmlpHcpXWthiP0G3DrG319KmYuF+F9e+r
tqElqA5HGeqo3v/Px+giWd/OUEtuQjEG2QdBotRWlJbs9y5w85ST6irVPXS6hOIz
cGxUXhCs3otlTtbmSb04hfVHcpuBFUmwQVq1nEo804TFTdLsUyV7pMVOw2hVw0+G
6S3ecoJbgLsHj+x/vjp8e4MqqiIHUM5DozePZ3uWG6RM8+P0gv+I2I7xjrBhLsYo
Kwyl89u3tfndmHL29B6eqJxljTyrPeh+ss2W1GGPva1mKxsTA6t/jy8oS3aaWbF/
Jv3CrO4Lwz0CkDkYkWRR7ypw9wM4x08YooWvSMuS2rrpmVibvTjOo9jqCVqcyDki
CpT4GVeyi3LtUzoHFfBc7YYmtyfv0ArR8KuYieZd3s0asKomkmtZbCZDPGk7BXvi
8d8I1ktc8A20ebZad9b9pi2lb7opzTgHJfFtAJ7mKeTHEAGZ5viIBW52jti0GxeN
93+pyk9Tw8RaU5otZhuu8NVyj/TKeNKHyN1hDhckTyoGRMWgr7BaAPpIjlXOO2De
wa4R6He+6Bk8YHy4wXj/+926JpmZS4Y06Jpxbv6Mvn4=
`protect END_PROTECTED
