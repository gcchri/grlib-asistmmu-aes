`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LhwY9lqIdnRsZ5iqf4dC/71AXBxKXgKqmVixtRfzJKAnfIYOI9kK1cb5zzqbjgGm
/yAyeRhrosLHPS+oBzLxab608rPS9bwOH45nhWIuevURDTlseGv/XSd7zEHJwF3a
Dev45eZcOGm9p85DH+qwjls6txkgRT5Gpnsnz5ttdZrJg0eOtb8CpasWHw58vdbL
fYBdGIs4UXw9UVCI61JCZw4pXTxKgqcQ6Xgwpt+quVE6Oh/wKmSR5BsruaeKOVHn
jfJa4wS9q/mahUyWVgkJiMPq2lTifxGfaLkF0PTrtV8Pji01GBpnkfU0r9DPpr0J
+WkqculDdy5cygk8ui1Gmo371UniuL2S+vhSbICJnVflV4VdW9lMW+K6d4LCaENP
sJVsWFyCVQdQTpiam+t88g==
`protect END_PROTECTED
