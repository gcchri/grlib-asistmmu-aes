`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olHZsDt5GOESjMgcOcmkAjsKGtrY8n6uW4Odad5M4z3DkdYTwpPgjzNFpyPVLrt1
fNH/0QZrkOLNvrzNFbzTL6O+wSflR3b3ZdNikiUE30XFFrjI25vesvDX9GgbJbQQ
fPsFU+cR9VHYgpEhqV6LrvEdqNidUMrahOxbmVyujDPBe6pmOTuzqzMWZPTIo9/Y
J6DuF/FR4PX+bTGz3kb3HvMgR9jnlm7EdZsP96DbUcAjYUCgsAGAQcD2qTWoE9xd
ZopqyTRI2fkujWky6dqmiAjWZVzzdPWo9FZi5pvUzQouDzxfQxOqqk9ZVoT8eKuo
JRkcA923GYXbK+IgOs07MFpD+GoRJbeDzhSpzOx538uLRptMF+rJJXju9WnNf9Bm
iZDputRtOiPHyrJJZqBW8D1i4NMcRVRXx9st26NhxSreXA66Gd5Q5OL4duutFQJu
893iz6nSWnzTChNzNfi2/Tel7tbUDdOOmrih9cDIIAh+mQ3LrTJC0dM7ECWvPPco
ngAZz5TMa2jwxPUhXfOK4YLHkYxdB/Q7RhnwHM5agwcGbgqZMRhGtVRSY7CiDtaA
7bYdsPwiZDREm7TCOWXZLf+sDWyugWVLRrtYphDDtPuLJfm2YEsvb53rgbokzRtd
qNaP3VSbLA0MN9eUMIPuFLD4pmBIV40K8NNNPuBGgeAbjIWadmsM98A0nK/jlNFi
LW4BFNzvCATrZLwlLfL2p0Q2KfuUg2Bg/6YImWvtjms6d710sbKL9pk/G0xM2GTh
8CeuNedOFnrgpmQ7LAOsY2hbHC0tyk4owdOpLdyxqlGl7cs/CTgWYsLmZxoRCZyS
8zz9yLyJmQKVaBmTC3n90usCVgaEX+N3YppCfqsiiXU2MtWDpf7mexVSXEuFSGB2
ZlCZTX2dG00ZDX7RJvpOKHdJwMAc969CmIoLE+Dc5JWheFsWOyJ8E6J2recRh1/W
H1RJbSLvCMhBV0tYOiNOFqhHM8WPXAOCc6zfXB2h60zLZxAbMgYNvlSiwt9Cv2v+
4qx7TxJTzCpM8AkptAT/eL9igP5L2QleOWbYKJvZI/6JkEvPVLX87ZzVFMJGbFcQ
jsh2vxaqp5mE5BeeVkYzVLjrX/XfToOZUzCDN/8a3c8BqRookNlG7KBNRiuVbwMG
VCvWT0175UEIvPgoav8H7aPpntljJO3l+Gji5N0StsP75JN7l34iSzAW3ZKi/JfA
d0u32yK1Ex0zM0wcjl2MMWlqZXo8fdmwn1a3Kw1H3ZFcZy3RHzPnENUYjE0byZ+S
Rwf0BrCiC9kcQSkzFCOyrRDFIxvwIHx5R/34kQMeZYfm3jrNDOGUIS2Ue146P8XX
xIHFLiti4gBOehoZgHeumwi+oW25EaSSppLmJOPE7Ld4ZjiH2PHBEhC1lN5bn6r0
62XrZMObYJlXZ2mhSKSaFI1wIK+DrcadRi5MnHG7PAzVPupOmez6lWVd74WxDi1g
lfj1XjRf7+Kpu9IrCULzVR7qKYO8ekpUKNrpAIRIfDISSnc62h9XC5sUL7Q9rpkO
spSKyxMFEr0rAEWRmKO8y/9z1hukePHgfIs6ZOPYcOkhGZI4TGoOioX21MmPQQsW
RaX6P48vZVgSX+SPGPzgwYi1/NXfZsAPRSwy39ERm4d+ycYBmX/6AwKs959bWLae
FyVqpBttNRmrJCVtZjw8wV/0anoVg5tsRSnfsMY/qyAK2IMitOGpa67wy6Cz8Gj4
ZzrBmQbbIo163+Fn2KKIUcCF0kgCDUT83EBl/e7sz9LkkP7Mqv8QEMU5a1KnBhao
lTy6OZVPGyf+Vl8/hsn5P5j4XS/ap1dgF5RAgxIGIPD33hje3X3jcxlpMyzGzSbN
xh/HAYG7H6ntE24ZTXx5f/ZRE5aeznibj1RmtFqBLa7vLdu0FFFD9863iMp8hr/7
r1zlCl+eoCeIVmTd3i1xGI1mvDd+GhYm62Eh7qrkrzN6v+o/1S9Rzlij2FTTqjpd
vnyI7a7OLksNs+uvgJRt3KKQKYXw7RYK4b12drr20ime31W1CMBpQf1Ao64JXlLk
P7bALimBCsAh9AfDt8wnA5bCuNMgv+M787JpE1XfaSgt0j1CPZU6dJydiwUtXYpF
UiqJnRxdBVAsFDGac+72MER4rZ5iLG1FozyHpKiQuH4oKkc4cBsoeEFWGPd7a/Cj
pU2l14XWMeFs/PkNclLjQ77R+PlumEaIMTCviDoPuQFwjoIG/g2lHxLtxihnlA0V
LcCLDhDNW+C9WZGfSMsGhYyDaltQvEhRHEgP32NkrKeFIAqSkgnpFty/kjobqd+e
/Qqcf4LGgxhos7hcbzJpdmvN3P1P3M+3j6MfHPQYiTNjphxQ7H4pcSJgoObtbJa1
5v70T7m7e72ixUFOPNJa+50jooRaO63QzPQ99NoOIroHg7S96IQBTiyL1372TfEQ
nkpC1udx3y4N7WmNbReCKHDnAbZ1bEOsO7OD1CgQOoI0l+8ejmje6Kkr0hfuSlJj
v6YElpNN4Iwod1bEfaAQJQcn8IDKVJiQK0HsRlj+IF7Fe7t/w2X2TSvVpe6fwaUN
sVWLdVAYD1uxH0OnWCJ190+ypwnNJRCXmu0jXLauZDaUR1y6ze3wb3aK0RkwfILM
wfDW9WXOrCeEUPJJ97xvxSzr/6kUl8q/UC97uItZRth5q0GKGGa7Yr1voq8DnSpB
IMbwdhei+AUKrzIvapkZwnYFe67mrRmPUycxqGJzx8zQobqkXcjZdfBe8LYl8wye
/M/o0fwe9dxLpIiYwNHpVA6DChEX5UifJ2HLVCzlQVvG/9WeStJ1mD/jjme8JHQw
FpJbYLZ1iyIUe3MbEJiNio0UBLvEgGBxoeGrrWTAdSHaQayEc55+dWNsT49RyW1R
RSW1e2GVULqUhtRLNdZuJU7ifSV9L9CUWkLP3LG966CjJWhyIe8F3cm4yWtO+V85
JVRwk4kASy5zTM3B8VBoUQNSpOAN5j5wk5vWbWJqzRoMP7uRIwDJYp4BQ4mfWWbj
J6eNrrZyNnnV3rkJXsJqgfiPeJmCeHCmcvZLW9ES0X3x5eqYZNTzlwmm8LjuIhHQ
ciyMc1MU0AsRwFqyx4uJG0pMjt0tcIevbZ3/kBH/JQQyP2VvZtyyMN5ZDfwlc5uZ
WHWalj90BD16BUbOO1CLC/gFOslCy2I+hGoKmtPfkdbBg8vU2+nh34M/ap55wegp
vGEEB04eJLEhcsK7SYiMDamhv3OMo1G+K7f+jPofCxiyxhNaCb69fU4U3u4VSnlO
OKME4urKDWdr9sAJuhogiVYne6TeehWMAcuL+iOPRJFYtlJF9ZBNuQs6onXZ8MuX
QVAKey/WTm7maxTOkLHmMyoKJFdm3otFQGccGfAIHB71eLA4M/IuvcikXnQLL083
UsvWmbcD21FwGUvxJpDeGGGdBJqqwaMUcxWriNEuDOgfIFHER6S1fXdfxq1f2SOH
YtWjPKNwZdiGjTv6WNfB9ojDjpc+ouGUUwVfcq3/K6h3fK0Mx0juW0IVBM6jn/ZO
KlLZrvs7YAyADTDbYiQv7kKtXdhcZ5U6kBDUUOB0nH5Cbjs1BaioM3d+tQxVeoZ8
y66zv327ybE6LLs0Z3UX+N6KIa9E/DfwKKAcrzjmINRbM+OKmNn0wgmhSyJUk6r3
BLrGgRuBC9W+YnT5voSQ+gq320jKOBrEQ8/bbFOgoVSy8ByZxfJNWgky9DKw0iet
TNKClU3muB6C86Ww7Wl/AdXpHMxe4tRLbtLZ9rLHmittlotZw65RkY8krtSJ0lhI
40QBTIHTogAtRitG5YICkizezyyFOWaEfZ/KhinUlzgcY1Bi5ahKBYw/5tyJKN1a
JyT35BwI8lbV8depA4h88/3KV1hzRY9CWvF/nKFLtQaPFO33lVKvfS7cP/GDKh6h
qodpRL32/hM44Ow4f/wVgM6upgxfwi+vV8ggX39+1w1AMd/w4hv+fz9K2MltgXQ4
w4bYzt+CEfeicYOv2CI/XyN+fGX5iH2qmau5oFo3NGHSUf0GR3o+k9RtgVdDi+1k
NYeu73FH2cQSB0JLpcY15JG75q4hGUWI5kb9Dcue40PlYPaZRMpy8lIxqOXsPGCj
HSz6qGc7BubbfTw34t08LvL93hbifLCHd0p03jEPVN5ICCdBjqktX4BznJRH0W3x
4+JHpRQeDf2lEXkLd57IQEjrLwZBBsDEJxA56pcE8vLqjEpxMaEDNPlJHiJtSXqu
yRqoV392+Yq1rfmI34SpzElBawJcinlT/7MfqyPuI+gcp0U94ArHy8gkj5WkeinV
4mtN6KGFXSwXzzXQ4Wryg0/aGIIeJBXP2yXOdAOTwoeRmFmvl8PMUcPY1V2SWtHT
JttIehQbyxnQbQgwJEaZFXwPx+93O/0LFNs7Yz6vLt4L09Irjd+9Qb9kE5oKN5ZA
6/2X6PzA2XZNtyEPtHtFEY6PHWfeHbndLDlP/vGYplVtQ7LbqXjNWkFEowUM7mQJ
sLTK9ao6+vVdjcNXUDc2CJz5TFp44liFqSvEEARyyfeEtajlofjsD4nezxNctg2v
4sX1L0OUU6rDEj5KSz3ELXUVYrzyGCuE7sQIYHRue8FA+b9n9num/o03Ns+YaAg1
4YsS5U7Z6UXMzPJzjn6gSiLAwWU0znPejVwERp7AX3LXSpIwCY29Kg0N8rw0lEBf
hhO6aISS0qUeRH1tqfzTyG3ew9dbIsZ328ypYXH4wzbM4sgZhiY52Ut7NN81hqm2
r5D7GR0b2yFpS0pBVp9bFz3PbaqwbT2RLo5LAKMzpX+1LgxOXYuJt/6w1kWogGSN
xG6DSo0b5Ho4jezw7tQg4sbTHDuHlmcEXZTPL48QjagfnjuMoE4PSi7CNREgZn3r
J0Dxqv2SYfv23Wds0XMXgi/MOW9BPM0TGOK5l4nA9ND/5qTZ8SgxmboF4n31sDG9
+eBJhD6ENTtKOC6cgK/6rjWGo3tN6Mlvcf/M0gyunQBdsMw1gF7oBG5LB5+5SmHB
xxhK0BZ8+22IlM2TrIzpxAj7rFFShL+hOsWlW3zMdU4Y7zbiBV5Ld8IGcguilC4B
gu/OGjPQ9isCo4+KBgxvlvCEKQAOzaU25ytDGstAI4D6KOKkY2OrIYpCeoFfB54j
bXTKXsGCD7BidMGLA4S6NypF2BlJwoYntnjfL15v0hvNn5dr+q6+238iK0YrAB2D
vv38J/vPByVI2zpCgGqY+0DnkOIKIFNf5xZ5oJQ4QFplDJ1l3c9cUZwPcy596Fd9
3xg7CdjKkcykcLFbF3Hudk96fv9l4sQ2RiMjR1nV/7JbEt7MTbVF+ZLi/wtw/VBQ
KazZpFoXUjPdqMMj3nsS5EXwsuMcYn1mBlXCkp1a2J5dEDAOeHE0IXQTW7Jjqjk1
z/OO7ji3kmYTilXh7OF0Mgtv7cT++1LEgMuKSmVNG1pcWQURg1lyDbo7MHbrPbZ3
k7QZBysmPBaSPiLGUbqgpIYNeOvB6Ie1cu/OWozFMPjzPyZpHBvim5G+RsQf1tfv
GyOWtZKTEOFiJHLieXYFxzteEzQboTDyKUIZcnxeH7l3CbAQ1LYKZPoDQLe2WNh1
Jxqxj92ahKjaj23fIqb+SMzNz5VNmQPmolX3grf+6qWUiahnIlufcsvbv+f9vM3l
evAZGkdTUIeJy7g4tfBQFr/MdmtiYoxeziuyEQsLWrRG9TWJlOBmoiaF2ZnLxOtO
Dtfze17YiKKeur3jhIypTj/G3MqM0OgpHzqTXYR+f3m619jLwdqGVm6GbW6ayfPK
0UM/YlWEDQc1tpTOCp/QqBP5B0yAxW5vhzqtFr5EXj+L1SqeFemlZtRPeB6vijM2
ExwHbw4GsNcAlIMgDmE11ho6Fdm9DTB3mhdQYOKWT+nmDIkMeywNhdo6JdOCShZM
HnvAzonSbcWb3ZP9hHbEbomH/3jsORzXbsVEz3Bciufw7intk0MRpDqT8CCHNZaS
IAmBGbgqWGeOV4xOxrt+BR6y7DTPALd3zcv9l5r3FgQty80QpUpC1xHyIZx2y43J
XYuxUDH/2lZ/wRCPqnkc4gDP/T7UHMtsBU7OknZGP81ctbD8gPw2h8jpiCuxrBMT
IlkhdLRIFWfDYut1oaS8VpTvYqq9gEwnDCTxFn5BOkMks7YKIIMORATaXzdtqkQ4
srcX+/qJfVDpPGA5ahJcOwRouy7vMZA0HQ+wls6DXazw1cE+3GbD6Ze9DpILRlRy
wfGk57zIoNx++JAh8QXvOeKgR5uKBpA2XxTkBB1GN7gI3eSUnBiVeNnv/x4Eun8v
f3swDziW9nouKYb8gM11vM6CErjOsUtSjYa/phpnpA10imObzXqHBq2OgWRE7859
RbXCAUJi7TWuskZa6lMN91Q6dhkyjQfEVG2c3XN6QV4MIaEHvLoqrgYWm1IHIO3O
7RS+dbJoHAYHcqOPGzH5G92i76azN5M2IWA5fAX++pNA6PIqihzRZUbMaP/Qjq9X
yqOl8A++cnU7tAtQbJEjITnjyXwhkauaLqs5rFOBqFQLc3Nj431/quhDMHbOodWy
ehUGf9+Ry5X826wcjsj4V8W2Lb5jsXPzh4J+9hKa4OTukslQm9QmirRzrG6DFvTG
SmRJzPdpPYv3yLJo6EWK2fAEecMr+15gs44AM84HXMbqLTSeVSvEu2tFknFq/Tai
R8oCu1tuGERPnBvo4lBfnKgj3dnrTmJSrZdbOmEgoEvGuZEBdtlloaUuulVob/ZN
2Osr3B+iBfZc+IlI9KEtd70bMb+QGVakbnoel1fnLm/Xi6DZPoUoOPbiwPUHVnRy
0TvHWlg7TapAFQWm5+zkPwzwXs3ptAXkpyjSRdwPo4Ej7CpO+GFHx/f7tB64FrDc
SaIwOuGoY+/XFJw26HD7tCj70aAaU0ZpMeRDRpbAPD9amYnW6T1A+MLeTfEF5InB
EuNl0yrc7V/zlJpx1cc2FWEd9rdI4gWCmU+knzZyidyl0sO/y3f/OBvnVTi4R8EU
cXIMu6obj01NSTgFtFOd4FvX+FJVlO4sQmsvzvc3vtFB3EOfzS/nCDADBAKcp5zH
IaueHXUH0L6ObiBV8eOLEExyMrmBG7/ML/PfTnEfsIAro3OSdxVz6T0kOCKn4B8O
jitm6dX/o/P1Nqs4ble7e0MMC3/PTzPyq4OP0x9a0E8pYK0j0SHhTVwjf+ZW5mJL
p9Ca8SQ/0jISGd2Pe6McfQOz+jfeiSZK71OKuTmtlPgXgZ8qUD1+uSVJUtqqffr+
dHjtYYs8BqbrnUflprPnZcwGcJY+f3Eew0Eijtfp4D3KgY17xXozoWJDr/7t4hKk
QTsAs+FX8C1NejPhWI6QNT2ImLyQK4DhV72151LzlZB84Iad0MHPhCDkzG8N98Rq
FtRLFrz3TbwqWvYfXk+kmF9x0+hE8we4+mQk4qOsOr4FOqMpkpsawMmfE4tYKoJd
6UBVspgUvWyVeWBookbe3nrWtOiDuDNVxlLDL4Tkp7uBPXahzaFq+zFA6d3r+POw
VIdkTwxr0RxESk1ialIa0QVKJBQ9MMT96bCfnmQ8Z6+TYs+NNwmL4iW66caqSQ5b
GY6yptzzIZEB+ygTnR2NGJhgewlGnUJ20ibb3xsvLSwfgPcTGVeMwxLH+dk3PcKs
de+6t5aUw0c1zzRBqKrsKMk1oGdYARfQeB7NYoqlIqJS3jkaZYuWiYbHLIUadEUB
MKmDAafQexrp23JBXFwsFBMzk2ckmOwrAt2SN1v8F9UzbXucqkvGChlW/Q2gAijo
Gx+NxglTpghnE3JJSTUl7RMBLXEX8PdJ34pjOgRtSq6bCabJnIWT57X5yllrLZbK
Pgq81IjkQEI7vj2jY+r497WrMm8Ur/kzqO3VL6cwtWtWzqDD6HnxR3VGySR44wVG
jE0mdHaGw9aLHCfzQ3x247bevTnkcUkp5boGci3Tayzqo3mkG19iVFfWbajdIy5M
sIn9YTXBlmBGvOQQeQrzc6jrMK6sb6f6r8lnN7/ja2pDxzw7OLa4Ni6nyJNbsBQ/
isfEyCAaCl6GE0sJCeOXhKMCE65vwaO9Ly3QreKoa0GaFPLR0h6IO4HciWZBDtid
FhxGdZFP7WTEC7xVM8uERGbnw/HyBiiHecD0jpmzPzHcYzfVS12y7myYMAZsqMOU
wpnqZrp37T63N3MVjQU4B1346b1DTw0xkxVXH4RZt8Q/IuB6GoUehtRHckuGL/ik
YJ5XuPhbMc+868qsI/I78ADOprHFqWOrrAuejbhkG2k1QLHAulFJjMC+IxNN3Kcu
Bg+wMYfC+lhQ/eYBLcuSLicbd3MWjIkGPFQI1fCKQhs1GSp3g37nVUMzHAHx8FG3
4rXjEgkZ13+nSp5PVJ0eVlwc+pbqkgmkgk3uYgwl3adTYi20wC0nK7fu6rp8oWJM
e7GWuUUFhfXCHs6KoUKnDta369zscmvm1dO25sBqpq2XknXdXqWQ2yiI+qWrmZ7z
SpPJALnidG2mK8oSqUQD2CVdV7ZEKg4DtVtaP1T6gk6pZ5BzBP46Gv2JYOSaL36W
MVgxuhY/tEk4v1M6R4aiqNiqbkpy6erap2futkRC9bb028WifXZBfM64+nwzPM0J
vWUnaHj9IfTm6mzWz0ji+NvDJHE+zrWdD8XnGOYcLVlf79GPbj/ggCWK94pVsKf/
tJBwsucdy9QfnnBXCgcd7E6y1/CBWw1QKDT4agozxrWQxrIRL7zVPSSC1tlF4Quc
FBOmGiwZFVO4iZydxCYif/L0dWbh4syUz5OBfzCcdC/3mV2hEMlYQy7A7iyYKjk+
B8RdnJZ17l4OP42lBu6EkULPJztQ8WaGZ1jXJEPEwzWeWldnVqg0xmA2itrFt/Fn
x4cGkvJ0pa83/OpFH3zaQoMD7QPzlEw1s7SeODd0HwL/q7yi3C8stJ+puhIkiMjM
gOErd1+HYl9rR4Cqki3YKgAXj6N80J9MRza7jQ8L4aOLTp9QPSF5v6Bcd2f4m+8d
8lQsYGyq7ls1P1cu8TbndO9nnLJUpoRN4qUIyozv2/nM80NlxX3Od0EjjJ3Lj+AS
H4sR98EU8P5gfTalgq4CPyM6HdPr1UWz7mP/uG1VY+LsMQDJziCv9dhir9RvJiZ3
cYRvRWER010jY7q6BXCYiDrxgFFy5q7SK1AiCt5XuYS/X2v6j5/srxAzQ/ZOjjNj
O/WLk0V5JPHQ3BOu1yg0KKT8yyO6UHE+E537fE/bhgB6Cinn6rVionT8XD6aUsQK
GmEPA6EPAu/Qgipfac3+p+Q0DDrhXsFKBFi5ZkEsgoVyeu5ijmnOP1PalUFIR6Jg
CRfDzyb5LUdNijIYJYFr9FGHBacRuE1T296qPFqg100Nkd+iMMez+1HHdebVb/Xp
slE28QnGZ67fwC36S+SXffPUxuDpQd4wySwmmuOlzIdRB1bulqzX8nMDhPPn4fqm
h+FexmODlUbNYxXeaXNKzrmjIiyuHinbKmzfwROXvzn48EOkC0T78aYw+DNLHUVF
NVsxKWQmH+ugK8tjG2kYtmtx5elXuwqus/WSw3xFq1G26f7Ut0FmIqFUTYPkMnxI
EtF4hDDvGpaYqEfK7yTiU7gff2Hsmig0aAdX5ydhkgP9rhWKWbp9EoBuiGAt+ulO
3njF67caUCThy8JxzJiGGGYahp4EoknawgY5rkKOKwxukooX+GIe49hwjQ49l4hT
OTeIyGqvHhvVsUEDauRZg6gi8r78yJHr6rrP24h+GZRVbeVaNkaK05A5oBej3OJS
p1fkx5T0ZTKauwZpSIx3B0Ps/SMFHRKcsn5H/585qhJxdQGlnBF4Kq9npv4syG/A
H/zYB5Ah3CAFAh0fqvSLLmtx8wESZYzEhJCB0WNWdzjA+bkyV36T7NFVhZOFkLqj
ucQ82KrD6OmKePScdAL3Og3pVWrm+NS0mB88QicHXmL4NJzSdg6YFWIdS+uVlSRa
Jo/4bN8vvPSEpqbOdiejukjs7TQa6nI/5q4EEb8foNOGnemtNlPfwq4rjkWnl4dV
fyiEfw6VpFOHc68suVpubzn6bl1ACR2Wreze+w3qxR17bDSd2yuflasZnHuQHKGw
l0LU2RpMX8cExXPzbmUrG4HQafKnHRFt7rEGZ++P1pan4HQylmSS5qIPI/1bIJyp
ZwLq3b32GHeJ9UNh0+RKWzNPDOnHKKZ496e/AKU4zSggEo2m5NKoN+mekXLGCGTN
7E3QTtkToRQZkcXsBE30bQiODrSJIuBfRugVifbMLHqqkopJQaT5IKrDgoEcIzES
sr9gH+P2crEh5xjKPwYgrAUC+kUefYtku6TIFxFtQ8QemaJb0GK+Jnf+y1HwGxgA
nxF+jPxEdNcEERw0VUVM+w0KHdWikwT/btg41B1cGxeUOcZveBSNrNHMEqspO1VA
ZfGogteUMaTmmUyTCwCdqXjQYOOdo4EZJMJ8Iq9iZ9tGLs2Qh0RdV0cV9d83DBnQ
BZTnU8vtlTRvpGP5WXNxiz4q+B10NUIKMkGM2oVWN/bluYenVFYAD9P41RPcGSgY
lPQXVJ05y4h9LAitGyytg/NGpp283jlEi1exSVoySReq40hx/fzW5T2+eMChGpt5
B7Vp9GlSAHIXChTt4XL89Pvp39sRe081vIJIFxwZ+6+AoGi9/ssBDB//Rj00JtEn
74F03OyPID0wR/4KWx14whoFzC5axNB+1zudKVOq7kd8U0idjEMtY9lzjEG5HjfN
X8PmYz6S0hIJbxIPLMAp7l/MW4Ax9R2Y6NLx5luJHw13AFT6UwSUOU3K3hWodbUu
RbpaU07MsIQ1fyfdFyclzGatrplCSqFoSI3csKPOR0I6OhhPvHAe6AAtUfUUx2cs
xRonSduk0Ze1Nq69N5B6rD4aQOz8NE0ZQuHPKz8GLzv0gPiuAdsluUqpqyJ0EbZY
BcxJYj1LNzcZSZquvw0yLDNKuhNLFgWHdo3vDpulRbmmYpw9YMWzdQGTViiBV0mu
k/YnC3t1KylsZl8UvXfQxNzztPf4PLqNTzdnuNn/+l3AxJI+SxCacrZi8pLC3Mg5
R55rANjCI2fc49QOV7PqI5MXmnptUuXLVZtLB2NBQSEkd02tfCCKSDiyLMpw+CDO
CeusLP8K4Lcqv1lZE5/YS6ZMm+eIU9KP5CT/c3GE1goAEZQmeo1RYBh06uMgXD3v
fDGSvE/LuYMTpGLkhj07KuhhFDe3cjoG3rRIPhLEfMisQq2F19Df3wyrmbRxdFV0
90tZ7g/dFO+1nn5YDOx+5R2EeBO6fHq+IpYlwuHs9OZE1BWp8+EoXw1fQWMCfq+Z
r2MuKP1Kg3FPTubMzVB85pbmSVVNfQxeX8DyUvjf13op/6qjAZ/Gtl7hRoPN1hEH
faBgsb0sFJP8Ey3Mok6iJ2RJRHWkEQIyrwd519Pg8cDtFT59acVidsaVIsW9SEDV
dbZKTPooCMWBmsUkAweokOtrx+dB710YtoiONM/17SVkE+FkoLVHWu/rTZPEkorO
Pwdc/HlyFsjZLFbBBd8sUyr2c/gGpGpHvIXMRBwL1SVZoS1IBO8s0NV+xksQVEw8
NOGDkGtqF8Vnk6U1YqDrIsqZTE2L9hWdgqGPtNqk/h+wo+cE2D00iCYoUxoc+8im
G0xAYMm0ZLUAjbIZtSLafEac/DLARMdeoEDmJCp9t4xMLffPPyz7ihrbTFIl/tf0
WECx6vMs3fUjBgKZANDhor7ZDzER7jb5CKYC/a7QcpkWMk25b3dpMKDqqDPHPn6R
e+2DYVvd20WiRaTIjbdnCe1EyheJ9zBYVHJZ/NnQuUm8bg1t69vzKjfNFQHmg9oK
AN4w0n+m7V+Xfiv7WKBX4ZD4RxIvPVs85f2Ut1EFVbpDC4jWIPKwp7h9GBRa7rKG
rlEGjQ3JQoPHnqThr/b4hy6WNvDifAFfsIxsbG2Xb0FnYT9unY1bFYuUhZ5gO69Z
AXisY3b3n0bqD5GtngxUOj131iBhB/lOZGN0AMszdJq2xptbrihLYK5Ciz63Buio
+NutaC3JdM+9LnBTvlkQrSWhfjnUb+h5M3+LDYXvXsGm0X0z7hdufCduhl3GhodJ
QTxoVFkHCOBR8nrPFqhb3KzN8R+PB/uxMlJTlZaHh4ORpHDQ6jv8zvq92BtWg9H9
/lvmTfUydOwTKlwvckEtKzX0+UHg2+LzQB9j0ZNLLBVHfdElJMHKta/wYQhJlV09
qYhaw4y+YjdXV+KbjuvZhPR+AgC8L6Yd7c36EkLyaXf65Im7baYUTaCtElhQSV1T
1+kCGAiDTNuBrdlhhdBjkGOt035SeoNb6fQwdy2p8leYOqoebfTilZfgNAJcE3sa
AeT8q+HmW04TEdw8X2mTlkQPI4CsHVPoZfoRsnvIrNEZdbvuUNNoS24UYbkN6h5r
JstS99n1h2ITvDBUlmHpJ8sBeZl5TzM3rCqaQ2rjAXz4X0tgbqyQgiHVj9EQWnmw
ekOirLUjNyjIRdeTX/aBEPpfPSJUlkW7UUe2W9f4Np49ay//tu0EoHO2QP5yXt2H
NDz7ynf2Gw8xscyymR+JzqrSh9JqDAptr8XIVp6q/7T3CeX3jeeIGts34shDRXQZ
piJ2gwVpZMN71xmDqZNEbUO9n9MOOTRRAwbJfA1BdemLxFVGfJEBklbu9zR6OuS3
s2+/IFSCZW9zS77oXbEoC9s/tZPEP5JIp+F8+92vjuI39SyDiRC9ylZU7rkVMr3i
wOSf7KsMsTu4F1EdmsDRmBJWvf+0HzBlbbh3yVErELiXF20TXYjN5BY7FYjhdGOf
3u1MGExF5jVB64udj3fFhIzf5OzcvjoTtprkQHkj0yr1DVQ5r7b1kClfAFNcvZbZ
H2msT5QrdDu/ck687w3zaUVZtc5p+javKdmQke8GfMLR2mDJ0nIpYuYZVuFn2vcG
nKvkknepOV+5PRarMkDBzcwrI1t9aqk+anGSh28vNT8/aBJ69e02noPfkwiWhNAw
iyysXCHY6lP1A2i75wONiLZoyHqrvspgvaAofXtM5QW0sRuKmaXtzWa5N8smxdBQ
5Mg60KU8XPFpJ8iPxWJH3WrXnlF0JbXcSYq1xQihOyjlUfHAeU7eka1Stt+AeOh7
tIDSb3WB02sfgWt+zA2WPTbJWaOD2RKd1hOBmrAQoegV9Q5iAI2v75fehgjtsb8b
ofNLVhhyO/hNvitW8hRy23T6mrO4AEtXuBm+N7SED6A9LzkfEkRX7ZKhJ1dz+P9y
EhXvJQFWbU1YPjLR8trGKhgXbuZmUdmeIPoxnxJQxgCiX2pV3+1Nj4TQFvFrmF7q
qffvcc56pAcmbKuPWwTCET3TaD/vili78e/v68+QP8vPVOFkEjGm1jGk4KF6MfMl
cW6fjQ+eLszskt1iTowMkk6Hi9VIRE4F5diOXufaZwMEMU9EhFouv9OGTPb0Zpbj
sQVisRaFjGMDOlDM12fWQU889CPQ+KL6zb82SA96aFzaSYaFyNwSv+dhB6Ma9fgR
/v7ZW12VYqYoIaypitmyTrkF3WPCT3frH4CC2X9fB72hJzcBLb+PzGWOE/wbOYOn
QuubJInbtpmin7IDmmRsK7YGoomF3j5Sm2I7qO3j0vrhrgsqnTCHFS6HXBvDh+zP
JO7VUgzHhHLepqVND6iKgPD0r2B+L8S7jKLYtEjN9F6CfgzVK5eryeOnhAXJ///N
sYjrtdKWASyvplHyVNGdcvG0rfmWQ/lbwDk3AhcO1xL9weKnW/43w5BUeLAACFs6
pxLvnR6pCX4ovRUE1fxejlaB74eHIQgQjPmGhXxHfy8tfc6LJnqhKJBSGr2Y5KoO
5bI7kMZJ3rz2uqiJ36BvfG1K8f4HKo+9uF0oB1h4McIzkPiDFL1ZgjF5ic6jQSY9
no8q4L2PNOTBuqZW80ahNwuCVTJvkNZxA+cScuFYHJyG9gZniVgGOWbyaMGoGlh1
m2UWx+1/QpTXIJXGbXtod3g5zohOPAW6qUbl2OEAu42OsOGRyLk1Vp6aXYonqR3T
nKNAYlRXK5OhtKLLtclPxTqlajBYoSyRfGpwnOvS3tpttw5g+A5uJuLwghUWq6J6
HsKE4lalb254O75gu/7J+geJsp0QbZC0LIbOjGL1pLfnFBSFrqiAnJS7stQey4co
Y63fIyJN/uGkmfaePefDJvliLlTUa4mT7sephS63rDBrFPO6oKyHoRGPdJRQa6pm
cdccTY3yCbupSTBV7/vgQIYbG2v7lpJN9UKFdUEk5CuUUkGSshsf3x2j3Vu0v+7y
JCQW9UBEEtOzqNGKloe1mtMIp/oyonaF+ODpkaTB4b0uJIXQprtVZ92PpR7eKe2G
KKrFpC9US58OlpN4jcGW4HjXmvgPEYIcglyhgBL3QEvH2uB8seNFmE4wHrOkfWlJ
tI3coCD9b1wdb5Y6rAicnIb/kq/9p6IgeahlDILcEvAzwmKCIFLMRO/o2u0Na1jq
SF/aaNAC9rS5JspFxxYznOCj7HnCBvcgnG2siVI4xtzB0tz93U6QU45slzK6ftGY
txmJETFJHUtG18xgGPhAdkZQ8jy0rRPt/5y3qdosppFQquzWXagtlSCCDdnJjOg3
G8CyDPGStU4D/YBm/Bbgf7K/CaQHlSVLvZRLzGGF2Nx/kULJWsKS0L/NwW4aX5P5
s8TT41gh19Wj4qdSX29leTs7bcqWuwp14xcHfn6BxOczAlaGcZBNgNIvcox4zKoG
mL/d78YCwqKDwAASkw/VrUm2woPu5BinKFF/s+XFPaUaj1WkDyFdb3X7GHdGppR7
vvKce1QWo7p764jslXgGLl2rLzlSMD3TE/jAZP3gP67jIrxDaKvWI8z/2GmnAriE
+Lfwy8+CmFBikFV6F/6MUB/ENKYBQPi/e/YsNfBrcNtsODYKl5DabX62pBiDr2us
A+YAzcTlypWHOuQiO6M6Ka6aHpsfC1AzZskshpLW//cPsS6tjNrL4E/VGo3rKN5D
AoFfFsRXcr2EwIASco4S0ySjawnx60uHpLr5xBtmoG0dnulzwIpZYoAsQvnQOPma
cw3JMgeIV/WeKEbrUEYyg+ERMyK8ymOYEEJHpICmpCivRjV6cIuuj7ONGT2N4yNe
5dZJ+0TgdLxqtrDbUPd+vfhVSk6s9/DPfIx892O6hsOQncYe+qaBGyekIQFxpZJl
gdRFiYP2mN3rSYaLV05ZtSNqaTib7BcKbEbv3WONNAIpid73SyPKPCG+zN33+vID
j3bl8G+001s6i/gHsyZGOXnx5dHdkg1fRRFu2RIeRheYTVR9fEKNpIPOd2UiTxZs
62+ohsk97f7n7W0DyoWpBtassDHSNaIvQSxoqK6sWvXpJXEZSQFTqKFlxF6NzEGt
rqsYzmVEw1dwaQrs8XhD6oHDMpySpR78GA8ldfewDidMp0NsvuBfPBahZ6c+DD+Z
Z/cy9EWAIIB8BA5oCFle5k9n+dxM76feA9mmW9Vrza2ebpnVejJBNKzqnQQogmkg
h9iG9Phu8wGj6Ic6Fbx8Jz/FSmWtzIvrWCOXIIGrBWkKJs2JXJXnckmwZHbts/ve
DlsmBlVdMikBTxvb6beYW/WdN3myaS7Ro0hBESZ1mJadoUU3UFpQ/O+JSAmlNb45
uB+uw1pzZXN+NeUJig5RbIwgKk30LjZcqrBRTR3V249CEu3H6V0+0Q5/bkt2MDHn
wmLtCxeqUpy8luX/jlr0W8+iJ4j7KeiloRiKiuPf9DcUvOo675Xi6p9Wvm9lwaNO
+zfskX64U5FpGnxSt6sSTYLBBa+imdP0TkYXigSMHm2J1aogh4IeNLTarCFWQZEn
3xAhjrp/rEsVWGh7G1N4J1c83TtYJbPQTkfLu6itHPEyYWEcDqgnbPWyCi4nEH7x
jBL5OCafkhOenN2UPgV+//ck9EIjvDPxUIz1VbdHv8ycMiK3NeUARZaYBmWKp3zn
t+JChTuY25nIHBCgGYWws8TX/qUoFA3dGSo2inblYXmMGlLKzUGISKN7zpwmKcLo
HMkcP5bzPb6lnPBDa8b1tHgW4IGm4Hgrv+iVoedKl052eQ2BIk3/cYScYMVRRHoa
8hcBZgCYPm+2kwPLYIrW95BJYCKQquhxkTaKwfqL9x2xvEAbxuKhC86FctY5z3tf
fU/1Gkd4cB8SRakWM7246UEvwb82pmti6ZiAvvt2Wb9qRz6KFZAjGb09lGyWy6DF
wNpraUeF6f9N+avpox002tbXfWpvqbP21OhSKc1vH7v6UE0wir+ouTq5Q6V297bQ
HMTFCtinhpkj5S/tluV9SFp1pIQnvT2S0aisRxmJlDQEHUysFsWzXLMiM7Iub/7L
lrv/1X5gtBbDxCt6Phf9hz0fv2vTkvygSIHIkquHHXHip7B4/Y9Ny5sQvURU9dnh
ZucIck1ZPa60+fP35KPnwR4sguP3mTriIMmBxe2Bci3DkhOrQN3dgC3Vwr/cfiF7
wpgEGmdV2ZOZ8yiz0Jn86mIXXxR/vnv4nG4T2DYGPX13Kxf7Sdu47X37WvtXM8og
FI4V88H8vEFIr7ua2gcxCjIDMei9zEJUk1WPdijP2IllY7HMQXVTYMsSNj7t7zfv
2YP0SCAgC111p0/qX+2qrws6B0P97hpY+yHAwg7zt3DIV4P7RAMrW3VLo66Kxi9y
R6fnZmNzEkWwgHgEAocMTXsrEyv3oPM1jeI1AViBBE1VLT4DNq2Kpgg3U4VGNCui
pEpUVt1mdV/XoAMwph6vy6+u1Wq80aRt8p1GH5OSGWgH7y17Jo582JC7pNwdScXG
OEkQIeaeAhNDvYYLtBspkSvLtp3JTXTteYsxxYrS2xZrug4dU8tx/n/MxvaoTvCJ
lGjt+TmGbBhO0tVUkGwMuMXLQMAiuuiAFnvpvfBUhicc2X64U9fSxhjkJqHHY9Cz
VO5bz+fm88l3dZ1A4Zl4b97iXMbQuVxbtO7U14219pM+H2L7LDRjRs3yMG+QfCXw
94v28zi5YX6xYn4g8YPAjQe51CuXggdRgmI1tUFBOy3XebwsX0DhwAYTQH6U/hLV
jqbGvIvU/zFIfDSd3KRUA5ztM8GbSNcgq/2PA7Eg/S3WLXple+/LD0dPMuAcFIc5
Y7JO/rBkHSU2/xEKaHh42IR1PT60DxskedFeIc09ZR57EdufaL9BN/5kcUCTmjUo
QtOefhHjI0qbU2ZBV7Kf3h8sRMJmeDUwiupWHJzPtkE7HBZpI5AD7lyZV0psNNAe
+0QcY5n/PrfZPP7/z0Opz3AbV+OZieZYQzvayrSYZUsexaEKXXObg2fBzUM0xM60
yO+Tv8sHVkj53qBJoLwqskat1AZDxpnopIgA/qtZZMWTZU3XuV7w2AxnChG5fF/z
X3O8cjqMpvv1TmQARW2KjtCMeGulWL/43IJszpypFm8TDmlOeKqA5KeX77R1k78d
9VMJeR7T7DiG+jocw6Xj91rYXT6eYaf8huqqEvrNzWAPV2LDxSzkOgYESF7hHzEX
qCZ/LEc0gOppuZBu3LNaIUubT95XV3lH018AYae3oNLGmi16hjXCdU9ismLoNUku
DPMLh9/o/2/X94tSWroUNzVyh3Mc/lXHZ+YRvhe4k//FLfLEmpbHj3B3f4zTorjK
d+i9oWceoBO6Zu1UxtC1DWBwk5mS1gY1H/k8O+me7DkHKQp3mH/6UMCOh8/h5obu
nNzhGi3VxudNj159P/VTA6BVXtwfxOppwlIZAbPfPrX1gU5UMg+On+4fQjWJNmzA
vSFerTlKWFCZCXl/aS+Qz5PKCsoy1/dvTBC/A3v+6WJ5yiZucoRhxyaDxSpsIasE
IYAesuC7VRNVCEMX3VDjv+RaRMdYPB0v4isSskMBGDyq7izU59Af7fzbUejN2eSl
/dhRECZRKbaIvak5lTFHqP9Xz99a7r9eQ0pMAoTgepfdM31KYDLJeyLomCUll4NQ
b6YkFrj5cBWfI1yr5vdvh0UxRZgA85ynZt8pWGnmT4pJMi1pjAvtfP/nazGM3feU
s00FtTIFVqmRE1dm15d3mNPld9DLaEEzLleunM5xCpXjt/miTbcLSvwZrsqvbU+h
X5kVidZnGhUqgGw9MHKuFsxCvJm55vv+dDud452oVIIxXj+zphgJooIH5chr1w8w
dvRCpqZkdufI3VHWm/Fx/lskDomOzZGUN69EfqEUopS5eGF6+l9Y1pC/SmqM5UrC
r12vwbcdy9SBxhkc49DRBIS1HxUEvqDhQfHLzL1j3RhVVNl1Ue7FpHIxxdrvdy1Q
6oVJXP5RFHhyLpqqZnUshtcevh6SjkMg9U2Rz+H3TAr4Je2a33Ii0dBR6Ironl7K
ngrFjkDlOp2AR7c0a/JXnR4DIGM4lBEj1NDdK8vcnqmHYQxzhSixpbcdpuf+OOj5
S9F69te6c/QCd+1KzVxcfnoIUJTYabIqRXZ2uxF4DmkXbsa06UQXljVsNdLmYhTD
hWSjYd1+ohcfah/nW6XY6YA+F/vftncNWLJPL11Qx3sUbbBqK9eN1EopLOUNriuj
IIGV8LfxaCu6amG6qWHop+RUARH2xqJ0LOXKC0JepauHrw/q+PXNbAtAtgQiNKh6
frSB+Xt7J9J9NHzbA5oeU4v36tuDgm9BxBl7byVpES+ViUm84ScUa6MTVUnLQYWO
7V8CVrfHvlYFvZgRH3FAqW67kujTkW7hLTMbKrvI3BYOjr2+A0duK9ON4gUB0WnK
FPR/IjkcfStuogyMCN46AtUQAIl1BQa8/fTHibpKydvAKQT0LY7/ueEK0Aphk2Yh
kceGStDwQw/j+QXVIU4KVoXSPqOJiz2iGdDZIIQ6PMegrNGrZBb2IhJo+Mf5ZaiC
lYkcwZUZpTrJIp9gDsDo5b4ZURfCywezYP6IZe9zkvLatbWvXJmi1bBn4+Zws9Ih
014XC8zIPdN1wPJ3mz3z3N/hGDiJ/DtMVXKwY0C5E/gN5RHZk9ioAhW2TQrfgGz1
5+USXTFqKZgCbvND+pGIaY7kOvX+bxKkwot5l0yWtcCbNcAVGE3a81OMpVlC2wid
twlcAWFcleV7TVd4mXWMSInJ7QLrRr6GEdZpzac/WNmhj3aGshYV8Ult9uL9YxKt
OxXL9tkNj4N/lPAMaFe0X75gBxj1ljEy6L6mrQP1tuehHrQIbPoRajE9iMfrjCwN
Lh85xxOaWhlqdeP6lZJ11j6wAzdAtS+VtDMC45jIRZAL2HvjYr2XxnftD/ZxlMce
d7Kmsfk0MuQDFTlcksuXk6nn82ijS1px1lru0n1/ojjG/rqnrJyiJ0xASQDnYvZ0
4fTLQe2kxXXXJNQ9eH5bIFYlUYeOJXz4vZj0stUeaBuFocEUTrnKCQomBDAyrOAc
6wMoSbSf/TXvdCokQDkFUHCrIvdnPc2Yz0SiF6IfeKQsCL5Q26yB6hZhryHXZiqY
TKnxsY4dky0YGdkxn+JZ604bO4M0luNVJ5o1f8yuYaUOQ8iWsCxPnyjpZOixRyDF
Ji7ko8YIHc8+nrnmsmO+M3UYNCTPYL+kADttxDyobhC5nWiNqjgjk0Mz5ML34B9f
OulqieWs9Dixq/0jbOWaZvurnH928fHUT07MPuQDFKY72L3QR8GBJkZmnAg3XdQd
SzSgTCFd7TANQo4dqbKw8YBL19nJQK2G4xBrDT+x/XR7w3nPRH6rKgg2xRT2hzIi
VtedesERNuoHRkjR3/RPUDknPKhB7YEedk+zD6cA7ODom6Bz5Ho6b/n075A0+TtF
U2l0iHcAA403Ln++//Pvdkc1+LUFJa/LNm8fA5X1wJRGMz/MIq9pyRvy8I6wK8ME
O8SvW1rWitBC7+tKz1FzJDtapbC5VOQm5FTSiPwJNm5DDIPEo599qRaWWJ/cZ0P+
XsrnNwqVCTvU9e/uj1Bz7yz+vJN4W+uzSJlSgbU1Fe1CdSk+jmwfGBDbm3hl50t3
Vlk71LRGoY21HYh3PORM7fKLD0htNu05O5O0dVu2dL7BC0nFwoqIgFaLboaED6hf
/Ulng0VI9PNzG6PgJ0T6Jl1vn9+2uTOx6givVGMzweenXI6KtRAPDEemvtqEDh2s
HOmZwZ6dw0UqPVIm/TyLr3QtkY6LaUdOtq9M4E2bGVaRXHlzJLWHO3yjf2MdJcmI
cgg62U2Ts6/GP1BFqAPhdzf2pwKJAu6M8DNGK58c71VQUn6VAUGEmy8B8MvbTCKI
9SgsMHfvnyQkXELpQN0FY7kzq4sW9OxK1yyEL0eFjwI9K3MuERduxkGR2Aolzu6P
e5MG6vO9v1U7t2DlPSnuLuocad/lr4vD+FW9Lm+/InoLwD6dQcZ4I62nb83u3bCN
4/YMzOl3iGgVt1DyL3YqERjDukmJhQ+AjUv7r2+XO0rCuJex+JT9/BX8U8ZrUtrO
1yL2wqiEvuZHpSeEfo6mmVqLYMoNl0PDnDZCAXi7XE1vsiTB4cDCqJFUdS2lxxx1
k4hWhBbFm09cTsoIwEsajRhVTrldpCZGoZh+19ZgdAXCQWXg/kSRv8aXmuoEQaIS
vURnyvYmOH0IH3FNV4q5RJl+lFsaJ42EC/7tJNcvNS7QD6j1PXI0oHxMW60UlgZl
Yg6hYvxwpmCA95lSpc/iyRWofnglEabOwlGg3r6FS85rxEPaseS+QEBtYC6x3wPr
sCMqIX5FJXhmXWFPpLMFgX5oH09Wt/4ToONE1m8dBVOzHT54pKWWS/N1JyKGBPOe
fk4RVA4KvFHg+6wF3IxAdO5Y5l7qoy1Dv7poTFtAjvN0XLH/38nbwJMVy2VGXd+g
Gw4n3zhKeyPMuDpuVcWhIX2l0zrTwui0ShZJqDGe594Wrf/Mfx0M+CINLLJR4Y+c
6KzrSefErC/kqEYKKz060yilexptfX6WSyXCcoeIgrFr5Zccyebng1g6cSggikKU
GDuBjpdB3NUeovJy9rmFahpI2wUCt/K6uZX5myQsaBr+Ws/QVewKjf9iR3HCfr5K
H4LNdk+ZS2rabq1jQvLg3du4jegJPfNYpUWDtPIpcDz9YhHfgCKyYVsrSCBV156w
kX4FG13KIgVzR3Evh7w9CD7rTWaOGkt12PbjHnivDq01a/IlnOQSZdIvmU5oEDb0
daVbBcHpfK4RU/C1twjLEqaW5tkwaoWzTferz/F2eDYN3Rjp97JWd7ypQnsOw+Z0
OkdnXxx21WIvYy2si9S3LwHYIijUiuf8A+XOmjyzjwinNmSA7crNZBZa68kRaluK
MiG6K6/JEmoRpRP9lRdUCx3OYkRIwWmERGszXtsq06ubGmTeq0jYCXRWb8HThGkJ
acZzgctfyotNUgwWm6egE2t+IqF1kdeIP2deY1moV9GBZHV33Hb3+zo1wV9qHYIa
8DG7xpxFPoF1v0bwDcCDbHGBd2gqMYuWcGf7+mxnC4dVwVlEsX4TE+L3LtFRTph+
BxP1GEzoVH6ChtBfGExvo0JNB3Rg5Xcjryhcdehk6DuvRKEyneYzpruOqtL+dhE0
HuuT64Twk1gRfGaMRCeWFY2FaCQBRFNjRYYRsoSjROEt9Vqf/5aD+0IINGb9Pvvn
yFuDSpWv3GGR/PQdt5rLtcPWpAdnC+MQ/5Yy4QdSimHnTIMhOhZzMNRGsghQSpvc
5oVaPo8TS5oWJMJVyy0O+MpOeGCKiwe5WJQb2maj+ken4vfTeADdAMi971HSg3Lu
LyD0t2CCLPdqZ1hheEbSTNLx87gKXnTQ3wP7+9bKTBhnmtnlrzpKMIFQFN0xtQJx
U0qmL6QVlORjbvNuTsN9ea+FyJxsGv1hWoQuFKxjzSp09o0swpZL9iM5lECBu8h/
SYQ3jRwANmn5OK4B0eg1PQo7C8sYz147UBJT+SstHEGWy+3HaT76gsSAmMfRPGDR
0sZX+IS76ieDiHRzIXQgQ0PsbmbCZx4zUU7JaW3lDnyRybs8MS1S2lhfFjU0hNrP
6o11ZGh7eyxxZVsHfJPTCi7Ps9g497eIOEF1/DD5eMO8pGRPzuAGmmmttDxmwmrk
xMN7DdW/23DpIjggQFDEAkWBcjlMfqBo/jRTE7Hc5TFs5wCxAGLZ3xLyBlzAfhPM
mZMUqzPT02t5Shjn5cGIaWdLitUp4OsEvnX6h1ezpwDn/hG8JMsnUCTVu3+GcXJp
AGRibUohV8S3z6HTU5VCS+hyGD2QoTDTKcId+IxEYF4BJWY9E/4AEFiLHwhdIwWK
AjV/57z6x5pZV5HbDzQ4jh5MUXjVmMiElaMN/e3rLKujZxC/KonYxZ1pr7TJdhKJ
+zbigSkO8Vx4AW9jl6pkkpbtqpvs1CRY38CAUDd9i/xoRLOb6Mq3G6aGXBkyEXV5
loW4uI4/YKFNsv71F5oW6O0p3kEBGKMSZ4oddMRvx6Cpk4cuhRnW/mkZxq/qphiW
yq98CUF8f+y2+hv2A1zv+3Cb9olntNVClNds9Xo8qoU4P/bqPaWtcuP+3N4nwRI6
9EIGs0Ynp6nzJcJXz7wcoqPC11FjO8eqMUTHxV9VzOCSreweQb+Wrk1pva6hkqhI
GSaQoJqsWDEaXnj7BNrBESGhLCaszQm5FzE/DFt8dj9fPGuHWfyOXfrN/lR4PIDJ
Ri0ZL8D7xho6Ul2H/tfiFRCqNqIb17T2X3X3rvGTHFJHyrCfuYnP11c4tSSD/loY
evF9pZbew/VQDyCHEl1z539SHK91D+gComgyA6Vl4m/4zy1c8qKP/5tar3I2SHhU
gB5bEOFn5k6aDBHuP+JYPYAcPNryIA1BL1NXuox09H8xkHcLM0HHTEXA6BsBN8/J
nZAVkaWLMZRSKHoW+jgbjnTkslQQZ5SOzdpzmrYoBTvBT3kj8NV+5+w4XxXMxw+B
Xe2u4wO1Zf7LNpR7pIUpH8M9hms0bXU9cG0bqZZYr8e6vIRboRqJxzCoh5r6rB1r
TPyPHeUK67JbHE2o+PVvGfOQU+mqwE60gvo/0nxh+fuVFUIDMz+hLYuDJqyu/lwp
yypi8hi+VXQsQPBwcQM6rEHM94iXYtMu7GCQzNdGyeb7wc9pS56UWrEEKiZdK6Oo
mz20qb3fAcTLQE08RG9wFSLJrxJDIQEw08P9gelqu9J1nWSgBYvktZJj1MCbvDZK
OSN5/dLVNis0/ezJtlmf4/XgxKddIgch4Llxw2tJ7MUxjkjy3hvWVIffqf0qcD0U
E71nnZba1znAob7I5+R3eFT1F3qSBLAUDWciJnJISktO/BskjjWXp/IkeBW5kUni
5P/Ruj0yZagmJ8fz7vXofIDVVPsTVLatRCPprcK9ZPTti5VH8I8QzbGomFpelzL2
1hc+NgOnZBe7jhHcohwROw7jt4stc8hfrbqIrKeaI9QifzcqPJXZFwu0CPdo7LdV
klzKr/UwYeVu1jWD0Lm+7pa5jria6XEtbSNyMu82NK8iB0w/Id4k5CDZUa4qnZiD
HW4o6uKF2EJJ/b41YpLr2YxPyHwXS2fuYcYHqc5lwWs8OVSn8kOOcjReWQWqdulH
l+fl9PabSBbZoP593pnA3qq06ch8wRZUhq1GFckkoqdkOADDjevSXeWEXvvCnQfb
Uu+wONNGplPM+b/NPzpFQvGVGrp/viziTXdwBX5zNeWzjXxonkEGrkGQZaf4YIqv
yud28Bk5z+CHxy3Ym4UTPHaUajKX7OrqqEPTFNOVgLEpmNcXyqoKheEbjBkfeLJs
Wtvrx4gTomn8vVRBQxJn93u8XQ4Ls+iExSylSkl/8DZYy2a9IBZYa/piCAkWdTej
xoNeOMITZ4RqsP2ypdSMXl9HqA+hFvpgGkUXk0GaEW1rTUf0XRtMQO4ESvra0uhG
CoGrSoSiUL3wHAeuCy3HCHPT9G9m1twta93C5iQPVofs/Mw0Sqs1uutwKXgkYPot
YqCpjsEVorlOgNPvfq1fYmfGKgYA+Pj3PX3wY9XarH/ppwV2ueZ4ADuAb3fnMq+A
EJYhxrE7/nxOeFuoxxy4Y59YuOCCeozFxiIfWPsUvzTAzW89bWIpog3X98OMV9qp
U8yOxM/sFpukFQB5l9zuXsLIi0d6rH23F8QfqlTufxh2BJHU25o2o4DWqfQrL+Ax
kBlMGhwBjmzxoa/CajJ0OvwReHIjdcRbF5YpUIA+7QsbvlQkXjBgvT/vZ1gwDQez
DmkXCHw/eV38ld5Vzu7Iqp38emYWFqNfPQT097Z0b3KF6Y4Le5GPiFifjSNBde1R
nKS4e/zGg/+yxfaFBtllUw42NLt/1uHFlcj9TOlneoJ/s9x/0tJWT6w4uiHg8esa
nfxe0ijgCRsTmyG5RVPwmcBKH25chFxw1JSevBIvQcMKwEMLeytaEt8Wz29lbOYf
Ob/pcRKQ/tDYyuwBxUekuN/fdmfE1byxTS4iMbdoJOZ61Y6B18rhwcubJZKeFW7o
BOM6ts43RrwiOkSkqcqMs32IEeEX4GpNPOm/NEqE6jKbwjIRrBHSD4q9CUHrhpWx
ZibOvGiB+MngOKfcZzzVDIZm9oe9LaFj+n+beNO2hhw6NUL6SKgtTDcGnC0dhT50
sgiMRdJebkRfttjXeCW3mu69iN749wbHbwHGyQCW0OGE5qj7OyW7nyOF4Nl444ZA
pEahMU9FvR12fEZDv6NCS2OUnyCibjFb2C2YaG9Ahbx0mHwE86RyWLAPVpR/Ij/y
egWHiYaNizbfjlQwyhtR33odB6ZVQe9r7EJjG2ZrLpkXdoMJjM0TmkMp6FjhAixn
/soDnc4+i/QFbKF/RyhVzCGNdXlDeL3SfGlNxDzUtMeTbBPU4qerK+DtpknW1nIK
zeM9H0JSFS6MhabPTFUkN9LrHIZh+wwX+rj7zliLpEBm+KIaTNqAEuaBPKAtZ2DV
0b8CW8PICPz3nO7qT3YZHOAZlYJgO6DjACSH+LHiytIvCyuqBou7abUPvNnjDCiM
iNM4vWNABNBfVLePcL5OsODIczrIhTxZbnw5YGBCYCWk7dHjCNKfBsCo9y0u0++4
t6s76ObZN2iBf8IhdKbrOonDFNiBSdeyMYKcDZVdVy7pCqBZQ0Z0vcK+5jjg/C3K
w9LLZOEXt2ywVAOZXExvsfPhu3ZwNYZ9yo/LlmBFD1oDsvV87QbAEQElyRiVmSbH
ebleZ3/ESp4YoEjdEWofR4m0Hq0APQl0i1P+mvOsBlqpx1GIe+EjQjt8PAQRSQpS
0KvKQx2bGANRFgDTHG/MfxjijnzoXyqrXSBHsi3z6AjBFei29yXFCEZBHuQivssv
SuQv3gUzQcZprXrMeSLFfLSam4T3JkagigjNhJ2q5f7Cyp5iwXC9xfhVWO/s6uch
xU+z5IvhOQlfhFT0/Q5ihaVKGye6Bz7ZGDlR9uKPBWRdBEImD/PL+gy16VfBcmLY
hoMi7fhhh2pG4yt52MlJclvTw8i7yxU8CadkhcLUOLdKVSLj93EmoTKc/xaBOEJi
qDb85xBNNoYmVbAEn1Fwjfg7ng40g7vmOoHZ0XZSSvGx27PjmouR0/DCckxQItKe
TlC1N6IDwUCgIe50uflcRjkxA3CVU6lJmEwU5uqHuhCOnkUub4L+WhIJvD01B2UD
p9z5BwVQh6qvMn7OdMq7P5myBUkuviAkO5/x5GeTPI79SZmhY+2zqZymgV3s4L01
1FE2iaxwc/ay/8HSWyh3X7dnexkg9W11gqtvEUHP92t0gPJ6sbWNiDG3ZX7JVWA6
wuSXyPOwQZX5nijnwaSeMAKJYAs30DqrGY6GWVXw47I7T6pfJ8ywDZyqwRbtQstl
o5vj+rDruCt958Y+FSHDm7NVC16Q/rs+rAe7NdnE6GpC03zm7rwGSEcBqH2iCyaf
K8MFF+IlnMNu3jZJvWBeUvoAKeR/B1jqlCwzimLRwiiMyJEW3z5eyBwDDO6WUU7j
n7u5sTm3p/5AR57iWRZPy9kAhhaQOlN0rTC8he6e6sCzec7yEU39qh1xW1iqF2Zf
RfBxcb5jVLOcpBBX6/+vnSG8rBXYQTzcy87YLoF91eAWKsDNdAbr6b+ernpz7PAN
xXWkKlg4IWuUkefZc/wPu8upVOY16sA1zzHU1JNYcO8xyggWKsc3YfBeI0xdlEOL
S+ksCaNkLYKeWUQODQLKZW8vk9jGs3a5kpUofUZ8NARsao7+wvAXU8jRJUWtMi5X
xI6CdKrpgyLeSEOK+yFwNi1czNc0PErgmtOlcJnKINAl7Eqi173g+viu5FeFICja
MRaXtDLafFdvzWOCzsNmDevMJbK3UjjdulgI6N+HD/pD2+OK5y3FlXoNt7aDKOsk
PhxuUFcM2gwmlbFCjW+Un8uMyrUGoEkpM67i7B2+4e9A9qG7as80aUV5WKIeovYk
7ODVFIeKDF2FAe5gBzk0CSZzdZsQRL74rGLvg+j0nyt/GVRsyTtSma3PW83U8wnQ
aYfb3LSwJ3JlIdI8Tol8P0sIgk8wkTyKOMeqBh/CzW45r+LUhakPUHgclZScsbqM
hmpJPsn8FWdNtuWbbqhd/AfcfHn17UeASyabnVbCbJ2zLRX56yscWE5lqvRbp3Vn
kPCv/8V915bptsDdQCVQwJiYJC0Zv2dWueZMwB9/3SzvrAOePg1pQk0buTNALzZ3
h7Hu8pg/7gCwsx/AnfT8xKC/Icw8DuNhqepaaeU73/rRTW414wXj7xBwkGqfvpU/
G9xeADRgx917qNwJSFnrQrWCGM8kf5zi5vF73743k0eFjrdDYU099UQUsCut2QQF
t+N6jYCW8OSw/yUVAUawGGJ1v2OTyw6a16kCI+VBWZP1kksE+Kg3tQ2ByFht6UjV
6YZ2ka7dy/L5Mw0b00tDNJdmcrtqcqzYX4gt8TEaLGeLTdoOPaEEgoyRqrULEOSg
jaq3zSnyiRFy7wb8SmENWN7/XDmF2KR2fJLcRfqDlwuaFJfkKMK06H/viiCWfBDP
b2KtTfCWISJeieNg7zMGr/ThlAT47mH4kG1MVPj/PRHdT5bhvhQ7J65MvrEFLLQU
TIdIydf99qGMBpZ2j34pc19nAvqE/OaxCnuXujOMlUVwZ2FiTXNIJj3ANQXCY+RR
wR7K6vQtJqRaqdLaAjGsPO5bzkIseudLwhqueGH7VFcQ3VIhV60bBHg67y3Oyz75
GeSTA5/rpP77bKznJZJlGI2ThYjaYD7ziE6pUT4C1w0REXe7oBQIOjkjb/nWeZla
CLDE5rm3SdAI6UsoxQa2aDcKJixMNCVhzEWPKMThj5ADuX+sD1ZwjvtTz08L9rqJ
nEv5Fmgp+6h8fqkbQfV4swqaW7EokSy6r4lA0+O+9QEe+REZAqu+bNG2KYC9+l0S
8SH+FuoIOugivKyK49HPM+tXsWum8Erd6hNMF36tRi/2syIY2jUwB6Sire0Q3stJ
0F8sZW4r4Qkx1AtE5ru1G4UCqugIBZyHJFg9dbAimWKfyLH93DYipq8tWvKLyR0t
mElbE/yN+3PzE2xMry6qObMVurDryOftWfw+dO/LGdfe1YxfvZvlms5OlHyvkqAJ
yldxtNUeXKbVGJIeyVYspzu2v7cEQHj26FgWofWzT+T2hureb6pdMlrzm6gt2nBX
mbq63vqkzsN1AS6niBy1LQsv5lplrtiGcMIJgaRgS+FGp9cVGohb0pgYo2pP/8hJ
kKtGDL7J5RykG1fD6/vMX0dJDftsr9CbeJmHVgTbUNAKNA+CQImiZL/GJPoPpsrY
odO/NPNMy8fIau5Hl8uT+fF7/1cTgJGtqWVICuNXrAsvReo0EsiWeBVAa+EfRAzT
CE3S2P5dnIe/p/xhiaVy7mWCkoxQIw1HlBkImf05iVdWYWBEuwCLYSBABfTsPJe2
t0EbRYN9IXmOlTdExaKn3+N+Gz5gmbMk5OebU2wRzVllJNWmAfHmuJsdbB5W3IiH
v7qTFu/UIKAb87v4vy/wQkO+W5EETjp1uD+jUbiGWeCJrS+OcMQWNdE4lPXE+iCB
1rJ/iHhYkmHmZtAap7kZlvnsOo8jzhOFV8Q0AEYKLJ6wykTzdG/Nfe/CQZn2/l8o
UbZzzVeO9rLV9a0HwLK2SFqDBq1ifLm61k9Ru/0AZE3uvN1R732pYuJplqqqFfnI
emv+WXDj3zC1uDCNN23xKJH14r3sAZs9bD1Z/n3qvBGYrLbqK3bRJKil73LWEznN
M48x7xp7gFAQWHcL3b0JVe6icQDaUt7hgE9oO0YwMqDLQaELKA7gyNqR9Jkp6UQH
uKa/yfghaEUPGO/+pY3s5Osy3SBnOzwhcv+3+6MlWxg8YExA61LXR70hnCUeZ5WC
kQ7IVTtCTdhziUlYtPajFTt8kuFTxH2m/ddF8em9Bjw4smel2vlKuqOLbDAQapMM
9Ur6FEkSDI2K2Itm2qUJlSso/04DHIUTHBgb1QyJSTva23FER+IlaOGdoE2+7upv
IiEIaJ7Jr5cnwcjj/zhGobZgugFvLlknNGezC7DcXzaK0EaLe643uFwzecuP0u5D
PJqRqkM4tqC/Zrgc5nIKQveLfkR1+Y4eu+hHe72cx0NVWA7cgT5JQpfi84fFYYLe
B1B8LQuj1/0Sg1UbyDvXumApLwKT2VzWHZJKg8F6ualGA6Cxxp34LwRWqoNMVr8H
jm1RqhJVjWAvXw4iiGKjcfn8yzRYJXVB16jwCMJkjPd1jMq/SA1j7VQ2gfG/umXq
eo/ClcWckI34IWN8p/u8WCkjEocAhStHJA8pC3Fp4nCaUvCe3IpN4dMPN0vcZ4ii
/HpbEIS4tjd4/kiUaEJ9uLIaLHS5BRei2TEvZAiyAC+X5d8eOlx4KYTodouP4pAE
et3OuQgU3AWrSOG7uE8WueXJ5kD+kQ+AvZZI+a4qQ0ub/xfPIMgb+OMpNe05Y+gk
g52KXXnI4w/w8UMMf+Au9R+t5cCl63IHbT6L6c5q5cqFJZtHTVZ4LCZFn1dD1dbj
Er7x1nvFGDtOzPsunel9abnOMoUz/4RC8jHW2NsjHzI=
`protect END_PROTECTED
