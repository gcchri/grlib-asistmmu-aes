`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O4Nwty5p8A+0Wv77//f77ds6HsJjxhfN+P+uuUrP983a2JOw34jKfLoJQkZh8YyQ
aGShk6s0hYap3sTYGVfIbWcq6wEBJ5iQFbuhqFzJm7OTbAbni4Ej+bgUl+yaPvZ3
q+h/pa8csX1ud5t71DQ0MJ+4ageQRNatHLJ23/YmAd2SKIodeykVITNPQD2fxj+T
tW3rG7RRu/S2zAPjgloyyeOLitWL5lIIw7yRbxmUlhRXUIdZ1x4SaXlnuH6X/5lh
7kxMc+LKb5wXrE64FDQTbtmEb9alfzjqGj/wB3SfyRFMjax71XTfQYDXw2bkn81J
`protect END_PROTECTED
