`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YLRIiHwE+2bRcUSQltMMiv4U31l738qlJn3+0CTXNORJfK/cwJASqckCl9SLrX05
ep70GnnZLiJrwYNkOAVrziWctGZFopkP+23W/hIf/Qk0lZ0KvULtdDBZK4jALLUY
8pqUetuIVVJbySK2DKUdXf13ywHdZNTafgsgQHMrnkOywvxthSEZ4L89eilsij4i
RfDFbdAeSew1Btm6LULfW8q2X/IBf3cp0dbkes51lHLvVikd7f7bRS44LWD0z+x5
6N+Y7r+WYkcKYq3i4bqcYlQPknnINjlFjdWL1Jw2B0RjYI/84Pj/YZMCm8UF5hjk
2WzA+heoXhFywn1YtYOD6Km16quuG+EOO8WmxhaQMiHf0TtDyTNMhk5VZb/TgBV/
UQPIzFY11pq6ymtgKk31qBgwzLZJjc7BC2ZnHkZHFfbWkXSvmbR15hJc9fkF6Tqk
vVBRDQB03HYEGXouIMdPOeqU2rU0xlRPk3x5dJPAoUXX2DvSAo7HdLGOp/udGtid
WqbtPQv5x6Wkryy8/gx9afbEfChle57dp8K5I0O/HLSlptPmb1PFy2vNdSAbp79G
HOM/XC6fEbhhTu2Si0w6Ey1HXYHPqJ+GwK0Beavvbux0qftVQ5VRJT/a5q5Wxjrh
E8WurLthQZhLxquZgrnTrA==
`protect END_PROTECTED
