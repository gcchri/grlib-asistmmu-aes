`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWRimqI9/y1HDqY66HJsnxW5su3KukftoOh1vphao+N6l7GtZpgn7eiUnp8t72Jt
9lofbBpHa8h0Xg68sItFSct7sIAWa7gY5WYk8CAVh4YCSvLO7HdffawUK9RsLhuI
ymiHF35RM9f26ZGBxptYly4rO+e/u5DPivJy0qkeqiHQ2qse6z83dvLrTIo91WmG
BV8JCBP3s3ITK3rQ9tiIy9VaVoFKRUTSOTIT5LrfOPXaC4L8MG0aVTsfVQZK9R/x
Bc/Tf83XK/jNivJ/uusJotgORSGtsuG3jukXEXwx4tosSG0/6zIi9zjj49Uu9z5e
/EIF7ch1cHZ3dSY57i+n+3LgDqpjo2CLEPBSuvq4707v2N850L+XcuuWJ1Jd0u9R
ihsqGcICWyY4oKJXqqoWAxhXRIPko8HOjFU5PH1z1TZ+EY9L+BsBjmSXga25Bhre
9AoZ/ELX5oUjFalMHuZWIDQDpd+8xGWWh+rD2hvWaf+EUVW7rKY6SLMlftVaSqON
`protect END_PROTECTED
