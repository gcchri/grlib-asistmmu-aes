`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rcUc6XjbJGzr4MgMlRqZQUWwo5hwDQ07U1Ri68I8RHrXrFHbOO7GfpTXVZyV8V7r
yhtmn6WucidngA+i4uJpmhNGEozon8YbEu+yI+L1OKMfTcg3cJz+TOHkZMQMGfD2
nQVrO3QaYlpDU1jg09DGcMWcbsJopU8fT4KeTihBnbqCySvZxo8cLB8cRgy+rBLM
+AsmzdsR6RwMCBPMTAMdJ0AvkaGZeoI4ilOYR9B6ILUyDHb1uCnQP6F9Cc5iXQVX
EfMNCvW2iKzzlA76KLPNI2Z/rMT3zf0msn0WOo/zPfFCk9FqSV229Uy5CiexYbwU
nEE095opD75CBtcVHu6fUSVQixrUtumVow4T23BP32jh3glIwPh4JEfBYdhY+Xep
sZhccTNGLR+tm9e1xYlbKHALcvmhwxa20nkwS7O1aGcZVN6Zu8wWSiUs596ETDk0
g+RVeMehR44y3synE5AtLy4j6KtQ0DaRLZtBbXU5Ejh5nOlqcBDKXoWdZxmPDrzd
62YgQdXhtUnWPMGtRkZ991DE5Rxmmh/lMlBjgDiA0SRMpl3spZyuJmx99hg0GcsU
eJOOVrMwYgDO0rORwlzEY/Tky5SKwRyI+BL9stg+KrU=
`protect END_PROTECTED
