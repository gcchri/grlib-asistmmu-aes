`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zs1NBsUQkmxFQ5FZDGdFFephEBpKvwiuj2mWym0t8luVHOetX0V38lNqNas8kLS9
OIk9rpl4s3yJyOXYyQxH84NalyV80/HUvGOMFpJz2FiV3/Nd4PuSv8+16+XpqaUD
L+9kPwC4pCThysHD2oBQ6xwdVZLs7+8zL4PdtgFyE4NIuZHE2OSyNACvCRiqmEwq
ZWdKWghV4SHQe311NjxGMd75NwKYc09GEoYRzKUDw0ZAOweTsU1Eys/L1CptRTZg
b6RnjLVpEYCLY/vJ4A8a1c64rmJk5bvBiWppNguPEgAQRR6ytg1DPZs1h16z5Uva
z8R2qHkWkGElr6d8sDVYMsUvL2leFHvOXxuIXoYURcDAzZJxsbWNvl47cgXZYqKr
dSFIEE9+EV38RI56IBMtQbugoIrNUjNtbUmBxUlGKSvxWQCPblYlkvjdeefjF1YM
JLifS7462I75GGs9d+QfOv3Aeiqc6GHkh7Bfq+7HXq0=
`protect END_PROTECTED
