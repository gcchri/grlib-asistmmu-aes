`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hb8I1pJSP3nQUrZISZ0anAC9U+n+JM0c9+TZPGma0KgZ+LrErMucx9NIyn3YVB/h
FxSKWcoQMqEli0nRzGphYJoOZDHSJo0RxSvmoNgx8ghKRykowQ1XO/0O3ppDKHWt
/z2egAU6bagZOhCuQ5Zo8Klb2pl2BDxQjxO6xP2LyBgmHZIgfKW+tUc3RoXgAvM1
IkfpyRovrXGJBtQqi9Ji1n/zS0DjrHyl6PT7DkapVeI4aj3t9leM2aGbzN7ULjdR
eFDsIQgjfNm4x9NeTM6b/EDxCreMnQn/2kEQaWqqQdX2ENGPzoRCQG0X8nPkS/QV
4Y1xOC0q+ujadkZYfqQmRkoasFlimysJGWFf5zUpCCbjYkDZbU3Z+k8n37Rq/w8H
KPA36Z1/yIKolTTwOeBZ5uA9E49eamfvacu0JTN8Di56ttes67ShboNvyLTWmwVG
oHZMUyLxQJm9OKCIU96znTNGn/YPTQw1+8aG755Tm7SJsQRcX+lrT9ZdFLPTwPzS
xbMZAhBbArAq/6tWoszbvOaxRjE9n7D8n/weCueE8iB6mfm/qF+/AzyhziAaVh9t
WJ+3xN5f8OLEwTBbx5KdyOR6Rczap18wiwNUbsK7jlfkLX88utufa0PwBJyVOQrd
`protect END_PROTECTED
