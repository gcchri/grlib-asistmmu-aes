`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cx7uccowNJXzFeuyLfQqL/An9Q1f4kaa9/l0ZSbzgIiG07leqQzQf+uhsUeOHLbd
gnjRTZyfWQ+SIoKk95aOPmE0HLLMRresG4ZRJ0qOQmSUAlwjKAGJXBlODQHgJJ+G
jqDuDqba5n2vMY+zMXwmlHmT7r37hQM50DCijtflBythT61mp2UEmUZGdjklFPlV
7n7rrPHFqzex5+P6CCAhZMrEBHOdffD2Qxth0UBkCY8S0/Aod4Gpa0TkcOHhKezd
EJgeoy66eVLwLmZ5b1GlKBnLKR7eqW5X3wdIwh95rJVc6h3dX1TIYdKWua+4KEFR
41clPMrG60rFIfz2i8j16qukOH1rMHfj7oZAmWUitGas5yyLqYmcOpNEImoete8r
`protect END_PROTECTED
