`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hA1wEYLorfPTvyrJOkBpOJoMXhIdY+KLUtE9t96g7dvBYuW/wBS9ZPXns8z3arNc
puPiYY8rtT3fadecPg8E4Oo3wmWSyK1IUHuRc4W6Vwkd4wDeWsQeUfncrkrf7OaC
5/28oVfkh4Q7Z1DWqpCtGiIRFWOlN4xDiPMNMwNe/6MHG1o0/61sVjgss5Glz9By
cC7zR5g2PTXZKcFBeQDX2YbJ1tmf1t3RAASeusXaECgd+93Ab8cMMbO8zCX7NxSf
eCGiZ/NvTLQMcZOeoB30690kRvvEUDOjrUFuSMvx+SE9ayv5fabQujlhYhAsYWlR
G343V44zVijPjT3ObctKTWL/iF5RzqTCsqCN0W+rE6W19gbTqq6pBsV0s+Mq94lM
lnSZtKCUKWknhBhRRgzaxNmZP4oQwVUTNZdnPnKsjlYtPSbtjII1mK8ck8IsGvGU
sYTmYNRNg+77DChskHAuQarcma+Fa/RmVaZjnX002L6f48PuZzslvvwp2unAAWJl
yGUzQ1CsnfrX3q8qhNKzQyNBEaMp5mPULN3kk/vxU/HASCKLHQNHXFFkMW6ux+iB
90m3MPMrd2/jxd3sLRrep2iKzR6ktIaAlC7Eas7bXKchMnOUbszmcxQ3fAVoAkXO
OYht6bkCdohQD7d77V00+cC2OJ0z7O8Nht6O7qm+bCLDSfd32ZVwgvOdLpyAbsMy
fKlqLDSbxPYDWOS/DsIzznLyFNiolHoNOiFiZctlm6RahdCdDuU2+4ycCdincGzQ
xrxLuH9yxObT20XEJRoNMKzZbi0+rVbbEKZwrYorY5mblZe9+FUTm7fLuLgY2U5H
6X8c+ODufV49c7B4KMsW0oCusVCTdM2RhFhI8uNWp4vn9Yq5XfC1HjErAwjifnAf
IOFydLHAht69jzE54aoVHEZT5ujhdTnzeCize5x7isQ3THnlLvRYb1BcD+s6Rl5W
U0sYUuTs262FLnWY1nLlERRLxqgapfUJ419U7QOSI7UO2+56ipzyv4OJGRenOi05
8ii0B+/pRGcNdojqG8FqT0Wf4TAKh4tycctKdLGMvGWwleFqIcW6iHNqhF4dS3DL
Ck5gt5pD/WpGS3ME6AKJgxRUArIwA3y1mRUMgpQLRCNZcaEh8Lcl+as3fZVJQByg
a69dTzudveTczfsZP74e9xZpSTb+LhmnRTEroJZdhVvqv1Y9UC3OLWkMEMuub4j+
UzQGZjlkRz1Cm/dfyu9m/QQVvlAnCrtq0FQwJYRDJiOILGg8Xm1zFyUCNkKEqhFE
qphcs/l4PC3AzKXCY/6+BKfX8W4Bu7Vwo1kzz9vMhYhSRifzCc7U9pWRULz/Bmd0
RV+r7ORjiTm6NUwJJGQ9WnBit8qCGNXRV78iu0+nznUhUFEHkyQV4moBWVkNZsmV
uXy+h7bI29ixYFYbcz4fIA==
`protect END_PROTECTED
