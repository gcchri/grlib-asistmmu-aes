`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0LAjM54fQRph0Wzb6Oz2qDFCYryI6B4oKDeeWs5yhODjeC1qVBHHnumJAVyZaon
QpIaUZq+2rb+njc7ScWM5yC4SGiZUUKvaRM/5AmPzjU0YOtECq3xtA0x/gSfYpMc
BtWxw8Aq3pXcDQiMGWEawSkmWjjQtDvi4eHWsQATqpUZHWJVi6xd2KhMDdi/+zYn
hQleHjiwvlZIpn0mvg2UryDwoq02JaeNeF2QOWUnE7E4hcg9vdB0D2WkZoNw9pqv
vPUezRvdqGp+9QsRVvtAphzDmCYuOx92BDE3I5ETpc4gnPAcergF5QoUvrF/elRg
fuU589800zuMEyn4gyJ8+aqS0rf8JR5KNeiYlnTD0nVQtPUQ3X1/cCcftHfEvMFI
3XCiOIhrhZzLr1GWwoEqwyjoBNEZbigYovM8ZDHQwpg7rdrqe3DZ++hItTn+DB8h
QTFuSKBATzvmijYKhugD/bG6BJRB9owq5HHid8oJ5czIkNf6ZfzeJ6wN4MkXbfUa
`protect END_PROTECTED
