`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AAlmJLw8cizHk3VGN6XJYX8nq9eDr36eJr1aVH5kKb1DJeMkvmk35VedZav4VrgN
vNp5wFwIVpWFP66rcAs4NoBGbGuqrGsOiD/su8yUMhJ9VWjU7tq6Y6t7LM4JsNy9
8H66wYGPS/drrFUrIX8WV7jpmCTZ1IoZC1il76/aRYrwyvogktvnhlbesqpyGwP7
0+ufXRyK+jsr26m0ZuPy5hXv5gzxMMlx6Da+RiATnU+Mz3b7ozemiB0AHn52j0ke
0W+T5lKZGgm8vBG9VugFSvhKEzHyJMdVlW3bmCICCiPYCZElK5uco1sjBHFC0Z3f
DD/rg5cgoyvmpK17crFZJwbHDJNTi9bXI59h+fpYDfsDjG5V/0AmhyhNmjJ7/8aE
YkGtDP7YLSk34TwZ82kevkhwPCgiCwoSjagrW3GdvJ5skyaSSlfQ+Y6TeQs62n/t
xcTCIPsslUM6Y/6jZTM7p9XdM9d1h8HoejulyvPrWDdlfm6KEbNBwulrT/g2CUnx
9ega4bEakLMCTWoVQ+jzxRY3OFNXSUI2oML/dGR5uppg0K9qxxQcxSrQzRs1O0pZ
yyFLvhtp7oQp/K7qlb/fsw==
`protect END_PROTECTED
