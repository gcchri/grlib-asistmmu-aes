`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Q9qhtBH1hAaYhsh2Hh0Hz0rlRl7+TKwfQ6+VuAr22I1hEqOoQ0ZRE5TMzNHlXm2
rnyTjCc1oFQ8ltwaXIeZ0WvkPK3sBLowQMjrRzPJeArz9qlJ/xoGScenZ1jbOESW
NH1SpnV8x2s5aF6v8xmFXlb0Z6Lm2V/YkBQ03jpmVAarx1GRTvx587jHvp24fUyt
pDaBir32Mf4sHfz4l18Fgh9fCBnsRjIUNCXOLwl4+BzfJ4uuU7FDEZIodODCMeyM
hc2hYkbRo/MLy2nK+x2dhJs6Z17TZcZkHzJO+uFiT//BEz2gsiednsOb9FNT7Rf0
rh/g018HhbpJ03JthhKM2guIAG2VuWU+tX9+E9EtQYJouY/7bbyEhAGl7g59d0Gi
96zg/XUJjM+BlDyI2G4bvQ==
`protect END_PROTECTED
