`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+yKWFLuYvE/z99tiFXVI8T4lDZd6W8yi4txhZVWDFDwQ1SmjspPjFHaN19nJGqv
KhuSj5etqHzVRTqE6OabY1lrlzKZsRLFO0V8llndQ/2iXSYDI/4dkZHPCCOwMqvo
jnZZXuUYVLtemGGVqlDQbmUcd6ACveZewBlDTAb1rjGIXdn6TT2zC7Q53C4CAaNR
W+VgEEf3EvWiHqo+83RF2D/DFG3RZIcCa2jwT7dWYvXAb5uCM+qTLURvqKzPgh6D
/4c7ia9Ohx9dtYxEqiv4JQ==
`protect END_PROTECTED
