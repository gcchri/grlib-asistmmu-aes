`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LKfVswFYtoupnaFuKmRkPIqlp48Op9A3viXvsi40OXd33I90jpv5LF7Vv9TGug1
X5QKQP6ICby01XrpJhJmNQM6erIoaamio+oKHrNhE+pdoQZah+opr11Fx6YGPqgB
HvjyUXA+oUsrM6bupt6EwyBkH37j1eTGcTvHr5+OggvqXRejxx6mT4E4Uz6XTqPu
4SnNzTaXLau+kMwS7eIp9WdU7pqDKRaJf11+pyVIgRCKvMIa/rB/lyyamesuHIGM
o8JPTph21gAXedfIcnXL4ALXoHQZyB88UzPa1FPClL6Qm0waHBHj+fQlPkOoMaZA
rzSUFWKni229683ziyVNbOLaGGYriqyc1T23N00GM6ab1ZYbW9A9qOk9OPgQclPj
VWoEpG7f+AtMMmvCOBVoD6vwkna3vyIVHoqvaYLq24hgNumXYNVhhPoV6bBd89QA
/bGmvOYA50/KVRKmFzVPc+u++Mn7yFYZekf6MruVbfj5lkvuiRQR1lmo6YWNGnw3
m1I87XmXGwEJBTQsXbo8lUsIu+qKImYHvzOBwpUewEwK+kOcK++g5+syHiQ5EtHB
IvvU7mEqyn0ZemSX3vLSl/Y71dm9cb+nEg8mkf6Y1U9AoiYOtraMmEaq799sifm9
gvZ8I4Yr5vgAlqKznD+7hktSX6XPvv4hgkzMYDGL0woKmHt46mqbtRx/iAlLRvc5
0o0ik47c24X0KIFingsYFgDwNapJ73nSZKh9KhJPD0nHqbrJSuzwMeiKXiG8RAPm
+wt3MYbAn0mYipkXan2kJuxxbpAtVQSpoKYAmvxJKCbhUuYHhXEVaaHc+Arp+y1p
J8BO0gyhS9orHMlJDLfNX+IPfZ7OqbcxiXQrjICuHYJs8nI+J2TWR4gceTN+M3wz
fgOFLNwghQa3F+Ai2F+Vr/FlkbfnrhG02mWTu0wQ28ByA4fUwezM0epgdJXjjpwT
gCUM9Hrec18oXbBcuLW3gd3bB2xLbVwJztDx6VbDSZTuA9hUsTbLaYTedK+Fbua5
JzDkWH0B/jc88SAhvFRrYBl2NSTUmYuXOtkTanGDTKK1xg+Oi3Iqs2S/ukbBGeVU
ccKgRfgbIZzZjsDgBKhH9oqMnqiDUh0c+NsIfAkva++jGgxBIzB6AUHmhgITWWto
fBCC9Rj93ATP0ewD/a0vLMe1vpyyKZxv3mOny+Ekd8JvqRJhWR9az4imktpLl9KL
yfROIqBQd+m9IN9N1m+UiK33q0VQCvX+1xcARgiSYlPq2XtvgQwX3G3t6am/p5IG
36iPmR1LctgSi3kH9bCcMSllNWd3bZmHsqrF8HoB0rUXJGMcx8q5d1OudiDABvsa
DGgwDKdYeQO+EcpWZ2annD55ozYwGgxVeNOzArt8wCCt9rjxnTwywK8QQA7FrKH/
g8btqwuupOHZ7ThzO6DcAmtieiC6xDt/bdH1JF34nKMQHpqdo4hcBJnx1C/N6nqo
vlTTlwEV+mjQ8xtOVRZ87rSb7IHgNlA5vpInrwIn5dkgypvJa+G/T2Rj/H5hl7ck
dqF5VPZydj6E9mmui+hxTwgrQtF5syXIWDjk9LYGL26z8RBX9ivdJHij/b/+YHsH
9IkUhjWrHH2duBk0ejy239dKrmXKWdKVlJjojvEXIZf3wDADy8dDRSpKeg/n5HF7
Ezm5CwovjBUkJ2zr9xUU2ktcugCD3crrfKjSyn6Z4dpegfakWFYjizvvX2sElAUT
ghzuToTrSzU1B2AfeiipLZkt7iv34DeobmyaW5CUcNMx6gQZdwNIfUET5JrqWdF1
mGYdBB9mchRDudpE3D9T+7+NZqvutBR4eMX/NqLUPbC3rWc6Rputl/OBHpE/dKpr
2kILgaMymuXRh1aVG6IVHaQPMcuaU9atEgr8Vpqvx0ctIHdl7XnqdDfHZFk2hmhc
gRyj2yYZwknUqP2s9mmTAKa00tGAXxyGSGHuiwukFu9CTZJvhxb71lXFMIGoF3X2
LWjumj9LOIBPkHhXIZb6wmOFC12zb0yi7ZsII8fzphEUCtKhpiKYCQS0hpReQ8ro
7chxeo8rC/idsrvi8m4VukJDn8hsEwHFwJr8ajvnzvbLU5dQWrL7BPSoD6yJ6xfV
n6QCPClf6BwkUD4xBiKx1bch5hM+4vNCbgq4DJV9iLcNJV/x4qM3h5i2O2MvWSxa
2vHc4Kqi9xU8pLGVAjGA6htMJa4FMJnUWXNh3lenb0foAvqL3+Bc8qsB67YDeBne
71Aa6vBGUXMaAWHAMeD8zVXmKTDHDhRcK2thQ8HIOnJHZY6QNI/HHQZKFZxCdrIr
K6kWye+CCH2UJGk3WLK0qd/GsUJ1GOIuqPq0zHMA9rH4mr4+aue13+S9Ku9OWMy7
zFx4Q96MkMg3JTxICmjlK5gojjmMKmb9C5BRpfQhEb4z9Qon2SWzDApyBcX80p6t
ecmSlGZCcs61msqfxsogmQYYI1Ue666Pegs2L07GLZINfsE0PHvV+fmJxge0eNrA
q2Y0hZAGhcCnY+4CzpCCybMHYJYHc1NdgRhtn3MchcxDjELHhPsXQL7evWYb/KaV
AzN3MxlqmxDCpoQycEaz+n8FVxRFy3k6c6gDiM47aExQDTyBqshJMPTF2AzA1T6b
+Zp+QnVy3Qj8cchyWWsjnXbT0zRhX7MavY8f64GCSmUbQmrjU3LnllZ4ypbyPrT+
nmK2lIhOvEoNxoeo9VBKGSLj18CExVuYUKnfLgxqGPhXXwuMgU1AgXYXc3C4mdXB
iqr7pGEgRC4JU5ZhfzAvjZny8nb7C8hUJJnLYIyVRGjUn6LQ5HVFICBH+Ln38kRQ
xyeKq2Aaq3hbznmd4N3dwJ4OgfFiBBGgJz23m//00ixF75kRbLoPSMT8ZTkToEcJ
`protect END_PROTECTED
