`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKWrfO7tOCB/vW/nP1+FDoV9VeRX8Fv2J2X8LK4WVo8cxgaN8tWsArGsBHdKrpuK
pQOOUp7qS99D7En0IlyAgaz8mBelgSNC0aiovaYLyiNJOFh1lB/BjIlHuj8D3/L0
82NEuyev8gaIU0y2mq2yeTzIOE/pwOwVAH+Rmk+T2q+0aHigK+McpgNQ3Oaz6gHG
Yvz/xoDGR05oFFSpQrdkY6oCF4L/J7Yl/2nN62yPW16GR78Af873o1IRSEhVmvjJ
MrzAZA1Ye7g3921GhPzqjogTLXT6cFOWtvZ4qccHlTBkgEzefJwBRn44IZ3UTCSj
FA/9s4F2zzN6CN2yua+/B0DKLSOimGQVUCfyzLL4qryDqzELsRFnEz29Ara+RI9h
St3P+gX5HBAL20lvFNN6hSVbFEcIk02DEGIJL8V4GLSR+3lZ0rGvnupAweo93q7R
LnGAHCeDMGpmRcSL0DP6qjMwCf6VohxmnLkgPRNRubeHYoSchdvSeq6e4PJnd4VY
CFVrYr59225OwTwurmDpW/NFDX5XmKuRHP+ytFATYOMIlTVR9KxeYijgoSdGcLEO
TTLgdojgDeCuJb9IscbvSWalKNSB4dKn+VioyA7LBPorrtxC1+fxhY7QbibF9yvL
xUYMwVOrzp5/yj37wK5JFT46aRh4AE3cH91pCDw2n9bf+uw7fc7rc8O5Fn7uTOCT
qp3sAF+/MohlYrCFzat8aHE82AK6VA32l6UeSYwlkEtlgBLRfFjLOK+uf5KKxRSE
/7LQZWoGn/oi1IKTmAupwGPo9qkeNMCCBoxjk+xrVi54FB5KOBvA9P/csYMqSCUz
IuieJbxHlwJv3DPwqTgToxYkDnNoYQutPROT6w+8/F6RVhBaWLE5Bc1VfNcWIPXx
J+Hd3b64tEjAuwuXn6de68mOihAYNXWl7m52EBxhGZnNcF8K6eL53rGM7by3lT2h
y3xxOc9KJfnzA15vy7RjLBcp/6lRhpgXh5FpQHzJ7AEZIEsvrckye29uzXSKH5Ni
/BgvQhjwUu92MZStcHmDZU6gbjnxzBJPtRRAq5ATOCLH7uy7w/QGSog5a6dSdlgt
1eI1VgLHpHz/11wv0D8GHJKtpj51zpHWUeILceMOR3mRkoedFi0RnbRMB7Us2Lih
JFr5kSVQKL+GVbJzXU6Dy+O0gVSPtBvIgKIp+5wAi6GtpV44kHcSALhxeCQsGbHQ
rFpSo1EyYO3uiWKDdnf8OKf0NNOSAPEspsT3lbF4J/5gwQHQyQH8nqK9C4VLucu/
N4VdY0cJN+ah7rIsg4nTeVANXay18Tpzsi7zKCrILSnYKIugjJLTIx5aYYf4Ntpq
T55Me9dS5GaoyRinO/t8b5pW6QAqJuSSf7NM1YeR3RqE0IIflfIIFxBKK/uknyin
O61BT2poBAhm5uLHQmLuHqK/uzWYK4C/ANclSaOJ8Jfuto2GIA4FjfHG5EDLx/om
L3Lb4sL2KqXbvalhjBUnEA==
`protect END_PROTECTED
