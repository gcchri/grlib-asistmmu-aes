`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7BsY/U9Jou5yJZ3/eggf+zgZAHucxaQsZJOIpXoHP75jWluKpo9gTO1ZdEGqjaen
DbD2ZN9t0qsr1IFqFdX0TmJQymDcT/kqH1b8JE4xIFc1ocn/+9FyYo//f+r41FOB
LZbGCQTRAY/EtrqgUiq/+ZXwD7QwX2eImwOi1Ry2MsEMlYnT/gq2hJstYDxU01/7
L2I6LZRA7/8VrfFtFAilXDBC6gxIBb0iqcYxPPidJO0ub/0ZeyrG4QbTj8vIoeHT
xNzDghrQDo4HSxwrj4elnQ==
`protect END_PROTECTED
