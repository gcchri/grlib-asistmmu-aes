`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Me31n5W3IE0LzT/jzUsa1Uxyq8OXu2JsV/cekg8v05R6515gOte9v0VnyWEevWyI
9i9Szp6CILO5yZ0OA53l3oQtvS2wUzKbfQwGqzxybe6s1k6S++mtTTfm4sXtSr8K
MfPlWOwcelrDKPpdFOLo9Ik6asIDWnGC/PoOHU0W+eX4I+IqhYSoOqDwa6/FWIfw
1qCxhV0h+6TJsDYPVXo9os4eDucrHWPWOFkutNj7aqMGwoC0Ijsi47haKPirO/R9
JRpwXjIflL63ZmkzFV5KK4SKKTEKpsBoLBGV3pdYYYHO+kYX94acDjCZEBK8W/ac
UekTtq7AkCZS4r6/CxvfPpZAK8aPQ8UUhVCb7W/1FM7+jBaot2Q4A+APjcoy7fX7
bvQlTXhL3tfufTnd6ElvlpYcC1X7cBXUl8ufcvEj9qOz/7744CRXsK5Ms60/tU2f
bfMfIcUmI10a2m9bbFg+kPXO55642ak7kf+IXzyqIsc=
`protect END_PROTECTED
