`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDd6oWu3lYzEVZDAUR+zvB/Xhtz5gm3t7mlkfRRlfCHpDBttgqhcrahz1j9QeMKx
UxQqktwQAVv5yA1CZhKLpm7AMfaaaGduS5XTNV4746TomkbQcDlk4c0x3Q9JwIZM
+lVWrOQVEwfEVGN+HbJ3zhvyuILJOkxXAqfC6ucu8Hh0JpUSpVPurGaOpjYEqiz5
+WrtAdzwbSjngXlF5IwlNvkcdsacylu78buVbrcxd0a5H8bGlJXvCkMIEQRRlFt9
Nwcr3YalSjllMulk3cFwY6siYriFP9zCUOJ9WeEgkexyuFw4pi4voSbCb8JHr8IW
YuZXpyPqx/jJN7jla1ZJkOR9A6VFuxjVp2LUsEomGqipUxVDB5FY5qsadhi1kFLg
likthN9DrmnGqIPTLUKCJOChQIN34IFY44IWClD+W8xY5is71dEos/xsZlfg6Q1c
iWVznQZc1M4i+BVSvWdc3AEt1oaDHDFNyKwb1PKEUGwBn9I5vJC+c6l+gkWdgRWb
YHZgG6+SV9koVA670Fw5H1DjyR1XNYLyvLocMq9od7ZFlZgpCo3CAYDLfEFDWUba
rmRQ2C5PJS6hiJ9XC8IgLQCH9HLi2gzDNFkrWg+ljCedXgulOj/Tea3NeH7GiTwQ
YIFW6QY2IlmFKR7wvBh7rMU9RuBP7T7LfU8I+M4zUrrJfsDlOZ3uLwI74QOaABnG
P7w/vDF4hdW2DtdCCtIOD/+cPxzCWym7K0iRwZRaANFZN353lwRXpamkTaBemEKa
GkuZfUtsOpy7dIHhb5F1oq4jZtuOfHpcN+2p9w3ruKMSwdFqSsJ40EbhLFBOk9n4
nxrnl5/CNd7zpXOWTofN8oXXDpNWupETNX7w+9PVROsv4TyAK7k0ccOoegIToSR9
dq9or5/s5drch9MQPQUQAJQ8j+6JZ/w1ekZO6oZLCY7ldyOIVkKZ3NrG1D42918i
eYaSR/fIyAqGwCRoQJ02RQ/XXG2X5XBL4jympSFPHnxtzJzf6DfvA2NxhuDAdcU9
2kWcmkl9qBRMweTYSxK2sc4aOV0rQHt1CVCFxYfFW4mHA4GY1PR1qoEgWnD57Ixf
3Z5khk+XZc2I2yeDDlnGLg1DuM92w1uYfg1po+Ou1R3ICbEzOfDEg4NRkS9PgOpX
hJDPSxIk0MSR5Vw2ojSiz7rct7J8Q6nHmmKM6vML0xw+5IYVqHlnjt6iM6ZYAk46
NoSwuRWe8BifV5pHyquZHakpSsRUmoJ4MIxGRujk4HtN7m+YC6uzrVSy2yt6Ccs4
hn+4I68U15jYs7yrUPunPjunA5TDIr1lDrrldKU+n6qpbmhzugrT1HVuSoFpdeqA
R9uxEB+BMdcEDvEf4oz+VugT6Pph7ENiFbeybVcqQE+F1sdJD/UlekEryB6TNk80
nRaiy3Y7vve1Z7jDjHMggGCP8IvosgNGmAvl0xvTJnG3/ty+iUsHs3cjitQTLLjf
F12V5xsQz6qxD9FMWGrws98s6Vs4GrtN4bWkm/+cQSWwxVTVYHBBRlyqaSM4fiVJ
4zn2EvtaZBBqE5dOgXsdmTGbUoAH/NnNcYgVHKSbUa+ZWlYz6hnMVNW85txLEu3E
63zdny85llUFLMivEh762gHqxIBTbHh9N4EbggIjx0YaqBJ41BVDmQja2J5S/bQa
hwwwuXQMS9FH0pLeyfYjH9niLToNhZQ+qZyR0aaNJrB9C8i1l5CIlVzoaXi92unB
u3yST5gm76fQuS/ff5H4cNPGt8vJ87oBFKoJNlUHT3SACD7YEthAPT3mkU3YSGjY
8WUqfckY10GOF6Gk7P0SsKNxjeT/a39RcFFaQDA34uUxId6Q9hniqyBwyt1V/Dbm
gOJcippeGhcCaC2weRl7NSJSx7fKt2RdzHYrBum920kXyY4MZkjd47frMV8YVxv6
ZX13sK1DTnZ4Nr/UePUMbW6YxjWKh8pj/0cd0OmgJRrKwy6eT/x/FHDRp1hZpWmy
66pADWVPDrq9usiI3PgG46eeUcKt8zBZNSnXkWS4zsm/XXTL579lEDje1xD7Qd7C
qjJXZIY5nOodhlgQmcE/0XaWOX3nJHiU6PPoLUabxugPK6ur3Ur4hpekkUY2HOUa
9YWpz/RVdQdTUlW2sJuVCY0QAb/8dfSOsisUj8K225oVg/TyFjohbflRMym3okTY
wXKDq/9OXamzWDGudbAsgXOdTd0dRa6LgH/rDSkLlhBi7ZU2xcyWXay61DPJnGy3
mzMqBx6ZTOt3EIQWcMgInD8hzceJ8o/ppBcV6+OVKSmB1iP7De3KEkV7RzOBnTrS
6uyqPJBwxXzLqsCj9V4EZYzCFPVSwDjOg8zssu51bNXQFpgghfPjPXmg7akneCdi
xoleq7xDyRhA71LT8IHUUedjc7i0iX1RSM70oC1V7QQc52KeVNuCOFYdvgFJAHU5
8pT7cxAx+SWWuQKRQe3YGuACBZLhI3ATPd9MaQqHu0TMQThsrllXaXOsKj2KrAXR
ORyFbwJIspSNOEDzokDbMr7iQFN2jM15bJoVTI0kiTQciypZvP0qdo1QPEBxCptV
Ja4gossvFUFbDhSw0MPHz0dyRhcGL5vAlc67/14QmNxBeVJjdS28YNu9zazZhX6y
6FRnMeC1TCyHYUiWZlKJOClLy8mH5HWTjbYzmMqLrcbyheTIln53wKg0wLmspkjP
UkXuBgJrjpIetBgChgWq8E4o/6Sp+Gv0IDqDpEn7SOjLUN4f+N6u29rM+7WDV82S
4e4UUPNI4C9uyFaEcwZ8SqzWYsI5SmWvG/8bBsu51OE72yTaOS3WuSEoq/a5Zw0l
sgcVUGNkqXJPmMW3DCBsgTIUfyemxk4IAHyNy4T3E9n10Ibv+nd9ABCxMUZ41pq/
tvy6r36LAKuRqbR5YeasvvNtR4j/949WAQpPW3WzrHbzLp70V3MxRWvxhRAf4FPW
PxjFaq2Jdcy7vwRxfpQpbzww0G5asSa98UX3z3N/L+el61YEn5JJZ9kwxEXIiZrd
ndYPSGIIsTm4JsPMithhXD7xd/XCytzbCMjs88njnQo+DOfP7VbxhEOowXebLY9Q
ZkTm0E7nFlH7XY8Al0i3Kqr6926rfZRsfqGfjWDKO6VEfz5HI4RkpcJHepMLtyXN
T8Y8IhYMiwMmxM89yPx1g/QuNXZUmW79v4WPJ4Yu1gnfr+w0i9pqNrd2ALSG/0ym
qvl2SQlUrATWSn8bvhSA80kKFSv9ES/+EyJCDiHPVf14s4Ae7xHlauiQi4AJz2Tl
nuKPGBvpXiBe7DSg3gFY0Rl+SBok9O/k6ejVLOpdJCEQP/2HQ1zOa+rezg6Uh3YS
jnEhED0QoguQ/ZhxvgeAx1NQnSeMBiYvSDsYR6wHv7rs88O4JME2IFykMRWcadcS
b86CXPCoZzgH2iPJRPDQaw2g5zoZmoI+tRduJvFAQpcKnJX2TUE+1jmvn60l9Mvo
zc2Um4U2kbx94txXfdbmEOxrwJdWTbi/b6ePPWCPDvj4qpj3SewnFUWOo0qbIUbt
vOwaObTlscPJGKo778NMs/LIGamjk3ezvTp0B8TJbguzwdHXURUZpBT5++FrA82N
Zt9RK5YJ8uUhSQsucbWOifQvSxAA21jcr2Ft8/LPC7yB4dTVpMzgZFfjzJXLvUxm
nHgXNENm1NeY0xbey7En36msDf6cJkKaiYMDDeIylxQ8K4jbmqQIgHCxUx3HoCCD
6p/c+9YW+sxyNYmbGaOVBIq8CNFH2WiBCp0xx0Q1wP740Ud6NG30sEguxqjYI73n
Pm0EX0WdR8iS8S5dJjLY7NZi28bTQiNnkqhwsZMl3YcsGPHvW9xPSStdGMMnAtvj
pL5DWz8LEEdooYdg7Z1mm09g0QlfkuwdSld2JtfrONbTbPpC2v6JiouChRQ/U5Ae
JBnuWRhHkAHB/DO/sI30UwNnl/Rn3vg1x1NjtoBU6yb9kfxBS/y/zbBQOm8i5agb
o1h/kW9QnpYXEivKbmtUPfnkLzXX3af8oBWcJGAMjY4EOWGjtVVtfVIjoU79ugX6
TnlSaGOdPSm5zJQpvvozZ1gc3+R9GN6uMclE4nmJTYzwcXSnJOxce9i4oOSVZixw
P1+BUKkhvAcG4WbPGZhzrjZRXEqNoJjKrCSi4U73ZBq2Wpbri5lA/mipxE77jisV
N2J5yOh2CN+m+RRqUKvvKECek1W2GXzkNMatpe82rKcgDW4Ru0ZWBJk1Be/pFo6/
U5VEWE0goLJdhIDM4ifCQhO1w/FGIh3lq6UHYWNr587gb87c1cKv2wlO/3Bhq9O5
O0A5lzk3lNf+6Wlr5cI9laKoO9hPNItDlGi1w/ei/LsqIYD/U/foLu+Zr52PZD1v
wLA0fBqLPkODEUvgQ7rxXkPC/P4p/huUrP55WTpG18Pr7dA2i2K2DfH5O4JfY+cW
OqIW3VEwnYylBGQhMokLmoQaaK2rxHoDByOJVIhMHkqIpgN9wonH8Ike1uspX1XW
vvc714eaMTOUiBVZaJ33Z+27vq/wyhLqbF5XnXR995K1Tbb+lWDUnHMHX2J6GkGP
iez/egx0VbPiQnP5O7zE80A9px2Ypbx4Mj87wmuNN3g86jrCkLIauPxJjKqJlyvm
L2RoOmvtWaxoxt3PRLe61O+XfjPZbeBFXajkR0zRVUwnjXcr4msANl5JwHmY6fdo
bXZZusi6yNlP9S08hZaOOnH82qwQkKBw+GqC5Gk51jzH1SdoKWO2i0vrvqNsNjBt
Ijt9oEzGuGtS1THR636jYXBsJ/sLcGqO+SDDfF3PwZ556pgMB5UbOfjfyGx7CZHf
Af/q/RkW4ov/wnCC34L80Fl48bXcYVf42JZQOKcMBjWxyPgur2aZ0BaJhwwPpH9N
+MQRorVWbOUffBpRm8XxrQK8fwNLktVkVn2UViv7ezMPDTbkR1ZS041VZwe8JFXH
OR9XLUte/dYhVELvbx31Rp15kRKoIqgp2kZw123zss7SUiXkiBuTrA+m5QMXAF4F
PQTF7YlowPKsBsTzLEeEaGp5/6YGj+uBjOD1OFEDjXoVtruAfek6OgotynV2n602
gAbPwlZbu55qrRgHrEMYE3DjcfeEHGAaCxIhReudq/TWeHyLnhftbxJQgVuTlb1Q
MYyjfDrOno6ca5QVPdmrcwPSirSXI30zBFg4nOwLFlCs7jEwN4NEphNmaTB+hNhp
3AqXaAKrygCwHGJAf8SdvNN6eS0wA3uGn8Q/5dASFyKb+0cL6dGBiLRiumLBmMCD
T6ALhC6ihMfPOvRMDEPY4AKzLAePCcNBlx2yjXdQTViEr9DJrQ5V4Kdv8mAj4T7P
y8Pd2GT5XxrCR5y7Mn7D3WIMBZL7zmsrAC9sLu5dA7sxBjJcT6PT7/sTfM7Kg3sV
ifJgWW7qssRlHOscUVeLVMq+4qE2qnNliCIKrF1C9qaB69vEazHQBA1uFfsL4mmH
uxQFdlTC7rW350lMRIiLfdmAq7dzPvA7lAGM/Z/4TxaQJnrd3kvKnq+lgjA11Wg3
E+UUKp0uLVWBI6UCd3E/S5vMaNx3JUoitizIf3l336r66oUchFQM9FdT8LpEKGan
K7PKE8pAN4M10O8nHZhowfYUPmeEXIsNmNi+IB+1dlijw/lnYk07QRl9d1L7H66c
iV/1nMEdPgnRE0BH3/9gvuDx2gOOTZdd3zcqbygAUfYegpwEFV26T6s4IkOIm8NG
V6WSVuaP8c+wS4MtliPY5RTwc2CT9p+VlLkToj9n/aKzyCPJheo1AYWlx6AkewS5
AR4e9KaT2yVNpWvd5WoNrQpaNjDfYNgVhEnhZmqrcmvSO0kvOk+l+HFK9q5xg1+i
mCJIK1CdNPnhF04jULz2WeLIoU8awOAzZDGtzCuKuw6vG9C2GX6gIfQVAoVOiQWO
oVJYhGLglF1/lg7v8zsLe+pjFjvtvPAJS58k+jGTlSzgBbZTzcdC12KQfbkdZZOu
6vmq37xjJn8DwheQjAIAreq0Ct0XVX14ofcIljLNS1J+xP04F6jNiUq3ZQon/1f2
7kGUO3FyXxA9s3E9kW2y9w==
`protect END_PROTECTED
