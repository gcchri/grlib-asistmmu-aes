`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJSAHQDzhfWef+R9WdOXZo/AEi5bErF/VRMvKzAvuXP+wDyqM79bDnauwri82r2g
flfIaeQB3fyFetrk60fsM3eKaWf9LffV6WA3JzizTTyzDqmX+jXffnHbtFmAwXx8
Pjk9oUoMj+KzECUTx/01hdJ4olIj8sD/b+dwXI+tEfjUJfD6O3QI55vkyKUBlTHT
/j0C+aVanSNfCh4IDPbkzQQ18Od+Dm1pV1r/f912O9hfYJOaQt5pbUhTXVH2tqoa
hFCzjNqU+kTQ/FOjzIL0GSZKr2VpsEYoxvwb10Q7zWrobnZo3vJXIYg4ORlzEi+J
9m6wHIxAIx/j9OYPwrRYuT0ub6RMdu4cHjkVb5Q2xEggdWuide/wMrYy1qkt9fbJ
q2TmIQirnwbF/h9mjuKvSTs7K/vtJrF8OSF8HbEM1R0rNxQ/1dF7mdGf66K0DnTO
6ftPziN57qkfyszK1oHO9WH3P+PW1QpR3Nb38wPn6Q2+XgajLe0DUD8md0WPqO6i
iRGKfIbT8kfkwEUqsy2iTcIoFWLBHki4RRWgBvMXWxbWwLWzGNuaV8Xv95lVN2VV
TRCKu2WcOWISorVClDVjIr+PoHjsWfdWdEiYDawYHNiKqhIamRSrdsxHnpasDVB7
7kdEy24/TIrzsckw8qVAGA==
`protect END_PROTECTED
