`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/3rKYtn/ieA40jCUEPhof7Hj52DW+xiQpYDDoAScyWYmfkhjkI3g1LP75V/hil9
NdOK8lq79aNX1monXns/sU+BJf1SoM0aSVCL+RTwwFTgv5dDrm8hTULwvR7PfrKw
b79O7YNRvzY9u+uqgbmD9b+KQR0sU8jXSi/a4R9OKAR7rgSZCe9J/oQsMK7i2gTF
jSljO4tCJRIMRKb+pUv6MeNlumGFO+cU2YtKqrZegzzklzcWfLcyqLvgu47ejOMW
CqoUc36NV1aVjGO/ghUux8jjLg45ptxKhSi27OZsfnseaCFzb5+wtETQzstqRsHG
nIJcwuFUMPBpDJpC9sDeK/C+GyJ2qM5VCQlFkRdo0oAzxSS5yC7bmeTEfDrvYt8c
jm8dQ+BwpptV/gWnf7b4nEGtvdgUUHq83VSaPI30UZ4=
`protect END_PROTECTED
