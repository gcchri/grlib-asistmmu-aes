`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ebn9KTmmi2tX1/ZFJKMr/FMGMn/ww3yQ1MComAM7PKhQRpQmrhpicXSq/C/pF7G
UolzyWGM+Y1sMuLgtUBtO6DoLmBH4O3im/W+zQtie56QxxGVG+AwaZBY6jSRkdyk
wGbP2Ev+vVUu9I/BdqakIqplwwdxzOR93erIPsFwWVk4B27trKTpoLC791ukxtF9
DzOJ6BAhxjAumXW+Y3J8IFonOHwtna2KAPL927aX7+JRDk5rVq5vyqlhG8nFF8Je
iysn8oH6z4K7+6pcq+cdKhu2PEeG/x2wEr5HOG6T2Eq+zDH7W1nLLLjsDfx/vb6j
8BYW+xo5x/xUrRedcz6ax5I5mfzNrc6oROXliidm/B6inzlC5Y3LwG9dPOZh+v1M
czoua6wqkezF1pkP97gPyA==
`protect END_PROTECTED
