`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NRlQNsyNWdN3MZAJ5TUyZH1WlZMCB7MAAqEZmWG2cHeEQ0nCaR6z/+wE/4ELTjj
ID+2M0XkE6/ayQ9Hq3WG61/6TapJp6XWIJlrOCuQVoI3qlXFmDr1WoJWzXhmVIuy
bHhlXKTXBARm42mG7ZxRLqvF3dMV8RzA4YsbwRyOtD7kIn9qRWmELOjdoFl2Tmre
3wQX828+pURqWdtmnQmz6YjrFNjPYOSpa+sKX7N3c1dDt2rhLhMZ79U3Hsj2w9wy
L1jX3c8gEun11NyHkcVWDTeD0XMP7eIch19J3bUU0n6jav/RWubDJ1VachVMZAyX
UaMMQEdp3nZ3c2+o2vH/UyzHX79wzTrvAFgypMmatv0EBIJvTE1KzYTcMSzuTQXq
1dX302ZHxj6jUFz/qAxU8+R3JjlWIloVdwIh9VIHR1s=
`protect END_PROTECTED
