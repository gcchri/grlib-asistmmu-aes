`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9IpWpXJjxSgLBpUnuGeluWVd6RcoXb2B7G3H3Hmsrjm2gAHdVgWoxyEfHOKizP9
UhYXyrs2bBpE09ctO/sjiqXtl2ZSfpPAn8B2FyBvf0kzMjR+WpDHkY2wtcCqq3LC
oW2KBg1zgvX3dVVAoaL+OxzXRBzJsUEo1GtjOh6PfNSE2OA2aFISmFN/NMjjsIjM
DbPiw3chqy9sQ2EoOtGBjGoyl+jCNoooZm10Z+L3I9Bt02QI9gbg6i26gylgfL3Z
Yed3qR+1sfcGbfFHm1iTW+eMVeMySJesIkvNpnGQuIanFdhbHFIeWKhxYDWEas0L
JVGuazIDqhLZ63/vPZY8uY0il/XX9EttHhI/Ro+8my1KcmMXiKCh7DJEqUnvA62k
hFbbnIGPhYctADVyJLxrBpl6oRosY/SDfMgVDSLmoRA=
`protect END_PROTECTED
