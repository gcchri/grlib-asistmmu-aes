`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GYbePfdD7FVB2Icd58TYjVT1QvqgY1+oYGiBfQeucRd9o0dfJybAWImKDtYF5afe
+kqVRsqABPTOOKBSA7JDzykjik7ezO4WEfsb/WSLssVlfypye/FiH2jV8qIIB1I0
gU76ixZD/2DRpfzEYZFMs2o8lqa7jwDqcmhVYEwNsK/LrwMS4QUl1P7sZCRR/2pw
p0fQbC+XSwmttrn0Sg+vjm50uE2JjOnPCvAhQj9+n5K9c07gNd3jhvQe4y0jzKHd
qpeN4pWheeizeSBRjEqL56OCKmrXBcZA9JwCJzybU+AC6wu9vlaH6cLu8P7i85Jg
ZJJMKovxLbHpahQP4ju8UVB+3wthxJOIEJ+Q3cxjFOmWx/6ZRAhGt2p/coLtuPNC
xXpvXugjVsyJUucpPReauwIyyWlYMjWSlkT1DOY1a4zmp73phKeT0DXbfY+t8igG
AC+BWWUDIPsJr+cbqgZf84DxT0eZu0kutprRIssh59cjCtNKNVPHysD6ixG+McxN
5OJJq6rw+VMOQ7HDYhqx83Ch3jac9moKxrOVX3DH4LqnGdWU/kxrd75yZYiSdgSx
CrZ0NYOXv8SI3RDKkcSkmdr00zblUIEcjhnmv/NpFPRkpGsXb2aXTgkNf5iw2c6T
PknSzRKhSEdfRkj6XqXuVD02ryyQE/1KacCHQew3LMxBHGXrJ2gVVZQgaBIjuzSe
9TPQnN2JimEfRRuQReuE52ylNkfsWxw5lSkDgz3JoTtvAIu9kqJaWQcLgQXjJysd
8GXd4KHLt5KtuURd7Y5Xai7QQVdwveMwd3uVYvMJ8f5TtHsS+kIKYFsNmHR7UT5I
EfPSo01Dra/XDB8Kg/R0mRrAeMQT8m0/l1d/9l8Ve5cJh9d5zRPU2pUpeMIlgD+Q
sxigeSdrVzPRkIIW0TrYfXIbO6wX0o7aPDiWOZtDBrIHLVaGLYq54pX9O5I0lRt1
MS5mHxjegvAsNXXQ7JWsbBhZRHW1T5fICrov7aHIMKzR/A9XPk2lUcyiIyQMfX9t
XZ4ZUQhVwKri7w3DgdHeM9fcbwlARGc6NuXC6wYkKX5w1Uho1l/GLty55vYgXvDW
etHCrpx6eGD/SRlqou3XAxSk8iHjtEMt3h/6CB559SAZ2fESa2E/MnzoxORPv0cn
bLTZPcsTq/TLV1jNGdnATp4U0XBCjXXkGsav7r/VBKkZi47konieDTjMJlct1hTf
OnG/8M1ihfjWftdBtO8KaBXINv2GL+pBybqdSV11xX3oWW9AVPyLVxB3SxKb1IGp
thti9rj5qQ6QSseoPRD+/VWOha9CfIug+8qUI16jXa1ndTPqrTgAGIqDynczKuTs
gDh9QM9R2/n9NuDIGcu5pEYUbNvqlUG8KQTWlK6kTeZ6y7iOtwzwq4sUpETHp+Wg
FeB2noOb8+mSTCLaQzKS0g==
`protect END_PROTECTED
