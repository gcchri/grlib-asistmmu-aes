`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f9uB9qRGWGP/hA6XC9gvIIdv2bb5pyYkVH7YTOUyVUa2ePHgKKO4E/2iXw6cbRpV
E6KRMwoJBAxAmNCy9daf01W0Ncbk7AQK4LE6csoo+7Tp4xMX9NjSGm+kmtsp6+vL
/iXeIahs5fQhtAuAkfJjnsrziTQNDxpzE6Z4VQtdH1ckSEi/cl/MYk4Grh7Fcn8+
FEBAVTt45RNBuh6Wmf8/3pbJJA2q0t1LEFGyMAm9oWhbx+qVJqnlEZG0ACVxOwaz
pFcl9A/HM1fZoAmpy72lmqeV7ofIzrCMfUX7bAzY8ectg/ycZHWnZJuIvYeqHCc5
2/5FImmUGrylWsHePfq1D81XRTTHAUfdJb0z5rch/VEgp4JHm0Nh0apSCjiGGnzs
yFWlVxnnGBhO4vqs9tQo10GXkTAcdbKn6Pp1jve3YPvicPT5c5ha2NIersKaQ9nZ
`protect END_PROTECTED
