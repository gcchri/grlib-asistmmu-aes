`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3RO8y6WD+jxw5fOx6XFbFYCcVwN+BBJxLn17SFnRAdu83aINeWdT13b0gwqPMtK
S9F94doPX8U7FlLzjoNwbCI5+akiKpmw1VEs4UAgPROIrzReKuDEGUpQLjVfWuUe
JP+ZvtEIh4AQp1m9ipyTsqUzuov/dKk0jNdwag4bx96PIrK9wRyUFeVPfNCeDs6+
j8ESR0Mqlen6YanfTn1ueuyUzsrsOMob5WpiiMx0fppvLbNECy+x5s1GvNhzEfBt
0l9XL4HnpfNZc5dx1K5a51FydBbTI5kVmukY/jcKGFR+jpl4Wk7SrRcmZZPUkqvA
eNbq+sDmoYQaY9sLfF7woycbKPfbjhIFPiakl+Qn7MbkLzgG4em+uIfNtHSoZfbm
XhTmZ6BFI383ZXHT8Lh2u6bSq1QMGzmLn2gNI7hW0PujFniryCJ4vkuQJsnaLWF3
wbtRXVOUJeYUIZo7oas4BH64/KTc1sEc+2kIrsAdEGcDOi9X9b1mvt9ee/9T/OOy
shWYfvrtkssbb1LGeEV6cNvDbGsLjjZQ/Qr+pTyFPBiyQYmT0LvgsbADgrCqWrPJ
WmoPg913HuAMh7ofx2FE24o0jrP/++JbSRjx+OUSQaenyU6yjqODtbVpeFgFx20Y
EDq2K9mSgyB2Ijgno+RV4AaB3Cv19FZyna3VWogN+A3k0ZfU5Sp+1Hc27z/07xSc
bL6Oyr+q/oQl8vIe1IY+IIx8DoBem0HfshlDP0OC0FwPqoSsEaGz9ednvv80HF+B
OrfC+Y7KxH8oA9kYN0nv/iC/EMaX4SYFxwdVpz4aSFPKQiKFVTyV0/I5ndSC5de5
l2WQT4cLK0hsX0B0W//LahdFlSz4HFq6OlR0OinyKAFv4NJXeIZVu5ytIpDloDz0
sHdDxDz/QUlPeOtXIWyi4T3R2c9Tugasx9Nu6HMZQh5V2wjCQ2hoOv0BPV2xOTwq
`protect END_PROTECTED
