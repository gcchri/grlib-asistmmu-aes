`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tryc1PgKQEjn6lNnK1j3yEWkb/GrB8ezleUB7TG9V2Pu17xLX8dT3mm4SiAxvosE
xI9e35y5otzeERE0FLHYFqdIN9hAKHRCuXZbdtX112WTPABF3+x9XkjITW3bU1s5
Kh67Qs8rvVu6JNBSQIDYQF/iy6EGH0/ptbIWUgMzwAHLbl+rMHxbFJo+vSVKpzcr
TNkdLqnU9kE/7KbfJrBVmnHsdvabX1LRBVv1O8NUOhW+0jWtqEaL2v8zdraVyhfH
/SqooCj8+FEipNh+F6fkpc0851PofSyLrgsjTdYaGSkExZFkJNcNWCMqR9JBxhzv
PEBHlKpQWf11DLHDMhU3KKGn+vYaIe9TrhCQdfhIqgZgkfk1bWoceAHGT1PXG3ot
43GlZSbKEu6ewB6qeE87GVtaZ3+iVSIi4lfzjvWLaVQ=
`protect END_PROTECTED
