`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wyf0Gr+7U7ms2h6olNTMZEUr7fgErw00kAlaFJWp4pjhXkzGDw6RZRDiI9443Ki
IjXnP0tIvfEZWZO1G+t7RNCluUHxAuHXwFxCaDFkgZS1vu7yZZiT1cSeZQglG9mj
cd8zLJSz7crdbtJteY7ikMI/LD7USY87xooLNYpXNeFC4ZaP6dpZgPIJ3QDWdpik
yj4B36Jz07o0sGTA+mnM1ceYuuPcIaKc2MHMk11UYYj2vp8bx4w/ttz4UcAoAJnm
Nw/Ll3Z0v+9xjz/MmFJWGGJJiZRB5nfLkkxRZ2/QF2AkY/9lKyuQNCTT/k97s8zJ
JF2Yy1iXOqEPec2u3tG/ZQwhYuAoCg4fbU5Byb1t/u6ODhNv08qHzT6ImswtQQCB
7HsNW/8O8F9nPKOyBk120OnKdz/bZI0YH8UacJeY+yIWLNvr0TYawOBa6/djTs9+
3FNMNwfUlsKLTS4kqZ+ySUdJxqUCrv73GuLI8R3y+tvWBjMLNpvL6IlHErTyLMU+
gplrzvB4N7SvdEpc4+HYpVQVImT4B9DIF9tm9VYh11tHq5neXtI5DDuyhGLYCKh2
ZCrZZTqDkz74pN+mvwA9LJe08lvmVE3aSBW1Y3VRgK3oR2jZuIsnbLXljX/5ZD5I
mNyeVYuRvzF2PX8GhtpDwsajjVjIRjw0LoXGRWD9gb4nbkYkq5Xb/jIb9p02+eP8
REhqToJZI41PiY0hHSK+Y28JPs1evKAAlVU2+x0vRapWE2BUw4MNf3e0BmyuoJGX
w+m+BXDJXrj5rWOhRwlHvEwUfyyYb7QHcd7WbKGFubF5YGS2By2jS16jb/qz+5qn
Pq84060rbLrClQPJUbNZPgSC60PWScEBJIoo5tkkHXMXrifx7aA3JUvyoPowhhs2
ypCA5VK4iI8J5zNBfYABfY9oBzcoWauF++AMMZ8vF1cOTuf3Jpi3NKF/5+nvDYHc
K9wR386O0Z0c0HNTRr7YkqwKBFbEwO4pM1wUv2bkswL48WGbj2VePOzPB4p0BEQZ
LdP73bWr+8/VYxxOFWtlv99/pbdl8QF/b+7MpTCuRBo0dWfMp8qN0nUApP6hU3R0
Sq3JxgOXggLGJa5WPVz1Lp8YlhZRLRWkgtLzhDr0EGaXnHPPvYtopdqN786keEP1
DgVrwCd++eJ3uY2EAIRczm7cSmyY8g4sP7kklyWRMe/4Qkgbjm8hnaE8vajnZOxk
iqwi89y43nQ+VavPgpTdLyWYYSURsGs56HDfu6NdyZ/kR6QFfDerUb56gPyklhbs
P1wvVQgPLKAD/zmw9G9NSLIisZvWPZl29Sw8CK+hQi8qm0NqNko7GU63D16Pxr9O
yDydk5AExgJJw9uw+0YgMHtbuvrkxsfytCR9AxU2vLjJzm/Lw0bbVFJkc9a739A7
FiH6yk5gQf1KZ3Gu+p7ACnptZkEyzvIURvPwVzpqU4JKLUULzABnjoARurwCTZnt
O9d+NghMUp9Ai6SGV8KVv4AJSWKxkCaTthS+wE4JAP9S5BI67rRrGX/UTzXhhKwu
V/RRFd8qt/CW36pF069dZ2E7H9v3ndXOEX0pb1SoOgFDegP+ylYqzv/++7zcvnZn
mglOAvw/SGtYDpLXLK1i04QEpFWdP655BfqS/JkBjcptqUtQoL2ApgnPKgFhlt2f
yVq4GnG8RepzgzJhWkzwy+QOsESK7oxAciAoUAguBiIFYer2dnxs7CJRAj10HBd0
cMklHGFAqYKi1M/nvP3JxuIxeXcCpg4rwoGuyl3zMFH4+vs7N+F6ZE/3fVBghoj7
1Lzt28XUGzdJwFA2mgT51dRrg1rHdYNEJU7NgGLCxcBieslq52nwDSFby2X5C7LI
wKrUcwR7WtdMU6v5PEFmg2oeDwgTWnU+W6Q+oDSElez9nAAfdNhpDmPAA9KOlkM7
j+ro0S4ayOVbnl+I2kuPcPtgHCsmAIVI6lJqKFRxr50201LNvPR8zfRvf4xmKMtL
fZ/QTc7RnqSiRnGLIbvswg5stHowCQfp8Tzq79EeKWE8IWWDZar23EZzuSjlzSnn
rljfrrx4v2E9EAceMzamAKmvDtqcMd2z+2qqHDRf7T2MOEhVkQ0lZPc3F8nduTI9
4rtqCP0fU60y63im5gGZ0LDJ3jII2YO5CZxdlgSAt5Pv796sqjCBPKdiOqNQxagj
M7Ty+HWrBjb68qmwc1pktn6pT7994EadedXLZZFHbSuuDfnMw9/R2GrPgPxQ40+/
MjmJoGvzjfrRanVFQ8mR2y4DbjOph1gUO4UT9DkBETTOWs3xrQAqAfoICHP7SpBl
8i+Cmhw5h6zhX28tTwVQ79rPLhuHyn6Of1lS03Ks1dPRXbPgedLM41aKU25U8gE5
D577hQ2xJ1IqylDlVG64nuR3RmLqPjycuRisIhWuQLEXPSWbU2BapNh0gDdHuPTA
WoCRY8cNYlg8tWy2BQeS27ZryNdvy/o4EsCspATC9IignrrRUqVd43Nz88bMswLQ
Yx5X/FGha03QBFZpLO/KkYMEXjZiYXIcpijWntHh/lDQWl3IruHG3A+PrDE94n0R
Ctcp8stSsgq7iDk121GUD8XLIfCHXBal9tpiW95opPwfemEPlASxpdO3DmW9X+pa
Cqw9d4liGKymy9i42RaLx/UEw46+im+aHpsh/fpiNriiMHF0zXZdrF8+8DA1fX7m
V6hgbPUOkdv1nJGvw2GgEEpyeG3s7C8ZUfZCDiqjVTAvn1jhE/0UEchDJ16J0+wP
0/pgEsUxQPRraalivbY39omwzcypt2lqP1R1otvqQ0Bnvz8iYeCAnyBsBt9HEEZm
kxvTLwi4qBl3tfC1PrT6DwCulpPRngDT9aq5zBbox924+PnsTAfGObhi+cdKc1EZ
9lUFE8SRw7IFA1YS3iH5gDsQJoAO8wwY6nUY3LpSufITHzDW/+9EMesSJTGTwfZq
1KKoOY/kW0uW8wGFgccdmz6EtzAUM2bdcHNqMAUu35+bWU+JP0+3672CILzvBqqr
uklxAdjxyS9nwGtg2nni6qTg4Q9eCX3F8TuxsAVJ7vHn5TphZz6XpIC4tnuQEzxk
NF7zhZ7PFvmMsQV87XI9ma2Vq8yyTi4SndymcmZAJL0YV/NJ3qPuN2DyaQwjfvg8
DyTlG3naQVYpncSe29JXsrBPgu+P8n/nW/TqHzsRT8avOeT4zj/Z9AxtfSPHyrnm
mDPP3QfiykrF3x0sG8ghRE5uEhohuz1y/RBxdXsJgGy2avPsUHuNv/6Z5hub6g5u
QHcDKKp6ayIBJbWxQswoYQY30X/mTM6DZNUjhRK1mHx0AUY7WECYbukkX95uytV4
WtcxG2ciKTZEwd2fzMc45g==
`protect END_PROTECTED
