`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzZ54Qa61J0mspx12BwSXAK4Te1dvmewGs1WlxymHVpSjU3sxdWBJrur6XOXL1q0
tXr9erSXJyT+1jZjzHqnXdqC6ldYLM3jtUS+ABXnzBn/gsHLFr4x/bhRtspDGFdc
6Rm5m2BkT1a1bCNLyyl/YaDDfv1KzlQj6wT2paaCdurx5a52RPCQJi5jFy1vpHvs
SzsOE6dbY31n26zIWZALtDVVNu4hCAD1utaWi86ohHzkSgNK+j7koo0q6QQnVbud
8pjqtZh5el8QeLH4oav/MBw2RYuIKnyFCDHDGfZCtOVkO3k6Mu4TY9gVzqeEct8P
lgxx8FW2d61rbtQA/oS22ApBtw5FjQrLb7Kq+oX9UfYAO+WbUOf7UpBTKeUDFIOB
LaRb5U6ZLIOP80s9Mg0J51HiE1RVc2532SCUfJIw65tSsZVRNJ5HM8fn+24y0VAb
n1kSmYfsbSebGzEpanalVK+KgGiOAQoSy+za1PYZbTlZqa94K2rY+iephTO/CIL8
5C24HvdGexvc/cAyXhonwpZljmmTjHJAB5nyrtTryNKlr/a1IGhMncLZC+CID2dD
rYSZZnSd2101AFnk/Ui4HtuNSN/dWHI6q3ZuCqTA3dEljrVWUV8NKGhEFm5uFOqT
EFlIlxH+Bziu5p1ThO0mboKyoUG2whdYVr9m5fWm+91tw/PW2Ecm/VRqSPUHiHyd
yfwZtGEA8kex+azmnIsdnnjlhKAtOq8Dyl6/+iIIYEaGiNhFjRil01fMagNRuvnV
HHyGtuRQlFF1Y5AHC10xxHBjktkLUkLmzR0RSOsD/gTDGSmFbio+jj2+Z8vT96jY
E0ZOfixHDmWmTiHJVYYQXSDrrG2gktsjcC4dgGGkvAfyH1ZEHIw4tSyL/ng0eyh5
JvX1EgkaxQYgIoM/kODNBNwjwUkpDfmXQ3X4qOEzwY+pqp4sYNOgNKfp+BViTgPX
ffflUIVMXBLSReA043L9jtCl+Rd9yy46re+MXLSxO+2XpGKyaJKW0R+bKlAIbkQF
aepEPs/l3k3mQnQPx0Fp0SaEYw5Is4e0N5t4yG6K2e82iWVHh93G/A2KsAlNuZ0w
3HnRl8XNFKLvhuMnVkCdt9Z1J7Xbre4H+tlTguHbEbACwvlwlO6WvOvDfGuoe6bp
fgBdS2exhHwzDQCTn/0N3AWvvHWjQICeFN7Ot4LNnyfZTJSj/LL1jOnLLedTj1tH
PYGuKrbzeDvqhrdmaCYt5fW/98KD7LATZDGD/ZGGyuDzQy7qd66LtpqkEXzpaCYB
S2NfvgTto0vQ5LbOjYKbRoPUYIBQOZXA5a8/NojclnqXdMqpvVxXRegfNWwfyM6f
zRq3DZLAdjxvBNYfXv9fGdxihx7W7YlnmsSgnsmZYiHfdBTz+n978nLyUvL8Mz/t
p8jSwpgmI0vHgKQY8KvgWDxd0XG1dd7CSn7JagcQ4u6miyOFiPxgvMK0qtXhg3AG
kUCEIzfFx0pPiI8F2WTG4laiGQoiBOWdVrE+OEVqoZorpfmkqaR7qYFqBuF2bjkX
EK+B9Z2M09kCOhna267/sCoy/5DTXH9ZlyjeAANEQXyjO3IC8c9wrU5svLVUsnGf
H0H+Us4wMXwNIPShavaUQqirhgXL1OCa3rCH0Fs6hwGMkGTSXbMmkKWMwJcGnptI
pbvkiTbQrWOoqbJE3qUckH3+/KjtI0S9Xqb2KKd57zEjc+qnggxkMJdE4coZ+2ub
YfoC268TUJgY/FfSHBs/JqUL2hM2OAg+kn1tIH5MEVDjyOZo0xHCP5i4Qgzulxk4
6yWrsm8H6iR8qVnwf492SBMl+nYGQEXYwtCBpvx5bbNpLzujWkuD81xpp9F2g2ZF
aF+v9TFDe6DvWfW/7kEsZaa3f45/1juo1t9S80LeL0gBagDB/MYms79nZzdiySjC
EoNnQsM59IdGJCxa2pX/JzHLVeo0ikZO+9NaXAgOknXghQcjwA2NMPWhuA3BE+ZK
BQxjpUvNvajTF9p08tpZaCkZAjwLzZ/7s/nhZ7kWSsje1PYvc2i+les8W6vPiu24
j6O3jPP+967XMLbhs5YB/ID7Bb88Saj3KOGJxgi8l2/bstgDDpWqH2ccy76sLzqE
zRreOwKmh7pnvUbJ105FCVhXJhQIwmh8Rpfvy7vAALBJyCUzxml386cYKPgB+zFu
QfWWVrh4rpG+bw2qf5LwiU+Wbd3iTpdzRaqTgV6OLDyLmas/Uwd17uZ/YQUSwH1G
vCjFQ7MZp5/0h8572xzlt6ByV/lIT+FuNL3ZGVeTEEt3+YtR+LBwJi+57F0RhsYu
ZQR8T738nUCyLtVebU4Q9eVIZSJK+lLE11VR2dZj5AJSvYtDVPjhpprZq6sVsTpO
RYoA0GXLAPWEsulq3L34VUzpNfNc/U0BG5C3psJR0MHZCblVD+a2BGPZp0CHynAA
jVJ9nHPZQ5i/VR84RDrmLsZ6ANczD+SEFVLQRTVVNRwaWmxD3H+GtykuzswCiNEj
lheNDlUENt6A6nzZFsUg4dx6aQmCCLDL6szGOrHNfMgn4xV6SP7xbptCAMqq/Mnm
kOWXjLvzs9CwZf3AGdMTdPQ83F/egFTuAOJQZP/qw4gUPH3wGktSyUIRDxW8P/4z
ylrE3ZbLbJmpAF48lYcIq2fAk8wCMsYsx8tZwQ1e3u+m+cjMbBMFJPUoW5cRXbPm
tS24HT1FB/oTazGhcgoF1Vnj0rbOMdjIeZfqf5EzzQgNwFskqcn79rCO1LQKTDUR
zQytRDWlETNm6GY2cCHIiIoBk8hQTjpqck5FzxyNgnycul7XUvubPZSDK+kGItgb
xO87wnmx3mbT0XHZLKDMsvnpa7vE1UTvA6773ErUku9fmMKwP6zcvzvGLCgBQHoP
peateUjvokbFZ2hv1CITgLuzOTZbP95F5x9GLXjugFj/GyvPHulOCYHvnyGW1q7r
QmICxDs7egdCkmppAY7p1t8hwjr7cZuPWTWyCeRFO+TdGSzseUvuMo8lsoGGVDTu
VOOQlHxPs1CZNjp63rNShrE7PANRbqPi0ApVg5MDEUbwO5jcDIOhDcRfzIUMGnaB
sfKMSZrWndPM9O2CecmDL2iVVt/rCAJaRLjle/Sazdw=
`protect END_PROTECTED
