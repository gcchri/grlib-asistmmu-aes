`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxgiJsI3qBfkwUZg44LBE3FJp+GE1yHGEWRgNxKElOWjpwv86Q6JdoC8ZfRZXy/x
ihDLyh3IShdtSJzWUPgtf0YnbDZ1s9wjiLCYixkRjmLb5c2ybSV3kRK2HIymjB3o
J8DCUMbRBp5uH9jvXn5dPUrLeTMQnyKugjlz8tGwK7IosQrrAxBAyDQ4ua8KaEGd
JgGTABsdmlhn3UA89rFZyFmaRfhwt5877NUDdbdXAO1q2f5e4cCcZz4/Gm+AL49M
E1EFT7N1wf1AKWQrA/EzS6lQt1AL0oNR8rWxgXMOhZvfFepuBmLXyVHrl8bI/bPO
RD9X1BisPVbPObVDZS0YJg==
`protect END_PROTECTED
