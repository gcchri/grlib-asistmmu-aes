`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yRKH+gefXsi6CUUA64nhdk1R16nElY1M4PCEbs3iA/c3eWiPFk3XpgEAxxWbUB8+
fLPu0HkFyC6PiQ/qbpCwULGGMdtQ5mXgNnZ+dMUw80R25nB21/vYUcFkxZwLxrRv
xzeHtNxkQqpJfGdLahh1kFEikj2L2Dm0n5gQUJkifCxW/PAv8e/8L/OQnCDoHqKL
+hd2lFVREPQDeIFq6y020fVCCkbAQCr4iw/sbEMOBJUAgE6Ld7abd7OarW/NMQqu
WAhkdq5IifRTq8WoTBAZXFtPuGw5VncOXp1GffoB2gqJDoiG1gDqgLyGYmY+6OyC
xcdyyuywCX/ZPvfYVESEsgGNcNIayOA+JqFEU81oxZiXeCrwcSdgLj1JSLcBrytL
2LZLcC5qktCq9Z3erRJz6CALWOxmAPeLBO50dKblwwIH7YEIjyCBKocZe/X9+n9u
0OZfErLbyeeooOkHp2bByEB6PFEhQDW8UMKuQqE3/AWOpkcBNhY63CTEBgvzIPQw
8HE8KGq4l21dx9EvKWb6VdYhrTSl5cWuJmfKnUWk4I2vk95DVCBI7bVd8sQ6LhVv
zLPO4nuaAQGxUr4uUK4E6BJNgl6x+LAxSnr1vRYVQvNHi0BF4Fj5T4g43mow2PDe
dCgfLgxCL1fGXOYoL5zJo2sMB7LOqmOFcng0p5usEkNI3V2T5k/aBiXrh4FbHiVR
BtBwYG8QvF2wO9Slme21Vg==
`protect END_PROTECTED
