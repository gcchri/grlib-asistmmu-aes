`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjxgMeX+iQ8PAMeedmMklSS7zhL+LlHGozUA4EC+Aci5ONl3l7kdWxclrhp+QNbw
1JewKJ/EVqJScfHi4A+7/ZnsFPMBimK/cVUjH+WVPuhkAVyCNyFxwaPZXLHeTeVV
DyTbnENphPldblXSGpZPtAaOGFQgG389YHV0uIFgKSyGyKfjl9f+QoBth5zOMtFU
3/GvHh5VKtW1Q08z8KanQ0LvfOCRefdtGyMZzWMhCyFgbUiNHbfXB6cKxBLGdkVc
r9ywmiJherd5y7zNQrkM29cHLMK4oe2x1EiS6LvwWLNSZGJZlcH9ym2s1S6fdysH
Zva2nWgcH1gw0zdVAY/2IJh85vox0FvQmAt4vJ7aGvix3mTvyubs8Dk/dt0tUvc2
NthfzxWJ96sR/eMMhvuCJYlYaVAXNSSnIs+Tz/UIBq7e4bKuu1JKAO9Wh0DXJ57j
oDCuXHa5iLI5CXrueVGs1u5IQFDCKYmuoLDvIRYFUae6CvrIsp0vyMbEOeSAcCJs
`protect END_PROTECTED
