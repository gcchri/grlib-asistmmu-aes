`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bd23/ggigH5cIjd4X5vgD73d6hzXAQCLEdAudRpY0EQ7gkK6PkhXJK89+WFaDV/K
lnYDvA2TbVKwwMfMvqzrTVyzx3H4jpue3113cQviFG9/foCpypwWG4YxgT2ViuJF
o7T+ABF1LCWoAPkfm4pkNXr9LIQXPX1ZbWhN4t0mkr2FsHFZBVvdFUXEBp8Y20uc
KRAAw0FJQu5STe6ksxfiua6ttiCW6MYWPSmnRjuCrw6s1i7uOLpekDB/tnERRVbK
qIizJqgDi2JWpc49Mxt2d0tf58ncjvBEOrJSsYBHu3MWZAA0rwGcZC851Er0IxVa
MqmYGatodApIhQWxT3AECrAM1xllxQdQycr5mCYrA3oezeZwOKPRjWmc00oRsXxe
w6/yE1OfDQsL6a7S+d9y0NA5/ja/oxpfvwMr668WE7c=
`protect END_PROTECTED
