`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MQ6uBSD1HSIi46lPrt57/UNIWKfqr7D/YyNTt81331dpx2uAtaNpLyFAkXDww66S
UVYrWqqS1fS17LYb6vm2cMUd0UvS4k3MClsNwwVWdqIs4qT/A/L5QjcSr7bBtFyx
yUr85NXGOybH2fnezuuSVwxsbtPtJi1u/55oZcJQM7+wNDh/NqVVp4X4My63bCkP
4GKL2vR8+G1Z30nOsyOZK9PmCf+qDnr0px6XlAlKh9rGcg8pwNNUpFTzTGMTH4/a
NecUvd5He2GXwyIhd4bASLeaQvBM055UzFKjgd2ZysXZxzRZPaZDY/qZ9/YUaQZx
rCIto2sRjrF+U4NG6KxFvzi33GFaKDo5l7lGkKCNEIAQIzZBxXpQmeyugqkes6Qa
ATQhXbdOkLYkD4dj/TKH6Oddjk38kWkJx+LPbI4CKOzJ1aaKqR4KmgWFDCZT4VRg
u2yLOQE+V/FyGutCf3jDkqtKpjaE1Yu7nYwi6/mw4meIRywlsXQQZTkoIVRcqvBd
ShL4voBqVKv1XD31JcFeLI+q5hs1w4DGe8YPZlvYiV8B+uO0lkro2MvtR0hdVhmz
KtZrYoExS1MYyQjGfvWA8uv1VALsaswRNDXDLvc35qqj2pcFfDYzcWDQR/mdOPkS
WtioMPJSl9Yrl5tt/LtNWQ==
`protect END_PROTECTED
