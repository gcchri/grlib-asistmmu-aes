`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/DNuJFuw9M0AlNXwpj0OBHibqIokC89ZcuZE5XWb/9MaFK5P4NeSnvNg5iuvihie
LmfbkBh97rKFf88cj2M1DdzD0b+uXWwOzDkFARSsoreUuF8j3x3Av5Szk1HJwBBz
38fSySi83RvZT6Jt4+TaRzYl/h9h8p+SpoS5Lut8hFX24FcurIfgBAxI68E54I62
HHhmxLP32ujyc5oSyhymyHtT3nhV/j/C1vjYn0+GrOxEYYgXacbmFfUlAJIvx/84
NT0kuc9vsKsGq5ccr+P0PWtkPK8vnZKHPcPh9jp4CQbpru6TMuA4NORqfrvTTPum
McqIxCJYmBaJGmkPzWnKcxL/f/igmVdoXaLnTJb1XKd/Ozx1mj1sMkTq/v/53jqu
3Fon5X9SXtvt5lW5Rvqky5Avc7KYNDiwDVFF8CbbhmW0s50pq5iGIMxuCP+wgvol
6zAPSIro6rTnum709SrPpQ==
`protect END_PROTECTED
