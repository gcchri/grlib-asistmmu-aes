`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xPYHiRkBtTCSYOWebEAPKHqT9cAs9e1+hyopuIjZfHJIHuP9GgULzcYPg5Bqquie
dU3fSwaBVH03SB+KF/RE+VE9EjXnYMxeEKg5njjlwAv89JbNXusDqC4CZVxFZKWF
mBBRMIKhsmvRSv8kwpO0vtOPEsocvBL+Il8Uhh5MN7T5NAT/Q1bon6LR6ivAepXD
6XvgLl5R5eHKO+5PhfYYou53XbsGuXPy5yhisyo1L/35KpyLL2FenGWRxQi1e6zB
xQDe6lXxdsM+zvHNzkPJWKYgcgp93+NIyKEP8uqY/PsSXaX6B34IzHe7EICvWk6b
BAK+UNiHODTDCvJIYUCSfnYSDf6BSa1rtyp1KFhyHVEqNS6tp2ywNjURbRZCdVCf
jrIrN2zfvtbOXSzeizAT+ymxAys/PucofsSspiz+rQqIzy6Uaerxxnv5QvtBdNRQ
`protect END_PROTECTED
