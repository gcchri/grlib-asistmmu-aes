`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DuupLg7q70jK1HZ72cableCfA1sBAHmQtP0yQwI0XYdWPeD2TVTo+O1u+FtLAaQo
1jdeiUmrKGAdoL5FQCBVha7IHE4cgZHFLIZu8Qb+CUo9F+pekkoqePEY+qd+QFja
sXqv6ldgMVEWNYyY/AW8iDUBok87Mb9jmnvy4k9N+z0oMsrzQhk6H7DfqIRfQu5v
8e4KkYoLKS7+uvUhl54npu2VmCu42i3ocrLG3gGnSSuAjg6fjh1VkiDZO5NNzpWn
9ZokgJ2/UQ4JGqkynjk4pRm+n1y6T8Yki1ILl7ZRmesC315gjRLCtzZmASsPevAu
XDgfpskjvSw1/HXsep7B0X8h/mHqsv7h69GPbDaiSvMvveYvV3G5Nfeye6UckiHl
eBcEsaFq3bw1iJPGXv9q4ESAN61aCHl/+/0mR6LAvgmLpeA35/ZdFVtbexP46NhF
AYst+AGMyHC7q8SH8gh+3G18EyConSJDKsbbdeu048sLR5/QfJXUGVAyblIQZNW4
vCmGIxkzzLfy4GEUqC5q+DLexrzT7N7hNJ0Fh6grbsNCakSCPVKXlxDmPay+Fhgh
4b0DBB/lT6e9aVQK8kNn8/ZI2pMKusaYRvJdPXX3t3yf2GzQV8FV3NNr9BXt/FUq
`protect END_PROTECTED
