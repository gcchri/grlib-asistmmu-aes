`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TM75zFpNtMiy6gdpZe7U50Me9niTBz/hT6oXl0RgavEDKoDevrxGC+Dj5YtwBuCl
qvurR+XEYS6+EXHmdtObrVQv7Chpv17t4XClbwMkLwlwH3eHmYo/0vg9UX7He1Uk
fyHNLqM6/2gVSCOMgbTwoHWE360eloxqhFIhaXkf1ahUBDD9NxBsaYt0XRw2fJNz
vSEslLraIqomsE3vyKgoYuZWd6VbUdjK+TMWSeBR/zUDtD4oaq1OCTIRzth3PdB5
wFL1RyEcfeuAEYA+jim24+7b+hWNhNHG6Z/hfUXoxqVxQRTMqG5i7BYxbj1pcyo0
`protect END_PROTECTED
