`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gvmaiKpJEjG1GuK/RURLfa1ZcMyDmgm1fxaEiMVWDF7RJfpsNb+Cz2OAMt2F0IfZ
MeZ2809g2wMXCa86LLLNAgNC75Kp3hjIgSnOMB9kdt35VtUs1I1EWk87w8mhQM0g
7bywReqWV3+i3WQoogpJUN04iLx41v/LAW92ExcbqoaxRxcaMTUoBFEF/StFSn/0
hRAQSyX8FzZmIVzC4Amp7IM/2kCBBlfd7hpyhP/pjZ+bg4kFyISzMEj1JILMCwZU
SM09p1rYkyaldOjQiu1MscNML8IfSSZzpyOtqW3ExMr5Bxvy3B17Ms+PDcXZs7kU
z2EHYPXBYtN8pdIEvyPjms/TuQzV/KpVLFMD8nf3KHmmE5hRammcFE4UBLYjfUie
YEOHSU2Odn7tALxvr8wsHsJSN2RpQg9qxuB+WjEgv0GWn2N5aycGN5rA30vORels
lf7+91pDihu/ZOv9ppc4rQ==
`protect END_PROTECTED
