`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5nMRrmSXQ0KDdVXJXkQegw3gbyhuYEzCl77vvJIJGH7R8myKBVR1oDZkOtn1af4
+/FQvSql7BgA79d6WjOLaElDTm5FdLPmVVp3q8WrxUhGWAmzHX3QSTqs20v/m/te
qiqvaA6dVPAijWv2mL7tEpqARQV4bPdLBDTLVZ5039CpuHbTOe1U4zy2tkWER+2M
N5onRyWCfD6a2OGt20wZ7/aBJPKaXQqmL32UxfmB2j6dMiBwCv/XeDAYQUg7BPMb
MZqlC0AyC4yjqCODv/patHgdWigo5Ydyn6mI84gHf6DdixDG/zpwqheNZrEzg6WL
VI1j6+Bw98ipII28QcrQ+WGKPFOqeLqceoqB0RI7bsaeR75o5JYBnxQPTCUMpcFu
zoMSMYlOxtXc9pIUisyIsh+2rkl+hCP83iCrPO184FZIEc1wXcAqW5Jk3/tDlFuP
PxBEuNxsuDzerHfZJmRkX7ZccLb9KX5X+Lv0c9Dwp2cvna/zOp6okeCvc7O/HJA+
VmlcI9l/EuhLBsRt+s3UTrEOwVRAsNrnPYJ8/okBo8xNIEaSmYGsDBYquTeprdez
307rSfZ5Mt+TsYouqaARbNhGZc6G1TvgpdkH73z/yCaq6Ei9o7JwfA2anLZTBXlL
zFv3uyVnVSJQVbtNA+I1aA==
`protect END_PROTECTED
