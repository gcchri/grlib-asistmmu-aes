`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
saeT8whhcZdHXyBiBEJflHadHJpgJIBHmtanOZ43C18yOImYTFFBPz3X9lbwZJDJ
cOxsrveou7G39RmUVJYSQyogcbq1BG6RJbwM9zOGjxPTy3c0IgcpJFpFG0o/11+4
3FHTwqhCLB3utNz1VDFeGAzAcOc5VIEp+4llfZyl0IERZuhBN4+pgH02rGnUIGO0
Sc+Vqqp6OKKi/x1+/E/mH7vRg+kHn1shgFHurHIwgZ5cRNgSA3dtMMQzc4Zj9Hx/
LifMAp3UWyBw63WIVbj2neJCKA2gYF30NHy/CWtBcqHCQOLr6rsBtydGfecMOZjE
B0kQJYqBr1DEx6HdxBnTxYryzkwfR0BXGD/7ujnwXyViyATNgeOZvsjCIZqMgc2B
+zSEjTb8KpNrm72xo1aCSuVoCFFW+qGtRfbpx2WqzLhFXDfvNA9xRkjTQ0/U0gji
UFum1YbG40dRvYNMBuafPCMSdAyVM9i2Z6Whgkn4Dkz0FEjcy4unLjW4StLSWGwF
54PVE2Yw/BRk87DqUawSHPOSoo3v/bpyGXPFSNZ+qDSjqmGBF6Uz27EOmLCBntkI
qO2OUjX4PNhZ1XC8ohWO9t+TMgTAq+jnxPUD3kMiC+0LCr+KhNhj2YJDs13dvOp1
4UnG9+6GHiQoS/xFtdIQBBHfej2997vRFCTHETdCc3xKa65GVHRgpZsxba0GHO/P
0lqtG3CEQStZuTR71GYUdV2IoKiyk3a4FWFZUUN1Bf3fopMU1EnZHYVJBd7UEbbG
MwzFnTbRiglL7/k9Ol+n4Dj3ENdm0BbnrP/1C5ZYBQUdm8e+quSVKz8IPadLNekC
sqXvCzmCylyPncz+On0HSBMMftwj/rG1R+KmOt7OynCwGY1xFR5Frqaq6LDqU6Gl
NZdM/r2Pi+gdAPzPZYLEF8EJowudvOv1lcWRXji5G9mNNQgn+W3bUv92YGggUJuD
DMSA29hIxE9bF8J/OC3kEkdPwcT3S47FXwaObqcH0LzBZVcUSB0AWLGtktyUgwqs
4nCQqKYcvkpa/3aJD3L6/LEvLlaTfg/eBE1wFtSj+df/MYFyIW99pw+E8YtDNvDs
EuN3yZqIypVGS2IdGf+drGbnKs3vbBadhi5MW470ewi+oMpEc+Yf5OiIdRnCk07/
nK69aOcVWgFh2jY41ID1NP7XP3nT3EgIkDi5h8PsQX17weakiAmNTCSIsNBD15Sd
TNQHb0P6+RrDUhvOiYYNRGQmHPpwmEzmkuCZ9IGDS5tst6xkgNBBaddxo6oV3jqy
2eujt63zJ+aOhNs5+aot+WZBicL8bWHezd+Pv03WcYb7CbSyKn6jGk2JFrLebXu4
Ir90GSKFla+JuuUYStFwKlTIotlRUB/jHH7nNBfMroR9V2enqYskKenDAtbZQS8t
oswEciLZpj74zSYQ2LF/5VRX6tSZDwbamh6J2J5+HYg6o0ySaFb01gW9lBS6wQnL
ETaOp2/mHheUf6Vef/gUpdvmdvT9YXmIgiy344eT6MZmpd4IgON1+sJSRcitjKZq
zsTnUvtV6RpgXbr2bMJLmvyC3VkvCR1ljetKckXiscnIZVNKxvH2LY1RaoOUqMHv
FWunO92fAmWmo75y4DesRcugcayhINVEU997HwSmhqM0vQqFzcm83V0waxJrXld4
bYpwLJU64gB+REzEJ1+2/9lhjwd2DU7y5/d6GUphPuYlahpXOjerlQp04Akg0bHJ
7g9BPX3PdWRmHxLGPl9UaA/7bOQWiwSjlwjbMYeAHMS947xPQUWwcRklaBJmXtUy
sQXPPkJhQ5tGS5w0bs42oubHAgqoVMrDjE8BP7F2X66wZwFMhz/dyKCuxQERwWmU
h2OkR/IiYvNPcQdFGU1jMFzNdq9elc0op7g3zij4gKH+13E5W8CVwyM4cN8EGi4F
rQM275R0xbYRLawhZ+B/qfJQKTmIEhuB39O51PUmgDDjM85c353sV2DnoVx9u6l0
qrv5CUFiwSC5CvFTqT2grKbZICF+3USwsLFrbnAMQJmKHSLrUZ6HVKFCoWqGGYtg
DZsVv8GhenZgaLZZMVuv2Nntoo7OZbzHJcedhkTWfIN16gKrSQHQlDJry6Jv4LM1
yWWXhEd6LxD8hbcWQYYwtXjvs+odpIzGg8/wNxZZPZVeoVwU4F0ATl5mnwddUYDi
`protect END_PROTECTED
