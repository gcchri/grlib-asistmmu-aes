`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1ckpO79WZTW3krA7W03kotNXjZVRUKbPkosoHXtulg15TI/CmHhe6bsuFeRgctu
bTjBUwS4rRsk9FWnRrULSP4TvFj98s9TqWK92ZW43u0FCEEabBLzvEFzqgBGGqM1
imd5PnitamJ5eslOsAC49ypL4JeNKvGAFVJwtot2ZS0N1nKGUONxJHUzK/rwRf5m
tKpbam+G4IwMUiOKXt99xH90f9iHno8pGTvMr4lCrrycZX3sPkOOnk8X3Ay89mGe
u1UyPcKV46h3t+W9FM/wYoK1jH56Q8u/8ijJxu15NwpuYTvKTbfWef7FpBjNmzkG
iyJzpPq6od9UppAJ+ZLkBUUr0Vh8vpAw/xcA/MYpS0IU9lZ/kdmgFK4lu2wcqPrf
qYAw4Byq2DAR7iCF95Vi3WDWLoaalCnLFpnmmXO2H5j2iOiG2KvBlpro15oChSN5
a5VUsVPmr4i6anA5fYIFGg==
`protect END_PROTECTED
