`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u76FZUp/JTMApc/HUsjWRPhs3Ktn9tEqhZ2aDnDmrGVWbJDOTnoH0oku53yrUd5R
yo9GT8DOGgiSzaT1/zWxBhIHrnyBf+Jx3NQVeMt64ziVKxBdi/Qpnlzmm6bZEJCV
8c3407wzFtqDLTPHGm57hTW15O3ZJf9AfrCRKhaz6nNxuRohbwkmt1WJQ0O/5wv0
SXJPATkoc+ZAkQKojsejEloGFo3soo7E7/bq9jmwlJ8Cl0Br0moWfOAKKLzI9nRA
SuCir/gsrzisdIV8I8eltQ==
`protect END_PROTECTED
