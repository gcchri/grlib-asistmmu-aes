`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rejJPaozlpydScFFzWId1lz37/RzAGaKn5bnTTicT3753isPguBYlRVI4ACGvo7
B7O2iZ2SREU6FV//2jhx9af2ZW156gY74FY4JL/dvSJs1vSyl7tKVp62vS8IG7o+
fmQDYGke3D8NITc6qCQCKCItNdU43zetZRChRI1QteYmTE09iosUYCt0aqhiYhm7
6fmbFxMVKQe8KSkCj1/3FrDQv7NQRUnffDIFC1Xazs9UUb0l1yRFY7Cw3UbJRcRR
y7QF95OJGGNmWJSi9xQU7xLn07/jabqTdOcceeJSJSl+Cl8bUtyftwt7TLJOC/WZ
ORfPEiYNTRsL/KABPRTsIbxoUU++QlG3YSW5XIjoPAASe4QjxJy/CyO9dN5nUlEK
q1yo6kW8bdZ0CHyIW1dFDphMptX+mIvI9rHYXPXElAhSksca6SAS6OolY0AdhkyL
ssc2XuRjfGLNlbm1c75e08kEwlEfqxv8ZmI3EQ3PthzEhu1mM51xJ0ump0cfGHBN
ZaNK/3sjTXjcRzokIwCxq2ad7aN1+mlQcoXc9N2IT6B1mIYCmoJbme1T5lLfzac5
hW2sNXz1ZFVDeRl35Ju+A47AMXbCAbQWncHzi8vL6T2tLpImhlpLf5O5FWEYIuAf
5pzf2/1R0hBIMSI0mgRmqQ==
`protect END_PROTECTED
