`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ZqnFIAaVPWOLl7K+ntsBSjFXwcmcrMHEI1pCQG90S4pl2COIlXi4G9vdLy5wCeI
CMWBD2BsVnhduzP1kjpm6CZ0AHjPTl0asZJMqceg0aNwM14e1oSZClUSHqjV5o02
kJgffDQQKpFxLQyBIIFmYUE9nxqbQCOT8ZGdLR40Zlm7v+Z8qrWqf2JE4FeVqa+i
xAWLJzbGA9Msi4JhQ23n1UDu/+mkDByvdtDtHrEb+2FTNEXRXWIQpA6g7kVZmceJ
6JHUJnpFHf2hu/X2cYY9YdyzSb+6Z/KjRiE5UmN8GM1IF/ALiga/VX33rOR1QmZ8
NCDMve5gV2pD5dzR0T0w0V2iy+Qxs1bqqe29k7ppFWL5uGpRGuTzBHk4ScF18xyv
mudWKxSVuilUT404uQ+56w==
`protect END_PROTECTED
