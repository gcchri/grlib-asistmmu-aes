`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRzspsBRNOHlHoC9tMBvHi2zj6lj5+M6ban4B47oIiM2TTyJkrY90LTqvVN7+PE/
Ud0l1UhOwXCF9FvyIwYAFXsx6Vasb8xwJuTPoKYU3M/kmXLarxYvqkllPiDIZgHU
GVFPShdURHOfSz2VlgprNpRoAyiQLGll1pd/ua/YWx9vHFuh9sp2Pcu2r/8dnRNn
ZVLqahEYRGmu6bvPIZJiZ1wkGJ5pPLvVdlB8ZFeCxLyzEfYTnd9b+MYIjg75+NKW
jtCZvoieniJk6x7tX9sZXV7n4wEDUWB1Sk/MvfuplRaY93LYd640zFCaCajE0Siz
`protect END_PROTECTED
