`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pNfqatzwazUVrubcQzkTOo1OOXi4oAoWOfQAewixqEkOu1sBEW45um3+mwFFiZbD
S9AwkQ4HPF36Op1grNGN7Iv7GhbAWnCXVSApROR1kMiHad+EjtREYP8KRzuJUXJC
BA82f+uIJgEsKLL9LkOwsf04E0GGkplGLf7lEj5tk+0pY3z1/+ZbFDRpDH+lmM+V
1amggyVGA864nKkmJY8mRGcB5lg9hxodH+qP9uVRuzA3X0nLoEbNygMRB6CE9XW8
UzNWDB46xt1Scg+rvZU1VNLT5zFDO9IJaAfkISwYgtiSlOjkxB6q5L/kwpqew1L1
UpHkf1lGOGf9rMj3RgVhQ3HN4xfEPIbTOVBWInxRLHD8Txk0NkGwNk1rC4WQMLxg
nyIdaxj5b2w57uGTwyT7eg21YSuCr4u4AkHOHze2IXdSk3/+++vc4ijS2fFTGbgK
4bXeqhEL5YxI1BTMZoHKruHgBm1BdCHSeWSmvXsIy/8iEtqmYJB9+li1c0beuh85
i9ta3W2oucl2FOxNU3xdWYg5k/wkQAflZJApdxJR0WJCps5bmIDZn2ujNmScTFEo
ewMwjrd+vpAg4smjMQHbtw2C4wBVqx0gWvlVZOKqoOmpf7Qn8Rz5kln7iUl3CGMI
M4X28sftinXRBlMicHEzRZ8ARMjHblNppdkkcjEK/Y2KozqH/8uQkBEKknXC40IM
ySe/ppgiM8LI+4zR983crDekpB5t3o70Unh0AUODPbEWcAvyBfWAwuWH27dofFOO
3v5k0UfnbI3qyK3j7S1iinkaJrlZEj28RE4ff583+zGLCTUAp3PKnxZCLUeOSqAr
WCbk9++O7sz0W1F2A/AjZ7tulgkhWS5HD81S07cGGX7T+v2PBViMrygsvMMvK3+i
bIZVKAnTgZEukmBoUlnbqUi0CeTyPdoJ2XnK49p0pTZ7RHHG5VTVCM9ED9Tzffh1
NbpwkfCM5zoThKsLvijsqqai7FA87le2lbdFVUX8NNtwYagztLxbRiBebf1MSc/q
hZQKgOjKyTuiI3vPbwdbOqni54Ih0ucTgHSp7BSh8F7pkxeQlj40eECRYgqZADTz
l9EqUu3TNwE9Sg7JdsXu9xVXBAw/FqREc2XMRe/CesvfoxOwMkW82zzw4EapUWpI
/QCwGUEHjZGUg6Ok6IWKOOf8Td84ibf5t/1VgnvDLXkkSVe28BxkFVX2uzipPiBH
H+TUrD6nXVnbH5xHRG4lWs8Mc+qaxfpDtMjEssF04aBYiF9A8YLL8cmTNU+sfuuR
0ACiYpcf1xgYL4WRZtPZTMbZrEUjx23xOv1UAKV40/uSDYmypNG1V+qZeVDDKiCL
panqiczs72Iflwq82kAyw8078mFI4osFFj4tYZvtjZK3dj9Pt7hb4E50olx0NzR5
0Ih7aFkH93R5Jptg/wXKa33yXMGCCdJnabIzirftiIFyAqhmVhsKKssx9LHxV4K4
EP4cIs/hv1A4vBDW7kYE6I3g84E4Z399SlfmLk6IX+TvjEqgR4JChNxBwC/tUcy5
HGhlQSekPG+06AIW9RceI6qHYJIiLha8PJ+itLtIZqrDyZ77NyNVudJ3Hm0buWK1
uzynugH6aVkgzvCwLyDBh2kXkoVkn2XU1xNI4mDWGO6O8nDgyzf2D5SLAoW98ogh
nID+Lb3/ioRJ2BkRMQhxdfMBPjgH1qnjO5Bc8pTJ7CYaPELIoH+HYixJOjDLHAxk
ayfCFs4mEutHiPr3HJ1dw0UDPhe31ACJbnAd4INgFVvRyrkG673AD1sMDs3uDbO9
`protect END_PROTECTED
