`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XT+JfIUkPjUdALsIjOvL6Khyq5s5Bpb7/Ngcki00vmD5Rcr8vTjy1QmGo45auHFc
I12CbylZw6xPiOcyZVz/cavqdwtz9vYMtqhv/7czdIIXd0D5/olGj1GtAFR8go8x
WkKTCLNcO5h0kS4SEhLXLJ1Qn85ibIiZYQCPWiBQl5oKcH8QXl35wgHnoD74BsGi
HX4v23JlGLemomVjjbvN2q3Ud40MOfIAdTuGpv3f9QioX/LAOBhoJBhsVnWXAiWq
YWvlekTFwe3QD+pI8tYewyIVxgX36CfFpCiGlPfQqRiN2Ta2yLzG0sCHi25mgB9y
odEaLX2k31zfWDpJyHOBRdJLdvYRkGUzbp11+6m2qTZbE03bGGH8FAJ736AJN+4d
sxQpCqOUsVM52SP8zgXb3j6cW4tT20cKSvZgIilcBQMoZjXdwgcfxCA3kDmWLHHL
290pXfVEpHHpeEeqwuQvn3hX8I5S05wdqGYYGbMINHbRY+lkoiap2o/F31HBgfx5
FaH+OMQcJ/1DDysVxMnjtXaJyKCQvdy+oo0UlB+d9B3h/tl1h23RuL0ZkLAf5szj
Lc7FSmS6FimV8LvrrIYs9nT0rKUjaycMt31zGel+n9I=
`protect END_PROTECTED
