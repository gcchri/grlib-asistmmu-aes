`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLLws8wkmpIX5IvI2q8bYzzRt8I3LMpYt+TgmpojgxL277IW71C1YbMSPU1Hizjt
S9mY+jiSW3I7yKZuf7WzK1mBvL1+fMK5O7DA4qw9JdLl63ctpD9MFdQaBdWQpyph
UM+ensqOZE2OnB6/vIXeN6tH/0ty5cXuE27AbqCY6jcPBtsJhyMU9jTsGnM+tHey
LmJFmWg7MfrLg5/L4867vBmtSrsglyffyU+6Sem+Hv+3ogcsEGCXhmFeYP+4ey8e
pbsmqZxJeQGKc6yFhYv9m2JFEoEeVPtwUV0s19wcHwKXi14Rox6Zh+4dKe91aiSB
nfl14NXvctQgl86Xl+UXR/Tgu0WCe7VhvdFfr+X3EHqUfQ8qbKwqc65HpFHmqBxL
bxLX09N53LsdPLLmmnwPzijkMwvNnYrvFkxHh8271AQempnEMZ5hHLS+w8iLl0xl
NOSCED5U+/uCxp+8YbwwL4Nak74ztTwowKaaoOCnF58qHNDuCsr8nWbEETD4IjJo
KSfB7y2/HthymtG1ntyr/SCX7NIBPEDR58QLp1dqPZexGCxTMB49OdViTHtGO13e
1G0Repq9whPJTQHhPzIHbOgKSfq51Om9fqG5ioDPUzV4gXrexd9cduyoWdLYZxDe
qB+6UO5Nwt1O2ZzCV7JqfOdCVpzN+hFs6LvbDSYEXnQf5SRONb6jMaoNaMKiRiCI
6j750bckr/ClBthEyMM2/ujxNoCutUYbh6phiPNSMIbvBjPks6NFsWJ+jSWoKyYK
Z8BfsZ+KKk6JwuB74x+N9HjARNn0XipKwDIb2gkQ0nVjmOSXR6Xmx2pldHoOEW80
y2+KYUJ0SXXBFsqEJsjtklHYHblaxLegbrT3aI0/Rn7xW/OnZ5rE+WXBzg/Hlyhf
YtOMw89r9U4NkLBhy5lMleQipfrdhgHbmnHSkqVW/flRNJxGlXXsoE1goFVytKEx
meinAPFklakPsG73sFKXOobpPhDRcv+eNMbzhixH3vA=
`protect END_PROTECTED
