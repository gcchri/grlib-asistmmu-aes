`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uW37REISaG/+0tHk34N/NEgo8IOYn/TSffPJx0/0KThJmzGpTA9BkJMixuGGGg+e
FZre+sq9Hk7oKSeA1CMTO9GMjfX+KiaNl41jLIaf9d8Mc9eliIA01LDSJbAAtkoS
dW1drqWoe/1izUvkBDd682BM++0zdcG5pMy3AemO86oLMI8aLQYpaawjfAXKO+3D
QXgbK+ei6KRElR2Hw0cLuPJqst9VGNP5SY0dghuhsXZ4nc1NqRvUkzauzp9mlgB3
shBrik6KL9A5Es1HMM9DTOXKPcT+T85mtYTrAoXdK9kd80PEH6xBbUf1wpnVA04N
ux2O2WCnUo8dCcUbu/q3lX7k5ogn1kGSueswStQhe/jPDExk5I3uVem6rMeyUaO8
D1v/IVDUzlfHOTxZbSA0h5edEuhbahbYRfMhlHmluoriXekHS+jl5csOB2r0q6P7
ycQEGiTVYY6Anf/SnAJZDy5LXGiXlHInPE6EW3tuTPB0ZV8cgDjPG3inC6TzXKQr
8MYtvwXrDfGHDNPLpeSzzp5faYmd+N5x7OHxPEI6ZM1qDCnwYZcFsaeYIcN0fr+V
Ef6lNUmTC/0bCRcrj55kXJZdsPr37/DKYaSkvppLP/WTw8hu56k1r411IzMDq1Mk
/rRwMgjIpYnzDF3NrmFi1EUDcm9bI3QmqBYw6gsM9EYWhGqBql9ccn3MF3F55V3U
LE7Qkjy+Hawjz7kqCa5pPkMH8uxZCfuXV1cBYrrB5J8016CylO78glH4l/0GIBUB
m29lVFdfB7JgL4E2TVK0vQFeA3oBLmmwg+Q0IqYMW0yKj3y1WqQgopI9OBNFtbyc
`protect END_PROTECTED
