`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dnvrFT1dmzDOBo5CCpL0Ve8MR1iWMFl137VdRPwqtQjg8HAXLUmmwXidAw/Z9rJ
L71WX/ZLLCopcPZEp/SY0CcnS7eBKKlVPVvwkiZOjIndNMAQLHMkSED3U34zEHP2
b9EbrqhBYLiiywyox/u6sgR6FNsgO8D1D5IV2LCm75ohFCVqSRQb6s7cDcFliBPy
wFVmOIqrBckXQ3Z9g1G68MYC5xxaK/54lnB36+1bhbrDpD0w8F4ylli4bhBFoMUk
SQ5uRtiUgKIRlHmKNcUxKg==
`protect END_PROTECTED
