`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjCwjFxVMD9CE5vnwsL8sLeQfOLCCepfjjid8Gp0NtAxmMUeHZaDQQEztuyKyA4Z
Pj7aROWhhwzXGQ+J4oNyrcAL6W1C/Qb/mP6Jx9ck4+G5TMOwD0/lBiM8NTWfqhtw
AfuTnagslLaVpiDjfxfH2deCr9SfQQ/uNyLyUbvaoPkbxKq0NifhKM3rr+b+ltlD
nMzOlrkC6jwSKv8waFZEopfjcaLUv+DkbSlVoGA4Zh2BM7kTr3N3jojbAV4Edokt
R/xM7VJ5XpjXmMm2Ur3TmXZe3nD5x8xpW9c8WYvK7ARTgnXVKxuETMoKmfB1KQav
8g5jicRnn466VFuprh+TaeRre6yGcwNEDSJzG6xon36ezR5Q2hPQTFze+QqyQJyR
ADa+ZroGu0Jb+kgt2fxUqPk0EugGuWXz4otYQ1m1UmvYySsGHOZkyT7QvYz4c/Gp
9Q6gQLexI6+fvPn5ZzIyzpljX+x2XWNA9b1xtQH7WsRQEgAjBNdyp1klpKqYZHmm
6fGFPpdscYzLA+luDXcE1IY1QKFjGs81LNQ5yQTejqy4IlouPiHXx/L5P+N0SdE3
n1lqHyj+LaSwFLdop1q4mPRZdXzGERDr9nMJNXTbEJoTedGSvKQGgzk55g6zd0OY
nPy3itMQvEUHwHhu6VNfevxoUIevYRVzvKuZtr8pJo09HrCARnREaXBcamLzZTub
UKy3qELL0E1y6b16J4NOlK0kVGNZ9u8hds7IJWmKF/c=
`protect END_PROTECTED
