`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qZb5UVMlfsNQesX1jImVd24cZoPLhnkt6iXNe9xVuX/f9CNjM6LpjOq6eh50Ou5H
699ENk8xaRLqIN39vR8nMKy2zctEzAz0zW5aQsR+g9X0RPoPp+gtUv/iCWWJzhbm
6lZNvG6WcYtKIIJQJmbLw8/ePW9tc8pK6/54rIBIW28bEc+YYmEpnhElnzJgmoxA
saCs/Tfum09EmRth0NB4p25dR3rtUx8rpj37vWDoBZ8BkKy2KqMOSU4jV25AXZ5q
5MK14WVUTgSZhSuVAzg7pQ==
`protect END_PROTECTED
