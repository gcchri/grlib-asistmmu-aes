`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J4B8fPibAdH8OMZBi/k2y/LTbg/xWihGKuQGhg3tt+2+VGCV8b1zoXmwbiPQle9w
6jIALmT0ocnNTVLjU2cnDmjXmi4vwdQTGHphIm+8dOClFA6IxHm/RbpSn6F1BeOB
SOQLeNpP4/XF7UwC2TNg1A8Yv8ZG0sAz2cVC9oy8uiSMq6nYo/0EIU/YoB50dnto
glWNiL90artnbL5N2t3ZnY/F8FIo6BKaosFkcqieMvLfOctKcKaHR/h7ArJb7lLH
0uU0cZ7smuMbgtCoLgd44j2YggIBpvWeeYz8dq0+j2QcnS9jcVb7Ew+2PWEyA4s9
YnJNxg92PzuXFPrZlcJJMZzrfA8DuPYVL6FSlUkrjRndNLqCHdGLdlcJtu1YsU4t
cPyCGPYYWzT/oVP1Epe1txlF0Z81NPjV+WYHU+X4NHAwkC5Z4cb45M9LsX48ppvT
ahj0UOdpMr/NEn0Ln9Ve9pw1Wl0FH9RHNmzLJZpJHWDKeqA7oGT9fNFUXH5BFsKF
MPEhNWTwyUa8SHizDbmyK++Cngc17AyA6Zm3dLyZWgVSkY1SdORJW7YNXSvrZu4Q
b8N94FDpiXOHHZHCrfUlAQ==
`protect END_PROTECTED
