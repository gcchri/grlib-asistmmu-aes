`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yRY9HQCnLFe8N9ncU6zg5kXoNPu7lci9StIusZXGR4uQ+f7zt/ev7oCaZp96AaeA
+vc7R72HFUKmYgstmCmAMTedrCdc9QDDfHeNXD8TY/byuSfMBPCm0uaV8RXv4jsG
YqEeEtlAu1DmHoIkL7UlcATKKkLTee+C+pf2d5Qkp98jlSCU32NITIFyUQt8pzf6
lJmMdmc2K8FhQJXuaGKrgpOBMLhV9BzjejcsaKthok/bmBVE5wD//+opQz0GEBAr
HFeR2/oXkIWoi4+hxBUjVpWgxe/Xzd0sQR3WRetCaf1q9P2sV1VZ2bv3Bs8oEZxx
/WtU36swwk3XR7NBJPpzwqdCqOOMPdVSB8raIaHY8yNFUNcDJKZ//hqiOIxhVSTO
UwJVuU3VCkpiSTZrK5O4iVWVJhLOGE2+FHNZiSeapw0DkxSDFAJhjO/aqUNbZt7M
ebsGZg3jwUZwtkT7Lihw+vxBxAgO/RDoor1ww7AhKkQ=
`protect END_PROTECTED
