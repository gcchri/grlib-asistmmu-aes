`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vTJQhhWAnuI1mET94DTNGjdOF1VcbrYOqeliHwX9QMqljrRskJRiQTQqqm84w11C
FwGmIThLAGkLQyKxz3YXvl2Jj3B11x8KAleHZbwQOeFxlkdMBDuwtj01HCfNzHQH
NS1aGB8Ytn9oqpnwtQ6hruWxCHDM0ttxwkV6Ax84zcs7C37Gg6eL371LbkJUUGcI
pqclyIqnYHwG8SOk7D6kYzsdar97tQCFG8/mDBSp9W+NNvXtRJBmKL3bkcQ5xbfF
qlFreOzMtdiveCRKhlqhZe2vgCHmB1vcbeOa3zchHufWaJ5uWadEP3wdMu/o4d/O
xDxUnDhxF6kqerXyQ1aW2uL0F65XtLCAelWH69swsI+Url03MquWi8zp8cICYgdz
tbqsQadPAbNlz+DmRkzXaA==
`protect END_PROTECTED
