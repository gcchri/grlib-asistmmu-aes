`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DEJSkLl1KqXXEiGPSAlV8/tLc71LGgO1SyN3rAvwnmF8qNtgY4PO/tH79xhfWgl8
vfXGNzf1breb4wVZtXxfORFIe9eJXbj5ncfTaCO3Wst2iQZlyVKxvzYUTtmefpFZ
Opaa33GWwvwRB5oLzitfhmle9Xl7JyEtLVzPx41Pizm06D1x+HsV/0lgf+WGGWtp
vElontNXOjOCE6ZRFNWXj6RGfnvMdivshv0dJ81axwj1L7GC5aWWAfL6LOpLFwYc
+B0lrPDaRqVWe6Jzg50ZJ+J4WTFP/erocmCSEz00oZc6mb6AIYckmDMv2ul4QYWR
Q2oKau/QBmu29RgqbjeKNPyZ195E1a2glZZbVB9Qaehw5HldDmViwTp7kYc5VWgv
/GDPiqFxV/fZUjn6yl2m8RC1AY8lP0DznGAgFOsXrSzAwKzhcLFTQ4TCgLhBLfhU
mmzXbipIdw18QauATn13viFO19rExUwV/MPATMN20s8OKuRfUnB3WjG7F9ttZnyh
RV6SGANcKjoOMp5ZfhvaoHTfHzAe8MlYBPBdKxxLwOqlSptKKlIW6pnNDD17jKvd
`protect END_PROTECTED
