`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MrPi51k0wN5EEPqEZE0ptPISKOt6yoWsyA/GWjVBLhLcNaXnnJEdC5d/6QvuG3Q
y2xCm1OXaHF61kb3lYOIn52j8MY3da7Hp8byjnnaj6z5XsN9BRQUqLkPfSlays67
JWJdIcjKKiggtTDFIY2JdiAJiDgikZetjTK2eakPoi5icActbGG9QlURc7J/asLe
nmbFHU8IFYYnOvEs9/3J4m97rlUG4NL1//DZzXmZrwME5MFYmL+kq/Y7P73tq+cu
YC8cVjR8uNgx7ygp7qUPctpxMeGL5oFkFxsq3VaWLCOqdnvXoQhR1/gMuAJ3JxSw
7vY+xPzf4A9eWizE/TroUOvuXVtUZ4t37bLU5She/If0tbcmnLkcDbDjOJ8Z7hRq
ta795SeWjlvO0UjqvGGdKb0mAv3uIsr6bZMrZrtiqPmR+7wtFjPl5Yc2nAmmKSrs
hHqlcyoYBHkmEVgScr0quhlbR+aX1bl9cikwz3qxbfLQeI3u+DFt6bibrLT9BlWV
FhzJqCKgOHF1H02YdV4RSY/l+d7pYk13fMai4jZr/8b26XcnPvhBTS8f/KkN2C4O
2MpjMx902/cYHNo2d5BEzCijfVasUX6fwLvKPB4QjXthor1Fk31Mtl76FJW/i4wB
YFwflg6XdpqVapVd6dr3h6LxLgyl3agij8g9ZwzpoMtrLmEhotTxqkMHhNdNmerJ
dC6la5m1eV/hWnTGC/ZxmfRhmTppUwLjbEm2DzSHBelgKuVwu69sj0C+AW+BCcfU
bLdKYjxINvDOD894gDRL9i5YuV1ov+UVj2/km0pnh85hSz3bOV1ffZoBDdJl2G4x
HXrOm5ikv3cAxJLKhH0AsMGAUc+NhBnM5YxsU5c3nuvK6HIMVyOAB+d686DPZQxf
7UEuzTEEqg952T8aex/+3S0KZfuGfCxZlNlCE+dyoWAge6ExZ7WZyjJKAgV3zLTO
UpGzv6ElSxrye9bmlR1M+OPJtI6APPx4gMDr5N/kB/9ghYps2LlU0od9bHrbUwJK
AmB6A9eZBQdtfTtb2TP8gUrcpkMbFD1xgGSN9TAJq+TNTCmYLnuD9J6nJZvnCtS4
zO4DsNAEGK7xTy+yDkRRz2jfJJ9veqZ1HST52DCW7LSChfluDm5M/S3BYnAUwj+6
`protect END_PROTECTED
