`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OryKs5XnngjzEphrRaf7ADxa8T6nEBPyOKxU8MhljpW8jwaNeaHgwJzGmKmgmQTm
wmSvvFPuI15Pb7yMKBUCypA6pdNVqHBq8BMyCSncjF/gqAWdGkNPGF/74QdnPcHT
z/hV6c4CxDckTwKZUME7V0zSm+dCT7/VpaiNcEKCZPVoI/3KNqpbqWp42NeQ1OGY
0e6DoPodIt18IuCvMPl5HFykVUgA4mYBFU3njpBzV8bosKbA04SdjyHNKU/6wJTQ
m7K6L3A9tmb0qp9KWOxyM/zpeJ2LYDTIwukgWZijpOIO6qRZxPuYb392/7GT7Q+b
DxDZmNp38iOBt15hNSdbmfAvANu2TEyFRVB3PWqYDd0hkpW5HBu0+c0NkfepfHb4
Y+KcPDWrBUWEQRFOX2QrSAciWVtvDj1jFhDZKlrTwTE=
`protect END_PROTECTED
