`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8QEfk77E6RRKDeZcaIpCWnLb+ZAnyn7LM8IA1Gfj4f/3TxSLpgNmYTXqubjINAY
uYmc4EZsLkT/dwW6EwCq0vc8Z8kxYrNLzQ6fo+uv91vrZ5HqQLFJz33McrgvRlvQ
NWNXI2emPK0NifD2DMcYbtfz2WG0EKx8n93vQxAqFsTzpxls8/35BwOuswmw9dyL
kQRYWigPydzCrdsjJdbfFsBDA5JMZfVsCjA8m9gZWraIJbKfge8khOkabCk8l14/
jXCBAUrCFKD6H3V6BZF3Jq3JtTRAbrhblLVV1P6Zd1NuOPRPWlVHLDrBp+xMeJT+
6vL+yAULZ+CfPRgOwaqtcQ==
`protect END_PROTECTED
