`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIVFbD0oiUTRbTf/vpU3i8w+3rQt0nP1gp+Oac8IHnu4xCXsmENCbyiq4L/I2u8F
iR9EJIo484uK8ZB4DcFTOsCYkmozmJin0ka3OVImNiw+CZ3r+V+RV3Huj3NTZV5c
atUMFnTpPf8q+fdiXcVu/YZXQGdxrUUTrg0ZJLPAhYcRSI+J2pXSfIABVSh3u7ls
WoTCj+jDyq45xnkSMGlXXFeA9w4ZHuuWIzj9WcOMqL91ygC+Sg9XFNvbEu6Yx1+5
wcTfz+aael0mZod0hQXtn34FSkLpGWk1Po9lR04qq1k=
`protect END_PROTECTED
