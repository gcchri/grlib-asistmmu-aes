`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CUs7BDaPOhlQ0drxhTbgZEhc2btaCgvaOUBJ4eQ16EHkBDYXIJZ9IIHfAP2ZugsU
3VW2lscmL8JKcEz+AHaGYqpVgE09TmopiTqCAc42PBaPo/vlEnKaOvcfRCOGWX7H
4lIUYoXM9D6U0MYcE5cEfb4ol8oNpMkrJgu6t+KQeH/L0/bguhWM/3DbCFTL1u2/
tDZ61WobI4nlbwJn0Gvsj19SDgQ15nlabK0QCrrpGqDEDREqF2VNn+/5oV4YNG3O
VgCE/5lupetDqsgjwjM2Ts+zSEHaNoK2MhSg1S23LqixZZoj0aaVK186RUGlt/lR
CyE5ZWOOBzAmNoTraGk/FGsGBBxx5abdNItIpdcN7m0N2ug6Nh+uGNyBjzkgRZFO
nEcfZwUsF0ItmNdWY5wN4Eg3F/sPa7FZm2T1iJbWRbdEjSL+x48vGLzKTM8qQCLK
loRx0pTkflccjWEu4mVaWIb4oLp/I3lbYpVOAZtyZxYZ3cHwiHzo11nYU16WyLj9
`protect END_PROTECTED
