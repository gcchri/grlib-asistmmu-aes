`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fzTMw6FzBkHurXoQ2M8cHE9OpxUbTSnlQJjB4NDd6iW9eMfrMUnkKb+kXeYe00oF
HVbMYfA9kwoqNPP/DsDj28aCd2gWsbLBhJSPYR8b+tij0TtrB//6bXY+48WwuP7r
XWP6MJbiS5yEoZoNzNOPxVvfVP14esfuOUGqW6IlBYFfJlkF5tKwFLqSVVJcwVz5
dKzaUSuJAo8+orPDTF0lRsAcJyfrl+/DK1ep5nRqkvbJlvLDQ0rwU4iRAzEW9mAu
tzOczoyEW9qebEVqahE0anFfYenU0Ep4buhZbhPM3CYRPANlefoE7j4qlXFtEgdK
tsgpRqIhOKKNOnYUZwetYBhX/oZVqMQv9Ju7lcc3xNEO7KTg92Kt/nrnx2nRvEDL
zFxfRb5yw00XnOKwZnRbWWk3oxZVKe+AF/0magiY7F4efS4bKPJJQws8KxrRnuyS
M1jgA48GVO7S4VOWvLAJuXscbG0jnDKrDue1OIMRUbrM8Ijf81ovKw5Bg0h/gGda
ln46d0ZvJi3VPGf0heW+9F83D4Jr2F6iar3lwpYhHjHMB9Z8x777tns+1qYExW09
G1aILBGE0W9SoerJcHHPCnB2J92whv/EaZtA95BXUsorvF51U0i1fWP9UqVYG+Qy
da0MH+L9+DOlhHeNIq1IHrpjJkdHcdRTAI7MqJsJ5kOSgWceqF4fp7EinMsclbHW
FthClOqQhAtaEkXf53MKRJDm15Bzoiyz9rh+toRac2ZTaEt1h4Z8FHHMhQyRe652
6IsfX5gHK6kdm5BUVLF9Ktjl09sa9u6n30TQLl5CSgh2TgVJ6WGnQgnCMLsCVcZH
DjNVds9WIJrRGYr+3fl20+Y2MyVhZl/CS27jxz/aTI8kY8bt3F5HqZEGUZQE6IA8
lFVTItZSViYOGd21+cRd1663V3Z54S4VKzjMUOImJZ16UlxwYEioop+l3e7JCZaA
`protect END_PROTECTED
