`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MsXn6VpWUgvTyHHEpM1VU1tuNfDi71noWdNoHLwC931joj90sFbVrszp1p6Ub6iv
pi9wlNUCUl3RQHAK8NSGH/JVD9d3VmJX0XMTZiufpS4yX9j7wazdwTJaUxGUATqt
5HhoIaFmqBdAXmgwb8rOofvdU4AwX+PQp/0T/ZDVNBhY1Yd89bG4ir3xL1Gmiyfg
mktlnTyj/aRXeAX8zVPDETG2GnXe6LFEJI8Gw7y82QWgNVfPqvaXj6X1c0G5FXh5
PaAZ/73AYtI59R9igiQLd/G0+QZ54VY/ew3jK94AObCMo1QVdYf7k8s+S0iJTMJx
PnkPM6KGapYLgHyRBXXG1B1H9KjfVgY1U55dl8VoLRQ8JjHo8FtV2VR+fheTbp/b
3hrzzehlccxTnaruGtpQ1xaew+tAluYuNZuy4HS9/xNMfBd+KpL0zgNtALaJQPXM
JwwxaBsK3Io89wYL4pxIU5BHuja5idu/jy1KulW0cG9nHFmH6PWM+Lmou6lZO7CK
MyN7vw2OCakbUYVGPb3gw1LVHIsK0Ed4jkmG9MNVxk0KW5RGukGFi1aGaFvvZ4wg
zRKwQI9T5/tJ6Ctaw7xAc8XitVuE7D/GuuEJQRIUlUa4Ips6Hb2xQlF57DwlRHwU
sz0M0S6OhUAfgLJAItVCn5U3EeBsXFuCUZtcPPfhyovcbwywcKvkY9ujm/Uy2gDf
agNE1rfxnXal82hhB4W16MXXv4m6S0r/b2CnEgnjhf4zrZCw2KImSodYcl1CAnhE
7INU6NBamMAF1dBuh66M2BemBlXkKOYCTE96RTmYjPjHG/HRPN5AV3IkeaN+yTmY
dsMBeVzfbi7CJIq97hm28/JduUT/jxo0ro07yvq+7lh5TLo3tAjxaVWkm20M9Y/K
jtpObTdxvG1IarAwRWL7miNrtaZn1LHB9VLp8XmXe8brSp3Zzw6nBQSaat36GKgR
`protect END_PROTECTED
