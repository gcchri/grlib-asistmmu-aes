`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4IzvhlS63iewFvyzvujUS4kH5DwNlU1fGdKUSasONpZQOZrj/dpSk7YkidU03pa
sPAsQMktwt6AJCPG/uPuH/SK3vlTMX/knNaKaBt/nm7g3wK46kbezejyZqbK/uu2
10kTTk1fgzBsoHmq7ywXXy8DXgS6mQW6Qi2EhNf5i38ib9r53bAms3UhL0ppSabS
I6bnXbhvvgg0q3vRfvVUH1eUU3PqyAwYXm422oJftC5aUF+i+yqf3g6gEFyXsVyi
JtPe0rKmRJY4v0zRBiYOJS7wMrHjtnmtUl3nYKa47Ut4yZ6vC4TSJWupCUaZEWZd
eW3o40WtyxAGgOgYZi1pn2lF957bc/vUewzV1TEF9yEGrexovmQkAhyIcZrRAMjA
JAIAPE9NWz9ntMD/bbxHNkRTy9f1/cZ12MH4YoiNuV2cc3Hxc9xS6Rpao4NvB/do
6ObxVk44Wsio40mnDhWVc6k9rK84lrc5UKsGq5RP0bXVW4QopSZuSxf1zqdLuZC0
2a4D8EMw9slmQm642jZTfQkLjNtWXhZRW3o3sGCVqhVhA4a6JcweTMe+BXp0re0f
iU+MxB9SLQlBoAESvFIvnQ==
`protect END_PROTECTED
