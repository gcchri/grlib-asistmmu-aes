`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRCr+6jm99etgtBqci41gUHCdYu68k/oMWIAONpHgn/FY2FmFFycsolePxrqRRwi
+2KdP9kX835d43o5NWhN2neRXzt59IWAk0ejAmQmZ+vvrgXmDMGYL7Lq0qe4vxgj
6uxBN3vyLpHy1ULzNrk0X6z38IimGmh4oCB1t4sDtmKLEvAGH5TEpfLqlOfYeZLp
Guw0lk2eGjDLDE7gTTgZanNwNQBKLzF7Rw31fWH5PjERY0j+9I09KdApY0vBhDrt
hqc1FsEGSqyMaCU3JwvmHi0XmUYoNGajzJw+lh0AR/V3ehQMaG004zHDcoMd7krS
fWxJEMhg4bMMRMDHmAoD8mkRVCpjOQT2D08x1iw8Rn/hHywFRIn63jpImQkG3jLo
WCv9l7xsqz6M9Rx8gXiCk5RgLjJe/r2dACM1GI+WrYPaWM3Hvzx7UIyWA5Ns6dZv
AatahG2XMdZCO2L9p/ztZrqIoC/YsBetiwqVyOOQ487pWvSaz70mx8MLR7HugkK7
3kIqjKpqYkZw+sfeDXtksb8TBGROZDlXq3v/0r6Ju2mHq/Xgl7w7tqL5xpDuaZac
tW25eFLZjg/NP1Faw53M9dV4JhwY0vpLvlJJnIclEDaGlfVDiWfaMpVjS4XN62GE
J/CddmxZocn3hN08xg4/TjCKfXoV1CmjJuEzmlLdfGrQyIBzW9vd+wyW7orJU8eo
YCtEHkVvjJi3iSq1m7mffrlvxbXHU4yXej5s6FH4kyY=
`protect END_PROTECTED
