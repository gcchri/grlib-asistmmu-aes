`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bIffhuSYQ1f35krN5BgcjkrsVj5ZxhSAkcdYuKptd6Eeu0+h1N6AhwyJoA5MQ3MZ
v+te783aCCxbZirr6rgBvtezcl82yVpB8aurWo+1fGha86EGIXPG1kWjXPtg6xut
sDIOvZP6JoVgFde1FP0KuFvtG/ELnLPFaEzpBrDX/3QdOv7ozK7+uU5Xcq2z5y8A
Y8Ju4XBtj83ywLd6r4NB9jaZIOdMcPLMJCp9/WnYmBkPR1UsP5WL5NElNnuFtgNf
nEIyjBwmonhKdbygFsINHQ==
`protect END_PROTECTED
