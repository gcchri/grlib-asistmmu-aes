`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lkpi1yoIXG711ghW4exk9B/t0HLAks1wQHqOYlE/uaRY1euxc+LCeYyKKQ/LjE8l
gTkqeGnOY20E5Mxo8CpPdlVK6IAXfkclHe17qD0Uubjlw3dZMjFLNV6pp53BLnD6
tcTg6kyllOTLuClcSSfXoQ6BOIBq7lopy0j+giE1NyZ2/F6DVsHito/rj3fa3gsd
/aGFaOW5ifLG/aDBB2uoNMYxekT+uHoZ1ekzjurzluAjoHYi/y6hnfOc1f9knUlI
yIrRZ9St7LWgl3T9SYggtEhNhGlulCwrumn36XynUT9cSMCN7eY1Gic6XkvGKxh3
s44JEb9xqkB9QExlQjnSVkjelOPdB8+YXX3qKHEl/uloqapuGvbHO4p3l7hRqCjP
quBT1rQng/C6KT20FO+OJT5p4XZkS3q4q4bZki/WVsKKivFyT9O1Wwvs+fGfWFk4
+h7zP9GSJiLzSbFTZXbuidJALk582HOJUsUvjfYgstS/wuJYwa6CIBCKal6eIysy
MnUsj+bCWBCKyIORO74jZSBzECMLUOXAVyuaTrESk6POYT5KMQAZjipUG4V3WUON
M2HRKPiRH4yTAVCwkzWl0Tpj9DfcNZfq9g+g4tYopCLcbZ3tlzwMvXqRUS5tSCe0
NGIBHwot0dAcAHUZVIGy2wI+N+PL+M+qDXQAFtvO3V3uRNTcJ9lXvxCxWEBV8oXi
01p+aUfiu/3geABXTChTUHz99Xgno+UiroaKX55YhN+IzdOZdGVkdN5K1pGQE+Z6
U32K3fM8mnePzRWm/x4hUnnfEdrYPFnHzqWRoxK4wLO0nMEyO2JPPU7WwxyEJFax
CYLSgjarCg4FXwGplbKW04OyIKtv+v4oVxHYHgws1fhqMh7MbJCKJWeaViH7raup
8lxFW8yqJgOzccagLKhED//FwZvCF8EEaPcMzH3VTB62KVlgi7UgDAGDlNLgGeJ7
NjTmh0uV7R+++ddqL2ngMM5ctPZeWq26nxK6qyf55xtLM+6kMathGQ5L/ZXMyU/Q
`protect END_PROTECTED
