`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJplXXRHqqjKHB6LxXai/eONTsdqgp4oxX+soWLz6Xq2TTpYbQukwrr8XOiiW9pO
HcaQC3sUTCYuNrhq4xqF+6UFbaWoAXYEGicuKOKnDtA5C15w2l2SQWYAmZMgjEzJ
kbOXcvvgTwCrXc8o+5UpZDMTtUSi1oeJm8m59Q744hzq+zSahVaViZu5CY4ezqnR
hQHqv7Em1vg687S1T7CZUvWUx6vVCQCDgRMWkQ3xWdrFzSngJBxq1unTth5EJnWN
P3nmCyVuAwe5t/mkiLoWBBg6+CS8xAlVN9lqdX4V+GwE9xRZgj79dZzCzDtaVj8f
1AN+4Mi9X3fwmNAujI/xT4OCocMHQiH57ZN2yI9HvH35MqTFlm0m6o9ll4dqNtv9
S7GowXt4pbQpFVFenVLX9xy+haWkUcn2gk5mcciT59DnmC9DMMblygB23ymYV7t7
Kjx1L1qFewufgxKIefqJ20Dv4h8M2Z2F0rrc9tfepj+pIlIkruePCJJjOiltc2qX
a/4jCqNpQhi5rPpERv1/adfYkTT94A7w0KywZTv/oxFYgrwbsrtKEQzrm2/lfkUU
bKsNI/53XqmvPm1Fe8NHXTFtuXKKj4I7XvBnLE54XcpLqwQZrWthB1eQ5GZvqF5Y
4jmcfeHtte08p8FqHZ+pOdoVeZkC4ydaaii8Njw77OIMqzhLQJZGTNtdKv6lDHpb
8wXxQaeOQoMhVQ9oyHu8FxP+PZ7pYO/i7itR1QudKJR4osYy9dD/xAfZ3zTkslHM
QFMwkLSdly25HNKbFto6McnORazY10SUGkDN1PpxEZk4/4KXlawGLdIA5ZGwW+Y6
gRrrtZstqF2fZSub0DeVjAWcKniI3cnyJhfZUxbVSA4GHv8rNQltPWV+W/2yzUXc
JygKuByimd3h5VHPFBm0yFeezI4HEP5aOWK6EoF5pHMdlp/wBjEIdXGJQfiK4FOb
Wg8aDEnTdwlEzOH46GVwNoVnGOsk/n9sWvwpDcAoOGE=
`protect END_PROTECTED
