`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8STAk1uBiR2XOX9jb/Fb6sbXq3+MpzVmz8aeTltGabhszW3WsVFviNbXLjfndqaI
Rg/BadBGcliVAM9FNypkK04rw22FclnTkm/bvk/H8hh9/qM4dka1OdVPxX/X32XY
hI9dyXPUoJpuSVkXrchMaC8TsaGUEskLCvDj99ZhMFLo7fevdooeSbHArGovD9gR
uBEXzcd7vOEfMQTmeR5M6uIZmj9DDVX/RcKrSgQ589Lez0eog47ydba8jsEnBJmE
9a0c+narXc9AObegGej39Dk7ha/uUYrx8dcNcSU3yvDuGwa3Ad6wFE3/7avqjShz
LoBjJb9+6NDXjL+offgNiFoss7Q2lg9SIjBZCdXX84x8VPShb0+M4foIkBne8ht5
ScV+4U9xC9H/JkEQ3IVmrQBJaliLK18fdkM41hW4+l5FLBOMPPOb93vccpEl3/Vq
AbN52vgGI75snaSGG1TctTg+dY5G/oJA9vvGQwKHOk5Xs5WiVEYCsE/US9vprZOn
jtR6hb2Zfvb9gr4ss5dw6/HGictBi45dFWv2OdwQ+kqwnkDskzEwjOVpapAhOH4c
7DcgsAP6IbLjbnSoNxh/9Bgpoj6sz73QTOJgmt7/fiPtbHfTo2604Z0W/vuZEJtk
zMCHd3S6wQsxMeDTY0OOgXP9ViUsKFBfgEh/3SP82jJHQiUBXXYbOjIh3gHCUAo4
W+VbBO7IF/esK1lCRX87iIPTeT8YcoomYm50VkLLoT2zBmUs+dYgolAXxR5eiNHK
oNsn+GdfOd1NEa8r2vouJXWGUzZ8UAzeJiLWr6AljUWZtt7LVuJ0gipzQMEfEoFW
Idyj2AbZlaQS8v/lGZ7Gs94Lgg+i92Nm3OggQdNbG8bHyPdL/YOWsXhlKpfXA5JW
ZX6v2wbAQK7SC8FAmfbWYNZA3iCT0MwBlcO3YmdBDlMGCHgg1/G1bM1qcQeRjlQ7
ZTsZHlS0x2sXZW81Erb12y92v+Uqy0uTij977iQ7EDhw4MH+eYn2ZBKzkdLgeFAc
q923dr8m8zXd5EVSOI7/gZp3tHPt+lT1ntpF6kJAa8nxvQYCf3TBVWzUdG/ZuL8V
C46UCdz7SbL3Tb/ZanvBvsj8O1+9iS8Se8jp6arQYPJvTlgDXJAxTZCREZna0SXd
2XTyT3fFd9vakF/9KgAHdGwVtomi1dnvltbip/xoQuyuleGzgB4CN69CVbUgCZZl
Ih5BYW/U33FV6g7BBS0L8mmpcfcaPcw2tb49pAJaTyscXIlqAJZXQoo7tIv8AY0U
2hj625DNK3m2bZJVH2WvD5G27alBcqsPz6uz1eWpUqVZGMgmvbCeII7Xd+Ms+2Kj
QQBZV8DxDiHr0EOD0t1LtRFQEkDABEG+GLeEX7EgLOvjUXZCRs4jOSWaiRuytAn7
ERZOgW0p1ElJolfc2G7fJqcHjOwpwG1OiqL4Jy3/2ENyXir4f9K6TjlfhHWe40cy
xBfsCcU0LEpA8Z2lq1HmznTF+XOpEt1Q2Dk4jD41YGeqXBVkAVWyC+DB//lh3DUt
DtROR4FYVbIeBQYRT8xZ80XNOZMLAQr41fwwHm/RABRZXBLRQRBxOPNfjiHzHJR6
f5LuY7lUjvgSCXvaEG86BRUDb7YrTQ3wNRCOAN6IFwacmV2gbRp2ha/ly9iF2YHj
fHAn+QRHb6DowVqDIF2fuqvwiZPO2BCXpm3GuqV6lMGCEH9D0Z872hYpIglGNzGL
JF4NYIS2o0Lua2yWxR74ChRtMOIGr5c2UG65Lx1N83pFCUvMIr7ROD1Vs4cpivKY
CyVB57mbGwcltsj4vnPbIY+A6d8c0u+aPg78M17ZCLl5dzBHk0mH4Bk4wEAbUTpi
9fAz4yMhLVGu2k6MQsrp0IGcxq9wDPpCyGd8Ubjk9g5hZhy70T5t+mSnHivXM1PM
EHVtCnEDz4/e0zFDgYHBCxMZmzILfPZbYGnViVmychNWA16PPTlfMpaUvM8bgblR
1D6pg/UQXxDJQu+oT+/vIyWhSPvEgmlB8VZDJOQY7irWs6ZN8l2pACqpko6lVsiN
Y8hR/1dFkNKzY6mnua+F2iGI9UW3whINdzuGoZd3AoLtsTdf8I8BaYFMmc4Vzooy
N3mfTJDEgi+YEhMx84Ykh3EVX554Qj7df9ht9pimxq85pqeBTN1h6faqKo3PcsdG
Gs81BuDNXv9EBD9qpjhRjZs1obzWq2+GSrmkAHejEJA=
`protect END_PROTECTED
