`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzLM13e3WsBE2YqXeRGuoiok8uFtD6iMckHp9Q38Fgi0UYXBw9zmGue0ujS7EC1i
2ZiWbeKS79EFfAWUPK4bAqGeLbIUx8DiND4+0PMGn8fY/pIt6AKOF+wJzYzN7Ev6
jsOt9zhxtZZa1qPc4v2KUKTqbxEb0O7Ic5y7GXhCdPcy18t7e6yX1jQtvMLxbyF9
q4nXi9WNQJqQ0MHgSmPI3Mr422+eB9YOHMItYZLKv8QueE8dhtL8EHDP+oauxQAr
kUSQ6LKA/MqoXlBZNHR4UMPkaaaUviTqXTajZh2Q0/HflMQeOvd5uTAQ6PQfEY6m
JdcODE7qGyg0C44zU/cESLDZyF8zlKCnEkmgxbjl312uEyRddriqJAL6iRcgb3ON
8ZJldhC6cfmdfdBjfNU1+4GfgG+xdxvzEMr0Jt3bornbucNzA1GFueQYLVFETtpU
5B1d3Ce0j+5hqCD+1y3v9mgczJzchW8TMKrZ3DMDs0M=
`protect END_PROTECTED
