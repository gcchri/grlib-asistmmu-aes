`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSbqv5EbsCPAWxEWzlR/er4MsPqIjjHzS37xhejkUGpZ69XvIKK4et9KQlgdXX1r
Hx6+Q5b/nUfddF2t41zE4Z/g4mCqWHX5iaMc3anNG281Dath4GFbB+khy7d5eab1
/UeH5rvLmQKfVFrjtvvrUlbMS/kj4Bh/wFMQr52rqqdMnDO1nPrNH1tsxkQB7CEw
T1TQqRq6g9db/m2h16ie79Bn15aRKWl/1ptnMKEdneuc5J3w0cmjTWYR2Ylcr5w/
G0BTPKOquD8qiKJinBYwgPqRYUDKrb7TL8RXFOnj/+qfSgjNYUSZ1sxSa049sUy6
TzsSC4PUTGH+/QWxi+LHwb3VtfesiZ52yLUltewYq4dISOrQYpsBzoPh8F/gOOPw
WMUNgK4ZCPd+u/xQEsNNyg==
`protect END_PROTECTED
