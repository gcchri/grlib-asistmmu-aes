`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eq9BcN7/2xj2L2qrYA00QzjXXZGADQmi3gt7UBAlcdHpTzbWgFo/RcULvKcT7HdM
EGj2eomYAXZ45tbQ/7tqvQvrjoIzZq3MpZ/BP9edaaXj83sv3AK7Kjww5+4HMoCG
Qqbmby7rXkfFtYnPs/mmhl0lUgXYKTxpKGNpHNV50wS7MH109yUWlew+2LE7QHa/
BY0vFWON9B6dsrJ143IRz5pbmtaAbGAZP1a7KZ2Pf0QD4KNvtldrz+hibnrK5KJY
ltoQf0CM1LYRIv8siTRLvD+x520EtFVkRWoJQn4mPbA4QrcIb5giT4Z+UkyZjYek
zfOnVY5KLBRU2+NoMobKHGf4faqY1U6UBuae1QrvCXH7z6TlH06+CKCg3QU5iltP
kb6nBit7a5tbcKB392MQlmn5Vsd4PEUb2uKFgojDbnc=
`protect END_PROTECTED
