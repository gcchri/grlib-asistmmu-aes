`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDZAHt0MoBg0rAW8lH4lcsGUytYEG6vay/ximXKhXJXVeLfCiOzzYl914W+S+nku
PcK1ZtT8zwDoMq5o6j+cnKElxtasXLTSy/EEEPG0m3vfc2iQykcCP0Ggwjfyllmo
XKvfnm7tE4QMp6Z4RB8kU9tGAGKvgBx72icvp3G8a+VkXaXMdQDYOtf3BzTYoUoa
SRsig5t6P1di80mrANciQOcac6eLzWRIff3jbagMFpp/ayZj860Jx6fJ0uSMsFyE
x2IwwoEby6irTrerIBFbnw==
`protect END_PROTECTED
