`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zy5PJJR1Yjr7UbEJDS0i1X4V7KZwOpjdJ+zy3km7NKkRb+nRsZQcarMDAZXaGWZ+
IIICZ+YppP9JDgExEj42xhN22W6N9z3dy/6kMNlZBZUQxlj8wK+8OFMWtiBVJzmc
ep7Ws7DtoGiOaTH97GN1+qTM2e6mPgRqaS9oS3k1HGWwGVA0S0NER5nZBFp5szRj
2sBhniL9qH9C19+mprrw5Aavc3MJ+gHvLflHg2yCZ7/skri6CftBUNaD1oHCQc+j
co+on2VCTPeYiuHDlYVEoNRVfXHIxT5IIfLlFEs+nldQu24Y8NGnxeFIsiTh4SrR
a7SNFFU22KYsGnuY5tpcHBOh1nInp13c/UtI7TgPdXYkv0rxJnViwa7Y6VSbZZjh
pTGelHHb+EzIRtGMfK8fsU+R3PDV23ysEqHu0ceYnbLvuK2xvV9YPHygtpO4FjRq
o1GfAtYclCwyVKVEGJ8XlPt02QtdQFmP2F1zx//4LMZKY5g/tvCVCvhvtAzJ2N8f
02m/DvCBzP7mf5UX5INCGnwFTj7u9+vc5ClTXhZkLIPnRkbchjl8xVHx50SLWrAo
thuT1aRwqXGD0rEJbT6EnedV5ZOpXSYJSS4MPlf5L/5c47XhObXmAWNKsLaxfp2p
F0WH997hHpfiHnQbVU6iP06MeWBmMYXfR106+S9DWv8=
`protect END_PROTECTED
