`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmgK0vBOX1jHXiKEcfz5h4karvk8G6wkWzjrbDyoJRpXR41bGOwHctuCN4hvG9vv
2g+ELhcK/jLbNFFYCQsXDZS2NhIfG6KSwB4wQbrlFpCgbmn3q5x21k+jS/A28Pad
88HXzcP7CbYhPvNnt4yzuZxheqRt0C4WMkJqHwx4EuqSjWcvkIbjzKfxvTj1nwaM
NkFJQTEM5BPCtREX6fFriLZtUMPYdZYzNkWBuBvPTq0vadit0b1ZN5UcJZf4J8a6
ZVrwyQZUu3iloJZMbB73z5wOJ7Jsve9Omz5rhVsRKsfmD2u9oe/FCzmNPLyrUp3C
tp+KV0KnsmVG/0lYIS54UezxBM3wqGECFNdpeOXitwMWj8lMv35028/T5UA2YE9m
gtQs6GRHVDIpaK///a9aJF/iNL9Pr52A9oYn+BCDinGAmL/eu4iSI0K2ILaxm92a
5caaAJcvzOT6Xm4QBrCW2KGL8KYxdGCJiYgbZmUNHwUZx9HwSvTfRDmO/H+ojd2R
UCPmYBMyBpfTmjCz6ps4FywyH8mNB2K2bC7AfLkBGVDV5Rud55TNT6J5K+sjpjUW
`protect END_PROTECTED
