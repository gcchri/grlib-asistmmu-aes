`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWaT2TZ8awFQezgGvEqnN4zBzCxN0Us1+n+bnTnuuMxC7v4iLCIzNs/UPkxE0F+u
PwoZuRuNladFA8+GXo9heqZC7ARiXSD9bHrL4zkydLtvY1urnvVF8ZM7izx4/Wqi
h3Q6JVYItUOk/IDPQWQVQKckTbA+OEj7OcX/vyuC/EMEjkNVE8PJaP6hM1VbQDFn
ODFTNBau1s/MyX+HxI5uaTh0+iOIql5E/B/3AxMHIKb2wy/8OXOkIiGABfJ61txh
F26l19IY/8BlbtzG2RG7RU4y50XLvopfNG9SjB9jmK01+C6DvtnO6lAtYUGOAt4o
/gVwA/vIGR7fIPY8oZTZZi8Kxv82ju2ctVypfNRjvNQOFXXoV1FAV1lbDnK/mBAQ
xR8WrPkBP5fImGPXsMDEwCHXDv9BR80pJe+gl2ektkNh5ttT8/QPkMyMvqobArpJ
/Lp8VwmBwXy2bapKEslC2jvvrn73lCONl6FLjsyouAcdLyhWSAkWKtgC19Zvb0Qw
`protect END_PROTECTED
