`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
shdtdmW2nOgzQ06XTERHtfHHXU2ATtcRX1JDdvy9WfP8necPWIUaw38zuKd9PR86
ky9RxUSWiwidVml4DD7Wd8qr6wJIzgROCUiQwmLQv+3i7mUKFM70jqBms+KTY9KN
abM0uSIUlJ6Xa8ui+CNCEo8+npa9qzAlNV/0BBgtggASgpJE9BfK0ukdzxD88IGf
7iXxNZ2iDLTt8Cij9ggRNyKL9ccb9jMB7kTC9ztb5MiCnSuJo8lrz6Or3+CO5y1Z
vWm3pKOOvXnxantlz+2SPHTqNQFJazHkTAFyr4oby9BO8FZ/F2hCUJC+OT2sleH4
q4nfBP4vlJOAvGoVwDpE++UYo7aniRZR+rvqOwxJgqnYFfou1REbIjpJtf2tNUvf
ERt5TtIIJLoA8gdf7MPRvIo173nQDdX2ZqaVpPTCGw7Zf5IugXcIiMVWQvoTcfE8
Wr5yv8Hzs+2PNImfxoaG6PuT9gr2kTvQv6/Ts5iPSCul5oxNZbqdthvudfeDRZTV
Mfik2Tu1HLCVSAdPOTdzM9bI7f7ocV7hHZQU+iBK5Eqo3GHeSPNZExqzkQ+bTmTx
PikrcXV7njddbbNeWe9ocmqhpomVqIJsUGthvyxJWHClIm003fCu/rj4SIWrFaxA
znD8IP8aKC6QgJeNVjrEAuPL/w0EyK6Qrn++O9IKvzyJueBkswG2UosvJk/D4g5h
gTQiUXrxgVHymqFTAaeBaczTlIH81Pn9VGKkopMTJWKvtA6fmZgw0fBrZ7jG0AsG
ly8JLD4dbTHdBIT186CJMLfcX5VQq4qi8XENtTvWMRkd1yOrt8may5SJ2+pNWeyr
UCw6FBnzroWxjHLeAOVUS0PrD+NVyqyELouC4RBOAZcSXFwJuqUsQ1s6nvFrEvOZ
B2r1BCVTQa+mIprRtRjIJGElmc2EWvaVH65+rqYpPDuQEK+wwaBcT8G1pV9IP3if
vPhFqgJ8G2/EWHapt/C6IvA2HNUcpQCrmhyp08kerrq9YipsENF8sFUS0f6HkY05
/6DdcfrxoSRF3nxODTkDlal0WOhdy43tqaFSe/P4ji9BaAaFQNk4wFvnl9Q9HljK
9lMANVINsc0X5eNtLGiZCFGq/BNDZcrlGgI8n1pUauVNI2GCgz8AypvYZVO6Taob
Bb7vVujUDJVx+QNjSRPvvX/pPDBEfbMjMj0fK5pNCPgdxEExzTEy3IwMCXsEfqNi
aMCXDeHYFy2XoqNyxelR1+0oZZ21P9OsQpdark1zV5P8xKMlrStMJSys3toU0WDJ
L3qyaqEPVeWio6SiWQ/W9QHIKT6xZ5T3uM8bZksoxsZRXLYwIW21M43XmCImlHmv
tyjPIe0w24DCWH1BFBn18tBBeeMrl7Nd4uZhPB1mOv07SrlTFdkdW4XDthyXSxxi
qoFBdIM+HorwQn1s5GPuqG/TvIy4wJEWIv9x8+hPJSEKHbPyjRomWvCTu3FDL/MG
GSkr+etllhPR1eBQw1g4Opp7Mel3fR/C1/mkKXZBWmJsudmwMbdCB7x9c5dr8N/U
eOuwbWtnYu21nD4NjTIP8mN827eQNlh/Eq4gsRVrpzuKPCEs6z+yNfvWQFRUplR7
GZHRuPsToBacqCKu1S2OpZPjFE/iP2q8wbFUl45/vseHRh9AGYhct50aoH0dFX9L
XXfnLKEFN+4IZ99qWPQtLMpRrcgDDLJ5WUnp7SBTGH1m0BchMKaWCUDGNcu9NZbk
JeT7qZjedgnwggn1r4rSq7OeN6bvQiU5dt31DGMIN3Q=
`protect END_PROTECTED
