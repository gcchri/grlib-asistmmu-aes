`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ui8ZzvxJEvWypy8v4MdEWfuT21SP1e8wFqx3BEEOZRSmNs+SZx9MPdljWobBLj2m
cBWquyMlEyvktc9DU8fKn/VS9Xqr52p3EtO4zO0nhzQ9e0zyuGREjIBpBcJzSF57
xe5wmQ+kx0+/NxNYK8Xjdnv9e7tPa8lWWU5HvIm3MsSKEGKtndRY7v+ACTGh3P7S
Ul9bjBR9e4CwGC7a6w9pR/LDj/sg7ZHfdWpaXiA68KahbmnFJnoEHs0jyCzgg2rv
L9J9DFhPxrmkqy4iZflgoGIeMGGozgnsDBWRAjxsJWWlzFgDdmgL1qxiJSD+LFzs
pHxp87hSwmj5QYbyhSYBbw==
`protect END_PROTECTED
