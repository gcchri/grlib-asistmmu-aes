`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
flRbiHvNNtYAxuEjMac0mtKTGPu3SDFPQ4BCMdXssHEYDV9AMHjy9+HBP/6BkrEU
wBUBl2zVJmCViWVSVkCt54pLIp2NQZyqe032WvRamzwRllSwFcODzPJNqfk88vXO
EtJ35s6rhWEGaNTtItZFu7tnv+zmbkbX/zPj9aa+BtfZCkuNQmakTUCpjQOWsaCA
7o5lL6EaeU3iGdaO9rWwuJ+Dqaa3omszv/gc1h7wZ6HWJXWZVO7OWkUr/yfaaPaw
zbjXuBBkkcFDF2nl8hZBKsHgPzsIjvRaTy82Hu80YKiX1U92nlSBRohHSVQx5vjx
YLJUyTblIKeRyt4tX8GGyB6znN+nn6/JTaZv2DO3rUZy5v9h0MV5gg9bMX2Vy5zy
FuSJPRzro5IE561aMnmbIo3FNZVP2RJXIk2XadK2oieKMIMPLMAnoF/N5Lyx1uj4
kYabo6STPJShdd0icDpiak2N8Jsj4iZQccFa0Ioa/UHB0Z751N/7mOil/FUmvqsO
fC7SqxhMzVKE3VP8bOZ1lYki15WaZGdKhn/GzmhWdUwgstgxpmXRlARbzTgY1YlY
m3cxCrierX+hO1Os92Iiuu9QSMX5LyTHeqd8mVJQdrcryD0Fc6T5ciiMQLHsP1LH
HdCxsZZeGgYAFZakoKlvHsvNRyvSZlwqMZhy732zBR01stGP4jHFmae5EyKavNpW
5d0Qp1hGzP+KZSmeN95+uobsfwULs76f9YyFuAoFJS+bRpsKNlYYe1wZzZ1U0UIP
1li2olJKqwiFI7K1nZhUXuYa4RkOnX2M/eYezC3gliV9bIcTmHcWu5AuM3NYW/CA
+BdWSjhlXefUcv5J9Qc65WHKcWCozE9WMCkrNICow+pfV60z4nwPQREhdjLbF0Nc
UNqUs7TSavR4vDC8sH7qpos2yYn6RbMo2+Je5hlz1krM2T2aMvnjNE9gU2XhSmnu
`protect END_PROTECTED
