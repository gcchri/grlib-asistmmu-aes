`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xjG2FXV1DCzk/tYgZHLFbvkO1So+phLi8iHGdQ1Qf6D6q4EOoZN3aDn9Rjkl3rDO
5Kyn1JeewWlaAKUI3QbXVtEQIYwOcAhY1ZK6viXR5EoCZT6ZVU80T012feWkpw7T
erVa6Xyxu4vR3BBeLLWYGjoFZTHD9dvLhhlKGEbZoccpPv7qSHNvW/mvnlQtGWLv
QC4iK0mvvZVnUFf7/1tSUJYUxyUviNepgcF8at7/EOdR3c9OA/pgDjOGbA5WRbwb
v6vnk9a6h1ex2HjW+0ih2g5kMYwNVff7z18d85tnD2ln33t+LuKdZTfvBpLOXecp
i3VOG9LVqbsGpa2dUwsA1fLFH73AbBCFtKs55S99+9QUh0aPTAPCj0IUlkGWG8Pa
E8PxR8C+Lvt2ogsbdsJ0HRuRWRgRvqs8JQLEbedj2zLNYTunYRY3mJp+/oxRRXRS
qpa8f9RG1rO+N4zroMr7ktSKzeHDp81OiDnquena6lk78QhdbEZy9haEwGmdB2aX
4ZblDkHAxueEI/FNdicegzsXp4JVGzGDSmmPO5Ar1Nw7qRLSVQrPvx6ZjfWxfr9S
TGXZaWx/fZcZXTztc9kT+Q==
`protect END_PROTECTED
