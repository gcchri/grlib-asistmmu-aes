`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiM3VNUpd5o1zB7/6O0Ktoelimwb3FQHA1y/gSCctxbkgC9gWAMGJmysqgbNAqCl
HUtbxh2/7secNlNgIxfQzFQW1GaXSgrLgVMcMJKsgt3wsMAPi5pOKHKE06YuTEvk
J3mBORf5I080OeKWpAAE/WRLimCmjxrfqF8SotvDOLQBxywsMQQIBWhpyrddfypF
3tD9AAO6YwCDOrz1LhEUSJAfiCdTGowNtBXTLSKquB1SjdrjpjJqyDOSex7m9qWY
OrFCWiKbb+YPHdA++X4dIBkUWf0v51/+Z3RPin3wstvhlHIcV6kZJfQ8VhuzDjvL
SXMV3ua8SbCHcibySRSKSazoZLhhrQKfqK6EBCOC8QVrdKrnZWeK+2i+hgMaCBWZ
d7/PKQOey15nYRCZtI4IXqJm4VzrIkKwwE8RtdchG9xZJSRe7Lxp3M26UvLU8G/i
D93L3KPcF2HgLGf+737SP9RC2I6W3Q6BIIX0AYsHuHBe0/J5qJCBWAfTL0MGY3N+
Pd04nKk6KP4X0XZSr2gUAyFL30WKX7m9l+AGzVcayAapJHQm+bnn18jT/cU49SvU
OX5/wD9x3sbYjeqYS/r+Nu668ocDXs+GskvpwUP+AfHtxZ6oMNswz3JBOJXroKn3
xDhgihtLQZTzKYv+XySuHEsRwVh9Nz9bt+lFwI4rsUSZ375SOfTiMkm5BDQYD44F
7kfIiSIKT0xAakdLJQG1pVTpUFrOe7A6p5x5oeNQUVdexgT9n3gIw4NfMQndsRTu
WJdgKI4QrBiTwtZXUa84WsNw5ZTfVrFT0E5fbm7Ke8+7/LyK2oNNjGwqpzKbo81w
KVM0FdUSqu/e6Wd4a/aByt6SQbpIZB4/A3asuXYaSiJZl4BKxxwZQ7N5AZCG0oNY
0PdEMD1q97WSyVMO4gd/NXlTDRmSMYvqhnawCaxILBHGcr6C4S1HEJ41f/QJIrGM
Rw7wi/dr3ehYpzPQdESsrqpPL/SGfjzD2JfQGNoKG6/EhJuu++ddtPr8e7NScU2P
ghTEkupTRvx9z12nUEkiD7SpJyEwj7gtXB4kyD/rIHPpymzHLc6ygvUeRJXtaYMC
7KAyrrMhuIlANAkupKeHgS11gTKtltZmb7W43OejqiYdtplF7VZVmktjAUtOuJV/
FExIgkR+c7oyma2Yo7kAngH0TIeHcVXavX+qfUH9tQDMazumW7Y7LewqhV2D9489
NQxvssFnxQIqTlKR2PqRy7nTL6pQT3xXHLmnksWYMHj0+jDTuDRWwwkwrapSXVK2
iYEEaw6AOC+xhUW6vNC9fI4B7va7gqfml1FUPGH57XqwTXxuBBF/h9BscrQ9PvC0
FGBCOLVH/AZXJ3yD00Cl7ZrE/FiJMfRKO6D6RHGf4JUN91P1piMWQat8Tm/UzK30
99JsxIbG4Auf6uC/VvjtkEaiR1pD0icHFgq0R9iCyEnHczjW2TJuWUellb1XVoNF
VfLfRvTL7xZrLYRZ1dw8rQS3O7rm4mZaPbXFJK8k8BXfVJtK8XZCIlZkZx3J/Ns3
ZWitqsj7IrUh7bAz7RYoZfnHOKoSUfI/0GsES3RTQkAaAtDhysNZjeGDnV5AuDmo
OmWN1zxPYunJ4HITs4L6717Hxg/+XmL8JLzH5f88A33tG+9Xw8hGDcTztlZMe3Pb
Cwut/afjwDAUZOssXxHsae+kVhI+Mj2iKV5jVfDUNWWpjmaOpPDn6xS+0o3qZ3at
rGkUFIEP5iTBsXLZ1e9Ef7JR0Vfr+AgUzXSH8Gd2gBPJ/hS0rROQfqjUP3tRpRyZ
77BluSDIIUXDxEM3AKfEQ/F8SjwTDNZDrdCaFYOKHedhDcAJFHrEWn6xSV4EwUvE
gZCF8JjiJ3P4k86zJFAZc/0yL60SsbC6Vey7Amuw8iccaFvPGHm+sw0V7PoeT7HG
AAdexubyx3qxbBsx4erUTJUpy0MCcQ/mQOxMYsQ0yzAY/zPEMYXHmpERJu0A7y5Q
06tMhi1OT329GGEkO5L8xbi1E+2LeCwDgDZrSPjHs/xKC6gflbUTvH53ecQyzWci
HeaWGNC6LaDiC5jOTvgezTzHboRESGqbBSmiBeJE+8lJHHTx8hsme0OOaaylpd4N
kDhHBtBDcuYJPnCWSnwNVKtilP+05qF+MR5YEAHJZ2G5fX5hzRj4gHTn0lbgibsX
27s7Ty9qECVPXS9jvziiLb4rYwzQBnOZu4VP4G72vRH/EMgxIsJqZ/+XGmqYzFzl
kv9NM3VknD4rOR1neuEu0+SBtpEOyPng8QtF/yzYqkB7z64N/mkNlzQeNwHHSocn
BIxd0whXUUrb2XdrO/fuzJ/xEeAvbVc9jjO3Lc5ndm+rysW/fyllbwHw2b81VbX6
O86M0l0amfADUuIm/s4jHL6BAVr0E7kWgZhSWHpEeWDnMGksY097KVtIKyCDHHc9
bcIeStrUmAvOMwDtDhkiMkDDq6crn3E/j7tdgqbvXVo6/xDfHz0Wbnc02cCu0/3Z
xcuzDWPxqjWQRN5Kt8C7F2TOGUVDl8DbnN2b5894i99Qa2gaNr1dqSZCjqICqRpa
K9CJj33kOH2jJp28/YWkj1JuLoVqM4LxRt7DISROieqBAzrTvWy44n8RYKzMfSAS
LUj3c3FjV1kv527lCCfDjQBIRirg4+seivwRWLtiCabc48OlKjDEYVIWgZXOF2GH
h5MHaOVCrLl4XdO58ZwwiosJx0t+D/lY5JXOPNqOPWRm5nDzXzPgWZUZeQ7g2w2M
Y4OeUiS/3WehFyYBRVZQJJJdHQdnqqT3I8m0xBx3igVakYw6aX22cojoyma+vfWD
HXaeI1eMNjDkgFggV2LU+bfMqT4q5PVIAsn6eSgs4yMLD9WTzFMnde1MzxFLhCtj
L8ke1hjjJK5xW6CvVnq104CcR+wX/aNa9U8UVIMZkZ3vXzTgbSwdL5veSEtQlxzt
0dskCrg3Li3SltUSV5wkfsfiuxBn9xrzi3BfKb84duvYo868wyQM+HfS+DLRTb+U
2MlHB6TUddjLuhjSCWCq2t4ejkV8UVtP31qpUrs3BuYv80d7acNCkKJlFc8GpwmP
sLQf09etTMRnAQSDyx+JtTocOyf3AjQ3Bh5eV+QIHVMyOgZATzkv10Fl7rMckPCj
l0iqMtRAaQUN9+Opb5eG+vSg5X9rQSZnAZ7gB2blhcQKs0tLH3s6Ao8A/ZEPofA7
y69XmZwgZrFWbKTOt5LjHVZxhuI7pkZszZsoZ5rMoaRDiGmCEoBfcfvbR4s4Ev/l
NQX0NawXNG3vYBY7GssvMlZgbjTzqlgh2dtDqKXAxcldIfxF+ewOrt90lnSSfuIz
XDi31vp6WEfY+0k2LrszwkuW1KekMwfFMKgkcCu/S+Q5F0EFy5JY2QMgi+jDOMbQ
B7QIr2uLFsbO3tYMzrUbeeMAIxFLImzroDD6S+V3YfL9UWFeVw2QCd9K7kMdC1HJ
R5UzoMDYmHM/0vfDyzntp5mX9ZVzfch9VtIZY4G6TIIaudbdBhm0qDMDB6hiwVd4
FsmotouZW3ihZW37mZkgbQJAj9AOFDCpwS6l1M3p13eWbBeMMinyArw6ugrpljwI
1MKaHfVGHSyPGc9T4n31EQNVgeKukuU5ge80YGLl7RHqudqdFgyNZxWtt4Ud6c+O
JUCIUGWa6jQ4tjmUGTiPQUJkAQr0I7tVolHe2stLgrdouG4Poriko8yioU1EDoTr
cPwUDBHA02a97OgFrwfVnxOBbhvg6w8dPgSLv5h/wwZIhMCoeulnnYT4cyNdjx0Q
/Rt5a85rZWdPbdlQicU2vW/osZV6PV6R5gkHn28ohJMx/x/twm6rBYdWayFHWHhR
tZme9B48A6zGuX4yh1sJy6UHJXQcA31xSHvLgisK3RzWF73fy+9D1xoT4IHd1HZ1
sg5v1tufyU3IqrKywrZveF8wIQzy1ttp4Got3McVCL/VYMJeRDhTNxVySEyeHCJf
n79yptjPybMT6L4jrBXlbiFV2Kk45GRBtySaL7aIKQcDGvvd/GuGXBr8gffMBZIC
mkG1q8Jyb9wSRpPWl+TQi3z3X4RAyzuSpt0AhEQelav4b66eCGkrCcvaEWLYDQEM
OcwoEryAOYGBs0FxkYmTnRv1a6ta1ZSCk1yiuWINw4ozORvn9S+GjKxY1S/ElKQ6
f4ohAptcKYvsmycv+SkkFuyWIHQIPJoWgquXTyTdZDYKEPTZpqfxpf833aJFm6Ol
0DSaR4ujlHXSnbyVbpqFOKcJy76CNBf2oAzbzkaGKmfQS/VfxmWuVFbVBKO7dWyR
FfNIbwvMh5YVguJD5PjnpANS7fPlaKt9nLhs1fvb/R6o2eEHOtF/DSYxvMR8dKk/
7K2anyOt/uq/33qwanuWPVVIGnzf0wU3//rHiDTLm1+LYdQ4PqV2juuIlfxOd/0m
pgcXA5+/XqNMTTrr/1SVqiE4C7HM8l7dnhNcSkiZ+XJ/7RrDOjk7siUbi5ZeJ24W
2FXnjUnVX5z/DarCktQrnk11sP3ql1oFlYkOkHOTIxISW2VYIfqAkkdbe4kI8XZY
/OyUzdEoJEqfsU37a8az+5/ndI6hDrVZDwkGWS0luZXGLJ3FUkductFkmx9dtDRW
5guPm4j208/RPWr0oa/j2HBKbZDYtmiXVEjUvkFST4VnHE/ziGsIpVEKzr8m1H2x
CIfYxt7gov3zB+EfQS+WVLL2zEN5v7on3f8BESt2vnhGoY31hKmt1oCanuwI3S00
TclEyZ1TojAU9lDWiI7/ASBAg0WFsYpS9YyMGLC3xOBXRLssFX7PVlf89K1ivBm1
9ngiXH7f0WSJx7ZW99wvHlvE0xK51VxNU9Qtk6whuCRAqovInvBVWwf7a31w5Vn4
DB/XLtOjAHKzgaFBi9FTaEFZeFVKDAJX9LU91CRmRWZmqLiPutkNYUKxfNNqbxF1
/KfXlQQcttAyVQ3lrSJxTE2+j5q5t26a5aSd8l8g0vh92gPszWfl1+zdKIfJBFpd
mhXxAOhUTVZFRQPMFNS875c5xrLOj+AEAMb8ZKvpPE+KRW0e/buMlYJGU7Q0zsAY
V77+3xTiYo/j0vCnIJnmsc3VDhQsOPpMXiibA1gKyR/Dl0YdP/oNfb7sAvvyOTdv
TvODNZ/pNTFqlWhAH2qNHGPUTFR+nbNwcr79TDLV0YjpdEZBdvE2gUdIXJQC5uAE
B9G2Y4hXz6vWDuxXgnNC7XLQZdVn/7bwiq8O62yh8KMWfz0udicARd2X68KYn2dM
4+5ozdtTPk9Wrw/zb5+2LcwV/+HkaHd68k0zr809xJ4ehcqtbhOsQjjzICbfKG05
el9S0RCYk3vXB9veU3A7O8o9dFcjUSuiY1Hf32olHYiZMeeRxdGRPBl7dihnL5t1
u4wR96Kmb1rAu978h/NDRlTkc47GWWM2Up3v5g8xzR37i/YDb92DA1rNXFrqhjRJ
HWzrYaXvHhyguQ7etKvZ5OE9wj18bpJsv1oPLyTzsujC+vzt/RRS6wqwl4RsWEVN
tm+f0QLPmjNGshCvqCFuK+Wikmp4ppYtq0QJRGeobJ14O8lTdd9F6ZTCH0WAYA1Y
4lcEErmDVv570+cxKkDSHW7kDajqT99QO44A9EQfExJPXlrF1mqwIXQQy6EPgOsA
6MEbitEspDOLYNhtyuWQgwFs4U3EhN3Csr2dYR8VUshQwdhtjCbGgIBa0DrJni1q
4eyHegV+Ec1yZduqZVlHLfxM3Cok2gZo6bRfpErAZv9NCtd8PCLvLc0XT3ROS9Ia
ZoEc9VYe42tt69GAWjJIQGdTzDd03Q4K2FnZMpKyy6f470CkHrmvBEe0+SaaHrjd
w+l25PXmMP7axrd29Jn2ez9xzDgy//5v67oInMCjNIyDp/aTizRzABQyCVFzf2La
8kpqBLKXysxSVx7UYHG4XflfaZcBkAgR5Gn/cazX06W5Tsii25R6Fv7T9/p5/a1E
0Cu5/UtozijjMD8FDN3Hg7FbSDYtNNBJn9GISM4gxUm1CLpfAU/DVbQtVIsyMAyS
WyoIWuiFgf/bN02QBSWo5FlCx0nO3L/bYKpq257xiTtP7kH7viqOzGoCyfRnYpnj
jj2EdlEshKZOFUnmDBqhfKdpPKYIwodZvQmxp95mfp5l9GmGh91Cewc9fHLo36mX
0DMd1T7bo8pbXjCv9ogvF6d4x+e0fF4jtzJSB+tbFzSs6KPTlaXSelh8m4g6pv5A
OakG0XC9A8HXRh+fpKydHAUTeXS6trA/Xfqj3+j9OSpFg95+3iunsaOPOMmECkEt
PnMaG5aqKSkaVqnwAZuq1vYrmfT8mqVAdpE3XwQ2n0mtbbyabDgHIRzOAr3z/h2j
VhzfTcmtAp+5Fb/t0lVXhs7I4I5Pe9YqUZEl5DA68JCq/+fWUwQt6MLpO4K5vW/y
1JKPEL+yDuMWi16pOqfKKBEL1uXU1MZ/HOd/BbyLIC+pzbv8iVxd6O+VFEDVzclW
fUe+BpQjXcMLnSSS/S9yfHZm8mFLuJn6eiKDqJVtku35d4uNRSMUIDI0Cro4Xbea
JZXmFk5vljnmggbp4YBU2H1/M2u1KMRGfO7sRAPU3QoOp1KSPOcxe4ptE8rSIjUl
0VWZOY3AM7bCMo+YcAGSPgne3faUsaGhBRKxl/tN7koMoKtpa3AVO6mwktLZS8ld
ryhwhMXpYSbu6PcRNokQZsNrLq4+l70H0Dp2Z0Kq7QvqNhiA0cmB/7Pm8FHD264h
cx0hVoXBEvvphg4p9ATeIXkAgpE7KZfOOwIz7p3MtW2YdXeK+cWl9nNf1IyjxDxA
picL4exk/vXovlkNKe6yu2e0idFg9Bz3rT9uN+jG0GLm/X70XAUzfXNkWaP5XshP
5JCT+p/Bp0qrAkXCqatB0pO6jThebBialTSHI5n8oNpecycSxnE/+PUF7GNziaRV
K2EJpNws+YYu3mYdNnJDFbgYfkLwR6K82pXdYvZYTB2ohiPS2bdUG2FedUOc7i7f
jM6QteuEthZkmvs7ktkijajJ/ziiIi+wDH7MNOAtXf1kFusVsbapADucLbMo6bIM
U2R6vVqLEkOCMS4i343cVbd96lPgQProGDFN+eTT5vLVJ2Zqwf6k5LQNagEfrAjA
1k72VIMBtxvJn5MctAE9BNMI1Uy54NgMOt2/Dj2RcLLi3hPDmq1SYD3AGT0ub1pB
fGKwWvyCFlBTopHILVW4ctPKivKUgELK6qS2M/A/1uF2kUL5FT85ajVgx3LJN8YJ
uONPoRTfHZFW027Vup9BrlQMSPIikIvbpUnn4LgItlFITLKO5VEWT4irISqWr5qt
F5rOL0X3WoVlOYGqIfEJ2rzsgxIqdJGtddBkV4Bouv7kr7FehnBriG7I6RrEvCXS
+t0bP2/ejaFh4bv63GXJea4U44UuEuD3d/VBh3hfx9rA5qgQB0BeIRAgt/o0Vs0x
ZuMVEcjjGBsVEW5BukqtNmeK28C/yO4A+ov9bAYALbw+8TfDC9uWhOlGy1Gf9TVX
0CnX7BbLXaWY45MJznkmjsbwKBOtt5nQ35jNesP3i5oJa/8a0Vy2tTqP99yJ1es2
joHh6RinZAoJd2lb8egOPwnEqpopBG/gS+dFIV8zdvm+z8dLOuNbWpSm7DV9KRw6
C2fDojKli4Bbn7xRNbJcZ0r0v73A3jXS9UGMaGouGJA6RSULoVUwIKVBMdjm/68S
t8f+wNIcI6bbE9fxDv3jj0ZBRmx41zv3coTNXaD0fKuJrQ0Fgsl7sGJGVuqXXUd3
8oWi1OheadyyiRNKj7HLcVxp6zRT6nR7p15Loid4VUxEfAOcQl53Ag0dSiRG7J/B
wq+KoM7Lhrl77LA1WS8ZqkZCEcVkmi+m5+b0zyMnEcEfmWfZoxm+7TU6DRdQTNGM
X+Y7mYMPxiXiWlu0e6DdFd0/AtdOVd/VMhp2emFZ7GlQCcIpkApWGv2M2lXxqFek
w7qZHQSs/ldq4Wiu+mx+gQNrHQ57l+bgW/CwyjmO04nhj/10FvPStXQiZ/2bLkrO
G/nVoPrRdaK/5dfORuaPNZ0UMLpotdKkMUVIgKLZiZFbM0KPlhc0lH5aSZ06uLUz
cKLwz5Y8JBsxIw9Hz2V0zbtdo3Whxywgh9cwT2AXrgYsSYz1JEhmmdN1VjT0fFXO
cZLEP3USDgc2BEDmRQCu2S4nK8aiiNdDCZIFZjsclLahaoQwv40wKoDu4kLKFjqG
NTI0mOBrAlXbi6xFzkz8vG+vZIZHQZZ3aJmAPCtglWpw4CRkLcoxlxNV9hBkk/dO
EXVYpBPH60bzxfAqx1OKrT80bVHh/irwOlbAqxvZx3xyvNgT2ktBdB+yQOtAUilj
ssyXuqx3HoAb6tUF1Jm6YVZ23va+OYZLRQRn3xwfXLdJHWM97ObbaPLMuwhGMEZ+
4jcl14KEtEAGk3HVH36wMJbsAGt4vixbW4ezsO8Z9Djodf/kqsrIYfhERet9gVGC
oLeUuUvkpymYbvPTtdMgSr3shnJBq3LBaTjxVkbujE3FH3nOj9dv4zBQbSv5BuJc
`protect END_PROTECTED
