`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w2j3ApAi8H9MhYiLs9/JaFkaM0jnvu4cM4mNCOCHMVmGoYRGell4Ll5LRt1qAmMQ
EBeYWdwGoQB1TFsarbpf1kBZ0CrOmJwDboFC9JiAvtdKZqsf+nbbmqRmNbr3a/mL
px3jXSAEa3ddddIZfzkWUaClUqTHFzDX5Js7Cb0/mr7qjqd8xJgl4c2MLmBxRKq9
qmTNVMep34aRjSHTUacO32KjuzCAATaoFTJyhlDFW6z2Im7Edhc7EHVndQSEqysd
yVNe3bN+TTnLXMt334wnUyCGTHCeBfUCZ3olT1m9k5SomCGGOJ2GCG8jgpVSbGwP
VmPQBtlIpJDfH6DUdQycxehXqnioHFrmbs1b/Rth0Ks32YSWZ95hDta/gJYO6dGq
zuDOOsKHAUYBxK20jKRQCQ==
`protect END_PROTECTED
