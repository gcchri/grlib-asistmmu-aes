`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2AG8RsRJzQRZAvrL+0hXWm6NdoA46aGFW0K8k3DgF8ZFqVHhs9Gzdw/bl5NMopEg
BRUUxgIQgAXg8hkZNH960678IvqCSunedOzXUr+H+GZYPuLqERjyr7A73jxcUkXh
6plXt7dSuQuRuFdTPcyoEJE07SpNDlx2Tbyrgfhdb22V3H7+2eeHJtCSESTQ62LA
diJYZDqEfl5VAwBnXaZpxu66oswAbV4O9ezql3SDwFKRUHE8Fm7rSq52L3M7gCDx
iPkpY0r5ChFvs1D0iGMGiveEJfYQr70AzxkpZOpMICR7wMsn+jdsSTMGKEhZtj87
eRsk7frF7ktp+hgIqeU/oqrRQrxKUE51jKLlL9I0NJ9NjXax4eFSY/clIZebUGPu
`protect END_PROTECTED
