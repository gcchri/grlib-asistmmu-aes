`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9K0h/S0jM5gYlslPEtPOkErjWPKr00o7bzIwYh9i+vJT4n+Gw/UbUU61/C0NR71q
ESeSfzvx9gwSJOhr9MvXqgAMXfWOuFnLuaGkGABeLKiLK91nB/RofWPrq1KX1fe/
vf1qwKc9mdovVZywW5jXA+TtqSsOv204PsvKwR0iwfyZTVwVxWakk7RQJkvYiPxl
jW9nJvG0W5r2PxZELo0hEuxEV4p8SOENT67uN6ySoRtLAvsqiNVoVqZu+luUWMln
p3SaGTNdtooossygm0+E9rUJeY5fgAxQ+6J5cF1EnYXREg9lPZuUiPidk46je5Rx
MbjyTuNJC+2rH0pxqvgvGncX5C65QVzqCo99ZB0Ne0nXPnUgoSWHDGEEQVX5nrJt
KyDr/ne453wofTorivzyUEla4z1TOUXwp+to1/IekHE=
`protect END_PROTECTED
