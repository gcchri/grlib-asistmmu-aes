`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBgnw6dRYil2n1juLmtaSBddeiS0UnDKEVxXTqxK/jlOUnqewvTGxhI5FOZhkUiG
CH2lqsgex7bC8Q7Is6Og+UV8W6/y4yWPVPx9MfkbmW3WYq7Labu12WD4G9aen05H
8h8rf7eL/1lZCWXEGCe4pl/ngHZEBD4d9RrXtLO+IM7PMr8dzAJI7xUStNBRO0TX
02H7WF0GHJrk3i27S1tx7FHXBEr0iPEbSntw4i+NNRjx/XtHo8rrIzwSrya33W6b
fi/ty2TvfD1S2lZTsRVlydrJe47iMdTWaZCvW9NdwIBgv7C6coMSaZVvHVtexkQ/
j5sN8yvff4G1KXBWRGAST7ASQ8qmsNMwkKrY5q5PybJtwiZpZobCg8G2AJ2U3Yic
gHb1oWqXb0om1RoSbMYcAA==
`protect END_PROTECTED
