`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCe8V0xfGMN2J726H7+dDA8UOSLsNh1nQDkN+UxgeBysakpqyfKa+p8eO3ZX34Bt
YeW4Ma/C7pFCWaJUDhVs9a2udaote/TheaVlsaHkjKRMvWhGd8K+ttrAWFy90RF9
2FH/oJxCF2qZzeDxRUCSGGdfD2OSvTBi80oM74e8bLfA3nofO+lLLHIovxwM8AUU
23x5TuRRYQZxjta8LFEeiJl+z1xbddsoLKgQtSfLOJjt++SnyPrTEf43+a5EiERk
JuctYq3XoCoelsmIxumOAcRbdhPtHRz0xfAP+lkSngauJ92Rv32EwDjbZI1ZVPfn
PioKYctpBMCmZINl/TEHqhntCVeIvkVEaxRBpxO6nMGLAJCzs7XVuUm7/PUSqf+5
L5aQhuK5BOIISL/S8xrELGmxTDhOYzDKQM7QVw6BJKeeB0u8Aq+l9N7wXfSc+5qR
yuOWCvjoERuDu3kwjAahIofi3kiaVv/mVeIcQXaGyj2/sXfUrfisAEBq32WbKpDA
a4upI5cNeccyLOZjGWhsqxswh7oxEI9h91yVddgHQUDMVKtiPOh0ynbskrLIjeaI
Upwf1jR9W7jtZHBQEI99zc0nIga8DK+OWrni6SGbuHfaaAihrOy1sMQoEnWwx1og
KMB0gcc6vSAR7WFUkZvFyywslAC4/yAv6Dos3uRxmX0=
`protect END_PROTECTED
