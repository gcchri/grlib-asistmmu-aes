`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dK1TH28JKS9N902Idwb/z+4+ku9FPIm2jjufFvrYBVMVZNWvssG5eqZnBfliBiWZ
PRNb9zKnL139DjE+TpqRMFUxmZ84IfJkSiPrbcT4Hpyg/R9a6IR8WGPjGQINJ9c9
oP9MXyYRVBNpCJSCM5qIFuYasQR7zhsi06m8znyxzsA4boc11hCBarmPihFZYCvS
btI6TmqRhygfZmlNy8QnLDglWcgCPQgxgVLUZxhk0YSkgVE8jLhkOkXwkbqIL842
prFVKN7yqiBOSKHkc1S4tDKFvad8wBC3q5AxJxvaEbhORfTwvx85meZvJQJR61Bv
6+txfHtVrj+iTFWDxk95QzdukbTLFbwgeE3k+0IZKfMMLEFivPC1VCiGFDeNfuGi
h8YAL50EmGc0WOlYcc9HIBDp/zcLghaGL7ThyXCkSTJlG91+Qpb8Snr0YnT1pB+c
RU40ZfHFWCdKQnkd1j551qy0cq6KHRFWJImTOSBrrbURjDnijDT9DsF8AYUARDlH
X4Vd+H2j58o9vS0cYMHp79b+z6aawpRazs66+1ILltkCFq8svlC1QfUBV8g8m90G
kqGYGLIS449Of4BsC2GpQKxZdKcpmb+vY337t5/qbTbvvozU7AAcaNvu2dpzZC7R
eH146zQKMyqVdkB3NhWZfjYdQ1NRwYZU4zKqBANpmtAEdfTK1RRBMiMp9KhUXstb
n1yqYrn85wFqVnT5oVEeuCCy7G3fbrt5s/FX9q0Vmz582zbuTTWyYIDkmnKQ2e75
rrSAHScS+Lnh7w76tSTPT+UetTXF9jUc6oPhq6uARbzcqB0+QeF/IvanCNe3a/dd
yJTGWWzEG03kEmmSt4iLcw==
`protect END_PROTECTED
