`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6nvuAdMyMUK9pyIirSow9ASy9Mtz4x+UGgAM2tUZ/a8aucM4tH1kDfQWI93Myv0
r8DAcelNnLgR4JIZpJhEfTpCHErpeYDrC+Hd7wd5GyaIKZGtkqRXoVlErJlUvZB+
7nsS0+R76R4Ym9zz1GnGGAWSChhD8kqbb4sHWnwgS/1epcS+K670MneTjOAWSDhW
bOE+7AxYZPjvTSkMwSdY+LV2cX7XBR3UacWDwUOwHu9kIsMC0GcWLbT7eITn+hjz
ZRTGzifZE0I/dG72RIugl8HRqeJSEuVWpmPBiYCIyaAkKEPFNnsxRvZImEZDBhLp
K86eMVi3UxWOpCpTtCNe+X8G4KZQzhVbxxsOi5BEcLX0mjiVFGtPAgdq+LyxlLTa
JzVMV3+21X+VUmLDWz3MzTFMooDha8855PgYk9wwdPuuOgBCnU1Ys1Acfik+W09l
7VntPFBjmi/eyal7B+H6I2ZVtfi5Aw+Y60f2hw3mgo9rVV7QyY9BfDitRJqFnXow
`protect END_PROTECTED
