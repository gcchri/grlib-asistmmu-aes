`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X5P++ijHsYg4PgFhmHb49TqfANL049aPmlHxZsIdciXfceIQCcnlD3hmOm5neN6k
mQW1RHd2Pda7lEl04jHSuGuNc7XT+cOKATwQf3IuvBkNbSNus3wcZRaZD8OlEVY+
QNh/5P6kxany4iYYO1+mpYN4c6LEHQorHp7IkaGZtzd8GEVIG+kU/lGOSyEZ9z8e
Cu9pEx2UiVgRTaBKTR4V4bX+MbL991NW++wgjgUty2gb/IXQNuGvjinxJbs88E3j
evpN27l6yfhcD3fd3QGJa5p7eZXTmaUVgMq0PeWSXGjsTHJanFOq4fR15VNrvDB3
GW3AfZ436G9xjpCw1hPLAH5K3KZKZqq4v3I/sGVYPvio+0/8mh9JIZ3qdqM1UDm1
BIAnlSPlVZMjaMq+CisD9ZC6K6XP1xxMO5WwYNKkXYRRdY+Jx8fhXkicWGiyrzxz
abpEhjBXftJXTShRwiAUlMZxVpIcgd1wMKPlC9Gi5J8HPdKxm9aiIOmM2IME+q4p
cE3gincsgOUdW1URrm/6qg3G+eGsquuUbkTOAWu9DWMjr+Hx5F+2CwoRkUVr7STh
`protect END_PROTECTED
