`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J28zzGa5o9QIVXQ2B7Hsym2uxiiT6ipGXxIgeNM3bwx+bWryQPtmRnQq2RJc6N4A
kr+HWC/i0FQUtsbqSGNoCSVTVMMUnlAKv72kYa2ms76/ozrcoK5sYYSzBa2jwtue
o3oigDDJj+zjN3MDN+3+ZIzzF3vZvCpMy6T5wvJCSDdFc8cFXzSaTqRbqSlQVcB5
JeEiZvbr0L9kPtm4m+k1y7B15fyRN71jAiPFvJRBlBWPmTQ6Rxw6DKfPCDYo/kl6
BJ67xiy6wG81tNezZms7ssxPLgTBpVYpmPEL++kmefbYTHeWHxzaKLQwytGUNKk3
3noNueNyp9Dp8rFDtDWn77okpK65bAkN2kZbmfvzSMmg+c11vgWkmrfT1F/ZQHKU
H8mO+Ose73Sz//JgOij4ZKToh5OY743zLSnnskfPQ0NI9F91w9LDPQjJMDnZCKEN
XW4YX2gnsfnFYNGWGWjlQ6C3GFU1O9o7tJJuOqdfNP97Ok6ls9goX4ADJn84KI1G
PfqF5UW4e2gt8x9Z/mt4fc+IQD59RcD5PyPnYgYEEPdqMqyRRyY3ZSdtbivRwr9U
ZXGH/VOBy5rblaqY3V6C+8qSTBd3T22OgtMpfIvSq/QDceuvMlX/00W2+B36XhKy
4EGq+ioEmAPhBXl0qmuOkQ==
`protect END_PROTECTED
