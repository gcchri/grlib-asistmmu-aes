`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OTOaVja2C8bN2f8WwigEvTacu1MEe3EcoHTaK1zzQwWQBmpt8/AYCxyboyFUH+6J
UWYwWB7MQZov5Cci2jb8RuiIidrRDLhSZNYhpOn881aCE5+H4Z0wmPKU4phzzHaY
lHXPYuAsZwYkbNZHUIZg/yc3YCrR25eNrimxC2B/ypnRK24IXkUeNhNkhZDzXi71
GY6WlMLQ5RiLrLI2UopbM7jFZmn+8656lwIZocret6trVsEHZq3za0T1sGRHJEXm
yNVfqtq3DkGeRt9GFa/WpBarVYRJzyIGp55yLZn6woJKRtZc24m+1/x0FiYOWozv
mNNkemCgSKX6D0EhNKenLgeaw/oUUxEULb+PSOTLepX+sMbFYtg6FvK5Q2v6gPdT
aSxKKzljibh7UAwZO19BrtzZQAwTLnmUGy4RKbFXwWwx3bShr2RLh3fnhcx4FB3l
k8TAp9bTtIHXeLKR50cNTRS9aIuwIzYnKFmJejDsVFWj48sYf96hdEtDpEZ3MRFq
V9VxzkCeyr18pXItmsi6jfcSFi5GNHehwFqjjPfubk9S9MP4QoZz88wTNjJTIHlu
CSC9w9c1OqWYEPAwlNwH2A==
`protect END_PROTECTED
