`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vho43y2DKF5RzalQyS1mwz0c8/d4J21Lua9Gh1xxuur1SmCJjsF/I7FRJRJDXQD6
FiSTfWYT2HgtO+H4hPO0q+0/5ZIl+KJu/TIkrIBnArV9vOPEySWHLzgKZWnreW9f
3W4voib2kHZtBAPZHc6oEWkV2Y57FlopFVWTnw6zRDUGKqulFo+DLWLEW5Qhblxc
hKj7SBoVI1Uh9ttzZY/yFvgNUIT22pnk3Yh+5njLRzhRO4bXIzAVD48ky95zswsP
V0vqe6SDJujXtcGIfNs2pNyoVs3sDSOLOiFY09yUlwJi42irkLV5vs7EURB646R6
2wbC9u25AFH8lbfMkJbyPPfFDq6FEJ6aAff+kDWZpTo7qFKkJMzmiWPDsM7ieCTC
MIWY1S0/ht5qM0ASen+y6D8c3uw3zTjgpGyv5iGYFFI=
`protect END_PROTECTED
