`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3XaHEbdqXWv+uQv/Gq3JsfTER3d2va6LmbhmEH3y1uYwE3BcDGKJB9mdD1sHLe6
BiuhlQplelbYQryyWWSby0K3MBG0Ra+sbyrh+w54AKn3/h+fMU3cRbIYSdhCLL8S
Z3kBWGzi726a68GRMqehu7WYW/HZda7p5t1eRAFmUiZrKhWw8bSQXY43gimNmv+8
XHlOzjK97aMoaSVcFFcC73JFFWsKqEh7ZudPciIQsO1359f8w7RY6Y3rzrg49whP
`protect END_PROTECTED
