`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+sByU9YyP7Jj2QnYJW19XkxpDb1HLGAirqeE4IODEf2oFRUzMufGaAJVL/jaaj0Y
J92pe1BrvktvinieTxy9w0n0gFXE13RQ9kDAPYZ/KCsRl2Y9wsdlA8Lv5hKq/u0G
PKvkNGEvVI1EQZGKqnZ0UdVcnLMm1Z66yH0KDFQyDgfxSUohhm2MofDJ4cvex1gv
5VgyE2zlCsanOKpabTYvIJRzqvqP2grBC+/ivxp+naWUAHPsd/RDTdPGvh7bB4qj
BdxDiPalM6bQyx/g34vq6jUf+6YB6Y+H8K5pJ9oSC8jcKh53JVVCfUsRi6MdIvAi
eqN8qYWBPA6/n9PzDhaZSVwb5qhJWxUAB756Erg3BMQE9KGWTeo9WojOBCEN0lkr
wdEnu1maGaTDL49TXDbFRqvnVtFgscTQ5L8a3jmvSm8XpwRu7uM7GZorfblOtiMj
sOa1gX9lXPQu6KSz8Y+JyHpCOZAuvZeB176KBc5TygvbnGZp1GxmM6w0LbhKvV1b
evkYEt/AXTJmgpm06/JhIthe0uccmZZJ6m0xjb6vXKEpLNPLel7sThbpl9Ir6eAb
tpQLFl9ZUgmEMavQl70EjJWFA91gHmTVlusWwjkH9QfI0BaY2uFvAxSFBmY5yEbb
AhaZ68vdKpDVG2+Gu+b+D/E+hlPzj/QIB7IoSwIT0D8ZgbXbT/5y/TZRjrGeCmLs
u2DHgUhE6938N2SOTF3sa19dNY0cft8EY/tFVQ4xmoiXJp4DA/uaLSh3boWhx3kX
M2HXuNZ3HGvZM6w/y+hHTn3LjJZHjLW9CDw58fSH8phcM45e3SRy9bYD2DUHmnL5
aTeqUp+T///hqjPzeEq/1l4t0EKXTjl3VnNubSKEYims/9hA0av8tPtOo+uYtfjU
i6LPPH90QBbieQZ+AnJ3Slmmxl1Je2UYX7Btgb0TXNbymm8QT8jLKea5Tf8P3Elj
xTpbxnkq8/vX7MlvP652F7QklVuX08fq8CNznYX3DgsPOiISOTEOJAL8ZEkqhKSa
TGfRjU1dWd5j2CefpihP9S1g1qsivtJotsfUoHrNGF5qhyPZfBd9sjRuiL5MWXB+
EaTqNIm+MdOvQaP+T2IRZCRJaqzRib+Lfd25oGG9HNE03zehiXfPlNqOVwoPUCOT
zQSy7sldqqQjhCX1cwsX/+FBY4ilJNKqFEbvY1/ABpWzi2ULbw9H3vWMHLO2xeDm
ZB+fAl721kP35UmHfv/bre+ecS2UqFDCXyQiG5/2KFBJgNP1y1nredXRhiv9lU4e
lm9xKyNkz3raFWady95zO/fJu76zlzf6wvppcK3huk+5g2Y48xHWf2GPpweqtK07
R/aIQz4vSBSPOtffYMhwVXBv4jZqiCdgs81lQuT9Qo32xb+VURjr9T8+7iWHWPEn
dAnY/ez4lFvv+p2oYzjV1/E7NtEdNVPTIMbBryUfJxs13nx9sHNzY1wDrIlLv81R
dw7+hjTXN6gz1BKEN6ugwY10gA05Z5+jYat7MFmkkaHc9KTfusDi0oGOO9aD/0AX
NIwcor9Pj44saKB7LiAH/DLZjkMw9VIi8VyGcGeGCRX2wsqh0kGyr4aHi7nXtr98
o3Op7NpT7yKCLZBFtru6lcqxBWPZkBbv9BUWli7QpsbrCUBkqsCBJ1DRvtkz7irY
2Ry/SrN2WF7EZLHz2b4whwRmAnFEbo1XLzl4sOaVkT29HiHwPW0vQS6sJheuXvHH
BAiMrZksf6KGF07RaesiS9BnDn3ST3dnVnuKYJbKcMFGJb6ycVaA+89OeHHlCi4X
tIX86bWkfc1XPdmIQV2zFBm0Q7dVmZJSPYpnEY/0vHYOpgbsJV3zfO9yRAKvUKqR
3FET9kaay0L9GejUVkyA0zbHhkbVNy8gOclwQG+/burAIujSNYkxmvkZrrqDQtSW
EonYqKKzlzajl0h3dVtE2qy/eyFYLUWG0gIFAm+/q906vH+SHZhauKHQyBx2Xyjc
U0IooLN1NOqziItBOCY24dGOXPt/A97aKmNuCTS0UdQQNZHbayH+usLooGpQwr0G
Fz/3IjtMfHHgfOsDTBH8ZFNS6GuAzf9MPIUrqqI+QyPHrs58u+qPySo0TyyzDzj3
ytPi8JPhxkwk/HsRx4jB55Tt2ehpIEHeMe87inDfVpZlRL7rvuzeOzmVyGmbCh62
Aa6ezrrM0JDEyc8LEHhe4yZ6a3ACW1vd5Ij6EgY/g5WHBq1XPbI2JPoiV1OtY2KM
9TnDx/4W7JPaO7fry7GYQ3Bds+tqs9qWyzqCO+JpNeOJFM5fjaPMVhHjOfeMrwxU
bhsf2HC4hS14j8d0CiDa7MVWpdEmEu542Vhdizu698vP88zLPIJxvol1Q7nnF4g0
NojLPzoFI+42oLMtFUAgucL8tRKDQ9fqlpZhV7AlScPo6EJu4dSvdFdp5bsS88zz
OeWORXPv9vZIlCFR2Ji9x33VKzn8TWe1ocmx0mmzdUpIlDvhZvmKBdAe0ta47yR4
6PrGJV8DJJpl83iwPGmIyw==
`protect END_PROTECTED
