`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AQgbQYjRACVoCma+yqk8Rd6dwPPcApDS6qCoMWZcobvgVNVvKNDcr0hvnhKLyfEi
F7WboDAjIycjJ2BvI81HL1GO3cYq36ujNuPojrJg2yEKi+4bbbWpCZ7uv/ejPzne
wTXO5gLPvn1RrFUkRUAHTcUZs/JaEuP99kk6M+d/7pvkguGhunc2lP/cIWV3mNQA
WataPTc45ezHZhQ2ORXxUCje9vMOk412KJnbaDdUxDZNJCP8lQVFnscRUj5I09KB
/n1Dwi/5RqBWQqRJaWeUaMgPExZDunmtQMu3GjMqFGagmM4sKI3G5kWO6JKVTpih
lw1MmiDULoqpTiJXtAfjiK2LerYjVAb/mX55FWnmEO2ChU59mPLwsUksmOUxqjTw
Mlc65h3WkHGipQRCVHaSuMkrUhaGMNs5RAKm2qHX9VBMsxp3pRD2ypo/fRb+pfp9
1TLwDIevLxjok8CM2hrJqGQBR1KCSWk7tJny3WeZDu0=
`protect END_PROTECTED
