`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UbpLp8ladX1H7r/5FeLq3h1kEuMqBfQoneGGujqlFMIndB35Lz/r1RqcpSngFBVo
JPOXhQfzitbgpqFtGuzJaEEnl8+NY7n6IFtHc6UM1W0FTfIjq4zrJZzNCz4tDkG1
kiiCXM0JIKRFbesWwwhRU5HnvJj62K5panuzb7eIgZTVfMp5PzRCkWUnp6jCKLs2
NBRYQNtSQunaofLplZdJdkyiFzIo2Qho/vHjkMCHutDOhVj+hSQutfVoCu+b85Nf
5ib1D9z+aOG/yu78D/UzZbZPEHNb69FGIu98p2qYUc7/c7QOBLzaV5eXGIfaGi2m
k5vjxcpPKShI0DwBsJrIAeEJwiG3uYihz5aSzb0O5TS60ozIP79h04gvAp5WZ5Q1
4r7wB8sdThQmhV1n2A/fl5zmxQylwDsGGuh9IOZj/aKCZEG7kYeYwUIMTHYrCAsz
yRRb+ssNFF8X5WyCg+Q2+1piakhOwjtTcgMVLpx8+S0=
`protect END_PROTECTED
