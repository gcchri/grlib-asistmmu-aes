`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Ie5m4rCklBtNBbjTjX/duMGZwz+e5nwsUEnUyjq+6bG4fql4t+WVxbQH1V4Q6bN
wTIwFfVu0LY1u2ro5UM43N75P/pq3ZHEzQbPOhFXQPsKmTCUH6ZXon293R/WFOFO
wFO5V0eQaleibuYr8MZSoBWkYh6pQIrgbAH9sIMV8He7Zl4T6aQSFim5hbAwC0ut
rba2Sr2Q9rHL3zrCSU8W1hRRSpgaUkyMr8xoPTrpMXaM7XcLkTCg7V6G4qktbOR7
D2S5x15iG2H8eSNJY330sF0FU87zqFSPR7N52f5GxxlYEe+aSmo/ReVHjWE6P6kE
P3KgaOGytIxXn0RWwQJo5wiIFbGfF12nLWAYcBIZ/UMreAWdHitYlCsZAb7M67VN
hLhFFTbsSlzMqrQRPunNTZmsVamAvklL/K8kIBMDbeBuE672qBTNGpteFuXKb1tH
PeKxv5zkwvvljP86fK3r84waW6RpSRpf4wzr3/dpq0JMmsJjnM46Tt0hzPYdNNCh
AAvo8XGl4W0Pg8h3fZkFZU7VwuTR+Kgwdg31oEYVv9e2K+xnD/vdDi7SrI2S1Dqj
LufW90bePR9UEItgwQXGW+IGTJV2wtJKG5Z1QZ6IlqaLX4cZuyRhg7z2J1tUyjQO
jieDuxZEWT3pu6Pcy0e+Rv1HLlu6pIdDVOMdOVFkdls10TkYTMRJAbg2Q9FE/0i/
l7zY82p/PT18dV2fW0W/Q1y75duPMoOxT0z1chjmauxxQFkpmYoW4SFA+WS1sW5U
7cAOqYHqJd0b73Q5U2ziZazz/toddiv194kDyt3R3lR8nY6NDzDjkhsBHh+SYOss
IFwIH9vvOuK5Qll1khicNLNcJzbodtgLp/7xOb/2RLaklmFMHkDtUf5OdVZb8mbe
GMIQAa6moW4rlufSXXLMBRZLMYratFzxLXugFWliqAa1vbV362zcJZJw9j2pJfZK
2EAuFshMePR/9IfS+CYqDxctV7Pk16mfAMu+E7ZRu9d4ufqahm5fRzUNj/8WHegD
dfvawjE4qkIzJLOVy8VKzoVTnFVfnHBuRQT94vvHNXM7AuQdyon4ykN4agGshbch
H/7+syy9LyUiPpIZkR8wWXQeyAj4xQZwf0fXK72iZ3UE1E9GguDFQZO0RO3iKChz
zvBZsZ5fsiMzDHVB+gEmoxwdPxpbZ3Hlmh8xdRtXP1fxGhX1EspNKN3edLbXSxtF
vqukcs8WlHVFxtkrRD0cFmeIIhzcdG85mUUZOoGMIZX6YVRp6pOoNiCLts6nxpyT
rUasxL+JWFkwCSDgviD83H0HlEHKXq9CXlH+XSRNUfsjq919BmuxWlco4Oi2QZsW
7HtcmKpAoNG8L0pYNFv82KmnjlyPAByxBq5CajXLWwvBjS9zlaSFUx3gWuc1/VyI
cQ2+x0ZP/3bhCSRbf3cdjKybDC9r87NjS1zQsmhs+pJR3dYpWroPCFpxY0Z7mU13
ZMdfgW4kCodyrXuzvpTTJadwEUd4tumfId3QmL04psF4JtgAvc/cpeWcnTYF+jSK
rAMVFIYUVd6PWMsNlqjNnsbesCW6qbm5vGhiDN6D5n4buV2NrZOVoU7gkraVb4UR
ErO/hoEpgGJO7ntEzz5071hnFKHMkGWe2fx8Zigdny7xIb2QD6jvN2u7TumyZbNl
6XPsUrU1QPziTI3bCEdo3s3zy73GdSOSo/Tyz7oNsubrQCalmdwjwx7qteqyUc2v
ZC3dkk6LoRGXVYeCD7oAO7nrqjOgXF4Mgtr3G2eggYt7rQ8/iBjVZpQJuMcV6zeY
J6Ji7Co7tCl1IEEjCguSJLq+BapfV4ZL/TmoHw03EThPfukLoWFqAb+81eSzQqeT
4gv+nfXHnPSxnRvhQT7zOL2ZQfo1DoGFuZXuA1bO+9HvEDykXq/FwRswAv4RwevQ
8jN+GkgGjFiIgPh/Omqtd98yLZLa9O/MlT6Ut0x6sJurPe5t8BEWCKoBlyy0cztt
XioEthYJ6CKUb2ZVVQF5WqbNW8MCDlrG3ExHaymw3SB6+jHZDYnTySIkzswjoX3Z
jY7B+SRTsg9vUTFAXfLgXzzumt6sWqL3jNhTxKqcbCcPHl+0rKSx6MQW4SahgAHd
wPv2agS9HtqA7i2vsjWlNL1tqWByagqGrVBxTSbh4suFvjZL+LTVtEMZrmGpq111
YGNu4rS9XmXR6cpsJYEXgNYM5JcPbXQXHiMGpLx/2RWLv1fqwoBRGosSziwIgBUL
TJk1cEYPdZ4O8ZXvDQKfMQ1dxy5kv+LTumID0mdFJIhXowlh0QrpevRsoiG9i050
ysJMT9jTITZYtQTjodGuQCpVZ2EQymlfK3Mfgafcs1XsJrBhnr53wP3NiOHbaFMO
CmddRRSSLw2CvziPRG9J7k0NU6t8Mxu3M0emsHsgxMd/DhtDugc0K1uqRaV3CS2I
mjTq3V2TEhN+uUKr7gFGMOs7o4NJc+jHFMV6SfopZppGdKMdS9+YN40zgmo+of3Y
fO94UURad8haV60T27U16PCMBSP9qjV5gnEyDDirdGJcLKihqsdnBID0XjSKsoxo
qJWYA2ICZWuskyl+ghtECx6k1nunlqOWDQ9fCBuWa2a0g4SUljn5rxfehaCDEdEK
sspXOtW8g5ym/gFVojt2SViEr7wo82Ndn7VzATO1T1/EFPkWqn+Rb/PfaVzV0jl5
4C2zRa22FuqpFmc9OGZj1q3iU9xSp/6EarRQTER2Ks2PAvMYxZp3E4otIIc2oiqe
im8d+dvknMFk3zgFw8MvLPIbFKq8VwiCAQ+wHTdgPmwlBkg2khQ/M9RipVvvUJwM
FwDcMZiWpLZDMqwlFrgCPfAwThQ3bMs6zsBx9VfMESSnaMvCZ8AP/Q/luRM1auPQ
V9RXpe3I7j5jELvBTbSfB0fhqxtK1ZXuP41hAGxRpsRpuRIy4LAKUaPt6Z0u3wPy
EZEKsALV1WZx7VzwTcZ/McLwDnud2zvQCj58UsH94fMlnsEya/mFvc3tRf1+dOTJ
smd9iXZKuK9hnwUtBJYmqSa4zfJ0zvbwV2OqFHkqm5+HSujdKTtxfifUTOGMMV3W
cLmuCdZ6oTNSbvZD3i6s/Uldhg1n6o+n0PksNeZp6DiHtENa+eQxWFpx/UYwroCr
xPGe5RvJJK5EY3CW6SWy8YSYqjX42RtimWVBcqhCvwNWdZyWIGk9+MtaedfME95p
MErVnfV0GBtQb7/sGdF02zBc/mKJFjtvRLNxIBMZJUMxbhaFa6jKGof6oWOrmmOF
U60wfRsznPkgyqzrre+siLVV6ft2Wu+2GiQa9xAsCxvhKPiVstINwR9mLIx4+33k
lgVVoVAacLq4mp5Alqfw3A624txJ5KJasZtKGEg4Qlw+TOcrKmSB+nKGuEDv5qga
4ScI023y5ocnfa5GBHtmnaby9SSM0vbR7SrcPOVJfJPdVIGf41xuGS+kdtw0J4I3
xneViFRBcjUfcb09EoqZLDQUPQ7iDUbhMOGm920+ZnSizqEQOSsP2f8kZm+Z2Ttw
sOb68VbC8IC6jB+G8/IpMZTeAaSV8qLm2r20RVMbGZSBslVn1Y5+C7yAbWqMHbpQ
aYgIYDUmeHv9OkCFlubCWR+v+wXNLIpBcFEx04qaZx5nVGKnxga9aK6b23cMlmjV
bVJyFyw4bMb/bWeq7GZtbXFGfwezOUmqvmK3j9DxnzN7iBlAej1CY1gOJGM4pGtf
vkHki91yJLpzdBFS15YPzXZkMkx0PWXmB7GyoNBvvy3QVyZIbwMrO4zolE6WVv5C
gNegk/GkHW72P7JHZuGMrDH3AKCylLZgjKWGPW9ABCcYZP3AWhn3iRsDWgzWcuyp
Fj9jExrA6Jt5c9m8zF9+psi5X+GVtYQ5KstG187fO2TCg65muZpTW1a4I6NsOs1s
g+9IpQrAN3mwGa77GF6a7G2DtvCbV1wDVRpIM0wAJi4NX/Fh2ib24HvWEW8AbHDo
5EZO9HvhlJ19uVfjeF27XBvGoT9xSk32G0PR2x529RJjlcDbze+bHl/zVDUr6t4c
BlKrmR00Potx2pRWJhaD+FdV/+HSCPB5qOPjhPP60kc1a7lxjIhTW/HnVB5XCqIO
GscKGcbzJ7hMRLzjSXe2f3GhvhzTPYyv0MCKOIQ48TQXpXdfNl5XTKmMWrhRn0wE
BcfbHneZipTzum57yNiXzQSolBUXWAYYIwAvbpmubLGJknfkjYpEyNmLAaOn4ram
AfzK06/nR+OFdObVABR+VMvm3HU3dbc+6mtLsyEHJG7atPzUGGh579umMYXLAz1h
LlaBORQjjCpD4molv4ZiJENTVgydZfdYFMiJn0f+pmeTvnEwEMxP7QVDwgJOx4kW
DxS2GPpaCHeigiSuhykfW4hqJwOGWWsQubRGBR4dW8RerVMlF73YnNq+0GsDYkj2
++yhbJqEuckIYNhlUxSTQoyvYorAU3u6poEC1wAejYQd3Ui/5kTVCec/Swsum15Z
mcINxByStnApYlH8qwQAXJE/Q9D3Lp3+IkWCsE9tLBOvHmSLiOpDvOVhUaOkqeey
v8xRaXwPAQ0WWyzLE0GFXwrQeFEMXkTlwvI0igZA1K1pGorMboTarCyC1vzPMVfB
puw9s+4NKyTKc6VtgzXjxX/cRuMGed8FrEI6VQXQYUuCpw6QDUP/p8ZQHpX6p3CR
PcQe7rmNPl+wBJmIH+gXx8b3Gwiq7rnMuMLd5HXeV1KBc98YKldZsf3DGEjnt7cI
1uGZSvvCIJbHL+zZrD5E+/hF/LQ1ml+5zKgCM8DzQgaYpqmDOnCRMwChLXyWUiR3
MooHAmmxKsozeLyHS75CI2vGu49udzFooJZRYFVdc3isXHV6Npln4ielqvNkFGyA
a2MmbtvMRSgvxXDdfUGoKH1bVxJccdd9KTFkrgz1vNp0oLwo13XqNm8/W/W9KMe4
tppuBbjQQyUAzFIAoeU8dhdu46ioQlDWUPVoACVUdezwl3o9m8DuXge3BiSnFRBQ
Zs7+dOP7ZMP5j4sMKgTfu7SEKDzjDUGSzTCNaKxKAxLDmO6EO5nI+ilaPTi4JtJM
3QedgmvtyXkWbaPPKYDWiHSYVNewmy/GbrbjQQ5Xp0zTqefdnoxwEaQwhMDrV3FJ
k/RzULFnMjmDCvXgWH+MXkfm47zDsGkZkS3WcIcWtPRagBhrafk003UusEBGwtlX
zMXHJvv2kV726Q0TwsM4VqVnH6wr2qLIGdiCnI4r08Ny2HQ2wKtjctdP6GYuP8BI
5eE5sAM7CXMDo0VhtDgpcwwai3OMER9JUrIuBZxeN/lz9mj30N08iv/pnjoSHXlV
JuxMIy2IVieRpVCpvniw6XY4Dwz1N6zhXM11DpsEf+47ifqNrpQxUCUPDSVa/N2c
DmV7OqpbD/vI1+nD9b7prt41MuUCDzJEEnWb/iq/gIT7MUaP9+zCsON+q/tI//aW
TbL7Ogb1LuHTZM9uGpefkoGGDlJqhjGapbM2zZLh2MDahFNni3C1Vp3zhrWw2X49
lp8wxJUh2pfFWp89ybCH3puQAbI8niKyb03raE9xAmEpM0nnoQ1uLhZdtNNcVnj5
C55q9nVwyVnl1SYS4xTrLJwRRylhr89bm1Q9Y/+1ymVlU5gTOzqKQXE6KQ7Psqfi
0y+N/MAgZrsDTifX7arwDTthhqwEuoh8kwEJoXnwV5W46irtU4v8ZuW7iIMfg+JD
mpBjiQvV39Rb3cQPXZdzwBTqx9lS+7fLEg1l6zveOPpL6QuymL8q3g8Uv1c0+n5C
exAnlBqwxbihGdvZRLwRV2PZFVTVqg4eKV0zlHDCQ3a2ijsXuciBHhjT4ObCESgc
mOIhQkhfGlAFqmCLLcyT4oWjh0jwUxOFBAmfeWf6yWFsDBIO6GevnHnKQbCK8XEZ
li/ZXYMGbBa5SHs1VvbOA8nHjlN1PpPHHcodc64+Yn6yJ/flKaAeW6/e3AlZ5gcI
GGzrW2Hn+3fJ3Y5ALJYQnjRYInjObkljmwXjz9ZO3/nhftITfIdmq0CI1NIHdNZt
yvhCSUeXoj9cp2aJdHb1rb880yXD+Og84/uw3CpEsTGf6fJIz8zpfJ2rMxpBPaYt
qFFifAwRwvnGxKkzZ5FHz8P1TQWojuIFCJNVOJEjoL83jbA+fjXWBsjSAHDbH/2J
v+Z/i1nyYZHV14R1GlqJgK5sEILne7CbB37Zxi6AKw6vkG6Gz9M/eZGJH07HIJ5S
8UjjlpkC95aoBar4AF65xIDwHCTNUMIhBalxQEAbj3KlrVYwZyucs61VwRoHCMPg
QfLeVn7d4qSXKLUuPgv0M1tlK78Rgk7FDwa/HWylia0cY0iZYM0AH0YGuGOJ58A9
h3UChQwLZ5nGJ0aYa18cf27hyw4AdGyPi78AgE6smMGh8XlkDkQvhtRsk6rWUslt
FYdnMcM7TtOW3i1SMgcTxNcSJXD1mdmPCKF8I/Secr+fGxoVXKYQWDalWAnoUWBR
dGq/HOm6V1Usgj61wZZjOzA2v+17hTaRouJs1j5Vm+Gc0sB1j0i8dRyzx7GDcnjc
H8UoaPkZDXClRmdHmDSKOATfmWnY80kMU/OPFBMGdcOSvHIHIFnW9mXF//k26/oB
COwLn+otdfawAW7XMM9TPjEzld3lSQdrFgAYJKbGEnc=
`protect END_PROTECTED
