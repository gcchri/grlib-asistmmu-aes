`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRhfV4Dc8csPQd6StMLs1Om+Au/oRtfQ+wUF+wRuLZyatnPMbC50ZXn9pu2W0K4U
IMX0KpafA4QiTFSTd5t/7mwRTEC+6/d0LFkbz5tEly83txXR6AcgbxqdOuVr1ABB
e+6V6aVi3ybyWyhijisym9KKRSWUBwiRgH53CJsSt0VDyD3jkLe43AvWVV4j+nLN
TWKZvRd0+jIvi7I5y6M05NOoNWfLihILU1gS7Vq1tqK0ZXCB/+/Fi6DJ+5aAisKq
m4BkPrGgnqlVk1FxtM8ijbd9d5+k3L7puukJ6BmbP0HO49MxCR4aUku8ghulvjnc
23SJUGagzvEHI9+ppWwiLrZxBavVuXxGGqxtDq7h+IH6F6veX+eXPVophm75z0d3
Z9kUtF1209l3yqV9xpFI9KZWk6EUXDUDNab3O/6oqOJ5h/Bf1x2wQTF80P8j+QJW
eU7ZEe4HcJT3X7PVvaGLfpuPFrOMHZyMQXN1qo5Tw7yf7Pc6zATUwOlfMlsKMDQH
0X97cS/pncz7h+5ILcdLEeQyBTUGEmcu742tKlz2BxU2zjuX8zzDR27yFVauqH1n
9l8or6fIp0kRxGZwDfra+XSxIC3SGmjzQ7/8HEYV2h9fD/Ixd9ADq3farMNpLMoH
mJvpTQivSiV5fLT6cIuy0HxJhyNumcNcaawoPJFWM4SkWVt27+pX061iPxlMQCMd
zPFA8WApu6KGMgPLuntVXbQRkAxo2VX2VFNXonfYyChIvSieHgWhqQcGUhUHlqkO
i7lXwSiWD7U9uVzNgvYHQ1N0w8nX75MUZRgl1odQWo6+5d2EyNi7wt9eY7KYiplo
lA65HkrBGqmI1HikWelDSPTSnNFTu87A9D3asITG3t7WshPsfWaI+J0wRDKzAtB1
VyhIip6N7jSLUGKHooJw18srEMTs/OqE/JvYXNe6XivY7VBGzIA5iYPKk0bi8NKt
`protect END_PROTECTED
