`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wZp28AD5wcRP8G4D2mff0rb75/9iafaJYnK9r6JQjH6guzxiBTkGxVo1sFVyU5Hd
Hs08C3Cg+PbouTVfqN2j7LzTX8UHPZc7uhOlO70MpPhea9fTKcRdvAU5zLnLKE9T
yUU8h0q5FsOBC3MIQwthjiw50L1KGlPKxMQGp6hBaAxJovYOYH6pEokCaNQnFXGU
24X4aOCpRmJcyq/VHyv4DOD9xS/oRl/sVvpMJXhqBpqLfvhBjf23EgovSKZIezsz
J49LL/D+665lGa6dhaCFZ2JVSOqFFIC81OFhqHm2P8FAsAiKnLl0C+87a8CHc0Ia
zWcNGHBqb5/ciW0EGWP35XWYCxonSFdn/S7+57WJ6AGygvI1q4sfcCQUv1ehhRkz
9c4MQOZJgEs82ikJJncJdoqtOhvaupEBcuNkguYxHABTUaRRgZOU3/ubAJRmYvkQ
`protect END_PROTECTED
