`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EO9MKhdFlVqyegacFK1h/OGR7KWzlyglbUoyP8i4TWjwq2I84x+HDmRv+/kkwhXa
z9d2XMQ5x1jxlPyZ6PLLKSD68tgAxDBKYytPTMfhQKM4YBPB2bBg7mayb6HGf0uv
+MI52wsm7Knq+sKLVdQpg7wwJvodaRTr12n8GPtrzxYap6MaqHXSH+m5VxXjJ2hC
RHD0l0z7KPLYrG4IJs/784GJswmY6gOpnH2OQGilxvMgh7mx88Gei92iDzFbPolf
b3EkuCJHQrg/ARVE+OsFfb6kz+0PFfJ7hzVo7IZGI6VUb4u8gXmHZtHkMWjv3vk5
mZeKFJ5OE1SR7S/Y/afL6keuuLAU7eppzRSe5L5GxZn3cMDwGh/U5NCrR0yGrnA3
nhDY12ZM36qzvUjc+wP1pSSBPqxXM8my+gFmhoUws6yEMdMR3+qGXEiaOpzH2Shf
Yug7Bi0ARxFQs1xn/2KvFOTvCxSFpsAcvI3+EYCgfRZwDz+cNl2hcAGZ1W3R//5q
IIn2Vb0qdqcITls6jLxJuBJZhQUEiEyG2McakW1EqoTHFQXrHicUlh8o3jlxRny8
qauMV/1/rNjqz9AI7uavZtX2KdqcCFdL3DzXVbivDBycGdaeKfA09uwRqXcE584c
FNZ+m3dcKVlsI/eeXk9lzaZjqL5NCrii06zAW9LEltprFKPgEEsx1ucSrroYSorh
P2SKUfMod0cVapvW24xvFKZ+KjvpXDFKve7astXAxu8syqtIeR8V32lwuqCT9Yax
Tw2JxIYewKS4J0FNdOeM6l6KuQYm1dmcUrrTCMmmLFRZqUxTwodAk5swTIWQfMPv
UP/U9/y9tYQ0HHNvfr/uZY/m4Y0iVJsGngTvMzqOD32FQtUPNXtmhjBW1cFjdmid
htFbDpt3R51cA4hjyBLthy/B96VeYVflmcIir3ajHf3pP7QqtUkJXmND93SNQ3je
NTP8SfDy/xCYNP/zDnRu4MR18f30QPg//eZFPQD3MgplOXYPRduT7/QlMjKCZ8+m
1Qfho0ysFmAL/vkJ9wCwCnRdI6LteLdrGb1ynVHnD+P3bS7dcmfWHLBHhhuYogNS
Cx/7Y6IU5TYFHRvaBSZ/AfIOgBWeNO1re9Jkip6K5r7r5dlSOc18xT6a9RQdVeqy
TzXylT+CTJ1yhSUiRvwlda3Kwys7DSIUtffMiWgqUgo+ir3XbkgtNddunU//Xq+u
MAsEwImDnA89oIwV/ggX1PRwCvdOqAL9Ubkzw/3rpD7J21K5nRbhxTfnAHD0DUFP
iOaBphc9hrICBBqR4hVZbhSZWKcSdt3Sr7NzrF4UzGvFb4To5Ua8H16zt8wtmLPp
iuW+14N+y61umhjwY2zIWEGX48JgH6l0sJR4NUdWqtAlXp5CYBVt7a8k6IaQNEnZ
7q00RQyLtewXEEebrkRNsXe9trcsZO837KzVfIuNwJCT8RqrBPSqFa0JNuZOT80j
/nbXQtXQ9YqlvU95g3U7YtqRDFOKBrflhNWG8pzTdmFQN4tnAswyLS6RwsX1FQxF
TuEzUaV0wo1ah9LfNgHoSuBa5xyU2FIlTKppnV6uQGJBSNWCANXURvzChjhJLJuV
9Z9ruTihBG4nl2Hy2W+YJ2fzTK2i8az5vZF+ciGJaHmPrivkFKgENGkAgjioXDzY
V2B4NOulSsS2r+m0/7buRsblUldjop+X3rWpfll594If6gJkAvE0FtqPWKfpA/Qu
GoJHY4AI/VHv+UU5EqDcoZGtQZKMb5J7jov1rC4603IprCZ/9Hw+9V3Kw55JPQrf
52gOVJUc2adnXqJ5w8To28x6kHVEhne9y0Z/jbISfhRWGcrcjB9qhCti6BTWFFQM
aOO5LLjiFPiq3c5y4Qb4dp+JOJi3Hhp1cVBXvFvGgqeoIpByKJK+wu+TxFwVK4Hm
zQzb+rBxgiaPYhXyPykMEFS3CP6G6kPI4Ys1hEIuj08YdMdCIITiW0z60J5gnqLc
ow7ihJRkOrk6KY39sV9VsXHBjzcTdudh0l5McGYktF0ajTtZ/MQP4QhlkOgpsb8t
nzziDBq1875fDfEGBgeJW7WgmjNaiD+hcIGgfc+V1zmcIpG4BveYP6X5HXWUrikh
Zhsjhb7b14G7JskY49pOfE/5QO2orj269oRgwfJ71m+4DYIbHG4wm7VGbbTn9pqF
/pFyai/PFRln3o3vNSUx6+LHLj098XKOnV8n/Huv1aPsqyEHRpWYHe6dz1zawBxD
K2/uTdKWxQzHvmVWliHovlxk0C3JwQdlIQPgXBrqRkKX4f6GNs5LB5L3NVI9ALkW
4iisX8KIAMXNhv3uGBjA2kq9jq3iy4pXY6HplgQc3PlhkQaMOisI/Ew5P0CC3x/i
DHLx9h2hBL2xMHDRup/+CCfzjAoEWyzsUOosn0drj7pLO5dfs6WOCeEK4hAk8f9d
zAoKUWWZ8MH2em7+6woQln+rOpvk09oaIJvP+P5zmbJVjrcmc5PGKhFlC5TaAzCM
MS5trxxE6p+B0dC8B6qnNQUhjZPsnjjSUsIkKK4XdYcIbm89SqRoRg9xkmZExhtr
0dRH1fEeRGGmCSMKWkX8rjamO0iZIV2YuLiQ/qx+xHZc6yKSgbI6q0kS5ww5mHFy
n1treRbrtmhyS+1vZ2krD/Liw80mybq83ujWmirp/GpEi5TypyafJUR+alvNHZaN
zV8O5dr8N7ZoMdkcMdoiMj9CfLq9NJKbIHCSrFyCdGfbAxvEL3jFV2IcpYNIXS3/
hOJJVEBYaSQlaVMhz8gPNZIdqk97D8jt2ogtuQXVqfeMC7F8pflJ/Iw8x22oCpbT
jzQR73RHltj1MWDqEQ02NCRUwh1GJVY6R0sATJs1TPGPOcFfdCKWVJhPr4YvjnQL
ofT4bDolJTSBw8qEfK1q/dFJx/bIi2XAFE+vgmiEPDdhrkHgxSoUtKyYNUyB2P5z
Njwi6IKxsClSl2qDJ6a8om8a+JcVzoV7GZ47rc4KJvDgo9NASMMaMisPbKqzJOxO
G4dWkmEw7zcU7ige07j7TkwJHE+C1hOpXspd6f/kXftBTYIxg9TJXSg/FEFeElR5
EnK83os59RmCVaWTVw3c/zP/4c8pGWiSElm+9JyHJq5xMArEqhscIYqWhIGd9u/e
Ul/PuYXeD1L1HbNd9njORyhs+7mxyZf8Xbkly6+ZGULU9Eve0+xO3Q8Z0sHcUMDV
DJoMk4mrMCw9OQJkhI6fTTGOPGkIGxSLry3koTnyefAWsCXhYll1r7tlfztJjKMq
L3VBp8Jlua1OnCdtPMzoCSHju+pctxpmKMl5PqsLxkezW+x3vmN8C1ZH87KO89LY
PmNbMS5XKPrUf8i2ER6XxhrR6YGBqybfNwzK+SXXchmC1CXwzefo0WZdUqj0sUY+
0YoYykQuoH+RLxvrl1syyEDPmxPLjxB7mB2aDSRiWMTGGMUZ3D3tXzrzzBroyf39
j6aBgZf9S+5n0e9JtIDBqJfT4tOCL1Dc0FY1Cy5dXbn1xdZq0d+HKktIwyxGjNh1
hVzpheSkqVb//pky0pZ6nctMtOvaDKocxkLnj1LdO3J1PMkuH165EvlAbdMZliFN
HLUevhk+dNKV3kfTOscysoWJ4tYs4peZZH0inN5K5KnPZ37XqVtMGjlocHXLBzEq
kFtxyO5TjbpCl/erp5Khn83stEiZ31WvUXdiibIcldLZ3TF5m3TAgHauKkhpRfhC
OkfY3tyT6BRT5QXmDlwznmRGNnUmo8+PA1hSyVQfbQFGw3wCOijkbp78380IEHU7
zNFYETATeLq602iz2UuGJ1Tc9PIFwvj7RKaFiQvjJRyxbINlx6rbGTNQjQ5HvvRF
MFdHrbG1mITQjI4/+D3O8Kj+8pAyyyGilsjd8gyFk1Vowgv8TLLNg7DR/C4DlN/8
RLtSyWLRxP+sIe72TpBBN5+bGkk56DFsLMXfL34o0UjiBeDe+v4r2c/LvrKvAQaL
Udeq+NlMeT7ikk85e0GZ0kSD4WSgy/dQbckT0wKY3pOYHmUbJwuBgZVjiMNv+1ip
UkisGYb70t2bndawp+U4haIez0a/Y3GGEbqaEZp4kULbbvMRrXBN0JUAPWhEg0g/
T0lBmnu0wN6pW6mMN+xjccx9Pw7+ZFeCZF6u6l4CxsV+BqFCBthxX58EjSKDjZ4b
GCNqM8Ipuqm02bGCdVQLs0BR8D4AD0BRbPvvyKSebu77PAsR8Sg7t21mXZltIoo1
eeAbhM2CHYgw2scvfMq8Bn6zhcBo3HKY1GH4hwOB0bLsz1f45kKLsASrF9IU2TEo
zeefGq/biQ+pxMLBVTGkBGzYd6K+fUIGd+8vcrTMC9q6u5enP2LQsJv5JdTm2QLp
ZpaPZmO5TcQhVTSKUzIDcjFgE4mbyr8OkdrJWLj8wdk3uOKU0wBb5Ga9BzLc7Paf
tUjKud9K8MMAsihH6Dl3Fg6uAkZj+HypEJfDlpuzCtuikDUxxHcHVBOl/XZK6Qzv
vaJ17gMrd2iekc1iu+Ga1j4Yi6cXT9k1dPgbMa+JYH8K9+ZhkQTvPLBFF9DK3NmI
O7AwXP/pPn7uE47ZFZA0IaSPLDhpBAvZo3lma/UHkERUwBC+6+MmNXum4mokKvxs
AWoE+EXPlB1aIqOM/NYGVxwlWcC9d3axL9xZwb9kvwzKnDA5tWEoK7BMUya+IFZd
1ERQiGYhA9Cuu7dFpqePtxAaP9jS/4V/+9vhLtoWJmpFEahQwI7dX+aulZKC5V/V
Zt/K0L+KEBfe6rUMLMqulbqn/6FHWlpaAHEgQWXXKJdIp+uCFSmL0voWAUqU4kwD
7GhKOIntPxVxV4aNnA51yAIX3j+JH/vYYzn+UBjodH5wnLtgmZsYPL0lHkkTE57M
wghYGysxRcs0Z0Rc7cGKeD+5Le1HDhVWRnLMWneI7wbyu2R9IWDGtni/ZKseJnZF
ZPooUgO9IE3BDaKaNY1j0qIqDPM+NnMS58Y63S0wbUMQqNqbVWBRg/EQ3k5TVbGE
c3pJL2CZe7Ca6u9vXtrR0tamc3GhPJrpvmjdA7WuFKNTPgrl0kiaSLQkUqBIy0Uo
3c7olTJm3zkm2c4fyo4LaQ==
`protect END_PROTECTED
