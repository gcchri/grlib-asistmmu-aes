`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uko0h/NXXOU2NnrST3HbJcNDeaht22BAhVI5cbucrFsOvwcSKnUEkhJtTKsSYiAm
I5q2umdUb9IEdaxg0Yl2jhXJZoSw4u/ABuCe/3OmKW1yt12EDfpfAjcUihit5DpN
qdYQCfs4DJUaMd1owqHH1L/bMC/FsAYd7XRFC43WUZ+wy7G7JvAO6bJhKELTtrSe
g5/Qu/Jtl/sTIUjZIK98hiNnfzQz5rQLIqL0x2VoAskNgLwSsbhFVXJ0nDgJIncV
`protect END_PROTECTED
