`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gt0cz0K0FUJfK/mqHWQOCoxcr5T+6az21Kq+oPkQtCRu1Yx4jBBlhwYgI23gAZ0v
dYAqHOVVwsMJmDCb0ujPoHpMCDeA6i7ZdQRHTW/TpoJ9dJp3/Hqkj7BbsYxaaBSz
hBz3w+bFaIOq46xrEDtWVbGZW6MT54bqxiAAFG82uGC95I0s9V5QrfWXjXddU1q8
su2/za6sy4PoETN20l2FmNh74Ph5r8HFnvHOca5lLeZHDxudGndYSn1LgCbnHPm9
ZhjuXiLCyLC7JfhwZ+/lUOgKFUedd18vVzNRGW/JblBLCv+sEG4+ewYpfSaz6UpI
OCtfYbJMB7wIKs9h0RrhCp2mkB0sZ7zkRK3XxhKLXFpAApgpOWw5mReZ1Dp2/fLp
+WGzgHl+oyRfXwbU7NcCS9jZdiQfTek0A4GopvnLTtNk0Fs0OfpxipyWj7UYabv6
DCxTIEbOZiTenPUHd01KAguwD+Qq+3EVoT0H3IhJlA1zmYbMiAbByrQ9PnlKuJBp
3AO3Zb9Be/UgWSe9GL4EVukMihAqchOPqGKIRiy5mAU+9AOtsn7tbY3RyTi1pvEH
H0KYYmw/lVGvYqj9VFWLKw==
`protect END_PROTECTED
