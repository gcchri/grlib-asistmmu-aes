`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJjcXBxx/PPh+BYeiM9HJBpcDFvj4ZIf7Q0cXvOEzQjt1VRCvyzfLQh6OQANgRzG
knYjjbJup9T94yApQS+q7d0L27t8nhm4V/WtHu3DzM3Ybr2m/rza+VYT951bhUmH
wH8g5gnh/IdAsO28hCODT5PyU87GL1RGT3KXeuKPt93Q10o7zNkRHJpqGJY+Sfg+
RAvMwF40/PZzLRfRjFbunxIM9YgVFw93B5Baj7QG8gbSSalj3dChVdGSeNPU/WOS
Cck+UCogNli4cAR/dWJz0EPOfIAgQ3d51VsgvgyNwZQhsDn4IwY5dn2YBLwRc8Qx
Vk1sS4EY4LJc1TN6F2YXOdEyTuCC98D2lkOOnCuxclFnucr/XU9MR5pwxzuMuzmK
trRh/VCu5qi5aLG7cgAuUGOaJawpSVvMwd75t29R7JSz3vgEgauEO5leb6ySiQr8
oaBkxdwjwWSozVTM4yx5h50bxaW8S5+23fzdeii5aziJjKzLzoouNXSleeMl/IyB
0UtSCgrCYO9Phy/4h9Vp41wOuxL3NoXUfsdW++8vtzLspftuY/ZXUi4YR9XzBYq+
/gOmp4b5Q3KezOZI+kZDjbrIH48PSpp5taRsXewZ9V6Khc1kA9r7bQmpcVJJDzJG
bjiT+wA59nsHhpJ6jClk/bH6XkZD6c+buR3mQNnvua+PwlaFKAXRzd0hqdtQjVp3
ITqYveQx2B6/Jzv2EYslZT6XDAzvRcgD6R2v+zbrTJcj7/tecp6MlUBFp9hAKSZv
wE2+v/jFoqv7wVkvno8C7hcj5KSZav0DebkpOSKmlgxmXVeIavP2WZBmQr6dyNCD
UrZ8ZV5YqhlwPnV2cStmfowpG5mdV6W9WxprQnr8q2Ht79kpIbrqtggh4IPStbMo
FmF3he7SovWEWL+plM+RcnJ5Dndb6b9eemnz7ig4yLeW2GjRBkUDb8Pn1vDfvpPq
EtRe9ae+eUjKDVRLDbgIHw==
`protect END_PROTECTED
