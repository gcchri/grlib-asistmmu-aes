`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0TCj7aF2IMOgSKwS5mPLhXHY4By9X2vvMcS3wYYQdzsr7K8o9zSXuOJD/0MVzv6e
xpVQyXfBWHn6FUYNH2w0bE2FrCz9JSQnHo1XDt5+pSb/4+EJ/n9WpzxOaVpmVjeq
gHmpW9u5NOD2R1+mq5n+tN7BUXQgzo98gvemTDcjPytzfucD8NY31/1YS03675Xz
P5N1AycQW8wOAxBlqoWTDJi3LR3ifP++EUvFXb3fqoyJ5mV6MA0qVcWFZ10pHBwf
GEoAVHY+h0yslhRVmG6nF/RsSEuYXx01tstoFsPm8jynPT2Ix6LloRbQrhZnunGE
RvjHIZ0XE5+B2DgqVWEYMd2Jywzj/jNj9iLKnbPKNWFo23muRRCKYfTGsy0QmPpO
AoXBZYMhca40DWEyBxKFbg==
`protect END_PROTECTED
