`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+w6B8Kg6bTfzzQkoxvyLvw8j1W+DJnaaDbdho/nMxNaNbBOIGHC1Sif5e6OzkQl
jwT3Nn4lJs8bTiqWv6a2QoKNTezNExGjchYRSTZANMC1M5S2mMBUXg5oV1RAhPhI
6Wiq13e4wdwWOQK7MWUgf6kup2Yqbv4vUsRd4H3Z24ZfDh43HzvmA9TBYJNICXWA
+bCEXp0VJIc2StRH/QsIsF8ubIEjxX5QHW0CHqu59DVYjoBxvS3W5Mt/gSP4Qif3
gBS6UpSE5y4inAdjMkCL79wNrbfqu+BSJbEfDeKzFhsiX2cTc8hQkhc4s1xBE15o
XFgx8Z8ga4+0xfU1qCcdNTXBNscbUBKWyGWzcT5ZtrzWXmuTPl5HUI9PMYfG4JVf
ZDJ6LCt6g3E2DFXy1+L3hF2VhJA58FOC9hlXaEv/nxA+GAK02F8ylec/jRJgu8P4
wZwKy5bpTiVm+gjATiIAEBl4C9LAJBpEjK3QPQypebGA6g9HPAkcUZ37bxWVt5lz
ImCkbwF1bTyIE5+u9+HnXBSQjqj17w/w7CLBDpvhukylDpnHt8DoKdwT1o3pFpfa
5HD14X8I/nVVNGrQQ89urCI8qa+IXC46pVLV6AGeTBe4lR/E/+f5wybTBs3I3eaQ
MJbJXNK7nmuakQpSFJHGXlGNIelMNhGEtytNCabvP4BNJI+/t1Xg3H+C2G6aby+b
cX06Zksyoo52J2jjkZAeLjXvHHicYdGi4p6VMNsOp35urKZfbWSeow2jzJQGs+Wl
`protect END_PROTECTED
