`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rmkcI+izJzOG7u/7LcpY/SxcDBpkGF/eVZfGh0rF2pu2nCp9Va5QvEVdgEk0uDs
/ngir6+3TDQNFTrKwO6ysM/KgmMisJbTe+a2yrOdDp0ZWKIWQkgidWXIbTiPgTnB
9fng3c2FLM+chSBZLh+47Dh24ATyyTMUlQqGOYhDIS+81R+rxAmh7PMNAhtIU0h/
mNMpUOAq+Hm8hshScx55sUGZafpBviycQ43HqvdnuApGlVSq9e7XUsquFmV82TBX
Bad59hGIx2JUB25mt460837etNyJ0A7jgrUnNaxSWY03TTMpqAc6UOlHNUisX5rr
SdNKLZBJFc9yNJAooLnRxOZukRAufOgBUQDZ91Oij2pBbePIwvH4QTKw3+tHbbjF
uDdknYCC8u9ei5rf+8x/zxd7dj38W8IdcAsnXzuCRE3JYM4zSTBe795HZrY7jY/G
8l75PpEaNJRDJZHMymhj1AGvp4gEGJXfwGu9rs1LFpGI4bGYiKhMgEto8kVhzRGH
jPz5cyBN8WQRPs3801bqWJ/GtRPcxNRZZA1SMpXu8VvF9VFbY8hJL64UfMWV++RF
qQhyLnB1i0uxE3L2+W05uoTWejpPxz6z/Ae+vpRh31c4QPG0ni48buwe2IjtpTya
GniE4UXd4GxMSZ7db7+zmkHz4et/5m4AImhPbO6ckBbulmo4AIGl6hrQDxDvHYqa
x1ofbRnuhCv7TfqjCkH++o3bCMIAShZFw1tVstM6lcNqG898GDMKhiIkpR06kVnq
CqsafDFHoNVwwHid/SWiTw+PVQ1idno1rKFCFT2pS8B7TAWjO5FIIWDIm8NKF4M3
m5JLoEJKeu7d4ZsP/TgSSmY36s9bB+V4KVkNu8CjCjn4YrNmSEaovaVN5bW4dVOI
zE+BYbR1wyLdzTzUHcPm41Y2M7mgz4SAkhoQ1OuxcpvV4nRUIWVca5sCrtmn9wG7
CIFFKxL9LVKoo8tJv961qse6+sj/eDzt2Mdcgo2/zA61YZOAUZ8OXjYYVczwMrGj
9RXZ2hTTrVSRAvUKSYaALX236DbEfQVDnWd2ihAPKo3RVmWpDyl0q9kgOx2Nm7xe
sR6tlBqBXRzF2Qdd4+Z0ORcHSNKWyhpej16zL88j+sT23wPUbw7SOQSFGZyMKZ+4
yMl5CbFXH87VnbGVJkwylMHUOcv7SehsOhppr5VCB5X0apYbuacrpVT4p+v1LR4R
VKBaqdiFKCFkLMUVMPubYpzVknXQKhiuAM4ywzAcxVftM60wVZ3ndlZfmIT/1EeY
l5nxf5eRx+2WHabG8yP9My/zDr3HNBb0LLR7+DbKILs1p3bdf8IlX6S8hgsVxMSz
BDyj9YEpm194dY3pJa909wLz3efy9xl89Qdon6cRJnBoJKHc5DauBchkykjYJMff
Zo4mXDo3MQJ1CQxlU8EssbjMgJHfs0Z8BeCfiGPX+awmtFL0GLtb0NwWENW0sd8r
FL5ggLZfsazaet4nmEUVW7j4oX8CC/AIaQfMJ4bIlyYG8VtJK1+sWWDjP5SJXMhK
L9rAHmlJBksqEIXtKqFju+kK84YumA/EavvcxjKP8bxbdPAx/Nw07gtEt9g9X0+M
zHGZwrTKXBU+C2peGkoE/XEvhnef3GjlpCmiYCLEWt8Ds0sfJMlueOWUyBck7E0I
WHOmH8fiWny081DtTihCSbYMR1zk8VqRDub6cLH2Fc3hFBpHaeW6UyYS8XfLxDCG
ntgVibPlaJbNIO3xAigSMgyG6Yuf5Q1qcTfxmFB9OAeKErEUvdfHwB2g4v0TFrvC
AbJT1+gjJFwS4jvBTA3h2S8y/gwMVNccLLh13o9v4Z+QhmKCv6BU6uOsbafJ/Wd8
UGepE8++lPLU8hsncn58H7itgt1uZ0B8cPQhjEttOmn1iajw29zOZX3Ejzfjc6p1
W8DkXkfw5JHTlNxAzWGFD6M5+5kPHvQqONkdONUgnWnjUuD2fqBNcZWR9N9VqIm0
uAeY/mObHCL220yYV7tvcOqY/v+UAJ0VAuE9T+v9vdCwOMr8kD7+HZYxwpxdwSOg
UtJMgW4za7e733dAD94gUAA7u9TyiNWHDbGXTljVdgPWDJiKBx5t9oUyUb74mwou
hkRumeL5XuTQkQGOxpotCYz6g9paKv6fwMZYWmF77dQaJ/35LjftUGOB2TJS08tQ
VM4a4Zr5tNn0b02VLyPiqBIJPWyC/Ai8oKkhY/ln+Tpt2wzUgKcsOWfu0F8fOQwz
mwj5BZk0Ub0fB1PcaiBSnLe5BDlexmUc6ainZ+rKbPWAp2zelPeyvIE7SIvxEuCW
9sLeoH1+9bk3RZy+XwOb3XJeCfpOQAihSkGHfWh+lrLZFNj1D7Hadq0nYML6EH9W
OS7908g3LaoQ88anTzH+y7n5r9jhfILBGSTaee5zUbO1Y9BmaPKmdlZ7SgYji4YI
Ufm4l4294sc0/YHtK9WC5aE/yZA0P+DG2v4Gr+QJSCLzEZ8V0bJKL0UXwFp7cP4/
fUlavQpJDz0i1/TyfPSmglzcQmdtAZ0PPhpJwyoY4LUNvQq+K8GyfbNAAvMgiirH
TgMA/HRtyyar33pJ74npetDlKoWb0ir6IxHoAp7NaZhjfJGUMdqqPL/04YXX84lW
aBXp9Z+Xc5B6b5xfBSr2dR8LXMh01ociJbW1mG7J72MQAkik4E0jp8S6y+4g2hiH
Cb/AzobmiIg7lqmc3S5Ypz1iI+lltd8f2sdQ5396cUkjrkoJ0eZVdrdDCeTcj10R
4MtVXQmdSyTs2P+C7Avxtsg4Q47T8I8l96UJgUNswnxmCl7qo8GeFOS2bkpyx6+a
h6d7Sh6YPTGGJikZNG4LyVq0wWbJp5debPRoZwyfu7ehJCFjxpBxzMKbTB+7y/wX
KdFvxyHCwkzHeEf6dA5zMo6c0Up70djT88urQ3BH4amzQthuThc+e3fwgD1qMON2
RPHht2QI3WJmdA+NQpGodk+tI6m3zYu5JFUkTW0ZoCupZchdB6qKUQezQts/+0/K
z+Jr/qUyLt18kJC7dJKQIEy1WqpTYxu1v5wQB2hTKZu+rI1/m+z6mNhzf+FFgp4E
g93+ibjP2NLx4fE92Q6v1Xf1+cuwpkw95mhHzH9lXcF0ImL0x8xHipPSQjvbjkCJ
tNxr1Sxpdr+O96QXqLgI0HoXgaG+nnj9I7jf7mt2y2FxV5Kk7a6uvb6oeeLduhdi
Uhqq66Qj56qXFOmK7dg5zfQ8T+g1TKklVDrKaEvNSAP3GcVrv+intMfRBLbnVfOW
RVdPgF8OBJDG/4g5BZWLAgvmbmJCyUCB8N/mewQRKzkwC81tMDbBiqQmrGurIdco
+EJX/v3Jayc/BRWaSiNojiYnMH7LzXUpogA5psKSDu7ZaSwCXmAnYElAge7Dsgnl
04AGtxo7jCmWpmt7zlC2Xipj7Hiyd84EzYbU9GbM5sB6EoqputcqVKiyfWfigT9f
OhNgOD93reLb4REv34YIHJLLI8P0UnBtbwoKfjrcsEzAaaQgdNkBwQKLj8RIXn/Y
9A18pXA8Rh589PQZDyRI29FnUlUNnT9WGcpnGfGlZTYnx9kBpVTJAnM1hT21kdkI
uA1Of8udM1Bwd6v/Zo86jXgKzhyDZq4/jOwfvx0QhgdTn+wQF77wEHT4hngqdqiG
+fPSxm0D40BZS8ZHVcPmPv5SQZ+PeftieYyXCVf43emn226Kd7yq8k3/ZjlZ1/sC
0MsZll2CufzF42VvSl8zNjVmeFGNTLEkif5SEGNmMUHmvCcVUfuf50cgxsTDOSCQ
zSUkxcHLnZz5udVGfRy4aF6WI0f4uAZKjWnyZZ/6WTg7VraHdq9udrcSJ74C4Y7s
LhDkVsxi7Tyc1JvqLmi9rB8+qizKU/Mg+tEQOWAHeRDWxCLcBrK9ASwClboa/S7L
/xdjbUuPEb46OEr6riorHW8xXCMlPiKU3CQkQ+r49lI/CXaamTDP9j2ZhE+NFXa+
KqGVoKMarVSUulwsCUdDzL5vR7nxZiC5EjvFYGrUIFKm7lNHIKM++BDiIbPvUV4g
ocqyGgSAynOJbGZhZ/86ujkEfIYz+ruNUGMzJVom7SNah0AqkzsbVe4a8kkZqIyP
uSO30/fRv0+7ufmgzkWsvBWw3c/g/7LMINQLGkRW4gLvHoIaFy6IcCMoTFxn9Byw
p9w4fxXBrS2WEgF7wW9IzX1HSh6czFdrH1Z/EB1aE+D0JpROyYw72ZzYYpGWWapJ
ZkNzDRNer9nEYtUrzVZoePDiKCpTA65Si+szSkCypI2XfMRF7rU+7kj6uFremwQ0
TAW0gYfGNvDztP3sBQTPmtXMEW+fbnFyQrRAwUfM2twjLvKs/c+SYaBrTPje30wj
s1dgqqJGTtE9hTS6PpvEJWDnG41rZyXYX8m49z6DcEOVtcB+QlYNhKjSXome086q
UKbyJ6HMDpA0pbcTXiFDUd3+n4C3zgEVDOP8fjCp4EBB5nkWdMzvYOGg8nkz+5kS
Z67rKKUAMpXarGUN4c6Tm6kIIabMdf0RcMXU0l8rrTz+2Isbe37MtwcFxFyUCezg
tWj8+Vl7qf2w0X9PH9+elxBj5EetCbPq2CEmTtJJB3+BKn6Zd7VYdyR7IbXs/V2u
F1lD7pWiax6otBnqXftgkJaQ5KSUPzDHn1LjBgHkX2R8stxtxPCeHwjfPth4cCk7
mgmv9JUFJovzc6uvufZJ0CIq8NQVgwgDigvN53sXHaDhzVDHb+/+MTVGQZiTFPMo
ycSHLL4v1+eaAxJUJr4aZpWI3fwTAA11s0xpN8yJIh+Hk9gQ/kBC/2Nopa9LSSUk
k1jiefh3t1qjeZzDFIxTj4sFsdj2Cq5dnhTP4+r13l+m2a6uQZZURigF14u0kjIS
aH6B/ON/m4ATLQbr0rph90OXyTNYDPDFes5RjCy8PJ+0LK5SdoPbbIZztjygskwk
iuSOJoZTE+re1kdwMtc3KslrLsXq1U3AVDsWxxzdNugufrXLM9kwpiqSNOZHRijR
EVd1X3r24PXJJaKjePxDY42NBqHEfPV5+I5HuHciOWBHqxHtag74EBu9NxXyXR+q
C7xZ2obbg45uMRJ6YsQZxwXoJI1yl/laPur6HbZjgmyO1osSB3gz9UQQrci3fNhg
MHiBFOqZM48HLFxCRcjWxRZ1+dZsQ/K7LOJm799Re6S/n7YKp5kOal/aoXKJ5qND
XVggKgzDaXiRT8qX7q84XQWnPr4X9eM/ki7nd4JDaxP2UXOYkjadmPBDUhTjAm/t
bM3hs5RII7jDnA5/l5G3un5uX4FQFFQiTynI3H30oiPmjaVcuR2iQ5JRrJL7MvZa
7USzw50wfKzMXruCrckzNZVGgXDOrwAX/kS08boQBp61eeg54OMbo8jxqXr8VJ1J
XYNdqQaWqW6W1xyCOD3k6M+hJ+45hXP0VRWKNJM03+E/dz7o/LdKyjcvKtJNFRP0
f/0YIoZRsVV/T+u0fqpu70Iy7QCloiwSaiaAGs50GI1xyleOA7IWJusLPsVQNbxs
BL3D4osPUg+9kvu97LOXYpt8wciNbSAxXVrTWfmXB0RPKF4rMhZ//FE5UdKLuOoF
h3rcqiTewv+PytlWVshYdVmRzX9QkhMh1KaJ/teMdwyroyiXh43iqEuUChEjPpM6
n2Ho/DhOjZfDwt4CZZ1W7poTGH29YPlcEqo5US/r7RKNgWCxE3isvoTxXG+Asnwf
4Es17lOd/XBwXAVQYBujNjy2TcFCBnMzMED+UlKzdH+VuzjLHnbJ1PDGH5u+ujbi
KsaaxwVnPCvBl9jvr2u1lfRZDmXTE7drLZXaHh8yaLu+BFvyz9t+D150ApGMp7jv
XhKihuWiV/xTDYSfLs6mcFqimIKZ/c0SW1O2dVW5I0NBpRxY6BKjIveR/DRbriDN
H96pYmGsvqAz4UBIn6UWXduqpIaXPwApwIWKs5rDoHpk0wIgTV1W6ahihKT3QXa5
AkctodJsnzoSWcmO7ZXs7gcDFGYXX7FQ7VLQP716tL5l3ulaIItWQhiLnH17SoOw
WAe1QpFp2ihNn+naEt8jowogUVruuNThsjlToLyfSH9MAiDz93XN7cBr9+49nKff
SFSgEQjXZuJ6JBgzjnir8Q==
`protect END_PROTECTED
