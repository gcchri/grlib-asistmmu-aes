`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uSC/rM8mPZ1Mll4pNgiSCvt1ve/nY+gjqnrvj03ZiKGufUpoSVmzUOtoofS2AOpQ
gA1WGl5msXSVxFMEpKW6nNgE5OejrymiwunVsY2JvZQf/E9HAZzprXz7wdK4AwGd
l49ySJip6PNJUB5r+MjY3TR+ld3cWYqh1f56o6LYwyQmNhcKeeT6JVoFvsuHVULo
n8M3dULVzPKTkjNbrHgzXhelJV8K3yD7tDy470fnuMUIUENX+N5qV1MoQkKiO3yp
oj/XBKeuQQh3zO/duiHVaJ1K5yU4rv5Wkr1CMUVC4g4ynqMKihMy5jIMvFri/Wx6
e7aNJHCeXJ+as3lbO9BoN8JlTBLk9M5+XjRZI2CRCSjHwFsYL7+VduGNQWGS65Jk
wv3IhPkUCrIIMn5DFOEVhFL95GhTFFuVsjvq7DEJ5N3cQSowunny0zkBrnkjODfj
`protect END_PROTECTED
