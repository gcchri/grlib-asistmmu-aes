`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zToNDKimpXDD/P3IaoQ1Uo6ezXZO6qMVsbqoTT1Kgo2Jw28WLbv8NKg6MqJXkOtq
2NfkRnM4SUmJGVJezZpmWbDipfxpexKwCtZYSKsVv7egjcmcUnizeqMZWbYdrcGB
yE6zI2j78/K2mkrFBAa4SeasQsj5sHqdFO7Q2BvfE+7pXkuVMl9h9K0ZjE2MkhRC
Cjii/FZYtBZn0jMKT6EHgc+W6EXaGmp821bhcr7xvT9cckiqSK8wSzjHGbYgSef2
5YTFKM5uXWEd00Ugntk1vseFr+dZivlte5+N2V46kwD9k0c+hYYHdi1d79YhjEDB
IKEuxQn0F/aq3WPksu4aqKtl/qWkigU8uU/Zkj1ehTJXT9yE6iSXwkrymb8h0fpK
3dEixe4kvkBwjV2GvmR6owrofpUwquMtcgtj3YG07YE3f5mF6TaTDrxTpPPzcEbD
D3SOoej+YAMHfEaA9VBFO4MyTZ5b0w8x9StANpmlCC119fJBJkYpBKVcO9jqhsSL
yoiEF7RlAQ+/4aXIvLyxHgU+B6A+3sIcgtfvTNcSd5nKwuJmnAwkvWNOzo0+1e87
1k6YCzYHzjl9yO3rPtJ7EEm5z9tLTU3LJPUej+xtFfpIXNXpJRT6bllLPKowwu9H
IeJqKHeV2wVqoraH1+P59wzdAKLEPrz3pEdQS3SyrE0=
`protect END_PROTECTED
