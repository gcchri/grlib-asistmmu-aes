`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/n6gUKJhYvbLydJc0khNGALC4kyRJ0sFe+QHl2E0zAMYJNBBvTOA+F7qNI3y+tD
hMAfGju+FAkX9VFPye5Oqc/Vh/lMMIo6pQ9uIMYM9zTIk3qFhyNxt9Nvt6yh2kq6
lCNicHgwAGCXZSCiuYwDPmN7/hhYYoKeJl9Qe7Mf4VrUyLtELGkANA0XgY8wcNc0
L7nfDy/quZbWIWxzjiGGtJO0FEsj+22p8SrLATbGXyWRpj0YcrP0+D0AW5a8tL0m
CBSosLtVENhy7PKt7hqtpaMjs42Hwuqx8OZm+kEIft33wZ8bplvncyMmnLeTGJw6
6Zr+1Izf85TgMgpCPQtoxEcHljl/r+xl/iZAssX+BEy8GWRsmOWYKZvKpKSbZJa+
cpjeISSQzeO/Fdss1QHobfTNS073n1DYN+xtCx5eMf2weB1va0Hi94YTdMPsDfKv
iQ2b9iIZY/5a50DqN6Jy1Ts/gvR6RDXC/ozlx/KIO8Ppso4M3AMDGNkJmIrVReeA
A3I+ABdghmKNgrMguneKucInyZ/8afLkpA1Jk2CUcvJrh5akajuSM+hOUqhshBbi
b3iWD/fMUit5331eHnHD2qYwescVpHjWNS5KPO5qhDzmwXXddihAbV7m92Y9Xn7S
eA9gtQhPpEebAIrgtyRbSXvWKg83sdUOGeOLXFl295o2wHwCSohmcvj8pk5UKMAE
zj6B9ew/arifb5E5wsXkse31CpJwmdV7INB596sYRiDgpDsU55+S4I5+6/AgMOws
9LnNYZw0gslHQ3KRtGPs6RKT/0qtgC3bjcAKTnx0EfD1EajiYCsVwAHsEWCaCmZz
xy5Et+kD0imPzHowtGfbF2v+6QzAyaxXDlZGTI+f9gEdQchIcbEfGeiKIdcqVRmx
k9RvUIH0O8qTHM2rPfS7W1rOSxOvOedHyDOhb39tPHoYTlUXLE7g6cxie7Y7LL9s
T3zC3tNqYraG5GeH6dF/OxMu7R9iN8MQ4B1aBSMy6UUunBy95q0DDQ4Jwm2kOEun
qzbaiqbp+ofs65ymzceZUymdPwoI/HK+DSe7o2YeKrvmlkL6d2mc+uihziWFpdcg
cv02fq3JzVPXAkXoOg83MAqFYvzR2Yzc1GotzbSCTHTgkBSSfGy660sUpvN7rOH7
MZWbWrOc7fG6E4mQpMIE2cCh4uvcbwLuCMpU1Fr74V0vhAxI0K9lUxrVCR4UIz8H
L7qnOM5efoI7dIwYCP+VKPipo+MRHYA0nI+rTSDM1b7GtV6Ak/RTvmHQEaXs6ZDd
kctE/gEse2hpux57yFPGce7Ai2qDBHE6pPXrrWb3GVdNqQOSO3AbyucWNn1uQccp
9a2+tpNLZrbVRYUBfvKKc3sTVoH/8WjeZK7nCfBHAiEWizp/N2s/nFgUKAmU6KZB
BYVr4E7meP3X8KczMip6ZYdRprTs3Dwb/Y6ytAVbB3SZT4nzf/foPdJzLa8wPHkr
PgSGeDhKuHY1eS3/C5Hs77BkLXhFT/7QI/LAelZw8pEQLwdTYkygQskT36IoM3gb
38JKmfasbgaP2TjyJ9gfC72N5TZGZ1g243cyTMiVg9saE3e+sSbVbY01H6iQwXyt
U7YcD/XuqD1+uZzvr4l/5LGwfvDzm2ddeTX9tgbuMoRduIs02Vo/ewrix3jAJ/Qo
EOROQENTSzCko6JVMAjARdGfijP+8RT8RnVzy+tyymr7R8/a8nyzxA+xidxlWHas
+b4TrPOY4fu3c/lxxCktURfz/E54vDLtBdK+EeCtwm6Xqdpxs1l3E690g2UdRBC9
3lvqn1PtztN3cs0jBU/TntEqDJ/agHlX7lL47gZQl3FiPoJtp0s/UY5aJx38/MC8
7iqwRMgsyzSlQiSr1iVnmbr/PmXGOLL8ZuM+WJw+WgJQSr/mFGeMJyvV8bJ6FaN+
a/dy2oemWYJ6OoyFZ5rLiYhyJ/givkeTmPmYEHS4qXhutADRU270A/f/JC8B3AfT
ppjtUKqjPXt3IABWM+Kz1B9f1rgbUt4n6BLMSJ1JM9xPU3QHWWBFZ6QsLk19atZv
FBaqAaWUxB8+awOMrNtj0KSwkg078PY/L85UBYudIZ1hthRHi1rqtwkbQ2ZD+i2q
15QcD5QLevqNeA+60EhpXTUVYmJ5zDFYhuhRSNg+De1ScESinbLp0LuzKZx9pfeN
uR0IVntyol+s3HwBc65IMDkQyE1I0E8fg7aMKAwBhW3ItYtUwSrIcYURu49D6BCT
GMY67zy8XOBghxR90PFAwx5oE0p+z1JoEIORe1f+qPrCfLFltjguRVl/zmLcqzlz
iaVnAxgh1RZFCvOqI4EdDL2nMV+W1/EYxxEiHAjMboOO1GBeqWN4buVKsWv8YS7y
DvunxNTy1Ufa6KhghurFKZro9L2e7rYvTsb5QcvUfXCWS8tRhuzR+CqZikWnLEVf
4ZgaH/1RuzOzFXw1wMY6Yjdvq+rb4cNBVwik7TowZdIWqFHNp6fEUhiVVFXVDAj/
GLx8jRrrXA88abr3IND/yrEhk2i8hXVi9cH/MpTNaABlbryO2yOoUeYvhKtRyO0n
dDi+VKBU5MZqcIQ2SItZ2Fn0XTBn/oVuYBmlLHQdG1ksZCWNXbIiT8ilWpBgV6B/
z1foW3EilFEaPVmsh05R12LnUjUxZ212pjjqtkgRJ+WXZene4WBQk1BTQpApnxyh
rikKy03ByfCPyRuLHh9GYR2B9/wGbmtECg+QZ7uk9lva+t+W5nctp0hkzpyRiujO
l02Xq6M4Rh6f8uRaPklzCBq6yVtGt0NleusI6nxZ0+M002kCerUaQQiTM+ZNRPqT
KHOIGRk+FnW5caCWjwbhqjGQG/TLOtkKLcbeAtNgXr8TpLlTjcwoTfpS4OPavqyQ
H7Crht6aRPpFqRiXWNKUcrJWgR/MoJMICHtsftcPzigrSl6bpfM4FqByaiDm20sr
T+f6SCO/VEzH4OKxwMS2nyuL48H4a15ELmwVrb2glhEJ7cwlNc7h2InLTaHWA4HJ
Z0EQzjGeX7Q5UfTSyxIe21TRkw3+jj0ek2e5NnKiMEoqudgANFa4Tm9ffkJ33cfR
pmNvampaB4M0atSTCzuETbTXlYb24OlXe1zrW1onnoPe5SDiM+bGwByZBYw7n4TW
plbvsKCdmCD4d7lbul/wD9LfIwSS2zuRWEHrerXhxmpgRx3zdIVRInnxSCD+nbgZ
aLxFckrCaIUn0STop1FudCmI0b9SDBQoLDxVAGPgwE6GMtefoxfbNXRa/6FE5spz
CijAo0AG4EK8IQWW1IkdEgJl+4M+98F/jJJWqv27xIkzCZLraKMeYZUUEeQRC/dS
2HErdkZM7vvX5hKPdg32CROdjjNwJRsQhmB3dA6TtO6+Qh5/0Snt5bwI4CQ+MEUq
eOceoksP964aiRLBc1E4q5RnEML0+we8g44siPH0KAmvBaNEqrXfBKLLCmVbW/An
p8wxfDBcDX1jNXJ+T74kbgcWGeS4dQgQxOP/c2rJM1w4uxTypuVeaexQG4b+dZSG
34pLORFIZ7iQjxsXSFpnhkjX3U+j9vzCHR5IbJZwNSfzO0//Sgj+QXkpFnfEkP+H
kZHw9ncn64ToDQCvGVmat4QfSeFlcu8ZGhOE/75akFxpSo8wCreofSuqO74uo0ao
YvdkQHGQIfKPJE+fc6Zt6EsT71S9nsn8w12yCxR26eeYexm7Btb4SQjRHpcWAu2J
3FWCf8vPlfKy1c95m2xHV+j4f9jpS3WVQ7vCu5LZnciDm0yoJEi5UrywyjpFTiYY
sdlFIpgrJ9DcELkqcMe6zAWlOSRqlIZlFkfleQEoDQrvhhMw1I8TxQGX9NW7d0yl
0UDKC4NPD6NJPbQFQSnVWHVWHi90LKP4vS9FTl0enlrhSERweOX9biQ1goBMYkVP
jXS6TBhhA4CF81ENmtDYMXGGa7LFbSpSLbVcwWIBbv2mKpMkrzklOxfZTT/LQhql
7/LpT5GLJgokj6gChqyDyfGJHe1cg5/n8vGATdaPWu/qgyQ1FRKcDx1DCpuTZ0vY
eyHNZBR3ADPNk9fHAp+vkfujTwdeFau2QN68/LLUo+Rn/hj3KVuPRptX8SIjkFgh
ur/62DKIj0wY0zTwgWXiPECDbpPyJqZOSrY+Egq0axT1rRFUnv0ZPSr/916haQSk
3c8HJSh8MK8+yPhxqZechbHq1qno+OUMZl7YnMLVLMmilbn9IwWsdNSH8dmjpgTE
kvmM9COj4mn0Q++o4e0meUu516yD7+rFQ4PVTJmSZ4LzQa+I1G94zRbDi/BWITts
/vMZiJuZ11sluQrngpq5VvGJO6KiYG+gwYAr0gfHNDzGFIyf3LT9oFaPS0OG620f
4d688hVOsczROPga+iJCmq1m04Z9cy02GQMFhYVpGR/me8Rq+SnFVWpQvHZ/r+sN
jP0IHFXn/1lNf82A5+73AACKSCrALEhzGp9Gd14DGADyt8nHvVBKRC0wmO0Wyusw
qPEIZS+V9rVcHP1g4sKhL646gayVKVOhqNKaPm5ClissH34uv/ge8E226WTH4q1t
LXsEf7rWds0GfHaldrBQ6yeYup55edUlRRRmXwBo7Ux6EaQKN/PDfrkvQWhPeMu/
QmdgkYmZTb7HT7cWw4rbkBo2EoHjVoM1Bj8zbipgggd5dyu9w7Xl+k/XlbqFB9x7
dfL1sUUnrP9cIqobY/lFUrz/A8wwi5BUjenXcBNmvzUJQ8w/FKrz4cpu+g/ftLGc
DiaARhbDH+E8MA6LgjslQiED8GG02y+mBtco5L1XrEAoGpthYxbAFiodFd3Hk8s/
MSjji3kYnEXcb+H5+zSDwywpVI8mREhnmRhGLSQuHwZ/zvULJXHGQa7pwNypB4YC
h0HpU+zrWeH5xTPfgurcWKNypfne6Ri17fMBw9C554FeM4kK83omcTh8DzWRRXrj
yjF4Qpa0VbrswH8GpQOCEmqomjw4njojvzNGa33GgLLmWainlLB8uuna9qMCwQG6
des4Q+yQbR5w2VV/FU9I89wVp2vgllNB2E3KYE91RcBnChC58BcHTKekAEWa14kb
3bT2vDDkMOCuCJMfJXdV0G2b2YToSCSPBzCmpCA6F0kmi4aCeNk3nUfuoyNnPyXK
`protect END_PROTECTED
