`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dpa2ES0Bsuy5wXTqUtK14AmhZJGU97UlG5H3IfRJWFpzm85PcojPg+eza8tUf2g/
yw7BMG+HFgc6SNZlkH9Gc817lQy9XU2b/epjyztMu4rGTKtyrn0Ts844M7APHO8c
xul7llrgbVpbBzaXDblk9IzKzZz3sNbQppsd3yMD2uEevGbM3po5c8fb9VKVs1kM
wVMKFVA0eL7NEvT+5/eTVEnxy1GuFP/6bqMlOiYnE19mCJ9BON0AUdgD4lz5wE+U
StooLdfmjBn67fBpLozpeTz/CsDv3XRhgX4JgsvB6DlZUa20kWUvS4BJQAzW7/wm
rUFFchb5ta7lnWgtbojGmzvT6XNGkw/VTeN2QvmKCI0dodI7j75Fw4IHK9JtKRvu
OS2gaS8q4kxftQEHr48SS5KF2+jl0uFEevWBbIVPUNPejXcUyHXg3c8rEiIsZnUL
8qGunk/CsExs0ADqL1AGrbPiuJsyNaEkkXmdO9pl7Gs+mM3HzTf1RmppIi7ET0CC
QKt3XhcMKWR9yVzz2RQw0HfVpXyO+h9Bq9CST42pmvU=
`protect END_PROTECTED
