`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ydcJAIUjPwrg7ICs1LOvsRpuK2hGZenb3RMbCfe2zXAwinUMBzpm0axFY5i6XzkZ
bvqiJbHclCoZZKKPfbR9QnWah3r6UKWzNDKnVfXr+lAe6yYX4+9H5EKMdOIlakPT
H9rwTlXhQSMWJZLZgaPJnoOie0VXbmi33ojOZMVsU+nLMmGm4yAff70pwqCa4k7O
4Z8DyoEC3LdAobXd3nrx8tr2+wfimPof0D1XoPI81Q6/vNtyY9FM109MkcqTDSd5
B/iN9Q7fw7fHpaNpZZfzouBQgJD7WHxQiH9GVeL33WcobGcJNByJgiPYTEMsLzN3
ERKDHN693ciyFp2sKMeiSSrBPohzRn8dq0WbezwyLfHGoYLJ7hxoF1zwQUSZEgQx
LVB5o3IFM+jKrfh9S/Vy5M/IUYqtwgwcaFjzOGp+UHM9s57dEh2ZX5QOr75k3tNO
JCBO/JuLoH+edVpWsnsp1mu9V3zgju3/tAMYzP0QVMhfjuRcLRnrmPyxmLXRC5QS
rNqbmdJclFH45NtcvpZPdXxzRST0iiQPij9lCIBJH4KvSXd0VnZZ3oea27Qvj4NC
idUNTGzIIO54EokXJhVj30RGXRK31Du/LfQqFOlFmPhMXhIcx7kL0mn0re16DBNc
GxBMqXJZbOMe0UV/tjsYbOc7JXEySV+rrNWupfcoA6Uljgx3rYAIArJ0CBC1JCNT
h0kOSISTNflx57iQSLCNvUjly9Nq3CvXZzVgORpSUDSBM7eYJUtIfBxMLKNdFp3b
TmxrUiar0bu+F6ucxLCKFMGUQyQk+Vs9C4Y3rWWi/+yanCcEXbewfnfBsphbJymD
3mcypFOJZ8qRkTWh3CIk9ApRevZ77VMQZArbVd/9ryMlbCxHwDYPikEUlXn7hIzA
zHMkAHxolPIeyURZw+9jGZ6Ic479sgO/tc7af55v5q9LQs6atuTKSY4YHCphf1h3
G1448rgeEIKIouQMUmb0biOWGwMCgCAwDhg0MuGZr7GDMLvC5o/5KVnsncjI5VR8
fY6kUDc4pp/dmCBw8+XXcllenKY90JoyV4r73y1OtBoQR2E7nRjT5laouWPPYp1I
O8LxfymDrMNe2RHwocn4smBUX/MVsRLqWIeDNZTn7mcPoQ+zyFEYcMjEm+g7UsXc
cvcA1oVGC4h8O5TtgL5LtLzn05mjRT3YnUjxKGlt8qBsapH9cMGs3YX3G4hjJMyd
MaMipwsGaIXWabfDD3sifEngXzGGaAKjaLb5NFmp6u5fCmbyoSt5hvEf8qAXLxlf
x08psHhTPViy94JNkf4LntS1hxnlIXA6e6a1Lvaj1WMsoxwDpxgnbD5J8usG8B/L
n27KqAvK9QjgOhQV67aW6kWwte1x4eegA3eu1SKAp23uzDwkaK3dPt1dmwiKSxvv
/0GTnxvaG8dm+ZoEevCd+6Ss9h0ZPUDnRzSESWNVKErAqJ1y21LePF7coK4D5U8h
Q7FY2ZgOUcCi+dh1Gr/JkfFsHqBoJgWCPojzY4VpUYJQ8nqj+Cx5qaRgX9V/v2eX
erD+EQiehNIrrD9eO02aTCodKDRcf6LEl+f6hndmX833RJif5HAmF+zWYxhzRVca
jd1+JFF9+6vd47UBb6+IKYZxQAGks0zBhEc+yx0Bb2PDX+Kwv0z8S04sl6hse/Me
8cMV72Fgc5a1Mbld4G6Hm1SWD9xUi2AV++yQF5Hd4Bir4x3BbxgU7s9evvuusIox
zxiM6sM68lzcbLntOLLbCihZJnKgjzx+E6E7bnJhWclMdXZzWTXS2mC8y7AjcLSZ
Eeb+B4BR+pO0xUL7TAGt8Kul44LzUZJTpSM5Bpu1oslZqKmZ1NcWZBLQQbf8ATsp
uHWm/NnjVowwxuQKFE4cXngXRQ3u75hIcbuxXWFH9gl0n5AY2BidTe2yQCncJG6R
Qa/ljCfqOnoTukTMtAHeJzSV0oHH1rmTxzCCOoxtRMRRaNPAtSRB59SGEagobVB0
qknGE9Tmwp5TgA4htHIBh05QV0jKiK9wl/nq4Tx7Q+Ef4M3ugB64mvYpiO1oqqsW
TbPqNjqx0qI0FYF+czlzT3IgErn7HZCpdu/mF0lW4u5LTbZDIW/mmCtPfGsVmgQ3
LF3OJAyn29kpW8HGt1SF/yo7w9qLLSZyWtNTPhEa9tTplan+2bTLUF/GLcoh5BvL
ev5ChpRm+q2wNGzfDnAWsItkuf+E1eUcMtuCjl3EMFLV9jat4kHmZJieYcyumk8i
F4WA7xf7Xh/7P1QiyHseI8NL5FVNmxiCvs/96mHwd/fq9cVFhzI+lDI68vsaYYpo
VcFmD6N4aeh/aC5EkHslVB9fiQuzx4rOBtMU0zPqSRkg8BgYcwiWE/5/tcdYNGA+
zq5ATsiQTb/PuJfxv/abggcEHptNU2ApdUlG4aFw/Ba7HNsHujslZPaM1lrKn9P2
XmHXbMTDgEWeOEHCelBOchV5JWgMzkYvRFWIxsseHlm61rF3/1cMTlBVZNYkbpXQ
pVCw9pbpP1Ceu/8ClJ+/pAzM0b5x+qNCfv1gtbug7oErXbR6+txwtO6Fc9e51UYr
izgKwHPnMaWwN6Ec8sCRuUKHNQCGnyvXfiQcWS14SiwY4NGcfxxGj2Ypa98NRQIB
6n5hxc/Tmk360DSXbvqrP9rFFsIzdtIwPAnzQmezf8W6AKYqyuJGgGmX9vQovRAP
J7ql6PNr0so1zeo3NCLYa83L3qb4P+b/UaaoaNAoEZHNtr5IyfYqWnsrTWVIwV1y
XhFj6ArtTc2Pjx2ElsdeJK/+Co4DHzxTLjK8WAech6TbxtBdnwLHPpwfiGByuCoA
FU8uSkH56/ATZfPz4u61UyxGglt+z52MJ/qugRmtBWM=
`protect END_PROTECTED
