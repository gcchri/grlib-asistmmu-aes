`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/6qLLQDwdFdBEDwwSA8yslhOWkbiVketvvyDN9gB4wYovbMLpLHPmDgjj2qa5jD
6zvP7GeLa8RAVNcJTzkAbU76QXekIEnGamB4CcT617ZI9Ud5ygfUGI1NwxHDAaB/
Wo5aAdErjTan09nOgS4Efr6DBsX65ppTW1R044Bqq4iWmIe7t4XVb19m7seRQ7bf
ijtTDFT1tR1TQhnmhSEgpLrUgCh3vRPMKcuuxm5VWlhw2Yf6sPx3lROWL+k+VhJB
qK8NINAOTr+J2cDvVRbuhe3RheRXYigx0Cjw+a2vn6/XxjurTpjnlabOa8mAA1aA
vvmi5zYzg25mUrOknAfLt2TAabROfNwQ5Ou8A3fYBaFNGflAFjwcutyo1EdZQr0N
8DW/UPMzdQ5zTTsG0mlFO8jt6BFy1O0i4t0WGGzxp7Um5hZSG5pwdjpHuZiD+1yA
si2/6/TnM0jMgHZEjnahtNNSSa3Pm00GCtVJRNgkvjTmpO6RMooCnSLvOq67aty5
hG+/oq4qJcAjvBVUISwHhvSYsl19Jv5ULYq1c7+fA3Ea29dj3g9rbrMGecKE1SjY
Lb9HEjCYVAKoA4xUxVYqmODV3rMnXqoxCa/+W+NDqX4=
`protect END_PROTECTED
