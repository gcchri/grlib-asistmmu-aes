`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mOVv9FnKWEUOQMTq2b6zIcmuLslOpnc4BDPy4s+NMdDUfSYeesIC1l/SbVmS4YM
CvogJPNo1zGvRis1p3hlaJ0F75LVP/Qt4XnLoNR5tvAbmkbnhwO6OTcToWtw+AbQ
Q4OJW1lu03ig47LOnDzN+NP/jOq/kfQpljTy9gwfwMtF/nasN7IUahDL7e9k3GTs
BNnTRsTT3dWEKxrmxSrs8WiatkrgSPct+28T91E4yR6zfVRG7d7bjuiXIvb1IN35
cs4VTzujDp5wqDHQ9FIbGCe5FwmPDsRyMJGjiLxQvHsoTNNTSpMx/IE3gM6OnpSY
5Cp+EMz6MU4/R3qqpJYDwNcmLmKx+/nU8Rv5gnRZ64byDr21B+kkAUIG1e0WBq0/
qqjFtHufGfd0WOUJqO1Sn4RaF3GGEefwxhArcyHG47nqrSBmo3vUMZdtT+gZz3oo
8u+n+u9V+f8aUwwWrp0tKant0t4HUOHQe54Kr6VmlNBKPHYDM6iYlvIo4h7dueeZ
t4Pw3O99NPeJEZMvW/wbGBQxYCwasRxH/NPG6s7xptwz4oKbWBFocBF0sEocHOMF
Z5uJQNYRxHKz78lA7TLF6lzE4k8szPn8HuzBWfYP0JMF/CIYv+zXCNFDdsPyjevZ
b/HZ2Hj7dJQ5u6/rMpYxWXNlO6fiZx0/1XiMT/D71itxdrg8cjgBCsbp+Dz3HvU8
E4JCOFtSlYwZZhvyfveZJH8vWhxcTTQ4N6pb4pKGsYcUAkxCmAhOEMUST5m7f2hK
8cEdK4XzUSsVtix620U5jWNMg3UI8qY56Da9GXqryhSkkdPXv9deIhz9ZbI7LOxH
lW/c8XbwBq3I198qlecpK828sgRaEj15/lHk85W96XFL+C7EZuBUfkqW3CoS/KYi
fRZkHHmTNDym0+lpiUYmNB1chPdS5SA3NhCG7Jiqj49H2IBBQ78NLztBEX14LeDu
CFYD2ITzJ4/JxkrVr4bxeK/D8sNcsOBCaXzeERNXEmuwU/nn+taHeN5MHuVL8yjY
5Hv0uS4nYDsb77VhH4vpk2vfZvNUMPtBdU0mzqOVknry/5niZtAbH2RgsvS5CFEe
IVUvu7xt+yi0a8bZ7geLYiVl1GjXrl/G4NV2Wtd58mCDJk+4DPUKweQrWN/QcMAy
QFQ/NP66TPwJw68cCMhgiOie1ruwoY4cnvzlAD77aMLYUgsjt68oRqLz3QAn7cFt
vH2+6Zeuc3dyK7AfE57hObmMul/mcm+vDyumaPq4ZEULiTuechXLPPvzsIyH2XWW
FlLYPljR/xxVGjou6SJGl6EaCwnUl5jQRf2L4D/0SrrzrehIZVQ65+h+bTdK7IrN
qdNE4AdzHilYh0VMxzNDICGMGCdrJgx8rwSeMsedY4dEVAHuBuVV+LQCLEir+IG/
KgxIHeV85507DVN9sbgGSk1FkO9HXPEnCAfrji03GX2+aOV6++EqumHAuuRJ0t7v
CKw+L0WCXxlJjg6+FkSP955PGa59e1yEH42OskZtv3TBY3wsI7Pbg5ZtY0rWzhm/
Y+aw4BlsW14roaq5Vlsj1vTZzvNUac8xTD8ihLA1txQsPNMJpWLxlA8XuwDgf7Ju
iajOFTIgFIJer09C86JvkSXcB5OP3WkxNgq2m393ShXD6YKedaw1YsOxBR6i1hXI
iZGVxh2JDfCbnEUheVKOgyvL+toDwvfA0BBHRWgOBqtUfsHECY9JMvxcLLypKXFc
A2VUwQ0KcPePrOIg3aw9zs77lkVUSc2gKbdICq6NFqT2S4CRiiNb9r2lRf7lFnwt
omvjwgHVf7OdDvnaEHUqptPm+T+ma0XvbmlOoCbkLkVKGTzT1l9/XQCInftKqwS/
dyWONV+vM2uD9UYRj8Dt7mImldQJ5FAtRB+XnRjBEul95HJwItrsob3jzXP1e3c1
qfwOPikfKcZUFsMeAf9jnfY80ur9n9aX37wpk79kMv/Iz5QmoS0Ub/zPDsEDKObb
5rscTgwE565ugzAZx5FtGrSc4jvD3phQ9Zk24IbZn2WmkoT7CfOPwk6uZgVCtmUy
OSGEE324rdGdZgCl2TsBPCWPC+Ox6UhrkQnKMWSPl311ka61ZpUfRvpb+dvqciO4
lK7JnPGICHIDr8tSbYP3+5bagUimEenJq/NIG44m7/sMMhyOaxb4RdQBhvQUPXZ2
efM6JfzkxLu4SeY75jG5C1LQWm2cTPkp7jWAEJ/f/WeUXn+ONmjzEtfX5Mj5WAgG
9uAezFlVUyqYJG9zGxZZ/uR+iPCUUKaCFJC79OkCwgDGMNZLEl39EqNeTSyCIbWd
JeGWZRd0M6sJLt6F7ZmINlDU/GuQPdNMAz/ZIthIJ/Mpocxciq0FZ+akxYtC6faq
HQ7aMGbAzEfxzGoL/R9xwa/OjAi+lCupSZ36JRrHehWd3c+jIo7oE9rQ3uE11VJ3
EJPJpiyuSdIIHr+dx2CGcyVni8QtuDhtULslEIYZKVa7YQb2vkoanRjo23VomI35
fBOmpRSlaiv4ZvR/gu1MwIQ8CCc5neYbQiSErmHXbmlRzc3uaDVfIqfjGOMDkuKn
KxugNABVX+YBWSjSJhEvteyHMeMwJeygUXC7Ga0Tp5ZjHcUepbuOSnAHC+uPb/TL
j2WEizVt2LAkK3XeIjgBvVrUq7+CpjS9Gy7wJ4bYCWp1YF5cPQx4+jF6hrrT1Oe5
a2a7Zg04xb9d0W65xEpzpWn2Bdqm2EOu4qYz8/bEoCtS+vA4dsUtzGTZ9CeuWfYc
MRjDoHYc1p9eZEFMOSi+Iymfnw5aa7QdRCDL9hHHohyV77fZ7sIV2ohcon1F7LDd
M8xCYTbkV9noCIAH1a66whARPU+o+EB4/Nu/Xi9nZ6Xa86v0SFfKg2GXSUl6Swiq
DcrRLwn16/p3Irx/+1AOUqUiZX0Bn121w8yhv9+3aheyfvUcfArP2JZ5q5tTaIXc
hKj1mLBQJKzIcqRCOw3Uld/wtX7TTKnQqlyu9AYApA65i548lEu+d68GsOFumz4m
UdgwWTbpKs9Lv5TTCkbj4qAavzSv7qbJru6Tj0Akn16UrCqo4XdRWxexH0nxYpzw
+7MvvrbYqtCxWPvrV9VTUG8CHt1n8y+jgG0pT1gQoNAQVthD36Ou1I1uf6/zSBvq
EKq5E9pmmG2/v+di0+5XNsZcg90hZ/HdcJrXKiyUPNNOZ4Inr15SasyfkhPvrFHY
U94+bkNJLIR4zVg8Bly703P8/iqfGyzAfZxezHNtLUkBu6nf8f9v/4Fx3mZNCSA8
9cZe7zH5XlaMHp/uL7GUqeghgyE3HNk54OAWI06IQd3Wbvo82xqSd/Bq6r094vmS
TZBPmtrkMIYNL3ykidr1nWL9B5l2My5+TSYARdcJ3/mPHNxW47s8BglUrFxml6Kh
WRUeadrJhbthZs5knj2GR2u/bLzsIoGw6X3ymoojJMTtg6RSEhBX5KD4y7//3ayh
m+I0HGqWOWkGp/WVQXbZkbeT21dkDBubYV0PA6PephL/awOcCE2uVQwQHb/94Bir
UHkdnyXC84VinoG9ZVJka6mPQcBiaZmiLPN5IOG4QANkCBAyZuLELb7LqiH5ve2D
JyzhkhZSZHpqb4x9wZMj493K6JdxV9ccmWlxqnhTxTdT6dv/0IXDqi/Bfr6VjMO0
k/khVGBs2Yenjqd33Zve3mbLKLkp8kfudygrbceYqN07fvWphprxi+WTSE7lxV1e
UlCIK3Tn9NMEqiUXk7/vmCWVSChDGVMvf9ljQOury/w9rgh9tRSZkg7MWF6OKEtg
lrnAHFFt2BXQahopFyFH23aMbMx70kiG6p3dsFTQuvK+SMvcSVnD0BF+N8X9VtZm
4GiGxVg65auRnNX/oOMXBWe1n2/LKsadApMdIVsgcjgo3d/mFxvQFqbpBbMyTDFH
ilzB/DS3BXNfONDfIyDZbsUnsQUnOZCSQwZUEaVqMCGfM82R6Z9jrDCrdT2CAQXG
5usPI9LrHR96w3/kKIleBE+DrorSatJsFeHDmUOHWRQ4fT967O16DBVTXyABZrl3
rkbTOcI8bnPcK93tAE9rtIyDv4HPN1o8Cq87txERGTRoOYt8r7tDRTm8wUrIS+v2
y/yVTwPG0rvV59PG3nuxIcLmPw9vwje7CbNLz7jPSJvpiEJBY3IqBffQsgUS7urm
huGc8nEYF6/iYyWXC4RFufg08JYgiZKz1st+7WTLGpkmqxOJog2YUf1yVP2mOKv3
Eoagl11rq5G7lsQjpQLKwYFd1s9QDLPOKhD5Z+yU+L3G+RFLWzuWr70quc/93vLx
qDf+RC5guMC+EG3KBzLmEhM/IMgd4PBLPWVwaIBaNqs9paLfr08z8FIAbE+zOrVD
VCujr7MtZfP4Et7huybvblmfKYKi8f2AxqHh1odvSjdPGLQ36JRGvgmcaOKHxVv0
k1n1rhMuhanhMfb0ELEb+GQLRcGY1PnmASPxHxVVJbcmwfefTM9d5Qhso36o08kC
j3ILDnsBqT1wiGYu4ZqF2Zj86lZMF5ICYmLsDI/mrG/oRbNSYhDC9fhf6jL0fn3Q
1O0eFRMIdLBCGkvf0COcWjm8rnaEuxWn5weSvLrAb89P1lDkTDHZF0tyHpPt1oAl
57S6ApybZKX5EtqBl11Mk7oZWJZ95NfonnuBDVMGFm6SvUZuBKvHJUJS4k8a5V8e
s/YDjx5SwqOHW7ZWY/LDVK/X/8PGZ2VPs/jWOa5UIXCSiK/IhFa+iUQ9Gl6EcrPL
XIkjBSbp5zaZac0yBUhZ4zwh7+f8bRtfCdpqmlh4cPv81q1K/yM6YWftU83WWtxf
YTJIdoGgdzm/APR279603HQriIIhC8ju8hSVqcdiNtn/SzZiS9Sn7/JwmCmV1lIz
wagZgsNTqZaeis2JGNbeeobyOiQjt2grhT83ZtnE3tSqDLQKwXENlrb5gI1+5+Xv
YnajJweQssY5rrxMWMR4+6TYZE1UcO5AjqFgZ9L5Zc+vGvjb01btjPdaFsU5kk0D
6fGXHXrzRAk5VJe/lnmA3PuTq3XyP3o+Ul5nOJC5pLYROIp4ocQVQQG3UvZYSIXf
MIx4huqutbOVUoukIo57fxisy67m/azs8rzlApMxR7/G3/0TOyR1OTGZtEU+YOhy
C3eWQdTmKoe/ziRWbstHTxkqRSbnjXVoCLWIcoH0jJ1fR03aw2dcKncsP0P0Zn7/
6OJXc+ppGuQhz+5DbJLOxF/Xz3Z5VUiq0yiHU6w5csp+W++MTmKEsB5WBAamtxd7
tDAcdzOdcfsSPafg6+zxZSni12nhc8fdqh+MhJUIeDPRs3V5mjDEV2ui1zOviC/B
eb8lZGMyAvVrCf3+xq5uIiBCvQYqZjDgAF1wgZjzkbRHUEbSGY1QpKcGYLQOzeyR
qZ9TOJW7oN2KrVaw2YaogpX5CBAaJpBi38UD6waLCfOe5NY75FV59sIIi48XHt5b
Oxhd/TWHHC/pzKUqaLVzDLYg2zK0a2ikRh6INHczAT26nVSHAr2xdny/OiznDB/N
s2ShjKSTH0raMo+L0kdNons50TrqE4TR0p4MykzBL1SAs3CUXG9EyVWL7Vy3dYkF
2ch6Y9onWV7V6PLHAXDG9xqPBtoPQY7tcmtSQLhn21y01IZyAbbn1PlVZ9tJOWCa
t8pQ+tVPzMCYHLRmhZSv4PFvOQN4lglG2DRmxQ7/zrXF6gK6pUlR177yAPAqMHHt
mfhxE0zZijawKAsb6WGbfeA6oApTTALdLFb/x7Nn1RbS91jnnxFpmircwQhkHQfp
HyA/NUtj+v69viVE7Y21NBGrCaC2tc4zpy2qs5deF/0MiItr0uX12epQqiv8X+6P
vjVBgzp+Jgh6qVKMIdrkWu2SMYjL8etSjF1hdPlXN5Yd4NuP2i38aZ5g4v6kk8OW
sa1NlIQB/cXxJaWzpe4/mGOaXRysmtMgY2vIuAu5QGH6RYDDHuQtU1hXWdLHFh2N
xzX577SOiVe8KeAUZ0HnNVfzJPUO112cuuFawNf+G2JIN9YE+IXLErMJ2FwD4vmM
uMORhkAPDHLlPtbMEngvCQ==
`protect END_PROTECTED
