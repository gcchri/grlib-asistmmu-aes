`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQ3REYsk7O/4yLDLOrpCkgKMHf/kPwIIcCHis7yjzjT/Fbn268MuT1qz97lcd0jW
Nzkjhvwin7zVFTEfcpJi0SiiSPzEkls2DA8u3vdn4M6AvqrZQDqzao7V/ExDtnXq
DySBdAqwhzhmSeat4rW/D/C4pDqCesKuPl0peB2wviR5QaCcWgyEb5p7DDj+GY7G
VuRtJ4oLaE0LgbRHxS6oz/pY0i1JaG9kyPBtRsRs5BZQJG6vEYEUA5nsMMsaZqLG
dBo+kXfSvHK5WuK/l4cHk2XCZc/BzbSWnyul8j5xGUuoxOlzToLTN37SErcYmcao
nMAxmxJGpevpnvQcqI8TLdQkxYWrkKOs6nOjv/aj6cvJRaybmQKUZ82Ncg+1RLRy
L2GtJT4Y0zujJRbJEhel8+b/61Fsp+wvG+d7B/Ba6NjiT9bIaJEJaO6uckMR6miR
GeEp6Id6orCix5ukYQ9BJi8J2TJAV5zUAhr5ymgqibcPreEjRZguUHUrA4s4AVDL
`protect END_PROTECTED
