`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w8/d+zojb/tavNvYCVAXe2yg6IZU9bgG1Gd5+pCUpLXOue9BMw321ufPQJObxjzl
W+iJOi11jpppPZ6BFc4FXCeFu/71Ez86oMBl6lRBOrIzjcY2pDV2Qg0eiD2jLvbz
9B05axrajygtCbnmPOrIxT9eLwqMJXnp6fEWxxaitWy2Qeiz2xN9O2+PrB1Lq1pP
221a6iqvGxcSJx2mkbT+EleuJ31hPRfmD2HExUnOOztQufBRaDTdy5kFvqjSt3/Z
OvPxTC7mp6Pz1feQvbjaT1IQ6ik58LHFpog4opanvPrdvCo3RY4mtSU3dOpKhL7j
oSlDNt5LeywOnEbcEzlMg39OWYX+DYjMNk9Eq7rYiyd72CgETFBBoy+ZACcBpXSr
4+UJvHDPMnwLJC3+s2mE8+BMg8bWS+BSqxLh9ra+vogZT0h4ZdwN8a14nEXRMdOR
10f4V3hYL8Gpusx4KrGMONmF/HKYjgO6DxlolMs+DZuJJtZfOZDlTYlBorWHdPTc
0uL0+78cLoFiqD0o20VYvYBtIAg35CnCFS04+FkMYRr3lITN5RtWtJhS4B7MLWf2
o37ifMGfTXFuuGYFub4RGobJ3Xs8K7y0adXuA0faWcambvpWqA6kAyEoa0p61KbS
nRSYQX0v9nNbKyxO4TkEJX7Cw9THFMGkBfPzJc8Fb1aHvt3Mm7hZx7QV6cfR/bqT
2LhXy3UmiGBsjr6Di/LaiEx5wKpJU612yaXc+KbFmZmUGHuDGoe/ceCSszEG4uS6
5xNQIfY6RPSDMYViPVzktA==
`protect END_PROTECTED
