`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tuBZMJYQiSk4aL5w1amXfDnc/yvM2PygPKeRvA1zRvVPs268/GPZjtCKspJOwZep
XAiRGNeOx/FHA/uxt9uLyMKtCPEv1YvjNaf2g45iIG6xZhrANlqW9i7U/ORiqmXU
+ly1+e9r2KyAyba434dXrg4dhV9uNGlS6v+PTtp6/UGuIcoT5+UEddlFYN4N52z5
h/RDPCF5QHTV+p0jEnzixyXikfrw90JOmPZE/pZKxhRPuMJ0fSdx75dFww+DKhda
yZt1bd81QfeiT+MAVpk4l09CNfHniIdTq/kofyI4fFm0c2IeeanV6tvQlSGjgYjA
KoJfDCfzM08HR1hfLoQNvw8FN8aUJubNQvabWBmzL41qharpdNAwC/Gsw5trytfx
NrxdnI0cBJQepPj4asNg0KPwIZM86NEJTHzOsULYSoGotowqjer00Ib+2GE+CTOV
UjClvczr8UhG6lJcUmBNieMm9aB/9RBT7Gv7F4OmcN2ULmRNcIr66Dqmt853uPWS
`protect END_PROTECTED
