`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFUnDlNodcX2x8xvraR9Tws60pRVTtexMMGQbZWmS1Lzw9bP6sOfHPL/6/tLqKUo
HlhfpkMQDakKOJ9CpldZwPyBeFKGJnxcvxUp6Ega7T2VVVMYorXgxkRpo9dAToSF
GtaasaG8jxYDjavtuUXBco9xTzuQgoA/WcKXb9rfV11euZzoSo0Cw5xX1i59JfVU
+jLpVmPayi1mkWmChZLQX6lJRV4rJAO30/AbWlFrmrboGj/Owq6qTGC/tQco6MBZ
32JbEVFNpPGRZwUL0bOc+/OvYzoP/4WvRmPn0x/N2MI5rfowjHccfc+JFbdUQGiZ
K6zrO1RawEBsoe/6ayavMxC5qTA0bxEbvHNUVIgPW3B0jkS6bMwWC9e/zU4BRqG/
yDSYzDnEeApKyE2CtyD/40sUdVEFkKkcywmyO6+GcP6Q+d2BLWuubmBZwy9jJ+la
LPD/9VgwYzIYLL/tes3tEvOYpWnVPET9e2YAib0AJss3IJtYFIIIsE9tWpiUlvnw
`protect END_PROTECTED
