`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0m45ID8npzCMlQJO0+ePGuTnbuWUjX+VH0zIBxK0wltvW2mG7liqhRMsIsHnlZhQ
CMmQ2+1sAsqYfZ+o6EfYTyw5N1vnUZJ8Z3UuLR8sY9Ooy6aP3iPgPWQ62zxK50K6
nVsWrj7aKpZVouQut0zXhbBBAK4I6nLysZplZdnOR51Fp5ippkk+N3nTYX91FWnF
ffpMBilcToL/1VtP+ny/Zhqp/l6KCHzSvr5LWiOL5cVyX/hPXq8k+erwo30xK+L9
NCvmDY3KtgwdCA0d/A6jKUCoWs/5FELKxFtmQFOP3lPfocm+5eKujatcn894qpWM
AboKLWcJezWuN8RkZ7xHFLSlmMKfJLeSbkvu55ZwJyb2thlgHOktZpOuX6dAZJ27
8zOSh3LzZp/RxiBLQXFjGS66iXXVUb8dzNy8YraBwbB2RaK2e5/L6P7z1WWVGnwo
9w6CpqA5kbXbxNyGaNx3AEtZy+dclSdv4cG/JMky5YxTx/MildO9+3ijssrpnIkX
`protect END_PROTECTED
