`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xasaeQnBdOH0NZuZ149DprZA/FZEMw4AgPRVsz7PrORbck5s+ZMyFVNn1ncFiTCE
Vy7wI2I5Q+ITgT1i6rUmdBfcoh19sp6R1MP7Ve/sq1a95HX9HIJTotNmoZV3eu3y
0+bWAy9yeco6A+Sam/ZsW17EWh8ALcze3C7wxvJXWErfFel3gPf/dlxUou9r9pr5
exKP0sNdor7AYwq0064hNVFRzgHLg5yiJ+uQWQfuk0zoBt/55XIk+hk+pNU5HyZX
EpAKZhqMS7UErL9ozKbee02QBG9e/IWfi1BRgajxheUIfESfyd4EXQS1d/n4AQsF
U1x2XkSsRCG8rzOyIgz55Ui6LYTVUcbVzEjIvJK+XnvvqCRyZ2ue3jMk6PzZchgd
rK7n8SPIXwX1glHdMw0mJtRCQsryDRf5cA9PU12c003Mjb+86pjPW3boNOxz+TtW
my8Lgghq090nOxCYZXZg+Jqce21WMQS8voeGxK/i0i2+qvOWLPv8z9BcbjRc89XH
`protect END_PROTECTED
