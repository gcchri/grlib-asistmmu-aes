`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fj/55Cj7Q6mXSAjSUkgCXx9gkyAnAKH487IFcRyMYRFWn9bY0eXf8uw/zgPjKVY0
QrFesu7OMMA8h1IlzV7zx0B9VVSUPOffgTVp3LQntVQxdS4Cwclr5+AFknTc6Ecj
Grgt2WRRCvoV7LyGHmDROamZW4lHMS2j6gJcySNzrMGNwpAcsY+D/LbZAqSqaV8b
BEHnVlaqX7ZP2ejVZlx7WwTcscr69CmY/V9X+yJBa8JnERnwmpncZagQ7HIJF+rs
`protect END_PROTECTED
