`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ulbNqAmMhRAZWNAFqVzG1jaroeZVKeHy1ATq1g0KCaRkRk21top4lV8k+0jtKhG
1Kawhj8U9CzUvjb+SivvNjnkdUHL/CnhSyPPNprDwWACuIGdZo/DCaklvqIAX+QW
eiPtQkLcSizl+vRyQBqjEBXFlRYQ4/VFt/EHKdO9yJma/dim54fbDrSrxwBE9AO2
x4H2PqlKgDu++Qjz1b7fmPCeuO3Pjw/ycENIsn14yr4aVQBw3IuT1RLlV98q3iqk
8s9A26aB88/AKXFWytIQaGK87tIB3eL5DlQ3CDU6phG4JjSSyC+JO/m1VBrSgoQP
XPuqzhnoOD/oYIecbxT5PxlnkHMWFqRT/MXHnEKq/W/Ij5Yrirwl6eTaUGArL0HJ
CTNPaMUb3wE+XpoiQc2Ru3RC5hysUHMVzUiVXTPqw1ypfjsXwdbipvRMNoLC5J/r
aaSXCH1Iuf0tqohliacVrf+hDQNgjLNwKd0Wjv3tUJbbNhcDiJJGNbQEM5CtLmxC
9VmEaCCj7BSQzE62cdxVkaYpGQ+wlMWQDqQI9Remps4YjquvPR5XC15IYfk5VQDL
wxb+PQfAh58J4sdM6g2+w/nBmJ/EEZ0APvUghJm366HxyVH2hf8BASM4j34B4RAq
B7CG0EHiGx7eLG7gesl8wienQf9Dt3cKa9RjScUe6cLO10nsS1Z6B1VlnO2S0Zxa
Fbe74mj57IoMOsCre0sCb9/VwggQyuHs26VSGp6hDKIn8nRGZ/xMHMthDma826/F
bTrFq6VIjUK7OSl36yUk8dNkhf0L69ppnFNeFRUwNPpwdcSapxr50GW1zu5dJL9h
zrdFIlZgPmjQ8yMzhxJwbcTw0AqY2jwx/Wd+cUIEdPcKLRjhMi12KxDyNoCmJMCG
/jsylLi/9lN8ECLtpJVuDXuAK+YObUxsZpQNtFinNqg4RCVyoYL+sNBWU44fr6WB
T1GwyDuoBZps46Cco01u5wc+v7FnoYzCyAyidKpXhw06/GqA2GYoaCN32xGmRvgs
zkcf5o8+jODxBZJhEW2yDuiLjcuJOBcryVEEtkQ1kCR8v+dAbi73Z//EOIRIZQ71
F0qnAaofbqpQgC/eO5EAmsdgraweW+G8qx/fwQ4NQCR0N05MFkuEn9klnjRFBs7E
zDYPE0I0OPDmuL6W91Iv3uXBCFhfreNICviF1hROJwnft25Y8f7z8UK69efI6CrY
bH8qGHqWKuhaSholBkAg02uo75mKOiilVlHke35g/V/hvgeN+MPQ/jc/+sW++bem
70UATAdaBXSJjAq2YElgRG8a81mZ9gVeU/kychCsrqY=
`protect END_PROTECTED
