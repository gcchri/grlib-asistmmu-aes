`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6lAquKNJhIWY5rWNQVi8WZmEFV6eTel+BFYo5o4Ko0DUy3kaiayvzFuFlL71p0+Z
oVEmjf7iXfXaKKojg8tj6U6TVMBmqrcwEmNht3Y3iRuLxXz5VjYxWXzscICOEblx
ZiVSuqOYqjbFk/WThzZCtt8EfCzyAOgJYbJiVFe4jennSGUm04AG5IxEr8EfpBby
rg8HMLDxwxNwQNTFn/B6+/DnKXRll+JxyGb+rPculvZOsLYSL+gorB9D48SC6wXZ
4jejlC74kLL9kOFuUkBpjT5RwArLZrrQW/3OwOYQ79md8pJyCyP2M36gPGEZK3rp
m5dAsmzQh3GcziNeb++y7g+iaEbWYVbPGiGHAe1zhxwfH4kz8mTAh6Uahv4t3JVg
hHC/jYRP2ojLLEbX+/x5FTG+3Gw5UehWvIpd8ItYbHHekm7vzVI78c2h+v6I3MYc
ztHMwwHNZcUnBxh21+2CSgYPy3//Y8O+vwZqrTNwy9rsAnUWavaF4HSByRBdJ2+i
PRD+tHt3NkakYVK9fG9K7Cf8yiA7eQWgpuTIWeA7O3yZYla5CD9Ke+sVUN0X6kgU
ovS494/YcEMI2eUWFIMDxKHxQjUQYMwPRLmTTtPR4JR6PmVmg6c1/7DTjRru4MPd
7Uv4qIB5DuB3H7y0iZWfPyvB+dI/LTN/iCUMSVVUR0nX8j1NFWlMVY6zJDtIIEL1
knT/ON4dV7+0cRMj47ZVrh9hwe8qjs+A4wogJAJ8OQLjaHTyT5Ob6MCD9XLSqEEP
iQwhacjnJhNDsSEOoyLmWyAkKvE3vL2RjjM10KOXXjfXBXAYKwuOpA+BVCZiey/3
Uan/qF7bWRPNPOsaG5kpOZ1Ag5/oR2ktBx6/+lrRXe0sCvEXVKROTuf3z6ikVCRD
ALzf5v7Ekp1MrCrux0at2aEcDJAdtxiZJ+z4n+ZS8CG4AfhhTfsSPN78zuw5Z89+
lWSoRZgmWscG1V4bKK6eDI5qGUtQur0e54lQUS4YV37xJY0vuI8X4uQMjuZ3PQ1W
Zqe/wrdpwQs6/3TVjwddr1m5aiVzwKXKUMwv9tBQ/VQqRbf4B7Y1d6mtgGGt9f4N
CBXipuUEV89o9D/Ha/E8IaWieJqjojUsTgMJKkBNVYY=
`protect END_PROTECTED
