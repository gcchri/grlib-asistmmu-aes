`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IidcVXBbso7n9lHfxaK7UGlj00UM176O9Q1TzipBNJsS5ucjn4733xgevzCdw0o5
S0/jWVchXtaL2Iqy0Iuz9K6Cvpl2TmQRs1+xcYPvKMP96E3ZePaTl7mFlH9afQoQ
kcug/6YrB3nCCMJswaCwkNVOL+SuK24HfT4ACJS3+4iyFn/mzrERMw0PxnXR2bXI
G+l6KJTD1h99mIi2bJIj+bFR+eM0l3EEQhylIKi15UIsDFP+cRr6anVaWi6Ks12b
EbnGCwolSAhs7H59uBRRy5c231i5m86F9SM1/jzZDi4wbZVVL3zNS3i+Geo9RB2C
dSOCGXk9NmgYznGGSNS457r27TYi5wtmxAmk32euAuo=
`protect END_PROTECTED
