`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/i7PuSq8IYAvufO5y0myBSGg5CxflwaWqGbr96poUiO0Ax2VgQN0XzUlR3NVQfMQ
VRVH/eVtr1vEf6Jmd+BZPVzZMhYIDnp1c/hcnDVmU7COdCouFE7+pposeBTcokWf
dRthdJTkOMMcvyESEMqFkJ9Eg3LWg4FBu+m8YMlVgsqXxi4I4fIR6R+szYhsAHNb
qAUoXwJInGptIRSnnqXSY62E3H2KKE5465/L7DfNgSnyYwPt3gL5Addqa8XPY46b
IBDw6eruQO/ZrI7Xp9jss56jAwvf73nI2T/jKU9ivHVtSnsoAA0EbAyuAtSSR8u7
HfLFXttBbZ0Tj30hkzXwLfHUE19dkw146LfGvI+XrGZRthGkO2MJ1omIZpxNVHAu
BOWjW9R6YVdFuKmvkMTXk05KnQ5IzHEadnvBJiLXxNgeC71BTzD4+4yUAAP0nwPN
dZWE/1KCepFOa8UXOuOTLAzqMQ58pQpFnglnPyUp2xc1fm8X17nFJrsDEiZMzm0Q
0VdmblENf+02Z6tnMxd7cM/slhZe0d5ny0HMHDhKgKee2D2+z4pyCAauCr63tH/7
bxuVkCIUjEUSp3c2ZPQerG1kUqNpx4HRpHC1+2YAONEiJCW7SFJCOLeRYvqHzQm1
Lk7A6yftwjfeLTXfKXDzQvMSvgX37fRLpfB1KIa7D/7nTg69feESj4agBrf75Z+u
l8anqkBW93PUKgIyCy0zJQ==
`protect END_PROTECTED
