`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8X3i/eb5SsqZHt0flf1tVMmk/4j/e6Dm/83654hhg8iaM10MRNspH8/Xt+4Ue0/
YOMBH9SAcXg6DDEj6XdFVjkUzmkIBMvdoN0PDJY1h40RIBpFu7NsZxX0XlbblQ+4
JlZRWUL603CU6fTmzID7hmZxv9gw9/cxnDFLDViKp3KuAJ53hDHV5NdU9URWcm2u
iQBC+zfeL2PqOk6qvfciSeZBaxnF1op6bIuD91QsCa8V+u8slKvhiF5WGHsFsBM5
JfMHsCwQQ6vGXqRkldm/1VM5TK7wHr5fhG78WQS2OJ/aZ9K/BTnlMH6l6P/jlP1x
BoRWs2G5DVqKSvh6YFhpMb+Mr2I1b0fg44iJZxbwqfFW0JFXJcO3Xr17KOP4Z0Yn
dHKKuA1te48uLLgjs3+xC8S1kbnOo5FkQX/GXxhT3RgnsV+OUfXjw5Dy/l8zaXyS
bBvPf7irvOIdJ7AzsnusxpWW741RC0DU69w1zPXckHU2nWIzTRK4QL1Ud9UNuBvL
5t28r9+rAFeHwsRQxXFI4WBa9mxuQCJHJa429ZAS7WY15sNXhZlA/4VqeBX3JeO4
e8BKeNBAUQW/ATZ28dm1qYyMDyInDbTToYUUF0z9IKgeP733fkPTWjUKf7B8dJ1S
/jHPoAIYM0z3rawxrM7R9bTCNPHnbVlLwZS5zXp2ypNO9aJszhu9k3k5su/fztRz
Q6b4qTz16XngFCGymU8I1cn7r/hRP+HlbMphmyjmW64QaKaxT8nQXi+/KWzdY9iP
nCNQu5IjaMXAxamgN5PPMotyF+lxgl6Ccrn4Dw3wIoZq6M6jMf5swTx7sjp93MRe
3wNukYz+XtoJsyrR9pBG1EubmmgRR2nbeYR/SPvyvE7l36OO5k5QdxTr7F4aUN28
fkqGyzZbYJLoq/bx6rnIdXyETngmDog+Ka90LHoIyj9VdhW3ArBdoTvwLBiSMMIa
7ybwex7EUPW7cobMAf1MhrRcFAEM9mP7lzPK4BXKqMk7Sc5lHkPE5j2gz0UqrLum
2Wt7bTQXAfUOmTldgYxDs2Y17uifhKmlAX3fQIF5Ufp8HhCn1iRZsXsasYc71jiX
l3t1OYg5vDB2r5gSUI1stGIscTM2JzE1s0/tz5oAbdT3D6JLjLfEvsxGZmWgze9w
OGf0U8kaHHSazJzG772fKtSruk8naRGxTkh1o/Fg8sG03wtiGTtuvBC0uhWW7Tbh
xrCntrdrSZeSMvvuAtpIKD/vEH+mddkGZJRIIPpqAFMaRJ5tmoRMUFMq+PAfr2Uf
H1//PBXuH80g6JfrLebIukKddFyzILeh3dkl3V4ayng1jYiGJs4G8W6M2Yi4z7me
/iyTPvMh2Utg4JsC5IlbxuKaImqEWGsRzO5kAieT6o46up2hLK9IkzeUX4VQDtBO
SmsgsSa2LuPrAuM92jFORk64okPD/RN4Nzppaxl3GW+QIppfaasjmkGliCk1Z7xB
wWbnb69kbHy2UnrPHdUwH66UuQ0luhtExfxdCHh02Vp6Si28S18/u8nttCD2Y03s
eMyAdGPSTMFjybAKRPV4T8r4chzLmxVFAvoE+GbgfqxsluqrNn8HVXrf4UjVU71m
ZIgYiS3YMbxBpU7CbpU3tnoqkv+SPJ3D417Piy0hXHEvY1hxlCaE4cr29xvPv7tK
8ma0QfJ0P+N5ducM/+8dWwc7EktGaw8rUSm/Sa44vYnoEJNnNeCvoQleSRaAoto0
q5bS1tx6om3VLH+S316i5vi4YLf/BDv5J2AGuVJNXZ+lG93WAgVI6/3x2ckRcFgn
HlQEOYubc6DKu6aWTP1cIBMX2uMTrNLEgvFw0RQJR3EZrHo2NkCSzcQPSbibM3pp
+iWM0AmY5NqyGl0zwlS8zqOHwAZ7SmfT5Ffw7/rBCrI2nDRPfdu92CRL9EOAnlVD
VJWODA/zHM43X4eagy9VXZ8Ml91/0wfarm9EtJM+M+PZTHVDfNbNi8U127mmgzoK
TPQAfOgvsaVhzF7feYFKr80G81x7THnnta2N0OlOkOsXdIcfFW5ON7Ebpx8+Strq
GbQbDc5VBMDAeqw6zc2QgGKQCyk8XcYk/ZLOkYIYF+ywCNBIV5jljAQuXFteT3Z8
u7/AIVlfmnP9px4sjPAQjHsYrqCbBaz3BVfGmZ4/UpIoZO4Yxvy2yjsv9R7rLcjq
XGFmwmPKRN7UZTj7BZfjn6UYj5Xkjo93pNU8HXMCmgEccPnNtqdisSouH8n/a+jG
zSN8FG+fs6MRhDW2tUZbntpsujM1RE5QkgVOoOB8wdMzDZNyQHY//vPF8l2oeUis
ss6A8/EUOOiJUvyx/UxLt924/jg8giZ/MAHrkQHp1Sh2K+h4SVJYN9f+6364YTta
MEfJvM/3KjFnsAigKxYiOTvLCIVEUFso5QakRQ9FFRBldgVtsLBa2EuutGeIcg05
kMLriTQ/Os4kcs/Yc2rIqNUwrkVxJMLmleumZhrbmDFBf+m+ftr3rvt07luDcyfl
BbMTGANmvSF7Y+cnJYRL2TlJfcwvIO77cBOLo6VIxYilwVCunzDIUvVl1mW9H2kj
DCql5Jwn5cm7u3s/7xUkgXWtEb8HPjx7j7uIlJnFCVHxYJb9UF7e+2igZdD+5sOV
xhcCA009ca7WBbBXLo1SBalnMhvPxE7nXJ/oFAi6mOdb33P0451hUyh+SiUS1zjv
cy0xGzSK4Zf8SCWRzxvNlX4uSkimaStaotAKb6gexSUNmYB6CZer/ArffxA8khoa
kN9A4nk62eTA7sMqFnYvH5DED9sx3fOSKRaAYbXlbszkCD4yphhMOOALU3xDGI/1
3k325NOBo9d04/ZrBuC4ghN2QUoZHGdIPrZHROCYR14H2oDA+uoKsSImQf5/8+gl
HwUkyAnj8V+9je3U70Khpky1QI+3qpQS2Oo8xtm/KPXlDpUe7bDZYlP77/0xoTs8
TLBHpRmmTIPaK/fl0LSw35KmVnC0Kh2R8RiIY29D1Aea/tHavlYcb6XRO/f/EOAm
ZEgmVP7VYk2xPpvZW6ALir3Ryr9Q22KYuFGSkFqd1k7dVcGrSxnAAHhk8DR6jx/f
R1crCSxi1aPFq11i017+0yRP0s8gRRrvJ+j4eog0qEua622/tSpiF0EGyTIAk6GO
GkgMLUVhecCI+fvRWG0V28YyszqRrf2MtoYQBAySyOkKVRxQ+5ELu3v/vB3FVZUe
7IK+L7lSoZUciHszA2jIoeU/tQbSuqaKpIyCYf/RP3hjwL6RaTyj9LNCEUavV1H8
B4BjKu/jNhir2XMqu7pYJgEJqRCtgI6Hprd4mi4dtcp3Y3mhDqwoI8GmASRoctFc
PEjqZ57qc2GfFM2MFSrnU+ZT15VblujoAlQdOvxjSEWZxxJ5e3P/EOogwgeqhPC5
Su2bjXGydu//pjzwz/cgtYugotO+edKnqSR6BKeDMKUvFnoiX2ToGLM7s8QWZl/X
vJSLH/uBiw4/13C4SQyRSr3CT0FyROdYNeGpLqQsNXRw40NY0wTtvN+y7/2ML+Kr
R4Ud1KaV0wOV3nLyKFBItbu8XcnP4RvXtXGjMJzQF3t754PY0kMSGy80Ue2nK3x2
XpOZR2B3/kN5AlKpSIQEU4JngMCj0BAL5w/P/snT0lX/wV51WvsJvaUYTW5n1ZNV
BuV6AANKqEjXEfm7G1Up7cPdC5Xm4FruQlnnKtiBhvBqEsRZ1PivG9uMmOmDggH3
XEd4em2zM3Jkv0Tdo8MsSfMlh+ON5bHZxxs9J7HFBfCCx+gIl6fGZE0499huAXaz
sbZ0N7FTQRx7n2nwNoNaClCFBwReWQydRndzBArtu0x3283MQFnptYMM8WFzElDM
XuA2N41Off6gjN3V61LBelJTaAW8vTPFswZ7FC7VF+uUx1otTLueCOqxZTv7z1I8
RwCHGB1nbp2LTOpKF86ek3cZI+MW2b74Cd0/YOfRde44QyZJJKrDahpx9zeXw6gv
F9zNT2laOOGo0leEy5fBJFn+AP/QqEYFvBWMsw6BaU80x58H3A0Tj2AED3xKd7As
6IN175p73szIWIMkiQTtsb+q+BcYkFQthwzbQ5pU13qUCV8c8Fv21XYib4A3dT8s
sA+QjLDqfEwTbvrpCDfSKRNmhO9yq49qrLyYL3211/+m+l7CJaclMvav8Dg13qqM
V8MwubQ/eV37ANYvEPnZYGRWGahS/lulgpTAJdQkGCE0ISP/uUShzh9RHLVSfWQ1
OwRRIHyRCBtCwmaw05sKZOezNPUcMmBEYPMbx1g3oSuOprNnYN0DrAdW00m7yzc6
UM60b7LqXQ7LKCb4WXqsddJMP0GnoN9+NRV5hSkbGpCHCzasid3TyTv+kpDruZJq
k7nTEwyLgNKnZeTS/+lOvxEuyiwGFFvuIyhtk1KsqZCIDpu5zOs4Sp0yV6bk1nfy
QNEMQcLwG7m44SXGcoLO6s4P6lZ5+bzFgtcaapR8bFZ6Uvbd4aE3i40UaCmdzd93
nWCzJlveJ/fZPhWnC5WulPsc4eklofXwpLEQwt4PuMEQqYuURWgLVyLkzG1EoSDS
RofO/nDlPMbEbh646iVKG5KdG9o9epuBFg5NX/mNezoyDlEdg0rnl6D70B+pBj9H
dzcIAQ58cED2a/9HJrRTqFecfnqe7e7mCadKA3x2Xd/nXRBzuKROtY9rEAjM9LAP
NickSkDNuhrT0FLpR37s2laeQDKuyZBV4HHjjcA67rcV1iUG+rnI4VwWviy7OQ2V
CkA+ODt85VYzv8d9jTC0V3EXdIneNZZbOCIDT0nAcf+Oa3U4Q8ykaMBCtsp8byfB
aGWqt8tEbc6T+daj6joVhH5fJ0Ef213IQXOpl+relX2mLXtMqEYi3ChSag+Z3LYZ
vlijmQHc8NWE3E65NjTC4WLWT71NdY/1GQqyk4GogV6F7s4rCzyjhdQxdOCR/J5w
`protect END_PROTECTED
