`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eDMZSoZabEAEinniHZ9hjPTujIEAX8FkVlktncg9SRJo/SokUnUz47NKHq1U6N6L
Qhj4WEredWls8KmMnJoX7dEsfOlXQOUyowYALpNO+9D3HDX0pcp4AhIOD+ofX69z
8HwVBSAFFwofW6Wz2U8JB9tPRt1gp7tYF/Vtfdf2T66xVMfIzyalxwOIi18ICObK
r0CLLh38zK1mkKOafsoHWDbbpl8eBpYXdLezYhqPo/qVEPu7dI0ytAZCoNgmpgQT
jUvsJ0sIO1tO0b2F2c/tv68B16UPnBV6SHjg0AFf3m29BFK0K7kQ4Ab5uqRHPFPd
0YlykfU9A9PSTqMcSnHARR2z5cVkO1b4+v91727lncpGbY3xuxF/w2hMELdAJZRX
0Osq3fu6+NI3Hi1kzw/GcAv+rvg9HIokWIxpcxr1w30xu9b+mCCbGvlfUkVeGObd
PGgfXOuommA+NGJTb/Z4G5anvcyNJ+OLydkKXFzxLb4=
`protect END_PROTECTED
