`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ov/dFmLZ8d1RdJ7BLbzMq3d0/odH0q+5xUuwvZsE0QpribNN/He8u2BjVoUQu+qU
YGNzyWfmG7AFXRtMfO3wJFCAN2H2u3WTV9rxdFw54IKr0GXo7+elP/X7F4zY2x0f
fN1NBmzseL0HYXuBJw3BYp/UDzFLAtSdvu9PI2Pmzp8LDAueZYM2pXLovaTemMdJ
pEXe00OU4xuWmzrqGPb7P2eWvz7szbQRXyt3+EOKi223NdPCOsD3gwFZm1yMWIjk
3X0LBTLuVN6Et/glt1X/Zkgbb66O9VI2UgP6dk7aABUfxKVxHVaZN5UgRBJMBDpr
EM8qZRKh8OHRwtdTyGMF+0UcKJkcjof0Pdhe4muHPNYvHQk2lZliQPVq+WzYIasC
jqiNYl9bbGse13agy1euNcdnAz3FmTTJ3UwHXd/cAl5fcVmfRGCg7Eya+mryf6uz
yLabEuv7s4RsFIwCVAW15pGDsR6SmjjfAlAgG1a7ZSk/ymbUOVWSDBbPyzewD23d
AS4DoQLbR04GeLmIprRuiWdyz+xPTNPBHV2ac/pnzDLbaM0cIu3B6VCfEdEIrOpu
s/+azgjGn0hD0MrZ2xv8I6YqQAPWErIMgOGshZvFdHWiBgSjbImgXTA89a23qoyn
MkpenAlDFyM2dfCKuKdQXQ==
`protect END_PROTECTED
