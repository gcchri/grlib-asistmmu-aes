`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OXVye8fPjygQymGpIeg/apKlH/PI/BEyCZZhH+NmGx6JrBNBtMCyTzNWGw6tIQ99
lK4U2Of2lEnRTv83tt6qDtHOeDpDPY1kaXI/PYbE50q3MKk/zhDyBRqGyl4Q68oH
mtw8dLbIHwrnnet7FFC4IOgfSYXV0Wrvm9Cyx+etiMrYI6yy0HzuOIyHRun5H1vJ
HcH8C3JFpekIMIb1KDkD37YhoHubrdPn9cNtPZgnj61CaP6xtzzkqPaCxaS0SszH
Y0LDgM7nv8OOMDzd6wG8xg==
`protect END_PROTECTED
