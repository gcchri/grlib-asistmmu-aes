`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMccY5cV/i0XsXwfvoZ+wXFftNeAOdyvC1aVzNeJg6LSTtVglWC21aR6aZB1D05l
bYOOR+APU8Pb34+p0/UoFpO1cHNZBCPXrlIq5kiBcA8huPUjTn2o65lQyz6ccgta
12/g/Qz9sxC3V1eMumunPZcqHJKPLW+RtLA8hfrLyYq7bS8Ft8CCQscgrJa/5bM6
blWe5g2gwfQ4UQltJ+LEVHVE/5HZCrlR2egxeVzhJvx3c0sRoloEeOKkPDKkvgln
eyQXcVDPSneKlFMAJKEf9Q==
`protect END_PROTECTED
