`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UShkATYuX8mgk8jbEupCyeNNSrzl2F6Sy2E2phNb+cL7Qn/9faIvkvNNdK3qxVdQ
MHPJWfnPz8gMTZEvbmDr+k+joKpL8eOR+14MPb18C1dV6qjsx2emHxB6zUgFTyPz
czLofwDUQ0WQA3g/Swj6dXZT51FJqJ+ioRq8CLYuhT87KgsW9rNSAmhmibeOYduC
OMlht8+le0B99NL1BFmbuBkZDiZ/gwIU0hOO3RaV6IBfI0wnKgl2EBA9RLIJCW74
cStHZhs5cfdemiI22hxBJpH2s3yK0Xr/BYv46z4Po/wMBuQ+PXURDvvSmsPl5XN2
8mVwb5nFyneXoYXhMUk5wpcd7FrruMNbHLYXaKM/MztgTJuvUsdYc74sNJn4CTfk
aaXKcvVrwgHxUYs2PhtAmAT7kZh6EBv0hXn5P0G54XssjhGE+Y6ukmFg171QJSP7
CuO2QMUO9SCgyR0OsYpkiEbNL0lYw5DmTIZSOiISErAdA3OQp8sBmysBO7id1jXn
bpl7aDMRm1r7otEE16CTkXa0cEG7F1XiDXP7sWHj/YUy6bJk20S8kRGapfMEI67f
0ry+/vztRQWN4pQZVKniezie93mHt7MsB27aI4huQCW+PWV/4BSYdodmHYriHJzE
jbnvwnpStW65hmLflhenJfjUMff/3/A04ky+EpT+ViYBWrfM+uK7wgWDCQz9R1XH
`protect END_PROTECTED
