`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fX+KjmI18JEiI7dAnVFMfoKp1kPJ8YXMnnKhbXv1lhdS5gei7RaacSjU0fN2cc88
BgNK5v6FEm6frq7rNjEZXXGWjJ0TpRiO/eXhV8HpgbnFG21RP6i9Uaj1kB+Ry6sR
eeAuU5jJHikGrUKju27ohWsNGDEOuxzYf3O0X4zXpWYVLAXbg7RgpcMJCE9ncCyF
D2wcDjLxGuA8+3gZKLhVvclnOXNjd49L7DCf3B1Tq3c9CskbuUWQVLvHIyrwFd2b
clLS/Bm5NcJtdM3V4UI/Mgp/NgjGvIet3P7qIqv3r9sxj8ts0qc7+y61y0Lld0y1
Ya0HxC0g/hBzGVdr6dZsuJmMQ3ZXkgSc2cAzzwiicVmrV7Etjch1xKYq+uIJEmgl
CwpWiVq5vRfzQ4hcBHfOijVl3ayxXoOUlXUd3SYPbYYU07R9IdsUp2dAu0H+GYAQ
`protect END_PROTECTED
