`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MtOOaeoGdhefjFOZ0dP00a1HZ2twqr3ITR49nCxOJssreAlEHxOTOkZDbw/gUj0B
mlp5CivnXt6JdUDttMO1Ysi7YeCT3CuhJmdKK2Qf1xpcjhmaIH+yc4qreWDIuNdA
7LFbuuT3kxwnTzL0uJFVa3M6AsNoGNSJvd4BI1LMId2UVPVGZOxEMuEpXeYlfrEK
443F6a4i5I2PfDFsyc0pagG0FmuOrpc93CgkiqnlT5If+q8SZItcwNLPrguwJHAF
huwM6aaUgFdtAYfH33vq2g==
`protect END_PROTECTED
