`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yjvRv9pg2Vkt20vgSIwMLXj2KP0w7s2TDww+vXiUORUAj+FSFRWxcEgFU/jKrc9w
iltYopPfa60QMRnEoajAMUsEPXNML98STr6Si1v012mp5WMvdK81UZRw01DkCUon
s6vXZzJfFLMx+gkKwmFeJvkSJGMOn9bd3uTpVAj1TabDP6iijoxtnp4gwlYiOaO9
Bj//28keSBO0RpBH4zRotckObxd+Zsy9R+x6OIPcE+pCDLEbJgUmt0u31thKKw7/
N4rFjIA4pAJKBV/lXRb/1cQ2vVxxKsdBMV/wpKxO+liLELu171/glUzv67I0njW1
mE0KiixCGBCYpgDPae86KIsTmi/xxrnjyi/7kydXxpUuezpGMTYCNMRV6A1khygy
WjT6DnhPGxpn1CPHhv23oWfTvgwJR/3r/3XTFibZZLm6vc8vdfIl28dOxNMHIpOx
r3h7M8FoHFLabtdat91Oy1InBA/gO6+OtLUg3yVJbqPmkDKA1yPlLhV6W5cxC+34
J4rRv7gYypohgBlyH07y72nFwguHc0OWblNwuIkVka33hBkmIbCXZk33ljHpr7jK
502+jaryNnN+df787Qvquii5WJtmewfGLK9mwLlrp8D1ljOZf7MDjz8Vm9tofrSF
eTJwoTm5DgjuDP0Yx3AfEw==
`protect END_PROTECTED
