`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kN0AWTI01XYDr9Rd7ymmYsh1GGwQiRfzUk0W4DDEddkVE+Hj+AfN5VYNhIucwjKs
3N9EZz5XeR2Yyw47nHjYXktKPgBwnSFJQAC47LXeMFHJ45JKMfprtGgt+8cIZQHY
5xRG+bKD0OLtRE4i3MT9MaJNmqAqIL0Aoqh/ppVzXNVp2Vm7S3EMaPB8pmQoSz/g
gJIw2z8AoWyuNowTv3zKOVK3dzTXnLEEHFz1jImu0VBRvN1jjWtpz1VMUe4Ej4PX
dZwD20Wo6ZQUmF8QIskm6Nfa0CVL+QX6aVg5vLorh7US/8YOIKHdy3iRw8SnrZaP
E7dkZGlSux2Ne8cesEIgBQ==
`protect END_PROTECTED
