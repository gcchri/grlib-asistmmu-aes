`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/voVsHRGGeshbghg+y1U6ANWsOEy+tIj5m0qedunB9Re0PmynCGAiBGKNaq2B/p
8z8rmEK6G73UtRcY/eBNdXsfbVnuReHr+66tIWz238KYyo/fy3WU+OTKZn2JreMd
O5HXWG/cUxg5wx8KvZ5xs/t0ZbtXEEKkLV3/GJOslOiX7cXusAUPfNwzY8u6Ou7j
ZU0dDmEMgxbOBa7jLORfVqgz/yF2wZtv/HDytnb3ObIVJeo09BYOuMu3L5lE4fOL
yEN2t5xhl7zRVW8AQZxL0NWU//exRbEGOgKVG7mjAY1Ig7RPdNIWw1lesi2SJ/YM
WlKk8inoG9ucSjnG0Jc24WpV5FaN7/EPJt/8/SWBUhBKoqQsMF+cVNRncMYsnjyX
Lr5Ofe3Hs+zgasiCeSr16Lrz8q6E78xl0Rx7ZyJMtVVlKjdcq8wUZYu1P0S8+f+U
RxE6jva9HSKWquHLHie4/aZId9W1yFALYX0tPXAxy/1M8ctyAiI2QHWX0tZAToaE
iAzDcRD7UGFtrStibIVyKJkVNogasiX+5rxZMckp1qQ=
`protect END_PROTECTED
