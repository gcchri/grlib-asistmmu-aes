`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SbJzeg7iDsC8G5FP6ZDsBmMAPSrMfMpMHBepWOFdB6LLfb6eB1cPulSXLvRaJBPC
JNdWxkg3kVz+oeOyLSRtrZIaUYKTogOhCDZ92RuIMvu/rJJb7+0FTkOf5hjMhTmb
DNN3Hs3aesTrozh0QvtQeR/hYFf0p1+X76/r4hsU6Y7q/9yvbfvJvqHW9tAUQEMX
1ywtRmvQiAM/ROqCnj8ExBLcSziBB6UfG1mTjZF8YDOinjABU+hPi3cIUCZp4yBZ
qNUhw5rSZeIDb6eU7USAP4T9gyXbAsJbdpKpjAv5RUdWZXT6Tbp8z+sKMOlX5ObS
R58tq7VedNHQ+Xql+FYWER4auw9orq4WEKlU5opAMV3q19FwHjB5a+TH1EKZbzIX
NsGAIE22oFnioZdgFJUVVxwW7un/dtdmuAwdANzPdeGRFkLndN0SgFsAJkhrHKgg
qpSQ6vi4NJqKtm6NYmuV+48Ybyz4TpVsSwwXZ8sf26b0kxTdjWameeB5B8lGe2zy
SS6hNyRGdjYXU0jhRdp6Ue+rYSRgCKEQsTFFsd8UsBO2fEDgdlKJ/GSNtZkVCZ1S
5e/zCXPcQORH53I/W4v+zPUJup+fdX7DgFBoa2FptdyF2cGg/JpaOLjmez+z9SN7
/kFBwVeFOmyKoDCgDxrv8s5ZC14AJ2Kv6oe6XtKnKCU7lnSwH99miblIpzC857jJ
F7GDYHFDJYdSW2b5ETvTQQ4y9JripypW0i3OCtH11mqhH7nCtcwpvdDHZ8/+sckd
ukWwN318ggYXgnMDMnDYsWY/CUVghMobOtsQS+1LMnQ=
`protect END_PROTECTED
