`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7gnsNugGWrk5YcXFjY8LGJvD1c5KcCwnxoIovbke494Q0Y2G8ol1Fvo7jk1ODlMF
yEBleHVPAadSV46C7VR85iB2hnOprnSiNGfOs/H6mzh+r4Uw7sDeXsEC4h1RUHXA
AdFylMjO0dAb/KzPB+MsFYGv5KLFl3jK7ggrum2oUmj2Fnh9Ze5+pMCDlid8MGIo
RA3PUKKhg05lRfH4NtOglwqwwG1SHK3uZcWq8oa5isjsMkJ8omYzEY4yzZfyuWem
z/uJhejKsfoEugLxCMnsDgZ3517oZ6zsCLu7gjooVql7/Mhj1MDyGocjQxAJKQLs
RyElxpgPyzeHNoK/L3eGVurIvtvDbxaXiYA3022e/cwdCwcpJlCHYSS7RnRY+jUi
m72dIRC7FoUtf7+ly72Z7qHh01OORdIjEjo7ipi34iNTWlXooahXy20PlqcOw7AF
rKNdJIOnQxiBxwa3/lY0lWM65VsnE6ApNI4UoRoIrxs=
`protect END_PROTECTED
