`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfNiy0zZNKGjlPD8/62KjoOsmxFwBVPzmmebbDKcYVxO4wyX3I9tRfWD2NKpTcdx
NPpHka2EwkiotyPJhb/zlVrH3gzuDbuSDFRnqYnmYNwIWneDFh1PaRWE1fKps9a/
Pezkbdp4iCY8q52s5p6ZP1UhGU+g8yyZmCO1GC79C9fdy0ygjoXM19e5IDQwN3Db
ddlyKv2ECwvQsVNro/Me6Vp5kn6yQIajU/jMeYqzd+x/TNi9Jou472kNfK7jvcfJ
Lme9r9HtJMM69Nvj/ECZRWN5rBMMO2OyjLdQfL0iyStwcRPSNWtfoWceEOr53NFx
AVwZcvFqI7nASlh983TVaw==
`protect END_PROTECTED
