`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nv29aAEUXsQsMKu+VKv8qUThP2jUc6kTvDqGtC3sdZ9eNvs4yXNEKRHtEaRLemk
aledvuhdta8ghzyacRNZkMttwE15EMrlNp67N8OF563o86QuYRuqmgDmjKKIqJrE
hNPzqZOJPbdXOleJgL9BnwF6MM+k+FcWCzyiDoVBYPZvIAOjpwwpOzSyEzNppjEO
Jc39jRQc7bllhKnWjiVTT3KWfpkTMunSREojsJP4zjOT1NvKqMqb4EqF8V6FGm2R
kmFJgsw8ZekLxRxqktpn6/8EN4hwIFDlHQa1PVat7tOeguMDV6QYtyJgCxMzbOyg
kOwNnlQQTHOOgJD7qRSIBbiP27r3Nf3Sbvcyr5Lgsho=
`protect END_PROTECTED
