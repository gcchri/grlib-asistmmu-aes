`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AtsUl7GLjidjWm3N5/wgp56q8Kkwc0ypD1CcOCb0DihnTbDoPzRo7KuufKmxGcGq
sr1pxDGFMO78KcS6SPRZJx82Vt1kbGsEO3bYht5MFSGOgLXhKTb8/fyordf9dJuR
bGcOUR3jEnW2SueQEmyRXZqP3bAImi6HpgKBNexDKfgg92CfYV1jI1BbJFpEXpuT
eknITTBjMh/Tk+55hyE0iyXMJHZarRcEpMGwhvfBQTqfdLq3SvTukVfNNAuHDcWI
H2keOrcUY2BJ3KKvA+bd4nR48Lv7DjXWKAgBdbqO0RP5ff2gGc8EjeO5bYrIByo+
+n//Eu/+LaACgnw537boP8XMbNaPKWl4MjO2X7yj23t4aIYrvz/VotUq35P/p/Ma
WdeBThlJaS8NLVp0jG5Y+PvVwOqlpzAOyKVHDy8mLYUWiWTkTlh3UqWVWMfM9pIO
6lqThLTbQDrcss1kKFC80GiHVfYiSdq12HvNy5Is1recxXTuYin82jiq4LOS5m2v
`protect END_PROTECTED
