`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jOrPPy5sK/i38MyA9avIElvNIXkqRZQ5d2kWur0uvkzwbbAEe/zMqtKYHIpV6JVM
BTgtgqaGX5aD9Fe9omw5RSzhd7hZ8EcBItqRLQDwolChtlDOQdjWKxbaBgCQkTj6
AKktXZroHHePUfmWnPyj7pp0pJmKkH4e6BN4C6wzR0EORe7bmjOa4Hf3tSBByLmh
xNOIH6zylU5Yn2LEHBd0o6wAELJHWtPzMKBaD+RUf33NGPKEHjwliu1mUvayvU+O
6OVdRNIcVI4saAQypHo3MnI0y1qEecYWrHgHR2aSb3mEy6E/7YcHihqHCbdFsdQQ
Hx8CR5+I9JJe0kWbxf06il288Osyvd8hafxWfpEuv1kJnMmuZVv8Zh6KR+isF8gx
DsznMbKIMH9nlbkXidz1FsVowRbTYX6aiSixnAAD8qfVU6yEEKKtFKjKgqy8H/Kh
Az53EygMnykD0IrK21uuJP2f/uyfAB5gu5E0nYmmk+ngXl4WIwLWlzuMLAVzGQQD
zZnZwxB8epUC2g9sCXpDud/EwTCxjpEpE8FdFBDqDfra1l1laaJC1ScnqPcm6fuh
I/pOZHYKGFRQ3MNUqrwx4g2AqaeaIALUuoa/EP8P/Aq+Qr9J+ruilEFfrGZ2OQac
nVL9it2Z1i+klrMBSrYqnIDU8J1+3dt/8TZQ4Q7qIwXXA+xjzlROvyeMM02RZUrX
mXf9+EUvqzU/W4LdTNNxaIf/lUzjqjyB3XRBiFLElbeUTQBWJHxLTyrUN5q0575/
hjLXuduECrF1CrXnVNz3GL6H8gdAwVNWVTKZ7j+/ovWQdG6hsrPPeIZz5Ej95nZo
0l3I8to2sgWdoQRyYSXAv4M1JQd17RxK83rkqn/CHrBZUwJ5CtQt2qeZ58BNPCYc
1ULCiGuDkLhJaoDhkcVOdqJddA65F02dVeC24R0LsK6prX0fdAKc/Z3FO7AVvBl4
VigTtrSL5M0XD04Wj7kyyBaWK/CAbUKxUf6wuI6qLqfIhBd7a06AaaDYRYQJyQ6Q
aQSEFlx4nGJlsxnhU65FfLlDoGDrlm5zwQL8rohoHBY467tKaq5JFL6II1AHpPwk
nmkhnjgMZcVcV/ES2SJoBSpWA/D+jugaQO+SzBlRbKmuBe64t/HwTuGn2730dFwa
p80QPieePVZCCs8617lu4+GDEP9Jg2Uhd1i6gJLkfmj+axoxvLT4jZSEZS0sAA5D
UVC6tcV4RzspkE7rhj9eDanS/xFsKEFVVjnktJ7abzbYnoT54i3Aneg31BkwCp9/
ByJKVO+R/RGhpqyUgWltyxcqfAAq1/ZdEoHnHqvuOxvF/okj/Du/7c1eN6aC3cdq
`protect END_PROTECTED
