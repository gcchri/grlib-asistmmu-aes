`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ThrZfo9PElFSWt1t8QBVeGKBsj2A2i+W1Af5kfirYR3XNk5KdR6jOrVgi1B0MXDA
zcQRo2a87cbi933+03poMfnE7S9eAk1pUJI/C1GaSp954LX/+kHNBooKHl0cUcur
jcdc/UTMTDBMo2bmF/5ehIQ4iruf9RYKTXw2bME9JJepi+FmypkGm1hOgjxegNDY
/YKV9nbiOJstYb9lajWdxKDXkgPXudrD9CXDhuzYyw6LOQtK2FvfdMwIFsZxnYSF
d3lOv8risR/PkT2YygHle4i8jxSmcztuiwahrFmb16mtoqeGnPbUZj/ikSYEdIJI
QxIdf/LkXNin2YUd7iFE8AocdOCGU6sT0B6ZEIn6kI+/cUxPiWSFBeMhzOn2VhEC
f6mo382BT2ghbV7PGCWrLEsU6inH3144lZRu+EH4eZ/NCQcfKCQm4surgaeGORmq
R/rsXNWCCrYUvXnzOSu1YIkJjP4IBwgXPiW6QN3IgNwiKkRjusDLLh7ea8neut8T
1b7LKd8/Oe7GMK7d34N8gyWw/N3QSCOIf4KnC7kYt4aznW3v3xapPNCkLHDPdWci
QfMcMz8Ny72eypav7hyWGuyyN4eykHJUogdtHmgKt56jm/Ln2QNu0pEx86DC+EUS
lx+wUQ/5RJ4l9pGMq7g/VQ==
`protect END_PROTECTED
