`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x6AzRPXT2FlbPJCVoYMEHpfOBIliUP3OoQXJfDA1v1aAiuFUVmZ+fmj1bwM9Pl4o
/2PPwOnbQM7bImWc2/W+JG9T+YRgcBdxC+KP1TOBLYVflDTE7J4eJS6qdb09Tmv9
chi3h+Uu251TaFVKs3sOBWu8lo/0t6OGwsIYYUDFkJzkaYbDi2NbW+2svXjFRSVf
RQxelUvThmTFWZU4hgBkHa6IMEOLa+nMjdPeekfDyiECQKdph3IaL8e2JuImf2WH
Klsx4k68Zc6A4yhrQLJ9HrT9Isqtwauxd9XMbo76M8fNFECVTgUF9DPy7mnZGXne
zQGdMUILjQ5nD9y8FBpBSVGe9iZL/SyGpfNcDWl6LzrJu5iJzq6aVpZGfl9FzaM9
I3ofYeFxIuBEXwRhS86BoxMDKt1BGf8S2hP/D79nssScvcNbgqh5EVZR27aYffEG
289aNVQK3nqAXuN4dbzGO9cz/6aCriVHAe4IuUGMD35qphsH49npC3z/j5Ws/5Jj
7lJfftBVrs0hWuV7krlb8mtLG6tz9jXCrpypCc7I3oWvqEPADoyu8JDAoTtRIkeC
`protect END_PROTECTED
