`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NoU8XN2oacoQCAKjdWZspJAUGaRibCJMO2N5MMODNWKVhe7lAeAuxvE/ypHhArk0
iETHuRDojSJ0B9Dy85k3xwZoHxPPpo4ZmssWe2N7CF6aH+XqDIhH0PxVVUUA8ZiJ
n3EBf/xTBhMI+RBuu2te4Z3tIkPaZ7NS/2U/K3HEi6n7ulnIv0eZb4upmdaXkEqM
3eG85wG4FhMohAkti2zlYfP14Bvk+x9x9gkGxUgq2XtDqeZF9VngBGHCdupnslXE
1QP3QPg6OElKMqfYaBv0/3JaKshqeiFaNJJQQTWpKGz7Jkg3j3+rlKNJnjQ0YxwE
sYM77N0y/klUBmYXA/HkwXQPq1pW2XpvrIpgrvKdyhHYGjJx8Fc9RTC3doGr2JW0
KTH/KIU+1DSDg002ivCXaIz5CB6/wrOHtvp81gi7iymT6NtD/RnJ+EMnmoKtacRl
d8JWUX8MPaLaOcjgNnxSHPNnzQrtAn4dDQFxAdlGxDhFulB6gQqUiKYq7A39cTCN
s0XbBXgQDvta50xUuDIGmySEFlfWrShMkv6htBaxzLWoNREI+DdJkMB/Ki4ct+NN
Sut0e3wwdS1+eE5NRzMtSPZPQ0kVbcTY/0XeOqMSewxXH6LfMBgcRPOHSKUkVt+t
aBBs2flqzIteoomw/zAJXgNY2g4CnEPuSyZa185gvlqScPKDzFIP3d2Ls4JQQuIZ
YV/O6Va/zxOt2+Jd81OeMhgTeZ8dFkpk0f4Z997h6hYhdJDSJfonTAk3Fl3sv6TH
g5ZaCpx1Hv+qCXs4uk7ye8Dvy5Km2dYzmCMDvc6d+Zkb7Qxk4rHJVgDA42Ss7han
Y3eLy9GyRtfT+t0UDtosnp155yt4Y7QgN/Di6m7mN/8orqhMQB0O40ob4z5bjz8u
20QAFmDMW96QtGOcJIOkOLuqF4UPe0ZjKUb78mE4Psx6sTRRPnhEX8qxO/C97lLV
OCpY5npMdoEzkC2RyM3ifOvvpCXNtLXJ1ORlmkE9dagd2tsDxenPxyakt+BWm3Zq
GTuXIgKuo5fZG4n9x+lImA2ijyH6UebdFRlFVxlOn/Zo8F2MTCeQ4/faqX4382vv
H112H9K/YhwOcRwcHyKeQTQ2zzwmbSFNSsKPB+4qqx/4rdYq7jK6hOS12qoQ+EWi
`protect END_PROTECTED
