`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EXnGV1Ito5qDfHqLka4yAmRkYcgAiqV3VNfEVnB0PsUzYDDpiZbWLz62Kl5F85TD
IwZqEV150pZYFQoeBQwh7v97rr7HWdRgvKtI2ZHIfsBhCNmTaCx0Lhxg0sryOuKF
iT6PgEWhoj/nzaBR9SBTYqmT6x78dCEWzo//trJJV9wGpmHbYTOacrAjMiBC1SDN
yY7dtFdeLVXUFSMf61f4wfhwnxsMrcOeuy2rpMRSOtROxU/kVNuewYJwa5AaOUGU
g2W6P+q6GfXa2jie0R/wnG0QWI0l0ZzI4h8FBeINJ+QTbfXuOB+7JJtAtmmGPQsx
kjhgy0Sg4kzwoaDDqKzt11SQpU3pVr5KSvXgcRGIIkrGklojC6pB977kBKgHlkSk
gAaecZEeF3ZnE8BZwliGkmnEu1QgoSwTxfJOVq4K3IuFFMC7J6CrJINyXj2e6eFb
w8rrPOwx31sA0rJNRfb6UQijllExdDypwMbEIzPHnBl3PFwE1SFc8blkjokEPHOm
beDgKf8FQKGk3pi4FM/HWDljKfFJbOcw+wdFhKdVqEf/kd+n+6GQlWT++7xuMSxA
chU8nC4Qvzd/qrKWm2mHc9aUfkBvW83xZzZDMoFwUl/BHf24RX/GoLtv4/sEzx2z
HbQdMzLoyBQSdXmqlCvdL4OjS8At6De2gtKEkwG2FbrZACs6O6NJg48aPMokbeKA
J24b9sDlywLdTTRhBfBWLH87TLAd1oIgpdSsuBv80mM98TQnvAe1iTgLdkLClIyp
ayFfB3ZlM1w+qn5y1DlDW9ojRuxuztOv2zGDphSurl+QMpGBu9eq1RjHgl4yuAtA
h6klhlHcU+Td1ao6f+o79wEnhgtxyQgmtLzxQtjfsjUVgZxpYCTnJQTCVGyJAftl
oY4B0xOY+Zyg49Bv1oe/dX2ZhrZ4fENbvO7/B1ZcU3X0UugrH3onXmO7T8sc74As
3znVeCbA6J1m29u2jk9c/x4yHGngqN1nQh08+zyskkXuzzl2qNGyDT4b9Aa7rIa7
814PTZqJp3t7AxZfBBMaemt1Tsgy0QA1gL2em15nr4/r7Sv8BqclxKN5Iswo09Qy
e4gemfKbIWRd21Rq0ADL14rMLE5CkSmR/Ii7lRN6aKVz8EnYJFUP2A3vc0enGjDi
AIssBccqcPzTuU8LPrEkIM/NCzPmEtqPlK8gBf77eHki6FX6pqWeR//7sB76SnIu
Oo4AQUcUWVW6AFJyUXkBHRBhr493ki8Mw7BM0zLoWQJTSOyEEfSG3qwy1TqcRPbL
jxgfP/2/GpOesSPxrsBWD5GlNWYcy4P004mY0zaSDgyMhbCV/CFNAES3rUC76e1U
s0EZHO2VoDN0PJud8DNAwhwKS3ph1WAJaIEe720P9fa5CdgAjqPUgR4b1JZZfjqa
eSXJYMg2iayFmhTFfQr9s2bd+bJpn02xn5FmAGFs93L/sMPjnO2+hBTiRclbNWI8
BZS+vexYaZRmhIwBnUnhHgbx8x6jmTkC4IGfrpiu8rR3/k/LQTBsD521beopDOyE
oEXOPrZLWH+R4xCexqB4WSEhRgFMbgI2QSb71K1X1xCde5OVOSNqgnECGysHiNT8
6av7VbA8iu3apfu+d7DIrXs6yjtMKwBT8R2ghyhwkXap3Yb2Jxo79aQO5GEdyIxY
HnQ8sWxZqA+8phopybwgboFcpu/zw8H0VbAzShZJuvat47X1WclIj9raZVf+kBms
Lqr+Z2o86GvlNBMcI+AaVu2UpIjv0RPl18r/761Fs/obMCMVATW/iDaQSdgFDDeD
y8WMjFSgOpW+SwQ4hrlOmmEBpuOS/x6mG3+bfOz9zbsI45R2lxtvMph+cNjbvPrk
UewZnuo2ERxs5Ihif+DtMM452L1hTlW8X2O3LWKTq67sp2Zsprn7ek5fRE8TkA1T
I5etIi3MMHPKxcS73tQTnTTlheDPxlL6HhN82YUHH/7od/ni426Z2mvtzZoBYLtb
AiFg8VFpFHIewftXhThed8A283UdzGDKU1jbg1tem/9ao99xzmEg/eFjRbqXUSQX
u+8Gn5lsmMF0AqOkJQJVn4uZQLpBFpY4NnegUuXOk5psT9nh5AvYY0DqRzBl7R8Y
Anc7FWCSb9Uzdnz4uRzZhlhRa2cxVeXJcFa2CH5Pw1N0Bs+p2fjqMn6C0kF35fxd
mQtcY+AKhz23yM0ldeoV/dBc9hfHWXvPKmyUuakyWZLwwuLVIn0Dhr6XNM3SeZOZ
x+JdZIGqXHe4RvalzZp9PsIxDPPkTTGRNYFOMh1+/krcNGqxVbX2sgle6IgY+q9r
Z0SbjR6IXMBVwkJDipCmlcgycbMBx2F7KngSQX1rLkvGXtnTdH8H69PkUYYH538N
QVEmmF7GATq8N52O3Pt36PHYgHmm2fOOejiEZj9COmqQUURtHPd6luD8x3CCI9DW
nkqnCpZdWhrUk1US169BS8AiqbXN51fOgxMMczK3xUYygXkmdhzsizzo0xLfYuuJ
fbFsdrvGNf8U2t+X5wekRNmxNlx38XxOAsrhS8DprjVjwCepfS8VnHJ5/owO4KHn
1Y0X5TK2svvoa/tFndLcavz462yemJXAkcu4AUt+xQFrWt7vqYNwGtbrbS4H/ADS
UTS91TDODRDDg/msAHg9yIUiF437pv/0pjArslQ1RJQ52YIaijVdYGJBartbuBWD
8QQvu1+2EA1md2JsAMfb2/peOs0IJ9iGAr8+KBz7/33yvB1OUrwASfnUFpikBc7B
Y89ne/QAxYu4a1LipT5NTZGkTzCdR5hRnmK2iWmuCn/aXhJ7SIHTkKazEv2bVAXW
fjDxxRVjj7QsKeeB7Km2dPhD3tHZVKkyYlxL5mIoJF9VcJjlLfO5y1N6ODpJ/NQ+
t92bW66ILWfOPR2mGkptkYxQV9mrY0QWMpu3unbjdosf5fpmZsb3mAvObS36SteC
gOcsV0+InCX5QVkvIis4MzjprBloaB+5Ycgyr2mq6eAfKNkDI9wdd1esckH6ntit
9usJyi/7zSysWsKRebxIUw0KP4O0AcuQpFCZVNxRRs1T2rLZyt02vs0Tcdu9joLu
8gWTE1D5IGWzup3+UAZRg+sy7FVBobQVyU7x41Iu8FK8FlyD7w61S079zxeCgaX2
qSaDFYTggi1HJCJAn/rtjVol2/r1Lb3kbDwh/nLAKpb/BtWlzaFiYSMEvNRlptIX
8EIFLuLJkAOAcfcpSdTe5v+Qsm15sPVXZ2WTWQpvt9H3PXgyZc6atcrnFO0nQYDl
4jwhiD+cGTQijTPpt5MrccEXZEw5Fiayc3YMCJ1ssD1hYltrC+K2fix4vIhPl5Fj
EYFtgbv1IQoE1tU0h6H8sNwvt5ZQlktCmgjJymT919qf4kghMnL7N6PZWut3neU5
v3CVr6C8ID1YsBHGoSpcqP1Xq3aq4zHNFxsRoebuqZN6foudhjkD4PkfOp3K1/AD
jIeQZKnUz5U59XGb82kSCQhUrew0e2B9xnTcATUhrzpPfBUXgURxIhQWtBBMTpsC
9iVwuZkXzOlCN4ek4Csg9Q==
`protect END_PROTECTED
