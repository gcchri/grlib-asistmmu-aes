`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYptfatpBX2GKlbtfZwEnSNZjqBAP5WfmgaIRonef4ZfIlx+KlnZ9EYo5jREFMwg
ReulI1WEse6wWB9sHpGeOzsJiVi3yWdP7HawRjJA/RtVoN+abECzUMC91UQvM7Ny
RyegCbI8wvZho6kOFE3mn76XSmmm78WCZnsELS4uscSMbkyMJxKGFVckdCrEOoth
5j8SZyaFDkomFiFd30KoGzCueLW7miZ5+hpslkmWp/JmENi58t4R2VcB0l6mMF5o
Y3JFlGKeoKgqGTaBJvZZjBuB5Jwb7XzIz+m2AZNcdNHTSJjfwffDNi0x2KF2eP22
lN9Bzcpk580YoY8qqfk0s3YAQBIR+kYvuHENOdou0QPLheUiR/9/bFM3LPOlRNhl
yWqrqRU5bhgU+Ab3nYJuJcYHeyYEpejOUJ2ilt5LqJkp4wHqFYNdG1+A20U4ZdRx
fJ9sWvE2EmbqV8hw4NPThOia+dvYdTsIhHsfSkws6nhHOagmyBJfxVh9USOJi3Ij
QRh3ivieKRDj7kGbQ9HFbsvGIS/HBFa0T8z7JAKJCM3GyXmHkP8ZhSkDLvOzUftW
tkAVCQ8sF8yAs5FXXYUZPP+xcSpz4vEiZr7b+aNfZSqVbjtOB0F0Dv3oJRMp4qjT
jAiktEvT/LgaRDLYRWm9vgFGgImmh0J8YoQKHzxeXfA=
`protect END_PROTECTED
