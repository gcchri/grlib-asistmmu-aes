`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3EVJ/FvcgAOiysukg/uuiAFbSbnO1U+WqcDsxb6pk94b7Wf7bYJh1PetTsNCZZF
9JVtLccMhCIFer5MfSu7LC3MbXZyuiNcvcHPwuXO5jVFfUNMJIw6tyC0wxvnPzbz
9O/tTxTqkwP9q+tMsKvustEQYvwGbmi7lLL0cW6ssfnPIhKtPV2b2S0hRu3nHHK4
imUDSwb5D8PCJI1Z84gYpZtoNC7BoDjNgNDJrMuys4uIfF+DAYealY9dcq9pNfkn
Accik3fnXc1m6gEmVxnOr5lDoaNnN4RS/vSUuTfkV0exiqCoTiyvb7Dvhi17A/Uu
PFAIgaamRPxUh9daKqjmoI2wtDb859xkLfYyK7k7TKQmTgQG18rZPMRlYdjmbr1n
3t9xyRTTq40Fewx2OrXH+xDdlTe5A4Z5lbCXYV3L2nJjXt9/2MYSSiApbtzcdmcW
RiyrJemcqr7DGoEjkfdQfmuGlTipjiPj9sTh0x7ylNpt3WFB9XbnR/9EalIN7dyt
WVKhIdbbfKT1rJkYg1VY6aAqK/njV589vfPaF6IqlY+sxlHb0/kq5pKdFaW7hKfH
qP4a1a8xjFuTaA5nNhYKKWBirGrGSxoiPL9eByf2OI4=
`protect END_PROTECTED
