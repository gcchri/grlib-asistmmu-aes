`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kLNcM+VZH8VkzPorAUHBXzP9Yn+rMyqJTrWWpiVqBuMb0C223O6ZzUEdd1MhmmW2
ebXCbQRnulbxXPbnvXVw9CuM2ymNHfxNJA7v65eRZLKewNnx1asjEUcMpMxUzbxG
DZd9z619IDWe1uEXoMGCY2Fw2uJXBOKSl108IEPc4KX2POOgBLwl/UWB+Rhbu2so
PFQXudCvEbWbDVbPHGYBk4w6qviSTOEjU/cujboBNM0FM/fxjT+pqupuEHZA/cQ4
pjiz7vgWRVecCIk5f/SkF7GiLCPL81WjH41c7VjYf2izdu6XV3LdCKQk32PJnv9j
TjXRRP7nOOmYgY2NWSTLFSd4Jacb6ZwE3uK1HS+t9bIc2RqhT+ou68KgU/IZXSuo
yQcw3s+JwkCMXdpTeP4biBv4DtF3Wrb7urXDuymD8pI6HNt1vpZpTCnq5XKH1Gbs
si+834l8oPaQu2cjZMCkaSX4f1z2oR9eg1XLbbKq9e0BhTS+N3BHnsIcvzEN83dj
xegHvQGW/pbA1cyA554foeQwCk/LGDSMgq9B8sUiybz2eCZCscBg77/4fZPClJs/
KAISuWTGkhbZM6GWiwXqoofv9ZaRDhhVjs3z9WfV7ugeESS0qn8hVVUsFzWbSCyA
n5BX3FSWfrZqEIQ+kxLGCodp0+3S24w5nwPZkj9PC/Ccc9i26i3oml+sMw+0Or16
XfYpxbH8LYlJSFNlK5WQLNQ4ASF93Kj/HGzzuxAfQ/OUGqdyM06q2hSRHQuJE0uu
7yxJouLNeneZiIU0ZlDJwqnhPFowNqYv87X1MTdz3CygLwd/r3k45gGKuZZiC6nj
izED5+6mOnYhr7EzByxyPQYUnNnQH1iOL8cQhrbK1wc+5067kQwthNjkHX2FnWUY
QcIZckBnQ3orKIj0ZNVToK04A6N4MUPh7VXOQS1OyZzyCsuPaju+DaoduA6fn1zT
OkUf8nCNHPtFffHwj+F8ZEbPysH2NpM35BILAcpx5vABw3iX1Um21afBhzBVgl1E
IZQa0+gSjNl6IwM3g8LcRy11qc88nkX7samCsSHbu2w1bs0GlHFLgEYSACEIov1c
Ykhre8S0DyG1qg2RkQbxir087ijEro7AAhV5yjS8hw07VQ9eOC/IJuNhpHROLxt7
Vkk7zmZA4aRntN0aoHve4z0n+hwe83LrgYBNwemesmSqeModWLtLJln1LLGJj2PP
ZkrNRJoI2uMGKPZd10YEcKKZtc2txxxyPn5Nr1cE+LR+XV4dZbrgKDl9hgvmSMOL
7ipK9tHFqtGvkMCdxNQrmqEw5RRveMU5ANE1HJbCYYuI+LRdSMUC33CruDLhH4fx
ns2WjPNPk+UNB/fGJc0UHdTJYmwfkEBVDflNBMddMORzgj7hFs/+w887t+NJ90Mk
J8Arjxx3pMLuEMfTjz7LfCeeKXcTrZj/xpTBtS4ycRYz9tIMlr6mVFqgsEzyxSxU
C45LkR0mPgnOnM/OrKovdK6rw3OQ1B7ywUM+d5XqW30+uMconOadCls6Kq3KmkQP
g8ZAXbTw2l26JjtJYPDsXgwv1AP7zLvtNINCZstvF/Dnu/Ouo7R2+k7mqtX1nK+w
uPzL1gEJy3dlOXzk8W9wrNfKAGtxR7GApVTCg03/6gPA9X/8QrK2eV/KIcezAUss
SViLVLobmcebDYf8NFjwqdEGmOWbWj9Of72l54DxM6FEcd1fVBJznoPfCBsRehaA
2UKqrel7bRJa1wIDfbzmTjfmVJoz2H9LBfMPzjY7zoaykYW/fPX65Sn5x5HSnpyz
F7LagdWYEnpRiog/5rv2vYv6VAjrqEb8DbxbhLT7U/SsD5ROldyuHL/vcGUTnR40
ta0JY3Sw92NSSejs32u6b/rgFrhoKXHZr6WX0Pdg5w9N6mS3t1Vhw3zeV+9h2K0t
t7R46Kz4gzWIaWVce9KRS/Z7I7j198uEX3K6hjYhg0o31nrEL64cNgpOU5fIZWZM
vrjGY60r3RTjOQ5eY9sA3/DwM5M1kCdhYzrMEMppdGcShmg+Y0ys4M4VJtWzd6x/
4G5hmC5ZrQw2KZiPeOs11ZVajsYc8aClQsoQmorKGgx790SmwqPBUodrGxpiiM37
vXeNy7fVsLOXt4+isAAMUCay27BarZ6CQt5gXQ90VxsjjctE7tN+6v1BTpqfdHao
ec4w9OBHT+LCU9fphZ33Ck3JdEPLev8JN/XnsONNqdQfcg6VNwPSGpJmf1Ndz4ly
itKEFCHccHkr38Ts6chVs6LciKmeHuAvUwqHNADg7RKbwCykdQfmA98K4lU/t1uQ
pvkOHwxoveiEX+Vw8m4AIUtT0AsuT4dBW2pzOnG94GbwqaH4TYOPalenKN1148do
sSyChfFj9NFi2qrWzevGkbM6s7ZdeQfTKeKh9+IqF5VK14f/uRhfU0HTDC56cJNW
wvrQ1h1hqq8TaghYj3A0NWwfMwqkxSB0C7nfCTG+8FMYSXx5bN+UPsPEj4+hGzDm
JmCrqkMmCaQ21DiN4r/eDn/9ZiU1mv3abY1dMLSinAZlYoH62rVmdgZvlWg9+dAs
HUQO6cr8ylkIUO5RtJM0c4MaInnLvHj2su5RPnIqVzDeb/rWlgWBRWmogVOPSnHL
AvN7FaBgDjZsdAyGM9E6aRKC3VmRBwoWsl8F48rAbTngrh3kpNwqRDazghk9xEuJ
wh9LysClHYv26fOtDLRxrA6YurteiLqtdZ2cFpdlpq5kKVtvZ+d6VAeUVMRQWGnr
fO6ERFwHCjnzBUS2lAbAMaAFRCogQ3T2iXwrEP1rn+5C1fntbAzw19PX5ja4aWZy
iDQEJBPvzZriEEEcmmNQBw==
`protect END_PROTECTED
