`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pl8h6DRWodmQLnZj55orgtML/3iN/3C3ET02g3qrN41VcOxSzoxKnsDUIy6CW2eL
gSFktB+wF6r1MUvbJydCOC0nlQAc4XhEzFlyqVOMqfvByB4jNzoSyehjgdQhNV+W
3wkkp977DqHIB+F7xj8rz1Vp6IJsjO1U1DxCqRmvbrREXLt2wbKChNY0a8gJKiGY
Ta2yB6IoPDcS9u3wyOHFbbf+zr4vXopuEEgwJMqgCsjSbjSK6WmTPqwtbca84KPO
n8CsKj0YhRyGAGGLHogTQ8ahlEguF+Yoc1EeLgQHujZELE/xSnPCSGIXsMTsGl0H
UC9mMwzW/5kgSpENirc05rDSWdElZh+/V0Div6Thhm7marqA7ffdiOlqNijaZPrp
frBy4dhs+ES4uZJRekVcsrp56oJifpghvu/ecldq7jrlALXn3mVSN1pHFLZYcS6J
MFCxKL/zCcnwpqJx9jM1iEdjzhon96ntD6S2F29H/ozC1cSqyUSjv5/YgLZh2FvW
3LcWvl8LIB+ebsqEIojfxZpD+qkFJxakkiyYH/Ok9+4jOnVxPFJEhzhPndSpQOC6
UVGiefl7K8cLUCH5RjuxQObIKskHocObvVCfDASaRQO94jk15VL5+DfvLynSctpp
vPF6+7uymRtlr3mJi5d10Fi9LjQkwKTUy487LCuV9SM=
`protect END_PROTECTED
