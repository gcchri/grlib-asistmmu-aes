`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P9gun7/R0DxwifMH//xrnDiwKjZcp8UXCT66J/88kiJykYma2oY1i+hPX3Re5JyF
LVLiv3RFlKhd12zR4p1GYwR6xLzKAWyQ7pNSBpyqJ5ExXIOjKHuECiGBjsDeD6K7
lf8QuhcH+tu5eEhdyrz2FLK9LEoB3AFV6h7AD7k2Fey77nM9E35iijanarsSvlXf
tGHXklIYd84K3JJjeDn/sNTT2Z2w+ri0Y1OBVgGW1YMjf5fB20DhwAzku6nLeD2i
Uhs13v1Pp4BLqtke/W1AIz5TPLlcfglk8h6XuG/WTio8FVFWu6zC0enHcFKwZmTi
x/HZiq6UXQpjfOAzPqEq7/6Cul2jDPYUAPqnnkf4WIwaAHXZ4X30oALpR5myqgO8
EZQAkwHnyrFtk7nf0q5nt9q8XCQs2bnlq9eakiVdy0Tu4KERlBvV7RVCfwjB2NKj
RXqDoAeiLn+ZJ70VB1zfzlEWA7RKNsO7qxwHyBW1Wiqcnqef7Pd3tSyK+SKaeuYm
`protect END_PROTECTED
