`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Xgu0X4uzfHs3lk+6oc6wPnCMzkINu5bPJ1GhOVSor8c5H+/xLbCXMBQVo/RIVUE
nI1oOsQ3MyYNcSScfPqEUfEaoNZHlL8RCqdEQ9W9IdVH3KJttPU86h3jxY8jbnQo
8AuWI5IIOR3G9cRntEAnzmyAePhqFrilSjVWJU9rn5dNP2QJ+lhy/FZ5+9ISA0pb
nAAoSgoifh3eb7/OKq6MUQechp2w9XZfoEqe+M0Dwk3W9UNSaJH9Y3Pm+vsM3EHP
dVIQBpEPJeVQa+7umFOdENOaL80vkhJPsajtND+FkvGQid6981knGjWeRKIaJOtz
lv8eAu+zS2iyplZpbDL1Nb1zpn5zWchd608wOgPQvEc6navUYu4KE7Jp/1u7Bp2V
jcxsG4riP1BAptQGggiwZ1TzjrrADF7FyOYcEhco97WZXzBXRVvo62wAoUjp4Yhp
qRoOxQttxErHQ3U3qpIs/tw0CSBAi4/ln47Aioo6xu0SejaTkoyVFjnytpsxNU+h
IgvBEA5Dl+t7PThlpK9cn6pb4jSTHtNGuT0JcW9sJO7QsJ/TLDqKdL3oLnJZF7R5
W5Ryvk6AKfWjd/TqsW2JosoWMoOKbjWh3qf2tPlhAEnNpfeBDGlc0dkGMWCpcbgb
zO7Ix7Ne0e5ZBdTYH37Hh88XV76PmkQfDYQ+9w31jnLMz46R3enIiTSqtM3HolnT
dbQayrSpRkkT8ZUc9AndypjMxk/AQSuy8c6r5t5vi2EFKWju3x564hiSYWvnm8wC
/Cl1lZkTXXnxhDMzWpKMpTNcai1BKyNttb4Vo9jc+1FQGGhUjYYc0+whHRhT1kYe
DrJgM/jMpIkwcSvDQ66H0A==
`protect END_PROTECTED
