`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4V+rJhsBlRSAxOBpsICojSqHGHJC1eG6QsZ3rRSnEyqyYG5tEoKoYXtIinpjUCGs
xm42OrneqGb1phTAv8EceydNcvjvibR4uljtp+rq8FYVRf0llvDmgxff6yxOXOZL
MY0yDHAgYQK+zcD1umpHvVEEAM1GP7sUKoF8hg2zJ9iLzFmOxxN4INjR7dBy7IT9
JGQ1tBHoJVdODhv+l4w6Dj4DWKjBq152RN1FOZyQz89CtOjjGyW8Ihl/L845OOic
eAEzGwYSsbXUhJiOg26FZQF2UqhqCx83Ylv2QBaotChHorXCExsfZdasmKYGZmIB
v1+1NjJzRrUKJqN5rOuRLuIxW+CiWZl6c33qBhdJUi0v2JDdvrQJ+mkW1tn0Cq+9
T3aY9rKczLW/DaW6A/Yybg1/jF1jd7t+CGdrSgNApaQBMMcoEq9E93Ucm3DttjNy
xuvkLBMT7x7xFP0lE01veXIWj8cphNTM8dLI0kjztGA=
`protect END_PROTECTED
