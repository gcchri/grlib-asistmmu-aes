`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3OQmSNnNZ7gkfiXwvb5rq+xcBlD56DJsz8vEVbOW8AGTo+eG2o2a2jWIQt7U+wjx
s06c7Me2ixqhIOyMBkeixqnYELo8hb+l0ICrZZQMTxksXJQmigT0W2VuMxeVIUv+
4EWyze4xr9i3FGgfsdRBiFNq6ZqEgymYoiO9hqE2cvjbYfLTIO64K8w1+O8QktRE
RXmVqShorOi9dHw+OU6G1u7YCaZ2ESObP7sJCs9XskADiVny4roNH0zcx8/l9cWT
3BnQhBMaPGSHn3DW91nLjg==
`protect END_PROTECTED
