`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fhxyYb6cnusZpkyAehCJhDPhxxWYYJcwhk1v8/KXxJWvzTIgRSg/UnXitcbPjwvA
ccZlluFG11lL7baaCxho9BlybIK+v/ojE2xBTuaXt0ABh5rGWFr5catewL4ZtRVy
R/adRY7KlS2El6plIjP92QvC4EODw02x5PM3xNI0ChkoGU60CMhpmBzDnciNzAN6
M6qXUhHfVGjp5G31w4Utw/Nk8JBTfiXabtwWaS70nFiRDxbwGcPTIl0VgvtHcbgk
L0N3hD2WadWXW14I8zlPHvDgrydwNnNxzvZXfiYv4AwzKNUsThmLgkOGK7KoL95x
bC+9lwp9ry9gdolvG+FUOgqZ1zzkRfQMw41f40m4Tj2pIqbQ0WeLOyrgH1Vsbswq
ep2OzXeKDS4B7uKuAdWdapnNX5TOGRE2IgKEYl9sRyb8kuBb5JcMD/ct/ZG0uf3R
`protect END_PROTECTED
