`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Y0hMlasQ8biZ0gDLdu5SSbJYlBlUTBdYdtr1FzOB9MDdaOVkxY2Ro7vgH3VpWg8
Ie3Uo0ERmcsbo6/iszUutjpC1sbOjo1ZyLbVLiw27kjxVEUcXmZ1VBQbFRo7JH4W
wrlNUMC4/6LrS1YORNP01wudxERi0P/cHvdfc7uSbHjoOzxmnMRn35HKLRyjRgRZ
GcWStuKQ2Oo5TysjGLuZgKwlnxRPgWPrxsjCKgIbUAi+JUd6xfBu0xc2GfcY4wJm
vVOU6Pu6mLwZVwXzSAhvC4QKgyiolcoOx8+oXlTXk/BaKthIOBDIk7/FxybVrRD5
cmMmnmfWnV2Wfa0W5x62wViaTytsv14jBq8GTDczssmAIcHSn5yQ44oJYEiB9jES
SyCH/DtjCP1EG90Xlel0wJnr+NNpqsGgN0w4zIi9T8YQ6eexZ6jHpLFBN7hRMbsf
`protect END_PROTECTED
