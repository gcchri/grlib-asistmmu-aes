`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
90Q+q9qjgrGJLYMcl6Kg2UOrG0wisY92435Qzro7cw91x2EHbFYzhto+HE6kmDRi
mBbod1FzUfg64bZtNcxDh9gzlbVzDcpp2l0Ky5/AQC6IG5pQ4ItDE+q77dcwXAPY
+0tvpug+SRql6+18HFjY4rMDrPNeH6pk4h6UY9TQ0KbzXx5FRMpsSn5/bEbgbQaF
5MtPK8TuWB+bdX1+BNwYDBl9xU/m22QYt5g2P1QOr+rjraRung9Lgy94aZY2uujK
gGCz628mTP0aRL+eQ+zsIVJc72nqTZpzhZ69F80rCZfb76/l7yVwUUN1nXZKXwHu
Tpe6CYsYSamWxJQrm3bNDaDhPHLqerGA91L/FjHIuKFGXWpMJjBDxAJmfNXOCcvr
UfqTWblFLywke2DgBe4NGFxKvf8MMTk9gXKlU6SXzhftkHvof2sbUm/g6Y0nA3sb
zM0gDVXWerQ70THPxhLUGy9za7b2vNW6Beu83VtPvkjVp/df98uBMpBo4+FJSIFN
KmZdlXilV04INDZqLaCAppp4zGYpQ88zmBEK7a3L2KibI1pNBoBIDonr9SKjFvsj
Leic9RbYZG7ndaKNXWbywzV3Wy7pDd4e0GdZ9nn9rtg=
`protect END_PROTECTED
