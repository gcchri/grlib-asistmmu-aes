`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
trN1NnBNpPaRBsWF/ehIapwq7WGtooYVPD9VAXi3tsJn9b2U7vE685DJty1h2VuQ
wKLsU5gA3HXFcGBZvP4dXsWBiTTfBenErUr7fPDP/9ZARmdX+vCVg12VtzwrRsTF
+KDutB/Hk4WQ8U6tQIW4yHfz6n0zkKZqLYh0aAZ5GH3ABIrU0nRlX/70aSg9AhbE
SWWESUtf7OBWRtSVnFVgbIA9oZ7papD00dF2ZMpj83MnGHsJzxywgHgLxKPJXVHW
RvwgCwvh2M/c1cUw6AeqQcNdpMWFclvcm5LyCqk2IbeX7Uq9ek9rwd5ERDE3Vb4u
soeLNIORHcrMTyAcowTZLQkqeY9mJ7k1jXTbsfAlTGZ6lKYrf92wT1aGEfwOx47o
GCS/MJqda/habPTpLeFELnlHjKZeg0gBhAvvZA19RzflLkoUCbjs4W3DZ21nLvpp
7nQ7O87CZOvbNJMnwt4GU9umFcim/Noc+PKOYHdRJr4=
`protect END_PROTECTED
