`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqCA3HwI7snKPrV96rH11J9jbDKCXYtNNNxvUVBc6O4Rv2GcvHuKvRJ/XbQULxPm
IuDh9aHWlrtQFTh+1/pixBtDw6zdHhIvzEvntK23aCREmmNnqf37b2Wjf4emAaKb
7q09MlkhePa/HgNtJMwRijf4heqR3b30h876haVE+ZnrhW1zKrBHeofcyd4bT+vH
sabAMrPEh4oVlM3tvZvAMzR/oDHU+zA0LFmSQM0EV8nOsXV74/oAdmSAbscT5Tza
d3ujF9YQzza7h8tv2rxCaab5/LhLo45jJpFGF4fw0FcjmK4+l/10qpT1wJHndU6i
Dvg5Xv7H0SRYfKOH6uAA00LYwRZw+7HzxfP/RF3Mq0CD8rMR6KuXpFY+Tmy3adO4
26qtvRxcFfV+HAPTlF8oVe1g+1N8y4j70alEsNqYoIseNLrBDahFCqr2cngnN24x
EJ1rbEWwgUy2yy7Icob72Q1KsifyJHQ6ByuCY0h4IV4kiIldPS+e+MBxOx9WwLYV
DIMNeTmpQclu1MWx0lCp0j/94JcY6JYtYgKqm6pJrN/GrCu2mT1Qhaw+I9rBjT4D
nh/e7X+VZi2Fso7gF9omt6DhFUqIy3T4boVvb+xT6+3RUhi1RPOADeZ8vmiw+oNL
h9al0zA6fwOi/uGtlOEnl5NoGqUon3VRKaLZzPJjTYVEYVXi0QlTj4Q91fZ8UmrM
fpQFLoMfoIKm/op5gPuC7YiVN4xxCsztX6HH88ekxw+hSurC5KqFlxJ8aafEtZFA
OXMKjiLWQ7bESN6gOyDDBXDFUAIF1ePFYYbobod9FiOln+JVqkdUjy5b+c6q5mK1
+OUj9Kpi/eqnHMe8b7T70HmleCKVb063UhQgmDsB0Z1JLxqMvrnxYk6TYESMu/D/
oPkorVLKElhqQzaPotVkVskfRkMvBe5Szno2oO3Opsqwjci1gbcZSgFyRekF43l3
e/5O0MSTrOyTkH/TJaxAOnkwte4LLi5PNk6uOdwBXZAFje7Bu7Ky2fUc6yW8/7BR
tpdRldd77ku9Jx+jtu2iffjTbdhppK6PWW9Dq1Kn1Ww0OnrlSjrvf7druCXrgLn4
b+Ve2AvS7TbXUg7gooKpLQHOwI2YwI+o6F2XIRjOt7EsK35l45Zokd7/e+wEGGXv
1CRO4MsLjr04njXPrvbzkH63TJVtjum8nWLd6L1ubcAyfe8mzn/2wLMH8EXKHDlQ
QGyQ+TP/dkL+kaZt0WQGfkPKlYYgVjw3p8Bwni8It11AdeP0Pn0BfEO5RTyCgOen
s6aNrqd3Z6vVsT7MdFTZ3ONVXLkRroYOGGPXqUrq7muKbp0mERhPy9+KLxMOxSVV
Oq++gD8Vap6u7yUKuB8LlTReLpTD3pb7+PU1ZMU/r7lfa1eGNEItk/KxeWqdWzVn
3zdBVWQhp95qpKeQMUGpfBBqoge6vU7A5MeZp/NzwbY/4XsaD9aqzmRK1+nJ62HL
eYDNEX4ProBei6tXcIu1l4fkmY8NJuKODZ8u5rTgRdqE4AGBNvvv3FxyVp6d3Nzp
Joq2+RVQNiz/RaIV+7OYDRzFjGUx+lSshzby+hlMIbJ0Fljg8u5NRFUwua6FrJUT
6vfcNNiUw0AxSEmzl/VnhjGtGxID1ENHm1Wjnp5YGTykAgmiQmKTplZw3qbVl7de
Gb56WXKmDznU6BYonLksBFizVPLnO3KZHfRShfNI5ma+UfEVC57mSuae/tvgg9Gu
BHoXANfylZHMbWSNr3a8xga0zCeXVfFDDDl2ys3/bCVCNWaBYzv/7mFsGeJsLlgl
oGYPM0tVQRhQnMrUDHD6QiFcXXBtOF2eCHEZH+yJ+q4eZcf183m56CZyTmHQk4JJ
`protect END_PROTECTED
