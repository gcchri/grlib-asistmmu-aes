`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zP8xj3DQ5rRWOBf/D67Zj3LcFIv8tuDNSkhPAFIdXptXcO8h2k5rKZapHa7/UHTH
dS6GvNEybT2Z9D/lrkorWmHQ8I+bT74OLRICFKRYycC+4BY2rxGzRYQUhJNmSmDx
S8ZdmzDLufVVQ5Q+7ey/P7GcjNBtomS0E0fSWQlEz+yoVXA2sYwWpT+qSkFlZXrl
ILb3TRKkuChnHxXaXLwEMnnBapkC0gJNR1xuY2BMueeZJgPxqdIormMb/Ki9bAPN
29GHJBBNmBluNTtUuaMaw+WuWBZFs4Rx3h29J5xXaNOcy2125uVX9b7hjHgkJz4M
HLvD5SSyKN4z7f2RBQuVMEf1+UulRyz+K7QoQ/oktXda5+bwakESmoAl8W6IagPw
sV+uNc5UTl9rKVXKLgLKiEvmRrqfaA74zcsRF2cdWa1Eym8+zDSbdypBtmBQSe7t
un7732ktLj4sIT052+XZ8F57KVSwLKx7+a5Sb9kvQhKIajZFRm8ToAdKB3+bWrc+
XLPy1UDnVQmlXses8SvWN8JnvINAOlaKrKNV9N/vaoNVSsBawI14SwG57WZTXS9O
v2nacrUcJCqxnpr8J03nlliRzFnnRSfJSxh0hkdI+eNMyBXZZcE19fcPkHoaM7+M
mO303nxE73afpahPM+eSU0EfgdpRe3+0i444Q9AXJwea9b+Hv3Up9Q6Db6CuEadD
B2jaQik9GUb5bLCVuTEXBivwKH9XwVs7gJvLVlhPyJY1VB2z2qSNKGc1Sw/5AdJu
fhk+PhJVqyhm7i/9M7FNMX1RQdPY1WU3f9MjImAJ2h+OJpKDLVzSmQ/Awfyx/BVu
6fNxmuaQdZRlgQRS3qDRxeOjU5APpvHO9ZP+OTyAGBAb/ZxSQ0VM+DjVvZ6o60ue
TXmTSjWjkMPICME+xZZ1WdLhundVi7i8WIpUyNcl09kmiegV/+XJECaid9VwQcnf
DZLnmYGZ9oeexqlHq2Y4FprJAk67ZVfxjMwROB+GKClOYf6pLPMYGLrbTbKrsAEF
nnY9Nf6XXGo0xwW/SNq7zVdoQcvwHz+qnxW9WidDeSecNtslG/Kkn4xshrWutt+t
bkaLRgA/x3CH6F7T5rzRWJmCTrfabithhYoHb7OGykgENO06dMtqt/HPBqb021XP
wj4v/EUZ6QKygXKbfdZRi8SlF3Di4uOenApZv5W0QUqutgxhOC0DUtWrOliZHW38
PTCw1ZXHuPUdmdV4jOCiLzVZNPNylKsJ2ZdkivINeMG84afXBD0CETtCa8Sb6dm7
aPFFBbDLAi7Oa5EPti7827yH4r038+ty5lMhFoK943LEhJW/1LHq1F004FVFMFBs
hlVCE7oKx04msDdQdz4mU0xcX2gmpORZ6xesYVGPfjhcl/YPBvyHarZJ3z2Wk1kW
3QZEacTjLC+ZoMAX634BkRbLa9xkz3ZmwaewqdYL6yCs9q4zuuQ5Ba0gz4zbPzn6
dAl/WZ1uIekdcXcTwOghCsbTNdDCvrxX8JZknsNNULaKL0Qtner3IJOr71YzZILM
2gTY5SwbXbuNcxQ9D/r9TgPGlmGFOaEgKEJlV2BKB48/DymArFB7uBn3RkMxEk7E
s/kqc2O1pCxGhBQ6wrhjVX6bJeVBBQbqXt4YvlgJrale4i/fLoz/r8uNEMmwXc7w
VyqR5oXmipPNgUNIV/m897sZSPK/rtAAHUSsIINPS9vIuYn/gQxwLvBgrvvssAm6
O8ApFPjNhthIpp0Lpk1zT9C10HXMS/Uietz/kulOk1gk09cKZ6z63LfFu5G1HZeh
5FJB7Q9KRCYcy9q4VPok/TYQSn4BWkt1+FxA8IJdN2UdSrOT8iznfIIKJqa5dEay
7QIrkrdqNEdDw+X4bGrsvviXtjIgT/r/BEZvXsQvcpKvj8S38vDH8O5l5PQ5Xz7l
9EwOrIwmRU5l5msJ0qvfWU+W8w6lSNw4qRf3rfRpbFpKpjTpBa9ZKQCOGBjerlbH
69DYqSYlq7b9hfh+i13zMlgs6+ri5Y4DUVLOO8cQGAWZ753A2dr/Kk5UolvBsVzm
KC+1Cf2YdOKvxnm4MPQrB2LHb/oT/F/CYT1JeIacYsnIJbstr2c6dt/imo7MVlCZ
EGJeLZtSDvOapOrYKdkr9J+3A5470CZmH1kj3iwvyXRvh7bu2DAY8OZC8/1rIlVl
l1+frRsNs9hRGlejNjKbwbtaGysztuZkx72mVRvi/TcGukD02Yl+f0aap8RONFch
T4VjbmR4uZ+GfLNCRUQYC+/KhooyqBmUwecOaM0yR7QEn4LmSd6rxBj8lIxksMwb
LgpYPnPTY3jNcmR/UJEwMu6UpCrOqDk2WYpbvKLePGYGx7CBoJHQ7sI1ypBtSQ2e
Ntev4E5ijIvryS1P7iOmfhAkfhlMuXzlprTzIrsGFJvbfHpEM6VQCGdwmsxEG5gf
M47bfOsYErVX0js0lemS8v+/p7I0R16PmDrw9L9GLujGQDv48Q+7fXj6EtU3ROsl
0EL5BOFJWltkpowWa6f27/cM9QdcfbvSCUz/mVx1VnntMoaOf3+8gQMOpMlAoObe
Xkb+HkLwwgzIXkmXR9brgErWY45UJUgj8n54B2G3l7wKyMwc5cxQjx0/6/CW6sSX
DGvKH7w7vqo9ytJYQBFbAoekiF/kUn6Mxp5GXKMLipRkBlSEdGgwhZEfNnWyzwXK
or8wegsk5diovt7JItcbuQ==
`protect END_PROTECTED
