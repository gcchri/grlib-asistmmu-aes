`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmhUDdUl+xRkcmH4X9Q6p2hl+ZfWGwmBRa1Hcel42omJDClOFHhu2NY9wBtyReZV
GMwqf0FXJbJJw3Sc2WtZcQwR5dW3Tj6Um5EGt47g7U9nvfN1rhJt6+Y/Z6h5Ix/f
cM4rw0GJHHO/KZG0UEt8k0Bgw5c/7t82THQuVNRvLpUWECu4xNoBT1X7ECixw6mE
8wZyaRh2UaIjeze/p2/KSsg6n5gvuo3UmvxkVZMbC2NcpyN/xj+7NfDTDFI3MsB/
BChR4HE5Y1VKo3/QYiM84/7Zu5Wag8ndzPAyyqwvbWaw1ir4vUSlk7dBh6EzEdjp
F1oep/fYYBdO6w7e5msVaqyu/WweamOpPgCYUesYt5w0KrLW3YI6+2pNGvT29UuG
KEraUtXjr7OIxrvYitKCTqiH8XfJs5CSfAOs3FTcs/hkT5kFpm4XmFrekS46uvDG
sJj3HYahwDg9Xqz4JezRjVVOmp7lbcWJB/f+2FK6LeKW/UHu1MhjABIlaOuflAKk
hT0t4fVPacRRY8Ya/9hqg67hwDv9uCSm/qp92LXoF0kwsHWwb8uJrwnA13j9LDaF
yzVuLfeeXV122SGGnHGKfDfp0M+YDG2T6vJglFvG4ZITlHKlexBYBPVQ2kEavsJP
sa+PvhbOSxyDN/VDyA1o1vC3/YK4x85pb1/F2opBrEkC6oCI7PJILytLLPorUGfN
b5t79TEiKvqy7mLPzG/Z3u+Ko1qCQjJUuzunKE1ZtssVJavxg4rElP9ud9LoD7Th
uDADEo+qiTS8UqytCfp8kITaePLSj6nl70Afwms4L2MrXj9R4nzaISXw2jfqOosp
IOLyhHTiJugrSKZIKmpJrTCC/mKDHaTYzHZbsGe//pv5OVTW/1mU3sAImjX+00mo
rJ8qLd4ALgNlzwxMvPs00ETeYyu9ab/xgWfRFnfV1Fuv+Qj03fHHoErFPKeMQgx+
K2VBM2Ek+7eGZGBU25FJ7s7rCSLtdiT7UiCs4lSFcAupms2gTRjZrYR1WFdM5SfR
0T3w41494ohLJZthwMSfhfW2q0MN3aJhQtjwzoJdL+COUFj1iXTU7XH1Y+fAXYmI
sB/N73I4b4gPpKCnEm4TC4D3pHHZ85arXSdu6b/c9VPAQmn5gnEtPOC9m+lTW5vF
MdR5xbRMrsa5spr4/LIr7ariuNtw6NbjK/XsS/dYWg2JXwRU0Ortdh8UR7NphCIb
7Pmb+QfkNA/0wDGEjxNjayoVpRDn4m1MGidMRTNEbOY5s9Xq6Jta+CLf/DpqwN+3
`protect END_PROTECTED
