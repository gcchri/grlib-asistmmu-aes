`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jAx2l+ZqmhT+6hINo8U8QA6ljDI7tVQwYpWiTcMy+suLHqBDfwtyJbEeKqdCO5Xe
NCaNDjDnMiHwjTFOxvTfiuikr2v5McqSJXCQfJcITjkc75EJxo/Tb1QFWXjxgeoc
0yHxfzH7CnVs6pODZmcVMBooFzw0xWiNZcoZNa3z8qZZJrXyp2QrJ759H6LThPcq
QCFBobp3OgDVgyYoARzEdG54Rdbf2fSer/01GWq93JunZ+CaDnmRGyALswRzacvQ
jVrMPI97DDK4KORk0EzuBw==
`protect END_PROTECTED
