`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHfVkqjUBwKpFPAtWgLL4KaVHzAAxiYnFMhlUE4gmxYZDZEWxM9WDc1pUT6r/Da9
uyBc5zqds5fhoPcBp3lQBDReKY7Wja+5NlF99KMF9Jfsgfg1KMDePxRM+T8pVjdT
E39Hqlp4eNK/XMXSHeO1Ngu2umFULQnUwApq7dIwRaw9lC1H+T8639mDpQAUr9YR
c2tbiRTvhMn0AYcmH6xrVxlcQYdOGy/eGoV/4lfsRauP398IZr4bDy/T4fw5zUkd
tGq6w38OVsukIldORjhMGmdmD52tUbAuvQ9v+0D9H2lxVajxt0AIHMYl7nsd/D6k
ugfUh3ZIBPxE2gSKqaksAg==
`protect END_PROTECTED
