`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JzJIqydZI46GDM/qPvsr7g/oPmqJLn9cy4ff/aNSgpPYT/IIsZ7ks3S8x80meED
Jre820bxCiuOZJ9c5Pu7UEYQpxE34ks9iOvjj52+qEqLjELf/wkChdf/jnNsx8Q3
dG1FIKUx/yb6bsa3DAEgR3InT40xDNYejJ+HepP0Gh765ecegoIosZ+0KXTn8pZd
y5fwINo/BJDhxgRXSnd5BoxL2OSgsgtqlzxzfDflNAtaOqEmIKGe8EHDv/KarFOz
tstPuYbQT0dyIyTZ4G045iYPp/7coleIinNiuVvH/g1hnTjXRDVvh02uwKbkfJfS
6+HTuyMpJBOljgqZr+hcNC5dPpuNqgMRHwMCgjpg9nQrVYSERWeTsGH1/il0bI66
e0cUT63FII5m/jcQro2Yccm4chmYT+0fhJiOOtaxrZrWJ2LmepqWCdy3KIKrL+1W
3280wbnB+m7VSkLkKLabfEIrb1gnRYP1nx4uEbZZ7fPLM3jZEtn59GyAMrb92da3
xcUeMaQB+A3xm1IFYhw687lnzQwNrt7zC9QQ6HTDglKIahdCNGMDfx0uGIIKyWRc
+W/keeIxnPXhjvVCIJxrAJRuXxmxOEZfSq+zOTjPNCAWRJ0wt3vaWvypaezeYmT0
hwpCPwqg3R2o5zrp8Bz6OywByROl351P19Tn2IgaEiqiMIpiO+OCIJlECoZK6eGQ
ii3L3qp9FoEAJ1i1fyYw3kvVfdVWRf1FKZiT3vduViv5IIiF1uBuwhpUQfjLgmQu
NrnsoJLHkJL/J1gE+oUtRmBJU3LtXFtm1W7TU3cSeSh/NH94tZZil4AUTlBGzQjR
CpxlxC19aQFyvu2FLmCTRh1rRo3kNQEgk3YNXsJVj/xNZVJD8NG6zCkbEnkXdKDQ
yg0JhN6Q8MrJSLkrjuV6PT7bg5Lkbg8B/3ko0t57z5KyhUmt/FPe3JxQWpRa9mtG
NxLcjVlMIO4KcEanZSWQQWu6aa3KKPSvMmph9eIZH9grWjJ+tYAGoCmi7N8qIViO
TRnZKnHAmuR0cMCcEnVixxelSKLeJuGbJd/IuNfdAPCs3o3cK+z38NAQG1qbZN5u
oRzEkt24lTNx5M6dRiAmo9KyfJEvWnVRZeN9KipRYDS+mU9wuHJKprBStKaQRdAD
I4Km0SBIN6HjMlcgQ8iVmPK/BkNGpmAk9hm8X8A/7Ali7w+YL6Ed8F3MvPw41TBw
GFPJibcmOhIdqa9LmIvglcokM4hTLKz3r4VA26SjPTpmC/wMUpc0ur+6IsFqPutF
`protect END_PROTECTED
