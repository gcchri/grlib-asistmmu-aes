`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKO7g1evZhqtERe6SOsiYwm64cr9uEZfp4YNuprZbD1xdEcH/1NrWkGScfNAU9ME
Fo1VdW9OxvllX8mKfO/dSTzNSUFvr7WDIvayOjaCwM90lLFMjO2NDpFKxOOLufET
kFEdEwvAaY/+wxML23c/yCUm1iDp8YzFgl35PudwsjE/khWEmqK08S7D3HrVmzD7
SJG3HfFqnDFVzRGcmPmeQiVQBdnnTw+itKN8h1EueU0IGOBCPZiQxXPEBKxvpTy7
nNFmEcDV74yqrM+C/r7Pa2/bA0JPxpa0/KlMpZO8xKM9DbiKQ1l+sjm+4ofdYPE3
tDOcMnYyzVOM59deX9orEF7Y5QHPRVMS9dIKoFHzBi0SJdM9rudLgi1oT9IuHSJN
e6LBSWdLTXQdpS5LJG/l449b7QJXPzY3AhZDEHgg8wRvkq6/cHhwVc7/C5t32VvL
mAopbimgk6rkJv5hDLwrfAtdon80C14s2+L3eO1G6nlsNCLtS26Xg1LbdMlLGbxr
IfMmj4UNUw8F3JaupwLcj+1MV1bmZyS74dglnBihKYz1e1FhzZbcckqmAMZiBPMe
8JbCeRZk2LO/ST4qvREtAQL8MQirSwYSAapB7U+bFy5mvDHRj2TVmut92T4CUMMt
CwDU6Lheue4rOF+wsUEbzjJFjC5QhwYYfC9lJ8FQfpVu9CAjJcjmzbkZR2YZCiWI
To14QfN2oyizNJeMuLmewPfeb2Qn87n2+9CMRRfFf54iwDdb+8JunzP1F84Wfjtm
nozoPdoixei8tml4LqjfFBjHU8HmUjoamP67bzxsFR6BR3psmnWnxc7JPa7VC3RP
jmlBulVOZYEPHhwVviHSxTfzD24lczkHh6WvDG7CVTlfEtAbn21rfka/8RKJCR8h
SAw2ZdS1OGKWxVsjW9m8/iFmMp9W/eBpHuKT/8jxcabO7ihSUlx+SAM3lCNM+gOI
Vzdx86OfFaoy0yzRtZ3kpopf1FOsFybd5yJXbFEoNYpMLCrnim6TOrdXSepdzWLH
`protect END_PROTECTED
