`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlNWQurEsBHqVos/dMXyH+V8deaj0QB1yE1q/Tysg+DdNGIFYalQSdpOGGV3nxQX
NtccYKyS+Y1V1UqSCwN6EVddH3rhGhZm/EcKoorMRA2Cdcno6Wfq+5hPEDK8olCL
b0SqeYXf/sCqUbt+7tA+JtefzsrrP9x9lgl1BKUMy/+/Kf62NZe7U5hJ7MoNg6uj
cimugqcNiZHht933cN6lJSSEgVLXDFKD1MwZv+6TF9ciCKJPyTeQ8eTXuQq+8UfU
gIRbXsSk5c2L2iL4331Z8ZlFgq9QYifDmAouQy3v6RQlLJFsCNTzTTLXJv5o8BE0
cus/1k+I3r1Z9nS3/PtNAWIOGvIYFHsOJq9VIMcYitj1DbL3apAWxb8C2PkG1xDf
Bj5LoyP2uKf5BZ14kvKmFyR4OzSwmo6tEXC6oIPMdSu2MHstVh/wJ01p+JMV7Mf4
DCp9TEx2fchz3zEDFrLkHvV3vkmzQkCQVgMMCmMdvR/I4sMmvBd3qXsoFtutiMfr
`protect END_PROTECTED
