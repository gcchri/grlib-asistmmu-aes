`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mTEYljkr2LElVNmdmRSonu9hCKXULMlUK3XffreAG0WjzCOECWdxHfPOsD1EIcAE
H4d0i4mzvEyTQUCxBZI3s/p0SWowKIFCN3yvzfrlUJ9VMxLclSL8si/p7q5WNTL4
ZgYoLfJ0Ee/+fpfZSRFw4WEDJS708KHlN4yowuswUBhn8hFCBj2OkcKKkuOqCKvd
jHos9zm+m+dmxO03Mw/eml4Wn3vCI195btfs3J0PWsd6/7ZqOXGf096iFQgHTLq6
gJvBd1olD+iTIULhZpYy5+ggxMO9Pc6CWfTmxqEG8KBHbclafS3n1B3hZvE/M6zx
AMlJPjvk2/fj78w8pk3ELXMxq/M8UdFi0ZFf3EP8vWUuN/i1leesX3FcLCnr9SCF
x3t3qXTovEBSDh1rClrYFhVA0tv0FcGf0xS4E7ONvhGIGOuMenT4sbUzQ5h3Cb7g
zNYflCbKStrpSXcZ4CQntzz1HCKPd+VXtsspynI39qBI84XjDVZtKGSNMvVVaSAO
0oyqO2v2/5U/ujYfigRHwtQt6k3bcMr/Q4ArWaIQ8NWNV0LYJuo7eQOzI6RamXnR
aNPNC+BiJdSPCoUeA6fRqwZ6m/ETIzCaGTFxGtH6K6LVXX12oDSj08+3W2vLmHoy
`protect END_PROTECTED
