`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ma/VQBJEsPshAiFDNVgF+UQHa011ssF09BjgZzXJ/kMAPWI4+FHu7WCOcA2Hs5Sx
lqiCvAmfp2anwlG7fjraA4fQek9f3eoN6Ih8XubVTCPkuN5OHVOR7rad5FBjOPiD
Z5LstsWysi2IFI/mLdBStkS5JznFkMtDPhG65mv5rQjGbryp+IweXtV3a+HggsfY
IX64YCHJUbF0zH0C0BNhgLxPgbgDQbqLsV1HIGCR/EQQ/QyW9CuRLMUtSl6iD5CD
Gkn+eI5ZhTcNoE4NApbMLc2fvfV63D5kRkJ3yHnwLr1XAiUM4uoroln8pWXUpu9v
mzpjkikHlra8HDCRGf0+tKacxF+K9vDtDZZArdzlTTpvrLDl7ep/EaYFvq15rKY2
5rWgKGok79zC9mw40sQlhEfnqLXud0UHAn4rDhFakNFu2q9FdtbJBVnIu8R4jv9+
`protect END_PROTECTED
