`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+eryuScgZV6e/VCxs2Wz9NPiB2wLuyDav9G7xrZPpXGCL4fq712sljAhMd3q2gMC
C5weqUvanjDpG4hOlr8+DM01XxVrHDVyM09aVWkcPlC3oIrjwx5mWMbKr5WKgb3z
nO6inkc5HJr9a1DIhEdVY3oNbRbfDtVr7xTBDKvePDLfAU5V57mMxBEKAaKtisou
/3Jq0uG187dw8mygd8mL2DUfYpnrGjgmgnp7cVjP8RdW8Hvw8tbIXZmMKVDWMSi/
/2/mJSzNq8hXZZMdcb9Am6y1yrk4wQdr89s/G1yAR6DbC3SyOGjinl2rtX1vCAiQ
KerjhNb0mEkqZKEV2lG+uw==
`protect END_PROTECTED
