`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
22Qz+wRmxj2cBvAIt/7CwIZdMqcSfI7RQ7aNfp9ZEFAbTiJ+divxS5+PWQcVprvp
mFowGKfZ8WDTtyKHPcBubMDnsmcOOi1xmJWxuOklVJ7yy6RfxHXVJmlHQuk0Mhy/
+QI0QsoRG/+64fX2cT4X+pVs/ijaTlpF6VgeUEywxakVGSjSLfFmfqftf9Oa7hAI
S0kPlb71rqgx5T62HhAJHBFDO4y+BxoAXzqLdm6gjG+vne+ePURVlTiZ+5ev7FwA
IM69FLht+yt81zd68dIgvXsC3MPPTqYnJp9SAoOQPQYaxjpCi0/dWR+OsVfn4WIW
QxWUGg/7pSH+fDrHUfX2u3vqc1bLOI7ISXbPsziL0pclaNOJgqojvcxLEmMv8R2u
Xm2Hjgx9XxikBwKlJFEscYyzWVCs12/EsYNUdz2T1J/0NtDu2G7Eeh5EtyvlSvak
uNhCEuVDfJt6LXgKS98bEo3nPyUdp/SYxdSvyG8TfJWltkM3PlnMMJa2Uxikv11F
QTQkWdN01admVWe3ILPZN8jHflTuKl4ZmYn9QuRJQXR86tZElo1l2+wbZKvM0Irb
0R0Jvy3KBLMohvVQn6yEI0Y8EqtdW68GraSepnKR99s=
`protect END_PROTECTED
