`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v8qmwahnBZJjNyqagybcOXrVcpB9qTgM89BHXFa5zJujgyGPnf/aaWDLKyr/NsMQ
3/ekW5O8XY0xlV7OcK3/xt79J8mnyKWs7TO2Fs6Cj4P0UJ1s9JggjxMfyoZqFexf
CT+tUkz2XK//NzsbFh9iWCOgfF+wEUIBg5YxXdNYF+BfUqyqE1+OCB4ScQR6D+wk
nl/m5HjuV4ZvoOibiP1X5+0kGS443qPXmZBZY6nsg3ueapQivdzh+vIyn6PMs+vL
GIhtEs80WUrJOvr3XFjmqicyz3G0bwypKCjkqDYzgw4k9w+8g/ErPvPntpwNdAdv
PiArdCRACiKsvXFWrARlKWmP/1D6fTIpqH+M2h7yFkzqufUQ3Jdp9ag8/s/kvE+K
OuANOkI3Byfq+IRUC4AIoxC07Hk66gUo1m7U4QBbuuCV/zxGIm5qX3/xcEMEzTA0
AWxzCG2vV9lNGYC3zQruhwBg+B88WwkXzeVR7p+ojjY0Rd8cAox2nMDDtOpRkARq
iOOUIOchWn+2Y7pm8KbCPxcH+ss6r8ZNeCSMlgVn2gfaTKEUQny+wvTZxpPyy7Lh
jbzoAmF3zYq3Kfb4EzUprpKZacWEnsklT758zxfvnfsbE/tQgm3nujgcjvcOB4r5
NP7ZgiGxUbUWfGFsqdfbDYNlRnqMN/vaDoSVjPQz5ro=
`protect END_PROTECTED
