`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6dU35jyXFiP6ol1+sgfabQfUe5ogqas0ZwFdj8YboGKMsI46J6GdD61D2LEEWtV
K99+T7phu7icwhdO6RgMCbFeFuqJBilmDy4udo25Sh1hFLwgk7JBVmTzUYsRVphp
JFIZUTc1a77WYIb3vzbeNZ0xTjyvXPZ8Xl6IFNEm3kr/qgCN9w1BC5NelN2hJVL2
wda11Grs/bR0F+bbzchn1mJji3JWocsczbVBDM6BElu0oDha9GAoUprUAGi9jWMA
5u4caVH9t4OtE7h4MnfDNwi/sx+nrblXe16DJ0XLbOFgEkUMJ0aeegBOYveptga+
1g9+ojUd0MvqNaiaz+dNLD0OOgfDSMv+QMF3A/vq/ZN11OzbLmn6v+Q9a8m5bmq0
ZlSqGGcqYwCWg0Nihvmhwrz+8SLW1cm2NbppFLCgb2dB2FhF5vLY9ks6WnwSXAdd
9u8DkbfHw7ucHWsjQObn981HuIMJYPC7rT53gyWS4P2fEyKlyISVRZZgdz+Hikn+
FE/Cz74VW+czM9zOjMveUgDN0ewgDJ1RAXeRL6dxUZ8RkpKGJzD+rInqHwA2iB9T
zIsZMJ+QVCmmWpgL1EqquIoG8ZIzjcxP9EJOFIhdV3nN3FHwLlLcQsdrVtJxCPIu
KwAnTs61Olo1rkMOBbmBVQL0krgxDqFsu6We3uTLl8Suyl7b4bpvvWXDEshyT6xE
Y+a/WzUVZw1y9zqcVOKR1Sm2OPkcmil34z3qtVtJrkzZaMAXi2i9aOliahUHIMyG
rbnYV7eUzcnUxloOBONQRBUm4yyq06Ycr+mE+MKYdNb6IqWnu2oZYHZ5fGNde4mH
4mWPSq63nmbA6bl7QyGmXRDa8bPiYbADPWySreGN07YyQswibPl42cdQ1BM8CMec
r1BWywsMHuAoteBzEH3l3u9MHitW49aEX2HVWmRNohL3kUmwVRhGQkwrRjY69XGS
eqGNZqYBy/6VFppU55btI5FUE/Ie0doOoZeYIcxtgI8tZ59wmwgMph4HApyMOhOh
fv/fRrpBo7hFUXq0aPel8/mTKG1/sGG55D5+CMQkB2UiWh6iYD1VF6cZVpzbQfWD
KjV3nf9/9fyqJX8Pvg5GFLWTFEEBB5RPbKKpgzN+jRPYi0AsU5LTKQvcSsbt0lk3
5mzlThrQn8fcmETClkWyEdrTAtpAWBePF+ZPVkNHF2E6dSVU/q7Bj5WWR5VuKiEQ
XutW6PP20Qp1hMtXwzFgYZ6Yv4imn8UGH6v0audjHSEOyDa6TzchBQSdqxmGmZ9B
wgdFNC7aFxHT+ZCdmZ7p4RvUH5TNi6cE4DWR402Y8S2HkV6K55St3PnEAMdBJCDo
v6xVcw/XO5kFtrd/NTg1Kf7a3bOPDhgWEhbybY/VFVZQ1gNobD2H4vEGCoOEqaMM
xx2+pH3FGZzbMdOX33TvqRzwcwL48DpRUv7AmzbhPOAd9/f+N+fEIXt8uxcOkQnd
MQyK+fd3NQ5DkVBAesIIHzK5tgioyuYRe1Ar82ngyJsT0GL0KCClN4/RKQ77Vlnv
1XotF5tMHDubdYXQWKsoRPii1N69LrrDZ2AC1HXnMZitEwTdiv7eLbaDLs3uqEgL
VlNaI+c7VfOWytxs4ZB7vsFhHN6SXTx0I8kwo64ZNeU5EPEyiuON2MqXOmrELD95
1ZNqorfbS4n//jElFDPFxNMTNUg6w0KxrAusd3zDnCSBGiL3YWSReE2+Fb6WcRrP
bcav2ysL2sZV7dN4qHI5dg7Pn0xKIj66P7pmEU0E4vaf/O12B728mIj1ITLfpsV2
mjRg8qESxamkswmQwyCw8pGkodVGjHjaVVx0SskWjoXzqY9ZmS8TPZ5kmZ/WCV2X
JLplvwfbAhPYRhyLiib15u1NnhL9D+MK/qix2sLyGW1u3yzml5jAYx/7w+TDjLr1
QCdnxlSVAH3Dm7+5PBBaYoMGpsmWKPYw9FB8dAp9LxQK6ARYx4I9RpmNyujVdiX9
aLU8gOYap7vJFhtErvx4oZBZ/R6bG6YaLZRwdwUDjm9Q8DtqNbw7RJzy++9nuTl/
65VkRqlct4EHrzceNlnEUWcVfp24OU4aoAVHtr1ol8BeLQFrFhO5J1yzlnC+ejHQ
5690x0ejxXzhDqdoq06aNvHOZIBa28l3xF+x535J9SZVT04Hf55sKaTzz+tofIe+
HLlAwZxVyg0gTiJEVbVUKlStAfHsHgrFKh+jra4n7rS4Z/FPpybsiyOe17HhaOGA
TK9fi31u2RxcaybpQIvzrEyt4cEx8TUMFouxfcI86S4eEXdQRznJIr74DTXgMQ8x
87MHpof/dtHaJsVzKrkEuHF+tMmldb+xcmNHqRI/bt2WXBPQE+oGW8xmv0eaEyMZ
PPkWY4B3ZuyDJUuKYjnGvLXIGZ6jN7oSIgKOt8yAHW8802FFQwoMOGbJWq+HloaS
hkJehrqvCca6ZskE/8MFJZGwkiAN2/E5fIJN0UIkL27IutQsjMyBzeo4lLAjrsww
vSnRQ5paHjsk7DQVgViSPxiuR5zn4XFCb9o90tTJOrRTI3aiWrL1t4eLpWI8B84W
HUp/o25+ZY8ZoRtV8z6d4A1F/OZVjiFYF4QHKtnjlFrLZ+KT1iFa1c5yH79FZzh2
2vgoDnthiOl7iktXscgFp2LseTjpdK6pyRwUNdmQruV3SNKC6R1n1Bt6dqpHH2TH
pmnEMUQK8nQBAqnRbvmqk0qhEHZf0las/INFeizifXXQ32zGo29eAcpPF+U1cNfv
sgWHu4hLCK35PcamWz/e+wGDvf9mkBa0xRzNlCDjSAyMOyFOl3OLlLxGR2/ySgB+
RNwJEpzsCZcg/S7koyZE/29cp8jBOZ1UN6H9ctseVAqQA6HocKZf4n0J6yg7ZvMW
hyamFk+GSgu5d0rZDv5PnLVWRALh36SbQpLpG31Bc/q4g104DD0RAP5N0cM4teHQ
Qk4DDNeOnav6yFuBVI8Z9KvnnTjx2UmtVdACaEPBkdN74n0HWKqSXwusEG8Ajur6
/DCnt3395pX4sWlL2ME5q9qPJOZTM+1tJ91BdaTsTsSYyuEqZCKS6KDK+iPn1ZaM
9EPC5bjyNOlKrZK8m7V7orhKnHybLMG1WsO+0TsxQ+ZbXCF+6EpcPfJ4j0XxiRPp
ToyPYrjmJnA9NY+xv794VrIqRMWTdEQzooEbUG8EvECylxXmNvrdciogAzMIMlsM
UGabvUsfNY5ViT9NR6DoxV+1ap4eH9ULMDy6MW0jgb/8HBy8pLVZ+G4LXw2LnbAz
/MAga/uCxWvMYMpYg3gBzXrbZkLgdbpOwDg8vO/FoAjxHirHOibzMX43LFW8S4BR
ZnwHQZa0pWZ4FllYYq2K4Jehlqbxd5yZgWk1fIgkxNcEAdCoKjhJL63j6qBIqP/G
Xb9D7JbPCwU6rgPmSCoZlMbP/HgztPiA1V1Igx3dx3+TpEnfVPCrzTQb6J8FHBZ4
7e91stoZwgvCxhNxioWU07tZJE1Jzaf8M0siLcw57380HNXC17QzkDRE4pKmorC9
1za1gnuGsw/MwqKGT+9gU66hn2n+0Od/c80kBwt3hrA5QC5/LmU/y15VyRaQ3O+r
09rjrbBX+je0DILkdIfgw8vQPLuz+DK0iEE4D051V6AhkVfhYUwfdD046yU73jpZ
Dn1ega1S+if6foN3lyXsS5x2s2/uBSSN4rcPVKM3fj7NsCYYGOgV9pOyfcamwPFr
Kms+NxlDTSpTWmBfmkL46zNaO5s399AbKJz7NZxwlGEJq9Wkz84JpBW89nuCtsrT
eqXjDVAA2WB2MBlivdlQuvzmWy8WzH4+41xGpkIGU/UsUE9kS2owpG+SxJ4Rp66r
s3MQjR6/t1uygeuumGJemGc0u/mEneHvBclCNLYlBarw9TbRgazgZgccehSdTiCr
NdoaN4NRpMTMuK6pnQb1vhfG5Eqjfsvy6Y3mZG6OTNyx0ziR1Aa5cXtxBxqeCWYx
1KHXz2tOCHa1G1Z1Faa+5OCXH6x0VYOtIc4TDGnzYXMvSThcIDIeCFJuMasIWD+F
tD9a3sSfJ/7rcwirosk4x50j+FyB9Gi4+9XGDwvIm1zQoD6EWFcX0eE3M8JqH1Jw
G/2Q5vnlHW+7W97U8Js4K8i+IL84F8Cl/crHsDaaishWtHZZSxK2jJVX/LA8fMjF
03/1hx+wvhG/1ceTuHitpm9YAOTr1B8B1ypIXzAJxSk7ZufN6CTu3vLqgKagvENx
jCLYfPJgpYZ9JU2fQz5Q51oL+xXXBFmyGTQa38mXqUiOc6PPR8JxVOoswXJkwkYo
ToSE0cCFIknWK6Z9nR/mEZHXwYfCerFXoGibB/EVJuZ1jLl9v2xambpNzlUDZU3U
Pvj9LoUmxTQOkKrbUno6zuTJDLUJmhtjUgXrQkUJSPJoRP2rb4KjMhbIOPMPSH79
UVXjxO72NCEn+vfmkxHnIrG2Ccr2qc/nH5KRP2lBCLApMFIftKm9Ka8EqAO3FQuz
zrPnwIgip27BWweWITornSvtoOqQIoq8GwCBxQiBJrlFH5+x4jA+pgvfTRwBU6kC
JcGQJ5twfjJM8+SLKGJuFLcVRY48IBiuBCVHLX0RrAbE4XTb61LdM+xq6wZTXbzr
tVJOlwMW5Zty81GZ+bBhs8h+0mYs18rHc+q45NsYJpbE6omMS/6PXn3UUdhK37RN
egNWpZMSwBMLFhC8/4q0BYivhNthTVXC0WSUswBlOqLv6vP5I/zbFcCuPlqPDygA
eDTq3lK6IkvtFfNKLb/7xUminvan4l0w7Pc5Vad6jRu9O28zhbfk9cr8EZ7QhvSY
BNaYTWLpBhNlwIEKKmrtaIK2XD+2nmFey+SqQi1TlzidZUxELvAVzILw0f71J5od
9hbBQw9vBAHV/+CP19RerOsNqRm9/J6kBDdSLIK9B4Ceg75exhVDRrBPypbB8ZrJ
uItHLhenij+63HnWSfaaxM4WbM5GD4ju8Xz3U5U9yLHZ+MAISWqeMlUvwsm41qae
JaBsiYp0S2vGUnr2jMafXox4W7eulXScJqJ4Hbq+Z18h9XZX/jgTz/5E3EMT7wNx
QUUVeE6Ex/Rv5YqGNx1B0RmnxvVAgIwTi254136KAUBJqcZY+BjbyzlaZ+HBo3QQ
jUp79QdYkTEmrvAc4z7xBVaWQ8+yr/kvpoLqRqh3fQd3QUdfa0JaHSx6gbACykQn
Kyg3dfAIcMNitN6uPCyE2HkwX1+4pdZzI7wW4a64uDi5t0mGb5L8wmwUF/JZjUUa
PoZ+WF4m+1u6+mPDxggPGZ3VggtwlyIJbw8sTvPBZp4qgpXTljxpAsvzjRAfN0vF
NjpiD/a4UkVG2clckfoY0mEjVmTZN39Z8KdYJQeQ/wr8bzxwcROVyy91J3bfyj61
ph3o2wq4t8+MrIj7UFwGOJvXX2EUmKb+4sLMvZiAJdYqMcQKeDJstjPk7tvndjHL
daLYYFZom8tbPdL1+HUKgRkv54aQPUDqtWa5rdV15DoY3FIDzaqcQfUMRgaFt2hw
RhbFxp7ayQJPJqbGlq2eI6a3JvgFX7ozOPI2ZB0fZXrwugcxvCyi/rm8N8U+ACSx
t9NbxIvitAQPbTyJtp9yt1Nf7vzKlZO2lEySJjrnqDgrCfXWBb1tAxS62knZf25z
5/4BCnR8NZSSqa0p8ursrPDZYBdycBnU0J/80rnnL9nvNiC8XX8W8vyMihDStaWR
cePtjxS8Qzfn2yfJO948d/NuEg6lfCmXKCynMaj46cEuH79o/zS4hSK8B+ycmJGZ
7jllQ+k6KXMxZRh2KJVwVvF4Oe5q511+4/dnfdmZ+D9I44e+gsdR0N0KtrTlZwXF
K/QX4/9xMYI4kMa2+bquSHnrp7pHg9lXIDh1MpE4XMBj+LbK8EvBlDWQNU6oodAs
la+pemS4Q+7jzAxqw3hko9LmXevPx/dt+cwIsyjuSezYxBP+WYC/NbOVsN2vOPBr
mVhnwEGoxGgJzTCNC2i0h7RrSCWagmFIzlQ9j2jozQRbP0+TIr1441HdfVbmK7UU
Fv2n0dwK3/iCib7QKUQ7lXPg/GEcPW/8pzKsL1NXa4XDPZ3ExcgHlk6nJOS1LAZ1
p8Dr9NvOlT2ZZU3tcEKN5r+pU8zWxY//bPwNsB0tXUSsHPLDdp3nbWh9ITPMgdm0
Cfd6TMsY+ncyCr0bgByCK1rZmf9PP6+aOZgE4TUr5KpOFS5BFw6Ef8VIZtJkvD4e
Q+nyw9FO8VbKS4vU44Luk6XM/PERhzgaoO3dC4LKTu3pR2vzKTxUbIxG9cWJTiTA
ygmKne4yibQs9Yq90lroLPLK6yUPTQnjBBtYaUwlYhu9X+iOoCG9iXF4/9KfgyeF
jP80rp7VzhzktFGoDall1mCxl2CNA2zzFeFhOMniMLI7B5vp7A5Ec48cqU+2fn+U
QjGdVu1LtaAKphA47/izAzfcqVQpIhRF0lxx3CguLh25Y+woEDQfiyjyBY5DdJ5U
ET9iQMkbmJHx5W7jXoBchynDOXUlMGL36/E7qY+JPhpssXYcmWfsLn8qIZEbu71Q
tjTP7KwYi55HzivrWcsZnazQjkkYDUQhOa8DcuTiDf1/lbxDATeMTd7X5p2aZ0bW
6eu2jXKTRReEmuTuKaqCjVfnjxr9q650f9B2vIf0mfeT1a3fBIN/j59391PODATJ
cpkrzd7L6n28WxIE1RnXjNDBsO5BIbWwMKzOQ53BztQ2uUn7JvWLHR9Z7Oys625I
3H0ePvRE27piRO9QmJzyk6B+OAgM6wF6lJiA4qpydSlMz/cPVCoRfxgm8N5TTiWP
7ZIWzGduoyNDDw3geHhpIPJexxiIKNDWXnXw8bC6WgmVLxR+Jy4KXlCeFMRnHObJ
GBXZMt4aJjxSFsHS/d5EOpXYFeSgX5Lzc3B3xwqeReptxKY3kd800oQHT/4J4L8f
wyNgJhKuBFE+00clDTRNK24YR/KTHto0vXBjkT23QgoHbmUpOvpZAil3zWpL1iqM
v3hryoDHVbp29hNYTKSANEpSMjgBylPyEwTUogBvsj3GuxQrP+vQgypylwHxSMK5
Ea8ZaR5G2becZNEXpPwnIGk52TubBt6zyAMGkcIBercOAn8uiLbGLjXk8QJ9L3J3
MrKtBA3Laf8EdV81iPw5qd1rmeqi66l9nbeMUVKcOxBUlmvPS/DaIYHavygXFtv1
DMKSlefCKTcOv49avLMmbrrWAOzXvG/Z9A4voDHMknh3g6p89z54tNoEgvr5LtXY
evFCXc7oO3dvwB8xf1/cbdNWAHGeVPy0JraQr+ud8nVZMrkG8TGZrP8nV/VupHem
/ekpo08gadw2UgfCNgP2jRD3f3Yt8WWYUgT+rdmMInLOn1/mB64oLviu1uDEAhpQ
IP/koc2fWSdTdduHKddlV8TZUxgCfcEBjlSAZ8BWeYA0H4L4Lq2m2O9stdFDGwIO
UkxqYnmFJIQQzGGhTDbrisiz9fIoI+KCRpitOKnyqLWmTodi+hM6rHLrSI5ls7yY
FoaDZat0XztdYPprs+dtCIry8NB0Mq4WpHZy9euEWjFW3TB02g+64SWbbo2+1enG
gmeq5nQGCBAgU/9xtntu3SGVHpRJ+Rdn567Iu3ErNWUlUoBloGaQ+cx4cKgWpei0
al/+glHqMZG0wRUnXpE5aOwM6LZZMaPV2ia4iPV5eG2jfI9uGgMnL3kbFDZl1mag
z2sMM2MQG/r4Ho4CSGLjAmuXhtMewrT8bVniaSCXepa+5angtBMNvCG73z4t/xmd
iLcqZEkg6A+SdXVHfp69i6ZaAmlm+I4riMVgSj9OmFVOobEqPy4jRBK4+ERInIW+
1wzxu9SDVZtc6h+RMHWXckWR8JEKeX+ncL+sXMMtJCxj6tv96jDlRhIJixpMfr6X
xBDXdK5Gl0b8AC9/bhinV+wwMfOclx22KVxmvRn07wwXqvwIrpJnaAL71lHaZBBV
R5mBRTi3iDLWtME4o1DQoy7O+M0ZewckUpD9aISDiX+EOzCEDi3UeMpFsQaxrzFL
lgY+ehOlqvvryrt98TZa/MAGFHY4gq95Km0/q0Wg09MqclTbEA4+cfK21ajlM8sL
G67hoaDgw7QpQJUFAoG/JyJhx2paIgHfCeKGNjDXuLr9qmevHrsaB16i9gOneWMb
k9oXNU70DdickRm0ZaVO8l1f2QYRy+iHj543uVQ8iMDiFfyfj89fUgIRLqxWSUQ8
xGF2nmE0I0GY8K/5rhdXRpO84t9+6vWrHeclYRc7n3rjQbybt9kO0xR2MqrhpPny
nNqkLXvvrJmSYMIE0XD6OFySj7LuYgJTkERtCyCU1HOwx/A3dyvdZ/exz1OQi/Nr
DSagYCU9BUdannGg8iBTSRaToWPJ1MBjrUbaJEH+BujlcLZwmmkZv1Qq5T7liDH4
5m33QurHc24KEZgmb1z3AdncGNqk/Pe3hhObGhGfvaZADpjWT/ZIoOspbnPv0/Mu
93pzvSAeWw7VdO8jhR8AHRMNb4qo4hB++uKjW50exuiE47jq9L97dK+KrzwbxTYu
4196G4LPOnxLP2meACgAx1U+Cg6vI1f3qWojiotivqrOL0dExxoCk8RgOrW2vwWX
Pl/fduKLUHTWwubPtHb+2MCEx9UZr39P0hQ5r/+Qngxm10jSUHuoBicpIna5lG7C
VkNiu+dAQU4MzjHkrkzs4vE20kNIPmBbEFBBmuHlWXayMqOrezdpLu/WpmCjTDv4
hJZ/oKn5u0z2kvCZRNz2dTi8KG+VdIeHKEx/wZT1BGuiPYpZRsyPEvVr8higo7+J
qSU14Q6xVpNfoU+WHv5tAUNjfgwUsT8YAGbSEFZbWSxlHHNwc1qClILcu7+DnNbr
ZH/AXv4cL74FBgdTz3iA1nCSXoy0/XfnjQnWkrgop2dq6X/lWd6idbcNhi4wpWf3
ErTg/e29xJ17gaBSU0q7oTZKLfONZpjNK7R/4eXeV8Qgc7y1fbbS9m/axPSxuNcL
b7hISbAoG/4QTXe7euSxsZ4h2AakGTv2ozJiL5ooHBZ1/w0J0SG7b07yn96HwM8V
tZq8ZQa0tqfWgoMt2XA+1O7KZqXWtLVzKa8ZP+/xsKLdUr0hjm4gYptWVo96opGF
BiTFBC5pIlsF1LSLjNZTEYmmBvvDG4uWUNe4t7+RjA2gd31c5CU/oXItS4scjtp7
8MBcvcu4FB0iYXBwGs+ZtyiW2SSRr43XJZhMQUhrcpvJp93UiV408L/AE6UMQR+R
RWzdmQHGTPKp0hypblUUF7dCv5d1wd5rdg1qoV6pUy9L5SOjAJvpzrbeewaYVMmT
/Fi5Dbqzk6rCzoKKNDimp4ROt5NxvgENO5egIA52hV9dcEsLOd+YiY1+nYRH8KH3
6SQ2YRP+w2iPTuWNdm55y5XK8mFi5k/FCoGdsZXRZDaycdbIbLC5vSpBqOatSPlA
FAt7DfSTEZZOr5NllPa+81P5QYvqWvYOJTe9qayBrJHUhJzpJdSOZUOjlgdY8RZ9
fTOqjf+VyWIWjxfnEvf47cb+RcVD/RlTXtQ7k3f1Wp1vX68ZIkQinVHCL6lg+UdA
4lu0hw0PAKHN6HRQQEQLmGrwJmkihivk0PquSQbRrayaKwEETC5k9rOXEozs1/9c
B7iP4tC0VNBQPt2HbHapQWRkiX0vQ3SRkvxbGRNEc+XXqCYxz+XiKjIczRssDEbp
IOm6t+rCVOM25bG1SBdBckvvFgHzEBpUUQhhb0xA+knfwXVuk/vE4VepOcPCWvdg
E/6uf5v7n5Mc2kuCE9LgloG6rMaMvKa0O7RAnaveHewcb0b/Pvhjy49YT3iqUbAd
mAP81l1SZQl78SrRfZQHZFL63Ex7V2001J81IB2Yj6HjitzVWXUIW8TyhtI9+N0x
PkkQx8xo0ghc7KpnvTDHS2aGwTyxKxSf3D3Qd354KnCTCm/Hy4/wDDiaOqWYJCpE
YSI1IJauj9mrwhqcWpEPGb+bsbj/S0QvXxdMe94pwC6a8lzeJBvWcsnuahJydEdi
hW7lw8cauv+CgMkjaYPT8C1OzAkSj5v1Yuld6j/eoAD0PhNxJ+4yNumFAH3rBKG9
eHcoBjssMyVrmBRgOZAgnOCOVOqTD11RUtBb96teJevD4a6Smv4ZksCWYLXThkLE
z3LvsiY1r/CuqcBBsfBI8GVLpunlYx8vj0knCfOLtluVQJnczTQL19w/9zUqvUGO
iJh7PdPas+PCTAWfzIcTDmNxgxCftHCS96iZ9f5H0uY49jNGJUFK3/P+djL4krh/
zia8oMoG70WqjIDI5WHNGqkMq8maLsQZApcYSMFT3+3SeFInMpsnKtnH6kb+eNVB
eMOjx0E6BCzBvFVA2nVZOgfk8D0oQWZSaALZz7qzWxVaeYVp2bjeRPK1cdxYEvhh
vNNqJmcHDfkCnocZoO0jeGQy+gcFFCVgD4g2aKnYX0ZhF1tTev2cMKRJ0SpqILEI
oTTjYdSDl4PbHeLdcKEV0KRHGI9zPQpOZTfrcoT1YwfaWcsY2w1tw38QBkcBx3Wf
ACNr46rhr9ywXSDrcxNe/O1k0dQctJF87t9jf8Xg25DZxd0T+4aqa9SoZdKeF8F2
SECNFnrDn6HSvJg3IdxXLUDTbLRdrorHfhpfkoy5XC8CCuVnjxhNn+YkwzxL+SjW
zpNScMbAYEvyGxmyahEShC4bDOKnAurJNFVhE7UAeIfGDap7tI8sBaINq/v6M8lk
Z927NgLxmL+a3nKB7MlFqx91urc2mYrC/tq3dTUTH9Y92cxkuQVixSx1OKuM250n
lLMFfo4ShUUE8y2IuGh+PKkdj7YPvHKjCUfVjehen8XeCLZebIccT0QZ2o3PHlys
v9yfdrbgQ5xW3QkTej4dYFQIZy2lVe6ij2MorOrXd8yMTzymbeBEDbRcGbbhk6Xq
zB1kfBjgTCWixmE8ch3jiW5lwlx0GCyVabKoxlWwsjNz6BpZR0XJYNKvJpxZAGaK
QdsiZl0QGJRJJhgoPPxhdzPwSwhMuglMfl9bgEGCDka1MHlt2BFDJEciu8JgHY2P
kw7AkMgHnY4h0cTbSfLjLpoA3HgtVHfYHN2SgfIFToWoaN6+UCWqfw+pSQjuHiYu
ARrr917STQ2SVKlAzIYYVRf+GjOty/jVpAflpzpHCI5hnyO3we8fniVI7TuPePsw
rtimfZhk3R8YsOP94V9NYTq258vk16lg8uRFX077IT9xwAz6v3VRqKObo08TK1/D
FXJ56zp6JTOyVxM+wHCbmMom7YtiONZ9MEIvt7z4HqctcjzH+U7tZmhIJ3wLn5ow
36kZLF41I7bR0tpJugK0F1gP8tsXGVEUWhafVAAzoKGVCvcqOow/ZXLebNh4AMu7
SPGcx2NwIDg7BJunOVCgmsC9urK0Bavi/L7ON3lE3LbjPaNkKgqzdfRMc2tnLWNE
IIO+wmBNvYrykzeaNJ3IZjPTAMJz+BjFlZRQAKmP39cdWICiUxnTuitKVdHC1IDt
8q3F4MSFb3PMFVDEFXaMNPsycbdQX86IeLNWdUw7CQS4B0Na22Yf7MXZrkIap1gu
ldO+X0CA0buw6ascB2ZO9BQrmqaPrFFR7bMDKnzOyO3UyhGLAMR4m5bzLPCnyiae
3TpvfOPSrZsYUN5F8GLt0PGGFK08FQL1Aaw7+SJap2AhllJ20qEgvw6uRAVCP03G
/9gkkaSrEZgdkAyjOCLS4QEffgsIhd2dT0wELXD3xxMo9jdcPbR2h8191RDotWEh
jRSqtSlBDtUZvWgz7OaAyAe2uc8DPz4PE+DLFgNpG6eCqMNRlxu+yCRmGWmVjAGh
hSYp3xOR0B5LMW8lXXRFh/VIWqCtclN+ZKtR9cvnprqnkbgQ8zcgSEhQZABQKx+d
GeGazPeSSHT3+LcmHb9E+pm+w8nf2hE7VtJo+Tc0QwQHnoJxBpdijLiZtnymizQN
uWxchoimA6pN7n7kfZrl6twsQEmksu8WRL23lbNV/9/wjWeP6aXvteSZmm8JitHT
qHk6/QX1XdRcwPHGfdFc26mx7XADHuj/va5gsCsW9x5aJHPdyQ2PxT9k6MSOYgib
XDoS/z0hHrZfpqNvDMJ8YH2OeM7+qZfYeRePnppcwFhH1BIQ3LOgP0jo3zMXBIcY
fM/gF1QR8kbfLMyEuUm0Z0MMZ1envmfFyNSQJHxEgfQk8RxdA1OdpWmls/cMOCLv
U5GAZ3rJugvp80if6aqIPJRcKlG/2gpm4rlRKRiof5lcj66vjqhial6H9ytaXnCw
+3A1+NiZn88Eq2YinPrKQcxDr2gpL8CAgEtYVO0Ay2N7r4V5rupFx7UlzieR8mnk
YqH9aCA5e7Adxla/pAJc9LFNSpmHDDGwcdjmZIzNcx0Ux1Em4ZDnUo5zRZBFEzfG
lJjqL/nGYrFYWnG1BLXd7StNgHmWMk9quhsbYbUt4X4aIVvzjVa4JNNrf4zvGROt
3pH0fzlRll71aPMwGThZQ7I1PsjuFrondBPjeCWGe82HoTOuLZfLcBYBcPFIs+6R
pvHJQOHgprjQPpmhcXU9tvap7Nm7NE992DKkG+8IibxKjjiSOaXYlxlPirQtPmiT
hfDzZxuYi58Ca59sx7KHYrPsBgOTNzF5t06EJx9QMmquYDwmBZb7YCDJ5EgJ4p2L
XGqXP5Lna4sJBsEKaUHWZdvXYCmRlowdT35Kizqm3irRoh9jX5rzlkyeIoV1rdlk
fFKD54AaxsL2DQnXL0TBOu+T5xneDQSBhWn21hIopWFBD4rrmUZMVP/Hj6we4z+7
h8pmSiQwotfhjttwpxlyTJDgzM3rZtvqY7UFLeiNZxgyL/s4OD6dkJfjxu+40HTb
odYaUDHI/x5ALpJ6/mY3aGa5c6+R4wEmMpO/8aEiPW1KqoLmYAUrf1ev0rI0VAel
Y1iCO5uqjrXfF4kIlKFfenzsITt8HHm5FZmTsiBSUsf1Y7zPgmvZ04HsmqRKuCZE
QFos+NlfPM5EtLOVD8M8areD2qu6aa6p8Y/2BvxpaTmUP/+lCEFrm//cprX4t4tS
7Ozi0cK/vlQHLXEiaWBYhlElBaiG9OtWGpX0aeH/WyK2d57ntcBT/hACwPGwN315
g5NVdFlNk/wKMnIt/vVqZMXWXkiDfydNFhqHSFm6suUfksMKLZbGl+Pyh9UlQ8uF
V7EznPLtVuGazRlffoEehRSQUFwob6kuFUXpQnkBh/7cf44gdca6un8uel7IQ9U7
HrIv1hUgALI7ihXc7DffVFhvH9/eyhYUTRhVcNvyHiVlYE3bwiMqLIMj/MkIaoXX
ElTPw+nAdxQNgj6KDmIY3rpz/ktv9Q0OgUEmR807GVfmUc2xbuvAGny3C23YpZXK
K/lQa6zpYPMPP+SCHrDlHIlPhQIO0wlYpJScXm7nsyWlrwN+eV/++ihE0WU2bsXV
33z0tyf7YKRRlebs42zCk4Ng6KcA0yh8EqXwrg4wnMrYquwD1TYtEL3G8ZvpraN7
EmJ+d4LR9nprDDiRPxFjxRmm/2qNgM4ZPVUsQOP5g1eiPZuqg/sXTPlG7wtJXdmX
i13TmA+iF0j/vi06wQgRYopMvPbeHjEWhoZSgcL3SjlVRh8GVsy2LBXoq8OXTfpj
5Edxq/EhQujfXt0z42hkzCceunFJYqM/kjFh94sLSXicchbyJq9+xHBlzoYg551q
43riloxhmImk7dMuJNVQ8jjRhQB6OY2S3wAyeMdaJv97zipvnjx+fnarypn+TTxr
OLyGO3ZEDo+arEAJOQ2UWRvnM7tQR4Hr3cfmHgAc70ei8/ak9vdSYCjaGGjCfktq
rOOedLNQlym1/0LhpX2W6ZjDQlQKqvaLE8ug9ScphaaReZ4MivSO80V8Yk5ZeYgd
yJKL9zHhvZpRKvEvDw8veuyzb86xBcBNzNXbr8RLqouo+T0mx3bPZa1eilJai7Df
AjiH82NQHHHVQILpyeyz9ZLqOFqEGLV6KZo+YJd23K5Ws+Ld2jTY9wlNmQ2QpPGf
NTKTpqK9Z0jr2csEsGmYYO25GqE3fjyszUPZFBCehl0Ifb7Ya1wvrtgtCHC7k/DK
mW3dGqSBcxXF6XuVGNRN65/EzqDNQ9wh5Fp78GDTUP6B0FO8WmKoXEC9UNL6yUi8
O1hrvgULcQq3DuSSD7lJN+dqOVfE+deqVhEVYULl1KG4xWVUGbR8uYjaVSlDV4Vb
ICDryHYmtqEs4CebjhxMMBSVDf5MwVFyQYgnmyb5RfxWFxnadV1FHgYWIRPPAY9a
cAFRcFhx9EGYylV3ue7sz+zGf+qiAYRyDumQ0IaijUeA03t8gO+v6P1+arv/4eg6
lSzF3cB4EnUtOPavjT3hZxdEyJ0yQUAB3zjHXrvmqmn/bhAErU2ckxsM2+HNUjM8
O8hHIPnXH+JDOGHww4ffKygxH1rQ1qOAW4Puh/ZaVKJgPp7QL0XBaW+FCw3h/V8b
RppM+1ONpRSUM4r6YXwoJF7z7fWcGSBSIsTv+F5NzXm5KENLk307/d/SklXcPDEp
0GxLIvX3MI4jD3URYPeZeJB6T7ujWb55DfZQNwIH1xrhBEVN7kl238eyhXzwUVkR
lJoaYpPlF+Z8raj1SiM9xDDz0nyBLfpsCi7ZYLQeUHNMz3um+X/iUIqfD4avvHwD
ad/6vIKJ6i97s8rK7ynLj/IOMbRKbem5BWN59JKjEykxFum3naa21gcbeu/gTBBE
wfrLtXVjHoNhq9f641++MI5cneRa9IQ4qv8bGpvMbfwcBgu5uhCk9wYTH8rkf7tp
gZjBZi25FXZgXvD3Bu054AubXuRblghVp2fdC7VCbtijj2vDixyAd9VZLsvBxCr0
/yvA916qn21Bkm49z/kgKDa5sb7E0LRL4bDvqZddThbLq1CJed7oaQUAT375QwKo
dubb6MIVQGWXCtPBrGCsoiv1DzZ9lQzkh8RCv7A2pA+dRTKLE6G/FH+aHissmYcM
JwXIdT5MyO4YhC/XNbM4E9PMv4ypgPNFKJFcbYQukpejqp/zz7ACAfYbYaCGHvUA
Wne7YAPG5yAec7OluI736vrRjGuRpIxWu+k/PALSP79TD8+HHofAwNRQ/9Yj6TAD
/ncvR/NG/Gg3QthZxMOwIVJLSqzf7u9TK6BqUivkrEgYWPVSxBqiDLRGaob2kZOT
4H66h7Bi+KbQnLl7eWYaHWRKTKqIeK1ZAPRwhGhOQNe3EPzBAHcXIRgdLXm7LZ8F
Veh9vAvJaZ1jsyGMjOecCo8lPZlk+h4ydUqUpup32Gjz1MBGx5o9HSDLUi2KdLOf
k8/8SyIyOROQIa+etRl46WWd5bzaP/bl+3xuWjBdk6Zulm9/1NTfGBo419nFFh1f
7pJKQWYRv/w/TxPf3rCw7BkIDdTm6vFndvq3nI+JX8uubgBdlC2zPsa17rhPPC0P
vfH2LPM4JxZM0IGL1r44vRxmE0ZEXxVAuvx6yh43YxY3i4aZaI0zmwTKnMbfx9iQ
NbKOihtgWtGZcwa3sLuTNjUD6WTaR4+vOVYtpJJeMrcWXfy1xBQxaDzV1kMI5Xng
iHfTC44pY7LsQUTLG3Lgt5KC9S5ADARbUWXRXJ2kdZ0A6SM4lO72JageA9GiGe5O
scj4NLOetvqviPwmE8e4jJH+4fWRbnZukG+NN+/hpeyn03rv3l98fSEmpCWn8ChS
zwpVypnSP/hOJp65QZPUqp6YANBifd6ATP1Tw5fCLAKHm7S2dLCYgCIQDFUXXEEf
S2nKGfKDdjgOyxkQl4fZStzxtRYdLI+3vjpOU7R4cKTPYhzI1Lkv2UzJI2/KqyRD
n2AnXIca8eenj4RPueUf13DwT/JvPhs2TK/+lOay/UxaRxCU99ss2diNFiNDT6xn
pcDj7W4CkOxblxvDOMHIPiXSqkPSIP5mKH0S9Syha+0u+WrsSjB1ibQwkzFnWxah
cBTAZROlXcIABkXo86Kx9GiaBd8k+eONOhR3wdhSyGXO0cwEfQygxZgGIJUrJclA
5vrPwHdXCiyoKCAgKH8RYZQfDEaLz0atuM/2r5BR4ExIAM5jJ8j0aBjx4iq+6h/I
bKPmpyGn8PumtPxEVLk+dhnkTNIATsEh2kjI2ljS4xZdmnzUWU5UJeIMefPzuwtB
qAmhEJUUh46Xd70J3sGunqtDYuVFHpJ7c077sh0EQtf/FzesKkHahUO7J2IAUl41
QQSW2GQIKNJMBflnH6+LiknHTC/iiZJp+jXswGqwZvDoDV0d5hUna1sXOk7QZXA0
WQhup30YY16Hy+4lW2muipFFmY6Ttq80envi1gk544ddZGUAa+EVluVWlbajWvMp
tEPH9u41qhE2O8efWOc1pSQoFtmPfpuMAOXgn9zN9zTK3yODBtnbLRZfhSCIjxH0
eACanqff9E1Civq6TaYibMHiNedtWEpSWaix0udNv0OCMdebqdN4uXA8hXZD+1Ss
RDL9A6874Lh4qytpj+1z6Xeg+dRu/r08k1yoqO1VS+e5V2WtKdRj8ETlPbVxtzeT
eMzUgQgaDIR0QpnsHmocFpTrcQO1SSqwDVpmlDJYU8Ek58dQT/eQp/dlc4uv4Ql1
XUid7cfwDsIEGy0ZmMD48Dvzrc7bL85eVOHq9roLQiRznzrDoV1UNRzf9Pf3Zxkr
QXGybMyEuLEBgJGOwIqg4jMPhkUh2G00rzHHrDzpgWCUZ80b4TBq0EReMGHTHmQE
NWhzeIFhVimH09BM4NhRFZ4U0pJUg0vwvSaMdH/PcPzLNA74LX8LnR0Db3USOSf3
A1Ih/HLf6IIvNOKmVM6rQRwn07UH4KEQ0+xkWhYd/L7YhhAdm8KJxuPXajHpiq5F
rQ+0uQmhUjnMKDD2vDTDVA5Qe7XSMUdX8jTL1mxcuI/g/t8KNTjsIy3I2SwMpOQM
He9aH8U0NmWODDoV0r7GbihporM3AvNQSbSL+ctOPIq4RU3Tmku66FGcA+4cA71I
Mgg0uzQRgMfPIS8dJRB8p5Le3hPJHVNG6iROSyuu+1VXFYFNeD9ykAryRW7eKyO9
WyTVCgir81pfniO9U/fLInaV/ojkpt6zss1WmDC7At7kGfwoCJgNu2l7Ig5nDP8s
QfymiV1pqSh30WKsIAembh3ZFRLeOa02oR+L3ArLoWUdJF11ue23P+KUshKqtlUU
RhgpgVw+dGmEFV6Xwq7QDgY/UhRDahhjIE1s5Qd2kmHdbbd99mu9oJJv3KmtDSuZ
cLuOHhz6C3g3WNEdjADlLmxjhI2974m2FJpPkCxUGTl08kNh0NtYuCcvdK/exY+F
GHkuqu/F1sfec88FospGD9ZjLnFGkf8aiWZIm6m9baG2S04ifoYIkGgMROtHqF9N
0WO0qWplZPD74DjStlqSXgxc6yOBCySNnj2+BABvxEy8QZrcHeyNOWgLRlP38kD1
HotO0zy+h3NwUOlCAKwB/2inhosQTWCPJho401qLhS7P1wy0mthueIIE8fTVDz64
/yjKnmIm5P9qTuB0d1DwYjBu5Y+y/TtIP/aH6mdYP8K52pGhEyOzZDHcrw52gTxH
OXYEWq1i+vUyD+ZRg6CoEwBvPc9btOUKiDRkzRAxh+3VbnUr/RXMDdGb/HVLpTY3
lw3n9G8A071+kiIcP5xFU13ZiNyPbpKyqg1TlEwohKe7oiJZlwW4OgcIHXyhicCu
uVzEPVPWRkFupgogno5GxisDlV2gHTuKQ3U1X+H9vjUIYAXS2bf0qUqgyVaxesY7
8Oqxe5CQYhR6ttJ9sAlVKcNxjbXWLX74IYnR4miNCgwJlkRqSLgglfqoR4kGQA7Y
gsmJdTFWDrl51MybKwk2Q4U8WWLiKjAtSQ9jQCDDEdgxd/Oiv0tJ6k3Z4GweBf06
fr+Vd2hMTuenGM4idllIIYHhNCS9/JX84LyLGkGfAj5MPTBbt31MWufZMFqPNW3/
amZOMwSVAhIcIQL1s/NQT0MdjXCPvK0ggcsjy7YFdydkmiGE6TuXhngLSs+J7r1E
F4eCQ0XF2xJfC+lTkWCn1aNuENlce+Pw/oY9mIUjWVM56i5mVDVHc3txk9DYvHTh
LqDNUI/5jUqGHlaX8jqTsiQRkrMtarIls3XSOR+s+WuK1jRcSJe31KaEmWjyP380
tqQlEQCRgfKuOI9T/CJMkRv/hgvQkPsANY2V4606pbfZD8+A8WVk93fWfyFaQlwK
emJTyn+3m47TL3zjJWQ2ZszKzMS35P5V25PWMo1pbL1/kfajwJX6bgfjO7b9FqL3
IxHFvaIKFBltKl2ftS3TPHVL+PW4DFZ+r1ThK+90oMyw+eVdDTD17ze103ehReo/
2CLgx1Z0XsOiedyoY29x11r5bbw2oMriMGZYJTO1z7kNsJzKabbuWDI/TYPbt0Zg
8P2kLx5VNTpp5/0NnP/4NfNMdzeAxBjdYqFunZHQ/wv/y6IGioa0S+ClURAW2PAT
zQvY3CV9x7F74Hdkh4vsEBaXBHciyKCH/YW/hiInF1R/d+BuPRx+TMgrYb+yvGlO
TkWCZdlPlZK1/C0GozqAeLGnqHFcM94P9eZomTKtWsxGF4XcUydHSvQ3cQi2infK
dVGMRRlKQu3ojU0ZmZrZFLnH9stDmiTKjZrqtrXSHNZpArA2HJ2VFZgIgxuGxW71
TMpDsbRh1sQD+UQaVvpkhybRMk5suk7ums+Hc3hjXXW6A13ShcmwcTDqc730fHhb
W5um/1R0AyuDAKB8ak193t3OKYE3zQcF5pt4iOkpIIJQiStzIicNQJ69dvJN/4I9
VU4ql2IWAIExbjSlCrBgbh9EobAZ0XhvthTcmK5WeZeQkebzItlsAb/gmf3TFn7n
4Tg0qsSMgdXgbbFpieMhgHXKTzNvVwTr90qlZjxVQV7XgzJ8zffOZv9lNLEqPEr6
ooxTaEEqbIP+d2zMPeLlFUhl8TsGE9fICB6oYaicIIlh+tS/UzR+dJd86BhJMP27
pEAWPIVbED1E2SouTyMecNQRuTtuMd6r7gbYhPr7XYYGmrDpVzLrtfNScMfRKvJc
mBATL6fXgIkgS7ee5a7Uzs+XWFdiJVFYhHFIAamhJymYlRaVNIwUgFuEpfHjBW+n
iCuarDu7oMHIZ95uZOjmkd3c5JS12K9Sf29B5/GYAqs9tb7FM2Uijg2ehpSJ/zGf
wO60shDqFB6gM+DDxmqEVrlTy10YER1mrRNd31vUADLae0PpjrjZUE0nEIbSmoZ0
EUOq2aYEd4oCfZS4dE6KtmB/ANrxg5u2/fMIqXdPxxINRU4DUQbjXdLuISnfLhsH
vm7fcqw13p/VQX3BDux2bwutmoIF4dH2+gpnM2DFTRNJ0aPI54S8amUPvh4WByLX
NHaAbiJnWBZVygV5oXsd3UeRKJhNIUztOoura29h2I9CEajVfhyv2uWhTsm50rIh
6SomJ7ZLQDct387ZbM12ZplYKHXt45n9U2jH+qie/ACCJLz+xBhponFSLYTBWoDr
KYyUKW8dbHytJDdF7lCEqHQ4PP6sb7ErkXS3ni7j+awjgHc91Mgos/oU9ytZQ1qu
OuC6JQD3ofnDqtSdAoJEKHBIfEpi+QG7togRNneXp/lDHOt/6l+WlP2ilJB4V55m
j7yD5VQH4fDxc5VuoQUXXet8yf8jF975DrDUv2B1Rc2pDXiE7yBoDkUkbLIGk+of
nkFVGvdRLeY0phhvl9qO6gQULCXhXo1Rz17LvJ5Dqc2fGu0CELt0Lzr4rA4m1RwY
M7Sq6MfRiR56OL2xUCDihpDTBo+hgmftwNsQeO9ihQ7PkjTpRsLRS7U9kM3M2rCL
Ej3qDA4u8oci++OfiIGwRv3WagBk+SBqJqptW/9FhRm2o1sNGTtm1eTFCYGgFc4T
z7ghR2/QQoNK7LuphlG5kOL58DnsUpuIdCOdCIJCdmZb0XxJoTG7aP/FAO/bbz5H
OBL0B5foc9q8p78DqWCMaJ9vyaEPTIAWrnSpIS4BcyP7on4invU8xb8gBHGr2V0n
eK54dWzC6VLuY6WnMu6mvLgbbLAqLbzC/yZI/OLWeeSKGMvCBI09iXGFXKgeLGHH
NuwDNaxfKo6PF0kukuuQKS9A0fCj3Uo4xseYsTX2gyLeP/pmgblSFWp1ZPDyBXJJ
7psaSV/Cb9Stx3gOe5Og5gLbXqB01MvH1+gRFOzfZwVxFmHV/fspQsTbNY1IIZq6
hZZDWGsUZYYtUWaQbnFeSTq+Kc2PfCJqDWr1WjoA++5aZWAwPaQj6kr8UK8UCl5y
2mszDrVQmbXgDiGsMdzCzp+YmdDP3tXjXJsOnH1J00DZSHCIgVYfANzmkfNMU3Vc
1i4bTCE8MkrHEAL5osY2nm/f9OLzksQvEoG+mPZ1AIkVD49ptIypvDwuGHpU8nwt
lA9xhj1FhZUp+BDba3pxPAljn+MOh633DVQEld12Fr3UPnvZsBBs/GJd3s5fXn3I
711r/NUM5/w7aokoqqcBlpLUxGBfaXIYJtdY+yxMFDYH7gJuaCt2aa5CYsd3liQh
hAFyNQg+NMt0YaTpLIRUluly+Cbw6uFe8LuikbObmr9FFJV5ExY8sLEy15/dRoH4
XVZkAyAA2HA29C3/lfN3Vwk1WHwWAaVqAxr6JhKN5Avhh9XrwLHbsqGuxS4uBduN
5qHnX3ask1tdHcHcXuQyxLhVThnV+hPeiKKeoKpczJam0y4aaxBZ72NxxVK3rMye
xVPCbGiE9n+ugY09oED45EI1wxBcUgVZ7tBoL7D2XdvMDzDSZ1qw38EoFUKHm1ea
41FFtTAmfAkvRZZWMudIM7FKkpVNchPtEVyB2zaiQ3/PtPwcn713LSX6VLwUvTHa
PKyCVi6+uOZrbz3sBD8v3Lt+BIOF6OI8oascAxTS1EzuCiHvcRjm/YftyBTrxhHH
mUGh2xK8eCbhPS/J2Pvt3cUQbK7sN0aQWv6G0umiYWdiFFe0Fy26CSM5MqBbvwwD
81GjJG2fSrNI2/CkmQ5iRGY9cbLJp2XkmN16VxOordqGicy7wrda7PfJtY2QEvf9
keZXrC0KXTh6W2j3tXFOKd3lENTLZBhevtQnrvgFbgiYuSeAcKk9ZSasoRaZrlgP
Pi3fbg+VTDN44jpeWSzP34VmfC14i/yvBHE5yDZ7SnTZxZYnZsUxlC32ZfvRiKlo
Ec/dwZdUmhK+ycfo9u0CLY6YH8WR5r3aRdghA62qixDCSekd+LN5Zdwb8BOHa7qK
gP9ZEQef3xkSq2jkUzHSvuI5k22mXqCSx1QqoUSm5NZkCOMpdAebC6W8P3BwHVVj
8S9jmckHCRgmXKa2WzvATWYGDRlLCSqfg0t2rlNwmsIYKayb6EW4CuN8lD/C4AAX
plao605PcKICYNDKn6B8uBkRVSg85IkzFfaHUDfmylxzYjzxdB8KKLZEcMXnW0s5
GLMLDwtQJvHVpmYijImJ3EPsL9nBFeYyfevjQAM72NAQ3GZ9ye2uvpuVjqTDpik6
j8rjP/0YCynV/nhMTWUVLk1ppXTF8U8T4eEE46oGi23NRT8b5x0cFFgmw7iUUccW
h+TyOhpIvHs0DVi3QBFC3p0EWFSC5X7u0S9DVciAOJ89IG8AO/mv4RGUs30b/zeR
J0IXWPdLEcRnmpKkuQ3um9EtoeX69CmFykXLKeQDEWX1aiu6zgsUW771dQ6CV1Ql
Z5muSvf3LVVMJe2Dq7T8sxOAxWRbiTLnDPKqndCY2d9kN01IIS/ET6acGh3kpxjk
o/CiDzASgBZjTd/zVa79ubNWrQY/L4PfvcBtSRqAab+L+ThvkLlrWXqPIOr5ofE6
jXmO51loc1Wb5BYujMV7JfFcjyF8YgwIlYUA+zbdL2rcdGw+ZFn0x2x4+lkIY0Tt
QKhZUuvL25qJWR/a9a3x6HHgFLUtTWXFXjGgrUG/yrg7fDekgl+A1NcIyMADT03I
h6wnIeQ47uU8gCPlUZC2niu+UqQwuWrjqa90+w2VD4BxmnZbndedjtOjSB6VwcOO
Vu5dDhP955JuOpfT+gVyFaCdh0+iNdWnGjRmLNV7VMxsTysKAza/GZNbgC1BrvBp
5qArrmJE4oI93Lx/pVW9W9sEZzz83ELqi/rKQ4wp12Top1ZVuT5K8Y+V95d2DYTZ
2QvlsYdBM2kifdo+mS2kiYvNrZP1i6GI+sPf5zCB0+31ZE7+0IcC0KC2Pp5UKUw2
i3Un1zfL39dTu8TW4MdVx04iDvV5o8DHyfr8BMmUPFomu1HtloGNsWR0CJGAk00C
m4BoWrpaT11MJTUcv6dt22oMArpGBywRt12reXxW9WVntmH0dE9g6MyCiJSNCC9A
0Yq6nWb4p2B9WVHdLBRx7GBiXHanPU70xup0eN+2pCC1Tw2FU1uI0kl9/1uW1BGn
+JuQBAbFxaigiSYTmsXKBUqjGovqHtRlf7Cywu4gKLNlYvSqzsgq7Po0IcWnXHkS
8HTarn5ZT7zAf1Ox3THH0BUpR8SLjrdqJ3uwYQpng9nGhM5SseAsj0B7c2Zwfl53
WxNp2PnfExW3dXKDERpNcTgIHm07O7ksyCLLe+CHodWm52wrcroLkGfpHKByhV4z
Ow87Xv1CY2wXZEx46q8tbieCsEeSLf6BI49MlIO0BrWDPgfsejJiLkLcZ1yGy8uB
jIOqP5C5yikAktT66iskImG3UhNbs5cyZcorPa0yOpTYRM81x4QjhqKc3mTLFjQD
wDiSB9s3Cv4ybxXtbuHnlie8R9wzC+PRAhY5Y6aAs/RbkvrODABtVxVPqmXC+IxP
2zWhDEtoJh6p/kbWYdHC5h05Dbv0Ht59tIfFP9bWf+JH9wVKfMhfe//aw3ypeMZ4
jJtZKg3pE6kVc3MPZGPCJggotzDx2O9sxE+YbZwbkg11IRsCx6hVBQnVgXizi887
ktzXBX5ypixK8YyO4R+asba3D09EeMmnQALx9ND9c5MglDrZY8tNo6e4PE/4i3nm
fgD9xDl7Stadl4C/Rec4KV2Mb0NabjivlntVkEs1ml2Yctfk3KUyljwVjQKAhqdt
yF7RGfsTlyyaZMpB1HsIUfSzKkEeAUZfCRNLdULqK5fxFy8psfmlSl9v83vppusE
B0gmyMiEY1ov8zgw5mxHTbsRmURHfwi0mEt6UB/PjgKHFwS5SxLmlWsq4dlOifB5
pYImOVlLPcWG/dOM1ABWhIrVKytCPjhvPRQrP6CYK4sBCs1LMUE3tan5FrONBt8t
tDNsHF+gMpJWyLU2M7aJzVr2cIh6XDfL9WoUmwtog8JlE4yIvvyVWSWNdkyYjsDl
knU77ta7bUuCGaCXheH77xx0I7+fZ0DpKrIw7tJMQ0ynssVvzDIQq/xouAco1+XI
FDCmGf9XgeHsMSrbxQ7r8bcmHoDG5+HKvSjCM7QWn187RBLuCIXjqtJw8RTsCSf6
VxSCMDkWuTUis/1Ga9F2W20UaUWArlL2+zkYTiEhQXk46ziFfE+Up9Tlo3duVmTx
mjL/F0Y7BE/QvEh6k/6v//i+DexmUAaoCbDY6xjUVda/6uZILvNuDh7y6gkMrXXZ
yWwvzgjpkLhkuu0BIkn1b3nlKFhURZfFDeIKZSWQK5eJRXog/Dv5PPgmaIC+stGH
h4s4ZYFLJJ1LbuMJCFxv0hXQclk8zoBXnBKoFm0QQjGyBzfZwgUF7TKDg/+OnMpK
ecS8xgNItJNh5Yl6ZP7eujSbOGi/VPA8MjBTjtAaJXeVkYbrqosNqxNNktR9xZ3V
iIYQQ2qAJi2YTIcGDCXeDwZe4O8FhNC91A1jJIF+RA63naiEGgw96yJvZS/kyRde
h5REsrlquZ3pPNtxBZYPin19fGCSaXxUGeZ5WKW4wGqmRJ5IRsRD7sUSY3xS3iyW
ihKvOaX0+2sthiciGPomFlcd9tNRkoZUuubg2s9A+k26fi+KkLgOZA9RiymO/iGn
Z37bskIlShqTX7msZRPj7gIpUBD3vgRdYHbalbFzY1sp8frvBSt2dSUF2WEJzM+Z
sFBKOKxVQuquEqQS4lJx8ckzrOP6P6+n/kQ+HTIV2pHts9hQOkHXjO61YaB22fgj
gGHj3ZkcTSx0y9jS31Tz+KyANjBH2jFr2EhM801FgovfwATj9fj89qE9WoXdAWGT
coglwvTY/qb+odsD87gczfK0tRTyASUB5UqEL1R5xkkuYN632ASVxFqBDXGHbXKa
4BkqaqXkfny2ZjXBud1cklI6HdE0txR9hr4RbqM3YNYAojtv/VJKywUGRygucm8D
8SLmLRESvb3i/UDBKUYdzWUz8h79YiAqTU2ASO4OihMGBDjQY3FgsR+y1Frtv33y
PfOLkECVDEPHGCn5XQCdFt8eR+Vai8F63sYl3+C3MnVZUHElfW8r3CQGN4g9us5w
tpmCcCpxTYAnN1+gdql/8YV7+jXqTEIVYGkkBhFzQS4TIbyQUV72E8PDLMZe7r66
c8FNE8Xgoi0qN8Cu6LqInWO9gMMYRoVVyFriKEXQdANmHPXslA3AwFG9ACYdVmXb
ZlKAB2+KAdIIbzrBeSNzuP5pVsvpfnxYBvZJ1xX7/SmqduwnWbK060fYR/GvIVjB
CM3uV7ySoGedKDHqQuGjQ+4f5sldyXtFX/qHJnsEkhJWXCXcOBamui6LF/T4qr/r
PObbcUbSqjPmD0/KuNbB88ZRHlr2iOYDiKNkWr9PNYGBf6yd0y+fQipaDzk/NINp
waKXrM9BbT3TuMsMJcNhxxsk89PQFIeVWpnZ/vqn5rAKEjlfygIT3Cig8FV+ycD5
E+1bpse1FS6Mweue4+6BXBGa8TsT2MjkG487M2w5Iu01szr2nkJlUYRGpn3dup+u
FZ0uxvLk4MEpakHgmNsQXpt+w6KwbyNKyGz1HBt63JMNolEUgZuzV/PoJ//dYkRE
0ftwokEhYoBPv3LGnP/AAL1OKDUdcKqSCSEJtgp9QOVLWXqdGXAhRcZncVPjPIHT
R4U5fvIOn/uen/lTC04Hu25lxtQlWicZPp8Ies9MCID5QJRQLXrRxRBpuMfCF1Ol
+RZ53BnGrwCGWCOfg68V7NtH9gAzDtd8bg+AvCKoexXhZm8sDx/LnLDJerCNHuzK
1a/+10+T7yFaVi2fhpU+3dzBwt9xry4kRDyzv2KYX7ZzDPZKlEcBIsupa4UuTkJT
r1No1lnQevnCxK8Amr501y+xTtYGnwPRHjfNUlvnLn4tg1bxZmwVrUJG6sNTIRvL
B+pMNHCUH1G59OoWwlr1BXv0NQarXNMHuStcMI4By/tLC7fm9crom1rB/QNKRrkL
rKb/i8sispTLOJN/eV1c/asQaS1QeO2MvoTZHsrAwxD75KTProd5MQus8Tax83/r
iK91HfvAToGj0rvo7dj92mEKloZH7Dvin8QvDYQDBW6SkHH+gKIjbXEplD/xXO0M
leWepADfzlQ/Ne0l6ecCcCNTQSlfLWBP8UnWXzptBNIxGTRx6meGXO9w/cFjRLwF
xyAqpsZFrF1IDrWkXUtkZvHehbBgyx4mMJ1wikD+zE0yArMIq/7ZRfX5xHsghSCJ
UxfzkDvTaNDGdmbC7stYnPUpPkV84cjNXpLEpuWEnGeILJe04U3pCAegXBEN/efN
FHlBFu5YD15LCrBti47fcKWeKafrxVRd+MgIAucbtnWWgJ5YE7YLQOikUyAahsqf
fWJmBgHWfM1keoEiMbASWGMkbnzJj7WVAk0n587f4Es/k4t8uchGxHCmDq4W6ty0
kj9gvgZzqQsE3MThcBTBStGiOsnzq3KYxNu5sv03HIhBo9Dpo/94Yb+dALQQKcKC
5YitJFJ+Kw/5GdufFJETnbedWr4+kOnDdaEoTTd4Pw2QZp3oCT9UQsxQDtkyTPqm
hUtGD/0azWLGOt/mC9+2k0ccSqzI8DB8yZ5ADblS9lYYTku5WKzlxJgKml2sBT0g
rPSKd/GG1GOoxAzoDu7iid4ZkSh3CRyDmkA0bFmCvkig7qv365k+Xt/O/+Oz6b/g
J1jr/41pGVMHZcVQEK7XD9MdFFLe1Bu9jfcLB3SrzL5+nqowgTJKQK+I8td7/zZb
xjYefG+//hNM2YJG6G3Tc6fMDgAKnz3z367R/7HfCTszePwV8izh+tKHZXpp9Ar5
3coblHZ5HQAjQ62LB3M06Tnaomk+gB4ya1wHKoj7LeG6GIw1gFgcI+OA41DsaMZA
s6s0q4qLQ9/Azw3EWiSYa1vyMtxQppt/eGdiLNuCYt/iO35lzi3v1som+KJ+vLfw
X/yaKLJlkox0o3szm3/Lp8O9CNJLHpWc3VyoZ1Fq/5BpRCDwutMJoYNZ9xYnZ7LW
9Cvs5eCZ6bb9BIpR/oSS0F7/pInyBtWIGooTlZfv7Agm3EELjyBVH6ggqYJWZMVZ
aGZu3jV8BSa9V0calCcDuVuaYpBr3kiNprj9s1pL0JEi8RvqNJVb4O8iJvLe0DZK
ikbPSmed1pTyQO7OK20ANjmQUJqbZ7I/vt7Csu2Vnd34sAGFjZ/IS5drGxSvZHb5
icrJDt+ZpyCDKdZfmO30gunJQbGIVaMb0RUbAn7ONz1RWHgvab+jqhksx41IMNX5
ZHNHVkvmWChiMznJpYyUdQT6IX2J1csBD1TcIJU6o4nkELJckcXBbil2L1pnUw69
oeU1n06WoWGoWvVYees2bE4thHa/qg0YEAu6clPoamorl/VLoI7cKQ6LaJ4YTW93
gK2b5WecKBhOy1PJlu/yLEcR1q/v5Ay/f+y0w6uBv49Ew+J52euKF2XfnVwx+RT8
D0+TB3iKS16irvwWLulRKXMjKreHXGbmUpCNdV12K3l8NGZPKOhgRl24OeefrqWK
UamDcoDN+ZRy0dTnIN0JB/WsgtY11yW3b2Ikxb+++0cQRGxGs5lhcBooV+cE+yKQ
B0oxBvewaA9IfDtldP0YMc8z+fhYqKpNnQWWUqpL6FLN563sN5xf9pUf1BXW2P9F
kdZHEija2Q7BMpXwmIk4RsjVlUND/DoA+ehOdZIA08ke7pYu2trRh0vlOnEHkoQi
aBSBbU3G20XBGANRgLzkIHSN8yZ+T96ED6leP1376PlQVMSuZS36r9eRilD5LUao
K6Px7H/H7hZUxxPOgcBhsKO7nbFy8b6Dyxfvmcs4R2jC/1WmOo7oB63qGREUoM6L
bXAYKtueTW0xgjvqTAUW0BIgGSYaYOX8MfWmgScA6DgXPHEitLwkDnm8d2B5G3Ym
svKDIpliVVeLylh/mL8duPr9NGZfaIgs7PggFE/2YMkoXO0CIvUObYpHvpZFe8JN
ytnIlEX+I8/NjMAQOiHEALdXlieEUZiNrozXgUwepqZrS5YlCy+2QwQ/Ha2G9wv8
h3XMHp9msHhke2mUe5/O0Bem/PSWHUFzmhL3Iw2fTvEHBY08mVpssJHQsA6ef4f1
bogrQnYgJ6wbRYMohGVc6f9Fgw/9pI7MDkPAs5c44AzaxS3GMZZWTy71y0ZBi4rs
vKKqXK+Og/f9KocAig4bZlNXACJp7B/k7lzp3Kzq0StTkN6hypprgXs0RE6okQn8
nF5dwz6nHAiBSZ7B5xgcSW19ix1w+3jNcVI3BzONmUPMcYgUa93wcSdrViQX1yiv
ybiCWlKZp8ijTtDA2u386uTyqE8iQE9fyiCcJAuUCuHcBF1/OzI8sfS177vwNFCH
wi9CDN4y1/3nNkNCxznll4xhg9Jm+/NVS6AG3ak0YGenUfwccnzdHObCu9D7gDOQ
afe6zGd5E4sj1jWjxGldcL2/1d/0EpwuAYa2n8X9j3UQN10oG6VeQiP1Rz6FvZqL
WuvMTGSQ3cSoWuYaYvneTaBdqWncCER4pI0dC0EvNGbbjsabaIsGDv+7KtZg3SwB
skWLu2/YmkOOAoJ1V/oghNAjS98jh7HU0cTkHkDODqBKU+4FSkoRv6rbo1Tl9Tx6
iSxb0RDdAguR7jiW82P3UHb0nDs1441UXNvr/IhRUQGJhS4LxHpuCKzJu1y68JfM
OZHegghuM4tCWg4mDNBCH9V9LBSAeQlCoos82d5GJUw77WSfhr2YAFsJLJdwmyqS
JYgeHzgmwQeaL9GpOO+Ymjm6tSwVxQNT1FTa/D+TkY3s30CGBDYpHn4TqHB9BiuU
1LcfdYbu9c8btmcpzJHtK8/mUtDnIi/TKqXp4WLf5Tauxpr4lTdMLw3Ur4Wf5ewZ
bo5sK8Ifz8m0ZKtVKbfQtJtHq6Q9rhLuuTGOvE52WjP8vLY9C+3GjyZla45i9d0D
XBRsjWhPTPdCJceA7SSPdnUD502N744kN933sINgvRe9NSs80q3IPv9x9D1B2Xst
bKEMkJsZ2ZxfhHgiobl9Qi8GL0VJ7n6bfUoaJRDIO7XUieuyzsK7BHDd+yBmJQHW
Sy2K0UDGnovVnJuNrl9VgY7mAPT/Egv7Z+TsIfdIwAEZQNN5cHf9t6b8O6/Fe85a
woxpvzCPKJnSX9JsozAmpGVqg6HJrqiFOR1LVIqjW6TJP4iI1A3VD9SOeg7z01Gl
9nUFzMzVBuo6N6/tRlCvCAfinj5rhksU8W8Nv3tF/AM262MN7xL0f5g0Eoc0eBLW
pxPKzz0INiyonWIHj8US2v+c7W8BikC/hULJM5VOPnoQqEb+0spz3dk8/TbBBg8Q
GsS7nCJ7C5UCYkB5uCSwyJmrIG+JFfuaXlm+XmgzNb1d7m/1XjKRLKHzArzNVOFp
9WxBwAOptWQ14vB24qoZDK1dYb7gAChnz0cYJgLRdz8+6xVmCdXih2+npBtEWdQ7
4aMerXAw3+k8LBOnr0ca1g5r010Dt6CxXeADu1l9YsknGCuJvl4CljII+Rkf7Z00
pSWJa7n926JSAAWuxGQ5Xaqf2+R88RAbyRuzuEGNlhikpEpB77DCrJrTP3I4xXKG
yd9iUun6S7jifgjd7sRJ+sBFSI0p4IcQc95YBCjqIvQ4/PjcxYxF9/0dg01cvFKh
uLRgbQm3AAZyOiZn7BUxjG7shAxP5RLA1W6raxYS/SAxeMz6EHOZwdHHy0dbXznG
aOyVc2/brR2DXdTsvRqzd/vJ9C13CuVXkAYLgFGAv4uIKYGfPzsUZOGbIE7CH0AS
KNBDSrALgPdnXuD1BF/iXYLgutDvniQxcH9cRCtf+MvGMVIxmMJU7mq6+ff/1oZX
IT5CUvWp0RgDmaFpmsAA7olzpaysqNiw5VwgcZUmytJXWW3saKNMKGjUKcdWLwTq
OZ5n0ym2Je9YWiM8WT1keMaq+eIsUr2sVY0Hc44fEBaKhywaSsVjm8tllznNq0vz
gP4WZyBk/b5n8Oau1Z10clMKCZm8gOeKOl1kWphteATpYsxOdc83lGmPkzA0/6Od
kOiKjftvdnI6JdiStqhEwpDcdBWMC3vVVQEnMhWhWz6aOf0oM++Nfl8cIYSrgmd1
TBkeLT2Bdj08WxJ2yjGbBpicjDt73gYSizT3XVYiR1zniXCW1jYq5z3tLTKJFApX
GBEKaitb3F99DN3HgmBkcO76OpL4QkHcPOtQdhq5AXd9VHDPDWAoP1tPUdvNxBId
5SQrFipHOjgfKUODoVxjG3dVqGncD3iGXO1O702anmTrGaYs6RUdH6/5oIJbVZSL
R5JUTrXPNdS6iKR25jWAvdabxX/6vZxa0FSulnZmbEqniCuZ5YrSxCjr9cb4DO3q
VdShUWUdQHaibSLQWjCYR807nhD3NUhgP1ZJ0QyqfsrqJOo6UIEzE5FtPJDR8Jlf
qTJj90ZhEuyfS5vdAl7BRDV5Qgv3ylQ4qmvxq0FD69zTTC6Im1ffCN5HBb3MWh7+
KdFDVrbRc+NHEGwd92MXqGkDytggYB1JXG4y+efc1AN8ZEPYJmvDJ44WBcG/5rN7
bddQsxcFHwxusERhMZsppUc4QL10A59gez27su0/zSmdfKqDQs9YgUQElBFUcgXT
zSpPKlDHkNacYt7nHJyZJ/cFuyHxP+DpCYgAUD/c2mYWMtwgcsx9IlnOg+nKTouv
tbcHLMnNy/5/uvkLNQFSPn1tcw84gp25WdmJNCeCxI9oi615hANyqhxCdtP3Ve/c
XmslV0uLEad4MELZ2CIMujQrQnYCwlwmE+sp82aBBZduummW5tAGfRtoRFzvZLSj
CFEAImbdh4Mwdo1x8dzGvQPeC8+7uwxRwWRcucqmHLqcn+0LZfARm1/Qm0i+CcmX
AnSiASX1kYYEwqeVuSxCTpE0F5Y7MOajI6IOD+OG44CAfHQCHDAI8XW4rbB+rqZz
HBLVvAdeGsOrQA1FUCQpfTYJ+1H8EN2bWcg/A+f1jzcAeZuFmC0uYtjtH6U8fHEq
7Ng0KMsHBJs2hCp0dn9E5gLmkDsSCEX6+mpqxe9hH9y9SJ9yFRU9Szd6ZbENvLWg
ug3UUlJPQH+8Blzji2i7zk1q1pk3/AameIW7YXQFn7vPrF8jhI/lQ3gA4SnOUMmy
x/UaiW5Os0vHkC172QAQbjALQT42XywvNPS2phY4H0K8PopJ56DrieB0/841mf/G
WSWLuS08l2V3LMSzbov0EXO8slXQ+P4H1UpvAH/ie57b0JATXqmjogo0PSxAKK4n
33PJ4yJ2v2hWWIUtGRPm1I5r8zuSw9OAW/Y1Efp27slUaNpZSa9Iqf7wE01AWXC+
JI3ASgFlsVpSLZWh4iXphtfkULQpLB5Msyx2Wn2S+M3kdMoZTbWrC61qY8dVTqtJ
ZfqwucQYqUfsaLwC2qZLOTBx3nyk1qWaIkdBwrzgxK050bm6g9hIe3E4MACzScqj
QwfaJrNjYRL/t3tBPL6AZERXb/3g7PPM8U64SCq3Ve5+oclpwFteBM4sdTTtG8s+
tVQsoFMHq1QSbBTzUHV8YF20+YsN/tPlvKGmiotD5tKVyfEOvZwjfLc2jnDpx+eP
jAg6tppvj6MWirRAc4XwezNzDCGsle8kWeiNDyu4KbzOZrnnapA7q+XDCwPNpa4a
daO3u0rTrr7BYHEnN36SYCvvk+gKWAcp9pvSYjLGhrHUhWfpjiWDcQ+LHcAhsmGS
YLG3dgMzVh6mOutZcAsA7P3EfdliKa0t4r1ln9gTHxw4ExTol4UdXBqaQOWfIZvb
Y+1pY6BIBk4bStWQeY4hPbR5SzYSPM6y4yhPdGkLcwXvNDyRfG4Xh57TzxICnAvj
lz8CMFg6h2K/XChAp2wPJms+xJ7uXEP5L/KNHqyF6osoNsU/H48+9GLRiZCuMohw
Cn1v6nKvf9OO6PgC49svY204jZNAPVD/NMIv3uo0lj0k/Nj2ad0CQy923UpGtE6y
+UgjMk+0mcSX/ykCNrHGCL9KMy4R90xPa+BgLx133PEeRNuyu7uuckGzHcEVf+wL
Vu8js8RP1ID9wXg+/hIqDTG1cwxzWVMenoxVn/tsZdE5NFkT2J4+05zFvVgKHeSn
/k1Gi1l3GcPO2t6BuWtoZq6bQgZtfLmgo6nNQOnu9aEccv0UlS9Y/lkKRe9BKXHU
uMoEVoy/TLPwN/YCcMzpQ5GttEj9wSUO2/4KmCU6DSkXN9ZWZUhN1t7QtJW+ZEKU
BerSaKmUPEWolP2XV62ugVEjnv64GkC5p+A1cv5tUAND+qZswYPokgKfXiN7VJ6G
osZVe/8xTfTD9tlfIkuKVdQQqpMC2Y/dZ9IwHxfQYjYxN2Es1Qepx7N4Bv8xmM6Q
6ItXVJQzIxK2qqpI0D/JPyuHQIiVYyT0uNWsSWhV1S8K5c1hoeGBEbwiRLYJwl8o
9JkBRIKDuwm7Ojeyvn4FRn6qIHxcELbpTH6oWhf2tFcPPL7CtJDCA5gutFrLOgvG
2OVWZ0NAsDKQZ60s7XTQTXogGZN0lgeLTIAV2EtolxSmigxZ5wY/jeQ7+8S8M7AO
nnagT3/8hqCCEID9iNaTDda9k3SUxwewMbW3jy68mYY6yDFAIUhV5gOGAKUViWjj
XomX8+pUSJgeMMleQ1F+rIiLAqVUwfEBW7mmBxdulaKvXWe7nH+ZrvSO7OdZWj7W
Xtba+IxCGWQJj50tTgqRjnRSrXwB94onmE23s1nPYaT3yvOP9Rb8fj69N6Dy3GX+
1+VP0L6ZQe2S9Zw4pqqPy9jNYIY4qUZRJAcS3A+40EMD4/wFIdrwRXUFORJCL1hs
lsY8WWm/i9xF8As+hWxkDYgxhzTUFZVQgIErN886gHAlMQ2j9c1942UYHLmxc7lk
/z7+ZM1RkRN46nyxnknQUw7mpqIbT4AQPsZTJWe91kVhXH2RSMI8pFMZEQyPoSS7
a+ZF3Xngc8EKlCrgxQeUO9bTdd8AD6twplscO2n7ootHIJBXXxOF5csd4m3CT3tw
gzwLKam65GMpPDlQ/WwWBqAwGv6S+uvFbqIWniBh7gitwEksJlW/ktElq5WqEeo1
m4Ux3Iwe87j2Bjgd6SrWn8/1QG8pbe6e9vzmg4tfV21JJ2/YBYnm0vgC1WCuYRYz
yUJg2vowIlCmwTe9OPTLYa0qeXgWnahFeTn3FCVz9Gs8I+Crk7H+Q53nM26tjMEQ
gmz5layprm/Sj0b347X/oSA7nUwUqPW06Q/bPEnMXxwWxgDvyA5kf2+DqdxU5taV
uHFQGHeHSp1ccA8xBqDCKmVVt8U0uXZFcglkMllJkzJboy2w1xnMWULvXWBFAe5W
AlpycPQIIMII85h2iDrAAspdEu3hPo8OWxIE/T2+HoUa2F+q5E8Gtl/u8SnJ3p/E
zzYBY13YGQ6JUNqhKJCXfYoVXbfpBNYPb18gE0MjZYu3+hWtsrEM6immNoTZkJHF
v6C474oW9tc9FcUszK1pbSieQcPXHCkGNJICiS+EW4qvsAArAOTJ3BtiHQX2W4bz
IInuKWR/b7o7TBf4bTWZCEEP8nwvzuDuGUmfxod8KSizR/VROPeah9q1lacD+mI0
z8J0VTsqqg+1hGP6dFPiAsTl9yDrH46LAeN3QpYMVsv3kKFq+lUobHo4yXKAZeAo
VqmjYU0hq/rQmw2j4ZyJEExJmQxVh466eSzaGunnQWZ7IGg9quk2VfMGPqLlD5VK
BlYmPS6kdiLk1Eq6PqLoqq50Cr6etgdh8B0AmmVHXcOPKmrTGPW4u2N5clDGCtKH
j8aWqjIzDrRYPsp8PWQyUWsXV783fTMq4QXaZeT9brXJLLYTKUDxe2LlSJYxY04Q
wfn1iWbcB8LLhD1axd9P1Na3jezY57Z63XDnD7iE0JKCsV9l9Wv5z9hqbnxo1nv8
y/q9o8zI50h2NDXxSX6Y8Bh/f0vD5pTorEBQObTfnK7jKwBDPD90CX+twN5civHD
dAPo0e/EFLJnrNMa3rcmObSYlWsPOrYFAJm77dd10hU6Qyyg7EiK1pExfI1b9LOo
a/feyfvSFqmnrCKCBtcuplVbfXYqt+aXaRhvFCcUMv5tG3cq3fkPawxkklzUFEob
stEABi8fTVXa5Q3HFliLiyj/5yDZOWIuodbkjZHEF39u3Gs8xT7oz0o2BLzat8lZ
zAn5TZTUfM3gNiecbMduOHkbDOMoWw3SNW21VqCEsHz+hgo4BPLHbEHMegU1fPVz
sNzt8YWAM3H2a/GPUuRD0lhKD0d0KN0/cmQFvRNe75LB0FBN9EKg/ViA/lSlkvfw
/mVLu/pEDjecC5I8D+rAttdpY5CDNDz3nzUTes3IuJNUe528oIRdxYMTmmti3Ifi
pJQT5heYwgp2/7RjluOl5Pr2bF0R8zzfwJVeAcbXdU0CqYI6JeGcdPXOnZf08F1x
1KAPTr7epsuiCRDQ9zsBiXuzeFcO5KAs3pTuk2a1uYfPSt5xkkW9Qbp55CfU+VjL
HE09Q+MtPg9BFWQKJTWnXEZcY0poqn7KWG4Jg114Lw1JB9PUZ7F1VAP8iFOjjPFm
U6FsQAo58Swj486yD5Myv63tcH2zQP596BdoWLskNAgeDA/RGT1VrLDC7tcGhx5K
g5P1Z4LLic+R6d22P54mFRVqoGrh6jTA+RZNm2L7rSOprDj7WlazAiei+MpJ0wTc
vMNvZ8fRCj2R1aRcVDaw60FoHyrofJtbW9+X2Zkac9DyByRhX/gxoiv0b65ym26E
DeLMHubmfjmsVzvdBgS2Ip40w6FlDWQdIqGgrmwG+XSy1mUdfnnzWETlL6NXGKxy
ggpH2s8Re4mlHkchRLIcP6ZrHD/VzwJRrFRZ3Sbep5lJ6bAqMzDL4yF2Z6k+RoHx
0PZdDrfDiv5rFAkIkyAlgpkihyV8gC3E09D9GIkMSbaZora7VOa5+we+K9U3v97j
H9p71QCHToOWLikg1igzbwoPYY3buQNSagfKyfRu9PZgg7NBbX/LTEvPyjkeF0BJ
uPposglDngg9xE93WxDjPfOjx2FQ5vgF57ErkJpHx+coR3iyYi9n9E9P/hwYXtKq
8wk54BzvfrY3wBsIwOEFcP1kj9Biq1u2/sEY6sD3/vAZujpfdd8IKXLWWfQ6Y5yu
5S9uO6F/ld9B8LWlj4hH8LIPjPKOD4RST1OgLeJ7iKLl8bnnhoQzNnNxqFM7T/El
WE5cyezoMJBUXkHphYfkVngeE4ouSjGG9XLGAZrrJjsEsKE/QFU0IwGIHXMGkn3I
C8m2evTZpF3qc1UBtke47+pJv6NsGieP/joWGOqUixHrs75iAOY/Dm/SHQ56sHWh
O0mGyuyAYtsjOb2LrgTJju6HMu8SlDanjAhLzYgRinhHnJby1ixwJWM+uQu1x3l/
ny/9Uz4PkfeT4AED3TjuKOmpDtEP1AuXmT68Qr903SG0mVg0y25eyJN4jUSuKLX4
1W8zmPKdRfPj9kW0yFHy/FJj4SpcW9qTcqhmIc8v881i3sPXfR1w7GeEQvTrqXTx
eMdBYNpK+QIwLQEpgcccJTpeI5kkPvME700ovSSCWWub+FRrcXRE40AbTLgHdDoD
4xzafYrDJghOerCzM1aBnKvyMDdgSGkzjVxtNRXZT2Yy359xUSPLCMI+jk38xFm4
1PjTgklGF5j05jyYY7bF3k/BcHjdTK+TTWVL0Jf0Sia+5CQx8RHnljlFlAVJdOTy
av7hx6RmPdPHNRSRo2uIGiWY9mmcmtpFC8LzJ9z65faN6uoGotbD7VSdZ59IHd7R
d8orNQlzZevALEKkqbCPsTuLKkECklqZTha2BLH3LQGihKJThEPFw42hQMVznBZS
nQZY7qMa7SFyKvrp760DAWSX1Vfs1c9HyEJNwIs0B9c1tPWW7dBiOcUj98a9Fx1S
DeLO4NwM4mIE9WJGHJnfI7J9vdlRnhstBwR+7VoHFJPBYXQ2zgNrB+gAYG4j0beo
IKSjVkKl+yes32WUL8bMAD86puyqDn4o0taYdWcgDSMOCvZfLWoMh0x67tvADTe8
/Trp5Ou7LaTRyfZtjTOFed1vaR6HGyJI42KXVLNMwrzxzdvfbYVWZE1tdno1NaWz
+SDHp65baGLyeV0GuJQDpDqToxaMjDBoLoDKDCxmaLoPeAqWHsaylNSYQcfTsuFQ
PkSI1IzlCttb0SGnUJp4Z4v9wAe0b4vwFpv46cBjWEwFpl79a0ZJj9yxGjxNxG7U
V+1oThg09YPa0A+3/cM8E/4B9NPfC78QbMoMw8duE81kKHC2coEvBE66PDOfo5R0
clfQI5Cps+z2edV9Ek4ENzM9VwPr6OW/HDBzaXJGpeiKbl3WALlaatycvjBbX6vP
jEowZCA0HHUIxqu93gLCSkF8J19daCk8Z76Ul3nE59OlfTgc74akpShTQdcWZOFc
GHRtI1Q4WE/UnE7Wi19FRxTwx4vsNbcGxd1l5j8euGn1P/YjbQO2Zd34d8rUUvj5
KpVYAwiJ46nTY5eI7PUYrTK76ap/g3loe8rE+wC9g4jtwHCTVK8HkyWSs7F8c3jg
OnOTUDpEP2zTE8IwvYbHTMOJGZ5V7OcjpOnfOROkSyYo6loMsTRRBQXC/5Rrxw/F
xgaCc9SAjbG+A9jTz4xsON6a9kFtLV77tYGNnuyfsOKga77SyX1eXeocAInnqgRE
wzXuI9pQFAGNGOVhjFD/Cb8QslFe4UMJrQarADrSHOHVU/lC+spsTFveT7hEkQ1m
jgmYyYhS00ax8dAhIkPvVHUXQhwo7hAtE7vzCwivn2pVwiCT0OnT3rvfNSyKWKPT
mZgg688zWILNLk+Sa5k7ycOw2f9ERyiXHVJM1qQ9jyBj5TDBRABHwMcmkDO7z31n
brZXiI7SvcrXw7ViuwY0epNXBYUwN0FMqzQLSMpKKv0LixIrpqeqF6dzeq7XtLeQ
62HY3Yw4sPVhfxfHoDafoAwC/z99Rj2R3SaBAJZYoSIXwPTTnlib0x20JP9HSyVj
K9LOmFNfZsHbwDbL03VcC0Rhf7DpqB/PNP9p3s8eMtzubbnn2gwjx5s1yzSO0Ywi
mQs3T4RWXOzL+tm0rHKWp1Zy7IcmTwQ9oaMzt5X7mW46KYZxi7mAwSSKicH57IIB
NgVtAFoZZl2UpYEtmYRz7QGpwun2aBkacSW/JcbrcDKOQgDnPFfgfrQcEYCVnReF
uNK5BwBL7FUxDRyTGkFBs2CEsjzKCteKhaEilx+9lMsrWfzPRcIriigIa8IXRdaZ
O36SSOWZ6zRoNWXxYzS3kX/1hVVP9FdLf3lIABwTs+kXKXUkx3M7sw5a02RwiFc5
1opq5eFMrsjCt7hi4WN2V2Xi5LJKQZ/RV1nRO6Yfjx9ozRg4Ckw1G3CME38izSki
tuFFDvHEiGMlOYpGKns8EA3awiXoGlZ603UpeWafr5VnWYYHukQMNW2Eub23N5AY
kqUFD8xmfi45pGklDj0czzUYmF0rDFc9fIZiVLtVedsYMRCdky6w7mKcjO7aRCDm
eQKmRP3Kurrmxkd+wx55F/Vsp9pMNr/pI3H/LkE8WMx1u8VAEpWRpNcuIYIfjR9U
8Fod2oAlzdp47hCNobTWRu+lFgqPuQyxMx9nUyfsPyIMnLsD7rR5fAs5+Tj7GZ9c
6D5sZses0c3icWrHXg9Qqs8hfJ9lFQRmXHVNpIndCzFXtKH4afrkTEPHOJ8BS9zl
QgdB6AUZhwzuFZJpQ5XffTyON+X20qPkWeft3Cb1QGQbo9q4cWTzXxMY4oZeqjOr
da1A9sqowkUfcmJTrXeO/VKwo0S41BhMdSC98NKR4GHkcujUlb3kNXlS99LbiQkp
6gnBKIt6T8kFJE0ZV7FDls7WcAhPhxpsvqIQLnCFaC8vkciA0ULd35/wd19g+eKt
cN+I10J5hW1/zVypTYx2RGwlaCtnJNOypyw4ikjzltWiJpZ5S8g1i+GIGJxYcXon
AEDU2steJ8N99WnAPjTtijpbGj6VJ/PRz85CQuBy+MSoKPaJvm3ZaIJzWexr1bN2
5ntFUitZfAtXawFOAr6K36h10M6uwSV8622jA3Pcf3yfxy64Gs2X+ZGUPGBHojG7
YffeMauSAMUIxrNGvseNxpE3YxsjuMYCaifOFII8ahf6f8YHtsfIzknLjdLQoGJ3
/BWh2+tlrq+QhuSGxgbPuGkhz44TVeD2G3oxNpt8S+pPo2XPJ3eO4Tq7st4ovOQv
DSGEihc6UB16nHUkyfKcA07OtCbTz/5MIOicF9+QXzFmPGtVIMcuvOaBcGbyPURP
EHYjEKONLSfcomJkVB8tSw5zNq3wbE1RzIjfgo968Y2W58asTVEIcZctD0tYRo9V
vvtQhNuQzKeYmt8zdG96uqgc7gLTVmjPfPfBa/58Ul/ExGDTLwkWM8FsZ1GnQ4zA
EQ/asxWepkzNXUnoXWQ4fRUTX5Jdtw8JayWHnM4GzPiIVXNueVZniEQ1adU5cUoN
WbpIVsZrjw4euOkktFVcH3fNPIlTIQWgkRWjWc609mLiX4cohEX/wvoxGrWvTdcO
0IH4nrcQgdyjp63k3lzG13AnPT+OiE0x/ryeOFLX1oIWLI+/B0iOQq1PtFQP34fK
MtQZT8JpCqEwbqVKG/vhfV4kyxopYMdeub3cxW80m9t+lULBYdQI9U4LqG7QYkND
vmYtr+KvKkpB1xetuJJBn/0jFO2pnW2dpwh2uR0eonC4JVgQ3YBpukG/vjs3U6wO
7u7KQzYpWJPM9WAowwhN3WpHb0QbDJWqiowmcDjaKnLaEkvewbODz+KSQBLkdh1m
oTve6sUhkZaXrXlZYlpm3ZTBRtg02SgO3q6A0KKRXaHD55uorgubpHYcVa+uRQdM
8HTD2T3CTnJ7BqyVdzrkuKaCqEAy6E1gOxhrJ+AL96/eMdozo+tVKg8sfe1rt9Dn
EHTSsTu+2z9fiGUD/xpN9g7t9h70wi+7L+5GnH8QjD5YdTw56SZpjRJiMbCM08Y9
J4ZUNBjZwPOwjcyvWfTU8OhYq7VE8GoF9TBliblU2vAIyLzQGjYjpwWCCuW/yXv/
h+f5bDpPviMfEf2iD6aEkKUdap2klK4UBiMTb6zh8O7RuV3Q/F1YDWTQqN9rOSpy
JeL5EPliGAwziHJjifIRozmWZ+IYqUlyZ7xNrgRcvWYtW/Vqg7CLhvqcoNX21djC
OEP8qtdOme3dF6kasziDV6J572XI34HB/QUKna9j4sKzgo4gMqk4deHD+oOY2oir
Cx2cunE5CESvqWRVcp9noacccZHIoy2cp14lThe+SYoVA8CVczuhITWvxNjok0sk
KsL/gXbpQUfolxyJij13Fb1P4jaahVtO6D0HzpIimMxbXDZOAr8aLMabX8OCtoj5
5mDQOef9JxG/1jK0+rUaA+NZoNxbx8q06sUh8qPQCaTyXBTKBL3W4ZB9mR87u9zY
gVre5QCE9FkzQELr17goW/G8lF7wPTgBWiqJ+KV++eTzITBKmC1NIP+nqkmjqNoT
lMa7ZkUlc8wfraNB/7MB8qTV8n8jIixhuiZQJZHLGXFl3dkOKmcVuwlJ8Ql5WX56
sJjCgDUJH+aHo+3/6rugc7CU/xekxOdhvo9SMhvZJmfQiQoiw2no2ilcu5O5MHR8
sgW93a5X1l+6prPR9GAXphBkZdROFNypiiXVchQQ5V3PnDAcF4/urWDbNPZFr7EJ
oTl7TGxqE2w2igtqoO/YMLUqwTPDIuuePkBNznu44QfPOeF3TVczpdAXu+luJH97
Kg7rX1/nPMEtLZPB/FcVlv3KzCjlD438VRBzJi7F7lfTdfwvvj3nymjYn+3FcBAY
fifqLoK9LHqtXsEbwYvold5/Ew027pNNWfJSuaMOasv80C0Q9bfrxnHR/hiadfu0
Yp45Y7tuNxDiW5oSpcJ8S5gMzRKrpWmi4/sCMH9dnby8HqvZ633uaj81l53WJRai
nYLvS1abbi8byzKVLuU98EswNVKnf2Y3il8VA4E0+n3IWm3UU+0C8BhQNAirw7Hb
n0sRX7kj+2cztQQv84yqcgqtdehtUj+OwG9Vg4g2M8zyBKa3e/EeJCg0UgDNOUjb
rocV5raIS7KV8o8ouYrJSUe4fb+OtQtrY5J/xmZ/yQSrbgfwOZOXPdl2+Zr1dARJ
r+o9/MXtUDfTFkLCIIG7HnSjy1u4SnQVLU6UheqhB7tnYhyI4Z2CksAmkd7MKes3
4bsTrnZhu/TMo3JyGZGpCEuaqROn9/5CRsZU5Gx41OJBu0inJOCo1g6hXVnOQlml
WyLXr5aGrg840s23Zn0vn3xTuhpl1qH07RlTtXvdln3Nj7N4euKO43t3NGYf3oXU
YGQ3TOXBBxwiSyVjXPa7AXhtcJVMXo/blE3+NgeqxiPwJ6LNLS70wEyjyU/gfOig
fbTcP3o+Z1EIGSW4lnC+qFQr+cgGmWZwZMPLPI/AzwCHvRXikXx6XcPDvlMTmV43
aML612+itkGkG3LM7koaUG0GH+cXGh1ST4DwsloXsd5AjpR65bp3uczgCygNW4TH
4QoDwuMJYVTLWsxUImFl81tVYt42VCO0g2mD5fqlnFaK3E/QdxUUmeqJXYsn55Yt
WHlU9dMq7aXma4gcQsiiYL+vlbj8aAzhnaPlsezoDLVFAHRHxTZiVtcSs/PP+jzI
yPQRX2aEdQer+IxwXVkY0sZ99EdcVXYJnpsodHP2TzhXiXDkBBDIkacJHXjoyPe+
mspPjRp0Aced/14KOKg69tjCH/j4byT2I5COVFVR4CNV6MIFmQqwd2n6zLop6A9y
UtyxJ17ko3dS8xCSlolai33JKA2EmGJ5JCkQJY89X8NxN72loknqOgG1EhEm7Qi2
dRr528yc6yzMBtpEfBmHKz6Vrrsg4QQsb9dd6QWMdH4gFEBP2ic/BEHGTnh3sZ7X
dI57S8vhrzi1dpuVvRau6GoEGwpFlrfY6D+e3dvlIyA2WMYll5cqIvVa8E/xLVZq
P6+9LYWNK6b2z//ycQCRYdTbv1RAUmSAE0dBF6C3bCosR+t8Lw+Fs0p0AbHx3nww
1w+mmYL0pr1M0Fv3aLKN4PC9+0uWAtxuoesI7VLkefQ4X31vNFRTwz9hWsYhsNup
8PJPmRzVcc79YONDvTr5sTyXGIoPvCKSGck9SsjtyEjgCnllH+bPtkcDb76M8gQM
xuKymlNUFs+gTWA2wnti5cEzJ7kEz6gp/akxrJOXrNuRZDRR+vCSOPjf3fFxvwPy
+lUQTs5ZOHSm7ixCjBkaDyaUfUdmD7ee9PUbv/MF+Q7mKHWAWrTbpHM2Hs/T5Z2B
hJQdejm8iwotNbht5Yus1s5YCZjp/2EB7HBQpiCKUi6AhMulKOriv7ts8z76Z9zO
JH0kcZa+zW97X7GWLRtmZseMsEfqia+T/j2eEq0ZY0QMJgcwDKRea+goXIOhTTb/
2wgay+D21un4gkePxwBw2ldlwaF0cS+4G4ojmbBKxKyKl5B/UEUUTXMBRt4ID3nB
Oy73ukTJw6P77MdjpKKv5v7wIhcCgSbHSlnZvjU8OBwbHdkcUrgoVlfBTC2Gcrn3
7VzYXeGQdEkDnmjg5ALMTU25QmFIYp6vjEjux+U+JcyMmOlAuxVMjI0XquKROTXM
hraj/oQYd7pEGJtslADDi0WUNG0Js/g6MoBy+IBh/26wb62R149c5YGLG686PsYN
qnmgvgT5L5X8VvdgMnN4mxv4+a4EkvPpVPcSQ9PUQ85q5kQkxQ9qMMhPExfFqTZQ
hNxNecLiU3ZqoNsavRa/opVE4xFfOh7iazddVGir4qZg9wbrJyqHwQ/kWq8qzVov
ZQVSB42aQveZmOqvdOan4YZtYJEUlxi1wWXNPtd+rg9lSgaluueSTXs6zD5/ymUp
qA+0sPq7jvHuxeP51gHCYbmwSOA+u9SsV7djPXyn8cvTZmsy1hayPPhJBnwPdCVf
VmS9t/vJgahH+N/nHeCSUFXhsBui0gQu2t+lDJA0+UF5JaH3RNxlO5j4srcMS/t3
8aZNJ3hnf1b3YQZRYFP+Q0lfJK57GsSFKYLAtHhHDq5lgCC8gzoU3V6s9Jl/MNmQ
HHUl3wadF4ji5LoCJe+MWq0V1JI9tk1F626g/jaM0uRE/CAZ0dBnxwee5FctfcxE
wrvFxmpwVegKcZZ6TDF7DD2tTThVckZatY4w2ZctNRB/Vachqz6PayqVqujj0b+y
/VFSSsxNKUGXW2mswYBpHzuEJ1YODD7cvqFmnZOgjQr+/MP4ousnsk3PvQjHpgIP
xMAq7kwuqFlRB47vPp0EI7md8i65NMhASLw5R1S+ZuH12Vk+MM7NTD1ZYVgHnqbH
hjSeiwQkcWbcnt1fEtubUFNdwk7Ud0+TiveVAHLWe7MMFx/6cfyouSLlVbRTYFJS
aW9+WfVi/udwaIaKVM3ieuH8dJIoxuTZLDEBmF1xNIL2ZgqNIITcyhQopt+YTdoj
MJwe9A130mo542lghiuVgyo5PToYUNZpa4BgTu5kkUIZHvHtMrv5olClPXIbSXjw
5ly/n+LSCsjbQkglFCrIex6hRgi6U9uL4wN1Aa5zB+PpwT2fo7od5A6NR4ZEYlez
G09D9CnSkXneoEonseOhKdK2iZnwqF098rw4DC0v5j7/rhwCLb7wa1BZsLEleVzi
kKcOs5TtUkgkXOcvHW9cRuLQ7kludQZQkmrZnAVPnNBWK+haaSzmC1zCXPnH31Rr
4yaqc6/BkaABOsDEexKGppJa33EabG3SKHmmp4DYiAGioT3SQdTe42tgZ9cKAJbY
LR//DCynavpnKNeDWUCTL1MQaeDq0GEsNvWgYYgqS/QOEjW5kK/vbePkNJUfwAZ8
2Mbz7X5JoJ17U8LlahRsRv77/Uwdm1w5gS+U1ChjJKnfTS3QP/dBxV7Df+dlxh0N
ETYMPKdflqQTTQs0BhG5fmXvxLjDKkd5HAFUaUHBGja71nM2HQ7cRK8CipZpDKar
lBdiNp+7/tJBwBJRWqFe23MfSwt3FI4YdqnpN4Be9QdbiJH9B8orax0DWmDmrraw
twugGIjHUWpp8t4xPFowcN/I9PAp6gghZixbLJqwcQ0DUKfl3liUpBhw4hnxEkDD
q+2egl8HyTlEfBUTVskgygJjFqBgCkh/qMZIHsTfxyr+70mTecdvPQzzM3G/ApVY
AgyXt2lkpXLpKQ/0zWmrpoZOqu0JRIFq/V8sGQfqqsCiZ1SJ5+kfV73bMUrieWuu
yoKv+tp34xQQhMCs3mSfD6P5PB85JXfWL0xDCGfzRXvQGSssG+WwCMFRqugxB6me
hsjd3M8NTMBnpkSYrCnK8nyE4RqkRUiCRnuQqX6zboUT+R+9UiPPy8ZUGfNJo9bQ
T5EMlpWunwRJLUg8+YERC1hoEh/1XtxtofI/U2FTE/7uFwg8px3m65gia5YuWElI
drPhkqIzT/96brgta6CD/h0hAaPqZQS6s1pbr/JbmETSrBNTflPoSzixSBONMz1m
u2IaOOtIGVIqL5dz3A8TahmcBgY5p8CVJIN9P8FGZQr0/MHno7nuRlHvsgah9/jT
J4VzR37g+J3qWepyeelKqbm1ESQWmroEx2rYGZNSKM8dnD+W2JsbCB/TvXQWqhyZ
W5cpc3VkCGHHgREwIXbp/WJfrAFQJLDUgYyT1DlUkv5tGTuxlcCovWZAIMYqRri/
8GO9GykIFcDndkozXMdSXRgkpx+i46GU0c+GNH07dV9bdH880E9dtaUHFgFFC0Es
TLNPVMYmzk7quSU8UHXk6CH8kLPoET2CQ7LNKimC+FKUL9MQwWegV99FPWn5ew3x
o/xn95wxlQbj116M2/UqGi1Mhy2h670bZu/Wmh848VQoZOZ2a9At5mMOma2j/N0l
6/BI0kdnINWC6Hq8g1N4645/bVkfKXMYmPTHKtM0OQ2z9ljMAGjPUDvWRxRH3DPN
SXzDVSTUkN+WmWj5qC/MEu0EdWf/fSxUTf8apTxdk+ZxW2brvu30XDHWj7l2TWf8
2PB/h7d6gN7KkQin1RSZIhQpKcBnQ0+cA0J1T32qKQCjLfYxIXZx5rTlrd4PnH2W
tOCM7073huqabRyBA2BE12Jh8ddX4/9KNvg7EtEIM5uNMbu38VJ3p8j2M+H+7KgK
3xzPapR/RqQPv768R2ar3q12PMNDHf6tG0S7cIqVmcHaRtalTUqRrKpZS813aKsi
f1nO7GlTtpRmhIb4lKyoD7qOsu1+40Lqk6r8P12BgKoImxV0PoIlsWWdg+v3BKpw
KiysOtym1jt+Mv1VUjZt+I4Cx319KLlxIbg8cQEeCVI4JHGXu9vlUf+cdR+Fe6Gp
Wz9+vObekDw+HELoy4inUwPLRHOUSGyyA7hH50/HmT+eTas1cQM/P69jeSbw7KWG
mcdd3r/McHicfC7ugluUIh/rDYVujFYeVRsbJlqsfnMA+i78jVwxnkZj+pjs/e0J
tPipIiAduFQKBel27voRVfPbKD2ClPmU/7DMeSzqiQdYZrg3xOJjMXh9BVbVq5DE
IHqBpmGubEu2dRnhyTOUxQQDMuMVvToBB8GSnKOka1EMIdFEqdrL+Zr8bwftPv3G
Z4QE/Bgy3Bla68eWpWiprIvVVXEeQqm7UibasuMYcyPjnxTsiqIwwHiLg7JRXOPe
HLv4Ue6+8l/V+NeACO2+yT98QOeVofdGDHAGyenUr39Vfopk/1FkFBOIl76yBdmf
WvPX/O5jd+rr/I1e6N7NDDcTJnp+enci0kH0bMMyHDX2FlcULqCrRkkrEa3l/T8F
L/Qn1sEIEq0IFCdJpUkdTEnv6zRBGZwA3+S11FyqyD3UIy5hFquirp+d4SqaSfMp
1JbBPkjTiuih32xd6VH9EHoWqGFUdSNufl0MKnAj4DKy/vHyeTNBDxTS+IkI8yDJ
78XNNGXhQn7kHtiHhCfFmSs09JgYiirpu9BMIe7yMRFbTVb7uClCQCU9d8CzMXfa
p/KYwlQL4EjCEqzOWpHcyvWLQ0SWKIVdmnBqTNWkLrSjTMHP3HAUNkLGlCccUhop
5cgqgWJgnxmwmKG+/VzejH6UhKUjl6Kk4aZ9NXAamWkV7K2XcAY0R3a53YI8aAy7
HR52B5M/z3FkJPyXz2pcC7jFdHOA+li8iKlQZGrWLyZkNNAMvq4GpqM1Lpw97L1p
/Fp5k5W4Gt+2gtTdkWbCv5UndCDLQXSDASJ192tINj85y7s3BQd4R6gIp6D2nx1p
m/BRhlMGzjE75nIejxTasJmRLfkDnef+JlPsfz7sNtxRKMHYC/yvy8sbjhqmtS8X
BBfUZSAlNrcR9fWQiRz5JS4JZiHMbdwy2I1P/d92ndMP+W3kMidIQhHcP0aCWLK8
dgy+Z6gOwU3nnaKO2wi+DpnuxY6XWNpttuE4fJ7AoQYkfzdJgm+SxLPjGtbESHoO
eLOZA/wzsdCbH3crgUtpSBn+oxzMmTQGIaMR0NNDMHr7inbPXOVIcgQ2HLIRcKMd
3skHYJsLm6vlrnXQJi7XyU9YbEKmc0ESkG14vTQNV74NzM6H5qn3OylVKt7m081x
PxhV/J+DL4um/S6zApVpGDI4Amwcn4y8Ppc9hlmevgAPP27H/PaGMfANar4uKnaY
y27PM3n/IpCb9cf+oB7DyRbpMQOS3EEyhwsZoUIgkP/9i3P6qvb+C5EmjxRy/+vh
/EA1KPSw/wF4NkUEagQf19umukMfvw/MaAUpsXbG6DadnvjBwCeKy4nOjPrrF82e
GBDTHfa5+LtrBBq02ruZNyfHHtsYWk+fdB8CozeZcgqKeouQW/akmyqyMB8/MlMi
Iml9Lvj5e+4WdVXo1pKOEivTIPpwvYQlVKckpilBUdiOlSjvvOuLu4TNargxBOZ0
gCUO89R73CisJSnph7KVoTV5oW5ILTkun77ei9fIlXShkurUL1C85K/WEol2osp4
WQg60AUvznuNDRIm0qN1DibkWPAJqVTbBC9UJXr65X3ySstQohWg3gVF0AX04u+/
t3WVshUFSKUw0o8KAnkmCaLwgYHs/klBGMpE82YcHuVx1u0pqe3SlCYUYcKBj32q
vVUZoCTXkF119tAR9TssRXVxKe3h5mP9LEB6sT/lhafUdVvc5TztrNwIPlOeuz/w
P8y+EztrMjms0MOCCkwBHhjPAVfCjI0EZ1XXkLonKIxyekuU7TiP5S3XFnxeSrEk
IAFxnDN84UoEpO758ZEXWWFZ5Knq1TfKjMCWZAx8VhtjLWrbFMKtyh9nP3z/iV9I
RYoP2xlV1WhTc7pjHH20UZVyFWUR/hJp0BTkh3Awa18bcvZDCN/3zGGbNi3c7Sn4
3HK6qp2HOSwus9sqUFXZjB/jjQdflwTSYbepnEaE1+cRXCFz7PUd3Qp9kGWB1+vB
gQjW/FG6RvFsZ5hD8CAm23WUlw7yzsTeriYDC5gBP8By0xgMZ+tjuBIDDFvEFP5N
F8mCwzDslQKanGGBT9aErqIpHwb7zFuvU2VmOqVO2vTAoyw50CuhfQgY7axHKvQB
HAS2IkD/jBXWsXP2wkY3FIlqlDuzPyeelFqpa+B/FN3bN9qyuAsTfwuuGB4lWSPG
2fwfYrXxdfpieo0Ei4qHymz2vWZyB2qiHBDIUbG6sS9AxXNkiAUyOYYi47PhyTpd
mtHnNt2mmWIgf5BZOuymJYNvARXU3b8TK2OjFo0bm/Tc2bHNRekaW0TmhtXLMmYI
x3tbH1vIPS8pO3WK7nUW3NUDXUzgKVJs0ge2jFet2ux/QI/GpAKpjwBqKJAp/7ya
CA1tDbiGPC5Auceh80YvqQdrEfJ2iKUyXeojyhoa7iWs/diHFmkcv3xBEdl6GQI3
8cDHEGZYiWNUsF/c1s+BAebFsfejm2/XR5WtDb+UsQBiDOZHiHHggZIEFQf2TJiX
BBGHtEPb3Vja/sK9/OQWQW83cNqN1RavioLuSkS2nf7MXUHnCBiujLNM7+1U2An5
nVxpESSdpfzeyPARYoUoe4eCUFZ+euJJU1MMIH3ilkparzJG8DhjYwaxS+ZVQ6Q2
11CTU4c9R3RiZaJyGk6c2Pq76RDJ89fyAbCvaTrNg2PvgM0AzrqLCrVhHf9A4DCY
B9c7KEMMI0bOEoZY9DqsTy6tZhwj84yo6CGghgb5HFuyy9m//7CpAU6awOC/GD4B
1lHIjP+vQd2tr1y8m5FcGW7ll5+N7GJ8ync3Dv+Qdz7yjVH2hNH6ryVGcril49U3
P1mSPTLXXVfy7f7XHYKAfXm8xKjRHW9pU6VpbKfLC7r2Dr0l7294LvgueLCNnVwb
vnMU9xHQT912L6Ifa+bq660TyChHOmdFj/e10DCwmAYjf68+EYd0QkDRxje1VNIM
TlWQ1QLqs10dgOBhxL9qKqnuMevb9UXVVDz9lY2ZSUSG60ObQz5kKVoLOFKIKvTL
w0k+bpST3ukdcSBqbtpw3O9R6JRTuOaqJMQYhlbqAoINPv3YmV+ogCQWIFsWxh+H
rKCITfnnzkI+c72m5winL0zQkYoczksWM1WF2XPYxxZG7U708GS1Qrx61QY9XToO
+CKvQhSzFGnXDua+kW1UxXrC9LN9ycUbiFH1zrXyOHikSap08cogakkdoAb0o15G
KvSE2i69KBdKVykcdma6R5mNpu9oPheBIDJ/WK/3tLgOBnxWrDgAAwtCbvyPOKPs
hiqIm+z884LPiP/knWlf+p/B76ofHNCjGlNwxDIVX3AFrFDhP1yWmw0gx9vGsVpM
vzYvQwVfYzbPXprqtSRl2Pxel1fVg+5N3vuynfwU+c9TPn9DyZBkkDtEbQDI7pUW
g/Dk6Fi+IVGCZyLqoveeJMQrwiIRFRVgxMJG6H3PGEzVhY4zKz5WEWb0Z1hPkaRI
/6KPFx8BTz1al58yEGgzmmJPCKwmRc8RRdCzWOhcVRLHEHaI8iZ+fiQXZe8CdMTi
hzXhrIxNqI7wbK7e1slNtoNo7cViSuCa7Uz9ftcDKslNy6TgdgqKvuiJidVOjO+P
U5hEEBdYnqGGK/uURKaujzA5mxvOkWVzFEUIygtr4PGMNskCTG0HH3Ljy+9YocLT
ws7n8uaXqDBW9TLUjthX00bKVyKDYPVC6R60hQitmN2h6uI0Rtn2Kuj+tsYgH9IQ
N/ErhPilzzWBzQ5f4Un7h6VaPe+s9EkzKD2Mzqfz5X1TkGnfhMLbiC9g+MSfv34j
6NokwDztfZdH3dRSrlWsrgx7AEM38moteBtM3nnq2QpGoS/DwkpOuowOa26HfxEu
1Snetv+r7xJXmop2wH7cFTCiKPA1yqBsOPi6KUeI9VpOBkHOybRlLRPI2Vv3Br9g
rZU4nFO7ZNX+cuQ+jBnkDXbObijWSboLUmGFvEnkaAAzbcgZYm99F5rEPmPzVce4
HcROFV08QNmfKHH30W00ciMsZEUq7OPFVwogpFyQe0+sRl93XUe9wFMI0YUe89M3
xrlWK6LpTuRzXVEPy7ZeYD8tL2qHEPi1JSj/aDMoST0HDFFl6krubo2PZY5fu1bD
gQDyV9R08e0/81eZHTcDvIhum7KlsgO7ErH8CYnKTGzpjOr944QhzviyvYThhMpi
xh4kgk1hxesO8ihGB/92AWoqX2OmL6Z0zk0FQ0LO9Zwj7F8wLcuqtsUeg9uKG/fD
Q6uWac4E9kUvGdvN0yi/R6AxgQIEaUpDPyCM+IVpDF5KFcuctaUuukTXCnBWqiIR
I/Lm0MMlmXft1Ct3DzZd3bNOyqYKtjth8XZZm5OP9RxMoLix7lxMyZklOrGo4A5V
JakrPT5H4yZTDs18draR9SHKlgJ7TIwa7ub045rekhP5mUeZh2kpq6JgeSVn/6Jd
da1FrsMpxDCVqyiJ2IRThrHss5IkyTW9h45QpJKcACSSC7SIH1VX2rKOkRrdq3mR
+uq6J4qu23V7q6u4zPKjVkVQ9nthdGa4wuIItXY9yuSXCCp3/hc6VQjk9e9xlJ/5
/3Alm97gIszqGgWOb3vrRatlnJh9YOTmBYU61pphO+uJejMTCz0Fa3HbFZp1Z/61
0e9SJsvkxdmyjQOlswazsNC2IQUTcp+CQbxj2JOQM5DSz6x/tCrWa/DUhzNdXZuc
ePNm3G7JCk8T6/7iHTOfOUK8MAHcHDJxZdyMCWXz/AfMbe6/nm2+cNj6XwpFBN33
PYG6tj5JnywQeDEM4i9/nJZmFGxh4IrkB94kx9dYud1bOMUoJ8RRvs2UdFysMYuK
a6495g/d+yWOMWl6QlsWLM9twnXorhcErVPkUv0KAEDYibhxgrmCRB2Tknqlix4k
8rzth2niT4J07jaACUTrr2rbX8yc4hR0qORy5sGaswS+V171OwJFHVbvLc+Xjduj
UwKQcU9sEBabZKCACjlpCrCoZR2teq9hdSRPK+2ovSzJ+qOUeAVt4Lg4jdGDDwZI
ok4To8wA6tB9fBFI4qMmLwYUJfMZkHeK1nk4fiQDTLEEoOHqGiYNkUsIy8DMV7zB
qOiM460Bh+Ik4ULuyYl6UhShF7MoBmdbNhhU9Hm97euwRHa4TgcxYZQIQ7JSTFUU
CY/fEZcDcHyBUUmcjpITakZD2Y8/59pNUpu7ivLHV7UAIJgUegKIqxYFLD9jlTv8
Slx1zkoEmyTl+n3+4pGocFkLP7yO9UCfUqBpGtf5aMS7f9Rp7tPQLaDCMDni+c7k
dj+Cq8BKm7rDGuo05wO3czPCjcwlft9WAK9scz0ku9naS9fliUYz6w3s3n0WRnTr
m3jAFWNwhwITg4MJ7wPc1fAryUTkc9EpBC9Nh7LRsl7vYXB2Xa6fMe0c/fDRjJjM
e4++q5EXuJK1uMGVllazk7vXrbniyeEVF0Ke0IuxL3OxA2H9EUTVs8jljkZ/CMR7
09q/iRb57I8aQ25+kAAGSrBGJiYgL3ctLx9J0rvqH3MaOA76dJ9qVkuvkU/JbCwq
ovBWHb+I7SjfKytwpTdJdKp/fiSA4PcF/e6WVn36uN3kSGuAuFsElzPAjnxPM08Q
d9+767jtv1M42ihoMBSaVVFAfaR66Oc8fFGSb6Ax7d05oQR6rBA2h++dvtXyOhha
VFCkxnJjaMfnzO/PNtlYUphv6jfRD6uoyi5dHmDRtqKlraF7ZYaBUylUNmSDiqzK
rqrtKLnmFWWb0lsun37ftPBPwkFyLWAZlYL3koVEQqkoONCLyyZHtk/epFOsQv8Z
rnUPcc2n31pDk5SSKU0sYblbwuhUEm2Yoc7gUb39ViCKDE+r7KCeHvxhZ6/s5xkN
FHGYfEdgSukLSgO76KUst0w3Ny8KgxywSmEmEgpZkBwSS97y4Plh9fzWwJtp3ih6
aT43v4kxLer8ro2veBx9E+n4bZuPtYXk4/hqFZbABryhiwp+O36PaRlRum8Gg7e1
VxDarkJnWg2BUCWRu8pQHIuw31EJIfypcHEOTGft2OtFwv4njOkoRWxjF4aLUU8z
2FnjWqw00X/kG6ZQEvRA9KLi23cqU7R4Cuyi2jKIpXnc0GqRiUOukNkG8B0EgebQ
HMrPe7p6HkWaP/i+Jnfl42c7JUweSl9Lo8iJfNDa1JkYbFZD55rIG/HahCRHoOHR
5YNvpc2BAEHhNZhhoiOWUVEIRFztw8k2x8wf4OYWbtbK5W2yySWWxjwJgWb3s7Va
FWYjIn1xD59xS9XmELmreY3riewF1xIpLSQYxPyUwunR4OI+yvaX1pfyNTMRrhp4
ODvvyEPwN+KTUVXv9g3762DE/i38o8Bxucg/yFrjis5vA4/2K/R8DmFpl8syHj62
C1rK5MUxFTbUFFt1PJpNZ9yngcYSUWokqZ9rWX5jrj19LjbensCsHyVA7b3Ngl9R
wZGZOI+jiaNsZlSsv5aucBQgKbvoEeEts4y8g+LKL2poQ2wnSq8SC/X3QunlviHN
mOrmVpfhZin2RiRMYdQ0YFPQeDvocn7MH4zEo9Co+oNMI59qAIsr3KMy7y0Ao+zd
zCYSR3j83iJz8opIXCKW6He66gk07Ckj7i4r4dT/VCwPwJPWQjG6l4MDSwlw9Kiu
vjZOY5c5ZRPosm5GeSU4kodsCDpztWz7t2GzC1/sqiMS+3wB62cDFWzFbhVEerDN
iJFU74sUsQQtLAZLESqKi/PxY7fJUU44hSqu/2VX1jqw06aBWo96ImERH6YXDbew
+DeRT9cF8k1xRJsGuHZTECJov4Ea7AafoYVAD4qEGfrmtvHl+rsyXHi9VMhuo6Uz
rh/LtFXt6OW+HW5cEoKgjHs0hUWmA0Cpd+2+t9A5IB2pthhwQ8ubHmhr4owT7t6h
2IdpBUCydEP5qRBUYzQgRls91LV3/3RzdAqKwrWOb5DSLHZ6zAGyQt4Y5s/Yaj4k
hOHHHf1X54o3jiFflkmg7OUq2+VOaZOwW9ZwjRI1nJ+2yaXW4pL0e4R37yl9zMW8
V2GiaKegTH7jG0NtdslbIqIgbrYPtsObDSCCdETVX3S68BnqVgXJXJGe2sLaEOVx
XfStErmxaeozReHaki8ning0aildE3+icPc+FHiV6vTh+7MkzwDs+i6Vs8Kx5Qj7
8xt5UianX8skT8ZfMls9Qoik1be2NTifqcSOud3wQKQfk9A8435SxBcXmFrKt1kw
03tEWI0VkBS5u5ELDhMkm7OiCpn4BwjNfWH5PadFDZ9965h7mMVpDIM5O3DtXL5F
GH8/WT4m3lh52l3vdj0c7Y+0p7vTfH5vCip5WI/s6ZPjFalyFB4HnvP7bBYlsXc+
Jm4G4khHC5mZLUeLnOmUk0/EiaPwDsL3YzB+25RfcM5cZfd4HGT44tDTUGuWn4SY
h+R+mem+y93IkTt+/OGfEMN+o7LwsbDuH8DjJfbc3r358Si+W63j46+hd37Gckbu
d3+9r2DdVt6nbLZIOZH2RpHyhxbyiudrJyRZWCod+8/CHZW5pkgIuZnBShuTT84x
U0L4SM+jObyh9J0fse/0ZkzHMctSqKwJ1YdwvUi2APR/D9SepGcMLZw9AkWraiIX
bZnNKBJlbsnKhmTUHFDisGDo1423h+db67AjlOHTTDIwMi/ZQ+UGSxYpQdjM6tnW
mOC2Xf3HbQUZ5qPMCf+Gv/Q8vRWiwRFbmlzCsMMK9ebeKwrtrd/d22kPkT0swXz1
BUzqU5g8z4W6fMrX3325z5yNHJveP5w1GwADZUIsw6bIuH2fP1oBWKaU5YL7h2n6
DdxJW2sRwia2RNd9j6wiNopyRF5jcYubs5jI8HfqRWy//x1rzXwUUbqJ1yVudjB/
1Y2OQj5XlkSpru1eGx1b4vpQdoPfEpXebqlXv/HdDLXIhnan5T1zmR8EFAxEIWqK
FyAxHFm49Wc6MZ3G+RmHWuDblTyzNcMoFTzI2OW4YcxnS1I68A6GtiNAKHpaN+o9
/POoDMeC91oYT4N1yYS9I/1hLHqwJOmWBuuNaCS+ePIYLJ1yi7e4qf7svvjk3JJz
qjJgICfCUmOlTsO53jynQ4oxiDYpLstwFAc6oqmKCw3kkJBSer8Zb/Ck0VSqtr8M
xII+wl/AltYfYXxK3pUzUVyBkybmHkMqpkOxet/shWQ57UXfCQ4HJ5hGVZ/cbJKJ
8bU8gDowA5jLtiCQ5W/4FlcJieOYlB72Zu2GmQczhtHqzPXOwSOnBtCYMf7/9Xou
l4CW/cYkeD/vSgxQu8DSRw5AyXBW44GFajM0nm3mLugFJRfQuA1+6LuBEPGlw64C
vanMezVbKSWzYRJ9GwDDdxNWbKhOIHTOfJeCBeBGiGVSzbWDuc6BzTeJxJoy1iUl
vB3uX9g30fqvKdmNgvQ2J1KuVGOw/Zj4rupUYVhyNAZ8RzkHOBawUCoLtI84LihM
hr1cUT6Tfje4ip2e3gOjCnp+gCatiSi+GrtEu+sLmLa6IPYElS8nWbwSBJ48IBwP
ic2UqzW0exNzs9JxGlpJYIuCSkOpb2cmzdsvfyaeHCXscDvXhF03MT4Jj26CuAsq
PDsD8ZILnwpAEgFm85bOuOSsgz2ZQq35c9DBZz39JrRJ+kMX15XfcsPh+BabnrN3
kkS9RC1P1KrYGgOavMAmWBM8mFPhrtF8yiDHE65Ax06flV8LbGKgd14dCRdmU5Bs
qAd9mXFffYX6vhn8eSFsYsrTYQGi1O7dLLutYgDsGNmOv0VPsofrHWsAdh8wdW/N
WAQgxn+UFEz5M6O6hu+4FZsR0zmygy65KLJJXpbE00IgdPvfCDuLzPnK99+KV36T
n8MWh5vZR3Pu/5tqfqW+nSGzmGRVryYNHSX07N8etYmHPWVhfpO4BuM9td2ehMwC
NJ2LGbHpNduqHZBfVP+TwHH8jIx4rOWWpkF/cUXIaf/1OrvYMs1KCjozy+DnOwNZ
N+hgac98QMEUsMHENnlwETY3UJ39JrAis/i+izMVw8lMr6HhLTbzC1GnhkeRnQBs
xE0c4dzXCHffv8vWSaWCanJrI8Ta2lDR4cF+vTwLtLZU1lu9UCJFoyRYAz5lyaYh
h9f5f8CVU1RJE/1Mo7yxhNmL7w1qYPM3NAdp6+V1vTfmCjb9y8yy+02Yr0ilhLTw
DGhCvS1Arw7xbtPXrh6RnqizAq7b76l7JjBeouEF7yOZeNwZuhHo7z5oVh7aQpPE
+cUQdxhJpF+AN7P/oHO1BiUMgT8xlpT+kLBb8J4qSFz2gROw1h7rBF005c25W9uV
AbkAXHvlgShYP3ckkD/6ba1q8DY1EtF96ZSOYwd2xxL4KMCrDOD2i0eF5UOqNaWT
94YzHW1tqGZzobdTNyLjBzKOi9/pX6QPFa901rpy3SKYCG3y4dJPQIJfwUZvWBOb
jW5X4GoA94F+yApzzwdxRA97Dsuyg7verQcSpuEUaL6QK2xAM2tICWVtIziQefqm
RtrVG7zT8NksahOf8rBm0TRMDcgK74LqwY4tJP3nbeiK90CfLoD6ac5iJs7UqMXp
n76cfcrK9C7fxfq6XbPw1SkdtoADoJBKhIo9BwbTHQi/hv4qBpYNjI4PcA7n+anS
jRSGBxiHcNlFovhNsci8IUADLXnjagw6NRm7giHZCdIamarO0gph9DLFHgYimj2Q
lPIc1rLS6+5oCcpUR9JtzaqM6eimSu5Ui1FFtchV5d5Qbn9j2sF5jKnqkNvoZ2B2
x05ndKQ2dI5uqek2iBzEhQjk6Lq+MUVOJf1Kd6CPRla+9dX/f84ckWYwybfhHKXv
bOFkaOUBD3IYt4nGaZam36YX8fH/p5E6e4abGMlwd0EswLTHc5b46E/78HyfldFx
Kyd2ibJk/ZuII4HL7ZCGFsaEiYeArl6cNLYcu8IPhqptvr2kTwoPFI/HmHM9RZtv
MoKdgZvJ9SgFtlWWPY3l/0M84drBoRCAbflrfffvOrWtcB1vYMqTDFm6ED/3TDxL
HaYHY1sfu0kKvWCjukk8gPDhU9Q6VwJ7YFcdPuhLrwJkQ3T/ytXrGFScG0DkRsoQ
Rgq/vS+jOtheV5UItfFQigDv9a91YTlh8Ck8/yORkO+mc4N+lWHgXzyE+wQjgfmh
maVuyoy4yryeRUhg4uMQrKbF3B37kQrU0MUyPJ+cYQLjp7SpaTdGoQU3ZlHAC/GL
7bYVox8Jj7ybxEfCR83C7wQ308GyRdIj453MUzbYd28kKd5eqWHgnrfLtG4D7QA2
pInSFn4CZGaPqMkrCZQ4psPkj3ATV9iECNqi0hqbmJHpXh0TXycTFgYETM1vY0xd
XFAqSR0V35NCCGXLEdRwtcbfA1FIdRUHRjp+bQRNBBw39b5vAYRwfy22AlVCfmGm
QZJ7sIoQ77yc0lNkZ0E2WUp+0S1KFCyBU2TSP/6fdH/EMQ4JAkntmXM9utdOcVxW
yC8VC0aaaV4q8CvUYWPOFw2833+ARuii18V5td45rkAugmOWa2HjcYi9xwJWf1ow
5mRpuXfXPkjJoLG8GV7kaVfy/9gKMhK4ElT0e9rHEEzg08FV6BKEkX89gwUPvRM+
fRLKuQFiuuxZxk4rxz4roSEnTpuxfWLee6JF9x6uV8gNkqj1SrvGZtUqhSgd4EHF
7uIT/gHV6gmsJ4nKsd+t3yHA2ICQ8U8G4EzLNKulryIyhb1khVLx6AhLZw4xhRKO
XNnw3CzLGnE2TvSw5ig44cpYgAczUfSJOlSSToaQBqfvVm+DmHckzTPI8n3eD/Wa
YDHMhcV1qe7DDrXsYNKRggWBqvVhIRgcX3UuxNwzVeJB2CSJpjaHMD/RogcbBqCH
aDLrlWpYTjyisO+kEkd2JRKjAoVFDdq4TrYurVteDW2N2sud19KixdNb0F6oT3OH
hYKpBEwxaEcfueYTJTplZPY/A6f9XOAAg81K9T+b/Z2LRuI2xmbi8NikzIoRMbMl
k46uIKQYMD2LWwWyQQTsFEKfD780lHo0e5l+EhdRd6q/Khk+5kVOtYkx5rrppJZq
hdKdLrNxg8ZgJSUkDGbhIaCeTpGBWKywTRw7XCF2QdQJTzvT19QYKobIW7P+iYQU
IBF4nFgQngth71TFDk/uvwdw+hzr9k42rRdMA4uqHBETcHdfhvRAaR6Gj96cUDXU
GTCQjPkbwUQ9YcEoZyMQW0Ku9PE8WBINVsCHLsNua50FcU49SDnzR/gvWc6692mv
eFVQpu/9HOzO5MWFnRnGHKHaIg/FVH0CL/tqQI40k+ob/jfBMPZNzh+h1LcKcdNg
TglYBzhTiEuj8aEoEBrhACf17ENhfbY0j0d8Ww+PwqrvJJGqkTkzzBIpbm3WCvap
wCYJnc7AsTqPKnNWQcj7WyIYQnl9nZwCSfNwfCNUILAqTmQ3fJ4u1y4VgNchf/i6
rfRuukTVrv5AXs7NKbvSNrJVq4to0GKSNVan8BH2Ao9IgrqEdHkHfJNSLNfsd9xz
RBnhVEJphusfGLB0Z5TmWlo96yxZjhVyu1GE7I2Aq02bu/uswlwBn8TPjj9MvtpB
xn4itDU3pOcQx1Dwo1tFXVsLq2tgYtJqsovM96XVIR9mDPQuFwpmpL8thzlt2C7U
k/cwJp+PtlE6YgMyZd5a4nNqluWebYlZO5/TICk7eNnBWsNKfN6aQUGYv9hKtpA3
l/k3GvikywXqOMF21GNDCfcBi2k5HkmqJ99Tz9kNGcg8P5Rpl/UYQwDwCLCVBtbE
/BVV4tXx9pifgu9DG5MfGim1lP6FDAZSWx5DvNdEw07GUleqrPFkoUeihsSAgxP6
o57WKt7bToGY/PVwrBr7wnnyO7hG2QMvalUTunoc4vjW/I6kmXfumnQ/y0oHivSL
qSiEMUbvAseqIIAfeS0dkIvVruttEheQK4N6mHr47TZtOqAeYE7XueFIl4GSNRFH
gB08tatY45SdvT1I29m3VcMWvxZ0DotGeQF7GenYC/BcWWXgiNM1aTbLxjZYkwSj
oHJtyR5bkjNWhM4b3z8n2qGMg3mvNGI/CSWSP4941+rkNwzp0y/fy1ACm8uXfle6
mhD7CDmBXtYrccLZD9xgYgy+EhiXztFLroC3KxYKEr30BBOUZqthnzjhdw+VoIXS
UypQH2WVkVS18avMYNNR3tDq/Uft3yFeY3gpVbiRAnFn8gpZe5RlEnmd096lQTMZ
gWOKXazKtrXY/FZ+5O4bUHU9YLlQPYgPh4ACQNFLv1nHD0wLj4YTdrnqEAgAmexb
NF2lPUGWT1Biw7VhPPtT9sffRnp788IldPss7H54Khnto2edTGiQMB9dX+i+/TXk
opgcEYR2s5W91zdhGq5MMqlJ6K31CcbiSRN0LdBcWOO/SoJH24c9+UxE7lh8seSq
7Aufahf+HL1x1seNGPWSVf6e3UCz/PhDdIoTHtEeTHIraP26SY131hGUZR88RWvS
WiqVnTdoVIVuSRmDGo6zFh0abg0sx+r3hZKTD/84UBhz2oOyumFIQ0FtDiW2+wc7
uRalSkH1LodZp4sudqMyVtaPLDkBkhsBBilBvZln7Zv6FDsclkQYFGMlUWqrzxZF
io1FOH9kww0YgUToDXNbTupIHF0gJjtggtUWVi/OJp+AYTk20fXyl9l9E8OdijMC
hnqz/LvQcppL07Kg9R+EoeLtYL3VSFHv8P6rP5TKZeYG0PfAmUCq0JVRqrWoj7BG
Fz6LjjNRZ5Ovz3qS65GM2XFiTTmnmhPjw/mu3pbcCHHwzbtonIkQrNquMFjINSa8
/m5ssffrhOPja+yyl5TUG8iMB4nlT1NpR1Zq9pWgO+rH0n8X+o0lRX9iBD/mitAJ
7NCotJfKoIhX4UbJ2UDoUJ5/mMk8kIIxQ8NEAfcP2UYnPC4ZXVgwifonfu0Ph1SI
Kh4lGdAFUt7yDhAOFmjvkxIqzP70SaSDOaNki9MONTemuHanQs+xm+SYt43UOsoO
P+MtE8+PRixYufxqvwWsXHCQprgOYYaN78NJsLsFwwVwnj+K4zpWToqXvLmTh6B7
BuF/kxrCmfLlNXOuaugJ+OGGd4vu4X5fXJwpZWigxjRgC9i2c8JL0FVg3HBu+WpH
e8ldqhvuBxY9eqDW7MTkP+3vQyFCergPfQm+BGkZEB5CKxQRRLQxOiWKMVTKtJpG
3UEgevBDrdpi0q+DM8yDFWA881MWoF5THgGJFuUwI8ac5LKFVe4NhPaDH1VmsaMc
mpsUDb4JYwhP7RT3N1JOP/hBbiOgQWrRD5nRzWkrcx6Nx3HFJiGrUOMwNIpCrl4M
YtgpMNLcNi8LOcrrCAJCEODYO5WPDQMoDJbdaAPhz9UbLihet3u18N8jlo1ejFxv
v0/qHNFyoKTJWdzzuhgxSM1Lr2sKMjgRMLRZ5Penf/3NdIVyeQtv/HFi1DjbX/Td
dgzsnKGR9VuaNqOueHwcnfkPMeFSWSvLhC5DmRJP5e7fFDyEy/+turjjWKZVCsv0
RtMa/NZwM9PNAwkAJXx3Ynqr3tFeT9i5bsHpQbVlDGa8VtAW/3fzQjiEekr/YwJ4
UTTU5/GkawyYyypcCJdzgM9Gk8Lu6dev86iiLf9cOMs1f+LgRH+I87dCb9Fxe3AX
Mx3jUAyVyNKxZpyPpoISPECGJoC2FtbVihS51tGjkixu1PgXnLbBcDgvD2lKpQJ4
04uLQGgxRMnbKgjjRwx96u7XD35nArNuwPRe6B1NiNew7UHE+X2wf4ndquU7XTe1
hdI5HrRQVlQXNuJ2D33qsxb3Oc8n29ILk9LlFHy6LwZURUA1iStOc5me+hSPsSBk
XFkG5OKXsSMxHWSUfstbNdjcmYk1PIWcrPACeYgAOzyDw5mc7u0EwVHFfUs/qyOo
v861Ai0oiGvRqNr713pYpj5g2kVTFTxXF2pcii1oAw5h31B6qLedSmv5gzcHqoLR
OCv44H3J4R6U+wL634fdrZLZwBcQN/0yn5Jh6TX3AxrLCHsu7wCIEPLj5K5hZq8u
a4e9pNHK8howEwQ6//Id08wdUWUKR9fUHpC7Lw9lj3Lujv1d9zS++6ewDPzk78HB
YaP4yf+1DJ7yzH30IKi6j38QXoJbvjdG5WrQzeXmadzRmAoDhKIiXEqpgmq2aKIJ
AhD20RL6FBSb50a0RBeIQwyLiAxkaCWkcgRKSP8NQOaRS17mbFFTrkgvfnik14tP
JkmAsUQK8ShEFoJJMnPWwWtBrHIgKb54299Lbs/qK3hRb5OsSZ74n/yK7ReXfoMW
1IAektVuR0Bu6tYY6H+yGXJeEBWdUT+52B6MrIweULRWGqO1nw8TKsVyMfoJydoF
KmcymILBy1eoL+rahGU1ZY/hWCM7Vh4q3n5I9WcXrsb0RVKV8r3J5LPE22USdASI
0m38heHN9pphQeW3IqCLV4jHLsI3aU/KhfxrP4pJ3LgylfExXlKs8MYVvvgN6QKH
/Xby9S4aG+iUAruyYZUh2Tqbm38i0iASpkrrKkzyZyQGL794qUZjJTcU54mx/x62
+as5OMSNvxyBKVRMpdVCtLyD1pV0VaVzwigstt70qcOUKVVwcUrl0TBTKg5QzOjU
bWQQW2X9kpf6QznWjdywPLtSecv/3jlZqhs5CDBKmbaWEQzSGl2Yw4hee2yu/FQm
zBiL+3a0a/q/8tOSBJim7cf5mPdFkrpEdyyE37RkL10e88/GJ7Kr8IS9QxMfbiZj
tmahfT00ICQFt2tW/g/YvPxDSj2KU1Kk5PKcqS+Apz+xxdKQQOBszgX/c8zTNYoT
g34AxG/9at27GRjWnOBTisZdN4BfERD44Z12oIRq7CasMF4wktnG3EGrSSeT3Dof
tRV8ZHG049zxpiDJZwPP2ZHbmfyfABFQf/fml9HGXSUPjdTMKE5chggCUw/k3hxc
KTPT+j1L0c+V5z5uFtK3u4bLr6xDYrB7LGvNxFqyOHFADdfBc2+JcsDtYW7bzrET
Z81daTojrtLVzGI8BuQG+Ydvs9YeNswk8N/Ady2kZFWwpEfsqiuAoUUn2VoQTxo/
wSdRV+izEYVzNytMStYiQXxyxeDVahEamzGpQVa49V6dh/QdeEgpewCs4LWg+M+4
Oqb7DVjBrqYM9jtEYIuI7365s49dCOeULmc1DWOwtb66jowmsoKhWplMwJvILnkL
bXVxN4Ag6qWx7BQKSCRc1O6kkbwSBBY+2qFYnp+UPbuwgLZuRlj0IVFHhVUoKU4d
wXV5BMQ47/mYRI9mc7o48O0kZNAgAUTfN/RwsusR8BSMoLzyEZ+/p+ORIzTmc2dT
0SN9o+XqeC8WTgXPcRUPvSF/qkAkythhdUttzu7jEAByZlKWfrG5L0811qTD8BwE
RWNFOgpqSkyzctjU+zgUW5q1GLi7w8jmmCFHDVNPtXR2IodQqpy5H8ytF1OUZUvk
z8e5aOZ2yJr7VDuG4Rh64dyKqFfMLCV6PEUXFEU1mbRPrvkNPS9wYBXKynmZi1Et
+EYc4XSmfjryN04ufqIuQFIRpXN68iz7GIj3OSb/33wqpr+qaXaWki1piqXhlLyU
KRXX+t5nRrIGR6AXqwnKv234inDxRDvMv81JfQGMXu46HG+2ge8w8zHBo/8rdMVg
EfHLGvK0TEYL5qulKG+ZGjh2Sym9BPruNJRZtQBmPaBo9Bh72yRDD7p4OuKTcSwc
NE8xeuMmZLFlmfynjhLNR2CJCPvuHltKhwBI/mNoPdw=
`protect END_PROTECTED
