`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61hvQf5ZLrDfHM5LhQbaa9mITu5rcZKuU40UV/tdlldQ0W7uwFy36Mmt9Tfde7FG
ha7za4soHdBUPHIIpRRuDqKYlrqR6M864vIztwUERedJ+eLLhF1WrSYz2cYcx2Mh
RVsAVAo8l/gFt62WUVdLrtZGuumSNRRJl7DwlTwtWN8qrYfzjeTXLKzrk6W/SYAn
PWKM/AhWc2tUCkg/1LySGkFkv/GVcmtww325AcGrSXLhFjtloTkk/yNdPoIWmGPz
/Ny48BDQiQgv1pxq8kRWaEEPs5MYwCE5s843TxGjBmW4Nx1bgHzUKcPfkFnh33Jb
ZsAFBbTF1WMWZhv7O8z7RmtyzLX1JAwbE8AKb36zradH5zOUAZdL2u8o0Q1YngFz
5o5NOwlUWDEEnXQYZQIsEw==
`protect END_PROTECTED
