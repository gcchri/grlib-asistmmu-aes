`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qAMfu5qDzhrTfvE0AIdN42Uxro04214NiK1WUMOUb+n0Ux1zVHWi6zLO8EC2fvd8
XHR7KRKD2LFQmFfshZoaDqb9vuf4Ku04MzpWOf0FAxMksXkCpY7EgmnaE2CjkKxd
2O/tA/dGwv22i5xvYa0lhMZYybmRQLlzIbujRd86hMQfKWi7eMRO+97F0jI040iC
3eW22VnovPl7yabRXLu8bU7deN6e+3DStPP97JymRkk2Vabtu0W4z1YtNBHJPm6n
nXonojGt1iCcL6HyKzqJWy06lWZG8QBnzC6kKzQsjSLN0TJjGscM8Dfs4ddXOZG/
/DWytZzpKFWP9LgyzLp0HW5Ms3wBPAthXhNkU4XsuFKI5W1OLHaSEHAwwsT0IRjI
6N8nR0kP8XK5ErV5hBYYCAUaJ3pMIvjvoHi0Y5fWBcDfWbOaOv1+8Ile3GquPzHp
6f30i+EHvWhTjHmLOonGol0tzPgUKAYC/hGOXJsZy/0=
`protect END_PROTECTED
