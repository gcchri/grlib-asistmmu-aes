`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxRLshmdHbidCZpyLrQWWsm2nQ4wOXEsEKqxSsE3rS9X5dOC7H+AgGB0TWoASGWw
dXTlV86q2HrHPOkTJJTW5zreMUK6EsABM3TsxBGxvwYtAXzN8o1R4sopWNQyyWwZ
fdN6SeP995iYB+Wt41RuGpX7AzBy6bIF/zGt1WX76qOJ3tJgZMiThT+jWsHTeJlo
qxmVmpuhDTxgLRtMkRxRWBPtIAtZEdxvuCWMHsVPG6MJXpYP6R59YFF+YOfOp+oI
Gx5lp1fL3llV89EA2OIhIA==
`protect END_PROTECTED
