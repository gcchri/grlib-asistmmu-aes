`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvAWGS706NKtT9YEBLoCkrp/zrSZDRzKTbFBA6JFUXMQ33G7J70wZ6pzDwZZUVKD
kE3VkBryZsvR9PStnTwIuWwq3mCp5IyWKgLcN5o45pe6z8YzNnloG3Y6+Gc92Ucw
sNevye3srdxQ9ecG1NJxP8ykgxNLyKPuz+CzfMZRrbr4s7EOjYTkpZV5se5IG59R
27l4OLQANa9rZfM9Wh3fHeHbVMG7HwoPlGhLeZixoMDYLsbh3GI3MXOa9jo/VEfi
6kkmwDfI+f7aPk9tWK5mWiOhVM07L9SlDTrlwOLUtgMdY9/BPID4h/+TrDS1cXTM
URWoV5th77Z+kckyowApE4KRivUJ2wbsoeI+JQvfGhLYdnJWQzdwiBvhaiTrWdl3
JrbOSMNzs+NBd+weP9t9/b8OhHxLPZJJabP21LRPwJ37Q1A2P3GTTWbteFtgNTLr
OigjhqI4aTo4Z01zz45RjlX9z9rUQJvQ2qcHnCRLJkPJPXn5kKQWxRoT8SUMuiS8
`protect END_PROTECTED
