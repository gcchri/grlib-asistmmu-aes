`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZab9V1SWr5fhRd3H8hIe73tTEiHMph4YCSBowZd0rFpDz3Hnh2ofiz8nFbEQHa4
DQj5j7uRBjKEi6MoBTsPjb8QQ0VOxAzmOi/ItM5BiRsyoEioSLRYZZmiEeSZUUpX
1Jde/hZRaBSTCR32JPk+YdO2mr8r0NFM25jZHFPWEmSBLMQImSgD0j26ObxznFOT
XYlH4W0u4wdSE2//EkHngrRELJiPaCDBz7aTtiPFY7Uc24sdg1DkziRPwNkgdojR
dsIGm/GN1Qmn/v6pwuoJlMQqsWKU0lgVV0jZhCW3baKKIpJiNBgkB8jI4Uyi6hw8
k0WRcdBCHkaKxbtVRy2US0GFpS9OyBpuhM2CnEWvKZraEOyQ70HZlrCODdfTRzfZ
uKiDgYWuUnP+5EGTnceyL3WJ+LBDRbDs/NwLspSeVYQG/FC5SLJoNZbFmtZYff1A
u7xANXHiWeHcIXu4MErOYIWYBg5iN1JmfMl6TvGJce8uDEouleYcsItL3dNL79BM
4b5jrTe7kFwISLcFKkyK2wBCRwyfxdyf6MLL311wORRQibnoNs9GhzHYjPjr8vsC
okmegA/LAE2BgsoDJ1XxblTqDnO6xzScyEwJ9733eVTFpHXPkbXWtb5pnrYYZRfZ
PQv5Z+yh7qxAwsMUankiwXHFNd/NlFQBHi0OXcC92HR2EV/GMZ+dOem/NSRVPp8O
Ayf4V8Wm3Gke7jEZYTq/vg==
`protect END_PROTECTED
