`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bigItXmfFOcg0glD+bkiFsQZ/nlKgRjWhr3gcMXt4r4LqXVjPdB+VrhKDXVPZevz
VI2Isaw0akvuHxcVehQqu9wAn5BNGsJt3BMCwX3U55mKj3pIZQ7JMg7rZ/HszboF
MVeLp/dvPR6VmP0vJSsOSsHddyAArNmauo2EA6nNLWCj8ibcM5A29nd1FptQZo3N
0Y0wUMLkWbjW59cdrBCK9KWDorzY302/qZd0Vnk6mJHC2Lp4O+6lM0KtnQ7UvvJy
Y/YL3EzzQwVXPLjLVQ32gnDUYCj2Ex291DWHJK3tXMjbsSn4Pqcfgzm/kaCkjg+K
G9y9OJ2HSFIxvx4p3PO55Uyo+wjSezsVc4t31QbrUUh8eWGH27TVJ8tZL9BrgJqd
O+gwIpyKqWHAN3CgMyU8gi7M8lDcDCttxVXL367HojAV3l8oo7sabFU/iHzDVSiu
f4z7kXqhm4B7u1V7sd3C+bwWarmFH021BamvCUjnNGlu0XG0g/7IuddTIpT5nwUT
uqva0wymHfZcgJEjTYGm9oeAg0ye3wKIN/UHymviHlpS82fAwPz35a1I2D7fC0Xa
Vlwo/9JQRX+PiiGdIycV8g4iFehKRBl89K7pFkfj1Y5uBfGqT7hZtUkfTfmb5NQG
gzC4g1/rCQfTvekwzzh0p06zHguU38KRpbI7x6T/wa0pIPHH/RsPbh8InWvj6WpD
F5zGyyswYiN8jgP+XPKikGThMtiA5WaXeEfpEW55xVZGAq7K2F2ZagwST4KCiSqN
hDgSqCcdqV4a9DCsub9cs97HAqA0Wydtd7gJdKGnWLGAIZ5osvpl74cQz3g+5u43
zorms8NPKhS5h4VQnKL1QMW4L2MnB0kHmJzo0KnYzc02PCuWKJGzPOdXZhABKDVt
n9RXdrCCUcNEPGFsuUjYG+EQfw42CfuKpfw79cpdtlR8fT5skL/ZMVxR9QnPEddy
amrO+H8HiRvYxHTcnOJMWV+4l7qvHguhNnMdUpCGMKsHD+U/90LPX69N1Zx2nVoU
`protect END_PROTECTED
