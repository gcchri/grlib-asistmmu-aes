`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+CdPX3C46N9514FHltW/SGnaCDVZGCmADwqWZ+IVfV+WBULA1BktZW1Kvy+7n+Pv
Hb31qTHpzEy/mF2qchYaeJf+sVzUmFHeFrH+1ZZpj/tepqLVjpvzteKGH9uCsnia
rJn2hhfLlhUM/p4MGKM2VIDQ8Tu2ZQxhLixsh5bHbn6DYFN0c06TzH+s+WLuTAzn
UVclkdmw7nGGkVxwFZYD5BV4nhwPDJ0EIK6q46woJaiAEtGoKiO1wr9pusGAFwf0
UoKdj7RARVOsw+bwe0KepQ==
`protect END_PROTECTED
