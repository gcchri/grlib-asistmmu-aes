`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
luzzJq8QwHcgkEslNigdDYkoRGvfGU3/z0SzKroiBcXHBeQGe15cIwAYaGOlJD/s
kqPD0bjk9f89VuCZASR7uCv4tlvyLXTiSfugOEVdVskGwny+kTSCD0z906DLExJH
VpfhMQOdccazSM/zW2AtRKgc8HGu5JlboSrVn8SnK3O8G50xDasT5B0cZ7mtCtoC
NCc7LOQRoqMjIoxrvIdkC2jGwLobEp+5tE81Vt26F/tw+QRtKgHc+TxVy17IAQbG
J8l9RbeG6uAzkQQZjB0Q7yd5rxxid6wr5bK99VEEzS/pnQyYirvkUUIdVN+EHDWr
apFuThbll3g87liCpERlIdYZ1JV0ZSL+DKmTRjKZGMcO+5jQNXxWlFOg2InJvKOa
NOqveeh31QyjQ1mPFTsOM3nf+MBqS4/zT9Y3yxpgQ+JFWehFfNYbPdZZSe5jrZ4R
BFqh41b5dmJ71gaHkAt2r/oZ8Z4GuWj9YoVXci/DRVxawZ3dhGy8svKSEJAvLata
8LvV2hFWvXOHxcZ4V7TsguVrPcHSwajH53hJ9L80DK4hlhM9iZgyObYrdTUrV9C1
y9nVdM6AnoiLd7yuUJgAY4zKHzPtwPQG3tOB+oVdgtmDV+FsBA9+ssHigYb3hFhv
S8iVqDuQoHscXN7DqqzAZz+Oz0jw8dCgtgOoalJCHAVIF9lciNiGzBhvalWXB76b
yPXr0zypxuozUj2/9tAR+gtuZAut72PKtBuAAbOunX7Cg5fF2bW7eZi7/St4vI8X
V76ikKpEY1e3fG1qDklBoLD+jJUiTP4xLUXdr31mO84SR3MVYLCQ6vjV9twZauip
NNyR3rlwoettUJQQ6SLkv8rBZewZ13BgdrbRO1hs0CSCZ2TdEMX/RH+fZB9yH8pt
VpFLZna4dBlSPUZUpNCbPO6zcJQGCerv22Jqqu22alwCHeLvvq/tVptWid+4XSpT
jhvDJSQuy5XWOBSl5KdPMRA5CahPutVJ5jPKdblx3pbRPjauPQ9whsvecvWwSZeO
N/X0ZIuMJVLJFNG6edGdg/R1R4LD/650QtInDhLCe2LrMsLtCXzMxaz1qqQX5Oei
YHhmHPGxo/fVIGAUtid26H4nShQvZ4+uo0Qpftj+l7IhQsfzItXdjdAxYZmDqQ2R
XAutyNneVFaBzh2S5kLtBVHm/WzlT4Dq7ZFw6KJw2fBTR9KEzIKBukTFKhLnr9rF
N5Kwfdj957wADfiQyoSQeGMSCHd0Jnpdh9O4PQfwcYh2/Zn3w17Ni/Xks+OzwBZS
6MBppMH9P7TksVBer/zHXMK8oErAv2iV4ezz1un5pK5yoAz3nLVWE8MVbwSEbHtl
crT5CgQPMVeU0UrFjrI37Cgc9Zyk5M/ANmpgLb/eDHDV8ErfZ70fzinTUvorv6a3
GQbthFPboy1Q5sPaJwxoz+uMbqAzecF4bS02UBNqmtFZgIoXjG6IIU5rk3OrXLEP
Dn9mz60M5Zv8xsQrLZ+BlxWPf2/ZTE1alXhuVFf7GC+PLyVPiOPowiybctJJV5nl
IqNHcMB1z9ATa6JWx+z+08eqm8eFBMvgGxRJIhMi3vuKnrpGGOqV6/3RVZLpbN2i
oy3Wg5gPc0/bDwojsEtQi4GrqXGIFt308KIPdYwJvkLDiCdALV3bjGKfO4MIY7nY
IQSeDyeMIX8Ak/KSZnq5tHeLpaZTeJeBqFrZdcZzP0Z8MKW3aWNlmf5JYM8wd3v5
kQnxb6sfEODqq6JFOkcTjb4BwPDxBTZXv319e6aKIahVb2NbmhXepSVfsyNRAMvM
0lcTzl2MdagWPLjyqjLFax8Mqf8hzNC8CAmWWzQ4P1mrdy83zaeLJFu8GWPfcmFE
kFQ7KQ0wKfKrKyRXXFyWpForSb8N1jX22PFQANRJf0UESpCrXVGGL1IwQOhtlEqF
MxV1848r+pQPdjk0MkrtOWct7J/z3PSmDp7i6yYpjO31dw/FG4wpaQYJMFVyq96P
50Bb0muET30ss+M7KqI7FN0xCryRkHfDnphtWh8+WKnsF9BjgpL897UdTrZmASvr
40HCKlp4ZCuTHU7bDZnft/51a3vhyUiwkgRVlabiz81q9QRs7e48uH5CBV7RsILt
+pLN18hi9X7DuCPJARAtETABEAzt1BQb11Bz+gWXs5dV3Kby2A/Hf4c7xkGEvbx5
Eu+tOnLgcR3u82jiJH3NDKa3iwnLbnKLm07AgunBbvZp9VF8WhGrIY3kmrmiLHIQ
puDOVxC5LaHRnzAXm1dtfw9bxDYcrJ6WjZArDM/4k3zaGA+YVRjkpKLdlva8z5db
f8LAS/Hz/xq6QINW41MK0VzXKjXeZ/ciB/SmGE6CUbGcERa3s/O4K77rHdSvNxTu
xznRcKkQPkzedfUTUqxmcmSFz09uegQxUMdzeOGVPcjPNdY1hJXA5hCkK94peFv/
d7vh8pMEKZnBGe7/NMMBTqMu2zN+xvNivF0xquA/vdS8EeIst1e0FT7B+b+xzDHd
8q0n3mxTowyMtdWysqNb8/Q73xzN2E4c7u/LHU6DVkrtiXzVH8195VqW1Ur9NQwC
LxrQDjnrUo1UsGuyg7RaLR4umCu3EWb9woSdkehtc0se0UP1QU7WZlWlQ3jK6ypX
`protect END_PROTECTED
