`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5umwCG1t0EIHsqPYYGaMRETbElvXRJW2XxUoe/xRmbM401btOiVJy1AZuNo0FHka
g3DghVtsej6Ky6HreObCdp4DDh4347qoVX7wL6/PkkURlzFKd4lMCDIvYe+AHFJf
u8oXf8z5zCyndGJVibXl52sUxXcsKZjgbgnBrpLg+Gfm6fg6r8X1fj0AbB+EpwRZ
nkjH0LJ9lo8FrzOMDJwe1N6RyAT8s13k1TMl+ggth9DPbXFT6NoMumR2MG+7dmTl
RnyjhWAkT9AfGGsMh86VPkGt6x4Tbx+MeQvroKdNUeo=
`protect END_PROTECTED
