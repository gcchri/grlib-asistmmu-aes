`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e1CHZr+Ku6eb6bumRZZlsHOFwimmq/X0QZm3nq/M5xr3y2EagGY/eiA0xlZE3n3J
y0irLjoSmLrv8S6aBkpU2sZ9f4WuuclfSCd1jq3Ud9CNo/TWtIK4fB/C5Ph+ATEp
nHkhQi2+uIhmSF6dY70VflwStdJpiw4NO9VQCN3Fnwwcs42I0R4iSkzM3FZHlNnh
hY1Nmo/0/UXS/iYm2GyrfGRLRfEBhbJ1Urrdanz5z07jiiYpBXeNUIpyH+5aSQTo
WJN1SZsQMnabLsE7cMFcqFi/io6rgpC9zQR6SPQmIo3ubg7+4Ndxew5ri+VE8qF3
JZLEye9bE/A6SSQ/4tdwvbvJCT5TJNdH6mhXZd9X9huV28rRDE3w3cetcCJlsRDz
kCHUiTz8+HSdbr4aOggeM3dNVtT5rFVDoN2LEBcz9x8pqB0fh7MnQ6jffTzL5GGc
xny3DCqXc6RYuoYZ5+dLfYiGgbGYWJDrTaAeR9nKEo+mDvcmoVNSK5RjlPdvUj/y
NaiqivfQ6whVgsOmHCH1R/YwR45izHefixcaTwex1IbeKi7sr0kO1/64ijVMxU9t
8cjLttPDY94wjcthTFYMpZQKHvAhPfSvJ4lcoeGOPsDCsK2z/Qhj10N4pwvIFH8p
tgaIcRLNvdivLvt0V7zE6lzXizq9K9R2SC0qAbNmZLTja9ISQg+XD/HdTj9ah3DG
CVtCFOBchggv9V0MaoS042X2vMpdBC/Qa0GgxdxGDZtw6oKVGCS9V3zOBpGMF8wV
VCjNuZH6DYt/i0ti+npX8a+5rAfpTVn7YXfg1PwfBGkqLoOnnaHxTiUM5ncJIWzb
bTE+jLJmBHMSKh2tjlxRvHXzh+cQBoi0/Zsx5wet7bOAU7QOwUVgxIYZzK/3iy2S
BfKt97bFqwijlJlACOir6Lkf0bmhrlpiMEjX0lupvm7qIAdw2uCELApH/4q2eteF
tt1iMKGFRSHOr72yuke7p6t/M00Qo0bH4OEZyAkWEhIEliQ0GBR9yLWzc7RwQVRn
YLnapyG+m41+kRaSfNTFtUfgSsll0X2xVGVSGDNQk2u8QaQDIQIToxob3tp+5lSH
WGZJZEqRRNbwuVXKFMLigo6HcNg1k1ywne24ibOf8CtXNPKEkSea7YOmDQA8w7qt
qHbIHQETEvndxIxOvgFvjNPFRlbs/JN2rPHQ0y2zb9KfX9u73wKtMbZ5O7fEo2RS
oeYSR2Aybz35Cvo/epKejczW/AI9W6791qTqGIv8lsC61fwJIfnyYecURwnJP0OU
Dooprff5t9mgicJg9Q1+XVaNPJpmZ2A9iO8eV6+xy0R84slfiQuChzYbHUWdacGq
BRACKW6SYx8Ym7dTDvG3qO9gEi2OJdm4Zu7SaiyVewhntaquqTCnfN0FRrzuiwO1
7lzlrh8e+flJRvN980rvb4dyghQj7O2NxNjjiKSjtscsuMU+8ALJw4tmPulJj4KC
A+e7UpewvjaQusQ7CAXJtKPxZEE+Vj0s5smAPpYw08XzICdH+k0Hxn1nwRtqgEqt
LKkwzg29a3vrdSyCSY0bR8hgHl5vaHQWW1McIhJK3jjY9bCJrLP4YZ4DrXAijdfi
SLmWGuxWQQrFd6reP53i0pMsq7bZWDpcZoyRo2wpYwhoemwd6277qjd0JuR/wZ/X
PWi+wY85HDDlk+MYeVT525K5vhC01YljTE4hQ+JXqVF4d21IQCilw0+CLNHM6snq
hGaCTqJF307KGoZNv9xpz4nIQYgsg2Ches2pP9JvG+VX707Wn0rdq8kHnWZn/grz
8Zet8BplTC49IWqAVnTAsYFAzqu5+DNuWwO8J2+/lY+lkPo0wXTYCWQeCsRRA5KK
nMOa0D3HbgOwOaK5muS7vLUaIR45U8db+glAbK99cIuM3bZlSFCuSvGN1pOLwlWb
ZrISNVYlRL4fuaRWnyti+MTIqtALGMOqWCDM7+9zfvMo0aWt/Q6CGwegJaJHJjW+
TXub7BLk4A/I8To/qy49ckUrpqp1fAXDEkZ90GP4vz4SO4dcXQRxIEyBJK8cvlWP
xhAp/FnOUGAZ9gyv8Ea9BaT7hJDzgobxRLfYUziE5GI2Xy2hlNLaiCBxQj7MbHeR
EAoRLhimyVpW03QPiINXE+GE4HV9ysIVGwAylx6MdtdcI9yRN4Zf8OSDkDEmHSTp
iPW0mDeN2hlxKDCJBHJ4JcGIGFwkpWz1JYkNrCRKGsuPUngXABzJ93tr1/YtlVnW
V+pM7owHSfJylUfUWL+fDzREDDRnZERSW6BvlkpNBhJgm5ASvSJrvYyK9uaj9csa
XFWmKtL+bfBeLrU6W0vPFr++aed2OkgG3Z4OZWsZOr+PT1t2OJT9vzZtwDdXBf0O
0ga6husBK7x1z7dq0057orM61gAbJJPWSULBqe8RKLVcttDo+EaGzQ553oOEsmf3
f/ldQmozP2M8V95okS1/UI0y9hgLctCG11T3a8Eo/vgZtZqZXLZUCCf1Ae+4idrY
J+KMDgWoRO1Fhf2ytK9m5YqH9vRIwwWkYrYu8DjgUcFPAqv+kmZ+ukDV2OYaU6CN
nV4p2GZ+u1f/TsGXRaP1vtQsGo1wKQ6pp48xTxDSmNQ+GFfWdeHEGXIjOz7yC1hx
6pousp5Cq3Z9qQ1xT/esrJIxG2a2oEdEF1qHtGlPUGlWPSQCAuKUBABzhKscdFmB
azpqY781hohTQ5fO2ZYbEI6Bwe84Oj2X9h0ocgt2zuIfr+iaNyXI0jmq8imp82Pg
xTz8HSEByHbObU8qvLtuoogOITx1qstlxs88edMxt+dBoJ1jCFOrpztdP7GG+wzJ
vahsFg/NZgojd7Sslzv0rce4wGg3j5nQEHDi2OP9K64gCEEpxOSHtB9KB6zZnAiY
i3/kQgjzsoWKAhp3zO8AGc1oiinkdoQDi2aBwDxXXxWL+jzUEMdBvWP/apGk/O5f
n6jMDnUXmjLc6DvDOY4UbWLjxAX4KBh4qdBeW4X+RzSDn+D/At7Q7YY8mK/rBLd2
R6I1lcUROoLpy4msrkPmdrlF1uVM+yq5evpy0qXjqGPwsXq5d3Ph94JzJKr+x8fC
ujy+L/4pKdCp932aLgevQdjtz94i5eMadCaoc38kCV4W93HBYra5BPV2ytAnxAZ6
d+eo4UEgvW9wYpmnbUowCL8yOT8Zgc0L0ec7QEgwbzGRnWNCc90MCEfdpRm/i7tI
8O2R6OToFyr+6zDyqAIzOq6cIMoA8n+Qx+rdxL4qbGiOCNhj+VmlJY25HZx7rJBW
6FhMGAv8GKkzOtcGGIrfXkRpv/PyM37MMOLEq4yNCQXAuG5t8uHDjA8vhg3a+t9a
JYDCj/STJzMyRIJLJj41hyczCbAZ94lLjWWvPksgCUFcdVVbHw30UK/QkCk7UMx4
TzEuaHR/VWVdzMZDYmwD+LyEQNEzXCJzElYFXHwR+1zlHTn5ci00bgmb0HiSUZq+
/I/25cZFSGeFFSaisl2YufV1qA88qfSDXP8zSEPQfVbb4dVwCHhXNMXfr8j9hdih
Ei8OCYxS0u3OWrLRKgl1b8QtpzOYrlf7TdyP5E6aFMfnFxtzikyIvz92AWAOPDxW
bS2/eYR4FVERDWbs71+E9xOLlhjwwQDgWT06bGCwg0m9XJWO+dl6r0SJAjAg9VyC
DT80+zsTNtCBSl5Y9hRMlM4IlegUsqNLmJNXlzIqXQhTX0I99ykRX31Empr+3mIp
rVyxdx+8ojN2Wc5LvBrKLqgSoS47l0jKKzS9Mmkme2tiLYe8l6n3z02BiiD8qvSB
uJ8nb5hNxj0jLGMjsz+QVfXEOxJO3SGVBJz0ZgZHAwGs9RFA0V0a1dFZd7m+/YaY
o99QVH8ji7HK5bMMSL4l8wNwBibdcacd6A9xReUQz1pPgkMgTBX5EAeX4tect0EB
MMT6db5Irih8aItpw711P8KY5tmMIE1S34+UvHPciYDXsJyr/NSHA3U7/GAi51Yg
Dv/C1PKyeUPNDQnx8HEIz8+272SuGoKCy5+wpggcWg6UYlc4uN0VXFmFCn8FYMAh
eY6tRLdCmDzyPYudImfAJ4tOsOqwqN1KJ7TRhjeiiOGNVutlcnDg/5TVVQOjYanW
163OgEzSps2Fh7Gu4ByI+bVI2/XBE+/DWzo+ie89AmjSReXu34lJrJ36arrEDlyA
wto/Ox5fs6YdLLmCgDd8Aceta2JoUmyyY75z659vVYmswfgsQLOpJK5iQ1MlExUt
bmlNPpYcCyXs71+wXltResBZ5E7mJjSTGb+b70PnwhG9+wHGQaqlEII+VC33JinD
Uy6oows83uvI1x6GY+0e2sPKFImsE/GBwfypaYWVCdRHpBNJ2s6OxUQrXkMv9y/D
4RFOjY8ByuKZXiZ6yTBbmwHJK0KD1SD4iYMtDnV0y4SCXRic2yCvlGX8Cy3KMC2w
rTjYsGWijChJGn/Z9p6PdjrglVKCu50JWXH9MTsJ2BrursRT1fP5WDsQRGYjVqhj
8kdLkGnRiZ1bAdId4scK3AthnqPilxg4Ii4So6PAobqCiNx5fiSrAPLYlcbCnvVL
m5GRjLF7HCQuLOdtNT6Bohbosd6bDmaqKHzMGf5Rw0xoh2RaEEybC5F8sC/UG8Wz
GsqpIvxnvCCLgly2ODnGs+GQk5s4qRmK/3yHNPeXhSD9Veh9SQeWLrnPgc1fOp/6
oVArBm3M4wAWdtm7wkcFlUleuioaqkuQnbA9+4Bo8o4KLBteaNyGjEcbyCJFCe0N
NGoya0z0UtBt1miHLKibyE5mOmFtODMYBn+qUsVlUc87uYRe3ZzLyxCr24UGg2MC
2jgoqxh9IX+Pwp9OaPZ7i9yR8WjJvSrRjHdTh2wAaUwxFWuwRF/3gAnk4Cn6T+Zk
gvTi7Hd8MqqG9e+9xnzNSlSlYUG5v4AqQ4XNVm0tIK5OSgmc6NiLdoby+gd6wOXJ
hPE4zzH+7TICla7NIt/fzLUeMzdimQj1q3ib6vCdmVkheh7E+yRFxtVZLBxe7c5p
9HTg7W9Kce4VAs5zqT0RqPAHSO20LuuGenMoqQj3GdJyPO/BAX28KBmdTl1yudDr
rWxe270nwd7JRJgpASc0GaErgFVG+CsAOfoDPNqcTp8aPEjr8Ogox61JNhgJ1sFg
HgN49jx8FQbkW3LYIxJWwe/DX6MfJHi/pvvWV5N9F6YUDIL+xc0pnh0jmJkK0mWG
bLp8c9hWIIWxXb8+Z4Sr3uhCyl1WIBPhbuwmV4Cv1E0CjBP/hccVZE1AabsZeS6F
gaMH/POP6mKGazPbmjXrqCc/cwCMo4NREMEJRG1Ya5Ar1CgoObAuMEo1+dT+NaKk
mBU6AwYIp1vQd8yBMlhd5j4KZVMi4ZrnFVHOh6pcPxsApkB4EujYJLh9YHYwWIAX
PId1sIW6be323HYKm0yM1Ku32WDN7Uf5NiVxPUf3ibRDy0hWju4EHuRvQP13U7CV
PTqCSKy8R4zPXJiIotmwhkBTEY/xUHRB8jogohP3PZ4spaNlsnDYRPT2LZ6KCdyn
qzc7NzPePzllvOiMJxx5SdbOZfg1dh4tWyioZ3j1lVs2a6ZbiU3adx0x6I1Itq8g
oZbDuZ2ec9h5mJ+rNUngLDmND91zgcifLWtoedWb3vVhhWN5RdEYMgUdEO3cG3wu
RP3rSQORTyONndkUeKJU1p0LANOfJS7E1J6gRxu1Gcrfs7mVXOs2QcS1P0IT98zl
5rwFM0obxotkWXCD2i9AYrF9gaMFjtU/qcOgWVGdoUji/nbVRCtBT7DcyTM+iInQ
Nc79jkGkIRxWYCMV/fzgxVlw0J2JDhW8qvhn/l7DlUS6bYbynM1L/kKleTacKsp7
kWslO2olD+alR5qy1SlD/I9EwdL0mq/rzgpZ2T87mbJ90MjyCz7ximSianVGjKxl
XX7RWmals4jVExdrz2I043EBC0tqDUeXXqYFH1TlkT0oQRcJPXkMhBiIzY2JyxwW
rn6G2zH64IWJCK046xoRFD1EZfqHS/5tjfb/vdhlEDbPf/jsVVce/kT2kKZdNOsV
7iyciRvruTU8K68lROAy7yzSMV+ckJu3ZjklFOe1/pdYqDYXdt4EbAcntFBaUXCA
zDFxO9KNrmks0DyUmFFgdRwL36kCnScgcFiO3uUAwdVmaNWL3REGskut9jmXwXix
tWST7iUTtFDPjrOjaD0qEbJtTBOwrbXjM0uuCRy8UlIAGpT8SnviwVbgLxHpR0Aw
HefDjPE9pGgAtfJpxlyLxCwVT8Jx11/VYFJroZgesWz0oRezKUp06vGh9Cc4HA0w
w98A8HYkU70Te6+WbMLMqVTq1mfupewlu/P2M5sl8asLfoStBulfgaHAAjbduftE
UDjdFb/03np1yL+XbPGCd0UzK3l1X684wg/Ja6HIuAxSxW4VmO9xjl3uI9sCrK/q
qQ67G0dSB8xAO65ykQrzK16NEFy04t5XarznFxN00JF4OgSiaPkAU6Dr/1oBu/Rs
kVYvhqDMd+lOvqj/XZtpvHOOUL6ulfYKyyg0MWvk/7oThxSHD0ADFXph3DS2k91K
3n7gXh6mSHosN0QKTEHyBplZjcaC0xKIGxgHo/iSxhhlMcREUyTO58puUse985mD
OhT2gBJCRosaGa22nssVaEXaJg7cKx3C24IfmnD/CIfK2jHZBXPRV7EW9m465WFv
In2yYPkSDJEugXuNf9hrJvsBQHdLjuDstura4xN/tvmvP4CY9LOJrnpUZUsySUc6
e/Q8fkh/Qbua+5aQdR7KFdyoHPMZ6FKhMuKOGosWSDN67hp0fWzDJeUfZbfVyW75
3BUqjwB9zuzXi39dfDEh4/DXVHy3h4mWbxLzRQivBSJh749Fo9pPAofvo5NBPrfx
P+pvw9kqsKpO7dNW2z5QeNZn0+VPC8cZfHjYOjO/y9eHUsQ7ZdvdNoA+RZqt290X
fHLbGfEcl+a/E3YQKqNYONOiFFgwh44tUniXewukCZCsJ6QOqsm25z3R5u63P5Kj
79FnDvtRUz9we83XaBMTmZ98PNbXFQqIzxsjb4qzHqen5QUan7MxwrEQyV1fq5Cc
JOcc/3xzw6NGP14I8Y5HYI4cUhHjdQteg0vq0MDh196Nf+WaGApJnQ3+OxTo8y72
kE9jmrkNJOxxBailIrm0UJ+2OtOSGkR4HfmuvVmLnoRc3qV//ehyn/sLd8Y8d1Rw
6m5X+acnFEo9BwoRR26CtiQ9bh2lDou6n2Y63YqIjvk+yHpUda+bjve2/TXEjM7+
ZsHp9/N/scdrdLAusWUCAGInZGZrwQyIYzAO3LmudidG0VXXcLZ8kmYzIvBcwlCH
UmBhrWhR0XSHNpAxVmL5g4+U04Mi2EunSlePvRjwAET51Xu4zfeRgcr11aUMKCa9
iLWveZF/d8sPLIleyneePNwJPN/X8263eccJ/dkWSYeOgi8OumVowyBvYkkKm7u4
KTSOIcEozYDlCGB7D8ZlWf+XRyH6MdkPS5uP8e8dddyu2e53DPAON0xTGC3WkrKU
DZSk/w2Lfy1cpw/7G1C1cB2qufKaB8pdu3oCDEzeX16iFo8NiJnf88NSMuZ14fNG
cn5rBdUdj4mZbLMV4l5RX3BaSXq0ocUdW6tZ3COxzTJS0Jz9p1bGDE5tB+TUkWj2
HJ9t7d5P20m3+INSjx8q3xApErhlTzElnOWqxHtz8uX3YMGJ148RfP8JGkXBSuyL
vCf/khthUWLciN3Naw8drP0UrXZX9t7MRmFl2Xh7Rp0QAm5/5uKOWXO3V5S/Z2ak
FB0726fUQvJVOY0Onyd2tcAnKhAvNxsoHI3I9TGR7P6cm5CfIqJq6XZVfmxj3rq9
cijOMDJAZACK19x93awL258LqSQlki5c9pQj04cyZ5BhhSKulrHAx4YmPiZzdUzE
oAKtUCLjqMnOyZDuEtnvSerYewVCNFQISLxH3TIMvR38mwKGQl1KoIQxfexOMclW
ev0UNvRNww/fVmCg+DGZl3k+3wHkifFiVNR0vNCXaqKg/Dgz5p0mSB53Yl1N5zoU
87rweQC+jlAW8XMW01EJDBJaU3KoH9RXy56V1BL2U62dYwqYB87fEVtnGUxHh76y
4JaUWL10Km+PNdshQDO4gfl23OJOpAF/D4ivtmKDtHVUwcniFBJQStAMmH2fAPe2
yTkf/i23r7oFVBMhoJ7f6HBOaLFfmrro4AK+CBeKdHZ0LnlBfRvjkftK3v85L+ZX
rdjvwXifKUmvfFLgdtn49JoKQ+XFjdZbTY1nBe/dHg8nmEl/d4VEFJzoWAuiCLgm
cpkQKyuK7ceWahTfH/kheWtW7SIgxOel5syhXzgVD1EZrAHPwy4Fbk8qOO7CoHk8
8K4SIYauyoN0RHK/R++Zwvz6xAg3pH0bvngUtsRrspJ1i4IJSGbcBNWSjXwrdB3F
kp1Qhuzev2A7bh8q803pzbdUPAsaxc4a5seAFxAtD3lgLRJDvxzghFbILXqn93h0
t8gKLp06peUYNyeyp4ViflCta0gRmNfj0fFh2aZV5ze4X7uoEBli7HnFAPXrZITx
ucuukc20RjGBFsa+Z51A47aPAja3J3FH1U3GF/kYQDzlImunV5JtkQ6MuBkO/beW
iQJmDVqx5G4HJq78T9ngRS6bg2lWKH6/y0//KeWIRzK5JhRNvXNz3Cek2O+4Rtej
W3cIy17aHpXxaazuPfbuZHUm7r8SKm/T2VAneJjJ80llfRx8yNzvMKvvu5F/D7YN
+25xr21jdv9XUDdxyokn7fHogox46O+ju1+QEQSkjmhbkIFkjh++Nnjiwf4RpO6C
F6BQtomG1VD8F+iMmThCUu1dD4DkUqwl747lEzwl2mhTKbPnSBSEFy1Ra7PVwUQm
K0YtRzx8I5IDTgtacCZEkm3GGvBb68jrNwW3iX4PPuqgKjCH0JdyC0S7Anria0i6
ElfElax4xWRNtTzoxeOfkUb/jzo223JFqF3mzzQJNFxeglTpSalulACaMVk3q7r1
CYGzLnOqxt0pfDstCHhljZbRoUa9G39NSJKzqImCG8u6VBj+yQpbtIC1gzsTVqy1
dbgHv4e4oT69SjFNaPZGrwAIFBW+RRceX7dygKjzFjnEq1u92us0i31E+zf/1ts+
nWVBhIUhbwN/CnChhEDD0mBVHqdvRw6CdTyKFzAcoaqOg0tuHyIoUvrspzYRHC+d
RjQqQxBXL9d063mf3aE4vgv7KqoeRBqfKa372YwZGopp8FuZE9Yf3zYbM/lZSvC3
olzijS2NuXphA3jHc7h9+edUSsCEBJ3XeTNpUbdDCot/VebT6FcBVnJ9NIftTmtz
Q3+e+jD0C9+44X7sD3egHHvtKV/f+AFDlibFFW682YL/VAH0nwu9KhXaim9jr4ep
rhSnMeqwc9JSPYfqWza5v4bSXsKXNtRGyxNiyfKHvmoh9tEBNTveJGho5alIBE9p
AdVjPOUW/fpLYWBApZoSYMQSGf3z3XCSDP2bgBISo4HRLxZBzUWJY0FNLA/GVtyT
WJ08tMHWqo7EYfRpEctYM0qyAe6HKrHxrXovk08cseL/IgyMX6tZrDDETQQjWcdi
3vGW1+aAEetyZuth2dAACTurtvWVvNa8qe6wZ5+gZPPiNtJECmkzcl8vdr1ad+Un
Z7RMtHVOxTKIgAdCkbGa0+FACtiHHNAABeSwFNZjee6aBs+xRkwo1SWZJaJu6GnR
UeLOMhjfEqerj35iX13vPAdcIQ3W/Edxin3kh2t8UI/HRXXDxv8hA+dkf+8rIWVK
NTfdDpm29SbB+726yQhEdvkJdfK89sNZJOtLa9GDxblAjpfc0oIC/02dkyKp/NDO
vyDAs45fyQts2t4SSdAvTpldnoCADZFcffr0C9duOtA1E0QUFmgM0FPrjXNRzZc9
R+aYcYGcoul7z1gOznpyIXFEGjuetYYiy021YlmrD+f60tQp2PGkNpR5isScH8H7
WoI7Fy6suSmMklmsLWwDjwMvKFkE7luYG7/HncoWOhb4kwdBNYHhP5dTaqCWI14T
kqBMwYHlq8L0/4ciiTcutkvM3uYF1YIGULxSwQRtVt2g5MkfxkIy0LyQyQOHay10
ffX8I5fTn9hISLM9Q22nMvuigAxGvqbHHtyyzAPOA+R+8UVN9B2BLDr2XLqWob2R
G8qi9FpbBhCNNfEyz/NfQYHLByGH/rr6EE/kZdb9kK3lyJ8GSoUDRkkvGsxDKO9l
TQntkcFYkjO06pu7ConvO2D+L8xu4xcrpJ48C9SmQTwaw29hEnZ/MdFMsGee83Md
c8r3qkpGJFt4LfzIYERCn8pGh1WNGpLhDn3qfrFm6SRlToP/S2psfRZMknXkJTIL
FzfNH83ZwJJbVrZ91ZazCz/pTu/YGYqd+5Fc2TQYmJlU2zNXG3sNogdeArZoMSaz
IMzBjANsad7jIUbhY4hqj2Cn8BBfske7mSVCX3JJiOuuzJ51iKf/xrfE2VlVuKSO
QcPdcAYw5pjfDg7af43iNF6uQ7lGIWEHnS+Knjxwdz6k81ZFF4jruygXRTraXE2+
Exv77zY9eFYFPv2kIEG+GvpQpybFDZKJosnbTZNdKpyM/5fdwbrb2s8PTT8VzlAS
EgBeObTL8eC8SFeBknNWQVAaAkRv8fWd/NKA6a26hPUgDJbUoKnPWmJSOR5/nyt9
iqz8NGE0xtAJB2yqgp4kEt+Eli54u0BzUcZZ9UjHVSPTaeItQNL34Gz9MM7hZDTJ
ZUX8Wrw2kh6op2ENbg+wet7WrXmu00ji8NPBJhY6JH77Tde09X/BkibAnXMrr2eq
OCD7UkLYMFvGzTn63W+KuTA2KD5mC90KCeDnykJL7/LJG1d6uattq4IkWLHTr25x
xbobtGC5z9bSn/tFTR5dq3xZ46Hf139w0zRIIeyF9snqEtMxWrCUbwb5hu2x9MyC
LSUjD4qyBQBN64QR/12hCRaLPIqb1DIyzMRth4H1PLeVERaXe7GBWgMw4NUk5RJF
z8by3ohBpoNknOtpZTU7c3uA3l91rzAcMrusVTS25f7/amFW508oNiJx1NCAXR+2
uS6ZXvgQIw46XJTX5obvdgUmuegF8UsfXpBJ67Fnl0dw7LQblKBHIAQ4x0dwd9t6
ifAA43KbQV/n+vwtTcIw7/htg5Yk/5+oWWYAIG5TMU8cCXoM89CiSanY39scTUMb
+w4eMAM/tE33mKexWOBIqtVDviTHI+zqSX+tEQ2x+NR1F4TQkCo+9JXR/GPYZVlJ
VPnOTqQL7Hr4Dr/+h52+1IKQYyv92OE2/P7AOpPkzTxPWUI/daunkmj3fO9/4Wco
3fWZVJ52Mdx9ZDnS8YR+BbMzoyzhxU2aE4eaqbBklOWVU0KLZlbQnu4AFoZMKSLy
Pd4CtZebadYyzvyGIe593Zr62zFomNpU1llPq3BchT5rOIdejOZspRLMUyjAfYKU
LsQ8VlDhfQIWfizzHGVGx6qB2UyYDcmD33ciuhMKQfkeCjCn0XcMlgUB2ODvoBbC
wscmV4jMGcyHV+Hv6cMMHAhbTLgk7LJ3lF0gWn62BZda9pKVw/aPe3Y3LVgj8Y0w
pp9OhQZeZywCjpTdQvqj8WW6JcLDyK+oEpDVTUZtAJZOBYmRpYhrFBME0q6Yuk+Z
r2Wiaclc7weIvAFBV2ruAeJx8Yj+gJ8zy/8fhY7FjLSKXL1q9z+YiBypRecG/yeS
Wywgt5fBHTg/oPcUHfBJTQBNwLDrmQCOLKKdfSrSxshgP5bEreYSv4KcsVZk+sqZ
vgBqQu9RPUSYjVT4c/x10b+55W0hBByky//X6q2gmOXiXLB/tA3nvBabOnkH4+gk
YPJohByVYJoMSD+xe8uTL656eoYAEnBrrnSNkFOhZGO6IRMy+TPqwnTXCeZmJH/p
S64zg4OST6AtXJqGoZJsmBuARUpnFxTUDmPqxdE0E5az1R4+Lw1FQcnqQC1KooCW
rCmuST45+0Jj6FIgap34ntX8rhL5mOsuXvEpBscv5OscmZrePd1X0SMcqTuDdVsm
rcQvnCvTbjUQL0uYx9Sk2/Rn3Yxt/up2oclBrlqqlXsy7kgTJ+GHR7fXOTU8G9QJ
8RkhUo3/WQ/xK5yPfe8M1gRirUmbaCeJnbE8B6fhFizYUsagEIjRR/v0peyQaYk2
Du3JM73P0GF63uwD/44WrP1SzRqUWyaVo8CiAxue2HnJ4d0nSuo0l0zmhi4rYr6k
GnNtbTltZMotknw3YR2ES2xXNcqX/iwcsGm3kBjqfVbAAWNvpofN04OMzqMn7F/d
UjCeseQUqZtIPz7JN7h5+uX6PJKMhOmh8QiQKjdKSmW713HZIh3vHIx+5+8VaS59
Kqukm/pJzPt4XbIwkUeO/W2H2ZYW9UHrt303sfC/PEUOI+MWKU03ApAE6M3WLQcT
HefmiDQ2Yj/xuRlw1W7wTWImNlScBejM5NkbilLmmJePo36Y0EIo8ltvbLFQi/dq
0vSN4IFAcYwkq5f/IxN8V7fdcMi2pMxIMKS1GxEv0OefwmQyC4eIKd29Hcy8/YJm
+zT6CfMsv6ISON6SgV8D1OIBHmCmC8W1n4183qcHIbwnBRPUbmvBiLNpHnsY7qz6
Xmu0FPzr5KtxLKyqhpXs0sz9rKQ2wZpXcubJvmDMsqs8HP1NlTVyLq/R72/d8F+G
`protect END_PROTECTED
