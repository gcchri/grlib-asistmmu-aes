`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6gihPvFCNeg6BhHezpGz9LIL5xBzQEElTPGZrZy4L2+N5nFVRueUAX/S6T7HX9Z
ux2USjFiFrVtgMrNY5VWU7IBE4kAhC9p5Iidj6JwloCekEcUYMK5rO3S4qRP74F+
sN5+9wB0lu24HC1T9rBKDhK18MHPgCSKob+GoTE2JZUvr5CAASNylv1E+FDkZysV
fMX+RW9qEtcLOIcHCQCnApQ5JZ+17zuLSVFdYBtadTPpWj2X0LebRbmkdS54ybPW
oOUbGzmGMPq8QYe0M20Ptk3ig3Z85fR9F8Qb2j0U+2op6NXZMjdOxjV5YJTN5U3N
a/R/yFHxTMFz6TG2IL83+IQ3SRELqoc4Wk/7Oc0waKJlv3ITtDZDaxMtNWGdcn1n
5ycQRj296M5466PKMOmgzilmWkVXN5HZ3X763GxtV16rfdF7LiPmQeqtdLF9jWWg
9w2JblXUImX3QeU8gX6y6ZmGUpgWbG96mQrjaCRnnssccKjOi4lBELevmi5YV0gF
WG1T3lT4gocTd+qqYavrhjX6OEXJA6Vde3rac+YROVoCB6sw5xBeXXN8wo++ZNAu
7BcpGMO3T0yZrnAN7PlKDnlitINCpjE9Mrdopc4gWTaOMZumUxJxS+6Q33CGphC5
gKBebk444lvYLUbsj+ZRS6+o4trUqVQe/uZu0FT10Oe40XtKVn87qoKNUW/lEw4e
FcAH890AJ05mTs9deSI/Xf+AelSOI7ZSIdiuPZpYFNalQnYC2SBYmOYxTU6MU63S
fw0YC4EchSIghdeBDn3aNvQPnm00gY/b7FYQm/F5k0tCrCtiIlPUmr6/cEMBT/90
PgbSCl2H6bl4EJ/77RmM2RkldFfMuVgxyFFqKAQlUsjnGEIogwCyH8POr1ilpoZc
7QuWQ1tRrugw+DQNhQTN/q6kanJv2SEnYactlwqum6eGanzEbTCOSgb6M1n+WvBh
FOceS0CTu/1y69SGBCFTcDVebFHyVTQ/kYdI0GVoP3l70t3Yw6tAmbc71XeWagEk
SjbKblUmvUt9RjSGB9QGT5iw2HzlVl1nu/iPnGnqe0hAQ821O/Q9WpCK0WYUTjW/
/52mPog1BJLIl6WDAqs3LhoEVqGgTvUaPXg47rNdoFnvbBpoaRTc1o+fIx/K1ggf
/d/P6y/OXh6CLEMl0uy0a6VkBMun2EzQ9gezxhIrksw2oFr61C2HV8oUWMW+s7y0
Bl3D7amS75Y9JLTPGxhKv7ftTe3jMq1P/4a9VAYsK4Kar1bq5B7//Idy5dFs9dEd
z4djRgefJfBahVTkKjhUChvw84nE/sFJYLqdfCQi916H0CGwhMFoSLFg/ntN6g2U
rc6lzO1uLOheZ6kQiiJvctTroir1UTN6A4u/nDdxCszZ7pL+FP7SAgcpNHOP+NAR
`protect END_PROTECTED
