`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHxfhVC914TSycHztvH+sRMsIxz/ItLS6b9YiJNNSI0c239ehl9oQUpvgP52Ltsn
eXEIgMPlTnVrL7P7to1OabnYMy3L7CY8qlLekLNRji8ABdX2Nkm+tP57xgdHD0zp
2muyvGGJDIXlLxjwUjTX/JPqxH8pppttLbR3K9sM/mTEgvz6o0n65bwS/NUPhWHi
i79K13u7yvpi3CL5tXfqy7EyXOA4L1B9hzD+KfcUswBJXKs/xC9tDSYW/7qyGipZ
Mp6hTk/q0rD6T4jClVP7LiXESJzhReGPip/wGiTC8k2InTG2Oh0dvwF+0iJSW4V9
eRlP4Am1xJ/LIY0pFULkAbMJhzbVbC6OaOL5lP4WkFf1VxYhCR7U4bnl5gbPUwGN
dnMvC/c3Dw3q9V+bZFj4lfQkpnnhbUobIB4gYoNVKxxHc/yDKOgBkDpra76N9XmR
yFM86Hl0KB+shws68SBuOeazGMuuFAiZKbx8oDWBOYr6m7LA1uTgiuaJ3yDMa4tn
DQ8+/Sh/hiofdc9IcA7GZYZI3I6BAY/qDkQJDRMVhQs=
`protect END_PROTECTED
