`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q08eC0Pshx/LpQHn4E4XfNcegtXrTQ8WeyAmEFdiKW5LOsudiHG/s9zV9DWkWQ7w
yMSNn8YYpG9vCxolYpEvrtrdp6bR6DzSZGVIQ+Hb2hZmjDXxqMwzSYlcBR5fhQuy
K0cK/OOTvVRHuWG33rbkie06tAyLIUHOtfGCDfYDXgWiecfISjE8nIspwslPfUtX
c/G+MR+XuIhaw3/ucI9TKYUnj0ooSejJIqGjc66mHZjyTzmcu4eB2revTJo5BjBq
Fxrlqpumoi9h81WE9pTeNklIcsSHvBNBXsHiqkM1kILwwgcGvYdjUNBqSz24MPyJ
4GlYW/Wf1xCS1Q0GoUsacvKhjfbp0aga/CZLySUOy7gfgZM+Cl7YQ3dx3cVmLgz5
GJuHl+DL+8Mj4EqZtVJtTnAyGx8QwjBBSuo/FYpfzsvCdZGkTTHwJdg3n+kY45Bk
HyKvVGdrj84rm2TVtFEBSdql77wKMjS0DN8hf5Q/4WD7e+QKZZSmU7zZkN49+MpI
ITFHNhIybZq9VpTexIeOwiWrYNO4NOUwOMpUI+wIBniPP/fR1PPjiGSUGXWZEsrn
GfwU1wozfUmyHJ0cqB9KVOG5w5lq2y4WbljzieAxRt8MO/h3NhPAc38ieBfQY8jr
7TVmWsWpu5oZVVjA3eLo3Q==
`protect END_PROTECTED
