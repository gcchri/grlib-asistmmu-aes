`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zosLzTPH2ZSwhuIlAjMHyAIbJj8+sETe0P8H2mv1c/g6Wc2P5rCqiJ60USUTjK+s
H/nshr/56SfvGB4laAPGWPUdSG1Kr0dZANntWgcjWkterBl3ithbd1LMZnxa1mv0
i5tDQ0HQXZFfgccblwjeC0p3hr6mjiHFFgFbOXQT2vtDPJwWLdd6m+D5hIJNxzAZ
SqtCGdqzgU9Yrp89UjDoAmYgp+TubSDilwDAnzt7Zm+8iOjv3PIihoju4hMKrW27
KrxhK5z9cZWf6YrWoSOGL5McYbLG0k7xk0Drd4WJ5Zl45bTlO/nVHU6vBYeFfCeC
MBRbqRQkw5I6Z62ZmvD01jJMHEi4rdGO6q5m0ZQ7qnFB62OzuT0qr0fTQpGC8Odr
nY6K8VBJiBkM2N1Rolp+k2z9QGgW0Vw4irePwObxKQF+1gERVvCo17pIzk0qxpnp
8g/5O0vJZSgk3HlqfzBVQ86EsN9uyO+t7aOBWq58ymjiCbBZr13zjXRLAK3h3XmU
V6xaoqI2Cuq7E0QoqcDS8Dn1KODJUFvou0Gzz43geV4nKpO2UHt56EZNVBihurci
hJQycQczGywJLQSYrt86++TtmFteRdWeo3UqxnCexfOlctGR2iWEOc+VJHW6ftPl
u1SyzBpjiATi3oJbInO6ePULwoTL0SV9c255HZPSsPY0hdbX/yFoGSR87XiG80b6
HYwWCAWyoV//rgwfQ+MX0R2NxzoqXiHtLUKKmdMwGk0LZfkhcCJg7ynxIYfwlp1s
FyIJfLwmppKLb7b2p0r1JZnImhRbt6iknrEmMqh0nL0V5p7quxo/6ueYIR6jxSmK
bdKBidCon7YzE5BDGa0NziUn+Jqw52IabxLGeEBsEOpmMuEJ4/eTThSZRxKdfeoE
9kfeYRWuKOHSBE0RA9OfEwB9O18r4B1OWHNJDatSUOSokKlm8ZZ9yHwoT5U/ohLH
J483p9lO8QDs5M/Ulr2NC6SkDewfiJuQyQINNfqSYA6LSgyB2KSIs36Wox6EztZv
Jg/y0DL2HwNHt2+2q1Oro0QcytuOLU64L/5yX0R+ksrz48kWpUCJFKQ13oUoM6/7
idn7VvhoRDFoYb0VoNTI2Q9gpK2JiWAoCjz1ST/A2Ode2JTvjwvZH9kwJHRji43W
RaHRv7sYGGcFMpv0mQn5lJXo4cKLC/3xbdP6+lKrGX23faYgSfXMShFJsEnEeLfk
ihXuHzqyGZs4zF5zs85TGA5RNm4I/beaXeyHgEylY5OnfZfX4t0lx6GdC1tV2GOg
K+u27EW4W4wxXXV2ex1+IM3wGzJg9EvTitgv3soJugnm8lNLH/Mo9ynDfqeRD5b8
bbZc8atmSmnQFzl+mRkYHRCxl4+h/2GsLAUYlUkgrdcGCMauzy65ou71jmF6ud9w
`protect END_PROTECTED
