`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PMKqaX4Smpm0VgruGKStV51F3vQmvODfYDAognbo7308THHF7XzGZRPSO0Y1Txl3
FHMKUoMnPVGfu8JRWwSijTJJnJIMV5cNIpaDpC29TCXTUOp6PLNeiMNArw4tDV4P
pmWT58iwTX6dqPSLh3qSwA8bfY+lGmoCt0AofOGYWK01vd4oZ6TF+Rxb8urDGEvj
Bamob5XFCfvyD10DDC/H1/shPVrUm6xMiPX3C0LyDnmgfj8bX6rk5SPm/SHuOQ1o
QQ6JWwO0KshjQvNYWxi+GGAPPGupCr1yVi+D8/pTUpwdhX0zPKBDAKIzsdsnhORy
zxom+Vq2TzII8kC6aRN3/yXpJAz3ii33xCOwP8Ndr2jClK8inuV7JGA60tFaskkY
obnXwZP/7h2FrXHA5DFbGgOMIwBGCRnPbpphhRPn8eQQMCVCkJ16/EEh20TZhx9V
ZZxeRpHVcgZvQAMBezxznr2x3QPUfdwvUNpoW6aZ0VzTm8x8LaV+hoVwd6yuk9WR
`protect END_PROTECTED
