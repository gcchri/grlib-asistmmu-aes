`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgyIbFCsYrAFhBDqbuztHkgKAEnUG9n/IL9h1CM7F9O1+li2k7OL5fQFJx1RAQ9y
Dm6IzsizkOzOryd93LggCpMEwW4vfZafm1Z+LWlVsQVaxtPxHPieVPTG8TrEoZYF
ED7o9786m80zlPLx48ks0yAezXi2+rPaqgaHFwdzfN+EA2eWQ89UAB9KmSNVrDuM
yaSxKvPuJ8F9JJzrfefA2yhsnd7HATDGs3j8iEw43pu4N+oYRxXQFae4Byc76TtV
HjfuKXAvhbYpeDUGduYcV6ZqcKXj2GLd/+Ryci8W4dUIdga4AEEP8QZhegX7yjGK
B1OWUJFOSoEWlp0HfO+K+GWuhM/Mn9toDh9qFMTaJZZScTyu25rA2UFQIQokXIyN
Yoxi6I5hsRaMXDBBRNLrkYDA3jmZZKlFjzRG969LAZ7fxURI5NlZgnvrWOo/Pds0
m+NaUeT3tyMPKWNwuHuW7Z7ICU8alvhrPUzDrOADhkBfFh3qj8z4HyugyRi7/pRY
YGe/XpnZLjeX91owh/B3dku8JJacTzyrB5PcN7WZsYCin/NT64QAZSCKRYy5FAq+
RBWT5nXSWZayb8oZW4JHSuUu0HerbeWt6dHS5wxK2aVPXHBNuDSea6Dpc9WsAetN
s1daZDnmMWLiTmSzv2i41JtPmlZLUscsZO3lg+//VfaHF4gIc8Du+QMTP255hfdR
YuA3jk2MaQI/iWVJkAbI8t+jf4HkIx098f+G3tpRTf+rWNV/3mWMh5dbpFjmeead
H6dFucswogXy+5C/iTm2aSdrYmjdNSiuvpMpnn3TwNCNBB94qRiJE6HC4+rukIxh
r5cBGRcEG6y6oe/WxO98/uHj3j8g4aHiYPE6ZWTnD+paZC1UIrI2j2oGs8/WgG2F
N+8FSwrJ96OsHTpvQQV3LPLX9Ft3rSSiqeeakMaN50k1rMCPrsUa22V64c7dICYh
TQ+GSWrqJG9RbmDUrVHZvwbO1sMSmbrgql/+YyANTpdmWgH2kLjmPynwFpGTyZiw
yu0Fyr8ViPMm7/2DGmlMn2Jd1QrGNhYZG183yFPwzTtwK1mo5OFtkq0TTD3KgVu1
1JBqlPlJ9B5p0d2f9ftSDMVUeMSv1o46enqDnDOB5Xa/ijcOecSrnfn5eZUy5uEU
d9+uqrgCA2ITxawEGqTDJLrZ6UEDy/OahqzGUR3thuuV3UVLa8Nn1rG/G+i8CxdQ
mfYxea2E0dt1cbZeFgQ1mwNpQ8dByK7LjSfEM945Gc/+iDlMwIKDBvDUXObIU9oZ
DcEd8iBEF/kgTss83mkFRQPgXcX9ZDm/C0JMlnsBJAMTt3eo4ixdRFK8QLbGmoAU
SEU1OP3Yx4Xgol3vWwQyemJshV0W+6AAGviA9WY1rJJ/oo2YlMwWfmXoU7GD8Dlk
UGfPGbJGb0Do9ZnUBDGo3Q==
`protect END_PROTECTED
