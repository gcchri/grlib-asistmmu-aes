`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Vxh2kdCnQlwCZd9Jy983FCSRCOCpij2s0RtX2WXIFujzKLKjF/ynO5eyqKpSzFc
0WKnpUxWyq1H/NfJrYCwml42gnHkXEMJDKTwcKXokUTetKZ1uVrO0e3dEmfZ1Yb2
8ACDXa0VvXnRvOxeeUWgrmFobxDKMkH7dME/dTmMGa2EswNf/kletdp2fpMmU9FL
fcfx20BN11c9tiQKFxvL9thFK/o9t/U79RsspEuTsvVA09dOBFaZYqrGhtP+c5PK
btLA6tcrLQ2JNGF/026fMVscOcQWaOuJUBg+zjdUXeGF+Be6bVG41KktZsDeaSFc
EmC4LkQYvEDZRGJCTlomBP38tOiPwCC1S1dtmuimkuh0aP1uA+ZWcHp5RhydzDR9
rqSEKahZWt61EQI3YjcCO6Cu+u70vr8MP9l1MXN0rTAmiOtWkWiW9wWHbmtZt+EJ
`protect END_PROTECTED
