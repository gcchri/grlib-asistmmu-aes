`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EHczp61w2jVwVUQIT9lRybrhEL2Hfcr4wszFsz9uLd4aveG68HNHLwzkCetUu1TS
t4P6cPjBKVh7/+uNtqp14LZEm/F+TJxLnS/bKToqVvf5DECLIAR6D3sZ6yK4dcUp
V5Nn6wFt8EDntk/IoxRg3UsJJDeph/oB8eAQjAU9dWKjZ4v/pDpFrwqhlsOQ1MrX
8MsVd/f5pBVacmorJGQQuZkrhlsUcTEu8TwlU3amviSe59sKvGEcswOVUv1XtqMt
4yBVyl3xEHTSHFmDPQVTFk2jzJGMD4yM/ywQ7LakUV9FD84o9zgy0D9ECOc9Vche
2LUvVRSrM9JQxCt5QCLnN23eUFgYbQlvcVovu65zy62hoTZ8g7IB2NsrtjHT25DI
afXmfeAMAyoEAdrcyVx7MFRB3dLVUXotpGCSFLIpyy52dggwGIzXXrAybcYxXD3o
qa/hYVj5hlavectCnrvqZg+qRMOmAx/wP1v+Mg6mzmJTak0tCDbLeGyYse+eTVWW
UMRILKVsfZV/0szuArUob/phttUS+SDduaVCUbGFPZ3LadW8diCr3fkjcijsi95a
Kqzpuk041TUbMJ7TXdo7EOkYtjpPA1MepuMzgA17rWvw+9JW0vo9+3L7YbCCGN1Q
Kc0p8Z1yLnH2QEQYzO8yaJn17IH+ScHBTJ7imxSvgVRBmWs0MODBi+nwSSxKrDBc
u6cZ1MXLkY5MGypx4Gpke3q+9cXmgcDzVqJqUIFMu032ZSpTHgXtYPhthFnQTGfF
g17d2RBHqJxvBqz9HZxJzHDkgXYI/+F104MXAJPEKWQnTuD40Bn4sDFLnhxxxEQF
vljbaqUxWrz8wOCLLTzv9I1zZ/mcWoIZcPtEAkgRqIaMpP8NlK6bFAYNiEv6KceP
qFAtiL2Uowl8CSctXy3XNzvw6G3JDbRegy6gVgPQ+iEdVuj/LnDrihelB4pEFnxW
0xqqARXd1R1GCxBTJl4RKK9uRHnNoDr6TxcF5kXsnlUy9MX9C6yH6sm0FRKs94qQ
wmSooYDf3qE/bjvcLROH7RGF+fzlxopuuQ0sBRe/9VnZTs3NgTzeapNdap/N04TB
xOQJ6nzzIlXbrDCvgs9db3LY7dpzQv5bZ6zcBaqYM/9YEDrgD8vzanBtYh9WOiuT
iCZAfjFgBZPHHyRRtFEscUmSa2oJWhyPBM4kmwvxoFxLdMmOOFX76P+u4q4puyxa
IbsJvGXJRU7vr1W7O/ro2PS3dxNN3jFrRGnv9mBGM3Iwz2rZ7w4KBD3WVIsVpbJt
ipgrUcvQg+cOJNSL7klWA0q902+6rXROt6FD03FGK/ZxOdlz07llcWmDwrXXY8bC
//fxriSchPYl0hnBEXViXCDthYwqCr65PuXm7blgQu2V9B8zw+yFANTuvWIHGeHw
oEihCRpgloO235O64bfW7vSBDH9mG2vQcMDE9WYqLgJbrtNFvenTmPTPwU/sIfKx
nwMXwJDisgQCcWgNk4flblserT9g0us9YVlpeoeGygMD7aR6jmtxTI2PKKWA0XgJ
VopS2gDSeLPlglVSbEK394KiKcCNUqS7ej9V34nhm9b7JyQPlaVGf52TaWdLFDWI
1sYuFBKJ8xlls4lOe7ceCFmcdITbWgxrwdgUYgpAzf4gwS2Z9ZNg+uoi/1Fs9dVl
5cYlNQKy1ep+b0NZRTkmKQJJWjx8YSxpDq/q0P2HBjqxCfzEPYDp9r5oPtZEWH0n
VwbykB/0s+iKYKA2DzQn2nXeMDM1TaoVAIwWij94Q1OdkbhLkKoxaHZr+YtOFrVK
rftGnKp506VESpK58XbOu2vwg4P6rokHsVaj5SFoun4/ulkzvq4LRIwL10Jy2Pm8
nZQFMSKYKO4HuuM0obZsEzgHxhozr/MLIfwFH5BQsVY4chzf5t78lI/wLcF2kDpu
2i+pdYyyolOiv4hibUPiyiWYt2zWUhPQgFjIcmbItR8l1QKY31W7KPTQy4bABepn
GmAEzjn3Qd11fk+x8imYkK4bC4adhmGv73T88t6UvLIfU+7eCA/yIs3WyDGV6Rrp
0ecWGOb0THNjKZaJzMeKTleDdIkrfnVubIr7VMiZYh8=
`protect END_PROTECTED
