`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QPqJskpRH0EV8U9BACz0ZR5vHfu4XOdFT6y7aGLGvtSE5KTdtM+wj40OigEAzUvc
IiPRvNz0a0x45FvdmtQcEtFHoArzlTfmPPUJuh4jyzfVjJse5Br7GBOk3++0Xbdt
hFLjvSfAWIrZHvwldPhWT810EzwijHQZCHBJ787rxUMnVk/9PWy4sqybq4k9SFAb
ZDQheHsG6rn+aE2FdTxHCIn0QdLOknZKGlmb4S8Ta/VLxJ49nsHdftVgJuH2qCha
DtOO60wUGw5KlPAGjCqClhXzE/AnlIiFfyVhT7G4nXOFfzmRQD1OeQsItEo1qph4
FBwCbrwg6NjLsFY79gUVUyQkp0QUwcPnXkwBOo3LjcXrwKDfZJNfk5IJ8gUZUiE6
FKCsCNPLl+tTvpBiDongtf68IUyCnwqfv3UNh5Ql40ZBWQH0WxbZdydenb8L7pJL
`protect END_PROTECTED
