`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CFVWAoqZ4LoYG3v955oU5Mo5a5/97uQ7BTbwyVuoo/uJBazZxwZMREz89NLjH6ai
I4qc3BKk220kLM+VkIeVydvpj0FoLds+VlnFEgkyCa0QzeYeUeS29XQ5IiHUwQKD
6Fu05Lk92jic4f2c9fQUCuqG/uuyXURRYjFJWATycnuUx7GdjPnMNK0GmTkqIF12
5E/R/URn4mdeWVPA2/YlTkZih8bIAnAZMDVDpHxd2vX65wr1Dhn+pLDBca4WWh4h
03Nd7+dboYrEl4r9wrRV6gPKtZkzd4T70aO7bXHd8mr4CSK7EFjiPo2+fIPSSvpf
vtEKQCkJAl68OCpXpwnqWO8W7Mz/SnsWVi9D5jujWoeo4XqoDFOYXgIFFqSRjLRg
IiCW4Sh6aetWcc8YO65QynmY0HCyNHHhVjsilsWuTB65u9QYnBLHVILCn+M8nMVI
GS/BnRVkbLd04iKP15eNp8YS8KxG8jPGTKzrzAK2DfA5w9//SdM2gw28Vl6hJxSv
+jGVnPG7KCFYSprSwy0rgoJGRrESvqYKTZHjHQnWQNRSxuyuDqHWGlRfA0QNOEaM
CvMdnFIFZFAgOlNTIxug9KJ+jLQT9Ugco0K14jmi+L9rR7vr+Ob9PuJYP0a2K3i1
+bVjMnOieTmBzg7anAYTqHu4uHlxLwEQh6kFnkGUAwupFjvruZvCAOXzu8WpCA91
zEBFFONYpilCZwBG0CncEsDWBu1Ec62Dkim02wftNc3rbFY2GAiAZrp6HA8gNBDX
BHg103nkfutZg4FCgRuZXlsAf9FGtYF9Uv1uJj8AiAD0jFP8T2GeoVaVZdPMDJ/m
uL7ylfXPheAi5Q+Q0nIHXYEmUJy4QIlxUz2fjVWqzuCVdm0R1Jljq1YdifrAnCp4
KIXSVpysr9QP1WVdFE6WXRYMFEWG4dyMvq/8lUQkNxPergxBi7ha0PsA0CtKRlmh
5KajAXLcwNAsvZFUzayYguLJPSdBNzelZOvqDmLCn4BH3GVLPUTb7OUEuySM8GDN
`protect END_PROTECTED
