`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jnxV7Q9v/wOwiuTHh8l+gZ0uAroMp3HruYCy6xAwvueyLSwPDNIuq8xa0dT8YGFb
cS2AjngYzagvGEltCSNDVdMFh29vx+kCP0Zcu/Mm0z7sE/EEmAhkk2LjiUdURRIi
b7V7NkCcJEFRd35o0tGr2ui47C9ncA/3sC/3ktdxhyNPndepZLuWB0ijCtm/WxsN
b9AmbHrUJobTacnUG62U9NKh61RtfJTlbA+0Q/q2yOeDfApA5giGltaYoQGEBtUT
+exFA50AWPnVZeWVdi7RD7a5+9hmzsoel3y2rNn7luWKxiC4mJ/JnZ2TBMvgplzb
3cc7uyJBTi5Onop0SR4TiyQ96iszc6FvRUFT1WPnvCVzflgd7C8ml+J8b4j0oueU
r10B/EHbb1Ap2GQbybBIgJNR1QNaKkyqJjBoXpEQDUfsGvpx4OoFU9jOygnhpuWQ
NLvKpU3Ma9sOfoqbdoieSmrV4XE+0z0XiCa4+pdSCAHwOeF3DqU3NnLtJmF62rUm
`protect END_PROTECTED
