`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmJZ/xwXul0Z0D3VWVXe99mvhk9TU5aeVmGE8Zc1sPRhQ8/oCZGH1Ma8JCUxAhGW
zvXjjCOIaaxYKAm9/7DGkvpC8JpA5ENq7yrJR1C58nN6cEsCcMQxOjRjInZWdLUy
o1fgvxMr6HHJ51Lr9IUa2NYnaANdJc3wd1LIK0O5B97/r9RabCxeQX2Tc5dWFFpQ
WwOABJygJHN1sIyMX6leAuFbYYU7rywboiGHYOgsXAEYasH3ZlOCkGLibLz+MhP/
jMg+pg0ty8323kHEVW1HP/MB7T7TV73B0jMEGDF43z6+nBkC2NkXMEuYxMxMqm6g
Yrsnri/05+5to6HVJesjr2eCAOpLneigHx2tNv0YaClHMHpG8OdnhoFGlZcJJiLn
QjqlG4HA352dFwbb6aFGiixX1zSeHbMxo1PcRrRh5rpJyylNpLYwNkk2sNOqArDj
vFuoL1P70lj38mPJI27XlCJ78VGd+hziefZJFp+QdlhNwUo12gVyAQdDjEUjDHtL
`protect END_PROTECTED
