`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zqx8Sw8seXi7HRAf4+vbDknk4kC62MB/E/nC2eiThKP/dzY5FaR43ZRbi/oIm7pK
o/5sBdTLDHBYsxeqGNCOZu1eovI7wB+jY6rIGt3vJPDYbifbmj/7TMwQyParqoxo
Zel62KfR+9/4ozKkO1UCAyTmdha3Q1kjsQdcLej6Mx+idibfJnLnJ5NLq1jGXLRd
oEyFq5XBykrWplETO4cJA1qLvcCSm0oH5pykohdHzXnQOy6sPrYtVZmqLfCN6Y1I
vQltdHwSkyOv8vncpbqFLoGv0s5yqx7T7I49Tu7SMajdcK7Q2dqpzs4sZJaOe5EB
EjmvqFMO+4ED/QxuxgebYsUhiAuaArYsiDW5MWFxJj1mNZ6JCU/SuHwLn46fm+OL
ak8L9L6fJxxn15d1WXGpq7intwDTJ60JiFC29hzKoOh9wd6g29fFtC5vY4ryoU/d
3q/BLtk2DPGdGUmf1ukLWlJmXx0I6ydG8WM5ulvRTYQFQNTKRyoIQz9/VRdaGtKy
`protect END_PROTECTED
