`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6N0fKRKx1mxHhz9VC5hbgIHge0Fphgcej1iyy7u3Ooq00TrZa0aYYOqj/iGS5v+H
EHB5Fv24pjIEbOzGu2O4Ki9kmt5ZFax/6r4fYMk0ClbF81PaztKmiTfRsjjGWCTs
X5tX3ONwgZ8cuLoGLXq1cFOXZ49pOU8I3MF6v5nhC/Gxh4t3jzrJSnTvnlfjdW/1
bphHDr9Vpn+mlPbqglNaDQqYDEJE09XsPYQyTWNamVfX9fj2JsF2nxp7yczSrHU7
mZORJC1xUlXmXW9fv1ooyokMm7tlFBKjPJ9YNYfVeER5Bt0qBuYDDz9a+JiERLmU
mkBTNx7avkytnjgDvMtqTZFSYOwOdOl3j/4seul4SkUQ4EYusabs830xGEjMyATK
Ps2rxZuUbUEEzHnz8c3OWg==
`protect END_PROTECTED
