`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4vQgTPBoc6g9+rK4MT4zlrE4OSOgUL8+jzE5Ifv3ziQPCjk9VSu7qO2FQJVm0Usy
7bMySTVEQnpnZ7phwx3632Oz4+hQ/ZKA7dYVgNCnLZKlv3EKkJlRjfWXLPVCSQVa
M+6e34bqMHkf1UgqbhXsbUhwLjYc81jc3kvRPiRGttQBpV/0gQ/CG7nM3ZN/JNAw
LfecySs7+6voeBclBGl4dw5zZvmuT0HRmKx68yYO8iIvqbCQxBjVf5qotnyzfA7b
`protect END_PROTECTED
