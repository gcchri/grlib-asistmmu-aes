`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrZawbsdsH/RtTIZm4Lmm+p4zAjuHhei+IAPW83X5yHTiWFsrl3yHREfpObs4blI
3S4N3JePugIr1QoujCBTU7W6oEvtHi38nFgFIoQhhtHitN1PLDVQo9sKHK4HdoCj
AaCNIVFj9VQ3gPhuIDWmiRJgE49hjqXbaOSvANSE07zQPYAhphhhRihtEqiWVUMp
iwS6+RUf94+pmSSOhLU/+V+KWjbs4VWzRugO/4AQ4yTD36fQi+YOMBXWcK7eAOHm
hK5I+Sm8mNQKu9VSL+pLg9HThop6NY3psp+i3DpYvLubVliE00zbfp5EIquqNeWg
b0C/MmwApGtgzZsd2dEEp9fvppPEqxGN1CK1ULrDR7RCgPrX7yYNotYsC3XIHKWM
meh12XaBq2XiTzBF62G7robidi+vduPfj+OAhDwTWkiR9w5QNEgoLtdGz0xxGVtB
zIFm6SWnjc7xs9sztYP9RVR1pjY4RSA7cC8l2zt9x8nnGIEk5m3JmKOxYKz7aRJ7
zX7AB8fnmCkEDIrC2k/LpSB2hN0yWvsfoZDFxAlalIYMe6VKFSAcmNtzWbOQ8ccW
paHh6UyWPRS2OMPl5ZCAe5sGUasKphDO2hGOFk0xM8PpfGB0Tqcz/c/SZeJtw+Xx
mZksh7CaZTeallN1l+WQEc6ARFnK8G/WjCSs6rbhB7Y23BZls8+2IG7lDxVyGMbW
Mu2kmurb9vupoSmmjLg/SsYeYGeieODCxw5O3iSISuOvrFQAKwY9Ji2ubYcVx6TI
6ERwcsoC6NZ0u6CEh8uWXABcG4Ru7oE5R85sjmhLQUtWOVg3Q59itnumHEYcL53/
sxb5zRIHiS2/FblkYgFgmIIWCndezvWjeDwxsI98Ppxz5WnXLtoLEbTB/vOmAX0s
RMK3QlMGDwXDGRTYzakwIq+AQDPOeseDHufongyRj6RrC/3gR3Auz3CJGInewFJM
xEevr6WZjaRy4kXCEPhCIakrpRUg1WWBiQve0EtkZrQAS1WuTxklWicCX/M920Me
850cla7ZSh01YRNrlha67yCSbqZLVX9FK6CwPownOGXidxGV+4Au5+lpAv6VKMcE
spcn9HIAA8Hk+9Zfqc0xLb9LAxSntBVVI/3vEIx4ejKgnFYGGYN7E6vzfgaf9eNC
T/krQHsJhMjzcq7tRtDv2+CApSF7COG3DRrrimTOwPjdO+LuAa1cwoOF6wv9NEWy
PB0X/91t45JbfstyhMDSPbliCNR2uwwl/emqH6kFtzSuFr1cM5FoIVMpnl+oDsPA
mFW3PUyKPUGDPc4R6xOPt5flnsKbPa2if6ZV4Q/qFV/xf5bKlUPr+JV4VZ8d/zcm
qy1Us9IBDZgySEKg9C5rCM1QzaRuM3YHhqpliaaQFkU93PKN05aIXFPU2ovZMwtr
7TcG64dhpUhbld+lOC9K4ga/lqAkpZqsy+MldvfuvrSOhD20/7EUE6544CYZ28Wx
3siupz/f3dM6/OScw8eVdP16CC17GFDuFlpcb2g+3kCfHdy0ZIF04CcX7b37lO4r
y1MpgEWfzx7MBq35iwW4cN/K8I/CR3K15g//aJaTnilNPx+g1houxv5c21IC57VS
l+zxFgOg539hNiRZEWUUciL1FNuIRntlpkGYGzJhK1/IG3PsMnl+rUCSgq0gbefm
f278bR2nPmtD3YiRPOegadClR3Od++nZlO+yVzry1X4cqyhud/Qxa8d3tms9xr5A
aFaBlnal+3PiPa/HyFs7y2s0RSVr/yabOzGQ7/8Dt4zm8P3CXRTvRgtjnUXFeW32
qaEgIf9UsjV6YBWId88lLsF2066iDfNsKokEFcwPWoCX8DNnxpzS67UQyag2O3tL
elT7vYW1/CDXdFmNd48XlF+r5npbHHAu9I7J9Jd8AyrTXPW9PjPyVvMBpXcOVps+
9eiG/fISiDyz0hAMeCy89QX/mMCvV6mJZi23cHcKdjAdmtmfBq6YGvI2eYBVhYvm
489NHy0mrodainvVcqNjNwz5TCjHY2+2e9SVGD/gSRYLhffPojCk6Zt44P1+j7VA
w6yqNzqCDNEnzSg25wiQraHwPSmL2hngxEUKw/of7178Q/q5HPdVSShL5N+dpwRY
9AkSNFFOTh3a+wxaZaD0kRZRHUmFSvlARsGkiQ6D8K0JUwdBs2lbqsGNsW5+GKSn
t4Ny3QQXS+/R7qcBuI21OzrL3MCPRUyqJNJvKZhc7Hju1aHjQHMmWejvXqPgPVIc
J0OBNeyPks1/l8PS1QJ2SXBUkHyR0x5JnCci3ReBCcH424u+7rtQcMAzMZ1K6Y4q
Yn8FequzK0GerexJ01qJi08Dd30M4+XofVihoc/LsoJ9mA7WaVNgoDk8Ad5Y2auv
DtOzTL8kQ3FWWCrsUDwAajAPkah37DEvgKm/ebGrkOgYQg+1s3Be/ITV8Rzu1z6k
wRQENd42PWBDY9YcDT20XC+/r8OsTnJkuv+ZKLCdymImr4V59AUt+stptgMwyplH
ELZblHxun2mePypBYAWH2JbN83KOrIKlRUXCbLXVdhM5TkY3sCNmUSZEq1rbsOMT
XloLmutoP2pwfK9HNTIkJ1tp/fB1z7Lt74sqCT9Fu+pHoN5R9axr0mkSbKcv8Bg9
mJ5hD722DkZi9Dxz/Ck88Ag7WTtv+22oZYMKlzcQk2Or05QEKdaldjXIJ1FW7Qph
nptgbT947leLAww6uWb4GDznr9uxHDHHPd9hNoVbhnf3Fey521cOHjOPWbE+YXOP
Eymqga5tvviqFRHa30/SxnvsHA9h3NtdhCGBRyfscCa1WnV6s/wlv1HYr88kHsTj
y3xkKpG5UIAbt8SJ8WRx1yp8ChtfLvJe/hxuM1v7839DI0Isbxiy6uiVfttZqaZl
LIGEDphEEiBe7qqwSqWj36HXDaXu97nUxwFuZBCe+em4qH3wVJr81GceYwtQ02ub
ydeZtxGq4QckUuavefWPpg==
`protect END_PROTECTED
