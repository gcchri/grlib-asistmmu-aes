`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+dqw37Os0kBMiRYbxv0VvoqQSwAXYbHu4SlRhJadedh2QLYsanLRp/+gwMi90dC
9NmXKCh7bDhY1LVNVeRCOm8jNNoxwN/o3/fq5ofnb3Fm+eeHdNVpC3ChOhYGzQ9l
/dKDkphMkyzmw7a2ED/EgMK1z27VxquiiSvLa+kUOEJAWdnFvsZ1kgjbD/57Nwxw
hKhaVFnNZLEg5275tsOcR3DFJFZwtOFfh3CecXaHXV2fz4SSplKkbql04QIFi1DD
UJvONhYEUV5TklN14poqXpqdNZ+LrP7uzANs5tXr5vS5+pLXNwJDgq5RZ51v19Ba
J2H+bT782DVKdfmgg6KTtPHxmDRqg8aNMmJWp+NJLXwS36wA/R4BNJZ+/X/S6ifL
1IVeTnkrnCOjXyxSURSi/TwGAt4TAT609+R3L8uTrIBLZ1mv+plaC2YiRSohIHQQ
wpOOryp7fFSrITe2zAizKLV+qHQbgrMOnyJ2j1lc8Cw=
`protect END_PROTECTED
