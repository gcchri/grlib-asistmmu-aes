`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eqnnjz2kSwLx3rh3yU9+J6kxh0C+xzQuDN/2teS1jbZGcuRIeJ5BxA2tDsq/o4jP
freK4O7P8hcy76t3XgHKT+/gkMv6tFa4h4qkIeYDkT6nMb0TRkAytusBLvYl3KIQ
TgSA5fU6yjzqRh+5nSu6w60pkraj0TuOs7ohB6PN2Ok7aHiN62wjm7GaXboWggmt
Ncw71gcKftt7+UDPNt4ZM+mQiRVVa5todnj0//PgppEU2loSTg6/tTzs1AG83D/L
Cp+tGViOOQVY2kqzs95pscX1nvOTv/O2i2XwhjJnxaRId3SgbVGOx+UwQh9q3Jxe
iIjGbSLejdLy4hMy1rSo9uw7vDpxvskBTQFpw0inMmpTuT1gses3gzmWO8cwdf1O
96Z50lUZG8IwWg7JUImQcCgxRSQ0WYVETRgthq5qwQr6Jb1ob7t2SKzTJuk8cVzy
qC0oNCF+RaCedOirkFGpFx0iubDd8vwCLjnAdpX/NQeeKCvVgla6wc5Ai7bsRvWH
UZgFub7v+jl+02VFDMZso6Tyc4AF5eZ3tX6KxVFDIeSvzXCXEUbWJmZ7f7J6M8cq
Ebr1rmtEJmioZIgeXkr4O3qRxBv/JAW5tgzf0XlWKgWXDrSqmnbtyNHt2q/VETOR
V/e+aTf77tooA2TvNkfzoGNcCIPjc1E6cSau4S2NGHxntL7pWUBOQdiBOZo4R46Z
B0B2jq72lgmmzHxyfntSsaoZVl0x7trEFh/HcExKG9edU7ksM/Nf9q1K8YvwQNYX
fS3I3md1v/EsLXJYmIAp+Q==
`protect END_PROTECTED
