`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZ8QZ0UkoaRLnw017whiYztiy8cUrlrpDEcf5thESp2nX3SWDS+pFZVroT0D3m/j
WWRKjKbd9ECBg/d3yGtogAp+TyY/8cNkUVWJ0t5cQwZYbzdYqXytidJnAmTv5kB5
CleWLWLFpJAKGt/tabf1qIo4HZZpJ48Gk5Cozyf8zw9Ipunv39Q86dG8MP6NDVNc
1zOit/24Ejxy8DpSFVjkiEmRtI+dxaggygMgY47vA4HNHptvVD1d4G3grH3Ev72I
odHBS491aBUbovbcTv5KDPRkn3isjfSfOMr5vSxtfU1Un+lgmePTK1Un+yDtX15t
UC2ISdy5KB+CGYJjUvtwMzRyELOb/0QpjGAH0V9Nk4KsB1rLgjTVBUuCNgi+nlLg
o6FcHp/1r5MkDqEvRA9b+5OgXSCfAKEAnhPSlBZYWce+b4sBL61n+bua4488mXst
KlyvNp+OoP63/tFgbevY8qNx47tV0pCaQkkADQpfAwqi8GL4K8fEdJd49XCKX4dd
NNzOvS95aMnIfVA0GdxRKCEtMW+36EcGAbuuGkY5j6haRT52bEwnEk8b5JPE5N3O
HUnup1IKjT1Xi/6u4KfGD0Yy25yspDk/78tVpmdQXgkssTeqCYqOIsszDwA8tqri
UxweSRp6Su8Yxw/25EsvWk79cec5Ej2JTFpo/yW4F2h6Dakc5rXwk6AEysUP/3X6
8HguJl50Kaz3KnXZq+eFZy/MzBo5bnL3gmnm00kg3eub21Zy0Z06lXTrnayCAZTl
t23lDdBq5W1FWNc6s66NWH0KyTZGBuxE28nZsysCA7ZcazOK86AN4QmLiQLjzL8k
ZxiH8xdq7dd5HeH4Vj3jpYhO46dwPspM61WAJ21qnXdy8KPQgRLJh47H9RqB9VD+
EBL4QNAR8KBogHM8H6C3L+4/v1QzTE+mm/HxL60oeXLx+MQgNmzXfwbIbgIb90Jx
9eiulHNCchs4vuwssd5QXBtoSqMJXwu4pmmNUnWwk4bxTFRQIzoOoKYt+5vWX0wH
BdH+rx8CdrdQOr6OMBY0SylIooe3V4138UESDvymI/jf7BxAfpbFoQIQPjzxVXwK
vFhMBm1zBhr8Zf/BW0O7eWC7S1YfpaPiRqDg9A8fHGBWvzBVXWcrx7AWKF1WKQLL
ZUiuSuBM7U53RA/UEXGpqU2NV4TSm9spnkPdrxe1a1ALSi6WnbNbKSzamwBzGQZq
WnT4onjVzHjNQ70kYw4i3Q9XnFn9VWeVWmhf+9jODHTVR7+yKbXRVubeh2tP37dQ
YpZHq6RuliYCz/GeeZUa+OEeNTblLmzhBlx8qpRk8VO21cclbVi8WOwNTii/ctyA
xiUKvFQbktQMOuSi9vQdgbSlGUcr0T8X9DhBze1AALj7bjMh2gR0+VygFE8BFoYn
kNDNrpTqPT20Va8uIU9h6StCLVKhdmoSFj/aYfpVOWZDXZjC4lO4niX4mxL0OXAe
P5u+9mTDaRtE93K28kYKY6q8/cPKjA8Jm0HxC8YDNUtfrzj0Nio4zvDD02cFom3D
9vtjjPq+N31zwdBRHjlVQZAJuGg3VcPqsGsXtGWTs56mHKhel7blx0o3S9FKXrDu
D5lC7QGWJcrgUFxUl3F7QteKnXe9YjvdhFjXfOr6+XUKLQKM9Mmv4JX8Y8EQjoaZ
clGkP9DHUci0IRxd7FX0yiSq2CZ9bf892Cnh1WFqe0pBatc4wssrUbWT7ezwrGm5
ZdMqpU4ptxEJtoVz0NXBCayKxB+VOveh1a+1cB7vG/ZmkrpI4FR6ePuZJsiQVGNc
0ccvOX0ia8HkkNOwqYPTClFF7sJv2oQyoyK2jlD7MbIvuGqJFqwmbxdZAEGwNNNn
GtiSy4jCOi/bWz4g2B6rfdIhPfWqNMjRGW7Tjh4MMFybuJyG7N1r0YHybvVOPNqs
ENJFKwYdp6NdMEbKz71vuH3OOV0VCjbnirkTtqGNOvzghQ8LtcSAtKqnMLWmn4qZ
qnrXPXuQmMxGzxBO43go03IBdYFGagwhGXmum5pkk1XHfRIngvyj5D1GyO42Inqf
y3hTHheEPJeRc018VEoaL2T/6KFuU3ijItupGwGcsFF7C8EtIuRCcTOl3gp2Seb+
aY85eTB+MgSCNFeMDt41+L7kKkJW2BAQejk2/v8YlAtSRgzdyq+j0jvvmqerBvri
/mlfrCXmgav+uxtneSMAgumMeEYTHfFWJYt7rKnNah/BxaL3aGrbLBPFXq0Yykpb
2giBP7x8PpTuq8xZFrrZTgdLkNstBWULeU8M+gO4pU+FieIIHjyafsvjREu7wgJg
jGKybG8V3VZPnaLEqX6tYUJbIuK49qHkOqj+g4ZPby4=
`protect END_PROTECTED
