`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XX8Hh1C1JT2Dxw8deBv3BrnrfdZ4k2oYAv8FpRTXQIu7lN27Pmqjl32gkZF+iqjJ
OTsylLMcmMBZo1XPJ4EDofPHxfY8r3sc3m52WTHMI/wYjBgNUPZIIqKKQt/W73eo
Koymx+4C3eeZCplXegwWjbJ3OSrr8Nppxi5ZNZufO1D8uYlzJi4ToqCFEmMlpKBH
i+fH8nOUQZuIIzgjvSLpk8/ly5rcX5/cKWcFkIZbZgGxAtu+nCpNfpPvRiFEIbPP
dX5bM84KSRT2s13ZqyiKtC3/J5xdfjlspTKpHA9nPGJQZXRepuJux7RXfEQs+Pl7
JoW3sSRLYGkl3H0JRD9cXOJzaGVkryWT3Au0fHasPDQvoZOraS99M8vZBigZtPwD
0J4+AHZ2xE7p5wZuwaYT+nLO3IPDrYQFQhI0Kgaee2aWK2iWrKSR6/TNsn8PpEYk
`protect END_PROTECTED
