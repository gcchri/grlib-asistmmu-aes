`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwm9IlUC2fgjVR1hpq/IEqE0y6qjtv/R0r6PdhQlHeO1GxfnFaMSZ2zb5DFz5cUV
z+Gcpx2O0+azBOeV7Yw8jdZjQz2vs7tTWC1cUH+MjzkGDZjb9NhWqPBoxZEY5HbV
89DLeS5/wwVTPOPsrsDWRiKSUdlaHUzzxCrhA9h7QHxTnrNvboP3MooyFX7/kTpN
wGPgIdNbddKREGmiWK1foRA9pw2kvmLio2rgVrJBbNNEFQVeSQgULfpQ9yLS5XZM
eX/dYeCtpNtIBeuKcUmKm3enQikOM920pzhvwx9HnlPFDGu9qdR87WlZPADm3G9B
YTMc6WFwp8RkCwEj8T12wzPs5GVbEkT+8HNzlroauDz2wJewMJlphkkxRG8E4pB2
PTJgD+hvBYBtkZoHrSNNSdWRsKMq/l48+cloSb4tBg/ebcfRNPGIClueJIdlOHA/
1aVqAew+y7RDqV/kruvFlc/pOXbvGh9x1WSYtPNCQ1E9lmJ8BvG8VxQyq4fja7PU
mMPLhuiaXoKTZfXCOk8Mc6MuTDjd0tBMu7Fo92wuOJakWUaFQTb+ROGfbGf9DfvW
fHwRjLqCxI5i4Eg7aY3puIyc03xdwSjS3fT/l//fIro/bm3amBBldiSDu8pWX+wT
NqwlXudZJITeoJ6EHUUVGMq94uuGphF6tw3GjDlPyllAhWjYIK8Z50oC9UeqdWgn
9/G1TnrHnePygXXFhsMRCC47/zEQzbJnUc+LZG65sx/DrQvTVZekDI9r29d3mDjR
XCMBIIrXCixEf41eK7dCPr7+BVAuCNBV1fQRSMFlrBrMj+/8G7reEb2jC6s65uOf
idS0ff9+OZaiLLtbS87yXg==
`protect END_PROTECTED
