`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6T1h/+YOpBMsonok6iOxSaZMKF+A418hEgCJZaZYHowFViueYNEpGAe2z6IYJkvM
3ASmEJahE6AcO3f4N/kfj/UaOZcML8+TEi538hDZUXLN4vFGZEiewAuwQrPPPom0
TMoJb6j44ahu70VEsc0c9QIjrEXwP5gF6Rf+FdhpxwfldjQz0uqeh+wKfj79B0Hi
2poFdeUFIZHiz0AW7peOQACT4oaLSp9Z9LL4bQ1r/qVTzMrUc+RoM5oqCOpC51e7
/k0Rh9zts7WcdPFUBpm9nMk7NpGERMxYMs2C5jy03hrS5H07H8IySgLb+Sb8EdID
6OeYfpzbKJVCDu9ncPis5R+iTeckYUbbo84I+28PryTMAU4OIYsQ63gOux3s8SLX
Lbke522yTmfZIvP5Qv0gQq9U97w1eAqYZnw2luWK16HEeYf1cJK8gi1daz+/bTDY
IUGpw7b1vTV2+SFs6pdKfv9Sku6LaX4naL1Hg7mKqAhvjcqGAXxbCP7YSHCi1qsP
m7KhJISqwNGLNbhnDbaaw12lXDU5OdPg6fds8uvQJqY=
`protect END_PROTECTED
