`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBntWk9qjMCkGf8Ws8kNjUCQWHQEfaqBYzaqxeJ+83JGpP18p7U2ai1mJChI3EUA
47BnvO1nbi3egSRUaNIcJy7PIKfeqZWQdSz3pTQKW0619KypYVrZsr27O20kty6d
Lpf7C7hyllZWykwNlg156ugTW5umycXTF+M8pQDdPQC1kFW3MwmUhbXwQhTlJ+PA
OgtgSFsgHE+5k8boscqKhQM+6IdmbimUKZJGzpFElwsmLEZkSVZpPwpN+lXBZGZ2
kBL7lcimkGpiPUoAmOzQHCnCnG75EY4rbZ/2peovnsZXfeu8TTtiXerFeYWUwPyl
DkKY/usZ10KS6QROrtLy4gfR7cujtxQw+6YRJ0C99+0+w25dxzwQnKWuNvMCHWnw
DKCBZ8qXLPSw2EAGf0z6zkfDQTDxQ0CQMhJ2XjlLSzlJv4W8zJLKfyUirodOrMVo
sRfRNIneLZP8682ZneKU8EAONRJeHlDf2NOuGoK7uBWDeNdV3i32u/aedO0nXZh3
GyY2asbAkl6mYG833zzhgnb8I3qQ+LFbeUVpBIdp+vCtuVc1YcqElAoCs1zMhmlX
NRiy6b2uZXpc8LWzSWAERicOT3AikpuKCJqJTSU06b7zRwgVpdY43Lt/hWCqSbUR
`protect END_PROTECTED
