`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YekUcBp7BSpbb0EK7soI5BQwwge5TiDDhRsVOYmwzsxyaKpmhp/p3KUKE3gjUxY9
ra66qCmj6RhPvuZCU2onLfk+AbHG4SFMVwFfF8jGd0ke4KplCGZeJCfMzd6aPhEW
BUZiPvlj9ztmYLA8WZxloJViT7OTGT/yH8skDj1kCJLorqQgQIzAgiP0wJFbM6X1
stxHiS9rGTUhFB22Ckz9aN7jEs9xxx/edrYKtH+knjJMrenh6OsgUwgvdaIYpiYd
HnjKRvtPkyL5v1kwRNQzpZzxhS7DXJBROWo8TXtGSKuyZ0v9tlhy+QO4Bd32sSP0
mPwoHz7+DzBtEgPe20r9jGAo7gamj/mJqbD3Z1FReCqzQy5srfCDuOS9HE3El99q
5aM5PE1hcVdFi7SWeJg8uu5I79qbAlzySKcPQ+RMudlplGJtS3gNj0KKrFJBCg+G
OMfihLsIMusz9nS+6WdaM9x4UpToKcgsilMDRr/dVyBW4a1iF++zu8N9q6rgzM90
inrpVLxGP2MDrF+Obvq9kk8tKb25yCjpcViOpDn35gxTUc78K6aSSOIY40uOLI8K
mYDd4RYX4szPoxvsdtWa2iSsis3ChKmIDmbOWLf2dWYLZ8EwqzV63FYzn6HG0zcj
L3NvWDky0z6td231HNUBciATFwnUXcO4pvhSBxOqKPEAGMwvUER+H9Z+zJgKIQpy
/7XIMQd4woQlROOkMBm72rMH6zmbcPvcXtZ5Y5fIU10=
`protect END_PROTECTED
