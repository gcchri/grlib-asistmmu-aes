`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J07FfMRBajfnc93u1IUi6PRVHI3FGKE1JMh+cw2wffHcfJuRbC18sgWSSaaUCQwQ
TlrxZowVlkO4m2ZPG9webcf6ByTre3HSQ3QDikefp0z8Bc4H3pOvEM3HICjZdqp0
FM8aPgOKdtEHCALPT+3pIjnEyz+w/H02jWT6WnsbHIl+InSwgKLSZsNsgoldAooi
VcRBNMT74QFDnZT5YAEUDSzhXMtKtO1iy3W9rC7f9GnnKBmxMMnb0FE+Bjeoo3B0
vN4o6lknNUbvWgoJdxUeZtUWCcx7JZvaWLum8yQWvHcMBsS/MaHKRPhMwg/c95ph
n/IKc7z4dBFKcG9oLoVDSTr9cE1vT1qbUFZjnH/BCTblI/avE+AH+YEupjWt6GsP
JYCPHovwTvBg9yrvE66zqQ==
`protect END_PROTECTED
