`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JYETi8X8BTN7XIwH3d4/Hox7VUZEYiQeW3P7mtlXis0fVOZ7f+WMf4xBKXfKzOn
7VdhmYmjKTYztB4qmydKDtybRyPUxnzDZYy73WYrsDdJKHq/Xed8qLGPzhaT04OI
Yd7ctOgOltfTWMLmHbzrh+rHCnpMCZDNvSxVdi74PpArbpqYqGQIdDPs4RPu4HbB
QE52o2itVYLiXmYLEfUl9/2P1GuXpV/ZH4AkjsQxhamB7jlth9ajxM8mwKjnNHEF
Z8AclKs54FhhNE8KY3iw3xOiKAFHSRxsIu6P+scwqHfumoj1Ie1KGftplsBSN2yO
Zs9EkT3VU+nAbvWVLM7rA0vZwte8bhr6KPJX3worbLHayl/VbTUcC8V4bJL01W1n
j5cvtzFFgB7K7SSvtzfN2CeBpf4T5AG3eboPscSCIfmsXPCJ8FL1jZW/rt/QmeYw
ckOauBxP9Vr/Ux1qCpIEXVES9z9/AO6yvAPBCLBzoLeMym0E5WhQiAOHQsEEIQwp
IC5/ryR6Xw8QOtUUcFMwmRXlH2THHvqyJEJWGrSqI9LO4WQn24Ywuld22KsyoQzm
xKDchsAJXYFNNbei96NN9i5IdTdUeZzbbF9U6v6H1V555OhTPWWrcr1KsWAuBuUD
iLaewcLXiJNwOcB1GIYzZe5jntonfxQQnc6tqoFKTbaFFnTOCsoASWosnT/sEkWO
+i7z/tS6IEslANl3K9zcDRfjWW/xyILkG7LfDAjBn7K2AC5lUr9wB5CAp+S5O1GZ
qx45RVr0FinWgkEn3EsOa1KjBNKW1+rNArMD5zn89nlXT7jc3GAn7EupzCF8GD2w
URfKqbMe6fV6rLHoKM5jjD3NKv6eZzXjW+8g6ElDrXqcUROXa2YBfDfEtDm8saxO
yH0+We9g8HN+svnSQR4L15ew2Adq4umaKEOT2seyiHFf4cHcV2OHoP58CdFSKzeR
+OeNk/INwiRHi2BNuzsrfPtAChGLcWNa+uK0x9YdvU3JvS6tlkd+oqZkGsnUMYCq
TXxptE0UFqQ67z2+nGTQHm7QSCmXJrMeLpuc3spvEoccSmiKWljAAY7QN/K/eIEE
sDOdWWQXrDg5Q5nteh/4ZcqUPlECYJAsjVIUHGdLFGeQC8MZk5PhGkFOfzD45H2r
RMtq65xvHhSgIBqPwNU19XhvovqjLplMuzcB77ttpUfc1nq4a6YAabIAjNob9C+2
gIrqftPq1OxhnywVf9tEYMFecJ9zbL20xYVe8VPNjLbumyRh8PUxvTk1SzBiI3J3
9x74r74FKV1y9MrRBrwsqR/pnn1j4NPp7MAkkkT1nEUlWVdr5XpRUUollQvJ3GYr
FBW+8mLHi2UANiai4OLC33xhxpkyCKKFwvmjKyzu4cg9HrUVnXo7GVRSZOdrWShU
Y1suC14AZkh3+nGJ5cMcf+7lAnBsS9B1nhj0FGI+gwxdZL+zkKC703npDCia2dlp
GTMCGQrwBmBRf2fwB5GxlGBsjn8zbJJqIFsmIMG/H0ohJFOZr3OGoNFN8C31qwpi
oUt9f5ZgRyzb4+zxccWIruL1oGp/DZBHvQuiI8D5LcSL4aWRsATwhzDmvVsKYSU/
J7eXKmbYFfn+DTQ33FR73zeD+uZxvPuf6yqxzgHU7/CBNw/vrp08DssZ2CdEzhEu
wjAGNPwUzmT7VU/wkwW+Nd6cQUUZLdljlj4+JyNxB7Qoqmtw3Y4w/xSZqBnmTH6s
fynDif8iYMiWih6japOPN7Av5sk4uGmNk48sZCukBjLa+hCfNFd+gxPGVBh9Ix7b
CDir6S2V//OdEr5dkm/p5RFhCOBBYi5BRwkokCdNpsquCucJlW1F1eleZDbv/FN4
nO5Itv7HkfqVYmdngV5vl2QSYsqOsGdC4le64ZnibtdFnlfc7lm6FMKsNgKZZRGk
8xf1SXaDJ/a4h8cpvr1qSKzI7zWs+fk9jRvqPSYZ6NJD+Y7L8Hlc8w7SEpebTzNO
r9XwNs8srNZe2Cg/tuEkuDSGFyWZnQlrZ8S5zgdQcw6y+mfrkg8xyTM7Yd4b+RSe
LQuN+VE5G1UOVVkka/OVpDVaVOr+L00twOVn+2jhMPBeMagrwURE9cYbK10dR4cQ
J0fPwi+k+pK5QlIWfl3okcMltWrLrSSnn/BaLvrCtora0t4HEbZw5IJsZSA+MI3I
wHyzNgFL0NpZZDz4dHGYbXLhskgcA+ckLE0qSCzodeUlelJml20WlYwpVlQ1N4ju
lyj8NsyCCUwsc6HLqw5grFqhM3EufAk+x3qz5oWUpb5I/JlWef3jmLaFSg4NoBYS
SA+TrJNRGlvvS3LX0Lt9dP8k3KeS+My13c7/My+Kbg6M/DOycwE/UpmmTsbO4m3p
CH7RVpwGMwHMINUefEhF50D2tYxRbkoVRKFtJrcmdG/LvclG+TVNcwAvEMCg/VZ4
8Fzi4hoF+ojQWRCMgE/7JCFK/8iYLFsR8pISIGEu5nncwUObRcFD5ljuAxX/gGmS
InHSwlO5vOXmq9W7Yl/NzKmHUKxZLQEwVUxPpkcCfSf5q1GKtrg2T+/72nUZ86dC
VZZU9UcuhAaz51/vppT88DMKbXW3jKFLZOGJtb5Po7pHwME4CTTg+FMut8WalkvK
NUeMz61onX0vHw2Z6oplo2YBi09oo2lOLUUDPxuiJyKfSY2GAsXLGHif6mB9Q6zb
FY3PoNVjixebcLFcfAyoKvRP4PIIc3gNCszGf11eUIvGCqeEiz3vKLWp1k5kX+vr
EXWsvb6R3di4TppHdJUmfiaVCbAUfm9aX/ToC1g7TpoAx+gOcmdFwYtnYQO0eG/E
76RN8D2UOzkR1rodHAKk619UGgMiv2qDH91SQv1aCaB+Ji1cHIpMExiLfg35VrUN
HF8xi9Ixy49xOB/JXaHnvg+L6Wq/X5VVezxfGUqCMQvvjnCoJ5RROTaAZhrvT+9r
fcKQOVUyljf+Rc1uTwb0QoXpJG+oFfsbN466oF74d8NyC5bcr3SvamCwTylZVdvQ
L0ivuNMQyDT/73TauoGkh/7I1GyyR/dqXJk35XbSuWghjoQyzdPueqjQKnZ6Shej
+uwUlbKOJDICNMqfWbZKofEYHyEC43FI687NE+nrDLuss6JxtGWB4VKE4Ssz/U8v
EXigCD77L8kVHDDUk+Dsp+rEXFLkcHGs2io3yKE9dJOK+FHr8d2zdHkYKHSv2AXG
uziQ9FSOPlg2Q8ikJMPJqJDZMbOQQpKQiMVetqNPu6bidHW7h7zb7uYImv8kG+UQ
hclPUYggdIpKRMtB69pRy6uuO1Rb7WjTWRKzJonb5brkz44j+HjwuQkwn+Q8+vcY
bn5ANNwhFgteNGqn5L2cRdhRDZEj0YVvyQYWmtYovFTL4S65w/VNJCCP3C6H9Rxg
aOj3WuX1DakOjIsLAar9X7ejDv678T9/02ECBXYODrZ2mCPE0hFc1hpCHZdN3Bh4
UbFOAaO5zxEzQZh+bfkHVe3T89sW6np1vmr44mDxT+MH5xXpCUV6Nw3g8WGdpYHp
DdMCaJnnBfBNz/8Usp0f4DT5bHR0KUCTn4Gg7z+sWSFpB3UmRcI6667JWhO+MCxv
IbHz3YFPBYGxWJfts44JlvyyM7SjB24OEBKLQh5irGZRci7i2qu7kdnr9OBGDWne
cfeHlHwVFvFcDiZEOr2ciCn5G0E7jR8ZKF6Om++bk2NENS3JGWk2C7mHVgnUY0tL
zuH08VYkz+DFHdK5hTCtu+YJZz+r5g7F2dPM9E8Pzk64LgMDMs9Shw2Q2cYMhd+E
xyZAPTkWIgZQrVHjq4a7hr2eJm4cbjYoI21JD2jC9B9gfeQnRlBqV+WGsb2RkPRy
hjqy4fJG2bLq05+8dn3MYGRHFbqjUQ9cUmuevBYuibMjMrqI1rHY4X4qFHMi5Y0X
UcEM8FVLy3xE+G2zz/C+Pk3IPYYCFVcR+V01y7tOuN/jYr5P3fczAZ+cIl9tPP04
/LWJ2eGrs22HfuHLgu/KgCkJbBthmQz3fpKfbR9ooHGqVOEHEggr69W5x9dIH4QF
1hcMg03dIQoIukWOWu2OcmG+6FWVA6gUJj5r+VkCm21EiiucGJy8DCLpjEVbIVnS
j7Oc+W1yTg0FbAMqki7lAg7oVrb1gebUXGTmT1UcbWOWHKCdiSmqROtmVx1dvIiz
y9P403/gTdZbVIGvXEiwnf1C7x6L4nsi4tErmLLn8YYc/z3iFyaaPdRsDELcWnxI
ir4lN5zpUDP3pwwBY4jpaPtwHRTeKdJ9fFEjfw4q++HaPXE/8rYp/ikVEMeb8dLv
M24rJb6S8TvtelBVB7nJoQdbtN+btBT3kHKF15BFO0pCzlnqqlqEwfvbAZEz2d0M
HFfQSfKvxeevQxvGVV/54U0/4lSMk/RtGwHLqPV+7Adqj5rAh3TDu4E490PYf7Og
hzPs//FKH1XmkPaEHEYJSIHalivHRFRumdkZi6Lwvf31D1dLPYEf4ix/AgMZWDDW
G5dse14WaWxr440EpHjx5f1oppANKGZibNJNix23AeOFhDJmE3xXQBxJcznUPxfv
gJgEluOD4WW6MB9qEc+ar+KDtC9txDHMCfMBhL3BoQXv23djb0a8toUjwc21gTwZ
3AXOQ8UIMHQ77WZM//LA7Hy7XfHxiTNfkQLTae+6mHINVFm13jWDuwPlH3F9LfSs
DG8qCgdghC1EsFDF4WnEJfa65vOzg/ze+DBQLNC4QayOpfSAxQWoArKRAdfUrYSZ
+MbE8ronb79/1PUUei7nIDldH/PphjY2FplUbk+DMelA92wXb5O3OXaajzVonllO
ZX1ECgWNtpvOHEn3rIv6eFshP1GSP1t4WC1PCprWFAfk/fWOQPMXhxZVBfWK1qeo
er8aEzLMP7cV7s5qu/UCloDjRCvPovKYOe34l84sE5Zd5yLo+g2nbqTY9f60uh2+
YtjzCKwu8dFewWLe2zMdUuv1jgBt6h7hF94lkVVcj2atySZviHkjl+C73eWxPiDb
pZ48isP0mW5zbaNbmJtt4iiP5QaFlSy+I4qWKPsQgxHPWvRxEnVDlz9yU4rIyss/
0KN0h8talzjdUyLLjDL+vyVNdq/5EXgTsgcyq6dc/k+tZLTViuK7c18TZY+7CgrQ
l5/uUKsPJOmo+k9oQ2ppGGrGS7QFtleYu4FKsKTKXP2ReHl4Eegb6ufqOycckhQb
n92jyfS3HA1FS62ykS1gTN2/irLe8SK8fHVqAKN738u0181lA5bnCX1PHwSKWLwD
ukh9QpXJQdy4A3tZismQGh9S78fwSwvmfTSBHhEZiv3cNQ4f+E/XUzM2ckYYrZtU
zkRWhTkJpcutChWOj8DG3UoGCKRekRIc3q0y6bsddfHyR4lq5uX3LIyqp8zOWaDP
I/LDycLK9fz7iarnR+lKUPDrVpI078yK9sEy+Z8dZ/H7mhbqQrHqHUAgqs49X4qh
OXiMFW889tUkxwW+7kYekFdtA81sfTOYvuzCWXAqP9/2EobPotirb8sJ84UC2i0M
nYxnaGRckBhh4spSUIBe6kzLz/Y90Jhv8fskKTa6leD56LJhcf6rexISrKO1xBZt
iQmFvl1LuuYNVe5qV5HhjPI7J71nIXuFPNHjd2Z4Kg3uBcQHPbS1QNkO1Pg1IQTL
Lob3QDBsG7HpRm0tdbxcHzzsoXxXeT/rVwmzkuXNDbCP6cGhhowK2hcHw8RIZtpr
9uEpYlM6gfVhWvNuZeb+xyHXaAVF8yAlO95NnarzimPPGvb33HzzF9qJegCyUVfi
sxXLpQtqGkWLnyOsEwsSZAIXbKu1Yyoka6jwOOyXuOCL/Ae3xQ7QJPy7s3DO15iv
2LswWL4GkECk2aliK556WPU9J4N95NCAj0fPS0QsK9dh7OzNf8qMSxvDk1PWxaNo
3vff22E5iCPzm6G2BCnt9dj11B/IM5szgWH49ck4zrYLA8AeEOnCSHECYnvcm9Yd
sWv4Y4RqXQuR34HkFJoWuNFhvrykHkJrZV2VbzL04Lip87vT0hldICovW9LUB39D
9Lp7kRxbj7h5QPEaxlFEm3FsrnsqtF3iVUI652CiZL6cAeO9aGUYGd3ItOvltz/P
BJeP8mpqq6HAynFzLSKZeJUBcKtk1UXpv6GqKi6iJL8ABem/njVzc+xzuPuT3Cb0
gfZigUrvzfbXdXVkKjhLwa+AjgrmRWEHS8e40fxuzm7UdDe6d4YsI1K5GoMCvlIh
QZ+p9lHRDWfRNJWQp5+2A2JgLcn3ctos+hYLllpwZNBRDz+hSmIhObGzARtQDL+D
/ZsVEsno/2nICSbVcqj5X1okPrwusus3ghQjd8reGhjInElAAFJlosaQ+eJKJFUY
jHQiN0MA6OWSBLbtloOql5c94ZcHwXBfilhImyzyglYd/YRUVqF+XdeGDlkBen2G
HqBfL8wSec9TjwDDkQJ+gbJ8ASx070cW6dBaNquK1PQ/xH+SxjX/7jN5wRjmvQvy
AAVkfeDDgfm1T2zAibXre4QrHtfz39rACo0AzmkuHWlmhTiiQ7k/GKS+arlWVOlX
obPzRnLFEc8DQKIYRDLmgVIo+WSpK4BRzBG1iITpOnycWofXqUjVyxwq+TckARCK
flDgiajDwCSWHHYL/U5d4GyQequh7jGXDGkp90mrDYNy2NPLebe9Kq0sqiBUokua
Mhswf1LzmTlfyKWVxrWIEjuhWSfDIJLIflXduEfbQuXnAyzM5Kc6j/G9O2VI6Pqw
8NFG3v9odp7tHBwZ+qkPwT8vG3kbbj9MzK4O6XQJnYlY2lNcuFG5FTJgk/zCoFMH
FLr0xjmx1qwe5SRJ+4awaKoHsWG9YjcSrs2yIqWIb/1SmKGNAM7i0LRYu5bWMocv
b3JCaIq/LN3fIGQNW/s4iJv9XkQ1GnMkMCcB7yc29j9BC1+0qG7ZGHEPCrTBd3ku
vMrXuHxGF3Hz+IUSCutTDnZax+6qGDMdFwyPU44kmKm8vTtrmcIxtWwv+YXaaon3
Mug7pEhXE5aMHA3qg+yjliTI3eyWzdF8i8kKrZM+aA2WnWfZw22pjtBGDLJFr0Mm
SHTO5t8eaFSK++d1NdB4hNBI/RmNUFsiAIQj8nkECwFQ/1oTqszcLM0Wg7JR51tW
pAUXBAnKsjdgkoOkyixt5Uf/RdAWr+LBzYeCgh+KtCADY8vOMLBZXMVGYNuRHCp8
n0Uzuz+jm2AtyBmzRQIOE7EK98DfkolQvyaLSdnrk/s8zDBqmSYtbt+YoCGtaMZk
/HovLFD548EqRNOGytjzKDuHiXMRLexyJGP4ymULm4HRHgxCsOuPnOu8kpP8GFko
So+ZqAXrhe/QI3wkxigXwrjkUkPZVogs2TqvTEMkXCCncWuX5wL3X4ZiRx+RRSmV
GZkMTubOJQTRCG8HvCNSACzXg0fWub8QqKIDqNypk/j0XX6cZskgvWfW0QGwpWed
pC7pVZVGysg1KNGQtyY28aNMtaXP/prj4tI+9Iy6+uNnZ+OOp3wtDkjUwCdn/hJE
NzBDtkZrACmCjbyBa3xAocrqij3GaSsFOU/2QNlPQbHX4gXIS4dm5Kon4V7pV1fq
ZR3EtlKbPKsRBDZvpllV7fF1R5Y00oH8wU2Q5/UPHEj1gUTDhKso/+XYXWZbHefJ
JqzKGZ4IqqUL7P8N915GKxMeTPGGIg+7SqulAxwnMJrkIPp9AIjH2dN8PTJ5pQUd
jspzGMWnWA1Cdn2PgHevf0xozQ5sdnOeONPgdObWEtc=
`protect END_PROTECTED
