`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TaJOuvFGwOllEpHMDRXiNZYFseo9/ubJL2k7NiFRuQk8rEdnR/D4cVfBVlspFh7N
3io7MdMlhZu0PX0K3/sIjQN6/gwnr7oNO7F4d1CpzXbVlDkYzUj8K8BW1FNB5NMR
YBVna5YlAA/EO4R1lnl3RdWAnIizPNnmXiOBv3es01atwoSON71xO5+fdSjEW6Rf
jP5hIRwx9y22oIZbyWHZqtd6+ucWK5jBNudCMM2hglKD7A9+6KeDYoIQjmNni9hm
6Us+Naybv6seV1Nyqn8xdNeN2SGovnc07hC/lBuqihTg1xcoN/7lVVA/T2EwBUQx
D2pTsOBFrmnwCtoYaaF4gBBUPquinxqovzCZ0CIjcEavUoWI4AkJ4yOLnbA3Toc+
NYh5+WHK49zPJKCgdcGVDs133bqEUzb5469AYsakDrTxoWEMuwS866W/U4ZzBpQ9
1qPJJQVKcA8/6S4SvuHjewzWzvOed1bBOS5nM5xLt0Bk6Ps9whrDObGOs1Qo4EAf
fxcwJ+KLYP4bhI5ntx/UwbV+vY7dUG2nV117jxmikKyOmW2CQZnmXsU5E4qA2bgV
YN7EFeZPH7rhkSEYDhmuIToOIGMu1kCSYLAoybn3ue4YNNNXKPVWzA/t7T0Mmw/B
3FL5d6IVFgB5pC76vucIUSnEsd8uTcAzuFkkd/ZQ2qmVO1pqo1NDLoS1WfKA5kiC
ZJnH/lEK02nhthrHyzpOMZ7pB6rt4Czgryd/OWySGko74E6Hn2YMDoMzh8AUugwH
8DfoYzxoLG3IrCRYhntE0n8oFTTI9b4TXznNZPGr7c3AUrhTAoodWGDWFsWqOE+9
l9bz8W4pDNsmnu7OnHAdciwrIvim5X+3Ped3ENR6/njMzd27yP1DLnv3mwW+HzTx
xpTsDThlOWPuKFNDZeclXVKZ/lbVCL941U00VBoXIh2N9yLr6VzisxkmZbcfj4rk
9Tk4YkAU3Aez+/lHjti2uWEA8QGvVZAp/nu4qIV/308rjWlyXB+2YdV6FKBOgGkQ
Hnq+0ekXfghp/x4tEkfQmtIvHdhNji90WK4PAC1qBAMQmh02jbR3YueqX8VPpidL
FTSp+stOHSQO1T+TyD2TUn6GfWFqxmUndhmjiOgF9wwzAR90VesDd7ne2xPRUsEI
jtBSbwv29ldEo7v6MB9Xt0FVVCZQZWmCr8xAAhJD8vWvTO8gxu9Es6CDmj0eOprT
ye9kKMvUwrpwSlVfI0zTQ9ZW7H2oS8L97eGlO3F3y0cC5579KVDbPPEUA7NM0G1E
iTm+KxnEtZketOS1XendJZ/PKKpbTqVZDqOFf/hs4rRpygM7dYJrjsyBBmTWsyiN
fxZ1dUMJDLZup8f6J1jYvKOkmdga79dLObk9EA7qrntVvMJ28/P2dPgdEwtKYHfm
N2d7SamdKiJmMgyIufa6CkGkV4MJ3HFtlGI12gMgTlrHlxl7gwIzQlUvIWV+QfeD
1roZfa3mhHa+iwg31Tyr7FuZZCG/HJQGQlYt6hrDMyc7UfyKHojRUFCMCRmqvkX0
F09TgCqeF3rcDD546lhZVx9CwxveP0BDr9ParhyiIJ0GMY9rmPHK9GIWBugLe13X
SES+L4Rc5AmhKCaTsmCtQt3SGxzcQEKTemu0K4n7E2R4tqU6q0LW2DXbo3nLYyPQ
ChK8pmJvOhaqG9UxIfNWkXT/OTWnTlfDGnxa7WeqwAQsuX0zw0ycHeYWfR+KHzBO
sXG3VmWXl02hAxQUvQ3qavcAtUj+ZaIBmprZNFywL5MqCtmVgxc1RYi4vZFK58UG
SlYC5U1OlgPw7o78rwKBG0da4PPSUvMo6oKJgUCBcPh5q7oyyjRjGjGE13n7g6VK
gV7a1VYSpm3jJeXtsiOssDlPjaZ2d28ohz0q8MxEYUjmW9WFkeYWvv2Cdjks2DVW
1gGdh3vhXhigTfDXSmBFxxU6pXO9KLJ0lhFbI83Tz6EY+WhEsk4dyzT1ibgY+kuv
H/O3gLOTPLOqPhCqnLRRwMY91FCb+UbGcVXOiL4elYet9FKk2iWGHi9zP9KD7a2s
8HxK6lL2rdauhR+Xd789yxEjkjdFTkpfsekbVXPNQSQ5/V9/8WQ7g1/iOGFmvj88
xiZYTtQwVFybT6ZL1aCsq0paGK33xBxgqROEkE5bUy1zRJNZZHt1Lc/lJHASoRrT
tp8GXcRgMCD5XwvxIIQAxAYrZrGVOHA5px/QCmsRVcSuGZ0Zb1qVuodAs9ofYaQ1
P/opazWbgsUGzxi4c+mYI5vFJqK4noMEA2sR+9Um9Djzz4/n6tYDzKt3KQPCNdLd
isPJFLrVmpbyEB3obmoWXQKJxzpWxiy2Th0xiQpY6tQnnqgNDN5m5Zvy1Ov/4osE
`protect END_PROTECTED
