`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aV8qVMa8nkjFyq3roZac6QxqfsJJIE3tjzPlmoT+zoBSctbomIKih/kLpPI9gTAu
tfDq/lCfaSpzu/f3La6e2/nty4dH16DR8kZbKTtT7TJmFLdlaH5JswegTLvWx8lC
bAeTS07ku+noW7FeZuvJeNYkXd9Rgvl0jtK2UHPASyviKPokd48wCvAn5Lm/mtwa
iCi+k1m57lJ/6K00YnY6v6gaGWxVi37Oo71xyoM0Kf/yrKyZzJXk7JdeMUUAnwkk
1hPaqIRkcjfeetxlFitAY1Sf+sKxPdnT/ck8F2gkbauyo0EMmnSPcYDYIFVDTjI/
3oIxlEbrxgFkHNxIKLHvdE4kwPD+FiDNxoLZTvHmI73KA9vyyVP7TYRhMXIMzIfP
rmI9oBgnfAQco4yOC8qpCmvs48KPd/72SYZnbGRWjDSxFQPAI9v3zL1neibSSdt5
`protect END_PROTECTED
