`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sOB/Uz19fAUvwUDlYJk+kv1T0vWO6Asfo8GcEK2t12dZpFO18Tw8wYy8FR0I+SM
ybsd1nIi2Jsfj4qc2I2IVEe4e4au9qKlD0iMFqDFRfH893ATtGzlbuoacRUA8Acb
6uwhDzGKzXjL9MercB4akXe2dCckQH6YF0oxET/r7ckNclbVGZ2cbW1CFTLonnJd
bLbA1nXvgw1uA/AFvGaJaAIFooJ2UnzrXAB5UW4fhvnXZUDbvqc99wPBpZfinum6
XmntbZV0faRrFswYjQHhJE2X4unhoqcpMuHmdY+xTQhv12/PtplYQqr0onaPLtRT
4BiekLS09kXN3afQCPKrV1tsgQ61Tjj7ggYXWl94EjieHXZwkxNFgn+Nu0YPCL+a
ItC2V3G6gTLinsYHJ15qsRIXDzBijAnTHpf8XlxDhgNRXYtlFgGadmKxzuOUDl/j
6wZVBgLF8ffocyGmHn2JiynkaW2ITBfxfQiUVST3A7EITOIeroytAd6UxANOy7zK
ecdfhsqsvsDHLhfyeABljWG6ydmi+PWw6z7ccnHf9yDyV6MaptpVVzLzcVgOR50i
xm8+mrMbdpqYYnRWsdndNTRM1RKODAPu+1LHtVMMulWd1RX81IEk1LBm/i4YM07U
y3aG8r7mgvJB9yLiVtZmKYYMLHORuZb5ZF5rN1YfWDuMrM7QHNH/wgHD50mI4mYN
xRRCppEs1Y9Nc25kxEMtY6SGk58MABiH5EBLLd+IABPzeP+tlCYUSVuinii6qZ2q
ozcaEv76U9mcZhRCd97ni4qlh5jDokelpbwCUTBhJG2B59Tn+lchBZjRGySg7a/P
+SFXXIEJkQQ3apO5O8jXP4WMkwBqbTUiTM25m/oxnyjP3iVdeAjAO6F/JEIzVr/w
MRs2wdIRvHwG9+STX0FYtXU3DxS8liXnCqcOGCKQ4ZSrHRsUgBLlsFcZy34HDhws
Yk5bgvKyJkGZLGwE5i6HPTlOHoAQP5Ko3a3GNy3qzfTK8NgGQGXxCoFs8UzW9L7/
nF/WWVbnjcCCbLXmWDJfWzWsctdMcWegA1sRZNDVRwSNe+YAvx61j5yGhe6DndBh
FFClH02xMjgekSPZfxD/wbpv0fBvBJwKSIOeJCSVzGEDFR1Lt4scPFYxBf0vs0AD
A/9vTSTOzVvnYq2Dtn5n1ThwTmE94eE9Xyqw3cqD2cSwvuNA+O695X7BtZmFP+D5
itdC/qAfA77GkD14ZLX8lO76yZeZRRmNzoGHzd0cHsg/cZv/NOSaZmxWPd0eLBx/
vcZWBuWaNKEp2qPnWYzPOFe5F9IdXvpvnObDw3aMDdKOIg5ucMKWeRHHKrcFqwIq
7J7aRCf77crEZvOSlIXZFB+jalLxYu7aEGxq2YuIzysLEVMFtQ4i7j/NmPfjRINi
kLRlUKfNaBwwgT4nsjgNatDipwP4Wgfn0JdEl0Zkk3zpAnfUws60d3IscnceN3BF
hLvci/t6jAzvk/PZAW+PXyp4GNtXlJN4qv3F3kVxJs+ySDsQYAod24Wfj5mSudKU
5yyPqOzsNmIJptSNG39/kbn9/qp44Wcw6XU60my9aVkr6fxTSB6yqrSi7WplboAa
AWOGtCepWJjO8pcrSc2n7EU4ZmbWlpTaiVbAHgFIWWNzUTJIwPi7qMFAXUmoFLTv
qxpZhBCzjOpMfDcsjeR8XDF1tVguOigZ/hSlOYtleOFCr4eO0JfA+UacUc3B4PPE
wQaJISm7huhgsg6LKU8saVvuzH3SH8FVFJ0yHG8pMGJIWa0UEpOg8c7JwnxpC85U
mhtq34QaL3JcbBoMAcwH0fZIiKyeOJCNbIiEFBUDJDl+oEwzBUX3i/snhh1L40Hu
+KL9UM4qotLzE+itS/mvygoBwtzQObEMJq/vvYVOLW5wK/svgV7jP8yOyRMXCf37
wkJQLFKSp1OrLjIa5XFvEsvrVEFqWjISZo/eHnYAFux1QDws1opBlyboJ0Sa4xxT
3NXJ9WtFEfXCwBrU6FkvrEA5nBSzol3l+SfVZ1L2BVCeRi9e8o6zAtkXxG66w39y
CP5alH2jHbLFrsNSS4w7lt/gM2OLSE2zllbw4QLVaksVyH7qQPGARnzmU2nc2Y2K
OeQknkjHhanTx9aiK3QCgipPpBcMg3eurNL7OYiO/vWMKB94I9QWaBmYvXCws3aU
`protect END_PROTECTED
