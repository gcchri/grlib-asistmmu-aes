`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E2fz4ib08z4Fxj2qsnkLrNhV9i2xBMmGKU/dK9sKF4NXmmerbnq7V3e7BbpwUMDb
VnvFge13ZdDQv4oY+dokz9hpcZoAXrZnlcSQwgQ9i4qnnnrPimRnIsEBrPtADxGL
oqQkEHRbu6xLD1dUOYMXrNsecZVl4+GW++WSBVhRk9Du6juCFzMpgat5wGgwkwyr
tdLM83WPpEbyDOuJUSDzch5w3z6txclD47zs/DxALJ164MvZgLAxoY+VzX4is+4l
tb0FD+GLbVorogqExQNomMdIipoehBqAP0+fscAoc2SBO7XOO9xYwthPk5+nZV0q
Dn80CS3CQ5uQnl88nkYM15na5/kJZxbg3FBS0I1r9kvw20yrnpvZetUXXUdmhg6c
W0+rGBK0P78sVn30Kr1HeMZ0ZVvRaORMpoMQvS1yqaoT4tgbUvKVMLKS+2ajbrh1
SSkQaqNAgT/P/uYZfwb79P4WOO9pSk+6c0L6QtJfY33x4y4MZ/k/AmgTiOyDdhZo
iIx/UTlL0Iegk5nZ7Eu5G2lC6Yty1mEgOi4aE2akAP/uC//22TenMrY3esfTbBrp
PMNVmuEFRT2HxwbCGzM+3w==
`protect END_PROTECTED
