`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwIveAeojdbdyxJAe76C4ioUR6k4NjmfIOOcV2F9wJJgA3GSargKZMkx/C7O0nVS
AUpQV0s2IIFSRflRAyBnHdjPaJ40gMOCw1odVamM2vLBnBWxqjNaUpIcpP7q4d9H
wT7/ryaATWFRe7Miflh0KE3jZYUi02oSj4h9hPHSbSNaRtI853Gjj2nJ45Sy6XRI
XVTD2Ht6VA5dde+/MpRRXPxWmpxHBIfgqpVkG7DwV9gwTyAH55SXKVbvpCzs1cck
wx5eCmjQvqvPAMAUVB/kNsXR8WaBz7tsYDffjenpK7FpIW6iMckq7fliGEqYJ2UM
z/cDgGYc9Z7S1172TOZ6l6yVi/EljWm0GklV/T6W85Fl0MK1iyt0ArZ3ZWSNBkMR
1dC/ti/8PzqRxy+Ni7sqseSal/jG/oBOMvT/2aw2paJRbS9lfyVvTKK+Nt66/X55
CMuVfPEcCmcKqvk+ckhD2Ra2w4yQvRs0hHn4aV9qam5RjrT2SOGTo4PU+FtQwanG
v86y7e5sOw4ILeAoPv0UZLauVGgDef3ZESk7Y2oa+FGJBO4mUGuCc3NMUi/BNQ36
dBcW6g0CcGdoJ6aOmH3CfbuDRHfUcTHOR2wc2V5rdDbVeL6bXHccaxRSb6NQk8cE
Jq45tBRl0F3IU4n4tHLzClF8NTDFVmASt/qH7D6EyKEsu8hRayhD54telDcqqhXx
4H0FJup+ZDGFFe2neuJGVkt4DTPsoTpNw7qR6xlJIX0kvsZRGWZnOlanvS4V3oaT
P7Em0s3l3qJyrs5v/EMH2a63soIBTyJ30smWPvCzHFyZvHS2lCmk+ZOB/CqvBapl
gmsHvSpXU6XdwYVvNK6W20akdXpoAUzhGgPQFWXVppkc8QDZpyCNIk9HJRHbiiow
vGaUQCwnaoa3s8sPXZ5fJ+k1xLJKxduuVqNr/t8poIZ8IyFw84l3PyseI9i4B8h4
0770RUaQUuq3YEcz73IDICA4Wup8aKMAxC767Uniwb1xnCp+6l4PxLU8x9TDy6Cp
9Nye4Qqbs1lQGvhdYEn6faD+wPYdElZFodJjp6bPsusqveER57i6G9SwDuxULNxo
6fIKlHvin3Y5MxhMHlLGbLsLY8oIGb5FYqn6Lb43Hklc59diFLsWePM96KnQeVFq
SA7KcIpMw+u8k8bn0x6HN3wShZuycn13YnhEIujl+zPXQK9t142unwNJkhN7wNbS
zcI9kQxxcWJD/F7cb8kbrcLk+M7K7nnor65EccO+AYMPCwjnq9gBdCFUVy3sDdN0
SLTa7mQ4ZhMaf53wk/PDFO02ICMn4MveJmFUpV6AMYTvXhKWHhO8fgAHO9R6N9O6
AD/F6wRoUvcNiKHCoGZqHMq21YAaJzDMPWqdRUCf61OKeaJ0KW0LTnDWX+1IK5Uw
g7qzvIgBckhguYm9e7Boj1E2ctY39HcjknfKOUoW9ymEqm2tWW1xA/gvWleyuDnB
Zer4dVlx5cqRQM2FA2j6QtdzqhgrrxjU36ujaCD+UsOrQnjtQnVRKpS40d22UeZy
wq6njHYI37I9p/5atnOn9YIqZUSBrVaXBFRLnbVTpJS/cj3All5CTQiU60tF3sSd
MSZGnx4KMbZi3KKE0/sbAXS7YPjzPHScDpDupd5reVKzk9L1oiaaUZh3luIgTjKW
IcqWu7MfpHEwV4OGD28ydXHmiqLycYumyrdnZI/8sjTR9+IaX0A9shi1g01ZmxRT
2ObGuxhQDPFVdkAGz/5HlAukx7OZQhz4BxpOqjdHDbxuErLwrf2XLBybGXcGCAP3
xihSZyRWCZOVlKolDWrtbEQV7NgDtFyl/ytNXvDiPDuH7jQ+sRkQvwy+Pi5LN5z/
M40gvfHpc2ny1DWdiAadZujHGs+nO+NR73xEOZBPK3NQdHBLZ/sJlqHhRAPO4xUC
Cqt4CJmosCBGFrCbppkMAJOJW8q4SD1Wz7eVPZscywaWa7eDEPoPgdeLZ6tKdtM7
elm5/k3qaYlVKg5hjbhwcb5fxs38I2WsNoSPuEUQEfdmO9AqyGiWSeWMoFrgUEr0
QsCZQ9CXqyHrFU6zn8FhZ3Epv3Abqk1xUbv1OzY+OPY4QJU6o0U1u2gR2IIkdHVr
qynXmUoyrTKkZKuW7PYpgMZewLswRJuwTu/jNOPsEYDjte4imqjnhaYYwCjMZLuo
n88jpixoJwJyti9/efCuSB9i6JZzaoiFw78VthIJlLn1OxyVzh2b8m6xw5+gubxk
mD30zGFgz8QTbGyuDT5V51vCf4VeIjNuk5p/Fnn11Fc/1urUAR1N9voMNF0/9Hde
0rXWQhFstwYTV3QXC7WnU66GNS2BUjHEH7+krm/KA3UtzQ9EnK7mqOTQSR2elOpb
5CWh82JJU00yH8aRwrPT8BiuKaTeMB0CAoRfUzL+HqSgd0uAkg3A8YVbub3Ng8wc
SwRxgI6pUkMLpVo7lOPxF786YF+BoflKzP6x3X3knv34uChLH3jacrD2fkrbReA2
KfRpaYJFklMGcUMN7RovxOvHGnIlkHb3GTNUf72B/5XAyOpBZ2oE+5vu8/zAQh7x
zf525ttzmRG5dsSG3CBNiUU8GIsXB/gRv98iJaB90ezXlbFvQC2+dBOV3n+f6CyC
RdWfzPRUN3T7oGBYRlrb8M33ywD8TB9KJDNpmnHTwGXoz2nR44bQy2Cq53/SH484
zqKk2LVEfWzJ2mWHmjCXUInSwU6laUdvjjwrKvnPYBrRKVbKHVbmGkiXwyrYaumi
tKGpioBXgiClrLxSdQigRnd5GGq7M0od1RQu+s5Ku0RRuSdiRJsU5RCTChCstKqP
AyRtb0ezQ93Ru9+SW/PDS7drRJ5Pe9jsLLIXST1TCXkvWxLUK+zi2j+peQy+i1X+
LJOXZQ/v2yYhWf1n/DCPFvYAKZENEk6AemxS9mk9hjOpb3l5hffJOdKTK9nBHFNe
h4qknzlNRxLzFYhRD6iabZYmLUzPCzAABVX5e0vOh18SeS0X6ELzQWA2KSFTy1Cp
04/cNW4CHyCokYu3+kIcEgdvYNs3DCg+h1VNWA8jqBKY40jAcUM2yAzr2NEL/NM3
5tHfcxBLTFAAzNfIfTlmKHp2hdqbd3pxqEqGUhrPxyHZlzOfyj4gO5mslmIzAnZR
Ka2IGkRnNRb+XEkpcnQRanILQV0xJPsVsHdGjblajbTVoWJeTYvByZ9/b/fiVy5K
n1kbHENwFUs1fviP8Cm9iqovvA+URpggPu8nSV39RdFJhRTA/f2xAAHo0RJsYRJ2
ODNuxhCOeMJDBTV6OA/GsDS/A6Zs8Oz6KeOqbPOJaroOjFBA7cybv8P39OhSM7Cx
aLr7e6+XGhpOy8mvxlwXcPkbBr1RaYeqyCtq4uukAAfC84xjfTGn4BGdNT6ivsXV
0p/hBair3jDu3uzqtEhF6h6axPy5a+3mWcs7XScioufDuaic3Yf1XsyDtbGYBr7d
nw6dtXhtV6hXv6sHYZuckYt/hze7RICYcFsN7PcojSebz4m7ZuSE3IVDLDP7VBNu
OCPXgzY8FvFsxOJtcbitUSrTv9V0hUMDX1dv0EVRN4QW8QPYDjaBFEQJQDI/LI4Y
6tZwcf0IHiBb8zYt0NmRIkAyhYzBFgUEXI73P24+bGX9UdYwxc1+gzWUcPVS4yWG
`protect END_PROTECTED
