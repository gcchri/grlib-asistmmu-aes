`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M/c0feh3f1DJlLP0K/SptAaWUC01wmNAJMNbHTUT/KQ2nAHIkwtcbdJVkD5gbZTX
bsHpnQ3gSXiKHM9mVXRmOyIdzWi8N0jsnAXDoSXlLE1bCHVMtB9KWR6v9ryZKKyN
TP9wsZA7ZMk6wPDNad19k8JGdx2xqH1CSrj4KP755AHOdiCSFjvyAqbQ4NAHwNWv
39pdMQDdmwctVu4rSdgIupACFhbtqp2gIQffVZLWkF/Dzy3tTW7iEpvkmOfyavSi
ezPKCP9vcZQRbv9oa6XBq5opg1tcxieMArCIy57ANSGRHMcbowx0eBT+d2E3qeQ/
GbMX0jEfBH0mZC16ifIfepB9t/prWQvonZs+Xq7yxcmtNZK2nZ698gap3ttHxXxf
+aS/MdFqKhOeJthfFhdDtKVzrgCuyPMr2CjuVIEx3Z7N8JhsJ/W0Cp3CnOcLsglL
KKuEtwJoDVwhAVUrNx+KpEQzPIFw8USjCVgGR01TVobR7YQpJH/l7bMdwICZdWdI
8dgx8VVxUwpYHcnTMv+kWA0VQTXpL1RwR2k0UOnqOMViR9oKpiC37A3APcLK5smF
T5IrjbSKAudCVufQ7g/VOj4J7A6TuStUKRhN1pkzD4c3dVR1BlkPWFzmDztJKXdu
x2zgsJslo4mIiVyRznV46tL0hp0UtnOKhZiL/a9HXxNTLAw4W/17CcitqZtH5y+l
V9tyVc34l+aggrA4aLE7+7lew2zyTFn6+E0qYxZyHvgBMzOu1XgTRekZ1cQH0KIA
p3isnBx1CHMqeRQYSKv/ILSsJDXOvC4tvtnsAJDC+rdFosePXw5PNSREthCc8RbI
+h/jqtzITpT6rt0nstfJLBfkwMMXADJZ7JtRxXLdlO0rS0OxO3y+l6ozYqUnnF8n
MB4nGA49cZ478aIe/OEVog6Skzwk7rUM/U9rOlxEKXyeMR+1njz4Y/c6wiqNH97E
p0jzVTpFxUFZdoPLHfIHGakcke6m9IXuixvT3uwdkvW3V8Ail13fo4/m2CehPFzw
`protect END_PROTECTED
