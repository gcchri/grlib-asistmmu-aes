`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgGJdoMVG+cCGbfJ9kCwV33cC/hA0ghcR6TTFqTNcf4FsdodcAcv0STpt64usxsr
o0bzijNa/yJuKbYCFZsJRCt1A1bJadaeLVN9ndMgHyWRnFKVn6r9DKR17GacM9mW
OvQ31kS6redi+DRXS2qLLvWRBQYPy6rp6f9a+OODw5oDzJf20CR4BIDoJfw0ZwXS
XLzXG2V634XB9yM2Y9t/DWgjRVgAoSsI2nltpID/Oeppk6Y1ytyqU2j3fpN4NESt
Qaw3VszEThg/63xaJGjEtPg5L/KA9NX2/1QsuGstMC+9uKSw1TRpDx9yxp68Irz0
mY00XGycZvzuUviG+31VPLcuGeYQokXajuvTxWgk7OSR4Xgz1CK+uhOqY9ALDyiB
1DHXeUd1drWYFOpIoBtYPg==
`protect END_PROTECTED
