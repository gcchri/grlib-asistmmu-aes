`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+SKeA/Tdj1jeH7Gm7J5KmGIDl+On75I+V9gNNDeaIRRXMzlscT/z4YCQNo9Nwrik
qljjs8A7QwEEKjaoeteseHzBCfE6zRleOQiQTS5FgHsGff0pvUPYyM9QKFGRKu9d
hRvvwawODceJmMc9uhZcAA39kr6E2dhLakOIuKticqZB0y++MVZLTbmVeWW5gQlD
QYktytNWrtn/TkLU+I8d6rP4lTgqHI5VWiSkE3/6qI6rIgGuJJ1cuaTWVDIGujiF
4/g1wdiUqSczjOfKCGfitBOAzQmnjQIw7YzkBTkU2yJBcDAYEzmDiuNeujeOXpFN
1mE/Lt7+q11iGcCcM3oVdvOxITPA4hakQjStqzFtWXfK9nQr9wdAiFFfTAuCQe+B
mZgjSQaTBKh9JxD7ZDdhWzCiq7o690iReYN1IyVxt3L/Z6qUOAESxqc4Ignoqrbr
D1ZuiLkw6f2Rnl5fZymRadF7S4XaMhvP29v3m4LCd91KXmQ0T9O00ueaYpc2RQuX
dZfzZ9fjz6qPkgzgxG+yUwVPxy/SC4iTqeVedXb37bIFtmO9ACu7G5sXJhdAZ0og
lZ42/k9UxcC3MD+maiv5ZJkcJ1Zu0JOVQt4RtkEohtaDGyeNSpNJewcdRDD/U08B
JY63bQBz2cMEKIXtaZdKkBsYXx1qr897h9e4HeDUuRz0q1/5VyEvM5Sgo2XeMdOg
SzrwbLihx7o2gqTxqo2c7NMJ2u8HguRJSgFucOBJ2b7F11gTUb/Bsh3N0e/QmCeY
gGnqF2qQMkdKWAzwAIJLP4fAX2KhEU60fBJ6rz645OmpiCI2YT0TTk15eYjUYRrA
GVlyejQu6q07Ci8GdVUecSTKmT1bkuquJnTxkWK0LafjRsL2v9HxdOQhzBYEoL1B
a4Ff9jBxoKuL3bkO/FlcGjqTPv4TcOZ5u9rLHqxxrHGhukym895Nwmw/BZkrblo+
7FRxD5Ww8Z47oSLtVUsZwSisFkH8uVmETWny1/ZD/QtdV8y9xfgvTxZUPQK386f5
`protect END_PROTECTED
