`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+cuT2T0lCDVtn/nrssLUG9p8Ak3JqPjDhLvkRG/Em9iFqL3W+xjS+0Nr7EREPVMN
0pavP2mm6chG2IRqTz1a5lRZOBiCYQKJEUKd7shJMRy7mtlLE2HObtB1ATZ0r+zj
EevUTWHiB+50LICv76+ILAAHfQRRb0U4sEgRSvBLU27JMMcZPUjLm0csTn3at8lQ
r1qvJzM4U8/UsRm6LUbva6uTQfhBtI/PGxQqTd4wb/wbg9kaEAv9dwUjrZ7SH/Sk
Wwfb6FebkXyJ3KBVla/B1W3d3Me4kMP20qFnjeDzRPYjeLsfI4nIvVFxdw0OHL8u
j1+2tnMJad4uO5Q/J+TGUadwyHjli0M51+2/glW8LvTGsLUCmrrrDqWNx8VUbWZT
2XPv0VaMNlAOjlFWCwHrERnFGINjEz9enwGZZtLsEiC1pzcIodBfA0A/dDxx4McQ
6OEgqk7Um+HP2WAirm28Wv1/h8nlypB25qTdkiG80tU5LyK0eSgjqyRxmT3SXdIZ
mR3xty9QAD9wrUVAJXuLxxd9SduSYJYr59Zn0ueZmLQglGX876Fp7Zg/ayn5oW/S
1NT03fnDv4ouaj7ayS7O4liJKKZ2FPwNzRhkUim5CV5gtYyaYF6YFLlcRo6RH6e6
TS6bO03sx5BDXY6j3O/PWw==
`protect END_PROTECTED
