`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jf/KKmtFzgyhyVnLXZsGmwvNd119mdQ4dQE1kcsr7cWhl4k9sz6IXsQEFG5zDJvV
8Zu/nr5aMdnNrAdpo1BTdYnEgIxLDZ6y81W8ftuWuHdq6MzBjBBercwdV02cYMuW
L+kSix1mDHVekOWK4hszVqy41Nfy6Mvb2WIlmduCNCVeT1rT279hp64HxSrUI9Tw
+/D2gLo9sVKTmDDNbUx/0wc83hKPyH4mH3/3ZAotM2azwwxBPSGcK4/9Kjs12qWt
QStwPGT1cxT2UVnRKJ/xxO7PVWHrdKyoz5eYmJ8oPo29sg1m8GzIQAREvBCbRX5u
TnqC3aX/cX3rgZLi/H9RYvJy546awQrTSC7ypd+owmdiEZXQ4rsfp3cRA4h0fsnb
+gV/CRiNzFsrSFNOhX0xLMci0eeAyLJi2j71NrOyUEzi8SEVbQYKaIv3jDRqknO5
Xy8GeUUAKUuGh34R8rvuIfyH+G921KFe9RHmDgtEzY3CtIXzMMH5gOLlGFsH85fV
UYS/CaK7VhG69JM3nHtF/NoW8a/8RwI0hlZZvuFgLEzF2W6eM8R+6reNhSWSuwzO
B7ekABInI0FC0okEQBBZx88yu7ooT1yjiUG8ZtJRubmxzZzsczVSZkAyJ8xLv89I
AVJ3T/+KPEpbwuz5o4Mw5WEY6+zUf0c3JBZHzZVXJNHpQih0wLmp2VBYvSDNhsE2
3DcS3azgnb5iTXmHZwRRgo8Srrzk0MzuKheQd+9uk8MGSei+mpHzemXDKVZFOGur
krGkJauxoKKT5+4KPEwM3f8REVwxm/2W+XI7eGf/Y+KfF4aaez6WYalsJd2upwsM
NsAytSbr/e+4gbF1idNYK/r74q/s58BbuqgWIzd5RhkxI7I/019N1WrYB0dnrMO2
g26Xps7Q/KqUEBCdUdYRqo0XTxVVU/bAWnfpabNggfTRWus21v0zSbaKyNKGpm7C
8+vv7e5NHEA+U+tgzaufMv1JX4mgyiD/6WXqWoNkKkeokUv902IjVsRikpZs4PnV
`protect END_PROTECTED
