`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvIvO76KnsnuyxkVgKVbMyzP60FHFXtUL1+xZMuHX6F/KH9Rl7oXN0su6tIKAOfv
/NECA7ID+YZGbcc4vrbbI7aBpu3DUbxX9WtE0icw/yrf4hW+zKbpznX8o9y460Qp
XFqSm3BHci2L0FPraxxasgSGJEwafxCheoKIlpJXVbeOXr3pIaSdkeeNRUJGOT7u
MxDuOPXZI/BFPjObOh2vDrhwVVOh8b3ke7PzzfgDpjD25q8aSIOtzB6kiTCYPzHs
A5iVL3Y3D7vDy8tWosIhc6rYoYuV2nIg5/sAXlN2zFhuoEtmLRDz4kI/UshtYP7Z
RVSuTpXNy/DjvSFCjPWWHFWodbAyFhS3YZRTpaAT+jLWNASerCRPnLywt1NcpDog
JH3Aq7VobSXG5HuEVaJZQXIagmOZvTrXOEwgGHBz/2u+zzxen1nCspJ4zSMf3SNs
svgFH9foXTTUL0LMXXDelj1ipCb7EAk5tVWyYqDQCte1ucY7bRONvJTuMzj2PCXw
bwF/htL/5LF9WkAPuD5Y0gyOQau58nJyc4Scv4Wh/634e1Adkrtd08tvLFc45n2X
rFKBcVu3vs6O+E7kGq2JcWrEFtk0VYfrG+baWMvYQdpD9McprZ7rkPwenzwI3Onf
KITMgX6GWdaLSOb/YLrBKQ==
`protect END_PROTECTED
