`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50yT0zxLmSCAfmyNwzyG+9GjvwxXsecZuvEKSFHisD5+mlEnYor+pLtAqOed3qTY
TK+V6XRUdERKxqqzqU1tfViezaiYTSMyXRhExDQRVaNN0pcfOS9cojS08tKaz5/E
qtbOMz2LHEDbtlaAujuBBiMDUv9RnovYJ6GPjFzNF6qJk7dWKnjysZrI/XxPTAn/
YVD/DJjqHgOWgDPCSukGcyRJiASoXTd9rjZ8KtLkmqjq1PCEsL7jQcOQy1Oxf25L
7USub+BXoiZt6iCLv5pyljEAfRSi8Af6/UQQptE0ODfUzTPPTN6Ki3Sz0yfQ4Nlo
T70GeagHAa5qaooajcme7p4Gii1bKUl5t9ssJu9sDdbcYKaWzFSkQ2ywjw1HFVnZ
7M94t+nAj8V/uBTBrlITWBKBd8mPS1JSUt26j9L1Kil9Y5q4IM+vVOYMa+8c/Mzo
rGzEXEcAOUTx9yov2i5oXfxjKwUGeGnMdHlrHycq4ZVKeM+ki6HMhXruU2vzy4Sc
pL3nF127xFYtOopGbkTWaszgWfwQcsP0g12DGoENyqMcMY0K3GEplFromh6Q9vYo
dvMxEzE6vjeNsSqt/g4RmREFmnNnBsXhm790PTWWKFN3S5b3huojixVXZFfeh6kU
7rHGigR5ob8iV60lllD43Nm0diwNcdmi7zMFYWCfDTlFqCIy+4ywOSl0X1tMl5hk
bIzZVDv6jtSVROg6Ag0jnjCb8HA1W0Kbl5K80YDahJfout3/TxPWaCFBOumyW8Xl
NzPffkYP7j0dVhWvP9V8P+fxnJpc4pZtDNbYyT+8Foy7ogVV5ESgtRpmZu+EGBJT
/R0b3Ew8g/Yek/tOW5tNtt6orTIT4p+VxlfeL0OS1/933JwyorFuoV4mBUMmI0qp
1BvgQkLq6896Va5Bk0yyYuJ6UHPxgzKUqtgBvNGEIdOlhkEcbISn2HXudlx9seqH
wZBjSrLo+0liImtwljRNr7RO39uE0bI4HHltYsX2EZhvc3Tj5bx9UlnUvkR0+yjA
69XJ88UN+oWYsnAN2/fRc8xSS1DUjBNAAyoKgKS89CHcnuNc8X/eJTrs+q/kdYdN
B6xWbkOVSMJairrsaAemHJU5j6hRyKgRj4u4Vbne8GH28n/hP03PRUW7sl/LaE0l
8o+PGsRbAnokD77/Rntj/s7yjP4Gvs2ezpvQN8MxvUdeJadnZkK1CbrUalX/g3Kn
RxPMTpF9r35QAxkmlQnLl2EV1mmHG9EWNApfPCfIXXLd+Wcr+XeOEzgHPKbIZ3JR
gMbRAjM8dsO1Xal4NdEWTrqeRKXHsfdli+eqv5S6AyYVbmdWmY7+MzRY43ifGepd
euQcxrgA2MvlZGsiag/I6eUJDTPImy/w7tTC3UqWoaQkXNM2GtSoyHWIjv/RKS1a
CFcGxNr6Seyds3t8bSJGqat3tOqdlXWB2zIeMCPVoeb4amAQbDcuvvPgwX9mGmR9
6kc/UbVdPoArzSXfxaL1mQ6801lkVryzUoAiLuPv25riPVaQ/m2p5vv9YiwvOMR2
ElT/LtUF0RYE2+9X4fAu1Ihq6VhMl2OQIzgZhAlCUhfbgGdITYGeRiqKTzTMCYuX
E6l5SuEflNy2B1rrCrC0q6Z3v13H2HfBMtaxUU1LgtetB4Ll7RnpdZYpQvaEjlby
+rzbX5umUODJpGjAgok2KFEscrB/0XAH8SOSIfKjcuBiWtuNP6s4whmKNiM55rNt
GSpyW47BgyfSYn26Nyva5O/hhdzVnjytMjpz2hQrTQHrZ98EnVodG9CqhyUyGEja
UqytsWD6dKoIB2PLHbpK5pV8WIyf8Do68eJuoeqnuh7yzzl/x3DnuCWe0z8UdRQ6
V7ADp1qQxoHGRBSQ0X1Kd3OdjEelrPiPqby05tY9P5QbG4Wim72WeNgt2/tcKENV
hyb66ivYXykPXq5m5iDl+WhyuURH8pzvmED2N8+kcupUbTv4+oOVjXnl9WsOuA6O
ADzrFnkuvpw3+hiUPvn0PcRPbBYCib1wEh2aQU3SOeA2JK+1ABP05yQcCOy5RuMq
yzFugoKLRIfMlkECVsUQGSSCS8iW4+afe26jZVFschbVoO+Y6H1V1aOSHVNKbiqw
dyn4akuJ8+eVPkTfEvTZhgllugX5+JBo1GxAJ9N+vLMra4nCbNK54byhvPsl59Zw
HIwa75hKUSlesRdEiPNoFH+Ak5X0xMH33wcROc+llnYz8mmSjVpU4h5VXzf68tGp
u7oWyeaUlncgDuhnfoYeQGlZpJ2RIblKlXsWQxWdRPzbSlMkGjk7aUraWG04MpDA
3R+t8peLk/+R/X7FabzsJsCFCJQ7XtQ9IwC3eGBDmIJPxpZvo3Imis8PtZ++MHGt
lz6nRG+s73qaxC3LtXhB7wQXxCaW4ivJgmirZWXMp4Amq1VKxPzNFkyniurt4rmn
koTIIpOP8oqi12zA+V/XHTJPksENYV6WL7Cx6zFNwqRGwTxAoiVs+sHzvsh4x995
2B1vJZFMQcn5UWJueBy5k3zEAcY8/AqQiVe85oTCtJbHi54wOFmXSIq3VlLj58we
qSnz8Ham+J0h+TxWpnR05s78Nc0bWuQoRVlRbqOgBiI20QKPOXdG5i/fLQBhs1di
Mr1++KuzguNKJh+iOP9tbILY1t8wGFxehHfLpILBxyaMlg4rMjCMUdYq1mVlJQKU
j6qyYOodqoXapShGKpEmzRj8Ig/eZlIOPN093VHk4gYxEZiYtfPytbCNF/XulI3A
oZlmTEWQMqLSP9MkuTMLJzEErg0Skj/3CwmYpCq1JtAZb/IA2c44JZst1ctse6PV
Aw5nVJmO22FZsEfCFlfNIlLIDM6xDZwS/B+oH/bY9ZYIhczJ8GQe2/A7ra9mHOqm
ZC0bZtizJicJUicRjL/QjV5KQyEm+xBQuNjhGuiS0dqmTXl8LoH6Zx7xAi7jgWzB
mGDE6FKSvPwIuyliaggREToQNtMqDJh3G7OE0AodmOdP/p0pltL6M6LvOreWGEjj
ZOP1Ns5PQeN0+H4hrMtM1hMju5edBKFqG/0CJrs9Dh8QXkoNYySgM2LshaW4aK+0
YKHNB9h2aUG/UxdiTpH8vSdBtkHbvgFLl4GS0dMrUfjhsEK2yrmlRUPG8aFnQe3h
4hZUJz1ihAi3FniZI46vpeP8DHByJCrVjhUzqRM7SPZbfs3Wvqwn7wQqwChWEDfI
sV3bMiUBZNujKr9Cl97z0VjP80vQHgPlTGbfSsdYK3e/aDoiQ2aX0QDihA4Q4IUk
KsO5blXUizobyURcB26rq5QVdKPns8yWsKCo81n8ioCH0l7NcB5tO8/RV+DZ1STG
YA0r7tYVHoVNXkyt+d2xqBXM7EkDrfD+9geLgclFmekCLWEwGFs+Ketm8/YjWnsw
UB4MRhptCdqWv+gm3d5rBF0zPVZki4AwmPed3+CMp5cqgtVJDGiuyyrlh5j0/2AK
va6VynJpJxt1m7liG9dqqjzyqwhI+7RUuPW/SNXb6Abk/f5/5EoxMYm9D5HgcPog
kbOtcVbmwHyYdESF5ONcZBC/c4dtB8qDglW9xhXBr7ZOD6NMPMSTnQQxoEfvjYnZ
2B4PJ3pSYCnUJNGJD4KLUmYq5zTYSZQzKkk4yUAjWgHR5F+cZ0U6+nqK6YW/jBao
tIrexnA4YYuwwsm45M3mFUZJTDu2NcgAeIRIjoeF6gANYxBUVA75E/pDnNFuC/Py
zgFIVzzl7AsVe7NdKHq2pgfAzVq5DBrwdjVRt0VvHNKNn2oRtb6ypUf8c0yEsYC/
+TbJ4WJ47oSBxfLO7HpcAUK1+Sqjybhw6a4tSM72Ujc7q5rLdHjTPjQ3JleZLmJF
tyaFTUa++OwTaVLf8ykdUGm+0/dPxAV/3ttFaLbjqurqXAZagDWqC+V4hYPoQpwl
q6q8kT8ALsLZKJJnTvkkL3BCE+e3DZxNXtjvVvl2o1PvFV6A1Ec8MG3UIxKzAbb+
uN1DISMAKUEOP+CcC+yNtp9g4VjNj4i9PH6lWlwzfLRVgG7bbhP3PaQL9/Lj4Z/z
MX1A34kem3iDUX5syByOMo8QtLCYFyYRzaWVuN6OBGaAwsZQ9YpUQq2avXGg11Qv
LK40m6Z+FyMGC3YZIHh/9cGt+GCQz9IamroZ4Vw5cTv/OlKyyuJjcjulId/chq8m
WVrQRJqOd3NqPMmn0Bw2WecWCzLVfFUcS+er/1QokA/55cevcsuU/E3PxF2a2cHU
pJqKwJUBisrifJG8t62UYfy8NLpJTI70L5KizcT1ugnd0riwJhaiRR5Y6Mfvo2eW
ZoJ2Rl0mk310Cr/u6aD2deCayofWpOo/RQ40fuaKN8VufSCk7KGujzw9ClxOWVs9
0lGuVOnXqnd543JpvttvZECyIHhBdOMfrlrSHE4SCuswrXFw8OD4z8NhDKRGwB9w
D1fid0kQv7lNoQLIVulxkSx57i6ZlzVnAPI8wv0NTMa/tiA62/iyIYhuxRKOyxfH
jixSdEkyErF82W+tTOtjk+NoRCiuGQw7x6KjC8r70cE=
`protect END_PROTECTED
