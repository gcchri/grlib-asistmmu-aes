`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q94r9bjmfZK9CyRQCi8RPdtqF0l+mgz0kEGCqSvGoEoLnZ/ni3MGl5iYxvRLJSiJ
zncXkHJoKyXg32qGmWPrneeQC8+oCzy5ha1klYfdofVmtNyEtV3IqeVNH1PYnCDw
veXs2U+U9Y84W92fQ+3nBjFZnO3tnwcBoryFlUyyOVUKNceDjnjOzECi9L7+wU71
jw89Yq+bXcYbkkYAL01Xe/TvSyMQicth+6ixe+dJM/sqo7AiMNBaQk4uN10VXEb1
ip3FXvbwLzz5V5Pb+6NkarzAIivG3/UmS5JZGAU8gNsq+LIT+fHQXI42Q5Z5fYZY
+eGzKiHO3lDzOyXWxru6VvWXiUBXwwpI0kD9Y3Rde6Y1S1zWq7h+vxys57RlSLWe
fmjG/CZexANk/O0uGdZr28BQmceVpPQPsFfZ7WGlz5omvCWiGj57N3plG0WZfa6s
`protect END_PROTECTED
