`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3VbG3mAAWF7buXbgJDpNqBwgb8FBU0n8bk32OO1q3sSX8eYOkihX4CM4LiTY53Ki
fE5+1Flc8oJk3hqugrD1HTHOcAkSPQ5tZaBWtqN9ADOUqVI7iEVPwBT1NPEBy5pS
Vb3PAIt9PpN6f91Czocu1orhBeMXYvJSMb4LgzATP2+L8YaI2JU/NPqrb7EjfObV
A0Sp9f7d3iI8/aQROvhn6RsSinX7YuPXa//AaZ2FBplx6TNo8NEYKWpuHRwVOnHw
UkAgwEEYJ/udX75yqmwKaU2upGo47pUUyqUb71Hidr1uq/spXdyF50+IMKEwOJmf
8Too87OeQ8GVWfQkTVO6uOrG8E2xJXGCPzpAp1X7D3Kw3oP3Yg6R1wBQvDqLzqIB
oD1RN/txHu2ELG5MgtN1kk1oE4ZvmDNRgE1+IJyRPSR6sz2aqpyoeePPt/UlHFbM
FXXurcHsKO422jGi/bhcRv3BKxFaFPbbJjgPUNui4gKvukekq+8k07ysy7Gwzupy
7weSrLftQjVoDKD0fSo4dxWhVOV5bvxY+4hv0XlzA4W8yzKUQfVEwVZmF0Ax1yYE
0ItEngCGCe6BwoBOKbhttxlM/WkfbJonpO3xdi3hK7T5xE2cfMzMF4jMJagCpLL8
FZbO1r/kxkvrVcC6mY1RMK9JUzL4HqS1MQHbRAXaMi/Ho118O68ix/WwqH3s2Snn
N9hHJLqRhTr0hWJ2wibtHVAFo/af1i86XbKJcPIaWSDntTw+4HXh7ZCUaL36Q6+o
4agWp2sUTAXED5Eh7UAJDeUiqpg6u+ttD9YQNnlwGjGSkZxzW6s7gTCdVrqJVRjU
Ppa0ScAWpwI9xS8IYTLQ7w==
`protect END_PROTECTED
