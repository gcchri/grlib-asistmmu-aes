`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9VxvuMpRY+05RSfLQdQLlaWloovylb59kPooYP+Zni+q0/rwusu/5SpIQaN+qK0x
cDTgkq4E8aS9vBklPvAqyM2UNCulZ9n7zpLlZQzs/LYtvoR1sdIlHiUtdDDgZL0p
GWcnFq9/oda9tNwQxVXopDAcUw+sLGwD0+IQXcJzZrszYgkDxPQDLEOKC6UHQzam
sdmcMf7fiY7+ounPalv5OayjSSevDTaMO9GX4s4cVp20OhIvE5R0LdkhDF3fLH9Z
s76xfsSCV1FSmdKanULEoc1ktvs+wkVHXmVCr38lQvOKMg3WlZEYtxUa4zn7oNpV
TRkbA8sgq1iUA1QAPIQW6VcsXCHxAj6WXdHF9OIfOcrZihp8kLZJ5P2pEJPkLbGB
gpydtWP4X8LeZYulkmfBYIAUlVwWl5Jl2jsESLI2TzvV2DwMVhU7j+07Z3DajtM/
ORpD29LhStSKCH506IKsltXnupzn131g7YsuxMzYyRYW7kLfEbVYYQpwN17hYJYU
aZ6luIp3rkQ5jOmrzOcOFifJPbd9Autci6PQMrAX3PvvcpqRrVvaPQ667694/Xqb
zDdTS/wTOkm+n3sCd5aiTXEUcFlI+wWzsnIjlumKtte7fAVJ53WoiQ4xT7Rsc+r+
L7aqz9VtfxpzYK/pVRXeLQuq0GXVnjduNa2hOKJQlQImnfVNA0pdvgCj12CiMme7
2oB3KAU6tv7HBheZq4VNLVUs03rhLKdcMfkw6YeZuvdAy/LB6oP48mYjHOBPifK+
sZYhUChPyxsrnM4Mg7mkH0/dj22FaBabUspolIH1RUHqfzy4jgV3orciEshoMKVo
OzGjmIf4gs/kO15kSguxTK/NGT8pxHOv4VHkqDiaK/Tn/G1EU1J3wUkoirLEgOOO
iGysgkfMHFh4mrSFd3XAtsDJc+uMLdsmTdj+2zb8y0Cepp0bo9iZoqze9Mj0hltH
6tB8WLGLSEburMu/bB9ggxOyn5JKltgMH+TyRRAWQAl1oUDVuZfVHDLciqI6vOBC
nOngPSzmIzF/hHE0Kj+PvRkuWjIMwxbn/p/XN5qWhN2CzgtRbJVxGnBsxAoBkcH5
crrsUW96TwtYA7DkSWo2tbrTlSgSl8VTgR2Orp7SGdC0NuwtUJM2TSnsCBR2ktwp
PSMdhZ/q6DR4yVwbGNU3g2uPabkv7xN7cws6ITdT2cv80OmBt0wZ86Z/UZo2G/+S
FwahQJ44+dA96y6uq0kG23ik5jDxH+WZCGmKVBjwQAmBTJpvHI8nUnTZr1lfIYeR
j3JXlrD7rDjhXU06tE74wwl1DQhJLeiLdJ6zbEv/HgSPbyGoIGDy0sEQ/3lbNCHT
XFrrTk6nRMeKaNuvBHwwro7/Xu3kVO6n9OiDaG8mRX9Xej1w206321td6rOGcKl6
`protect END_PROTECTED
