`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TBwbjxIT4bOkhHdgas4Pcpi2XZ4Ycaai763zp5BgpFd83DOM2i1A6XgA9Jf2lrBR
s7QhBxbAMdqFA+P+KyP2fJn3P8t1aQjHihJjcGF1TLy/535bd5PYkR6qCD372B5M
QfQaXKHlOa7KwP6e21bQFtxZ03U2GyOo6L+GxNxYm3J+8K2lU+b818v8mZPcjrU2
Xj9PmpqX0ofJQt80qSmWch1W/1e+D+m95Lv0PDKo1lm25C2SNkwSGQ61qJdrHC8C
j/8N+Rltm/BZ0vB8LQhUnRdF2Xo1yeVLhia8JlZUNmU1e8UaIgBhzoCaQryomoj5
otZSSRARPaygUTHfICmQSg3vuza7Fx2ax/cEZo9g3DIwxj/WVLwO2g8KGds98faE
hpG3HcxV306LcqX84N2uNrYcV/kh+NGhg3yDR45aou6vBvHrJa5vra5nonY98Uaq
ZU98so5awKcEMSYlaqmvxd5Y765MGqucgadnSqgjLcVzFwfv9FY6I6/vLxdZPEVl
9qOQHA6vUct7JiabO6haA6CLPcX3gCLiViLMPH12dczXCnCoLXDNYgPvDNyqy99N
Y8zuK0V62X02PbqQqvBTmNOb+fln+mpV96y0YK7MkqG0K1KYIf03V68AAE7GIrE3
pJnEFkRNMO8uI+2DGOIQ67znASXwzwqaQJA8lOu4qb4LCF+d7yAnDdAZKMcaw0Zg
hx+ySq+hoP4xGvp9xBVt866TxhuxYXdDcKurSYwf5c+ZRnwPOeJMqCgBgiVHQ4/F
ooXHVudGTVpHIh99mSQjVg==
`protect END_PROTECTED
