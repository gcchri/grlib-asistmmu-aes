`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TDXINNKXprQ2CHrpqI3bt9FeVW2ejKeXBkxRD9OJJKb3ANUSF8YLRAT7t+RDTQlG
hTyqhRXjh1sNy5MAe/ZkLCJr+egHV03xSSdSoc1AZc6DAhEwj1QO1KFnWIvR/tvc
WtxQi54qbg/HhahGES9575auXUsLCNfjqh5TI1uiDsUpPrpopJaSPmQnEGBnHXar
RHFCmwz4C6gDXgDDwzDCaFFZ6A8eVSKfeMifdbivBF6EqMdomrcJvSYS9zhnoTyy
kv1CQ3nP1sLF4H4ew24uocB4vnYxBdIc64t7bHC6ORDk55aaahF4SBknwuvsUU/6
agaTNrt6wc/wt3HLnKeang==
`protect END_PROTECTED
