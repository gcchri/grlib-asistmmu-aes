`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+LSe587yS6nPVM3FTo48uZxlguEswyxU8Rb3V5t/iDugUTV1Hz4w5X3uS/rqhL9
rUpowYxsIojn0ZhHbr/tV4z+hK/ejQY8bLAUtgey4J9+JymN+kD6X4psFLbqub3G
EFmo28WxS5lT/FfG16TyteL0UplxoyyH6P8gblFeoTOnp2oxZdiER9sywd73iQlG
+uwR/nRA3YddL0TQSejriqVtU/wT9lfXEtJMGlMshRr0PO3hNTraKyGWGWjnHfJB
g4LNHf+Aa6rCXJOA41Yu8Xjp3KXrek23LvBiT6B70/YxxwRduQ3QQccSM7iux2J9
Sk4VqDgjZe8/v1q0BFdzT/L/rXrJts46eaxTs58D7ZcYZBj5B8pqwoUV7ehvd3Ec
r9OlGKQQwX1d4w793jPkO9wjhgW2eOE4xz/jTw/j2ck=
`protect END_PROTECTED
