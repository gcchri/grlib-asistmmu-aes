`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xo0nh3nLbRQP+b3yFYhnt/gpvHE5Lg8hGFW0PKSSigAUg/iDjf4VbNOO7jMJ2LUu
gvDClrhvG1DzMYzS3EHfLpD+IRS8bgtMdy9UrOl2Tx+OX4QETtD/B+o0qWJLbSHJ
zVMwlQGMtsT057wGue37qeTP94syfs0/CnB394gilPLoaI0BCi/fuvlHIrVfIjaN
F/MHf66r5mSp29DAR2AwqjEb+pSC6QudhG3JbhngGJm4KrUFfyfCDF7jbc6inqSU
T4bKNHRyu9d8BTz0IdDBySSE28IAPkOYsnfWipIpHnSHLDpLKDCfqtdexxbgO8y0
y/hP5p3w8ZrGTgSnhlwreV9Cds/Oc/tWN5ky0bWO2n7DpKQrTmkETh4swAI386Pp
GrAqoki2mkczKRNlZnt/MgiUNwsqeuuKcE49MX+KbeM6O0dztYSErAcrwmn8yTDh
RbUf80SAFOu1Adao/c7duQzH6LyoEmGs9YvU0IB/Vj6v47VzoCjjKA48omi2X73f
mFMWzWetMn8yX8jyodgws3cpo5llUrhOSyOw9wjZLvO/VbIe4ntqq/Em/Pb/Fnh1
DeLHWqCDae2gVD4DN3QxMYmh8gAaEWBLx9MQ1tN70J/AjBcCk+BLGW8DstHjzT08
HWyQy/e/bDDGLop1DriT9AUhCUnuU5MALTHUPUWRPq0YNi7hC4Ynd+z6nW0D1IHr
eMJMa8cFt99MR3DiDZi3DJlFoMgT0LFExyM27HUaAIW8ccbSMcj5Z+CFAIqgU95N
0SrSsQAw28rbKDowV2nLR81dl+HEyY50N5Z1FtA54n+OTYIGOWmhESOuO1qvNNrg
3WIUsCxWfyb59Em9Z9KELidZcN75E5IhYFWs1871SvcddTb0ARW2quHCA3oC0sxP
VDr9dUCiLopdhqol0eepaVfFJIfYojUd6pN8uX60wiSLPTtF41NU+pXmXLPLogK4
u4ErtV8XdCHphuFsjZS4iLzyANGU42UzAeTZdrNWbXdEERkzumDIjcCfACSZKVFM
Mo9R6fFWT7/0aJ4Dg4qBGnNsfWjvpXpuwbVD5jlovjhb8w/KwLegqVrpV7tfi4ZM
Vt3VF2oeDxCNg1YBuKOg8VVXDTA/+YidcaVbAfmQvY74bbmWjRFgbmmw1StVcX34
3W1vOHotRrfCv3xPLZt+icVzRXqCkVUnZJsxexPLL+NT+n51aKCdbUtaNUpHuwjy
+j/K4poolOmvoSAwVR54WyDZa/Lpi32IIQiMWIKAfxp/KZpwf3lZC/4cu1oekpaF
FYCWU+3/4HBbgiRP6b7q8h4ukmAbSJDtXplcmpCIwF3RotPhUin3LFUQ+AWIDSh6
JluqyTPu7W+Ks2a8fXPU1nwRtDgeGjLhx7IYMRh0uG671KH9rHEInq2HAOKziKOQ
V9gnB2wflHrDzKIb/SiRkJY1jIGuC6IvSfcqC0f/6cQKD9hr8Jzl8U/hBMMtSi+H
DP2Z2tYRhgCsJ8hP5gpZA+f3klO4qMO0umn6FLPGSehSmO0aosVpjZqE/rI+mcZ2
TcH3fjBV7z39Kcp+6iaUVBTsLs2ipIBoEMKCKKY/8bSaka73pQM/o+jKlxoD1+b5
GfzEh4gFXXxNgABKJ/eZf7Jkb8F/gbwHAqaSGrtWHQ7SCVUSQFt4OpxhgbOj9wPg
q+9uKFxXi6wE1N+1blEGB70BJLXzQz5vTpvN6mcCWn4HFbCYE3cuaQ+wk/GrDg5P
JgElwEBd57kQXdzatsvAqpzURvs4qxD50npNX3Zm4rsq3BbRoMf9jAfQr2UJqNt/
x1+1NaeZqGcnZ4iZT44K6jeMf3Co3qKGe1gkffSSjJ8VMzhO+tlQDZV/pVb5cDcL
jCQHv7OZoUwCaNNSzN9uhHAVWSuomhnLc5+ipqXt9He9qkrHJc6zAQVtL7riFp+i
/P0eJbebxMMSiNZcZSyVyEszBZjQ6FNEs4dtz3SbB7WGQmjHDS8AYCok9wpXysQd
r0ekOQtvFL9agvnNM+FkDbiaHSsFIuLaJBmADkwNw4mnm1S/TqMO3IHKuDKlHeJR
qw9jbmbQldLpaA1RpjwXStiNzEPphfZTRvJsi78gGLEpCR/foPyRAv5tfCiBRdBL
Z7agx94GTmJ4R/jb7q0BAb4vzGxrHoW6kK8539E+czTjQfq2Zxiqw4BzA8evuFqA
NbxIxCNgEhadFW4WDh7ymDRh0cs2v9eGBZgi+6hN9OWe96+cO6wrS722aD9VVCFu
Z1DoTHfuJhFnGWvLY68kp/adaMEyNzJpgmajD/pmppZ8qYC6hr6GbqmyNohTXLVw
`protect END_PROTECTED
