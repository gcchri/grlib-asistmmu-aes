`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cjqQBXahLnkMgLNPhZB5gBXQ/L+ZFncf+wkiZxhAIJRS02chN4E9orcqFl/763zx
6hQGR9wo/eX5wOjGkzkAxAs3a5LftSyx+V3gvZmr8AVwPkskMrKffUz1FieNkQ0+
t/bUVTo8eKN4sdDfsl98CpxjZl1BrDE+qQ1NfCmdsNa6Um814lwPloDtWOS+TRLU
ZPAIqC4TvzOsrG5NPBsNfKc7tMNwFAejqjVlt+01v9lNdf6UZjvS7BHrhKC8zcLF
MeuU6shJHcZP9AzN7DcpCFcHLIb+yiSUYCHzR1VAqnOfiC7OkZ/NzzOi5FT5642s
2+p7cS4UMvIXOZg19iWciDyAn9GJAEJO3NgipZx7PoS2O1iEZF8k9Tz6r44eXnUE
rzrtqkWYgGGnBYSBmMugwXO+jIRo86v2jMQlck7eJmmFNjbP/gZzw5cBW6abBeYi
1IGxdJWca+RYVU1aAyj9CcTE6rE2sdgkkwYL+NUWu/9TOEx+G0Wm1ZWM8xatXCMG
1oOu2M2Ly8HR6JTC4L7Le17mi8Adls+QI9g9flveHE2BUaHbZ9wXjJVN+3yg1YWp
gz8TOaw0udxGnv6XHbk8bhl9UntDFc+m50UAXRfuX2MPYoALl9FBOMrhUlK863An
qIx1VA/qAQgF50glrnxZGKWKEcXMy5PQkSQom/JYAa3KulXFiAh4XZIhLxIJWR/d
yjld0Hc/JbPCt5re4PnerBPOaxHOAuxdf0Wrda/nxtzdf2H1+J3oKGxmYxra7yWR
D7vjcPQTqsUU7rIZWmGPVUXUKxpJQhktELiCTkqAwZLLFQMfedISsDLPI6gXhSCM
PLwVN4UxR0ZjkXD0HG3iwDrHpaFZTyrmdwcvaYNegExVVtTpulK2Xkf9P3bvHrHb
ZEb8koFNl/r2uDGJkps8n6iADdOk6zMMAZre9OyWb0IpI3d3F2KXrs+7OfpMXmvU
HSVxgwQqdsZG8e/PSMypXNIdsLBp64OTjpBQVBWcmYujUJBzwoYEwC6zoTPbivVT
qfLnudGZd1EPTsF0ck+Tjih9vQa3y/F3Z5vi+xhgxPsi9w5Uysky+HdC+aq9S0nF
AC3QRF63um8v6mP93TZWUV38pmqOxHrKUCJ6nSERkV7+rVqtMvbhH86p02vxGljq
cRKFtLMknr7NAxHHMSvZdu5J807C1USGGLT3MOFsfJ7WVnPdC232COLjlpOXBoXW
NAxJ/GhN9iIlTaz5m+57DSXNm1thgdftI0Ds5OkeGOXaz+2qSCpk9RQQtxJ8b9Ps
JxoDTwXcGthykDuVrYKw+EGc284nHhC6wrGi69eY4upI/fOocBF+kI/R+aDu6yBv
N776Ict/zeyTYKinyzNQTZIgWgw9V5TYoIt2NSEP60scuEPmNG8aTnohH+efVsn3
bcMW6XsMeNVCqgof7H4txFrN4F6Z2a/lHU650KHLR8HgYmv6QPvuRPbtLNGQ9Wd8
9d5UzYLeZ06gtT5CWJZEUBFJ7T2PP8mzIyMgul/Bg8XG2pBnF/1yYNrJ9bhykv4p
PhUnu7K9wp+T/g+yOtW4tQPdyKvlY+1jlKTkmlsKnXbGPSmoNFGEkZaD+JqmCvgc
8Lgk3Ne1BqIguMfXcPlhWHMlc95Zd2C+O+VpkOiOQuWYsS1Nn6+JxPfmjRYD9N34
MQWTaHN50IBbnjdb19gQhp7DArQIdYO/Aq1G7U4IymaBvrCgd0D0fvjLt4QqIdaS
U32nfNq8DKQkCDKyvHlf8/edy+EGaUYsLGRvCB8bxXNP5+51xvRXesZIQkIqbT/i
8TNRx9sT6PDXvpxEqjD3HiDNr02FzR3QnrEQUhud33EjgL2yLiw7F+pvxPlzmlXD
AGiH7UCOeBMfhRf8WpX3zk2+/1zKuY8SzTwyg1fNscCmFKJ9c76aQ6I32kNxBnZm
3Rvo7DavjBr/PpBXy3uFElYnw7D2+/UW7//ohmtYGovFvjbpWz9EWnO3MZsucC/k
9wNFb4eoUYliJfPWYgdZZypyL6X7zalZG/Ebb7FKDVsWMDc2WI7PMfXZcSLB8X6X
xoQJ7I05icYuukz5Uxfcby48EqAefQ00VN9uVLrz/rvsh/5fEtoJ8zkditTKu9Q3
ma2MB7yKRzjWaGVYREWH98XNIlYMWr8xLofFx9tzqdi/aPW2rumxhazZfLv3Cd6J
NNHT9BeVRUmQY0mpDd9c//2G5i0VHp92qvPAmyAUuLxV+TSaPACK3kCLN1Ng4sE8
Th781o7xej5lHI8UUjAJ2C9TDrg3UN3UU3Ff+YeHQthA4hvxVvw7ZgfaCeb982w3
h/esMbB8cufN1neHTtQblM+bWzqPoabtMVHuEWE0m++zLoSu2387OCr0XEwGCUcj
jBGhZD8GEcrQurz8WESHh3BpYjjJyF5h6U/plKNSGfUnYdqxHLuoT0Lzwf+PheFu
KmsClpG0PsoaUeQ9oxeZWAx9T2d/ZDFLH5M+TCmHUo/DfHakF+ZfMCq9eR8WBTnY
j5sZxcRSs5SCB1mT/GHlc4U0sYag4Krhz5X/AE9H1Bwr5h1zqs01FEcD2HxJmkBT
3k2/9eKvOs/0hjdZebrRRMabGxybjXHZxehgJaDC8e6kMp0PBehz+9koZkhnCuKD
kGS5dwVh+LHlBezAAlswC+vWOiEbENgVU+pWILN9+1cVKeNnJbyd81XcCA+Vrgt3
ysOW3lqIesLrwEJeBgAbARa+IKHUoNzc4PkmOWTn94eTrU5s22xJyTTv7R+sJHDX
U2POmNQFziYzO0knmdSe72qxSKAYtqRVFrwWMvkzIN4OLXgJAL2UOYGoiYyVVN5u
`protect END_PROTECTED
