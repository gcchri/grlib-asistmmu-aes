`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SxLFSJhWkknyea+Y3sgLDwt9tyru8oZWy1OyMaZmsyNSSbv9d5vhOa9W0twfKqmK
MGS2ZH2vQkgr8XKhcv7EadJgoyaUpPFPdiBrWle7gXpEpLLGt/m+YiQqZoSGsBIT
/yC+Pp8zH3vdSIm8vI3ivak+NlMVDs3fqoctBU86GYKPPdWqXb/Ruty4ctKzQW8/
gl9W1z610wTId6X2tBk+P6UvCpv4SWsOAQo1Q1gP2beN5hRNOLUH/KlT7PUcKgZy
dMAgJHtZ0PYlarvJNr1OCUsf0Loe2ZmfIPQa3NyHGreFrZ5fC4SMjx/TzzGpKQZm
Rf2O1Xnknr0qI0X/J7ZDdPLgKV8W9B9xUaRwxUUlRSbkcKvhzyTCz2IvJoSP5YcO
lfRPZU/iTV9+ketQT1zV1GMA/GsVN3fGX8KMid+P0Vy8kLCrtX7HA3wbqEOVGNtZ
VAgdA9ZRDXi7CjXY0AlLvB5X1PqmQMhC/Zga/4JuePdRdKEAhCXOyt9fyKm85Ga3
NUDIrslGCSr8WEC0x1tWAwJxQqabbegLOf5pWGkfHWhcQoTtOlQpMpVaG0ZdgUZW
TlAMY9iubvEkR3fL6d1KIKJPXn/4uVdBqcjR4sF4L6K1gLs96IknwvecGwzU1OPn
vuTc984SkdAluAi4t7sniA==
`protect END_PROTECTED
