`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eaCrbgMK6Udmz2Lb2iR1VtZCOPAUp3pVyCLDZAJSK6m5V7J54iTM9QXAVvD9G5oM
zdJlHDLPOcrM9VvJbUxt/DjvBkvsrhiFHQzDtsUPv9pnlfVyPbR8Ga3kbgPs2q3p
FrNAoBED2h4NnrJf2fUrlX6FOqJZK41ONA9Fh3IgVieqLhyuRkDPbTpMyS4WEpzV
4P6Sp9UTnALo8WVtCnegJqre4DE9UvzWKjbmJuoeJXznSzY6LRFfvvj0iJ225hO/
R62w/jDq6JaUixw5kp93BDoTH1SMhaCKno4/SYscIfhQ24plT87plMBd3R+4uV//
vmcUw4uQ4CA6mA2ARMnAbmQtvlNlfP20YU+M0OQipdFsLFUYSCbHm5OqLXt3ro1M
or5AZKaklygSQBJCma06dETKB2DvUw8Sc6Phvrbz0Ox4f7rfL3Sz1gWvaNJOTkG6
PUIB6heJXnNU4UaXYUMnIro0Z5dUzuV6Guzt1JTGk+kRcOZ9YBFjgTmYgYfgJKU2
aicuu2RIcGmnLuHO1VNAfB1Rd5xnN5zMV6l4AHL4JKgjWbFZzBNF0Qr2WHhQXLuZ
a9L/BPyTcUIRlsUTvzZpiFf+iV90ZyjDuDrdMXvFysZ+cBar7itEmVWQMba8Udd2
6OnNL8CyKUbatpRIQuTU+w==
`protect END_PROTECTED
