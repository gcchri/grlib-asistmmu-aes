`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovwqiULnvuCifQOotCp4rR91BP4dF1gVmDp6bzgWubqXpkApIJ+8HuyyTRJVaEjM
816YFI4bhPgAVioSULosGCEpHDeraTjWwZED/pT0qsBsansnMo0TztZzdedo7o1+
8cAdnQVkFvHTHAjNoflDin9WABupwCzwDWmnXK5X9CJQHl/+cDnP0xuiaaCnk/x8
ht5p0TRDu+zZMO1/LUwPN+hLIjwnBEjWmQZbjPwPPk2l2JLiOjLCQXM9yL2baXBF
9rNxaEo7vkRwU4XLKXhy1T8rK9AEpa0+RvD/rJzhW899tbhH62kJscMP8luVBUZP
utBsjGLKMQ0k1ZG2ouZrTA==
`protect END_PROTECTED
