`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BG3F40y6xRyXLhC/KEQo2XiF59a8Kb3NC7EMF7LJlvCv2H3TUTNlbDtQaX6SOp6/
ay/PbRC0KwHPWrmcCIDwWIq8c5bljTdcMI3V8MjuZFtoN4KhrvFbk+EXMND3d0VB
xXjk9ulsgZyyciWZu/ciC7W5E8PTR+FzcavidiPzGe4pKQCreTbxyNWeo1EaXBhK
2xqS02lTHNf9hF7ynNlor6DSXdFkJp1VpRudKF9MV3CAe7cLKipCt91E0iFaj7Hk
0uzrkssGUAAuaocpdk3IAygqo5JGoKeF+bpWfvGZSuZlWrs1F8Gn8mLT27GVRI95
XR81pWo49daEb990ZsOPeePqtYux7eNhTrTQ+LOR80Jh+IU52FAxpjeEjtUBmrCF
35Cm1mxASSBg5AX3CfqqQOtxNChUkMbcL4+XFUHqzB8jULA9ya+YeuS7f9zEnM2Z
WVFA4AY0bblmxeAfc4AtcYr0vssvTh5vXxIqYTYwj4rUFADtRXSvLHTFyXq2E1CC
De/3bTgpXVEGOKQw/knWzrrC+qgP7d18It/o3WMZgFK9BP9xbK1AEkHC8acfkXae
YJiFhuinI6WsteTCcxmvJyB0EOU8BKijwjilpb0x3vglvvCprAvSNNT9reHLEp+6
nowoJArX0nqH1ojw3GpvBDdpfhJ55UVmb+hs/Rg9CotAY0tGKErFfYaQO652zlhJ
8c9TctnMZ39zM5ygzz4ZHHH21Kmy4eDTSnkQCzo8xPp82uxqXAzJ1x7qe/C8KWRf
7ZzE0QSzTaXryoMaVNLwy56Mn99A2mYWiMIZLUQiXh37QaN5dC9rz7jSAirrCh88
hj/QDt+lSiCGaM0GUY7Ea8PJ8nq+bXO9xHEufQZv+gwdY4Pv48omUahMVny3iWEK
yH4JMoREP3Z8rhsVtEjLw2IFqBOe5N3zXTS0DWQosC+Gpjafxgr1gArS7SIW5wKz
bY7f1sdV/Ggnz8/hYmAUttQCYWdKT931/gQAwFGvuOL8NrhhuJR9pBdCa+bqecqn
aJ0nZLRc170JmclF4TfXOC8VIBmg7YfNJtoG8SWusAQHT2SZm+PrntP8DJ933hpl
pBZf0koApBCdvR7wk9Ho+u9pCuF/zxnphfwhjRDWLD76xJAS19fbW2DFUhy0Z/8S
AplWOGS1ttinph/9Zv4Nufb26vj0qXFhPLrvakXtGfYZwfW+PfUJ00SnfEFwJhe4
yVkhHcC6WUkO6aI8RMVJKTGTw20KsDBWGhi/bQOvqplDcbmuLuX5CIagGWeASnCS
Ql62bBMnZIN4UoZCTrvyy2Ech/mX8BixBPpgtkeKI2K2uQ2QHIFwEk3XaSNhd8A/
nJAgzaF+bqdfORrUR+WM2c13J2zlLqJv9yFS8ENWeuxti0mMY1fU9HoKEPqKKD/w
hWELMvTMftDlc+9IXKBI6AmKX4WXYweizfni+75FkDsTNEUbNbVrYjHVJo/RfVFb
DPFW3uTSHyPFs37zyTtm22pEG/NqYpQ0atcIUpAgGdlmFs/OCNOBTQwp/vJY3pc9
R+hSntHi+jLrbythpdjzsAlM3WVaaf0KPEwTIu1mr/JZkgXkO0nQP1TfgA0EEiHa
so2nEPpgSiRA6fsL4AxuP5AMWG8MjDizH1Egau2hm1IxvRQMh5C4mpKmOBEJsYsR
cNLR48kKCXPWXZGXz68iDOvzgNoj6VTG1QtW7QjASk9SUPTk6J2Pv/NsWge8KN3k
mWOS3kVnHSEvmCaifgdgTIP6XvHbxw2HCiOKrL37PyxSvqO8NZbULgNU+ygSNU+I
zkLzHcap4FrA32ZpiXkzBCT8r9cH0o3N+qrcOr2d9jedR36JSCpjT3a3Cdz+9nae
AQQA0zGfSAfbbKNTFVOp2Z3ZRSnXv2OYTvsUEsUSydonWEme8NkJPFsLdZLicUm7
+P1HRIFAHicPH+mugUdpAEgoTfmw3vtunuOrvaaR4RZdIr0myADX/0p2IP8Ay6uZ
0bnknM0x0AX9bu9x6pwMTIjc/BtTP+ue+JtM1cGWiS6Au4BY/FlTQG1IQES+B58h
sAo7m5JpoPeD+wFb1LXmA/dWvC1Rck3BSMe1yxsTWalllVphf8RCHSgxY/1ImsgN
q8CIsy1/FO4lUhsjdR/wd3t3K9IGKyv/3soBTvuwT3oZiWMOtEICk9jKoBW3mTEZ
s97zXdZDQ/LU5cTjcRsHGOAj31DkDI8B/RzkZfexbkM=
`protect END_PROTECTED
