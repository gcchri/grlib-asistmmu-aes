`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yq/AxHnd3cpSW8gMRYAvXO3kz/0UDZlU95LPC8X1Nng32/4Q0qnPf1/TQCE6wdl0
0EmsOGgQEP00OVQcxwZLXzGWXxsk8T1Sb2VECjhLmPVGi3Lzb4kn4CNbK/bzjyfe
f8VoWqda0D5em30ILFJtNHs9O4Ik2k4ouGep1kk+2RYPgr/7/9JM/l7zMwWBrDI2
nb/yaJ99v1uYsyuQjlSA/eWEdssSsF2z9n4Iac0v5QdRnVZv+cE/l748uRsOQU+D
LBC9N3m5cLna9FkgyPBvR25nLW/LraQO28cQcSJS4eHVUrqDn7ncT8Pe1Dt9n0Sl
ZHZBLsDWB2VWZNRfSvw0zhgbxWV6WZFL2BF3XGLfFMh49Q0a6dnyj7n/r0ltWmIs
`protect END_PROTECTED
