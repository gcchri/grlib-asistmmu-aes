`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dk6MVL3Rg1sAXlcCejEt40DyZN48HN1XXQzW3SRNrsoF6FEVCmdPyI15TnRzpWas
TvSbYP4FOZoeFz/pbl6xQkVS4Bl2q+4u4Z9gTCWzw4Vrfl1a79GiWAn6bKU+KI7k
96mAQxj2KShlEvXwE46VKx/DlKtXgR5uOdpXv2CUgL5DYaFJ//W+GxC7zbAkfGtu
dU6jU51ct3kd5QeHHJsuoPVDAY5KSuMtNUyfbmI2nqEAWTdce2CDCOzNr0xt7lPy
VpsuPoQzhzXpQTFSGxs4zPHl80LS3jvPxWswwQth1TTnQcn7O2tIjxdSNbUMCEB0
0w7Lgt9h7tzlB5Yr8N4rO/viKoHT7NzjNdcc70rVwdSjjffp7M88jibgOiJLYDCm
FD4z53OPtrXFnjuACsu9kVdWqUogzWKdbUYFnyKG/2jqrA5jEXMgGNc3jMh2EMvc
`protect END_PROTECTED
