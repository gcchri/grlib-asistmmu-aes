`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KyhLXIoaei8vTMofR8TrLIgQRiQvQHVcu5BnW5cvgJY34T5teSSXo0elijkuZ/AL
RXd+8ZpmWCu42yaY0yyLRd2CgjckDe3d/yTpfyQQ8mEgELWNzALbMDN/HtW19zs7
GMlwNKnRyVLMDISsW2V9BV2ammWDtwsA435rhoHJzJYxLK9BkZwFeW31eCmKQpeZ
TtaAGZVKUAmNDIyIi9AzFfr0roQmPLS+FBXE2Sz65MjAeO1noAt+CF/JcKwEEGwS
ffL3dpBpTONULU1Wrs0O9L4yfY6SYP+UBfomshCxPsXbpZHqv7PI0luw220oTY9u
NPYM1ojPglGoWZxpdjAIjw==
`protect END_PROTECTED
