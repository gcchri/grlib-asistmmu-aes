`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYh0z/kPGkjngrA9VaOTyBsbhgKBY/u07An++KsJ4bcGRMOUilmB4ve4vsb+bFTB
sHFY4ZTlDi58lAoC31tZqngL5GNYIuG7jM9g2Sw+XncV8jjyjBp1VUcOXEopWHj0
DAeQb5fO1OoYnPbSJc7fmZ/sVq7Tx1kJCqLlHn9FOTd4v6LtpuU9AP4AkAxNbeG5
al4bit0zwy+vO+BHksr9ZbR6nstrrZe0jPm4k8M3ikFLN1iDd/NjkV+nUto4qppC
P7J1PJWNXEcplmMcVy/VC8vPysS/2pSTgek6O0XUedlCX94YRNjcu6Cyi0ZIJMkt
+xA06K1/r/bSWdQn0IXGFfKOlfSLgNiIc5S43nLdzEBeQxnb4mVzb9uR9TEFRXE6
Ij0x9WcNn0qg7A79gdwW8JDEjaUF+FoI8SCBmpU3an1YXArW/Lx/O3m8C0TBXhOx
rChSMoTj5ElPWJl4Qrf4OUtTt6dX9LRAMF5zfzCcHKcQMR56ScV0v21imflo7bic
C6kP/gnah6qQnWnJjY3YnmGoge7AABKDv81lucyWxzXKq3OsEo2PygHv/AzeuKTU
V90I1S3SuGCXP+zTgG9rwXRs2EFRKy+Heykdie+7XtUL5h2IUYaYAt6+jN3vD+fQ
`protect END_PROTECTED
