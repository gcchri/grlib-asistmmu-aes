`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ec45GcmTrHAVXSL9B3OH4NyvL9QKQH/xldOyJ6KJ1KKJro3nYftFMh/xpnmqqgQ7
jMpAcMJcB/PkusaKICEOkg4VOekMxNDmbBCZzStTGYQ30XifthMgnJlKJ9sZEaWt
Iiy7uZTIrR884lrVOLY/HzI6rd50mVNV530MG2aIdWGsmxCOaRJ7mCIjgxzqFHU2
Sqm1z1AOktzc/CAILC0VQCFUIZ34kvDYAyGvoNts5JveSulR9sQ8jDv1uyrBJ5+O
`protect END_PROTECTED
