`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/l6WJBMbvnAGfQoto8icNOall/RMG0TTXoQpHpOqTVhOksLSTcGzlQfhawIkFYia
IHBQlrul0Xn7PwcYzoV/AWQBmh1fBajU99G6FQAwknreG+VR9XsDAhgbps7IWhEW
t7BtEnEJ8rkzE8B/zrJc9sSLlrMAMSv4Z6yWeqA19WNo5O4I+COV5lYnEgsQ4qgt
ZapO8jcEeJnzqNWghBF181QK/B0Tt0l/Zt5rBcIiS6KKgPbekV5SJ3pRhVM/tpyC
yOzaM5EoZ+TNr9BCYEuITmy560NJpAeGW0n819y5t0dWarUzdiBje4vuFk8Rz9K7
q8gttJE9/rC/xNzotjcbk/ReIW801Em2mbwTg0YSjmW5+otqHSX//0q9qQnUpBZL
Jvz/D7hYxL/L5DFuWaKBXeE70Xma443yzjAwhDM2Y5U5o4pIx3VnYxb58Nga1rZg
P6xVyg1yqXO9djBV5Wdw3tT/u6tGeWUymS9V3y9bTBfCi8S3GiR3D0R0osxvN5Zg
LPeu8Bfoiz7P0iY/hApIv83gYIF4G1qyiCy2Z67Ob5P4HkzFAx1N4J6mPbYJUgF1
2GdfHro4a9SIMxdp1ZMAFc+5VRiJwGmrwAK9WPIEWat3NOw2pFGdFlpvp6PZ5y34
sweLnFzHqMZbzh8kzVOmhaUR8ABun/Vbc17RlRNzZRsIOyqg1qWOk3L1Kwn6ad+y
aLJZwKydbGgwJjTedo9rD6KVFnY1PkRGtnORe7pbANNnyvoW3MiYGBwk5sUAnZar
oRu3m1+MC7pR1Tb85rIoaF+jN1eUYY4K49I2+kAF12ieON191BTaZYgDMxiYNL2p
3mPm/ifSZgA2+vb9+mW9ZwiPSCvgMx2zP7ru+DFPK/iG+yJ1LLyJrNufxXmdl+LY
CxvfmNU38LzrW/qYqLwDLqFGF2ge9hTlmvFgqaSM83DjCJ7jrvjjsHtuuH7l/UKb
Vr7yLzLNkWzkk0ewgKeCf7g3ZDKr6yvPqYwsyZ2Tzijw/+0xVaF0qvbYLtwRBV9J
o78Gk3yf8yp3KLN41oOwNQ==
`protect END_PROTECTED
