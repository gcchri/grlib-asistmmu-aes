`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9n5SJ1ghRm4I8zjhYHR/sFb8z7m0eJiyq0HlIU9T0eYhizBfvh1j8omg6FumHbBZ
NQV45o95Zv9B6WSUG50Oj+QR/HKFpPyfWY7QFaHCjqJYVG2H+4SmgNqTynWg0cD/
D8m96juL8BEEeoMaJ1TuhOuBsgqhsj8YuE1yQK+vFgbcDKg8tZGKXuFe4meMkpeX
2SDMbbQoqhHdAKZDNp+KIs6NHh0kXGEr4/zmN/cqRH8QaetudVABkikHPYpMq+Tk
pwrA+Nbqy2SgtR2s3dEKEpKILyXZ/JrmIRGBipzmmxx/2N9XV4Wf53wwL7umJXut
rWFEUX0mBMiShwmN8wRf6xcFvuKZpsZasX/ltGP3dFw3Wo5l8oVeGRChzKglZ52g
6yyQ5awjI0R+21IN3y5BEZy6i4fu0mxHoJdK08RFbPjxbRTHShVribM4Tx4cdNFQ
Tvxin5VtqKwPA7IjCQqe6hKw4Yl2KM6JX6cjc5hJ04IZqQbyBI5MjlF/ENbkKRDZ
FVmuuNugoWEIjFE8DjqACACaPd4COlIvW14Qr9mHBl71X9qOyASewnz2E/pClHzm
1b7g0WayUDkd3W1zfB+P3VyNX/DwxEJ9fp9TEqtiJPxNpFpW9U0AdwpO+CBjHL4Q
05T0C2zGb9OSXhHKXaAyH4S/r+Q9mq41sN3cjD9KhfCI9eIdmgUr8HYka2RIXl3z
YhAGZhD6UA4qrMKxzVUOAkTG0VWiccn8w9ExqyMsJEYBMbbk8oQeZwkeLds8KYyS
XP1GLpup+gyJdWidbF3iopvBviPLzfqQ8f1esy4Zc5eE2LMoPwtoLJvGvQRf7XxO
x+Lw0ip5RlmkcJH5638kFp8AZON6BlSYoIs6uis3ZC0t8Y6No3RCj6gZ0g9/kAEP
RweOxUpBNGvTrNMsMReSvHfxq1Qhk1i3UlXibP0TiHseAgtHG87dQIlxG9Ujmz4N
qq/ZuZ1BnMrbrYl13MgDTc3Jquy8qxGiThIpW2l9NawO+nsiNlCDe/1c9PyGLfFy
GGbQqviVEDTVZdhNgMFlw3tJ266teXn8VTfp+SRGB8OlyxJXY0DGWhOJSamH2OAq
fq1CVDinxyTPtJ3ez6XrfRueyqDQrE41c4ZNM/8lhKQv4OfYRP3Ky7JUialnUDEW
Z1S8zuLD7XMEOU+8ca+kth5iSaI3BZiPRk7NzvuvKl9zNISTZPcciyFG6MbskmRq
tmt9uc5RondEMaK2wbptCORz5LrGnR7tRvyZEIdfju3Ek3whRUkBf1pMwBISBYw1
Q/cDFKm1EYrcum/+P3mzGNnqGTX8Fs3fYq4Ry4mtibI9Zy4eZTfB/R50y6loCxmr
YNl6HD1uJKVJWyUb7Mq/ZQmZ0WQ2C3rU9DoVip3UWZQnbqhhkk3Ksyn+1QbxFdFz
wWBmixax7eL8xHXr7RT2jYrmGmpzH6Q7hfvEW4yg7UksJgV5s2231NgPNK9nkvcW
TYtoW3KZv0pT9rLOvfWdR5jtrxtOxnzKsZKVnEywB3BXrP0olJAPk3FFg8tbjlnw
y2eobzJkn55XAFftwXa/0AJgNnvslS2j7UTt6wGycVshMKZNRBOZCIIjLQ7YPYPQ
zZokUY2AEzLqeiC1c/evIzdut/TFQXYDJmFMnK5+WAae8poGhwrvG/rT2NDsx+Um
BVMQ2+nmg+7rHWTR4vciUJvHPUa+kloZYVB7b2paVZgE/iUSHs7Mr5bEDdDpFAWN
fNv2JuVr9i6ngLI1EsF91Qen3kW/W0jenyzTYELHjleg2rmwL+zFtIZh8iMF7Plu
zWyFgQUAt9KXYLPa26qJMmC+PSFH8FZX6Us5FC/qfpiWaa0CD23u4KmLrJZZodb4
XEsE6LtlJS7fMhTTDrLZIqMONXKSfa5/kp5OJ3V6b8vfNY7wKs+Dusd+JC5ntoad
XcDbZ6RY8jeApgzCVuYt33kexBGMR/x8HV9i85C6wQ1fjtxpfEkpZDEZgVBr2sBT
/1o37RFoxG89PRiOzLAMrKDhUzlVhHwt/l2zhPMrLKrUCUGKdyxNOVHYU+teLYfB
JGDRz7VfJBvIYiQv+dHOwBzuws+/XlftzxB+Vz4zBXSg0bk3ntb9vkHkqNtE6dUn
Jv0euD1PWHKNGdDXKpT0ltMMTL9WXye/pKN0FL4VRVCY92ge4FCQlzDkZ0a9+vig
wTgeBpW89tTZLeLCsTylWLoAS5Ha9K/a6OwYbk+1spA=
`protect END_PROTECTED
