`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/3kQIVCcOg1k/jOjMHMBr/cnuccj0Mp2jyWDfFj1rtGp79tHGLeQUze0lOoTizo
WpMGLpVwXo+50e0HYkBROPZuSZNx1LriJ7QYLfQDjcwXk5VDbwGihyu5VtZCqh8F
5HT5XrgEOmN3ZFOfJ2JQICyacw/kCVZw2ont6T6usRTr/ORW6nwzNM2F9Yrx7bYC
L1jLiwUPyze8qp90wm5vrm4QtLn7Qx5+AC1pDqWmI+l/NFAyJYIktcNGxxPYHkq1
WtN0xL0EIdEgfiLhMqxVoxNa/L0tyrE/gNGyJsEkiQGPDhhGdmfE8+p+AedWcRj2
GWXU/LDUU7OnOepdSM7DamEPy0ORMkc8ahL+c3ArY5d3A1I5RpIPfdlwKmfeuyVu
zdL2GHHwSFVavbYs8ncMD+oxENR9//8W1hKXqRgaGtpESoGwhkZnlwzoal9PbnOf
`protect END_PROTECTED
