`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mGDsOjHQFAJsK01qxoQjFs9vv/gmQrU5dso43UX2fn7fUm0S5YgKQKi3MQ5qTsLS
RoQ875Aftat0dybF02xn/qpmzZ4+LkSRzJ/UVAkGtCksBFwqTU5vfDRDSfjSY7XT
b45iv/AMcIEsy8vA6Zx/WdZvUN/q18HKEfWxSOitJh7XwYzcftTqSKkR8Hcrw1Y8
wkpaY4oU0//zcvTbFoLDkUErHYDJXtTytIjV7WFnd7szTKmLo0GyirNYDbduTk3k
3iJYjQeSRWtS9nCq6j5F62TSoLQ0AKA74/ypiIFfeilH0hKhsW6x64MQ2Y79YZat
zMt5TynbJHzCM/d2AzWH+pG0SPmn2sTQFptW01JQi66ZBH0ah6Xw4xHz7952vDg9
`protect END_PROTECTED
