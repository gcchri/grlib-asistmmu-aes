`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0M0MxqtWC0s81vNeRHhTc8t4LrMn4XV7CGb0FlyObV5+i78J/lQBk4OXiTwQlcn+
kqWjkPjqDcOVJiRwgzXrdF09Z1Uy6qRXIqilADHMUEeSoFHY0XppIvpNbqwkkC0M
7Hmff7b4Kcn8RZARBx0v9wocgitKrbzilDiakCuAHtk8O3fDprSdflkQjMCKVs7C
TBYf7mEwVgJWLq8PgLVE8spCnVTz3TGcQtoFxk5zmMWjgWgAEtBeS34YrA4uKquD
OAvi2SFtFjd/fOniidW4RbnYUCM+b5Af9oxI9jqlAGNdrkYtrE2Q+iI9tGTAMRrw
`protect END_PROTECTED
