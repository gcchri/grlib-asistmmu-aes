`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PLgKif7a4YqlwD7nLBwrtnryjPSom++yqu46r2fL/ljqwoSta/PUhNPk/WTbtqsp
tqHsLnXVq17jeinMR4oX5STyPSjGQkp/UQSYyBgyJtNNBzuQoeHFrfmqNEM7l8rM
vWQ78dv562ZrpMiM4pvXjPJcKk8msK7k3BLOCaFQ1pWVBCeTEXmmSW/zZeTpEjwH
NWs0e06h1iqAeYyuan8CVpV6h9NbudQW/NGotxv5xIWWELuBV8bIGAZcOMcKSI30
C4FB1iXyhc4Qyai08gZjltykauv2xtYuEii7th3lYyxG4xOAu14YxWQ61XmAXefR
Ys8x/ZOrvy7aDl3cnSPFv1vLrzKJ5F06DMad/xTA/fra0yMmUuzbThRbh68uMYvQ
AcDnOKKlcXIFvDMTTXAGSY1E/yqCoTSvJTgnaKXxmjA72wXnJbi15NA9hVdwjj++
mLggvsXXouAOVMZYPx5VCqvFGOm9yaZech8LVDW6lwGtvXpLr1M2/gY3pvCIk8M6
LqNIkxEfk3fPhDjPzzptNNM/tiAMzOpzigyLBjcHTKE=
`protect END_PROTECTED
