`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3OGmfrepiS7pEvRJMOYeIu26jkTm5tbbReL2jpebMsl0vu9yaGTX3yh/1XO1beyU
KN6r6WMkFDLTpQkLYCr6O+eVHrGl/mvrHlNJiv3sDlfNd74mUGyKgPaGLtdzsZ7f
dfaciSxrYt8l4m+FgITybuExD4MENGg6ofVjKCmYo4EofZRjSSP5n2O5qVcGUIeH
z7lCjy80cTT9ebw7TIu0LMm27rep74SPoHrsgjtQGNBdhH0kEprEaD4ycU+9LPAl
+PEyxSQycCmtzg2iPs620jBh/1VV8leCSR89G8u9P1K34MNjROuZZ8D+VMmHg9kY
HQrh8Mhoo9SvVQgO6WKfvw==
`protect END_PROTECTED
