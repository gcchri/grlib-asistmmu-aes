`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZrqL3FfB1Rc0D1n3MZ0JsawOGIf/LDzvaoEr4WtZkli3nh2SOKE5cHCz079MLdR
q0sKZ+19YFFdrijnswBQnZ7xArCJAo8QuBWkwNIhPq28bohEStEpNRRrNtYPs+Yf
MtnWY6/yb1Tslb6jVXxSlqoB4J9sFFXgFo0cUqgNkFIIMio0gwjGR88qJexlBmxT
eO4eAuo8S8L4BmUJeXBxz2d4u7rS0pgyd2BNsTBoCJRMhRTAV9VywQFlhQzTgJP2
eIJ9J7T65h5aY5QX/pEZUZvZWWgtdc0zwe2ti6/Aqc4GMG4Reh7OipjIcNpa0Jv2
aLU0QFf1zOLDiSspuJt5gE06TCGa/SpgykkZK4AjXk+AlVrSQjvR/JscsoLDO4rf
3vCRRqVN1FR4dbu+UdX7DxR4iOOoov7Q6nytfG2A8WA=
`protect END_PROTECTED
