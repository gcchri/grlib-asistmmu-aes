`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1I1cBgOn5sqio0RdcTjvYjIkekwQ45W5RAetBh2/qU9M2OQYZONtyRIHtkEniLL
6tltqsaYanl/UnmiiYDUUbJVFMizxHtmVLwSfD7IEJ9j6D8oGdp0mcLj5manLtEP
owiUiTFUJL9Fyw7hijGCFsWbw2OA0WnfwhsiKwuj2GC6y+7WPpEELlTE5QtdHPto
uMeXw4TPUpBuwKoCmMxRd3/R05YxGl932t4T/1ccBI03NiOMTx9x91EJDt+U+Wub
iW4n88EnjMqQZfB2BObj3R/Xyl+L6QS/LDdPK3CAdmQoEX7nVcllr9i5u19kITKm
AjRGbx+suoCwsyy19mrdXdQHPBCU0PPSumvzil0oN2IzJfgla6ph1tFy/qIYg5Hv
Dj9e0y7CS+9LmMAk21sUyPAZpZpku0SU3nyyTskd861L+E8Udl3N4ZD9cj3VhFlv
A9EVlmYNQpLxYKoO/FBhFfWW548cb6h3pBPnI1giqRg6Ocu1FgciVj3JBOJCJ7OQ
ZDHNVISYA81wH5p05JceKaoW7f7pUOFpx3zlQR6fIqwk12Q4jLe3fAXmuusTb/Vv
7zUyPCV5y/jEdwkcJRpDRcbYF052FyOMU/yCKUw4hI1XldTVRPZVFD2yoMDNZuSB
Pf+2q6Srg0eVLGD14QTeJg==
`protect END_PROTECTED
