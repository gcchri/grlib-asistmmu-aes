`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bRUtgNxp8XthwFn8sd8n5So+7Eu1Jn/JFMevD/T2EvWGxpzIFaE7NPYw8HBMnJNJ
92eJKWAiM4FibreQCWXiDoc51noFZbaseEm442vqb8aXZGLu55CITHP8si5pMHwP
mPSOPykFaw1nWx81Ihj3yuIFkNPMn5z9PGkKTsnQHvBZSlvDWK6sBygsx1aiCXZ3
M0X0kUVrH7CI1xhrZ+Y4RntaE5yR0e+HNH+eG+82yEIcoLYNVgs8RrKLNlz7NPa6
dZOR32hRRLZpIcFqrJ+jOJkcXD357ya0BJXoJCbkSC8iCY2W7yJ61uTqUdQ5B4Ii
9hCc9YdNgfc6Fms1hSlqbYeBEwv10fVEniuGbEznYwgOph6F8OLaz+LKhF/Q+vhR
SlSknnEbPI+9BPTDwIXNCVuR6fdX956iD7BChq+RP5BhyR4WYI3/o+/GpxXc4+6f
Q1wfOcFko6DE7G3oPKeE6+IpekeRmoo6FJp8C7pjo1E=
`protect END_PROTECTED
