`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2juNpwI75wMsJuBeTupFk8ejOj7Xh68HjtX6YFsRSnBfTiMHcQb4mLqGNqztH9Qp
naQW6OZH1g/6oim/Tw4u2F67pLllgmYaj10E/2lJtHBRIBaAurapqaawp3dn7mud
ZbJxYsxmnLM5N+SzURylkFP8xmZkjezLQZNRodi4wm+fs7ViKeKTW2Di/r0WlP7T
B2TC2uFUmc3uuU7Bxq30Us9Q7pZXlWmXw5Z0BnUFp9HRNQurNm1r2Fub7143vDLL
/L6nEFvyCP/iB1me2t+la5bR+r3vQra8dIxp0Mnx8RLrfhrxi6ecaBZKYaAg1qk6
X3mF8lJgDCE95+GqN2hMxR2zOdrUxANFF62oVIcvdF87mUXlRRbpoUtCULiLA5Ka
olQmUGWhnbtbyfiStQM61gK75h71p2vL8gLZ3LhDGgTwOs7I/JsLa66747Pw8oQY
fZVUkDi2FRDFUCeUqNBwha8lxRHlHbPmiEOcxVABH9KsD3XXprybSXCYsl/RLpa1
D0tbcb2Zr09rgtcsnIfhMaoxHujbdw/AW7Xf8nTrt02cf1WUXUaGoa0iNJ1LQZRB
+Ly69V7zjglxN/NJbg6owOMOCZOXUjys4OCw52+vmG4fYgFqhlbAvDp/XRuaL7Aw
nOAnzXhoVkw6alQwswqrZzwPfZc15lXIdX6bOe+TAFaXuSUUXBdFMXN3TGzTQ/yy
gFuJIoS/XXzYVWjA1EHmogf/J5h/58g+iXGAcxBwvXuM1YWdrixFxA4FK65UwYpq
RILjOugeu6KUzuib6SNhRjFt7WSePQtXoLlW1mMLz3B1KwoOOxdSD7K8mfZTP0ZR
ysUUE6qcazyNEBbeEmYdnR1JNeyjsI8XhyEGKrezctVLsY2yVqNcbCPYC2EEdKIT
Npc7SRIoLDzFzc/pZtaA3yrXGpRDzM6osMr3trsVrF2NtGuQ0FslrzowtooaNscN
TDEoOYEJUSAlA5Y2CeaRfLjDqkyAyGbxQZlBtM1CmjN6xH7ut/nO64dvx7MvH3if
LtgI+eAQxMFoi3vYOUrQYuxRyfOCI5r8aeRoWttDtmcO+osVcTPKIt99q/cGfHnN
ss1wIY+0pMaR4VmHL6eJYwix0CPfbr3T1qKTG6fXnT1ps9MZqC9CP/qD6bBGj3oM
7EmnUBDLugKko5uxkbZemF6uiJISvvHABvUwu8ZJyE037GmQLSXPHR7ftwdP4QhG
UbienZvxdwlNnHWBI0UF1iHnwhz08p00PWrEbjb/1gv+Juv3/1Rrx8Lhxf3HcYj8
6G0CNtzqvEk+fXUTS437SEK2ESvdU2bTUwmz/dB4Mcc8wqCGs82cjhWzE5u7Knl2
k7Yt49aMLDx1D0uQ5DBS3IMDtLu+lGDXqZHHjU9EpSTU9FKKK6+Zr+uaIxF1oK9T
0onkxLpbtJReZbP9s8ILtPcTubZrpL9nBMrVeN1iHY6iYDoBDPYTmy/zCx0J1n40
Y/QZ/BrziIIude3XoMLfvl7inH9M0zi/Aqeg6hAsWMnLmS5cEX39R/KfTWZTtHzJ
sQzcu6uxk8wI9rQPlsDd5eSoUvlGiD+Gh6YosoxX1hBMfEUUBr6xzHlGwFFEbKsI
weybDgN440F3Q6XNBpfb6NKeFVAfVZhF6KL4FyYp2XZeA4aNpaQFEU/dTJ3D5CVq
cADVI0auPFxDSaJkHuswRDVfQi5bHMqMiXG2ph+m4Ok058W/Emj36O5ASu733vYJ
vOoqGyfxQOW3prnxFRmZnXkIqWu8oTeJrRukFFLKBSWdcEwQdORVikW1MqJbsGaa
yW4YbRh/JcLUhyZVkKuulWbDv1e6dyE6lpNV67moYh8Qrqw1hK20NeBRdqsQwT65
r6n1YPIj/b4mVaaqBO64uZ7ucP7ZhldPt7LBABkHYGo=
`protect END_PROTECTED
