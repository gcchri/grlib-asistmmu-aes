`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HBivPzTawbXTqqxcqRae7O+iORnCnqWO4P440u1oMnbXT70b3G8x8KZoZg0XLXHo
YK7klZaIa6y36AyI+aicn+RYvdl/h22KHXexkRMAicB4GsqIuRRYDGUVXiiYm++i
oEBRBrGMFfB0fzfk+/5hVcbiklyYIyygHqsPv9WswC5Cxv0/7H8Mi0FaLsRnr5Qj
dT9UHpJ65bQdEUHTLSvoc5SeoWjPLz8AB1yOJzvky4y0a4MgrMUvqFAWZPqAW0QY
BNlXWjibSSUqKWfJXvwigd9vFwtr3WnlgkPx4dUtqL1wMH+cT+q+aaWR+AF31cqL
D7Ghs4zHWbe3ZtQICMWFNNHtm0BuSb0EWCnZEmLPXR8XJ7vrW5lopkNUrH4DTEgP
BbAGKU0aatFRyaP5dCTPFax7+zWhm3oqcDJxkRJ/bCIkODCXr5gtL+OPVlrnHT7x
DXIgyX0j55/yNcZxA9V6f0/R6WXInCCai8h0XTULp9XFYQOdiCJhI+AU5Kl1r81E
xSlU9KO4qwmyW1oATXuLK1XhrePk3NLXCL4ey0ROBbgAybhu4pEz/+AGB/eaFUoD
6ta8UyBBEW4hz4dcyBxTZyzGTDzo8uaLBdcwU+n4SRZOwaxoBU8VLd5ExFptnq2Y
FbuC+0yifW7LKYqhfVNZuhOGfHIwWDm/OSJYLxMUkIepX1kBdQHOnpPxRq/VE77/
Ce4FniJKtmrAo0kxTqrc+n2vy+HHyn0ivGv5N1vvgJufwefU5hnGVLkdwkWmPIE4
7X96ySQNT4q6Hylty+LKT8+0t4Zrd4YY28c+KkbnZxPCzw4EneLuW3bzdPY8fYKp
hwr0NMUFlx6WfdOhywdqLiWa0yAa/YV4m5psOKg87Ru4jRqWRkLczsR7WlSsq1y4
XP6xdwPBhR7bbe8x4jY/81iOXC/QYQSqWfmegLkYFT8E+ZFnT9hImkmntVMgYZae
gdkw7+NlDtxReW2gf7RsAcE1O7u5UkzyD8lkf7B9QLrFb76zgplSm7x03Dlfj5vs
B1owyEBn0r478iFP35i8f9M0EFMUKupltFosKblzUvMLdmvajwlQ/fqs9ZXhWRaA
lKdyhWAaZZc7nQwMu+3mPsGqqC1qyNOGRp3iYNMNCAho5xAc0yQfOpmDyRsEa8zw
cn/gj91JznHilChFgM0uajSg+C/eCs8e2bwEYOUMLa3LB0q97oW9LzDvJuTnXWM/
4GJrmJyGt14yOF8CIQrlACSW+4LTHBbmd/hWHB7UUs7GdLMOwOJBm0nw6l1tP40E
fZvCnODUYaPneFbaj0waX7DERlqEyYFZINm93CxCMOUPEwugDqtNlhuiJjuen1Uc
d2PWk4QlwjrWHID3DIDq5pKNFvV3W+kDWFVF5gs7Q6PRe6JGMKdI0vLWos40aGv9
1z6Eh7eFupVof2FHjcRLOAcBvtC+abGcVQg1tCSk6YHhKyynru7697epR0lp0YqX
eqxGX3Kqj/EJ43teDwleXzXOeZhvmBekk65HFgqBiJYkVHgnrshLaJ3/KN9EXRCD
P6FfI8zOYuMj15ZAjF+ijx6fFTIaKauz41iZMp7HZb/YY56m97ZA/OYfqb8jZQ8H
kxc5scdKKyWByIkFREP/J/9G1rYLrDFlOFplKUkaLotCAHSqv9jMgx3T0zV8rlHZ
RyR9wUXZcMtHlQ+1IevtqV2MTx2n2JK7EtxM9VeEMJifblqz2OmqdqjIxlnizEvG
UN0QvJYriyiXhSnBdnwRUnE4qGyVCJWu49RUYKoELMgT6FVofj/4okM2HQAekPMB
L3ixdT9GGt7LkoY6bJuAZih97THnk7apWbluTTHwg8RV13qGKaaO/2AMFmNMrtMh
3AEiBd43ox+1RHcbnEwQaiOTxp23WJzYBCCvVVYZB6wqK434qz3uQxyvsDO6c5na
/36EFEx1IxlsbzTCiJYhooUoxiuGZRx1jFFEW/huWMEzH/ygaZNFKnrVrcQn32bB
ZcRGgdX61IpwqFyjFhYoXfk9JeJEdYZ3gq540r5vCGFRpyKYpfMYo8S/n4l+Vesr
0+C2tuopc+u12Cp7DtSHCv+vVKf84YYlz+leU6dBYLP7bVh/gixnObFqn5XFSxDY
HT+8CZqD/isoGvh1nTRlRIKKRteCJjhpZnx+MAibrTDu3DT29oefr/tguNhOs0mu
2uUh2IOMOnvem+vr12ItcA+jGIKk01e+hSQ0MKBo8biAHh8v6BDbDS4cW+WecD2/
eq1yQDEoRq+VIG9qXLwCZ4JIFfiY3h23sEtkeTjNBz2qg/AET8EyGVq4s3Qj5NXy
3emfvycHXRryG9qbMQv/7Rp2laMGBLq+OzhsQVqGF3XNOpzB9hefdeb84z5RDNpu
xXkZX3XjSm0d0EL7eQ62fO9FGHsKjfYb2sF6TcY5SronfbRStb8g7nfCs8ZVSqVk
DZHSn8grd/pABOTKx0My7xpylE4hK7gm1mWtDlOiSRoPDkGn8ZHVF6UvpSW5Ik0r
3tbs2MWbrKqs6A95EM7fRcap3xgPj9d5Vw+W93UWAZJ6YP8pBC7iW1u8g7dozjxJ
Pp1UVyUF6DnpsEMLifo/ww0g+kGDtb/asdxIVOTiybSLDAsab2P02HcQqBXFR2R0
rEEkvv3HMCgB2rkZ4FOC7nyrh3lDrXdE+ghjggB6nA507QNjKUNwMl5JJxNFh7tO
j6OSVmvs6waYpjCzbLsvtRn97zdo2Rw8WqVqSRGwKLQg5oepcd8ttwHYwEPEZ+AQ
YsYbuoPyDnSvW6WHsNiA7DnQyhSpxc6XmLIb1EXFmoQjzA7YV7926YNE+xn9LrY/
Y5Y1f39He4z2/R+ygM6z/OlssRg4iHVpS7RBxC+Jkfju59pZRbqtkMvCA7itj79a
jqJPG72+U4yINHJnWphVVLQsezrJLcDSBDpzbNMuuIGOy8Y0TSmwI2hF4sSFz26R
ZUtTgnBwboJkGi6WftvHhQE06g35lQI1bYHyyxIM3UWTNnR9mPkLkNCqTehM9UGm
czXt3xVwLyoKCNl5PHckOm9EIw12HcGgtQZ7/q4GX8WGVnNhEK8913V3uQB3A/QS
eoRc+VXVNxYWk2jCJJML+LlIS/w6LGgpqaqL5ykeFW8cq0VbFMpxTGB7VAgLeWjA
mAhiH/LLboWZQiRHzIDp7nUxY2zHDwIOhYthkzFPxOA2klcEAe6WMOPqgpS/h7To
/PEc6LGWkXxlXhwkXhS7EA97rruv5Lpcb2wpxaQq72ufngz8COE7rgplXFV871Go
VMqHRdRdp6kvr2tghrA1Qm4zTL9UhBgM8DMNi2szZ0vmjUZ9At0SGnNFiKdePzXB
gAimmyNpU4GbKKFZpM5jii2kTUcgJBmhd0QRrsy8IChdmK7WE4LHsm22jxOJldiz
JZK+0bpKZO85uqc56AEwrlLWVcs2kUAQP4R3ko+WlgVjn0xVYgupV2eLIq52jSAk
jK2GAYFny4rA/DenlWzGfdlygcdFWPs20SthlUuYND5yBAbFjo2Fq7rg2Cw5tgTZ
RefHTnmXmVcMdC8ZVy6IVCpAwVV/O/e7YLKnTw3q7nyeGljnEdw75k25LcQCmtYr
CgyGxrYVPwDc672aGxZqZU2SvqdBaFW9jrAppWHVLgYiTEuXYesHX3zjca/9WlwA
lszBo/XaXHJTUNmYxjbajci6emwGPV2J9tTbsPm8cfFmauVqvIrjl1EoxNwL7AQE
/NwRemwHumsXzTDI41z9bRQqHHSu8LQpcLl1put2D5XxPktPtHjPQAhJ9lK2odXR
kWyIqe6nVdrv4j3N6rY/9ALBEMd4vrpGE1WElRB3r639ZePNU25ijGOiAdEtsx3e
l/8DSLu02j/8h9Q7PT/4nEN7/vF1eRXpRcSG8aLNvZ7cmBWtAK/JADysBF0kKcv3
DI9XOTc/egSamGIsV05RdUVz1jCN0hi6vQDdkMZ/oh6z1wY3FYoekVJ83uDgIraf
spoHqegMNTT3+UMKp2g0FLRmoWrMG3Rt2Mwt3uIfiPd6fmZsStmeK6uHPsnNZzTI
NY6aIEm1loqSJFk9mceD3Okoi4BZCVNkBAfsooeb4GE8VlavR6/XgdUncdeA3lYm
rsx9n52BZBgCS+9E/iMhtXuJDdhFoB7/7ISd9ycr2NDeePNgzi/0LmJvvcVex1ms
W10uf4epVzOk678mjlJUVC+lqhw0VneRlsFAPD+scte9u3jbNRGZjNIieysGjVo/
xRrIQbtCsW52aPADZ81aaxVsNiauOpNh5CckcF4P7mJ2bAyBfa4X3MgNr45QY+ex
7Q2ruWjvJzN2XE7VOWvY9o198lKVDO2k49Bemvrn9dBcLvDaAPQ3W2R5CxR1lt9X
ucdJgMDiJerDd22ku2Hs/y4anmk1rNz1hH5n981Nnj9wkSpsuQAy+ui7arp8BvUV
lLQGKy006hu52GCHI0pG++N/d3vcyIffcxRT+PLJ7KsH/rjDJ0gochlpMZoaJMdr
UlfOeYXlBYfCRSDBK91AkjqcfkEs9GwCNrqSr0Sz0uirNmymb872zgIIj5S3MbQy
pxN2FXT0Zzz18LYDEay3/RqmERTtHrmVMU6hS2oh1LqsjlDvLw4RftRgpUGO2g65
PXExTzgTWbPKpAPFpcfY5p3kI5nwVUFPdFpPC/SXlJ88JHLi13u/e4LFXA93kZql
j3sQwiZf1A4SbDOYwZQHzIdXu6Mz1nAlE8LI2fDA79jrF0Q+rGU3noOkL95tl0eo
pqZYNVo89qRAoy3qh3tVfeMNEFUJEvMnFN1BaN1JKgNkEVzQQQO1mLT4PaMjPhBt
lAq8w9AjmB1igDuMK9GkPj4DYwZAd8UpWrngjFimZFkoVrEJw8SxGQ0PytU9JKY/
afe5tMxJRMRd7/s5SFCeOc7aaVxxLv1XnhTdLZO6nLU2nA/M10m54SK18wuUwDD1
Ja6XqYhwOka7iqrT8sMk3YpogUToJGBZsk8wb03Z1ifQqB19wMhfxkLb5Xct5i67
y7EZtBKNV6Cq7IlgHXEgery0YPkByF4tVvRNNcFpGf/+RqgA0DXlcFBRJq3h0t2K
a0UC9GrV9QxHrRyWNPFAHtKY/t6M92K461gUBIvG8saPJ8I1r2+n2xm8D3u2ZMbf
7ZvBXcXCqd4NKkDRD5fKasxIgOxAwT+VMVKHQ68Py/NEGV3SbnyvMTps/tLP+V10
1UYiXT9igVkhL/WcxK2xbQmfx2oOBdrN4Q3ZXziYZk6e+o0fLcDeLda9X4WC8zm6
H2usVAhNENCUrBvwj2/lw89QIclRqR4ZbXyeze+rZsySQisYIq8xQunnzl7wFeJs
1yJmLJUqQmnWthoupa2j1WjkNXcY38PrktJWX11+FZOy0iFRl9a3zNzVhK+bzDjK
DeweL+aBAFDtGj08Ko5cDaebIvBCvooqMxvNrQDJbpFVqmXuBzmLIs8fiyiiq3mi
8pSEd2JGwn18B/H+t+a+ImLVyNGmYbuAx7UdN5mtbfsaDBzd7YxiG6qI7TGEFfDk
dw0FkyTKhBJmME8z/6Exj0o+lGRc+Q7hBk39QDMqxTeTBupsUI6uqCUQyj3CR5lN
Tjt4pjXYg47wXdq06/eWlCJz8yRhGyuoP5wQqaTGD/GGZe9/J04qDyZyOVO02ZD3
7/5K+crop5lU1V4Rv+APtehUc84baAgwVxoFNRrgitxztW26DGgMUba7qIbL7tK6
8m9ZJlXOLDiCYuzIT+z+Tb2I1uYprPyg6YROvp75gc2S4cK3fs3zEnTiWNnmKO35
4rafvQ+kY9La7aoIoABw2J+apDL+i4XgOdNrFQjWfT/9nd1YCy3Vu6v/IIp74A7P
2U/HAy8mhU90wZ0mmnQMPQK4N7T4mL2H9jmI8ZXL54PJkO9+VeazYhN9YOfiD9+y
SnRBwcDdpAtXJBVQsEwvcUpCxJgIsTOedRzBRChdc+56BCa1kwWFdtq4/kJfgULV
r+nuLeA1Sr2axxQdqAtfiW78iXKiZSB1fhslV7f5goxq/YzGCB+Tbd3p29qgh/hN
ekZ+8fD03YZPyz1sQnEFgbDn+nQLnt9EanyHnwrQTOFyu1n5V8qyTnwhwK31Icl+
UEzi+CovGDR/qWncDE7NE0BcZtCZ5YJ+ewm3tL/v9MSyOtXjJJx96jb361qr9kD5
LZ0u6JAbTfoLLHcc/7YzRSEoLp5NmPLf5P2omd3ESVhfoZ7QY920QFhjmGbeakZB
HWIuWtGV/JmxiJOGLt7iK1a04qH9oOA+Z91Z5toe+f7Ky2kcpETtLm2Rdi9kU+uY
ygiN470OeAUYO4LTSiuSJbUNv1DhZvbZnfMAiAsieN5iUh/qPmVuVtbKbxgY2IJW
WFKhs78mxjAF7cqQOtC2HKszUdLUWLvjhyorU9+qDP1UX6ggVd1ljqYs32a6gIPQ
Mj/t24eirwLNP4iyp7mooeqG7BkIOFJwt/t4JDhmfAKm+tRMXM4jv7HRLkErlCPA
/7UDD/Fjt/jI5ohUbyp0EbWwx8ouxV2fc7SF4+KyK4Q+ERdmBgmgIemebl3bFINQ
Ru7NGjUZ0oMsdtnFU+CiGfllgj7gvCsO6lorjx93vbztUM0ULYKLaMOiq4ji8nnI
rc4HD7fFT0mhRITDWApmMwC77tYZPQEGZVftAXds0DAgEdQJ4mPo5KfyOdZw1Vol
ldLHQ7KF3llx06yDx/vXUam7BWS4+GOMtq8X6F3S1Du7vZTSj29zrN+Av1hGLjP5
RLXp/9hUGR8lGecJdoXJaObzqPYU3exaZsLEj8pdkarA/C621v6HUvv/H7vvQKyb
ojn1rF7A6uaFnmhlpA+2HGkTxQ6z8kUoPxnnYQTFPly+7J47Y5M8pyKOMiMGYnRW
kQ9XJ9rsKHApE5h1oShNSTzbGzba3XkF0gnWTwKud1zaL4ZCg07oDsRIB1Jg7g18
UlSD/BMCaZBGEsiGqFC1u6KBMkAYDOm6ewmaWRfY8J6FSwxXUwbKx1t2w2WVrGru
4SP35J0nwSckCWbuwAUMUT0DahEPL0sRw4HIQ05lYAz/tEkTwEytJtgiKN60tG+q
X22up8xbuyWRM5dOgDMYPM8UCOmmZ6YVshIpaq/GBNLxc3oZSIvqFtKqhRRrbQCl
FVqlbWQfwcx5m14sr+6qB5aHLB4aRYmxRHClR/GL3uU6or3aQbv0tHEXgbIDXlZa
zqD81VTVdTPZGgncwESTwHjg4od+fhAg/bd7YF27eBAPBFpak2TzgFCjzDWbCAYT
LTZ/KWw9czEQ0khkE+MLZz2PX70abgw0yd4z8+6SDjbkAxTjDiZPi8lmKNrwmxiK
uW9w2Xr7/5jB2LBErA/6A65F0YBlaT1v9Qof6jL3g7PIuMz+HlHPMdE3gF8wCmmB
n2no15W+LHm/hFtuh11kcK8a0Q1e/uyoL66QzatVfqkFnSCIRo/ixWy1tLDIGXUZ
THY5QbsEb+bhis9rLgj+ND8NaEPwDzIB89onuStzR6pySKvXh9d2AfvTbrPiiUKw
xT80ue48K0RD8QzVEjkqV/3lefOc9D4sW5eSLOQ9NnFb04kR4r6nLOWMEPf5lYvH
YjRma+R2GUIYNt+bBrhq18Ozi0kOfCLY3x+iHegk2Xh6kDhwtf7hRi5dACiumNJ6
1ZqN7ERlNHd14SJ/mWwd9xxUNJrxz1dPAQnM0atfTXlJ6DotSLcnIUGreBYHFwUu
2eNys7mx2KWHIy4QGsZC+S21spUX8mV+dInKOqks/DVxys3FZGB5lISVmGH5P0H1
E+oikJ+oJWwIZaew/zsOG0qRMFgqzCli7cB/wk+OEAxBYy5a9A3lN2w+McRr8D9B
CNpjZBLzf/ue5JiZfYFtAzfwVpqIxMYwkYJDlLlhkVl9MfLuOtsWzfkFUyWjMMmP
3ThB6I217n2S7VtqJO4Oi1NYn/9oVHmHoThfuJdZY/0xjEDx5+EgmAR6QNtqqPLF
NqVYckEF/IZ4Fp7GVI/M2Fym+O040Qw5YqOvZWBAqaRrzHak0WGx7yERD9GvvVid
yKu6DZ0CxiHVr6AlF24HZaVROka8p2ArD9V/YtPhdL8qSXYEX3XDuRRmqqoxIVMy
6PyLQm7+nrwuLaEE+7ruY3VsulohXEzTTruOo64x2z9FZUtnBrkv/YiSp/SVFgx1
XGg8Wy69R4VglaaGqbQ51FID0O9AqNgTedkMkkmN/80DxtPvoJrOx5wwbGXzOAFn
qsuDLKKlWbGEsdNU83FTpVyBb6+Rc7nmRV3mCMt97W3m9KB07e2+5k+yLbjj0Pta
+fnEqARiMQYXfo7TLjfxTkAjFJsCD/hFiXYK8hMD7lguKhN+KzIlUsA93Ak2db+k
XCFjaphoOdrTqLlHX8JToZ82BnoZ70mHt5hA/Zfackyamya+HcZqVsK34G+kvqv3
cNhLO0O9br7V0YKpAzlwv4jeRVQIQz8aFvGZPWMDJaEmlGh81hT2jHL+idVRg52N
xA2nlhGTYYKu/ad/viag2OSBCjGPJE6UsSor5gbZIuii8xVBTCqbRbd7JLu09qTN
NRSRRtuhTj3H2uI3zGCTN/HfBR1sewFMKhOb7bW6wjMqvXkuqM2yWWURa7LFbk/X
HYODpKdrzwx/OESiqFZ4HWUcSaW3MKuMG7jI7CN1z7KDK6kTiUTFuBlS5h6oWx34
d355iB4tTfh8awOoRAtRCN2KxEl3BCh7W0Lt/uA7ny6cgYNLQAgp3Uf/7+mKgkjB
WYms7P/+27fI5HEDovj8OBQHrCjLBtL92fTiSV3cqOxSIqeBV3q39ss613zK5Riv
9sj8HV4MKWuXoimxaWdHqBNaOebkQxKOztG/DvHgSw5DLghTxyItFd4DWx+X2LbH
K2lJv/ixSbQFRElnrleNPPesfeOoDdTTmd6J3OqT0HzyE5dEp01+myXALschjVT6
MBJiVZ2kak+8gNsb/QU5XJ5EhJrp6LYEOnDe5R0lgnmeIgdTqygvrU1pLmCeeYHx
jQZwTe8ntmpyC7T/yBwNh3GrMLBnzGBiuf+k3RQqS4kXRdk+czqYWG1kfza0mK/m
DCg0fFFroosKyYwwOPXkpQupkyNwg5v2QPZhCnBNTb7Qko8NavFrZZTfkTndT3hQ
y9zrzxBVwxdZt4WhgeSbo24rURwGN+NsBNDVH3PbOk5A3P+k60MQxNr4BhRHaJD8
yUqY9Wpad49TP0gYFrtf33i7vcUlo5IEwBaE60ryMF4d+/VGkWzj1k6Ub+MmcP7N
XfEZCrePriNUD2g+hCq9+0MLKgFWasH03yycNpl/QMYDxwS7QI3e4W1p6XIMzZSp
4QpOMQ1deqUgC7YS6TC4QZHDD12q4tMaJ0ApxbmKUDrSOb390X/zokoUz4UrVGcv
3CkqGfbOWVvSr+TF7uSzAGc5SXkKQZE77KYrp9L7MDvf8HBmSfVJdUUyhoM6+OMA
MEdkhCK4MxFL4HLbtpzOmd/8v+hUkwCmnawwGbJZFA1wDSgumkmXRctoQnXa4W3e
5bzyQYfnsucu9dpJC2cA3jE/iOjV1hNy3H3jZ7Jvat/b5xRf+tERtZMR2pA9jJ9B
s3teAsKDF7JxpxtdtYLyXqGwhreuYPj8hMUhMQVDA1mz17POqNtMVHKAl7kt8rLg
12DdPA6EPDZtM1A0sl+5d/PjlCKH2Gez3kkMxPf4epeNVH+0k8eV9+wyelbLiNf+
af7fh54OWlU7Ogva9vBcKlkok4iy6Q3Z3dKQq/EMbZoEEqboEL6fARbE0YOak/3j
+y9sazs2KPvw1T5bKonsmL8QufuHyTynv3ek0HCinN0M0yv5FVgl7aZIi0Ii1BlI
lt7uvhVaqQeQJbUbfdpaVBf8G67keOPe5TfChOmW4+K4Mt592Ql3YlfUzRCnn7ZF
2yNtWjyzfRofxUIyQ0iM2iNzOpLxLb7dgi9nIIHBfEqL6PeDU+2/Rcen72vIuBMR
7T8PFGNVCR4wQ65XKJnWp76RrcwqkuhbfQM29HFbvBCFiEUHtTCEV2XEdQubNhP8
MV2KRRIQTv4P11HD1mq2mBRSMV5BfG8C2flTepB2YXZZIYadaGCoTRIsKmZyEGjx
8sA7Guve3xxwTN6yXzxa8BtY7QDHqN/UYnfw3rVHYN4gkg5uCH7OWJjmsezKIynQ
YzRg/C6eeus7u98+ppwhUFD/Djqj8PAxRpDqAB8eRmIP+Ht0p8pid05Z3k+aHy4F
ORAPXJnqIqIHXN/wTJ4sqSA6aRCar92E89xzTv7fa5NC95Z7Jr8Q1m1yAg3mIQvo
8pPlFPOVEwsY20nx92KQ3P2IPGldT6IyCyrZkLXP4QpVO/HbHHGxw8oALu/Y1ymn
J7hq5iHPUx/FAY6gXAbDPnbH/HbPYYwJNVpTQNDO373vUk71c9RqJuU7ZRM/VTWN
PQ/esrVEb0v57q35A098lGLJBdl3K1Q/lNbXmici735Y+KzIe51S/J8p0JBnTBJT
ejeg2P3XxfvFqsl+pdnBD4cEc6C32gpzbr8QynRw4b6T357LMKZPY/9GrMIottpK
VcpyiJN+Cm7W3qHqqyHYEguh82w7fLeyl8iHbw/h0/0Gaj93sCqBZb4emP01/h5u
VU2dYG+2UL6spg5Cmsw2JoBgowpPEPpoHSSMaQeMqIt91BiDTgHXyTAR4PAm6Cms
AzbN6nnDmoCABqC7lnfxTj09Y1vrfFRyAmzofqypddn8WLMNCNfjvsoY2yXlXPan
Jt8rXhh335D0X4rJKvj7AgdzKNrxZuULJcTLgLrk047u+6ZpxJQnss8hyn/qtz/E
HyQdV0TAE8y0GWFTHW6EZaffQRIkthc3+lLoYP+k4aDyzUXj7pgwiJ+xHdWSVtZg
oZFeJJiQ93VTDiul+JdswmYiKs1Izz2YmdfYTqLyMnU94GLOGNwmj4lpsqZcFqkN
qctysGm/8EoOaMDQRdGAS+U35E1gQaDS7n7ScHe7Tge7r3iN4q3dUplWuQaV2Toq
RDhUzsbIMU4uKTnw8zIyb/xh+L2E/dWJzclJ6Qi9LeeFUfg4DUt/Gkg7H2N3QfE4
yZgqM28qAM+tLk73djdknGJm5Y3kal4694rLSyj+m/tO4lWKHRwN5I727BXooYQq
rpkzXoeftPZ+71yvf0corobBm4VyXwvYSv5FhLiFQjCJGz/SxBjLK+pgCE51uyem
85grDc6rwssXC7ZcjdEYPUqKYgj2PYdPohnb09Xzxa8EIf+uXcrGL59YvfdPccnU
EFw1vX6D/e7MPgDIxfz69g6l0ZU7biQkq9P4tzw06OgUvKmjkag3XTREMhv5JVSM
c8qrbOBN9CQ60XY2hA9dafgmX6CBEtGa62dd/SUrSEJmfdwUx8rjxMQL5j/PcUm+
yJpI6Y4IqQ7FIr3W3gdWgZGgwmpNVN6ORQ1ake+8ulUJIGRRIdJvcakrHkNIfNgV
fP/jrRTxckkJKsqXpdUQwsbKnHpfSW9GFzwHishTnqB0ccYAIq3sKs8bvPBTnW+D
DjWiJxKyQKcBLxAxNhw65bv70rYVVsolRgy2kE3+jeNlQJW237R6Uk1xBPnN84fX
+YZuPqDDvQ5AizzQLWUgtEeykmRUQR6eVvD3dRFkPPzHEPlzXO/xyiM/FxEG08KB
LK0RCAcsJanAtXvLjVIAd74ewkQ88qtvsCCRIpRSgvcZ9784TN5ajBKBokU7IrOS
2EHzBvhHBAfRFaEAVQAjQmuUsgkZZNkoZ1Mt3E6a9UT9OAkvYDzRkQmGAwph+qv3
slv+/ScaIf53yQ7zXNmV/kkGCzPXxNBxBnmwBpCMdJdfPX+TqsRSN9SYnj3QX+VO
Y+7inymD+FDsxdZqKHB7Awq9gE7zrGe1SC+lFAZzQ9PPRcbOImgqFFM7Q6Xyp/ye
CGi7NjlqVXS1dPDZMDT6y1BBkIokVcVrYjFdA7HEwSUeOjHFMQnMCt7PMV+vu/wb
LTQK+zgYELOKDR5TzIU5AMs64WkeAUNrPvTocluoIC8zzoSMn0JypBSF801YUIt0
HjivjDT5dMcgkOoB0IrtAKTnI/9sSniZcVhA5kqRq3pRDZHDoQA1aIz9USJZcmCI
+FPg4IHvVEjGbKbzKJbZd6ac7pjqStOllPRoNldiqmCVr381B25nLCuEhBg86ZaD
C11EuAR/JbUEWt/LuQAgggfkWW2ArueGQG+JCntDTFlA+qKbOpxthdvC1lDeZmdA
WA+ScgZRTLdbpu0sY0geZ7SaGp7cAmAirA3kB9iDyxw/Euln1WbVJbvGSK8nlTKq
9To8Wm5VgbO7V6vtsQ1PpRiVABq/vc8kK73QJVjXr8FDxZVnJP5PvZQLE7VmErFD
uTsv/pBlfrKRoOBPYwIDAN5EBhz+uS419IlxF6m083M044QWI1PD46tTewzEAAJB
xFxSn4maf74QiervDsxvc58cQRoEd06Mk0FqYPkL6vuc1b3MVysgepce7zPTwRvP
9MitoZzyYVvWpb1dj3tBiVTa8OrG1VDenALbUFQ2/kqnHsYy/KkV/PtEPHf8SS7K
nZcGoyIg2KUbPcDPEbEOV39Ga8Ehr8qtNYxbi68j9FePTZG7XdSaT4sG0FZDxveQ
o1VGlbCJWs6R6aA8qAsmCol5JIuQZIe4/z0bAVcL8s7rdmWAu70D417Js06pD0Kb
nVpBuzBn4o+P6A2QATkrGsVcpAO2GvyuI0ZJ4y6036SVWyZ2s75t7BxAl1cv/hek
eJjlwihvnMyGuRi752eTCxBPyuuix6BCD7jsh5cf9XJ5ODn+Me/p2uDK8rAAc5Au
3BRWhHJoFvCseNS611bMZ075NxsLkoGcYkYMB8mzQbcU5p3qREziGORmSvwXokQG
w6NgPvzSa9/X/xhX/Mzy27NzGDwJvnEX8DVIzrCh//4HhUCNXJfzSid5MYcq51xj
Poo7x1kgluh0ehFIrZqUiavF8rH0NyIgduAL7zhvX0dkMoWnh58HmEOKk1yqK7XC
nGXjIw8G3K7UXlPUcTG0bwsB2Mgl5VTxNZcIxnX6n5fHIBO5pH3F5XMIFBdnToKr
84F8I8H74ki/LZzz51KQp734g98Qz/uvyFkmj7H7sqFrKXCaEHzSNOigISA5slof
ouSnaRQLZ1Mg56qtLMaB16y2mGtb8ZwZlZa2yK7VQcmhVSKgvgsDsHI0Q75D6nfQ
cH3zyzkH5PHQnLa1bROUj987ZCniB/IfQKfRELEZBxvc3PNfpOSfU6/nWGhv8Sk8
Dj8wQiFGQD4tD1z2OMSnBuuhtyZuHrM8JUUAUfzTIRYPWVSwPEkj2qz06yCzuEiY
6BmiotZ+7Jt7OXCbhI2kempZ0h1v4KeyudTX9/iSwDlv9Vxso7FOpT2fb27Dt4nt
2Eyuys9EX/Jv032KWh1wExYM8d/iGHwi6wxGtwocnbm1eg2DZEPozgQ66YYw6GwW
NQShHuua7XNWsHcHHdoLc10qNYaqptXCRKZcjeP+u0t7KcEifWX9lkB5OOEUAF2Q
LBcEZONSmtc2S5D0qJphhEUb8RMAtCGw8uCdvQ3VynCQBxJVxCQQ3T5nVKPbBrtF
VE3m1fjv/wbMv9c1bO5zti8QFci9yj3uabXlN74XHWwMcFKbPWZ8qUEnNYZtB+Ye
BtHTuJGQ57RTJwK6Fap8kd7J87VhkdKbgkLrtuBeevaKmYPNO5uB9GseoEe65EQG
6ZisxfwR+9A0uueJ3mMgR4E0ezkN8JU6UL0xwd/y2JVcX4EJlSSfUPTkNNmk2bxx
Poc8xmQDSOWKh1Z+efhBn+rzMsLjFK3XISTz8zmDbi4BWSRu9Ca8RX/g/FMskr6l
8NRg/46MaIjkTLjHiBKnPNxagvXHijGvhj99WcsbRT+IW9emt8FSWkru5rl4qsHd
w1fLhKGe340tSH63OwFQ7liHK5Mi4FQ/EBTd2TNcyy48kRSR1jXvwM/p6feyuS2C
2YDnjCPiSp/6n/X2VM9QDWN6IjGo1V6t9fJhv1o18CI15Qzqq07fq/sEmxOUZldT
TYfpQdMWFnY5RuguwEfHiaKB10uU0bDOs9cmL9XeC6M5Q80/GM6ISVf32GfEfcVF
lXh/xa0O19mFb9X8tbKiQDXXNb+EGxJe2cnP9Mr8V4AyluirRV9nVBZpsI6NqAmi
cMbZml9j7hmKuSrsE9jpnZru414Y0r56EvcFHstCiEzu0lpKitaxxJ3w1PVX/6Ee
rQ4tDcKE8kQq/fGfDKBBzwLIKnxKgAVhx73BF44iTOhV6CbQIVVlgfAuXwOexQS4
JoHpQg9Vhzghal0stj8Z9l/bDvA3iYeLZS3ip79N3YcQ8CMnoy1Y3c7b/u03PKL7
WKCGJJZB4Yyer8n0AuJhprdp8skoKIjkDr6lLja895wxxn7MSlJkC/+GGTxC1EfS
+Xm2ehS1OGhbXnco9AyWqegdj+IlqpD4RjCpFwcOjoQtnYMhoITtQf9YZX3w3z5y
9x3Z8i7NtqIg781kblawE6UIee7OLCgGWVtMLJfSBIBN8XCsgpEhnA5K03suIoLm
PYwx81G44Hpn56mYISA4vVKGD7kik52aL/4JD81nWqZjeWXw+XjbwYi75Z+sCSXo
aUvFNT87lYu1FCtJFdLHsvrB/HjOmZ6bTFuJcBiftf+NcY6lpPc1JiWxzqwT+6lX
PETsH3OhEL1loqXJq9YzP9mouojqRp1f14hqJSVjzvweehLD1rV0ac1t61yxyIhC
7asB8asYUnIQ/sWOb/46HiMu01i3nZKxTtlPKQEW+7J5DIImN7d6RQtgTYPcOIde
8MKsLiOiE8r5WAYkJ1A7jAX92uZjXgWdivnRpvrQjv47yXAcLJ+9q9uYTEdx3xZr
QlTGDcpp6o6wEhhtAbEL++PvJGCQFZr+Olsh6Oi97LCAZ5c+VCwcco8hne3fRcMc
mlYiuyq0VTAm6+OBQhpjk75gx0ebJNLKDlbCRDXkEXx4rR8/CFez0RmAJNjQfUEh
FlwWzjFmZQEnSe1cJ2ENxC0nmn3MdrpAPDIs6kjy3RoPiRzaH1vVWH4kCEQjQHpn
Un2lJS6MG36m/1UaP0LsVlIHC/YgD9naSDoaAw/5e7aD7PJkefj6ZxTzNPxqScio
GLBnfNyGQgNxz2YOlt/3UOh6bXQ191vM3mS1Gs415e0bgpVhd2gH8kSw37WCgzcP
R/W9yj1SbyE57JYXfycA8H2icdQMXKMgSgV/xB4zdr31/cncZtimvZAIvB83JG/I
1abtoGRBOr/NQx1bwKiKdDHkm47ebnuyYji7QBJNQoZPYRgiSXuNa2KTWhgYpGDB
f1viCicXr5bFDJoD4RmjytotVK5uLVKpj8+zI0YIQBnmx8/9EgESMxiQTdfwaW+P
v9uQoPJ34/nUZgCBEjL8vcRTZmAibiZY7RDVjr3FAmcwpmK/UPhWn0r0bG6Bq0jn
hXYYLnSnBhjQC/e1YUkBqnkV+UzqgrGICo9GICbjyj1JWGxn+x/Xgmoiljb8rHbX
Kdpt7qcLNjn6s6/02QuhePN6K70xyyVXL+oymnvgxYnriuuyJUlG932c+YMqAjhm
QALft7k06b2uCgEPM5xmVVYRgCU3kzgcCOCRxf2SSkO2CcJ1ekzIdvC4S3Xy0j0a
3QE7BK+tVCAYYmmE+mTsEx5j9O1oGI9xmTCc13y9BHZkOfPbAp1DuZiy6KQx69Ob
fW/VAg5X86M6u8/AS94ClKB6og/kmWiksdc0+4Mts2r1aBEIm6nw6YzEksNlxFv5
xielQUI1+dJqw2s0OaRw/wRw01Pq83Owf9I+yP/29eMHykZh3m7830C7VQUSyLGr
v8p+l8ulUfAIdHOHAbn3Ld72G0ZyeonYH1xLBYRLEtX+4j3eWxpDfyavs2qN+TdR
0P5vkocj8hmFmfq3N1r39wVJF8KwB6XzIFUjhLzVB3jNjRxpOKKNfTigY4BFKYOg
pp1rOr8ChccUOPuGHLIQOXKjZ2FV/Y65m9c8MG8zilaTzvMRJJ4o30exfKaNCjVB
iKG0Hg/Uw70aeqIVUzC0FU4d9uOO2OSS5k1wa5yhFNjQKLqLsBmsxbTQvSfc+6uA
woZ+a9U3L5MS6gUlSs+ymaagkxcAmVBw3JCQN8WL52rbajvu8Ln+ZLyQYz04fc3b
QIgoG8kBZo/XM9mZo8FFT4G67jAdZY3YYG+5Fa73pB5vYKRb7mUGuXNmXAzVBvZ6
q/90Aqb/A33n1YkgNCtCWpNTVhedIQYZhEWo4TlymIGmvIfjxB7HpxDU4J3TMyMs
ErQ3UT4lDg6f29YGXHU7tOWQ9KdI6cTzQERKk7n8d5EitJKgiquXwsq1rEuC26Fe
ButRh6iK1F3rpP+HrL0fm9mHvLVVb63SR+raBf61M4hFqszKg9th8GyWxygS9nMT
OfP8ur146U0IcYLwICbCA2DVQ3fQIShThfvWi+9iiZsjmCb/Wx+Rk371TnK6cJpM
j82CoNrnYFki2R9yVqiQMkZ2fuLuUhooQ+EjLoyMrkmHEaHk3sW5hQUJ5OkFy5GW
8oB4wY2IYUIQpjaeMAHF+p28id0Rvmndo2UkFXngiMCG25VCMkx4g8WaZ0tt5rQ4
ZGWKnNms8NAFx7ltNIqcgApvawLeybW/lxm+Y2j9mupDMJ4dz2l+tadEFX88cZwT
iGX+4TDW4dOckk+pBJa8a3ks4mg0GJZK+5YezcnbdRQI7dLqcxw4+xbQDCyCsg/m
ATrEiNj5SiFO1f2NksrJa4H43wKwvz7yYAGSJBzepoy6OI5DQHmTQqSDxUZC9NBJ
V1fk0Ssu2cypRXXKVRQvLzdrFPYWOEml9as1fpW5KIHtY3KtIHBAXCAjMIAbni1Z
GbZ6kisKyzVWrmjkQZNoEJZdr7tSrazA8nwWqGNq0/0u2DzAxoZvTKlvA2iren85
xsXAnvM9HUznVaiW52Rgw2q6AHKhJuzFCqUVSC3f9FIJ0cHoyXNWSNin02J71DB4
FGP9nfGNabsr52lrY9hRR/8QQ+PJ+yCSeWkcPOuISXRuHijN2Dj7PQAD0xGZlohU
KjyBsmfHzr4IDxsRInZn8kznkndv5txP4KC2sOS4GSc1o9t+WYPOOIho6mO+cIdh
sNy0ztUzQYI7qpIJlEraxYOLWKfIcV20zB/wYmFXdrP5Wa0RPRkgPxxcdISGpYx2
cRGlr21BYz8XDUtZNi0Je+LvNrWBUM2FePjExHdzb4bH3KNYCdsFz//CeYIy7J1M
4hnTkQESv2lC88H1L/mpLWYxOSW37JZTtWYd/OXgFiTxQJew6A1JeDCuPXvEhlFc
VLxEdyWKfzLBllvtV7H/5aZd8kzjF7EGAw+IZhBWt79ysfkJ1SlvCq8n5bJmR9V7
P0YVJJVbsCLllN/Oh9KUftjJWy640Sdgsf8dienHgeH8xtqRtg6INqTQFMwYmMxI
Gb6oTZQ3kljq2/sONFyq+LreSl6W7grvBMQYMchxQu0J3K0rP4oKflU3Ob5L1ajF
6jPzBnFSNX/e7poebFSPMq6++hBJTOaSdSEqt2kwAcSsbqJKi9GcNZ97HHLvjqUM
NNANjXBuGGcOpqPg29wETY9uvDHoFhaVbNFyEwsc8IjBw6Tu7O0lgSZK8JFWfhQh
q7jT9X0THFyV88iMTZa4jdM76vM89abV85hmcbVcWLJ1QH43eQL+WV8Ymf4v0VVo
eCEBvxzWs5RK8+9tVDsJTHNcCV7hZVSENyuk/h6bu9GA+mnsM6ahJKXfLlhF3qcU
OmWFCr15db/J9luRpF6NTUiGJmos5Dp+tW+Pcbi162i4IAeLtlsp3oX9nTn5PeGW
roQfGKgTsWou4Lc2NAoc2yGwTzXcAOvtxB+3SJWBCjf8d2k4D+h1FKHAIKll/27r
ZKweC4HOY+6q3vEzb7bZCKEvakLZqXsccIyvCWXe56OPXoVmbLKGi9Sr0Gq2pyf/
Q8+quvPgDe1QOmLshCMC0Dc3poMVNUCYjAfvDZkDX8CcjfQfE1FnOvYsnWrTgPYO
AK0gDxY63O58Q/+Vkcx8QXjqKEcChwcPdvtO66flPTG8Y9ttdy/ZlaF0mA0GlFF2
fcvSxRw6F/yXiyDUAT+gkWYmhwKyJYdNf58+KDhlxnp+kHkhCxp6KHtY1zYHicYn
jHQXCCSodUlnoiB7UvpIsB4UrAdXcNpzLEhAvk8yl2pip0VEP9t8Toopk5TT99XH
ZkJQH3CCYR8UxC5r6/H21OfWvdXhIVF32BgzTL08VFaEuMLO6soyOm4PkbjKUVi0
p+hSssZ93Hfl/OJ5zH7EVaQJx1ZII8xNxHwjWN6Bva7htUrTkaY4iBrmvwadZtDu
CZ0M5uYleCxZl+Ap+nXE2Lk9bQlpEIqvVU3aK1ODY3B/E7Mv4n9sHsByJweHDM6B
YjnARXAKjSVWOgymHh+3UPzGOSoCKeWEEueA1Hz4Q0DeYBLQzNSAbDwIHUmThSZ8
F5DvpYR1k6iEHz2wDPJhHP59fEfg5zMfVUKW8oyhTqo530fao+jDZKESB4/h5bAa
2DN5da23p6LoI8gvyPQAwCw04DeCW11KYf2X787bCFWPVr0cwdKXsPBbK5p6UhJp
1BLrlr9a4MoDcgClKBrJAMkGyl1LLtCM4td+EQqUitx3LecIo4tGN4PP9fuqUXQY
yGgdQqTNv5s3gWmewUPshZfifdrRPKzdoT528hZyNDPyDLSBm6zscon2hG7YP/K7
Uk5xNquV7uZUIjJZ+4jmHKk92DKTamFtgMhan9eLdNqOAGU0qY22CV7OtbZTP9jP
bkWuOFaDxX2rEtTbxDokQhosChDaPT92tOku4wWUVYtM6cNOzs0rR4MBBmvSOWHL
UlV4dRDCdOXbReFY/2EsLdq3sihIHjgSH9ECG+DlY2xhVJ/I0LAssDk6m+hgYY/x
GqUZsy6IiXCGzGvKPUAG9vW2mdBtg7b74e1g6D9fXtUH7X7b7DU4Bwm4Kikul9ln
BDHDLsMnVbmMX3TeAt1BXNBD6w1RLuw+nSNMOMrOqNGrF69nX9h3pD0z1453uVtf
go+1e7wjGLlSqvKNcloGjF3viisPfQwM0BX49fn/WuCSmvZ3dTQPnsqra+g1vqPr
6386wYv2i8TtoZxG0ADRGZbl0M4RoWPUVT79z/1rKKDyjTSOoc28v+dvcwynjCtU
LMa6lOqVO7mUVOQnFog3EKi5xi66UaaaV5qU1v8szrBAGSjhpZtg3UXeq4y7ys2d
uq3xOrLTR37RJmQjQJNutc2R6Dn1Z3tcz3Dq4Us6CRNWIwZVup//416ETWm89T84
hRyt2B6oyvdv5UqDjH2Lop3vO4YA/KxM6zs7CogQrhCoQo6ML/Ufmz8H/lY5+qyB
YfH/3AJJhd2wK0sXkBA4Cb58Hl0Pr5ov280CNWcnFLtfA66w1rhcEL4JpnSFgN6D
LqCphzBFMH/m9IHXWWdillimP2nvCAOC1gUjs9KntyzrGNlDhwf6/KXSSnm09Gj+
Z8lacb1BppWu2aD3+l1l6p+VhmmOtA7SJgbvASjxvItLhHHBWYJkSKvhTPGqfj1w
ExKMC0KLZ3XAhvDzVtvT8ifh9D/rJqjZfPwCnQ+Dta0Wzu5NXSNDs6ScQ40CCkvS
BI490zqriEtXFBsM3fl88ckgtSTdwcLF33p3Q4tiLhdJNBpfsfqA/YA6hfqFDMc0
GaC0w0GLWTY4VGPxA/zxQG1j2xdRn2u8T0y7dfeG/65P4cfqXHPGQIQ6An2s3Jbx
OxUbF1d+7hopf2UmOp9b8dVQCJQ34+5euqfwjpzJEGAV799w162sgE0xs1eocUzE
ovOJtcPe7VFjd59sUAN0ZbG0SOQljvjk7ALlf+kERPUj7R58Fk7g0OyZUNZnq5T0
JoNDl0gDnZ16qUUTC/PrAGHOqRQkVwn9DJhne8K/eXi4Soc9/JihkIKdBksQr1DE
xzD0b5TmRUKsawSzUOuG1lRcynDsCVUrfFbR2Nw81yXu+GGPjm5O+H2MGFCTKvpR
k9Od10yKbo5JpvmUa+apw7RVEA2BcIT0uBOpBwa6dzg1l2l0Mue7vtDx0kuPGXZ7
Z4y5G91o5r+oTlcXePzfUs4ubPfHjiELbypwpRJmLXcO+PZ+i0tz4xWN/eJD1pc9
hC+J/ROhJwtmbb43wf7FukDqPaQQMLj5ElSi/saEjgiPT2s0TDx/Rx24ww9FxJ+H
ZMxO63inZFjhLiGXwT9dFDH4pT9JDTFhEgEApvYKduJy2lJKc8ym2FbIHcQFZZ3V
CzMwQzKWRrZaXMMm7VUQTP+YfCUrw/qaS33DMDT4aPTXzv5ST0VlfVm/tlexGi8K
V8XWNx7VhA7NguDajNDlfdUVhNZzMGiqaraPm7RF54RtzyNz0iBcCH1mEsYYUbDZ
3m+VBTjVmuLrOqiLdjZoJJdGLYc898at88vZsO2p3qajYOZBP+dxnTIMaX5asHFI
NGNKpy8JtY5qivcSfEKGbSD414T6xAAg8NEcK2Ps2W5aeWtjOBioAWFxaV1WqQ4s
ZdQsUGbJOfBvTGhH7qZKucKVZQP4Qpb1JwnRUDW3v6Nf6MPDX9HxYzRa2zWCD8mB
RGZMZZFCCUNYHpt6pbitdAqANvhA3DBCynlirFxVidz+QlR66tMKgwrzCz33n2Xy
sXm/JLM7O7Pc2j80ueKuva22n4vTOTfX4d6SL+KFm6g3EMwnDgOLeYaXBykasEKk
IjxMviXk6RmQBg4eNTUuQx1zMCe97QO98u756opIpuDnCxIZBhDq1nzvmaEr9vnQ
wwFi0C49/nIbcM/rKA9qzR6IAl9MtdovQPqxyEqVtVLP1v0M0mGJZI+YkiyiWUoB
G9AZOZAKbk+lyYWYxI9skgxkc5jtlpx30xvWA8mj+f4KnQuntLiO1wMdinNXi0RG
P2NF8oBJpXy/SwDEyfwCM/0VrDsJA7BD78trquarohqHkARcWwTJJ3fK5tI7kbfZ
J1TmS23USmGiho6KW52juXVAy9dzRnHGGrqKdz3KtqjFXUezBCpC3y6SUQ75TQdC
sX4JlM5v8bn2zAgyJR71uM4Jjz1R/h9/l9RgqXgCAcWwwM8OK93dQTgdMkbZQvaR
s7M4ENkDLfJ/RfTQbyx7e5gynZKxsA+vpwqRzmp097aNA5jn0B/VdY5HPBC5WBop
YyZRhmMzZprMPt1Dpuz3CP+kexmD1Py76B44LdMJL79NibS2agNltaNd4oXGrT0V
hrM43yPJdrO5WWSf4MPJExkgZWIsAVGhQfxXBiyIaSy2ptQMezmWlT8TvV1ZgsUQ
oQchbJHlJbqNe5BmdbsuN9lWxpZdVyQFH/6kYleTjNKcS6YDvKSoKtcUC2Taqt0n
uzZJAysduql6NboUaLHOVxQLy5FmblLnVMFExnNkhi2L5JcBZJeBtfu0g3Q8ZRDc
V2Ab2xrePDxNaXybC0xJFFykcNkcckDvLyGrGny9ol8EimUmgd0VSYSUkEYqtGWZ
UBODu4kZrJ3Pd9gayAW1OK6ILQxg6Yc7rlgyAv7FF2wfuO/7gQLzUNNIcHs2oniu
sAoKXM0RSPs6pM8ypgN1uyRQZJfaK0YXNyIV+iTlXXa4GwCemkNSUT4gYeRWPnwm
6OHKlHuDaGXZtV7UGe0Vgo5szOepCXeQ3Q1h4ikd+ub53/oLpADVdBeD2kBfSMrl
v8MF30dyg4SX4t8UdeQwJMDtEy/Iu7V8OC82cXvT/w1++XPqRW6Y8nT1zL6pUeJG
qfypQjCVumpeuNM/i31bQ1tZnucsIOjQiUeb7Maqp5Dl1HMJnWIxsBroseJDE0l6
mhhQ47fx4uECHkIBQJM7nuWZWFjlG+d8mu7eh5p+uQFgERuQi4HmgGoZgL/tFWEi
xT2bGdx+P7OXcfi9YNoIwNUCrnpodJ0iOC5jRrsbYCjIH3TYd62zSXUH/bwpo/kU
qMjaS8b1EVuRqtSlru2vUOSs4pzwbdRfDWTuFl+ynoOno6G3uQarClWCXO62ilnL
37BpLBIjGvt+4R5E/9yVSXG4QOJGxWGgja37asxX+YgDPaxHfLnhCDLPQ1T3mXtr
ngm0y9BMwxa780oyBhj0Gko5IrZuJ+4ud2AnEQKvgGp5/ifKulc40bE8yXItd5yw
wAuvMUbUuX8KTx1d8c8TdsjeUwdNq1G6kbtGGBCF3gXhhVq86nuRIzbFyCs8qNMX
macRECRR8d1W1Rq94R24vrcVRUSPmY4VEDar3V7vZVThb7gJfLWlyZXztaTf5xRb
isTT2jmcJlP7HlpvG0OgV6mA43TC01TGBjWbr8Y3b2khXTyQZBFmQ5euOI7CajDh
ry750gxYH99L5OzTifp01uPshE0UES7rtAAPxuDm4Uuqf5NSKB4HqFJbmt6qN+gb
/zZSNmtBWFfjK/HL3OlvUAb5x5xxVTZBXTBRPUquy0FylP7QIOglvmwy/VqJJK/u
R/yC9wYPQc8KOnniTT4AajAbBcv1Q1VbKaYVuJu+RAHkZajJvMSExKWDOWt8ZWhB
voyTr4De2hrGYl+fKimMrPE6f/sS+HK4UidwKvpNtvJln7VoMjKuSYL6JwbJQkWO
PW5cqoGrFlvHamdSI+6neUaVEeaczcZT6GBg1J2DTL6wNqo2hWCngL+BzhggDFK3
kSWrgLQ9wEwYsthZNlOGf886hncDOAna7UFAbDjWlhtezMW97itMZtHzL0+ytPJN
HYxH3Ei1nss7x+nzNz5sfyQouQVKbMCgZG8Ki/dmGXsyXX6UkDwvvCcg7hFkMy+8
jM7YOZHfHnSJLEBtdcUrLNJLOjIoWVby+mpzXCUi1KL2dvW3zjtUxLPzk0qlmyqd
dde0hnQohvz1+DcHyMiQHf0zPVTjX7TK2Um+p1fdgkzzb7fQz1afR6qDPCq9vUi5
B1nj/yT6hQhKonvGG1o9RCoUk46HNWU+qsLWB/dBkQwFTefyuSOrk5+36Z7GUikJ
PSKghlNr0bzETcgLdut3lH41pxDuWzOGb6gKgwX2yNnMaMvY39D6uKx22uY8PLra
Y/1qQPC3lP7gXEV/IBADLkV3bVHN/OlAQ41I8Q0dPGT+udIKh83HVaiZVEIPKM8m
ynEGgYsHk6klnnCwMID83i5T83SfiLLb9S2LxZ+QJ4eFdM7JzkQ9W9n/wy5mfAJQ
QNA1/5w6acJfY8mgl6X1IKGeFa9fNU4PZ1tY60EJn6tv5ZEBCdutmfo8fh02Q/KW
9SlrBAr2qsBqcl2pajL5pszbAfgZ75keYxodzkea7cOZd5KmdNom3a+0wcZuASce
MCLxpOZV/bYeLYAp6QPguc4p6wlo9ak04cLPKD+I0ILTddLF7UQOGctHLfuF+GU9
LL1xzVjEauRLgrQjA1JJztjobEZlDvWrqDTnffDBo8qDVyz1cG1gIcIAmfv8WWsH
7oD1qxCDScceXzGFarO+jVvDA4vVZ44z2tR8sZjGrdOCyB+EOoYubJpu5YERprZb
gvyMl/X+MyRSLz0U0IFimB2Yn0FG9YRoJEnr5g8uCk6TRLkq4P9Wbcg6Bj475UVn
wNlEf63lm35OwLGxxaScAdruEBNHMeXWN8lSQ0l0zTJZ1Y2xUA1KlSQPdW1TaywY
iueCrDRkdsVjZ4DpcmNpIpR5nKEe4Rr538qT39VmKULHz0rMd36SMpLynr8GXO95
QneH1Isv6AtYrvJvyy6PhtMAOmeHH1UAiHs9uXC3zWAQPrOQyFzucrzR4Xpzwk2V
RyXCDDrj/ObeTZIKGlLwzs+xzh1Owl2P4Yeom7kPDGcgvMbb5o8Ng3Y+MB72BvzO
/NLgQsrF+QWHv4UysckjajnAY+pgtQoi+SfyD7v3RO8WUjz7PZjjZC6BxQ76xxqm
aM9KKIMLzF8EeVMJlUBMeRBr1IizwrjX6jRwYYhpRTS1yZGbbwytdvHmBMpJ/s+c
oKz54hYXWDGgOJPVdxQB/Lgtlkew1dEmZ4ofoCAg4f0hkdWSENK6rOVhclwfStST
7Yh++S+u0RDgPNMlpXC3ozG/Vi4ovYnW5EerZt7Dk0cJDXCkOrKABR787hgipDxF
Fr+OVHWK5kDPy2sNpFIOdAiVPtwPZnKSyfLvMk/pXtDH3hWAmzemxw7FYmzIckd/
ydJDtV3JJslydb2aHUmsIi/2L1ORxAkLQ/bMCsOttOaIiSKBjMxKyNZ11C8oeOfr
vexoIGW5Cag3nmdGNpGFM2DHMU3VUMcj6a5QyAJHVWb/kSTJvDlsJjXZ5o/Mi9Kg
zjWW6HG7BbU/FaSeHnJANIqEJuyX6q/dvcHulyp5E1jfMVF4y8BTen5Kw1N9s5ya
4Z+mE5o2vTrwx6Bxi9Ydt9hEqy5nMc0Gs00sWuFOqdbgwMKSrClrL891RpnO36pr
9AIHtbNUTLckn5nd3zasHwOu98EfeiTZxRRBIBy/Ky5zdH5TAA3C0W7U9pbxGT7/
VlLVlGFfenyIqRaFLpFUWNFDiunScI/VFVw0oH5znGt/eOcQ+QzKp+sDIQe8PW04
AnUC0M3t8iHNttQSdqf7rl8xxNB2P5+GBwCy3kJMUBT/L85U991FMewHKLwPxcOk
NfEh4zv2DuuukZ9A01DDG+2wwdgnRyBC4KZE5Y7BZF9IbXu1lmuDsG8BbBM5kf/W
vuJx5f3ugkgYWKGySe3J5N95CppQkovBCUTTNv5dvcZH/I6a3Z3lV+9scWgLH0aV
N3ht4pHM1W1XqrpeH3Y1PVCqo+96p4K03zQ3SjQbh/2Kds7LJgtlkQ82PbQz60Du
mCAC2kq6MEuPVMTmgaSAAswhrLvLmjPKogA7RyRrDxA+CrKRMMQuYoLr4dWG1USu
fXByUKzRx58tjT+e/GUTFeOBoI5fBnJz8X/t9G7W1PPVJPO2/GUJRYSupUeMvwLs
cfMp10TS0uLzSsHljWpRI9AsCGgcbEJcjkbZ4lWeI8pl0+biQnIPDNgtvSK0YYMT
KFDn1H4tUnTa0bj11Gfqgp5Btp5rKISWdInVVD/8S6sZWmC06Fn4l+ViqzHeW+Jd
o2lcJB1E7i7W63hzKYplGU9f0VJr4/wvq1v5MSAs0iV81GQqeJFHhUDld43V+rNh
D76lJX69egewrKSGjbntjOUipKuuwYviIcuJLvq2TwxDw/siCOqhJUR/Rwew74jy
4uBI8wohCLgWeaBaBGmeGgLROG8+f8J/4GSeI9H3DwzWR7ysVQlfwqbKQsVWdq+i
XmT7qRE58mHQeDhNcZe4JzAaedcPnPdCdPzTe8HpLTjNKAR1hrWWwRCWMJfrVxja
lbDsr5vY4dVFv4iNnS969Mr0kIcuajiuxTlb1JkYXMlzSHTVzTOh4wD+z80F/dG3
MgjVd6y5OyBue8fTSv1QFSbDXOuPTOmerCu9/eRg9Blo25V0bNQ4siRcP4l4WFHM
aMHd0PND//UUt1wkGrjm57F5Hw5pBQsIBVF1mdoxVPSg8nbQ8Yxs9KMjHG28iLDX
lDwe/nalrNLDPp6A5al7FIqD7k8mYlbtvABCDu8ynWwlgQkmGI+sIHIBJrj4eRKM
iQr2XLR/b6JkMKeCjDNyZo5h9iZQ9F2NpWjb74+ZphBoHxWGZZVdjzPxCW1h5Sr/
xQI48grdDfI+lB9e70mZshlHAPN6KPGX/FcXQeJ14XNytCIj1CFNE5Tg7S6ZAjZh
KtZv5v8wLkKLATkLR2IAgVSnYC1OzXUaEU77KofzSDbDXwkvhpOxIXxocgXUBf9B
fqgGVkYe/wgXxb33GD8jBcIas1TUIYaqKDyksRqFStQqEnsrrsJt8DQfoSyn75qw
YMXhLcrTyE3nTSP+eW7W+MUQgU2uHyJAa/Kf3NpQzsUdF+itQynYU3r+Pv1cFllu
aGYr1E5v3nFTT6aGOlrEzkkokQQuGufdH7O3plxtpiRrg94z10ap9HMAEOWDhknc
JKj0oBTYXZph6KUsGAN3rbi61CiFB4Ojave7Ns/sf+UDcKvv1s37yfThHHr4c9Wj
+BRHlcVHCTyDbFvH2f8aquyVtF+nFehG7DiKELe7oux8CL/P7XW6cP6rVEu7dAdE
L6JxXIvUtCnjwT+hdvIoZvsMiDcWnVDiluufDa57cmU7RI/53o8pSrOJLzv1Kn4J
1fre+rhSCFMu6mSu3UF68KHEtZOCcaybbUWhawi3Qwfs17fV59VKWp6L+7u4LCWe
bNHGNyuTYbn1s8kZ2fdRtyjtDuwueCrAhBV1QtjVB5XE3LWQhiFkXZ+6jI6v9HGS
7qGY+qkE59GeTchPSrRrFC+SdfBoPXnXlINE3jm3659LQ+mlxfjpL2VFjPUUThy3
ZGVN7PfQktpDOsHNPui8YRCny2f6XO7mT2I9UTVQgCehAa/n7je4gzgyoBZOVuU4
iHsoDkjj3miCPjPb8wcqtq31IrLsaWt6dtryOGyz1X9RzMb5H8waOSqOo4vn38BQ
tsCVZEnNVpeLFvcFOvYEvhLvJv86oW15wanGBjBCWMwnF/uIOnUpOM54oq470uJt
dJSn68afFOUM5AifY92lTsMUzLCOG3nwTqExnrEKCIEryEs4rQwmmp7sE0YYWv0W
ppsIN/CibfIcPIYDOICi+fjTDZ2WTXiuMSBEB6ra0VmORVd7AF3FDm5dRkTlWSsl
os/SZ6A8hZ9KheWXzHyg0mbHM+w9ZwwWUi6tJrBh8ypDwGSI2z5b8enLDaP7dlFc
FArDlEX0jA7iKSw0qfUcq//BJsCZ4tYfBtt+KRa2AYGw8g5N56SJjVoA7sieEgey
0j9A4LVS84UbYnE7qNyc7AIb/JuFMq42rHw/GwKW0PsCzAfWKFcqdNP/RzBpk5BC
kWIj4n8HiKfaT95S8ayCkQzx13AwKtgLDrIdkwOvi3QqeMpbH5TQHbs2GLelNdlJ
SdO0ZGbxYr84rYOpvmdHafuT7zSm0PkfuzOTYm9C1j5bOkCzlJhgfW2gXlmXLA6/
2ZbgXJVKZWyNm9onCas6q/Vmqxuq5UIfWpt13wR4ZcjjShg7+euv/wnI8ZR4RcWA
osmfTWEu+hnnvmt44t/wBuOvyOZHcpr0bE5xNw2yQsZR6GDFza8XALv6C/90BpH+
iWMZgvixwkA90SGMMjgQ7wV+FU7deysxsxQS3NMUJJQL49sOekAJMypVLpvo71De
OatGoBRqmIhYdC9IOto5hCFFOgXbRq/B/uIZaG/DIeOsyt1yZ/H3xpuNhbOn8fJ9
/zGZaxr39q+XoHk0veuhOtf2YGGDXK+QPA2Vyi/f9o/9NLsKHBuT8aqJWPewDPen
X+5lQBfGjCPW1WxilN+sucQUnRzjvRYUtO4m+UQapWG567KXX4shcBq2aBfAHV17
mbUtpjs39187Fr4yuttX4p9p7k3KBsLDzrZGnSw9dfUfhYaL73kmaNq1OD+XfcC2
qBY/7McwCJXs9JdL5Jf4pwrQIu4LYvF3ps7ewVUzWo8RHUfX9fxzASZSzW7xthLs
2fbNs7Jr3yJpklDBz+p62aovQ22SSDz3rQwhN7jUeV7rP3eh4/7CWl8mP8TRU+JR
qVaByz/en9Jbyqi82Et4+iDcNigYfyea2b3B+u1BIPBSfEkRmzBAqNNuda+5en05
LxrSGIIHYsDs8MRXZSEQPRithqRrs6uh7ljQIdo/XuKIpmwCdyHU9UjesBcj5Bs+
pt5CVidENWCONbON4kenyKBfpR50Bh1SBqbPPY+A/S34WXf9gl8S2AGlvvCQEHea
cyGYI6sP9H/tAoVmFxo0XMQL61fcSgaphmzlpLQDP5PeSb4FdiQvKYhBEWEvum7H
Zo6ePIHqlmbvpPizP5TRCGgIoK+T1sK5eBwoWpqrE+1zRdW2szxxQbDvF9Yed5Q/
4r65nFBKUxgEJ+alVhp3E3a0xorcQSAq7vBGLG72/HPeQUp08cGr9wQsHEayNEaa
AVT4pkfB3rnEFMsfXNYv7MhZFMTUCe/mzULK6Mu8zNiEvjeTns6UBcBKucgvsj7J
ZEeh31MAsb+up9X/sqZteVM8p0evNRXqq6EST13FY3+1g3FGXtrd4qF5olD/amYl
KRpx5In4jUxP3sQKvmiNUzJ4rTVGKaM6Mrsz1V6YFJeOj7txnt3d5MCIk3Bdm3kP
pwkjGc6vSsyQzkkre3AHEeAippCiRCAPVZuv8hbA36zGbbiG8/at8xz/Rd3IcGt4
ZKwaDuXbdrDGziDuzwTpvSABO3aPOuPAcV7cfmhXZfcQxduenhBsPJIiTg2d835I
7vdadVoysaRoheF0hzoS9uTJbEW48BrOyPVamQd3cNFRxwxVBCvmYIVmaqlUgj3l
PM9XsEzqLjEjIx0x7D7dTTAsO/ABhoychGPJ6JhCNo/Zw4rlrEDbSih1PmoqF5yH
C3evOxPyjn+k1f/ciLwJfDmL/MfmpZO9PtwkR7d3dKjlnBKrvwYcXjMrOGuznhzd
Z064g4lzzhcciaPBEYBalimBuebBLw6oLYwmcLr6N2EZwo4xVDpDxlnzyHySe3Q7
fYQeYnqIOhZNPaeXKmk13MeT2eGlbOTAEefiHNI3zC/yOsdNC3k8yZH9emG/XCk2
ugvE1XOmAoFncYlE8trEGUsN6NIeOMG5hFHa6INz6yoF/GSZsJtNgW4+N7rNjvaT
OQR7xyBd+G9IO0DSSA5Fo9H2HXL28xY5b8hPVir1PFeOXfXJNCCemX4cF/XR83+W
F0Xt0zhYinAK7eOKh/xTdtY8mLLmfyglca9HP+DP0MX9NHg3nuGGb1KVuN0EQvKn
dpk7anzZhWZGtRUK4CsNxMREcyfnEPY4OhEX9DfZAbLIXaIx8+naVDtYRaN2g4tF
CXdpM4OhsSZ7dSkbt98JHpc4/wt2cI+/DKSnxtRaKL0pKO2OmeS3Bc9Przzj+rdU
zWq7vxY9IjRejH8Ey30UfADpxXivVSsJvlZD3OBdGSC8RnR526E9UavraR6cVmKX
WCeD0uPZqoyT9rkKr2efmHy7xWSlBB8z2KlxHxbCnFB/kwZExq8dDmHKvameCMo3
6iK3odc5YsQ3NQZeUMc7LQFTG+jCF9OZdIaCcxQnEDFJHehOSCsr5hQWxnIU9dE3
1yidVx5RvKE7mrfVt2FxQnHl+Pf10RR3CeslqBgJDF+mja3rNcz8xpARzStXWUG0
WOVbDeHJasx9EAfMN/P1xJ3FW2aDCJz0f6vQgS1xprSFVo5pyoUExA/o0HViAPcq
lptsJwi308eIq+54PAm9qQk98jWvadgttOxjDp19xayZKOuqNasnSRnyhAno4//Q
VbJuAvenI5zfiqneXlE9505KpR6IRc4tzxp81wmzk88Tqc1vNfXapBNAhcknua0A
FClQkzfVvsILy3q5SQjXjlbNt006ZF1W7+nsBdrZQ/byT59SoMUJwn6XDQawOtcy
skg25ERPTgCo/YzwlYjQUXmUObfPQgDlMs0+oS2DOYFr9dA3+SQWnexLKT617xoi
UQEXzDaxeZmAbpclhXT2uXWGzAlIvo2nUbXDm6m9ouihrQVmgfRi5fiyAoE/NpU1
scM6O3whZnirp4wnzv7vdVm/Rivd0RdFzZvrIwpv8LrZ9jjbMqrrFFFmD4SI0ZWd
ZBTqQI8s8EEP+4SmnV2F++GOmzOdR0ANUSejY9n9M3GDwrBa8c4e0VTHNOgtInTV
cq+Ab2m++5+ctkQ/Ipv4e/NOnsDrL99zCUVP40aNrRlxL/IBtaqJ6GWgbrFQcyR7
q8kGAGIdjthHNLkq0DWezb6dEkKcTiaWRvkL3JqsNvU+H8egJN8pcePrTd1ChOSU
QX97KMzJeCWEKfWIUvQCzhuV4Xs5VM/rIvXsuDBjL4sI49d0EQRHRATVhfYj6xKe
HL9bsC/EHhGiKtEmQIKpMmDFFo3txI/wcTAiuN6MzDSCCExnZZrbsy/1c/Ydk+NR
ztnCCYo+SIVUQrhTt+i9KYzVUkFhkmDoBSGCtnJGvKWFW41knokAVu44EjdT9IsD
Okw+enndcjECZc1XQFirMTSKZjOjDIO8yRYZOjeDbpUFNGrDLlHPB8yfWBYoVuLh
UhImedu4DD9PWbPDpiZzaSJW6c5HViPDh3P02FOXY+gbudVs0k1T8cPMIh+5RCQp
cDzTvBlt83UlnYdw7toDW0RDKkNnsLvMe4NV9ckZHdndbyxmVvcGhg1Vk3A2cF8S
q9U7H+K+nik3D5lcAzFepJt7aNBpOeFXLXjzwqKFK3g/jyhdHQkoahBzzOG+/XEN
Mz0lltwy/V7Wqj0tYsgP6yDo5a/Mj3rUWBQjo5kJbdqynBM7/lIymyJxbGZNuCK0
NdpK+FdeRapWVnw2lghvBLxsKm6hg8c3Od9tYt4Z5MvgRGq7LVAgKs7b1672zXht
87q/OvBevE9iRfUd74oUhDEevda7blKCICYuVZ8MYUvOGsU/tKMHRm0ZekYsUDki
6wtX5jUdk8WsPFQBCALJgDeB9sVYmx0cyqH87voJiCuq2UcuaZOcryeAPeRO+Eru
8oCJQ1JZ9tzuEyg9le81XTchFtOCxufu2PYLlOh9fFDANjEEMiekhtCekUgDg7tU
h4GnzHnTXfYOt6cosPCRfn5SEuN3AVTO9p8YAMXUxYFkGX9hOzePno/ZriI+/ObC
+n3a6jHPPdkgEZj4/OvPk0QWDAE1a2YHVIt1IGe4ZjYsXBgVqc7P3N00bUQXD+7a
l9Z/wA9l2EWEIbN7YC+cEtGxh1qw1ITgCd/Rp+2IaZtu00co+z5Bb7R62BjdDpw+
OQDRBpU27xeKyYHntoG9DpU1Fpz+yy2QM0lJ//oC3GgLBwyi+CWH1HDtTZWnj6ap
DN1c758UWP+YCMOXUTn24UQQ7VG/6dMB5Cg174TMYFGkBVZIcIGg4RlcAOA8XLUi
limxc42vIvnN7djS+0LDcLtddbJLJ+VJJZivBN+VCiLudG1wlABu0qoKGBBrV1LO
BM6Zy9vifjhUM+Y2BjbTiANca7zheOO2JOdn1sC+x3IyXKv2llAXFDm0k5bghxXD
xm6bliao20Sv1T9xmwtpr8BTq7PfNFom23hn9JRND7z21OvRET9AY5y+SosE3z50
sKqjcyfvah+oEjY3FWuBATVPM2zeeqWteKrES7CkZxbBRh3JhctCjZIVi3fscbPh
cFptujr2Dpebe+ZuQPCLbhHsQOeUierNJz945D6wexBAcFGCaP6JrW9galemUW/+
TQ04pJrRCklVUrgSloqxKFVMQPMPjpjiREkbOeBWS8e/JCqTS+AoELOy0sroV33W
H6ZFWG9+kIuDVsgGnL8PWTfxiE/DqHw0/hUcsKd2bYrDlTH0hhbpTq6UWGR1TJhl
gEve1jndACOkiaoXq59I11tCuAXgysY8uJyVLA/UlHX5xBN/gZjx2JMGb2BTzMtk
Qt9Yas3JEv47ztE71rghq+zEJlYE/rLO5RtmLI7fRV3OZ4Ar8yfi+36j16oiNgNE
MepgeJreJXXad1+hXrSTmUgLIxhZ2LPnv4gl4RK9jso+jnycmk4ALBvkPbbReB3o
/t+xtzHKODyCTRk+LbCNDrwnaxqt0abSnfMnugtTnlDbzzDTsigEbURZoQbIp5jZ
WmFJZV0HaHvrT9xwPggNaXs+iLk6TtUKXK2C7b2l40/u/sFiJie+OTs4CrWgudse
Pa1EdQIDDgWgono1k7BcsZu7qwMxYT5v0ulW14TsE/FU2r7HdsXiZAILoJObz0+f
/349VkJwpdEtFHLTuQETEi03T9bTc/W1NR3H8Bd++utMXtAAoXlbkwfdon/9mefm
iVwBV+jjeXRsrzT7evdkwjHRh93mXwNxkKWm+gfu3yWRHG3Ch9CH4Tftb8/1Lfwt
Nqh7jnxD0niM1/QKS/xYoTO4Irx+kR9qN29rWOgX5lPtu8xVRwFOgxRdPuf8Fjal
VTD5xzuAn5od3KMi4rAR2GbwdEqUkSjQSpUAOcb9jy8XeOhNTsQVjokrrCSKc31w
N9oUG0w1Fb0bd7cw7/08UOIykIqrqzPk57FL90n3wogSPZy31NZDEDp06NLb9vRp
Yc8bPFUO6reuIweWTKoe7PlcwySEd9xDZzd8uAofFvtmlynVynF2cUa+VVczX+ih
WRoSu4HVnxGycZNp4MWAc83hf+UAnPZ/ta0V3vXiW7nXItu+atrHGx05OwslsBom
DJu8XExorwordAOwDx7SqX//cTLWbpfnoQyELVkcb59jysKm3S03HyKpR70Gtd4o
HzmwWJUiJkEAc15QmfpYAeYN8EXdtZPBKSIR4JiBn1zXGkd3eRWXVBd6Tn2TH/9N
weURZkVVr3YgkSMyWOYgUgbAuY1I/eV5G+PJArAUDAZ4y/zrwxBvAdrAcZRhzEwD
x7l3BPeSZDW8/+9Q4tFLx6ThFHhdcDnOHWgVyQPSANXjvrFquRIqhWhIShCnwGCe
U34NJMshTS2pEM1+EhKGe4AkDsqYGKSvf2TgY1Q9qfCHKkbaysHpsj3Wm/fIGxZh
9AAbSV9zvF9Nu6v4gOytECf84lYkjwiBjsGL0ufmzSk=
`protect END_PROTECTED
