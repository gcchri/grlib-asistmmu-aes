`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hqfzpBmY1upC9uKYR30q/jvca2RuI4kQCXqkKFjiIQ/z/6wXYjcOXypgdSXfldp
szb9fwfTgFTvGuVVYJJ8Qa5PKpHrhcWq1WNNuBIaSB1v6J3EFl7S2QKIgVBZz+N9
IivKJrZ+d9c+Y7oQgIMF25PYk2Wd9TDXF3KJB7hObPsPFkg5tiUVzJSbercBU/gj
hOvixkKU+Cb+i9Ep38213KAHGBesw3qYpxv3iE4PIxE4uFCGKe80caOFnyrgR2sm
qsCrX1GxPBsMRqLtvnVjHVrW9v8c1Vmk4HtAcyJOi8tpuDshMEt57vxr6gg92TFn
XnhooKyrWuJ2Z3lOzSoEkZwJQjJQHb5r1wI/P4LQgyg9TFMmeUs5T5IAs4l1z5m+
oYjZf1QfBeBp2f8dDGZyUrErjaDRg2V5k62ewqxoJA//b/AJ2Yg6r4umRFRFRxA1
MmD5BsI1MpFRbXc/CLRBMeK7ssFPfber0QjpRlsUadjMoC3c5HedRLHuZ9+zQ3ZE
ZEqZ0BlAPt/+A/0iMZtl2al0LzvgwNBw6cb7XpMJpcTr60OjoZAG06yZbZ5fCYRu
VrW8WMkrZ1KSUunbh0qX8cGQ/RfA4oMLRQdrG0YWqGdB2iF8MZKS7uUieytpW80p
GhFrlE+h6erol1hVK7DEtw==
`protect END_PROTECTED
