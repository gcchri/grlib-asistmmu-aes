`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJlhKR3SOb2Zo1IKnl5GJqISf+JK87yPeQ2lyZkvVa23DFs6hKCyC/InFtM6bg9b
rMHSNHWJeyKeSKnOO/g9i3qONzx61zlyUGrPpWyfHVQlu0nV4jSMue4OIFuuUReT
8xbRh/UPzWuDPmDjJ/FSXT4KXD9o/BkJ2wH54XMZ1/vKWk8eihwEOzEllXGqcxzj
PtFI87cYBy0idujw6AoFTz30ywh3FFjl0o7d7fdUYpYXZhkKFh7oHhOLtKf+Qjl9
7UlTL2mvdFq1JTsU+0AxWF6y2BwH2NNsDQ2iiIj7cnjUhEIEOlm9jpeyL1tIhbB9
pv70jEMMAjZkeHF2jexoRRUF5Kl5n7PWYnlG9PBYpmrlbCTXe6iOa4+iJ2btSN9C
6vqP6jjrUlTlhW9ewr86VA1VlDg3kGMpcyy0dGqD4utHpW038XWXeOl/PJdFu6g0
JtNYVUXBEtWTVA8esf4yhO5qEX/bjlsH/qzqrkVovY3xPsCm6SrX0pUdpsnJBfNA
bCBLAT0swvHYkZCILAsZYA==
`protect END_PROTECTED
