`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9fb/NZCpuMU+alhckK65ieE9ix1S72ynCDXv4YPuqNB2nUv55VPMfQfkMIcEToN
8cO+gU2IpA/Tz2gBnuZjbXos6OYGwEbNnH4NygNHfQU+JcItbk9GEeW0I2Izja7z
UbZPan19AA/1x3KcHuWirqFaEKqjJMpA/MU2e556iq7nQfVugUTVAFzRz49kOUH2
Nn6hlR5h7u+SAQlagi6AevQR/WyIf7bqH3f4n/Mw1Z+75wE3IZS65aV/koMOafnl
di6iPAGaw5BrQ0KxFhtFvxC4iede6byQYvppMVAF1mnXKVA9Jse35lGFe9jJ5liS
NRcqVDL+ZunLaAzmIsAMUR28bYfocIbYO4txFmnSrR2WgwSSu1QM7wz0BSXwU9z+
mMowTdQx3ln7lZjav+yV5fppo/sXk94YUGNGAJODXjkBC1IftMYCYQM4lXt6qyQT
v9LkIJ+EHdKsprpVuC7ufT8vnSj041UBTH4ZrkJ5mSxRbuOiwkwA2z2Y0a6iHJ2b
Q9FEiFgKwFmu/9vlC4RUXAQPKOCJ2k0I0j251/D22UkR6MhZQ45MQVAnYTQDVDgE
EVmczciF5D2kfS2oEw6x7i0kr1IEryxMNqj4AYRDwKnpSiKGBbZGlkyDdUVvx50A
IEyExXAFSkUGWlSY9O4DwS7JygNjvCCSMSUQQLPgkjcvTE6HV6+o2/mObXZgdPpO
rPVrDOBL0FY08hPRXpkfNfcD4XqvoruGxklxBweeuBDl+ScQNvfjkZzkiiD7+BCp
Qmf0fskgA7S10PKO1KrjMcV3JHs5pp1XwtAhbSfojozHImapS9vUFQKRIjr2lDES
Lr9ye+W1mihRjblvNCZisqK0vohruOj6jsvLppJpQPvpgxkFf2Bm+7FYDU4CCt9c
+03cf6m2Fzb+8o3dn2L8NgHU/BQQYLY+B9e8B9PaKST1gOzx2Swzj48zGvLdspiu
70MgCE+6ZgfahcKxpKrtbqnuTmfbhunsCXuWNL5zaYcNuHHOnHhgnLvHJ9qwVpu5
fZDwZ7Ark3dXSkthbPvE0Kthjtm02UYTS2EKoELCnh41grU+rO9VfpHA0ZKLVLaV
JqABwVxFORM8WTGxj4XKbd/e5fKxUI49/INz7KcZGsREjQu46rX89FrdG0jhqkH/
w1+/7iXM6ailoO8BgRj2vfIu5BMUnl+2fPjbbm0ISYYcmVn87TshprQNbOpt3Zvg
21lv8S8GFzStVn06uhn90eyo2iEhgjB2zKsHzlceUxzcG3vpzSlLwIET6TwoobSA
gdXD2qNqhwVzYZ2NW3x0f0I+O8ACP+FS6rwU4iI/uuPVRKn9jZFgsarShCwabe7u
7XT0FiR7Ss8EIi3+gv8pyXCcxXJ8r5W9h3cfGRilP7g6nbwfdoFejrcxffDorQm+
gp+Dq8+GJLY91lIK6j2RovUiflYkqNELqIfmH/jONgVe4KlcUHraBywZghd68fpS
vXJV/DKiJ7e2lCq2Ssi6ldrBwVu3ZNWZtl0m/csR1L7SfQP3FbnoFbJWRD82PvYp
/RmmF6UUbHjXKNiOg3GoRhU9nE/Ftbp73g730jWnrXjru/xsAoSw+6vBeCPs2vfH
a3gRvQ8yHBsO44Qa1ChwOK9PdMiH9WnXOKE/UfGqwfdBqJyqnxdy0y6M/n/PhsfN
fgTcDHlcswmmJQGUJyTrdVYNlKsaRE3vzZQt6iQPFzKy7hIKk3yBya67g2aFpAj5
2SrWbSNE4EG18CMxxsTAnNwOb2h3hD3OBudUVJXhpeuFOeNtw8c+GsK1TQe1zDwg
cOuvnR8C4j544qZOvr9Hb9g7ra4WuULidfGbwGSvrlp9EdyEFoFQreBJOjF9ra7T
wQ1qmnapzECviLNEXviLp9dRflYQsTtWE3LZK+Lvy3oKrp0opeyEwEdKHv2DMSpT
d1e1qewTw+UZtgyhSiQiI0IRwbvX0hgOzI7Gj5ZETH8FiKAxsig/ygQ4AzYDPoSJ
mT4mhLuAlMw744GtRjGL08iLErk9409QWPrz9GAWa1heQQkNO4bO0n4KW9CI507m
JainsH1Yg+x6yI8ebuiDxkJOkmN1ceY9U+icLpacp9GFwcgkJFvPgrxuEaZxXOS2
quqGy0GY1b1kGSaQ73V1yPzg9Or6ZqK+cvYb8ET9JTZcHlnCr2gST1jlhV7o6Oiw
+odk+g2799PDBleY9RKKPr+L694kvKFqCowte/diHpJ6g1OyYF5WXo1ardUXqOGz
namJYvZb9owaVoScSN25kTef/BRZFIovxSjVGwt4mFjiH+jEnJNBOcUseK11fjro
EPWM4DJeixfs0zyYDmzA1Eju6UopxzDGJIleYfvSgKeAFqjezzKvcZcn7IZQDKjI
mUVlI1cbgzUXohpWAW8ECeq2b51G3H5zl++S4Cw//09PO/95miWJSwHOQJKR1Xkr
2EkSMFdNfYPKtnTgTgAgdP6tMXxfpoFXfPFFyh8yYEDkCfS7TL2n6vLQZsfJ1oMk
0vVg0xp+fdxRlzvnWzvDf+BroqsF3BX9mejcyKx7Z/GEZU7jp3vAsptASdM/fOV8
SVWqrFj/6G/gSHujISAluV2HWoLOP1mQadkJDsDEjFwbmkG3MVGYp7tDm9yzfBFT
6quDpAyStlnYEIbxEMBy5vWHl2CiJCTIfMxJFMnWzex1bW2EIAGEcEiMeyAQUvMv
v5stYBDFYlwPnUC93//3RF5k7dukkRNeSXNkHufynw/vnOHREyW/E+1fj1zpdvjE
jyHAN/TlX+Kqol+tnNfpEj10CjvXicvd0KhBPLVmGNTEEB5PSkupy7/MlDHcyo/o
np4ungcAp036QCZR+TyxR0gdF22Zd4gosBFMFzN74OSVu5DYbAXeWS50ygPk5ROC
VBION7AS422YnVQp2XGyr/yA/aiikYGrOcWxulCamVnM09HGFtDiFmqmJ6X+UxCT
PEVzk2HvtPrkgdCVTH+VIEncGf4z/M1OTdublZ0bj97p5fnDC9yU/ygW91WRop5/
Jdcxnul6qYgHt/yBTIzACLANsiYII5SI/DK0ZHsFfuYUng9JPMjrA7vvKr44oeVR
wd26glq4gpAYGZN+b2jcwbIr4wb0NthtOeHd4G6npvG2omwr0F8G9Bp1zK7P+Im5
S5VBll/YNI4Q0lq4whYJ2vqQ96cUebI+XEZ9w32T+bwJQZ8u0sHlZnqOpXiBcDx4
SJI9pPOC9B0S84ciBRuo7/H9/gcQMWsvA2b1HjqfhzAbCUL3Q0GBjcGWUXbLgzce
TqkV8KtaWEzXy2ZG3JhZJJ16DsdYZTqSJtEHkNJf5Ogi/KSJwdd1Be2bVbrmaa4j
u60FHGcjZHbUW65WzcCM4lAz8/EEwzBXqkUWbCsVk8saM01p2R8yppX4e0xtRyuE
ASlbVjVR3APlqL7J6PKKEeKtxPPCEU37CxhXXrxNkw70HuBQwSFGSwcOR04YBQ8g
lQ4NiP/U1nUUXSSFCsgUTei0eyzmG/GfapQDT40CddTujHyzlapCFh3oRufczfqr
2+Gs7DFj07gZt191FOrftgYee3bNXZ3Z6p8QqmKBtE0BshlBpAtAf3EIbe6wVwP9
0SWWyhyrCJBvDBHMzmVGyaOr1sZgRTgKHCzpalpD77hQnbss+dggRnjgcoVQe9uB
t7H0A5lvwuPlTkJ9qZMGs9e+aCtqd5UwctOb9cMRGK7I/0Ir6b/UVnQOXc6FdJRN
JLxu90SmPTNvKF4iTOB6nWVGZUsf/6tsRhTLFDd3zwORc59z2D92dA2FwHaCcPX3
lwcFuSx5LJBw66FA98fzk8/0ZkmSGeLdRdgZuI9ngggDuDp8Ct13zcLa1SjgGRqH
ve/C79+pWoDQHP+vF6rDQgQp7yhlmp5Tsupc163g8zaHAH/R/BoGnOEMkiICQJ8C
o35zdqXBrr7NELSVIhzP/QRyNkjIblIuRx7hwZvBDkM6ZssMGK71GAu0saBY1+qw
9A943bc1STGxfZ1H2ylE6gB4fIEso35BtzU7Jdxx+Dkf6pPTYSwps0FbnUjrOmEU
QLYLbaDQjOkYAxgbnvMrZcL9E0ykL6KwqF/NYf2Z7NKIlMCE9FHXW5Z2o6xNkaeS
rzqnkWYHjEdxCPDhmsXGXMapAwyd0zn/V2mTRkJUSG065lxLFsM1KJ72UwETBQK1
oMJ23OARnRzcINxgDNPY4E2HgU4w2DFjD6Oho9qTvkwva/Phdg+llsMl8BZDhu+T
qC80CuFxTpc0+bBjg4H5/dnZ0AsFP7esL/UObp2lvFby95MdT0abBekbBxGz9iQe
26PQ/c/3IozETvrphsXER3/HRcQ5jGPz/DEMiDRQLx4Pv+iR4PeZb39leGky7vpM
GwD8S5P9FehZnzwq6oQJhuaDffYQbdR3iYW8DsBiicvtYEjg7DonWqZYxS5ceW8i
I5yxQbmqf5pjatksG77cZLWUjmWiyDWULXOQnRAI/+dLRUaiR1qxq/yKe8s82CGI
nfIL4Soze7wbUfnT54thrLzd2X5pCe4GxYu/mzX6dUJh30akL0ByrgZrrgJvU+DA
i3EfJm2Zku6SCDDEomemj5S7LLWojwuIezBELz3M19G+24Zl7lFYgntPNaqBnyF7
gYPKecXGZ/rLuAbD3m9smjxcnvCiwd0kEHKqxxIFzDFvn2GWfmLDySYVMpDz9bKI
99LsQtjgJhZ7uQTXAZRpjAvt0Etc79iATvjhLkoVYGOE/mHZJR7LUmDPcqWnK5ZG
feNFkufwxy8tWFGn1hm6KwG8OO8UGi0pyPznvpRs0XIzMZbqLhnQY5y4Y975RkQ3
DBZhgEevL4rxDPEV4cuHH1S4Oi2oYGyfeF2pDume1bZ9n2RBMQe61p3nOXxucm5x
cYZ7awfGzt11QKzvvUOFxl7ZQF8LP2H/TTV5EECFCiEZrVskkGMc3jNAowbgUDqI
i19Bg0m5prwKmIJ0salZLwfm01+7oGSYA4cFHjlPPR07nQ/6K7HY3IpFOBGvWDP+
870kQFXIZ34JfC8zaRInQkyaQQm3jw1XKKG9k8aSXzYpnn2Qhw//N5bolZtljBad
2u8AlStSLPGTAI7vRmk2JGRJTiYrlaPgolI/6FqsEJtRoYBTG6qcbhe/GH7UIdUE
hJ0y3TrZU5P7DS8d54d9AQ3SglHOR9ZCDIm06dR7+LA1Gkp/DbvPp4hbNZL0uuNh
XB131gukUNkCHImBAIXEGZLEWuaYaGuo2bOcqkvQXGSr65sENpXgX9c+OvYiKZDZ
rs0HXq4CKDkn6ByFJSbFQlf5XTxNXE6j1Nump9HzOhRHv9oEo996r3w1B+Q0uQQV
Lsv9ak2ZBn5xcRG1zojyv7KMXE03okh9UeRJKavoVuQQmqCTWBx3+u7oRQa1wvXp
mro5eo3Pej4oeLsiZa1khApmQEnyH9S8kLBkMXKRtfHbSJW9PPIq7zqSPXzpxDB/
w3hry6U1qdJAy9Bu4K3wDVKMoTNg+jEN8P9dGr0rkbKtBwbVXLE1Qxchx13ikpx3
`protect END_PROTECTED
