`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v48tAfIExDUfvr+0vdlCs5VqQ2Mob4LkgU4fK57xGTlqP9bSes4TDOb1JbJ1FvLB
MdXizoybm198Qxcvj91Zx2WlH/nQ0GpB9I7xKJNR3PJMvpvbD1nxdm4cP+HLSf0m
5uZr+Nw2+THghkfMeAKHooSzd2FEiKtBBiOALbewCMLrmItlj2gMkC1jEdFR0v19
wHMjAHoPMy+fq3B1++Xf3L8Lxpk6q/FqMHRnHxyZHRYnGQ5E+BrdJQmgR9WSkVoA
Oj0sy5kHN9M7vbxVgSq2sgx8mjsv9ZuhdXVDCqz7dVEY0KjDYXPnC0w9UChfAiRA
HAYzX8Ec7GeSBw59hkvfcbzCIUYwY/D4mNEYkVwSOcf2/EJWytJazqhbXmV8U1OR
WGBuPvl7W0ZhSi7/7OXTOmeoq8idy+mnihJtjoEF6no=
`protect END_PROTECTED
