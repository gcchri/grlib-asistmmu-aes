`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SrSYqjv046UuItpVw/b5GQB8qbhfOl4DEZKcRej5GaKU/wDvVq6bKAlB3PZZJGP5
1rvwub0HQm7aJnTpE3qWkxVAs1YgTfNFxxtrCYubwRADb5luegKS6WzKHxK9AYSr
eTc5c2suoGjb9TrUfuhTPwv+TAYui+AE/QcPTqXa3atiWM6+wRjFdtvyrcXM5QNh
+AkDWqI1hZmDORwqR4y39JqXFsEgiMvsmFT4YgXPG4spa4gPxXrZEVV4J0HKOmiw
9ktUtDOLOaUKZlZhJPl4oG2TIYm5okCf1FmetRh4Un+QY4o9I7+2t9xch1nx15YC
7oLwJ7uL9SRsH0WfJ3Mi5O37R5F8aKIPsFvm0xs1DFXla6UYBqtEW9O5lUwbR7fD
H5q1oEfoM739BOsi9bcPE/GF9XnucSwLimAWgAG9kVOOMFNJFJzykoSt/EQeZFjF
97UP9vs/KcJ3kCa8MPVYaDRNLoxnRu41YomF+Akz5z+KabrfxVlH6b/rMRt50xvw
87GCzJslhlBdCDYSN/yYUgZkoAGWTe0sYN3FcJjgjdLoXnezXPPRZP8odxXNhi1y
bbKjEiV7QrwkkPpSe7TL4MoIDJwE96sBWwylbD1VVCdhP3gqO88zze/1v7vzgoNv
AI8/MlYCeEldIPNUJtwAgQYIHbK2t9zCivPyGSjmyzCh61Qmzf9XebxHk1Mp2gqU
2sVqeaCykwKL8KQ5OQVdbCLKvfunTx4Y8dhkmLX/Zvdzf4Th1EPSOkbSIdjOSsJR
9Ku08fOBjasmsDpNZdND8A==
`protect END_PROTECTED
