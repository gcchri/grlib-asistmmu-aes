`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTw7DRy4Q2twBkomNHKRJH5kPmz/JcSnBaaTYfEq9EzpAcCzP/XkIuk2l+UxmisB
NXiuhleTXHKRLmxj4683ObyoXvQ0/KqO+OCtkjdLcf3F0zyM4uTHsHqdhgFKPMOU
6yvuCe+OA9p7Ny3K9pq1uCxNwSYEa0CNUdrGkYF8YmT8y4IFC8jPXSlhHc+/o76e
cJpVqYOMJYDDY4A9oAgjBlu4RPMEkTIRdSsOJM9IyROsZfhw4Bm/eVTWZTIaeCpz
888dYknck5IcmPJY3hqa5OWdASVKy7onTa3nFSLOqzgWsB8+tLLC4AIfROxCo7t1
a1zdJ0lggv1m3Q/dRWAj55e081kHdGhBqyQ3IW5+YNLcnPNxherRndngn5NP6LWa
M1W9+HIsLOzt+9H6si+1P4zYfJYYLFKlAYJ6qc8Oz+M=
`protect END_PROTECTED
