`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRKaifl4dUYndWkLWHRoOXmvCTOp5AulCQSXyI6s/Aw4hWsJBGgRAwNxrF7KqfDH
LBQ4iP9718NtSBUoqNWRfo1g7dOOLBx2mbyimnynHEAv8nJD3Z1fucJR+7IPQoDI
8JCl7zE1MbAbNKh1UL1IVzbe8a7l7mWOVO9ce886Tyqbc2UPEZrRKCTO+ooE/7Yg
0EW2rE+byp0Ei4kFzfAMegmxeP5lkid1a0pVDu5Bdn3sIzCE7TXOBwcE+1jJpzlS
jwl0CnSwQaufLQbtmXTA0g3v76qym+1Rx3DYkQh+08Jc9CGEExuFzhBpVPSGoOep
D9WfeaWp6uu2XUw2a+IBg/PHBElfVPHvrjzbABvQw7SUgtrOU6iKnX5qceucd3yG
0kKrwQ/15k9dBclEgVCATfS3syMZ699lpdAwQFa/HV3TlcSUEt2yNh0CxQqXIvgO
zdy+7D5Ksv1SDu9BHCKAQA==
`protect END_PROTECTED
