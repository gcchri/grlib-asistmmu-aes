`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/nzns8XGwOqmVltkA3FaA5+imQ4BIPHR5CAyxuhggpXm/MMGA/KTLW82rtFCukO
EhOrRjbz3TbNah1wpzOdK/VvZD5nmHtZ1r3pkEFuDrcqtxibKp0JtOFzxamVNKQg
8edKTByeB6vt/p/qZy0EC8wDk9ilaLrrG+EKGoWykeH9SrrnpAZerNIIPaOvhPqy
VofLeMY05CANri4LeXQTgK2+r7LBC+JcGcG2FiEqsjM9z7of+bbRBdC5A16wHblg
5zfuYNG8KZqxlUaQpM9l1gaj5JLUuEun1lRZg3///34KRlDN1B3wx6sBLwXhrfJ4
LnUdKrPBNtxiNjNO0IAFA3SJRxKKuey60VfGg1EMpiF5MidArlSN0iw+1W+6ZvSg
TXwYvT8kAM9kFsq2qSk5mPB2ghzr0zTWoGK2/8eSWIXFM8J091cF0wy8ChTWw/8i
4eX0OYog/R0Gvp203wuATbBdq/IZxUSSw2icQGruQOGJWXVOSRCD9WesEZLbbb09
8HLfp27uggxCDDiGOnHZBXAEZDMd7xVwCwnVEXpHsw649sggn15VypJd/2s7bGxt
z7bOkEi1c24/X+KQ0Jf4di+kAxxwpW+T1dYrLQdLpUH3kR7NSaMxBaRtPEUnbg4F
A2qPnKWXCMCVU8XgqtBiiJaalViIU3VpSZt9rqtZb+Ra5jK73c3RZCKklI++MbeW
eFWc2tv5205HZ5N6eP88Sk85hSx4qU9G9guSE5ShutRVQfPunww7RoKOEmrNEWzt
1GcmEjGf1JmFn5qodiGiL1bbFdA7V83Bo3pT/zcT7l4XmUjhnl9AMWMXuGgys99i
ZjULyOs7LYwtCgnv62v+6iCVX96FxZGDswXMwqnvJTWiSiTKKnp/b3P6DRI7FM28
LEf2RZBIjPyXxHXs1MZcQfuvdPfpTXkPMCkL5AypK8LU0kfq5KiD4F1lXgYq+P2S
OQp+LyYo/GSz4Ml7mt3X25Oz8QssBwVNefUJOR3CpX+VfKsgJAkEoAzaZyzqy8NY
lS/PtBdCEb/L+1SYgjqRzbRqy2PiwlCpV4qD0Pv3Gx6iqVJdyoAYBmznOBSAxZqx
MnHfuhIkdT/rPf9q99D2zna3QalaIiJOKznbhfKhMTCIANFE6mDTOsZtDCg/NVVR
AqXsCZR1gPe6WuAyIS5MYUP7BWJLO8rH4337NOARz9N59CEnzUhDhKu7Ys1EcVV8
fDpSwG1Qa9fA8s5BbYxFzHUbKzS/UN9v3Mpx95qpyq5q1byGPdtTMJC046PHTrLr
Tv2dKB+dlJwVMizgD9HOVr8x4qat9IVASxUTX6mxTPg=
`protect END_PROTECTED
