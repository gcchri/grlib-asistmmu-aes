`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKczjA5U29Jy06sya0ZNy3tCMCUMV9xn3CIOzLVkzfpuEICX4KeMOfdfK6J+rjPh
Tfn8Q6b4VcHeMU6Unjp2V4bIfJ3Rgr5pLjuuuofEeEnUb+FfJmIggA721VvhU92S
TTuIXFCF+yW2jZ2dVE8wy0QYHK8yaNUUOaSH4FiiBFWMMSEfbYAul3oHXqprsDAF
q3aPUwOOzpIzohV64+wQixi7UHghf+qsqgh+xRke95GvNsIQpeYWgneYhjq7WEyl
RF+dWXjKxFL7tx/sJcDY/hXz86QcQKmybSHecCwh0jOBqpxChYwAEFBnyuRl5jJm
NyzdxgUZxH360uZ8AKsE3LFZrzp4oMtyxmdUXhKLS6rM3AwAKI9Y0a/gWl7lHFqL
lOUi8B3NLdlT8I2bPsmdGOG/ajztS04xZInlvzOe6kd1IeEsWxS2pKpLr00x64cr
UXozbgkJU/ym+JvvOsSeww==
`protect END_PROTECTED
