`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHZA4+o9dIqgjdeTmOj0uRvZbB9y+URfuHb2tcrd0+vo8j6R3gyEF8oZ30KA2ufF
cW/72Nl2qIPnk7Y949GXkDUUl2NDiT+s9ezpKsN1aAZJgNdvYroEOmrFPj82z2Xg
iT7ZVnWrW17+CCJnQ4lAeuQp/qHWEakPFi+W9+g4eVHdpolJ3BjNDodq8cdU0MFf
Jcjk2PEtFvZJ7xh6mOyYklj0IhhScV7gsz2Sf4Lkn+LYi+l7KPzJLxhLvPckTUyx
TC1m/DmqKSlSmmGMX3SmRJTKSuOBUxZVI4C1fbCas8PW4orSCjfhocxPps+kG8Bo
bMXsbPVROOon1wXmkg7HcAMmXWbMmqL5RfQbjgw0JnA1a9ydQjU5m/VJbnvuIWwe
87DBmdJPCatoJOcr0j17opTvZzk9zyq18dQX0QbRYn9XNJ4rupjFozbc4HTeAcY3
UqlFGZ05IiJi9/l+UM2/MHVKyADW0GS5E/TTEY5+F4nw8+gjzweDRzorWhFBO9X8
EcOcJpAH/qmjlbYmuDYXFZLOSv+1oZaPv5ZT6pvnLgjxxzhH0+j+gXUefkaYmMS/
eY0VJApbABBmv+fFbp95KO9PBe5lOf39QmydjayiIcDAKqXODefWzqudc0Bi/T+V
BeMdk6q/5J4wZfEL/kp2czMneF7eDB559y94x2WH2o7oKq07CIDhMEWpzY9+0z3P
ai93g0+En8JzLqxxRBFdtASpIEEc5ovqJT9a86JnUHVXWL5gjnc2ZW59rl5Fb/uS
e0Rk4J+NMHj1+FAzY6D0OesyQbxHiQ2ZJIPtEWlTOEW1jOST+secHSE7gQ+qw/ZU
frmBuBR6kF69pP+QsxKGHBF+VMDsOADk7nkhg8V42wclCVXEMfrA4/Vbe2hH//Lb
5WknRZsj020o6xTfHyLgQoVZMBrC7+lINwDnMomOUDHAJZAhguTcu7gcaqYUrMJA
aZiOjPcABCFVVZY1rWRL44MgqRAuXd7BXDQ6THoBkSTPuvBw11kh5SP8/yrG0TSU
9JDeyCbW4gLFsrfaiyBdNmUCsQJuctjfNgtI9DF+7DJvzYiHjIxJp17O7wS9uhjR
rmqz5YKepJ7rbRUdI2+Gwae8Pt8GPgpJE7TyGZZWW+eF7jSlvBkuXLZ6X1wQDHce
a2asNyHGH3pkaSAfMAv/0/h7ryfviW2JEvY01fKxU6QGdkULq/V6BhzupZZfstsC
10X3l0DOWYjYS6tE//dB/g==
`protect END_PROTECTED
