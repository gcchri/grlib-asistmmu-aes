`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sNUziN4OOFuA/3r5fKz/t4LzQq3DDzQUDcz381Wpvr2cIzXnTtd4GR/NK7iWTAxh
Az+xXdc5GNXGvTNMbZqwTWOks7bQTueGUBbDCaAg0ry6D/xDsnAKkdvd5b/8wMHP
8ep5wXwX8ZnLRozfppAUKJdM1Zap7QxhmLJHDElgqql2C2dg0NUInLAu3jxHroOm
ZmSNFRHY3PnBYCysA7ijoh6H76mY/kaHKKOS7FXDB0I1z/lV6Spk7Q6+FR9OWDl2
nLtWvFETpe79iuuX85GcRF7R8uZlk4aXYKtxo9y/lhJI51wMWu6npDyfGsvjxLhF
OQSrb6/E5cc+f7RbAtxkQER9IRTgpPqLlOBBwgrjiCLT5ah62DjNED+lurpzu2Bk
`protect END_PROTECTED
