`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLQu/hsdFILlseobEVoRkcMvKyf8f7t5W8tHUGnYLUJPj56y0vHEjzEdMO21bxrK
e16yU6GZd06bp5Pw5To3IgI1u+3QTJ7wV8zyXqXYuNDaNJ+q40kZazzgMlESCx3I
F9AULBC7xY049c8Qcn0Sn8SaS20tHlTldhnZiJwYxxKtxjpT62ExUHGLD+vc9Aej
8BP6YpBxpubeuD1j6GiJ/X7gHpVBQiCOw3/X/VRddB4QvjNOmY3aTHgm+KxEYQuz
vuVwCvgu8uS5dT45qtc/xpLM1DnTK+J/MaylUkkQJJUT+vIobBASErEdUsAIlQ89
EIH6vQYJh7JHE/jo8b64NOc4qUcjdD/ZshMEcqVxYIQML5409z5vrkGu+x9Qw0v2
kmWIqwcP/fic0KkhiKh8mgxqdONF8G888UjCtYIs3Kg=
`protect END_PROTECTED
