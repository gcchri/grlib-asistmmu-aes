`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHhtSTf3477UK1Adscwpznwl8fcOv8l0Ejj3ilKCzFA/uH8hSWhC9xw0YCDQDcGs
5TSJqwIri13MQSos+N7NJsue0OfMKTynmBr1YhDLFBac2mfY1s0wiNLEM4d5lAmG
f5iRmVC6i+OJnc89GCggGoDpMmWdqUmmQh0Aw3YYvbnvDzPJUTg5qxlWhtouXoRy
tIgd1BgNNMYOuKBK4mfMXVX7mP173nWmKxJwGC/BD0kEnbSxhG56k3S1k4Lymcp4
Kn+bTo/OzYa/dyTj5zHIJPmQZ8f2x+FhEJuUYOKs3N7iHIKMLWRZjfP1xE4uVS5a
DuWPTXeQHrbv8Tv24lUmGQimVtJFfcxblcvA8myPkrKWYQggYxNQ0tClPVexKXXy
xwzy38Kr561YMNk8wbh4B91YGk3x4qFqImEGG/nOOVbXB7ZL8pVtYg0kG4KwQcR4
`protect END_PROTECTED
