`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Jqsg942Lgrh97TM9HNkD3wlud1FUB5rZAmXuu3vOBWCkp4SgjXejBkpbtRMNhF0
6jo4VXFnUf4HaZYLyrYUJAA84avTZ4fkqktKlnL4uHYCW2/l2ucNks6styjQYnsj
NJ80hJcdg7lStyi0/VhJ1Oslro8lnqTDPwnEsETk1W82kTmsfdHZbLSv4HOmp/m3
0t9w+GOTYf/IAPxXyPr6lQ8zk8O1i7hK1lu9xJBS2yqfCPZXn1mllpXrCrnONism
kj4x/tN8JKTFSShykoBsiKmFEFbQQKFwQ61MU4HqxsempLfOipstbgYGzOfMWqqs
3jKhixZjnezojf8PitotlC8XTeuiVQQ4wGJqnXpigjex6ZkXBWHuCVN1E7xAwzW3
WVoLHRE6TojtPFuF3SB/Q6ujWxwZpJ8LsdrH9ILCK+zTCONnRUMpYtOaJ1anE1yv
S2lsRIWgIIJDSsNJft4g9GMqb6TVm2XBBhHvq0j1gK8+phQXDnxDORd/1Pybo94P
+HWk9q+1CxiqVWw7ST19KLLXuaN7xRMRemIfYI63hbQ243Q+aWN8ZpEChqKNLcRF
y+lqT/auIqrI5iknqZ/6QeL7bqueu6Ta4ab2nVCryw2J2zBH2PYKD/iPlDpHre3a
opCYZpQVa64x+kJKeY5VlA==
`protect END_PROTECTED
