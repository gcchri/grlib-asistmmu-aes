`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/i1yxzTNWyWfMueqkDVzB6ZU6sHzPmAAgEAaej6zpPlLtCBW8jHEEa4wUgDUx0k
rihAngw6MVisXBHLlac4GScqlg2K9q1r6sEZjFiBrhlF3ZKf7SCSAy8IT25ucXSb
huUNm06XdcX3x5u5OCBH80JJxGLKuxefV8VDml/oT8HFw/38jIgiMCpHxeF1wgrF
p++fagJJkvbBgAzb885KgPXS3AvEb9FKX957lJEFiMknRQ0UzvY6q06CBUN/879P
uROxKT+id5hVSFTjcYHs8A==
`protect END_PROTECTED
