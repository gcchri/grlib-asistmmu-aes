`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rlDoQZmIAlLZzLeoychyBKSxjstSTtzM5hackAoGrdzcSHGh/Uuuvaiq0GJLJPYq
VKVWAzK6z9+VAhkesK4XFqz6WOtgECtUsuF2niJXutzzdOpgRCIzBA5ySviGE0xo
SmPecWOJMuK46WB8flyYGq9Ol5B63dckWXorEy5Ygw/zlcRvQHNkLwZH0ED3hU2f
o0rHqvgZgH5CRVJLRp4/uuoACJZAZs7QoI6mRQM9eB6Ohx71X0oeXOR5BK17J23/
+dVVylrxXmJ/aCwzadGKbb3PyyKyY5q1jT9CO9NddlfBnpLQ7LUDl3wYhgiGZP0I
tq2zb/vlo6i4nP1jZOqe6uguPQY9lrT2xkP3LFAwOg90KxTIJXr5Ak8NrTfuZ7+R
k/Z+6/8JXIzJugL+O8PoSgzKQSayKUDHWQo9oubDreHK3Cnew0iUD6X2/Kv8fwXI
1sQ4is9y7i1RF9czYCZZbC4giOWoqAdibgXdI54GekxJJ1fdjvYd/XlSSYbctW4a
kyb/CoQDsOs4mVPYgYsWb7olKvYKyl0ieJfWw2fxpP1INjql0cWVnJJwTHWA3fxH
mZQIS8U9JA8hdSf7cQz1dSXjE1AVvkqxLF8XKUJ8MTBJqgZEtsmJ4ZF6QYbMrWXo
4PgtfJVkyNZFOz+cmoa4HacE7sD83CMS3mJ0Dy7K2uJQP5L24tJdwpfFMHGar5lw
S+CDApTLuzwOle/o5VcoOsOKM5zf6LlviINT6Es++tumTDPOPxOQjmyH0ChkZt60
UUoqUPxne0ps6MegHs1KS1XgzaZ6t1yyWUdm7CauiVW389z0xuAqaJH/m0A8Am/z
1X4sMZnsuvzVEtsbC7p3kQ8Q+HOS8gLVrq8kJzU0FIlvj8zi5InsXxFmQd+Ze/F3
rF1tzPGYaxLrMOby5LuSx2eVoky1rsxVaCqspQpVVptNbm6/tiEnGojyNM5ax2Bx
/ADOgU/pd7J8o4R+Chm/39IoX5RJaIAvdFklZhzWcggwTJi0ujc8WLJPQdi5/DQw
uACvJJ2laCbUFZ8J3ilpoozlOBHe7YAhfFAez/wge7TvO0SeTKjZyJrcRJKEd/Uf
vdk+IoaG7M2OhDU8pHgCLvAwB9VvFuScF70qFdRYM00RJwmcWecmYup+4KXS7Br7
uuCxtlmf6bRVuYarfuvB+UXqOa21/nv3Di1XzUxMNI0O6nUGapC+foF5GvLZHitJ
9QNnCscZxDMp4DfJdQKA0rNNk4851tNvwLpDwnqns5Bz4l9fdcisnNHdGZdBgY2h
ZGF1FWpIO1wTv65+dg8ED1ujaFqfdSigiPT6Yc6UN6yfQprgYuUoiuUa+ymwRtRC
QZRSqSv+wI1EqmADL8FvO/4F3wOkgQZjcvZdSjIF3voXy8XivyKRFAdwQt6Y18XQ
jzsi7ellyjpMcUWIuvahbA1VJt6VyXYbsze9BHfApV+gCHk/xVyAsMtNNZ84bHHQ
ZFdONBSB6hJkcYzgrojezPjIgqnBQ1cPOuYUU883QLiKs+AYLl1KQnj2RTefvLUV
7CzrVRZ8LpptEE7xneiVxh6gj9SXMM5nJ1dJU1UQMByIXRXYtInDOngQEDaN0KCe
V6X6SdXP65LHnpMWd1KLL6LUNhRUf2W/AB7I7klJpBDSLNGNz5JiFTbqltLL59O/
2wrF0GTaE9xu45yB4U2H3ZNEj7Lj8LzN7TibT2ayF8FiR48b45NNGkY3MyORPEAY
BUV57SqfjFaEi30GOb4XJqAABCxpsRcW6hEabT2ypgi+ZxWtpjuwDUHQ2M3QIEL/
Zv+eHnOJ+6YAEkWG01VJpNgycQrI3zAoSIyUkBKc2+vytRAB6D/4/LZZgFRdfdJ2
mAlyywRWY+S/6AyfPFbIEn4W4CJ7vV8IuTgYMV9D/gGfcfHH+UTjPRfD4wBEn92S
Z/eB88k5m/V5Bzl85mpid6cRMmdNZI4fv8tnxPFPuAw7zc1mldqJWz9/Czh/z0KL
4ZWCj54NvXtfujrkU7o/PA1FTJYwl3SZ9Q2vKvhK9eZ+6tNvU1oK36bUavjcAR9m
hRq0Om988UZ9MZjk1abfYNnzenVsqQgloDIiTY9PHJLboSLi0SQguB15VWNWTghB
MKTS2DZUcry77AFYoCfkOXBamBrwaJp95Krrf7u38j+HPydPHgCv4ZAvTgFoDPKP
wCDC9NXto6uPqI0wqRnI1o1mXaNdkO8ZDzJziee2I7RAHjdkBibg/DaiMMP7Qsk/
0vAYIcGiwLZ8aRwqUpZGJ5sO0r1kdzT6Qdd7EGdb/PdiAw5uI0UkiP+3J6wIUNN8
V2Ehp0RgAhRQ3Ojyp6NyHYX5LLOuDEQixUY4pACeup7FAsEF5Z20cdBl+CT0x4Tg
oQROvoSKdC7hRDKvm8R6JFuIMrcRfhwrey5j1fHa0bGbAoN1eAB54wZnHYl2BimX
i9KX4/AIVWaCotMjgM1IRcLMvUBIpYTds8LIkK7/IuSQBZKhFh40xJNHEntC88q1
OB3ZJWzspzQ7FQylHbHgePHuZtD4jwu5gUmpTDy4oWRDD3ZaDxkfAMJhEZYr7S4k
vhZ+pGRhrza1p4NDNdN5srx4dH0oThbHV2O83sgqdpJw3ICbetDPD6hvjT76NmGN
afApALkHMg30PyNdptLCpEDoh8zcNzmxXAeWAjOMVDBDRak8L0m8PKc9DML69J4f
gzXo10o71FPGLrZg+I8bLvaQjjbqoE4RnKMvA5P6KiUULC/2hfluHDoqkqAMoAuC
3zOIf87Y26QQa7gB24DGg9z0TeudbK5A2OIsPA0XGb7kk2ygr1poMJHVIbONoLie
hJAWx0YfxQ9gOp6mLKN8+DXwdWfGBU252Lg5BB1jEaVUvwV6TbnQri9Zfajv5fYa
c+jJPoDOjfPAkKIbZfYhDExCK/fft9Fx8IS2dHYCxLp+wuEWPC/ibdvgOqIvFXdR
ZFAm0T/EQsGa6EX9IZZGcwE9wzeKg03V0HSLw9y7J+S/XpBxcmiAkRatYQPHrjcY
XKX8LBMLE64IDeYhtyA8KDM3o3jG2uWr5GBKFaz6Q3shrid48tdRiwF7FDXNbTrL
kVSf6MoFnt8kT2XdNqMxfDVBpUrflyl0X8YeWEMShuUdQ6GtASP3lxaoa5Ia5w7V
QCckP6DDrVXyZjbTezvd78ZsIkPVmQS6UjviZCVCC+HieeGgIM55y81/xRtKUatf
l0CPyVmasmUvvTqTSrAKbqzGBOfdejyfZWHvGEDVco+JRu/AZV2yEuTaGPLm5bsy
fZKB85aF9Hp7dKrq8/rWl+SVLDWQ2oGngtfpdj8xOz+USObVqo/11QumbVy2WXlG
SnMKwkLQICEY5j/sdaGllmkUzP4bSerHeKA1pAgTsClplj3dCH1MhEGRhXwSYDk6
/MmhDNs7E57uLGJNfsqrUm0jt5LI7kDmkKkit90e5DeTTUlQlSGxEob1KUKvX/Sm
MHpkSCJ+6FGG3b4ntOzrUKGaNJkOyJUf1EIlSPFxi342l0wlCdJQ2RA0HCbCehx4
bRqT3jEV+4ctyPNedsmjfqke3AnwZc4GtBNA5Lro4BAzRQsrsr3fT6f/1icShbvh
IRSQ/w711rBhA/zTr/VBLHrNjbGJtE02YqjymbkW54uLeg8QY+bHhSGUwOCE2ZRZ
YtQTyZqfGOnv6GTQaMDAQaaOjk5mCuNUvzQ8mBszFzBTrwYb5bHI1RkZzJxQjDBz
tDJTj+7wBOsa7HJIDXsgJKeWNlRDFBYia8P9HdHBR71LOwf/rMZ91EvqsL8vqxE9
18P9lwMATZi4ru9ypWqGBjjg+AnwRuaMR6WY5Jp8DcbWC3in5ec4sfVwGzJ3tduf
wRAVQkYRT7yRx/46l8fIFgtLHTxtk7chQFtEgupf/z9pcOS9heEjdP4pbtrvK0Z7
qV3KmyqSDlS6LQZMU4AiZYZWx98ZgCvcOJuA5R3hkWKd5sml5KV3Ay0izuDPqrPS
NwljUIzlryMTaXheIlQSYmNgfoqBq7pmSHJU+rDBLWt26DvgLtTiTIepo6CCGshF
vwL2aYAaGQNh8gj3J99MSoHkQdKNw0cDNGx7HvAK7Dl0PJD8EvzwPBZRtle4XHlb
I7L+r2S4lCx13BcAkvpYoc7FsjM3L4yJ5bhSR2B7fC354iqf7fRnb2bMuEXbD6Wa
qCcOKxEEoM1eDNHuQ6dFv1iYm1ThZ8ixVYeHT+7Fwc1pNqf8q2g3OIdBgc+N8a5w
EYlBpEnX21bmGJmL0PtgpiqWVrONmE8WvyGd0cubwLF6g0T1IK723fbvqGShCYOL
F55jaqQ5eWxmyQZksZv9Seckvn/gwb3i5hEupGMpzEI/QfqdjRjsB+kT3g1C78Jh
BakapLvxVkWMc6mEHN+VcVNkbQZD193G6zyxC0EW5MN7i1/Szmlcnjqp89V1DNOD
RsB0c5FT7PgcszePFG7cLyBE2Dkn6ym1yyBRBqH356VIVvrjMjt0DOhZotfjKF4k
EEklmg/+dLQ8fjO/O+Fi3E4Lpv+FtZI/EShEgWUbuLyol7Dhekxeg41gyLDpF3nl
zeQyhc/7xefHceu6EooZvcBtqH1TCUGsNzf/8XQhhvdwsTqAz9xcrGlRAxjj/XS2
1q1khNvezTE1i8e2D1qNLnkTGL/TBC2jSp3UBsWMST55qcP4uWeZCKex+TbDwCf9
cvO+aq8eQaGYzzJQjrOkwpmw7196RyVs/fotrzY2dai9S5TciiGly4VUHYNkOrzl
ePAz/1vl88SjgRfz+zjn25fWdh4WeiPlKpcws8q6LMcQjD6Uht1fJSQTHyFvVxVJ
XtZg0iXmKM685y1AVl8r7290hTfTDblD6weK2kmegj+03C8IWKFGBmuQRxXOubEa
maFeYR1UcOJdyVoTUWtGUIkV+RMzxQCMOOEBhSBIGPJeW2FF3Tns8/0g2QCI1F2L
a5MPhuefO0W644q4U4De8mFaq/50sP99+Rj8FCtbwdYeRFuURZpQ/5oh5X6qghra
zEfzsKk64m0J545wBlyQViXPGTkxwU4iqFZ3yfAmwSkygO/MqSsK7tcLZaRZHZca
FcrCwEv4Kl07+xygoljo7pHnKRF+gTeiKqJFY9d+InNWyQPwGwqs8Ndq4G7gadqo
lDmEHhC6epRL4B6cxuKGH7Sf/N1OXDiqbwcs2RVeidB6P5XWJhSDCgUxOhb7Cqw/
3QmaN8bfKgS18q2N2uJ4m0alqnhhP1ww6+g5fvEKVz6OG6I3uQi/hjFvER8C6Rpq
LC1ZbQW5BuS5RP+dY1PatVgTDxNjR25CU9iU7leJ954dLrvVImLTCbDM2Ba1WuTT
d26Ar7H16DoxOM2hT5TueSQdI/MkoQCd9iXtxulsJFJqTaiFPc2ddF5JprkUnTpu
Aar/qwRyOJKij7WN0Gl/iPwwtveSBxztHiwgc3BY6wlC2TA3VY3mDd9NTc97tkRX
oTc/wayW2fx1bEZTvZnyfJmdMg8hztG0lTcrhiWoQ1RKX6MPd7VzjAC9d3pLSASH
L2hqjKCCLK3txU7B54xlwt7ilpum+Yx/u2+tkYSxqjoF3TFfaP5FZO45Nl6v6zHJ
RZ4s0S0gaUQTvAGzvHg8wq5XUzRxezZFn/qsGX7SuP3KmzXXzv0wj3PHjVIJuE7E
BA2OI1ITKZLbpyAv1gFBcvPT2OKWluXvHWfEos8IAWHMeffxOfcauoP4FsjNtGyh
NO9oB9bTY4u3oRiT3cJPMWjx757MjeP09roH0ZvL1bxE8y2+lL6BSjj1hP5WvmmF
iGu8oKN207zo/po4BvPqk3Y9vUWhdACEmRj7gb0iWOIrZm51peEN7eaiBiheBJSR
t/HyRWazht0Q0Z9UXeeZHMahC7liNhb8HK48UzCJhecrmr/gcVkMeZCgM1F19bHo
n30N+INKEGwAxAvw4C9c2lAwSn4F6MowEPLrToI0giZPfUVERnQBtLZqHmYLjNHT
BDHQ9WYADJX28k4rLY3WBz7KE3KHPF+6/yxTrw9B3tLPYO/ApFr+4DDiCpgCuPj+
kqysNmiWaXwpI1BNZL065P4HV8hox//MvrdyXU1iM0RboVClNunRNw8zSZroaw3J
Qv/40NI2ncv/xIGotWQIl3VcaIiBh6Jcf1gP418ItAZlXSkbNZzAtHmfbIKUL5RE
RB0KbgJ0Euq2sDQ0Hf0dRJze2jdP2Em+vgH9lLoUTDNTEC62Cxwwr8nTJrMwYDIB
2+8NNASepQ4CRFpYVjbUE+CpP8/IQnROkA6bMInh6ed48GAwWYJbn1LTjBUSEkzx
7TZF7GcGk5Q73uA/pKnMS7mjszPBUPhsCCcNvSKjjSo78B8ngNxbetNqNuPvGvC6
Lyu8nM9m1mQoLTq3Db+RxnjnCyeKE4LO6LfS6nANlYK7xASuoEL7nOo+XwiqEV7Q
IWDa/uN1cFFca6aFQoz0c/L8ygkAU1L+Kiyxm/T2YjDRND6WV/fdxWxvSV3tf3Ys
38F4DU4W4pmf+IICJVMJ0mdhOfA1DIW/zlRbPvLoqqkdLyH/epXI0Dkbb48Qtm9P
0/O63nVzvIczPAL3dtT8OlQLJ8WKPlqSRcalt4ly3X1BD5wxYD3FJgVyxo77AsFn
jpEDKmAPqN2ns7bzvgsN8t42CqcVrxWS7Ypah7ohrfKJ5hhxe8R4AmDU3qiYLvGU
MsQKbNEWvaZpQZE8RFqnfiG4mnHtRsBldIV8g1M18SqVSOZWfarE2LxToyJj3f9K
BqdLD+bgulPw9lMeijPvNk9i6/CCOFUUl7sprjGI29yIj5iuEQ8/lMC5QHFoO6X/
w49D9bSjJlryUCuy2Z9z1WLzgM4bnIFyF07VluyV/CubND9ga6UiC75bnQalLBHn
/JgcJRHSTIg26pTh8jg2b5m7HRUoZuyWh/IJ2sygu/iz49l80r3+IRylJuj6N1Sw
czW2HmnySUe7ScHo7R2DWmnhPUDJ7Um3b2Qn3r7oAZngjuX3aRYstAkHEfGEuSGg
APt6XyJ+M/Nc4zJzVk2Xcf3wFIp5Wshz9b3HCrY8AWe+ikO7ffC4keUw+N96vKFi
aKpPM6X2oaJjJ+M9YlEK+f4Cb5IV3nwr8hIxQ3LGNgY//5jloiybK00tfVgT4BYo
iLsQ+GP5Xkm7v4ygWv2Lx1HA0e+EX99zXkjrU3wYlJAh9i4Xynx0Gxz8R7hzURMo
pkUvIcT7HPE19mW/YSW5Q0W7rosSwfyUl0qtUYP5XI6H/iVNjseZ/FKAfPOqQ6C3
sCx4ir4N9i3JOzfxhzZrHHnPdc//iiDAik95r9ks8V6pbztrlYknHI3VduPyuPn3
3z0XBk2zquVC41m7pdUnpC5bhIETgBx/XqSrbNSTLOd1XKJWh3onnex8YnVU7gfq
9ZNT6JxZmlhphb/vaAP8IoV7l9wJdbUBoq61HNm2P5GidIaqy68qByw5fO1xpLoN
sFKhSJyk+JDXlE9PG4EUiOqNY9rd8jNsE9mZsgCS7CHv2iGszsFIuK2kofXAvn8K
FOp7KlY3mC8ixarab4jCkoTAD5fVHk3ePkZ4hjd34RPhH7lh1GR4dXK//xNKomCt
wfT8veL/OlJVby8eZ2BuRHeY0CaWTaoxxx86QjpK3HbXF+hxOaERGT6uhfDOTQzE
T7FZeMwYqI7Bk+wEZSUP//OhgaQ5JWmpO4dlxLVOKFUkya6fuw3Yv2WL/Z96keTG
fyYeIGxa8JXCGoj2lotqMvRSxqTHhX7ooHmzJhIKbqQEu6EWyG3aW8FhhPTG3XQD
O2TZ1HL/U1Dua57ZouS8H2jVG2Q+FXxDJPepLQxMjJN9dmawbfhxDQ5eqiwMntq3
D31gr1S1j91X0fDmvQVejd2q747gzPxUdbnaXFDIzx5b5q1DRmD1nMzLeQT/5xqW
Tt21hDpPnI9AR5Pe0wJzbJlwgPGXO8k6QpJPVlz8yHJ4QAjGIshcGxIX4aSsx01J
UI6nqlcDPP8hFC3ltmmY/Q78YMO/rv+IORb+WcZbAcH4hWh6MVevNMywYHENb/Ov
ecwlpMhadCXKaDAmc02e07l/otUNz9JAKLu9/FI/E6O2Etd0xyopo+EWYWfvOeJV
T83wLwSr4VXXcACCgrLqimiF+zwQuk0wXTWfpwHk7YZ7hmR1ZM1zmT/uYQwg4QN1
PFVmbAkJCm3qsEkAkstdyNrte2dAWyuYYAUDMutZCe2BDdnerT06x697CqBjJUk0
F1aEHcJ8LfYoaCDziLmA2ENQxvmd81ce+ArX3KfdYU1OcXVNR1xbXUuVf3vhaDrD
K5xl4xWh/Qf1qZGZMLiQysxcW2TYUdyyOxAxe0UD1dMA2uHKlcmZyzXNIOWSSrZ6
NWUOTf2Ra4Dt5HAeS1uA1IqRSnuJvTdYEyhLUP7LTCTtpG5rpDrzDZR7QBvB3DCe
IDhbtCdLSe40SFFmgkt/WqTPRMPdhxobBLf3AnIyjcKRZxOV3KsvoZzKnUOpJr3t
vNKO3O9cHYqjAb13c5FuptEGohKzYwm1WjMngICXmagjIrUfXTrZaiK3MqCkNE2z
J4+4b+ANQrdR+QLtkgQShrKCZJtj01S+PN5u2NvmQaJYkdU/GQxkdD5+kQmcqv7D
0smwJkSvlx3HyV+iht+ML7AolYfgKSsISaqMu2sshLo0m4LKRdERBgGQhqPiHIjn
yH1FbZiDSQZLUjqJayyZ9NpW47QpBzVwFk9CN9ekTghfA21kUxOXH20b9j/Yk6tz
e9fcnjHsy07OTe3vgwGo5XaxFgKmOGLzA4DYeIGmcxDv2gToAoCiFXZKRkIX2sbf
F1BU2UXf5IijJYnL14EtgZdpMI3CzEnShaQV6BSZO8G7REJOnCbj+IjpbrSd5yRG
IbP4aXQ1jrLnPjniNST7LdWC55kebcAW1hxOf1ZoneUgs76eQ4+UEHNCtz87ipJn
sN+GQ7JobcBkyiQ/18Y6HTR6PBbNH8FGKQmRYB1xLtFmHIUHwi4CTWFPIoLUA6sf
Qmni97fKY6sZYXk6V6z1yTFVXxLQsIrnmmLD7rhCqeC9bUV8J5dXDKw/NGWm8aut
3nVlBIy3UKYUANjkUutz0BytfdHtj9SmBsCAIQLSjO4cjcrCzPVTBQ/EUNIYMHoJ
ukCchJK0lACvuAy36FzDYaM5RCqgyZC52aDkjsF/jKc2kDINrqOHQqkiNxoL+OK0
J7kE25oNL6FUgKonv1aY/rx7HZZdTbVO603jRkdm2D/f8n8A2hoBO7omuTNx/NVZ
KtoTMRaTdCrtCcm9syYL7Dh9kgg+iWscOqt7n5Gtyj+7BppJEH12m50xEGhMVu9c
/02al2uEFmsbXZTM4y/DQg/Ls/A6OstWXsyfit1TYJQb6MvMAu+Kdsxlh54orPAD
s9SMsv1oi5WvLXPsG1CcQK0bkDDJZfF2G2yNRTHvq9B+9+KWIXZiSVvQAgsCwZQ8
cGiJFX94yzGVFqq/vUcnqnyEhxODuqiDAKnaXHDWgo2/iFhQ58YW/yZr480ou0x6
eiKCEx7+Hs7WMcOH/SSqCD0WcdJ1m6dUqludjsEMsk21Pdu3c1r+RujLDk1T73fD
sCMg1ndP5oMRD7JI5LzH+8DeErlCuTjDErUpBdoOw+QpoucWTAXObTbCMVnTf381
oBeR6qOpX/bX7b75s5mtK3pTt5wj8TMbFkr4WDOpSKj2j9mbPkkmU2uRcOjxeXaf
FOPP5jZzOtWtwWg/9uiq2rtl+QNaMML5xfDMAd32uDTDTrtOzPaBrKL78U4vofng
bu6RjA0wsBC6xXPaILgft0grGlmNmd0RYh5kdzkF82Ff/JNh+GuZNzTvNH0lg3S0
mJlWMxriIanvUuVF6bmie/fNZaiwcehKn/lc4eDWii/wy5Jt8JJc4aqmFGxXVDCc
+PvTg65TsXxZhs7B1lFUHnHT9pAwizjYU9XKbJDUGFGqHY5bi7485crJC2kfvwMt
qkk32HQTIQthMjhCgBufULVWsqP0d7sZ2XDRBOM/jG8FidtcW4ZJZ1O4cBwidxpD
heYciohTePZfNqJu/XH79JNs+Vl0Kak6eRrHVe7Leo10CFtSuqs10RdMWmOoheld
90AktxCyzyQKa96cQPmsQMKV8kcKPbBeO1KO898siIK1JRkGZQCrGcK3E2JnRZs+
IfwOTu7M2AW082uUNGvc2QvxDUjLarHXOmHMD0ll2z06Z/lrJtVg1Ss63J4lEcxK
BEyjzpxjvYTg3LiMgr5sh9uveD3NwAoGHOSqf8ACOr79na6fvt7LzOsK691nnHXg
CG+paDUq7TrXjmcLA0MAAYuQ2tjB77gknyLRsW+mFiMXj88nkmKL2Tc5+lZ5gqKr
gMclwOkq5TIMs9KopZfHC4s9jvWvtz3RSsgHtQV43oLPWPQUpFGxaopeRohJ0Whu
IzNPnD4fqle6ewedhicNnqeYUieRgbeu9/D2AL8f3ira5i/7K/Q/3LESLdQCMHWO
g6Tcx0f9J8uZ5HS6QLaaOCOAbYZo4vAZHjonVjqEkMP0Nj4wklkSFyC2AVhrE4yb
1wz1JHG6aW61vLr9Led1eyXbZXa72IbIAhZ34uO/GmWnjUbBm7NdgSjFnOkJlgx1
12fgy68FMMb6xZPGO0DHurCxti7D+UuABvg7vMw8kfxWvtGZqimsEYi10kDEH6Td
HiK5Pj3OXA98rfMUQ76ve3/H5vQdk31GjPgMuQfUVFF50g9cwH1iZQlBO3NE9Nk7
Chrl69VooVf0OhNeMHnLDa815nfBLxYZlrcvdKPUq3L+MRxa3FQM7yjq/OZbtPQx
t3c6W4XybV91xxfu5u3mho7sb2UNqU/64rXSgpH5Z4uRV2HXAMA2lvPi4IiT8af2
gyqC5tYGV+z7nyjOv9CtNNdpzXQZTjLnjFmSX5CqsY3RL8eQ5nz7OGcRQaPEIVZ7
Z4PE63T5t76shP50o+wVXnMA3RK05/lwCY+5LbSofekhgrVpYm3ZAnJRBpV13rjS
0xSEPCjS6qdH7w7eT/AlwEtHezpSkk7V1KKXkolquJFsEYb8MNpR4Oa0sTOW7ftC
YeB7E7As6Ql71bPC4W+auEYH8PcG96/E/w7KqH8WjjovwLkLkolrXPMkYTOm6iAw
sSAYYd5+tNWn3rvVXZ3o6yfxNpIAw3fnc6TdFdVVvTX//nM4SRo1SATjHATXqgOa
v+fjt3HR7Ir3DmyZUB/T9+azVQxCiMYte8kbwTioMxPu73f1pGgpYbfMZNufJnPI
Yj2CyaE2y4vCd6Vj6uYkai2N6vI2jB6ZStSN2K0ykXikgshoDGRWHzicZ8Yur7Ey
LG1NcOkjIu4MPQTy6reUfxxLSMvifrWPhZV53bZ4rsS0zYccVwT/5LAN6tukI9xj
qDna4VBdHlqXl2oz/uBlMZfgEnGDicRaOUhZYXL+dQIUJkplCAMwRMBhIN/j/+S1
OBQ2v8d39NmZ635llPUwHCQxMqKsgWQoissq2LKDBAfSfNo5VM7xK72PMwrh/clX
/cGnM6Zk2s9Rv9vy8CLrqwaJlCSJVw4rH1Hq5+n9rZ6dp7oJHrKBi5oMv5CAXj4x
coKFSr1/pWIgWe9VUr9gZtJSgahoDIemOCn2coYKP2JnJD70MF/iaWkYyRpD8Mg+
uAFJ9JHOez1GXFGzWGvid7ewKurmhdiFZ9c3atHiP2cQSAj0Wtz3ZM+JcEM9PYZM
8A2T1Ubpv8frPoWY5vuDRxIpAYgxfGn2RBwjm4zrMd4Fnwsz9udTA5/VlpKBCcDv
rIj+FQX3UzdhHcUetmYx+KN2XRJddpSkgAhgY3Nj3RImOh7X5wApRmV1z8xi/CxG
499Ref3x1Ck/GzPUAptKHLtd+tmsdNnldVCYEid/I1aYdpeet73owqu71/q1EyEy
DvV11m5neNGAGvVqtAjqXJv4Dqbnpl0FHMG7sSAAttFCmKlqnTNFgiRpRldPbo7b
8VgidUrLdPMcecNLcpR7MVgVvHf8uieNFemHgjX3RGtxxMUYfE9BwSnnvUZ1i0fj
NoL6TWpW9EhCJ7mivCp8iskgqDm/faZ62XKGFXU8FmYd11/yujPvEqbVYKq0RYDT
AizzEbxsmV/4qBNfSD4qSx+iqJN+oGwVfwbnjAifWcEpWGqCCliMA0lR+dEywf3B
eH7VB0rHDOg5y0VsaP9eQGPA9vfgKDWMVJ0EhTIPcux/m6HKPdWsa6+FCSFacBku
kGq90jWG6uVYVytfbexKrCZkjV8i/clralWdn1wc5naoI54GAtOeaTPsGNKkalu+
afm2t8PYk8L4HUa8hi0Q0OkojAH99OKOYfwRpor+0UTxH2FVueqpIuRZi1BNgjQN
7CZ3ulTtw4BITnFt7TD9nDtx/8vWA/t1odd4Gr19BbLwYOxb40EXhRJokIRlF8wH
jxAzzWnsGn41tdc5vZiG/Try4wY0u0LcdW4SyTnPugd4bA9Lwd0gHsOOpiw6dbqv
i00ehAZ/n8duFOMQpDnAg7pD9A2rQfEjtovVJJvcJIRRq1IMacbcZaMzm67bdwIQ
afbfcV7Czw0wRJtEAarc4rLCbzvB8kP7tRxuzrTsuWphvFhk/eeZ+2UwOnUZBlC2
7Ifv8054rpD+ZHfTqCZ8j2CgNxkfCckM1UA5/jsGNISbWaHjojXmDsRmANVSrCSs
3/el7gnluYnl2P6xP21o+KOrVxGa3bx9OCHXmjTg2264BqV4l7dF+d4z7KJ6qdLN
c3XdO9h2TS7uA1iXke6QWH9cO+WW3G7vt11HbdZQUxDLNw94pc3YLauREptmX6zX
mcUp2sJ5NzjAciI1s9fsq/61O+w0FTeLBWFkzd/xw1ZN3MDtaNsWyTtDClRBgX4w
O11Kwky8GwLc/Y5hYgT5JsAs0eHAxlljDcp1wu45f+45LLm0iVGfD+nVY3j0BNCF
H8hvS7Rmz1qi84jH9Zh+2IZa8TA4VISPwj/uHcGpx5RjMua1NJ5wh1Rw53FIwgOz
qUBwCHlT1KJ4WaLu77s2BY5coxBQ1QLe7MFpzh3l6m9UkBqZTuPlRMEPaenyYhXm
IbIaSTx4mVeY0OTfK8+bS9LVsK1P8h89vMDA+u/tJEFbx7EFugnOI3w9YWB41VYi
DdgfvUd5SBIbSr4nEfRMQlQxI7+3oyPbkIyGwZOrdODxwmsNvJ6Y5cXXBIllx3Gb
Fh+sDBWI5iEbm4Zc/NCaVHu0bHGVAMY0GX3XJgZB55vdZNvdNZmOyjpUg004dLjP
dJGcP/hkArN6ApFko6Z671rcAHRFQUbH6Y6FihSDzzaouYUn6nnryHtObksO++9N
hQdxhlq5SYm8xqRgO8uchOkskGtUu/NT2glzCCU8wxYYbqRUMNQb6nG5wpuvLdY6
Jy5DMZFH5L8RNGM2A59RJQ5CcrwLf4mG8SP2Tf6qOTPxnVZkdwnH44z2+e3OIguT
rzSJSe3xl2iAbmZNaOp1n9ABz/0EoP5nbKbj9bQS7YZnP0bXwBfQ7fr5mQ3rHGyk
50UpOZ+A6fIBroIdVBl1DoeiqyZjg8JrvcZbf3HifT6t+Cpx9BmNa9D8y/vp/Xrl
x4L8Ks6b8Wc/1zhiVb7/FggeHhOIs9qontj4/DKzhYJFHWfURTMora9i/28OZ4kA
mLOwMJhNMHByXVPgBnQPilMj1kswApI5XYJ3v5gzg28nYZvkNM4q1jzUXoCf4L82
/+SjQE3qOSIVgmB4kGVgj/NMknzHDaeCQMebXpjF4h3LSyL4ZmEzvgYD1E9SxEgt
GT29cFoh+SL9tU7V5rPvQgMUWd/uJAnfd34uGHMVkcYe+t3A7UxPs7AqhZ3DQCjU
HEmYc9FCGUqlqZK07pChWBTt2j6Zb1xpyPV2GDA/rbFDlfY280cSPHCpFlrJ2MEs
Xxd6Ru/w0+QwRXz3/lZnZlcdH+d/999DNMV0WcOVyeQaoya6v/SHVggVd7Vw8GUk
kMXcXrKhzYcblmvTXdJNDDr0Jbyoxsopcuumsnm7tNU8IiIhBiI83R/qrXngqKIz
Rl5/If55kehzFIa3qWEqsRz0s//yMMIFrYzSTkjke92GSyEOcpvz+CbfdhAu0kOr
P74O1+/Oqh8auVlWxIFbztZhCYLu2HeDB68+lr36RyMGEqgVpBS2pbtAmD+6ROe5
7g91M1UAaYfqimokbG3nC8VuFlXlR0xvizaIZBENqOt7ogzBWqUBdJU1ZwFe0Yhj
qLTANbJItSbcmqmbTSFOI9ohwc8BhfITC5u3J53o63T0BEkwW+MyTZmMwulQOS4j
n21NPK0+8Lwykh+FqJDbxqGBY7OGPHStLhaJwyoxCyJ4FaqOnN58V02AES9Pps2K
/GdB2FrcZAwJ9ME3qpKduRRNHzDSRqQZDbphmkZXUHUzmuZT8MjxXHIQlFKm2edk
rANxbUCrYup6Lj+jsFpRM7HoY3XS+irZ6HU6pjTXE4t0ysu6RQ6P8UKCF400ClGK
xpFjT/u8+B7LmKeWIOEgV/m2QLJtKsQdErTHQ+pJXhGCbuMeBCqizj04+g8aXctn
15GcJEkS9ipSJJLmcz76RCpsSHNzxjadKLCaeCWKzUrjYmEIHMxBn3X9ex7mY6xf
YvFE2b4b9eD9a9XJuUPDSyfrWehslZpPSg7dGnwNJvPV3lUlgYdciC1mLqlWi4Fp
XrSVjF4porhOJonJaDgWkA0mwa20Jzk5OIe9gJnY/GS3ZUYrdOlsVZ9Xw9TrSQDF
VxekZxACb/VwiTg0zgbeNMGl9BerEDllIDDcFjQRKv6grsCmr2Cijhq0S8saHrxa
brUX3YnMeM1veeX2+FJZVl+5a42r4ieaR9NqOZo0irVhWswX1imX9D4qvfGactPL
J3w8c188AsbhqkAFPa486/iygpWWOqyOWdD6zyxZRpBb26olQ59yph2b+nCiIn/g
94aE/ejpMHCEBei3n7Q+A8R4C5McqlA+kJAvkWvWof3yIadkCfsF2EXbEBEtubg8
lLA0esvmcO8BYFvqVCqRSED6+6Q+UPlJ1JXlsI9Blwyj3u4e6ecEGStSwgAaPz20
Ehee8NarVr8ygAB8nI8ndZYCnG2ffkhFUxZUCC1x86mTRuuafla4gLKKixhENfiA
ls0GO+3WBf8zp/9p1EOHgyWhTQ+h16pzg0EUAwd3VQkI05WeVslPwGV1K71/kyZ5
2T4s9amMXw3YbM6mEZCvnFmnGa31yNDqWimzo+HrihUty5u9jMRJhe5n4aBfoQje
i4vyca8KDdeqD3CCYfh5DyaJT4/eGX1YEsQT0IruACVJwrdNuikHeQviTlHQRKh9
0ohvrzUQAt3yO4Dza0F6A5KGv+zTLqEvL406m7/Ru36iD9wA4LZFuyBgBOJRLiN5
A0e82hXwqQAe5ZBk2bx5deTDlhwe1zvtKEsjEG+gnCgj8wnTnRxDBIQf1DMJRuLQ
ykArANv61XiZUE3J9J9R5ugubZKWcSlKspWACh00AposYXYdwho4EYIaXrqrLS62
J4KVJGApKLGm96xl89VD3XavUWw0q6SPCsIrn8Qarn4GORBlQGEknoRroGaZX5XW
7pH9CAXO5hYzBI2zVhOvCCwiRBRkjoKUwPVVQKYH4CFeweInElYEi2BVTqFnJADi
A4F8o70l2CHNE3BFuXjh6zqVT9dOhaxzrvfksUfqeuedn3T4K1oD7A4skw76VADe
SjGg+NGhXPaZIjvWPneSt9DUK6qURx5FgUFS0OW6qdZQHp20Nzi+Nvd5U5tgdXYa
U2BRAM4aOitCwoKsQiiKaTFiDHTZvRI6d3xz6SzRPUBD38kRp6O7ijqMf0SDidC6
gFS61CXY7CxZxCgSe/oynC1xqEmItG3hNtR3yaSZjNp5IgSbsBOHA4bnm2f/ElJl
hkUaipZJTtm4agfMv3iyZRaKC1cJH5lnSdj/3rQ2z7Y47jFICYD5RPI7te0YLg6e
05EcsEltZzGFYTYYlOBwkAWE+BGCWJio9QhbslpAuYQmNlPc5STPxlydYdr5QQLp
8uKKTz3E1C47+xSSQ1PjFtr7QIPD161yRlqrOVUeng4PWg1rcpCw7lUaLDRRBGcL
isn5FV4olDOjjy5Lkh9ckfjZ/BFiAQhRIz1t+ZLjZGjRGibf0HCQRtGxFdu/robO
egdlpUSd993QfBFxvi71nYSJIdt/eBcGLa6GvwaEBquzvJ3Od8AfnwUEuxoYhyZE
ieFmUE1kXjwB3T/azVf+lp9hEWp+qzVtcZgVU2/LPjWZ1GdGeYojwM5qfJhzsNqr
1h4uQEKhtO2GsChqhf40aOoOjmDHUMBSBduJDxH1CxZo2Lx1eHoZr+KJmo4oMOaA
KLEjYHnWefPX5XuSKbdQJc3zgbM5lVwp1Un83MCftHGvxeHNwQr4w9KNa/JH8DQl
I0Nwwup9yMhb1qY1Dg3kmmsD+T3NAjsrgpELBH3ZkLfIP2s494RmSFXYCobfRY1o
WTyDWq30Mme51Xi1AwBhF5NbiWiTvrVevBp0BUbwPjmW159YFAfQ2eA/SKla/I4V
F/cPzbME34qITt6Onlc2OILpBd/gYbLwIQXYLkTMrWyvTWfMAF6mJzZr9UMvIPEf
s84C9oD4I+ry7f4aNEmrVI7ZcabCRV6fUahwxZyIuqEjFlK5SV7V+qVZh3rQPmw+
tSrPyQQugU54ged0FzMBwbTldfqlwWzMQ2It7ZXFcTjdDBB5BZO6U5cdqSgoMvBL
ECq4O8aq5dJefxDZD6wihTLQ/hPLxMB17l4owjTAYLa6MrnO/FRP2y+KQhr6Cxkr
sfU1wwwLbsOgcQqWzYcnopoobldUpshvKIk0B/RnT2B3TH9GT1hHETkXq5JIk9MO
8lZckW2C8QOFDlqmZdRX/+IDBUIdHvNc8uAjcKtA+KfAktv48lJuOJkBN2z7uRR6
OBpVrl2LRGUCEstt5HlC0WfyJepgWDznG1WvVk082uGtN8rWpQaWqAaW154/Z5Cc
+9BZyqwNuGnvr50T0jneXaMyJl3XuPAXYND4niycDYbzcdlf0OPrRYfTd9Cix0u2
+fKlIK8WoqfFh90Hhd1XCVOeBLKLsAD3MwuowbK2N9tbHd4R1RMpqdkjaI46C2KA
iAtZAnlchqSaz2RU9hW5pL8lhIXDD/coMug7B/+uOwDUHeNa6M2+R0oC7YzHwF0G
ZWFUg6xk3Br8ezCPqvpIXzCHH8J0HCg1id3HYof3kzJp+BnVbayd81fz55LGEst9
NfOPCyPvowOrJMRkcZK1pXWHOzoLsXdjIjcQzxBTySlOlEZOGLlDKnd62wXIJWCc
g+Ds5US4kW1VlIcnAjBjPUXF7HLpEKIflTngG6457E7hL+wXfQblw65hH/crBP3T
Yikxq7bjxSBgc9rjiPILWKBr1wbEkEHXiXe/1sSqGbtL1mEScYYgYzhgoe+VTMsE
tJWpHT+ynSODrqPIOLaEVVR3QawIHJll2GoUexaitbNAGXfMmu63LCdg2RfwpQE0
X2Jc+ci91CL0VkL8jIX7ZsmXFVvxaWbpLaVO08mhnVMZjY8Hl0TmzYOzh7h6hRe4
gqoEFOTkwPbncE2gCEqbaoIhHfp14Ad5nxmhn2abdlPt3ONnwVYoNIY4fUZIgFRU
r+ZGxL+6Uk6Jbsxjs7ro5aZW25xYRZu4HCLbNexkZl3rd1xhn5usUKFaSTbQT+PF
o8J6O2y+g7meQCVgjtfMp52skT9UrNjqo1NSAOwTCxX55a4tK1uKO77tT88Dqxpn
wkjgml322nmKiD7xITFXG6Frywu6WezIILM4cju6MN43DmsWJkKg9xwYiy1OdTOh
3/P9q0w/v5wFS6+dQGoaNwCyDpzQXbzS2xBSi0xdBnjcXXu8t8l6F2K5m1rdRmFD
YhgMlRggEYmY33KMGsnOlf9anMoXqVfCfCNb1DeZolNygx1zJrt49EigUQ3HEgYI
LAKXT9wtYBFye/+onsjjN6B9D73YVMlQw6PsJyBI5wBOhY6q93PFMhK3DCWKpA0n
fz4roi9I+Q+ho59vtiK/FT6Eldh1xPtGIyOxKRjabEPeIUR9HO5OYPNutxhxIO//
VwDGv6I69vMRPRtNKcx8Z76fwpnklYP7ZwKNW+2WFbQK5EMEHjsfhF90HJ2nwHpB
tojRKEf7sqjdye6VSkP8weIYpQC9DlJk4JctiVKrMmSrpeuca1W4VPBnU4EHLqjT
nZiYhaoqX/Cc0SRXDxZMbznRCDYz3JHCf2KGSrBGXCk4UzlRuhm6qZcmW22hDlm8
BIXOTy0odgbbaAq0dOr6JXfz1PPDaebIpHVRVcIV695cTAu0tW2QQN0EN5fHT1H2
ynhVD4TNnZe+H/yvu8E9LdOg1ogRWECEdXUtm/Usnw72kGp5GOVDnrZRD9VigVrF
OcZBVWrVyAISor93AtqA5hPWq0Xf+BVt0PL9+EPH0Dswc+egm01K4pxLTLyV2PwA
VjivAqdyxm/yZYxDlPZiKwILJq0GCJL0b4axF/GP/YK32VrWd75ZN9m0tynHo1hM
rczPITNFQLa+YZPNIvBiFSu41FtFBGKxEnOoyQWARnZkIIKyLpl8Z5shTwBtShVs
iS/bv2/9az9M5ZTQzvUFvWEpgFS/5xUrHdbvrJ1RGa0mF/lyVWYUXmyPHltXG78M
h6xKo6iNiJnQ0x0xlkU7zJts9lT//ym8xG5rDHeG/5k7GBxOcrMYFQFPbLNxoMFU
4a883KiUgZB/NVwRukJRGrawagelDMm/NNXl4TAwh9IgbXB4K2QuhX0ugO1uLtmV
q8i9q+q2hOy5uWJFGo8S4eu94Xtdv1tbeErGnM/qYYRHCJpXR5fOzy2f2HWBr/Ea
IDQtwZ+tdZ3VDbpbvHKD1O0CMwURnHFGia9bdPLK5CugO8E94y4EGuKIIjk00Vhn
3xpIQr8PmZ57M6NlvvyGaLhYE4XR+2IXFtHpyGtP1Ss0VpaSH3JCb2QRn6JjMZbU
SSFHNXb5slhvQc/84x2Ev0lH0xvNalY52bQBKQ6isRY5SumdldO8O1ByUCsTAlcz
yuU6uKW2nWX7iDkmZI1kDFXK6F2QsITTHftV5XwpskjFneDE7YSZvO/PvwkyHL9P
6hCM6ghV4tkJl7PcE58K/035+24qlwyM933M2Iuz/cPpPUmqc0DN2E7HVeoYsPYi
vzpoxhn0x4CMZtgzA/7bbNC5BVmd0U/oSYf/dN8aiZYRthLYfdxGX9lxBhTcnuIh
Ft7brNmL/aE50Y6r6BkaqcWW3GN/SDZ4+6As8i9hH9pvQVcVKqEOTp2sh+s5b4iJ
GBeqHJaApstK6fif8sZSHxIhz6hXNqJ6HOBA68whqJIGp9RHKx+alk3McDbAwDps
6yqjrPeXFPQhZ/OrDxEpqkopZ/viYc5ESUz3Bfole8QGgVgeeRlJI+Ek45BcH077
qF+3A3m0bVvE3mATj/kWd2KXhZ5m9dDDvsS8Ds5RchL9QkC3HB0THU6r4mFFrlXG
QO4+Y6yXYmDtgnoyBxe0AVfI+p39AmwmRKj9GZb/9wtAdjCE6+mI9fZ8sixw3BBM
N/ETxkEFaJgqZVzhT6JskyL19MrZQOOB2B1ARduX/mxSZTDELyS/mLqDYnol1Bke
PA6phIY9qHkiJIN7SHPBOaGYCMDpQSgiJ/I9Xnxvc5Bwsz9KKgYDbyae0IDsYa4U
nc0E9xEic5BoS5DATNa9tTGzpC0wab58595UM9dYt+NCoAIZgYKyagrn2ImaZLjp
ZxH848lKHpO/dQEIiFJHH9qKRK/GaOezyb6PWAopeBb0gZPUnqBmJ2jVzlbeA1DC
1AfKK6aVa1jjC67ENRxqf15bpStogOFR11FkKFXbkXuoEMEXceb4sM2MSsnoVYBc
/6G2jGX5nfCuPF7em2Q2pe0Dy7pRrSghtViCRHntSujAQ9t9bRApUNeOk7g4FjNd
QjcY9mHQ+3kF/V8i6UrpCtdnuihM83y9VrDp9DRUnXzPbAeAdpKhGyenxmXoYSu9
nIpH7wc21wzrqqqGJv+kzE81a1ELPCMUeKDzqtZYpSkI566UXuHrq9wsrHSzFoKi
nk3e8CFBoYPnfo1GI21llq7Bp8PU3DPZNHMnvW1Pele3XjU7KEU1/C4kyFKbPbAd
Ya88MnMFSbhCeLD/A8If6ioPKzWcDsvtVOKt8zzcxliJMO0tdQQ53kcyc8c3dktr
5Do5KTQUONmOVoC1zrmjCi98QM/gDm1gN/vVPscOHo8IGELCw+iVcIZD3GAk6ViG
7fmkzeUa5mX2f7osfDtSqYMjy8gpcvF523xfnY6gE5QLqBzmajVr2RNmEDrCgAFv
qPInzDiKrxXdxRUrCLbuUfwqc5jbzK3wmhUNeWVr3B94uN+bI2wxDDqttSp2F+3k
AyfpzMCWOOm6+Nf0W/Hsfq1bDpSmOedhsCyoVLGbpffKzTIQiGVBI9Gi5S2KwFPt
hxuuOSwvuaOKQUslzI1tdcoAD8r4yqr8kNvuFiMcS+1E2M0+aKQdN8SpV/ysvE3l
0Q2eUViAYZ9NgNa5G8T0QcUZK7ykbISSajDaoysMD8aD9gRNxBuzY2/xI9JU5M+8
SVBkcgGjTeH5Ybw2KaWT3iZIsPlFcR7wKTEvwAz859wheMvV7NPb6JaiK5C4rA61
Fj5I+kZ0hY64CgSnA5s0pW/UI4+uQfbDm9wfiEUmxTpFzScMlKTcO2dUjzrbpe76
nB5Y9MVfgevUub9LjgFlN1ZR2USkBxA9E2cNkNcQ6l2GB4j3lJBC625hAAzjGmcC
h0pcK0KIdmjQYW850Y4hQH2B6mneGlv4vGdQSGgiJ01i36m+po+zIlRUSBcz92YT
Z3kY6qIqkGvvtYbiQoI+K3LvoCsfJZSk5g64mHmBQmgyTcMql08pzj9KdTBmEZTL
AhelUDG6pE/7IWqV5WI/iY7jrqYu0P/aGmeUSat3RLkjbW1BPRH0sTMp7u+ihHgd
NRZ5nFf8kDfPF8ZYbzidupYStuB/PNPM5qiaDaLTp+Qcp5jsP8aUXxM+1fvIOKrl
blUA0+KrrVO7l/y4XmTbNcOXB2JZ9DUIePmonffoXHo6f116QcQM7ne8lQmhEzfj
Hicyj7f8CBZXl2mI/NDm9MKG4NhHbTgxu68tETokmVBPC3PxFlyPdu3IYVwA+aNn
EgxrEvjFxP7s+5ZCEAaDq+f8JKHtmGSbeGsOk2+Ypqcj4ThFMTwsJQfltDZEi2zf
aHFkPKZu+eQCU+gpkCjIjgUrN8c9PnGB2OXTkHfQFw1lNSLDeevyBf0ENBA2mJaZ
+4WpPOnG4uWrgUZeQOVOZMBFkkdr6I4te78lZ6wQWnmL+tkMUZUs6QCKK17dt1V+
SY79Q4KU6oL+TopXtsduUULqRcexdpklmqQUh8uuIiqdIFURN+ivs6gqPSAnV3jw
R/k5FUgD5v5aGJc+Oxn+WgXmQq9T8hDcLuX5bEsm8cKf8DE0mvDgyzNwXGWUuYkt
5ovnATla885PZTDWFsB2phnk1O30NbiGl+RUH9wxkwGwSTpWTwJAKv+zkCsonwhc
OQYnIevSOApWeeYMH3gnsE+kkIE30dOHctqSSNlnTUpbfJ+I2PikF5/Onf/HhTVC
4lwnVV3Rb8dfCvmNOjo68PZeULGfUGuEFNvdoc+kfDc3nK0CQcGqXUQA0RN/nqf4
f5pjbkhpD0tB/DklL3XJN3p6sR4whjp0FOryyFRYn5AADRHLF/Pf7HT6Eo0Tg/Dm
6X34OBoH922RZOfnRiu8f1C/lkceS6ANB6lCahzPaAGcTM/gopqfBhNvrl48sMrU
Un/dpfZbDXM0+0r91pfV6amEYgctH40EoKzDAlgWow75X11RXYkJlI4VN6tryNxP
5n7m6Alzk/zrWYbmXmskscWOGL3BWM5anLFkwRE8zVChXgydBQhdsAuWA7rpXUUn
Eda/4cKkvqrJ3jJRI2qipS2GFCahciUCMFJV4BLStU1u6/6OV1P8VsTZqKR1EJIU
G2oJj1PGkYSGQsaB2UfEWAEVpoJCOlVN4tfpHwAKGbqGoDqAhIA9EtAw35CRoAyq
HND6c3w+YD0gaWD0L4VnFeR3Oz30yMl9CFaW3KTB0UfCa/hER2AIwLGQrBusF3Eh
YNS9tCUhJxtHkcwjBvZq4ZGv//NECMCqqCEvP1YsP57Mo1ViMhBtcs8aitLFiwEv
za10RIg4Kk66H4DQGHgfvecUoJMSZsf3QNUUgercRqTiHTo+rUiv0I+2HrnfkfXm
+3v+NIOF/UsaG7ZBEgzjPEKhSdU6WDfs9JdBzJPBUIZFZQ5Wb+hwGdJXHHObw/h2
5dQ5uO4wVGbRZyRXtTGGoiv1LrNp9JIRKUwctZljyOSeHmfFLOe1sUHSuGcfcoZb
4XhLdHwLnlPcZrhEi59TdqO2vfuACCNCBLKMmKAPxiV4tHYaciW0zCQ654uiDF4D
fh6nHFnCANRY0AFnDP4y+irZJucsaOMLsbcOp1Z7XUTSzokVvfwZ1WFQZ1OFW/Rr
B8Iys+HKolFzan53MsiaxMp68TZRnQWD2073h2wrJIc0K8hoOGQ0kBkHadkH375E
LByxhciDl+Hnz4ezy3MYyErzNbzHiCuLQmEUE/KYzb25ed47hiBprPL5vBRUx1s9
/9w11hjPWYLyYXq+PuaWDAQR+3tkrVecEnWlDqVQnSDROifhbEumwW7aI1VTQsqo
DlJGhaEnilb7Q5VQT3+1QBA7WH8uPREEm20r2XOVQEORAsctrJIQV+A+PmVugVJV
9LuhjP2JUU40v+xdQbu9r+2qk0OQ4y0wnXZeeg4ROa9B5PCq31lZ412z3eRp9wEX
rqkLBxDKAWg7/Vgr1eT20NhtLlT7pSZrXD2CJ4UE4DAyDPvzEu/j25bsH76X4GEF
qB+RHvY45XcZmUWuf4C2tE2BpnjsgxfDuVYGzGLx8mxRfimDvY4ZqsCo9NWjS7Qu
Yy+GcRkPnhnIADvLgq1s9AKWe+gVwmBkk7oPpXeePMof3OrgwH64oSbLjx54sFhR
S84bc7qvp5itppnaRDqkPZvVdLb/CS5PdXQbuCU8gvoD6P7WLEZnWPSh3JcX9ibQ
EgTcTvHWE0BJrXYr8FHEsNgHGlHTpLw38JTJH9FkWCoVlgGhMo46SlZuguzaKoxf
v80n0roRY0XgWurTYTvLVo99eK8PvUM2b4eOke7ev/W1PKelgM1aMbYpA5A4yK4p
KYT2hqikPhl+isLORHbo+ssdC1JeEbs/IiU+DEirzp36pgb4Qa9i30Ih7L3epkwd
dBire+eMt++BNRG1h07ZIE5byE9XMK5g+QT6euAONSAE7FQxWxhZujh/TZvbTcZd
cRngzT0cgQJKAGK5UhCgWp2LfGDJGj45iaxIStDcXQwXQtq1RI7gw9lmEdA0nXmL
kzk3/yrKwD5vMtOCtWOihXGFTvBDjZA74boOoDGq0lFQj1fUIHZIbpGkA+mH+HYt
6EJBKsOLzXikpKTsO885BAZJmatCkaTxRRrYpCj7RNDS/3KR+aePAaAZpXAGhATS
44c+QIb+YSEzHRb+iZwoHTthKDbhW5MlYwUznlSmN7xDcx9C+1rkPzoijsykoyXP
sG/p0V7IC5wUGvgH1xnHoW8X0ft8DXBNwPJA/OoDPQyrndlxG4/jRf4pVHKe9F8n
HMgRvbTFmf6YRGnXE/fsXzojd6KTzsqkE8VJ4Tpi8G+kR46qI0qNwYDl22c0k84A
L4HsRuDkMt8eoE2DemlwAWNHWP3HG0YKicKmGGz6Xpv+SznJLzNGL2lhYQzhDsb7
gFSkeXm0/ON4jJ5JVJlenvrzh54RkrYXxdvsczmjdr3BiKcQQtYizKQsBIRk1fPm
aHFqOFwGjeRLx0itKNNGI9jt2S//2Pv0eJc22o90DEi2S2FBmk1l9ct1wc5HIkto
KqTtGNRvf83AdgWAKL2zRRr6v0ekDwcAViBSrSMozLPILB4wR8zXiMafL3hgEBS5
rF9nM1p4QWMofdR2tC4DUu8yEQCs7bUvAehpmdrRomx05Kl/43ww81a8JhK+fER4
ShAed0GOuJ8MhOiW4vMhrgsE3avP0YBgGQrWj8a4vtqHDHe33yPNDUUPUivXCQ9e
J+FOQcVBy1JDbXL542LFqRIeHj7dKPzQNj4OHmxgLqglBd/Bved3MtRqflP6f/8W
h5Myv1ZrFHSWF+FgNebo1nQahMLf0fQdHad+9kjRBFq190ZsY0IcyR4gMpojDvIm
xvMuqjWnlm2JcKOBgA5iBQm43CVRwQprXiDaOPYG1YI1ol4rPvdUJaAOUM7D5200
zs9OtZy2Qul69e5s6Z6May3reH0ZRJR4KAi5w/DSIwPvSJV1BWLiO2Fcpcf4cI5W
3kxc8rT5P1bpWY4NS8coi/chK4LW39qMlSa0huTo6gS/RABxQkgi2FNaAR2G80wN
t84lQc438YMRoAREKgGFGGv/HFKHpOGPy3S1A/qEGKwtc7uG/de2KccXitFMlyIE
zYHmqO45BPdd7nwPTYpm59lQhOha1QSu4B+J3iy+tsLWMTXMeNt4Y38J9xixk5fi
kpiZpbSg7r1OVnpfjj/3J7hi3k55gUq6bsRkRGJuhYm/1IE3ru/iWuN6NVH7Tqu5
iTZkCY8B0XkBna3R6R2GX+qHaxurOW06fE4ZTeYU1RQbLXkSUEMCxrd85MaRsJl7
yN23aWZGruW6AlM2clkmiHV/+GM0QzkmSul3z+mlJWUzCXabQHbyREycG62L9azJ
3wBfhzrkIEtxLjdx4NbTWneHkgPyUj2nPQcbl0CTpmtFKVFNI/Kn9HLzDHs7FMXE
CV0SBJZ88sfLOFC40NZGybaNC2p7AXGWwL0rBMjAZ3VtAmFO1oTqAMp2CGB1Bboe
3/m3tlf/cepeSCD1bhrHJLDWzqa58He0sMEKpnPvz1imbGMUAd+nErJx9cAoN9tD
Q2UqpKClRwgZxVKfTiq/u7WqcZQHhAipom5LgOaZWEWIRqg3bynvOz0Gxrni9zn5
h0wD5dVPNJkgTJ4lSfWlC5GjABAzQALRF7UBTq8A8N72UgnQIlIlNt9aafFQxpKk
ISH5MB8An7M5ZxsWWA6krzcu/5XDryhfkoGB0UFjDel4nXe91A1kFGOzkU5wXNr7
pubVaJIzVmgJNrVV+i5/H1QeUqDUYqrEY0SGP8ioZyMtAdBqg16vSrflV0exxujn
Xfrw5qsyQszhkiUN8PBx2ezs8Yi1ZIKjVUNQfDO5HB+ls1KaJDIcMJ/E0sjT3fbb
83PctIeaSpNcSKB7ZYHumLoYzVnsE5F012w34r/xfxor1bPXdBwKWeLIuaOhZsXc
WZ11rVdfMxNAlkzZqx7Z7/SY4b5mkK8haoko9LXVkGigmnNK74D+lzTAKGQjaEiX
ZpPThQsQWnQUIk26/KrMpzrMWBhm7oUhkAFc+uWqkchcgskoI31ZoG6z5SqCiDhr
Ig5IenXfM86HkVr6JruEbwILCpHNlb7QxY30J369PjR14iBRyNkUm0ltAfETxa93
mMeId+V0sTlJ+WdMaBd8N9zbtlmP+qCBIqH4kPwz0x733afgIXAfNJNKAweELk+A
Msa5doEkiR7ZXuJg7Zo7JJ3WNLhuC8A1zCpGhEDpDkiniKZfYvIDbL43hOUmoo2E
S+2hXpRvbtwt+0toFmQjGMygViyYCTwd4Sdz205MYf2c9Gd786ENaI/BqRt1IUQn
cWY7t9yEDCBEvrzVBHLxKGQT4qM0jSgKxsQAVdvxnXKaXfbOCOmLaZxSeeC9V3ax
KZVOC9RChZ6EV0FVEszmkDZUZpTN3hX/aIdEdug5siKvsMrW65kLiPRVWsutsij0
vFsomY5DkJ/pf51a06dG0yTNNl8lojnnfWZ9t523gQxeRIQqitHIiQ043xKo8a46
ZFS0IwF8rtN3Qu+sZ4ifgEehy2ZLC/ya/Is6lAobHJ2Inw/jPMcvnQ1izRO3EJv7
6U4B8XfBT/ygEcnGwaHj151LJIHrQu7byyLWaYrP0817Dlry8PBxZeqWIrLhWoYX
ylxnReJLhPaiCAjIk9t/6wMPEHCnxL6JVG6+faN/bkBk2ssawXRnpoEX6B8Cvut1
1EYE6yNY+lzhSP1sHP9pqrOvGQSExiYdUpXvmZe62FwuEBEkVITyCESUasBwa49M
4ItM96eeZZMELJzhmDBNOXn2H3R71AB8/ulanojwHOD4Gj5w7ilBVqRjbE5w1jwl
eoUw3wrjhTgtL0umZJif7mtwJBaKu8CW49nJ+FuBJtlmymSOHhfcGZ5V6U9Apdop
WpJNPz9m6n3MI4l1MICV6fJHnoNxS4OM/LZ0Q1X9Lwk3RE5NZXdphWv3nzjumlrT
Xfk9/meNEBQJmlD0UnPC2lLE6Cuck8zgA5ARE6XjteDRIJy1q0hskIs3XVQTVJdW
UC3+A4KCp1cdulinlu/s9FHH1b52Q41oIQ14We0Aj2vN7PKGOfJIXscPWMtrbFTr
bQ55g3pqnTz2tTw+0jf5hrWiKAKtdhxQleDGOzWBzR+nJeW5W5cE1tiMmD+XT18s
vJntGq3P9+e3WqVFhMFrWQRvuYC8pYx9Qw0QVaJSEi4sA1TYlIyr/o9vHjmKEGlB
XAYsrGq0/dluP7MxXlDn910IuxbNUkQt+9vzAP/rEMpI/9khE7VkR1BY84xW4Cpl
KPvbgKVel8PrJXyNCuBH8d6aFGcmKopER+IEvRLx99as5OlLEkMsd0Qjfx93KlB1
RMHT/h3oWjPoW/f7pnKdeoiiojlfXCRE+AiEu6JMCh/Phuus5fmXZw7GKHhtBBEc
FMtr/lXYZWA2uy90fPD5+OcWW/NvWX3fPKx1c6L39hS/U89yteQ3w+bUEWmUSv/e
e51vKmP+A1mfnVoxP2m9Zo3P4WxMvbUqsn2IAYlPB/+gKhM9tNWLaeq+tn/uM6hD
uL0hmCOAH63Pd3xz/6Q8XkqfMaRo14BU72XxZOIRRe3apIHKKdrWYQ3XcOfF5Q7s
6t7uSFX4N+RDyuYjovki1XBOa1YBL9U3OtiFX/gFQlPY5n+i0p+gUzlX9dri73/+
ZTttNn8XZwZHneHa+z+GADlF23JX6WdWxVEcsTsEFEZV292xZCAQzsD3hmXcWQt4
KLkLLChmSQdDJJsKg1oNvTIX2gN6348gEUu2EnXH+pKTj00Fdta1Q+//YRkuxOsg
QeIGl2RKJtF1JMziIKMVPVjCd42y4+SNcxSeNM4phRNXuHRwlyvWaRxRJgOxRdGN
bBe0giGbUcdhZbSFn9URS80nwmLkvSPqnoi3jezgm+Rs2LgWrZjOLcsh/F48EFzR
PIMXn0k+wHLsAPNELtEc64fespaAYyw3dpidpRGvALUP2A+13omUTYdYqIMs3b1w
uiZFXhtFXSuBwq2diX/eNv6VYgPDYB+dIVhjxpiZZzjbwuBieiC1eZ6IXmEvM2GT
5yLUbFzOFcruI+F4SZv51Fyt93a+zujyIAmudCuojOwqqkxwAPekz6ADI5LJnmvq
LnyyY8sATQCXuwHKJHSYsBQQ+MozaJwY6LvC9rvtu4DzwRxK8pVjyrXAxAscipJO
CuICLjO2xFa4YSnqhAdbDwYBgFdjGxT0m6cRwkqauWCUYYdA4o+9spkmUDIDslTi
S+SaX2TZfdnm4zyJtxz3EZPGfJHVvwWIuOvIsEBidzRMhgljZd3VTuKOX6YcsSU7
ZLtwQTA5jSleZc1nuZ7W4GzLaUnFeTRVaNfFSTRLd3PYAakmN8sl34hm5tqQOkOt
Rxs4KuHUpTERr2lfeBKhQ+BUBPbiNXy4wbZFNKqNim0TNRYxdAJCNqsP+4yJA727
WD2vfP6pFbQIhMd/+JnP3zqj+8Le2yZZWrOJVMjM73PHg8PhMGttjFJfN4UGe6DI
IISl0t7rkkWHtTNXYxBfL3FDVZhneOAZrQ+/URrnc0RMinWjj9JzMdyBEiMP2128
8IAJr/6Xb0rnnX2/3o3m0e+k7CJC01tEi7v5BNPyd33/dmsQWMnSohOQPY55wjzO
W02YXtEibqvGPEDQ/NEQlIa6CHvARtHuHTJ4TVzpqs7d6gF2LhvzoFIuVjaxo3nX
eJqCUBcTG8FTIRp/9My7R4ofBXwNea4uMuW6gn379WWZsPF31X3Swb07NHoJ3RUU
drOKXYeYSLmzu04QPvjQbZxNNTtlVNKI+N2iPZIk/y217grcFMyt7UGsJt2xhyoE
dtplwHrmAlybob+eSXrI/UF5m2WFNXdEwYbAknSlKAiiuWEO41CbakSeXTozdLBg
XkisbJMnwKk/fRIGfc7xmgmvRl8woIceSERqwAN9+7IH07LMcKkHkxG09TEHQbIR
sj88AR1ulEx1vkTx4S0sygbNqPXUM2Zp5Y+IJAp2p+w4UnrQ1Cshd20XBLCoMWXQ
FKQ83vscUYnhbkmFRnTo0xRUAyCDYMbR6Q8cUOV0s3ga+y1pVpt3dHr9H2OCwQFh
vn1CXrmdM4MyiefNDtl6etMiP+S1EHYY9gVMqNmcFFfbHjhX9QCUkl5d8Zlxtevt
+FomMID+4hXyDrlAryJlqXvpa0FBJnSJL1eT/Wfg7dlt5GCFaH2O9xOuT1bLqfGw
ef6N93eLtdhhgbXNFWMEQYXuYJjFDzlKaASL4+0DvquIxcJdWTsmVCuWakEpUY7R
scg+61Es5bTyK6w5u6PRstdwiG0MCgwB2dCFU3puiJ0KZvjEhbnGw0a4NU9LBMsZ
BWZWZb31VhuRoTdARZ9dv5nV2umcHPkXMtbXjIMF5898GgK5IA2bfqrO6lKfz6XB
pQbCidKvoItEslzApKsM7AhoRzEgatPNTnxu68HYIIEjfZ5dcdX2y2/PCvQgyqwN
U/t4etjUqDFYbj9h5RGKfQx0rsFFZwWFSxYc/d0yHKyGN62ZPGm0sPCZnpQQL9N1
Vv+XsbXrcgIxn1WGMGWHp7f+jkYQ+Ztv3WpKiOUYrETOq7quRCkSdKIioed3R3z8
1NMxX0Yne32rLEwcceVNsMGwMHzIvGSJabPvsvTbNprdsR9wMsoR3p0wcT5f3bit
dJtwxZz1MNUPXTNt5+xIf7cbK4INO1n5UN7+XRy/ibwzheug+hJXnJYUWIxmuzu/
7kXWQElCQMjKx3cwf3lyqR4BdTrlvhQJqFn1g5FktODGWc2YQ5MOtSCRT+/qXLLh
mZb0va/zaFNGr51f5Qlg6dC+QXiInuJPIez5CTfbqxmF4YD+vv/gK9X7OYlqLgXb
370cwr8HVsL+PAp7wBLvV2+xRyeM3YNWP+VW4XUJob3fy6bmLt0bOTDJhLzKNGmO
1+KcVVUMN48pIuwpt63xt5HoKf8zPxpiBNbeatcH4X1n3sIE+lPfGU47vIbG3sI0
5JJfeQZ3T/HwS9sZbigfySKxtexaabAvQpeCM8wvJMfSY+Xu31t6XtFf5tG9QPnE
B20qJa4zAztT6wlOKGaGbx2Qn1YGGT6gZrcbTSYczeAMV4B5jemrPHtOUkFupr2f
EVF9vimFh/RYgNpZt2J+qHXsiqTyATLdf0dVBxcKEqGlcWx1EusxsJ5GHrgu6ATF
sqgWkJSrsKpWSmLTPDJb0JoQJphXEQ9djoDh6K9NT0A42ByQJhWWsQRJu5Ma17ZZ
nmaoU9F6AqPBj7jfw2XyLJfsOC82RYAG5NWok2mmHjxdvdJHqc92U/3wprnrIqX+
WBwGWgqYWXowoq2c2zLNfNDcbKWky7/Rm2H0MliTYNjkhOT9IEUFzJu5+x2XOsU8
oBKzNUyooaHA4BnGfG5kZoVNLVJ5x7ZfGAmwDqpV30+LpnHaUuAEbfiv0MajR7RI
wsGMKMICQWEPRWoXGIh11Xgr4V/SpJbPuLgxvad3kLYR3JVEEHCKJq+wPPlmH0xY
MJlNNUQlEcZb2HQIoCOZKlBRrp9AzPDIvmW9EBbZPio/A8KiaR+cAjwMvMblL0Os
nW8H1jSDqYz6+mnle4yY8x/iB5x1ohLnb6OfJHinftszthKP4zYWPJvSWkWk9DlW
iaSgC9ZlaaxMctwVsJS7IFGkuVVAuLG5A/9mvn5WvxXaBjUKuodr0TmLyzTmw+FU
euQJLDOZ3FRzudlc3yYt1mdZyOKoGh+O/NwQwfyHx5hEMEx6dz6P7KsMFb5bTO22
8lT717ajwr/i40bEcsr1VW4ugMNrLYkiY7e26DfIMWU3F06Gx6lWSE4eS8e8D1Gm
1LLLZltsX1uPMTIv744RFE9WNaWQ+I71QkUzOtydR99Om1JpIrBWjgEVw5iO7Tcb
JB7zvNgO+oEYEjLbtF150F2yis6Ze2VRAAPD84YTaW6oxcgqArdn5s3FYzokT0Ho
NcU0hIgx5GxEuy/DtNUraEfsUpWkvxYsJbF1CocBeLJubF6JPDNQMMOjeYuIW6Aw
sRyMGFopIycA9p51EigL6jtmEJtJAeP1pEvUQYt6iLRqxu9CIP2idhNWfY/VI/2w
BcxGMSsVE/0DLPpmBhzY0nhbz92R+qeW8QPnAu58W92eeotc1b5TCzw+k+ETysbf
8X1wUS1qVkLRlGovt+1nwu0ZLjXYv/vwKXszCq0Rd9wceoPJEQkxole4o9tmOevI
NsKlkcWb4lO7LubJk/KT0h4W5EBMM/2fGMHn2t+lrZqSlvQhiw8J+TILBlr1+OaR
w5ZL/hiIzAH3A0rnwhr9AaE+ela5bwGcUUe1/a3Ev1Kz1IhbUeVaPBbNnImOCjzR
Lv1DA1fNetiK4bAStRaSDheL3xgiFyZHVgkucmi9WYeyhLKhUXUFgmiW/5tlwEZb
+Aj3qOYkIypClNk+20sH+qUSjugPzL2vBzfQdVwYY3XL0EbKGsltFz7oB7/a3+I5
1+TXA4657Do3ixY7hUNdXuHfOK3UaD9jri3oe4Q7mCB6aNZ/yBCqUB/6TrSoh7lO
Ic7aMneBfge5jsFRwE8m0bJTfkYf5s906UHksSMATOnf7AGNOiXFJ6yvoHj7itKn
W88OrqA/ZblC+9n1k7blUtO6WGLmwtDctqmtNrCap++1GKd7TJaDfGakCSGSnGH0
+qGl/r4TIK5hiIRWo6qxYSS/oGaUW3Fd/eWbktPHiweynA+gW41gRqDNeAkgpfDP
k94eI9pMXqgP5whdq87itTy+hGTBnGe7pd7S6QbvvKkozixnq8u6ENT8gQ5DWjUS
EtF6PeafKnf0gNpfYoOM0xn0ZynFR5UiwNg6GoTLE7oe3RDR6CnLpZ4p/jU8v9+H
4kiUnURU3VGI7ZGTYc6Uj0MoTleDRNlOfBBhETvRn9SoNvToOsl0+ESpfBluuxdJ
K2BZ8oybZSTSF2uTnOmyxO8KE3t3MH2i3ZtdauH8D2w9UQNyOLHUB9XOeClqb19q
8xeoNzcf2RI89KYiZjSrGc7o4yfOkd/YuNp4rii3T4snTXEAOQmCLR7KZRrLLneo
WQr1sLNbKFxQk9P6fepjrWc/YIMoH05YzKq2XBpDsjPTxvHIS5OYqFL6iGHQLxZP
7JgzPd4J89RBKt8bd3Ci2L3bQnoI8Hs9aRiMrREENHg3B6L47CTOr5+lnchCIKQ6
AP7HHawWT7wk55Neb6k2L/BWs1ybzTQJa+bsYJM8CXVBUcdTloL9l5NIbpf916oc
pkMs1oucsVOGH8vMo2PIGR/8x0Erv96f0H+Ie97YBCcai0fBeumDKkbw2A4+b+2f
3aBeyiOjCEuiyFaGfV7S6rlCe8R1GlHzHwLMsqj74YPKvWQmVQ4lz2Yf/Z4k3FAW
P7Poav2cuWsOus6aFYrvudipQA4Jihvr1JTgmHMGmbPUdhK6BNiuQ8bZDj5P8aeF
e3B3xVne0m1HqQ9JNaefgytbUBXO8v+Di0nSQMdC62kJY5BTWMEwQJY/zJ6DXvCQ
nRDWsIo8VzDuuvXx0TLRrtyeaPxHvis9gHxj5ZsJ2Syk7j+huRL7RPBUMEHJYvWe
MF1kbeADYOuHB+2c74AcpJEzo+Fnu1ljY3dZBClQXnVTroQrEKR9qWzdVJJc1Vdd
9ORgaHZBuT67dQRZIYkTatyIHPCY/af6/V26jBRNd22BP9LPfWH3RpyOoAXRORXz
l9kfstOWnwEjojqwlNncqe57OUa5927cO/Gw7MabrG6VbSetgFAJOEpcMozaS2YW
vXAYHUiBOGcN5/KM/I3AXxelJ2mhHN4GBaoNqRyxt2AY16Z+gzgB6hEAqp4X70Lc
vEE7JlgHKErP7SwVf1ktf9OJxiThPi+2ijemmi9+u7dphDECnv3EKWHEgmdktKlE
8ZpCERmL3u9PJiH+oyNG53nR8MuSTxczxKAJyjyfvxMjiDnM9V0cGRAbsmoquove
78hWGR1BcLE+m3ODXNSBxtjnk1tUfPVxfAVs2SinJuHLZsOeFDEEuGPG27af9Co2
TNMQxfZIuxWVtom5baZCbogvB2RlXfRoOGQE4APnwbq1hZn3jIMeQ/s7T7MKSts0
apcwD0rpYeuCdEE49zcciV0rZvg7K67u8PsGpz/y8VGB9Gb/FfWqHr41z83HsCNS
3GBziOdAtgFAIcertjI3uMJ4Ng7zsRpB6pajPMHcNe4gSoltMSW30HqTqqVRp/wa
7uAASstPxh4FqhN2xTOE6gt+eS3PQm5GZtuS/C4tqRx6nJEiKsHFfmxgKEJF4U0O
cYZGeFH65eHKpTl0fx2BhZpd+YrbAihaDtg1l2zoA8pSnhruMI0Yt7w1CyfVQn2p
xEwppxV/Uh68JjR53yJNWkng6e8Axtm1tHtUuWvV7RXyrnd1v05fP6KmpNWmrXcZ
O02N9DyleWeZcE6kYHWNeXCbL+AFY6OseNIpvFGqHFn1aYconJBSKW/IphFb9wRX
2UI6j6VxNLyejUiiR6sU32s0+MFk/faClZneEq9scmviIqnWgvALmjIU4mub2HmQ
uHu8CN8xWhPoU/yZlqG7AL7K8uzRZiCtinQO4JUFX9K2VLY43NTvtU3Eu5vbGpaa
JzWM2yXQlQh/hJmjdXtWLZossVkj/QjgSx4iZxz324vETdKFPGMBcsNw4Z5FJDsA
FW8N16v5zdnIBsgqoKv6Cmt/+7mR3Lpg/ii6CuPYp7xvK2X4jjCgkIId8Turq0A1
52KHvUlNBUU+fuUoWCk/A5T838DxjHt8n/SW/I24/p8Oh4c8IbUOyaEU3FY3A7kZ
yzQkqTNLNRLXlu8ZnthyHpMplpHnWBgv9eWSColrRfVyC2pek922jJO6vfmrtEPe
rc9hqe7TVvKlQ3Ysjfm0OLKp4CaxBGjEqVnuhzLOrHckYjlpdVDSVlVgxg/6QXqA
9ncsJPJqgu4JnsLg9jACkI+rUcEroNn+SvshAxQjmbJf2zxbwtdEEJkeCseKLvDB
/rC60KOgLzGeZBmIG1hAPOUWEVrjQPKAgEfJ+CVlxgRklah/dsVIC51/SSg1CQM8
1/ooTA9hsJE/q20v/L1opwixWtiPRLK5GVnFSw+z6eckH9KBKwMa6nAMhVf//IQ+
sMhMxOXQvs7riBzqbNuUZX2vcEYE4HQHlHM8khAffK8SOb9lJ51rKYZeIM4nH/+4
Kwe74X3t+1BiLtxiLINMC7NhA0CjmR60GstKb/O6JnXO8lXcm/Z+fP2Qgfce4jft
qlPzM7Sq0CEJwDhPTCB1FBTnVKpQGzd1ScojDvDB4gXzY+NbpBFIOs4kJfto6bgf
Iqz0UOSBTiMQ0C2NjRVDcEtuGwSiRp32C6EFk2SjKQnn6HFYzffwzDT7pA5NHE0P
y21hwLFq7x/TxO2GMxJmo8Gkl/7m+TaZnaWrcXN4ne1GDSTjTmLXGBGAcUEShey1
+jefuJeJNG61GTsn8/nI5P1oHOTYzEtf7G0iD6MO2W4IwS39OIyzdDn1TlX3vD34
h3YhUN+EGVRUHrriEj8l8e3GJmhQmvY0XinZ55pTFNdK/Zng2A6jO/ezJZg2ury5
aM48box5Bu0bFVVX4RK8fVuTKcDBRal4+84qqeVzOtzg2xr4bv/nCIBJrdVPW1fV
CulJWPcbvE54M7mRBsJbWYpYSKmFDJtAyZqCRKZi9xDi1O+wTxyxwRjJ/1oWKdMC
ar1BbNQcMUNOyJ9u50NPmOGKwRDWNySCuNxYEAtmqzG4rz45WQ/o3u/u3zH479+9
r8MBGrdlmT8mS97BDwjhAgBgNdiMFou3H5rPbpurNZWdax1gfDOhIBhiEwzjAvd5
Dz2WVcDfxKSt9Q7BDbOibP34J7isXfmP3fWh2RjqqDw9j4G7Akr5jcKCKSRVijKM
N6uyGNUbpzYIyMjA8ai8RcgB07e68TwwwtP02d1vUbbXEyKII9JNVsy7lwy1QOkq
ZR4N0o+HvVCDMtLhDHMUQe3ECEMvZxgvvHxwu/rs9zaH0qxK6QrYDD8KqF3JgBcA
X2ayl+XlUW2Gq0k0CBJTG0iuRVgoIlxWAfn6qrmhnt2gYpRCW6a3fB4/Fa11zY8A
I17Rwu9snWxa/zRsfZjxhSQMqXX0yQYvEsUIuL/nP+X81DZZBVC7b8K1laXhJx3u
BPLKK7nGnAxQxBt4VGr2/ewpWY4+kOpSRq8MloTUEm3wqcx4CMz6jzegIMqqabxn
hAYRGIdWLVUEPXDSyyFaTqx72dpMJepno8SZaLoJetjcRdxzK9NJ3Z6Cm9Rw42er
Xb+9IhmxbUd1Qa9t3Gg1dcD4RhuwvHAvUSGvn6Pth5qcD7wUHMIcZf9p3H+JGY9P
kNA/LwPFFTIgu7jeEf8aue4bh8rySq9b+VD3a1N+r3qsI+nGeQ2t24h4mP7dHJAN
O+eFYaK/XNLt/aQMmgkQbZkXdtfV+iOGvunG2zvERUA89Rqr2j2UPi5oGB7iqY5T
0xDJpho9tmyadnV6Oy5W9zptXeTVZoK+D2ceKGLLXHHKTCLszzI2KmHQg3ahQZvc
fT8FeCsgMkh+az6vYe0JStVZWkB65KQXpU27adraVJeh7uk21fY9kAncBXMqBGB/
WjCfRv5bRTZPGe2vtAHUS0orrq9QcxnBa0bSYfKRGjfW08m3iBbZwF8Khjk3sArD
v47ghukQ8FIqxbEp4l53qBhjiEexbLB3UHuWpzMGDL7C++xNgMJg/Iwzzp48/R5W
MKl8GKlRsTeGS75V3Ly1E7wZ2hNAqYLni2//GVkkjkJ6tAdwsG5tLrFUZYlz4mr0
IRviqKzhxIoOXIurHNTZb8b4AkhTft3anNhl8W81fsxsZUeZ9e0Cd+8/x0rgvV1p
h+l6LImittWNXUxmyOWo2fIG641NeFNibercpReWNtNNED+7cfwvasmmjBVlnmZS
H96kZKBlQtNBbJ6+dOCoB2sORrrd1O/iqSgCx5asIkF/dhTeiSrS7X+ArAUfmu6+
06Wi6KRVeOU3ioEUEfvPTlI/1kEJRoJ1CaPviC8RaK+44p1vM4EfVhvPNIhVFEoJ
j2met3urbTE/zFOArSrr10Agx7vdTidAk49sFSGE5e7gQjtMqNTXtIOi/IulYoPT
kT7S9eVyHXguuZ4iO2Lq6i5DeS/biwi4M7tjXwQ/PcB5aY54+2i02ptJOwjqabe7
AX9s5sgSOLK0lGFpPS4q3cat+bxGg4gNWaNYEEkIojAi3zYeBKz0DcwwiC9kILKA
122ikNDNk7hVBT6O8BFAkh0JcQ5TI6fSvoo2I4jEHJu/+1pnA+mQDA30K2wpZiLH
rONfaWeE4Cb7p99ru74V60n2z4iBnl0+lmYFYrOHu361FgWl2DUJl24/psN2jTva
WKJBUwJ0kQ1Jn/5OmSOijxDN0ZULpEjs21P8YWtj+BWB08h6ii53KbEV7iSbzyzs
dvDc9aB/7QPy7dU+1F1Nnc0Af1JJ2C3RBJCygqIcbF0EfvppyJXABWMvVY49fJvC
KHL2OzUyeRtYNdhlEkmDw5QJJFvffPXTXK8hVcAjTSZ8jSdtWLaj0lOGrzRfGxmx
jmdgIDXhC1LUdJ96ye/Ff1L+lLe32Li1f5O3fQ32CmGt2JcuChTcALxWSmK3SquI
Nbz73PlnNC2H7ZLXPqYMFOpNhsqKaJbvqw17q+ZQoUxBAjyoQ6Veb6DBGO+Qkygz
fV8x8krEYYJIu9+KGZ57sFAYtaxWkIHtXL/WKLYjxnTjTL+UMGf8Jimt1DOXA1Gp
zZSuycT0gr/hzneBtY4qtD4GHbJXp8q441LHPmvBmhu+ejMyODagxv1qZD/TJcLq
EBFXCsmukvRkR1TzV/4GOeAPuPqPyn8di0V3zlL2ziiIdzPq8D+FiUCrzofK8qNF
HClwO048ZTZTQ7EL1y87P5wKW1a2Fef4sB3kuLpjc5S/aM35nt8lAp+zKDOXyyAe
obJOgxeFL4f1Bsls8ClrPjHYah7BqzUQSnwbXaODEOoF/mdCDnOwAaK91iFMGW4Z
AlJ1vZjcnGMF/xZAeMSSOLY6X7MoRU0M4HCqIFXZlaxW7R2A6fz4ablCbu1Ritk+
VYaFbj+rMJVitYtujyU1pZ3/282YBK6oUB4c4mRxcIAEv+C5fzCNwaKPtev721+d
75x3YWshZvMYj85T7kypOk+4nI0EsShnvfYNkUg0TXfIo6hdUWSo8sS4em8wTFfl
UpCKaGRqjfGGFjmkRCCXAMZfTAuO8c4houKRqAB9VlCeV/l6QOJSgEmcfP5P6DYf
ikjs/Ywyp04YzQfQMTyWxzn1d0AcGn5wbKGBvTW2B4cNiAprV+Aghf43/4GuIZWo
iEKCY0oL8ezY12T0eFinEl6r1JFxJsY5tHe6J0j3AMKMhZCPUQm6VnAXwdxcWHnu
+WpsN4GixvR34Zqz0k4+0/Nxlw2eH5kwYCGTnGDqV3ONH/CTIcmQZxokHLFqc3CG
NSS4BFS3vrHv0qaRc1chamYtpF09Gr5F3Ct9m4Pt3+ZMJUuQ3uFcadD2DJB11FJh
e+1dqV648nZsQpcZjF4MXwq3Q36z9PSowYlGcSFzP99cWFRTOBdoZx5qTOgKL1V2
vcIRU02l4HGqGAIxaZ6ONDgZMV0uXiLbRFSeW+16mz0D5NpjN6h7D/lrll2fWAvl
syI/3npsEWX4ou8dnNTnthU2RpdZecGP32vSq6dz103w9078ifpAnbat1drOqP0N
zbYLk/0LUQ0G8VfPWE2juK+xnYeIVbBJPox8qU1YGALAG852YQiMIZCaWBatobg4
N/K3k3NFzQ0lITjvVqYePaex1rG3ZqMR7PqCl81YrM2fdQXOOHKipkBr9Oi0h/V2
wfy4xQ9/Anjdd2xzWo54MbMTnQifHrLXWCg2I2tzSkjvkNPVjdNMGk/5Mb4cPHlp
N7ZtZwLRClFeGCoNY+px0bGGAGi2dQa3fg+LM/vZPoyyRfravpFA6IX4msovFt9N
C9MNI2N0u7htAeHKQtcZLmJ3HaDyl34LfG5nFAVFSc8bafkMpWHwOU14lHurE0rD
h2vLDtJhhtshB+KEpZsgYeAMR6oEuPKaJJZY56UqSypNl6YJTpay/z48s6YH2aPW
gp2aEOj9JpFJqwXS4Koq4TsRQi7PAG8Ox7GixewhuZVD2CM8Szm8AqgOxQCBkNGK
wsKBt7hsLUja9DRwq1PECxXJY4OKcFoT/BwWMeuytDfQqgklvTge/b1dUc2pejs6
+maooNaqQSnF7jlWkYzsG9O7yNyIagWCHAfIE9DyBfze6ijhNgaWt0MxjUNtuB0d
2EFxsgn4N86kH0Y8Hh6twqr/jefzbJaJlIte24LauhMFEt1YrOch2/tMwZoiPa5c
EfUdEtpiQdr0Jtuzn1yJqTeEuYOEIs9RRq7SbHtbcKjNsIUJpfE0bk040caHo2qU
vJ8fvvwPBgqtn/f+PxNpSEQLCFo0tI/WAY52NrXt7VK9xtEmoDd9sIEGRT4q5ar0
+oHfEEhBlbR3SxF/XbAg8sAP24JQRXVfxIucSSNj99iIN5GEtfnZzcWX4aRzwMDw
+MqlQwAn+fE1A3cVLAm3wR6itxbx/wyVBrIfWXFgdD5V5ea4DWk/EBZD3vEqM8HV
Bt/TFqV2cFdZiJ9NOKgsNTqxb6caXZ3uWAcXmcxKjvuAWbg9U3xU9Kj29MFxNit+
pRmp0evMT/ru/wSKVTTdMsLWFHV+Rvln1whrp3e1CGQB5G0foMLnOW8/1Uc82vTe
xMMILv2zonuqUnwYHKPygBOk96iBbYqvGDzgpxFqgjo3HGfBN917nPLZQo6EmLfd
Mm4hFuBWQaqdOW5rdObfGkF9kAK11SqRvT2eDbEUZGgVCx/erO7GwBhW5bak7Ryk
/JYGRJon3g9MjwtWJiQ4nYYyqxfM0XlsyUANjT5fvLKkfomW/ITjcqwDQlemY2l8
iOAZMLxigyGv0FHYOYmBR0RrytA/W3xa0hhuEj+s9tx9OvMcEJWHr1BFWOp0JEqi
BRiwpJY2qiJ/Kmj09LCRJDsVOMD3NukBEbbrY9K4OOEsptgd0rUd8ncj8YFpXFCS
uuxjLziPNWfG+tlsqG7s/WR79odWCSS38GfuUNfOE7RJ3AFG+bG0OvhV3aOFyQe8
dbo60dd5UUIL/6EbS8+18jj/yOLPAlNtT6WyUzystfcHBhKTBUOSXxt5wTAM2x8a
sCH+IuF7I4dnqw5J6w4IJyQpNW95zbGG0U9QUzlnfQOxPIA4nZApolD8OKVxP5FP
m5tDT/cQClre0aUzhRYPg5SDjlZB17jHPP5TMnSMcYFsZLlatDQrMpAbTQZ8qSds
5h8HG2cjIYNJatp46KUU56lZoAHksW7eA669KJwPEKvOClcNvRSlrUn5Ye8FVS2Y
t3kcI65E3OXfzvuil8iQn0lzmadRQMIS5omFxCLyyfZyty63jeFvH22STmcjk5Mk
khzIfHUeoZWQaKsen8twrvW1PJzwc5aqBogfWqyWdPmAmQMrL0eA7XSZLrrNY8Fg
t55QJDL0Zp5CXCBSkFHLaLPP3AiOSyU7m8dLmnpOK98KP5mflXhNeOYc4nBTaFIt
I0xf1AKsneFG7MUEXEXNbFC6Dw5vULId/N25dPHXko42t/G3gd/+bH7tfPk1bswD
q1ngXfY09XEoDYaiE419m99aBefZTJH1TRO+o5JJuCchwf1QrWznLToLbRCW8m8r
sQLQp3tZADBchvh7/jk2NiaTTV7IZQ5vT8j9mGoUCO43WU6jP3OoyKvmvmqVQLpI
XpV3NzXr95VBPO0ptOFoLNYB0ucCm7XW7p9A83qggpRQ0VoEm4n4QsKxnkn+ZXx2
p9CybQxYLFFtfaaKDtzhVVj6SrQO4uSaUTNmbMBGV857jb/wIvkvRoGe5SWxOaea
dqvxt7QQ5zIF5esLdouWYpHpmNdlIZ4bIrTkh2m49Uj/BGrBI6YOduCr6Sfy7oD1
kCA2THLNZ83Odn43DvI1KthR5mJBXALuIj+TPN0F22eokejcxSJoFTsZqeq3kVCL
96vBpXAI0EntZxxzQ637CCN/fDJpXyVvuUkFljDae7EvWUUv4eHcflnZzcZIIcvQ
WgE6MroTEQFbByuA4wMXHPdeKNNEfHTVCMAioWJfH+vvEgBz7CffeEcWdtr/a8FN
LiEZx5TJIMPQB449B7+MLlu9rD09vA9eyOm9/OS1PUSHu5+efzIEVT1sGU0Ddrl8
Ct+ua7IrUT23+cf8i6XeZntvAMZZ3p1J/U276nNAjXKNEQb2t8gnVeBx1si6O8r4
BBG1aFRRmRhY+83h9REMDbRMXykowky4VHpejWuiDROmKkq2rRLg8/YDfxssCR/e
w14hUkWOJEEDZDhkfP/w1DPxpTrwLWNYIyCyrjC0Z2EAEt7p38uwn66MCB8VGyH7
keoUvIMBgRJsp+3gEUzh7fV08laQilqKWonaBE0ehVj05AdOn8j+3iHlmIE4gYgp
jpY4iddmUSyLwIgWO5O+Q7qoBzkdR60PfdITKTOiNJym2MG9ykXcC1pXg1sUpMsZ
VXHsFWRgI1PYm/fP/d9WSQIuiDEdAbbE5LzMzbrzfiFFX60PCGS0u32aaftggkpT
mUMMot2k2Iwfs49txExr19v8pXmFGHOmmb4/0pk6iHt6j3q5SPnnzuAdRgPXjKgb
Gv/g1TpBCOgYl/ciunsUthuwXxE2MktW17SJntBFsMFAVj2zrzG531+clGxaSlpd
A9C14WZga+CbozauH6bPHth6RJm6BbwTi1LUma6jlauFr5zcn+pYksqqc43Y5nWo
S8a10CIn9mmhMXPmCRGgimc9CEVc/djDqCtaqbJFMgYE3/1dy/fu5v5+tdM9uM7R
vpm3WiUcPIk9d2ZYyDffp43EMgtAIl+RdK7V21rhUZvVR4KmHzCgDO5orgJZgYx7
ZgiYM96aFlixd+9W8NdL8MYgvCnieglLQwsMQ/1h3NXhDoBOOp2FCcyeBUjNFk5s
V59k6uKbYI86XXccw3U6iFtOa+n2UyEZy1y1v410WUhu3c6qSoQxnHq6EqBugy61
/53j5w9iZOlHWdgDX8nCKGdCOjSZXs1YEtncJfc1mC52KoIAh0r/ACWqJEBE1G3F
AlRErjjKheDhCbC5lgxv2XcNvlwl13pgoalIZt35e52DZAuZ/46GGWldhE+ENbfP
pecdtKoV9vOjRyFdpJwWnO/ogG+qaCTsqOTfOcMYaqP5I08vTKVgMms9Wov7BQ0i
SJ1JoY4mCTlHVoFIeuvCaHZfa4aS0/ZHx02fkiKNKvWnaUXNH+sqveincRmRjEgL
Z03Uccw/7exJgZenRlAzUguz2aZiv9PcqUO1zui9FNXA6QhBMIEfPIg72DahtP/d
5l8XToDPPhDIm8vj9Rjy06+cnU6pN5mRvJ72DGGtMhKhOTmOVY/nKzIbaBR80hXC
69L0e6FJS9MqGKYsZhFf7OmYebwKT5w4ivlwi7j8NVgPR44kM3jY9t8Tfl60wHAs
q2vuk5l5Idm9j2y/3OCVHc24mwwbpgvt+QQszV6/ZXGTI0z/MPL/ccNtu1nBqDwW
Hn2fgf+QbI7EOvSVqU0kqJn96eOW7xKrMPOxBXYF9/M9tLz+DtIV+NoKGVzgLgZd
EZLmTgs2vi0ElkLfH/ME00hq0+zJ/bZOkvCIubqNtyBuBsvX3cFDRGbZrjOTL6tk
JNlEsCcNGzErtEDVgpHXzS1a7Pswq9e6Vg5hUdubYgJecYe7ltHVQhfor6rPps77
XRrIvwCIuegQHcXQvd6q0zn0Yg+aOIGz2OGQt9ss3SG30RUe7ugyUG7ekGXO7Zqu
YCkDBySCmBTaPEDph/llvuCiekqGKLhlRd5VG9hcQNGv/+/bKsjCl575cUNjMj6M
rc3F/FMr9RjNnuHkUpSuUUmnQ2+VPW5hOuluYJHVEqw+5mZLBj0LUqpeStsw9g4x
FGWOklx9bZWZ2mz+2WAxIe0cOEyfXpBfCA3nH5Dk0qT+8vw/5V699qYPmWgo6Oqa
DTYhHJn7rWwHhFgI2rK0gAQMndKrmiaPbqomrWEJVyisOu5cHKsL060uuVol0IgX
hX1ZTio8JF1yF0wAvSTIQy6tVFAQ/8Knd65YdtwGT07sBmPtt0sdsxwf5xgoB2Ge
zsJgBnY0g2zW+tIYUzvIZiNNoLTQHPoa3d1leqU0+PcxZH+sX5qe1qzaZx3A80M3
ePxLfOLIEuGAWTnBPfE1amhcyLy0T046sO/Hw9PbePdAO8mdWV7uyoBujlfOO4OB
yeuwEGF6PNffs6XGJZ02z/0V6fLBjy5RFGWe5qa+ddKvB1XDSZoYKjdfYElD10Hc
gMNTDwg99KCDNm9tPezrtx1lJiIXIMu+XLQgGKu7JrodfJjRjy+0+Za8gfEI8TnQ
e8MSOnea2Q7442kQ/oTSWHTj1d6Uaj7cKcmpr6WcZXk170He/2POQdYrvBzly7W8
2RZdxOKgZ93R/Rg4FRbaD6usmpKKAEmE+XpLoYfqVSz2t/xYFlCKAGzKmkN5UxUd
a7INHFLDXFaFsPd554Efhm78/yJwdLW61IzVETpSz+wxjwTp2kO+v8aQvvdXZqFB
uD5CI+oNIMSrUxsTRUq/wxrdJ+7CJiZYK5q+5o2BgyKp9myouIFxdHFQkzuIxmwv
C/5bPmhlfJYZ6kUROqSKdx8MoRXVrKpWOxuYO9XOZ44PTh3rJTQhmT5RduwKFacz
tXMXVesEX+Rm18HmXdfKNG8UQCsRxmcNTRBOEvSq+E7uaRPxAul7HZRVgZJt1FXq
+2u4Vqq+W0Rv5pS8+mRJi+zrS8iXWLhzm3MFIl2WgBKte+vlfyVqO8AoT52KUaD7
XcZPzhYOmT6g0kf4rq5wFJAl7XV8ROFjm51TWsfJjV5GD2Omeq/fImoxbgpdejgT
VdOMlKcxDNLsC5AGfTkFYw3YDFJ2R87EjDgKx1aPO6ZDMA7Y1WUZebj76eMUf74W
iFN0nXmDXrpD4XPEF1NmJ3EAflxb0dqnAriCRmVvjdckUwJbxlQOkalPeQwejiQR
kzmMx26FD16VCAE3UdUu8aqAg/m+phaT0fc0A1Ruwsy8kj6aBNxqZ7LSd8M+H2tX
THqsk3m/B9y+EVIpgNAOpEct+dtlsQxxaY/rbrz3cjcIIs+cxUTpKwHcKdIjoSvr
kkyS6/zyhVBeugD/x9OIIdrHNdFYALY9FI7ttJYdJsUzZlbnIIidSTyQuXUZybtx
cnXMGAPgGJQkFokqP4y6S02s2dQs0GgBYVQj9jpnL5ml+2klPCJgjjl4XVkw0+0c
si/5itCvoYJnykBWFdX06C/X+UiO2Nzlw8qp7mzx9TR3AuyPj/XtKy7DMBJ13xdC
tqkyMbHwOOvXOKsJMpGpOapC3vrvw9VWsBxJvXxWl2d9LQ4Y81awOiC43hzN7h5V
jcapLcvW+0QDHgKXi3vmAF+IgNKDAIKNz0jjU1Hgh0CahJKgHQo/h5B7VV8boWnv
GWd++TPmURCPXjdYJcsyn5PDAn9ep0O4o5QyMHQS90uJw7IUjm7BqAeGHSfd+zX9
QpIS2mTbqCTFhsduQ/gPk+8Y7A7OjKgjj/niRBdXGIuVFGDE42yCiJactyuJNjQz
XJQsZXdiETVrpSBV66AQNirxyl2r7xUOpOn1onnNxNiIn0xh/vFNFfHA8C7VfYff
DeBw49ME59Ig+o3Jq/L0AL4GzHvAwxFq8tjRobMRe4g0WXJEw94ISrMqfNQ6ierg
9FCVDCku4jOiki9ML2CrFrcXkBmZBKAkNr7AqBZ3H8SN0fCOnF/C+OwmgLJ4TMbE
AYiOahUdKg91VMiBrjObaIZYKwGS+iwrk0Zf4ASgaHm3JJqJ/amYHK9S9YZZU0Av
ONNuLMIPUMfwuBhJ2pKpmKnDiZ3gp/KUqIU4/T+yT29YVeYvxemJgbtbm6qdzfkz
SbkBHVjvPj1ySLA2g9qBWb29G+/1x6CLtDFgVAEtlW9tie7Akc2PSs2q/dZHw2Cc
RsKtqqk0nVTMNf57ywsqLWwDqL6XmSiR9v2lS0k1VCDRAtTBzO/5Qi7+MlK7LwSQ
XP9Zr5esjE+hhSQBQZyxeRI4WhgtQrLH8E8shMzYzor+ERkY8nR2hFHZf2Dp+XkY
MGU5qyCWu0MzklZc6nxaNJgVCnhxcVmZrbGr+bhX6FfNwmRaRhppwMRQcn0yJqkc
uBz1bKFoLnSyyLjUIMckNpBrm/hfKuPcXDmff7eJjcw3vl/DPTy0OjyuRfLxj+lO
rdBhzPLdGb+zlJb30K+XwLJvpaZ4ik8Y3zQdhCM86518DJ6YBxu6VimLpP9zi/vu
2+2jaYs55BC6ib+z6G4UmUtCoAIClQ30o7NG7U5SMNjCCFz/BQWxHS2CoSI6RWLL
1VtG1jftUIR4Cokst8P3yZtrzUtWDYoyxvqOlIEntB62zL43v/SOeJRsEdYyPkaS
ymi3gNF5FWL2q2EGzexi50LgItmpFpW9b/Izy6/O8H3ckXS9aJEaw61jsmecnt3c
5FYeJPVt8FbS96EQ3tfJI8ZH2VFwCTd0TZXusieT7i272UI8IZKgSxJJ5jgJckJ1
dEUItkBu93D4X992PReemZDaWpOqbub4pRkn/E9s7fkKUbwolwFkWIYBgRY3Yb0Y
vpYZ5LdW64EOE+zx+y+Tq5KIxjjTChiQG+nOoJKj8QAFYzVW/Y0MMlTrP2uBxRej
kWivyo2Op1bMPc9Ck/gA/tYGqnhij7SWJ408MOuFP0EPZAbtHWXXCL+fjzLWyIVu
y704JWt6KjZhUF7rtIn5AqdNCMJXhrrR0nXheTW8qyXwYtzwxvJwGNBDd0eIzRvZ
xlt7mXewBm24X+9OkiN8iwtyglhtF5Qd5v7IjNOPyecwSJ/DCAXSg9VKew9/0IlK
5aBf7BMHyuIbLNBGamX4gaoFHxOOc3B0fX+THNIWarqZzm6fUVaZGfUILP4bX4xR
iLxXEbb+GOUfEL8/QD+scBbaFVG8h26SIDAZzzAheWKi4byfpiRzBBLIuE2iW5hE
t4C2EkYs/7lnHYNscmF8HKXYYQYWEtV4H82yboHNUWUigxepENEHfsZClNopB3lY
XbHHanjzANAsHhP7WzPpKDn70zBXHPNdRmoZrK479IN1ELWgyvY5NHxk1cb9QGpD
IX2WGu87R/J8fCw15KH34jdrHAlnLXDptyRs2TKt89rjxqnAlMxoKg9KV8h4436W
0i3/LUxIcSD0igydMHZnaFoH3Ig/mAWAujkkAjGRtcc6/bdnWvalzS/hqSdng/6L
sAgQ+wrl+GVnrkK9ZBlWx4T2ClU2T7WRfA2qkV9mrPpRhmOJq3Ycrk+Na4/kpyqW
CRr824BWab0qZd+QmoouTcnHRL9CaWqRp0fZqc4ZpnQ4cLCsdN1SDrjpUTsqdTXa
k/0IQJU+jMa1fSacy2pMoa9/4oQym/26EfLJmDzkCL0Oy1u5NmsyEdBMwSbhkjV9
vvYkFgk4PVah3ePlQJK6C3psSPdNkYanBZnagURshhs8JgS4BBt0ik9Qxm6c6mAm
dZz/I80wCiYXAdE3CjvWxzciAov8VgDCinH2y2PdaHOHOA9y1JfBHUZZE+E9g1Tu
ncTDJIxh20AUZTHqvkAisJedIk3MDfPzB0BWviWF5tP0disrl7MLIYEGzdpP7/6W
xAq3fJc+IyxCBZGNmkqNoODVJpK4Rq0B+0qF2XXip07F5Olufrdn4WcH3zWHY8TT
aoIeSY7hksHYR6k4dV1e7ywyl0mYWpK7BKWAggbWc7S9wumeK/Y4tZeHN2tOI9+x
xzIo3SKK3tokSd0Vjl20h0JBvaIYO+HN4ZJwX7eueu0lXC+RrDmlC/4nIbCWyTJE
nq1GwWcVT2LOfoSWQs22ZgONJiDFmde2DkHgPmjKEoEmh4xIEnWht+/DDsJEHHSj
nPd0oGfVjMEWdJ00NqJjcGq9LApeV9AqHMLW53q80LmfvPeXcXzneG1OCW/B2NqD
ySVYuliw0z78ePdlj6kYQDyspwT2aQ6OFdiwyvFkdq2rbKA2hGFfDN3acQ9SB2R6
h2iSE0qrBLvOPg4JAncUQd6Z1wA1TXX2qwiwS6kNplWUUmPBiYWotRUSfUopgY7B
Tm6Z3LRRQDVM2rVhteimqPm1WBiCWtEajGu9tZZPQXHXdQ44JHvOyylJFIwWQPZT
i6RTZOo3LnGueC/Vqc6ZHOPUOD6MtgTnNQcuT+ROXt2GGZ0YH3DiGkJOTb6m7J0c
dYcVUsTr0No7NZk6NXIaMEwQgm0A8oRCiKu/rwcruRcCq2yihQ8WDfnKGo9t3F0+
ieUTYjWKjFET3WOAgUsVunzdadWCbcC7azNMp5mheUJ63LSSpdfeWlIc7NRJWylh
pqJ9F1JST6RI4BxveLy0054FnzlnGzliH6L5mNk/xo1vYeHmnQitceN16URtDet1
MF6VrLYlixZW/5+zdBv27UzjmKUX7aaI8OXmrWIu9zgIZo3KR+nKf/YE95YWd6DD
oGLdCbNTpVVgjeS7YC7+o/aELxX+W2NgtZWLZsF5k8rvoAB5QM4WEZMQBFj4/ZSS
jmw/JrL73PKAOSimlmLvjDLeYNZ0F3nn40ieaWOgIHS1a+qpBwPPwiOj1TtPpsiF
1eKgchJay0O9JJd4h+bGytX+CbkNNKQWLoNx+X70J5glhs6KEzQbI0oDNDG3Nkyh
NLdV7VVZyufMwgg9zx4bTovkZeBHeGz5ewYfv8gru5MLMsFvLf3eTOXNM68pQSeg
AXaAsmGt/vnDQChC59VLLgq3F1DnO6nEiyo6XBNJYJ8HPLVGuu8KQHDcTsuTP+hT
va+rbjk8Fq7GvrVA5355d1L9uwBBAavJr9ATC2i2rzVeEUGBg6POrMxuJR7BqCqO
5+ZVTLSPflyLtJRHOV/0J/0Ri4cNJ4PolxSJAdFb2YJxie+975Nd7UUjDUmg26tN
SeJMZzwIv3Pf7GxTLM/ZLY6BRa3wRorU44HdGlpx5gzPnfHAb2rJqlmGMRnyD55I
SpGvqm3XL6gOhAbWG6ej+MpUYEHnjdKOdWGil/5tlzHpNH5gMfNx/5zH7W9dr9bN
tqIsZtqeE1lqsPD+XbnzmJkVIXcDc9i1gweJUPrZN8wEwMEOuVbcyFYf0v6SBvJK
ptYe5uEQu7cdFmYUUu6V0giEuw683xNm23d2HKOv3POzzksV0eQdE4aUgTlyBuvL
gVhvyBfJRRa1kUX9B+gzASN7/jJ9c7xol5JfLei9/IRUJcfTH/T/Am+8kGEHW1Wb
+m3n/JwKXkDzknNKzew7Fiy7j0fau09gHLARxqZM/G26rZHySWv7cMUaqci5Z9ps
E63cvike0jIPmYNmRfMoOxMA2ELeOZtlRyIYdkHvp4IwaHGKsdaQqIYDbNy38e7q
06/YMDlxgNkKAWZxoXP7hhkpWXqzeyE/ewc0HIsU70mUHwahkmrEMaxL+LKbl+yM
kWbsaEHSGvGweBO9JnF+gugn6ky2HVVcNQEfhAstLkJaCoQeBMuDjtEve/83v/XQ
/2485ZhF+XXlgxwSaTCwp3snetjnY+/NSp3lEbN2g/m6VmWkCvO1IzSVCgpGhq7r
amutTHfo/MSo8TgIXBqlMj5X6yHtT87abyzA7bCFxXl+/WxK/4GPxYWR8r8FzI4h
8v3A6RyiqZAo8ayHNFiRuBPSkbo7wOMSfUDIpUSTVO2PV6w58+79OEU0qGYeBY7l
RkS2HUpMI6gPtVPfKDg+I8+SUuyyxTptClTBtvU1dxKw9QaE+6Yy8Git61eD5S70
a4WWWJTA3etaTzdqx3R6hva2Uptrb/bjcS50hW7x/hKpPvGXwTy7rHYwnBdbRccG
LcXlWXjyRiGKXQcY1bpsSwCMfpHqDcG/G7VkeF0F5tq1B6S2vpmBlWEMYfjgWaR1
hWclN84gpCAqRGcbNHTtDTZ+lqBorQSvuYUYYyQkxKsw+aeDVpHyEn44ZyB0NJCs
qJsAvo8TBHDJECxUot5OXN7n/RcV7uHBPjltgkc4Lo/11GsoHAPSbGE4M34Yg8wF
n6Ea/2Rfh6ltYH2XHVkKit7oeXLT03M82W1YVgXqkAnAYXRqGQXp2llWo0hMv7G6
WHx4SuOnfztpmmN4BLV6HtpUHfcpRAkGV1lb3R1swbwV6bk+xuSxrjKlPF2g8bGB
WmVQwdaVhbOjR058m8T8BczItm8sPjp0r2H8zAwk8MIBRUww3lROrxFuu4iFcWaj
0wwGY2IjJkoh/PlW9vDcnmgAYQOaOnQOMX32aSQsqPz2jMMIn3hIzUMbD5IdYWJb
sOUc1a075mqKKCasWviN94FEkqE6rxU2ELSdA+/fffT/MR/dO8f+SPTabWHYgNHy
FL3sJ1WDrrWTXfrmijQx+g5dKipKIStsQjpTqGI5+oPA2dNp4eOnXGJxao7yHQS9
SJKqpaiMf4xcBVdFYZlpURhyerC0uitPtX5QR/PoyMOm/TlXeVrfjeP+00AuYS2q
mA5/XvwZNIvGFZoFy42XIChzQPiuWfUeHhuB2153fNIEmuH9ZdRtz77jQVXzvZtp
hEgvPg8jg6fnuEUgBD5bc3Dc/jepxyZAt6HC8+uYq82YE8bpwb52K0ZVMPWdlzu+
+UcbILRWxiuhGoBrHmMsQcrEf1OjxbnrPKnhK+V4DNvLBocRmeYxHdRgjVoyKlvg
ft/7qsP5/idbopCB13xBPNW+w2lPa18ccWHO2B5vBNMyhBLecQU1phA5ejmzksU2
mmnlZM2A5zwuAPW8XfZP7OedXZ4PGTKLcYeb3qjE8dvtGPE0aI6Q7xv7YhWxYf8g
O0qrbLq3P1WaXp7xmvwHtnbE8RmFMh3JjXj+V4M5+07of7AB/9j0kHiZWv/cnSc+
xNfPw6Bnw4e6vddPoyqoC9QcgNB5VuBEqb+b7iyV3F/9GR0qOtO8t1OMKiQqcCJ/
paARajAM/OSyX55qurTLGfmXUjIFnNpEn7yoUjh14JG56G69GTEAuhzIbyDKOH/x
UoypFG/xuyfCGC4fnaiEK5kiXdnUp6/4diXYF9hVJDaftWRWnYeQDbP0AdUwoXcK
tcJaWaSN0V2FCTlD/JM+TggVsf3qwTtG+RYYQosVuffJSbuX/q6Gn2Rf0cB7WP/K
jJ/lycR2L4UmUUbzZObZ6fLuRP/o11QFm2WEHPiADhSjhNwvpTXi568tes1SQl7Y
2jo5VrdKDu5bHODFAR8uWSWhcxiLvKd1IGIeonCSM8+Ch2nFZMwZPYYJ3zDteJbR
w7d1aymM/M299xD9LUKk5FH2eT8uxfPq0B+VAgDgerEHtbqDVHQFpoq252bhCpEU
UJXkNHOq64L1OlA7THdYIen7T4HUPVBrT7jPlkuZbzeNeE5TvpW//lRXHm1HRDm0
swsIO51ljZybQhZnWmvEd8RuWruFaqRmNen5awC52DWM9ZvFFcIfqgA9BvxuJG5u
quADWIJWAi3gyp9QkVcJtI6u92vNAWcNknU3euZnycgimubB1C0qDs6lZO8Bf1Fh
c7YbwdcLydA9hsvIacakalNaxmE1z5vTF72hP56LvLu6VWbb0Yz7Oph5mTAI15U2
3EPZnK+rKYSHpMz6gGqY0EacDYAwrYHBz4RppsZFy2V2HDyoAdaotHUVbYLOo61j
oOksmy7Qfv6Vfw/QIY7vync5b51RYeLoHuC95a3FQ4DMXlLeT8ChL9+hwQMFNkJx
I9o4k5+WFkHEYx6Rc1HUcqsmB3z6ksr1fQzztQU7ganMDWH3qmyH3nly0vbAWflW
a9kwSnosjgUdWQubA7KKxzTaO2SBBxHQq0sRscIiM5n6L31EmLfyCLHkwFt0AurE
6f0FNw9l04o/mnXLN7SdDdc163QothPlU3tziNyIXnUgr7icUC0/DqReWoKmLQlW
SzDNh0QRcFlv6cTW41497cZsGr1ggpLnODUjwuR0lluIxoo4c+9dEdOd8FYghF2v
scSM594+tGxrTG5wEiiEElyn7YlNOIFn8HQTJ/+WPFaHH7eSMOUwtCmpersxhYPf
swUQR9/L7TmAjLcv/SZ4/RVNHEFD+fR6ZkNpInU4xa78rmhS5MKHkabNapquu8Tt
S2Nfc+GIuApU2Uvhp8PXxZXi4rQgfUQixzYLYr/xUFGfsxo7JHrK2iZKR1YccdBU
MVCwYBKqgFDn56Yi7PTAcPpWA69FrHjNiLyLe/HjBL764K9/l1dYdyWGdODaSa6n
EgaOeOqtyJCSFkby3VEntNb/X18ED9pxuxNo74ab+7MhtlVnMf/AMVZqIzE45rRW
fJWwrE+Cz9mqUBKjT6c86vgUyB8g6NoheuCeG3gW789cQiS5GJVst0xT1/D2ZvTl
cTu5rOE1eNa3ODImhv88r9HG1POGScvZ00PgeHzIK4aDraPlUGjEwvkelxpzvX8V
3TUSieh4WvVu2/NSe8qO+Mh9MywFkXqsmwCy32h9qBXi0UUZrdd3h9WVvdSFaGfw
EDvRhRGbYB7MdNx45+pZ20eVNsizMM+getjiqFjH7hAPpPZXQttoHIf+JGQ4amjv
6sEgXPn2ZoPltYHsPgo6h+6ZGfoqfyMF66jCbwVGVFIEc9/8mnhEQD8QAsOQQBhi
9X4qaP7alp39tqGdtQAbgNbpHzlbQS2uczaf+oQWhmNKNDuE2bSflEGO/9ceQxEg
/4mO6LCI5iZ4/ONomg+ZxcZWMcdiXHzqPV1bzfH6/8TIabhPgxxQ3Zz+EAxJWerz
4j2UDFEk/ElTsIkY2q1vJHZWN8Of+1QQZ6YmYTqW9UTNxzWdfVlu1Fh2uNchJxKp
idG0SGfIsksslSihX6bAiIgivK5XXZJggoXQLdfheZYSc6syvdfxBB/amU4KdPC5
C2ei99neMf7hYgGwl2zt0fOnCPv963dH/fgBIJafoJQAtzUb33Lf8Cb/piVxFaxk
4WWHi06A3VC0QKPWFSpGOzJO/ZG93rB6eEqZ1nqJxZCSZitwj02P7E8ygVz1IO1w
BpIO8j3jQMBx9iuomEOFOjA2IKvuKg5vC40a1s6JeaADotsCqVBeUFNf2A0+XHAY
7JBYN98kn9/wJnQlUYgCuvjI/0PSCG6xjDerz9YGXlxPXBfVpYy3coadIBl//Nmv
7DdR8GTPPfBh/NQcgDrpihAQp7nR3oZyd1XVOsKBM5A8OAzTd0KqB+VohjPNGMTm
ff3kBOnxS355f9fmf9NB62xItdTeS3vA3Q45W740Q+qWkMx4nRJqN4lY1qZR2lqH
lBcc1Uh+Gq4Yfl+GNn8yYo7hxKW19yu/k6nE9MSscWi2dLXSwkDMB2bq2wS7KElm
BIwiNweWVoJ915w7Zmi2jwJctCiWV26YOaPQjW1M9EfxXY18DLOw72MRmkx7O0/h
wpNl/loc2hNL4U1l5Sxf/kVJJviwyqi+P8SQWSBKIIgzM/hrYENdPzp6xIvXh6Mj
/hEpOuhZzrDbOK1QlEB3cEPuWqCPmzLxwTL+L0VQ4WMjnvhN/BywYq8TgoVAe1/O
co9Bt4Uez4CU9xoNhwOD2qxorAtOejqplDylX8+Eb6/j2RRq8bK/HyrfLU3Qzmsm
CN+agCfO0zFcKAR68G+ye2oXyLYLuFQlGsNWltsgUuk+sywcFyT6ui1dOzVtSzw0
Ep0GZAl41ZstKK6nxQogcmERDYW7/Qnw3DdUvvk1fDEC2rUY7J20ldFr47Idvst1
l1g8iQLv0ymqyAtdFEjpdg4OchOBTRDprzKKr66JHDx1m98cK2giPYkm/8Dq1dVW
rgo3EsO+9KJkYucX7Wk+D3S/SZWTKrmnxbGKmZmomRgPploZhcZtjoihMMOszoXM
IosRgA718a06zslmWvgsk4srYwCbXnDzvY7R781bftJimfa7qgYRzgn7hRosnnYM
67aiqpPS+vYEOFDKSOOukPGlSWTI9AboCrsIKw4SMyih2p0pdr9vebN1P8Feku4i
zPDDkWAQWBjwSpxS/TrMSKleEaWytRy+MoeWamIeRd7LIBVt0NsNqKkYG+UPG8HJ
BdvU7T6+6/vG9IhiBdTdmn/KJwd2AhsQkysbMnH0/hF0C+qzX3ohnwMdG+MaDJp+
OVGyldv7ZA0XCcIvjmDjAKVB/RdUwcJycxbAMQ8c+oYxVJP5u4Uas6avRtOQwFnz
lPHXl/NKJAsW5W4QrENo3Z6WyrYl2yktQEUt1cBcAFPjAymY1LGCanqrBw/zzCyX
D3iJ8t8XShoCesK6g0plYcHyXgVwZXzrtbSmwkiCpxIo7SEkC1cfB3CF6Xzgqlh8
0jLKIbX/nbqUnGDvHuzn4h7oTjfGcZFXa9CqrldEQFe6bTGgxGxoS5tShatn0Dzd
CLkcSA2ndVJx5TnfFUQQUg/ouh8gTnI2H8i7E1sXKBSnbNNVxCKYjf2Wf7hUQnTC
W0KAwHHSiafkWFxmtWJ3MaKxpYn+gCl5Ec7LSydANCvo3HNVDoQrn/vsnAEoL9Xj
z5ZQJHISLG1ot9HLNsv+LDQRh81CaBb15Y9aZxUyvg0W2pepZXDh8z99DSnHwyd0
fsagBhgEM1xcG31dyXxlrRYnxbMPTiq0ulsEeR+bc/PBv6A83eQ93bIuiSsdbeX4
wGFldLe26E2Lu7geUWgUjXa9ERV5+t+iZo/b1RoXBLaCOIjuuX1n6xIhbnbg4I0Q
JYPDAnIkTCPWlq7kx4wbe+X/zgpaiHD6kPDTyGro6PZmzZHsIQwTbgKzoTrr1zQ1
clBQ71tFyuTvKGnbH1VaVLIIRu5pNeWydTmt7DzCWvKV4alnbOQhnsExA/4/4thN
NmKPTyb9TzRTaI3KHvvJCZQ8H4rsdYSRx4sXPDUFUQLhGI26WdC1jDVB+V/DldYP
jKxMCFOF7BnhMOAfzcEBb3h3S4wAQpFK4H+Wj1tvtvjkAagf+L48SLJkKf2qRSrK
MWsPrkZIMw7dIwBFiNfh3xK9gBJisbIcK0Vf+EL5SR3hYJS1fI5oVXj16dB+YvbI
J1JpDvOaxowTwQ5fW7C8ZnogBKMzay1yg+OPcsi3yo2tOQYdzJ1rihRHDfCVGUez
ebvnRPNTvyZCq6ciK1kEDZwISZXZGQeOwDoSuqA5/w3xTisi8V4NZeTjDhz22ybo
klOT2x2HSLuna/BWe4DdwYNaaHtqPPOavv2qdCAeLg81/AavuqdcYwmme4Sp/wpc
+JL1WVULW8Gq+Vo2Hg85RoveV9UtgiepiK2NiZnCSM5Htr2JxiTZ1zo0smhU129n
n5x117w4C0AYwOFVH93pWH5kvp0BR/cwoBqzQYorON2IYPMAgXYnlkfDidClo6/s
e9HP7X8GvDTdz8dgErhd/G0Pg2EIT5DF+ItLwnEbvXeMY4Uk5BEyf5CxYSkjQl/u
BN/R94fpArRDt9MVwAVKzGp+CfeNHs3G7wj0QxaWxAXc/GDdOj9WiynHIFfLhWqW
4tZsqEVFnYrzzr/xWXzav+ssc2u1KOUJiOwVoSWNPQo15LTmAGHeSYtf9FS8tffV
VR4NQwSBo3MgrLtnBNsi1zob084Ij8QFKzgAZHb9cIiTRb4s8INYDO9IHUNoFYBN
pjdaPoJ3bAgU6eet+hlPoKC1hR/2crhmWJxY76HrSE3qhkNm862vOu++FPMl4GJf
T2X3zrtduEA/FKVTmB0DmDDW8bHDk6yQx52F0PLgw31Bxr7kHuaimkgr9RMHQNem
uj7+Smbtt6XftLdk57Tbam41TR10GlAuTQvrBQJpxejuSYzqrW/FKjEwpsllE8D/
e09MOR7AU0ac/n8MRDQpCmBvlw8ureb8NKKV35j2rgfAe38v3biJ44RzPRSFvKTJ
RIPe24NfhZ3zLA6L9NR/k9OKFPBkwuhF4o8uW5qHXgn+CxAXkvpSPBmJtwxHPWZF
OnekhG7foW+PBauSNgv07suJFJUD7gtlAHJ81qcLl96jtCZVTdIKf3SlmNaNu8nl
wVleyejm6Yyn4vSnItQ8SNV6Y6T8GEI5v4YZiYnOx4VhH/UtJmCW3gm68bpNIwGa
VN2Q2LQzXS+D0nizaNA8OCKWvxWGFo20FHsgy/QaWyQYf/2mv3PYf2gkSGjpsYFJ
ZycxEHMWGwxyFB8yjaOfD78z8QGGSnAhFwQKzzTJK2ZmoF++1r83LGUnElTv2DMA
C6qH3octTI+SGBkgBoYChtkJu0Yo5E2jf4bAwgmqUNC86DiZK+aW3bYdQz9m2Dhu
XqZul1C1ryBul10zfEJBGDrQu6M1kcrUbHGoORjAU/hAC+fDubU0BC2GtfTZJB7K
ySPNFJ+N9u9wpMKTopmGIiY481COnAKGPvdN8MIZsHpVhXnSknup57t0WlHuw7Dw
+0UWiHFGyrJRey6E8Q+sLZEGeCUkn6s+G5M3h7n2KxlM5VDtCFJzU+phFllM9Q/O
Yo2Vwo6bzGlWJHXUAmuxr9VVCHivHEtU8xyhucRUu1L7o0tbQkZGG2QB0ug02VVO
B70QRamew5d3KmPDIYZnDzhsVNTiJv6+/4cmVw5h9Gi0KgGgpunX+qIQiPt3ae1A
KTbcMeFx7gKbNYK2gjX8DFRINn3fmrTEe5+gHL1zFcyk8NkyzUb244x08d1cvPvq
Lx9MdmVpFUCMpnyvvd///ZOF1j6OlNUI+ssE/Smb0sJPt8BF2xHSpQKCpIHujL4p
MGIh7kk/H3SkMC9kPa1XQ4sPRjbTUhutQ5ZRGPVrNYug9MGeFul2qadZcCL1I9m5
C9RmoQQfNkBdbY3J2c2rqNhXAqHlPUIz9prEN1KmEg8pnFLWO2qexXoMrvbxAXku
KKVpMO8bLbvlAZAofcbCjmdzEZMz0JmluEunTcK+bSh/1ImNa74bO/gptLm6e0Te
FVzusaMlPfKlFB1yM821SyP2EZbcCsOElvdMlvskxIhCndYiEQBbkdZPHWtmKl9f
ijPAuz5z992TNHkWqHT5+bPALDTuSpn9bzy0zCQE21fVwL8cCdfMi5EsaReU9pQK
AO5884HjOhtVJP9K2QJQBtjiwaDujFHUf+Lc32ow/2pNJQ4ajpD37aBf4Ho8g8gE
CwH4nI6FH9DUB1hy/T5hcLkKyP5CVNciIx+cYu96nTYzWCOPnhHdoZjTwOikelXu
vQc+wuQZXPQRF04TdeaYqR0cW5yBQCD0PsCbXfwVNFSC/ybIFlA8Mfk4uEOwKQ5Z
hhXGc79jSME4j181omhveTaDs/BJuFB8m5tBs2+jeqVMCpC2WK7oxwhQSBCDdz/j
qpQRBEumN2hTm0MgNdnyGpa5kesFxLK3DulsEN9H1tpwYK75NR04Q1GacmUTQl22
CDvpeEJJ7MIFoVed9u/2sTWAxB+9120GFdJdz0fLl6zghVgJPkkUy7FO7/qu38Wt
uvr3P7u0GeRR8I6b0fIFEgBfMQ8fm+gRq2pNS8m1WAGCazWLe/xm0krWDTyW/B8y
KSgZosH/m7xJswSq8IwZV83YAX+ZiOx6rUmO39pnxTXvIHLNdljwjqZ3cE4ciYta
zO4S9jEHF0WMxToJoRC/zSoqezUWu+24d7eRK3+eT3mQvfJeGQo1l/AzFLO16UMu
QDHIPa3EFl0vH9rLPB2Q9zzH8mVM8z4/KVA9IQ3K7cBHVx1P1g4R156EIOsDg5jK
Dl/Oe8xhm5LOnV/LsKdHX5ZB3oYutjWFfkCT1Xjx/Q17Wpb3N5q+5zjKTRP4xkGb
ZKGNrmTf4iBbbnoAMbAv7Jghh7W7xO8CLA/ianeoTA4LE8WDwxRNUwV3qD+abvXJ
xUAPhT6L/YbwvfFfBBEUZuNm7XkbIYnQC8ewE/tO3N7zm3uAkAMr3kH8Qs2MVMqI
figOlGB2sbQmDDMStSvJy187wB72UCSZZpXkIRgvv8VU2ESQDGpkG4X3C08C0+/E
4PXim1vFNfiP3H9EmpcS1mJgWYc/S3/MifxN9W9xROqoOYx3wANleezTakLH5RZz
KOn/X2eIzUK4VzEjo3R3GJO04JI82IrZfWX5Cb2lGbRE4y7Da78EX9B80bhgje2v
2thh4JwAbY9QkVgIYKTee4Tr6raonT8QK7VtH5/CmDwLg4kn5IOYPQG8UrtEyDUA
P9QNAmVh6H3Ptc/wUUc1DuH2zUWAdrwMmiKQ3HmgVLIlxFGxU4pCEDBLO6TmTNVP
1ozjW46suoFS8NzPkSG77WAqQH7J6zun6ydldBmUfFIYOBvIgr0aVQFXqaIxc3Lt
HGn3poDM94EBPrNQCrvii8ul9XitUuHCUSJ8+eSlS05ad3Izl36EG4a9HrZmFAYH
iEfmgYkobINj32sOwdR0f8KOAHvXPrijsbSrS7xgOTtbwJEusPjOd49UfSRxwLp6
0rNkeYnZX0U6U1Lcd/aQwDazbOeevcoKpxFNb69tkgZg3lyJy1xpfGl7iA13BZ83
mrrkir58WyVb9Tz3NJoxDBAmqLuyvblGJMFAzXFObSLvlfw95u/Mt5teaza4qVOJ
dN4gT2rP4WnCW8L3BUnuxsI+T6Vaa/racUWQJt9LI9JIp1QOaMJl9gp6j0nq+ymD
gA/xQOlQHlSLWiFMq9zhMVynIxVCfmFI6M8T0cXSjqVdZnPlHcLFuGndLY0tfC29
tm4RzAgqyU2d5JUUz+fsuV4uxWyHKa4Ib7UUftu3CDydxYamiMUy4fkTDEwqhRZr
zhWmTh/lHeH0N109UTMBbM3sWTDSXrjCvypKD0QXAucDGKq/xKVUECSblyd0lNdt
eR4+fPNsuMy/hE6Re1GndwVjV+8tJcMOJeMken1zl0QVpbE6sft4OluHFxcQ6OKX
8TC5NCCKeileuvyZlb8Z0r2FzyVvUYAgFVf877nTd1ePSVfvEkenejWM1ZEySXUi
PRb66n5+wafZI8GUGHWb0o8OtxxvdmTrpMDySE0SCfCul7zGiGiX/MDaKHb5pVku
WTEo5O/Pp+u4Ik9gb7YkXmcfoOi0KTtxVaRTbeDFWdbm5WiVT41eKgrDZ9R1qHIB
siSX3YSvuPg0xrDCbE4CioVLxlq+CUPGyznnz41ft8u7tltZYL/jOhZdSyO8Gy1+
99FRkiA09wC/q0foHUqdzKEQ/fFDaoW8i8sJXcYxQrxuJInBBercLCSO0DZBfFnb
XvFk5yEjsLcoZhtES3vEQCXdx5NvtHBNfjrQYNjR5XZqx0wUl9JpmHd5qLtXHlbz
EpXgFq/hUZrJUy3BkHrEfDraQf7do9a7kJpi3eD/D3G/qi8QTaqm37y2R7HhunQj
h4qdMQwc5/GYQF0nuFYegxkiUZo6XMPenJnIFvGVG/xE/ycqWdGamws+HMutnO5j
5DvcE9KIveuuYpiqwqPXT8jqH5JeK3omN1kaiI/n/wvYQ13zZTfOIabE0JqSlJFX
HCZrToWT98k10obh26aBMTa7YUFbviYt3a7Dgu3qqBHAfvkiT06+LK62/JM0ixyG
tEGBS3aZ331oWKipAl27SOBhuaBf2GB0Gx45FvmIfoSA/KPmUIdL2YeQaGrwhnNJ
brR/dmlzowBrobS07xkNaKfEf39PcD3xHTOggZJRYiY0IV0p4/0mGq5oT+zD8Wfr
jIK1UXLsFjmJjkoVyG/nhGCglGojKjzDehwJX0UR0Fj9Ru7Z/k9xfQU0HfnOnkLL
yJjDyl18++ETiaVUxsTkNnfBROmRb4IQTWR0+ObUXAt9HB3HlnhjwPm5HiAZ36S/
n2zHiD7sKoc7OWJtNXtgIw3SF3nyFf3F+7+k2ga+kyyxQh2Zv6EeeCGoG0dLaJ/F
NfveSu/3Mnpsz1Pjj+8RuyQxsZn64Y/MAsSSvI7DQhZ3cpsUnePWQUzeaf+TUW1O
gaiyK6y7Suqhx8XQSv3ZhwErncn9SU3WgxYVUVBWlxul/jMAVrgPuVICYdouvCam
GZcKqR43m1aNi2UqcC4zQfDIetuugU7LFp2wVzQXKgr2gzAJV4PrKtQTmxZgcThG
PuvVTTnSCmyQWNcGTF7ZfhT7lliaVBoJh+10r1Z0e0RfMXrWI3QmSUsA//PRLO1Z
Lv0CY+N83uLfZwpumZpkYXGF2fW6zeUCVOgZ3fJnkB27uwmZ1qHeoOyN1YoU6kRk
CwO/AZ5lzTMh9EHZcdqT7eey8gurIQeSFFX3oOlmosTNKMP4bQqgIKOZIenkjLvk
Rler7X2MiW97AWfoAbL+toy2oID7VKc97aptCtI8EJKFY7+0Pw9Ps0MRYodQXkN5
PyFmRMv2nZqbH35vNrrd3jjqaRDI4IMvovW5PWYuet8mpxYkF6wQ1PTV6tS9br0U
yj2h85XQJVaMAy6yO1OigBIaSHpWdgeZhAaC+YciAh1Qgh5HDsTaF2VmgRs1z1Wr
cTZPkrnRSph40cmufnhf1hN3n0CR/5CARtFLh/Ajg8CVJBLNAreDF+qYv+PAGY+L
S7VYLTbHklems8JEL00rbag8o0YHdNbb7UP+2WG55YpJ9/IklthfFp9CaxdMwIzG
l9M+JWv7+hNDz0boVOXJvaADgT9AxZWuxlAqFEK5ZldHnl9SLCEVXe8h2DbVY5FZ
VcJ5mBKdfCwkgIa3TZdA/u8tT5glDsLh+wf5dN/T1Nc=
`protect END_PROTECTED
