`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0y7Ajj6fC4ByNII1lLGWhk4WBAIzNcEwE+TcIB8vjlYpM0om+LqCAdQYSs4azYTT
5EodOCr96XtKNCY8ToClFsKN83sRyZARi399ZQBKrXwXzvKWOALMbhYxYek5sMhc
VQ6e/cii4BWyWqFn+kRO6liP/LgaPIx6MUMlfRRKUMY=
`protect END_PROTECTED
