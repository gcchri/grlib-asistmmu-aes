`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
So25MUZNAYtUTo38G/HzSLZBC+YQjOWGzZOSalsNQvZORBtRTnht1yM4DWnwKY43
5LnbNrUigME4W93t9b47Pq5K9p01l2sU+0oSyGrvpG46fcFPqKl5AtuOC65tt8KW
1cHJnzRieynH5lmZwyORT9+EdJL6KXL5DB3jI2WS7khZ+EJ660sqgGm3eW9M3dvZ
kA9Pdgr7jl2g7RrIJ3TzNEnK4DsulaSh/pLbaJPMQLMBapoGV00JnH1gQUiqyQSB
hK1QekCZtB9psCLUkgU9KUZ/9qUSHG2vr0FpcZn5yL1Z3S5CmLz6Na77GMKpGKld
d24I18ARhzfpO4974wwOW537d/9w8AJzhBLa91CREAYJ21axh6SRTPIe/LmMxK5Y
6ica3fXMAdoWK/V1tZ2UXNT/zSER0q0gIyedt8I3PWUqP7I5YHFxNyot770nOeIZ
KOfrztJyT/amax8uHin9OCR8kIalfaYDSdo+4F+mX/mEPUTes17ikyufjw+MK63a
ivig6zLe1oretqw/OalIjYii4OOH4/poDlU0HZMtd6M=
`protect END_PROTECTED
