`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2rRriSbObJDoKT7zXVloSidiF6sZMg6UGKF/+QrJxv1wfpbla4QXj4S/cr7Lo+W
Mvcvz+u3XNpyeYhyCecLgobdSGbFOjlBLNhGHCEpsIcUTJuXeWjbyJUohoT3S9Fs
TgoCqnUhBpdkEYmkBX9+gl0Omxo0huG/PtXH568ZSKb7ZrKNE8y9Unikt+TZQoxs
oAfqRdX0GRndvWXA47ljTGXDlyi2SmbbxjCx5Qh2oG1Og/NJIBlJ8GgoRuM7GEF0
ioF3HpsmuG/QSaI4qiiN6/FQbJpSud4h1GOFo7mYnJzcHripaHxBL3ooueN/wDOr
9ORu80ja1Y94aTbu206hnxl3FI/21rSv99PQqEWulHGCCX46UTfyhvgCTLLqJRIa
dKT1eQn5dkqj9LYDaF7lY0ZIdMWo0eqFUzhU486YW4hQCTb0Gj8OsnsDoAhXbtca
`protect END_PROTECTED
