`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AQb6ZOMCV9ncjonbSMXui+ciyHYaRG8Dv/VrsClccwRQacWMfNdIMYXhG0istY8n
NH54+zRKA4VZouYO+LJFPcQ52i/MpS7QYYxSAORVK/rIuChF2zQ6SHwDCkuBBeGw
Gk8Wgx3Czt1y6cmQYvUNOfcQOSW2USJFCfoqKMlNpk1t2oCUPUMWcVVEcVZT1XP+
UKZUXlfQMRL8EhaFE2xptPYPdmKoSuJoNV5k8Q2O2H7aKt2DiCUqjRj0AF9C319N
67FkL0F327vgNH+4pw35PJ9yhgezLk8XSaanbjtnMEjfrORu9AXdvkNoiino3scG
E2tkKs0RAn0bCbkQ2bda75rXipUIuDd90QWBfoM/7wkSxrVXReg82Tfgjf/id9kk
k4zVA3BUZKKTrbw3+wLcmhdg1PtajxX5IZpZg0kUwNYq4H3cNgAvgKH71gLPoble
x3CtWffE1QyC98uALhNizu/mWR6rjqi0TlQzp8tLxc0+wuhfXFzqA/7MvFc48pyL
ghxzJv6aVUsHSC70IbVo3DsFOjx73FL7B1OXDJ2v0f3UceuBY4jy2IM0ItLD3/By
YrGs65B/Z4ir7aKlotnF2N55YuvcB2kQJUMr6NmMko5p24xNRv2buDt3IdsYP4W1
UexPYwPHPyxgOe7J8GYq7EjvyI6z0L9YZ8UaOzPCp9b6W2/z91P/9osGy3zHDyNp
4Gd7d3oLYER4XZABjzSoEegx161913n0VvZ5aT4YxwP/Qj8SJcjx+o5bySmxDiAX
UeR5HwoI3wePONY6l4YNo2SG9qVf4pjhHxQrk77kTbKHRlZUa27MFh/tahql4sNC
JTtVQqEEs6+/ZV7ky6NSdFgEhvXcMIEShz1uhpQxwJW+rYV2IStrhM8cNLeLEqGY
BOMFfPDqUUD2UwBt48UZQYMcpUzvgXVaJCJuJHj6lHK+HFrQIhLY0H/Xu56SLirC
jB7PyHcMFOLC1MQ5p2qPsTE0uUQXlDh/MCRcZZq4XSyWKIp91Z5rDucW9Gk01D2c
AmP1fELXZxI63zEvzijUMJlfPtHN37WHvjivs1A1iDbm5jfiv4PlTp6kSOiRFJpU
IaVO4AucR3hCYwK6G/UAzstV2pDxYcK3l6lHUAQsMR4pahtiCiOIGXOG3CSQ5Qq8
v6tJcDwN2KHqjxRam0wzAu3rwONG577PLHiOwdJunVV5sVbhSU8QrqTbbcuLr7E/
hoyhZ9pPXlwG9+uUCg7TRVbnJTu0OdYRIsvBzrB6bjq/dlWJFms0PVn8F0749sAw
htn1eFScnGqFcyh1LAVwQ/gv2rketMFfjwFVQwtHlucU7RGW86x+iRzOSVj+Mr/W
IKlsxtBfxTRw4UKEqnHqgHKBhQZgj6RQ1iVoSXMMtnc3+GNhJ3KRofXClEFGMiAL
+dN7iLhnbqSvovP508atZyKlm0bKH73OaQnLMvBVgbuwuMSJeCe6eD1Dv8gi1KED
Ca89QACHTwZ/EuFb5QHyV269Wx22eHm5zIzDfCmDpgoSIor/5dNCLJRZMaEZ+lTa
JNQqhp865oXqrf6gQf7+aCrCwA2z/NE7j/nbZBY69RBwizF23B+5ggRJe2H+QnmM
9iYza+Oh4l2UWDK0BuAdSDK83CFS4+ajRkavOSiJ91K59Y9JT3qB2V9NiZ8M+HAR
OKj1TRqiJ0KoYXczk3mtn0fvCMpGuewbyhoHfiQqXqFzD6m0ugq9PbC7F6WAiW69
tlC5B+xHIPd77OGi6t9hPejKOZ4bGx78u8SdsDsKaHg35SaztrZqsSxUVo8U5Nmb
WkPiOam0R/9yfLuF7U1JAVkzvNZzcaQCTOeBI9Njk4TBmefL6fzq9o9Q+QqQJp5w
6kUUsAkKrplvBbZ+4G79qJTibybYNMBJ1KSaMQiF/8cMx5zgZgFnhF+4ngjE2k8D
KxaXzP8T0lkRZhnPuYIWKJNHLtfmSfEMKO52tOqRAXJKBCuI7qoL3kh6ouKETL/N
tMsJZQICkc3KI487VYisrk0OpYay1zlR9k78MwFCBlpMDnO524tQ9htBDSeTG8/p
nj/5/DVF3SJyd77mZ7NtO/w1/rzk1tt+YVs+/KiJK751k/d+vxA0aHdLgH1Pf1Ur
bX8ke5GkSKGjfrWInZQaoQiG4y8HYL5flHVVkN8mcBIA1z9CRHO8IRt3yPuy0vkn
`protect END_PROTECTED
