`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zrpqo5ROIBRFVMt4lxEdF/0/7UAEEjEJoShZQEl6scg4E4MJIxK80I2qH4mh92Qt
RHGs8eaRFTxCj+ys9FRv6cUZACEmcr1QlZxBASAeiL24Pq8VFDhZTjYDq8BIXe0L
Ent50QG//J4rELHrogvyhEm8kYYFAXEbWztsPYhBOa3eh9VsaBghq8DeLNvs0mDi
OiY9BLkGDvL3up+FMV6vmtS8uSWtidMd2fbAqimw19c2Xh53AieIXR8hsenUIqID
AwrmtJ6YqVcK/tP6FRh63Ln18Pzh5zGuIrDJFFPY48nFxzEz3q+aN8ndKCR/x1sW
v6xmcjggWXmtv66ZRHZrbRHJ7hB33J6br+d/3wrYerLGl3Cwl2uE3Qvir+KYTuFE
`protect END_PROTECTED
