`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZGYHtqyFwTx7ze5sBdSG/6vT5tmpaaN2b32x5iw+s2igFfLWHKI3gTJ0vva+ypd
GLISTAKwqQdHN36a5GS8A9r61ELmVBbfVr7Phl2uow7fvw9fLOC8rZkfkyy62sc/
/ckdL8Jv5TbVRMsJcR7DoDsgbx3fzY6whZ2HxX8vGrCwfiumX1BbU8fdyeAEw9oS
PzYksFRQlNS/skz5eV31nz2fwCRJvB3+SW35VbCukTqPxXNVWLPm8zG7NIN3jX5k
PQVZZYJf7FP9huNHgwjEcbz75/WwhKA0DBjOLKeUL8kkOOaaTNt4e0Qh4H7Cm2dV
yhmAukyJh1KRnsuWcJRwXxjsjw/705yew+kuDULIIFpvXyELEgWMUP1tHy7+In7o
MzGXzrJv4IbwofoYGT1JY4kblHEH9uOx21vjcyhcbixw6uziY/jJAVFZJH1CJLIZ
okmMUHj9lNkWiRVxaZrJHQNn/VRv+ZnSFY6LHJkZjJo=
`protect END_PROTECTED
