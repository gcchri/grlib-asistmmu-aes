`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9xOKIG76cxyuBJ5OKsSv16nGUA9GGU1vtGcmf//krFUOAAG3PYqiQkNnX7pHBN8y
Ilx3D7tE22ijGtWXpIWwsa41w2FLN3ucwHtkYfgVSAyqFY3uU2OdczcwRuz7hu6N
C+h66BHFlsjH6Zkcp6Lgb4xNGFOcL/nJdDJx3btFlcupUPL5Ie7EHPhI0ZIbtjca
k7Fa83sDuQsnjBUu7EUJasckY12YbGSVe0uLrC8cci+qcP66GIY4/C2tvACYq5A2
Z7Yc+X0UKfVP+TmQoFBpKT9kNNGXMMuLvY/EnQ+e01DnhX8N+oTHUlG3Vq0IBF45
t23Vn2O2drx0l5p1S4BurizwDdBVnPXPO4fxAe60CExRvQT8sxFKJ8hHdu86AU5A
4ABI1jR/wfOAtMdHECl9SQyteaBbO4GsK0ql+2/X+uoi7xkmk3jLrE2w+isUXYtI
sVKLNVxO0C/tRw4Kpc8iVZFDqTEXmhgmzpKogGjeqz1zrRtMLw4Os3Ee1oEnV8xe
L1lfBZa5fbz3B4ElUqeh6NAac5jkPzi11nPDqQ7unIlxPQjJbdP/dfpbFWX7fdIF
xYwCPAHPNIYfOlwd6mJxI6to9zGG/rmLZ5FPeUkv+7aTs97DH/hvslpAGr6fyfWN
uMoUxRWnwp4KxI5/NO28hGeFXvxvm83k9tdPpaG5eCm/LSldDmxZC6g3EpMeB5s9
RGQxhvJ+Y93Tv6742/0xvn9kfFz7mr7BK8rb8Kc9/K/h75YA4vKctEKRjjIHicjA
VOv3opOKBfEoKDN64r16YWL8l8nxaql6LfnPRpHHhXfhJiKcQLkNUrYbJzjvrzPq
pwR6PWesRuEFkmf9JUaxghxpDBxOZHMlunwV3KDktPOtEYOiCajcmhENfa8v7qPf
XZd14IcxhG384t/cpq6ceXwwVV/CXhd35/rIMWsmkAo1inCub8NYJmr59mwblAyp
`protect END_PROTECTED
