`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEDUmmogofBgPEyiLLOJ9i1fcsMaIzUi+Pd47f0XKyrKFW9jfSHe/ndf+IrJDTRx
ID32aAQuJ+VrioDNKTQIUlgFTDB0Jz5MFyl+rpNoN7xbrhkpnfnExg5qjfXfjA43
O2hQYBvdyygBjJO660+lULTI8jLJn/aCElxPH+DM9Mn15kI12+ReHjh26qfdBoKN
YxUx2xLkcABSfE5MKk3kIaSkfhqSnJPEn+WL8iGgCdo5tvqZU3o6vp9kBM9fpDzB
gc5KmAhPvFYd0mJsxEq10MmqUba/qwjgr0RCXMv3JpbV7rzZxRJpI/qOHrJ6AG1D
/lKWnCYion+7L0LOulvOddPKcynw5/3I7HDhAUZzYBtg6OZQ7w8JCSwBbDOFHtF6
WfP6SuQZtf6XWJ9CaC9XjGqhIl1v7ix/m5k/PSDQfJnKuhiHoFynCnnB1pct8KZz
3y7nMWxTWDw92lh7puXpJPJApUgU9+bTDV7pEXIHdfywKmg2eog63oz1yCJNZf0p
7vzPSL6eAVLBHgF6NH1Ls8OERexzRoCb8ttzS419eezEEP19WS7vcFEX36IY1hMc
SgWw2O+ahLGmEBVaU2cZFW/zJTiKG8E6S7JxBqLHAhe0lbOrd+Ehq3e2pbqRR5Ak
4SabBeY6CkAklFdYgVXRuXXYZa2g1CQl8KZ1WKDQzw49o0S4vOjaS1+eROER8VYk
DyGGET5TyazRY59PU17ymOa77Lx0kuumDAhTADyFoJwhGsGt1AP+LquPbbiNGtg4
OJ0XgRhrL/G8o0Vga5P8a2qAgQORh7uw+lf6gu8VraOEyHzlwdyc/MioU90IzZru
L5F0Pq6KNcNTMY+9ND4wx8fdqOMdaNyiIJ8hxJsoWGdquIj04sv4y2NWBeeF5ABF
Fufyn+/P3LJQmZORs6l9LVi7KQEMZN2MgnwGIvbOqYGoemoxr9lz8UOzDudv/74W
gjoM1glR7nRKh1OL645QlYBusCA4s3m034TEYCfKaA6zwyojWVFxjHV2VVnLNVP3
QVm6xaUCxsWh78ongs1/uJUpOz/vxG27iUzU+ZKFOly7y6U7EJThx3eqA9twOJFD
FVquQBszintwMLtsTXK+26r9hN0WJ5Rvr2NtiI27q/iaZUY7Ga6kH6xngBIzMmCr
yQE6YSnYKNM7PKG2tHDgmgsGD9LuiCeBJNKW6LM29nIWVsLni3JJ6EDVLOxv8fmd
CoDc7f75sbdoyU1IaQZn711habs/00U7IRzA3zulmChkIUqyMBe7hr2hkWkMw+Jk
YLO5bXeRWESFMS6I/tIqkddL4NMC12J9/O+WfHN96X2aInC2kuYxz/frR/RO63Yp
jaeQhYgAyUjY4Nk4O+ss2DsiIeotIWbWhFRAY6sZMto18eAVw7oFGavmY8unWX13
ua4CwUg3IfLuFkc8cwjSO+XTF0CfSj6SUH2+MSr/VUYLKJ6/JzReyMUS7iQzkj/T
9EZ+72Z9DPaFP0i2aC1ob2ydSUajQcWc/KMYoLEmxDtGjqOxW93M96CwRDbnWgGn
rGpQ8wXpnacCheLIi9b3J9RQkIhHFVrdL6QHCHop4i91qqv7MOHGNrn9+P+p8Fqf
6Jw93Dnzbdc1GSktf8jd+1CGZZvrEnq575/UzETWPI9hmOVUEb3eBFGCb+AcCwou
cwcDHoz/1qh6XGl+i75plfTgEUrE+uiCIIPMJzSox0Y+Bb7J6Z1O7W95pre+zpks
E//wu7A+PVoFIs8cK155wRRBmCYX4FTYF2BwSxE01vg40/cBarVVU871Yz56LQA7
ReIxZ4S/7kE4S68jaWoxC/b3hRvLR4OoW5GMVd7GcS10lOYphNsPu3H9Pp/y3/sv
hCs0ka88QEhmXtv/D98nzAzJZszVExQXMFv6huQ21m4CvV2ffIoFLzhreskonfvD
b1QG6kAG2QQ2Shx3tB90ozx4CqidPQvEM3paN1RXLURaohnpqIwMuJh4hPVX4XZC
lb4qvZnkZ9Qjk42RsqhEZBQB6Y5hOZZxIKUzoqes/L79lB1TgOl3fOCaSgzLhkLc
HWHvb6DtfhFkhWNm05c09BwIANOGS4LYvqfUE+qtCeoIUXLis9DwU0GxoikIefyY
5l3X2DicS+b7IygHv4OxftMxmbNGxUn7PgwrCrO+7tY6DuxW3mCFJXY9nHCvxRDB
V4K/jSnbtfoO4qWtfXnv/C8wfJxNI5RR4KS0xGCc5ZGZ0dbCPzTf4szkJZ7j/JM4
HrXpoWm5FOzHgk9oUz6U/YSdke2GNB4e0rvTOwcG+CxziomOE3sKZL3FpMsOtM7w
U0RvHiSvxn9CEG7GErlJyNMMRMFqb7rGR4GQHG3gPG5eByd5HIFT+sMwXjpuE8+b
FNnw6POqYErpFquZJ9RnbNZ/MuVMod8UUI3kXhWNT9zpNFgsabIdZONMO9EBDuBd
eqLiYz0dcG+N8uriZcWmSA==
`protect END_PROTECTED
