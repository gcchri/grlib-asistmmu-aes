`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97pLqd1owH3FMJMOIDnq2GSlnsr/rckpyW9HvMv93bC5WpYCkMrs0k79pMFwKtzl
A2r5zajxOdzOL8XUGG8kTxM01EX0m+eoAeX1e9FKm9pXKpkFkBZtPJNy1EWP4spB
QvzWR3SwSybKTRs9pAwvZTAlPWOaXWEXiUVrQKhd4hk5nIpQ7oH4zdOnnMqV1Wtb
TZiawf1rQq24TNL0VMjpJY9xIIFOAECs1ueaQbnafWRtbVopiTXq4VVjggA8UByq
DMzhoKsYeukYvrE+cI/zXSD2Gg2aWY0xAQM4NUCUwbaGVCoaCbOARAys8ZdWGwbO
GHfMjANBnEM0KrqPfUdRZAQqMEczmmGwqzMNS1W9t+xmGTHqlalfu68F4suYFl7k
fJr/5n7jQtSnhhr7MIwP53G8S0ew2mA4e61zD/1Ziqd588HF5rxDYReEeWWdM4vk
to6ranwn9BxAUWYegRfGP9ybqODzbEiaGBaEqIEin7jKI0mJW0W4c0RByOTg7MSb
aSaAi7u+4wD0peB3un1CsN+I/10oLhzkplK/vPFz2URvQOQSfqc+C4ogrJb/NrAD
TQGhjfWtjfLGygO8znOpBpdqSsc06BZyKXATTy/G3NNXW9AIp3geJgiafkZyEHAg
L3NRytUr1pko8nKeXazQsGLIuBdqi0kkON2ilqoOe0/2qV/1BTmGl3H844nPY+eB
nYO3x1i3q1IuWj2e1d6d7XWvDpulWRghxfZiADmoUalCotExA7ei59kNwReqxZi7
4EXDm31dJ81zQ//keeeg2wSl6Oo1jGDrO+qfYP5odSLObKRiHgwOB4jlP20pwTSL
LcdYf/A064C5CcUvRCgNBEmNVogZXAPO6FeTqGdVmCAyhNrfGr3u/Rnh2O6Q5Xnn
QioQSSj+N3gkEIJEPQVmOtyLG0/RI5sBQqXSW3g1me24W8Vp83qKEkg5cc6zgCrB
9IpPVrgajmp4FBCQ7jAuAknDYPcluHdPP6GnK6nsyECiL5XV36HNcbYQfhHK4OQM
ZoKmNSlRRpN4ZcTFTr87kN6QhGGo28oytiPIIEP29XdQmYjZM48fQWOZtPHYo2I/
V+O4E3kUbTKOzGOpfUMpo7MqkPLH75ZXyGU6SeZUZhPX6SrOs3gyBI2H/BIlh3Ol
vTP2I3TL9C6gzHmjtYYYdjiPX76y3yrC+bsbvhlaw3o5YVXSTthSjgQUmMsXA2ba
NJDTsFhqzieFvSUIM9JukLO2andi1fsLgR8jpGdbofzYRjpl+KEN46xWqq4wTU2u
cf92ovMI30QpohPW/DtXXMIHb8wmsK8Xv0XRV/NA4Hmdpveprf+znAbA9fCpxLxV
d/y8bpdOBmsTRSzeyPFWqNHz2rX1q1HDkQQlEo+W45Ky5Zfm2dBjvNjYeZVfxgv8
zRTj+tNQEEnquSwnEhwbJBoFLDB1aBuJytOTY6SkkjuzfOGgPQhMbxsG3uyukr/k
TgTTL6O3g3+XaBpnZHOw13Ty+hVYKOldRt7xgZ14TP0=
`protect END_PROTECTED
