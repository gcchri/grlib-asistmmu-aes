`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHCcp+s0M/445C4mnZPBL2YFonk120Eu+9RlvmZInzqeAW0EtKCTf3iwHoursAI6
UFGZNrxArrKYGPxj5hYIqhu1mn97tQAa2HvSqRpTe987y5AX55bdnAPRtt6GNLPl
wbjHTD+pYuhPMbQ2kwO+ST+I4zvKjpLiNiuI/aSuBjfg9TKDrX2fVSqH3MD1YZBm
Ky7T+sFjxyh0K/xltolU+L1hgAsAYPZZDjzkH01GUPcG6HaiTl6SJAvzegSU1ocb
5l8BPoaySai02yClVpp5rIzbgE0Cc7mPeBdVlPh0aj9K1fGj90Rx8T61zxfakWnu
P+BLKU4q2KNbCtXIyib0TSVxK3q73VoSDIsIcrehOL2PDXGmbUDAwRjQbweqi9Xb
z4qrKLtthMAQL7ZR8fnyIuwTiucyVBMBDS5/41l+0kqBPHyEBi7sVD6X4XWLyHn5
jb9ll23BFQMlesT98RVazhs2/gQqNrhb/Tt5LljFjBRwi0zoZ5HjGONSgTwQuam8
B1P/yYtEpHxJpdrESgcCunR/Vsq5IxQ18vO3egq0102nqCFLMhqRUoexjD8OWKgy
zoaNEGP99FlQCG2C1EvKeEKEVNR9k1Mpl55ygVjQnQnad6p8SYXy7wG2JcRc1JoZ
XxN/jc9hscbEi01SJhlzyQ==
`protect END_PROTECTED
