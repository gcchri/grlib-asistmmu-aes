`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqtRwc86rPojCB+/pSRmlZOb2dM2r7J646W2I2flGgxRxW9NLLgE0GN498ZuHg7q
HZq8XFylLImnevL8noAaTtFnjTvv3Zifn8KlyxldPb6lhz4TFXuZ/t1yfylz+8dB
fbpke1rsk/r92vq0GrB+/PJbqVS4t7yIGA4Vs0XtJBasUhPpQSXxePqzr2FwQVNR
TBjs+BQnQhL2wIHH57vScWN4tzUzAcoq5LRCvV+vH4hf2zsZ4587yG8sBXGnoh2N
n8/X1NwAkKESrcYgluEVi8WI8E9ctfjJW2YD/Qm7r+KqqSXGTfTLoC4MSJ21O2Ci
Q1Zi2acqTd3/28mlHE/qo5vIAwRX3VUSj4AwAsATupOl0y2VFg0h3REzbOCEZkgg
PR9xro2/imumEgSfCVnpFysR/QGVgMNFTa7eKTbaukQ1yi4cWe0+WHjISdYZOyLB
S+V0LFyP7midXuvKCW+VwW7xmLvJD5L2veZ2an7chpwn3aTb/QBA1cLc+1tOtFXj
wxHSvcLsAdb0LETlUjAazxpErGXbPfa4kcBKvzrzgs2L6TAG8Wf1lbhbldSxZ7YR
u4lhDC4gtlkk8epoQfvWP1r2I0PNgZR341llUtJ+27irTNlQl4zhZd4zoIYftO6Y
OvN+DgeT53C+z4qrlU0WEaMphQLjyGxjGq5flEHPejbzfrgaHKCWLaQmUltG4wVk
tKjJ6IHr/mTiQbmNgE5paNhefRqpooJXIT6Ho2GeOV5/vExFCfCHo4FKHwyU5lPo
f7cFSc2jMEQKLI1NgT6sFObSgAV7NFRo/qHGDAszn3Sxe1945UHFLzNLdw2JYjb2
dSJ5zNHp3uAMDX01jrmDyfPeXN6cmqnXFhq0Mkz0X9f8cZ+yR27kU+lPIBHgPfs9
mYCYcfrohOMykQdVfrtgtk9l6+boRLdeeHTZbiywbQGR+8urqDbn+Y8hPxjVsJHm
D7cMVR0fz5wRbQZVoK0t/fS6lDeZWKdWkzyaq3hDAygcNpCZeeOIjelL+Ez5g5nX
xhclVK+p9yBIOEqfuchNOGV+KeY8sHPVoA8W4lU6uS1RmvxTeMzawd8+jIeMjO3x
jV8RcTlpFo907+pRGKBTVR77ReM0ZxUVi4TTzAtBZQLQ5I1rPjh275o+RCqvTMN9
/YUA64yPxdKXF8uy8ktmPnSCEgB0XZsTsrxEoIv/P8XynwGGPsxMGA2O0STg/JkW
BsNkOLPlo5FOsv6SaN9bq+C5PUys5B+mhKltfi1ZN9h2feHcJ6BRY1ViBf+k7oaj
s0+7DTuyGkf7+JVzsqSNVPBmY8GNY+ZfY4Vu7UbYmlEpp69cgVaDSx4bj74yaVxt
EE/h6rMBPEiJTQsO/PD8D4Jt0oCu1yf6KbwwwTc71FFtuDCxdynLiNPDvhPMEPN1
8jusVHbLMRLYJQXG4+scN4tJii9DjebosXLi3V9MG3586FKvylzbiMVSNRGKB7zF
O+K+8jPkiteLn9x6BWgNFETnwp4nQPTmzt3IUarTTN07YzJ0FteemzW/Udp9vPaj
ZmTlgY2duNCjWj1f021hjTBy6lc0rHnScVVkgzHSbfXgYkz5P3waBNiW1yyWMoVn
acW6EWDa4fmF6tw7dKE08DCxuuhZ54SAx7XpbRQq8eRxtNTmmggvEznp7kToXykm
EAO/tVAMyfY/GI/r5JrzoeBfTos/p3T1iOMiSfciafsEbVusVltebV4yQfTV0eGK
Ygvr9JbcTFYPDYV8SK4fLHairpsk2UVhclrP/S/uY+syKDWzE0PYTO7cA84/gFqP
BU/H2JQi/kgnS447Z7M8qViaXrvq02adjR2RQCJgumwvKxbWgitFW2UvSE1RCwhE
DdulwgC4Das6vH1b5B2se4ngAfQXlnPA4vD5CkALOlz6/bVmHe+j480ImuHALte7
R+EvPm+iWfZTgWqMV0xqlYMcYtiSRX1K+GRMoQIL04tPIgw7ElmFqz27hmh9HajJ
May0afDTSXYD9yJe3Rja+vuK0ZBag7wQm/ABrCQdYcdxTS19v7Eg8xwm1SwwkEzc
csBXF179icB4AOiIqMEWHIBptNvOLZbBKgR/CEkCh/84qupcKfdKrCE1RyPNfCY5
E/pazd7gjaL0bo6kW4V5vKzHasHyq+oIF2G/BHlIL4QeCC2b2zoBpEVY69F/N/tw
ixxT3dRS3CNqkKogjrDpSaab5aBf1Dq36rTDMRPTAW1WD0VL3590F7umI9T2rN62
+1/CBSdF03pAxedJdXNTCpCsmYSpmIlS6erQHQEyehWKipvsFdQUELpPd8uJzdZh
ZVVkZ464YC0Q9zgjZj2MyO9fNlAjX3GBbFzWl+/ik8UGDsvJKrK0HK1WrEgGXq31
SPBnAX2Epdvsjoe1K8r07WcKqEK/VHRS8Le9yVv/rxhh5mi5gk5CiNs8lK+ZajxG
6sxYTA6dCMkvM39FyyPDvj6Tct0FelEzh6KR5RL6g9OFKZ8a0FQ7ABVespM8pigg
AkNRdiYt+WYdsn1XE5oIgKJBWnDjX9GWgo025pPBuIBDJS9dsXB0rdFnitDgBMMb
z5nL4fRyaxexW+fr3HOFpdGyihq9RpCxtkxut9t8od6iy3juQ1Lb+RGPEUcvh6Tf
c97wRHmmf4hxU80EEYJpBG8ndeH2F+wz13NkEGlakdGL46UzGkf5UMERG+doz4Fb
s2dt8Q4UFntizBvzZ/fqhw==
`protect END_PROTECTED
