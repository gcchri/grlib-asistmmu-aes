`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8glCc3Re0vV+IGDz6Gs7z3WZUfTdN5g6+kPNPYwKR0hKSQQ2/qzhyFXLfcnGnQ6I
0tRlNPNoztqhLZjWApNmLzo8BYJUAPDVlfMbPZGb/ObZrR9D2lXwaLALp3RMok1S
eiYdFvbFdBCzfUu/b076k67tqVSbV1mSDLdu2PQyUbJuRrSoMo/ZZGZVDqCCyNKs
2NncJs5r7dCJFWaVdKladq3Z9ITtbGdthxmbzPHo4YRdQhEX0/NgWb1wz3XaJlYA
HVmwZviwhBxaSJKlaRreAu6FiTjR0aD15MSdwyW6PbRQtj89owGHw8AcNjW0O9dc
3mEyhyk7j89rWA/tqPtQrZL8zeWPrl7WXr0kuudTaBwJ9QAICcOjiJ9iAhdfR5hM
MWCWNDsPoGZ19Q+OcBSgy3rGtPQir8Zo9HSGQoxTl6bAeFr4JNV3/uW9smtMoF2m
b70K9ztHzcW2ch5wQa2Dy8rLZ4ITRCc+YMLdkdX0Igs0emQyhgOs9H0bWZ3URPfp
agejtL2jmB3ozHs6q6fTZ74a3p9CenkA4sm3MG17TfIaIszldXdFwftTYrm4vtAk
2MOM8BBnnpTQ03Of8G0imnMJFQ7gRz0Ey0dXvP6cSFQ=
`protect END_PROTECTED
