`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76IGVmbR8dcrt8kXnNWGMexAzTcZ8e7HjOBVtSntzMCkp3JTSw+Fb2+GDmm7XkZk
53FCKd9SkM+jecNkFf3dE7+dS/tK5B+DhrT7G2INpiudtg4l4olc6piY/sGuCKxZ
7o6O9F8Ws8HAIsrhXsA1eo+PP4GAoyQIK2bWWcv/NRnyrFU8Kdv6pqocORWnj8fb
2ZIKn1Q14y7+DuBMMn87xgVpfLJ9c0GZkvqoMIreehuPlw/taQu/v1BZ/OirC4Xm
qW0mNwHEOi3mSiTHYiY96vXZN5IBjEDLh76CpOgTL4fjCVIhLU+E5l3UCDLoO4f5
cAG+gZmLb49Jpnv5vAQmotB1GvfLYD0KyyuiDhJoH35PnPyEdhkt1UhOP1Uc0SCs
S5XcF4MUqySO1ILYlIMph5XPDRBbmnWvEtGgKiOuMoFDg3KgIOx9YPAbgDLkR1ur
WXSSwTwyuX9sQTtv5ytwVbg/VmWGGfYx+7IKGMVCBGy65F0rpOQO+DrffsvrvJpP
`protect END_PROTECTED
