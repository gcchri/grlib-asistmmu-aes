`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBQiZwG/cAOu55bpejz5ECNPGBjJK9NcCWGcszfCZzqSUCbuSeYB71jY7OfL3Bx5
icNiDNuRU93rcLLoLBfUg83g5enm+Da/fFMPDCDRMmsvKdW5eXD6rNxlT/+/oUHC
fb4JqWZNHKjoI6XDV8tdv/X4EGyGzUpLr3oLD8rgbzP78sAElzRNmsgk6zZkIVmQ
L5EwFK/TtyGLQWs+CoXRP8I8AtjIda9gMeqN+ZHTLdE4HI71JtyRpc1m48VYuBWJ
J2/YUvXtPjqjMTSUtRjE7naDhqCTU4GWZz2UKy1KWJhInKocLmGh5dKeQoIlW1Y4
arKOw5k6u1vJ+lT8pEIzchz+c5OqUQS+9Zyi7HwNlLn57vni4Qq35ZzaKpqO3I7o
WlhlNPIT2XBpZqYubkixJDM4MP1XEvu4WyisYpAT5qaV4s7ffqVIep2QxuZFMW5g
cF5kSpRW8zcGEjUHxfG4Qsp1h4EzMScEwUXtbPN+6oHElCiXAjcWQNKmSHVNdEg0
CV/D6GFaY39Ep0q3Hx7OEzzxKQ6mbgtV9NsPFWmZG4C8QxyloGCBXomA7sj+ZTnb
oHBdgEiMX4wEvbs8CLW3MO5b6nLSpnDtt7pr2UEShDLO4gvjDBHHzbACXoZ+kCVs
AWHo50QPkrBIuk7E8ZJdV2GP+wTHu6Lfs0+mH0vpyFk=
`protect END_PROTECTED
