`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mt2RCbM+5FhmZTtOqa1W/8WozPIYDNcLAMORkyKahXZIUTJkWWT0/pP2FvjwBlLE
lqpZTzwTe7xx2xTGJSjVZzsEpYLARAcOakxYW0RSkPAUWczOG9zEyX/EbgsUYbuA
RqKN9jlY0Dc38Fm5nRbXtqjAPow/xZX52gx2tRj+D/DyxBnu3rHtg7uH2swZnhWH
rLarUoBFhvAGZaaiMz8DIR/1FwwDF8jxGgpOc1zAofyOIfjieV+QaFiCGjpirgxY
AA/FIqLhYqgD0Hib9yKXNt55gYSH+C25wQxdJp/xLicq962VkXafZa76le2br5vM
h0rv3Z0f0aOohnIkMDgK3g==
`protect END_PROTECTED
