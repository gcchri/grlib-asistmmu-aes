`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Ha2wT5lLLfWV1TMEDZ5NmEzpa0Km3fCvSMdZV9TZO+ark3CvlhwJQVZxaFhQa51
6TSeXximUDcrjuXVT68wX0NyA2mlU3B1SI+Zp4t0exBtKZ+kXHUBrXOXdM6hsBrS
dxJGhXCFg2AMBV0WYJM0Tv1/psoQV9IfZ17iwcKZ8niakFCYtNt/B8cfZXrDXs3a
m5Jddg0s4xSVX2hVgeE4IcdbtUOHufvEwt5iuHqBINREQcW2+Co76XnZ/cb/JWAC
K1i50j8Lq2o7yyl9Zyxa79/lKd3B1e3XFqOH0f9M7H8Rls/qxn/NDwQZw+nQ2rVb
bbh231AmY9iFzISNR15rx2QEBDcfsYO/WwH78PESt8+8AkIud6wikcbGOBjj2xfF
H2juy5/uPfuVPQozUljrs7lYvH5nVBKaDl5pYNDC1kGDuwqOewLQeN+ja4MZwMLi
`protect END_PROTECTED
