`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mymXKPt65vFyF39eaHT7jIb8Q5ObRnBSxhSxrmEsSaGqujWpCjQYGLvD9sVBtPnw
aCZsGVQPR6E9T1TLEZRERO7uQJPsxtLII0zt5LfSkR/rpli1jvCcPQ4UHbc2zkm7
ISC8bBfKWQK9LQq4kTGBOQmUQGg/y8Ad2jGMt+YMXI7L91yypY0BFEyTgNPRJ7f+
e+0EltQguvaYXshP1EHdLg==
`protect END_PROTECTED
