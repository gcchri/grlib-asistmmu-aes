`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwhq/hDTrY3xUQKCmLcYn9xrWHHazgQHDKh3JyPbM22mWy+QYMR+1klgDi3gZIrV
d2b/fNQTsxOPLn3h+F65zBJ+7jrPDtU+0CszSn5eNCRwo30sT3yYhyW8hSdd9HAH
Bpb24UqMIBhnyAdlB3+BfC1W12i1XyZg6B8+RVr5PbqCTDcrpemObu6QyZZph0mT
Ei3wjEwXiZl9lxl0NAB+fmu8OyAwDncyirGtgS2IK4TIVoo60T4XoAaDVhzfSCt0
ZYwIQT6kpoasyTRVK82GlBXWCKU3+xRnAYxl1MR0AAr1uzPE0V4KK113LbBqpuXn
TpkVuaZe/FGlmBVI0lUUbLPjI1IIgpmVB3pv7DmFcNFDcxp2mXjcEM1m+dm+m7ko
SbchvBqh2jpL6RXcpU6HQSfOVIthn2bnafyTY8rnDAuMsHO4V+olvfoXHBqs0mI0
hLUm6dw9dtrojrxAGei6WzHA2qKiqieUsR57V4jhSY1S6CXqkPBKneR8UCul5owm
VW+m+PC4Ipi9uHb8KhIQUbN1JhFVJ0ZdlN5xbrZCizjl8J7BYZ/4NTAJGAwZY1MU
atZXEWpLuaUeI/QwZeHcb2g+xKKCw9d0wdlq+id0p5JM0IPVGuc+vW/qvQM+m/f9
c2DHuBoMLKdL1Iz/lbOdZA==
`protect END_PROTECTED
