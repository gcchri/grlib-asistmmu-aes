`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8IHR6igOqRgD6CIXJUuuxcZMxCmMWGnk01ZcXBKAFOGaQY87LNBRPDv/SyYrtle+
Qf/D5NEbL+9Kw+VzZIDChPpTgNnLrtT390l+hOMl2R9vZiq760dZVjtx576TgZ60
0s94VaEjJ4RcneqQ/r+jP4z2xQO62Zbu3kbrP5cJy+Ia7RQgTbs91SRKWqo7KnKf
fZaTxeSL4AE24TLoVt+ljDFWGfY2Ezbq6xgoVRTFt/S77/31xgnlLBjoijoTml0+
4vF5SE5gPWDY54NiVNF+JdKQbRBGfgZuQHC8MrCo71k=
`protect END_PROTECTED
