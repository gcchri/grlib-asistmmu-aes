`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Wy6Ln/ZwoejLh/Wi8aXrv8+7Mn/QaN7UA67D00/5NytLXRHHQ04GfV6YijiD38t
G7DxFiLg6IPta9vMEiwWXhPzMVCKuyaGxkHEtZkdXBIHASZSCewAeuAa91obRjtp
Db+fIdreSMZAZS/cimVgk8/U6MtKx5UNTa/fVR2twVnlHrIEGObPzWe4Ganx3O4O
4ohFOQ0Nqw05q+aL+bvsmau0BOk+Bg/ItqFTavPnN1Ny6/hTcmmS8KyyR0F43z7O
GxUlsbpFohVXiLFfMtFlWraZ6M7uc8lZkAlZl/dsD7QvTB0cP2OV4xz2/jB/2+XB
CrL6tj8c5OW0ePZpcLnqDrJEWy4dB6wkxVB9fcb7Yl1n1A2e7qESMgh50ArWrIQd
`protect END_PROTECTED
