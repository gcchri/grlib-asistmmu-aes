`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UM2MTOUkWOvyKSMubNfUwUk6r0DyVSWHR1O3qVvWc10YYyN6k/nsqQqtPwGMvcUL
n2WZSgeCOCyJkceNrJiLx8Y+g8JNxAU6bTvQTGAtreOzQq5q/BsGdSVEAhatWXq7
ho18FyX/g6uffzzscqlUN7tHWZlBZaX1pBmWCTsE+ZFqwJL7115tPBAatAW/lYtH
3Ht6JN8bSz20lll0eVmbIgHTB5uQt7CVFIB9iTJU3PJNGz6tRYipSvLrX1dKLIFF
/YOgIaan75QoYH/NYfIb7pZrfPwbO9pTM3l+/Z7re1rHBSkI42d4/b3jK8A/Rhfi
D/Irph7zEMe8N8D9AS9SDP+//6fS0MuXM4edjD5EIwbq9GwNIE+Gzm9LkRIOie0V
y8lteuG+ZH/QUkX3iRDv+B2pNSvilU8xBZUdldzwzbH53LOz87gdUgY8dgvN4NEu
GysJiQyAaXCbmqaRgzPMgKQsaMm+V8mvzV1la8IJ7SC/P1Q6ieIDXSAW4/pS8XKG
FiNdMOpotoEbSjt6Q4hFyDv/zC1ttre+wi6Sg/JPQLzVdGnV2dQkkPOrIcO6cmMg
Bz9DSS5kE9dnezVYx7D8jnRnaUQ/RzcLgWBGTcgadAES+wFC084wSK6Rc8XhTJw0
1q95he2+uFZVk/CuM2xfSI6eF8vk6QF49VinXP7UUgmSetQ1riUsIs/Um1PD6TGD
DXGSfAZ3IeD7m/Pmeg58oTQ04SjdRN08rSZyaXquEMKY5yojg3g16a4Ad4RWsZ/V
yAB+ZnD6k3b4LfKf6hB6+xbpYuaYbf8zd7TG05VD1swMl/Ob2ljHNf2F3GcdlBYS
8I/4v+k77kLq6HcA4u7BGZ4Vud0ptMK0j6hyV6ULkEOyCxLN9Ads3/xUKNnNGWyq
OubKbKGgifi4uUIHyMwbnbs00Uxlq86nHe8dHywTrlrT1dtB9HFrkCEwfvlJvw/x
`protect END_PROTECTED
