`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YLFLTkX2fuODwPoQ3+C3qp8YUoaX2QYTF76IV6eTawfQSSzTASpyOgzbg4AJT4ge
eJvQOHOrfCcm+pD5KHZAZ8cLhMamlQDWkssZa9fPX4dtICGSZME6Cc0M4sRbbpXx
QWn0Z0kbJGEaHdVYEAfz0scvNTR0ZdRE3sBfCIEZJZg0nzdSooyJn7Ox0ZMGJSsK
gzFXule6VoXEg6wWAebxWGhkv5+TJUzNK/zVmKF2H/YlwJTAIfGXmIepPbJ5Me3w
F+AsreDIb6uCpp7IGWTBFsdk3gNnDgnP16cb8wvW9LF1/tlH8y23BqFXYlvDoJSI
xw1MNnfHaswVQ6ovgJqmnFsHes8NChLVS0aHtw4cKySbVJEdXiDzjP1Usk2fCbbs
1ZyVvHp8D4nfCu/uaKOAQXSeSbLQjTuaK6+MioSbowVFUBzYzxK3e4SjmS3JH210
xbGjC31yNYmdFucvtsA4jm5j16P7ucA5PhHGh7/+oqR/Dd9Q3ckL8yAQvy22JGNB
7lPGmPdwseuw6qNUefrPyqklPyMW/icWKsIheRvqmNGs1odp/bSJioV8D9S0rBa2
5KaJ1yHGYWlE4kaIroIOZJ9zwNY3qtF2BZoAbmVil0QiSgGTmKHveEF/hQZ4RFSd
9NqBTTFwMNi9k/zy0CsnnkAjeE0gbnc+2Kn8L62cjMOyE7W0pq4JlCa5NBO5l2fz
CVaGm1baXDq1WW6yW3Zz5plByo9owNhtDNlqftDTgLF9Vhuf6sXbvJbTZTX6ylqR
ilthS1DuIEJb4zeaha3JlWPuEu2DC/v/1Hm2U+EqA2acu6sOIUGxm5q7bj0RzIFf
w97flAnL/HtKsun5GGS4Txq/ttUVzlY51o9wtuf98er2XAa4/t/2zPQX5Q2ZtX82
R7ZFSclKHJXUWBktckeiYI6bKMAsuC+lJnwq+/u1liJNwg0XjFbO8+6aAHSfubyQ
olaEusvC0PWFDRal0HvFnIIQIpRTKWZ41r7yTlsUmhD46rynG/+QcL0AB2rN6V0R
JzVJaWwvXnfKjEUBUSDKnW5OJ1lwtX0EGAf1oKg+sGkBf5uKZV4ev+JU6SXYaA+s
v7MnFQPPGIirmFYzG2mZY3ZFO1D0i0JYCsALJ1vka5oURrQBfod+bl2W63bLdz0v
93Fm8GDQshdOuZMeMys4LYXofFYaSgtEMAAYe/SGJ2aT1ASSpmYiE0IOvghvpjtJ
RutYukqfIZpq6RokRPHWogcrldoOLPCaTywpCPoKalngUxqoHUjILtlu+bJzBRQA
4MWEVlCpnlyYyAVbfiDZWffuAj8RN5+L6yuhAmnHdzcq0CeRmiUJL45PrZGiOK0K
wjW5I3MjYhVlCCzQ1CkVCkkhEx97ATn2BLacRnR1Ll1vWwEMMIiQ8+OJhTKVIo5O
nJqs8RcKGRdfL+t2kg9PNmSx7LVFY/WyDovVFwRd4jPrIUu3Av1HmzVy8LSG8qR/
m12DR28WICOexv5+h3zB82ckMvNzZgltrgcN/n4mt8cL8Vw3awM1SXBhlrp0gS74
6HPmT/kIsojp17GggkBTXC/uXfUWyK3JJUUR+fY7T1E0mQvJkbkEl0sTiaujtOA3
B84DM7BGyDY6IlgNb0FpzFHmcr9M0ZnrdIJApqBY26BByYb/uFaDBuwhy4SG05eY
cPr8EKzvRGa+JuBlx5yz0T+fel+uKrIeEUhlUyzH5CrkcT0XXBoIKjjoK8R/Wr5A
n/7Yb2u4tifE+qhJnMjxoS9t4Ydjd4/9j6kgvkDeYDyk3dELOtneO/CSq5h3mDNt
kV5o/Gc1h0YI1rH3+NlagBIsxy40UqubbJebup5HEjFjKMuzWqk63cH4aMr+zBhA
MHeYvDLGntHntSv3GufJqkIPBOmU4mZPAmGz2aKnZfiDgOLcv5958KSQqETIKk2Y
gOoIrgaDW7oHBsgTRxSVFhOxFMXvQ7uvEfERrZBdEWo9kSxkHJrpLg5/HABjjvmp
JBWyilnxRmJ42VRHCfjg40+pLD7b+12TkBPynLcuRzXqaoBvre4y7XEU5VxVTaJI
gxIYcGDSGErLxilSPM3S5D4PSZFpw45MxjvF+rn4jV817OMClvhColQCJMUjhrpG
nd1NPvIbTj9OzcvbTuLfQTemUl6Wea6sXYDlHz5KplKDNAn+hwDbdVUODrZ07ZuC
6+dYe/Cv87kReU5jkJnr+ikV5jXAtvSDs13gmGxSjEV1RmnpA2XYuXnwvKnivp3P
9ih25/VQrmUQtTkT7Q4Mof1T4cMI/dnhiMAY9jAI9SunQfd8mO71xFPy6/s7KOJA
wwz6Vb6pdtVAt50Ozx6oixjXjfqwjdCUqWs5V2cOdicgD1RTWuHmjhKoNHs3dXAi
QteoW1yZTpvfEInzlXtRozblgZsws3eqqdp0EMin6TLlET/ItvWTpAh5MqdgSZV5
p7ZwddkwrhNo0sWMnHbVQMPfgNleP3ssSktSvE33p8gg6XGhnphaRMgYzLI0fc8o
puQhKhukpCKL9tLyTvh2PY59go2T7lEapItXqCKpoN4KXfR9i0IhqHQ3P0zDuyPI
hvd/gU38rYtXfcAO3TWeCghJ/nXMAXkK3nQ+GNyzyMs1Be98dbIsBx23fONKbWaM
Yd8YNzrFX9IOU6Uw8/ULHTDtuALgnK8zA31KGkYau+/K6fXBJradizH4q/LlDkCZ
kEMoE1X63sU8SuzQ/7hRGVmJkEty5gVQWR1nN8Zid/9iIQZowKsYXAevK1lPACDP
lYMqvKlHYohkS3Gz08Z1qAqzESuHIzAw+tRVYSHv2RioXudA/Qis36TL0ZV4o5XM
uPcxBXJfFHoa17qnvTgA7eGN3Xam8lfCB+JTkPEEIH/ychlowmdqXV+AZXpY/Iho
5FA1Z0zQxDnu9BvNTrA+a3s0rvn+ZgDM1aeMBsMGDU4LbGNO4zzDFtW2217aiEj9
/8xFY6IgdUOGt77YIBtXmqvFaSm8Hs9FPW4sV7W8EK89gfgV/kVGWdGG2xtavVk+
9f+e4x55Mhs9Xpm6PFVO8/1aC3L6L55GamlzRO2WW4OC0y4K2INXHK1NosgEum8J
acT/tK23HXvomRp9c96u4YKlyeiX84WBHyFrRtwUBey7W2M8U5ICN2IcmrEdJKGb
COE+fxZPO7Miug0Lp3bQDh/BvplAraXqulWUvTSFjE13bxM+NOSF2l7FZMSoT9YZ
S36sp0udPFv4CXEDwBkaKykOfuSXshaNzFypRSPC9vZwevAFu8UWimUrGi0TZe1b
KUSv9ivZp5Ry3NUBczGROPOM8VRECTTGqIGAzyIm01IsOHzDHn1OIG47roGqmFyO
Dsg+uJWoCSWR8QSNrtRjXPrmxCQBLbSyAW/w3Mn0kVph31azUEJYVhYh8uITOhD0
GBF4ypJNJ/cOqwlrL8zICzdjwLGKRsBZUL6Jdve5DT47DzJK7BZ1B/3KRcn5QxLz
iQCNCEVlkGBkeKeK1qK5f8whQ9YASr2OBP7fRrsRrRlDRoXQdPGZaDwATF8x5Y5K
gTWXSkX+B2e7pvTiZpamLucqekUtVNJEYrRuNs2SZBgKjIqZlfu+OiOjagAPhuhw
LhduaDYqWGs3LgMW3TH32ayenpbn3x6+OYlwZG4GsWg3MD0JIFYFR5gN/aNPJ50E
dBShAsz1tiYL3qHDEglSxjSSmePGysH5pQhImkINgz5Jvgrw3AOk/xXGcbTTOgZD
OWbrQaTGY1zxCzE/H+kW4XAJdtt4o4QULDaLr7tITLkFImzg7tS/yju6UKQoz9Ez
RdJvJXoMf5cC+QS0zI2LJqfu2B06S2rC+ZV+SKBUcXWPcE2edteK3+3HX2HsEp8v
mO4J41Hk/+czg20IdJAUW7XLwDiBTGf0Nxh+kNIlAHOIXvLlpv4vqZ4xgYR8A50D
Tsb0LrTVgp3F4dhkVj88hgCQThqGP5xQo4II9FCIeYF8nIrMXLByij1WKMMvsvrP
aZ7ZLAH5jCMbvmHJUoh55TdNWQcW5FvVEhvRJODtn71Sx8sZjJMeSwKDdU0s1Bvx
O9t+GEi4RnUAT7/XlprgS4qh7x6wZO/7/P3fqVACBPTsnqR8TlWXC2nf2HONW0Qa
xCyT8XieOlanZyC6uVadiR7DqSUVGUkXuFUYq8cyAwr9iVdy73bxXuKyqVIP9TpA
9R7WuTw3cF2+U28076SvlVWMABYeTwVO6yzptElrMIkWmrggotKnZmceX5ho6Qkx
JU79qvRGKaOnOWnrVa9ub1zWO+lpC/R6Pb/Dk52kmV8R+7BIAj2l6hz/RMpLjli/
a8l6AjlYTFP6LTDhZ69gwMgHtAk8K8OdbSY39Dg4Oc2RFSuhpaR6YYgUO8OO0eXp
jEq7N+onavi3D2CM4auHF1wLjJczN1/iUvIjkxtzlqGgFwx1yegxumrENnJNPYhF
Rf5cl6trEC9yTRbSWGbJpsh/mFSC2bLaoVIj1U1e6mU9VaEHXKCclbKn4AJuE65p
YPTCr15pMyKy/oTarPeFXYQRFQ0VIJvmMq1S0I90lwatq7QUWRgQpNDu8BI4NN0t
wh3qjsjTo+UIFjuc35SChE6SmiovfDtMlPg8A/ji5FLLr/e7warcgvl4yST6okiu
IpOLygOLxIqA3WZdvEY+FLMBR2a+Rja19w7pZhtMU1xKRWrQJ4/sjq7AWn+hhLHo
emHinpPr5gnHPg+PBCXiAk0uxN2gDVIdtLjZlp3s2QWvElfg9rzgtdJIkcBID+fC
qyBCQmq14vB32hUX2fzLziUb5kc9/3wYuXvTaDMKYx2aiivQeLEj9WqEtiDKvTa9
2+9IOva+AAhJHFVBx3vJPFdbQk6KYUB5Ofdmtr7tP5Zr0HQCw8uWrzBuYN+Wq8Fr
PqxoR2vx+Lt/I5b3ApnX54FxSu/hQnqf/S3XQdRNW5O5ijIrh8yea/lUKHWCVe/2
pB5LvcBJ/kEuagBv94i3lXXj1E27x9gA7uWBff1t31TkRbm70QmURz6Ont09bGKW
BiuaszFszJ8PWKwFmrhrvr8ymZu8HahC8wJGJXiu6xr76OJ7kRErx5YjxswowbHQ
h5NJOr18HYHbeskTyUbz0Xr0hVdBAl9OnsNsCfBHGG41t5HwjcQCvc/Gn7ahgvtx
9G7mUIKceIbK8KFxpn2lORNwkI7dF/dVV2f/CBWlakBSjcFdHmwowU+mcd2UYSVZ
P3Kt3FPGofdcdCjaZUxf84Noz32zFANVi+tQRAnx8BNmz4hgquG2/4lLAXefPItQ
P/jRgY2lQvZv3qoi2pUU+mcRdK8ay7FSPXsoQzOLOtVhE0qj7LP42zKl8bs/udL4
qhEffNMfy4/nX6kDSerw9eoTUjdyUtoR7bujpqCGqHPeYkUr60lhVndHkQKDfWq1
QkYZ/SRc53rotwNY9bx0tHZa8kSrD42R/SfRri638lr/qWqbfLbv5cu7zYo7bIQF
z4T6G46tN19kfpp6CGEfm9HrnzBNYHRzkpGryTpjwhorlSgVynCCb60hnKfBPxiE
014ExuQHlDjiMDjZrIfN0rziYCZqXmZ+lUMa4PU9mRsrebZxRcEnnOoGt5rgT3c8
im9oGASxJTGd8eCabWCVW92Tv1ep/NKPZDGVbWZVmmhEMASkXf/lIoUokZwuWR9f
GboHIUQk/aypTVzXLLov/y2jULv+9r5gRKE+G++cNMNXduvr9UeGlqu2w2xgutIY
4M8IJMhxm75lSuTLKeuQplheb09tT+em+m5JRpd35j5vqblglf0VB+WYQW6eGfgm
I2fp15KS/2ZroxrNhFy1P3InHb9Mpvy3gqBhbNaK+b5s2OVvTnK1crotFBVhw0o3
nks9QkHdiuKvZe3HY4Kx6Kf5EjpKCZHzKZLpRe/wO8GSfhsRHE5TEIaBFvic+Ktk
iKESNQcF0EcQZ82+s1ruX0NOmZTVccNvCNx0taaQJ+AxLp/srdJtS4fgNYjmThJk
bSS8UH/aIERIk95jKLwERs+kXjn1J3/XwalI1nyfkF6TmLF82LWIj1PwNqP6lGJw
qm3bPUGK808LqxIPSSiKsJOdZXtm/7WFb9P6KDGup7WuWoXEm3Wn0BOWJtF8uq+k
NH+ZqUW+87GbLejKSp89oLRHeBR920uDaLHvrZDdE+GxSachLEUmzTCtEDWEDv8H
aKjnOUEhuLlAQ5Nu2SOazuZJoRC9Er2KVrCNzOXZ7zvTl+bPeOO1aONTCTecbheR
j8tIutLmDYkZbhBFlW6xRPum9bUK2Rv7uMr01WfNv5UVoQjWNPYG5cLdDhxnZpgY
V9ln3+znSOZDi3TtirPJtkQwXRQy0CkciK4XRJYuWWgTN3AIMGfZT499ti6Jb2ao
3KKUfbqt6MnBixCUkbveZTHKQjWoOVQbPhTmwc+Srym3O+7MHhxLtI+5rQu1hlS+
75ecAv4uekDsN9v6ZKJ6Q2Vhk6zXuxPPbfq2Oxg1gkbrlQ/hLps1U63Ac3+7WrjV
s9BXMmumoFqY78uB5kCedkmW6BAYCFRR07U7BO16y6fKerRwSGODC5hR8SYj+ibq
HNfjhYQl2RX/j7KbnnH28fqpLZINEASP+6MfGzAJ1KiMzYDViXf4r0CCZNF8xbqz
4+C0+7M+FOiOxo7WOr5dszMVT2mS+Dgm5+REHtJF770Zx7h0wWi3EN2Wd8w3gO3/
bPcV+DT4g6cruvs44m+4iuNHRp9+JLczKjXN/ib/spv5iyxTJ7nin/aeR0AnSpLI
oOieaRI+jOfVnHZchuohTMGAImfJpHhvRHRXL7trgj6cEldcHbZshWQ/jPlJq86T
LGE6R22G2kxKCnNhYX9RugEqzvIr3V2y0yx8gybIWudGQx2ald4wtLEFJ2qg2YgI
WYSPn5wrul7n1W8Hj80DXUaTfaBQskm5JMLq92wyyS3syw0CLn+zSDUN+e/ctePR
e3DrzEHkHA94vOHvFwg2Ol4cVCCyO2gipSsYwN3k3ztupNkP2tE7ksgYWJ7R20Yz
8wGrdSs7PzrS+qsTKyoPFz2jadtJWUQI+wKg4Pqo01CyedtXXYnyHA7RKpvXYHfS
52a4iijn1AwDENoQWK2InyOPxlvTlemw6imSwT+itpq5QKQlaQ84i+9OyMZhoa/L
MJ+5+s1CbEc0qP1izYLpbcb6+jzvSgtlx39YCg342jUFsfRiXecvAkHjJkukefPq
0h9Uq1Wa+Lv3l3iJXoq5JbW/gl3ihpCTTQ/b/l1jp1HTlDxr7m2xnFRcVV0Gg2on
dDpmlnqfsmRzuQ+27+7u0NLTCsf/gnnGWu75mDxeFhQY6UDkIanhpGa4g74nGNpE
aMLCsu/+b+vSrgBdXQZZyjpjMTFLw0Sj6/wx7Sh9GalqJxk5J1cVh1az2B3W4TtK
5sFQgXCaiOcbabWooul9UJa8IA7k5Ka7qYc45h6AH70e5WLmmo/1N7XwDJoqMI8/
dmCTwAgkKyawK/nbSTyq3EFg0QIJ2u1PX5SrWPD3Ixrjw/uESHuKifaX6UHcfTGk
rotBl7SYDC/x6vPUEVXH/xl8ZBvW5/UZO11F/H54iw0uiD9Ut64NL2b2uYZuXC/j
tBa2dyb8sRuO19WotDUj/OXV944Sl618jaJ84Ts12KZGkdj1D+eZxn245DQRDv/3
BchmOQLczbfwrmhqF+7hxe6MPq6FOk/NOZt4ky3OJAG4krb9483e9EQOH0FU5Xk0
VWKeemq3MpdnUvSPCF9EIttfOZb50YnfFG/DmMhqFD2hZsOEbd/TxLSh8UjckB5E
UvtGzb/J5d3KrqCEnLhYqjplPiEsSTGV1PJTBwlOjbbINsqSJi7bCuyOjtSWleME
QXVlvvJC3f2m+ivaH9Ppo4p4eN1G4EYAVEVJ1g2uhiuW1B8DOykNw6tw9ix64epA
9b2dCQJqnT8W2ErySL5kkur/d9Y2/OmIsBLk9ahAcS7FqScfJyZdAIOR6BxlxD7y
7IfVc1bZBOXKUENx4a8qO9RpU2Q/eRydEFWQJqNFENk2LzCSmKWNZ+79U5EWy3NC
cmq8XYrFyu9bNGik0m3z7lgUs+rTTcuna8tTJOLMvb6JGh2wQRk/Qc9i/HEjQhT+
+2MQMeGTixFalfp6tYUvnwDM/LfSd1BfP1yGWd5rmOVf6m3neNSf+uadSC76uSPt
NLs4heV+Yya/JXnup9ODIY2nXcD8ENor7aj4ObYVuV+pPk/Vb1RA2enumuYS53Vk
rPhaf/KsPOwsoHebYXYKqQuK6764iw7t95FlpFfjw4q4u490P3oPXKKr1XmpXwoY
DrJbZVFPZG6VHA49+zGn+L0J13ZHp+sSP24zSKTRcwDV+HO6ZijKUBR56vwWVX7m
HgHXjTRNxU10GkG3RkuEL50IZ9QLGIkSZDtvf7JYra/npEjEfDacnx4jZsWRyLhM
5DTChYyomWVaEjVfqBg/kj2iQ5U/dtoIynUh2/ls0D0QgiS4scCz+oaHNvLaSaNZ
SJd04P/zaFKdxBNB5b8AhfCjykHMegOhDIAGtit+KsX7QcLEzj0ebW1vN7cgNmz7
yUjMT+8w1R2aeZENVzQjFMQIEp2Q3RQoVwrkrQXCO59OiwjyTkr1/3IM/hvUUNAk
MVLUjmV5sTv7d+aQJetdH1ul3GAA1eycrOTwnVfMe9Wh57IJEG2+s/SMWesPRQyY
98ZZr8uZnqqa6n/AR0/3JZnfkkipuOGFIOGJIUlYPz2fe/797NyT4KmWA1DFGG9m
yFD3l6Z1RFEJkCT9ob10YQZV7wulPShB09ahUb5prXC/xdJ6uUK48bIVkPCFuzoQ
IcLEgmd2zFrsLHImPSr66Wq3RSpJkyYR5WegbuFWfPARzbBERjmHhESGSlUh2Hyk
atFKtB40j8zf5Z3kh77YGq47OVdvexUglU9eYuE3t4rb26Qckq+GGYbb6Eeost2C
fLhVWgyyg1vSZ+350fYMlNW1k1o1EmwGObR3n9CT7gnyf0+BBUw/Fo646ZbmtYnM
gafqQdeenNKi+6n9zQsdUYjJw46zkpF7wsFMNGhJ0NZP8iA2S5EiazKucJWv1eIv
uycqTSdwi1cMD5vr/7MgJTmygipENtK26AiKfYPAagC0n7MrDsHclSH3/PnOPSdr
NH+h2OJhlKZOs5KzUWlUeV0r14Xp2uuTl8Y7AuiUkDZndUsmJJbab/JvqaMIxgdJ
hvdB/H1IVMpQzz+XDH4geXvB8t/NLd4Y19PEDpAl/JS19HRZG9w8+aEZOwz9KaSH
VCdBKOicmPqC6rmQmS4gtuJFRUXcozUaW7Y6IwnNY0pdnxo/phxDywnWI922Ffaq
OWNMxI+KpbJWRquOlUvo1CAih0AnybBpBCBXV7dHr07KwBR4AukqKnHMTQIBlr71
UO5BedNpR3Y0s7AWJnIIXbnu9Ym4KWVW1/sQUXqWccqqbF8S8wVCT6IcVRF7N2M8
8OZLkfzUIiiK3R27Nr42T95ijyUALrGLbGA7YiQPPP8VkrGCkGtzI7IhSwy7rjBk
tz2WMaJMW6sKDeIvvEuwEzT1iOIzqcYFptL0hfuF5y8yFaNW7ALpVi3AWzVqWfSh
aiygYAfSzzl/W1AJS7wQLy45HcoAANMFADsvuisGZJZ6E8fKzHDPh/Pn8UPZu3RG
Un3l46GuJi5L5eCQ4N0L/ygucUjNVhwmwPhG4U8YwP694ejxdo/vR6GTon41LGFP
3LWimfqYK4TkjUNjh3zadwVcsMOh3SuonuKWHlMNBl0fHCNERoC+K7dx56MX34Rf
D0dAnOJu0tYkVcMd3pvbBPS/qnNVRlghP8cdhzdOrNmcuT33MoiQskP1k7qAEJBA
K8RzC44vr45d1axYBE8pZQ1fnaG1ZpnA15u9sYu6/Z86hufi9Voo94M6X9YcWT7w
9k8qCPT9X3OziF/h/DmqNdCvOouwd2T/j+LXFHQ/rnKR5Ka0jJWtMVTPWeWSwQEU
3AyBewuFtcwPo1DYwwvfbY/IVo3uBzOu+CZfFKa/Ldklb+ZDzUPrrZIfTXBG+B2s
FA24WzmJnuZZN+6Adx7dbWLEtU2JbzapGEcKiev8cUIlBkd/SWsFjZ0f5HgAkd+q
pqg3qAlIWvnBsJJU/h6mWUjOiU8RsaNWsnqhf3JjSVOEBu6G+dLDn6IpS4etX8o+
a9XXu8ngiHi5nEg5fj9f84Ew0yY1y617HONojJuLhMrLSbhCsRRdl83R8dPp5AVW
VtgP7jQN8YnJdcb55aOZkQGCPZQjZ3JRWkWa7Zmvgt3QILP/mZts3tVtE8eOgNqQ
meAkCuBpet6RcB0VdhRBLI4f7ve3w8t/A+gRRAwqcQVHEp1MQAGy69opeYpgwTAr
1+/lxMqXNs6WnOqGXFz9oGZnJuC1X9qNcIsOnVlwEmbsN5hXHLZWiOqi+mH/NF0V
ojAeSRo+u/Jd6kL25ELDrD65vtlZCsQLx7m4TWVZqPsuUJGxpttLTxmmKHc0jvsj
emFtcrUd0v9BwigO7qy5gybajlvNpdjk4OUkRcoQKL8o0+zQUiUHCAl18UbcK2B/
rXP3gzrJtWWrZg3yQ6DqROVGCSL/+5OeWX2xOcY1xIt7AOZm/DuP6LY91dDeAkUm
W6vZcF7tLSZ8xI2EiDCjj05oQZR4oLzFIp0p13CdtA8wq6w1LI1CVw2OpawXxI+M
vqOxk0NwHD9thJSlwvttE5Pu2wfYWJstcBYevfS/R+6+IT0EFkB0J5eh4Yv3J4aa
P1eY1I5/bFH8+FqoOPZ57k0qAXVmQniZp2jUTYA+1QI63enviU9Lu3WpIqHaAwBU
ppErfvQ2erfOgz3+pQIwwifXsP+u7Mz1as8Kll800vSyyy5J0JIUfJdUU2K2vNft
peMwsJ1fvGhoqaWEAagMZX+gx5vjZcWci6y41++mHVvHQIk5ltM0dqNuAY+PMMBt
jL//G/bfAfI4BcpJGnhHbL/VxfEHv5IMZAax2XO3e/vgktHZ15W2aZVK/p8hJIyw
98mNbhyRcVMAdtCJaz3Q5JMjnE6nyqw+PuZRHmA30RZTMo37/4KdI9SLtNs/UqeL
xa64ygHjCCAYzZGYFElU0MdneYR1cqATp+Yx+Y6dPz0LHR9oVS1skTNt7oY8e6P0
uec6SmD7xJQPuJwGSNqhGP1Bxiq25d3bgaaPtNCT6XkwKJT5GcWBvmXXOM1tbKQW
x86334/fooyqEK0MoQusseNG4gzRHu38kHntAW7Vj0dEu6pYpFYpl0/QlDn+bkSh
ofmp4JB/21VjKSXPiRqeOPZ6HJAl1hi+ugxKkLYKJYo8Iy5VuOZXlsjph290CxLd
PXFOvvNqvcAoGiiCSmeETJjAXlvh8+3DKcv3dk3WO8f87C12TnaOdy9h87s9ZFQc
va6fYjZH9eTlJEuZNBR1Xtyz0pT0qVyofoxHYK1qmVdhMYys6smoLq3nwSuW4JCb
jRVmWG05qtcwBKAnsgbS1Q03WNH0dwuBQ5yIwicrFQD3e/sy1FQayKLpTTyP2Hsw
GYzGuKmJx3RcUoCuVDeBxEnTMUWucMMRyR6or5kFR7FX2mnqNmA5a3dnL4QOUdau
rpfCdMd9SyKcIyZ5dc0XAdg6R2YKRDiutoqA8wgp7vW75g3w1lMhLt5/tNkTlYMI
118sdj18YAKLMKPZ/ZcwmN1WWFKTy1iF48L5MPjIe3v3xpvzv8kObsoSOSgDtvhU
OVUY5cpDLu8ychnt111Mil7bRIjIm7emvmE6kEL4S6SWJde40r0CWu4mzEHCej3T
ut4o0iATCXIpjxoa+CR59NNkia/nH9zXXQiIpJul6Jhx6c2K+NYOsR7BEkhIo3ui
IiDpGPvR5ceLEPt/E/QYUydL2TuhYIB7rPiXxgZ7p/qSiBDUcICZtQ18Wyjz2dsT
8P9+Vq7IvEjK5felZkZ+8RrDg4E7VjwHBIgAWVp7fZAs8ollZktpik7oRO86/C7P
MuMpZ+pA9zLA/8dA3dkDUGGWgPZ7RouI+VsMiQ/sBKzp9r7vqqM9ZPoqUNjlqmv9
ZoqcxfMPuPBgFfDuJ52+YWXvaIFBMYx2E+OyDGxQIjlJsCt+3xbRKQR9uGcFIaLe
qsmVbDpR6nz9y56K+jBfjlcrRBJ9rLFYNwiOG6sXRlV1WCtrm42h5JIjoPMaYkjn
mYDM0FWBg5CwKeqaSAtslvFBw3+Hyc0FK19hDPafs063zUZ9Wws1hSFa3u5Lk4DL
nbVsqjOB3sDZPUfLwlsTmnWjJA40vnQyYkdEw3A0dmv7T/XPkho+fJt+hUzApRgY
w4VJbJnQABIja6xORApMwfOENmpRtDPZc2RlGD9WopfRVtifSlu8olwWYCMu/d+4
`protect END_PROTECTED
