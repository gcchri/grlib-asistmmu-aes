`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjsG/pkF7MysgkTWZLW4h0qxBgIybCLr0nvTqeuvvnd+5wQs3ZjQPv/oId1JPLIh
+nR3aZyP0j4aL9Yp5f/+j2ydWE09ByKoSEaquQq9SNbiKSv7ujJ4k/ZveL0pEaQr
LE+NifZ8Y07/GDWcVYcIHXg8B+FFnUZG7m48vbBCRrTO/Lr0E1xXLUifqAhe7ksE
aLNyrQxtCSOpQ7Ck5MsBVO7/lPa3Us6fzuPrYFs15D2LZINSgOd9mzAZKr/VZZA+
uCH8hZe9QX2XVllnaHn1JTYaUDKgH/3mHz9/b+jIje1db1SZ5vPpoU1Lr1Tzqttj
aBUHmkwEOefCpk17KMvWu5Z1GWpJpkQVmc1HQFy7/uIQNqzp+lsRZ5dGHqtNBj6B
YDYo6G3tIzhsA91g/qsBu/sck9teN1SxeW0cH1gSCAz9nidAPMGeihiNUzccqNdw
5Ds7upQAucbjxF6F2iFEJU9SbctAOiuwsoD4YnKK439gCtey9UQpHQEBIm57mAr+
4aBkIn6kuw4JbO6Vv++3hBJiHUR33zfqyqs8dQ2RB0zneh6SuKsONWBzEPIzPgjy
FT3P4ImrCMegbFifGBoW9OBi3DgZ2R5O8vwTaB6MHJB/kCJUuF21WGRq9ccHsYWa
C8E7YPJNiNR+Yy6D+dYuRQ/e6RQgxa/AVUHJ6HfcXFC6bsRtFVw8zxjubC72gApR
rm/s5W9oD+WwdiO7ObYRNEY2kvOwG1klRVAfd1mu5WJICd/El9I3gm8hqDBnF4r1
YJGATG1y1C0RN3B9py3jIt6BE3ycZKCwf7KI9OBx2NgpX0k1TJFyPykb/cYiM8rR
8S4o7KvXhtzDgPNTOHKAvOuWp1EpzsSi26JsNKBBb4vLyYD6mn0YYegaEGrEvhPR
k4fWOgmoLw/lV1vFUHA+aQkp/w8VMATviwsL+U78cWmN5dNM2FxMTukKtMduOc/k
`protect END_PROTECTED
