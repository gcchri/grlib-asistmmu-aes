`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fSIrgK+pE8YJfI3f3FRmsHY/w3zEDB5xBcsdxFP8drg72F0EBbVkAx1XisV2+zmz
5dulGq5lcjjz+5Mgeyk710Ko599sRI6Dq72ELZxxAy2e7MOIwlD+vFeJ9ffD9UgU
7jHRDETeddTYO5QF4do1FeOGqTQwDjYReA/OVJdb8VXEUBMSXEbdXFR48sBnm9NN
fkD3TfGe1bXF1WQVYjr2D8X61cPRhoxa0PE1Y7SGMlBtCQgCNb+t7nAa7C8i/RPm
haJxm1LzblceoXQcaoWg9Pi+AL/y8Dk/UgG/YmuTL8z3NRbYxL0GrU+RtkL0ynjt
IwpJ/yPzHsButYqJwHqt7LXF1V7V5qv9MPHRrUO5ZTwoDrM+6Rda5VuOwvAqM9V2
27cHF13AcMZ/Vpfd9EfDActOGa2i7IEHQo3+9TnszFoKmSsUZH2hgbCOy6WFDW2Q
sSrW3Z+1Z+iY6uZ5iVbO5yYKW49jR7gw/9/P/hGii5Y=
`protect END_PROTECTED
