`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMvNTHhNw+K4Ni1xC8spW0L7mEKHy5B8SnvwaLQk/9j0KLQUOHTFBCCnz+ZLrWOo
md2TdzDCKJbyeO2KK2RZXOfxeX3vpiovJivgrP+gmNPc7IUMs89hHnORGiuyUd0B
JdXo8XJB5fHwhX0WxBXmXlo7g+VYNchk25oFtXcuvCFI/53nE8b4LwSFLYQmmhAn
pf9Qn3iHzYZU+QVgloticaSpsQ/Y9/j/65aqdjp4bCeVCZkk//hgA1XPOEby1lKN
Y8N5pFxTWLcENAEsZiCNtNfxxGXuCxkm3xTujs13+i5t+Ik+1nNGTUAazRCOY7os
2wD8o+Rr+VaoIATbkTAnN5XOAgHe5vHYYjc+Ei/1t0qSbjUMcynqCLoNWPzqThtS
Mx2CWUVOEN7YtvefjLxnE9buDparOQH3q3NkvB1WKVzIs4ZcBXtmOPB0hDZjRuO4
EC8qyYsv0587ksxYau5ZuF1CByYGydWUF5BCtUqo3rfmaLaHCFcERdcy6ICkVbmi
5R3MtsKHdVRpzPXbTOvoknBbTplAZGTmsrXLhr2KWuP/NpPA0mF+/UCYOQaimqNO
TBOSQLwpKWEehqoOo9K5UO20n5tRXJbfzxUKPPs6m/ZuLScfdAWwOIy8drB5hAjc
+Q1hKORVYpm0ya1W5WhvQvVbS64jb8rw3bXNj0Uxq7KcV0t1Mkr+MzRxfOqJbbXw
oIGXhZVsKO+2EdBSZzU3kUo9md4MJrGBIqjeGXkuDmoGt5Ne0ExlzVZeumNyqVmJ
`protect END_PROTECTED
