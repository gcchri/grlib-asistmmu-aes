`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGqRI1GJi9ne3qrCtoZ0GPkkNX3bRyLl2cB5xPaD7sin6Mk7bTSKIBrbgq3fe781
tDQz09AYZqJhNn26qoCZZsu+0nQHscYulRQS/yL4eZ+gYR6O1U6Elr0ywrNgztqR
QINZ/GDdtK/iqi1A9jwgZq3qBHdXrfnU4L6F9G64Y4iAWjQZxksj8vOgbN79O6X9
lca1weAMenUNi0bbPDR9vfwNtVoCdE1DWwO8Kjv/a3IE8shOw5uD9J34StpRGJQ/
m+L7EYkrgBoaI5m0VtQKleBMDBHgcU/Z0gn/F5OyOqt/FfnTNhO4DIfDwN9Sbn6Z
MyAsn62BZw74NhFqVz6TRFRJZCYQrrC102Ywj59xOQtfgDofktTIsGSsmBo+7tZ2
LZTXgVax6zY2Ze1Jj940a8bbmHwZCgHPbHU9ZgjWL6S1lHK+5I4QFYt3kfbKE7BL
zN3WRKXX9uabgWPBCmRmT0apZcA2OTPBTtdzoICUCvV/lUp+sjfIKeRAK3XI692c
3aQ59z82zt0JjL1Om71h7D5Nu05exJ60+abnr1s3bA2iu5V4wXyiPEWBqZxrrz+j
4C6Z6pNlyoalkD7NsvlCWrGXbzP4tBGcZaFHCZnn8d2JUllPpUMkv56gDEkyKXg7
OHL6TjRiZAmaYhaePmCGEXkcv2yWqLb21/yjYyHJ6O9WX5eX4R/na/kSjyqPjyY2
For+Actn/NsXmCKWZyD8RsyiWyN6NRNPc4EcQDY903snDO3BKn2TPALMzCrlCGGo
cWhxnESns6Vwq+8qUyRqP6ABtO85a2ZcSnArSj3tdt9KqYCd+/scwPY5Hqb57fOJ
vxRcY57i8AfIO1i7GIx8f4lliusg0pUQabbc2YIlgJxpidziqlOkHCVz+ohFjyRX
4w/AjwEUbqhMjxR3hyLWzk0KJiW+IEvnXRBbc3ZWycEuc/KWyKWWvHKS1D6I/wGY
UakJ/u8b/IGK7rAJFAj/faUcJYgwOhB9gzvQlobYx2ooWiNma0dPNCOaPIetJHrX
WiZkawHTSNefl8sxx6GadXUQM0wKqFq6QV99jl7hL6ebmo95M5bvujtp5n5yHnDf
WPki5RwDXfMFuj6vJW3M2IfHAoAsvAyXt/9AVePD5VkyM8Cot+cHwgtJjNPPcN5J
qOUKBKqlzIIvIllXdWMQm5osSM2ZZWQudxFeTbV7jb17hxDfPGAIvKSKW6bmfN4q
5ndSKNFRQWSQ8VaOg6KatiI9GT/N9eFp0qorP6JgEe9/huiu1AAWIBC4+QEH6Fbh
xYgUYlB8tE9jbv3HQAANVaWKPuMOYo0d1xxRv1bGed95qelLx7W+osmnO+AToz0k
TvtxTBcLWD0BXAVWl4bfi+Id30ck/58tN3uA2HyyFV9i+Ww1u8b8BA9U85gMDtmx
R9lIJx128SvV0/ZiH0MOrZSFUOsKFzMBaXMxGtR1eVxQu0QDOOOQ8P28tXNn1OA3
GAvxEfA48e8n0LY5Et/iv3bO6xA6OTNrC+dUyR+th4H6t98VEJVbC0kMzyhFq9YP
zRjle5Rfj7F8e88ASxTN0mE2gRXDzu5URg2ZyXFj0HTJiLkSLpL1LEscg0LiOxMG
OURoo9CEr8q1NmExYC8vb2rNE5BIp5CgqCN14aGltHJg+RWiKAM6rqKOR+1rRIxp
DFFBDJQ6qn8gmkKT/Dgbnvrv3U7BsUSnfNdJlWqMgaZnrAGTUdbrUmrZkvjLeOYS
Xej5uag1tv9SGK0sx5LcJnHh8RdArDIzKyxuqUd5NCzGMKnmXyVzqir6ZXlOW5Ye
Q5/R8ED8336RLLXn4SCCRcMIgjkzYS0FrFjvFVM7+oyVPVDEOa+uiWPA7fvJJu3n
N11RodSBBJogHmq4wBugALtEhapjWrM47xFArK/yvTerhC3o2zjEkuVq6VVGvQw+
4As8sKZc1TwL707Q3UGuEt2rPN7qq3rAUE+rPTyLcvTPY5zzx3ahmCaFt712+RzH
mwv/O1YF6Et1eBdCchb/ykZLtaeT7eqVLHcGa10FIPumaZG6nmLwcGMRVFAOATCv
FMn13XMxV3ita/ZNUMtvDINUfXJQ7O1SSKJhV6xxPpB+isfJTocnZ79GphDaVjLZ
c896wHk0WC/i1Fxv2cL+M3uQ3VG2ERHkTz7XtGFAELEMyi+avzqMYRfWm/m+MsrE
1lRNk8tBsfi12J3+MKwdKQ==
`protect END_PROTECTED
