`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k1HjBte+HxHBvdO5X4gBMkw0qkdeASLZVEaWBqkmSLVdB0OHrAUrUqaA/qaL4thu
YtDMowG2h1lF5l8hbCzHcS+42W6kKyg81gCh/o8wxvv25ud/KhSE40bp9w3RvDxN
oqOPE6V2qViaR5bHwMGkt27rlh9CBNyJmPJgTT/Pq2RXck9IYt5eQW5pECeWkn2z
k0PN7k3SPj6gpAVGv4/bVe+wvuDAJsSuTkeZBaMbY3StwJYbPm1np9tYSwG2G0bU
Wgahdwwz6xq7L3TG/kwPveliyXLn63Spmg5x2XO6Oj4ttmYt6m1dfi3eZ7v68rtL
7FgRsEY0AgtAH4BFKrgg6wOOJS1UonzG70SmSzz8gC6cmZX97XLqVSNzyQUYAX1j
bzMQl4bitAAqz/m91Gu/2Q==
`protect END_PROTECTED
