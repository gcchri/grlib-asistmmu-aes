`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yMhc6W8eAvx45uyJ6mLlcmAo2p680g05pQmGCtua/dltlV6osphRNm2G++cuK4UZ
MiE+xwrpz/wBTtwzg835jdOVww51G7MrTsDCUvRaodrkfLrhHksb5WOZxaEfbTQ0
vKemmMx89FiE0Nr59rCPw3yynBlgLeQjo2V/z3e2zJxVQ+d80qbN97dlC391lxhx
tJQbKqQI6UXoSYLZbIMwsWXFngeDjkwrcBi/1L3NrqN0M3ZsNvY8cNKLVO+OETFO
w+WaK6BYrVQMufksobApxD2wtg5yZDTyV2PJyJvfQY0GhrewxXaMauOXelGymo52
9kURGYLrSt4rOrVDWU2wwh+ChkT/EbTwzNCwDU2mvcCj/Kz291BTVR7ECuNSfFQw
UoNi2DIcAmqE7ZvZ8B/vpxabUEQIWQ9UZLolF6CgvG3MwWP7HwpREqamtyBrtJFp
rYG9Fbva4l2BHv+0SLRiIZwaDmet4uJKWp8wlLAKHfGuR61duHMkUlOwwiVDa0Fk
CGXp4NS6GHl5v3NtDkMXSaEGGICwpaEy7l9sweKuzNXGWcSIPhZzlgA6wMH1N79j
Qtg4wZK6ZbQUkf9TYI+WrZrQHlda/HVXD+9g/TmBk/OF3pKXZ2fTgxfRwkKbKGuH
MPlIs4qp4ENb+NQ21uv2Ttt1kVmKZxvQmp5zanyvaZGxLG7uDcjmi/Rezs5sDHd5
rUmUSLINnv0f2+KwdsdyjPOVnSAT8bMiacSaUe/jUUCAWOPvaoZ81aUE2bOpbERi
wlhYqXxGJXQhoDpylHs6wg==
`protect END_PROTECTED
