`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oX/QlkKeOIRfIZ032mH7+HvejGUFM6WGu/B0vdDfRqaArOs5ELHmAnXz+adYBh3s
ChDU0WNjn4qWzmsrThEeuxBKDvYP8WhbtfqoGnapKUYiGaw5490jXbpp6EMk72nh
bv7WoBr0B6lFFHGVGV2lyYZcubjUv6Gp9UpqXnFQbLgzyu+QMy3/kXUNbAatudAb
bnaql3BAYPSz8cGNc46eXZx+WLxG+MwcMeTF3mcIDmpLwJCDOFZU7RcCDbS/vkDw
DoGRqRuHkAb3ycxIdFNWpW2mpflhzHt+Ods4lckOHWU=
`protect END_PROTECTED
