`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LyLcYIdOn8hrwWWe8B2lvKnUBtVCsyJQeH+HFujCZaI49Cj9KwT1ILJj/n5JQBuf
tCplQ+F0Ce5Hz9mMo5kSYyTW8gQ7SnMCmJbZEHF4GxVKCGE7DVAAUYrw0uouFZFv
X2GPagMnZPpxCC0g9Plh5G//ojJW41rVAx1LUF14BUbc1fvISz1110jrkPFekb9n
24x03u74gUXA4Q0nQ0e3IW/eOi+JvFe90gcauVbrZL+vfMPm0lgGtwrGQuDJlXHb
Fq5xMyB7yXIfWt8nnVcffUHnm3QP2pzUHB3EZXFGtQrl8mQDhM3FgJqFD3ks+SzF
YsMzhMUXfzKZ1klV/AaUKw==
`protect END_PROTECTED
