`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0OP3I7e8X+FPIx6rR1+rZyVsJ4jIg54VvuA9GhTf6xDdGy49Ty0LPdyTMFKIHq1
/xCUOU0NVy00Hr583d7rK6KjfglQQhbKlYzSLK9cFPvwZizr7UTrTpW2Uw15iNqy
+Rzxnf90I7zW8u4bdhs/OiuLpbLN3t2a2bYk7bUiYo14weHAxPRwzgpoicd6Rzz7
5FUiOK7C0AsbaPtwEclpykOpCRAOS4jjd0vZ7CeZt/SjHCtajbK8YVqGneQbpNwh
fmyYrBrTcz2A2Gk7evs2w5nEmD51HFMsOaj+h+vYIsr3vLqjbK2W+19I0RcUmRZk
6leQMTvd0ok9wseyPDGZJQ==
`protect END_PROTECTED
