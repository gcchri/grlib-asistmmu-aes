`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pd9TfET6sLNr1hjaj5ROri+cAYgpHJd/bEzUQ0dyh6hZCewlPwVT0f4smklrlflL
tb8Ox3DOE/RzfOgE5n2unnFPmIIulAA9wIU6TC/e6vaxXdAXwOj1iuPgP8Y+Vh+2
9acvBoOl6jwn+BMXT9bcFfxgkF1F6NXvdTBS1h1xcG4ewwnWB2CWQW83QJLs2kXq
pz5/SB5Cm6R2SxVNzUbLxn+zIFB2w+hP6dhnxTevsftwSaIUK6PbisCJQumfyHOQ
DvXOzhJGR/zmdmxedkprQ09vg2KmYHRKuOXDehIcjrTXaM3m00mHpHDwFj6O2OjB
NDOPeC8JLLlo6Ep9cl1oGKPNV9HOhshz1G7ZnJWmdhkv1Ls5nAwvIScCrP5MjbJQ
msxzlKepilCRQ/upBjYRIgCfyWNnaFtrG0xVpgwooanG6gvzTBAHbQd4twpHSgBV
wiGF8bkikinWuOS4WPCByCaI43SKaacDiL0aLBffYQLL5lirY/Z8RAXME1rN1+RC
hS//eYJiZ80uVeYYODKVDcaH17BUdZ7Hyyf7c+W+oEyKqrsxZMwGboZ1IHfZgJVk
qWBBx5QX4rIBtX3ytZslr/6UT2j2oV9nLLgpj0eWrU6K2ezLDeTvF56F+feZjIpQ
Bfih0pELntBx+6DVSLcx/yCDajXxK4ZkNf4DlSOoH1+kW+LXKn+kUWby4L3RMObO
oZzgpIab3yNHlw6H19KS9rjc7IvWsoC5Pi2BNBSGvjb/Y+Ger0XeXfBvyN6E9gmK
5sVoeNroP0XJ0AmlzAgdkdaaV1UDdP6KqokjgE8eNEWXHy269lv9iW5VuNl440ni
FhJnUOpDLbC3Q3rN83FQUbWr2V4G5NmKojIbeuVtYL9CyP8vL8fYcVa8fyr2ob69
l52P8zkx7Mj+dCorokle84HDA7Sbbaa3A2WLntQNdOVzAsS+54dpqKuNwFiv/ah0
ZRHLglLsRuO4ppZia3rjPXz79hMFS/b+L3kF3wnlxBY7c4MnNIWuT656V+i3Zr55
5gp5vG36e9pVWuOavw/YEHfszRHQSPUj6yNb8+s9dtlbHQkH2mVWCDUk3Mlpaoxu
MekABG/J880LEdu1M4e/yTpP9imK/qwGZxbrlZOiGJb61G1/nRZ3MKimhYqHJa03
2oHJzHCHl/MpJzbjtvFQNAK9oyl5IYTmM53n2Eyd6m0sE96GIeOk3z+3RuLf+jKo
GW0du858j7l/uuGVvj5LEVwIeu69LLqKotIKjJ2cocxVFxmrcgTqx7THSsiUG1BQ
MNNcyGG8lqxhUcq+X/LJpxVoHtGMBmQbo0mqbbI6EqKouFof1Wi2prWT1jH5LGoz
rpzn2nDFiTe35J/PPm9QLBK1jtsJ6HgZDly9EdwCCAc8hOs6wwM7VVdzXr3uSBnR
xsgBBMnWlWqn9oNvK2j5JlTTExmW6nFmKyMWFota6+ZvoN8N/lDTV872AhDRKYKG
zyJww8Wmk1pGI3CJmabcNRTmBIIh8CDIhInxEsIfXU78YACRadDaETnlhiUzhSFF
8SbULKE+mTSFA2leAVQIbEVeHW6u4k/2Zk0KYr9QZfEQ3RHlWddcrA902qQbeQNn
yANLoUO+uHor43vHGs8hrqJbXCjvqAllQqLeFg9ahRArSoWj+W4HT5ZSigygnwD4
vsJyAhId98QuII9eSAP7QL1w3r9h6EmH0/R8DTxre/XWxslhufiPueD2qZsT+eIi
dlWcf1vZKQnbdUjj8+gVBsz2J+6CDAoLzRX67qNkvOpINJHQiTgpKhAJPmKjduDz
bnz+PJ7EV8Jr1OQvtMjLisn0BbXx/irHet3WEyrge/EiL8GOvWTQn+eOIbyD93pi
fS/tVCMwU/DzBY8DpQhh6jgVVJ5Xz3h6g/wZS3W8ZxZs+sGGuD4Z+uiydLnd2qgv
gS9SkVrJ5wnwThKsrGEMHpd2vgO3zISFtbCtmDTemjsTrR/x4cjg0Qt9FDSW37mU
n1TJ78KFWNy+VhrA3p8eO1LtVqVqr5nksUDXmXOd0giNNs1CulIAwbe0EdUiwmfV
OYx7pjPqqiVdxDfQRbpIMAmvlS+rTi0a2ZeOFuCECCfNNb5FX8vZsyGT3nvzRV33
whUPurtYbt9PnQYOjkNjG1/Ly0CvgQ+qonCn+5afhhUS24Bk0/jBNAO+tCzXNB3J
GavCIb35aNE2enmvImq3GIfHXxZ8UZulJOLfnBgORH1jogNiE/5nhHGFSnBoufHF
qadG1NRH1oOddSMfInXThFlcblH1b0SifXxhYK25pil24SG4YI52i5SnysZAqA21
Q8s5OPZ6zSycYoflq853SLiPkCpxrijPHtFgDrO9G8m5qBGF/8QiKB/IMfqGq29i
SSHM/vG4rSDen3NBe5f6BZSWmMAFfmp5UKa7qjXwaljEXm/KciHLHvpAidJLjN2Z
kWhTNqd6dnxQ6xQj+kGIDldb6RSNvJfeM3Td0Qtm8VhQEb6D6lXDF6uZydxEdJte
JZVBnqRNU40/RT1RufFfGBeLWQZev/EG5rLn0lKsZyppTxDG8hJykPeYLXUzyjpr
`protect END_PROTECTED
