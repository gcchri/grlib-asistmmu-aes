`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XuHX6gjmm0Fl2y8WVbUXEYQUmCIwl0CWcBKI1a8hAWj/MYJcE/D5zJbXAEK3IJ7/
8OpxGeJ6SfZie+5W8gEKSB74AdbUnpD3yf1VbYtQ3hr9lLIHeG5OZjo6M8BgOQYg
XOP+QsFSk51G//T/L2tesTbEjE2H3BbteW5bpkXvb5IJCndGWX+Yrac18kaCYNgq
YhL5UN0R7DpBtiPXdIo56MGTJ/kW4zNHHkjVNMxeMuq2LTJxpJc/4yzYTLd2PBQH
N0BoUD0/sTjwzXdfdpcNO87W+O46YnDdfBv4+Z8alfFV13Djoau1Gx14F598eQdH
wcBlZxEK5idwXvU2P/IAU4TBT6lVrBcb/KlJqP0duzf2lzV5fldtbbRmIn8sWO/+
NY3P1ijnw1FIqqlkfWdzkw==
`protect END_PROTECTED
