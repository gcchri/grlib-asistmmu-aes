`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DXBkB7OxwH6TmFql/IuGVnvU64M+dztZpf2wSlV9BYGqiU3p8HQ06zdPq32UmSjn
SAUuYpv6JFcOrRbJuGWYRGkRgwVD1M0vxUKnFu2o5VTOeyXILoLUtOL9W47fNePk
Qu1ZzLdm62vMqsiu3NQztveFK9IVIODzWrxl2xyW2GXqtdMK3pVC6ZpXa/FpGzv9
jxzbUf98AoxS0dWrxxRewHqpUfTZA20/KwoqGKEf4umL38Mct0bNGZUtCiljgaM0
FC0tZn8IpX4jNOH9j526HXzUDJBVW4pFygJKyJSuJxg=
`protect END_PROTECTED
