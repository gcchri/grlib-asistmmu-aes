`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htHkncRsX79jelFGBNyzFgOfc+Bqx11BXtshP1/OYB6OUbDLKZI4nSvHBfKF/yBx
J6LcMRSVOMQXLKB3ZrZowV8b7UgfNmfAK/rDIMWUQrVvDlaZwWW+5WWyXA1NVkpY
JfItZxo8sAHfMvTLM4CVHER+REH9y0vkjFum2+gCvlm2w9SjkzBL0bVrJeGrLnzv
og3bvYfkhjUpvZAphtcxeYVRvGHykvpO7+IWzoaE8bD1VznLgAeYLeYLj8SNgdWL
UBKYmi0OO0cQRMJ+lVeim9TvBfx8mzfBQQWY0C84lyU9KOIahKaO72Kpp2NNqi0Y
7nJO2u6to1N3KfyESuKfDLxkFJxvZ5V/Z8QfwFKJ7JJ+EZj8t/SuTh3jvWPqWcdJ
kt7JEpehBmyTXNgdHe2mvaxo2J5wgpu5Fpj1U0iSdfa4CMy5kS8bq3j5FluNWtzF
`protect END_PROTECTED
