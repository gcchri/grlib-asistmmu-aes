`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCMBYHFpHE2zu0MN4xlWBkCMI7TmXuzHhMUHp9lMpddUvnl7lgmUedToBD/bnYIZ
fqe/a6isldSMI14YvrK2jREO8PMDUQo5Te8z4OD83TTe+Q/20mlGmiV5Xi8FxL1B
Nb4B94WuzyPSWZgYlnjKCWU/TaiTg9BnfAy87ew2sS0J2MEpTIsY20y9Fz57jFtI
l0pC/1ECxvNsVUbCB+v4ZJ0RQPMFONIjpSYA78yQ4xXLX4/jJ8nOgjMGKRllcLaW
+Ku0ptuPlVgR8LaTra1Ut9y+O/dZ5fICDXPYucNzIWjxEue5Q/JaB77wCAPwmbfz
86mhBOYZkrxZsFUNsE0rHg==
`protect END_PROTECTED
