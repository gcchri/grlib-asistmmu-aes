`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XlfUK3+L42i2CjWyQ66LE17qi8m8qX9kg84V57ABJ4ztSLiSnpfCXDA08aYLsUse
T+kLmik/+PPBDiA8fGkN1sVtyxMbdKJUajKZL6X1wjVZlTbtRqtA4DnL3/tM9+8H
A1pnOdVeAs3vJENIRlznrkG0l/OWkkO0SB1cBfwChKg8OpzAiBZp6T2WWdNrw0EM
VQ46TFE1HlsKmVSnwOAm+R03gidf6oa0Xigmx7vnke4V9MO8bOC7v1HansCOap3s
9/BqzroTNDOjakcPKappQ0uDJn3uZ4KgXZmk/A4gR4XQP00KOc+JysHnAtH9+GxM
bfanIfAPdR56I43xE+8CrpvvnHzPVAHvuSZpSg+GavTrCFREbiZyX33kfD9kbLHe
US/vCjqAZqUBNkk2jtSX+ZcDULJGW4yXNfgwIEjUF6ZSOv7MY/Fitd9LT3I1MGQz
JcpJNauCw3xllQ6QfrO2+EPVu1DCnj66gcQbOIasqSaOG+MpCYCPQx4c1AX7k3z2
v4LW4Gkx/trNDTVmbGOxOcy4jIzcySZ6Y22ZqctIZv+20/8JjXa+eMyLNUC0pHtm
+A0kNEhJG8JBgoIo4lunE9SLtJj1inu8ET2fZbUbv5JjXUCRCefnxTgHrplKAu9Y
FehgXusodV2xRjB6uycTB1O6m2XuMCk99ExW1o1H//D6djCIUciMXhaMndzL9LHV
JWFBbpDwJ3SI1Q231uad8fSgeq5vHQLTTxdXbbLA6iTrR2svPxZ2XAzWW+MPkvAl
YVHfIXQ/Vhuf3xKxdcvaw7mpgVHKcR6vrVQ3dEWx62Ng0OK3qhq6VyBVj7rt3GN/
9lgsxzz9KWkyG3D1Aqa/e9vKs6Qqg0MrpBq+K+yiXF0S+DsLvYnnud6KdNcCWKn/
G/bmCbmpjKeKxBlQM83JTXmJU/8bNJxDgsTR288kB/mDuS5pBO6hns2entM/VpLc
GyQ1i0/75PMG/dIBtW5dBnh3qY6Ia9lAx55Kejep8fd1wiEkO9TdmCX5ad+NMXoS
KI13prFR0jZ63Q23efR9dqjwxA5qasqpRONGOobSt5ntrgEO0xKOO7s2Iz5QW/rV
GyitTibGRqTqOOsoYFADfy4jESOL4O8HZRRCBasJimTp4+l5jJPfNnNsqhnpvaaT
UDaDMEOG3pJwNTtavFQpc2CifhozRBG9v5347KSO/fV/pTMAdE8bWvZEfPTCSe7M
DUc3QcXQ7DVwksAlh2vAJlll7IFXRWZQpGmEgLgRbmUzo1pntf+JlDYPQhCffxUd
kvHiJxOVee4KWXPw6onS7VTCJ6Il5M/xN00PW8SlM9AtEyhSxSgHw5FxbaWgivek
rBpKmbVS0y6LmKtoLg4P16BO6nxwOwMHEzr9jlBT5hZOfl8OyZFPzaQMnRiiePwh
gxF0bzkwPUKYZ6ZBTOkgEsmiQdeB6EQueKL/Vjb+0emzAL8b4BcBgRfJPI3AsFS/
3YKGGX7izbqDScYr+6sOjYcRjBAjfzEfxCJgRNKrjY/mQPqMMWM4o+UI9zCnDMYX
J5AaJ6cXblakFjaU1p9D4kdSYpUNyuLP/Jjndb4AOpKlV1vWum4zMqpcT7C1aKm4
QEbv8ccbfdffTKIdZaCiziK0qFAgJOh8fQwm8+6BUid9V8FHmc6YNKY7UKwEombL
DmWGukwpprO6StGVAB1C1IS99coztJjQB8qfba/50/eaT9MRG3mQuqR0cGctflqS
jIcI1ZsEfX8mOlZXgtUcLdrEgSsoUtT35Rxm6kbIoA1vFjm92G7YhsvwB2A5iD/p
k8YXpUg6IZLpu3gAit3jtpA7NDg/NZ0qMcqmC17uisGbveUJd7pkf386m/jI5YpT
9W/CS/i6IkONH90rIBFSPFqWFNGkgjRhiBIODTKQ4Ld46BcsTB8alji2fJr+ZpCo
T52CfOsiCOzFkq4eEPKahB+ItyFx98qSSiDFQ6eG3sKoFvwVnCllp8S+OvhPfvC/
1D8/OYivhSU4fKanpXc6WcdZ5KRiXjBb42vg6QiJLQcaxRF0a/9C6Hm+pOyLjPtL
iyF1JyOoavoQzQvdDTwqahTYnyHgvoTqLjN6nJAR565lmSifZNd/FfVSw65JmTCz
8yzrs9CyxoU7ovYYQ1GBDEqx/LzhRhe3U+VR8z6QKhaCLvWszq2uin+wUoz4BZui
R7hmMJ+kK5rw7okFKQwVrn+Iezbh1di0hB1srsRRyAI5w5VpLtQaw6t4fBGDcHTs
Ws3g+5f3keV+BwxflGW/wokd6kTuOH02xcrNZIQ7NxFAaDKcjacrTDX+KvPvunwc
34ZlrtA2psoA63+CBLKkBEYFa8qf/zLdsTh1bfJbiK5u27FmqNMRaVuuIpC6/0Zr
1ROyYZq9WguCZ9/CVHT1uW/vmYH5NhLkFtqNtSyo9zDa2xrnGUT/3L5UrP4BZk7/
OEIa7I+a+6agViyTm0I29/DIgv6VsXOo11kuykvNi7gwjVBcEUBMCbOWcAJ7hLiH
14nSgrLqmnMy6W0CxX0mepuzMBBe+fQxMxubzU+vVevsf5RtQZYChVwTw8pV5OIN
ixi0lydZM6P0IhoetkA7v8x98JwsZCRGH5DvzavsDHUz+QrsyE6lt9UxRCozTg8P
oafkgW+dwWak6KkpcdgxNl/S7dmOKX3gYxm/O1mTw/Duo6Qyt/aIlO+L000uCe2R
qpqqhKhJ3ipaHj7361gmjXw9xyT+7HCdYkRz/jo+Qtp3v1oMGqmVK3IWGoz+pNks
VL7jwyJ+iLjM4k5p9Tux2BE/LhMsMADc/qwIwuiYWNK+to0MhRIoOKxBjl8lBE4K
2li+CVl9we7WfueBs8iUOFnZ9pI8yr4wdIBWu+JXUlIX/eGtWWJWPFEocRE0m97v
0RtOz3u3/Unhvwwp1ws777QprapFp+ekHKQp3j/tz4fjSsXW1ogkOT58qf3V/D95
YSrTagX1knIYeg2oc1JBYuUmBXUUecZk/0Z9W4tXjGQ3rnBj0hg+oM4Xu5iYXgYW
E2EbKy6plL2DViZh3CD0cVCcTNQm9sWsgAkfKpKxGML7JVghtg14+45VN2RWKynu
fj9fA7hMCCFBcJYnj2j4bBogA+QI3p6LyL3yf6EP75EUP9L4L3p6gZhJ4w6LxX7o
84l7XoJYL3RYI76gQ0oaHyi6F0ZqZil9EEoMKIR9UcCNziLXecO22shZ/In9IgMq
gJ80B6tSOx5rpqpO+BuWKUWA43jJXrrC8Bc2E4GvM7wR8ZSnc114zCeqldjseAD5
DkkQEGkebGHh0C4KlelXAeehuuf2JW8itWnqH6ht3za+UnO29NRIrrWFEjPPQmds
sLQTg7ml4rGpY6ijjZzJRtt3rAkrmftEEGO54iJ3TPTJ2E9hfQz5RhYwXE1fKl2l
rvvpZqqX8/1z2WjI7spYFHQBGYZNpINWJq5Y9LXPmrtTVsVltSQqfqQtuoezexFQ
RnH4z6Bkr14fwau/SoUKshqAwxZMD9q8hIQ6/FzJYvezL6+ctshXwnArY7OLl8ek
h/K233zgGOSIOlcBLGGMF1xoBP++8bRK/8UzLlLC3g9sBglC+E3a8cZ6Pgx+xoCo
YGLfz/HAtfb8eSPYtEZ7YKKwhGr/MZV9xUzRz+zxlkjTDhKfHiV98cGvlpXAtBmL
hLTKDzNaww5m7JmLjVDI/0x+NnIanmWzqhp/5/yj2L1q9whsW6+06WgI7/w/URP4
L31CfABRfiekZdGmpG1P1cQLSKFkMXSATZYdwcD2JUCTrgZUdXOtKTKj1ak7n4GX
TJ4PDatvpsi6rLGx42QDhbMX821FILwFrh9kZrsIJF1j7RNB8fh8Ng3CGUQQ07gw
0K3lcq0rCulq7YlHQq+dH6IImoFJRDfOIGERPEtotfylUAh93YwszJoXKj5Kbl/g
fqBbuCISOHTPB11a//HK9kdiEY2s2Xp6G+XckoB9WFE//GLKhivwmDt9/48Rx+qo
S1Mm3RcGhGvw8tamIMkl366HnO2YFVlNWOH3RfPHwjKDolgE9PKT2DXQZZ4y2EiS
2ZeTwTi7JwC3CxvNhSe5+aDI9slw+V7nVa7fI9dJVbiG6CV/hCKcg4lLAnb5gVQo
zpObBY2U5Pq+aJrCkLewAWj8ycYQWoZ17bNdcpf6kby+hrd5pyszjfmTUOlalkk/
qUI2K4jwKReVftkbQ3Iec6peHZLylQ/7R1+rbS61FaeQOyOhM71COR+vmJo1X/gR
lpQwnXcsL8WLMoehKEkyJS7Vuu/c1ltM6T4ACOt5hMEK+tYnf1yg/PrBcVuGGbh3
nRuEEw4bj4umOFdapjMBdLPwjbY/EXmrrSAhhDHiK8C81YpQDoPCBkYhOpdkz6A+
bEWCBOpp+Zo1ufTTsGWLwdYnVo8OI1ZK7sXMw3U2IooL5RQGS7bE528wjomDntyq
5AccIifezjyDG6JQQhW4HpLlc5FdjHVPWUs2P20DbTiAuQ6BWh32tbn9DTNaKGUV
xNlUvmqiX2gSCerJ200u/eCTaGMeOyoXSgbPZ4fokCe4pjHXb9UUJu1JGVZXByaz
iYS9T0nrYp8gh5d6A/V8OmIkgheSKKqR4FUtO9frAeZaLMqxQphooL13IgvtbyKQ
xnjcTkGm8PrZSvxuRzR98OjBNumqkcbxNoCgdg/vdlVqR7I/fbaoaDeQTaa4AIZ2
sNBmKjeyMhxYpupnZuEMGTPeYZKcg+E/8dKEyWLsuxefKxn/Fhcq18Da86opZLdZ
U/XHt2DHGWzP0w1XEvngiVQhw1cPIoN1F4AuIX9cLcGAgUFVaAYOjmKQAgvH0Clj
agGOaW4JvbS0VIyrLzs9MMJ7mcl/+QCQ5uW4r5xnQQTh+GxBIIAnS8mZMMFwRpcz
4knfHjrC9b6u1F5EajkA9/pcrXDMDl28JqCHhRduWp+BTVxbpTZ9NzbvhKYGavoH
T6TrPy0KOle+vn7VLybmW85kpC2ywHwf5iVwQQqbjn0EGY4tUoviq57g324Y3C+j
ydE3Pl99/MmZSuQ2Rjvq9xYIzYVG0HuO7bYsQ1dYL0+0iCroKneXVf6WGG67DWYn
Q+oZL+Hw4+8xxF7Abl/OIsKEtNBpuRJTj/YYSJDpMDZhfRVGuYF0ltwqaYWGlHJS
tSY4xIBHXwjDbN3pH1CPNgAWYL5Z1Lrpn8jZO1YZCtYAqEwUuIxR9KYeRuNnS/1A
Scbvo5QOttIhasbHTpUc2AiTwcPAlbNyQb4S8SJwKBKrkYsFf1pJJlKFJM9JbhxB
9OsCeLEQ8OW+RwR2pL6m4aVHecUfM5ZH2aba/UonU3NfeYRGka97kZVNf2oJXncM
h3wji3dfwZctRWiOn/8+VhMVF7+jRvS+NxpfftGDMc2cCt8be10FznA1noPbmcMf
xfi2dNg5O9x9DNa2gRykTqwMJMMWtqB1GJCURH3n9rKl5JzgbDtXf0t/DuMQsL5K
yBiQCQIub7nJVVxbaryFbDPVa0Sinw5SsgIc61agfcqDy4/BbdqpNuJqKzMAe1pI
2ge586OM2E5Cz2dXm1cECnumE+pxv05AkgdBDB5/PIP85m5TWRAbVNHjht+wqkfW
/U0FLzHtsObbGpz4xfld4LgZaRBjKAY083Ko1Gc1jnGTBef73Qe0qlv7G4tHpWvv
zon5nMD4CifJPbnj+d9s+/hUAGaDYC0aKk4hKRgG1hfb+kVL7nIBKo8N+8eZyVNU
ZmKDkiyUlwTb4pQJhyJUoeHvmHLJI+3ZdVEPYwbp38/dyB5eTMfOiSANSB9Xhzrf
/g4qg5/ltEG8oSC74IhLmHjd+p+4a+5Vxrve4oez+QSl+Z1Ayl+EJJjSp3Az9D5G
HYtAP6RsWDOHWTHS3+GZToUMcZMd4DT6S+/BbWl+NTv2C4nbIZgosH1ukC8rI/sP
20EWPzbAh6ZC0eLlVLRHTjyT/NFoOahsntWWUdMhpuzhK2saLskvNix5uN/51Zdm
6RKmVHtN67EJa1dDORkJK5CjjNtg29V67lhu8ZKaM6AQYZYS8qIWRoJHFoUUgfWs
91UgxUKZ7+SziCRZcGyDsJ1p3MFF6DQ1cmBx9JO4yJRA+d3DDvo7uwAW9O7xVVZx
g+k9jhmXRXia/mq4tsGz0pg8v/oGZz1z+bd4Z/6nxCI2hbB+2oJqo3CNJ47Ka36I
0bL945MJG38571NgNZG6mlHuFjICLU/YKfBHObKS4Cp/RYn+kpvGihYM6+Ky7ZVL
P3Ui4+RzuOFQ8S3eQ1cpR6vmOucRtotm8LaaaWBB/3GEdgQG9hjQLgKY/x/URkkm
Y2ACTikm9Eq/JUQSbGfnNi7Oc2P7AdMAyNReMVqSdPJ7orI01JVOej0sPKtQ3OUT
Wki1W3SaZdIkp0SRetXR/YnMpwHSkiZopv+dmQkRaZwyVuaRXJzynOfJjGGKoEir
B/sS6B6bjVkQA+fNbIUHIgif6MxEGBvQ8Oqdxqm2PWtuEEaBq7H/34ZVaz5Xpw5R
so5163N6dur44NxtjEOyLx4TWSETX5hclw4nQydGtmEbtRO8usiTLuFjkrRQKT2Q
VVRE+5wvlNYqCTdgBK/yEXy/JcgdrJi2IsfXNgG2hbNmTiJiZ7KcwQaPsuKysZCV
s+10JGV9kkkc4tbpeBNx6iiYmNto9V4spLEChAKgX7ilAJix26YncLS6IBLSf9pb
6FsKa2gMO5qzsSeone8f/s8dOJ6CejFAjpedww5QekR1i08c1EXEP/uvBphIWhQc
lMVYYVjSb1amtav5P/pLwqPApzOWknN6fP/un720eP+I9A+2h7pM8+iQMrK+aCx/
wfRPi4oNVBmst+9tgXwio7sjXBJCrePmwAxeeFwuK86oLCuXdj/zkSBMy1GkeYph
7iExaZ2MtATCAXkpab2Qyfer7v0l7XGZ+QXN+mpn14V9LUO0AsMn/zosH93Ms3Ic
UScSMzB5KIany/9Csjkbutlm2qwy9XDSpdw1OGCJ4Gx1saCdLk2zUrjISz5wN4RK
GsURpt6Nld11tbabLMTacUXCyRcRRN7tKThfbuJdH3riHcKNp/ghH3gJNvtwvOnb
QrTC1fX7CLfOOpr2HTaAO7CK4otP2jfbIdW2JmAlCXwH2FuYN9rw70sYhecUZ/5g
WxiA2J3GwGoxiz6Cof9kd3t2Om/4tzwVKCDjC/i7pxNmgKuFZtHH6vscnoGDz5P1
pM5mDtGDN59NJBGHzuxoh/cpZnGIALjSHyWpC1YBJ9sF21nU3VCX+2Xiw3pmIwDW
1Kt1LCRlC1lNz+otWp+Za6cNqY/STU6++SQHBxk2yqQxU7c0pRQ2VlLCupPMo+OJ
73Wy2Ib+hP3j60+FyR2KBkU7q5Y/qg5GcbraAd1RH1fjJf4meKXxmtBEPUrHLoG1
/2qmjoH978mr9YS4tJMh/cAxV75VtIJNs8iPItVjdz2WDJBcWxz+oA6V3+Kh2TOx
UNB9HpR2NdcqTRCeeKkAVqkelOyhgXOkInqdts6DPcdr+peY09P2tqSnw4kJqAaR
pxnnYaw4yuyA2diNAvSwp30sPpAaL7ouS3Us8smAyPGwpgTW4Wug2iHn9dBeh3vd
Zsdfkj0qLnFhU1wYUdrkUgcLUd3DMb/4zKBvhzxByNnKGkTqw+GPl5z91ORbtxjT
2A4DIHZdiOLzI4U3NOTEj3GiafB2O41vRvt5/D9osssQbXpiVp4wIyPmRS9hY+le
59ADeyV5b33+E+yCqPvFTvQGbDtGdgo5Y/RV2oQ2Me6kkbQsFz5D85uKHGtaitks
sGCBIiWcl/d6YTGmMTMlQCXt9al7wO794JchvIIWFi4LAeOYoQYTLyGBrIU3xlZN
vvv/73QBkDaz5qlWQS9SwXZAnWrdlV5JGt8lYxC9DroeTpHYVeTbeGCmPOddhNNI
zmf+Na4QavFRxLvEf4SvWwXdTZw1VgBWSnGzcOEs1VBYmzPqnAhiK4bnvAaXr8Xa
G41iVasm0TtOiQ8Fv1084XxtWSb7NDEfDDtU458wnIgsB1ZM2bbnAoahyUt3pj9l
XYDvakyMcooGpy4+fvmpNs4NR6hrZRWK5sSuUDcpaFyz7e0dAmW37iYuDqeV02Em
q0UaPAK22MqMi9CX6jegwLsq/faNxDKD5r8woT1py5xB0zoZhN1M15+/VSF+uYsN
xDl3HcmoXTKZdOZSSCYHuMRHPvQtueG5VLM1P/Evc8lDhecwRHSHytdx+VQifLZc
uk+Z3YytcJUoNpBAFOWIiv5uvVWOEF7Jw0WsNnUoxOKGA4eh+ek5HLBi9PFWIDfH
qOVvgYWI3yi/FBG3zM+e6brZFhj2vKsGJwMNtX978apyrHBy7v94TbjxWkL1UGme
tA13RHtlxdIrM5zq/FtAdml+ipBpdr0mF/wKyEaGIWWlQtsEbDI5LF+vRy87Dz+B
dg+U8UMsHkHffPdCX1EyrDekNnhirqNIPskWx42Ll8DsaLhuHNKHpaNdFdbtM7fj
WJWzuAL+Rt5HS4BKcN5PSCySx2AbSvh3bD1v+/KUc/kl/v704YTfryVoZlrVidAa
E8iB/UD1oJujSkOuYkVPunZpUEq0qogAv2TeC26zeSb5c4G7rIAApKx/hOhoL5zx
Tl5crDp0Wgn2fnNs86QNVzrJGUWC1ri2albXJnGs2jeCwjHyn4g9gIbUJeAEeKmA
Cu0GBp7yxB8Sb3amMlu7ndbCnFKGhh7tQQvjebhXDfi+TUPGDNRqEckY+ZF/aefb
PdyPp12chB+zmT6a8Wu5gorr4UsdjEjXmD9DQxx56HWmob3kZVfv/gDfn3EG4L8j
4cPTrTJly1ar+INf/t33Qxwm73sj+1jnZhJaT9roopOfePrTQtHFjE1ZFMOnz8KS
V/GxTnlHN8sOCsIw9XI62xcFfNPQOtFnQ+1S3wnqjPRUOlrUsKLaelFNMJHoMdFO
VNr1C6X8EZNbWsNazVV27bPwc5C3Li0xGfvqhLc6yxz684NW+SfPZ6lHX3tFqqcE
uzxKpX0YKZ1rK9UwlRaSiipCmru5IMmECODva04oQlSFsiLTXZ8IdmfsEugt1tgF
0jqAe9nOV80DPxEi4uEflpGkkczhNCAxaFQAVy45o9L0m4tEGwG0LMZ9N0omVzS4
yyXq47GPs3WXtklWhOoj7Qzv4buuU1y5fZsApv/bQ9K7L7HNI57V3/s2Z+aMQoVp
lRJM1S2rMNpwqrWptepvSs3iNFyohDdgHeZGVNJuThPHinAjOyu+oIB/gVPoK9Qx
D7GXFWRM7KvndqOgJAB8qb3tNdA+RqUTOdbd4U+tkDuhtU3R9BmUCv11UWoEx7er
2hC5Frnui/YnO389QEctGfY8QJMe/qan/iWVRpEfmUhH0G5S8Zm/3YXo5TXZBOHg
AX9S5o9MUm2huY2OwgE2qBbR8RoJA3pf/T7jlRoHZZexp8Y2LigOI+45VlPnGENs
O+X5Wqn3+eQzypKeTRh35kL1x5csesLTGfWNZgqflsNtXMVJ6pKDRWTAL4fI5O8F
sQO229ZUHws9N20ghgaNx+88njxcovTjYo4yPiGLB/pHAis8REc+77jkcZilOU6g
98BsGwFoBtC24DHJoAtOLqcfFXXxP0msFKt3S1ZlHoL+HTEWJW4yaM5kogyI0pbI
Ws4aZNvw5NjpR6T2Db/Pc9OVZTW+x5R9JbOmuIRHFzP4RbohpywDCzolMvN4i/1Y
X457OLUeGCyknK5NfuuKCLn35GqwSUAOuXZzzhXCf4LdOWwB+zVWiTG2iFABsoS+
/9tEBCE9MKnm9AixZSUreWBrctoAwnZlTRUZRmUcr8JnX8YDjgLVmqpiUc49EE2a
lUVmyFxcMKA4xyO5Q/I1ug6iQyB0RsYAoUHd2VO3daUzED+UzCm5A19DqsNRkUjR
sp37QU+LNEQRICrweq1LdOwwqhpTXwPsx8bZRlOLYHyrG10qk4+RX4j8/jcrZE8D
wgQQeFRodr8QxxSEnHM2/ViaxBe2UfMQbyraU6O7YCD7yT4KKZrWNRe11Nps3+K+
3YirxwDsIABlgIbjoAff9vsAExRUp6NSKDLf1asYCL6FLTb7xeodX3DLKRjqvzIa
paR+Hn0ntLbdLtKKelfMhdFq6NeCNUKdiKOycV5nMfKnQpuas1BZMavWhyh/3kMa
vVRy1OpxVWVJTahaIMdR2l3x92RZDBODVcn19DRgR0gCRKoODqB2DXFnXEBpPv3j
ecC+pyOb75UnSgpuk74imBb67XzUo2RaIOa/8pZGPngmhk69vRTO+2t4gvOhYPQj
52X5uGiQVuaAr+B5QteyUfiJystUcf4nbk/jupJ3nAlWv+klbafQFKeYrvJBQAFC
2Ye3yIpebd98lYM/i2+2fJ1/LJuEupObZwLp407aBPcCaKr3O7l5qaxA+yveOsOy
uN3wtoKt/dN2YE6P2bCBjOfer2/NyQNuBG7EEtT088s4bfB5K2K+Wh317dtflSue
3lhKDbMZWDbygaO+Mnr1lEB32a8elRhGUTkPRfOGGTfBYz/rTaTQ7JJWuYAy8Aji
1taes2i7wUykVhm93eQsK1hYtyoqurUzWDFENt0pGSp18ed2dtu85bkjPGOPnxAv
Ogu2M+3AzAR7AkwA79sbqFUfdKx6jcMb5+jv1k/0jRItyXUGgA6ORCqC1G4jHohB
zQz+Egx6gbHKk3B1sE/4k/WOSYkCMdcveu1kfCthWEYEdonGtbsZ7I6FgtEhqOSU
5CIzwjSoZjn424146tco6tugKCoQyPvGgRrjg/2azG6+POw/hRIzQUTvN1sx1rsd
yh5t9ycK1egXBDBUUbtcbAnqhfysrlHhdQtLvGKkhv3sD42gws0p8/HFZrs2bnC6
x8ZZTPwPcOAiLZ/t9Bho13LvDNaleSwGWexlxFvNshGiwPEl6dinpHb5Cvsf5CdB
gQcbM+tOtHw9koKecjkI25Tgz/IvSGAOwlG/G8MJUVRKTHpk5cGbJT2UzLWk2Vjn
zSHtnzYw5k/lSojeQhFhD91fycQL/WigGlS47MlBxKgUEHDjsJ7bvvmgV6G4qsFW
V9Vg+9PoB9xBKYr3gwjIS5g+VpXTO4lO6/EKIqMM+oMvJkczfu2GdIA5G/ZBVX40
xEF4UXkuMRSzFNPjTnZiD9uIH57P+9u6SRni0BkuJ0tzz1STTuboOIoTIlVSWT3e
EkxjQJuQvGeWLcBYuFnMIMky9vjzcnZIdEn5OM0sj4qr8RFd4xNdJyoxOIRM6Yb5
yptBGKP4+dJKgXS3aCekUjHIWxASjKfLMkOn1o16biwns59zSX86kZApyIcyOWjP
QakAgcwbnk2kWWbxekwzH3QSbyud797WzJeHCjVC5o9Rhmi9AZofeyKzuWRdNin5
RuDaUOWjtMw0L2ZwCGQfxJFq/dKTUWhXGwE7I+/6RxKXvp4LBSzURVsE3WO4H11h
+XlwH7Ei2qOwpozu4tO6Et5KHBdsI/zmVgQnRzkURZV2DexbmFJuFYbRTJX0/Ip/
Yi13724BQG6Hd/LM01AOqmTzXTlLJiwB2bQsnKCe43aD1hrnczUY8Bc89MxM1J5z
H4FfJv5FxcObjwg3R5CImVp95jTB0f/7Hh27C+e/miqL8ksmO2xBzcJKnbaYdbsC
l/SoxQYRowxLKzGese58CUBtbs/FL5dKOzJIsEjXondF+/gXyiphybMfkubHZFFy
/uDkX0BeyHBw/+6VNCr8BAsdoXA7GpEKCx2V0yeb/wS5VNZXOWahqlHy6mOG7IYH
tnME+HsiG8Bc/T3fQswe+E46/KzmMA1LeiiBU1JRupXid9NgzLOnjb9DWWDDQXt/
5LoE8kgpacPDGwhaF7+duiogm7205xPf8HnuYwhJPCT6imCEBo/eVd7pdPeXde1J
zxW+P7efmk/f+6xRir/HrQhPDrbgJCrd+LA12myyf8IOzhLSZSoj3HK7ie1m5Bx4
ePKfuQKjdxkD/R9/EpOe5ezMY3GXpYGP8+0BJAgjdu4fudBVmmm3fuDvCKS2qm/9
JNGVcUnEcgXNiryuh2ZxeGgmUbR0pOfAEF3YvSl141mKs3gUwY11GpzOmEJnowI1
ZFTV/Ko1DM9qs70Cp7OUBeCpjd+qKhGR7QHN81NvCBQi2RJ2Q/vhinFGCRGeJO7b
cRHn0JR5mKqc6fZ4CvxwdoK5BD1AUYKo44aLTeqTvqN8/eT9uS5QQwhvXr12tH25
WGRQYXJPGQcPNRIfxIUIdNpd387ZCZICZyQULaxLIfVNibfs9MC3GD0i3H9Z7JjY
Lw1wGJqAip615q8BaRA5RIfvesd6PegVEechWrtUjwJs0u+PuXu9stFobtewnKYJ
f87gsMKagPjpPHCfyQugXOBbh/qaUnKbPmZJ/Q3bLboru0pww0o8T34muyTyER9O
LKCtoaYDX+5JCEVH+oR0p8Gpcfgv+Qyp/pTnlE6UyQBewGQDxRUglC8+Xw3uld9l
xy3D/BP9+EbQ25oSu6dXHD7p/Mq/ICPMWIl4WoNqiOuabq7CEPqrQJz57FlyF+M9
QT4OwjZyfRxEnqoz34lhP5iHfd2XiSM6Avr9/ImjrmGE2s06FD3myfYzBamPFF28
9tDPXc4BUcXiE+akfWQLqEpCUCOGclWhJrDk/nhblryOaL2CguweAEluXumiA/8u
6l4SxKr4MiOLg/vMG/5Ib/3nnyfwq+xjYUUDlnztwpemNXKu6YKtYIwVU4+akpzY
Qp8xBFX30q6id5F2r3Z+J04vnCYqFZYpmuMLZ3rBQYpo/RX7vrpqiE6rUq43+Pgm
s2CpD6u6I4/qLQnoRdh6M8iId815SYbuaozWp5VcWMG9/3zxycn9rbBRoLcrfRXr
CcPBsCCzhr3xLrX49LMbGJvGg6cJ+trT6o/d8VWgmedhEX6g+dM9+GhoKBb2nmka
vMDBOi+ahfLs9Xpmt1UNuYJeHyNe4rNYzbErh2uNY+gNNnMPMfHA1SPM7cb237Ii
PDQvVbR8P+oXlgvlIZ9MkVBp1/Z5qHSEdP3kaNsY1/SuoIavLvdkmj0zaXgD5UN+
lg8wKdLp/9ZXxLAGF4GD9ux+7NdQBHYit1H91KEWItChh5vOWbhaS9zF/MWf33Ex
21u9IoaL76VlP16YH2oKEW8dvwmeenhplNqSEFNoIAS3CVtX6pMAe+Rn+dNpGSi4
GyKZqiVp53CIxyyaNovszWsQ6BVj9jD7VB4/81JGvg2Tlky5JuHM4Bg2TDhH3LyH
Owx+mlLravWE47wEJz2uPkYYDKV3SuQSYxuKuMGgGBPVucj49u6yjs/Fwh2oq7ix
j7vHlYVGwWp2eDE0QIjNavCOB1O4VuM3Y9dqg1d6Gx8ELhNu65vQh+13AfzxDUix
KCSFXX4HLgCHnLkYYjC5ghFCmDXi7C2/Myk9wfIvFTdlmz/pbNTyloV8vrJOS3E/
/d3e5qwY79QvQoavwJ2Ba8Nlo56aEOXU74ksI++Jc5So+ZdcfdZZeOtoz2APmUFn
oeH2om0kHTjpvYNhxnshgqmZcueZcFNFpK5tja97HSdavvoYqYzs/L2m1R42s25l
b0xI+H8vWyoOkzTnyBHd2GqLspCPL5VIAWUjmqu71pMg+IFZTUB1OzQAUkc+YqeW
ZyrcHnwEiX6HkZn+PxQck+DOOG0tDqCTiMrhcZM7ZdGl22+eB9NKEqKVY1xKDgIc
cHqzLD/FV/NkGrdSUrBfvlu2LcE/+cegj4shpZVwneG7ob26q6XE0/4Fq3ZuXZwl
2lxeNhOeVO20LqloALo1ufhaS1jc8jU4X3VF8WiFYZnLqV3vTQUIFrso8qLoWNwL
EK44m6/TOlo1rf/0o2I0dgmdkv+1zpajfzADpx7WDX2D0yKHCOLM0zsdgbeOctlh
i+MMx6IDUoNrooAWOtqjJocmExT9JxDmgX6bi/xk+VA5Wkp4STyfkjH2x/cjjyKe
cdUnS8+u1kcqbRMXgKwNc10M5MZloi94l2Qyee/nXCtaU67HNXdsgLfOTc6FMIVI
0bHH/0vTT7Y25wZP0th+NdAa/dUznWYCo1tnSAJpM8Ncg7QP6A0uMHtsfULnKoeS
hR1TFPZ0D2DZLtodu/U6P260E4ccdm9Z1yrmR8T0Tqphfy4fiB36bPb7CUECer8O
I27O6azR6tO6i1DSGFGsIu0Hbsv1jBf8H1bYTQhRyzzktpBq0rSKBnO8jnk+YMVS
Rfx5tZNyjBCO1pdZDH7saaO2hTDKq0zpxRadyGSYx2cbkDw2DjdifFbDME2qi/+V
gEQAcdy6FzFrGxDSoyyY6Ox1rDtONbtwg/LmaS6yE82Eztww3u0MZAJNico5ld4e
0QKvKwPsDH0ZlxHb4XmTDCfNAhaGw9BL4wveyMEIPULlLnIk7lojr6gRdbfXxBRw
OYHDAL1d9+uKFutKZGBp+LxJMH+/rX93GyKuYKcMaXJJKhaRbMe7ar6tJZt+0aZ5
YqbimdyWWiwcWe+WjRiSPHd3A4/d7rGRi48nAmxFeNo1ptluBBXywulQVEkGYTUq
cHrh733WJlzVBu/VkFckLrjZQdq2iq1A2mhLHN+8ArDcy7FDhCQO53MtC4uAku7E
TaQMQEO1Pz5ZeE0pvgdNiN3BwKfUsi6lJXzPDncwG4t++YxeescE4nMWFZ9x81qS
hdRl8IBGFcMWLYZ4OoOr+vuFY/iRk5SrpU2XlFHyToiVnh5s/BoZ3NbbMpJ5nIMq
TQ7e+bJsPxTZe4u2wO2gOAjf28V6ETA+4VCuEVC4K+Ll6Y9W0TfFltlfbFINT7nX
izTVn3UVILSYO37CMgSNQsYnIGU/jeph01kmIooRVhdxy35fbAmpM3qbEmMvQVyb
L7E+X1OmdMTtzqk7mGYbmn7KK6xBC11vWhL/cAdWXbW8SBCqdehKYsOMxH27Ewbb
XWQBxBv1G6ljpwWH7YQnF81FCDHdmp8phJBvGAFucSCTKFI1qnWc8fwRUAD6pf21
uQia7PgK76vUxWsu3veSaGTmzKKDF1wQRyzqbmOYoGWwrxVFeDNbirXcS+OsbZON
w9/9es/+bO1LlKwKFDIzRmTdJun02+Y/D1hIMWWtOayLH9G7DWGI281Tfzpa+BOS
idKSiGrepMuQv5KLXq66PH09Outtbbxo+e6Mg2x0qxNcW2CzrctrU3euylj0TL1w
TvR3zJ6DGC/mbpF70FwTnpgbdxl/QSncZZ1jtnqmalkXiSulqkrAUooDOvtmVEt5
6BNlb5UDHft7aJ2umJgluI8EsI0l27BH4Y2z0e1UNkg=
`protect END_PROTECTED
