`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAjPXSkUZqAMEz2NrP19DRci+MEIIZPOXaIRyWf9XM/8S277yekOW0Wpuc3JTLze
vPfJX5Ody/WqYtcJCbT4LT2aQMWPC6uGAAbFtqwInuabS1dnWmIwsRPWGOPLRF4K
eL92Rl2WgW7QB+zkqqtGlL1T8gUQtIExo2QCmUD5AAI/Hrwb/Zm11IUKO1Hc926U
SXTnn35Peam2MyffPAF3gMPkoEViz8ewgAVcgOh1vwLpmPC/RIwETkkbphqlxuHU
z4m3O7yruav68G/dC7QbfB0UC4JM0FBilfJwInb71fLKzz3StGmgpABnqcYeTnF6
UlWigraP3isxTw6PQsDk86vYez8YvKdgVAcsJHgESH/FMCqHlne3UfqXwR8IVjzm
l/n2Z7E+1qoDSl2byBffRxe9hVjV7JCntnquFNQzR7gSOcCCthcySComlA+izGge
treWAjYIYkq22hcCDwTtLR3rpUnJ3GLICRWXdFOgTA4q77UMpXEBBD4cdvPYu/k4
wlhRGgjzQRHrblLT/iStM+10WWoHjsRWNgwT35wOPR53Fvq9QWNNhg/7704SF/1M
xGQCxisgTq3fgZPWELyUFEHYDQXAUMXbpNVBcbNXZCrcf5cK+VokZNT9FypGXsQF
966iAt/g2vHZ1mfXYxA9yul7QUK1XXtA+p9xF1+CeU8EsYZzs0LmtAzeBCNsMpTb
p4pDXVD+z5p0+Mq/cqlXCSOMzwQ062JfTXaJM4nf3pHpLbMFLa78E1wBIcYW1jSF
++InbllLZswWLnGJMuvW5rBsYNg2llTDwLUMsre66Bc5uaIXjNLml46Z1GFFYniv
LD2TC4PXMspOzQFuJpxC1/9KWYyQ3Me69naYDPN6TKiOor1WrJ7puKXu06dXu0Td
IMtPe5sa/FhWmCaABOzQ2pIoOsOs41kBTH8fFELpf2g=
`protect END_PROTECTED
