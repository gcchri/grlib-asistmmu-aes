`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bJv19ytmZEhTiuuGvoeIi9HUxvRm1u/LS6skD7jQDa6PALbAPx6V0aNTMpTevUMm
XQ3rmSX0ygNbvmFYOk4rfFDBHhfE7FZwjqwUXgh/Zin1UYaKVgpVsvgxUN8c7yuD
mwx5Yos/qKFH4dzhErPC08bImxBG5ibgbQxK3kElfaLPuK81v5theWtJhPn6FVZm
o05vMwSpqd8Epa5QVtUQxGSCKs8JMX/ltb7/mm/VrxmeibfmQ5xa3w8wN+Rfd5Bc
iQ4AAcfndXguZQjsZuhfNo34wqXzIcppX5EO9vO/AO42GjwXUr8cj6ctPMGkkjPy
j6Xxxo4dBNpNlNhNHRS09C5RDa2nSjOy28yMDL/QAGnuyqNs0wtHUTUw2yE9SAYO
`protect END_PROTECTED
