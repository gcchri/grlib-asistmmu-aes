`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tqr8084kpV5nlt6+0p6km6m9A2JSrjkqtYKV1yHgKeTZyYTFRzE5p1FvGuu2OQL
VDRcoeQg8PrjHwSPEQO+NUux0SYkkr8UJXXdWiYQoV1zXECYb4CWdxgCnFlXdraq
3iTyD1AvxGEk7F0Q11icWp05JQeXboFdQJKDvE0rq9RggvkdDXcrzp0yFWhl062q
UutTe7Rd2TKcGxW6n5cr1PGwWCFsM5hK5dVl/9O2dtLZQg+4s3ieoH8igvGr3mOy
5wEQ0kDXBc7Yu+C/0AoWZ8ye6Z5wRE2igTrkBXcwVOOPvUcP7LtVbbiAHYrSRUYa
os8/uwRde6NXZqmvVUbgrOugTASMw7fWBE6xPKJxkKlMVN3wPWpGsu0N1OB1nd7W
H+2JQrDT+8FiKAaWBE8zKq1Nv0iAZaUZIM88xGs6u+A=
`protect END_PROTECTED
