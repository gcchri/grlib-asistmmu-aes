`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yrrcdLN4AoJ8TJbCl0fQOz6bl5iG7EtKssCs0/68dZRsij2UfwH1MZuNa/HXfEWU
O4zx66aDcOapVCpIai3wg+kGGC46yKUhE4kUuv5GoF+Ls41EEqfkdG39rrgsbLXE
MnjC4Qz/zF74Tz8xrp+cZm1WxyFPFAjqqDI6k0VB3E258wnutwmHis5Ts3SKmgc2
NNHb8sAWRi/XHlP1/+ZPN4kB9T1UACCOZqiZUvFzIFwidNbvYPqYJ+2vlmsB73tU
s6/T7tmDqUfQ53FQ1bXK5yJ7auHXibE2XwofvMT4iKCCUyhOh9izHXzru9Zuzc9u
JTiB2bi2kWy5cN3LmhYOix0cTDfenk9FM9FIO6ogAWXvr5RTqJXl3pPzkeAvrAnK
6jK79WG37Wfb77EXWLg/tcDJx0hvLbtUvs94c7zBuAt73NADzlr9p2S+KVWl2ZYg
kdd0n/4NV2Bl09eM12OXY9gDRbxhUUjhBg3EHZKw4tiVwculGa4HbHaseYc4657j
ceq/EAs1zd3SToYvJ4GtvnxC64LPFQw3lfI0Lae2f9JuBNZmE+30+2/MgFDcMuFD
7ey1qe3SU2lZW1/AE8V1r05UvgqfkOmoOlQIhF2o71OI0fqOdKGAucwkvvyALGnH
dNh91vV7h3b1Gi+Fd/JkWSXJpiqQ6FN1E4Fu5kS9DeZ3pzXpuw/F2Do4mU0xaSJE
`protect END_PROTECTED
