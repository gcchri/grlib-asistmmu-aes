`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k1W8K4ZMeycihyzi7fXy1pymfC0jIPzfe52/QbMTMNZ6hF3m4q6TzJCB/svxjgZY
zWFDynJjdl0m0obPTJPhE0Ohetsdep1vJAH1tlK+VZ+Ufs+dKAGaN6JAkRGrf88H
0nCRu+Eehgft4fltRJaPK0jSmEAKSfXkNAZP/3J2LpNlKMMA6OV2SW6vOYfSFsDQ
/kg77OUEUfm6ioHJol7pQnATWF+e9RGR6VQdcCovnT5Po/krd2xqcytW+XaK34YA
nNXF+bmaBRJeHgnBSGacuA==
`protect END_PROTECTED
