`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+i3pG7AZOxkLQsPn86s9QNF61Ru+lZORpM7TLiwfrWrfimSO+Lgecp0Ezxd4HUR
52F+eDh4HwewieEfIdk9yYFlEBjUFq534Ey5mm0CITcNCgR/WpYTtZz2VIbH5SWc
13nLbmMvv7ChW0mvbGiQFXs+Ax7Jho5ZTrUTbXLSjDThYMKw5PDGbw/SOBj1GGZC
aEnwfS2j1nfy+KJ5Xj8G+ql1Of91c4gX9CC2i0q934aEDZzckLaN8vV9fzeMuuak
J06R1bl/uniXwyhuJdki/1EnRnBDkNAyefmSqLyEn47jN+CvDXkDql0Gnmisq2jD
P+9k5AjwVO2C9/zPArqvp2OTthJ0kKnYo26dv6rm+eemtt3xNd4+CCoc0gSLz1SS
0yP95wqdVnFYrTvCX1w+USsTRrz3xILDCIGqAu/OuNyFXoY0pDhfYHO9TCGGIPg+
QK5qm1fvNsZFlsZG0aHDdtts2DUyBBJAHGYQzzN2WLvaWc/bmGvHGY3kEM0eFU7a
KnQFqaFGW4gIUq410EQyi8Zpk8lgy104B3jdwo0N1ooIpuWNOjxD0RYaRTfokJuK
P+JQHNzQGPv2iFE1kQTHihD+wEeY1JJUnCl+1KyQDqMafs1M6Made5U4eN/UM6Qr
dRw4W1w9dGLC8ih6H5Yw7Wv8wLFJ0AZxxAQeMNBn7BzrYLTSaliw7C67EdI0fKz1
OPXxlrzYmpv7VPYyFovQoFXoRBzgPbA6OZVOp44orLHpMukvGNgEBDsrtZRrYJbN
CYDtMI5WIi36yb5GmUdU5rXR2v1mB4ZtAX+qC3KXvIIIO5Rm9B8oIp6ep1kxrgcA
JRKb1OL3pZ7skfnC1aK5uTFCjD6ia8YllCJBT5Ur6AynZWUI4gcMxfk9md1dAQGv
sBiD8N0j27i9dzJ3mqZnu/r3TBepiOZo6lZsXVpHLaTVQLmRuvPK9dQAcjQD2n6e
iL7USj22EVia0Ag7hy4/PPJn1nA1a4WCy6yjzI7wn1nKl1hAOZaGriws0W0ts2Um
MeupS7FEwR1v7FJ1JyySN2bu3PEy0bWsTmGMngdJwIhwX/S+hGztM+b3V0KhM3Ia
HvY/BNNKnB/zmZhIKpPAHSh196IYcVnGTmzp96U47S0m64XYIl+9kPjulDKZQxig
f74kkQJYOhIV9S4DEQ2F5iMgI7YQLY32yyzX3pH3klDi9wDPRKb8hI9jBw+sooe5
FlNQvsqpjEi+rTcoVDGZWB5KWI79ZeTYBVt8ZjNHBVvmQ+eW/K7FumXQE17dhCOL
zsKVV129od64BIDabFNAMjD8VU6CwW6ngXqeqvKZmjuGhYquDkQnyvDhsKn4I3CA
MMVrGRt4OnIfU7j7eVM8yq9eeCXL4vNub6SrcIGSuoy+Y9vzWM7jf6EJPhQH4OHW
WN9Gu96FZ1veSHj8MmXKO0wOeYeuDWU1HPQzN9tmvuQ=
`protect END_PROTECTED
