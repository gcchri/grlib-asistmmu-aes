`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
trguhGYdfgksVZihohp+GXQShghBJkTyAnP3W9qVAeocXDEazmIt3X9MXAsKNjPH
M0nzgPQ50C/LO9mObwv5kzNKe4AKVK8FTGYlCXfa5AAMVyGgjA/T6ud+LI4WKIeB
y+ZJUFvlSpow55r/bt1pNpL8H4/x+AKIFm4iLPqUkyaptPiI7cLxt2hP238aOVv0
tQCtFvp3Hy7e+AZXivi5c+/QUN8vk/s0SsVR9gTYSV0NsCJdHyQLNa5f3DboMKOm
juWV+4XJeLlfcz3o1PL89Y3PFo9jYxZKPtVgIyQEFxhADe59CBBxVJFDPHK7rSFb
MIz6X2iDj9cwXlt9ebNMx6lJwFUrtIQqyxDIznywn89lDKkX7tvJf2GTuBHKDbV+
OULbFqC0hP+ZCCB7RQguLY3KwYjxbYDeCiKeLtH6YPaBFzsrVQR71bYXKHVDFD/I
LnnMvxxIE+ZejpBHi+Yqfu7VehPvRCLlT6jV6OmA74Wjo3l4QDtlEt2X2eRpj5OG
sKXvN8lUPzCYoQQUq7uLYIHrYODKI84MmeFBKlYUu/sCGTXNw323CJZ9iXQa1Cyd
PBZRvBOUZirFcWr0Vn7NoXfXDJBM1tx87TEIqcKOH/QoHR2zoofVykPpco8ktgfq
AFoBqaUHwJ9537op3Fvp2rGEunhmzL4VR0KSZOgoBjU=
`protect END_PROTECTED
