`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJQz+HXJH2vBNXFuobGoE2joghsvm82MWQFg0E2oIX3DS6SBxG5TPqMk4TuqBH+L
5GkwgMdqBxm+K6yVs3Jvt+Hn5R1AclJaQSRm+QVqR6qexuGzEbN0BlAmkeipoFRN
+ITfCui/FzxkcSmRH9J0NLR8fat5s3C4+N+K802oct76brq+9Z/GSPueafm5JkoX
worB499+Xw4Y+6HG6LFKIXZvByGSIn1CnMRxP2fhaSHcgrS72lay5yp1ea0B1tDl
10XM2YobQriNkCqnoctB2mZ+zdOa2igFkcEmf2EjrcKBMaun1jvmVyDHjoPBLaQl
pJ8xuMJdUqP+cx0T8nL4vypMzvzZ8LsCx4rO4KTPON+d3vrvty7Cf79dyKbc3AEZ
5on2gONyw1HFD5WIwkVyjGw+HPtSSqgWC4dVVnKS7XENymUue/a/MiXowDz7JTdW
WeiMp06WsdCQgwZNszMyC251eNcNXlyxNfCbslPD3fBOlWNoCptaApnpZudJPxFv
wvRUjAPprFpblY9piuN2S8TNlxWTvovMj3LelVjDJ52EBI7p+iQi5PQ1BFJivsFQ
9tSBIwrCRN8uprCNJym/4KYZDSaoAw1ButaFzfMHX04qCdmdPqM7WsdZZzy8Im/B
w8kzQkv5SNy9X0EJ2W57DR1lPcLXk9HVNOBgk2qT/aqF6HpWQ34De3/Ww3eiGE2/
iDnDQVJBSQjH/7trQyo1bArAcV5JymIINFOEsqqNZx6cZQnoXf6NbYfnDF18Ur+6
ATB8bUfNyl0do8lCLlDlIxRnQdNvSw5jwboRGD02GEiiiizc5au5OqvbGBfBbTD2
66lkxc//2dCAjaFgnACJdGOg9iJ3KWoqnUnr9mEM8xxgaHUstvDuccsMl7Swyhra
Bwzi1NWbsx6lk4rza50PIHVB5cjuQiCL2TgzMJRdx3fsKR0dM9tKsyNytXRNAPZ4
T/+Tf0QwUAmKnFVBBRwu79Cpql138xwXZI9II7+eO1SkYP+k6NgVMlYraWFsSJFb
ubfOyQ+qtrt7H7oCXoyKAF1XzwCU8bicr+oqIxELfRHPgFcdu9niivHtb+DdCE45
sZoHsrEaAvA6XoHGUMtqm77ZS0gNCtDVbNTGFgPEc6KuJdaUTlvMnqI9fXMYIsdj
jIiRHl6pPxCn0OrL5R9GiJ4e3Xw1KhLhBhvgnAWQu/UeL0OvRHCqSF3mYlxPkc+K
DBEu42q2nifJXr3Xcq8ItDBprt+8MvN4xeohL08IV8b7f8BhWKJ1sXDTZSjgoYlc
GdTkce//ZqSLZliqHbVRO3X4l92tQScznZqqhs6Q5GEEVdBBH+k2lhIGOF3Jgdkc
/p1f8L7vGNnYIDi/OAC4tcDja0gTPKAYAR/tjIgGpM9mhdnhAYHp5siZ5PAuO1I4
YBPZNjmqhM2kLLAtZMc6Dgc2crKRhULO84VQvBR+OLIbbXX6l1jxo7VyagxULFRg
F0oHhE/4ta6ZSAlTbHiN+OHsvyWsr4MFlfFEn12xkJcNTD8Hmf+fQLWn8G4Ro0bB
j3WXi67+48Qgjlcty8neuFwcTYgpN8Fkfhd/tXgoeVokmURFpz3IvoJnwgFRi/pN
F2lM7TujSlE5OVsVw9ANhKtRlkMDfJcVIT6I5JjPrs6pChqKlSIwAfeSss8iFQKn
dHqe/f4TaeIEABXTIZcM0wVl7+jFJBrBxKqiWe9kSOhS6obhYlmX0ljl/s6KG/7o
gBqznCbkwN14z5Yq1oGJMOZxoUvgxZtPR5KDHX4p6pg4GPRZdvrn7YRj8/YPn/Bf
BDmaz7VXqHSOKehIPdeparzTBKwI3+5e4JZAVIJ+IGBrbyci6cwE5+iaZobEmS/Q
HoMBrTDRQvFknWAwUCiM61JhN/tQagpUZCJAKV/jm74=
`protect END_PROTECTED
