`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wb6J54OUTCxNuCbEN2bZseGTEhSGtNT28Rw+ucHJ85oZGAIHcQjeDB8whRzJJdqY
kW4HUvb4fhqpCj7ULCgg1xe35rZE3RZ4BlWLVDstQ4ZkadN6UfXp1sCT8TthvUqq
Q0Ljy2+HnBJdPwdpHxMIHlkanqfVQt9PT3XCzvwlP2N4VoaT28h84F1+ZhDd8cp3
ZP9K6UlyYGg44xc6AT14NmL50IIU/YaIAHEFbQ4klIrjDstHuj7NCdKE1Q7DwH6W
FUhBAOxq8honog5G5F8oNwWutijRPQC78179ieNSXjHAuUUF7zJs1dYTErCsSUe4
Eif9KdBnsilxjmZfCHcJ3U70sznBODCJNxew/NIocjSoo2reTTnG1Sa3EewjaGBx
O//Rn09Dxd0LlQ2DyssFsAGKZUQFc+FmGtateVqzlyeECUPMT9aHGELgDlHw5a6S
Jew8OEnMH4QRKqHk2lYH8qBua1QBWRBUmLJS3nFBwjLzXnYgDjFy+g5/Ui+u+t1h
A859j4PA9l9UOAwVqYl9Ts4aSRs0T4IGOsBGwXUTLV5c1LzSQwFPJ9SECa/0HCAr
KOeW8wJuDnDoUzA0VyQpMQ5aJyFmU2BpQZWgpxxRXgdD50rIPOoC/8puGTuZBZT5
MKnw03wJJ4Ef41ED7Yfq74qDVaSIN4+PwWKZT9vuvwtVeu1AH+7Cfde4hMXC6EV0
P2lt19sj2QYsnso94CNcljV2PkHgbKMYvguLOWAe/0/ZgZmUCXExw3MdtZQ86G/S
YbsNTL+kFQ0D2l+rdBZSkA==
`protect END_PROTECTED
