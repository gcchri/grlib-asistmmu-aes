`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eveBg/OMqcUJmaEyPhDDfbcntex7kGjiztrYWbsVFfftjn127yuYaOINrSCg8q3N
hbENoF9Wga3CEZsHX9YkD6L2HXnmSp4qEJIy/j2dvHo+kkD44VYEP5Rcq6NGAFGD
fvpYg6dzHm4P+QC2xdPqm8k9HtbNw6fGyxyrF4hWVVJyoUV7JwY2SuDwRqYyHqj3
nb4GJBQnpP0fHxhppyH5XXhfqNU6S1bLr7E1P3CYX6dBRuMUuZugay4K47+w9qx/
uU0aSovC6po+TiTmfwFH23lDzwQ5QXOgEv1FaJHf8jVJcSV28kRtqEzVHDZzKHnr
J4K5EMvpkZmNB1sl7th7QnWt6EaXAPb5BQbRoEN9M4tgCSHJkU1c1n7vu8PYd/Hc
OdtRa+rIEsXa/3jQKl6RQg==
`protect END_PROTECTED
