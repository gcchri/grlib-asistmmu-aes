`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Db8/Qd6X02I9j7doyBxVNJvLvwItw3zk8XcX6qp+TDpytWE/9SMNpl8lMtPp1Rto
ucdjzFitAyOV4xrIdn+ne0fyYsb88q85dsXpXC1Q9x1rzkWPCDyJvfeHmeXPjw8P
fog6pE2uATv/SDAWZiWuHtb5tKoZmUdnYR2AnQInpfW7SUEX2Q/jIWS6FO4U2H7I
oQHFEzW7KRQ7m6gGFLfXFuo/tKXtboXbvcMRMZIuUUeubZjxOhFIoQ9rb8NtN2MM
2WbPgOG5BMuxwfRDhFgzRg==
`protect END_PROTECTED
