`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qELo3k480uLQo1oDy7g8TzwNs6ksJpaor4ks/gh+YThjFGPM1PuIDr9fapr+mit
RFjvc6IBUdVVpCfMHItSCGHzgKVpQXLlErf9i57g+MT6T+BCVLPo9VbFNZenERDK
CZR/2WL2m6W/axL7QI17bJIfiJUsMsmpAHet26ZaplAthQ7WIAp4kOowbplK+Bgq
tM9xNY74MsplngybcfZZpgH+pnlOJ/OQFujDceUl4L5Lop32FKTYUeTWvyV6fvZQ
wWQ3ZEYLKmniDJ8czmdCMJkIBVoW6kaLR3BG/b6C+4uULaDCmJnzQDs7SoIJtPdC
PET4PnPfq9f1Zr6uBLOqWWNa5a4DjpStUm3G/V38ZcCZiTVElVB2TBQTPIXtB206
ltEcCBaipWI8MFcUYQXwT+Hepn0VAnKMUAUsYKz7XRWqsmN65CLz1vuucBUszH5+
uKwAEoawnMzJzvNZLMuHXWTBdTp89OtbhYz01CXZ7VUyijRHM2P873OHopk+aycF
CfwDp0pOv1VT2hPO6s6GTAUqXnLNNc2LBzZfisOECtDdvc/Z3mpcB15n72Wn7biK
9N05bhiD219++CqtKaLIqnbLqp8SPE4q4PhtVjDyrzpglBhMd8WXFv1QlC+B4MYI
SuT4PQNc6xy2AVj4A0guuLce5BslObkj04QVC+nV6vQsS0RqiIKb3lVfxWmsKKbc
jgYvZi80I71TlrTrPkUPzp+psPLiCTlu0fVux5nezovo092ziNuZQvDSTlKhuEsi
j+tANMvwFSHqQCq0KTLHljF9N2+aqOIVuBMhptBu1IrWn0ISH13Ymf6Z2u+kdtn/
zow8ZbpakdaUtpMSMP/NzUY8+5/a1nO4IiVya8tWO9TWB7kUEhxyzmk1lnjPv28h
xvGkHdUsiW/6aepJ93SJGXk5j7Zt6embWS8aFWIX6ZWFQOepBuh5tS4QyYDYMVcO
z4hxMvHIJHTaJOQAdN7yijnlBvJIwW/AY0px0+jyUAnnD8nFOoMGVoqw+NFD63gF
PGaNrdL4TSp7DcbCoINIZOEquLbEfor799yT8g5t8moyTmsnpzv+Xqq1fvnKDqKF
klEH0cxZQAxSPwZrsiLydWVxLJYdnzjUWe7UVsOVIzk+3fsw44S87a4SMLuuQMSA
a5x2J9alNgSYMzmUe6hJbHXJxJSTPUQuOBLuedwUYgfUcp1/83E3FBwHAyBlPVvE
WPBqdgTs6c9E5T1VrLn71QzV5vBly7r9TqUuSIsnzximKPfFsERV7jmHxoyn0fUS
HDNHjJw3ael2bRnLg8OrcGqj698q+LrrGmHBnbZDq4yNH3bpgn9iaUgL+xG4Tw4x
NSnbZpp/QTcNus/FLEFkXRPnXMDgvHQ4Q/UWeAf7WNAyOvAVCh15lo13e2c3FjOf
8d4PyhtRGH1utUprM7ovndfX45vEfQqhdoeMVNAcwXZ7BabLQLgpjt0DN7NufSyE
puhYU6NGOnqp7b96TG7MjTl+YGtLlO5iTXddtVxkB70GW1Zp+TO6E9IK2E5U5ENt
Q418GxN4UdoSJ2A1oOx2ttGskCwfGunHmCSYUyW4Y66cv0nRMWd31xhuNogl/SbY
SHuddH6FlCDsUiATxAokTo/W4U7qoyeV4xynweTjds4GZddxb3FZDRZzLKS7Bt6P
qbKyx2U1y/1A1MjvpzPuLbDOXezy3lg8AwMPeZZlsj/jg6k3QO1Ca+tFqPmjUJ5u
i4cUZKHqVuafUOYrVRYKFPAJIT1+Kr9XqCP8Kk8u9uevo45AgAkGBo23CG0l3rDO
KiUCdMCi1qwq2f+DsRRZjU+/irIriz3S/ubCi5om2kMQsPI03eV4u4cPr/jzCVl2
1AzR3GIa+ii4OQGXLT8PGItS7KpLZOTc1utJ52Tu5X18cpmlULWErqH3UWExGGCI
TLQ9Iun7MkKji40wRiZuzCQrvI33kpcRkaQAEGbYFXfP304ANogdwCzF5N8OV3wS
Y2HzpB3goGWecV8j0CDC2aDNRfNfw//C1dPqg4I94FnuIs6saxXVblkpgB4NTiHQ
tHcSZVZ9k1xX08OXpDrEQFanM7FYnx1Drq98WL3VuuaZnao3wk0j8t87Rl3fLL/4
saDHAK9AszCRQLoVtvCZIE2CFRFElu1z80ZdepfWkUWeYjgT9iN7VbRr+DalIWfk
J1107rNRQH0CqBRdM23wj52XnyuWevxGVafyUxB6aJOTxP44wHRx9Tzzo4vC/2yK
fAZrxT+LQBiw0oevtUZCNYQG/SxshvzeLTi+eQJj/+u5QDyOQbbKoWOs5Cl5UEwB
3fPbWqmnDpVMArRRYy1IKJ26ACFnqb458xKNzctYGFwJ+/SxpVIn7EIk3tfzgs1i
dEXVtCpxWWLdJHonl7ILmo5P0f8J3ibUUqTRUX6LX2MHvneAawMcvJwOu1RL+Lbw
xSninj8gmzSRkFq405VmRSSfYO3ej4g78aKay4Kwq6fR+2wdlRe+POFhmo9p+VHt
Tt6mtrzTijyiE5tbsUYME8BTt7bVm+Q/SkP5Ef3c0eKrKFF/kx/0r8wwEald0Ic+
/EpN5qAWvEI7Wbw7Ni5XKYemdb3AcF6AMzhI0ChQpn9VMQXPYJTfxN7OaivGIKgK
ALOEqmnpWmPBfOQt/eF//6KcV02Rh0D/T8SZbL09Ssszcj7/nspDEiSDSwKqLSZs
pfE7dAoDnkscVD1US2PCk3NVb2Wq/RX38iqs5S5VIYT8BeNfrdaUMX7uwtch7xv6
WK40R79p6mtq1aTdsTG2DlnTZ9tNIo6/OLzaR5eM6xPUf2SeDt++No0xGJJp8gIa
mgtnoYLsGL0+AkibTpvCK+RtXu9H+zsF3r6nVdfFpwQYHmvPrVkSaVgzjRNZGHkl
lvVp5rvTmoifctNuJYEqOX9lAR8qWXnGUNANHk9CIIETZ5in2GHXWeZXy7+1CAzT
GdgFy90OZopjXDkJeWj7EZJrPS9EqkdXOzPimkezq1SZLnnOqSEgLHzrpwNgEEBW
1lq/6zLTrEkxNLDkeonRNS7HmGfpkhPE4vDmqFDah9ORfKkn0JT8kfJmhajyapDr
5C02nP53xf+2JOWNaj2hXulBjKwzGoFEB0YBBYu+dYOtUO5EzGW/s/Pzn84kWvXA
DvZqsbrYD6Y+thI0AOc7Sga7uOnaFPHkXvmi1EJcg5IsNUpzGRSiFJP/696xNxxe
B3Wv9zcpVTsBNAMNUFDgP5/YipY5yR7+WmkqeaaCKY7VcxU70aAwATcHZKnv8esT
Y5JCQaPqhMzAjvHhyEahUS0Dk1B0etoPXd0ULwGbuVDrLTNEo84rCatQsIqOhTqQ
HNmw6A8U8wiisYLVauFG50NEQkcQ+cx2BFwKz8+hZpAwoKAEgMf1kvHgiCxEjIHw
dApJoutWVKSts1FcdjctVP+K9z6bdmkR8SWESmLURvEnZoyvmIWSz+sJP0AYUdEE
Tn7dB6mUPWWyDHvX6EVuUfaOGV+smFnVfyXxLNt9WsT2Jvgghvn7LlPpsAin/yp/
O3mISZLjrua4soz+TJ7Xejva0uoqNxiOqI6IyOyiMa3D5gDIFY0eEN+4AcFF++l0
G4jDVV5HpiKIg6AGgkeVqGa5/xwDPmrNw0hrzaU2V43+uR+biOBnpFolbZfQCf62
6RoRtfvkgFiB2MkaRMn2scJ7JKN1jXsFxE5XQDIB2doKLkF7R0lxvp0eqKlWCtsS
t+Ph8ZbAPnx298fj/rq29RcOnM7figMOWrJ6AzT3YkI7x1MNuYDkKuKCIdp3KoqS
fFcTl/49kQ6BaOvX56/DcyT3abFfzwv79/jjYWyeTni8aupBDuX+SyRTIZpiO9n0
n6XA7pkgtbWOJjfjygDA5Iv4D+NiOZ1PqDKxQ9JB36y5ac1E6YnqE4vA63VoLABm
RxW2U7pRHmAND14GGBZYbnczWA9z/NFfYj2RTFEiW9BKe5d/nEil3rDIQzRIt3hd
IJqsvRNBS8UYmi9/8LMwhoCdHYjIsCYh8EBlQkK4AzDedAe13GF0QQWgRY9NsS0f
tGUrjD8ca+MiScjGYNGeFlcwVIBIGGaZSBWhZpQPkbcaJP1zYR6uNetiv5Ke9CZW
SN2T2Ud7JfF+5TWf1NyIhxBeZb3ruSBE4OPvIAbyAHcWhuOIpG2spQkXeTZ7gZcD
F+E2ZiZOLpTC3gB7bSUQAhFTKWKGp+xL3zVnNpqpbFRr65hs2H6btO+3qdbcREA0
jalUzn7cjO+tvZFwqWVL2xYg92DPn/PpFhoe1rtkozn5kRRyHYqe+Z3TwNRW1sof
EVBlCV30CmJbvGH+qFUPxiAzttI4+PJZa8VaFCu1LA8l9jR9wt/OW7Y4nIk42QgT
7XSmuxrTKtyuX81LX6Kxz6xsPW+uVrTDHVEgq4/A8ABGqL5ST/yQhf76fvSUFSuJ
KdYHrITOjP0gUdMUgqg2A8MJ/7kn10IjnmupuebxHbPB84xcp/HtZ2HV9JVvdw5A
dRYJCEL+tCtcIYFS07yyjtB2hWCRFNuqsagNtc5mkzBNRHV/1cG3+UAO7c7wXoVT
099ulfwS2cgqE3leva1vEoZhDKtTTq+t/F1Wp/3zyNx0YtSh83vYfnM7v7g0naz4
xMF5E1kPn2jETUbgz/Nd3vx/q8yM0vgkcFSFpu3ZlK70IMQ4WLjLN9WZeTvCZbe9
pNz9MOPGPrz9Xas87UGpaGc/ddLrTm7xM90Tui89BmJ8XB9q8RixggOC31q0uRTm
e3QD2Y36zK/Px6MJcfAf1OY64eCjQXEZFEntv4C42NZgpD11Lt0TRYBi2rPnPH8B
tnuqUQvKQcqOiSjvaBvnUfmkK0FAQF3h2hYd7xFWONuAUmQxa/IuqZA0ppuriU8U
dE1bu7I68RraaDDYopVBUIGKI57feUzKlYyUp/1LupnKa96YQn1whVkorE8NzgBd
TUkwq9XJkpLbWfKOqvP1LhyI5kuVyx83o0YqsnUM89K56c0XzzCUKx1a+AGursor
GlWGsxt1exIbvPPCi4aHGbx4t7Gs1zK5QfAlvM9FK4c5o6PbwtWGgJrnIb9iYNXF
GYFZZ4tlOzS5HU3b+cCzI0nPvxs9jEtoQdzz/vQX4StTQztCUvQQWIIbokWxGlBi
exTrkmu7XaohCvwRHDLPCg6aKarZfU+n8mxvPHdRBw1Uh82r5xGoGLhy+YpwnpM9
ErXcoO7lc+gnhezkSpJnHqqCh4rALvCVcxCDAJowDJgW+8kCjFB2H5DrVE1flqjW
UWNOS7zeGTA3EhZBhFvxC1C2HJsN7E/2DPFRcemJFEqrAP1klAERHC9/X98JTG4U
8nnlBOWFkeEy2s7dW6bdIA1s001QXa9YtDt6a5NMB9Yi1aaQgD0YBeQvSO9qLtLV
mS1bhq8lnjwDAAS73UCsZE4bpwC+EmliUNWzRtz57IGMUv+JjuUQpxnaKharilrQ
nP6c5f6YlyAudUxGhUw9ae8d2KQe11EZDM2XAojFhZke+1rXvKBFHRhnabzMRy+j
wdZXgHikuWj9h1VMQXs0MOxzTmqsPvTkj8Xyb5WpGBCaC3+pvt6lSh1x7bTVVzM0
aS+WbnAUk/W/rajATonOlfCG96E9dV8E31SeDqNhY6GB2KJOtqTIT9jsUkND+mBO
UMc1fpEdgvG7VTiw+wa38tkIcZdHQky7rEbQ6yhmvDNOy9FUoWaqEJELe77MoYRB
tUP8OviAhtxCqdLdNnxyMWrJwQ3ZPxNe3JVBcSoaJwdjdZiXNUR8AMwf8/eE7Pa3
RnRU9FiTmRv5a20aKQPaa/ipSSjOnnea3WzFmLVqoIi2MfOR0kocmdwN/tvGljhq
X/ibkIidZRFljKTNPgxGeX3S7aAxZqsLRO+D1rOhzXV20XPSm6bKamyhM80y+Owi
nio2E+Y+a45ghE9iQLwVuIjEnmfnyj6PtqrjX/2IXQBG40jiz1iPQdC+7Oux0A7R
7S+WirhwfVXXkEIo3Yumc1m7CXOq1KWHIbfRkM/qgCwzWk6ksxiUhRwW65z2HPVJ
HJ7CXOMSf2vlFFoIeNOCqvYfIwLwixORnkyuK6ysatkZP/S6A6gejN1eo4enfoFQ
9vmffEtTdwTChHDjjeJs117v2xEutZtQ6lwKUHKMUVIl+FMTf5RjqHLIJsB3516z
rsP5ikzbiq8ezVdCQjoYJyfSdkjYRnUWShQ9ccuDpHxbtG56t2xKtl6zTemXZqSa
MH40nPWRur8zWJVmmoq7S12py5sIUCZIcX1iMlzCLMUUYoIQqqKDhb1PNW74LKCH
RAc3qzsWtIUA1RL5n/8RY563EpnC6ijyooesimWOBDcNTLMSzLQ/fUHYwSdKkfOg
BiEadMjssCA2KgaOuiCngKZynoSPYU451MiNA8nh+18uz549Iyzt/smZakmU+a7H
GqCeVFgxPj9lNlDgSxnN+vAjGU52avcnDlevcSXtjZfjh+bX6X3pHCBdZ2DUjA0e
rTRHX6DoUKr7+eFVJOG81haQH6hRBanhh1QjG4C9q6qYPHEKcsVUYK7X+2NJ6Nj7
DVILC0vbzM/jw+s0vgebzuvHaFjwPPAN9ozYI7rKLQT7OofbsdTy9KG2kN3O6C++
9orUIhL5uVXAJ6f1CtftDJXcHfRaTitj1wwmiU3guspOWNTDZkDxQkaD4aVFBGct
LnntBmp9OOQQsaoxFcMn+nAn0AV1NUuf1lEaKfzvGELYUbItNjbMsn71XofF0V2d
pzLRhawJkKLENwk/MBQXlJiZ4MsendKxnIc2RDTp0KETf3bCIjFJhaKL6adKVNT6
Q26bsf7XFBR6gxrOKQNvyTVi2VAd6lYtwLCITSu+CZmE0378PCmjOfNZOirWrGKk
xC91znrLUh6oJmBZXpeAT4Dp7PTmPiX9/iky35LfHjTQVEryJlzdureIpkh2ldjn
KSEgYLf4ZhZAV12cfgInqFn7NrZor0dQSNaWVkI4INPkLlqzU5WrLwb5QG8xdnuc
OuDAr/N2e8JpSLU0V4pWKFGqaFDVfvZ5OMp/2s9bGZ+9obr6FmiGF2H6KQoLJ90r
aszOy6Ndy0JnXgAvZd8s0pM2S3/0u3mKJptPD8I8q+7Ws/jF00TYDXzdbBrrAZet
a6jfqKDJ87JnYDmmE8KFVGD98aSddfntkOcDFduqXkz7O17853SB9xoZ2ar+miFc
SyKqbg1ag6qrO+96OeYBpO/GRT/NE4v9I9/orUkqLRmCNDIlpMVNGWYWXXlzn09b
s9owP0USH2SBLjLT97BjmFjk703anbxT2Ce/6RgbAw6uzJQRkpY/kVWGQ+0pi3bo
7g/JLa8Sv9Nf0YnJ2vl0rw4zBPwwJE1hXTmJfViRtvF9eZT1Gp0Cr6VIPEchKrx5
5D0Jie5eDpD8KMogLb7+5D4oGtlRZJ4hgARGJOvPKsQhyjg4KF6sHcxVUBQhO0RP
V8SYzwXNWl5I/mhZBoGvsYIHvjc4Iz4fiy9McWliwXjJYt15yjDgAFbFasW0ByWU
jx75eawr16+hZrUbG27iba2A2x4a8V2ip7j0nzM/gy2W27VmudUXrbD5wLmjw2Oa
SRAQV5BAjuAkp6Qu83iivkh0SJGAhR7Pku6oHjjRFZi30D5gszt6Uo8s0g4p07pq
3DapPdBMWuQLoK0SiLxds0rCF2UzwA9Y5EXqOzIrvxEEGrgYfH44/nn7mnBmNwrr
bjZlan/k9ip0puOtirpESDJYnvkJSRX4Nq4NSNsDZL8M9Utl9Gy5u6Qii44M6nf4
A7MqbxEiMwYF6giZj7qqbasFA8zsUZ1fyMcik4qVQG/5bFBX5FlKxtwIVTPWJvRN
Zl0VNfQd1sIGlO4iGX9/MuH4dJ1mXA4PHnJ9tUEdU++RmoIFIvAlSOBhWCrC/opF
MgpynQx2IRavxadQYIkwuT+4Vqcja751JQ7fNcvl1LIS9CNnb8mYWyOQz+Z+hoS+
JmK9KF+CWqNeIMVz6qgnpB65y4aztl/LsAhXQLUH40aosFIPpsWTQxHZdgIr+5cq
G15+NbcT+udWu/X3eT4tDJI/VceRqUKz6RiILg4qDYRaJncdYsJmS9u0nhczJlMi
QhMg64ICDB2SV7skNpJF5V78ioRzsRn4jHrGzpk91oBY4aiI+bHOAlRuqS+k/92Z
9TJqoV7SCB68W4z4DG6VkCXpDeAwUuvUDI6tWUYZBoUzDY498UCtMw036wUnTSCs
Buvd5aUWL0yZr7VX+WzjvIivKJZYjLdKtdGIfYceN/8VS9ylsdWBRfYc9G2yUtmI
9yckvJQQaZAbbOsoeEWzvlQbOmdIplEP3/L/ToMygdGyjndsDv5hXH+S9N/vYQI3
ncquFE0z6lXkcQsxkGdtCTUJid/ivR8yB6wd2WAf1EzlxlVF33lQbiiYQkveIgh4
+LRCTYRjwQaSvkXDcfKT75ElKIW6gZnByOZg8CcoQXa/9bUj2/fNV2jD6xderOeL
BPALH0Hq8aV1v89NJcHEkyjjFSftg2Lq6kXLQHWiqbAOMEGcZ+1AU4AJhSG3fQSx
RolJf9N8subhHyBEG65BZaI+HHk0baSQteubFbkHjVuK5vHPVixNRcfH53vIWcdA
Y1ANupVqM3OB7xemvE/htlWEUguDeFTaokttleeWhHddilx+rU5t3O5xaByad1nC
/V38yjas5D9pVX1JDYbPonQGmPVhGsS3iZEGJA9xicKOMJe7sDTQUNGq7zZF1Mu0
X0UsaEt65gBtWsIIiqDXjSEBxxl7TAkk+dbN14aJ24GbAgFos2C1LtebvZcq9F94
BXwanPGOu+Hgg9J1liAE71posE/PbqO0aPaH3uBFbia7xM/1ow0zAODNgor11t00
IQ6Sa7WX1477knYqd+itNhu2sGrlPf4ah7MeTA7Pe7UM8fZ7riHWINCHujqDccJX
LPSo7fc8ZQPpVlzFyoYx9Or00TilhLrnpiJ3HTSL1N/2PCqlnn5jXc6D4vlw4yuj
IMoxpRu9RVryjJu8vdGx+2r1nITkHBcseMs1TJFyDm51M35obNBzj3Q88wcqyMY1
Qa7owFesBjNbLKdM64djamrbbmavPcDz0VrmadRbY3YoU88N3tf9k6ChG6iglFYy
A0aq9wMDHhveCfW1EmxyeTuoXdbRDLqNhD1pnd5zAYxKzkLYoqlmtsVRkd5FWwO7
SNnuAhDQToOGm92dYrm0P/Ye0kuEo4mq3FuCUj1P4QLP+4n26uLBe7D//Imi56vy
1ZHwnphhsdDcoMS3pm2CjM5o0mioKFK7Hk9rYGLMP8LOpY8u1ZdgcYowBnfI43Zq
UPtW/AvC9aGG+qhqLa1DqLsJnUmnfy4tFJydtiDc3P/1vOLK3rdREqbVl7JTlSJQ
37FLBmhJjpPkMjgRnNl+6HJfE99GhrUAUUjiPV3KXGX2MocepS67PY44VcOvARnm
33ZdS8J+1rVkHdJ+enUrIpeeP3kuZAKC94oz4DG7roZ0JsdxQi83NW0Vrqw1oFDC
mrTufnrfCJp7y77eaD7aEiyWxOK9CbTpdS9+me1crjXTVqJh+JXnR1PmS5eHZJ4l
j6CHy3hDhuvS2S7pIEF3Brv8NGRw/rLxrxzevD2mUEzv5GdDgQL8q8ZXzLN6euGY
rbHtUT35qDXsF3SEVh0TkILnW2m8oe6UgKaRuJ72q8XEebhBZecVQB8tzH6hzpW1
RVwpITETko5xSR4hWssFerKFkKUFTEzsRAAkSFPfPZqRejU6Q+PQhWJZFmKyTUmX
gq0WumRDIcIM652UFPcoc89aOEZUDV5ciV4mhlf5o25GzflamFoUDqcp01R2ULMR
Id6gRY0cZruMdoSxGZxhho8DQKHc47GawLz9fvPC8WKS14tOKN2yFCBjYKG0qqf1
jXuY8mu4HJgjsUKzrFvO8sPOf191j9Bvf7LjA+cZ2Dwm7gaQsosndWtZLvuEliOc
DhCJOyGPO5BCkqiHAXAlq3JrgHeg7LBhHAsa3gjU8qVCmUNLRYOkijnxbk1QhNBQ
xZS/s1mODzDYNQeESuEVGo261dWNbaDk3nXMHtLfdaFazOMSeT5h9PfU843/5J5M
IxtArHkynzOsn/RgyBPnLWsHWPwBRM7IwLBCg2Spye7DfNJ/o8d1+0+8tRmU2Q2T
KLCGvBHvV9ktKLl9dHIm9ku82iSQW5dm4ZpMDLKwRny2mwdOUeChMSZY7zjMo0vz
TPBHvnOLFrIE8TfFbLZNxQpNxiqMX5Grb5CaCIivNNG9ZZ78hLiVTCg3BviPd33M
c5w80MPHlGZZ+stDIo07OICuh4kee9zqfemx2DwecuM+HSGYyFG8ROW6b4/Xas0e
vbPIw9v7yy7SchMku+uwReUFUqlt7aA8sNBw7TS0RJDVwwgrkK+Mg4pCcXnOpYCo
i6gx3e4HxuypcXXeWiJKV1cvB9eG/rkpIHHtHxRoVc7ounGZ93HFh6rFHNmyElsF
gZ7u0qY9lpGo5ncz11sKuX2JQ7Dkv9f5xJkBIb3VITj+kxxxDGWqljaLrT/sJYov
oOIUGi8JOcFsfRId2ki/l7KkCzwsaiuNd3XPvVjeeFx3K3iMniaiITEtOfCpAXPp
cttkwT291K1YhfYblcQhSZ+49zWMKIRQrYyOHvhp+0itzWPnmhWjBjiCy38Q0hJa
S410Pm9JHkG0z801hcay6+pzAybzA1Nk0ohgwHoBnkhUbkuGpqmg7QQW07pSvFBQ
BcZ1uPxA7EYvPWsBzciEbJIyOntPNIVdKVOPEFChifgdeCriMW+srss7NUMRG/1L
ibzlG1h2WEiPdJMcwEr4WVtP0CBt/seSKrmFKktQceXvoygANXcRymnBPMn7rbCh
VRkxPl+jRU5bVs2aZTB2z8TM/n02N6L0N1X8kh/HhyW9UuzWlNsKMRGR9b8ygKZu
nYdik+UMO3MRbr2rSl187asbf251vvQsplGkKgqwMm6btQkRfU6gGxP53sraoGXw
fZ1m9gCpT6EmaG3P6qYb37nPAMEj9a1JM8mY7SeT5YlzLLoCHWogDjdCdyLc3BkA
zC5QPOMSsHU8wzLBeyZmveBxOw9K3ujIVOrJXG3ANpdj/HLg2y3dtwbhhN68URWS
ybS9atjAkA3yhHrQomg/1tqDtOFPUE/jfghzEWV1b2t0rP657nhuXDr2UtiRQp17
cRfS+IfAb+HUOKHmxMhB8cieyzmhdV+GmNdTDSJm+Xs+KOY15boUjA7R9g28ofh5
RwC/lc5ZyqqR3qEUgrAw5RM9DXc//wQ6hTkLcP1LdP+ieZQhngX73q6fkOavR5Qr
zsadxH3BlZ0N8Gnt0w16WUIUBNVLma0v93uODQYd0MKf/06hLflhg3YDy6/erV+n
FzXtQgIO9u8+jmGJxQZZ/ubfiWTKh6byEWVOaUL6CGErnKzkS7n7paPWNsZFEYx0
jrU32BUHptioWBPLWiLUY7wlZ5wo0tbvj9gdLftzw4Pgbhd1M/hIR9BseKDMvEoe
/t6+aWDdlwD4Yh5oWWrEH5de8yObcqF+cTQ9kDLWbJRaT7eb2Rqxy38WdjGDQE2e
7LVYbW464tQaqW2D543LsrowFHvF4ruyuZAySVADbWYUsRhMFBrVVFK++yHYHT0q
Vn3dqvTfGUQ4Jzs960Hv/p/ZIC7MokkOaB7MZI/a8TRLOHqnpgbHiEZ7RhSkt+lj
HRAZaObL8c6VuJ5v1v6OXvNI+l/b4lFn/waLA5QQghYGW5BUfPKLVO8a31H0l73p
N0iNMIHZyLgyp3Z4ULp46nW3QTe22Kbc+LyuXC154KRMZ1H0HZyiUVGywKwhm9Mw
W07ySQzTNcrG+0FniNxOyDlY0GURqhQGm1t7ig1r90CK3ibhP7v6CvCNUD3b6lVf
l282OdoSUMKP45WfKWoI5V0tCV7EG1vgI8qNj8S1rupo9N7Ugwrj3socoZGPWIRc
gcCngd+/oic21m8MHzbEN4wxYQSyxmhf437quYLfrUFYLXPE/AWs/PPKdImceqCM
F+bEVq+LqVi7eib1R6/8g1gnqGCGaXI371DtSytXiNQ4a76iuRSnztXK2GVxnqX6
shDdIpFJyKU94MUomnvRRx0O/FujXb5AG/JV5ZJTos7HcJhgEjJzv1KJ6u5Zzq2T
nYApg5jbdCUZ9NjErLW+hR6A91buWdcztVXNAfXQhKWo86rtNUBFxW4C41WbJ93l
ZQSItL0rWXynmTzuzXkaWyeNnEZCW1Bh7vjbo7hRSz75DdFLlUC29/PRlsa4s8M6
1SMV4gMs8245DkSWBJ8+YUJo3W/sMz9Uu0PPzefPUV9YprM0qUYLdFfb9MhIrOyM
k+aoR1n8G19IJIiySO7WlfL+BCA4eXITUCQqupkR++cLDXBqf8bcU4LWGYOCT5Xe
w1o28JrhkS1DnDruE8dL1w0l9POmrsQq7r8p+Cg0zjdU/23kHh0oLyPWtfT/YSLP
17zY/ZM+Vre9/b+3n67OE0fqIGcrdlSCkLZHqlh9Vmxl7K+SibcZoXHXKLhl7PYf
8Ss/bQbViyxYl49oUGUJZdIITIigTMDCgdqGgAKRjy8hopssUsuPabbhlbqCq1j0
ty8KZ+vgqWkk22xmUC3giQNp4ypQLB0wRTnufNjbQSsCKgMvvQZs/+27iw5nHb1W
RXsUd7Zc92h/Sd4mYHWwtHtMfC9jiIKpiZBTnUAZzKWQkpvBsmhnKI9ab3kkph/P
mw3mCwNWLVnaAma9O0ZF3WiT4/2v5o9+gPJ0SvIUN2MFrVZ8Fa/MgU/1f6FZDYYR
pmFK+9tVhaKpenFZpHyk0FdCN5iM0ETXR0ouAinAWuw2PFYGRIwpzUQqqa1erM6y
VeCklBZWfc278HKhj9RwJzyQ4s+IVgpnte5HAP2AxJ6NPSbAeNuWYhCtOKyB9xM8
yPzATldHH41k5rWnQMhJHOWls8pMi5ecrb/yC0N0KFPWfpUkB5Nn1yTEyKQ7CtlK
KQvbWkhde7a2iE86eSpbbZr2gT/XDmL6BpR4GkSmsHYhF7eFv+2HSywOJ+eQm/Nl
OA34W+zVwJEPVl8ij+tfNoDtqzY8Tclrda3d4al95aTM6sk8/jftHFyqIUq4M/hZ
u1GIrMQSMEV4khHR0++oCDaJbTWWt44NeFhOVEpQq1RDwJsf31JrJka9YuZ5DCR/
VsLMGhJNbez1jNNHGAcDRxQe1z8NhNTd7YTVNfe0piKZmTBIZb79/KR4AuOZ6/V8
kQqxtqE1ZHnCznFRM+2E2LoM6XT0rwC93y0iS7UROj7i1dfCx8pZcafQdL+t4T1n
HZF/dHfdWyr7ym0jKRpkRDLYJIwRc2FgXxKUYJJsLE4maLHU4hInfspGi34Vv61h
c6OUYtqCwfGtfbwmF7wwV3A3vHZ8t9Wmpb1QzLG7jnjlkXTDoPzHlPQuyQlBGj6E
Hf6izaVxvE7aCVBZr/fiYtupYu0zPy1ouaDxCgLFzfofLABC1xVePPD3B6jxv3mR
4EHM+UDqxhL3viuoecTPNmWbVORD+QGA3ynR5jAYp+bh67KLL9+lGOF/lx3XcWMT
nOoWP9IjOjKuosCpN0tSt1qyXAYCjf0NBTLMQHFjSomW1KciVyzgDdEAk6EpygXJ
VL0UqZ0ta6e4J3QAuh1/hokXY+07ivLmAVBN0qIGMdnEEANZTKsSF1jboKc9yGb4
0fb7nsFNkvJmbkaKceZITiXKBzSkCLgD0nTKOACwnwwhUJzzgp0dQ3dx8tpjW19Z
M+/D6a80m3dPiQQ6Rd8Ui6pYvNuLGp08RU3nrbB0CRNXhmd64s5PN6+t3fs54FZK
og9JQLXYBVFG1z//RG9Vcn+Q9rNhoZYLJBujsIbpoP122YQjpmBshdRfzGUO8ymJ
vhZ2vsEH9zZBdyupwOY5rTqoI4H/zTxI0fNqwSYiKk6lASIVwsDJUSeHpaHXXQXq
cRINwKgh4nn3Amrwj8wCIFv3dnXjcAeCdKzKR8lT44gQZb7rucGju3Ny1aB4jIrx
VWQibNXHp9DnbfHS9Kn/mm6HUQm8R4QLuJrK+QNlUDZqiQjr4Y1Th5mmnKAn1DNx
noG/PKEmVI/GZLQuevH4j1kkYN87GxCQfjj3fc3y2SiAfSaHJg3oDaAZs1esMNLi
t03nKd1awsf/am98iqgyiJJPpnCaxIt7tk/hgaEoz1FC5W9HxBLqT+mf0WTsq4SR
hLeUdWmwQ2fUyJdY+hR5RpQ8ymh0IixAacDVFXumUfX9YgoGrVORbbgOg/oxQAwv
8slh2S+s/ny031EWNvtzUljXbdVMGc71FK7A0dIrA2s9224obsv7AUPch+oN9uXn
RNJN1l8VTgfCJwEdJOTX582UI0lDAN9snzSJCZfPYxcFMHfrBh9qiMkpUiMXc7bx
qbkM4PW/B8QYlyvQQMEOzjC0DPbeYursS7N8xT9nv680fHLrlPIY6JjlA2rJ32+o
av7DdfbJsk6Gcg2X7VYz/8sZuqG882a/MdZYVO7p/d7xH3Ly2cHKASZ3ND/gChJu
BhfcGrfPLkIMG1KlSbRKPQxvkTGXFvhEaBsvvUIcuQfRSRgb2grd1b3xbohqQfxp
W2MyAQDSmrmoNY/BlxBc+LMsXxgQBPZI7wbSxuVuY+idmbIwWqiJSS0gdPaVW6i8
suKNeVveoJAheD/3IKq6qdO+JLeE2F1xSH0OzmlJz2M5cbLR06tDk+FPA/6krZr1
jgqtF11vVFnXVZiCpViD4TqSa4xlBf4SUq1djVtmTYgEN2u2xkXUOyCtYSWKlUPL
+vWxet6zcJj2Y6qUECR1oVTkMOKKTzh9geTHlSHoP0cuz72SDPCUvUY13KWTHeb4
CTabtnnhlt5Nht8Pq2Rd8kIg4LUKTGqhSTB+GPDW0h086UFlK7pRiC8goOIeozK1
ovaTBw9t0yE+IcVdRL9Dh08mNqgAk27J4PVUNntsNQ6J6sImeCyTdZQwWR/g9V3E
kv+ceJXVTHw/5PJfksJNDSO3VUFfFzvQlBJBcFWapsWbahx156/aZRdPohthTRZT
LrzQdytaNS7n2XqX63eowSyAkNbVI1ATX1Hy3LDI3MIyvUMrZYTVlQVOSRyX+KD6
CbTJpYjRT62LWwz1U274GkZcoVMmz0NQC16UgqJdO0DVm/mgbx0/85abz8fkW0+N
lZSWxkeIb1ZvPFoDJEjRDiyq8DGTJGMtR+84BZgyCpQoMfa0CX2r+8aHOqFZDxZK
f6Sbw1DjJFuiUh1IiO2Hq6T931+Aa+//EUwZzpZaMuUDxt4FH6wYHvhaCEq3jrbT
f4dapHAQWk8I0XPrvLkqSCxLh0iF27vnkZCC7GnAO7jBgnNSHxLWH9OV/BS2Jp8h
fQXbVNQPJ0tK0Qg49QYzcO58ZG9/VkN8Er5vLCjuqIZoP7YBZi0ecCHYwWe+VPJE
rJxFqIXW55qzZT5RnS+XUiLLBd61rCNBLi6F3CuM6dlttUHyg1ey1WNdUTwOlOGZ
cbbL6+ih/RMFLR4KKlC/DQm5monraMEqJu0nvgVxStW7wSjq7aGol/3lQhbLnhOp
EqG1qNxp47qDt3s7eWYSipOEX6WHue7Ym0nnSx0HlVHo7+CxTniSivTjN0urk+/k
bjKVJEBIJLL5L4rA9uwCXQH8OnKNTTAicxsa7uU02B6gG5Xi6UhBDtAzdug3g+xM
bagI4i2r+CJ5Ac8VxM00F400bRjmOOmJPo4t9B02qDg3FbAK/bhVucv2E6tksMYi
p2JvbmrHtQy7xloRARmgAecNC1xPDT6iW+PJMTNo2UVYgQsGDaTZZboGHXKcylGz
JoUO+qdhHDc5hkVmAlPjAsdjr+/aT3UYTc8YpjkBwpSwKvkZv/71eE1V7O5ePLaV
b3GKYZjuV+z3bM8Qlc8kXy7UUfULWAroZB6ecmV6R7+eHPMm6mp8KsJD9/7padcX
z3v4a/tN337tJz/RHqYBqblDF+pjNV13E5d1uBL32IKgp2nULXf6KxBf3Ix7NrLc
C/NRrthAbFbBsBpdfztvfzmycw2/vpXIg5hvUbq9S0WEnfa3kUvBruACaUrQCKNr
LqQZ2XNpnlui+7ZyKY4SO/Aa2+7P2OrmQSYZF5o4MHD3r9o4xQHt30StSxOnZ77h
lWqsTgLiYAyI5YjENCa6rUaduDJZc6LJq8smTd7deouOkSKmiBsn/mIShtqNRSv/
W4zKhDanAvlcPnUMnPGbFgqcPSIiJ+hMbS41kOkLxj47crxeRu7PZ2+Tzr7+TQN3
+W6xu3OHo08lDpnYjdI88Z4CwfDElWPD7Jq5RqcfLYLhO+hYCEfiJBWoLoINtk/O
Su+GjqCXpI+wYE5yZtgnTaLs7Eto4jbTJbdopFYQ4wbAe6wfnBR6hkh+pKqB1qEc
tw0TNy6/BOavmgQjjUlb6kxSkdWQ6RtGsGzqMDEbCtMWN4okcl1iZvKHR+Fccq4v
+vZYaGC0ASLgH7Dn9L+KYQ==
`protect END_PROTECTED
