`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNFw9fPW6WhW32xts0gfRprT/B1WJhEs/Qdj4xjYkF95CcNETkipYvx9ApF7qu6I
S6vE0eSJ3z88S885p3ZJtRSbByv90DLVkevukv8NFe6cfTESdjZU0rq7CKX89b21
shPL19BtZWpeFNsM6EJMZEbSmDqg4sS/7u0UeJZESYK4xnOsajP27qIDnHPADSCs
G4a0SSpSZqT6xxhPnZ9Kp3ikiTTYTZSZYtH1PSbgDYOpOBhaq/BGmiozUSe2LX/A
3AiaC7RMynfsxJK54UWYMNsCLcURcEffe8m9x4H1gowBqdOGzI3v5o+vLXK7xF6G
GXTtdWZ+uvtSEcatNKX+c7JscYMFfu2QV4PGeLXdf6KGO106reidc1cJ3E0OyJtD
eLo9V8rFc3mcNe8dzi+Bmke+UPUP1kZB8NtEJQaG0rRFr9jBQ/HRCgfO0j1XLaGs
IsaSzKlf/vzNVHlZbxBZQIQneVvdKCEnGZwdw5tSOSk34Hgu7Izdi202xh3/EfFL
uC+oiLiV14GeFaLaFo8YS078RqYHsex2ctkHkXFQ+0SaqZBwfq9ucwFudGyGVvGh
zP6L8wKSGUFBdQq/7UFnpmGk8vT7zmHavcbWhDy/YFCgeHvJM8Z654Ir1FEnNvmb
OozHwXHG+0xYraqxGJzCWMeJxN6RCxYntbHXzric2PcLOhIGmeaSiw0VJv56zOhe
jkR20+5s+oPJkxHCXYOdLuqHTO/Gx/sx0Pdc/hpVERB3DIMeXQO7EbRNgk3WuZgX
nOiVUvGpCoMsYUnk2z8bKfvDo/eR2lpwfQwTb+1EGMA0qHLmta49igLLPr6zoMkB
EdPi+u4rsha1zCYSSJtHr/X/fLLZ4gh6m0EtLPFRl3J21bPbJxU6dmC6t3/guSxM
QqN8ZgUgk4ZegYzArzJjOf1kHmtY294KVCBSIf1eeN95/Y8MpR7q+HuolI7PSXgP
0TF9hp5npwZU3TMQicKTmW/yBDwUoI1zUkWDTBWQXIU=
`protect END_PROTECTED
