`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EysMZtlK+kmuv2aBw3bYPNLuAxVnyeL1Ifu+aSXfJCUwVt0rLfNtjKoac2niNq5f
j1UspLUJhCHwo6GiSeHvKRrsFP7Gf63HLRgxlsLUCoW4IDEYnyDMrd0w9CLgo428
MRbJSpDnzN6uJ/z7DSiabX5VYk1pqi/htMZvXUKPs/yuNFjPjFQ8xofoTtMONZ3b
2pExAYkb3u1RklkK7OX84VZtZCmVGW9sSogi3z8A3J20C89tLTuSFMZqqrF1MYpr
h5eMBcpkRmM4B1NPU/5prTxaKif5b8O6cO7dYoXMA1rNJuAAKt8sjCkbJOz7vGxK
pM69B2nhWGIZhH51M2zgWXe8Ca71R1RVDGWhhDHbzEkvFbaOMSLHnc2GPTyeaLwr
gkssIiOYV3N7NOLJ9WopRR3nNWirRDKtjH0DlVsYL3qrBaPk4rOWSgJBr6QDErRG
OekQlpFsGPw4/yk76SJbfzBrZSkLiOkXdfYc5U7ME5WdpcqrPeyBXiHuNZ23Jnrg
h9HpqkZorIArbSQymNmhxAJGwdwrssB8Ip8AdXVltNi5CyYBtLkHLOpsuV0aYAsf
M784fZrjXWXtc+iQu3aKZ3FQtRxL4T9MWp0SeJyW7Hrdrwz4uAMhT/DiG6DLw0lT
rqLXrS7diEDxhYHocIzBX5UK1p1i7H2KsO9//kzWYZOyeN6XFhPUVUtmp986QU+7
bitj9ncOy//DSkSxk5ic8gdIOxjmR7oAWrGg0jfPhKN/NUOjUmnT+qdiY+CdM6Fd
quB28ISaoM7ilTR0pPUjfTLzgQ96WiW9cAgioyr69akeYqD04g4MB3PXw0a+1F79
kaZxssSspvOc3leOfs46Tm6z+cAu7s2Ud8SWwuYkHcOZnNZRDsBIXGH9KqaWSSak
z7uga6MiyIgNaBv/KmXnjaAUT6oXQiYgGU3lsBEquX2lL6xG27+j4e/n2lBsW17W
vEGLx0AeQcDBDzTwQt1fgaFuo+qkocisrciqHSavtpUKCKfwODHSuV2OQxNwaMQb
Ir2E9S2rYbp6xRVVp/gjKWIUrbkEBvfNcTPa39uiTo5YrcN0a9unJpZcW9UCNbAt
h3kd/seWXBGrGT3I2cy3R28YR9RzQtKDZdJzF3HCY6I=
`protect END_PROTECTED
