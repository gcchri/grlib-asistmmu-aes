`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L00BJiA52HKaLryu3L51ZU6lrS7NFxF5qftV+u3YqeVu0KZaX+mVFDNquzSUcwmG
6opKK6GzEL+11jUg8ASvUxbWMbV0OKaIlXBtN2qQGk32zsS5XAFacTyntKHyda9+
Czz3RbTUrvavv8E4zcFqjCSrrkohzHo1pI9/ZxS4GyTD7mQeKVLqE2NFaYq0Ntwk
AvHVUrfLNi8+DRAlKRdhJ1PhDAjFFfTI2ULdiEaCXgcR5oSsqXUdELcGQeBPhRqC
ee8/eoWcT0+GKcz63oCw7V963zMR2aLasuV4QwuY864IpNNN3dfeHutJS9VFlBJZ
Y/cVUTuqK6bHsAzyLCpR9baVH62+rdYu58KnlGBO+Bwm30Zd+tmB0btT3uGxL8T0
ZlDmbRgirdEG2JNi1csRM66lVyw5QfFX6LgZme9XNnz1VNpMKJzcS38CdPb/moPq
ByYc9anMmBDw54h6ySFYtt1SRH3mAs6MI8B2fiL8ORU2mQCHz07CUCj9uJx+f6JV
6X/4MAduxBfZsfmAcsJu9K2Yjh+hh+Ac+r17PgdS7+4YLl0kxTckk/LSDhYzO3M4
tmPstGkZEQLCDICihRgKiMrRWEtNRJeengWseU/zcASyfDaCPvHMGSG9Ka6kxX48
`protect END_PROTECTED
