`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQr+vwtJ8zNJ3QUWjpXpAFTiE3TDlOZXS8xwkIUPnZYs0zJ3KCARNbWVP6O3kAzn
vki7/yaNEvNj6pr8OdsU7bL/K780Z98MaSSM5t9SF0eHMhoSDa5RKlyzK+rePX4V
necS3lJ7vPU8vVEQh6ctI84UnrtWMr+gofgJWwyFoWiJyE4FludEIOl0OE+UpiSp
QVECfpv4LLhmwbUTlsbuVN3V5KyiyXzQkkUG1EcItdZzS55bMRyP30mn/leapuoK
0s88yp0mXXCGDxiIC2VduO5Ueo02FN3uMapSkbdghk1qChsNSAFeaT7HzEsak3xq
oe7j9z9PoYBtLFIFVCpl0klckHjTGbY3vytsti3C+dfMlctZiWh/S4eYbbkqlHl/
srZ28ED47M5yf03nkkt+Jg==
`protect END_PROTECTED
