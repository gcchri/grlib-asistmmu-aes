`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94AXUajHz3yVELlmFZVXX8u2t/8iSYOYTLZgnioQ00O60fIdQi3YKMiOKvmiPSzW
JGig+I/aBGilQACoyuY03BzLesgpyejcY41x0aySMxGAR+u6xFfYKZiC++3CQJ3n
IoSo7fl5u/FKJ3GYPKYKukPkZdDAeOe/G/1G2PVaqj2gmpkf3vLTIZ6EnUdFMLin
qGOxuUl5KmU3HeMs9vppcaMSjKxS55fM2v1QtFEYDc9estDyRfKUrYNOTB61b0eR
GCSefTSsKkjmzK7hr7oaW0+kmNSfpinqTCpUZKH4XZ/yoCV7BUTpKpjuNiBkOmr0
o3MjK+I5Ooim0vevzeFz7UFoEmIRe3tMicy2XQqh2KZSIop7VjvmvmM1E+846Rmo
sBpESvC9uoHQ10WHBNCJtA8Dme5RvpHjILe2Y88dra0i/SMGXHctO6aqAt0VkRoH
CDuugfuo/8t1xVTvJMz3Mww0HhJsnAk1Q+7dnJtL0vd0RKOkiqyBrJOcuCNr7+VI
qepr1p+HfhAFEnJG5gOJCtAnPLjKhlHxB0Y+UYGHuOe/oBTyujkV0K38lMwQ1F/F
bg9maLiltrJSc+WEe+gZlMB9RsdzJXli93zAjPN1+1xoXYemaFMg1ss+HUH8LsIz
DcGs2EirdMU8S1wmh9OEDc6RVeJlIkGQ7PWO/xxSKYkVdI5aq/Hgdpm9ux5qtmMP
Xm/QPCvwC4eIWjOzAULIt1Ewkc36Glt+qXCvWsetV930MS0CkN0XC/4Oq9Cs4eQW
44N+RNSKFL3AQtIJ0iccHvS6+e3CUupjm856jM67CpO5PDKMUrEABlXoV1afZXmQ
TnC3VLo4GepDQyR8wZpFnToEngQCWu+104k1RbeB7QS1DacuLDtgCLFvz6mr4HAX
z5LkvKymEoUkzBK1xK2c50dzaGyrPG5yxFh1hSLKeiDDstIVikGCLmxvOMGufVeY
Lj2FJwjMATTZB7hxEhrdyNwrbH6FjP0y8eSJS6NYQkhjrOkw9e9JIWPYIiF5AMes
4RJniOJ7IJdUWHUtuL5XVH9IYrCktW4h36m4hh5B7e5QNJaxzII5FPJlI6khWKPX
EGTbuQhL+B9/KL4KcEeSDg==
`protect END_PROTECTED
