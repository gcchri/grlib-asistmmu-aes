`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PEsQeD1xwjaZGHnZc/4hdVzw4MliPPCFpHO5z3v/3Wv3/noTWM5qSrQYuXR993ex
6X6VGQEZdFlehbCPtLgAjA0g5geY/FKyHIcBzk6Qk37eBtAf+qG0XDwS0RHRnX0d
CAaHR3X+lZaybmNM+XUE9tX88vDhSdmk+a/F8YYgjPlXlTMEpJkrYDvzDA6q52QT
3NrNTu1BEh7tOt6CDmoqC4lVZSYdPqrHhxqDpxdsYHMkrVZN12ZZMOGneDcxhZxX
2OgeW9DWLMUrHhhZe7N072X7yo/gfLXwKuSytzSNgPUCCyH/W/MwztUEU0Jd/L72
6R6CbdRxzFh14LouXn0cJQ==
`protect END_PROTECTED
