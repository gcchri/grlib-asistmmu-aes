`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vuE6yKfKmtNnAjBlOPW3n2lopctDP/tyRyOurTL8i9CHxNfVu+BAsoisylfuSwdv
6lsjvVHhGC7PdyhP7EKWfGT/TYvHb0RxTq3PJTlnQbKFsEtxJW9Hx/j9OgLu421X
rXET4ze6qB33CBKzqKbJcCkBmeAcNwmekD6pPejtK2u2twBfphGlHDhm1A7/K1yV
GS/u5JlnIhklSc9jj60Wx61Mn2hjgY/hA42Trk02cy5XPKEGUKZgLOxWHTrUF/FB
cBN+TMAYmu+FvPa9dERZjb0HYy1uIeb2Toh2Rys1F85AHcSdArniAxkbywu110Vd
Mo79errorGkMgqT2W3K9dPBr2vuigR2yLnXq8xFzVBKqFkjtelc5QpNkGmjAU9i0
ll9Va/QZ35c/sgdZ+unAU3f/XdEmASenu6smpZ7kzY2O0ndTe5AZLbffVzR0eFrO
9CXZ79gYOrik1m7Gcrn5wropOMXbBNWTuH58HBH4098ahHQi0nHl2pLATrCVjJPp
`protect END_PROTECTED
