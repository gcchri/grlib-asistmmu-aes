`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJ0KrCRCStxtZ7YKuHpkLX7jN0jDyrF15ffbyK7iK+C1OH86uH4guVT8Ce2Qq/n/
7cfzLa51CJhrXgfk/MhQ9K1pomEzTV7ECLbIUeUjpaRtbocPDvrRVG5AXD3ir237
0YANIR7TwcDI1z3/NmElypXhwSJSQBIZMzA6x2KG705V4IGuE1pEzhvkw5YE1ov9
zVNEQumsmQLOpJ7ztpmf5+4FBJIBFfakrYbbFSMhvpsRRiGWNjMMopQicEoqPqVw
zM5qvM6p7LzXZiwr/Lr/30Bs5nuk56OO/klY2GavOBveuFl2l5E1OGIXdshxGmcz
nrPoykIzxkxrXmQ2LABdOQ==
`protect END_PROTECTED
