`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLeoO2jfY1ziGIthNUOW2FjTnDSy19XrdSZzL2ZuFZhobfrNPvyqOKbppAxyCRi9
0zR/QKLdTHJNrMyRji3ZoyRQ2DguCLA5zYNjZC2DT41K8rcjJqdhf0T+nQcZub2c
z3auemEuvKmV1jN0FbDVfhEL8avKbZg1wc+CpZCRKrWEuPf4Rq1+/2yNumVxNsrm
aQKuAFPs64cGLeFGqgYnvadYeH89ySP7zvLJ5hkq2/lzE4LnuSJRL160i1vfXbvf
6U/U8fx6HCbUejfWq6BRwJ/Dx1reCpr65Nmthb661Qf9JWg2xt2Wi7crnvzVA67N
`protect END_PROTECTED
