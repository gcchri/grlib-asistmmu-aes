`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xh3QV9Yu1KdSFzTcwXR1Fn2/pR63TRFZHV98gFbXpEuLTMKWZJ7xfmTqIctntFfH
SdbDw25e2XWYnRj3gIfZlReu02Bnsd4yGSUW/3sA8ACAcA1g9uLogpZl9E8SiYKv
wum1LJvXmO3PLdvw7BV67MMg/q7h7skWsR/kTaMy4gRMZ0sbaW+XqSqpDotAMyeJ
r8AU+4HzC64aRksp3I2SiTe5Qk33Qb1ASGJ0tZkoeaGZNt8GSEWjWoS139G0ZNQ/
fsnqkSLd3unvVEyctz60WgLRiTaYoe6vak+l0g6nSqQH8hG58n4RQL6BcV3NhnFS
K6ZYm1jRMM3jD4jp9EzHv+X7ojkmB25izt7DeQA1pf66s5xa6e/bbkmGwe2H87bB
x4Jl8D7FQ1iZjBdwKOmOdgn/ixTL8kmlwc0yw1RfHUf0V4TdUWwNl38uu5o/ev01
pZJ3qQb6uae+ULsw2lg5NrtEgzc7zfW9/RrazCq08TX3KeMr7dUERnZvH5MFnYaj
KuXYe4vA4qKdnhzxEjL2GogahXF9Kg9P+gbDAm/Nw/hqrGNmhdQ6mub39dg6fSdq
68eE4MXAE0jks+HfSngjAZtEBmPJrl1KbaeZWD6vlah7l6FUQ4WKZBGODBElcRzU
rt94GuuZcq6bjG/f4fOAS47YcgpksFW3U6Sp6+IWshoO+t/Sd15+7sy8YQTe+Gav
rDRfgb38cA6LQTgc4/ocrDQERTkLvnoqRVTk12E4JTocHgo6hC0ZAchqhHO/N7S6
mAx6fEeGcFVVgqMI3Hwb5sGLTK2EgWahmeYd1yyHMzx6YfX4FRh5vMW/3WWCOgCB
YthQZ75akbDnoOpxys+sxm6PStLWIfbig1Z7chFVjOliGQXNsJsvvM4Z9vAw+Lvs
v4mHUHBNKQ1mtkTHBbBfEdbafFDYLsMOKqCEswtOyQMTg78f4UcNNz8EMMtU5Vj9
+2t8pWf7MtWNr8MRcCEEPN5iRd30urJZGXCQFMXpBq5zQb8qYMKHfP/ARL15UjGg
k9l3Ac5OYM9igoM/dS4+3ArX7JQZkoOVRyqgmK8X6jBX9XoRYDNJW3HFlb0bPlFh
F8j4XTyatJ9fZsomu3dK/WZk3S7j6lxH2d6bo0lMme2rsJZ8kh3zCPuemUsBPS8M
jtBUfqdQiPNE6cprV7BXYECXJaPfqvHxOcGcehRDxPYxdSLJ9ENMR7fsEq/UNFE7
OTv6Ab8ZiiLb3Nw0frLqLA==
`protect END_PROTECTED
