`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3B0CnrcK8k1U1yo4o4HN6iewai7lIbpDmssCde2LZ6V2IjOi+cZuMNuDrVypbMJG
VigBf2RvzB4vTcr6qxQgg7GsQc37T8BZNBCRifbWB9wAaTZ89h0mvo9bIpwUXFP6
UIcO8qJzIFIIuSavs2mr8nDhbc4nGovXsyMLT9N5+CV8lN36JKid6lL1ZameqV6p
w2GNRUsGp8hevbYV2TC7UAINdQaGzcLeQIVS6KTS5gy0eJvoNp7+ROCQSJdeoa6f
rF0xiEhK+gxzcbqGkXAQgLJ98i1nT+M+iSuAwqxbxdan3WvsBwcBu1bnKWVF4S2d
N7ThZC1cXaxgQBmSRduqKOa0NwH6/yh6n2CcgVcBxWtwD8Xy2EvxrKZj0vbAxYdx
zdbTPUh6dxxcSrX3F6GMxg==
`protect END_PROTECTED
