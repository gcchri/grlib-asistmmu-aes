`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBU56dYCohiVWwLHRJAMK7z40bZiFKe63rLPq825gfcZ5H1hbRKIxjeQDy+Hq7Du
GtkkXpUnsEpajSOgRmSaLDtjv78Ue/6ArlEP5dNqMl51W/UKSHwbErfmWmVm5qKH
fu3qneFPXhPHzU768UzPngmbq4xH/GnQPmMjA91LKYaLvmktNEknM/H8dgYsqB3s
aBmzbGk1vlBrQbbv1mxf5BtaO7CjKKggqq75p3/6E1z4gog/EoI5vy9FjQD7/hUC
`protect END_PROTECTED
