`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hO1of/peeJG6TJf6KtHGdmBxLcqvtlgSlAtUxjG9CoSfgcd7cYyAxezxytN7ucHA
gLi4DMlEXxdYkBe8DC/5z9BpavI+cqqoCPPFL6qe/GB2gv6rHIBMhmNXhrhE9TDV
Sij2k1jgnlwkualb5cxTrlGxXguD+nvwcmWf1r1NFeidVTMaDgGQN7WKdneXqgQ4
AMEAFMX+katdyAhoXzd7lsEFooolAggb8s/SV6R0VX5PcP5NakIqj7bEsdVX+L5n
8P6ZU2iAyV37UUAGv4XITlmsgMmzleUFYVddbkjhv1O54mmlbaGhD7u4rxVpD5rC
z6/hJQ5toRpqHBuzD5+qtKVu4Al9Ob8C8JE1/o5pDqfYlgdkriD6SECreI40CAy/
H6xNue4PRF5FSP/xjGXs5w==
`protect END_PROTECTED
