`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NKEHvjkeQxNbadzuEdDquNR5OL5aJAAGzpeBiowMlhrGmbGvaPQI40B6wPsavQ7P
F6XQBdYpTxMozJJx+BnlmlbePp8AC0tf3QxKq/vYlpoei2U0WU9RESlpvhBVrsH9
vystc1tfcN2X3j9Aw9EnjxEW1NQfmTAaWIFAuWDUGMvJaqEBT7ffZb+YTr6FKzPr
U/sjIkD35KK5c3bxAWUm0pPUuKAaScS206fLkXxgf+fCwrWjieKagaad+qIRZyYR
wCQszcLk82qBlL+/H8wwMtF9IdTVddYB2e9Sx8YIaQfil7nVYXks97OqPwDJPO5A
MCN8OQC3STqVA3qsvC0xsQJam7G0EC6aaIT0DqIZwIL9vP7TTk0KKi2VbJHWaVqh
og5mPS/02qemB0dJVOsGJBjqraiQLy6KOS4ZALx5E8ohAIHiPM4yYigiVnZ+4NwE
ICeDAzyap8BZClW77xhb9IifUAlqWAbn11V+eqE0esECmDb2AB1zeNZAvtBt2MEH
xMNPeBPa4Do15JU8HnszovVB4gEhwM0no66xhGPGkAbVn0kkVLY3tZQarCnkZm6s
`protect END_PROTECTED
