`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rCCIMHSZbOh3GtVmLMVFc2eNb1aBNeBURT0MRB7fJUrr2Kt6DV8EWvMx0eQsIL0J
5y+BL5/lvn0hOhlxRLCol7uIuG/GBxpM8LXMN43iRRNCv9jIZp5x49Vn/LON9tCe
4unip7TN4DgwLzTqfIY2IOJolckJv2L5Wb+kP77tv+w9gRgZZ5oXpPCmmM8rom66
RlK3HcIMid7v65Ya/N36Wp1iuPUiLk1gXddaxzVBHT6HBmnl+SUnp3gmkNMst73G
sUfBbG1i6jH7QvHK+e1ol4qz6boOA/5xNdSTNUXZveRNdBY9ypqWR3w3L4wXVbGb
UOqlaa4RAexmGpmY7Dst6PQ6lrfPPNwhFYvLguxj+WCj/HjTNr8T1HnhBDIwo/09
b0XqBLGaXlbwvYowNzX5befGlluOHRb2naKm/L7UKQxDoAr3peK68UZslSqtqEkI
`protect END_PROTECTED
