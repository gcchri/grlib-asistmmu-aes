`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bgh8IPH9UuCLpyl6hSuEGXbwwWp/xHXh/QTSsG1TZb6tj1fVeVot87CtxrNXQfSV
ZVsUK3HdaG7qJe9metr2C9Sce8uoqXrqCBmienmhBOVqrkGuz22kUxjY6wkSch5B
sIUFUd3+lEdICF84p5E2K8fEKLvt34ArLNLmIlZblgaksRY+72ah7khy0+macvkQ
6ACRIXahdtxR6jsby9IBoUXdZsHC4j6HfNNdBQ8inaZW7fQuxM1bjiGTL3hgbIJL
TqEqNPnK2AE1nDhFgahhE854h3cKgli9Lc1lA3qKNCInwjn+HDwhWo+EjGrVnyFv
ucQUXP+jF3fC7MGAQ9AQLytJuwOXIA+KdWciVSRtrCEqgLSeMjd5XJC+tpIrNTYf
baVtaicx+awQiJAm/r0OKG5zE19JhyIw/sozrmfPb2ZcuduEE6lHSKQUqTurZqCa
r3DqlevbeKjaWFnMfVOWldqKKDHIRx5eg9UXXyVTBtwd+1vaUMht2CBYHs4Tmk6f
kkyWCutNrsPPyxvZk7D0DTInFaW4tn+6o/hNQQMYBFCc1OgSn7jTN33U49rq9KdE
DCTNlsnwMw+60Ju5ZNew7Y0zqvjfwXS89LHhg5yy+u4H6RCioWmyKPqJy9QLQOwi
QcjOj2Hkt+XiQPrSjYXOYf2z2eN4rmN6IgMnr4/XR6EnK+/TUw5+sQtfyOb4pt0G
Uh68lkTp4pMyX9WphuvThndngp7oHogegimiixn3A24kan5Y4BfFCEd9XMNarwEy
tOU4qxDOxT58uLxrlmGhroeXniXDG/Csgn4yThRh73MCFwmW3t8MKfsbtDqFzxML
Pqg4lxcqZNLyx6aV9E16vC2cFzmg3BiNcsW7DkiWFvi6NzEbL/dn2h39xNtL0B69
U4nl2lqEb0DyEHJVP1wAgA==
`protect END_PROTECTED
