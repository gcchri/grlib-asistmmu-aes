`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
soqj/k6PmG2ShhF8QR7qW4lYRXE8eVj8ofnM/KG5/04ujoDX2dCiz/2klv9bqtU2
/hoFHnQXDCgyCwiBFeBwOE8LkOW0/W3qxKMMLURopevLZRoWq5CGkYSf1h8Rsf9m
bMvhbY14nMRn+97kWHFrsKsKYIB8k/DkYuhBi98VCSr1ujWOFsGVhRmdIVPxVl+p
9fCG5sHYsrGGZKwHTOzjV3bCdqMXK028ZUw2uHxuhU5KgzehzwZ9hQHPi9V/4ZRX
wilw2tPbGNlvM1+XNyTlVjDN7tma6i4PwNAn5PfBIfZpYEesfa2DxcaC7k/lUhKR
l/M3Xc8UO+czq6IP4HI0N+9V5lYCpdskVVWL7kfNDgRsJWnSMe7Khb15fgpDF1Oh
GBwGapP12hqk3BIMxw6l70oH+YIR/6w9wk+DFKAhAsZoxE3QGMHZS+eY5/oFHXS2
`protect END_PROTECTED
