`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1i+4JNZSnjqdQMdis7Rf+H/jBqh5tL4IBF8Nt4HwoevqCpCiCJdYwqCWEM1aIuI
+6IzOomuAUsHkm4aslNGIZEyHgH5+CVVqZ2V6zf7wvNnC/PNPXVVutQqCSeMtyk+
SMwuHtDl3dwyvUeVoSC3TNk0LkUk4WxIE4YnYh2nR8PEMwu30mBOU+0LA0n1fzTI
npzmJ+iyszcBJ6fmGaGUf+kJ9QM0K++YQvqoqNMZ1+nFhKitBpkhLyOdE7UAklyu
77Lhht7aE/bGTvb2D14XT6AKt/tjBByb3QUkb+coRHIg05r4714d5lM/1Bc42Xfz
riKA8FTzox3ZFbTPokDT73xooX1RhuLrKM+V661p1AsbWfKlYbDfNNGRuAhglsGO
9V6N9vqEpth7kdSs5ECxwFxblsrlAyI8FCIum5iW4l03zwkl+9J/SJPKPHEuuNnw
/c0Nnlv5FT4GJZsx+2TDNnifwNXYYnQ9xiXcswSW1of9NM2mUMAY1kf2C0AKgLwy
`protect END_PROTECTED
