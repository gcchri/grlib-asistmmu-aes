`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2eHLOwoigIxRZkhmr6kVmU/64BCNfinL8P5NLhUTm3la5RwtW0ENFOcagU23M0TD
I3dcMcyiZk2z0Z6xoN5drXE8wcqz5NOvacwmXbvI/OIDyFfIaSb6VkKremMTeO6K
d+iaK+bNO3Ud4G5AKrP8SdakdFJnoacvHPKGk/xC4qKSMU2h7sbQk9VNMsXEx8f3
/KZB42G9zS7iItl+Y5Qn6CbqPhODRZqX/aoQYKJ74+NybmQyx791VJJAfMMO46k+
Jx0nx7g/0ikUw5/QlO0ezCFyYdjIo87RPNPL0RpHTXKQK/iVw4FDYzEERPE+jRcR
HIvn48bmcPD39IfKnUg9xgZp3jdVLLuN214GC7Jd1SC4cfbqUk3ukKAzwEq6T3wj
WXqIFUUpX4pWskwzpOSmqVBGa03nuMZ8LeTOp1flPv/5o4Y/clFkE+dtHWGyxG75
KNKXDEWwxMXGmJf85M7suS4fG7tLyiUM8MhvfE7JHpteL3kWBqgUuIE6L7qAl5EP
R7MzBEWdnA/4zrODtEXRp4DcEr+p8IfQytVhGuAICLKzawz87MvSiTNWvBQQFzAc
cRLe07okqCQZJ+diYmUrEw==
`protect END_PROTECTED
