`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFmVrLv6jI8e19LqubPj7i13tUxe/e+ZEr5lyfWN3y9PoBqht9+cJZ9Lz78eYstp
/UVqukb85m2bq1E81YdUuXJSoDtT2I2CpThwRqi+9SLJD7H/Srsb1krnhrOWDIOE
kZNNCFaJclmDaC/xNxTJeZIfbUBugLoPfXMK4LvGAMQC6GVyGn0jptQzqWSupj+D
8dKXDQrzN6hLYd+S4U4TXhEypFPj9g6SQ7up1LWqUFaLTMcTZDqGvz+lcQSKL02y
DVV3Wiy+Ayul0wH9FkOhe9aJ3HNWxYj/TqBlsV0QBV7orkUKzD2D8W5l3Mk/R4e1
09CRFYVwHu4Eizlm5C2SkRsgC9fgtrz1bbKdUHAxYtlkqDoMAKbQ/XDewLRXSsnF
i64DHOm3oE1zRTiYj5M4wyDb3xJcfTL8MKpL4PZfsovHidanKNajaNjLFOgE0VPk
`protect END_PROTECTED
