`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJaJXMNg9BgScJCHceiApKKYEBk8s+kWAgNUV4ScbTBTq17R5xypWFim7AFgez72
al+3BNwJ2j1uobDtusIHwaZ6TBlXdETZgrYzH7B1ap4yjwzD+zL1n3yEtrB8Mqa6
aJ2Hl42IlZK/44S8tD9XR0CyO1nDO6DbjSL+2IONyvk+9rl46SLZBCU1UmsYQP6H
/Fpj/NVrgLNoM8TVoClC6hz9PchLW+owf7/4USGi+Apc3/GENFb1g+jAl9/xx7hf
k5CB+ee9bAjglXb//16H9Rw37hygnMdqRdMLDW5lHLOIDkaXjoeoYhsThJmi8IEN
6Kf5gbkGQknKohkLBBQ/ivI06q0qB64eBRsc73MkEJ8mKgZ9jTMw6C5UOdKVC+zz
UEj/rkEPm4/FQlEO7ZXHIu7lzZrLQju4l3EcIXC68KoZNCvxB8hohPaOkt9uqIh9
ahnjd7iusvsIo+tEpROhHqTkCk1k5Oyu8GtKUN3KSrWhKpLL0GM0ErFCezqA0Opl
`protect END_PROTECTED
