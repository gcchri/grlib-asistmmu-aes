`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lu2ALe0L/8/E3gAkBw6ZixkBJuR1fBNTD5h66jDJKGk1n6wqLn1cyNs/bLLAMNFp
EvZQhmLTshVEFdvhoV2+qJCge7cyf1YgpvWAw5NgC5JeJeT+qUNPbiKaYcEn5qgU
TQAv8rpVVETPYvO7mYPndPkfdv0qj6P5XmlyRWiUv8b5DLZvEy0+EfVYu5zyYxM+
qtI7BejSVU8oU1t05CJe5EVHxW2SApR9weDAcaFsceQbmkgMJghCdtHOLg/LMu1z
xlq0wP0tbhXLurqTsN0iR1Z0+29KfqceSTuHYhJrIN5RYC2qSuQs0F/XlPxqxfjT
t1AnCVtJjqfpopQBaFhxKCOhOx1T+YS6WJvBD0gsqPvn10XMO6M6vgW2maNDKgYN
SXfn4XwJKfI7F5M91uPjR2rrvyCJf8pcy7IYGM70Nkfinw9fiUTJNWVYpKwronP6
B/0gvXNf7anRhVo2JhRskaPiSn3qJfu5WgtpkaiTi36R98NIyKypDSwbSo/+p6iQ
CQOzsiIeH72H19Zi+WEJf8A4opZunrC7WV6dbRr3YHNQ8GK36qHsNI5Ts5KiVTrj
WBFd2ZIIVydVyS+GYQKGTjq3hDY5OlrchDBx6KlrRwp+dcfFSkI315UYjchFfaYl
qUdqItpE5AyBNcfhZzLCO29bFktWs3g7tXWQ4b9M6YCPvSHnSOxGOaiBoBAT8taE
Dlghy8rhyVeMCHyo2OFOE6Gu4MtLqxA4xBnJ4EvVWaB8Vo8y6lmznqP1XPOQKd9x
SPEMw70XQEmruvUiZWpFCguPdH45zoOlu1SuE3n/mAodBF8aJ6mJUT0mlmfvBv2p
Hx4ZUyQE15JbK8jBM4dajPhjWn1ZQVHzUAKPM5/RUzpB/7fiRM87JGa4Rs2yQWzf
INcLRMn1UajhCk6KNQk4L44gCxFTnSKY4rOc9ZY7DIHQf3KbgpW52ernFaRgstNS
yI8pJchUDo/0zHeRFF12IEU1ZqNXTpnuPVgNKpAGs0rLDWrOZTnGBECjPHckDmwU
Qlwk2oEs9gZ5Ik11gYeCXkw7oWHVxArs/yYwQbdrt9GP0k4dhkeqpPqW4jkc8K96
zntYmcuy9UTD7R3cegfvj3i3qNxEYPqZQdPsB631vbk1rw8fj2488W1PglYNzJJc
bwHx3ieeeoFNj4aDY29hQFMfYx8l0iCQPdtrne3FjL7SPjXo6SyCSx+p4AO4Vm6B
z5kngZqv4fEQmh62YVyeMryILKmtfm5dMwRh55XAnDRJhEIhulaPUTwf9ntnzq7V
`protect END_PROTECTED
