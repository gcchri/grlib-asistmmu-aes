`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMkVv7JU9aXhXP58BP9UxaD9NE9oydPg0YJs/oc69TcRz0IOngymT6LJo+hy/o4B
h7Q3pPcTPwQeENC4aQKa4qOwuULHPHLChwh1K8KP1BVysZe/mvrf8InWRQU9TNNK
l9Yadz+e0NCg+CqJPxyjcYFBpKo+AKe2wdvv8yxHSMCtuc3NrC0uyeLONiSe/8Bq
de390gK2qsdtvFvmnTvmCrHevEFozmziiyt1E9MlP0Z8DUHrn/DQ6N8Eyni8kY9B
u4xoJsyyHWr3IbhtXDEayl29g+Cs7uP5fgId94QZRappyym35NlsAmQsOYfr2lI4
oGNDhF6/wMu8A6XhryZdJqVf6MpWvBFntyAJFPO/3XvvotQBtUKewS/XFEhT5p8l
CpNGl8dNqa9HPOCfUfkztc1mzMaV2j4TcA09pZL9hX6hEYcpHKkOKR5fBm14ywzr
p1mVSeKTyaPKEpN2tdcYo5+Uap5nRiL+H5GsWXj1VneHLZ4xi7Eany+Dqgz93BKz
QJK9WCw/yhzV7Jnbj5RYEidl36bgB0AWRiv2jfJtqMRa3UKSaFWX16NHGwt9nQdg
Xp0gZZaUKl7dcntY84kafL2iWzEgx5AngD2tb0AnheyD3OQRFwkbYLEtvVeJTBLR
7bGiqEaANlkE8XVYaOQpYspmkuG5c3IeeEwvnn0HyhMJVnB1AcMEAkRdp3NLhv1g
i2/9yOoDAonMGW8I0VDVB2Drk/x4co6t+5hWWYRRD6ViwGP3ZXkePEeANKF4c8id
dFtTKCIGG7TsXTBXvkxnMUmZXj5Vd5TqLS2a3TEoI3s19lYWxgRbi2MLjl1njWbU
9RuzPkJLJoUTbksCXY6eSKTq8ju8BjzAlnpF0MC6bu+SAo6GHTtEbTnWTjPGzRwj
jNI8RlyfMg0ImRkl8W4w79Jf+OPvgRyFxmjnilvx+R6unrVMzQjl2aLguZNA2diu
Y2IE/XMh1wCYO1l2dhIouEwh9dLVyQcRwjNcyY/TFYVbBg4HPEDvtwzn+kx75/Wc
QASoq9v/ng58ArixNTQLHFo2Qnm9ghcnX7QI96+Xn/tDPCSvK3TcwgkBFG9qowYu
Up/6yhY++YpQVfbh1wESJ0aMO6NI2+kJQDmNAeAS/5M6W6eYam6ZjGMZJO7JoMmp
HZifNE0+dJE2MJ1FX5Ea9nrAnBThEkgxMRI0y/4vfbufao90AzCEOXDGAgcaE+gi
Asg3RjqBwdjTLSYfr6Q4U4BXVMTMQ4qIXmT/RIWrerRkU4H+B1QjPHpukv3m9uM9
bOIDUHt7pSgTUR/HV0N/o1oo27++NWQpplafAFbQwcE84CaD0v8Sy3Y6s+DgZnSb
V1mo4cgRCvxgFJ/7oHx+LJJmMb53WAFJw2SLITc3fQKLx8oeKiN0pX09Vduof34r
tX6dJ1od9rUSDdNVir9ofUi3X/XnSBTqHNZkxH2QtVCYHwwWrGX0dGWpIHeTTVlG
3N3BAUoMiaI/7Ox9sdWEbSBm+zENIbsTRoYP7OPpJCIOB6BRm4EANSoxB7o8iGse
u1SdrPps6/L1p/mB2SdlG311GMfOQDk/ryD85tGO9AiaTV7csym7hYqxOWD1T3hj
XP01g7S4iF/rqc/LCmiRXP2LouBNohNNCScPC9nm2jtpnxVsps47+Bh6dbV4kbxo
yZPnFuS2a24u3KYu+r80k2EjmCN/k4jcpYmsfHlm3gjWH0zW1/vsIpt1nIoJ5cIf
nRnJIsx20CO2ObKKzOyt7rrIhWZe8HTKPlxhuA9KtE3EzgQQ2GTjPPPyDjgbISjH
PA9eoJvxIL8QMnoR7m9OIJOwDNgsoFVqUUgShZ8f7gGUC9BZmB2bWD6/+CtMx1I9
PZsZzbkSiOZtWZ1/qK4XTgOD/gw6HMNcM/arDLbQh0ZbhwXFF97CdL1pB4TO2Rgj
rmmmQIW1bPxFStHITpTgcrFeDmrLPbqxjZYSE/oIn65LbyrRARvsScK501cUBfNi
IU4Psa2pupkAWNyZxHccxkMx7g8/h4xg4UyQVPvG8NQXiNwk91iA7PAx9u6wai7N
y1j1wriT1EuXnx0zkp0DRsOV7JHRRWslSYB0qMjgrmU=
`protect END_PROTECTED
