`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uje7qWbKOFQq+A8W0uZBKdMeOpgq6MvossCHaVZAhahESp6n2EjUgsaX7A2tVwDM
VdJOVoQO7KYq6xAZPwdeeEcmTDPgGC35qjd2KNM2iuPx0IneKsXytzEKI4C37CPn
aBUriToKcCbQsuHQvEM5giNJueOiO7fNQVOHoFiEwlbbKkFuMpdia0k56Vet9MM4
y3BgUOaKu0c902p6iqjbUP7hLTWfGsoeIoKcauyHrpF/FfK+F01fyEhRwwcqBQtT
yi7MT2ab2XkfOn8QoLJctlyGE7qoUG+5knEj5xGNQNpQyXICW2AWu02gCwcNa2Jf
822by2HjqJ76LTWUm81IyIzCLV1d5UIvoNyHpVppHr3Ur2GQTLFQV7nlMwI2nd0F
BYEHr6QL0jbF7kBT/06ujhy2taI++Ha0F6wf32wVVtaG/RN/KwRiTGHspMi1115y
nUsPwq2J3d5KLUmIjoUny8NLQQ8bVvS65m5guKprZAY=
`protect END_PROTECTED
