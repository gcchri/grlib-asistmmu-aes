`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iaGuWoRPbKqw43xv+qCkp8AZN84XuFcsnZ4XRhfJzYBJ8BsTUYRkxm73kQsLLcyM
Jo+wMYlWKbnEXKQMQSye2tKz1X6gy5zQpQWafNTWgsEpqe9R/pp6bxn80PMg6J9L
zgtYVnHYi7DodeNWLcuubW3VbSZ2m+caKdt33ETIBmNQ1Li5cnU5idNcKZyYdqv8
4GD1FOiFfr74TFtHEbF4IeXvUOn2r6WFxEyC0upOGZciDSIsUG/IziC+yN6LGyE4
hwucqaSHXuTSilBiA7b1a/3Ks5uYvPFx3vIjlNofnI4Re7vKrrkU90Rq+4BMCQZ7
Yh2Xh4ZGQNNOYuvXojPtLibSZwWFjtOpk2aTCp5ZE01+Tlh1W0AnlI/S3PiudJyF
Mc1ZmN1VCcdl1Q45V/QhPAkIoyyrxccY5kBr1D59ySSu/wS9S6bkphE7BCJGhR30
XVYMasX+h4iTvYjhr7/bNVL+JgHpzno6xhjTokcHCzHMAhbNLdu86XpiwRfYCIlb
LydZBk0Q5Lh3u+Ed8FHej++5zDs1sVTZF4TJYXx8HysL8ti0fwWtTBF69IQpih8y
QhrG34I7Jj0NL/tbhbOfz7uu/uyJNDjvTHaWDGIlEk00AGczSrQGy4NZkptmTMcD
H2QWKiu2ShtMNGPl8DXVgG8754JSszZ6NISfI7lKew2s1TY6o6X+DNE+vuW2jv0i
6rC4SdJz2NcEB6DOvheK5OYl3RPoYHt3KRZ5tbj6pZY589iMUW2raVPmTryHyp3S
qL/dhiR3c9P5c0/wDCeXwetg3D+42/lnAd5WexFGjcQwJ8vFCm2xhVynpGlR2c8S
cNrUejr0N2kX6te9Dowd3YWtvMIHB2D3+e0y6eCFYYRuJRHeWRTDBtnRVF5hGhYt
L3AhzmLrRKV+igILESCM9R2l5AeA3bIJWkt2JwGkKn/srIsSKm6WzZmMIhfVv7oS
bNk+sDGnxg5ciFk5j3jhdSGqWIn/lEU7TwJvxRiHOpckhaU2oGOSW3Nr9kCAhBzU
Q1Yiuq4D0S1lwnq30yShqQT2Qi/UqUmyZjnaJPyPT9a360I+nuggJl/ns+umpinb
nBB5RtzsZFQzrEPi+UKcmg9WcXMTTqLqc9ozRuTF6ETpNgTKGoqo8hianPCLnGm+
Ul0OjAC/qiglrSWhzCNVx+Pb2SocHbnDrrdaEPcL9pdyNsarYIpH/caAC8aVG62B
Tuz04Sg/BzYvg1p37bRDe9sllgVukfec1SgEyZxZ9s/dpMLCJImjd0qlJWhck3ct
OlJgOInm2M7Vl4hZQCma1J+ubEz0WkQ6YRDMnCCwWdIxXlW5SOf+rtcsYNIzih5Z
i3Bu/WCtQ7OuzcR2bpAhPK2QDsVHWwSoCK/MCTip8vy/N7zACsqSj/goudaJoYxW
s25wIEfoNhj+COrOoOQZaVQIPSpv54Lcw3YO2cKItsGfG9XWGdUO4WsrX/cZ/Ih6
vT9i5omASaik/7fdrLpCLVVNJCRhMSv1vPVpeR0d2IAu2fGHKpeCdNoIUp06cAUQ
DxODuDU+rlVtbh2lebbd9SIjIJPW4bWmn9qkwROx2yH0mW2H5gCfG5sQakwwok4c
OiKtvW0mdjheRC6lvRCSK8oWKner1Vf2qqBl6FosYd22NBkTFxw0bd/9LpfAUhNN
2Z0TzYlf1H1HXyTv8S9qeEbFTWiFAu0UAgyLySbGHfEDO7Lcc2kgoG+p+dJcdayE
ge8AJZvLadT1WKrxfHrZTGToz5jG3Jdj4xkelnxAFOI0tb7pQuoutzu7ELtsVmuC
6swvp0Ofa/ExBodJoovFFJU/B0LeK0KHDbHMk0s4m9xhPcCnUwNBMWEw5nfSycA3
HNSaEP/Hqqh9tnuoQT8sJbGvinSvF7OAG+O4LSSCRR62AW9s7J/OvWzhTkhlZmMq
nlu4v+Gw0OQuwlHhupxXO36nZ+4Ng2CEkbGfcCIsGac5zOwJT/M7qFQXM69Y+40W
`protect END_PROTECTED
