`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1LEHKZO0E8Mgd7nfBH3fE48qFZvbrGzNNNoVMiyc2WL/4tT+8S3BZimiFUC/VOy
p+ZC9xJ7bn0IsndkRwvHae31gG0my2qzqXqMW37csVLkWEfnss43zmD1BnGRhyWQ
Mz3PnI69XIPYEncsgrdbkyoM9V6oMy2NK0yukrkpL0/SO79qvZVL9CQpo9wIpQl7
uqWi1K3YDINLLLfWZzjUcIkXivjHYSElhYsCnuEqQ27oV6EXQBpnbD8FIoEaoFSp
k2hXUemSsaIlj4PhocYPZN+LPhYk4g82J9AZ8tsxYDFL/ieE/isc1dK//TY5dDRg
MHPZKOmGGIkss/ACrBHzww==
`protect END_PROTECTED
