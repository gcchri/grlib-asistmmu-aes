`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBZawpupla4hqAhpMUQPq4U64ePGAQITB39iYGuXLrupXjZcE+Y8ldktR6VKhKMk
yOAg3YUqan1p00/lW34wVHzk7k5g5wkZMLIotUSI7bRCSt6rOi8hwbtTy5/skp94
ISUnQcMf9AMyg6KZRQBu8pb7JtY7WSnSidY4QW50Ov1iOBSFaHYecRkIQ5b2k40r
eR1c8KUAI3ZU3/MfWZqV6tIbrX10NjHybpTZ+9mBpM6uUDp5oEixtwLSfs3DM1RG
B3I3HIkSAON9xZtSNZkDdaJYgQ7/n/P8urpSYMjyB4IPUKuGgQXtDwkFvBqHjRk9
8yb5Xu5TRmxwpzAr4Fqwd9ZEetFcQLlFLByOZzk/LYjYD4HlzP/mQzFj7XfzH+TE
b2a97qxI6Bmp1Nhlf77RfrJPn93OxfkmFI1LQCw2PNgBmEHICO2Uvh1RI0hdVmOJ
yrqhX37Ry7QvMo0mPgghbNwJBW/nO+TWvEQtu7xylOc=
`protect END_PROTECTED
