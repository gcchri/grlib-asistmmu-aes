`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iOEl2CtjhFGsZ6pPSumeHGGowrTv9eOabUdhr8zAlZAQAxWuTI7wsGAIDiT8Ct8E
KG6bu/tNR9wNhuAPMSWUK2a3+noJaglMaU/JXz72cLHnkwti2PJeKdjnlSElWwo2
kBXXttZpndraQsti72Gy5fulyjtlaWZfh8c2crxg55Gze+9Yl54L4+bCmN2KnJpE
TGGvEHgp/wHmwJryVWk602I4GKURKXeaNWv+BA/YESteoSvTgivd0LON6vII1WXo
xC02PXppStt+LEoOilkreatNDELryynuZhsMLPYbIrOK8PPNcDW7MWkMCtrsTxiy
Pyy7Pg+fjStV8YRCcgUZUNBQ7Ucq7dWMlMHGBuCrtEAIzh6k2UR6qFhwA46lk2c3
FcfY3Kp5N8GW5BA5BVEX72wMMU9tvnHqXQfI/wBaokU=
`protect END_PROTECTED
