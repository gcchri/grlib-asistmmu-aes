`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6bw5y03aSYjuG6tAfJA3cset9yE+jLx2n8NwbrCYO8L6gNAB4h/Sczgy0cNu01kh
id18TZQGooMJqOyvhEiX+vG+i3m4/MTjyfN1UviULXakqfLgFqR/lpEN9/RQt4y8
Gz8XYgV2PzMULO4D58tP9pL6GBbu/TzsSno3YQt8irCX6N+VBBpF9grgY4nPV9ip
qMCuvUJ4SBd36b88j4rOGgvDVJnCQPLJeqX2loo6PDCO33xiAM3H9K52cUrOjT1i
Xcg53yOz/8Ph4fGY/Q7dzmsOBYD0DE/OdunlCjnw7zUGb3fa9VfXu/n/vHJTuQbK
ZTuk98tVFNVNPt7A3eZD4A==
`protect END_PROTECTED
