`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2HHILCzBjC6WOAfLZ36lzzKJVBLdP9yagdDXmjNHNT8cV7Z+tAEbx8Hh4fOX1Ie
ej4Y2bypSOKZXh3xi4XW0YRkzzLldqpNha9CZNC/cNcaLj80R8gKIymjVVWQLCvy
ESkTnxQViMzOgk2wfvPdY9vfJzAvoOIzPOOzlaTvDsbPcy3XLKSIlt5jsHzzrO+v
2VqdubDqKSCXYseyj06WdAKjmTDQhYPo4TffW6C0ktJ+LhxHMEsyesXg/Fny1X/T
vhvpZAQ8cqfzBOG+6gOWWa/uXdBqbDdiQgthr6SG0GpFzvWdlN2RjoQ7hT/tHt0y
nHY4j+1OXpnkPozJT5WTD2AtORkiSl7FRU7+emOsLzjSC7O9SDbJriPjUqbhSWWQ
Mr8ys1W7yNd9VJD2JEbr3MStIGqM3h3zBzC0Fi16Jn7Zp7FyhPNeGn6Fg6uXfk7r
rmqnBjdyHsHAhMqsyPi4HoG+wYa9XcRKIPkKsc2rFTIS5DlnoUG6S4bZgUiV9fwU
WK84ZfjdcxpkaQ4KMN9T4P4f3dPjMa782beBkrrQrnUDL2MePKSkQi4uuiLsLJla
E2kNUPJuAwOgrXsDqHqaBg==
`protect END_PROTECTED
