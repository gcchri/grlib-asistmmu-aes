`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r96x/qktuKMiSZKloZAZoKcWBYYLS723K+HYY3qRdOl3OYZc4IRIN3gB1AWYVBSq
XldIE4PEVmVtAOIdfeZld/eth3tgfzZtPR1ychpCpfLsH5ke76i8OFltaSRE2qer
cjeRsZHuhQKCmWgP1YFhIo/S2A+/8L43ssVP4VR/FP572yeYn5XJBKqduNfSe/m9
DN1HYsTsnm7fEK8f5ZdFRgwRihX9B0HUwMjyvXOcsNaErxzKGKVUi1PCjD2tTFxL
C8bmU9kK94BVPis86SGPLRTVIhJsOIbwwlkrzRT5NeHk9n/KrEebdG/kuSpUg4J5
8Wy+PYIR4lkzrntS/4bWVY3Q4oW6PYRUVtE69FhL7NNmggiKHmA/1cDHFeZ3s/ua
1t7ZMOOsa3wZqYDLayVRGxl/PhhyVwazP0nDHSVT5aI=
`protect END_PROTECTED
