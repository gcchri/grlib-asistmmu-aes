`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o7QIukw62kkm4fleM4qqJ1XVG/zjOzcFGK6IFg5gkM3oEWJFo/1vHMwTlHv7bEtH
HRjkTetAleYqWuy4uQ6kw8F4ZdRKdihJGXX1JxfYdSx4lT5cvzqsxPMG819w5Dc/
5ldJ0OhbJPjvxRapxPvjpu6kZeu7fedSpNLRuV+tkfIv5sL04z/014t5za+OFNb0
xCfkswMLjEI77FjYpO9xAVuz7lRHOnCX8Kmgd7r9bPssU8uFCeyFlHcA363RiKRD
v3w05ZYJo8z0SPqQvZKNheFRHHRmfypyNdL5wSM1lXgzQApSDn/gFc8IvdayJw9k
KDl/G4psJfgpuE5f+rh7PjVPSS6rrsTw83OncgWlfuKOeNgqvmDni3XqaJ+2t2oY
qaIlQ2Xi0WbFFaatcdaSxAVHCGZVrBMm86oixcrQwCSbLluBoEYk9LE1GCM/d3ak
Xw8/6VqVzCsWIAsHjqf2Qlr/BziX8FPDiZUKxoOYh+gyiTuYgT8ujMJs2Q4j9GAF
r/bgieV3bY0RtU62JIbDdo5849JxkIFGZy6GavQSpfJLzUVhm/wBUVvLbYvemnQV
59VdCWtlODusag/HbuSPOtzjJrIq7VA631P5Df2IlW3KDCJTE5liZZyxldav3pxu
anHsqcZffszy9B2eJT9b+fAZoYqg6eBIiFmda7TQoTp13Py+pw5KrcY3iUDy1NZc
aXvq1DqiM9AZOqzVmdNrKS79tmcxHg+aDhkPqz4qUvfA2PnKz//DAgNdvvqFm23/
t9y8DUc3CModhRraMJA97r4CaQujdNoEG99C6SIS/PA0q4onMpEPxSdfwRAr2xBc
Nqr6M0MuLP2d7gxUFdnwDdug1ejvEc6EZhZ/JN9HqppJ+qjCJRMae6rW8krTkGDU
ss5Btkb9TVpYEBMUIWYrQIH1OyXbXobYp3cA7k5o3SIuKNm8jDmjXUAh6R+UfXc0
O/5jKBsq3Y59JIfdwFoHWJpJQC69hRd22uWns6MI506c35CPTPGhOSed7CrbWehc
121aE6m8LiLXhH4+A+rgV5g2zl93Z3AUahnJKS/ga+NiUkS5lj9XuF2zDWtkx3+x
Ub9zvVVW3zQy81kvxAnzK8GKJMUkI96WezkMxxazLOclJQcqInapu7BVjlWQ1N1K
sTGu3sw8XyJ9/lpY5YT7noIaedZOaZ7FTNNSWumYGQb1iym5Ea/JM2/NJQVJwhLl
kl+tYOyS1w6+zFeci7nDzBV4YO2wx+8ObtzMgBOjkoeB1mnMBxU093GvAhXJSn9k
tdmF2zlxXRia5IOB2714jOROm4I05fe2P34QqQB4pOulGLgOiUL/4UFF7Lg89o5X
wBkgzALL0aiT9rT9GuMFT3jB4c04YjQ+3fVldXOeHreXRS3oi8kyL5Mglycebk9n
hC85s2EbVdogebkz1quVbIj2aRn9DpFlodNEVx+6G+kh25q4w9LgMCiGfuNhIFuu
z+I69aRQq3fCJsC6QSggqT0dyPYBCiTgdkyJDj/h8lcgjZj+9/V94QNn+0BauIyh
cq4Wzu74cgPnm8ePDK6+qlVZIB2ngkgY+NO8/Qb4TNX6XZ3NCwieq+JiztGDkrXe
xl+kSXIzqFrq+BXvIxhq9SBwHiJmhk8x6UC1RSjGihmj/MSD+GZffo3ldQic7alD
8DWEM//OQRkuu/Tp08570GLe2KveG3PdQdcZforKDdcPtCK22akVsmwH07JBkCpk
coWLWWyxPkOLapr61rN8hk8Avm4nnnVkwPsHmrgydb4=
`protect END_PROTECTED
