`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0AjLE3d3n5dIP+A51DLXMPv71mdRwjb2Kc7FDTQXuOn+31f+09hZziq4jy/cvgg6
gmHqN8eQ/wu15yA44DX4L5LXh01jDDa615j6Su21Wk9jfduJb2NWUTzn2Ialn41m
7U076cACFpHsjyD+xRMQgbqJFt1Dq6ZZQZFB1ngDS2spyoT7IYCM6SP4WCI29amF
qQbcI4YxDsr5BQLN3bMuwhGG/VJtMbsROwJiz42sDfl/r7Q6855caKfkyoRz0+LO
IAsZo0R1vc0TELjc/wT5ZogOh8+2b7KXC6tnoo6fxU1BQdtatIsasVGbI/zaPNmL
aKbV/1GeJtQGMXdaBHtX0ufNKP6K/e2Gwl1qq9VNkLxPBRcJyLgyhx3C1IdsMVZp
Ibq1Cx3ueGf/vcJcDIy07sBr1P1SqW7679apcEddIbBz+xD2OyssN5ZGPn/8E3cU
+9pXrF8TwTGEBQ9k2xgLNA==
`protect END_PROTECTED
