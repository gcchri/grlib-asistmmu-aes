`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GqWwgPaRS2AWgIcZFDRMNGLSfICiEAgtd8x6QgA8YoC2QR+XojDZzFZrw3cAC3V
go3jrt9zU6FY1jlSt9hxqrasZiUMc0YVNKxqLxeJ7tz/S4cuABvSoOTRJ1TJTwYl
loq1Wc9yHgOVY+ydivaUcvaUEHS5Ricj5djKtrKAoANHTsiRAKeUaEfgZoh6hd9L
ZE8fnRMtmQLyLOQjG/eFSoLy5EGecUAKvAlKkgVH4yY6h3oKYeNi28NuE9PEZfZn
8wbEfCxgySHmKduc924ppGV0bJ2j3096HTk8t+wgTr55yzNPPscRGbDX+SWhNAHP
Ihu/I35B/kkx4PigmHI2uEv+c9REplZgFjOHjsQLyk05fsJL5wM2shgiBg/yR+5G
TIVv47fJpDywB2DgjJg3w0Ihp3Dro/p16mHsOdoU+zZEKPV9X6SYEYi4zDfW11n4
R0rQJGGYDDd29m51U8b5BD2+6+fEHKL3KoGEgkXbdgr7Nv8Whmdu6v2ff+zWtxrs
7C/7e2573PLRiJ/0cIvTEo/hc9gKjRm455h5xFLHrgxCbrY2DSkP3Oc5RJDPy5aM
KjHJOTS5JGuSz0NNcZ0myNfWSQcYgPLo51Hg0NEDAFlZIaJouSNePBukpboJ07N/
i/83eDkiFdXGbZMKaKCaS03rOzFsG/CV6/TB+OQMm5jeoQQtclVY3YYwanGc34F4
B3RpTxKvYd1C5yPcOs9daq5Y/01eHKT01WS0VUvxaKqXMI8aGsWbGRrvU5nGSFT+
j1b7BaHlAh49bGpRozaxW8wrcjHGKUDqjdb3ovgl6HEFkUq323UgYhcIXww1WWdE
+2EQbLfGc7K2aNzlaRVH9VsAzls1QR6dsOOtiih1H2XEywOmt7w9ZKlsnHtqoJns
`protect END_PROTECTED
