`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tg6A0a1lhcYByF9e4T3xEGZPDsqBGG1+rmNcAxBCdo4/PJDZhzcR+b3q7jwshgBw
mIjv6P22yAC/vrC7XdcYa4XVIaRohIVN5pzJ/64pm7goDYd3PM4msR4mMNelS6t9
1xa5il93gcHQGBsGEOax19T4AzgRlq4JKUkWCTTUxJMewtg9E8ycN/mRAxaQ9Y/+
quD1Uj2KGyFT4uw7e8lWLU4CwMm0OoSkAUkk2NabCACb7+V4BYAifAJF89y1kPUE
MP0+wQFLkNht6u3hUzo7E6pabiQ/W18OP8qmdii2nkJpMlwcGKp0yJnnBpM8W2kn
zP4HZFmDW9R1+0QqAzwvc9b3e0ieRGeR7qfhPHJGoulUBqbBpm058iezd5czhpfw
/JBAE58H/qZqeFGWgcJPsPXi6nJ3EO3MfuhDPKNvB2we3ibcceVVe9zaWVzE0S2t
iDOo+HMuBO+b+bFHQvF4qw==
`protect END_PROTECTED
