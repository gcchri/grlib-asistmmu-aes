`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uSDO91riG4sZI5TWQDrQs4N1I7PX0qimwZOthBj0qxZkoFo+Dh+ReZqbUY7rIfIl
kmT3E0m+oRGV0lMYtD14meeLtX1R1KNQP1dnKcp6HRin5lQ/mItD8h/nnirfjn6Z
Vo33DgnJknovlcMFteJjLW+6ltY0LndauPGdS6geBUsqIgRVnTybR034M0lq7jZf
WoqZqvS1AgsxaYcwQlMsJuYg6Vw1GipdHV90wdyCz1Rjl9gpFVwVkkINFKa0wigz
AMx30+8/VTscg6TE+vjqcLhrdbgaouBICiunkm+P+xokK8s1idKAifh9ljFSXeOX
Jg18LdzKbu9DsitWe0CVWtLMECeaqkr0W3oa2LenKiRYCoCrCf9u/k0xZWXFsXsZ
FOjTG6DY9uoUyd6y7N5l4w==
`protect END_PROTECTED
