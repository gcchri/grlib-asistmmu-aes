`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0fk/CN2t3J6c60iVDNUCfMg3ANHw72/T2dkIC4eO+4dLmtRk7ODLj5jysp4rfvJs
JnegVQT0hHuh4PwHU4fI8DDNBUg9P1aBNQ4tCsZAxqh58SSHXMsvNSKp7PHWxvPw
nR3TWWmZIKRu3L4/neJfgoFheOSESWnVbuLDTbIWdUZzQUXYl+KJ+gvzj1PMzdAL
6kRfOOYBCtgMz76z47LM/8AfzQGNGNmENLzWh4525MlNgfaToVFYMTRLqFBJxZAs
kag9doCjWj+sb8787Q9u20itIm1j4KIF2llI0i0iFES40n2vOudYHBSA2nghLS0e
V1H/JPkp4+6Shrj69qbVt+LOScXWHKb3/dpj97MAfZWiTPy9RlJrR29Q0OzPir2P
v5+E/o8V6Hr50fxG9mb/MKSewN5MAVgNg8xz+38jiNnvmQzgQ61c4OR55J5dtH5M
5yZFxtS9LxfW0d98z4jLy4F47AbyHQ/Mhw8uGmcVZ2A5/Ve+LJv4wiNQobNBsvdI
EIEwyy4Tn1K9uZAZC8rzA73qIPhZp2b2JF5H5g5v/Ex5uoEogORqOwJ9q+urDnjD
Az5TzWeHFWmEjgZndcb/D4FAUerLEsd6pxG5UdKAzb4PJuRX+yg9hEvUsMF7K5c7
IeZFYPptsfZ4Xgx0W6mkixbupqLSEo3/G0TZCoinDrviyB6LPX5jaCS2IT45A2DJ
mEl8BYBYbcit+V5Erj+2frp9XZFHEQWoS3yWMipwjALaDAGanGbL72+iv06r9Ncr
s8W+2ViI1W+LPzbqyG2xx7tmJdj2e/pXvPt6sgqxKk7Aj8QSZMhS/tXEPC/txx+n
2eAjQBFcCKwNMkNCWi2TG6l+IkbfqGaw2tYyY7tdeoavwd2i35cWYlIrM0g9t7Oc
4QFk/4Tw7lAlO7OvB/1a6dLgNDZWYlm/lfqotjn1ySwCIZMNWH6Vs1olAB3EmrVi
7PWHihg4nJObhfUjk+2zSaJN0hp3HO67p4HLXvXKR3ODYgOuXIxdC3pAj9bqTh7z
jIx4Df206IugN6JO9lA8TW7OWcEXTyE5lrbfVRlrDMYuApf4BcTFvWJ8LWdZ+her
H31yit4CZMcM9AwEopz8omnJr/JFHZF45if8a8MVgQ+ySsdXCVyAAI/sRroUFgMv
JblmteZEUgftmPlDE/GSkj0WUusYXdumpzPDJUj3Onc92LsfHJg7II5pO+3hTvlI
8ypZ7V1+hP2w76+JnbRMUlI4COPY2JBor2BAVAGNImkwxKgjNsxq2ZmaxgiLNP9t
65sBTJhrvwRLvGmUjpZdlSuKHRbC+Sz5lGGZYwMGM9UCtkWD72NXptxQt8wlQDQt
h/MZT30mj/aPhnxsFjH2inXAdLQ0EIpifeddNlOU4jO6Y3VS+yl8gRi6gif5pQN/
6MCZHImGk7wrQU70m8ggEQaWWo4+TUyeswY1p9OuCbDb3fZRA03POzkwfpTz5eMd
XERP0EKxIg1+cqt6eAdodr88XDCT8rxRonOLIT8oPwe7jZwtSWP+TIfF9GSkNjbs
hD7vFveJ0lKGj7YGJabGCzkHdj5b0ADjeUQ/q0/y72hGvVKeQArhg2rWmjGo7Sqw
ohR6uXlJy2uVxUKB8YEwfdI2TdXm4pW48zOd/BnQPFfgHAJ+/vDJJTfT4HjpBEs2
RcBBu3MS37X+Tl2XlAzPdd3isGR6hBtciwWP3U9PcEBpk8RBIm7no3KEGHHIlwdj
PQNwzkl+gNamr03JyJOYsqPES+Utc993Qvbs4RoO/7HVFshaP2ty26Qhikr3ZZXS
Ubu665DXlUDfgCmsiojIJm/kSeSjxAFXXw6BT2dFioRJ3mFMDpy8nF/Tp1E+0Szb
+amwnELauFxH+mJ8fy2SB2Z7lpl9h78YD6GoDc91JeYDOLQ+8uoGZD4XRXADlqqD
1KP1wRswXbw2rOUU9RjOtr6/Ity/KhM9yeo49KeQuO9KeP2JToZFEyocjKX9iwn5
wangyB+Bl/jZKPEAZK5xu8pUmwOK7yjOkrICqtL32Le90ACJ6v2LSJUtqcU/40+M
g6OK1kUr5ifTBuY5HU6u8ORe0Ofa/9MDgCUJyfhf6qHgvkb1FP7iUSDlrt4wevTF
/DDTNZP3HXPdqKKtjSB467PmQwujkDgS6bMiGGuzv86KKOzXuN45dMaHJllnYEvx
Ho3pbUxqmdnQ+DHEJS4Uq5ElK6muVaaFWhY5b9+bahNeqCB58MB2c8IbZyyQHB5Y
q4YMYEzazlKa3u38vtuU9xj5HFcFMfouxAeU5XqS8ALZSoyVB+GKsv44bWR7rdVv
g7eMU8NzVgrhrPsNN+nJrr3LVmRTmPpOxGbUGo5J2kjohIyUHYveZZGQoEV1hV37
qTj0CezpuusUv1xSrpXretJa2khzL/7D7NT8vPQ7jNR2hM0zQQjqTsnnFb/QFTsT
/IChpGDZSaCzggvrsO2kkt8UohSWCar6RC70pQ2ozCfWjShUlHF+/VtoVpwHYIy4
pv2X2ZqSrzCCEjgM8V57v4TUGkjNB0AfB58ctaXqoGdtoai2Z3VEL7yeBhdXJfDi
iUdGCIfMkvLtabLn5NQPO8TyMHXRexmGxEacuWpumMYCiKwwXKyotpnP6CAUy9Vj
zfypjdxBJ2Ldhwo6+Topzadd4BWdSp3n385vMdYRb6Lj3220FlpHMJ5bFs+S2ipn
ub8wx4hF5d0V16CrFXf/1n+4MxKaZIQVmv6aTYTlS1ENAwqBy6SHfZPXUvI5AmKQ
JJrMjOS2ylk3IBgMFzkdGgFSdfk3SoRgFQ3DaYcN3Z0D57QIPsuWEFh/z+CYmw7C
q8BcMxd4+DKASuRbH3keeayDLMNg6B+CMaT4HZ5ZpvVm8poHqT/tCkTKOHeBL85b
hlsN+SBlY4ORjLcthG9qTEYw7WyoCJZGUiPLEgusn41tU5nqZchLJKAZCFbW37w2
DhA/3vByhn/zmMVq/WISX1zYoJvCm2nfhwXAtp7Ou/lEPvR7XpS9ocqgmHq9rrL7
dc4yJXRQMy6jThrG6VBhDKXVKTXURrqu6DW6hPGdewJX6VpM+RYw/zHLvpkpkYht
QoZFFvfPRcbr4bmmfTGDP4Yj6YGpam6dOYhuAfVWugKdGu4u9BySZZCyeK/i89E+
14WIh81w8Y32lyKmhOFGmgDQCjcyLew7/HziPV4Z/nnwFmLrZe9qxiD+X72tEmEo
iYCse3sumdt3D9/44z+LhCcSOX0nUGLZch9n8Mj6s/4YQMWZb0JGdBVyVFmR0tHO
D226mrdVic5HyiJD+Qq14XHap+T89RtrgUtsYzTjTVcqd43FqT/Zmc+kSgWFLXlB
/IF2v1MY6Sfa34UBCTHr6ze+PP4Ag/9MlY9bVzdyb3FFQAKrRFMnVwzo2vclZkc9
n4cZWRQNRTEJufo/l6mHbTmQQNlk52OVoOXOQadR2g3CyR22BLdBXyWGmd8sSNqB
C2j+RugotkoLk9Yw892iO5KlVMUjdfFhgVRM+zxZS1pPxDDB5a3FRRGs/JwR+iMt
GIRwK7F4Mqso4cGMJ7uximgjBiSc+zWn0vLHC3qcDJgNA/8F05QOjomI/7sh7o+5
gAqmCetuw4rzyuOJcZ5aiMiEq2cua8kXTpQT2K2t6CPfAlGAJGJOLkY+xLjGcVks
rd6iUUd0HuOHplJNPpt5pZ5tBRco4/XvXOaa03ENvqLsPzVlo5yrlIDb96MzGQYL
USOAV1j0PGJXRi/VruaHrUUFzf0+BMe8veMphEFb4rYszFskzt4Op0rmgwBBhrPN
E+R+WUDpzFMsTe1PPK7zmI8E0AwQUTen3nENunGBvRY6SI+LlDasFa1SLLfKv+fy
POlXESy8I73v1813ZGya5tCczrxl8emBA8zWwjngJ4EopZuvYDcRQcrk0h15k0J4
+HSIZ0kEih4QqYa2oVlHnjTcV8k+VbKT+mVQbjmuOM3c1wD3ZB7FHVNXi2R/HLwC
B3Zce/XBli/0Q+TkPMAAcblXCboApC/M37iKNrsqcBodQFip+MKEdhqESLpDgXM0
ZZS1wT/MpK3M0lY0HmfFhunuUDMxCWDcGU155SFWlwmTFwi72bXCxb06GFVCW6RR
vLRHQPVAztWlDUdgjIKWpZ3nO/Q6XWGvaUaZG+LJcbGYLyQVJgoOPAqpuuDplI1w
+uWvilZlb2L861KNkBVY+estG6tt2g8aNyD5fJPgPnZfyhjU/X16cUsWmiedkP9R
2+Rqw1RtmLTcsoAAsvOnW8aHM2cQ0v1eN8RMBr51p37ftn1zxy2Q6XyKhG36Plm3
gwfPeKR+d/YVw/3dPxu4AQSjT8CFYWQ1tIbu4eodmq2iWMAqSV4JDfPpZa7NLiyE
Dv5/hAQWUyD3Q8ADtwd4Y3I/5+eCPkRfESPL85ql4W1o4DorKEJqfs1sqVFiAeH6
g8OFgt19nyQL9M/08aZtxYWTSxGUQFJ8vUCsfrsPlBZxFJ5wZkuT6UFpDP5NxBad
edCHVQ1KmHrziL6SQrnKk+es0ONVc1lBvQiUX4P2K5KOvpTzOufBMMwRBingWgXD
KWqUg+bBW064g/ecRnTgZ4k0NLYiwZs66Uf3EwvghFjgR5IwMdx1KZgvtzwpoMeP
EtO6iLzNG3eheG9HsdtQAZZQHHwLr/VM50EesJFjCx6FPvusjJ4xppHT3Yjq0K3r
NVB3WDiMGOy141hRrpCm+DemKL6caaDhZOkleeoJuPeHbkSTz0NsoKpic+aJnoTi
BiOhTyPbIi7pD/7dR9Bi0bHl4UR1IPBVLOPa1Wy0/ZGlGechuZXaOF3oTu8EBhXr
Q6hcSiY/yqrIV9GCiuPeYjVca8lHiv4q/wqjSvxXqu3ODRSfUgAQsGXzpg0DYVm1
TstDjiwj9nFp3EZbWCvxkLHeG3HDRTJb/DP/acKWd67d4PyVBsMD41d4eWQHM8tn
A0ReX8HY6dK0WewINziM6ZmFCxFUzS17SJz4u2jIsZTuViovnDci8pOwjAtvetAl
059ZHtEH86qQ8jmtZQUH8R3sCZLWnUemm/4ctGka2UIfgauR0StHEPFlMj6IBKVq
NfJcb+IMqv61GonBS4GfpLfwp/lrAD0Gq3sZNKId9Lk7iOtAqiAxhB3tsICYaIoI
5HjIAhNME7R00Lh+5WzepVWPWeCUBSZEHATMasuo351Q0ITnEtgFqTofKlCvByWf
23L6u2mP7cUZ4dnRQjYIyW1KKEbbkXuNQn7inqLE/S3wZqx5iwDIZ46XBAne25zW
8zsu0suOVRuBr69KAwOr4f2m1fxNp5kxdLW3Q/C7gzoLY/bUSuoV6+t72QbgiPa/
Fb1XnB/hKXwrCfU1IXwOvQ+Y++zpbpTakxCaLRAxc94Xzv6yv1foGJFA4845Z+0W
q+SaDRqgXeg4wuY/vYe+RefFr9xbNr1tsqoldlrdo8ceP7tWG7cvfL00/gMvG8l/
WqszjVJS3hL03m7R1Cgxr1PaLUFlDk5P/LayuZos5VN3pZIySGgnWHQ14igknoIF
mq+cA321GZRCRTbUVn/nJAwgfSDHOca1oj+49FBeE8QW7prtluGEneO5F1m3bBG2
/j57d21BQfp11frN6uMS3NwkJxs7KKARMNjlrqzlmWIxhOvwD8yDNlRb+nCPVLEe
nn6xsREusUerUWLw4VI7CWPQyDY7dP6Xp1ALPOUyGM9hsOalurbz5SX1rsBaKwKm
OR1kPBTVnOJ5rXkzkSG6l3CcUJIEQRhe1qB9MvC2By+6PKvMli5R+f8176sakvPp
H6twDlxczOs7ByJxDRSgJEaYH/6y5HZjphF22b6sAhKi8X7E03F21a7ZGkF/NHLD
t+C6TMUC3BiCQnng2C2GZzeDlXf7poxDlNioRGSBfA8TohYAcKAwDsePpcAuRn6N
4Wn8BQhN+9/rCxUcEDygE5Zlitks+6PoWqZd8DxuywuMMFx8YJ1G61VjVNP1oA8P
sX+IoOZZMZ1GbaWZ9UURFmdBgt3sW8tCz9KNXFMC+HCXXKHXw6oAaRyS4hLEz56Q
FtaO5q/B1bm/0QCqugeyK1CGWA2b3Rfjbb/a3Kan0E1bJi44nIiV8nxc2G6awKnR
9rqchxFMbgm+CIMoXlyZ01FAzRGGXiPLCTsFp6fFlwP++g1tLG4JDuIKkP7AVZy3
4ULvRurXQAO2AgTTh8Abjo0M+k9C4T8myLt6+D0uWzWLnGIWnt7EwE3jhkEfWsNV
B32PyZqUsSx2Ux8pN/Y73hBQ/5DRQlgwnzSN9K1TnQBfNIlgnyafNPqE2EIpd9x0
rPFyUleYcdHsap3yKLPaG6nfynvzNwfabgAZShh8ZxI/V8Tk08WbAZtDzdyyAqiN
ECgfXVVcDBdOYbFSoKVTrfZg/WCdB8XV3ohu6gBlAFg5mF050nTNhgpVHkDUFkr1
KQ90MvyDCTPHJEHChclEuqvPkGrvjvzehGNz+c3dbHC8IlNrv+xmOG3x1yX8nYu1
ngeyHAlBPkJRdDOuNh6SpSZ5ZjRHPKwKGrlnozfmeavDk8PjzWef2xvvumgP3NF5
gR2NyLP8jefwZsWU2mcJRk1zfulMhn+AcPymNE18is1Y9zQeU+SMIKg5FGK35tXF
N66tU0+bfo6UIOq26sLuvTB50Kz+FeFcSxI4c4NEAqV7PRZtOT4YMRheAvCydTl4
UUHzpTKwoB0vNFJAQ/EKnyshiSxzCEslc4lt9Mj8fDjAHr98S4TxwkXuPt7fLBqP
rQG4kuSb3fYjn0zV/TYTQd8RBrB5BZTRrap4cNDbmXH1RpclO4ectauuOjGrvzHi
Ppil6JsrMhJ/YsGeCUf+JXV+Q9o39fP0vjuf7VVMxAxOtMxqhdTN+4BtRaO88k6/
QEIHfFpuqoSz2ldpIJGY7AS42DSZvzD+bG0brQWQ/2a7O5Iu4wbcp7OL/xSuUuD+
wXoBXrycF2TATtyrlhhRtCWN0+Q0jOOY6N1he5R/5JYO6gXWJNgoOwl9vOaksgXr
B3EW3/Neikx3krltibv3gjSjE7V6j0PUgMVL0B6ElfF1s2cS1BYkggOh/2bsD4OJ
ov74Bsi2XAMn6YE88AG+68+MPwlQiu3sUKgT27saaQ6BplZRZ5Mk66qgrcMJl7tD
WaRr1YNp8OOqEVBf5wu//n3DQ3Z6g67MrsXVBPNl1LTLLCTb3IBozYkcvVj8kj6o
BnpWsoyWdHTuLcnvBJLOIv3BCWrhI8NlWcm92MrRj0avZ2OrB26Un2S6T+eLOtmX
LlS1ptqzGUZqZ9UpUdVOmWeVTE5c3bX7IyHIcuEtOz9DnzTzjzMJzd9oPLsaUz4Q
UiI2cWHeyuhGhI8ncbUqnZVNdSHB4WZpN2EuysFRGicYo0PEUF8ICX7z5nDt2+hN
CFJ0o3/y+vcPoV6yCsmX7ae6saUA090NqxK71y2W+XGlwzY+7pahTYPdRmbwT1J8
+Wj3/vWPSdoP3J+clSrs5Wi7Qh1RAVxszUhNWXNnbdagJi9CikNiqyUOJstZegyB
s170jqZwj5ozqiVy49zZTvEyBS0fYuvuLIfpWCyGLsGTkPF9z4Td5a7X2m30LYsL
eQGNcokVEOxTdvSn8Xxlc+NGWeb7cqch2ajS4cj+ecJpLfI6bEj9q0gEJhMnoc04
rQecmntRM8JWCdKxS6m4bEuTUF0m0SSf/O/5ayWuUeqFuXOOh6N4AjbtV2ISLy45
CxM4g7gi9Ce7lW7Wwgs2DARGwaMzinFL7h0e2GksfTWoOsPgBYlpqiK4uzVb7/Od
/IURQqV835eJeJyRlQu8lnRw+GlG0j35nFLSsG4UR5pGBwn5rkZWpnbFhtuJCNP5
Q/jg5bJGsX5mVZyyLx3qVlyhAp5Gik5KalCyDO65ZjpVFxMzPZgUd+pC991rSHgH
yzpBbxJyuE88SRtGNSEMuEg1F9KCgdE1gPsm+0YWteiXNDwPk0EqzDP3ASG896s0
T2Fy8FHHxm/ue3a4w4uFx90fV5LOsLLNf/7rzQm/YtQRw4OxKGzeIQu/BadQL2l9
NC2GHvW2X66M6LO1yc2LzrZr/2LJaZkaDIP0+yeQ0UP/QB7SmmoC8w9WNGvIR0+h
065fTUMQNOwewpwwmqH0brNxGTKT5gxkQC9PwmWkVAUbCaFocDoAdh0Q5s0RY67f
qtcK8d03EQF73RZXVRrKPeQ2IOh+uvQ0T7RxyC7/eZ0NLagjj203RMgXhuOJDiNX
RrDZV16NbCZNNREG9lrPSlRyGH0x2GECrX+lkMmA5vn2KYQsZF0s1upQFqhqASWO
x7nzHtjc1BhlgRqLIlgNiXhaENM8dGWLddiH6OmKymXoG1t+TohB3azfl99zSGIb
smC+4BHKfV7rXBDy09HA/NO2jMipVuIxJtY5JSxYbr89TxiE/Y+ZEaa+nrMuScQm
pg0IWGFZeZMSJpn0MzOlkuo9nHBJLg3UABpRq9KY6GmgcZVZZPKj4fordSZSkDrL
hWOnb/6nfsY33l846uGyrjR/E+vH7uo/JZ+HpuJdUic/90LBbD+PpMPnUdZdyx1k
khKWK76pHmxPfHLDxxKpS/Afdu1OrGFbj/Nsp5qEw+00H5XmdagbFlL5ZvELhdQE
Kv7tZC7axWSVI7VA0dNVH+34piKVrSTpZX7PBjjLtbzfjd2mZ1tbY2+pjWd77lvM
nItse8s3ju97C1Ek+QRHDDDnwXPlmaHMuqtr9nfre/YRYApFNNzEACmfyhVBftPX
cfxt27ZPaaZ7e/xIpAo31GjdppF/FyvZFBFr+n3aatznj4BUNlh7+8rmrQ3hC6HB
ny5sqDsL9oijtvM0l7L0xbT0m2drwn/+MpVejgz1Ost6l58F090eK2XRXjVnRLMB
dFBf2KDBCuB0aQ4z+mCacjMrjSB2a1dlXZ0rtQBDNQgrcLbQ/vhq+lJBdLfmn0So
Qtc/1FkmsmPUzXpvbtLx+JJ+pYfjSzb4odlxQIo3y7vCQdplyF+wjg09SOQqOgZc
BeLiIGnFf6FxYDFUsqXSCpELdGlKiqEMZkkG3s6olUBsB+m6i2at7plaSq4Y3wMI
qabliCxQSgBkyOUJfDAsI+Slpt3cNo/L0iA2kX/y+DZPKUCwszRoio5U3pQyiSm7
O++/F5mOHFu/gORv6I71wfoCjw2oH3GEDWIbMswhd7QYJuYezbcVmb15+8cFp5tu
yNFb7noxTlQsAPZ5EA72Bayr7Mnyc+UddgkXdFo9LaQJxrK7M0q8Ig93nz4VgNtZ
RJOL3dXv5r54ZnOtJS6Ouu1NvWnDx+HjL9KVQdYC4Fg6AcT1xcT0poLMht4VpMsd
5RFHcOSrDmuaJJWMBMgq02kHbAWagr2oUQaKdYl5jPMVLJXjcWS0nlDOqFt9a8vQ
ZWbM4y+J7rE+ly3XpSaWMrExWIOto1trH2ReZG52yS7mChPMifaH7wowJQSrXmgl
Y4g4X0wv8RaHIE0kKNJzAQNnKNAPVM9lEjSPCMfc1mGExcAIa1U14nDFkwVfOTW8
d9css4nN+ABCXBqvqlzZJHkdUO4WBmZcnmfZW0F113FmICjNkTQ7y/XxxWyPyM1X
/dlpHibvKxrwCS72v9IVVnqLHP/Ssdj4NLRSnxm3oU16gacXZwsxXruy00iQAfuo
zIwrwrSdOv54zbJYnbQP4v6FfvbaXe78kawFM9rB17emw8RHFUxzei6PDLxOXegB
T71xvimICzRueEd2/5Qcx9MDUSqViCobNy6ZVibf1j36i1ZHKdHTCUaPjSnwZUyq
EhScV5S6qTydvBidqAUvrVBSgkyMx8KUbfd5pVSFfjq6hddM+Q0XOncsu9Qe3iTQ
e51dimDEFJu1SUvlLFkIjmPIpais4DaJqQ8gLi2Y0ML+4VIuELC7SlpUJgNuffhJ
u2VxPrj+Nhtj6xo9fdgEQQuxnFibn08wJlojIHNHtWYS2+73DNKBq56Rdqpf7O7y
1Xo6W5GCjAM4UtlH8bCJ+N8kV+1lZWYqfwpFMPvs0PbLIHof5YjCCmiIp9FaMgd3
ymrLLOHsXVZuTR90PcnN7s8ECbjXIZaYhCUNNtFWaz+E3s+xh5O+zJEh829RU6fY
HZY8O0tNy40hjrs97GNsHjpfZ2CeD6Ehz4PTv0RB9HTwpIWEGFCBDTdji7YhTRi3
l+yY9xot1eyDUhqQ+1cJkxm/CxmB8c4Jv1ItwWYp5W79bHGoa3wn5wNqf2PFbhFH
qxnubOE7kQ1jQ9RdtKR+d4seN6vb0evB9ZQ93JGUhueDaA211AWHFtJwpCY4/LlJ
+TDNJqJXUdvBB5yNWsNbpdgRmDNwshO5jm9fYElLEhJo1lUnnNA8A4mPLWmesyB7
kH7bVTPHEIkDQdtT3EdWEGldsMCgWZYN45ecrcMRlTBjwy8FOU6cvu1McPm7HZKH
sd1IKf5sXZdIRxy3cTAweJ3UauZyPJMO4Zs9abkuqXdOqDCE4bqDon2TSauSYr6a
uAHuvMPOQGkag+Umxk+lhH6Uf2CQUxKA1UotKMENjQoaKX9ZFd2p7JW0MACdfOsF
FnjCHkY+WiTNkeETR09D/f0RI46spUu+A4sCPOf4LGE69yaZh7TmW5zWYaTMtSZW
nlRIZvITqQRzhrTZstsHWFuvg2oQFY3WMfmmOtkU8Pm5ayC8I6zczavZ7k94RO0b
k5MK2NmhcG6zwPmvw19QitiLNPx05Pp+N4o51VStBr+YmrSG2uG/t17HTjy56NGc
mE4DSULQvyvQl0zjY8tKPtIrFnHpKvmo28vczgjuElc7+mzDAREC71CySgTKY/r3
hIzeqEDYTJXtrLs+eQoqH7XEjHgCh+BOlHfEKLEuXEm8I3Z+UYui20nue0TUUDXQ
Q6CHZHojdSUhb7wVuaF3VGDKOYxs9grHKTtHnsm2fE1XiDt114Ci7EG+2t4B8sdy
Sadr+PyzXwU47d3Y/M8c4YyM68TW0QBwR/ptyQoef/+NZXiFizZShLh3N5LMjbuq
BVfxsTHGQyXBoLujQCICZf997xweKYhd2U2y1WemnqkgH57E1G3Hkr0H4B/cFsEU
K8nPXrJxScXrvdWKEjqqk8RtBZ9/kVv7eIR25aojkpWTLsOeRG94ionf45ktDfzv
2RjZexfg4tm4fw3xUG1EduEixbIKqsrcjVQ+lD2A2oagrBHU/0eNVviHrh+EiCIW
QM8QF+1gwB+83IbEd/8yrJIzQMPVCzki4nrh4tWCj8y1n/u53akjQJZ50l+17EG5
CTx6t6n1TMTWV5z17TwLfpEY/YY26/MEmajoapEQEx9PTZxfHbu8BpEHoN/i0nSP
ggArfoi/t7Og6Sp+oI2PlRhn5iHDFz8e8N8YuT3EjleJea2eYBrJdByotIQtyiW4
gW2ANzOjWpXXk6Lrb4WOqGQnP0Oc14x2nLaVLxaEGEox6Uu5ktWbPHBnGgHDIAed
xp+yr0vthzqBbeh08iCWRH0Qgp9U6GwIT94kCJNKCRSWrd+do+LSXDXtGaseVCgg
LvAl7fTF/82wEjS3j/pu4x99Iy+gYojAQyz8AeWR6LFuvfAhmzkuMpEP7aptTksp
W6tq5uzHcJuOgCgU3cEDlW9Zdjub2XvWTIjh4Ukybce8qv+7S3soPzI/DNVxHbzW
U3MeYEi+xSAypYUXsOnfom3Cbn3Q+G/wLE0ogYsWlc1iGDImAS6GQr4KSmr38z+G
uRnohb5Qf5KlKfBGlHfpBqdRJmdx6nvIqhL8dBJD74z1Q+nGRk55EZpWhnbc8AlZ
1c9sa8u+y2QDLLPeG2XH2rUlrCMhLM5zR6IthWqkMeO715roUznufiC1L1iYUFlO
dkwdmPRAnEja0ZV0f3Q2AA55MxxKhWqHaQLXgRuTdRhy/Qqvccqu4oTPCJ/GBAPb
xOW7TZUCqbqCneqI5PZfwUniEIY5phziHM4S7DNXBSMcal/vrNw6TbQRyMw9GSDu
jorandR3gsjYkJuYtGTjUYdAYd8Gulda21jwVt2YdeR5QLg2SweKt3NB8fUA/Uii
FmzOVuHyxB7giZF37Nr4h2L4bUHEyJkHubMOHypW4ynQznfesnAp70H13ymdpEuw
GC+O5zQMNkriN+8r9WLF3QV9Sr7Q64NqBuqC2snJMHDLrJZuo+nA9+PTJf3aP+zL
0vKqqQv2mK4nKHEjuD99hDTPapYcnKHpA9YyPUqjuowgrAX/JdMTNgPM2SORadpx
7ugTYuh8G7jmRjzXTLw76zX5f36Cml4RtOBXl0YsjYCEafydU9KvztocVjqDFF35
JixHjzqw5+/BHtRWwSjLpAUJKjGJnJqjjnYtcxDJmmLNKGoZeLZvSmEaNGpFwZSZ
41XV6CxllGrTGC7sDPwiYqWYLKv8x9OF4XFHGJHmJtlfZOLrug1BOa2q/tqmFS+b
oV8wyNfmmVeOn+FkJzyXEG+ThFpJkK5QYUvYBWB7FJSuH5skU7tyoXNdnmsac94A
elCIPw58O52P54uwuu3xHTdV6gnlmx0sv8HLc41gKeQYxX2+T9YY2gv1FK1Z9N+j
nqLW/f+m1/GNpY+Fxjhb6yOPf1FlHr8UxjWzI+RbYksfo8E0pgThqPW1VnBxLoHl
MS5aSLujOv/OoIGc/R+rbEbnohlzMyTBM0iNtvQSifLG+Gkux5ZSCEZeu2M9+SC9
qRr02Cb/zE0PsVGK13tE8fvjg7/KVuU8EINlIGUu+6s9NlEmCjkCnZGII6QWfsmv
R0BEw0xrtyxTsv+TXctTHatWFDlFCT74h3/bzENnq+ncaWZoLVOaeEAXepZHgRVv
/7oxB9ZdWa59ZeCIukDlcv3Xk9zDmWuMeZj150b8L5Na3mUvMTr644lOgQg2GYz5
1vZKTZa2pJ8XiDVmgBqwLRBckuo/PM/Ue8ddx4+R0f2t5LgbyBuzYiuqx1qhqUeD
2BsS4XM2wRmttSLzcOsy6wDJdfGLnv+LDwQ+ABT86igcpdTzGBydWWXarXwZG/4W
vJy6jvJcBEJtSJ29ZnGYxpvo5mOJYkfalZmmHhZaw/2AuYTNMQGlHba47nkBKddN
7MP7mMnl7Wvoi3OXbAr6gE7aYD2wd7S7d2YcyAMIptrIILLdrdKYfRSy51FXqC33
bZC7QIRTrygRh15UM+zxd1BosfWmGz070AoV6qOJURRzLPRufnHJSCQtUPWgY40V
F3jCy+SSgXPo9bUPSg0ty4uIEaVEfY39DcTxdIehvPiY5ld6SAd7bquzxdiVeOrC
klqSxm5ko/y6owF5qsTp9B0SC3Z++1+cO00W8ZVnymtq6goGLh6KrYuq5Mtf61Vf
Yt5mZkPyD3ljnWNjEhaQCZYhuBw1kmS1Uo6HcqCfaJe42InRmEtIITNb6zPDeQum
aituip0XyRZM8HWJddkONx9hk5AI07+/LtKm0qVdmrlpo0SgRa6/4T71dT1V3Ds2
kMzTvn/H1K/DTGFZKDUTGU8s9EFLG8h726nlJVkhXCNGKVAH2UXeEJSmAYSXBboA
/cAm7zp2+EGhNrNaEnTvLxyiOe8h03ZLPNBjF/oDqiWjcEa5bSEEH/60vPPWwdkf
tXFXgUx9x/HrSeoayJ2Q5zCiJXrrEmSiAfspLpD9iXrRY+NDvGTs5Btrk5IZKszE
Vj9B4Eww+Y7MLk25OfLB+Po8B9KKvSp6PdR1lgnbM3gSH4Sggv/igg1+E5sE4tFN
RfjawZts+u6+hDyQyf3Q3QjhWo//iCfzvBxo2cel/VuvwjkGKHQ01MV0JJ69MliR
yKQGoRZm043WvaAtsM8ADIEuXQWfaZzuMqEas8o+AWgPFwJtyuuteOo45/SwZt7J
dr8yuh374mMhz40dHH8uz3gBkc89feV9ZbmIw72QvE8CRj/DV+IK10WUzezh6sRF
61bZEs6KHSj6J3lQiQYor6YepzPLYWmPdzPBCQgmkHFf2c5uB/fx/G4jM2D0Kv+d
ZN4F8NVxuMaxR+AyjPV8ldpPbb8JCy0Eizc583bqmwXtleEgj5u6+4Hpc8zs2wFH
0MwpNS8TuLWmLKS5uobB6ejPuUY/ffzP30GR6vaVwRAcxmEebdaSWmN9B9L9vFme
FXAqEWnDQKbzWpiBAFjBpfhnG+dprYdGARdrHlXljMO7NQy5iqtzZ9iMIcw2Ixcx
UtA9QN4AMt/1pED8TrlfuP4si4ZT0bioDmsvHEK0kKfKdq8KC1y4M37PTk451w5D
wOtjlJ8vXntpJqOVFvi9gTZ/eG8ozzMRZWpSOSvDl4w6h5Ifh68mHspmbmhH4ECb
H0dpFRqlXkp50oOvfu4ljBzkAaJngcGKeeRU4K+PR3IOzUPSzl7IqwBhq3pgDg67
SfUV+32U3q34yyjy+It7Ct/C4HoQvjCdEqxtJ+6DNfFYh431Nm4RgvuhH8dwrp56
YQfYsuCSu08k/yMiMvCF4+7obZsbkMq7bPr/KFDqKLONVf2g3LNwoIl6WRxB4S56
cN+AIap8H/4f9miNq0v5/aCOb/SPLWZJ6050XnOG+sl4kJWx7zO0kWgN6WHmZx6m
bmEK96ANsQbZ4qx1cZoYZznH0UGWDvZilVtgbMKFIP8nhFHzY1xHCqDB+u1UHzrj
PZe/z8qYTip084OIJdVFemdH8YiRous1XiAig8yJVubBP+YSm7BwZxiBiPi64aDA
DMWsbEaM7MdlV12hWoGcDA5RLWTjOHU/YoKS1tX9QW0nnUddzVdv4I0myWfE5OQY
+o74H+kPLRZUNFjablF99W3OalnvSg5ejLec1BhtZ7LimseVo09pPIp6bKJ4PM35
+7Yb2TFhqcDrL3xl/EsELTp+iZjQkMUBQxF26Ke8HPzv6QYXn2IYdvEIfXrkNTpG
TFFGUavtToOa+T1mTjry8OW9whFaVLds/FWCCda1feL6niTP+8K0pB76bKGHGTjJ
OP1+P+2bu0BSNeoFafFzFNHbLcEOLnpPEHsFNLrdPSegekJYoH1hxHoTVnJvMQNm
hxz+Ov54z0wKHPp9KEFpm9bb9qJ+B0XMqrHG8dgq9R+9ExXJ7b91AFvDh02R9xl7
Ae01xgCeHAmhukfVpx/lrZ4OgSqOpAFktVxlcbnGsUPm9DmI0slxqAF5K8PBr/cX
7E6Odn+A+MUn+l54VF+aAETmZ4PU/NaM8BESUYLVMrxmItiDqMjnycYfPh5DPfqv
ySAiBKp1fiEeehAlqrnSHUJyf9DULa+o8UyS/rfz5p4iAixsGnXdzxhQ9nmAPDcD
7nIHc4hNx+jU3wLurYvIK4V0AzElgxBc54fJ+2TBm0vvg1WWwuX2WhSnXmQq7yHA
j6u3ssTFWMZ9LnFxUrcA1LRxPayiZ6+tI6nrOaL/GGJZP5FDQgzbtA6469lZ0xF8
m45ozWizFGLl7CIQy14PaBjlj/0ITkib6k7ltyCPln/eKahrisiWFBZJMqJD6hiO
/o3afPP1VZJP29PSODJ1VeoKxVqJNlvPVBwFYyGxPuN33U8e1B1XONbBBrHj2YS2
NiTiV8XwRQQGqdlodwbYrZxkiUP3bEki+x6DmmvrK15gXe2qJvCrfM3SS+SgWcmJ
tRk+iNH0e7bMR8IexNdkpxyaAThl45Z9aeWGM5DiXorjc+5S4b3Nua8wyHqdBeJg
Yz/DfzknEnFg0wC7OoEd8ABm4nNauZ7EBLj13SNYA+9LTmNP+fFV1Ra/w2SKpuB1
TLrid7Ep6n/y9Q7Z+pXlmmxSY4AeEi35Yyqto3NVIN+9DeIfyH/QgxFmpMOkVjSZ
i8KipidxTXoE6ZEIEHzEm+x1TExBbzpHaGUQPT6LcATpwsnG7OKobKXvgivP9B3f
JMuKNxuwOFtroqf3d34n1R78o4UlMKTdoGP41cKGbFE6zjO0q+6ZfunIfZtqIVTs
sdpPvbxgbQ2tLgDDCpUc4vSDehh8iYTSyBr6stJm/zSuS6EitiHuz2BhknUyCLA9
UFcWv06B7MWI6I3aaGp36q14ZfYLRZq4XdJ0Yvsc5rDgUlH4w+PsNq3P5AVBaksE
Qh1+yHJTeqeaCXVbNemIDLVswSoeWRgRwgdWrpLIcl67dDkgQTUryEfJRJ8rmZLy
uGY9rIECbm+f2K6BuczexKrqDKwQTwJx7ZxKXvMBX+lxlOY5PMA0U45VD85ekeCR
8LSR+7Ece3BWEm7v2h+DBBtWmWUkQ5O0/0mbniAjKihnPCpNRIdp1WUhsMaEFpMj
vBAuXDG3rOozdrGbzHDukg5f5GU7/aBTklBJRutmdG09rooQCwKF93/qZ5G5RWxk
JH0p+9RrbYp+LmPr+2ED6MA9FyNxnnpdh/P2RJxV0wT0CWo74HSPnmQy8/j5ItmK
va7nNnL8mkjGoUIoLgVvERpKRup7G9ax5DxtCcwrvRxbr1QHDwA0QGX2rVAAgz0I
bWcRqbupBkm3eB+WcTwVoXXljLGB8/WuqSqnIPtr50wcWjS5Gidyu+faOM9w6KtI
DUdJUuZzjUhnwVwrlJFBlTefnUu8XiTm3iw04Bh40yVYeQedL6f1gLvErdKM3Djd
BbPksaUHDz7XjNZnj+4P2x3B0tMbiyB6s9KJZav7zWYSdOvbhC7cl71JL4HEucmc
1wyUa0GPunh3cdiY6Nw4u2MXtEeztTd5qJX+qTu7vUUNJNX08l9pmzu2TFSO7yhA
EqR1QerSZvlHuyut8o3Xr0Nwbwa7vKKkfN442snAy8SJ4wH/cTF52UrpksLeOWoY
FaLp83eCAgJolD+8XdZ+mNEvDvirXi/tj21g4lwic5v5an5tuRyzYXnGYetN2aK7
7wSLhIRs2PLQUS+Fh4qPBoPVZ/TBj3oP8LBb7up3u7qNmyghR2FrlD6WgxSOvSlR
UAJeWJtsqjfxO1bQqDSWcRFp8uTB/7ITZw/BVNVA8gLXhPcmdUFjj68NHERBQd2T
xLGMcfnGff46EIArJ9Sq1iIftJ5+eyMnbVVKapvdx3DV6pkXgv2b1xd5YN0AVYx8
z79JzWS0Pc8x38QyXDLSlkj2OoHomwlfxojtXLJWAum+OdpM2XX5zzWhw86fUv0+
wX1F5sHti5976hRNsuuZ/xNTouSznW47ZuTOkbT5BK/JPLc4YYYdUZTqPi0FumBS
EMaRmuiPOnCQgEP76FBanB3AkAXi7p5n/hnTPtpNW+CIhB5E24sBdi8QpbzAMT8p
Tfx+Jh2FMk8BLcRmXe62U1lZdfslDEa/6mPh4bO/4CD9tlH8sQiuxfFlnOloqb3O
UsPY3wzWtrBW0IJR6+c7Z5cN444K7t909SNHuVp/TzpFQ2GFPcqpYFy/2CFsvEMZ
3B0toPNCIYjdCi66C0LHyf9z7hrvmkttDcfGMNbly6SAHTrX/2GkrkXkCnC1AtQR
/Q7TYYGIlJZXDjEhbx8nn55rKXzgKYCIuTTr51PuUrUQGHpzkwKAiTojyMTupvdK
av3OZAuF7jo48ZN5p7xgX456xVM9HU+MtZSoZ/GX32B2/pZOLwLHzjoehQ8NP/K1
Uop6I+QXfw+kYfseYRDFfWaprTJUhuwon6cZH0mvsHMLA6kjnBjFPykArWS1ukEc
g7QAA/Gu4fRQ/vY14QrAhNx4rrmb+vNmbm97mW/yWuQw9qlNBkHVawu2OdzekoBD
sj3f0o5GHzKj8k400e1BZPSMHv5vqyg6Et6Lskvxyree26BUiL9JJ80eHbh3Dez2
NpiOTpZxkmmjlLDMRT1n0i+O0d6EVBTJIhYG3aa0yFg/JdCA0v7sWYfJN+NI+UKq
LoxJXoi+Wo5LXI/o27f1T6uCP5RqfEG4hDAcS8gJGqxCT9yV4KiquaR6oPnOrYAo
gDpZY3FVyhQomIPqPmOCPAOc5/BDeYDBIYxkm/+4mXDs4rwYxu1TCwvmXGQ5fxFC
IW4Lkt8n0F19qf7ExYbYPuUysCrn/HMOOwoUpcsQFX6dPUf4SATJzfEpULeU0DHU
rK5owfgCLc1HHzf1UIK8RBpYMsnN3tQFiaBTHkgArSbmc7GFNV1U372wOLJt448u
63WiY1gotSU805TyutU8P6l/PZEdcVmAoGdoC9zyh6BPCrfkzXSKa9y7/81yLWrD
BPH+3IK5bMqforg+07lYABgRYcyFMNNwNYkDIcwiEjEKWJM6E+cBaV5mHDpA9y82
O9s5q5SPcT62R3MV+VMXifwfdDkmd58RAKXskUCg/eF3LRYiodvogTLpm0YSkmN7
2AnPCG21BMn3DlQ+JQ+eodv0puxWL1q+AfznIl7tVucyxXBs3kqBAxYYzontHCQQ
h1u+EiucKWQDZtEEmqsWjdngQlOcc8PkydHjobAhBMo86LYAMiYAnVep08KOqM1J
tImRBnOAhDGMKRrEVRaDpU10y8VBg4YrrtWxGIQrIev1GX8iDY28L2PzeKYW2TEW
VRkv7Wb9YLPm08FvtpSYMaJWToyKHnrLqewCGw06HUUkkMx8/nyW9cmCUaQ376dG
Dz6sFYktcXjjwbpR6rkasfWRCotIsofo92ZiwIBx+lEDFvnoZT3TR+ZDFaq7eG3/
xQDbZp4htSs3X9ceolOMdVF/gkNQ4RYjtvjJVfi/mLDn0PCHr2aBNl6QLGWlgEnT
VIM59l28KUcHOF9O7DSdnsyqQ74LDvI3+sDVkGHGqwOLPhiHj23UCRCaOXjiH4e7
EncaaLaFKdE8VTnAz2cTgOH3m/+de0hPpEC9ISngSDD2bR5uAjtehU2CkYcgH1O+
mLN0cheLOZoj3r4B9nyxgIuPMbKA9KV7IUBHMeprGDEWUYtMMtEaH42vF0m80JrM
JTXfYEyRuxSiLZL+buDmbonI7wJAoVSDyEyYaFKeEMpwhlwLnEOwK/FSeHTvPEEW
K2cjzhed4kOzsPxRqnGp/zWq8bPW1QMvKh8ZihDl9d5/DJ17+FQNmKDy/5mpfXEp
wdlk26HasOH2C0thvSsW2eWTlhzYCMeYxKkyFzot7ZW+ZNBLxYLt64PPLgL0awTE
H77YLn4B0AOvjMJwa09Ol2QDBQWEVKe8ibvLZxfL0smrhKq4odpT0YpRWkqyHRI8
dt6v9r98VIYzu+CWI4qV4yBUgx/RI9EWfleBAv5PO80lJX9U9xMFA10N4rfWiD3D
sPM2BsUw/bDJaYmqp9DgeNuiyLxeWc6GC1+6MjiO4j09RD7Znlvk2fFABaLHwfp6
L/vwacjBUn9Zu6ZeIeFtgT9a0ZYgStFoV5dQ7SkX4DOXQcREyYDo5R1lpfB/GtxJ
A0632wVlbC+KLSWvLPOawK1OrhgOZsSHEP2mpWmLNwqdQRxAjHPCJmkpOwh2/KuG
AeWAvqbAZQZ9KZe7h11qIxh94jXRg8CxnXsGWKvSbOmAyo+fmZnuWIhgtowk9rBt
DCdflOx7piaypCPWtjazRIVcBSDBvj8kvdkMBNUmS23C45j8ShCOWnoxWekHmbiw
QaHLx0Cgk6mhHM39kE1LA5JRp4dz5QO2ZNwaVna/zXuJcurNf5hGCTgCthPu2Vu8
kcf0zP/quzO5azfyg/IiFasVWck5/FVE3N+Gtiu9fYLvBGaKqRSRk++hT54S0I5Q
L5HoKcM3ZS1P7uz07s8m9ZJVrsumXwAmOXE8R0xfGcdg124Sww4l7jYrYbWY+QT7
YF37vNqyxgDFBUpcZ3wjofzbl2S1ZohK/OkkWlN/zfSJWfhe4gcjAoQxq2R/VpPa
W06jXuCdtkyfBpUU+EViQolTLOSojVTfCsnXDBLE6gzYZ/DQ+HIlzjB/DI0zbHA3
p5vrQZ9vj/VS0NngTvP3Lg==
`protect END_PROTECTED
