`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QaLpNlLF5rBWOn8Nfu52hrqlX/h2F2Yli4sbK+ItEig4wxdp0O68LjMlnV5+dxxD
a/r87pE0Cpxtc38pWCPy5+hFYpRH2VI+NhfMnGGljelnkjlZff9VuB0DkfInIsq5
SjFHTO24uQIVCkpHQFH6xndARi5rcJDIkAcEW8d0fZnFWVvBcwL/8sx63kpKD7cV
1rOIF6IQOA8bfA1FNDnnibdSASWlJ0qQlkzXSdk3A5CZzHYRIo/MRbupi8V4p/PT
NotSz0BinYQXB4ZU+qdJuj4OaUmUboIYayBR+OeH00w9dklwxCoe165/AdSqBud8
40fkG26PQG4otBUGvEaxQWQbDFHHFfRiUsZRuzv+GFguW+YPZ3ye2e4EfQXTMbBM
`protect END_PROTECTED
