`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1QVdIMCSmq8oLzixwYJmjKf2BPmLWQnuWB+w+MhdcW7NlANZnLJST9xHrYjW6tI2
TJLVzLHFHh9VRTonhHs13r9mBXW3kHVRLzxGn6FSbC8u5ahQIH0kXCm0qgdFtKtX
VwnWoPjg1YDsKhOrttauSbpkKXStK0uTwKS+qVdN3uE1Ysl5LX06oo219Dn1c7d9
JhFSoKtY/S00TvEavD6E70bgrPanDVznJG2ppQpV1/JJo1xMeJNftaRsCnnibZ2X
zLI8qYicH9stn4xA5qoG292EoL5j2NwfhxEcGTsRolVDMwXwhBFoIlCgN161bjtL
nMLHTeY1lw4xGifRe4nBEq0lBdWI37avRj2i/tSgA2A6QI92eF2iK95UjB/KmHxx
IMTmdkpepQi2EEMBhLfczuEboeonqqa/QFsBlfXRHTYJqBeJ+GFs1PIH5LlsJta5
zv5XYF5iV8603p8dDdHtUx7Et3j0rh1lY1JHSLXBLXf8/HgB6O0tHtUnxH6CLU1t
xQX8LfEUqMxvrtEDB8Gd+Mh5UrU0DrmycwQsaZih+flW8x9JngZnyK+/WRkqixht
72ecAqVjOvmeymu+IGCIWenswgsp9z7ih4movvoIvscDguz80D6qFtG2ZY2LDKT7
3YOA4MZsMCqgXwpkHVHpbbpD6s6py5yESyvJt8jyfHBr/GdyTRInmetyCMe5dzR1
AfajB5TF9btMlZaAD19UaSXm9sJU+CZwkzkYWedGghBmpBtJohKZoY0o+fgrbvx5
gctK33LmPRzosNYV7RbSEVDaXxCkvj9Ip7OZbKMFzoVFBkIB4cTUGOFNGBdDRWLY
KaQBN3tPwjOv88Zoqen25US4r4F0Pxmx7EwNgqiunCOW1JWOwDrTFLaw6ZtAq8lP
QMjjsxGUlA4NQ8CiavIevH7fw/CSMYNs61tizXrCtL8FwIUrdh6zCmVEJ1prBTVV
S09E3nUuUm4xr3DQrC0dW1O+uXZHCjfEkoZuccU3U3re9TJG+RyhRn9kwLkQBmv1
1mo3FuiPNidVaedeU29Er7H3/BkYJJXYtw93Vl7lo2DB6m+kaUAQcKmHrCL8+HBh
7cS68zBEC0aaMhsQKVu0dAV5nM6HFLvQRCFuufZbbd0oQq12PRP7/xSl8Rp84sEw
TLfvKHzTZRq4sYUo2kns301drZcmI06E6Y8fMRbVXIk=
`protect END_PROTECTED
