`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QnrpQc+0ljSrEmuTqtGEs0d9Zwnf1evCP99KmbITCKMco2r7uSR3bJUThu+EVlnm
/dS/62S03gGd5sTacROCxeALbPfABcBwTeQ7sCRN6bisyfhBCIDy7X9cP9fLegCc
2NVZl0ucazBqVLoUlkWZ8F7l26WllI69FKO75HLuQ2LTZQXn1pdIDxnFUzJbAF/t
qddtO8+ftkNzlZ2wIPnzfs2ZvuOkyl6Pr1DYRwWPVX1TKoHqpqNIklxVg0hwmXHb
BBnyALHSMAza2GQ+bdPfisLuZ3gJbFtDfa8a/WDNEB353Wxueow/bF0iU3XaIXrb
Sg2blu1QQX+c78A7vjbf9g==
`protect END_PROTECTED
