`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Avyd6Fv3Y1msqTKRnJWO41fi1WkHji/K2FbfNFJbjyvHQJZ7DmLdYb4lGE0z4Rlj
n+kp3/nnRiu5//Smt4b4yfrFQeQK5LGJYTh1kDF3KFSE8Sm6pc3tb2gDphssP0h2
GSnLQueyVfTpH/V+V1+wT4HDKQGSo9lWCwjIpuYpA71DDgZQa+KZM96NQILuOS95
BiF6CG3cCsIQj5A7CwjVl469tvUkGlqyxAOqXDbL7JwvArNYyTZntIPdlJw1yitQ
pMlz7EW+jUBD3ATZcZf+1hcFuP7zF8/sG1Ycabe3LzD2UpQ/FRZ5A7lzwk2UT+2E
OVuJrCFW6qXSL2yXTvHAI0AugRQLpecO/OgBl+hi3GTYv47w4EP1wsBGm8xDu3iH
SHHEio5zjiD9dw181oy+BseOxJjY4G6aQ9bjbbrQ0ds=
`protect END_PROTECTED
