`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6vyAD/zXM6DXdwhDbVe/AiECGlVjEIh9BPwTp1Y1chURUXfBhkxj/k0twI+ID/N
n/LwvtBHfm2UwqTZ4BnvE1j0nqTQ4op6phZsUK+s+ozuyL8vez5GVRsYohtC3b7M
7V/+hpFO+5TRuu58PUzfgt+Tz9hA1bxBauw7i0O/eM8eh8Ll7GKpJdO+7LY1KUPW
4MeEbDall1G6156mhKzXJrfCRcUQoFN8FFglgFfR8SJuu0qZQxUlfThBgFxED3VZ
jVfWJ2xYy76znfP/2IVop8pdTblvNKHrk5C8hM68CAZtrl14KsHc6BH0o4N3FDfy
BYL9LOk8vUurm40EBPasbZ8d3RGCNseZVeuL2SB4o0CxEcEJpRg2mIBNt8oQsCBb
ATWao4+WErfJHpBSGidEMWRMBieYgIaZh+BvupBVS+PwFBYHCZ3PTi+JXO6Bi48e
i+LGyEsGJNov7ugTOgP+QLd1JgiYOj7fjBYsZ1gQPIw=
`protect END_PROTECTED
