`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/PBnmUMxF41qhY/psvP+bDxBdY5+6vBp0OUa0k/ES2IrnQwByRoT9ei0kzMwp2mE
262dc4eGb9rhlxYSaf6G/JbXxi4jX/LOFeOkxmk5M35f/RVae8BpnJ4N0sht73km
CyCKnGsVm9arSK/ZtIy+OEKeS1e7jaVge6z49Cv+BMqvWqFAQXirGlyZ2DiE9Jxo
cq0Ra6obeu8FcmGZC+LfaQ+5MrxRK0mIYEQRuacdnY6vQkLCVC1nspVq9C0rv7JE
WPYzKB9taCenQdsMr7NUTU++34LxTyVuTCSnY2f2ghQYVhWuPGK2JZKRQy4fpNvl
URSzG+SPIciRI/okL1GykQ==
`protect END_PROTECTED
