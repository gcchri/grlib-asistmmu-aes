`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E0ES7sskGv3HBlVGuB+qJdsa3oKfGPNNq23yfvQlZ0MRfuhohk9PDhMukgp7C9z5
Yn6ha/seUwG8/WQVw7kvzcVAWbog1Ykq3Qm1Far4/0wcUYhiJgQVn7b1bp9ATReg
16E1fqsOcNrNlUmNJRxtwnYAMeQ4D1FTGn4dFN2zHYCh25A1Vgt1sPFx7ssTaBt/
YaQ6EkORjt+prc27O72khqXj5hvUxxlaK2ZwlITgLma5+n9eCdCSPIU+oKBDAAWs
R22FGrmcGJCwh0h2pcqqHCybT5CQoXw20Kpm4vFJrLTLudjMV/EdLgkTrgrdXoat
xnjnrh445scmHYK9ygteWozn7TRXFtTcjD8fcrFOc/lsyKhcuWGcalDixi+94GR2
M5eQtZnDgTzB+I37tZaakrS85gotNkoYZFsWpajZIJ8BOtaF2jxE6rYEJgRc+KJZ
s7NotC9ihM4iaxMKo+ycyBPztIRcXAHEc4ITo7Jp76yp1PdhELv+UyiEf84q3qsO
`protect END_PROTECTED
