`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uaPY5Kf3LKYMVqubiGFbj5BTJl4DDJkQmL5gfVCFxh7IUeQSR/+vEfZ0kyU3mAL9
EijvYiBMIABAsHaG4/TEFub8uBo2Ov6z1AQPEcfObE0Omv5kPLpcCVi8ASIu9z1z
O+6kJqfnuU6G2IMlHjpNAI/fAyn5oxGCLgrVONaasWVKE9YvexSakX/vEmxlo9r/
hhy/+QSpvVrgdMFuqSjRt0ceXXMy2hr/Z3dznrnSkz6Wy/qYGa0iea9jSSgs483F
9xtAIM0v9DddCDVKKvyQiyYzgWP6cQbtVZL/X4to/pwDthj/A0IUSbhCU9RNe+D8
eUroD7Iqr9xP0Jo9oy/UY+zejZxtW6eGO8DSgp10t9b8fKasp2uifJh2sC4/zafz
wmETsH/p50qepHeUltQ+zg==
`protect END_PROTECTED
