`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2q8qfuGf53ccvYodx9XQq5ERxu0Yobc69UlkB5TlWc2oJycbtqWKLnRDB6uvvg9r
E3G2j/fTud7JphNikHQCkFY44PXNwiLine1uuHSYrEPVo3ubQhrNjKE0aeKie/Qr
dKCbshsE9EFjfi22bI8Wv60I78P3cV/oSx+pJTmvz5RZFV9/bhCVpKbANPhyqJ1H
8x9CY+qX952yYZQPhhfPx92WPljvMt3/0A+R4wle1kx4MAQFx35KIm/MWxnMr2Qy
ckcfGkt19/+lXi1wHkEeO7xznr8fD2VYyl+g0qOPmy2jqTraa42bE9qU+UdWpxwR
xCwYCl0wAZdqJXQsqbrAG8ZPnexGrcjExgAL0sklUw4cBQCcf1p7NVYufKjGX3au
Q5jp/2m1dPbg3afJgYoyy6QQKdft4Mh7RDJkhtmv3+Jqr9XFFtgHgmi+Hf5sE3lR
H5erHD61eTYC/fPPRIj1gk6zH9Uc5IYtew8xIO++PEQPkj4MvSjPdgBloWyRRGLr
OszWEZz3sd2MTD2Js/06/8jCa6au09ilZr7aiUi7vT9RTiQrhItGTEVew9EMqVCz
IfSLv/13v/D+grEbgdVhf9hRN9oZuPyOALsuysJYMmp8Ija7Y8YbHqT3/EhW1TVK
gBWwB4CipvvNRJLdAElx8oJyA8yb42+ebKrk9ePZVZWSJNoWoQoKK+qs4KFeSqJ0
RZBhdFoyxKT1MwMWO09V2TxPXsLzYS3JkmIdvKlQjpR+BNrMjQ+o7Oadfun9MjxJ
rNh4zBn6hhKU90fUkJEd6ZOthiD/nRSZkWeWfMz3wktehplyrXCIs3TnlHedAYFi
V7Cp+Gqfioi8CGycE/2F7xEugTHvYSIvusI+FN8z7DPAGPvSNsqJCEBnTaIodTHf
Er68Xgg5jt/uOVW55pTprA==
`protect END_PROTECTED
