`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SfErtSN2EUtywSikf5H+Gh3K6Z8w2aFNtsPgbtDmJFWBmcUrGrflxtUCncQuKwfe
GQrclCocBB8NKn87mFW1pLF0c81Rrsn97Wxdp2IzAm9sW2YYV9LbdnSCe+2jPrqv
oJD7Lkh2CZ5NJzBQ4M+0vvwL5/Tky+C7+jy7WVT0gUPwfS5PLSvQEcDYk78fThji
InNeBOvm4tgeWy/kPsijUV/8WHEKl984i0Db+P4sQJkL63Zk4lGoWCVrBhUWnyaL
frZ61BC21imsHqm3JBinV80AnCRWqJrRyMU3vTAJno3HEKZJ+G2aLOcgfEqrN2yJ
VTuhaLHkmnXx45a0gdsAaet5VJiyU+Mz7AQFXUorjgtqloQiHSerpIGfpc4/z7PX
62O6O9ICgQ2N9BcpXF449lnxafw703DqgszTV7g7HKh65uxvdnW1lPGIAJwXsL58
acBQqYe86nHlEpFo8lpejXokAVj4P3sLbMv1HV0sbik59lYUqTL9doTv+EdG7n7J
`protect END_PROTECTED
