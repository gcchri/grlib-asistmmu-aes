`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WFPH6w9+0rn+3o5deA6tnK2TmJ81IhgnfkkbSjU2/zBCuX2rFfkbSvfiq1EPsnnd
9+/KrrOii1L6PC8mr8FwViL2yGRtHG3RlnTBXNqjnYGOYY23j5O0q1uuIWzfCjy2
sw82Ht9iDxHBm2r6g7MdOqbiueaAi1YHoiIoAveMSWWMRfC7SF51Tflwud3Fa7of
dsIXbt4kDvDwWnOXgeMLM9SOsTEyfhxlE94rVxfHATN5I+DdqbtDpZlT4WlRUDPP
`protect END_PROTECTED
