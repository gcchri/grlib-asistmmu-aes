`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EGrYMrSPogtXuNTYIjJcEzlIjUfqC/TGkO2pku4H1OvVQUYByxdEcHOAMzqcUNIi
I1jYpf6kfsmnSbB42p2KM8BXbLiu8O7FiO/fXZgLNtTwC3a0YcvUc2iD8cdHEMH+
+7aDIKU4JNgSFSXdaIBtGTfALlYVny7edMou2gTRdIuHvKKC/RGDlFvJQVBLh2OU
/cDkPwAjr2CndYWkI29xg+Y5cEMwYEHe8syCm7mOA1HR8X9jGt2NMkqmWRHR9qee
Da6ZMpSmA/pnI/N0ZiebXiFInTofZd6b3n03iAqBzxYExMxBAnuGU3wbdZNOQDU9
UAQmC8NoMCV5rTWpWmXJpi/gaSl92ulWbZj9uRhqywzt/1ar7Q8JN7CR6eW6Ax2y
XwkaIsLJxHsN4zjRbhw/FHsgE/dR1cDhz5EzWUwZ28UCbgROlTcFxfDov30OUoYn
NXBG+wFfB6BBwjTMO8GLkMlLzHXCiklZeAtTzYf1VGRKnGdJrAwEq+/SCK8JFdzx
OozkIO3cDpWu40HN+jNba+TFzF/Lt/hz24PEZnW2lUx0xYwEqAZroSIiZwst4/ce
FTznAWEEC7LWBpAfwqhdNPuu/KXy6A4xNUQL3Mc7C+ixKD717tZUZe85OfMdPzyK
2fOJNI5vqNSZeVf1uADDH+28ADx5lAD0pKLRo5YmEm1OsJSJvUqCce+BaSFXaL67
uLJc1mzEUXwNiijq0EVdoWvAXvfzsaQ7Lvbw22foqvbz0btNVhmVWwiAiWj4jTUR
7dYEP7SX8kTua5dXAyNF90Iw+6ExjuQnmv/FnPyWKWzAMNeLMOKKfk9slc8ebcCG
E7eCPVmcDV4nUhsul0VoO4xt0g/H7DJn3Wc/t3qWdtniC/E4xcmuIg30I+cKyl+H
Ua6/yGqGbZMd9Fnqai5yWBzJRg0BVcRgLum6FingmtCL8e+6LXa9pUzdJtSIVvrV
1bZYFMBwHMwKzGfvX9GXYjm2sX24I1iWwpCl2Vl5VNgMYMYOjGTAonKiTjcwTYLY
zSrxmTVJTJE+OD2Jv4Bb2T9NI7IYL7RYxVhtvU00SBz/DCvawcY4+xK2fKcI5rIF
bphXMqD0LBuzopEE/DwBQUsuWc2cwdIyeOWEuYTR1XqKwxhluoz8zPjToJ8bPVwy
sH/fur7mzAKRno6BnOr/I9R3OaWhUOqOYKVp51Jk63yyXBVaKpQL6GF59om8LUxi
WUSI0RhvOP6u7MkwDUisCuKhhgcXz+5yd0ry7vEEwx29sdUazJ08FRSi36DONrDd
5IpVkI566CW6kyJ5tluXmaX8LEYD5E8Y2jTJ10mY+XJvReOZO+IDW+4MrFElDq9e
wdq722yZ0u6ogce8JklGq7suN/NqYEQa6nATbOw4NjPBAe1QGdDyZ9m140BVDtye
vvYQtPXZ3pmOXDFniz6NeQJxLUmEqXNZrt438nRQVWaqVCglNHr0FU9pViPrbyRd
VcmwTeZZzer6JiNuF7a3C+kvZaXhHjD4SMeBW29XG2sYd3WBc3I1yO8CTJyE3wmh
RRI09gn0zhuvmkSZPPGEf9AX1aQhOjnOKVYg46ORurdwgYnTgqGiJSPI5VoUC+V7
O0Sem8wwhw06G/EeG+qRZ5D/e7x0H9ZYgg4Ktm3B9HB2tvDpyBTK3GOGV3XI+RsX
cBQspmnF8XvPk8jjjAAJWCWxrkyETwOAQX97YLuDQFkwL86WftNmV+JYSw5emJZI
5GkJ5l3oKHFAGjTdq8SwMHzqHrZ7Z/BGp39X0XleVP5stUAlKx1oqbEzEcz1n/5E
2wa8mHZSkdTNfAz2X96ogosIgkDsebItbQA6tqwlrAD3rRqjylFJc7FdcBzND7YK
EEVRUkOoR7qqT9wbQjHvzbmRGUOIA9uN5ViO07EZ5Hou2ifIkRkBbdGW84z6UuL0
XUKFbudWiQTMnt7YRbJomReW57qwbatrDqauaaDWzSI1v+VF2uQImGoXcTOK2YE1
YPKSAV/r+vxQDUO/ngxTWlcoUwwG9hGwHqMNwlAqBxliT6FmFBT5fLhAqNMjcQY3
zs/Gq/G+hho58Fa71jIRux2+jwCpAB6+UTH+TSO/SWzXlNL0Qk0uCNL0xtppOhMz
`protect END_PROTECTED
