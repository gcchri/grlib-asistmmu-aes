`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ll7f4LeAt9IjgcSCUaVvZeOzUq1Wh0/JIxYSPtqXuhQ8oSP2Rpkx/GRl4jm3hvjY
mT+6DPPT6DtVpKx/aLMBzeSItN/6hEc68WLJxQ8RgKEX19jDjyn/NY79lmDQ/JCn
WLHogcSB2xOAGl3NFqnWOHHsibAAP6zUPFo90XqDCRJNqRxgHPpcuSVCnYfNHuqv
WxDau3CCtZySvN6FoiqBsiZN1wREy+mU7lhsZQSs/MvxVBop3sKCf2wZaQ1osztw
98XRgXxkzR4JVBMthxzfaUUFwb4MUeuc6iiYCxNuRQ36ciQ5YGl3OUTRbUH1oh60
Hjx4T8V3fwcpm+S6zWMiTu0wUeib8QdohKFzLCDd+5nZ4NP1TFz1aWk0GqzJ7pbm
fLK0fZ5KSokOlb+C7fxbPoWSwXQYtR3pj1fz1CF9y2L+s9H/P6XlJZVcKE8OvL6M
05NiEUs/6nP6OTtobESwnfpBgPHAoFxyVtNV6InfPgyM9AdAzPTKOBB21qguCvsO
YuflI0ubvQPDZp2Wq27WDFDdb6OmurMrylkfqzTHkkSCcyst+Cs0a8Bg7H1SqTYO
tCb0pEPQyv3a41UlCS9xE0kdOqaoAUi+zusSKvc54LkDZ4WCV5LFCOPJMCd2hbUX
urI7/2GjD3WWfoAr0IOBdG/j7cQLbQmfxMvHUxA3ZgY=
`protect END_PROTECTED
