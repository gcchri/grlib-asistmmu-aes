`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H7MW6RvAbLfMEfzwAC0kU2ucSLNB+O7zw3drAyRk/xNiWAOZZkZ1vw91THvuyNh6
xKpiVlFtXDrw7ST152AFrJVbtbAozZJA+yFJ/sBHKAm0PBjp7YBYSALqpJtOjQGx
NV9+2fh446TVm5yDATvILGOUoxzzM7t59OunyLG9CAmX3coNa+UBo7KR6kwpS+9E
3wYwP3V6gh9q9bH8s1yz75EzT7MtR1rKOPTMNBET24e4a+Vd9RHoXVPAbHfQ43oF
CjcnQYrXXfGV5JOxNbc04XFeFBTijMC4rEq1gOVdJszMO+U8zALusKh/dgjflLGf
YSjb4bfyfxe7rxbXwyEzgTABCCjSqfg8d0ATBXJaMQN0FvmsYh4aNU4v8t3CbW9F
hiPKS5h07Za9SbzMq5qq8COpzE/J9P7QpKMfiL5GS+RJIryugOWHk9yZjCS3Wgiz
h9plA+uU+V1xEy0ke7zlwwb6V6rdvlqcltG5wtlMq+yc0jXu0+/fWbBt7w6sHwqX
DGTNjHSVVUYQKztaX0G/I9UA6pc0MEroAeNBifqwXNNsem1RPaF+M1hrJn90a/e/
lSXFP0TzO64ibVzAyij4wVpNHsG23TvF9qgnnSsqhwGV1dIU0/u8Kaxf4nHSE2d2
GUSdRT/+BND2poYG5pkQ4fOVq7D780pFPI07MBTVImVVFsvLovvJ+y3mqsD1FLls
Omp//3oxmi2xj53GBQJ4cxwgjYOGNmjSZ4xSGWLJjvgI8ceoqozmzStapDDEQCo0
JwetxtS3JV91qW7DJNv06nmwwKYj7RQ2xQtdbK7qbHje0GPoerS6XHlipNxxjlRQ
2KO3EK1C4LMJC8QLJFS4LBFjcxfBf1TQdviVfa9xOgiTzD6RrFAjFFXL+hufQmml
7+4g+kIeEaCQhyLPKWPWW4JKZeBoGmtHccruvx7ekplmRRKrzf1mS/RK6M5zBQ3N
SLxivZHdO6TBeCO75tznuOUMltICbIotoDQpFs8M561jXQRTzpx+6X14wrJeFeqb
XNS2GiEuAGPpHy3lOo+aJCwuEdldQZsfqL4QmwRnBEry51MyxdgoWM+MOSRMD/LO
OK8ICY+W+DXW5LM3w21WFcxbgTdtpy022xccJanLYk/IDNf2muBj1QQRp1/0GmWM
gM0F0f2wmwX4D0EsAL8UaxHXKXpXTXu1RBU8nG/9LNgZPiZA50GEJq/+sipFyVLe
+q6icro1mrER19OjXPRr/H20Bq9EhUqYIhxEIKclit0D40xKYgfnDPTtPEh/Ssw+
nJuDLKDcOHTZFcESXRagvEbaNUg0BtzAXa5x9wYe57/e331hePvQnlSje85XrRfk
xGHxJLXfnOnJQ5g/RRC+lvrLBgJ0CXOb/+4VjACq6xajJ9YjgZw3HyHs88maggUc
WuD9rpeaaiVm9s574eNzFyk8mC6dExBFv31z2GhWRcJ1bFmVaIA5zsaO1tSPQFKR
m82gYAxeKjZxMVzC+SWdfGxl/As4CRso7JOQQB9lMxPF0+8aA69ZnDjbtv0xUUki
45amsTK7QFwguxRtLx+hQbOUqAhWPUvP8eGf3nMc05DXzKwslE9dfrY3y0FK+EK/
3+5QM348kooAC/TGllX3hvfHvQkL48f4mE05NeBK131ED1TW5e2I9llbhK4eFzw8
VZpqVDh9Fhuc0BZpybKRA3AAIeYDCTcFrkzosm6sRcPqyAZt+ZI8Xi4qPnWVJlkj
YQBh0AzLDjpD1KEMe+dVJxsi5hlxXVBtsDDjnr8uVC4/d3M9MYM3ujPcqqAZeeiy
4Wjd2F89GzhEE6UooILVDycX7LHcL8aHtFNLIWLoKPNt/Cnbi10hB9B/m8Zvi+ZS
gODQUheG//uoLjrBUUA/nWL+KpmWDgiN8pTjX5+fLUDtNAEQx6I32wvAfyebDrXL
syl0K1ytiAhlgVWT8QzzWRjs3qEXBM3Ky7PEA1h1de3lWPjYi3FaeoT4maFGpzob
LlfiNq7+DUMFMS/MvdssphHX287UTK4rZjmjlzmftdVZL29ZQMmylVPzK5c2sAhD
6ugB6rse6Xt36w4ZRmVrkKdfo2zfb4kNGe/vclOz1nLRxn9O3HTP8S8ddW3p3ZZE
LF4oyufnzl/0PimSgyYY/eZudHi1wnG9AdfauURuOQJw4GSUtMczal4ioR0ncIYK
U4/m73q/qYLdtGaqC47Kzw4yNgawOiwgk9SR8/liC8+SMQQbjXObMiTIHCzZ/u12
vWoXaiEMa2Wau7jfpb+PENCS9z8oL0Spoa1jhULrRE+fV1RYA99t/CyAbPt2xEXN
q6oJgVT40SW81i4MadbHC8ztwgJdytF0a2ZS8PLc3QtNDIrqfEDrpXvfEBXW/J8S
/RwGp7OD47risZe63cb9eo2UD8CPvIvzGFJtFuCymmYA0FX48QaU6xc8zLh8/Uos
/6Nk41zqc5zvDPAO3PrFZ+/KDsvIvn3OSCSUtW4O0Omk4s9/BuPTg7Oxy9xkePZR
y9BTM5tusA3WPCDM1VezsUmGrYO+fpIqQN5DqIgAfHyR6yCu6JX9FANnP4vteTNx
YRG5rlCgUHu4qL3DvNrGKKrMvSwrZ+cC15seaxrREAp//keAn5nMKzV651hXBXEN
U94CjrZD/dHvQ9XaRD4XGpKURn/qYx6eDJQXdxvY2KAgOIxgS873ykVRRO/2XYrb
TfyfaZxlxhCXP4fyWBf5Q4/zcZMtAxnNS1++eIKzvzLIuGp3Gbv+fuPFJCvMCkNF
ULw0xdSYM3O8FxJtJKgP6tmyw6ZBxHi7Ij/2kXTLrr5+UlCAoI4tkgJuaeqIhHR7
OhwDh5lOFuTg0hXLsLu5GJjhGbRQFaTCyjNFv9nRODYS1TW1XQ58F9ZUsrBQJUpB
iB1QOspNsfYGEMf2KfFGj0inb1+SINvq1e47WFRsNYq58QobxNysLgY6IgR9sQK2
MM4UeDg8QJdvgoD/KlWKPRuu1YIZJfHu8G2e9y1aSYuUUzODAlZMverIQD93uqn7
9vqhYxkFWX64x549L+R0ef028vmUl8a7EBijb7xijzRGUXxOi05DCTPaPJ3hxnpM
aMK0NI5EwOmz3B1tKxR9AunEvkSFodg4RcxwfXfGsWUjMFOhN1M30bkXmCzxXX4e
hS8Yu43Ohf0ZyA1DMjxwtV0NNMk8wvljvrE3KsuVmeRxGF8K+dBZCtPq8zz3Dr/P
xPQmEYJAM9eWZZWFO5C5c9Zbf2NMTyBEiBI9bMLoCrOVTfajqVBRm2ccuvs1rMU0
SG8AEEKdV8gVUZQfWLoBYLihEqkFLJzz+McnfwWbz15ok0g2VGpF6Xq46ECP1ewb
DWVyHsmo8MFykEaMwdm/djacoak+XlhlvDFx6aek3zT2dnAYqvFbFMmzOi0IpbLG
Po3t+o0jzeOCftFQzahrW3epJbLe8ycbhFi4p6Xq4EN/xyn7rEcUaWX8grjAhe1z
uwvc0s3erAp2IhkofVNfEivYhCce0xBPa+vksk1ahVuOIAHh+k+yFbHPZBP3N/sF
L3Xo/AG692QFYIekvOpSI20LmYDU34w5BFPkHCaj50iyi1I5ECvcZkJdOxw0qEMt
+XW4MfE+g/8259JcYiQv9u5Jv9DsS1ZbSsF4kK+wwk6DMBRLtA/MihzysV0rxKFo
vU4dbzgwAxMRJ2oz4+pKE47ThyIp50qY8iIFWLiJTgo83GsceoRi/4hrb3w9phr0
fdJiHGrsuwBkyIPoDoIFIg6vMMIuzQXSaiZV95m26IEo3td5Bi6pVomoyjSjCvQm
RyyxpyHVBvQv44AYdvAb4zCoOZYRiH5Oe754YNZuo/0m5BkIl0IHD6Tn7Dr0YWg+
WHRpMPZ/QEXfhymkESMcO564mtm1kOakpwRHlTx4HzqN++2GIHEeXkgldOLa7ieP
28Mb1529ZI+Qj0fZMa/w2ANs10wPoZqsTeQ1jf6+CpAePdmyjsDWkpLHeiREIgvP
OWFu+FJmWLFsj0Pezsqp7j6ut6bzD6W1m+LV6bUUkMMaGYqIcuTtw1sqkwUQnAa8
R7W/ugPL+g2wrDZAJiW7l7BsldeMCFma3TNt9YYGm6gdbAcdBy43+j9RJuafGJQ7
lm33PTTi2t7qFmau+TqhZb8QCtdJE4SbuLHK+YmxHrBtvacUgFEmdOhFQehx0Lzc
HfF9YxKJsITK+fx78JisBAs/9JBbDglnBa2QHlR8mARzldGtyUneUfzYrUQqkxtF
VO0qpqmDcWNSRz8PNjW1RbgneHwvI9fADh/UxZydhQTcf8HdgQLCEk+CClY0Pim0
GEazlH40Ipj4Zxl8yQ9B5dhEi3LFqoTtRnntlgFFO3X61CUIGB7P4bEaNJp4DC1Q
XbU8mO5nP0V9biwsYNXuaz9oK3/ZdtC0wXOmIsmcKCMQqsd4fdvyexdtlFoFHWL7
GkB/Lhyurg4IwiNkXruaNukGu3AoyogF817tJQGE+QHgJDDlbNVe6pGm+Kx0w23C
qbvhj+8DygAgAGeMJSl7McwAkncsZZpgeTXoOOEsPa8=
`protect END_PROTECTED
