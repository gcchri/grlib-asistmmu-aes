`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yqzYRBEwns7/0bdA7J/OUPehAENr9JpsVnYLEB390c9xwBccaaJuHMCEiMFNEa2
kxHhkwtEMoMFer8T9JVkQrw/oXcz0yuVF42JgvNpDAGRDpMibT4JrxgbnOrbeaH4
9x2KW1pxWUqR+c6nflRWizc1F8Y1JiKdkGOoRhlTlusTCtteCRwkZGN5sgodaA3o
FhLfOfrXhCKMGOVAKjWrxvvAWu7lF9PeVzk0Kg1ah4DXdTyuKStdpzQtLBQ1/hNk
XShgTvZvf3gRcyAHBBQNeQEa3u1fYdAVcSu13pUf9HhdQSBEr9ylWic0j051ohVY
9ZdFFBDRzHPoXwIcFiWKQ37cgi+5n4ORIqIY/M7DrFP9hA5sGdFiYM6FkJ6ZC0Ff
RxuOOXKwMul/z/Cl7UPbbsH3uLmyEEBYiHBtXJhXiMy4D59r64maquo1+XZN4ZVC
XnUPqpVFRq7Lt/r/wkqQhcHSdEOH8DwvoW/EfvmCpMlHsFVEFRUUNvfBQl9ZG+iu
X6quMFtMJrAZW1wC38qkuHjXxI/PllHWd+7DqeAxezbwlwtWlTtX3l5NxhC3NDMi
GbHrbd6/cxjltyHngyxegV3/9jUdQIH2nQT6qYH8iiWlLqPTrE5PPINOGCcYO+2w
2W9uokUM6kkGGKMjiLLoRQ4kJHDm1cSs8pyT7k0e6jbpdLjdi7T2IBSTBYOThkPE
Y+rx7PPk8EOC083tYKjwouiTqSu978gk8K9dsguHZxjRnJaqZlvy+7FGXmlStLNv
iEQwCQ4GEx61QSQ0mfoYFctA2EDcAQIBzLpt+KBJKk79+UzHWPGDDVnzPRHgIVBE
0+djaYgN/xZBcU9DT3hB1rTZP4dR8nokn71JDzuuWUnu30v69ErYJyGi+T+cmfE6
4+LSACCrrpCr5YIHpoqhxCbQlvCm/u3zRe9hsN1n1aOlQCNbU9Z4JGm3hSpLm0a1
F9TCK/H/zWVy9GNcwCMP/4sm4wJB3SUAwncS39P6LwmXB5LRlt6gfhTsTmdvKJUD
0ASh84oX/2frmGcgBxMB9qCy6psnTAV9qPKuDCqCJb4P6t/DLjRkD32K5JRa3MCW
ayvpubtn4gYN+U1sGrvQRmgNd9Kzu/UHDYkBUHoVp0j0C02kVOnCX9KpE+Jod46Y
JjaZ9idz4jlSnoQYYWWM+Ziwy7DtBHrFtlwy1fnxwD1C+CeVSG5T/2YFvcKNj+cG
njV+VQ7xbm5P1FI1MD2+UWY/vFyDqDIuBQ4jT9fmADMSNWQjals61kWDp2qBDtNN
NXeVSDRg3Ml8Cw6gfOot+as273lrhEOLf1llJVlIZzwLBnA7Z1/aEGVSDtBZOqWU
GRHkRh1cHRfqxE8iJJgZ1ZYvHUnBa6xYivHqH/FcNQs8+O8yrDdbz8NsDCmuF5uo
bPtV83M/Ja5s0IgvgTRbITdmWFM31BVWFLYVk+5A5kR2hnkfcarwhX9fb0n3g2fw
0X+QJBcJvoWOjyqNXn0ZlzbvIFqFKqRcECUNtaOBaLl8osUR/s98J8x6BqyCOi+V
M1J4PEJjVjN7mUBUNMlBfQbWgyHJTXG41q45LF5cQRYoWVxUtASn5g/+vES5Ps/h
VxtjyLZW2QAlA3VnLJw24vYfuaG0zezSAsuRYTXvJpvyxfQSf7KMbPDBEWLLTGsP
g5u4bYwMn5SjyIYCzTr8D3oTpW6xuxNmxbpliO/LzcO3NcymTwN9Q1DOAKrInFD4
a7pTVeO1HwDM576qhCMJcqFitYccR0gNnNwPrTeK+UFbeL2tXKNT0N0ubGvupc2L
NpitzFYnV7xSjeNACZxnQDDfcIDJwbdbMMmf0JtXsyeSgS3PLQuVQQykNVBMRUIM
A0iszsdntC1gAzSsyfRq3cp6hHSHsoDcH0WLcpDc34/C2/u36MUyGRAz+le917Fu
bV8Sr/FMvkB+j2Use5bIbfReezqku0MK5tkKsSzaLPH3/X16000YrfF9Bmyl10WH
4TJlRUthmXs9AGjjB5s9LMPlD5Sv3bKHWoZGtQ6hH8DlbxaClxLjFMk0ZiAbsRbW
cYa/Y693yjfw4+kEjftH2iSaT30D3jdcA6b49T6xENbcu5Umhy96rIgjfuDEJEO/
E8dTl/maWQIBa14KCoKzKEKiPziAnExf0xKB1yFEb6mnTDGC2Sq3Yi+5KVkUQu/K
fgpjAnZfXsX1FDyNhpyYfWrLoOs874QF1TPvxBtl4iIvwhT9DFqEfwEzCFgidY7D
40Xy+760kdd5EF4CRN42zeaP93fqnhTYrXR+5Z+8ao5jcjMScz+1yss+nnEtWiW2
w69WKExUi7VQW+jlSSpXb1MIoo0R3KHa5NvhJFisq4CSYc/eMxn8pkYGGeuvjs1a
zRmxkj1172V0zlYyYd/ToY7icuv8m2iMP/9Qu50Nke1f3Eha6pGr7T0FL8OwuZVb
2yJuYB3/p1XHbwCanUadic8XFWaUTYcseEbf4zH6FfXSyfOeFCFeEMnM2PLJ3Tug
jbeJkbH7ExCdlfT2EEhOUw==
`protect END_PROTECTED
