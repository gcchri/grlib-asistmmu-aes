`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f8e78V0LKLnThF9MCxCjyGY4hNtfwVjfHYrjRm43KoOifZNp65LKhKRIJW9En04A
c7VEBG9pT0uiVGEESCIUqIDvpqKo7YkjHdLp/uXPahUmq+sDeXham5U8TI6a2TaD
ALxP5VuFUKvNBMov8aEUQiGWH40v7IwA5AYTgHwiHhvCT8C+eaz5e3deqATWyML1
HKI/VGvK96QuWhfB7smAew2JY3KmyguzhlcHxFPzQ11pAd84bzievy519wTQphgg
p/30pozT65y9r9y6Ao9HKVL5II2hjkLSiLyjl1n/gG4CRuJzosMr0gl3HJkXWZra
TIP73RFHDZ6vvZrR8kSamyvfWHKMo+vWfiTNIO1plNmFX5egDgs8Leop1yEGEWQI
xANIoaH9AUOtnuPtHTbvl8CvZZAax35gc6GeUrIOSkc=
`protect END_PROTECTED
