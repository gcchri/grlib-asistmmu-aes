`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MimAZ7hnFDvYjhIGOlkgHNIz8kfm33NgG7OUq9PYNO/4yGOkkiZn91W7Yqgbsb3
PytrrZ+ec82I2UQUBjUVJWVuo8fDsTXzgi5P+NAppXlh6oEGuL2m7w3d5rjFwo1r
h9IIsbN3yyhlXrkMNbR35qrA3yHmtmYrRlit19UVz4P5/Znydvw3jSNMNMdaGSaS
jDo2rQHtfYhW2taKPLBnV65tFs13pXMBFQUWkhnklMfwCwVZLe/HfXimVOrvW2HK
BNCBfX3GgzGWZe4trhBFiZaXaCsjCybteUeufdByWeE4rcudvPvJ32r8F3N2Riha
LRxy9PNtPhxrbRVx0RMPpiKRSzqyltS+ly9t5dsO/IHxC2LaItTLRPMygVpKya5h
JK/ajQfvjwm/4GOvuQveyKNr1a9i4j5ETgeVOmDC2pia0dEV38VdIDIwBKmkgxiE
Bzh9ECm51pK7waQEp4+0I+QzjzazDtdn8sHCV8/iPj0rsXns9huUdvPiAqaDOqqN
h3j68+9boAFOQo0xyZolr0X0JY6GOrRLkjqFIb6YqAGzedBx/4KLfBasZ+oGunLO
ZgyuYLoN3ClCVFxKWcyVWd2119a2tTLIvmh0Yitenz1aWesGhUHfkyuMFrVq/DcZ
t9TFeYsj2AYuNyxG8z65ikl0HnVNBgpCVHGk/u5yEWP6O0DRIlx6HeWUvf3CdfOl
rszWoR5+XkhQsuZtLctyYdaaxT8jt2n4cxurBZ2zleQ1TA8xJQKGRFKLWW1Mgn8u
JKvvamfqGOZCtYLbBHZyb4puG+YXBKQWLJIrmsn2a27ogunvwbahoTOC7vPHhnSu
SDOU/oTlXrTKUWIdnhbIPKvBivNGeDJqxg3g9tqP9pZXM++InIGfX61Gz3eeafPI
p1EdNC1Z1gJVfwaQ3TOjqFBtJlAKfe2PHp1HoWuSHtIa1tbRnYBmzfCglYVjU7F4
UEg6hL9R1qvhOS6+c7B+GW9pKdAjw5I46wKv0mIMtdCtRamRPvk1Vh+E255Mu81D
8My9ksTlfecypyoXMnRhmF4gOCVJ+vN3FdJQpbIvCvFMQxl0v5j+330E3hhHFsx0
NpZOJ+f6J/tBZ+/bBv0geaUZCfzeFehVhUR9gtDjpQUafPecDJ4pajNx3MPBa5bP
DxTzrOZDr2lgBGJiEYyaxBaDQRWBzfU0LlJ8vH6yPWAqI2YNobWhkFn7vta62+FG
xWMUi9IeD2rODRkMBJKtkKQqDiPsmFesFwAHQhAbNBnyZOOJpY8dpX04bHvb7WBE
VdCL3DIZzUevEXrduLQ+0O1IiAa/SvkgAcoaNqoP9eQgsOFmGsJ85W1eJlSnz8UX
U40iHlSnul08nJyG8U2hVKfHNDWUOaXlDKIKhJGeiE5R9JgGe28aOcEeBYghLK8N
Vp7kIU3purrutI4tydNZcTlfKS+9AQiI3yjEpeD3AWdn8AnmRIi01z+PVC6HT9st
LKvNyHMbjROgdxDFqXEz04SpR1id4Q9UDnEJktIRINoppQpzMiLmba7t1AF5+Fe6
U2asFdQVxo3cBtGiDcJCT0RIcBDa/+eYjiOO9L0K0OwlEkXtt+Ismm/Jz1WQ7ggW
+c4GZgDxqqDPCytiXALOqSvN3tJvEzMoP5fgNCt1FJmayhjWn828qhKQjFVdnUvt
Txhw1rjiy3EEMSYpyWbZeZW4J4Sm6OAeTPxe5bvYpUTuLR9vZaxjieQrs7vFBQvP
YYOEVmuC8cw/AHckoWi7loBKYQUW5Nt3WvI7IcFj+yQxACRImA+DqVIUJuWIDCy3
AMwY6W8q5E/e21MyUnM3WzcgOMchirZULdy49atlDoh75lQ/DsebbIexPyUTKk5d
MMwsTOK0ioPAVCSVZsTTx2JevzphvKjBK1fTYauQXAUKcmpljK4kqMYVpAnD6YwJ
o9RS32LDlS+4DlbNAQZUKCIHoz7DpIhwvAQ81S5uxZrUr6A2tLgMeEcw0mwDMAbC
m98rFOZ9NHgxiLh4Ygch+NIyDfOPD+BL8RZ/Ff7Nk4xur/YAiaDU4qqfJycMafiT
Rz9XHzMM7c3DzrbbdM7qIGVW7dD4FdmDuF2AIfxM7RkYRqFl5jahT3DggLG73dM7
zss4yCpJ8xJHoRtE1KbVLkdtK7DpL85PODW0m+fBAkFUTv7X+h121PBYGoTxpWtq
JeTeNsCw2SeWDh47wKlrpgK9yn2FHgQIEgP2y/U4ZG6MyArrQfHsEC41Gyx2JIYi
DNJ8azZ4jBko82ccVEKYGmf8Rt7i4GAuskD57cStaC9XoxpKRE8Zn5MZ3kUfCVSn
KfxhMr8dEqUC6m4E0oN2jrWPYPek4Apup8ziKiE9XqvObCfw8rYiflZ8Ias5hjKO
coFLa3cNIMo4zsSR8fKcrTF7f+PqyT7z39IUJla+TqAP310Y3T43ej7kVVeD3Elq
WGg8wDTTqdMyNtM0Bgq3AInGEAGIshkXxn4JltzUf+YJvLpj8groaoUDU6zBBjFs
HoWxwOk7i6Oz0ihxKQq38LajmrfFqzx09FKFipLAr+LeePnjO4FovILf27rh4rDK
GPGRSjjJqnEAnwgqJGo+UUJUpgqA7TAKLHd35wyRpbmlZfDhmL+EndTsI+WBPwwu
4wMoe3y6I8RYlahLjogqHi9masY2Ba0+91Qxu0qjMS82/22AG9LewwiquJ8IdOep
LfSrqRNyd8kNp6v1zwymw72mpW7hGLA6x39kAQN85oVyMcmpQsp4cyUs8Y+vzwyZ
tfBFHbJz/kzl6JK3qgSIaF/vdNupLHQQSkU6xoMClyBsfnZln0KmeFkvrgv1056P
vG6OzpO+FWMIEQA1KqSPatJ/pYXmlzKgC+IFtICxkPAD5w/x8Xk48Qt8lRPA6m+J
3dgTPYXTx/hkmhkeesTeYyONscPj7hulPjbPwSeeUfLBPv+C5beFI5cRw2yBYPUl
WRjEbDECQeOItMCV+AzMENqQ9UUQfZxw9Jr2ZEs4IUcvutAUX5ZRTuZR/xQ/LfR7
VBlh0arEYwQZ1l6saxNFbI45tTRZpuuWDQ+w/ZQnPP35ySXqbLmHEkpALMFC6Fh1
IeGUTfK7qyNsr5BIhpR+HW5o0dhG7YwwVEaqGyanQWg60vb3i/hiCU8hWPYc/5Gr
VHbm5axvqPTDo4mA6kplLCiH7XJYZlCjnyt5+er/lNgXaenf2HsiPaKyQma/h1Ub
RpbHfj+HHvYM7M6l+Hna1J7foBrmGCaQceA15PW0Y9fCdZZ7ANXt2hapcA1uBc8s
hvWzDlujwWaYGJoozE/ICzeOcYXa6s1iM3vSQ7JHdyfI6veeihaJx71s12qLBgwR
GBgtXxa6OreDP5oaA1VGHZbv/goQg1Tj6zbmCCYYYlR0nZjGPpa84LtyzC4vWGxx
1N7OHMfl2wC2pgsKQibZVUVWRpm3Rc92+Uj8fVo6JO+tz2SGufmxamGiVQtLdbo6
MtvrXiL17yu0xlbu5ZJouhlfmnqCypYv9wuwdaMNOeTOQLvDo+OmziEOV6PSYnfG
yJ2+TErSO+piDAZ+73mIah4ucRUnfzM+8bp0FId2dHf1nmKhsAH3gdlmC0KFm7kD
VSFYkaIuCwb5lCA6o4W/U9oCB7Qg1QBMIXHLzK8F7c39REVyRJ86+Gh2Hg2S+UU7
hMBNFX/wDvC0NM/GBinrAovNQ0o7M76Dfl8qgqAU3TI4qTe3GhUJF/Z5OG1qlg/B
wXeeXTiifk3wW5tSuBMMZdhHSD4190eAfjhbslB7DiMM3IS8WreOvE6tM/UMz3gy
J992aqoKSsvrrNBziyEwN+aNXQmyUNdA6sjM1syucN2vodnNb2mgYIP4E0eTL7N4
6A/qLQ1+PuxRTUoIbqrjEL75MbKX3vqCYxI5qDYSEp5+L/dtW7QVldImMpL3DdaW
eoTuJEnSYDtTvvy8f1TE+U7SkmzIBle9wLIqbE0skmGVIIbwpFZJB3/Pn5NzoaWZ
h3Yo/FuLnlDKMByxPHXZ4d8IDMHXCSgWJILgpUetI0cBfCoNn7dUuJnhpdCvDoJH
o7d/AXQMwPaa+BpTyWQ4Fmk0cASOqF7aXAEydbTyv7nx4Yxlm0dwXqM00KZ0kdHu
POgC8PQvs9P7EK5LGtaBUuAHul95unEdULfDeNqH1wj1HO8EZEkhbUou3/57+1Zi
tFI1ameHn6X14v5XzU8mQfZqwsI30uPGXH1IPSbnmQc5/vaKzu1QWuO7raTOGXK3
ukiTXioNXqpRYeYmVag+YxRGUIUOzyv5HcEYI6J6CPSY5hJIwzsaRutq2bagzYRc
Wua31Zct3JgH0PgON83YQTZkEjqRSCJ7QYvnl89923o2Q+UeZOiGTZLZBtxxCwss
D8rY17Jplil8qKYnOx6P5DWZerHCBnB76DiOAbAphW7JX+psmAU2QdE79ua3Ub9E
kYUyDLOWgsq+NCaEvSKRoJs+aZFoUJ8kEyOmFPXsEwG/ZT3/QZmXpvwxnNCQZaa9
zklsyfE7BTfjoi0ZJp9eejYt5uXA4c6QVKlw4+SwddGBXrxDHxqNBNAg+CivW2Ql
dapAmoOsgyNoma1JToHQTYD7lQ2ZsiiicA8VXGY1v/5uDufY20zuwxyfB9Sh/rOL
MyxLFV1HlC+5/Ae8xboyQPmqrwlbkYNunsobt2G2OPq5Y8Y6jJS4Dl7NKjwB1bQg
8iqgHmUui4+zrNvzMuuUyFAJAlJMiusWTRgBNQ/YbZmj6GFA4myHwOCCwxnOr2bd
zYKO6/GNphS+f3X7cRsUBzOwbF0ffdF8jn/xqIwPj7LecNIjxG3rsEaUXDxibmXb
vIF5FlOJY5G4hZUIuYvspb8ctizOcMwEaPzGeC7iVSLKmkqaVqflvp5MELMwEYUp
Zocu0WrzxbD5TisGFEoHCexQ1SPNpQdvLkb7GzU6w5MZX9fd5a3IDgvgKMMIwqwi
6g/2h3CnrG1iq/SG2DRKL1TZy36aijOezbdkmjv8fjGOUySNksuCN0hg0cfH9vOl
ksS1BaxM6BfA/7dZaLn3Q89QZalBvcWwrBX6KwghhxvbjNG1unhikLMS2V4MTA3U
FJ515xjH6O52NmXFouvY6OS17vNQi+PcvakJBJ0isiZSIkLfVQxQxt8evdtIWaUd
q6yo+vr39t82RraoUlyokGqhcH6VuFttqyY5S+aAzxBNsZwOPKrkfT5yyedx+qhj
5F3PEMbCwrE5y5fi5DUShXA4fjDil/pmTVOuIZ5QY3Vvkb+lRb+ofrz2M4waMRuE
5g45uw2RQ+343jEV6wQkXEWv8JhNDeby+scUVwh/Y/Sl13g75qEEWaW44mIQ/55K
iTiYZLCqn5yT6PStWPve6DBsaJltXngD2xJ6TipoFC8fLUoQ0BZdqwc2/FjKd1sK
NwV7yu7MkgDYGod7/WYcNVVEQtFNU58DyUI46nL+eMrdyA7A9nL9CCPhrKgXZeoN
oPVCmnTbkZNYEDDegUrSfMy2Y5G5kj6zEJLZlRbqIQIGrs5452cMlEXfSpGf4MvT
u2plwAWnH/ZCtOPLsfONXK9vb4Aap4oqUH0jLFskAxvtboBWV3EybbKRi66bSQPu
6tNQnXMesToeONihihXtWyluD3dksEeb/lpCt1L3tOmSCOY96Y1zPEtKxVMkhjpp
yCPBWGHacc4m3MjKj8z81Hk2J9iba7NeieUluly+CXyUcSZPCljmaaDhGjLVWGXZ
18HkLoxFe5cKYRHvr7zVqtksG6PbVEVcHqLrtTx5kPi12J9riYdbDtQAabNGHCVv
d3Xl3tAjwBhTZaeCbnKCnY56nTglZKDBdrRR+3VqCpaCGBAmCmicj/+U3CWH9pi3
19268lRcb4IN8aVJZjm3QSO4b9mH/vCnz3YdCoT4nuRu2v5eglwx/TvSIuGEh2pB
nn8MDgGT5tRSB/iAMcqkwyp7lx02eiReDwbBsFSXsFB/N1Wv3ljwZrGh8UOSZOZb
2245LvYcxQ2KvkM7IhvSVZwt+aTaFNiHH623mc6Hz4jBmW7YrltZ8RsDsLnQwijC
U+AxDl0Q5fW2yx4gwdBOQXPbGBaNHpmJS3jcSPlLTSltn9Mcx0cHQ/+DE/VaJCes
lHRVPW8cFlMXVfoGLyX3Kq8/6XRjXf0Epk/oQ+hMa+NXanUkvMzNkPYaocdUbljr
C9K8Wnlic9mCMwgKP4UiS10t6KpwXhfcUvGul7vua/jMKT11CFv0GIaZbp6OXzoS
w8YElORNR6I6ARcWhB1V7yDa3sHqNwxJZpLywqqk5IHLxZ6oQC7GtWfGYPMcKRs4
U5Qb8BYVXdI2BJqXedrT8GcM5LHan1WhWHJ6ahYZoQjMMmV4RyzIUv/2RrbBzX5N
atLSH8MZ80ba5pF6eoSYcK/OuTHzFJMfgDR9mvtbLPDZLZsrJWn7gRA+HHMU74hR
cBFToDog4Wr5qW+prbNK0zTw8MUQqw4ywKOA8YaR40GAAQ//CyKJZOeNNZ69VSsg
e5vWrCREAhXeicyqbOZWVWvZcFwIi+fCE7e2f/3uD6iuJ6s2vOohlM/ICFt9oxpt
Ug0tRrIknyl4bHwz+L/sXjPdtIYZaqQUgmh0D8QrTlUqRtwxr7MGczug8PwDMwb3
y8AqPl8HXA/6afeFSOJNsqjMPLDiG/h/Kib7VIZ++/hV0ndl+g79J+LBS6i+xpd1
vlT44KvlzwpYY8PSb97tVFY33KUeWH5Y0aqS9b4A2Bt07REss8OnYKXtoVzeWU31
xw3o5wnDih/rXeYEWqeaCEn/UvYAdq6EoGvlmpSgKXWcY4b9H18rWvNxTjMwhbnL
tpz0+va3aB4QAcviK9rpFQmwomdslxRB8QRGpgT4UyleNk5pcbHwWaHTJT8oWfUa
buA4VzlsbnOfQo1HSY/ETKKyGfrvKG8J7gu5bs8xN7lj4c+RQ1i9mUGDpxb9trpt
torgIxb6dIbNkCw37dBH/LOO6c/gf+ldYo78T8aBi/oorFc/dYL2CvRdG6Y8bW7Y
neNq9ymI2CD9COVDPBUn0Dw4m3suB6ojyWLOylnbv9HZi+qpiambtoQF2l87vhvc
KOn0VDBNBulo6tmrbTpss1kxjM18h1ObB3JcdE0PTAg184yurgfmMaQOsQ08Yx76
ZIx/PrGxcggbRsvPMy77jm76ooLgqb4obhrS7szLZ8K2K5Vq7ToTNi1FCDkwdVxr
uQHOMaFmU+5j7VxQFpCCQu9W4b7pRf3EyW00TSc8dqqJR9+JQfACZs7ZtWu2DRwi
zP3xVRS7imvAHYxLNioxJNsXfAyvIdU8RVh9Z0TQAaSc388oxjnaepjwJcldWtm2
/6tpbItkGJMQxxkbj/uE9nTc0XKAf7coRSL08UfkyZC6v5BhaXWPoFYCiYGUBehz
H2a4rq+ekeks1L6L5NPOH6A4lW94IlO7n6T2KXIEln5cDh7BgKegJeDFlkCmPsGi
V5G9pChiuo3sA8DMY8kEfV4HrOs8ZTVQMPL7DkH6kTt9rvOi6e7peohEFbxl16Hl
jNZGKl2aIT8yFgVPRhHj12qxbRWl/Ysv3Mn5C9Zg1E2Hz/VnuH7CAO1VfJjD37tD
AzF6E7Vvgf3AheKAJJwPbSypPKqMI40xoL078VCnBYyyWicOMSukgnAULaIbLFGZ
ZQYiFrSklc/dxmFYkNHa0BZpiXjzEjN7OhAjGMKYJOH9+kP4sQq3Hww2A+nBja0o
H6eHxf4fChztsOxy50H+9fxsQgCi0FzzTm84N/FuvPqqGYYtoKjbT2XPdSFIK+AL
nCOLO9VEkrNaZxPe47bFQXtpTZFcLObnOr5ziI7ko9BOx7kk93CdpUlBkV/PrbZb
Y6jVzI7vTJGLlSQWYUlqkswxtK/L5gMfid6vNs/cwh77Gim6LmRKOM9m2AAqb9HQ
oGO1EhwVBT+dsgEG78kTpO4Od+/pg0by0H0mLWhn3d8FAXH61qheF1wVfXQT2s04
e1RB+bEtxOhE2hbVewekEsJnUuZWXKvdsDBwi/8o2KkkgpZhrOBRX7d8sXEqB7Xy
RZaopL1v0uGvrDXuw7vzGxleyPWhm7TKKpf9Msa95VbmE3B9/azJTEN8Gj3O7UTD
+4LNhlZNaAToP4mJXUbdQzwbwBEicAP2PGFl0GimsdzfGMVtctapxw0U5OAk9KYG
uOrNhA/qpnuW0qBzbS+7gVByY0fLaE0uymRZT4RrFTbamG0Rnw9sgM3KcSxvSvxr
9iY86UwSoGIt7H1/SzN5dgN3y3IDsqdmNnFnPpmoruEXdyxyeDMBEEFDte1VeQTe
9bDbTle0EkhuZ9j66WlICP76Q1k+htfZOZGs+/RGOMQenn1foIt//ghrsAfS7N+I
SNIx8sK7cNx/ahbhY6rh16tDq900aX+nuc5o6VoMHNKTqwQJT/cKn0MQqTjEBJQJ
+jrkVpawFY9BfiOfMUe5ucFEeDIHB3u4zKxjlv0COjqiSLtC7TcRVzVDsciaa3H6
+my+z1O9jk5Go46y0wuffDvBIvaGUFt6Z3ypMGGsF0UlGbAEK5Hgfp20a6hVLqZK
nKfz68gs7ZlnXYTIfFLDthKVqjahGEErHilPdVC52EXv51pcv1wMG8X8gCRRHeKM
N5qETfJk6gEsRJ/JLKqTHZ6bw6QpKVaNT1CaL2BAMLl+G0LgScUiOnzUqn8vaSIx
9LVENQgWuOS5wYl5yd3ftlFrfv8K3SdJSW56Ofop9ITvfDVgPHj8d3gUnGY+FANb
9HvoUQhL2K0XfFJ7npe/f1GYPndpUa5K6hE1BoVZt2Da29E8wZZBUN4JxIHwx0sx
yUMRJrL6CIKMOT75eU4exzXBFK3m+DOBpN0kmd0wjE1cIHdN3f4kRTrLBO4i4UVa
+BLOCZowkEbPFRJ6w+kHuy3kX2WZnezlH1V8ub9zO4H+KkMCO3joOT00MAmaQOdg
ZdfuHSFXpIwWNWjHfrAwPF5/o4VPlY5hb388JtHpEeQbstc0hK5+UoQgTJegGiaT
Qrx5zT34qRDcAlfAx/Q2PHXmvf9Fkquds4vpJ9xCc2zFQQQmCEQnmCGtiVr0Xu6k
zwE0E0ZomTHNa16NFqSnZmTl86bidP7J3hQAhoVYCogfTa7LLTWlAyhT+jI11iHc
vl25+jfxi0uVUrhRSMYjepudNKzP04KuV8s8v57Aq1PPXPNkYwYQM3WkdZAwMgpw
260iddWwcih3Fez4HopTojta4g0fGh1LQfsviwHhKuBmOljKOIE62TygvYxkBqnz
rZeTTEn4jsymG8Hj+lgCqXZ63sCaxHLgpPpb3i4DLZSP8D2BJRW5OkQD8CoSa05n
bQ3GNjc2x+2Tt/b52EQJqYZmVlpMDk5B3hAuq73H79ugZOaNtdUj/L1bfT23j7fZ
xjL82P9oX3++xicb+dAX2MtmjEhEa7Qx5+PQIpQTAqGfs51nJfO+i6oMAuxKQ2qY
ZECGb/2jXmCeZY6yefLUc7PaNSW6E2dD2Z5F2MGC8Y/K4WGR6aG+CyQtL/QeL0f3
t1daYCFJdFFOoqUYfiGgkzThk6Ntn+m8hXBkRm9w8EdLESn8hQsgsQTaKODXs+7S
imRJu7DL/loTxGODp5SG9uMHcrILoYETqm+5pOo25RsaaEnN2Kq+zzzL7VWTK8Zn
O3iIijNb9oQwh065BqphhuZIb8VJTxMP3JTodVnmJ2XTWwl3A5iJCgmc7cNGt1fX
yt/uep0WM+lBNpOBmcl9jsVo219k+/fQ2b6fN+YVICZdc4AJqDZJ0lrQSGxIcDIT
y0DzteeBPUCO5XPh2XDOg6BNvVCctCvx0WVqFmpMDiQNOYC8OlpKUqrYyYd20Gcf
Y0lg+fgvGStxr4YVFOOLHbvDtyOR0eG9XG6FIjLKWPqzHgbLnTfC2gKJA23Irpg2
`protect END_PROTECTED
