`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i2EvI+Om4aXvU93V1gJOsnZHB6+a3mrkkNR1Ur18DVe6Zh7PcV2TrOLb4qHZFQjm
nkjLntPWnfDqmNDWc9lszOWZAZbHqtEiuCbfiVufcxzaxuzfX5O5bFABp/Ye3y6Y
QhzcwbvSu+gavD1Q3vCxThe1q/YDNHojXhRGSFk6oZEGaeWTT4Vpz8bxgZHSeXgh
Ax+Br5gGgPLf0lX3sc4XckWmrFPt1H38JLkEznM/wau+tKxGSPjhqTsMFSSxls6G
+88aM6TtCmxzRx32OOB1fzcJ8YuFzDElIRVq2vxaogVlXCOTBjQ55Lap4rEHWl09
9uxMTSADHhsMaHouAXBfNWxmcq/1FsO8fBS/ZZ6fsSp3mI93eI2EkpAhyYrzuO+e
esDA+q7nENjaOFSpgxwy5MaTWe11O+2EDglBXEPhnjpX8EsZA4NGY7045HW1BSyT
4d+AtnMVTLfdhAKFCEKx96I+M372lrl4p1WszXwX258bAvHXpUI+HkTc8R2iAJQN
oZVgkLvl3wMaQpIEnRRYq+o+ZuZsBx3CotuDe9WRTO1pfN2aMVN0Qb6UCntA4VEB
DsmlYmDz2engfvXNLlzDonfz1xDng46FPVh0LKxgOP0Gz02CW0tF8MVzHXlwe+9I
E2cRjrgzeg1mugdlM0lsRBWGYR12oQAYmDJFghvJvKRow7e/m4VfqMTPd1GTr4Yc
mVm+RdjaFQYIbhuJLZDpmvApypcd1yqjBGV9vUhUBb7B/59pAHcyIYidP4FxHFUV
o1csI8kWoTymzckbjgy5Xp1QPri2ah3gCs1/43+rEddcKumIU7i6cVstJfivhnV1
NF+ron2JIFdTbZbGQ/845y8QQPZzeAlc0EGZZl5Rhaq2sEpnc/CrJzRmcDheWyzT
XdThzbWW4E8lMmZjwixVciSmT3EqtY+fFBA5ot9suWcOp+X6jDR9gYpoaSdqwoxS
ncieTKPrzLeJX+ZoTKkkXZaseC4STJr8iqs365sP5e8jeK9L3B7D89jSKXuuxrWn
yKWACxwXI8n3WR1YJxQ1qe0oPoYAIpFV1PjPl65sSE08I9SNw5SA6mcEEnzIpuLn
DRUE49VInl2T+FVdLQZra+Hx3KPk3Z5gmyxEYLzo7ODvKQRy4XHnkLjCnmMx5f0x
zKJaL7RQ8bCbpM7PbNUpY9lSfr7D7Fexh/Rv5DQZFqFPmJLp9OsH+DwIFjzHfu0K
Ngwic7M/U05U0S3+wBh3PRLIADsZ5CtTVGHjtrIsVeiZaz5EFwqahV09z3SdHWH2
zZqg3Ryfbr7LMA3MookSMml5RRqfCPkFaerKe7d/hHOHeQ9ngz0CD/ZDKT7im4mH
95MiAKuyYPrw+VQNfNd0J9j/fILbGBBQdQMSX6mnwy2NCxK8bqg7JsbVCD04l0EO
r0l2w6ooOUr90vu/2weRKGD/gf1xAGxVm6E8I6yHBlDHunIa8gx3kY0ksT5a3Zlz
FA7qzm1kP2p4qnKQlqnUWC5D5ngq4RraHuheGu1gPoetEm1KafGbuWCJy31LsQ0u
Ywr12njYZytHXiVN6yxT3yjwUUnPMi5ZAsArff2nTyX80kdPLXlXVxa9wDUUsaua
tHFR1VH5hiq9CrlHd4FTE6T+t5ZRD+xTBkcKgFySpIRohsOVACsSuyxeSb3ob+cH
BexlXIsdzAO/thiTA3W+ZwTXzr/oOtXz1JRnC08qicCTpaWZQtVg3p79Cn5WY9Jd
sEvxjNKG1v5FRElwLU56JYWb7vpQm6eZHcHAVQI1/bSZ9piVIpDUmWed2Zn4wJc0
lPrPqIP1IIaZ0ftQkm5oIsYa8DUca9O5Z43MoOVkxCcG08YhTPNXDbkHNUiyhyPF
zdfckLBh38MX+4uRLfOHNgbE9JVP6qpDaL1n4OIaEYyV7XSPY2UaNvBbBtyeYEAt
X7/R+eqeUKk9Ebpyh6bKfhunl9Uq4Xr26PSR4tr7VAs=
`protect END_PROTECTED
