`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4nz0UiyLwen7P6CFSd9k1ne44dv/xqmSRX1bD3Ox5WAvi5OmyJ80O5i2Mt9V5l0
VRdH0wIionc2pSoCvEw6a/SXtNK6njp4fPdHA0+5PYB/UcuCNPhYzGl6dHL5rjSD
oAXyrCp+4K28jFSq754Mo2QOVcfmFw4u//hXtw3eVRl5E8kdb0CPs9EezjCXPIGI
icBz3MPCguEjsHSzYWjkGxE5ALvYviKrTXx4qLG/FRFbzHITft6JRW/SVE7Rr+8s
dRVBVUZOlnm3T13BpiM0RN3qFIvOH5bP4sqh6j45J+BkPnraZjWHtfv/z+plA0ch
HytKLG/qrKcXrIdBqM0iNJPkeFT+I7Ag4dRRklL5t1w=
`protect END_PROTECTED
