`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iL/mVmY5EZ2rkhqLHFAQqLyizZrTqKNrMfdXpDiunIK6HTPlBcRtVYuPioX9lrKz
aIuEdgxLLJjvdAIFqmvpvLl5N2CannCRKd/RaZoLPIaXOwy312gZf83hAP7sldhG
p6Vw2N2IGYjfumjA2CtyDkNMUEvnnpw6Q7RFZa8pcCKRg21OnQ9iuHaYr1srvXQC
l1+tqP3ntXNhepAgW8w/A09G6WvzWzoZuFdVfupyZOBdn1PUJAHhvzXA8GoGxiJt
nM+QImM1k+vdBUk/jAp/FfWpQJuCpXAlBFo5G3dVUSJ0I2oYqxR/sPL8qINVptOS
f9EyAr0TACUCUYcKzeIbaVrqFIcOTZNaOy9A2Spa9cJDKidAW8hz/85+2wecErAE
4nnfDG8KvQRQkAbgBNY2JkKpA9UbTAzmC8p2zdRdWauzBAyV+a1kEwNVEw9V6XvC
389wW8x4azapAD7sFuWoBO2Xf7qoE578sZksJmSjBviNU9++GxvcCTLJvU84Mqre
5NlCn9Sx2nMjdkC1dBoWuiWZKpHy5bKT38fsrAXd+UmLbE63oUcQIRMBDWNjbWGe
g8Zh0ekbxwO6g1HKBcVlehLwwbl3v9XBbzzmfob/F8l5+qdU6P/EPtNBuqFLO53B
9S7IAHAoDt2MsIZi2hWyxlHhaeCmFLZTZCfyRtaHo3uXqUMpQ2WkXe2oWEcTL1+V
wRF2iLV0phv1N0tngzRP2WoMZxizKO1GokSZNaZqOvyZK3yru1ZFc7q67M9A8JTJ
QrzQxR6L6+YdmoIBnPWL4wtF1whWr1h2aAY726SUhLTjecjeWUaReFgBRIpVWBHv
10LuQ12Y0EpU/1T/b/yizAJuQCl3ED9DBhTQmnAQNqwQSao68rzeDulelRXqsWN0
IN3iSwGYHT8hJzGC48o4A4cKNFE8hca1CZ65csZbOpamNbIIU+qFtKTIETZKDr0u
iLH28/VBQcfpsG/cO7G+aJdZavTZOcFXT6M/REsOTeW75h1iRNY8c2SxZddWQ5cr
fwzCCTSKflmD0zaGaxT+wCRtRtj6Si3s7BvQZR3RvKudhKZxaJmgkHJkJpb/28T9
7v+8Fli6DXaDbOPa2adsr50YtGyDjG7AvoZrDxshtgdaH37BM4tjsD9F2+5V4uAE
`protect END_PROTECTED
