`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/pE+uMWlRo0udKaWaHUAYiFxfoIKTCcnhWwvrcxE+6u6ycS3N3oJNVCBLhEq6sr
ysMwrAKbQl6+9u+/cJ+dF2EFZ/srZmD5HfWYehOm42DnjnPB/Ya1Q4uZwb3zJLn+
T0DHvXTiF166ExKB/XtLL/cfF4RgwR1a7J4F1ULnAbnrwA6w6177VzxoWyd3YQMO
19X9jvFSmf5gx/QKnG7r4MYScO4cpwVxDGqEQY2GMnb2DC2d90CsJFffspMJvWFa
scK3uB8/4tdqf911SPD1JVGuBs6/slbl5aSuXLQ2XUe164b/HuED04HHfx6jkqjP
yFew4KdE2SOrhEsDcicoU75TB0V6mIGJVp61vCqwgngDIDAKCyaIPiICGfQ131PF
2JR7jd05OkwLLF1rjVj8Z1ock9NZVv3iilZYwFhCIHMc2jOsScoQoiunBnOP0Q2P
1ZRnr5bZzhy0ERsnIgps3xoHRFJ8zngYu9Td29nt/bmf6WLsz+R6+QIywZIF27e1
wMoGMTjOebVk3nxvytiwS3JKbznDkdfkOnULSuIhCyuWEGhrp/ggWG5SbxsTjo+b
u/VuDotRQvzRzxsDSLLucHFICRSA7LumQMKdxm+izd1ueHstjeQhvCLgs0Jbn5ki
VY4LbI/t3ezcbnEXbdafI8ielhjaR/LewlNOa3VMC7wNf1O+4sHMD1C9BLz80RZb
ZHgx6tn5ZE41JfFk/b+4IaL1jzohaSwQ4igYYcWneiqACVjFT0xstVMehwkFEjNc
IB/3rpkzI90ZfBpFhBUVav1NHOn8p9q0VAJyz8gSyMnOgrdlLpkYz29+jeChApJx
Xg0g4T2y56t5eJN9RCHwG9kfD8NduVbOqtSQjOPdMgVZvdnqMhjirKGTeIJPRn2X
UHZZ1/mY/Q/IXxjwb34+Cr1mvTziL/uWxuQ2TExJLCxKftCCoPDpIvvhwjplcHu6
HFTY6Ab1iv0lgbSyTPq55d52Qgf0niLZ8SvOsPSQNDPp/LTy4e68YK2+odlYcoNz
2Bi2bQjV2HP5ttB/okD76b2hCPtao2BKRph5IAtcVnkLb6N8vSCtu4BHZ/uOQ2Vd
Zb8uN+8OfhLMzYAXNsPMR9hEm9+66kJjQNd5GHWZR0ijK7Z3CeymYhDuBZPqELKa
7BoMXDBNb7Lxp3WldaEJRr41nYaKy1t9ubF1GMUBkJ9tvjdb41krevTP0mba9k9N
7Hk7uM3PP5Eun85oMC57I+Tb0JvwrGebBQSLSsKuXUNszldRsu9vjSh1MwktmR0G
V4Egv7k8h86mj3mZ5Zs91H+AIrpVYIhX9XZCg3f4PV5uKV+pKLkduUdYZczWaWug
KJ7GsLrFXHIFSbHxIGiKxRFdrZPjjAE/s7NwK8JgIE6wTKschKMRjfLA3fX/dBkW
XZJ/9oCu//UV4jxdV06i+XHpvlNYiIggsWa/X6n5D0UNImsSVwY7Q1sqAEpUnvQ9
yxMsVo9JrHfc8HMCEfdv8sa+NKoLh56E2N+kSYSdymLPkJYqb6pv2JXqcRDh2PPG
95uPUrIiyujXo93Cq+vvF3WMEgKGZQfZoIq9oKUUHJBlmcT8QX2ZnQUZZrOKZyBH
/t7VfT2+L6ziVIEWj7R0un88NAyHg9kwWIMb4/CGcWvov8e924GsDqbesfKnlGjW
14qftbhGD+02G3nzwaJJNPALM2CR/jUM0VyzfZtJ5zcGKabR5/iv1hIsr826S1tf
NAz8ydJV+7Ei74Bw3roLrGrKvmHnM/VPY7BER5O9u6rNk2d9lPntTsBOgmm2FHni
fOJv91omgyjSBxSBoHKo/HrZWBKeN/poWp5feX0wHmhv2kaH710HXsMX2VsuJrKH
XtVWf6dC1AGIxFbBkW12OnCoGsp62Ah67QvrEKfCF8oVarv5KU/J6PwO+XQwziIC
yJl8rqY4pLqSdouWThUrRP3MkBmK4GVTeDJYAzltKbSLCCKRczRJryVBRuldYeMa
iTOqG+Wo7T/H6L2fZzqabDu5pkJ6+QH1cWQNjnbls0Ibs4ZQwCdBKp+Erytz3Bq2
n/hgOYZiuJPMczy9Upuy3uJik0A7KVXc7He/IXKkP7oeekq+5i9NpYojDr9rDuqq
ZVcDFK5wd4IVXfGAak8KbbGolMmw+zHIRGkd4xfEdUwKtptEGRKrlnwQg6faMTPN
2XuuKYQtHgcofIgYYo3y+031uD5UFSvfxbqYSpJdwJUfyD1bhUKic79bzA7xh75W
VEU6GWTJkNNcgzgoLU7yOxskAEZV6Mql2dqYO705hv7uSqD81MXN7DIhFCSJUXHk
9LCPmjoK8TnCuWDjRmhQaGAw5qRcwPIwudr7sJw2wvkSJEd76dx7cl3qSr7OyX7x
954jHzq1wUYW1QaHVDAonpAQPP3uulhyNbsTyqKyCJCdl3lZhkrLcx6EkOMRR7F+
KUblQuhx0MSdMWwKTO0ffK7PpygHx/LhFpTobZfhuLFqOvULm5uPbVOK9GzcHj5i
TTB4cGCwWfK+kVbSjXRJ4iyC/ifJKQMEz+GbfCgxRdDXp05YoI17yWjqskb1dmAo
p35z1Zjmk/2a8N6pl1mgT4FUvuECA6RdNa8R82VjiNymyNIwPl164ux5g4YSfsrb
h8DppSi0QxNdnQwV9ci0RfjzOkBTKHhuGSkNBxSz7NGHGHmQm9QlSouinzU9vKSu
PbGIEejZj4TvCRrSybBs2arycPd7VZ7qHzbT2BatD9BDXorjUyVtKlJBbKsF5Pqs
tgkq6vZOJTFDD09PiSGH5isB5hmADj0FGk4WDGUpR50yMTuyqIsP3VpjS7j9w816
GxDCEyL0mhHYHmfluGpsT1S3HiwmXKKXhYr2xEox0aPtmcO3njADJj7HZ01KE2uQ
9B4oDnGYANzswaVHLpWRLmiHYZ+uoLv5tZDg3BtB+yzBNzuKsXEe73nfBEBX+8j1
emJHtI0AxS7XHPjynOzOmTCI82GVhToCE9L4e/mHsYmmGVswYRO8sSUkHDP9zNBf
OxvgpBhGHfh7xaPxunxEva81FuWHtKPdqgNn5ZEHtVyv22XWNmXQKKp7B72gkLMz
TTG4yw2f0XIrXUSoJB5cpybRSI5on4N9iYEhoeUIBtfeLH/tjBYUeP1zdEhrxLJl
cQYm6N/cd5mBNjg3bLgc36PkbhoNBcCaECC08btYSPrBvzO6Yfva7lxgDh8Qpdf0
UuMbYQ101ptxtHsi9Gc38IeoVbQJUE9GNJ4X1GIaTRy67gEVM4A3Z8YX020Q0moF
2HenvgaVOSMr4TFpqVvGPBUQbUmZjhAOl6a1hy2ou5fdqKm4A7IWMJd2xJ7vGPZ2
3oNmM8ENuB4D+eSIwfyqirS+3wKJgdPzd3t2T7J/3vJSg1xTshCwZW4/igmXtib5
RoaO6gUOLYyMIFkyAUlPrrGePWc2N1xxRqhXA+tzLmSczoghsuje/eLqk7B83yao
auOPA7dBQltyZVFct8AnUeedtauo1uX33sw5pux0xe22qW1zAsrOOaz0iQ5J0CC+
NuaZm1S13FPSh3oJJpU5twdrR4HqEI3F2n1zqBwFK4EhZ47t+zyrL3n3Mb7y1wg+
Wq2ReW0fTIE/posl+12HShF/hOeKo+FH1ie5mGwmDtP7cjdET3nLeMQRmFR8/fOz
ytCzs8t6rQbD3sSks2kKGW5vj630TH02ofwqEtyvWJqskDnfJ4oZ+vHGV37cQm7X
A7jLw1Jg9BgW/t+oqO2pieJEdBODThnPnYPRyUqCkshUDJtwwLO7SbnYBPXl8TkI
JWFQFQG5VT3k4JgBQ57FlMt7WTvBzHW8CTYgnbI4G1XkOitLeZwpsCpTmL1k9OIk
XRGl0zqP0D0snnltE4jpaJj1ULN7JPuucA1sG+fx92XCj2KOeK/V2CPq6ty3Z5NY
bZdQqZNXeX4aNcFajuhApLQImCvuv+0sa6JN4WAoGe+zFmo00/YKhk4JnRZBV9Hc
loLQyJPo98gmlnEKrCztF9Ca2GPOIxFwkz+hy1w2CnoEPKlQoeYap0DkitEfGc+Z
i8VuQZ/riqzriT/XNkKkWR2Qba5AaRg8A7pi9ruo2XA/X2yJab44fDHkCfCB6Cda
`protect END_PROTECTED
