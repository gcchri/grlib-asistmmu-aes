`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yvb9ajtSK8Z7ofsfN1Qn91uynjWtTnDslTWkvYcLd9a7YssBp5W/x3X9ksuiKiGQ
t+hrRk9rcVHazGoTM3la/H4VYjBOnbxjU5ag+CEEe65Fd8KZzHvpYkkDVpp0k/z5
DZj+P7y4gHfAMUKK/SKpvAo+kvc5Xu392vaFImrsLQCngrvQSVtScfXcNAT12m9u
JOMEGOzGnnYr7sGR0XSqvO5UKiw6urjqBlg/HOxNA6IxcRxpC6wPLDQVCVK7RDuW
p9xSRYcZ8hgwBXcTV7xUmquiULHhLc24ddMj1nXz284Q9S+VxhowfVIPe56QslDk
R2mNKgtGQ6ovEiYZHCisEW/LK3klsbO4tEIZsdYxEXqtF66rwAUlYX6p1MRr2Am8
c+Dk/XEmw/yojclfDRlNnU66MMfnWJ9PKabqM+/hoDM3LrN8McSUPnoLzS/LMBXe
5CdXRIABaW+scsn8Ow60VI/c7K/9uwPz8QfsFTixOo2Y3L0vJpEpIVvIAb/iO6K6
Ueoik3UNO52kEQzxXwjXSKC/BtWFQcr+f/ymmRJef/pka1Zct2ZUSs+P7JLzSZoh
Rwz3yP157hfaQN6AEYUis93aJdLmGtdkHechqqyYF6Q=
`protect END_PROTECTED
