`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j3ixMGSK43Am1DZX8VRkb/Px6TfPV6P8m2zKlh0MH0c/8jfi/enT1DQhG5kl6Yce
ZGftZGS00d12H/8wU/4SyR27tb+HL/5znwlZqoEeeScjGqphk98DkOkMW26ccK2w
I5FPhlhYjKCW9qozA2Y/hijoAJ3mOllcsALQ0wSSPi/SraSZlleCE7UM/f5vSIIo
A2o2VE4c7dNsmx/n2bYHx4PcPlIsjmqvR0Rc2l0mC2n63IyTWRF/R9mnBixOp89m
kGmZV0wcb+/syicm5LtaJcyflRktIrbEMDoXQ8gTXroaCTgKv8elri9EFNYNQyE0
wtfX7F7moXcrjtxJRcUC737rn5b8A6DNuW4DOFNkWGP3ynHYHSEV0y0s8MW3aTaB
jJi5BHIqzmGIOJWAByc/ETPxUEcz4HecLZz/ATfbxs8e5Sfonel0PfVjXHWTlj5J
scjvnsF8Mjde5VjYfdMLb0LZvPA1iDEYKowAlaTTQcX+KGwktsNIP9NMo3I+VulU
eUNufMYzgmEFP0Xs8ygDWdmdJ2N4vtkgJPKHgWbW2036lDjIy+Q7cjB4ogvl2BGT
WIovPdYrzBQJkBSQXliMeUIPIQgK4Al0AHgYp1PV/MoG6Yp/t8pq8QKcD3YsI7PB
P+vI7MqRaOYf0dinBhEOVWr8nkhJNsEha/gsTC0/0Wok26LZhrjWlucvONU2w1Py
Sw+cfQwBs/JaTByjsPZKJWuwizN2Oa9CFcjYrZ6qLXtX8vihWiU87zFLn2oZT0lj
Q8rF5OdTHCnpw354Ewb6pKb+V+CFQnYywvtlR83FT10ZVspEjpO5PG6gWRAs64hj
RSJvwbbilPCpOO1xUNkzdNWqsousd4WREgP8K63QQtF4LWb7QXybwaKMUjeVqXB4
/ampO1JDLCz6FJ5+3Ca66xdxpVEZHg61c2QU6KEk5HmlvGDjvNNIIVN2UEQBoLxd
83Reg1PqyWcAq0dpm+5Azg==
`protect END_PROTECTED
