`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Huwk6Zra9hVF3DvF3EiKVqPauTR/ij24NFgNc5T3kcnXYXykafD/+fjXrgJ/npY2
7fIFv65FtuPvYgyEAFucAaGEztO1DGOdZmOl/GsipVxYrTGJnbLxAjLHNT1lkYDh
TC7uouVk0vPUl0xO490eYLtpeowFh/irZlfmGPy+G7SYh9ga2fq9fVYOQ13zcX3G
/yAjDH8NfAHP98F7boyRAZb1m6AMn5d2JPFGrH84rvZZWiq8nM1B0mVJsGEtG30I
j7MAxpSP9eVOYzUSJOGUQxJBQRLQGYSOqwtnCii1pGampDe/2f4jfsK5V/6OzLGV
b2Y+jW+okpXAouBmkCUFHqv+0rKdh1LEs5q6yytFMsb9kwB30P937hCsMhhe3jvq
8lrPECmCahZOwgfZ0NvPBiv0/pDkTapyr9cdg8iVfAaKEePxElEDu3cp9VOoVDOq
oDj2CZPmo48ys4SMBAaCBHKeNy6ZszwQGFLeD5IinYvdboSIKA2IS1S6UWP41y2K
HHF335oHvaHXHlWPXa+ORForN/6frbne+mGrhDLzWA46zKpG/W50MslZCu5g5Ysy
TnaKLhy8dTCZpWnkaLkQNyAtWsTfeLK08kFTLoVsniHG3Xe4B0fkxL0xAhIFXozI
87tvUIWX5eULXn4YzMAtA8ug3MqOdKNPyUB32V5meNMS0ac+g+9rOnHEHGagsyzw
zbyM1bOptXtmO1vhbyomrWBAX/0zbSEr67T5g43uzKpx6orcL7vg9BkTcWSaOFlZ
gA9OwcXUnsBX/BnOjd8e2ccP9MLQd0RQ2qwARswc/A0V8fDLbcGNi/Z28NI/ynCT
Das1fPFU4Et6qNRXqA5HfSmHRGHPRVDEo3FuMBKL07fIc+FPBw+gAC2DcKxn+HIP
lDnAPFB8q49i4Nnd1f794g==
`protect END_PROTECTED
