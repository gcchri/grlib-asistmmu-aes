`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PuZw3P3DtRPFK4nkZI0rj49Z+Qmw3qWAPaGYQBOBFvEB2gPmeWkUk8p7IpElxLly
fN1W6wpcOfnrRsStClqigOIW1NshmQZDeH+Cl4O8XP1t3AKszJcvffx3wjyCMwNt
H/bQrrtcGMuUxe81jZM2fQ9xwWXOqtI5Koy4DWoDcaX+m4MpEc72LlUew75Om3mA
QSCPk8unOO58m4l4yROzhYQLenyb9HEkqU4Xvn2YUyfgNqjHFlyN6ITeERTEkz4m
S6nHkEFTKN2GTtZAjsOGKQzNVkQ/sRPYApl3dI7Hh+kwlic7Lq6npgyf8ALqfmF+
mlILlRvPWXszJ/9VqQPAipwtuAzAatfIHABTrvmGSgoL+brIdiIZ/xF8XSDVnQDW
Vxr8VOJmTgJ2FPA+EUFnSq1PczgPy17ZXoyjU5/+/fqxyjIo+xO8+PmCLsYky2E9
`protect END_PROTECTED
