`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmQg35FdhxHk8AFbF8rf7jB8ZhgT09cDv1s3uc2DOjPNuhUZNr2B3/lOktMQLtad
QY15lkD2bL5VYUE6mDtEb9uJHllUyaXorMlj6yJn6GrQX+iS9MVWWRvyaT0bF5cp
u9Tex9uYqk16nmtDNaxHaN7R1GX1nfJ9BH55LdB6Fko0ZXlWL3NIuV+U0UDTfrkK
wcnRjGgpZwEA5GJOC1Xc0Va5I0+ZvS4uiPh7k97Mo2Xt3bJR498b8GYasrkiowue
T9X0DGdfKAIzGBiyQEeep0AekwanUH/dXpD2r0FH0dFGNdNdIVuWGkOifLlmTe60
0B8syeLfmL6Xg2lgYhzRDjHJIhkA1Co87qYVfFeExVK+KaPLVMtZzxT6qIjI7BLs
Ct0TZEZmdJzNAwaW8CbJ4Ra0uL38TMwlgzS7HcIA1hMhijX/gSFF/hK0ZiszMPOd
6do9TjIozIsvJglandG7IaEmfzPupGgSVVKvUvmvFjGXmYhDmjHoI14FNFQfRLAc
eq/PcbUAEbndK4ON2/E4UGpmCNtIAucDrdW+7JPV1J8IBeBoijjq4y2JdOTqMuzt
ipWtPHtJM74TmCUn+vKZ5wsT/Ohmk/BoZD3qu0q7UhoxHD8mtD6sRtsYeu0kCLqm
O91XEWnJTxluUp7GgpXa3ujOdwOpaWd6lhe30F3SCVdcEFeYfyJPDpQsh10ft/oy
3eH+HEuUwkkedSn5jr90g8w4JT12L4pp55Y6F4PV8hmyVLbf9MnLFackMpTMevaj
gRxoCfRQ3udtOU9Rb/zn8/FdUP3+BKnJhMwKDs95aCbO/8sK1BlyvZ9mBuOT2H3a
Qr2fdN+o/0qDqpVat2JsTOzHrhltBiZrLy4A1epF2wuPwpv6WMyHON/b94Lu7idL
fj32qhoKyVVd4lsMCTNsDQ5Q/v+cGNBPzS/56g2emLQR/pWsCHW8oorngNELViKc
h1SkbkDkcQW96Ucx1Ny0/vCPprWNBJ7X+EX3/5NuXGnWEAo5ThXJi6V0syr5UDVb
a4kdgqbPTuWi6Ddb4K1tet9/xj6hjDXVrupHigQj5s+fai5c6V1HO8eW3QW4H+0Y
ugAzIWTAMXvPOmi/vBYJdtOIc6pN+IEx4ZVbnHiNwGe9/5+h0uNBa+tVfEeOl8Z0
W1BqjDMnnI0fiplImmnzVv4lPJrp3NQKCH2yDI8va2dKp1vyA7mEot1jhaxTGxX/
1m5qWKDTE0rJ+Z1ka5xm6WZiXJFMdIG4dBpGLUkgV55ERzMBMC9mqrBC4AzNQ+ez
H8ksrAm+9OORG3tcTN8MpRsgzCFnJpByxv2v7xWBlWVhEw6UgCL1jxSn3CNv2+Gx
F3ILX+EzLg/TN8f6Ny6TSIjB1mDBbsh2+xYKgzFzO3kf+H3tK/n+l8rBEeg1UoLA
rVGBUF5wAoinR17f/XlYIjGaNpCMrfBEM4HBk7DBfG3DgKGi73SjVBbMl7qH4jCj
E58Cw2QZHwGUOUFpA5+LDsTznNpoaBnfP3zFZsEg4reVg9+u8sulhGhQw/n96DTL
Z6GAld+MUHx5CxbYtEtjL6U0VLSHSHf1ZIKr0jVWNg2Buv5o3GmvmsHBkn5mYLHi
++Q8VjUUnNx2+EE7Mfd4YQWKsxymdBaRvf7uVZyKKxn0f3qgXj4pqlsMsI1/F7hj
1fzsicWfiV7HUdyQLhJpGykUaJ8rCk6iXcJsourPj1ieHT71/PlzNab3S+PVZE/c
4k0RZnjEjLJit+H88i+dL2XeNiApN/9wWbgukbiYfNU8CCp7Uktd5xXIhNVXpWjG
hjpe8fxB/k8VTL+6UKvtzTndh4eQeWcH9FiPbInrdyrgujjAm3wZLK6pSM2ArTkp
nTJddUaRkcWSEa2SxoPkkAev1IGG6BBFuVw1muAGcXqO3dN/wfpegQ4z9d4nWllE
oL9Oos9t+LIFXP8F/NTZ/G/IlyR5ePscNmUoGtTrjjlCI/zMGdy98G3UXEYKA/dP
dekGJUON3e5/MB9kpda8MuB6N/NvmxAT3hpKBwRCgBV2fmcpHLv6GM1dA3BzF6cB
t7dCPfK5lO/yWqCltOqT0SDDdjuMTq5HiHEusDJ56G6wAb8yUNRasW6VJPUQqDYB
sPzhuAddgQ8tJvpDTFZ4QVl4bz9I7DPuRKYLQ4GezvlPUMeR/xtqrTPy5NRTms+l
ji3nEH8CtaG8Kavf78VEq2NWZxidjUqIH1Nq1EPz0hxRJ/YcXqGhjnRk0bneY8US
QA8fz6w2nQWVcV/cKzF8gi0ZZ0apWEkk7+jyK6STPpjSibMZMOQcSuqrizWgA1h+
DUSaZ/4VNhkDbOImd/lDC5Qdns4fyQXC16aHvPk1h705p6KXPC/+BUds5OZQ0Zv9
rRhuwHsbIBCQB2HLyJGENoBYqrXUTkZA3gQUhqXS2Zd093LuA5DJ8uCHemCjiksK
RKAbElwCW6Bg5RwvakYjUcW55BdA3N8ht4hdtw10LbfVMDz4wkSjYh99uJg+jV7c
vgoKh07u4TpwOG8X1cFvGw==
`protect END_PROTECTED
