`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzWKv9EavYYnx9ByT/NH9Zj/hTn2onVpfD+DsnmqbLR5rgzfBGzEOOb3u8KeBUJx
KDJHnI2MwBftL9n8QHIftU/yhsIbHLx2TJEf4cIOtIXU40EKLYmWl+CAupayBLmN
PvtPku6Roav/YFydn9NxBrwI2dY/l7NeWh2oSwETSW0idwvaWVL84XRzXkV/8wk/
u8Qx9BUSL2R8oyg9Jnfn54ZhEdNhfwQcx87a1XwmEq9JpzejNoYbRLHwlDCKm0ZG
SmrXkERL8W/VcxMOW65IT5gv76azC8zYdx0Ajaf2st6KAH0HfOaKoWEKdGMo5tdk
mmuFtL9O8wN7eARwdYW2t7BYQQLa3KHsyTQ5unZpxM9xcIudD3TmERWk2KIB2RCV
RGnjmXc/X3xmgfD/9aiYJj00kLV2nCreoVDjwd32VrBDvmXZgPTmK3UIe6eaHwIW
VfsJTRIn3hV/rs6vAZvIhDCYUFfhEJMcA6p+DHp21bYGbr6g0YZNrgcp7Q6ZGNvC
RhzNsNRc47D9gBnwmiEOjtSjh/VPhzeuR+ghJxRfBtli7cyB2lRLt7Yo0IQeYSuw
`protect END_PROTECTED
