`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70g7atWXMtdbeJYlxSPcrbrUB1GLO+srFU+N1sO4Z9vfxfqZ464/tFp+hjSlWJ6+
y9j3QCfcI6kTOaXInyKNVB1wM43SdnffeQJEjG2Q6pxBmRGGHjwVX19hyiys+jet
i2Z8xcDZjVPYth/lo2vv6iJVwzhA9Zc/t0enj/5eLh8xyka6hES3bzsezJgpYqJO
6r5MXwmRRNT8uFgGZ1SJj/Dn1iFFvP+ddgh990B0MEJ64X9Zj/TmOSAQU7uTe5pD
5MtZve5zC+PUTA48tXDh398IHZYhlNj9f2xpSqHMVdxP9yeUB/FvGllLxnng1975
83bUGy7MV5tZ0c0iwBCcs/Wvu4QNQX3wyfL0ePth8bTLI0QYlbikOpTIQyXkMMBq
7p6jQQtT9fKlE955XDddWsnCVjEFa7i/njl99Javg/uslLZddeT/YNm0+FrDcRwz
APDwhsYSDewSGfT2giYtJq8lL1PKrohEmU+uI1NJjfp9OFqy7NAoRtmviBinRZFM
ey9z0ngWEMHVbaZffn6suprrA9vYvyps9MdcYTfgrojGICJKLeDJsNSV/loMwEdC
zRBvR2n8GlyDn3+JGJoYVZbsXN/skO3A+YFmkDd7xNdpoLVU5Ts3mwaTBwGmdcRR
EH1F8zFxUk5xtJIUI7jjHe2CYcYgKYe4M+ZStKKz4LLXBwvHC805XzuiMI0Mno8l
jAovtY3VXr5q7UFTbf1sgftvpUtIY32pCX0blYWY5SA++j7iiPGHwynyPgn4tsBW
w76H7sWUieM3g5KsW5jepoSa66jubE5l3s0ejf55S8REhHk3yzOCXlZLf2zCJHGI
AIwpm+ztqViZsTb8J1yRpVfdAunVG1XVoI57RuXCVXwFzKJTwlRmBjJSqrUnOYdV
0GRXl9FK9fafLGVyWrADe9fhCsVkj/yaEDG7azor9Kxx/7+m5fLOPweNN9GXFTnQ
zUBSRd4dv+RU78QlSViR8kVVehPruUCe5+GLgqOJnwZ7vHap5dNTtNy6plLtXt5s
OPUcGRkmg/ziRh8j9mwOOzAqXsCxJThGDTQuRNUz9RuWhzymBbi9GsIccSa1uX9d
PhG1nm9XBs6eSUGjdOtah9nXS4QMgY8feYd7edNxPgK5doBZl89JFbLlgTJzei1k
zPMum5uKy/gcWYrMCOv3hdDYeCYrWj3mzH4CtB8s6WBES0qLoi+MlsVPyPwRYXal
1JPv+h/2XpR6/CbSPjoQzv2NzrLxtlGw6kVjEezUwt76iVJRm5EpWKtrsmmmMSxU
fh4DHOyDaSKsIKswxZ0Dxi7rasiYDxa0OLFTXNL4+Ww0kTfEPcacWbYDvk5LtzwW
USmvw3sV8yfTLjcqXMH4s50gOoj7WVpsGDcdG4qPO9S7HzNh0zANnve+YVoWAU3x
tnJDE+3ZCB387zO1TdUJHNb6AQNVlKPtH4CwGy1951eHFRD1Rad3BmEIwNuANJ/c
12k5IyZFIskEtUb4CvIfTY+zkiQRogURZ1tgkkvIcfysab0b/v6huWCy974LhkTG
CwJ/3v3/yAXxeQSjucLk/o8TbdjB6PnwHbb9cNQSuVQvByc61bT9QYxODP4vKfqY
AdJIJhdBXnF9lScp1R8jdls9FSwHpdoYvJGbxkKQUTxX44uhy5gPqAFWvsRAfqb/
ZNs+tBB7NzoqZ8J2rEw0P5UXFNHXISCacK2IQus48JPm97wp4LJsjQYnVq8iJ7X8
+SnMbCsa2VJq6PW9u2o6OQ6w/JmaMqdN2q/06ReZSZwmPr/sxzc/AdKM6HPlCoc4
ivpba9LH+DgdBkrtQkMQiqKes7DhdT/L7U4/6UDeErNyET2IF2GP2fEE3HYBS04h
eGDmD1aWBQCCuCIv74lNg4S/dAMuFNm9jy0FmtZ2ZVJa1eb5A32mPYgmPvzOF4rn
xDzvMzOa3YfnlUsE9zmGF1/IVEjnJRyluAfhEZI2D5FM6/+kQ+5wV1yaiQvhXIAy
aFwzlYtrGKONcw4fQTN0sOc41UhoWfGAeBKjGqVhqNygbrxceqXjWKl8thWBBBXm
MO6TJJy8zE1Pu7i2zQuX87exx4AbeyCsHCVbNbPwQZuNa3MJJGY8gGS9AWzpsDfb
`protect END_PROTECTED
