`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zvUASW97rR09ipOMT7VUT7Wn4YV/RXNtjIimkG5sHLr91zWMhGDP4YUdxnoQU8kY
HUjNZvaRdXli4fjx4TKxaLZPRjA4BzSckAPGphdSH0YJuuuKYSCsDzIQmPAwhp8z
m8Qv4YFTb4b4/kyn/b7JW2RvBoKCd5tuykkOkhq9ScfkooEiEqLvWh+i+S6qp4PV
eysdy9DElnEhWWnSX0CUn6dX9M9y22XxEOcENJ0l8cwOVjIoyX7aMVJX+NAa0pL8
HGVCDj3yW0sLmZamlvBSvb86r6BbNjnfYY0oEIdjIIxuU0Zo4XxbRoiIgc1/AjJO
/gQGh4PPMCQ7AhWLSqJBPUELju0HZJHPLUkDVqBvI7i9o4BG6id///YXJiafumDF
+ArN2g3vVxL59y+7PJUy8WKJfQPBTZ9rF6XDn1Q3bgqz/CGv19QBeAzdGKqXBSqV
MFPNP+9ajn4Au+9fbAb7nM61z7cfk+j5vi33c1mDs6rWrcn6ztgcHK4yVSX9i8iw
tjetlQmqU7lYEFBeurhwEDGxhEzVUsu9O/gy86jLiEbnk4WPrT+AWzT77N/gDOv1
lgrCi8I0YKE7iZwJCxu0cRQ9ulhpuOcKo3nfcXYnuEB8TVd1hsEbMIjguU8mCcPY
TJ3T2A4mQHvOD6MBjURrYjPjAw47t5aFAxabJXNqSqhtoDkMlOqTT6TwCwvgXbIP
HGjkvZaZvFOtaECMYwPcWPhsveqRBV+dYMr4xmYjbcaAYmdZVFe53azGZzprmfhA
tmsuLy5rMcLwWqRfUiwqitY8nFfsJt4MG49FocieTw5tZQYAQZSH4XNd6u5RvlwG
Dl2pBz1s8su5LpyJNDayJdd3ByIOzPPUXHbMPo4CTEY=
`protect END_PROTECTED
