`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEH0OWoK4vtmEv/NsDDFZLTVDxWQijjEJgimRTwqeosal2OXLyNcFrCye/rXTkkt
GY8ruuEcOWM77GLyOzzVWDEMhAkuSzJi3UVO09HbOh079QWedmql5zsNo3UniKzt
beyxmqGQWY2xAO/GIgSQul7Hnaj+YRvHEN62DS9FZzcQu22qT0VbcQk5SxGSyPbV
I1kGisxunCeDELPraWJxtrJ7e3Sk6NETaUhnEORxnCmFXBs3HWztSaCHuuUsRhpE
/zQzr7ukiT/2TkL3SdSx+aR9ao1jONjANUCyLMWe0hMwFSJeYfFQOd3/gbPp0VcL
VmpwkKSKIw/HjiU/8daN2qZkydTmNXmvizzxAiYtG2GfahfaIQ4duCsXo7WUA7jy
`protect END_PROTECTED
