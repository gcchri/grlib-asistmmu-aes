`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmnaZV1392D0qDUt3Oai+Lai4wwiTlr0nnWndnWGtPtx8RhrXuQWvvG3pnk1GGSr
mwplQminUnOOkELZEKr4roxrrkdEz1aq8DCWSXeBW6XWN4xbaSJgmUx2Zg2gdktE
u9oESuXGB6OEFWnWP/uX9CWenX18aFJrS2Cx6ig5X/2zmNfyDV+v+i22aUI15WDT
7oahDrUNY1iaYRBu0ADMwPj+ag110j5wIJxVZ+2hv+e8MIT8on+n4l0HOpPuW9ww
4v2egjRiyDVb7E3IsGvutYsT7yia7lNfAdTCFH7MAeb8vEntvPz1szvDskaFheNI
JeSWHTqaf8jtrzCzyQlSrRY2vMzuZ31p2nH2xBiISGiRion5hyjA11r/nRz6h4L6
XZ3aWp1sMfWOZUnbw2zA6HPj+8mxMeLkXJwNkvbZGL0cqchV8L9SsBLdH+utcfel
a2lwNICSuIVkBh9TBhv1XTixb7DFskUFr2TzKyru7Y0rQVfDWFtT0GuSC4Zoh4Hl
8RF8vbcxY1AK+Jg3Cieok2tYFz79HdKJu53RcT9LB17JEwoGnUr8V56hIHl0+2re
iV8PHcfEycTcxDOuJMUZB/XhBeelkDja4b7k07LueLG4YfUSuZw7TR5ZnTG9846W
5e4ZhtFZtFR3Mv7oWn9pSOwd/goyJ6wZ2ZukCOubFqocnPioxrqcUqFH/i52d+Mo
megXU5m0sbngHl5kb8SqMwR/QCIjHeMjdNaBCLjh+FhFqGFhkBkLKgnVNpV594Yk
rNA5UHl7LG94xKP9Aysy2etLJ4cpUdhRcaZTkzK98y/Rvl3r8jVirpKtu8rzLH2B
W7rUFlamDqPF+JYVzUGHGxHgVZN3kG2eXDcKSu6ALfYw4xAFjqkGYiizpzAhvSSS
XWj1S3bYhlknr3i3jejQ2kHYGKnVsbZaqKgzSuqtShsJyLS1wthgkMtu0m1UL2QL
rSH4mxs9PWs+4DpoXL+mtL3tLNHW44bAFLAL+IkjJH1OnQ+E8KaZAomOVfpel3nF
`protect END_PROTECTED
