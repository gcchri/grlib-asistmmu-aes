`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yJcos0g4mxOqjj+HEdlX8xmmhzumC99ryxGHixo95o4RI9uDUOtK+mvsRdBNW51N
5NXYaRL9JY91KpQmHhLFv4pAg5erAwvAzbXbhkXRLmBNZseZbZSOzdCdeT3TSF39
7e3K1XYj+HISXmh8dnEK0YlfXQay2A38pXybnP+o9SI93e1g1CsLZlUwPWl9vIQC
HMOMvMFpLbDwx4mrRmqh26ee4w0Jqtta32HcpFdVawmIk9qzCgO0AF4PNu3qUfb0
Um0YPJLnUj7RRwk6xCB/csifvRliOckFdyTJJeUVcmL5uDB72DVOIUfrFsrieMr8
BNZrp4nk1U3COxnfeRJIX/OkUv63wpP1DixbotGUpJQz4sCvWSbMPi5OgfxWR9Hv
`protect END_PROTECTED
