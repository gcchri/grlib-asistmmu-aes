`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8TQCUbPRw0PPQDnoNFA1zVGRc9H3bT5S2awa3hODmv6fjgHYmm7NZVr9vGBjpdR
f2hthsHhzDZpA4JYVjnDokk9tGNeCL4D0/U8tMySpFk21FuxYgUp0ZwBNTDRY0XJ
AaD4HcRyZFX7P8rVKs70nNF8oxw0TmFCVWk3NjZ10x7ssOhY+w6O74uUv/vicqRo
nOyo8fFUkXHeWmTe0eIq3u0SzSMPLSBM/b+/TZqIVGWtOp75TY+9tmbQYBYnhWdn
+1FIje5QEcE1k3RTLtKLDUgLtRparOdAakuqje4dMKgh2Lv0HwzwZIQywAbACW/c
erPtFkPDVxo734YQV/gu2cnCfZyRlX92qIdbih4Ir1cGLskZ7TX1q2o5iQ/4W3ui
d+ZEaf0SNWTNgVT0OdUQETker44SQvpDDCeR550HobM=
`protect END_PROTECTED
