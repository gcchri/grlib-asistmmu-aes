`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ylo+ypFKHJCATL+TpKO9KZ78D4uJXVyVd9T3PZd0FD3z7/CH94FG1SH99g0h2AiP
GOry3W/ovHK+Nw4+2cscaqz/eKYHJhmsPz1EkjmCQsQtcccP/BirkHQnVMSckrEQ
pEcAVqZwmSM1L9Ru6RFN231wtPGt2M8gI3R9Fhsn791pDIJx6r+itXlA5C2O0Ej4
yEAoqZL3goXx3sr9UUY/G1TlSL1eC+KB48XL3K4ozT2ETc7QaUq3JGRPulSuOJ4o
6bs3t2SIPe7y80cEf3WWXp27q0TjmzauOL04SKdGG/deruZMVUqwYangNgNTreM/
P12a+SPgrisBrCsPXXQlkKSLPsWPH/5iESqwmu0qPhdzGrTJoXr7eXybHxbePImj
+EgKPCumTmUCdIuSgxaLxLn1OhSGTVlA2+IE02ixMBvew72buQg6cIxajyurHh3d
8o03AoIeqyTl0Ugcvh3Kpu0Mg6Z6ukdkWVJSi3kruuZcxYmL2iCzSlBO/zQHQgb5
1MGESCDCQVx33dty2JVOS+tgb3WcS1EmLt0qs/831RGZoI4B2SLvlBd70mA/s2i7
1LrtWh1wZnG/UnP024x3loW0YOOXgB0zcQMHqqS3qsQVzyiGyzrapU3IM//1ljyC
pP+7VCeiyNq6iP30X0hDR3e7gkVGswLucrYt+y7fafomkF6EbyNA6UcPDXhO6KEQ
IAqCCAq1z4C5rN5d3faR0FM5WLV+XQOa8PdpwBuIpGiDL0zs29Wk5wSQZld1nFi+
f9r2+Pe6FLsx3iDPwQamoliNWicsis5n3YKPz7oiINcNwsnipkeHto9KOTnA6Q59
giaEguWx+fNvQB+EeoHZRcVaMr2rJQTH6fmpWPYowH7fgOvks1VfELNt2kLjmAq4
gdPtNDndJlRqyC/StZc9FegXMSrAvInrIe1J7qkWSxqBbS/Kw+dRhHOugZ5JrcHv
gZhtM31nqw08/iVlsM9JNHWVrqyefxXmKViKBSD56w+9hlDdO0JrzxobbBpM893R
QmKSFwPoxn06ryPgTb1aOzjRO7Dhlr2e/dUZd2VSNCyI8ccwZAobB/uByCj0S2I3
Pdo3kHjOQwG1RupTPgCzQz6d2XulY48U1B/IthXJafTpEeNM39K3i6azM0odsyzq
Cu2mag+khvoQIxOSBfPc4AXZX2A7RPe19FQTuOD5zEsYVZUMvLYZSA97c/31mapn
RHHpOObbQ3QrMFn1SH6biiH3LCAfr5MOdy7GJ9MLczLTNZUz2eZB5/Cc3eGy2kHq
PIv1GzIZIv4tl8soKS0uHBr77d3HSdkIy1KoHpATpQWvVgk8VbNiFmYwpxwEYFzP
jMkKsvsKtHYYxKjd2LtZibIDAkxXddazKqU+nrmGh2+DvR+U9MNTgSRGP2BN86lS
dXxkiSvhWoBxx35aQqI/x4VdvDg3V97dqMoD8nIidPSZDZU24zuH4E+j15D2JUQX
B7vq6cqaTkPfiFJ8JCnxBTVMK/uQe3fWyOEQK8hcISGkiWUIf5J8zKKCLeY7Ys+i
pVam7nCe3fG+sRnnlMNhljj8Nfe24bpHsKif+5XJQn3AgdK+zu86whd7BcMfuWqN
vq6m8RtuePwn6oYL3Ixcywz2D/yAba7TtpLp2k7omiofJGHfeDNuzrbU5hBqZ9lI
dTOzXjp5jLXZkXDL7lIJenyenDGThTAmVrY0Ie42yKr7kxc6LHJ69W5+vw5WMlta
VhghXg4/aDyg6Cq5AF5YaJ4OnFLlmk0HUf7fQUAJgHanoRRcUxrzZ08Zw6+wZblp
Uasnnfa/1P+k0mSsQGcOr6PQvg01KjIoGibonuZplqS5FyGJUmnRp0EcW1PuBOEW
orHBngzTQ9Z54JkwwKK9Iqx7+WEZ71ZVLvI3q05FKlpP8O13QT2qlb2WkQpVurdx
inNIZvTfvfDEdcXNl4NL2rCUnnLJ729qSnAKi72ihiDGEg/QxpnykcUYtaNvvlDY
G1mmBR536rfmzS68EbuU01ujYWxhCDmpOLQa4I8r9gMgsoCg+NHRmAzvwvAt9M8f
`protect END_PROTECTED
