`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bjJoyDAGgG2tsWKK308KJx4RKWRmi4tRjkV1+VcUu1yf03y/T74fSrjArteVA7sy
pWl+bn7L6WMPetNvDHXKHxatHmIyK73voleCsTxLZlVuJZj0waP7CHORogkiGArW
2dTbOj1Fvev3C7UrszMzTWSeas90O0+hup3ekyjkIzO/JW00qW7fzJ7ENhuYJxzl
+EQ6hDHyR7Ne6P/q8kthD7SJZk/Z/lP8XdKIB9vkvgG9xA4i3KCWmWPKaFP8ufiu
7f864Lmkhmqj+cCisWpnL1rzomppY/wNDsAWEalH76M1uWR6wMmBHlUksi1qPxmi
QfdZYiHwd4QVqXPoLf31wrCoI1LeFQRJN3WHApna4dyTuy2LZWQhmLC/k7qjKTnj
n4jwNxbcuE4tFhFLip5a4MVPX4hgips20mqLS3lL1l64q+AEGp1pDuIVUa3x6z/P
lFYjeiCnWi8k7fmJkBlZTx6c1C60Lna18Ru+Q1/SjVJQmx4daoFcftuPZ/XW6ql4
JRd1FxmAqQ6MOPxxgWB/eL9NneAlkLqKYJokOhYj8rEJroYHQrCN/S+VxxWeLFXM
J0MMJDIgv1MBxZ6n7moRm6rCQND6L9vfZewsAiLlW6bMdmRVx/H4uV4aLnBdkkU7
sUMWIJv4X8DBhPs42UeD0QfvFK/aGD4oAYdXm3Vg03YUpK0wi7/skX6s7tM3zUzY
Edq+4AFtPcgpfc4Rtw50ONuN5YXykoQmYY3KZ2/UcElN7E0C7CVdaUBaf6LO2ex/
6c8eU1MIq5IPoeP/V1zkWDqYTS1+hOA6Pi8oibNDwWa6WXnspMD7Ixb13ItE5nBb
EZ0qqDZrHaL7l3qQiDACsQSydooSLDlR5H/Rdujrx/Z+RI6Mdn3xspDlXd+juwCg
`protect END_PROTECTED
