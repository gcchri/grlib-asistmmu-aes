`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8rROQaxIgSDebp9JL/XkmbyjJZGzfxYIz4m4B4eegAKLujfS2uW+EwUrbSXkzVe
31NCak4EQ1hP/1Hfx0Y10BjVJGoPVpic/2xocAdXirDTMsLDv1ib5riwvCdyLERI
abtYixRj0c4PNBDyfQAotxWgpQrNitZFM1TTEw3WomJrWRZ57f697M+BIEY/N86e
oXVfZrhQsI3bMjTT2RSOy+nE9hW+XRyj/msuf5AQkzUtk32p3TdfZLErBz9KblD/
Bgmmjeh/4DQPEB1Mx/4tpwQpTgZJB5VuFUZHn5IHoxU3w+2W3srH1JhxsvGmCIKN
/1TFMEW7isKdfl4+kS1UeXjTe1Ofj7yMmMkQV+azBL0KGlCYkYnFxS1pSxx93Guk
7gfAdizBFPkgDo465QW7G8cIgdhtpJ+PqAlwrT6/EX2c07zgwXoknajDhl+e8tJ9
7J4hra3GCNseurwiaepiXz8zhhVhTRvXOFVfg1b02LshciK3hl6vFPp6zqkBDGYx
6i8cRmgcpdWKRDdteuWeUAzrItzIVcqVcIF2ALyn7jrXpxmwJwAB2KQIrhTfOVxF
9UR5RqRx+NeHZYCWlL58snrrHdTbm5473q0iysrBCQbm7jhcaJtihLVBBCkvjRI+
VxjRiSQ1S7Bg7a3dNzaCDml8+sjP1wFr629JusjmB+qHDN6jvUf8QCP01qCQ3h5M
hW04KpgNL04B/LLTAOH1N0ki4rOTdGYunNm0b4+2Q7aiC5yB4cj1eISmuNFFEhtH
qVHCfETePifhEbqK/zG2/XjCkkUQSYMl1ugwUNl7018K5MXuzqwcadlX2OY9dEeA
mJorvEyF49B8wVRAlpXHVux+Hrpaf9qXvkAGfRGNtOun0HO8fBvt7tllC27VtjiP
0wdujh3xPsd8y2VYwSTZx9A6tWGHdE9rX32EZGAGaH4ZesR3lx1kMjXE3Gx9vtkG
`protect END_PROTECTED
