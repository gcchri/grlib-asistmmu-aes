`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NeiZJe89gO4dWqPD+3/qV8miOU0puAcGY0sitwFNRwzKSGihdfLo0tSqXDNhjenU
J/PRrC4F64mHxWLcQkrnG+qCLORc5FGCRQpLGeZQGVoBY4gLl+wDg1Nmjh/1yt3f
7nhJUFq70sHTmH8XZt8j89iwWwoO5i1UciJqY5PWtYgKu3WICjczyOQDVindcqgw
19Y79NoZTm5x2VySUeuIsWCguRyh3QTNxpY806KDYJ98P5GAeSw6X5QKHJj2ydCE
KwLL9DXzVNEFUwvxKUUMqrxcBYUCF6NPqgVlN0Xn1ph/QMveagFeXK0V13JCaQsM
Ap/7Err5pGwwUHm33gi3arM+ikenqxgYQ4y8ciu84DARpswUGTQNZV0Ed5Lz4KYj
JtUR+iiDvF7lyTQtN8UjUrmzd6D15zhC44EQiZlU7aUsG5sHkazyTpbdiaf1Y+mL
SKo8DkSeVWsAi5ER0cK5CK3Vt1sRdb40qhJ8k6YZillP4SuJb+jsI6KhdUOdVRbB
FvKCFWyqnSxajQQHFKzOSuYT7HBl1Va9jAy4CCLyMZXxxQCCcY8PA/B+8QxnsSVI
EkSgWfY4ZrdWw07v6eSv2bLyDBqMG4Am6JtF2qJZHG2eYXEJT/NPC3mq/nKdtsmm
SMRqutTGYs47rUbFPJTFIBaE715GR6ahL1ZloxxYQTvBi+Sz15shyBkEe3/wW1x6
eI6dAd5+u7KkKru/1uEIhbqSBGQHTyi3TJa+TQaLP3GKd/kMorDXqpyH6TglPsh6
VqXhrBa/eeSSxBEO+Ut1RdZIP/A9GT5PjXgcZnfuzKI3dz0ImNKcro0COvepUKcQ
vyei6EdzyvCe5zihelFByXPfKIRChxlPmiMeYfuDCVJtwB5cBRFx3dJI14ovCiHG
wOySo8T+qTOdu6kxoHXyiHGxYhhrBWK0XWqMIOn7uxe49f+l5ey72RN+SbXvQouM
9k2L4XMUm96XSTVdchyxB5bE6w60P7Jlb5eJPEBPn8cD8ADyFLE/gNlMZs3ffGyN
Xl2c2cpsfc4rDJ6K4Ffj3KsHJ95modBxg1sAiY08lyCBzmEZXNnK8+CsBWus/Jgh
vwoD3NOIUxoU/SjprBGikDMykRc1E1j7Y/OMMa0rYSyO2mvreAJwjPDrfr8WjFDA
Ca+NIImCAIszz1Yq4VhphsWZcTd95ZJRcShYrp8KvKNt2aSjKllMZhI7SKFCBFGv
9gJsrei/CieA3/hSY6Lw2ckVhzr6kViaOW6SJSdv3WQXy5pLzO3Mw5LZiecCvoUM
6L/1vG8f61zDx07ugGT9RzNbTnhpyXREzEJoxbnBDRE6DKI5BUqDH3PdsSBTvODF
aQFdmgxDfiLnIlHXegZSJbvSJMJ4GNFjBQ2eqVfkU/aqlNUap6rskri6D8sBvGe7
tuGLgMHw5ydsZvROyG6VDVt2LSCemDTyKOQTI9v0Z7o7I83eggXrl+pecJcKCVEY
eKYgOiBccF54uUT14S8cEAEgqdiSfPNYSMefdObGa697GoORyvuwMoUqPcJyH4Ae
R+D1FfK4EquZDEo3jfGhJWfSLTFleK41j2nqmx1tYx4/zd10TdHXchrNpA4ML/g+
1HNyamd+neNIF6wGvHZgG+b+8zDag2zfYN5TTQQh1y6d1bif+FcCZKApjOxaN4QT
GiodxjfBxRj9oMdv20LRDZOuhw1ZsC530+buWqquc9insiaTYzSBRAO62wm8fjKp
TF0FqZuKyvBPNzIfVsaITZ5RxN070PvdPAor8YtRUhXiSI1pW5ebbHQLjfcHP3oK
fGnFfVyrPJGQxV8SsbBI28Xo+zQtzXC52uTsztcB33b9i653RcfnMhsu7wKiWBqX
2SxZnbC+veeWaC8PMKCKpvjngCgRWt3atB7OqdABBDdqI6TUkvkOk6uLXBu1oxd+
BIHfaj/eX21oPIdka0DzQGnpNFykiaaCCmqicKDJ7QjY3ApfgpP87aLkDSQVsncR
N9DWND1jOXv+IN19k66kx1WiIJP7PRX4ClTczJQBWv/RlNM1rbgW6C5s0HFoY+SW
EtZG3PpiLShjCiqlZ39M9ey7TYvlR8iCz8WSHmKGQ6aNLVpOBTfjeAVoEaKDYnZG
`protect END_PROTECTED
