`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4hUMeMfJqQE1OnI670bRmoNeOJ+xk+04ws+UAMydsykjBXM0lAcdYfsHJOUhm5g
zZCDgVh3nJp2FYVHOGPMuCEV+Bz4q9d0lQ9PV7Lm/DpioobLfnYg1TkXw60yyTeF
RYx5wZAymOJVvO7lq8KUpBnC2LUxUTmnBkQTrPa3JRAqLgyHF3klut5nMuKmc5XJ
BuQbs7Rk2FAN0y6+f7ufeW6icz1ralZVdGqjr/YDLs4kF3wGi48x8iq3ixPdSeJm
fdsu32hZBYc/o9GQ+YLeYwFQTL1NsbdaUkmeacVTsPmnk6tpJ30ks9VD2HLQYGFe
TDuuvLfY/HQXpqKRQ4BEysiPgc9rJ9Wt+eoSv+8UZJkPwA+ECr7wniDqX+bXhM1R
/LoLWq/1+v/WPy2UPvHnB2g4uVvhy06De7fuWwjGete8jgrLUu9DNyiPhipyO1+2
mlqG3Iq9U7XaPeFd7EImudtkL+v4TBKXO9P8gH887qo=
`protect END_PROTECTED
