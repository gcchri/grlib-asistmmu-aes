`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aSAXAgWRQQGZo+gM2T5Pb4Xhs7oK7sF7ekX/PgLsQg5soccu94W026dlKcYfzxSg
Pc7mEoOzE2JoQlL/ExOGAtJfHQ6EUdIMtGvC+Gox4ROwCENpK+55YbzzlhksmUS4
0+4hTatGw42LDn8kY48qDT6GH9pGPN0DMsw26RVKC5/ukAHyrQgezZqqbcDLwoHx
FtIUUgqO0NOHWnHawkBaG4kYsDHGdZYxIPaasjsKosytxw5orHYnswsQD90lvtP/
xTQDeBmY1iOgJGwFrtDWFUDBWDlDRax4hrWWrwByviBJ0fzwJbTD0KdAtrn0s5Bz
ULZD/SDDuAEM3zPhpq0EW8fzH26c/HNrY31dGqi5cSI709s649kILONe3QmWzhbp
Xc1633X6mSt02bBF/Df4JROX/cYkLBCIuU8XZMFiQwCu9lJFhmSn2M6wjAPihiEY
4k/L+wjzZZqRpb3/Im+LIMOrWqFNoizLe2B5tNtnLBfFQZNc0/WeFBLmR0UqMlfM
hS8bxCHpN8G8Q7pSE5cOCdb0Bna95QcGCf2O80tntPz6gLXA/WdYKApBIJ9bskuC
E9yuj9w+LrA5ykUaEGLW/bRbWNRHTdbC8z+yXgbDGu1OUElqy6+EUrEszfwBxEQt
Xaw7A0jQRkQYzXqsMcmwczxE7vnU6CRYrhIwJ74XMYqx9a4XuYkUWuESz50M/cAN
5/IiygauulbR4iyTDu0eIDgamIJMvUnkRqGjPPd31DM0nsJxEKWTu5FFcF74Dt2z
MYqZx9awbiQ11yUusT6LUCjtPJNhSkXSzc0rjgjVu68jZeAf2PodsfMeUr2VhDy1
3jmVTV6qMk/gUy5qajv7edg/WBFkm4VJk68upWx5xuE=
`protect END_PROTECTED
