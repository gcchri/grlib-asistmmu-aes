`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4s4jx3vq84vffP+1os7BzJgADo+hq8G892Pl+FXOkDu87IPRlQ0JepoAihxBYGMT
I8tS0RNZbbRZTCa6jMHc0BEFYDKXU3DA1xr3o/A4bJUPjuqC9UrtH7CFFFU+YJTO
CMsVHxhLWiGq6BDyP263+DBOMDn9oety18FAXhUOjkjioi9stthAF2Iz20PApStL
Ed109R3NOGPi1DTO05cR4opHIRS4tFssYH5LIBEqxmuGzD9NTgqryggF/MWIbjgd
Lp/5AKIJvBxYxcOVje8LfWgKnp/fwNLHYsNAzRafPM24S4vG+G1K6tQq6Ldi447a
8R2X6/qHZlTtytFm4hyj7xuUVRQ8D+2htVJxRuFfopa4czFhp0jEuhFHcF+dX1YU
UlpHv7v3zNVaBTauFXh3h2gJuqp0emGpcg2uYgaFb8TkpNRbtLyQQCsnEy4iQ+pB
2WnK+7xASwBiaxL/D4IvFBTNUkyEwy/liI39Npf7UOewnnA+F4L7ny1IyVetH0Xq
TIC/emidbuWbcbOx+8Tdy45JJfxak2qy5dl71KcoGEx56FUvM7V21wbI+OAihG5i
iXyrGGhLi380ZPlU+Qw7BrCYDQ6sHgoDRt84ORBEYOWUfhJaQdsxz0HY2DFISOAf
098aOuLKlZd0SBL4H85xAgY2D1Ubh1Vx7t7vxwrBuOZYChXfxn6eNQyZ4de65qx5
IN8CCXNtVRiJPw5wQjcYP7LH71aReGg4K1r4BuvCw/1OPnqHZQwCK1EMxSrDVsHz
/sf1Ll2nEGGwWISW7itniUH/cSOOQgnxiNoSb6156BXLzlyfB58NJBbVEv1iek9X
2VqRRz+1kLbv8hhZijgsp/IhQ4pMZuLpmXuuGVY30VgIj0JZMwQ1JYcsrf26XIw9
Cz1+rt3dVPVlMRmfTb5b2AdXNPgAhlWcZA5Nklzkwy/CZZp8jkQju1F/HikOBXCp
0LogcX28oHnTS+Bq2JlaTdAFinckE0D8UsG9kslQdTDVHSheUsRPqncjV4QmuOVO
bJ41f8+ju1D24pjrnFiw6ibtjMjBjTpQlKcRvNsivdMAnNxdlvmh+mbdsY6S4FsQ
xytRo+4ZImIsJdgfmcqpx6rMyCgkDUQb0yjffqkpVRGOOmjOALA+PTANPEwlPswk
eQZDGzDW+OXr0IKksCB402aN14nJXRfTsVBmXZ1EZEr5s4iFtUQxZJ0oz5X81j74
rPfPNtl3fd72oGrKlxZaZMNDRhoUJTHAu4oEaMT/BEZrjCQCQLfdi4X7gvC1jzWB
`protect END_PROTECTED
