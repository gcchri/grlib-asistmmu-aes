`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J5JLKtHOIkB73OPrBdoKm7/W5ID7fpBRNx914Rm9k7s3fQepDZxZf1x5AbVp3bCi
of22eFkY6DP7KpTjEmwZ0Xe/oMiP+lSz1X9GpM+U4wMNYJkd3C6XTkOkbxKrFC8R
GBSbyL5M8vezSOFeIkD+g8Tx2MW85atX/3CKojOBf5mnwSFKE+4qc+zs+KKjCOIh
OfzoRxpaNMHFyqYZu5EWeCPQGIjB566wEz+yemyUwSXKrTsDJp8uGHMLSBpjMei7
Duc0KOjaxGwt1r5aVcp2w+yT9j1MJIKoULLZRF3rpMLAnbhKvD3nix9341OkQjSf
bzZKYoYKL7Onto/jmSO08A==
`protect END_PROTECTED
