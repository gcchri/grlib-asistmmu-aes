`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCesHWl/rKC0s33VFJEPcExF2rUZ1o5LAtJR6r3uK1RRh+Vmfz/6Rr2e22n4On0k
G7+H8GF5Y7De9OKLeKGIBo8Cj/tO768WJxzJJfYSTyw1Fx3/8RIkS84MrMJPZiAE
BtiNFXBEorLTzHggh/QyHz46l52wCIR9244QabORiwiY0Sxp6wDHvoyFzYtkg3/P
SKg6nWMiQat3vzuPakEv9aZWN7IPOu2Zvzjj13hMBxGWZnZN8xLg4K4VszAdZMz/
XwZPaT6DMAfFOhPwBYgmP0Y4VOO+XUsj3/VXsKrQL/M=
`protect END_PROTECTED
