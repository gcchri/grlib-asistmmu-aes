`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yVortq69IRRmvccESVE3us0QXfj0fDSJpyD1m2v0bvhmPWfZkX3rVBS+66/4Na56
V1Uhwe9o9YFDymamujjRXzFPPOUfWesJAjHyTqXi6D0Hp9QxoDYPV1p6wt4rgA5U
SuCoV2XL5FZdD/XYe90eGXfJRyVw/zeKBspssY1O4NmfndtSw8AVPEXeuvvDXqQ5
/rPM92wU5SaWe2QKvISs86RqTa0WEKr7P1wY1De+xPMqRR9OyCid/xGZxSSMeMMR
x/Ad4jq4m3qqwSXn7SunGlTF9PVp7xIH3Tuo6zOi2OEvvLa8nxSMHUVzWvUdehFu
WOo5YRr2xc+pSElt5MhhF9WgNQmja60OoQ4t0W1y2jBJ6qK/35QNvYCmf8uJxjmk
gg7OitQTIEPZexaV7nwNOsEvogoYtH+86TGs+KLaBRkogO55tnWuO5PKYKt6Vmg1
76nrCqfyxxz3KzRyRDPBm7W71ZpsJGRk+vs/F9ivFltqzAMKAAiXx2QzhqCIC4hc
yPjtwxRZiu89l9MPwUcuBmiCd6jFCi8+WY4+Jtw/jvITTxUS3Ob3kZWdcsxJozh2
BBwXZ+m4V0jOfLchJpwoDg==
`protect END_PROTECTED
