`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNvjI6D3t9RHkIaGxL/ZI/AFE0seSAhF1ICg9anbFdwFNg0nGRaBMCEOxY+0Icdk
zBPkJHTNugRtWlmSZNNzDedXgMOKE4k92T4+qag3xuWKT/it+gtC2UA15+0B/UAw
YADRODyoUIiCrrwjlWVUs+iesV0ZLmfLtuqZawLcKdGXWVO2in7qupbDRxrQvmZ8
lxGmVAruWL9y7VVupTrQnPXbrL1ILbhCou7+oM447RjMI3nT2th2Qti0jaa0Miri
kHQr+5REuG5Yb8E+tEulw9oTcSRRO6klqje+8NfmDpEMTsCcOQ6JjAJm4C1W90cV
v6z0xs/ci0fcr/2QTaYmEGnzaitSACQ3+vokbOpQbPYqcrhwX7DabG8QJ2DNR4mE
8Lk+HWWoTglye2Nbh/5Yww7BZ5Jm31Pwsa+n4zEe65DOIHCgG84WzUyvPz8DceDa
C/hQyBDN6Zy/T9MOK8hkifyVczVRgVV3uP4iquPCBYGpO5mSBe4XDPjGHcJmid0T
jBtTYXv3IDd8he/BxBzJLjafs3cCpgMNiylSdW69+jHiQVFxWWBEiJGZbOOnSBD4
Dv+VHIwf9xUCu4nqwcSYnTJxhxM0v/uZSsW4hRSU5DB/ZI35AokoBGpUe5elDJid
lFci07gZ4uLCPGWIZnFL9NvWyr/iIuBEH3lGi1cs+fN3LK2fTEWnRexZMQJ2C0+q
6tuTv5Sv8G4LUwVizzI4lg==
`protect END_PROTECTED
