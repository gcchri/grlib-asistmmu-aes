`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wuz9SIursYtuhEopXt4oF6DNDakBJi6uiJrfUvWtlIj7YR8T22DcUFe7n9g3Mk5Y
6N/7S7x7Xy++2ez28sn7NKB4Kc+ahYGGikxT+JBgUMk53pEGjz/NffwoHHfGPGSx
1lLDmLYHEnMWOYsHUkDChkOsUIJMmq93rTpwrbFG8363P26a49fj2jhkuod+Kwic
mtIB01FQvXSR5XzaBtghOTtDVMmnBPvFeFK/mmpvMVa+iKGXb21fTqd/sFXI1rEm
lTksabScRCUHtFII4R4N0CNsbb3ulEadR//dec6+M07Y8BNQkHNgETNMUza+hM8U
`protect END_PROTECTED
