`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vg1VgXmbkTwXuJL351GRP/zFIIs/ftUvxt1R27B7+gOYvhEmUzkN8o+OE+JrnwOn
UPj715pwRJL4i3eBygvp73N/PqbzUDSujOzii9i8sLjv1ataAvBzeX1f6rt6G6Uf
KvqsNpj2F++aYmL0hV1NNwohyPqsPIwLjEwFSij+Alc8xnv1d6S5GBaB9Lq8H9+v
uNRcM1fr+4hQgSqZfPA7SAmdEX37qB2MWHhZbmrTyFRMAPSPDvpCpJHzs62yVo3i
+DD3SuVELMP3664vMLgsCRKR2j017renrfC69HBwPoV2647l+ioVZXl8O7zUPLz7
kXqc/6rK4Z6SYM5rjSVqgq+dRZyA96x4jmHw1bXPBaLTMKuXIVifKE4CyFSoAqjM
mvsFNPxpEFBhoH2fOpRvkwIUgsGGOz6+bOU9LmOIzN4MZp3lbuE0ABLaYvVj++Mz
MqXf84itQceaIFfUC0HXLL+gvJpYvE2OHClHs0OcdXMbd/iRTA1Glj3Cf1pdsjck
0k10+A00Zwdw4d1iJ0YMe9xTSe0LDLmGOpr64jiAB0Sdb4tqlhGgzkMqMtRj9Lvg
eJrCSmeBKxl+kbH0137IEX4CdMrFgZKicR9xHZ8eqnI=
`protect END_PROTECTED
