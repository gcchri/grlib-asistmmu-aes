`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQXnk+5yximx4nmC8t6KUyhlL6cxhaV7xW2fwybiSpEo/z3JDvmKNjH9KI2JhLxL
w6P0dkLIo0QNFq3Agt+rQ9k/H7vvFFGY3bEczVwMBSOfjvX1XqwI/DRu+5qiy4ST
+JDQisLsjE8nqdCTa3wRIK6MpqJfGtT4obG+tZJlmQRnXpbzrJ/ELlyMtJN4C/H7
Ol35BqAv4HacEbQNiwbM8UsXeX/pCZCeFCdn99PRQCJxJnQ7dmKtO7sPOmCx4SUx
KYwkK4/oSRrMKLZDkEf1ID+ljHJm0aMMhl1ZM17/+1cGol+Pls6cqqtSOJ40Tlq2
tUd1FMGsg+EhXZlRFs7VY1untDWPkXiZ7xnQWNlmPqFIRRwFG5MBiVte0YEfk2nK
TdiYPdLhk8YMPOTmP+BLFRGhQjotR2GlBG3eBb8Kclzo3GfJSm5r/01pXEKVIDsC
bmc8EeNL6j7y3FrbRQm1dsaLRUiPlbSmVyjTOLyVjik=
`protect END_PROTECTED
