`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0rVez4s2meEQrne7glbT/HGELzM/xipraRa3R7hcIsNXf/EhAmnbeBMwLvSc5iX
9ezj4/M3REMVya7NSh4EFlxdEYa3MUolKXOLsrGKOVvlq1hptoDR4hjI9ogEjO51
FYGEqgG+TO1y9PaNOhUjapvIWdYPx2LDRejr1OVkE1dlo7fbWIcJxhPSp8r205As
7vAGLpDWytXstqxuBAuuFsII1kfNis5MaEKMr56G256BeYMZo72HH8TOsjZYX+ta
JAg7EIqBLYFN53nQ/3jumZD6SCAgSsXzlaCtXvAlvzswJku3pZ2IuOTmES9zZlp+
OvN0HCxzkTIGpKt84d9vulyr8ABebgMKaETComTYTG0fP5SPLEBfAJZLu+gvFB6e
9igTd2b8EFNly2CGQGh1Vuy0awyQw6/LyFsoMZFhY4M+T0vo3YWVT4XuXQkL14HU
HezizRyPvM90vQSF/ZReEoAZsfVdB71FL9Lza180a+RJ0HP8dQaSVaw9r7HGrZ8m
D2sq7sznjYTbGh3foRINQzn6sH2YaaHw2GJOafJA/PUNEL8L3K4gkbk7fKEZAzAA
oEYrIxysqdtZ3s7iAN9yfkw4TMOXhxaW+HQJX0KYR761hJAVakvidk95UCfM21sm
ea70abWymFYVwqMO4TZuwnMNtL/IA6tCefBxhAd7tQKJqb9eJvSjoLpeAIXpD/vP
93iNavayrT3lSrRdS8RFU/PVeNiFcVN059ORMdQc29fWBVT1IHUiC9416jlNLKFU
jfO2RkDFhuuPIWLJwk3WO2eJXzRJDi51hnVS8WJYeUGcHSRdC2iqrQrZ1bXYSHKI
+0AdUcgGov247DngOvHOWvAf9tUsRlPeMjO7ZueztZ8=
`protect END_PROTECTED
