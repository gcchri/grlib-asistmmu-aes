`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ChMFdN4Uw160rL7T1l50M7Do/nf49OqFFrkHlsNKDlCZpBnriBEXVLBwBzknmH7o
o9vJZO8dl8BDJzaNH9mx3BlRuiCjkLpScY9TR5VSvIlFjlTxs2L0lpJnpKPtOYaa
QPhdU9ElrVHS2NuG0LwrcYWRfpzOwMYu8yy36rqQEAn3dmaXKJ16Ld+iyyXWMEmX
yUhJX75bQfB7KqZeyZiQ91zyJkXrgZpLoPCw2G7uXBCpqtKgWSixoDTLIHNzBtTh
4QPxbSeRnpliBj6QdCi4KoT1u4LDJc01hFW4WTPzYAHvbafwIYzmxHScatTe6RvS
Vt8GuM9pSQic+BuEnzlbaR60QR/tBq6stZVX86/zKE+IR8Zo+ws0J8pT4luvY9dE
UmdENEk0ttRxaCxQFXirmgMBNO6KVMWic3i8bdKl+lyK8nsFKQZGh02Aa/YjU0lT
nhP+O8pov8nLr1veyVTmeMXWazDi0HDg+12mYrlkySUl5j+VKSwuX8rghgmtw8gm
IBpV1cKBwh+8wvLC8+aql3jW1AFq7rQEwptaKVkQZkw8SBeIFHmINwezG20XJVfz
`protect END_PROTECTED
