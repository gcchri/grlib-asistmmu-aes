`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MMl3vvE8SPvIKp7qmtUjGGLQfwHHaaCl9FoWlkrn1vgnXkluUN0l48slfmtODPeD
wTGdcAZYN+7ZEspeV8kYUGq6ZySokSD3gUOwGgorFBLF0h9BoRM+FgCK3SQBTUYX
BUKkICkYk82eR4Ew+Mt6jtTuCz8FmgibmTnJncM+n4z+2vitY0XQcKhvFCjS/l06
QcgUzeUwkqGw12dPRWBL69KTDjfmpHO2dwrqrjt3QF9z3QNlsUX0jq8BlTNnh6CN
wERyu7SEkFJ1ppEHLoEqT+Q0ToQzydL9StaeCALDO49/6OEko/UFuuqDEWiP7bft
NzaTWS2h/J5baAXdCC5U2D/0YJqopLkFyuiyYZ3yyZdsLlDzUuqNkgWx+sgZgzHK
JLtPdDlCsN4MRjTC+B+foYA8zVfrYbrGGeIDyFzxDkWZjV7nEaPav9YJVqOvqBV8
269+uv3xAb6EqjjiUjdA6UuLIZoEN0lrKMlA8Jf3RiuygcGLEYy5PCRgB6mjdbBd
NPPWFQom0EY7YLSD0RJvsTjxKSqq2BYHfau6AGgiAUV84Tzq4cvPFUgj6CZKAvnA
j9ABX4Xw9timHiFJSEVYNYiCFbOrpRULtTZn+XBFo5ZQq/7YTzYgcTzXy25bPJpo
ffGlsbL/opCw3UjrQpTQj2M9MG6ebe335gTQrCv3CGU=
`protect END_PROTECTED
