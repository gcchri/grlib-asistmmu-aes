`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0su1YBc26ixzaoripYbxKUIQqwEBi5f8H+eaiDY5QUijy+FGLsn+NM0mu5ImhwFv
xu023UpJzptu3pyYlxlH1L8mg8tRzX8Ht0dL+J+lnf93rKq0bpwzGdbirDfTN7EZ
u/MY2PhZ0v07X7H+YxB5lhQkyrr1oXyTY3Zzo6GfD9XarMVAR4c+EN0MXwFVfkkO
8YlZh93IEqGoY74RwPh2HHpQmQebFLt/E3UiRVMMVzl92oMT1boURYAv74vLrUEZ
gP48b7k93DXsS2ZG6aP4/XFjRoxcLNjC66LE+/hYsYpUtq2RZqxBWw02fQe0aCZM
7/RzxgNJ4KgGnhusS47CCeKrXEQ6bmqHC4HJcB/wcZwYQUBPKuFLEMe7bhzg3YC6
/h7oomqdEP2Xj14e0O/JRiX6xrTWuhoY1/e452urIaBuQh1OdrxOsiLYR2sQJcqv
Gy/B5fyb4vSAFt2L2n/TCwHXEymoJ/ExO5ecKFljK/rrDismNfZl5znAOCqut0oz
iSd2TcOnqH9Yao9SO5vP3yVYXwu0v5vyAoHM1k0Q++GpxhrykXT9K3iRLdMjEkdb
lUIkvgMeTiJLUFUbDtvBc4VmUoT14lomIi13qOFJ9qHJWQ7tHV6NX0eFTpiGW06o
idDt4+R3FgWnLtS5xNKGlixLHsqHfk3+O5lXZIPvm05Xe/81lrCYGoSoEJ/LdpBd
1+TBNYGThk0+6SEa4D9uJ1/6zCW7ZxP7VqfdqbbEVwwVoTqrdqsKBqL0r3Zcu7hV
XI9G7uaS6ZnQxu7swd+bXg/A3vBKQUzXzVtet587qpeZO/iHxZ/r2uZQ8FZ02drO
kBPuSNyL/q81tPVZHUQ7rjo4NYiqsu4kqeuzXcpuRWS5/TbP8WwUKbySXsEraiNs
3dLl55fgyKguiUPJLl5YMgc6A6JZICpcuV2AssKvQBPbgLerw3bHztvwPKgBKHfI
TyzbiOAYUUhlA/XrzYzXcoWS+gq2AqbpSG05cCmg7LXmhEeqKnNSA3Yi+Qo58Wvb
pT5WGCuGHt91B+hvqb4VituTFOB7CqdwkxfB9nPY5JrdqItdrOjSPzLuRkkdcVS/
xZO/PWGcplaORduQzsP2z90gryby502xAaFk7O4qWT/2743E4BXfZzBtK1EKynFo
b+6zIiiW12VYkl4swsNt4uLtxfVqEdNu/gN04mQESR3qYJd47q8MMYFtrbywWYPs
OTFA6t0bpZlHlaAVcD9fkNdtfTsvkdqtT/4kL7cUBcu4YM4RCMw8CKEY1vvDslkM
9h2m/GFdc8bpJ501VnAZVYbkbCEso3gvG0sPPfxS2a24CGpa2N8KU6l+cy8emUxI
Wd2bTXL5ENWom6SDglHOx8C0/VxpXLbCEgxl+py4xQnj4QeoqHiYsQzDXVcMFinT
ycy74pZDpufTPTEKXI2c4sX26mM1ReUFQArGa5RloVs4JBPJKwr/K4NR5fpRtydD
b48q85JrqxtsxgtCjMSw0B+PtgNGs9KWYVCm7gw3W8qFOrlBEB9654TZUC+r0iRZ
XfDIudtSYfmuBSMc7chcIkHyQyckVOrAMF/KmykjGkO8eKeZtDGHX5ARkGJhNdmE
HR9Bkz0BWRmRB17UHTW5bsApmNdjiIa2LvOSD3ALeGuRcX70fJUlJfs0YLsSjiDZ
NJlOXXOS0nv3ZzlDdR240RWWHPM1WwRDxcHb7Up8NPleBKk3wg2wIw7usrjSAK1D
Jqry1EN+4XKpgXPSfG8jFsBq+R9n3tOU1FQddClQROycMjGNFo+MmyAYmlAVGVZ/
FMDWNoOvJUzb9fpkXJV3ANKE8NRTRuyWK2oHtSmxoNWJl5RsswXCOuhxaotOjSs6
EqX80SHyqodAgoitOMy31UGr4J3V6ZDPelWwpk5PeOYBkOn3RsrGzBaiK2P2hbyn
6KnXATA0mRuh0Dz8joRxfzzd1t1dJruCk6Brm0xxTD2RdREeWRcaJ3SJdpeMoU77
cVDpKDWY/cF2Y2WmdW6ZGOHNCujXLugAxcVBtJ8OJqrOppgQmaX3J7fd1aEA70V2
LL2vjga9D8WHden+rBILqaiFOPZL+I8jqHBTB/FYb8ZKadXeQVY1y8rnGCbHgWZT
WwPMrg+XwZ6RpozrmSKxxKQpkTsrL2QGqKdqbLoxPN4TVx+kE8ukx03zVGRwQN3B
LMVSf+hCYfNhOg17SdEk92VhTglVxvmL67FYAuZN2KzhPfjNAvhC8KLCn6ugGUAn
JKjAKG6rLAAatemxUkBivSyX7KqcfS49SIM81DA60biQsVb0IsUFLjojVVkZpspD
TrxsI/eAG8zgKvoO/ilgwlSLmOpHFGIz3djbCqxrgnEGEtnK3f1uxgyv2xCGQ5p+
j8sQD2Uzb3jhfGTdkpPSuzuWaYu18JdDX4XGur33CtZt0t8qiGjfvAl8rTim1IKc
wMLd673etGI8SjclOgvEJ+Gba1XFBus8KNY5lNni06XQZ3vR8Kumvl8EPMLeqACY
TRIpUvyfWequiU5BaQAS2wZ/XmyHNQ7TKxJUQLlV9b7TsYAqBRi566Vs4Q6nUWGy
/sgh6SEkVOLqtQz9UuXXlNs5nZiyG2lPZOvG9w8RGVDbc/4c6MPapQJoK3RE4vGP
szuO0WRSZTJTB7s+p8mF7tqZ10y9ZlduFmr54NcaQkG5DsNM33/yqs07u5TZVJEH
zCLgJLVdQIvZaSscP5r9Z90Zfd17FaeZjz/iYCHUjTk2bGH8mlMyVZx3shUNJSwg
Hnw4/IGJs3ZAz83KL4nnCsHEBKUUkJ1bYbPGTGnzILMVoJerpnhoTefe4cHsEkB+
WfhwJgEIzSS2iq1kqUVKJ5OX+htkqjfwSVFc81lH6NMfOnd94hrhvSHjm2VwjCxU
KE5twjtfu8IKbGo7Jrd8lx7nvgRZ7dc9BCbsc0/R7t01H4HT9RUGXxEeUbpbpl96
Qv/4b3+Din4yKmFLL0SPuiKWA3+qsHyXN0SjEiyXbNyhOpatMpb1la2+/eQXxpxP
Gt440T4MYAS+idUM5a0HBGqakQ2Glq3FqoIWr1HaoVw+VYBwThXxVsUj/gYgKYT4
vObaDhgNqtsA5RfmG8znjNqVfp3v95td0UGfsgwBJFDyaQMlAE9I+6Zrja+a6m/T
D4A0RZEiCnxr4j4SAZaNl9AnxR5aYkhAFpYZ/fewzahP57k8xi4JjfG81JE3JpXv
4fZ8GuegBtn6mZfbEmZyWfkOTa2ZbDloaZLuVQM/FSzwKeI49m1ZW5hwYpCH+5tt
fUD5EUw/yC4SN5sdhZHB3zhx6/Q61yQvWRa1xqvl6kQb4UUGE50HWxYZZ0jtbv4U
WqPvUpbOs0mo+NbBTzjsGFQymJ6fs8pp1FYwYlJLwUalUM0HOwe/LOvx5k2ZuRN9
aB1981ad6Kisna9+r8PgFUh6bOH8o6fQRnYVjy0dPZQt3YlOsB7dmwJtteNtBGTA
UGSmZ1MmCxZPdBydEjm4wVUT+iAAuxV2sa3emRj+cvo=
`protect END_PROTECTED
