`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e2y4SFv/2gDnFCTH2+MqjepvmUn/RPP79UdDdUAQMnqzXM1EiOE9oOATHo58gTF6
0zbexzekFx4lwlycdZfrWr/xxMNnWWhUlhuNLJe/uJ3/GNlwfa5vn+8loNTmgxx/
ZP3Lb1UH/8QK3bGrgzj1w0Kne/yid/z93YhI+Rl1NPrtvrwuN+23M/9b4m2v0cFN
7l5Fuy5h/5eUpGqZWud96YgxxIE79ZrDxWpCOWXtMVuraef3GNQ4hXA9q2IEQM0/
ehCQUAnIACE2wZui/nQckg==
`protect END_PROTECTED
