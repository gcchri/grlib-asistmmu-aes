`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SssT7C9XCxHBKkbQAZlfQsfMmE0EtJ62QecCz63cEQs8VWhLBCOGVHZVXg8Xkv0M
xQHTaZekJs0a2PpaIcGkhZQi2ydtm4Mh/EowKFTjkNuXUiVr8f4y2+13SaYbfZB7
oBfZ1lDtabG9szJRI/vV5RBLJCE0/57CIev8JghEitdeNWCFmSmaErRZ6AGEZS5X
sxC7oeclnDZbNZS7OsHQPVzbW7DMTKZYmzn0LnH1HsPcE9V3y7ieug2M6MjpNqhI
vWk1k8/j4rPsrXSpnanUl3plIOIwKFBHA9OurQm34QGTvS7wT2rt+FyEzfDSHUWL
XSuzxmNQOer0Hwyh7BNQIWj7Eljn9f1muPT3WpkoKrxkqwughkuhh6d8DpaRIvPn
Nhfcqi+LBHPztbm6wfRbMmuzDmEwmiTRRPTH/b0U6cWH8/CCdQUXRK0NkeehCMGw
Ca50ViARwkPeb8ji5ixCG21/LB9iC+l/PgltGG06EmaMRbJ0V6WbUZMvppeZyBZG
QNgwTc9JLLCLVE68T3P1ssFYWXferB9NzKnm4Vrqwdjqg9c8+KAVuQN8B4OKkfPp
cXmmo4uxvKpwRtTxze2oaQgR4eznlRdpuh5mRIi0PobuQukj8CjbH08km7v4+sYI
qMrVA7O5spG4TD8PoNPAiiHL1E4MwVOEwDRPq3TcNUScyjw52L2AdtYzNZwpEwcu
obvnxPtSPJf/m2ufiDZikiLXrq22LJ030N7Ds2HJfuUdMTerS88RPcJltkD6wGho
6LfKaa+3SPx8k2lknDCI9dmqTCu0v5JW/ktTr9p9OrLM2l/AV6yYeca2u9Ydttqu
QT+DAOtz/D+sdV8jLDe0nzw+tZRdd51/Ecv+Ju5JslZQHNoT0W1Vf8pc1l8woYTH
pJwbbKEgMLi8afLtPVs6la88MXE5mBwbqBDAfgVpopQ5vBpWq9aEKX8VEf7Phw4T
MBTFLpurUa4alnb4Yvanya5rmOpsxJZAuteELBd+HV/P8t8i3HIstHUUl2VE/6GK
yM+vKOUYk7oMH6xutaSfF+zgOq2zmTs1VLuRU+rD2Brlh/FJWR0gdLToQDQTKuch
YQFQJ2CC60pa1LrlagBmUSjmhp773EIdZrFPfXh9HrOuEyDimL7Nfz5cfWLGmPnX
`protect END_PROTECTED
