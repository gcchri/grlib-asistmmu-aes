`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0kyIZTx805gu3HPVxr8W3zQM+LBd2W3TwWEPGvyebSWI0b9BgUCBDyJVay81g9tS
7tuGflsNXNrtrBvolrUZN059T7J4EMliwgHlVklg4tcumv4JJHaEbJLY7OpQoPeU
c/HtO+oopWVrXSa0A+micrGQS2+Ah3x8OQoBPaSIRNchuEMadj/lwlaJXrhHoRCB
NmoxOiknK7XWx6U4JIOUqveGYvwt0DzfiVLi1GKRBNv+lLkEIZ4lJEipPfb5r69i
7SX4r6nwSyVU5RaGGeBN+yqRfvawGhYvgxKjw7amGhqHOtmrGEgF6I/dxzg7zfOA
`protect END_PROTECTED
