`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mbftFjHp1zUUMzA/Xh9YWHdhs65wXr9Uph6FLRkpY2WwVgd6VrPvR63hVD4sJnxf
DOMjTRMEFPzLeuMf4MOdF8Ve2psqAfnGMVtv0T48dVj3iwBvSu7JDxOFiTPsg+G9
6ls7z8CUlkYpaxY443OAKqRk/yILDSMHo27XEneoZ851urJZS0zUia3urujnIaMW
5ZZkLawrHfObhhQJxkMwtTo/yvDWn90bCcIzZPNFC2dhnIlwsJ/LDF2gpGNqwT5F
uQfkwNyIdHfUD999bLvD/Ps2HSxML3GzVHeGziLYtR1S28BtbFwPVpFrlXb+1KSK
a8RiuAcokYxZJmXahNT35w==
`protect END_PROTECTED
