`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hqNHNim7Us3wGx9/E6hJgdhIVlckzcQyL4uYtZHCkKgOazr/N5NY+WpfWKFs8D1B
Pf3oAILLxP6kf/rmV9nPWLYYtE8yaPyem+fjbyj12OaLxuXyhd6mzuTkilG9sP4y
EvavyYPoK0CN4eyxJ2M0R/67Lzq5Pj/qbzyx1S4WVGCFqqA/Wf9hiPvHX4fR5ZyX
JgLz6m6iyrQd6A7UxqmbVN8zDOdW9nbFN4KcOyYHrb8cKcQMF7DMYM7+fg8Z4+de
VvHo4g/F8rwFV8mAUHqsVcwkbKF2cWBMmgAt6nUS1cU=
`protect END_PROTECTED
