`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7oenuaW0CshLRyOtIjIOFLLqOCB2sfPe8XNkGFHXpsrvtaSskdhs3qvzuFJOu7XT
LnVDyIxjVY55KibhxhLHVpARsuKcVEDCcRRde2PO50RM8w+PVNZyj0Ow4Y6edsqz
aU9N5MwutPkTOFDSdl1ul3bcHdVPKHGmQ9NqbvRvmt1p1X3lCn+uxtz8eClKLxCF
GemUYn5Zma9RtjV4GSPuGwztJC6r4OJ8L8JxcXDfVRzQ+4PltMGzH0Z5SteHhf8T
6IXI0UNok6oFoySUMmAH0NIR0THYwIZDdk2V5thWbpqD3uhBYQXkzt+JqRtoxjXV
Lpq+UV5TvcpagOKMyzr13VHIU36+6YabV+KjtbA6mAI0/UCqCICZMQc1QuZj5bdB
FpxzdctwwD1ySzwgZV+R2P4wDe2pqHXmWTArlrJC7lzmNZPtZHhaig3wbY3LXeiG
`protect END_PROTECTED
