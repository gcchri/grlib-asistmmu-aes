`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fpLTCdtvLkfp7EEhFVMW+Oo7iISU8orSY45abvGH8cF+BRVna+S7D/iUwa8Bhuur
bvM2Fw9HlZ8jgBeIPu0Oklnt7+jK0rwmTq3AMwvg12MX+UZ64JacHQVNpvjD8mQD
PfqW2j9VKheuEXHvNKtBvsQvuBZs3+fyGOTF5I1sjtXHt15tySlUriFJ5mdusvWB
75JydI3+1Zn0O7bniOUzNhMfeyzWNbgPuxppr+sNsunQONNXSMPc34U6b5MWzTqk
JNKSODPGYqlv7zXmjhux/sGtgXaCFhF6An2XZt1nPdLACmrhGKfs/qnUaBSD1/4y
5L8ME4e8OVnLdbgysJrMSpShARfhwleOVePJTpybb1PKGZD0SBOFWmgY2UdH9kXw
YtccKBBvXx0tNya2Xat1QCUyGiEK0aHo9L416uFca+3nM02jsSiWTUrIf9QaypY1
rRs7f7qDinzOsRcA0o11KKgycqf5D5VBui7jchdx7nSzpb0jewq4rnxVCHCJHvn/
v2Er8eFJDHypagwi2FRmzRj67ZFeag1SKKIvrNj9gBsOoX3GzVZkWhwrte0Jrrwb
DMVNPqHZFAiHq+KqHPtLu76rS80wCH03cG1tMRl63cJfliOFP2LL+cY/5iJ4kM52
`protect END_PROTECTED
