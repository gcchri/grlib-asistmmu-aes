`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyfwyriXSWhhTorhyoA7WJf2KXmuz0K/Lv4HoCg5Ii32z6lIWK4c5qtJ/wEmoa26
Y6t6kbBmNxmF46O6d6faL2rbiIg3iBxTHDp8TtNGVrsojieJo//r5E+OBpwUSX/u
k9dkPylkOhhjfAF1PIjHyheC/GQnHvAWm7Tas4WVD6aTpsEoEF82GxNu/D7o9GRn
Pa1rrFPIzRo34/YrLAyCOWkCgjhgm4z6Oq5bYPLPAsAxg5KTpCoN/qsEOFTlv6el
lzI+zMQr8G+p9hxrsKFxOUGX22BfCHDb/c5tV6lsfem9MHBQ65aWu+kGVkZvyQ0d
a4KFgKkF+We8wKHiREUc28Ae3cc7JQdHqz0raixyJRyBCH5LXd0XBlDi8QJZO1tP
JjToKLC2niDv1QWhEe+5TdANRCIkyANJ9aKpS7CGjxdjYW4ZxBcdM2DhtNTwkT3J
XAUTRv9dkP3Hw+MG9dEtU0mkSDqOagOS7N6yFQu3ONY3Ls+Kik/14PU3V4NICC/g
Yi6NFZWCylsISl89RqYAcGUyUyh8y+uI8bUue9m2+uTW9FJsK9VoEI/T4IVA6kL/
PszBBZCO2+oY2VB+0QjtfhwSE2pdLCncer2zHTBcqxrJzPd1mQZoB1BjKtRClFQ/
wiztBhxzkhu3liddkNiUD0I94qQ/ItbFtaeFJAp2peblLx3nRwbr/xh/8haA2Be6
6lSjQa9861hOTPy+6AdwcX26BQcrad6eYO+H+5l1Sx3ogXh/FjNOE23SXrsXFZtU
MJyelAzEZvGq0nJ9+hJaKr+fZldNkBTrSZA3fHRPOmk=
`protect END_PROTECTED
