`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vouQuwK55RMBMPdl8RRG/ppI21He6OGBv26hT4G5sWjunrboraqT7nSGyggcbtTw
d8wEy7q0CpGHw9nS6za0Kcs4RwDIP2WaY40OHLbszPEDo0luWK+iGZdD8Yi+wfe9
UkBsHkdyUHuR1jl0dg11yIczCMPfFU7pZAZ2LAYe+z9TR1XMdDlvBksbs2AG5gY9
VuIM8gNpLZbAx4mekFtXgaWUfdWhcFh4ADZibnpBaRDo7y1+7TCvpvKczou6AMpt
kfKty94BrdqPmRjcvjP61I2f6bnVnagl23+onGkGPr6+EYU00hTCefqWA2Do/oaG
Sv/nCmDFSaCjIQKqeQisxzgzEgeYCzXCdWscViYQGTIBTXkq0Gi+vSz7RAc69VeW
JLEriHWsGtI5K33grqx4Ka8dzhE/QIw8sDgjUMQx6n2rIqkDpGl+8wMdlHbFobGL
l9W0ZYYr+WqlrVlKQL1oXow2r4HRb5PPO45W+HJTfio2GLPVYzDjpEeDvWeFw963
OGG4S4wZ/xCOpJmGju6ClnLuNq1iltU/UtO+CN+VQ2aoCIPNJHn+qPKs8Dye8mpa
Nuge7vFfFETE9RHgQ7mQI+lxoGHWOt/TKSud7PvlqqwAjrw4sOcsuKKS/zkhiHmC
l4k3x4ObpcnnpHZz5KzFFFkuhLOj2rGe6CX2LLTZDso2VvhGNIgYXB0h/KoJk5tc
tpUba4O1kcgGqUF3g9LhLhRgEtvzSGqt/O+GtcCUNta2BWczzH4VK9CYwdNMxh34
/IBOgQinLwknsHg9r7xwzcPh0ak8qfMW8vm6NFx025PZoDgC2JAYngIJZKr1kGE+
c6M6zienGfA5Gu/y7dYKj8XziDetC5YG9gCYIVH/e0klgqbRxx3Su/jjClu+MxKm
NDe3+6RmZekDhzsScb7HtrZ6ux4yFNPhC7QHqT1X4CrF5GUMCdhwHZ2Lw33sliBu
8xDpPAphdQ3IRUVV5/6GLa3YBCLZM5UswuwSQReR0MA=
`protect END_PROTECTED
