`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2idAB2RPAkotUjGP3E+/tkEyCxfLeQ2xv1IcLxDzVmSLQ/dvV3q9IXQXurEAuoyH
hYz8xzMZ9ZhPp93RSLneYSLakDchmGe811EJ8HRIEVa+Zugav17gAAWVquJN7wKQ
xzvqunTCvpVX9Q8k/tfu6DUnsK+Ygc9kjXaZ9RTh4o31mM9hjtx5dC7yyVjdObnU
mmKzczmqjhJIC6yN40VnEnwYjZj6qP82vQ+LWlyo+BGcTB0F3a4xCMHLWTDdXgBq
tGXvkk7Wd9QF16BbdrJ3Xw==
`protect END_PROTECTED
