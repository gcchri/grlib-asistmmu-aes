`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eO9i2mrFO+xVc8TtlOxlQqRZITa0u9YXIZIennbitoqNUogfiSuAjvREDBGusKHj
jE3CwWHwlKEzRcSbjlVS+kJnDeUYpspTxWHcWt9F39BFJuINZye0qfwBJV28SLTd
dzCAzJvvBzc+wTWsDhJaoWVz36OGkOwCO6B77uBx5EzmtyMY/iJlP7cS4kH2n0jb
E9etsKkMRcLl7kCbcNkHCUvPpdkjKcSSBB1RFFXtHVK/O262TcZZb/Ebm+A6XnpQ
icECBGpbDlwXd+C/CvA0AqC3iHkYvxQ2oEtzjrUmqAzyeEXuv6jC3WHn2el2nWJb
7Om9/wiVJgZridRlRbSPMg==
`protect END_PROTECTED
