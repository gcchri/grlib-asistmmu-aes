`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pICheWg05xUwE3rotjPGj1b4tv7O6HfqJaUR+6/jNuuW1IZtSRxN0SyV8cWxa41r
Hm68NqJGZ/UHUd7kAOxGf5AOTfvEhMz3Hi5CDIVEJPQWc/rHiEkWu8EEZHIHLAhL
PO6LKVspywEDbECiP4TPfF37NQelz2fElxlgcNVEc9ML47XO6OGD2INF145FZ6qU
2izrqOIGwZr+u2SCH8crsy9IzgP31tM7P4MBtaQEEGw/tKUUtd/IKvhW8dip8CCl
JR3CM/ZRIGbuyu3hq0IvTJFcAJFRq41PtlYYlRCSDCTamIqnvbnW+fHLU/zRGSkl
feLoVOGPVA/r4vbcvMhLthkjE9D8z9kSCdRZMcfSqu6eeZGd5PTu0pTDscNm3P5L
GlDX1eVkEVywNnxvoFAiMPi1UAGgGgcinmuPk9eM11pA8YJMTq37g99CgEsHVGF2
lKVmqXA1Z4CHzKDtzq101LEfB6Qv6Zxlke9//Gbf/Kp8HAMkSGeq9jkKkWY/McbB
J9q0AIJvZozPdpzE7QdWeDnu3V58eFL6vn/tNeZwSXCiN/ZOudYB+T2kzMzZq8qG
6CvEDnoLIt0z26t+iO+9UcNCJYAkpNYv5ELbwvmscA2uH5Ep9v+6vQekLG5hoqes
Ir/tZHwQLSQZjxCdIBjP8FwXfLb06+7usW8fNuhjrkPJPDkJhacvaTJNLAdjsGmF
AfEMj24Tc/AXzSfC7KR617TcTe61US20VezdJ6+qzdm8RQlstZD2Q49SgTay42ic
0UHa/aC9btuGykKAsWkGq0J/d6mkKISJROagL4dC46ns8ZN/JmWFyqHak/dFU6M9
o1MOrbs3pF/WFSRi8kYOUttVKvq4fO0Z9GY2CTFxU+VRG59fStIBxFcRZ/SvEj3N
S1o9AFR+x2Csn62QjLk2qUgo+QGM6CYCCtbN3XEARA6ZqDXG2mG2he82iY2CZba6
B4nhGiUyqhOCzNi9K0504mkmCGJrB7WpBlYkLuUqtwU=
`protect END_PROTECTED
