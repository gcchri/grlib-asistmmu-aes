`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWAt/o5FkyKSazkX6lL7lDi3W//BXiSFmyqUZg0oKHS8soLZkdo71qR3ivueBdIS
eQNRLksZJ9vrVps7l7sLI8hSwluXGZuDeWpD834pmFVVQljlnJtcock3B972Y16F
xT5JWOR2Dei+2nFsejHol4tzNXhh2iPuN2aKK9Gnrd+hdiZaKA1SHaTy3V3raN8A
/iWep7s05ymJUEW6U4xFMTCIN5ACmZ15X5dtc2PQU91M238KJTm5cPLssY2rZ5C9
UNYtgb6hXy7BespO70ez1tI7HUY1ecC9eX6CYIyr5FNB3WjyaY59JlAWLrfjLff5
yp2znDhWijWN6rbIJaXBbxiqHJ+ACAm/FsKaxGS5czQ=
`protect END_PROTECTED
