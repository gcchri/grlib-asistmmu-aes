`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RuA6NhNDgyFesD9GCDbiGzkfW5Il6i0laBwmQYJTzIMdcDLPLNmCb//jEfWuoLQm
k8E+FR42FAYYY7zUwWODWTghdZTrUnp5MCXPP0Pkju3UQ5WVM5gBdMgqLBFEmM64
chwBp2o/m7vT1u8AVaHd9qjr8ZUrxHuSIcdwadAD2xPm+LyArSVpEI8ggVuH4t/N
GJW35WAbz9FJv2ZG9ioH/SK+iE/z6AHwjriLbzgf4M6tO9+Nu7rC2nlS/NDC7p1O
`protect END_PROTECTED
