`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ujPNz7s+4VJ8S023MW8wDw+v2IbGmGX0eDvzQfBgaZXKnlp0d6suZLTCZPniaEYf
HHk8GmmJBIpAx2r1TqwCxBZ+FnvGkRR4Bs+zMPB/cKHQ7Q2TZcjFqMVPLqUVUhq+
8/KbM+Qo33v9g2TFVQZlW91qCvSSfh+kBuHZd9nKJQjVgC93QKbI68wwcSVBwwBt
E/ys6pA05v+YkhQ6EVTgX83Pv3ppQwdZQRRa06eppMmxoBqdvVlSTGRJ/oWbaKQ0
b5Jd8aXT6Q5vjRuS7tTPKz5TIMTx8TaLoN/3aJBQ6oNf8/1gdzLwBLeHn11Jrao8
sET4wSwDZRBT/CWckYO7jVOL4tQmh554Lkbpe7qahHC1RTuMGbiuzSYNl0A91FSX
zu9QqgtjyyU84JLEYk5MHfF7sYYeNubeuCI3Q2Sb4Ce8Vckd6hNCgwiOP/MWdGPR
0+CcBXKjQcHj+7k/mvzaxGRHJaUJAbkZIpYP3u2UKEgQjpEI0DTB4OSci1+ccwLS
hDGwmQgwJsileWsjErC3yA==
`protect END_PROTECTED
