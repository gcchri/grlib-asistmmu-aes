`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rUTQuyiI7JXm11wVpx780ZhsQ5NU2GIzUfj2opeg4sQoiZ9fYAnxsaI/znUkT+MR
1N5a9fwggOP63bLsDZe75WafC+BSjuZD0FPh2HsbofxYL7ccz4PDAzZlwULj8870
lLVWpcBcmRwoAnFPcxv0Zy5u7vRCZjcU5Be2uec2EEWBGuBnWCjJL6Yz92mJmBAc
mmoveJ/tIlfi639/CVbA7cRRTVJFckr2WeYxk8aujSeTPyzlV608lewl77N1fGA1
StoIl4CBUxk1jsl8FIrFDA==
`protect END_PROTECTED
