`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ypwgroj91zf7qTY51GNYJk5Kzv1jc8+kmvxWfXiG4rkBRbcKFElo6zJI1y58uHVJ
BUgimVH+eMJhr65/cBxs1c/sbAVzXnIGOAUG0GXXM8FORAjhF1Cqz4FNhPqSCkjz
nK8O1VQJDb+pQ1HitmD89TP0knhOXVWbtETiH2yz4ZS7tZRFA5OP40QZLuy1xleN
PhAxIWZYw8flNsrhyWzGQZQ+/q0wx2G9DsPqGhEP3EmsrK4lAstvDQZMzSjwYq0p
o4o0wQp6gkYpPlOAlYbciK8RYg8GY5pkCsPToT0JzaE=
`protect END_PROTECTED
