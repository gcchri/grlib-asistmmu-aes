`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/Dut9a3AeLz32cDVtF6T1wU9Kp+JPrbElwRr8P6lErIBos+dNIOWW/nP8BJuezX
sWhTI3d/5ZWmV+TEXQ7E+eLyC44Tpts6bggSGemLOPV/+BMS3lSzSsi8mXK5hd7C
bLo6XF1Ilb4dUF2c4CY8VtB5D96Hm4B15XXYUP2CTjbAuNcND+rtRAqxiKFOW0Lc
IXp6VNQ5RxAWDdrjP9RxeZ9SYcTpKlYqbDrc98P6XNukqikZeg+QYvu1Y95kwAsG
eGm6pI4Znb+9j27a7SdEYICaMgJnTeWYlGb2wdsazu6NgJ18wy4ggdrppMuFgfAv
B1vdf5EieKbySMf/eNwZpvA735RlgqU+ld7VmHWG0t6XvAbXPSR/8QoFqPDtnWWo
ZHvGAC7gL/TfM7GAhYFfRN5a2fUbeK0BwWXNgr4LECsX80wUqkTgcXfqJB60dim9
`protect END_PROTECTED
