`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b47quX5ZmF+158qZ+biQrEzXyQY942VSFO+0o7ON0i/24iiyZFt6G1iweAKb9UQR
VoMMjcFQ8dWk+NSeLgtaVXfOjqQllRBPugrkPyfARQe3qvJFDyBGySX3cb6nz81F
dKrIHU72Uh0JiqsPYXQj+2saHzBr0yr4ApTXpnz2oB8CxlTfAvHNPQkAHs5IOVr2
G9blqeGWEszmLKp7g92XwiRapc34AOJBSJmijjxyYm5kK854ZN7Jx7ZFj7AQafl+
pDfkFGAeWukcz86SxAkphtbnHMHQXkyL4QRnIxR7+vVvlSkPSC+xDQZy8DYCNoWW
E012K3Y4LNU6QtxDIjSdc9yZ38FxWtN6EHYtytnhmiRL/HUdOA02OgtOmAL7R2Xt
R+YdJSmU2YrBb5372RwRlL6Cyf5DtAH+mfALpVvrtuQ3cty9GfCL7svT05SCTAMD
sgvOtHnW3+p1dLYWOQNkpA==
`protect END_PROTECTED
