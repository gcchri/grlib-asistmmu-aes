`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OnnKY1TM36o7jIFtLRlVBDzllUr8LkdpMqubOJO211mdMmLmI0HZ3mEvwGLQ9HKq
Zl9dJwbwbm28oKdPKZeIgFNGTnp44yZvBsl2unr4LWM2Lk5kebC75yA6MBjtZ5Xu
mQxZsqGMZ/uUVC3SvxOVY/k2Kb1g/Pr+AsygwI7W/beeXjMV+z3/ldHbXLmdKXXG
+1YwDrkaJcT+hoL74n/gzCXuXGo3dtftLpvQwB7nGt3BrbO0ddgVGeaR6eCB6LdI
2Sy7Zwf4tWOR1irRbuFB5CZcGDT5bMnbVzWo5Z+K+BO0W8EIfCzrxDqHE+h+E4OM
9gDeidS2C32YS4X1tajyWNzclfQWOphqoojJSglGdYU8gnjF66UQKVVoJn+vFCCw
6+LV2rOgqKGGfHJIeQgIfeO+rtL31XL23IhCUJCFyX0KuTISZ0djIdpa2kOOZSvh
8TqxxPbrss0h71eHGIQKpXXj/hBzEpvTo9sb6lNYFCnddlePf62pyOmKK3KQgW7Z
Yd9bV0nFvkHir0zrSRbyOVsM/uQCo3eSSyfn0/fzAN+eN+YBHZl9seR/fd4MF85L
`protect END_PROTECTED
