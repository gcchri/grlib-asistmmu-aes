`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cRugKUkby4AvMonVV6ncGdVIqh6/pd1hCU8BT0Tr0wqWnO1JJ8vLNxI9aVBZqRMY
Q3+1K86RJypfIGhLgkRFr8l2xWge0Y0+HJEKC+bpBUZehfMf1C0iEOEAcD3OstOP
bor2Xcrji8R1Awi6dcz1Qg1sh1GoaPyc9IPAfYAAUkPQPL6kSp7xZTT6rF+eMnPM
cOG4Vx/h65MmH4I5BVvlDHHaSoLMbxgsld0nC8CGN4JREAfxqYQ3oaIOSWNuGVWh
K4Fh2G2PO9mMjSX5sHXv0PCoW/qJg0f3+8TjLDgwjJgN6ikJxJ1bTiAKw2+g6Xhr
bu8begju/5m+qBq5MvqR9W1QyZ1lHYjO4UZldHnhskFuV9kFn+70J5V0sDr4RiyB
YiHXQZfcvw/I1kguqX+C4TOa7KTgV6Blj8xm2eaTdAW+9g/iJs9fKywrZXFxlAIm
B2M3SlBWex2UPPmUvba5LzXU95987rm269qU2isGzonU9uq7LpdmDDFiEiVirUMw
6MLun7KNakURN36Uae1K+TjEHBAPjitD9ESu4qiA16HI+ZQBKcAh1NQWbE50R/nD
`protect END_PROTECTED
