`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sss/Pm4oaKnpYn+8klXdNKcAy1QOas2arvNpdiHxFfx9uxj/B5s1CAPDU0/7wGOB
5EER2tdaCkqfSByIV99AzlNUD7nWmoM15apLOqZLP23e47XyjqoQVuPEkAbwHaDU
ztMh9h6lLJsuctUAT3jTdOE2p5y7uvzx3472L2kVljvFTRiScgyUaLKFc9ij14ue
uePIu7l0rthQ/fry6eWgZ1/nGevp54JJhzr4UGxmA/mrqS7G82/2G6HOykza82Oa
nhU/OArOX+S5impfnwQWz4+8yLk2pSaB7weMw9hNQyO6c6JLnmTdspgnuFnde/TA
T/FstulcZgje/6vErUjGhVi8Hlu6X54yh46FWsCHsJLnECwnzahMsNftRDirr1jl
8cRAsQSE4zFOu8XmCtzVfeluDEusLWEzHo88miNxaoM=
`protect END_PROTECTED
