`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
auStmDSa7TOuI+8OMN/p0DXphkzv3o7v8gDBbj/tO0AudXuEBclweZhXu+Av1lIc
u8sYJBpjGY3ithMF8984HMmRaD44SkNbDYL0581QWxme+Qdy6lLXRnwXtsRgKkQa
c3PMyk5jcerYLUH/Cc+DkwQ5Xu2jiI+p9Gsw7H93OV/3ha9VOoyZ5HQbgaWdQTLC
wXHaKksIV5hKvEtwCCI8yZoOIi8D970MZh7S2tITKXk8mRkCKfQhMg5LqGlCLxEi
rUu6tpUYgbGfRrh8f+KmAa9p17gwKhBG3ShjtPWbDKZrQqKeXF0QCPjy/a4BSV4I
rUVviSFmaIv0eMrFFQZ599DU5SQIINjSOu3bhoh+8PJR6Lk3R/cvLj6Af30/kALR
/NqRkN1cEps+RfBf3JpjzMLHPcEZk1jvn/efWy1Bp6s/9naMfvWhUK17NTUY7B7x
/u4xh1un5jNlepDCxdNGq0A0vZFdJ2ggTgqvkjdYCsJQG4buYRYv0TfoLOo+0SwK
9idsYUl/WDk6b+s31f2pLG4hw7t+5dhNRgw1AGDyb3ljVc+FbP/oSliNDmcoicjB
5TGIKSfKZbcN+P0eOrACy4+9h916SiZIf+TdSpCsX7mkoEkNAsNZvk20NhgkH875
NEqQGcmKhZSIaDfgbOtBtj5b/NQCC/gGKZR39AlK6Vvoa7topXgv74v+Q6Bdsivz
8yxzXJyrAmLWEMv4q23IRz/yAU976j0Qsc3VNbhfqeyAIpuDydNCHeonS8e5mQTt
DIgJeUKgSSFUch6MRv5Z2iE3qds/7w2KmL+snoNdipqrGiQAqEr2FavMwk9gG/lY
ge/jL12dQCXPQ8E68EvOGny6XVEa9hb7nxUYcJTsS9I5pSt9E8IMiHV8X5de3daT
z8qvS/Z3NgUqCV5a4Tprclp6kyDyZYQbuopXa442fQhBE8QeVOFfw/f6NZ0b/oWr
dGuuMeBCMsEGchYP2Z2eFN5W0SLT+MV6vPl/oHBla1+WU9mx5ZskB95ZLXvvtUSo
NDaUqijvj43kqAw0p1mtTiJ6c4XHLBad5sajzbeGBb3mirdUAnkeBNkR29K/TIYl
29AH6O18mS4HxFHe2cx1F23vrX8gc0ZGqXiVpZagNjdv6oPLDjwpZ3vwjHptjEqa
ppQqSm7aoae3DMr11ymYS96oU82igINeevrna0VkC8bTjuK75tPy2pkD6HgrOFTq
T1LGnpI7aJFCm4EqYGRQKoOeIkeSG9wh0GgIzG/R3EF+lC3LneFlwnVXhiKmN/VZ
CGcpoXSGrx09GsZNVf/DIRDIUa/w64MN4zuUPps0Ck9+UfXyiddd0oImds0AXLsC
9aeUrTz4lGi9PxbdBt5d7WHSdb7Di5j6zCiS/NqzB+UujLmk5TMz+C+z2C54NTPl
sQGmcagKygiHvaqvbMJSezHF3RgHl1cJdSO3DdzFOv/UulMxNYAx0fEqgwR8uRtQ
D9Gufl9WoDSwlSUPgHhubpPa3LjEfXHNYI1IEN3wxFYxqIVh+LPbs4TNa5Z15Bce
swNjVuFBwY++Q/ToxNIOwYGHt/G8CZGpphNqPjLEqEmDzrdPZSqcXp1xOJb1zSwB
7g1ide6diry/SxxZyWtSZd7kGL82gc2fpcu2AlP+JEqBYPu3ESv3UuwqPCczoWxS
6ZcEH2AradS7nfdPPM+FPeWxM0bV0SEW01NBKuSVB8PVO9TONB+pt2evnm84uqqO
opayJmM7bhZD5epS5PFxdGEG/TA/TL/r4mR0xt/54SeKk09XydcisJsOS4xxLrgR
optmrA74GkMhbfENCJiB9AtnX3z/yXSKR17GcCbqLkLe0rZYoFl2lby+pD+wSx2+
DmibKB2eWYOVG1/s92vVc5aDJtS8Lkv3yZb4oaMqMlL6F/ilCEurSm04C49Nc3SA
w3gLV2NdlnpRZmEuXfxwj0OrCpHpOq6YUbtBrjiaY1+5hYZS9ES/j8BJ94VBTdjk
5gl6pRPxoSQTu6TVE24kly9fWfa02AjuOHNJDvAooRYd3nKWBXH/U2I0KkggY6/p
fU/n/jdwM5enuM1Tbw/fRA6H/SbYQBEcgJfdZ8bJgaecKaeLN6/TnMDZ9QTaFKee
iAl2SGqZudt5X8Q4iNNGeonCwAL4F6F6n7jnQsZgG+rBMXZkHC2RmLC9mEhWAg/2
hIqZqMrttw+vlsdJVgvsebhHud3GtgbFckrnD9SwwYKZAo7izyhre5C3e6KhWtq6
5JP4BwEIoa7K99dYv6DVxMvMzx3TXb300alwqdnFiIA5xrDUh6lMeF55DfSoRpV0
GhzAQnbfMpsb0+IR+eWUnVlzZ6iIAnCT7lV6eMdS0xO6tVouWTrXiGyzjoonqya1
5JjctU/uEJY9yOLUwRYwU4j8OFvZfpqNUB8TgnReOpRFxYKtQpmvZi2V8kc4Jg9x
MXyVjFZUrlfHTiKsNOBjiUC6b/mlJTIxgVKOTW2hqsEP31iuyV8iwHxlrtfg5fcq
+TTDr0z0YFsNqb+QWBZnHJ2+r20/D7HKWf+ef2YhpHoFq92lBfm7iYJ5GExgjNGZ
bpYKa5cctXk5kwAtOEJQv/5p5jhKx7nNW1FVaGbOwCsfr3isPOFvEghOrsT14uPD
/bYwutcHSRpVQHQsPMUG+4B8/v1MUI8sg9iV6Kq/dAqsZRg00uF5+fT2Nsobq/43
8wq5MW67o9dzw43RrcfXFtuxlREmh7q9Z/nVOhnW1T1U/oztMHI1hI+tqQKU99XI
pPES6gaaiJ4YxEmUytoQB0wbENm2z0FL/7MR74AI9qdvSqKqeUZ558oSEMAZ4NAy
8QPCLK4mZXJOKkydWon6bV9gRY7WeIuvtJ5Am8pCap4I/9qjF0v9M0YEKgymMD5/
sy6R+FxO7qob0cFkFgjIHy6EFVrwT7OOF1wf2EW+qbiDtdbXr5xqfRbmeTVZLVmQ
vwpTHMxn0GpGw1eajN4Jw2cGZxd5Cb4Ydhi9k/Xb10JDVVSyvl+pN5Lnr3l04iO0
`protect END_PROTECTED
