`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pB6edgGUVWof7w0vvYc/QE9lCzmaILA7ojW2d4hbaV5HtXOTUemzRMCqpQ1TRJW
mp+xOLeUKtQV37x2xd7vPH4VezaGnUdNd1xahQDp6RkNVKPMmREoEcwKLXGqxNvO
e/6igVUAccKdloSEFL4ZxP5IQq5FT0cUHJhMDu5AsIA71a9bVinnkxtgVIFXmQ3/
ezlJMJgibtZdRXye7LGGXmRVnjkwRrPxwHmG4LcwBuDhbv+DkVWLFQ+80HfCb09H
H4J0BdPdaBy0wj2tT1X6ryMfwLUxJ7O3kvcQNU2RC53cyEeO/VMJ3EN6xU1rZ1V3
rghQkNXHSDvoD5RvMIteLUppfv/YFybO3qUjoQBvO9oBNGkROQYduyxtTRtfte4U
VPY0TWW2x70pI6EmAbevInEBTPREZPxy18awwAsUQTmJ34u3PwaqoLmLWDVP7qny
jg9VuERe6qPMKfzcfnuPHbE1EoNoPYgMxvqo2osLGgJcyZPjySCaigxELsLtE66T
lHLGmv73xCMuB9/oy0EDGSBbH/A0OM5YyBxHwp86aWg=
`protect END_PROTECTED
