`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NQahK7dxmmifQlJrpzyIy89XFFlorsW2YhpetL5Mm5CzOdxIXhWAu2BMNEwZbvv
5PjDjz3vQ1exYTk4bhDxXCi1vugoNjAFgYUnp929+J3HK2NDC8CUkVNAPWUq4SYy
1siZyRipUEGEcXtHCa8wiGLnr8BRkU5qGCyi21S6dAPji/NT2Zb36jj3w0hXtGcV
b+XvzLakfPJ6mcWR7e+ck5jRwCxKjFApp0aqUsHzgyG3YYl+46erqL0AfAlhmIJF
Mixj6KqPXHRIBDSR3EXHIvE182rhxtgOzDSPldvQRMlv2fY8P5rMRrBxnjkAgIiB
FVaFjpSr5PLfA4a6eX0rdCydoVhGuHlUnkCAWEMO1C9XY1D30Evx3BOSTmeJ1xGW
A7JRhvsO3JjcnG2yHGvdmO8nNAsC+Nup9KPexdQzWsMDiCJJSRrcTWeZDoWlRroJ
kA9LbIn/uVUmGzaLUiUlN4gXlg1AnUfeKo6IFX87CyuMT0L+EAtmaURTH2w32j+O
g94EzOeBlAthF5AwI0WweBqz3xzjk5MFuulZ5o3N+V1187SZu9ZVN/cK8qZHxKiv
Ymc2eH+tGvN20uGp+3TuWA==
`protect END_PROTECTED
