`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
on213nvzb7Kqt1QPWSet5GnZxGAooSvBlo4C0MxGfDbzrUAsK0pKOhi8x5plPT4D
MpICJ1/FwUQ+ndOpf2dIEjIJbj4+llpuK2+RtSquNlT7IpV5eRPQgotSeDBtmhh6
iFd3NKN4T1P1mcwnN3bHs2Nni4qaIw22CE3k6+PVdZCWwJLMXp2rUXA2misYAVME
lEqk8CfsXHUXSlpyRW6em7Khl7cV8WOTCSCZqn5e7kD8X+TGWGr2JZsE4t1RR1qC
QGPKubCnZ8XBa3fdpGiQvi45YEpyi6UVUgjbO5wjbCnRTyULGWdrb31a4GA/rHGI
wDPmS/r46o/euMvxqUItCUAug1Fz4U8AouSzS5i5Uk0/3y6eiW133FgdA1SymZ6B
GpR13f0crmYQELzVkb74R/a5hQuvDcUC07GXVseCYbq5EVT2G5HxmeTvcJsPUbwM
XCy4fVCCiCTC+w1RQ5qj2eXQ4iewJAlrT/sEWdT3FAE7febV4+xNbuQpdDNwWgnE
11wE+CxCJJQGTCe4XHjlQH9rAURnNlSOmTvFWe6kqDM6KSvj4VthFfRlGe40QyVU
3oWTaebOx5/V0uaTzLn64U0iDN+UXtVXkX7FDp+VjeicwSAeRxtkRgt1TUq2sqZY
mHEBvJqc4dFa8wvjzcJEUqReUMpgHq8QJGOKpd4xYsAAv/DIhbqOL6hyb0o3EGgv
uu8FjADA6FNyFMiUpyzF7jcbnUl26Knae3fiQR1qwcCGbsuOZ/QvXFE4fhK59h8e
rXIFW6nMH8JXsqK14Y8xVQ==
`protect END_PROTECTED
