`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8LhVCGUp1tGkq/6zgMfRWkDzxRZ0Jh+yWA4/uBObooydIBCDwtxrewrmhvUvKi3g
ZlueOYrPmr4dPavO8YkWQo+/+lrlqwxNA5MuAfZyWFGrQamqAWrVYAf6lCLiHSaG
RfniS7nm23wkjfu+SAxcQqhod3eJinWFd+ihJ85+YTgWBBcBCVVHNSc+lNaI6m71
pnQ+FmiT8X1HwiRIOarM4iGmcInC8eZGWGBG19zCFPTEmV6746ZK2XnS33CURSp5
Exre33tMIRoFTxojyWT/t0crBtLN3TKT9gx71Yut1XPjyI3Cyczkkrfb2VJ2keea
2ZZdjjuLfUFQnZ+APB65KtYVegYPUUYStrnRs4OVHj6+29lYIWF1mo2xZOkwp5zz
Odv60jH2xsiCejSgeQNPGcPjxYJDY4TGlhOWy5DRgmkaroKVIEl7zvGNQ8iY4iR9
lZ6inYUDeQzChwNSJKlCF6MwHGaBmDMPW1gfd3LtjrOyIyIRcklWnmzMa1AZdxih
LTbkWzPxabxNupQaD6+cjnWbadDvfnvEP8Fu3J7AYZC2T130b7Hc+o3LlV/LgdWV
rUfPOJNHMyJvSX8MBifantoRsUrH6xd5vvZqrFIeVCC0WS2ypUjLDizGSc3o5CLV
NxCQRhhDfW31yEnESBpe2k6Jp8l4gwRWx0ISDrClUlmBfC0WMj3079e5Vq3LUR4W
mcMzML2B0j5+4b/D5E6c11TWqkWQ417coHBdYEb2JaKF0Z3fl5axO1TbB855iz0T
bcRM6+c7k+3gDco/xN9ifuAfxMOJONIw2e7e3EnRf3Y=
`protect END_PROTECTED
