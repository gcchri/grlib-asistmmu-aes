`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ym/g96jEdKZbM/HZeX2JOvUiTd432TRbh4Ozz/yqZFmRJovn2wrdDUUqmos8RhVE
+/FphDVmeC2iZP6ItboH7QO95mVeunlveC+8kQBYN4p14QdipnOkDnL18DKOkgOd
D/l4OdBeKtSLJ9ue34OeEB6BS+PnDj7LuLp3U5FI43Eh0wkTvVvO7cW/GVAb0YhU
qOsdrfwhzRC9MUI/bQDrFqKgvIoTDce7HrfS3zWpWrl0nDI7a+sgUqMm732w3Eqv
E2Y/WqkU5ScwD3ZpssT+Gu7YfTGlIiTQZuEQUkbzGi/nQmGOaNTnRF+vZQbdV4Om
50v7zjU/TCH52GDZFqqRuxpd1j7Kj8rx2Gp7jeG6XojjfDd0/+0dwKFtOIZomcQe
TKyPx+5VceaCf7xDhKfTN9sCl5qljP+Haw+MbbMJgFiW+pGIPg0I/SeaIzGT+1ex
zMZM2Hjy24qnBDA9DVhwCvTr81HEUeY9DpC7Sbt6i6Mps1OUNGUOxJ8FX+Nun8Pv
Vxo42IxaM/PvPYRC81LP3fA1MbV2/FyiXVwrFKHe9ZZ/WQCHnNkQddSewSnqFCKW
yk1b9pKvbLEa3FQrIa0yW9Hz51hTlqYzmyfqlNlsOCc=
`protect END_PROTECTED
