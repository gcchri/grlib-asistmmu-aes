`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P5at43sIi4y2Y/8vHeUpMZ/kBzs1dRLnpfw8UhBXe4TuUtE9HM1nc4INCOopljaQ
n6sXd+cqEY2t77xnF7zSwCqvXx+nFjKqAUk+jxR8WXIJoD+bE07+S5R18STxpXmP
wLJZpcUwdoefXxHKWQDqT9fcL/PjIs9gbgx/apS/x+iJ/k6i4XVV0hFEG15u/m7J
B9A48KMblHnkgW8Z0Oej7hWSxRYJNl+ocC/FEBIgeaI+dOEQ83r2nYCxxZcE9M7G
fYZzPNI1EWEqaPs4bGsOz4lqua0B3IYletMuGaBsyw4IlcnjnIE8fy8rFqXbjMFW
gFUc3szbNdNjHxg9ZoePHefLABzCkd7VhOSFu+MLDmWRco9NAbfZ1fCmpG/l0LfQ
0togKsHVRQvueodh365TytPNAaihCtoF5m9ahMAsC9Ok0l/HBMC1cCmd/Ib5qiZT
Kgqw6tKqO56YtFgUZOos6KWB1fynRh7pY0NH6udZ8Op2OuO4IGLgYcLJDc/YDIH8
vPeWeu7+05PiPejAxd1DOCFSikSBycgZqeKmEIsjlPifIkmsiMxK5VaN5gg/lWEa
0UyeMk5nEEehDo99brrtNuA6hmVUFR5p1VeURbhyX7hVFKS7nRZ237ZRL+K8TgTX
6k7pNURXTlDbN4JdE5aJtH+bv8AVSBwk2wStJZFSGvhWacf26nscSnFxp1DD8jx7
wwO2/5hM2hI4/POriUCyvMpotawupS8X+beO18EAL4meXj7Ym1hVgkX7nqqHJLyK
E3JVGPBKTIanPlYSy0yA0eIL+olqLxc2+4VZzy1fdyNgE3q6kUZq9TGOyquaz64y
vqevTAbjcrTpK43uGBnwLDJYMWKvPMGGg4b2HSGcu5uZuDhDK2zE+fjnE5z7FP/b
rS+itepa5Ds73k6d6h6ELHneOCJdsFrGj5tFb9o2rHNEmMOTq3gUFjZ19WuYid1Z
ZWgtiopPHGeY/uE0p5aJ4x4Bc8m7Yw8Ka17nLgIsnff6uEz/ftPhLVO0flS4zxm8
9DAHccBhm19BixR1XWIzCAELL9OyQ5CVLcI7UMmAkiZXNeCIzk2edvVwmBzVGt9a
29W5IgVQHl7zvIV/TcM24Da7MJWAAjvRIpWYzPV4UJOrPPVysOpyeAb2/AHM+8qU
0d+FYcoJT5jv9YCjCRbDVF8Ahy8ok194uJ6K5mP7NZ6Xd2aSyHZQw37hNmS22Z49
mMkEfTRnTr2AdemDiF5dY+eH1KTCyVl85w1t17HaSB1zNL7ljqrlFMW9mg8MC29A
FRKELc8vKI+QU2Y4QFPNwzWj4VpIe/xoM7Os/R5nIOM=
`protect END_PROTECTED
