`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dY9ftL+c+DcDjhQMM6Kky7FMUi1WM1yTUWPnkwTyXMsMX1bc4h9rSe3TQCeTghIl
Sqmlzh5m4gKVtSA2/eXZTFiKZWUh9u3VYFztB8uLCRJbh24J97+Os+OA0ZdNtUaN
9zSskUuq42QiOAhvPI6XmKr2GT7FPPasPC5PBnUCUoD+ul3sfvUGdb3SdesLYQKs
rMTZJdms9Ycj2QZcpVQByPXrHsp4TC7UZv4vd13IBMtpgd8eL7kY4QNrI6t3U19A
pSggURoNdrVsX7fysp1LNXqRK8EECzkQ4J3B9MHkW/72ZLKUv39VPie4HrZg01aq
FLctGGrDle/vut3xzD0sTSdro/iebDf3UXmsafEC0WnZFVmL/mNf8n30HkOUxQ6p
QH8bS6T7JeC0/pdKxBo2iCOrm6M17dbIRqapLsytxeyu7CnGaqCWLygqEn8bzzvE
V7U5pC6M3ke3HJ/IeL6HP7LJpVw/fjVuE8MOEzTRCzPMcCaBGIxdvVTbaAUSVLrN
`protect END_PROTECTED
