`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJVqxO9rgKd0h/MX/vHOIGkMgJUluz7t0M/8Pv2uoojsQIEPJkGB2Av+11Lh3U6i
SK+COlBkofLNwLx8LQX/XwocYh653uLnvRZlCCpELWk7wKCfpvyv4yVAesXWSPmu
d/l7mhpbZfNVa6SO2iqVLILgq/eum8TIklYz1T45Y+qBpqWR8IsrAlEZvBH1swFR
C2D4PxbF44jfNK+BV/0oEQezek6ljAaU1pvyCqMl1i9mRlC6xUJFcBTdWCnp9JDk
Ggrrgas4t+R4RlZx1uXMXkfOY6xl1YVIl3A/nYr1GLE3ZSo1VS4t59gipRTeOPkC
02J9kwbdpXMeuOfzHrzrAzqlZKrYCaUJaKIEyGzWH+c1Oxl9/AAujudLpmEgfi3k
RQH36E8zd+LxDvBKoLCgC7FwswCU/inCiYeL9ZvF7IRDYDF9EHQOIfqmFdoQTlmR
ueTpBwh+/xSng6iBtHohxnz6nWZie9BU+xdC13g2z4fIAKbQ+olpw4vxGwcnrz+L
GvEb0Ky3WloL7kqsPkaLzoArgTaiG8zhiDFyayxKEG105DOeDVBwRGdux4OwL061
SxjWBbuBhLBHoWxgsMWooi43rybpI7Qn/IoxZLAXXko0rIHABpEQBYXRRCG7EarN
z/VMfszXRP20RM6GtdO7xXZJxRZqbSmJvhPVaqlc/p+JDOuCEb4NgaiNtnU4IOIi
l/XT+NNxqw3uz5qt+MLHkDiagLwSYJ7NZtIS9p7ALFA=
`protect END_PROTECTED
