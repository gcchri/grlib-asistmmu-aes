`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nl1Vr5X/7aJy23gYUGD41oMqMLnaqENylbZZmRjDW50WDZED0HhyUyqKT8peGooZ
HRSP+wOmvKtgI0YF3XiOLig+MVJzaaiS5Z5L1XpwE2vtksJ7S46Qt+micKX9bb5h
Fd8QecD0N/7VOvu23hGnfUzjMn32n2KP/mlQOLust5gbvCGXh/Jzcvgq2gEKlWky
A5cML1quimtDnAtKJDcq1NykBt3bpwH9b9MyFgTTgrAGxc8uPtSZwjH+MOYZ9S8J
n0qgM6lRC3XPh9P0Ojvuej42iqZwNOBASvVqL2RjAVP7H+J7jO3KN0OUaZusVRke
VbeIFKTZJJ4RcICi8rH1ssIhzpHQ325q0mNiRuC3QNui6vgn8t0ubrga+vZ0fcvA
FobqQhjTYN0QjIj71lqwW6r+jP/2G9rPHU0zgegplfan3njLE31VeIIJzDf22pLY
ISecpCN60LwCXiBWUXJw73UHMi3jzSZlJddTPq/Pb2FPzOkMYpYttJXnRRn/YTbv
RqCSZWjLhyvqTt7vuaHHT4SAjC1b1vGG91Bslro96PZI9tb6JIRKpETCiSa1Zxxu
tirRwQzywTKNGtzPa+bvfrSyG0ylcPX3W5wxf87I5m8=
`protect END_PROTECTED
