`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jumjkVGI2by6ZOAok1aVTNqpxw7XNEJoUllW5uAU1x7OXfih+MmslrpyrIFeB5z6
UdzzOeuiLzCMuanC5UzfYC9adiL9qHOBOrNQqgFZybhs2TRljCEUpTOVE1Bfw7RO
syqNVnk/Knp88AVWIlssl5GzmgdKqhVNK8OQLwmq1AXNNA6FyFsXu+t15hSoCquF
HTN/zW4hLP14oDl1NM6UsbTkRdE1XAmX48GqTc777/NB+tiJU92VHv6forNECMsF
h03Qa6RJPC1B1gFhEC0XXw==
`protect END_PROTECTED
