`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0vGcYwUwoFQEk1FzWu9pnnwIuxFvqi4mLt6sA+QwCFjL3+FOGcHLzKoCcwGz2EYA
SxtroIUSCLc7xiADMFTb6qBm8W+7SQu+NhYYGfrugy3e43enG2n97IJNygeT3CdF
XfoP1eKUvP8Tel7ZnRqNjT0oKdvdnh9Eh6UTtRPn5wFMtaA8RX0J1mi9mXc01Qlg
VMEVZKbuw4CFl9iFEGjBrE/XamBPob4FFE5s6AUyuBnytVy3VE4/U1+Ga1o0tjRU
6+iTJfoyy9EZZp/41YNo/XicNQRG4tgCSsUd9NXk4H7xR/4kEe1n7bQHRttDslRZ
Ga6rQWmT76uN3U8NUz+JkZJT6KxnMIp6HTeLUCPV8gqPplUgWMFKzSx044TFRZPy
X5RPmhTNiLaNMXShOXc1T2jMyhhVqAjA+TalHsnE8sAHFGW3fQ+Lf3WZohEcUaWU
5akBmG7d7LOwfoMhGnCYt5SWglBM7htoAVR9rlrAYKB+1vYxrcabQDEyt5q2pjmY
d8/qEiMp6SpEq3tupcaDVP46Bzk8CQAxpnjQV64bkhPSKrm1OWzqYpfMWyjdG+eM
ZAE6h8U7TVtsybbsB4WdyN/YiPj940t0pue17Mn6Wnj8039j6SRomOfcpM6N1s9R
lxPUzRGgD4GHqd4F7sJo4M041836E2xLAtxqmM9bha7xGjO7mohjDzAizk3ZMmJ+
JQxPdTt3AouuKduwa4kuBIlDqd8v18HF0/IPqgTOL9J3nO98qe68aVMjP55cNThr
QpalWwqIw16WXye7spXD/OCy+WXjPme356WoJ9DHOlilotXscnPdFWkRHktZNbBp
n8iIIIiq+06OcPKbi+pkbmUn3TvPqmaQzanidMxn+ZcCNjLmq7BmOPOxmx3d1Cfw
pbr48b1Ll70/460oA5VGSvbfQ1rcoiFABEv0FFB39ITW7BYoCTSuMb/P57NA7r2w
tmTxnBy5BSpKtENtsf+QlPXxab81AVF/DBgcatISzcGujxvRZrQtbotNkwbULr/1
29/WjbnIwa1OsTxPs53cSFUW0UT3ZXLm5974LQ5ZkMH09KN9UXK2pt6d2XtOqvcc
MAl+jawlrdWeyethQqUH96WK1zKxoe1y8bopwTstCRpFkzytg3yj8uHNh2wtqSia
c6vnNzzoQb1Ora4HYBkDu5a8yedUagW3IjUISyc5+sksixLnoqAzea9EH31sKak9
jeTV5tWsVvOTa8iz/iAwqaNgDV63X4g607BfvOiOaeNiFgxGq5Zph/E6wboVzyJr
cvmay29aYT/4igcnQ4zP4IOHa2HGlbtw1sp/hLPBLvo=
`protect END_PROTECTED
