`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QG7Z7sWPZ8qvH93dNA6/f/zJtPC7rGAOOmt9AfkCwBTKqWq0voOVuT/STXG5jD5U
Hi0VXDCp7W2p4o5msKHeBL5bvwKB2OHVSCZdC0GpsiWVcr2Ur9651mBxRhQZnr0F
5c6p2mo6+B94zz7JanPNNRu704dxMThVwRGe8vcKHIabcC+jXsoPqs8C77EpGtzr
y5ZDnQsFjUOmmNXF9X+LocShdOgY5w1N7/1AyNBuTvWxFhnwjxmXUnO0XP2gavGR
gIWvtnF3SxB2vbRTUusPKXcrzFP5apKdXMLB/VLHlaux0DqOFKdCTFMHZ0R1z7CA
fnU4mKobicVRj68TEISH7r4Qg+nN8Bcx8pqhfLqgykCZTQIJ4SGrc5gD1cs7Y5U8
`protect END_PROTECTED
