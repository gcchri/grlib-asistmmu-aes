`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucNL74PHz6IROdLTxjJ97drnocilQjYqFJvTgG76pxio7Sr+NN+QRL9eAy4trdNw
NR1Cn3e1623+VO30QfXOeigH0Muy4uQ7V4AUxi6wDipFycGtKpoXajprtbw1R/3G
9rB+NbODBmo1ROZSEmLrPO0c4Uq9/ZSc1srTtq3ZrE8HUI3aXVcLukOXcFWsQ/nd
a6vgT7jAZRS3uQ1sxaHTNYr3l6z3lZaaAfFMojNDv2B061OWQu4HoEgiAWR3snb8
Zw+a/6VKOnq+ZPLmdFlO7qwXTfOJL2TA4Sl4oI80z822GEOXOC+XZiAhoKcCbdTQ
icXmQBgLQkbwEGBXZAj+TJFNfzRpYWeIMzSSvvdAOWGzpMS+hbaj9dSAVa3LCGGp
5WV+REiGWzyqHpbjUKCdoS3wtC42KU8rBk0ZNsDX5p7UUFpX0MorfySo0V+alYXt
6KKRW12M4Bl2hltYTJT+fxxFmqE4VBzIrzzDgj+eGCKMPpfYOmePpECGOVIgVRwN
Uns+IH0wQCVeVx4cVKJwwjVEqUwWQ7vL9HOswLDzO6LCfSrEkX6HhyVFwiCIVCJT
rfggU0KAVk3eNaia4y0IYwReg+9yhhfFeqMdQYvEOz0=
`protect END_PROTECTED
