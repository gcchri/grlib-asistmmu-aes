`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BsKNJC1M9rBk7wUbSelI/SypRhgNo65PsOcxYEXYyDbHtwvLXEe9hjOinve8QQ3u
XKVDp7DPQW6L3u1e+yuLuDcKNhaW0GGtY5DwZj8FvHypW70WXARxbUnpgM59KEEP
czbNwjDMOjY3F4PLRP+6UsSnl0stPW7pz4dd5hK3Q+bYxpPWj+0CYo5K79IEZt89
GRVquDb7S+w8+LCiyvBYDvShnVLWpTSibgi09XkwIWyY0RXoW5HPJVf7kzNwHlJF
i8A4MiKAH1zF2q3H6br80/fBcxNXL6LTYq+uCdJwMr0IReorJxJwg0YYKDGddDab
b9NJf0mAJ/vabr9vRu4ZQobBxt8IKE7balEIkoIIPffaGG5d2vbD852k6Q53pShy
dFVzQNN1X3OhQbZsNe+i8+D//q53Qu8VrfAM+CUkoKauDtHK6CcYPr7d9g93umfV
GXrshFowkvQzyb2OTetRxjjA7Nfmq1rHX1FUzcXqbak1BSoFNUvo14pxLPUp5Dgh
s8Y5SsApOV8FAjkIKPbdlIvD8NEG5082luSiAS87KVzJBX8l9S4q03Ly/NrxgeOk
`protect END_PROTECTED
