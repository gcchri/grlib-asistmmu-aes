`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xz7+TvHBtb8jZAQ9qlCi7dpp1f14TfvOFQW8zN7xEROAjTkNQH19EFXVzy3VW5VJ
psk6duTuSD2ZNKia+jITr204XBOyau9wESvUNDDzTxB8W2Yi8faCBap9lnMhg38i
Lycat/uH2JtJO6M1Vd6T2fQ1sqHhTQPdwZ/pEFzKIqSRX32R9L9qkBvcI6nLuBo1
VkTbrj01n8gP8VYlH2Ggu8Tbb/VN+QLe05cq/CY1/iDahO2hDGguCF8a/qLtPwF0
A6FNvjCLl8nYVfNzer2oyw==
`protect END_PROTECTED
