`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
be/Eyij6j4YAUO+AYfxdQnHIKj994ViuJz5AlXyHhc0T2tRoSlauHIGMuIeHYvXR
H3ABxktF94d8Ti+iVvX9FwODZnEVdDz8027uH3YsjTQ6LQPzC23KbOzMFgFHxywJ
KWire8S/Dwm1uQAFo/sEIsSUZopd5+krSQitsV2N/gctBCQHh9PyBF7621XhdyHt
YuYn0skDmbZM4DX7j8A96HIVViA5RStk3Rbdf1ulLSguroXYzlrbVGyP6RR35Ep4
aOoexeUbCNROFhS2BOBuCmrdPRhrC91UWAtJ0gpW+lY574xCJ6MGt7rRScendIOR
MDMjVYT6+fiSSZS1n0+dHApVFhXShNFlTUqC5TaZIWyO2dUFNHyJAF+v4u5Rc9Hl
t/gTDsYSFk6CmDVuHMIOl2rQcUQinK5iGSpRkQ0Dt/0CHnq3jzZd1vjC07n8Ji50
aSjh94Nn7YKNZ3Sc2+LiYJ0XpxSQsFlD8zb5Q12U4JEvUrVCYXj3bcezb9l6qCo6
aU7W9gBAGcTm1jx5c8Cv/v3tgXgLQFvycH/yNVsp9JRMl0Zejm8tdMGSRTDD0Kxg
72uQj/X+UnI0QqyCs7NPpmCUqL+TV7uZ1832cbTwys2ABSr02VLhD9zUMKWhzEjO
ClOnnaECtSHPccwCoOUbuGghKg5Qxxbd2phT62vbNfnFqvPdj5DCNa3l3glgplLU
nFklQM/LWnGid2Eg1Zt4OBFKTqUrs36y98kN2XK5PhwyEfEY5avwAk0JNRam6OoF
0oOB1C+VQ/lSM0OtsmppvNO1Wyf2zG0EJ7vHy6FBKmebtMUE9R4Xu5UKUi3+p0Dr
b/u/46h5gMS6QmCs9qGTiB8yKmh+1pWySjavHsWQzwK++UArU9qTSPls2tDMf0uq
c7xLiVmUjlrwzm+9Rb84Kr5EnFVif+RiYuSRYAqEsTLa7CYphrl/CwikKWUcdN1n
+q+7FNHrqbBZ61wDq9B9d4SwW530yN9g0CTRDY5GLYJOBoHDMCXH4pNdpOp1Db0I
fDrstG1+tV7GTmljWRk9E6KFKP/7r5PV1E9khgRPA+OpIzOyJrAwN/rN7Ye1R2OC
dm6XawIoe25KvJP3yYfK7HadS0iD9NYV32lSD/r4Jks=
`protect END_PROTECTED
