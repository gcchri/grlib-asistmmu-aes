`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGeK0CqcbCL1+Udf10mjRpq94WiACvqGoDIGRecpK25KdzqUfSUbL42a7dLe4YkF
ThlAkH4yqR4Xyjebz69FTjUxQAqspsCF70e1jBI9kWD3mgrU7A0g8a3JnwDiQNOX
QIvVfrdgSFR7DtkNk8UP+Gi5TMQhV7zP4XTCt3u0q86g0uKQhwm+jNGfT9+TjHH0
BjI0HlvlAKoGZpbg5JvNGDv3vF565vbwkfK8W3vnAKNqbllUy5HTfPJKRw+jKS9T
s/12Lzr1xwTxoD1irz+zHg/nwfrypycT2rOQjslSQS0h6LhxywQB+Qv+JV+mvaQc
LTqY2ZNmxRjwVUaxJfMz8qLvO3fsoxVSKLIWaxYsPLFRyFvRevyGuALDadeeS/Ix
FwZHAUZY7kMrmCbDLV5s0w7Q/8qbGHinseaydhfKcJvN+1LS6DAJ0d8fcBO64G5q
0D4O7DxWjAZNpcYkD8mP8Of4UcK9KvudF7JF4Kh/E7QvdafNl08vsAEe7JreCRcC
`protect END_PROTECTED
