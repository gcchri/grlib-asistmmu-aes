`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6rUgDutQvsyg4rSHM9kIYku6p+MwbuJwANjeHzZxnKa8RJtPx0FRFb2kLxMuG5xU
fEsnyvtWGREFn6H0sDOkqAzxd2QYQeEYVBSWgqnZmgNdn5kaX9T9+VomWqfDcfht
W/1DEl5UZHAN+hjjMHTGe8x23c9P8Bks0l136/iiz17V25u0Rp3/wUFNIh2jdSR7
hqKNcIvHBn09Q12f5f2uRBhGcRx4sZQtiHnkuVCroToB4dwK4RJZncKwbR9Wwfvo
hviLwsR05TARzyeIn4sOJvAcAuTIJ9fjE5Xii2aeytD//gIFruOZE4GV+VbqEGfm
D+b+cQP6ggHqD81NTdYn3OZnQd1p1ZXHWSxktO4cEZp8oak4eQ6HwwbS8hNBBVcM
upwjxH6aQEG+b2xSFK0QszOB5KBDWIr+yH9szwDckIIIqKI1W3p+Sa+04IFvGQmD
4ALh0DjTqlNQ9nF3v4UvvLGFb3jj1tCRSj8cxQIdCrK1SUoEHCcNX7MvzjMmSobD
RP7Rq3PEx9y3hqLI0x5HCO19VFDSER96h46V+jSDmeI=
`protect END_PROTECTED
