`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5KOFL03r0cwmBlL/G3v5h9DAfSL3sv+s432Hj3QI1BydnSCtg1VOBJ7L2hS4GiZN
l3tW4nd0Gt3VJnHSU7JvORMS4n1z3fs+2zWsF9KWZ3dbmnM2j+ub0/wqGJoKtKlb
r3HxkYqfiJQZZ/zhloOcaA/kX3pmsVgwYCOijytGvWBmbAbPLePCseHVQQtFTvDu
Za8poeNQr7rHFYH5J4IMV98Zv354cHj6kGy3hGjVguRLXsSOIbbya16EIJAa85Jk
mt3klfPQEiPeaD2SMoLiI4vFXK0gg87v7L9iW+VTJ/zy0FMrFemDv0BzgAawuzGe
JCYCO07/jNcCcG7RDKOOFRZPDf0aDMiHBWSgQ/otTkE/iPLvO+kXckwMhKW4QvUU
GDav5vz6gaABchdjCtrZEgMMGVQZr1JZNB1gvxKWlQJsY4WIJe9wPR8aIHTIhGvD
WkalrVjHhOZ8ljU2zLO5CGJYH7Ndgyxmgc1L9Y/P5vu6iRLIolBnipTyYUWfXYs7
hIVXmUW1gvy3GTD6YtsZ2Be7s6M2e5gAcxRN9EU8TCGIP7K33KAXcSXSd7Iq926Q
Eg/QoQ0reJvHIEVXkiWlcDWiM0xHiknlHIvnkHRo0yyxFSj1n2ky/riP9F3k8D/v
vxlNsSnQi3rkBHyIFOeYDc9UDhV7/wWmnfeFHiCT2HLf7oF7NZ327HDTUYGhft05
Skh0dP0LbCxrcnaKk5udHMX5xrkwH+W6c5ztozEqiD0fCuAr0BICs93DvOEyWNOg
429D/Mefr+Aj1XIXkG0r470xBms4OguHC4oUvFcrItOCx8786ORGixcwoYgb0lV1
/plKzerHnzUxpfc4cTpWvMnCiKD87xPoJNqylEvmvLBrKY8tl1+2+RbwpUeT2Qhz
t32mSztwtqhCQz+tC7j5q+6yxzyKSUyCEUdi9Fm3FfsrItithIHMaJTeuKp+gf2o
E6dcSp9Xhv1TgR3zX4cd0HtGyk3BuYM18XwY68V8W/JUfKngV+JbzzGQ5Hzl7CWB
Zut7+1W3M661+kHg1LjgoSQ1I5EVvim8GLIPUU0KbaiNAV/gmEF1AvW8OLeBcNEY
ayXAadk+QWcfcKdqII183zMBxLuykytaF6wdpWu5C9ul3El39Sbag0Lf2kzX/M6d
lgcqstRcGJWINKniDvsV3l7NeinqSYN1unozZ24Q9ugGXLCVQ/XBsycnxkdlVEac
xoSBUzHkzcH1dHnSQmqNGN84ibUmAssoLv0yEcV+r1BSzv6oHHdH2xoOUuDmPX7u
N06CWYVWxDyOgiypXZwPVGVVYYrKwNOZIWklFklOgyyuVqWGBKNr69+GJud+un56
io70tGbCpstWPzka3W7QOrFYczVh16aK4kalmHvlsNII7EkLrucROCFEOxXmpWHV
OixBTFHPxHoQStfaJtAZSjJrQtYGy0EqFZFW0/tCNb3p1TDMhg/TwORW0wDMvava
WHsviFjr/Tnc9zl5lbnKz6LRw/jRV8Ypj0kXnBUjhXTApZZzTHAbncZs3PsYWoRG
vxhPlG4D/AoXMlQMT2pAZAu1MP6oOAdUr8G4ZMd6SbKgeB+9dU+gXtlxN2/W2LZ1
q/XNdWGBolUGwUhoVCb+5ZB3fVJLkNRhHl3Q7Ao3tyOKAG9jSH+daVFurBkroIYP
dcRUJX+fXJOHGBnjBcx/l2yfDo0zzwU8m+rdvQdHYdkF8q9RzLO51R0CseMVe9cm
eUHFX8qFNFvu5Cc5PrTg6JXptSeNEW40Rq93zHs7cL0VazT1lPN0g/YRTraIrekz
ScGOtn3oWz/0U0mVFQz2FiBgQQrj9OquJQ5moUkQOsj8dA7Mm9hcOsEApCJe9VQ/
9jqGkgDXWKKQrW5xKoGl2FGrU/u5qeqIhfI3npOYh6LTsGEkgNaYFOy9VrVpoNJl
0zM02hit1A7ogOEPEy6Gfqcp9aPcKx5v8Lieeovtbqc8Oy1XO7s7d8lV1qzhAMIp
SL4j4WN0FIWLbbXOFqZnOon0WuYT1teoiniqhj6fJ7R+OsRfKkHlpmmOq/eINmUg
Yncv/slW5Be3UeIIV1TWIL89LjM2fMkAJAcM71uzCCPzWhuZoszMb8EO4vYvfLz1
QriU8dK8/22ZFCx5ip9UjlNQ61AHbKA3R8byCJGCaJE2qw9G7LECJOmqGLHrp0V8
QTJkW5PrimRwR/jHYepSZHvd7J5FQ7Vfwi0+p1r96CX8dDjDqBYIZhLNTmEKuG19
BlCB8jcGKTHqxDDjyIfzuCqRRSDmmdX1+hMiT9dDVrhAsj2/2L0Hy/UyE5Yzp3yq
E1OGI8iUj+BupaqttdqSec9FvkQaN72v5/26mcEdW53J+QPpLsE27Rd9VvR+58GY
cF59h/rwVOdir/hJNrhlmmIVCW1D4j8t2bL+BL+HwVo+fxj4/YilveOGFXk/2QAk
IlCNm5WePeAtL4uYuCT0U+iX/dPRQqwfS+C2f47JMmDqAGhYiHw5XWEIkPS3xgnw
1+ujNeAV4EsN3PTMo7a1PACv4IrIcuHjoOrBNKREceBRXbwsi0SZwDWP/lSCrAt9
MYtie1GIfYK2onrsJ8mVqqxie9ZivhIZf60trSIa7T12zngIJskZNsq/5sPdb661
o1PCvuVK55sDLKWfb+h59lysjAzId0zWnxgh8e3SjjOJH9EX1HorGxL2lG0uyan7
W0J3NXqMmGayQ+z8kF/cWLopiiGWRlF/oh9kJP7IXKvXx7+/b1LNJSe/Q0rew29p
F6S107ZY2XH52Nkd8kWoPcucH4SNPuCsLUvPTkRjeDLf6Yh2OD9adMnrk11Eoxxr
1x8bN1wdJmwbRxQHXCmoxvxOKjQywCctjwFyUMP5m5yDrYIG1W4ef2JkHpr1MwHp
HIavGo0apPIsZ28L73JxUyMgc83Yz2MJquwwf3q6bJVHztd885BdlX95lDQLHHhW
MKB9TCNW2UZYiRLU1gdGVwqpf9oeTzh5O8Str6CxP2mT/mo2gZ8tm5vnKTO2pRy0
ezSDzLCdfCrjmcbEy3gG6RsT03aH9GScggwx4TeU4FWe2oqvCfeXCeWLFkKx1+ci
FONoINaNb5Ys9U9OTebCBOfRdsRy/kzouSjPZNeqST+yLPPBqPcgd8+D0KoqIWER
NlnCHtcpUh72/vTdsnHTXUr8aPrF1NDstCLkpvsznC7j7LFYUlvumSqRmuNI1XnJ
ra5dr5h2w3KvRj1ZHyyml2o6448c/JI+J3ICemIWW8oF/iLGi1YXVe0kvw3mj5Dd
N2MExiIq7n2NIRgBLflgJXi4vrEKPc0BWHXl23jnLweYmKlWD7AK4NBOi/XsTHxt
hiTTFmqkan3qGE8ApFDRe0GnmNkaJgTK5iwM3DH5Se8hDSJl4HtWPn3ZGaUn19e5
1HkfNk51lHezNnmnlIHxqT9YpeHOrK/e3OAymTLE+Cqwu1XJ4XoDh7y3W6OFhb+P
O716Sbt0wXeIuxJg+5LeUrhOwM67+sVLJx5nLmhVe8jExs7LrgQBxWaLl5Kneu7E
A7Q9f4ImBBD9tTkjj229vWL41q1U7glg257o3GTy1Edc0V8wn+lZ7Ar5YMF/7F/B
iOE4gFWFNSf4YjFAtVrw/6YwhzzWAiM+2D72/JU30Bd2SyonEovpeKh3KW9dKzqx
6NKvEPOIe5m4cmHCZ3atsaXdVsBbO4ER15121QMyO3Va+VlqUEM4hspmrP/finhk
gf3g2dbDWPjNLJHPhyA8P0CKcJqLwoajAJW+BYyLquWz94ucaFL6K35RJLfcgERB
i1misLM4R/XzbYd0AD/jDl3Vi4uVYB+khk8cCfDfcEA4jpGbB8CJOZWnoZjPn4qY
d/MkcKTy9kO/sz11aD/CnJKNhPxqdf0jOgy8NL5Uzj/ymNAczQ6eK3qbupqCoCg/
0xnXa7E9hAHpX/ZAgMvyX+MAGM4kxgXIliZbvmIXwfumU9jfSQLQbA/3NwrLMo0f
yVDXjJvDau2Wimub+TUX49TX5AGXcZs2EJx23z+pcSJvYewqASvE+P5WOWZURG/c
JI1H86aTAssb7w0QS1/zBRxgQ2PPms/e9Yt2O5GwVCIKhiAjNu0OSsoKVtazu/jB
Uuo4lYZklq6tpCs65e9xaqUbCcJwp68jSAgfXmAssTe4oS4oNDcj07UBDUH6PeX4
gJzTTDSZtTLw3FEQ09jH+0rPnk+VnBHwin1lsMdWGACyms4QFkfLLnsHI8y532Rc
Nt+LPCHNjQYCDmz8FHgLw5jATasLtWfSETKZqHfLDBAjJ6TDJdGJSfa7QEkTj9e4
C/78Gbea+4LV1pjPIkAQBOU8ZOiQ6TgJ8mkEx1IwSRDpTQfWMSYWNv5/2fnJwUgF
XbgqPRUrtw7ahRLyw4QmS92dmQm76E2cDD6I7DetCFwRruERNBk8e5fiQQVasVCs
cBLw0embk+vH8tDU9jGUsTPWt8+RhsEndibmy2JdQuXyVvixpCPo3pm6CgkT8K8L
U/wyhZ+GtwwmAxDvoj7kIpKvxnMNkLIdlbxobMgDZ5XA5KDtVF84zHcj/OlpMejQ
oB86Wt5/6LyTZaefRg2rARW9FviYU5/70b/CHsvmiO8maxRsqH0rw6oABjitGqO+
cJOBet3Bh7Ghzv0N6JJhygmQvAPeVgVwuBSg8AhQI23/2JImzaVAY/KfTo2ACLmf
dAYI5dHpkw0nqA5xxOojIOblY+c26JyPl6bGBBiCbex/WtUkGn62QAEvdPfq0n62
oEBDK/NPH0bxrBHmdtXJm86IAo/UkJHe0eXxIhdAu+gmAH5ACIgMQlsMyX+k2Icg
UuGVfEoOeOlkR3QqcnLZZl2J+9m29GBKVv2hLkFFlfmo00vk8J7k3mLGpCjYQLyi
vBHK7Zj2CBA2DtJVP8By1MICFT9UAVXiV4yoLu5mP6GB/ngUqToCs9MSPaaoDoCk
iXr2zb4CLeRcnJKr0S+82cjMuXaTfclSHCt2TcBj6U27DbGkNSACMox2J2bwRWfZ
Zz8naw/BKgBQFus3i4Q6inc4blEOOwGYI0IAN8XsZxqvyElo8OBKO2P/FnPcMg9X
R9gpCH0iwEzVQXHp5zqdlstkIESJz3JylhXzE062egKXGCmWidw/X0EfyMMk7m39
Y9izDGW8WYbn1OAxyhKYWMURgcmI6xtb3uGvsSn9VvNibCvPSios37hBHhxuheeT
Nz9wQEixnnDvPbKtsqLq3jg6ZGsVqCsb/Rso2t7adHBQR1kkzl7/MLNEypLY8ogz
l4yAsNWDS4qUww9J//200GY7ZC6L8u5bp8YDbfKdHCM68yZYir4io8dxoICBH/x6
T26fOh49+zcnRETlE3XZVK2oO174GmHx1kf/dpHl7eo9TPw9qo2IcuXGgVBnQKRo
71qgkXnilnewYmHJvrMR4QPTRo9k0EOZ8Pd0yFMUK4r/jRn7QMml3E6DVr16Cdub
ffhPdrwBX+h3WZrx9fRsPr+U7Wn8vIoO9R8NknM0VEjR/5dU0X7W1irXnxxPE6MA
9jFidcVslwdQ25Am3M1kDHGOfDsX1vFGazuXomYjwmvCVOLuqTHFeY3fWfo04OX1
GMBwMprtH9QWgBkRo6dp9oHIHSDG5gdYg6AUNKh1ogGgK/on4zadbQWGJ8vTmKlu
LUHPQq9tWJ9nJTRUD5W74BIMQCwo/e6ffBBQkRip9VUrUcck9cZc0gkyiLFJW6Fw
KxByhKuz2+eVB40QIGVBu5kUGVDZPPd9005TFNQ+QXb+MGaNblkqDbjHzhoR1mjw
iDam1ukVbg1RcTUpapGnK2lkxkntJVmuC/DpB+I8/NTI6Sv9IQiXtMArUa7rRKIx
fY81AwsvFGhSzh5flkCPxZiQqPu3sdvZtod1joDcdx6kBsBmq1GSJZX8gxCUGwFl
UezCZLzHYzxhJy2vFmfgsHkAo08yIr98AIX/p3u05PSUdooYWSPKYnoPOXzmqcja
MPuvk6jiSuzNMYbhy38bIxhVTHD5Knr1lwie5VnSQEAku5dTz+YyRqZZST68Reke
8WgBUHmDePGR0LgtZu9mTEVgtvMvOQe4QQIzb8fDJtBIYFzGGvu2ohESjyfa67SA
gMzm8Bd//KGi65GPj2vUcvkL1u5HD0mUGwQQ4W2BMAt8mE6spUA5r7u9n1oXTmVr
ZhEvlzbg0DsPEPMcpO+uIZk1QTvRvvWhiAtrOc65zvbho+g4mlOMs2CZn6XlEHbk
GbPJiabC64zgEk2d7EtH4s4imAFXJqyP+yyf6ytjPsXdsPH3pgouaxPZlP7eLx7o
9XQtVlykSIUioPGFaegpRRX7WIR+NyjtPzFKGQPDWy6asqQfXYMMkTQMTI3H65Rz
Jx0myOgaWpiWYHv17GRxio5alvBASSile0vD3Yunb52Eh4MwOFJZ62nXQbp0JF/M
`protect END_PROTECTED
