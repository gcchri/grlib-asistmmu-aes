`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdKS2bno/Y3yYQ6o+acfAyGIV27szD5sPR1VWm6kJ1CuXjB4tirDPLp/GOxP5uL/
kwx6i01HNLbTEe4ToQuNiYIEsgyOER/pU6AdbAAho0G4zXo9wrAj7s3jvz6CSXRN
ubid4Fxg7QCO3jvtDqHFujNr0IkfeNDYRoQrx5m0o3X68ttH/68sIQ+3muS7VUca
ii5MKy+NvLF1FNecsGVUFcJw3V8193e0j+f0TuaGV/cM6qtQGitEhwIvUvUW7mqY
IkqFrAvoZxcTZrMdtII6AhkzKpNyxenZZBZlp7MF9mP9Xr88od3dAtKx0bD4A367
Gt7LZGxOt2dVDsghvG4WMAOR/qdoX1coen0ZYP5puXD7Ac8TU2FXx077DRL2m+Um
v692/+ZDi3FWR4W2yzQaRdqo1sfuQ/DjFeUvOrjJDoAacBtjyLaxmyg11YBJjOzC
iSqrfUITB2Yqkuy8f/S/caw4rSc1XXXNgexHsbID2JmLtWoahdf4Pi3p1+KhDqLK
F4uLMey0vt4EolWylVucbhRDafjYRGqFVRrJ8byulkwmEsBLp+0YoEAyCKqwe/4z
IV/TUNx3XWpyhyN3H4T9A6UE5zm1I7IuTHiK01vyYF36njHWzg4mvSQ/WLpb5015
0wOQXDrTgU9bMi4IbqDN4CX3T9w2Oo5r8lA2ZXysSpI8OtpuHKMrrPFm++T0NyzI
JbytpuE64gp9aogKWa6DpV/FWtENX6PLb8G6b6E1jRnyn5tFWpOWN0BV7xGELZwK
N74iZyvt6G68Smk4dak42Q0kr+TigjAQXUK34F+N5tIE/cBNWMlwAnXaomSZyZAi
5X17M2K1ADYp28r/oqu7bx7d4BSIPspX3vAC+wvTncvv8gFo+vi84lBb6zU3XEp7
ZxRAc93loqXCvaIf7xYpjA==
`protect END_PROTECTED
