`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLZxpZ31sF7IkO0quc1ozAZlGHFx6h7Gx+SUCV9+zOpxmOlklAERLDV3o+2TVbGP
L2DUg0+/RbEGR2ufRGu9ocSP9ax0Y3d7unXeRhkoNgMa1kOqCIe4Ci4ROLlc5Urd
/O8mXR6SqiuT+FUTXl1jVEJ9bBj9d9KrXdZGMbqoAUkOf7ukszdPvaRmKJ5kbvdd
oP0U6mjlEUGFvd5f83cr63A8geeHWH/OeZbTy1bJ+eF08ryXD63rDoXoKMyjA7+t
g+wNhsALg3JP86/avtVs0UwMMmjkpS/O+zPDIsCPapPPHv5cK6QB30KDVRCQA5zw
G4BH4an/BtzGoQM8IIjtxfca9xK4ve4+Yn+40SvI2IGWhbd23aVBR0bBy1++VJwJ
qrmsw39LIX2irciy7+BITAnFuEkqKKxsldgcEIJnRp4=
`protect END_PROTECTED
