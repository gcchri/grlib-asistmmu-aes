`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4NIkaQRrOFOLqQSbqdhFnj2a6hOgSzGMXuD3nKwRP6oQNPvgUQVWxCkd8E/TI1C
wprmWCstje+SbzCCYW52C02vo/ZWS9F7wCrR6BRijK77RQI67x+VLP0CTmsm0Ysy
EbNXhRhApnKoMNS1d0iOcNCLuiAep+JhOxih+FvDH9zHYnLFqKjsiUKgpXtAOzRQ
J3j/rC9Vrgx52oRWPhaU62r72uBsygqEziZGEOKCVuWkb5fj/0uDoha26Q2tDE5v
8PsxVyOtGVgDnZpqDrUI24shWkU26x5+gfdpvR1mgGU0ft8/EnCtTl+EIk196iWJ
D9gd5IoOzdtRtLvLDO696BLPley8oJKCYvwSFSKZFk+st/fpLPPM3h/25+JJaz7R
LBReyrDjpryYxGqLYMUm3Nu7lBvYW+N29dCE8pBleHpxrIhUJeiowz3BrfQhHMbF
TSoMPLCAL3KtZzAwltR6peXcnRPACBm5+QkAc05J+7ZRkxMG60zBY2Nq2CLAQxb+
LGnpHkhvlYJPhzdEz9Dz0kN2N79ydFQPx5KrAPPiYgIQCWSoz9pmLSga7IlUylPa
NLxdDHH/1ZrXveczDoDSF1FOeJFFyiddMiaFZX5hcYXeTqRwKyg5kZoG3vAPxlnV
CHgpDmm7sGLrvajWDDbyGzMavfT67My/gGKjX7kQMVEIJq4JM0EdXAsllCSQ7lit
e5uJo2HmHyPRFZNSbgGuz/5lZN9Yfao754/tdgG8bKkcWTsbEpjYoPxU29sDkQEE
fj6VBbpTBo3pZUj06K5zfntKmiMef3iQp++f2hhWs3C11vbZn7BkWXhiSGOZRfwc
FoLbtxL7RBp7pRraMnO/+gcpXLCEpEAQ5/zLYKHevxooJRFYT3v6apsUAR/vchDa
KIpLnnF1eZwaYpuDdGP7E5XQEWVpIS8KI2QhNLzyTXvSN0Kxd1qNTVtc8dyd8ctR
rx9MevuKFajcfS36Rl/Tei9077ADxUOTZwkgrGR1YLmc/JCvz0Y0ZVAdkeKqIHyd
l22AlXEUHuRafRdQkrtz5pYUD4ssLk1RaOsqqYFlmFGYvbxd8xkvVOYa329HQonU
g7w+Tu6WX3FZ3oTkC/Rp4elPVpZskTHmn+ijZH6eyJCKS5YgNvrj7KerJue8wwiv
YX3Vq0EcZ4mMDD0jciUgmu0WZIsO2HN8rFAUgSClvU0TGmE0gEnnGbEBGg+IHqKL
1Fsdon1ZOzl9yxaySxNUuVqXxlsX17lGweXLJNeBfwKSS+hi7MSck/ztnxeoTR77
rbuXm+SrUBdqNvUGr4iSyDr9zs88fy3834PDEalZBSbPTesmCpZFJrf9k3DNDYs3
gxc5KiP3bjIGffSRN9SzXqNCxPJ5eDdaA1JEQbqsls2CM03aQ6b8ZKPLZf14xS/w
Ih1aRH8ZCAo3ir6tnGiYGLHhVOt6o3bz59ENx4XL7+KsGZO8W9BofvlpB7bvwVJB
VISTDst3GIsUhkvr88hUkJ8XR+bAjpQwoqoKICW4rIto/sv3EO4PaTO12yOUIH73
8DMdb/na/V5ocoxsbFmyFaJ3kEHe6biVn0Ti4+REPOrMkzV3FyE0ExsHaFFCdMwU
CbxDkFy2WeSLmCJ5v5RMlFDh2XJYULeDs2Nvw2RW57GKha68Vv/jiZS3axsTHqgz
qMGgCt8AjMne2+LwbhCnIxAg14RkL0w+Js7GqqJibn6CZs7s+Rh/3HlGYPwHX2vu
0YqHsvB8ERNAzUWgDTboHKedIi1GNz3Bp808MHWZiJhXQusdXLIn4YimoPaBGJOr
FCMQxtcqFpq7E2dGvbTSXCk7qtupDe3XCfY7YwyhNYoyqnsBlN9vvb1XL31If5Yt
UTI6VeZyUWIitrB/9W9LqzeWb7hneGc2fEGzuHNjr+cdUO28xTfIycjqLDgs30re
7gd29916WNJvPJ1DLUJrArTqP0CdUV9T02Q668wJwVxGwwflikybtz5JpAEURHko
x6UHhNWHBsFYjGgU07hy1DmBvHeX36r/AQsbcUTwAF5QWHSZDbGxORjsbBtedKT9
pKjMYK+7fdm0IXdv/H/cBG/paNOLaaqXlvXPwgFcpz/gPxqOe2Wxk+I1l/XeNTeX
ePatJ/su6YOSFEYYPFFSULtW0371UYDYBvSOkoURo29uliZ3niJkeDZNkFmi/5YI
sMFYTKBS7CnZizK7ydUpjrHiyfTzQW+hCt5NRRTkivtn7ubLZpu9Osjt//jxSbHi
4O9JVzu8ihxwmz6jd+8b2sIwDPOvHgQ5aTURAbX8fvM9yzOGoMZbcPJy9e/5pBoA
o1qo9ZgG7TTjpS3/CIF2R3pFJU6VcZ2HZPeATgQuJtrwt0zYqopLW4dFHYYAFt32
mNQ5nd4lNunt+GP2rvE0PO6L4kmrEkJ81IpEiIE5KZHOCXD1tSphv3oPiMQMP3qb
thQpw956dSPB27ZV7t+gQ4C4qWzcW3om0BwHvU5xepWfXDbL4cja+l7eRVQ4VI5B
CqXJSDTGI7P2k98wSiPSnlpf5HjXXDyIvgkfetS5PDNpUP0Aq5IZZtIQaGWXSMUu
7W9HEH645+A5haDLiF3UmDLf72VpPomXqomrA/Vk5f1Sfd6ZK3UE1zRhUcPIqrsM
+j+HFsrAugAq00km99GvNv5drJqKVcIHkY6v0jgj2quP2kk7LEvdtWJrAuosVY8P
M+hHTKQVxK1owsFOJJvGL2qYf9sAuC8Wqdm6JxlQOuJBX/enMm6G7z/Vo9OyYvOd
cUHpGfPm6a0fXY6kQqykABvAURjOZnIQyBq7RHTeoAsCsKSEvZwpAajvNecGbt/r
tfAZaeQ8uRAYNsYWsCkT7JcREwrVGyRLZ6AkfLMywQVeE3RO6dVwtmj041yzcuE4
nSzCAXXiYmAPd61KkC3cB/g2JfnajHlS7a5ousHMp/F+NzwmAD9hJ2pCt32iKUkO
cAfq0B5FuIHXYXdhOkeBlAMh03u5y6vM7lGTNhYJS3QArqQeilREcLjrIyV+sMU7
uRtuGno743CmnFAz+osgLBI7IuduHgJrWt9E2+hzVCmfICtzqk9h5wAUhQCVOfFY
MLbcr8BWTjCvEywXQ7mSKpn3Oiee063g7v4gLbSdJq0wU1oOjN426MRmsesitNBQ
6DjdSY70zLftf55VJp/61AJH9ZY7cKEwEivfRZ3Jn0U+G5I5TZdN7H7OYRRfJrWF
Ijfn2wSx5iBO3p/J3UZMqzYL1nwxnIrDOKzv73WLR8jxCPOzIN4Hu7beJd+JQHun
KrQqV2DhiK/dkwm7LAdo64V6HNGY5uGFoijKA+GyeEWajW0a1dpWEma6kx9nVFBD
CtPPmBzt+efxUawD4gsnH4Msb7r9sbeKjSOtB1rL7Xi5vWV8ig5ovYRnBy/uqpVK
QyKQnMkSM6X/vqyIE1UGYZxsI6kzWm6jO2EP032Y+UabvezAKhGUpAp5jAoSHp9l
JdhzPeOBvnBwYg9Coo84BKPCnOfvkBeDnySV0h6yfMOGSwuPCuflv7UERRf6lWXE
BOUfBjdjx9hYmwvhpz/3nHB6QNA/XGeKAhtYm5hNGPsEAnjSwymRQzDPyeez+Vjx
4b4AKWs0vEUrePCBV06BeSM7wzW0HoC8bCEDeD/H9/gP9ummrlw6Zid4VDHtC1z9
m1vjYL+VOh4Rl5Xj98W0v7EOjt6NmjaGi963dAc2FH8GJ25Sgbmls+gIPKyod81z
MzYL/Q0Rp7EmdodlsdWiVcTyB4EYDPn8D6ngXrqQpJEA6W1EkLKKVk4E/fYJSS0J
YS2AuNlUD6xbAO3SYL3s7rGOsJafm2XfsISCsowBZkzTVeiNk9h0Y6RsYUTATE3E
0bJHF11E1l85clW0D4VZhryl2b/k2+hQHREZOgebTcPH29Ywg3RPVMiL9cv1KP+d
VTZV3KU07Gif6Pk+5UDlnSQ4bD4O+yP1OksUZmkQXll3K4o3/g+Z/S8XO4DryRW0
WA/zQL0cTLnsmX/Pp+ISug1+C50BqgZ0LhnYgAEzQUHChGkehFLuQw3stcNTIw6s
lw8J0xO8G1hOHz6Abu1aKi5JKtx73oYjeLokHw2vY3Ldhe3/f24qJ/mpurRupA0o
3F8mVaIINAQXcGb0WUpgxgjghmMl+VNEiaPr7muYFi1JdtgjGp8Zzhu7NBafHD6P
5jTzPidoo9cV3WfS3jjf3NBZfL/qmV4D6QJLj21vCHgShm86mapwqMt93aYVhDBH
sjOrNQKi5zNLe7XFFJ/iQFYU98jU6F6FQCEVnVrodeQLioIGqGvAn1z9Kf0dWa/a
yUpqLKYvjY442e9JihypdSPAL/NP8qMLnilz3sJ07/8CLmYjKyMD3l/cQ+Rhcq/h
cHu47UQetc9fAtTZ5L+IAse8l1HUcSWkWvu1RcBvBV6jE76c99LHF7W/8n39tsEI
umBJ9uTyXMoVlKKQxpd6b4vBJxHd416+IGy+s6XsvBh+1cRAShlgLClBzZHandaw
7U4JQC5ATruKBfFhAG382rsEoZLM0t0gyE5M2ahie0gJ2h/bw6xX8xAHGXtvEbPC
VkfUpzqu5Yqg0NfwsmtBXdm+JR/Xt3I2T+iUQ4fscpPqblIs+m1NVInjalQsZYTq
R8h1KsBWbDT18dcA0FgIc1XJcX5VOIwF0TyUvccKFq4KpQHnqKIKP38RxPCPZkpd
bO7pzO2ubGD3yY8xNkmsQJE5MSSjcT/TmAv7ZXOGtrtCUlNkSQxCcdKPBGkoCtnL
iciYpPulUP8QkRCdSfKgr8AfvWpwhH/ous0YJ/htbVTRZnlbAnGoj7sqNxUNLpEM
jCNQX4YHTHy9X7F9QlO6zJj56aQM08kXqpT5t/GMbesFHh3dK3FBe6xim0U6J6xI
JJH0X9yzdrkCAXcIZqXgDX7HvqReSJD7pM2CE9CPe7Q6JzZ0UWbbGQEXaAVVIHgp
w815vkcGRXVcadyyQ5mD+YOyij8FZ+sVLU99ExjBrR4jc2lBfrq3vuAVfOzMNgNm
B3K/tAQBksY8yU0czmIbClrBt/0reEhbRTsQkzE6nEcP5GqP0Eg/4Mc5YgzsG8fs
ENb/n0A03540ju/Fw7OA5TlNROf4jZ3ET+th97kXyAYOqVOrHk0zDyE9llYHlyqe
xzJZ+8GhkyXRrk0eKIDsZ8ZheN/woYnDh2WK43Uj1BqIy8nL6gpDmSCSZFpohOZJ
d74hmVkLtdmJ5kyBZERXCBzdSzw0VXwQle3BZlY+CcsnhFLczjdcHFEROuXKBFJN
oZWY9B6VfeP5TM9sQAXEHOiM0olXasJ8QBytheNCwNFzMX367S/FkbUEZeny2FDo
mPc+FNJfmywM7zjfBWWqNKhheysxt61CxdAFWu8Iiz++dstapFDc7XAbweY63WQc
RyxI+sbJQt3oLufk3iO9Mq9fQzUziVKpA8hVrRmcWY/fNeCrLOFqxzNU2wYRXAPV
9vtC+7d+Xp3X00rW2SjY8rE2+j/cIY5boHF91bPT9JQCnnC2mQAYxg/ZHtopuOBz
XjrFBG9fpbrf6eQQ7+AVk8Gx2xOU6RTkq6c9lQE06DjbiSxwfUYG0dvHShgZiF0T
Nc1TSdUgZTrNWSRmM+nX9rcLmDW/XZLnU8f9+2av17OxGToWoNnB46oagQXR4Y9x
FKtZyOFjPWLuoiJVDxYVizaag44YK13PNpQy7JJEsGOMB+7WvStPTfEWoWQpKoPo
9ksxFL04gOcxUbPpTHyqCnzXQiCUFfSzWJi2itWqm4sKlmozpzpQdBMVaDF3W7S8
l7Ca1aGD3Z1Nw458EjcpMz+eo1FUjHy9jhAW4uau1RlsSTOVE1uzEaDV/mw5Ht9J
J1XPltXPgd+7a+PnpwGyHxMJBStITXqEaxy3vQ6DjzVDp2BT5mdUJIVYGjC85KNs
qC/t9ftjOZx+dlM+WbDAS4i7GmQqcEsZhyu6ZaaHY314eROp5nXZLoLGOmNFnXPd
orgJIcrwzaY6kGJbfFAKeoYfRXo/STesfVu/KvQ+sPul5joVJbbO1ypfYi2zFwqk
`protect END_PROTECTED
