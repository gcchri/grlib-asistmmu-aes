`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gHFhU2G7Aw0n9UfaaBaerUFR5iddw+D8kNP0oNAakWtRi9bGpvkP2orjhEgeGmB
mtTptDJZbfOj4m0PNzXDn3Xnbma30sNgkqi8Vez7OQoBfmiQc6NB2vo7gsfMqtN/
21x1s4bVRge3jmDWDdy5SgWN7sei8VsSoLGaRs0mFTxN/UzXedNoPecbF4xzou1b
q+d7BCpKiIkYZja5fVvTytl8m6+VqFieUz6xlnVLLOLR9+myLiafD8kGA63/3Dy1
ivcgP927iq+gB5vcbkd0sYOiLnjLcBsRZGUAWEWr4JoNNvR9edwK6paTmLhETYE8
yae7zX6e108UlSnaBj7MVJwF27ovgaN3G5PdbsvKfZElOBIrD4Mv1Vt4kkoWUDv6
prDQWcZ7ARlwmhOWoYapjJn9oEXuIDEwNUPnUI9frLw=
`protect END_PROTECTED
