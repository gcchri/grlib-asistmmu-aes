`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0OThKc3jiEUpWA4VuUL4kY87964WXyLXUvvhPPTa3yRT353Rh5NX6+LLIzNR4aSP
S3EX3mMDCl75TuQKiCbjRmdZVxza5RkTr64YTjG7b1TN7vw1MCQ19d9Ogwz+ENO2
pLd992GUsStRzbhJ6ILZbtM7O62HDxZHKRgNNG27WePF150ySXKwG3+0z9YOjn/n
iYnqTsaC2dmkV2/jfA5XwLtMfSxxwBb9p3TdIxKS1sSUhDRYnxftfqoMTtzXgcMv
fxmjghxilIX0UlphWo74hBgLQUj9M1o9jYj0CJSForbR8QM/fHa4eAob2DWW2I85
kWObWCWy3mCx+Gk00BV0ANpZr7sw5BcWrbFBO74ssKZf2d0ipBPMwmjhdHUI7QR7
YyqDkwKdXbLxZZaTysnJVIS7JeAN76V8MFA5Rr7KN81bW1JgCE1tlsHLOKDwEvr9
Q7UEV9zd65Gzeh72KeHL/Hev6V1BYXJ5BoUxXJnFq06N7wp0ngOhqVKYVGgCHX7n
wY0RScqyOfUV7mFyPJ5xid9HcI3/yq3lPosABo3zXQWopcCNKIBUvEgxxdimr5lh
nGhaZJmS8WLX6eULEp+YOx5Nb23/p/YmQD3bb4A272jUHjB7cGUgWKHz6/0GvgYc
vYxXN/QgLDwYFIm3e0HBsLuizdyE4f3wmNQsGgMZF+rGhGy4g1zVEK/3leyMk5k1
c0PV8rLyx1HyZgAlyH3xuDm2OtdWTOT5JDmnSFHBGZ6VDzLBv940tZdWro88D9F4
S6JI8tqfCldXo8KWiwGqGqtxPdbE6eikZ5lfl4AQT6I=
`protect END_PROTECTED
