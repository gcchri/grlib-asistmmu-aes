`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGC9qO4G8QbGpZ3rT/IzuACcWz/J+hN087aTLNx+6LcADFiIsFdOx07ZZtUh3bLK
QPOeTsjVcewBJbRxj+sk6VACzhdb1h55tT6yHdF4o1BMFkRca/Nxh/OQ4nTegFap
YyP+bzEj8s07dde1SriRJQIoC9ISj/OdpenldAk5AE3nmFCc1t4hgvuaV+DKbzuD
o2duGIFMuIV0D5hUBZFKZBFlU/fQnx7AUENETSIsRG1YhQXwutcOWYeMztf9g1Tb
U/jLpM+i/5rCb4HNoNODbv+RPLMQB7iZ+MwR1eTUuUsaOQiO9re0+tPopnH+KeBH
Grs2KOS7lFf7TeKDsFv/wgoCM3f/FeBU3rITe4a+JZGxfgrrPfdRhR3wtFrh+vpu
CYZ5ME26eldojLULUZiWtxYCYLRrmRC+0f056xA6nCfs6WZy4MCPcQNZQ+BmW+EP
6XMrCAi5tuO9iu5GrBfjS+KAXi8UfPgS6RKdDmX18r12tDJ7FiwwaVcttZ14/u5E
8Bsy1ys1zib77AJsLJIMUFyuWmV9PJuK5vJhjGPl34aoQOqLBEW74CmglViUNKTZ
xwAHFVWzzXEv8xowzbAuMUPa7w2zU0Iew+nCVX7k3rcWLHbbug0wGd22NyuD8BL2
kmUgVupsDnDL70gxbTQOhCpuSAxqXM6soLcmz2bzLV1kGAnuYs7CZoxCJxHJFHOV
wrbdngjAt/sdxbpRTdLxtXi3mUGbCGqF++sqQhFxKJrdtPjygal9QzfIf/U6ss2n
MLlOoJAmXgjXZy+J8ukuHIabcaIXO+xnLfJKY0At0P7r0muMLGa13/0za3z5ibsD
YmH4fBEE44Frxs3IQnoCWtXZV182t120vp+cPoZ8zwe/0yqF+g6+cxnMzD2tO0cR
GNCChIddWzEAs3RjxY0IhdqwCqqkvdaK8cbkeUWdRv9i8djP6EjO2sG6FMe2JRGe
7kwDvUtF4ft0NKCCyKZfWbcPLbBcYkjszeNJB27DKlFBkeIPtEiorTIhTbpg43qy
WqYlxtD4AUAj9KDXn+M95APSnZaHKqvdQNhadYyRcrbS6sbvUiQ3f8NwOTMVrSrY
EzlKMHUjA6wEP+Ht/y4RrrpudM1EZerK1ateRjmsPNU/Ta/3+WRnfZeE0I7EtC+j
lJMjcE3Vg+K0GAFoAXJT+cqKowczJZKm4ECofswx5tiIgj9A9wq9kIULtNW2f5JU
0rQJugno6kNsUNtEd/2zhHPeERCBsgCVJfT1enbDD05lIol4qYdoUz5ZP4ogWpPc
vLUleD2vd1hBC8ziAFhT6UAY62DHcAB+vqtX91gkajMXGMgu24n/CFClWTTdm4Sq
ZDqIvN2ZNh65/S0Z5lRkMP3Ms4ktOx7q776CwPQY37Swn3fyV1/V0zobi1NY6u4i
wySxNXtmXDqUGoNFMoV4sabvUn6Lck3egEnrOWxTHo0y4fO0/1jP4O0WubujTxA4
C+yVdkKPWz9+ua1l1YT5KRPX9bHKXXGn+JZ3O2DOV2RoLYTRz3MwPTljARhupgu9
rKwUOmdNNINBiY344nz6yuJMg31ELT1WIhwF4tfNbREB1BT/HpjOI7p57W+Skw2s
qlCB9Oo3qiAlbL3uukQUyJu6Lp6c/wFsMTuecTdlZD7kreTRVyPEZJeSpUllTIVh
IVIyaDCEwkreXVkWqPB/0HfiZPoJZb3Cux6f7Iq00eImLFYeLIJJzpwHwRhvowLd
0e6uyFD+EPnKYfjUwfJh1h9aEIxrLVbUcpkcEALjnTK0Ar/jP1hfRhG870Wls5SA
/jJ9FLxZBCvuye3HGwaW19ufSoN1Y1rb3Uepqi8mPhuPVDhXKQDdEOKhxopJlIcE
yNR0kCGaPqu3JcpgLgSDsFRKl0BDlKiXLvNLqnBRZWyWzD0zEnewA2zZLcc+9EDO
MAHpeB8DK+LvdT0RfJm+WQKb1bFi2lExvIN8ZagkiOHM8gXfwSV+DSfHDmEMTYQT
bq9iARYiPEJikkdMGlR/uYJ8K6G4WRnt2Ruf60t/5RrRe8AbY26qUjAdGtwi7DwS
y7PZXY9c7rzUB5HvmgAhpAn/QF7wHZsOdJWLTZW4L/PeSuQqnEe4JioQv+IT0Ste
561yRK5ExnPrW4CgUFKBtVBdzZdghaIUO+kzKISgkxawpGOkIlsq2imH/Maq3Wy0
Wni5zlBDQasMm4AV5z2d8ifUr84TxbmzTXHKMM+r6feb/4kXOvYDPUAZevyzoCy0
yC/wL1uRfR8f0lDdFOF8E+u6ZC+QtMeJ6XZQOF2+kik0yvLkStajp3UQHFCA9a9b
/nSPFTR97GANKUnJ9tjWJiHqAgiH6j/A9k58v+6Uf4NtJGKryyBh23rF4oxr2jWX
ZDCIyr+QltbsF7hsVTHjUNcc0/+CYh+sraAPcyB9Ui2+exL9+2KmKcPI3Ax1IRB+
p8iiCwsg5qRSK84UNpkw451ljRKCe4evHduJr6XxneJqwMwUd5IQ19tfWkCEisrC
q4YlUG9PMihY5boPk6ClJc2qRqTu2zq6VA/sYShOGmIJuaLx3BRUrYiplKpUag7e
cs4p6LXwj5UgFLlH4LX19u7halcgNEayZ5N14GzzcUeJ2xrdhwpC0L1upbraq27d
exXIZo5io3G0iLR/3Lvdq7zBYjVgJyZXlZIyBwx+ZJaeUv7doBOyhd3cZ1BryC58
Ne1VydvXEtj7/Rv9PYT3asUISryHXFDRq1HE0LrOBd7U12aGsfychUXr66bV6lXw
LVZQV9PVHP80nnFKMmKzwdUKOfSIEhz08SpRp9TS/rMf5iJ9bc/qWVamHLRFtzst
Uih4mtcX7ECxxWqBog6dq0cQMkqyglYYS3p0WiEAZeMtuex9ItFq71aoA/suAzyy
JuOpJrLR0PXZQL7dA64zTR09yOJn31EKCbULB7rgrvI8sa/Im2luygGPGZ7gzwKH
AKd1rkfL/l5cHJwHfIQ+zJrtg1yzqEByEtSBwz6KEqNKhEiuSzCC0F3/cMxVQsOT
KOWfEq03au15j9pDocJSamilIAsNY6PA+CmV6JM4eKaW2jJ3LLBv1vEyOB6V1zZ8
aD5IUkVKCd2xhXfmIjZZYI91mIiNaAWlM/ZurCzhXY54Fs6L7oGe8qZ4+Ezi8zvD
nFNurJrlUzHjdmAKy07+y52v9N2bYay8KKSM2kbOSE+SHkIkdQ8+hWc4991TuzUk
S25Vma0B+t6MkSUmBhCMHx6rgbNqB4ZqQEkIW9iiy6EN/HUi32GPGOq3cK2uXUxo
9nx/kQATciwvGdha3YVrq2n/S/p2Wvo8Nu3dImJpe0vzCURiZaUApJd5e/ahJCRY
1UUhP1xifiYlsJ6/eh6VkFbeT4Cl+/BkhQY3Lwq9k1RohKzXd34XoUCaXPfV8wfs
WhuV9WH9t7+QYbcpjdcSI5ScLui04Wm2jW7si0g8F2WLTgZL09N7CF6Rv5AMhRPE
CDXr4VXlOAs9SKSYc39pauwjuPplzyzc8L2Bzm9lSlVfKk6Bfg7R2ubGgMZFD4Jc
8HHfUViTtJb4cr0nuUto2OGhZUJ2cY0eyLQNF7ch3ATVVEqUWdw/ef5HF4/QxGkQ
2sZMAzdtLpvNKLS5qInNhUkoR8iVZQFoG8sqWEnArMy2MhpjM0WNC1fnH03mC+9Q
mmC8fNoQegPH/UCI/rWZqJlc1CO0AHtkLer2+hSdd3ecFfa/AFFhB8YPA6T/+xqM
DJRt4yKe6vNaHLYNWupwst2vd3DwqCUq6uUjhSXqOYJJ/wV9mdAw2As2u8S4QfhQ
Ev+A/eQngsRqTWUxiC0YmBo4hA079HTh3HAoaDEqrUiCrT3Ndj9z+/lW/PpjeKjy
qSlANgHK3Ew+pfYjDVSIoPMqkOqH5nDHsr4/nTjKyYPo4dEIteUYxQ9JMnx1WB4u
DguyGG9rbrafNCKRyJIbXOpIqLcmwpLFnAILDxNfoHdogOgVrzM7GqN6QKKeWKiX
rcM1QTYBi35YRV7fcmRm+mjC5xIkx7WMfdFC3nvpss0mADYvntvfYyiwOvc9pvxF
QZTnYaqyWElD/c58lwJLs0HpNRZpA1wLbextA9a5PgRzrfrrQy8bQu2wi1H20pZM
CQYMkZAmcdmEa+0vrhYHHluOmT+iynpGoYMiLJmjONWx2g/4SK+hzWEZGx3GB7DF
rtHThQcakYPgtCrnofaw9cQ1vfeNYUB9lm3kOKkiYQylvlAEktTLvncYQ8lex5ef
aBuGM+ksQA7FzyTXo5Y1UQzxBnQG6IPuKImPI/9KMA3l+yW0z5jgbsrONhW8yHac
C8Ylncv2nmzZbi/COVd1fiXSHO5yYzt9O3A5noBqyvS+DKjEVVphuoKliLzmdULZ
8xeM0PefFM9RtHCByW4eFDvAdboHfp2kRLbxaXJOWp5WZv28mK2APubUlboPH/2u
/rcF4q1vFHXLBszQszE9WEliF/znGX1CAfSZAVIAhXEHYcrdJufV8Vug27EETFD9
nEhkn2izV1lYOzdDyH5w3vITo0srgfJchI3tHDBUr7mLdnjyKzOe1B8taINZE7Mh
Wf2ZxGSgt4c+75XBeZsZGvCTH4SppUDc0D3QJ7TfoSUTEpt04uYCFDsnMn6DCajP
+/WmmUb7Me7Sq8D4S7BiC3EW1BTJ94/Pt6K5rCU8ChLLsNAd2UxA8QE3lnyO6ClU
lcCCco8MyEBdYxG2eTT22re0RDJwdWuLy95iJxzyp/Nx8fCphBatoNH9AX/yURoW
uazBP7sShCRIfMKs0Iif+pXzbsyqsg7pyBDxzvzH4ILU1qNS+QvLf929zqIvjk/e
D33/oUVHI7mTlxfosjcIlNnxXEVpDAgxHmvH/UYfde0LkeymawsEg37zDamuFdv9
PgVyk2uXE85OFTMI91SuNHXlMQpUn/fUCVy1gQibf6LTWzjgMG6AUoZv+tJRU34X
Djurdgrnt02giHqEBQfny0t8d+Qbcp6WygsyLcJfMLPndOa9Wc+Q9kDTSMCR/+4G
nodzqsn9iI+otA9fRylKoPir7LYUQ3tnLYtBbdBT9KlJvQeRhldqhiekmU+IK+W/
N22IXGHoFonfTc01Ft3FuGN1sFPjqhWUhNVtkyiaGRIL7GLbqYDKlRV/i9oYLtC+
qqEon4bAWu/4GpBvLHZ54P80TZXkednOj7LVxMHvQLAU3yFyuIK6mcfcPQZTv1Vu
3NL8kINZk9TfvJkF9aNW3OsMyFmf0Zi7cp2gLZc/2llJ8O2LVKPccEcBAvHuB0GD
sDLOPr+k5KEKs6rbNu0o245irLNJa5M22pZh7lTsE/UE0oB8H/EqvGqkECgvqcyE
2CQ9Np1RMqjvEtbVx/gNDWvlF60F2J8iNSYHpjjKOwIfsLJh0QqU4DAcKp3X/SIX
vEy+tAfFKy20Pdr0b1agnbPe6NH7aWllWxlBM79zlZEkZ6QGQhRts7bvpDynbexU
CbUmZPhAUC/vDBS/HR1a+go3+VB9INywSQYISEC4bhQj0kS3UAmjswCAS3QR479J
CEtP3BlqnZoq+2u7fPNHb2qR1Y1flqG6UQFjCF2fmjTTD6hyZadi206bTicKD3O4
Nh4nvoPULGwFxb0XTOFj/jxFLHRoKySxoyxs5Phx78/gAwu5n0mWMK+jSwiIfci9
KviL9eicA8dXcCNqW46FgqQINmI5fl+BJ6vjGxcmctxMYHPq3QPgrQGTimQ/Tq2N
IJNhdMdWAMa3/OakMPl9JDTxUvU+vwjfh1HIDhAW3vbwGEeoX6nUFFPm6LHuhG7+
UpTPIJ1B+mfzuPJiHQV21qckJX/u65tljXMiMk9EoM3aILwCMBcVL5h+G+B66d/p
okhkenUKyM2v/+cBwFX+XwTd4jyQp0A2AouPTE/Zj6OnH0issrQPgSQqhAZuWSJk
LNT61Apul84bFVg6jcj5mRpkThsojhtR4ARll5ZwvZb5SWMY3Ij4XqG9AGKV6VAQ
p8wpyVc6TRZdpwauzjPTb5/2MrgvEkjvP13sJbqoRszp1AMuiTO9CBgx9wX+0cQ2
AAy3AXeaJDerXahYFjKc8jSBuHgtbYIHZ54gAILDMCKVo38knb5liH0SIVi9Kqye
KS2XPn2yNVnM+Wo+p0wALBC6lo0A4FCBju/HXOcldsGOCuPhfn9vTFW+TgVkMn4G
ufxjHFzO3VPL4Trl4+N5LVnUkVj6ryouT4ZnjTsgvsYlql1kWPCRjh/6L/9wWbC8
5lYji1lv6p1gglOt94LX/gNHB+KmQE3MXxENPaM0ZO4fkJlZUxy726BKTU1cxP/b
JofQ2oyZHghEeYAodU9Z+hNz+7f9gSxqbxa5V9DfnH+53I5i/0ft4jiDt4wsAaEz
FaXjsAyxnotfhM8MIICy/d3ED10V2eBWWzkOlBmy1EspcNBcH6/kYz6baMpNEC/j
uWrCCBoo3Kt/Po1OFJ9ez7c3EDw9oG2clR3KKZ9ISQf4dB8oSj5dImkcjqBOWlLg
kmezATtnPcA0YrqUp8eyug9++vmJb/rhI78mi1v6lWrOYQ9i9ppP92iJNX9XVRXy
PSNosXpAb7NmOyHVuJwnO71YP7bmvzUnXiFhNBFZTOH1O0aXUvLWuGkFNaiyMOiu
REFbI98OHCDn48MD9I3gu+hRKL2M9MLWYcJNsmquyzUjZz7iSpCojkYNMBO0lOVi
mV1Uizt+E6w1Q2LXHUmDvjpcdhD7BtdBWUZ1mV53vvBNRcmExT5lJXAvN2iNj2Lt
vKg6fVCnYHqY+PooWzaNgI5YoziD5j6E4bEGVvJQgXMwhJ0iCwKOjdopbT+8L7zO
Awy8kTNPcrCvnjEdheyHr0LRGdwIVrKqMCiRNP2jvcliRl76uI+O13iLUlBsZv6i
S+5Cp8ehAvBpRCA+nOIlpRN+1LuzPFK4kDunD3mPxhJjxZ7yv+c5MOZWU9HFQiyH
kmNtZgiJWi/X9iWf4DVE/T+BX9iUsJEyqZ7Rrg0dsOZUwG6T9QG+B2tfGC+WrPaz
ctYvNcHseuXF0IizA566rJyJi74bpI56xHYs7mo35YFxPkE0WF0zsFfFO3XR2eRn
d+UhVafQcT1wZdzv+o2sQ+j7qxTKWEh9xwnC5UIal8i9hx8pzwf2pFACZ6e3NVcO
S3HgOdC/Zk3jOrgvV3bNUKniuagwrZWwJloW8gPPkib04lmKLoBH7Gm/eHiFKfPE
umlS1NHOHYkNgWWcNnx52VXBQ1rfS2ouV/AxakUrQCw8ZvFp+AmQ5QY4g0A7JeAq
AzKNt9qqzPDRJgSt/JkDe4g8Is/k1hw42JxE0SBgByFCJrMoBduAaJL6CHnsQYCN
L2UBg5vYBV3z1dK+Cw4rqx4D1ogW24g9NYOkkQMibgtQXGvG38I+EBz69WB4udl5
Xr6JrKMq1+pJOkQrQaCMBWQ0gzzZII1v2RUWt7C4m3X+3SolHipjit3rIFzxpWBI
k86wSlHJt1wdPztgUnIXPKirc/rdz4hQ2ha9/WShANJilqiJBuEGOkh564LtXc1h
i3LjeqtdnScJz2CKndc04P8I//w+Li9uc4DvOdGtJ/sT/u7OnWXSBWhUhOjuUTMX
xElCWz8wVThvXqOAvcHqHKuC+pkT9r7EiD7fyj0sQNJTF1MFyPCfUALhCWvprAzR
vuOP/0sujL5BG2nelYKdjro5q/n6ZMJTs7uAJ7wrz2/AJZL9/iU7Zs2ajf22ydKK
/HPmtWWT2724WyMcNBObqGT6okEAI94MO0xJwTo2c1jWSpkjLvw6deYcCWQclAyL
3NmDxfaZ7q+doXVkI5xuP6j5P/McmbJzxxLWujpHQK7Vc4o1Td6EBPWdT0gX8vJN
ikkDPJiiD8hyq5nRYKg5cr7Yvw09ThjHz/uzhkHpA8IFViX9KATOfUJaiCvSQZ1N
dXC607ddXJw1RNTFT18Ed5UXUV2L4GEPgunbTX8GYN9nadPZsrSMEQohQZAqbkh9
tFl/nk095VQ2HtPJF7Yp/xqgP8qCXmKZA/bctyK/p/UfPeP8pJCx3tfvBepLQ4Vz
PjMi2iwo2r10/B6Q+TfHpqGgDyjrpzSYzM9TcXDRVW0zqpZ4PRzUSfLtSsh3ZJZh
pRl98NeTjkFjezi8EVTIh1fmDHn0PYUIaolAGc8df+chtFQvrh/NAWeWL9V/RKyM
Ij+2pMdvnaG0wseQAuLLnYsmU991/Wr6TiU1YLVp2bhWhmy9IMGqcgz5tJMd19NB
sa6/8HHuB63Pyoo9iEYqtGYwaUkeFezpdeEKgo4nrPwVklI6g32Zuxj7NunmXfS+
EqFEhf/v8UqqYt7MjDTniSgl7gtGUb4X4yspvl3M/PAcJu117lfD29n8mUrsOjo6
grm5YbVddSmgbvFSVpn4tlaU5MuP4R3HdgBuZku3oeNtnFUWwUUCOe3jJwbyevyH
Qhx1EFUIF0MXdE0dYfcBCnNd4DUD+dkPfstDTZW9GN7xQ/5AVWDjZKB16nLBvDMy
hw+9RJX++IqVgSW5z9weJ2pgWm0vHOKdQIOry7EcOIil25Y+W+RKis1M2RHaBtlX
Evipo9rdsPji8Cncua7TviNaK0C7MXRs1nOr6s/l+/H9c8x5EaU2oMm4azsh4Sel
5L6577bNfL78Kn5clAqalQRgwcbowRPGKuEdu1fgYCYPJYMxKxV/En20eX8SJFmc
5phzldSBrtU7fhfN8gFZB+SAAbI/++0ne0jxN24ee1ebFxDXkXCwCkRSWanqZRg1
3UMuKPqyx9g5TRa5/LTRIJHWB3fggUFjSVXGhG4dk9p+/K9+u/qVHGbE4IdqMv7S
ilwlBN2R24DCH65ah+i6fobS//fC3goF0vDy734s3T8A7NTb3dFRPH9ImBXfWcPh
KcRHhCsDhuVBkayT5TCalhKgTbETOleCGk64O5m7Serwz4UpunLQXizgmlN/ozBZ
PXDx0ykAlBewdsPlBKofAkh+uGepwnFU5ChpZ7ozQqb66/PbNBhRQ2NkBAtr1dE6
3jJXt5mjyeKoQm3iCXep4yhLOne9INWHd1Z8OaweuScf7z/r7ow9GMzrqrHbclWZ
TxQ3krTaXjeHu/gJylfUKN3kU57620a4iC5Wg6+gdjFoqkWKM/7b9MghTc2rmObH
4rd3EqNMtltDOnQXRwdRqfChXaA4tZl3u0Q3vwc5t52VVeRg+Nci8NQ/cO18vD/J
i6D5PGC9QtUpxfD6XtliPkA7ExvPupDUhtHZslq4lSG5RJMUiD62O4Sw1N626d/c
qibAopOSM0+++6xERU9kz1ZB6kcxA5DPl74PciOXkkI/qNZGTYVPn56YPHO7U6QN
QzXEXA6rV8CZsvqrRpaugxylewb9vdIT7Og05MZQ9mqtKBlKvt5jsbfQyKfQSsHG
eqYXnI6/Jtg6audKT9tv1nFlF4LyJ/BIQqPHcWd68O6RSFP+wdIneQuNQUcEsi56
8PG9IM40nGDB1WQgHLM6FrR+zv5TMoRF642jPjkauIDMfLHdaTgIjXHjnn0D84lR
KUa79uzbpz79CFwfqLal2zT1y1VgjW0wsBwRlhMM5mYXlTkSAH3kTKtTsz8WXIX9
b7hZf+Na9X2TkqW1uK4UTg==
`protect END_PROTECTED
