`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F5xImYlZXQiA0OT0ElBixs2mubLUCur/qEubQIcKzY+98pIn2wzx6TXFKRcNcsEA
g2WD5zStvKmxXp7W8T+M6EAOhDj91ALgbKJiC+YZpbXC1Wl4wA5iD/MX1C351mtu
/9WI2YzOZrZqnjz7p76sTyFDdqI0lSKCiUHg/38Jpj/1+Amrwkva7H1gTq0oEL0/
b/RzKSxbTwKd2smSM4E3aWA0XUjVSvsI8Rxl9jKW3SqwtOklqrbopVqBhMmnENSu
3axXIL4hw+uLMstl1YY5rdqvoGDNEoA3BJMZvI91RjwOxyXY5nKiHar7MsLjqCKU
y40/4ZuMcIDxRtw/2d/SpiEOgl0R5103mSCKqyvjipZSbRLDWSyB4nw+buRTdW+c
ep70+vTD2EtwrkeKB+AEHulCaSBRV1H20olvLrjhFt7nusuUxQqa88ZNn7sX1qMS
JVbFStccEqDgiGhIBP44SiA1r35WHgnvr5sV7KzD6YvaEf9sBp/05PzAT97bcHth
TsTzrclfa2vf01/iAx8s8nrSqu/3j8d/ChYdM+hkL7mN/U8sM9mhKdd2I0uAOV1g
NaosGE3nXsLYVxhennuVP59lyBmD268brz4noZjEcUGBdUVcaMPImDnx+ICvtYrK
N/oefZLNc906Kr6c1CXX4ewzvCqrwslH5J7J7d5QeMXZVUMuYX7C6VkynkDwMb+Q
Od5Ov+eVPRmg2hI7qk/kZBuR5reJPIP9cIAfxTLz6Q5BemnMH4XVGzdaA3UqsZFK
EyZ7cykmhlF1f4E14AE/Ga4pE/RjlU19EYTurk4MztXU+bGdMhbXHOhUPaYThvbi
fESx9UZNF+LbDvVaQi78373DwcDUY74AbEctjVSHULGmhRdZPaxPTrvQjbxv9Ydj
BOLnHXXS8EedMuj0TwVHVc7e/IT/GSoBoAtPTRubda3sqr1grvWv2Rx4G5c1aVQJ
mpTFM8RdjqKQTWPwfzgpR4Ml2iPWWH2k8n7JLmoSDCRxpleMQruozo5yNfOU3utM
mMN8jWK7CzY20Bq+3SMCelaJMFVQsWFy/t4m6QmBoqkw5O/HrDG8CDV2PlDzMe5Q
Z9v1IgvcpDkb6xZYUzBcvYL4xHYE8qrgh2RruSQ4UYPJlgoZDOVKun03UHZuEF3V
xbhbOYCVo5AwB/C3ixj6VQG/DiVd4rtviHJJ52Xe25LXS8NqmW9vi/uVu/FXKtwQ
+SnU6cCoP1G0f+o4qsbnEpfTW1DF8IU3Z2o8O64XQhRRD+HDQylgy6wJBoU2ZdAc
O5vwIj8a9uWqbS4pQbEI84tnnenbGHRlKGPkC7dIpEXMeBR2fhhAFq3I5VLQ6RdB
57kQiy1/adAwpTSFQvDFu9Sqn9GlegeU6ekOMZlRHu7u3NUUVbYJMBk+krkseUhB
LppnasXVvToMiSGz/v9PBCmL35tx3NXja7oIHqOI70SuK7PNxNsIBskMzT85/Pfv
sHtw8cqtxhCQgqOxcxnjHlOtkKXDT7rGte7Y741mW6KQzaZrle+GPiC57SzQJRO1
QOw7ndm+/Wsu8bq7mJVHQeEEoR2IVkDQGQPYfcy6NcLGAqsotr9MsV+WwaQTvVqB
4Ri1FDAd++fMiHngLKX8WMKv6YfHmSzKuZgh6EWc6wnCtst9tXQwwxPXk4Q/K+3n
4xUmtr0f3eXAF+BVJOpsSRmFuqa/IXWZlVYXOx+GzdWNX21DGvc2tiEyC2XKD88v
Ggi3L+mGBi0MQmHZlERgPA7fLThtV86JxT350hgIreSMsuw/3vOfmjlErzXjqgny
ngmJjfKAliBtE2OeHFG6MuJ6HK8QCdTRHV//YAIRlHSCZ3TX+U84TuuNxu7jVJOY
xPM9a7wAmmqn7+7Qcg5ayZVWmj01R5ynJlaP+uJfzbjS3rG7AEmOxZrorHumXLmE
pGOPXj8VOIYhpKPMm9Z3zFxNlZCb4nqgCxuiai0lGK0WB/U0zoLQdT4wU7BeLPyh
S/MyRExTswRish5S1sM12HEUB86ApSTsdUOi9+PA27xpHTqj7rukLkendGaYahR8
e4i8J5j7qzf5oL06UrfHgmY2auPxIev59bkIyE6MP5GGbrtEKlYBcy+ESh1s5eV3
IZuIkfCLrYPBozjvnKO8xNYEWUYqmMZrK1tVRrEPshRHC9JqnvUJKSB0q5NgDmFk
/baTSyFa7MHFtcn74l98yh4OVvGkgDibQ0JX4yBCWGWYSkG9+f6LtDnlWd64tZIA
YYyR0igOKTRiThhKuko8SLDJYW/ZE4DncutrpffTRLx0m0z1McfDKnAq9v9c4aFz
fv545SHivadL11UJzoiY8Gouk9fxyhMo78S81BevbIpyQqjkRIC1wGzRxk5CGYqi
vUzTmWmGDLu9V75RzEnCU7WLNz9z5idQu69D0PKq8EtjwV9hv1CO5PBZwbmxSbnH
DO3wYdz3QQpD+hd6h87H4pMedg4/Eq1vVAQI7rbHyGi/ONz02XJ/uNUtPZXxAlfW
k5agdJy6+D7cfxllldkURyb0Ra2sBRBny8ynARuof8zqBn+d3SeF3f2JDBIb411m
rpLeNiUueAlLiTGDEoif3X0e64cRpaQUa/pnckzlFcfBmoG//ZyLlQ5Gqb4s7wgb
n3RwzvQJis68pS3kuVkAphJ0P12xqphzu8pPUiMgppe0l6oKoK8zwLNr5mGR0lT4
FvbhEspitB8HNWcSm8NOH81N5yajyHKH21cgBzKb6vC8R0WIRnrIVC2NIR66s84K
5ztsSECMyrYX6nHmlb14wYiSCbcJ8AGXIlrKdkXI4O2RkzxoIxmkgDEKOE09BAzj
gdgVnnUnwKj4F47qjePEIAJPts+BSfbPociK3rzZcGuHGSG65fFtCAa00C1nQLhP
O2/1HU/7qY5oR7hOdEsxBEVE0LS964h47Cpbe4ixsGgCQYzh+F+qrlH3vyxa9Mrx
I8QXNt734ZSq5FMXRIJfpCYf6mDNGKOnVIZGJlA//MbW/S8bwYsN1nVS+vLGXO5s
6m0jwH24RcLIU3ULl1UKFra6F3NhPTtJiasiJGxHuL3UQG+z1z8n+JBZnE8LQv+2
tIG0Krix1AKINWCYubq3KeW3QlNRGHdx+mIGNknhu4fqRJcQwgbVC5NHwPCxnOW9
vnnmEp6LxNEAa2S6x62bPU+npa8smae4EkJmTKpX7688dZ/8TQRc3d13ZeGYshh0
mQzmAMzI2VbUPyiwFnwbISBC12JYVx7YiAyBFjASR7HCczxn9MgYkA9UPT24twvF
bpSnWrIkvXJoJZXDbUMaecqm6Null/fuOP891Yhy+3NmqtsZgxP6xuplZREsu/0p
7tENZRWDYePQtymqFI5IimqdAQ6NnlDsfImSKC0XsofAWjDVTcirAFF/vQPOTAJ/
FivcpdxrJeGU1Gj9A/a2O0eQvYIH3iE0m+OnygVkbTeaOg85bBS3USmJ+6yyrcLn
s/LMiILwXGKFHGUXpjWz5qdx7QbH/0DNFiGmOpNwnC1eGN1a8nWrDM5WsU89FNBP
9fqFJtm3Qw0duegND1FGfPiGVv/0rbeDrYnQ/QS+OqHXsh1KiWtakTst5F9kmRNw
kzSt+k0jWCRK9QOX24o/lap9BKl/z9UPHXCMAFCPv9V393KQWTpdIKEqwMJGEuz8
GdVZWdawPrXXUn//hP8gXhAz48hbjlptECJuYOI4g9I=
`protect END_PROTECTED
