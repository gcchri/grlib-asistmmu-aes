`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kksiP1y7v1WY+/VZv+aeCGQ0uI58SjD4uEFwCThzjw01YWp7wezAlOQSvSa5Rp8g
tatj7nawBiyLXHRqiDP8JK4qY6YMzZ1/SSDmy9Xm1kpVqbu8ejY/gVkkkLZW1XK8
WZ/kycf+vh7hDSkPcYh/aZ3V6r9cPHfn+ZVp+pAS6ryiTwLDK2rOHVQCUoFQsN+I
bdmC/g/7m/iFFOP8PQWz4oaF8ltAfUoH38C5V6Z1qTfC9zmIl52sVQnCpVbEm+4M
u/tX21sXb4xy+Wq/EFQ/X+/yf7dTU/HHFAW8h97aJJ59NDwRQzY5bVzl2jhhuTAc
sviQmHzKEPSubxe3aNrHAOay+A7SWwcOG0VqntwVh8hjArdlf76imYMYL/BWiZAo
RxIzA9qtCQiLSC1eQB63MGYTQHGvDF2r0VsctRvrusELPTkzpgJULu1OcoSZAEHf
0fWK06FD6djNIXqC+qChrrHWcHZAxCsiK4Mpu02tGgK7QJzAite9aLNwK83ZhEsj
eyK/7Pk+tyzEMt4vXhMt2hgFN3CVTEGfP/Y2I4rpJs/D6S22Mh0nWlPSlwUbKkTG
OLW7lhycKnxWqBUHMbQWNQ==
`protect END_PROTECTED
