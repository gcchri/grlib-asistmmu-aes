`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TlAywi90/ah9pmooJ8bmwQYRurIttjum+SS0m3v6aPqNMm4TmUIU8+klZ99pjQeG
lhSk+UndRLANk2zMHHXb1aMk950zX3Wddjr6gWwuWnnzgXFaL1RbwvCHS70MSWNO
aWF/xKYcLo/MUtmxzCey5tg9KKP6+QZvtg5VygDgCXkEH/w9Jt3jTQmTW1xChegg
/3Cq+Aow8Wa3zaRIEs7VmuVG7xkFLxYismLGn0YOvr/DztIydjrbtMQQho0G1TIx
DjKkKqwZavBB124nNLG3KwxUspp0yTTj6MS2MGZECsGykpHKY9TOSusw3AR6qeyq
dJgmXRrSCzlIp184spmgdThNeT8VWACJ8HXizdYOepwgLvzB7iQ3JAWfqxeNRipN
uUsVAHdG84633U25pgWKyk79Cq8a3fT1eSPluCFtHEK06oKeBxBFuUjJM8AnLd4+
Cru2fl/Vb/CggpwwqBvZHjF/YtgmiXfAGEiI02FdOfhGFIMztQy0B7uwZ6G1Pjy6
DOsXJ1nmXCTg7vylW7EDxyGxNJpOYCQP+pIemeiCgN2zxhfV5ZrIO4A48G25JtqY
VdDwa0Qp8BdSiX/AfjYqonO6KV8NgiJB2KBlEv3qEtX8sWL3f6xP14TOuRUkimbn
kxucd/cJv3wRojdvvhN/4w==
`protect END_PROTECTED
