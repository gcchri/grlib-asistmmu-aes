`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVZBCiueRBTPki74YcLNCFKp1Kpg9X6uSwrz6pkgIv2nJ4Rm8UOLT3sBt8ygO84h
CyXOv6OVTXMPXYeemO2v2Eft4gC3unx1lqjkJpJWwjrGOTRUGGqdY212egF2EzTa
44vhsk7jp49gwLAMU324Y4yJmrpZV3XI3Zt0SWYCnXkszleLudnsBI7ArZUbn9Kn
tYJFx3xotCVUsBuUM7rJxhkKrTPSIFNgv9Z2IrPjJ/1biaktXNis7lsiyf+oGzX+
Uu+lcsyBfv94m0h9OUVhW+VeKlPFha19E/5mSEFoJXaWRK3fdwRsdjSt9IWrW5ty
CqvNf+CC37rcDQExRLzFHpeV8ikooy6sVFrJ5062OZjR/9Y8dA7I9rnZ8KQEO5bG
Cmtx0lXEbWLLaMUA2JwVJr5rvuKOgNQLnpoKQld+o8q7cPv9Cdo8YyKmDuJmrPPQ
+L/CFkGJ6WcjTIbowTIsLOdXgkIkpfxDw1rfw3oCQnDlexpUUsRC6ZatV/j3BYa3
TlIGIfuhvJdkXi2QW7rEnGvbp5qq3W9G2T9RmotrUv3f2YibcT7sHCIjtmL5/Vy0
39HqdneHud+NhZxQ75JOjp5NFmFvS84u3I6XKXpWQ6HIJEvI6eAmX6ufT9N7I793
`protect END_PROTECTED
