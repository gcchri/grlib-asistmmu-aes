`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kCpxpRnMIFjpy5kVfJEZQMIiG6zXf4ipGdM561xCjPpXQRv8HDaY7QEocfCdj/GS
veLYagrHVZKCyb8+TY/LpT8FD9sBcNJn9zNbl9IWoyjhqGrXJetuVfsnVjUm0fUT
3X3gA4L6Idup7n/FC7MA2q47/4B+iQuwYDeceFrLHTSxe5CL6dBGmpzG3NvgZOgz
q3NTlKFYH4gjo8kNPXFkxT8sZvmtL/TeXi4LtTYakr/JWkIiqriMZrKb/eAxu/Rt
S9/2QuYT5SlUFAwsyW8tf1z2lmxDakoql9AQb0w3eYVo6EOwlzT81hHGMhdUxfno
PokcSI3c3jGlDtQXoHQdEqIb+Zl0591M3p0EV+ped+PSgcgTr9j41twfSf9LpNLp
Wju5WCfE3bGAuLoEDEToQm/QZIW5aUWrI8y/qL1uQLJIjDT351JE505VURls/fyB
hRYRXzW+qmEvBWyCobbkLOXGKHZmy3mvwRQBZ7IMNmM=
`protect END_PROTECTED
