`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9l9EbZU912Ctfj8ZSjmbUCHRr/dqf0J12s+1tzpERbr22V1wxfZdmAxpW5sepnu
6H9r+ZqpLpO05EIAiOmjuCPXWfAs+2losgHA7D9XmY311s0tPegKLf6d11UB1qFB
vQmx7CQjC66nVvM+tq8gn+F+FdFDV9+Mp709roXh+pdIJ/VwhEF3jcH2LlXxRUiz
NuxSuwn/Gle7lO+IWay0ozAY5tNiUUiL4ClvZ+9JoNgYMIMSLcwxItai+ilQVVzJ
QK4DtfdtH2Iu8CyMh65V9YhIgL9uurfdmm4O0s+/8VUWruu/umT/fkfkMQI/v09G
92QIiTbBLIJh3R44Hbju09Qrhuizo4sDbecH+maQtNY0JOPoFFiGpIqz58z5k3Uj
`protect END_PROTECTED
