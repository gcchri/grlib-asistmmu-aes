`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OM3mPiAvcuDCp8eV5gaRKT/11BeIJ9p5teX19CKJXbsVffipQSlKrKPwxVTj+qkd
iqQblTH/7D4ao0MQ0+7gvhhmHf4B3DnZxEoy13/wEO4sdEwL3U5fcZCbvQJ8Na4u
5htIF8Drtc+20/cfFoxVhkvMWK0KGbZt1cF53Skx1vcpeg//pudDE4dIElN79oix
YDsHaEqOI1AzP4i2feEnTuZC/tXvXsDCNmmclHNXIArwFto9FWet6l/U8uQqHeG7
308ljtXX8XMzfCFzHRjm9VdZCjXawzfSZQsX/x/0blM/eANtHY/3xuCOK45P1n4z
VmO+bmuiHDlvdi/VxWSI3R0fTqAYbPA6fyLnR0FmHFwJhbsP7g3Y822t4j+oSgFC
fJq9/u7SN/4soT1vrSQn37IDmIzc0VtWdACMe/Bx9PVAQsPg2aFxDTrFRcBqeuCn
CDKXrLuZ89R6Tr1YR1OiARQqHpCghgov7pIXOv65zyxdRdQIprwos3Hfh9yNHnfi
OgRMdAZfz7vtKiHw/FWqv4+9motAEas+f6qjyw8WlSbWX3w6YGJ7+a1cGQKkd4Ze
ftmd/TYWBXOj7g5eHoILr+Ylyn1yB/6ned+1MM5cthvkIXkn1k+4/u0g0RB0PG7P
+YbPNpX6DgusGS4nEupcDvm1cC/AbQ2bHqh1Cvy+wecqiwxAkiWlPeOa+uaBiH1S
psBE4be1eN9p3471M5kguP0SoIA43kJn/lMgLBXlLzjh//SPU4pF7e2LOog1XAxA
M7koZA0sdSq+MgB69gHrEzRNc5BteJwqFe8gbEvZK2bB4tX6iYwzEz+CYCk94IhM
ZU9kaD250Jq7RRw4ga/fYFgkNWPj0BkFBCX+Qyh+k5yEw44tNt/0d3muV9w53qTm
Tz+dV/1QuuUxBOWxOrbUMrtpx5Jhyxt54/kIaaYLdIT1SN+2PCE58G5u7wNrjO36
oylYtu5MYjS1J5pEMVKU4w5siOnreC6EbrUA83nkxDUQbUmLD2A1ZVG92TCurKbF
fikkZuvcYQHICAlVYb5C+t9vSTmmNh7nI9YGWOf/Qiift7KteZPjv9BoaL+sRiLf
n9W/hSejdVag2slbALbndhoOUcG0Med1m3oYZZQenWYBssh0F2s8TMwW1iQ6Zdes
8t/xPZ3NnULo3wnDtbWnaLsW2pfM8ldZ+az3ZmYeW9eMd0+tMSa+pFgrwAL3Y/U5
uo9k58clbHAiXvbyx4xLf15u+7B/rnl1P5BO0qccvv8X854tjXVK4Sl47Dj8p0kM
9xtc1FaQAJ6G/BwGllsQb7dL0/vUBYkoW1NjuqklIgZ+ibAnojnDfGB4V+LD3QZu
+3emi9nE0WtYLvIJy+/IuiuVzmdjL9NY0V6Ko1Cqh0bqD6E1cEFMNJqIzkcrr8PU
mdB4otSZbCnZwzaY+cBwkjcSnJjSPihZdldcBz8EmkuqtvqvWxVRp1VMmW9rLtoV
agQBEHZviKibeTqHJaEGngDl70nO6uzUuIru8dEuoC/yXwoulCcFx/Wmn5mDBRDd
W+vGlUP+hY0tEU4bVSKb/pf9ZRYXpoKoLbsn7zWCZShTSVcEj23AJERd0QK+bQp4
J/DOLgdVfCpsTrUBH47YbQzpK9tFBuQeBOb3AGLXCDkS23s4QG0nfQXIRCy3l+WS
M3FnANwSYFrO8usg/xyNKFQ4nJb5/wLWgTmnrG9wbX5n9OXfIhhVLjqeW2Xyzd6u
UnTwPgIVuDiK8rUwTGIklhqKtnxeJ+xN86Gcn8us8diAqcUCVErRymCwKXBdSsgB
YGc1+hgNvg8LqFrcbH8z4BkLvbgmMMp2dNDy6x8H1OanopBC2oyw1473VbHcD1Ci
6P4RAwa+zvrjWAxqRswk6+I7A+fAbAOdjCLU0DsTfRSVVSN/PJaYsEtKD+DrzTrm
HwwMKPYhZx1GaMib6X8wGtuMghiu1mILTL4JimRyNu0fPp4u1zWQIxNiRckY4pFr
FMKpuMkPsV3OeRzEwzExUrL/3kTDSU4iMOhyorAzuixQ9OnZsekdVdgFm5JPTjP7
gZ7H8+TYC4f4JPDZ8c6ZkWOey4ooOB62J7wSIl1mxOkhUD419U7eoqhyZ1/PrgnC
OamFskAQnPKUdpKsO3ke20zOI+WDc9Irmxq9Kzbu8u5BDFXTuAeomgmVSfFKyUJ+
uuGqjqNM0rtV12Sq7hz75tOUi+ewp4KSoWyGMjvCWEGpxPspKN3FpmHRJjZEjUkg
rA4EtQaTXsl+syx8lHy7F943ueILo5HFlD09CFrgJ+VdS0FG03TGzQEnlE+6TsA6
bid7VgJuvZKCDaY9QxSfC2ZlI7tYAbgROXAYlaBLRje2HbL6DmuDLaiuQOuj/1qG
LYYC72J1smr6bYyRCi8w07I+KQWCp2r3pE7g7XXaDcPNYYQl7p7z9GavtEGPlfpw
aMG1zvU82cCOHAlMAI/3BxIkoUBlA+GlgNgZh2H3sGq+5aD8L6eSx8niTwwZ9/LP
aiZJjwVws2VQ43ERzFlt99/mKtget5BC9rmT0ucsW0e8tWfcDBienHyra/nYFgET
U6WD8qYJHsMRiEJBW7bEhHO7bgQrRqhG/6gfyr23nc+Rhi62fa9PYCiSeBeLblim
jTiethHR5558G1bUflzTV/1stYCWtWsHi+2/506JocKQvp9Ys4AH2D6AVGoRCl/D
br9F1mmS5SEpZu2sTWrxK6m5PauKKhCCwZ3kbCsOlKXFIrdY9uttXwRGOnHBVHtF
5NC76oSHiU6cOQM06LzdriUlIWA6O7swLSdBXMMpKB61rdef/lL8vA0DMF4wY8hl
EZ5Ja/fqbwnHgFI74yqJFiLpOf7ynGE3W//8egag9qS7isEvGLjLZPONnfO76J8Z
6FpzxRfBeRdp0b5JrogCcNU8+oy53fw1G4lg6+pp5eTY0yj0oE666dD8bVzjHzU/
TpE84hIP0aHhma9RgEhKkBEWptWOhLj7SL73NhV0ts73R6stusmu4xbm64p/sQiM
oJBlWW57bdP3qzOz1qh8eHwhkA+Xf9jmAk7Gt0d8t23U3yitbAx1l82mMFSs9hpK
o/7+XvG32L2jCVdHWbUsYLYOb4JCSRH946w0HfwpZm7c0BXXWQ1p+GlpdWp06G6z
sdC8plKQHRS3AjWMutJNQmvvN0qBgHh7pkFYsVKqpY/eJhsP1QdJNKm1OvdoBCYN
RspNmTvILwmBB+JJ6MHTRhA7ldcddDUepOZxguUWnm/ML+T85AZCZz/Uy4nQeINM
v10uz+wvmTNDGJ12gDFcwAvKxWzozPvO8hAVA50Dtc1Q1JoNwwbGxuXbsh7xvbGY
jhZXGs460xH2KQi8uVQXeO6v23xzY1s0Vd1KaJsGcjYhjBPqUPhGdmNTCyRwJmXB
arHV7A+WhQ+TlX4iu4TWhauDADef32JQlFHFckJK84GiF+y94N1uzyax+Hk2YPsU
TtkrP7MEQzDEoG+Ijfqr580bdS0w1mBusCrOvxKZoJcLGWJxBiT2twxrE2hKXwTD
DmDnYt580EPGAaqM+F0JW7bANsbEdw93kcGrl03luQ+0YCW66X/YosMbM5CjcL2v
vZC/R/UiBWGBkU2X/FmWGz7ARYu4DcH491sux44S5aBJQ+3oCfsmIMw6F85KqwqJ
ifs0E8nqsRxsHioibfhUw52TUdLxQSAqsXOdaqFl9SVMBbJs3ucCscWNiOrsqzUT
jKdy3U7lC/Gnw5LSW+knj6q0wgSpuSv6XxPAHoIdw7ANL+Ddjt1oaCJu9kR7+qX/
979sZolR60Kpp/N/TsTyUABECxbFj6Y2S+kXvIAaBeLknj5m0NG7dZF5h2wSn5rj
pS4zyfyj9cvXsUGN6DDbwQxlgbnCR3THomax5bAd8wLDAswxk86cFpxPX+RHIQTb
OJ80j2ZpVXux6UjNyZvCCs+zICQI7a+tXHptJyyP1unq93spesnySpr8xPfYxCG7
wD0qkN7uqqiskWtK/ILsOUuaHChPx7pKQNqipdAiSZEJ1eJ+sgZ2Zl3q1BL/6qiT
IS8sfhteu5V0QZ7Gflp36IuRqbdac6kYHGDacaHJb6E3qtGyBwXy+GZU1jdu3N32
NuI/dj9y7JV7T4XCAg8y2bu5f3onyhKqf8B/P6mJhkJtjEdf57ASgaIk0jNx0D/Z
ShU5ib30iZWekWJpNHdwwQpi0HBU0qeFB6DTVmos2voFc64yeu0WQm1Lu9LQkiqD
ci5qyhGJ3LfsopQkgo12CI3IZpBBT85/eGsfcxbxU+ArTr+SvyfDXOnRM35ege52
Llus0zSByXfpurKv+/bwcbG+fPvwuqTxAZavKYKXuaw5ZNAJYhUC9THsYovZAv1/
2NTF7iwI2C3zoy9mKJVgG7Hm54T3nzd2PHldfejRsCsG4lwoLBxFJeuNDNg6LLTF
rMXJpW9xUYIghgRkaB+C8PgnFt88Nhs/+5N3zazgBSI159unRUOmtaZXBK/MtXGp
XavecNGa8GHzl67Q5EulhFhk4T7n0cbjRsUOh8o+F9e29HW8ZUpfnvPxCmb7cXG1
RZMnGd0ax6Ut2l5FWz2pGnpZ7r49oWG/H0XKWTie+yDmS2ICWznEps6KvVVSlj9m
AD5m1plOL8fTg3+Pq5lc/bUZuL/oMs3N9y5BbSXqreX1ZOEq83JUyXJO3zqSJXDa
fla6dwhLH+cqMfAs4Tki7XE/8oOpybEvOBOFfA/YKUVoynNJo6SGUkcwbIRhWv80
xSCAwqYLLvMPC+FwfrFp2bCE65IY6O8upQT/n8ojGsXqc5E3+qfmRujl4a2wZwpB
Ltl1IXn6Xtq0NLHn+IVpEd9EpzyhAmYTXYz/LKwvq5b+WukySRGZZZF8kDTU6Kld
DH9PMInFhkc+VHorZ22VtS+q4/0WHQUX3uSlo5j7QMdyHWD9Y6VbxHGnuszjQvHm
pzgXNVc6sSEpc2z4M70sm59EYAlDfxNfLxUU39bqXWG+24vUxnYstzi5lM61iSqw
dXYzlKmjkmbrQ3KU4FzYjjhEmmXSzhiQKPmleY6R+QqwzZcOVoZGTCzjY/zsIZlw
R7dEZWXpS1/bEm7/Qs5b4gT/Nk8j7ZhAtgu23tPr5lGcjkSjzvGnZFCxUI66QiQ6
f+thLVvCNZAAcaA4Aw4QAaTXKD++gR4Tn7fcJZrSI8lb6RacSYYFeWuWlq5sbswN
K+k3D9aLpDemkl4XYbpqF78hu8Bvtn44H3OTicHXpOlQP73J0C5AWelk6urv5ebr
wA2OYyuahdeg0AfABREsCiyRUJABQkxSKx+PmfLiqZnMeHckIno/zDQxHshQDbCL
NmV6tmNlFCezs+/cnfGp926V9RlyX5iSmymndnv/HAnubuS0RmcJ1LY0CMjC3wey
1lWOl9KLclD9+eFF/cuUvRqqJoVm0te+HLfjOy8rMosc5mVxvMhdGn16GmtW9Hdk
NuZ8ttOjeB3zaJYOXloCPyHojDK1PVF5piZ3C+vDVwYcjFIBMi4183wdSdXx2jtf
ap598SczhO7u6XThQWTyh1+Z0Vyh3eyQrHcV7A1DHsxpCXprBOAtEOhILjTfPjfm
28TNlBR6YrKrKtEOVkgrv6la3fppxiJbsPrb//nOCc/XrGkMdpBSlaBMwBCkB4HW
ZihwN5oz0vuf66FXC5IoqVnlQ3DZxd+qFOgyZUm0K9kmoCw1ryogvzmnoLZemiYe
fS1U9okdmgdL6IEHESL2XbCP/F6iNy1oZGyZUL2+KRDZ9RgTj2NwQzuHSQhRe+rV
kQWYIfJ43Aq2LscQ2wDTHDjrybBYZYxlD9zeumC/5NBaynlpYJvSuNVZi6MxIu6n
Dulr/LL7NO+LXiFtGwcnLwEYRbUuSTj1M8xpfRL8GfPuHGdPj+Gjc20aHQumMo1D
JxNKQzTdo9l8PU3PwXAflxzox/GNq3HO2QhuYbeT+GueAPMFlXNjAvT4aLbN/rBD
Fk7puBXaprn6I1rtQa2QBkdSIBA5xsrAUJfH8ADmK/Olc8jkD/kHTVIq84he4exh
yYfxuNc3Zl9mauDgM2KLC8YeYBNK8eCaWVDzKodp1Z9gnrGfrSqHsUR7uHbmTTVr
WfCWtaW6bNIwDNTPyIBUGoWNoIH1wNixscUJItq2f+M73shxrRsRHAbWEaIF3i7j
DeZ99aAG7Mc10pr9WNTotBrvs61WifcP2s49Rvm5+zTjnfQnN0HDedt+cum8+4V0
JrjSd9Tm/CAYFOkJc7jqBoaB0C4dKjxdl52tf7073d+p9zLO0yq+drtNYC5HVImz
30jhJyQJkJOIFL3kcYrRVXU+2NIoEjYvp9EqfZixN+y2i/7PARD/02SvAc5aTvTy
3cju5AFhO9sYPrkjmtE++yPnDXVNQXQduIot1w6Z2Yz7lMLDyjC8HiUQiSeIpuvI
h/QVVz6+xT/YW55k/hssWxfy7PQUJ1o69JkiE9GE5Ei+lL0K7nPpQ5TupFeWqz2r
LsjRkiirN6BsesIkVeAtrlZeqJjNNb/S0M8VjQvwduXfxPCML5mW1igSF0nNeGmF
1UhqeN/nfcFs3xdgOq9L9uSRFN9JDvnqn8nozhrYdkxRyZiFuf1kkt8zwK+vnvgQ
QwtbxMUe3e0NqHD/wBS7tJerYq19WhpHnP7xQozWz3KmudUnW8N1t2hdeaMZoZ1O
93lPtwpzIYGp3SCVRJzSwj6rzAaXVan45jmz+NtkDnwIgiQZGdzkj+BbFyZnSAJy
KkYf4vA+nVPTJp6xrXNF4bHU9axQ4RHJE2nCE67an03Ky32g57tGoOqzDyJ/tki1
HIFT1BUS41Tcg36QynRWKcdO2cLQOTsso1+4ZuRF+8mrpBMVh5UbqvBtauceSCYE
r151o9cMgupnIPj0Hie07huZfJE4aqz0qKtcdgbPDVPU2XqmQ2Xf/2hKGtr9e0Q5
aP62eqEdsecGX8We4gapxs1n/THjFiRYWu9lwZJTxvF6vDZXF7KDYvr2dmWyvqze
rrsZWAkStZraIFb5zHfOQnX0r4eK8kVqpUbj4WRxXcArKths1yI/DNGV+4YyybSS
eX5raCOLYuV3NJZZE3Bds5nuooXYRXJeh6PShWEXfjzyIhVZYZQPcGLVwl0AtqBF
tBoCnUmDyzC9HTKa1W3/EURG8qXyVMem+G9z6dXX6GAH8bYr2U8D7kpyqlWgzdgm
PcJCRgk4qoTkWWubzUurwml+taMk0nEt0CsShzQ1dyVP0kiS5A7YHS+iL108FtCI
4QpBWgoPjguBikc7lByxyIthW+sGCBGJvmMQ6vGt76IMGeF3iJzqn/diOU9Shbju
PlrC+dxBUmEIk/gzIolFaGh2pVJbuJF+dbroKcNIjBpAYBor4LP0oQ2Es00KXnBZ
B3dYO6Yj7d7eGKnVTiM5CJUj/j8cCfdWHcPhuTChCecOnZJ3tLr8SOOScdUvOnG3
u4yI34qN7Jc40aXgVbqPkHifVDKZZzfBhh3+o+qsLfYhFwdiEkJIdDrbrQH//PoW
Dee3Ji+ALHcaow9FTFx764RAvUvP1Ew4v7wx/mnCE3RydtX+7c/MpKGO69mPPq29
yqazUuJpFze7DG6TMEieQ3AAPX2UCLJm5iXPnF/IWDfcDWfstcDTP0ZW5fe3Firl
fMcml5B/BmjFJzdgD19u8fI3Kd4pFS/jqG+YJjggqQn9OdiIXCAZ5JZ43OMLgVpm
LSDty2uMBJwGE8QMJ0EdkNjn+9DRKr1WgRMnfUsEh7jZAUa1zDOtF6BB6RQw8gYp
RQPc70cYOluMW19Zf0EcXrT/KJdOZh7Hett8zfaL5ptvAbbwD0NUjMsw6A96vwRV
NZQL87ASpsVEefmevc3FwWlsi+S7Pf1H2LzOtZT+LBv+lpj9/Eu/rP3UU8PfMBey
7RHw3aPTRPCq8NkDcqIkD9jHuOCGhpLm3x57ogXbiFjTleMbwjem3xCggfwx626d
uwFrsC4Hskv/+wfWjoQNYXjaLiYkYsr7libn5FpqkA8aYAhKDsInRYI70ht7MOg4
kqgDMZRNHCp/ymkG9H4018cZ0WcGcaqVpJVmr6/cxiUa1Cx4PqfgJIb/0nu49wUT
ZYoQWoipD7iCMT5zE4mvhhsZAglHJ5wXJAJRTldMXX1O5OcHyx/7YQzHnoWiPYxc
YhfjiSpZ/So4qn0BTuZwR3B1eSwz0R7plLlOiuCe2UCQR62YUot28qyc6gt2/Wi1
AA8jSH7wu2msgVoKqjk/VcqQYsbjbTBHKrDBPUDogw1STBBZyz1cPki2sSipA5Xc
yB1AA8XtJBnHAEbUy4LHlWsleKr4cDWiaNzdNpbiNkr7WXkFQ/kropoly1c7WffR
iQv2a7tvCT1nXalnuQ5U2ajtqznKWDvQRR1LqpXpS4eint4o3T3oZaYSH3P5uCu+
vj2pkxkJmya0AAbB1ViCZufymzU2I+6YnyJIIVi5uMmJERdHZCpY5WcHrZiPbLrP
1FrTyglGzOEWRnNmIUsnB24aAtf8PAipTh7p1yZHhYrnb381T1mdAtC7CtA5RTiB
SzoM3Des+yhzEryQtq1KqOwlc1sKdEst1orapjuzYIutLuJhxyr+M2+nokIAdZ9z
HEqxj4XN1KYFv6YW610y5EiZThL/Orc7pvAX1KB+HxIKK28OgKA5gSxniWB/4rPV
bSvBl5Q3HsG8tUgzCUgHEiY+KQh0YmnEngNEf5VHLi2+/x4Ffmo8wvePfdSr2sHY
hTnwUOARFH078XgJQ5CzAGnm9sIqkWrls4DYP5X6ladMBiSkR//XhepmOkw+YA4V
ppg0KaWH1GqdLVuzOVUl81KMsGxIEWO6Zm7uDkS2uNYFnqKQ0xYXhlOtFG/ewUvn
FlRFpYfMIlnxQ/+4A3NSRyWoBJ+VTEd3uPh/Ci/BaVI6wEToFW02vogA6G335SxD
A/ut6lhDLi/kDXgWgAjiniY0a0D9N1ACV/TNBXlSlwMe0PJaYGTpBxFMJrLblA4N
fIQMXjet75elY11BlgO/cER8S5b7qBNt47EYSJ4OT5C5lt7qJg+BZIVOXvPv3XwT
DYnv/AlSOnhbm+c76QnunrNDGES0GgdXDsrMV4Omss+E7j0Kkf7YlkFQRDCqP0M8
8Kd3YE/E3ZUTfnwI/vRKtOlxpMI7pZswhb4lfCgMUf1OnbK3owZiKiilAFRRlewV
qD6HOFuDdH26UOqQS+/sm3sX1iUztO+yO6df5zzf0+WqtvtUCxPAwQG66C/HWQx7
Cuon9VMUWa+T33IfmCqe+wYkr9VB2U748D8uQ3H15UFkp/ciFu6fAtou0p00JHjb
KwNOKdo5YnaO4XxEcIzRPe7wM0Za5bKkDMS5IPorz4NXah3iUGL/+zfDaddPzrTH
3dhROrISqJmLLa8JF6YGGNjZkcdu2+F0U9RHI8OEDoLqDBRduQqUgJNxJub6K8Fv
+41198OEf3eehg9vdyYANszZvUVVim97LGzaGriTOqxHTXy6DbMjl8VSfa9hbCWG
RUAuhKLJ2kUKKXc++SJnk4ejD9wwmWzc7Jdqb12bmccVKEd1cQDBZIQVhg/+bKoZ
htetmHIcIa+vLZk8vSm31lXyeucIV+Nt1FtJgKNkXDBAUQ+INFIVopijeuyCn3Vy
2wl8+ExVycsTpm+MGde8CsYbASR4jK1yJz6IC47X2v1TTuLv1Jxh/LQ/qJil7hYJ
qD+YMFt3GEcIFnWiVllEKemqzf/LZ/T8BMrra7K76FfVr2yck7iTneUXgTF/msjk
fL1UyqaY3Qe2J4PaQFgtBE3sa/fRvETq1oSbA2iu6OUqz3UMyvxh7WG/NM/pNHZa
nOFMpakBBOD7JiwUavxJZQ7r7awAuyNoZ5uAzkWCYROxBQU4P+gxUwt6tapSpNKy
Nzf3iUGz1LPXJhuVNQPO8shrveNVSKX5SZ6RbdVMfCnEt4Njx+1r6k2ruZthrlCe
ePJ4ngr2Pna4DX7zDZK6WaSbF3rQk3pV1DjjqC4wQpo7gGvEgDt744E/WYBf4wVf
SIDReFsDXB3TuzA6cgVASI5LXJtfnl84qNRocdXfQJIleLq2xhMlnsjmSUpuaPd4
NY18eyIkClPkMuxUfr/gGjsKOBaXWmWTozljVf/drZBr+O71yFuPZM7IruBUSFTq
9k01vFdQaT/UhGOmtPVjil4Whzxd3zRSmCn+kv8CQWdQ6Q995WQqCpRCABr6UeTV
gw523MZr9K9HpYeXhBJEkWEwN4x167b+DgCcjI7qCQrrfCMViTcDpttlQbx59Wtg
sD6Sfo+jINhyEc9GCLzn8K5SsTetB9uHSbFz6vMEkaRDBmh1pXGz/EhIjUSxQ/AO
Cy0kCCIn/eq5W2uhIR1zicIfmJQG3awLCbywtxgb2gDzH6lI8dwwuukEmLoD8eVH
FO4KR65rXz4GUL4KZ/1a0A==
`protect END_PROTECTED
