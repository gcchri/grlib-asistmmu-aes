`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evkY4ns+l4aU9fnU8PgKb+HaMm9gIO8r7lJZg00+VhZqZrp7A3UbdQxBrHdHrgs5
8OWodVACno+HY5WQInanlNLL+x11vuDch4pmKIYuAZfmfgDoOP3wmfnukp2Bgc98
rAqIw7zIVOy6lTdjA8IOmv/Leop/8ywbVSvOIUPY0yHgN2EbTChkLrTPTkurixhO
a+FUdwNTgZxe36jx7OT98xAG0+QUZ0Su2n1v5bWO30wkIhiN9fPbTDzD+ZUu8wBj
6fpSdoQ4Bwt6+9ecZC5KBnLRQQkOLvnlq8pdLpk/4FaPvDaFRxcGSOA9InfNQWem
Od6umoXtSx/eIqTECqogTDaZIhlAG67KlJQIx8Ykl3gzHdADmX+yoLAPltWONnby
OiREFiO9j4NmFSK9wKGyupJw+HV7MDPU4B/Qg//34GY=
`protect END_PROTECTED
