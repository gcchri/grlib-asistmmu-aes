`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+EnHRDRHIesITY0fNy4yJD5w1vUiYJ4HhGsUo167ZYKkH+9phnTnReVd9BvJpWP
SzTu+RUv/MGeL1YFIZrVO7faI1/LVkyNATyNTmlq7a3wwhC6youV/GZJVKfT5In/
JVbGSOZD6H7IQFN2qOhntbl26wxZaWSaIyxATNoO0aT0azNoL4GQMDfwHhg38Nwm
fB1IiK8oDGLxk68Dxzxk3RLWHSfCnAsK7+B3xk2UV2y/RsQ+eKznNUMrg7/RVnU9
LgshI8roRpJ8UUtGvcin9zLqbpfT1LXZEH50DiOz7XYx9jFk2PnbEZsxLlM+EFKq
2xq0I8zAm/NOwOQ+CO7oBCYOsMXDwvf1gyoP7DKVnK+thGt0jglAuAcvKAAjAH7g
0kqXzomrVrzszqz2LMU0IC7IGi4+MRWL2WYuCneZcgI9yrFrRwE5Wu5Wya5dhU6D
ZZtJmrPfQ1PvlcLmf7gso3ticLUbFl6HR52WOw5U4K39VfYc6bcCnfD7xV2GU5PG
ESdoQsJWUIesHyTElQcYf91Z9ntZn3sPoDVi+mBUmDR+fZ3c85UK28u1/KQmeE9i
O8d+Z9PxKLZ7M5+S7zpTrkh4lJTH9ORXStf4g8YeK0YLYAaIF8DQU0A9XqSThnK8
YrKn8Uqn9JM5VTPhsLtkc2PVQ8OesvmmcpFNM853JcjxDxs0MMsaeGmez7r5Tr+I
aMESAVfMdoevWlnEv8hwf5q+ShynJbAMkUCK5ObpBQk=
`protect END_PROTECTED
