`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qLWpapGWVUOtyY9U2MMe5Txfqy4PeYKCD0FVA7MsCB+VwACQ8muHu1rDrlH6112
B6C3Un5mrWln14SMFnZMxLfMPhAq7SZxgUTdQwHjW5EihuseTP+eFyM1DyxyYV+y
/teGiO74NtMUsdgH9Pc0ODv0RMVb4WMns2F8GgSmggDoR4Vt8zgwuZ87YKSYfiqx
ycOw8q1rp3njQjx7XKVVcNQOhQrtTZD9mV2FQO7ijYcdhI2GVlEb1eDq/JsN+iqS
lmejHxuBrkEwfhlJey+RbRCds92/qdrZ6tcvwWzP4M+tG+GEqW/mKedctuctlU5A
TxkzoArp9TXkezQCWSzum4QshQK4j1ZiWpi1aMyAJNUSGsKtr0ThhFDj9yUGk1r3
CjQFoZVuGmw6QNOIr1QK1UjM5XiMmjQnup1HgEb+cCy9FWwWshGTwPMgyFKjM9Lw
KoApvQNrfFXMXCXqoFKccj9XDA4CmRe9eI790MTlpcYrkpNA7giYnM56Lsif8gVl
ktrpoiau9hjQttHdlLhUMGDaOpTkU1Z81Fl8Ur+VQUs2oE+rsCMylxbGRMqIcV3H
j8ftarjwOxo6E3xySdrJWYIzyTn3/w7eQdpuECWOfvUbXDzSBuoAprzNGOVo64lh
YgntqY6eNPaf6tksxb4BYnbJeal7q2mgUFOmt3zij+NtT0OKKiiCv+OhjxjhnRCh
kin0el6JK801s9kWPjgtLYGL2SenADX1M7kromF+PC9ZftPWD0oHCJNFCi5OWaY9
0McN2AWckYv6ABSA3rDyEqrzaPozZJNCxI/YvUG42yFiafwbhFkSbUxsS0guXmfi
4bPDikks57PWFI9ALQnFfzPoVhD39bJSd0XWbfru+R/9HF7f6afxpXaANGCFEYbO
UofD2sPysk7etASaujkUWElRH3fLV+Don1fBx6pJnQH2PtE54rOQT0zmBGva+fVI
qBJxhKY4qnrGNTia1y1rw53+oNgZzP1ERkNx8S7DJLTrKL+P/eceKrkptDl47M2e
3zMIj5azDbTCYyUTBJp8MEHlg3s4RJChwDbVPG81KRqYLi8NJu+w6JNmlSbSw1ME
9K59X8t74BhGwTG3xDPH6vsZpXny6pz9p6mdwMY8GYY4yva2m+gq6NtdSxRf/p2K
PPbEM2kOEF6mqf9499EXvG7jN2vphV3LVSa+fJ00CARwY1r0hQgENMUZb41EmIWe
qlo4pn2FSm45LvlnM+Fi9mRCyrIujgVa8XVjeBkZGKSwdQqwRVGusckNoWc+76EF
FnDJmF2FKwoXoOvM/BhCXsI1ad0G8rVO0Ii7a2xp/+oJc7bCV0lg1INECWi28xOX
PwYjMddy0iqx64jsYQP0VftT+j2xRKgWe+cck4JgnAYIUZE4mmI75BS+5r/tySe+
nlOA9TmAvBN87n4ik/WPpJY46bpI3sRlVf08gX1vd8VAALwH2Gl0trz5Lhz22Jh3
HNfxE3LNfSk/YrTgcGd5soD7oYb8f3ZMkb3yj7dR3IrThg0fB0T4YArzaBflBMdo
9Dpd0i2/jByI9m8VQCHOfvXqJW5tkCLnFhv++Tio209EFkEdecf8/LfkNRpyDQHd
7k6KJ62Re601VXY+tqCeSRD7yPnV2dLe3isMNiuI6Lsnmbli1ywlZqN95tM/Qmj0
BsaxdTCOMjyBFJ6bGX72SgBvzgUc83BH/jghfG/sUHY4YBuwJV3UkgLyq2G8iw4x
o61U27J8XLPLQTAcMzhtdQQ9QSo2v8ZiaLbv7TWq49zy1ySoihys2QR3sskmVn7O
M3nN/DtCwZ9R2m1n6yv7MiG9K9kFwbwydAi8SH3X5Pv+H0BTNaw6gGjEuZuJdMEh
zwuyHFGTobkKLbOM1D6Wm+mmvmtSQoTN0WNiAhT2dg+Lv3Veplpz1MkpgywsSM87
bGKmj7g4qaC28QPiqJh01cQyZVgsikxLXXEUQ4HywPlzWBMHogrP8CdaAR3HCvIO
obcrzfEg73RCM5DQoUuT5+5MiE1OmmoTHlmVr3rjTokOKzwpwpRYkFUlb/fJaZm9
cQdL0STxxR+NNj92/PhB3hbHMsC1AHdNbS7QLpvDOn9kufklvMVJS5Y2ew7j/88W
seqN5TAcjwZiYZkARsI4W0I04RssreuqJY6KNG7S+7orK9RDwP2qmrBT7beTJ8JZ
nDPd7y0GI99zKmBL3VDvNmbvbnmpElNNTOxNaxcMg7kOVAEYpQiDFmJWUEfFOayB
2or28WeDNW7C+W9hy9SbBkui2CsHpaDJhUuKahGrE8pmCIxPDgONKYL847R2CJBU
MY++C8Djejk6JvOIa8Xo3n4S/dGacHYFPGqzjp4AbOS8pac/LgAXjwvi+ng3kRk5
rT3tCof/2zK3XP6i16Hkg+iW2KXLptIZJVwQJ7aeQ8fo94+UCB+hgGBGHEvbPk/C
8tq28hKkR4Ce0BSXOvfw/yQQuUi/KKEoI+A5ZFOSuJeBitSQy8PYeDdZUPrzWkFN
IhDtzUBP2ZPQFMz/KekCg0kVo9TcYSE2stZ9bSw06NQ1d4U5qmRaqlUICUYpVL89
WVlBfu0yy4fPiLE2VCUnR3apaRGmpfFvq7pg7ZbpTQQYhPaNHWSl5AXLesyq82B1
uChP6VKeYblZt6jPNJY4Ah6oAqrl7oaiWQjdsiG0CXLAQMYWxqauog22JGRf7YH4
Cly02H8pwq6Zpi3K5AzXLIYw4aDVgrsz/N+eeL+GY9o4xzv0ww16TL0jnRj8oE7w
xAMS99DMqjrQdNWwTJcny+h69J/pFrhvHSlA8a3C6g6nM9DiwALbwY22E/UBeXFY
4Q4e8ztQGfGHodg4xw7/KJ+D9J1dPH9C1UNJNbr4/4S/p0pX+XhY2pZlkelleyA1
voud/6c/s02P9Jo9zxKA/EbCf89d/1HKqTw71E5cmzQmAZdEAEDbuIF3aJ+WWQS1
nHOsMs85euOlYFXyYJ6+QFueHEFEji8qo/pzQC5elJKA4BiuqJuuXSIkmbXou/G2
H7CpcqarQlquh0cXXhGj0IwjTrZRNTfXA6j6FkqaFAc0FSg8/NTHtg93yeiSao7l
Rs3i3c8QhmGLxAW/km09OkbqQbMoidvTVR6+/Upc9KLiX2ctJlpGgRZMExwvbIGC
6WKFi4d9OU+zMDyv1ZYi8mhcZh3yCzL3HyLgKP6IXye7Pau0/RJ981q8iFX7vPX2
7lKhs+Xf1GWJnP+j/ZP9TdRCejKuNgU0OSqMAME5cq9JkBEEBU0YlqYsGiC5RSr9
kY/ydXKPPKiN3ki+7vWp4yTp9jN8ZHV1/Sggl2VjbKynxmbGdZfKaYMYtEhQtsyS
ttBJhr5W4h+b/O1rSJdizJtSwpX++pPMrsVyEPuBlT40/c6am3ATfOXNRrQkU+5d
+zg6iOh+k1SQigDKmxLzucZM16r8EAjzfPOBRU3fpWlLgsdDpwQ1q3sNJcExASBO
aBe9uGD7ci/vy6hae+PW+IGQr/peljac1UBTKF1rFGkduj94PNb/QmfybdUMje4U
Ist9g3YlZ3a9Dl6/v0olJ2oCnC1NXllftrgZIDJLSICYe88k3PXjzHm54DlBzH9q
kOqxNBBS1b16lPS1AhM6u0gOsfWTYbyHZz/D3XBUC0V2xBHx5oHJY+gYYQmq1wBK
rYG2JPjHuu3y7Khm9+Cu2mDrHPyJ3phU21QoLCZXBULe3rwCZwvduCU1o6+sODYt
24umGoVPXSlj3woBgBMK1LHy9U08B31qP09zfjWIq99AgljyvNceDGhvMYeRHm5v
fX98ws+LcRRZr1VZdY/l17elfk1s/ubitFLVv3M6oS5AEG03w/0fsg2AxctXhoQH
vWrs3utvDMiFtUzz6/DFji/IUq35TfWaoWtC1dZfP+jJgngPKW32gCq9ow61gpyj
SHTxUfLsSjrbhFcVjLXfARm1MeFLdwCNDV6Oag6CTk03XNvIIP41dsIv79YjqXY4
2G53vCl50lnzqb7HZcVE/r+IKPFWjO8JGbBKr3olqw+KZmmjTkm6ePoF0Pcfc4T+
AHb6FO21XpeKP+Hzd/OmLXGDBY0nBOrQv2ZvLquDfykMqGysz1FQOH2L4ijE5eHM
L6FocpEm7r5LdBvBYk5XIPeCGUhQGooWmBUtRwe0Hh5U17cPko5OV76BwcFvIUnf
YuiDB4VExS/liV3yVxaNNwUFrLNiirE79L+ApUtdZ9URsm+nnr51EmKu7Od6n96J
JXH8znBizPq/F7dG08qyf3PMw9Cspt6Xe4clKQ8/GT4TMF+Ya1YRQiw7p2erfiki
lsNjT5mNdH6UQ1IsuN8BoaXUDamRn9SJSP8GuVMhp87ZdiQv17HdkYxLpaxpi9ef
SsDJXUxOpVY867zYHvN4wEB5doJI428RjM1MlEf7Qxo81XQzBprFZL/fpWDIJFUM
ejehCrsRSkR3faiHYCZuY9MpKs4rNncrBWduosRwpSzFHJoO+mEgsGPVn7rd2YJf
XC7RWwRhNihKkiuqpG92m28Y2VEyJYroZHHrjo+spbIoVmturFTN0pwgeC4HXfD8
9b6QZnfHzwBtnHCj0aZzUEnns+hkI1wEAT7i45G14hh7XzZYBg8r9tBIFuUShFjd
JhJ+OO4M5gvAC9YDYDKMqxZ6dNLTmW+Hl7bpHyAwMRi36aKjJKCJJ0hHHEw/Bhgq
P2MioNlCMh+0EombWfRB4oe8zuO8tMP1KD8tWqIg57v3XdSx0+RHQmRETPIBdODZ
PRECOYCZ49U9Ktaa3u9HPg==
`protect END_PROTECTED
