`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WN8t3U0N+B3tt6XnykZsVJTqV2dnJ094oRnVnb7JkkaatCRROMntbwebAGP1rKml
z9jstIWulsiFRVXYhP5jLnR4PYhhFYA0cui971WGOvLKRRKLM4ch4iN7SnPE7EEl
iXbJm6SAbg6WKu7zZMIOWwN/y6t4LBEtL6Z0z5YY6548oKnhG47RCRypT6as6Cdq
n7giC4Z1op8GXa8I7m7ojLFOzU7IS4KrgjCgjjDOhjVjVRIyVjC3IRHhh2XGul4j
hAHPPoZ2E5l7mZtveLY7Qrv19XYyORSuGB2H69duB9MWQd+oStj6sKibEIkwmReM
Bl2aARj039fuWuHRud0g+bLFV5TXE0ofTWqatt/0721AEXCH3uTiXaXKngtmLpFb
bw/nRLqiJ8oq2SCcm7dLuD2Vvz5N5Zj8kmfKoyAJqbn6QF+882gmqjPWltKCbDXa
mYCmzIaMY7Z+WRMCYEjPm6PXS/x5ggK6RbVm8psUbdSZcI2HnEp1UEdeJfnqY0Pd
5Ok4wOCj9fvj/Yazr7GfGP2bPF+GV8/p+LDpzsgsUePQwoLLwZkSBxkxumZJJbyx
QNzkTVAsUgaZaPpPfb6utqO/m3gOgD7I8wYLfiKl2bA7WasoDvUeCrh1bH/pw2Sq
923x+HVAKoV2w3mWHcUPWOvndBYLtp+X62B+Hw6oOoUnW5JmiKBzvjLcmv2bjPxt
yEU4FaqT4jl0dDoMwLOzyISfg9Jlw9lcYrLv1i0Nr/NwsbF7jj1AuEuJN3t4ADG0
A5KMhOzAiH9L/TJ1sLS5RsSdqn0We+SU2YpVGelkjFNNxRsim0C5UJc/bMOMrZWR
3doUw2fiE08Q8qitQWg0nA==
`protect END_PROTECTED
