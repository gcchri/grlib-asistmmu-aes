`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aqj4NT2Jj/fR6zdi6wRi/cEgT9CMsCbYRn2HrfSM6wNk968nJrD5E9zlEtfJ8lXD
OgerJhIRxdLifdlFSZVl17TDFVi0TO5uDGO5XDTMTd4QFv8eDCMelKxtLMW6e7sg
Q1Z0pSCACkEh0NoKw4yrQ7G8hrkUqPxRW/6hDdaPslX4FytCl+AzlecAF8uepwn0
T3AZZ4+0h3Asyhg1rSTdCJJ8wuGRsnyHmAS/F4USZUM623qToAC/OjuxTxQ6KCDw
95063pzBQZIJaWUCQEhA0vkdr7x11inH0Fl6GuOKp3N5fafUyoPApYYuxUidlpzL
N6VYLt/txIv8H2Fwfth4PYW2GaUMeC0NmXg6Avuthm2+G0lV4gvqBf6rlUO6xFYt
0yoLcyOhOgnju9rXhptOomf2GjCXdoE1ESodZhSOz08KU26raUIWYY8eMGJ3n4J3
rr01WyBSrLnd22h7db+C8gCT21N8G1UVgiuN5hf5y0/owokFk440vrylzdRFm/I4
yWlZ/OMc+YF8DSSsDO/Lk50XaThL9QgK9g2frvV8vHnoLBdqJ1e3rqqGFe7jN1Ui
HAEUz53hDkmMzlG7Gol7wcjuZc+Add8XiGQb0DyrESCUT4AQ3U1OaPWs2XGqQ6nn
hD0d8gVuaXRApCgSgE+ynsiTIWAMK5qOGFg4bdISvqQ=
`protect END_PROTECTED
