`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3MvdD6WH2d/gBpPPM6bFBd910W/odbMqelggfF0/yMqsPzaR13ZQtVVumLyQPDvY
DrAp1/AsEkEjngZa2Gbte1HJClNgAy0MH+64O0E0lrc7A8AD+SA79+yvkFFUg3hM
EDV4RcIbZ5tOSAGznUK+m62FvVJWos/xUE4D+d03R89jRUQQyBXJtrpQOg/KD/4w
N9v5RbIqy0qApM1KZbqCqav+3hrG4kQobBWkz/jj2bkIIyZyO+GP9x32FXUVNphq
ppCrt5eNFRPRl7jOIdAtpYKlekFw4tKQ2+LkXFIN1j1KaPTKixuZ1wFiv7xEk1hD
vl35QX6K8etUEj6PjjgJ5UpjShpyETF77Co/0FGO93kn4Qyt5K3gTDUovXd7Fyzl
iHg3iZeSulN7WiwQW6dMiDmS25aSN1EmlC1uaQZ7/w0RnVdqczDNoAMDdMZGD/nk
ClImk0/6Qo34m0a2nVGQ3H/Li4TyZlkjNYQtBiDFsMqd82oPAQNeUf1JZqTM3SN/
/dCNSf708Xg8cJhQGhPl6gZsY2H/txViofCgbtLxjLB/+CZvk+p4MFtXODPrhe6F
61DJzIMYE7L6GTNHVGgaQoqB2tsUS+8NaiNm7Fs+aBnXABE6FeiNGl6/ukv+8PJp
udhBtUlXv9WX3t6y3Hxb5t21Q151FV2VahGPIRADtk/0DT4C7p3eJNi/fYyFeTM9
ZlNPvpd0BoKaXjSXk2Hf4cZW11un5PFhRQMa+5974epOW2SHdwBofw2fxJurAWxb
3qydtss32/oDuHckdm5iMD6iQ5XphT5QgGREppa2lwZJHqjh09vUHiMAzBtWwCvc
MyIQdqNRxlhtio0KSlJ62tcIPt5rpbRwalbfyeVOqxyk5txxtbsmb7vmzTzXnAOp
9g07BB8AokuoED9CojwVgQ24xiNM6Olgq6SBDCTUmR9pA6SvqIiMnVAKqHlkc0Kb
Ae+1a05J0tGxkaKKZe1QhFBk6/8y6Wtl0Di9JDtd8k6hN/Xs8/bYXRGl7sS1sSx2
Sb7QWoWDBBn7mx8Tl3I9UFeTPZcghDsPXEinTzktFCqopgRIMZo2Fzo/an5yixb7
BsHwW7DnfazFccPWcpAeoR3Qu5FkM8+oLUY3WYoiwf/2nuE8EDXqxAoRHNP5/PSo
0syjxG4KaTOdaEDEqzXC0z90mpxjAcLssU7ybamyThtM3tqZVn2eRXRtIgGcVzOL
InBHfemKtOpFK6lPNRvhHNFX3vQaalVZUkoYJWCV1WhQedQ356DKhxZxBVi/uNCr
MRbVRaZyHnETEwmAfZUhiBRKHSEEA1nKoWerqxmi9uQystApLEpI5iFC+bdJ4k1q
fyJx5jDElDp8gwt5dnoHLdDBbwbqbV/7kE71GzdiTX/ol//CA4xeit1RBXv7+ZFW
nFSeeO950O3KPUWp8yKIndxgZZWcrLEoCbu5xYsDzb+L6pQf2CLuAOYmHXRly/Or
TNBxRb7tUO6lqMWVc29Ktohi1WCPqwPcKU+LFfPYnDj3PSW5wCCX5A4gvQqSEzf/
Heh7KTjKI86b5/W/X8sfsTOn/lfrm24g3FUSwdZCZ3JX/KShrpFu12gSzFAhWFC9
v+mulcBdzSKZabLIuuIASesrIDGEPT0OhgXxdQBKEHuJZZLlH//xTSjBZ6Ct7LAB
mSlO9eHfozm092C31NOqRgvEdowJoGpdlw90LO1r3dxH8lqKSZIxmiB6hFmW1UPo
sPwgqkVV54jWumTcmHCngECOc9zacGkGcnTsftOe2HezACfmGQq9DdSWuFuB7EVw
K5PWof8ArFB7oj95eUQsRh47xq1ribglPX1pl0w/pwT0UwwWnoMEX0EJrucdo2+C
6ZQ4/qIjC5G8q9rQhXtAOe3qnzgSTUEcDh458yec9Lh114f8AZ2rSKrJtzzCKAA7
wuy3TaJyYUvWWBjvFXyphEfiK1G+o9QrWYWtxsiJJl6GWi3x3kK9R6rqUrkMSEen
6ZFgCYQGZrwDhuzoxNMmb1hR3YP0Nv/mVTR83ycV83nGdRl5mxtC25tGqhDcYOR0
Vr7LSV/+bTcqW9QBPSQmsVAobmmvbp0OnymEcG0YZIbcXi950Q7K7dw995NGi79a
TrsjIV/8O07sVFTgvylnTgdDFCs2blH4hd+9Bh8ttjgZrXBCNvddoVku+QLJB5SX
XDj7hpSlpsE0gHAQtrVVNiguHWo4JomZiMKYgLWh3anXGx9DF/KqzCZ9mQ5Qsx4m
8nrGzomVnSgmK/torKo7Ir/CQvHX10g0aBxcB7OZhB6/PJL3ZQucU55iMU1J7Q/y
hgYghYOwa3VEiNQ+TEqshGzGixBvaeWCKqj5jpgNqTMOHgUtaPv70245KQXikN6/
aM/8bK/6LfS+w+kViE5nMEK5Tt6Dw1s2dc3NLyz2bBkzeJ+x7U2XnqdkkBKqMsV0
WBJwnO6pZIHsQ+L2OpNJfr3PfCa1SDIHwEzx2GSarccD6WQK8AkjXNBfV21/Qns2
LVP+Zw+7bwxRF+OLfYn54+AZTUlwVFoo+hprD2wmlqLTu8ACpvo8QsKydw0OYVMl
PlX2mNMpS7vMJU6Oo3+KTiZOtDFNqW5pe0PjScscn3N0zFZX6jLjlO6zYnGe3P6m
8874ewyYsBO+FJ16PHDYD0cFcQ9+KnVMCMFjjTVF392Ih63urXNdHwbIbzbbzIR0
wUUTP7Tf71m+Bea8jDQRhpmrXr8E9oROJHBsPaK0G3Vx1m+84RnBloziascmDGXh
`protect END_PROTECTED
