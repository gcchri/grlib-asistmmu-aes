`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JroF+VfYeTqwr/tThki1rAGyoT9CyuB7U48W90oipZnkFci3cmTIn9ngGHyy7KVK
U0co19ZxOsB8ZIp3TggrGuYj9hzRVEgQl3PN7XQL/w1nbzCnkfZA+cKWGhZScyMR
KX10vjnUCTTPGMgLf8ROuIfLMkDeD8Gn47VI4fp0nTLpROx5E5EFYri48fnROcQn
YWJGlrJC179Os0ByOQVCnUYUHskkov99U7M9zeUyV2T16WCFdZl/5DuX+pVGfbgk
GHF2tZdUE8QiFjar6whkhH3DQBRMeos0pzZbR3D6y77ApmpR+RSab6NIezoPEw14
bFnpMMFL/0s7lESafccKu1+lgOqJ/3dSblh1KFfoZF98KJHJ8lNJ1qtC0du1cmaT
2ZuSJp5oMcMGyDOG+uzGj7NuBrX3OynZOnGN+yERam6Y0eiPhZdplYq7S2eK6YDg
i3frW1AirZCNfbu+s/Gbk8Z30CtOGmxGyQqdKkheQSAkP8eXMjNrz267yYV+9QQz
`protect END_PROTECTED
