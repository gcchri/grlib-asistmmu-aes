`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2s/wNHOTecCEVD7NakoZaYQZG5Gx3mmnzDSJyKYU0IbJkdWW0Q61/czF6/Bu9V+Y
3eoPvhvwGbfQ2D6MpjDDdqoNRJtNZ59NyrOJH5oUsXGPlO3YylNK+f7bNWVh/khZ
xby4xJbUUyZDc+gOcD/G6DmW8GbfSibxJyoyWvgHzIj/qsUNq449pZDcaz/Kg8YH
8LoB6AQzy/Z1PdhU/agrwsynEJOD+I9ddyoi4fwoidogBlh1BiaIE7gWj1LwIgAm
1jfBN8IV4v2NPS6pApm9fY4bBJjqb+ZKosE6MYCMDMQ48u2aOtwoLuAJM9z8ZiaQ
uds//s05IMEOKMuTrMmZmbmmGP29b+iVyN43PfHR+tPYLXm6d4fxgFBS4kr6nOiO
jPJTM8q7TWHo3TjCyE2a3g==
`protect END_PROTECTED
