`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wvRP6eVmvWgWduQ+DCL2j9S4OOEkSRE5j645W30AHys2qosU2hp7pkmI2CLKILSP
NO+zjUAkkbEDIJuU8lspW5Fah26rgph5TxTAIu7wDs4H1+tsbXztNNl+IawizePh
cu8RKz2gJcAo2lbQfGXqcLO5zTD6Q0pQU6NgDsYe53351fEloaoBJ9QThcOcxblt
3q9/AE5WTAhBx/ip7bEIP2vs/ck+TPBSbf5QzBozzCmfxn+IrXMxBOATTlOvG00x
OrT3yso2/Khn54EtWkwFlcK8e+baHPEmRM63tWOMZXvT5BSIPNiEv1coUaeaNQmz
`protect END_PROTECTED
