`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7VowreOenfwMFYUi/2jiSo0zKcHHMiJLs2Thu7cAqshOE+9v39Q+fZBAMhgEqQOy
iPv+CDbSFt2YQOSGpUnum2etZkDtaVEazkubaSIB/ckRHfCsE6Iv3uIidCuEp9kc
J49B4YGlK4DPHryAug98TAdoy9OoK0BWn11m6VOsC+etIEtxBEcD2VAXvj3fRKLq
Xr/O4FHVFyV92ACQvg0qoOEG2RqQwPASLYNx8zVON+bAwDltajwfJnApyOdVWdvm
6iiwJQWNHOdcNboMCKbaQUmsuIybsV1m3tv2irEGdXXm68X+Mo8g/E/tL2R8B7c5
hrBf6Q0YARFtWRSc0aPtdx3GdhPbbFeT/4mT/JUI71mjG/Q4JUyAJ0lQR6ZPHLFC
i6d3zm5a+p913ARBto4Li7ZOC9gKTgJvWeepMfBZna8=
`protect END_PROTECTED
