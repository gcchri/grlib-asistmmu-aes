`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndnoJsbp3V6GEOb9r63/faiIanv1EBCAcwY8D3Ek0ABvAnSfRA3L2EAgTZ0Q2vJ9
H0sc0t94UpeoxlzzagY0uSZQBPZRK1hNvtICSMxLUZrInv2PuJUIhe3MJgY4b7O/
02KBm7D3GspOjrW4yTjBEwObamhaoTd81ic3pZfJyKzYw0/8wB3UKfd4mozCLept
Ux36H960KdstG5uSn0FMLvM39RhjUtn69DaXm/K0IMbR7jV4lv+/vBvMyYDQEN1o
NadIuMZF67IR8wHXUhchMO8yyKV+KB6jAJZixzHoAq5xzjsQFfU6uwEuteD6kO+j
cU3fV7LNz5y0yJeRPkqUZBGDklmy1u4TzlB+RJ7vkemgaloUrGk1Hcp6Olk9to3L
w4u+rCWKIOlqSBzFtETuJXizK3gdmxueUiuiVWQ0lzc115s9MSY6qv4kS3pbRQ6O
faP4tLWZyVaDFlOfTq5xxDIpFglwHBaCTjRoYjEXOv/FNCSVP6aroSOwGE9xZ3wU
277lBxVdYaDZIWoanM8+9AJONblpo7ZFiv41UDCwYN0exxTGsWeVXVns/Ry+zojy
RoUer8AC8C1+uSAdD9XusaNRHxV85H05QdPuGsyZwIyZQqzOlj31tp9ZoxNATvZ2
FQhstE4Hv2WMjJ4emcUI0jAirtyCyxuQwQkAYuoYVEkTGwFrkFTP3llg0wvGVDi5
`protect END_PROTECTED
