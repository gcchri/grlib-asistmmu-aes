`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YI6qQGM8AK6k0K+FZHG3kmeqA/+yy0jWvp9wgfG9cco5l988r4kLmRK6II7NLVkZ
94JSeSqHszJHQEirhQ51Mojg/agMwE59Ypss2L8t+H0uUZ+9yT7afsHZB8tEtPxe
RFYkPuDgNlKKN7xMLcov9RTnQV76B3eJlD5km/ph/wR9TSp7NBMyRC/t9kuRPAec
ADR2bLGhcz+eBP8Tg4UX4X+nZ9VZluaXmtTFItSeFTA0UldpVDdermjDPAmPPeNV
ys79rDqEtZZoFqO3BFFt8C0RxcjnMNekFTNq+wrfWQrk2wFJmrPkbxjjrgBIG9C4
II/wZ7vlI3v6ZXqVIuVGUplEcvdoXe9/rQsRKmpme/TyLMAYnT0o7wfcDpKIo3hn
mxSU8Oc/gOHUlLTmADsPpufW1asskAaAN4W9IOTgJKuEiVpyTpkYlqFcFjlWwL/K
huUloyWv4wj+O1Aydui5i0Q0rT25atpDmyp9zjRXgy4GzVIKAwhelbQ4smoTFCBg
14u7BE5qNykAzvIdglLVy8kWpN6oITtTOCRpgyPylDs=
`protect END_PROTECTED
