`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R9n1xKI/5vsZ7sqNUWuUqsvvJslJl3T4VL7GIQzdZJKqA1TrDJmFwBd2hLnoEZMw
cTurNLWUoZBibxZPpFQN0C87HaCU2DeOv79FpIQz7q0WVNKJM229q+CfweInc/Go
E7ISwjmolGktcEDw7CqLUO+sNeJZ2Sp8O+/LlEElmatMfR0b/JY7kJG+ir98hF1v
9w+ENr13ICI5EbmBN3+UN8vOQn2imO4mRrPDYJYQwdDQPxJDfOJzTSE3YDJClxOh
Y+Qc1gYmiFpGjDIqPtbsCahiVHIxUt6WnHywdmkygrFwOo9DMpJKDXR/zFdJrRTC
I6MF4FRGd5jR00AIaqSnTpW4yWPse4ItL+/4Erw5i8JuRPg6amUIx0MWi6Ll3i+O
3gXfpzzBq3bQ2D54OBBEMdBCWP2R7gYAeNz3AsDpTpz/H/jg05agD4KuHsX/y45F
OWDdhI9KS4/s3CozmtErkYTyAgR1hsh1CtMdel/yW6H5uHax45w+anWMUeNqtbl1
e9O0ENPfZqkg5gO+5mj7Y2DM0IhPxXOIT27s0I3FJPGXsvT/zaEaYFKxDX9XwpuS
nz9r/7U/dLYFHcUwyUdTbskQb66aqcTjtzL8HBj8zhuTx4mPHJ0wBmwpPpxjQTKK
/lyosNWJ/ztjfi5VWzT0HEoPwpc5j4srO3MKEtN0oqETH6/08FzqvijnoQ/SGn9S
IEVOCqS1Q3YTKCmkasy/F4geOUEJnGbx1oh9i9Z6uZMIVHWfSPKhyA5iAJ1OELuu
lfQZuFyJajYunnJaJy8VVVGaO8xleR8TCdJXEMrAHsgDmigyaxbK/0GT2kHJJ8hF
RS23IevET7vvlezD2CumuQHAVIV55UMWZ6Y7mLpAC8q+DbYGY/wRQFJIjTs0DfbX
wQwN8e+HA6WsI/xmfz7WJXlkE3rRZOAQegsZiID9R5Ua2vKX/vrxxbWDmKOghkEp
3Yg7r8pR3PHk6s2FZ89DmyGUDJOo0JVe0twFIhZBuW/BnJI66S9uLDIl1J1hChgl
+QFcA+jW/YCEpfz+7IR3WVYyjXrpbwc+iZqflRd+NVQGzX7oPlrPL+819D+yy4YE
2vk83InGCv+nXCIupSbdirShf0H8faVngViUIaZmzJ+2RDuXxZME+tUpB+p+XTtJ
/uAc0k3LvvKGF679KW0PI461RA1GgcC3RBOTQNTRhC9y/s8x5CIE+zvZSY2FK9R3
QoVvMNJyYmnc6ijbbx0rTKMD498nAQ1fyYeIg4e1wrHtv3Tubl3YY0WMlnG7/nsZ
lwbND+1LC5VmUX0oJ+wPBWA/U8a/dRh7lsKV2PfqIQhGRH0TXutoavNP33pwoo4p
ZNgNcKixZ9kBUZGj9XcrmrtHUW/DdJ21IDpEu1ueR/12WFyb5dGO+H6NzAaesgAK
WaZya4RNhiSlhQiwiMldPK4fKLrWZt5F/4L/4utSw6feaX/WP16xYiAU+TWFrtEA
VUb3L8DOs+BiavJ8QMVmnuE1fapyuxsHRle7cDsLO2Pqg+mdN+NaSxfJj0Cqws0N
mbTdYT6t8wjkermuMln25cNRRhd8kRoyVovbMHIY7xSYUtUOJtaOkpdjk6Jr2PnH
rbVEnsUFB6NIS3Gsw1XA1YksN19yTKap1fhxGLKOIoX8NYwH3ZG8ZfvrKySgG/lj
Jv76YeEPFjf7pwywv1ld4xbLAKxJTQZIzkNTWsVg49LSWwc0utnrfE5ErHifJ4a6
qmVUX+NHWFN+D9FdSykylFDUK8lg66d70Hsd/vwVQZR9g3qM4xPtl6IGzlacvwqw
aL5BCrjBCZSTXzih3RmGnPNYwjroCkS018UsaD47ZNI3fNylNkUbYJl+JdjkgMyG
qPtMZmmgdBhFsNRQ/vhC8/irsBL/RAaLMrQ/e/AynlteceDPPGREuf5LnvtQsEur
oXlk+rr/1WmI+6CjsuFzLSYgmgFbbdh1fVtz57/9bbJUa9x/9kUul+Cfpev4bZBN
ynjuVNRrHuFINr0Y+5Tv1fsqg0ZA3lXnkHQ6+k/VLwWN6mPUNgwbLivQIVWd4BtB
U4bgI/U8wuYTQ/1wqNtKKHKp0xXFpXYyTQzvRsAfaJkpQRc+Fe3RfLYlK5UMe3Il
e+DuIKacSAhq1Z9A8qQO1srv7pN473pwRoNq0zvAqKlhqctUFhJ/30VWRrMQtyrS
TVGex68rA7TYaUjs+miUusiaxLH/EuRl9sTrrMnTEKmyGPkKbP7V26yrKumERvaU
3sVcZEMS1fsgbDs0yPbF9y5UZLzt6O9+BX7zvi+evBDiNLuTH9xF7aQPt96E2dPr
+bByvP13JiKnAcMgy13kibF4mOMPDNnrG03sRoYHa3QfJQcczW1sNOvLC6c9fCaN
RNLL1bD1bD5M0KhBGonzqtObbsNNdbno1D9Niw5CpTmuifk+Lr22xbrNCry7MiJZ
WHbB4/QiQm5ouBBNgD6cXIH7z4m/r2Bk0qsv9HQ2ZRPuOoOm0iFoRLuDwEUqHvqJ
YJEoTrsxvz2LRSqCsxHtHABIRo9YvOQz9UK7vz+MgnCqEFwdrT6uRy98fL7bzt5G
`protect END_PROTECTED
