`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UFYo0UQi/3qq7daPGKWuEzmluNmHHXBWMmWhn/dvYUegbqUFAX9ER5eKBSS93khv
C4jhVWssxPrvQONAwrB0cHihUqdlSG2lOblCuuUlRoNJu3NGWs8mQm7EPf1eCxWH
k1SMJ98cV+HklSh5DryeY+wIPmdYU6SsnJjbqHFtXdMoZxnZiiFB3MGes5Od+Cii
MP/BIQETzWOUFZ53Ka4LW/hj2LWx4lPeYxxUAVUfPg/VpJsY2ftjOs1GabaFm5+c
4L5Fuy10jzYXafDRqRT68OM3mAzwP1SvfPgyfiaJZRZ7xKQUNiVEmzzJjd5nhlNQ
wEZV4YjB9ETS6z0huwhyoYwvTASTRJPvH4jU4HiqsBZO8y0AanRaz6jFar1PKh0v
V3HWfMpPKaszCwZWXPs1GJkprWBUdmaQb/BH3g9NiimLod1CQ2jZJC45Dvz4zvtD
4H4dPiDOaH+XcZtnSGxjdVibcmVr0NjdAeSGS4w+1fRni9bzL1WBa34j2qnZ1lD4
f2I5Pk5KvBEC9R01tRJIbAkKHG5D1iAKafixrxyPc+O6NXIkqJ4zhs3c9cTz3G3F
ks+NFsF9vrb7e8a3+XcZIvJN38aAkZ4Q3gW/zWh5cixfC7r3Jx08Qp+9im4e9oNJ
foZ/k6gYVvmbHq2CLR+G9w==
`protect END_PROTECTED
