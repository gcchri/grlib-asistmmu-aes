`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1NcrlP1DDnPKkP14WIlcr5q1rb/gS3y05z4p9727YELv79aCIKOkuI12dqmuES9c
TQck2uzx3SK/SrW34uX19svhTZl9W5881BOPOZ6fwV6yuMHPoIMJSafgqGkSUOt1
BA4f4R1Fudzftm37AhwsP4raD/5mdaDwGgcMuNfmQdQ11Fn2vHU4MTRFBt+xOpnC
gC8pJmVcp0D1sAenQ7J7DPLkOoO/cESTM/6LmOfh/CU8yda6A5T8giUr6NsKuYGI
o4lyh4SC1Ia41FMK52EniD2CpldWA+RIbZD4BthaBqYFN+9p6JkvRw0eTRKKGAdI
XSRzJuWLjJs5arzduhRwhqeKECx5cKYYslQDpEsETB8gyB5DmeujRkUuMPLXZhTc
4iEEnAhu0S7IdKVejZRSuBxaIwMv4d7ofK95cDd2LLEW5FlsZRinsO8CIj98kS/6
TE5nyAZl0tZr3EO1343smoOYlA++yglChCvcoR1AlF/rdAJmLMwywzispc2SgQZ6
z5xQnCo6HSO1QbPxq+NHqBLSxyYwMQPGuyBWAeXNpIIX8hggnn054DUG0peAjhtZ
VPzDF/DDrQnOU1XRp4ZS/Lo/zJWDLkmO6S9alofRtN7nDybvAjkxm1vRttbylT+z
ZrYhODfr9FG0vYJ6xvRdaAxigX6f6NDh3tRlOLcc4WwGJLhD/pjADrRytgC3JAkG
rLuIERFyqnDw8qCx4NCqbaQXkqwemWKbMolG/15YNKfN48moQkwMoPlcyq0PfQ2m
E3ntdgRCQwYmqGsckDe1VCMdBCR/RhXO5bQ0fcwVOhM2dPtFAiw67Sici4vpnBDw
Y3NH4ET0Sim9PYUYzHncoUbal6zP6fV/KsV/Ow/sbXB9h6Ex9C2CPWwg8d+BkRv6
fGrtKK732oCa4G8YprAJMenzvJyzcW/lz9LC37VaY9ii74ZiDAbudgtpFup/Q8Tg
ylsI0GSOJO8DkzATn8/7FhJ9pIHJnWKgVCDoJRw5/zA7socykAU2Q/LbwH8l9v9v
UjxpKgdiIAbpOOGIxpwkbO6voVVOnzvgb3QWM/1YqxkJEnS4qfhmB5zvxV4QtaJc
Loa2EH1LiuwFSQjdDk+XY4rbsa6YeLzAybcDRgCkLfa5s+GqAeB3oB2uepZ5VLmc
0PvPl+IU/HxnD8jfcLe2fgnjZBS2H+5D2wLwUiw5sxN7UK7v6wrmih65ho9uzZxa
Cg41Bd6WWm2KNEMPbhnRHNQiSHrpFJtjyoC1RsshQwLzMVitKkPS6dwn2Sp/V/YZ
SYHQgRHw35VNBRVLy3Sn+jKBNAOSSBenAXa7YQUYHy0bDw2LG/dxonsf2ISLQr1s
Qc8I9ytqNj9zM4HyZTMZmG7gi9xzgzxJFT2aTEI/hJa/KedLRBE+gZO1GF/yxLLv
1CwnSpkvSmO4yV51oXuuqeMCLx5mW0f/hCdwdEVywJnklzYdF2MNj+M+3xhm8GIf
uZlkQKRDS/HsTmaKXz5JqcOqlu3QDVHphHYLrildYBNH8NNAwa0tm+sqAGVgmM0/
AS0kvafHEJDKPU7Nu4CPQilaeVGQys13ZKWSXYl3h9HGbAug6rjDKIhQTyyMFnd4
qCXeiyaxzdSCIkM+Q45QDp0MNjM7QP1HhXXqbG5Qf17OZcehUbZe8RskCOgIcoPk
ruwHUFvkOqk7S1Z3rzhkGNOFSAHjWIa/Fkl2J9jfdPihPwSzoZhUPMua6JUZDzf0
JHsH3Vr84+uXK9b/xLwdFS8w03wXzycPugRcKe/Lk7BM+2r3wUSwAc8pKfYmN1+h
GkmsUXmHJVzscxVTxsm85Lw/GZwHNVcQ30a578D1Eac4uPJstvaKuToMtcNl6vRm
ryuNiHaJc8UJp+R3+u+n9MpJW+sxpYBwdOkos5PASHdwMWIdZwElSIeWEaqugPY8
2GVMkHnRItN6KMZoRuq5afMrjRIDsd8p3e+i/2kFY8E8soBhFFB4hhneIV0RD4uy
ZW6+L0Fs2xC3n57usHF6aYpTN7xDwMuajkaIflfu+s0GWnvAlVBXsQ5+7FrNBjvc
FfDUZGpRWEP3AaGFEPsZw/LB0njpk70FGWnXhOe2+56IZL5q1jmRk3JM1GLYadGO
kpW/7rC6R5qs0hvPQTLdTP5k5QLJU06Ba4m0hVXjx8uFxHh4LTMapx6t+0wHsFRq
nRVnP0iN7cBoFGXy0axr8HYKBJtzGBvsKWZd4SIJrfqsCVvguaqAyu7X93ZQ4Dm+
ErK3QEUd/DixXsERYuUKnyxFyB0CDIfSIj1+kALHf5d/5m3tUoMnPH9O7pR6AzVN
lhFiK7jTL+5VzqXHXd3OQb2VPQP0KDPSRJTy/VAhZSM=
`protect END_PROTECTED
