`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRul/vHfSlenDki+qDFzpnAnh7NA7XshzqoY1iQfwPfd3VEJdWkGROWRnknL7qSS
1F1rpTfgVIhCepEGza2+DCqaSwIReBnOVgCRaGCwzSKohE83Pc7+w4YLUJRZALIH
/6/yuDAlnaBZflTE0Vg3h24pBj9L5vInlqDfRzwVmSX47QktY6ovORuhEoa188Di
VTj5CTqDssHl5uNlhJsvR8YHyKyGZEHfYqCH1vsUyfALTcwEyiDhaeXABozMJHmx
n4PgzXF8l1YNgHot5fDfb53TSq6+Wqqol7920wdPUJNPmyRm2e/W9gLnqwrsSbjn
Hn06iBY/YEJgRd+B8vT+m2MnfmQc9kwnLdRDdezBfanHco5pL0mxBwSdx9AWz+Gc
y3Bofho+AnQY+CZEEZQ1682DlAK3Va/3RhJw4QBRbepWC9E+dvEMQAGt51NLqFY5
Cg+uPfKSrrBzsi8/0U5Ol9fRyIaXZ6oNUAYq6Ddi6fG7tu51UWkmOxH3tZtGeY31
CGwJyDCmfz6RHWFaaPzfbv1p8Lv+jtE/F5Ma+H5jmXvaH3V1dcC/MltIBlYBuYAS
i2jSEGi2fytYprz0kErVFuHIiU43exvySLyZmjhwodalK49vl6b2e13MrReBP4fs
v7svYIA1ZkvFPm3sEyCD9s28zx0suxtJyqr9kdtAdIP/O5+0BOOs8nGONLBqhMJN
24bxO4au4dnEFnuXfiR0GM6q2aAqv+rrojE+16QizyK73B8KnjgiXLqAo/ZT+kL2
erd2N2c5BAje/1cl7FQaYwtfuzOEH6q50ZQmRNxRHrOh9OWBUhdF6AWjixcEvjWi
zYpmYyb+5ednv8ykkRqLBGPMbnABl4zWCka99oK3aYhtQAF94w2tVK9F2ytk5u/H
f9hnyxvonCNGznlqiOLw+Icq2M+ytU6OPA5Ul7McRbts0SXUwGSZyE95NMFg4MKG
dQ1LDR0RltRXpMD32t82Wmp97oXNazE6+m65Hc7hXGpwoZ78sR0ldA/xOwNpa7ol
PDKDdXjWxJMZdgoLyWErNjzF0zShYiDvHnl0t5NjgJcLM8zw7cYnt+cZhVcsN9I9
/qcOmiEOMIRcRyzhx1NEag==
`protect END_PROTECTED
