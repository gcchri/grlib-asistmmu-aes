`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJO+YtQ7wXO+ngBnUUwicfoyF6XBw/rNOpPIG5KltazGm7NDVpwQ+zEnAUVo8cPi
J0AaNLwhbVsC/VZBNnFsFHJRfC0LGQ9uoBH3a8tuRgOAX/O5ta1pZqLe8lu3+wds
POInLSFTH+ufYnDbDMYvUBzgeH0SQ4arw7J/YBgcbG6+sXB2XbB+S+h7flkXPlqi
iFN6Iu9aLOpvRD2CZAiUw9BDBX1DgxnPJjhY9w6yyTGgcWCTzyi/jZn+yc2AGSwL
nm4ExUoKiBJCcmYiyblYsrmGwhs8pr1ewX78RbVPxy/dtIQpnov+mm8OJSSEtL4e
7iBp+GtvsseLaiIeI6wkVzizG3slIjUO9JzNz/ht8U5R4MRzsgTxGitE4UJjC0GZ
`protect END_PROTECTED
