`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kobi8DdSyYoJONon1zC9jJ3lz6gSCNeJv8UkHgAtZoq0cmU5cVsWIeYWzXBXIais
kXbfOXVDuRERP+Az9WXyVGe37KE0xRjGFyvLBY2nqGcH0pPHm1az7CfFJhyaKhC/
XopjxYER3RtdXPYFOPMVM1GHykShpdcSX/oPboP65kzFGKtQJUN2bOLbt9KUJrYk
W1CLQtM3n0QMn/mwuQzjaEDqEFthtTlSLb5u+ktOlWb9lyY/h+lbLrBUwL7tKdaz
lwH6XlUjPTsMbHsxk0Fxx1Pm+Kg/g631ckYExR/nta9Pi9fedMuR7JnChk50uU26
kgPTpd4X55MjIeIR8NbyUhwBCexz/8d9AmYhtTfJHsgCo1Xui1OXte9r293TSk1k
uesWRBx38CZDe9geM5McCcxmgmGddztLFSSOGVVg3h4dvGcIhnyJ+y2bHxA35jpF
sNbgmYJZ6CtA3vCf+bs9UWw89vjIEI17dxPY8NM4y0vUQceKE5xP2rZdHNAMkuUA
R0Dh3LSo3litetBRuQdPe+pLA6AgfDkq1q/Qp/6y1IL0ARZ5DD6J7qFcb5vK8CNK
cUkZ/glTT1s49rKcHq2dNGbacs7zqeu9VknEHka8ZRr8gnziSfevD+wMUPjg9uS3
FhGtHigFLoKcvLBmAd/uFw==
`protect END_PROTECTED
