`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uh1DD4Reee2TGqy4eLym0U0/9YJ3siPaYEFG1uhzouLxggrQ7d6l+dbvWaN0opBe
azZy1OgUM5z8STJUCc1f0IeWuzD/kQ/jqFX3IkZiqOQt1HTG3w3UsmdVwpg+ia2q
M5N1DyHg13X9f0y7ZI/Pz2ez3Y9QxRoqS8Z6mG3Ys6G0SbwQ70mKE3zsnNzbZAak
mm1h4R/DIzMdWDEG3boFfi5E4Y51AtLhzEJCta1zfuDGMVuDY6gPly9mmBnwrQUn
MVxNg3T0ExeJRJkQyW5+9Q==
`protect END_PROTECTED
