`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QdSKecYJTeLGyQlq52YOs0VykRRWNgHSyt+cgkkXIQuyf+jZSEO5WeikHfKqzV3H
A0thXpy4KMVLm7Ihcp6DEUXxFwi9453CVm2CakXXCQ2LR4BAG4OM48Nr5+4hichH
T4LSm7Z9PBzYmUdfBWJxTGH9NSqYyMg0ZHpEaAbJk/hUiTmPy9hMJNVMY6yKWRxN
eCXeujJOcGIgVb3dYK9I5wcuXxhbQfPpmw/yLBGqFaRsmEgAvvcT2pi6jRtBbl9S
DS/+ei0LeQJXmQxx6OhIhOr6guEdI2L3KcfzmCK+2jdxZqWYP0KB9qwi8QTRWbiV
hXHjoc23Y+2eLQ+A2guPHwJ+Try2vAHpehw1C85cHWssV+GI4iFMNA4o19rOxneP
ztqjzKoxxrzxCUtdma4aiw==
`protect END_PROTECTED
