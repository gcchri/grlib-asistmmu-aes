`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJK0w1ootYhoRIFv8mjvmhRWzH1dGglePyXHIOkAN+N+UJKVVC9vKoR8RPieqxAv
PF/sIUjW93GdrirmlY8Z9wBGsgl3V3r2PPLEEuz+btMyqJyr13xG84LMMjdqJKEq
yBHflsjI4QhNHHivN84Bwi0lKKthUv6AsYODMXME93pyjheuUf7Sne23InRghzYI
XrrGK/Bp0VsvOZQ0oqEpSAN4jgoQSS1YicEjBpjFx1fklWOWQc7xQyGkesQH+wED
oris9nwtLhlCOMRJfUDd2sHTjywJZLvWWYHnQA9c3ryJYoeD5XNHGMP7PzfPgrid
zV4jo1noPCEm7AevNvSc3KeJukYvFujXZlVnQXIw1ub7UZKgvCg50+ZfbHU6Py3A
5giu1/LfbstnB4Cud/kV5/uYRT9aw4qrgoN0VcCO+iAwak1T21R4A5uQZ+ab4xi1
fpQonZtG/T1SpqP1HI8KQ1J6cjbrRIv/rpLms1vZhpBnBetLxjruUSDEUwbf5sJG
Pu4UMgo2dLNNbJ1SJkC6XFtgeuCFiyvwuCuZy9R9IyHYMsedkXGFsLEP5hEgjkH0
w24/D0p18py7j6neyBXyX/VErrNv7U+8H+bNaXADq2qqjEvkkgipxhWo/fp8oIlf
UZSkek4s1CWjn7GoywWqXuhxSA9fwsow79dO74H+4ctgDC8wfkN2KDIxbQlU02Y1
Oro4VmZpu5SRuEnIAWSYEGxLgkuK+5JBMlgPeX2TIjF64vC3XTYsekALDU8r5jje
znJdp2D8UAcYQRmwqDEa9dG5SgJIsGm990q5+LsTtox8YxhiwMIFzb+KWaOYjVUf
Z6rNoD9zCCxg2/U0aivrT9VOZT+krfciYS1NBRfOIcuy14icK2+fQd6ZTIIQtSvB
yy5RbjCAtbIegjFuG4r5uKvkEW7IfJdTCyGvscIixdmTLbs+vtWnKC3dJuNRM0P3
`protect END_PROTECTED
