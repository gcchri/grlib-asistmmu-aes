`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+ZcUrn1WZq5aYm3V1tVN5KbKJc8731t8UzzaivQZUpvico9MfRqCLl8eRLYAzdg
k3FUFOOcu+njWyrtAVF3Kb+CETBb3IiDhIZRF21IO3C20KFk1Jlr6wai2AgIyspC
X6LCZAVlXpG2LdcUh4WhPrjD1RuXNW50FmLsaFdcSceJre9qDepS9+BlTZgfiw8K
/hXG9TJnT2N3JRrqKojsL3hJFFpkl+544RRkR5MVYtl0ZuVLunlRE0TCXzy/TDDw
0p0kPtg6vZcjE8a56OvVrV6Q7InofVj9wGfmU6PXoOTt+ugM0xM97JJlkJAp9rtg
fSv8dPb+GASKixNjB3TuSwmtDf7/KFItgkcAnN4uB8N7u//pI+nb0IEKzf9KgbE1
kCC9IdEAwAfm3yRRjGmXCHXOTPvvQo6Xn3PBTp/DbKWOkWPG1bNrcnPWJwPmg1hZ
eAnEcQRBvw44iuSBRd73Ic4Lgk05Il9RCuVvjJaRRzJY2uQqscI6Ihusr5Q0K9g7
1vGzoLhhxtVtdsmzEvYNU7MHjkIBMkXp72XUMDKY9Q6W9H3WGuQMWyuyf33If9qK
aEsMxr81HuAVkiLKQMKQciteLYp7/IKpEe+bZ77BXFeOWzE76J0k2ii1IfL7rzxK
3dBDbGZ4Bs4yS1X6EWbGYw==
`protect END_PROTECTED
