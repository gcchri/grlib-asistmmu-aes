`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4cf6vFDyyKuWa1RsWK94LYCF353a/vFtlByuJfk1/pTeuCginowTi0V0gBB95AI
Tu8PpaupCO//YjF3yizrKiZrx1dxH2jd2U+KoGY9twu6Y+efcrb//L+UMKWNeSnZ
wboH6pjuoDcFYbAl1hR2chDCKlPRcHER9an/vZbZoely0UYg3BrMn/eT4ImyrczN
DLkrXf5aO4urS5puLsTU7BDT8cBckfyMkAWhahFlqVe6f1sUkKrJesGk8Q0Vzut3
sA0OtcMvQwoMGyTuYqKckcs9CCdbRU+Mdh8RbIOzXbUc6eX6ui9P8DHvbGnFxWGp
L6zGVLmw+gNb+Wki6PblXhAzmP5cW/cnfimUB90TbwRYtE2ZM21/jT1f6mAcYQU6
uXCxz4G7KEnJ6NNn0jma7N2LU09XuY6vOWYfwCPiD0keYnGIxR9MvNL7f1/2OMVf
g4PBYjRooghua7ZgMFAip0BfMaIz1tap0S5ZtUxFiMflLduADr+f+58UKQ/o709F
9OmGLHbmPwqSaNZckMtl2R4eWSvxR6ODrWo7oK54IMChXde6LlTcLlnwQoM1Yjm8
nbN5fXW9caFVQr2w1ieSbxNGQrl7veVu2LuxcVbe1mCMzb57psTDTOLCsB+cOaF3
/yyl09rSnWSqAHYpDIO9dUTCuDZYKlBEQxYvDB++gUpqI+TJeIEti1PUPupFeSWd
H+OpsEuggxl/WD5sOR9zS0yaUc0AZVDp9TnXbaknzONmouuv6S3QW0M5myOF0Sur
d9UTDx9eYwUGV/ppB7KPIOtgLh6L4j804lEcDyuQIHLrI/TQUCzW5/FRvCdzEuUp
g/zkHrdWU8z4lgUwQ+abb81a4LUtix/aCB/vL9yoxh5eIuMUdH1sIiKsPrXj1Uh3
DAbeeQGsvdAuzqu092viylb5Cebxj//lqJpB+n+Dx17t177K+cjJMuoJcn6oKcDb
QpiQfvelNll6CrsO5bZ+kn6wnzL4yzIzi9lxS5crT/IujMOPl+Xv3kEcUDum3e9b
tZ1UmMj/BirLMbOC3NGp9A5lZCerBeEgs9mUHi9h+fCVo+ms9PuGiFS02yuprZOb
yE/8nCLyK7iqSrbH3MJcG+AnTGNXm3gFgZFlLTdtq34A/4aKV5OUyMv1Hb/5pXG9
vzJ/C+xZIGX1L6cA9CFlrPV8pybjIvPY4w0HcnxMyzG4ea0jekUyYu91gQ1NTNYd
Vghec+iVLf8KadmB9uXdEXajyD35SbjbwP8yCWabshum8c9fMJmbDROpYQcT03cJ
1bIPOmtOgcGgueq4fCNJam04kHLIPjwtwLdc6+ufyO6QskavYxHvn1qyWO3Hxz5v
dEkTzvhnkMkIyr+HsfuLmXKBcAYzJfy6zNlQzEbb7EYyb5AhuaGgEhS6sbTptdA6
G14yaCPZb0vcRbA9gGq0Wel+5cumP5XUMExrZ6U+Nu0i5L1jTBmZwhA87IcE3v/R
JRxh9EpNxegBGe/ecwXk1jiXxcwXI5yNTwo427XLvdCeWnbO+bK9692c/Twby6CR
HxftCuwFreGwH/mvrjJKCLALwtj8+b2QIlSI1HmxcTE2B83T5bGFyvbnC+WZ0nZL
AeQkLlCn89m6q1dB2b1rB4KP/TrP5HNJSjm34BmJTK8NSwJLi8sQhyB3RnJPrPBI
6Pk/q9hhjR/AW0wF/bmTlkbFqIl4u12uLWo7mL2eQ8uPeZcGhZsJDhCIwyth/9tD
h60mQCgxI1IHy1yDNQKk4KIG/SX/URsgGd1vPr3zPUXc/v+COQm4Stvi7rcnm9rI
5zLumhtfwk0cMfU1giDfBHV/3fz04Ke2C8C3Y4H3QywTsMaIDKuCYBPSUW80h7iI
FgNdo5SuYTuYMhu7tJri5PcLcIyceLZ2L2GO1ZXdy+6n9v20pyF2M19C3Hfyh98G
pbbFvvdjNBZ7BcuWk08Rr8/z1E9b4Of9gkjhqnCaN83X7KBd2ncSPzBfXSvN16FO
Ol/lmaMleqG76IfweYMSb7Y3POFVZ0Z4CqpGlabB1Z1Wut+tpzeuwqhRefenTf0q
7ws4bte6SXL2bzs4kndrAdECmsp3r1zo34w1myYVwx008hPwQQcOoSfXFO66S/BR
6yO7DsIEbPLoQe8KEGhLzQmJDPgccWV/EnKCKSXlfhClIYrKd4kVG0FLHClnjYsF
vcotEL6YRN6NDHeVaPOgtri+h+h8GGOvLULgs2FdpvdJ4EyYiO/qkdEpcoZAme8/
JZTBpJYaOcBJoe9kGDY84yhtutQx2D5ybDIF1WqbTmBeeb/0547Y4ySxjCQFA6Zu
L1IgIRMQLdmwhGIoeTNK3Tg3b3XQ7LR6nXIm2QZrcU+7KaacfyfTGE2vKara+Jk2
CUJ3FC9924JEHgMZoV+/ALmDnlAxwxi+NiGoGqUugy7tBekICc9lWKTkWREv1/NS
VYPTAIUGN7xr5ydIdSTcT/16Y51DMErWXZl5Kfs26T2MFEjvpCpaMPLQ+/+uvKGU
MWt8EIv6qxlBx/hfV8j/uyVSe1OBE/X/vrEiFEa61Dyt3eVtdjxgLjkfxhFjcvK8
cusQc5Oe8OttpEfw0rbAv7Ji/uxSlBtCfxG+cZT/oVSlxI6jMUv2A2UsJ8SyjZjY
+hxEMlTHnHoLUmcGiRlYNPdXx6QJTsMg7XJTVyuL5YabMLO05ueLQLZlz7xYgVGE
pR8mBK61SDz3Y2+/Naj4yraW5BX0asQpsCOzWHBOdIJqsvIwFdKGVpETLS4nT8S7
75Lq7pyCfHr6KuiIrHR1dXq5vshKukqOezYmS1VZAiqAuYZa2KSiPrvmRm0lizwL
glx9mRHH2H+31EINeX8Pl1hjNrwY3FB9iZKwo322/CmskQWFJ3I9qULrxiwyfSA7
bgGFn6CR0Y3LDCkeDbyaJnBfiJ6LPXFgIf97RkuZM6drDcuAPeklYy7SRI3IUTmY
PBv7gKcFHwy+bWtkkza5jaNjyyiWRm+zXc3ChenOcpHXcspjjJvyQLUoOaPm8Btq
n3RIM9ChnWd+sxgBDNGe8uzCywWGExlQRiTaKySDYh4=
`protect END_PROTECTED
