`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UcL0GMBRPHIIfxfBy+JtzbrZ9RZY/Zsh2Z6OyKxiF8UlQ/ADku+EMKuH/5l4Uy94
fE4FVFYqyh1hSoSRz2+zDwhiTiK+XU7xbc70FJJ+WCg4yDyjQB+Auzcqv4Y1VTuk
lUqff5Xtz5TjIPxnXj3ah74jiENosGupFa4uKpllpCE2gJoNn2jJXgdfS+HhcSIP
+D+Q6X/vWuvd5rQm3Poq1bq3HXdlZX4mcr/PD5f8aAyMF0sSaSLbiQ1aJg44TJ2U
p/eBiS/5ZuU6RH86Egy0Cw==
`protect END_PROTECTED
