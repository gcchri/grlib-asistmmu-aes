`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VxL6+l9beYWDk5rnza+jNTIf+jQeSUhxi8MycJvrORAg70mxJ7rNs4zxR3HxRXfZ
MqExC1x67W98lsuXyBZqVP+GfQ3Z8hDRBRZQo/1pG+iS0MVcocpIqLBMSjpeTuPv
AL/mTUGMevTAQTcJ86U6CXyz/SVrKBLSaQTjvXEF/+aeLu10ROkr+JEn9UKsOsPv
NUMzEkjS3vBys0il9xJgqxmzgzCpM7lhAfUnAH5FWEiHv3SNcxkvyUP7yh5EP2I6
k0E+cfAY6kJJs0g4S688ZbmFN71R66bwEslsqBAo+8Z0gneulxEDE/cLFPHG2R9D
8FP0slKkruc/aVAk1pbcYdF8nw+cTqlu+a2kPu11+T8YY/f2JV8eKHDixNnU0Gdc
1yVOOIm398yDK7/sznWJhsMKTpoQmqvt+bfloVQoDp7xRd2ll4l4yiaDBSdzZjU3
1fGdWXpCvohCJRqpO9hiw5XsSC8UoJB2FoXrugDcrAiJlGK9kuaS2Izw69CJLtbe
9JCUkShUOEYKvAHitqDLMnNVF464DWWTYXpHJEzOTf/jXKkXDD88hdNDRoBUSMQk
3sp8L4OpdY2ssNNdTWb/voWtOpsL3slG9A+xaUKS58zOVb5b8Y7zajiH3NlR9fiK
9EFrkQQQlGwJrM3m52AFtA==
`protect END_PROTECTED
