`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5I6C95npLgSdW6/yjYGbGC6Kzowkcu4cIIz/dfb5URjH/nnhfnBYnTXnZHnlulXV
/qa+h1u9ZSy2R3gAdPVkXXeC8Ryy7F0YERwH34qpZ9EPpcAwTQrOTmwxHhdPfile
p5BnCiXq0Ii0kCb99mLrSrsbL3Yifcb2NaSUGiKEwOE3JFnofZDyBuMztnTPWUrB
lIy0aRDkL66zpjSPxWuEFHgdlqwBJ5y5IzeFdPB8ObYfsVrT86uLU4yZz2xcmnxe
CywGVI+l1RV2K6qmkKfGZQ==
`protect END_PROTECTED
