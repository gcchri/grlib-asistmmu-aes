`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMps0LOlw/28ntM/TxXCfhdj/kYeZM+wzd4AtEWBUQAngX+FJqwt1GvG2C6+grAh
y8Pdrlj01S8j3w5tfX3IwCPSc0mZLcEfCSVybVLZ9KJlLLNkoqZxxYO0TYIKaQoq
sDe0H12ZoBFeiTJ9wMBCRll4LjEyPGcaHPE7HJ6nZ4qSq7IfKSuOHE4vFp/JBz/y
A1D6nC3PGJkQK9PwDQ3TMzJah0/XsO8j39UBI1rAjxjMguZ2xjEaI455tml5iH4C
ueTzbufjbPSfz+t13soHaYPx0kKbYQHxQGPmQyFtXZ9XFfvR+YlnZkz/y11TAJgK
tI4QUgJCKmuI/rEBcFVC5MtFmXzm7EdYAun57dfCM9S782X5XNWWWPhaY4RDHH9J
dXWAzNL82/DnemJm+PJm0PBnBGoDj7l8dbCDSKbXIXx7yU6puUcjP0HZvmTUD9YU
n0Z1x+teZZPyELfcJa0kIOq4rJEYufN67AkhUVvbPDmZoE/LMJMY3yM0Ks+mhE6E
5DYq2C6SjPAgxvONYVUMDKN+Gi1/nYQXfsrv+GjQ3fX4+PXyzN9PYhCxRqfFZMJE
ll+v/qpi61N5MlOTPh6/fmphGKKhYAI1I3B1qoR7NNHAvBYIjRmiN/YdlnLfKX3N
rm5bulKwkpdorR4lZUdBxKIurL4h2x9eFUtw+PNOUh0ISqbz72JgTZOj+aWlswX6
5bqQBTFva4CeQF6qoKX3LPh45sgdYRVSeF+CylwJH+rCJ5t72jFSfUlxdJXyxoeV
zi5bG50029e0PMwLYx1BxJZsyEJM3P9W930yvp+uEJ5KUuHvHqbGKC1pI0WyUDDl
SAf88pSvCjGopJZrZ6LJTBhKhATPjaA2SBpR7I1Oo9uKnHhtWvRqaLSdbS67gRaF
rIxpxDQj9mCY+fEr/sEqxVJ+RCbc5x+5vuC/GkXfXKUOHbjda9zaLAHys9/eVzO/
ihB2O+UWMnb1u7fVhc9zopuTK5QtcEwRe/AnkGV3M/PXrXP+RMElRJ8opDSUu/HI
BLpEYvpW2awPxgZQBfVcBDJ5RTnB8doJSH8AwGUkPfiBNQxhc6hDx0wLXCdbB8sL
kM5T+NyEw5HgRPXsnDdG0txMqEKw2nyROs3Dn1kLr48jylNGcWiNy5CGlVPlCCul
/4eXZXUaS3W0uhi7h9XPYlJX5g0sBxsDZWsDZbwJI0jmYXFMm/zPHRQDIMrUd0K7
/t+ouKKR4rR1B/FU4+SBuobIKwSn0M8LR4yr7qo0IgDurRaEPK78dgVmNmTKA/Zu
UzF27n1+epQ/IDXzYfcS9oCAb8NRHswIHYHBb8QQldeP7syprC4nnc1qI5E0vtxh
yXQ8E5WXcD5vGrUCtC/eJO5N/lNMKFgxt2WhcuFuoOoxmM43K7uAY8EUGZ5Vr945
c6Rfl5/OKHVO9R5D6d5xnsYitAJ0AfVZd0rJ67Bj4w2iJZtXSV+RYCstsx3h7F7G
F37aEfUMZSQxnh3mJsoAuqFK6RU2tzIqk6/ZxslvZyReXAXaztkkMWKd47eCgMfp
64WLrkLwO1MYeKyEIuYNWd2fsYibtwEe1XvYhw2ogxYmbPj0ERR37jQlkWCOxQVe
1oW0i2BLFp/95CzqAnS73v56smMv/LA7jHSIBhznjqIVIO0lSzHJpvDnhZgBjpxe
t+sweReH4TfVjjVlTQNhWyZ7eMSqUzY/umcITXwl6kI+BdtTKWu4RpRQpKtax5T3
lXGeTFtZCecELlXKEK3VJZvubfSyKbZqExEzF5s/nshVuS1QOEW1ogx3OLkjSo4q
gkVOHBX6VcZEuwDs4eV4xVIdXadEgRSl7FgLeGqPWdapI1yT9Kd0KUTCEjDI8pnH
xV/CZx0NohJThuuxWjJfD1cOjdWGv2Bj17nwZzGpUAqYjGQwuRpTImT7UAv6I7e1
vgnnPXKsjJySJ4RcgGTflpZrnIBvHeDj0Wud3e4O1zciBw2Z1Y1mq4xTMy63kdeU
M2Zb6hq1LwQ1KtN2iNHsldLItwIBSkcKOesAsdpYp31IBE5KHuf4Lyu8s5E1RfZn
nKTv8AplFEM6WztzZ4k2Aw==
`protect END_PROTECTED
