`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/1jlRBUU1yqFv4aum+6f/7MgXm7fql1Ig0D0QyervlOoQ2cwhB2ysUwgm19Fe0d
5b/aXBsYxAaAfob/Z7GagcY/k7QLTDbAZtT7Gg732U8YXChA4BKI6BpYHmpqM0YH
z/4WhMSwdwhsh2NmdScvpni6OURNX3dXruYpcunDqYex0wpqJPzZsPhXsYRCy3K9
iOWok4pNnGXr2i1xuWUdOjJ5z/m8Ri0L+ACQjZeXKSXs7AzRAa0+aqPbFxCEib9f
Z68w8FP8bQ4luLAccYfDqI7byJRQW8xNW9cqkjCgDmHK+bEFVrVYqOFbKLKnY3pG
mnqjvSwDNcFDGLgsVVa+Xd8mp5AK8DF7tO/p8NWHARZurx/JhwsXmFyuoGEQHwZ/
`protect END_PROTECTED
