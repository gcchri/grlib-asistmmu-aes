`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F7a7UrPnXRIDgbhZficorZ/wI7cY48DHTsK+wnbMtYevLZgLhF8h5ya5WACuDHnZ
vClZVe1vAEFggl0lzo5+u5TWoVc1r60TgQA6WM/FLqOtXnRRkt2c/Veq4juvPhG6
q5R8B91C9DoWR+HegzNN2qEmGGYyXq+9dZ9pghu2tla8mcoK9ufnZiauxn7NxP+z
+56zqIrT5KUfHZGwdAK8q+IPVU8RX2kTTWxmY93QY4tRkIGbp82YukH7xmNckZLp
6YpvFgK67+C12e8nVIg4MzP5LJb8Dn/8CqAY8lXOi86RVuAc8mhuskkA/C8NEWzJ
o211X0tFR1V3T+LlDqmpDA==
`protect END_PROTECTED
