`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t58GynpAARbCn69rVkN/cdteZ/wZlp03b5qvWWuazZgnWkHo+wSv9YHerM9OM7t6
JNMITlm+Hzga/r/cyeOwKus0OPK/rtyV3KezY/cDeK7I/fPzDrLRsRN1dLrAuxRl
MMjLNLPfTXESKELg/uPRajT722JGjUSSzWW9njuVul9q4//4Y6kAZ91x11F8GM4M
La5z7/nMCpKTH7NyCPoSvhm13tqndSjwtqhyUywC8ni2LbXiOVvx85ausdqDJGLm
NHrezgknAvTyVeJziaqKjsxuFS1W2YPIkPqpsb7Jtztll97uM8/aEN65OSFpoKux
VZGnG4b7rpvLwaQtioRqiGi4NkBGP0X0u1LdQpF+GBGoLM50PYgePE/SHZbDKib3
CDLJDWDtGt/NU9SU15v5QIxCMeEjH2z81gxMR8H5WXXuQKlZisVA0ZS0Gsn1Tyq/
AD+BlNwGtCLRSs0jrZSluwGRDzsnAXJknZBfxRBBozLDCKyxvcmnsA2b5i1ROC4c
qwLBG/I72KagrFzzNuSnr4tVteWSyanuDA/Cm02YoJ8aAe51WoWqbZ4GqxgLiyx1
fYOqyqhlc28Tgm2FFqHbHTPqwMvdfhwIVUK59+IpukLjbQLKRd0+finJV9YR1fOy
3xY1fid13cSmzFjmyLjMecbusgqnOopkqzK3ovWDXlwpA2hoB0DwkaBWECI6jDgk
tL5EkGXvkXzonO0X0AkRupVCqM/LDmxfAJYLS4xTgWlPmml8UJNl3F+cFqomznA+
`protect END_PROTECTED
