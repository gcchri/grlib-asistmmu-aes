`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8tTLqXiMg7vLqTzHAbyhaubvajbcfJ0nitiYeOAh7V7Tq5Fs14ux/aiXiY/tYNDt
ME43UgjR57N6Cs5blLoR4izkbY2+8Vw26CfoEVdNQDsqRNk3jB48gmjmbT0m1bD6
RVdwupod1eVv5bm+ro7B3a829Oy3Z2FbKPkVQrQjv81GWCPMPVgpUIxrIBcSa77u
HqJMXV2+jREU7VBT2FyPiTYFDhM+Y0baAMeXBRozoZ+ZBy20tJCEgXo4C/42MvkW
R6aNDZPl/ZzJ+cdsKKhKBxT7xFd6korDdSCgSjd86MjFYBTyNbPUvIkbTWeKZFg6
cv0Dgn2Bgr/vSIsyX8QnouuxljK5XXNak7ryPYYAWf1XNQaGk9GraLs4my/cU7M7
67t9WO2+8hRd9/J247l8fStuu+JsqLfBvUyc49X4q+aPvZ+5o/Jybq2Z9Z3RAAH7
1wQDhABOtQJdP4bTLd2xVt9MeoKvmGMoDi65KmX3yFK88mzbJDm89ZkTItO1xMS0
Q06Eful8DLZJPmYObYEEuzuBnFKo4CHg7HRs7I6Evb1z+xN+qLG6lcQ0pDX43Gbf
lAuZPjtu23lBTglDYLbDQL/CHrOcifczmt5dn/ChBsnokIYCPD67Gj46iuv9aQEh
OaEi8zhw/KyUPTdCxbSRBqC+ZcRpQ59PmxzTcAFWo1A=
`protect END_PROTECTED
