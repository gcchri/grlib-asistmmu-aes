`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wRObs9lo1wFu+H5/W9XE3dbUM1HRwKp8MvU6YBkf7cawmz1URtoHEMJ6zswQU32d
hCnop2O5B1551YT1C895uWqercyCrs7iCWp+NjyWQ4ucOQrOFQ135znw7G6HH32S
6ELPERDh6l/XmssUm8J63sM8X/6aZNBPXUQf9FVODqaRdmYpCtq/txpFY8NhgS/H
Y4aur2A0uTGZmTwMPEdoxdDgAn1Tb9R7A+bjWXbB8yWVmacPrhXqiYepTt80DwVJ
EhPnbbA8pnH/pDzoan2V0HyEDuu0jsW/JmgYXLtOX1T2nI2mwRiJ0sBsv9NVT/7D
GUZza2MyBCnYtJz8guAnewTzPrvXPzUt1XVR9cQXtzIN5jtus8HSNkSxhSzQym+U
4ZZuf7W3QWiPGWDe9evWvMsLFxu1iBO56expPb1u67NehZ0Gp8XdOEtIHfbmKBMq
LQ9AjDyPt2NyuBdRnkB3SkaqH9BGgC4BtanG15N9DIHrCppCJtJX250JXQH+ZpEU
LNzDTqhTaMZtnE+QEG/F1rcXKCiW5SavHeZRNxiVj7s49tYgUrrLoODASds9699I
QOB+XmLFsRavj7e9Jg92DQ6E8rNtvlkyzZH6MpINI6w6faO3pMOjFB6g7/2wYh8U
sVduF5dS1kn+iw3FIlBwgFTTCDYWRk4rV80VfzKRPE+Cr9Pys1fTaa+81o7VxmcU
WV80yveONxQDx0i1tEPob95rG2xPfum0iNkyfEE6YD/PJObom1eUgeET97OwknEg
JjnSTm1qMFmEKanA6PnpM06LUErYKgtorMGXyUKvHNFPYwpEQ7Hb7g05eH6XDBfb
IPmEqCkId0irSXYFVC34VmFnXP12KIw56EBGlWaWYWp+CFl/j6PB4e7LoT30ee5P
nS7jcBE7LFaZPGfl1mYmzsn3Kww8L/Z8RzhDwLXq6iI+Dd0iVtyTpLhgz6Gf5UZb
Ne6EhV/T7dae6g4hJG4UGzVc5X+2UupJAeQONo+KwNLINwV0ix5K45vyRgB0VBxj
+Z0sQX/guezjEvPq95hvwFAKZBu2KKj7NbFi+qYWwqN+P0ihqKf0p1VZRr88VX6H
ne6YFoPEVvGHNIo+eFvn8I3OEj/VBaPTVdkbBb9VpXeoQ5X5J2hIzLWcgOVUezpv
w9Uz0utxjFQ6YUTaTrVEvDZInzfeBdsfPLIdYjDVRoFSw62kKjcRQmdr5gy2ZW1e
6LktOiA/uok86gnywWFwGF/9BXcOyQ8tdf+nfrnLBNJKdkm1JpFcd9JhJ+SZRYMD
/eqy4/auHoC4L1zfNLN3/cg3lpCqt8ErSw/gCOiulLDD9mIi7QypeAtvSFU3+wpQ
IV2rHwvmxIaRnerj1w1dYSdtNHLSZRp71RByndUvRvazyK2OO7o/GPFzAqZHI/Ox
`protect END_PROTECTED
