`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JnzLelX8ROUJ9DLl4iGr3hZ2IUY5Na/7Vs/NCPzZ8nr9so9BZYpS9XHnS6/78cz0
tnjVtHL9+jVd/Bcens+T2h/O7UZC9oWZUiMoAN0czl/LqWaa5d+Nl5NXmhwsg7WG
4UshX7rDB90bLCSsj6FwhX6XRVCyB64+QbNqMw95guciGmtRjOcFmWiUNBzjl5GF
pal1GCMMRA0e6eaW8hIUUH7Dhgmu4VGcV+qW7zKHdvRowHuRAInPJjuyRmlKwYVl
MX2WH+gC+AQBkP6Cmh5aa0bJgZKXYkXiai0CbcmCl79ibMpI/b06GnEZpZSBoXXr
rZbglw10MDa50rySu8S7GTBkCwkquSNWKUbEJ6Vk2yCNnoTD5///hFHIsicmTaRl
LpQdTWDowN18f0NHhgX4he2ICFWvN0vR5ArecZ9hly4Eo9Wkp/d/Fr3H+oJDBh8i
g56Ve/JJnf0WOPgMcfdGZooi2rtSjFytYUuM04JPoPF9z+n2v9QGdwC/AskiDugg
Xq/8fUgCb54CtpD6kxvi9fjcJC2tm42XSENVSSUVTMJKaFVTX42lGw4s5l1cTdG8
Tgsc13YR31KO5Led5NTAoVRC8EC581Z7jCtkeBxk5PbM05IjeguEt4Vm48YXw+xf
tezwxgzNCZc1EGbVgLhfbw6/MiibLE34mp0CMKSHD37AMfWyoLpsoN7s278GKVqP
dxMoMYaLRbh375AT8aMJPRG9tq5NRExd4zv7WA2D8PPo/wDcXNsOUx2GHdUaZdGZ
fl39vlBLrNXkwdgb+xHgcjU//oFpAFJIZORK7bokORpQW/EQk5fVIGPkJGiLklU+
tgM+QMsqIn47ALS4Q9vYgqC0g7HlY8vmzha79OiZqVRT0ZLH1aNfhUQzRyyaekyo
iYPK3lKcl6KFtDJDQt4w9sDEopBwVJ86CGEb5fp3d2I5ZhimHYaJMpc9hlIS8hwq
E5UxWs+4q/0E40q/CWpJkOgvXQ0rK2lvRKREzPRRdot5rRrvT4Rp0P7xD/m7KX71
BICvisDpmdK0SG+oKUUrvZnwyCTMDkcbMN3R/O0meQKnYKK7Xj4XjceJ2AKsCXKP
lzRhczmGkyHEaRl2v+p87kI9K0j1h84JO1jOV2B+mLcC/BZUmZyfcSEORb5xfndW
Df5bInbP/YSf3biqJLwvK6TSkmroLPeWf2cunHUctSSvhqyUamEsUTApB1zcVYxP
kUfi1AcvYSdQusx9nPN2+cebNC5Du6xaI6HIxyOo1gjE7KJfF7e8wajr1UFO2CNO
99Kmdx3LLJJWkt2FCnAgQIPvj8Wxte0+ib4D5FAcCw5d7SQ3EJ2TXpyf8lkaff03
hm75kE6TMsxoLfa+9twrrM1xOtaH1dsLAhgQcxOshUQdv3dIe6GJiByrhC9SKqlC
lpsO7avwXz6sAbgUuqzPmbGAyXQumVxQvT3CpWsPBmTAalx2MORASUBr9vzfuSCx
NgP3bMHoNAM50XrnNGfyOot0ZCuF/6iHCwNlk6a6m7uKra4hlHgF+jaq6TtXDxEE
avFJ0GoggV1n2NxJ57dr1F4tiTNyjPisJuLMUZdcj+7lqFyCoSffvwLRFT9CuZEP
lUQYqHOnOW+UePX7BFEbTtN8ylBhFbHjsreVpC2PKiqkEZ4LXRwUlUzoVIOun8KR
qyhjkAt3Jl5PVyTuZU142TzIFBaiaifdNqLYY0QMNcHgBbe6WgHcglSo7cug8A1J
5ubH6OW5TfDwoJRPaKMv6BnuJion8omPAWWPNXdW5bIu4Afumh9qW52yFpF6EhDz
shY9I7CXcXD66kLvouS1pHClWxeQGz9SZM1OIQAw5FYu9K+330ttkPtG6u2dT6VA
xgQKKLlvKuEh8+rltsP2pHpqtWZvWWNjb7CWsLfF6c6BGSx9sYZfTsfg4LSlE7Qt
KxxJbe/ecsBut76Kqn5ADnrm/N1xDz/NtdupPmi3J1Ryzptu8HsIEr2FV16YZprO
`protect END_PROTECTED
