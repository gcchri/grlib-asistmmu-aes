`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BjGlwDuJXpTWtmOhQVUkelaOHKD4H5nr8B7jn8ePtW++wKdUmzZ6h3KULb3Abz2q
8Uq7FqxmLY6Eet9lOwy1Zd9bGtwEzhvCrcDAevaO11WLLmH54qeTaIzzcDgYtb5X
3OxBcLRKKUY4TjgTIkA0F/Ou2FUSMel2M0sLRr1eKT5XTVnU9/Zj6RQoZVUYQLfE
8Jmo3APWrV2Eza1Lgn9v1pxPvih+BsAQX5bhwAoHLzfE11R9VRtSc9hpgDdcXxwS
FQoPpnUvxljETk0nFQK8fHH9MyHiH3GWoObOiBAGk67mHpi/8goLeLyKW90BhWjq
P//ryE8tdKrqCPTQxg1PdF/ax5HBXSulZXFdzF/c21kLxQNPgj9oSbCk/uvOJzEv
+s8B7/l8k3Oef++NiBPluXA9+Vzox2Hu3iSZUyQaCIH+kho1yscoIFVnjysdSUxd
RZ8LtF0jWNnN1/SA4aVDfwS7GsVSyc5JI44Esbua/PEL7Gz64cXevstgbbfJdRD9
c/1nKYKP9QxkFBGq4xAcVbeoj1XZopRrsVnEqi7PUAk=
`protect END_PROTECTED
