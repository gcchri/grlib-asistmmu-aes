`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VvdBfdzNDoCXE9Ugs2Q0lFbG9msberDbiz4C3y3NqX1U/jVg8DP96lvgzixVST+m
/flViw0+rj+YyIM/9JJTW/pFVbkfxcr2RgL2GyxAU5LgP3KQE2fRho/2uzT6O6Ie
8M5KCV5JA0eChnollxw9A2jXASk6IleGkg3dtP5EEI6gkhUzyUkhhISjzybcJPbm
c9twQQUkqhEcP075lE0GsepqKnZIEDVZ4fwWj+Ls/LOzTza7jhtCxt4Fioo386Yr
A1Dh2TDB+AxR0CHqVatRQ54o/8zFSVChd3cBjoJBCIMmUe/JbgUEVQDxKetw/6Hb
Plo+EXSULrkCAvITrFo4fGaZMAykKoo+af8RfO3+W3oKAYVhU0MGN08Ne4k/ruvr
xxyUYFbXbeNW/5aUsySi+FdJIi6Berm9ktqqaBtonW+E7mnNb7MmOjTIedCbyrHn
aJPdm8oqhY5At8+OgDOURo9xhfIxy3wlYW6Lc2XY0SazMKvDuw2JV4XSGfWNKxwY
CwojRacfz83sgDERWg1DpP8+RNfW3Xo/EYO8Kj+TeE6jnD0pKBWT9Qb89HISyL8s
b8MY0Gf4safgS6ceZdEsBlMs2jZ2TyYllRrda50iSXQ=
`protect END_PROTECTED
