`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRCZbzECkUjXT6b8MO2bE5uQDXRBfDo3uE1ls2yi11xTX28WxK9IkjOl8dfZWk0B
guokCIHpWoIBPcUBVlJog+830V5YHxIm6G07jY/dvSPxLBOpAqmHIwXkwlLAEGa2
wPYMnznHMBBAxFBCgrvW6NET8bapSdOA3eHt01UsniW/qBwDNoO6MHh8rub/on7q
gMWetQb65aQ7Y+ZkyWWQ9mxl9s0qTnjv217HtDgQ1y0SxMeAzK+sKMWHp8Ue11Y6
GPcrykE59UgToxU9+xQvubrHHEJgvGsCuTWm9etyb3sGzWaZsJ63BFgMWZWM3kCC
tpMSkekzdMLiNrNEEcHOAIM2m9D3X2sjcJxh5vK/Jo76NJ3JrwTyVwzwCg0qM4eg
nipvmp65IZknKaWh18w7aNoS3lshu6DQ7V6Uy2vqCwiWKpdoAiPuIMEu8f0tyfiO
KpsZUYeJwRGBsQE3PbiMsmn5xzsb80Akl45zrdxE0/7abyWBbSkOS4iMK2zPLVrJ
AWMyx7Igwxd1bHfd7T2XFZtYyFnBgIlkgqhCawKSUHp9jZ+sPchcXgwDv6N3tYD2
`protect END_PROTECTED
