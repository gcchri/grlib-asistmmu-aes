`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Wega/OmXnijyXqbJXRENagndc8qxsaWOE94IKu5jwtcviXEcxp9aAAMiYuOKHRJ
k2Mdf6aLCuCHLUgMFj3UZxHU41JZCcYt92GL1VV46OL60CDcXnbnGb20vY9R4NGK
2Erq6w93yBwXDIRFToyLbKrGc4xGGdeQ1z08g5F1+jc2HDlt0GeV951Bs8Z9SfuT
PTIcyoaHyToh7yxtPsVo33Lb4RlolPHL9TRLdpOkojIWQT61iv8kMQzuRPOt2uKy
fY8L6BdKP+wZ03lFGBYb6K5ZAsY88Sb+xrep7UNf24toUpRtaqPznFgxuGqid3NJ
HlKFWBMVQr6osExm6J7w8C108XTPqUWe2wwxpvW/4VVr6ixgJI4zm+OmaqlVr08K
lV8+a4OOJYnsZUMYaezqFbSW0LXdIqI4XDD8ub7PG2EXFm9GWxQNsIgrkCPh6MfL
D0JAL6YkBj2+O/sMy55Ca3SzFkANgAJhYP8pDRyiEoCDrwVgtkP+RCgXe6w5CXIJ
`protect END_PROTECTED
