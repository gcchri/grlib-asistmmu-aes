`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbpN0Tc6T01O8oBcE/b0xW/e2Mg54w/SQO7AIIFcfOP1HmDfH2Sv3f4DmlsILiX/
nu9jTblZ9EOuw4SLRLnWSD78sBUk6fUUifqbgPzIKGqTW9452Q7hp16GbM4Afu+p
1qxaMNYqfc6MCZ/YqZoiV29S6/KgsmtlbxYyQNJUu0nwwB7zctGJufN6WKsD30Ct
TKgrPu9ORYM5IMCCU10SAtyHdR57nOntsLhsLurJ6I4sJ6kx4ERtjX6H0G9rYaRv
7igVRa+BBJ7q8AFF13iH0Yx3mFp00VwTDQL+9PY87URQUVDwA7tdw9DAXFc0HkJs
2wU22bbgOKF8T4KDSUFNBeSVmsJ3HXmAhv2h2yEroSYHeGMEox1tdjAgF6OhEeg9
sRtYEz7Fc6XBH00erUszaw==
`protect END_PROTECTED
