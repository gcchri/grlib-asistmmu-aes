`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Otq0sEyXZKVQrEnywx2f+6Qbm6zY6HhaZiewYInIPGsJAlu2w1ghIGxBvGfNjEPC
hmvOxALSszqCRhBA7d09qu1wcU1gSPXMSop7Hvq9S9GyP15hYVf/n5KlUSgRoDPw
1EK/aQtSiAXzX/rVl8Roq/fzzIfqcGpdQCnEQG6YrKcBsVOmRUVeHyWiSVAWGOMD
WbxVAHnQoigWf9mDAwvjcrQsB8LI3zMCIndRs5ponAJnwy2swbuvqHlQNqCmJQmo
36KnR4RLCabTmjE6RpLbo/8dky8cVSsmjnUs3xdyLU/Gss/26zow93VY8ncdFeC2
J7OZi5kI77+259HLhbkOJHO4OWYspCrr4XqD5+kDlH9qfhnKI/BP9euLXqL8kmft
K0iV1UxQHBhdkclE1MwkMg==
`protect END_PROTECTED
