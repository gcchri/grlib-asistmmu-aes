`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TME28R+teRP4wfeW9opkwdrQ1TDb6WeKo23Rt3Jmt9cYkOzpXOY4mqD0G3Ij4hXh
Hdy4goVEDKN2Hm1pvb71w6V6XRbtmEbQlAeSksFKM3FeTaVi2b8xXOyT25XnVEmo
F9boFjvbvDXnJiwxn3n3yk0E0mvk99MWJPEdMHFK/NKyLOrdoTQ3qbBOhvrdibtm
Nh3zPj1mcF9hjyxm18Nbitzt6B0hmD7y31xUHjb+vTmv9ClaeN2d7REmT3jxLx7w
y37jdRtclGLYLox0i3/CXbHvPk6988u21eZrOQgqDNo8GdLTINNRKyCJ+NNHlpf6
qy5lJVUQl8CM5w83hDdjEhOnJTvoybMjs9I0e0XvDq22v8FAw73QVBHD9Ama6kPS
fOd6GC74+rQjqxIDg+T/SO7KykoexcG3RiR+u5TMiDJAvhZrLOwxS/Zlv/Ch2ezb
3Ubh13FksPza0X6DAm+SGonw2nV/giMmAzudxnFWzY1wRN/TLYqFU8OtV9j87Fen
zyg5sEp1jRcuurETrKSxGyK4a3hMw9u1d3DKRVoW7IBc2249uwsN5EhckZckGRyz
5BF3CULloufnny0Uouttmg8TT96Y4HKTCWyt4tlh169dpiynOVfME7fEs6bcCNGg
3URTfjJblkVK+ufm6SGH8Vos9QAU5ysNByv9NhVZgB6S9em8UfNmY1uMGH2to2eS
9BYJsew/P8pmHyHnn+pieFFE+FnYFgS2eoQoYs5iH8vkXbNB+2pl2kg/t/A4ZDGD
0JvDd3xboljJbai+CejUmEj/bKqG0sJyqj3cQxt5fRaVFPOHbqnUXXiSsezNlcpl
d+mavlEyYZk+mMEoy0W305/Rj5Owl3SfQDlfenQX55ePvRO69uKXc+0zyAPIKe8/
AJXOr5GJynFNBsKfxCHJpw==
`protect END_PROTECTED
