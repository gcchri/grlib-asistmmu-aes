`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WLZ8lHo9BGXAIzJA7OxJgLOnTwWGOjN174tvBTuyMfM0hDhmTBsf43K3Dpq2D6Lb
bpyFAgJQIR/vwJzFup3vWHQbUz3OcCJUCIye8uyZOcq1JiThresdUhJPiCWLtqGq
071kkWK7D+zM9oxa0N5Po4Wz7RQ0JuiSR8+A384i7sBLtLwfmOeLBEgsZ2qZLvX+
SS4kYJIUtIeMW/VNh5kbBLjheuxid2cULuR63eCMLASNLu93driTYmfo9RpWX5Ik
MEmTuEv+vbWthGNv2pt9Z+SR/q8eRNEkKnloxgsDFzBAjg8AT3rU4JjffbmulMMD
2AD6DLQgG4GiPh2e7d2hVxyJgsqo1DIgrdeYRmQY0PU55b3Eal1FfYvA3vDsylib
+e4O9CehZuJYY0Vq48OqRZ60SLQT3K2AQOX8nobmRZjkie4j5kQZYgLBYeH41OO/
o5CXEBgsqEYvhbc1dGnkwSGqiz2Pd2iPcX9z3qLzrZhvEmAR8Kly7HI+OYqAis+V
kn6+vFWaraF7aJfeaNShEiHxXErNwuIOonqg2UuY83TniF/D1jvP7KeHrWCx2aWU
9xBC8HaUzMtBtonwJBa5+lBRUD+7bwt1Rm3R0Dd1FbUtuebYNk9oYy4NVC1UJRIO
zZ6Ios98qW58S1QCbmYNQIXaTeuzfT5I38a6vNTGpXaetdVzhd891/IGB2soht89
vqvCul6UtciLlLMGol5s/Hi+UnEtMoNK4fU0SwQVDx4Kj2+5s/KpyOTWOuyzKzob
ESM3+uHll9usD0UBG2cvci1aGqAAC6OLrEj6bZAYkra/m0+JsnI+IZewkW59C0US
Av4ygDmUn7Frd7VAlWDfoMmMAe3y4BHyc3cHi7SDDB3lupFAC+bwVTyqeVE3nDVx
NVcsj5GDwkN0cnyluXeprRuOe+hyp2ikCr4RueCCgDkBZQPxkmUffeq18MMAal9X
`protect END_PROTECTED
