`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1UGPamqKGTinurOpGluH/GvoNXkyTB6uMe/iSsBhrtvKL+xqBDa34sGNE5xPuI7I
LLi5Rui5Q5s0ukQFVYVvC1EmCB5Dy/gGM4cYWaJUq9EQzv4iZ8ML3yvmkRWD5KOG
VzgrWUpFtUXWD7QhIAgHYWz4xuC5ktHXAu5XNW2ldw4Co5p1MDF69bjexn+wQVG+
vm5+0ViUSLSlflGu2ONCGuVQ6n8hkMNiFiHeu0pDZXYCtjqbSzx5zUgF13RooYyM
WRzd4a6G4BG04z+ZpU+N/7TBMVmbIoK7P5cjfGeEI0E0MSD6PZlDqVCCAphetuQi
tXpTf0XXCk4HEa2aNMdind4ZMcxzBcbpQXnj5E+8Lt1lLo9R1hmhl8xvqO/bkL4M
znEmUBCv1D0tdnEEcjsVQ3wBYn/YNQpNoiJ1Ik6zGxiKkxMtPYdLYQACnuO52cYM
8vU9/T6awRKTPDc30Rzry3IaPqcFpI/C8xT4Ss/oo3LsCDXHiHZqdsNHYU9JiCx1
Eo/yVK0eYaLkvzyCZlX+HRbqFKi3FSoNrPS+cn6yRuDOlg+dcMBpqu9uiHvgB8PT
74FX4CpeWlcRecG+qoZMOKAt697LNQ+s5BEM+jtIRviTm9f/aUnISWJTxji0L/9F
`protect END_PROTECTED
