`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXDBotEW0E3gS0lz1uXnPXTMkFNkMndJvual/jPgnj+wMA5zqd2g+gV7JC5pFREL
65RjklSdDle6sXjTzr5YuYsE6EwdvWmkvOtiT6VoXAX0xxAdNYiQ5gyV9XRpiHmD
ihcCBEfw8MKRykzASnC+bAcb96prWuE8I627v18FC6InrSn733k8yjpwYE9PuUUv
NbPTnBK24owkNjsp6PQDV3HLv+lHgnbUVfZyLztxH1eoC38SF2ZlEXH2M8mkX8kl
Vq11sZn/QoGwrBcK+31QsF/j4w0o6wRiUy7W1bupi2+NOh/2pWYglNqa+4bqBSNV
lge4LRmlr+t6G3Rot/Ou9T0vYPt6XQT1R7pdvaWxMZme/zZlQJM82ZTXysDjKQuT
HYCTu+j4vtIztjfyM3JBoQ==
`protect END_PROTECTED
