`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gfrgYaAj4pz+NwfFEIatnolY7nj1au375dLB1j4u/gwgSB5gjPqiMcwzjrpH7plY
Y7R7wNyBjVZ51xDlitQeQ8Ne9wgKLH3Z2YkENAHIKBDyD79eMr5AqcwS4qmQPz8H
/G7ixRqxOjGkWQnTp5U+S+BjGv3gAR7imCHKMV7GDqpK5vu6vnJ7OeKkGccXcOdz
ZVM2iMB5ibO6ReebnHXYiouhIV3gY4UbSkvHCsCJyv3d3fWJCaxKGsDRIg2ei535
X7W40OyDqmY21bC8/2lkQ9wwHxSmPDo2eN40iEuXU8LCN14duBmlHxZ13I8Oj/XU
12u4kaaVFnTUIG9p/Vu8symuZBOVbFgWt11zf0Qt2NW9obhIfN3Nb8EdUeHk6cm9
2DYsjhtJK3b25hRN6yjtZXTeJYsxLAl414qey45q4EQj//ZS5qZIc7V8sf98xJrJ
jm/RL0uOgh3aVjLjC7tDuP9OAiwbAyStOyxwJyZ8/Wgt0BADeNmIV+Zz8WYsGjLn
LyaYgJIpkWSbCqt6nxbUnbhZ4OEWHRZIJ5ESnjdf5EWDA1w2PgKpy9c5Dq72qaBH
EAbG3uzA7sb7K4zme085VqggCHdtyxhU4YP8ZHgV5gymi6as2a5ApTkOmR+z278P
uriqRkplPIA1oWWG7bjJp9bwJtey1weyp95kwi/0adSEALfhPF9p+W2vUBqBfjVE
`protect END_PROTECTED
