`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11Os1N9Owm6ALz0bUzLnAlwkeN18dFxm7u6kbuVAveNrpIQf3xvfWhR+QOrjGgvb
4if07PxSMQJH4k/kLmVLDT4lMlz81FEw231TwGUfMhhWZx8heorgIooSdEpStg2m
7WZ62SvW7HAe2zCGDgDyu342aGoWhHZ+5NwyhGsvszLqt1EKew2M+mfD1X1N+jcB
GDnTJ7WFNQ6L7JEeRzUzZCInnP7XttQw4bX6+/DaCNhOEGgsoDEk51u0PVi9IJMz
jNBsMV64NCsAX+3+7uCMMuN+cnYJRcy3CRTwwgu9CrI8PCoBf6s0a0yPliSMaSY6
u/TN8HbntZx20wmrh9DHbr+v2IbYX/G8ClQ3ZDTF17kbWy66Ffep+cI5jcKD0t+c
t0PMYudV70sdK3qKdEbdI/iM1U3t36s5l+UfYFRNzgE=
`protect END_PROTECTED
