`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4YzyFmXZBVOHAt3sGOgJZcaUlXkwwWD2S9NKe/h15FRmEofjx6FUuqjKNbC3P2/x
24LyFof63XpdiyV4PK3n37WxIOTri94KGCaTTY+Fb77y71+aGYIlVYlQANYBIkBp
HZK48Ya5+z9jBtBT6L0UUizjMx0fW0vjNqhc7LQ0HzSireC8hzaRRLJhkNDOjgRv
MTHgrh1+fq8p1a5b4N/g2jqwSE5wUzX326Un1un97DVTH2YDNCRXjUwHinHtDHUE
`protect END_PROTECTED
