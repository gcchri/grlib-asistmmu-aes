`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HU+k3Jv0RAS2arMWAI6M6cc+eUMdbkKEyHIYZXsYfS+oRIt9VrCsiZ0GgcQFNcWU
wusy2cYTpIM1wRQGWdDWDXGiVScHJL1UmmPmXDlQt/TuTbNQJ2aFwww4+7EdTiWg
V/AmzrWJkiV1GgvJ4AYMRrqWzeeZLprznoQnyn4zfa2uZaO48wAL/sHU4JjExxzd
8VYvR/D+efgusvwf3nKOvyy2pIy/xAQFPEUJGSo1lU2mrbu2/8eoUXaJfc9Sp17i
RbYXdErAN5sO4j3j3RZpRJ5+MJCP5KBhWK+MVwPWqj1wWAsOnaKRWrtpl1pT6BQ3
F7YCT6fJfSupw0qRNNP8vOHj+XXpn2ZAXub7gkGilOG3uYQNRUMpoXpk6M17gKBR
nliS7Z5ne4g4N/r8dNod5CXvA8f9bOWy03qr1A+8qT1VD8eYgkn/5LJolBbmo5Hi
MRRmePNy5mdEOr7Yo+08CuJMK7THEBdysxKM2BXS0YNBiWh4brEdAoIxmXa7KGhl
inM0ruaem+ca/pKA5+EaQkTY3oK+SGYsj3XGfJZzb/IPOKFQMF0Jq817koJb42sI
wlFC4sgJ6vNBPQTrB36TKqTb+Sbc4+q3rlDFAvarddIv/sGciMK5Tv0jCmOVbbao
w+m+EZS+oggLtfEsEC/o8Ih3pVajcOX5yr6X/eLiWvLqaKFPkaQcmTBvq/eVFAAI
1n0EFGezyILlllSfDir7syzdnKOdCJO6O909STa2S/U2mDFGRQUIA8qPnEc6Vrrh
FLVkWQfSt3YNzz5dnHIHNN6E/GaDI0JtVAcGmEGd5M6inc/xCrEUlWc/HVUu0xDQ
FdBBbuiTnS1xLVQqasmMJrg5mJfPzfz11dZ0e2xuMhvri/EM3U61J7N9+x+7LwRd
`protect END_PROTECTED
