`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTQQFKUWGEFYoMB7WfvJiJhv414sVoNcAENWIYdjuB6km+ub47xqmEWP+iX88f3b
Iw/3xDjuvyalstKRN+SNLlRFcCAVfcJi3JRDNF07kh9Tekg70Vr+UCdLrBJCEU9n
CXrEXAhIiiIwXDrkDocThAzKHl2SccY7KVaUV1uP8ZM1FJN3jOccDJ+x299PeBRG
f/jwwhsZUJ9Aq1NBPoslIakNHCUBEkN6eECcNRQOrnlKz/L9tjk3dHNNGNsec9su
MGl5iJCJUMZsgNOm1a3GAH4RMq8imQjbSCLOEORyTzcE9MEJosjGYscSIY2rHr0C
`protect END_PROTECTED
