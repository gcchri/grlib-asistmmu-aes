`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F1cSfzhps+L2+agkebq3yoSyl4g6hnWJ1VRhCl0nANrbSzeKlHCnflZn21fkjqlc
pYS1/eH7DfvTBQkd6UazrSC5C2El35Z7XNEQIaS54D5Y8it6hO6FaO83YgXrlJUH
BME/o2HjdtI/MqHr/r1+yT/cwtU8oCL5iyEjWTHVSrDxp3LXFmJMIGOIB6dtlLA5
lJ+Ybg4n4ceE0Z+5OcUGxU7/jpZ+DkbbU8uNvz4RbOkdj9GzEOoGS7jKR58oVAK5
LsmMqURCf0Ia57i6sETeHGUOwSATMdpKY3oM2J8yVYpq+BSbGNraQ8vnR3kmr+IC
C/tMjHyy8xXFU42TnmWx4bMBEyqUSWIGwldWOS6kyS9OzVtSxKudSd/A2HUKNahn
UWQbkIX42q6qCX7sKSAUYQ==
`protect END_PROTECTED
