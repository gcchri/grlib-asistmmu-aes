`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYcHr8cdj1RpDmQ83c6PVi327czkpYTeF13yeIyxg5PdLtV3pHFvKMovVvE9Amm4
VDiKRYecVdZQZ6yXHLHURQRQeskH1NLL1wGQ8QaMMj9HLHo8meFKRMFuLmzGVv9I
zuF/rG0EdS3fBczF0JV2e88GkzJKraQmyWp35isYQ42SkT0jIl+fjot+e+QXCHl6
uTBWxpfZnreVP+guOQ/dQ0D8VZz3jZ8di4nRSWXk5xg7TfiYCJZ5auD0R5XxdUZf
qa988EkUI6C/8FbuxClHRLGjNkU/qU5Tjw6nEw+1McSvt+MvihdlcYGKk1+0LsQL
U9jMpzkSILU1FClRzwZLS3ptRheU9MrFxBXLIqPHBb//vAK3ftZJAkY4UYfMoA48
ENNQsPztQx5i4tPvoEZK8D+amnfyOeA3P4QckiY0mzwHEUKqs7mPR8wFjRaqUhDz
k6rGjhWOSEITNUOxQR8ILY4Ra1b8VfZkbjqjVi87n/aQvwfRnPP5kWBBpctfduWu
PCcgYLVR9HrG+W/jxf5prjer81+/wKOcmX+4MJrnn2nROagYxceNpM0fZWLr/5pR
ktpztFUWPYyAy4cPUvi2OQ==
`protect END_PROTECTED
