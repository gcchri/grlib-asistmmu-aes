`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cscxMt0ioKPIHH4Apzo7z72tdb4lgLa9k/TJYaju0OLwkd0WQlsd3hcSia7O6D+f
cWfDo0LKNm4EiCMKHRuGSsw5fot0Mth/WKI042YNgS1tZdrAAaguWxAxGWG4GPn/
qZ41OGGcXwdPfoBQ7I64QdmrDVP6M40D/tq0FfIGItt8xJtytHt3A+DFnwjewZ4e
tzbROQdkNfUkiIQdb420GKvytoz6dSOF3ci+AzLyiQkllD3MXWp//olN30eG04Or
9XjNVGJOvyswaRYeOQvjLso+G3KQ7t7/ca+Td+MgNWOd/KkS9em7pTMtgtFuTjfV
B1sMarrzqvgckHB8A84xgROyi5A+nUUWvBD8SgqnZfCQv59LTE0gdaElJ/576J6g
Kh0hNLXbel+sGUeUICjNzYn0/X6BHWwc46d6hF/LfbNEXIgUAdNSTGIL5UhWerKQ
/YmJwnK0Uz+FADFsfXHTiA==
`protect END_PROTECTED
