`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQlLsZtFdzMP0Q7kjrXn+lYwxwbS0cLgn8FH5ro66AuiZzlD+ufmdX8nsLPl6voz
wvyZgLIY7iEpW1JYBa2ZYPITy/s++wLZwkPXosB2uWtmTgqguem1YSXsATK/yeVY
Mg8M+mID14kFMrcwdffUh2TLgx4ZRfTywCFTryvqLFoE7FVzimap9ympZXDlv+MU
rrNiLJxpNO4ME7PaSqNADhVaqMo9zkY9Jmyp/K239XYsUQo3xQt4MdLgzpU15znN
54iLzb9iCyEGsP7yxSYBKZCZjp/q6ckb5gUw9PDDEIRoa0fyckQoxy2Xe9Kc5d4Y
lzDNIvHG6yWJs8lGBPnVbqd2+z/VM1xVvBYJ8kmHPytigQGuF/aqViZSm/J2fiXD
dhpy8/c79gebDq0H362+7T9LiZQn1w9P6X0NXn2pY4/Biv0xoyvI7B08mOSk5XTQ
N6QxQ6ck8rrBuUiCkCbwwQnXQEPp2k9/5tR/1qK6oMOhnO+cS0HzRxzJBLUW1me5
Ao+vl0wjQj6pLLNKD+ndmn7Ck7xSIPVJDIsTGrvEvKR2i2q5WZ9XbayzfyHXuyYA
bshyI8lmF7DbRFIfXZ+kMNPp8ihSBDziAi2BM+1ulhJk16gsX8AkQ/lUF0NHRXH8
xLIXBonB+hDcy1bT7v/S5of8uIujarWK0dtMVe/nUqzEplpNWB46pUwrcBjk5bTJ
YYOCgcU3HCTFpVPLCABgymgdyYRfaC0i/G2SaDzuzoWnWM+wVEWPO70nzhBE0bey
ISRdtD9W3PkMP2HAJCOIhXmT8S8BID/Q8VyV07rPPHXwxBIZSvnZeUoqIGH6xErM
EDD4DIXIWtiwlRGpO9dZSZItTiKwfmvP1pCI7v98HUIlkeYZ4o8T0Z8kBo01i44R
ymYgcPnvsbcibSHN3NR3VkVuEVY9aQaogIEYP2+wBtFuUtgDneD+FR1Gwc+5xWnH
WCyayKSrZuqRZ8RzkT0NbfsYvfE7PlJ+IcJYGBJcryMYdVtfteIHiPlRcJseftKB
BBfZKAsGTPZp00PKHkgZ9NQJ58QOeQtIqyyWeNhQc/JMYzohvMEMYqpy/uv2PnGF
APtbPFTFkhwZy2GpQ8t/vE/WghE0foPa/KmgOdq+jmQSJ4FotnYMpfpI/ZRVF/ic
TfdR8MxUxLYeffGlpVF3y2YsVSu5Xhip0FNEQc04T2+2KYjD3B0NYI7TNsXiS7nE
M2Kvuq2yIbqFwbPYFecwyEV6tQqp2EeO5TWZgQQLGwfsnR7ZE3hCZpqvGhzvhb0r
tfwoJE4bDNyQs4H544+KE/LwP+frgj98CRF8KOElE0Z/3A236qtQYGds4iYMUMTq
WO8l14GWgUvqDAOqr2hxTtqfC9IgSVSyCaQrp5ZdLO0RSGQyNZYMuK247W6m+Rfl
ivDJYBXfEjMnhoo0NeEkeDWmtKJZHILFGVLrpKe2gV3cKYzBqYmgI/2Ul5EvKjQh
9Za5lRfQoF3nC9VL8OEiNQ==
`protect END_PROTECTED
