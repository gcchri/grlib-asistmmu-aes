`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TCtnTpUZAkTmFu61P+nDy7SR3+tdhFiSv/VQLXJamUlKbkmFHcGHePwLjYBSFCR/
erDpSVZ9TkYz7KhaNbmLecQ1MBxJ964RIwWi25ByO0HmK666LQDolYtKBZ0JpAUA
JFZZUDnB5FbGos+CS9CPM0122hLQQkHie3E/7SQI7UlSlv6FaTv44KiANq/Si99Z
mDrcC3jDBY2sxCcghR9KUdCOMjQh1V/BbBvfk/k9fdM+FHX9KsjHxtdP00xnt4H4
wZMZT07nPmCsS2E/gveVEaAZuVPC6AXe4lGeDdZwJpaIcqMVnJSwIt3InicV55h/
cDXtZs17FUmtwbACTl+LFMQBwF+0/p8jYNf2WoDz2Prp+0x6ieZjB/EouE1EGqPl
yjRaKWIU/hcsLXfg8aMhkoUFnEp/kdpULPLA1CSYYHWaAAI+J1usqpJ8CXq2PYeW
rFB/1amZWhr/SteI2nxTrDYCmIc1uMfk+qSsoQE1GCHTjJStux1dDFVvKtXoHoCT
ysW0KcLvX7OsRew9UPxyhdvDntzYUj1xo+48EkCXUhnY/SXpdDkqYocJlAhauTWB
QIR+76QYNdBGqFSPzES5utk12ja/uR2mBkzVuL8HEDQ=
`protect END_PROTECTED
