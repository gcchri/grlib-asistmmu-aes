`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M5l82hL7R+3/DQK3b7E4vvAESZtNkHqTM4q0Rd5Fa7SFffu25JqIIlVMCb8oC7tB
fs6pqjz09Ld96Sfi9FnKB6aTM4QsC+PzfbvnM3Eq7AJG+XJR3iADv+agsYZ42+zI
AhQO3w+wUEyY5n8FiSc5G+RF4bFwgqTNpRZ+jhr0Q6xCCetHbH6/x/DgBP2aAlIs
I0zPlNORQqVlNtGTVcCXVh6wBpLktWFIk0THsI0gWduOMiTIUksJlDran46qQFOb
vEy3gzPbT/uzl+J6X8XEt9D5Hf1Ie13+ASHPb7/fBx1KqerC9lZhmmxPljUhdsM+
rg9h5rraEOTZQQiH3lqVGAFu2mNZbYxozt3KbqPxEMKxjtlM8T6EJPpaJkRH59cM
xHK/1Oz8dt78NRlvKEAwXWabg+KAKm1DeK/tpZa2Ico=
`protect END_PROTECTED
