`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFJuWcGzqMBK+6mknQ3/M+Sf2NuKpdm22foKH1twe+BuwKbsXtAeE/BOOhMDpxVn
sMU4vCFMzSEvE+zq4uag+f81e5ZVs8J/DVwJ9y7btOG5KKjsJWqcQjlchnM14cb6
DPZSETb6fDaq3Y1OsKqNatiMAv/w7OSCJ7gHJsArl3vitJZ2exAsJNqC35v0juqB
L4MVprqzh0BgdyEPXz+72gG52PjVbahHR+h28eLSPVey9clcZMIjJ9SIR2PM5n7i
r4XFRW/kXm/Z2LbfbbVGxr+zNQHi+xHZxOIVrj1dUcuYs0dwMSNOy40/qC0mp6+L
nkSAZm283dWqaABGfvHYaO22x25ce8oHgtI6LMVEe2gHBFFPizRDPJIXc1Rb9N3e
pjJb/690r/fzII+znHNrIR+N0JcXFFID0g4cQTwODOgBuk8zmiVFvGaJH2TxCBe8
yh9m3wCU2euS1UwzsuflgWg09l2pwVvnO/9rwIkvq0ishJoGH8dnsUVhzROkyYXx
rnZqg71ZtB4RudVLwK0ryePJxQ1R9irT3a8FqbdA6oF5cPXLgAkL6ldgxA8U860d
2t23FdVErmDSFo+Ko6ie1TR/V7Jwy09NO8PHIF++NIbpQOlC9BDAZMjnNWHcZlRp
hc9Q0RGyk60cT1Rt5azhPCuJkR1it+pcjMAOZKrWZWVDZ/XZKjjz4Vv+ONuTZryP
4XyANKlghDuF1l/4+tod4tfnaHTEvk6CEVXZljfOVsiNv6OYNn6IkDyMV2g6A/Ls
b9Y3vHU7eiQE32m0l6HqVSBjvPqaXDDA109RWMP7+g4nd0we9kvteX6hIgVvtF8N
88tI7v4xHHqpNCf1NMBHUFvZTQKGD2YvH4uuZhooAFYCnq4g87845oMi0CLxd580
CGTl75i1XZFdch1mXncoSaHkjlg35dtOXWRJuwH4+9uKhxD6wrcZ5es8lCwo3Jp4
DByrvNxxEgsCQcIhHiAH65WXRujL7n2T9lpotxrlWXBl89PLZxVjWoYj8A8KfRVR
07riQ/5CR0RcVtbYWcu6uw==
`protect END_PROTECTED
