`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eW3RfwRqonn2Ohgm4Fym11mVdppA4x+HaGUc1I2b/iSCDvqI6B4ZEmE+1I1FuxSh
enJujY4nebJd8kG/HM0nu5kdXjit/r//9W1gh/19s4NR2X7o+X38G/HS63BxsY6a
QeTcGtqcSOFXdsQx+hDJjMBEiT5ikxmorJYJTkKyL13d8UFoCjJH0yhxygbk2koq
FeXBJgKxzTNrIs0KgNPK9FuW24BXEok5BU39oFq55yAC/GJYXqQ54H6MzNC1iB0C
LrMGvEWES0uggGThLE8LOFY0Lh9Z53JM+UL8FPpbA+eKqUjNBwVOHa9yOVmBdw2F
UshcSoNC6tLv8TdvEa6OqiuLjYzErUJOURIjh6RrxLldaORk6hYLjkAaI4GoczCx
VU9y1ozR19orMlU905OGsM4izcVZ//LaTCi2CsxjpdjDVWWONLXNcnJ7ilAGOofh
/sENrcGfAJcvGOC9hxIn3VG0B0nzfmwztDX4lbtMZywu4MGC6PtbpZGnPXn9lqnE
J3rRwrooH/2YwtP3iPnrQuzDQ2MViwepJMrf8kwSzOdLyyt881sezJOaATBKxh25
7qi9Eqf1tW1TiEGtRDQIK2gIC+jEfkRPrQiOe0/3/ey1mpiXi0TxXh4K37QAqzFn
k3YFfFgiGt69ulr5LOVaxCxL2lplvIXv/4Uuky589BYyGry07xEb+ITM6Fnsbqa0
ZBuOcdhO8Pap+tCDbOr8G2FDwpuJfMDejwCh2MUJnGIWKhjucLENyTpucjrYJOWX
OgZmoyKHlwiEUvulYs6SDkp6OEJPiqzZKSHQoIB0LTmTMAUsAwsbwy+nj/PA3JdU
IYrEJQ8aLqokgRcXVgGDJbJ7DLpWxewaS410XEvHFSLFVu60FTWFvuWJqxsM6ZBB
b6LiNUpFjPMBlNWIyXtIhV2lJavw9WfGAo0/TV/bzepH28KdxHOnTOV9+y5yvydn
QCSRF6gX+8dx0C94gsuq2WD+tg9buM8+4gobiMyQz0aFM7N2pE4ZkXh8dVEdYzTi
tZx5nhpPqX3fw2yRr8GDFsLSTL+9Os7EyWBWqwFa7+dZrD4nsZTUhtpXHcGs1TBe
nkjZtEHcwVcrBUCoBOtEhnUTNcVXUzsAZTv1oio13HFOl4NW5n26YAovkLdf81wd
KYf5JtySPwdooY5SR7wyos9/OcCQmr7fKjQHaK+A3EC2BqyCbXrGHdgWu5ZS8DHx
TZMswiGdTbD86svchyUHQbp3j6dPqd0QHEb2jLrx7NRhMauawJwT8aeSfUp+0EaU
tRYFMOwZ1oZVzIU6g4vkR8NHdJH43m1vZNyOwrgOsSOVyqY/aSt6fSOuMl3mBRYP
0J19CLVIEogNpxb79uSpy/BfgeQu8cae0xpn6UrKnXsB7qvSqefCku8jo4X5K2wO
ItFg3Q1e4atcj/dXFJ9YiQoaGMxeLBlhfv+JXsBnNyHr0tQdCjwQjcF5ptQJP0i5
Rwg7IVzRIPkvSTOJu0JV3rcx3x6qbSYag8faFkSexUykIBJfmQ8A9nQj+ibzkIrp
5CuMCYUL57wlejd3yELDZ5LSeR3rpynSSHCCtCIlnfj0NmUKBME76ebSlWdDXZJW
joM8Lv6alelkOpXS0qcs6XmR1C0YRBPOAlg7JVX9wp93W1a9w0jZzddMqd1JXfma
rK5QewneTSmhxoD2tAkkQOKEOVQj83yboudzOyKCdFhXet5qY/QfB2M+UDlYTA54
itcx0g+K0KsvEEpZBRQoLKn8CG8jy57SSgEP+MRAvVm1BM5v488Ytrw4pPq1yjmF
vL0VLhjnKVfv8gXmwbustv09scnCqnSsYiTOIVMN6Do=
`protect END_PROTECTED
