`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7OV8XKS2R36eAx1KvUSfyUA/OIMQ0PUEV/3YqFgHdgyeCOxOzZ7SEdFQte1baiJO
b94UPqWGDiGj5wH8DnOye/nO9WW+m1qCu9RVrFna9qREGEHSD1WPDb4KnIzTiK7n
usCUEo2YVlOF6VfaaeI09fagxBWf5shVWdfLM39cVY6FqeSGLaOakttWhKQUm66u
/Z+YKuEWUyezkLFBtCTDUZh0/CwpISfkOie+jPuHV3y1PqeRuQiwoWzJoaD27nSp
/KVAFZe8bHnNxpZcWClEUr+56+3Ml2edrtWFOLUjxrT+eG81QP4sRtobG8ZHBbJR
oMeInO8kcx1b/a7mIxzD6R7B0osLi3EuAFKFoHvEziGIl8tDgE60qX0oifKr5MG5
ZAxukRGRuPC1sHP9KE58WNnqqcUX2x00Wlw+Nww6ls6vLOi02Z7DGogmWjjQnrhf
6LbweQjWPaMmXlYQ/gxbQqEQOcfxliz1N49zBz8yQYBP0cMfM5hO6ggq6DEL0J5N
BDI2DeTa1egmIEBrPuIuCqODWYeZ/mKSoSQHdeKmXiwTTeEDciRYmDzHsY+UtOX8
3jNyW42eKowu/NvV/uCiIystDDwL8RnPi33BEifSOaoscg1iK/IvtfAmnf2Wbklk
gJXb3FeW7+ldgtx1iL/7Lm1L8ppgVK+nUSCYoJNWrmQ9WaiOLRAIhNMFOgUG8vXE
pMdp3JgySY77i2UVWFhlaWGPDVqC0i1tJf8CD249+QbVq/HT3PkVT6MhhfDpxZLo
A2W/cLecqzLL2F9PPieKnOCWbDvjYCej0MzD+Ospqj9YwX1sYH7gtCUqE73KFnIR
+a7JI56GRUxFy6zCAC+17/ygMIQEzha7lsnEJ6SX5GxuNbFhTZWtxgS1JdzFxxhi
eAvZnGdkBDRuYvxD0oeQ1A==
`protect END_PROTECTED
