`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7UNRz/dRCYqgvQA8lrL/fsIJscKkmNPmGjjowE+QBJrvX0ubxizWiUb8BXNxbELG
cPUmWdghBciV9+fVXyQGzZpU76lot0pf9zx3xHpD9ncRnGPEdXmuxpj5dCp81Hkh
SJQJGB8I3CxQIjxFZ25v0KK2ue0nj8IZpr6SznBIxP+p2QSBGuivxvY0+ZEj9j90
PFBhaWB9kMUUdONSCIv+cq0sotMUE+50IIPWAMbSQuhErzBcpfvjPHNgoHS8VxHT
KydhSq13tNZq1ufoaiwWAqpqlor+H9xwJzg49miKFh1j+9/9UrHdcUUnRMcwxmrf
jewW7axO3d5YJIWpessGTxAl1Z2MtnUswmA3vSlMH53mhQoaKs0Vlr8nMFyi8nIG
RJSMFja5KhS7T8GGEqQGoh9E1mLTdegGz5dvoY7exRUy8YrMGfpWXsS6S0JhIjd3
s6ZuRYbKROmiIWn5Db2ta2UU+EAfvv/y7B6Z2Rk+fvrw8gNExT1CpAFVpj/LRQ/1
/pdTk+gD9IKsf6xr1fr1+TR2M2Iep7Ud4bsAQJwGv2P8deIWijqgzh20GhICWf1Z
`protect END_PROTECTED
