`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S5ojOmjEv6Q9au00w6Iu70gWJOXoiNJZSdDEcE8TuHMqWfZgIq7eklCcMHqFCHb5
UdhpI7ygxj2mTsrGf/HA865xvFR6EenlaDDjyfANWbg5q5UsLf6mdaOSj200VyYI
G/OsAKUpjaxBfvjeGiimMYbf1ThNbn0nF7NOtkxr1tcaNYikeJtEgY9V2QkgFdmZ
RT53daKxKwxrIh4DSDwl7C+Y+l2l6k/0kSQOm+PpxplohVLx9lA3XiTSmI8IgXvc
rIdW0TY0vzMYzqD8FInDlJK4C/PB5XFvTZMuYJI4k75dTBjrAVDBW6P5lWqXITjS
cd1k6g4ekVhZktVKCxZf931z/n/5/iIcslwOwVjqXgrMeOyfAdQ4k1ynk7PxVpUp
5WetW8vz1S1IJILGKtTHrGW0HbavTPkzg5lSy8J3hUWHVDW2ulhJUXv0RhUoVYJp
VJSMbJoXg8pW2EyaPqC5Qjwkd2B5ePJie5udBWLCKtxgyjRy24ghsdLAMPYJcrsE
7a3ZEGKPp1XRY51ltceEJ+4eYuwmdXV45e3KxqLOPcy3i5c07bVIVtAaZsOEZFpU
s0gzv+ZD2zTUjXYNUC3Edp1bH4MDLIrldgmqRBDCpu1/2/G4yZsaXMjWpQ0F6nL6
`protect END_PROTECTED
