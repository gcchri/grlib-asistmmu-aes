`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VVwS+/fZfNvsbsd+KU7g6Oo0Iwoi7Kp+Oni3i+QpUDJ8iczCyNybMNpFFahOfxsu
oXk0MirgPlg6p4zQ8AQe+7/PqNMBITXgTO3M9Om0dEbQ08kmLrUemUIKPjAlFXfW
jbfkax62l1WJJY6FFAtS4MsPj75RtMBkvJcpPSX7cvWYsomi3kN5f7J7rKlR8dE1
h83dsivyrmY13vRu6asEPXvqp083RUy+K8qAW9zoeO+81U5tFSkMbv/L7fDZk4V/
NW7IdkOjnLa33Zk5kY2ym/gXGLYfop/YOjCndMcqnRvGGLth/sypHBgcn069MpGr
ZjcSGHg/GlBGC5txsmTVmN/slvF6YrZ/BqAwI/A49ZbaqfeWAgVFCD3vY6gFOyvg
3drNOV8bW1VBfE20KJwZaQ==
`protect END_PROTECTED
