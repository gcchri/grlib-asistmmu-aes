`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+iLDCLqSN2di34LbWoG8fcAP3X/hdeGyVw1zoym5+BqyGerBAvqJ6QYz6abRUqvT
9athxfTzTNR2CLrjJ6O4QXoC54CNTstPR/7uwlSberE1EsqEWJQqW3CEmaf0vRzn
Y0Cq7mxwhTVQPkuvYGLF5cCPYAAz53/LJuYDsczh69l7pYn+rT30mNkdWTk1KCqd
/Q7Hj92HoTcYwYu2sFSTlgSkE6fh/zjvPDrXDjQaVi98QLPM4c/90Cf/5kVZ3eo/
OJ0PQOa9Ogt/q0bF90iuwlEVek04dqVvI3gMGKV3hTkgjcPDlIIHpNcYhZlZSB0M
Wq9smIB//0HHSXqt3CrfgAnzRQ1+3QiUQ6DcGihuuoz32i0NeJxb0AEAAxSeXYEp
yVbVPMf1Mp7E6zNm8f2B4E0UbqqsppJOPTMU0m2MgQg=
`protect END_PROTECTED
