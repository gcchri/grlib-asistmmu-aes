`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cs3FgYNDXJtG5a9W7FCW0I6C2/5YVIOWzqkKRnX4u7R6bNbYLg0burbSoaTSK//J
FgtB7aoBb0nv95ECKszG62R1ws0zUDS2hyckoat32I84TukvbvxxHYt9KWAOLP+A
59Bbga7aoz084+ceDzhyDtMZ+q1bzp+aIeM4Vuy4Rxi6Tm7OmBYQ5hbBBKfrb/7u
MDKcxpKL39FNAZwsnv2ahpNZl0BUxFd6Zq1oT2LGgFMPZpni0wfuOfCXJk7zDXN9
BADFqCFfL8ji6vyapLk7SHXP4qwUHEKDchQHOUM0eW8tnqi0GXJZundOuwty8jTe
pWvnBA2zhSQIJMYkJMq++CuMiSQKGsZPven0236HEMSmjqCBW7X2CcOEqBPJzXG8
PzIfXs4CRrNsk1WEaq0lPBK5R8ny6bRSdSDxAvauFAyXZIKJKhPRyCnvOd79JPHV
`protect END_PROTECTED
