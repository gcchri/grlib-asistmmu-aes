`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZNfjLrNluhbnPuOvWbA2i27oxzjzSQLk1hwSjrq9uAY48ZM0NmT5aMgQJ6Q2YkNw
n1ST81mT8dO5BytIrjbDD3hK0NpDlRUcGjoDkmK/ZmgdjeV9tX0/K5/9yRyYlu+y
wKEK3cujEI0ovYxGmb5/N4V/m1u+PBJPp+zaG6YvQNsuATCsT5zj3vuj8ncFlCn0
SqFh1KnFzPBEzJ2CjfT6iKPC4cBcw7jraNb0QvLhTog3++ccdKSB52LMnxKScFzh
VyCvOUfSgZp8hqz4STu+I5KWhv/uZptmOoqQakKuHw0wTD9CB2TiwPGVGTKTnhtU
LkgLBTIsXX7To1Fv110vgJ+DzTerf5eeAfzq5QJfc3mGqjBixypHw//vbBub4iAz
jg8pXGyo+dWKj6N9FOYMDeDBBn7wcQI3inH/D18lXnXdj0ONKq+GP1pNSO+AMJ5O
hzHa31TTbmUG7h1HNF6y8QwUU8JfIKp1JS4822+mpU3h7Ra3HcBnALWduiYWUQnn
ooIiiac69DSlUBjpp5JHAWSrnQdDNuKD0PM6QSCDMlYbv2Kt8HH1+owI0yp+py+X
ba6ieSqcaYVGGh1TN2imKlCy+G9w2v6ROsryA6YINvA0IiVq5UfTAgtN37bgAtTL
FKXgkwGsGTtqrym5zgtsRq22u84j2jWoGCNhndYf+0AYxaIe6AsgLhcXDTku/kB2
U8zthqQytzBmJ4TlYHCpzhSrkyJBoqEGbSRW6Kvq9VpAJZDCmeB3vcLJFCv3ULrE
P+3TqeikFFm3SWfrSB17iAQn9bRnhKMCSt/5G1H47JSwGp+VygMTYDzrY8bcMkwE
wP2MppTpn2eQ8Yo/7SsVzbrQlUKx6BPRT0OP4hKUNYAScEtEaNGcygwy8Yj0GMl5
S01C3zAvopGSRDLgeFgUJHbDL+XMXcZm8IY5bH037kVc0eQhL4A1vQ3s1a33aP2R
Z6RdLi95VlaN4lYVsbCh/hAh5pfRgaW+Ja4uQE4mWtwbsSIgVQxwdgMuCQk2aOLz
s4QpYuUhp0cxyHFGw2Q2Q45xL3QtynXafJFgCuDy7pkbr9PtDyGY1X1UQ+7PiHcx
0AKpetz79W3WFoprAM4FHVZB7cEUmOfFk0WA6xzeeXmgkZRrE/zKw4UAV8wosBR+
f9eZutz7AChoardkRqgXYVuZ9d4bq50Mlr80nIczc+Ivk2BKNGY699B3EYk85OCG
pqiYu+4umHYoBofS3s2R7kcqxOA+/oEZoQ247mS1jA5o/xEL9E6IYlIjhsxNNeam
oMS3zHt8yHlgJt+oCLhSqbLtOobwZyG3uf3+EhZMGHUqW5hYhWOQbDC9fjIDYnsp
C41ZO8K3cEwNJJ/Yqv+mHkIzSCSjwSEfoBmG12gSFoDubzoKZsJSNmq6CBufRYKL
Idf/8YU7PIZzfbkCFOn0/ucSgiixdyUVuSEC5W7Ks+NZpE9V6q3hBPHYioeel2vR
irJhkB3BDYr2YaV/bs3wmsLucijLMdp1aiS0poANq+NBCEWp/SWj9D84MQ8ehiQv
qjB7tdvUfor7E/atEovIJmMhsGg+TIG2shFn9gGzqnvuZABVHGAI3eGosn15cJRa
SvjPAFqlp9Y+h9iWMn/6wLfMmHEYjlN9g+j1yNiuxw62XRdXFhpB9zamDmVN43yZ
RDEtO0d0iREsDJ8fJTp+aQAMgDHN8UDL3Br+kxXV5AV2Mc/jABvf/lCYY9ucaTLB
Yl15/8y83Gt7jaelDWZUqSnJRzKGtKcPC78IJ9NXnlGFwG6yrpFK5gCXB33qntho
j+fEk9zFxttVFLjOMulgpXbfbCep2xGMrrzlPwzeMqknP1p85ZO9WyX+ME9OUkft
GZAdTcN8b4o+aUFIm1bCq4R9kHezGWWt5UUJyxnid3GavVLvFMXx712hQziwjxbM
kty8krgpzYd8fsB7oUQoeovYQqqU7Q7vmuazoFMV6Qp7z9nzhYRLGVqavLACmVY2
HQ5xWHN1OEm6cpmN2Lpcnr226jegEwVCvGYTn/F0EBJnZ3SCquH73Q5DSJFAVmA6
z/lS2fLuXn53WW7PfaNSl33yV+Ngk3iw83VpmbcIA/WhbYGdPBE67w7h/248WcCr
VOiueYvrcZDLvTDrCImu9ZGSVZ+/yP9wHFiM+HCGcfnts0hVSQVEZhqYbMQKbArq
4x87nZFaGL867Cid2rWf2y30zyTiRVhZhfcoC+Y9Rz1eg1w/15MkCHptTKM7EZ/b
ygmPzO0Pi7KiEe82Fjr1x20DoWsoo4LD93hkHvdSYF0Gxs+vMVoTIG2yYIYvhQr5
7+zjE+fMlh9olGPOKmDTDUoKQrOIyIzvKpbbmIGvF66GtUKbQs9rsBzng54l229A
vGu/1L115iB6mWlaZRP6d6RScEeo+u2sVXaHR5RuTvnJDsg8fFxftYvubpp+6Iv7
+0tp6GZBm55tPPAWS7T1B3OGEGtbqu8Wzy2mD+ip8diuCCx4/dRAcIBDqKMSsSJv
7rktSIbv2WqivO/aGG9/C/+tAS2aM6r3FcwC63UrBwjTKUUqPxM1rzZYAfmtQfJw
qldu9/o8CQIcYTYrzBOaSWR/yHl6W9Pcb8sx3ZGA7rrQUbJ0B/tI51u/G0f/wzWi
gLwvk9z7q/G48I+KDSb22560rNwqDeHmUieCc/t63ICVk3w+iHDQ7xBwdENeKRhe
Cp88CIqv9RkXwu3uV/nDuklRnqa2CItvzgIZbKzCi7jWeYj72at/NSSEvsJDO6Sn
LhCwTKdE9rCLqvrlrBgxMIL4/yCAfg5dpFjw1zt8+sW6wWSR6aS28MITAv0zYUQf
7MJnqQ+idNzs4qJxy4tF0NDhsfZRs89sWTCDjYVm+4J3NXP2Er/cjEOnP8bzjxXj
s1TSFLZrBYVuORi+09xakF2g5OB69Lc06DqnQyEX5QF3HTuBwrk4TaJb1GnXaHqA
P2ODvJ2pKw+tYyggGLV+Ev7fdiVoc4prfm1zc6depfXUX2uarSnYyJ2iuV6JDIZv
1Arl3hGC6DST7f7KOfPnAnlsaPReBt8NQDCENhdJh4TnUmp0PdSpQPyVe7Z2wN4R
MOGvuKGs5CQldLBMP/v5/vdatazZJLsZL95JUPp2PWoSVl/BIUjWAQljzvcXJ0iD
aYYFqN2A5VFWUs7A1ZwhsNDKSArb8/31irJvhYIzfojPJrAMnfVQAM99PeeAuuNB
RxoHbn5fkWnHxty2MX2dmeY6K41mmJRoSG1hRxwZ2iEapZRmdoRPAKHegH13MEEC
oIDSs3Cb2gkhknthJOT3EE62JHI2TvHH8sv9drdBkw5wI3Xh+L5C1KtKXj0B6qDL
Qqckc46RQmkmhXdU5koBSbeGfbG2A5av+Td+TmODGUOn5iY1V3sryeU5zMuAPutQ
Q7Su/Jpeo4jfGdUXHoKNO02qsbAwbS+14dScnrvUs7N9efk5K84/enlG7wi2gRV2
LeWnyw38L50H5HFYDn5GdezD1S/VKZGRfKYwCN6WORpRXk/Eg/nkRFcHFEMOwT/d
efL3t4k0mZ5GVDGB49HrmUFFIP4aK3KwW1H/jnrc5THIaXVtnX/KCWZqCY2S35yP
FyO6VKA4CzlIlOighwX8QjAaPAEa6Gnv8GKrxT7ynT4kufKyW0UElY3nzDfAnOsi
5HFIKUPTI4ER/3icVipXwLaMrsoDS+da5kPwSCh1n1JvHpqUQ0v4aDNgyxbS5RRC
RpRO5xviVk2g9k+Zpq4O70JchmDs2wlqoR4SOjPSvZwd8tD8t8rC79zkfqma/vYq
+oTK48UKV8z6ip1Mk7c7zw==
`protect END_PROTECTED
