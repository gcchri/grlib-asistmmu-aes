`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eSWOpaNRsG8SsHNDKmeKU2Gs70rERQh0MCrLNXPIwHzE2dSEe11Rg50nK2Td9U04
032Pi07GVTzujveEfbodAfGNZAagQ93ivVwd6HcQdF80KIRiOM3KdNxqbWlvhPh4
3kLbkXImK6Clhsabj6Kdl9kqBP9GjkweRKf3SBcgb2mEJ67bs3iMcLiy6ygNlohv
/h6TJAEQrD6B/mleuipkvr0acfRJ16LJnxTwY016nbEQRadato/9Qf+Uxq1tnny7
/KjcwXYiZ7q5+yDuwUmFtdPomB/GBfC9HBXghGu0H1Zca/yaCOyDKAg/fBsP0yDp
RW/Jk5j0CL/PJA6Rm+pbVZJFizuD09IrhwrwzgfrLFeEWTMSFsdIarMoV/mwWEeu
wJ7NNcV+HENZ/ZYLaUvNNo++JMPJA3b3LY/BjdtPcE4bmjq4YzTEIfENsM++QNc/
yyom9LG+Zzotr4pjoRzcvXeoCYcS641OtkYF2UEc/Y+wWT0JhfhEtAfvEqybxfHO
d9LiP2yCzq+t7P0+igsOL5+VVZXf+YmCGK1/jGg4zv8yGu8Rcl+ejC1SZhHUU4Ak
ifLk0Ajh08ZW275qZbfmzB/HPiLZU6Fjpqpdo1PbYmbrMXdmOT0KiyUZYrCtyan+
HA5vahRO/U3k2jPKcdtZ5FadVPcbFN78/472JlEKDPJ4tJaRmx1tL2OAfKUIyGZV
Kg8/ZqvauPIn7Q91TsZAJ2lIVJMgmyyp7/eyyOhHDRA06y1rbittWQwgJ9pMXQqM
1YwQuf+/bSfq1IC+2E8+ZUGyd/eqQs4x3phSovoANDxiIZZHf6dGDF9Pv7wPQi6U
HevHvgdmPtORq+EawPGAezoK6n20HPn5mIuT+hzsmHW7MAPLS0MSaKPbLFTLjWdb
zeiEV0845rsP8vOYB8LvXKn2eQ9qJ+gZ6pikx4YAn9nPWMEhsSEcaMRNlIfYMIKO
B8CAbCE0ZMogsHpO5hbd56uSSPH0wafVApZB+CjVFKJcabi5Kug4VHOobXx2G/m5
ivt1Zcimq5N3O0yLQ93njqI1BM/KKxp9siVkJHFHt0uD4eDF4pJVBuz91I1QtCu6
Saz1qa1NqPjKfYD+VwCmSh2MRi5xM3riLlb8h4xYr43x2I/hR5//uMIEb3peQ8RE
mwUTCk7xW5fagK7DXZWxT6riO7MuQzF+RrrJ7/YvQsm1tM5AkR7ow9ZTOQAQybDw
rCiwSadQacZ39SnPV8uZlw==
`protect END_PROTECTED
