`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UaxjeFVxv6EmNFsOfH140M9aW8qKVNjG1iQXe6SFNTFnyPJqPRqUfSNbAuQDGjMH
zJjhiiV3E6eYN62D+MX5Sqr9ZDerPbJxyo1WXPf+Z2yyLsOT1vIXa2J8a1MICGTM
mXeyH3ISAg05mDsOuscdRllY1JP+YPk62uyqEeY8EeXVVYxatrPjVmENMWPzt7L7
LZvOQe9a6sS2BCVydrgUd0grn4gb2dofn7EFZctFeyOA+0+4D6ef98hQA12q/BKN
DD0F6pgyR4KxRHmf0t3MZ0RL1XtT8DEJENrKVLxMPGA=
`protect END_PROTECTED
