`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NRnn+8mwQoMBefwulZ8u1H+7pajM6h9IOpmLH4fPn6rBBZUjcR8Gqg8q4HjyN4dy
A5WLxpE42dQpkWmehNIMUiy62qTymeSz69BTsF9Yg3nrWl55voxJprLxJScGMD9m
VkTjUKujLODwj21/ntE8DCNtytCaXSaICrZh4gBkcBytb/yob5NZU+x474QYT2w+
GV2viLkAnixXUn2CTXLehTW1oJv3F4KkXn3RyokQsqzjhF9bugPxWoD954aJFqvI
ld5TPXrlTyTlTHKOcK0O++yJMdY/KRh+nH0BGXxm1VeFLLcKEMhFaxzVZAf/zLMk
ub4ej0zGjHECFDQa1LLL0D0M0k/KhplqCeGC03mT3rOrBDPXpfl3oYPriK/SgblD
UcG7z5sxD8SprpF+owm0TOLNMiSRen7cMvnV1fOX1A7o7sEEnlsIIKZskierxOf8
iHSziifJVtGHIjFFpNJs86FEvXDJf+hdylGOd+zZfr5W/fUPRwkLTT7OWRMdwJVc
vSzVEuYE8H49YSjGRuuuCd/pFTGZrTA5KbHgXD2j2QAQJscZ+m2Y8HR0DF5L8Ylj
kNqeSfTuHD+mCfnpGa71lMKBdrzJvUdT9+8kIqiRqT4QOTtRzxs27822lg9mmyWD
1O7Mp5ZwPU3x7hd7Sn3p+ERmaVaF3lnmaOLIZXI52ltQAsNLRmhslcdFzZBhQryz
IJ/awxweSjuVKQP1veB6rXKT0XQJPOIxBusnLphDrKz0tthS/4b13J7Kr8yNQvx2
CeVFR/THP1zn6DaMZp+f5Qe4nnnLhhXx0sJmNt1LbgPLkKAnEovlAox2RKQktJKd
ft8hpuiX0N1ax8f1QyajOYZWON1mDkQj7MC4xvkNimXNQ6lasCbgO3JcHRHj4QMr
8x2k8YtT8eMmR9GerTgqHuomC6xyKuNLDJ69b2rnYD+IL6MLaZP2Zxedsk3HsGS6
PvrVPfYXEwisNspxwz3KoqCIDzHoLk5NMhwjiOMKTvu9fRlHCnOJz2q6T4Ah0h+E
O8fcfS2UoQbSrG8yAkazBQ==
`protect END_PROTECTED
