`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
05tHXdMojwvjzNTAHrzzKyQD9XkemlnstALOxn9AHha9ugze5EvKxPHgeLkaNVMi
YNVT24nAoIfIpYspBP6YoTVylZvndBvlQQiEE6Dii2jX5WkFNYex3yMc+8Zvx92a
58OkVJDCqdUr8bCAuQ0O3c2C7H75YFwlX36BBZf2V5p7oiP9dHOb4iVOO/jbfPyW
EF8REA66wXQV2vTtZCbQLUSYNrhU7EZk44R4o8QiDoA42s7kVkk6NYKDjNpfo3vP
bikpNug+VLiEB9yN4cHD9DTmH8hblCHQn0kM00x02hBgPUD+QXmI9DvgHblm1fX4
3HEtilGlT7aZjp7L9d/RFJQ4bSAUsD5XMv0gBoYpLl7WxpPeSOdWyk+NUNMU/W5l
6wO/HtlubBFrg6t7JVw4JZXYyz9N6H/9YqoWQ/aHBZX/24Ee0JOQi0USaqi2owmd
w/Bqus4W+OnW2xgwR8oxvPjpFz561YWqxFCIcFMANTy/SYhxvhI5Kr/7ZVzSkxne
KQaAMPrbgwEOu1mDxNL+u7FYZQGN4XYgF9KE+C6LKpEEhrqjETk1WFuk2d9pmi6q
PVBPS3gQyne5QRcSLv0yYPGw5i/xDwHXeB1jwHDza3AlVgbOe6+KH3LFtdKCU8fP
9h/wvfzu9aFYQ5PbaVH+bxiY7McUrr1lr2wWXVyA4RdS4G+EWZB9O+bapBTaNClT
RAxxuLdnTw8ZjDPB7llKnz/4UFKCOWagC7lYE0THxy6gR2wMweS3hxIG1mwqJa0C
Hxl23x/O1f6v24GjHcLFTHXPq5jQbCQ5WA2jG+ITAhLS5jXo5N2PQoazIvZUJKGE
aWb8ED24iYsHhCvLb6v+IETcqncDw4KTigGFAe+KrMjlqMPUku9lHuTZ+/8GcjpP
vDddjpchYiiK8kgMU9TClrsUt112HFOBJfyItzDjkfbHmpeGOJlYmN27/8YTu2lL
i+4nw/A34+1iPsnc6/nDgzo918o9ydlclbNyz0/JMMcYnYbX8ILYrYr/NHFOEDt+
uR47VlLHNz23tm0FOBhfDmYZXoVDksgTiW85TqX/gWpD/xk0mnNsXgdafyq/a6So
3iJB4GGiQlCBoJzHG1ogDB96tmfPaVol+K19IeQpdX6dqV937bc50Ybvh/NbAkoD
sGPeXPQaVOMeunhr/oFd1AE38aNaBHCSmYgOpD+/vqveNHMT6Rc/UPxKX6/OcYK3
p6Foscq2Szv0aT21kSw1OUqof6Bn3D9J/EQiD3tBRDHDSokdDP9duXD2UTPf2qGE
KXhUEwrr5I51xivGN7RSjcRjWyvafKM3oylak+lqWxJNUS07GhsBTRlRptjP9+4Q
cI67gwG9sfzu9OsIoT5aXkPfm6zB5PO7oX9jZ3prgRg/etjjFHOvX1IB26l6FTUl
qNrS7ttQo4of1NJqoMTDAOfZCvEZyDTLxDUfDNQbaeSeJa7JsH/lWRzfr123/xRf
JPMPMD5iMf6yZW820YuRLrALLTL7+T6vYKU4Uk6BBiOIXmlSceX/nL7gJhaeuLsE
gIe8NBI7GYEayPJ084YJlejPqUcpaxazLElJFHHX4KcPFQ6Vn1idi+An9IYh7Eu4
HnTfIdsbkgcfPdWxSpQ3j7Zd+0f7Q83o6uuBQNqpkSA4KEGxE0IBPlQECFR59aq6
MfpS35aRlY9PlRkXRfZLr6v2Q4+1c78kKrz/jnu7giNG/YokCi2Ge9nxsvtfN49k
PR9Fwu7BeV7Pgso/X6vEqzfoC8tF9htzIAd1HmSemhVoWgQlnsubtx25ywiMWW+4
wivebuo8DwGER+9Y17M3LKbdG4U4ehI1oV2mQaxYunIR3IKuabpJHZZ6elnNqjLR
Lc2pm1txfqTSeml3RyF+WgIxyst5aolWsMl6ukuksCSbOt1smOWRVm6magEx4h+n
3yyrABVaPe+Fs8bMhITjAxIbkBWf5HLbGkxAurySbjOmLqwKk+EQ8ckmJ+eulLZM
8WBXaFN5ttPXYrbSU9niNLqhp07O3EPsx7SShN/kqCAn6ZNzbWiWI4jK4CwDMz+m
u3VjKTA87dhfUsvxp9S1VU5z2xWkywftqwU4qyinNey0a3wK1I/EwijCyFJwlyiN
Zu1fSliqb3Fh8qEhJK09nVbRmKk8U9Rexe3qtF/yO1oHDMZF0yONaFyBXZyEtNj5
/aTM1xvE6D6c0qGelmajO/K7GxoVdb2O3ASUdXGFxQMMXjCBIq8LkOPUMASKdG3m
`protect END_PROTECTED
