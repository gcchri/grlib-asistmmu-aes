`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGC3sgNFyjEiFeuq1Q+KF7OoUOEn76RzxqTSvhia/CDdFzZxTRdMYYW0KCm6Byb5
fnGHia6Z4oQViVmNiOFzFLRWrHOU7k3CsDRne7P79Y6VQg10ptiXTfulhI9ToTqd
JDGusla+oAbyzwp4RVOE5rIQXHKXIUsryCEtktSgdR5dcDZ2xfmCcb1ttbWUYlbf
Fxl/Lp2VdxO5CVHso0rbGSWrS3bS3C34MMzYsCKCOj0liq6xoBlUGOQu6Cdji8MA
vkGazbyiU3/ZR5bb2KelKf6gR9T4nSNzXaJOqfnkr48FYUopNKrl0QX1jtuWQzZc
z7nol/7jjou0sQOliIzxu0JFQOIpejIjp0e526xDErSEDySxxVnJC0PmVaPzbm8u
xI3o3Tf1eaEMrmVwW08mswY6ZJ4WJrdYYpi6FfhklghPhV95+vdaKXdtsdjrK0e2
zy11SwMra5kN7gb5VomnOUNc+ep0pUqjambT6vFov0gx1qvBxJZqt+H/by7EXwa2
`protect END_PROTECTED
