`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
//U+eWoNZtdB57wd2zjOlz1BiboGt42geHP3OJ5XeUkbJu313LWj9PwW2ookJuEQ
FrEod3dzoWDm8oiu0Be6zW0DcqELsTD3Cvj5gELmPljIIIQhJV9tybiDzBW6Gqlk
5MfTDNx+/Ed5/iBQpddp1Sp955lqAh+XAS1UOnjxK1HcNhvNBfUFRBNsuGzmt6Hv
bDmpfU4ciZJm81csZnPhaae+vUqj61LcmnVfvHM5EgtCpBENk6NMOZd0X7w+Z/7d
eqLKy9ueQ6QQ2v8yQG9ommfPFhY8WQLKsM5auUzpTKPtGyrTsJeFu1S400EdzaKK
PeoL/kZkJHwN8PThS799qP6JjkbsgdVMby3T4ISD+sTICM0qLnDCTJSfpAvRMP0y
Tr3i25/cCB0JpN54EPg10PORSHYpgxi2At6oOA0QV5ovlsWRDt5++auSqm/V7xo9
0fe/KE+Bmt2GESIGddDwGqwFvM61T08iZthOCeInOrSBitWnUmaD/LXXzZtpLU3L
8IQD8CX1vYh+4i5enRdlDKJCgtmWGJTx7USb2Qk9UhQjs1/AOnh/jKslkjgBkjnk
en3dRvYdf+YP/qw1lQAM5xUF9LgTJgxmjvyud4bQ2ow=
`protect END_PROTECTED
