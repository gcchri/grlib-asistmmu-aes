`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Gvh/eTPgDVGsZwyPcyAA3DezNHw0Up4zOlNsnrxI3jDOPWRg/UCMvR3BuzLCL9N
ZKaxAJ1wSHIaU8crqZ1+KfjOpeGOenUFJjLaOxDmAa3aRonMcpSCxJjkkdfv1HSQ
n5w/U39HRG9YtKba0JeJKzu0zREMpWMMQDcyFsEek4nnc13B1cX2jMCvYUGUNpSD
DXgAR56tzxn1YW9NavU0crYIhao9Ru62+4ajvp6qGYy6RtPkKvnmuXr5n69ftrfG
UpLo0+dKpeCh5qozT8SJMjg0gtXSNjqjVT5Mm5YQj2uwIV17vlbktp0RnsKQde7e
SWZ0+feBDKazrlq37CcuJFN7YaZiNnUs1D10aE+Og00FFu3R8xquztlUtlfcwsyK
1hfmk0bD1PjuKf+ZzxUN4gT/wDj5SxEeyQ/QGmGj5kzwHNiTtq/b7onybftR6Jao
YmFpj2VZs4QmJH9hi0Y9im3R3LW+GQjJzjcAuWL65wIs6gELYzq4hErZNf8y6kPo
`protect END_PROTECTED
