`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cGLCk544FUbw2WO4u0PkQFwmqP45lRZGazYqbL6tX/DrTXAGcUBHAan42rnz+xkj
WtG1QPHRXCPPlDdsjE+BRJ7pi/BVryvxY703qZ5b93+cssTf3pY5R3QXkdjWPB5W
nwVlClJDktSiGBmrwEXNN9Fxc6pNyDHB82YTLKnieWIMiSuHjUHfB2jppTXMyERO
cF2GMBhMMHQsJ1gjk1R2PcFcE5PJSX9gT5UugQg6LAy1AWFh2bYQOqiBUkcvrrIH
SElZHM+TecRI2cvsdMEkqPc8FVsX7wGF+NGcrvJN6mqWMRAk1x7OuSjuNNFj9g/K
pRD9PBtbI6PIKrK6a9rKvyTLJxTz6k9MdS2Rkcr2UD7g4ogXuMhbR+NRUlEH9KRC
E+HlXvPYa/5FPy1grSKriOegX/u0B+ROFLNBoFgHf1gUXwfIS2Rz2SVYAlvKdhi+
Qv4cdG5bbrPEkj/Lc5Ac6InnSs/1CJGKWlfHCNo3AR+YZY6PXNDqDT2t47PIygCv
OLcYnb1nZKW2OjXtd3HGGj/lSv1WcbUuFbDSqj3l/UDUv4BwQtbFoqjF+iAInTKq
8gEWc2+fE0PZNsnp+z3zZ+NaH4srgpPCLwQ898M7FJPkpeTuK1YmyXFHdfcFlvRT
nnnGIkucOipPTuC2z6Mda0rdsCX5uSd1LAcbFs9VkjPWtn9mJT6oHsHHT6YuzFwr
Wgzn9otgVnijdLSgu1vfKLsX0yewHHIZaSZYDTyaDISM2xWKJlGH8POcq9rNF53O
rNiFU27+B3Xwh3b+WGkR0HFzdiabqYCwAW7GO85itqrzidPwm9Atbd/3cPIt9IxG
H5Tse3f1MONIZxWoR4rBYBSTkRwXrByZTdgqjwzEo7ol++V0gNPT0ShOimTWDW/+
tqsyD1OVYtDGaOoqwCt+CcPaoHAIPN7lR6CWsf08gudOk39GokR9ugjz1yRJ1rso
`protect END_PROTECTED
