`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QFuF7mtLmM/lTNkS1UdmWjyGAJsEEc1xn5Ek2xhNNRv72d+wlxPgFUVpK+dTeqdu
FLQ8lgG0dZQBJ24Yo+cQAL3vEb+4r2Pwd4RFkVawVSFKGyOF0LHnF4Umorm74TSi
LnOo86sHC+CTXUfw/2al8r7XAogUGjsdQrAjpiYU9MR1Oo4W53KijC7KLWPKD0Pf
Cbnes2nNbwgGJLRpYlHmiseMEnKNSa54rYIoNxC9kyPUN17czYqwOin8+TXD+hIh
htuNvCav3M5S14Y1mc6UTHLqimY6JnaaEaAvY8nPNsW1F/5x8jzbkn0sHPL2Igj5
tExBSBDaE2ZPvLUHgLeqxQGIlrUHJsDMq0YOsa6fW6mJKeNJYPgLcQprBpFKY9IK
uF97hzxXWYHqxReXXxP2MNq/7pWp4Pp5Pd9alhEa+XXl/+dyGtyS7YZiPriWi8QF
pxPas9WnoZPR4WOf9K+k+XP5owsqFDCVwOY2nuhZWYiNV4iHzeame3t9jFcfmi9M
c1ZVYeQOuY9+G3qV4B7kAlCwY+3uKsvcRl+480MF98DCK/ko3NIJR8wlP3/LV4Ge
3GA3gLqR1tc45dqjbCcc94fWMo+/BElVhth2OLBpGdiR40LAKJFAN5oOZhwuMjGU
JSD/ROdezHShBcYT5kK/soIh+h7AqcaT6J96f3OHtOwVY/6yGaUqkr5GawXKqAVe
/RhQ8kWLo2sU9uHB36iS+X50Qh/Z2TCEhqshNo2+ZpAFfEdkAUBTvST/nwY8Dgs1
kFiFIXbalp+8E3KjvNc2x73M/tdssz+N5LktFSfazCk=
`protect END_PROTECTED
