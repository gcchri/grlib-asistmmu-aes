`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiayBl0Uzu0YY9Rqc2JtvR+3j6Qv+Q+FL4PqRmaQD3eIActTtMcysZ84vlKoPND8
Cc3snrHP1NdgtSwdJc3lUS5OO5N8eQrRCMuVeFjyWmATI1d8fOwcCyoC+kzkgg4i
Jl/Lx1unyxbH5KnkhCFWjtL6qGGPIngsKRfRK/VrvRWSRmUXEGiXK95bu0LD5LSW
3fRl/OHbVKBRoTCjFPyvREf4CzZd5VWNH5+92iHit4vv2vyfYmzDEuynLTqWN2yM
HYQJK1PXs/lKFghbu4S4E8dvHWer57W+WiUbFrYaU6Rboj7yZAZuuDe+LgvUuSB9
Y2TJIobPpeDL/lK7nvAT7vdT7jvqcvOPRBgHowifSbcX6yZkQuSVCj02K7mF7BY8
VDt5bCCtV6MlpW7eiWIUyuyciPR7Rkd5NFxbI3lRMCw=
`protect END_PROTECTED
