`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BENet3E0mIOspvzXuNUnGDfd1f3ugI8+58ugzN+V4b28jXFp1MFaVw9232SdAUC/
JlNRcLxVItlS4vpP88dlK+OkNRejzRVFRd07yeFaeOl7aYi8i1yfTjW2/7P6AgDL
/jn4Z/PbRsIi4BtQFYAdUNEAlTSKFPz+LGY8aKcckdycqqk+4yXbkIKVNcQtsph9
pLVlD2jL9TqVH4uDweUAv/dHUKPk4svH/QcOVL1Hbm2kSh3OgB/Al3l9RoJxntCA
ufxYolCxi8LleR0dgpU9oa2ZOsaTzkBrVMOD/04Hhf3B5kOvYQqM2ea2h69FIRSh
KtvTHB7ha0jX6XFrBQmYfIL70Q8c5+XlXbT0kVxLKG9vKB9LadeVa1ui75BdB/ra
2vxg6F4Cngsyomj2uEIrQgORvKbvcjAOQ67/MZ3cET6QceqAdYjH2Y4zwY5aH7WZ
3Y23WCVdMarNP8VcGJda1FNoSKUPyUXskZHr6ISjUXV3+YUsMfT1PJX3XCxtR3YL
wQD9icZdq8tlICLb+hzByWzBpXciRPooNdAGOddiwZwaS39xaLD4gklV8Bu3qgmf
O4rAStzUmUjh9xCn+1eiLNqI3awt7604rL3Dq2BE4+w1CYjFQMFZGHU9wD+XXE/9
lx3jZ3tAj2er3ftlA8s9e7TGbN87dXiLMYO2GIJb0dcKGS4PcoonZXfZwJiC/k4e
sU+SsLsqkA8u4+HB4eYQORt9OSubdohgzGTH5+b71jzHDv40EA+mO+De4M29qS9Z
SOjCALvMfxVzTAC9I6iDS+aj6PX0ziwyRUgLBRseIyoSDLrWFWZFs1aHzQfUP/VN
YrAaTvXwlmlOfhogddjnySbYI0ppw6QJtzcbTwrpyduezuqYuga8BhXHDbPpT8l9
pUF/YdhgAX7IdY5nMpQ29omdLsz5uQTeYeyX8t/ojhSyx3XVAVdsGdKe1Y+yAywo
lVa7g5PnCvBfbXp1R/+l67TLqt5wCGlv+xyTfO+ZNNr1XFXMLB/dKvKbENYEetPY
TtX2dTUUV0z0REGBBvAM2N/UnqnKNTDTh7bKSscjeZMcqdW6yk2/wuMdgT4Q340P
KqoShrIln6uSi0uFPn3qB0iHb7bAh6kfjdD5Vc8xG+X9xGx/PQqKUTv15E0hUEa/
nJqNDvFYt5LpqRda9xkeEpzWkKkY16wCNN12rJRiuWdVG7sJSTVR+lBkF09vH+b8
hJcqYFnUuorpfZCmOPtDGR0FQCgDmVzhrF9ApdYVbYh6zjd66/ph1WSeux6fkSbq
+IQSDTstlTAL/riPGAVFLCGql6W8zWue8QU7A9XO1DYDG2oyaISlXo1Zwz9MguYg
Xcqwz0mnbB4h9ceR64sTOZeXprPH5NAaWfFVLeceTOy4RoW4saBX+wUJb8Yxuxvs
SYEvplHz2wch11cq3gDitJ2/gNRsOphcJWg1hFyBHLBGSmJPKsgOPh6pWsHWO8h9
`protect END_PROTECTED
