`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCGc2t840ZgTuEK15FfRpw0Tg3bQbWok1e8dlUDY/xQF8mBWQx/TfYQTJezEeIn0
Leq78pocTgC5rKiH18eeZAYEnsLNDzlTZBmngCl3lytNVInte4Kbz0QTUnJ5oi6v
aL2c0SY/7NLgg3aV/xo+Cxf9KKa9Xi5xgINal0DtaeX6t0k6cNIb8P8n9/6VTH9f
d0NPoRiGwq+pcnkR3qMRRNQSH3HvfikxTWqdZN+8nDucTk1wIA/vydHQ3j5SmH5a
2/GQv9KUMWqv5947wYVK2tAg3OuHe3qq5vG7ywdO2FiXY2B29g60ih3QggVEXWXL
AuzEsyFxIgdEbnGDMHrarBuVjyiWozrNJTuvkMuX9x+UPylP+YP1K+h52s3obR1C
26jI6x7nJrRC2MzE/W3NaQ/oTR09IgnmzW9609BkJ1c=
`protect END_PROTECTED
