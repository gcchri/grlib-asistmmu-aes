`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NZShRHpbzTY30V4oaP2jxM0B4lIKbihWL10K4+0sN9FTknwu3lRSelA7Rwbt+Mz
69ca8HNBYfTXUxieNsx1wQG/pNSFFzSiU3ktbGU0dno7FvzV3APb493Ffs+wxJUi
mYvvjKdQb3zvMvBfBxBRBSfRc3cgyGbe7fVpNvmjbuZHvbjzgNIcOFphPl3bWTCK
ZNnzOU+YkuwHji8f6h0W173gNRbqGJfl4OfUsTScu0G7bUqdjn2TVc92qELk/8Bd
j4FgXzX7lbIhZOmo8ZFSVt1Orc1UtTN0fNV2wy7uIZkW9/ZTOwn8QZ0GjkQL1Qj0
8kVchuR7+ziNWxLgNff+uy0iVVhyUfdcJcIDckka2jpRNpsrMAp3I1Pz9ga2bM1i
`protect END_PROTECTED
