`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Gaf+C4SfQEaPcHaxzzQPxpnhwofvzohL9BMyH0p5YzlQCB2oAi9EIMLauJuXV+P
scb7wRbq8MWT9MSRZgBitnxhXOVFaSq3kBG0WmRkfATj60WQ3OdsEImHCVVin03p
Wke5xDP1zoce98GEsP08dzCGCCqWenib4ckQgbuO760aQwoOijFZkaetggN1nSZW
oFV/+rmqeTEzBYmFM0priNSygC0lUvl2ZY6ssoZ8K8g65axMi97lKU4f46zAF2s7
4Ws5T9E+h5lrwA3enapOKXv+ASg3968msEp5X+M4UNTQkLBxQYAYAkXcZ5x8FjiS
UiPbId7hLkeX2Qy7JhW5iOB4khXn9SJxx2XhzuNaWaebBYjdhvEH/rnNkGQ0tyLx
AYblTTrXBBK/sTfq7VlYXaWwauqMhzGj20rxMYbRvls=
`protect END_PROTECTED
