`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YckHvyNA95yE68qjuZrudRhraCGVK4B6l8gZP82PLktNln+IUwI/n2Ecdsb09Mal
bjsXZ6hRUE8gfsWu3xP4YiOWB55J7mbPr+uJ0QzDnipHq0mP0y8ZXDQo4OuAsY2q
SW4I2H+qpmSPetyzDEJ5lotJECtllndjP3cVFK6FToxL/8ZJxPYZpGj/OU7xz8lq
4+5X/TDdyhtk0K3mY2CpAlOswl0iadZ3QyH/wJ80EzpqrrZbVXtTd7Vi3htWogfb
YNWYUMlc5lbnUDNgDKWF3XPbG2u2reocvW4yq7Bd3ZDTUZMrHf7hSwv+Ho1gb69g
wBHw6wDdFGczVELNnzXHuzlg1NtMiJxuxZpCLc463lInLeGO/zB+eVqE2jBHq1s9
puwW+zTkXCMKdk8V/2gMtdQeGHg1CtRlDr3iTxttGjN6AFm+OcxaAN+PvrjdzUr9
gB94tySnIh2uhoF+QNhIEUouifj2J3nalsFIccwCVptA+HP8po/roxkEc8vFPrDw
hu+3S7U1xlwYqzJ5kVoOH3onyrvr+RZc7FZCCNtQ7gx9asZDTO1Md7HEVAmkKQFO
1JL/jA9qnH78wxZQX/WVWezyRsVySQp7BgDyq4qqrcx/WZTd8yK54B1Ni+E3Opj1
ARFpmf59sO+xb7bepYIuZy7kaaeXrvbTbwX4kbRIZxpNlnsj0uxgrHTosWYd5hvi
9d2ssphBP8ehNhRWt7dZSFZKvJAXb/0DWXZJ2hg+IdEorpm50DF9779bjfW2COxW
B6YY5C9k9Q5dtXtehSMVwaHyGwnWqtSZJ1qQwAMHEn/mhKLFqvyxP4IJaxMj3aSx
PLwuae6gaggoCxCXqPW513l0dz2gWctoJmsOR+DZta4UfHcAw7+iFqsteWyttxyd
IQeJF4EOxYXnVN1W3WQuTVWGsAOz6rcISGNtRAOQDZIwMCEMQu2fNwj23N/7UknW
fAEwTsiBFMPkOOY9bpcVzc8x7CUDwCHWbkWcQlsQe3eXj9mow+GgyiRE2A4ZRi8D
6he+zuM1Zn0/83C8DQljGM4EflflMJlS4GwOqONuMep6LU51TQP8BupYPlz92/rv
jYAaQxPFHUSh7+ajeMI1ukK5KM0+hPiZXNMqSR6/jUhcSP87mYOhlfzCSmZ8Ut/z
9HPO48Dtx6fp3BLWgl2K/7zCNX1ojJnJ8ZnCZFLaha/kTZ1a8Cnk7EwysXgSLjG8
4yUSfNnFDDyNFYkUlC6O/TRIRfTs7QJ9AnyKyvRtyz6KJZSnNV5Mo3HnXPoiUj06
ReshjIVD1XP/89IxSoARd+xr7Yc6fLd7Ry7FRQBHnkF6o0zG1hYPGcfWYg28QG1P
72vdBxnxTV6k0S9rw7nGsIGktJSzfA5wdXys7f9rKm7TBk2tZAbQkZY3Dp29LCaH
sKZ/lZHPDK9XH5BSZBbXRqJVQuXFfDwH6+DOMmpUfnCDgpFGB+I9bAkrM5dnR53r
jZYD84ffoKWpYaj8gKZ7iJZ29KzwSmKrLH+VIzlS/peRLofU4fWHT1P3r/ch1+Xn
yfCzpKrbs8x0d18NXLrkc0R+Htm+B0Hf5yTAldpuFYB0IogxT78/QmuB9/rzYdGY
5ODiK6kgQhXAPTGuA3si+meDbZZIPllEzWa63VbhXlRZsZIZ/ZNOsOUWzlsQIEaT
UcL9NJEQ6vPXhAOt1CFS68nssYVddH923rq4hmPDUzrPz07JOvpoS3Mf4sO98uyJ
ki4yPjbF4dSobwoOSkyZxS5GlwRbRylapi7429Xl6m7+u2x6uo0wa0R7LDdPx2yd
F5C3VQexkkNy+WhqPcM5s8kv3po98fJGFWg+SeaKrr5pKrDbofWHZ8SwMJRf+Ilo
VHaNlDUMXeLh2bMjcCuTyQDpEbguldaoyti+nfaZHJthnIUA2psO83jGKEOHx6yf
TYIqnzqbvf/MhjzjdbRDZrTKJGeFRrBh1Ed2LBWGfiQQ8FtSzgroE1YzvEcl/qJ/
0hNKI9i7WBBePfFhntR7VdI2tnrhhCY640INhI2BcZDrPle34prWF2qp+hUaFnrh
s0aHp3IhJ+mKjvxL/cJSlrhMLSIuH1QTHZvrHhU5pYMP2xGGSx6mTIs2DHT6PfNt
SeKB1foAhZpx0ZMspoVPds+IpuBwDmKLOmY6JJsjZKzjhqnwvYdMrvLkaXA1hcy+
zH9Aq2LWO3mnKt6d15U5uqLkcxEbOq2RsvP5/ifD4Ab9xKBfOuENiQea+sIOoLJP
ALSfHr1h+t5A8S9qf3Tw7IpSah0S6GDm1hT/mnCHPOxpnJahCNBESmwmCgf98DLh
OBIRUXWX6wkNEUqnL1uRIlcxZAI1o9Rl/kG2QnVNvU7/Zt2DSl7XFNKGJrZNv4Rn
VVUEKFrlbbwUFvslHbW1m3+WbOLYhdBf89yxw/S2bhOvRS9L0AJW009jXU38+UGW
9W/44iraPyL5F7KvzVp+QFE6Upf641gnVBxENXZubcuwPLB/Y15XtHNrXN8dgZXP
C9iCTElwssm+HJfSGG0rDpCv5P7jgPvaoCEE2m31L5uiWIsnElYZXWYztEx26sj1
Sf7dgDtRvi5/xOIo/odmFnPVJ2wRb8xafXFMZVSldbc2g15iWmIFuvuSI44GXrdZ
CTXwjxxzOHk7IlwwakJlpWoQSekLpF5sGdusp0BGIP3ijgzN5i/syNuITD+PSVFG
6pTtT5oPjq5cQ8r8rWLvmoNpO2GtF9R2IIA2LkmmCGHUs6Jw30t8qikDl0OnMZN6
XVUmtOBC69f6/N6Mbi20GymlkKqvyWdZ6EgvVebulO+bXs+ewBxwAjuRRnmBeGQs
IGM5EMnRadBOG4tgUab7QvoBjZUgBWFkcCm90/XsaUGlGITXKzSBWiZvR4mQiEmh
1ywVJS/VnnSpiDoUdwOrmC5l8UMrAzKbm9sSqR7UqsZLTJ6IfTlaPtRPRqwXVpAO
glybi5IJ4WQfXQnnsIwxzxWO4s82k5H0+nGBTtz+tBp5lhrhFe0fklQ0Txqm1dRF
5/oWSSTR8JP1EELxpMNsgWmlmv6yWTTtEBOBLtVH1c5SvxNy4KDYZ5c6Yua0uMRS
MqraXK52UPeFna3Yp3PlZc1u4LmqVSVJfDEDGdrr/Af5g1KKw1J/2AoaOHh5giHB
G5zkroEkwKdeQrF8/z5t38gEk77ZWot+Zs+GP/tPbrNnayQX2ohb6telVBIdbp3R
m9rHarr2mopwC7sZcstavgCTvnFoXm2ElHwc4uxlHlKVzuWJ3WPH48Fy3xZQvd2b
vTiK1fyC4R6s3Xy+XifVBdYf1iB3ymgCl8cdrDEbm8TShM7d2CnBP1yu/0LL1ShM
61or7tzITfUIiUU3XQTuQXYooVzRxmvoQA/4My3bf6Y+/Zbs0678unpPUlL6BDu6
7/wihEYn2gLloFMdyTFO7J5tQH/54wrK4CeAbR/0NBXUJ9JqIb7fBEyiqpB53f6J
LFM9g7KC8fXef7dR3NYnEEadbXnboztinrff4+czhBZ/2nZpLaV20kwvwaM1mHv/
ZnD/V+3BRenkbsz6pILYthJXe6NmJ4smt3NgYlw4yP5Oop5gLGf/iPw3/hVwZhpn
uBXa0HJwD2ETVrwpsRJf/lDiTMRryudU/o6Y/hhq9a79dNN3qwln/pMMtCdYfxS0
KnrPDotWjluFOnASCfTIC/BXyMLr3fbmGglaNz+Tsf1txcmzrlQFNlM1ftjvv7eu
eGTNVg2LBp3sLrklUyJkxlLccM5q8y/mm7+lmJNZjOMgGdVAPmt5DP7FVdjxyp5J
4VjXGnHOPEKLCK3maBIg9n2XaUThQBv6ZIZp+dMx/iZUshQMqvA1SJ2RorEc4o3p
QEudhxl3ngAHq6KGrG9c2BD5pxXMyOIrzipyRZaaltGvnbazXYM5LxY20EI3l0yg
Fq7hQMVn3B5WEfjSCcwu1LUsIbRbwcGqJbmvyQhqeeonO1LmyhkTF2U1pxqC7wK4
drzL+t/+7Px6tz6kQbTNJ4q4zEygfFlzAOq7znlkT/z2UUYD1vc65a9hCtywW6kg
1oX5ZRzLwJSECgJ1dLqya16bZCBDK/oXzuqkSHjwxsfu4CQQ3032Ssk4UgMtM2da
ysqsWLBPXgZ7GY6bH6irJAE0omlcYMa9LlWy6NPtrF/smu9zQXtDo1u/34ko1lWJ
cXbNwOemRTPAwxBIoJprCxBYeMwSnF0+REvA1fQa7Do7YJSh90QDn39tptDVVbdH
zHwBR6KuUmyQz7evOcMJ8nBa8n9XaOj7OdFOqatY/jau1274K4ekALqcZfj6peHP
CNkt/VPwZEthdY5vs4av9rLJuNHhuiGbNxz02EjM2IjzpZfXJXLw5C3nh3TQrVbm
+ahOlLGUzH3qD62crgYYhjVN9BmI3trMzwdRseElidLiCev2dBo+4UnyT/1c5XUF
bBNn4U76kOePg6Qm+WM8vTGPzZVNK1e0QATKvLR/mPrBTd4+YYMiRwZx8NlNlTJc
oznxO7oUL/LinicrTRbZY6ITA98aLZaqnCphNwM/9btFbYA9V+aN8PFg1WMPMi9T
rOomlt1FYizOFME4tafEOusBtahdXVgA0XjKjh/JjvKpnVLT7+E2TjGIxnn78bZM
bikiuXT3I1ma2n4x66jIibJCkq4szXh5d3F572CesQ3cojSacuRvUUUN37HQGDDF
oOMgTJsjxWJKJEpNjpSOULyZ9xw0TLfx3c8KbL5CXcyKQRd2U1cjl9BR1JFC9L8p
rUtJUStRtAQURaGo6D/9qXknCpy4taA67aKl9tOHiRpNImK83DpuLEODugIwBX7B
P0JPK35bTM91ICFPsTGkDNG44/z5kswpJMrXxjN7nUlWVjPEyn41Ao/Dm/Vxzyae
5jGNj+/cQrLlQP5T/0whGAPP5LMKrw1CNqYdwPFEKZMqht9R645MvJqD6/FUqcZE
7jAOgF2PypLWftVIADQMbfbs8gLvNjZPDv+HzSfwmEkRyMsJufzJqvg4w9RyrF6z
aGfKcAArUUdk3L8AjH4vW8pkrtIiZOURfJ+ZPRNSBUjc1klNRxjS1xccADtudgrl
XSnGWVXgyi5Hp+TwkfbnyJQtENuk81FGlZKU+ShWGkO8lMljXHjXtQ4vPeEzomwU
4HDPAQCA1kcUOiM3b/SjxdGo5lkcDq5ay1Q5sHAvHq+CkTHbTTQJAAQTTSodhpO1
+cAnU02S2b07AVcnb1Q1CYUvAVOonDUUy67lazW4lmwpX/i9x61NQH8hZFoXrRGJ
vt3LC6cJ7xYZMDfXdObVS1q8bQI+bvfk8ldR9aJrfkGcfyp82fO/9w7zwYdzyo8N
dX6Bik0WTJUVFntoOA1OuEdJmYpo0DdvlTxtKSATo0tkTwfexI8mXAz1vAGoYFZx
nxu41Vwl04+sZWJuyM8UIX91wr6J+XNHsI97eiLrE0EEUH8cwBJe1Cr4AGQvnDnQ
C/n2TsWvnWlrBAYNZMMZaE9++UUyfnrraMGeEBq0WrYHTlYp49+bu0ZtYACv91Cp
mO9GcaSCJjPsIXaXdpHlmOVOkMB6VdOH1ASQsO7twUYUxNmI3265epYjkScJDbn6
+mbOAlJkxOY5QqWEnKrcft06wqhi44oH12wMVFN3BElQQaVTT/uD+Rs1zF6sORLe
qkf3jbWwyv863IldPmeMFh7KxsNbGbBAvKMw5qVsLy6yJ3E3Nwb9uj7wLNS6idb7
mVpkzhgit0e1o7+d1Y+QHqm9nH3jM6Y1DGYQtKOh/e930ZXMSkYCG/mcw8EAF5Ap
36RO2sffiY2htjrkW92J9EcbbQB59SNsSh+qOrrZASnvCFypdvYie4qQ6BqoKq2E
AZmKZFpmPOn7VhEIyqsz9nko1Bw9VP/CtmagDWU3PUJtrsKhLeJ2S5+9IVGeuqCV
opZWNRYuA6ZhGmdwTp4L91taEIyNsVNhBzDlIYuFbZTGlpkvswz1gHPEBUaaQpgu
GdroabmXGeSGVeAF/7sWlyRHKP8mBYm68KEXqKyn25U1B3izPoRJdrzYufTAs0Tw
9oyroZ8myiEbOrbuCmuPIu0sE8+bUi1aWv5dq+q4JxzTGRMzHjuFjqtvED+QPYdw
wn9cEOsAHse4gpJ5QZoUeonw5Dqmnn8/WM7Dm60fcPwQp1xCtGdKEEVXYBqfqhJZ
XqUXuycIDY4vWEWDDFanhNEO/coqZxfK/XBXTsXCI7+2rQ3ldhcMOKOIi2F08UQU
/Thkl3nc4T3AonScjXQ/9JSVOcTHizsForeAAMRSqsvqYOSuA6+/+zQfXqUnoPRz
dLYdkOnQ/6lCKHCU01mzlUKZhNkKj5J/R92L8DDW9W2jF/qmOUXcZijwo/D54u3S
sYCulc34TMCZZwE7Efg8WpHq1rJtGLK6XKeuP/d0QKGN2DaYGCdUFpJlUHqNhBUU
zRFz83xMMdraiMtgAUIOhfjqPi3uOBESDIkGDHo+laiR2ZEgaW1N+ODwHcgnLj2O
2SwnhYsTydFsnCAdXsBhQld4MzVkmgcqj3DoPBr+hz09fO++taGYz9WcGVKrsPe5
daImook0Ao2dph/5vDnQOxJCnTDKcaCnhg3n7gmArdJgwqH9+ymrFwokRTYzBRBH
xQHq1R/OZibdnk98lZxcJ5ZYV6+SbvQqy034qWNCd1DA2+t3Fq+RdZSAT1El3PnU
MH0Xjx6pxaoCf0tB6DtZ1bhniz+ulxLFAH9Bvw/tSZtPmqLLhVd/yxLntbuR5d5V
wN2WZkwMJvVeq53+0jNJX2sXYEqa5Zl3jNLRUZVWs9TuaGBsLbBR6IZx9aefYQT/
HjRx5Q19kMwqqKV6DTx8swDVwRYEGzcoCXRHu8TiDa4lQY6++KFgY3thmBf8PJqD
T1+nSRilUStSIax7TG35OuUM43cnVFKARTps+f9c8w6cENZmYifndbkAz/wDqmmO
/JaRDp+e4MvsflAekl1BczI+J9xuUQskDzrLBm4DNRxPGyBgTyG9d4wZbSzioA4L
GbNzbaaumgYRftVxdysF5hzY2Bvij4sHToh/wx/J3s0e6DUV3ITcGuUerYkMGutL
O732EX8wHHL6xfpQZ8XXIMKTfdnUQM6A2QCBhb1NX66YRbeldie1oaRxxf/7MPuH
2fPgonV9DXzWYYMIM1Shxh27+D+oWbzdFICWEVjBmbEPk6wjxJ5HQDQh/GtYKS9z
8T7zce9sSHJm8ftzRGgEFZ3ErOBszmB1kpBkMx8qQaDKUU554TWEC7qnINaSakuf
IemHT5d6PRPIuU1VYoF+L/hL5JjSXNi0OmDwERTsK6onk79q4xAObSFr+uy0zC4v
w7Tiig07UiTQTNUjM8X2IO4GbQQGf6STAdgafXxKft71hief+4P78T8H/8jvG5o2
niJ+UF4VrwWX4Cf420BKzBGmO83wr9Z2XEUx0tRj9bdoENqiEeZD6loX9SiXZmVk
1FRI05TCI3O3/NsgGsYhLuSGp7aW9/vZyu3238IQbBK6HVv1+Ezf+6IPRxOhzEyN
/PuS2wY4NrqGtZmxQlJ7etTVJJ1To95/G9HNekUj/1A/Ml1BQr4OAUFescC+KEza
kO/TPPQ33/eFMQFhnn8kxIxqXBf/hSP2dT2zonDuMACUiXaU9gPNYCPLqXCARQsn
hYdb1wNFenB8xo168htSEfFIGcCAqCv7nnVxhI68p+i6ZMRYGg7ex2eu8UptMT/4
aWM9NBhV5NvJOSu7crIhQRdU0fIUg5EIA9yhzuCI9+E/FJgGM4ruLgr19GSxvrGG
7uRaoZ5U+hbJJw55No3mrkqXbyemIZLruM1WdwbRwww5nixapyETGr5qIvTsDM+y
Mm6Jq3CX4KGp5iKJjc5bmhTUA+JTDey+WE0xt1lSdMxDQfYxV10ijDX3ksThuNoL
21vsCoIgynuCqBw6l04KUURrhiFj+wO6Iou2XD5V/J6IoAAAHZKi5e1S7XoWeBAU
ZxirqLhaRzkxR0AmKW85tcxENw0BawrrUTt67z0cX1+mhH7XMr8o/d4wIywu5ZMW
4LaO4vDFQe7x50igQRYM+6CNMCLtCa3y/OrY+5tUigcYPLmWBJeGbjFGOfc1VMXU
0cNCeSxTYuGGWRoLn1L4kIIomNAopTImmNwdRhTvgTVyliM61niQ5gBaTJb7IFTs
dOWZPd7Elu7mBWC1VkZalybiFiAC/XBJkgEPP9T6FA0o80yMTXxcuMf4atlG/jl3
pLRpOHTby/GdpT2rDoEcKr2QwWKikwmKT4nOexatEVGnL09xNnMI6mInHslYCOYe
Z5pkEcbSvHd0mMiqdavmO+6HVIbFYNGVdGHVwx7tZphMp5hXu8iggi+xxZ9QLqV1
V4voXQ1B6WvYysltSvIbCf8jseb2ttq2MA/zCFd5ER7f5Slf/FjD8z+i/tfRdWWc
9tWyxNTIHmqTlb+Z7MOEReNXzeb3inwupy7VL8LjUS1Se21cjEgkO7FjzBgZH4sl
selHdmuBpKkQO46QsMq6rf+8qX8U/RejprmoiisNRXjnIMCT0ZW1x0Vt0yAg9I+a
m1NeFAmyoxI4ApabrgQt6T5jsvgAPgKJt0kGf/+oS1bz+KKxW93EoqY7itiRiUkW
zaD+45Sesxq3//m5V0yFm3jOlsYSVdg+xqgrVvCYJO6GQSuGOnXrXZqTUtKj+4oX
iRQsV5IsKRNkr5q4zn9uueMDiqMQxSCvmbGY6KzUiQLUyHZPvhbQUyvow10e1xIF
XLIUlc7rYMmLbNC9Tg02PYtjerq1LxFlwKmFW9DyVhdHgD/9dQd1rNPrcPHqTJ2h
haBq6uNVvHsIZACNxM3oiHLhEQAPHf4WzAUppfgrx155VhFGOXTfZ4EoU/ttb/8B
MhvOaDVDECFzx4qrwHFLZMwh9ltdiREmtPbt5xbmLuw5MYBeqliKkK5t/Rl3C01Y
tBH5IP/APO2Df4NfuSsO1E2GUNolWmq1cs2LdVXfpFBFgsjZ8Brd/LCNgB3f3+K2
qpP1ICoWuIDb6h7fsRRVcYg61BI5sERm8xpMm+WSevmoaN2c4UTMNT5UB8MAh4em
k7Rw+0vx4xF5/QAyD3tDIRur3I5EnLUcgmqb3RCB29EYTv99mlLN7U4piKUxL0vc
65E5+kV/6RbKKLHuc4oatSfaKU6PDrVdoizIPtCpny6IwV1OSvZd9OlLEQpT0A1x
nCm4nqKrTSR1MbHRUtz62kmKn9JBrPK5UqYrsUTWosh8JhyfmDLt4kj9wdwr0rop
Aaun0hlfdzaf6WqmPnPevwRr4Kjfd9qu8y7vUfAcsIeU2/KXmw+YPVge6jpVGL7h
C+KRr4Pa9Cw79K+J0xDT64XShPD3Hg2GiIihKHVTVKLYbv24idwlvqhZpRXuVkdi
W2XxQ/plZ4MQrcXDFlu/geJqtX6cVbilAqXFgDg5APefOpnwaZbn68nqyJVUvr+Y
fXJVz6ISUpA/ugR86CSwIGlq0TSujgduXEiLxqIyjGAkc7tcYz1lncpbq6GonBdL
8KFr/TyKFKd9I4xz8q0nw7Ykj7n/x2LEOxV1UuTLGobbkEawYRxdcqTTfb5tLIux
gLuJQJJSV0h9/JZTbQ8CcmuHK/HGvvtE9PNf0xk5rzFpsX+64z7mi/Fzd0ik9Zoy
2BCVcAB7GfG8M7MfC8hg06lfR5XSA/pRFsM1zRdsPsSnqWgi3ZC4kwXgAaIQCDxh
WhbIYLccJqXv16GBQmJeX8PUovKye6iKQyANkbQuYjBfZqrtMMl7G1liWXsTucvo
PmSgUnwMMmT/qN25xsMHXvun5T3V87nOyJ2U/P2PTMTBuVQPK2yLmWxd2+aNf2Oo
KShBQDFr1g4JHqSHT4Zz4B2URN5ak4lMqxCc3Szb2BZFmTlpT1CWMtxFcNttKg7D
d6DDOdkkU8j2jNyQfpSS0P06c9STKqr08jkoE2PoLF/oH5ol2FT8Ofkve6GHSMbH
88hZHv5w7JUyA6X5QFJLtT6XP2wJ0b+zZbAyYZP2WzqltPtfnUb/JdK+LPoM2Qb9
dto2UQvBxlMPnyxPtzQs/UOwm2ecmLONkYkFVSccroAmv9/UGdtxVXkOHrlNYlgD
HI/qbZkWPdRIlZOnjsdHnxJ/ctPQ2j1mrN0W2BCYHAfmlty6Y6CO6dChnj2RoK/n
wAfuCPOs43RDj38gmCd7Nk2seAryPpGrdcTPbg+uRdFi9Ppac/Boftw3nTC2wsJj
DYr0+6dXcWDe+GH86RMq83KpUTWlbeqdyo7GThntwc+LBwAyrItaz4JO+OV9QQtW
eysr9W1EhFLXHnATbdCiGs1f9vlyqD+QIBdae5+iBd8mdKpYn8jgus9doNr5VFIC
cdFqKN7hdr7q+hq+rMGXbnN+ceqa9uurvISTv7hG0Zk8PXUkLn/zBOxvYNConaeL
dpnHc9q5iRf1gZWh+114oWpIGktG9gmL8kURw2e/tL2fw1AL1z+eVH0qSVjya+UQ
g0lnKqmCZgwJvAh1DjbfcdxKEZFe7mOzUS9i1VBHwfkGn0iUkgbhJ3VRUZ5RiyGG
BGPCXegg5aG2zKcfc0emUzFvy4kGWSfU7EPpAVmGFH5OCVXZcS66HWxbBq5Pt6Sy
ohU6IF4Ge1NHnbMxa2XPjCGzq5oSEVCcMrCosdqUt3TI6618d/7CymQg8UCFkNvL
+U/dILQ8jZxc/hlVwI4mNYumfnXg/sb9BVyWg0vbQrTw75cHs7gRm+oSuEC4K1V9
UQjXyKn8XdVJD7Dk3c7zWM/6iaf9O8S9fnjpdjxke1XgGrzyJnTBPtdtbN0vkfFE
jO1eUiieQ4eDK3U0mSebPV4GP/yUymRENAkpz3iA2TryB/gi+8v0Cgtj7Q+wa4tC
kT18f35QQVAaQuQESxvCrwRiDBc7AqWRiPfytLgt53smk2a6iiFUYfyiLt0pwNOF
GvnhhURkB9mIEClyjETrEHzZ0takPRKcl17xGHck6+iga3PwCsmAQnyWT+CtaxNL
Awz1CSfIww5gcUjaP57l8sX8tqGdyDEGiXF7wrMYJtLuZjSNftQxYHbZG/O3evS4
d7N6T2t6PxoBrc8AMYsRHKHBBYCEvGpvMDjYbZ4djCGuxGfvNJUnH4p6Yc7CGi4s
mpcvchBdqeoFBB43gcG9w/GSE6fYK5T9/46rqgrzxB4LgjblWq33ll4CnOFKicYc
mc+8ZPHELv8zRaaWRakIGcO0hgNfWR+YTba6YwOhE8vD85xooNNcsWUD5OYRf5bO
b/zikKUm74AbPena6tAxBIiUVbXzGqU92008Fxhb1fxF4avDaxMaYPK9lpR1mp8m
5ib+TuZzanW0OGAuvMMr+/CJrCdkMnsXsAzavngN86UOMddWaD0+TBy4IHvpgw/J
ZEirlr3QppKFaFYPTBsR6I0DGezxuyNTgm8MhUpiEpocB3r3V4UDkx8+op2kVbfy
AFQwKghzb/Ufx5i66IAe0w3RNT4Q/WdAE7Hj8UYwefr/fifloqhwMMC1jQj5r1P3
ggSKe2Ehyx9d4iP3Fii2pUOnU9MvnonFofGeLqroCEMIPT+TRJoHmXx4S1d9eFU2
vr5sMwtGfwq41ygv3yvTXBbHgY4d0CZ3Z3NYRuaY0IyQszeAqAYCY73TtMr5bvLn
yGZdaxmXtgeRPk/vbp3YrGMGN0JBYysRxg6rIQEv12Pao7JThvVCBSqcTyKq+5Zj
zh+YcDHsa3hYzHIAYecS8ogcSubMby7mHrRaQAROdj3uL8U2g4lKIZlzrKTslv+8
sb5euJL6ByvpblnWZW/LlexR26XXOTuPT8Hg2A0te0KK0LiFbEvIiK6SAuJ9a9r6
95vR+qYxZ5JYCm3mF0mBRLRV0IDyfRQIUyOTHbg7WFYjXjcQ2PuU8q/V32RTYhd9
S5hvpEFpntTHteQE+/r6oeim1ieoot6/dtpYXWxs71KVTWlrXqTg2bv3X7LPO5K6
bSAgFtDxb5Y9bJ7UvofQyyMvEBEOcTjCbKfjAX9I0LYsZrAUqhX/FVdCt7R9CJtk
suSIGo1x53ij9+wGdsofBWNHRLrLhTxeX6IqwL41BVxhXQIbxDQNHmAcWfDjI4XY
wuqpy+qYDw83zztIEMX2vI/F8veaxoYiAt1eaRO4wXzmhNOEd1CvFScwVPrc7ds6
BLke126AtR8hRKZ1QJMf4MZT4n7gaAD7T3Qv/r4qia/yU+JA4zqSYBBu9SUBBZQ0
JYS8PAShgASyIoqCnAOHBJMGfY+TmVDiyf3wCrmqLfCqhJBKFcqwJrZGAxnhxGx5
cuFbywhiSObcQ0so4JoFRB0r/TXeA6DbM6K8ktXjszrVWxzAFVeYYzfR4TR52gVe
rZ/60zQ5D7nxUU64yQ0XnGRCWVEgHzv3FkT9uyUWV2OfB5zUuJjY0uJrklMv/3qE
/+ksYhQpm7f59DuKNC34Zw2XXf2h8R2Bw+m/BlbSbAG8KlX4qm9GRMZFIg3jro9J
yjMcV9+fzEwhXPv6jf+kT07uNtnEpoRJoy/mLYVZAtzN6j6lVsokYASbgIgAL4J8
DdXFI7Fz3kS4MEJ6xli923GsBPbW2BREWxlC+yL0B5qPFmYHnnubQt3GkNg/8F/G
ipSgkPUB7sEnhD2swsYEqmo9PhRZoXmpVSH6jtZq0tssNNkQ/FOVv6Disbr8wmYV
8ARQLCmc5j63tw92GDWsWbmljWwqgdKxuBcHZcBvbcnBbMx176VhT+XuuxbaPYsu
JTRH4EugS9DXevG+XufMzXpGoRh4Qqb2BDr/REWfuvPzW4NSyP2kAoKNURPABGlR
kILVUHoFsZLdFgVOzb6T8ka/X2rz1doLLaUFbjMl1mwuYTe9Fo2PzLLt6zZtHbop
0OIsw6ddMiEaEFJmtrefd1Piaseqce6BgV5YX2edd0PFNQUgtpvQzjDHAm3NpVpz
8O0lkiaoJsibMwX1w0GE7UoOczCPg9SbWUBmxQyQBQWRErJc0d0e9c/5rJVucYDD
HCVbKdmIa6JP73Ng+G5J/UDyMH0ecwYtEbS7VWinFl8YdFPW9+HaX8CGRajTYLwm
V/3K3cUeWn6+QD7+kRdfYh4Pl30HBXtKvZJMn+hkoTbN/rA7sVtUr6/KnARRsqA8
JcgqPfvwfHSgcRJGRwV8UDz8jepKXhHsKauzEG2M9S0VzGoRTX76yHMx9MS1rsDt
ze3DUo7rGCjGFUCCuOMuZ6PKErlaggsH3RdN4YoDWTw6LoaoXXHWQkFlasG/nVnl
WepVwu2GIhi/Q3Mumq40wyEY09ACwegFxc20mj3q7fE4Rx1DoyljMiI/9pIxtnb+
V8+jJ339ZXXSL6RgPZCd7FCSgzGqXE8CYrqA43ZHz1eT+pArhQG4HnYTuAGR88FP
V44s+WA0tTmoDmFBQ03vTmnd8AZ8n7ar9iXIH+q3PDdjy7LQdFtN0zZ8yDDa+EV+
trH4qB+/0fp1gRvi92y+aqsIBe9ZpaySPTm4+HcB3cwYHywxqJ8H9ruEmNwiJujH
iVzT8AVrp0eNwBAwoMHAWwB+r1ynNY/JyH4urRcUa10KJxpscDon3EYRiFiyvI2l
Zbn7Cwh1HnRN5gEZiCeLpbYBARQgKREo2BaMTNqlBGxrJLS+BPyPpR/dw6SEaT3P
c4GO6LPp+p5m0QjJUFqcTpoSNWOjBlfYuMUjtuQVVgXdk7A4NCg2Tp3iU9Z2lpET
shX2PwumV2uGJqoPVmcELbt5/GRxFYkVVciQinaQ3LqJQIUiDTHPXil0LKjnu06Q
z8wg0X0qs5YJXkEdtYfSxpfFYC1ZlKT+vrtHohMb9+KaF95VabotQppTryeoOdIs
vPBTIl2VCyapF8WCVM5zVSXzq2TRtR82H0uL1H/y2rFFnMvhYtMbUnHpVz6qndJk
O8A5qZkD8jJkyyIuz+g7nMfQw8nhDldwcXRIKXN+c3mWEXF5IRPvN+vMpQAVW9D3
jqDfyeCovjKX5eFsuJ7lzkSEptR2mz6fv0FcUx3jC9+sDqT21f5VleLkLunh64nI
x5i0JWqWcMzx/J7JlTpanM9lunI49gRYaVB6ws6j5BZqzF7ldTmfUszihKhj2zCv
CH1p9JvN0LbjthbBcRSmtQd2z8vjXyxYhqBe4VpX1Ykr5cCztkr6w5JIWllpide4
EzTCEkK0XIh5htPv861sfd2DmXT1R0I9QphpmY81QqYdRpYwlSukGXddXNDHenCB
oLu1ZPPU1G7/A6T+5vrEakzKrb6pxltQJtWQvTmWUKGcSOJ67RLAyiwBaKFbKOmg
m23XcYwSD90rC/WGTJCQPc26ym1ztW96m20cmzmdK9pQizB8REDoVR5u970+I2Hd
UlY7Mgc5e+dDSV80vjxK4BfCUkJrIsGRf8zCrV+oUei3Hqf/9V0qjujz1lVQ31NT
QwwEg2waOzSPXH8595KFMPTkRtbykdmO/zCTHWErlcHJ5IxqC95GJGfvo+hOb7eq
KXEB7Nbmr5W6mH+dXFbf8URNidetV8TsjtFJyLjkJ3jLkXWpJ9kHB2eVztr0ULhC
0ravhTM4+Ld1rD5a+Jz7CXUKGBziq8SlL4HkzgdjZjhEayekCWHulIUXQGbZ6iLR
vVBD8nliPseQz5LDgn2zgU+VvJrPAOnCZM2KSj0dbsWmq7tlgO3Ya3U1UGZ2wS51
lwztEufARi3QciiUXVKe5a5EYBjv6tWYB10DN8LPt3JWtxTA9oPkrZFvvm6XHfLi
sZv3fjETZmA4xRyGSaJzRUDPjA2EOrGyqjKIt9YIFRNp++aaaDB3kPaSl81qkZ8u
ph+XI8u9GOxbwKw52Aaw86o96TttwdAiATDDKZ/+fXt0TFF3LQlM+rjGLjimg9eR
LldlUbGYU8S6/BbGwkI+dp+pw8YEZHZTFTflDkswlTvKaZhlUah4F2ONt9+CXCl9
nBzgzbIr802kFia78qrQsjRrWa0tuaeevLSAsjVy2r2GOoFP7cvqrqkJpwFFyuZc
el9WoZCko9sLOb4DSWGdU+mcJnkxSRxaENVTU+OpjvH9BmpABVkE3OJ+ooX7ZHt+
13HVzYwIEkT81G1QfUXPZCjt58NfF1F0t8rEpy1AON5kZGilpdNa7zpWTk691y2u
tCU5YZaXAuisnPUvYn5+1wPuBapbv6eGIQqvi4ndvtjgKnjelxE7puLjkT0h7zd4
oYN111Yi8InERWGk84ukDjxcPBFnykZXSh77J7KoWWOWVCCnlFQIbgLh7Z9sdC78
6Rz5MUIZPn2Aqw+eIkHdJEgn+ov8n+I+Df1g9i4QngeDpuuBf+6TpOmYeLv3i1if
UnG6KF6BWrJJZf4yj9V1orHUfTdlYNCJs/bDC4JKe9eeHDDdVaBkQHkI4ubX9Mrw
bPno4+0QtuLt6TIC//X75G1kG5ggdK18m74jlfy174DZwql2Rt2XRUfXNdx24Ldi
53ar5MEV9MvZ7GOYwrfOC6bxZiV8hr8Lws3YafzkdqWV3W7D07MivL+JBRm4Cd0R
V83am/cNURnB3KXNe0vGpG6Ka1hBYNcEuAkwV6zwMPkVkNbYDRIHl4wDTzX1rizH
KMAD/alrZFuJR2Bu012LDRzyUWO/np6owvA8JZylbGC0u6T84OY6Bu0O0DQR7W1k
z5xgxY3k+yZFAlMDtzf+jX05U6BJUd8Mu9WQJXG5bxIBp8/bj3XNNBZejFTndZRw
yz5EFEJDyu7cJMsOWdXn3C+vAtw+puHa5ecOd07czuOR8ZJkaYkJZjwYaiqGfoiL
g3ujWfS7OcesXH7FYsVpcsjyXK+PrnY+nsnqVtuYsAtmAF8YAPwa87Ti7NTf/cNT
qrjpPU4eOKChYsfiSS3MY0eOsB62QocEiYFid5Sf33jGgAv993RAoIF/DHA0nCrx
y/fNnfGTU0styrD2oH2fBCxnSQ13Qa7q8NIvu3nkr0v2hacO07wvI+9JSvF/WgYc
++Qby9Kf8QNe7GcJw4HrAF1C6e2CyuhzS9alALBzZWt2dkxI8k7Z1f6ejCAg/ITg
Gl0gNbTkoaIeNJ0uaktJ8UE0gMnzo1Y2YyxXNEvnJHklmoRxSbq1Lp/Q116x8WNA
Ti3ncFZoo4n5j1e9SQrzYcfZ81srGN7lS6swVtBg0WZu4Q8U/m1Txjx9tWgSMmAR
dEWdhMjh0GC4BeXaab7BG6PTUbduSu0QC3gZCnGdtHdKDBpXCLsFgqGc+5g+/cvo
Fj1tPqtbe3Gc4QvznZIVP7kfTYPvCRTaqdacxyDSIOixrni0o2cx0jnRN5USjBhW
+BQ9z2oY6k5ps1+28XaFDuIFL0CN0QoFbQfgY15WJ7hN+rvpdScGaRQwTAEMu2Ma
W9i5eXYGrUH3LNpPDiHRuGl74/Zs8BthZmQu4sbirYlOMc+nzVQNpro3cREWliZt
kWtX+XrnF/bjsA/SjWaifsUNzS75es1JVp49Hk2oYjLJsLjpWyVQm89PO5D8Zv0k
HfnXNPp67sUJry2tkZ51PohADonBUpfmR+VhS1Q3O9yFqTb0JLtjiB4HM42+YpHW
qBREyobrraOPc9p6120uUgkBm3ZT1QwUKRp1VB2+LaEkqjBeJMxaKEVLJhhm1p6P
gMkwGkEy/w2EmH5cjKqmK1DBhj/6y/cZH16rm2zkPVsGQTWNyrmxtcBf3TbJlbDZ
vrGzWiYz0RuMEz8MrcxB69CjmqhHGBWF7og6d/w7oWCA9PO7pOpgbEViITntGcC3
NwmsUj6brD9p2vZjYfQR4Vb0bvYCJu4e7fp5bGwvrNkPG1MSVCSoSzeU6km2EkOD
3ldvv9Shhrg/cLYylc9Kclrnlu6Ucv2eygAP1GjMABpBreXnd3c1BGjBPugijuhU
ye1SEqGCIKdXPtcVY40sofQIwCw0iAoAS4xHfHta9h7NvjeGkG9cVrUJoHDUP5/j
OeZMy8MT5T0tV85ElqGAY1s7nDUgtcnT9bS84yehEXWp2KmY7Mv+NFBCmVZRxSjo
G/Q7RekGEmXhl6wpBasKkGGkghkM/gy5+7RCK0i8Qpo00L43ODTthGop6au0F7WB
LiJcOyFDD0VEKu+eWDQZowj5zJJ6AAPCmvht+d6ghFnYen49Csh3SqzvOCUNd/h0
SLdyUcGrN+D3GRHA4C0qRJDltK8bCXhIusi6ZX2tODhXiKQNWbElc5UQrXb3AQ66
6AY6eyjxW6Cn8HBqwUjg9hsPw1pvKYKo7TtSZuSoNF+gj3F3O3jh2lkX/kLJ9Ftp
LYBgu9X4l1B2yAnoVRPL3Whh9Bkv2kfZ7ipWyVo97O/t+Sa1b72Qvc4jD+zqdxhQ
HbrSV15lcgsUAQhgzoMzhpsnQnH8kLi5LS77nBl1tgw7jLIZD0gh4cVC19Ampco+
q7sXB1uNUVTOH1idBuuvmTiIProEOcxqxvQ5o/lJ+P4m/sxAbhuHrl1bzkXOUMhG
ZCq6nIzsVgNUq4tfHCiQZNn89jIgsqOWgDVYHB9gdLy4muZyUry2JgCE1nzF0nZI
C1eHMp1MpBzW9IGczydCbA/aWkWVamPLAQIBv8ZvmKqvp3F8QHa90eLNcWWFomER
RvNbS9gOi+L9dG099mWc/CVFhWh4xsvP3E5DrhnSrReiJk5xb/hFS3eqT2uXyLV2
JXKWhzMebXCf2IPBE/7uLqKBd57VCq1pw7XvLbYu3iAict3J6OKgfMQYSs9whNCV
WVnGdDIJNnB4jOkFvOemdFixzNo18jemh5kfkiIVP2s/h4XsNAXrOAjR7qhcuoA1
zImaaU7t4SOpg8Vg8ZZ2uCGyjKDiV6rSH2MnYzGBQK2MSjKiBpQTC3ALp/4O0K+I
a8ZDsrhP15YUyMIcz225e19FHc5PdGtsACkndNt3KEF2AYkRQnsphLbcg3BQBi0b
Myf6snvYEDjMoU4b+s4qIkUzo9ZmsyqE5RE8rDAeEaKcXHjgugPRckyxTooOc6xK
Ui16XakKIy5Qe5W1lwZxYPXKVDq+Og1vaFyr2A/OnBQOrjgFIU8QcDGQo+/dyJgI
HTi0dP0+HvHIy1G3D5MuHUvKYpJOfFbwW/YLdR9pcP7hN7XkcebV5g5AZRgHyw/2
zdk/HaLpGY8e804Tm+XQS8p2uwnIL7iZbiMTauACt1lTBZyKLf6DT9SLumq7FbYY
6soMrfxYa9Wl1bmtOWqZlM9D6hJdQYJBIkYJUwUDFkO7Y33glUO/L2t5+zSuGNfM
pkArNpl6RSMbTrH7LixU10rZDO2FlV1rDccLJTMLLaajm7yeWKr3T78Q5+kPJD84
IiOCev6Vga1N7E3F5E23Bdzwl6xARC0GNIzkQQ1aI1+VcuWFMnIBfFP0amrTeU8R
xazcg3qQNfa7uEVKNr38BQfb0EpnIgF9xkCGILN7AWQgtn3b/D6DAxMQLFH9QXCA
ScRQ5wHsFZr30R+RUpFbAjYrt26BK40G72Q57UQV5zDPaDQPPAlX9Yw9CA7mpze8
O6Gebqp/EeiM7V+sldlOMgcPCu6zCC05VQPAEnKlq85ALq5XZqX5IMHaHUgP7+Cr
oF8HxrY5O6/NDYTqv0kceJKDI5ZiIV498g5YVqzO0QHKhG2u2vEzL8Qw5tdoKpb3
gWJ4bsN0LXywu8GnNAUiP35Dy6A3koNuxnMFJNOqwgvvpEQparHzqAtwrW4Q5NfX
YLf0qSplW2wbRNJjJn52wOhMJccN2BaoAkrGNZVfga9EiTE3r2jKOkIx6ggcB6/i
wa9gjctqjJKxX9rfNrB1Z87bZgRYAHeqp+PwkneAV1NbKBenY6JoGEAKAWuFxk9s
kef3OmyECXyfheEMi+MEbWWkJkx5I46qruHzNzd9+c7vFthkJxqtlnsheqPPwCcX
Q1+LN/7mrhiRge5W5N7UVSPxl3tEJbG5TcJPZ7V2xQIHLGwSLSmP+gfyxja5ML1u
aO9h1O5JbkIeF4WlvrmcaakOI0HgWH5LMb8w/Amp8k6go9lZ8+MjH+7MudJ9NHQo
zD+0bJ9QVgrn+KQ9m5vNQMhtuPeBD+7ys+rkqAl9qiGJke97CfHlIdao71OOsrfK
pME4uWEhR+MUNoe0Rnpn1IRCBlMGj0GylWnzRNHF6Irlhm09l9gz71F7BTcxElqq
M+wZ+PnX03EaS6NZszrr/kP3v0itKD29pgK2JsRlGHOc+arBMxmri8B0zJMNwg3z
bvXoecelx8kzYOTBBMl3LUnQI2c0i9g5jrXztYcuv9V2ctseaYrwZJCv+QIWqaiT
ztt6KLsC3rB2iRfIfobE9FWjaiYThUDJ59LPimZIz26A0rYZjg+Zwx9qgDs5xqBn
1FYtk0DBFRl4vb/xD+e9DC17rFWNDl706piTcYUh+/Y5XWZwFcuNEbUsvL2gm7uN
VGek9knk0H+JbXs41R27uKqzy5EX5fd79imPVgh9PE9E58R5HKmWCwEpLL82r/sm
fhTjFpSCzdfd1APi86Y7rs9vG77T8RZ8A9oCwsjZtNzmRZnEB757JqH0AxpVgvIn
B4yjfMCG9m/msrnyO3rxvbR04yve3WcEOiwAYo8QMcz4VgWpJPHv/UV4JxQLQXO7
C6M0CMpRoj1QXpJx/LMAtTjCIJW7JYAiSYHKKag2ImDoqqHRi+BL9TjxEFjJOsp4
xTdTrt+b2tj5y2STJErSNiDeSFAcBxshgjMX6C1RolHm+Hc1KFDxcv7O3lx66x7Q
zf1PQ6BJBPN9L53iB2PgTcL2CzbzK9h6IgvMdwkrZ+3ETsNYBEymedoHL5emKQcR
wAFDPSkFyAanvnwktFwNZGyeP75M+awGpuayLNKaChrzz293Nz9tn5QfA6+ZdqeY
RMk/G3ahKU/31qY9tBEga0mR4Ca9ON3N6zFPU+DMdm+qvf0kP0xs1RdOas3Kx0rH
UN1swBemenA5jr5O3WkyF/UbfXpTNzlk3irXsCTwIsCdIXdtvRuSx5CaIVqwEoZR
KShJkjYOBzvFBT6LSro2G0nx6+TYwIQHRQdStmA76D367fVHZRkxeDqPwcAZ5MKK
mQq8XKO1h64WszOV8/vsvQuJKc498f//jmkhtJGGZUtsHZsOiGfDO7xe716Yq5e4
ofBoQcL2rHktA+phW1euzomEOIjQN8yYM80msxXa8PcqJTmvra0CrCYa+iyzouEq
DOCNlV5D3DTEVQp/ca5/OfQiqtc3fJmJh/dMsQLoPfATx2LKHNhg1RXO596nmQ1S
BYi4GK8L+llxS1mzpktg+jATIQ/MmDVIYhnEaaAJmwfCc+aRdOwVRJenOmnJKqfe
GYiUpET2EOGkiQIgVXwz7AJzLo39kysf46oxSUAS3wogEoPKnmG1KB9zENrFDygA
8ASasuDE00P+UAJwCGQR0TgMFf/MIHP1wu4tB7RmHATVvTIuntmQp+MO2NMaQfsw
F9wGIVwOU/eK4XohHKhG2m8gqlYusf2LAojhSYNVe3An4I42X1uuYfTI6pnu9dne
v2CI9N0aw0pLxIyVjvJfiZbowc++KaWpMutYoYHRL40yB7i5bsJOeNxw9e5UuTI6
rGs1v7MVum4CXDyxvYenn8cL6nL78BQp+t1Lmk04gSPk3VSs7yB3D4TROYiw/Bnt
NzMPwtV0nKYnlmpcU4sGXwiO52grNSeOch43Hl6yVFyTdXa6F1uuHBXm25I6dYb6
PpzKneJ6sfN1uUumQ6LN16L1l7NBzR6cTxP8p6aZQyCuk7p1M4g6L1jCMno96txi
C4GWyaKFD2sv4VWZ1ZXX9WlELTG6xnrT978ZQ7ZNvE2JDPrIR4lVzDFKA8zPyaAc
Wc4ChMtY3nI5JrXFvLniFMr/gL2cabwtq6OBRyCh8i4K0pKu9AXOY/XlSQGGLLxA
3Nxj1Hr8uJn1i6HuWsfDhDsNtAf8ZjBe25858oAGPgxRh2jW7OgztjxY9wNIK0Un
0+itQn3Qq7y05JWuGaDZzsetogMd9Artrs1gTavu/87hfebWuwNA1I9lyJAsflpl
6SyPa4fG9nOgLnJ6nLa2lgPD1smT+vWM3rKWYZO4Gw4hanaX7igBDL8WowJj8NZm
IvaTpTDwvCYpUNjom6gd3FV1C6MbKApjSajBeObOJHoBrpHTtkXAD21ICaNGPMrZ
hXOjhO0cZ3I6bb6HHdKXrusW6ejMh4bDJKZIlxrrk2d/t7shqWiM/xYP0m2E2/ow
ghbm116lxwfnu+GDzF2r7xVfYuhM+yXheXX1I2kngoodWyWv/6+o8/5SJHbSXWT7
tcGLuMieg+IdfvitbmjIuzRUwNTwQYY+apYGOigq3teOo0V5lIfmBeOCUg9iUcBf
EYLBjofp8YgOaqPeQIcQaChqH4I6CTok+EQ2Jq4pFRw7CUz588KxMPMAkWmDVh1D
nNeF5Av7rPmNggrzFpO+Zkbh2Q7qXOdRZE2ub4B5ltNCHijo+87u1GpDu41OF+E5
jUh/U1UvnAaGlXiqnZkYeQHO9NJy85pRTMJaE/7qI8/hNu5Zzbg7SMv8U7CdQVeM
SaJKTZhQhudoZP5JOqvnZ3sBTSip8Mpa7sf/d6Rt+si0thwhTmix7UBsZoYhzCG6
lAO9fYCsRutzN2RidgyLsdwSnpSbZ/o5v3rMgUSkBuU8BmUn+/xNkBAhWQODOsBO
Mixt9Q+nts6epp78MUbKaKvPmbTnXCvUaFuXGs1Kn7gxSPJUh3MIV9k+ogFBNYiN
iDL6hiEUX6v3A3xHHeBZ9AeGQgY9sHPJjnBqMlZvAI+Rh5ieStVwSO8saW4uqUUg
2jhmKkzV3t3ibWVAFUL6OOiFxEIG6BetG5sNVciqtV5zuQOtsPBsS/VTdrmC9Nyt
UAwdI5oE9CQkMaOPrv1frD4iloqS2F3TITc++zSKDTgxUSQaoMkDGipGDES9/ggq
PHVLMb0XzYz1B5pqyUC5cgpgHWJFgjNpRUzQB5J/UBqLPciV/QbtqWblpFtocNVn
kIvSQkvYWI04zdN2LUrRvUIz90RrrwTsVk5t2dRSgz+f1y5e/cDWsqHxeFXfi8yv
SEvVwVHx1p034JISjIF9zkVGXn6PO7ol81o36YuX21YSlfO/F93FBKR3QWpW9/6/
RpNows4nWMjqclUSetL7wAiuhA6SHgM6nWlFAyvCgdQ/cBGA5rK5eW+KR5wdjEQb
QY6QHLV2R5siYi+owq5CsE9n0yLnMXH2+rVxh+p9eYlxRK0I8plQoEYiuU7gIzMl
DdsmSLCFtmM1B9eW8j65O8bWZ4xxIk/ou9bL9FwDVMjyzAO8gUU89IOWVK4zr7eF
fnK3HNrSUnyuDoKkSvvmASKjw+/CJu7iZOOM5bLmbW1kQ0c5+Xjw/Mo1em32TBj4
5xeiLo2cO/XjJ5PEQkbskt0XtG0luPU15RrOw/BouvwsVmIUAME/XJOi+Ow1KSeR
/omhHcWB95ay1eXl4hTWktAjA/3Fmx4JmVKH68a5GtH5HpaFqcKOZYflsOugc/Mw
cckGvu0m2mqROkX2MGzDYcvD7ecMakQLH7h9Aaxhue14bnrhKLM9Ov4iW/S+uIxo
dO+mUtqkuwwTbAwNVURzV2H/M4br5G0h2lMnJlqNYWRbcVwOlIKMEiQRRCnootPB
WPYnTovkIXFyXEgq5QvG8PSNEt79ZHcySzZdCTPx9iN/3pLTO9JAfHJfjWnK2+o+
L6IehU8n1jAifcUVze07nYSNVA8FrSNOVp6BkcEqrzngmn4OC76rPCsyeBRzSqth
MIfOElef4aJUngf54Kc14kGzkesSXk83xTSmP329zkCNT4RpVxMS4GCK1S+gwfJY
5jvwQwfbJW1rlJdPteF7U2su5o+Bex2PumwcHAVKMlvRAl43wffdEkXM5vpXKuWI
LnJE8Hv5a7dop4siQLt1taYhfEY8kIaWn17KocaFQPCdVtwlpBhDK89Cleg6/5W8
3CFJ7AXr9PpVc785rZyjNlloyuYlTqmpWrpwY9/2vQthmJd+Mag6RSEhgTHyFaq9
Elkv3ONfsyGfvXPRzp9q31WDBniNzmE2AtugunDFc9RsxxHBwz4B7R1GXGYbB5ZQ
bV2dZchp3l2iJxsnozVioMeto5TuJr2yXe+nkc/840fJFfTb/nkXAqSq4eN4QuzS
KIBNEjP3f65pKUS5VrjWvZxp/zQxbCtR1boqKxRuV4Wy8zXYGr2IpkZHNrGZEiJp
XMLEY6ZiFr/ze+RJ4/dpiI9UxqY2qQmYqIIbxj/qLFUS4V+Egt0SaBVQEEqhp3Wu
OHBpPnXqsCD6cDGH5mlfi9egR1++be9O+1blq8wzMiBHJ4e15XnZQMppfORlyICx
n8vYDjuRg6vj44Q30JP+EbKRWBexuNNQB49wqDmfUzPHgtKHFUzo2fZZRtKcUgYS
DZogI9bingnr5Cm/+65Usje40L9e4UKD6niCkJS2eV1aHrdZst62cXlFBQm9Sno3
eqzoO+cPRRt3lYW187GQqgZfmukkT7HD8EutYpbtXSk1K6utPjJt9GZ0YpmsCpgj
syMR4xwfZf9gI4VIPg0ObWqtqqs79ozK8jwTFNV5dVJDSUDQFesS6mZyGDMf1ksG
Pt716lNUggrY32PqVHubQnO7XBlIPINsEC40IaAkbtVkJ8YB/XMA+J8Ee0hda4yd
sp5oj94uUZOYF6pDcfQnqbBCnPzUQGKqHXSG+zQ2W7+VDEC/qPWhfsMX/QZfMC9D
1Sn1fLP8IQvMPUX9gjAanAwja1ly/+Vdy1Cvmyh+U24ExisS9x26YcuwMDJWIe/V
AR10pzKIKnDP2c6wDnGc7HKMvY4uAkcDOiNXQUhP9z2H34tArBLSnSmCBqwNR9HX
9ZchZPbTWQ5WaY8xxvOUjz+91UaaNL8PHbl41dz7TLTsPI6qHr94tog6/Bsi2y8U
rfaZsp9tXHtLKhMBz7sgIqqX1yxrRBb3IoFj7Sw4Rp1Q445MGLRPzLbrNw0FvEgk
xjRtUypVHQw22gTU5t7w4nRnkfUXsU+zWOfxl+RkXHt8w3CjVgHsHJuqSP1ITBOf
XOIsfnxbFW/P73V7MTVJ3hMFxlLvjUBk4pRSwevtW07ApAscYEqTsl+qto+D25Yt
Prkq1qKMlF2MzrIhlTalzIr2GdhmwKHskgCEfix+CCSc5u7zMRJctmqzRPk9rNmU
UN85dJKn1SNC7vvrr+RMZrKU3YQmbOJNR/uO5f/7sahxnK+HsU6bjoWDgaVUTbcB
LnY+xHZlWjAE4ndH5CRb6X5zS8Cc8Rzz47RBbHfGzoiD+hcG/o1s+ah2TBzaQapv
xhrSRdeAnBJjFHJp7ZeVY3nORwOuXrU8PA3e7jzf0eXM7XVW7uEx6WQ658y241Od
VB2iUk3+Ka5UDh5/y8LSxDmkH114yNTYUo9t3neDNCaMJ4c+7QMVYx2fssZQMnsm
GxMY6POxBEKtEIo7/UMu7otJSFmoGDLSEIUMX7fjHxoMhNlTcPst2wagl3GpttMz
Isf4j+1q4qDhw3v7Qx/vwMtNZLByene/hgT0dhaqdFbWNhqgR18kNjzuLTNCZ7sY
A0vtvgbHlC5RtVMD53EQ6Z5SivqjKhq7NUu4cWavzcArL25iIKw5KuDFa897TjCB
zw6duHCr5R8CVvcEs7uiIBgxkyXoSk+RON4jjeC141zdU9iK2GPKbP1bg3xXGJQQ
NKcAbn3h4IlVCaP/mV3Y/9NVR0V4SBchRavoqM5auaKTGZCUUARMYagwIi0OmaHQ
A7P7U/KdVM/bKcf6kx7+veQRAlGb1yBjss4dQ5JQn9zOg0tUmtWrRanm2e7YX2OT
Dh4wht6crbEcsyppi85HxD+R6hzU58KdO4NgHS9y/qgTviJ20oZds88BKgl7Lzln
zlTP0XutI2MJhuJl0cxHDhxLilfUHgVMbz7u8BYoXvyt+tdoePUA9FYfjejIGlT4
GTiSRevXwLbfd4eIIZn/VyibaEfj7VAiNrUh4NeTviiCpX8HE75yffqRUkujWyn8
SZ8Ok/KV6WljDHiC3OPJsgzN+Y1uEj2CrqHaBhQqPBzqISoUrzPvBGKiZwnDUsCt
LyWvTfB6yvXsFDWA6RlXUEqMy8kpzz1eSzDowAXcHj4lGaDgh9HUSCwxkAd0YJ3k
`protect END_PROTECTED
