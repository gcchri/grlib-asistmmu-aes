`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IA8G9kLZpE3RlT9jJyRkMWp1hTIZgyDiz+nKrbU8pw3erpVr6KEsz383+BtFFpde
uruWG0I+yosfHGIy51w7dzZJAlnmqODiFspwSVSIbTLEpqvlwdwyO/4o38x44z28
6z5QkUeWEQHQDBUYuPGfvr+Hiv/2SRrpqwviKNFFFFwFhOhnnOQLNy25UHt42+wK
sZWYnH9QkjHzXOMgHiGi6O6LL2BSPmBJqjKjUquawSGpmsftTSFNsxZL5A/bxIQV
4BbxoF3EMIiVodlGOsRK8wqBCofFIxcdrYOAfycMUwJNely2F5K8o4nYh72+ges0
Tw2F7kJ8Mo1EnUWt0RtuwnJecq8f0y5skCv7VlZvkPiJLLZrR08fVMXaOZpwzB6y
Ske7jFSLEtf86E+yioGw/FX9y+BcRkX4QKJ4rPVv01s=
`protect END_PROTECTED
