`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a61avame9KL+0pKX4FE2t++z4DSCdvtEAazpUM5y/CJb5UZgST2eU1H93SZ3yEqo
UPQCScV6/3zupXTI42JC8eJ+h0dNbpc8fFzHR6nLSX6p0jvGBguuauef0i8A08Ti
hX1iT26wdJqZO9XfBCw1c6jJ1kcRZRLPHPVkXFnj9I+g2BC7CJWlHXSC7QkFTsBw
dbZFAkFCvDTIDCpUpggeAs9h9feOmfjOYn39oSlSv4WfsT7UX85WaShPrGEZrCX3
wIb6LvQkrLjyWHrLxmDbN347IbTa3r0+bPoiqEDZ3LDOSUWJsc2l3bew4IuuIJck
/LKn2pNcn/5F6W4E+euIo3dJMdv3HBowQzDVTK47C8xKhdjvwhl+irl5zJy8rQaY
YFpCFlPUEHpdbrD3zy9z5Gle38hKJ5zYN4M7l81z+YRyj8g6hVpyd11WjkFvlE1G
gPhWzyuGbQ2ay9ZQrIdLTbv9ljcrzlGJB7egK7MtsmgLKHw4OT1OjzZpeeeBMrc9
`protect END_PROTECTED
