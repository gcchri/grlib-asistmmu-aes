`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URVMlma2UQdNUcKC3BfhoiTxOetftSWN5osXsOJT263GH2oDFRfDffVjpDWEQd34
egfBA5smwX9d5aQpC39Fr0liivbP7j1A0ekuR8f8BSQgEgkjhiu1p3zm/yY5TS7x
iIzqeqqLErMAyV4qwo+I12U8q/Iagkz1GgCG5vC9Z/cxJ8QBMR7eNWI7iWiXsJxp
2U9C6wKftks/gHVqc6U2zdv3FvTSxKmL3eheW4FqZtHG4wxMFuOYCHctjTRKIfYu
r2NCwnZToWsvyJQbXX4FkR2HD6xvbCUWGqLSCjqgb79Y5iRVHEUNK/lnAyVRPSBr
NSqByXD3hRcgvdqRinmp3UBm5W0Dd3qD4YdvM5a8MTrU54NCzgsC+YgzvuVi611I
AQ4TDtaYIJkaKeRA5/1hsWkjLTMvUgX1ogABUEimlBJ25nmihEDHP+qwIyIuEF6b
+Wlhe9rTgsUBz36LCcDjAo1pyhlwLXoB83ljxo5DTFKVSN5CF0mqYxjzPicn2s44
rzvkwlbiEZMlilP5+mke4N1ywhg9xGu5vioUKundmgY/YEF9pKv1Gt19P45tDIHK
iniLcBmQPS4TJWLozSXVvc+MiEdB+oVv4J9I2GCiFJmfQROPzgfnfq3ek5/cYgjq
/zxY8BPQDlomIlVE3DQ8Ra4sDo20LbIAb1nNZyMozDn3m/dxbtMZZrV2bIBZ1vSb
9cQ7XkWMCbaTRMEBGNsD4JFrsRAIdyo1ZsCrCQh+FPIjgOkX5oR1219OMi+YsQyS
72HvCRbZTCqYeUIlaS3DzjldqNmTa/+U8Ln4waPgGJSbz4wP9H0pQaj0n+ywyd3F
fq8nOaqtnia0k6VJ6fBQ+eZftCKFkSHBtLW5e9kJkgEXBw9DFl7PQYh8tEo6h9iZ
z0IOU/ayqlVDcww1iVw5t71gKjEyyiCed9X6ToXXH498J0KwLrezXedZWNDnAcpJ
K9xw3LTjAxQ+aeTBZTl8OnwneJ9/3tAIAagt+k7cNGQa4GAkJmaQbrJpkhxywnAV
klFvzL3OXixB/Z43jtolTAZcLRfWMtgvf8sMFJLwE1c2j/FEOOecLy60yqXaQWdW
TN9rpvBxtsIqWTkxbVy0cV9LUvqHr937Smy+meuW8gSK8uplI2xqpMtq7zpTZkSn
vlMDGAuzoS1FsZWNIl1KWzQ7wk2nR6TWYB0lLakcEQxyqIKY+yuXnj6xDLHa4vAT
rCbnI7nGUlt2vsuWOdyNHaJutjRivy/m5cOiOsxZqEN1iqP90ryyrMFdGwU/EDY0
G+daWU1EqlCtH0/kNLe3310Ki0KtbPHGxvnHS0zvxSo=
`protect END_PROTECTED
