`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFC+LYb7kfFUnldv63aSA6rgXLUOUQ413RWEXSYXiZspVehqvYN7tFKh4GspKODU
OWqj1rWhQid6N9Vo8eDbPnIDBp0Ghcr3+MATn/uGFv78IgiXmUwoynnSMezgkS9M
pVHvvuZKPWPzpTKVnKXUfqC9atxOYPsPdCyI+r7YyVChUn77l1RTf/YeKcpJCYAC
oSsGNmtzEHNOkPO98TN81psU0H2c8UK4Gz6l+R3b+sZKEAFyKs5zGBC+htsIlV/y
MthLlZUh5TD+TV3HZKDF38Cb8OI3DCyZ4sg/dALIJAuIjJc/S8pZ41NLSkf68BQm
+kV7raUXBbLqyl4narwHOdmVNJujucjNh/JEIVeJ9UosRPlwhnAL+HjNB8JErzWW
yGLVo1k1F/9p+ULxWXfwA7pVuSQ4d0SKIPszoQxq+TCUwMzUAUr2Uc0o69a8+xGz
7gWP3VyBqvO9lDOq8ZshsAfFgy0qzj+EL5KwPTwmZqTMVezslNg0i+jfAs4CEeYY
5NQlzAF4zhnVSp6ToaysoPBzqE/rJ2uTCc9B2OlQsoxgF0/02Qn5fgI3vFLgC31M
WWpiQyfKw96uG7urCVsVIVxCLbDRwG5K36zY2EV7uUJtbTJkeSQouuY7MbdYSlZC
tLB0KXgI+OHfRAtw1LV7L6VVGY0cuNkO+czteQwh8HkEAaebc187jbFrPFnqKuTv
wXzxZC++EMnQXgcGVshMjVVpsNuyIwIwuRLr6y1vjDnMroOUVW3vQwy9fXOX1kPe
L5cwpjmZBAS/h9EblI+rcSpU1wTfEp4yadrD8luI5f6hJkZkwYtLutPJSrwODi2d
UIb1ew53lgX2VUc0VUQ8NIF0nEaIF9fll00qV1TC0BwnPMfPf2ugM6RN4uvte+8A
PAm3Ak2T82mu3iKUa0gBuQN1+N7QHtcgj5XLasdPTK40BndIi+px3RVywVA96IdW
0AqyEgjaWhbYoUVa+LBmTheR0YSohgrwFJ19Vxuy1Elv9A9aXVNdFYzfisnUxc9k
WyiL7TGnYqSxRvMSVezJmMirsd4mDBUovFhJKuLUYWjxLlTM2Ch+utZl89qanqQx
XQABC6JCPDA1GtUo5q4mtz5B4gbkKrceDixJ9fevcEwDpq8l/TdB2pp7pSeHQ1hI
aJZzoZkeY+jjxx5MLhLwhAYMgqgTgrDBOM40IXPkAdTNV0CFJrVHiLvTqs9pIMCm
HgSF4kBLhBV2K9GotHYdEFwYG3CtnSmIWd/nbU/qO/HsofRds+QwuIKJvoVQwiwL
I2FOR5wZR8sj9/HPo+AqNqLI2gLCIWbO9ycfzIkWWvmgEdJWwFb3lfKpaUgIV6Fq
3GcvhJEH3MMpM//6bz08KHVYfTFstRCJQvoRcuq04dfiOkvKSFv6+XwMzMbFSolC
65w6dRbWDl4uX+soH2QP6F9D1oH/qdUcmL2MPeX76AkxBEj9SvFVaKIVTrhWbdWN
ginbuuumQ3+YkdQknrfNCTKqIo8qSruLgU4QQJ5XAt/SLzMouTzxP5CY3uB0iYvD
FnntlG/j8GQty5cX7GdDZQL3FxcThRzyT+52JTu/45h8h+GgkqCi16SW5ixljRPC
jMgjLyOIWtRyufU2MChRE8y/PuWejhNxds82ceamLxkkDYRiFRCmoNrqxjI1sV4F
BkSFweru+xikvGGklDGSt4zVRstWVFP1/f0wiBcWHCw3Hnf2rXKkpu/YQ23w+h2Y
m64VY05FDPFHv511f7d7zHxgzzeVbxbu8ZQA8PJ8D2FPHKpRP3WC91AOLvdbs+fq
2s5OAoOcHY7gYo7gFCmGUB0paggqkh7Ozm+fjdAbN9xVGeN2xNzQ0/VM81QVfm1F
wAVS/yUqmIFc96AE+HGm/7x38Z9YqC39RRv3E5ewuXxtjEncQDnoCY8GRkficg/Z
Rm18imFECKsF0kJmGubKXE9O083xfrSV9GDuTZsa87IPfzUf7EEFmG0UU2lQTled
3oMtMtCdiljysw8ANUtvWfRoO+NeirpFtCJ2A2N6mjZlXbLdOYZzb92VgORk+tuC
cxrmU173npdU5ws9B5cafUdnx05lC0kTkU75+j2MeUIjLGOxtBKbKwg7C4d8eq6A
mySk7wVMxhbfQKceQSn5EPyMKDu2ILp8+W5zyvwqQ1y1mYKzNq2PI958/lHhfovz
5REy+nMQiUGavDtqOah4miOaa8zfVWyqXIdHLul7YhAVN60i609/s0I+LLK/rnjd
8HCW/9OW2yoa5PiEhRaCvW0UQCWbzfXQX4dhrGqSWksbZl8I/wb5QPLRw5iV4FSE
TiZr/FUkAcxRnf2n58M+bQEC1qF1StHmKDaInsCwOGnHVMIR9J2celIRFj9Q0Zhz
Iw0GV1UXMME4YyaM4bXyYaLiwD0eIr54lvxbr1tuWK0cDmvXn1o5VJDX2TQvXBug
FlyyRPl0xBQTykM8PVt1LjzxNDhfSsU4RcZeXBhijY20Gbw3LOAFUWcozIodj7Bn
+3r4U0GPBEWaSW8eMgbQ5Lc2D6jCkdb0o8IbUzNJRDwKY17E/vk7/kFVujkDPBYQ
QtITnzwipf/d9lbozc9bkHRL/iJ4lcD9s2FUhsycM5ffhJYH7VIbzo2LZYRxMotp
+OgGrqYh/QIgbhdhCvKHOYIRKrzd/LTv2VICK0upnWUDkoeyYCU1foNTLBj1P+ZO
O7TjqLHVJbsFShqa8q7T6up5sR8ma5SkaAVg7LSofs73m145ySU7kO4A3rGQQrwc
pYAE00jEMampE2ckte2ZpDQJ0BI2KyAnyjS+obLWcmVBGqCxyyKgylQNsSkpOwgn
9+vQYAVbg33oosAdUNIsgq8SmpIDLt/SfrlRRbVQTOXnsPldckfjasybuNnQdI47
F5jOFuqS1Qnhrz34KQr9ZNooopt9QY6U4KpNUsfTea4uXbOeKck0TEpUWXDGgSri
QZmQPmfyEScQZkOOoMGnjMq5KJNTye5OeIJbdMzg2gosZv0sRVyJuBxYf1qOCGwK
+2YTUNVlF6CajfqCfouBnbDS9chgPcAIdmMg3yxfOeku0F5/atOTiRVHdOJ4k6NG
WA2B8Ue6RYx8cxufh47sjQu2zqfQ176uIwNM7idokPzRFYep0U4kipdEVaH7cT1K
V9/y+QZ5AKCuPJ0UI5ydg3dXFAeYxr9ZQKHcyrbCjbMq66gYsXPXMES87qC+TQC0
K3OisCZPD2ws6J4C1esqQSOSqDDLcEyv9rVg9gxq5Xjf7TTTPkgp/4zs97FAzVex
kien6d0iMorws2WntipG+EeGozErFkiuuzbKLotrfFgg4dCpsX+i0ZeHDPMnPi7l
fyBhMPtglrH6yNCiJTD1wBApSOE+ZkQrfShyXQt05N8Y1hvc0b1ctp6UEpCsmfdT
Rc/bM419bucghTNOJt5YDtYlV4XlJPgyWWnqpS0tdakilnveEyH7RMlqaxXc+Icf
z/9Y4LpP2Fb6gJHnVRcvRjvtzJJtty4ycUz1YeBgPcU/ukovp5HPVuid0h+/dvzl
o4RX5FOtQ4KXeL8x7UMkgzDOJrHftnzo1Rdj0r83H+d2a9emTiR2tm9trrLH0KLd
sGHGvm4jWTqvaMlqR47q0EHW+tfxmGru9xTjAWOrw18OBApA1LUEl4H5geG9ETqk
szCz44MjxC4/wnL3TrdBeMU7A2e7p0OXRxM6MA6Lx25dengoNFcYxCbnv/CSdwdm
9Hl/8ke5ojGElBjbhkMrmi6bemTw/0BUermyskIK5fyBcsH+lzSviibH9BfUf1Ev
NZmvw8ZTv/3mjjB0FopA8zv4Zl/ZLFCe0xms7J1hpOSDuWruj7AckgY0KTmkedzt
QeGuRx+NIm5skSSBsX5U18PqjHuMKji5fjX25KVuNvbNwEz9LI79uo0vkzsufLAN
XeeHH6mnm2lhyt0RcpQzggwKOJC6iqEdJHu8IQbezpUUOCDMjMzS1sgP2d6Y1zXF
+Fr56NT7oa8HLgobskoztJ2J2s+YVBqdz0MV6TTOFLjhXcoH2xxk+aQOpErChMug
KYzC4kF+WJ9LtnVR791RfVQNwtVbtZuTfAWYMZPiVBe4ZfYNLJ5pdPiINl5RGYNq
ZyT4VwYe1FFZdR1hRhE0hQmGcxPMQIb74EFA+eAVGrzAQnFEMvHfXTH48Qo+xQhz
V3LFvb2o13CzAcNoLI6EEcUCKMUwiYCkERq92UPIQ8Pi9xIOw8o++2Icnld9a+Om
HHdeYpsbgLeG5Civ+Jlu7XWfWfqUf2vXyZtBHGd/n7pALBLlCZny+NCtBwOt/HM1
F+AzeftbWjUri3bLkAIEW8uNluqmqxuJ72jh7bbxyeI76tywmzXTjU2iMyp/JCpv
kxTrG32DCNYt1OIu1BGYy9EaIhxxm5NAQyLvUd5drCc9nzoJUq0GdZeapN9yxKgA
vjl6v4GSDxAv1wM7GSJmffoeHhXeNptcotKOlMIpH6ryTn7774PwxRIleNLz2W15
St0NTf44wh9mHfBxSYSAuobXZ7Jr1oc4nn19NGYMJPInuBp9ODn3Rj325Vbo0DDC
h06owtnWTc1OUfDwlLZXPKy6jU8TQsqmMP+CM85/7RFpoTzDueQW3AmQSWpxGkTB
LkW6UrY3bhUWiXgX0wJf+BM1c5n0Wx5baVY1aS0rtXjMXuKYq5nVjq9l4i4Y1BhI
yy/nobqq2jL26ZWOz6RPedE4WPA5QsH3s/hU3EiswY3xE+8Dqjnwcekhb/uekVlc
g5XKSpdzHqimiAHhD2F2nqEjBhpXB4KOHNCWV6j90ugysmyXtyyuvVS9/uZNbnm4
fl6q1hpHPlJ1SZ4OyRCvfhQyJIzzVnfoR5G+9tRTQunzpdCYJk1kO92v236OlDQK
5Ql6EhV5fwUvdGmckaNjpFOlwBYj47Au5oDJT/ccuIJuQy6h2z+5wKgzfBqNAylK
vFwgt29zmOmoUuKEPf/EsE7fkz5TqB5Gd48tnNjLyXJbDt0epPeNAB96Ww7TSoi4
BVasodv5ICCG33FdcyQifmBKQDBd89JBZ2Ko3BQ6bFnWwpa1MAKueKYVpDRQbrXB
EawQ7PRQynlXzEWeBYNM4pHWVD7wtVV+gCx8N6DhtsQmw2uwyid6Nt6yWsAa1JAA
jeGdKnM4CLQ/QWaZ4Uqrc2w65BVHlvYfBBjH+X3beGARvfrJxbmFjHdtqWu6OapK
zc5AUV1lypSFBIaUE3hR6DbFTOeg9b+8zhQEpodzxZs2b82ka40KjIKPjw+1sIac
kMC9HUlCZ2aAaND2h3cl8QASj1+zyuviN7nyPG6D2DHX/E9cQfyMSHvEtihLZPvy
qqeh/87kbjhct9lMrY6m7W8u+JoCB2oA0/FPwre892kWmjvFRTbfdPwL9xeTjKUT
N475hcMCFBCIL5fMnslk3BLwgYwPiRa7yV4uQ6E8QqaQNo0Y6ns0ZMvIARaZnEwM
US6Wru1wCcvkgDDHG7mc1NQbGeSAt+vntV62asKi3V2qZsoDCckSUQ/QCaioYXpG
jy0yaFdzj8z0RI97hPrYAs0N8TZ6ZjxP19QIGS2oz4uC4zdKpuRm+ecqL6m4qUFl
Lnw45n3ZEQBsEAHp/oDLNZ1hdgrb+/wpy/Wsp/L+EhPhWFPyL13Pxts7wZq3sEmw
uKOvbYB50KORQX/crW4yki4mU5/iMUTDBlcJVcqVimjzIRstZnuZNx1Iin6IGTs2
r/OCP854CQYT6YeOfywAgckPwUWOe+KBj22K3RuoOFhif68lBnHiNW8IVgyxouPm
UcazHHty0npHAAx6FIrMpIUtzfTmuh9bDkRLaVV+kNyE2q6LDcX3hzUvWVVn1hWe
u/sh+WLUmkQeuhqqZ2ZbcSW++pjrJx76RNTjPeZsJkJBFPd8Z0qS/uzcb4Y0ebD1
iJlzMyW5mfPDUvw0WFLeE1vCKua1qtTbEEbMXROqd+JDp0u8olLC8DjFkCWZjYTJ
oyNxsLMoOyuB7CIz/TClKOakht6i+YS7BJiyBcf/HDe2pjL/UYs/3naCyJuf319q
KhyzSANNjpwYm5129+t9xrBre02/yhcT5flsRnCruaWnz8BuzXK+rQct5FcbM3Gs
zuol/ReAdGa4mLW6/3zID/DnlALdsVoCFRuURpeEXUkNVnyMl4y/oWhQCq+Z11Cq
wwpiPuJesd4Lhea1cu2GiBKJpsBmbYtnJXLAeNEf3fEQQRbTtWd/fQXiBmKuZR9u
iGF2Hmg213cCm3sVXXiAopUjp+GfK9XSL07ynituSpqKCyrUfSw9O1r0ULqOxD5J
xF8VLtbRv7kuQ33qC/S+DcjF472rbYLM2nz6Y77P+5m6DoZH2bUhjEgbrZcva3iZ
2/R1RPctrEXtHcNJcT7RYS9xwUy1mnDTr2LF3qmTWER49nqlC9/e2BGLi6iN0Ijf
FdAOC90OexfLjyqT1rw7DqqDjXRR60fCvUcmURwWjKuZ9eMLJilpdjICyguiP8jS
rcNcZ0w3I3gPoZDeAAPsW0So7i1bT8c/C0Qwh18eY/q9Kqm2wy8llTgL6RXwWmN1
CjUrYEMaFVx6tb7DfEotGnT6XvNdQktB8iIjxHbr1ElrV53FThTX9cAORz5YxyZm
rW1uLXrr6VByqTU0vA4kf6T99aueGW46AwWo8uhuqPjuY4LAO1+8gV2oHN/zHnnc
rsBoCuqqYWR0dRlmtBmxhOBkHqIaiMMZcCIgG2XCOGQ3yDsZGnm32AMawmY2gBay
hI/swUFu8lvcdE1D/xvKL+bQESXLlKURwF7USkQpJh3NziiE36fMu9h+U4MTa7w0
D6UTEWcEKVU4VVKVwTQiO0+JBZiPOnoKgWy6h662tP0I6FeG6HibJAprSbzuYKJr
2fNyfNSpniizo4UyHIrIUquv794UM1ERKA4JDuB6YsTDEVJ65VTSK5Y2gGSYzMdb
u7WwPtxBcNvjyrg1qfhFCpHilWTv9POLecBju2+eyg/oR0RToMFCYHcm9cI8es2k
k2SPvdOHyFrcHJ9fZJp6+yelH0k6puRwvqVFzNhsiZfhNdvaX671H7FEDzBrSU2t
3yj2+MiWOtlLkJSRrQV8tOKlLS4nfArHVZl4gZs/OdTnqCRXKWLf713GhbdDxvr+
Esrn6mIf1lOQV9d3cDL3meJk3R9AQu2tV4ABBjdwJEXdIpKms+OAI9/vnGRwiE4J
Q8Un0iVeTy69azJ+wi/dSc4akFuFLa8y88IU+XbexQgq7/LkS0mNulpidrdV+wiU
kCBgzEnEBgWap650Ac+WQloepoqHMkXuKYwP3Zx7QyIfXYhNUB7+Mjh/iUqtWkI2
OOEJsuZrx1Usu0r6KzXbpehnNvOtqUjSiKEM5ArCXP1hh+bY6pgwd1tk3frPEcdq
g+3cwzHVPM22VyQble14uEpjox151ShuaHBehtAGfYafht3wHv60W9lj20Tv2IAw
Gyn/Shr3IsvkQvmSQsqSmMOdipgl0N2ivRTgeXoUPyUuv74mStNLVzwx9ebUaNFv
4Ie3khz/aIpPrLPSu/W8z1SnXAK7MAQXBBaB6dAZ2EQlGaDXoj2wdKAONJspv7xj
B9AvXqsaRVGBqdg//crMH0FMqSKDw3nToT0aY/OFDyt61UIzBvG5gpRfQgtCD/fr
IXt/r9uQB6lfiAe9vBe+lvgvujYamcTk4oDwWumreOBuWlYZzilJxyn66VQ0ayz9
JFrZ0NHFMB9db2ufccei0L4H1Cu2sJqCGqRHN78kkTz6F0HQ57KCmieAsvbZ6PJW
LY4n2beVRyRdzgs5h997i/ZWY/rVwxSv3Bku2XVI6WXSXfajZeNLAl78+pmxicve
oQR5Ue6W/j/iXqzavrcj0I8e98C5kAAeFPHefickJADUlvZoCc7aoP8pk80xTJkE
MqMYLmRLuOwoTtz2vAo2AIG1rlxAcdbBkh9XNaXyvw2MKlSN85mAXPtBrJBZyslF
nDIWDOFijMHuKPmpk3suULFm9sTnKdyfXBeOM49w7mrSJE1bbq0rnHmnKxTXw9Hd
3nDzeLrUtwkBEBvhyWXo1svro2vVRkWkqhu6EMzHovH/ozgNvzT7uICEai18ivQE
ShpwJPvLJW/Uiod08f3qYMMS81Ng4cJeROp/N7WKJ08ZiEh+Ip7LNcGMBtjdiW0T
x9K9VWzAJsdr0PHAYZwQFGjipavf8spp0B97rkQK+AC5AEDlsHuNXeYLBxCbdKRf
pAE7uydguaUxm5KkE2MVk8pcBmUR58//+a1dfR//3xAXJkKrFSkRBVjFFA45QfYl
0yzAqMkEadg3XQGwhp2OazMQWvaNkjegHCjM9i3fHwdpjKG92RggljDFZyuZc1nc
0KqGX1sSlNQIn4/r/DD5QTPUOSqRmedVRLWJ68zgHR7PZDwyxoG6qyYR3pt74bEt
4q54p2W1/NSNcG9r+TV0zofaQiVO9D+uV6Ah1aRlGHIpGQNKeKS2eMZ1UGyk6zZc
53owLHP/gVDNtbPMfgvdcy9qMdUzBUom+NxrWCqcpE7C4ZMegMnJ90SYnNG9mDGE
LUgcKNWG/b85ObgelPHNBnbL9wcQPi8vxR7Sr4TLLIqYQrchNKnXdazDxmHVRPsu
iDb3Elz9R1aKsBYnEo9Tdi8NSxeDcch7dvQ4SG52UhYcBDQvFEIR2XbZXqSxzyRS
1fjG0Wok1K24VnLwEcucFYLkdikTJxWKsYvYL+Amlgu+yfRPAofiL0MXZvSEAzPR
0UB8HuZ0VxB9aAB/iS9I/lUV/OoKR/Z3nWkPSPaGWZaIXg6vVS1XpIKsB4yERY9Y
hiP5xdn1qd/M0yvJjPKOBSPMU0rJoLXuSEXd9GOvYcir6iKQ6cQ/DpAb+pZRGGIZ
6PdXxkx3OzOGQHNCcOLrkwrb/Hnx/RltZ39QHfz/uWY79570T0F9YCxE0r/r6rZu
ehXd+sL4jVcRXyqESWAj8Z+dS4/LAKMp/AFOalecBAp1UdCR2TlHsHVNdQoayxZW
fLOC/tv+2raT9x0YPzwE3Z6Rdbe7qMNQUXyVD7R/1CAGa7F4hpGEZkUlpsL5978q
7oozyOdrr67q6+iVLqs44sMRBxzNhc6hJMu4E0owaONq54Y9RDM30rDupltrtBx0
Qe3HJpdhazbyy6ncQe7gdUEUhJXgA0nODfliW44pdS3E+MW3/xaje8tvaWK3D4VW
tkgiYFqm0BQrm1ogHQUUf1X+zLn33YY9e3GnOCCdQjcgzfUKLb6PpFs1AAVSLVdS
hYhldxYY7hEnoTqD+pr1WSeZ2kQLSI2sO8xkH5SykNykkETENi3B2s7cnpIJ6uUI
6dFxVubajjZK5fOSwQJtiQXKtRUX/jl+3H90OiDXZT/4vYb8y96Z8MFcEoOTPAcN
4PjOwAN946/zp32dS0YVKKxbuvJVzEtM1RuiyQT8sKScc/7Ws7V8zWV63XFTUzpJ
g2z8sNBmr18uGAsE6nKvGC3sT3aMgxsuWo3jBAXNu3DbOGR/eSApIJ+kZrv1RKZq
d3aovKsONGttviBC9ILwgVcKjA0srRNFbhv2L/IFy6o8RgrmOwz1f5CLbCuokqpP
GlrUWjeXW6XVs1qVmHHqN++h5AMjfvP9kEy8WMlpnDyJCPvMhquN6IHxhc9RqFNW
aA+cBzjyDmzWXh/wGXURWVtkbkimGdqZjr1UB0HjoECtdZQuRhR+Gejyth6cuDQ8
TW6A3YjjylDGpc6N1ZbYZI7hI4DwuRTKyv/prXzK+iemimLyQGHy911gXH8F7gk+
m7U9J3CtLGlqT10VUZWcLxQzgiY6BwDbHlDyvG9XKBVMjutcng01OXHXzgk6Xck/
WTYffkMvFK05nK8yrnq8foML9quhpY7OMYizxkl47A7nFkeeTrMX4Xvc4DNucO84
WsBLiH1JMzVripXru6jZMprJkg4giYCHQUgW39ZnpPV5M5/HmDpgQrJZyLVjW8Nm
2nOUken+qQdixIVuYimYJT6EaAo58E1U4tkxO2b4sGyUhMZACz6oLKe9/I1sLfcj
F5T31w1ONRRgBCQVYqIiiu/2+7+rEmqJmX8w3iatCCyYGpUzOpcOaqltp1l8PrFI
4QV0fmPdK3C0sJjXq3NVAOx6OMySDnxF1lRGQj6rGMHP7z7ZzdSjCnnm4na/wu4D
3jX/a44JB9Z5BTwpOAP9m1TIcvtuKY3p8vv+GIfqQxBJKZ7gu+SzuOGRKdDNHTX2
FseAfQTO+dCrDsDdD13oEiFJUFsq5EiCV+/4mVBeQ31TmYxDV4voKEBMDn/Ug+6t
AurlmnKIurUm48YnwN/xF5bhsGHCcIhdtTfm3vYkzA31FXc4PI2D3QK6malLPckf
rjYHBFybQrV0shgt6Yb0RcCzM4JbSboSCKcVVE2aodRwrZN5xV2teR/f33t4Dbyj
gpbTJmg4v8By2OyHS3z/yFVvy0x4heFSGuTkCB4vrCXFA/hO6BpPI1villt9yt1D
g/wFquZnWUT32aAOKdAWgoX7yQods5KqAEmeKhU2cZ+ROPwmP9QnKtXElHyhLQuS
oWWIlwV4mpyPvZQjStFqM+CqurSWLqKu2E0Rqbv2TdwFdvbg9t46iuWieb7D3Emx
1QUMhQGQIH+ywQVZTMFkBM6zPeAARtVbFETvvqhX0Xsh5/1PhZM4xdieZCP0l37v
Xz+QvSoodN4qlBC8C6kN6axwBn9vr8UWozfflMCwnJmCwv9tmCEzRJLjFq+X6Lx9
8WrrnldKRMrbR+CbGr1n8Pp2jdZkYj0upq4SnY09d9yVpwGlhyjEtNXzhAzjQ/ne
k/F8GL5TFQTxyonT6GDyb7G0zkaKh7jCKm/vIQXBbvwF+nTzEbGPUy7hE06SKs7j
GXtCn/kLENs1puCHkn4TS8CWGMdP2wVFNAR4MwCew37X5/QL74h9ygTmThc6NLKn
54v6KsBS2QgLNTVR0fVbmx3hv7bRsUZCsxoVYPz57RBceELfVoHC0IQYbxiNFol5
A4h+5fQrgR+X4fPWZiiKQi1RdUk+DZu55FkAweNcmldK3LepAFg3+5Mk1uJ/x8ia
2QVeg6UkMc7fU+/gO/9qSxQvsBit1ewV+ty95+6ttjORF3AR4rNcXrbYWubvtcb8
ldeCcxAJ9Y0Pt5Q+T8nl6Ks0c92dlPlWOkGfit39xOFsVhCyoC1Orn9c0ZNjN4Db
BT63P7uRoP/Amk+tJ4w0aJSKgv2mw8GFDVqeKB/V2RFEz9UWw6Kl4ojZ6Yd65cZs
982cEp/MitHgSBmvESEGWlPuFIBXZG65cgxlrsX5EoiGRWw3JHYtMr2RTR6f06xe
OjxRzGlRhxF523YpEvtKr793IGZRnImcq0t6tI4yVxecxm7mg/vXsbSlrZ6gkVLs
lemxcNa/Wrt8NbLbwgMeodcHpoaGGLeSLDJFMtF1kv6xICa9PmBhVB0KOIOB5cDA
Dlh2opj6O53AiCotQ/nROmeoWU1JuJTZs6ucOzxv+T/mtBHYvr8umng1BR71tpke
DIVpgBgKVeXaa+wUugFC3P/6gz3xOegIwvlSjshcj/8kVlmN2BEmcXld13F+NaxO
BZvnjg90cQH21/6yv/vydNZHAxB81ourD01FyTjwubtarLjKN2T2sMCcKPqTBUa4
OtUSw+jrOlf7DU8RU4xzl8bQQtrS8O9MQgqljx0W9gfb1c7Pk3AVRXve9tigHP//
AUAbGJcazkHhi6eAvrscJ29ATijz2rtj0dUEKIJapkNE+K4b/PwqTK+IwA49NNrN
Vc6kvNV+43iz4Cf9PA3CP648uE3jUNT5mJKHIJnKzSstPPhEXsdNOo1q98OQl33w
BWT+rr9ZnepMLV+Ea5FP3dcIFnANI2NgByPMQj6fiS/xFqvka+qFA8PVtu10Ik1y
ATCRsYQfoEAs9LqQgfFmb5OLig2kVfKIfh2xoRVlqJFpUveWa6xnAa2sqWOtwlZJ
oYGgjS26C7PkUSUvCxj5WCJUI3i/4dsgEQWwqEkHpiEdF2SVaRtEhkX9ed3OEunC
9SqyHmTlvpnhWCbDod4r1UxGljC6kKrDlEKW/CNQ7fKi0YO/7CtUUbbM59cO8mzZ
PkKPD4IrCqr5Ct+2NCX/NGhlLllpUQvQ/BRt9jqBQ/RavFnCUdQ5RptDCveDUm6F
L8/U4QwZnan589Qy7ubk8II0A7PB1Bx4kARAyZnQl+of0RYkjoXO2Fqd6yQSMxNa
sH795NHDSF++B1pNFQPtVy45JH9GkoFUWQlVJoXEV+UT/zkJgZpB/0QTbatNA2wD
5uvHF/VvG/quUDK0Q/aMutA+/iQGcmmV63eP+PCgVy3Pg+gZiy7lPiNsmp6dYkRu
pTntpD23vOd6UogFFGPeQo8jp3vL4izV2ZRnZoYdRi2KHFEMo4jdpOfXk2MKq26D
eBe3oA6NZGdHvYd73KphAurOmb/C+SS9gtVOG4tQ73XiA9rO8hGEl5b3d8MKeIPm
3rLs8wkY6qJXugMfHdgRye5vPZUKMkSSEc6OGn8GydRee8Z+wZvioCGABIxOvssL
2whXgCa/8aGnTQTrdCTnYPnuX0K95HsWHoawPTSkpnF4S+StMReEPCDGNjLWSzTi
cyzjdd53iQHpDh5qUDjhx1Fi2EraXc7DX0j56BDyaGXdR8BN82LWlj/BoNFdbk7M
hVaB9V34oftvgS28IleBZW0pKqPwItZv9bfkKa8lfCu62uFcb+Z0/wDkejJDn4uP
EpgfbldW3q4a7pJWvUGelpFpLov0i3qG7yL8QA+zqvj0j75F5n4Vbt0BrNlX2A2E
P8jVlS6cxz8bcNxbNehT0PYoKyWPPi4PHwiyPB+tB+ZXPKGoeHXehFb8t/Z/l6Z0
NTYKm6S0OkhhYV5QX85Rm3e30tOGEyqrRfSHcEe+sJcEvlb6523Tw6YiXLCsHs+E
3sTrnbE1JV0UnZ+6918SMIEhPgc5H7ZUkb92PkrROu4h+02xdGI1afM2wbuYDXSt
qqEGJ6FrRC6dTbzar+VuDdAuLiBcOD0aUst1DmEcm6IfVxrCKIuqjJv18NoW9D2w
RG8F34uifoKa1tZvGzXNkPT6d4JpW8FrTolnzSUT4E1TBFjZkaTTgWMzlPaQRFCR
KAAksXxNU4MEs/H7X8AQQxpjVBkb92IlvMBrFpdrl2c1lxGzMCBOuePkehF2jbYy
/SEIXw6Kg8jobBY7mD66kdg6rjVE26G3jTsyXo+2Y+WWorzLBOgvuEioRq42DPBk
lzf0H/NosbxmbG5CvTJKXGmmnTq/RGUK7PqGX7zNtpaMPimtLYhq1fo2O3NZ/apA
W/oKaWF9jhXXh6IpUtKR3jkmzTJd+g/vF/dxNKKfICyGXSgbbOcDe8RqlM4AaVYk
LRiYMYduuCNBHbZRN9T1U2WfuWScctY9Isa+iuRb+W0wF+j0+lTnslLLc8D1Vqld
8moVeYf4h38vSdkITgs4AG9C/33A7qY45LGGp+j85OWjp6iM6k983vLCP2X3FXw4
+qESNm1HbZJoc0OAiDhO2GszqVdYDuffcZ1xgcN1SXyoFk6aFyC3LtFVkQEQ43/e
LnbkTfDr6ZBL40DZdpMFWD4NuYw+BsiP8kmnwk9EEMQym3BPSrFaDMrv3n6VZWjy
RcPIW3MN4uIZlrZIE1JOF18Y+A3r0EW2d46FZHP57PfN8g3pH0YwntbYsp8Z1tWQ
217P0DXNWCpN5zqc/rmttj4cjrDwqVK/f3r6mbjv36trhC7z6MFMgcjFDreKnyX9
XSU+Vshk5b/vy4QmYUOCgJc4gTOy2fcC+knFxLPmSL31aUXToTNBrJz3Wt4JfgaK
pcqzskPgod2lzPJ1BsmYGiGfSESxClXmdaw1okIS36vV8DQzJcqE5Q8v/S5XUaj6
ZQEAWBPX1xMTFyd7wtfcH0CUy0ZIxkj6XiA7SjCW6jGjYGIFraLWRGGtNECWG/Mp
jZhx9kGQrVM9DXzWEkqjAS1Q+M3AbZ7ZNs2WuyZ3DVK5OMRF9FcCk9wsyf4xjlUz
KWFnSfQyV7ryfreS0yF1A0q7GRtBKf2IW/ToDa/xfPAZSL2KtI3pnmh3TNb2Hdv3
qPUA8iUkIS7lw9M5h3tuVWNynl6+jkniJ1fDKRj2WYj/cFqFL3EWELOlUcaTn9uj
KqfuoOdn2tk7irkCcvsz3QBgilwkx6csHNmE3S86KpsYbiOcS6EySzmnH7pbJeWH
BtbvEPuMq/vcoyehKMcpRv4toqbvCYMct6h+4eH56BzVVRhbXCAYbmXIHHzm14wL
LfnuUB8pk3oV0A5bnguoWh9FbJiF4m5tUNLB8XcY/pu45PTc2cGDREVXJg5phXq1
6joTCip/INSVxL3C6XdFRdMVRiDIx1iMUA8AveK7K0pb9MVFYnFWmNodfBLTSLNZ
e0MRyE9feyqNAYFziyvSNE7HIletDsldvmQ1XUxk7czCKFUhToDBc+VkommXg3y5
1uADUTTxbOHo8As8+H5s1ztXD2GucVYj3+gN8ZKxthbBFvHayTgsqSckeMekYaFN
VsTkC/HfoS1EU5STBE5VskU94BNX83h4gss4+llPlJrvwn+IwFXPz2lTRz3yOIlf
PG+k1Y1P8siwva4GohOqDwtcrtl0ecntfZ+6R/zCqZIbaQo4WFqVVYyoTUAzzvhB
D5Gk4BYK4WKnSDqyqGJCAwPzIxCsl7UXjOD9kVLPE88dRWRLnfcONsDNBiu1JuVP
OLZQ14D0CbygutUaenRKk5ujipn6cJmpKo9A2ErzyoS3P7y052KgCVDtk6knZiPY
4ua8PvYap3qIr48UvgcAyT/x2Rq6g6gbWr/7F585gNe2sp0P4MU1P9h0tUqiChXP
t7Td+u53r9Bw/LLiocpa/jT49gCxhPA0htHj64gbiLz+CCbI3uEGBLrnj2cojNXw
tf2f/JHnFRwd2Yql7gS+LS+IIC3CCb9xZ3IOEcJcIC/9vqoJ93oQEVo4Rx3ElPC3
MmMn+HWSGsBNaZAh1FYPSAWkXuyWSsFALqc4J+lREaEbIFvRoMWhLCyepKCzoeIl
Kzp3MxPZ0+7HXUFrDCYPjc245VQzywclnDCynRvOXf2/byPpuBI/JVLhCPuWJIT6
Y/WUOibcKzB2+jLjNKDf470/mY8tAywglQyeapPg1AdR5wIyPDrpMLXIsijSsVYM
rsGP76inOnMS51TXZjkkKQqazXtQkG9Amap3EvujsVe7ad2jPQB7b+f37OIqoJPb
Q9hiP46nYCjgrio+/q3DZD7T6J2Vk7fxRIbIb6e98u5PGe+ushwozUGOHowMIAtn
3Ud1WNWDbFX8loOLrXgqBQSJJ61r5pDLboR377cx7ZFf36sgA1Saoqu/6X0CuUGc
eyxgdXgIfGapXIhvyKJEzhIc3v1HOQDjldluFxy1gaRASxsHjiuphpl5J0M8pGSZ
Tigdq3Da0nDCKCNf9TAj0ouQZR8rpEeVG9NMS/tPsLxjbM6E5sICaqNh9EZPBXrF
Jxx59u9zbznddl7NfGEltcEKD6HhKTJMqLxfEW7S5Ur6OTI3dtg4e8UIEUxb0pqd
io0DyJsZYFdUbdfKv56UOXpkfLI2lc1sJz0XVtxm4MsyUzyleTatAbZNzdinrnn+
SuCsM9SEx8L9drXHv7pQEVLvpvc6KwjkXs6Z4L0aoYKSNoYLnQq4Y7g2SGAGqHNg
MPIv99USaf+ifLFDtgznZzguA85o47goi93WmTBgKcledIw1FZxreiKH7HMt1G9n
PgOmkn/cGK0Ho28XIsNuXp8cg575V4UGnBpm+rjRvI2fXecsbBprrMts9+2NMiYl
qGxQ+yMM00rxZS/UHo1JmVTK5n4QzmdRh+1xOYP/Ge+hzinjv3ZcHzcuMu8Kj5sR
86Im37t0q5ZlHS2yVtn6EYXToZ4DDJM2PI1nhRL1xO7r8zaEP1aTbdDpJNftr2wH
8x4OSPL/dLafWcKIfYBm8Ws64RJiLy1e4++ZgKcuZGZmr8QrogeRZoFU0OZc7N+0
1lC9tXFYRI19vf2lGYdA3AAnYnxtBKgvQi9lWdF2/hpg36qmo01NfQXY0M/LGfVf
Lc7241VeGrC4NYRkr0skp7EzdMlLB1Vswg4S7oQG919EOxe4qnaJKOsO59sOuN61
UY2bDV0eFn8XgC7hpxhyEQxmDKI8n7g0Ui/6Wr1ZEjSMsAm/GOe5azKde0TP5prw
1SQSZqlZSGA/e+6+1xYkO2fIqTA9g8NbW/GkBgM2PPsMm5kTkbWLEjQ6u4tWD28o
H77wlfTbhFIeOFLVaG2cSLmbzqCD+/0NU5UEIHOVlJe/5pfrvI7VfQTnXLZDeZXr
GJdG83mA7Fpnq6+iTB23hiPUfGlXM+UlbIxqO2Fwl/HHdouhSVPt4x0FZXlkjyCg
+w0v7lBMMua/GeBJcOAm1hGj1u/njEDV7fRvRcTccDwKceZywJH41xyZq9DO9vHT
eXI88ukB06fZxSlccYhk6EQ9hOe+nXipoJtNTwJfoZq2BGuRSc5Ww3j3XxOrMOM1
Zv+Sh+qT/cI0WfJsuYMsWVxTJrCS1HcUcqQrCNCOhM66loo196AiuM8oonFvCfYE
TvXKOkmIt39zi/ptlvqxLgQ8xRBB0D1PzXLUGg8X3isL2xRO0YZr8QlsPbjGAErg
zqA5b8x33kjK3QzmcwC+cdUhtg7gdyj2W8PJ5bDOIm14b/l3A7/OhKRmLVwa9UqZ
a74weJPYHkByiB6pu5fXRBmlKmymXekhVwZMZYgnbpkGjusj7FdiHOw7yPYA+YzU
pXOCVshJ/L+kNjN5/sat4mwHqwcEuRwPSuUpKRtirWGJDSnYQ1CFSzyXuodX+Ysm
KIscDZsS7mqFMoig4dOGC2vNvzcw1bRuJbADnydEUBZFd8H2c0H0kliQB5trUlMG
u9QCHg0k8sclw4uE1EHaG78w5Be2OToI9Qq6Up9ElOWEuRxZtPlcp0JE0/R7lko6
EwNgHo2luJ8w3posDiNvEABjzEMy0/WEGo3QbtbHlADpufHu3/cW3DdI8X9XOLGa
abYEoW9mjIYkw2ttanbtcnq45b83c9Gyq90aH0n6nMlJ66fKBMy9Mq7oMXcYnHxd
Fi/adxaht3y1qg0rViqetoNo2lKvD+iZA/XTXcEBcGeLo2/vD5ZK+YFsIfjiC4pg
ay2cBntx0cv2FfU4hVmNUDPEQoNXunHqiAIiDnoBbdLeSuuev16kJ4iKs0Y52tl8
4Ex2kg6cszu72N/BeUtSFcoTxP1+uLhmGnK/ho1eBLOFSF3HPz9omAHKgM0zRhqr
mZagbn256TQu2jTaMALuQ75V9BHcAXYOxQnxATO8CUlGyi1sexpmhsM3LCh3HGuL
ka5ugDHuDRQTYsw3Rn6jE14ROLK6hlkM1vcgYfAYW5k1s0NG7YQPxz1IVq7ver8l
Bwgy4IQf21+xFjUOYo9H2gwdMofWprJ88LpMPUNLNa4prFOzJc27OlHOlyGVcb7F
JmxfiNY7j1B64TZU/S5umAi9upxD83CuoE5Vbhg22n99vNHqF5eZUSM/w+tC++W8
n0JmKUexhxNXBjoqlKAEGUh4DvaK1w3wg3Ti1Hau6T+Zey3mr8R6DF6aH2EqXBDO
7MTn5tIxjQoHZ8ToYb87flH8eWxU83BgarxpYIxIXGZeL4fMzS+dxsVZbSLvDZ+A
q7W7QpZQUpjvCJuS2V8OmtR0xPQhLJzljzIOnC/4epbb+qIo2hH1v7nrq5tNnpDe
t4A67UfRRryAEHGPLNP5a3Y7TiT9H3oY2ZBhz2EYg0V7W0Lo/4b1DYy8cs3xSOez
YVp1XiaYg15c/Kx91y6WT/3hJe+BHoisdZ12EBqKQy8u3kBNDZ6TTeD1GfwbvFhD
IRTV3davSFGb7QljdPbPAsfB30lFHlmCuHquQBp2reP57vVmmA1YiZigXauGgnv8
NDToxu5x4Ki588RU18xmrN84ONOIVHW05k68JqlDZ2TFuT46DawZXpEUDPo0rFAW
2oNbjHAOM7YogmLlNVFMDwFCfUdNzX4mtY+DRYRd/6Q3820EdC43ng/GbeBGWeED
l7z8JQRornsDrAie2y9taMQ+nGEB39pOSjwqeX1XzXWJE5ADuSy39SYT/M2SNi/E
xFgfM4NU4bnAId6PODtM1wL2TeDcyJKy+iDFyE9pyi1wNuzrArxwpMvdabeMldFP
Qv+B6+1HG0MhpzDsl4HtWUmbWNsKRxOJ3EX1K+dJI2by1TVXINXZr+M5/0qBg+eL
Xh7GEwa5vcV5ZGdrDc3zzhrzo+GmiDinVH3CY4nDsqOsl9yjT6jlJtQELJIIcCaw
F2kM4D1B1eZ4gJB1Z5nr02h9BzSDEp4IxUcCRufw3pvdH0zi4YvHpaRPdBJOjByS
n1Fn1zJfe/OSGCBgFJeE32mg5zlDT8qpUB/0SD9oSYmcmfGhRKCXBnr25Hu12+zu
azKsDK5npVfaHzxdQ0ULbOj2IARUShq2kTJUsGnxjpGPr9lYeBB/5TpGfmxENgFB
rqGOGY73tQzEqq9Fy6nrSKGIgt8pIr4G12U6pQbcED/L20Tq7E28FIZYcPo3vCoO
nF6kb6QEKilaX9wk7ovqOWkI2JiDlpRBjrhnVtKewk+qACKarLUSqSYPlzMJX+IT
MwKcNRX19ZDudF/e60oQaqkfR7MEo6tiYj/no7AGM9HomK4pZEqvI/cYlUPdF2yu
h+86iHKG+mSWLfggCzGr4G4wCZfgmWzf7MGNH3MW2dGnsFyjOkGUWm27Luom7Kpe
HIrZLYRV5YrEXO0faJfrpcOLr9eWB1+yKgJBcxQ1P71/mS8EP5uWgI9dPa8GpJnF
6UHXfay1gskK+i9vrYHsqLxQeWLwnyzFbLgObN+6J3C/0UWonP+pPSwbXd6keXS9
7irdloPR1I6abzuOxD8gPQefFIgjvLWOsGj9hH4Y5lAYD8fghHrFh3GfOP09DSq0
fnl5Zd1wemIB+fAjfgcTu7XdBntnxeLpMBD0O24uznT5UEmMoiMARFGlRuw3VskI
f+qnMpFYk9NzRqdQUL00C+wGFuJ+wqaYIjsq2ygYyb22kOME/hSRpeBWroQKnFav
cePttWv9e0TLEPOgMLfdCXcs1SfW+AQ278hNvL1Loexl3P6cm4LDTNfK2Td8bz4K
Wm1u5F5mn47Dr0C0fvPK+yRTPh7XwoFhlmyzCmIkUKs08PXEscMxMA602HdnS2HL
pOs/A0ajgy7ydUEWBx3kcHXNlaVBUPw2G4MJEh3G9PowTr5HOLeJBhpWppthouVD
CQw14vrg+SOMbVuJiCjs7B0Ivp4FWA/Jv5uQJV593a2e95Tpu4QSm+amR70GH8sE
6u7lrt5Jh3TfDI8VAGCtJANuo4XblDdDxKuonPYssmtISph9Cj8YkKf9p4yLHhte
9brC1T7VAwyGM3h/SxViI7o1qpU1M8jw9WW3IZ9to2cKXrYUlMkY6k0ZcPHgOahv
0OjpH2d+j16ZoDSjvDpuRNcd78WmcuUVFsqhrnhiptDQRGtPOAOqyv/XB1u8y2HS
eXG0+NQjSVpxATp51qV36iRfNIvHP27rzqR8bJSbiyaAhZFtsAbpd9T+8y07zFdM
f8FoV/QHA0VEnjmdj03of06X/rOOlTCSmkUMaJAP9yOeXcYgh9juCpQdBY8ynijy
SaIOU+V/Gy78MffDPTjqy5WugbNPruZRcs72FdufoTG3EjWaglajehIUMtiZx6oX
gsrE3WFIH47SsFDnR23oeSJh9aqvWIJw4MYlXgvGwlCp/HPE1Ugv2e3nZWP7wGBC
e51U8G8nwixdPnWACyjtMa5Cy+hVeZrEHIml/TvkVolQKKK6btTpJjMVslzF9Ncl
S6q7ZkSxzkI9dQ+T45HIkclTy3K7rqdXFHSWF253KYJ+HNsX7RtPyybpkvSin1L8
nsbB2mYGOduX665sMgQOU8Pzpg5rq12Qodv1wxckFob4+2bAj8wp696MvJrxuql1
uilYO7nxcEIt+wbCdlsqhPq3xh8R+Sb15qbxkWw1DBmOwnFEOnL1hcvRfBdx/Ffi
c1KN+Y/29W6AhqxXsGm40qSIazEpXsL4rhnLRQCNk7GItVyKinAsCrgv+e2c8uxS
O6Gs3pczNZRh88QycouCQAqkiPI7At3kBwnwm0GVSmcQMvBk1h54eyfKPPfCrKWa
3l48WTCtmVfrqOBrkN3gXEfdC3qpUNW3vgSoDWvlrVwbNEUsbmjdj5GmCZmX4KFp
sRt4W94JYj+0A9irgDbjcS6ytXxYp3rdJbsX8MxF0uGBb8i34ZEvs3JUgImsqgLk
umGamoWLyfsvoWpZMojcf1VjuDQCu7+5w4RNjlqfYtT2gBwZJHJWzK/itb3HWwea
SUWO3b4TmL1lWrCG0U31FuQ/vsSCUKd9hn3Ez4iMo+GHOjneqtJHHTVgwuAB+Qwo
mQz8E0zrqAotbrab3mqI964e3WTiDjkx15zfroIX7OeMeU6Y2o4u7Ywsdugq2Qxd
wydaIKgo8Xw0pqsrws5vtbte6s920MXNTggDsMT194ay9aO8AnGqszrsYba6npMI
Msxg7+0rhcHDo1ExjM5Kv2SbAWA8KpQIxSAoYofUPz6iVDMMDLVzR94iLPD1zpJ/
zEZq7XaopPdtrHVP4XdGFZ6RDpSqBYzWBiLncvofdlrJT9vooq0dTLS1ptnyVMmX
8zfu3eh990LDU6edNi6EfUEz+UGFo1dzKg5wwWsBM7CBH0i/AN2gb49bCKtqJwk6
X4rBtfX8sT+0k3yex9VIYUT2y/G6+Vx5qf9RWpyofNMl8XvgubxbrYHA3mCIqN5I
ghrG2yawBxtK1bPcLMIPLqP80kp/Vm2YdOs3kcYWQyX1WUzkq5XBVZEqflkiGu+h
502ZaMoe12FhyHmO8HNc7dxacROWTWNGSzZI4kDgCquJ7LsUlFM7IsqqQf9pHw9K
GFu+CUsNJVqTJLbZE+HiBEuuAQLebcw5Tk7cZvu957onehX91lUS0/Okc3+XcK2D
6ro5MWxh9zgyCwM4DlWvoNTXBJ5Q24xUqPl0Tj4hLcSsoSR7vHZB/a9LPc2LtwEJ
J28kZ+QcEN7L2dcgf1a1Gts6TaKx0m0ZB3NNI6uikM9PEFF8Odk+12VMJ2rqMuyW
CuRflSm7Ah/eDtsqv0noRmjoduURh1HF6jr8kWUZUmhXEl5+/4KOyHqg0S4DEAAE
YPDUb3XPisDrDA5ze1mRVZdCnM/1VHodY+y6kzfLK47B+kU4H0ufyiAUSHo1XcO1
HvRScSudRIGX3xIu33aEg884oNhwFNPw4OtM4H1P+/fOpPbgni3vQVmH4vkvPiS6
JZANGwBfoP/xUw5wRrmmUYtaVaaR0p6Sm7XDp3n6wNpcYQsAh/wHrEcMnQZHbYTY
mMVI1DYC8iAyF9Oh5lYcts2t8CmnmdoN3zUaeNHE0alHJHhXuaImadUXlfJqrlb3
89Fe/dW+M5oxE8ZPLI1N/xRutCSHb5kMMkdGQD3uiyifpVShd8BMH4eVOdf4Vo3O
bqdUb0oklbpMVATF6wTaUXdS2LOmEqoQBxs4m5hR09zshJkfuoPUJCEefpGGmdSk
cgwLZfvMDxIGVmk+2vPpHdlA0bhUjN42kwzrr82HOpj0DnI9OO5c2CP1hyJ7mM+J
8iv2ZNfweJDQXIOrLOx9PG2OK40VFhUfTPojrAffS4RnxDEbQqvvZEfLdOwD3oEk
WmE1dPTneMwiBGoxSApKi5fBav/ReQy7jU7qeQk1I0HDSr/+4LXCRmBBDZ4EuZH5
KTVnXYc3F/HgY2HEUVjM11GyOelyIO5RzX+UVgT9kdYZq4bFBRMiWhhbQXuh2FQ1
WrmU8CuoxTah/XeoI4VT56kaggXDAWAUi0fGZ9CIMQtINfRe6pMmn0FteVl8f8P2
+kPOPlPquLiNtBT8pK+ibjSnbnuYD3+Dxt0ETbFLD0CcssugvMEDlwTxi6L4HDEr
8B8E6wATFTy42ZI/dAccLDUV5wM86YUr8yR0gkhcu8CN6adxw/3PDE5U2wg3biRM
7jdXZ46pijSNe/93mASQ1iBXJvmNDaO6eTSfAtT0B4FnNqvL4h4atT+7qQfEXu+d
5uO9UZkC24w40jQ9eKOPmef2paDrRvE6H4EIgFMrZwcYW5IaswMCBnnyYj192nL+
3QPacTPIcvbuH0TPlur3uYYhZwP6Ubsj4OxawNA7X7qeG7I7k3SC3hNm4TcTwmqZ
UVVGrUmym34eJ7nUcjhtSjQSLMnlsfCYmyonoAxx/IFZsCzvLeu49MZruIrc7Jyk
+CNRpI+wcZ9+htaExNWdGt8yj3jCqVoTRuvmh+luQFaUtN71ZrXbMt/Bu9jqdmBn
`protect END_PROTECTED
