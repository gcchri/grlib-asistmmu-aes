`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RxXzkcisVQQY+92b4O1HuN7DMrEJk00t7axQCpcI68cQ+CFGmyvFTfBpFVg207ZH
RzNHpXOmCZB+OWKFhKRaHKAxGwl4H+a2XA3/maCmVZKpOVMm3kTH4jj8oXqAALHv
f7aJQmnlF0OisYmHmfKP59LWIoQQ3VZalCIcHZY70GjgUuMcRTU4dijHwnk1HSJz
j/wwW3PuD1EX37ciOeicEOOFOVtXeYBx6V3uidLxZGzIswZSSXK/IavnQiis7FQy
WoMsNURQHhdKcwHRSgRYddZMT3qQLY/4X8YWD60fZz3/zM5SKOyGJGV6wWM1/Hzg
PR7Yf6OyK9mXB4KdI3FN7iFRZxxlb9AMj/4uVxXT3Dxcc2Fcar6vapLOnpFDhAGS
uoKNmaE9Tjj6Gas8jJ6sLp8D8FTb4tH1AaYybX79GLJal78TgjwFa+8uZGl10vCR
QG9cpNAfV3VobX9vPfcD77ddmmfZ735lAhvRvUQQRmKDGn04DEteVBlU9bqAcz3a
nT0otfiwpxKp4O4/nTZR03LpaY/wmzJe7WDIFv3Oc+WIPRsJH13ZWcixkxgKHUxz
ldHuo1cJKX67Nb9AWRcfGqwW9gRstrjdHuJ9AL6KDxoTzkhjgduqAUt/6C1QeVAD
8wXyyUTS+PHJMgEpgZklZ7AzGzn0qqu3uqWxOPujL/tiJ4Js531I+mDxRwbOk6xi
Rmk6enlVhEs025p5oDsTx6FA6Bq3ptVWSr+p0Ygnyq7W8ZXvQNgPNDK+HXxqvenq
bHSLfxvokmps6mEYULcpvvaJGn4Msx8Xjx9Rz0Po2NbYqGszZjMatK2ATXo+CyCo
szeR2Odw8TchvxwZyiYBrPJx77y27XIA5VAzZjSlCDUB8Mo+Ah6II2q7vY0zpw8h
eTV7YI/cOhZBDNHkco6bRMIHrhBGgkZWyT8cjlQ/iX1RYDBP+f0VXDKKFj8chOo/
wnbsFVKtyQmPHp3qGuUyQxv5lP+Hf08fG/oCn0Y92L7UM4dZEy+KAI3I0iJA/5gT
NxpIeviYbAORZ41nzLz7Ch/83wg1xseEkT+743Lppjm2kZnDUSQ19xughfKIdeH1
ySAg9A/gNg4miROxQOtmKmYHj5H5aSXWyqxcpk8rTc8BxqLceyIJdIjHveALXl/j
gx3/aMosPE4lPLNclS9KJVCxkNiO2fhhMV15ljo9NrsNeiCA+AtOd+LMQzvY014P
4nZ3WXO44HQlVAP2TgQ+7QzmjqwtF9/Nhk1v+AGmLbcNEecnLVAPkWORiccpvKVV
+FkP9JkjFSJJvunkNL8rqobx8V1XdPJBy9kUSnmDKTKyOBX3kW+fLjl3gTPyM/5p
AQVueHR9apGBsETvAT6sS+uy3PPy8wM2TV0Ej4REwrfVLOhhvnOJ1WBCNDec6Xkm
s/aX9vyJvPaoP/RCaFSySsfUSDMPCyjgI8RaX8qh3SNdYmA6aZRuVpTWMe1notyy
y7D19do0mtqrxldioS5923msY/ebva/YBqP/ztCwARjGJE7gc5RyHkHyfyuKPURP
KSzuswcT9ie10cWJ21zaTGLTeeWoNmYjKVpH8ldzS8kZ9ZZZ7HpbTCPaSWTOpOys
IGXbCpUvgivOXq9dC9ocJ38+ddBjcSVZ0Af5PWn88Q97qz4bBR88oT/bT9Erz8H3
YD9p26qxX102wO95Q4jo6Cbo5Bh+OuXrihchEjLEr2mIRM2Nc8pVEbNzUJJ0pp6Y
qxE/o6V7FV0adAKnL9qoU2IA0wp1+exhbryBOQC6ke2ho9SKy/QT09TgZEgXe37q
Aldove/Ul1uhRCXIpTPmBMEwipjMZVk1Gwa+WjmuZwJiDdYwjo9RTq5phTRiV/9N
cE4C7QJZcJ76fwKw74pGorUal9sVMAvsd2aThBXydjqSbCKH3QWA+PGxaGWfqbM6
JVbQc1HQGLrCIq1uuv+A8ZGDFhcRDcEKNssxf1jw0i7eSPbNyBqNeH6MB4w3xHxM
ami8cExGV3k+gFHZtpJSOXJkMVwaVlfEYViYM3UwhKuL7Y+SKXGiVRAcDnpjPCPA
T/Uq1wxNtzzyRkVM8LmjOY070V3UHhOUgvt/ys+GzI8ETymQmHJbGKbRs6uJtirp
TlOFyEh4P/vjT4dJTZT+ihU42zIyOeKb2P+cLJ0o96FU5EWUtwyen3l3s/YfmeDH
KbIgatfxHwt+NPt+RnroPxIpFEkyL9o0Xp69GB5z++KkakfQ8X9VKZInTTHa6gWj
NVhgacMOsbIDyJ1TWQy1kJituhWiRclPKxkB2QWicLNxiZzdpH/l9agdcNIpdv9e
Mc/bRhYci73R0QCcpHqFDzuj2/0zX9hNruFfGuVSF1XHhci5xW40tx6KtLZTMIsW
TnEyW4ywtQzRmhi4zkENiCkcHfSt0iIq62gDRnKjmfFaDj4gmh/7X+SyEBrITOX7
/SYAPqBBY/pb3Otn19Vvq9tUe8Vau75B5oZc53Q8Jhr19lto/DnSUztVXydwimhN
ARaczrkGFJ3JelQFWCMeGQp8hqhNNdFmJ/uS/9TOAQdgMoZkvE4hP5OFfBaf8bOW
8NlxhPZGUE2YnMwPAmRTo9SesidHINPfX4vvZlWia7rNhBLZyiPECy0pnqIWOq6L
kSYEXj91LGc8RKfWekKtAhY5En0zpfVXLYz0rc4VKrMYqUgb9GVT+qYamex0HZK3
F3vDGONjKLCVg+vSd/JPOEdZ1bYcF5ioC42wY0IzMaE0z7jPPnPwykc/1P9LEKJo
XKWhoiHiGnxPs//3xnoWTZHRbIbpXeUQtheWQ2LCHMzzZPp4Y0NAvhIKyA9L8tKU
qAVO/9WQXPiELeMn0lO3RMq0ReGGFzfyCDzsWnw0hBQ=
`protect END_PROTECTED
