`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EV0QjQMEnUqEFnh8qY6Q9BfuHLQ1clN4wK1jHbC5V5JAPD//+MxOu+RYOk2Bg2Dr
kS0Hh/hqGNV7CiE91wlciL83cdeJplx4dAdQjEchaahUTirwxL7qAffs5QIvwFg2
Qkb20Zny4Uew+/1DCCuj4qr283Li1HSglQwSZLE/+pDMxgLqUwFpvJ2bmmkiXEKP
pCnM5Xh9jzIZtlZhhSUDFzGSS0siZNs31mX3jT1JdJkjAZGbSYitnf0+Kq1rPKWC
p0mhuWCWZWjpqCWDzSSmoe7VnkCpf4qAPgEjwYnLxT0=
`protect END_PROTECTED
