`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AcDYQxKRrZViIIB1yoalNsDu1igD1OfZ7eh9NU37aySE2+mPOghGKtybgOzS03Op
MXTnnWoYoyWs/aDoHx0XyQfLxv2mEHED+iEE1qSRDOjsTs4mAhBhlXR8QVmAL1ks
YDHm0goN1tK/irfPnfGLSDB4MRtIOeQhjtERc7GFFfWl4jD35GLNNA0Ok+6EfRF2
oTAn4Qe6krhXz+8P9xspq1mp7DSifEFaRtpRr8oKn2WnihZMB5qfTGKtfJgv1F3I
VXLJ0qhKhhrnp9lHECZ8lozTdKpTwkLqrIS9IRnvXQy8cEw62Ul4SVvhR/qRvubT
8afbZxv4/Ii/paFjuqG7/oHzZTIWd98AWBG58m/gC13WuINex7UMF6Pu1kQDcayg
7DX1LxV2x+Folo5AOb0C50SKxKNhlR1yQTURlXOl8vDsBWGaTAXhaieGBTMR8yof
2ibfiFXxqtiaU984+i857CTbGhVIVKUGmT4fozwobITp5+o1iJXg1LHe4XQtG7PD
gIRXxZNe9P2aGfOqEUp490IdSDBxInJ4eWvoRtaTuwbqIqfLaFVHnRTg7L+IpZSz
MntJlY4axA2dnAD6lWfk54YlBRtGEkOMfNVx554n1Yb3bRnTZl1Poj7g8sydpCQA
nYEfcpatfprX/qTPoZ+dviKT54lVSPlritFFiByxt80=
`protect END_PROTECTED
