`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TzTM7LSPvONHwC1DKeGuQ36dTKeQpCLCADV07tSEN06uw+cjBSl54Fang/ylMOE3
3piP0Bkbx6p7Qt1sHQrguW/gdhldQ7Z4eH8kh0ZCknyziUsem3S49kvmrrxcW4fH
gwM923pAuVTjyCgA7nIWBxYn3+vcMICVrAqNnadXSqQPl49OEdWj+7SdHQj6yL2Z
crMgdRJncmb4HXL71DaRHNuJyeIfSXEVv4+qwvLki2ukyrI87i9iHrSSOn1VbKUk
bOGKXGO7Fia5Ns7NOZYsgtLi7+QUf9OY2rba9U988hpE6r3NiT0H33NiPksaA8Hd
WNkARBQ3mOISWgJopiEUu+TESeaS02hZpZepgNNHJq1SWn+khPJt5CSZz1tONd3T
NO0Un65J0JMXwtnAxGDZ2SvNnj/W3znHT7ESAhfxsrkCIJ8DJimYKyYa4c5LYwxN
QWkyuEkgTorKjLyIcblKVjKug4/Fc5a+kPW0j+yiMwnPxpStvbLJLvwpoZBMyKvk
vfPYQ1Np9Bxxg87NbTVTgxw4u4ZvO5eMXheiahCpAJ7ra1rSdcOMnMLS4q1zgsv1
FgJ73fDFltO0NgGasYj1Wdwb5Tym7gmJcMsXOUy9vxw=
`protect END_PROTECTED
