`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WdmzCVfZQNkOAeD/9oiDpeESgzV8BNZYZ7OluvEJNhAOu4MQzT3sFdJcmC5xRujM
VSpWCRFmMtHukngQUfq6+syYRxkSs1eCfTggIN0sEmRITdDdH2mKEFhjh2vfIMnt
bWVBEGzAojtSw4HuQZgQP9mziWuIIbjzipyNKz1lfkwtDtWRXnDeP9E4v+kHHUmB
og7zP+IjvdZjQyZnglIIcHQCWsf3EMDG6M07syIAcA3I2WAMC1s5RaEKnuGNzY4c
MIEvnPwVc8WRxRCbZlSCigNHXOjiCY284GdvSZ5bdeU4i+sxZe2hb86zZApcwAes
3qQSr/pQ+SBF98hPemWiQ5kzLw7JKivrLEvBl608rpD+jBvW5bhyFlO02Lu4Pq1P
z6vuyqpBseilWCrSjbhOE0/BjGJm+BwssS3wnUI2JCuT7bv9utp4n7+vZooJJziX
ToxwOexS9yd66X68kaXMNBuP5Ki+9iE6fnSmeqqP+b2vMSaRT/+RAuE5MywZhwEF
2BRxXjomCqYBKlOZ8HtPivfWsqsfAYC7GYZ2cs9ocRo3ca3i2N5Z/YYIKnX7FEfe
t1MF0UckZD/COV7b8LhWhfiscy4BvrQJA787GEWvNI7ShIaU8Dcwi/9Uu/rI2ySU
lH1EStrXZFk6cyDfXAZRBj4x5gLyI9tt3YqKHs2MGNpR/WxF4gt+3ERRZh7+XBGd
dyViJlAcWpkLRncdGknkI5QN8taJL8v0mL8fBBb7AwMterZ5AaC9kFRR9CG1VuFG
PcmSR0lcTy3cyvG599W2ox2Tq17xvwXYlJyfBCqWNHKOOBZRwtPqMiaesIsWFJnh
oJZ/d1VFt9RnqBXoN5NbW03x5Xd0bUwoBukVEqrCaQVSHDXAQumEW+Ng2KxyZbtd
YJvtVSUowNUdolSm8zcHWps0jZHKadF0tEzxAK3LMnw9uSJb5Kak/lXPqj+u1D8v
WytS06fh9EF+diWZePPtMZcY18ZoFomg1og+lx7ItirnsSMzM+M/bvhCAV27PW3m
unFZY6ID/WgGn3xLzMmqevphPJGkPjv5QWtUNCmwukapiRGwfziVhEuMQ4A2LIWH
PQWYbld3qSZjmpf9JdLlVOOkEuMKH/gvjwvtorLM4pMW3bUA9Tn1LpvWo2HFHDk8
rb1Qii4kzq6bX66B8SQP9qY64JesiSSHyUIJgrJEcFI14/El9uXSlWHUz8RXLhNS
GbEoi4smQrjY35GuqibgTx9/BusQM4kTRcEGiLlAfVDxXIj/zMsa4cwCUJSZ75P0
8OJgzxgwayhJRmaBdYCyGuQB9Ioic0LKf1+NRIFYLayCVFSL7ewzEKwNQ52X4q5B
W9JtTtECVCSPstAeF4RDwEnskBI0Vhylg1OGF+O6zNHYt8/XmQJH35laAgzxhpjR
sdJ34h1mppUX1QT+FCWBb6sDGdGTdd+ifX+ehMCja6lbERx/Mhm/IgxzAzVesbZD
X5FRborZRuY7RXOkOxOcbFivoivYStylr9jSKa+wtEDQ3CfOhS7LusW5cMRUgnz6
COodRJRMGHbx8uOUR7w9T+T4+z19vHPWWsu59FO0+lV7+7O0m+kZKpzaoo1JFPIb
TWcXs26tfn4aZRtmNeRYgLejbR1anVtuk3YgQNUhD5NLo7rKQXL0IPHxPlbAWMVI
kYibMzAT2z7vx7uNJkBuYCQ7WqWu1LYnGWIw5TU1W3PRwNSgbzo94PMbF8NGYmcB
WcWtDCd90nyZ3Jxa6UNdDlidZzIXKedxj4SKzLlwJBs1KhpaSI9tygRTRLdIMANZ
bGcec5/elRndoU6D4nmR8Jtgz6jpAcaDUDKfGvGM+rblEGdkabt1x37Lua/OwJRz
jDx+PPateF3wKrMH1ua6tJ8VIFeqhQVpOULtf4QM2pRBlvFr4l3+egS7n42b8/hl
WV++SXTiefKrbbjGijGvJ3yySIvC6urCcPM03cWKQNzCF/MLh13LfhH3LKoP+sSs
gdr3k+2LgiRIL23wkVUYFClmfRIdhiJ/kWPrVBhJfPLzXFlel6oIMSrUnpsTaIvD
ov43RA8b7rvy2D17+OXIFXwbEr2Zf0k09fv+jU4X4qmUx3vUSvMM1hRh4bvyspgB
paZ0DVXFgdv07GYJdDfgfmPyj9UakbX2+QntYt9oOjU/F2Y8J2Vw1/7N+ijQpA9v
axEkaeUk20HU30VFLlYflO2/mtdnvCzUCAnqTlZD0/L8q8QUKAkBe6icOQ9jvu7f
VnPG2p0JCI0v09GcULBMgxCnixDSpXPdBSS+XZlRvFMSyoi3Z3oOQz+iopg25c6Z
CDxjfjgLQVc6UFkXWNgUH/Kt7olBCEorahpemi68F6bQgdmdlRx3sliWo8fgjpqD
bOeZ4Elq1mnLXOKv2qVxx6COC98TENvmg+Rf6ekFFxROU0SPgbtLOXIOHd9pmGrf
hz9Tg+9etjEoxnwZl+hj4ZG6fX8Vv34nKN+i+Q4KVLYJK8G86GOjvNUd7NYVZ0mJ
6ah49vsloIZMCsOmmqAtjp+jAgPtsUOLiyTzFvBzNMnjGZNVbdbP1dMLWDCqBVIU
Pae2corRgdodcUvBZ5bHxiKCpJxpzOL3354x3cAhUA03qnj6yi6R5axEn2/BjBfQ
I2jsgFQ/uZik04pW5oBcTSMsQDCZnbljkiqL0Gvtm+I41gykAIjlfNjWaLWS1DdR
noR9sEjMcnZuFenmiHTq4QIDJjxMsEFR6VYfd/rOjMdtFBmW8UPtFkPkYkTuA4vi
nEqlpvfbvzgBwfdi5pv/ZOJan4d7AhVK/M6i8clmaZLgBoycUe/PAd5q+Z2bKrK0
nVSwYBqYe1iE7yFUfJ+E8gcWdgAiWx900ha5qf9GBNgMWeg5AMX6HohnMh5NjTVU
6bIsReqlJELPBmLSlfQowlSvMv7vvanoon6HQFzWJaRzuncyBFXziIqfUZmXtR+C
xVc6wB/ykaKnrVgCSw/qjJ45/WDUp8z3ahERj8Z1EDnUAG5gIC+abELf8FgkZcYI
gNW1ShddCeMguYDxXVTycGhRcGShGB8kg8mydOQRo/QHGtwVAZV7l0b77iChOkEi
eKstqvBbnRhz+h8EpwNARtx2MbZHLOLPbhclRMKhZUneMpcmvqezEBO3ieDRDN2Z
Zu69nUUt8eNGt8MGfMZQy2tq2Kh3N+wcyXmPbRCyKb6PrR8MDVoUWT3V1tAwSs5K
PcmPZi28aC8asFjXaJedjmcowsfY7e/MTli3Zti4bhflYkhCL4DvfYg/3bUR+LZ2
qpHlpFOpVPJDkOYFwFAJB+ROaC1x8FxxfKSAVSJ7YUS3OFj6gcFwQYx6sNCb4lZS
5/2pCU8JUWLxgQjUj9DLAZ1hsIYxkN5MXDL6XAcATzD0YgXlY50Qifs+cB3r3SVw
hfvZSl6fUfsivChwjXJO3Zj4pV4eRjnEVFPfdunMI0Eyw5BR1GutMc2o7TnuJy3w
jdPB8MNNVGcnnAOEdp76Ivds7Yc0GhIS8CNA3UKmSmUCgdoGp1Gw3beIFUMUgLC6
6nvT6TkX7RzyZnuy3THYifFUK3h+ja2oDuNQ9PfjwLDSiwjQRCk7zuULC0ZwRx0M
9GG7egI22ngqXZs3ru6zW0ZngTUlrmN4nfxHZWukbW/Ig/DmI7gzpEsnxpOFm6+p
4u3Joxq/SfXY8F++JLB0jgKwaVJDxjhj04EYcmWEJbZakYZoDdL8NXab69CRdBXB
JzukZWBP8T2nkKhtzrS8hD3D0zs11aAMZKm1P4z74dWwatpdOnEAspUiV85YSh75
bJCD9xzpJxgOa28tRGHAvlcQrOvJVWdkMzm+g7mnIAq9PGnM4PkBT4YYsZk4+5xW
iQHteXydxXxX/h+DIkXMtG4ya54kQEaJSQNc4sCcmiyYgH1NbVQZZd/Y1FR1Y/9K
sQLpzCu7oKZsEccoWxlM3LtRIVbsVHjhsLYLsvjB3KAJKPYc24oWusAMs/ohaHWp
Fm4+NHuTi8hmSwrH1H9CEsiDi3HcNSHzInTq7ricdW0=
`protect END_PROTECTED
