`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjm2NDisQ5Qs3Xb5BgLTiCdjSakL9z30k4WT3IhB9VAei8EYtwTMGKuYqPEey6U3
lBcw48VGwuhMd7TLcuhtwNbX+TiACs3k/Ur0JWv0WjbxxcQoUVpuCwhEY989HFc4
iu0T77by6tBT9/oHnKqAkdOmX306HhM1GaA2el9z9EZDcunq4ffSGYifdHA9dAYS
AgvgrjJm9O/A7IvDCpO8YkUMp9xjgTJbbHRlKZW43lMdlDqTBqlHv4nG4ClPz1mZ
GQQA/KWzmTddGfTBh1EV4VrzWcuAzPpA8wYivj+uiYwVnCHcUGLWJTvMPcBOC4lD
S2xu9cMGxgXGoxuu1VMEY6LAaEmTP3QGhEBD1NpAqRO4jF/OcKypoKuWmP+ybhQm
/fPjoDr77AqBsEFfr/jE4RY8a9N3A9IwowXR/MQgJbRU7DU/JaCwodPXISnhVEPD
G9e/sjNOrh0U4uvdjGvTb18VfsGRCeloZwZvvpRnL8uYI4sFr3rccRIgGuFAx/lz
o4fmvwpIo1Y4izoO4lV2qr97D1ygeTVOUyGICrcamSDB+N618cSsAgKQS8dPBfEU
dOZkmBJtUY8XcNZrbLx/2a6OFoGfozLEzTPy4bzZLoCslnxm2qHgrvmUAswaBX6t
uNUrQ3t8ZK4QDCA5Y65qACVKW+1uJ1uqSzZP+FUwAMisZ6PB2s4C+YrSjYQUIyQ7
Bm3407muA3eCoBKAG2sRGL57/3B6c0JazNtiBpMMkwt4jLjZigfIBjZY+8Why0Q7
OiSWmEYXwP9nJcvdbGcf/X1POpg1qTSmje3txAfoM39g45LSoXEso2+7CmZUWgk3
O0SQogcRB7Euz22gvywhjJWDe+rpKTMMOa4u75/msv4wiSYa+WplHSI4cxSuaty+
Q1r/nTq3f3zR7UUWvjZWM3djyP3JEqtmt0tDui8TaQqzTM9ph0cRb1mZlgIEEo9L
3X8ggeghftbAg2rSc/GXIXpWZoz0hlkSELQSUpb3NySqaZKmQXmbXo4bFQ9qv0UY
pDLwZteU0JdJhUEB2v7NBJnYEG4gLjZp9UNJmmWUZIDvm4ODSNrkjaI+dXYTMGoc
ZeHEgEkR5UWMuqrEM0ITlFv3pU8fCdhCEBdbSo+oRwej5ryojXwZCHpv911qPdrZ
/+G1BDddDSAATNEH83MAgy7iClDfIgVEsLxdOI9sZ/pZVtPfz4UaR8PsOfNYetOA
8HkQNX4Z9KJ7/EJlFHcps/UEUtD/Ve7MBgd67x9tDpDnLO/ShpNJS6v/PGNPqtEI
cdBi4/CjJl9kMNmaqF+XgT1sNsanx2Z/jnE/PHGuG1c=
`protect END_PROTECTED
