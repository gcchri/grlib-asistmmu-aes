`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ro3OYrmm2TqLPKVMPiHrvcATfOevLbQVmbClOTxGfSZuDikZwxjdwBq3uIqdX1VQ
Zi7jxUK04YZJ054Yt18U6so0QzyfVWLWbjuyau+p+8/kc6dVLlpInoGmVRxj2NEn
02dXlC1HwMCQOi9xAAbwbVv2fyD+pd+yhZVLVWfiG9DQSQ0C7dOEExgfT6/1GAtt
FtbcoD6UmnW9llWtq1rrTj4ZCeI2T+GYAT/qrm9mGQ6S/K7+CpblnNm9eDj6vca1
TxZF3KX4EThbJZl5MzPcZ9Vz4XEH65NddQ8pMskvRIIjNP/YlAOW4Dsnq/61+8hD
mhACh2cN9J0XHlEjblkzh9S14Ls4206jqH5tG79rMsqos0JQhRcp2zrHX0OR/V/y
cCu8vT8Bi9eoQksdMLL06Wbbvt4i9Q1NDEcH3fYcpARAUencUozhb1MY6DQbFEcf
DeAQrELI9uhNUmg5Sz9FHOAcnmruh0UqQ/E8Vl734iGoxb4VqY65pur9h7bqTxtz
KMLAWjsvbZPOVRfQoDcQyneIScoGxGiwzkQ6+nqGYUsUhXkkBKLrek8R3TvewbTH
/E7n8Gf2C8jeKhDo7Yef82iEkSZXIBIXud2dxWY5g+eGsrkgGCdF2ookKpiFjFkv
g5f19Z2C3IHdCiJBvaZUd/KUKSEZDYzM0lAsyd55cqtI8tb2EzdVPVKEiKgMjP6F
wWtagLP9N1PVT0RmAB+/dZLNfs1XJ3EBida1FkuKbFIkh/z1y7D6bmXz9pvl6dOS
5PXyLIW6ESOY+Ug9XICu/MYMTMcC6HLeeHmF0+Ma5r08mrLwRLsWiaMu/lK9S77Q
iqUNDjs/tGWRvpGd38bMTY3PqgsdlPyA2s/2SdKRtiX2Jv+c21SqSO5eZnr+H0YW
HuGHFnNpaNO5x0RBVdV0QRMJi7uH/4U88QyNheKrWyHxfriNmMBi0bdSOQZZaqIZ
yuEnOkGEEvZ7ciiUXUp2lEDdN8x/uFP29nPhT6yA8TSv4SOoOxSPPOunkdrViGxT
r/ThIepkPC8hrpHYgv3kK2hDD8j9dGXEy0hWBpAKv6CbURhfQxO6MROTU4H+Q/Kc
I8CEh1owA41Vfo9Un5yFyXqz7hmo0g2dZsbbHLWFVdWf6sZ6/IkMQLDA+QvYP23a
eSsc5WlSkRca5Khh3wICi0zbCq1ZM40zmTNSGTRtatZakZpBNq7tdk/KgvJt33Z+
51bVGjNL1XL0PFSqjfBTR3NruszLTtLc7NuwKieJf44ajyxCH2d+qIIr5sTM82mt
6VcOIAdKQnLi7FKOuYpPPdiChiCkPinZqH7x+2eus3ewDdgFIV7HgCZY5n9rGg8G
MusfVMbioRmXeSL32go4uS4rFFfx38ID+apqYPcYT0IcZ70yzfU3ETsGG7iiPk76
Kys9wIxtRCJnacjydMo8W0a8qKjhjYUGsP0kqt6u016LvLn4ny5Rnzi8KrMuCj6s
B5J1j632KPpyvd+PFVXAI4h1xUT2x2WbA/D1agUTGSQD+mgnzWQAEz9izM0OXOip
aUX84IdDCSbERUreURhTrNbH7LT+xUPTeiPpOoQwZVMYdWpsQ5j8dVKfldyKGLB9
w4Oilt6jztGm7/0BNjakzE9uhGsVuSs2wM8sXcTMrk3zfZg6u3kCcWXgylXXTchx
7niM0TLIlDfPo6G2gL+dwseSf4k1AM1kCmisoecK2piqKuVLUHY5e5fS9aZuZ1kR
vfR9N2688+6NQum6PfxZ0qri/I+cXYcQ1YeaXCtV0pXk8QLvCYDt3XTm3RU/ymH1
NC4WAS7xH5HUSe+MvGpbRVmP4mC2wSqX88pWj1HSRNgvJXOuGAjsraO9pbCosabk
dJ3vkeRkQiFkBgtFYb5Y3YUdhfAVKiRRpNNi00IvtJytQl53Ryxati0Uvzdi4qJ+
ZVhBTMisf+Wb6itKhbgxpxn26B2sgYMG20zHjoa9X8MmeLXj/oBFalS/VbCuY146
wzk0yRYJYYrDbyln1kTyMsLmVEmhmtQUqTvwTav8pdtPhjm1sNZhrJrwxnpBmIpB
PjJ0S7f2WzsNx7dj5aR2CqAJ6d93kvYe2NQRmZVeExVw1LLL8C4JuhkfIt8bTklW
Tyim2u71USGk0slJa0ukCLrawQqR0diDIrgrsI3+QsW7tVIUjHTJfWqwDrvvPX9N
wj3WBbBYZoZ2b/PkCjCkC6N0PTy0eNv4IPiMyacBDP31Dzw6N3n8QIRucMZos0fC
+kD0M/bB+cwbg6ZS7/UF/SH/DyHx8h6U7ksQQmmOnJb7Xhqf7Cq9EPFAKKPXvwxL
HiN7iZtpO8upnAkTKMM56/4hwjHl36hY0BECPeFbsYFAklpCmgnWgtfUCUxDeAxN
RO/+PxyLJvedk1JeSGHdYCl3x0g++l7ZcqzGCmVoiU6b22T9wW2tDKp+oCE9Hfrf
a6KgzCigUUpEWoBR1h3qTAzqPmaT+x1D06Xk5LOcLaQ6UMnOGDAmfZJLnz3kw9Bg
7RokUHfe6oquxFkx18Hm/8QkZ0hJmQzE+d/SZXA3orCg+vYo5TEc0FnX+LP2sawX
386Kw9A9JF10IfRBQIVtpPavz2+Y2nT4kGXIii34ifLBBqI40AFs7CmsZNtdRmJ9
5bNewTCY9faJw1Ppl0DRnSkMJgiGBlbXvKMKQUcXyEJE2gS+w96B5NASawisE2xA
/bCTLuFkQZjUK1bXSwdI5gISb6Kqtuqfzed/yMVcGkKYSkQj7ra8qZcIBhtKWD+9
+cwV7R9T9EC3xJCkrZNm5GSntm/UQsjUVCboj5BtBZ2nq5baPq8pONcmHZTy0TWe
l6wPV95vIc5rkaR5n2Eaf3W8SfJFUwF1b82Pe9qfCEqx/fNIL+kWPN88rM/R+5CV
p+DO2TITKY8iNmb83HpMxOKib4sBl1LpJY8m0tTMbvk6R97bIly6WdCyK/RezoAG
LfBEXvUfSorTQrlWZq8Na8MaCvlc8Ks+/jc1kpyj3o5pWqdonmANmDM7NHFQHcmL
hJ1ANUeDHbaOBedMdHMQ5pLfgEcxtZJz3jXw9TDpGXrtdMHceSGK7LBwc55CIPUx
PI5wDarhMIQf2CKDdrtZDissf9Pc6jz7Lt/lKID7oTutndTQ+mFlgWQu27GG1rcI
+e8qTj6iR+kb49SJBxuD9T6gn6X7/mN4Xhx+2ydLhpP/Fk+oy841pRFF14DxXkQf
i/hUtiQWsrh+0+y32YxqEwPQutKPAbmKKIuIOj8sC/Jr+7a5LXndzOIjhFe/0sEF
ZeXjOkwE4U3UZtLH/xWBsgsYZ1L++GkKbhV0Jn8MRY9HieNq/57otL4G2eBK5LMo
PqrSn0ykQjfsXHU/UzyK57T2Htfrfne2ySDwJGqJ3XWeyysGwJB66hao+5ofZpVl
Pzz00DYD2AFW+2TST36R1O9O28G9iDNvPOXek5wcVDOQonIpodkFUM6mEjeP4DOq
ZkIB9z+40ZQMmQ5rBOU/mGZA/RbW5y8bIygAbcpN0ij3uV2RdVsHi/hHFYItOFBe
FYP+c73Eg9JI/r1OMWZQ/CMniqbUYiXUJ0TvtIyMOyKv1pDxK2LmDnb0ka5GoWka
COf/GfvXC0CxbyBFngkFwCasiZYq3aXffEeLYxpU51WBou8V8qe2IYi8lDKpxOhr
v+AXLWo6CQ74aCjYP18BXwSKZdgzrI3tIx69/fUdOLDrPjuOSzanUeQaEwaR5aJN
7671yakM9+0z34uQ8u89ix8fWy259GKLARjNYyH5p0q1Fe/4lB5zYWS+HAqAF3uO
W6XWkgcf8GPrMRY+GpKFiTOm1ojXdjp5fPrDFRz8ObsMFmSkJ2mfLXiwmb8ottLy
qy9xC2qe8X3Oj0Pe9+vKQnG51Hv+5CUzc5ui/f3E8sUNwcOGPqydFauY5arAw6sR
ycUFgLJfLtA21UaQE6UDN2sSXgHKOLaAHDmsadJZ6c2GSKETdJfVdp7M9f4LOuFe
JSD4SO6T+g1QyHWfjhd6qoicYdZzIQYstdnMM7/7BygEqyOykCyeAxj5dBu1Bjkq
JcYRSdvADtqrzjTzJJDvFnMFhBqnJfQFAohNP/Pl4mE4TiRMIa3BGtVxJ4Iah+Re
wdbp75QN+3q/GBREUQ9sWalooozdRNVCFzcesI1UtS6PumFVvprsoU64o0wY1xlY
uklzQ4hL9Bh78hrAqjM+42vZGTc187xVPBK3DUMPeUoS6qIu8snWyB7rxBPIpRYO
H7kErif2odVu9JbOsJjFsG9CtcWj0yo/BNLCpeVlm2NPs+uY404O/ZEZ6KyK8OYH
K7XYkHcccU7T2XUX35eNssj7o0u1nBPBzqFj76y2I4Vi4BdG7lUOIWGqx065nQ+K
oZ1Tbf3grSee5io5HvFsFOce+L3rqoIBNoWITQpk00vqdM6qaHpCwXuFbSdqsKlF
fbM+NxqQLcR968g3UcRXUEjWjqdgoq2gohMZMIRVcjP4oBkZ5RWHV3f2jbaEakP0
DAa0vqGnPmuzrHvR2viWcv+x+3SToOdwXgZVlP0LEPQGzu2+2fGoVLQLFbHT1w3B
mnfa4vlWwtRpzMobz48f9Q==
`protect END_PROTECTED
