`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIzWUT1JabW62p/j/HngiEYFonznXELKufrw/P2dikZ/BonA8uC1Y2sscGkMmJpU
spr6dV/bCJyUET0QCDIaNVj7++lw5P42eFMTD5t50y9kCCqmfmFAjPahwnVyjesS
JyhrBzLCf2b3JThx8ST++/zW/fAAsezaegXVsK++pISd5/tb6+ENR41Q6LSsmjYg
1rMfvoekYi8VbgKOR3G9u1ut5IYOE1CdJnFSuZx3PuEygSLtUYFix21371wOjXAz
hJne6D8uGuQSv0aPvI56SNRk7v8aDkMhoQFcKIQBrG8frhPOhMTCjEAwlktpC2Ne
tFyWvHDqwuQ1zV8CueovxhFXpp1ujwZy1pB0jSbcCQ64C8ZxkO0qh9UAacIZ2H+3
q+HDl0BffY9on/N1N0AmVs51+VREyj060OJILfSlb58egYgbGWiJ60xeF3n8722M
`protect END_PROTECTED
