`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KMvV2TBYelS67GqIuEUMoQbqwBuKdh3JJds1JtdTKb6iaWwJuV+gqcsEoA2RiDuL
86MWHbCigt3PrLNpnHaI8ESijL6euyaAOE35VsMpwDp49Fp+jXZ/HMDDFWWl00Tf
BhA/M4UbZDvkX3+v4Mwi9Bnrm2Ys0H1d3ayxa3K7h+xvI98wavMS3RiYr8POYH/U
fIr9WqOXGTNqOSSKF/x1vkL+ynE14Q6w1PBpE6mlRZCp8b3ueOkla1vOnst3XVcU
3FqCi88lDZqp8JTajS3Or3vSqRYAhsmr8MImwsU6AzJZZPihONrWJ5HQI0eBpl1w
ZB5xHmoakJLXkA8OU6ftqiDzBFOd3k2V2qZmYrxUPs1PSCNYf79/dzatgzC4vbwP
FB5gWo1Eci6COM/jwfjc6ccFKHOv6J4I2H0/UWDFEOU=
`protect END_PROTECTED
