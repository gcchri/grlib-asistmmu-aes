`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eEze9OqsqzKOR64rrjUfiQUQjgd1yNyJRqUtySDOp2wA9ZNdazdQK+9bKMp55A3N
V5H8qhzYP9Db1yKYgwAjDR0UCHP2RGTPm8hLUMZ5nkWyMroRze3f6dtgj8fGIzAx
zqRS5KRtFZy0vXLCQtICvhrs843ByWeW+SgA7Gl0J/ttAeUSXA4DuRKiQvKPiS8j
/3TixVemBY0R9Uc9N28WDcLypB6bymRbsGd9LqtkyrH+zRg0G0RXh7pfW72gw3G/
OdGPilBhtTEKowS/qHFATf20g2CiToi12Or5URtYvEHF0nOZtXXkQMJZiplO8y86
kWrFTH4mZgOepgPYhOzvmRQWMLLnqQ5i492pHozudkwirgJVV77kjWFw08g60UwY
mzlgoRZAKTo5b+YT805Ko5D+iwhWFptp9rGY0jatueuUsf4/Qh/s5HMzItVgqsCg
YoivEiCPA71brjXZEbaDDbu9IX4RMNO5zH5ZCJsORBcObSClKF/5pPNUrPnkK75/
AOZxDKjf1ylLOQhZITKv+eAF+us/itEBJDR+F/tsvYRxrGUXf/V/JHEPvEjw5WQD
nymF6eW1eABHTHDcNpuKYA==
`protect END_PROTECTED
