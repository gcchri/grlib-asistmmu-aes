`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+TBvrmXSZXS8Bp2nifB39GsDQWjhG0ls8ZHqc/4QYM9MdcKr/0n1IBgvFnRoNdl
4yNqgePK8mi9wgLbwTIKGuUYnRoyu+gncD3aCrGXj3mEjgeRxwrtKAMrpA+q6FjT
uv0QcRyWLiiY+Ijzp2R1nbtGABQursnpC2JS9H4sndLDd1UpeH1wO85XYGrr6eyI
+Q04DaT8TiVOXzgy5X2qnxTZEioZI/VZe5MaeSJ0rxmFEIDyNl0W8+JQvsfiImIz
Ag2WiYFjjmRSz/F+fCzLk9FAvyOxVOpLFYJ6QbSjqVH4v644/bcw/gA5kSDNOnGB
tL1tmk5N9fir8vMgm2pByef/oQgf2VCXyMUrNqQersv5uDvIYENouvuGzu8BPwuR
Qy+lZAJu4Ng6+9kksmrUkGgbGy4UiuLA2ElH40UD/qwOal3ro4wYIhdsfxOBatrK
ZzpHWBOMVVBZjhb8ZLyiMq+JX7Vtp7BevhtaLjjmSRZXlsOn8rKo4iHmBJDpqUuj
PAOMPRbu47Y5qJdd7wGRZSz+vEKzQ8vMTlXbFFBMRCA9WoR5uzuCJTxdG2lngZ92
t7mK++dUzRzhVBHM9Qyn2Wy4dgn+Et/9Mayvbh3NMmBKyuskKFw2VWBWdIg5whyv
m+7g0gs4E91XVy0slPv4ZQ==
`protect END_PROTECTED
