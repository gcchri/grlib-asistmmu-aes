`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KqEgPyA/fZDDxfqUl0+kYI7iuUd0eTuKvSBOqJDBqPrnYkhNaMt40A8uHc0rccYx
YjDgrtS03Gf2MAl75ut4etKFdmHt8f3zQMTtxgsz4kSQrAztPkXoa7sQcUXl6ZQd
Y/yqJLmOjRi4TPUaa60fUb8LSlmueWmDqQNJvpl5JaNwiT3ehfCJdZ8ki6I15m2r
23II/6wMJVTMgt3IkJjAdiSii8jeC4lzJuDGn7LPZqosXeif+xi4U0BsYW3qmJVd
cRB6ki3FY8UiW0Rzarhv6a1YcjQnUgOrbiL3aNeCFshUqV3C/nC5PlqijamT4830
`protect END_PROTECTED
