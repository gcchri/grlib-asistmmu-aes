`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7GEveDQ0JrxAJYgQkUCGbBfAY4kMdoNpscjCVvgUMP5bmfSRaCXhEdO/kx9RFZGf
bo8j9awwrixmpfUvBM+BA3YPikrYGAj1cBRKX4SrGMikvPo77E8QCI8fWQx+/A6H
9jjntmF5tqVRdO17wz7kMGK38sMuiooNsvBiFinRfB3aR9irYmIVDKVNhPyFdvqU
kpj0ckYaUMKjvu6xaHc7Uud67lvZjLhYh1nyLwCqOvOXBMOSxQg6sHiJwNpODqs4
46m4zCbhi6eQm6+VEAMUh4QkZg4fllY5QazZ3ImKm5s=
`protect END_PROTECTED
