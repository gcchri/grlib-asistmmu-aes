`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8mNA/hL28bW8rTrEaW6241GriyjYjMyJX0h9+KFUfm+ITyADCs4CiNKGihHY4H0C
XDRyBcsWBFNzl6bznvr0dOaXsIH+aP4ofdcEv2uEfceIS0Ldf9K/GGcwi6f5c62Q
nYi8oiKrB80Ly69wmsljF5AKbwxfWsyY0dsmPKhGNtb+cQtFqEEYIoCTJQ6wQpci
ChfuBWvqLOwRGRoeuXnRpHIWFlCjbpcxE9/9gjn2VudM66F/UIPeO3XnddLAY96/
kBykNdnJ0cYQmyytzeo+tuFBQZBrDX+8V1ksdF9YBTKnZWYxFMXpxjd5AvbJP/0q
`protect END_PROTECTED
