`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aacTKxtMZfcM7k0sg90yBZQhEMQOHxQMEx5Uc1txdW7kOoGv22BExd3vDeAZj0jN
MsoqEpWznRSfiqbD1SmqmOzTYxeltEej7IT0u9gyJwsVclRBBixT+78bqpz1nomU
3PkeqOPixKAbwQ06OJTlGJJhVMk1nC6IdZgBT9F2PL0vwnJ0PS+n6bGVet9hWC0C
NIhqk0vAnSqORe5mfk8hJbtNIdD9KREfQ3pYJllLUi7vBb8kHXIwms613wx7rLiU
WirwnY0+fLTUNO9Y3vYSpA1jHnM5/671Q+4ABOLZ86PY/CJjvOXnKdqTI4jG9Agk
OFbWXx86/EsN0tPDIdMLSX493/Eu2T7PDwFVPTdd/5Qe1g65FVjfuxZoOn90N9ld
Jn7N0gm7FA8wA+NiLjjk1v5CkYm8DlVe3xA5ycOPH833Jvh3q4RhBG5l73zim+me
j9IoJ0qlKjugj9mVQB6jgYQ0aYaZ2NjU8leSUe5VUVZLC3sOeFgIeIsJpZNfOjU9
BaVuBZwhZxGDI8qhq2enLKtU/bOWF4upDKymAEHCkRUpEwP87W0k/wSZwIP2ng2c
GmBc/Jr0yZzz7FQgu8BgSoliwUduORVCq6W2dzB7eq3vibohwf4a9V/tvScEkYbz
G8KcSRLWvX3u7Mtb3GPGbOgx5DE36i1RtbyVtpyZWZHdvpvkVglwj49LEOKyAIA5
SZN9tOkNQJzBGi5Wkewz0rbqc8iInjBAESdBsn/Y1qcAIaRnFAUMWCufa/TREvwS
7pwgqgtTwohEwFEMOxfUflCutUh2I5AbHodHTATY6oJgPQtHvTmW3s6wkLo9mlU/
KxrCLF1PoRt0zecKMT9Dv9Xra8yYoJ43/Xk4b6tIcHlNxaY2ogEnr87bqS8pUIU1
8FV5GC79s/KlwmBiDDUbb01rBwKxwoAeb8qSjEshV/lyb0DZXiqzgdC5VlQwICRP
sUuaDAnvnXcbeqNe9BEfN1ryoK2+TZizDjgRzGG74hHtg/S/q0/IQMaBUOl6TZLN
v3Vi5fXUeP4ms/+j7+tn84VNx3FKxZHVS4UnT1Lrn/AbhSvn1reVOYJMyJLrR1P+
Bv5WbxFeDvVUbJbu6AscKH5EqDaksscsMpMmCM8J8DTL5qLaMgWKaXT+pgSXZtvS
lTOvxBfndgIfWVJRqBjBkrMFDr8mnk+EcnE1uuwpDP2rIj5qOIrjJ6xU7FOXsDt3
FpYde9FBGH5tKE/I0NJXUWwcbjUhtDFnp8k13uuivcqAL/wcq3W0zHZh0pap4ptq
`protect END_PROTECTED
