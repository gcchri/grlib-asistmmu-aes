`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PLOjtYxg6YEJD6efOBX22WQFa38y6/sebgbpgBrTPwGLll4ytxWjyV4EhDhTkz5w
EYb7DpzoDGF7A6N6m7waBopKm9nCJ3vO6EXzgIrI42WFJUJwPlb6ng0waMx+njuo
0WJUfi29/KilaDpvdEiXxMHNqvNqPls8UGflKoOy1qlSSQjvNSvMi1g9PUEdem3I
a0ZHlc/9mTXkzSGZVWOz59Xq7lf9UDnkd/RC8kCNTtk6rxHsYgCSImaX2BhI4sSu
LtcMpMs1/K8q6XMSDStLFcN3DsKpA43+cJgsyUWOJm0731epgbeK/Ao1ddkv6k3V
xF9yL13TzFO4OO6F/4aq2YvFJdSoQUPraU6Yi0rSbxUQrjjL1F/X7s50CS2PPJTs
nhnSGQaMgi56lsu/dGaDym1Wc5Zzv4K7BwwdlXy0o6rPLoKDx0c4N0pC0Z7mMAkJ
QXqMSrqpXY09U6l7YEWaiD86pKeA2eMNhx4iDGi9FbSDHdY/B2AbtdSXvM3hV6A+
`protect END_PROTECTED
