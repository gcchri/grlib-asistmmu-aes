`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RfCmqn+EXYx7JxEPOfohhkdPPaYl16txeCfTPL7pZWSR6LBeyB6HCreVA0Ge4yWh
UeQzixbHoO/uhs60z2GoIiHuzVJXn4OwWH5/C2EaX0euEZdZkA+7ysC0sdeQxp0j
t4PvgRjYpqPQLTHOHACoGOr/eHgjrYKmUZUmtpZZ93k7Rhg/84GTEXgoRTBu8E6M
xYXIMCDkXWs8fLbgDDcK7tmZjq2hnBRQ6nMuxixcaP7yPITnD93yr3Luow+pNSp4
0ZUesy1oPGh40cNBfCo8gyLk4hfd2SCQF95yPR0JS0O/V0bM/A4SCzPWBID0lkTP
ADH6zAXrlTtDgszv49TJ2h+hdd65Y3OP0XYlP9UHmeU3NjCNc5qouXf1fhjg00GT
SbaAJjNqKfVoDB5ehNHjiB7IXJHMP+Z0BIpMc1r/8ve4wumHpO3i7TgPuChxMVEn
`protect END_PROTECTED
