`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LX84TptDe1f7uLk9rJlCAxQTaAbArH6Gpnk/cDaHtJ3WK0af0Y7WWvjLQBsAoMFN
8mPAv896BcDpb7GgWRW48Gme8DjdgsuyNjzkUw+RZ70DqQSjfPyfYmvMbLkwuWgL
jwmbi3H9E1S7Tq8SddAtBIp2Mf53d/DBZOGkk+K56H+j9kEvtHvFtd0bmYuMCnU2
dzrt7zdgTScWatXsD2nZ0Pvk7SPBvfC+/jg24hlTVrewvMZ6PZdisdtsaT/Zw204
k0XUVUbR8P3iRbBh0cC1ko85vRk3DfrUEc+zf9Vqal+ZlQnZ21wNy8bDZ1wx+pDN
5raM6Vdutu8o8zSp+qHbB8LEnLiy7n3AvfJsLopo8ygQvbtPFVD6d9R77mh5zvTl
r9xL4AX3t8k0oiyDgk39K66jtDyaMnNbP8fSvgUnHe8vBVwqEpzwno2KLAoOseY4
`protect END_PROTECTED
