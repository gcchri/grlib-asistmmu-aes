`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nLXsQm9ZeI6nios0GrkU8JmBh/+f3KpZSPHOtfW5h0KySH7i3Vxe42omR5Dmt3PW
RwJ5L3DE0EUh2e4UCPJc0x7bugrFMhyVuy2XXQryPBr5Twiv1fym72LpXUAYqAgM
i6m2rampHhuDz8OKDfQiS6G/17gbZ3LpFq11QnDvTYFtFDnRqtFjhR1AZ2DH9Nnu
sHvihqDj3o6gzRGoNmA2nZkh285IQF4YOas+JoSfGQEPRl2PFYIJk2FEJyYmBUpR
ngs7KqGXOuCeOAtXXH8fA4D/VhuH6Z+63RQfxupivShkRp5rrL+S1yWI5h1JlN1V
t/9Po6as2Dc0Z2xbnbHUj0NvDvgI1ZVO+jUWcjGe7v8m2TTqbZW8WZRzfBIOfGTG
PW8NuuMlfM4VCIhvwt2W7IZn5ryjNrAAxKV9aJR8+Llud/zofQU5StjQlWVe2wL6
B9UzW+Rr21Om2r09UwTGGyxHsGs/JRB+SYoRNApJ+3/kONtuZUhFM8BvlUGAMhvk
`protect END_PROTECTED
