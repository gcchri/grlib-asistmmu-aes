`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FW2mERziiSPUS/toZmDENY1uulXQg78dz2xy+uTPN+TJDtTN6LXxaMnEwy2IbVVA
IDnw3LUgwDd3efXHqKayNI5BLiUtUrPE3Jr38Mj+JOpjHa+QueyA2vjD2QN2dQhh
OqbjXE+EUziW+YVhdMjrgTDWhaTwjoa5PJVtpyKyAJmGQmYwHIL6UWz8RifFt0go
gOby6h95TmTgtmrt4WcY3vfnp6DxSYBZDBhrLI5SJywoKGgwiqbZR1Ck8EP0Ny+T
uOm18DpiswfdcXBwoL0/Wrvk4Sn43ZDAcsfte+5ybTwvb7SYB/AcRZQQdcACe21Q
snR7vl05xs9kzchhJe/AVw==
`protect END_PROTECTED
