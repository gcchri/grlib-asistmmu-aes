`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cTt67D8F2P+EqLcTVBvchuTFsVV7WJxfgSJhsD2ugP106qzWX0bSW0349p4/f3UM
tj5Cygd0Gv3msEiJye8X5NphoZMArTa5a5+TGgu6gyQ2oolft8wJZB17upbbz7Zb
OdB8cH0JT9WXRoIttOzeQv5MnZ42OXQP9+kMpVnUSjITe9249tiGqUoXgBxVbzaH
9ULxjOyKidwhsqbQrnMaROgVFy8vpM6SZmULoN9aAhUWdLvsEKFO0hkV0LEubTnD
7SEtpaDKRr0n+2QsdTuT6iMN3on1JsFDtqhWkzhZ60YMXGFMQ3lKKI5+k7nSwQGN
IhX+Yu5GMNeLsMKyVAwc6oUGXISUu86svtgGu6kwR3a3uXL7k9eR0EQttZxel/7Y
`protect END_PROTECTED
