`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZDbb+1y7i47cZYnxm6i7/x7OcaKzmHM2yMFTxlZLsm0McKcHGyLyl/T4/jquLYFZ
A/nqBd8+RBKTu21TPlVr+wJby0kgFe8JCHO6kOffZIP3n+i7TwfLRYCEpU+LD6l0
ydwdXrq7Ou0xsRETiokqL9G4m9132nS7unPIapq/TEWqslXCdF2NDbnAuQY+ilLG
Qybc8mwG1fjMIGR1RnDaN8MEheV9ILg5F/U8fn+oFF9dJQ1l6HgxhxoigCUhawEO
pJwLHDz1C0IjP1acGTUE6im5T1GL1Oflw+T48fRzMGHq1r8YneDOSfi3EDLBjlW+
AO2qBKxOcXq3xeszx/pkK0Yb7JyccIncHkYsnNVIui+5PCwMEWH8WUKStXkJf2lQ
HklO4sLgPh3IjSxESINHBgiL2TFOnsdTbNCkOwgO9F3PjVfSmn6LNL6PyoGvh2GW
S+axsWTwQJMFR5ZJzUAHmg==
`protect END_PROTECTED
