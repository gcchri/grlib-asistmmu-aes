`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bRs6RIJbVXECdgwKPmxiZJbT5kRVRPx5qVh8pdNdg1Hhv30qpymFjRSgpaVWU41Y
z8fadiXhZqZq88H7egTPfy6+wM+s2nrgoPo8NICZNGAg+OGlXczphnymalsPs/2I
Xe9ZpESBZzwLE+uyt3rJWeoB9GLY+m8UNj+RmbifiWk+WT42v2NT4awERhDqQhE5
srV7YkALzAEAACexKw7oY/oFU9YVxv6FEaE0IjP6o9IDsi/mVGgWIKAtbP3DlJCo
fmlOB7E6Q5sdL4FsAnDe2g7BW2IZgYaixWTyDIKTHVogrGCpw/RKatYopRhg6B7q
YRVhxXXwuT2v/RkwzQolToUTtAYdxt6ed5ZqXmQT6HC1eXfXlGZcgqorX7v57SR+
Hpa+TbaEjDVkXN5CTcJjcFH33u0I8EEm5uZ9Mlb2O3gMZt6Ip7BTydAqOdDS3RIH
+c+/MXbMzPoUinxJZ/g8dJkrkuhCD1UNiwdruYTE8zsnk8MZIaBpZx5lCdXisaNa
7J0dsMQQnj5cShMhkqO1cuZwQEHalWtivXaAjkecEfj2vkb2PpoTZg6F5MMUyFkm
aG2bHhDbUcO4vBrOQXlRg+Z8H43OKlahAnxo1Oii042G8CD5WEF7geB+VVB/73JK
SrK747PsqoOs/GPm1j6D2PUcGE76kVE7f9DJq173hQhJFsyzL8RdYFgLwFV8oTby
tHV65e+kwWVCKchsCRuX/zMAZ0vtNHtQg+u7CTRw8f3a/HJAFrl5+OPYOBBQ9dxx
w0Ua7/0HoMJlxMRM/0YcGS7OBoXimB1lMB9c9MDr4x59srp6OMUmvi0BBnfnGAvU
8Ew62uTZYfAZe3r0xkyROkKM7RVgqU/SrNovrut9ysfMmDo0cfgc6KT8O3UQlIf7
hzvy7plltMbwpOteYZaWTjkj/82RqudHDCHAyB1z6k3OHrxrmcr/IfeXeGsTeUhG
zfFpGARYOTun7Knwi7KI3rX11uejnQozGQP3JDvlOHmwWoDUt/L27usHqBFx+k2+
MyvKoKl6XA8MoxOTOs4rE8xWB0lHjsZuU+IxU8TtlJ+Vuk/zDGx18ee3kppLGzKy
GRoaLOUcr2JKTYHy94poW8oUJqJYufH+TTVOQCUQauuuxe2xKwWaKI6nK2iGQCxV
ul41XrYV7/jEeLvLBN5Hhw==
`protect END_PROTECTED
