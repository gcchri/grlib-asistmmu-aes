`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A67WQT54pwAlQoE2wqXG+nIyL3ChcSlhuGvxq48+slzIPn8jyupI8jz7Vm3AoaRl
v8v8L7jCMj/fcR1DBog1fvKp1j1xX2CgQtMMaLihrcTt0Ucu09Nlff5vc75igb9d
Emjetj8U7OjTBuFg44EUnqOfCWYUDK4OQw+MF19UHllUCr/uxcxpvDAXHm6D72Ei
UZ0f/HjKp9nUBgAe9bOlcs0YOdNPD4OvmNToioSJclhlo6WLKLJZApcK4EttQ+T/
fMQzJ+QV2EqxnTVkVUpWXItDPM2wSV6tcmMzhETuOxbHQpvnHhFOMsxycTPQGCQQ
gdECmUYlVRSEPdisElyR3g==
`protect END_PROTECTED
