`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KtrFMW9rExgWWk/ZeA0rj8a9pDMvaF1NLQKQ33CPfcD16ytaJrH9fMBW+74TmlxL
G5Gj8LG2ZMfo0hMsSSnJQt7jAo80zWwpPqc/iOTeAroGYyxrSGR0dqyY+xQuF7uv
iALW0YBklwND7isg1PRIzb8i1b/JQPdcGpENEJAEfFZnq05Cmqj7rX5kzL65qlpN
AblEI6pDY34wK2GnVKWjF0jXH55si3eaHQsu2Eg0SCHkc4yer/qMHxO7753upeiC
3a/bHPnKf6vGDBtNYtaw+oEIWmkuss4RxiLJzRSMvy5CLlVbsmV6TXs5xGlvdq5G
AcS5qN2xy15lX7FgdiFLZGNp4o2RdBNF8+oFZzQQZiEU6C7Z+pPoo5ljX+xTZ6UN
T/PVVlCgLLtnyKZu24M0W764rFuOGn0uwZIj7DFaCj0=
`protect END_PROTECTED
