`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tYO+gVXzRyFTfIPpaE6BUIIcH0HMMXXBMDa1c1DJrAb3psOfUhUvslAiQ05XXWxR
1j8dPvd4lNbnNxJvnlQbqgEh/L2qP3GJo4sW33vIsRqIRhExBrZJ399TlOs2WX7W
C9YRyLgz3JiD9cagIxZax/1joj4tIWBbKNC71P28aQGpfM81oov+oC6fh5LEkGeP
f0r3vMgyyOga/Te8shEDxBDZagcBVixnpnOsdtleeR0vwGbOXhuxOw0xUK9k4ZH5
PZRJDeQEpoH9LDCz2bsdb7ZVUYYA4vr26aW+bihxvbTxrHx3arHmfp4cRV4kFzlw
Xqau5UIujq+2W/KU0KM5JFfCxXa7Nn9UdxCHHX0cBiXHCPbtDE2EJWk+iEAgMyI5
B4Dbk1pyQtEv3wck1EoyPA==
`protect END_PROTECTED
