`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tgfqyyZJdEl2U+PuowB+qqVo1KOq2VNSDGpPyYDFVrRxlJXE/laRoyDqE/cWLhQB
C185Ryez/0TxzMvtNxajk9MSMFSB79U9bhE5C7LWpzF8dYvP1f0i3BDM5M2VCigE
zFgpDinUa33VndPkObgNbqiM8YniUaGAKeCgc2UsHWYz4y1DOhw+66t1MOJGLmc5
4iMeHspd1hdO0R8ez/NpEyanUJA4+7eZs5PFeG6JRXnB9yMNu4sOBj3RT9ACM0tg
vSX7EUxgRbL5Keo5aNHJ8wUQbG8JkSsiA2mjJXRSMpQ0PnKj99xDwuAg8CugIWDY
ZXv6fr7qlHvizhW0bqnnT3+orR8q7sNsh7DkVMYIFB6N61bJJ7xQfkMPmz1yceBy
xWtlCSVN+BFehi933dHqbaKENU8kYqGlzeNjFHFazo9sR2G3LsLqadC/Az4DD//d
6WMyPLDQuyMBWrfX4hfPR6EHpLMI1rybva8xyk9FNGWLcDVqQOmeoVKH7DIMqF7o
5aX4xBUqeU4Chcf/tTfOXWTzDq6YB//RvjSYL4BkcEPmGIRk+iiS+DhZpnPdyPNu
7uRB4X1HokuVjQbCbk7+nMKYbiJFFgeEpWkC0TIdLIY=
`protect END_PROTECTED
