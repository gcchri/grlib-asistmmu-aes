`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pX34rpsJnHMuKC/GzvdEcdS+KkN4LP30D1wumd4BZrPXyIpy2rQbY1ZPSU7qb+o
LYb1YTw6qvLnGXB+BoEIrQ/xKr4sECqlhx6GfiRV4AuuxTbCLOEjrRdmeVhNw1DA
eMKCyFeDhJS9/+EyF6jwpoDbx9iWOn8M40CoZaK4CloI7sJkeR/Jy1wdN4bLoqAd
45yIXqTfLQIJzzKMbYzF+fJgyLvfauPW7CfmeGPtlyA9JJDLbGs2wkiov9uC1jC5
O8qZQ7ItTfn0cNLAasTRLP2xVgKnMPIh8f/eSE/iF8PsF8Z/scvjviDM80gJc/An
F/sgy25wD4TdjcRZt6Lxvw==
`protect END_PROTECTED
