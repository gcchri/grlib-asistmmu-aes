`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLXeQUIbDgx/OR6Dqvvfu6+6H40KHsVNAojQjjkyqQ+5seY4p6W7Q348J42PCUhT
jRlk74QxCbihCTqHPZxG3OXKjJ8oNM6lq/GfB+jlCSixjEH+dsI5CSm/jqwXnnkh
8iPEmIX+XuBnn5J1MR/xks2lPpZpLtOfUhsdqAid+0uFZbuy4KdGF10bke0Kr7JL
OENpqPiM3QlBsjwimpDR+g==
`protect END_PROTECTED
