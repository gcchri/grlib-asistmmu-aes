`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Hnb3W8Okv9l0SY/sUChSOrYF47NzmfjyWpTloHFrpKqflxVV/z2L43LSVLWlaKM
aIGqtRkdEEAIv3h5j3yV8i5IkGGY6nQCIQhr053VH7MlF5rrK5A0coJfcwn+AotP
SoVE8IR54dEe+1I7bJgqZiNNYeme/+MSfPU6KuSB+BPu83HI0hId5KZy/3QnjHy9
1t1YgKMK43HZhMUMZbJub79p1e0I1rmnGe/dCxA596G2paEdOA+Jo0LXmooRGuFj
tAJ94i/ZBD+ZrsuaImt2bw==
`protect END_PROTECTED
