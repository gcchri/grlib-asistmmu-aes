`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UDKy7N5bV/It+52Dk9i/QRU4xhTwOQSZsNzZjYnZzm9B9mVf1mMDqJ9gO32GlZ4o
1KfTM3l0S8Ycd9D+NkjffwXpAWagNCPu73kcC3jcj8llOsM3QZCfBoNX9EGXKpHv
vt6ACoQxTotD/eueGzyok2MTUgPX6CurS1UyHmIglH4fZrCu8v8/wIqjgIYG+HQe
21exPRRnaYvlWOiHcDQS77TSw+U1vzeAHyxzhtsr3TNY/mM1HWnLB8tEF0qvTgRx
su2CwzN+sLdu9LgiYQ4PU0xfuy8pFnRY79o0m8akwyvDF6xagIOJQEyaK2IYbF4N
wRno8F2lPkJq/4m9keT4rHBjkAt/3Vl3//jWpQwTYGx/Pzpx95sq1ZLBXf1xFu95
6kCt6+X0/DicCR1D1KRxPekYzUH6xRrrm1jnghLMivQKs6LxMHocM6abqVWySzI9
DQHtWX9ZkpDprR2lgJ62t1eDoy38WrqyK7i1/hYnMnYLHMYW4vOfNNPYEApk7Pj6
jOh0MSMDlem7foCKAXY01VfpLUsbW5EZaOOiTH9KqCoOtEck1WNRzAHnV93si34K
XGQFZeTRgpvSs4mOMklUeCiB8NRPhRzOvg68u4SEOXtxjGKslkg8msCRYl718ikQ
K0HZGoSN2d5DDQdXYOEeqZpvs86Cn6mAJiDgwJJk2CJGFAeWqNNz8vk0qTF41tC/
M51cXho/BZenWgzTjmEQvE7hJyhpu02UV1ZqaWZoH+92tuDf10VcaWj6tWEoCgX0
XrWWInTjPufFg9KWiii0eQ==
`protect END_PROTECTED
