`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXizebQ6RFuhn1z4/0VWkjWdPDtJ2xccKN0IXve+2NvJgTlwAz2alxa4RYkIOTLE
sZlXs04kwa/ko4yybciVIQdTjbgnJ7bSygql7Q8GplInSrrvDz2MmzL6BWePc9rT
tBBRauD2BSA8QC2otkFB5Sw13u36rC9uO5VGZcNMNxbfaowy9JG7dw67PGXLXBCj
9NHQNQvAouB1yvgySpjhcIzcFkfKDyS204cIoeIZc5EvcQ6+YetCY7pLwG2D6HcC
Wg1Vb2t65KF1yJ0OkUBk50YXhmYBwLcc33b3sCNhErc=
`protect END_PROTECTED
