`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9nKELp89VwDbrFaZrN5gwJJBG59WsE4HG7LKEFHmsPzdUuaHwr/ovXGtzioGyqOd
G+OHxRzPp5Dznq6/qzaRKAX4SG59Sy03frJj34rnKf6Wi5m9AFf0GtzKhYjWob4l
uNVy0PRmZsYLQPU5F6eQuIiOoQ4wKdHXOdRExyeGPnJdHZ1efUEhNmiYWjWUg3rQ
1jvcwVaZFpUby0BbrmZDVoOjJlby5n9Q+qNQG5y/B1qB1xw9QzTZlfZjwUNhY1BB
lCqCLPEom80wm/y5aYa5JSVL4DcdVZlZW1Tg4ROSAOrzJEezbDM1kMEk4FfQg4K1
zZtwyABOYNgMDCDGayuJNtnhfd2pAStvKKSbcMYHWvMbSciGVIBXXEPbAlk8uJ0G
8SuwuOAQ0zJUedYvJMRwnxmpnwePaRXsJ/LRR1Ri/aqyL2PctQiuUaEWourV7m8i
`protect END_PROTECTED
