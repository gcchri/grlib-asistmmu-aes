`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1AwHd2N9VB2SZi85TiuQH3lgyVmZmJ9mrMMs73fL28ncphI4Mxdrld8tM6Wx7W2J
cqD6Eha4P124rf1erL5iXcWeAnxA8AoddHoUs0w0LyXvD2ouJUxj0VoWbXQn72Fi
2EGVqsB8aG5DZGXYzU5Qb8Bb/ARFjD0Cq1/fHnUxsw7HHcbuKHlvY7ijLZBswCJ7
HTrAypnOA21Ip43hpDs92VE6xw1Ly8TdMRrqWaH+paENE09t2ruhg3/Ivs8qcbfk
XNMeR3MPFKolh8xrO7naz9Y9CqYK4y3mhSc+h1Na/BOJgMfw+jd0R3qHdC4VHY4R
Ck9/cKcXmaglLbEyosgwcPalrGGc81mCesMnuahErRkKCoXxGOx/ZsW5otXuVB0i
zw6/9ictvQGbuTnAJbt/f5lPos8hXKhJ9QgkbdUEOvo=
`protect END_PROTECTED
