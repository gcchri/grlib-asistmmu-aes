`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2SHr8S7oaM5q8i7WES+tPljo70d770m+DclvoQhyAebpPsHaDKaDOUAYA7a4JEQ
wD4qTpbAtr3hSgXa7aPZ2AViCXpEa/g95GZfcsUUAUQ/f0L3m20QiK/c8wcvl5Vc
Z0wNG0x1j5N4Hk7MnGIUApOYJupJjvVsKvTX5USiXpS/xoxC98T8GAc6VO2c0OTL
EErKw7hP5aWaQmQc0TyJziY1C1FUPQ31v2m6nGeo744VdHSWRb+JRvlBWS8RWPCP
`protect END_PROTECTED
