`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1QwRpDLUUiTIBvYOJKHbQb16b16M3KcVovwo0gmTWcaj/h7VADMmBi2QnBiAK7Ru
0eGSppiHf/hIP6Fss7KnOBXTyBY+dJUubTzy9TUQ7J0PZnFKBdvFtPxiJn4ltd+M
w+sGipGVeAI0hCfFzLDi+SMzT9wyZh4Lv7lpX+sWmvL9/EkNW5rhusZEsIPb5XIH
4EtsfyNWLZi8Pu4hid27qeFXNe+tmmMUp6TyAh70CI3StKN46F9J1hltOyWSl8wl
zRUl/s08hjdQS0XMV5Wfyd1qKOJHXielcy6XfYB8sv2yyzdIP2dvloaxzrppR8GG
UjBcDbFdVZmPaH2hZpZPYg==
`protect END_PROTECTED
