`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Q/3fFqNgNjbIfiUMbTg6gkq6IC6Dch2mv/gDBxn2YimngEzwPEe+gXxRtNBTx4Z
xetxKZcz1x22BHstQ+6GUKyeBMdswWPnJprKV0XVGGuXgMkStdE3JEpQf+UKrb9W
CNYfb0wI6kcp9mL3YgMumQgCBkwIGPjPDdWSlYLAsBgpTHb2WrSqoIGYr1cZyY8j
qu4WLpqUaFuDoefd49dMezJfhoPkpuKoJae7aUW1mhlJyCbqbEbpMV4v32w/u+9S
10EyLwkNlxFhFp/TW6W8BJgiJT9/JVHnBNudCZlHJF04h9vj0qQm97AnAZtZ5BGL
LaCMOHwK3QMdORhiADh67I2+024JJsYxccbgHKSrFEdLSmLQCsMf6GfpR7MUSfhn
NXOT8iUKkCRHfGrHCTUl0ZmmSWvK9FjDFP56IZPmq/9rte3xgNCchiSpTBriX+1Q
F5F/m9ktPge8djrdYWRoPn8VyIGiDhffOPxsY/TwodDHgb338bawcStzulQOOYof
iJmZDZiKTX0hC2A8vWTMppr8ZalM2G5cxEfg/p25ZphRV1JLmEzUZMk/icZw9NyR
`protect END_PROTECTED
