`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EMwz8jQuN+x6GmfsYyS2W8Oyck/r7odhd4fKUJErySZTqezUMgAjex1iERk6D7M
ueuMkUc61ghbx6i0W86iD1wyzabF3YujFEmnR2hC6vjvdaxh0PeDxJwloCyn4piA
O3JXF7OnuNbZFq2oUDieUT7QDBZIZnf7sQIoxIxvqYS6yjACO/pnGOJ4ShfJieYV
ZxFOtzFy6LWhL4qsP95AISG2/hJEjt1qBVqIoFGBZ2D6xFZJ3a62OAKEPuAyGBYd
d9RPQvUbs7y2TgsaKi266Nb7HSlLLG0iqsN7K5lG91lIrgqQznliqp/Bbj9GN8PC
qhYRFgAoofKO3oBDhNMN7uwngocCnDITUnfJdGVoqgKkcB6gveh23wCtndKstw3Z
C8dliYups/HTzbidyPrCWLCisbJdnDD2EWPZ+bRJFvYp3gFMQqGN/F8JA11UA7j1
seVo56fKstLUsLuOmH2YOtrCYJAENKy/DbUNKDOAwVErn+czmgYZPskn1a8Jrnub
WyBDkHaV4CEGRLUZGR1GObfmsBw0fhfVfOJuU7yQZf2M7gopKQsQAcF1I/Selch9
BJa+WhtqTncNoagCkKFyr/wD394i+ctRO41BeNsvZpYQmg+PLdNeztf/SdVygUun
D2KMfVSxJaTgepc2Cx5K1OC4PQPE2VwW8O/HZ+V0+P2pdP6A0ifoyCVjFKJv+Frl
NrkYFI+wj3iXTCLKWRqTu6n8aGZbD3cX8u+R/T7Svwy+pkodGVyE2TqZ+Qmbwlk4
fKAUCPezhQdAT627Bj6vUFBFu0YXUhL0Gw5UicL5Sk0wYg3XPw7Vh1+zJa2ubNx6
jbR+nH1onrYwss37GcexD1VkvY+BsCfRiw/ZxZA40bVsYN6SKWEhoxVzyMI+rbkD
KRC3MRJuObKOXcaPVpQAYX7qRZ06tj7xVw1CU+kd2d7xzpIKr2aGb0DmwMjjeeg8
am7gUrAxW/qW+AXudqYs2P3axtFLN46ecXaKzC1p0PEyAGtUgvKolB/JTV0F/sRm
crqXSZvYwtRqDXV8cNOZEEHtPqrZWnODrlHqoZP7/vllNZ/w6K39QOWMRvqIBrHt
/ZtfOlGSlp8LeFcjyOrMp6PtclR2WjAaH9M4nqQ4UtV2HTw5+fyoaXlVKlU1zK1Q
3LYGD41nLA8i9AhIh91NpTUxkH5biv7AaJ/5at/ROpWKhmEaau2bUXstH2fj6Kkw
Ryzwsd2dKEBw2ilVwEUEMm7uANON+zXTLt4R+V4437hNtK1TaV+gwwvTtyOBT1ZH
CFgIY8XquPtZwx7TsbNfaZSBlxuiKwc3aquUB0Bz/XeV9OP3WYWaiclNOI15PEOZ
8D6EPXJwncN373hc97Cm22j4x3ltSiwaid/jhZZwGV44oA21QvWPrQyI/H7/or9m
M7/x66EO94RI/R5MMu+Q/D3yaDjC5z0zAGvPo2GLa+kQ8JDfvHhUo85fHOzk0qN6
UctzSi3HAdDPAmM0a+JYuyLss7wrhXEtK459fBimaZ8XsujXiXUtVp3Go+UCiAVp
Z1crmNmB2bndJJdwSHvhNvLoqFAisa71FGyNyws90sZatPm2/yRgVab5/X6OL8w8
XYSlfHLujJh0a0VQOCjjR48VF6iwfaRayEUh7dTf10W+olU+qPnAqS2TNXsM5Moe
F6y5Rz29Jl6I1ydZj1fMJHyomUQLOMXwCKoyqDTlwjYxuL7FSlbpq0T9FItuhhGK
vB5glzeGz6g/udEDOako39MBjnLitTvE+edrGS/6GtR6h4XCPATSd5KJPpkEc4AP
MCz7OJjlDQ0sMizgUyBkdmlSRQ4wyhwes7Gor8l8UlyEjxltSXykBg3kCr7IIeEl
5CZb1ZOpPD3+gjxOZPvULgOzqmYX3LxPPG5Tm6LaGyT9veCWwGLKZgHOdxgoSX3L
pbvSi3l46k/7VBs3nQ3PC8ZaAAy80OStp2ngFeFyc2MrCqBAXAi2PZEuVy9OCKpY
Ypx0RLF3CLFYMm6sPVZHiPojxuMjShm9AQ9X0rydmqDp4P59Q2ft8gFQXeeEu8Ei
WZg9yv5DJje8v1H2OKP/gxribJmz/NKQVen26PE8/NgIiT6OkZh/PpcXkjAebc8G
EBz4bTfy2UBIyp0i4zajB+6djhKHPPRbVdZ0nSFTJsQ3wLJ+RTkRjR3r9AawNq74
W3hjCP6ZNSh/aJEhXjZRQPKcRhLU+8Oiol0+5Ad3huqbtZpvJGHOdMOyCTmEOhpu
V1GryC8+MsuqfbII0HEPsus8pRJqEL/UnXtzm+ndWEfRePUz5crVD++gZJIsbgcJ
1tzQxYCbcHFlnz6pkMdAh3ayCHPLrVTIRq7JowpzfNTzHkaRPd+lhVsEko6sHn+s
U9dBaP8+3NXPxdBEhQy1MUiQ1Xo5NZA6VcqDw59DNQSDFH49cw1x7WtG3tQN3KOI
Qywcc+SVs+kNetiSL2YCwRYOFJE6ELHewFKayWY+iCy9RscETVG7KvbKKtO72YnP
gP13sG4X6K/qzreMLBbJBLCVEAZtWtWEmme7CMsnysjGsCqu3Qc/PNHlSFeJrGhY
TCz/wOX9jPBZB+rnV4OawxFNgTQmG6504xiEMXvLmSAURoyBRNkTtDvdCqEdTAr6
Qk0SDay7c/ylV0IBvswB/cEeuUhf+bZECs/wWzi5gE+xe9shnWMOmqTKt5ftflOr
CcEADndzkiZng7dM7dWRC8TuwsztXXYq7KeEyNv6Eb4rxnpUwI14AV13hT832KBW
0lowmmBulTqW7hQNWDSaoct0N265FtUwzJUhFRiVIRF6ChGj6f9g7O37W/E7YK1H
J0NcqYRNvJECoe+iyTzIAiIHNal3APzMpBWU8b8gTN+Nt6UlCcMXFJCpdqWLkHQO
vSMZ8WC02sWEEui7kyLfbOTA1owWaqGuvatKIK65QX2swp69nffb8r/EqeNHCjAl
4vS16lFcv7TZbvcZGB1ntNSVv8D/Movrc+d1alMuddP4bs3uAnxAltCavV/Xx33Q
bT3zfKCBZEFPCPerL1NwzLZw0ZKdQmBCBl/RuxEmMmoMTbFMCeMwwaqgJBSmPHSh
rpMjNiIqbdw2qeVxr+xSciAXIx8g/fz+zEOpncKi1hEUj5e94h/orPdaxAnGMN2T
Wo0p6GdMVjRyxx0BD09Lv3SeOqaJ7iYY+T5elY79leKLHjWT4mcrLQP9LawOpqlb
erpQ3fC7LwRcARvh2uZv2B/aw+oyf5ERNb6UCwJN4YPxDpXHNy5XfyM4Yo69iqmE
Gr+oO44ZkHF4MHvWdWMjyW7ys4FmMcVAzrUj23JFVJzmOu59s4M1r2Bru4PeFa5w
wuvPW5YJU3rKEPAzHGLaipVs9Z4pMf27CiVvoZ3Xntb0651blY+lJRE09BvGuthm
eK3arzBwcisKQtGztgQDORVJWejFlNE15Hyn24Pv6DLiyPAX2Y+0XPd6+Kq1Qbxc
CoJq0hqlQ2eFWNlDGXeRKv8lJIcoTuRdJ8QqNf+j/LBgQxt/dX3nDxFS1KMqAVdL
uRLHT60GgmlpEpX0FfInAdwfyLbHiQEOaVjgchgLSZLDeKyIwGo+JuJoSL3DMuZl
6f+3uxeOY1Js59y0BvWG2HypeVE7u8gW6zkmJINTssUijBmLJwPyfOluQcbR+5X+
ffhGLRzU9iSFeECBU9MZKpKl8rGeBRSBxBtPusifoiZq1CUJnNcgEz5onVIuwaq8
7rkCcXl4pCinDEM/SjHJRCzlLQfT2XSSMQ/UP7ciMTRjE7cvHG7thieMpBRtEGSO
Y2w2DHZU1a9jRSDNaeqMRNqiKgsIxjwl4Lvk3S7XckDTO4roj+NHQrPtkEWmTZHy
T2wgfzklMqwveWH61nLePx9Aok6v8Pq0cKUzAMmg5qo94CsAPzgzxOBQer5vrYjU
7DxsCBT2RnXzWG9eBLYZoxGBJwc1q7hnzf6aSlk/sJLdl27MP/GbpTlLBVDu7dYs
C8VBC+xz4JHdBf7weWMqcRral7Cymb/MEfpnVhGhRzHkElq0ob2iLgwUUurIBED5
Gl5KcVNItmPEpgukRweuXY4JFNVG6OfylfTxCXyKu6nFQfq5Ur7Ani0OBTm/l1b3
++l1nUi/KWQsjIY7urL4XNxKm6kwcqcTfmoNPpKeGM12jxCulS7ktwVp2gHgDQOy
TyRU1buU7sP+y26eFiaNx7ZAJ7fBFrQ4bOcS/Ghpqid0LncoIaZ78QXHUxlWzPk4
QclIMS2V98ktiGAbtf4HECRYB5Uj8LLrh5TZJnco2Lc=
`protect END_PROTECTED
