`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gaUZtFwzw5x88ficCSSAAH5gfhTS10Q2+fqkfsXJRZ4T/qQDGOIFvg7qoClOouqs
RKUWlPGFK/Apbulj1HNHJ54NEp15icBxbbev3TXfuEzt3/jPU83kzCpLDcZsqDA3
pVnNfgVHSLGpu30yMCOsFn68n890ci+zXHwUpV7rbd+XcOK1NZFXDvBV2CcB7Lr+
vedwn1Rft+FE++ULR9rlU4BVT1y2Yv2WBy5o9I2sb372vBxEMrvRrvQucapJ0d5u
q+Q2p6VTyKyf7ZB6K3lLKWQIOlaIzq38Y5181CFTMs0RZmoI8bBTjf3IOL9iogF4
ArKyhQp5AJUF8zLaNW4dM7d4rQeLnwP76YQdIzwYAbA=
`protect END_PROTECTED
