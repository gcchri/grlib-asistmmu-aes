`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8EEFieC+PsPJr0mEqOREOzYQKMWESq0W/idZbW086IrCHH25tOoToIZJtXlocAdw
HR+5ksV9vsnsbtJyxhABuF1TVEA2K43EcZCzNp3o+ox2xSq6upQxfStkgsttnFAr
bsfDWpwpYhJhC3sqpN9e05kemvAzdy9EICNb7fBPHpPWlDggTUPyOBR+3waE+0Yj
vponeKQG6f6DSnNgn/X1hSe6PI7zCG/hr9oBBHhYQf65F/TPzi2Lm1EHxX6YYVaG
/WnbBhqCMMcfgVnzj7LAsRLlN/tI/mdOrKIp1Ay0UgdmGD+mgW6fOMcBi2zENFn5
Eb8HQ66oprZBDQfVfU96SMeVhSwiELWG31CX0fXk1w0mSX8PlRFNrHNEmQonhEFD
7jxn+u06hHMiVBvFqmJyliLxfVfBt7zGTDpcFbJD0tRMJiesokcjOOTJFv823G5B
xbA8hJESYnO3SWQQtITknCsCehTfBFvssfeEWEXI8o77i6vhuqsRYXePjk42pMmh
f/qCFxCC6zyy91Fz9Vbqr2gyTKIlk2k5h/mocWC99WU9q+Mk+jpUBXyjQbeyQr0+
7grxSCUC54IkNW4jMRB+ipPJ5tqriGD4T2knhtW4Yu0=
`protect END_PROTECTED
