`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8vskKn3eqhkv0djw07KnmeQ/LzPEAlnJMRXam3w+vxTDDBa+JTz3TB2Isd0NhOV0
jLnDErW5Ncr69XB8VGxCDtm9RqVxhyAvV3gx3nITMGOT8mkr1rS275d/ySt4T5z2
DBlKrRVT0U4u7kyK7nCvOONvUuDDyzVQu+yUcJImxAMB9gcj22i9kmZmekgMPnI5
me5GuQhqTLhzJrYoZwj8wJNqdvKHWjRtklVFpPf5yaXWthBfLVSAQGpB9ybuy3SN
5iNdh3DzHhI5CSusBJF5CLElaQ0aqxpb4sFrMx1+PtDMYSItZEFl+YTxZYE9S6kG
sZBvkZR5Y0f/ysarr1N8MimtkmBaGh8LuhQXjbNEcaPD1nY+zaREzax/UIyv8p51
Oq2FXB/O8WZ+opyvlBEXOAfWGH2tWi3indoxjLHzKxtnqNM9t/nZeLhtJmVxdXOm
CxNuDojgUslTvTY5rcetJ7xNDBS00/XiUd7Sew0fG9Cn7rR3m/o6Pm7Fvk1Aw5J3
XB7zv+ml+uZ4E2/o7qUxRHYWGwZgeqSCWGVUhaCC46uut0LRU7YR0BuxSNT+JTC8
7MayWi8DKu/ISGIEqWE5dDnefz6CaXcfHhg+aFI5lMw+ap9PZTduwjKN63xIgDUu
3rQ7MtyrVEET8Yzs1KBO0TVku3XZ+WZ9igmJ78usdAbhXk0b3JrlCgk9Eu1ESu1r
d8t/jmPXTIO7P8FxhYdvk6ham3eoHeJcDtG3TX7lO41ZpHNnl7YHtTg5rWzVAKdG
Sg4fdWYN2Uj6B/g/jNwEgARw7F0h+VjnXDfQNzgr2fd++ZOQ0aiG3/nyKcEH5Ftg
CsQu114ah9lY7ygn0G8Zg/ooiXVwPsgsUoeb9uaTAaSfveWMuSmul7spyfIv6xBK
ss+EtmZdxWTunKhsJ9jycw==
`protect END_PROTECTED
