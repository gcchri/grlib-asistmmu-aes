`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zCq6SJi7Gz0wxbz4R3SSozoqv5iKp2AnOP5ys4n+5E75VavFO4aL0AWE8IhUHBC
FgYWC2PD1Fv+o7sRuXziRlyqsmrib96HEfyN6zHtvdAHL5ZChkzs/wS9783K0xw1
qq6VEk2si9180EscZ3wPRk0/fAQ5GqPr9aAk9iTQIvAw3w2aMnF3lZd+8A4cs6HF
eAI25Y9U/gEtabGrt6PlYBz1275Skf3kek0hxjr6jKhjmWPpgh5NEVOwQMcCNwBO
Gn7mc3PHnFOkONXoeET0u96waOuXvztfH0I7M7N5DjsOFFvGpZJHohQEmIKIjwNA
xK0ywBEA8bwJSlixh2HkFU1rhD1dc33ch+MtN8AvBdhGy1ndOe8kTyd8/Kaih8zu
j2ead8c+9pIu2VkcYK7vmrajc8VsiUF4BiK+7ic2/IUMZAYAUNC8qrzStQVTRhvZ
`protect END_PROTECTED
