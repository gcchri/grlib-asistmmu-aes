`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rdI5feEQw4+o6ekTUW6riReCXOPvnz1PHh3lHUddFfMlwaKc370EJQ0brKNQeu+9
O1cjxSQ453bhrAuaCluh5xV+wf9Z8cPsuKzw+HtVhab9uw8ILuy+bBvaSc2KGyzB
5VLKfcmVnClsuD+1/mCoTcS0pylbgFIqJMi9rHBczVRsiNELj2CTNgxeRrScMUw3
xkHPSHjHcXh6UfjVCCxG/snsoOF4yGsZhDO+NbtOvHjau4dYE4OmZeyGzyijXcjN
8ZWfQNmLUJOrtTfKtxmFx8gGPwfhCfQAvddOzzIpx3fUFHt4PShSEBIYsOV6Hcty
JNSUmYojPn/kgnPrOAF2hDoKYPHWmJkKxgqmVV7xUGOQJvNJFJWyNUOyQgwLRwuS
gcVgCzBEG0l1WFttYIoalMuuUmWc6ReVJotEqhs0YL/gfMPj/Q+0rKufNiDkP88V
iR+t2MKiUsUYmBnWQvn+4KEc3r2l83Cyps2CG2NRwXLkpIJ0jlVGxBipxKU+Kcyv
jbqwJr046P2rOqAxhsF17g==
`protect END_PROTECTED
