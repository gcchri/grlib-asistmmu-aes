`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46P3gMOj5KOIdgRigJpfRjGUgyWZdsrjXz1iooEAiGZrPthhexLIjjOcaFKv2Jd0
cXg54aOUYfTvCB88EO8DixHSYtMl4Qk0Sd8y7Cm2+vPFLsMzDn2vQNGqAWcKOFLm
7vG+2XT9NswrE29yif/46Pkuaq1uLn8QQS/u8KoDaJtagqjoEhpVKoW0YYrB5coZ
80tRiI71rFyuAdakj7yJ/o8GIRBjmS2u87NsEf+9QuFixJnQhQA0VZt2dXpP0Nl4
1nZIg0Ge/EOa7JIYkcVFYIcFsZ1hmPyl+tWtUCNJ5/qCoCsgMJfkIv5xyfxnwIFj
OhBLqn1S7RLxnGDw9XYSD8rUmsYugg7eZwoTHUVu9daJy53ArVIGBGWF1vLwZ3Mt
S6FIAHV4n5uro1/5salcrVfzIEEgAZ6Uc22dMT+IN+/3p6LNI158qsMubIkng0rr
3yk31Cogj9HvR0evCQ1OOUYpFsRKv/89PB+btlvRD+t4gGOkEjlcOj4JJKId2w62
HpvVqERS0WQ3Y2wRFj1SiKfAWAJhWIJ3mKbKwl67+huAAJRfJfoKlBT9HXLlmh+e
lXECqcjf6hrlHKgDCnaSdSpH3LVJafK6Rybvt5GwqUAjoq7exXkR6Sj66wiGYNFB
YKP6JQsQ0MhSa3R9aLRLufdKzes1PbSd9ERzePalVQKxwmPdSaj39uoAHXNBbCgj
YoVqjYOX3RpQKJkVkHhsw9ElIySxxd5UUsOnAD+2b0mE9yJF1FScqajtsR1AFm6h
DciHbknxHkRG+ZRJ5aNjZLihGVo7irgyhQS4yxcnoQ1Xt43uVA2+MXkWFFwGUxcG
SyVZ6qZPA14SZ0Gy5sUGZKQFbnCBoNHIw3UjOZsEmkaqs37v/BaUSgLcWjuzX6XJ
TZHAo0ve3ebj5RQHP+CPuZrL2xobmMnix/isuURuaMla/pck4ZA9UVOTLhOF9GMO
zuiRVp60dwWBSOMQ+ioXhy73nWpx5WHra73y9vqMElg8ZVkf0dtlwJrGVv4qogvG
7G5xBcxfXDpyQ200dZx5r1OA2oyTky1Pf+hiKrUf07z19pY6xmKqOgiifqjbqDLk
JUYF76FmioteO3GM0pttVsq9m2qWUHGLltFdH2L3bj/HXO48nbr58CblUk1ZRNr2
WVxEqWjDMshLeQHFL7d//uRJrRv9vcDVtOFs9m23QF638oZCSV44ZxSyCm/x9sqJ
9MnlOcAI6lenY26Pt/T1gJUZEJUliol1ckWzEIHDWeB/jXR0QR6IwBymYtQD6z3J
Pa6zRsPvyvwvajhWp8TIXt5mPWEqGp12WKVoaW3ZWqN+v60M20xnY6SGJ5iR2q8e
KtDh2HRyYPRR2UE5OjRx3MsCGkhepsLPf76xYIiPGW+arKMwxxwTsgK+p/9KQERa
OHgBNf+uqSSsqUwrwKpUe40mkfLroi1U2ST+eb2hoHaiQHmrZ6D+BRuwX3g4TtYz
LMOtGD9fY8rjUPBQ4sIjuwsm6VTB65Zavk5nUxGDUPeyW0KYh+pqIcKm+K67hEbP
L821UL6Xgfzxtmi7xbrhmAwJm6iZgL1fGFILnS2Z5hiPz/mZT/nPla0BatW1VbLP
z4UObag+lkyLzYqmM6wsGr8SQ1g4LpNQKmyg0beGc0BYmoarSPiUOj4gb577/qcT
xxlmpmIBjaBHI/ps1xFA21YzlIucxGpPnoxe0srHB/9Hrka1TLxpibNcljWrfl2d
u5w8wsyV1eF5vjL0b1CInGva5zLPnzM2omjqZgPHT7khCwiYTEU7Sc/KvNkAjhrs
xsJwAAZsTADc/MQJvbqAeEWDOM1W/3E2EYn8IRieNiiYGJ1CGpFCs86P929JDemy
D1aitkoo3hH4UjaEsAK5iWPx4cizW4nKm1cX8Gde1dnycpU9DLdVfstyLIKoAN8L
87DHBO6XJmGHJ/mRTYce9EGkTt9DIkT4xv25Q0WbhD2HxdCJC80MeWhsddg0suC2
p65cz9D6DiD7Zc0zqn7w+2LuD9dCd9pQGdrrCIhryExVYSyV/Vx4bR/bwP7kzhqi
teWqmVOfUtazQpTqQBxuUDp5x2Uz12UVyEnRMalc3HHZiWWtcm3aHiQMrU77GNx7
U8to/v3xUM94hb/sSJKE54cRqUoy6obf+234uf8cQ/9Bg4l9vHZY85dqLxhW9SoV
9dm1EgvmNeo6vigDQa+XtTjajakrfBuJwLVh/FADkF5p6dJm9wh617x5bFZUu0VK
f0gpJCpf7wSxX5+JvphaSnaAkZeGl/YHenlR/VRzHMlqZMSomRAUwj2MsIGcwEq7
Oepo/HtpmcC3tlFAuQcFdj2+QsGaGgsXwyX/rno89/PKYAe0MkHIqMe2k5+nTtbC
VJR6zbppFdpuV0sabqI9QloS1Au4cBX5XeoaQau+y9PQB+TX7SXkbEUYiITjSNe4
a51et7utDhQrd7WCaPzknrd7p2/4jBQ5pZEe7LIUOULIm3iHSujgIbyBxHEGchgu
QmfyychflXvah/3GTuNQruuxe4xRFNR+aIEEwhgPvFKtkzAVAAMhwcnApBmw7LxJ
Ve+xmniGossH4kl3zF4GiNUuMgVXJHn5da8qvHogKXidG80GnQ6e244i5+07X1AU
tliiZl9/FEh6iikzm9J+UU52bLnXp2bHWNPjlfJ5FYX+IRBLvolJWjPxoD74BQ8l
qOb/ctoZ82XDXEpQr22K+S88fGLZkGCqTwILm3mc47G5kX7GHLGjNZyU0VEzd72C
hw4oDtOG+hFCk4IWbxfQ64MSieoXjiD4eGiIeSxmu+tCsuCvda7+umfOJsqxn5mU
gPtkMT7WY0ngS12r/nLVdDjy8+L6gfqGwWvR7GCiO77+4mTlZIxZ+b9k8zIVJz3z
+ScaF+i91VA4I43v+Ds552CF80VBZQiek0byeVc/XLmPtFkY5miFqUU5VCHJ4Q+s
`protect END_PROTECTED
