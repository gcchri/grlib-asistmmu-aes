`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Bv9Nyw1HHiAIJB2Od+ogfumBMsuTRos3dkxwvgPsAJZ2avpXAFBr5a/AuI2NRhZ
2n6avF/m6OmU7UIwMi11onNHQa5pkPQs07vIN/3F5QfypOSAaFvDLzDQ3ToKt6ud
2eeA8PAK1UP4CYNSq2vgckPiA832pftXD+U4dpCfpqQwdEozo3bQ0SBHvX2lwUkQ
0RkCHzmEB7o9kjaE2E8aZROm/5pQiU81YW1Xnv7o/qO7mX7tc1VZCg812IqG3Uy2
rh3BThSLWg5POev2be8UhK4hSqNMd8v2oYj7qqT1oYkmJ95SoataQq9xD2iLx193
sK8f0j/hyGsqaCB5m6DxRp2UvD17RzV5c8PI5LN8HEglgOQMrXnLUimbmPDOaEul
kVBseBso4CbaPs2PTXa2Ew==
`protect END_PROTECTED
