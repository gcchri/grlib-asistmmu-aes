`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LAwfLkIl89Xzfe9BCJBxP4eQEEwHIQ6MgC7PSmqBW3k8yQC56cxnbubuAXuLKN55
MPBbFBEX0uNVQlcTrSdxJY+pa7kysO5FbNBTz8k0vcT5oaagv8of065+EtIV2qkU
h04ZWoCDBCZMdiBH9mfL6Rkk9kkRaMrUvy9ByPHUF8nzcwPYCvUbDBcTVyrCd/C8
okTKHbZsazxvHtame1tqu3Pk90d0dgBi3vJT3jMp21a/axpTF6HoVdEJkNQ24ukw
A0jq/hpQFCheusO21ujd/2vFhmqzwhCI7RqH9GCdIG5OXVOo62XYRdLnSiYYqcXp
WhjoyGbUR1X0Lh1LD6iFLwhD4BtcC8RraBmBYRPOj2+55+8LzhvFtxKh2jh9c4eg
ufwnJfhZ+LU1uLnTQ/Njh2wk/uA2qk4BCGTJ0j+30yx8YRNz5j8U2I80W6rZjasf
MoicaTNqK3lHhNvgRUJ3dBglvqLsHvFcyIUvdjzDJixv6HVGMjFL1SLtxunqpKSL
YGqn6BpAoCR2AMEpTnhbUQMf75p+n+b009g4gjoW878g/7nw3wNDzumtZp4tPg/X
3FMdxadkhhpjHgvHekxYplsC/iTo3MmsMMXl1anmTm6a2HTux1y1A33w9DkwGohp
oRItRUCb0ilLbEKFFCsawAL2Y0z9CdzwKch0IydGTl3scEJe449zCXzyAhSJK5Xp
PUYUdsfbPDdblBCMEn0M/4VVEyyP2jlIeijUaWRaZjw=
`protect END_PROTECTED
