`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fGuTbHC6ZFWNWBGOUnn/nghR+pbBWIs74WfFzP76UAV8AIqsBVoUZzPILwotZg4+
WkIXYcV/aFo0oJ4uyqhy7g2Mbqo5jsFkkbPFTHSRJ71d9hWyXc4YOy+uYMUoE/9G
nXpoQ122PmIqRHJQcKd2XjJM94+uepRlYTIagZyGmXGg5VzNCGz/DhNeCmvbWxA3
HkJdOkJ/7fZmfaIonPjmhmHD1gTRog7RXpVmgbGzjHCUqFbWPyjim8hQDoYxz8er
lUtz/5MIwF8TUfbWQSpSNReRmYM4IHaymTKnhVQ9gBGMQCqRVoHIpi4f+MkhTywi
NZP3eyLtyBHEPyGG2/Ojfe3bsv6QF6YvrH0m5wwZa9ucPwKV3dRESxIDay8EF4pJ
kAnH0xPyQylKRiM9ME1gG1KJ1pmdA9DqGqId3xtxm8qiO7+XjYwwerTCeEhB/svQ
az0phDJDKzIDgk50wkhS9BvDLkXcKvs5CG7YozYKR5urI7o1qlMMsWlcQhu1p5Me
`protect END_PROTECTED
