`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LgwtTpxdGSYSu90ojZoIKogNhvdUADZSUqAz4lS29EFUPIWBVcSw4AOVX8CmY0vG
SR5TZ4G6QSSjwurhBBfNI52Diye5l93dbOEVL4I40F90NOP7R2wiaMDoQtRCLqcv
kurAJIFYrNZ7/ywDOZVT3TeLnjTALCqssJK1jclO7cwsb2BoI4+fCFNha6htpjso
FdIVDf+lDhY8pftaWxE2oObtXib2v1UBTcKog5HLXpM6ixJPrj2IvBPxpPyglC1/
UHYvb6xVE+nMm0KuMr9KyZwQdvyYe1TvSBlGme2AfQuqxMrXSwTtnOCeSAeRsJid
TzJ8kayY3C3SV1f2IXd4W0LB0m2p8YpQMdLhTMHf8McTnhyXYjVtxnlWNqEJb3rA
lQ2XrnfLWLzU/nkdK6uw1MtTXA0ilBj6DjHG8qt8G4/d9vWNuW2VV5bDaLxqvoGv
7FzzTjtqJLniHkHgHJdsDXkuKrjvLoFASlULW/DRauQ2J6LP6a/S8cGcbU9PHoP+
iJMxemLDCrDdJCY7+k2SdkiIc9KRDJ/9R3hE9+x9/1mqMVEs6PR7TtO3Dvhogn65
AhToAcHvaZlh3pmsrpCTuXckEEiGKmJB1igkVNnBWJOTC2hC1Lez4ENm+nWdl3EW
Hm8AgFraIYiIzjFTeio1UqXqulRGSF8qUjCvWIJF1i56Sh3Ybaf3lFXgx2oPrgvU
WiBCkUASdAW6tXXrSa6JIRXai2ZJ4+GvZ0C3S/TE0c6p9Iv63f4qtSapMSuRCaYY
zU6yFPbksTeFrz4QluysN6LJY4pYf4mwes8L76BNOlhdeCszlZAYZQkLCAsw8X4Q
iXr0cCDPO3fAUYT7SFmFYuCPXeYUUBIHlNnzDHzGgSPksJ59GSrVZVWSl7PRn8ew
CmFJ6FBX3/8T+g9P2K+jwPjVCCYiTqqr+pJC3XwRLixwsPfDeEXSsJXEddlhaw9M
vQK0gWaYObIRMBt5wyvCUw7Cu3SxL1gWmr8Vz924PJfOOM5xsWC7bogOSgoLisEJ
7/iuyyjt7i8KwZ7cM30p8ClnEAX1d0UWLTdJxXSduLHpNrZR8BP13IYkP42XwJJn
gYFjBnM3VSv0XebxAw7X7A==
`protect END_PROTECTED
