`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m6N/1MDBhXFuij0z/LCC0ZNlGc/MFdxddozdSNAQ2WKk1vrTH9hYEyaS12/joi5O
bzlncFW0AX2IrS4SZfTlp7l1CE8sFQcDV5Tmq1R17aN4ED0Z9DOF3bRDbcV2VJjg
0b0OeY7HdjoxNqcKpjy6FdMO5QajD4i12IMMVbDQAtSh/qx7gpnJTh0I84vnKGfZ
4MhZOqV9J3MHZ0JcL2YpesPKDCyxC6YvvehzYYDBmSMOiQ1NLodSLW6NHAUHm310
wHxar5z0SlrICZ3T9YsdA5Mv9pxiUzgDPF+ze4ueAzc4++NPIS34gPd5SYdW436J
pqIvzXoJptqnN3LokGdOZ5tPi6at5RD9SrblXPj+9wMduCg/vg+4emjuV5riNDym
LMReHA6UytTsJFYlEYvlheIdJcGEM515YVfE3/MTkaEoNFb7cy+S91GWTElv9kya
gz0yUqiOinWJm7CKYkYfejbM3tRoY6RtnjMpYGe7iPHZtgMZTjKtTdggkTGflPm3
7dzEkBaXRJkh7JRmKPEXakhCCaYgDRL/BL1padiDQJE4u8V6iWaCyQleDHUekVuO
ARBvKentW5D9Kh913w3DLbTKKqRMH8GBQCGOrwsaOS7m01Caw9z3xFoqs2GFPVkH
jgrEBW2dc9JJ0nn4Szfm+0tPAesRd2UMo3vrRQbRGR/Dk4FOwI0s6GCx3q6NZMlx
0FomN+q+h4Gqr0jumd/qW0E8YWS4U+RFz4xejdBxFhLkBguhj/kSMSLOStGeab15
Cmnu29oJDfKBrPCI2Ku6R2netMxCTxHJccRcsTDf1rv59BlLhcswse6tVrtZewvR
X3rJLvsjfM56K3xBhW/VtnLodA632z3ZVlBPFu96DOO6WUHIHvAlFOzJdhxwjGl6
aTbDEO8fLDNO1EOEBPPuS4Rz276+eTgnRna9qoAm1+hH8icQPnc6XQtHZhnu2Iy6
JalJMzWGxNThAc/NnKZW7pj5Dj0oVWbQBuL4DT/UnLT+XrZpcFY30jvNZ4Ej8RRA
j3nFFwVILbjHwgIWhmmVTuMukVc70OdUym+P2RKKLZHi0/1QrnKveBu8+MNfRA/6
IRfuWupMvKEZxV90LRgzJNK/8LgVZsASpbzH7Est73tBLOe0f6GKqGnyCA3aO2Xq
BNo2thoENq0xhFzA1Jkn18QgZEUsl7dPgGe+qDQmPiptGs+/SL9ZDjUra01WR623
WC3Wt6wTrH8LAgCm3yAU7Qx4gvigFA52SHGEYxflDN/9snHIBLtu8yxPGU67lnJ3
8/txdM+fb8B0/POwzXnCi0XVlXXG+S0NpCTlRJ7bPnmTHaVVfVlQpMIEt8YX4fNj
y8+vNNbQwBm1ol0bMOMARZ0X4dagij/eklRoD2t+9p00RBC6p816yTUByHYiZM1U
Gow20S6ugpenS4v2RydRiMl8+8vY05wNFn8umO7OIlyU/q3BwkIHEGUR4ExmI/4Y
O1NvAJwtQ6NEMKYS97CUe/l8AXwMrstKZSgzHgRXd4L+4ujRWEHzfDfowV/0O2wW
1Gc4y42rPDIRX8BDDXd3EsnI8c0at6H67LWzVzWOcSFtrRgsOFjAec4xS7lc/I7l
IKZtwElnSlt8g6xE9wJwGNxB0LLeK7RPIEBO5ck4/5IlXFVbxkKlKZJwTWl8KGXR
tZjk3LGAklmFnqSLlSnjuOmDKSUiBndY/ilguN+d2av0vNRRhvxseM87IwR/cxEr
aZSs5vwjWG8uuz9LQCu+oWEEgfYTMwCy53TGdoN5jjkhqyy91o6U7p2EqeF2KKQO
0AUxCKGMhJlLBNJA0IkDydb5jv/Dy0UDyzMK0UfZGzPbHNBvz3LS4abEuKCoDXLF
t8AQ0SyZ5V3/V1+uqbpTmb1hoL6yNdL65xrYja898dnopFLEr3Hi08FmlmpHFR6u
hhQzexiP5bYihzyJj9Mrcr1qGxQsO6HlZmab382vNMqpP4OTvq6pXZQJCkhgHfDP
u+HdMXbyddwBwqzxeI538Y7BNQLf3IbuelKiSNyRXzI=
`protect END_PROTECTED
