`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O5zesXtjpZJcp13nZCUYomuLZTWKblXj/7kwoqktvLR+MdZ7vZqqvhiXXIpF+r77
U5aJrEhgWU+9eWCUbNtcGwLi8UYPv0Jj6ZJRutsYcYZT29b7teYMiXFqcqJAWfg+
j+mtbkg3jLkAasQ8/SWlG34NeQ3qSxJ0E7NktLe0ZKKLSuiwZm/PCD7Vr6uPsixJ
I+4iXAwe7ZD7l2WZdxjwCVwU/QoLp0an9iRNVNdHwePtZp5sVej8nq0maMgPLa9O
BXzSviOb6iuSqbfMziwz4Q==
`protect END_PROTECTED
