`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiGWTn2w5CL1VS0ZDctzLXvZELGnrQ6/q8t1cmNCknzw+my76ZJ2Jgusl4BvGfVr
ooBySoMcFEvx17y4LPQ+EAJv0Vp+68NLeUP3ZEofajazdC5zzmkNwxUE/JUY9yj7
ub2XRIriGzigAig7uahJ3D9g3vIsIdqyUX0BBvY5nrwsvvAt/ZSWWs3zJYSnJOj2
BSghi0CliuYgmEMxT3Mbqc04qaygxSrd4nPTA0/RMi4w9h4HhSxCtC5zDMRAq0C0
un1nGKlhP1joFeIqx713XnPaEvUIVcfhIlyMjdldaZ3Q+oA/wQZxikWZemdsXkPj
7yvwmWPnm9ICVFwMarmdD8hendnm1xd464O8n1fB8LZQlf1TRwgVaaR9WjCPxrTf
`protect END_PROTECTED
