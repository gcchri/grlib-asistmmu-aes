`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6QD93uf/+bH2NShynlQtVCdk8o9lDxygcaKTcIrqEACjj69fDeWS0x9NURNMso85
SeLy6VakcV9orbC2AcCaYj4WBXan4D3o75TV5sfI+4JpZuV7ay20FTiJtEdzRjMd
27WH+qMdimmzseTJIdSeRf6r+tHBcKezMain7D/12FUp6f9EL8dK6q7PDavA4xyr
3Dj3venuQx9JjjfFHyMYcsydpvUVYEmphaMXJDywAZm15EkE3ohlWCRoKhvJL9fk
XMHB74FBcF+rI5iFHA37kQ==
`protect END_PROTECTED
