`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hijGlvnciLAKmH8pOjxj+ukCtqLdka2+6coIdfvlmXz2AfPIa9H9BiDA0tuBdDtb
N/JmriYVBr5W7cYyyc6XZYHqeqd5ZYDgw5mDKl9G3coxzHCx9ow/3wnQVnciQe2z
26BfbfwwU7qPIl26VxZ+kaQZc5tOgnGfMJ7ZYkiKCxiDmWLwbkpLmoaLS2mE1jVF
1rkQGe4jLFMcrHK014A69W9rFRSMom21NAh37R8Yr3U4bbuMwwD/JYUuMLox7FeS
3GsoO/vNR3QCvTdL9XxhEA==
`protect END_PROTECTED
