`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILOr9xDEsDORx0f6yZI+a2wOraN0qEoNOMT0k86daxLr3GbcGV+EybuHosxclL3S
pyMduB1tlO88DUsT+WzS3vq5kJ35DhbR58DA70QWuWoUYx9uRY6Du9A7LLpyWT19
0cJN8hgUUXgAG8GYRSUk0IltqQgb+jjhJewCwb1cDtDLPePlzKQAgbBZ/qycogK9
NnbfqDbnFxkMqhJ03qE8wXtwMy8Ur2ZdodXvBRrPRnpIlLeREeQ35Un+uQUX7Cqx
VP0M3lX3fAOJpKSBG8lUjdYcMQMWlS/JeR87o+AIRs9PRW6usEz34HlVeN3umz1b
`protect END_PROTECTED
