`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
181kFk+PIJVCXiXilZ8uL3KD62UJlVDEllclPqa6PSaxT2996FTO91Aq4Q6Es6eN
mtF5+hbWVg7Xq8BXcQaPfywZv9L85qSgNcnGa5JZcVB8v+Fq9/nBRxW7cJaiLQZ3
NN6ducJvEHPdk1tmjk/kxZU7CW3G80EG3pNT3zjGV/n53cSVpEyPRsjaAkcB+WoP
HeuKB1Kq6X1kTUUUMRrcu9Oz37B3dvJw1GQapuLA9jLyZXw0qJxmLLecCNNOWu/c
yFqwbn2cVwZdokh/VFBX9+Efj3OrIraw0vYaJ3IFYP8A76PhQxlROawe1EM7bWfb
0k7S7tLeCahWt78SVP/P4nQYmsfKrjC80/FIVewOCQHaEVJOYzFDcqUGLFIAYPsK
oirJdEMkidKbqJRyAmpfj0ZkuvViPtxGbmNuW8aS3GMpOttVERQSKHNmmR6Di7Ij
rmQ4iIvJyUwV9hGKZLGRWYMc2wbR8wDlVWyqgL74E7DfhZGCbr7RcClC1uycp5HK
tpNvLf1DxQv8/Yt3rEnDUg==
`protect END_PROTECTED
