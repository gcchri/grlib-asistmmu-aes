`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cTkHmDZwVr/zOo0S3nQZNqvvJXkK+ACrffKzaM6lzugow7ys5Uwut61G+k+Eo1js
n4WcWYmAfmgdl5bu8nkL4CWUxEyZd2L3ivgWdHoeLTw9VRANqcSo9ZGPqj/RhFdy
9unbsJU7/uiSs4ukk6Fba+oBFJd4jxMzZeW3EemrX66E880nvQgNNtSAPJEifeVb
jVf9FeLK4skp0lUotiwj0T0K2Nw0WlmPG8obQdm+L2mcxp2QNP+zSZTytVC8qztQ
w4T+LcesUzIJF/vMuvZ1rUzTQfVCz/1yydeVpGNA5SYRe+7eYyfsZaLYb6CF/k8Q
ycVWkexvekp/eHFcfOzo9n5IN+4a6SVrtLaMckTtWtEu9cD9HMoluGoehLmHl3XF
8U92rF2y3Ld+k36+24ICNDLzt+NDAgyIXH41BO0tZmJqieI6Em0hqhfHAC6LozKi
5Ve0GxTbystO1WhCko0PtLc6xQZEuWEVcCrHs1JTachRHUCEp2y0JXXSAYoxCanu
1CEYRdKjnfXDvlQ4QmRG/g==
`protect END_PROTECTED
