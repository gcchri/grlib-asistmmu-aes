`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xlEtgZGyja6gsr2bqDUliVuuKkZ2dsUSnzfNL8Bq8qn/ZyQHFspqBsoUOgwZYsfD
N5hXq0UKTwAfGhGdMZNKWWFRDKZpzxMAFG6w88Y77uwgL/aVmyeDf7vES1KYr2OP
5GxlEaHaFs8XeX8XPHMupaUwBiwgYoRH0wNaVgaN+zXABX8Os4XJ/mSFhlnToFu2
/DHrfZPdUBpvURzxLIGt5Kznt/tl+pDPkznGUoYxz3bPtUAu7jfjrWa49S8Ok9H6
LvHVfqpo1+3bV0bST8RK+nstbQQhBBGQG/GEU4ohy+qqxwD11H5FYLqVLi+GgV4t
AgHZQW8E7k1DfOHk+z0wVw==
`protect END_PROTECTED
