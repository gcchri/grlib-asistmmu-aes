`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vAigcgYfzfMZ5/SkffPlZ4sofJif2Zgwdny211H9a6cNJ1+JWpgvH85hDgbfUZo
Xlt7dJuWw4CsaoOgCVa3Pp7InMdCoB1WPDhgFxuI5LANzHVO8TLPWQTtTEldL+AT
I8Hok78L/Cnl7ZPwimZFlbPH7/8/SVAQhc3+IFUd55iY+aNKvGmnp2Cyur3s28Kl
rhYqFP6QBHd4tQLkIMdaHdGC8vPdZ6VNm++yHn7bjvdgqwVfU3Wmj2+y0amj0CvU
VARkLbW6Nx9hrCxFrqoJeZnk+9HMlucqUBtWy0xi/F1+RgpuLaeAG5YfaNeBzljp
Zg4oXNzPVUkaArfONxgtHDtDXDT+blzBrUD5p1tcjDA1Ka7pU2yWzB+RQ3Piw23p
/Gf0U8f1ZeJhabkbo0neLYabWPtlvvjOwTJuBt676y6ob18Xk5OaZoSGGvJg3exC
dB6JDr8H9l9KI0f6Kkl1FRmz38tmBbGdt5F6L22R6RM=
`protect END_PROTECTED
