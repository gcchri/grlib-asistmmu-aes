`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLiViIgLxoC1rb6yYMYdDXegT+CV2gFS07gvzG1J+92BS+FyJLXPH17AedAqfbF/
wKhsZj6QkueVZWynylEizAfLoQG6IDHpMYUtDezz5b5I3IXqQNiLBqutxf8+WwfW
JGG5VyO3QKr1Hb9QOr42Uw0KKBlk3r5I4u8SjdfG2uZ/yW9icOYOq5FelEzBYSi2
8qsxgg01VuZlb/gLg423r55L3GgAVf8BShbObtPjgY1r+WZmy7P5DWwNsAa9bs/O
caNFgO+yHKoQPkWGxhFs3EDt5j7RwrUTgker3KLGCz2UPxWTFOiKON2517NNHsC2
junIdiS49H6zI1QbBx5FxqAcmcYKOTWDwCNvjNK4fOMbuIiooXsPO9FlIVF3X2da
Jm8FBchZl/CrT/tZgjLzgqaOYF3uIZrulICws7tiefrTIVUnvavNkisqUTHsC4Ul
sswpntxQFshyWexTRAQqoh5hHLfef82NVH+5mFCD0+E8AFt0zUFlk1KcZ2XArW/m
`protect END_PROTECTED
