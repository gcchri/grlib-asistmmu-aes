`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HypfcNsHTzSRn++1axQ/H3DmKk7yyt5rFIb5z3erVyI9e5sXeZQPnTbQAPXQSvNT
Q2ZUbAybuqxlJcA6KS1UMwVsRovyHuYro+spu2yrkI4m4UqgbTQoJV647U+0iJeA
sJuhV9e3a1qw4Lco97hgqx+sHSeQDWx8rJyJuS4WWTX4M6TmPuG19szHls4TGrvi
Lse89HfdnXPWjayfF7qhGJlIJ9Z80IiUJgzgCEd8bpi9oVuZiSgUi3Q742rXkRlP
KJBlw6aMT7J3sn51Tmc7lg6JCmih0jK8gsZatAd0FGbLMG35uuaGKpxg3yMxbxWz
`protect END_PROTECTED
