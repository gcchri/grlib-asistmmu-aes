`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+z75AOiOZLaJjtW3945L+QckZLY6PpDGAjd2bH4LjxK1HnmF/X2xn/IiXkwAEhVF
qyRCmERtczH7ReRkD0eURgOJUE0U+Dn32ITB37OKz6f5zCbUgrb6CY4A+19W+xPD
JTUr1n4UY4skReuoF5y5Yb8CZQyua8ih+TfmGhxK+gm0rYmuVVMtbs10/h9kv1Fb
tIOz0S4sQghLIXGreOFjYkNiSl4yXbB/dsg9MR9fx/3Cg5DW3PZOP/xgkKKKvybG
apPVCwbWRPzkG/kXM2fFwwGjTcuXoVrpZbeE8rYj1KMoCWLwy33214iW2unJRyTt
zbwJb6FGNIuRbPtNrIUYbWtWNLkJ0iXFylih4Nl5n8Aih+dujGQ2uxjh5stOtyFg
wmvcOtVgTtuh/deYUxiS7tBSuGf0KXSAjcigLqtVrrRbRiMXOk33e0DxmM0TPOcp
z3qvznfe7e53+DbUICbKDcu9JJ81yw9YrPJBOIksbh05jSeirwZa9DKqsXuEf5Xz
U/Y0XVL/xvW5PrE0sreDXL/N4aD7m/r/+vWQ9Xk7XRrVxmFvoEJs3Hk/ODGRZQV2
zolmrujtk1pGwapB0xts0ucFIzOuzfU2TB6v6rc/oPl6bJ2KghXJ4e8xq+eli9Kf
Kqnmr5B87mJHEK0yRD7ks9Mc7huuAte/3PhLN+DaR1FrgMEks+BhujZYkxtf83X5
KaUFcUffMi3+EypYTPEao2YjymLC3enT5mqKdzMZlZk=
`protect END_PROTECTED
