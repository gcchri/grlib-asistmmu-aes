`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p96oj23f36AB9dunpyOjtKTTo2lF/M4PcgMpAetmP0kl4dRD4UxqVDMVWBv1dL57
XSiLNbmd7nIozH39Z2HCoY0/VnNh7iRCLeIKmq6y5Fi64ismHpMl5wjH3SuCb+8X
llPKIqJv0LBKji9vyZDo9I6rUS0H7HCHQgTEFAb2nq75+wYgpFzbMhZ5BVRSa6NX
Z1yNjYRUe0INK1+PXrFFRmgfEGnOjygA2xPauoOcK6CzSEjaw6stgY1Czf4y2eC3
plaMeo6wxgl8x1pZBLh4cd6EAk9oBGGDqrd4PR68iusThmbyhVlylx2Hu1VnSlHK
k6rs/HYPWmeKpOwMcWbjBBiNlFk5f/Bg7d9Lqht3SOXTBi4yTTttUhB0Kysuh8wk
5s8wxJgafZpVzFWAvBmF8T4QN9p20asqpuduTFKWMQmam5AWxYZHoxruI/IrcLLY
CNCtb+J4dUSYM6cK8hfJqLjr0lJuVYy1waxQeu2wQlaj0R1wQk/2Gq7use2LWGI0
TsgzRkg3fLf6cHmB2oiNDlesF56AV3E8dlB6enJdNLDRKz/6XOEf/Owm/FI2KgpV
LThNvvt89Jq+UjPcl9+1X+07wiR4QHfyZ5xO5f5OqS7tdKcYRJqM6flGevHYJq9V
k02voINTJn0zRGGlmSUXLQFcf9bJDW1R0h5AcZ8qaY9IKkhkarBmzNE7rHHl1WbE
NUIf0iIC5dhhU3XXcXD7V4zEAeCvD/1mKLjTLWQHRWy3lO/B46/XCgAIh8e15rLc
Pr0N68yBr2C1pNvl6LssRey0P48UtjHc0RHbC6djJXa6PNbZjSesJAYkvEX2WhO9
xXZOBEBGDRf7EiEiCS5Keh4PTh+gmJjP/rOPsRZTUJ77jiSU71CWeTyhS/J9UA1t
Zrd73JGJHnFRt4k4I9ba3x5G/0vY0XxJpyecDjjTQrxxSBtb+EdegSohJxYDTcBb
Ojrzc+gERlL1UA0x3yzEukCNfyQRpSiAZ/lY/PO5xMecBD5s6HWBax16qD+k7Ta/
rkqt/q7QiaJs7GtCkIKnECON3bSMgKuMAaPQ6k1BdtF7uQ/Vatx1ac8RXTQ64IVr
K+KhsYXvE/KvuOaXw4PWRWBKgYq+oqwZndny3kBF2kWO9pQHeodgaZV57uTeNnCj
AZ19cIc9NARKnsIBOBqKka6cjdRzIHGW+lZoaRPorv6i3OVOcDg4Fkn+TVBMm/df
/hTAls53UoBmz1tLmCHWsjMtG01AUPU0jzJvEnYGZ8+MIXpsByuCACd/CM8FOlVm
Bc3bsc7WCPdVDlay9gzcSu2VTM5v9iy9hNhpngB8pMlQwyQ6/xKPPFAB/S9IDGX4
IufglfuHB8nOVSW5kMi95SDSZXPhacN26mlHzvS6ICybJH930+ulSHTTHJ8Y2aad
AQt8wBInFwTBvWdI497HnLgoR4jxO8LlKkhhQrQdGMiI5EKGmc9cw8JzcGGihhqB
`protect END_PROTECTED
