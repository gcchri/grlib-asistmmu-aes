`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i/U6/U6RDbFTajNd4oJjyVm63EbCiT2GajyibwBWbRg4rAK6O8gLpsqM2BsI7F4X
mdDckh9MoA/7voAtBGIU8fYdz05AP9vo2Z3u7f31CdGBXnokF3NEG6iRLd1pHsJ1
1NAebXzEsClcZ0BK5w2vYmy5ZbixA6eyKDATTFFEbpBDwYd0S79uFy4yO9gBAVBF
mbxRYQ3lBR4dm7hSZLjWxpgpEGZiLqfi3l+lcOjGuYXCBnF1yqHs2yUWiraqG08a
lbQ65s1n6aoCmNYkLvbiiMgJT+ujFxNcDpIiQZVBhBMENqdGK+F92TMvUv++gZ5Q
G4WTU/qIjd+/cx4JhGm4UqNcdp5vgL7FGh/9XqoPbn+bGjePjB4Js8x4OqyDRoQh
VuNPm9/yH5sk8b+nrSIZK3Yi8Qm5WXg2D8X08dHE6dEQerhM3kmPK36KYqVsdxTL
LREhoVzpuW113qNcZxvd4Ffopmhe3KinFbUmCvkSgZRaDsDqlBmbDzKqsYrIL7mc
nTrGRiWh8t4lqGtCuOiBOBOY+ryne94We3dAg7EYtZUEB61FDkjoxzmcyvqIRYLI
eEZe3dmGbJAYvZmUKzadGenhoaBrUB1WCMTvNIIYZPhrJXPHHcbgGwjU7yqMvO7s
XxGsm02l2HhKWWWHp5c/sfnzKtur1urQtk72+bW4kqFk55fAzUfVF3yflrJupfBg
RT6a7g7OV7Z/S7FDLsDzii6+oPdZJU78tZQBBxKxJghb+WHn6PTXjB2eq9o6Otzi
VuFrhNiC4pClO5NxMW7TqlzksTnWEmArU/O23upCe3JkLs/f5rg7UcO9Wfs55M/6
dU5Uea6tileJ2C0FhY2nLbgYTCNZsuvOTW3Lql99r2jQ1Dp3Pc6GzHHJ9fluMa1D
1OaIYtIYXFQAaoMwQprVh6pBDlCfOcPvVVExbEHW9FYyqDJXtckH/Fs9y5eA/0k5
3md+oFMpFtYU2I8h5cj+TjFm3qEPavb6IOJnrBCMcs3MYN2x4T01vCPOivjbLp9K
2lEjC0smxeICQE0HYAOrgi6oVQgUYXOVSypUtc9GjJJehxCZYaMMVGOATczQ58Z7
MZdRkg4HyXdUMDSjYDiFhVG44SYhfs3u7IuNg+dLaEN3Kt9lhKSf+OIf8FvAAq0s
MJTezqUbp3f+L8CXG0EdY0IXOQ5TGwJAcikK7kHZ/Id2P3zEUfviItETmNgYewT7
GjzbpfResznTb6l1z0+oom/WBCQ4jX7c46ijJ7YzHS8L+gc4z3vxA2Iby116OKCw
MBrQhpUGmo31eTsFj5mt/mH8paDaD2Tnhq+A1hIcFevX2092w7T8Wt4SyRtBgKru
tJsKzF6xJ0cgg2k8E1suxeUWo+HIKI50hHqrmS4K+TIzm1My+DmJbX/xKDHMhpdN
MuwUOw20WsaZ7npUGZm06Rm+Tmd/ZXkv0XQrUNt6aS/zxDlrT8Tm4TqYeBll9omK
Bgaa1V+3RvABE6vBti1ktmrXQZS/EEM/TLlqigI1pHON8ugkfWKaZvjCsuFrtmW5
m+RLg3yTqhfnIceMiSg5YMfXRRBspHUpw2Dlr79eRO5XC6GR7IJduOwEiIZpoDdl
+bI8QFnRRua2Zea3PlCTo/t8LxEDiR9RVdNZVfvE4JHuGaPcSxFX162lZRl64IJ4
Rqc+yFrFu72cZ9Smgx/lTYyHLghdkg2dnK67WnY0HyawnxZ4ceytr1RkEML+Rwun
4LoH/kMWeL47quOggQQ8MqJh0aof9n0egrWhrXV4CpiXkCCXdLiwi7pNkvU7VSUy
qn1twVRCL4fof2y+4g626/hwAkFo6mIDXWNJZJRUUGRzSgAYr8YNU/WQjF1Tm/ej
m1o0K/ET7q4l4EvEyYR52VMufwbv6TPGcyKwpC9SV//f77ONLYxJF4LXjppraxgT
W2HxoY3ZJ4ZVa8QqeHnxMgPegctDOHJsp3xWuyZo31LSclB3sBMQ6fyhBGkPET7N
lZMY6FLT7pQK71JTx6+7kbK9ipPAN3Qo5LAxmTEIT0tfL36ZTJSJfMZWb5JiYJlC
JtkqB0HMGOmNHI8r0K5XJ2YNz146Hw34ZdqHDlqfxYynApDvWVmWHm7pKxLuU//Q
7uyEqCLfrO4ojMDih9s3nzSMjJ6G02KNLqcTGpo4LJR45/Q/NA6IABDrvlgwH6cy
DlHfBgYNoaqasrH8143GhniVqZyV1MgN2yaKOYzr4rQmmx/F84UN2b5MsEmrVBLU
WjGQOqTBA4YrWgKraLMTMEJQUaVZU6u/JvDGH5Rl8zgsBSyyZ3Kt0rCcD68vEXan
LfcnsjZQ2qVRTzHwX+oKlRb+kIAZ+hzPT+6DiJ28lxDoSgFev5w8pL2cwEnTmCbh
yE8g1FlIjZ83hOpSUvNApXfS8J5kFBCToOX3PxMQavx2FC1VrDlh3dDaFRc5mN5X
MEGrT9xvHMeaoz3zFjNKL6TEM7Q8rHf69vdfBZOAj2pJTl8IDsmQTciFBLiy6kWI
8uo9wb3mBaIe1D17xcRhwDp0tWV9sYpcC2wv1v4lLMN4OsgV38V0wSdNrcUh+mvw
fkf7p0UpuyZa6Ki/ZiOcUqdcaW5/qFXo0JRJD5p53UB7hQOF4+wgIvKcU+cCvJ+0
FwRLMkwTF9uXqzbW1qW/sXLVdxZeRznHhveZxcxwm42gG6e9v3TkoQuLyuwH/yZC
AbwrsRthcSdevHV9by6VcCoXjTjeQDHPXjBsP4XSJISZi5YoAPi4kSj01Ng95PuX
D5ZR4kwE++pmYcw4hAwFzQUWPoy3ddpwtDfNUH9rWP9NY5b6UAAaHx6hJFe7W73H
RCz5CaBbgkUrGVHYM+lVLAxXSXqwXqwj1+81bgqkKqjUnleFaPFQAdosO7iLgz59
k+h5JMeHVRuSP8G/rU9jnQ7VmIyBgs2ezyf92ZDoN5I4ABZQLJD3ApwNcDL7BzIe
vJRUqHe7ppgUqtSemwJSfmor53pmhUsnzY6U2I8Z6rOK7ejG9HheKTQsS+k7wVFj
EyL3qLszQRrZ2K+vrGjqZdYhdTTQCO/VNthtpRg3zO5JfhuTWdHzBzEXgqtbWAUL
q05RPhjlGSa92YfH6/SJGk6jRKShzfllJedVqSYXUfbIo4cujCUzBlIXA8easPaG
CpJ45CD2XvJ03Nv0qTMJv0xxh5U5FQCcKteMhdHInPMqiz6ev/5GRQ5SV9oUFEWc
TRtQGMb2cUDbIHomidwN4xJIEmZ6P4kyZdSQGNr1KRObBrqB1ul7akTXDRcq+6Mt
j2+KRNLB8j2I+Qd9pyI/d80OR4qW351uX+9Fnq2HkCcNbTy/4dbJNpTiNnVyO4D7
LrceK/BtS2nzfd7LRxwK8cGEGKfzTP1EqLEJHdfoU/ecFNZwFLmZxt+7XpiRBQSe
nIN2s6Hh2C06shLJ2+xoBZal1SGLQ2g/UfUlqVKRtBjLhpVW/O4p30CcE3yvkxqU
hQz2lp3+ANY5d0QOF26zBA/b3TGm/BzT1Tta7qOhFJrMGRUGeuDfeuCVeFh/+HF0
A/L6kGMt7eR+e/lu8MCl+DYN7yhNRwB8qAuGKPgsdJ1mFBND8D9oNp6WDuHGhQ0r
foxvT1MX6/TDgLm+xZ8dUpuLESU+znmrGCmpNW25nUicoAoL0FIHrMHk9LXNMug/
rYN7rbv7IPQTj71Eo79QiI4rUz+kiYdkItWsLs+SAxHfFV+eWN/+hQBrQlTAaV2r
kMzSVBsV9WSyGRDmw326TZFZaJvkz2pmircEHl9pFBLsUZCP1wTcAazu+Hrkxn84
EZ3qJRlC8uymBxP4y3z1JfNJ10ytDSO/jLNVT9wzCduPScQa/ug6aTj32cpgO8dy
WNEgQUc5581T59SBHkT/rcQj6Sgfnkq2BFuAcoEmJShGNTLNdK5CTyC5l10Dlpi9
e1NyUb8IAkuatvGiPLpdIeoYl6CIu5j4MPd5vyWbaNv+ls6Xj+XVsSqyOUmPJfyr
HDTjlQyFPS2h5OPkupnXj/+iqRQblrxZMxTUSFFmfBLY5K2+lJ5GN1e7sULN3350
w3LAjN7+sZ7UP3YRNC1AEra6zX2Oi/1ico7BNvz61V54IUXgb3wt+RZPtaU6F5lE
sK6HsgyPq1o9XOAvVjHB1PIs0X/mZobLs8Gk11hDgiBUxqeDU/Am2fqALl9sQ+r9
JLrspevq0UyARKAuHJnlg4Slq7BfYT8cNS1uH3mAG9fvSvKF1U1Tu2aYgMHllTed
BJfcLHOm4Xffg4rpNEzEQ0TV7qmV+ejTm1mIVxffXhcxq0T6vUUwi70Zx2ujQ0cm
qkQuPn4X2xUtjtyjMvLmuIVb7/7OcvDdcNrTt7w1YSL2p2I4mBxA8BIRQhHdD8rL
9Eoao9878Pg2YO9Dx5hMnSTTl1JuOlFKDX0C3Sg1iywsqbFSj551+RpLqvl5H7iJ
Rph9ZMgkSxgAXsYHu4F5hD+olmSVX0yh86DCIPsaUHvrRViE+KNnHDMw/RtJGEkr
HEDjCFOEhw3NCL6o70Joi0DiXYTNGcftmWPUWn4jM8CEzaB3s7/huQqcVDjE4A63
+2Zn7YnB5IwNYqxwQxVK6rgaambKL/fqyv2ioDA3Oazd+/5gf3oZxtne8exrV4I4
gtfGOPpU4hmH4NoEBN8UlYti/Vbpyy4It5AmKaxCLapw2Bo6B2sAC88RiW8Ov+Wc
RIfWFjJdXDxdeFDDpQ45HXf9HmxolDz0SvDMCZy+3JptCFKZpYcW6dMZ8rf72mAm
GzTUmg/sNkE9mgagieyIijx/3LryvHTxcIJI4CArWO3tt9UbiYV3dYuzpWfTfORK
8+2zqKJRfiHvqRNgMqn/GXQxY+r0CQ0IRBIeYbeI6qP4MOIuvP37p7lrZDamPM+q
984TI580leKji9X1OaUNqmKtg8sthbTSWcRxRsWgMdoa2KH5pIHEys59MLFk60mR
B4EckNro4tEN5VFDljUjtnZFu9zf6FK0WyOHKB2c9qpsQkSOjoopslLhEWdOTUTI
/7MKn1c2TxvXckEBjWP9XsB1TKMogDrhGZ60iZgWU097DFwq67lMqE6+6FSFw88M
8xqgxyy+X/zPSxwQ448jLJAs1+4Xx8c7kgGC54BgfjPx4XRmuaxRPxQB0mbfbcnv
+aRv928J2AJU6b49Fo/PiNH3LbqRhdWhUDRZY5R6oQVUT/JO+SAnPsyLH4w7NmB1
galUs7CGm/d2X9sNvDdYcHxzDZEVkTGck95ezuDynZg8b0fBMLZ3avZ+R9/Mri/G
qQ0EBgQvIr95mWodQtwYLZhTGTKje/lM2BDXxzIoc5f4uodGEBw/98h+bZUxDigA
gtVAtzgXYvPWbVFyPsle1Hdh36eOLaVa45GuCx8O3/M/51Fgnv3E04VEk1O2cNqB
qapYAandf84NLDMdm5GYbxqKbPwOY0gFAriyQy//JmWosPcEWqP0ehAxWPmo/6f8
qd2brPGNzfRI8gseSfOJAI0lhlJARzRynjsDV2nUM/30MXATnmeISkmgVTgWLuyJ
UcenfAea35K+ttEyWzYCYWnf0gZFr2ArHf1qYkqArno9vZ7v1z0+ddn0gq/OMSty
OO0I7UQwn1FvfRKs+1QuqJF5VSv/lfCFTPe0LB7qfDT6G8ezUxSLc7rZPBfZlbKg
2Xu5/Za1j9C1O+2kqfqlXrqm34JBBoVyG0uOY6HQQyXYMCSlqN1964wwvhJz7yvE
PWG8L+zCKn3uUE/klk8Y4qJXT6YA0Ks+uwvYB5uzyzsQ7WuaV3C8K0ttLe4cVEWK
LKIlXlnVKX/YbrZgZauN2WmFXIhGHhXP0g0y1dxCycwoBinWzZM0oecP01kztBKN
STRnHCln5naRnp5UEaxrsdSHlDjkclxkUNJWdmu9RoWgrROsNW1I9bvnDV8k0PyE
WxwY5MZ2431O9S7/dzGizXR9JtnTEPgpNTRuP0G6JFMPSuZPBQzXprbQJzDYPVBl
4ZLmetDVXfbbXA1hYgr/Jik15NLI3EDoPLnjyjnpbaIaXa9sTJQIGeveYeE8TxEX
CTQOpVHxyNFLzeS1WVXM5qoa/K0WppI4JTJXbaw1oXX9q6KqaEFXE0vMkIkK6F9W
pHgnkiG7+7jLjG56tVRIS2WRQzagh6SMUnlxNXP8clWusmxet1vmelwhcumEpfXb
6BoOR4t1TWG2tEPEyMMxKb8DaMz+IoBHEkwTNvpyGhJSxYJHdG8DThQXs9ZJbbqY
gVPuDYB/ZftHfBTzJS9yLtWmNuu2+tNSPgm11uzuWK4lV5BoWzg9dhoxzElrIq4j
DeEa+XxJhduKm9ydAmX77/sXfE4dSh7gJgHaoeNZieOQbN4uztMt8GmhCeKX57Cn
tqjakuUdHyfvxkPxy33t0cToPIkHme0eyP+6ebtWE8FCkyjuQ4qFKXh5gtbZKdwE
LMZzjXrRL4uETWwfhoiQaihpWbo/6Ueu1/sDXpuMVptkdnSx4SaV1aqK4+tFxeWs
C1ivINI1KnHlxafuOkyAt9QR5rTNNd+svacaSWCKyPD3/9KrNtIeGoMt0VC2+YnR
8L5IRAS5nqlD1cPpKQmttdjVgr5ZgqUYEsYiiwwtne9uZnNNqdNfB9FnR/YzZrRa
WPAyMYJpToOJH+h+2Mvn+OUHZ5NW1d27vN4RWTgaCJHTwYuiJEA2tsH2FwAff0LE
YTstO6KakWA3rW0Qii5mpFkAOAEjdCWM75kBdiJa0D/K1alc4+raKAmS9JSjqt2S
68P3xqnVccuT2Ea9GH7RxmujXxFFefE7d5rb78I+AtFTYDmlqX8s8EHYnVp9BzXw
uCZMseA0qjVu+R2Uue0q9FAAU/8HbNO2VbCv8pa9FvrrqPVg+pc7aUnIUtQr26kC
C6VMQvKAhRijlCFmY9NJI+r+ZfCO2AHQB8QafYWsdAOggrME/R//Fy9pFHs+GCyJ
iZmpqGKNZtSXCPjZHYsnuQtCV+ppOhzbmDRUgg9b8YYzcmfmKJfVzjVRFHlYY72Z
GjXMyqDnvFC34cbQJxM42wUFFmxHAow6Yglitk0G5vFzIaNmKTVJ5xScZxB8dALm
M7K2q7XHt7DEHB7hxZYXY+Aecw8+l1YLoCcRfozelQG8c6ELhp2XDYsoaou8t69v
JPNHb/6IuyMLQk8mhoj98b6BKFksUSsdVEWODGHSPuJ9/MljVGsE2slNIkELdCnU
FXvw19fLxC/j+yJc3soO+IInoktsJtrZemgQyvEJRu2/5Hj49TyrpCfgybHaeleH
EqDbSbZP97uKnwKKbNqmr64uO7txHGwl8JkUvEdWn4/eZX6aEsRZc7R2uhPWszWT
OTxOiysQ1P4NTH6AY4VrAY2HO7C+aCmj6qdc7vymPtYrkgwJsBycdkFzEno/YeBc
kg5aQf3APEmJnvl4uLMbOu9twAAOA5CFGKO4iEZbwkrVS9DWEkeo7Cl01QEZ+iZ+
vXAV5B+xLeV1odkZDH7Y8QrzlVltHSqiCd4fOTIsOvS0NsgCKAyKK8mkLkNpDkIv
qICYOnXHbhgXe2WW5P8ETJD3CFncgBJD8xzVStUKSfhRQXz2/obV08wQfunqSbZU
CLvnqi0DqH1drDKHguOROdiKpbq3GilrqCknC13rlXWAgz01A5aGHq7VTcq6k+jM
UvVLLw0ZQn01af4jZ1uwMowUj4B8xYKSNLiwL37sIobKiMk4RUqFURdMlbCqZFac
DOOan5GBUxuQVy6Ta6Dbdt/apzLsT9YIujD9AFDKh5oEkeyjjbS766urshSRrRMu
cp/Tt+sM1XgElkNdbya3YKsCJk5aS6Kzok0SCNqg6dRzG0HUgOhhPl2OG7HSFhCc
iZawrE/7h88u6TlqkQwGb4CGIBbfzbk+jpf9JgWsBvFM9jU9Y2rpGUfyShV49V76
E5uF0IfzyAZVsULCNk0WyKFffS/O6qQAW9Ex53Laytcj8OXUtWtyzFIikwXs2TlZ
CH9DKKsFElUD2P4J6k8A/dWfRMOHOSoNrtNzCHt4N5yVxWEHvemiCD4bxSIDXey6
hkl+4wPPkN9U/VafAsqz8G6tGRIiqHKHAjkEQttOh+BCO9PKsXS46ht7pWa6BT6o
4/2xwG6llgU5O1ocNwl8SuqoqIKcqSZBv8oH5NAiaFNJ0DT3tiu1iFOH8HMp7SNd
DoxCNb8q3uvIiOedCFDFaFvw8x3e7WnqtvXOj3DNy6/P3rp55kkVC/8cSpoltf3Y
9U9HJWnTYFy0SDMWTfC6fMgWn6lckoRkIW4KUhHiPorfoTi5p2FGQQFLLDiaP5BK
dGdaJcnlxAUgcHQk4aYsbmbBJzK68DPVylU+JogDGftQ9VYRwaZNXpuMFlTWmLd/
N2VbKBIKjK6HPOwac7zkyPuI7KZ7fV4WUkibyW/f2FvK4p3KHs8GsrmZwM3rtkPb
J8Ftsu6WU+uc8Y+UtKYtQvnaxu7oW5zkp3Lpxrtn9knFY8jMK88srhwfCg3swieT
onHWNqt4iYBCokFbSNSPOn5CKFbegDV7u7f81EP3IWzCfg7uiNbNyFSpM0ARR+6V
CbVaKLNOfh42vGbA+M+3WvMe5vg5ix9wbw6ecCLa9+EmNstHzs9kHSiOESPm/lfs
D9HG5tHtMUesD+RLIPugZRdftl5hRLvzji5In82/H+t5uyu4ncj0Uh+Au3EK4y6L
aYaQ8Sazf85pS/Pbd7ScXcPPmOoETieyYY6B4rGvjaM//wdepSuBVbFiSZo+Gvbf
6yGtae6TLc0gc6/WyLO9oqme41toLZuyUH7HlpbEqBa+whL7Tk2Ra0lHtNaTlTZY
gvqcYcJBmVQtW1ZikwXw/QApWlTApp0uImRb2Iae1pnAccbCh3uDhCxTRoBXUu2x
DeW+gD6ikrx2EF4xw4akfSlmlRj45Zpz/v2Wke5GdpxljmvckghTWYKgibrAEFOj
3Ci+JCzjgb3ST/TqPaTDjMWrVzTKF5gfbT8o53+G6wKfrPbIcDJIdj5KPYcJETSq
d2+05oQO5xp2l6meLy93RQBWk3bEAdXenQ9lZ8D+Kp+Rh0Qbtnm97UtspL1TSykU
ZKzTdKlsRRy+VHd4BLg+8X88zP+2ISZ/6lk9RYWvqUpK4nImBlvg0oecMY2zS7It
YcX5sFEGqvYsdM/WKxq9h9auFge7wb566ue+6lo4uu2FHEBW6rydSvIXf/8ejK/H
IoFuViofdNqnqx/hOKeYgnrRJH2U+WehHyPjdwZRlZUYeQCpkgXqNryaT5mvue6z
GTV9Jxo48nOA6BTfgCCnqe3LxZS9jsAPQ+9j/DYLYvCLO8T22FIKtlwZ9Zp8RnFZ
ZRvQcZeY93KOrjtYGyvoQSKcRs7KcmWpq/nxhlW29WJyJE7KDJGMQmuSbbT0Ejnx
blBNPWmdht0kxkuKAwWNp6YTsgSw6iwTldjNyj1VUSdz3xcLDu1/2svA9R/So4kw
Ym24wm+M+XhJQy4jpX8QcUrgE+ei9BoWOXxxGinCgyBeOBGVVO6uFO/ApT8hrP/J
/j7g741Iu7fIYQs2HnBDhtaM44tHbk32IJwVH9E2eFFp6Kpgm2G21ypPp1tk5VeH
1IeO+5mM8DpWAljRsV/HGTDrFz1Tmq+1FZVhMIdsKfg5/psjnCUBMxFO90nMH2bH
DvSspU8IExj0jIip7aJtJZ5DeKhv6uP+RPBPIhwaddYmLkooqzNsGlS3Sz5DK01g
CIDm72teQUMau3JWRZu4eBs5oNn8cQTjmtXlPNtm266KsTFKNo1Gvh+arlXJE0Bq
zLbLjxeqI9A9GqgdfTOVxPUVlio3FlkudKCxJ93NBYAwbtt4OzKZ37DOhuWOYkpo
6SAEo5IjXwK55fsYdDY3DlxwhU4tbNZAAyeukJcB9s4jPzlkBCaDrTFf/qs/v9kI
csy77Q3OAhWbr2zSpvMv1W8BO8UL7NFeohV4CjAi/fw=
`protect END_PROTECTED
