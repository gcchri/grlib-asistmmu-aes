`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gLU/2ZMc1Sor9lJ078PCO8U8C1R5B56laTYBZNncq2vBDB03kjbtjsJ3HYGw1Och
yHHx9jN08vAtJqLJFtOwWp5DLToskXfRGNYTjVXL0h4/5whPKN62d1m9iVkUH0U9
y8yI/7dOLoeVSMduv/OI2saRSu+ki4Hkl0YLiBUY/z6hqGZuJk9oqhKxTfXBu9JW
WT/aYo5IWrJ2virdi3klqRfKbsjdYbPFdEUFbZklDxQ2LA4QWtd5ZlkeQ+WQyDF8
Eq+fH3DKAzBejWNfpUck8osPo71xiUArLOg6P/hUoAjEglYr5Fn+ZRIB5tXCDmT1
+3PJhpj1nPMyp9D8nNS8JrPWmT3L+gQUGf1O6ENVukg2yTLkWRmPaUwO/0BN1tqF
3AOxwIuKS0Iaf1iXd3RIjKAAz+qnNnrsAag0/LmGaE4NLoowtK+EgybcyCmqHko4
lB06/YH0uTwC/aOIrs1//qGPDiOehtKjsuF7yW19zQwQQUqXYYJI/RI1WwQVamyH
nA69m5K0gEsZg0KvRhH8R7EfkhVXzJJRD+GIuGBc7C6LglwWYioImmkWXuySoLy4
WlXYwrkFL9NEJCvaus3rPSlUBcw7Kn6N3IJf5zpymuUYkZSz70wM3WNjrbU/0eHH
cDUzWY4dO6jk8TxtCN98zqDftMPVO0EZ3+aOIyVmFUHAmndSkzDDfws0RFh+gaZo
qs6LDoLugR9xcN4QRK0cfxG5RxCF49OXurszZ8QUt7h/mPQHqMeFHHp7Eb2Kr00Q
WGkIPXPJJr1nG/LQLc8cxwAqNQlz3XcC32n2JXa4clrA6yZCTGfvIlYMdFjQR4Zj
roZRi3HQbxdfhIUQxg55R8ZoLyILJMhFqjgGxGh5bJFShDR5Kn1H28GD6NDivZdO
441FXIhWHNlZi8nfdRiHc5N2ZRGaPaYgDEufpe+ErWCFp/TqibIQGDsypoyjrg8T
FNbtrNYF9xPSpbmNHfmLab2nC0E6x7XZsYrATsx6UCYQzEqWOpTb4D4vmdpxrUwn
2wsvhe/PvrO3ILmVh9nKLCS4QRYQ6lVWzCewWgIudbaOJ2xklLN68YiWSJS8y9GD
YgTMlaT+AxWgyd5J+/DzSx4AFSfaqmMfjx4BlWwcThDk5rGv4VDKbMDMXxvMQxIl
`protect END_PROTECTED
