`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLcKSW5IyzIhs8aXq2z0hbA0RyskyjfQwZfXbtksce0dMr70h3wqMzWIBN7zM5iO
gltWf30/+qQJ9eGtvSzHawmnDV599o6KYr5PWKSgLI6SRp+dgDF24w00Lh0Sg4yk
ZUFgpANDUg1pePc1CIg/LJyck4xrWFafrw43LiGURXtSSsjUCQqUcTmCX6LPzcFr
myoSzE+gFI75LTG3fL9gXHGXT/PgH9YsbplXPMyMOGqeZKlYob2ho5avC19FdReE
RihH48xACJPCpt/lDPlaXFYEBy/eMyUASgvyQCgfi0qm9p3K1a/ul7V96mIsbHvL
bAgp7SgoJcm9l41+wKe18Z116TZfyY1kgK6cMthcpa8T/KZCIfBZnXjR+2Qlacsk
vqpHquSpe7vlqbDrr6e1EolMqFQ4wIRTQUbcAdRH8nX5p9JJP1ePu6Xo62wqcoTU
jtlVXpObfW64QI7iUHLJrYAfeN9mPT/lRKR6Ea+bRjkT9p38Jg3YxOA6ki/XWaAH
kNBAnnaHh8CFTp3g5zGSHsPX09Si8Q6Dzt4+vDsL6HVkj/nKb0ceOXH1BqgJGkc7
FQwMqpDEmcOu4/H0QARWMMXS3Pu3ghbh7GPOkGBRYVpYfGikvVwp3XV8xcB+Zgn5
NaIJSj1Lmey7q+ITS13bnzn/gr189kzWwhyUd5oWv9chVzD3BgOh6monDPpwP7i/
RtoffBRl/scqn5aTevpjRUovzMABHe99MUR/CYEJzBdqJp+157stQoZu9TjXOiAg
4FV5Ao9NajI8em2Vu7joAW5ulex9V9zcuduFxZePMtaPuHeYlYwn0po0T6tdbP9E
6bVc/m0beC/e8ODOXHmu0zTvULSlQUoRTBFZy8IRBCrXILy8SjhaesjpblJfMtCa
Xt2Fmy+WwF2lxFr2+JMxDvdTA0qOUOjjuycrIduxk8PqtZSs7ZcIR8pOaMhrM1FP
W0flvPGIEa7yu/LUOT94Bg==
`protect END_PROTECTED
