`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+NhVxbTKoeYkZP91gh1PVj+brFpcehAnhJcCBC/d2CS6S1xssz1gl4h4q2LOC5H
am0vLTsgoL/YTNEk2tTTtlKBoECAzZvy2bSqwi8EO72Dnq+ZWgHKu4dqFT9I6Chd
k5ZfdOv9OkY2yhTnqUfQa2viEw4NiWAgWhuMx44RlitaOqIlIcoEf/LUqHfJ2NZX
aeO6fCDfSPjv+j7beLreBcVgwipmvLQ+vqwL/+pedG2wkzMH98E0T74X/V7JWr4u
MyzkEIg3i/u1tnwglGKVCLHWFU0pR/Z0eSv1O1ZNe7PeM3CGzxuDhK+wlrKVfaex
CfR1pxSzPmbhMOuSPwSvPMuTxcT4KSIFYv3Qto6ZVRKsJ0iybZFX9fC1bNCBIpJ8
`protect END_PROTECTED
