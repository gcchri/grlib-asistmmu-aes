`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C7Qe13aJqwI3YbSVJqydwqF2GOaO/iu63r0z2pQbUtlPLpVrmSiUgXdyO1u2M+H9
hO7ptvtCISO0xMXhPftrX/ojBJJjck+epB5PclspNTf7+uLPm7M+1aXh4mSmQWYa
nmwyToR5KXAONJUYjDsVYfEmRVHIeJ6PR8s0D9aZ0RhxLqys7qPjDlIW2Eopg8HM
qMaOIEvIhQNsooOiqjJy1dq8DMZQ5Ln1bdrhgMNu5W8XQFCN6N7U8Oxy5WobodFr
fOQiEdBZZgJUo/tiQSWaqVxqhqvy9lAvI9LpNBFRF17n2PN8wZRUV2IvdK4+jJxp
OYnoK7IsHyZHDLQfXR4zHHqNQWZf3nK8gkjGTqya/hz/Vw3wF8062IIJMXBzYWpn
/Skba4Zxi+ofiDb8tb0k29GPHiIi7Q+JJUiRPN9VSvB2Z4N7aFnac2bgNwFG9BB7
KvHobpwMTBgVFOQLjLPyLM4Tel8QxYnfJlFd6NT0Nl/t+lSArmYezBZ8szZaZ1+A
Rh1EeVb5h8uDP0jDKqDBcFJs1xd/5wmwx6Q4Cmg4oY0=
`protect END_PROTECTED
