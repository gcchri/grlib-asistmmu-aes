`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTzL6OEDh2YuWE7W89dxlfCqXLV++e8aj8AuZtAIrYCKgFsfxNNL8f+8YhLi3j8J
hxYW/8bJ4y5hlsr5/d+vX9wyZFpzg3ztjqZjJQue8dMcYlSCD5UVTGi3NRgdDaBs
FK7ygjscO4r/yDKsjdwA9LVHFmHupyhl5DcZCRTnbIjZuK06tCQ321lzxDPRyNh+
drI/DZB/YK9041YIq59aBL7ySNxBHtptRXYeK4RZe2s85/kLuzbVgyEoYhoPAmdk
++KQHvle38K/GNdkIEGeguAAKymLSrgUy8OpMa4L5/c=
`protect END_PROTECTED
