`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B2sC+zP9rLmpXkL6I/eSyAwZWSAOhDoTh0AOZqCkG8s6E9AAbZrU09rsPWe7DoGh
ZxNqUv3x03d8RRjba99/T/GRG2UQG4LMA6hFIlwbLyNZX25hNvyTBYhNOIVxJJo6
hZl97eZ1N+g0eb+XNxajG7dZS2aZlKjmWcrM8eawiuxaUyiWXeQc+HPF+izoOCQm
YSatw4l/Wj03SuEgtoUA0RTkB0FsvLldlbpQovpxFfjpPeVViRw1cQ64aCdgItvG
UN9lo7kpDi1hV2WMRqpdy9txUMDVbqKtsaADACXOpHgSJPD+RbE4Y2F9SSxD/1rP
PH2IJZoBSWEeJ2YHHI+iwQ0vofEWrAGXmtsSkY5Phm2WkbkWw76dOIzWeCGY9oNK
Gsn67og6JocuIt1yWLsEKCsxrERhOvsxs007itanWdiiRA/V576ZSX3LVZW1AZSo
ApQYC+W4L3pODiuNocekbkhi7gQL/P8wQktSHFepJOXNE65mtMdr77/OVux5XDkf
2mrJ50zh0ThWt+WQvncfbsnK5P6ajIbxU1Z9y916uueTmSmeNmLWqkVjZGtZTPkU
V4Qx8s4hchKdxJJSNoY6tA==
`protect END_PROTECTED
