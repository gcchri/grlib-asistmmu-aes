`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2w9+95SNyzsb/fe7o0CHa98t7VKARXCU8xmXy99LAZIGeTNCLyb78GMKUI8kDKh
zNfiOV4bgZYRLSFFNdP8lpyuNLlC/zIpQsQOlRMhiVsy5+fUfURspnC68dyqFL29
nBZK3mmSzuc6XXqO9heypf4GGdeXUUtF9Cn+S9wDG1Jid80NKnXOZIDTvzIgjaFs
R9ErK7saahrVchatH9fk2ojDgcBjUGagvQCNxPOb1jU9nkJ5jtJyrxyxVPJOzNyD
LKdqElMdh50lR0yrmf3EHRnIJ6NKBIvFdy+FjD9vzlLGw/KBWYRIgn4FRs25GOYg
qSNVG88DG2VtgF409CbhdDWYY34GoRG66jsqN1mkFgl29CXCUZi65efZYY1dKjMs
SkNUkC7CY6NWuYz90ElP8EcjFYyZo+ibATISB312sHkgA6RC+drYsIfjDJ9RS6n0
650QbZKdrP/lHfzL959ZKkeymJfqYPOgIuEfXONaXWzoF0rGgZItwkd/+UpeBdDc
2tR1UDpVPE3YMvWM2MFPj9Q1Hfo0h3KPh1AhY4T8GOn6H7DGDMRl9VOsTeCkxtmJ
ZqgQl3OFFAkA0R5PfsGJBAF0uCfvAGNouAsAuCAmXg797sI/BVgwTmBNuz4EDLW4
sdc5D5UNeKXu4IxPsbiQyXJe7/JaSmfqvPCqGKoJzo+Da1vy+PFe1Ic5secg/W6V
q4ZXx4csXhBThJH2aG3V/StgQ7caHu7FefBqSarRgwyoICu0z9TJaSrvCmQPwFDJ
hv1GJe+FV4Lri1h3gCoXMSN6Ms2pow95L3YtLhH+s6V6n3CQF76iLzj9IBajoFnK
mI2bYFQHzcHAPCk2HL/wcR6ee6K2Dtq6EUfcSisx6iftO06o4b7e0ieHz6gbwicX
IqQXB3TkRIqMBZV+I8XNyHnPVKg7UxymJ8Apv7kC/EY2wnrrEqpkQzykIW98Q+Ke
nkz8Rd+5nroszl6pVHULR4pDARB512moJViHCMA9e3/ZUNThVLuvz+EkoJAaF5H4
VKzVdBE3f3Gd2zAEO+36MXdaTXm+CaADpf78Mzk/OX7l4+MmhG5JwKojXxF0Fu8c
Xc2QrAX35wbhtSgtuX0t1lsqu0DbizwDH+Uhzt6K1ZRT6eYzXceoAq/VXBw5HIxK
01Szvo42MUobRR9ZQOheYBe3cWQF3HMrtDim+kYUtzsYQcGDDk7LQSvIbCWn8ULG
Sp8tmzPVROTuiEirNfnnhYx0HjrjOwbvU25npa2x8xI+zKRvmsMDPJTd4MIMQbJS
HCg2lqHt+YjyE4IsIUtPSWRBk1GDmbm8ekCCNIh8E4nWhygl354gp+1i19l9Y4Gn
EhP5wn9KNbe1gJ1r5nJCSauuCp+rzsPkEzBoOshTVaNNPwymlUlYCsLEgqenhZaw
ekCPD0YGmqqIldhUPypQmxgAqHatEFb3xNXaiKHFJDaIu0rT2/12t0TpJqgaC+oT
2UQFn8O4v+mmxsw8E1F3PoiEpG24bC7xXQBo7ZYKVntJvZX8/l7JZacG7BGkeHu2
mD7brzIf1kaxLJ4+UnmUdXEt9aDzXi7COaE7Xhcw/qbntqlfnglWkucT0s9ld54m
cByDDCnMqaYxuCnAWWvhQVgRXwTduRl7h4EYwjz7PO8it2VelV9Nqok9qgWqWyTh
+EoXbClPRsy4hU0Xh5WW65kHq2P6umVrD3dZm4xe7Wsf/tWj+sHtBHrOV/TSOlKA
sGIrEcmwsAGO5w10o9XMH1Bmen4/JkFWT0L8QEZHbZcvGXMa3XG+9/5wDUGWt9nL
7vG8gwdkaD4df7ue+LeOGle1bHGxLpEmgUXyQlFu6cyksx6cyNyVB2zhkOL9rZjw
ybZrDf5Aionut7ZU7R1w2llPzGbKl8Xb+Pu5urHoiWyfpiMt6qkzWJ1A73i6JUsX
bnpq7214Zkr0rh6YDmILK7iv9joHqCpoOCLMfjZRM9vVX9gdiRpcxylnO3UpiiUn
Ec4QGv4t4XlOZytwur7v/jw9SfR/sGF8ber6+szhO3ESybr1VBER0a/TyYv0bBar
FDqHIcufMj65ZAxWi/nkRtIsgkzU7jSp5cUPZIEKjeSNoUeSA62Y3vE/eH58hA2+
dJym2QzircIjfaaH/okeWDJv+AnaPaunmX1nXLgCnrAC5vNMfqC5n9yGLLLSkOVi
AJpdEJDMD9lks7Sf9/VnB9go588d8o2JxzbOjCh/p7kG7fEltEe6Rrs5RSsw7Zj9
0FOW5jjCYR1RBYk8b8N07YwKW7U7gVS8JDqg4c747uh+u/JSn8+F5ukE0Znp1PYt
E83gy55Ul+KtO6qilbzjhBaX65M1Bs9/juqjABm74DYyiuL8fHb+htWGz+grMj/G
8yUf8iKEx5aWwEZB/+di594rPnPhvp1U5XC6u/PaMpdqe2WhF70Ee0BPqaiGAhPX
IqaWWTxPX+WUPmSPCj20coFyct/xVO1nnht8M/zziAPnewjvtIVpgZiFpKW0Yk1W
RY097pr0qOAjYF8OvveZn15BR4WNiq4Mmo5QR7yfv41L7LwcZSdtrO3elSkyjW75
v8S+XQeoe4MtImBSydCLABqwPtBvoVZoipk37CBTGrBN4SgrY/61/b0CmTh1AUNO
lsZGwZAQRRPshBB3EqezDytsiAyc8cDodBD+p/OARPNXGB3SeI/VzrvBeniI5DLR
X8/+NeUABCLpDYAQJjpD7APrB3UspOJT7nffCbcDbfdv7TNCuKWEzITNXqSY7FCt
PbAP2yZcrEx/cOvQHcbXHa+sUhmx5OD3jDopXazbuZ6/Sv4zqU1VYfGsngQ4+ehT
i2Q8U/7AwG0aFH086F1unsE7Q9c+g65SS6cue8TrwV41kYXqkaEgl0mMua5Q317G
WhJMUqEzGMsowSjDGiyOd3Lpxg9PVbCaySMQPTK+5Wh8aHchxosC/OfuZFr8dfY4
VejmugnlXXz2TvuSG+LUaue/EjxSKHRRSkDaCQqSdkMiQ6F3lIiY/Lur11OYR9MU
v+YQ96lj8yys5VP2VpYIeJNTClxokQu2ZGn8oLdh0XAYYsNLDbgeKUMPh6F1tHZZ
RU4VtzYq1TdEqqUBHVimgkgmXZufihg/AgXNCGXgepS28kpVuXjvv8FcyIxOIOWU
mqX2EfNh2+154X0aAWOdsiFQyaOkAMoTUeF48pLqpQz/h0tr8qCbAcOROBVecVsL
IzDbX1VoKvAw2CpHmkMw7MvL16Z25j0k+7HsoqTYTer9/xALCabIsS5xXMHxoKzc
i37tuH/3uHPSQ1XG3ZVa1X1MgGZmvrYuGDGIOh/cX+8n51t8+1N0TrcbHYQf7mBC
LlIXuQU7IlVDW4H2OcqGNhO36I2wuQOSisS5P7FiKcFiG2G48XV46TnzpJTz/cdc
81sqWAD0V7kmGfdiGdfYiug1FQA2YyI5bVr6liqnCE7/pYIMisAnS3wRPp4MtaOO
MbKQ81eY25oY34nM6HxbY/43jxnWSwqNJMCiilK3MwFseGT4wo8W9yHfOyXHR+MC
RShmXlJoPfa+E1wN+0AV/UIPy6VyZDx2z07pACe+U8sLwoRJwbcMnctC2Y9KuT/T
JZGfIuzfOfQHx6YsIx5f7hHK3fQ+o7iKRGgobsy8wiysK5eL1w9NSS6x8si4NMhr
NneuHGVnhODkT5wdBx80ZhhFimCcpkB1dtqK7r+9ZpunNQSvLyhASQs5zxbVzyn8
IizAJBYTANDiJcZNg6MZR1DC2yGezVpzTCCld2h8+GIHgPrczw84QISbT5JDmxWI
wjc736P2sadP3AJj9e/bBdPXQHdF/TzvBMRdCVN8x6wSgYSNjFhA2tziksg54bR8
Jb5x1eRYGRCMXTWNQyn5VVXEe1/feaPRcwQ5cJIOAYWw5txQFvJccQOwy07bVIyz
3+/nlr6DL1frsx7C6AaTBvpa2dTywsShw/6s+mHfHIairhjYV8ANpztkXTEh9KKH
Q2CC1RXcAkhoCbeoWdE2We9Hz4xsXuQCX9I7Mk5BcplyqCoAA51R1ncBIRzD5vGo
pwneJexphXMy8GMZq0VF9iUy2QwXCRIj2IsvbltarFJQ6t8lqUEvyQmLQEWTyCJo
DEG9ZTTefdjdRtO/WMNKmIYpzCkgEoWKS79hGzCX8DwmEhyjNN1k2+rdo9lPSeBP
PqDnwV7BysQgvf2EQiaawiz6ZMyPCdWScvFMvX2f5aJX7JOAlW8Lf5sdXEXPNXnY
PzC8Owtu/3lfEcJASjr1EyQ4e51yLL8F5wEx1grVauUunExZb0p+mX2pyQvXyQCS
H6ctE9FXBpsQBVVCZ7AEMxNS8EDYO3XGLjRiTSfPIy6nUQbEZaWqzuI7JgCmVI8l
7bcdJgx3v3F5+yw/s6a/F2fZbXhlKStUVPzeEW6rHl0rAumMI+uwGBCNLCnrFjeg
UhsQm/2s6cqPEXErkTT5mZh54Q/i11AKzZkWJ7JfV8qJ0OnTJNMuAaT9VmejQt4T
UQ+bTOelaKvYj7OsGuXNfF7dqbVwOIzgseCIUlnpraZoswkxqiOQGUiJwg7KWgfX
OZp0nO0GXnFUD7OFBNn6LhZJMq9mp3XVI0dhOw8JzhbVyeYAfWcuK6P8OIJi5xT7
sZIqhd/HEPi2gTQnWfpC4h8s/3Uo60G3vpk1iPwrko8Dt7WayMzMqBeLLxtlIu50
3rQ/BuJVnPUwpZbzAk+pD70HTYU8JpbGCHY8AOzWa7QmXT20jtfcGKHpaS/mvTm/
yb8IYdaFwg+XhlQblLOcDMC/KCzv0NSkkXekriTw6P1mJKgbk/SyweC3nUbx1SmB
uUrGszt+YITP2Ce5xuaG+ZSEAXFdebTmMod76EFYEJU9rmIcmAXLvWCD6JFsvtEu
mhlp/efT5N1lnBOzOhjcd+/3mAuVXmhWGFYk1/7Wm3VtDeEYRxq21JXpb2tbcR+6
tZZMfl3yClmHBWvXVMxq+V2WEFvueB0ves85Q4LKNBK1ba/+S+sN39Xjk+msR6Wn
hzWtHv6NNTMvkfCnsaNMGF5wxFTY+R+gRBF8M1FHtX5R4LcY40O4ucoEdwBSJV/D
1BdNObucT+WjAuJanld5HaS+Ct6QufbTPKBBlkTGsVImmtu0wjMfovqE4s+kFa0i
gyKkRUmyupXz1e/hY2RNT+GEClAmn5dH15QBbaxG+m2tnOFQrM2GZgEHJhfWgksu
AG9kLr4z1W0KbDOHAmWrW9vgByjY7901+0nLwNumPF3C55vX0fO4PpwCDaZrT4Zb
j1btoSHDht4MZaFhX4wL/9B/1n+Il4crErFh/RqjZTqU2yEjHFv8IpYmNgAc/qAB
pHZbCxSBG1jH2W+13Sg2+JY28IyOLSXVvFM3D66nEanvXN3w7twomkbRkLP8yMyE
QGvMPbyYgpPBRJMrXbpzgjZjAqrr1B6anN4ZEVfa8331xDZLxJyLxoUfYwmTKL6z
PmpVHJHMBhQmMUoefcz4GsLzf/jhu1PADRSRV12wzm3eWsK4NFbrAj2UlS4YNB+K
cBlOwHYaq5qOEqxWiopSWjUljMhoT1XwIiSredatVrmKzsi/X82Ih+aUUsx8upxx
ciTGUznx/+dQiwe2ZFXgjMBw6wN9FF6i/xEFArtxy9OcxAtFmXBo+YxENhXCjyzP
yuAipx1yzzsjsodXjpcJHazOZEbO6mSBKZrgLJ75FM8z2qy5XOi5rDo1typ32Koi
7Li9+GWz5VLm2O2jrqz1KLNOEbWeYAtvLupGvyaN83otHrf1FWER15auUAH4z+tD
uob4HWJN4LZnjJOG539s5OzcLmFd5v/KlcQ+J73UPlRepyVgCDUvLEXaGRpKLobw
EccrFZzG2I3ihgZqPhe8nB/Xryg6U0BL7Yn1Xt7RDwqlxEhSyXlyo3ypcKbnkb/A
ng5gT6RQyqCuBgiJPDIqfe5dxOJsTpm9qJYQZ5Q0pjbjDcyk0LJLIO50VqgpS3GN
HOazvujNApcpo8dY83f66FilZ2dcj4UfuJDHALqVPp2WzAGSYuJVDoL7+cJH4JV5
gdgsyv7aIIA3OpNjpt3N9XcBFnS5JHeVFbCCt2UoROSpkREWDxm/KWzmdlk6oZJB
o/cPBbeyXoE24tAMdWmYdNoNN1NPlOh2JJfHeAnV4HfNRYPgG7DvkQieDu+4mK8V
MvfuL+O7xFMR80SEwZdm/kLQ4Jjb+eS9kzi9FhJUIYQqfAG4kQG5t3yzPgCYfAW9
I0azgjh1YUYGi4ucPouF4vuEExGZg2OvylsF8hOJoJ3acmZnqccbGA5yKRYlmyNb
g+jotcPqLv9yOvH3CgYzLAe3oiCnCY98jm6wivNdF4PhX1XP5ZSUIg0AtxTOYJW6
YOMAhqDMr0RfTLz3d858fotGlZ2JM32QBEe7oZz3nW+bPXjYKb5GQsUTAwcDtMaZ
I9GiQhz8Gj6AThzsXBMGk3EQ3gyuF6hHVj35thXEh9bZGf5gBi/tCNeidohjPS2J
Rn5xPqWOGbYf8/FNeS5xwsFBLPyHmwBC6/6fUmqp+cFg9+53nBJD0L7dPe+GOAiM
qnAvRLzMNdDuSQsHIr/84lfK1FFRD+PkWJf66gavaEWIVC2m8RMxfC6fIcr2AfJP
jbV+3zYQlw46GCb0Z100oMGv9hu7xxY3VGI0CnThb+ys4zNEr1FpoEY+/Qjjcspr
6GTT8FA+adKIUFg+a8r799SU5JK4auIfiszZi1K1cXtBTgYr8m1n08EpsZoDSlJ0
N461TQCJO6K+uLXyRAKks7pMg2+aJxuryFsMnvtNC5Zg4Hcsd37saVPOMOmD1uJo
pTsiElEeMZKyqSSUP9N68aQ3uBRLIUoH4u1mRMUxiJpTGcoPAHW5QuNytzTQMsCA
N2f4kA5b84b95BuoUedorPVx7dv0FFQwRbr36DcfnL4ATStX3TyME3wvl4VfxxD+
kCkCusAHSYsewIMpUHUxG3fpqlMH2D4Ilxowg8DG4GoA29evUJOYBoHEztBgnE0h
5VsLG7uJt9wtghdl/fZ5neLQbRq4lebC12gWK+a33HIqZBs4ZVhC+/vSJJsTNPot
BQPG6JZKd4ruR5fZW5JgFq+Crhf+PWl4cdAqRZ2tDPt9X05n8GMCtGsYA3etFQwz
fZtlwJMRCgXiBfDqIZeAB2BATRzYj/Z2tTJV40YUjqEXzmp1wWtIH+Of6L4iAjt8
aV8lJQYv84meF/nomjYQnes3Lq/3nUkClcLdwcA8nqnhA30AHqCJFywmHMtmdphu
8w3Vt10ORU5HFoRaT7Dr718hArwJf9VJMMhcU2YCgRlN358gwD3hgQcMaoLentjn
B5OceeABBH/M9GVPsyNLCNzDnRq9NJrtGcM+CajKuCIqLxMoI2MbL2aDbimp2Kzr
Lbqox4/9e0DfJMfM9rZWcbZ8aZ0XxEG2jTMhi4/myTdz5ZpgAvn/q0nhdNyqyNpo
NlJD8+Ch1SghGEZANI6151v2YsckaMj+uyVgtIC9rxhL4V9MpTTF975gZa6H1+DD
OiRI3UPkEXclIb1vNBc8kvt8wXw4GyFtYSWXABZm0kO1+4vhM3CeKVv2PyGuy7Jn
RklFN1xoihGvldMg28oLH/KDPyzZtXupfmhvgVnCmR9tmcDjCaLBTwYPGzD/sUt5
UGJ8jMnNVAnDnKea/ZFeZ84Zei0qRyHK6z2pEHf0A1zZlLRHxQnNVGHUc5zv9QTZ
aPaOZHvQxInPWKv7QooZBTySJhcPAJfiSoh4q13fQ8DD6Y3xFsUvX8rye4GGpPz6
xzb6+Fw5LTCkb04htWmrLA29B3esTwRGrEoA2cq+jy032pbiqfdvFZoyFNsPOxgC
vMrNpuDd3bJLtcWkaLGfEu+qFXaNulJu85GVgQKmn9b/x/20UN2EcVvbHW11+eFm
hTlvHMV7IY6+8RXGLlEmXCPbhJNfI+eFXwPL7kGL+pysF5gIYA35U8leacNwufr4
nl5qs68ewz1zlAudK/qays2cbSMulpVFDVK11dWTcFK7/UCkdbVrQLDpE91oo0ho
znXL2xmS250Mn3Yh7d4aHsEzqm6zS8jm1h5XotYqYCmJyTPvrigkbiT0utj8dJdM
I7BPFGdPizuBT2okEnvoKmm0yklSIQeF44Ll1eaJo0cvk/VyE+ilQH/hcFijOmtr
V+r5Um5pAGbfGZ+Fx9U0dQWV2nYBdxKS/aSth3r9ZKL4Wuqo9iJgIADtD8YbdjOd
MEworGqezyxxMGgl6/UIA1WjJT0e6iTYZJRZc0VPkjFMwXRbz3XsrK3vfxx9oz+3
uo9dY/7c6BrIzujwp1AqJME5uX5nctFZ/HcnNMRQspIt+Sb5P9gqz71QkEm90AMq
eK0DEoORFzmqT/5UtAYfbLSTkI4Ay33gj0M1m6PA+qMKUaKBrEidD21FFguAdtgb
6xLEgK5BszJsurRoAnPLRd3Wj+v07fZxl5AV5T9QXnq9tp/6j+tAKyL8EXhuUYvc
UliGsJUE8CkRTurPdCcYIUTR6pnV9uLM72cNVYgt3l3uVjlDB8kpow5iB7ZCJ7E4
tYRgdLou9ERIP3s4TKAJo+Be0rZECvUO4Qku8NXurbTg0bSxqUYPtqYDnSUeSr/b
yeAmaf72PreFxCxB7HYqrUY88jgs/SxoHN/gHT1w16rYlCa9P3tUy2J6wT/htV50
luQjSvn6fnnYVdFAY20yHHGxEITbsWFhtwXk1WhK16Plx/Uu0Gxide/BWRbC9j6+
EfpKFg7BJVu/BdatuWJwcVOfHks+QY+iWcUlHomL7e/CSP2KJoXbKHXF7OwJw9nw
/1sfqNcaO7yk5nqUwUzEr7Tk6shmV6Q4IWsahngQE91G6zbJSkB7jNwpAQOI9yRu
jqFbEikNaqMzApQBvBLl9ANSyD6W0bSSDRNmamovU2DrfOFv/16zDMm3utORIEFZ
xrfr+A1now9hv4NIYSBDtwH/mzFgsccQsaDvS5BosLyMcPARqonW8G22mKIJv9Vx
6pkPpUbHmp/kvj4bFdYd0hSVN+6R7rVzBpgBYqQVAux/xd3d3LT9RNnifAmfipDx
qurnuh3Fbaago9hFmo6Du1/DecPLyO7NbJDgo2ROyZaRCzDGNulZTpUmNbMw9umX
7R9MpM/B4U1Mkw0x9vkiU1oDseigLSNZHFz+YtX9Ug1jcMTITbniO1DSIeWmbYTr
03IquA/T7BEdR8lGB0Y0b//v0D9STtCnUF/pPzl7trAmTxPYE8oTBnFaSzrq1aGr
/FFoah7c8YkPEGuc2jOkxCc6henFzLxffsQ/PX8EpYiRh0JnHkHIV/yKJrYSrACV
2ZcUil+mjGQd7M5aF9XewQOcWGQCs4oKkn7Lu5Z+hWNb/8o6qwXmLKxykmCAtbYt
AhQ7VRshTUyBWtt/dce4ku5yugcpbpp1bw2tuYGMLJSdZq+Ktt4Xrajk49aG4iOK
F1ab4Nlx9xav86c1yobqOtkErX3859/7xx6yr9uQoOX/TiGALEXCvtT1OmxPpX4z
cykxcjpKHyJPYU2mf9kjQqtgrP5HCxzTKUJ+mcYPNyGh/LMizpH0bLB/MRFndlZO
Rz9E2/0e/xAIj5ymtY/PPgEb/9rziZvyKe3/Y2pmqJcbq1u2fs4XV4WqfnzxXBLI
lS9mrLQMb4P1XK/uBhCUQ41pYmh6myqRoRWn5CoYxA9L849B4+v3BBXP8B9dsVDk
hJvUba7jBcq3G0ExOOfswC3id5ecypoGvU/JheXuAWZP20YQGnOz5pDCcPVu7qeG
6d2z4NgzZcVwYXTxSKWDNvdFMZJDn6kK0E06FiWGfenpxbGqqOcF0smCvef4Q1Yr
b7MyfXrZl9jHf4VEnOJkF++3raH3g7NdzRxo++vMJkTU6KnUuDXfq6f0cYHC2SjQ
GQtr38oXb/haifJF4ig3/+7fPGa6tJrCYRt6sPj+DKp0sV09ksOssvH7Wpq6WTFH
mhUD/NIKnDdo3AYi3tGWRjMxESX8MXMxFVwOEzonsKnK2ApI5hRSmxJfcbgWoFpT
sKRJ75nAw2+UopL3XqYJjOHUqu5mkHFu2hz8gGljH2AiUP9U43fOUQbZDGCVofQl
qxTmnlzF4Zl7b2LpEN+N8VuS4t9CGEb0HESXvhMyLWrqJQ6cnewvwPHlu3OzqlED
rlmS0mpVON5iDSK1ebMvSQChz8Tap54OoVdwggS5CFyfgilHbkGB9JpC9B24Kl5O
RME6CYAHc9RLK10UNHK65OofqLy9QhqPxh23FtqmK3tstmwg3q7Vtt1r1ZYafLaJ
Q3K2i60Un0TtN0SSavqMKIWAsNaImB/DBp7ThySB/gg1ma5THSX9TkC4pbYvGedd
s6MCjOdIme9iPNNjcjfdv4JYIggDljRTnROSHSCsl6o=
`protect END_PROTECTED
