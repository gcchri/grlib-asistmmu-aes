`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GpbiYoqu6sk3B2i7q8oQD7rGPWfFReA4dlsx3tTm92pEnTHvEk547T6FLYzYGVhE
+dSo/k+Oulw22SggdbJFmTOAoaDqOki49CdnXCjT7hxJ86B2vdN+cz5e1X82FvTN
9E/2lyMziqNUziyqL1LQCelSNvAI+nUAzszbJjjVmFrCnlJTHCs5GcZ6yssus9FC
Am9xCo1wG4LyhitNxU4BTJ0CO+8rehyDL64WT+q6tWAUDxtDsp8ELkisQ7/WENv3
GtKThSv3YW6o607jF0RuCknMR6bewJDHKBvudQQZAnBATXmSOp30nunLG6Yd0TBa
RdKs/9OZNHkRfOa1RYXQO0mqai8CkmmCDBgGnPqfXLAqzvCXumh60N2whbrHolZ5
DSbpoo9fR+UJNe3S307jk+nw95lA0vxG68VypADlB6XLJ//xzGdWGb8AVQ86tbiQ
CylbALFxlt7nhd1bOyytWq7nnp6H/OMlaTTWnIpTNTrTCX5ZVryU948vWrySZVMq
ft/EO5E+LjZaGnVsPX3wIQ==
`protect END_PROTECTED
