`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x90Touk8dkkDy0mdMoWlypQp9zXJj3+9iANyfJ+007O4+YIa/6RNCeGDvoXWFftB
4Qo9+Vg7qj/ctx44LETvAdIByV2AGBpByljOVNIzrjun23h/dYpcF1oRZOFZ1iEh
N+N+lZEbYVFgJq4YpYlAC1G0SPc9mY9PuoBcAca3+Lae7mAhb+WqkOpXdmgF7K1t
1mKyR+t8fMQVtQbMRJ5HvWvNdEnoyuciD9xQJkLCZj6nPVh5EeNiR+s78pgop3by
xpsNn0lBbiKFSNmoe/DuOe5pJbD5gpfOODgerGVrCRkM2WxHkkgX83/UzsN/02+S
JbrpL3aL0ObjC+ciKw6D+uCQhKOMUZoK1+8qYxg/y59a0JzGze8RN7hyRIiJwH5C
YiIpY7mPO0XZs4ilqwV3t6dUsJ/iVuLx6yKgmDfSHGedwXwyirrpn0W/ESGbJZdC
LNuR8UWcCmJnvoH1+uNIm7a/CX0iUn2r7JtMUogGqBcwA13esknwi77q5GvsijJm
/FrWCXb+SAh3pnbY4ZJ6EpU9pYXMHexWiNq/olxXMS6VeTMbUEnMntqwtaK3JO78
PxJ77igwBP+ukhPZ/4MrMMWgrcJoG82UEGbx78DYb+d5GjWfr+oHyycnhxmwkAAM
9PDo3e9vC5baW/GRqNuu0Q7sCior/W1NAWxD5cdodaqIT5FuFHLyvpkK5Cxf/yEk
QEModwi2SQGqRbtRG+9DCRRqWY77DNb6zqRB3AJ5780o0V+4bsGTzQdWLU5qJEZz
cWTgF7Uq+8aNcxbBGDypdahO9M+sQbjaZ0EZAuLM204EMVyd8lVSftf9wZ9SzyMl
ULpB/mPERjr58ekJl34HtL1/oWqMR2hliFNJb7WRBWD6E7rs9WTPDREbeic28s67
odRUDuun3BkRydFVmTv3Yb1z30NazBgXZNM3ab96TsYm8Z9wXfH78lj93Mx11qv/
/Ybd5Qf5VAjfzM//9ncNOizGSGRDYCyqKMBTMgow3jdjVk9TjidbIhUUIq3l0ek4
Ns3w0P2fGKK6DUyloCabsMYxl1gVegZXeFMQpDZpUy4=
`protect END_PROTECTED
