`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TK4VkWYc40czMcUUxIrpw7HAopGu/tGrhY6bB61pCpR99pqOAL8Js0OWQUvBWKII
CUQaKoIAN41BtTPFHrwaLb2ypRbviCJuveZCOp0Q/DKrEryViph3BauD0kjfzavi
padlXrJdLCChIUfFsOOaKamTVAiPtIUIj2raq/f9H6dRC8M1XL3qpSJz7fOJ5+Hl
rT/PztIzzNdUtpVRgWqLCcKDqb2D2u2oBy21n2dRCE6wPqvfOTbhU2m8nCjLGhQN
ZdtyHbwShos+Aq0Lm3M+HkD0prTeKFw8fVS35Qy2N+2rz9SK+k7CFwJ8w2rZYi36
7y0qZg8teJr7hXI9pgaQ4dUawS7LENEeL7Zf964H8PWi5R7lM1D23zNw2EkCdQJP
aSMKmM1sRahVWO1wzO6sQfNRpwcr13EKPFD/Zy6LN2cYH98w67FUVDIBStlZ1PKm
wgB7CajdiUQDJwSWv+Z6qJhpsLKr90vuDm/pD+m8UcI=
`protect END_PROTECTED
