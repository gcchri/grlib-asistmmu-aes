`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wh3eH+UHdYEeiamt89gcNzqdzpEClFwOWPSQHvQtkxNL0s8h1Yd57B/co5DUndmA
VUmcb0To0ePlWBYEo+ewoQGH3wj8epo3OtO/6r/w7A22QXVdqF6qTMylG73UQbKX
cqL2EvBqrtdqQScNZR0OUm1iwN4+LCNE/OxQUcX4+wUa1VscCMbVktvV2XaW7vnu
hUaUbnZnII6kVjg+gtvPZGh0tCdYEdv1n+/WE99vz3bUaWa80vgHUl+Xq6bCl1HJ
Sw+NYRFmC95p99QO2cLkHFuRS7qKQoCeBqZspPSPr2CslHdqwIAJJJlA5/uNBZm6
PSIQtV1ZFnf26IuqtQctjAZ38wGD0vhE7oUe0t8R5aJJVAorEYnfcuvKPztlYiv8
TLdwTY8YCAhWi6exzoEGKtd9ZofhtyvBeJtorjo5cte+a9Zrd/2vOPMbhjAerMU2
xPEBd38JakpsdkcOKv1VddorfE75169BM+mmee/Cz58=
`protect END_PROTECTED
