`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9N+RalF18eDjuFXaJTBYmhsUm/oomcbhIo9dIu1wDKOfwdyBLn/oCOtNuCe5Ufq
/ELYdG3Gre3lcluD/DwkZrbSpOiNhbU50QZNduXhNUXfXrBLG92lAYPiL18YrmUy
DLdv9e3Aj39dyGTts+Xg+x98n8Z/ejGXVbInBf054pZWSH8BoG+PLFfdCYooSIac
I1QWoTUfzu4NzmXhXTlexytYWWtt4FHOn1tLLbPV86nag3ylzxwKUBBNNoyKnkWS
S5NZ4oAj2+i7uJXT83DpU9EMtGCXrLk43u5+u2jSXWMRyVjtjRo4kFj8Jpwh6NeS
okqK/V1KiFv2NjywTjRi7m0Wgi/CsRdTxaWAGH97ZULQqk0rlAhiYhbIOfRjKEJs
Tjeh6UMER8EMnRk7AHKDZdr9V3zYWfffeyZypMFoQG2ZHCeEsycillDdLDbPMGTD
drCZK03YZkf/0hU59lwkCv81oLQhL6E35nZwrThHUgV2M5P/zQdKEwBnWftHe7gV
hef6kwo9zQz5DNVBdWzVt8B6LLTQ6cs+pva55ucNXl0QbWRepaKZg7UUTOVFZbMo
ltMad38dd9syhv8HUD1JQuwpyCVBv7R6zRw+O+6Yax1txvfVuI1us2dfgzo/6UHn
uhBOmIM8fxwDc69oO+Ta8qtZS4M21oMqQM6jPihT2Jk=
`protect END_PROTECTED
