`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oKFlcCV6jR/NenDKdcVPuhcBxYifNq5jCFezz3uF5h+LGZlbab2BseyeKUdC5kbs
eCyuNIRlVJXPrzQ8qr9aXInPo1o9NHVnYPv1K8pge/eryfA46vyvE+U8u6sQiM3X
613/4djbp6i0Lm2b5685YJn6nY8zi2v01WLi1l1eMjPvjp35W89irGOk72cVkkwy
MF/DQXb4znbet3P5OGkKkL8I3rShsA7ATCCSo1fP/ec3loA39yMnk+GLdJJlmbzd
GlenVWAek8DIBIdzDIbqo0h8vgFkRfPw74t3dgMlMwVpunvH30m5mpQ/seRmFjfx
qgIdkKPDiOG8s1i6AqrnQho5GgGdJ1wbh8wkLBhvIg/c0cNxdrqmWho8L6I3pM47
7FF3CQIpCb1n1+aV8qjiou4z5rbinGKao5tN2UAX2bP2L0/ZRVGBwj8lk1NSkep1
y0fa1Bpibp8hHYqJ8Liw5eYSxrtB+nD2l8Du72v5u0NxMv7kJJ0kxsEHQwLbdwvY
`protect END_PROTECTED
