`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4tE2c0qYsl8k8E6zXmAlAXqpKlWCxcV6U97x5uE3O6M4HTasNJte7rRTVKQLs1C
o/s20WN4VeS7i+1KvLdXWWwFUs80gI9M5oNjUIlpGZhdWT0PdkNbRa30BxmSJKEx
Lt5Frd5LGhFBFhwHt+djoFZ+1NJw+fkzAU7gKLgZAIBoneQDWNaN17WoBrYFFVWb
8mWasDq5gNDVJaNdPq92ovYnmxRligpTTvcH5JU2H34ZP7u37PPNaonPLnM13Bse
zrLtP4Zo/NtMfjdOn7bZzBhBSM3/YtHSZaPaRABK9t0hxriMHWPBRTk4cgmewUEm
+7ODnm/0lGs13VUt3K9Jlzr5HVqEIL8kB9JaOzq7fGJm5f19zELtTI7OBcycrOnF
hhx1rq2PB7902xpZB5HykA==
`protect END_PROTECTED
