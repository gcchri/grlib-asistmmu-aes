`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vv8hprqsiM6lXskiUNZ9ldMKHNI/3FdPlSE4TgAWUwFsrpYH446+HpuZgRQR3+jI
0Zo2FMp5J7Ct1fUvjSNwrcbIw3J9prMZEaxzOY6C/O4F8cjh+dXZOn8rMvR2F4fV
wfZGLEiTAtjg9X3ha29m7Yfb1xYtLwZNdlZaXszA1BqQaLKUZ+urXCESU2dfLRZx
1FRcs9Y3nFFCy62ywr7mrn5P5nEc9U7pyflmjweVFqkNFHmp7zVREmGMcwInX5T1
+3CKZOL2PgobyhRVM383a8j4ZxatMIhmGcp5rS4aCL73STMN8FnrvNMH2Iv3kHi0
zfLNHeV8r6kpRXYgZo0J7GTAb+ILL5kpGx/OdGTFF58xIC/6K9tqGZf/jiufdcVd
aLFNZbkaPnOqcBcyro1vEnHHUUFmhDj+Y9XhwDCANyo=
`protect END_PROTECTED
