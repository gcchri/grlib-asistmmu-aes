`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gko5W4ZyUDjUAxFUdyTkWCQrPg58UrVjsr0N6QKSoi5xIm4GaqiLWgbPMjPevWQv
engQrSvAQ6mInlbECbdgxkeByw6q4ih9kJdTx0ZRG8j81bKi8oy0yt/U+ivWyn+7
xGr9GU+4U2FkTAP+g4/znQOWI8rC7H/GXJGRqfcratAc8REqsHNHf9+wOHX1vOFH
WUPFePlw7OdAaO14Al7THLL9daBwo2rwVJv+5/dp37g81Bdy6tgssvVhWnSbt06d
GTZr/9MnVPrirS8/5inptiIU22yd4pQ3DKQVngbvjZFdzQoVXnpt1wqDAOkbbrNQ
KbtUMIlMG9SbfLZg1VrtTj0qbLEnpPF2LHzPGxLlI5zpCp58MR9FDT3dYrzQJEiG
garb87twaKAdxB9G4pUW2gnE6p5DBiOHJ8hCMGyNN9K4CJwf8q52tExU1fSIYrKa
pQd2TDSfy3HWaaXQpLkljRp296V1PLRvvY9OhWS2JMr6se+9ANa4Tupk5yZnU4zO
vsmBhiVxdnKfO2xXPoZ+k4EVAXvjN4xxqmzT0h6T9yhdGsgHXrxbRjAj81qHB6LL
h/4mVgzBv8IdKacZbacoHoArdCHpSZ0OKO4kRtmKBpew/LODcPNIOra3vLl9dALr
G2BXVK2O45XmSLGr9opbkM4lYPHs7Q+RnRGdHiaXC+6x4EfNtWy9WmoOYajSYeEN
aJNy5y9bpyJYQyrXrBUz5y6bFGLL0g3gYxG/Scl9rJdpmpt1iIUdNeFQHYLvJGJP
WO9LycU1EVTSF+rFwStZJKvBvxrsegUbUuyGY7IV+OueEpP7Z6L6HHPABduHtdrF
n7RtBXLcPKJwS1hYk2xhizPEUKOBht4B+QitmQUadYRkk9HJU3ti649rRUpXTu5B
N1KaHVyQbjG2/xa+CqU437Atx2JOODMLXeraA3D6J2GHIq7IR9t2qQPyUbCNUlVx
Age6VgCcSLdmYOXfWsQvQyLIBFapc7ynz7wnFcZW3MaOqxvMTvIWyOqdYh1MIhBY
3+XPXSlkjvXs3wg5T/bRttnzZsYcvqqMRk7xRhqmvb4Rk5ptdVVfAmrtVZdx2anu
KjyIxCbGiXvwqxVjHNDBI8+lfwJQYC/hSPp8ikza8smKXdRutCn1h6CHsC5x0a3O
MHueXNDKBEwBAPM5QK0zgRdCIJxRGC/gehvk0fv4hnojX2qAKMf74NyrSCy+Vz4I
/Ql42swpOp8EE/BevTxsGzkhnuBYVwPuytcu9E2SKe7Ake4tGhlltl6S06di9NW5
iwepLlu4ZmouyjzKiPMe5odokSvX7PUDiwFpfqnIig8vkD2Vo12XsOtp096tbBAY
kh14FkF33BSuJJl2fPGp9YJgzmNMVUpu1fe7UedJgl1SmTMCAjS8ZnhSXfyHmXDp
PUWSXujZsTY8f/rybfFWQI5qSO2yFkg8LpeZWwB+favzCQM8pO3phr+6draFAmqw
tOJ1V6OT0aobtknnFEsXRAYYeXGLmEhdMGGYXAz8LNAMPZJCWPoAEFm+jJ1MC2Ep
hhqfh6XwfTauOIS2szOHIQOGaYwM2jZldeHm9B/LYahdqhkEO3vXm2e86PyDDD7A
vJsXeViAOuCCqh1FjZLxZ4iI7byvL6rYrmt+cdQgrZvvo/lAuutXnxXs9TZqGUex
tZHI2oMNzFQaPGNkwS8O4Dg2Ct7gD0L0KiMzpOIr7wX+8q36kcdYCpr8mfiuIyFR
67LbhVhW9JPpNUgXCCt+kjfEr8ZFsJ/UKFzX3OSX25qx6wQR4QMBKCgW6Nmp8P7u
VzrOhvt+l8LFQ7amjyDCiozYikywIdgAEB68pTIRjq/nlq/69/sX5VOLWE/mYlwk
EomuMFTBIYd+t3kASKEPxQShD3LPeRPgumoHT+UW2mnM9uSn5rnzFAslB3LrXWQR
rAWaS+P7bnXE5hw8zdBPKPaXCKDbZkBKj3cKd86wIVklsmLLFv96bBp36hG/GojA
Ste+oJUZhFxBPk3FtURogfkp6s39+x3NPCzdgzJKumZJqzKR3eOxi9P8gsW1xcHX
BoSvl2pgfrBHhkw5CrPuSWv1nvsMZa/+jqbIfTEdELDN0z6A/sCnj5yix9YMU1oC
53p88ss+KixSSFuiU2gKT2ydKknhNsHdEguMUa2zFvWPKLcS4/7R86PA9N6cedkB
JWIPRWx1tpslJbXqPay1d/dBKkoNNqORlQOTq13nD5Nz/V0NG5CpgUjM6LAeXfUo
enbwf66+az6z8j0ckh95syOP5MS2Q6yhGhEJbY83siaKQOtnl2s8eVAM+drDSHGQ
tyjATQcT3+kUlrwjxB5X0qLX6xnlNPMIsTEkC/KqjDKtRvYh08JaaTtRIRyF2O8x
5o6RMy4ilt3AySmtWGLE1T/b5OR/kftS6sPDq6V/iLkpdXaXn559XFNKu961oTZQ
hk0gxh1VkjBszRX3uo9neH7l7sOom/z3VPPdJJk50p3mCyk3kVlU2qBNUqpy4smg
2DPEXBj2NUOmqtoT7fBn1tq6iDZ3JgJwq1Tw4M4l4PZlA2PQFcLB+KMbR5WmjypG
GgZlmPQdM1wj81lPoDdgKzerXra6WOlvP1k6R9tGuT7mOpkvX0yk+hl76ZJNpDil
KnjvGA4KUnzQZuoSevN4PuVtiJwfE0ROo+F8rc0smk6FirKnVHLbexWUsmV/ae6q
GhRK89cTd5eAulhks/VhKifKezKcQw2vqn1dbRoIR+DwEPVx75hbaSNADgIQIrFh
sIUsNP/T2YeHuYnVy1tWV4GLjExaZhuy//gxBEjOWkjS2QLLniu4NuHG3O/fyUR+
3L0HS2e0O55bgYoi7++Ry8/6cYjYsIJ3yN+ack/BesXJh7L/Ny8ReYd+dhfDu7p5
hKP4zkkLD/RevVC0w4nZkbVkrCmJaS8jq9jBtzmvvQyk6L2x8Ya+SE6a+F+8+3jj
g0IJMZZOj4Iz7EZi7i8gWPo1PNC/jgyz/8XH2EIBIc/HTEIF98oZY1A10lQqd7Yz
NmgoSU2Vi/QVL2w1nkzTOzJj+uX2xbDisFHD4mJ5W9TaOiG8zPQt7VEwGqvutqb/
asV4GSjQrjer3xBgSnCtmM8bbDOI72fL22cLmPJzBNdyh+/roeB5lmmoT+Rj43KQ
lci7ObkimWlAvWbJ6p5g7gtYD0ure6s7glGfL0a9LCSe2h+k1naf4AwC35yETfYc
6cj7PAiE4DFO/92RP0GBEdd08IsOvOuh/cKo2yHbiadNldq5MiIQinexey8m8bgO
KUdq2xpao4y2QfjFmyRlf8O8QfqlbEu0Lkn9c/A+zQgpJkOxn6MypXQt0w5MrmTv
uSm48VGSm5iwjLRWTB2v6RrPkLHtpi6BgIKbbxGCImpPip+5CmrQ8OH+cPbO7thB
fZTW6PHW1nMUsllANFhFGp3MgevqP0b1bRqDUa/Uo3gln/rNu1wMZWK5V+U4twRZ
t7/fHIzHi7To8msa6hU4UDUvCGxME3Rq3ETExygObpltCsUo0nl+UnQ6D6eQrJq5
dv1+2nuWGIpGLrFIGZgCyI5CYlWPhiJNfys2WK5FONQ=
`protect END_PROTECTED
