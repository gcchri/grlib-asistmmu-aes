`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1Pbieb8Pb1TwDZf7oxzgtVtkHO8nMCkTIc50u4oLg8OD4ipXkDERe0zrg6ndTZl
iz7cBR4cyaKLLktSBBDjk+YDQPnCg1Zmu+tpAvwDAMjOE1db/u1W+5WHvyF+yViu
fdkTx1u/J4+9SD/Jah1RDOvIBSh6Nj/bNeE4ZM4rut766HP9CzIaAubXgkhWpthl
umWVNbjs4l73wNGLI5cgy9F0Nw90geRWUe4vTVcKEpCX1EIboc8tqOUPTfwcxR5t
KK+4whSGD87Oipl0SWeE7tecqnjhWKjE/h7Q47rxiIWGwFpFKhbP6Fth1zF838wR
6DAH4xMYFIO+dpwfI82ijtk6PL7rQ1XKDms+d/m6Zd68df/INrJwrvVdRCXQlm5f
+jiTAjMYzfIKyCPzLJXyKz0WpIkDSZggo+BL95Dop4I5odCR8iOCfqiwuYIitCss
RyYETzkin+YpYVbBUzAb16cGiiUeNEWy4c+H+FUTK1h0oI+6d0Uz9ZNUmTQ9Vd7m
LdYwWPByl3PEQWwHqMgwHnUthMP9k92mGqw8yytVJ5Qhp82b4R0lecWv9Xa7uGkT
czX5RYE1E84AJmLmUWEdXZWEwtQFLvEKwFSlK29BF2HOoKOamMh1OMyiEwV5dEpJ
y3V20VQfRg0ag20WoMDvl0pgj5ah6PBl7byi8Q2aFTJxLE1ISMm23co8RxQudrgj
GpZBtl+qm1zUa3F3NsP/2x8IIsee+b1/y2/AULY7EFp2OAHO+vTHRvmNP3eDsgty
jRfWKpts9gxFI1avkyXcStroG1bRcmElERIsmVRpPds+xuHLaQmvB/63H4bHhQXQ
5wkd7gl6JoW1iWv+1UZJHQ==
`protect END_PROTECTED
