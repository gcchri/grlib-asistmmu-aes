`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pOJGsrW8h1uXXZSkOe9eZRm58B8kGfzKNVvulxTxA4YP0feRlyiJRVPiQAOLxiKf
RY6gcncU2KFN9IpNnvZ6PsWbEtIITLSJO2tAPqkX5RlrNRtdZa/NjzU29R3shivd
lEvvlwVLujQV5NmHCz8rwesmsthofc8AFuhNArTEX2Ewa/MElpmOsfbfVZ8G+CfU
9BMcotujnoAaLQswQccWswsrli6KdXQ9qJtnn1ScrvqNzlAjhmKcrKQmAMH4eaT3
GJRTdlHti2y4DLVmvNCPmmKEtMWLyjrqK9Y8gfAm4bO5CZv5rC0FmHCrCc4MB+Zi
sG7FYV1qxFpwgSZVGRuvYGUR/yjNqG8FXUp8npUkT1485FWOmjX+9AddNpfZsAm+
JxY/Nr3BrIh6Gqj3lZ8dDhAUy060UU6TGTSXFngE/ur0ocS6dNpeU8XI9xvIuEmu
SALHwFU14JhljA/5qv4Bs1ARaNXO3lLC8YZ+J1+/oYwCjVy1vlHrL4Jc0s4uKXYO
drOZVRhhZEPS9M+lzDuttResR+2S3tykd79vxy7Yz3Yh0XlPjhi0JUnHt1/lNAVU
xFIP3fc4drBgfMFRA1sWAqjqo/N2FYtuDmbaRtneNmfdvmvRKfy0tfcMl6kanFMH
zGvwWCi7HifNPsfDo1BuRTfO4oqTE8N6to+kk1tOG7dca7NBijZ6FBWe/CtSvzv9
2/RbCEllt94mBNmVDH3IZt/hx44qgp2VjV1SlzyJrzQd9VerZgVBguCGgfyXlApK
lbg7/xqgW9UrIzkdFFk7BnJsnnIrwGLFc7vaEEWRArIWpykpz7YskWvj2Is6GyEN
fLK70pudGgjxhBqk/V4oZ/AAcHzJnHtNno4Hu+FGxO4B+v9HMjWJWEUKQ2MbQBpA
JFm1JHVdIlWtCsNSdGwZPSsinxfQ9PvNCJXvBRs3WMXJuUEbBfTfzXF3xYOXiDqy
`protect END_PROTECTED
