`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VeF74ZOXYJzX7wYJhxqCMvGhplk2b+HTDGc3vGriEGbVyq7/3NvzmEzU8v55tWyM
zZwH0dP1ApnPEWiCpxdTffgFo3OtXo2kbtbBXrZnpCgZ0b7GtkieHJ4VuSPM90rY
5q+UVHGasjnt3RASfUK/E0MpDIL7MvqfES+GrYF0nnAY6NleKqSCSYl8vcn+K25b
LQIwn/f0lnBEttzM0OozbjKhBv3uHuUnr8VZ6pMKb/bRTdGKEtqHgh+L61z2/mEM
JWsofLsZva1XlwcdI0OgXTipWK7V9nzJ5eVzKeWpW4xgzDHttPHwPCTeI+61jBYT
ZVg5m56Ead7tPx3ixXjyrKSuNRte55AMt096Gkc2K7zRhZv1JdBVzRGw4EXGDmTv
F2UyKky8QgdsB1xQjz4M25m6QLSaadViCI+Tep+keUkerT1Q/uaD7nXcn/1+vf64
lhhirJGNdVHAFOjOdlkKg5/OepVmAyTjdwpawzcVULVZ4BxXErKex/vXEs1voKyu
5JW1MhYnPhWegs3Ufi9HeuUYa+ka4sUMeSwpF9aYpAFWe8Mq+x8CB5SU0H9YfTPJ
pHSs0HLJor5PHlm0UyGBEuhhhv8gnXRSMO16voLaoQV7JbXdtKBuU9LE7alj/ghl
YCC5iUunO3eWXJReQNQMKjN460UcOSmlwdzmnYiH/Fzwy5cjy6qpjfJEoxks7g2X
4nze6jE0oV6CaSsWdaILTOyzQlwpj/ptb/sEeJzC8eU=
`protect END_PROTECTED
