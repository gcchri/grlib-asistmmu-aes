`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/zepPNVelR483ZGV+sQCLNSY/q/QY39bz8gPqQTKHo3he4TTX5ryw/pZu4cU4HH
ljlpMpDt/5rmtosc6woXD3qWk/rwHzapImPg3I6SKQZBmY5Kp29keJluNUaneS5O
97JCWBqU3Ka1NxZtf92aWdaq6HEMT/cASjp3+Phb1gXVun9+TWDyxEcTQHUIP/pV
cNoJUDEKDCvEMSiPp8s1aMyoqcgKZnZ93LIZ0COrClzMHnkE2OuLeQD41aJfJVNy
Pu1X87GDyoTGhCI97cGCI7wNycg+nI40xFS7oX+C7U51We9W6Tf+6hjOBUvVt2NJ
v6gO5p2CZzazdV1+t9DoXnRZ393Ec1Pp0JBfrs8AeTwDIGS4yrSEIW0iX3ETrFyK
hbXdsxfjTAYtrA6vAKOREK/bPh8Y+NLCzBhCRf6frFPny1bEQjNBxA1KRo7XQuao
d2yO8PdmBGc4v1YMXFngmc5cuiw21xLBP4VFy6HmgbT84SLPBrlRLvR2yfmk7kVt
`protect END_PROTECTED
