`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOMgE3Imd1o+XGMoqB/JUX2lA6/Odh7JgTkiUUNpWG28hyxVZhSKFWgkxByk2aXx
KBicRvGWdvxRv5DHGqYfc/LQLt4hYPoFuzOhg4L/arHtLO0zSBepNalQOtxSBOH4
qaPhpXm79P2BHhsO6vaR7jfMoQkNq3ZNU4FW1x1Xn3mgRoOB090tVP7OUh9QKDW6
SaedKWTZC4zmd3FkCHatbDk1ubyubgHuRDIVz14BDw85i2g7k7ja49ff/RUMUWZs
ZYX/tuQ6MZXPVlIZCtV8JHamKZdsOlqBqQS/e078KkJt9a7/maooGRVf0coK2l3Q
wfh+2dAoAI4Xa158hQe9enClr3KSsXRWqIg/bCgKA49W9sbTELv7BDwtGjWFwbJJ
1nmPLZe1D7YoZ01IPqZU5oVazq3YfEb2Mf6okti6WSW0HVD6AilaDqlJcOmKeLjQ
6o0Z0KGDoq1Jqh9Buwcr5r78zT4KQgzZ3V6umUKmJZP+0HlLdRn1ikZ+ZLmYQ+4a
BK4Z0I1OvQXgk8fTalfRyyvNE/YN/ceMHHxxrvE6R6qglk35PRzLbawbBCPKbiAg
ZHbPqAS/63ZEX1icidpA6N+dE2q1RVTdiMG9qBnaTWk4uFPmjaVfUTxHbEu8hU6M
z/n5DkhXcpNr2Rj9laldGQgEGZkF1YQb6nVhJ3jLtvdMaDFxV8Wz+o3n/E8Stplu
Rr7LbP7LWzhhwwP11/teRiRBNoO5p8zg016NSx2wxNCrhboAOVr3ZaEwnI0cO1Co
6iQobuwNQnOblpzifRbqH2XTjUkpkkUTUsC7DdYEWa0cl7q+1bA7FFs9EDjTarQh
jIh13pv3Ny4BSCQmMtvqYNE/es13lR0NF3xCk741/KA3kwG81tJgwYvjxgI/xM4n
pdfkoiIDGqzWDwo5wigxaYvO/vwXqtY1gROwJ0dAGdJ+c8130iGNgMQW1+ZQ7oTT
fPS9HgRlGqQ4UmYT8gxffOfPzF2eUrkk2y/QF3upnqeukeRYuwv0S7FqrDET9kof
/bWP1IeyO+RE3E4WsIEiyW4lvx6+VstTm/VRQVc4aw+UpTLDjjSqNJP4atqAvNj4
O1/fRrwCL5EZGCrN0bTl4LpBrCx+g1Y3flHvf2M4WrunD30+G0IUatffJnrdx6Af
hXyYoXhN43pGJ0gHpjgsOuhK2DyPSQlfYTNT+dVk8PduxJxouzY9RqByNjCKIbB3
f6gXUJ4UW/JCjJZN2LsoryE2Tipp6AvZ/nkqdXavTe2Vz+fa1eJQty1svJI+pEzd
HqHT6v5teKQcwraYCD9hxwqTJ+i7GnmdX1DWSS9Ys0XWuF33Sdoz/227LrMg3RQ7
bRH/RqI7JrvlLZ2UYPObBiWkW8ep1ZZdl8dmHOSEbsGVr5VvNSzXCWHLiG7QyrT7
dCmdN/Igty+SUB+/k+2xgsZ4LQ1qKtBA35Tm3VF41nZ8Da2BHOwb95ZsaaQrjzSj
LkAv7o9laO+RiNOhnAy2vA==
`protect END_PROTECTED
