`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQ20h4inlH2sEytCklx4dBVe2/ZY9adyIbuQ1yNEVqAre6MlNqidsvCMPXs6eKZ8
hc7bjiTqB8cmsB75uN0B2PEFUQDao8+8goEFyRuNLgNZXVR4iJD7m/p6g/yfVlJ/
pOSGACgapo1JDPyAl0mGl41P0XTRVj/Y2Y5oizzb8Yw2pvauFyasot+2vcRkUKat
QIvbQpoaBlw+Z0rDErCN1Ud+hRLG0s5dN3XbtlPvPVNvjnHef1CzbJyGysvxWNQ+
5dJzFE1RqwPwBnyCl4RxdyjNEcvIbt2WvICfGPul9VYWS9JenrsqE0aYnvfQiYnj
oJRB5YmqbhNygFAIkTbIYw==
`protect END_PROTECTED
