`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYxxcKNpPcJbHUSgGNLZkUXBU5+reTWzN3HBpW1BGIW39MKeAYe7oB6JX4U00N7o
ldc9Dyh69yQuyGLVkDKE370g00z14FtSrF0kkr6jtMODgvJoDEdpkQBqdSsfRua6
G9IC4e8ZVQJzprOcdd6v3IlEksYtVKCE0O7xcL8aJg7G4/oo4+0fw/lam2zZxpyY
ZFBCZtKToe4yzAHYRirrYJVveiCbi90Ezu1lWbKR4/hBpJq0jpfP2MP8sDBaj9x7
+4usesXS+3M+wdXQvB58nLaV+38WzFWmQbJbSoEczdTDvxJZF+yZU93N1RGB3y7R
Fn8THAGkJqv+THSdM6ahdWzxgzHGjAmZIWALhan+8NxoP+LdCvS/WTlDT4eCUpcJ
VfVRK8KYW4XGcTTwMtC7ipSWwVdd6UO22DXz1p/NnikcC37peiWSVQihxkk7qcm/
CgttElYazn0rgO6iXqkF3s0B3bxa7dyJtDf1/4sPkSBi5sb+2do0534im+S1buqK
/eUGqhgKkqgCw8Yird1iT1hHJDQvFDlM9js0B8B1fq3M2Ye4/M93xAwNCXKvipy0
MgRP7iJvFBNfqYuhjm8cBswu+iBYAas81QRFQz9FobrBpYjUeZPm/8+Qt7fA+gIX
wTFmijRbRUwgzoOKAN7i2aOGy1CiTqQwUG1IzWzeNuS1JP7+3Hhob+5SX1/Z95Zm
v9Mz2gzmqVv3u2Si97o27SG8sLiv9MaZwc8/lzHYNiG8BpcSqiwX8s7lylIfdDus
7KXbgHwMjG8e3wzn/SJgrmumwpd9dIcaTMaiIlNyxy6T8B+eu5axwH4Tx59s2Zv3
g6vstT32BJcA0RFODEYtY97T9SPMsNIHza/63PMhA9IBs0FORjDqb0g/06bzDUYK
zZol6LA6UEdiunOl9EEphuZZRG6wB+0fSTzknkeq5EwN+n7ik7H5LnCVpNcW1wM2
PMtyYCBsLys29Z5QWmahWPosp4QW6KRFYG/ziCV5wXo0rmPWw6BKhZUxDNENi8fA
METl+lkGLa7YnBFhEEMwfCyQZC/LnMP5qf1h5Yt8IUe9NxTA/Pxyw5u6eUBMlxSg
aj8XaKaz68+hcoUNGJIJFqT909SJ2jF4lt+BAb8dH4A8OZCcjlCQjRwujtiDVtl+
mzePmtFIEXuBupUQ2GkM0xdQ4yeapKvxN5jO6TM9zfRFo8i5NCzVM2ILs01WpvnD
V5BOp5iwaB4GqZwxaY+YFIxUBfDob2Pp+24u9+LNY1LhKiyQ5BGMX7e5/b+PUjMZ
WM4OL/cml9o7YWWAkYrG0N50KC4OXW0cNj7Hss2y/jUxlzWp99whVD++vG8YOOK7
NtHRZ+nEPOjlFwiELFdtNbdTXbPTCNiggEAD2CXVDW16q7If0dAC7agwKDnNlDFw
+JVeQa41UAxONjFpjLKtgfJOOAi6gkoszfYEAphBit8uKHWWz+lKfO2vAQ13azxB
pQquP17tN4+Nd62Vg5FX1KFSgLCUrL+3Wa1GPhttdid1dF84HfvMJzs4M5jmO6gm
zxl6tUiQ9IACELUDWiLtHSyyomwfvJzcza0xEq2q/v0GhgTNrxvqT5UdpzdD/bqF
IAYtMcIW1DjGA1coIcwBi724Po38ze4fE5gybiiJmlAWo0/fC/pNklh5OcAoMm73
c6GgRHpW0VBBRI+Mr6cQERN+qHgoafQEygd0DTiv9WIn43uzXVaVwvXgY2i1x5kS
lnXnO9MoPO0xK4tGxVS06btyPjH7g+IZ/DiLeEJ5NCSOWjRUfmuSYR6hhamlYHJ0
fiI/8Gz25Uv9tlftkRHG5l3+np63o0WjnWyvIxwALrDyDwfmGsW+e5gxWPWNZdiT
dJvBxXfSpOioBTF4Yeuvv3MmbtTVYewOkQPKjQ7neokZmn0+D/T25jRqVLzVObV5
9TAiV7Bk3TzCntkucZwAUzlpW16UCGoefYqc15BnL98ezvnj5wzH+kkdop+5Brys
ytVbO+9Ipt/AsWCM1j6QtDRdCskB3IJsMS3lgSKK6kAzvZSs1cpGjdOr8jNuStaE
mLKctyyIU6s0JmKzuZtEfvcO2QPLsqOA+ulUGK7aPu+wOWYHOw3s1yfn6KqVO40W
Ak5fd7lGvVScWsQHh9YxWKe3kHjWPksMOm7t7bk9/OXrLgdXcUNScn37Y4zGo9oC
w8lRCeG80hYwXRbiQknRzDnJjtHX9xH7u453DSSZrnUJBskYxI7BqfWOGbYNxV2o
Wx8ep0gyTAQOGLTXLTy9krBc2Ka1o+rhbjchDF6unxFmOdx+jBNUg1s+V0hKtqHI
1j0fmRore0wWl+zAlSxYCE+/6T6N8BODsh0ZJR6WM3OjfEPuFNpXffhfZ93b2ufI
/UBvCzWQJCXIgfukGwsv3FssUBTF9+KUHbALfe65lCZlL3pAsny4cHe817xyNBDH
qVgHCZ6Lrji/QGiKCqfz58Nd3/KBqTTHkAxVmjw9AJhPqK9YTiMs5rYePL4rlT4e
i7/xO2begWGqcA8Q4meHf6rZVLH6XOMI4h7KQ99aUs4A7rogbBfXBcUhpAKQM6V7
YWm/n+IY1XINwLvd2F92OTxOid9ansR5I+0DGwNbGKJVLRxuxh/Tq77HyLoFtiGF
CXYa7nqDcz2Oq33Vfd+5CzX/0h5zzF7u+sP/6JGXxV8LxO3IIHahm+2YHqEfRHjp
PjYNgKOAhtTbfOh/TWpRwrRxZ5HuCr1MlGRkJGfm+SHR0ZBudTeRMEOPSb2E+GRT
G4D6DT2wzg0oN9Vv5ZBPPwl8VnxiuIyUMEJLSdP73Kbzy9lfwDUk4kiEMcsKW+NH
OdXqIeIKhFjo5X8XKfOy7wWLLXeNzPZYvuaxJeqauhmuYfZUcEQFnB5vEbkkyJae
QcAipdL463C6JeIkPQzchiDu6WWdE0sjJ1GYfmp0TWSy9CGPcw87ZwTGFn3sQG7p
w4PWFVK+7iSm3LZXr1MiGE5RQeHoMM1aKols+mJtLYblNbc96UHyovMxdRbrua5L
RtWReMsDGBPLzhT2fOQmYYtwqOrJ+dAmjETMOnFdMS8TaQuA/6CSAyaYMYuxa7tr
a//psSQSOtDJd2y9uAUmT/nbzmLdKDE885EM9/IOzwYLTRYFAhV6OgS6hX1WV9xq
UI8uQQ37vR58KPc2LU70Pi/TfqNakwW2nO5u3+eqCZDE9lVPQvOTbghKQRkJQwJU
J2q1bY0ApRhLW3wb+B7LGlXNibouU7+/GNA4+TQs2M6+xcOaZN2rA2MjuR25VDiN
+BuoBuoxxv6bz4B4Ji2fym60RFjpi0YL00JxFf9GHCypLOl5BL6WWe6ScGYoY82C
uPg7U9S/TmOREzL8k+OqdHoi0huxWC8f8g2HJFJyD9Q/Pm28jvXahdFWLcXm2UNw
hc82EZccxEJC6AHuZSAx9z8S6F8q4hEFyiPj5WPFENqXFsyd9gjLAu/Vt1mAqrS3
Fy97+eRaoLR2XBPUhGNRGSYjc7Qj4PqHEzQD90Nd/mMyU+rRxvF6C04Hf6segynw
hHmYn0bVmW95KKFnmo/xtVOWTwogLO3x0+y4ZRjeZ45umsJ+6HUpg5skoRc7pNDd
sWH7wJxdFVmOGtBIYPYkXmgZkUsvIo+8VgUGzeJRszdQZDNPTQPPkt8HistAzRBf
WtjeS2Wk2rvbu/fgBLPkNbDCmYP4t8PLS0Hu4rBnwF8ePu+W+UPneS3zyd5wRbCN
MzJzLVDrNShq8wKNJs8KM+8HEeIl0cAWDn9B/mfKXrPl4Eh1ItJ7Ew/tpAiQKQw3
aFxYz+pV01UVPGAo6D2CV9jbMhOecaFhiy61AMP/PU2/Kve0pevlg6QZFytfd5W2
mHvHZz3ViULckRi9MB0Wi1aMVBj6nqrYcC+NHg3E9AkiyDfO7k6RflSMIv0SNCUa
LzfBTlsldcoCqstrlIsvmfOqcB4zgy432CYj3vvD4e6vO5waoMnR0GxZcuD2EZEj
WC8ooDJtjdY6q/sUBRibKdOWRYJGJRcQyqp2XHBBGE2Ib78BE/aQdjLsfixNWvMN
npAIpJatR4SFLN4ZMyiRVHs8tTmjmydbfl3y4HrrhswFsEY6RD6VKipG73ehpTuW
p0x4wDoNy+rbJt7ziS5ZoQig6dHPJk0bJbxFKuu+TfM83mPfXpn/NxDlSzybqUpd
xf27zKG7PCkoNufS0Q63A5hZrOoveV70rNhNvMlrbzg4HrgZ488e9U9bSqivQ/N+
UGDeo2N1J5wmfhfR+ojJqXC1+H/2I/PWBdNl0LWpByMwQRwIZCGhXOTL4yq4rn3W
ssmNXdQSZd9lkH6ZRJalPB4jIia3j+n8yfBf6s7cOvnD0HQRVBz71Lm7JWyej/NI
ZIdF3cU1tFVRHidvPOl8IQG6+8XGSTD9tUBZn5pYdhBxQPpQ0eC5JrU2wsdZaVdO
Opid+hpsSkj7Z0klHmghgpb32EaitCo7YucuJsCBsH4uTNgQM+JKH0D+OO90ak0A
EJMYxyNiayTpcCU39Q5kpnTMckBltdROTyOwCN6D1CRhy1MyH1B3Xcrkpr33KDkP
jexDOQ7CVxy+IX4NKf1GRtcd11OhkeRr8RzmrHNfKtERr9E3DEp+MhhVG6e48DD2
vcBSJqi+KZcI1dSBNXmPXXxRE36xRiKZU9OSXyd6C6k/bT5JFKmw675UdJ7Pp9Oy
NEQOJJDTojTWhzPNfvs6D047uZK69GOPP2oGrQjodf3gLXPscYoykGafT1FCA6C2
uxKXVJSulnGiFHzY79Ab4v8yBA5l8FGv8XBj/DIAfNZtaqX7Xo0/COLRyU0EDOE8
aAOpOKjC/xRqIxRQlkhj0An9yhHayQXg2QFVqhsP26rGL6O1uulVaVFPzUvCjL47
pVeQYzDYmBQEdYJJVpVNbriLXxCX0osuk8jTCgK9rH7DhRssy1ZW2vacI2gdwrdR
JamLGr1HkZlUZAD33EqV3nH6l6u5sybCxSSUM9kZD5QBUPG5NLO6T5P0UMtzSmkV
uZ1YTUSvU/HGLQPibK9jQvYs/V7mD6EuDe57rT1k6UHAcwtQkppAUghsWTsQjlN6
HhrNvHzLjYbu7sbBiOEuWG1ysOyYeeJOQSIdV6QyQMqtod2FhDX01tLAV7kHLK6j
g8ZMO+QKFG5mLOI0ZOHspbS6oPfxBrl4COyw6vrTljPLCqTLm/WzhkTyYG9zea1x
9pq2QCKf4BWYfj1rOTQDzuVqH620+pWk4vMtZDzZJShR8swrScGW5PU2XHPmsuPi
6ZtVnQnNFxcW6ILky9sip+h7qakjKnyIFJwsv210pHz+WqRMkkYmBi5iKfTS6FAp
k0W+lfXjCl++CZGHSo9eVQhpacWv5KC563CVwMYsRmRVEIn0F2W5noSXXhTKOq1D
ld3Pzm4SkwZXYmxQ+U6HiuenCa8YxUdLnxLyDcZnrfPc0gVYA2+Uj38nh5cyZEzQ
1nfV8pg7n6RXwGmxhRyVjl1uz9gmA14OvUh2nC8mW3eXejF7NnLIy4YT9nnV0yLy
GswgdLLAk6tCz6uut053Vz02KiprA3nBxLVCUcW2ehnrzUuuljOiMQWUQzj/2yNi
UDg/LlQboWgHbTO7nJXaEK4RyPTO9VDnCzBVZspCeUP2UnQatJ+dhwR5Y5wgKb45
XLCHU1UU4sWdm3RamrzORT3cDJ4cOk5k+P9x2iRNCbjUP9XMvqFN9H59vDxEZNsa
MpLk1HpJH2KuQAtF/EQU0nfR6Bg9qiKpmJbSJqK4L/X2UZmgz3Yr3m/kWgpADwru
auCNeBA7ds7ByfhXlZCzhVnVEo2qEn5zMwy0u674EkZShOwL7IK9mihfzL3buHbo
OczwUPE3y45aCjES4ADW7+LuxfVgHkDBfRgoPRfZxQnQRwXa9XLGLDDD0P3pjS0U
KGn4UbG0oW8Ija5wMj+592XCnWHQmfzmL1RUH+C5mL9vSrOc+W6p8wfnLHAcWyb6
ytW+6UySd7EbxmvwmYA9b0TtUcQNjaxfBDoSbcJk6Fwsbk2/BBYgarEN93g+3+71
QB3w7BdNOUNb390tnT3HBYhezPbwLsKS/diHLwIzB15A5bAWG2d5g0OopL0P1z6U
ArnIOWLzWs+HQJwaibbUDs0FE4qDaqZnLi3CFQlhC7GhqXmmI4M1Eqv1DifzAN2b
Yp7pK8Le19Jfp/WAxSxv5hjdA4it4Yq0aQXsIpS3VwfgFSpeN5z9fg6Q9J7AzJkK
1fV3kNOAoS7/6T3uwwdOZb8wi2tIUGLomzFYKw9t0vrjSP1Rq9ju79agCTWTkv1Y
hWf1HzUAUdf6aR+2IMZI4N/f0F47GNcY19rYc6iBXrUUCiVe8M5fdKilgR1DX5qA
129ciu2gCV+a6olE7oiuL0NzVue5SYDlvTWaKUJxP1Fc2q1D9/FVtPxgkbOrpaGm
Wb+UVGIOuEyQrIHAZUMK0fyl0moNIICZFGMupXGqEXd2idaECB3anGaogm6n0mKQ
rmgIl/OVWyd6vRDlaG5he7YNYlnWx/13hSCMT05GjCdo9edOwv0zYB3rZCNPTTd2
Zh3Cf0XA5n0tVkfpLNd85KoB0u2lvqR3KNp5FrZ7uSO1mb7yak/eomuwAV0Lhak4
YIrwSALF7nJIJxAMxNeuyb0IeodxBRqEH4zvBxlkcB1y+RRGhurKyTCuj3daZ2Ao
+U5cdi/DMoKuThWNkKIiD2Y4kX1ob+QDWaTa7E+J0FpsfYZ9QmX4FKQRYMWytIKE
tqSQlwhBiKohSVjiBIGORmvziuNDzH1Y3mTVOMsnj1RJ9y5QwLNhoYllvVdzFpne
Ma4n7Uev0+DlYmQ/FjIbgwwYyW8hUqVEAFaghz7LAG/qkHGT5+meW6zycm2nN5RW
LxEj3OZ+s8uih8a4BmSUTNXlqJUzfs+sM3m7u4oNtPZcoatOFsWigzQlL5Uy38Zc
T2o78FiDIbfc0Q7I+F9XZotm/t9uPE89BT3V7I5ZCGrswfFnUnb2ZWwvSu7JCiWv
Me8l+JJmjriibUKMuZDq5butIJlhpF8yUZDrhl9P/ZNmHILwC8bcbR9GKcfYvwgn
tMwMTRsF4bD1rOD3xKyPXbEs9v/35Gi8ZjD9OlThqEZ9kRVBU0dRPBh5oIUfaTwG
PeiaSK3x4ke3majxgHRqlpiC913K18ORygRft27cgh/s1AlFIiQgvywajb2sKXyV
Am7scr0IaDPtUPcmVv/xFP0EPJGPB47Qq+qi+78K/T8N5IPrV2s19Rs7xJeKZFUR
XALkyM622QIAu0wA4aIJgFCLZfiyK6cLCWdxrOR8flibDub5xUxPk4O9uoLi3Xim
nZGrqUSn+mxXTdBV69UJb9NueZYnx8TtZbTLKsI9n87CIXTE2qDqOv5IxFyC8iW4
`protect END_PROTECTED
