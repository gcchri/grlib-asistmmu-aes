`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iF1lAD8x0ADznKSxo3AKPiSF+yIRkUeTjDXQ63YyLBDUdIK/KHekNkXPbwQw2u6P
vHGroE6FqsQdHlAGLmjuHvPAVugbQa+fZoLj+Q3IKMp6cvo95eikCKMjWJIu3s+C
L6hsWE0jtp7XBva6gCrrm97s8rlIKF7W21+p99EG5Bmjpob7WYA7Y9YxLvzKsRFS
DMZbpGjz/382Sp00BC4bYyYSIVO0BvjkhC1bfLSw99oXtsAmDCG5E110+/3VvIxi
9Z39DrhGYgJ+gkpA22H9F7TE4vNk2NqVtmACqgm9wTjp5EtKZozCkKd8ZqnoDq58
JuDtNtD1+bZKBqZUKoz6jPrd1OqlM8N6QAIrg0j79zOEWX/8EYVIKolffUQegs3+
+PnwE8AdE0BX56j6IIj1Bmw1WTXPdzSAho0x8VZcmg46zjnzigtZgMXwLvsXkilz
mTYX4H3idWBOlvswXP5Luy8dnvh9pNVdOgn8OHugMHxNx3erA6OktqIyEFPpKDUm
EmPsa0HIQH/WfKOWAYz8pmkzzbwI9fBNAzRcZZagFzaaBhqKQpkI22okb0SVfvnP
1Kw0rqHgxRHR5FJpbVdirkh+wVh3teCMvMiKpzAaKy8SjDPQbUOgdnH4LNuueqTZ
sz3McxuwWp1/pGPLEG0FZfEFdlo/DorZCFm0Sj+rwmlOcuGKsCXwwKhdE8UcmM5n
Q4sB7+vEYV54ESVigmUpA7d9BTMzji+n00uhRZaBzcVD+7/xgjItbbZz/RYv+D9P
ni8E9hozEQAc5wTQqY6jkNx90uT+8C0uqseifcqBvqb5hFw0skfl7cfK/YWZ41gw
dLLYvHtiEpy7wCZtBi7Wq2jeOtF1gHofXHCU4S1Z62EPbVg5OegL46we4V3NLkH7
m/YULW9545To2mcO29yiuDpFxbT/W9XqL8RRqdSSe4RxjMj9kYy8TK5W9I/+HYeQ
YktKYzw7Mvph/aZ2KYklmMoO7TijRkxSEYk6sEzm07n5LA7KjnV37RTMGIW9Y1Et
cbJv7tkxgFcfTxtOEKHJC+mI/hcoJdZz6m1wyoPtk84e5kTXGNmxPIEgRIFw1hu5
Q2JxhotTatpqEjglCUj+TrDB3xaaNIeI5ZbaRd7TXG49a4o+YoMPvhUGTpABJjbo
PKyflCj4FeRxDoCztaBK395nmPOrNHDguKzaBjEYc1Mc+nlGSzodSF8yxZBKfgHh
NcFWn5pggwd4/ltMSPYJbUaYqRj10smROxlLJ83kvsgm0C4/qZdhI4FC92fSPHby
RG7ad707/VPcsJUXFOyXHMiHMeYqx4gDxJxWJ7O8OKz9fjr1bSpoL5SHOIr3/GyJ
tNmMDyvkLdAfbE4rcMOANQ3sU2NcpRwcfM59WxUGy8/lJdtdu9/+/k8pbRO0rV+R
SwrGeF9Cv8m8oBdfdVFLB0VlGyjxsMhKbqGwwb9rcH3MXSuLIT7LH7n6myX9bcUS
x5F3ZP6vjVLD4jhsRQigUBtjoub3jA9XtpuZKltrPjIt9ZzGzfZ66ZWhl10Nj7kn
q2QiRyE3WtBc7OToBvpn6Gu0EWxdlCCOoffSFIqFN4yr2vLm6Clv22xFIAL1rCyJ
5rNAuI6HErzIZFeg4taLAAKQldsKhy4JDLPlSr6bq1H/dH0UzDn2EANUQUuV4mbx
tqXHvgWXGNc4lF3qmxu4Q8HwXXUZXwhwmprugoaug3l4ewPRQBswnL3l7O5//99j
YyOh/7naITh7QjHQroSDwTekR+vFOSABHlvtecnfSEE5o37ZAyN6v5r7vcOCQLeQ
kk5PZdp8m2Yllbi9X8I6d39g70LFUvEb4umwoMp9rL338kpcq6MpYitZWa3OOnto
UpfHJXplH+FCowdnzXxIDnAMe4v1qVusDf+RZhN/O5YTWnvvEKsV8+jNOHGaUM7Q
ZMfX0B7q32U/xfPmsSzYkQ0Oz7mNSFvVD8Smm1Fa53dpfqNwVRN0iKRTNAPKIRzY
6J3gp2sFF8x2OcpoL/X6zKB6yr0Wj2vAs0MZzIYLDeDWAC/L8FeAsFv6sWE7px9O
hMqwsodlu6PsxUMOjYL3OYJCjPjdpeCWcUkODp+alrxZwZ10VyufI8bYIjS5dBSI
+9S2o1hysUXaVwCdTW3d3CkQ4unPOxOW7nMyrGXoy7f3F23IfRtnpb2wve/hVsVH
wh5YBEsIrPvERjEBOs4N/iLqSmVf+sYy0PdzeT8gCThJBITeIO0DdRH7HfrBin/E
SzLs4P/3hHkc8TjXQiMD1Tzmb6u4CrfnvRhP7D85kkS6edg3JWXvFo9P0VFsZEiH
SNzDWKGY+Yf3h/AcmLB1cN/BiOz7LseABC9iAa/uiQe75icvgOGt2qRLKmtXu9/K
/oM0pru3wjX7mUdNTaMeVUQ8WH0HfP/1WLB2v4u4Rdcrw0oCKh8RSXt90Q5WVTK/
uiOKvBUn9WSD0KDl4/FnLvcFRlZS6K6j6nP2Ox1jILpF9gTH5ZQAHWduQ2h7acho
6EDDZc1azBERCPE+otBt44xIz343CHQkuJByM5Cpo7zGj9nGTB4KKWz+ZLt2rIQK
pWySfSDZTBI9inUxH9NhYTinw011hDm6xtloc+lal8T/irDUdc/k10z9mxbI9hVQ
TzhgskO/M3F5Z+My4sdjTRd1YkOhkQA9wUvRtEvnZwLY13D+F6lnpQTkGQWRgrym
l7RMlLbKgGBceGFJiRVkbBmKn9f9u0zidxLqQxlZlprJeoAQS46A4aPbaDpTt++j
qjXnXNWI9KF5gR6wrhO95MiueurOvUQmnPfYZ+Hf8nh/+OUOuUUEB5aB3OPFdX3z
iPkygdnNB3QQ2W2wRmO1nqPZjtZlcrP0TscRomgi79wUlw/2NTkSDgMy2u0Y/AJl
w9JAHcq2Ai6+uJxktnsij6415SXObxmCqEUEJ+v1PRNblNYN0dLBEvvufH7UJZvE
83spsVBjlCpRGo6ISTkHNg==
`protect END_PROTECTED
