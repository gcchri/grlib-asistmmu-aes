`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRxDtyt7vCZ6nNNvMthxP0sBsXkD2uQzz9e7a2jl6HLmUmmmeMDlceiJr0iohoHO
rGQG8D2160Sl9oWb9qGbrUVHPTWnDKxU8C5A1RhttMYFxN+H2ymQ3X/Wek10chZf
7o+tfi5XWR0Crxf/OqpHpfqwJeXz0AeEYulFk4LgSTRTRP+Zkyv8J6F+qvcWRF2t
Z5XDfO9t8XT7ve2zNLQaoFLlDo60lTJzFC6zX+/6WvpuAJDH0Byb9GFDGGx+ARFC
yHCFhweFbmjkcF5fiI5CwZlnWPhJoRlxcFmXRNgA7T7m+pPw3KhmBVcmfxBxz+VB
pR7JBi+4LeveR/gAji8uDuNz/QqMw/onxFqb/tO/CnD2K3UpseYrTU7kUyxTJivu
oUFAQleyfQoSDaMB7zRujoaNrEbp67o+PmgLY5o7YvWJfFO5LzgjKDLKsYgkDzE1
PhlO7ciXZlzP2cuUhwaKSJg7m0ULkyA3XAGUU0NqqawHLCCwzBjUILGNiyzOR5Vo
NXcTBUHEbBWSp6KdmkX/Z2kkO+0O4SNPTiAjFuq2LUXlLu7B03WjyZ6HriWooMYt
wuQk3dAB/NlDZlROsvzV699suF1oRo3tH8/suygGlJBaoR20bzUo49oSWosktQsV
+F/jt//L985PWQLGm318Z6yYb2txddfA/XQNFwRGPXGCL5TVR+KXpN/p7kBv1im8
FPEQOz3lj4EpokK7DriJgWO3im29S/CjImEboKzYJSmFRoQyWCCfMpVclSgUMpqY
c7aPMLD88X+q+Ws+Vcd4Fyw31xhv5AMWr9spMcgjxA/MN9v2h24AWp9efdyepAAb
5dznefTBZIb/ed3NHiW3sFTrn32w9S6tenzMZk9n9Jowjbna0crbFagCLxEgE6z2
LjAMzdwqAVuInl6BmklRHhujIZRfgcPBBH2EU5Fdg0fNysDLNE3fyOgRY5ojBYIL
YftbG0TieipSBIFaOc60AlCCGs0Y+RecQY26/Cq08uLomZSGOFdR8Ge4uZeu8UZ0
tVON1NfwMfqypO/DDPfeC4iucU0GtXd4tm744kY1gKDgVyHJIyhcvUV9apmoXj4c
cQubl+bsRCioIPlxSDaheIixQpKvVvTi8aXhT6My1JKdcjJICEt+hVNoBjh+X8fI
s/QDfrIjjts9KMoLIy+tOfIagd5C9oL6StUMjBVlK+E0YeQkWT1J+Iarphov8sW7
I5d3GkHcQTryHzVtlEHnxPOuraexeQMuMHHRA0hufWOSzcxPkBAWQYFO1SPD2RPB
OA6eccf8cKFodh3pJ8MkA0wquIv10qVD7WcbVoSRrgu8XTGB7x1jxuEriKQPt8Mg
rvippXYOMZLoE/pFDR4dyrj3QjcRIXZNv61zTp7R35XAT1IVxpHNrfl8PZEl9UXM
tgswYPGJM3/vP4qizbwwTnvAe/3d1/hzu8xzvcNSdLHj2m2x2Xpl5dYceahRkufc
xP8k6ifwkC2Tt0Cxo4Mmsd18nWBgE7OoVFZ+kd9RMqtFG0r623aPODOeyBm6byUb
eTS9PG7GJhA4RpDN428P76mmNuBNhVK8Y9tpm3RClRLZZfU5OwrbYKUC/lYCKNTl
mSKkFZdX5+S3FAFwTzIQrQrp1RN8BdcS+J3xlYm1KPAFgRbQXoWfqMdWkWITlLqh
ewlPLpEw6UhK8Q6kDLQl0ZjRSNxrnEXrkS/2cvwEvJiJT1L3bh4gr7/6lBAxFC5a
kHDxshyveVIlzJXdwm9klfel6f8SL1Td2IK3On9ygcjBXsolXaM87/EYpNl/HjNA
nbOxBjcwpo/bw0rwvCyV9KpX5VujyR6pLBZA2aBCPub8GEcz9aEFZULms0xVzhM3
rS+cAgcUKoJR+Bn5h17B2elpRZdkHJrQ+0ofbZrmejjdMtHiXdAflhnngV+ugbO9
5yZ0dDXNVmO3fmbnDZWSgRmNe5RZMgL4WgT4QQeg+VkUIfTmJ8TmiAVuGxArCrMK
X0bRbXgiMnf1zsNZgf7q1VLob3tesCOpsBKUTSvM2/o=
`protect END_PROTECTED
