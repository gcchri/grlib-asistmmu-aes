`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTOIUbDQT66/zniRu5O9E0cQmjQPX6K+RqIcW5IvBwLHosSopcba1JJQc3tv+lJA
z7IR1ZFY5jm357WbDECfxu2py5yFYaikfvL4T4MlbVuIcRt66h8PKEoFEp5SqRUw
gAKFR8DbIkQiipgpQfjOiArB31sctSjS3PiswOFZvW36QQTK5LSB4s2214YvELJb
9hoMUUglrjCziJiNSLu6Fr6x4Wl+LnUuxnrc8C9LujfAJhQEfUUHUKwWWwm7Hn0M
SQUAM1Us48rT94d7VuWSQW7BLMoyKEgHPRmcBr1+2KVwlAhqfhuWP2Z4CcUNl/w0
O5gLB7iW1JIraFvziNwQI12j8X1a5e8DoeqcW9EQFCK4ucDPl0l/fU5dVdpYIBzU
/59w1sfRhb3006BMd/aUJfdoG1AgsWsZsgKZbQiYgM2PP6yFlLFW5puA+lom6lDe
GIwcmVYi73HYlsrv+06aDvB52Bxr+zCQW6uK1U5xM5pMg0oZbSCeLgs9WUyWPhPn
rFdeQ3L2uPlSYOFXrvlKledq5k8kyqZAllMPsVvQ4bT2ns9aWOYpoQ6LD+/pLR6n
l2Kyaq9NKUuX86ed/4o9QsXYRM701zZ+IIkcvcNsmAM=
`protect END_PROTECTED
