`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cF4D0dV/OtcZCA/U9YO3C/zhRY0zk61PrESqmqoCfjeDixxskE7TMW9YZwD3Yq/O
1ceYOdKviGTvXtnVZ3+rUWT7d7n8W97G0Cnvh9zuZPjdTaN9yNTSN9QC/J4Zg2VO
rrLDCamGejm09jifK3BbgF9bt4lJXiVDrzj7Bihem6mKRpU5hycobE/avNFYUdl9
ME6tnR03BJy22oM/sZYKWcyyw/Q6303xE3x0tz2Ii/J5rNgq4njdOhaPl+qU9/GE
FSO1orbpSqgZJGV2/oygx3lws4wXxYfed68YJGshPhHuCtLWmwxFFdHy8s1xkJRS
e7mJMv8z7yMtHkBwHNIqq+GLfPEooHhUL5PzVF90gsYzVVQm5WnV6mgo8Oa6VoeK
6ZUwD5MgdjXbF3IPSIbHw7PQlGOxWR0lsgcfVKFZTIjSjyzB7RLZUi/J5pjPy/Qs
TIprJYehINoDBCGX7bd9wPWBFJNfttfLdVQXje8GoDu8nj9nyQTrotrXME9oblVU
`protect END_PROTECTED
