`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5xaRXic5/1CtvhRpTlz3nFRtZWjNwedAarg8LG4Uzq9TGg04JUUMtSolUKNgan2k
wTWD/f3c7c8yPR0/BKPbkPthJw0bbGsmTkQo1MdlYxJx0H9GXy8Wjge436Ml9KTV
N/eKN8qaUMFfQWu6SBHuxoGIcvDvzrnjxQF+BTGztl6amggoMYDu2l1hK5WFZRCd
zrhVOE7kF2Dy07luEcm3PgMT4dR0/p4ZgMqLWf4inZXDQ2hrCdVxFV87QAdAXt/P
dw0y/7Xw6r83WMVmhdpUTywWaQO4eFbUFgNAttBBcHI8Tg0/vm8ZiuQguHt3FXaO
lPNx0eLZFILDilbTOELIDMpv2ATs3MyLeWxUMxSNnFgpC7eZ4n0/t4rzwvtd++dZ
crJKPvdRN3BHrbNHRe0K8N39OqXOAId0Rf8h8I0+miSSPf6vgW/jqBTAOez/5Iev
3s/effK1zCg4Sn1yqEq+J9hzLe2fxk9xcdlsYEjYHHxjzTH/mrV4da6KnFluggO2
kqHxhPgsL0suiFIopbadmuF//LdQnlCiQLn6h+LyO/9yidpZ/FqseWNMGWYwI6ao
etDMabmSwpV8vjgq9t2ky6hmIAXRJ0KcuSKTonBVc0rUcAVnll5lb3HURkPWwmGA
ldJBWO/4TMO2yuK7JrEj+guLfNxwKcxQPsG/kp3x9sKy9xhInfC7Ks5j7XWYA3Iy
nKN7aJEa40NYv1LhmV9/6g==
`protect END_PROTECTED
