`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3jw9ARl7j/UHVNorZnPsepPY73gl/rBpSu/GBkK1fT38F8CN0jaDPro/ngXv8/Kj
ie2K7ES88aZ3CFhqV0T3Yo+FBkTrq6N1KKRczwPVrz+0F/4wxBxlBMXQ/YbPItHI
GIz5/jMV9TSdjoaGbW9XsWCgdZaZteVhTMIYzPqsQH6kcUT+u5v9MYhAe92gBuQQ
TlgR0FJ+xTjdmQntwc3yZobh7V0cPd80opG7xIC24mEZrKgBUGJXfJolZB7ZGdkO
D4Bu5S254/xCy2/8DFAo2koDKtR67TXa/b2UbXxWN6c1Qc4UvzXG2ZnkPgZPjUdx
E4fH3vAgveeaQM4fBdcg/eC/D372LjGY7rksQ4PrtVE3Abf0HMoa2/fsxVXLDHPb
/wuDfSdMkyIbkxJUZW0k2IwjTPPgmAOo/nuFPmpM6zNhlrbK8tgiRwF2D2zvl61V
7EgJhWN/Ki6pTDuFfA3b/x4j40KzqQoi62tMNZRpAZnyjRNp1cwwb9gGKGlyoX5C
NKdbrtbW2GY9Czim8fjKhv+W1Y4D84VVCT2xLxVvrRphOAuEUe/o0fgFLfcFEhZY
/e84+UMf1R2RBN1+6bzR9ERA9qpOzSOkTrytgyvA28TEw2LDISaFobbgcxZHVzFt
EdFAOIV07BOQtbeID+lK2w==
`protect END_PROTECTED
