`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxIwnsDgKABN7u29H2R62+PuP07GiFvyTbfU03iDTY7HYynG/vuT+6HlBzMC0PBh
NIvwkJT7gpkw5xMd47BrYEiVGg1Ollt/1j9zzdqzzb/Xkpcqxc34vsYucohaq/Wq
G2T+rcTawVAATPPYilWURMN3IGQQYQVo/0/Ns+nxMZed4InLyt4TJ8dHblkUk6Rw
ggAuDwoH6okFZEjY1719a97Ay4WSAeyh2hoJCoYIgvnVU69FSKKgRM4huOspm9z3
BQoBb6mxNPf0iZHu2U/YIEnNv5nW3DNr/6h2b42SJbp5P4VQN1k6AWejafJ+1dK0
bEk+GN9jMlmDdepiK1UVC3kL2uiCPCjKIc1f71Cwmt/RMO3WXF2bfaa47ABMgg5R
zfMei7RWa2ONpUy1zpsWd62nLfw48Eeu8xPNRPkbulMT++PGhHKwkTwWl1WPccDJ
ml/eFf560/S7Shcz3rK7mOTXFf3TUUeS+IG4lVXFFIL/D61kf8suHSIg9Bj8lGzI
R/dbv2OHzOOsQunhHvdSwhB0PzR68v0ipVLNq7xkiKXJ5Jn2VKUEkpJj3qnpKHh/
kk5iDyCQ8NbwQi/AToNo90q9/fenJFWr0uNH+tO4gNEhL+ab4fpT7HITnW0/tfHh
yc9q1wBZAHoDEVvlTkxlwwXKos7ytSqXfbVqqTv6vUlCZViBhguWeZOp1KjHXqWO
66weVW2kZQPEJsYO3l3rmgmYTrmfWq0nR8bPie+lNhk3bcBXNccd4H7qh9OfsKe/
w4QZhgdgbijpMVnRpJj0CpeNHjnxcMHrZldt5YfDRV+yc1f9BHThD+uiyoBBGDVB
IcTl49sLGmuC4vMizb8GOYl338o+qHfJg9qvTYNWkPw5buQzxlFjEPzYyaO1yld5
w759K3Q0HCaH4ps5CVsgexHOjQuGhv43N8zk0OlctcsJtBbPKwoFc4l31OTFjMvt
Lqpjn+CiieohUvRYRvTjK5EfQEJcsVlmvn5uubNUgq2R+Vqx623ulFxmEXJbjXni
rhkQOUL80zp6AlaaSeHJ7kQUKdujUW6R2T/kOrrW4LuiWawut73W0/nFP3GcZ16G
kSct3Ga6eWyl6GepxldPpFAtI/a50B4O6eAzSuZoGLA3AY0EKmBYFSUPYwL1eVu7
jrIIhqfrMy5MAHXtvoMvZncLl9iTt+Ec4ngdHnjfL8SuTdjpZ7xa3OZrc1Kf9ePG
+PhnZkiH9dr7fS1pFM6U0WAphLppdfrPK8TtItI1FNftonhcauBdH1DdYduNu4Lo
RRuGHVl+if9bFXC7wt/agQaC1Gj9zOYFi1aW1LMDOIZAmHn8exqMzieSkcXmnbRv
MOEW1awdDCY2oRUi8Psba7WFBGEnZrWbGJp3Y1eTTTC/Dw9TUuYn/QZkV7vp/xK4
WzIgiNwkiSyDuqUmtVa9cmwu75I7BtSlMZYYFd8aLgF+EbzPdusSXCNhZ2UVXeoP
QZl16d1eoNlZNfueT98ntZtw+wtdGwc42iSkLY/gpVMrJYZ+uLnyZ5NYbvtyUcA9
IahxVhgXEVgbAWPMXvJogI9ywgqiQi5aY3vs8RYm9p9+fR+vSOiU8YiNdBpKhpCo
EprTXXJJuYFUN3eRyrVs0u01DsNZtAS7ex56kNaPXW67nkBnP/8XYQSMKciYQNiZ
vmnj+GznQrY9/NGlcnZOXOI2KW38W+MEX5k0dVf29azHQCrui2fYKRbJBE52ISY5
ecNwlHdE51uHdC4F7r3rdtTxE7+MocH+GUHEitOLBtY=
`protect END_PROTECTED
