`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JhncYToZghFD4Bv/GpWjhApbS0tDQotm9HefV8CJGqHlZtNjlSLN7088T33hS6Hw
tYGv2lGf6WW0ABUQXL1tki5Ot2qEoQHCNFlHPNc/yAv/IryM71dQhaDFLujaHunL
DKcaD001JjZwTTGsezpctZbSgEaL0ef53jr6wxJT9FJgrqsHv3l2N9mOlvHyEqen
wrTvj4JelPkLgdqzJpuyqDASfxZBSKOGRSP4XdsdQzjrGshM5SLQaNadz+Z2XEiX
YrjfO5+91LGYMXhffFkJtfW6FjZeQI+49yP2zJBOgQ4YB59Krz6Gg5DY4Ahd115b
z1iLJ/28BH2K/v+gwwfMJAwaWlmG+2MMlrObhrzuyY09tn23us4x1XKs2VV3jWkm
mA7rPlc7q/e0/FD6hyd8jrb/fSvdj2y5wgBFFF+Ih3Zpp6i9z+ssIpfvcbOlxv9Q
T+YtySmWGNSU9uP38z33n8jPxGnsKo099bczxFiRiy67uAnyJe12RNpx1pX0YkW2
ldTNhpfGsu1GlPL2rjVq5dWfBxKy25RYe+L/yWMvONQzdFvSkVpXkhS69oRkT+Wl
EaSeB+YgPed9VErrGesAqxVmeGbFQFX6ON5Jze2PivRkEZHk7qqwhXlj7HgdwBZ6
Zfu5b16s8RoYdfFV8B1SPT6cAIEoOMriSbswstCx/jZonPVkNd9EePU1bEpPcyRZ
nGK9lI76xOP40R4y061RRu8IFC4fpCqQhNwYjaQ5G7z8SBV78WPfzu8VhlXjM+yY
F+tHDFhJQVaLf4lCddEyG9uoc1VcjoWT3qpDCfXUcJIhaVCB1XDNwt0XiXwgYICL
0eFdFFCwtHZSD34L5P1UJsAUnhK8jxm5kfnJD6WF3WHDwuNWIrEw/upEI7IiCxTr
DYn+5rovfk97iAQZnglF+lXyPdCQWd7A9HDMrPp7+j2WzQ1JHrUcWJBFu2jw/rLH
Q/wn5ZmiZ/s6SZCyCjFJ0S0t0rErCBeh/XlDXRWjw7otHrvo3uwa8n2g8Dedlsjf
HLK1KJAtJAnj60UjopCRgSuAaoCidesp5IS4GmceLYpBwGuB3xPv1wSIN6izLTqg
mkz7+R8CANH9Jukl8rTdpAQr80NYEN715/j+PT61g9YfuRPsFf1cMWsj8r6ES63U
XKjKytM4XRPtIBRkRvq1OgXgUkBzR8xsFF6J6vDrzr5GFs40BKMg6fkKehvpkNQG
iwFTQNmjUulmoNkIL+tN4T/2GJEGGjpDCAcpa1TfBu2U7Bn7qdHmlg/freBolD7P
rLEa29lbXY/n9vsO0gj7BXZYKkGWpCRc9+f0OEWaxJIjGrx/saLo5Wc2C9nKIrKQ
fVunvhsUZeGKQukeDKsqP12XVgn4ISx/pVQUT4WkRuQ5dkZcGrlWxcwwP/4VMvdw
ezpGJ7hyTeAVmgofsgPO5NLcp43/ADZsoRwfriQJViezqZ5TcSqBLdXsoG49e1YW
oyGvkh96aYN43l6gNqCH0azXXsnUgLnhDIBMZHYsGkrJIPdSEkzr0hYSZz0HzUTQ
16fN/XlFJur47RyLxy0xuswA7uglkCmet3gpcBYQItUFLKbeJUZ02vmuetjVdmb/
QsA0N/Bg6cxxAY4LpzY62opgqBxWM5AhAv4f8joSLEPSdm0tQ4HRl2bfkyVBR57W
I2ifujDF10EJa3HTc3utlkfhSIkBfy5RGEGE48SBgj9wXY3r+3fyVHlqxUpsZHqq
GJXThEexPuqjLwVY3v2nVyBGrqq7dYOFGQ0YGAmoWLkl55fYbZUcXGr4hjpYoGpU
u/Siw1v2ek6Bu+c3xQwCtWgz9s5Vt8KUDvwSwlS6vgNJuMgSdT3S8ICoPFT3ABzZ
rrckLf7GUsTKrc2XxoE6YUgsTW2k/ILqTBHc4Xfbb1+EjYgwZXfzJTI166fwjwio
G2WgZqFSYLgm2uKrwLqKHBRgVVLT86mR06eDymvgpCGsviXQVJCrTGw9LDv9rNy3
pSaltGB1dW/yKaUycGn2K41Yf0c7nIzIpNZh8AWH1tuFsSSq4RN0dUxf6c+gmsnD
ByfJc41pjr1epU4zHQAeGo5S3qqKWrwDONQ1XJyDACKuy5F8VTtqHs34D08OMRVn
hlJPzVFx6RKB5bs+J2KBXCsX6nwgJgsvnd7leh8rUIfQcsOmQXiHxtVU8/yb+wIJ
K+iGRRNGReiEC6v8dItmCgFf5ZrC2zKVJ6mGwDUxiy+iEocbg9fpbSv7RNRuzvKT
YfPT8ETGIlr4oaXs2h6RfdrmFub0680mZAY0fdv8R1TN9SgoHLTIsY2vV+A8I1Ag
XKq7Y4pRt5Er/MEyCImWa7VDtfkTJYZ552YNZgq0EfonmvWjxfFe1CQBXIvUaUi8
gDvUkOvmL2y74Y3uIaNYD3eJFRAdLcHpgzz7Bv3W7/TXKsk4V8ItHXosqLcDzAg4
L9ljpWzd0yQaAbR3gifajX/SsFs9lKUSSN7XYMGuD5euO/hVIkFzCQhIcVbzmSr0
6SDlQrwsD22puqYrXEaqGiFO6wUmmnKQfv6GLCUOshRMQUbg52iEBB2jXkVP6hJi
fFkD6n/HUjn+JnUBjsNkofExto3DSMHamfjcj+RhJsjnQD5Ls1/MGhVuDSFIgbmN
cfdl8XAXDjoxEKMcx0SR995QOYsU1oy/bNTny9UaGb5R5DYkClKJ9ZMX1QTySp/R
REG1JZQdeQNfNhI8RoW65tHb+d40zyIrxZSxt7gySfWUKfL9zvOg4W+yih0gKf3e
/y/fMm9fYsCXzg73p/vOVD5TEYswPEPw42sbeJJR0UV33ZuxAi/D/8Pfzqs2bBlV
0psgDxPsKPYnlxWsxs3ZzzMarJ8EiTaTTxFy4pXTP7HU9fhndlxxC3LTGbfF2oqs
lX/0/tSTl/uNbABT9yx68xAl7n9sbi4bgRkV12JcxgK/hvRSywAoh3YSSuwGNv2F
fR4ibd/io8E22SeIUJKuha8VQQcz8WgdO0/IW2/OtLTqTQLDkFH8iaXs+fmtCTQu
xKhl0irsGBYRXKlVikz2BQjWRBd4x7erZ1sxEB7htsnQ9fNfy/BUDuoxeT5E/JqV
MThZEnsUyhwQ/UR9wE91NGJO6V9QBnp2PSeQT4mPSP99U558RAjiJ5oWm4PFi2D7
b69fodyvQ8owmqcTHjnN4nT/vAHIRmPXWgNxxXMnVEmc7W8DdXotZJwWt47iUgsb
xBCSuGp6VwX3PoQlHAEoNOhTY0Ghmu4i+r7ar0dcc6OCNtWjuGoV2KCavZicPWoc
N+Z158u119eX8vQAzpYsaIiogPyyovOON6TdgNJrwXyYGFXZg+Lb6V6Zy6F2Argv
r3iMS6DuDsU5suJz9kaahtgUmbe+zvLzv5+gfGWASk2q7QLHHNrYj+Ua/vRMnTxa
XkdJQGYnkyaCYO6tgAckdJegEeWbOSiXhJCubDtNlC3eCzpPGkRgSl2ROy7JGdp/
VS2mMI+Jz7xk/uJgiehcGyi3jZsG75m4Q6VRxMn7gsazc0qNen6nZUDLmForHSEX
sMA3AEVDEJg4eC5udSF0g+h6qST1WQbVPbO61snlmRhHFQ+H4gbyElBjHB8TmLbH
tA35i3mGoz3fXS+T0uzLQA==
`protect END_PROTECTED
