`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2xLXQcPlLulfY2MOYun5YW/GrMvS37w/2RZfLDYyqGiq+bB3xQ2NnERywyQMxNHZ
tGSAqwlyK5cFszX6ovM5jXhuOjH8uy4cqRvpf89it45/dsLjR1+4AUKr9fVLovUP
kX4x+rhtqwKMa6YdQp4e+PWeHuJ5IB+sLECkzLxli0xyI8LcKT1BpsMes1bF+CRu
WN8fVI+KFzgxZdS997TCzTmFXByCprI+UbxYJJiSMFc73G399DosFtrzL8WATsim
FdpyhWS6T7fNhhe8CBBoedzRaYU9Mk+2Kztoc1G+acxOULTzT9+HowCeO6TujqP2
Lq8OQQsAnY3h9NxEthRUd0Fw6OL4wAO+UI+2BbGXWsEphuCrF4uUS0vgK31SB43u
TmEaZGre4MpY+VQeCdguIzK8j6TqXcMqC5114I22n1eZOEq57V0HXFOEXuEqSGrF
HBtBU8VfQk+R44b8JOTTfS5us2DjsIOhzmdeF6/tI5exuL3zqJzIABm0YKEBeXar
f/fEXcb21PhZf2fVRtZ6crHEXSzu5jKd3zIujte5XST6IVZgCl4Qt4Wi6n3rbrXK
AWioWtz8XSBcxxlLttk6NiHMxu3Eb7Zh/drQVrSbq5LK58rbOFYg2rQBdHwIyz/B
E16Uzqunq0VDVmVI5wQLDY/K0F6KtqulDXYGQTrADPdhdsenWBD267xVLeC+OBVU
shaEKm7atrWzyTSKF5osmTjbYmLpQt4snmeriG+pdk9K1j7GNz5DmWZBF4TDP/Bv
YzfxZdA9pbfDOtR51YzS1r5KmxM2nYEv8WR7d5UBrF9hTkm+fFWiBd96CSmExSw2
6YA+HPudnN1iO55/sHTJjeh/U8brkRew/3iSoZPSfX70JSdF4tWBMt2i2/sajIgE
fhcTeW0FC1Uu3MrDNVL4BdIfy573od+D/3AGLGXIQw0=
`protect END_PROTECTED
