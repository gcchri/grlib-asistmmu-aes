`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zZh3IYHm2t06AnC8PQeV4gL2PbRsISgqdVFJ/hNwtsZj7vYceYRV50TfkQcRcY7
clXBi5Hp3OyUUaiFDJkUtFaZlCr0LDTMDP9eHhAtLw2CkaPnjZv7TFEpMvtyt6ks
k6Y81Q7UYfSqPX3FoCmUJLX09ogbC9KBg9BZ1/6Be1GHg+xB+8sr4b7qZyctolg/
kdAOH2zzcNwm8YTgYerPVviByZ+1jqh5+t6wtQNyaUlXVz9I23frS1k2Iw4BFal5
QcbXbxJmKHjokw5FQaQsNOK8idMnts3P3rX9cu2TC1KVmjltlXDIajJ2Et/HMZSV
ZKXc6FFr/d4MWzlagulfKMDvhDJqYNnJ2IihFRyuLjdOzFUEyfa2Z9wmvM4Fg7qt
KM+/byf4Q19zJzHsJA/su9looBYpYvEnpGRYVEpirgt8cxgIuR0CwRImjL4V1DL0
t5oOl75NNyHnNSqk7CMysq0A0HEJQQngZFVKu5bx7xjA1AEAO1ESJySNrYXpiWY8
OvI/U09e9bFkQA8iGcwHxNZ3Si8nChDbZPbunyNvKv56cMFL+IPyFdCpWExNLfMx
MhCie2Ik4mT3fE0jYCRm1w==
`protect END_PROTECTED
