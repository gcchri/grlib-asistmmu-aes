`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZjNGZw96MlydMv/qswI6jS8/VsUmQczaDI5jukrJj91DIjJFJbAFELpcUQvcYyL
fwnfRKFqq/v4uFrjYqReBuaGnAMGW35Z6ybGpwbMrpxuXmX1Im84iLSyYCOz7zSQ
If/+WXw4gUCRe58rdCV1whU5yIY9f5ZA3JbOR+n9Fr/ZxY5WpUkHl//X1psilqxt
vBkOyA8V2UVH5inNl6D936YRg4p+lgT9kgFuKousBkjc54/v4OU7nHjL8e8e4mJy
5+MqWBoRbWLpUd6nBwFtz88m3UDPUfeqZWgGmmBqTcghFWjnYDMmUjlKKJ9Gzvyy
ugQH9X4h/KFrEC13AplopAwQpvxRkVm+CXQWj+tqiTkEh2CRxIRLRbal1LU6QFLv
`protect END_PROTECTED
