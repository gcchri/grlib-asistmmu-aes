`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EuK+LevJBw0U9puCmiATCwWsRhA/mFB2L/n7mkZ+PK79p95k+Ga/zvz5TDIPwGE
XJFe1AJyh9uWKCTAcyr7maSbb9laxSGWjsy8M+3AxIwhkTgbKJCRYFnkw0Rg1Ut6
R9BSk8RncIjvMKf42u7mNCEXxou8wTiGrpI8ULfDSG37K9EkVPCeQy/Wvn4Cz429
A7rc0oswv3HuEbwKrBiHo3dlhvI6P+NW/kdAUxfLhDueoJX2HH9a9w1mQ0zntqLv
aDS6sTeJrIaqf/faGfifiEYn//rz3dUUogqa9dhRHJD7Z/ph6p3zN160b58BjoPq
lMaE017EFZg/tcz5uRcrIUJJ63Bd0GysXRcKOEdZAAv+tYRBQAvbRAoHyBk02ENq
b1RhdbXPfUSHarzxAJDbf9ELgAMi4H3d77QCTxpaWY0TNnwhsfGIklrOIh8mDvQ5
zc/1IcHgppsqZ/R3qjUhAE0gpHJo6T+CSl9/06mkVLBEdLWk4xywjHy5nAZj+QNe
haewIsz2vE03nvMhJfNJqaUzaMQ5FzLVjOHVm8waa0w=
`protect END_PROTECTED
