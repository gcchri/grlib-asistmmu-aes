`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QBpsgZbGbAb7BFWsfQWhPwL8R3yrLeXUX+52cdSQxLOHxlG3RVfDk2oKduzJFz2o
YoMswx373+WAsPbUgCPLpOhivJP9H0B8Mrdckjfq5IZNRaf8krEHKqrAbIfoN/9l
cHfjKI4VQ9NlJu6h43Js5FN9xka1Bnr+e9mCOlGdQPIB/pXKDtXLOcNJi8mzmSNC
KwVktsDPc5g5NWvKExhUlD726s4YCQWd/wamRy3Q3SCCVlXd9xwvDqDg2H47ljmZ
t2QlOgF1ue/TmL5bf5mAnQU8yyD38g9Ls2uXyTfGEuLlWc4A8MC4JuJ3K+jCg66O
0LcxcqEySC++/2ZTItDd9fsMwNCqS7g6wxUE4BDhFf7JTlR4YmatD/i0NVqZ5VL4
QCEJj106YIP0ayfdCkOz7a/qj4sKJb0tgtIl8oKCIaWp/50wcOCLvTHV/+mE4Drs
CxBDUT8zfgIE3BPgbKUAAuciVyHLFWfrLL0C8iO8IEpSIgJTGdP8IXxOPNv/Bl4D
S9QKZnU6ui7DJFbiCFJUIDCSl8496d9+3hecNMHAdGigL5T9ubTWM+i/6p5L2Xst
`protect END_PROTECTED
